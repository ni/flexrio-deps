`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 16560 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
ZIICkMu+S2rq/yOQyqhpupmJ1IlVmAI52F7eUhB0KOR2LRm1jdRDUrY7mI/ekrRN
hmAjUwZirwa2ZPVtNt3uwzEH+oaqEXsx6GNBNar1dfvMyBltqVQeCgA+5MdjlY/G
2Rkeuxryhe+00Iw7crERIP17zAbVYOnkRhBfkl1aL+dGi0QFDmkBYkEp8ez1Vfha
7nl9mo76555qxFBrbD5bNH38PhQ8Ralb6s9mFv7fTrGXAhPlcj9HgEiiDuO+Mv+d
Tdae+0Z/2k2zDfVeP50m9wk78I51XFX/b3E2wGC7ozN+5lS8kxvhld6QcZVEu0V/
nK5CPUmemuEp0ylC0ey3q678Esc6cC0can4E3mRfFmbuVPIwrxk5hDl6iaNjk+CM
eU9A1aZeqIm1PuXDkaZI+ozWymCmJjw3CRRMZzJgjz/QhkUL7KM/MBsg2R3DNkNY
Z9bzRkcLEVnHJ0R2ktv8NpASZ8iMtgZEXvxMsPPl6l26cJAHg1v2Ye24cAUoFuPx
k1jGUeVlm6JxTDF9Bo8PFMz4tnmAnKhJd23QIL+az3lhoocUJvkfRoPrvz4y9sh6
LG1+zzUD0NGHtnya5tSK+Q8yyaI18IFN2/Zi/ZujchsZyudNoCzaorwovu1GwL37
plTlJkQy4VCRQ+NnuXME1w9ue1moFds/lUDHW2DU6az6Cvq1UJdEN6VnsMNILxnL
M8dOx0YuUH/xW+gz2FyWP4OcujDitpg00iy4IK6M3pkUaaPkSfOCdUcccbs7Trpw
+nvYJ7VkF0hc9p72oRzZcMgtM4A9w+xoS+/84H30ve8lzohoFo4xXiJ165ghi6yq
c5U+ArvUVyeZYfnI1TvElx94R61r2p/Gn+5Pj6FTJMLJmg/9vv0BEimxb9781fyP
zKu1UX9saA1tnuDtjwYROFOiJUEPU7Pqxk6063fgWwxXnkbzclT3HarWSp1oQxac
aUCTVZHdwwCJFgZP00QYqVcywJAesgoUQETngahgiWBfCd3cgKyqmHL7HiqR8QG3
nhR+kX46kYOPAqa443CfNZwvGOeCDNiUhFUkJRPraN/WWXZLqchGoX5OdnZDr9Xz
DRC+fuebyp2aWa9mL1PETV+PQGZNigcofTtu4605aakQAcUWLjEGhS0+1M/qrhYU
YaaXPQAYFVy8IaxOVYSwcWe4j/hu22azAO8PLYnQbtUB2aEWoijdz8XfrTLiwR9c
ilOXj1Bvx4xp+1Rt+PAczpLLDsnrIzpxqIzennjf/ntl4DhkE/eCjPrOcHT/CUzz
Q51FVEj6uLOj9/cZJ7SfeSpu8UPj1E66XcOl2RXjG5ID2cc4DwwLq2XfYMsLIWj7
CRMUsD2+XjnvSSKVYaBrjWr1dBm+2WlNxlxxAT4YZYskGmSEiYvXoac9ZSfxiqrp
rhy2uSmaK9JrIr3w9uVSNG9JrNQqRbzSJSAQTwOQ07jHiwB67bhOYeB/VlwbGaLJ
2KQ+7Lm2ekNfPL79SD9ayR1mBvwQ1B0O2NR3nrHcW9NU+Zg4AtpACbnbFboKWR2T
y4oOLgbouI0vvx5n2Zxx3Kkl02jaunlZn3rBW3UXIAh0oggl2ATB5Q5o23UejBIR
dlSP2GdpqS/WRoa0GCCnRIZWxsNusI9EadV2sVaZlZFeY5YMachJP2/HKd3XU8wP
kt/Uc8tU42fsJaRUZHPxsokhoFfQ+hFB9RF/tW4TDiMPqof8VoMiy0podQYjpcXo
J/SBYU49FJb+EjLM/gDQy/hl20D8E8B/4n0shubq5KXe+HP4Thk2cxILA0NncUza
Gu4SfatcpmCMtxqN2lqJCst00FlaGJ8VHmdHkspEmoQRpL3YDxuzG4uk31Hmx4Cz
dRp2x90QiW+feRoOzyo/F63y0spNjUk3r0acPrZ0kRWLkrBmDSkY1Tn1Mn/gKlO4
kwVB83w/ocHftfqKfui4It9koitWNqbQ1z3aP1Q23vj6ipF87jcruWRFciEVwiCb
ubO1lT8wjPcsxsMIV9RL0EaWpTCfD69lpKc0f9AA9nimI1oxidhP6STK+Pqjbgny
7aaxhoftUt4pYq+BSRLNOVnSxyquccfmfHdzspN6Io99j7oneVAoOdUz9flG1FHA
bguoFwNwfgRL9m0GZv0sMYCYvUVrZLGFjXyW5IeI9FCmvcBnM8WtvzOPMZMnZMoG
FDFVrboLBM5w+gpygDZfBa3iZiwpMNmvBxFlmTQhQ7LcmaGt0KbwubB1CTloqHW5
9+n/fM3Tapqe0yr5G7EZmDMeU1FPeOwcDZIVqDdudGOzd4lns22dHXiuMAw0iHOw
if48Ool5tKO77TwGQFWsWbBVQgSyAEJUP/DBrQPSi/hpKTBzcGsubFVS1OFJrjAI
zvKi3CzbtQq5TOOUmViulJ/rdIcZYbhTS8v3+cfYo8LrD5Q8T6D/XQCI8l9GXVtf
nolY68A13uFeB68Gj9ZlV8DHSJD16UoPRfFpfYrVn8Cr/vL3Pd7DyF8wd4C+tALc
QF7YXzRj531CK1gznqqt57SNDLs/KXhyh9OOA1baXw45F1184s54kjXVE5aH5JHx
xQn7zaqQdCBfexsr29zHj63oeBOiSTyHf9+QuHFjoUOhguZviaVYsg/iXnLxOm14
/6AM6N5g9534axnIFSf7P6C1zNQVg6iqwGALA5WU9CImxjuDweE9Z05QDEjnWGhx
Z+UdulCvfiEJwR4saw8OiFn6Mp6qoOco2MXtZP6hkecBT7CGVL66oTPuH0qc35Nh
9cK0fO3Ni8sRtnI1uCZK926AVOrwag7z4+zZaV7NGDsQX2flspMh5EBNu+ZGYhl/
F4A4jcU/gP3z36/ABlfg80yoEbsuiApQmuC72+4ceuQ5GfO/S4Om5ofOVIQr8J/e
PCgO8N1eMyNOZdUSt1zEOsG+bKyEsmxrLmSPP/FQcADuHfY8Cp/zQZM+MSqxPunn
Bza0JU76CJZVXE/GeUDW+KmpyRMCActaUNYXRZM8r4eX3bJLWbyxCu2Or1wvWSb+
q+jjWbZWUgrzwLgNsumDJ3biLqRw94lbylGi0ntIg8db2o7OXbAonlgkGF6f1h4a
PTjmAL4UYuVYWhcBqQ5StvM22rGK/IKA01lttZtALxcg1JUlYZCrQ4mwDgumhUqu
bJLQZxxHAPCT310PhciE/aYaCCF61UvlNqWWxTzc18zgiFeWBqaBvalfhICNNhfT
IeW7gKxFReAtwhN1BS5mRnFHjw8WLlYLw/0DH/jxy2HsBjN01jwaUvsR0q/HA5Un
hwwuBvLAin/bbqKyOnmTRk05DR9xs/nkWVJBK4Sf/bqNYYME3BajWTrn++kyEaIs
HDw8GqAI0xpspfpOJiRJwNL3EkNnO5Zxy7rV2TAiRKyHoTJH+rBApnekg5CFGiE+
sBvGCgvXQ3jJ5I2nJB+Bzx48wKvEyDM7nQ5qafi8Ir1PhLXTV2dJUxB2r4icjgoP
39ozI2MmfJfn/4R0MIhg5rhBNRrGWaS35jdp2HkRMkr+9igqQJkQISTeV+RaPuK1
liCESkdk1tjvTX3aVtTZLggQl7EMLgnf3TI7PW64NcVKzMxX2qbO/UHF9mf+D1Rx
5V86L62fOa85+4kgTTVCrYmycgHaiV5YNLDMeuaaxj5KIs1bweJ1NYbKMp6dAoAf
TMyft8ff9EiX4oB+9RT5aBiRNZQhtczXKVRCmDl44RtpMUNivIdOkSV54u5RCh/c
Ug0kqmX0sy5+JlrYDRf1Wl4MB9Fi/tHDTGMNwdsULJhAEYWN1r7WRkohPct+VJzg
9ZvPjcM3+BL7ioOsjeZt1v9kCH9CilZC9gzi+TiFBdSHmZ0B+UFqfAV2laIr+JDw
WboXthFDzTlkE1FKnCT79am9vziaYG5zI6Z53k863ZlY+tuyIFTZl2ZmUHfMxlmt
pFCC6fMjdExGu1nlCp/dcgG0bAtX/QIn6//J6myfRqampsMJeLFpURg3HcVehLVU
nhi6mATYTxHHZkJt0ptJWWIcb53x0lVU0raPN2SFZKwj7fXT/AOe7geO9PJzFZBf
t79XpI+FhXemGlZ8l395LWbsurH4u/blX+PKAZh/sf/oU2c8HMytpOpcni8JctbK
haFX0X+DfB+n1Fg5rA2XMCgAnZ9iHCjWk650lxjOGggxiEqbVOmAsQwuhE96eDYQ
CaY88AT5A1b09QiolX9JDlv/CFqP5hBY2KHtPDrbOUwQpdjDOlURMrhAV/fOrFK4
PVZC3htNVbZmpMkEaD9a67ALoU43fWg8/lwUZhfklqmg0aW6qvuVTbSQ1i73QfTu
vP8/Hnve7usUDB+P/WTaQEorUnRczUpXjlfnj5IE8lsrDQ0CEiBrndun1O1IckLX
vmgjtMzRVU5+3hAtFt+IKsz8BJXBJFvt4c3u1elhGkw4kXIr0cMg6BC+pisN4Xs+
jUPxkkT63/avuV12iB1t7Qv5vR/yjOOZNnrfdZ+9L4g5HI56aSR4xOxvHwwG9euO
Yicgmjxz/blJKnhvq7W3mWtkTB/rgrkQuc25Z6Z5e8Xu8e1uzNAbMm+DDv1xMVSI
GQa61/ZBsyedZDyIpNMji7iyMdERHNGxnUT8w89VuqJxM2Q36CP+2QBQJlnTdLs0
7Vjh5ecJkz4g996qmsZpSAGUypfpQ47ICienf0vI5Ro+hX+kNBqkg6vvz47Cqb+j
CorRUhfIJ73jk6pjwCz+uEJ4XV5Sgz9MxqZPQs+9NBBi7HbQn2UYsqtZIafNTp2z
ti5gadlxCLu/Pq6ppoaRmIKTNCEz4qHZlxK2JpLf/m6Cy7s6E/LGoI6Txw3RTodP
8GN3mUyg++kvKxNcMehBCSQV5T47kTTUFihoN6fIwTuJr+xVwwV/ajUr1ixRXW0c
RZ05hae0Hkc7xWGHcdmBx4dEtDZ3SoYwP1Q9gYEThmj6nRTgwzoxhDji92bDr8+5
F+Uz5Fq34WtgZ9DFqudHOVcTlc7z28MRGVEp9VBCciB0luuUcBU6S9RUz+VQw6JP
2+8k5442rvyMvSy5NY5yAoctBToMRRCByKOVmc/N46t9WDop1b+I4P5HEsGL19nS
0lYqTH7RotleHk43KIw1bjJNzEAboep7S86b/h+g+hsAKlnh3nZSZRuxS0oBJ7V4
5fxkAUNhoKeK6DTA0BfoTab7LjhHmv6u5txaVys2mET+k0U3k8BtSmm8JPY3GiDJ
SeexkyOd05IRQ/MBvl++ZVSbf8jR/4rZc0v38C8BGoVDhp/7AsL6Yqmdcb5lDccE
Q+apOYyI+JGGS8LRClSvnlJjrHfi8Fs3oUECIMsnQQrf2za/qlWKbaaDC7zOfLnt
9XOWanyesMZrqjtrq5yIHUWHrLFCsaN4toQKYSDWIz9umeqb9+LSImssRKl9t6Ql
F41GikW6VAWzijZLIxXlKRp31gls98sJOi0FOGjpuDx32jivCGuLlrSK28OEeerp
bIItPabENLDGNttkUrQjaGDjUBPwerKtXcQAhiIrep8HUq42oSc007R/N+9sFed6
yRHcHvqruGOUzy/mlQjqUcRMHQuI4R9t4PFH6UkVGvXA0EbntH7Cpamq7USOLacE
3xkO25QtXzNMaM/ritMecUxjPQOKzt1ZC/WL4sf01azj9ucK2EBJXbfKq4mNUNp3
6eaiWux4rBfRUxSQSfJjqnodlBsT9qubW2wJe/xa94aO1xBmSwXaYwloJkeoEloi
wtvlBL4N0GT0Bg4LD4DQQsRwMRYHMbIUN+nZVuh9db9BvWPXwToYNFN5N09FI62p
UzMHIzIx4A3YUkcp5IhTnvxds+8efb0O8g/Wtq/uLkGo8am8zJBO9rib/DsOEJul
9UgqBeFM+rUVtU7zEcB2kCfSyQdn/Lo7fJ5HTWJh/6gXeHzJfI6jjMgciGod5gyj
6o2TEGdQTY9pyrg8joV5MhSqcLuBTh1fIegoU9bnn+M5JraVFC8Leawo6/aPfUj8
/toKitjrxQI1K/4a0VhhoObvSY4YoZWa3NvfUQw6fcJ8KfEH460+EUKOAtiUmZW4
yqTg4FJj1qMKrH8O6jC5rrQbofVgGoLG/3YmW08XG0gx+0C5uk4+kjkuq76hJJ1+
MCQWVRRf78WevFkIsVDB036QAXI2TaWsvute1Qx4qGN/pGTOaaeaw3qCA2Bw/qnO
1Xpn+fY2XyAzQa0AygGg35TCzKgrkHp8jKRo3CaGCyc+fApALeuw2ZciE75ocqdk
D5u19Lnz7OJSm+OPcbHxgRBlZowHec98qG2DqlgWIxeGYiKesKCZz8as87JBQLE6
SQV35XANSRkjeQ0gTBQwQE7FifiZFAm7zwIRu7Jx4OccdEfjIygonAxPmhYFbCav
j4xP5IXRS7V1kYjVDnC5IREIYU9dUeZCDzoO22iZmueN40KX42JH21ZHG+hPFtqg
BAQM4XK27pidrAKARWqSdC0HeCGpZWEKKSih/6/DfZxj8Ei6FfHZvlNW1Bofidoa
1ObyGnj/c2GYdYrs8DARbeJV/KX8GbvUFVyBvqLT8KMjIDul+0iC+qLWW/7wiQo0
2BrYyVafLS+uiB5V12+ZbC/amonoy92xUGgop+V/T9Tqt/QKKyQO35g24CkrDq5N
CV/ZGG8+Akxhs8/JOoNKadlRVj6RcdISxSIC2+E2Zn5zdzADRZdKzOs11mJj9esY
eN2Xb6mtFJ4p4Cy1GNCowrGP7E+J/Yw8aShGfQtbVFhfyGKX2LriqpR5N7BJtO26
OkcV08PlNzESpH8b91o6dGIkEYhYXrFjthb0XBJAqPvsizWmPRNUOJOPJNb66Au9
U4C9DWe43G/+SyNmqzHgNCEOk5C/jMRDvjjwJMetPI5NLDVwY4c1gMZGCSvhQ+4f
ie7XV2Lg9SRo6yCzu+VB/SHIE7zpBEjo0EM5BxcMRaEQ6UfpofIcwVYgjlhQqcOP
cZZ1eVqKmT4I2gkg9b6WC/3vQhcHddXej95oqByZ75DXPFk5nUtbwUE1LeogbNSN
rLn+T6NAR9M7UWN0a8zv0G8YP0e1f5jB+uU4f2zUK7xcUO1o0AkMpTMYQze6WsCv
lS8DxYOSvetYcH4k2ubeKAjxld6qMgwQ5FUXZh4kufAnKpRVp42m1siUEQ54Nd8m
4mYhnypIikgvQaCO/vyXr6KD4Le5evX4sgFL03fWolQqJY8Pc2TnjO5hNrvKwG2p
SuhJ1tcO1b1a6CNZnXpfnA2OftxkTj0OyhIEtLsJZu9IKSh4LrqncSckA6Rx0tUH
Ikw1hHtaBuxswcAHdy3peOQkUuU4mYoSPxfjToGTxkVcCDHR8h0v4KlkUEYyAauC
WMHI8xGvRZmeeF6+D8aBbc46Rt0oGTPZNFabFBeLbJOu2NWXyhXtiI4AH42e/75A
vx/yT9pP+5TiFB9DwZvRZqI+1UasspOGSvzISPCLV41DDwYCV+BSdDXygbiEiOPq
+gY/JT3IugcPfvmPmAVgja2TzMyznGSxESvo2Y8XLa/fi+7tV9Ubj/+w9fYSwuQQ
eZj9he7W9fom6O177fw1qGeX4yAjRUSEipl7zKg2GA87Dvo0ee5yF9/DdxMoSpZ+
FRJ8ib2ko2chDIfv1cqNnIHlNeJhVWbmePD6axsNEZV1EkVW7akSqgPLUn/ptbxT
fkjXOzG15Hjk3goITYl4WNBPgIF4BfhQzPGMKSVRno2qmrr9Q/s8/eyj6OcXdLcE
n9LR9WES37y3I62lKALMarySfOf9xUt7fp3jQRSJgNwbuD5oFC0P8zVqtbJM0Wm3
999PNaTQD5XYPMQ0xNuMqRMqJNi6xL3L4OH+qD9FqKo5v6pMV6HI2zEwoBVHJXpn
5u9hSxPzEbzgIsSFrxlj3sAV/a3hk63X5NUpEUvOwLoNHXng1q94mfpyR2qpdUFN
/WFkDpuVPb9wtTFdqHdB15wvp2iHBbrwQEmYjML1RnwbhI3G0JTRKh5alTLjXyno
NXKRhTxnEVIOkthX2+Zcizln9a8omI5dq5xPw1fGIOUXfQc2EPjqaWqUW7Z+G2rD
z3THJicU/2ta2eDiQIy9264Z3Bw/RsbVV24JcXEA4X/CppFdlOftDTvpQsnlridH
NATpOdONexiLabZcZt845/8q2FTbe1aF4Y7bIjcq40CaziHESkEu2Sz3ubp7ih4a
lvqTliCssT555HVOSlTvjg5LQXN3RJU2yOGwA2rC7cFwYCMSFtwhIaXVFM1hy1p9
04NCRr9V6Iupj5KNEs2pxAPYqmThFTSxt9/LOfN1BmGz9LnXQ3Wj1nVrzQDIw+Kq
9AXhxgg+8zu0yzKurOPR+qXBqLMitKQ3uWzfAORJcf8FiX3oyA4TsgBQAuqI6Ahf
6Vo0KAiOdbo/h/bQy/Cxm4KlrZfq7iEwkh8Rpdr3xz1Wj8jzD8qG2SSEkSVF5Xgy
afe958Pyv8AlNQ19p7J71SZ1mAyCPrc28R8XH86qAqZXe/KuHJ5MRvDFnQfL1DrR
wn7slwu7mpBEftvaBBD7x+tWP0+OtuOB1Ydlleyv48qumJWjVFg3G7Jfgkap1H2u
1t45VhFlWzVhwN0Sa/gZhK6TDNOk/h0jEMeVlWlTJiWzPMvvUseXU3Aw3B55lhc3
8myOuUvHkHrPrFRMeVtYSlVF6qs5bHmbv7qk03HwGanthCQXQL7tzh0GkjNlc/Rc
gF5H3/l1w5LHvPBcTdkoKhhXcJY6R19bAgvrW9Q2HMyz9u6eilNSf7WNvJYHqp2Z
NVp8IRYbxkFbXDcx1whNIkdgyV+8uKd50nu7RJmLP7Gphj1EbdpXU06vWVSe4Ag2
6ln74AhxwGqZ0XXS8V4ZV/GMPlX0JdoumdxXvqFp8pSJO492Y1+pVuBr0sGUm7p/
/gfKL10nZc0vL8cq9vWRE23+OXCpZ91Nnoeda6KVfhTlm+1SZ3AogateMNu+kuKW
uMaADqNWR/jpsHtjkvccIoLAbAMKW7XjvbU+IJv0yNgz4mgnpUSg781EZDeqT+eF
q9zPkLuMxp/hhj+bIIg97Ms2m6pMH/tuOmbk4qZhAyfjRNi/qZUm8n8Qj5Up1Xdt
sLetuj69KtMsC9BCfigXTQS9kVr+WBipLtNHebSpNwDT7KwihUgZD6vlY811sXNq
IzZGMQ71Us3L+a4WHUpYLebxol+YWN3TYCa+XTscXVglQrBqJITPAnT7eN/CwdhL
HOdYnr6DAZRQN+FJ8EEl3znLVf6a7Ws7ENXZBa3Yl+CXA3pUuJcIsnOeV8aSJwQP
YMfe7UrBfW3Q+DOET7FXbRZ1LT7PPoRgOJnYPywpRcN6a1rOAzTaziEJryrTYUCs
H8kQuDlBqywLzH3cvLTUPdOAMBBlT3Mz3SFdBCQSZzXeYyfRz9cQrpgA9w5wDWLy
8Qf2fEEydGEGyA7rfUYeGFSlps5WevR+70wXWDvq756ciP59BsiHhqhecwi2gbk3
J8J+S2FAUvbIfFDFJdIm+igzARtkqj5rhgW6i0LVMigOnKhg7oUvzgsudpC8YogE
g7UKj9G935D0NLU/q4ppHnYc29DIZdWqoNlGWvVV1loOXpVYMgLmXZKNjGwtFqrq
nL4n4JogI02lSPOpJA79snX/p9TeJfCfybuCGxlWDb1OcSGMFDnX95HEuVv9P6iN
qppvkcSgoHZ1CEGS8lT4JPStDMaJSaNS6CdfpuwY+Tp+wVjVIPkgXibZHaIC50x9
m5P9Wef+IAMs6M1l2IF9SuEbnkATzmYqJAXMOo5m9RNV12O3O97kx/lto/rJXSFX
mDBl3jhpTNjHs0AaU6qN5mZZFzboJxddFWG8DlQVjEKLYfgsMHjd3w9z/K0iib1O
pn1kPdzHUEyHhowGkAVHXYfrBD3d90joYxfXuaEsmNSyJ0syZT59j2ZQgoMA0vWN
daJGcqndPI12hP5sHQwHCwEG1RFPoXhzx2DXWp2DdL+D+cZRgiQ/DMOZ+W/dSdbW
ccqQGlbaq8XCNau9TKkqwqn0mVmEq6CVnqTQ50lDEhttN/SJWrVKzn7GZPfy1mUf
p/eaIM9HU5fMO5Wx/wlj2Ll4A9uS3pgCdSZIBjxbRdOEEeCv+s0nG1mhPoYuv9q2
3xraeXs7aE/XcDZhjDtLnQuRWUmnK5qNavggqg+ha4YB7hr+/bW38n65aXv3t6Tf
CoGCHkdTlbvGIzO5yhkqfIxiN9BIhydjbrKeKEF0IMRtssySSpyhHSnUqQPUZluh
tnIwssYInOjxKUOKfE2VfUKxbj7J5ytI077HeTh06opCArjeM/8Lf5IYF9dlupHr
GNaSXOEk2Z76a+vxo4fFg6CbSmaShAlKVxAoXnS7WhFz64uXE+veiIxiQKeBEwdq
7DFKlOIeCJ/UmKS3AlznNK4boKtYF31VguukZyVkHVCqGIJuYByOe62yxcQDDA3L
bf2dyUeX4E5BboSQyy0VyJsIqZuiPhQ6sErBnZFhXOR7I1EIeVzJv+GO4zbufKhL
2II86aCeF2pGH8tKE6g8UhkVPdX9IqbFCSpf9++A97y1wh09XYSr4X2fsuKEkgwE
DytKykk0sQM27seXx/oIocxBs64Vx8G9tfVcLd1IlpDbkp/jW++U2fyvzOLGPcuo
Chd91G6RLRU/x+HABBVtcotABCczBkX0wjvYfJJRSaDCnZotyna/LXLQZc9VHYsW
7QNvyN4PX/F1Zww6Mizsz5ozWlA2Zne19BFS/UBbPUGN0BUB0tWN+WakETBq3w5Z
fYhQzfgTdLOF8Da9BIhmGbkUbx5Ng4jg2pz4SsP7IcbpNh242olbHWjB+vYN+qZ7
VgPhzjcITFYk4LIJRJzw7XeAcYKEWWz+OSRmMQi0HuNPk1lfMHOL8jXBjigqaBvA
xGqOO4AatEhjKpSK8ny08Yu9yYO44alugA8RHVn9WYHGWE7PwUsOBFVI3BvMOd+R
p43GsKhCJUvxE6Y+Ik/cmVC0i+ZXw91clookmRL43BXsTm6+yDP86IryBxqmuNGw
mRf4sK7DvfLj/d1UY/rsGT69ysSsZSTycF7tjH49gBsKz4eI6VsTY1oAxUAFMInJ
rafkAfUiRyVeoftvoEsOC3Nwaay0TfmuzgbzTinFoL9Y0ZSDS/dZa1rHnwINwi/r
R+zumwI/2jIckshB9CTt7vyapc8zLzB3bqksQuRBlTzKpegasLXQ+xHCSq2mmH6c
k97qvrRYC9WCVXVyR0z26apu1VKZJU1RvIg9ck6LCelJZd8dI0Xa//NIomYMrBQc
uBy25/0QW8gN/ZX1z02dmDUGcDPdlgYVpWqWVNLH9vfFQCH3ZzNqc2F4ihZEpYQB
7j74OUl67+E3YJpYe/db98xOgMRLPSpniUxVsrCihZkGqpfxeXJcne62OjeNeC4F
9lRNjwwZWEIBDejkWWMfQdv8gXVEMvAT4nOH1K2JZjqZjK3uVvN2agumpQeLCXnx
80xr+/RANcWkiQvKbtkCZH1w1tqSSttfyPKBRzb1r+WHvglx6gplYrEk8NF0q7VD
rHCdes4udjDaCF9y6hmOM/QlyHH4qjc3g/DzzRnti8xPLx+WS/kCD8E7UAzZABkv
0peFF/R8jbDikNBZ5oZvLO/pRU88YYu6BHpnaTXbURRInwysQYRiA76SgUIGCZqH
8lnMOGLzD4wOGQ2dDlhHNhluhRDFWC1eiQ+y5xxzVdWCC0Jh2OVzmX5VwmRJw0Ph
FKW33EfFZNid1OTLhV57RG/iiro4oAXbqelh4LDZjisacqqKwmuHiWFUqbt480Gf
Rmp9RgOj1R1e93VZLtEkvj/ffGgrc7hVbdUdI1qqZ8o3UbErgLhLrn/yywQ6fRWj
6dyrNWSLQ60GbiLBFaqeZuPx6yXvm6fTqYHPJZOVU+yF7bkDPst5YEKLSl89koMD
tdZ9bZde2vw+IxHm9KJBH263kqrcbTqLLUcVxPMqKy2QPVZV3EsWi+mptAxjHU9c
QiRmaf3nU4oRCR+tpkK5/pC2LT9yDh3KF8IGXrYVeuoAWkYx+i767oNEwzj51X/6
/1uKSvJtrMnMzC42WdkxZUB66ANGh0kvH8OQ/WZzyacGhITuvd7/zJGjkTsiPnp7
9leB/lbPi2v27FOrta07XGSvcJe5d2TRlxNSelSslD1iR7RG2USHV9c51P6ui85w
wpC6rbZEEYoB/OXwgPLBdmR2GnuN60+JvQDsw/lWoMNKALpkObaMFoO34/oQ5nuT
PSozSrFLWKG85T4RI/2LBwMvMpshTRzXv+nu1+ey7xzo8qsyAnvuDg6S0b5Ry/J+
zdmTDPvJMTMC5BT4LX8eRObXJqJ76Db+FXKFk0aPf17ohzybQ6+k+3bCpfjJ/KVn
X9FFn1tubn8HuA9mOSRO6Ojk6D2QGfRCvf80TVX4jkNhwb8K7FxAT7+9w4HEBnBh
DlVNnIYjpFqjry3LuzDPPDZ5KSJiWkNM35upyjgqiD0F8VTQu6OhZ09oe8woLjDf
tx53G6DQm/Ni3eeaM61FKPO0+qgjqwS9LGVGBxv07ba7CAfJLCmUf4ik8RjHuu2x
Mvjw096b5I7IUQdHfZ3axHOvHixRHuUueFeXyA0MXiPBJpQ1LLhWTmuP2Q6Tm96G
K9B/JsV+5KEZlVdtZtixinDLmVLbdNwLg1YYyAKgjnk6w0dWtgyOIaXovajY/zPd
3ynWiZmtuYsZbTvVWjTycB7IjsJA6fLF3J6EL6WbpSCmUgwOAYF5nQYoY7+RfU4V
iEq2c70FQei7dQ5oc0mpbUhl10TizITDXeymYpqUebYMZcDLpBBwXegbOKyMImk0
+OZH1sWxeETEpFNqUZ8FxhjhXbLcS1VofFSvivi3aTR/JDwZCGXEDN9FzezP2srv
DNeIeJuRh5l6Bd71e+9qc9Hwl7JlPitFGnk2WLrHnx6j2888dYCY0QyKF0PpDkJN
MvIxHaGpaEvjMqWnnd1lXRCJRsc6cYScdz2fORUSR+ILiS/+MJpvv7YOiF7bj8Ek
sfpfofdnRha5zNdWGZphm1hXwF0ED4HqI8a7cuA3cdHD8y4Ul5pfq2AmZ5OPruh/
cjam2bJz7y3lwSBX5NKu0aIZAL17O4RZtMlgrg6QPiwCgLqDl5zHsZVIxGv/t/py
D1HydJZlVfLCIu0320s0PtgVHtvh09ORvAG3mJSsFIEHFg6AU+E11UUZKeiCEZNN
aU+pMxibTIU/JeaNTQChfl6LESVhIduFbCZ4DEi/NpUT2XQ8lyudHOxcksvdms4Z
cJvpL3EKtDTkfv3xSRG/mlL8vIq3I6GltoeJkum9YWV5XjGbXB6Wp3+75sTTIQ4l
puS4rkwBWXNKkjXpAqhsr8kTX9XOc45XQRRVFSExQUBbzGzTnqs0YcjWo1cZJCRT
e7A/hhugrxhNTEiTirAkUZHURPwB01ZchCNPtpHeN+4BN0UDtCEkJaFyzzilJsGQ
xMFb60jqzW4Nv5l9SausV3VKR+Alz0k/fKSKqF9kwJl+HPNBGz2s/Wih2+j2ENpi
OhGJOryU7VkxJ3aupT2DCrfceQ7qpYx9wJFmwnSeLum5EMp/erQT/TdFMtE4JASe
lOmfWDa5Mwngn0lGUzTFwv3d+D4YETp3y0olqVebYCfCLBX65dqFn7LYJDLrCVra
OuV4IbCBOvlgEKgVpTVPMYKhuVXAju16ZGPi7WxiJ2mZVDz3tOLLG7hlTlYTmm29
HtkBzu2eDZuMurdH++qcuQ66QiKeEXAiz6K9WtMthzsRbmcp/A9alPv3oh3vcaOq
/8ZXr2FWvsAuw4QRRqqp7lrlgtcJaRqY5gkZNMYnbF53yDkukRPyccIrzTjNQEJb
64MvTjZ4E5cj8Z6PumX64obpmaXuSz49B/xju98KXzmBd/2kM+HmpPqv4eU4f2iH
xrNUGeSQ7pqOsn3eVVh/bEjsealI0XmkAEFaDZQNjVObi2ONZ2SuJqzEzsLFr6Q7
18B80QWZwDpz1dZRBmL/Q+HiCn00ATYE0BUkQbrz+70TW4Gx8elpTy8u4jk3RcVu
tjmLc5oRIBBcwwvIZun8juvbqoh0rFHOA7jlby5oYviu80hv0u1WayTrs5DUyLmd
sHnxxV5U102UNQgVNRdrbqGSXZt9if1rYOTcIYgfAxA13Y3TaybiSqPx8oNfdW/f
OB+pwR7fHLDgtR/rXptwleXVMtmKKI2vCTv38OBV2/t0t4/vcwi5l275R3q56oYg
RarUFUHSwA6bQCoEI0LQvGngBV/6MCd1sgB5TKgU44LNIESYHzcHLRU9woEAXP7H
VbuOhvck/Klw8dJpYC9Fl0rrUVqCXbWrxh0Qzd/uPhBC652taJ7r/dAjHN5ZGNnE
LDS2ObizracKn2F1OemnFGakIHVAtZ/5OxQkK/KveN2QarmWh4pWur06WbhQTIWq
DsTQWyHbI5mGKeWGORijsqR+SMLX7dEy9s5L4FfXAYKcOw+lf0GpGx3V3DnG0l8T
bSyJ1Ah9FhltsefJg+NFoJ8kNhID5MWR8xNtK0S88JxytGgfSI+1n2ak/NoXLNw7
HmphCzTRlJohB+rrKZacgmTWb8LKQ659P9GbEhqfrWg59bzzzHUYXJUO08Udru4P
uryXxDi9EzcrieskyjPbJBr9EMgEd6pJKa3HFYE9P5aswDtCD1gzDCLzxoTPbXXr
+7A69V4OirUq5iTbxRAtzDzTKPW0pa1Ez4ZF1urxKUG1oNo+JP43ijKG0dFVEIjB
Tfwr2Lm1K3uct2LiUeYHgYr6GlOCOTQUEf8wpZIjNB7eJPKygwwNSNmYH+DG3ifM
RsmiROaL1WziKzSQblUVRsJnXKSUUrW9uSkEY9psuIcmYWd6aLwmHFfJ+l0rX05Y
9ph5SYABGsl9I2N6c/eDog+/R9I+2+eWqr47t56l5JfWIJc7ZhBku0yOFf5iuymS
2wVGzCWbD2/QMIfxCXjqSDVOsZcxcQSVKdfHrqU085S/gtTn0fgN41aCiMtrWnh7
LU14gefWg/tE6tOIe4aDoRI4JKGYtlgS2PHpDzJMgl1OHN0NwsKpG2baB/ofyjqH
iozgUhvH73m45S1FSp7ygs9TTTFh6sQMpxv+8kIlSlHKfhkne6gdrRAuc9/Tjugk
q8op9mtUwC5Ow/JkmRu5l9p0968uvogBZjCAtWjgF6tnX0U8bw6v8FycV1gVYijn
zQ9mGX6sn9Va+tTDiY9H+rq4Gpyy+GgDKHRkvTw+qmlUG6i95oEPr0eNvv2dd4RZ
fM/O0pbeU7Qt0VImohcukMcU4NK+Xuo+6RrL0OTnSGuccGYmuXNXhwNWIW19qSWU
kbdUFL3VUkQ886fl73Yso1eaykfG+XiAuT6oA9pz9TrkV5kCiq/ZQ7/EN3IJvq2v
PGCmueOJUG0sAjQFiTlpeB9hu9T82Y/G0ZLVXcgyXkSdmO6pEgxp9yGfsnn8T1fv
Z6SE+lfhO/hhZPPCCteuf0jkCtWi5/js2RhdcjXEwK3b0kgxVz5jMHR1wDmcdYlI
S01laGFTnrwSAjxYQtCBI00WWZcRHKQpsNLq01MTctK4mls+z0ZQWknCd9TWZD9F
CToiyuY0VPCifC6IxMQ/jHJvPLy98ArI8jYgaRk82f9qMKUFG+zQdon+kuX9kQjR
LB8dlettdChx000/aEaYTLFoCTHvqLXcijlOFDkWDDVc72YtEsXhVF8VBMCYmo4q
PH2NOATdv5dEyaWEuQFGCPz5GZsTGClGfHjYMQMnA+Iv171aXtHu6RiZTvZqJzlH
tFWzUdt6sD+76fIKXFh1Zeqn+2p1YKMEoJH4Em8+UCa9fss1hAUDrTvaQsg5D1Ey
FTzSe2SWhk5Ww2S92CV1PwCDjH1jERZxH1B5+RFg469p11QoBPEh38Wew6JcBYhD
H6ktDdGylSZOI+SQk49TU0bFV3SwnzY+AyupkjWuBu+Pke4+9A+EOzsicPq+R2yr
6WHp/H7KkKLw5B6BcKIOwsy2Jx0K4hZCl4XgSeqN0iDYncY+YK0Ym+ZeAV5iyiVA
a6JBmW1vJjrfMfWqujGesfVt6eUQdI9ejQsqI64VKoSK1rUkTNSSkShjB5Cz+BwO
bbcC2B62Pjn6bVTY7+sKUqN/0pusLkZZQVAzqmhdcPxIY4yhmQCdjkdGlqmr4daG
RfyErIwWKT/9YLjMg6tqVK/z+tngZbdOgOXobpg845Bw6CnFECkVQVVloJ4KbgLF
HMmfLpw8ygRz/WW41GMW7LLzaTwIPq+fKFZPy1x4EcJJ1la2bpem3Qj0ITwiZ+PQ
AGOEmvWhKPA2QAY1uWDIIWBsDgyMBBKgmwEeDaN/jpxTufX4hpzLbIp0eTL+3JBQ
4OsZWwE1SlyHcBlffkW9SLJ9uzGVVaN2KdLBv6+uKazhp8jzUElo2EpXkNOjQ0fJ
cvr51y85pRZ3Dw1dlsbajkt9QzyIZoaPKL+65patA77pvWG2kHgzIxbgbIRFp1rq
x3VC1p5SHEZsmy+VbVD//e7QxDS+40dPvEsiPOAa9VmBBSQHINnMZiTlDBxUyd2p
6ehMSJtyaJHzYMjVCvdj15bofnu7vLeB4oyVtwSt8CEOrMNPZYAuCmbAeJpV2qzX
PN/wvuC8CJ53LPoDn7bw+mmn5mix2rl0vD3iVuo1GsdoezOWP3OdwNViv7btoUbV
A5iw9Q28oCX7jt8QycudODZn4vpW8gKa5l8BrdP4hjBcpX7LBsAzI06R2wWbG5VX
SdGOqKz65/2/3qVLR1GuT1olgoYLI3v2Bq2ZZQZWbEw+gL6/eC1sD49jg3VOfhUV
pjYOx3oOnbF6FKw3m6vn+s9k26V33IKV5fb5/1G6iGB6rZx5q6FrZW9kYP/HCmPq
YQmTuyVpmz24H4LBPVtcR5kYqmHKMZTTvbZYJnIxBv0tuX3qcRNAs8reZyOPpPf1
012i6a8qDSBZCgAemzc58KZleenWlBi+C899o0BOO/ZgvbaXj0LeFJMkFiolXezl
Z8ACNucEZqga5uPdt5E1ilPxJwZHN6CCOGT6EHt4rtqupvrAP7sOz+dN7MFnednV
K3eR8Q6O0do5M3slENpZmQOYrInLnbJIGszSJzdDqNAQusGR8miDyGwkp8Oiltuk
sQh49cjjB9DWF9WH65L6vobHX5YfSRAC1zP9HteFKSDVBdCvkfXceMGaevxJH6IE
ZAnPpOEv/trkcfEnXJZoRJxcvBA+cOEnHrQEuqi2r+GlryLvRF2ArR0IzclRTvu6
bT2as5ftYukU4rR3UPvooncHM3cmUq02p2oSptshX4XzXAyRBQNuFE01IhXXZKKs
w1mzdc0Jo1eayTOmHSxPZd4uK/Xbx0fjCBSTNaHEyXokFL7vOtR7REHNQS5++D3i
mpyJQjsyxjC+JZAvUL6y+3XPxnDBN6KkodiPnqezvSkq2plaZ7p5EQcFXOK2FlHo
RzQunJVqR/Z1KgMa6XSdjzNxrF/EP95QtNBgKjHxOnCX5Fd0lkn90SH1uN2PmsVt
o34tliCgf7W9DhYFJ0UC5WH2JN1ME2nKacah9ocjb5Xq1Shi4nfBU9v++6a25oOl
oMsDE2PZT7JGclIx6kxY+3VHfm/aVZAvuFPfdHZfOqsKweMlmGeDlGqpWBMY6Ojn
4AzQPea5HGUBKbyGNDt53Ij5hBVVB5ITZBFQY1DfvPTrPl2UBMhkHXt55Yybs6If
2n3cdsoQyNRa27uxSI85W15225Rk3hJ13IxxucZu6qRjXzez7wWdCiya9Bb3LllS
BsQdR1qxR78ale5nFKEJ0HUXjFUUgifyZKfCH14c7FT/6pf9EdVDRSAgzLnjMy0P
UgYBwd+14GbgJ9fE3BsadeOTIMpnMIhnj8u2YaNaxEzK1muXjzN0H/W7ye3Zhqwx
xHGb9iX86Updp4RpAPzEoAezJKlrVj++EtEWJSAjvuWEd2iXT2xwDwU/W8PMa32L
fh+Bv16ED5a+bw3onHmtqNur+7LLu8EFHtAjClwNEGGcC3X2nxTtckc6Ppg+OFeQ
MkjP2s1b+SCRZc/46xr4oJKY3e70mkpw5PS65/SxeZud215tPHsPfXAQo7/Obr3n
kdZavfGIuZ1KYDhyVb4mx2USwEuwiQnx8lC++WAWU6aKtCSb3QWAfc812rg+d+cm
L/ECR4zflNPGxIAxsiBbXnpzQmq+qVovsaDIc8wQseX2W15/wvJYDho7XkGICC3n
WkwsJO12jzyp1h4qHtM5UfOOyofkUkzjy8KWPL+w/6CkI9TQw7T2X+67tUWYzCxf
liKk1Tpt59GDhE6nceT7Y1V94huGg3sONcjB8wYQVCEok2msJ4Ena4jhNLXdo6Zr
FJXqErhDAZBfEpMfI49DX6uP2eEgoAQ3QrG4mgpqvzI9CPOrNUnViXYcHqYruTHm
J1zHlaVGpbda2Ca0CPrlwCB2qPh1ZLkzCKYyk1sKAE0Us45e2aoU7OVka1PpoHPd
JJHy94fn/Kb1letku7a9iY/uiAyaUiEZUMfJryoembe6GULjq6o/EpNERaH3rU/K
x6au1OBimOSL/VH1qm32KZ/DBx00X/tauU6iZ20Mn4PCjuXw+cY9U26PxgwuHBc8
98SbOHC1S4lPtMYJ0HT8t1tGJEUl3E0E2XGqoIxjyKZ5DkFNntZ/0TOgLyOAwrTG
2o0ItCTqxxGhBIhSSWOlnQWlq4YB9Uws1eZfBZ4TsPROOPasJ2i66Uc0eyPCE1yY
AAJUC6q32ce79m9sIRfawXEAiitf5IB+YZ9C4SmA4aqO5GyvH90/FJXAJlA1h5WJ
Z88xCzBYIQnyuhlwV3qkykwYMJ990Zb+ulXXO0l5wplRJrlicbOlrUFGV3plMpeS
xI9q5rXu6O6urGfvfajS9o+AxEdM/a4xdCIypQiqYthNaAXs9hTRu1tewau3UoTo
qDmIreeEs4vuKMjaKSJb1ELpzdOc1hU8IvUocJ/ruSFWd4DLONyZaqoDa67aZA/W
RlZEohj9myuirTVmPflIJT101wKapgE+RLpFp93an0mjQZUaUd97nsWhdbVb8NM6
rnwSD/UX7zJdyVKE281r/XnyJ6L4TgzGdPmcQAY6lw/aVXIxEGAqiwftRadjSLUs
TMVYF+8gAnYltdmyURaXUWiUvrB7hQa1APnDkK34rHjUyvizl36HA6mBsz8plwT8
xRBsokwPrA4ocWaZnWwil4SHjSvzLCVsXtBvovYZotuZ+7b0j2jUPmby5E8mr3vk
Cbk7WOfTUi8C7B1fH5St40BQae8tKXlJRqb9JmSvW0uma1Iu47Lyy5vArK+EB08W
D0kjxAULgR5/0hdXWS1MRghLTZfojJ20CshLXPepXOQiwUzESK6osb93TS0K401M
fr0FDOdL9CCUrKRqGB+ePKxVrpKLpmALqeuI0i19/pqiLkUfbfZLyloxZM+HsO9v
g/hw/YVlxsElYg1oR/zu4aI85bD8rfMdN17Y2Bm6EnszWSlARf+VDoMdewe7BSV1
mO0Ijgrr0qrTxSOcTtBjT7SLo6ptUr2YcS3b+7+jCI4s5WDQZyDid/fPfnPGRw0Z
XOTW1cvjSaNTmiokbPN1T5o8AI7JF8C7A8imBehZvs5FdY+iwUYiu4jliabWlOuF
/rP/LlomVFslKNc+7qoKolGlewb7SYbLqR8y74kk74TF5lEXJab8stAOW3kKuRI8
jRXbpUXM7GAnyw9v8ZTBbcqcINDYK8/vrQ9bPO0+IITdGgDgu5HpnuKR+wtdxVTC
4Py2fGB+xUrRuVl0BIF7APVJRJpUvzfogizhowUESPKv2uujwgST7ytsMhJX07g3
W8x7ZVBG0ykpYFA9LOxYwC3yJKHNVBGacHyTtiMBCPp2a3dHUKLpjglNTU5bZuIB
tPhFJaFxplDLaTnv3ucY/0GgRM+ss1Wu6xdtezmm7AHONwFv8ibFBn4oU+Yd5ddP
v89Q5Y/NNjCVXxlcS1Bst9TO70ryWjw63q+8lYejnszcE0LdJuaICNQf/2DtO++P
4OoEB2K2WvVTrzbiYPL2i1faqNHSySuwpeY/vWSuyEs4xP5GYtTspzeWwWXUPhYM
saGW2aEeg9c4BgUKvquY88NucbcRKym7iVlf956xPnruplC1HdFZdNtPNHSirXcr
sxkWzkRm4I7DXMU1xUPysiX2b/bgPxd4YBA6rXZ73mf0cwY8xdFWNOG9OW7xIq6h
QBgTWyQMrDyLNeuckEYaBKTdRlyQVLukbTEmdxm67j3exDG5rTZw60s4eAnZANku
PVdqKBmaHILBk5XMQ+GEOowT+I4clGLvebYqTw7X+rWav4ZnepGkRbrMiwRu7oVw
f3vhi82WY6LCAXydGPt8jmhxELwsw4skG2w39uy8ww/RL0RJcBHbm3AAdY8Fe0eX
P+4G3mPhzHUbXwtsEeuBQmH2bs71UZqaxpLiqJW44IPkNgCy0/zCQp6Vp2JmsRWL
pevkF+1wXjMUI9zebEYvcioVEC+AVZefW7ICeSb9JwChzWtGA++hy5vaMY5zFQaT
5Y31XYQf6NYwE7XsV8UP/1v5j9FCap0/fg2kMLbyO569yzRU/5SHZuHzilX8fuuw
SoWIj+xLL1ejOA54Yvp4RWE5jAPPMSFg/Ndp3fPkt5P3pTdVk17xiR4p5l6pZZsy
3cN7cZD8r6gnADj/Jac+0t6KFBA5TmFGOkJmeKrWUpUTS7d/nSfDgh4LBTGrTo79
AITCJouZOyeVNJfN46NmHh+M8vaoaUROVHAcsX9Az6E2IfqdhXLzSSshSbS/Dc4K
w2538onivi7EM8cPxsJaJstjFg757xsVBXz+EoL9qym1jF9wUp0IJUdRQmIl4zVs
DLV5rpI6RJJA+cA8sM5o0bPt9FQcBmqtzZoWsCJeNvbRZLY+BMl7S00xgk9GkH2E
alKUcxYPO13AY8oliuf9RsCN0wNb0FYRUwSUn11agggnsvluI8uhfYhdlj2p4xl6
DdRXtXMgrx++mMi6rWJp7oXAdc/xP+bBstwVq4y9cJdUR4F7eh5/y6YcvvGZcchs
/qHFDo92/AT167r2ORWSlnm3WzuRGqJYQaOW/iymiTXBfDq06AB0FotZXE8hiiAr
TUQAkcX2D69Wb//MC9Fxz+AEl5i+rFD/kNmVs1z7WnNGhRoC/yGaQCl2AaO3/OmY
f94lT3oD+XuPjZ2l5vsqfpDD5r8d79uAxiMyiU6hTBGoYwCqgGohyIMyHB0VHHmd
5J5WPWnl6bEwg/SoSclJDTik6JxiU4BSUZLWckVXqjb5yBL62nYagiGZutnbJjtm
jDrCvFgNqBTao5Do+TiJYyIc5EdnJOOXOXBirhn8HLAIz6VqWUq5yvePG3F3ub4B
yVL12fdD2eEclzJL71fB5IQRQ1fmjeAkX1g4+hjcBtklTh103rQnfK1POOenWa3s
WlpcrgvK+YLZKS1RtQ5MkWbAS+h4RRtK3Ufl2Uc2AOigMy8fM7xrZGfHOCEWDOqq
5SwUXHFuyqXOOLCt6gAC3ljbMpMMZRL+nqVDxPxX+GSD2YeuVOxrkvlNLKaU3dRM
qcNvwvpDfv/jQQVYtk+crnmWHXOSt75ogF7qHjpMS11ROoyK1hs8DrFsszwHRpSU
xt6TTCIRDZ3d1r5y4E5RAhURvpesb+2Nc2Nny7DzB0++G2kcnl9waMT5E8F1xu0D
2n2O6cpn1CJAlJrXwnsE5EZWd+z9U5Bs+1sKeMVhdR9QJHSrqfuqc+FgNkQSN1q7
RAiOcBQhmj/pSrn+qbhzL4jFir977ln/aoX2GyYqddJcaPU8tPNbUxOdcORty7tQ
aH5Eff79rk80MrtjqeOaslYGj4Wdpzfb9lau+58Ly8IPjsQRW5aQzWBb7iRp4ept
kTCmByk0YlFo3TQO8D5ks6y3S1lck6SipeFhU7NDuvqzE/glRfH/Kg3kNwq+xtPf
EKLTe/niO+AqfyXqWFgNjSXco0ie/yN3ysEh2DGDnWgGkHAJ8HU61/oQtsBTBRqV
CfoyypdxKaBP3zVchzDNlEOMOOZSmjyCAQjsvDlm5MludV6L2rjq2RdtiHDj/ocG
`protect end_protected