`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4368 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
dnVBOIGMhMFpJZXzCENQ2LmroQF24v0GISR/A2R9ba/HnNU9CB8qeCAwcHTJZ8Rj
RtM4RXzGs8Cb9Gdm2zEVSwqvANlB7hNm9F/JwNl5o4CNc2uHrmCsShgN8ZsXWZz4
yb1OAMYFxcDN7T+eurng1AIAe75oRKrdT5o0fzCpR2KZEFM3AimKlbhx8rZo/I7d
h4p1Ukgx82qB6nVCWTC4FMKBIEVSrn52hxgs2uB9nLrvBCG7IqIyA2V9H1rJdtPy
3Xl2XrLqFmkxjXIdjexku7acjKrc3yteREFEltXEHQLfhy4/wcXbagaVC1DqPFuw
ZK5OarTfTw8Lya+wnLVy5ERpcV9IeVGRgiL1WPtnIcqZpgzJzNY3LPIxwa3j706J
x31+kuesjBu1F4VVDprKOXkXRK7RALzn4dFhNuYm2tdRPDq1ycyEZ7yvwWMYJyB2
/Tn7IIDrF7SuhXHUyBwN8axO3whIRRkjZTMlCMFvxJakhcw8UEwlRBC2OSw0fP+9
XPoTjZjcIIf8UoJjSQFE7UB60v+gtwMMr0r1+PWjciiIL88QnBDkmCZVwMNdLOwX
9T5+sS9YEuRdIWBa3zrrbRokf+7nDLkPtvCSfHAHtOOLXAUmIXIzS0lEsqmuf0hb
bqAkeNJUBoGBDOLx+beOtIKaLgQJO+jgLG7Xvy7Jr/EgKxpF78qQYmLnGxneWk9c
HHXpCfpB/ye/BTrbxP97YOwXNmn2+LiI3rb3UzUchAs3T6H29/74/lFtcpLCSqNW
qW9DxxYzWNw8MqqHYSXLx3lWvOurMozOPF8oAJ2+GL1O3I8kCvWNcugJV9+YB+/7
biN+F5oqqrrM4/C/S/JpZbm4JD8AawC5gwfGSY3/DOCA86n/jARTGmj74T78DxW1
md0rg81ROZc8bj1QAOE9fsGuenOJXtWuqyZLDHMpEu7WGfSKXjsIFmNXk6mB+MCf
eH2NRP+jfOS6KqHKXZB1acZ4XO4frbt/I3nG1/iiUBii4TF1kLTCsDGj587Svu/T
rSpTRWi4jeJIbRvmYttiHN2fE+AnMT/rFYgJo7sPRqRelGCsRfP0+MctLedYtyXm
iIfNZqAIRCsl4UhIsXI3rYE0StmM1+Zliqqihwmj+nzyeUJapUhXw2ikrX1yC4S1
sObamOWZ3cul5901Ud75pWUqkIep6yFkEWI7FCg/hTnS+IgZPvlmixmFRsiYaAJm
ZysmPVwcPOixTdPXWwpQR/EhaUf6BjuBc1jNsG9My4Y4/9SoTii8pob9rYfoC2Xf
jiXglWvINsRvYN4L8t+pRXnEQHQQamVFQWbsCnHj7mzihKCvFa8BU1Vpyp2CNOvL
TYajAg988WMRpJom8YEiBd8Jw4QdadidKaZ8qmvhN85DF5HzxXwqKaLgM2XSyBST
8WjN0CLiRhtEdOx96kMc+cYIleMkyRiMhfSbfDpaEKnaeyHe5QxrpFANkLjnxd6D
xy89dPTAl2Dcd4+SCzNq6Wa47ypxTdSYQ0q/7d40Vp6S9+ZjapuHf1G2KGlTuF+p
ydxufnRKl93Bv3/F1/aEyMJZIueqsPoTDJL6crKxx5IhXw+2qBgJJRZ2yu3Ix106
90aQx37ruvoSrw4rsJEXNEnh9XkqfPYmruYKrM6KO32n4XwixoUXqxtLtYJh+a9I
bviULGvkTP6ZzzkCde7J1Q6Udx2NjtyUoFLvRGTuqypkv5AY0aGionrm97WZVpwI
+PK54pEHcNIAdUPJoX9UgUsRPEEv9+EaoI/0wicxWHotq4pLi3Uv7TRrs1OAygwV
U4lLSwhXqK6OoUUM16IYcHiUcdwNse5PZfebeaH8VBMiJLEW+wzogm/X74pU9OpU
f17gEGwYH1oJMBXgazBh+xiwpPVy3ITlkfT5YJsQ8l0ArS1VjIjAcnW3PHs/CSj7
CyoiyEn1CAM8bW5s4AB8CUTEMBKCrFDWogEW/BtBWKv1DJYBvqoj55H8zUA1GRh9
w9CORJ8gw6QMzIy/Tp7X9MZrh3QzLlcJDklrofq4EAjvtQKxj10GmHI2Y08ru1HK
SEtQc6HUzdpmYs1TO77qyhJsEVBNrv0UxyfoKF+YhEI6VuYJSatn/O18NOqn0ia0
kWIgLvVu0mb7CPx21QeLbHzyt56W8L7Zj7fjFBNwxyV9l2MEAf3qWJTWrQuaQBQE
KQTbb9DL0L4px8FRw6MfsmWeoIX9ArV0CQJVjZJHUraHINn3fBBrpb/kWLb2Ykoz
AiGjUeEebu0aD5NKZzRm79xYVIu0ti1ZVkO3eX4+UtGpORoRxzsBxPQDV8wMKJHz
qM+jNkusoZb7Vjwl0B3NslJVYgRg/aBUoBtuaMg9BB51DzJtNRZ7av+AsL7ZGShO
tRgUBRlCDbQobmNL6LWh60x2IW3d2msOOL4GNXx5k8pSI1ylerll70lSavNLCYtU
sq0GVZPPsK55Xzm68GxGbwMqDRCikUVQNtWYOfe64fdsmf6TH/ZokAn+vWdJwmAo
Q2XtoedbwTIoqs/L+8kzQpcJjWQfjnZzs4RNIxoREdJ2kE8/1FrJQ5GpBAUQs+qI
YLVBVW+Q45XQMN9V6woh3P8pYkuF26A80gww8k+ctquQkzD5Xqv6mqYF9Ghn5qH1
xfsIeiLaST7yfN144jnSJr2PMWucSPocfkjPKtjtetbDgadKeAELQMyV5GMoUSgz
O8OGc4gafsBj5n/9OtQe55gYLmWqXvZC26ZBYfxcL6ubGJ/ZaJMIRt/roGNyqD60
Pblg5FIOKS+3x6FWD4NJ3/5ExDi6PSEz35NzOEfvd51WtWg66cvgOrHCXNE8iNOu
qwwrBGv6i7ddvEdOxNWusogHFrQSp/NMf3/vA5Kql7L32Hru6DjPHVRcnXZQoziU
6ThHS4CnmFczWSbj2zK6bJtHje88V46+Zi5KXs9k0sqoZMmiAB9dMcgqKn3FwJz5
3d3BrUNB0/LIKImQRGFUTSrmtkDhueVx7RkZ+7DF1TpQE06iLGHRKDtgEua91+9D
xPAs6tXuk2DDPjhr0OthaPpv5Mlr0KLdGNr4TmdEWs/LDd7Kd2xOmTA/ONjeUwdr
ty9/9TNX99BCL8171/632brV8vr+AZWab7druUpPrWIEJT62PyijZIjXjwDN6l9o
Ss6FS/iR6nPXoeMBRvxZD6+IUJmyVCYBMEteNAmoXfYvMu/Gl5gxvSqqtyluPLiV
ABCd+8YOvlKBSQJboWVw+TjRul/rQ204cDANDrkqxzQFXIrwfA0+ZNuFIfw1IBjJ
wjUHrlwsvFWRc1jpBadvaQrUGq26MQMCUWEPjvXVHwPi9fqIxd8Wxr7ff2rCprcQ
iuTq4EpJs/phVPLogqQYA0UcBeXsZpbVKqosTBBZQqUHVnu+dr1VCFfIAO0//y7Y
T7ftrtg3jRpwFf6rgtzAM4GoQ0wy5GYrpN65Cz+t0UPO23zrf2C9SzvF545xZDPD
TPmlP0xe871Hiyr22uoHCygVSNLwPRpih+4ahpxjKsKR26Yu/FCxXJoqb1mld5L9
0tEqQYxJUM14PJzMNT49mM1lUSojfhrjpqV6+d+FNdW2EeGicOb0dxxba0Ul5TSi
afwbzScQX5fc3RvUwEjdxtyQD1+g3mWpUBvXVYZG+w1u565JlFIKQo/O4R/wkYnb
VXHRzBU1r8fASxrbHX2MpT4Is/crdNaxv9uEoNYspok5G7A9LNp3+PlfO8q+9K5G
RnlYkTBeK+kMWufxeWsyVHyI6kY0+P4d+JXJDXujOFw3IacBWcd/b0jn+GMOxuI3
kfoILp5s73i/wiisl7k1XmWZJEcmv20hPGc3KHlDI1+wEUUuuexe68Sto/g0xeaM
Qkq63sJT/XjXsZil1zzV/yS65DQPt0boiMiRKL+228n6QdmTbiQ/81MTnPKvFEld
mxfEI6Hd7m25LvYAgTnSvofnsuDxDPFmkrB9cJrfSGWzmLXt348QZne6mz9fAVQf
YTbuuIwuw499H4AKbIpRW+69fUgxSy1qvjAcnVb//cOicU6eUgmzMYQiEVh1jHco
+ExjnLHYik6UN4x1KF2RkSxM2G3v9WNCnAfnVcIxvPOl6vvZa1jYufzzvJszmSKa
+FrxPpeEAobk+2Yq8waY5xQlpaJD57TlZHrQmCFAOfAMvSr98osxlqYYGqT2F+/F
hIPFd9QkpwD2+ZPq/fd7ibCX6km6Zr7jpZieHEJoaXWSZfj8mx6vvUFMXL9hmk0R
AytzB/VhNc5+rqMCUl3njJjripWUE/mZO5/gxgwW4lYSZ1fRoYS0EIPEwA2yc5Jh
kKylKiJSG+h1e551hfA+cptj1gziopjg7aS2p9QIHcs6Ohb3xi8Hvdl+RumjauUS
Xz/ZmkJtRhxBKi87UCQsTwAP8rqnAeIYhUMV/dfRm8jqLGewZKjbNfoDdjz4354J
KsOYIk6hiUR00u4xIBZ8GHr5YYTpJlNUaELJd0gg/E8ndtgutYyEhIvPF+LxjhQ8
hWUTWxtC9rhd6sv5jdvv9KtztTcB8Vsz2aPwqsyXdeRSAha+Mg6ABkNtVd1IbwVo
+s5xDNED2TEDo68qU3+ZgH2qawXBHRcDF5MH5PvCDc/WLY6hi96C8t5BBcdN4bIz
0Bt/Ruyj9Mqi170qcMIbzYK/pD65Pt0DW96esFsl4Dhi1N/n01W5/8uQIGYg4QvV
IoTSXW9kJZFKX39lKXVUzfTBfO24VmiqV5RbWSDTAduEngEN/hSGtcKAXpLrMkt4
G3XKipXHQYieHEwCpb2ukez2eNuJRONcSmjrO0IDQ9Wcibyi3ALJh7R5J+/vB9Y/
/N2VffJb6+7+kxI2D6yhF+zKSE7sDkoHE23vc5KasFGGvvSo5HKvXSo1fJB3ncq0
uwP14nK52MQvTfEFR+os+twvLDEUHU4d7sMPVzXo/8ZLTZKPdSlE3a1QQIkmzDn7
T6aFwNN1GRUMaz2zyVmbvTKfBd6zFDLuuq0eGKPi84w/pyPN3DpCsmHvSQQ5dwQp
ZnqbMBHbzZ35mp4QuzzdQAro/x4uv3xH/77aUXBK/9fzF0V5QK7mZTvqz5UHz9sZ
d4cF3+34l/5M9oXqegsYTrNvxaZxr/e3lNxVpOF1gcxHQLsVw4Hqd0DMh4VXrC4P
uTNveiP5K3uQLzpOfI+9VBK/jB+7bNoxWbzKS+Qb7gELfaRki4i1DppVi6k68O1q
fHpvH5tVrArtr+OVhMT241YI7tvWTiEYAsPvcU88teDhohbWs9sI+4slUIplTNgL
Mfq+70kUf5XXEo8i3F27aeXqD4lS3nw5MgOk1ZsuzboHTHs09CmJSoP4R9NTjXH/
4iW4jah8FGyPPgF1tIJfKf3MYq9IJC2CUJ+9HA8M/BOEqebCifD8IkQ2/sFQWmZG
0jyi6tRAUixEru6CGAK+y/h5GOWNH0sSlg4qZWJE1Ek/FVn6RYlnnoXZ04eG0R0l
4q5yNGDakqWCTt7eR/rWc80YNe0AcczUCg+JYTCE82i3PIdtoy60yuOjkIemLj67
xoHi+hL+fdCDXNLfj/HkSuErkTTP6AYVdksSC6PdJ3mgOout/+I9KR3PMgm5wIn8
W1vdzSomfuDIyq+f6gmlSgk3EQwlOk/11ZBUmbbjnKeAYpespMWI6fsowdkIcFC/
SNhyKy1AKcSJ3qCP3tfMb7E5+VyjDj50skC/dWQatq32M8U/p1dg8gMYrDJBjDm9
`protect end_protected