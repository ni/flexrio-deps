`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2688 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
9oM3kKfrWu/c6xK6HsCF4eyCFdVr5Uy5aj7+c6r+CWmPcNT8O5TIDpxiODNEez5c
kzLLqCqBROpfptjXFvo5hEcitAYfbLFgBNpCZTF0QF3Y8id/IW7uGOi1x0k2cORZ
/zKy2/rZszESbG2RodCYfM+ZksFBlHBSW5OEq0MipIFZOa00R36v8CRoUOoMOT5A
U9Zfth3cXgsqp0ecJk74GEJxq3XdOQCvqHc3rMYIrMxDoTaL9C5P3QHnc/t2RMAd
yx+y4rZazeA0HHzR1NLULzV4ieZZstbTvDetSvAwdXh78bGuiJcWc3ym9BPiC+vM
d7lg26pEI+spB3SPyGruJcFcWHTY9HhrlrmtSOWSqLnYv4FMSL+SYXUKHIi8hvQy
+CuE/ezZqH95aTt9XXG7L0ZFy3JMGVfZ0fgVc8eSIQTcuXhEIkUtRDizuV97VPFd
IJM/HPubO2yMpJNfix9nTbdyJW5MH/HMvwrUv8Ry+9eq1IoGSFUVHHVMmfmYKrIH
rlnzW5Ksb8YqJ7JxnZSICqhj8fAUzCrijhAP4IOpeRbpDVvMc/slAsX4sveHKkdc
gH0kHT05ftVyzKCgYvjuUIm0n0c0M1TpBSpI0OX+vGHsiC9JB47NIntpRIdK+kx1
PdlhGJ+2ovWVZQ2QrLlNd+falXg+FyGvQJdQra9dx7UvqMzpW/HjzsFLc9S1SLQ8
42j3WZlrvdcUy25yghXTRSUmqhWknnVU5gfE0zQXxjXIklyPe4lP/wJBTzi9HC6N
CnTBO1G+nvLLfXs2JEeVfTsoydlgYWCF5A1vu80sCQ0kzduT+pPtDDOX79K3aIHZ
0R5LA1gP7OaYS1oIWVUFtZA9Su4K+0eE7ncwcocKOBhMmGxEAhDR27ZCFDPn6K80
yg53bJjD1tRR5JUrkmzkJ+HlKFj9cgWCOj8QFAqUwYPgg2XRQtn1dH+yN1FNyKe3
Gi+jDIwmEPcjk8JO8XBs6WbOxsMOXkDy95qp8oY7BJm/HUdYTFcT7UOhvGQGAaZb
mwDBivNQ8L+Q8I9GvI4XT7vZ2iEc1ftzhPsZnvDJGN9hjgDqn917pGfSz9+ggjsC
wuq8msi+zio2GSkz7D82hgw5+8DQpcwEKtiOtHlEs2bcELy41ULbrGMP4tE9WnWk
SkWYHWPcnG3e19GM7nJokIRtdeWUAJy8M/oOkGhWEgP1jMGb1qudFmVIJXKr46kO
hDnUX15fPB/TLnHH+FbQ8pe6TZzhDcf6lysLEq478bcAuErXBqKEPRwy+HJbgOLP
D9yzh1zWPZMXAgMa9w8XF71p3PhEGErll095YQ3KdnAVHJdv4I7Ed4HUh3bGpMjg
7OoIgH6RRSJevwzSz1SB4mca0VxnVEq54N9744oLdTs3h5lhWmpJl78zbqw5fLHg
npo2RvCTitcH9lyYZs/Lt5ygLCbIKWKnqqkpkNSsbqL8iB9Iv+te8ZZuWlAPJ7q+
pf1YYFIURI66pQ881IDNUf3C3RFDWennm+JOzol47Gb+2O6J7pJ8j2MqPL27iZMB
6dXRgxT1Mfi/UAtv5XCJOtyS6x+98MCJ99E09XM/4jMduRnyyhK15Kpu9a8tmAzn
Gc73IGqgKBuW9Voau87/Vo5FIbELaAIQnCQxjW6QGuCYKaV58wiQrTrvA9E+5S2t
vsb/0NXmN3ee0w/8AsgbTJkAeXDZYOzzjorQEFSeMLv51tGWpCK0BZDs1IljQ3It
NSUNCCnLZHYEssvrg0o1Y2W66uTiQy3Y50YbkpHtBFEPPwZJEisr27mudgC6UMHe
OfOqciG6viOV6lsNakBjENFahptLq10O+p/5z/5m2SeK7CWQNvviYmajNcKeSNZn
7nnvD0uk4o9c5vCFI4Sr3gHCpdm0n+hLeZmgK42RslTGy/UUS7p5jh6b34saa78n
KaAmydnZh+UsLHPnNmKWj6gFWUTIuBXoeaDPfqAXFM8tFeeq/E8BNbeVagcRrcQp
yBGqAfmXXh7HAQDvkbZI5PDZjBjD+mV8KIWowTKBkPFQuSuUkTo5zkKLIfMEldV5
P1zQiKzb/E30Ur0ufLwpr7uvV42ktEsgmNpVjauJZ0wSIjmd114CsdqcP+t5UTyx
7gFB1z4kfr/4RFg5y548dl5awzSMUfuqcc9gKDX9rsXqI8ZHNhHlR9QMDZSGiC8k
5495j8FTVk+Mdkm6KOcW98hfvmPSqslkk4vPKmTTG+/V5WCnScxoV+pf8EHC0Azf
75u3cy2uR+M51N5pH1IG0RUOrisf8kzTKExSIhgp8K65jmcthl9Iro8JScIvW/oF
lAh7zn5mccIvJvxZnhYnnXkUnf/PCc7wUpnN45tucEC5SVwSGQ5RMpjijUjqlctU
naPzz8vW9ullupLHIUJIAu/U4T8UR2YdobdMt7ZnwYUdyCGt0K2iXtUFx9rExs8u
ZJMEMWJHM25EfCGpAXexScMy+zhsGXPommi7os7iVFiV16cpwpfiQZZ0um7aLAgd
RRdOVXPF3qTI8DmTgCYIZHHW/oL+UWkwK/cyLUuj+zRQ9AJ6zDye4gWUqYZ9JAK0
vWNNubVSweDLTjp8HTK47b022e1heU/Rg8APrx9SztxSTM1EBiz6gni1SJfEwFeJ
Q3L5Eq0+WsOZW7LAPnrmMzk4qUWVfiM8QnrubG2nY8tYqeQ4vBvrlJ6H/9aJ4KTK
nRwONfbHou8EQ1DCjR1XHj5+u6uXHHGD3d5OFGRud7eqtUm7nyIqObtMwBWGYZJQ
En09QUtEhGvSTNHGMfkvPc+ZFJvwVjle5nAIQNgMYIluuQ0kTpIh/Rc/HiYFLufv
k4ZS+o9/To/L4PV86L7WBKIjZ+RHd8c9z5xOPGl9kxzLeQbDm02HR+yknxq7pO35
O39TYZSYq9S9j4xpwGK+6um6wi/pAMzlpB9zEIlcvDL58Y7/YvRwBkBFo8S28Pip
gW65Q0ryFPHPrnP5VPvvs3OeM31xwDeW6pmQpc5VOt4po4+wvTSuJb70nXzZdT//
1GCQGdWyc9j53AJPsfXTtfxFURPE4xuEyDOQyp6ygG7wtvf3zeG9lnQUCjpY/DmB
daG8QNI5sUqu4+YCTkjsreSXKE1UZjo0XaShsVxpetsRi9cy7aeh21REPbx6hDfz
g0bB+g5wsEEQVITr1wfQxR7/wfERQywma28sp3NjXZbXb8xJJvAqWQMKgvbTVw/4
IsKaBKQfEIEb2L2FL5597vUi9Yo7UxnJGO2mVeMQL3C92XwKK+QlZwJno/Vo0Oqp
sX3mhaLbAQvDzmgcpwvmRcTRP7wAAKc/mrZ/f8BakxsuA+S3D5n0Xm0IsF/AyHRi
67y9WLmFvciyGYEH+shHxV7NzoqvcJWV7VWzfnSPgnPtkACqAjg96TVXZC+L9yT1
IuRXOOMBFP8BYnyOefLqWCpwZhML6Kx5ZSU3NR93y8fgBYMLFs2qAtjGOpc3rwUo
`protect end_protected