`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9776 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
/vEkqJfyK/81z5lf9X8oFT12/av6SK5UEbzlpHrYlnN+plTEcdcXhe5tXR2zaky/
oPxgkE7braOeHY2FFzQLG+OD7jjfBCzZmvG57kG5HKruBO4bu0rrcofa/uUc2mpg
Rr1A1jL6qbrwY0DtQMReQMXkQ8SFRj1YHpEIg572cCz/y358V83WuUoWpmVKt1Bi
JBQG3pQUTVVZbdctWDReCDPCYIJf9XGmZX9R8mxqIxtZUiTv20++xDYT0Yp0embe
AxkXrQUhlGmzZOxFJCDO5mNuzZFzClkhYQTgAjQuY5C6gQgeAIrZ2P5+CSQzVJ9q
Tvcgna530yNpDmxMNK296OAMSWOmawxZrcoMYrYufS18wESRyfkpWnTWbIkTHxuE
UhN0Xb8S/9y+adCbXJJxpzCdib44FCO5N2RtOrTthBP/Ywd8wSQ8kTJtCvWZKawz
ygPiGVwQc6fLwWgtpTCxreAJEmQH90G+rjWxJvgD+4Zbg3uBZKiu/2x8YixbHmEz
482VCzziuDZFRGi2xOJnQeaDE0cqsdXtTXm8bBMG7FQijnabWiKSZ+535ocwKof3
hYk4aOVwleKkOOGIazTiUafzm8NHLBhDCOEYt/3G/1+3K7BBuLH4/14eXj5ozZra
MnC+HFpR0P2EmKC+AfCUJ1oVdIPPqE6OCrxeI90/elUYlSWQfmevo0DMlNZiwTZU
vFUhRWETrjFhKj+tTOegxs1NTQzC4wiGo6Xg3muvgI/yd+nh7XpG0rRwUrPto5We
kOIXrvlWrWBCfoA5rgj3VDVMN9MflvDcd/+irWhIPfuG5UpWUG0lVH+C9Ihs2gVU
tIUSh9LAbyyyoyi5zE3w+A4JngrBEfIA9kYG/6l/xpWCgmwzmPmk9eXVThfTkRFp
yFoNanNVJFYWVcR7Mp/bl67t8/p5xJMCC6nEsFFUD7AMx86WPD0T2mAzagC/bA+1
oMr0jalER0m9aPIQnmKuic00RCcePjSFDx9gblTqhywx/7/JaMW7ceXdWeWKvetd
gNVS2qFyEkj2w4m65tqoH1ZFUI1jsa9DSDfk+KksqvCchphWuOIwxatVPhj099r/
9MwXoTM6+s7r9wb3rx8gjR74/51SM/x8VJO+5G6Hzf6UIpHEkAlpAw3j6XzNvqx+
lvtM5hf2Xao/mCVXKm2Q8Z41wKxGDiB7OTjM62lWTzQDRUhcvdl6AQ23RpwxXQdQ
SPftUQrVshf6JRuAUKuCJusQ9Qf6ku1kk/U06bMGWhLaoZuAKRoRo189mpQ6i6M3
CWacOJk61jrqjdhACrRVAgniWgmaIJLk5lagw2I0Urk4CaBxUr5YAtYoZspExkiB
574YLNVTyLMt28Deb9Ja8DSwTXiPCE9nPmwsjksWmqrlgu5gt0Tx9ah9E7dJK6mg
/izd2l/3DXnKOULiVGe5uYgnNZYbaSxU2Z/eJyKRAq1NVR4VsFvVABgmr4SEeV8k
u8XKBrWowE6fwjtnU7CJ5uoH7W2W/MqNH4k8odQzzNZ7cpxf1B3MxdaqDbOQb6la
ZMahmNiynCHZ2gb/eodlPZUNB8p/1L7ED2bXm70/qcQTTPX0rhqKVpSOVmaZjxQW
3qR633FBLHghZrTk3zd0ec0K0akSoyAfC6hj88DqtEqy2r1ZwgGIt6hCPpTbGeAZ
TX1ZqZ5vyxBSkSBGUabqPsUWLbCA2nJzGj+ob52gPXWRnd9oCFnl8vFLkQqLRhky
VVvy/5TPsqlr88+DCQgjjPbOSpipAIPKwjZ/xI9HoutT3PYLGt5364lEBrepKydX
qfR4UR9cDNaxKltDjNZkhWEaWAh5IE3ZKpzqSglAcVoHE1cS6JrZfszBSgwy9Er0
3K+AVPKl3nN45khK3lJHIlNU4jL0XLfdZuqyFzCh7ll+0qC8Yh+djWZLW7i8TgSk
pAGC92tEZ5/4IntK8GP4mkKZ290ONsEpWYGPC0x8xjxVjbbmf2ACHt7WgcBqri4t
1UPW4eSYZfw5BqgrCvVISux/tNCY8rk5wrhmBDhYHCt5aJa306V++wAxzCGNxVgW
ihgvDQXt+w6LXyL4bbZ7oTAqpHxBaF1EcbwYPRlDQ8+xF2jQur6fSNKUv+0GPbBp
4YVOpwfdolZt1hS+1ChfyVVKmabjKNNRno5Hp6qdT6Q0KaR3iiZK1WI6s374gEN6
FT2cZBKK9E094VDSVTlaevgEAd2ElXFc0q0E2nCey9ttaxXFjt0MKQ6H4fAI6Z0P
x5sUN1DSpsI9zGzG3cvdhy6ONeQGFntsS27/P/GWVY2mCQQJTcz7UnsQ7g7Ho7uC
ewVOEGzZcFEjY+AZOo1xHt7wNa0x2VeEhWSbDUByMeisFVjsihHWAMiQWNnEp1Bs
JnzL7P8ADt/ulK4Rh1yy0GtaLmsIjiPFyM6TxGaGIH/n+I/Hki3ndachrLx7vzEj
i6qM842hdfuAt9/elk17o2/1Ky+a5Vh/hv4Um86SkaQ4J37Oq7Bwvw5SqEOR7yhE
7lk7iBPc+JPGb1uEjHg6HT1XP97EvvU7hUCrpDPM9oESVbLHqYBJ7zEGwdU/NZAb
nmmSLK6woBwDZ1NBbw+lBEZtrST4wvNY15B8q5or+am7hD6wVwvp48QOy1XB4RMv
AoIsKFLNV0tvZ4kQWmS8ReZgH1Yp0tTkfzU1/B/2khJ7JLXonr2fiAT77TV7/PX3
HJO/WogsLRJMqwhR0AAa8cQ9TiFl7qpCfm3u/MS0K9w8kXpEDC+MUb7+pTDeML90
W3BYvXV2XN4hnCCFs8AGblH2DcdwQSrjT+i/zekUV2htlq5KtdMW+fRwlu1Be5DR
wTxYpNDoniJOIDeki2ps25e5RAU9B/BBGkMLAYn+kqL1mEbiB2DQ7E4W+bhUOoEy
F8cAahPH952ICuwN58y8fcDnLH1Kj1s45ZShfgRQUtyZY4i/BuRqEwe7EVnaFCSY
kEznf9rsBnvrLb0v9OZaFuaSG97G3bsC9jPubq/wX4lm/maPhRI1t9+dSDwxGcMW
r4lKgxX6AYyt9VDpn6kQqQnBXor+WeC4P3sljrAKi887KWpu2GXAetiQtKz7Tlu6
J4Hq6959vQFxHJlmlQ4aVGGMWKwAkL6LOEZmjnbPrnm/zpM/Ti2dUWbrfkIqOu0y
w1On8JgP3VcPEstKPR3JOcK1Mk2GuKpvi3Or/wWncVF0UPh6HSJgiAQ0/U62ureB
ZXMlchD7DpPwgrLDxZ1OBsGxhIfGNJOrLKPTjSaWsyxfIypO4hlWMHEDBjw/3YIt
MeV3Yq2pM1QqS17yvyKaut1TpYeZYBNI6plhJYqZ8bZnezoVhnCKKZ4TIF0AlapO
rfG0d2kAkgIbBe3J48+BIFGXp3ph8o3SMIpZrEcUYRE/dYHGYRhOtGEJr53Xs7wd
z1lqS2BF1YEclXCEUukEIyAfVojhsl/nEtAS6sN+xa3WhZ7Gj4xiI5aiLiYWcdhd
OYCxWxrjdFP4dZNBV6pwNImDQBqyMhYkA6kKEiuEiSLPwj6n2PV3qkP0QKwH7LVN
i2EncxzlL4mw4mHr+kfWfwU7epeK1UgWsCY+nf+ioGFplD9wgKj3N/6KBJC8dZoP
q95sMvGV+RaBqhen0I/NFf48wffd69aVPZiiIoJsLt59d/T5J3pcLrV41PXQ56tM
t184UldXCX8P48FV1fbLRmNbaPv4kmZrUs6GHSC/y9OIEHl4oUsrk3lDG8eE+8R7
PmYrFyq0JQC7tbvjiLYMR8zMrPBMvwdDDeVdLDRVX0FooFWbEvHzCdMqZXpIfsNP
gdszfHsFDwEi/NmQma7/E/4agYZ0LU2iCeJs2fBkZibMG9Uq6+8fTKX53asQxcWJ
XDJPiOkGKQ9rc1Djemw/Yk9Rl25h+rW2OqyN8yYykLgN7f/6XfthlwnVFv7Sp6lX
t6TfvbTi231NC17I/B7aBR52n2AwwL0k1jlgbEJ/7+5QVKeo2ak5N4pHCMZeWBF+
XyKIh9f4zG9Yop2V7olCCGl8+1pUt2pzYuLYq3nOzIBkX2iXx0wUtJV3lNIfG8Mr
0dNuoDNPV1sMUm/rEdKMqFfTwqZxKz+jNZxpGZjst5e1Sap8W96VLkjidmXmrkAA
w9MioYLmewfWds71gt3vsAfvX4b8Vp410PuauNrFxIo9XX6+SXC9YsQ06bUKnns8
tNM1f0ANzqK1Fn8BFmcTNVTNWtncyx/aEnAPupboBGGyWWucKojSoxkkayK3SRU+
UAKBY8PCSISc2MhFdjJsVgyGMKQ58c/aIpZBQAbwTp3qayZA8rDsLyNbAyAAer5B
8kAmwGUeWcZem3Dxtk21loUg+rHsSR8B/l9WNIEpk5OhHABdeIJ5UgNZUUTEuScU
GLGISOOx1ST4pd3gDQV6xVvj16+zMmZgJ/KJeICTzyqIfxZI/OmU/6g6g00umrTb
6Gu5eIUVP017uMYjbEjdVRzaEoeR6s62W3BUrlMHSNMsA3LaUdId398xmIH+R71k
BWwKen6n/PzQn8ZdGOEXvmh9whq/H9UkGhrLdlN1Em7fTM8Fz5JjOv1dDiV1L478
AMx/+XhW7rUH0+HY+94UoFa85lG0c9x3u5HyLFJZ+I/bQotUFTlDas7UJnpqzlpq
oGaYzau2f2M3M9V2WQ/cvMLVwQLDUha1k57K0/cai5r0n95+MGyWWH989uLjyHd/
Y9Oc4QzuyegAO+Q5ca/qhhBPmQl0cd3baYwZEzn/h+3/EjkUrqaq5NzPWS4JlqI2
14oMeaRjMo7hVE02vebDTD3Kqzo8+BKzkB/5VbBSVPrKa0GSMdguFwHMk56hupwm
teCYa36BkW+3Ym8Ntt/JtBVmRIFRtmLLnv8bFKrImLRH+6D6qDynaJ25rbqR4Gzv
qX93j8yRv6hnNCPHlMiNMF0yTvp7t7pY8EtW9NAkb6gGuQAM/uMN42PjzaDmVJz4
TwbznaUBbdFWbnu/DspST6We1C3UxpZp2/dhspVL7JowAuc2gDx4VEIgWfd9Wgnd
uJ2EqAS99odPogYv+EOOMiYGkqU2F6BfGKF1lHCJoDaANvTiVrIAn23kCz2G9trq
FXP+hQ8zw+Q3dYBkPLl2+miu73IavRxaUGwPTNmgjZnmnIxuRAF5B7HdAOZLHSJU
HFZ5K4I+vHmlnMB0L6C4Z1zOPwq2g9zTV3f0YtRq29nAE75r9ZTjdlSVp0VZ3Kup
b06JxAP46NX9HqDlEWmO1DezwsJESYWJ7YtvIyqFMB6c2vWzWHrr0ybg6EfDW2wC
Adyx3Ql3MIqI2Jb6Ljym7GhQhq1wAAb2DRmN9z4yess7c747o4+yNIekrI2YtK/7
VLmbeQ22DdxTI9j3fkAUZf4l0xAHyF3y6qKsETlguZRuWt+7CgEAikU9oxAyRTLX
I3c6knawPCRomD5IYYoqusi4PAaTT76YthCuIEUmMK0LPj55ueTk/BuqI2ma7IPg
+p2758XG4twsOTR7hHzIAQnax9VIzqyVKAhSR/jFX/BAM9crb3hcEQeb0rlEBTU6
A7gf1l71KK7xhLZy/d/KgAQ54PgRotM28ikMwyzL1y2tZ0Jr3lEIG+ITVKp431zb
u8sB2KJR29DgbijlxtIUiY5ky1aiXavur4W5PwNK2DixvLvDAy0cs6nFQXHeifEE
veVwC1yFbL/yWPUrlpVMHscT+VaoSvzh+fX2jjoZy+wFp5gjnhCEloRpNzgxzCMc
+DT5xZyyNt4508FfCqJ1pt6H7LlMZ7IfDqUx/8O5+4KVR/OxKktrWLE3HHRF9OL4
7PlQXyRge9W56FLlT9T8KhwU68TFL9NYYy/yTLkEKCK8DlOcEEf9JYqFijI7xUsk
9C63bbXHMsaWTjGP5whluhIu1zL/FMgVOf/aPhKhX1870kkCAjlC7s2y56Y44ZZX
+dePhMGg7NpUJJzbYc56QTIv4UC2gND5+crQvzc57c/BnthadFIi9nf6LIWVT/HR
W0S+OWTrqd+1mNRt1+xtqPhoYW5k2iWTebBaZQDyF+AM7efTYHg5JyZU49gNd8i7
JLWitZgKKcvB1mdW8rRDER+77lAFM6UQ/FS86eZn2FksZMTPykHFuO1CLmP9d6Wn
E+o2A2L0vaCS/C6BIA87SiVDAFsJqd+YUtdkYh7a9rAwDVh3Tei+d8nhBoCH43x2
B4jKVSSEzQ8G6cVEn/XG4tOvjSbXzg11nJCbS5DrPie/5n7JVVI0AZChf767J3RM
jXS8Wn3rGSc+lHskOK1uuWyWhFnKrCpOYQbShoafW1+F5YnKM7D9qdMpJAX5Tl8J
P3ZggO6qx/yDw5y5/fAAqaE7fefQUMNb8MYNvG+zfcKCiYHJAjLzxpE+VOQYPO4F
G7u69lyrPyd+UwEL1jFkvAgxjMvWLUHJZ5YcHpecdpRha+lYUcRKH5IApaqdSOEl
uFqC8yKQlleIQVsOPbhTQJWVcqG4FsXRvd7YjhboBICgdgX3JoYVtmnqrlHkO/4T
44qMcW4eTz+tIVUeS1vvnilnQDRzZ6v8GL6dTGeoT+El70HMeabdtQz8+cZVM8nD
lfKsZf5ZlssWymE6vxZp14T5BcPbUDnxoy3y6sHacY/IQ2uWK4sI+9UU3E47GdSV
ztVcqiNn/zvepw5nuDKn8VEkpvi8qQTv/vRquyNf8TgWNvznq7sQLPqXX6wSwOSI
aSWL/Hwt506LdxtVAqAE5e4p6KGTqReeqdMsuRp+Lo6EsvdcUzqpqtzw1YicSpbq
Dc9cfe2dQTKlz/jwFsZYhEDDRWb7poZInUa9jIrfTcPq1lHYuM5qd42O3Hdh7DX0
UEOSU5iHEkua9T8hofkJoNoQbQDpp7eLHtfpDYyTd5sGH0a69DSTcoS7/imuZjqy
iQyLnKOT6QtgnfUtPoFaOn2ezLO1oVxUZVM/lb5IV0znTCg6MDmbx4VLDYnwyeLx
NQpAVhqQwcUi0iHD7wsd69l/1T5y0kbARRbcxYVU2mTI18oyTo3ZmH47UNnFKgT1
IK2rYErUPIitwwb36J4aMDSNlHcdr4o02EMIbYSsG1XlQexOiHLnzx48gLxWXvsX
SyfYnIemjHsqW/AZSW+Lpti9HLHpBgtV0FNCkQfi6+MD+vEoDECjiWDYe8L6cWYE
Sb56CTnpJRfTp+6NS2rS8yxDW15oIVPsUUZbSaGe6SaWlju2deGvLhYYlbtbrOQI
dXGyosomviWQqXpHj5SPyX5MtRCExMJSet0gB4ItMil+3NOB1rZA+LYyrrFyeyWP
2cuIsE5RW5TXSIIcxaR7i7pA1/URa47PL1WiPUikBfLE2aXn9m4aO1xOKeFvcYcN
Zo06OhpxzQccmGbZEgn2d2BCj1QNkmf18NkjR1wa/k2BLL9RMt4eNqmG2fIRpXiB
0bEtyEmdEuLQWwnyofrsdMagyB6VGvczgDuQTv8gcdja74shKL2bU4JKnbAUJxGa
Q+tgSn6/2OLQT/VG23drmB3/TcIF1cGlF0O5vgrOAc2TdfcsJSpmDpsJFhjR7E78
ZZkEYZJpsmrIYeWHiGhtACcbzw+CTQkJHzW7sLlXVGTfDQgjj0AKAIlKiXexcora
RsHc80v6mwaWjJSGJssXS9bFwVRk8PC9XrRICo9XNJapoNboj90RXT0N8axy96lj
RRTqxvVnqCqJTvkByTgybWxwB1uvqmthj2bqyM1RfI5nhbbwkuEObcZU+GaeO/LP
2XwwYP0pFv9+LEKdYxdXUispfkTiE2fsSrx79O5MowGLucoU75x2EytaB+q4AVWH
xYjrOrUV4lK/rNv7HFh8BpLnOP0WrDH0RhDuW9owPT3SV85ZHIL8SZllxiA5rEAm
1cy+rQBl4Q9HDB9pZD+uFQ/+FY3x4Ari7BO5ZGcDP2K4NudtFh+q3Z4oJwQDgwRs
7kKCVqyHP8r2j+xGEDDTkBlnLEPFmcTGQQHCaoVdnosYKMpgsAXt35DkobFoRDsz
ojNCK3iMJJYIVz38LlXBNWeSSoX7BmGE3TjFU0J4BhC88+3Apc3a6K0rZv6YfwRV
OYoLkVRPTkBsHElpJLGCpwCMYPsk7eWSV7/YQkno6T8YumeMmcj2rI9A1HjjYlpZ
l50kT28+m5KWowGgKXP+ARHBc9wTJVYJq5PdJwsrkSfFpoGuPkL7NQeid2VRXQpF
DZsZORFMOidoHtcAuuOI0Rg3q7LsqzElX9NDdSqbl4wePHahhFniWu9R/yeuOvwB
msO+eJK9gQO54sZoMPWpuTNpgkDYRZq/Qbd8519H0SJFUrTjIBRFJWpKeZVwRL2v
wCGowOc8Li9Fldvs/bPNCygz5c6ZBqAZEp0jOFawYEjrEw5XUAftgZbO1gKdoZQ2
5U3KxYL/ag0nEixBfUeWXGry5lscOlHxqea8byvos/Ek6AQj1c7zOYwZsPP3rgPM
nO3xRgq+oW7e2UwsqcnbpPjM2VPROBfQ6/N3DXgxuQLhKFtBJHdybNESMJmACGkr
00kaOdJAqXyFVkiPfSslT5gUhJ5xSYhlFefXjO6vspyu1QULnyUzFKj5vB+e8lnJ
bJ5XhEu/eXpUld0+r7ZUiMzqiAH8XotkIZpadlZrrKoiEzFrP1xtUZ2dFMuUzdQR
cNkGq0PoXXMxX3FzHMQqSGmCNIpAMh8bP3iTL4NfcSGTWWH0sCxl2fsGspAFbd/o
rt2fN0HgspOk1PaFS1Qz4Dr36JmnyxBvKraq1kqlP8cH3TqkMblwDRDczhrCUWWX
/RwQ1KhOm9a0LOIcxNdMlZHb++wIC3WLWInJzN8REWo6Zcqkw4WJ7NgTvE9T0Kzn
sfrT0nRWXNNoTKv30X0RDjTMJfwE/PXnGMcMVyKJ3+3sBTa8+XDjRxgUdYWVobEe
kt6WBavJS/K26SHqL4J2d0boCJ3wsE4o3cYK+e1rijcrLfYdvKAgthery8hp6p9B
m/mM8jloQvpqvDhUnZ/6un4Msgv8NKNIZIWYReBFgeXr7H1MX2zX76+Ib8yRCx0F
ZZZGcFss2NHU5zW3kxEqxIjK4WLpjNyhpTv6OU3Y+tZY9tDD8MGEVMlPCrIzoxqo
BjpP0ta2wpD046btLag5lHeECCg1wkc2uvsS91JbKl4zNHMPbT9DTrvQzRMKVKJm
Ax+PbGgJ6jmHJP6E3TXuztAuaYX25M6E1G+p/Y9EKvlXNoyc0SnQOCsK9nfFtHfh
v1xxRn9Ozj/XHX/Ry51xl0lrvAjmOo7t1Dl/66BjRbD+9mPaT77fdioqwZHH6wX9
UzzV+Pl9b9wINfIBNSAgWiwPicJdLw9ukWwFHTteS7AAnHtkdk51SU1ivqVSjyaE
pKcqNarA67mCXVubCkEaBeMiVjM/2Z4f2jt16PeMmEXS6LRpd4TCQ46JIo5yukfi
h506LBfg0sthe9LLr+bf1c0rC0CsIAMjMWDqqNpNCwlav/UEL/PyqDSI1iL0YmbD
OXaJ/dUnjiPzqWo6z45Suz98RgF5N2DNxGmjdgAcbBnFrag/d1eOYvZlNJZvt60j
ZCYwQdAxfbS182xUB/Msow0ZL2Bnexv42YdEfZSNQjZlbqhCnN6KZz3RVNVK2HMX
i7pBEHpCc1g+ps4GjC5tERHramDBjmLzvXVoVg5sv0tmdTl5EZhC+SV97xSqUFsG
uvDJDX8Flgn2PNF+zdOQLDeWjRRSS750GR3jjmekwWYZbXb+Qcx9guCpP1BLknWj
Ol0GYLEYMG0AQZ5UCjWXAyOSx2Yjp2MscsU5NAHBdkH7a4GNbsawDhMztbXMrUnO
dKgJGfPsj6r3y6FvWKXqSyViNWNB1j2TxBwgQQTtTKQ9IMuy8Mc5T1ACw9+Aa7ih
RxgzGuDFPAsitqcG7CbizKNTQgFz3lzlH0PDmKJpFIUc6C3eE5mN7brYe9GJ9wOL
y61tkpQcRlPtDjoevuMwytJdeFDzRpa0MoOMDAiTZL91sgOQQN+W5I40yd9LMtL6
to65/40KZOCL/EzauWH2pr+Nx3nCfv4LPEd3S/la8ZAmf7xruTbUtD0Pj4grn7Xs
3vfdxtxSkboeQUnTSn6Ya34B7y1CiiToI1RLyW2NPV+EK7j/isCoD/G6LLzl0BhE
ec/LN5abdlKmbhkq+sax2MU/2f6QQ8zq1HuWictGsZ/X6XUHjWhloltGyZ6wGZib
0Tz2qabqmhdwCvF1nweRrFButY0fHrALen4JvnMb3ethPgiHRD6vyMudnC/cy2KQ
aQ+iia9UpwI9RGWPugUmvciGd83atoXiqN7RmO0O+2sn0bkB273mu55002ohaZJ/
jtcr76Gtlwbm/dFnKQD4X21xQjBgAHhVicIqbPMYFm61z/dnYES8XNsl4QhHgxhr
d6J6AtFN5WiPUGq8I/Cfa45FYei4gi+jjMddhcv35oZM9xnTqVQ8uP51jA52gleD
OeXsTu6yS6nSe649vguR31c7yMqVXw5AeGXg6V0gw7DC6VNiEg7nTQ8oyhvjDFSs
KngsmY0I/fw4JSQN7rtlmifcJtdGYVAScGNErP7nvI6F3HSFf6FkhAhDMxLzbofH
bCuWmZJNSupuO4dhMz1XykPtmL5dJLiawAGSStnh6dU+g6jZe/oMAyHM5EGMUJ9I
8q8aocqGiHg8geDX0ZcwvAfnM0/j6wd3Slu6o6o+aod6FI50Yd0bBMxfPnkkrIlv
2gLQ90kO7QUx8IRfPmFR5+EwfxM9wUXuu4BrkE66sPwu0qCgBxWItIsTrwFdaX/I
XshgricJXoFl2dI+NDGPf+hBY57/YlSOhUDCCI9anTS/eF1Bo8NHI3hhmTr0r5Ig
vaKEwDHchR33vRmErzPQjZlRpoQLtUxBAjxsQq/0fnhaR3iawgYgXK1uZydxzejV
EKmQ4eMWHG9/HR0ak1/SIRuZKZpLos2dWohEWRfl/PRfDiIAxKryeEhfrI0Z/u2x
5KSNIhNp4scIAowMqbAj3nZAE9INL6TOAjWpL9OQQN/hC6vi2ZA3dFhnVZSCaxVm
mhiHznD01mMVsa7BBk04pejpAg+KEezZEs0mu7/GahET1G96qtq7r/u8SAiPXaQr
JI0uOQPMWR9ZayUtM7ZTVSVIIW6BX3Pu8x1gYCRn7Y7IiLPaVvad80VzhkuPekpg
mw/B6HYn+bg6uInVv1lR2vjO+nzxNgcYw52RGKuAIdjvd34EAkkMvWBGiS3GJOqs
sA7KmC6X68fScNCu/kPBq2mnsZJ8fLhvyyHip7OM4U8ikjX3hWRxRFLQEvIo9e8B
KOgTCMic5EyAUNAdxsVCcll0VhupiEzOiiBjn5eWb+i6TKcmbZVX4m23v9RocHYf
gJd04+p/cref05FRU2Ydg8iPCcTMLNboLX+TWAR8mat5n57p+3GM2LlWBGsdmU85
2l3xRcj/oOC7ozWc3uujWpuHETTcCMjCz1cFsB8LagJKdg+/5w5vsrgbi3Oeuw+D
MZsuhzKYn1zGsSY6XOrbATbojApd5/3rmWLHWqs603t+hrLaExfP2uoYOSSX8uR2
41QQX+rZnNG1PVI89iyuHk5ore6+ck85PehEECJRcAvNt4tyaTZYOh+7bTmCTJSU
mDJUscJdpFNd7TO/Ap3ZXx4246pAvL/+cCEGuHhCVIoHHyAXeryXVkOczGGWbMs7
A4mn49S1GZkDLG8tD0ndK7bDptKC5AvTQZszYjKZ7tf9jT4wl9nYAt7uLb7+SztX
I27fPe7v+K/pHAW9Hr+2l1pqfP2eIz6XNnWE30YdcxU+Az1Edd01BBAlsdzXuWkC
qPrUPMULj/7YacJDU3TpcgvjJH83Ebbch/lnIektf0YHDRfbLHeveuK+JuUi9XDy
GJciJk65/AJ2u8PeSuaJ30miTr6SfSPf1qk7XxBR46YusNSGoQmFduSBL2zLetYP
qtNdTll+bnMWwa+cy4rAvivoeYj7cr7KPgkx/H32kIbzWwRu13Be2vgsRfEWRUFW
+aEiZUdeMr6YBxumrAg31PoZsoTOahRd55y/7g1nW/389e4P8ajzY3pMQUEKVohr
Wx5S4SfOzZB3JqWsGYZWPIKdosv5HkHrmh6IFly1GyxjrPCSjnwIE2E+p5ab74nr
0TkQWLAtNyR1PZfnBGE71qqGPcs+X44vG/xhAPPvZ9J5tQIESMoIFdx0JBk/zUJt
nua48NeVWaKaNOKuqEMSHiJIdqJHb57vLKVCC3BGfuykaXjiplhJoAGfyeOjG933
sKzkNKmGr2koG8FEn7kp9Tse+ERxALs5thX3ozCjSR7gN5PRt15glE49qBtiz0Yx
M1WA40dZF7cjUf04wUVWpAihhF2sB1+b4NFAEdrcb/o/PZY9m5orknIo3QYPWDy0
2xofio53wlDq2sx+utoqXp6FVVmeB3/3Bz9jRBDkjO/vZLQVkj/OjDxcx2C/cj3Z
DABS1kY7gmdFOhoREXNCmvH3+EPGvfveRY//Mxi0EwRZYqIKiVy2U+ZrALDtxSH0
xqeWsgF+NbwvvuHTwK7Q8DHwz6DRXK74U2dSBlriPr2vKxejflgF8M0xOl4WkDd8
eo87EyabX4TnVaBF4Gx7Cq1cOpaBP+8Fod4Cde46nuwdzLioCnzRYSYnHqp3TbVp
3izU2AFCOUhaBRHkF4G4089bypwe8cptHfyhWazSBgg4F1I+RIJC3pQLBVIChC0W
jh5cTIqm2iBCgjIb88SkFb6pxGALufrwVkHDErjzWBRj1itKtqenAi7wc3YU293o
NkxB/IsbZbCyffumMuQC2GYFtyRhEfsJor2yI3ayCa5KusaoPHEapr/adcaVIAcW
Bwc2iQh+aHodKhUxnaDTfdB3It/5Ifqgz4zgYxuGTgGDEu6sBAuCrlmUgUt7WOgW
NhRKfK94TARkYi+a/k+xvXS2JnC+7CgtETOZEF9AWO0+VFF1EgYe9dMVZIh+KI2m
Q1Wed/oaZiRlfwhkIEFIJJbjEsLs7Z+1LCquX/1yylk=
`protect end_protected