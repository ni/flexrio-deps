`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
gMcHP74wBZczB0bB0IzoP2xg5wC5NPjD/GsvSQ6VQgzYAsanETMwwsWi4yhFtJwv
5kY07u0WerSDf8woJ0stqW5xF501W3JLIS8KMiCOd55RHBOnavjYiaaLeu7oUCmB
TtTS1R4sO325rP2zOn9YwRbyyS5Ljn+PzFZZUmkt5xMca3p5NGqKtZW2dV6Babni
5HlLuF20Au601B75m2nv+ZRoGSrpkNElxoTibONmX8gBflpIVE7BehhHwaKSucEF
pp4QQ5zZAZjEC6aplZepouGVggAulz5AahlX5bf4opOVlB1J7IrgyjENtw6ysQ/q
DzybQ+ipztSXBGhmcCVU3A==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="jAI3OJE9Sh00Sic4PtM/KZ4WjwT98XM8AMZrZsQkxWQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hyw9IrFLPQsjvXplweG8O0lkaSLBN9Ijv4B5VdTRt6ipKJT9Kzsb5LxCKvkQyF9n
sGPOd5i74hRHnkHfYISGkfxGJCa55ieOyFShOsqTKRLxclm4oja9vTIey6yFm1BZ
54IDCG9h3PqfDiTD847UCSMRvFssyycwv+BRHQMQlFs=
`protect rights_digest_method = "sha256"
`protect end_toolblock="BnLuc3jxknmZOyxfJK70E5kp9u9O8IQ8cgkXv26kHA8="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24224 )
`protect data_block
xABArkLxBOK6xG+7CdOOiGu0zbCbHMrEntFfAZEE/xRFxZaAZl1QLkuFI77OC2KL
XxG/mrHJzO3taVHgwRXNLDdc8ePbxbAiQfzV3NJLBO+gsBjmIymaCa480cPNpHLx
0+LIRl85m3WFWTFxk3QeDeQJIb0wcjsyJ/NPQgTdGXn31ZmUqfbsEVs2e0AXm041
Ax27u/3QD2lMGpRM8w80YUMAjN5Zv76o/SKGYAoUJPBbqhaMHK7sjGh/rXMvCARQ
oVjZlvw8nkgKvTcxhwSyQBFFoXskpE7heglKX3yhq/ESZM+DV90vDhloJn6heeoY
dOY5TFUnMSL7pCBGZbWd5jlXewCJYL/Zt8EbsRwMIFKm+zmuYSVCdOnZrqBP6tr5
SrzRm4pxtmIGKW+5sTCV58oFqhZXeHhhDKhXuAwqUWo86wYKtwIyju06qQSETqjP
ykpLM8SsLwioY3qrXkouORsLMrozNQlVIuvU9h1qhMeWs+djb5PYA9+lkLxeg7Gu
5P1zoYqh0VC5M00cxJ90jFOgW9ntwEFG0aOlayuIfjJl0QFTE5yjjqRSYEGo9yrg
URjvYEuAXwHGVZi8jk10JPGGhOK7Mnyj/mMBeCyx/n0mhgCOd+L51EqExIfmcRkz
NOwKLChoivQnuVkc1wusKvWxcIaMbcQFXkPtfP+88nJ1B6/nbRTgPgbssLi47W2a
9Pr1I+aIXiMOlBi1B3ESFF+O7vsYgZzRC7zLAT08Z9T4ew3c0GtSz++VOGX4cTxb
Td9vXVWo1kTkMJPojpBbKp42Yo7UKE3L75a92e87oQvYmhuC1HhkukYC/BZWhsM8
1qRVxueZX5yVqHVWJ17sFvLkO8mhgehLiyk8gvVm8S9yrkjqO52/f1CIgXm8ie+z
rivVaUvQzmhDH73cCi3LI6keJkn3Boo5LIyFjI4Tn1i8NLxYyWqVmbsFdPaiq/Dn
ISQuHrLHhVH82otjsAX0jnhovlR7c8fD6tK7zSsja0H5d0roPVtT6rZXoIRxjBYN
HUKTAictSIb3qilR18W3CyguDC8Cg4T0PVMFgnT9Ca2CrvR7htyLtf6SJKK68QUX
IJNq5uPbqa2IscDB2eX09EbTEbf4/ZEtOprB8hYu3z/27ZJvzk7s1a4Gc4u1Qxw0
+sfdSIRL7PpOnHBpuH9f6MgOV2djnnGgbuj6JJw4OSnMlsO/9V3j6pznw7M3m7sG
sybpNr2lrkDs+V1TPp0B+CL0yGJfqtWaAc5Z14K9qZWlhYMvPPL0yPg7awTDC9M/
uuuhtZEiTCRRRlT3Pn9gZ6Rswrh8kg8W1rgqJeOt4XKxeDYot68UUZ9prpatK8w6
gVIgRRET5G8tnWIxMT4duePYt8XjhuJGW/OGNoiDx6xQdBVYbLY0rSnikMpuF61k
U8pNY3mqUv8Cha2ICKi52R2oi+2eZc0IHRxscC+vVFDrpGhgypC148vRhlC2vZiF
yvre+jABqWNYXeQ7zhVCBc/vpEJgp333nyJdvIh2DC8XlC1CBk8ckz/0ZumLYYiB
QeqlEEgMaHDgJ3gP3a2n76YeBy0Nqk1q/4AliTBcpzByay2CHgaXwJ1ETy4HIBEf
kxJkNPljUbfoauIBtjXsufX+gvacSLhQ1SByCDPi0UGFeMDSYRg+svze8omsSWlR
7WDltWjEOjRaL9310kh35qOy85x2ybNLuswDb2Vm+Zj7W4niw/SpRPWR81GZBG10
lFG/RasdbR98+SgFBBGmVE7rYS26mPTXRvpVxdEdAFQDG/hmkKEZGYggeYqXag3E
XK3px0WQINsZjf7el7210HyseSsmRxSQmr4LqK9EGYENY+Xg5YX2yV9XZQ5/2rWV
SwLNvwWfrMN3F2b9qiPz1j63IfVCan1UgAA48Drn9WfB36z6kOXdFuH95lWRf1vz
ydLjnH3rExrOOeDEeupX5VY47b1/1unBX+QIV0IK2AF9zToxrMm4Z0t2tPA/j0AT
pMXSVyEpOtOPBK9fjOXf4BaWp5wxVwifpB+dgsokZE3t5z1oODO3mFg4yTCmAowx
l3N+V4gkynDIkvqIvsT8liqYL0YedipMDzCUqjOP5w6VE9r+EQXCeAqcLkDCsDda
dAlR6TIIsPb7Jm1MJUCWZKBYXieDleVu12CDfo6OL3Z5udMjw+e5LTq9eX8gj16/
Tdd0SKuqC5dGoiu9IEyzLza90tXstKxaRu0QHPNNMA2JxX68+JNrjuHaCyK+yL+i
HdBenpex8Qs6nCa4Wg1XG5WKgiB/V4q1yzkXzcYD+ReXC+RyTDDZgoFoA4Oi+zDe
iuAyFmtEjwsYv58w6hvwL2csA6puTxt6GwEucGjh4giPjJ/cInZWJBKZVJKuvFPm
dC55o5pbquGEzvOKEpnk6wAisA0SS8CzJn7ohnmux8oTu2dt765FSQ8LGLiZOERC
AFYefs6qlpW7NZ5A7aJakATvWjreHN53YhIi/wVr3pMMkBNk889xZ+k8RyvLZmcf
nwm9NNiZaC0GMv/MQsaslpBpeLXtRHczncNEdXNccl7e1GAXosUqckz/H1PitbRy
qCKiTJYFAmR4AOPrqFIuXRbHOoguHd1eozNiERkpgDBtR6P8JDqvvOJe+3K5Ul7j
M9t0mK3UxnHqwsM9S2cObiBDEqyUqYRIAbyGmRaxTYSnMsVxkOYxWQ8EcCIh2lLH
9uCaRhety6Bgd4C9ABfQucyR4vTUyBdqjE6+l4Mnw7/B6kLoAVb4Q7cbRXoH5ibA
nC2om6WcCXeZ/3E71+UeknGGiqsxfHLMXc/gvLjlWNC1RMFSUaBQgL4qzGKIYScs
p627yI9EnGKXIHsLRHxAHQSwJ4ZYRjKWN7RJjPv41LBeucAo481qAj0wOAcI0kb2
vOUHcta6xnDzOXqYlZ8hcmIKvf2HuVUealAbGR2KB2gM9EFOFVfGv88MW/3Haonx
yyv1FapocMuVQIMQ8JXDpMekglIpAE+yxmicqxgGc/T9UvdVytSS+rafdzY2Uxtq
FOBuyxrxBv0uWOuZP67Sz4yfSW+V2mxUJAxiliCBdpChmItIu3SYhwsqOIdVNUiF
IZ/lyzM3u9p490R9ffDir4Egu8QdWopaqoL2aR0+A7Hnh3OsZJnQ1kUViwVxU3FG
tP3EQizXZviFt8Z/7GVQvlj4TCOQIRjxIikRCcuNzXCWzzAISf53nG6UgerVbHQh
GqX/aweT9l4Ym/XEL9JxuHfuJvh/mhQPPciO1jDo/fOKQophltCgCotEFpR7tzzF
tuOxIh5C6QGj75nDNfS8kM11lNeCJNVcuJ0FyH2w1ln3y5VC9SCYBvgudtj8RK4y
i5IreKUeMEdsJIEfZW+gwOdyotr8/KZYhdHOhvpy/SCNpRNZvHmhulV1HtL7H5MQ
5N0V78EUImspLa3VP5nN4+Y4hkXhAFVP9AkpxoC2Dqg/5HJc/25aH1DldCYpi5jC
C3dewPUc4uSiMP59VvpzubgGBN3LrmJOmLfssgVzG4K/wxbgzrxZjjW7Tp6u2skS
y9mB2+zUdYcZcHjkIXbh2FUx6Kq4lYaoc7fl2rmlSbY4NJ++ei4UyLcbk4XtqalW
/XsPeCe7CuWvE7GzGSdJQm757+3azf9l6Lr9vikS6SK2oXH1x9y/ONnqtYgWFMMW
FDQQ5PCtCmpQ4pXTX4jnSQ2MPlSom36rvcmuUzZxDo3Hs5PoPEMTU3FR/YXZbNuB
sOFOyX6HC0k6ZuKAn+xDGY+kZCBKmBV+jEpZaIaa0Cx/gL74TPrHYqaMjmBqQg9w
eVwLqns+NqCyfpYrimklvlAvOyljB1NLpCYz9jZMNqHnYnnALK1Te8jQ8bnTlhWf
UZtKa8shMfwI3t63ojU9YfvgcUP6SQt3ZUYj8RKMexRAbTY9wBGof8HQiAh1o89X
7AsMX1G+QGvG7RZYvD6g2BzJ0+4kTUIq5XC/DJrLjndNh8+oj4BDGtece1iBss4Q
YNTYp0hgTzKMS/fKTDPNfQXvoVZqR8VTSjkHsrCsLXX/B2kxl2A50VFvqpU2aF6H
uXrqKlJhVbct7/neSbD4oZZJtyoPspEJpo//rBEwVzFftkBxjBkD17cA5rZVqAaB
bVN42pcQHeBpv8S3cdztvN+Oowmbl38D88q3quUrp1ZzS3AX1rzJr9KDcILp6OVa
kcYeOHePUL7MNxelKFX+AMyU99VQu3Fg+Cw1tRfp9KOTNUHJhUwpqeSAomKt3iYm
jE0RAoJ9Hn6VPQusbNbDyVUQpDAkj7kyISGKDenQ5ESNjHxIMB1xMtabHFh5Sdwo
x6v2CoVJw2/EjR02lihneUJrHC7bsK1FPknoIDpdtWMvea77zO6gAverSneytNHS
b4uua6HuncmBQLHzo6AbnOwabp1JMLkFaldgcJVwOH2kWjUFhaMFYS5J2zMrnHSu
48mOmGQpSnbQc25oct/3tTTBx1GPgEMXnubUNHPl4CzBmkEfFIkkIbBrj3iNAsNd
YqhloGZZ+GZaq1smB6aem88N/OmI2/5YUeCsXhcYA36T435ImfM1i4U5GuwDg85P
vdtDorPlyzCjTmpGkb0XWQvO+XPQxUH5NdSJz4QAOTrUD/Zgfb9oGsFjjL//yKo7
8IoDoWk26uX6IjGgJSrjPXSbsziOa0PhlEjhpB2YyBSUh+/rNct4bmv1ySOXakt7
M3Qdt2rR6aE/7jEbyiKAPWvzB7mjBNrGiLh2kT1PI7T05GtSo/iUAg+3zCndjGEQ
EmQ7g8qiwOc+5AHkDshplDN5J5qhhiathMVdPDg5fH5bDXKQSpgWNAWBUHk2mSAJ
2Cn1CoJgiSEfHn0lSoV2WMo9MVogZ5F4/8kNnjb++CViGo7J7MRvFnGt5XuRzsfh
VJz8cRUESbkh+u7tKTttopdEqqWBLKsR3GKhMfKj8uKq50s9npTRnSq1Ugt5tQcf
9tVuhML0P5KaGzS4ONsLQw+l9Fc6wmXYeSW2tCwtFbT3aEC2X1hjn9JAcvFK+sij
nKkEMpuzO7e6eELKK5AwneuzDtu9jyroFg6uj5dWI5roWhoEBA1GtqrxHb5DOZNi
/virT1MzhzWvysn++9xlWcvdLHTZ45ywUC6kuqmiAvHnnFGCy+LIeuY7dXqkpjVo
VjR34jfb5vDNSjLtepFNS7B7DCgcBzaG2vD4IdMY4atDUwdjNOnqJiJrWitdVOsC
BXRlUWxWatNT3ZAfdSHI0Fdj6Kj6BpQwwOeQ0GCAD/+1DxX8ZJIZ8a9zvsZxeuAx
Obnn8a1NM5BTg42T1uAN9HPhhN37K61LqgNqPHlguLjlAr78M0NieaNHmbi9YJ/G
kLv2RD3HPYLEHS+QS+LjY2lWUg9EGzvaDc31YvGv/cekPRM7NJpqSEEE5TAYJc86
21arcWsrMmVRVJWR9vJKSpeP+idn11p2rHxGWHCgTG3aWH50hTdaCaY+7Buw9HWo
o3BZwlkWnfj4/oTBOiv7Nj8lzTOnDU0CQQ8HZDptZFGP0O4AoArF5KsBqznzSPKr
yKCS+/J3Nlds77gnd+4XATzM0A1LDrjPM+cvYY5BGpabfOi/A8p/gvoDrjZruttd
umQLs1el91eaKsQ1HkvVk7BlPOpwLa82MB+mkTegigY7zN7ue4+CT1HcFMifXcxu
NwQomJLrUpkdE69G9OsLkmf1MEJUO+qHC5RfdY7Yt0bVRNHef/dwqvbmWlzhmx/L
d9ljmuh5Q/+TQgFehg66byEXBryS56RZhUtBxg4AcSvnOEzsBXxc5ClTvKSl9lBs
MGeZWox8rEqxMHAX16U/k5KQ2IJ+eoCssjokCYSK/e8bamK6BKX9mkKCaFiiTYMz
VdmVJm0TfgdFpdR6/sCCfkXU2NuQL91LTOFn+wvf8p0DnWFCWhBiLsAqPSXpN8JZ
sqjCh6IAUUagvOCneGRFSl2gaXHTVmKIrwefz8pF84aHaii6masrvUJK0gS20vfj
F6lv02cGN8BGwEk4NjbjTrZt/pqImBcPRWqgthdZQ+og1xClO2vr6R5CMKpAASKz
JJtsxUowAFFM7rFWIkugoomGrCFHCuX2yP2ctriDST7JTjf3CEnPQ1hGFXyyhkq3
v1MiHe5Ji8z8lVjy9zSl4N3GDeP0vM4Mm759DZL3OJ//+ZB+Btvr07Daduwy4qQX
le8ajjrJK6tTlSCQY/RYN5c61r6Vgq5uFqOUCBqfVPUQ7cr/CaPOC9pXN7mKUMVA
wdvhM3lzli249bQ2YdJ4BKiot2PmsmhkrxPhchPTuIyfYwJ6OtMD7IAFEO69DTuQ
HwVIw75NSR7D8ZZzZ7DRZtL4Focf/t1qFARbI9Sc4Kkejeg3Hh7rBtb8TYSVWUW/
pnGLatuQwEwfNNnwEDR6n6m3se3JR1qWE0Cbl8uxyzDSdRE06gqDT+K3fU8A9gNj
n5sU/viOpGynfGs2OLZvxpoVXyzxU11P4R90XKT2Cf+cw2LZqwWHdmMUtr10HLoz
N4J+XpjzuSyN/orOQsXBn9hL+OHkMq9lhzqDkeiqbZysclHlX1u0bO77wxBmaG3m
t0IOHxlMP2X6v3AFkXIWna7K0/sNHjupojAEpYm/MuQheby+Qg9drPOmJs5u6BHa
N2vMyQzUl78cwIXwl2yyvdyPqd4ECuwm3Qz6EmAZ0supl+P3/jfKhG/YWPnixDwv
tkyRbs2Vtnb2YFQjrQsR0RkeidWsC2bUrDbiOaNvm2UmuDMAcU+JGXn+dTnWNZrk
WLQF3UxfT7lvElQ//dccVqTNY5VupqEPBgHTTA1ukVm1GBeOISxO85kNrQvFIlgO
OhrDhAgMb4I4NQR+g7FzG7OKz4Itd8V4J7NYJGFiC/U/v1PCUrk52vss2rb3Xd0I
ZWuInGoMbFGxlhIq2XL5yfvJhFXRCH9MOjXWvZKqZsWCOOKNWXBHMBTtwEjo8hiF
P/99bdxC31pH1e0c1G34ADejajFOAgakA7L5MO3sAzcr6xe86GbqdbK1QU8Jp2cP
utEbnUq9akRXKsn7F0MEzMw4+SJKaJQUtRJbUXmHcpBg8eHLlxnyuoZ+mgJt5vnO
QNBaYzzN5YGGr3N1dn5CLgkL4BoKlAQEthBPJmqQVq3+Cv4rRNCiASO1UDQwRyXu
V2qfcNkQjQQsqWtZwkgTnCc3RQpwdzj9Fua0pUHLmmvV2hjreg6buyoHjEhGetYH
F6aXqNAIth9gTEp4mcJ+QHp5Kp2SkLarsSwNyCzFu6ITNIGMu0iNFuurL+Wlax8L
ERYvIq7vFS+bq7dXFNqMwrQ23VMtkpzC0VFaroQJxjAfmyh3lHGUDuJj5OOLQtRV
WqaEYBcx7n2wdbFp+gi4OMx/EDNThrXwQ0UUA3cqrs1097GhWuOh3WHP77Dj4MGD
f9t7SwH7ES8r+ty8VyCMb0rA7BSswSXbbnCT5YBc2xDtXQt66wMdkkJn52OdKFaR
qtUR94xSvBd82srpHtX1n9x3msnRITsSgaFRhJxKXhaMPSpLafeyMPnYlvVatEIE
tTzkdsWeaK4siMKWoG5VLapg94Q3b8wyH/tZqXhNvaMnMaUtYG4fsrESWLhnFpTq
5QF/eVydy7L7upJAko9UawweafmSSuUYps6nCyXNGPFksLSnYk4hWIxbG4mNbsfy
PRtKdL1LM+pN5wnNuDKMCdR/+xgNvl1IaiRr8DmPY+PfeFQ5iEetdYETD9vRsJFS
KTmzbw9ICqxnR1Er2IE4JbbUmkfvm1uSMTioUMGipbg+WWLxA+/dpNqCql5cYsXr
r/bzVAER61OgitrVIYKkCU3l6h15UyXm2b5bzXqTi+bddJ0hsoplvztRXekV0Ii5
YMce7sgnHvgxQbL8gMDE13w5Mpt0GqdDil1A2jE0FBeJzWcECWz++bvUnPWCCFHQ
BWXcl8IfL9KYmehUZYRFXRLtrLFNT6nLTI5jAWPYt/eDUgxQhLtkZVzkrcTOqQnb
KM++Z1+cyhdGofYuPpme4dmddt5dT0fiMYS3F2K/QtxPkK0gATM6m6yGllYvsTHx
7zUYTipz2xHqjUp5bH0WufDIQkh9Ii+omc+tJH0nCE7y2ZSHS6xcwsjG8/6aN2YG
hYMpILC5kBtGD0MY6Nc+AhYGhaeaUOgkWW1CHCyHCII/ZriyBFPHVyvhbQaFTTmO
SED+awf+bliZOD/NJF+5bwP1CZRnSyqaTlIY4t7S/wpgjyIg9PKoPDdCOxmUZvpq
6Obsvrh+KNKiCK41tYzmTdh/qG8LntGQk5wZa9J6jBvLyBuIzi4Pc+cCHQFhwg6O
Zie5Bj9bFYq0EPi06v4ZAhSy6AoWtaEQZtVtxWFj9S1U+GLGQFdcXRLs1qxGvf6t
xjMVInAoDjF1AHT9IECklDG+tnMT/P68H/TZq0NEMolHF3+K3MrTklErr1h7ssd6
CPthh/P0yDnYc+xDArHFreOBsl/gvEf1qBdgceJXdVf5wMIRzPti4acWtpZq2U4f
3+dfd9E9Li7LDBmPSP0SUWHr/UIjUPjDQpmYPNjr3vD68+PTIU+QPMn6MyLrNJ/X
eJ8GCEfBkifc9gc0zKU7DYmMdQNy9DV4K3b5IWTu0p6/PKETaCBT6gCP7M4gQyNW
L/Xbeg277Vk5T15W/EVBFFazPdtQaDEMuq2WqbfZsCMJroJT5AL035rKNslHRlsl
ZOXwWlhPwN0FCXHmRicJhQcJx8xO4RAMYjERiRQxpmDe/CPDZyeAQq+0Ma60R/Cp
jSgQ7x/Pzu4ou99fxVlvkjKQyued6nqnE/EXfAvfSM7K4nQDJXXsSgOnoDRsXUT6
s1ywcHtEdVO44n113EqdCVuw4IlFNqcHQJFEatuzYvmNwlNkW62IiudCBUcZRXzw
AVz0iX9zzQIAmGlxLVj1Q/E+BQ0CMXa3GRPRjDctOA0t7vHLDFIA7z50Pod/dlpc
TossY5ZLAOTlCjGyYnft+neyk7Lu521qy9GbzUCkf6kCCJ67FeEyEnV/E2litRD1
q2xrWXeylh25Lxrao3N2VkZVPfT3rHaNWHPGQnBJGj6l1AfEm2ADxsGdc07Y57UD
keP3VNNuUoWV4XO8hjO3tn2aMYoQh3E88HCwML2wu0YkwIlvvbGYDArAKKFmzScV
uNcZMbNwnLK94G5EOAkw6KV+NAOZ0yxO12m5tAoK7vAOBEARPdN8MxZKQOp2Tnh1
nPRP1nuvEFetw++NQiTkRXilWmbBevaDKPrlgfeUJlUEBgbb6/2591ojjAPQMVYI
b257ZpqrLqHodR7PwIwa8oxUDQfxlnU2lVrbVGZaZjvSG2U7ZzqZFZVq+FTjAL6w
dcU7XImTVssSXz73gJBz9v+WbBlwvjF506T88+prdiuzG6cqok4IYNVYSj+MisI6
1SKT8N6HnuI9RV2eWcKsH5//uwILguEKb80iR2UEL+F/pFEeLTURAcC/jMml/OZN
R/acydQDPniugY96Z/OMWSfdbCVfv+lnSQ6WZqVDADIBQNUPvX6eHbP19c57r82D
3yrCcfa0vCdv2e8SqS1RCjc+Ml1O90wAbMU5Y7MyBaf64Z7pTf4dqA6z2L7HXRyk
w5SUDaRbBfQbEvOSR5wex20dYAccvL5jDBRYFEtBSahyaDcr1KIsW+KC5UPgj03m
EUdiCzyf/jGuk673GqQXPv78qjQKkXb8BBIeSEkI4sY/aFawxvBiH9vCfBaXM77d
XNad2cNPzTsIPcHzyoN5+83s93qYAMVDqlmY1Zh2k+GHLY9uA9OvFUAIlMGuOXP8
0fZzBhDLhRMbZ9pOXdOVH5OOKlW4sdbzmSA4nUngStmnmvdG1c9vH/QnkgxPXgea
L1S6zMx1zWE8KugTS48dyT56B0I2oon6Wq3K28tK1YVev8pP/etmyhS9gUEH+w/e
ZI0AmiJgxDC31FhK1lwEIXMb+UGRlFWdSDQfV7giYxUXiTPxEE1KnvjzFUzYA43L
pAgVPSLXWjJAQ1w05KtchJxvqysuxV+GO3oAnccB0qH7qaHX2tQloItAqq67AzHr
SrJ1GLhtmp0n0OMoLaXwEI5N1jK+Oq+1okCx4U8i2q71N4DXUE/ox+Amx6Iq0mds
32gQt3bQNWe6nyUhpaVxMO02s3Qx6Io03BorJxx4mU1H8djM9wFy6Y6mpCvgpIHW
HdERcTW2I2mAC1H47FAOqJ6aovi8dvnhHwoGfQth6O6ydoudna4MEr+5sQX4pEvw
Z704Qgfz+JWe7FI1azKe9K/oGKefnV+GKBqz7Avd4ilJ0rznwXzxa8K634yf0hJs
L3UweIxAzGTg9CkpWFTXA3+0lJw+V4R/efFi6YxjTdHFdGQfAk0P6ximG5fTy2F2
J68BW6wYKCWLkWPBuoolgzPQ9AdvhPRUW3kyEwO/Y04/QbNYoBAKpQ3U40OgAKxT
uWnnHt18RgaL2PzHLny2p8gC6sMulGwDz7yIK/so7qvFgA+pkj3AAGzgBwGGkaHZ
dNDpMHPb3k3wK8gCdK5KSk7jhJtRGYZscEXUVwYSdxGBLbXe7eRL/pU9ZU0x6trp
qLmiOAB3co+DZ/qLoQxGfJPIM1nD8R2yxhP8yh9sx8RtuBjLO4CmAFecISqy/2NT
DTvJxVU5qU/AMI7r2VPx7enUbkqEw6mMgNEt9JQlDBn5Jrkxg/L+/A/ZdDlpEsoG
S1IEyUDE7nvZFBG3qeDx+JAYWhSVMwdNXxsZT7p4+TsHFBeZCX7j2MeHPM+oSm7H
R2YM2jEAf+7RhM6M6htrgF32lLDdvAVKgeeeaZGHm/aBQT4Td2jEgNifWfz8MhGF
fIXAGJ5WwVB0FT9uPbne0v4TwKw8Mz+48zVQC/MLYXhC488TaGuyQiOtE1TcLBPV
PxalEVuWyMnDi+R8x/FtlVLAdeUCTUo56QTpsgICTm+kqV2F8U+5TNzkIuEAdU3T
zVEuI6F2qgIhOF5YxMpz4rIrWS+yfiMLlZdrrx3IeFuJma9sNRWIazdR8hM32rkn
mvEqD7HvZn1gO0Srww00hZPk+mDkaSlYFp65+HbrObQqZiJHPCs9groHvF76KIWi
0hpjOShaU/fmVgTy0lK21om1BhcXC1i6EVL4HWe3clWTVGRqd20KOkeG2mR92j3i
3zjHiE/+QErc3b6Jtn1TU3lR51t3IdgV/G4NiiCIQqDxYCFCPWGHcER9R0lifeNA
g+1uuVBZlwCSTUv6I253ul1sZXkraI1kuItTDFbBQ0X5/ozbOlVCQDz1bz0wLBSo
EjqSVQMV9xiAWJ6ZJA78USaMyNZ6LBKazbyQUplhBZiMD8JFNJQKCJS1UJmWm2oe
uM5PzB4ir1NDh+cXdb4klSCKgX0e11vF8+u5ClvSkkhaeuk1VkbM2egRzQrpV16n
HVqun63oVpoeKQYlYkEKKxC+WETGiINecSMA/WZfW7FAOy2bR42rNVimJm4s1jJL
dV+wY4TzOhP/GqiKeGpcNjWfrHJJccvZoGVu9GLsqW+W/UwZ/KxE2KQ74s8q77Cr
aQlPmhjCe37b1FiV07JZ7sLFjU7F0RxIP2Ld5vze7swBPgw8EmZuTygcO82nfcrZ
CAg907LS8K74SIpUJbHS/9BlQC/kMBgHpyaMKmAsIIncD89YzCA38yCivFgsGV69
Om7PuJXsHJAIwUX2Nk53sJgAf+Put/De4kCk7GnEqEIKop7+TTuc57IYJ7OjA6nG
8HUkrpCsTZhy3jQ7G0if/sqJL9esIbPNMjiMLzmKa1VOyYgYS4voEear0k+8FhWY
2sk3gXnQCILY5j8HWdSeP0huuQ6Il7zGTZNzZhsRm3mSINQSUPqRb2nbf645X3Q2
zI/LUMocK8bIGbRReLPceI++wuorBDz9QWoqh3VCi+Ywf6+vZYy6FzGk1N4kJQLQ
as0w71yo8sfvctyDiTGfukJInpeGOq41VgHPPuCIrz9g6bEkS4SUrwB3I+B9l76/
q4ruFCkOC4w4BuQyw7WXdh1V3Ik/sW88w1tUCR4qAi2Xk1sIuIT/sNpHJImF8T7L
X6zb6GHGoddpW/3vCUlL3ke+V5uwbzq5vou36mlYT7iatFpqf2/jN5cv+QMByvo3
3dvtNmF62YDrL9YUVZfg0dXIKpkyK4dp9Xxq+zn6H4a3MSnkMgsh7u8QNxabaVSU
DuMYFwVjDyMCc88oCxwGbv6zKeoUvfac9XwTqD2AnKj+yV85775Gg9qbK353Ezea
nI0lGsS12uO3G+mSO0iBJaJujVLra7Xbcz+QdJlV+W4ZgMjGnmKh2u4tYDA+mqAQ
EA/wxDg1ia/3UExTSs4PWJQ5ZeT67xTQyVX7P0KJpRp1UpXaiofJF/+K3VFl/sMg
fQDB3HBnDafrvkHbEFij51SzXkKLrMgZQ3NOr7GXWq3WmqOy9cJl8v0/MHujoGzS
ZnI3PdxfLdWNPlJyza4nIs4TNsFLgGnGnprp14AIsK1Eph6cPcN6V04bMPJcEd8+
mWD1LwUFKwsTNtkZY0NbBjvHGK3etP67DNPrLV8WfCgnmktf4aE87JOkwHvZP3aq
akJ11sdcqWjPdRAbTXrAGjotZFj14xft+z0ovzOcB7IkAi6OgKEBzfvnNYJwGIAv
UP3rZ8jNIcj092I6N3YhG4BXIGxhPIxtwTU0D55v3/CtjbDWXRenhr1cFjkj3UjW
KqJz5zWar79huT5zZIGXEK/aaZc3tYH13HLw2dnQgA3v4HXmn4y4hcK6AmWWOVpp
4SBZ1zqGrkGB/AS7YkzjH63Wqca3j69qAzZ32C9aHvn/8srkBT9vTSwlJBfgNOGS
NiQKGvfjimWt3fzaLvVgzJ3HBfvO2oO539p63OnzYIDfvJneTyXdADXPU/UxTlQf
Sdw4XfdeG+yGeu65nus6n0Z7ZKXKn6bb09z2BEvMl6+3GEDxCrp7m14oxif6mPt/
EXLdRMeOZF+WZ+coWW+1uQjkRmwNzYAaPUNPH3uLIo2I1lpebxU31Yh4l3Pp2QAf
zIuQqKb7x92BKZlFK0jISeQ7oM4GVRFkvKecDr+fSiTYKm2JjPPPNPtsyXOm0ZfI
Ph6izKdr0dtunQLmACTOYWOp0MRHdV4lHK7W2iM5C/I2Ufvq2fsL5xNB7vuYikbN
Vg6v6Ld0W4FLEn7uJwNLxQp2tJnaqOYBZH3E+3EOVJ+NVdkQutodagsw7mCsY/7o
EM69sdOv96KXnPdeAt9QwCTT2y8mqHpBhweEBVERhKB/eH9LI8lLLpL4SW6POHkR
b8ohg59W/X7SbUUXYvor+AQjgaxPZEFaM5LqDdmRFHQIMHJqFWhkjw+GdhRWYs1Q
HfeodcSfQbspgKL8BCz3kHSi43Pr3DW+Dbhk0KN1sgPmZqnUQdAGK9JrArMGI9TM
U16i67xgeCTb2sB6DWHbveBs0Hm4vUYDMBaWG4vSeHa+ZY98BiuwU7AOkk15jopB
hSGjQB0FlnklRBKNxG4BBPA+zyVNe4g8G2ybLhASzRg8SxLIAMDumYIkGgz9sQNp
2Qiv9+sfsaWtm0cb2CZ0JSErdT7OT040YoLEQf3lew3u88ps4FnXmfK4N75fm6hW
EKSrjytrqXShVx79BDAESSQ9bfpNw2SpWYXxZvOFUsvuxIXPdEAoDCrHCsICwhgO
455wEmyqW29rgkxyQ+D9C8B04vb+0AVmUsbka9XbSlTsn9KXmdg4a1SrH0XhWOvJ
81g4s7wSQwmUU+EmfWQOYb/iI7V4w2gJclajEesrybG8ttfwYAHjwVcWc3pUriOG
i+FkL+EzBPSWtmUAePLxIVZoLD5dvFveqUhgY4C1GhzHjJ/R3cJkNqEU81qIutX4
Nsy/t87P3ffTqrYtgnYkDLJz2KSlbD4BpACvvmwG/ZvLTJ1hbyCdu+4mXuU//zIG
OiromUQaJoCog9iIzPqAoBZ63xGpWcYmORBZtt4yVPXM2uU96OdVDfdSH/Dx9aMB
7l6i1xQW1Jf7H9854QWBlR7hYHbEd4xAsXMa52gjuYjcCmRA0/rxObb3asWgh2Hi
I6y4JL5hiXz0jch6aok/Kiit8mpgPvXHK5RapE9Is5+1affUZaftQFsYa1GsgIFE
3S57Gt1vMIzQ5gk7wcwwnr7sejyDNV5ZldOBQKmc/zqXPmDUbbC8U+b8Gn8gpML7
sw1PIRZoWLDAwk5+f5Tq+Q+nTLf4Oh4tn+A4e44UOlEFgCuZaXiUhe0vngpuybKf
kd1JXswJQbhLoEG7D/OkLFndHPy7sTtUCL3KYonc1cPSjMo7tJeKxV3mvu54gMkb
E3yW/IskqzYerAsuD7cQthERhTAx3oERqcgYhSc8RzxJ7t0kORkCYhL/SU5y4qH1
gJ+cAvjnj20h7497pacUegKowqHwsiCKxY4OLVo943gs7Odalz1wUFDlLKDZamx9
95NEU4UMlgHIB79IZ4nArZ2YLp/Oe5a1HuqKCKJ68soEN+wVB6JE6cMG0MVOa28f
HUMEX6OeCZutFpmndzzpmI6xs+kVMrKqQc1Wuo0wfvN9N8e3ltnLT8YPny4tuqAc
StRN7e86yicjatf+Tmnyw+ZIMZk1v3bPZQ7PpM36IQEOg4I7ATZLi4Wfw6HexqVQ
dhnia8yfEop7csZ2MQuB7KkUxfWzV88/1f59HWuoL/Hcv9RNF8RzcduGbAIUHZlC
PbEOF5jTmRnwj8qNYEmdh32cUTPz/LX1/GvUP2EGYYC3t/uA3Ff1jhj4LidZ64/W
v3H4kj+NDej69J89rfC1am9Flm7gRMKj7htjwsy7k5Smo9QoaqgLdnQ991TN7A5o
S0WJBWaXl5Up9NahobqgC0eaiaK4rzWJIFl5oVshILUnMxAZmQwLp8kPGx7O3IMQ
9KFniRNG8fNZV197LZ18eFDuF2WQWHmApMZhXHJZbahoE5rxuDhgwRkGUv2uDv0G
40zGH49g3l1LjxyrXmeNiocHtIsrlaG7Oqm2Q4Mn+Aq8U1rRpH8GZvLilf3/ne5a
o03K4VkRZlQx7MsC7iXpdQoQuNKjdEumgqx55NIhUsGdc4sF+bOXOxsBu9iznT5X
OkHhLVt26f5HngYSyybNpY66CV3kdZKYKMSnuaR+9j+wabfhX03Ju1p2opMYGhXp
HO3jx2Wd6fTrN3uo6duzs4lpCIeBRVa9qoF9T4v5DK1E17pHX26ynyeusDT2W5jo
ABNQCNZeHxmG9pc5Mnp9NyTkaHZX8tTbGzfk9PcJdq1Feakiu68KFtgct1ODa1sW
dK/GJLdpXPxBUaE5/VGBFVrHPVxVvYGJ5tn743b1Fk14cqrqkeGuwKZCZFPWRWDn
y67kk4+22LkiNZZbWoTFUFqVFhu0oC3J5OTUIsogHCTzio9L1bf9TRDdM3VUEaXN
y1k12sxWcardd2cH8/L+VQGE/WpghpB9tPT1bvVPN+LxeqQ4yA4UAiy/n6mYHvuH
GAX4DiIocU9Uzalb5OpgHGflytX009ov+dmQCN9B5i8dtL26oyseoeaJlepPYmaY
pUq1AznA3vVMECvV+coBNklMTeHs6GGdTkY7SRZFhe38igC0M/iYENbg+HgN+u5x
nZs/FnzmRARaVrzaDinuwPdyizOXlIwi/ubOCCDRQmJ3f0Uv2nwIbA5BEF9cHLxH
7r9Y4XQvWLvd33fJLz0JCWSKaSSPvsILF/0yjhAu/wKsZg0Xyuiq6nQ0fNrPTlFo
nWfXMa4r15EHFyGZRymZsby7IHObZuo5iKcIUDb40yJD2KdECfPU5oO3VyGlao5B
/ZP+1V10O6H9fDchsB8TQ1WWzzyS725bv7Y7aGJ5KyfoRz0At9uuxZwGWVeGYL7w
4vs57S3/6oiyvjWuBleQwl+oWy8Zn3ETXZkdV+19qYYBYkvA1Ik5vub9vBnZeXjD
5w50SdmH8i57iGWObgSc8XEgOpEPciqZ8k//XVjBRUmnx0274scha9bkhk5c5p2V
oSdIrwDhxCJ+bq9N053HAXhu49FtmXXovfgzga8Nyh0r5Q1jbWb07kv4EQVtJfUN
zE941M1KKIz7B3F/3VgLTEVSOsxJpbHQ2Zloz4lqB2Tg8wzJsqCcUkbK8bSZTK8w
J7I08geoQD17Ntw6+boWD18Tyr6zNJQSF3pdzsilADX37vWOC5FFmIFmrqRq7pfb
nmjuaFXe0fg3rAmSooSXXqjsjnSwsnVfFYhQgzfKHlgw21rFU9y5wEG95yeRzf4z
QQxEl9UYyznh5pWqsLgZrEXlNWy9zxz9pq6mTfxDa9gDQBfTvhFlPgBrOqnoFNx1
NbOdZsyMTgsb7zOb36FD4Z6c/jQRvPIyhIVVWut6m1GDB0qHagtOFCpwrxPXd+tn
nR+Vcz3XMuKfANymvlPiIkM/Z7as7VzbdF9o20GSj1ZeOC2edo7aIJWCAHu13R03
rQ+AHSx7mlW8S2ViI6SxAaU3eKG0xnkBGLlphGn8ix7MiWlFciB1KX4eUAj2zIJ/
AaSFTvTsm/bl95KULtBz97z86MtYHw7CHmRNXpDJDCor71gP2TTtqjvK8mD1GI7k
Sfx49t/lQhMpmx+ckLqO8ucXcyl3USqELv7Y6zA+MSTeVjE0jsEoI0QmLKhB6O0z
SjvhKcSOV1hZWMbEyAvgDApWg94z0jZXNUgxrTRZ9qzz4z4SnCxQYbbQjIyl+bEu
O48kK+BMGKhCWLK01yUbyUOta1EhATK05O3zyIKkZsGei8IACHNQBINOcVBD5jVO
2qdliygAhKsttn9cGGawlMFwy+x5Pa1C8WgVuoNunKXBBvHTYNnmQYoGDvsS2pA0
JrMBd98VNy/vUbU8Z+81zHaGjUXai6KBn31NjzKvd0U7Xsw5jw9VhLdUd2II1eKt
cSnMmbBoI3KtWEcMDH2cU3hgaZXeolxEE+OV4+xMKS/Z7++vLhupeQb8Gxi0Z/Z2
jFLQeTTX0EILY9Nu40r2MdUJsz+aaI7nevXSMa5E9sMX2z0Whuy86qkOdWU1SySl
wh/VPupWo1iP4+xhcgIqKcT9dA/ae8viF+4MaRE0jcrUpjLL1TYSGQ/viIMqyKSu
aHzRDEGQL+yGNHvygYfL2xudet1k5o9TZG0b3Ffk0N5yiHWqH7JXxvG5bAssKpOT
/huVCJUdwdZeHA5znQ8ClWt0zrxWniwxWNmk7pvFVSDcnq6ySHT+GwqDXKRs1eWh
ZYwq/Gg+JMWg1o23X3JRtSqEbxWDUJLusgFhhLALsQHCLvFYmrfM/Q2h+YeJh8ug
Nw0xUZEesIY6q81wf1a/J0SGbniOZ7oECram7JLpO3yliMRBUC0OE+8VX56EO6XR
jrGgqj7av5anJ+t/xSHzyGoW9mH6JkOjczhbzWGJr5IZ6A1X577Mt+vychi8Xmil
RS0x5Q3z+REI7CJIuZZvAkoku6k2aYVlF2Oap/iUPW3Nq/rWyDmEL3Zi7OL1qWPB
9lmv8TYwj1DMy1aQIqUfC35uaDwzaK4WfiIFxGjLO/9Ztn8D+kY/Jz0i8bxmZEru
il5A8u43s4frVouRQPcij//2uanOvfbfydQ/h5z61qEZr4TpinPUeHi+UNFM/hn9
t++tgREb85Pk22YRJHa1nXsRRq2qX1yAi024xNnoiuzMkV2dkw43yXsK3hx1Cru1
wT9gy67JBAyyEk6+UuNpIAXHGWrPqWSB/CBp8gsjn4sErsK9gLpuB7qLf5NeqV2Q
pkwj+j5cIJLEkzhCRDOqv5QFIPWcuw6NM65Mzc7i2nuPSz2c3/JrfluYKx2PPJdV
3kup6qqRzS8oasLvYu+YYykSwDmpBXpkMfJrf0pRfnFQyCAlDF+MyIXudPKxNvSP
cEwDFrYKb7Jb2C8SZ+wCd2xrA6oCWfUirx9giotXcR2kEBttJm5kxSHdmdhvoPTo
FovzvX9Zq/W0QJTcmL3AyAW5HhDISCTLA9qeZcqmvPV52HL1vs7IHa9ZeamyXxE8
xan0H13LivLQDK7kK7yd49V/zONLjHgPXjb2KWfmLaqyL9A2PaNu3Wp3p2M5/yog
P/VHuxEerrsb5xw+wftsRsw+ZPdap0ZX2vCEvuHu+3k+hv20IPW5PTcQZoEiAZD2
M0xHGx4WjBZ4m//u6o7uY58kWB8hane+moU72W77/KUxZSbaUq56x0ex2xVHNSwl
WzC1Ui+P8JjPS88thJb6EOBUAUCN3O7AX4b3dUR2N9/gfHIJ3fNgINzaSBYeGRxm
Re8TYr/jOCkH8DA9/xwa2VRlSyY7Gz8cY4gWXurS03/q2bIC7tvWE+sQX0uc+riH
GDjuGQUDzU+D+fDQdnjwxYcYd9o42VjoiVgyhqU8H64jFRtNHzFCQZ4bCuAQr48O
+1HdZQ64oIA6/lKsowNiJ1RSkvMcsSqKvEur4dHg5gEkONGfYwGCqtkEG7zkAjNl
YxIxfYplMrSgLep4PyWuN0Ghf6wZt7V9ABjCx5IdX2sSedvS4B7JjMClUCfyXD5i
Cn4ikXPm3QI3Vff0sQ2GrWOn9197DylKHJu0YgCIN/zjZrccaRre+9ojDLHHR4h9
YRiobOHZL+LBb6RXId7ZoGxoiEiobHRWrL06eMrs2ZyBZzYEKTzh/Mt9W247PTac
31KnS9Y6QWOj8Rs74MZLuIpD6P2dfPsSD/AnF5XBWL61fQOP7NrMuOmFmSqH6TXR
HXTlehDSXOi8ujqSGxTQPyouqDyA4LIA4WLQc65NEbTp5wKoOb8ndLWZRguy/n9M
kFeRhbv3Ok42rYNaRrW/pPeeUA7supc/yeos7NKZYDRsn4NfIRZiRYofyh+1a9By
RUzYfa8j42BHJB3IgvjaRJc54FKN0Qimrga6nNluEo246WTsw4n6m3DrfJmqqudA
/WgorGI0z56nmHxgjgZHfSA9OVfW77BUgfvtuHGF+yp3trWVlu3xoX4I9MYs4SRV
8jV63xbDnPSQ4+17FOyQ3cKyZ4g9Ln4WWUfXYsx9TkE1liZj9eIVi7RjRsrERWt6
lALQr6z1ednvzm8FC2SKVqdPuHH8PfulfwerRXkyJyRz0nrPKcBRsIFXjwti975G
2KOEZ8AHg/59LScxoBAMNxsJ2Lm/RoDv1nVYN2z7ujDEiQnfM0Ycau91jFXqZsp7
CPW98WuxyLuBIl5CeCq6uZbTpEfvP596VCb0dwyzG3hAWKwU2WN50w0LG5ppDoWH
yopKJyE5/lpbVI/XjSwKLhWwcan0PUGn2hLwesHg4fEFX1aZ4Tex47a2jPcLp7CQ
85YWyN+BAOiBPkpSAjdKCky1WvBxIcdJC9UEB3u4iutaGbWW2fMNtAwrfR2fR12h
Xn5BwCF1dy58GbNopzTuRZ+s72Qp9oGqYxyW1yYcjk+irn6RGh4A9itpyAGcqXKG
kdqKVq7v54Zmb7CtyrKCklR00to1ict+Cv+H/8cglq4pFPpMn51b8W0ouWJzITpv
nWhojeO/kPTNlZOWHwuMV0Fk0PuC3ZUctXIU5VlswTQR/QXn3z+hVj+PnVb2W2qg
3Ymf5hvly6cu6oTKVYW68FW79PyZrM3b+Ve/BsGuMcHnnzIvpIxq9IahyB592jxq
1z6JH4jzWPThU516JxSRclfKmH3PjPTMEg7F3XR6YynmA1tSCUdLj+g42QVAU6fR
YobaDdMpryCH9DeWC8P83zdejz6cR6cqpQKZT30uj7udYiHtFseCTGmP1gIDLVFL
SvRCUH8h1Q5tZ3oxBg+Ljm4rXF8CaZj9D5tQ9OZOY0SP9+dvGMWKhB7hX1tV+A0c
378OwqP8lrrXtG5NZ1gySCnznnOqnIQaRDXUzDfCidi8VSnMU+uo0NKkUUmtD41J
gLKOde5imUM63KathXPEX4KbrNWFd4lrys1MoKGop2PwTza2xnlOJzGMMIK+rqfh
mA33MRhvXfaEOfzanm9qP1AGDlVmLhQGYRxTsUkNkUgv9TGvKsFT0Ag9L8Ws7WWI
Kn2PSpxJ2/niXOodQggi3t0BPuRtKXX7BapMZzC51q3B7HZN90CfcEIDOQDJzG4l
ta91QlSK0CX07Zs5HoK6dayJ40OqaBvDAUuVIfFUD6DhmA1Uh2Mo4iQiUKpX4Efm
apdthXqbKC26bjfYmaA4OZZAwPGCbzYXNiWdnTMB3J1jxtRo0S+u85J7Ekyx3ZXm
BMfky/ZN9Kisnpgd5wCnUY4+JF1xrB75WWI2meVZIw5JXsMPGxM0MlOEmoFlzRGe
DFrjfUziOhlnRc7jAxhsYuQhdPykDZ5ZXDXWfXMFOHkKPedMqyJW/gkQ+fzjJD6x
aXLKtIgC5TV/aavPUHt/IZL/ucEyjThMSpc4DGW9Gb2fhZB2zL0XKh6E0klmuVKe
hlUaqoz7uLUT5/y6weinI/ChTD8SoZkMe6fmfZU8Lzar5GGSzwNc1tnDtr3OQx1g
TvtfaL1AK4wO4lB4g5ONqoRQ3C5C7HajpCnocv/ArsCRPAxqwt6gKOe47OzOy1UO
jTauttRJIHfDU1FBMVqEf0SKqwEqEiGaPEe5CoHE+Et/0BgG0CLAZHAEUNIpx39p
yAhST8CamXeBV97pWCRN3DEna1/jyKixk4hXfiJIQ/T18SCAuCkb8noT+xPr1xyM
Il64RMjxx7qoKphsngBKIaQDMegoZ94Ix/EJ33Z+tefoGqYN1+FBxYAq0mPgmbnd
P/NVG5l7YU01F1LPRtXzyvUO+5Ib1Jr6Hmq3pha1jWF5Rqmwo2sj7/cWr7FSGlBJ
WEpIHggk9XCDhbmhYcFbiyNJptg3AGug3JvJmD5cez4n/cSx9z1XQVx211DYfCH9
uItuxm9SX88qaZw3GVjs93T/qQob250SfaiNmpaJxlRwbhLZ1HLXSTdtOwTjXQ5Z
im0eG4Hfm5hv4P6IZaCiVppCXCn2wtbMz1Y025nY0tsLBRyZZMxHD6C+XBS9xthH
JkdthmXqKiXDupe7W3WuVChlMCPAxNMY2lh9XUoNNjSvtcm5+DpRlfEmYdK3OvWk
RlA1C2HZDi52IPcoMqgAi6amHB2ReLwopO2tW4cA02i+zx5UEFPO57uBou84mbCm
KbN6KjHmXzhHyJKTsxy5KS1qTz+/BbG5zVoimT4pX3qodTMy27QfQCHNAzuVJuh4
/b69ZqOEE4tUlag9jPWDb88Lr3xXUUEzuXRh90zCmyQ0/N5EuynoSf5ingbbDMtQ
r4+/3i7XcvxcX90JD2MRiKSLPyW3FyUrZigpPt30VXbLmjyMfGp+C3keqv8uNJge
k3yW6GjzyYFtB0QVcYKZM9Xi8qCY8xxtlRnMZpon03lqKktHlo2e2LOuEF/WGe0V
uaPGmQAmTh8XUf+XE8ymu3KzYRsdfFB26I6cCtSi157mPxbu0kzIilqaIPSA13Ox
5NqTFxU1hiqDF7OSLhYT4mw/sYXdAmM37Lr8uwVJ4F4nVk/QJw2QAdVAPq5epr8K
n3kR7jfuGKzmNLJXprwjt25kn9otH7GNQFA4Wv3+tVw2DI5IkV9vXLHAoLREMhg5
dyZStRQK4bjE1Ie7mOwa49o6iha4g1fGkuYNkWibiT+Gk9y3kUYTc5G/nq4M3MD7
7+2/In9oxXcknm974ryZA/zMPwel+DnnU9YpSt1JeV2lPKdSXcdgEJVhMkXy3qub
9ON/lw4LM9x6dw1lT2pwQ6GnLT4t9IhP+iJorr4HDpbS7ObTRUrm6xrIicDxlW/y
EI1QE/e2BQaaxprD6sqE5cGYhoBNRkP/ox8qw9tyXm5ephihlm598dV4XzpuAzAT
4PPR8zzDN5rGnyWjK9Z7eVJ9X6mayaLo35Ajb0BFoE0rt5O4GCR38+JwlEy0pTGO
Zf2FXdcsphAVcROXBcdtXri1NAj6pYHLRjlbezbG4yXGFOIC4+NXeodOQltLGY1i
lOYHFhC2NRq8sq/S7Ru92eT+4bCJz9PsvXfrR6lW5I6hUfDRx1j0+NobyohoF6/y
9lzyDhLYzjnOiz467Vs1kO9nKLBtWEl281L92ydGED1FFxl4kZar9or8vPPYYk6d
/izgBa1ATEm4Wq591Zlo9bq7akd8ZWIgXsd9ZpD/W7kYGztaUMYdpCRK6xAVhiEw
syPCuN46NxiK+jphocc2o4I0Aba2YkUBC1WV2TmG0MfeSCNM4KusMwHOT63vUOUk
TGz8DfLHpdhi0bOcrKmsXP66a9tx0j4FZbf+By/20SHu7PW/rb+EdoYT4ypEPBwr
ASZ2Q6m2P7Jl1I+3LBwHBgxGqaoLth7Fr5ZK3oesg9CiOjtub/4tardp5HfPsR9w
9GzDcRUSmA88UxXXT4dIad8s060wMstpOtTff0qL0KuxTUC/Fxb0DN6S+GzQf9hC
T1XDxroiXZdyz3wEnLvVSBa3YXv4bmrlIwlaLCX1HCXOmquN9EoLOsY4QQS4Nq9X
yvpCYyHt6D002XHVjr298hsd1OIu/W1naMkWarpuhPQBq8s9+z5/LA/A2Wi3NV4y
Cegh/OhyV/QbgFGHVBNEQhatssJrS/WPVFV1qziQg/SnMp+Ic2/oQseM0hTcSzwT
fFCUYwASfEEb2DGZdEkxBU649kmSWwzFV2kFluQBFFBiP/jtid60gFZXUoCON7P+
tlJTHJT67yRXwYw1OTGZse8DxDl/Q+VqGUyyJveQq8vZ/qNvh8YqFAaHTy6uxpBc
qGIsdc2OxuEoeBsvoFmG+p227kkZZli9YNkxxGWyhk6DSwtXxwG5+Tzfa8OG3sRq
fyg5/Eyn99do8ttFD3DKOr4xaWVeGHDdjTbg4siNj19MdNS+1B37smNl+kFjnBnx
+WyDDhGp810k53obN+RBfU1CL3WowrIpid124ouT3W9eXpY+BDxqdelIN5vAc8u7
u+aq7EautoHnPLyeSsVCwN3MQm3Tf5p9MMex2C6v4I4EumVb/AJiF618Ez385orj
Xb4xQPlLESPLE5rt9r/TSDAnCaRawQxai+1yHQh4KCEyAQMjbr6oA1tuUfj5K2xP
l8BG9Y2+Ew13gHLRA84fx5k1h6liSLJ5Cop4FS+hjc+JtiR+Y0qDZc+qR+rF8MS4
uWZqBuGYSCbY+eg59nLSn17/QC/0dpOQFDtlbOt9bHp2SamUV+ja7BVnoQFbT/4q
d+BelNfZWN7rYvBLU1YW1eYt3v2VSwNzsRWQm8yhcY9OM+ClSLK+3xWyrN3341MK
reMtkf5yRKk3y7YBuV+GjrmEFKQZFTAz33ou8EYX0QpoEl59cOcAUsqLNdSI2clT
XVTqdTztF1WPpjHeusUPi9OZ7Re8Hjg5CiTg4W2roKzHIBvsaDxpHEErUaEQdsWV
8Cbs4UdXSsbeUp++aMebMvFi8PvSmskh4jG/GaonD+6Rfxi+3+N73ou2ll9xuIyR
62uEL5VtJaucdlkUbRbtS6HCeB8XeO9BdI6k7ZFdyDHuYLQnH/Q3AM+nP5hS7AZW
S6DG0233KGftRKcRqaQUvf0njmu5O7PkioMI3JMx42uhsdM/m1+1Guc6iAWSmyDz
worNFGMbsbkssFsr6HHhwhNXJfeKsrxv+7FPsr3vz+NnsDoR0lOXXxwdYB09oWH5
rhPg5AIbIG5dOKxa6fq7tV8qQD1koOTkDO408Ytjy14ROH6yYWSaKsZxU+twmRjr
o/8xLVElNUBXfx+i1n2u9MRljznqDmlOfostEa/hlop/XzZipNlVfHEnfeISYgIY
KVcuh7fEKchqpQ7J0e0n+gXIsOCn4obDwSKN+uU//N/v1aeECihS3KcQFiVy1FSk
em0Jy7hzeVxMm0QWXu5HriMGBElGAfG64GdwaX4hL+bvlv20hyhcufH3LrUYnRnP
JKizYvQQ0DrcMMaZvzXKxZ7BPVh6F0nilfPTFftPvI7P16XAJyTPMt7mY8sJNgTO
FSH4TbBfgtQJhWPJWZr3+QcDu30nNG/cqdzzs5ngPX0bpaXF9zpPfUkV/UW/FlbZ
deS6PbyN0kMHnj1LRfttAuh+tRufiJVQFRPH7Q21lmQkn+aeKyxAcBHpvhj0wyv4
mvctXUHqz7S/I05uASrGfcPmiRME35/hdAD/GH1WfKMl78MwTER/xQSjIJbHJnq3
6So2aW3KYf1wRS97aoAVIiJm/leEqbY286j08cqAzmqOkMgf3SRonXoIXIp/aVmI
fRebbe3EncaRQqop1cQ/pWlyzm2XynMugB98XLU4mSAqvsMXfqNJZL/u9KDkMYHc
7+7GkZjcqSSBoyYgHiQ6FfCvPMTj+/XHtAsiEerXsutT8nUbI3qvV/VnMu7UHjKf
h1RBDpdIcjEza8HRVCQHpscR2nYGh4Vn97Bgi4NtzaU+9eChKispdU6G2K/7QB/E
1P/pj8zUV/yXVLVTH4RLXGrOgGMXE6OIz1ZklLfGEhVxHv2g+oE3MSwHHKwRiAck
2I2KR1hu0utzwbxz3j4MFwWEEKlk7ouwoYetyvp7WDYgtXy5++BZp/X+Zwf8vpQ1
P+LiEv4soikyN2Etg55g2kp1JT4y9um1dFqmL9imEBCWvU6KLe4CFCSRhz3n6ZJY
vRnv29Y2Js+AdcFsYkoA0LiP5kL8UyeBRARWjQ2EzEtMZSiOfW5LiEsHziiPX34H
Iox7KsIoGhA25sefml0oFmXn3ZzdOM8q6Qez88sddtxO3NJcxcgv5iOSNUX4Dge7
PaWujta95SZLNBkNbm/2nqUxLNXOHbgHc2skM5UN8A3QVMHJUDc1wo2v7CU2aLst
P27jW91F+vNCf4rTCJzG/cmRIe2pi16fWGoW4NwAVCAmw0WK6HFG1ZDVEt6d+ogk
YP7ttJBIKTUnRtIqr0TV7Mt6IKjSxMIoS3mQFpL2VpgbFCgJ6yQQZ7UdKNmGZtj6
8hSDHyeQkJ4QHXZMzOt3Yb1k4ZT86FKqGHVj87oV1PEr3vA7b5im/isU8/d79Goy
XCbOzKF5xtXQSfTTFlpKY/JhLAWDlSq2AwjuARd+D0dy+QzRoh8BkdwIqPca04gc
SdNklXYeIquZuJowImHmNKXUtaTHv+85K6c9wvMirnfQDX4A4jnJjXB6vPAvpryJ
XJjHvwzdn0g0aPvuxbL5zkNNmG54cbwkxokcxhqDeZ4Qyt/y9aFJ78yosl9c8fet
f55yBFsl8NXn8UI2Gie/IytahGga10u5t/BcDZD6I12IVPMjVLxuz8hVC0nRUypt
DBgIljryp4khJ9xDma1r88PZEKydNa21qJstr/4Zc8vIc0LEzJFdDveOJ/4OXiJF
TyS2+CzZAn9Maa+3L6Zl2vwEKGnsvs66/xKVD+Y2ZvUhZBrPesTQBx2qJIgBcqYR
Q6GexowWB8yVE4pztYEihIdrhhASiTRYJdNhWOnO7gcFQAOJB7GIfemza3FHKIrm
4C36LxpYo6crqY5Qy3zopC0ThFZso96N5F5fzsaudBoh2AC98gDoNwPKf7dJGcPy
ezGe+OykroryYGLlnRCUfeD9KG4xCDX95OEGHDTXWFlk0rkMxjVSROk8t2zlCpz8
dUPvI1hpE4GRDrvkdpzLqxUA8mMKUGx2Kc4ID+ZrV8Rd1kWXugKt0jn6Xd9UYu9V
mjOx9C8EOPywWULd3r9odIwvWs/6hiOCObcRqbGngqEhc9NpWcL6lqlcVIzJjWu/
/EM8WhIap8rnwQ/t4cuoXQ4tWsJzHHEbrIUmbnU6uS5TOcAHf+snEtSKOrBk0JHB
vnHm8B0iq0DxoEX7Gz1IdIxHbOLGMLZY03Y2zVh85alKWOy1Kqktj2pmfio3aJkS
TCMOoZwmVCEe+HX5nBZe9dsDIqrKAs4/quKrtvNgNpES7V7eeclnel43MPjhqOD/
fhRPL6sXEScy59AclnrNO7JNqBGI88c9oR6PA5MQZFWEETU5WXsUsprn0UbiuNdV
QwVIwN2BWi8vSgt/2qbNVawdu93/P4EN04Wx4xMZLA4MKyniToMh4gP83veOB0ue
bOFCo2NSoErv2WACHwT6L8I76QA727BQPBXsUKD7MGwN8Z+PIu972f35uV/rBjJp
qhCbP5Z6WvVzCu3v0KQv8JzfmnpyhVXLEjlZUEcbMtNqLV0b6VqaXO5v9mJb4iZt
sYoMp49vcgXfdP9mATDb/Zdcrr36yu2TUDCa1nHlaEd1VSw52oSomIjhEqyIkRcj
FBs6cSxeJaYi7oVTFdD5OnJ96c0N2ogJdN447oKkrGVfgAs0kp4Wjkz+K74oOWWb
/p6hA5WeMFc9GSM7trdE/2ILbqUEsrIUmYTkzT1Q5CEHu1uX/koKwzDnDfBm5AGx
egHLMzGhHgvSNJPcq7lEn4/ZuJGsVQfDQt+JvSlW00ylmaZ1YGqdHNQwUsTLuv6n
OGllhUoG6z3+k4+qNCUOizLhxpvEk2wivMhi/jYnFbdy6KoGnGfcg3wV05c8KeQ2
wak4ToC54h45ZPOsUAmBZs2ZCbGydAeQCoQ8w3+tReuWiq+Y43samh38rOErUM8/
dkbor85948RJO+D4C2GwaVwi3TIq9JKWNHDoPXjUwCOQ73nbC8xvYwiCFd4tGpeG
KMjufItbyIcjXHe7LJseZMk61s6Bb7QvWN24Vj4ITICCwnyKWjodiNEV72+OpT1o
X0H9G4uaxNGE2afeB62UTEiygzPMrw27nYZICcBLP0XrLqOzX2w3xWt9bifsQOcP
hiB1DGCKVzKRUTXXKdZFVEIZnFdaw46x8PG3aNRVotvGEa4SVLoDcAVulyd+aGaN
nB0EpVB0Dzb4MY2pwodFCHa9t2iG4I39cjQ3UDMziW25HJvEO+KL7Jox51qaYEa+
+Dcr7rZrk5Tuj1016gWWi6m5vp33e0zDM+TIzPWhxthFjpce7lfn+tdNA4S2kdiu
UIO5EikjvyQRlfhJ3H+afS26Z2pzOCKYobWbFcVjRgUvsxr8BqnFG88gATQ7xUCb
IIqP+nkcUnBtZ+k5uGSDU2mqCP2Uk8tusZ5C5aVD+cfnB3UzxY5ocabTMk3sTqYZ
l0gd69maHKCf15ZCiDiyyXa53ExMkLxyC5oWrnzqhD3vKZSnll/SYSXEX4g9/RHZ
maqG+7uSq8vaC5xNJ9VS5nc0rE8ul1Cm162fz2OI5Q5vonyT/0ot+yJOOmDcIeFv
r2s1FuZ0seMO/vzU5tWZoy3c2kL8iJWwBjVLcao+1nYqZGR5Q+5tGOoBFsZ+5iyR
bshsppPRi2YZRgeRrQbTCIMYC5zGJvnlX4JMxFp+0sQF6UnzPmqfpcZitubB/N0N
7ugjw0o04SB0qg9rN1kfA70jMY6QzBNZISykvEJ7cspSutK9cmDV3LTTr1laJThF
dyoWo82l4Alh9hkiCS9hQ6giJEN0GPoR9qaA4gbgVR8XA4WeES9GjFYKiNJZt4ut
CO6KMs1qvMcCiXf00t50g9UCOwJfOx165UCUDlrX0ZS+PT+giUQhexmXgXB6E9My
bJNRdWZuoV7N1+ZxvS2DGumiVSL+lf6Hm9p17diLxUcAxb9McV10WMFRpyezg8tL
GNRFuf+WRXDNIH2eCuNsirSqHQj0iWDr3GnLDqpefzPx78ZP2QYeMu/LJgC3ytyH
1vkyMNeq23GWaP4KsO1BfL2+G2ci3DdyeBMSd/VxOdTAMF1vIKOJpFrMvdUy2fvK
EEBej0nZqcNLgig5WefKQgkQTrFyKvKiXMnadSgBI4gBqLeLXGB8/UuY/ReXiVgk
V0hl5y63zj7G7FG8MgK6s02wsAJDF6I/bnxIcFsmnNJLN9NfdEvONgSt2zupwXTh
Dd6otc5pzKfyFeWFomoSQkHMw14ImzGeudIJkPNvayd1gpkmtlk922q820bwMLY5
fQca/MvHaqmKpG0W3jvyiIcGNC+DNktUjBSud4mJm9a7QDFjFNjXpz1Zps0e+fsP
HFpxHOpCRR4NlCWo4Rl84hWkc+1138VIJwBihHVgcQ9pWY3xPWB/QkKi3b+Lpqb2
wHq1mCep9qDqcJ4Hc4SU46CaBKBJ8Y8Y8uV3Jrx2t0eChRLgsvlvt+ZjqztHhvV7
6S/k0txJamc7nuV3z0IRqNCKnRQgNHxt/NxEGJET0p+FAN4XyC+7vbc2TjHTG9Gi
fCJWHWjgGmhoexpTvIq+LwyzhgoJH82h38s/Id6juwvaIHTKKY9obwJIhgSKH97j
Tz5PfnbN/hULOLOwvoK+eK1HCN+cCsmt/Kzm6ndunmixR/j1sDmFCzPCBf/O0qE1
1bWZCe1RcpQK++MswuwKWXbKuySNMkPqA7PBptBukcFj2R84oiqY9e+jdKtsz7S6
DJru97KB1WKZTMwS75LXM1Ck98G0PdmDjSkcscmE98k7GxxPlrDhFsijU8MQfsUl
deUl0A2dSr+4Vg4w9ZbHg8UvGcdco80nVfbVijpsqYsAyZ3xYvHYZL125v21zrZP
DxIvsBR7oZGlNJjLSD7f5e7yteLqmd/XGtsloVRRGKMCJT9mHs304RgBMIifvBRE
CAy/uumvXEXBeZYPXnIFcsOl7FNS+BSmYUPasrRwRvJgjJrVYkn7OEUpbaja9vum
gvil2LZkHEM1iLAu3lz2iTkFUqddROV6xDEbgT/Tr+JRUxOX7bG+DFJPXO9hqKkA
gedpiCXIv3m8enkXOJwpkcV48TSB2yc6PsZx3kXaBJZUt6RuoZMOy1rCO5wRTn8R
AkwUUzASWizCNlIsbC8EO2HN3VjZXMR1YO9lOGyi9wYYMTQWvnk5XIM0cXK74eFd
wTuKvxqwjGGmRTmg/btJjQowZVdN1IvKMJ3eEIB8SE7oUqT/5CYdtuyV9nwUVcjE
o2lC/iNos8DHkybfNPEZFgf9VqbRwcLoQUS1Zuc6Dd3++MIMGjcr2pYHnAD04PUv
9L1w7P+nHmpBCYF5/Qg+SQBXXhvSSqgjVTX5jtz5qDicVP1zZH3IQWd2BjsbZgHB
6EA7QnwGgNy6U7SzINCNUt9SYAjCU+YYUijrxN5ALrEFoJOSBpGg2pPzTulCowQA
CUHtMvkvGFGwZvppbVwv8/Orix1eoNymDgRmYPK+97smvrS52uxJ8x3GSh4ZNLHK
HbC0eIRpxb9Kn5CC4H8dK5j4xYcyUuIr+UZP4VTiI9BhxB9I7G0AkDY0qKZvbD/7
GAjHlfKG0r3xaUTK3gfNAYySI8zAoAotSaiR5+V225fjAv5pre2ThYcxa3Pn03/J
7p1gc4semF87ha2zBt3NEIJJRiSvVPGS+ShIuTWNW88sX2yzS2c9LJYMaW5sUvt/
6LNUjp4FHdSVgJSPT0F3R91z4I1NImegsvzsRdg+++hiRiOKALZYazubL4jLfPbo
lDuXbH0ONSqtgAD0XGMv1upLfjpXlqPG5PmRgSafswy5yhKMhvN8+LV1cWOAQygK
5/1osPPrnWbYO1ho3W5vJEJSAJ6INW5LBfN5P4Dcp/OtVo+SPVPqhb5lyPM5zPfn
R4iJ0RYR0tHFmShJ48RyB/Dx0fjFIOXmk9lT39Wq0Vtv68iF0uLNY9os1XhLlf08
5dUVN4/dAiDB/nNDYk8KHRMiKn/2e7swSCLd8ZH1KVW3D4RPFq0d0ZmDCxuWjkXY
lFPdlCswbT53YP47v0QeWl8c7ThHPLThONVyjZ0Zqkx/RgiOoE0btWHrM6aGW2HY
w2Jmw9uYychP4qpwfqzEmD74iloLas0HlN6t5ho4JGOxVncFNtPWW7VvPPgqJcWH
2tMBsuvxqqNl8WXkxH4PZZpXtly19f1c0NgUamZKZiNwymdusok28ZElwpjw4elO
JsEwxlT+8l4/mfPbrqRTJSb8ZRJ4Ent4Cc3hGTAF+ZD5sfVJCerhIa6S7aJ5hyxI
2oY5Cq8zzMkdl/OAU8TyEv3Q0DLtOxF6VbMO7V5z9Da8Ewq5X6b04Gn4AkmRHc0k
VvwkjdX91WOfe7moHgKAo14r8njR5pDxWkj3/OlF9g+P8aDXJ+okPgOQ4PIjGDeO
+OMoALsmpf6Ev542g5TM/xJI/WUfOrYaR0nJdhM23J6AC5ZtA7wjxNxZSosxTnqb
mmM3w6Tjb3WWjjGh4HzpQYIb0j3y5apTxt/DjKUtpozIkGBxYux4uuquT+Zr0ckw
Da5ohPuYyXI117S8IL+6rGMJZDhmYAIcaV2x/Y7aVeRvBiDzsIyJ+EbDvKXQw810
W20V7OwoUhZ3i3owPEeWe2rbq8CRdC7MgaMYX+xxxtKwEWbqqDvsoMSZvsZkwqRI
kD5m1DB8/ZhZgn4lh3G6dPrKzexTkojWZk7a8et8nbnKQzsdkulrxsdzf6pLpoFb
YSl3Px7Adzv6i0J2i/dqXX8uJ2/HGtEvd1WbZLZrsBztXXE5zGtMyDyLsoe9VHP0
FlBuu5JwYnwsvXm4R8lXTOSIHhkOvDl88xIESeSZqlAYwZ2tYituxJAVa6bcDWLK
nxhGRlvI96bdGfy1OTy6j4sICu89iXEjhegUUKlY3ivZpk2C5o3VJnwxfWGpWbAQ
ChWoQKOAB3Q8d1LRgvp6V05134NxwC3Nf0/o/I4ZyqsWHD5780Ti+7fzqxCn82Pu
YVRmBx0lBTjOG++GwBNqJmw5iNDBYUzPtaaAtVgiTaW5z1MUDilb5Q2AOHLZS/R/
5FTXfpZqQcBPW/E8Zt0hHijlGZHUp0Si5bKTfnL1tiOmHe07RCiIAlfQOJpOCUYZ
WysgCFzUZbti5ir57BHieJh+xVzHL4SZqOHM/I6eEU4E1qW8THv8htMi08wCCUi+
XDn3MUAj/58A/nMJKFD0Wsa+B7M0L5Ha6hz2q2nWXVVa15ijWcY2qPEbEnhr8q6J
dP6VsfuY3y/qaALnHYr9GuyD4ocIvNv0AyIxwcSOogNifQ4DZkJ+QJJfxUTGUyKx
G6BfPFUjpxdMV0QnUaneZtEF8JW5mNUFtjHsZZE0REHtnmniBoI64070zUFQnOcU
kNsHbjaaXADu3LR2IaREpPkw4vqFC84cNTMwIInnVdBAap+bvzdpBl3VVmBmu65j
3EoVMQ00XUlVw3/O+1J4ZgsvyhxluL1pcP3dQi5eibN57vIWNa/BwPb0mdoCFT12
QbU1Dx7cvtHV1tX2ryIXA91PlbDBw+pCZ/ROxUG9vWr0UNvDKSj9xRQ8Zvd+CRa5
Zq4n3h3SY8BzzmrJRy8Y1V0rJXEIL7zH+pqNHHHSdEdgL6xAUBAvT+8lXSvGPmD0
PVZrbI6EBXiWzvX0riExjXt3dceBfq1dL0lSs0AKp/GT0P4q3P0805xWBMKK7yGN
D+hr/5aWFd2l9EdWMQn8lyQmstYJo+OKCn9zs1H/4FY+ePfJa8Lie5p6e/Y8ktda
8CKH4zLwb2cb7iPED2zTsrMVJ1/K690IuF/ZKWHiq6+uOPyLA3eUho64ASpzX/kf
6EcICPkEKccaEpTAlPxJVlkpXtNNxDftY+5/IQeONdqqNQ1GZd39qONsMrEYV2e1
EXNBbxe4U6BFSKS9IhJ0nDrlIEHcu8RxN+QhBv1EHixbQxQb9TKzdHZkSlLdyAnD
PsyVP8HFpUeTKPcS43wgLc27hlycJNsbYcQO98TWuRABn//qITt6hj84fdy9DSE+
Fc/m9ohqQXpeRCT8Mrvthei7UZee4VO/fInW+YoWDEzoy/ZDAQL0cd5d3wuSPxAm
S5abtwoR5CPK4nNXDGJPZMLKVhCTTHcxfnBdCK/ec+TsHnknr7mva6ydDLLJou7h
PjfOjhu0bfzoxgXD7odwh+I43CB9O7UWEfICbM/mQSclp4t5xNOi71YuczdSVCBI
iAzAMK79LN50JfdzMhHHuoljk1TwboFbNxmXf5cfEb5QVxHzsw2uzl7KBHtrUj4F
/rUTLfwBxB0VMjHkSUkSB1Lg00R1BBuPuniFcKPS9ozRXFKje55kdCC2MACMn/F6
ajvKz/AIgiIRJ0QFjNWhpbk3g/VolKIA76I5XRBhShjRfjDKImihqp3gTWd1TLGD
XbGLif3KdjV21OMIaAI0pB/6Krxf/g7paoqwRVGnmo7BgRyq1hoxLJjmBsTcm9Cy
/5GnmuP9HKKYZbnMolXbPO16Ca8cgzg8bcRMnNKOuDYgu0tvIyr6r5MmwuwSvehl
OaQKEt4By4Vp402KOqgy1KgEiTuEr6JtUSbMxGPgMYiYFx+ppGUDcROWBoqYy8GT
I936Cbni+aUG9jeP/bDo8m+bi4SHW2+PyLR94NBi8+Kzo7Zk9NQz3BH1KRKUBQnN
paKIn9/YTuVFZIJj1OyQSr2eVgpR2ydRGlixWVPTc1ZemidwmuLZ5OxFR6lXC89J
N9S24Uw+OL0YrnG3Y+WcWiNafpB3cK3vv9/qVmanSjt1j/misx5gSIWnxLBrrmIZ
HURENpV90GHcsTRhsIG7N2E9c0zCuZU3uCmB086zLkBg+Wp/UAvrL9CLQcVfBEXR
C6CbEHxrdaqFryxjToFRybHjDZCCKeHVeXRzxDpJTuneHIhkX1IrlVFHl5mFnyQj
fbs1AWFNBvUlGGbBphQIvke95wPYcsVt+aQPA4Z9Vy0=
`protect end_protected