`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 27696 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhHD7FxlI0zjeeYUDWrEWJagv//6zojO6gjm5uu/XhsV/
xISvl++tlH87gO9IKcX1rjatebWJct+i2cfkKtW+GTl6La63vjG4dYPG39T0D8Kh
YllykwnWCQVlBkXQDOvWMYUHbzWZgbW/zsNLJchVYVdKNn4M+xAQRB6/bLoxAb9l
PlscSwq91d/Pz1SrJth3LsR/p/tvCFZSeQm4a6r4UxWc6L0Bjt0vW6ZWu5Fg09gl
EYKlzwZpQGeqSfiQL3ICm+7J9TP1UoiSTu92XH6S2K80aGBgwhonjkMCOsFs+MC4
sTsiEJbCeaz4qTLKbYgRedOY6f7lhETVfoMDcw7k1O5pkJJqHvPj/bm0U6VFIuA9
QLzBJM/9KEg7YBlgjkCYrRERdJWNt6Wp3yQbgRv5TFnTKiPU65GFqFGBQ+1Q5+wy
Wd0oOvHoxmBZ8J/l7r0VoD2O5IxQTczyrpWM/wpn9MKmx77wsaVXY2GVeXV8FpOG
+VdWf3z/M9pqb3/J0CEmJzTdDl5/vSgk2xUjX3KRinyBpXHDaqBIODlXk7jc5im4
BQ9X3PPX1cF127fojvCXfVdTNOGAaSWwoWyBbn4+D2cjrZhHqqq7eqIWvp0/TZns
cIk4odnAscQMd5n6PtGW/DhfRIHmtmNbqy5dC6F/y4shYXrK1fWCgJPd2lyUUCYz
tjOTL0kan4xbR0ivcXuysxlljxFdpcdg+sPevyczqD0Dk6W7pGHOGxUJj3l2pw13
zjJifCebAf25MMc2BtCQzkZiZ34Y9knHLG2JFkB90HjjNXGbTJKa3VkkUWCMtnho
RZoYCpyhkT3+tXP33FJJfXOCr/0DWTGUQ+C4fyna2AHv5U54Vo+B73Qwi7MMjjef
IQNOQZFaPZtD8OSgIg/uLxhO51qxq45WsmyG56g6WjbNmamHjRvW4a4tptZ9612G
IuwvIYfTlmLma8Y4xZJrCw8sUI6uxxrB1xREz0u8cN9SgfoKTdIIJjc8kXDlI3gw
edNtTyDraWbtjpsy0U58+YeuyiXOJQXbkvMjRbfJ0vcFstXDFy2RUc1mc35P9GZF
LbpfkzK4X1K+IyinYQMxw6YADFNcle3RagGHKU2Jk38yKKeJdH3l1zQGMv8ofAOY
IZAruQ963WnNMT3cTro4sjqkFBCqG4mu65NmUoYPUnjJTiBOKIsWP/L7Maukw5u2
/HkrtLjuzmB6GzSg3VsuzwTi/l3q+ya+e6PLWfpzxjVi+97BgbwAJ8ukB5ktIOmD
MqnaGv7mJ/aQIJRAMKtcHR6mZYOyL4x5LwgzZ1qE/pAl+BydPH3Ak01hN5JRbaUj
dXi1xZKbaurENgjtmjWR+17YI/lnNiW+JCBSesjQVk/PugwKN6g7PjwcoY++TEaA
P85mmPttexsH038S6mjEq90denf3YfSWYWae6QuDtPO+hpUs9H8SnU+dcaVQSc+4
YLijh/US2cRZ58lZuhTee3OTZhqi1VGtB8dm1xSdNdK5zhtw3dgltMktJHg4OMIC
5f+i0zI6+NIufnWoudMtAOFrOIgMMsWsvD8sswjRH1NOTZPy5CTzhDWMZlx+Awj8
/wMyN26fOLOBitaw7zDTSpA1rXF+NXPNqN+j5n//lJawweHJ48okpt+/78+Wa91j
syRITdXR8J77c3n5fY4X4R2E60LV5HEjxlpw93rte6099tfVsW0V57V0hjRxVHLq
84hgpIntoL5WrYyxraGKx99IftBsJWdOts3vbYXg9wg5EBw58PISJJEi7Vics6Ty
4M0UKmn6PfmFKtXh7WldN2CALgChtgNYUuFyFdqCZIHgFM99OfZcpgZBOjexugjm
g02kxK6/PRzJgrV02VIpbVOlWHUHzQeI4mLUTWXex5s7RdUriBOHylqo1onC2dqE
D2kSyTC19KSyOey0ajNEpk0TIawi6VG8QHncYuKT/4JL2R4L8pu3EaATqugyMfVC
wDJScN3LPeWCaSpLpQILRfkKt7gJubh+efWB4XyfWdLj8yXcnDQTAQgjZlkakC4X
FKE1whnz5Yp/rybJ+jFHHwzEaFDQJog7rqO2cyPgIdM3oA75Rtyv/+9owCQ2JYzZ
9e5ymPfq0iPAVp6SXoztR0W7DhrbH0eKEXbxObtRMZKqpi+L8UfSiKgwqvX+AgR+
RzJFjujii0WlHNVtMnnKJFfs3gQXBjLHhUooSFeMh9miNNYoSq62ihxYb/Ce/5rx
POC4m9ibVS8kSCiS+PPoBHUtsD04Zb8b7P4KAgvEZJZNFnxu52aAJJPQr8kXppx6
XyBERdO3/NStupfxYZ/xnZUWQ0vpGG1TIH1FtV04OEtFGgOkQDULPeGkfyvFeco1
KbwRLiHhxcX8fY9DQ0hmAjbhZgncRCYaZPbT4EjG0+FvHFdiCBOMwIugVw4mSW4j
GwzI2E6092T4y0ekMYUg8nQsKlvu6disWZk/XuTtogM6DEZvNLLmT2Jj6OmhFsrQ
KX4KO+BZ4swnTeteWrTcSwtfv2U00iKpjtt5L2qL4tsRdG+NCLXz7NqNYQL4d+6z
AvpEUgjM0hNyeulmYgHf29M76/BhlzmvFPAmGEaH8raD+9jzaTXMfYiqy3pAU2JG
TWzaz8T6ms2WgRHQmUFnJgdL8Zu4BgSEwne8WNzo7AHja+EyHXde6erke4e1WVSi
QcvI08m+VrDSWNJpXAL2ifp4MLSKIsbp1+YswK+W/d8cB7oDu1Ld4VsEh++gtonX
HmE2RC786wQahJCAt9zlNjSuLJ3qKR3vRrQwhBwSnz0Gv5LbSKDxuIyLfoYleGnp
WKtAh30DJSi4CQFWl+a1h5BFCXPu7xG3v2il6g/A2EuSYMQU2izDL0pvu8cOEd+3
XgrcM3KAx2iGHKDyBfWiw0VLIYpeWfkIpTuGt94A10ggeebdNZIp2Q4+lLypL8ll
CFoxdcdYO0OqI0aix6AXmQuTtd6SgvMwxcTRQq29DMNY5fijlW+lTkvh62M0iRxu
7M4qy/0tekQJ+hxYljZl2hema+qRdbdhsErcGXiuXGZ7paKkI7TMGFfHV+/WNSP8
tdbwmDRuDC6AK6i96+QBQDxITmDr2Dnipi8VYiggm+4DenQo2U1EnPyzUr4lxPou
Oq5dbuDwg38Cd1y2Czy99erDaEaPEm79hWyKxMD/hQPbGZ9PdZ/K3lpgMd+XzENY
1vNzLTK3Pj4N9TuuX+1uz+lo8ehh8MSK6HTe9pD5L5RSEx1DHiSlGV+LXGw5Xny3
skaGc5+5okWbqmtZw4NjqOZ2WIyN6azonHj8nbFvjTw7tx+VkMl0JXmhcMO3fukQ
zaeRIgx2uRCwAcEIb5meBFVdcsEzbo07CKLvgOdJ3Ow6m1z+5vso42eD/iX9uov1
60xO5RvaLcPPgNCtBkyxDk9eiH0eXv+wOB355tqXnW3FOFwIRzCw5xYR05nfET7m
U8lDCTDvinBetpnqMtSevCHyA/LFA9pFnbRZbeCwII1xO3MaWPnDsTKtz4HDNX4Y
FF7RXjvC8475/HXwrmNXoYjaSb5jBiBtFlWEm+O14EqMG5GXxOGXquRYZPQa+KoJ
Q3sgeLPTv6FNAcTygkhi7dbADXftA+BQkfGNMWIxYDmd1tHfD/QLG8IbW2QrIbH4
IPLkfYPKyQTI3zlDWaAMdilYnRtVAZt/VndJH36EZxYxGAppXUKu6TXdML61/9hO
iLUjTzTxcqV3Z33AVLDBXK4yThHJLzV7EN3/uPBYuq+aX6J8LH3H79pvxyaDB4Qq
/u0NZKBVM9g7Q90zxP6LiE0Vl2YcHIyo9iWYDGvMASMAojtV/3ZFGr0/HkkS1XxN
KSRW/IqcD5qoKPZ41A4XVKTpBJmAMY1f5Am8ycqWmMPS44hS3k5Hy8EfeaYnusA6
ucUpaQbfZHRkRwibm0+2bwnB/8GYRCwXltoXlk65HuX1lsEORYGLpq18CE67qmBg
RZ3waovjuGnb0InWngLfDieVCBEvJeKkWmmpMO+lZgL5BdeAw/ic/KLRPfmhu6Sc
5kYIYqvNkSR9GMHHaEtrxZDfCcW6nP3M1LUW2OlDRLh7WgH/bLtjrU3jbe3KcYNg
uQfcaPGFQxKUcFO3MY/4U3odiHzQ2J66oB/6ExCVVQ90/xdjfV5QwaKE3gwBytzY
StISFUr8I14COnvFlI9PgSz8fln46UVhi54SKTyUY4GF+3WW+qMZm+B2NErG4Rog
8T3VtNb+jEWYJaFXlT1KMJht271CY2fp00x0s6Z7eujTDEInQo43cybOObjcR5kf
SOrEvpmCKDN0lpy8OccVF55ltJRZ2fm5I3G9KMcXEyyGc0Pbz+S+jf67nmFrV6ht
lO6fMQHEDXVshNIl7gulNJs1S/rw1wP/onFadOHs3yjfhtwObQ7/F0A04XLmY7RR
INFxl+anRhI8uV0G5vn8zBP+oh8vzjybIv/oT4Z2sSvJffzIBYV/GCVTY6M+r3lr
baSsCf5sl2fjtjb+4zntqYcxdCps4/rg5sQvo9N19jBCMoFCg1D2xBDgulDVX1Hh
VeaHYAuOSG9dcvnQC67EMEzJumSGewUUTwZv/WfGNpv0EmJrVDB5yPmV5tGAUKXX
2LDYCENfxCc5LRr78hIq3GAlk/IBWGKIwNkFMtPT9r+biVRKh3b4jkQBzENzjbGy
n59yTDZo5FboYBm/yDvaLK/k/cv1LD4jrFS/w7kMV8OjX9Z+sxl6sI+sPLtL0dM0
8kaqDGYYt3MC0WKqZ2X/2/ngpO3SUucpZ7MlO1nOqeWdPjdV86/K4cUa1rj37c1p
ECaOSzRLJLoa9og0dEui7pppNisSystm/N+EZsqtNOQMHQk+B+QscfzK//LEkjZK
Eo/VMGe/sEDDJrnBvNgQMs1qkZdzr4SPWE8ySgv3+Cl+VtD8xLXeEiMAxroAoIml
ZT0mf36k3c4htNjo2NfhYRTtQ84VN3y5QX++lZwTLxWlxYZdcOJKIu2/KQBFSGzh
F4F7Vm4vSXMXYGV2cZVxHWwpvN779VB+VA/Dcskw0z3xRHRCUcCkhyqwADoqNp7d
vZWI2jOuOvckgwiaqnbXG5iMoM7GptkVik0N9bQoFj4XacM5OEKdDJ9meMLB2yml
ZcfEKhkyLiz85pjwz5OlWniK7nAxb2JlnqHfF50qK9zlLWmVQBu7H+YZxn6lI5Aj
D7FELkmP7plVCkQCJ9EBlvShzsA4WX8H1CxGjxl+iY1Hutttxd864m8U0JBMUhDJ
gaCa5BqhcMWZv3iwe4vAsUvmFwp/fiOo6Q8lAlvlQGsDee1V1VjLJlhZ/V7YzXCO
VF4o6rw9AIp3N0WRgIEz80Wp97KhNGD9OuWiXf2VuxbcN195UX0NScxKtYMR63iD
E58fzakIMpq0LjGLqghx1IF45KqDGIpM7kOUL05eslhFwcXEgRB1ObxB4UpNgYK7
phSw6TubqyJuemKhPycRccVuBUgc96yvFgn2J6NS1afoV/OhiVGFl+AH1suMOvIt
xnVl9qD9GzPSbs9IOAey1A5jhwLt9QjDx/ZV7AO2pJ8obmCsaoZH5WR23E8birZS
jFAS2oIoHJ9yZm/7Y8rBG/TuCJbCfkR6gz2eljWIXDM04uHTj1ZxRRZo+cJMb87c
8LSA1wOZ43j/FmBoKCnfEkM5Ydcntxr65joB0EVmzEOo0B+2emjGi17UcwzmMcGw
F1pbz0FlSliLx+W1PKIhcab5LTh+uqkdhh1chyxi8j1uMzC/dPvG5VBPMJHIAd/Y
M3E8Y6S/5GPXVRd7RklNv97VHw65I06jpPVIFZ0fW3xV2Dk/U7kELt+S7lDpnav2
2nNpWLSiovwHPKkmWkxelZ/mj+xNCD/0/sxS45p1fkOkR2jDdp+a6vnmlZVLB6sB
77wSy+8vrL9Nox8scTnQRl7djQ3mn2FvCmu/xIoeR0tb1VpINWy4M5a0BLoqvnHZ
ePcy42E7wyKkpHj208V6QjBMI8X3ayC/7TrYxNy9OrpFPWWZ4K+yVWs90avOiK7w
W9z8TH8PJuyFZXzV1fYQAttw2SwhVfGcMV6oGrV16VEthmj93PmHvVgiZ/RASIWX
SiW3ikxY5s9oRR9qFjqmzSwjLCOgAZfWmtPJjtqg7r4qmXo1+aIprkAgGyOEw9jm
tnRZXd5qEZhoiWNXT/jmPAiVqlVJZOtD+aU6tAtaWt1e3/q7M7Pozbi2gY5lTBjx
GlYuOZz1kM/mFA0jWCg8SRDrxdikYtdrqwok6MkevrgnsUITkV0dSu41AeZ9m5oJ
7sgiT/avowLhMWOc26GYQnld20eKFL2GpVAZhrvDJ2fCwkIywMQmNMcKufoXBmJ/
MVsfWyuSeNAyFwE0oQMauueJoP3/2LPwv+GGA/Gu7zKZPHyZHGOSHFeSZyoYXJts
T2761tei8+abXQEaqEqcNsliMHFw/RR/1V0vje2nybZxDC2Mfz3H2mYXl83zCxrT
07ciREtHTCJ2GnmYTGAEqbQoCBIB3PNrXyGEBWXgNW+xLJeRfBTvlWkRhrog57jS
YM5sRVVyZcKs7h3LAlKm5q7sBAQmMpifontwU8L68sI8brFbpnEq58Fb/e97p1EE
588rIfzYO8mzhEFbtNzMiW3JoOJHKtneGpd7NxA52o2xb0siuUPNq79bOSe2p+pD
jJjsdFkxQzcdKvkzSv31AG0ZykvAaKMgBtbTX3SeS3OXbhpdUivrz0+HyoNRq/fu
ZLkqB71LU25S2UwpxtVoe42T2HKVSf+PEJrzicZesXiuenDpv8iPRJdwI3+lClsn
fHGSkv+qLOkNUuvEmiLJ0/B3e/IaD9RtDpenHTSvo+RSCPBt+9194UaMUr57XV++
5GEx2VzCIikISTsdIqk0xD0aw5zcJgfkVeqbjTBbFrWptjktPy7Eb0CZwaWQ/IJS
hzNVsFE8tTG4XQWT+ard7v4AjkFbyIoXVJvc5eY57awtKXxZ5lB6xnnG4hLnnOzQ
uOTLzFvNNlgtofg+xo4a/YbuudFAu4Su1nr+ZjqO58cHyJMlt9hHtaWDMcPZ7bVK
5GgJTDLlGRziBs8zwcXfvB4w5MEq3xCa2lxtfjkcq4MhHeAgv9ZxyyEmRUPJZ57U
hzHvML5w6n8GSToI93RZDv8t1q3aOSIoTyK0F/SVXiqqzR3Zqaxt3Ut3zY4ACbrq
tri1/JQI765R1eTTCAzv4Tv37Nwb9nsBR6BUi1oqAuwxAvZBCo+sETdaHsKI1xkZ
nF+aTb+tvw0uTxGqKbwiGTBR3Lp0GNhyitldUr1EW7BEb4thd4sv4ME9BUbXqnH+
2HEpLT+Hw5ekjbvODDoiiZhYnaTKJNI1ySq3w+wACVEwIbef5eyWMgup4QmFwBZS
dBJ4szWAEY06haf2PoP6wY31XUOz6jZZnBDv0VPR0dzqsb+IArAcr50GAkuIQjHP
CDYGUguVBDNbS+lfYAnPX9SjLvHwsjYRl6P/ci8fZbhUDOThMHsOtdMWRd/KTWAp
RIHkewa4zlcrzDPbqiMbfFi1sahgI6cg9pMfFJG67hnNOlQgIWtTbp0otjbJc9Qo
2WPuEVPujtUi+qhGK53OR8qDeW6Kk2OoDnmiaVE+7HT1AOOPV+rsLWaMmXwN0QM1
puD/cP0HBb6O+mvdoNIoE+r7kn5AP9w3B17nriE3Cm8bKJHwsIWKzIDin9LDF9Bb
NyeE69wcU52G3YzmnoIAgPGhEjMjC2e2BaVvOy4cYBdoDlaGFe2VBUvigyRk60ak
4Dwp/d352N086f8g0ITDT0HAPFNCTT75pfAYWw7h6GBAONhFjQvRfOEE4fOvyDUO
zApk6b5E1velRpMt3BAP4lVXP5aGGMFE9ilcVBtfYdkZHEjV3sYXmn2aZtrsIKaB
iGyFfkNv4urcuY96FCOOTSw0G53tac5DMVY+qfrf6Pgridb6dvBvQ9vIk8fiEiqQ
EgDpgewXmbsX2rVQP5CLzbTLq/jHtC4cwa8uEGrxeWHKDJbXkhejxnso/5Z8TOix
Bh9JcroxpfQxZ4DYrtu672Dvr1Onj57LrRXW+i3ytxToEno/isexsFFqv5meERVf
MhJ04t2HsoxtL+DTC5/pmBum5AegN1LQ3S6lA7vtx0ekWnT18WSq/Z7Ijxhd/YlB
P32OY839oEzEnhhdOqK6q0RGdh3nzpi+zArhOWTA+1VZRRwT8zaS6Ha6d3zLEAs8
/uuaJDIqi77mGjlFywf1ILaDwDYkZNJXs1rQRr7P+Ked3J81xwd/yMVXWA0RQ+j7
4G/yUeUDKo2eJmTIl06yEp81/4OvSm4X6SycwJEhN0ytyctO+4gEIXbBAyOwicxw
Yo9eyuBZXy8ptfYQ2QREbd+5WIrP8hVOtK+a+Q/S5p4kdVzOaS5BtOgCSRMl/vhR
GEGsIy1vK82Ks6patdqAHQh3atqxYbCy7s2bEByIm36E/T2LxyP7RnYuUxkXC1R8
h8aUnHxAoOHMGTwozH5F48/wD1tajmShqJkqOPc3gqgptiujT1qHr2p+oiZDtY7b
TZNQEeo/kRNeSlgDuiv3+dKSFzZ5rmxq1Eu99l6sYlhn+BBONkjGMNsKFPkYbHon
R/q7NvY5hXsVZyDhzhCYAyDVBypm9d2spUIpg96692aypy2ky2MLXg3ezijHFvCr
iHiqRY2Kn7KAzU2YwHlXolxY+VMVfmMAm46ivhR6Fp1Tn+LBHBFFnvq/L1Bfs7xq
CXdC/ZPL9aryl4pyQWtoF3VD/Vk1dqK3lsAg4jlbjUp0Xgm+/tvYv0JjguIFgDOl
KA52lEleoqKlCEVkRRyzyxVCVnL0CdtgMeJqPhNfi6sKe2mmkz92uTApItbobfgr
TNfZTqrUWhzl1Q52g66waPQiia+I+a2hl42nVi6C8FPvHmbbdWDqiqhtUz8VMzHF
CfNakazJG/cFQcKBjZ6epm+8g7vzvNSmgb6IreWdFarYpBw47fed59i19achx0JG
48BA3jmjygmEKLAdXD7F2xfu6tMjBqeHZDU9OQ0rrTZ7ABy8WbP3H1sVXPKFVbtu
DFIeZMgIPGGt7lyiLFHDLNVUF2vjf6nJCWc0fKpSr4qQ3BA0UOBHUrLLufNs34YA
Ih3dx6wPmBz+Jw+0m12SWk0u7V5iEMebdCQCukwLk6PdOb+T8XdaaHSeIZ/WwsBa
2+cFr5CsiPqOy/mvtUMsy1lgetcVBlFAx8OQZGGHVYOGn/8mIYZrLXpRYgfcSiZo
aMP+hL304VqzIJoWUI7pYSYjA0PRzNJ3sbWGG+ca4tGfWdv3PIcl8yznnBc6MzHN
3QFa3GENO3a0W6nF4cpn9dJXgP4kyCdWYqasIzdtHr6iUgKiOEEJLhZ+yjH1tg1p
nk96vPShnVEg6beYCMhQVmDVakuFmdUHC6ust0Zroer2auFvRb5ueTRQIYBgbPN+
1I59ogXmZpZ2BYYpPlhK18fXPOMYRtccT8UbnTANSkaLoUIPQGspaRltIahuvPY0
1OT0/y8o5RfQligKzMKGykvKO6IDCobkSyYirqUywViYQ1EMrMFmJ6qbZKjowZUa
9DHkbseJSJF8pz2rtSoGRKa1I2dbARrkdJWwf6SW8ZEZ4dfyUL1ftrQ/dMU1hFFs
PttIMWVPmRfi1SmlKCW9wy5uCmQ5ZkusEZzbHY8VeaGUtpg60djQh1WjDPqB8PfV
C4diUACqC09D1XXFb4eRAJDeT+Hdq8fYQ9NdSsXMlldBGbVnINWjnuJWvSqa1Pkl
fW9/sQZcoOeFh3aGfL+N4NOaR5xW3NR+xwXe/kVrF1xr00Rpzfw/puNAnr27FJeF
LenUZb3BKoMTJBjOeBu11pZVN0p/8mhBrzP9jqZ5rTRBg+aRK7WuAJtCMH85fe0g
8NlphZvkVw9qWAddsmVIZytbX7q74UBAZxdMDkZ9G701X74MjL4Sz1V4KzeeAcU2
JSHvyZjl62HA/3ZAG2K55TsfC65NwMjMb/rzhRZkNogLsj9jLpn0Y2LA4OUY1ESL
mRJLW9rlcT9j3/cmyp522ImgKu/5xzwV5KhpTR08Ao652Q6FhIPtOaBumkF+POaq
5HHbsyV0jsskP1aa5kSMbp2edE8949LfaSlVnMkKYCfJ6TRi6aHXBVZIZqx7V18l
F2uTOl6SC1ah721lPmTLza91X+Db+YNrx8Obyrasy8tZrqbV/r4soB+OeRTzPA4n
pK9mdNBR+kmr1Z7jFMq3I3qec/i7na5RVHLNyRVGD5cdetMEud+X2oTuT0kgTY9c
rk4jILtY6gbs3dJoNfsT2T0qo5k4PZZoL30gbXqwdW4JHUjF1g9eUa3YJ7I5ZXsp
S4WrkayZHX2YGZWH+9iQeKz7W4IuZiEd+acD5WB8HstRnwVoZzSUECh0ZbNDlmRp
m0RSzWFoHWaqR7UsBya2n6KtSI0OjJ4l5rSvyLrQFrC+R5AjV4ytXoM/DY9cQM5s
LQNGte/Sg7QKVMV1UchaqKmCZmBBIGdtGOKSOUAyHr9bgFjiuCWRLQHyrM6AP7lZ
FoFIp6hfPVgQxwCK5dGghnknYx+mbKabDI6mRc5SF0cTRz03QNdqlUaTS3rrWpbC
TjFISY6hgUMg80nk774h908JE1Ea55g7cwawMea8uwswP6hwCxI+Iakc0FecP91m
wBTd7IUnBWn6dbWc2/mrakaKJpw81KFx3fVwOoEaRSmUy3Tp5FNH0myGHTV1wz2h
ds4CPKFA3hMToIJ+QQ2wnjncg5+JU23fCPDD9DemYAKolFgLjvyK4+Mnmh74aRJx
Gr2GeQB+qXhXk+nZkgVgU8iS/DfUytX36BfnGqGGGbvyPWQROY+uFUXT9oV2s/GO
/b+tDpE1fVr2Vb1CuwP7/PORugINV4ROtH1SqTxJA2BWrv5fjTjInDwSlol/40LJ
ruKTYDgb+JmZWVACerQM0fp0s9Mid9E4wO213YZxDCoYpsNf3YowVnnPAgkpy1o/
MvtA+I8MyawsitYVqH7tGKjb+Spr+at+8s/BTD9IVrUF6Uw72zURCsBTmaeCwBuk
ox61Eo5SZ9cwZDI+tRKG2PaaPxGicGflf7V6b5LtmMMlO+CRlY60jbNSP+KHJiCr
+A8RUiCShJX7XZ1I/mFh5uDBlBZX1JG8B+KnY/dIFiCv5vJmhJT6hy37ZS0ndKAV
8kp4yL+5hgC74yty9IRi1BTRn58qB1pxMinD4e6+4UQ3Bk+7jzLsCaw19335dAjF
AByfuhBatFvBZBt7uzuPfD1kC4FZJbGuIprDajVYPq8CmY/L9zR5Re4tfTe5cKOt
XpNoisXffpGTHZrf5JhmaNWbREUOsh2LYwGZ43okYKII1EjflykW87gYxm+HoMHi
EQL2zGnQhqbfZmhhWeJ+/GzltDUkED+Uc79sgtRFt62eT/JHZuBuxIfFQ4GON5SD
xIua2XVgeHmae5dSkLwpsTD4NbSUUB51rWZlYW/M1riBF8nfONlBbicCzYsglLB0
EflfwgaEKtEfMPlBY3FJjUBeOb4M5ck+TUrLc7H/rUqElu/lFZR2Jn1t5L31nlRh
+Xevvy5Fwvvn0DnPKJXfHeOhcY+23Kups1+LaPHXKxIqH0jfAa2XNaIjdPOAUXXP
HvuLyvxj1MWgLCngnTBzcKDc570uew8QQ/lAlft4aRgtw9GyYqx0eCRJGKUA6cS2
09HXK8ar9mfZd3OhIjCruFM5Z/N/Rr4w1d9mseo0y3CIXY1M2nHCxdrx5gCvucqu
OypjVbCw2JnExOat9004oi0u6md5UwlGn8dAlNhMz1IWe3gJPLF/I4QqeOvs+gEk
1sv6DQ3pdgFkpDQ84sRRMUWgWG0U/nm4/bhh9E6AEagl/y0+nZXGx5QzqKU4DeCA
b51KEVpCvI3NLd0pNl6YCNNujb1+bF6jrwJ1jIiN2oALW0q0hWzC7W6MSp13Mm1H
lK9iMtzZXThATDXXsdBhPAYCeHWL1ERAFoHY7IuoH/TQXGCyHiqxBkVegPNk8Z7k
a51O5WeTgdVH9A8+u+Xg2AP12lvY93zwe2OVFfR24KQjvhdWlxNyeB3KPzbiHOKf
R6aXl6RNWDwNuxm5AeCOl9uL0numiKzysBZMAjfstKVmwk0G98VCTnA+rpp1EnmA
BuCNd4wAET9pDcXGP6VcgpbHcfQPILeOT/KIhzXyy1YHvo1bBFOPLbxjNW1JWb89
MwD2KedSXop0vY8QkGC/HDbb4EVzDKcB+hdu6/897CVpq85SYydJhSs5/KyFUWM9
qI3T127+MKFVjtT8sHvQAZbkynpJYtFx/q8Vz/Sks7/SfsQCGH9yeZcR1T0QLMZm
80C5LFgUOR4r0+j/pYPgdw5rWKLL4sX7K/viMAeW4Zb/3up0B2icHZe40b5QCEzO
NFqeOaqLAXxhXoXSBPwSffulwV46QLDFIZw8JkCLVlD8BwqAY+PqYhcAbIwYLpfv
+pOuh2TBUklKF+NxWhLLttpNZnF5PBa+fNyyuOQ1SAyBYYMbmnhjV9O3tI5PcBr2
gX8jLSyOvvj/DJ+rBL8WlyhXujct1eYtYhnbibl/j8VHBq29ZGExglBWbGcVN/PQ
feg0dF+Fi5r48v8NPCLMMouqntukX8EN8H8kwuxtgAVGgBcoJnhnDO0EscFUiZk6
SureSTz95Hk1oGzanKNX1hJCbB2kxxK8YZ01zPKGYXgQjgx5muu3oYv/zllitZli
CnbJt8h//zFA5ijk24unLZM1jAhb+aG+PcMgWClrRxnjotiiLu6N5mrpAz7mb2P1
sYhCVqM30RH7mxgJKia5g3b2NXoV9OTIcRtbfEtegnmIL3O/0nv9mp3bf4aHSsHh
Wdx2FVXLpcCdedSvX9k8QEVKwKfMyFAz4zUMbcadYT/x/KZafCobA6FTYj17hGkg
IGucev1Jw85Zbe93T9c4S4Ln77fEdTkVrY/zutv72IfUGmE0OjIcJSdpULUuIbFh
UZITVHefade2DHvq0Gc0Rab71dC5JBEGS03WqSfelDrFTbdalo3jIs+q7a9IIUHL
fkXSj7a1Jnh+ywgQyBtMXe274oMuLwrdQHOmdj8hDhVlGxYOub89kIAoVMGmNH79
WurBHHqkPlvMSCmEgcpZmjOCki0ilVJu49+kdwfL4v0QyPWHMHdssINs3FNRKdra
bYXmf92jM74h/uS2QntJC5J2WI5gQydIexYt5F46HvivdfHzKnpb2h/3j2O334Rt
w3bs2bdbU45FkS4Ay6KSZzQrAqGh2qWOJ89oC6QjB4k5lrzVs6apavBaxE2N8W4A
EwWSPK3KlzDmDk6dVFa0slsZh0hqcLKA0VXknnN0Y5gxVRmGYiu4euOWpEPSqsJJ
e9UTWwGsi34D1RpU8RGLBJN5nxtyBt6fTnvROxaygfWYwZbaT3klDLVTXNnZvArd
P9M1gEMGN8EUSK8mP6ul/vmcPwlzRT5zBpcDXZsaVJJKYlcJmB/uPKjCbygjFPDz
Gj/c4P7vvZbymlHbmu4PzF/jEQXbG/Q2RtfhTcQO/VqGgfpWVpEbtJAGehLZmpl6
5n3uq208kpRi2i6Wf5nDeJlzS8MxgLD5Ph/aVWJOxe6bg8tFRzPB35Sts2Rg4fVj
bHn1E75nDZCAWEg8rPeqLYSJpIddHUPlq1/wDTPux1LHROn8rrWJxloyR6gBWaYX
tgCQXdfp2jg70zQFR6vaj+tz0oaJq/80vEO3ySlsd3bwNnrqNBiV0BtcIHUkFT91
jYZchRcZevi4wTOZV2OUxdHb1HMPQzlTHqu6IBdLsJ3ex5XSd6q4PyX943FqG6t0
H+tHn53yHWQ3fA0xhUw+P3Skv0lmeoFVle5p+eq866ecEybDsodlQh379/tXmX6T
wJlYeSgfwe823oqpvtNWQyvqmIimaxXRmMjKXOhou/ULIqbhZ+AYvg7W0Z02/6bX
0P45d23mGaSA+XkWBK6YhPMVI7VnnaVYQrRT5m9nrt01e0KzdjYgp+yUBZNn8BIP
NIG+QC+gCaRcF/ph+vBmAUIE8g/VDsfBGUmHQ7Clo0w2eJzZrIume1O26BZWr+9r
NVfMwHJ5+HllQeCc0Okaegh0Yo3Tnm8jQZDU1Jc5Ia29w0ydbw04Tnm5ajOlbOav
HPCYd2WkGcQDvzManwvl/1YzIYts883wmmSiuJiiExUBwu1z4gGkiHD8x7a4llav
a9P/a7l9Z1wTtoOw89Efy6I/TUXOHWFs0cTuQeAZtCS+G5dEqEFRycoFgPlU63nL
qFlXKe/KnhbL3QBc3V1l7pYyVEwKG94Dy6hVAD8ePIRM8L0R0M3AGGsCEfQgEugb
lJNDHE8a7lHTZvSn9hhuus3kvOaUMW/bZAtzvA1uXXrsDCF3OPqSByf33f2mtXVr
tB1fGnwOotKJ16QXDDykqQx43/haCR6O1hiNf/fhKECf/juJdIBgl203G9/9HEtZ
oXeMsPt6WBFWNz7nevvvPLnvOUOcVV5em7M2hqTypQA8BaR1VXcnaMczCk8M7ymK
3g5JYL+crkIXfBTFUWBhTsCDnh90q0J3u7kBFSeS6nHZHmxoj1gP3GS3rxgPfqJd
p1FUhsu3YjD4W8triZMA67qjwcfxjF1cjO4RNJ+wRXBSlOaOAS2zdRSImewKoFdC
ztN5cpD+2PA/UdBsArG1lYH1Ooir417bnjCR073j9kFxBeXjWX3z6UMypsdYlJtx
BqKihAWgmPYReWu/3DMpKtrsA7jm7L9+pFz2/XtvnheKRNUZR+EWXCkGq7gxli87
Tq0QXwDwlUyzECqzxElt8AabUBWMrcb7EYnu+QpZR8Bp1PXvRwgwXFJxFEsCbsRZ
Ks0E9K0xO4fSyp+ZKNv9uy8914D182I/oHjo56EC1ssR+207tl8hPFL8Hksmv80M
2Cma+5h0QFCTmEbpA/5B7JxY/ecV1LZGx6kQ69J+WsATUr3dROKyc58/Cz596zhy
HST8RFxKgAc6LiN0zpr514GyX/O1crRSXIglOP1aXz3SmNYP5dKk/4tp4EpB/Stg
ElgKrhRhPsUVaHM6MDwgfQX+K89pZzaUDPKyec63nQeAHTdEksycZ5x2cBZcFFmh
FtmQ85WfdTtMyoCX7xB7JQaRTBZQMwT9oHAnRGl6OMDhbGkGq9ATJwcEeB+lIt42
/r2lVAFwUBwgiqT6TM72z8z09fvaWaObFJ8IEwOPzraNLFRY0UyZWY3ng4lg4vjT
AuurESe5lWpNArUbO17qCP/ApHv/rLMmOc4vahVf1U4ShTQOznqv8jifKyUQM7Ld
v4s7acRUo9sqo9syMrUbYQDFk+uX597+vQ+P2/eafpfSzMDLHeEM8L3GD2Et9ikI
N0XMpZgAbRhsI6Er7Q6r0GpKEGx59yYALUdiUGEX2Hih5MzbbMwfYBTrviQVF49l
BK4yCXXd+d6yXqcHcc0izd1wuXtMCDwTe4KkI2t/V81cfeEptKZvPEuIiik6c3m0
ukqMb9qjlGJnM5EC0PX5Sfu5wx4tpi5F9ak1ZiNIg4WMrH3SRaAj1hsHJThArk01
km9M7bgKj7Te1I+W/EBT0sGZEu+LK7MQcaB2ZumdGJ5JYlAzagQbgihRpG1Yimwx
vvV1UbM+EWiJc38bTd0aM6U7kp6QTNRBTM7zqboWYiuy7fsTGonr/pXqDtKqUVUS
/oXbrbyAUqw6yDpgAYi2gH9HthkDewZZTv8Dxe2ZQfsz6/ZRSr0HuNxa9poKWeiS
+MAnnqOqcurZmEkGY50gzlacONQFh+Y5grzIovbanlTy5siFKtEQfzBoq7+7hvf0
CqCoDVAEPkBYoZSz9kUohKNXMakLoULCLwbxi0KULjmEwiSSeEsqnrYEz/2wCiZr
7og3IvKmemPg0xkZ2ZYNtLXkCkqv06tfGLjQz4YFvupKfnalNzkx85s2ApEb0gSk
D4w64PRjneFqtbVT4k7jWQVej7UunX8AB27z2/1GgyqZAsI4805Vc8/7sgo5mCTA
qne+9rv9ViyfNT3QXeC4mUcbE82H8qG2GJ0kaPVTv0KPYB7uYHCM0uyBmQE228Ak
arEkqn/3gZFn4gJCTPE8JU5CWFLvqa9xyrAQgukRKzkmdV0Mh/BxMMH12gVSKe+F
EGgHyMl0xCZOTTqHLpkUPBtobZj4JruE7y3XhZ+jkugacgBapbR5QNDXfRQTIk2z
+Lp9ZvC656A7l1RWbL3IGfSb3TxOhaTzCvQtm7ar6dqvdLcl6JUuQfcpUDshGPeQ
ujVUR0D8JwTd5SrNXvqVGwTqB9zvHYTRo3jv78Il2ijVj6IKwOFAs9A35KkcoRfR
8d8ne5I/AMVEntSVjFYfs4wETihDZbwJNXlvn7NkPFt1o5lJY/4t024Q3DL0x7+8
ep2VFRlfXom2bRUK2HEYG4MfNNv4BymNPKCea5c3Q3v8ZQ0iG+3Zr6MPb4g04FVa
6Z7VqpTeR63RWXEOzW4agb0IbLPvU1w6HUVtP4y4fIiPMkIAitCcuvYxmh7GNK1q
a8vemWQIAmk4gclb5x6Ut/xxPAwxLQUl4a6hOGhX3wyrMFM+WnTyS5o6Wztp5tV/
kf1edvZrgGjGBm0jK/O3d1squEhmTdYTcyazyZFyv8oQU5VIx3dWg6ETXj4ApwOT
vlcuS1nLV2mt5ScBMTRbPPRtGuNGJMpIDy5lzD9Q63h728u5KhiOsZuKJyWzzu2j
DVIANlXct/3JTxEhZW1ytIg+DNehVh3wntORyTbYp+0AvA56uP5ZAVmb8shwivKi
FC1nI/cppf49Pub3bzszhkcOHXp+ILJ5jn8kqLxVYhLmKNJubGmTtl6A/kWECAHY
8m9qa+cy5VSbOpyPwY1Z111khVFr8onNfNyYGtwApVqDtK42O0qNk4YmesYTwWod
hnump6lUnCQD4vi8N585OuS/zCl0IlSG39mG4xKfGNx2Eg7zWRndgE5G8lC0+Gm/
mcS3Z8/q43/BzrDbgIqUsnguQRoXUY8M76ZecbF+7fqKX2POwCNSYWsPTjISxH24
u0PeR6R931s2e3CbgiVTGQMBvv/A27PXAVOsupzD3y/jkNniM8+CAYiKiQ3JRsyG
MbKfEbd5GSmYT2qQBjPedy2sbrhpthK1HkS62doYTEqdnaqZYabFtX96WKBXIQy/
3BQaliLfgGHJJ3eEa20Nm0ErsCGFqd8bQ8Anizf+jPmDMDlgpRpmhxCYUO4SPSVe
XMAVMgwoUNXPaeJUzAIIBHrEXx/KH0C4Y2OZ21A5fX6qscefdAYtc+/1UUcit3dq
J3XBp0pmaiUpkyUgxUj+4lUULzqsq+BA/kEjWTFwQ1hoia8UPm7JMOKy7EViY7Ae
gP2TwknDTfyINKvIJAGLnkvxRv48zYZ8GdH2Jk5RThWjKCXiQnekC+hDshP31hfb
LCKlz9i3bkYhDwUJCWfjwjcBWHpaqckbtzvIgjm3dUFl4bPCuuAoZVZZUMP4KSdb
Hmikpig/UoU4TaiTc4nmCl9e+04Y2cdzoiyKK1CFnF2MXJk49Pf4XRfMbJJlOnj5
YjW/bxtJJ1Hact6IxZn7vhWcXrr6gqoFfYUnLrAbKdWqVzohhs54jkriTpOQZpAj
yrmAkAn2tDX+TJANqISGfCnrc4zQ6UUpZZUOsBRibjpCa/p8r/pnL5jdCPJW2GMy
UkEitrCOH7/kOKuP4ZehmyxX6RQATnGFJCQYfvNNOhN41qefy9+ZCk2szOSalNiY
CIcAjBaCXAXY1JfJAQhftC4Q/1vUe621byipcgJSwaUF9mUcBRKMQrFsOs44k3my
2z2Z0c5UgJXflqasMSLkh1/QX4GlvnNlEVVJlgODP8VOsEeVKZRjk0eNnG3fQigF
jFuOqlLWe7x8cZx4eItGaVRsbasbcQtWeGGQtN0cnpFjsH2QBqVrd6KVDiKYfBa2
H/VMn9fKiQxHINwTUBWEznMuJOznvmu8Srk1T9hRv278fIcd3MWcL1hC3szFomkN
K3Bos2aXlcrH37ZGzrXlUAzrSkeqBoH56ubdszgfUOlg6Wu9/gcHXMy/yDz5D96q
QzdEaOElAM2MeSFmksmpGBJHccjrZ/J5s6YaGwP5ptOPKA99ZJGGOwntslaJaTmG
m25J9Yt1jLW3aqZWJwallhRzTD55U8dk2kxgOU2hqOhEwrFImMvOFudDrvxyeigj
+Jfx3k9BQE2nVZVhhYDcB+xS/rvt+BTFlIXK/OxzdigffleONiLNEnECBTrFVke4
9vXDyIovsl2sXyMZ2qIERZmVQ3XwF9lVd0cdsIRt6eiAmvyiPZ0CbrNSu31SDGv7
RGkvtPxOariYld0Tlta26nSr5+hO9zoAJp96B3tTQa7fmtALswx5oqmSu8fso2FC
9cMtTqgE0081r2al+GdvUak7peKwYW+ldzAOU2YSY79ouj9fYPNhC5JtgeoEwGKr
anc+2fkm3bdlhm0Ve3cO7zMooHiEQOy6WLnSDC3HxMfuE3kCf9mwIcCatd7cD3LV
KZCWGf1opwBWFBlmOrFMNn+amt0qhY4pXXo1xGzFpA/gqDPDoY/NKr7QIIFuksnD
ASnXj0TFM6/fg9TH8rAy16mEf3tw5duoDtifjHR2tcKOO+FyGbf8EQnwuxRp6Ges
AB/k5oY6vxm7ytVd9EpVVcNY/3dgpqG8MAH4UbzaEKTzLQIX3L/pmmdnG2qyeQ2w
GzmlD7b0XXQaGZfdwT9K97r9Wq1/cbYC/THCvZlAtYsqO5IV8qfPER+xC8L8wNs9
N8XmZN+lBOUCOU+4XTC67YGB6xYH3Kv281lFGMYapdOyEs+U/xzAWM4+KHuPkYYI
ebc80GF4QncM3AlabxW3EUONR4C81ckTIlxWRgJQhsycg9oxDZAyjXQ6OgspdsFU
AANMy+FtIJA4jhgrAGmNXa17vfj714uCWGl2oungM+fRpraXoFfSeAn+Pzbgufee
WaDXwAz9qpgLPfj5bFH32S/tnR3UTCbP4MHjkfYN9kjYvqbGxIn1S0G+KX5dFTiI
1uFQ0ykNJZ4fKsLKFBewxrYpf15+XA5H3STS/C9xJjhxe1X0mrewIGtyEci0Vfqr
tvS0yQK+fM70g2ZuDKqgkMAySp0mM6VHOKK8aKQSjxyLT9DhS8+AnbpKrS1446a5
r6pxLQ2Y60eGSVY7cDU1vBHUXJw2QBLSXEdtcZNE5kG1oRWeH4SdCjhvg0rq9TIV
0WlGV1KDOZskcDQyQVb8+ZGWbSBC5k/lu20OtDDcwSsQeYfp+qHSBBV7LObiaKnx
m0wAbOjSuxJA6bH5aCoZg3XSiB82MRZL9qR/BQO0ULlsh/wljd95xh6UX8rFUH6L
jOS5UOK1j3HhVGU4WACCmlSfF8nb4ptIELasWuU/uEotUg75UK6oeyNtERvYU1my
v9aHCSpjab2ylMO/tE4hJni0fA7iXJw/TPc5J+A/MyKQ3+EpGknWxdGYmtnshKg7
dALIJoZ3GwSgUb9Qd5CFa5jlK5Mz/kdfxjnLkQXae9k8Lk6ToM7QD0xbirsqT4bo
MVygUax0lGYk2AMmONlO9LlRCCPA+bUb8vXwdYed6T4AACED3NVt1t296rjJSX5J
2HNq9m5/CZv+K60wEY+Bt0R8x63cga9h/BNZ9DpccMCVp+34TswLrnkwPt+CmO12
k2GCuCb2gEgHrrhLDOZ/yYiUhwVkCYqtxha6sSJcCpdR1ZXIDsC+LeD7IS8HQv9l
GU73A4teTu5B0VKc1Fl6q5/ZOva9OSOZF5H0BqrNGqcMlOJWhT2SPH1fv9cfUWc0
nusyzmMI1o623F603pQre/AY9Tl5wL4DBrnXWpMPPVSk2FfZEoZ8r9vptfvy3wtV
BZID4Pt682SFyu4//7PP9fEGrJE7IZ7kVU6Mlz45TyC6SONXUNHs2x7LISg2mF8R
WdNuox8tHkUX/FKPx0+3biUCUMY3Cp2pxIUGSb+JpW4SyLT90UuygWZAIP7XZTnf
awXkDvZrwrBtwHBgjhGyK7GdBHmSqYOK2CBy48o6yZPPas+JfKVmX7XWl7VSl3/Y
zw6vpBwX1FnoZfqASceqFuHEnUba+7ZmfyK1dlklB7NUZukLa+QMYlXYi0SywRXo
pTijieUbtxGgMC/EQX7wuBKeslSiDM8gQqMeTcL11uhwTDN+KWVdt2xOn+acKNNm
wLR0qMj0QVQgKVTWdTa8pFV838/z3miLao7SQ4BW7zKh+j7WT+ZzeThXrupUlAJy
H4OMu7SbU/VjPcghZUxeD3O0f0oTduWqME+7JxinV3gWxnBpO9N4wcKaweE6Bd1f
eza8x55HAQpDDCwYyWe5MT0KvWMnJu2yDEwqflDxU6Y1aTaku0rzVYj9DY+6T//o
c8x/NpCi8/5HKF+Kc+TRvix1qRYNrDGM9qofxdaLWDNja1pXnJNIa7qxWeMmp1Xg
tn0tMcUw1iHPS9SdsgeDFeq/FFUQjhH1EheOiRwRl1TLmd7UTi1Q9IqqAbQuea2F
A+pm6Geq3OZASLvzUu7R46ZL556rQXCXZ5/qVZVZlTr/YbB3Ibu2XyNaZWMXBmFr
8N9S6TLfYzmqNGrW/BalGrRkfAIVc896epgr0mwEIb4Fel8QBw7GrN6Jl0STht0Y
ml1ZHCVxTITRBqQ8B5ie/RBNl76j9m0ogxh1D2kkFLA9yulINtRRIvfv/ruFksOd
js2Gar/buGOMgUFSpW4iYH0rXjkPx4azFWC01S2kNq9GC6ZUxPZq/qVFbJChOiWA
4s+BHr6auxLesGUkQsK215cbzS7aIaLPlxSn6NLfofD9ZiyJ1EX6DRrEdRy6AFdx
yPhvbPsNm+2RyXnLqwkSwxqCM9IIoFCddZJ9Bh08OQmvBY66dpaD/64/4c+dQu3b
f5mDScemU4HrAAwYm+jktt8DtLtOooioq9WjTY5u6WQ+/L/25jvI8/m1NdzsM2qm
bmAX5M35v1WFen94oSiqiXXmqAKPRDBXkKcd5YBqwrTciU6tDdjSDb7tklygld2Q
blv3y1e3KL41m75W8SLKPaWnKvpuviyYefZOumEVh5Qomr7yy8pWblWO3GvD5IWK
WA5ehjQ8OwqzOkhEMW86JZ62eqrqNnLJt8eYpa1FAdGC8+LbWjt6VuGTLvYoRXfk
yZJMODXMKP78PQCjkiF1al1sb9qXO+2Xr0nMEftnGq44vYS9n5s61BOFN07JBf0c
5LFri5tm+RS+P/SuGTY4fGZ7aX1ZlN8Zf2egIBaFEqXdsdPnzt6gLSR1XmOFtTeL
pS1q0rAFowPqhHEc6+5uvDTaB/pjlRIiJR8HdEaKHUuHz5V/LZCHkS8VPVk2xqFt
dNRzHzcfDxSeJHwN1pSbBLsdLJw3NQMy2P64WiOUURPFDS11q6XGGSsG0T2uG8R5
7xMLAil4NQlloZiMAQCkxi+2l2abBxyi8l6AvGBklzzrSEcu0YOjurkJLiJ1MB2I
HaGivqvHWx/eCwJvMQaicr2KGLwHBLZkQSel5LdWPL0V+5VZm3J0Uj8dGMlrPU7L
cvJ9cOb4Z6UfR/cUo4QsGuaSgbxupnHYavk6aTjk1kCOlkMx0wdUL8MDIngL2tbE
+GwG5pqweHmDTU3eXiOkQTI4rA0HGgIe454RDLuKiDbGQteI8gigl5WYZ3ZD+GjS
mjhf48X3dGXwAh8heJwrOjZp735iNYyADR/Bc/qBaP9LBNruNZ5bCcP2EdBEeZSN
N3sX4Q8Lm0PRItHMB5RLU8MYT6rX3Hz6lzZ1U/KtFGNzVjoZHQiMrX2tbcu5VlKY
crYLEE79R4KA9npqXVvAQ6eCNw9F/Txsh3kdwvHDp3gzfteaautvV1rq4ampPdT6
/K+BjEGP3i+/DoPyFDYVjOW8ONkD4m3vd3H+ByAhdVdbg6DGKHugUvpFzucExK06
83hJTQDCddNafMAv2CklE7j8qJApMLvBh9W/+Ag5aMWN/eZ7pfhfVHVbniPZqrkt
YTDqkY0baKYDaLzj69uGaJxcy1JEIDhtoY0iNCr0vxDmjBxOWKt4pYS0zOh9HD/G
IH8NxmumeQ2Gi05nZEI1SvUwooM5WbEkYvUwbLvcTSDCOljAdIR9lfD2UYv2EdZp
j7wPk9+S9ufklo9XStGIQ1g4vkX7HHxPDjh/9Cml2CJgPF0pFVB3dVULD4jfyVGw
bNkvrX4g264ed9Y4i3uT94XL/PJIQwQDWgW1Igh27trekeOT5oghelNSLXcBC/9z
UZt8LQFYjVUsSjvVRFbSBb7006rTlGn5UpakCUcJhskdrAsROvDCFpBLoGNXGGL5
DQRsad/AXaB2wF3tmem8uWbl1eKLYcte792zwyRKe/eUxKnGt/YNEZ+BGIO2sO6l
tkJko4mASPEUlHIVtppNJ/0re1Pd8EqKFPGk81WVhQKI6luOLJEVGA0VXovOYpKm
bymWnPQHQuf2NB2Akr5zris88+alPCHZQ0y0QPhKOj+ivn3LUfw9WrKcsCFBMxUH
hqBzSPpGYdWSXtvRp0Ug5Vzi7KM1xnyFfUD1gmedea/jr8b56iZxshSALO0NIbXk
FZsmPUYCTblzbI9g81YdehQyQzUoWMwmR8UDMr/bkXUsqS/VNC61ktbcXaqeaX9O
tUNNGvHejlQ9iTfBhH89ILa6m90xScSM37Jnm6bFT+5SgERyv9QCexkJ0KH+Tkwk
SVWzE68GUmObIL1uglloL2IntR6JEYj/BUiK5p1EiWifK+bEpeXiOqGb5Aa0PLLd
bKZilQLC4Zzs1fv5oaw1UWv5HsEXJNMiv54r7RD6a90+e4esNoT8aPvBHm2jQVqV
1zMMNRCmD0w7ft9GHekcE7pUX4husftXtebPeCKDexM5IX8j8bgmKvAhT2SZVPOX
lGgk7iC4HoodflJ5roHyt/juY6zH4Wg+vvDjILliWPZc9HNbg2dhw3hKFMwsN2Ld
ttibo2F/cSgnN7BfEepbTP+lIpdFv5j8Sj8vm0sBKHu5nXjHMem88R1jK2Gv+peH
k0NtNVbFK/T/mrZWinGCCi5LfPcDgZOzZ+/O3Q9zIaWUmbJkOX6qL6eyypaspxmS
P2G+TxfqHNLJlIUvLbhSTy6EkZFGnVOJPxcKl4DivDCsFq3s1eG3/z+SdhETKJ+4
VcNCVpNf81RsIiPsZM8PrWo82U3jWP9W/lNTwGloHD8cpmTW6SvDkN1/YyVIXt2s
TitJKBJPY4MQROGExQnIR6bYmldsD5VIUzWK590rM4eDuCRsGtpqwGhcGssZQTV+
4SB7eS7BlkAhL4+OUK01T9Vkp5Qlj3zpqgZDELfQhstpA3vUTnXJBgH5/n595t7V
3HCyupd23jHDPI7qiGhF3/XYbTiKiPrjIwDWneOxZ1d+dFTezj906SDlEpSWDUxX
NTpKp+I6UXW63ZCdh6qA6cResBNIM6Zt+FDQkKcbci0cWsis6l9oiQwRgUOjtgY3
b9UQG6IVKMZ+QAvLKatg5fPP2cpv+JQPmB9glhmb6PT9qZQoSNpCGyn/BzX+72aS
MyVvmAJiTh9z4oIlmiLhyD3Yb5rEIQQ4MLG8h9jVRcyez0bDNHSVvSJWgDb1JXeT
+j5VNKFIA33BQB7NFr27Z6Qdhk5MZVRVR8tGMJ+l3Po5R9NfRTwMlgZ6M87gq4Sv
hdeUoNVyBro2EMV/QuUuDz0C7wY7ngyrmmEkwcQJ2ijKT0QGo+NG3Y4jFXKzzmQP
MEfaWawUMkueUpJYIqYbRdjoO9Pi16/oDU5gEtDhTp3eOQ+Hdwl5n9aed6QnFo3f
Lq/pO6hJQDlNgYnGdkK07jT5ZzGRVUODi/bno6zX54T/ARHj1LuqWmL1voc0/gaI
NU+WW2EACKB61DhqtVOQarM5kmbafGkUju0+YbiMs9igrougSinEdgzcA9m/cDVe
k9ch4mbNz3qZi4JTvsZrs3BAQ6HsQRrlAjBCJO2YqbItml8YORcvpZr08+g7xZ2a
jYYu+Y5NrjrvatrbFWtX358lJMgtlCJoQb+sdMXkl6vYfyp0hL1doNc8u1lhVAS0
rDHLi8PUgnldUF0m5lS9hWJFeWeyTWE6BCkOnqSDeX3iywcz7k6+7IudkMt3n3uP
cfKLvR6waREaSbzVYcFZ/CxbvpMW1zYYsPu+YnRn889Allfb+Sowj/+A9jIcUCw2
JccYnEX2bGfcUyM8URF4ZUNekmLgDsjx18HSGLkNMX4iGmVL4JYP1ndmYQq5IpL7
NBjBLDWWivDJmQgNuteKMp9oHXjTMbH7nb/tbvQMIVjNJChNURQEwX5ugtdWPDct
K7Ux17TYiRffaxc5AVHu+MDFMHTtyW84RFGEv2NXYfj2JZrB9v3zO9bDrucXHSLt
bj931dv08oRMMFbienghb3Cl7PZX+5duiqstbIb83wrP9cM2qzY9rmJPFcJ88EFY
Wg8G520SNpbSLYobrJwqTe42Ci7AUMX0dbh3tKexxvRr+C/pKe2nxCGa+XwcPSmH
w/IJ+kL8JHIa0tKzdHZtXqqyjRC0c2UDsZj7JGcAfPtZd1y51gUdKWWsOz6EkoOP
JafoLhjjlHQYBrKVbbdL3f2IYw96JyRlv8vy+lJWCi7XVVWprnOwqG1UGFQTqu3Q
c92I8nqxJQtP4qfEnwJe+Gee5SNW6LcpqAtvkLK+RWSQDdQmJTnof3Hv4uBS6O/L
Jxh295JtiOrcBaiZ8F4eLIbuZ7jW2t6lt/d7TFB3zPs4JsMlNyt6gitoj3QpWV7c
IiCxRysIf1SgojvxFGyPRzJJT73sX4aO1rrACLNM7H5t/urfDdKfsbwYaWrlNkQa
daaFQ997znTPfbE1cfbKuSUcJF7x087kGoQdI7PhrhW1e//GLi4agLZ4LYqmmD9+
VnXvBVvc/s0OiXspY0DSnGacULSkpXCKNmcgVRJh3cbnqYI5f/q1XB/RUnPCl+Bd
wt3Gg6aEhL/WYt1mbURyK8ipXkxVyt8Iwgtd2p8fZOGmZIYc1FzXYDDmAQFpFz2s
szd1UYCI1XcXMoNLA0JA/qzfHvut69f9MDtzzVyIQouUSED8t7u+dzt1KGroFVeG
niPkC1u8wMrf3rMZaCfLI/hyVWC4zJOtzymqV3sBbS5yRFE3cj1ybjOzAO8gctEp
juwqb1DrA2dEdd3tmNjDOaMkSUBq1+M2CDp3mDucgqz+qWAaaHNic213rQjvocqJ
fwbv2QoNoyh7Ev7Ui0HuFdM6Rirz9fSCrMmW6vq02o86QyTJ68l9F1q5RVf3zxNZ
2eUlcWm63RiNt+GA7nwr4gltfZn27o/MP8fAmR+FIh/EwY+ddpgsjqtM09a215Qr
aWDwPm4qWehUAKLvARMVB8KgsFmPBFbqlp2o/P4J6cVuu4NzrTEa15IMe15SVmC+
npzRiO9coMeTXT2slQtlpXUfm5z0sBqddQKBAppc2Uc3s2OgaMjkHduG6nYYCwAf
gWXUPE78xbt3caLwZoW03YIP33B115d2LUtc3s8x8nKK/QCOfm3r/4yHtP6/AoZF
G4xeXoTvqh+nOQBLiZ0KIPwrGZkO8L3GePXKTFbcHlsHIMLkZM3DvdlXH5jOBVu+
1jTxNBlrt5tXPzIB0AeLg3D2PHxW1N2cn16XN31omK5seHn61CtBy6IU6odlF3pM
SxPPNr+BaaIrPCUYc90NO2X6PVtR6i1e7B6eaEphvP25fOAsAMckgoN9eHZpM7Ic
6ArIMa79CNN/Vsyg+/zSQs5LhuFOcwgvW8NFy+fGSHIPFU7AIa2OfJMSNAgypHYF
O40Q5HBQkxJZ7UL0I/tXmxkvt1hPIi5lvIG8TwXLg8Gjf2hrkJ2S2oY3CIKQWLK7
5g9O2JuLvZwOncWePJTgd0r7QC6D1E8QhNCMzpviCFeHNppyhCVdKtUfPVLius4W
2CWQNY/+rbeUfhZ0Byyhx/oym3soiHiFjblBZzv/+5lh/AzjZpI1a4x/na5EgMJH
A2HhoXLbiKbmm+gz1uunj4o+8fiyvonq+3HUBTT3FZZrEPKVMtQt5fdXXU79y48l
OuK07pGQ1xq6W3MCnHwAm6mfWEWICrKC+bQAIv/RaIxl0ZZadLCz1X8m8/b/H5yX
AsZboO8Y38Hfn/oR6v45aZb2QpYCeXkTYMUpWjLoazIw8JiQ7XJAXquXzJBRccMK
9lUQuUZQxceZBq4E6QI1tJuhyMx+t/YJ2Mawcy3EdeOECCJSTnSoOb4DFeFFiLty
IvUiWqRMVUtcZp/jf2D4tDDC+bheUgMH5bO+0lWalIe2bmjqt9YA20yK9DvnnGAz
/zOS2qTMVFlOUWGtoAV3EcTmsSVnhNw8nXa4wRW1Xpt/Ryl9soyOrZrTEf8A373e
d+ffKV1Uxrdk3aMNnTZVUVwZt0L4MIHWm5L+EF/BbuigVih8IPV49dj5XkFFFs+c
Uf0PYhzD5E6EHlhXZft1KRb0sbQk8OdNBZNzlLrgZdEvSdwYRZwiYt17rOVw9YQO
hLlcE5ZqW5yDNkEh8ygaqQaJwP/1yKPClCTcwJZTsCzejaEBC/JqXhvnng1oLmub
RATSYRWGvcmSspfwp3ITU+m/AS2lxEu995NOgshK95vUMwV3HAS+dpQkU5eJ1bxN
/5BH/ZHEe8iPiDRoA1zKuahmMhXqHpuZfnt2DpOiWUOlauxGpalwch0jRh0PRII6
RqnI/l+IYPjElT8vyRviVe2HWzWz4HBLxRsPv66BAOhqcm7XxMLOOzBKwu0qeMdc
uiosC3Xg9+WFsC5u2x4uhGW7uD0muXA/TJsaxCfkjWC0x26vddJJEyt/60SiyaI4
MfPYizNpb2gVaFcguER6rkpSRSRo9shQ1NbMKTXnzudedEOcsHVoOgpc1SPyaS7+
TR0xM8dETlXJLX8N4eYWrM9fActHlrGLQ7wuc19g6O71pI/QI4u0IqHDOGnbPiLm
iCpj/jQLAngUTPuJtrlawZMFHgeaXn0u5QqVuRZPvJxP7zX5r/iocWg2ChIZNWRZ
3GbxyH8tEZGi7H7ckLnz7KSAfs2Du+iBPZnmX7DNuTpYBJRM7oWrrbfTtSvuKRoJ
OG5381/rQz4v4h0ibw8ZFsTJVt1sLZf++YVztTkKMeGJVacPEQSn3p0WcxzRdYMz
jIoAHvP1pxfKaQ2bspBaEqDnfLASEB2qGsHTlnJ/ZXGbdYY71iHjgp4iIdvooVVO
vmyTX+YgryvXb71jLtiQ2fQYl+S/F7zMECEyLqTrUaoIt7iz7a3s+2j0qgitMqMk
o1AKeJhAqsGOS582TlggC4HUCw8ZUGtUGPMkPb1IDwurU7ZVnGBE/s1ja9OdFb2y
A+f4C5r4PemSA4Wmd/juHUV5wChHGrbie44Out4+sAKV6oFCJHUmuCdRZvxhzSCa
/P+upM+gK7tXGYbVQ+Jy/bs+HvpRoMfyOkBQ1Tj/SZhTPQFTP0K9zETtpcNdi2Xs
KueWg2bX6VisZjQYHvOcd5Pgxk9uz797Ai/mMyApdw0hfkle3EZZCY5ZBd1XxWvU
zBBgvJFhtHtV70s0Pk3fAYNwkdFaDIkMIDZXLSjjMjKvAySfUjHOLJn6fZ7SuMlx
oHg6JP7XnGnw/h+FZsqjK5l/0U/8dROgcVf1iOCcHt2tE33Lbhi5puCiY41FYyEL
91vTjhVWq+QkEvDAxKNznDzwpxAW/CFzPIm0zQRrQXpErbEya2Ql7GRykfififiW
dQZh6yrejHvZtYw3b9udIxYFoPeJ/DK7KBtJbwrxg7YbSGwkHX4KzJpR7rBfpEci
GcCL9twUy8s4iEAkIiN79VIy8pO6qkFwjR+ROH5uP50vdpxdpmZmrzrqku7ciScN
SpUchyNaRiec0gG4cdfO5zCpHmaEEPlJ5H32rOozGXl7l63eVIB2k+MoT9ch9KaP
wQX7pKLt3NdtAA3IsFEvKoa3xUeXqUqZ7vx7lNDq8u/GUmIgPfWrpN7ykWsNxKwh
XWEKVcofKeVluGin1y8BnQyuy+SnVuTetZynU8kUQzNUndk3q2FaCGumJ75EERjr
l/llYEH7U7w0qyMEb52VNFZzmhcPEKt/fI+WXTu4jcako/Dm9EVrJnChQQIROdmC
zre3UwTAHj3DI7U9Kz29YndrL23hCMn9PnPcMWg0rT43GV4IL+qB30JxQ12R4Jh7
pyVO6AhQW8dcGtstfvQnffwMB8SZ/o/cG0NLeNOr0AZd1xBoV0NpxGl4HrnwL3KY
sLhGOYRi4ZJd7Ozi6sVA7oH3Ms2vzuXQL4HZIOZWe4VAaVr1Gc7xKoXKZNGGrRjU
JqqHgAQPp+47QPWf9/ZL07ZuzcQybGSPj8T9jPSASgF22A9KhoZ93bZO0KwZIQRy
xtaC7iIOwi+dQvhZs+cuGuBJjpkRUns1ccB9p9JMS/cgORQvwdBP5LBg59ogkPrc
KGmbytE9jwKhO55Kk1z6F6hrBpqLwaHm2st/ku8Y2rQYTZ6gU3q6v9W1l9YxbhBv
KVPxMc7drCxifc5ospVe3LLaVlw/D6DuHpx6X6G+vzqtOollOC+l8DejdGJWa+pB
QO1jDczsrexikf3IAslKugxilA7xExx6NG5rfYesq6vHgxQvk2djTq8X8gWGxcfd
y7bwTMYym0ZrTIF6bgCZ4ZpgUwG1Snm4pniVMaDxLcnw7xt1VsxGjYeEgxywWhW2
hmDpKOAZ4pjzhyFwrpQvw1fFpl5fnAWPbELj0tDQx927xS75/ZPQb5gWujteWfgc
HIhE1mguISPI6V0VG1BJkWSeG2v7J9fnNXhbpDLSrbBrRyZYAXPugaCqz+PXJQsS
1yUlaxyr+S3p5SIwrvyv57q6f6AIOZc3SVLi/w4YYniBLEHDMHIxTUTpia92sUut
0sWzqhuAKO9aGf3UwyDHLLqHnTrAb9F3wj3daOdYJ/0+trcE+qIL40gyb/BZe5Ua
XmPxDzLqt4GHPi8wHlukOVtoMDnCcw7/nI6j8MXCisAP9ttCqyQWOLKkyZdnj5sH
fdo3b8hyF9TnUMVFtWKrlJE4f/uDi8EilGnWnbA9sS3nd4xrl1+cAGrAzv2rB53y
kiyo2IDz8wCiy4VL0fmqUaJ3YwgoM7IxttJc5H0QsTyFu0pWXGLzVx+Uid8SGFnl
MzEpENdbYSOdZ037+ryeXSnbk/2amEkJMPmzZHaQzDx79OfO0W1Qq47Hg+41diAp
fIE3aW1/zBhAJQY8FGz558quvgXEucu9iETQyz1o60oO7M9Tk5qCLCHgLe22UgST
WLVC6czuERfN1R3D0I8EirGRaSLCUqkeMptg4sc9Wg7x5T8CWd7L5FRpfvDX2UTu
KBhWPezsvPcf+oG48AXYdlrTpEIsmo2JFyI64rig6gELoEFikUGYeZZAB1yuleFr
pf8Hf407Cf8VhgMcV53iyX4poFCHu+CP0IIXB1ZK27Vb+qM8J1Cis2uk8r3Z5QvE
2ymHzpXPSODpwNJeH7A31//RRS5NLP1FjrAyb0RVct36+UcXtn7dyWjKKxlyuYxz
V4KrmHgZ/xXxj06XtZu0OutpEiTVBLiUOAan7zXzSel/n6VwNoRzeQvxmOXZGT6q
YWbvZpT9odH4fNhn7//LWHgizLF8StkiJHgp5+I06SbfqGBDgr6alDGXRMQL8zf4
xfZA2Aty+i1yZhC5cj6fzCHd9+YPFnl0vEhuF5j56hAvICk7owHcBl5OrTOVKOY9
DtKzUqRNXvw6OlogMzIM5jPRVWsFEEg/cE+zYZtx8DW4Wvi/ZQ1UyJM2kmtrKvvT
6JuI/3kjAUFb3e9HXN8HHY93PB423T5kDw2dqDBXm0lQ2VhqMONR7CX3V+N3TNtd
kDeh9Me78zWkwLpARJ4KrwvdV6dcwsjuF/fyjj0NvJXHpVtmLtGbU8LQV1CIUDBR
s9h2Wu2f83g1R/KbHlkWz0yDhRWv6EHz6vy/98G1vL7kAgCLaruJ3Uphn4ZyumoT
igoUCmwz5NJKgFMb63R1tnPu3yyhTYA18LISCdf1NdlBDlDqWm1pypk9pBezr39m
TP3fyN2CdJ7RcaIfRw3mBhRNNNtQCqpSQtrLDfga6HaxRaUQ9pLt0y1/824DvU4A
kiuqD+YGzRhZP8hdqM2FL1MRWEPzd0IZiCV89PJIOcSI9ohA+BexHdhHV7xymZIV
8lNBaFpQQ1q5+rvLA3uzMrTm3BEtkjA09ooG27ora5WSk+jMq981cyr914sfE5Ty
7bVYbMih+LnUA9u3gq/p5iUr1jcXEHCe8LzIwGgdpXjHBL9/Z/21y6JDfjpj/CKD
466GaN9NltfLS0YjQSNd4LEmgFTkvx/Eu0MZutlNtBW7sWHvw7lfd7s+JnCGjeZ8
rhGIldgFh23K39zKbY1Vn1LyH1//N5bYgNkDXB97cfLER3B187rGFPluKBhTVM+l
Hd87Oh9aUCtjndSDJLm43I4eAngNVJ+kS0xOcNPdM8dfICelV1vDuMRRZXVvTXSg
Iqmv9AeWPQcS6ltR/shjOGhkK++8OyqQX+4ZuCRdrYHkTDavNbMhb5iuJF1ycUsO
q4LIPmpAJtIZD5JG/QEfiQg5VSVjpxT0eyR33gpdHgn8+o7ZTbTqxiPeHZAZY8sk
BTwCitKqtdBz+E2uZCxhxP3v4hNtzsYljkhibAZhcUfePx1GiCVnssUOqlsFMQug
YMB2csESnTPRwl/QdzpqTl7sOvM9gMxHkfRrQP0xoE8G7lHZtQPthWpede9Pq0sj
+Tu724fvVZjJpcG4txl/QaoTDQ2TFk0DDl4TZHeLq1KjFeppCKNLZDabW92+Qkfm
jMMyiDP1psTE+uigfxFt43g94ivLUf7Birlv/KyIvQbHXfwPOW/QUQw6LG0sYb5q
xku3CEJQNs2xtAmc0FlN8m44wRwuX4K7+hIuzNRUDtKTSMPg9emPCedYPbK8bwj1
N6vAdmvWZvavyivxO++H3VFSzweDDv8s6EIDABKVqRKoDdZkhQLnwngiDPe4qtYM
cpICxOB1wEdHk6t4J6P/NCPX/IWVLmccN7iq1WiJ1sgIjpTW4Vs8Wm6g5NEiyK8Q
YB85GUxGjHEwHdXzVA9uCo8ot0UbnYFJNI78QjVEFqkYDM7kiBBBvXJtdzJS1uO2
hBdv5p7kmAHBNLIHRJX+6c+Son3ggd70pbjY/CkUnWpbS+D4rTLXMCqEoufCsUXA
92e/bzo9HBXoD1uKr3YYzVMnGpdlPBvBEtFJRudXk07dNa9eWcdRxzkhPpqyK27v
FI5BiwBMn4D/96PNMovkZ3Pu2+OuzZXUOcHy0u0SaF9u7MjafczlkL87BOMAhMai
IhcNJ+oVXnU9qhcFj6oga0zWYlCg7wqnBIrkk0KA0eLMGY79rZVoDCEp8BeouKNY
Wr230Qk+w2aZmni3M0lJxR+I6aI8felcVUPQC8gwW2fJcpx7gOe/DGP484waCIQV
w1H2yxsslAmq6DxyCmw+mdPmfBBxPFO4Ih/RyF1HCnzRRwAk1pXPEg0C81W1Bj8+
GvqMuMqi+Lc2GJJb63KejWsY2wzMhdskQdPV6x9fcQtr4hVezXIruc8Gmqjbq6Nr
/AWfmYbbFHSlaMy1sYFkrr6FgNICXpjF/yAICCUi+qpk2zu0VnVfkwOAK3Bl8uzF
uASAzZbnaR8t/f4JIiuL/TaneS833t2h2hVknnJ46Jr31inToGhzWtbNoh6QCy3e
JalGSc+eqRwZx9fEGdOETgVJvUuwMjrXIn1ETfIUcRVfXrOqzCfhWfpjtYgfB0GM
xDrPhuZT+8TTvxl3ONzEG3SWAVywIB0QhbJotwlrvRaW3xaR91Zp+WiJ3ngpUJvj
9jtf/QCzey0RGcPTR5Dk0kgPpppH/1pzl7gC1FuG9GPfmcFaCCD/ajq5DedmiyS3
Aorbx7qDOFyhXcbhkYypcGSm1fAGCMbJvgpFTRRRudrmXZrP2a+4Its9Tp0FRP2V
xaLh9RempKjp27OoQJjHk1gBGTzIjbz80W5A4mlNdbZz9rd7s21p+TrzIVIowcmC
QuCgICvVakDJkX5cwzb7qBYC1HmVR1qrZK9T25NFJaaG9SazssWN0JyY5G4Bmm3+
urR9Os8I4vjoRvQFf9CwmjJi6aVOW8ACmWmsgBbjhXqJN52yPCcFltAFxCiHrDmp
XsTXXZMgTAqiL/HIOSXqLm4oOz2CcmOVhKbt7yQyW0Yt0x0mJwQ+Y3hL5SCeO8Hn
h0vktMb1o/TAGky1THCr0QjEpShA5/2qAKlZSPJNW5JV5a+eSKIvLYWdMZk/Fume
NxVUHSUFPh9xRLsDdBgi4/P1sm1D5/LhQBki0+j2fx4jwLUPQlVKw0eBJMVAYlGH
AUX15FKC9YRUzUn8X2kPHANMvABIXyE4PHludPcNFqPR4OHkDDThetQSLIshC0y/
wflugz7LWSXNVA2cikbSO1vuvnKVboPuaUVdMdrWSbmP3vAbpxVcxzcAEB4txzfN
+K9FpbTKcyedIQ3jdyfiUHA0lZoGnJug8AKsi0b9bcgeLCJINytBSJy0P3xV9sUc
RRPm7JcZ/4dx14LnfcH0VXbkdzhFAlliB1kDuSLNLfXgVq+tI8pNyxJtgJiUjn4+
7OEEfEuMQS1i2hBnKY7rIoT+1dtq/tFItvvJIYLsiB93Bj6qfaMLhtKaghvKlwu/
H9SduTkCRBGHdPhU0CD4CakeypVA8R5/BQmDUd80aTcLjI3BAU2ggUFSWRtiFZGo
2VnwqUqUejetkXSawfLO4UnSlqwgkls91xribRH2ZZm468Jv1N72TIsMjgjixXBX
ABD7ZXsQtd25tbr3yAjRS8prHCWd2cNr3Wr+927CyK/qDYVtECpTJR52VUweQrjF
WHP/hFBen4AJA8UuTJM+GCIXIL2u5dAnyOxDHEES1NwuNn1DHRGML2IFt12FiRnC
3jcZuVoC6pQ66MYCDLRuSXp9gHmpfKchVgTF1DBB9sW7zmslFdOsCWboiyn1fQ/i
nWRIRSSSYLKQfrZA7VbrDQKZl6yCVY99p2cIHSBFC81D/Lgf8DH2y0R6EpKWjwGI
I2ZxMoCVSH0zyKYIqehLAE+A1jYPd2LMfEmQ7kvOaWqOrSoFMlsTkRnkPFqKTMyg
Y2Zbjq5N0XYNMhWwZWzgZooO7+aSaSedzq7gNNJsPf5WdN8RG7Kd6qEq9b3obVbE
139SRcGauHFtcx2RiMLtJjuSz5L2cvOH/sKNMXX9G2Ac8/YdakzzGcAs03aWcV+C
4pEZ0/zS6xEbRb1mUtkZUkKt/fxOBbjKaAENFOzmXnZubsCMMdaHfxdr1LjRJptX
xUcU9oisIXcI2zoi1O7pr8R8m7nKSeNSXRI5r/t1OehVLdVjQjgIy8tdB02tPDXJ
U1rR/QYLZn+WH398mphhSqSZzxTBoL+yb93UOaojKHnJheyIMnG3bSA2F8jPE7St
l+IKhwQkm05ZPaoxYIjg0S16iJbTYSkwQbhgBwl2OpskKMGMUrItSCuE5fiLExeB
MjN6su5l3sNU0WTWt8vIVIcPiJsglNyaFgFgRHOgH3HO5ue1cIffh3ALQITyiG80
Hsx7pl54687tZjMLI0PqtgNyE7YoVhmnE/oLL05aBMClCcqPDnASRR6QylIYE8Fh
PGitZzDnG80iPuoW0t1O5Wjh87lDtq17y2bb683kH1GeXwCwhJlRsz2Te95d3mxF
fo1y8riSiRbA41IPssgNrlA9/jcpaLFvarzd8sPrjopyW7Gz7Wp16FFP9k7Satxz
zjcvHzcgFDwv4SCx1ElyR8Dyow8vZ7/WR6SfD9GNFvFaoyGRWxUzY1NXuc5ipomw
hceF31PCUMBWniMZV/Y9aEaiiIbDOyqxnHYEUu6qDnSH4uFZwxU+n1AK5+zVNhLK
K/ahpkeFiNqU0CB5rlTXkSv+B6633H75/tkJFtwQ2x3J6Z7l6TaSbj/x16OCJ2rR
ziDRLao0MgSCNNpMRKggq/aKHUJVMLgSen8/UJcFDC06jf/FHmTPJX1FYnVaDQ3F
Q90Vk3eIWKMZarrvjqlUCuT2HJdvI+6hp7Xsr0dwTR5/CqlZ6JBULaidTmDTdxt8
ASeQLvwGpt+8dvbcwaoM/d0MkI8YuN8HI/9AzsAq4GUU580UFnS8ubv5hSz7elxw
BqXMwQ+CS+feooQ/M+Qnr+RbL+p7uUbo2Hsm9pp0U9bCj0yy2zVjYwbv9IYh3dMn
oDUP63H1a+2QHaX46AX2gygstxvpfrN1YTWu4+IjBaSogTkNoFHx+qE+TwcK9918
6tsQGK+X6OnDU3q8Lf8VAcdKv+dap6L/WN/8B7Nxu7odfEAY31C1N8Vzf7xmOgUf
8tnE/dB1hV+sUUGg305UpXjqlUWeS/wRuU/qrGd94D+ObIhixMYkvd/zkflINRFq
kr5rBn7+2oACoUcz651T0/0wkWcEZfBtZ1plWaE65ckg622NuCvAEGNPMfPlrE4l
4c6FkDmm3y83RRLo6xNFZoydcqF4AXUf+kDgk5vFGYjaKrK2LiCBoCorXthUn8eb
ywP+LlyzG4fGrAu/YhAVIjsUdNx0pykOBvxGVseoB2TyX3umDVUo4LFOr7bzN8Ml
xZ322CMERU/SqUgU/nTuehM0GeCHbtdtal9LAc8VbDW7IoY1Rd5mtIIjDBGxLdTz
+8ROiousnIIHgl3nd8es8lnMn7+5VU7w+YjpFkvPa9L8gyGIovl6veHG91ki99jN
qpmKLU/D4wLfSlZUXB5AZWdo6m2asuo5XD9rl4x0awfm+rEYSeK7FF8GWvIklxfD
S0ciBKs/NIChdnBNuIlupvEAlTFUH66vFVY3ud+Ut2LILGTWJlgzDAb8HcRnfmcf
/wLEKfZJ5oZ15oK76lEgOHxfSaJj+7eeFBcfj4RpiSnU4nznQME4zwq7oCBCQK/F
t872TLZoiTahDHqWX4ol1wyL5W2975SIkYZ3dG0HlhNjQakAj+Sf1JLwWA+7mrWc
KCzBvLdA2EwokV1A0rlEBxtKhiVeAEPYfeMfFoJ5CkopvBSlsoXQmg+EZn20XkoG
+aaiwnFdAfj+/FEIrpFXSvpoiGtUm/F5LynwMFh7kkoUmxoF5BSXTxXN8YXInXfT
f1LsTcuakapeG2hfjk4uxRy8hTgd4lQf1U7lHz2X+yw90zrp6+2gK1KVNhvL2b1x
olaap58p1YAqqwxLJNwHJQ5Ztp1tgnROA747ZnfqT04WMsvV+jy5zWr/AWvg03BB
lEPJcghJ3Lq/c0WuAz+VHs319/dXUFG/bVvH7d/nUw1H5YJ9EywckgDO7fe2/hMl
9hTeFxEN3xb9Rc6iBL5FShB9eoTU15hRH106WiAei4yTfNWKGMrN4p2nvDeTXnrw
CXDHbAlqRQeJose7+CZsAu+qU0bHqyUHvDbCxibfPC+S/g5MDILVPmuIfYLVo4rt
6ZZuFfG7T0Duqeh6JPBkp0SJQdw/VcBjZkWw+qkIYLEhX9jMg15WsxKT805g+gbW
w4rr+cJIYcA6LCDHKwpLJWGTjJ/mtBY1vIUbmIThSyXQBzSFMFkmj8bBfD4iBwch
Q0KToXH4ILGlYhPMyt+/4m3MpNNRBmSfGqNb5S57DvY0+kcGGv+crdsux26S0ng2
isdZyCZEKtJPbEMLvK08wkjmATSlD27xr7n6Nf35BXPMJ284YSmJMv64jt4cik5T
X5xf+cMJ2Wjxfs8mT3K2LwBKGEMhIVxy01lcG8nZPfe3ZNK7oWNHrVXBfZrtXTCg
j/ml82W/hQc4BiIeVvIDl8abc7rBZwIExVrMqExYqIhEjA8Stm7j9T6CnEc8QU4b
2Ifug2YZIfJF0Tn/c1Ma25Yi6p4w0Hdz2ByznZOki8X8E9kjgOQ13geiPKVfM1s4
Mn1XuVzOGA/ruJFQL901ZfYeHeKQHLDD3igWWrsU+l463jOjHZmfyZWNeTkVsYw6
P7rsF3OyIVa1kFZ5ER/IiCzrQGKKq3RLqQ0T4xcGLeW+MromHlMDz2p1jw0nDKmz
8YldpUCtylsK76RFMaWSXbmvcIgdV0q0D10pfdFDNiAvhV2l8HmOHVWolkTKZoTD
eVs6+bGP5i+J8aIg0se7qIay488GyTeARs0DxC5TFZOeP4BXMCIq1a4VXSzQGEDf
H53eKPDPUvpkcxwx3LCgs5xuGSP4loXaypGbt4l3AmXeBXuO42QbtqCgwcmkrKHG
WhVODhzyIS6OlEVFC70bXV0tSsKpz4UENxbnP/auy59SnuEWXDC86ynmy+vlI+wk
rF+PXQXEhtiVnf8IMvDtuF03ESV2mgW4y2ABaxtruTDGlT27rukPGgFSNigvFYmH
v1RyqL9cA5F3Oq94W5V2CDktwldKvzPDFmGRa0sOugAicHgNhLCG2l7Wam/bpc/5
XyYYorx5NBDgSqN0Ug8s0ylNSsTRLt+wHYiaRBEEKKhp85cMTmEaBzsbr7OB1L0H
h2LNq/GXloC6PebM5M0adGBKn1SF+YS3HygJvlDm+cIDe69PpXfE+djh42W7BkOW
14t9Hi6n8/ynep372bL7jSJmdDIksLBUxZNHSkJfd4+ZLz07NTZqms3BPcZ2pDx9
vnDCxVhmOqkV1WV5v8grrhR8ATPLh0Km7BeGqz9Sux2QF5dfsHVuk/yWWd1MzrqZ
9KsoS5k0ZNwbmaSEQZDXIhJTO80tY05f+dStN8JXnoahGE82EZqprsOt/0ltzV/b
DFSaAKL8JaZxjHEBPe9frMZjmQRRHnGSlNoM117Hu+IR9WD8IFsQu786WMzhIBA2
t4kdfT4JIZC6/dB2k+y3yp8k7lsErR0YYblRdquHf3EE231jx9H3jczDJXE7sJ/M
k08aNZWAYQhK1J0oYqbo38/vPhf+ERJjwA99+cByfdIe4+Ia2VSVxJw5No0+sScM
sEYSoPjMMMudDzUPxmSyGQ4ZKYvDmcqv7j/XI8kIUgOSt0944NuQmEJkPJpuRN3w
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 27696 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/T97rZhQva68T7JOm4bkq25
b4BW57ADAHEm2yg/Vzsfl/MRd7M4YTcFnCytkyp3YRP8pg2Y22PrREMRYQ2vNcur
RtN23Z/ZKPFZVnt27HioHiBId9VrzwurPr1c7+gRNmOkH405+oEhjmhK6OhZT03l
TuVyLVdYv//fy5bruj9Em7xEnjZPOCh6WtPFOaVRjmjHKzwvTqz8+ruSOpAlkqQ4
6YIhs4smvqDqZZEdvrVJ/3l8zkgKd115H9Hx7JZLYj9/UuHzWax4tnGbNYCaVmur
WF2jtyVsUPFyb8ieV+Xjv6UAus8Db+QzUEuwIRU+Mtfrtdd2sIAN2Lw54Z2QHmAV
z7ZfSWUbxyrXHBWl0CUBAuLRs7OGs/h0Eic2n1u+aMdJdaB2pO52SQ7n6F3yzCdj
qxVEk9YvcjJbvHWnQE+i/B7X96wDeNK5FzyLMp23YseO7J/cZVbLQzlx1gTHsKhR
ztEF8acT5dhi3bgwHUUzoqs2K1CHlTOueOQoX6XGu4uFGY90rXx/Djja2nILL4hG
9AJ/1XtsyaY4sUtPZWNbeHv+TGjRHwPcUU3tARwlXSJRp9ZGw0f7Ja5Ldb0RpXjZ
G961zivSY96HUiGhtJjDaMNp1TRYL4+i6B+4jjgFP6Qs4Y1VqCAzjjfSjoZ1Lhyf
/buViISb5TNLdCQTsRrrulPQEMBJZGWzmSy69K42fquE1cCzzSQ4W4StfLJElGw3
LeuF5idZQOs2jVyTX/ldzS3bTzSls4xR5z7EjSxDHqHgM6+0nRthpQ2hSbbAkqUq
RPhg+n7iK3VXTZG4B1uBYRk5GS4OoHJ+V2bD9dV50NUaJcDAAylI/ZqhN4AeCRS9
JCXZe+1iq9ZWwGKowui3PWpIRn06Ch2F9fxfUyiG8iQgPo26LHhSz8iuwQ/QnxfE
sX9BBWWyS5+piAbf58rrIg8EeXTe/eJj5wDMA96PqvzTfsd0I4JHKhjNejbo4vbU
sWBPpcdidnH2W2YR5BKkYpGJT0YHWw9ErW5YFnG6kHtJ/aSgGzjSbaLQMPwJITlX
alcz58P/O9jMSiNEXAc42J/Lca7OYVJp1SoR5cPXaS9hM9QIDJrLz3y2P1nfLBn1
uhm0OuO56Yf1Oi0k5HbboOOv6OUilLenE66uA0y5T3/YUEJAnJ/EUGJOnSJeSoUw
bGsNY/QJnVS1Xf8j1hWyofBZqJM+0dPApLpVfS/ejS4M2E+1pq8g7fUzXxhspaze
jCgfWpVIQGOpIrpHvWXXb3xLggDD7VK9H/ZZZfPdNa15aVANhTJExYNKO47XVbKT
M2/aOXY7u+8FnsQDl78znFGjSu7mVoVg6xSyw4qKbNdDQ1FWWoIncrXz7csT6z/q
z9DydFB1Z39Iio8A6VY5dPVe0U+02z7a4Kkkhs7uHs3tI6wUDDi8WJXOASbfxTPi
LcvWVp22Wnxi3dOXiTLKLUtJLUQm1RnAAbl60ZXbyxK+iamrpwfFRhGJi6mSZIek
V++OJvpnecwriUxt35mwBN0lmW1S7qSW5MJF7YKH232n2kCljUqdIq8Lw7/S6JX3
+SQwQQLoUaWodSK+gLe4vHPoVDalVeyX4aN53JeKxRkjlJWvF+SQkUH9+PDtrlJE
znwy8cqZXq3JYp+qb6GVj3hPE4MIfVXZQyZ4J6VjDLItmOeWzrPv3rv8DiJpczbM
DNcTaxC3Ua9tsRn1Jcbjq1U1uJMt3OtzHcSvp7VeLNU/t7pGiZ1GJ+PKeZbMpw1J
ZR5kBm4UKFt5yT7XbcRiW6PV3IMFxxlVuoXunb/PVXWOK+vq4B/x2XaKwH9ww5Tw
k/zScrCznpRlMnu8/74OZ/pgY+lxaV0Dz434Ejhm7sl7cBrCi2ebx1OXQBjF2wIt
irKr1KwJI0GP7l6ijXwFXVDMXu1SGi6Q8hZHM7Xjy2js8t9b0Lbs7DKK67+V/wgs
kmXC7xiN3XuDN2wy8Z2N6GEAdNtIIlX7FvWEWjZXscU/Jl98hAYwy6kQdQSDKP3N
PCDOKCJLk0D+XXGPG75+nIzRRr9LqbdFR62/asQ9wtuyNj2B6s/k3poScgesjqQr
rF/EovF9BOr6jLbxlUYRN5X6r6KMfdUTH9b3I2p0+m4pVOAljCtwfb1xMxbO8c7f
ACZi/bu+iumKvJbdwTAiSf0DaqBOQHqt9O8YoPD/IA2puXRXDabfRBnedZ4qGp2O
DLJSWGjunRuxGPt+qcdtRNpEgmaKOxXGdh5stJzfkGCtrHT6sQ/dN4htc50CoKyT
7YzP3xG/yCoNvz6Uw6BTm3z/7zcsMgcROe2cmrzkCy7wFs1ORO2WE5v83B5Yn6Pd
0kZyR6VaabL6KUqqhZXTk/1vNL3g9OSJcOW8OEikUXC5C5uWC/nZ7Ad4kVZ5on6w
EbiJ6UjvPbCtvu6V0SJCV85pGxS5GEbjv5kC/KLbFhIbG3V/TbnTtPppjILTFpxQ
yNA5wGQe3YGfILYoR+nQuRdBoV2NUsQUjE/8MSOGMO6RYgX9FMCbeDWXcXDarZ00
yk5G8nF3qomNHX5uIRY94EcQljlBY6MJ7VRBkhYCgl9Aroypmx0zV6SLbYvtoAWi
MO2uirJCiSKVN9GiJEzDXilh5YKj6fCHgzgWpjNeE69rlBjrX/6ZJZPcNyCmq2me
Nq9sPHRbuPfX4dyhs7WxmdSVBYOvAd4vDJo99we9RmsHNwsbPscCSt1FKnjSmOAm
1p+fatBEKrEdOOD8AO8dDLqdnIAA9li+JJtTz0R7VuEGZQcOpjhm0JceP8p52r+i
c3SLkYo6k4lZ5kFsHywFQAOT+gleM8a1Ri0cmrMLMKWNuJPCks8IDR9uBioNBhOQ
4DS4KDY1WFvpvj85i6xtYXd9rX45JLpIfsCTFFDt2w1NI9OIbtGaqG+v4JQZ6Xvd
pfSEdzoLQQjIpkdYIpCvd1fWb/ZUTctLJjyKXxiGtmnk1b8BbT4Vs3igat97SLv3
UR5IuSWZWVNlw4xtkMiMc5seU1RHtmfzH93z1qCZTcuOjkX7MbqOe9mXRy9kSXl+
SuDy+WSJq587PvlFs0gn3dpGd+8FYOVl2ukx1wIyq13ePQ7vIC6Lr4XjODtEEOPR
zAcEs7NYI1y2DnfXPdGzBMWUXhKJUVmdyYmd3tQ/nEf//8tb+BiSL9CaHMcpvHBC
l5YLKv5PmsNwrLa2yAZgdzAULkOQtJ90qvww3Glp1m+S25WqMqtpHUgShikI1Tdi
mYao0WAUKnRIqUlVvc3pYIXoW0O3GNfsi82VzhMxTc8bxYigH8bI73dkBUAEtbaO
UN8E3Kgtm0emcmGqZLWMfVWrKgWg6jSXNu8RdZbfAs57NGesd7ijush2+080IBPi
4+zyHowdRNwLG3Jg37zrC6gntfX1EN0et3GYBVfUikUeafOB9pIPsKKzukyXOoC4
c14jmXbLhMsSQVM+KfL46/HGdgBdIFt4cw+V6+jVjyGW/OY0MhsyMfkrgf2/UpOW
E1yxtPbrLNrZIQBJYh3eEGgtQL6zseKmnc8mmbAGkxsOMejtCIInScB1bkjtlAa1
BBSN8N/3XZGQsm0ar2zycttcQpBEww9rL2XpIqQS/o54wg3ZG/UXnhBd4vQKnZh1
FTYrmWm1zIjHuki/NSWGtKtwmOTZf9bL9ITi/QMe6lkALZjgOTOgafj1SEaiOvgB
n5NsbDTbq3u4fbrmda5o1Mt0K+1jUu+2uEU8l4qiq8ZcxAFpc0R6nAAvAQF52wNM
xQB1ZSFQZz8CScGfWksne4uegf5ZvT9+gPbx4JNR8btNzjbrwLOM0CU/UJAeyS2k
Y2TRTSl3irxp2qfE3c4J9cFCKuHeqRdavUZjKO71p3+nU2ekWZsW35QlkBwdNMkA
YqGe9uAS9UMoriOxhaZN/mmUBzAZ4Vcg+27RAXaQsjILHMVeAUXMMvfVPVtSqpAG
nxHurUdBpuV5SPwPoQmo0GBPGehD494wJiWLC8e4PpIxWfenbSHnoJWnHlegWezy
PeIIHB+WI/eBWLQAa8daNkkecrn/FdE5IC4eZWQV6OXS6TErpyLF6stf0OEvPAwG
ntGCUY9uv56dwtI20kAsu7s0hnvPOJ8zXd7zL459g8+TMf0PPD0vfPJV98GOyKrc
zepUNid4PQQ8nGCWPeuTVWkHmHCf2ahXVtKn4T2+ElqnpaESgBfUhhCfqP/bjtPT
/U3ebkpk0KDaYJBSwDpONRk0T6oOyPTfqpMXThZsLFZfqgzaCATFJOHfVbWQowl1
Yd2UNAgadfIm9tJwV3UTCgoW0YZeB3h0BDsUFn5SlfakSfDylFzHsDMfaqciN8QU
cxfVJsQ9CcSLPG+V3hNHG1aCVphocyWtPi16LKGWBupVCV/VW8otXN5pjpDg5CKr
OcbQhYvp3dQayjqeRPgE5xDEj/RhbdvDjJp8chpV+1SHMg4VVnS9J3K/M+doXav8
w/l83c4dz3+WSwxTZjU0x+CVLt1Nkc9Fp239rQ119AfugFu/eZHZueaqHLYNuj2G
kmUoVGZLaIvCuYqFp9jaOOPoL5bDNVILezcgZ81KBuA7yxj467Iei6YFGukBxsi7
QeBzWATDeecCZ/q/OJlALioMvBf73+FJ44tmqKDvOBvZj5qHsLxF9cjlYKiSmerE
m3YhBNsy04tpZSe6XKBuCBZe2dTBIiklCHWryf1xdaIIf/OtTL25cUtRH7V/E1BN
GwPJ2PRbxhlMtyZydb/eNRPI6zPxa2dsJR0P6zHVsfXv/d9vKj1zGv6vb5cVbl5Z
qxN15QPdzGSknJgv0RmmJHJtMhZZlO7u0zqbEhJknZvQ8B8vmqNVuDyMdhfSPMfS
IKqQbJVJebqp+f7Oz/OnA+8N6fyy3QZJj1jyb3pdhB2pnrP7QRb3iePZhLeVvPMj
cv7wYqTIWiF80UZgZuWnA+vHAJDOm/qRIfQ7EVL5QiAIkB9vMeRHB8K1KVXpwPSn
NR3E8eeUX/kpGCp29jKD178uVbeBmq+jtv5dcOcMHkvCk2gEJ3Pp0R3bKfmYC0fm
ojBoFoo4p/aBbOtJcPWkY6sQpEiCvcpUJ6PtuTDf0DZia/POHFzlyUlCGZohXbXO
rv7X1dS9FYkx50zUxU3Bu0QCyJytPXlChJRvtttaKr5dnOosN+umEKuJXpaEgoGj
JS4N90kqLYcRUtkefCP0TM9Z8toQH6MYhXXtweJdW3S4XZS9zZsSMU5OMO6Zcrr+
O1ClwsnHRE80Opic7WfxIqasAL6ZcR7Yjkg7dMnkY2pxIvlaQfcL0+QbrdRHveiU
KOE2g5L8UX1iE58J9ov+ZYXhUJPqzO5Z2oO5Sm+maPU6aTKxj3UBnl969ppIfMu9
jbgJ2hvw16ebuQoWTgwCEMI2kSdN//TfP9q3J+rQ6FpG09t/L0J5IWXPmH2DCBcV
0jIWK9qzdtdJeaZhNqa5zvM/1iwY2XleaMej8cURuMIn6OZKiJGCt3ktZ1vrdV0T
S7b3g8Fjkey+58IhuvQsquF4xDm2vCVxiwPA2OUenpHxa5kcdEWPHXeOp1k/T2ny
UINFQaAXtWyDuphfZqm5MvnuWhR1XMmkN9IVhwJts6+NYyBnxJd69i0zCE+fs0b8
LGUxELlW6/Wk2aiycjhV8Idgif2MTbbN1ZvloY0nW6i2wnJgXOe1U079IrEpjoTt
9vbRxvdPNpD/03i3f40i+yFlvFNUqHv1asGmKNlm0ZUOjL55qjdbYjKmqs/i6gyr
qVGUHSgoGAuLHAAChwlGeZYD9o2I93vq6jqBD2WEnyfPdQGvt4XXbyrYQBL/hx5e
tW3o2HppU6qfYgVlJB6tua27eO2jcyGOqPkIwHROnNZWeOMxXLtrNBidrZ6KOc/P
pJhQ2OJRsxPMkj87Bn0phqCfkVC3vBXUIIhYWkf7gV9nez+ZLrYUgPBvDtbvMegp
AIQ8CKanW69BPySIgilkgUWUqpj88IjtUCmTupTpo5PFTE/ULA4oZwx4QGY9yE2A
jRnpu/o7o0TOptGzqylnRwg55Ks7XiRk6QDyCkWavWyM7rKFif+qT+I7CnUVniZy
D5QcMXAVkwQT/Bmvv7XYLAYD8WcDP+49IMCVqyfYAj/vhh1lE1s0Jx1afrWzM/ee
QerWpX9iA6DllRLrd8L4jRIhzyOfjUbFvZa188dSHodFyuptS54FPTxGdJ22koMu
zWwCsigb5bOLNo++IUsdXGZeiE4w7vxObaRRIgQwTiJxFlPlycIM3vU4FW1Vvma1
BLc6fR7NHnj37Xxf1kNQ9MuyWsD/8HfyjENefUtJmqyhrgvrkfkjgbv7BbNXZ9FM
bB9kQxv5HWcOSPfoyBcjhSjUvyoIkE0+FJG0jboGNzxsNHZfWLAAjpLTKnWFAEuQ
V2AmsAKU00ZpZwwv2n1Gwpw04oRrBwyIacLn2Zs7AdXv9z1J8mWYeZJxw5/4NbF3
d1MMHNG0yQRZm2NyfNqcKw2uoEXt7JOvoYzrlU9+/5wPt0lIJMtvt4bBADbHyGbB
Jniu41UZBSzyv/SKlb4Mu6DjriegaZham+zDOhpFfmyky8GXNLO2hSSCH1nXG5aq
+x+42FzLhC24aWrUlrNOTr2luS4is1yQR6IMkNXFhH/JZfMOIxb/SQ9xCtCcrXFG
swjizMWoQwPbd1RXib9beQRfrgT/Beo5ehGWNL2uOI8RWfvrRFTyl6C4cttTV0Mu
sgZcbaqtapnoHq+54RVnkcgCEdiIXJVFBBpi+ERUwR2nQWVs0gluBPdJTEl7bnqt
t4w78d615zfLY34AFAMRgTJl2QTToB3U+9TAa4jhRCWaytXhH2kK5ifRDSveMARL
hMNRECv9gce5bEax3Apw5tBmH1E3U7r0+NKCWQv4eaTqEW7fQCZ4juTvesfUPqUu
cH9VvTUJiNTw29jeulMguIPL0OjyCQOmqehMHPS3JMvW60aCmgNOjptuCanPSvyU
gQful46Bs/HaTN5Xldjx9ekXKKmhBMaRSbF32lDKFTuslaGgYLfwG8yOmtMw+leB
nCAWEkUgJ7wLo2QgSRnjGXcBAB//cbrNI5WmNC8NtTCww829nU39u0feZx2L2t9i
wooDE7uWivHJFLcOEvTdKP5qg2Sx5RJYWmf+//Kf7CgfURQO7pbtj81TsmGsUfrt
AjFlz3S7x2RU7vsj9weReMZLRJn1+iWd9gHyC1WOMTjGRN04nuzaaQIcX3AgAhpS
jiKSZjZinGrHzxTPNskPquJddIiqg238RXghFrIzJXDcn1DgLMneiQBeHcVZSfMg
/CBwHK+Ve3tN0NdS2xydYTChitvNLpy1PqiyXh2v493Rv2KJ7KOQ+T+n1HmzrdR2
yYhCZ9+hvEP0lJGTe9p7PvVaROWftPVMx7R+ciF+RQTvl/FqctXvZdsw2tAiN3cz
vzmQ/5odIZ+c56fqAGxguMnrK0HubpzdM99aLPX9qwggjuTNRmaE/PrOioWAUtUM
qv7phYC1eAWW8FwH0mG/Tfr3u4IG+7CgX04mSnqQHK5rn47SJQ7Gz/J1MnzZ/PKO
OcxIqQbm/qm9kujlO1JHlVPlW+v64qPrATzItDZBYirFwjmcbY2vGuzuZZrL4/ku
OlJmbxzl0Nd0p6f5m3frqpDrVEDzF0xrPJQ5WaAzgn98UG5vqxdnA6Sz1AORqeAn
fl26Hjv4piGF5Ih4P6chEKXq1s5vL07dRa8VvTV7uPd8ow1PGTcxLH/mm6lMo/L8
sUkoEKrYfkpsykqNddoFiPGRzDopHAU8rZApbnIhkdTruZB7+Ro/tuJH/Ex1qTLX
yLo6UlhZbvEb7yzBV5Ioh3aXapHUAz/ft4bUeTnGPSO0ylQOPiiz5DyakWgKIpGL
GzoMX700enyFmPtqyFLRapcM1b3bRld9DJLzVa9lkDLBJxwNyrgWkM7RPfXkVn3E
c1AFam8FjtFBn+6P9hbaUzAGCaxLAjmKbKAor2XWFuh+KBuB0OFZkktymsQT4imX
mbOncljvcxPlgahqER7A+78rUP2bda13QY+r2iWGIlkMLx9B0rmKI8FC2HbngdIv
St2PQ+hKP4gimrKImGA0a6WA3aYA6gwH+pnRoQw7kDER2KfRTt7XEnnPlGkUU3DA
BtF8VWwD+NQSXexPdNpwg2NDzNm0uX4/PKhq/PDYcF++gbbgF6hgKnVh9oVp9YMm
oj3H3Yfr1TDhTfaR92IYejcuuDT64HqPG/GHAr/s+Vtu9f4vr8+6zD1KPiSWhNYP
H3IqJQeZmdSHxZniyh1Z+FiBXVyexuB/hg5XMEylmxHj7TdDpIzL6oIGqokIaaPM
5GVQtgu6lzZIk0lGPZmsF1OSgbwHnWORWU2M2ZW0DmOm/2VN34PcmLDO+tj6hbVj
Oao9ncYV41NR0xL6PCbHG4jUS+pD/4cPYDs7lZ+W0QIMMX22Sm+iUBo5yoMDGao+
abqh8d2JjnIAIkkTVSSTAsH5+/pvYD9B24FHN2fDFsNyH3/i+RBqgRmggII3AOPW
3Bwp8hQkX44pQJtpBfk8XdU12YA47qyp1jNQy/zVlTpg361JO5Al681T1PteBvNn
A517fN/Ei0S2ZHLHidTZnEQfHQj4QPoR4Dn848IpT6kJF41B5huD4LpkXVbfVQyZ
WN4HbLvLa03UkrCq4YVwKLCBJpsnd28MyUltrdYrpOxbpQsWs9FcSRdzpYTKRsfq
RSM1y+I9ZDbvhlH8f2RJXYaaUZS6ZtJxIhVa/MfLnAbXHzU2xJZZHJqCpSokBsvF
iZqOz3WWX4N/P1tQlAFiAtWrvqpMufOXPFwyYEBU49MEO6gJL7ZHpnYhfTSd0F1P
oxRcZM6M4aOjsuOEMvL672/btshmCqk7SyCU9l/RJT7e23z/2iiiXPf89hQPl+Wx
Vs8b1AQIphIKRJ3AGPFD6Xg8HNOsIn81lJNMz6Q4qynwfmWMasYwus1Cmno6LB8c
EW32lLK2P0w3S/WgotA7tsW2ZYqVS3NqTyIch4Gk8XnhQShS3KGtOmnGZ/On5x9C
5ggyzNjSYAT0zsx3Sb2otxO5e7uSZ/kiQBeSEe59qxLlmioQbmNH7pmtHluRwHpR
iteyvWNJjcJLLdWTGyoweG75FB57kUc/9I8eJx6DVDS8OlJmPbSCgB23NtwAzKtz
J5yr0En1l3ET1UFq56sTV7j8GOced6oM9MBvumUwr37t1F01PMwIGFJ3b+YzxqM0
QE63d5IxKOtz9fqQ4tbtZYdIVN+T5P8JNVd1ssOu0hokWyRqIv9455OIM9Cw2fZm
jwgQWvPCIhOcYcTXUB8nelaZDiIRbKpzP8T7X3LgSKyOli/E7EhT886ztMakM90v
cyMPVwwkHDuhGz0wQ5Xmt5aWQAl3q5WyMEgmdOd4GrjvFDiWyEiYElkvmSgnXu0s
ihazEO6JJVqmHnLYzgvz6Ch50lOKGK3bbYCqnNO7BFpnL7f3S3C7cOsdXbCujxK5
fVFFKosI9CX7GLbj1egUQI9J0qgnf0pjIygd9lrXb+bZKdaPAQ3l93OwcjUEoSvM
8emk6j4eWAg4+crFVEPSVTBzFxKeGHDk6P+dqwTAxReEDbdzlRHoBivMkE8Iwl6q
cITMNgd5C6P0CACt+YdICj0YGkKWYGECpGZm0vhfVU3CmsaHFJJHANu6vle+coMQ
nA8gk1YYPm/K5vh5GPEL7uVt0cZ3U0TOzMkv1GtQLpHnUHLQYu7aYbOyYLAkF/20
aUNku3niOczV+z7bXBcS26xdrIXzfnxhGer4uP9z5H6sm7GW2sVfwrl1z/g1+QFC
sBTDEvimnS1dKAMF8GTHj0gbGcTsaZatnopKuExr7WtsQnBjzzS9Zqm+JUGQ3UYH
zfCKekJcr+ohuMsRwBxWKixzbYjCp5KY7nlT6s/r1bSGmEHRqi14trfOkb/IuIFD
ndo7mnrJfHBmOhCYlSwwY9eF29mgcOQhYy/VYMbwsZEZnpuM47OoA7Yc3GZhcSYz
FwfOPcfM6P/FGyBgQX5/Usa8hJGRpqAyoEYV1NDQfrc5P50cC833ICS75kEqVOk9
pbACaYPyubQ/dZDbDVAXtD2451+Bin43emS3c+pQrJMvUrHeMvxKLeyTAhPnxuEr
8vwzFFkUGNiiB3Va1SI87LTkPFdrzAd6jxeIZXa0pGDx/r34nQ+f99PvauSnG9AG
EienuL1Z1bdUro3A8oEQpGC7/D8Y2VQ3CKFFL2s+ikPjVn6VprRzD6t6MoWkkg/v
z/7sEtt9qZDpDQ/fBb4VGFvGbVuHRsqnMH1YlzjBXoNLyPahQRbcM1NqHcaTVkBe
n6ovv2MYYfkktkkxoNISIE7vaSQIMJ6MMTEloWKDjpwEIz0glJ7XnhxpBWMqzyd7
gk9twf5ouAoh9mm7SKAj4Lj6x4EVeCy1eyNvi92XjUt4kMd2xOkvQXPkwTZo+gXX
iOux0hdDV/qmtls6RQYS6jg3bm2uJqM/E+gpGBqG/eJZuTGd1C/gmbpOG1L54GB7
dPNE73z8O3c0hzwh4bE8QA35ZJBeLj0cL1vP4UcrDxS75Sz2eVupL97LPd9fYsl7
4ur6uT9hFI/bNCh0dWqLlv0bmNvUV2jzGP6NHG8y+3R1iRKb71ymE4MVJG9uThW9
vIUuMCHXhZlW9MmiXqAiix/d/urJYp7+3E79PuEdtl/8VeFFk3xD273UjlXx/Y3m
HeGlr7NgeQh+KVSzUaOuDCybccJrV//3NwDvepK66ADzTHUc38MqnRsKPsLvUJ5t
N0m8mVls7r74MCbxXQMIC8hqVvvmD2Gm+3F1YjVOVJcAXT3+6JCE4/0fhV1saBaw
TZc6N0hwfc0ZTgm5ci6K4vI2VF6eGbcJJrj54ko58air9oTWi7Y8wnt4LbjfSVSQ
2XwEe7pq//9Mcxu00Tmo+yBuub9XKF/ARwRFpb5PFl/T6ZauG6VIjTT6CPTvi72Y
sV0FmoaObCdY+VkJskWuOX/0nVCL3Uv+ukWHB8FoeVMukY0d1UpAO/R7em2BbaZC
IGw69hgfJkox+MiUyFEOrAKUSqxicZRG0y37D6LU9o/43MLXGMf5zglOoM/8//kn
JGxpdrfSOr+mUQbaRQBuNIWHNjxwETd6B5SfVpILlUjgDEU+k5iBj26EXccUx33s
RPnLdsxggBychcxTC2gnizbdcyWSAw7Mq7MxM6LdS/5C0yEQs0bGAGPH9kZsExtY
yL719o6BCcI7f+zs0z4/O8QQPImgJAZQT5lcjW/7FoCeKnfuOSbOGBohzU3zSuKs
6bCpcMzmfBWA48vI6hcb/MLvesSidKljankPw3xxKzF1n0l/F9XmscpRxL1lVC+9
q0IEQ7g7vjh7moBbsyAPnQPpAM4RKlfloOoG4S6kFvlppYmbx4xFFTfZ4pmQjnmT
gawRpUvG9PQeqblj/Mu2y4QHnDN5i//nsKFpPulqCDXK9pqy7XbdMO15R0igxlZU
fdaWcFctTVVfQJl0sx1D8rbbxWLDEkNYf9MYFdLmz+2BmLEbsnm0pVAtErp8/XCS
2iX7/xIzzpHY9fQBYTIZhDfyk/72E7+rCahImrzxhR1JZppyezu/AIISIBmgR4Oc
wQlDnwmxSjIRw4NqKXGYITMcasY4ATJlj82Tzw0r1kWfT8spMjLYEHSQ/C3Emcuv
XG5Omtj9nqZomN5ZiEe7/hYGEzdMliq5JsPTPQzhKtzGQuZnTj3xwdbANxrZdZr/
aXo9kwX0nWCgKTi14gvqXCBt1gi+JtSwVKsw1NJPzKc2vzTuNHiOHeQmkhkpIjBx
n8emuGAgIg/KWGo24+exjeR3QbvgMR1hpYDKjMnepVqzr5NmGVKTNfpNkAC1LnHA
meidAEg1yKc0XCtoU8fh6lYsCqrRPe46nyvVAZe9PK5dWnuIM6Ry3GQHzaRV0zpC
BL9iuzA+AEGplt3CP9zDRwYCKkimTCBf9RBKpDRZKSb8RoefF6zF8JFZG9mc74i9
KXM4+JPDwGkbdd2CbZ7GHmm/8cds7h7efA2QwY/TNbb39uGzMguDg7d11D+1zlYm
eEDhkJJgiA18sP8YYYjkn4s8ZdO7tZ8lOz2Wcuj/RqHrJ9EQYf1JqLYLDjedAB1X
aMsv1zPnTfrTyRTrprnsmg0UUDIs7Zu6cBzf2EdWP6xc5dlzIZ+BzpgDpPyERrhm
4UcG9bKv2UyfsJBI1umR73Bd1VB7cNKmIDeEn1t34Y4laPh+Rh2FS/sHITvvRp5I
4X6TtS5x6MRfSrhgbPeUrctQ0UUqXslJOkSFBgq4DiUawGfOQsEcH3PhYB8mALGk
eTzfjPCPJF5y6p/S9p8Rx+uS7+0egsZPmUnI1YiUtLwzjtsHMaxdL3HizPRlmoV2
lJpMeapFhzDdGSISGZ5ux7ErZB1PL/ls/+yATRJN1XiQOFhBf13YNCG8mxsh4/yw
3oFyvIcDFVg998wAlrLxDzz5+MxKwgOhHpOAEZxpSMQqS52mCvs0xjCjfDh8VPyB
0+spw9FFvk/zytrmrT6Su4XvZHrCYrwd7TWTyzJ6AuEIzFu0BuxKpBQgVgjAr7PR
Pd6u/rFUCRK5WW0p+VzZLBLJFWgeTD8dRUgDwAb7DwhEnRHtACLT3//S6V1J9vJx
OQ/NEx7yoGDrFwXkRkj/H2EfnWAT5uGA5z5ney0Yt11NzwidaIQuLltYds9l6Rop
VsUshFODZZg8OtgW9c25xfOLomhKgsPKpP2P2Wb9lReQpnWFhaV4W5hpAT6CdcZC
ZFWCd87e4am6yWBE3JNU5Ft2gKU73BJDrTiuEn8HGSiUHoVhLQSrN4SpGZZqZInT
8u3fIF2o3bjZWJNbDH4/XPB76eePo+VOmmq+9PX4UdDlRIjCQwSLMnWuBbdt4e5J
OzwcfI8zzCvqBZyQcExu2vgoEGQnyn6J12tjlipy8D612R0czKC3Jf01QYS9zH5f
lfXM9lFh2nBGdBpHxGrfIAfilj86IDfbpIdwoy2V2b5CUZkikQwBc4mxao/cUu8I
EjV7LpHh5RQjLTjSgDUdBioauvKLKm4Wvu+LT9gC3Am8QS3pBcy2rz63eyTcvl+6
kvDtsgym79oxwp22JvC9iZVPUOdgexiiQFRr6EknQM5Fg0w82lIhPpx90CtjSUM7
+jGsMwMlFbHTDMaX4cC0rbExcmvmlTUfQFqPyZCCgaCzqcKC5mQ5N4IBdfp9igiC
0E/XPAUdVm42pwBaeF6S/YntOcLDgLIj36g4RlB33np2n/vInBRntRRdvr1IR45t
EmYsuA37Eb/2B5DcIc9/bb2H/Ga0AOSbNrPj3Y+mwJ5wvArdVLfI5gid5oWvC7Y0
a7mI+DCPA2F/7VItOynG7TFxoRHtBxoJRAzqX3WvtLKgjW2weE5S87n1E7kTmPNW
gCIVP3s0asyo0/1FjZy9c1a05I6AVkoAxsrw7DZKmbHXmxYgMQNnnHQEz5yv4Pdy
HiRoilXpuQUrp/No9PDjzdRlQOOpxoqx12vMjW4Fmt5udeI00eVsopgA7qo+xPtP
1QFl0AauKBKJP8Uy7KBjApzw+vbHqdHv3+OmAL2Vk+zL0KfAz4WpGuK+acFGyekh
Bm5iQORPdyg8tZqO872fFxJoiogPr/tfYmJ5iNDCyTrbGCT2Xhi0DAvUarNgEOOo
i/NlY7UZpgn3j3tSxZJp4v+nC+jt6ytktLtkxtfIlPLsDbxNyFiN41cwr7s3DtyF
FIDulGy9w4Xt44q6ljHfWTMYGAjwSbsBFtUT0vXHsAf6IfcLj/esXa7fdtmWF5om
ftUYWWtdmAIIh8GpFQ+WUsfb8qR51qIS/6Bzm9F+Tki5BpDkUxD/qF16K2jvjBCw
9CJDrWo0OQq7RvYNil1S5zwVEqOl+nSHV8ijwG1QPZ7N+GJPY5YwD0yG6dwjKSVY
COU31qlIN+T7OlO4SnL3do5mNnjdPFIr+WQOGp247CTGSUh0UTO/q8fbcifp8jX1
+lIMym3jSBzD3+w/mQT8WmryBil14xH02k9n9K81Sy+9vvToxb+ohxb3S2G1OIWf
+hmIeOZ8+Lq3MudD8D15u1DO9XU5L2zBSCtTdvTWjtPdQ3Aol/GlsZihRPR1AN2F
DlpFT9w4k+MgA4r3Jch3V/fl2FfaJrhNK+sRzO/fJR9Y1VKfMWuG+G0T3diesgRR
Yms+3ApeaI9Tvn+8yFqQBq8gUX4KAPdpRu7ERI7ISpN4kqJjrJ8TMA7ol06aX9kk
xUIGG0hp68WZnDoWWThJJl/DjR7GbgMwBkd2jtvcKn5vvxFLJ68n4j0Z15c04iCi
Ta5wAqbo9HOx91XvE8/wRB/wPQcuLMo5/3fy6Apk5SR0JrCUZZ3/NELDW+iN9iV8
hksGJoI8GYiNcOccFnh103xFDUAR5Os1TEYAC24mW+pJVxn3pJZpcrAwt2a7UqIK
W3k4H+F0biwP9puz6StAoSMxoewhK2JDZCtrkoROiWQXzNUin5IJtN9Tfft6SW0i
o52dC9DFh+MXYTv8McMJBv8K6GWK4PkHuiT0LsEP2w7Zq5+jj2K0yfWjF8/sTb23
zOo6exnvJ6RHgZW9a96VwBFn85Jhqu9sDcPJJAkIT5UgfKoAEjaWyRzb2yS+5wa7
Z/9tOMY11O2LXsPnB7O8Yjcnl1tY/ufeyl7mdpB93uRU7zmg88yMfbouPDUVIdjt
xFZCPnPUpKXypnKcbkHdIKfNqjjvURMvO5mocYtIo5KcB8QFoKoHv/S8+W3yHNNp
ZdCmH/MkZO9Ep+yMZtCGPAg8x1Jye/tzndeENOjcBVyTV1RwAclBGHyBmfFXgc7o
7mCkh/nxj7lzAsw/jsF8QIVek9ftMW6qng3kIBI2HwitPbvuZuzYMwpGz0Yml4QE
XfcKvn5esn6i47qDnMNeSOkTJgdhOnL2CoKvBSVC5H8fi2DhzwciOSZnjlZwbklO
4UA4V2oL1n/sAWg6KS1ytlAkrjofy2cqbovfJr2xce18Sp8ailQPDgVQ5BpLAfPy
K0SEhf2HbpLu/0UkPu1zttsEhNe/VqyOHNJiePL7I587VKsPOe8jKlYbm+hQE4VY
C1f7Y8ETAVh+P8SWdSuUuONWF24ZDWwyjiYWKvuoGF9wv6G9pwJ7L8EbT1v6ijAX
J5C6J7zpVDJLFGeczs1wZKaZuP2j5sEPheNHjU2+xxKGo3kWVQoTOmwVfBHAzFjF
SCwvt3dlCdTiydBDd5iKWtRA5PbjBhTaWxOJ8aJ4X/5ziN/brROtrptNHzS5Jx24
A0sfLZ9DXRuxfHuXCTmiM8BnDS5oenaXVCwEveUmLszKgSJ97QsudSQpA6PZRTaM
q679seImYSyPi3gE/Ynm41UjgyORqiqgEP+y0vYk1CcqXpT6/pQzKZtg6BKI9QUr
4JDUIGYfCtNx/kV6d12/Bx2jVIws6jTTbr/k2pKqHWibntSOv0iVz46agIfz2ANc
QWO/aPqzES37zbYatwdOoNoq38432izz/ldi+F/LWXISroSZ4EVX15Au22guk6I3
tnGQLVkU3xgjd3H79QtVJ3/YINj7GPvJG0LO2cENbIu5ZTJbJ3UPEb6V9JZqIK7L
gaa08ZP9t1TLkkS5RVhmZETkmMmMLK11sPv5puk/Co/klvV8F05OotD/fDjDWfoY
JmF21JTNqKMs/3+bqyH6u7Go7mDTyAWGBvtdcme0xAX/rH2wf+gheyLUuX2UBb5i
14T+5Nf1PA+uCDNPGkumo92DndPzD8N4pzcbk/5zSYidQKJdu9e6/tfBRO1i9B05
ATatV8XNnFRAwnv0VeabgyhORYS2wW9rA8xlvlfU98tPbVvtgRB2fkGqMDVXIqqJ
wK9jdkVEkUsB2lKoBwfK2A/PxIZJD3iahjyXi1SLrmzFngmvb2uo/LYlcI838Npu
6estbpyf29+fo2ZPVfoZDSTvfIW9gpMmhge4KflIJU0RsrPcWH/RHBqaGBcnmnF2
JDvdnCkbregh/6Se6cDPo/uTAXu2CtSPcuDsUA5mci+JX4ButvF3PcnYfTYdX5RB
ETD9WNENKj/Mio1hQUKLaTsa65H41xNM5ftErR/WbZARXoql/+BznOBnrgTQ+TBd
W5AjdKsYCBBTweH6C4znEjyUSbKVpm8LtU0+eNCHqHFraSzIw4JFRTcLbKrawDf5
NCCsqU+dGE4TzjTv0fuR1t45HsBqIft9sU0RM4R+xrdyWnqrDWspi9Q7kR52W07+
jKfY34HmY7lmJlkTRjfJYUEPa/qN5qX3Ay0xmqaFdyhePDQu1X/ogWm1KaBo/g1F
Dznr2g9wdzD5S4r092kmDT1TmAlnc7J7WxStndyHeMOzS0tjFnrH4JKYRxaGsthq
fllR8UCH8xSU9PuPWMPvIre0SFOy6YnC6IV4n4pRZEloUw5GSxYKOYnPd1HYKgl/
TnDzHE6upEXHP0qhDMjG0mjI/iry4iHpY632OjY6hLRSoDanjjFPl/h6bgYclkLM
7Xy4UfMtEDS1mzUH5QvrD98zGARZbPXNDuN+Ayc0t7KH797PEMAAvfTrt556KVSK
lzpbsMyAQPWjAf2m20y9LyLkOwjMzn9FlzNJlFpekOaMrjo7h6DnPPNC0OUbUG6X
gcfuYJiTxdvtUQg5Da4F4dDUFth0SruJwzUvyVh2iAq9jKzfC1PWl9cF8Gb2VBPn
7WwnUw9ibNGMhCHVQsiKv0Ylmio+eLuDKLmAfs+gGc1ZZKYS5D3HXqadtNPi+xBW
rw3twzlvWLjg1Fr6Aqi0Nzu50XVLVKqbjkr2VVxErDUvLfiQJPb5cGChuD7EpUre
eL97znRSdEZgBjN49+p2tStk09+/PjeHXcYi3Lc8pYTEapD1JYy6qpdmLaICR6e7
cqSmmqiQQWybMEGRN8A7yhcOhoWTtbGYMJAaEIh/oQ7TzhphtijtG+PHb3mlSSGk
1t5h7ZvO1785UitQ85B+VNIsbPQqdI6FkALi/Y5WIJmJ9Ohhd5tIT+XLN6Rdm8B1
uctQQpLF32BqpUjJQeV4zqeykGxF8d8j8EaYUuajQSLlBodWOCmMvMhlowERjkoZ
TDYH6PjC8ET/lnBAcgOdeABG6P4gqZE7OWefP89MD11ihzw7GyJpi3dykN9JAjEU
5ZQY/P2Evp+u0JZS26mSvtnFz2z1CLgzeZV9+x0HoguSLf1QpgUEYnUpz+EY+8Wb
d1biESqRrEwkmZ4OwL7psx1JXZdWGye14ZCQEhuWBFAKNW/FmOj97YmG4hx2UbxN
Zpl+VvwmxOHaW+BdgAA9BQby0uPSkQLEpaj3oIt23hXwpXy8aTnA9sJ6IxvXP1By
aCdXastN+nEmSBfA+1W9wtrtzbEe2HqBVJOBEOtH0fHbltgpUBDuobylFptRY5Yh
bcbKp/iR5XY1bagN8PXfLYW/OX7tHqUtWujCe/c5T5BlPAYr1tzrMsd2ZbJ/wle2
lNxLV5jXJNt537xbkC7I6smFsJNpEBNdVFyG8puwgFhSupiJ7Uunn33Vka5WTyYx
I4Jl42x9A5BfO5cTpLFBXoYtQm4Og7OCWUCi3J0nP0oaDSgvDJCndlRYT8q+KiCI
vSeWKSirbNah86NQdsQLM8VlsejJMJbPyxuLhiOSuaje2MZJaZ1UxNq658HyCDAj
BapKLZK7tWUL0ogDsXF6xQ9yoKrcVtnsjOhVIH4A1NjG0qwv47aMZX0URyNiGuKT
Njlv/SUGjO6U645y9Qve6GAo0u6VJd97pJgjiSlAntb5Et1cv207nef4qvC46Mzk
Ezc33MLjSEKxNzW2dWGJR4bU5oP9onwGIY7tZp5wU3a59wngpL8SqYndjkC+dKBm
GTKxM1dkH/k4BuSWdwjZQinS9pBnwYAIg1XQpsQpU1GOQMSDc3WG01/vtvgVpowv
OUYW37/QqHj9NA6+6kx0gXQTRpKjJuntNPfXkU1Qg/tI/37SW5Rl39LICZmJmaYQ
FZW3e85Wep91mTbqbxQ02HR2rktTGMLo2TiW4TWx938bf8XS2xU+ZuQmz+dW/Teu
IimTQBtwHUFhF5xD9RdivtDprDONE84gbrOXA4akM2gujYaEWVxYFPAOidbkRXiG
O9udPBapv4GWwLv5TMJu1e5nxSSd/sUbWEyFIqj5fAbe5OWlOXf4C6XzgZRUChYL
qScnwqziG0DGhLX5CDcv+CYKr3BcOFEOs/8hf8YqO0k3ZlyQToC70sHjOkcL4eLt
omgZSN7zPX0VoIjya+eIoB2yDC05WmBxAaojDROexwXxGWVZQM5VewG/136w16fP
BmnLibMmPyh8lk/Oezuc7iA2qamDRULb1UpAjDW8VYr19/Wy5t39+gco5eZG1ZcJ
yN+wJ6Or9+EYkpBYkIWU9wMp8/M929RG6IXRpZTJLXE106wmi/yL6ToNabgu5CRV
aEXcmd5bl01lUApF/W4NN8A6CYTGtCOi0MT7hSNTcY5XpxjpqAkPxjTPZvupQ7qV
el0ZOsgT/mXTn3Lv1skuEkKQ+YEUPYId9jgTXK11NAjuG/aXY63VqDpKZdipp3rM
tOEvxQpEJGwAbg6yTtgcxkL07C29aIdNsuvjLU305RgyKV/IG6x83OxjvJCSrzr2
LlKbakbtUJCMum119NGIONDbdqIzIIhEP6i0jfBO0xW9oDNaVS8+Za1fmb7ufxvm
IDD6JhT/BO2isIJcniQdcyFf7/Jwv9sRBrFiu10dYVdSNzQus/4rqET2W9Gs9ke3
A8lYwMx0OvrLsolj7LDkAfS7Scy991zFnLTTYYzuwg27tba8F06j1hqA7GOkOy6M
2ndRkiJUQNIyDdv4ji3IaQE8vG9IqtsLuVd4Ofc424u8yZccioJDCrKzEOxttQ3h
n9ElE7k4HeqTFXvQx4+Cxy7PR3JmCwHwIbwwyrWc0kl1cuaIqDItgE7cCrjAh2gx
VmmyvTrJ4dSH3cNYeyfYAJUMWXmQNVxXrqNp0QjvZ2nXpUhacxc+X+A2WdO5pmVZ
BsqltpT2GUW0pu+js8F52PEChulCB71/XpldoUiE6NCz+94aP0SOmqnQ9SF/jfdU
J6TP6kx6E7r/+/VrqEKwOdlR9cxulakhPF4OSw54vFDy6YdZXiF7haWGqmTIMB09
igfA2avUMTphhaqENzwLxShUIxAM/V4fHCQgOwdQWfECsFe5l1Dz6DgyCRo45Uqa
DLh09a7CokYFr9mYFcU+eqs7KhxM7cwZB6E6DzXw8S1e7WmoBvEig0p1X2BEdTYJ
inmZVZlk6OVa+Ht/v/Lfd/kM1hVovNc/6Owuo6ukms8rKYkyIr/sMpLOJV1z0WD6
v+dxMrA6YUq7/T3qRXDPjnc9FtUnHehzRuaNMaHVxdCpgMYm8ymMDwMyaCJJFK3a
t9iuBDgG2kHN8S2ob19T++6BJ4Ni6hzikGqwabhKv1mZexcIv6Ipqzy5VgmMH38J
FTu7yY9LANeDecY91QpfYMoDpMVFfrC9QsBkU2QcVfo2XrJdqxcQTJYm9KaQDLVe
WQdYMm0DJwYNS1qPQ9OfKUwMhp8oiLw2XBHIeiebJu4n0xESQuNarEuLCKu8WHSi
zsUJuYSlU5FpNPEUnaDhvKS6O1wNDImcAvVsLiXygWiOxfJ8r01PF1kACn4y0jP2
RsvX3Eb3cO+b/qyYtYbISHain6/apw4wz3j5bVkTU7JprDN8XdzVw0fRJ4BRULyl
Z5M29JcNcIMH+PnQi2dJN0I8ZVRCA/f4SXIsJpmR51DQP99F2plJWLiY5mTUbLab
Apet3hMBmPoK8OogfvNxQaCFHfpdC3S4QLQWikNSJydJF1iAkBxFNn/OC2UjA/Pq
COsGRap+AjxPoUQw/1wO97tUX9+8xPiKgaKgsZohLPhGenFbMEAQZQyuRazDFrGS
flDwItxpcBOEyyZVaIcC6V2V5WXncqmRd8FyPVAf2n9ssrFYzx+yMbU+sPGYMR3B
VEDmhQ8JiSA4l5l2CdtGMai1haPlv0zcpdPhI+Sw+y7b8zgKwLXwTbABnPunpXPO
R1+Caj/5G5p5tabBEGyE3nuY3Ovk6KqW6rQ++NTrMUB80XqtZY1k3B1WBuTiqlk8
K/plfNMVBrcgGbrTeNNEG2OJ+ny/7QwQcbPE5wgI725LT9MdgAFthVXysZ3Jawpv
eJA8TaOO/tiAs6hWTUbpajG3FqJUmEYfDzIdbt+IBr9Id9dJpY1zusb2B4RYlZCP
Qcf09L62EbV5Ozb1gJycg8nRr61UGez43wLcuJu9azUIwcXfnIXvVqNGuxIP5glX
48LgkYmoCDw4vY0Ya66NxCl0FqPoMj3iXSAqlXl0jYUhzEeuTbqIqI6z3z5bOtZH
Qy1SrKe8fLcppjTrLA+PN15+65qCVzG44vSn8PmvgJX47Pd9egHZgWLLZ2rOwxZ+
MfwRqzGkWtk4UG+UhYGGVIfYUqS8dT947xwmr6eX6dFXy/C6D5cJBrJtAJIqv94n
Q8dWZHfskRiIK7ZPdwUrBPTCLCSOS+u9NVBEYFJzi/kcBR6m+ZhP6bBBNLN3cfv0
yUn731WJwJ8EfSOwOMWzEV8Hi+2wWt7t+DRUxhRPlvFHLKps9iDSmoU+qygLDGJ5
DglAZqfCahfsU84Bymxijy1Zj+6uYXfqLA68hswyYxPKEw8DMbYHfPwU2UkrQUf2
NE3rfG92G+Ns2Y510WvyHCDt2EPTStRlWqsX2hIYJ880AoH3xg6WGpbjNCyTbFNg
Fp2SisnIfAgokMPr5sa7mwChR2WzkFDuYrZRCgyjGHFEQOrpC7hs6iTNcS190pj0
M+pV+ScAWVXdTX0AA5efR8W3496WbUf/hpT/DcYi/wegnhm/Q9BAIXs4rydIsZBu
gHEqm/K3f9KI0dBpiYxsK5upJ/aHOL8JsVkLbO17Yrvo34X6Wh7NaGOmOESi10qB
9dr7Rrnp3tvfU0qYOvlE/II9bXC0KUkQ7GXHE2BQaeZOXSWMqYT/GwWAbvV8KUBX
cV3wCm5NK6sI1s8cksUK7tyGhvAnZLg817/CEohc+kaBFOE6PnF9CTg67gPbLrfn
Ge4gCquqaxs1fvs8W5Ff3pSVuK0ums3xyDa+uBVriso1CSb1dqtIZBGr+mLaAwPR
t4nRIvFx05v3XV/8drGhTJpe7i6sG5A7qzCuCepv/WMr5+MJMm0PC1SEI78C5/Rc
wqe6Q+R+yAjPwHQ/PQjL4BzOhpaGYcBpwr9jdrl0h96pUszlAn1kY8JGhhOENEWM
b3nR9yc2YR8Y5dsVlYUoBDi8O5COSNha7l18sOhpP3PjaqJpIZex/WS2LJw9p09f
yBjL2mCL/Szy8aKWCYiH1wOwBMneU386fze2xWA3eNbtUe2srQGDOamlhJ65TrRn
VIzi40QZxfeJj5rFgceEg4CU7FPwCPyoaooSIoqQTsS5vQr1YIedh1GDBe6tbS+j
r7mj0zHfHlaitwO9HuyBOtTPfhry+G7m2incEizAtB7/shabLoadY+BgGAXpBgFx
Hj1jSLDwkdypHj4o25KX8P9puNvrjCT/gZNBrOAYFeHK8nmlc0YG7Cny+egKYlIP
lLCKrDsripLmXqu9sxxZrq/sE+LVIErmkOnyKowuWHKaeVWmdwn1rPPshw1Spylt
IiC183flKfvM+8j/nil3EzAjd116cnzWRbfhnA3tGT4u3eCuCWd098yu5CvDEOUh
f5njafzEe6kBxFhRvmA71DvRPfXcjjgZWfnCYIv0Tw4bSIvVuYwwW+SOLQFxnNqu
vVp++OvJhmFFJPjNPZ9vyuGmqrTZ4uNVqEanY2FCVs1qR1ObeA533mIpHrfOTxmD
nNmcu/LHvrz51rnP7B40fxHajwPXzGIPFlQWtK5q5yFKF1usMd6+D9iRNX/q0fDa
s8WWQF+EHXA9Dx/MGz7xKabs4b8tCCPieankNlkyE/KJIzFGHvwHgbEU6wtIOu2x
a2FauzpIMrGr2ZmQztPHV1o0jzrPn0q5YpBEGze1UvOJM0EubvFpLtuKNziNU5U8
PGjqKkkldMDcJ4nT5cENp1zrOQfXmCdcxZun6/5gBir37XsWwdptbO3h4ymkitn8
6Rwth1IKpgxuK+GnNMsB+8alAi2YORa1212vDQoPuWQ0Yp0i93EXePCgpRcehTjQ
zBV4uaoh4x+TrFZd4jocMNusQxXXufYRiCnPPeS8wTJW7c9lZA9PN0/lb8Dlug6u
scezm1le7onbpiup4BAPNh6AWpqPBEXqmICPAbt0sHSaBmQ7cIKWZRDnlFISzJ5f
C1mGyUogzxfNZlFYMcX9QhK1u9YFElVJM/GnbVp+fs1sUX0rXRik1Gyf9dQ//5vS
VyvV9gp331h8i4dPLK9W9L4LQ1iYyTRW1KntGhaCvuOGuevVlmGIUFwGtO3Y2KLd
Yiiqk79WC4TQI4CSa033A17O+qsg0j6JkX+CNzafTqPrlsbS8lerg1o9OgoeDq4U
zWNgRFX7EGV4s2X6tN5WBRiw6BMGhBgYyzoa7vYZSLggMVNOUxqBkcr51+dSlWgO
WHtPQLNbiNuPqcym3ZpZdBAoPRhemDWhoHvqDso4RS0cgwrB77SQp1iPJ5fhgECA
SjSyhbNzmB2guAEJvCW1oZS47ZKeGGRQC/MPjdglddQIO+b3pWrpe4mO3yaQwLAM
EY0WYWUBjPYgSa5qkYaUi03cl5UzSRKFlvLTxQGUPHI8Wg71XJhXrmJgBF0j/Ypf
DMF296xyIPLPxNaBx84Vn/THW/PfKtN/bTiiJa81c1tQnbh7Okqec+Y/Q9US3hG2
j97UAOyMIBw7hddA9zry7roSpPCRl9g2AWhcuH//f8C98YZDv+3JOp2c3r+n2fIQ
fcqDa0yRkQuinnUOeaEW6SxMI3L2yJa14Y+nLHowd7jwFhS4Na/AVLe8XjxY4dPZ
he8306PikSpJbl+KOaCL7sdLDllnFtb9bzoE5PntFqdFJcH2RRlqlnXWtf0FDRHm
7vwoHUkJ/EYlkq8/nDT8GXAI5omlU32bAU4PB6XzP0O/GjUPYc1eyfRxAE5CTILa
huBzAs37QUs1NyxqobVCixgmYh0tS+LffUogFHb+6IrHwfdiM5FULLn1mA2E1c9B
tURMkwtJpll+1S2XrWrVCJeUY2Rj/SDjnkU07BryD3KHPNfi9uUDa/Jh1OqW5dPI
ykHkEWtAOKJDvy8IgdDa9tD3hs9fB9CqUgZA5N1ntSGBJmFGoe2e+8NPi+4ZDDZS
L2h8GBI4ndPs6SLJKyPL2dbBEdus2SN2b8dA44JDrYdRk5im4s5WKE4GgeiTOTJ0
zUWCD4h/azvcO78+RL31oIBK3zi9+67ouYQGef3mz5Ly8bz2giMl2Sr96ggDG+lS
HU2pjXwDFKKvmq7jC8+QA9O5rPlsT9EePBOxE4iCjPHKLO92OYBuWxti+CX9vENv
VuZw7ttLMcMqoY8OdoKrK5zomErO0pqdw6bSSQ0Ykj4EdHZrGmi1+8llOILne7aO
tNeZ9HYlMTs1jVN5KsQTRfzDo2E/tjS6oOC9WtZ1Z2K4MVE57rs+N8QTtTVY9611
Af/WQUruG75Yo7Jz9jpD7SveqcmGhhB6Dg8J9z25qsEUfygs1PBk1vIKKFzsyAz9
mO2kuCT4I6sOdrLnUvFde3fQB9xdLHc0iPGYtM7Ejm2Wf2LRfW531uDvh6BWMhgs
DUYF81tRBtf7J5xr1iNhaXvZRDN9VOrLuNZtKzYX03VpK1xxIcjLLJZ/ISBl+Cge
iI40rWblD91XkuzFGmEwVeMHT7Umt3QU3MqodVE3JkLTuppAO95dfxlB/jnvDGHy
LabA750wBzI+GsWhFroZPHm+lqKzRjhzUoTOtWdkvRa6J/4UxN3rIRpDK5qnt0rH
sVLpQsc2yyYjU1el7g+HiSWDd/DIMkx0/P7mjegz9+OmgyNRkWNXw4aZVM2XZswh
zabPPwsnNr7JQgfijWtNEKbn/Pab/0AKoAnTel13HX0aqW1duREnOEuUZsxysckQ
H49jimN0tPSQly5V/lJCN5gUXjJBnzvJz2AsWpYhkTIZDt6qWoG/ie+4KFYLolng
6wMtv2PBqZ0SUqZJoEMVHWhNpv/1Zry5CoQlG5nRRWuhbhJgNepPMsaeRqsUvyME
piufVCp09mxk2vj8q/HkCChfPftmsPLcdpFfMRdiDfvlrMqGGhs/9+8DSE235fUA
1VKs44IexYODHWh6OaNOi1zss9pedGsWN4/4wXmydZ0MSC3abDnItsN8fvbeFzAl
EpOBsBWr3oqTe2+qk/pRAEecim3KJH4MapxVU+vEBKpZ+l+eTL24OD1piPdbSlJN
oFytQh8DJhF6LJ8oU+wGrAAXljMINrrBvGDG7xtLUBZoVgF3JUUG3XA+9M+vL6cP
7mqRarJ+WVsDiWsfPDxFX+OB090JKuBnFbH/A+GI5DdKLSZPdCVNIfo9JOc13Dku
6ZkO+heClOR7bIfeYj57A0x0vWtBg95Sup9wEf1rDIHz9LOW7IzG0xgFqg9TLGIq
u1gqmwEZXFqai4rYqmsaQgtEmym2w7cFkRt/z50lovxL05qo6F7gDXojWCYB7nh/
uh9OPsif+SfW3xgTPbYNU6DdyK8N5IPwPrFq8s1jupG1RIkHuMBNBh7YALjOPX0u
X8nHrpaM3YvM9NzVeFJlBZeRgKbvjd3gDdbqRfz3IrX3FPR5Lh9mNrnNQbsMfxry
hzWa7n4nzUyUTqzmCJZiZwFqImf/kIWqjqEBqfwtdGuyRj2pL519c8MlAwwhAjKq
a91NIUa/6KQCWrqszx7dliPYsd6q3JESjyEDC0aOtJvqB70ztvPHKCVJoCgkkwaP
5yhbYdQqX/IbYpVp1sKgZ3TAKghRgYVKi/npoqA8ffwGM0AgrMOnZksdF+kuI1Ux
0V6VA/NwVbVAPeu0eteic9F6seTS7SiFGvQSd7ZbeP1QjWTImrAexkqN3rVnCuK0
C6Mg8VZaA9J80YgdjR6dRMMkgOlHaCp/H4xV3/orPbgHGVH5n+pSDl978dVQjfjI
De6l/xrfyjpZpzyS2RhRGpOpwoYnWwTN+x3LBaU8pvtbcQcwkZyeEqYcRonUZoJ/
N4HtT4DLLoTWRGzqiL1VaSlO0ufSirYEmj+NtnFlw1bT6a6hg1eGx74xKDat55Jq
47PX98MM7RSaiXXzQgYmzr+18rrFhW9mQt9cNNAfRNeqM507YKuMHP4R0PFfKGEz
WP2ugyqHAYxEsYMouQTF6dA0Cqc8pGPO7acwpWrr6r2l6tdprR0jiQEa7vjp82o1
6yVOm7/bY+OU+6AqjXb5IN9Knv3/rsXILrZvkCqS2qTbKJGU9NnkWUQpFbHKaI5j
U0wdjMagnviq+kJ2DalSZJrMcjAyta1GD75qBvFc8xB6D09XOoIMZ6S5G0gcLAzj
sitPgkowR6SVL8DA3OcejzGVFrJMC50pryiOzb4d8zA8fZJCz7QuGK7J0cyrSqIF
ZKeOFpwO2lwUwFkPxHxthSyU6pX2gQwGI0U7SYIMQdc5BSsPakxR+pxgu3ltVuKj
GwDKDLjCsZO6HXrbiARaf3z2c6uAi67LmwCwBkXYmXdxTYr0OL6WTQ+YFqIIVwRb
kNKfUwCbuNYIzT7WYAqBVVQACjmAfg1I4HCHoSIUmr9hAFA+zOkDY1ObiwL74owQ
5KccTr+On1W1zqGnvtu+/vtzCBePfKHFTtFdGLBPOc4JoUvrg9GshexESKotbiwi
O5BMid/2oTX0YOhToDCt7Cra/O7dhfucqVj97UPnGF05KnOAhGwJx1A+nQYt6TDi
taLJ3mI+nU2RXm6mLWWz5QAMZY1yYu2kZ9glxdw5EYkStuYxSk3KQdTNjzvJoL6T
p3QihPMEZeUaKxef9/FziRH9w8h105BCyr19v7wCYMRBQqq277F2WPXPYaDIv+6E
WTQWIOULfuwdR+35eLRnLtYgyGsSXiTXogwoKoXKF4pUd4q8LS1MjmGhT8mJBP6c
uWlmda7efjeXgFqm+QOY1UZ5C0ImNivmOuXCo/Lr2MIHPyHfwr/ISbZRJg61xkPu
z2UZgN/BnUrNSZJEdpHYZf85D7Yxglz4d1vzBEgtVZyw6mqRPHcLjjnRmrgThzAN
7WfKtDA6zgUAzE3t9nLJMDxg4VQq5y100pehAueXEugHBFsGQLYcT0PKQfUhAmo7
3AZCVLxn9GkTNa6oerK/QqWqzxMIcIfRu7XKv4ggaAYwIXPlaAd6ZQxFohaxLvfz
gakVJC4EkgHEWMdxEE+IKeR1knZTOZmCZdPHDOE9xGp5LfO0kyWxO7OJsON689EY
gX5xJ+C5P1ZhC/3gIAjDjkh1TXMW5VG0GlgiJg1tg7moskv+7DCRB5yubSCOEDv/
uJE5WlL5O+TVKNu/x6Utf8CRUdHtsptVISGTy0oyrtzpLAV+scmCuxiWfqPxvjT0
U0xTB1DrRgBksQvT2JhafSQcsQhjfjt+jHistq6PNzFf3iwZ61J/I3jromG2oFIQ
pxoLr78ZUKoYRFCEhJ8YcppAC9hSOOxprp9KVcRYe+4xtVcuudrq3u2Xi9B98Veq
ZQ7QAJOr6K1pk4XLjdTXAThTFPb5tkSkMUuP0lmCJQolYdDFnjI+APTNbFv3AMFs
2WBD156hT1C7SI5BQkWf1jVfoD6CdKv7LHyzi0hCr2GE9mezizIoWnHzu11lacgG
jwweVe5PHYK/9NUf+HoFJXOmh9nwFMYUdL2mssd+WyeQUpTqGad+LsTbWo23RpLu
6SzRLTJs6jFfTTK1qsPR2iYEmvSsZwXjRNNkOPjOoOrhoqgfhZ1B2tiq68hGDXfO
fIx+Jtj5znJTM62H3A9XUaMbOYrzXozETwa9YFW+lxrcXTnPi15IIE0PWOyeJvXL
ee2hqPY9k5LngQdH19ahO+bVxryRY+zzEFFpQtl4P8KIdHkYdLb0Vg07kh09AO9E
BjFy0L7ooLfGblXCi+J0a/JmEh/wE9QDG5vOBo0Zi5r3IVx7zRZUPCW/kJRoM0tz
91tNdKg4l+/5G4fp22ydai2sMfXtU2mqV0QKtksWsTkxUllMH8uTKt48eQ5lSOCu
dsUs+BikIy+MxMOvyvvmETKjj//3WoTSmW0MF/bAb9d+KNH43QW7rjp825prrjQm
/Ig2rwgtnCg8gsmZrU4iUbpxDvuVlm+eF/RyTzKR2dlJ4nz053RrYSeZ26pbvh5I
h9utHH7CnUjJELEb49m2RPbLm5Q4z6O6hZK5NMKxAFWzffMNlE5oA9SwC8BXGh1f
JljstniFes8JPQ9lYTtvFr2BJ/PilCmqWR5AWbSncdO/15sGV7wfB9vyQ0Ak0OCy
/Rc3G8pfug/raIyCgnpyakiNlwMppC7ZqDoZ7Xew2ozvsefOwVSHDhLbIdEDg5HK
pU5l877Zu5jzrUXOmD4h9kAnLTyDP1Myn5BhUvU2UOukoS8W1lBW2mjqEkRKbLSV
QBqdueDmbm/zgp9tzJHtWjFXmQNDKE5Y+1uA/TMD+q0+wQ5kR1mywr7Gtepsk5Rv
1kizJ5aNhejSWB94Ev/2fwm3m834eSIedhHryfx7SlW8W9P74zcKGDZlJbW4vBmM
QnYWb7468XuvXEVM2X0dnShqb+X64Gsqb4MJ/Rt/X31qJJ5HX4wuwZn3uwRwR65G
dBug3dETB+E6bh0LuYOoUKZ5Zjx/uolunBTR467+H9rtqqLdjWTL+R4PNIKihY7z
D+91mZNvo4wWFgke53qkAJEs5Df+ahXW6KsA5PuQiFA4RVxEkgMkGyfhLVsbocFv
wWlJug6mXNjB2yn47yET8MJqHrEJjhNEjn7mVgGDLl1+c7g7PkFeOUmgvyqzzijo
c7DwmA2Q0ulVSTdnQQl9IgDPk7skd3OAV67kdHop9aJzGumgy24YDeWGKxPnNQ/q
Lk/vz2ZXjBb7ctlRGVpWPu6I4SLMaAZJwFXC23ydY+nJsVPJcB7UrLu1kPTp+qO0
5AUPXvs0sbmI6FCRXaKF5VRXsi5VVAUUxMycg9Pmy0h45gQI+JqLvFmuX/LnxbKf
OgXsTIwJv+HyDStqX9wvm8Kk42TesYFHUaOx6A7BLc/cFQ2Jdgn0t4EqNW5b0Fq+
jIkXAzKG9fmkTfXC1qpse+Wzae3l7E8scsm0Cy9XN4w5yhUqd3IUr9Rm96E+6//e
UgbQSu7frea1ByLgZ4NF8k9lJ4b0BLzWtcCV3FRVJsIrTJ7rhCf/d4yk1/Llv9Uk
dDQ9AoMVPAbihLtrdwRxCEpj+oMdKiQYgcQwooGNiwFBA0UmzKmSj2GOoOpqfg2V
7tJ2NAHBpbs3mhWr6ChQjYvxQEQ0N2JjIVU1aDsX3EUDhOGWtsyjXpdpJS5hpe09
9DTpbjFz3YHeY8g0I5seeu/GTsDV694Iomfc+m+W5fDSfzJNCOpQTE7fsXylkNsS
csIedTBoCqEsY5jOg204NBh5UrANfbs4hIQz0smufmVtf0RLgscnAKQf2wAf1opD
QDq+Q0a8kY9w2ac8eQqxnVED7xSsC1ogTlNuLbJb0rKuHS7GiC5T0nkWBXV9nvic
jxXx6epI5kr8N6eX4K/n9QPM3smMGjz4R/cgEQee6cblvNyZVhjxIjKoamSodV9a
cDQYKhq0P4bfSxcPJxZWRydu6eyDi/eoAQFNE1STpFWiVLMKqmNkPo1PQ8LwtqQs
cduhdBTxc1R2e/3PaPI9lwWKaxql3/DAHRe5eMhpdG92Qd4t1p7GWKWCCNSrUQkH
AeJDHv6K2loN8ypJswiVVCgZxqloch3D8ClcPVc/7kuFSEWQwGObEjih/8R0Eaam
mbPVlvnbpmzV0Dirayf+Z6dQswBWRlN2SKDs0w2Q5KVf3500gKiMon7YbuXtqrcv
ih6XvDwPX5OFjvM13zOjnH1K/l6n8skkf9PSirJiicPrxMytFKiqpCg064ol/Upp
OSClcTOQ4M0J85WVHivr7VAOA9m56yTviHLx+ZXOky/Lks24wxq+UdACSRKpL2fP
Cg9tYKsUI74b/ISN7dDnGIMGXv9NAbT3QV43iUN/ow4MKwbU0I19qGdXOAccXNvd
omrkYQuhuleRhLMbzp4srSBHjss0afLZbRPhNhVhbwzg7O9uBNz5ee9+JqgLaUIo
GCAqM+9fi7WDedd6thKPLsqAvrWbYsECXdSPtYB0HQuGqiXnlSte7qkkJnZXPmb8
pKkhHMH/n3Rrgnr4TSZa7BTIZQas2tKoPAStlAN2mson4jHTW+vCrDvlSGtMjGxN
hk9eygZnK2JH8KfXYplc/WmpsMv4mKAej6xiFhLGJ6NMtTrsrhWaXzANxS44Pld7
yycdwrBaaphcnaYXxZOU+1Pnb+hiIwzA89gVxAsVzhgoQwXzKcWofpDiDJBZIJ/j
rIicLxBdyMvluHdye+Ol3XXmolR3P03/VHzlAiXoLupmnN7LfTSsUxqP2jkyylP7
7NfZMkP7OqwHQRdMK9QZhZOmvTHlnBlNZkR2mOaKhOrV+4rSdvrqxXcUrtOJm+nA
0q433val62f5oTn6Qj91cf7VwPMJwWhSByViKDzf0CLH+iV91qIVv+OagDg93+S+
dxIPazrw439BivxZDgN06kc2vhAE0zsIA/7L5KvfPjmRUcGjFY7Z0Z4Y2d0LlgAR
nq2iG70b65Ps3Gg0NwJk9pMX2bjG5Z33ReiXUOhLa7G9MDXHoUWfvNPVxmzQU0vV
VBTtL2MWg0Z7ApeGAyAUIOVo+61uoWA0otIEdeIHYa+koFNHG6QoFF/dqyQXto70
0dEVVsZivHHoocPIBFotouNUnL8PiWTizKjwAeHv9b6rS/AXAOhHveT96vxQnv0f
47SR19hdhP6TYnsTZc3O+ZG08wMVx41Q2wEh+fv/2thOB+LHqatvpEaBaYS5Luck
2N/3GHlNUJJRYITnRlsEsJiMGZH3relG1OxzxIsvNlEp1Yz++oyUnJO6Mbal6VJZ
QJT45bqgDXV5ic2We5FtUACjaWfMvd8lHDra+paMcC+RefIzzukhtO5xKEpPOIP0
9PIsksMmGMHf/7Xhr6RiWjLN1Nu/9v+nY3ZNlFbP9B38aKvH6kTFZyyRTquTgqC7
mqzjZbWJVr6qBF+HLSlvRVtC5jd31+vqVIF15pOWoN0vTnrn/5kyWlw61c3lghsM
lU1u42lSzA531ZPoGYMnutH0xHSb9ikr5IiqbDI+2/azjZyXTpmkh4e1tYdfSLwC
h13zMWRa0CbkyxeG6NBoEowUeW6JMxREobxz0vOehgjiWg9uVGn1f8hFyPmRu1MM
JxAwaAFid/rRvH6r0PCtzxxfmD3AFwLSrbr4C+vTAEK4+QWuQJ7t8kU+OhNYmvRE
VBV5nw4qPBsumu/KPYnzUYsY15YFed7lWByTZJJ/x6OkB7ciXFKJAg3gWQ+4a0NS
y2UMB/v7vBPnzqN1iujIHm5qxmU4Qw0myCLMbtdK5uQSrMrytjDyUo1OuMNrq/LX
ZCr5fBou0BKxVo6YnWIgxrsxePu5p3wH0o5NurlO5iGwRHpUggzFLIca5vKmiSP0
QluDHF7n1fTI45a6pkTzavb39t9CNHVjg+BzYzov5kq4j3zXerOlg2z19XmM0j+X
sPzCA5z5BLVRbv56t78qiYtea+gPK07WpDBsV/o3p3yxfLLsDc5ggW8+KsBvAz+5
JmOTqhEdCXynVFPA5dFb/QPfmgJJxyjrJzW3nfxd5IsiNWmccV17S1Lm7zbpINMr
9E85aThx2Pl8HdqGruosV3WE20tgJ36DpbiGVi7zE6iN1c8gNteoCd6I0+U3Zpqu
6Fo8YUR/hGwjAXlCx0NNuEsbygTw6MzTipw0PvVipnrKLS8NVt85ozUIp71tMkue
nI5AJVmULKm31I3gjhiyGOlBTxNR3/WqDZs9z13RqYDQpV8uiqHL1gM4TiaEPyOV
WYzwe3OZlg75/3U4MVlH9uVvFvxjAUJS8yB0Lpg6zwi0n8zV9S6nDJk8HelXVhOr
XHmAeDp3HqGCUXwgo3ltYq/xCBlBdHDWlanMwLlVXKh3Ckb8HcSEbol0Bo4DCWiN
DhsoDxawJJWk23W78ED8RGMuhc+1QGR/TkiX5SYM/yvKw580yLq5wGDgA+su+T0+
ulf1zbgcWuCSned9pi7BvL7czFVi1hWH714FwqBlcC7kNGd07xlzsrzxXxuBRdOD
MQap06zZXc71B/ysN/hU9Zh8zJApdoW+N19oKvB+hVLqt8EKDJIPmS6p5E6j1QOT
FqPukCcIK2iSPXE4fsLc8EPDmK90eUrg0Rzzm4fsM/SoJrz4K/32DqbbvvwAsvCz
rPf45OQf16vG9zlMLDKKZZhxT8r7CkHMLmahEAopqUqwQUt/ZW4wgFktNinFCDQH
gC/x57hLEgOArpvNPmvFaH1/TIskH8Zp0zGKg6RTvylhEiK2iWw06REW/fWz71QZ
tqg1PPpVKvbzMrKD4GWzFM7yZEEhgBYYwI4NHP2HDpUurUNhvUEaGvTho9n7zz4x
6ZH6+D6FZv2K7xecCwaI8EB7BaaqYnlKLfVrMotUoFN+7FMNtZ25NWOcaPVxi8Ik
ofuZwOSqq27bUmp+HPPUc3l5Raz3GGuDMXiLD8D+Gje6SHFEB2IDTPiV9n/SpjUL
4KMR7x9swP4fLwke20YlUnvyO2aNN79VIH3pL76bn2BbNpMgOi5frfjOIg7vxeo4
67H7yaJQBymJPQXse7VfM1782DEI3maa9k3lYTaSzx64Ij0KK0zR8m1leQlwuDuV
mMoErJ8fs5IbKnsYGM8cYkxv19v18lUGBOEJRkuQyT8/+7ATrdEIyUO2sAPra69z
DVcCbOOhb8qzlDCXJr0Md90cFIY3+7b5NxzDfG553TJ52QhqkEjhotxn1R+Anyh9
REXsTRXeEGT/NA7T6C+d0EfSXrrQ3A6Zy+BA6SDPg5A+KepS+hVK/QlOQvStbQKQ
kwFRj66ZBq9Ynwy9jqpoIC7IyH+y7XBNIwznciVQ4DlDb3hj+iWNvfBAW1NfGnfX
COzjBkjpTkJPK7HKWz011VxPEFLCyZaH4IUFzYKwapkyjbeptWMNgH3PZ6U35vRt
zkDqnYZaKfAV604pyp0FyhSElo11HP+eDAc1x3B+5q9Ilsh4XxXggW7AP0c7DaAG
/Ie24nxMauucQP1N18wkQ/V7rT0Lkdv0lai3U8U28MQ5o4TF5fGx/vM5m1mek3B8
6r+b42Wkv9wCTuvTW5DgoCQnjB7FJt2uwjtEhwePPWjlsZbBRY5dYh5ZbfirMUv2
cdxHNcxAKaAV/1dLuEOnAVKBFIA/KsdP5VhTvrPNKjS7kShPQNK/oFKtAoDbcqjO
b89+TmVvLWcOhKEYW697bnuL6kEVvj+w0zIqajjpxT9857Neh4lWAC3dO4jUnqyi
mAz9Uey2Cv4H2AE7oXKFITclfmQ1urAR4wNrjOOLPGxlF7G+VMZ76dfuG/+/6wLD
z6ZZZEHR7r0HsFi7yfjk59Mtezxu7lIoffM/9XhHIHPmCLnRayCby8vW0nVuWy6y
409l9M148AdTauCTRlww1xOwb9uqs+RY+oqNkSFfpXakflv+57oHEe//08R2c2Sd
zWZS5VM6yUlQB9wmRBkBmjhAaFunN28lftDGWQjOGEuQrr7qzay9dqIsOPBOjt7s
5Dq7AzizJmVfyoJeloiH+BPTUo3Itcu9/hvLvfsKdUTP0zZLdVdBr8O0T93iwzpa
CDWBMub/iTwnjWCKDqGIr9altL6UG0xGjftDxT6vNJITu/3L3aXaDYgjzqA0ZFP2
6kIv+2ERJM4T+m9UGMRw3qt56G2YyAv5DH8h/frCMk+cyX0hGCIIYPFGBaKQsC6E
WtsYG2p/kPTleOFgu+et3p8HtcNulqT1zw2F75OMV1A8yIaUAT2sTW4CfQdEWGKQ
C3bZ5qyQ85DAA062QZNZ428QJZJdFXlCCi1Y4UYl71CIK5/cD9/4ztSjzTBcth3I
Jx9Qd2mP4nIbr6O8vIHjHEy7DiqdoHOY5old6VVS/QjYFV/OWLZU2zeaQ68f4yCN
Wz50nyAK9RisLGLRbIjSeSoahC+6j/+XZbpMZc1mGCj+H7crGwV1Co7Ghebi8GUz
yl+fAbRsQzgEtt9VLaE1PbpWUNUDgpUc6ZA7/jsOiJNQXrXF3wXmAa3/oLIvKhv9
rukT7xkfqEk7z6bQcHv8FtrotfKBepQUC6GHEB1RbP4h7vJOfzPSbrxYw6y/G+Ym
7ZoQk2l3wwPRlen30PffTIcAXvcUBWT3MKo8MeddKEU7mzgGuSin8FxrG5AKucCg
HQOAXOhTswEV2XdTTQ4PrYmTeIsvRR4J9dpWuwqNLm0J2JeAiXs9o38hRx8RMx5k
K9lKQkhz/+AVYZpvLoVrjs5qPBUx/vLlrwLM0EDpm8IYEz9nNjQ28KKyhFvsV+5B
ULmYVtfaPq6Ymjm+lrtPcYlbsqsoU6Ly2ijy02ydKzaF1OFpW9o/QGe3ZStp8bvx
htGay55OqZaSbUT4IPkT6eSQccpMLv+biROyfKnCFwMyKqsF1ViZ3SSwh6hDfQMI
CpwFRor933eZIYX5KSJGrYUX2Yp1qcLvKXVmjuZgjK6mW3wYWj203u+IeW5o/N9R
L918KxvH64psrTQqkh/AYjzPCrTDT6kRjmicYzrZp9UrK87yx8BmmZYZS784rAsy
WeCWzHKRTj9U2c2jmlFdjK3J+DXuJnzjSvIgWfcEE+tg6Tv9taBl2aKu1TlfYtDH
AOeiBR4RnR7N7W2ocj3AjlTG4bKBSdwKv/aZ8EGmLSE9cZxj6UdesF6nzehJbUYp
7ZXm8fbuVicSu8qA/uilkoAnZkW7BrjxX7oXm6GqCNZIBCY2fsSrV0BGipWGWEo0
4Isgc9SCecPyIeFZvaDtfWZ81tP3UnfR43MNFJ8ovHu7Db2vS/mROBPzgRJpIqFM
2HkMdnTevdNfc5GjrbhnQ8XRe3Fb3R4M8zj4e2k0ZEeoWPpddk1MmGg22GVXcqO1
HyzaGlkk7ThPAnzt2gNCohLnJdszPX/R/G1bgkdtbiwKrpmvUrv1KdkoRxYg7Ylh
3+nvUorWCORiK77z7wrRfIlFFkbrESlVPXP39qxOpvzylug1+slYfkf7Y2RB1yI9
Tt7oQSIh9XLmtKy0ecKi3l9133wwYJLE2UgnRLCm2tjym4uZpVG5e/O65IBi95ah
WeBol10FqYaby5mBLdIxFtoIJhSSFabVzDM4Q6OzpL2WQxKG4l6QC+pxeGfQRVEJ
tZFk0KPGJvFXySiwoPU+8byh9c72WTcAa5SHIiIdSJ4NLiZxkujyVxfQJsJeZEA6
pslIgu4uhGweI8EFOAEWo6MxfnzyoZStRx9wtU0lZfMe+wUkPbXAR7miJe0fI5wL
vY5Mj+L9NPHE9vz99MfZXThndx0FELHeoX9lUqN3P3PbX8Z2ucABeQOqLwmqM/37
KxWKZ6hSYVKbkonjQ3oMbR+9vkJ2wp1RqTblsCAeRrTbvA+H24NKmfOdkcmIq+xU
JjnTtnUf9D6L60olx1jVyS9/YcrrEDUhjbQ/JQbP6pNu/WFLBKWxce7xXi2gnXOK
u5dhSztg7r+/dvNLeFyQPVFlUZhzKrJwvb6A0dro3QMng2WcSHLKGO8+axFAl40E
MnmWIe6KTDESccQCaZ/slK6sTCdlI0qmuAOVA7SEH7jndSA03/qWtBgzqYIP9dgF
Suc3ltxg6Dpvuzd0c0cZHApTrjDJyCnNFbNtgVss0FgYl8ROOnEVZfdUfaix8Dqb
KKc84007y2khAkDQXS8zEHeyEI25pyWjul+25y6hyeBoWAn1BC5Ocmqxh/hPmGkW
vtNAKTXOKZQT6tHxuS4zV98rCCqDsJkSy1Jcb6BDe2EURgpFcsM1P/pckLbNm6jR
hlurDP2Z35Vi2gWS9ZlO99gJvfhUmJ223Y0GgNTm5G+cOego9d6ExYiBTCD+iuTu
B4k7TCifyEO9YGab9iBOSy76URj4m1SbYnbijaWddLb2j9TZ9wKNuOmvBfIUH1+M
B+Ugbyyt9tioMtQKIp0URY+JmIfeZzdZWeakA58AYtI/LIJGZlirUt7nP26rCKei
sKuCxZe6CTwoEYL6pStEKzyChgDmURojivrZ5sj3taT3WmOmR4lhPILE5rmKrMnN
FnxRAeADU5O7xzD/C97FVZvMlLaNF4Bub6QIxx6pfhhTVxPi6Qvv6Z24bmnG0iiq
c5qegsco2WqhI2hEX1478i22jWruWVUDKl7zpRI3Jy/wo6PYgYtvOdnuxEQv7ZuU
kgl5GsKRrM0kRg3dQAact9dNZ0PmLbmfYPqmceF4cYxwu8RSNnnjiGW9lnK5yFeh
DLgb0V/u+u4gBdbd/1lOdBw7Wko0WXlN41lqNx1dPaeavxWNnXuJjXcLVwN+VnQE
jf3F0oeL6buyN35qce9hRiQl5cfzYDx1OxZjL+VdPaJwueWRhZJIFszvjsL/1x3j
MphpkDbwwJ8JxE9JID2N/nKAJZ8yGwMcu4sIXox0BOr7p4enuCa0sj1Ke2kMmU+i
TELV5ghT1hT6dSqfVhqpF5wNwQ0/wl939q1lLctDgB0W0VIRzFFTSyfRSQJXhiw6
3cRghLGUWWSi+9zO4pF3RHtlow+BLOc2iZi1U+arx5ZVx8s1fr8grU1AIzNCS5ry
cmQdWV1m+kKRWWVVx1bkK7c+0ghRNGC+jQFeS0N6iKIihfjW6GWE/2l2PeP4kqX3
KK4uXDMj4n4cfb6HtWP6n7xMmufmXvg8SOPRLAB8J7SJcsz0ia9UAlHfvz4BUhw6
q+DupcQz/tC0k/Iw+Tt5myDni5SyoeRXZnZTsyoaTg+KwU7sG7RlnVz6NahM+2c6
C7mIaO1+v5ZzloLgjsz/a2oJV22Ykzap32QK8A1GenQLUQgVkVyv7p9J+fBrpA9e
oULr0f8PAFRf/IWXNLvzYnFEXcrT4Rt2EV1o7f1bBjCiAbXr/7mSwnGPN3JWasTp
AO3tfZsFSyQzhAUP71b7WyWB0zq5kR2EaOfzgHStXCcxX/6z/gtvek35qGKteAGv
zGr0E+lV8V2Uz2rWYxWQdQAkeaetybUpBCueh+lV51rJ4GW2YGdGFyLhsLKTBjld
ZHTzmOfsj/TqnrlIZO5FEwIyRdnwgTRpam4QEc/ysBngu+PQb8OhXh2N0SFhia97
vJezPlEGHt/mh7NWlJsFX2TybmkhVBsi7ub4W3AgMCXyRGN3AlhkoS5sqCw2zFjz
NKAz6jNNlaCEjzJGkg2Gx+tnwI2cu2g+sK4n359vp+omOgxWm0v0GAK35nrFQU+y
uj/oZ9w9UcEGa2ehGDG8/YxmjOPiARQ39YJM/2Tj2rsJEYzlOEFal5dIvq39sth5
TZLIZ5+HLX9ScvceTW4HVuNGzYe9pNuF7OtwNinaAskUlrEZMk4eVgN+e+PPMKPq
Ba2dWFDjYEvfk4yZoB/ogZ5YKKEmWBPHYCo0t/D0UXcKE3nJXV2xRj7P5JQD9CvK
o+s2LvB2024CZTiLc+UnJR5VL0GHAXc8qnX6xwJdpgbQ0ePNAwAO6axf9Pwzy1wB
2bw8P1fdAkiEpwA2KG7gvysrcXeFMpbSi21MGmOPWhKPgjq/d0gfWFARzYOyrear
mSxCVGOCajzr/jR/dDlg2+k4vMrFkrmgN3Zoa1tabu5hkwZkQrre379ot6fittXg
Yzkrc0KoKlrFnM9+lLKOQZzyN1G8YBnLOesDIwfhQWvw2YF9aTL+m3Cbzu+XXEmU
8V/zOfPW6ILYLb1g96nBBAmIA3uelcAPN6fYYaSd/2qtHvTeyerjieTeyADXbKRx
ITyq/eFG7Dv5juvIFE9gtjKr94XJncUCPaY2gX1mMb8NZBjGhixsZRHdm0tRVmAx
ZB6FIi+7GmawhnUi5p75auUDO5552ZESG9hNMbMoPRT1qS8w1ax3xOI6lAmmjtVG
>>>>>>> main
`protect end_protected