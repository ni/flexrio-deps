`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4320 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
Ju3IpcJpVj/VshHyynUPTAYHkqCG+zxoaJdVRpY7F9msVL/YCMoGx023t3FwXRtR
O027Tp7/W6O/0lwwLMcG/3jC8DkGVpcf6PilS7yJbjTOtwz2SQy2tA3nK0b2YF9V
yRfxMZ9DFli/pii1c0CTTcv9CR3z7TkyRtKFWw+ZYipb7uxPs4WhVH65XAEMnd06
S9apLYwmyt1BTFlTyFukx4/8fKVUXVoqMN67a50KF1qsJAFSbtAfxGtx8i1DKSkF
uBsq7k70t8UMjGEQfj5xpvp0fuCIdR3MwFBZpCYJAeljpbSqwN+nQgmeQticKpGH
FtXXMkOWSJPL/cgYhaOeL1g56cbxs7Jvn367R2EzRQ2GqhlKV8mdzAf++uXoopWb
1po32gU88AHXtsRQyPT+BAQCoMrA15Xb5ffl0qKaWwnQ1WrAuSaArG0tgcM2FDjW
m5XMFKdigB+RffJV6LpqN/xnG8vKO6F6a2XN4k2AXbepv0IFRa7IJTx/W5NWPJGz
9ZfPc+HFmEOJdCiUxWnWlhqWC+q6NYF5wyJAcY09FrJiNT/dqDdfqFNRpmU8dols
DULcWDmFvjioaZM/e8+s/iDBTSuoyhPoGpx7REbr/2jnhFMcI0GBCcAkkC6fFxJu
TAYWhwLLVC2/+4No9ISI+BgDLrLQ6sZi8iONlcYRYKn3fy4iASMVh+TyDjT7NUk7
SoSkak1vnEFLNfO5HHu9UkwHgObc7itIUoW7YcJxr3bTSAK7WAOfCa9/79/XJeiP
TqXzqhSZos3hQcC0t+g3bnWc44xRkNCe45H1lPhcbyrYTxczgWzzrmKqyd5q8JV/
JpSCmLDxWVE531s/rtEJGyMLuqR9SVaw/RSqNgkyg4srsZQsj9uTTttqcDXeRnvL
xcEFWlcNJ0Wc8MAJDJwrnfUFwE2YJY7A+G8csJ80Vh5YKEGY7lXHr0EbbVdSIWCM
86BaqUnLFYi0uVX5OiS6upTsWSyP52IMPsfcDawrE7iGPbhYRHnjCA2iHEEGTUpk
Sp1PjzUSvRDqXzuoCnrveXc4y9yvAIaAHkaw2yqTgzMJ4AxIgDyL0SO4DxL/oo1E
a6xlPN7tMmfyRKp2gO8wJMNMxQANLfV7ve62xARDiwzj+hUPewzs7zinkIV5LVsY
Yu5Rsj2bux1fTglBwKmRSYQbV5qgsJfucGnigho4Zn/5l+2ERgqWIKN30JPnPBVs
38PKK/zkk/z17FptrrqBffwR/OQwu7L56ZQ216BBj8z46Vso1jVi1f3kprwcYB0X
w/USbQUU6dfOhHjYd6u3NhDD7Ryn0pVEGGmMZOHV4L2HTQG6k9JrFLvQxgP6wBBA
AnKo2ZKLmNWLYc/H6VwhCo+TBudQPZCYtS0HFYomjXp5Dhz4pF+JFYkC3eZWp4+b
lsA9aynmy3aT491Y4galoK3F/l77XOsJ3aDAQbCVoU9oBsJwIJfVAbXLOK7/EZ+V
ajFxloCkDQVW+8BEtRK1f+WcrXN44olhc/AONaWFPOjFctrYUqRhSsE+ccXiI4Yt
igXG0K7HUJYx0qKhn3ES8geeIdDgmG/Q3CXLh7Jj/Lqk5Sny9EiXjr765NjOoOtr
ZAYj6BU10lPTVL3T/dci55MuG+xCZ4QqGtauYCMflMvsSnmpkN11qpJkeQ8phcwO
I40tHyU+Nxjg0ZZQ68BN4PbqjzcaLduO/2cBVtNw8yAenu7Vey7bpZ/4Oo/FiDcG
iY9EOWX8Vv2HgrydMVcmuFz7TsKmxMf57fatkiS4M/flYDDEzZhebQ/6XFwBvJ3r
cpB9lG5dO7Au+IBBx05DsQ9vtDjGWvtmE/iqGCgvON8xntWu47Pa0X3rkx6QUBi6
ODDxN7GcThCV0Xhwxi5ilRJw0sVGhPPzJxEaR+MMBll4qKUVKgvEVtd4NVWB/jGS
8bCp1vy+SQxkVhiKWaoai1dUYgAju1GJKOeqOShWDw8DXJVzN86Ny/okxCxdLlda
xuUrycJxe4Nom8GgFFAv7CkcQ3PIG6k3+1cO0iM/VL0U38gpepoAlp845RHBnKEK
7qqD/LQmw0I4tY3VnvAg+aBUFKdFN8MtD6emkRjYx2M7M1ckkvZ/WnaOiox/r2O8
6VGvEVjkZ7CittHCADZpj7/NQqVffXRvM7WxRsWm7LwH0iPrRBHqklU/y2J3VNBj
uboarRKTAyt72slmlnJRfWUeEWqqtobITH/5wD7VcXa5ZcVWUCoWGVS6CBsbGYI8
19PaKWckDG++7toMdO9w4ISV4p1hAExT6beeFbgEqEpTLV7ZwegySDkzaqjENoNi
YoMBU5EcMMdRYgGpOJ4rzPx71OI4Jw7AWOCHPbCl53X593Ipti0tDpFXe81aBIS4
2zdWcPUANZeaqZto2kolZTdwYCcxugO4Q9aYwMcKjuvFuiQ2+u1kLSD5awsj0vyz
UczQKq0yB5IXRcAxph4ePYPqYIpFaO6XpSuL3XFt/pnwQFOVhLzP7dpWSRyIXwu+
OpCPGOnS4OJPyy6NFjYx9HJIdOSlAe1STmtHfVFEEFzl4F/quShF+Kjt+Sd3SNGW
asAYH19yzjWrv3WcvR+1dKhcwSm0+fd9SPs2AUhNM0CjeaAMYb+I9N7NjHmj1I3U
8TDSuRVleme/sVtA0bg9DVaL8Qr1OEL4HTo2jK/7BU8+piA7inRlfTnpOLsib+E2
ZD0/pQIe8EX1mDG1VeEAgegL+BCSDL2W3AFwuPZBN4uU26Pptkd/tbn3qMUEbMvI
+bPqupPJw43/a0fR7azhZyf6UXpaz2vqOOZKSVCekXqUZ7IGyTh75fQBE6kpuYsM
BZNDSMwb7n526X5KMjH55e5dIZ/hvGNIPnEXUyX9w6due01t4IjdJixjjEldyXGd
mi7f6cgdjvJ3rZDcWOb5+GZiX7dePoxM0HUr7LfDK6V0FPmXdp2zg2IQ4bG72Yej
WfeZfSp0sKfQ2ymreN8qimGazjpCLsduI5GddbBvWfDfAU83SIFOo04QJLcNb8SH
m7GfK9vjxMQdf4oZw1Mlf6P50u/z0jhpU+FximuFurU/pupIhKhNxmYoAgvRaFTn
fYozWtL48uKw92sTUmio0KvRB4nlzudfrQiaK5Ezx0bsigfbakENiqh/DzmOy8nZ
SCj2G8VjNNzPnPuIMo2cJgwyU0DO+MdwhisN8MCXhAqpCtz3dPVdZmaGJwYXMBGu
dzmTaUKhbMvwM5qo/wc2nmYvw7QefRh9MXGL4Mq9bUJBDuXG628/VJny8AfO+nSq
5fnvaeL5W/kzOrRnGiJrUwwFGjuvCJLUcN2FLss0SMd8dbBkL/SglXL1meAWNRsL
sHni5AjRkFyCqjjjFJxyJpEczK25HZ/ctgHOpwZP5vsqtDjNYheFTdHey7QxemIt
GcrKAecRmVTigCuN/aRGfsuFSN/xfukY4imhfOum3BJYA3nlhK8GsVHIMAZQCKly
cFV4nuoeuM8DvbG7RSkBZqkpcdbg194xBXdaTgaSZFeuNyyZ+PJcOIlD/ntkc51Q
20Y8HvIwv4wn5iakGsqYSdo4eOeRJkGRFQkuaSHbHGj2QCdhzzU2fzhR0NVMf3kV
ReWrfFMkc9j8TXcEr6pQqQ3HRgCKsMFYxvpVJuB3ktu+hYqTogZXcXZRLLRHWkCy
o3sAz9jCztTZ+lMrYgVnPXa0y2VZoCCZHtq9NURGsAbi+GoRnAqfcTJ6NKH9MgEw
ogvRVsWKkb90tdsV8MjpVWVdsNfhLAVhVfFukQiJDuAV5ZpasWWJsDwDi9voRE3d
UoKYON2wqHBM8uWuoMkf8a9qLJIgu03/ulH/AONlYdey6QUGLLy0M2UW7FouFOf5
mkirU52Shr4qccyJ/CAkNsw6Ybl73DuwydFJRnGV09Qlt9CXaZxl84ZvrpJdrx6G
fNQFIQ5lX/BLpYEWU/eaalrf7GG1xdDkDYwfH0/+cJa4lSV9s9KBcaVXzwOCM6Sp
2UIE4DxlafDflKhtT4b31YtoUWPIUAROySxM7Nd3v1988PBDnXHJt+RtdUcDWdJf
ju+KvvuQx+ye2rBndMYV6g/TVEVnjDZJY4ixTYimWW5OZyLGUxcot2uq8Md1B/2Q
7OaVdWpRYAo7a+5E1y/xV+tyRogk3mCYUXKlSwGSRJ69xjMk+76OPk3nDuqJmphz
bE5zCrgDuAmQjFUT2+IwX57RfTy6Kzqbki6K3WWEuiWjOJ5dqUzdl3it74kBAB3P
74HhbVRMv0qlq22EqWh8Scs7dEhVVCIUsi0Iu5Me28fjLeh/TGp6v0erVtahk/SE
X0wrM0sh/TbqkiP8lOzwmALTjt4McusPE3kT1PqFUwA5ptjQo0QJvF96W9H6r5Kc
8YB8HbmhMUSTZ/ZHOa+tktrExdLMetbIoJwBC3+5HnUEQzDCmGfaKwRn/9W0fkbJ
UkREE2FuTlzFnEbSkJAsIvMzuyajIUksBrNGI8VeKCphbw4UY7moKXs7Qj81tr6f
VZL84swu5ccfL9TF+YdrC95qwG5mriH4DTXREoroy3ZBw3x6RMib81t6Yv+a/Fon
rZyOmStlVFLr6Lerv1s7p/O5lS7wIT14VWqAwYl77JH22M3PZT7pYmCiYcPszr7q
ukI9dXssfvmYCUo66gRpJo/ROzv1FvtMxpkizrkNryMBbp7oQl5+B4vj3nODlNqg
pgtgBVgFUioKlKbjfO+HYeCGKuBhJL9W/W5POix8UrwIFMlijZk53cqOJjIythrJ
8/4JUW0Taw2myD3Lm7YMr0JZACAbVukL4bDwuiSKOUYJ5c7kewlb/MoHw3Q/sUv8
LtJd1GxVIloFEpb3j6LjimgdfRp+l5N2gXzAn667SSpNkx/6xdOHx/yNd9FKTWmV
WKNRA/jPWfGFCH8rMwMUMSoNtop/q3MskMPo5I7GstCkRTv7i6E3UIzHFNOc/79z
L9618he/NHTVDMh3gJif/PXiuq+uGqYJG/1UQZeLEHuK4MbLf+Fgfq7u50062Z6A
PS9IXAtTyYfbwbTUI/TAcWu0Jk7bmpKMMrZp7M46nEsGvNeomctpLEZ8y8EOcuTo
VTLkcOoxQOjLEsZb2ZBEG8MBPngDJuTWfjhsfqjR5b/RfiAo5c3xVZBbdvJWn0mw
uCwo2xTFcDp7Il3fWop39T6vtHehC4dL996htL4YZ16RochU6J7ioi3/9CEELa2s
bOqOBUzRnI9rwZi2wltT6MKmKbm1RHshpL0ytlZXuntZ0zfC9LkKMGBUAOCe0l2j
BkJFGIp2168GRI2Ee1mVFFnKTP4jted0WkaUtb6pzHYrDo2M54e11NI5CqT766nw
cVc1wD50a7pCB42KGoUBpr5PppdnBv6lYPHvNnKu9LEeyONnv5+CQzWAnLMyd2f6
h4H+9kvI5vpVwTxIQZDUC+60RZJTpQ5mD6GU6rwbv7LNcCxH41RFjieq1y2FmFOG
idse4atQpvG11//YtNYGtBKOyEpMY8QRrEQ5afOWCy7qUgGp3u2RE3tB/ylzz3HY
VTeH61QpfJy22AICb/QhdkccJ4bnwtOI/Wqy0pvL7wXD7H6oO3dc/2UcYDt3n6c4
mHzKWhfCEGVgSnWXTty4hTb+UVzvGWahYmrpzW6D1/lW6aH+aC27/NOnKn2eTK7j
`protect end_protected