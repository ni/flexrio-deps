`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aMReDmrPskJscpWYThVKVItA5gecPPZO1R595p0GoIq1TSTG+UxXhmmUXc+VYHJ3
u/C3EW5qePLufxmXxmhmDnr9U8/cYC1zLfk44v/2OPb1TBrTsludEDQZdGNWeV9l
cPUMSIfZ0dHXN7L1M1E2XtgoTWQxf3VDHs7B7lU2y9Rdm/ibz0fWMow7op2nWdD8
gJ4QlNl3f9Oiotp1p8vz9RFzzZOF5gBBslZxcTF5+z4qO2W7+xLByngthWm+exIr
3Pzy8qyUo/m2DDwOz3VJSvSNm7RUq+0/yJNOOz3jr3j7ZyCj5OqT/jDAWjJSMH+i
2402Un+wDMOQxi21JLo3cA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="5R6K2aWI3OdbT2A+sz4o9+2XAInTqB1/cSw5W16RnA4="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
Gm/2BIZF5/H5qen8uQizPH9RftTuEE9mgEOF0SqeOKegtP64CfvEUnIxj/ahmIpA
6xUR2v2l7E5duaLZh39Mc1GYsfqE91NCPU5whLaBPg0UuX4cgTkO4cYbW/7yvcrd
4wavUfwXEp2VSiN7EVxL8RcZTSMSI0Jr/aojiilFqVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="TEmQtJ1Dsm7TOzpJk/CeTSSFx/zKExk04H6I8sT4Meg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36368 )
`protect data_block
nvPqn26PC4XWLLQG0Fq8XsMTlhB4evbpiwGjZroFFLgtNlE6bBjdtwWsB89WW4j7
jNfYbKN4sBv0hDeMH0AAR+8g+TCqoX7yLdIUd7aGwBUZJr6FdDs2wTUxRkXFYNTL
V2foUCw8RCp/PMc5/qua/vxlpjalH/10GgIMyhDRgP9jRzdarXuvk+F/iCtI6bso
TZzvYTlDOn+9H4YCGOslxoiZ4aSrnTpZod55oKGWUF+HjlNws3grFujfdfZKdZ5U
ORcoOkmVSTasmazLEVen+pmt6OBk24AIlCNZWgBC/pqKB1TC9BhOwBTqfsuZ4Tpz
3dQR5+j04cL1tdzkXoyJ2/YGC379SGIouG6QXvXVP/LQqXoP1OghPaDTkihXNw2v
8NlK2NJ8ytl3GEMyCV5kEQsApOLzmQcgtM0/7pd8XxhH7fX2IGFr2PmBcBHnFJ0I
TLrK+LKDrR8SMPKz6RjYR6hd8TTvUsEV5knGMi8Ji4TRz0p0jBerNMqabFwkempF
B1QQVmizyfUpmSoZsDvoylB434atx1bIWUHlPC3G9ASmtmwdyRZkVPil/1n1Mzap
syYJdW3F60+OdT07BDiF9p5vgcIfejDfwxfjkgymt3F5/xcWwjaAo7uq5S/Oc4mU
+dYUMSaKZC7hZVOFQwk7gHJ48wYkZFBSB45oHvzAW03xoTdBEN+hdnNTixObmlqa
hvRI28akOKfSBpYKwxRWVXyLyPPdb7UVf9bK5SdZY2KMFQqpd6C8eMmcmbDfbQT3
MrdDD8OJGTpQ4AYHNgK5QdYm7BG0Aa4PPF8ABby9OK5T5n3Zp8ETg9E8PRAjWT6L
HJMxzg5Oh6eNSQi1n6B/Szlg4r/lVnlr2AHWQXFWL0tbet1mV0Dofks1Tlf04ho8
VFRwwEzWmGleLuECORv/hqk1RtO32Wye7SzHl0tScyfWfxveLEO98+XHikJaMMtG
8nbloR0FA2hgE+URvBNkXyiXFFhatcrNweebzrb0EU6vTF4GGNzNV3+cUfg0zc0E
v0TUVOa30SDbgf092pYnW+4+cc9uXZMq8ZPV0H0hVtEJPt6x4mEx7iSTpZ2k5pXW
uFhHzkSpccggCuxnk/wEHXqcUhvckBXmbtszXVduEBGu1ARvUq4cJBez15lp+wLv
E0/VO+NxvtH/RDwPmLYzv+i2F80YId6r5XqR24XZ+OkoWPrgSrf6G8tgYfYVgCmm
emhFBk6vy7f8Qy+yJ0TDQKbiI3qWSGt8oKObDYfRUh2RAyGwIiQjI0SmOKwRAr/7
JWFzz08M5CDR4DP+86PxP6z4XR7YBITgvMKI0+i5tM3ccxEtZKbQRjqp6mSMSFDE
H3/+0AWGMctSGdAqXuqQyrjIWatP+nsiYDEUTIeFDK6ySVwGNm24nzwJngoJ19t7
Cx8VbEwIdWk1YXnBAWJjTrKMJC86tkLoVdluhEdbwo3JtK4/KqksyhnL0NmtftO7
/c4mqaHLSr9+F8eJIpmYnUelWhDx8fIh+u9oRv+MyAMDXuFnGgbd1mAFXHJf0f4R
St8J+TB1Ix4U2gNz2Cz4LRsZJjRccL4+Wxrdmen9yZ+uhhYf5hTNZNT4C9NHXDnp
F1hFGefKyLtSts0a6qBFqnlxSe+Pc8UW6On74yOLXO+nwoAdBPqxabK4Kud7ExNS
uO99rg/3xT0kRUC5/evLqeB5vHm9bO5tj/6D0isESwB9yNusffoO+008l4P5ueYB
uCyrxiA9mvrvWIQ1tGb0rp6B42MfMOhbpIyYdJYB/91iG2XVCAAAQ7N3R96iU7lk
X/tEG4b3LSUOS2REBMkCL0KEf9UVw3ohG7Dwz27pS+MJqZBi0P56S5sdItIoeyNF
ZIfxA6Z10Vl9uwBIaoHGUBjq8VPPzE+hW/nY9h44rM/iEl6KxYzh5ohFEakiLjR2
RJKJx4xBTU3tD2F00YttXW0uXoGQ0BWYvOT7HDFYEet2cNqa0SBXj1ZdkVBG6BMS
aI9PSwZyfPHhfrKFgsyAKw1yeCgB+wEVKJbNBdvCE1b7hk5GUa0kyj4GF06Pj6Oa
FZO5I8Jr2nmn9nmD0KDKnIVgReVhoAjYUz+xziZE7XSLSrwI4SSp6qr7F9nU4tGq
kHPNE74RL8YOInwbLz67zLkOREQKpt6SpYsLJdA/zrryWZbCvqy9OA9F7UJN3ibF
zXwP0dKb2ugVJLIM5xR5gNCLfKzpRp+vvTcumnqEaBIGhtvUfAJMIY1I9WdzqHnA
321Ovt5sIyAOTQcUEtrxYsuAplHDuLt1uBv9RkvPaphLHUUwhq3DAf4T4670ilQK
u5p7F1Rb74usau9rCPKe4/89oTp1xScP7osYXjNxBo2twa3s2AgDktpTX0ynt9W7
o7wVySr4BcS9uKTf/MEm3beVjoByuETBghWjcMWtxJ7xL31paGM39g1kCIFfdHiZ
nAvWKto5gZ+Rk88G994bURwG5mTH4Zs1LHXdDHfiqT86cce+PixGgsbwOF4icwh0
HKq/OE4GBHMF96Tz/icnAM32yn1gkgcRk1LganxtYkQHA+38JuLNhbqH+OmKOb/W
ds/8IcdcjNgqFittdLpSPSK1vq/XwNJZKienELiLJypipGDnazT/4bzQWPLbH00G
a0zqpW/YLlGo011rUsr5WPRu1SrOhyqGdpxaaOqLNVsiH3nZRJ9bt6g17jbdORZB
txlj6mILeKAxrbMlN0P7S2OKFRmCqrMbOKBtDz2H3IhmOvYd1uezPq40IMQkTgWo
NTWnelZ6JC6izHR6CqMR9uFS/PciJco2nH2rPMc+TPhAB8LICUCwjiDI9T5jCutt
mrN2gayw7z++zw2O/AbEurEO+VHm1IHMsrYhtYchXtBnPTMM+HMP78dAjuv3yuGd
jh5krv3c9oJeMlhVM3iMFb8AOcmPnsvFhMd05+VSqED6I2B+s4HQHeA70HqTff9u
3v7qj+ze/oxKx1Oiesz1KJgYdx3n0G2eudejdF9mQ4qNS7Jdh9LkZLHUssuwAR80
YymnPXMOVN8WfecFcIYxcw+t0qNCl9Y87dmXoiBgFEuPwJ+z+Ix8MmFgyn0QRpWm
JC1x4OLuEZlilFjI2XO/qvbCfWbJTxqppQb0W4fmTBL8WKXRwV0cO4aAda8zmMTl
gzvNxkEtGqzyNrXIfcbKCX1oLCm8dyS4D3kydrSiWLVNe8MciU6Ko3kigXWNyyyD
4LLwLR9SH1u1N5Yohe3fTg2zAUnNR2pspMc7UxdWZLkLSqVfEeVUgsNV4xJxSeZf
ddiG0/n1seimFZTw+41FsQrHEnGjuZ6SDrWdNGm5KCnruVaz6rvNIjI9p897lYqx
NIKkndqn+71R1ZyXaFjrtnVKAHkfZBosCIrwI9Af+McLDdRZUdx34HHuJ6xJm+YQ
JIGn4ySFRBRfrlWnKCfojvsLxin81oN71euAsLm611fP/DOQr1z51doaGrFZbDZt
0TDqt8UTB8fesi+zHesALNCsLrStZz0Qm0I/pW3kEnxIM0owk4+VsotGmWfeNShs
dn8ngsftrNZs+W/ks9kJDoFHckNO2W4vh16ie/rOPKmWr5DymVsspjSqb0eaXITR
omnpKNhNe7epZoQNjcko5/segEJHVC/GDhAYxXJwiclswtX1pZmjm4bdQAelycJj
9BGZDAHSlYnM+FHJgXy8AovMMvMvok0lYtuhkIe8vFQlkYoZrgNZAKzhKLlQmWlB
KhvXgm6LnuE75RbGe/NhMqmLmg6rEX/jg37q5BJJvT0wMXWCq6dchNykW7ZVP7IY
ztznrhgdUVTddMkYCXuM0Jy+zKxjnXC+CRkXaNvwcDShQdLQmzRyMbmJYVhArdit
aOHeqGi7sLP2h3boQKjMko8/09qxBVXDZueeMUaYQwMQZYPc2uyPh6T4Xqkv0X1m
CegsH3FBvHXxmWEmrwsT4rdGMM+bC8HC5s7mmIeDYOCHf9kvCJQbNpKgG+1nhTrS
Ju+GmVNeKjpPBy7dTVnYUEDy3r/R022NCzV4qwoojoB78OyHzU/rzA/Z3V9dXOHl
8V8273oxkYEWwGs1ZEmhShx8Ah73v6FkdaZgldNDWU+pCZDOGGlvuP5TY83tW5iJ
LkUMUiOq14tT68gIfayQWdrhGO5e9WGfmCY+bmadPJak3RYduMmTB+zC9xAOOcCD
PWWYhiTB1gsA0uRgVzkK3PqD1LYweRZ4SYfZdMoJsWEfdw22M96m3gDAbjxfWsqE
C4gEmQ9XPt0JH5TmduU6TUey7GFtyDTCDd1XSdetp1HODJJaRlz15TZKcTxYnXUz
PX3S9wDrjx7tPWnASsZ2EQ+vwg5cbTygLPC+y/2t4pIaG16JmYgUIi+oYfR6umL4
5FmA5aSiteqKohiiN1ktxa8DncOi3LgUIU/EnQnsaN/mH9N4l55pP3UREbkAZPov
ZM9DHNuASs36tMhnOBGon4djpzqaEs3aDz2jr9ZnsxfQ9EYmpDpT0ziMolBdOvLW
BDw7MXgrTaGo78rj0ARw/lm/TPLYLw6n7pZ8bAPCFHUKMGUNIK2DS1MaE7RgbGz7
lNTI+o/RbQ7DidX0DNqLA82HXhDTVDdoTeqE/x3G02uLpD89NRyFxjGv36/Bksmi
Gu6vZZBIOPRDSNO/BBn9hwdriW3m1uhw4ayIF5W7/1x4U8uU5a79AUKgjR1hkNws
cY+bt1wmjMFsJaP20KaUIqCB8NzCoRZgQLs/rifslDBiPDGRR1VrPTQhxFuRYgWK
qnDRhLETxgMVSMoiUxE6ZQW80JNDNFnq3Nz29gNhWX7HhqFOOWdio/NEdHtBQZ3b
w4ZHCy045guJ4qar7EUGiRdi4GzN9eO3Cf0flFLkFpXKgKTEH2MMHVNVmqdahSRl
AtTWXAzhLCA0z61p0eJF6mGz8ezdJ+ehB3o54PUJFNQgljJ4/+m0SyXoSG/guXwn
0jhz8oaL8D1Mf5GyzbwrPk91cOtLBu0Xlxfq9bpIpilhvHnL89DGPG+df+e/Yjxq
x017wX0FGfBW73FuSGIqXyeW7fs+YqLheDNWE8Oa1VVUMNdW/WHCyG9nnNsycbtT
72Kw3X8kecSK999XqbzqUaTY9Ui/jTjIRPnGyQXKM2sUx37lSL/wojpfMEZXmSlj
8Dr/uclprTiOg47VRBkPivvPENhzG7/1L7B3G5WKvi4jZIgt4G2TI1YteVXer7Rd
85Gvo5FmOLrbjv/pAHUiN2iPNTJ0a2Tb967jzsAqreZyKh1ljP2SMvDA3HVpufRN
js6vYt1XbNkQWRsAsAvLdFV0oj11XqofA+cZc84B7EL1DEZuvw9kXflQ37VVSM+g
Ufx9d+TibzNJqjDFvLbdqAi9RMkKe8B3hCUhas4vWB6iAwuvgb45Xr+l7LLrAyLR
bJw2G9L43/zuEWUM22EE3iEp853RRNMBxuK6tkvBlxyl6vG/VmoiiC1Tp+C8G26B
xPjxYBPHnJE+BzxOLPIzwy43E8bbWciAdJSTY9tot8aD4MZXBxOWuiU8EvUX34hU
Vd9iwA82KMwM4EcpfqqUzBQen8TlCJ5N4Om6DHg30CAqa8e2j2g8ZFhSy1UHp8Zp
SRWxW1UPT+DqoaGPbMHECI/Yfn5q0tnjZ7luEND88RF4VhF27F5XaNlBjeVFaVHd
sr5SBA+zP2f9yWvs9hak44Q8Q4zjqbYa0SjQpXi0rpc+5hZH+D2PNW7rxef/ebiE
UzBRH8OWTzEDoF/A49bBgDrBErnT/QaSlOkXDDqQgRMb0X4GRmiulY4ecyQPEdTO
LX3DpZt0Smu6WHXqRhN93dq336lzUmnxAhMB4jwzrJ/zud2IUAuzw3J3ybIabA/+
55zheoRzdkPrcX5R79ilyDYrTFGiGvxsm1SS4c+vR+GcRy7nmB1BaKKGs+joaEhX
OxyJtczG7scWquvxQ1CHhGI/WkMC5TMrNisUigQbfSmm1yRq5npGm938YxN1slDM
43s34VzLwj2nOCxPcYfd6enQhZYwGCQif94nbhk+9bu/nP9V9M6QHJ5keDXU57E3
tOFp5KngfvGvQT2HNIUuu64r7bmWfxhusu6XXeLhKvdwq5ax3mDJ4l9cQTLciS9C
Q68/UjM8Ib6+F2sO3qg+7O4cAudRSFoKpct1HfKEdqu17XAuvwdoAPlv5D03zY0z
SNp6otwKiaWaIlAfEDUuEZ3tf5WLT9q08nCM7vhVEkTDdB21rHr2AzWTSffS+28/
EnaJq/OI5wRX9VsO7Xk7HSBPK+Nh/PkApCypiqouXCta3I2SrhkDQIDmG2hjyQyK
zcNEYC9j8vHHfEvVdDF5jkvn1BAVvuLTmJCPZSSpIn3+5b45tkb6qiZkF2ddGoRa
125frBgO/KGtZUDAcQx5gowyDMoNXTuFS3WAcFZiKQV4IoIRJLG2Cst2xz9Qnya3
2k4zF6JHFNcz/Wrb4LQa7seDtszH5R0fO7Rfj1JC6VxzJR7tIFy/X9udkRNIE9L7
yKgtPbhxA6jPtVtkB/8p6/R2Wx/ptO5HKHBxo0OYHZqfq4xPgYlYcHq0uWO7+3zW
nL5jvOlYVQY1ZAUk23QuAceGwVUOTXf3YLkTymaW9n2UmFhRL+8ptYnbJ6beEgZS
Cia8x2lngG5PKAbXUzmYo0rYHB02riwK12pxJ2O83LKKQMDmIuynxLkYXGPFk8eC
tASjhp8AYxj5jSoIpgd5pVpKnb7bAMdbqOwlUYwqOKQH/HFsiJtHlGnTb+u0pZqQ
iyjjY2QPJVz1/ycZ8QvEk8+dKoe32ziIvDlFlcmxfcGMo31TRIn2uBRkGja5vGGh
W8p/gI3c2ahFWMMlJk7HEGQKskK8TBsFKz2kMf3aQWxpYm5TJ3W9kIZAtfDbIDnv
i2ayVAUwLME3015NGdY1WxqrrS264dUzSkqHOv9m+3CWiWs4GleGwu/Apkgz+WZV
ybidbcZxnFC6fXPeYdhOzSfdTpoCIrx729STi6ZI0T3sw9MYiodbq9iy+pISw4Th
RJBiUlmRqOPUnbcD/f7NGTH0FCIjHm9P9IvjkhYb1SfWX6FG/FXmBD3lsjJXC0CH
CmyAxg14P6+z+9FQxLcYllMWNdpUsdTQFiyzreo0qRpeGBkw1/kOQql1e0xHhmJD
QKjzTXahl5v2IyZf9MwEt/NYLFmUz4CCrEnavYHntjDge0BAJQibAC0g7jbHQjm/
8qBM6Uc7O1+Sk3PD0DBsYPJySBFKbLMqQEBN9I9ASG4oH6F5m5wZohrWfy8px2QI
A2g6Rs9T7Vf0/xnqD0aohculWY5Tb+lWDKv4dxnvhOd6v82VY4aiNSwVT4p9LmGn
8cuTgGdXi/oBBJM+Zu7G/kL6sMEcam69WLA0xjOCfNCAUg0VmBIInTJ0HcBFxVQl
1q+yCAjr9n2sb0d1sO8lMLkb42UNZFOjukUglje0Kc86StCrRa/VZz19iG4J6SKA
zzUiHkZjObu1yNLlXYnGj33YewGfx9uvsntAi2MIapkorI2MAnj1Ko8sOAemg3K/
nzjMuEmcM43HuPspvXx9TSfJmYwLjJ1K+qFAhUbtARgXEwWltoIoUoV7qaxlCxcY
ImRqAVojQxfjAxpHVxjYgmWUsMksHvkT1bxuxxYursMol3Cz5G56v9C1CyYPuxye
T8b6wPJ3+cW6EF4JDF8FaPrVHdIuadnvqF1TRoGLo9AllPhWhIQdD/ihP4JaIglv
mrxekiqm/SQlvheGY0q8gpoopzN3mLvVtH7lm/iNup30/aDWll3N5NAcH37G4hXw
GfJllEYapw1O1dUD6w2lEzKSo3tJ62K2h3NSFYV/Piht6NcnVCJsXe9S0bHuP3W3
L8Wy69GT1QuHWX7r5mku8fE2pm2t72GcjuJpQYL1rLBunr1WTdGl/HP9AmLOy/Z9
1y4BYy66mL/kCvBnhpgCTrL71EO8l3WAlAL6M3ZbCTW42qcbgKXx7xkzfkNPs2Pp
3nAg9q/+PXJcl9hu13qvGQdJXp7jQ0iENcm1YoFenQMnFu315hKspw8M7DTg+NO/
e7mifkGCGxI1+wfhuoAk7LZdXu+Ho5/lKqh0w7QUe5/v0I40LgMrlUw67H4MHOJv
JICdqVjZFC5TeFP0taKIsPJnvuiFdh9jWM7/qLIJGFRhEKavBaq4Y66KOfOrhfSP
tEhCwqp0/PXiKchUN0u6qTemIdHCVMZ7U5+OCDcraJRnfxhjf/nHkvjwGdZOadBt
4jQC528sRE45iFO7LKvau6A1/Knb5Opp9SUfaxE3RoQsrsaHaRQZ9bHUn86C0DQp
MxvZqkteaArFMCKt/IiJ016pqbfhQHPUk9lcblibgnBPh5ifVMkwyaDpl7Qqr+tn
jocITnZejnB2zEDxrgNINvXUEKgCbQkHldsr0nQUQ4QjSchMKz74lmpA2422lU21
C6mTWGJEid/BqZyyivPNuwphyCuekfnmtZqEqLgxhsXAtIC7gbwCkIcqxPNryCbK
h8PTaaegvaC3uKU0ABNsu2S5HbK2lvTHKQT7UGxxCGmMTGV+CJ+wuGWIdB3GrNXU
K9gDerI9zPFAFr1/B0wPmT0H7zn5tha4QWj3afAo7rDmirOml06KzWy4Oo80Kkl6
Zu3LMGVvqEKT2Jk3HX9cPT4JBDyYK//+SPtLrnCOpgDAJy5uDtwo0Y1xaV2B2xcH
jTUBnKqeJifuOLovRMOsfyx6gncCe2yOLt2vTjzXQHLljc6hgDgcbA0YNGTRCbnK
+0u9xisfSS/8cMG7SUxY7sFxTIVFnzNfkYwKWZZmbCFN2QExnq94fka561bOikFc
80uBkywEAKcYL1WrGQ0BJDDmOZBq61jvGrTU9LdkCszXhTkBHlAVvjGthRXKhEeW
2sIrXGyXN0m5rrLAzDVupkY8BBD0YHKJefgCD1+sUNHVoJIXfGY6yb5eT7pIHCKm
moIgBfEF2L46B85SP/KZlkfWaJu5JZiXuRBvR18ca1FvX30TxVHfKNQE1FOzxzug
DEOTUUsz05yqCAQBAdHOeMl+U6VgGLViJLTORJE7FO3/KzD4kKm9T6pICQqOUNwr
tRk90mIi9BEsqpinNyceSwjM06TP2rTe0aqkoaZ5ptK1qD9Edl9oFNh60Le4odUU
IAe8Aw6bQ3sSKxH8xv8wB+pBc9Nd8vOKZ9Dx6WANJo14egT/YNuxXcrLVCz5mvtu
sF+b1l7X4DCh/RM60zQl3s7OV0KlSH5G5/327DmUoh6cdRScwGwk5QKzkX7LXTGh
I2VBxzA28YDTErniB91Nq9v0/AclyFm2AdQGc1MWQIC51seu7Pg8v5VJydkmks+4
7e2zSGWagS8dbpH+3GOlbhOWjkBeNyHB9Jz1FuelzkfGLE9yYM7f0Qq2tpmG1HpH
0YVdZjLFJ96j1n6fGD+JNXzL9y5bBVZlVsVRYYmA0ci7orjfWAt4w37Mn7mlCipP
HzGfXWtnv7HKJfJVx4i0a1c5w+JN/zMK8iv+q+nIXc+IzmhcKPII/BwWyBWFbpyP
ZT7Td2zM+DBa4wGcd7qtBZsosxAQ65F+wphRDuEAQuYlj5b9fBHbeWs2YYPy4K8C
q/UaN4wamY5xJjez4pBOLoTSawnzmWh7TWMGHVrlJJ9D9K56yz1OpTYyPGLhNHDI
CB7lHuOLxgl4EvE6zvQlcUwF8OVY2/n+653ObR3hLaTkernKcmM6yoaXGCVOFgsH
apGojoZL9zJKVAu3yPqAvyMpTnUKfwbwZjTVmvKYBzfHGMnlaH6jCh6RfogRCVut
RkCfEIrQt71MJkhcFwZFV99IoQOBwwlQJElIH6YQsoMzegvvdXTMZUIDwXHGALkG
2eUw0l7bRabTltZsp7kES5Xk2zDHhJGHalRCrsF19atOBx2RZtgxarx5q6nF1h9K
l3LeETU/yTB23ByiAbcryybQLYrLVLvbULkIF3Xe2b5Gwrom+QyHHEi4Ajb/vTyB
zLc349tQeuGZ6ZrndBUT1ng2DdOL5Wgjz3N5j8Uy4UEBY18SPaTI943vEMLXGFy8
/Yw4er3fqqpuGD5GclDpHgfNVda2ObYgQILIDVKGoVlZ8ltkXlHv7fZFB518QllX
87/gTFXcsCIkISQrpBFiY80Y2+s3hBYQUqT8Jd1bN/fIUiNMQDR0UeCEm1xxxS/R
bwIiyAiV9GewT8kDTwOhoHe1EzYBRzB6rTrCPvSt8tus3h4P6h9cd3c5NGW8LC1c
dj6EuZTnxi8lews+FVz93ajHSnhH+nKsxK5P9bjvgR9h/YnR++TielxYiWdPA6hj
Tj0+QhU6YUk8ExlogGriO1+GN05mjrmD98IRvn/3s7XqQ1R0bl1AS6YUK/X1MBdl
UYUrvg/V8Zmw2+B5gltGkKHmjF0sRe2fqSwxIi0hG+RMf4Y6KXX2A5GywDk45kgK
ZEzMy/UpMNHwESZXdickGksh2+jLSirmX/NZvDhjrdvgMtk3C3gb1NUXPqSaDKQy
Ge6FvM8+X6BvOOgm5PMDkIKIbWw5xmd66IM0poL9VZnGUnhnWsSnuWEH9N55h12k
GgOc2NgIRHDCm3BH5BWojnpDf2/rVhRJX38VqXq1s3Ge6kEPgSocQczQFWtRg+lK
+VhAc4VhnSslKMxLL4Jw3tmckQfGjRzpaEfs5965p9MBFABDq0JVPsIwoqCLwv9G
yg/nLdIVXbo2lrzEcjxw58FpmXL0j7WVUb5SbqR+c8AU9Nr4CCNaN4ejnCf0xKKu
du3512O3QnYD2XnsZzfXtjfnzKKiGl3bv4xt8F2KGxsD8/3Gd2ZyNZhEIIp+3V3y
bZN6dON7pKh/zd3ny9uvB8TQql2KBa84nt5Y0rzA5/j0nmozmmSqrPj4FqxlMNPj
Wqr9U7wNod6/NfdtxEWXBz+KvT//ZUuLAB3gpfVty/DwemGJ/9j0g10esdc7fskK
0cwKy0p+WejdmoED5SLbXhTav7+/Pao4RFzMZ/4HY5y88GeQ4g5UMeDJyeeg/z4u
fFbu/YOpA6vl1mmnf55NOJhOLDT6oWqAw99tcp/ny5JbWGmyptQePU6S8groiwyo
kaa2O7iz0GSX93JUTGEBkN6i8Daij9i8eU/LVkl1hx8KBoFCNCpXW28VbM/4t16D
7D5jpHmNXIFQIeB1UFi+ODMv0JcPH9hrlBCtc8o7R2Jjd+9r/+5NKRCLbidXNyvh
Xj7cXDnUpCC4xYO7FKR++i+DGABtX66PrgEUM9lUc6mqvjZm4yLT5/7KBgqgNHLd
5N9p90mr9wWzf6GsbuuAUZAdafjUuDjFYCubHEvpfAHpwrj2Rp0EcULxoBQw4O1+
Dp+sBfssImgIHhnFDyg1k8Nh0QdY/JYmDiUapymymecrOEneGCB5h32YUZ++3PL1
W0rp6rdeHMSqNys561tncuCboXjroRlFfT40rbMLLPQp1KaBzmefXvnCbtPhUvSS
ZuxZvpWQQI+dNYzCucheddMQtGGx7KDVInmrCr65k8RWTFswaZg78jSF5w9gAxbw
HMNoZPjhQ5gYTVDNOybWUWYSyDFhdPdxa67ZZMwz+xVONfZhvTADC9Dm1jdMc88g
2VK3UuKAsX3vsXSaUp2nLR+v4ULbaAnVYc3jOrGPE+kw1Rt7KVv/b4g0to+9ghUq
3vwONeq4UwTdWc+Ip/umV9NlcBakZhoPFWSTqTkxaBsdCg+Corrs6e/qHqXECM1B
9Sg0IlKAbuFQi4Liad63bCbnBfRNLSOoZcjM+elDcLwZiFN7mpzIERezTVAm2LCj
MQPtoDiLZWEi6p6hEMWv///7dOimTjczEb84JTcEJOv3C/J3iwbBbOQ1RLhcZH5m
VrKzil4CHreFLP5zNf39p85Z/m6EVFPCBdHs/cDSvaBHYU3eX3i/RNAJK+MZLknd
JKbbNyRBlGJ4ysSia42Pup7ptYUIdJjQCTFRlAhz1cmUVI+/whSwEv3DGeTupZMA
iswlPYBccHNGrBV1ll328wL77P1uyvDXr+uMoaBfzGkGDSGSYftMTgc/sBFRtFlQ
GLOPvtYB4i5JOK/OdiRsvyHPBVsIxXbb4nQIznHraNkqCSA256mSFccWmyRNvNhN
Z6JTsiAVBEGuFvv/CQMSLKoKy3cn1X7TEH7DZoqocSGQGXod4c296X+h2X27nxuL
BYLuensWIsgPeocmv5VQQ0OvQPAhl7u4xTWvh3jHnZbQireheZpd1NOWkEcBl07L
cu1ympUThU0J+rLI7NYFl3Wp87u2N125V2ZCOuV8+OXZztth2P5nwEGvCTYb+uK6
UvD3okTa/FnriYenQxGMDIkQ9Krg8pDt4jzhWtKRcQYXsCfEJXS7zu21Vybcq9GX
pdsLxz/Blh/I6eI/r6maKxuqp06GocU2xsEfLQx/Tccs5k8DsM8AYBCyUni1NysF
pEF7TdEKQR+oM3387Qw9sOfB2Co+3T8Bl+lxguxIKnY3Kkz3q4kvSK2j6wXSz4BO
i6suqogWrHmIPGNGTCwbBP05g24OB2rbPe1AGIWaKPRCOSdagFvLN56vMCLQZZpW
vOjfUCp4c+1r5jH+WLkxowiu0NktIE9kX84Ot9L+IgCr7lL2J6auoyUHv5etD3Md
XKZOgfVOu8zmQjSQMWSBylwEu9PQWARxmklFkkCfJ+Nm9vKoXbfuy94IqoYvqy08
MdVekCe1sxKAjHVHKDvcaxlyq5pxDPS8ifTKkuPOdAREaf0Vkj+9+Ec0DJOdwMeK
HGAPHG6l+KS2bhes2Z+xOgkMCS5JXagICLUW5qDlf0tn3/L3+few5TtnI/vW0FA4
XbRLuuzCnrWwGjzHoSNvSGRO/SVjVOReiYSkDQLl4CSeWrCpZ+gsaoBvGERodace
vc82E9Dm6Y1aEBibenp5Tut5c+CB3hf9UC+Tswh9eTH1lOvBJJ/ogVwKgasL2Bnk
tMS0m5pN/o2YTeFHiI3e5JaJq9jj83IhhHo1u6oM70euWCmWiFHuSJY/luEhynZM
ksXv7vu+JL5pCDr/mtiwo759iah4n/+GX0g6LO4hWFBt4y7uTIRNUMtDVc69JF24
0bjo9pMOLdwtwHKEf7RSDQpvDSXYhTPlR8FxGIe7nTbSRFrvOfqeqmKFGFCvoSaF
77/V+u//uQqc7ZqLoYV0BlYXYg40+fbC1/5sWe9deQP459lXdDji/eKDKVEHWjqN
ddYUzCUc5r1xfXl992M3S9ORBks7Y42qr4RXo1BZx1ssOUMd8BNpkjA27m90XLs6
/wJm0+I13//3eaewmqvZjFfq3lEkLPLzwXKCl6NtjHQITjHwSfdtZqdMUQxMdJQN
QvwNXXhAgIU5BycGg7e0C/h+nkfv95k+E6ZopFHIJ7pncaz0KWslXyMKqmfULd0R
S/2o8XOyipYzALCVq8hliqoPfpfhGnfQRZweIxczYcmA8D/8VK1eO6pQa8ipk0OJ
e4GHZezZnlATeE5JSVTSUJ7vV9rI0aeI5rQI7hB0nuJjRgFDES2aOFoTE42eOXca
RdlNg7DAyi6U2+vJNSTZwIE+TrH/ubrExwIFPi6iEZCfTNgcebBh0kUe8IQSPZDA
yvnw2cJEpfmhdr1pNcJBQ1hmYkJeO/i49dARLgGp7Oo7dt9cditiPRVDIGziTCB/
Twn1acXQseqinUcA/mIzx/9WzcnV4LXWMRsFvThNYLa/jvx9CcFM2xyFDp9Vkb4u
Uixvc3huyevMY3JG1oC41c9qLNpcu2DHjEVsISACZOBuj+R52h1bSIc/NRRJnNvl
7LMqFH+1+uRHn276/rlYitfX+rwCrdtf44gl7PMCoYilsFKrNY2N+GuO+kY7Rt32
EwDjOdgpP0feBnWce73cCXkz4bRX5Dqt3spNo2cGJGxaqtQfvGIYTzUYoMcMe/zU
gz4tlGWXNwRAIaVqfhXUdO+OQsc8/Xjb9x8ownQ2SEB4DV0dOiAcSMFTyQF5nC8V
aGD9Saj4rVp+OBFh+4mE3qaMvzzQjHwXWFa+90t3KlHCwFPHWrGRNBHdRTaSOP8P
6BE9OQstyHw41i1XIoXl116NGP0L61GQ8CPspfjTz4UdX45NHZjJBNWEbGzyLKLC
AtpdrMhS13bJXm5/2/ZONyQk5IdmZiNKmGCZXfjf0ahTBsTW82HedxCi/tmqYw5P
ZIrazalGp6IOoW9jGrKTxzd8krn9Uz3h+2dLDSsDtV6xIsdPTZYB6nbkmuddIgoT
r4pd4Vd1bmgzcQ7hN4BFPRUaH3Khtxi13vzpKOeWs4RbC4xuSdcoKZrJ292m5PHb
T/OJbGaQ8KxQt0hk1/9pyvPW+3nXOQ+4okPa42IBSCNRdY5ta/LRR0CQQmIfvIYh
eT3aJGLVBG8YUKTRGYDOAeK/S7/ImNqDNn60WTa0KiLPjCz1fVT1lV45RPYVeUm9
pDda6WbWvSQ5+nHRECKlPKU+4a6u4CXvT174ydcA+2xT6T2OORDDQK2YS4EkEPOA
dOTZR+qQKnmP+0pVm9lF8fJ0UOX9yqvHJh31mg1i35gfbi2AIA094iPu8FvtLClq
8hFqd0wIZgwVYjOANd9rJUI9jdwW3Cy1P1WwV04PbYF4O3tHW8HZDXYUoWV9GQE+
Ur8OATIujKZAAajyzRuMHcjngthp4PUz1l0/wNd+50WyYKslEJVaDSFZW1Xg2zMR
0pFDgfVTkHB3fmejU8VhSF4C4b7kZCQlx2/0wk+IwiVFrztuw0Yt9qFWSGOY6Fow
+Z+Q20Hk/CQzf3S+x90XfFqV8RqiRh9tNy422eWHUvbrWKI8TA4YnAAH+WTIfJN1
fLOstxmWPPHnmyz4+TNjxOCzuZzPtM/fa9C6LpU3EOxdz8AEAa87RlKztH4Orscc
Ry0IFEUF7aOnaoYzdZQ5oEwVmJpVbpb6ZkTPnQWH89P/LpD3wI/WgH3n8E+G66i9
g2AT1G3oI2qfrEzDDyEa/YsxLXsqbPFmlWm0pKE9P6AjKXL1z3YzW6n4tzha2Z3I
ZjgGmgNXgC7raqa3PJW+3QH/Wxp2VpNxdq1cl0g231zhv3nWiQHAQ2eiRcHgLhzB
CAEI0J8KKAtzbk4LTha3darR2rPxMzx3a6bzwsa2elHViEV6JsuoosbULdx4lZ1h
G8rKoIh0ra7y94jrDxjVfjTPVQBSfBhCj3ARo21CRMB0B2e1mlsY6edYbENR8lm0
yy9JjirqrwOK5LZQcUjcNsHl/x2dSYpDL+8CPicmE5yy/89K5iQ+HO9N17DcEb1e
YWTYbMsc0TbJt4uK0nFaQGbUfqWi/e23DSSIKTx0iSVsJJu6pWPpe73Yk2o30hjr
NsoyvWYexkj2PUwkGS7O4cTOU9FndDhwWhIqwWADHhBlkHCok6X39tMMFtkT8SPZ
kDQaDJ3NFS9kI5jYwd3gECrlTNO1VG/Rs5omyuiIal3irIaWnBxZbFmp6pD0/SI4
iPOPs2jvkfh55MAGQ+7XJheqgmD+tO9DKRbkuTpnNzB45Rb5RMwihIfreYCxmVCA
Ak95Rjibeoo/e6tn+HpxV2PS6vmh006zJi2pheAUfEA4xiHl50/Ea9fe9+kFoLGu
/uzpJIk8awEUQAdTgp12xxwD7G39WbK79p5yWJqfxTiNgwy77Z9wo+yjZUzTKhdt
Yj+FVIRJHl9CUMrLZWlLTF7aIccH1AixFHYBUdp0jheq5Rdo+q+I2jyWmKctVyjG
iyEhygg0kLSXJcDWR/3Pz0JdpN/i5slNOVGr2uSUoFg3xcY5AkJmw+/PrBQDv9NV
nw5QMKvaMJgPAt0dc35I3I5tQT0Rg5rQJFlSs1Qoh0Sdvl8O/hNCb5b2ll9YTRFa
UhZMx2T+ZNavshq6LAxY8WpFzJ+oNnQsLZc8SfCmO+3XJ02nOFdyc5hYmW4C+U4A
TQdNqeNZC6cm+Nke/hIzeEhYAeAYGSY4zAdkg+27JameI9r3EyRaUJVdRrGVOqYn
cZTNEMs/grlQjhrD/Xv8+m92c9AAKzDX5ZqCDdelk6A0sMwzxtdSe4NHH1ULRW5v
myp1hIWBTKWNej2Rmx3OCJMV88IFEWOjK2R6f0vbiBfRHbI9jDGCLssJsz1WnEE/
+pF2nB/eHit9ogxyhwnPYXz5a+BsI/4wTDC7xyIBv4ZuRwvsK/TtCu20r/OaUQE0
9qa8Ax51lFJe6OeTvaMLVgVqQ88XUmpDYGXwHtbv+GPkfxNujDBzAfXy3mmfnMrF
ZbPqRJIhHinZyhChvG7ODsIBKCHfnIrC1sCy4qnsYk8NdPjj60XabPSHFHQZItaw
PNFYo3QC+VbqYtV1PlIiHQ46SR5Xafz2UMc7qHaMbmenoZ0mRGtHWrKgb+eQi3Ek
L6WApO/I1mK21jX94QBVjglBHCQoLMzLi4NWTq2C7MiCoLHCwmyPcCQ5cLfA1Tf6
sbjh8jSbvKVHPU435eCKWAo63z95bXg3kSLiR0AyMuGHpWm51dC5HSOWhODX4roE
tDInx4xf+J3RgVDCFCOu9Wbm8ceC8KWvtUxr4XQkSlXIAj6PjxFbLfaSsJ3McvQx
1iOhL4QNHjIaPYvLbZvDO2i5dl/2wTFHFemPOYhG6zLJ3TZamK/b77vWFhPaAFB9
4vhdHjN+2X/I4LDgBExw9vBVGoufpd9O3/q6XHJJ+RFjq1ag7Q5T7LjSprD057am
lBaqVvjbNPMGQeEDRR49lO9OjoQ7RFmszGR9JwfnSApOnX+baBoMpVrVYOhx5rdL
rTz6u19bQ+4Supw4rFsjR1Q+uHO5FB06qOtrZjPJ/fnDZhXGWxMMZkYYVgnQ/QT0
jZdIKgygTM6+NzXqwQbmke1zczrI6NepYBxzkEj5dVQsoYzjc5aoueftQUSn1ob5
iyuot1bQtZkrLz4pDIxVy9pInjD+Sd+7QlzMLnxJRMJZ56hd8rmWFwBHekxSBZmQ
r2I9YmRDuG6EkYg06clR0CxBtnSpsIO+Tz9VnqLEDbq9WabDJCB9fYVceqGn7u4M
D6RuHZhMY27jU6g7YydDHx6ccTOdKFGYPhXGoVyOxPokEGD2fh/ANJ4ntORqIJDQ
HWIXDzErRIr0noVpUAeRXxH9AcrgdzOVmLOQe/eAmHqi4IzLPBrcP3gZkcVkYTag
H5LYs05rSTHZP6FWIGwlgJ3+zarlcHbRxV1WdMbnHJ+LnKS9O2Te078f8a7HE4qq
3abiUGSniED21dnbVkBbWqIMCt8cGsaSdSn7WRmdKZ38A2MzqzlV86ar2wFGyiJb
wmGbMxhE6aQqP/cQsG/gAl/S2lXjELgjHaL3b/dhjuHeh86aW8idO1g4Qzej95de
rNnDyBR5hqMcLAyV7Prt8B76kfw6SeBtIoTZP2QQ2+0046UX6JE19gEDL7ItEMhh
DEjlDKt33oqM3U76XxoavY5haJz6HwOa0f565DLeAbNoJv4Jl1kILq3hGv0bBuB6
Pn9ceNdUrxFLA/0k6dqIUB3wthisDB7zaDdKaLjngWZtWp3mXSHO1xLFNveUAG6h
kCyt9+6SM8KpKDqT8U7m4RJF17NyCNI2kFPa9UR6uMlgNtH4aw27qFM7M4hx3mtS
X9SicvDRdEyXvU+xVm8kGH5sgCQQOWumFg8AaeD1BQKAvug/zV3JIdfVn9StNuAF
s4pTB0ErhnHV1byUn9e7PHABLe1srNps+nL5wjgksdgFa1tNbKVAzUdy04dqZTxl
SNL+i4sE/xDOQsh7UuKckjeUpX1WycApFWkVONcfe3oeQVfPWBFvpoSDInWx094+
8KIMfN73gTJYstox8SfS+B0MFdnDwA1xWSr8EY5QB20ulH1UGZAyJBHgDBrE3Hhz
l8zm/ZVykYscXIQApJhH5EFMZVAYVR8sXibZ2PcJ/5Bt1KtikN5m8Zt3hzIRdQj/
TLMVkLFTamLKccfnu1dE+mE/e4/yADo/F1TmwAVr94I9/iQQTbeiC8sqVogvtW0k
UGe0SvfQ6kxOadRJiFIhKnDEJzLb6TT74quYyW2lxwe9mANq2qHjL05DMKZKwpwP
4zc6GKvVdFf+DtIrxNdy9HSM8gJXfYRfV09ZwJwkXMwPWW2KMw8MjAusXCM9kTk3
v686EdywXiesEhQDW42RIxbT7DG0LDjmcDM5j7pJeS23sH9txidQYdBgCJVV9ODn
GPosI2EeRSB030Ire7qtjYjHT7/BA2hdpaxHFNfpbf6KnTsyycvkeSf39XBL0VCU
Ci6IO4sMcCGx1HGjrVP9lAlNcXetUWdQkc3juAOOHU8iMupuI04SYmVeY8FPvGDc
Mc/7H8CU4Md9yA8AwTV6FHK62wxb2fR7K7xd0PGDeOcdO7fAVvVRpJ9hSx752YlC
pP5pnkonrW6eVub0deyPBgelEapgPYGww3bIxl5VXabrn7/DHffQvfdbY2+1TmKw
mg6tczYfNFKksTwxuQUm4gRnKM8fyBpZa+tV5sXvQF1P/nVPuvA/TP+vQdHItcAP
J7BpTep8C89CFIRfEGTR4fqJCevGHYRuY7cKZpF2SHHAty2DznkORriBOlOCoUMN
gBLgo+XqtoVeGiVLowdzVml1+qJ9yAcrIi8cfpv4wSk79ahZugEijBEx6PRUXg8x
Tbfh2rtjTwXChaVsVFe3z8TfZyUTwy5ZvUMRnJBClt+QgBgvjfRNpCi3XocUqLsM
2vrAocoQXde6BJ6PU4hY8ACRWOGr8vFkjd1b5lZQDerDV8Qeh9InvmnhaVkRdCpI
wQRrufSyTq7Yen/bEhrrVKjH3RJu91MB8tmUFqcVt49ect4nhXrAGROCxC0E6cGi
bCMFDP+E4xr7KcgYSjb0deM1G5k0RAB4X/U/lJg9UlJXs/8TDLupRSnJiigqgcLG
C27zQeummDprLwRn4w4+WGX2MsNs6eEMzxjObKb6vVpC+d0YapqImzmiztiT8FeU
zWbM5Gr/sEdGwmzuY/Lmz8VjTKjuMxc4zPTxc79J3+X5taiFTbaxhRZ2Sac3dCiU
70RPwfi1f+/O+Niv0nn8bHQPvy6oo4u4Eg2MuCetax67VAb+ldfV3X8xFTcbtCin
psOIqCYYhg9f6dKuFQdRsGAYdqm1+4Y3VpQXQCSimYNVBGCnxa7xor4TNevyNa2B
gFhpUnfZOyyGT2uHzTk/9mY8cIyVeSsN0YtTuUDXE8YDBo2FATB+SZ1IvgKrTRYo
96PM+vHR870/rDLr3ZQEOlCKQWvkwh5DsFCI+opq4XW4eej21wtBjCfRSXTUwkrx
5e7JTNrBtUXoC/Y+SG+4cFWNOPCcFOoJeZZGfbYLg/iJU7xKtMq1N02x+OfNAVFY
h2+ZgqZ6VfMfFhEj08Lj6w3tQjpjIyNfwVjI68ODJqonTG8OcYP3tcAFkeu07kp/
cyl5m7LJq2ItVL48OBJDHK27EW6XeTKeLKwgB+fwvvB+s4FuYn3QXag5I4WXcSGy
EShh8pJuBwS3QZNrLyqmGrapwx2wZF3+iFQ/9KF7dbTLrn5Djg7BmomKyaf0u+1+
nH/PN6zZbhHnhirm38yLRei8JE4Q+gInPq3ImywNVBFJe5sR0iXUVRNTfRNxWoYt
s97exg+fCfoNfdN1M0Yb2+PH9BuKPe22Yvod6SOvQAcq1rbK2oXOkGecma6UckS0
TXHUaeABPDbrvMOAnPjG38Gvx1KSJuN2qqSCK6t5l1yBIRwqFZ0cfecVExjA8Umd
j2KgLJoeNojqe8rvdxtqKje+D9HTKbkIPLGYd4OhPOhsmFFPL1UCRmH6sUfz6gtm
6mgrgJeQ8kUZXoz7qRVFSUJ/T5OMY446c4tQZyGEZsxd7emFrvKjEp+tUV4sto0J
WJjjZfUZsAjj91R4XfXIBLGecu/Rh8knOafuOIpjLXexwlS24fq6SU4ZSdoFV+tm
5Q2etQGV9jlkSkRMPiwky+3Hk0g+i50TViGYhQWxFVjU5HHhug/PCGC280CXI2MQ
/rCI0VDJ0a5FRu6F0ZCl6WpqbN+vXsTZzyL1znvA7RHW5yTOlTxdEZkYliXMs1Xn
aULY9OBofZJiFNnCEcA3Qt48LcyTWBrNU8zBi01ZcAccZfu0l1S4M4KqzBjNPZ7Z
mcFCZaRnHpFfBKJpA0+aYJOSWkh281e88dvULd92qL/bXbzcDV/Hcq2zOA+dpt9e
Gd5oV1FwarmQISGDMmxn+ZzVVcYlJFZilgLE7T6bGcclcCesb4ostiXnrW6hLgbj
bUI/IA/OidJ6USVqtBTaFTf/ieUH1nGQqIrpQknOUkXh/11vyxpD2pi3j2qaqDPa
djmVuKKg/m7O1qYm55In6L5QW6JleFERZUlnWmclQ0rrPa4C9VXHe6Ajif0k+MOM
9XY/a5NSjBakCqNcpk2x0IklWrh+D60jUbb32cdXjEeD9y0YzXpOAC7WIGcoxry9
IJiCISjRWc2xXS4UFGc6WifS2vUz6SuQ8zOr3m/lFiL3HiavuDPAI87vdAmCus6r
Qf1Xx+SoZ5JheIxKT/wG6mxo+smvRZIZajDi+3W0U1bES1SBLHVbyHSYE6plTDFr
oZwp6WyQ+TO63AtoZC2tDVeqV2lt/rPIWNfDUbLFzYJf+cSjnwC5GejwEHiFI2xs
jHlaMOu0TDFOJXcs7KZdtk4wlU/nsfogNDAVSRTGbcSfhry9vvqgTmNFXQFhnO9u
AnAa4k9qiwoQyHPwJdl8qiHDCjo36CSPeqWkBggUXXkJngQ1wentMbxtng/JRqB4
ua0T5BWT80zzgMYt/ELIx08//Ih/K5uFrMWfC32POnLyfQLQ1AnWJABnE41PEicy
rAZHyBwhUnDI1orNE7IQWX/ZHxnENluVRgVsTeqzhAMQZw3A2TtYfKHCwwNktjm+
4uPNoacb5XjCiWhD7LLv+tXahtCNTBEEQFkh45j/f+aMwXslJu4JuQ4cLI9fpD6S
4gzGDMQocGA0gspjeBNVPlT6m/kNahD/Vsm8Z5XwWSpnnSwlELnBTwUdbbNxmSkU
dpGeEmbX+Yg2gMUw1DwcLgtquK3FvFvMcF3PHWG6pTj2jraeEucR2drb3UMxNbQw
cFvRAjbyWojSnfJZTGIsYDeMhONi7YkmhBhZtBALFhkA6TMJcw8uWaPdwnXbFLZr
x82xCtVOAhAPHSkqxZxudxg1Sh+Pl2Z1QlqsHOFw+4ldZ1yzJ4mTPj8DqdLMKUj1
jYJScQeKCPoDVlPGNYF7dXIrdld0YE8KrKwXNqEbE38gRNQXphTfhHOy0z/v9cRJ
+M+ryHYdY3ZIT66fX4aWfYO2Kuu10Rq3uV0Z6KGLqDZerSUOAlUMwhpIHkh02dU0
VzOwDpaM8dUR4dl9faXkoxKCaIVklWaCjPDDOoFNsrz/qMkg2IhHwBL+gjhpeRWc
jO2LJQpdI+sLkuzzvK+FT5pAuon3q9ML43x/8PA15105yQqRiqTKz6IWdoiUAiRG
O3PZe4RljmBugsrLfAijqdvxe/lX0QUk0uWq8jIydp2eQsP9F6SOe1N6fq3ZJRyY
0kh/v/kAAEpHiykYPq8dQYfhb0nyS7QsdFEHt6zmcjz9GfTx2msSqg51a2IIvfC9
T5T8+fmtNMC/OKysUb/OHUNb9rom2sgc3djQV7kQRHCj/H43HKNOJHF/DUnXyB+l
UktRONtJ/QhY9k0t79JV7P6t8u57H7cqGykhU8BKF1cBErJyldU4WgWTVSQOrwxZ
bBGN/wD41ZGN1Mn9T6tJQPG5sg9BMf78+HBR5kBhwSOSe1by6N7xLNTn0pI+PNzi
36mc8pBrK68RtpTSObSJZ0NuWQzmRKvptm+9F70MutXbRhJGguutrFxkZ/IeuKte
0hPJbNKPDe1WODRyisCq9E8CflCwDxacmBSmGduGFH59XB0rHq0Q/7zh7+el/kf6
wLO+eAQkoWNYfY54fNzKEjEfJ1VogCM6/PTu94D/2QIIJrETIRQEviK2mpMjtmLX
HXCpyh643fB59WIWZeqAWdbtInVSysNyckPldCY7tBEzJci8em9VeD7WN/t7+Gik
plvsIjf/TRRt3sIROqtLV/x7v+rtSWv+zwdSv2Z8Q6BIv4/oB0svPzDB793kH3/C
sb6FsfWamoGYGi2UnHr3S3wYRPhxkfZuztFqo70Nj4AZ2TK7CCFRwMfzGqxzjNzK
tCa5ryvf3hlKpWIRIZ0yPSbe/n0CYB6Q8lP1clnJaXxk/quCbGZI36YRljLOXpLh
vjGER4300KJwrCs+gMly5uzTTM9hu1lZ8xYQJ712hXLV7PlLQ1hJ1iz1apk6uWJI
omsLO6zHWXUI5ZLYuaizcD1AlYr/I5v7cCtzSXw1gzFhdG9hTXfH1YfhsqxQZqP1
DXENkU7KTR8sPORtH5731vXOnJLDFFupJvEQhgFA0h0JXIBjp89R4Gqc0vFnpnH6
lv+cr8UULz2g4aPhZd0L5SLQ0pTpC7vRBcOu5CmcCvJT2tkt/ChR5Mto0iuyI2lM
Peswh5QHtFbIZdefTYDXCnbpfkEiMsMBKhOJyRzeTdUvzxVXZalnnMYpISOtFfyk
mtaNDoarpzQNXiIRyJ023u3CvU9YH192EAO9hqgaunekz3xvk0px28sAvzDZqACV
eBb0cqNERgawQBtapEvCAvvfjV9DW7Su7uKwYmE2pwAaC25F5fti3QZW2Gdj5X1y
fl2dMRGBGsEjxwbG4Em+ZyJLEapnHd0EeT7dnFa+ADx7sNsBsppIgQPozu/1A1BK
Wx7gTWj77YpksPd3h5klsyugQaMiWVqmaI5XoLLizlJndfhSyxixkvkP6ycV+lE9
VZIYVkuJ3Kl0g0lPQcNwtVTi0dtLCzAcA8sbQng7bK727Um7wgeWf/QMTWDMnTmM
pggfDBbvoEdDSwvzYetgVC4O2+qFTKtUaJqfIkc3dtgKFoTvlsyY/VBAo1H9G2Vd
1HPF91qLt/gTIrEkt7aUHbQyMOIoDJCakfvIIqa1oybLhi1FDasLigopUAUyEUMx
QwJFzF5YUwoWXQrXlOwbPTOO8JDZAhug+q37i3PGaju0Q0EBSzfL+klmCkqLsK+V
MfIjZ5/lOlhIR4ugaPPomv7NCJhCp9QKQERw4rW4GXgXXxTuRWjmcSV6m5dVbAIr
laIzT8JCqY31j6mpc86fIX/N8zvQrzU5ytDbHhXi/GmdmJpSx9dvypRZQMqJFWj9
Yl3V/ERC6StCMeMHRH86xo+0tjq7Pt3fVNGg0sWbTorBdR8unc2Bu0dNU+4+SwfY
bBEA8bIN0Tm6YQY11eA8bDXP/QPXAgfiCBTsIcokoOndy/iNK7zVW9LFYEOpd8c3
nPQHF5IyLHvluOxV0srZsCMwtU33u9BgfG6nsMjqyv54BLRMYILN7PB4PI13p1YQ
NCqmtjwDj5m+Dk/eI1J2cg5teWYmM5yhwwi7MxCButX0v66TMKpYhfTX7mnzr9ZK
JDtmNGbBDAKaFVMKfkaILrIwJD2EUD0Z4cWCmN3R8CZM+TKmRVj4hXTK4II3o2XI
Ed0TLCSsaYeUz6FrutbqmQ8UJ7hKM1aww1pH4HwVoMd6IcA8CIcZ7zMFUb7UzD87
KkO6MHbw440/+c/MSu7+aWu2K2CZikS+lfEnWe5QyIUqX13PBJhbyHUoz4N8c+yx
k3XNeIAhjjCJrFRpVV83Fp/jqjcylRX+/VemV7Fy3U/uUkTsIpbN5u/FETeTU6uG
UjJSiDRUhO9anC/idxPUv9GEYLGVtoUqbn73B8v2g8F9B5an83JY8wWdF/fCEKY1
GwsnXmGdDMCa6vZFl9JTp9EKULx6nOVJ069mfs27vWtoj9+akYI6vdwuTqTEBuLr
Ko9vP1lRScLC8rCcNvrmsER94sxsa25VDuiCc/9kiJLfsJgL55pnB5hAUJLJObqM
qTXLUssNtOGr540ghi0dFPvmLE6QLLxb900RhWoYTw5+/NSoqt4PfRdbjKbbb89Z
/BXXOU4IKWSePRTdNlAvNcYrO5AL8yKyLhNL2fvQrXxF97mRT2GPATbEBzW9N6Xd
tmt4VzJYwt0jByKQbSH/l+Tn2UPD+nSdpr6cyuz8dVjQU3BJFIo55XYbbb9GMjs4
lfNhV6/nGU6rV+MBa7kg4U92FrfZvH70pYIxWcOXtMomvaYJ+auOFJxaIzMGPxCQ
5ieAeuMp8gEs2SLdVe5n3Zr33sPPjXHgWA178Zdj9tPhYZFwtwpN6a4sWs64Wyqq
uxREPsUle8+nhWTrE+X2bq+e1+BtyMEmOMP61tAzPhQMIYgYObd8F/cfSLQ37dYO
gS+cExpR4o5PtcS+dd2rNi0jrbwpSi0cdHrgk3eOaKJch3DvTLUYsXPDYhfSIQ+9
PJv7WSJMp6+vZWaZW4o5v7MdbFvL2e1Bp/vFJORzM0wbZgmmQQ0RatGnEnAEpR2s
ydgLlJpEOcd8dIdHJx3u3Wyfv7ZiSMFP4QImOEGGBiKcqs0m6jaWs+Codz33D0dc
L0ktmLXseo5ZPBG0VXO9O9ND+pvx8DgAoUbxag0TsHqCL4zkkWeNJB6e39eOHM04
05GmH23Ijr5H8AiP1jANXFw7QzlBYzZr1xIMaYgQ6K1nHuPEXCRNXFVmCoI6ruSR
A2tYYWoJmzTim0/V/+MRjZo93uNN8YFZgwvKDKvIQf1U0C2Y/Fh4fNStUlH3DEvQ
ks4T1BCgtFp3H9e5xb4cSXHJM8GFQBv4pmrnbJU+InCXsAewNpSG5OAeC2kGuaFp
uUyySorTEEbIQ4d1+MSc7RptXSjbAhiJsMRA/ghlvoWHiKWLQk206a5nOfMwzloK
vRxBnxYBCELBMCVFnjPoumzz0uwmwoXzgiuBLAEu6wHrdec3WR7XMgpmBSl5SZOp
KlEuObJSNzT0JWU+t1JCrdYov38LqZ5j4egumKg7FjZ42ErYvBRUhC2P+BC38kQE
16ljVG26cG9PT+1n4tPg22TuSNaTxbUVmsj3tkZv0k2aPRqTnG+YCGR+P00ET7It
ccNrZTEyFA9z2Q47jQ6pzY8h3FVh7zwog+YTkaAMAg5YB8yzRsU9lZnOAnhU8PDZ
ZXDeMMxsNByMucnBBJ55GG40Ym1vHAUN4eqyn/1FPbE2dBXb6ii98t+WDiSm28zw
wOrvziYfy0rfTp2W3S1+DbLlsF0/kephBtZRyGqQNhNXE9DS7NHF9WUSriCb2eP4
FQO0/XAeEQcEub/gQD9jocwtvbttht0xpn9njp/MJNKvC99/myLnZY9P26raRBUp
mdJ4BK4eqcMXVdjECCxfwq/L2wcaL0TAVbMoxKDntLjf9y5B80jn0Sc0fLzo9C+J
IIrt7X7bwuJ+ungco/g2PklY6w/ZiM2rE+GOOfGm5f8BGwpUtKBKlljZOPJibJZU
jZELkwGdOPLYJkPJnNfcpcqswAHpUQs7uDqR1vTqr1Ki0+VAfqCqD0htoYggAonC
TVtyTxApzgfI1tCNJKTiojnehJC91hMnzl0+DidZwefcPlUpxkFFiYYPcUmvoPPB
/5zh1ZVQnNa8YS3BemG7tU3EStLmbuDA8BfN6KSK290QUWKFNUmMJQeIqRVBm4vB
FYdHXSS0nP4VWC/pBPDylP8ig5ScliIWOuWRJnovtnTiT7/FN02uDCUWKyQ95uY4
DJqRIPLFEHqafCJaopvdrQ97OI4WJ0hbd5Y3HsdOA/I+piMK/tO8oFMDBZphbDAN
Ak6vvIoxo/ByPH+jOFHH5/pZwIonxVXUXlJANZabTQE6eKxkHXglLSkM+LCXRT7m
ELK9UaomcZbFjQNSzZq6a0G9b8EbrfGdqD83+YzTXYunanDKoJ7j5warvXKIqKd7
zHg7EopZ27Cn331JkP7Jpd8P4NaIoLY5czxorUVpv/FGsJUb26vDgV+oTrWhbvt/
mGRTNtyjjhzVdvZkJl0sCIHsYOTrDrZXTTuy9IHlA0SCa8jZrfdC0yLibtQB4KKC
+vn9bxs2k4OAIDl2sSha+/hwTwr5whceYwVndQWtRQJb4V/wAESJtDAQV9LlLVAj
NFCm67VlBGVXn9XIS4BSQGgTwDltw1KBFBktiBcq8lCeJbUZYcEgbF6QY9lK/coP
qUC8daIJqU7QmcGStKoVQ8/a+qOWQTJZ/ebGNym4vN0TbkaUXNINCaAHrRhIQe1z
vPg53plv3gw0tn5ZiDVCSJcp0gikUWhcfcyG0ht8JyTvOiAvoEROJ5XEmYujcijE
+mPrJOg7Y8RbhZI/0m7MQBAj/BDKTeTR22e8qEUCtaE4bKg5UBorcwdlEqNWzns9
dOUpYmLeG5ieM6LMh43TayXRz2brYRm/EnmUXfoBM9K5YJbNUI4sDOQIevk6EIHB
KGGO3i93fTh3ks3vs/Tz2XWoEaaJPx9sXQJSSlJb3kbWOPlZzFF0jiKJIHJjGIv8
rJJdERAI1Pkkl2SUNAiHdPeCfMOLBoZJ7drtVzYqmaReqLiFAmTZTkzBfTWRBIyV
EkvLi9kY2azIPuzMSnzGZtELtiAqB5nLgzz0hCNSJm/7U4cqdOtaK8QtmfwlRUxj
WPadvRpRj13BOcRebR1cuQKQovaOCpTKRsPmW0j1BGZOur+vLoVxydIUasv+R6Yr
A6pJLs2Lz3ZOa8qp7b4z9QAyJKlbmGICebGJhY3aL3NeOu/h5eIA38IeSBlbk5Fs
eZeUR57L4TWm2BROTWWa7dT/xTFwHY4RKVxY2K7XJWzzmRikgygcyDj/O/Vy69Pu
RGSDoHZxk3MBLOvmBsyYmGbNSAoqbWJsGwA9dR4f8XK9Y1oUxHOBNn8ybHQSZu5d
m8kChueaW5EkXZBjbwOOiky4iMH9DxHnUg1PA+hYxVVMZCRop+CxwvtGXGYDgcsn
t815g82xoEzYR2FKS8fgxFtaEW0kL2m+6ZJJl9ooV4lBcyOp4tsoOhI5uoZVeEfI
HNVPAC/cPgSxZ77X+IbCKhuWG4ge30zhB5E620o+LDzdZZVSlxQ96bg+Wt7VWKqu
ofRVW8DxErklu340G0/jFoonpXVvWO6uJrpIhH0UHwn02dvYFOvKWaQHGTOLhWm6
RPF94zE7yiQs7yrHZ1EbbK1ibJujI5P/LZS5uYGRY8QmLVpPxqHwZKMhVcAvN9h7
h882ijyKcgBah8JC46nCM43YifAk3cxelWerAvzUJ6jSBxWCHnOzYMoYVx6WcfJY
BNmLwNh1UuP8yCCcwhRmaozA1o4w0VpOo6OOBWSDgqXvwq/34+gnGSnR0a2W2eZw
vdFH4Puw/hkaxvg5q9O7RbLpn5eANJI5K332NnTd82nh4N9lyI7zsFnDKSNZ81jl
UZZUi8P1nOyLhlLq2Ct7xWKI6Hgz2UEzJ2eQT2Nv6JyT8tcvMURGhQf1U2YqLTCC
KdG4Ha/v71egXaVTnxFMnR/jNtkkHtsylWoUdjtCGgMTUmLzcTH2ReqQu/dyMrEB
/ZMppo0+CNoqKngPmtGa2Ssu61R5IPWIo2UDHfyax1AUuv/6Ebhf2eFaAkwmXPSm
oVliOGjLwSZ6OzWMNYQcZq3lcWkW4Dx7ajLgYyJ/Jyeq0bFh6kvEgrgE3x4Wdwje
fjjOeJf2EV6NHChZompHqBOtk4bQnidg8IkN0xwTkSLaE2eTy3dH6taRJIvtP4tq
J7cnG/pu4hODk+kZQlwoJ2VdaqF/f3DyciCbJIawJgWlhfS+ydYGHEvSRDuUbSLA
p9hdVhFRabsxJyTf7DoExgqU27wqHeu4kjqBV+nxphiVhq8x9CVZjyCtf9/fGKM9
e3Qt2YfqYVAzr2K3yoy/wBhfNeDJLZUxHhc64052Oi4CSyr7ZfxSRs/ZSGORe+pY
ALkWb3iFXKqY4GG70c+mF554rAmjePczx6QjpowZflRY/0crLY/AdXCJPI7vwR9L
9/YWdV2LC6l4XeCqOsioYw0Vmkj97vjF9rqbw3zwYIUpsauqlAElEpVoqbqdl+6O
v55sxPBvHimo2xbkNmcNF7PhZT/Q8VFMlTOtNiMu31Kd7GSgZyjHN2fcc+JZ3o7T
I1rklqoAKcYLOHa6OU+yN22N+wd14XGHO0+X6KSsZoP6RGRuJK1czBo8M3YuAyXS
bPVb5w47LEVLmDvqjDIaEXCNOPOP/Bp8vUmjkusGi2utZQvILyp3PWLKX8L0SlfV
Uex5ASvNH+4ukmDFUAM2cet3fN6DtR2W/Wboz6k25GailRTKEt+P7DqVRC2hdNw3
ASF++PBHPt7oUtorytDFAaxrFCQTO+rNgnB60Jzksgbz8FgBE2YdmBBRqEjClyNo
Z4qS7Epcn9WI/TMWfbgYB4y0UXNriVXB472sdOSmDyqRxluaQHXVE1xtJkyRKjzc
NvQSlalV1VjcmmIUAA4GwKgbrhlBuaXT8s/Hv+ObN08LoR8TEaCxIIPy8eYhGDoC
eHmddjthf3ZuQRxdnuJOdMseDbabpJ2A5Rdz5MEBzhf20gh/wWc96LdSIwIBfILK
DPtPu6C/3Ag3rZR9/xbPex4s3F07Wj3hNpJD0OiyEhbwrT2mBCO8jl0xLkFrbHNY
QJ4GgBro8WI0oi+ZQY8N4zXD1/7nqAcAKGHeiRnTqP6KBMhGcHq3o8fWQN4heeDM
BRHVU3ZpRRmohXPmG/a6zTyv0exDofpXHf8r+JAceXgjZtynvr43Xame2IsT/rav
AxEx5OhK1eGurd7/DkJbAk1OOqWUP3l5qHcCw14Q2CtIokxn5gZBLueVnO5BIFnP
HK9dEZrx9qgtTUt3WdZWhCnXQT6R1NF9StPPTSA7TNgC5/aKqJCKO1Hj9wAJyEzM
QIAcMz7gvlq8UvignzXddJNS+Emin4o3KpL68QtZ1xixNgFWeW1gVF1gPP6ClB+w
h7sGWveBcXcSYHy67sY/MAJeYPkwZGlk4IbnH+RNjWj+oX1qfMUp/SJ/b3iMNVFj
zE5IM8zWru8DIIfxUJtP6vLGgI39jdteBUxy3GBHRcaztZX/5yXeO+eW3OD6xjS5
wi3U6fMJ1a9GyfXwDmUbmAFmT142408k7vWIngp2MeK0952lrN/+9pHCwen6yuFA
/KvSh70FVnJkhyUNLFn3DJJHGwz+dxjPQXZg060B420Ni39HplDNPn89RRO7uXPH
i6Ttc1hnoxWWqXzQEM3YlTEg57cLb6FDhmQqxjWpZdT3UtqAnpsIb2hu4yKTHHct
Fga/JVPDSNc0JeuWzU/M8sQ/uiUtzkIIjKGLB+CnAJ03uGoay7rGsfrcvcd7smPu
jnNi8+qeilReE69/z6SseV6pBWkIAy/zH/CyHZKRyq/9GETN3FzJH4Mc7Q2Wqrw9
scA0pcEsUVbdBDuvTsjPbvRbVVq8s5yeJA2u2YUdb1lA2AvMOr7Mlo4Xd0xHskJ5
Pjfx8tLVSlPd0tdX7B3oSgvEHc6is/fDeNUkbsxjSDYMvl5H8nyQXWtlKwUUrmOz
p7wbCUr8zgSjjnizoCrIV0c2iPmbrxBOq5sE4oHKicmEHsyTCFhI/fiVXX0HzLQP
luyhIDAj5Beyy55Z6EYWixtEBhACr0Jp/DJeNopKFekUWHMQcn8H8xi4Lirc2JeM
O/EtoRhRHJfF4hZb+2fzaHEtu5CjxIn8rzumh9jmAh62jbZ727kE+73Na7m/SkUJ
1JeB+IqFac6JH+e/hoJIKOFJ8eJshBRL2/AErTxg/gcW1p0xTWy1Ajqvp2qgjS0o
xWdRHanRc1oPUNdMIJfQSOf2mmsFrsPFFHqxOfI4LKrEWFy3VbjJKzus3hq3A3IC
BQOdkLByjJEk/H70XHpEwQPjVxzovP28GSXkDHCZgrAb6cUsz4FHJ5FebVg/Nnlm
qpV3+JAqugbawso2n8HyH7U++aMa4f1vSZnTsGL6MZUkCgiailGBhavjVgJbIyj8
GlQQUSs3CdyzIwgpZEpC6xZXp6Z2BISGhbxBPIKcyvkcs7FZwKVb9uGKE+wuIxfj
sG43XtX/Dv3RCHcSf3P/JIQG3MHBBhm3X5+SotK35wTRepyIvNbWBMhwO3x9pYnO
dnN/PimnVzgA4DsUw9GQkR01skxPzkvbi8eZbCE1alb6ykAYMJoc4Q1iYGOPRYjh
y5RPyCgbGDAcq3PDRniDMt9XUBck5doCrMGAexPW7MzAKp5fH+JN8+dfoXj+zMoZ
TyqCHgWB09U2bzTZwMEa3rz8Yh97JaJNj2CC5unNgwI+lKuyyF2Avz+vlmGxusr4
mLcCTumfTrZBIt/AF+JQdopCDPl/tep4gIa6CRS8rPOSkTp6vU/8kui8sNlPAql2
Q7qEVEGDvhSKHsjrCFFXBqqxGkSp8RH1EZFn1HsywAF2sahgBcOE6udfxfKgz2bK
nVRTXi1AbLkXOsFhX0oEZHJujdS3oF2RuSi7nnarEp7Nqa++JU4HOzBijt9yyW/g
KOwnaejMEs88QqfMJLpPD0VSWyqYuT57QDfyXK2aTJNyyFFT3RhLXvHYKWLLlUSc
viViiWx68R4w2rKbm1/FhPzflfhnml31DXf91HYPfvHZoUK3d5IrSNemtP1NIKp0
4ZMoowy4x8yOCu3J3ttrA87PcOxyvVKhkWhF+8m/fWPnWJqqZFusGKQ+ndECWySH
OGmBwugS0WeH5LiZTdAICDlGTqfegOwJ0PjdWn45xnpqmMYNnz1aeQYtQOEItFLv
4/tdfuuXyKdYlWZo2zZILE1zQluyZ4naumOz0XdUtpkuriK7r3Z46OSHKj0Va+tQ
zmUQqMjB8SmqBvCcPCapKIR/8RndVYESClgEEWROMEv4UlhKMU2W4I/T61XRiH9s
dU84DEucDiExoV98zFv5ZY2WDwsmxWaMeyyvV0fF7afv11GHalN9uxHZTE7JQrLs
PYUz9px3x0NUDoDGrPVgnV4hX1iyqb+IgikqbZkDsjxs/4dMAYA230aliQCbwPYT
Wj6XoT3XzOpyD2cGA0qPIWYxfJTfdDxgvrUBFbdDiCrrk6ZyS2kh3jbCJYLHvkHg
QtdB8jdX4mtHRJbO/Sb2rEOjbp4MJ8qykCAmveD0ZuVGUFzrf2SHeMA8ODwlBZxJ
EWi4alWtZB5CqIUTjzcfUE3VXCaprSKnZOpmeiHMfHk1q9x2pwdkkow7x6G6AI4x
k+PXBhpQ/08l+uWFtc2/zxfYAOgWyXNl07FXZ9zWpCXND+CeFFN5q1nmn+xnCmSk
0J7bkMSSgwl3Fm9dy4dxFoFmvUeExSZjBvYusQeyH+qYWXCpXG3+b7yCWV4yc07I
FGx6KDHH5eQB8RCGcjqC2JI/eZxZLWPV0FcEdsmohx4bmoLcdKtJfJdAfn5Iec+5
9OCJgpzC6KqB2dfBhHnvayT1U6TRG47P0lzVYLasZfIdM2VbtIgY03Lpr3yWZBGK
TPbZQwu11R8M2lK35icN2L9J3HxC8OAnqR6nlN+GQjoeJQK6dCZsSZxZn7cizBst
V/UKR79xH2sC0cc2/i6wfC3TTniOCXwcGdwKJim0FmvA47iuj87G1AIvkVKPVgir
UpbPihhihD3OWw+lLLX2b+uThnZC7+mQ1IApqPXsj7++KFE9QRmokFbx0kTp6d31
pBTgvo1MO63aUJcVM8Jcaqi9dL2VxPHtI/nTlRP7y1RQwkMEU5ffpg5Cl/aVdrpa
31ztNhYLfjTMovwI0BY5feNJ32vuVjdj2Qie2Z2nY9nAh32Fts7yBsk8573L0AFQ
clwen3A19Y/Lv4YWklm10LD1NNOdN/NbDW2OVKa/U5AJSJ6ED5wwpgA2b6LTQh7M
3BbXfbYBxE+GZfB1pnnL5ZJgcdnM//Ll+jyden/xSoHpDuIxqOX8IqvHC1+LQp8c
cGx7VeOrzgg7+JAGutYhlQJY7VgNA2LEMCRNnChUtHpxboD+7lSFIGwgFMjLzBkZ
LrqJSouYIOkS5BqTM+5gQPTScn/GMdOcxKKaiCt7d5GRpnWwbP7u21215poYQqu4
rHJoUxdTRxXIEUiC7pU7Y2wkYM8btzcDk7XhvZehKlyG7Rvw+k9UTr5A3yjGSXdl
5HldBOcwTDwiFrFDTKXDVGa9iKAzDvjplP8bnQw0+Vq1SqG+CZ/mwA0EkAi3m6eg
2K9U6tXcUtHBkJ8hp7RE8raw9DR0yoeKE5rj7laMwecPoX1zXfyD9/DMJxB3ZpZT
ohtD8d68CReb8DuD2/JrqOMXWkCY1a2jxV4mr56MFsUmwRps803Scz+hQs8gi1eS
ohY2+wtdzCcdEloOVCPp7/uVHqYszOjOhtM0tdLAkbMKVJoduNlsVAM+2gCmbq0R
ijTkEmCP8+cDRMsKnXSK966jzz/HQlSb8LpHcPq05kB23EjUYKXruw9FzRxb7Qr0
vcjKNn8ksr9zhFZ7FqhBMYk3cIbtgiHoqFFT9IcHXK3VzJ14JgRQiWvHZ3ATxI7i
8rZuBCdFWtz3hZtI2YJw2IZccVnZiqB+/sUGiLPorYdqjyOfFRQUtys+Esec6sBZ
Yw4h6hv4F2MTtSBzjjKqXbpHL0VuMF/JyP7Juck/9JyADg1CbQNHt5jUpjz1eFCl
ceSf/DlDrrRoSJENTgwZjQoS7eZOaFD0hJ+HSXcZ7ZPgdvW6BKWfUpgzBZLCRHO2
/Vi4npvhfbjaVuWWfMH7J3mGekEkUQwgZc/azxQtDYbQ0zbrQnrWLTxQ0f1zhtiE
1Yo1LPbBE1GUmozEUDD+y8CQTwu/d6Inxbtt1DKttQ9DRfpMOjB1wNQ/9JFj+44J
PYYjFJCRS+uCDIlPeoNb9ub8BeJ97sQ3Uybl56W8the9PLc62ueSMoVF2FjvlEmE
5w0dpwJLwE+tGIW9e2dNQWz8fGYMDM2qoQZhKZ10pqts2tLPkUhTokHoxSdB7Vuo
RDRcPbnEGku9il0IVbvf+cnNN4FsYmdJ0l4tFiGms8x3vYB5yCah7dAngERIY9V2
VPg6bSn0e1Nh1aeV8wDFsK40sJor3wOPAAJEWsJNVnz8gobzL2AZRF7t52p2SR/D
YhYb4pJFVZNX6CMO5WSTdYJHxpjAC7uxseKSIjh5fABY20XeekyGOhZuu9VV1C6M
lAVTmnLGnVZjpbz6R4dbzJaiB7p1hRXELqzO0ahcgXdwU+i3jlWWTUcbWRqhnfY8
g8Hj7srKouSFLNiQZQgvyk0X2fDPPhdv/3v61+k3HtfA9C15AB4Vj1wVtpnuRihn
lmvv5IuN0NU6HJMsVcjaKGbY74JXoeAfdi0dNKedhOhZBzd8kIAvDkawGjX09nI+
pXGZiokB7XS6Cpa8jlz5KAbiazsvlIntONlHsjn6fOFRCaTrV6mNiaxEo+uzvqy2
jTEqTCAIexQz2kBAzWGn/GwuxRG6emt1U0bp1ztRs4dEcg7g5pnznwxcVViwyCBZ
YbK9klHkhxTM+9zLHXo6Q88JSUVuv/pbWt0vQF8FJ4hc0z1DblZ/yyK3L3Jv8Fur
7Hsx0d81BnzNC+261tp22E/gaWIy4tH1EZ4+V4THgewaI87GZ/7keEHuWveixhsu
i8C7mgKN9wB8SdZXSReGnFEerpT9VpgFZ9MnPhSM0VX/UOl3rxGVrfI6Xgzzpp5d
YHoaTV+RFR1Q64OXQX5SOv2lBBp3womAmNyCkacCg0C7ydqZ9RASMCd5oF6oGYNO
Oj4O7CkFEQt7jqb92VyPpWFKMAykVLyB+inQh5c7SGPjYXhpox5vKA26OFDWGhG+
2JFCWz4kr/u1dTRAIzdlogC7zMbphGNBccsCK5vOScHda9oBMHEkFtGeTnqzpSDX
JvdfvOvMJCjkUN6c2/IRHBaa8MZ2ot2yv7DWEQEe7x1Rv8Mv0omcGIZfwVWXg764
g53nVHBmyoY6gU2RsCKDRQJmWKDHrHCCJp6o6dIkXCkunOsdQ+UmCy4Sv1qZHy1Z
vK4wJgyUqIu69IVC+c/W5UYY4SA30l5SFsXln4CgKhLswmbfwUT6eOsPimrAPCgq
FGJPsYDv1pOMUgCB7cBsmXAlsh2mAx/XDdfEj+l+ebR6HptArhbUaGoouCpH5QcW
eCYTQpH9J49H2l2R8GCYj0ZlqDbc1XxOV/HMneRO/8dkimc38nQG3UAlVW38HnBp
A5QLxu9JxkTcZMmy+E061eopwPhqWSqGoUQQ0Yp+R8iOym0sN5kU1V7D+VpRcBEr
iUK9E7sjhRgJPOUHSx4TaZheB1JfZO7qan6oGC/ypThu/61MpYk/O/06oFXnZDCd
X8mtMuRIcaZeNWniyKdTEQrsML9HN+LGsiEeLEXDerCJVqK4g95yXJmP3PkfQZkG
rbztcWT5tYJysEtDw6WJIv8/b4IvyMo67uObzJoqNLa37XDOfYXurDxkn/KNxOkI
2j/qPl6zixZ8ErhATGcFnmyNnA6dcuIAUQ93Y/MQlM75emMSSsRYpXbwHQCU4X1a
+zxVkgl6FBL0gpgkq+wBsXtD0bwqjTDSjmSKeODiugJZONfndVd87htAYb19iECC
xaO3qSsIvM4QX7QM2op+upIf4P7uqvN/Fii6SG9GZi9u7yhb6FpLKqElDc2feOmF
wFHZ+8iswFnE2L6bXRIO55eJpQvHWnXQzP5WwCsOCfv8sV0Bjd9Dc2+ElB617qmp
0DpLMc078WuTzC3nL9Iose+8cB9uh9gyH5/IbTgabVcyuhp8HwyrunEt0/AzviK6
Agh8AX9AOQmtsUq22Y1tsoQMqGI8ScB+43aebiDkV9cw0JXE0wgFSCye+69XkCvj
uVxVFxu6jhgtILP0dIB7Gkrhf5Qt+4kfyK7WZ0fy1l4NYxYb91+vOz17Od66Lb5p
sSuGwxk6/22ICTixTQgjBVGQdja+ixjOFytldD5HjpkCZ3z1CSeQpkdZVmTQKwdj
Komgf8ilzxui99ykKog32lYJG9AXGKBr4cEaDVYlMyIYbNxjRf1FKvPwD0UwLJGk
5sVUhXpT9hl9JinVKCJtIRDmViFDBxIicgDnwI1fzup0PCW8GAaMQUYQBRypMFJq
b/eU9H9EaPDWOlAogTAQSocSYG4fY4sECIQBsko1DyGcsESDWxrYDslqbwifz7ZU
7/WzomoiVJxBnfCgYKCy+sRha1zlMxr++IxyedTMgw8WokBVCKQDgdho24IQ2frN
dFnMZDN8XE78SwUMfqkMeu/Z9sxDw6DtnpVnBTlbYev7Si8Q7n1ubnSIWfFEr6mA
K5dlOqtQHgaUh77GXHRW13Og6tc5u5oA+bxS7N3u+++JY/ZNlgbzOFK43jLge8dM
/Zt9dhN7MxKv6OdtOlRag4wPja18tjEICuJii5/aD0cfYxaT9zwninPUimjr9rev
SJYKVbHlGSTtezV5r4n+PzJvudkraoypOT/yU/mSrvhMvp7Ye/L3eXa8OVBOIrQa
FeqlF3Nn1hmRYoiG3opW5JIwcm3PHPMAIOsQ9XcxAV33No6jUeKARfTxEad3E4x2
WzNRmGonO+ktWw2071h+SUfylYD0pqLgWRRaVO2O1XfMnYaMQFD/bvWBGVqnwsmH
2FF5PMo9QLDZQlcDxlzSHdFcgLokeXdvHc7u5lqNcNurYqdMFsaz3Nmgvp2iPtZV
wUyuLFrFwKoEWz923DDVb9DYcZ8BE6fHum3TqP1V2tiTI7RbIrGXmG2BRNupNx6G
b1IsK8MJT42mafJist0/Jt8cenD2D+NFhNwUV3TJ5I9hBE+DKaeD789Dzpk1k7sa
k0rFqFqUsiSlxpJ6BSwboheGqJ7kpHCy7eVwx0ThVxVod6wGdCvMFrOe2848qiM/
zU+62ekbvXVc2iFiN18JWRJbmz0moFRD6alghTMciTCyy08HNWL+Hk7JNAmG8b7O
VDpcwN+3Dasn505t/ozt7HHeYjvV/YtHQZvqK5KbkiLTXVNHbmACDLqt513lxCjo
GhyJIXzuugIUKJG9EYPYCiq3nPq7/RGSFfWtMhtEkcEr8EUdvejXm/tA44j/+XyS
96SiOn8vTuMsC4v25m/MwjuJDa5NvFVs51IXidZaG1b0DevbgAoW6D5Rj2dWqGTn
k0cYpeM3dRO+vAVHI+6i83QQoQKXltK5lAAAHGefzKpLUzOJQl3weX7yg6yOsxi/
g93V9gkJ9iFmIVwDjNrdF5hdpEIY5hapyQdgpWoULrFlK2PZUMiuj87LX3oK7RmQ
t84VlAtpA74HWvxM1KJKjTBnaDzaGS3vj2BmiuohpCz2CkaiV1r4FDH4RxaY9vTm
ypk81LqeugxhmtqZrPGySazN7A3Zoci1/f8VceD/aLNdKD7SjF8gmWz6Ell2ue6Z
UBvTJr7qRPNNTUR4rhHKk+geQ/1oYzs2WMPq6i+4LWBYpV90IxiRbWeMKyNhcPC2
lf+k8pr2qz8G9gOEU2VuxjzjbaqeAFCQMvu4FDRLaytQ2qamIe7eBOQkI9LF9cE2
uVLOeGOJjHpYCkSonmZY/6otYJb2v6k6G+fjNvlMMLxY8G5WINd02t1FCFz1O96t
9Z07q1DYc5WaNuCsslfZ/ZxgSphnm/bcqiIyAyha3MqMYkVsvu/Ktl2AtgE32hhI
IBefcaocK5lGaazN/7ZeBtI6ElYZ9MxdVv//YzMFLAUCMaANAIDV5gN3UgoBorrI
V6ZQK+dP52zfEfCRQ5MV0O7k0zvkBOqhmc0z2NJruwTvDMlWrBGBVc7SDvwrvyTI
BzTc3U+DRX1txPE6ZnKeIAQTrL9fES3L6YHkgljaJuJ5+tmXBH8/8yZc9yraVOzw
PtaINVr5bHhacJykdanX+MIDam8zsdR3P1mANAEGNzMWynwZiR7yIBBo+ZR70grX
za09c6qVhaw9W+93G2TLufSWJnnkFnYpwtgXlH1Ilvi+o+m68zdPrGfaqw45v5JE
jkE6utvo+UobuSqyyKwA+hgFdeQfpClNIzY1D7/lsbwMdUI8kHJ3/vU+hJB1AHTU
wKtOEpqdnthDePX4X4cF6a2xBuy2ga8xlgqM1ZG8mMZ6D8cFIvMOPctR9yy4Z7L1
aOupFOVHw+FvVZl7rNOmZdwoB/0MnexERwunjSuOiuPWeDJA3HsiId2qSYj5GLd+
1LFmj9dwjjbsbTnZr5r/0xz2edkh4eC8AUoPJmU8mqxrfSCbZy9NEWqMsJuG3yPa
TQXvRihPnsTKqyqUZa3oyR8kb48voY7lLj0NRxPXxSuYxQO3kR2ympe4Nvz2I9iC
ONb7D8A8rsBa4C5da/GtweOPEQeSZ+cyakuvRdzADzAigFBJtKIkIMu+fJmPrT22
zRjR0l35WzfSM4X9sFxksRhiPVL0htW54KYbOwMwHnnY30q7Odjl42H51b/YwW5M
McfQvxzPFzL3mdK6LK3qKfsAZSw6ex/CeoCl9dvJiApUZqIuoC/bpVx3WRvmc8vu
nMuwRdOPE0d30vhYsOWLps3sg/l/iq2abBRXSyYFgxLmftSew87VariCbBH4tXoi
TM/vvtoc+UuDdUbG3nWqNJ6alZLEtHGsAh2puWR3b5m/UXY9Q3304cltNY4GS3ia
6u5fh1LK3CohVhabtScjdsblJ6e9N1x4Hr6SGUgto08cV3GbDg+wFB0krpIUYtgc
rdnjc74HMphF9DUuRGqqNcurNJ557+3OtlHNWdnI34C6SbNL1v+P2c/9YrZFA0Lb
v1o5DHVUJmxMhU7uEJ7RWlR7ijMtlgrE53VClTF2dSBlk28OHt+YJbVqTVrACmes
cT3RxKfX25cyiIZEbgg6+i1+3g3QsXFv/ztmmpuzGDa+Of1qQS1heuu/DqOMIQIk
TAP18tyRf+GcAARXmfDNGPeJ5YxeAd7YIAIpn9TFftcmeT3Juldwq8EJztoQHqw1
MfNsK8OWdd/iGzdwCBrcVJb6DMbJ3qCZsjAarjFO7sm3Xs99KIoEVh3S5umvvM0C
6IWXjC+GLb0YF01h/v4zocLpFqW0E4/hhVGmGWcL2+nW5hF3BFkg+ixDs+h2vk9k
bwrrWdyTn3c6lLKpbz83upw9GcnyLepP7YJNXiKLXTpZmLib6QsJWsal+fP+yTrh
ceWX5CXhE3ke7uiY9Umts9vIwSJZ/VAl1Dvwv3boGsQ8DVlqJPdqEkqQQRVY3r6W
Ovsgox76U8Ihvt+OahHMsFrkFfcWXV9m3c1r8GyanKAOGQ8nYsS7R/hOmMRWtdWU
savMaBY/d7d4goKpTnMEd/WofWNwudrqqEu8ehXMqgLgcQvOps+giTKlt5rl1Uuc
eUiCy/opjQ1iVQEdf06TNJew4iRyeO1h32LjUiyYeigYo9ZMJ3kqDsCzz5ybZMjD
pAtsTg42Ks5nakGNZrwPSUnM3FqwEofZ5HszVxYTdk+5nrQN4J0kMgYzoGcdatEn
goWc8XRQK0QdjUhgnbrInv9Ui4DYCi6RbKdvwOlcbt4ddoHRX0omy8VD2I+yQG3w
oY1IuyyMCVqbCmfyWqMfEnWPlQAiiu86U1gOG2xjyw/2au6UrEFGITxh5ijinx9g
CUG0DvMdh3PZ28doX82a/SxsQ5eWsLfPpae/SoyEN1mBQ1I/0bYBeWa0wIc/J1KH
2Ddn18oYimQcz0I9Wz2nNAa60kj98VKBBlEVARyZToh9/0+fYso9/7ip8UIZFh2g
0f/nndDgSSuLiLZfLOMndEVBIHbLyp9oYR2yl6K9RzG/o1IkOYmAoUgqBSTvha1u
x5ogAYyFIdHwHDFO/o7Kd+XsNEwsuFPbr/he3sxQQRGXqGxw3Wd5E3nfqodRACPE
ur2NgTc9J34FLns6jHXWsYumzsACSOQ+t1XWjqBTbsHnQ0IIbwfFABhzSckDcZBo
p7KFbiwSsW+iquJ78WGdpPAgRhedpxFRx8Ggqm69+3jp1257eTQ3p/B1AGhseORo
4XUXb4HeWd2+a2Qd3By6sn7/OcDkseYlmY20W9QHM9DpN7sXEgpVUoqkrg89dHSG
4GizT74eyHOmtrjeGNjk4P7nhaJGXKA15znWO7b87NJTAjERh8m5t/2Pfor3U/AG
GJnsDpTmZ/uqWceoZifc2E6Go66qwVDvIPT2JnoHnJSGwccb9T4u9aP2QHN9JZZt
a8/YbfbIKvhK0sFOmb871wQkDadwUcMB77e1MPZsuNImPYxUuO3Ws32aJ9OW+Rp/
nhKaHsJ72tlGxKk7KLczVUvQhqR7Nx6PWFHP0wdj02roIXwQUrjKcE96FVEwhMHb
Gs/QTKDifslI/fMzQcFWct0gJ11QD2qRWui5NZJyi4BjQovDU4E/Q00Kb9wkF0gR
+4wMIfVHqHjDEZ2r2bWa2tzYLlqg1Nb5GU55I06cMbiFzMbPbt0rIlcEs9VaI2no
yDBVqdjcTrRAuhAP/UBayepcYw7BvrRFV8p4LqYi+CMqPpor9gPqmhqG5sNHWvJT
E2f3zw/gQeC9CY6Xv9nGSgWJUQwRnBH2HXLhK/PQxFKYWBInne2OgK8wQnlIx99n
50OTdBr23QUrj6OROIxs2eyZrtk/w9tzSyH9PAAHH7V5KjvefCFV5vB5EGo17nI9
TdOyDbhgGlYUwrnMNJh6cjf84cZoKQcTTjdlqHauKHqJwWNJo9PvfeYyQve6/+jf
uaZnz9VhFALRfbGS89sxVyz+iuYz0m7bJeEapldvU6L3ZRDuvpJ4t5Oa66adYgNJ
z97VkgwthCP1UTdoi49OkmOaVCfxzkoDzRMm0Yfk1K7rLPvaG22O0am0ap/ewnV8
zgTs7W4UtUNaSaKUX1tN6NxDPxtt+1t2WtvHjgdM1JahYazttLKmB5ZkchfduUrN
O84p6mreRtRfQHENVIRomZNcg7UzlfXhgtLhaxYyphjVZP3LzOFVD1gS0MEbQTNf
j87RSkra9vZ4+DzavSIX7Kt3lycNYPdAs9WpyODGM8I+C81IPYf5v+p8VwxNNNQy
YSJN3woeeYEWzluWxfjZTD1xj35TAqrYSxYGNgj+ABBTA7vUc9qluXb11Wd00a4M
1RyEYPa57ZTLnCIiD4gQXi4gZoHXXeYMxN7H1jYmqm0Hbc297/OKYYyCdqRP6adC
qJ6jefnsPFPf5rI6ao7JTgWxPot0ktEadHgFxZadDC8HBUIKwxPA7zVo9HModL0N
N/FITh+z0Snh4M6j+58rwDUVJzrWQ+ooYsjrIuoNFE/eh1+vCbsukeQKw+cTd9J9
1v4oUCzHlx/UxzWg58/iVJlB8vt4QuY79CaIoRvxWNn5uUZoWk0rzxU0IMn4Obuy
5EiihUzUxplFQZUedsDG3rUDG3rbmbee+gMmn7Co9ZbkDeJnBeyld6fNPfPSp8ZI
PdJN4uSrgci/9e302Ky0VFhBGNSUN3Kuw+Q+AcPx6xwosMXtCez/2SnMZG0wA1NL
ywKhZT/t78q/V0jNQ8dxVHsowTR2bCaahNbOZZ697Sm76PnddSxlvoK7gFl/SsiH
ncFSU2QMSHiaPztZZMK5BEfkTat7p30vbo3KwK823kjO820d3vhCbqykczCdvklE
z2e432fcr4mBVh5OzWZJKG9mBfqhSSMg6xRutB9IJqRk2gIK15h5koY7LjCQsd36
OCcmYLILbpxwwYQVdZZ/UAEkL4IJwq0Km2x5No7vUK6lZxJ5Wp1wsnJluNCIXwQS
0CJgKBrOA9vQxQKdEnh3lPXkcl1D6wpGR4wRRj8XM89tsV7kTBbBsWKP9m0t1zbH
LPP728+mrYTdFvmA8LQUBT5JVb0JvJY6jT62xnK3y0CaQpiDEXfNgzRhfr7/bb4/
0DSZXsZpfd83CS58L6RbSE2vTei41q/cR7vDSZkY773ypEwKy99SRXw72jseQYF8
0DI1iZbbf0MdUCdmQMzHvZWOEhq4QoZjIDOG7eRuhd5GcYJcADy/nOJ8nDiq4XZy
4LAEWRsU82FJOyIBNTitP3AvqkbkhOCN/wNc5Fp70ZnphHeTp4anC3Z5bmhMblTG
uuyFvIsT+EbmIwL6jJjee6qDpr3Xd4c4OIvRIlTShBXXet8inudQNY3hc8mxluzx
AJp69+BPOXy/PX9DSc1uTfbDMv1zyHXx1d/GJnGBL6F9XgB0iqxkXaUYmLYsWTIZ
0ESP0hIUGSLBGQWdBdENCr3sgrdp/z1GxO52je6tYDjvGvraYD/DSifDDpN7baSY
tYPNlPuH5MJbrLaTxYRzVUUS3VD6CkD2fo6Cuyap+uwClR8Q1ZUQR0aBAuB7wPEC
pcRPo+bJ0jB1IPrbvXcKCpSJzlZnhl1Qj1lb4c6/0A1A95zQ47Ui/8p9JOlp6k8S
N10cXCdg2y7ZgOD8nm74z24bxHIs/G/b8zaAuuprDhcoQ4FapmLYgBwd9+cf0wDC
g7bSmJP3XkRnbwaN8j5EyrE2+GGSz7LhLVT13XLYhpIXZXTIrvuU1ovIns8dCzRR
zR0vrK+9O7Zw6UN03g3wZizKWi0yBZcI4pLaDaS5su3OXUvdrZcyBNaXPsGtvBKT
5blbGAnpiIVhI2bbN9Ri3Yn5W+qOy7Otm/uaU4Dumyj6BPMnnn7gi3dxSbBcZHR7
X/TUeVBj84WbuRWWE6vGozu/O3zWIY3itQta5bEBVOJTQkUbzgeZmhhmc+60cBMQ
Az4k2JX/GDTSOVvX/56PPA2HJUbi/lZGY8OvKgdvajeRG3cNq+QF7zjUdKlpnGCV
/SZW4e1rntT8smCfWf39qZf9qHXYSmWESjs6mE5BoyTOU2IK51UTRp0kUqh7xw96
9pvlcFuxZUYeRoLrknL+eRIo9GcYPwPUsvDP0w+a5k4wg6IBZFOssifBH4ueBVcJ
1qOt/v13zgXN170x58qThQctYXqXCwkPsum3tCXGNA+lXRT2JQHb78N0BTag8zc3
hQHbkVx7yljEFk0NkFQEpAhXZQ6j1Er6HmkeS2iO+dcgREBz8YlDXBKZoOOATppY
NANHwheJQiFH0yDPXoaVLsOSRnMUceh6v7TPSU5uiceS4IDaf6og1Qgqq8LrqLSD
idwU4pHj6N6D5+9c5nu/poXx0dilOGE2pW6KEBytU19hjDHjz3G1qqwEr+ale4Qs
tyNwr/QcOGxlCb3aRbBHfJTYgkZOVxJgICkiTJyEjuSt1eX8gsyK+ugBFk2EOC4f
al4WsmX5u49/7mbVSnFvb7IzYkpnT+6zwY/F+543d6ZROBHX/FXhd3JMDJC0/srC
bsyXMqu86Dr32B42ooju/o8SnGcasGBMUIvB0FKEbRSqyieYQ2RqrBrAg3wCF0NV
qxueTU7PXaNOCmsI59hbLLGyUqwm7fREfwdwWSy8W6IiWtRV9SJoJzGk0n2rUgnJ
5Cp4jDz4zAZrXOPgA3FVJp33rYpeJxNYxKQNLhVWAAyY9SHXYZt8FYamDcGpaTN2
yFTozK3TEMg+5h5MiilY2SG5ArVcRmcy9oX6ggAeAQFDvZIKY5FleiS+ShwfWjVW
LXj8UVNp4lwQPYEaV9ffKB6go/wKyhDozGPS1Al0WlyrKnn1AweU1DAUacNPgDS3
tIxYKRPelyt6CBc5xbjjP05F2Adb1tlh1V0av/sDprJgZ/UGmbX5RBKLUC4Ch7Xc
MUF/ugkhD1AmRDpci/9avJiFEJ7KdnFF9gNz66sedlXGqW7noCpeitwyKiZ5T4cn
76nnG0PnBGcSSNVptIfGnJt2mc3zT4m+J6xWAggn+SLTXvyZG1Eq1FNV9XPnF4fs
PnkCfukWLXeXJMmg0yLY7ZJI00DbbChk7p60Admyd3p0KKg1A/iWkKem0Nrg3rva
4iPVv7CQ2pB00bi7FJYV9GIMCbLK+sQEekyCrTNoIy1uBVrIbd9jjTXYMODQXGmi
XtucuH8zsG4dq0e3aT0vYrN58r5+hwaXvM1Dstq/qrcx4ybaP/AMM6gkXT5612D8
spvHB3UPmn2l71ZC3s3dOn5DjySmZPGA4dXyKJamBEbb474JY60COptzSXTzeLGg
uMq3CC0GBMOqYMjJxJJuLeFKIOFj0AMblU20tUdBKYDV5YVNhsDzCDRkICBerXaR
kfIAlEgVc0APuou8etZ8iO/oIuMPgRhJtntKucqv8dnUoF2EiC0DJDO+L0vdwsHD
gB3br07y1vCHvN0IYbPzn3+V7ZGIK4i9yBn6k/29iJ4YWYD1JeHjUQRJSQQ75/7b
1RFZd5XEXQW2SpaQ9rmw9wfd6KsP5AQho/4NHWSyeZ6CUpBQSeISs1aARCg0k9ND
JGVAe3CU3hov5QtbQflrL++317a9MLJhyftf5F+DJI8rGfyKZHglMJCgm9D64KRA
W3dKgEe7gizbPIXEBmmOQZVpksUiJy3Bv6yeEc8A9IWuWAaGAxuDjNr7IBD3ojOu
l6G8GOfwwMJ/n86u0nDJnr/F5i3NZr+W/UghaupgzGZFWz0yuW2ZkUlUKtabknNW
x1iqvBoBDf1ZOaX7IchP8MbZFz0NxTwT7ptcZfCK1ODbSGe0mbQv8PhK0/jgXxTm
/u31JlR2HbmxUO0NXYrKaDeMVKvZdqunTnQAnDFKhCRnJjYcl0KYfkhzcPMiw7ly
k+yztaEHj2eZDiZyR7QzeiOW04hC3bbko3hwM0YHzHauhb6/GGfyuWpzR+0RHdB0
8erNXGGWT5vY6gYSoeHyx6Ep7zmQy3KKrPmaUfUxGT05+aUAtcxYPLLUH5A8kGJH
ke1rmH7dwtopElYXOMv+St4NJK5OeagYb096Ow5X5z0BPadDIyGsRtTK/BpaNnP2
3XQnZqSQyh3aJUoXsB+MF6lymVmK7xqrP+htlY0RVYRALr+Ua7bMfU24Tq8/9WhV
0acoDcrd2RiuRGJ6yIu1HXnUcYOjxCb6xlGnwYOFkaKA9GOQIKyoCt9rIE//OguX
lRxiuY9e+l9dhWcV0xbaPp7DS+lohU5VVFmjTEgw9MvrsebLWYinTICEKL6u0P15
z0ZEtCx6pKwsFJeHk2HiHVhBn7qiIdpM9G606uccTNT/zqXpAHwwsKRSw+8n32Tv
F+pC/ZMBDLZAwdR69/b+/FqcwGvHtDkq0UcKTQk6WRnZQx7ggOp9YlehF3faFcUg
npLWg1d0bSrNV3B0qgSWMqAYdIzwsOg1WDJbmltTNLQbC2NlnUqNS9ulpgAbGuwY
2rOsTC40e/3kgV4Hoag72eu0/O8ZBPATmVe+sOhyoYHL6b9B46QhYxe8WH4cYm6t
USxXoX9SjbSIlPf9QttIEAv4vnMCGZq8V5cT6uTVNqMpN3LDpAhePzGf5KZgjyaN
d2qvpfHoIfj/NblspErbS13yd32GkcG0yk8PEtH+Ej+H2rfl6PNtru2IWwL3hmNl
YpwKt1XjpIIHwzPEoCTxHKGWbf4ei/Hgoh0+pvb2VaPuRxfy5T8kR3oWKiOz3FF8
kE1rFJ30BA8I+hZi0FzIkfu3uBRS0Se6E8LUjD8DMNwTZt3jtOJAKP/fz0YPWr42
lAENYm0CVvxMZag896CbUIMuKf3W+zcSuvfOtxZgT7ZUzjZm6W3QKAYR7gG9Ra0G
d6hMv4BqXxAttYdk71osM8g8CBLVljjYIlyK3GyKkGi0oEPmJGo+gJGc218wjj+c
Kn8y2G/tgSYw0QTob+vjGidkI6d6RDo80DVzSA0yycI2SXYWKXRs4qgyyH7ogRbv
wnr0HK4IY1GnqlBJkdPYy3FSj06W1kA1y7BOqxX43xi7hI5A0cfnT9yYR0cgA546
mOkkNQ8kaQ7JcmGCbkHymS9isCny+5kZZiT5NO3jYlS4jc+k796owYvoIZf1KgCk
atQAIBGaqZi4dLbZ1xRu3dhOBIPmB8MADUEPO3XimMOvSVU4nKxsZRvE937A9L3O
xKdDVLnJPtlm5Hsa/lYs7bdzZ6gYnJu1lHCsC9Tuzm1M7XV51f7kQ6wCbf6dT+ph
BdFJBdlQW/NQeTDJlpQdYXpEtzbQ8ifYmvEX2EQ40ZbudHPEqOlsrOVg8Uze/pwm
EYTUIsf2DwB//HMrFi+uBDInWPlC71xfepeAw6n+TF+3rZgH2wDX59FkamEwJZb/
VkRa+1cLDPdVJXYoTugjDddffZ2HDME4BtWyGdQu5dUiqKJpnJPT6+W09UPoIVQ5
QUG/PlGhdNGst7KHHmLdSVgUyGUtlKUJopNUM7GsSqYlXh4Wop2OoPxNbiLIn65z
KJmUGiAwogy6oPlasY4utoOSmt6ykign+5Nd26CAcSUXFsScAI4SS0FqjU0XpM4G
dBamAOAtNnYeJkKRlIaKqSZvaY+qGGUnM47JYdi7fJbRvej+PJLU7LAVLZOGGHIr
W+uGNnCRwk+fuwRY+cRjtVnn50WHbnu/XsrTS/3+3TZxCc3cTsdWmHngsRbptrPG
izIfY3NkRSMzMsDZOxmuCX1uP2gUroBNUp99JPGMdlqiMTts/HdFuEG0TMiQ5pAX
YZNb0nWOA3/fKNnceOsTVxKe9zs/LULUiE+fmpT5ftNwkfVmsqvxKtLvG09fnSZ5
R0kEb3IFJZq2T0Fggo3BAt+qxQCiTrX7ZkDhfBbOEVd39iyPKL8lwcocB4WCrQRs
QoPtEcfaShSoCTQdgjAI+4QIBwyhCoDJj3OYyagJ//nCwg7BkXsIJbbJhURJztOx
gXtqn/Htw+0duIMLPOM9zYqJbo1d8iA0Ze9ZIlQmmEX2rQX1TYbxoRPQi3pbv6wc
04QAnYp/my+hwu997SnXQu7+ACvGgFK2hiioEMIQ7CIvKT7CYAz+tJ2eSHVlUJsu
O3L6wTWjfVHu1BKcNFZhoe7/f4v0mIKSlEZnCsn+nfJwtu3qyKU5YerhiL1PHVe4
gyE92k7dTUCuXFbj5bO+Ho7hcl0uDvqKrnCNiXEGq5uIm3lezlmJqfTMsZIbuR8F
f79MDV7bjXlUTX63XvNuS2yk8UNCWRPXetr0eJYjAeH4UsmxOMlIasEKgx5X34zM
E2RblUHRCjYJcR+0Pc1KxI2DXz6o2FNDydS8hBZSG/UMxkSgT/SDnNlDSxEU3KOB
elfhpAAhitJQODf9B3DjN7Yd1bjrXfBxsis6GIae060p9/CBNDNkdOGiHVi1MLvo
wgL02H5tPEHcKGRLY92lqPDJzgHSJtJsWSY2U5JRgIn1jgcRbgaGJVP5VURshMh9
AeUu35FTCaIivDvxkZXg9z6Z4Whj8d9CVgTtmENS6ya/0yS17Mirnh3b7lexwghP
TqSMkIO+7+hjWBeEe3Xb5Ec3IVQ3Wag+ZtoDMRwm+CXwoFgdnUeq+9TxFw9EPS7X
/T4Cyr3Q0PO09vMgOTDcahdluSidDWzD1V4l9whmnVoNHsurRKmjcAkfC1MrvY3W
0SitwZ1DFK3Om19nto6D3+4DNlbqtUTvqxPOS4cpXlBQXnwBsLupiSOMnfTxIuzV
N9kH1XOall+pHBvLNr/MkYURUmbTlfJOdkLiTPbQpIY2NoCF6myM9cwd+36DCez5
86g7ovBBID9zMYt4O7hnNjghDPaTt73lNN0TFRbHNIqPGeb+BIIn4/LAmWjIFvIP
Xrom2jP8QhAwQH6CDvKDzOeRs4cuApkqzLmZktf66EJUGFOtgeVJYsGYQ8K1OAlu
eCVNeoslSbEOFlptrTKDNQSZFJEgG19IqVqH8e19b7zBwMjodzNFNmK3zq0JIb1c
Qg9HGUA+a2cPW6cPvBaojs3v93NDuXtCwAVGgQX9DqKNRP9t6TkaBmgeVu2x/g2f
MV9iwQBRu1dgukms9sGbc+QblVeW/Eg9kV7QEHWf2rQqgqNhm/kV+bGztPkwyXi5
gwxXOhUOpTjoMibilSs2GjYh55rqAgpOL9R8xuWZZTbjl8sdEPvFM+CsWxhezAF8
DoTqOqBCPd/cPpvMJbLeorgC5LjEt6uIZ3xyPI3wvEvFrPOFPPeC03gga6NR7oPm
SsUY/hyrDtFYHOEV1ocGDnZ6AEPbnLWwIyA/q4XCoq/JI9dNgv/kWzLfuUoB//h2
B0/Z0SiPhmxfx5Lt25tb9eZP5+iwBkwI/q0wELiF+yK8Vpv15WPVbCwc5HeTXMbS
SWaVtjmpEQZ8Jb8xl0tTipfVCwBj+UevBdGCrAYwGkQvOIr4+0tD9lMDu/VlHZ8Z
aOLV35QigZ67VpylsPHG06vGRD20UtlSmCzSqNwJFjIJi0B7FfeaZa6pXY6sMUL8
MIrANdvJEijsLwjkOobenvhxWwvXE99v+55S5tq/eTIljzDp3Nx6x8K+diFyakqX
VCD6okHHlRx+1vzaodCjJe/c6ZRNNo0aZuhKwa/C0u8VpPzf5B41oBOMO/D6pjl7
H3PoQCPKeaJ+s5S18P2jSNhQdO3+Y7LrnewCPsBXL6YSs1OngRYCKS9LM4WY0NGx
cPRgPjTSKLrU14nuQpddzQLTRs162/9B5LNmPxSe3Eh/puW8Aq4Ri0wh8nlikx24
QEV0D+ExZS3nuDxovM/3of2Vf1S6X7FJTMjxDr+BkYzdch59L/08ZX4s9PWRoaIv
MfZVP1EyoMnAQNSROpxHxeE0dZytCMIy0oM8wyj6QfoFa43A+FzA+b6nRXgjWMO/
3tYITcpULIqX4e+JSlmluEC+icbeKl/JXQoCWs9TMwncXhogTyI5dledyxNdOWdT
76W3wQ5fPx4PyHXltfP4F8TWvTPTA7foFEY4KX+izscf4PYodYdhRVmdStz9oC5T
MbLuPD/Gx/PS0QJhBwbc6o2h7cCo7yQpaA3I9Rq5gjGVynGBik9SHOyT7d832Opg
sA/n16R5nOkBL1emwP0gg8uyhjudI8xS7jTKEMJEmUKduw0jxNTiq/Z9mEUDs4+3
/jN6wPMP5rMJvFB/WtHWiMhXLKR9PcBXZNlN9k+ZjIuwzPp30tBbMbkdIjQjl2Sa
P1cdOpPtDBpBifLHwZ5MFXKhYFbhA8AG7e9oeJS2vYFxoH/AS7oL90q0xwKmcyzt
o4pPUojCDWLnjigx75N44HgpXYZSwWCGeoVeMy7c4ctwlbaUbt/n7Jjv5xQ20rfD
5AD4snCGil1fYX9bQGp0+zccy3aVbQcQPP/vK3AkaEfqTsgffLJ7dtln8UvheTB9
jGVTcKfBP084Cu+dVdgE/t87KvkPKjS8cnRxjAm79x8p2iBRgQqlRmUFMbge+Uxd
azASwdXQXJ0Qk7HF1KzngHIEq21lclmtPf/Tb96gPQnfr5cD28A0tIpYWESvJA7l
Hor5xbZtNnDLFZLOtTqyPV0jznJB8DrnmwBOUHKMJvuHtTy2c4ZU/hdwJCtPLqeH
XlKTNar0xUNd/zQle1gsugB+J7q844Sl1iGlo6pz47PGpbI95EsmD4GPv6uQSrjj
il3n/d1LOdJ40LhmoP1eJ2RQLfv1QWGTzZmoAdSq/R4xpIXuYCKo2z/hVmyVqQP7
hc0pm9KQsRdKVPpvxqamN0XcoiF9zx3X7lspdA8wHlUXdZXvlqN8QW4a0jevb7b5
svKM54g3OmFVacd4S94V/Y0fPT9XfmqTxm8t61Nkb2ypfPkRBt3wzyxKdSc/ezzf
tDTLtIQiPPBj8y3p/6qM2qnClTtYfQDK2Mh29uDvRMT+rSNyte8OHAH0D8PpCI3B
wGZPE/qrid47+T99nuGRX7ElGCoiz+6N+RUZksHZCOGUGncR16cxknYkSOu8sxXh
5cQIBMKuSeiSfHhBgnDYRVou4iopq/j+l/1CFNeIoNVJSHW5bsNaKlAO+xRMRJxv
LZtWwdcbA6j8cRhUxcZFU+0wFPRQIEUmjGX75DUse10qmD+j4cx/75qIrKKMUWuA
R1cocSSthkSuN7MK4/zLBtypA2zXIpP1cpHrenInOaIxi9fubHkv4MymmHhWBwvD
71PzQN24n+q4tx+AmvCjtnE9wXLFtVzV6vx+f/ibOy0=
`protect end_protected