`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23952 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
hRRAlfE1xLfeNfywbrz10OtvJixhnWeYVQCxik57Bc922p07VrPKDp1Q3tvEuDXC
TLAC+7GpauO2e3rkOYILKAhWwDIN0zXGnU/1T2wDxApECnsdX4R/8oS7nwixszOu
efZTkV8iFpcvagSK2cDsaD0K77q+jfgNs0sIY6JKd9kghuw1UQETZ7lcH2uBZ24/
kwd4AY5ln8S6FmUG2/7DNtjh89F6bmNwTCwsoriwzFiFECAgMPFtgl47UNlZZdv5
c2xopdstC9A1VflHME+cEqkESV3Z/dTSrkQNS9dpSQ+e26MlfqS3iJaRAyMUoL2P
XMjQTIQZgX2Pmi9k5c9rz1zgGU5reXSc99rrU9+wusmU43G6tSwd0A/VI1k3nbDp
csXzIpPyz9O+89tLWfZX7KTWJkEVDo7gGgo9j/70JeVANFxQBVlogegpiwsi9r18
1ixHWGSvPIWMMVCUo6aDj3hAHnBaFnn7QjkZnsQwlhdFWXhUW3BUoQZuQfTVTS0C
cy0120bJP17x6Zn/pWPzW0gojehIf9xPS/yBrZ6jun7Uz6/ZHiJVb2098+dJUmbf
+B47KMf3DmwYDz/dk/fGWXOJWK8ByV0gxvGTYzyk7MI4CE25e8Ax44jTG3qcspEi
Kx36wXBnzZXB9EMaHqO88j0ynGH4kaKTMnN0+Smb84jnwnDQd6sk3E84Zv2B76MO
xP3cqDpqXjsZO6qe/DPz2Zde1O+eO07ORvLYL5oxOoBchaoLSiyDF/u/tJ8G2nam
f30rAz3zUGmAGbXomHsUGcX19xCpAKOv2DVxm8lw+4AwuShC93AJaZwxzpa3dx9s
HCZz60T/c//ohownvmK/gYpKCS0T+4XL/5YNheIWKiy0Wt6xd3dO3eKoZL33YRTy
Kqpq9PFOkhahhkx40ydyErZbJxVumhIKmh5K/cBm6wijtjm59nLI68eUoAyjNIbb
QU6Ci5ARI28Lsny0It2oDLpiuMajrBdVpzOYto2HYIq7m1piDux8wL10PdTUAX/R
biQsIRGtk4hH7Dio0yVaXLIyF2yEQfz40UAw9PKlNslec5XMDqn+1bySmFt3cMCJ
jBdAvE5OmOaidjhj41nWXMWthQI7nHN8saWfZsoGDsAfgibMjqRHlCc309/MwpjZ
1pACuh07guL9GatZdoHqYba0H5UJibihRj/L5NYIjIJJTHFu/VwjgQHO8Iwj+14n
6FZTrh/Y7t7OUuLkrAX+RfKaCmhpuWviaKlkqUAZHZobTsWT79s7dEOFMmuD/Ccf
0xgWN3X83fQkqrKyPFQ7VuzwDtNDwFYFK5CsUzedimoF+eE2WNGity+knIjTn034
ILmvXlslbylmzvfiTBeqjb0IaEZGXsKcGTDGjJMru5F/OGVjvGG/knSVqWTQbjjw
iwX01ClgXAlqK6itScRuHjtATmx+Pgl1CFTepI6r4n6eYp8p5FdIUVqH+gvgW2Ge
lYjaqueoUQkIY4ZvGKwpLGIQIRHqWrCyj0us53rkkh1gYDzAQBpOowiZ8Ox9m7kN
g+cHy3UABHvtI+54u/2pyIZ5XgEu2yZGoHSMs3c+w1YdQTxvzUUEFXZkhSl+0KL1
VqRhs/B/u9trJZ651V4efHvJDAz58vt8BH4SZMQP0dEqEbtg7hzsefS9Q2qKn2qb
1jfL580jwR3NwoIVbW5WtayfKsWmxg8WzUq2HGQYamGWGd+M2ccBo9vhUbJDIIFK
xJOBQvOLvGn38pMwoxkx9NcPJ6Hp/bHARBcDOHowsTX6kp+nccVpvj82efJgOSwg
uaiPBH5sxLB2QoddpCrZK34MgBWuU2FBBXqd2h9e4qNtbBh6gwSLzs+ww9exTBnE
JQFr4l+oI5kqqeh71PnsUZnvANMOaN3cpLj/3WEY55S2/OBOFLyGDlTwYH8FWrJJ
pl0S+JzHakc8TZcT/FQ7MLAYIXzE/zUA3rdSgG0ZBwk3tyu/G5otJuEX2s0hRD4d
LsRUxZhuMUDcDdr/c2c/Y2TYjDiiDi/yr+QGuoQAETgkqVq3EpukFn54gcVl2Fea
xW+MGAkQlFCBr8fsIBnWiXGxOco0GH1ro82dGRHjiwj6zFgHrz+Mw1N1lGC7GEMm
6VFBLGqjLvdRQKz+34skwzTN6fAoDDYvlOYaH18+c3KHolMouchx6/Pi5r4JYX6c
EZs35AyzCsRJKOFQPbrjGkH69q9bbdmEvMbJySQZAN9+KaL12RRX/bR81ccLMiA3
DBqMiAC0JHz325iW1Syqd9w7HdR+KmDQYe+NKCEggytlR3EvAN7HoeDYKjuH7wkk
0e5BRSsujARMelDbAzNcSSukMd91BKAZQccTvLeP3+HsK8obz45n5lbb8VPKos6m
44wT9QPnxZirVYjFIMT8NlorYeAR2230VvXxTXsWkPkmuFEkN/CbQrIZDNW+r4Zq
ScmVcw6CPkTH2WriyvPG0Fi5PjJNr1K+uCBZR8/gwsTVBw3t7ZXeyz19ZQnbKkLR
Mn3Dk1pFYh7dnBuJ4SIMj10izacvIjNb3I8VA4z5uUp3wnjoPuFk+1kJSF6ucG9S
ZbMkXbwjJJzMCBu1kPuZKiKrkjdqcPiKNjIBeinOP8ginOd2G5C67m6IVHfWOwgi
gCa3ztqJm/m5qOQu6VLQKKwr35BPMnRj9b/xCCCurdQXn1n/oFAt/A2NI5WUyCPu
nzD45Vohl9eZ9Fjr3zx+Xlp1SwFweZyL/GRLHkQKzDscjjrpczRuy1AjjMM7zmp/
1lJA1lpVcsIpzKcnQf2TZ/u5zEvoElhZ+DQ0HjkwP48Zz0knce5mpKbgafT90qlO
dpPKlIs6F8QuaEiAzCcdhCmMFB+W1PVJhqc4i6coGg6kjumeuGDSqELGudEgzqAF
h5PStPq503FNB1A8KUzsGqJEoQtoQ9uUlwSRO40AfcxfX0qARgbAf1NNdfSSUSKx
Lgy/vhKona2TErtNeiZ5bhh9hoMtkl0GS727UTZl+vJkn3fxmET8agbHhYABqmAm
T1nyIRE0MqvMSIAz0PCZFrnmx9a+CuiT/daCwxl2Fz2M658o3eNyjdoHl8rzz76H
PWMa4HZLAbwK2IpMrGBj6qtNGQ2l4oMATJVVvOznlQeeIU7y2C1BOqxitJGFT939
BBwYLEBWxHJbqCESuWSHELOPQm/xQKNifRL8sNf3yv3XfR/4QEIl6Ejboed6I9tf
hkdv9Org3YuJC5zMWt6XRIE9VdEqr0Upr3jk+Abk7VQSLUF8YJc3gXWrc/4mA646
3+rpSJLit2WFHoz8JWDYXxmxWoKD5eHtw2cvIsd8O0e2paeoieEeDceVfuxLmMiY
mxy6ysQbf1v1p+5Ra6oXWKxFBmPL2C1qWm3g4Q8XxJiaeqeIrHpbRViN2SVqTSjS
XIyo04Z9fByCm9cmqQztfiDFUOyE709Cv9lcgwgg9IKTjwV6tIfMKDcuEsPi0c0y
PkuRXTlUwBn9Bjuo/Yr3O0dC0NHDT47dBoTXfA3sZ7FvCCuanPrnlogKENIUGMC2
YUYde8Pe/9Z9j6+jsoTNQ8flYvVt8Kab8bFVCt2bv/tJANB+HdCqXtyIfK80haln
Z9KgPlshEgUwOV7ZccGzmlW8p/6MLXmK6AKJ7bbbwUYbQQb8Gdp9DdO7/wZuu9a6
o+8ObdkAAEXAhkC7o6uCJGnOW++VDoch7tHVS8WyZ7UxvlDL8T/dhh3rQivSD/jZ
i8Vo7KjTqW0+9JeAUdvsaU0cW+lpZA/H1kb160cagaihnnNUeElbjKrrGVIj2Gk1
WX9Lx29u1m4qNn6aowLzMY3Rh7BbcGVfwt7BRh64gqBWil1Wtb+imoMGdcpluQR/
FFWPChLxUZkvE5uHIPXt8ebPy5EtoBUOk3dxVIFXnhyk1VZc3iicnRzWA87jXrvc
d2FRSRyHfo2C8DbPt0KiaN2jjOq4LPUFxfVW/HP237zWVSerFImuwjm65sEa3Njw
PXWCHXBqFvufI98qtHY/rYTUDOVWZk/3Be+vE+ToGC1+YnADAPp82TcGRV7jWQyu
qR0LTuF+D9rrKicPdzPIQBrZ1csZPe8yg+LF/41qvdXBw7yFiioC0Bch/xkrq2Nr
6lpVXiIH1krmDr11wXJo2dHON5xJXHVEc+a8sB0C2n33pA3B0m3YLeTvZH8Gb05i
6fMFS02VHVtEypUgtx9zCcneBQ9z4Fqcuv40VDwoYlBFSB1JL4Mv3hJm1Ou3JP6t
C7WZ+xtqxBPw9ub6reAuWCvZ98MCWLSEkm1s0+3lqV8bHebyf5JzjJ+Q3vCTpag3
Alxm5YeZdLH+JB1HVtxUI2GI6ZBMKL53S5OPshluo3Lp8k1ks6cr3IV4swF5o/Lb
Mh1+C/cg+vD4zTalkvNOVWJQwNL4MZbEJ2IkFECH30407K2p2BiSjmKaJPPVHmFa
J2dHsM7ObvM4uFGumOHVmP3PKXFbRaZBM/yEB203iJh/1xI8ttioJv8nsw59LROQ
7fWyOut0CNslC4f7rYIniRSOYpj/mLWLMDgnpogUNqjfSyluuj+wKLj0uSy1WZ4/
MHFumgMblFDF7gzZhpFLyUJlIgbrrdqfsVKqf7x+v+yiF7nvjTIMJBxJejKhec3H
jgqfLcRwvyJQKip/tnYj3V1bmQZ/gRcUFX+NrSY3LF4pY2aQpVzztIv4m4BIw52G
6t/W8nuQdflgCF9AiyV6kUcLR0KBb3Q4kd+VA+y4yQCoXiXKVJmQrn6YWP8aRPB+
vq4PYUjcxe1EBclrWH5Dq/noKbytXCUfMik3Yp/ZI+Qx80StT+WdfObept6DKjap
hItiBjWdJM2NdDS+v5BNvi2RejoT4XznzQELbu0cEjWaWsKwjPLN2zvEnfaq0x4p
2I2+nhjVe1+/McrjciU81gAIGjH53/+DegfJ2vn8/lY5+HBpv1p5FS5oow3hkUpq
nsVAp6x6CabkRiE8an4QbfJ/MJZjb2SIIZcRPfUXLABFtzjSjGFhkBxtxrmVZWvb
ezy6QBq9nwjpYw3KpIOCCEVZyeX6Z8fx+qRBaPFK52/v5DGz9EvGCtl49zzPjWjC
+RCSvjWyweONn0AF9G9MYTQPAlzvXrhDZXOwJQXJd0KUmpDHC8SstwY8My+j7HLV
605KA2QDBx1JdktrMBu2wofzy7Xe6apf0QiEsEgrbqOsXQDS1oPdFhQnXlLvTRRC
/vGjAKg4yFMGh5phkMp/hlfOIG+v9JeVSwKz99Vwu216XzokJStrnOYQEKGCSM0R
8xLnZ6/4cEFcPZipPHAOEHn0OFD2VvqaO3M/CqDzTlzNbtn2sbCFJnmW0/oCPlFZ
IdEqcwwmMVjVwWZTJt8Ll4+mhdvB13qfIwcmJ1BvOMIy2hzvTpP4TO/g2GxyY5cu
fIKuzF74tZaoDX8gV36yyluYJlA4+7fAeKca8ImOwWKLgJduW2o+GAJrwBCGaiOA
OHzhEw6Hp91k6OSSYhDqvikHjYRVWDU61QS6BkoxvsQUxT4Yy1+/ILIA+BIaqF1V
wyuzz5PoVeOMZvY34+3XdVw6S2N2EE477XBvax6z6Oh3khR8T2CGsCunHYAnfFMQ
x39BsCvKJ7bnmC1yABH1dkrnvImjkaR08K8EcCNiBZRBjOzPTSG4dAghymg0EQsu
eEy+HeYxNqERTMH7Hwp9T246EQ3AmN4itspZ+bJAOBgSL2gJr2w06QfzHKolANSc
eSUYGyFGvCj++GReqvZdI7BkgwvLFL8FuCv2hxNSHo6RGf18agvVST2UyMz4JBhq
vnLar85OzDrwHrK7tcFvZrbY77TRd2n7F4sLM85c2bfKZYeqnqL2ab/CBsKQFEwc
ANEj5TgNeakUNZRwlrUSBtMn8b/LlRk5drqF/OX9av/wnvrdF9454P1ccntVpJji
Wk26y1VesiFDbzW/QXnAg1NAV6tc3rhu+J8//zDwVj8XEiRy2zTz5JyqUxQWD78L
FNXFqwjWB15E2gb6gtEFVCALTOumHkfq5+WdTCPdzLXFEsvM3ZPHPWAhZf8BAEbZ
7w/e0Wl+Fa78DNQwOJ1ap2/QcXNj7pgvOhq9HIJnfRvfrHievQwKk5cCrSYDHXjd
rnLGUZOYcz4xsEveEzBvU56mMKqC4W3rY3jIv1xt2+J3Dp0gBCOOyaTwR12JHZYh
sVElLvd9cpLhrB+CCamnBGwWs+oqA7Y2lNkUCc7Clz2rLV8kKAlWnfPN1mfNUe00
y/nkI2YpR1ovOv6hNzVUWggXzP2/Ng+2cp9t5sWpxUfGECiUGoOWJrTKZJvMs36l
nxqE2jgsVsdtyat7cxG4XJ39XvuRzyjH3F5Wkl3jgkzSrlp5Nk3VaSFjhql71Pna
myEUvzKPbJ17Cu+G6/AHAYdNBOF3xTCJ+QnhvbwSMTq3NMdW3D1n0U/VJkSiWa7f
rHStOe4qQJDpmWAbPPQI7gHFRQOcpkMKdY61JXgOCYlj4maYMPfxYX2KYoATawXw
IR3ulVfluhfVnvi/muWJw1lEgEh5oMUeKbrgHcPsNhUW7V91oDoOU9yVqZ60KZcG
0Rtw6ednEoBRK7gExtQjt3ESQ4Ax3WKxuwQ2wSuSGOEDXW0jDVVilwdXYt3HWcas
yp5rspSge548sPLUnCkt776cR4fQJfNkqrCEyR7wgxu5JOCSvfUZs74vWFvHngFa
nX+JNUBr+oET52p2oXJsM++ridSUfcHpmic/29165FxEUxhxhgFwtqmNTosFD8D/
S57SfA3shgqXuoPwLQjvuNcqiX5Pxu1uD8tQqajBKFCsgiEVOZ2Xza1D3VesH2TW
V3eBSUP0VubYr8DIJ/UpOHbksJzUEFTGGupFn2sQ8PicGuaj8RM5sEJ/sNJaShPz
9YGTJCdaMPzeIFI2w/amAf39K8MqDIdiLEgZaSwiYgWj0+sFA1T/uuoLHCUfUCsV
3RKIMAH7H9CycTKMlxuiysNhxgnGctSGJzseJuCuSfLHGOpepP3OUEUNGC3bs4jU
3HEw2wKrx+S/RAhC9U/Ucv8O1/CPWlCrhYrRwC8cYWUHCTXl//EY3U6YZ2EgHLor
SWJDicuy1uX5vmUrRp7nBQdoHd/7UQIBL5AYpBL2aDXJ2RTJogbcOXfeP5dK5+m3
ZjWCLbXTBgZYKJuebyPC1Oj56FWZb+mh2QKmCP2j3HUFHNAlu13CN3S/Fbm60Esl
4Dejk0EL2CZpl0Ngnmbw4Bf9wCmB4e/8/XCDc7yKjPzMDAJPqbPE63yKrbrwYJYS
b3eWEY1up3jLth1y7K1yuarUpiPxbTgBLU485wqleEG7gFMnjNXkaxCX7tns45vx
2xLomf6JSBeY4G2xhINU2c4dhJO8NXypZPR0pl3QjETAaCoyJYPOTtQ157RxNCdw
inll0fFZcvOkjM5l+8AYJj20kCfpBRcqdj1RmxWf81GnmX7JBq8BxB3gue5oZpLv
YGpIdcygOqkMpZMlJlPX6WAYgZFdADztuNpPmhhvxupcC1IsR8U7r27idtu4xg4L
xOUNeRlAolFEwN31GBy0RW++d+MN5ZfIUKWMzlBZbfonjTvxlENXItfn9dtFRi64
lYcFBPb9sEuOSvNqjBOA3RYUXO1LghcBC4wTQOA8lhgKNNM86/nys6T1YcBccdAw
QknFubIQ/GPOL/v/TDbV9lKAlsM8NpGPw+dxTfEqh6Jksj5KsAsUbI7XsOS/FbvC
FQ4P+WXTB4xj66qEjM4zLrnC2RDA0hNGwPyIkn+gm1JksvPNePfpOX2G3rNsOIEl
r7zWfIW6VSo79KglLjok49nyJ06h0BNnMr8kHMO7bLjMfsU8Avr4zipBpsvwrjUH
eyk0rg7MtrRANZBAGbh/QCwa4xViiMTcVtqfq/zHY84F0+tnyGoXpFuQUhh1wXc5
5HqfQwBk6pKnlr72uM0zVrlwKuhliBLTyyVnvZsgzkxMNgcT/zoxCaPG0M2APV3k
llNqKMP1bD1+OyyUAk+KV7knEusuNh38v3C+6sEG8rwZ2RVVzwz+m7FstimY8eoo
KKCbgpoPfAIlrzuBTcEPObf0zu3UGMvq+E0dE86LpJ6dIzGCK7sGG1GIt2fIY6tC
bQHgW7mZF5tfhc9aDYI+8O+1KVlYEsHZxkV/VpjtMZ5NETidgz3ChnLep/WFlMEL
Z7XNMEXCdhNOaQHMjfpu8eVkqLTdSi23uwsiQ31lX7tduwJ4OOIskpF9o6YO3sE/
9PwESTYMqtoDNZyZZzptQeT0ABzzFQg+zf4Mr+hLr4crfdEQ3uE81WOTZZiCjYSH
CorePCcyvvP/lqiGKekOhd6aeSsj5pe4TF/91mys1zys1BI9rINJZ8yyNiLVjtSt
BQBCkWVkyqf6IZ2w18Wtz5zIoMa8u4TYMWEvZBk4lFdjNAJwrVlg4w1W/5hHS58P
1b386q+6wC6YSUUsDczEL2JhK2cN84uRJEwQExSfRNcm8BzvGKBpIf6U1RHj473N
Mvkm98povtGyzk3nx5kmATBBiqEHuBO3lgrHH0/UpmmigrW/tyQTFAu4Nu5eYKLF
Tfvom7AoikIogszN+/3FI+JR86vhhO9V1v8FZyhLFQZ64HQwj4QEwCEHPeHJQaiO
kT/IZQ1wPcLYGyn4yIE+u2kH5qxmDR1CodEJT/lpcJCy4tWP9xgo4/nwlZYGzw5S
UbitZ+6G4KtaQvm52ZpPeHSgJxdsBUuYu8SAPLj+GE30cieN04ktHyIgOmZEMFVs
rLrT/GoWoL6MrpVYuvdonNBRWOpPXsHmoSKZQyhthy0BK1sZIqT2s61I0Yqhnu6f
cQADQH6NAn+DEOGzT0J/eXPO/lOlio6Dr6nTXSA9XWDNyfzXfdaVFQ9HGB/z8WkX
oz2qtZWeoe+IGY2tNZ0dJDKa708vqC0g6tbxY6lSnFZLA8zbx4TLmsMoUVrL2BFB
vcOw+eKXMMfKcaX+CuInAmCSUYYCLEk/NozlVkVV4nd+66Q4xmUc83Zhw7LF9F3C
wX0zi8iOQl//HwYN9dp7cwGGxpQWH3S+HiH6COhDxg6F8mqzhCgu5whddMeMPc4P
sehj4E44N0cPAQzh+5IAJJGEeSOEkgkuHI2+pclF2yayqLeOCS7Bi+1wJQ5fc3zn
zRka98gfbQT5sWtDUb6Zd+Ug7nDEECQWOcH8knoUiJ91pVEjsdOo8vx4FgGSUPet
Ma0mFVN0iXr1sd38PM2H5YCMUzCuOpr/9XSfYy51Qnm4JyrBuPgcVd1mMClXVHEQ
PKDtvsCbPQOVh7CwVA5QIVkfFRB4wD8WeUH7Snq4o6fXBbDUcjdHReMWLxp9WwHB
yp5dQXqXdq+ZJh3qBtAThTutesYcPy7xp68WFUJOoV++xlYGFT/xejieFiBxbqA+
sryD1/id+whWKE+L69KBZcwYzd6E+Ie1qzFxvhpfcT8Q65ve8CmSibxSjQTHvP7f
wgo2UkHN7r9ZP0vtzPvd32LBLl5muB+nbC3AvhbhG7Xp1ltqgshffGI5nRezCGow
iNEekYfZmK4IdehWqIIVJwTIellVW1wFBW17ca49BFM/DwiVygyLpzEw4eE3uKRL
1vgEHwmzy0HOSFCz25FQ+5lCk/WrjwxEcHcFkkKISPIcmpxKViYcyJey8+fYtBjU
on5wh+8Eqe4Zj4mxj2KKWETxQsaPbA5XBhX07lHo9OFEW/v7iNn00hvtSGokcjK/
b0v5CE+SPJIZ5b8y4doMqN1u2qhcl4ViHpwuDQtV0Z3WpqKPr2Q6cKkfWa1dYuxU
W8EnHsLJF7ytO+C5oR59rLmxEI69gN1ZZV2qK5zZqQd6ThA80QYY0f5Q+M7jOZzU
vR8gFmIzxxHxdvTbwa8HO+tiZ2ighDv52BCYAYIjKFpTlEK1nN9LnTuWkE/Dal1c
QqY4dZsjqqII+/4rCa24+q1nm+pFfA5XqygF+z+tru3aqcmAEzD37uuQMdyEuAND
JAo9H33QpzlAZvmEk5Z1xMmbsvNnE3bNu3nsIkEDEUndjOj4ncQCASqEpqgGL4Vx
kmzRxHmipubXAqkLVYqUi7jbJ7N/7L27FKYA3tNcS0mmSnWEX4uUACY2aZdIN1Pj
Q+KYNiFCRjwZZlGBags3r/J9SE64OntMTi6lcIAqEyuOVsq6JMC4NANPi60LUw5D
zqk2Y9vnaUoN2NTOBMl94xocX6mA5v6i88M5Y/j5bcrGQXyk6aiYgYTTyYv1wZ/3
lGxMfrZvwfeu92WKP+Ma8XMqJB0rG9fh0GImc57XHLk7xIOdgVwfxQZeLcd9kLxX
y6Ae2iODoSkGS+NMh192TU/cd2Kuoxgz0hWrhc7OL7uaWZ2TaavsHKUetAz/k3H0
DECl5x9KR1EwzeWwUjOapMEeXx0kbsnsEga7b1m2wC9YMsFmjCNS9i1G+xUAT9WS
qNkLLpVVcyO7IrCKsc3lkWGt7VprtUstPVvItdBU1IHYC0AfRCZfRLanQX3uRCIw
yML5N4B48XhT50AWvl2OPkn+Wxuuh3W4vBd2lWzDxQx7Gf/BnN5cOfqVkcVsiMnZ
gonTfAzOzNpyz+VmzI5p4XDhk29Fopv/VxMcKvXf4CY2okbgyYE298PLY1fp3CGP
3rss6e49en+Wpks14mPkkn7v+j2uxUp0BJ2717hTwlz7xD3FXW0wFekW5ILxPrxX
/IP0wEhoqPYK+oi/LqD42AojwH+sNFpsYFSwkIQxcMAS8HgTZycgFnS9oNxY21wP
6rf+E1Yj7skwbw/oQ9LBVKvi+yFGhymx/+9Hzt0LlZpoVNotg9iW7+dByZgrd3tu
6i5MBLml5H6YaSjD+bQugf7ghV89juD/P6LNo+fGroXRJ6Pxz4YTsDH9cZL02TtW
lVUjzT+ABeLXV8ji64OmHSJs4STq5Ue8bHK3vRkvoWehDjQYdQm6MUknnbbKYpey
HAef8GmZHIJ6DJs+HJMUMcIG2vi6jqrDFhOjqQbagCdqYWjGJsUAzUFAHQfm2+mI
R+NW2n1fKAIf4AtVrABcrG+RsUbh9fqG7iU8Yo8pzhOOvs6TVhqRbLX81FNkOks+
1fUh7PWd2jvKPNJCZ/EtwhTdoMqrdfTidE1AB1SC6NdRjCkMxEo9XvVRaFFQJS2/
GHp684tUohh0+K0HvtUBV1o92ckuMRol3WBKRrcXVn7303Pmb8GwO88GBfj/tTgX
NpVRwwB7H5Txrz6oi0zOqefLU6ylMwjia7ltbazxQ6D+QSDegldxkNXm7BGCtU32
6kVWcGmm2y2WwMdvVvjroLkMGP1v39RNSYVbUZ2BjBO+rk2qtIUi7baz4FNUUf+d
VqAzfnexKZ0RvMuZktaZJUswjMRifoVYJ2vw+gJLyXXOulK/2MIdBWeohwWthBv+
IFwBn/V3/Jsi7Z6/tyjWqeIy7w6XX01SVCDGv8sdWclD40rsgSraqzMZYag1usrq
RdC8d2WODV4YCtJc+K2mp3a21cGOlqjJuzzImilDoVpLvnP7NXUBts0qdF+Gm9wD
HjdM25rkzXdK57NLtlcX5q8pVS+y3ZhX+oxKG32WYyTc2eFaCAkBi5Lyadd8B+oT
74DMwHSmoGILPeDcQSQVJa1MPTtDLwhEVtSHj5hXWoeI2+zD7NAPJjQBseUgmOpS
HzNxFDoSKluF2tOP2RMIlN6kEQgCW9YMCQBtx3FZ6tKJLOb8HG3gAu+51AVX4JFL
kI4o46D+fWBTNC65YTTJMMwJgctU8YWRxnr3Cf0yYD6LjIWHl/ol6eInlLBHBGT+
EVZ2s+rs/8j9bQF/U8IE64SneEN6KQCxxPcLR6RgIrU+wOddQrp2L97KZ2WNcy7B
VWRphGewawJd6Iddh1T9i8KKZEtIrCzUXO9JAM3c59NF3E1RUm2dKgnXqinACinc
j/j37F44U1GRzbJF2hHXdBRHfmrWCyZBEkwfyxy3xpZEqT40Fj4rzAANNpomeUSg
+VYVAUvfyU0mwtIkO/mWBQD2T/gSxRKJSSAlipvl1Ly7jR/yWqoV2sXkFGb3YCJD
Q6+cL1hm1oyq+gkCtTiDTL6wgm1aQ90NkkX92guoSccuosejqBjxaHhvelUU0EN6
cdt3J8aKq5nLGHUk2HYaZ4PED1YIAET5FIcIkvVpDQocHheg+iZdUFJ4K68bKNC/
z3BfJgIdEGRgcCiAtRzQORjiizNEUrMnpWC41Wy+Y2bGIA1SszqfA96vPCzrhQ9Z
HDBA/NOB2vTBAorClUrdRp8yioYY52Blp4f1mvv2cvG+oA52eza69U+wUP8M/1FO
9hhsRcata3vnhVAoN/YlI54+lgQxVDxPc4swZx9zORggWQq2dyflEIQbQZuCoBDi
FpRC/k7Af2mePRGZopYotCd+ncStszPnJYGHyANN3mbM8ACJPRz0R9ENWNhDRvcQ
pkLRj/nQU2VHSLp8vNCg8ZhIuCniDcMkAz3FeIRLlO9U4r43CAZV6am4u4WfhTIZ
6uASXYBSRTb9HZgrxITvnncUAUfOsQz+hFoQZY0XkgMM9CS8aKK8eZB1v7Tq0rFn
tg4/r1eistqxqJmqT3wehf63Qex+/kG861gLPTauHGTSn6plchZY8GbQBflhPhe9
43SC08iiA+Dp/Lz5qXBaES3zRm9q9638CBY3SoTxvaDVbw7MuTfNJUvaD1z88zB6
5P9HyR954esVFuK8aQNU8ja5dRnEqJ1n4nhFBR4NF74GmPPA155Wb+UCCrPbxpMH
XTxS81d1JuhPeats4lzMVTzzUdFjoPYieoApPMbIegGgr9A1qndnQXeJHNYh5+xc
ExJSGwVVFrs9xPVIKtFXAM7/IekTAHBkMD5W85IrjnM/MqoOBJevcsiX1mtdBW5K
Xs5yGzBMy1uhDuDlJgTaiyYFZDrHUejc6ZEE4JsYA02HtSUbZbRvuFeG1mDHsaoy
uPiTUs0vOWDCWpWkoU3iM63VWE9t5tihQSHcx0ZRYAjii8Sh2mD5KMAAck/j89rk
yYOSWW2XPtGT+v8njDrFQTFn0Zs/998+HOYxzuMP2VX1/A/UOc6NWNHb5yXlBv9H
cwT5rsI+M8l73LhrCHypdjYBF0mtkXkEn1cVku8+hHXJ32Nub0ABPb9DKYHDpITL
jZpTYoYM0CvwcnJDUjR2bAd5cFWNvjM7ZOsJczHlbY+l1HMwg87aGs9KBgMPUIRz
wMaMNX9eoMQbIe54Gws7UcyHSxnDdl9LwjlZnFuk34pEAKF2ifb/ZL0QMpEKEX3Z
Ld1h3MvbLV0YjE4vOtfuH4+ZINQ5gOfTpdkHsWNr/YeuGCqoWMrcwbZl3FozscYF
F7PD24eJA2kJNP3tgS5GzcD3E728i9UOBk93s+dNKirxZpdgm/sZ/vmGbomDo4yU
hP9lsfjePWlXG4Y6PdLd4b9w43m5N1lumrOko26OcANI0MTymmvfkX3+Pwq4Rz7M
OWkoSZt0E2jFLPJVFx6XlQPrk9/I6e9e1MxGH+ioKn/6hvq9ZE0WL+TZxK1fAMMI
bre+fXJI7dUc7DsCV3nH7yIL5JWciL1f3P0+7SrDjZlKLB9zSXbHQxatSD5rFV3q
hfXx2ylFDHzpLlOBjwiYboPo3H9TJY2/vuDlsT7f3OnPWSPel492A0Z7OvrX4+1X
NKRmVUF9oqCv1ZTlneCrmF8qKRnU7XjTLW8+LwXJgq7M7nM/jy6Y+qs9ke1DCU9w
U478QPW5HXVe+onNnVo/mq26ovjhXNazyIwKlmFqTd7IRxdpNSt9y2U1CjjhTXe6
WCNBheaHHTjCUfvlbnuapOH4sXKVVvdGmvPtf/QLpXI1aaywGvn8IBidW1UtxBJo
yd8rYRPqPjjQcEQ/ELdtNIMUsi+2MVd06OojHU1hwKWcpIcrPl7etWdum6mFc75x
r0cbgbm5hWW6b/60IqZOPbzc7P7tcBdd2SkPYI3ujhe4jzEj+SuUIKLUPG8Jd6uG
GBC2JlfX89nVfAznpy0N8rp1Mpkf4VPuZmHy51QGtxbxTXUkkpJ/btcCHp+XfgVC
VKAOmM+Zw7/ecJnAZY7ot9Y8I4E2ztqnhhR6Mw/ENWcev987kwakZUa+o1/E1L2U
icXnE9UQj+BCkuWYbDq/saFlTG4x+E0Hu/L/G0wrbo2aEzbu3x72dHO/SdCvujFD
nWxQ9ISi7xIIo5G9XZ6qaL6mXWxwl0ktwwghdZBY4voFLRveeSx3+A8/S1vfJHLw
XvOk3EpqAFKBuK5Dq9tSrkhsMSW/ri78Yiz04GwDQ7UgQXbZLOEMgzkP2AhgSAnC
8wsiXJwAF2JuJErhjsx390AzfrcIFZhGNUdPdUNfRFRnbJyzY6vVtuP8zDUQJxpn
TL2wQuSro2o/aU5AhLE6lZ0eDALSbPFlaVQn7OoRhHVohGMPfDkrJuuwf6Kl94hE
rmTbaKIX/NprCdmnmi+SqeV6Gf/oBdNu/JRduOq+riuhZSeKM+EMRKyL3NC3NYO7
yuRRmuhUptLmpfGER3LTTeNpRhE+bmgpKqkR53okB3SbVWwnFSvBqoLoHodp/kCP
kuPVOlYAvy0Vi4mHakv9foibqHCbg5WI7EPAXYk4z8Ot/zxTJvtQPjjDDIg6UxOD
DBAWx47YuG87m3io5aoWHbZtg75oYmZJj5iPDI4SOkYXRptxiWwSp436wjaKH15h
y4ktUiqWlM3I977RVroFbET/sDUlJVsU0R9MAbRle3Q4hswF8gDIYxPAadUGQCuR
rOx3SHzW+ocy5gI+ru+pGA3Ir+AT3obhSnn4TAzhOfm1oLWrbvni2EKdl+DwXR7n
gTQjTJ6I8mx3cGJ+8ozSsvMIhJsi0JVPdZi8l3UWaN1HwnT+FNFSbskJiF3unxMC
2fBvkN1QUrK9ki9BPWsDasNWY8EERd13aNttcqLl1W78AdtQ2j676sOvObErFXWQ
4KlOD8fSFqmgfi2/yPiXtdJwCRPIs8ZrsA4gwrZHOpcdA/6tmHesyhXZM3MsNSuw
2lk25dUqOECNhTLXUODn/k93xkzTdtbRLN/33YRbMxZO6CSFZcrUhCcPALe8Zkj7
0Pho9JQy23V0z1eKc9E8wtDxUFFy7WdadRUywNuxbmoCD4h0+ag97WOprw6FkKO+
CYRMlUXqRNYXIZlsSKxDEcCb5iCFuXT7fjOaJ0NYQnD44sEJM/Q3m6BnGAlqRifQ
3XW4kLo/N6z5YtCUgmD6l78qtg1KyRF+1tHD1uW1GGJaEr4Cw4Itz/cTlOU4iQ8F
6QUagXr2yanX+/appoFKgIBVfYj8O186XOVCWAS9TeaQwOgcScK/NdEdYrZo2Ali
jyJ12YWrYBRIvFdpfQwWLSzFt2OhkFgyOGAXshgnSlhFs1/gYuUNYL9pulItx10a
bOS/H/jcD+y7k53Kj2kzwAq12C/vDouCXpHlXYC5T3pY9q9f0Gu+htfTrZWpFFRe
68BifmxSrBXNPmLd7hA6MCi24EPRrO9+eZHyOgPvOUNsdQI9eYJ75ssey/98Xfsi
NqBWbXyorcqP+/Jl/bVglrY0WbDpZR3xlvGQow4Hq+p8X7IhHbZs9wC08KCWYwvo
y0t7Tf+CF+UgbTdDuhR+P/6VAVuQ3L1NkpKV3EUJ+SiU2egob6oX0irohKoGPaGU
4uPdW6q4oTL61OH2GmCOcvBfpNQavBrxue3crheJuaWSIU59rHZ8f8ombUdUUO6R
Tp5Dfztw4I7sHD7Oce37Wjo1JZmHAexuBsgi76ViN6Kpmtk4w3DrSHyw7svb0wvY
iABlDnfcLwRmNy8E3ECcH4MnYOsvcWapjs8vJritObc+ytIUCfjYBefothr02nXr
eRlyP553FX3jRek7N7ucdmVbt7/sWAlDJkpIzX2rSzw++s8Nj1CB2yqb50Q6gjgA
tzF6F/FKuR5wumyC6byQLvzLrD1cV+7lp7cGOv7WHeOW/mFf0HS4UGxCLPcS05Xm
KC45aN2Y6dSYZlXdGTE2G4TLQ57M2d7ug1lLA7dESHoZFtuBE4/Kd3ivapuy2Q3K
2T36ZC0+LaMPoCGLMfyZcI2Z9PBFRR4aZBy5c9aHbGbc8njuwJyQun+PE+FBt4aY
XCFSCva5vgHYnepD6VviY5uiZDqBcde2EnrEzNpfRljMNtTuX6t4ygnAti0arWxT
pCDE0HZi2XCfsO/VuqbLaWhfCiqmReMSdm/MEB9OA+j/ahSESn7WEIMs7DGRR6aX
cCfLaxYAe7hzXReHiPlMM+0p7guHYa/V7CzETIZWclngTODXogfmukwNjfeBdood
g1hbdKbHDK1CdgL0gMj/sfyhvtx6+p94YejAIrvHADhGk1NdTon2h74U8ar2X1w4
58t0y0W78BSV6qGESop/kSl5KYozsI0kvDsvOxYTYbOHayZzvTDlA60IsNBXspO+
N96r794H3Gbq7hgz6+1uaVmvaGdMM0Q8UUgjFlWtlWWMdggwLP4BOe4pEtQIKa6O
FYeDwm+knLjgsEs6/34/rByKk6HLR+Ke2n4w2AcI98UuVySsUvxlnhADiSG9Dn0y
HKqiQ5PUrcBmhJY6M+0JkBdoMR4oyc49J4joZhRELL4GYi2k2XSsmWJOR4SpFchX
91NEWOzpWAr5VF3G/zQeD42lpxyVcxADtnbRPFNcIUb6twu3jeoj4XY/FW3rWcu8
vmSyBLCSpbYuomo66jqWVrFlusWZQ43Io1YTzGr3x+Vq3dEPjgJ24lmbCfHOb3Z1
ae/8CZEQPgv8jIKJWkMvkmkVGeYaCT0ds2ZPOnpMP1/7G7Z1EFOrxf5CivsOa4nz
SdteVmuCfoQ2FSIPCB6mQQiCr2lzOyaSkqepTrSlDhAyghvvMhTKbZRn6BaLpZeg
Nrh5JnFgWAiZ2Uk11UA2MRItfh62T2+H5ubByqjyWJSkMMVWMZO/4U3lqtMs9vzS
2FtTyoN6Cjc1LdRtw4PVv8JcFi34DEdbNUaQRLxQK44thoVRtfy0qEH26bChoFP1
QV36lgRE0j54hQqwaQ4Lat2W1UmsgqPtJt0nv+VezbNFdR4P+t663TrcTKwLfwuK
aV/cu3tLUwgB2U/g1AUTNMAdnLlKzfvFuNSVz90DsAhf05BT4Z/hXw7zYGpm2eIb
B0lqceOfn0XeU3Tkvg1gfYF3AkXxEwrnWNUBcRIWGNHfQq8YVjVTUkLCx5uxz/hk
WjX2r1QEQfJrMeCWZsO69vHjZBDAWxZzJXCvs4OV0A5NfHX6G0Rf/SaBY4EDeBPy
2HHrLplsciS4AhiFuH8dzvWQmnn1XhUhEvrm5bZQCj5Ll49F6oTYgppbcjWFPgel
XbvEtCp38YjSky8CoIxBfThGn/E/ZBTbGua3EfPV9D8dUlYuUOcBmzV0TfFTKcD+
kB/c03ueOxO8Sg2ZRRrz1La91PqIEKs+YDUO8ZltbPdGKIs13VZ09kkqXobdB9vk
q3Ms9kCY5NJ0Ld3GPw4SFvAXcaWTAmtiTjQ7jg0EYBOuzLkJZtDDShUAwaJxUHfe
FMbvqFIU/Ir3U0OZaQQdCmhGYzkTLd5mrfpx2BhluCUb6fZJ3L8sWZkGU8FrWxqM
0DnsqlrqHWdI+GY2QLna4XgLCZen3t7H3aDhzBr0cYKTaDg4H2mQOAAcUmZo1OWV
6vUsZnPJdSZ6UQfeWSGymdMOYZjAjN7lg+70niouQq9hd1bOpgInOy4Azh4y2LVP
t9ofNSaJwQqRHKXecF89f+AMgLVGFLxxJK08FfItAi6sokA5HQY9rkGUWs5sQBRi
GmF1iJjxpvb2WNNjLUsxtN5bPV52cSgu7JDZWmamD6KaLQ7nC/QVsvXenhiFBDVN
qAAH6+JIuWQ9f2hDzXHIOa0Of0QVzlPfu/I5eRXQBLlGRvTYgRP7rmbmUK81hcAg
rF7KVCmnO+3Lu8bVUVJ5C1mH5dEEIo3z2N9I6pVJQzhQALpOPjjyKX9NT2p/ZGjy
ZVQEzNJk+GgHE8l3R3VBIobtA8boYWS+SfQJzdeBquYDiWzxE++OoQtvcRIqzX4A
4myydn9vujuL1VZSjV2hbPaq6kmBBaV3VXUa5KLYyU9PvhQdm953IK3RJq+HfWhW
2U9wG/KyZGYwWU/BIHomQMZgp3WNqj56JWKE6h9tBna3tMIs/Rn8IC/5ZvebNDrW
optGIksin0A0KjM3MhO/2L/uj16GRkFD3cAl6Owqs6GUOyTLKMbU2keDze0X/DEe
ipe6Zjb7iQCwlE4vy2V3eJvprMxNqcTUrVPZQNqGWoGv26pZKsTx79As8zsU1Ypa
hHyzD7vSQep+EIIvpclsbp4Ytx1zC262QoinM1jaOd+OXi6CbQEajzzNBzF5AQSn
akd4wMUoMWOzxlJpP8pwMx6lakDCffp83xmLHyMUxZfx5J5l3bIaSY2mXCGEFJ8r
pJDYmshX5ZunX0opb22yF3epFm6dNcHtBDuzFG7xjXXmzCcXy6xGdHergSVHDaoO
qLjS7246FqcWwoGl7TbW2CUxTQ+xMceo4YqkzQk+KRtpJCgpuGQ6FmU6VdxGXZy/
OKGy27zvvxHqBLXHefLNH0oLZBU207ztQ6DNhCTvZw7jIEnEalYq0ACigtNAlb3Z
WNRki6e/uXBSY63dWEKfX4Q8rBYPNzMaL8fkLAzfKlUbAEcItLK52FkHnjf5/f8L
T8cFunQpilItOjohmdR4/sVxX9SOYvs3FS6riC9j8kuyCBp/eUg41Kv6xSVI4Ofz
OPSNy8bd/cAOs0eTVlIlADcWtnApZRjSJsGn8f+HqzfaIkmiUFWI7wLZ14zza1lb
96zFD6Voe+8YyW/gthRXCuF0lt0nqeOu/a+IF1Yh3ovHN2w6QoyalFKjVuAjWgio
zUzPoKQoXqqZEeIhXVCcB8eu1lUfbwSWOW6hpip1iL+JxGcFuviqM6qg/OPaw6fa
Xin4/R5bD6ptoC3xj9Uk4Lp+OkclvvP7XUuiqedMywzOVVU0OHzxBJPTPjNBLX7n
veXwzBzNLurCcZfQtuCApICPOF4HP8N3ZGYQkbLDtbMfa/MXhcUioU++IpjEW0IA
Y+RyS6gaAty61ZxchLmr8ET9mLBYUkVNm64sMABVe44o+cJwMBO30RMK0kMGU6X8
KXPFhYmA898WDe0FnJHQ4dDmor/1nx7v4sCKH11USuJeVWa0HpbjIiuLkyOm0IPM
RwntIUpni1I56vTwfuC9W4wF4MJTtKdOHXMNv5r5P69PnRlJ5N7n2L6tJguL/m7s
ccuIePk73OcwBkE1gsbB3lc1/YvCakDypZn9HzN4x+orljmg8uGuX5Ov4ASkd32I
bnlsADDl+YH662sUUt3tBTSKBPuUzaFD6dWsmLPTcFsOUa/6G+UDX2r4RO8n2nNL
urd4TAKdKBZtmKK3hP7D80wAQgD28cw93MqW6Q/HS8UBYoaSC1LjD7msuV2T0H53
cJ5f8fP+U7cSca+om7hD7GJbmnscqAXz/fKAZkMK+vgBDCO/ss9FESyzEcTLUvmq
d1UwK6XjMr9eXCUWDbQzrPt9ZfTGOgV6ofYTfLPF8DTAGZSBD/NdwoekdT0e/ZWA
WEoNO9phZaxOAnML469Xj5L0k+IgesOl1jePGHgj0/0NkXZORxIH6cPupucLQ6TM
nKzqL1dmDlD7mUCYcTb0PH8kHcTgtY120SlTQUUuHD3pp7UjZstotcfNH1cV/UU6
ppKXO4zrxkW8BCiGvgZUDilbGyD6WHzW6Yw5HgUywqZ9xLlkQpzUrxnKJvhtdlhE
8snNttFkfmRvjeUhDape+Qo9eeLXltZc0hDpcTAO1vTqiDfikSIcab9/McgMQuTb
iMaTlD4LMmZil7BO2ZIplJAjmaeXAdZ5Aa2pqEfxwQS83LUGk1JIlrmBWd1GldXu
qCi3emsd+B7kwzobEP7yWninATQFpd8rlmm51PkvWNKN7Idm4B8oOimrLENp+TdO
D3S8EBDo41XxBnCrlR6wMq4XI0RCGlEOKDvKDNrWW0fxD4J2MWJUc9IxSCAVKaAf
udmEROUmDNLiNhYusHggmsqxDHTiOFYs/yCuOM4QXdAVaLBBXl9iH/sMFnQF/fpi
RR5yoEvN8xE/D3TWik734on+MwlTZVvpJdDd6VG3X7noPCMfdHU0p4ouTY6tBton
asezbm3Kgh0KWFfggq8tMEQMYksYO0Bpya53i3T8sZ1xjnj3O+GHaq94zqzx7K7A
/Cv5WcSv/Hj+wLJndtq4anJxvTIKQPD+Q9AauOe8SRqLIBcDbzsjpwMtlwON9KUR
FWOTadagqYqgLskL7OAytKbsSS6H5C1nf1G7By4v7D+nEZVQbjelEU3AuXnNt1ys
M1v8uIuCyhfHmzESPyc7+2G0hOlDwhIKE5l9jvk8Vz3wr5bY4Bi5smvrg3ib1+Lt
Ur/hiPBmGanN3ZiULLyoqS3fC2oBx+vETdGaIlg1ILIU3i8WX5cdJ0A5iElFSw3h
CagGBKygG5zmhZwOAl2zFGp7LmFQaIqrr7e15Wt6nshU7BLZOzSq3lp31kfif0Pd
D2oLHvxBiemrnIUsLjkAchSfEBr47sjOM7kuVyvyQuCNU9qt0yENIoUx4HF5ldUP
MRZWZrUc6MDorE1/HLsex6nfCHZ6/mwKtbDrx9f0WvAtaYYb/9GIw1sdHjLb+FsH
vwiRPmiup9bmUZdp2lCzPejQs3wyoqSS6AVJjm3xIu5a9aY6l57apSayq87qMUIs
6Q0v0q6sziigW+yGsbYwSmG/pn5UBsH2bRcAfhCRuCdWsip9L6Mc0fEXe9xeEZlP
UIy7SCjrUlP/HGoXKC169pGq5VbBSJUlJTlBEKyaqtxwJQPIoiuRG8oxDp4P/dZR
fMKL5a7TfOYAH10X8S2UsQPH0tefYsSzsQhCud524kuuwDaQynIY8ElrgvCQ0Fqj
iXuEgmAGQ4CXuNcncuYnE4mrc0SZy4sW01DKN5GTmfi4UkSQti64LPq5bMZcbJO0
UbPPFkBkQ+XmD77a6H8C43iLl1A6HcyXvjHb0bbSdbEFjTca6k8Oqto/p/1k4/S4
yJhZLC9gQM7l28Tjrf5XbzlQ0B0aWSD/+uB+psJ28TxCwd30rYTWZ41Ua1hjhctb
lIH/ByfJivywBjW80OuFQk9HH0x+R61DLT58d8cCCGqzY5t2EVScdkan3KwHZ7hD
bFw7xnwmsgUreBGVFqdqftBjGUdFI2IvqFHB5oOUAP2w01+J54FAIHjka12PvaDs
82vjrW0PCumZ/3qdfZ3FCLEe2IGam+dODunR/KEhNFjJkox4zkkkpf/CjAgW5Xng
O8141Dv2SKhNmz+FRTRXYZCdP+AF1w4bTWNeUUQPdVbRnb39L0KR/Hn2XxL1gfz4
YUO074RKWVnWDCIy0kevr0YZu3O9FSVpHdH8jc26AUwV2rIGYwpEom7Wh/v3dMsT
oWUx3LPL6FwH+zEMQ39hkfogVyDbblWagqBsCwMUqy7ZbMgbq6VULWkASH8ovTQu
eLyK71wWaZWW7kkeEOp89ZDC9Ct0k4tWYk2o91zLClbflcAZ8eAvIhmowFSHDzyv
dtCxZbdE6Wj6hzwDxpmwq0N4O76CqQFc9WtYet9h5cOGHxUf8ZBueGTiNReEB/Af
RcaANDainWIIlKCg7MiY2ZmwiEci6gC6YUbnWAxvURREVN+EE9tUuain7tOfL6BE
3NTKaMO2XNSH0JRURP15RK1HsFd7DcKECuaqFYlO5kkvoN/gd+E3lrgcMat5tMBo
rxmyrLXRm5wLfYZNX1mmYa8QksgYxqBH8vfChe1tOxcqXJiNAHmOD2lrphXbtpE8
6eEkcdf5zUYzNsNbV04NWR/QdVB+GBdkL63fPRmFdqt+VS1xyE55uSICcjwOJTE1
9yv+hs/xzltafEBIMDUw7ElECZtjg1E4NFlU8Xz0jVfmxd1L1ve6ax2c+9OUVRa/
xJLLmhzyX7IElUd4lJM3mfNkp4QLugq7RyY7Jb9tm93dOKsVNTJx6Tgt7CLF6rRK
YQg4sxjIGZmHh7wr6XZEXAMLRV7PBxqm29VvvfUWYSxxZOQfLZ9a4eDYLZOJ1j0A
I/di/9b+fH0tkCyY/A73dEMYbvKSp3hMqSX2U9N6FRysnarF6z+f9yYo0CbCe6Ih
i1jJvkKa2YPzC4eGlq6SkSAKAgnIjyrNsnflC7CZQzyqmFnblXDimfCJsreJJAOm
MLceGV90TrJT2nXGkJvr4cLMOqHUtkIdmez8klu+GRSSWw462nJsuoWsyld/GPhf
7FLA69TZNKsqXB7OPpPahEnZZyk802mhlaI8yXDLJV188M0+PsUhLcnS/ZPXpzeD
/+iKVQ+XveFPyFkt7LPhnA2ILIJw5Cnd3vDdCn+uSlSFLpw/cLftX0Cdm6A4pJ5Y
XCp29jt6RFr/EF+0wX33QJLNt3NNmkSNcKiBFZGcrkgQviuiFrBd4SrycrRshGpU
x+wXMZtbjMM1v3PvazBdh867jHOdz/YNuUZptBpzLD95FMCr8AQUoKh/M/Y6iwrc
TN42Vy6+Y0GZ5whfiflhqI8EHVAPi4H5ADrvjsFZdl/o0WyV9gB2l4M1x5aoxw/i
D6GJ+vfyVFJWGDFg8F349bvpfG8PbT8ju0UzVUvkXUFGy28ip/Sz99NqaidTnU5H
JilWZGHiSDqnLbREF4ZCDktMETeI5EVmWnDkZcfj+FZYHqD5X0spM/2Vk1Bk9pde
uFZIpwwRtxgrU/oRXm6A0UA/VlXRfJ+mUkkdMMAmZaRNkzVoI07T3+IgDiL5MQp2
F4mBgyKPmrsJ3ZO2xKoDZpapkE2NhBJyZv5NdqFyJCBFW60o+ug2B3xRWw2MQGcd
OrUMGU2tUrax2TEYgWYxphS3ZhF9JPqBvtIu1srA2PGXFqCgDqBviS5EPSMEBt19
jM/+PPh/mRuit5gGiMYcQh20/i9AGUgqKD7RVCmfyEEM+KU2HsUlStpg1hxKZrmx
E0P43YTWAPwOYSWuwLbpSOsLr2tdJUAQqjGIAKSazAVNlhSYV5fPBxM2NtpyF+j/
BuBv4NFCBXP7qEv3fgHMQ7kA6uqWQIY85R25fUPxgbcYsgrc42sL8PRneQjjwar8
uvbRnt+H1OX9Q+snNpey1QsBo+QAjtigdwbRdt85OJPFTNzbViwil7RVb0YnBBiS
C99O9OidsIyC1uWvsqrI+da7nLThZ5lOsIWeazyvfmzCljPfxp/pWq2oihxDdlyD
Xc+xj+w3VMk0PFTDBKlQrdrmQpF5wropEMqoOsBBn/jLjGgb5AFMdr/sJi/0Ov9t
zjqmAUCA4RE+u32F7fyYng0vSh5Chbtf5JmzTNyCx1wRSnDhXDX76fzmxnmYIcOh
CqcEBPbDeM08SwLb71SRD9RqWmjO6o+LmgobMycbbf8X3T4RPMRE2z98b9JwuQg1
mXRU+7ol0Lvd4uTpqC4xGRtw6Y206GWanK/oR4QFT1wTdB9147WxOblJxZ7abteT
cwqFBCOXDfMLFVBs4flywdaSlmBXV2BdPnrcuMv3HH7aYWDv/P+LpSkDY9OdNlxJ
V2yqhNoHD7QdnvmSqmf/OdHOQalY7ndjgmNlWOiSldPR+EhbD0eRQbGJrGYJAFWv
0b/UbnKG7Hwg2g2GrNKuOqojJIP8PQ/b++DSQxt9BUriqPO0twO4UtTnk8pekTFS
Nwtz0GV1I+vUC+sfFKTmNfwQFZQ2lMiWjFrUhJkQO9G7hGc2Rhs1ga4YR+t0m8Re
YvDQA44B2UR4tkHSGfh4Qnix6iWzDBrjqemkNqApU2hqxdjhzJOUCH4llVg2sNTg
4GFPHyeGQaEQdrgfAxoF5Ejcswfo6XEHriHt2Zh/ByR07UC1pgg3YsxaFhq26rPQ
Aq8XmbaGpj1x1YS7orx8kmsMOEaNSXhcoAUhZBvEWeJj/weNxtEFg9RssQ8LiW78
lNM8Ywr1XuQj1vbeG3dKBJ1tOybkuVrkgKuexeH3uGvkAqdi8xLfMsupoeVbTsxq
rccjo2J+DElFpEDmhbdG9yvZzNuGS6S2oxjasdPAjkoQ7WsQHRg97ztAoAsrtKj9
MhmpPyM8BbjZMMAShn6MzJiVf79YBihMzDtinBULEb5wCykVQjjB3uS4yNFiLEIk
N8IgR97UY4ePH4eum0dVGw3gcv8Lx3o/inKPKUSFdvVxjnlmAhpEDsdBCmRB2KYZ
avjlZ65AaqEbNSitNcHKDbddvzfPxQSyUYhX18/k57KtkE7SA8sNiqSWISQE0KPA
auhzzuL3trc71EfYFPbc9NXqGjhkO/zSY4q8fV3axQTzsRRmpNf8Lt/T4bxWp2bO
r2VWCaeGHP/Z2qhf3lkEy0H9e8yGCt6ucsbR+GH7W70EXj+EvTyJ1Tsdl2SIypOL
ZwuFCg//ne7mzhjWbDpwQYDi6b6G/dRkBN8hxo8s+aqIa8o83w7GBlMLGvAiCiEr
ZyUNcokXtPCRobTSBXSgbaBfD2oPVuVSicJibaMg+UU2mfn2PP+Q8e5lBS76auDP
Lu4zswWGtC+NhXZRVwIH3hpo/F/Qb6g6OuJu2/j1iBPMBnqsa4EzEyxYk1SY/V2z
wLv4TBYQGR5lN5e+dOTsmWDVSjSEeTnlFNRUOwu4K/fJ/96WpCSyGeK3l9bD8XJy
Y/1Z7qNBlVp3g51cBdNMgrrYOiEEQesDWrjk5qlWHApTWzd+pfudhFusngpmf6Wm
41c3twJdXFQT8ztfom/dGLTGEfTzZ/uN7PA5yPpU1vMrb4FLqc81lyprp7FusPcI
GAptRh5oFITCIIvxQwqf6xLaAQ/wBK6cciheGxlYC+Ste8awf6ZdgyhQ80TxdAM2
uCPK83c++loIsnC+Jfw4jysX2rjbgoRgVy4WpMFZOoAYHp0sFMS82oLLcp7axORS
rdPiTChN7uFOH9NJw4dM914wN9OgqKBFKplJR+te/Q6UyJ6DxeH8X+AKzy9idZCc
/Uj0ygUfZtT1hswBDtZTkkmUa90XwVtvzqtTtACMNMsC+u8ot5V+K8yRm/c6g23P
uMfY/JdHgQCymS7WzYNpx8QRakKzz5E8oYDFj60+EDR2mi+eEKGbY+xPybZgjssK
AODj7VMNWTrVS2QnVecXEAbD9f3qcEaARrFF1PP5x9izZRctxCUnDILSoyNsmRab
s8UXP0Tp7AYrk4Eau0tycOUve5lNkGoaCp6ePf5ETr3TW2qAUmPwr7bXpOQIMSPp
bcsa9Fmqxrwj4/JBlxtwZjlhyoGl9eLOpns7ngVbOj+lZcL9ZGJI9rrXV2zZhqX/
Sm49PPbVjVbnoQ39omqVdOQn3iTa9S29iwmiEpHUNhNsXLS1vT5E5EwJgCNJtelT
H0NLxtXjBEE87meb7cK7SBp9hKOZE5TkxJyqn8+ZUOjSqzoyOzdjVwBSuvqFxIYQ
JXvgBxC1VcnIy8Xf8v4EAAvjnlrlqZZYJQf5lP3aSi2oPiAV5SRRnL0n0A+Vh9uA
UCX9jEv3BjXNMg90Xy4ArtDARW+77qryAYt4LPHY0NLhdwlR0/0GRbqc3XPl/TPd
F9HqLTbGOhnzMVbaOM7mQb0OZdwParWDS1Oh4DTKqBGexyAoEQPwgc09V8/8/Uur
KJIL98lo5x4l/Du2Zp9J02CLXPkURx59+zDR+CIutgGNDRd204qGR8yp2H56To8G
foeXF5JCIRs0wZwg5zsKU3sMlCdx2VN8z1/Z5fv0wb23Q6VpA6Ue6Ccu9uRmBtuS
Wf/hav6Op5jI5UYNn12WvrbQKSDxcUrGUtsHQsHF2yArIUcaS3gI1dtfozpWbRSR
MMEWpTRO7ts410e0DOBX4ri6W8KkbR0UEVI9IdnjyEshsVRbPpVB+hyQZ9r28ZLF
sKatjrZzRXGEUAD92RCD9c62778GWicuOqBY55bBvzT7GrrpdlN7hb6SZgr6qnCZ
Erk4UxUwSBVwiCEFfFrPMIW9XcwnPjakjz6jh9+pIvTVxjUzcHRKxdHBveQAtaHZ
LGcIYs9tWA+9B5smXN9/QiEWpeUYc+RZW6pcuPIEyDa5NkouMUQ2CX8EiGqie0+Q
cfYpxVJlNGKdFbblhu11o37RhmdQzNisMk6k2U6APJSK/t4siC1qC2Y7GuVS9g+J
Xma64IDTuXJ1IaphKNcVkhSzUgtu2X+HkRY+fjly9CoTTnyCax+WCYiYmAwCrNRX
7A7tjXSOXxPNSy8gKA3mHSUhQGtjOU61yb1uPO4lv9GhIdjzjmjA4NsAfABj3Of/
2HbRZqTAWipmMQTsDjY5umn7QNttEM30aaBNI3h/5cjSo1v1uvTVgsnV8I+w7tfn
9jDBV5+MlAgLRSarxwx6Tq/XhzuengAU8if3Hl9BLkvmg/MQ+zQ18WMFTQX90fPf
Tf4dN8+ZV6YtU/7pv4NfHaPWc6RfW0yDjz7vdmKuzM99d+K8oOeY/9DrCXwdiiT8
Uuk5RN78MOoMWUPUA1q0AYbplo8gVjvzKKdXDrlHHkMwTlb08IXzx6RT1UYq/avS
YrboGf65EQVRRIAvo5pFFaAvMP273+A3AYudZ5LA4xLH9Xwz85wnN8Mvy0GSY6UE
35g2dCovs+GUwNf2rEFVI04MFuLP8//7UEPNEdGmzDIRcWVhKVpcFG+UHdJgmzy9
c5zeIxmv0oAnrFdy1mH5PgaC4hvaLYmpwEG0rWZmOkN+X5Oe5mQEW1DJBrd7i3WW
4LwaOPYxGaQvbXngOY/ADlbgG9Pjx6Ocg4rF7wb0Ha2RynT1JhRhAES6io4xrfRc
SkCvIHIhJTKbPUHcv5DYB/72MgX5sFmaYVac6gqLeim/WyYDAoCPOYM76rfTqocp
utwJB7F21i9ajE4qO+jHq+hNrXIvGi1aRVbtTyypVA4AckalS9vbnJnpw2cTPeGT
aw+mVnoRFRWc/AuCDflZfPKu2+avWzKq5OvUDZ8wCYdoSO/oIS9W1NQgoU2R1D6R
CPQj+c5Iz5+cq2rhvaZzjdG2Hmqqk+e4PyMpy1gWyPk/El54Yq83EuQ9iGzUoYtE
XNeD/sTcxsFvti8taBoGJm9A3ijUZTwYKK9+S9hAc9C1PsvqaWvTHajXUyPRbOhg
0SJ6mwg8o3ww8m3Prpblixizeu2PfzmtG2wC4ugsvlZj5U+k/F8na6GPpCy8jOph
84GbH8OgocWSEWB0NA9wJONGEcAfF8/QISMiNuJDiZkiHB7aIwlcXWLecLAmP5+a
JvJcgnIKqK1upxiG6dwMPyvqHsxqEQcY4RXRXNlu+CvZWL0thpq9nzTP+sNv68Xw
lPUFi1WSZO1eUeCY+LOY0W0FLNyzN2h4i3t5KXvrH3nPJMtsfjiJwHn5Xe4gEOM4
588xAkLJY9ATXLQLZAeTUWaplr8HZzuahqWJ8YtWW9cxtkVqFEEm+lLFYfiNKeVd
IN7jB1Vh7KNycN/MtXMxtsbFNL+KktAO9TyslhraECfdGLhiEudcUo7fMD3XEwXt
VAzMBoWv8A/yfHLq5VGI5mRJu4fu+DwH+QDg+YN9A41uTAwmkzMLk04ye5lKs+iD
uDRV7XtopSzYkxm0VCIoFe86dD8nIzvNF9M5sGaFPjCTZvN6uPQyd61OIhHpDxz9
WHiLS61qd9UD0+utkCtFwhIUjNxSGRQAMxL34kiQgkh9ZjtJKd309rh9Apcc2PZY
D6plPI1P8Ppeh5PiIYro2Y4ShjVED9LbyVitAQxZgr3ie0YyI5Df7P8hf+e7A05g
i9PJnJDUxVWHMzXyxp7YoZ9F7qnEmI9p47bJxpbd3+8Yx4W+Hl5/ORxJAGQrrLTP
UDqAKxNcRHUJVJ3ONKgB3R0r2eEv81VxSCnLCEe0l7JnBM9h/uK6ONQ/XSG7rImb
zJbkaz3oedC6bsjdIXNqMv/ump2aj7xmigzQmuIefy877YAlqQTQMKuNP49Wfz0p
KjgOMZEukdIF/l3gsFN5jeOVXINAFiDFBw3yQlLViE1eHKFaPLLuKCYdteqRXvEB
LY2A1cMvha9djomoLom2lJmNLImutMJTB1UBaJsxL+IYOt1iVI3OG/5BiVGMzoGo
7yjsNPCwJgf2ZPuWliroGxFFQTbRjiSqWE0gdWtXI080HqoVez2XeYx+IW6X2eGj
zI/uxOJZcRuLGKlI9vIV6gMDp7cjEIzXCyUDX0MxP8bcZx6XwATuwcbrQ6umq1pZ
C9O1hkxAD9dnOb7Wi2Ex9yCvQa7Y3zjG6D+bik3kQzQ4cYSNivyFP9Tdgb8cmqOk
JSgvG+ppYZqnI98MgV9uS0UU33tpVMuoZXOf3P5vS/PLJ0TNpzERPBq1fmU0g9R0
mnm+vM/k79+hWp5YoqDxlTbP3eAus05Iu4zEalO7QB6ivaOI9upFpKyhllyTI145
VKMElGACG+721fwUzr9Kl5pQpOsVjBjdmwgVXterFS0MVHAtp5QO1xdZMivoup7L
xg6932W3qVermvZKEyB4vjyBrXwezP3eNSBvmMKXMM9sTntgh1sdC2XgEw4mgMno
hgD6SBEFniqWtpLtA33ljTgzN/PDeZnNtHRnBLfIvDYF53UzO6sYdxbvt0rDxM4o
nRL00bUvyCZiFb3FhBnbVGPc1hZjY5dDSfrZmt+9x6o4PSEGb/xAux8wSvj4eEGo
XnRsUL698txKYrio3lbwcrqTI6SthayZaaE+q1eSKpLQyOY5L4SYSoI2h+sqbDVW
+711kSPtgSKHeqO7ILXPaTVzA4Myb0StvEEfebqxL52p7C5b/ij7zYDFfEQ3s8NP
Ffs3rzFGe70jH50AJe6NZZQfHTz3ISl8gLGoL5gH1vxv3BRR6zluvRWBPbi5IrlF
PPXz7U0dryqiXo52Af5/8ccDOSDKAs4/A7xaGcrCRR3xxZJduw8ABCvXqSkBfqYG
lzDyCCN667EUsQAV+SLFNl+rN0oCpiaOgNmORfEl2lvtDFl1GlY0fphqwyMECL7W
jLT5HA6S/XdlnQS1+dX5WDAxEgP4SehmPpqAB8wnFXskUr0HTymN9Gba9tH+lPGa
CoKjTNFSgOohMQlGbXwZfoxCbIdxTuocO8M5/9tiSrTI2XQYr40e68mPnPj2Gjb/
eesjtb7kQ4OY2oiNA01N4SiRzb26vNUoV5Zn+wVt38kd+6GvvaHVR4wyHBsnTkfc
67Cdv9NaXtQYW/coCkFj3CQ3GR3KTPy0SQV8xHsX1WxamZyLSv7ttMysrB32O14Y
r2nGMhdTEXLEg5CImhjWT2BnAlQwOjZxnommMPjn4fYU0G4Wj6geET8yr+AENTwB
6ZDPeHXHHhgSbd7pi+L1t2XMcq+SsgRWBIvVEwxQaLFXSb9Zej72cHHEVVCA+qo+
fcloMINPTpkdp6XAwAfSgYjHhuZDuJjy92rSzRtjuDG+ZnK+aD8iF6wYmFlNWQkB
ESjRsP1qhAdB4vfM/7cek3f1qXNh7ygZF4ApW6krgR7EJhSQAMyImbZ111qSmC9V
3nyywkES/8gVjtiadzi1EPnEfZgWWE+u9YaqOvQfD7UIsa1AX7UvT8M+3gWKowGO
z0b1EB81LRsXXWdBZE2cmX/F7bog4ezmII3Ym21/NpuWvqaa4icZdhVk+z4ZRU/b
kG4nWpRtwU8tihThvMsPsOePJO777dB0J4Cu+R9GDC3doTyH/27n3DvWMKY0ZFew
DAqFhzaj/WcN7qo1lqBBvEWHV8npiMU7hJaE2PH/MDrleBWaJUDnqb7UBF5ljoOT
mYR5mQFywncmcigRF1I62eCbNM5skE0y40HmZzjpKcK5Xytm2wswGo9sBaDZ+sWA
o134sm8vw8XoDgvcCYcv7+Ern9quLVhWBkFbui9hitcLZSRh9OgieFOLD1dSBBqW
fF0G7gFEYuiqFb4irvOZGMRvy5jlohx4wwV5bm/YBMYJt4N6re/mzzr1toeZrl/v
947sbbrgDPfLgxTm+XQgsrfjRn8s2cU0BlqtZ8DbMYcjCBpkvfnWmhKV/BdDmEY8
VPjMVvBvtnZG2j6ggi5eQ453ECT5q29JohR0vgnM5uzTJnSjsaI5eMfz5pOsoMhB
ql2xHKg6cgNF2zCpl6zdTftJ1LcVa+wjYPPglFjSKkTdoRy/ZoLaHU9L3wtAabs1
5mxi9bDF+m6aiNf86MgMqtKIHNMvEyI9orU3+J9vkMtF1mbBU+AjNHDUqz5RDd7G
owkseh2WcRI4WzywTZYW3LV/sS10lkN1qh9ZhTa7HgoIG1MIPwmE8F7MR7Ya1iZX
cPLJ6+vVJ3Sm+nH/pvKa6T+6I0AL6jtGAkeHdx90sAGQz5nZ7Wu1/vxRczJ09x6L
7toQ9PemeXPFIIaGy7TjbblDwkqD2vuXSeln92CG8RWaFngkeGYUi17K0BwRxCQE
TiklEb7jCQ0RffjeLgYBC4yb34Js18YtAvxetqiNUyqAKlUu+ATWj40sTvmtukQW
Q26fnKwob150YkXosgS4c6tI5orfGEb/+HgGT9aUCJnx3Q3Qmz8EJJM+fhBDgcAS
Jb4D4aC8LBGRGr4ZELOmEOhDBu7cv1RV8BHuX3JWTGumA/a05vN2tw8TsbqyTVB9
6IlXN6vtyQJk377R3ZfPNQMn+YaaBzg4TXiGhszfzpAZRS8ieDd7FDIEH9JtumMo
slMV1t7rP9PKvY66N6o4PtD450qExbIFayHtSMcIZFZ3Amk7zUof/ATND/wEqxh+
6p7Y7bjFvnZVjYXR+fPu9JlKsaHXN7/IPWTQKCVtW+hzCNGqL8kv6aC/t9kWAqr2
GRLlYJotIRssV8ubzLFYs9AwOGYiw7Ph3qu9d4sVe2H7CwtCXZJsB8R1B5KIXo+t
HZsze4fhp4GTNs9j+HYB6cC1ySvUh0F9qczkCLf4ivVF3LFavZDcAx9PcB2+I4Jx
eSPLxIe7zCZagCizFNgojTbOD9tdCX8v5V16jgpGvujp+52wy+wctlIWgwljhFSG
BxFU4Cl1pjWfNLx1yyW2lyzEEWt20hZPj8q2eOSWOCmq6DQnhhiHntz8WQjLthqc
+JfPBE1JPdSJvxEYvX8t1z6VwYwSRWbi7pgeKeFL9n+ECLDKMsSem0SMQwfY4/FX
ffMSWy82B0Ui9E615JDc6s0hb13UJYUBofDejN4D4A/hnJ6UdF3QhpPlCMPHkvOy
aE3bM6G9jSgVphVMgcduIFSCIW8GZgsIhFc/aYlHuSwvYUxqLh1nSBDlDiHtI5LX
WiJmk3Q5ya7OOTwDP2hM7rXp1xXtF6W4BDaw4CYMjvg60U1Z2k5d5npsJlf2BhGR
sTUWRbCC9gQkFK8taa4VrfSMBq4f+Wy9qKK51KWQQvCvVNqCLp3L8qHyAge39OEg
TKWlKkADbZYoOb+3hGgQy3d34166v3wzpMX/XL36W8wEntu8vKGdWDgD++klMhBC
exy8vKctqo1TMW9HAhrlaQgl1opecpqCzPmxjNlMyMw75ad7cqw/FjkIZ0/LLNvs
RFihemhtuTommAdkRFNbfhGb0etMiPdREG1R/5jLCwFZ/fo1kH9vZsDwstrQbXLj
9khE62M7weYXAblSNYfj6e/OBqMcRnM5QjV7eTA43QT4N98sxgT3a6y+XMYQvz5N
1nskrEysWLYytRNBdB3omnORXC1S5GR3mDe2IgvlkdQH+TG7cz2uewmVeQNz2OI6
eyvCYBp7g440k7LAK/3OuDtd0exKUfI88ecfkEhS7FKX6gYfAlJ4JSfUQiQLADS9
aw+mE8SxslnxYcce1v/rQr7d+xPOsWGnjUiMButWOQFhPGpSy+cXDq2hfE6RcyLW
POUZXyAgmngBDbWnrEUifkKgepj8J64yK5btGqYvKOQ+lw8Vj+qItQDe9TOmDjPR
SfNJMJethOIZkY9m1Ts/QZMg30lpC3ELm0iTqSZLKxJSTzrZORFws7lU4dPHJd2l
PRS0LQHPpk9TYFEB52Plo9+RKxJH5+aqoDwmfteGAG5NF8hzX/SzmOMsmhCI9tZE
`protect end_protected