`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9504 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
iga4gzPKo9olJM7FS8BWzijZW8CJRd7NkwpkOIx54CYM/c8z0z0jGRPN0uehpL9f
7/PNxYXoXFndnKHcFctClpAXKKTvWeZuoc6thhbxcVTYgHsYn4YdxaJEn9J/zTGm
aIQqsvDOsqTa+yWdQYIchhXiZLmKAbH9KaVIXbNZPYrzOtZ2GR9k1ljZepMlZVpb
ybELWYW/PSkgSrLIiV9c+SGpQkzlX996RIlG7fZBm46fWsNhkl4TuODtddxfS+NJ
rQzxrCcBTFKSbW0dKBU+f/zjQJehqV8DmJZRyqn91a0K5+K36tTb11ki7M8CRJ7T
M6Ja2TfpJjlQV1J2xoNLfCr5Fqw8WRxxw60FTAx2FSKCMea234mBf5hkxhNHXold
Um0oqyNMoVjWxDe2YbOx2Z8lUgIxPj6n/SaUf4uD+Xag3p6TeB9WHaHihQbrTSTb
MA9JcUuiK7kpXc7Z7wOiR03LrjvX3cZIS5uFChPhVooXd2pcnbFLnGfRbai+Hx9z
pArlORv0Qej5d5Y2vX3HIHc9I65LyvcDGA9YW+78ZD2+evKEE9SBgY02TQfN1BuD
L0xviIYVu8nh2RryS6OuQkHgmmtFXCcZWE2xho8EZmVQmmgXwo4gGAxZFzLY0sNT
PLEfgI1jkWyz647r4Wvw/EL9qvRjU+oE6SUOcIqqPoYKCv3wvmXTQ4imRpBWDb9W
UiRGuDyI8RALguL06+6Y/D2cRcfDf7DqV0qY4WasgRCWWP7Pz2DFgJ6xRM/f0JYV
Uds+1fqw72f8gx6uqPAXmLe38don8wTn8nH6nS7GakM7hKEvU4ZVL8r8nWNAbxbG
yYLFfU5TAD7TI5k7tZrSMhOQXa4Qpx8h/V9p38+KSrefQUJO4Bvf/wOjxoNEebZa
arRthu70Na751uu+InYb5iPTUfcT5Giszvz7c8ZdwMBACxOtKW4b/Xpft3Eeccx8
MJZlpVv1zcaTg0ER0VK4EE/7lIveMVio5M/nSDH+3shtE2FLLjLa8mwZl437TZxr
QRqe+MYNLDncPdpdg3z6ZtdjO2HN5alhCilh6jZTQ1BtdR0tS3i2O21bKTGPOUaW
U01+QBkS/nQnKf5vbHnttpUrIWmY2x1mYqSgKOjlYNsDc5tKwao/FZav4SYQq9/A
xEVYyIIP4E6eUTkIO3Nekkh4lZwc7enW6CAMyjMpJ5YcJJ/PsDNbOo7vGodGAMrD
hkKjglRgzplONOd9z2ATy3il7e4lRA/30lri1WPef6Prp5leH93mgTVE2thrwrPg
UU+JkDU4yhi2+epRbfk033PIyNfE1kkxsxaKOJjc2VyGhD6Sma5syzEh0htvpxBf
rzFuy6z8ac+vZtBxrKEaW+Ep4GNe54B75OUw721jmeOUVuBEbuUVH15XlpWmsA25
LEtbsxHAPEiTlxqwIti0PNpK+6QNqngVerV3YT4slYx0EUgc11qI+HkhvnsZKXI7
5m94tGnj+AFMFYsc+kERsVEUvz0TDEgJrvNGErRqIRl21JP2N8PqYUv4oA4PRiYR
TUs4vrYKduVq6x84YtffacaumUEzJ/8mx6StAYqPPpruaGtwmzA27rA+TSeZbZ/P
8bVf02xd1mIETladKGuipPspCNVVwTSqsA69kVDee8NvZ4AKyi0nJIHy6msOT6xs
YUIJ3a5i5aw32J06ZrY8PdjLXiq/SVm++N4HkfN+EJUfyUr8Hq+pRl9XGDBmzXKX
IZkSBwsckIiD0nOKYQBYjD+ZkdeRv00kJ4Y5u6H27WHGqsD/EInmDspbmtvo2clT
QLNwlFwHDCunnaUOoVpdfzd+IhAu1MIYgaPq9bB8lU3HIobP4VzG3VhiOM6VhEzz
ryOvhKyBONFfPIaBa/JeW7wHiYAjqmcFaoG0xMNelzibxATxUqrGL8Xx3wGHjt2V
q1/VVUglADDlcKg+dpWWqSOLb2seGWqy529dICl0Yi+dUPgZULKT9fNKGCbvPbz2
gkJRX1QDUkUvp7O22QPH8DQphDdD0e93t9P+dUfgHrKCWKY8LFFsS8jh2v2b7lH8
PbHhb4B66a/9Q1fhmbspHQUN/JPKrAWIlc62EjtrIlDIK7hVGSZHWNlJuuPAvD81
DILNHl5VpN1fG4AruzyTc+cgQGXu1MQKg/WB8HyA3HuGTXpvGlQx7gQcCtUKJPPM
34OYBcKz9ZBI4MKf+FzqfK/Bp5R40zlFgV1AmeIhwRbUexPRBeP5Rox+99BRlbIu
88tMZKF3sqajxAJccohkQArgzRNd9X8ekNHAcOOf4yGEL4JbYvZN6g7f2TPLfvMi
qcpBW+bViFgSIyi/5BY6/cPKSFUQF9nPCzFkmFc96dGDhVoXsiAWFYOZ53uhM1t4
A1oJTYEeWlYxXpBPfg8JjlezCRJn9u/6LXao6xNCvgXQFnxdXILT502LrhYtkrMe
YcQXxZkllnilS5p8YW4VHanSQaLgT4DAXwD+hpEHs5cpPSRh8qADtxQc03ti5XTC
pxKaMmdQbSRCT5x9KU9UEyhlkQaUwNimkKe3Mp0dGN2HrvI+o8fHe2UPZ/fubltj
Y41vFlV2MeEYsccMAW3yAbgLv5lHbR9dwmRTBhU+8pI2Qpl9yedsXEqmkOxBAdRK
lOI2cPe8MsHOuSJTRQD4FdCCiOr8pjpQQjRC4C/fWoDwPHcl1PPV/8WXSu15WO3A
Qup1KBn+q0ACAPGZzC2icT10g8Om6CQPc/eskAkTZG9zUM1LNIqWT6dkXi9F24DR
jruo2iXee37y8zuoKvbW0Tm7b/eyIZafh7ixrVdz/x11zAZCAVjhkaCOrQQBbu3o
IipiYahKSqXR5baO7Qk1seLREL0Koybssx6x04oqib+bN1wMSi+sFuWJax1GoDaq
929Er1ULX2gUqAx2BTSSyIYxL4e+fkG6P4ZA4rOCIcx4gCR0ZOfJoBzTrkzGXyfv
C72IhAjUCOw5Qs8xl0OTf+gkFl0q9CAsMk5N6IRmLGN8sJZi9fqsYnsNfQb/uw0M
s5Guie1B00IcX3vsBqJCXodqvzXjMY+sy2X7xIxMdxfoT/0TpIcEXWnz6idsJxMX
gB48o5sds/jY3DT84xbLxaRHzonJirtNhvLnNNgy5GeNe5nf0TI7e9VMZ5MwqpIv
kKj6JlPKW7/TDi8fLvwxJhG3HJj3w1VRv76p4irLqUPBuMCE7BOwP4r5Qxq+CFfY
xfI2DPQnIRvNzk9S/xAQXobL8bVR1ZuKvQwMRcxjkg5qUBGHN8U6/8qH9TcZunb/
AVcLzJUK7gyzobVnHalVl4Uxe+nxrxqisqUFqIcrIAxbeci1QxOwQubmj6PmJViN
5XU2ixofYzq33SSjGhhCdSJaoq3f1HeUmpAYLYdu9fPcWRJ76vqVSdt+9mZ5hT1S
GPkHHvB18MGElu7CU2a9xNjfMH/mZVhxHnj0mleJ/hxLsR8QeTvRHKM9T200ek2x
d5okYZ6FlQeS3Z4COwB/UW1q1JIPpmQJGnfNEzSqdpon0ZNoBEoSu5ymbCCEuRwa
Asaf6oPrkSLy3I+1oXjvJcbzU4ynJm8xySJyaipsvIGEiLz4aB3gpp4zMtwTvd1j
IZYPVhKH2G0JWMnaZZOepzn4IDV6i+tlITEc6F9qaR1/gHy3zIegi95HSoG/ZNPY
2FSWcniYWLxeCTAmjWMFAsQ9UZVIyEPItEGQ0asZMuysh4xrd6weS09mfk9MHAK5
LTCQM3Dj3vJgtNpV/H8Igha+gdfeWB2XNYOBvhC9E29z1M+Qu3GwxiSEy3/BQU6m
e85j/uIooJzxZlm/IFbfRD9rGEY3fgXOlC3l3qVxj6cglCG4jh2r0n00JT3HAhKl
Gtae9AV3gyQmyZf+gveQ68wAzNCWjveYxbAc08WPRztruviagAIAgIOfzAefQisg
tsFCygaSJ3+77ajX0iLvp5LT0hOiaN2wPYsQGz5Zk9ANr1gyxT1JhE2vHuxInkGw
nIXOLqxo3XmMwFDpXlgpgXJu1+ou4Tsz7D0H2J1TZfuboAhAw86n1ZLrhGdLN8IQ
3svnoQUphfFIK+nFqyXOYe/WKSIIQez1v1LDoFjl8WWDOt/54sNQfat+eglZ/P2C
4EaLeqQLXGJahQwGGXbgW7uiBP4u+VTfZAtlY6OJ6U4DelfHyR/wD12XTdIX5XkW
jNsFRJs+HJ0LOXY1cMt5S7TtCf47Mcz2BqE4qWsV6dTh2fHz0DqAMa8fV+qo1Krx
BrGFfjO9NN4PEAW+BqD+8mtNPNKt/fiLmmX4CEV5cPyGwhtQAV3pe7ACSz+OMycX
kirHejWBNMLW+i/wgwfYaxex3Um5fCkKBXWr451jWQ3LPWGNNAtpv4SkwGyF2scg
WU0aVVUeGWB2fe/+ogUatcJmGsBFLrEPevepJwa/ZU2sZmEPPwctRYqQ/cOIgqI2
+P0b2nJ7RxjPbRCWVl4xiMnG44E9gf7PpU12RVES/TftMe9ebAaecrAjOhutfksk
iyd98DFiLEEPOocnMSdPZjLIgzBcb54z6K8F22txdE7FiLpi/ABhPtWEFKo2m7VT
NHb+SOc3BW+XhDi8+Gc8SEyEgfM5AsuXCrT2IB96SAS7Ho+wqOTs0zE52avjt8nn
H47bpdyifJxraWGUTtNC+VwLvTxt7j+XWfG9k1LBKZia5erjDcLKyDFv4z44x3l4
SxJa6PisVn1z6A5t8BlkuJC2it1Od/qQtopJ2yfPGyXpJSOfL2QVJfHgtvzqNo7F
1iOMC3k7ulT1nPhMAQl6MvpfiQK3IUMnVxeMAcVGpbaKghli/MXmmp2aOSQuOq+y
YRfwfV/oGqJW5P5Hcdp2UEzAg2lhTrbp720W/Tfyk42p1TDqgpIuK7dU7JdfNnZX
wRYI0xovv00JMgDI6shoB8o56XfTsKjPAhTbouKzxoDwEG/ghD8BpUyl0oOOizUD
aSx9VKumMctH1xX8WHtlYF56kO0qR+NDLuS8T4zTSoLrxaAo0Qd+ROb2LFT2/ca3
poVb3TqEQiehvfob/TzKhF2VDaqCZaprCRCvcO4xJ//aWtNJusgCI6RBZcBIEy6n
6nWtD29QmMIwyaavwIMLFA7GKGkoj3pcsIZJhgsNHSPFeaVJxyfdWRUqh8X18ztl
bGEcNO+C9WBBbVXIB75tX3E4uwlIkhqNmAfTcnUGF5fDaxYbFC3m/WSKyFLggLER
HaIdzkrV11HkgTXTnRTnO6Y6TB92HMDKHpLtY0BwPzGQzCgLLvP5ACw6He2DdWmP
dwzizos2yiZqXWeYjQ9dEQplGMvudgcgdKEle3/EgL1Q0/NtUDSCrmCFBH7rKt+R
4pPBrdc3IU0pbN24SRkZ+nOQMBVozfurd8FHJbyiKjKcnk2IUbQp5M50EhKeoAJC
v5z8NiOBDvaYWGKRNAuXEdhCMzm0IW8sY7flRaGuAwm+YD6/OuqSsKTuXh9rQdZ0
Lodh0qKT+EDWJuVFgI/Q/kDKE2qkRkp6hYmPItp8ZXSrsNEBppHvGrY3n6G70VTL
et1Vz7bYtRq6crqAEO2hVBFu1iBjX0N8bbmU4H/X9fzElTXD8uPr+84mf904o7W1
6/cSVuG2JnX5j/93rN6y3RCp3N1dVMLQ66D0v0EZgzoJrDzS9X69Hizr3DMiCFZK
E+myodLpjz/J8tTKw8YQGpNHY9VHDC3yDKZ6OrUk0EcKqDlO9AAIcFOac9nDNAAO
2o6kASsRUpaVP0RKes9tlufMwOD0+CNw6+PYocUaIi0Jq/cly97xfAQohiVIUAa0
hw2CO+kVekNLbBOre8B/F2g4hskfOxqLPUalmMUa4RYRlW9RUo1ijBEOFofgMnBg
Ges2usPxzjFTCjO6GPHCF5S8Ep81orPhHygxpCXRKTXK0qmE1EKfcfMW8U6lYkwI
BlVo8AU73WTOyf7x3hyN665PZl4P/39h8J3PDWeLU44UryFA+4WISoEhrzyr1fDh
MoB77FlaGnkMSbgpN7YCyggrh9t7ZBZA3o1BD8Mrx/PaWprGqb0Setsfd/vcUeQY
c/b5FYLbGcMCz43pyQVa/c6s0tICfkV3Nm4PMbS3Gzw0RHJAsfrY0Q8Kw4Y5h45T
DAFZtBjzFKU2Te6+BB0F74glL+nNsyz2vKxhM4Q34HJCEhtM0PEtd2apm4hibFXy
RvsLAf7/8ZtZ8gjOvoDDY/qrhGyj2HILUcU7DuGYaBESYaYdCEgrBaYr+8zR96L3
3sBkQXckLByX1JFUanIVoGMI6sk0E4ZUD2CoSX1FI5D2DeZ3ja0kFZzRjGLRgZKd
ciM2QmWnzAtjhZE0xgF7e1tgvxPlgtCk6Us6qwAUT/90bu9ORXGHsMH3F41NdHmW
U+e3pKKb1w+jpzJps/gpejflt2Avjd0NHMUlRX+D0GhkOAoTh9RHwlLX514+nLnP
nr03+JOmzSShqnd7DxGwZC+Wqo9zvIvOASXaFlI/ylQZrt7A6/3HT8lgxaxD8uWb
xqgYoy1MLKpvRWEVhG9IdZrE6qwhqPdIDGU5ierTx0F0YPXL4AIZ4i8QkaWcsM7/
/s1iA92HWcs2BfaX9TAvaumKqlvd3y8QEpEyON5+fxSp+0+NKcBuGhUcmfMQNBLE
FwgebW/ClawMGoEQtGlqLwth6kg2UYIZlgHUtc6UltPU4k4A5NTjmqDA7v339kHN
NTTYimreUeP9QQbE6Gb+gIR3xC0iDIetM3pf5AQTQ5halzYW8ZfOXsRJ0hq89hVP
YWv8PSbFdVouq5dm6vaFpdw+O+t+ltvqVzR7SDo7xhgKYBqW8mFuVDL4FZPHfxQr
N8C0qlOgLkrwwxh7Y3fWPpK5C/cOepbHq4DzTrNWIf0gM3ZzUAJCjEKkXrvE9KkL
+3xcq3yz8Rx+FrdY/E/imUYyqC78eL+np+OCEYp9f+7QCmtRuGCIGTEfveVOzhj2
yYVoMgzhysx3qO1xSA41absWIcRRssIJo72RX4LQv28MLnCqkaKN8N1EEtd3PySd
Y2fgToiHgCwdJx8F79fPxNcD/G4K+HDw3nWmURqMoXF0NlG6w56bA78rwPAgA9o7
AMbhV3L08c4ZH8756HqV+Zv9eg10z/nNl4C88DoJRoBqSptcpwiby9aXS9SmSPI6
K+0FlFsrvRzg88xC0jvEEgUYPiVKMmEc/PvaWzotDCCBSVDglRh7XSxuDbcneU4E
BTn7nHjFe5dCfz4mZVg7bm5dJ53mCZ9fN5HmmhcdirJhxZbWFSqsT2OcbIFf+izC
BICdXtG7+LRM7zhrd9IaEwccjLrBs8aOrKLOAU+Cak3EAlpNyMm+dasJaqGwetr2
fydeBuvgpdr9EHJ6eczYprqRZKELsibXmtumjytXrrPNuC74G52fFcIS1Qpwi7He
/rDUlAtAWxpUNF0wpJ8dEgItXzBUpcAm/5v3Mx3RD+ATUiKUXLoeVxYUJUYqwyRZ
xMPX6W7bI1xxALbMZPSiEJlBw0BTswBPgNmIdHpfdR+4synlnP0lftHMQBxfuZe4
HzhFfoBTPY46ih12s9bAJVSVYMZnrnfevCNXZRaNfHW2DHpKIbW9FEvBleyzKPlZ
5DWuyz+JC/xPMuOJGaqU7cjWBeV52bwn0Us2XiAKShT0jwYu1IXK+UxBwrHV87qk
SsyGr7ZTyzrdhpCImvzCb6mVQD4pMqsNz2j7kqakqoH+iHB99iHpk2jTfWIRBn4F
Mydt0Z4vfKLovBDbdnBnatlBcmf9YFZa6VeZ4QgTK7y2tGLSSUYT/ETwiNcIQDv3
8sAdajpjeRkjtQAcBWQxlVAd3buINkRpMi2XMjgHQLIInKZht9ion+Ty6F6bZ2eL
dHUKndVbs1rE1F0opgxtAt5YFLTC6P0X4kYLNLfAyfLqeyuhOsVa3z26X6NxwcH0
tZ/b42JhRhVGJxIEky5AnJ6vX/fp4vX/67rlwVy1gPQ//HgHMUkaEWAR5aqDJP9E
OsuVdBPYuWOYIBQPjeEMV3dYtQxJ1tcr9NyG4fkaG3TM6PTXbbscXLrQDqEPCqa0
QRjlMk6v2Nmw+ZxOeNLQPwFeWBZjLBvRn+nk3mCMdmh2GSutcXPJNTs+Qc53/Svy
EVQvrlVaJarBKgpD30lO/3SUTycSFLrvZZbIWhKBFdrMn+Pp79eFMBST34zs2+hw
mT+baRpajgLeOKu4/8QfJ05UrT0BAoFsqRil8oBL321jYPjCfR6zis9E9bY0U1s1
Q3rJ0QRhiF+/KZYpBx9pAjnBJj1XO7MbV8Kx+IoZpsvYxXXE4IjUXi63A0qRipP3
nRkxFtUzB0x5Rm9RRdaF5sb9qxcVqUIBeLQJkCiLwNbJtcIxGFs84KlEFB09IM5z
mA7Ain08tLf6YgkYSFWSDYsmuEMVJisu5CsPWXr6lHqoTRWlX0ZFYQ6fKASmeXdf
lTCDDJCUZiHfv1itfOgdEy80mXX847UulM37EGdEHH66OUNanCh/CxytTLFIsWyc
S+12pukimZejA7YWhdcMt7cNURrVZcHI5NbLOpKpzugJxST8WAO53Qf1C5yyjWP3
ON211JH2vVribiPw/j1fH4cbJEyLjfd73cKsOux2IhAt8pPWZuJxlCohk77u2EWc
wnG0vYQ0sI8X0UIKhoqzxeLSFf4u5+BIYwN4KfhOTqQA//VGW24nFUSG+11D+eMl
nBHq+ndI2UPxMnYNZpmSPAezgLCOfIEK+8JI9N3lr76BIS+yND8XCe2FqRdX96OT
CYY3+YjNUuhS4xmwLmX3/61i3zTDF0026wd9HogRMSr96ExUhiVUTw9PrasVeXVk
ducnmTpDW9NZyEqujv3CuX3OHOJocn8RtbqgFQsQiTipVs31fuFJO15FhkgC93oa
e1IueLTYbh0PRmmc0hDoZLx91/tEoOVGQPIkqv/97X9CiGO95zG8Xb/1g7gvqvQx
6yAfOa3SOyn788zzTrzE6cy/Mq1j2sofuc04l2O09BMOQhGzswDjdU6zQS5HjVvc
TEmY2eOySndLVimxNioE7hU0LnVvvnQQ51i/V8vVCl8jfeeE+qXLnKTEtO1uZXS/
XI13hq600Z9IYxPMpMMy31rhy4RVM0lEOVtUFR3ghjta8aJuPfpffBe5IDlUeX2j
/Tegcq5xyUPJJF3v+3FKwFXcwleiL87NOWyoJ3DN6W7fH8FvGhQvsraHYcZMo9Ya
ss9qdWG/g/iWHO94g1fmLhR7jyfEdygBjpSMQ4Qslh5swy46h04Uo9B8XwEIJzJg
njcA5R8c5hFGlJ1/DMxRL2FKjMKEpkN26miXS9EmJesXcIoumuHYRh8nKseCVSsT
7k4lCxCk4s0UtcBJCbDBvG98UP51vGr+lT+fMWRJjBEht2UxKdxLSVbwQ5kUGlXM
SUe5nDO0M1oTmKNiLVskZ2wbJ1NwKiKU8r3U3iGUWuLpZSSP2QOHb3YV/WBqgyXw
o+pUWGDjPBfQO2NayIFvglrmxKdH280E80+FF6MrhtVxYiQioNf05qBY82IL83zo
NUILP8ugwS3hgZupJgDPZ5ZWQm90kzbOo4GoebZLxnUIdsgEJvjCZhZ1gkthxab8
jZJTB4MOx1lnK8maap62L3y/mCBmAcq3tw75qjkwAiGT556ezF1hDiPfvn82PvHR
vcUbSQ6aJNY3bDt48Wl+IgAzD3Uz8xU9egZicbeXP+AdM6DrLL1vv/t8vJ8deBPj
gbNxnRCV8N5C4Vuu26yC/VWUIggGhpeSDke8Tfa2YcVKNCqKeyEZr1Y+PiKapelJ
qpG2EtEg5cwdT1slO/dkagxr/QR7Gk4YInvAHsZO6I6xaLFMi1WLbduzUgEYLcMB
Q62o0ZrTDCLMuQnPxX8UhId2MQi9G9jhd8ZzHP1dDQhQ1819MrPGC6+jDhk8k1Du
fF6RpeMTxk2NgDdqpS/gMbgGXjjhxeuX/Pt4a3ugsRa0xIEgg1XrjSbSoBRepqmY
kZmkzJnGLFA3I4y5bUZ88mTFLs6vldFTVihXkzb4t+E3LL9PCz1M9ALyRQ4hxWDZ
wDTKWttsjVqVqz3WO/GrIAorqJ3GLYLdfnKFVZxxPh4Kwy3FTSMqyJA/izrQdz45
pVJ4ZJfxp9lj/Vvxo/tJbb4RyeW9mncdPALop6OFexBSIzUM3k55pATsY7Fo2cLO
fAhiod/8hqlJi1nEGX+X+FmFBg9IWKvxBayp37B49TROdRpZG6g5uxKpvxc7qwiH
Q1v8WBALcsFg9lcEkwF0ysNRwHbtsWJkFm2QfMNQK+BOAufOrCw4jgfDF8q5lJ5B
6LgOILOUkW0/KDHDXcKRoq9W/GX7AIU9MP9LjpLyuSTFD+GIqbOi/nyvyIxKLOwM
p1Jf2Qlik5+uVAvYzMPp7ezvl1EtD5CwRLOP5oJSVWCwcZSLXY6nADyGtrG8R6h6
/t9YDMHQfMDUb/eURwHp0eL/yOQ8DgXr+m+U4Dy0xctPuOwgzb9zyrMxlMcZl1QY
sQkoeRGmNhnBqxGfDFsR2CU9/mCAnzO5/sGPmwP2iEuejSsYme3epHcVkV7MVEZ6
OkU2+N25QtldfWrL/m3Au3XlichySsLIV+3dbaYyqWXnKWHWNCkLdSlWI+3j2Haj
sh0ahwL8dzf3z+zia/nUq0PnQw2PBm09GmvAbQiydXGlSGePY9RkvZ+PfZZjPJj2
m8rbuoXruOb7l9IKd2qb0HR3l3dzMtWvxqVIUWJ7ubDLfRjLGXRJiyzH30Kq3lnb
6H6W+Sh5zN+4ztO5yPWAthaeLIBVL09oapXPM63WPbtbGcisQPtp+w+oZGpzNpSO
p8PLdm4EQh3Et22703Po/RFAFdkiooZEt++nAQXm03Qbk5s+qOGrJtsJgKp7aR5a
JinDFcocoqav21Nj/D20ruiYuHjp6K7qUxTtw8WOHuB5L/s8Rcsv9b9bsOBrmx61
nn+fzAxermyym7AU25HnvoZEluPHmLsAP52DkPdhZODcM54Png8N3JFp9iX3iP+/
LOiT8Sm5PjhaKeTE1rlN8nEot2sSC5XZ11vuQjnzewwYkBqyugJ7JjnQQSg2+o23
gHR2kHswx4KCnFZmjU0T0YmRcdyinhzeSTbG+P8mPYr8hdUbokG54cFd6i2NM9Dj
7JU5JKkWtSXzwHkjofP3Fe/8hdTdZ58I+UBxDw83OFccIQnPj4Y1BZsntlfmcf1z
D5Tt70Ohth9eR9QnXHcyNGnbUlApcPs+0MuLJ2r69eilLCs0Pr8Xg5UqiPhO/9cx
jzq2LDh4WOtp7eqr3QXBDSwty9KQnTtju5t64eYdqp+QCy0nHaQn72XDo1IiirTI
2O63Mv8kDpl4bE5VeJiqnyXqyjJtxZq1nm0W3MCSRbJnG05ucdqZJ82P1yvY0I5Q
6Ym/FvJiY20eBRC8aYNLvOzb9Liz5jlrH9GtN8BF6CqwHsqfUcy5deWudloPx9cU
FLsC7RoZjZ4iqqMPa+nSErywA0h9p1z8k7IZU/FLnZo3EbMpeIU75t7u6PVlJ6EW
OibNcxa5yDxROKpb8HwZvXvw+49W+zLMxyTG1JO2O/HKV4TCEDWYyno5an6AO+7k
oxPAlGhoCjgvzRAqQsUZ9jrTQvLePpHS6wf0zgOc7C8MQhsG1fg20Yqkc+xJ3RMa
uuvMSnCZ8i+zBrtyZYQDqVSEAFIJmko13BQ5Y+gFao2FhrTha3R0fXMfxCPQBmEV
oC9IrKeGxhAd2S2F7cvDaXCSxAstbOmhRLFaw86wDXyCSF0W7SbRRUz+jQ3bH/5G
xLnX0E/TV3wOCWz7s3zRvgIKoOu76JFZTDceP8wtHv60m8inniZa2EZirI/fVZx1
bvr2hhZ27aWbBqDlLZaUVbZRMCtLlJ+r0qyVimTpg2MkMuWnn1QTiaTSEu8NRq4T
Uy8DKDEMPtF5vtVdvGKKPE1qYvj1o7ORTdcBzatVXx/kFL0ioq3sY05PTWjHcOQg
CT+74YgTTfVyvHBk62A8kCNWHdNWXyRiPqm/LEtRmhesd5eeOc5IB5SUwKfzVVvw
wAYWv7aKlsrfu1ywRUYs+t9UWBOPmRtZ6sIfocNMOhJmro7lMQLLpt7aE1XTq9Rw
/70kbUOExygd2rRogbxiMKqt7vDt5uOYb6FyiBaTcRGKb2seHONubg+mdUsE7tBy
hL5YW2lmTqTdPQ8k7gwrAPw/5GGu7Q2sLUmZtUVSsx9M3mzKWW2WtKZ8N8bi/RCG
oKlgRJum0PlG+dVJO/xYcXEGdTYGB38hYi0p6bIAVapouSw+1IKeZlGH4jNzeev/
JuOTR+hxWKnTh3MlgYq4h8KxG+aYq4lxUEXzDz01AtP/gbrq6SY6PcRimPTLRaaZ
jhPn6rRDKxJf+AIji2LLcJ3h0Hwsm1Yi8aGpktQcCiaxUktpGtAcYLFAixbJCvZa
dS08F+iIPkqi7iI+NoSYYIAmpqIK/DJBn+Fxj6fPSAe0Ougj3aiSEssjTHd8/bTG
DPWGwuOpCzx0eNyRsl2NeQMFK315RyYnpfz8rBenlsaQdFlW6B0eJUGsJF1V5NVx
l9yhczT4ScjLvLVHoBMsLaE0XWeM6MohyWmN5ZRBPuy6YwsVW3gOTFqzOKBxmaNc
`protect end_protected