`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3824 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
DBGZtUPdvgnvgIFp6VMrQUj/VluHKKwbBPBIECETxmQhzWGHySgzMsa1bZUckjga
mw15ITdl2ZVYz8DPUkhZPf+FSto9rixiuQHAEexQbDXWpaO/PRyp6uBW5OOPQ8ks
aC/+ZtzuSFnAP0q0UZ/x0JRLVnJukTF1yadeQzun6oYkxLnhZRUzfV/105Gin6U2
qavtTI3iiuaIpvpH8zasmC6l4UHkuBWFk6Qo+JCyi5DUf4Vf8tVoTa3HZfSYonWD
ZZ04P1V2Ui2grZlSkYV/FBSchZ+ZTTKsFee4ptgRf6gC03tJeAr1SBsnjfunHv/H
AdZ5oCKNNsLLTqFL0yzz9QoACgAi6qF1jJl62yTEVinqNoKeHsC194cRIj/Bd+Zj
BsncB403yanKI5T7+R1PpB6sxc3ScjO1haDk2etS+c+nLOL9gyllMcAf53X1Q/ZC
woujadgXll9VjRb4xWqIhZsqF13V6BcGmL2nfb0sdVifeLPzLFptxmGHzzBryi92
ha4tfnJ+U3OhvhqaDc/2pJnkD/ZWbQP7e+ovqZ4k6NNJIbn7h9KDXJNZiNw7ShYI
TitKKVpj/7fLhYnH2EfgbErsmF72CcDikuLw9QMAMUb2jw0/wuJVHJpPmSQqzb3M
DUB5sETSuu+VXob1Jo/IWnXLCv9Vb/N4osb/RhagIKbW7s/uHnWUNb/N8jGcFY06
qhKuXhdGiCqJzVCUuz1tdVIJdz7vpuLXHxxLSQ5BIos/K/ij6Yc4iVJzyC2lF76C
pO3yL4FczRiglSb+nh3kVnnNwmIO1SfIu3du+dOfP8kcz6+0kB1phOVbH/dxwSOv
cwFpCvJgktwyKBj33O2f+ErX+EduuufFM+73QyntQm933Cche1Apx0ykGR1zqBSD
vMBceaOgvolJRJRng2d7NrlcI66CDQLrxORDT9us9Amy94/utVaUDQmgOT9gqwXR
uUU+914EscVLJrZ+EjtdTW8khgyEPo7NP2mLi+7IBCPbeVwaiUTA4CGCf+2iUtTs
PGpwXmLxDyGNzRVpa7iG3lRhSubjz3gOBXeVN8w+GRgW1R+xKDBJ/wUvLKMFHDfz
xv3JeW2AcxgO8syp3CtyIG1N875UjgUPHzUyZChfAm4pbLJ0daFWKUSTJ0xrfYRX
OP8RMDvf8KplqhZW7ix/jzb0qc09H+SzuxbeOEaQtJF3WQdrH+BGaiEMZqEyEPoW
L83ZdSwm0tW+1PntpPp42rgQlZfCEuJtRBF6rERs/UfsOA3QA3/5GpzK/Gmp3ida
ssMN5wbZRNqT9iFjCfGv2R4wRMbQsTTWrB0NKJunuZmB1AgeXvvfJ66byMdLmgMQ
tWjk4RXbRlXbZCYAW7CS+MqC8CmdnNx0cAYiZbGT2Z3eGKd68P/R8c1PsVWySvDE
kdQZjQUrKnJ7EDQoRtsq2m+TYD3qx+LcchQf2rrcOuSS2d4kjjc87oiQpHaSsne9
WSPLyLpoQ4WG/Oo0XUIZaTNimarxF8+6Rplns6/41dWnxE4N/0LvjW4pkEla2aH5
DvL0VmzK6HA9WxVdRi8CPg89K9l4yEkgRrn5AlwA6/FVVFuJD2pJ/ReQVpIJyA5D
4KUmjDXqJ/vssh0HtdlUNDInhbhLV/jWEC1a4HOncX3AjCJBQPts0PSPwi7QDQUv
3B/XpliOYQcSNSXpGNKxN7bOd0Jx/i5kcxy5qBgbw9Y0W12HWV88JDaeMvGpVowM
MvkcTBweMtOIvKSNl/2qmItMuc5+36OBnfV33PZzTi18LL1l7iqv/4HII1hRa/f2
U7RZ0whplkJmA/krZ+7XBuyZaMqbtqg955cvcqU4k04hxo9E0cdXu4uUCfdl2iDO
arv4QA1PwT8kRP68mMxnjOtwqRPoAydT268qA7rbPbZWj1SNgJeo8ToWphI+wYcY
Xkabbu74t1nODXNmCAEG/Zn3TzYGDp6Xs3RSi7C187eU9jxAGxeuvPpCKMPIEuVk
Kj9V8bGGBT+6z6JSeHHJhFMrJOod6LihLJTDV38lqRdA1jVXITiiiAYFDvAOGYVr
3xoKIUqBtWNWdFaJv79wLNbuAkeAYqJIXHwSRBP+eP3Phggoq77SyhtgiHPPQhdm
kC59WPAJWQVKs37FuZaKTauf9ugaoiuovCmE/Eggcm88cENnnrSP9/hISa6ozwyH
uuDanGLYb+6bC6nqXWZTz2/9kTT9FRhWb5P0pQ05MogNwnEB4fVIcaLz1MYgVdWV
N6f9t1msc1eo+LiA8Exf/IAQzOem1ycSpM4H79Ed7o/FZLjVGMKJiJ3lWYxO3ImY
FS7p0eOJkjgOM90Bg8iLp5dCaFnsx9tyrlPn7poVm6ydYctTSa6uGX0b76k2GlsJ
nwigVltvgZ0SAzw4LatmexV7x0SCud5zaFpDMz/7H7AdkHaA1mr23rp2M3/MhsGB
NF/P45/GVpMjhNMeCwpqXmGmRMFOzn/sSyNyfRF6Hv+mqMn4RelsRCu7SgKYpL2Q
V/Jah/5ehTQ8WW0KQuOg7+MCR2y/DkXqt3Yv9xC4lCQ9Cfqq74T2JB7psHCGh6Tm
Fab5lXKfDz8bc2T1NIgkT+4dSTsR+Rv1np4h2JQlpWQijzKsgCpdBMcbtQDB2Zrz
G2LP9S87k8r47xwxkV2HlatY22HW7s7TTXzTzLQrL6ZD/SjZD4QgjcZGWMY8vdAT
Cxuh8Ane23qejjYm+aRN1OOkdxVBbseiGVy2MeBE+B8fI9tXSpUMGKcDfEoJnBBd
LjkVqdcPVZGL178Wno3MBkAlJRgFJi21RsL/ieOFINXXZytc7KPx36rxOeGmhl+4
JI6OHz8UGxxyWYRxZu6UdSMvElYyXw17kCTacEc3SM4QoYFZHp4LAVJ/GCfuPhWO
4MYVePmKbhfJNyNeHGU8mPflOjPCSIER7SL9bv/TvGwZuTe6WY/6dOj4UJAR+CzL
VwfojHhDbiW2hxKX/WX0P8zVQJlh5JqOzNKDAM8+8NjTbL//U/CYW9wwW1iaeufl
L3lmmKEC3mEF8ThhHaz4WYEx+vfBEcwupHcc4hCiioFpYfF7RWCuvHjlNrebUhRk
YSHc/2Lr/Az2NKTNko0B7yfOsM+DoUE/sfQweOChEij3hSwEHofr9ymMbLHsmbxx
m/fQMfB99KAl7rAkG1iHLp626W1/OthdY7jkplSqKQFBgPQTSViZyFCVO6njBTW1
pi3DfcbcNmaBZjaBT/YxOkoXRDl7ouIi5daBu/6IS6J5JEB+2HLJh7jYGzYwji6+
vLZjRr0iHIuBajn4thZ9/BkOfhvTadpoAplLLnyYdDh0iPtuaUUnU3VGL91wIQj0
8nyY+wYDItKixuITaIMFZOwuW9Dqd2cAusoqFLq8TEBYPYX0hixfG71QFQO03YG1
yiPXyMI/BBoDn7v+qLSchIvzNpaCHBXce7Hpwsi6APgZ9YTEE+ftVFQZzIEPKWSg
mkn39Ks2ROY2hqFOLEeaC23YlFFKhTRoWDf/qVEji9QGBJi4MlP8Zp0Rawg5Y2gD
NiNjEdF5LNfZM14dC0LGOCjMoMu3TLeVvIfs0qtiFq1LEKKSgZ6dKzd2EOc76xr4
Fs0AN2y5O6H4gLVbYkUHB5pSLsxfJ9flr3Jdjsbp4xOM6Z52dnBXGhcKHTBpa30X
3m22Ox/qh67qh5VE56wE7nF6P1AR6YTUG1u2KfH0G9+cCfFmbT8ot1WSSr1ILBwu
oGNutvwtPUW8Z7I9yTQq8M8qU9u7w2fqakbJdP1VPevYnSYUXId+Ur6OSf+Xlsm4
4jLkOZca2/8GmpsDUbKSpVs8ZL539YFwq+Vb4VA2NCkudQHt9sjPRiwSPqLEOy/B
kfF+zoFin667wbDOT5vd3PDeqjk7l6VnKCGLn75HoIT233CPuzAQpqrlh7T7SNjC
PXZbV9wKcj5u4bBI9PHlGpxDFVxjFN0di0ffOWP7AS7EZJ4zZzBVaeM/3j66feD+
zPRmaagvFwH+rzfjK+zOwj2HoqmHKWFSRdDL7OXHLm3rPnFjPXaIyzT2gl4iVKvb
zt6IaVt5D0DBlwN7QPCPfW0vo4yqJOvEnTQtBHqFbt0Izcky7bkK3L0NcKavsMzP
GfM+PHVFoILtXJnS4NWRs06HPExppq6wd4+9Gtr/UvoEY9KVu/rANNphBsh0EEqb
+ELDB6RHrZrze8WJBMTfjWgV639K4g+h7rg+wPMWtYmqI6T7itKcrZYQZ31dzqA4
FcjefP+p5L2l7Zg+ATHQYD7joMU01GDubwtlYuMEhtAFplWU+d7dLAYQKySkZH/z
Tgci3bEFDUg1u8ZGLfIMqS7SQpvgibRJ3G3O29/vYBiJF3axqfdVfkAYP9WkPnUx
9V5Iu7+pQ6FRoHqWpbjHNwBKQOhbOO9vVYsIcJ6HHTmN+h9X+/HEbPbAxfdmJGRp
h9ZLiT8xGJzhT11sezlowpMhxmjab3MhTKaohgz16hNLnEbexmUNBp3gfZxMSTew
G+Iy46cxEaGaHgIJqHK9GvFdffiB9U+seKyJ9kuaglI9ZhleUIIEnXMjcFVpqkhr
JPNYvHawHaDsM5fLA90gkuaNbzqql2NoaAJpJJ1BmbVO04/096HM3vmMhTox0JX4
NWyhGxAQX5G0SE7RmyQm77drFpipe7z4OJtGAG90iqlmpE6zKf/eEuvKpYehiR04
JFQDmUxmJMBMqBwHPbAdtHV8LFlSo7kF8Z50frNMNFp71dl6aOXgdg73DPIkdo+n
XFYGgVEu8GwclmS7AeBv6VL7eMPjATuyrmVdmOEUaDGbqu7eF6bdYzQc7QvNbrU7
llmUZ2oKQQLycon2jryrPgp/UqOCQxh98y/+L/S0RHmSHEXrefxWvoB92bpwUvdC
0/IM/Qs10asizkLdCtfc9/vOswlCa0yjFtBG4ghtyPE6E/IaHMpQaGiFBlVX7QDo
Rbm/wB9R7800Z2i84XRGXdEyhk1yQiYNKfQDp88/jus=
`protect end_protected