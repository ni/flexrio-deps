`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1456 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
m7OJaCYG4D2XeQKzWhbYg4N2NWzc7cXmZsZj4eV0rNYclKusbFJfKFtsb+VhPWOw
7qV5efab93M1niDyU7a0szR4ytzpz4/6KxcscN5V9F6tibdxBLf5Sz/WPDTRQgWf
ZPY4mDsDBvE+sXIVjduWqSHLN6aStUYtz0dQmGGXpJmyDy7dkTVfZHnyEe1ao1GH
Z981cvT44o/Y/4KsMCKFYvq6xKvMbYKV65mvK1ZsLNnDNBZ2IUSBqH6o2n+1CMWr
zPwV8Qvwu2IfBKu6KoO9OkEOk9bPITSIqyGSDAsn9BWa53W536YKHIcNqBWFBDwP
+COcV2dXAAvhXUirTo+sTWgtF1IJUU+filTj515P1D2giVs1buZT7t9gYhwzadAN
FjcI1c5kyKdMVBqGj3F2kmA0LyFQX8KajxJaVYZBrbiR7gfecOToxmG7faLW7mcT
VIRAmGKrfeA1SXuVhSBBboWG7H7UcFt6LKIsI5texhwjpVgvV1EGZMnXyeJHkwyl
me8dZqcgzW5yV0cRbqqxWL3U/D10cwsxWjkE+jJJ+CtfGWo4DWq2+2sc5NyfyNLY
WUHz11seAq/woYbA0Sw1WBSpZkENvV912xw86V4jyXCnxQAHyudAa6L7um7Edo8e
6s0nR4iBCctwY0fEYRr6hzFFv+O45qvySRfbAmA8J2uzI6+I8l4Ic++CsBvhlMTN
op6j2eJ7WyUkxuT3TN9Gm94nRawTgHU7XRs/XFvS/0T1/Ei31xpAVIh+/X1CyRvG
5fGEaxm1rTYx7YsU1A6/c3gSLGLeTtW1wkvZDDHsEqQz9neHQcoVTSlKbWwxi7ug
i1wjGTxv91VDDKnSTG1HoMgPCykPZOCbwE362X08u6Plm2QhAeowDI/HMDXcnjzH
JNGR34xclOGVYA+i1CGS49DAnXweuqOQycXdZp/vlVFJnTf5zwea8F5b49UlgrOe
HrL3Vm/7Ht6rHV9hIVxJm3xpfycfm3ihXY9hXA2FvR3Dd+8zxSvTpwgYomk59wxE
jS5gsami7uax7G2PU0+NQNlnQvWyMNyIzo0t1kKMmoVxj+qmt3xTUrHMKk3pfFCX
C0gY7zi0LipG/Y6ZgEhuvLac/ektZ78jqi+NHLo8fC8YKVdD131apFgtESJk4oKG
XFwA/1QP/2a/vLcG0To8OonJa61h1+3xZ2OIfpRvjGL+a86u/6cbqRgmIyE3u6Dy
4YioKlInK/tEyMivkJSLjNDzUwturZ3Zd+fWLROw2Rhzce05hJIWmgovGNoIyc3/
Vi+49fFwCgnhXgbnN5GNY5Zu1djqADUjYm2UjOhiij6ACjPwMRH7SWbXj8VD8wXM
Lqi/hIj3JmH++f4NmHIbpqp6z2xPj4pYk4lR+BPXQ1ZrH400aF4ZQYzIwzy71WbX
+a74I+t91mu7oSnGQ+kRoKLqoF+6SRaQmjmaFMcvUSmajKiNBY/XX4FOLqOErhSY
iyrH36El/U38cu8QSTLbtd13DiYb6qG9sxPLPIV9s4NMKDOHSD/QfuOQ8eMplgGe
CHcL1MEF1JgZ0q/S2l2aK3to31wNSCtc8Njwe3PB733rsp4D4++4L+hl06Y+gIU8
ve8HzISHS6kzt2UR9y3eIuYqe7NTVefuC7EJfC+y2jSNo7O6rk/LTX6N2dFpvXLW
vWaGD4q6fdJz1SOAn91pXf26wEEfu5TeM0INWr6HlNbdgk6oheqeQ6jYMNNC/49b
3LBvw7MvIHeBv/GSKPTdrQz1pJ3tTnDnEukz9DmOWKhFPyGNkFnZekTAeEsDxgYC
skh4NRTY9VSJRj76FO27Vg==
`protect end_protected