`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 13312 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
ky4SiZwRIlZeVC0EoaoEA/sEH81dLBgPPi2ZfBb0EAV+iAYZHF2FkPOo96NsYBbv
itutRsCeUuJlaXsu5QjwBRD0735w1hohICQYlZ5gb+nJKzCuTjh/XIGU0J6TMxf5
OMQ3iJQ3qk+/c631GuVtf2pDqPAX7AN0X2BahRIBwZofJJxPIL1+EbRAZtkE+jvq
Tqvias+Z1VqlV6RuLV/bkF5uWwU8344OH8GJlAKfP10q8qXYHt+crQCGTWfv8kFk
ddSatA5PpEEAITBgyml0qlaKlHGS+3HQyKpBYaEAYu4c4TTz38CAh36bFjfOE0tm
cR0sMw3GkjtmBTWcC+RnS2r8d2YDu4qraowTw+2lbczGoPl13upQ/RxTxLJAqw5S
GRE5BGKI5jCHBUPvAgrkZfCqRE+ah9CGrhXp2Sul9Eb7Y8YXyqNjqdSlitR0+iy8
KWETjJYnBbN2JGZhnleX+MsFfYH6zyRK+rg6DfSVr+nn9V7TrdAKLnPzeYNvKs8d
XvLxh6MtLcwzAWDuP+ZTg/4IwxUPGdbSm/YvVLLNU4YvHhO70lGROAsz0Fehvh4o
Lgi90mvBtPb0m8gHvxlxVE/zecXrR1QkXQ6+LO4pSMz019Hh8nxrcPKSQHtLS0Q4
7V/Oj/Uz3KB4up4rAnTSK8dTLVw/4KtS/dyTFyFTp2HxPjgxzQhGD0P1+7nIAtTg
4taZ0hT0DgqLnbHiYB185iTgmekieT0a43q/bYH8ikGLgLQnbHeeGkrGLaPf7jHh
tKpJG4h1ne91ApkqCJYfdlhh/YYbdgY8XCg7x0z0did6KoDwpvLT7TyY6WhdFJuo
m2UuyKw207fm/aME78gvo+ynMaY6glxpYF0GA6RYe0/WL2z9HE/G856I9tAZfcXY
JhyZ7Tl33w8DdnfOGbCqBfMKOcH6JXip8ZpXa2gJPrf562Ff2pdtiBiJprJQrMb6
vpNpBpCyQqbxUNkdGDg0zWOEyNQPys1zwLpik6jW7O7QHFkCtm/fdULRj6hKnQGS
FsNs8bVcJGvdNzNbf8NLrTKFwzI0mJ0ySE+71SFRZ2fKCM0ANpunuypmQYBfgpra
M87lerh3FIulybWnlHiGbWTppMJLlrxVBj3zZjv+rPHaqCXyTyGj4Yj+yLUXgoeC
RtP+7Td81C287ioklFJwFNVHWDxypZqqw/BuzCmGb6cZCpl3g2dw5OsvTtGsqOxW
xI+Y+OEiP+uPGI+n/ybesoHF9pKZsp7iTdbfkx2Jgq/6Jf1gqA55jgUE026FvQvI
ZWCiz2oAQZEOi356bMwv3J8Nw9XSDWXnkZHCzJRHZiwaifSHTZhkPDwESruSx9FV
BY6JI3A2n/tR2Apgvnftft/jelQ5fu9/e7Zmvp36VKLEeHOjdYZ1kA1MK5ej7YX+
DEZOiA2NalHeBdrq8ndDljZXQbgzanB3BinBEPye1nLS8gou5JKK2N56mp+6oPAO
FQnDPFLipixs7CPSusYFqI2708XRiHj57mmv77EMPE3XZ2RjGhyHnrFGMTWHunUr
uGmg1A/MRK9/i1lpIgftYbzdugM8QaT/ZQgOxKBlT5E01841IjidTQm5+f/EYVK9
knfpv5fnKN84jlR708nwsDoxjtAx7BeqF5CM/KxDIbnxLw8VCup93NSlfk7ZMzMU
tH3kV0NvlhIMoXwWKrOVj0M4RnGF5yRZ1C+HZTqKwcWGIXuOQ944DTZqIM6q8EpF
fb6+aoJort21Eh+ZPWdbjvSRKlLvNbilJ9m6Ow3/CSaXJv2TeleTj5TOrDx3nZ3O
W5WS7txYS6n7qEaki1A1PrceqXTyWc6Zcd3jzqzdhR7S6cV+iY4/EbfnX69IIGko
/1RXV9fcpz8A8YTNyONcFhUbUdrRJ3vzxgWbNMrUpqrqMaO7qXRVdVWNWHh3LdCL
GbRbP09fOYBwC8waw8i+/AZM7NKV2wEZlbKRjNliR/nGBZ76+MH1X3qhiAoILvhj
oLJ3yyEFDf/AzGdbp547yeBbQaMsJtIqmQ+RyNiVlomxT7TOTnng06ETPuBMCZnp
SPgX4mjfUL3kA4tDKdz1mDGKPfWuF8KWsF5uEO6+HHYeVm30KLvMJBdzVwDWDSwG
sm9+K/kHjnhYYee5t7U4Eh0BcTRbg9BLIbSY5RU9aC2B9+7mGjXKq1NzpexJLBcx
zmmLZ/q/vdseuhlXHjQKR+UTloUm15jPrJToGjaWpyIqCKA2itcgReMIGNjh1WU0
pkkfHPNdGp0eRitD5VY7QSboGKaapg65Wd2avQIx6xQRInXaJO+z8YlAzm25gOd6
GbkX1R1+wtV5KitaH+rQGmd9mETrhvDTJxXjYfESfhjFZWAd3U4wzQvo7c/lqok7
mjKMgObruHRVnS1yM31A4G6kZMuLwJF9MWbaGL0FkGxd6FTI5e0vnC4d4q6/K6YO
HGQKfcPxhF6Sf24wD4aBc6/TESgqgLr8SJYcav3bLoZYN7IeYszQ1LfYe2JHONct
loFcI8WxsZ4JiokwvU149Fh2RzZp9BvCDGSI+fjonw1MIM2ppUv50edJYQ2l+GpO
XchWU6a+IwCGJvL6ZQCa63p7N09FX2FdmpExuBM61QbR5gEn4KNaWTuU/19ESh8b
Jg1YNL/Bp7yJjY1cG1Cnijs+STFaM95zIV3sFQ35+a3Wv/txcU1FLROG6C63fsXC
ut1aICkn9Q22ZgBL5hUESg+BkEQOvpczb7RqjduXkzmFAAKeg7f1WQnxhS9IoF/w
3bkS+Psk4jPmluOUHp3+/4eAjjmofaQKEw6EC+S06KwHsKBHJjkS7NhqAP19a+gC
n9HMo0fUmMGUzRh+PdLG/zlRxQIEZ8K7aQ4EGY9Lj+OOh0erBBE0dYMWgMDN5AVh
ZoNVMJf/eOHcjQfnkjAgv8nb006C4Kmu7Gaj3ZQE0u0dNm3m526IsOtCA2TM2NJM
YpHK7ltUb+vvvj01DA2uOp34PHzafRsWZU1W83uVHlXrOTaKvhPDzabDrwG4a/y7
yQGqN8EsVJ9CBjmLQ3nwl2TtpQHtGa0MRpniz2U+cwRyC2BquDiY8QqWARSg/YyE
11p8v8k9qBi9ZHBpOotvU/OrG0SC0VIbLEtbfeWIVj5VEFC1Dgk6LHjIuvH1ZXa6
A70ernlOtPP7YV/czop/mZ7fzUbafAB0sKysAGumZYWJ/bi9I3hZ5CzzWdOVcn04
hFcTDhpgsBhrlVbwcm7PGiHpNUquE4UcrJHA/6NNWmuvuQdktZjpplKzmZFWfXDE
uQfcSmIlOYCJmt+65H4y6w7L7T/v4Ay9H4rIB0s1suuCbFNhpqa/xWGFspM5b8B+
TI4cJnpe5qiRGkXEdpsJ3hIjd3S/QdbnWBAOZRrbhgIoJE4rMFHL7pb5ZDkdJ7XC
8Ky8lD7UHC0EBP2Q5ArLFZU3HR3s0dSYdtpqFt/uCV6yCsPerAUh6DqeLd5GIzgj
k+s75bat0HV5NKgB1itY1duiuE6USM3436jS6pCTabp4ZJSR4HTDtrLa4Fg5e2oK
kdVF6+nWAamUvrPB79Qe5bF3icKWZ7FvdmyWcmX0Q0Q7X3Y4BISKVwgg+kzzGCxC
WUv4JEja9DW+CNGx6PK+8mwWDcv7m41AgtIArl857vEN5zrsYjKuguSziPupfUVr
AZOgQTV0RbWL5HBAX3JMY6XKr4eXfnOTk728v+6sqGpJizMBCnjrIpnBPhlwgavN
zV8PC/FYMpLGnBXoDuf4ry2fwzUd2r/5zTe7cnSikbdK/tti6t7esiDcGcYMN8qZ
N222Ua1u4DUvY0bWdQcteFJW/+WvO9JU2UCgpJpESB/JDTj1Gc1hRWOSRfI9+Ova
ahQDKT2VxcIVW3w7XIOSEmel4leODsrvfuhnQp8cpwVpnWLnpbdqgZgfZzPepjj2
p5tfwvqJD1tVgi8Ob5UHFQ+pMVmEpTL2fuaEIDWfao5mwuUHTQ1hd2A1eqpmX+q3
Ry0vB+95pOhsI92Bs68WG4VOytpl5HZ2E0KZqFAGciaym3M1JFwxu9SeeDanK6vg
hj6wyKEX7mB3EOWzdp4eVau2d+/EJisXj7ZN7TU305ZxbLDf9LfNsD8IUfLXLRQQ
1AmyhkAibnu6AvcUq+G1uvOerMN5yrVJEZvKBJoEFOMuONs8biPO0JYjxAUngtqZ
A4cH3iFvmqcHJKbsKNNJBy5OGReh/w8qWNYdELqRprSk9UHURjs2WKKCO3ZHRESq
l6bkV9QAfbmoxyiazsysnAWDOjGaAVDfpyWgYzC5UvwSc7/LXRI3enwGDl4cyVgP
/4CFHENiYBQVNgWkyd56OzRs/eVngzuQsJA8SV2QJaBIXJ+Hge8z5kd+Zep9wSqF
BHf1fow4cagbrphWaZUIzmSMrLl3kJD/T8dxyT9Zy/ZmF63IHwxnQBZu0Od7SMXR
KuquYQJGSNLxYcfs9tcxu2EwCiAx/0dg1BMTqJ6yYptW0GwygM1lKfo5ogW2YmJq
mytoW2L0W3RX/sxUl7oeDO1FbdVu1wsNbbsTeDGrfS/p/af3DwXKT5fdFaTE5LqU
FgOcEktVXUQFiNeD7kjrd2Mxyah95ghiG2gOzaOeRhfc6m0A+p+z+LDcWvcpYyzA
KKG/hMLEOTSdfq0Vqr/maHDCU5LtT4iG4dadqobDRIKnIZDy6koaMRecNgpsCVLA
S2YKTpdE3vDUGKOOB1rD03xAuND2E5DSIrWA/SE4qbCpT+7JxI+LSE2jmmd8oWma
QfB2dc/DOVwhuUq/LH/2V8Yj4nQIY74XRW3+p9PSywLbozSd0H40MHXIXUFb63cG
/9QXsDZAvEyjefmtvg0Vj184Tlfalzh2RQ3829OL21UmWOzTY3SXVDNtH9D3ZQen
YvXUaCALN8oaH5+6NLf2j5RJBdHEkFoQeNH0pM2OGKP36fUxCpt8SUwrBJhkY43g
lTG1mSzuFoLqlfn6/YJXI6AluvG9N6zOiLjR8Ps17q+f1XonR5+SsOZGVU2lDgpD
Mkl1A7K/M5ewwwO4FQkQsOa3+dFjj1zYP5WJo4h4Khxh8ABcFcZfisDlhELjF5NW
VsczglFBQxaxXyvGaRY/8mVB/0YbH7LoB2hpTrhdOe/raA2CIHVrmpNFkmJksSq+
kZG5CwEgig3bN/5gG6F/Ken9r0EsZaczhCmT4rl4MmaB80LhSRFpBrZgazCwU52z
xeoCyVH4w/sqxY4Qc+hzn/rnhfeFFM+a3Okv64xbvEkKW3vcyjHLbfQf2QbpRTqn
JEVYLxnFXKZX5HUBEYGj7UptzHD38lIITz5ZzhYyvxdVngcBEejHz+aTpMaYKSav
0J81kf9W0fcKmWs7PS3cKpVWjzCoaSbPGyDMiwiOnypyTN0bdtYJuY2+AsqHK4sY
hceGuixya3D8UPBVZ95A0DuMbegE8vxZKTIx47qWXghmmTHRCh4EZ+WattfcuMvM
tSauRE6N85/8FI/DPw8u5z3U46SIczq91ncVUGjzVMdPHB9u5ND/K+1aB09JCdWh
eKhzKhduzKRkiWi0FEBQ9aiWyMsWU1szAxnT9ge9WJuMj+UwTfS1pd9nl55jg5yf
8jNP/CBHpCWZLFftetgrZOvM/llANPtgFoXwYhqg5gQZK2RKAZj3W5SnB+W4u1zZ
6y5lJPco9gZeQAXg2ji/W/0LdHiCdFHsybry6ss7hPUJby/nCDDunhn78+0G0nEZ
V/fcdSr9nEx8D6WWZXaJCahLqjpJnvG+v9OTX/qOUJNcyQ3qiKML+D8l0E2X90Jc
R3yE+UJoWJO3xDvYgTWZxJENESQ1wGwwEHJTM4gCZogvCe3sRtimNbST9ozG3Qwr
++b3j6XuqK04oHTe7T/D94K56T3rgBt+bpN8w4oOE+PGJ0xlpPW59CXKSL336Tye
Fg+35GNs2EQpO4CThd969L8PawEu1MxPE3VBPbhsVV4KKFObxdzyBtBoJ04nCpZP
SPt6I7A4q8glc+/ih5t7aoNfpg3EKzvJ923BBHK8XmKKiOZhiwjiui0DhBkQtoIm
TYInRPluPYLFmhyf6GrFPUyr/DJdADQcd9Rl1LFhvL75ZfeZEI/TTX2IXVQhczwx
gPNphCqiwJDUyUeAhvnL8KhRdtODVELxh8RccbKjDIKk1EEevL9oVnGVfHXu04E8
BzZ3FWvuOarLZXaIdjXLnZmqRmp51bFoDtbecswh9h7U0Lr9up90AeTRpJFvqMc0
xxJAMKWAHoHRPN8jnoX2a7NjjnYP28XrPAWxSoDLO3Pz6sicsJWb7oEYGLd3Dz3X
oPjOV3ZXfGHpLYK4rWEnnNap4YUCVVNxld5eO58hCl6nKyyswm1fgaIiHz1/rxuR
jf1wdIV4fAZLkuJkIuoIdl73QC1GFtdKbrqG+OEy5FZhvcz2wHf7tXVkQNX30iDr
lcElJ8jE1yYCJUjL/omHHPKZH6ssP/l5ZgcOAu807TjlMZyHs0DnYM20lN4bHIqt
5GhvUDvZB0uYLdEsCKKZqEzRGdmT7bldqVVsOmKATLFuAZthUnxkFcRRXioB894S
b8ss2VVFn7kginAIMg6NtJRSBzORTgMDgRiT7QiE6sg8zJr70wqbxYlJE3hGOzBL
InTkG7ulxCcFAI/jf2+IVtIOr0XuGXe0HOCDOhr4mjXVyQJS73RoimIvFv4yFIUf
3ULY6x6BTZ7f35w2pAEqfAH6/h/IT4D2irQarue1XtAd6yckeVQwGV1wWQmp4589
p/MNp4t6tLmHfCErt04+VD13UEsA1Uk+TIQaIUW8q7vYYCV/ymZ4B9Mq3hVD1K4C
+k/PI07EuA87a8K+0Go+3+4hrp3WbUO25PkUMaYSGORbYvo57HkmCVbq+/DWCRL5
Uq77kAmjtsfguaFgzhPBcdn8OFAoSgmHcnPA+vvpJbLUipowadfUOUdG0yAmvoys
+eOX2hKPM3wUC9VNXnEWFepXmaEC8xvoCAZcEPok13Mbc5jbL2NkI7BRZYxpq1kO
/n7HzQEyFeWeoBPcYjIDDjND2VtnglpMi78CKZLNIzG19U7FIRF0eqYpnEYY2N9a
ibqzjRLl5MsuJ5aliGF4bgn6T8mZ0JZCaj2AYOPpAth5e3eMG4/OutVnbzTJ2/pq
LUgj2KXVuHP+lJDsq7PyxxvUaejmgmrFrqvChtcRvtNm3+ZF0GGL2v1cdIkp27OP
lsEK600Is3F8+fVi9B2d8+mh0ZE4m7AFByLRXIvLQNjNBJroqE3kBOxcStGzy1kL
QECy2VKTdNy4i7aQGu/p4yYC6ej0YM4fB7bgz8lqKwyR6FYY9BVg/kGdZlxKaC87
qfnKF1JNbX8xwnVTAf4LKLiw3lNjYcUlahqaEnhZtbTOdmRuST7//ed+jBqLGPTW
5bR/dsp24UQpe6/aH1lDM+TiTljplS9dy0mbsLduXZyIp8q7jbjQCFf02IL6S/nG
T2P9SLK4rIGabAzvdCIYnlWOtK5q5jei2AoKAl/Z1nC/b8Fm973UG6zlyIfiPuCv
nBCqYWq9a97ZHDG8woGU5vkHSxE5rX/Wjbum3MMerT7sddw50Cjsd2vd3qTYKkCO
wQYHji5usYhz3B7EMwbxIZhbIo6FiktsBQeYe+30gdEdCCbT/gH+dPzyy9gU5z5Y
K3xZNJDlPmmNO3yZCNUmmKIxIwDgURb+NL2YazGJKg6uXiTlHf+xI3B0PDhP7vP0
1Cl6BpWE5Ev9VFUxdOB7nBW7zInVPx/KSBFVa3kd9j9BHs7M60PI5PlZm7ae2H4g
7xbWdqauV5s65EaVNhi2Hx0FRY5rwRiUvKY8MlxuFefwPgeRCtL26/cI6eLqkl7g
eVyen9nOjpVOuuwjUXklEKeA69vPxpO4cNagpp8DvQhoxgJTfjO4EphAzxkuoQJY
+wawb1SsUCl8lP79yU+SZF/Z3na05HVmhghAe+5k6k1HuBxU8d/X+PzoKeflTBQO
jvClXwgFyGpEtXjXtV2Pjb+ddqbLBSprTl3AMWVp5jzqR+OaLtQ6Jvp8iWz2GyLb
esBpCFpvPW74APSfPirDorVvN/XhmS7MduX34joqHzVGAs8LCD+RL157dc2F2cPu
56wo/1ivLq+sZ8uzev5wqsT1DvimlJ6QiWCZD0su09AL2PpKabABJ2UfssrwOMQx
qfvYibcilF2wDckMxJ126v/hx5E4fKxb4n14TJd7+pjxieqRlUBVEkDYcgVHZORR
Br5yRhlluuh/t9rJsbPpP1VrdSSY4EGb4h/5MQWmu7dJfaHaB3Th9IGEe271KXH7
o1xGbmTBX5rc3ae359fZmT9Qo49LsiskKKNFtK4bNww6JMn/uOIClTuEn9aEGKbN
+237RauxKDj3JUkTBvP9VXbtTXR+HCDW+w+p6QBBTJPF02gVAYT6XmhKK/1IXZE4
+zYvtCcXQulZIkJHauZeW2IfSvOUKkVqSlJctADUdV17oRfyHFYWPsq1CuIWqz8x
HhuOSL04ms4vAFfXGuEwlRkxXHjY2/My9Ze9ySN+Yr2nKG8rYaf62HsWkd7fduFH
wwEqWQv3B94D0MwxWvq3XQa0WJfovaLFtwEc9WU+wPvPvxjT4uUsoIdeVmMcsgMl
4HgIJeHBkknqbfvxeSDtaUSwljr540y+BxlnsHc/v10qZSHE/vPv0HvOpmN1BJlZ
yW5+BOs0eBGGhiX5IcHEN1IR3+iq0leF4Nh+W05lih+trnvdcdAoHiTltr8wVcH0
wri/TQv4+TKHYmwJCENKtVHdlF4h9TIJPkIhSB+4GvuYh9tx+opY+sWis0oXa1m7
jbBs/fFTwCnxFF4hAGo+/BQhleeeYp3U7y6ZSW7SUNSAyu2xQCyNa0l5HaxSkxMq
FDuKqD3J/LLkGSjOYy3JgP0LjHipxSmYNPuJEJcMZPMCKMffpzp4vyyoYKSQp6or
oY+fA1XS+6Oo8J8yeNPcEfQOkTlz/i6htY878HxZEKmdg9hVVmO0DuLd2SmzE/Hi
1csYT/wMfIK7jgB+Abw6a4uFPPqSEgt85Z0vJWWT7D86UWtg6OFVF0k12YdskquT
pO79atro676n+go3lyaKAqWsQmdUVTyVgOlHu1TE5L/2CoPenW+4teFfuA8akLwQ
tS7gBFcQfa6O6vYG2RFoz2gTmyTVFO+L1geOFwfcODSIA9NGWmx0I1Lo+2V9dioU
X8k8WjyvbNAZ+WWGgbHCjxjpO9Eg5qofZTqc0mE+xTo8/2L/IwHJZgpanLQl4F6q
c+QdN4nmNSRN6Olj88NWSZGv1/Cdt1GN+ArPMOyl90ODMhiREAlQ/FArohU7zIA+
q7Q0bK8PjNuqhFIjOVhlW522xNHIieNK/r9SmoTjV7PL4PtqvqsO+pOLYl6jx1cf
ZmV8g3d7F96o0PTJHVQ8ENwcjoES98N26NBrcXwDcT2XgfZ2GrdTDQbCVuTJFnlV
D3DlAVVHl5kqDOvPTtvGvLUochMvOK3BvhmdqeG8qCMVz556Md5lCrr77LinPhmx
oAZhSu/IOjJTvnwM/zCF92ZG9SOy+9BPXK/Yo6/YYzMa6Ca1sH5E4OiZNLhuTX3H
Gzcx+fE3yvkyaakuA1ZbwXOQK6IDJjbkDyvUUvqidJHDkSL1bJAW0/c1OkfTgyme
XBv7eqT/Eo1T1mlLCwgII3I9OCZqNygsaXpvU2xYv3vIeo33lS80KAqHFQtklOEC
Crm1ETAzp3Spp8HWp2DtutfoLTo4zlEfr7ecdQKn3xaU+8t40+wjVo2Xj3D13qsL
5jE/U9sb4GG6Mq7U5jF3sS0h+ToTbc2BDgI5Jag69mVGhFy5GEueFF+LIlrCSsq1
8ylrAbKwNrQGkiOlRtq1s9GBBBp+gCECtir0NDrfEPM+3pmCHAfPyc0fLE1PPtte
mZQtpKL4s6P8Ezfxur9BpijKc2krBRl2VmDBW8Kr9DXm8z/UePryV5ZQnpIeyHJo
cRuLFoXt3F5DpDgUyvDZ3mawAEpNuaYLyQ6BxucBlD9kus7iczw1mR+GzxVfhLFT
rI4MA1yKm2fUAC/VP3FWOpj8vweNbvMyTpOAEVNLQ0zl6dAOQkCAfD/+xv1Dpi+x
duo5JJNKPYMOrPvGHe3NGxSmyOOWxsWYKd96wwFW01j82MyAXQLaxHzvOEyS+v4P
JtQDd8kGYoCoF6Za1Y8t9hXkeExf1JUndQY3d3rAn7sRbo83ztivK4qnoSZUPEk6
PBaGtLPpxXlCnhtHa+kDTjqf45sGi4h6EKlhcLkgx5v8lLh5NhY2AjsMVUiFEHVt
nPpP5VfdzQVFrd5vyxi80LF8gQkV9kHTDPmp7shslweWTrAmRXEOXTly5wpSIsBW
y8IXC8Q0RKAK6sDpueGJaxMJYCSBv6of2dnXer/Ngn5TIv86TLGxBiIjRsimD/WE
uiFzBnA53r0K+/tEJJJ66WkA9KKQKZQY7VnT4sgUzVu68X3Ibp6EkEygVXNvEHDw
EBWisuSjsiiueQReFkbmBdTegAiv5hXybdmditc0Nn019v8kd9FJKTvfcGYXJQdf
aOL+iE/zeoge5xaHzc+y8DPkfD5zwMe7k8Qri5ykMjiewaV1XRbIjXaqQBE6qalg
refL1v7jc91wlkwZfHdzEsrjQjOXW1zPazdYOQVlSv/4dJmgfzWMsq2HnFq9qBWy
UlgDqtnccFk+ulBaUfCQiMwZNwYhBKSwvB9w6OCetAt5BbkTcxtl6EscWNrERmIp
25+w619S4DnLXpMuD77sMTfqhRzPdzdhw6jDoYXZerNPPkywahVPs+L6FxWkqqAD
y92Nu0rx4a+mIsgXZWBsN6drF1wl1RP0H7rOLQrwE3s5m0d6RkyOdoDPT7R6Bsph
EwRdZRJY2b9+8dq8A5n4JVkk3TeYTOACP2dqqAM9R1Ufy1QLpv6SPC/eRsvzwL9M
n9ounsV5IiNq/LLPSwrUv0JuJiaaSwsnfmClhhr1xFP8eupbK1zGmPMrodoYCqWu
NW+4cu1//Ze/sXMlbNWaS0n4eokjtEtpXbZ/6XC7kHz0EPEIarDR00uYR9yRlkRs
ISSyoz1vnv16ywEeiqIxEeCwfZ98/HJf5d4H8I9cfJpNG+BOK83hC/MrzRZIUUm/
kPWzV8IDT3FiHGWQqH2yiDF1TLwF/DhCwlVplM1kevt6tjxxaobROdbl9TPKp4Qx
FdQDFzc666ZFUdTs4boRY7lMA/BW6BnauRiaqBvoAPpfv/krSbMU4xJ4a+wOXIAV
Bq/jM60LEB/oXeT905KKdmqEWYx3t5TERlbQAS6zsLDbxaLW+esDZsWzJLEAuBB9
nOUfsYe2O3s2IeBtfNnB8FGeVMN80F8a4gnUVobgm80L9DBen4jj+PNgS8OyTcQL
I1q8bGeY4QoMzMqfxeLvxCpOoUPJicP8n560lAjTnKXlxBFO+Zukcwao/QWI4FOP
J4BFA5eeyXkiGBmOKfRGowbBTzUX8koAJPV/aWivkXSJkPLwwkVZO9hZ2j7PGKpb
pjJVAXCgtzfWeSpD0sBBTc4x4BDHMkEdJ5TFQz65cddaESCOjS7IbQHBW7Z5pTFa
55Q47VWw4R2TO4RBgrSt1onVDcb1obQSjmGRyJDzySp59LfSZ2SQQAkhdJnkoP0Z
oyOHtC2IRSyO0Acob5NCzB5B2v4WnqRf34vqBeBM0SNkI70ijy862KtxSUcBaLlC
tHXe1Kt0eP64h9i332eo0TD0Dc6uTCoOQl68p7tED2urOledHkL/V84aO8uDoiom
zqGZQRFQHHGKukToxmd+bttSh94r33aIQ8O5sanSk8L4/r+FJFQhD4dtInu0CetE
FjQzc6r69t6axTxnWM64WoJY7pI4gy41izoMBpODP0lPlQzCCcqvrd7iEv0LoyEz
0LwERJGg0lORgbs1TKf9fDyq4XKbjBbjtiQdwbNhkFRyYe3CEKGpiJCfIHtvPIIu
9Pqsn4Yduee5Wqzwov3rtZcVtb+eer+ffUP2Djnp3GO+LNsKIQWm0dbMkShvbHXf
fWH9QVXXgbYezoCnOawiAAPp9eGMOsVbeZzSwjXFGGV3OJFySLNtxYB8JpsIwoiT
1zmJ6FiHYuwcEWMwvwO8MT8/VlVSNm4sZ3YcS1bmjg6XwubO/AxREOkzSOLlYDEq
Liw+uzm8M1ndLhxK8zwC5XTd5jAtF8QsY/6dl0nHpVLP5lP+j1kH219bRlgFHLB5
3saJAiFLMWPCJYGGQgARPb0iDmuDyheBv3IYEcwc9765GZL840QjNXoBfpGj+UNl
tPJ2C0g9Xnl2Oz57BN+NymfA5abs16s8RVPWIajIJQo5m208kSknCEHayS8xiLd1
N9d1r5QUSFqcibHZkU/xGC8AGNdMxFW6dSzAHlQDPFqI4RIG1Ewh8FxqKDIJ9C/5
pnA4HncXbZtDbKKYDew204mcmuhgi1u7z861PbOn+Y/5IA0nsQPazo+rHG0fhMTN
k7jN+CnOMU4jiVo97rkVmj6+Fa0mM3D2gr4BPMcnO5Xl27RJ+tkwttpq0EDlJlsT
Ez3DdYZrTMSihU74s4hrzfBoLwHjFNAPccYlRbjN42RQHMYp8WWdQZRL3WykCBAh
0k0DWnQ8pXYemVp9vosKgR/g1qLsAQXiifS/ET9WPHW9WmmPJP/4hfSH9XWKX9eb
VOptBwDQ4WTe6RB+0SA+pQpZXUXh7/Rtb96nVfNgRxy2QNqMRUElqBtT26uKzisI
F0rWj/z8hDe/XomBrMKwbgjz2b9vBJHSdgXN1yIX/M3TvSI6h1s54B/mulAkLQwY
iMNC5N0UQAXLli3a0kiOYUdEsTb9NTip3QochWbkqHWgtoU4NdsIfgqcmE4+oY3R
tWehl/2iQQVVqI4ICgE2tZYlGHW0w1ijbjtJvBwYoBFj0lmk314ixhFNsjJuUPyI
FWYz++ezCIajTKIiNOqZLKkY/C6I9+0kiWbVGu4kM7oWZl7LfYmT7Vno1CudferJ
lilRrTd8zsCS6sYPDC3wwk2V4KmnZGmN7V8YFEdBjFoREpVoOsQKaAS0XqerSFa/
NeWSOlre0ciWMGz+5s+HotfTXJ8AinG8CA90GlZjHdUvuOyCupdMS9gKFVJKsaPy
U4cw9KHGZ4XRDbKse2GF80SYD7tt3U1HcdK5LrQarl8pYR7EVmHk4vmRYrPC89/j
0oLQwU42o1a+uCZY8b0y39zHUeBva96GKhE2pHHWz562pIdM3a1UlJH0Z4ylONI+
o5jezo8qdR2qHwoswKuMF5Ix8SFyD3wRs4N9tTIYrH/TC2lTIHMhuohR9xb6VpKu
jt/zEA/rhLvswcTxzlg1BC5lPCjKvwOahlMGPhvLPxQGn/f72GDAaRj/jogun37B
eVULOa9uJjoU2mbIotcwYwB50w8ch0jfhxhjO1Fh84MObL4IuZrjW3HAvrRwiSbc
07E9K2sEo9pwEwb19udIqdnasUtoZ9fQQmyQFQRrqWtp4ZCKjpReioWQUh0jJGqu
PmdotoPh+Vx0SJunu785PmZSDC87dx9iDdrcN7KBa1c0NOwn3awa9W6YfELNy9LE
CjbmsOwUQLQlWWC7lsWVzEonZh7AAwaImvyVul3QHDkW33xjiKDRFpGW2pLh0+vR
b/8auPZ0+Bn9+wgK1+anwchCd/C8maJ2FiPvqLLpXkyIs2TcXr5hG+bkh6PlsXmG
vyuPTD1cgtbjjJaCRAwFR5NCCKAFDoBkPpRfpFFUpoY3xlx24PmSp4Jo4dzFXO8H
IzVbeIJX4eQ7bFHt803JsvlPZQaY/9bffOJdOUJFLtHibi5T5zCGBT/Gwv8RmOZY
+HzJJOMAuveto3D83TrVr50qS4AGJJ4X16uotvN70CGXIKH3/avCHu/aKB+4yL+m
Ydg+330RMCO9RxWjj1mV6kHXTnTA2R6SHDPy1Hf2bi2nAT9WyQarO52ya8v1Slqa
D+pZnqhDLZeXiV1QKOH+3Mz3GM7dsKwFnO7LeaNWUajZifI66Tm19Fw5HHQt32Kk
1c18rovWvvY0fFw8yVriwrE9tjc1MD9y86ozZ8Z0HIAHT4NoO8hXTSb4f3iIvwaU
+Yipj3ErTKwVjWRMxhfl2kcvY4U0roPRvbGbtd/xZbN/uI5sQG8T3hDQNfudb0xC
5DJsIDBbfCxcBjo/7L8y0Foxg3YyIjCPaazIh+1ne+bFqL86qFUodVDHEJhCqFgh
OV/JIE+wfGM8I1UMqTqX6pCKCrb3jxiQ8tt60Yq2FTXFxH4p7T65Zrn9OHIOCWib
MXFHuYI+USSmceBqvLabiL9ObTqrvGykrwK3pm7j8brqJNCc7WjePVDOIXJMDtK1
DDRT/YZ7BpVtklOiXLDkwJgdxhTPJlV7U/K64qH07xdJ6gm43NWprZcyvmV+K862
FiuvECcoShCbVOaMtWLWDbcBRbSYrBIq/8Iix2bCvXE8qUi+4ngiHdA2AN2QRHKw
VpJGBEX1kp4T1Z1I+9ZBHgZY1sEuaWpgzHpslKND4esJ36SkqObZ2qdPms2jsZlm
21M0LRGSStMK4Vrl4FrLZPuHk2e5oCT1omSTRrnRtF079UAvWqzzjoM0yGGuApfB
d2Z15Q8sPt4lgVkRAk3qpIAY5kLa1EghKo0lhoJU66uaMjGHyBj8MubqRCYvn0QQ
jTPehIepsZyjURhAoO6fWfeZlzPARiZBNN1oo1fkllxTNx52Ixut4AyXaAugWSge
zE0Uwpdoqau2qS/Hutha6p+LvPt4fG8ZZ1md5YAVgnz64qh6gQ6rAtl8uRfcSPZH
TouN7pAZrQRKauiCr8B+xaNpCISyGEqIrVoeJzKVISNApAllZP9Vy1IQ1ii9KJ7L
ysDvXc1mvlc81EjG0W3xqFGRjPpWrQdqiniAoa62TtsVUlfq+F0MAcnRfXE2/fj5
zAscxD8gpKsDeIjdy5sUtH0iVRS//hWs+aKnyhnWe/BbQwUzkaouOc31FNqngrVD
7HZIvSCT9Uv/JEnJ6DvO9UWGsaKfPZdv4zozeIRuz9IGDz9ZcmSDWXdFdR8XzPUQ
Z7lDNr/oYSWlO5wG9mN4kMyaJbdrwq3FqTW6/xVOD4C7phkSW7zDicAECfJYKoDy
R+PEscoP9hM3xRCb0NuTmxqI8w5DXBtteZHvo6Nkdq8/U2wPxdOSbfq3AvnrMk2f
TIp+jndNd8r3++Jc1MdM8LZB7NeXlSam69aW1ik+P6AbnklUadDvg4F7h6EbgI+P
T5Ng1ly/IIAxvScqvnBSbqL/kK/hnD51cjysdbQbKmxRWWoniZUrXSGC1zYcvDAM
sAuJ5wTnCguxZvxyRhuYbac0CVsqMT88KXnRT3Nilrp6sG0raum3os5r84RExI5H
nyytkv8405YZXc+yVWFYsZhhccsRPbJ/9eUduJ1N1zhExrRJ/7dgSxIJruxUrQL5
bPpHYW0SU6uyuyiISND26+UJn9NrxBe3xf6PbFZuPDdTUF9Z2ObOMMdI3mmIOo4b
YoNzWgqiQhW90UousmdRdAT+xTWN65J5CrILj07BWS6K+pwIEkOeljuEAJLwTg27
3zQKUQ4pTt4fMCQYh8ik1UjlEALGWYs86xztG/uw/dqIVkiVDBSuGEc8C/Sorwo1
ZrPN1h9p/1WD8KPdcXkQFi/QgonCIQTLio3pvMeka5PkVMu9u/SdyLLADLj9fn+b
8f8XXBKCDQKnTCcYU/X1EPWnKNmABKdmZb8n5jCHuOsUljnNopA3KXqtteCmn6tO
h2nMMVCvzuF6xF+zgEs3TszHwPx2OXTG/pF6tL7SonOLIhbXpPQG0+D6Ujh3GUhJ
zFu2CbMgoEZjw6jsijkxGc7xbPFKErFGwd40BE97u6pu1jSGO71axYaQBHR2QIbr
ERVfTaZp5kwoQlVpOSt+WDKpdNu32JrT75NKdXp28pVGUjYzKTTKGiVatdJ4BqdY
CiezuN/9ooBDvCZSbXXadUNVHByTWn6ZtmXgyKAKaTy4maav0wFL/MwHi/+X1IRi
uLHOXwjJ37+FDVdYG7Oc97omN5dpmwwhDOrdMPjYTd69X+F2yj55OAskkfcmUVfV
P0x9nYOgeVQ2O+1Mn3KD7APuDTGOaKJ2TKWsI1SRmmCOe/ui8yvCfsxbpw2rGsBF
aUBSOXlJx/HT80HBJWLrP8cuXs9HfdVSu23QedwePJWCc+dLD+Sw47Zmoe+JlUsa
dmLbkBXd+1k1iLWqutXrA6SNuU6s3Bt4jDKXxLopGcl9wgclBdS30Kv3wUPzIQZL
vQZdY4sRbe5kDTKiiGoa3Y1z7QdjSmUdWy5N5BRXCpRSe0Qk0dVo/MS6FRCcJKIu
fXHdAdHylpGTyVycfK1TCFNa0QJ4q/g8RioVlE25luMKau66Pjs5GBwlb94/KYe1
rEPakW87JgzE18aKg3diOkDTflbzFYfVBf/9p1NITcGuCNZtwQ06yTxn3g9KGbhX
sUEczH6AOmgsJce8gEhiw7ia/rJ7brOZlqozzaP/dyP5mNZgDVh10JQvl53oXBdC
vSHCu4D6RCtj66PwbwfiL9JGGcLGFGcH/QTyfl4elxuHHbbZd8juXhooV4PRXzrY
y+7d7rPCBLmgqLG0nEGEGs8ysDn0Xy0DIC7IHiqDv8u89uNBVUYjY3qWStzDTG4b
rJAUtKAWvf+esp4uq2ze4bxRw8I1LCCzNd5bQvUVgDwBISKAhgE5+KSL4LMToVWU
7hUyMXCHPSqLWvgCA3PTz3xtxQV5+bgBPtSihgt9SyvDQz8MFSzNi7XVihFqbIR7
7e9TddO0sT9ePEoqpxcuhFeRnDMRsxhYGvjjXurTWd+gKkyEbdrsFo1CeCuskqUU
vJWOQp5H6vbQhvNR4m4GrYNauHS+vLx03pg/Fk2okK+tWRbFrAUELswfJAdquNek
dBfVj+1Tn86G3NcXa7pORVIonhJ0M56dYJvYsVPyNOMS1npDr50w1a+S7ItuQKGk
5hpL9Ehq6+lkJGwyi/NlwyqjOzkekdnqjn/hnYSEvigyMA1Km/vTBUaP76dZJ/1m
Qx8nETmN+mO3Yz2cKprIJ4w0OjZkLM2478XG4/6kNbOeOdGYmiTvsx7pQz67k0Ld
Vn8hyrE1puAFYgHRGZFY0UU9vcac4fYXW2MJyaJEwclNhM1iJsZIlzkLNqPwxTq0
WlwpxnPe7DA8R/NPlfXoyitiXDOs7e849tatXRaoU8Q8srHg+zOwmERlySqgB0ml
OlwU0e2P7r8jGGiqfbMy4OdwSMfw0Y4v08KNzLhaeqv/1QrG5ZqKVRM5KOeI+OJ1
KNNtP+me8P74ItmgUPQi9RUU4MY8EcFXMUG0y5MG5n5QxycenX+CzqDTLxxXh1iT
c3KZ7tCnC5BvdkaBeTnK4py8u1OoMDoE7XbVltiYqJyK4MudpbMv83ixDLN+8lHu
uEu0aQKJSDEOIJ01J/hzTCwqU6lFOweZYRmW4rRopDsLvsTWoK7uqO32Gt7dQmpI
oHVWR28ZhjTMTuAdbukrerEkKLxesDkuZGv+zi2sxV9jtIWxFQ5/oYn+Q7QzqXzf
K8tCGRWbgEdpaBq5x5/UvF8bSw6jDECe/CKgdei+TAUoMk16B7zOSPPUHpFlnjuO
LmqUTQtPEqkJI3ofuU43XThJqTIYGnrnRBAnObZ+LwU7WRD0uH3Qm67hrbgSvxQW
c8rWARS8KfiuDA2jy74r8w==
`protect end_protected