`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 29664 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
Ju3IpcJpVj/VshHyynUPTKDmui7WogCcIH7q/iV5KAqZMinF8qxCnlINoFTczA26
pns4UykfxPt1YPhYBXhgOm0F89pFQ3PvX2CWYZwAE0rZvS3OJlwLnQaEdW5/c5hR
vTjYuAoh4IKk6T/SWsPEpRIKo1vTpA6NaDxeNMIjY9G6fgo/wCKxSWBLX1hqZr1c
MoBKgXEr5z1pF2EJKLjyjNA7zyWuwgGZNxzQxv8W63VW+xRMwRYE+RbmPyYyb0qS
GdF8K7xyGhzTPnlTBnHM+ZMFXDUXCBgZDU54JbfmIeWsAI19jKdMwCDOiCWzUQnO
E1+AyrCnB0+elCK/+us69qRvPrw7WTwZ3ZOErq6tmANstemugTcKqnwhXVM6fXnx
/C4qrNxoRGa4tmnhfYBd31qzKTnz6doBVujGRVlB/Cejdbt4Z+sr+RlKS6hVk6DI
XpruJ8+liz0Uv0LUvog6Lf/+xXApcfj7b1qVq/3KmpP7VnON+dCssWksEANVEBXY
f65Kzg8JRwcB9r/lPToVgPlqtwxwG06mreoHR6gGmpHPgW9UFaPhmvkXk4YSAe+b
mluxU6IVthb+hi0V6X4PJFRa0ppe+ofg+Rdm3LJ421tYDy2AzDyxyrP3dCTN1hNj
MvMfMcY2iCBoHDAYQjBnNxTu9eorvMJvGfWotaqoGQKyV0w6Oy59KDRlESPFLGG1
IWFWTsueHS6Q96QPzZG0kpfgFvn0/Af976SeRxkkDKwe6p6xLlm+asVXWrv/28Pv
s5F7crwzaJTD3RZ2IndEm9R8Y1YXuvbueyvDkOG3/YEm35peDurOk3W3Pw2JTca7
5XjIHQ9ihE1k/bB+Nw21Pz5QWtUb41MOP8TRQ1GzGdSiA1W1xzmmEdRlFx724Z4r
QwTY3oKCmHboom5KmRPmjygy5tLymXQKQKgBIGgPTGhRkCZykwzLw9mm8p5mMM0s
lBk5wEhanvmASW80SAPJTf19w729xrhOn6nF8jSpOFUtdPjv+T48uouQaAgk0Ltg
xph/n0PaDK9yhSdP/7crDfsAqaf13Cq170kdYxfKKsj/QKnzQ2kMZw5CP7MYI5dT
dj2igD7cfdrirg7fVWPSbSonV8DzIG52Vt/5OAvo+M1DcuKlBuXfnpjtf6ASjSmO
o24bNqxtxWtW/cmMpifH5B+DtGnKqsJeqVhPLFi/AzIIskcoMKT6ij44+GiPG67F
EkYbqasGjb5p8Djy9vvtwUCPp8tsb6bov8nVQ3T93yNohTDx+8FkNS/2ynC7YvWh
83P5uE9h5eATXEnflbNCCyXBd3YJvqqKaYFpifqg4MRRm0Ie7JQ2/6m04Cf+f7oO
wxi9LnDQqVr9wUCmM8859UBuMZ5QKeVmItbyFdiO0u4VI+QQUFLQ4bJkNf0t0GUn
IzoymSQsp5JVgrEWQk6HZCD1Du/JkEd0Tc5yjzijK02aBWZor7pC6cdIskChAPnR
SFc1zxYN7p+WaNioDlk1HgrL57JvJ6Q9upsd4fTu04H7PQqFnDDvGuI10Kw1oTA7
rJ6KNVijwOBLcFYYdE4VA9+nRl5AeNSEN2Agwd5yW4F5C1HLS2O3u0sbTfjJepRh
Ucm68s8JTok9jTN26ZA0orC3OiXUP54vnU3t8tzxNo2jpe1psNcMZwnWJHXzGSBd
7ULEqcSlANeFjTOYMOe8DryKptdY6RGGX5bQVmLYq4oUzjMS0XuDUb25lYsvISXI
tdQHXnJPydzFYs97DHxLzMllSyLH/hvOGBbR++dWQYShj++vFFnISeaNgRiZspjY
8wnhaG/HAs6u2Cwsz+LCeTvD1A6fPcGiS+NfM2OT8KsybylfBmOyMx4g17rLwzft
A0dRSfB8QvqZ19WdGZbOi0P+2qxZjgcWmwCxK77DpLO4ze5M0XQevGYP4uq3D4mj
lO7M2JN+dVaRFftofoN0agnTFFoY2KD8sdM2v0THdWnbv6TO7D+4Qsw1hKqz7DJy
1HiTOlh3mUjoEcqIHYQMgaIV7xmpfZovS3qGg3+G9aqOcsNFLeQOiFe+e+qqVeyA
5V06XTiKLRj9YItWT4nK3Z1HYFlnh8wzSP0tCQXhGy8TuyBWX0sCzL0a5qvzatoS
TEClHzCi8TjGicW9GtrHZETzKGgK6FjrobAXTmWfjKa2ZxYmNaQwEH6wvrO9zd/5
lOwYwBNRW+2EF4eQuF60yM0XKWDNTPnH7cIJh9uDRczQfj4Qb6efg4k7YxbukVMP
gPc2ecuFr9y9Zd+1/cNZa5owvtGw6y8b53fKABXL8lLf45Ysiw8OlAZllUIK+XgT
oQEYMmfxg0n1BkPfuT4O2IqDq4pNL+JNu0arauRyQE68tjI8Ur9SOcZyD4dH6qH9
tLE0q8Z6yrLz4XPud1w9HtIHZ3q6BugPDH3QWE39W1yES5/gjHUEZ5T/Ftu17+QZ
byEKPq4nDAq90ZUngnD6v2qJNVsXVsrHkcP6+GsyOLjBB1foeuUnlaN55iX3slkK
zCRDFa/nRvflezf16vZRBQ/Cirxfw6rucykqZ0ZfSj8z+Rn3Vxgvwao8jhDsi0fY
6k7L4NPtJbA0mhhioJ0PK0KR+NFYJl4L4N8PY1RmyFjKuSk84rJ47o1JNFLciHGp
NXudMecFOkcVK82572J5rEqtXRja+Adv+hFeQJj0Cw9xeAgOSSmsPPj62FrQuIOb
hCPqcDWjsVR9etka9jpVSkV1U529zXf2oMws/m2fdI92KdHzjEc/YDzfdTWe5v3h
81xktIpWzTMvueyX2HbfuhFlhG2Z7A4s+G5zKS6Jgvpsio0H635ZWZkySgqDQcsF
4mrddf2/SAvAAAGmvaMuugiT66PaN4gPL5pFzSaqVTZOFapZNdVPYISZEH6tfCRR
5xdVDQSb1hYL6hF5CHHUFQ0C6o23zvk+mZqz4ggzGM1wQf21mwjtXTZYVjyHV0LI
/vGwXabK/qLWyrQEfkISoE1EMrRhLeotbWlBR8XQKpiZwHwPpyJO83qmWb30Xxje
6jnx5z8Euo0NwaEjW8bxTW5Ej9GVwf56kUdnVIl5xjMR1YoVTACDLaotPkQwiHpJ
h9uAZ8BIh/PmoQCvrtn7a/9OZmVjp3gzwjKFoYIRgd7RtDEHL/tDAlscbOrKNYzn
SMJ6DLndlNAq6kbJj65ldZTMwbjPVx1j+J1RvzglcQ3iQclfJpVv0bJzYtFsKin7
jGuMtBHgkFDy9Zvl1gLJzZ+WWPsrWwCyf3qCLObP6xg+mhxxkVieW1bPlsNIyCmD
W8tqD9zz37KLI8yaTPXMeMQ06wxN3JqHf5AwGhTrZfsBTW3Xk+M9oq8YyGW3L6kO
xe7mO4ccwYadrZn/qVV6L6Djgef0YjltIzFrxhVIWie5mo+tTX9w6RyVvFLci1nr
PwtoYWIgyWIM98qaPZjoMfcNQXUSapn/m7a1I4husdLHttWwYPQSKF/w7e7jtU4C
YIpgLZqIOc0fCr13o5qjWIV1dJKcyV3nq36ZWMXtUdCTJm1aFy6XxjwvGdKihZHD
wjQk1+73zylrptq2DdDzb4WBdH65G8pK0bn+UcUSoeqjJfsczIIvxn83v0KlPrVe
gHOl2JW8/n2v2zfcqiqORui0bx43C4RflyYmyQW8nsK3VAN6y/djFjYgZuZs9ys9
fHvqZtZbBv5iHBILwm7F4ndstVQmLA6jxbkBu959c9kGbIeuZ1/dESzqUbkDIe57
dZnHs115xKHpis++xZs5SYPBaTGSKC17EW8hDl4ScvsCeq4NJRQ1RhYl/zGFjj44
IZmMwhTqG8+LHyvibH4msx9vAowP3JqDSiOCMIPsJYYLzAzgK5BaoOIiNPOeZZBH
pVJoUCOOZ3Q7TYA0lZHgdBlTUK+s5P/p2ZvP/rxRMntUAu3zOu7I8iX2z187aR7l
mdd/OOy/D0ty1hV/BwsqU0wKbx0QrBqpnx6D2ts4A7iRtfMWgIDp35R2JRxo2Dww
0k3+VH7yvx/hxucuD5s73DGL+QGf0h5dH0ixsQJCPD5gYjNCgRDnP52dAeaOfPQ+
o3eW9/NImcPtTFyOXlLoPt8ujtjTZbR3CA1Mp5wSAS/N5CXBuSY+X6V6mBWIsf43
7N15COprRXVK2Yfie5oI9sb6cV/c+Bdt9dLz1EZ1OU9Zqx89LFVC5jWlyTbX4CRm
VsaWESJ5BPun9w9xGgbR7+AWkJR+IfJcihT4Mp50EI01SUFbdTUpJnyvfkMip2TS
3GSFF5JF/gwGeqqbKoEsQHIDek3H36Uq/XkF4gqt72Q8HK30BuoBBgk+oZCMBrvn
iBuds3JChaWvUQKWRqKQdRwRaX5NYBHCZrdYmMFvXayKEh9LBRZQIE0uGgif4HXq
pw09WeRYqOINdo8VDzrFGP5/SL5yACRe8CcWYC7c0gmgS11zoNGlqrnKZIdYvHOq
9Vz53OYVolSLOtsPsNo3YGU2MwKxbqyAUAYKRMwFGp1rT6KXK7sCXUyuX/b6E4PB
aRzu7eYvecidx55zyYsUZYhtm/ossq14Yt1bradatDg08lV4h75rMHCR1V+qTYzv
P/nOGXNjBjzaCkQc1QN6olHlIx1AasX1BCpOmojw4BeyLyUQA8ZFMp9HnjfPK4Er
5S+YhqJdYb+cM2eWN7j6qmwmUh80DxbMsUAbbd8CJkosNxXfuEjCSWFg7/kbEmSf
soNzaQChN0JhdZyUTlZ2L6fB9FydD3UhaOTGo1AnuUL2sE8HhGeGy+G/o1hagGmw
Cfq7eVd3NrPsG3PIQ65Y6bdhL98b7f1tEU8UmnSm95p/d3YIbFvLB8VH5kp5r5pc
SI8uQtJA2zfoWO6+zBiGmuOF1vl/9Ct4tP7h9n9OXtLN6AObW1bniN57WIow07vj
79HhV1ogprJ4TMUpwrmdWv5VCS/HQNgYnPwl03HiCXoW7yxHgcWFS/tpyW/b+045
wSTAF8towSKUsxSIrx9ghD0WONt+8h/TW58dhOkgMspFea2EFLaNlLqSgYwYeG5P
OEAOFI8fQXGU9MTaDQZA5q6ptHJ++I86zN/RIiZrYos5/i3+c5NRgyi36ikQKX1U
dsHF0sp5IdSk/u9w/AnwKInjMFNhizwibyJLtTMDUqAol19YNTnUUgfnXOY7CjCH
BUwtifZuM6GKMGDIkrkpq61VS8SPIq+Z0cDhL+qPG2lxOtq9sIAezvFl+QXHMlIu
e9ZqE8SVXB5a0rbZNUN9MCO2TDauSx92AqZIdlyJ5LEyGX/jGZa6BegPby8+EI9U
GiRZqb9G9rhlPawOKQYwyE0+TFOnq0dhrcvlvnFlhT+YSiXte+bdnjlZ4QSCPdZM
/S/7+c1HGOpBnCRLhDBlXeImoBLIVA582K18+EHphrPZE6onTQfLkh5daG/URRO+
dYuZDuGXUs/Xien6tcvchVylLO/HJYFU0ok3QDsHJk9GAOk5o/8S6jBM9WlZ4nli
HBc7RBm7KjP9M2B2yd5y1uaSs5SQeRgXBVyFPq0U5FQRwKj0SljV0ITLBKYUWQvk
FIm/hWweMMeV55v4jIJN/hv1naoObaLsZtXJmDGQDvQxTETKFlibizhQcf+d78d/
x94M3lJ3T7Ex2gQD0aydTJqonf1pYHS4UP8AKRecTZyKntFwNHobo+/M51sOf13A
k6evsSpF+PRpiFPbV464h0gKGeRmEMkBTy0P0OVI9dpcpZbAaBwLxF32bFQP34zd
zaSlsA2ZOzNDtOkLwK2eQJRsOktrUERAIYUxiCClG/Y/24qK+P1XWoDRMYmtuCFg
QRfW1fGMcUn6T/pfZuprJPn+EyxqF1RUP1JSZYNvqjaELdCgegHW95SvjGSRgc64
jzusV7MS8c9daeKeKfOO/RFMtQuBk5rdSwQOY/Fk7eutvoU/Q0CGjEucENPuuI7P
PEbEuVYyIePL5HdZjn9CmDG6ZfA0N+0OUoKXRZxjuj6LBnSR/0nzqoHnngtziUJw
rmX8VSFAZETCmQ0uhuzEss19bRLJFfTopy43IbuqAoi2x/3EzNLNxDbHxp8/DI3K
Lv6KsstEdkIIw2AzXxE09fyYoem2VUmiipci56p2t/KulvIawrOq7sl8atFXfinp
P41ZKOdqaQnJ3SKtF+FXxQtJKJLVElI38r7a83Npy+eoZsVO1Yhrjimt2V52dR0R
nBXJjzXaP1DIgoM3STkKAXYcexyP1MAgpw1R99zzG11eLOooRjhdowCas79vRb3V
ED5VUWsvbkpxkayk9l6rR6aVIcKUJzNgpf/XrPmPmkUjYqutzf4LkDZ6tPnYmmEs
V4kZ6qutXYg4QOfbdcSJ3ImUnV1PnW+j6Q8jJoPboMyUoc54Eepqjhq7vY6ooErQ
E44xcM3dk5kI8h0x8+E0p0qiXCHXIu9Z1ToEQEX6kAAzHLIfg8E59NKQsXYWBMds
puiTp2aqyZPxlnwoTHBB4pw4YaNqY76zyJii+M9aGYa6DOVhMaf3344H66fRgPv/
HROWLSoC+tcmw59FDt02wMFaqR12wWZwWv7Kf8dJFuRVaNPY8EKBns6s+lsSfKFN
NyTmIsKr7b4VZPbrJ+SoW/iHeszd7VAErhn2DtDUaBobBSAoMwk4Hzg7uAYrv5B5
u5uIarozq4pZKuFmPW68jZdzE45ubMgGmT/gF/oLgER4okKmFarGkR61d2tCERz0
63gscXCsV4OsoOKx0k8OZyGn0/qwfgOzD6d2mSMYo4gmBYTHG6m3+wGKhttG5gHd
jMfhZL/6+eQezpPF8N2Y/sgiOqE6uB0JHHJvRv++YJ+WXKuXHj2wp9Kxa/WD8Z92
I92AYMKE1DktAnfGYZ9A6sTtXO99X/+Q8yF14lrxPzPDmO+IslYEayiBAvmnwTjX
+uBvwSulRm9wl2D9dEtRUl0rRzBuugYlJOei7nC6FvnP1DNUNKqKcLXTTesnw/ND
j6uGJVOVQFNGmDmCAZfi/stbWX7lcr9IYePFsG02B1WgN2IGtAO38cfJ/CDphdAB
tp5uvtQ6mjhUPUG7XvBYKFzDELCSGEI/cZIRJFiT66KNfXYfhcuteOpgXYLoQIyW
W2bpBmMbyNfKYKJdUCwbI7xmZ154WgBJdxlRQ/03ZxVEWsXZ2NwzTHHdV0lFRz3m
bcMK8loLw/QtgWNlfTnEs0EtJ3KpU4A+738PB4DS184pvdxHTNjWmaZVtvFqs+Nd
GFDuTh91DOGHn0RC520n9AAbEp6DnFiMVtgJSgSpjvVx0MDmfMmcuJTEF6GH2ztJ
UYkm0gh4huUnVDrxH6g87l0UYgWGTb/ChsZw25b091e3BQStTBAwcl47+CtccGd8
nrMWeAlTNuDkUNZGeHF1qEmPDJp1sHjmL6fUmV6OVFZ1kkxB8l1HADpL9XI4oXnG
P8NVokSP+qQA42aazRbp9255/RoU526hEhwXzO9tbQcXCf1t/XhYslBJsU1wzECA
eb44bixT0m6212CKwOOJFkD+o4KgEALQpZutpjMauwJyqFaCM0xw2vwMeUnr2tmv
Vy2Ce8iz+Y6aGlBFpgkrETLrhPMcxGHxspJB9bSbVGgm9+V83/ORZiuoHGrf4SfB
2x5gTwIq6YhaW1ukvyoqZv+XmVjtrDLLl7epkoxVDd446mBoxumeIrFXuj/3KVze
i9VUytdqBdwI5+gX03Blqt2BXQoVph7kJdD7ehypcoWLmXZ2cPr3qARRdiud+z83
WTYXsgYgogF4uIIDWCYkonL75PwmpvJg8UOxW2MP6AL7aR1AhgWaSwtOzgWEXaP2
sAS0cHhdb1JgkGPTJSPxBFKT1+avgtnjLkecd8/M6QBS6PQloLDpU0XdTLmFwfKd
pmvdCp/iwsyATS2tIVdieMTF5L34aiEs3zmgNRZsw2bGUonqxYmK9inY+d5T2L+N
l5WJt7O9JiAJiLhs+gi9zGZRh7s91nhwYDw3PVeEJxYlACDnF9YRc7oB6YEh3+en
eQoSMuYAnSpHs7cpRK/0mDAvxy7eX4/x9/0RW6p2LKjYmA6Bw9mecR00Neiz1hqs
5Q3uPDbVzVVwVzuJNLks5aYeP+/JD3KBIpMv0Pyzy5+Gii78+BG/AY/CMA5Wfjoj
9yLPNPOeIurBLr7NWOIr84f6yQ19uKMdxsyHOKR7rnsJHKNf2oUgNs+mPxAkJnia
qnUWd5P9mVa6Y5CtxIj3xUB/UgDA1qQfwr/pa6H0GezC+UNt+hmBrbJ+XcmHPdlF
ZTkWLGRgBVxovyAnMOq/Hf/bi0CrFEWHNsrpWhdUxvcMhhYt7r0gqQVP7B+6mDQc
9jwhSShFdrtKwSh+2w5tn8M/AUdCTao/KYtR0o9GHwiXtcQF4A/2yNMyJ85Djqil
oVPE0UQmg1aiian+VWCj32iEs3Jtb4WkNOJ4l0EH/hcWD+awVtIQsfHHogHH7vsu
LOvQq4pzjF9sLHz09luZcnkgZOkxSkqwn34wMq7Y4jWlhhEgndHMI0A3c4cZRdCL
H8k8Nhi+FGQas70emTJgu/Zc+PckQ90fRkEYEM/ssTkf9ZA/QOdoasAq7WRCldiF
Le+Yhn0Riqxt3D8ApCNCM6kw0B0AtSJsLxg9JN9Ha9z+hbt8BCk1GJFQy0P7udMZ
DLsp+asDt/YLpoG/FkuyvujpvxTs7hobGql9edzML8IPaPnK7sfwrLMeW9RIch/0
NOVTSWnmjWjYXcsh+jCdFHKJWaYxZjghww68mJvsSTAM+c5tInK3w19U5/+cBkvE
GKZ/86jIOR4HMQnc7vtnHzp9/6ZoJD4Ex+wvx/dBO/Ci6f4I91/O6a61HHOR/Ry8
sIwW88cSlTC2RAo2G3AwYgWR0MV2emynbgKvcT/TACUsewTcQd3GTweQRDdATKRN
/YKK5ZzfruFVfI6thLhXDdWkOVrcVCF1+P0+onHSFF0m1YiHTgJXQ8mryBoXeMGV
8Ni6mabfX37bzX1+0LDAiHAQ0VoHH+erkUwXwBLDVqw3ryB0/rr7UA8qnHbSMdVP
osQsr3GHC4LS/fHLZ2vTAhtqP7HvJUF5uias2j5z893aW4INsJp+9rXivVqd5M8g
kbB5Pg+ibHp8pvDyn/7amCyXzSyOotccvgPlSvXXbYrZWRpdqUEaHs+GqK7vDlX5
uUykFQXaB1VhZNTDCnKb5Av+Y5bYV6w1/SQwuQpxgvMhrFaVevtx+gzPGOs33Vyx
TAJqui/l0qO/tHuyYOlPyVE2j8h36c881PS6zpJ4OKBJ7VfGnMjaE1MN1m2SCnYD
c9HHl6DhTbZ/XZqhKybRp+hYgYCQVP8+WBU3XAbsimJjunvY2xfaO2b9qY4y8cRY
B9eXKq+ox2d5yyE3HG6EWHRS+vduPXDIQTPg/AjjAuT04NKuM2uLwVfPqA3HKMyb
0I2McEPAT3tKswRDFW6sGLCQn77UhaDIwyny564MJz3EFd44yq5zM94jlwv4qn00
HD4p1T0zMtPsTK7eJzOFd4/NXE/D5OGjTbujLA+B7Nl+9GGmZtTOyOZDq81FjM5l
p2TnKoNqyQvzQQZt7B2cqtogroY2UApRCh8ehw7/FNkD2bhtpy6yayb+Z4wM3Vgp
KOTPCYQQB9XEoXJC9oLn6A76yAfftODVqrFbZvrGDaXLa6L09TBCfo5DHFOcRgrR
591vfZZYf/L4NJQqUpRodJwQBYYC6IwrbIW6/jocNALO/3BrVB44Oa/khp7zTJ2Y
UED+x2R+yXk89K0IyFH+Q0zWULqvSEwsqMKDYNPu5jplpRn7PCh+8YnUlog2uzoS
/GwE4+0kG4eXrafULe/ihQg/ZCxyXAC4NYeIIvx2rca3KN/6u5FQaG+PWhFAPxx2
N9pJ1+aTbMFteZayTMo8snkCpBlSaiAC+W7rHAsSkAdWmoIXGU2AaD1JXkHoPmmP
cJOhECnt3dwvhy3yluAtt6P+oqpaoQgw1/Q3UVO/Q8VuDrLbaOmYG/ZESX33Od21
RSdexKQ8XefY2NwEjNoF2Qo4jqIPQU8RaqhhEIscFIDdVnVhuykm18AWuZsqYqiV
VpGbO2cqxxnt1JlqLsX2HhM4nI0N2FFfb14KkF2bUczVvMBFrjH4Kw8OnQ/DQD3N
mpscv5JjSBg+Qzvfgt1YjGF/3Cua4FpmhxEQi5Au0Xwe6TtMVyenlo2uXb58fpvn
y0qkg2Kf3pEdUfMkpA7ZKbk+hTnzkEJ5tIKCLDZlt+E/al7HZH7IkXvLh3t0ctfr
Fgt6vZjRXUs0Aypgl0UQ9SY31MlPqCJ6h7szqhHjHNtAaWTIS1MothQ2ztm/YtoY
xF3tX4jRqrSy0pDfYkW50dsCC5xa0cS4jnHxseNdkKm5mmkrJIInP2drayWcqZNz
zAoGnaw6CzEh5kl/Ff5xJ3DapkzA+bpMih76hp3+kuvmbc3hNKs1KN66jT7+2lX0
5co9xy43ymMko8sFDwylewlqHyb4YiPxJ0VsPqPMRy/tCAj1bpq+Nh46L7+wu8+Z
1wmyeAJM5+uGqyTTvGcpVZltZicosqt5r2VSXqw3a5zvwsPWZE393dLQ5qKsFn4q
IRhvYV+vz7mFM44royHQS4frUaE9ABOl4R74Gz5AhrTIIP1WVSWsT6uOSe0aVbzS
3C6yl7fzfRbzPXiQ2rgyUxNGCcHESs4/OiJrXOhcb2hKitltUatWaRNtsK4D2R/r
rSJKayHffHTgf/QWVTVeL02QUIIepZMBtus8VS2DNDxKZzwyifkju5tEhn2DzRK4
4MEINme6Uo/ew4+UR5gcuyYQvFRfHxMEHxYWjcWM3lUARy40lA4JVMdOIBgqJPHP
8Rpn15OpnmZhFkhwX0tQdETZaqlN+CWDAaANdVbVyhuqigUCT6i6hD5KtmMaJ0zE
XXd0TDWZ9nx/Q74aOxMY8qyl0WsHsXbS4kIwMdEFuqxnrJ2Tx99USJ4nEqLErMEl
A/2i8J20S420RtKbFcWsSKg+q9ZhZ7d9pCA3Mjjjni4u+Sd49sLp7rlFdUPNyRma
5zzR7YwNdjEdpvomkOZ8Zg5rVrXgLlvixv7O9Mr14QOrdQWv2u/ELEEvEogP5zAM
nvXZSYkhupB/ohqJHp2KmWSE6tDVDQsOZc5/voFthfT9pAcov3HgM/28YMBdKAic
YukOCdR4FHuSdopdFDqYTmwtZGbxcxyDhnyMoErYUulgusySQyJWgU59efT2A2W/
q1bp+jXcfFF43D9wAlNdnUJlNTxvMPcvS0PMQJXXzoUjFxYHPRk1+6UoQpnH11rm
r4tmV40hYQWDJNuy2BkmysOjhKynLFnCBvphlct51OoVI2Zi7EqjZw44GvZzWoOc
GRcR56vYK6GzsuUw/RGAfClVBi8Tn3B/5HEoPVtkW2cpAh2c3lxExCrGVdMXZ/Vl
PNFRMM/LA25NmUaIHR1nexdtVnS/eHL7yQhk8ogNImsxwsX79j1M1kdB8lcbq8SE
dz9HzJx4cY+cbxxPJmDywmVEf89MxUtbMjj1OlYBn9JIpA8eMZF8guHOTXg6HT/e
UCU0neRTP4cvKS0gIlCi43Su9SKWKE0AFoNfFNqsPlRjuSac/0B4+MMnntVuAGtn
XYlyz75reLeKu02II2YxNBK4psMl1JKamPV6HfOtpCANFzw31mBbNrh1QEx++1z+
HXgAmgo/ZTd6xczumoXLu0fstvTDOf0FAT2Lv+h639OWGHiLNWrXJ7O55cCefCwW
AacHw9ZvQ6TQuB/0vStTiRBIYOVgqhRVUD4oaXcGQFWGtVeMZ8HZU5nW4me+Sutw
YL3SP+2eXKGLiXtcG5FbQ8nVY8fulpRvfth/TsxKepc5RD28qA2e+vveR24+WN4T
TcrrGRQmvEDg26e5O5w1I3FgvN8iIIvVU708iMMMeOK6dQSfYc4yD5x4uKe3UF7u
vuIJUqBTxwVR4vsh7A43wT+cI4Wc7VUVax8T2bG0K/FwZvTOKZcsCVCSIuyVwIY2
ePXWoC09PsGweeFXev1QiroJgx1adrr8ctyq1+Ld/pL+NIgPVIgQlEtmy12/dp9U
NpnG/yQfP5GgEF9acXOlAshIJbgZDYJiV1LozxPsCW5H/Kg2Uu0bXDOBajwyNSdm
SUlQOhNTnofzdeMVWoDzo8j8FTLH4U3G3LHs693uEInCc9v+uiXymQLDeqJv3UeM
rIkL28HPSU6x3f1GmWKbnXw5ipEGhyHKi+j4ASROpLpuEoYYAV07cg+GUj4pZWrq
shpPyYInG2lVljUxZx1KyEAJGXvxUWfUlz6RnEtXthgRy2CXQiWMltaHraI4iGCj
nUEKg3XcH78m1elTaeSh9CRSChyoyIfbWJ2lucgtroAx26raJWAYtlVo9DSsj6U1
ZMRes4mq4n2QijsqrgNedRGgV14zewpLueNSTQdC90SsRLBbt084yaZbUOpRngC2
Nw+uJl34S/5d5BdPqP6RMFiXzXlW3vJC7u2UzMQhYIXvHhAcCpoekM0a7Q4Rrlk1
RkjXfaojJLaDoU8UsQlV/HfY4SndWgBPMdYphxPiAQZNOTWYMkpV/XRpNp1QyKIR
0qhtM4b4BW2RXowwUKNtE0TsQpgqBkY9xDYg8ITKx4j9+2HeInqL81aCSP9n5ywQ
ThqeXZIS1u5IzTL0UGTJU7TyTxeKf/Kc+ZkYTYdfW+Eb6x2jKecNeSTGIFJ5KV8R
sv7w5uhAbnkQK9IhXlPSNoRiooAro5dnes6WcZ7yWiRerjAaeMjuOpVpG6bQmf+1
kGoqSrbZDgSbvXoZ/HfbTn76n2SKVDNPabPkTV3HfHE2+Fkcl9yesHa3MVE7f6N8
Zr5uklJbTF7i8BRPhlrmL/bjI0hCGQ5n/x7gg5Vkcjrv8iOGc/ssyv6vxiwLpMLu
wvKxyRxaRRo2A5fs2Di/hCyt3dgKo2IKRVH+QNPnIXbjR6keE8A+BIUIjg7CS+3i
6CBcEXMHDJ4tjS8ly+58zAAiNsrzFn687ollCE81ux61DieR3yd2RPShbcj8AB39
MIBLOua9LfYW5WPHFYIH6SWGYcYQKJSqplx0UkkqlvWrjHuWWj16IkKmUSFQM25H
efpLS9VOXNqmSPpQGIuMvPm/hFzdC/W8poxhCs464GkyLQcBjqGfLn8iN74B5pAj
9yA+NiQ3nL/xDpKHxWtT1ue5izcGUjA2AtLwJXyBBNHmaYtgO/Jdzqat9COQmM9A
Nn2RPH9KPG+w5X0J0vQe+cvN2ca9Cei9kBp3OPdWA75S5VLe04djtXwTLZ1YkPT7
kw7871W5ogFTZwt/0iSS81qglnMzZcsT4GLDPJNP58YlGKApsMWI12VPVt4aMgYQ
seTE+ISTE6/OPZRF8xLi2c5xo/Tb9tzmZRBVeKTcjCK+BlucQGiaGoWVr8l563Nz
eorYdBLMSoiUYK+5syzSdcogzgWR5AVBNOqp5COeAwm6SkYQQqQfdDPOp0j+RRpL
UX4UJL5v/jZ719HJGFzfF1vWPpS1jEmzT8Q61ZjWw5vHvmTJWRy+VB/IU2GwKHO2
4/eF1uI2hbYBq5oUdAyQHoFx8HeVLZ/Bw/C254HttGTYlKWE5LHhdxCE+NIdvmEF
Z17pnxKPdGMJ0dVcJupEfALKqa6TZ5vDlAgk7XX+Cx59iAFsCuhN5b02b1hBG5tb
HnB/KoIq35guSa0gY8uha8xCKDatS60IfepqAhJRHValppYEGs1qAPbNC5+YVSdS
FPGHoTYygebUco+pxmjnQUX4CSMBFXejV74RMG15/mHu4lfvmKfxkc6xdm+0OCE9
1PmEPmpCMk1875hPvrRJfAbmCjEok8+49VbM+AmD5qh5USrMwr+VLnCGmdFg7NGB
majS3sSuXaXF/9BNkyTug96XEiRvZoR1mrgVPG0caprbN4VvYM9ssBpXuCn7djxN
FfT3SEEksn66BVfeSgN1vVWAKfsq4pUfbGCpSZQxzIVjkVuxX0LY0PhdYZhlbWna
1JiS+o/49SmH1yT0sWU6TAwAEb7/5N/tTNnN4XitXTwdTFSpwupOxHX1owyCmyn/
EJe1zLMk2XXGyVG8Z3Jyt+T0sU4yZmn5z+Wsj9bStI2Q+EBrOVqrETI1Jez5Zj1j
KfLI01cG9ixyubp3cL634jsO8xbmJTnE+ugOC97o7ZvAVQjI7/6SDWGAqgZ84is4
I92tXKTTJQDe5sbGz7P1LyfGXTc7uV1P4aZ9OhRhQ5xePN3Vy9U3KkNUeX594ldf
yc7+5EMPTu53AlFWiwaJBRboQFAH3YTlySJAFYyVfmu2yaky1VSj2lEYrfynuFoG
Po4HLAZn+0ExLjWnN8JSKgIQ6U4wfo5FlyZTBrKbBXTBKXxFeb4iHtiKRYAJMBZR
9rbZcjEklUwAv78AsXfSXE3AZkSKnDz7D+9EMCXyE7ZB9oH8f/OHTaRhOi0BgFOv
sjb0LM6eBqx0Hvh3eHZrlJ4EOZysWP4uN1voOI4qTtpoQDZkEYXsah7g24B92KKw
1sJSy1CLnKhbfC/i2n7RsZVh2Q5MHiV0msAE02qAeqVs0SFadE7nby+2TuKKTx5u
cm5WxFpL5ANfXb6Wf6ic/jZHP0C/UtBEqdGRKS4ziNu3d3PyEuLBfom3uMrjd6KC
EapmV1ijlvZcMc6W/xjeKfSQxU+cC7io3F242M4PXimbMdpqMA3cNgbv45yKwRS5
wS3b6tu0dqSmZryu6onvRKC/fJbGf84tMYOEEdDa1COLH2ZhWhLxe/QrAfj5vHBq
cjo+ium+PS1fM4tN26UY9qrS130LawadMx37IR7zE1H+6KqFBapb5qBOM8Gsb+Ss
VNhSl7rbmKhOTDmMbMAy0V23POk8cAU0FMR2ATsy9Y2pBZYJcisa9T17pKTdGC90
LQvuqLdwAyLKj2lvmWWiILfdZBO+iSEOIl1DszhwrzBUA5Atj6u0Layy0n6fbCu/
FZPw4Qy533Ee3GLR6d3jPcPPgKKLd91C31iAKhcpljwB1ec4llVoUwkExZcdowBF
dQ/W6oQ8PXkkxIzp6Iscof9ODD/G/RXmobdQFSHlRcgAzvV8vO0MVPy7zLyhY2uK
xmJfuD2CuYTHHVBQRx+LjfxZQFOeDkF1QGggc8RrQUSi9w32KB7Yrl0hlu7UIfhy
2xnrZZxNpVwOjyADDchpbR10dMcFIEN9BFFbuLeaYKMaBzpgsCgIVUoLEOiPgasK
eRSBt21gfq4cpqg8AuaqXXeFZeIRbkk993D+L7cjeLIcm981xphquuvV3OZ3p+LS
ua3KsnKX37llZWJMr7Myl/IaFttn8OCICl0T4WcnyZF3SLf6Tq5rM1uf6aOXIA0A
S98WRK799o9IIlEa1SIgPsig+hHsmfDhBHGclEBiV9lDS+DK3fcSTTksocsSaPKl
1Xh56ciySZ7WkW5mJbnUYGpvt94SRksF8pqVTOQX7M8C6+nsC/1AYzU7yyuasOT7
YDadWclBDlf6SoPAFqfAxsoHRmA0SzfHKDVW4pgB9pVE9IZbslVaDND57vstmB89
Dsmai+63C2SV+b7/9v2txRivlg8blbraacEFqF7POyA7V9RHCQ/RpdQ/UzY3O4B/
WLgStNolt359m3khh7E8Uor5nVH/SO+vXpePx5KeSZMHGD6FQ/08CYdn7kFADuNQ
YNe+cXhyU5hD0hI2rRJ/2kcofQ1WniOETp7l999ZfJR7hanXh0KHu/c6YyOnuqYY
nsj1OOEa5RiHDFdPz0TTqo/YFwl5WzsQFNyFDMOgsq3pd5Gu4WNvCl2G6HDo6BpW
KpS9R3xYgCFdCxTnIbURQM6H3LmM7s37MDlOgelo7P+YtudQwHM6cfO6jFDU0Vue
/EeM2HgkQ8C10Vw6+oeWT5hDMOxKeawzUj4T2PVXTKGKxCBO50ps49E0uqBs4vl+
DrfMJdM/tlAduS09pDynyF1K2UigIn5mJ06ZaWrXdUPBBSAJt2Vy4sCV8LsHj5bO
QydBB9Y7jVV4Fbn1KcSYpA1qXr9ZP8owi7kdU9paNTdcZ9k0gm7A6UIfmRUmW8zO
4GZ/3c5YZndlJSicxzoCQ2s9QY+F5H+dMc8dPkQyiVP7qvR3sZ80bkX6EJrBCtxH
AahuJelZAI589eTHqFfJ+MPGmn/3wR6rB7hp6RY2nOYBI4DLcHT32cAYxzp9rNt+
aVXiwKzKgY+F6OYwctJM8Q600dIyvuuX+5WFJZs6rZmd2OlQgcHUgxkg9LfSq1vO
w1qiMoL+IHPivKVDrw9GePzDv8/O1QecMRCeRyaM51nn/lfhr1fEJPgcQ7Tq9l5/
qHEkJgr/Vr6V2QSuwVSrG86Ba//2/+RJCV5qOICeVFt4dfAU1vIaxOeuZ6pRiuY6
0QmAqIdPxWiH/KDr+XtPVtAL34nlsYCs3Dnax3GcrKq1XR8XM8/taU++kE9rtqOv
Pv67TTZkPONXdRrF0RmDolsRYqW+BHH6US3rShpKtNtjsAnN7zrgkPfYEGVGP3nQ
6bKcwbHKrElaTkpAsE6YUt7qhH88jpUk+4PGpkpxJz2X3ImNyHsuHJzOnYAS78M9
7cW+W/3qPK1Q3pDEAV55QBWl0difi4pYezKWmlquRNkhF8I5pMWRR/GwHWC1aCCg
LFMcCfMz9ba8eOtIUAutb3+YsU7Dj0sMMKVYZ1t6dIrbj2E+JUaspJCtfou2Yv39
tK7Q0cnV39DPtQdfhDSSrojRVyNCLayDAZro9xphajMe3H259237GGkR4s755n73
JQEQeTQF45Tw8KRQMUKCqgiXTMtNP7jAVwaQTmLk4unAA8LioptWo+XHP8AvSjaW
SfN9B/5rER3WjTYJB7Ibrja8W/amYkdZcIn9kCIBiDGwtobbMBJix/ZJvszPnBrM
NtoH7AOkLB17NGGaT2/n2zWb9tgt752iK+GHFpEGq3TqcCGONKcVstZ/h3/sLbkN
COXWA4+cxCzcALaofWXdq8QWM9A2PHivBi9tIgn0SJRV3LH1s4WyLN5/QvmkcfZb
uPa8OrEpV+2dRRS6LydqsFmt9FCrQ+VRuvcycRLt++1nQ92cH884KrMefHxklx1L
2zq3JViuL6FAO5ZxupSBgVviyzn5ux92U82KC7208APIyrtbLNOzIvM280sm1aem
+1mCH1QqP9gVDedmz0NNyQHfPsAHdTmpA5BnD68Os/5JAaoy35s8p8j6+oLqR9B9
6hKc2DCXKLDkQV5W8T5hEWizpRzD1ZSerTIzIw9lADJ8dv1B7uyRlq4Jw/6Wlccg
rMZ9eA0r7wg+UlNboj5p9Q2OUbeF/ZZksQdt0sj6AET5UgJgZJkajH34ADa6q4oN
cyJLFHPig4RrfK421cGdFP5Ruqm7eBPRS15Jexc1Ar6UXggbOe2YfTAf3NrD408k
DocQ1bS+8oAhAaz8lIqJg78J7OZ/LQ95WsSSew5cP3O9MMesKhJ9OEVQLhCujbri
hgBsl0lgglLOFpSNk3088hgA5QqVtd4vEealMMSzA36UKD5uKewIuJ0YzmUrF5i0
QFu4EBbQD39sAo22oCfkHN0ftW9p1mASsWz/r1tOyhaFDWeNPk2/RpzrrLnvCDOX
SnxUaMNRgWvapz7T8Nhtfngr7C8NiliEdbdr8N5TyFnuxsS9SEANijBgCkS6pU3i
vx9gEY/XjnwinyNltVUaxQgOmqDMYRv6naOonfdZL5nU5dlnjawzgejhdmFrDmsZ
gN9yyg06fuVPx/l/xuzgBGlkuGQ5ZfWysSMrcPI5fyG06wpoScNZBrjZozVgIu4f
7RGt0SeEdQb8XCUvZFilIbelyL2Y/9FIR38BYNMtIOLGsk3tC8XCNXfCY0WgfYXq
Y7mIBCjh5sbaCU/Tr3e5ylwvXI2UYKlS7Yn/XSxd20dFR5tTdz48BmZFd4fsUsaN
s9yNzI6bK1m5/nkn1jsyqKfpVQ77GO2Ux1vzAZXFauLcp32SNujSZyYl9JLxrMQh
sSReYgxuS06v7230BZpnoe3q69R4GOHtV1qRquXUjmdwzsYgMXP4LlMxu9vs7aWz
HqaVzj3Iwvc7cqsqOIMdDh1ylHqa5NR6ARPfCS5Kp0FBkjhbcz8oZLJCdKN7YDog
bLQll8gq5+vhMDf8TSgTwQyf/tMqzfoXZTTWMjLT9txTxnM5r8ljOAto8MLOob5o
0Vfiik05JMXuWCMcr3cFFHgpmXQwVYDn7ghTfJVZj3WHcHs5JKUnX0UEQwmVVjhL
7+CmpqUQtc+UyEgbkDpzS1roa0hFnbLjYm/zv+yELdCXhyBT+rz5IP9H9Dp7bH8F
2XJ8cbOKmnmXgVaFh8D4HkeSAL9FmvTCpTJWkJzLQxE1QevU6Z/f4jH/qUwSotML
qozN2gwJxgdRA/L7N27NkHPB2fQ/GOR2DYIc58XQ3LxXQ3SCEoiX+ujnFF3W6GnW
LJv402r1cI7JkZPwSh6ZIH8lbWq7Dl+wwVJWofFvNdrXhPN9qXPS80LWeAIHwL8L
5w/iBI0WUAFSB1A/Fw4stwWt1S2pXMzmLG2Yzf5yfCX/cArXznnRfm5cMHVJt64o
rQgyjLUzc1YD3STTTt0qGFSVJbvuhuzjvWkTL5ecQ3hO5dzi1MrCQy49e7MDkyVo
OsmiRiVRTm9up46cB4iAOU02ZykE/apAFHwfnXHngYt2w9Aa2WSenLd4idrR0D7J
W+HfgLP7HhydyaFBm1kcO1f8Jz7TWOvjpzSolr4gVPH6cmL1YfNxPKlYfHvNtoBU
8rNkzEnFaK+rT9kpB8xtFyvICwb/7TpEX1lBBncj9tXJhJSLl3rwyPNeS4qR+H7o
GaWCbVV7uEeRC7q89DnO6dwYllJP4Nm7yxs82VRSy0XlTdEPdotEmy/I6yR9Jmdl
pWtAZsn0v/SENRS5pGuH/YjyA2oykinYAkoVQrV3NUvBsazabs6vh1tqkDIFzGem
2DC/ip4+08U0T8IoddZ5n4SpEyoxhWg0XnnnKavhd1peiSccjXVGHJtYKRxWTjz4
XTC9dxr9Gr14WRT5Ef4HZOA//bGTxiHVZcYCTPQSZ0wS26+HHYQdGNtjFkcQRHtj
mCcYhEI95zfridlGT/SK7BO8fqrBLjhcWu6Nn4IEI9z9sPw9iiN58SbMVPMgXMPz
I3n2sxxzIslDOEcwmRofhgs5cxQwxXQhSBZ3FtNV1NmRVVcyXqMlk9lXs3VV+AE6
g1FW2uJ1i4eN5XHif1ZPo058diTtzMQAYRLW5RNsOvdPApYKWJ5+/4ni4HcJ5EkX
SaNr4I5XqM1XvKhcKVzzgloUh6Xf2R7ndvoJ9i0/xU5F9RIi23xKlZFfSj+gmoVM
8BXBfWX2wRJdvtwbsWTEwr/2I2pjLrd+aOWmo5veiHHTKLOFoYL4gH5KOsObQ82S
7XX+q2CKWzYWASJmY+ebV47LXkf6IQLUdRCKc6L9ZQQoLQAnGM0l+UuMZx20LoQp
WcEs3US2Qz12lJ7ZxD31zsJU8+x4PjoIB3i3zWzB21Fnu+X2W+VAqfh1j6xiylmW
o5I31YiU7eXTyewn7PEe3CpqsEFW0pHhUKaVop6OsSpwuBWPMuFgYIlQXHVSeUIV
WY3bBKaDEuWv0EkE2iTcQd5py43aUWRnMbh3/XZUPuBytZAAVLQPaSuT1vARu80X
+/s6kzBid3XXB+1lQp065I2XjFHSXGqPUOVoMNvcAS/ChidMCJBSotE+f0TOqPpc
bpPw3+SAAmsuYznggGXhXTPyh0DnbAoqjgeDsmQtDKHuSQjtlJZjwPZjby3YNDnh
e0hIffxJUO4vcqpy8Tqr0ja9HUTnqZEk6Y11i5d4XMiqvHgGAcUCCTj987cCsVm1
8gku1/eYS+6IMkBjgcW2YccZ+SiClHrGDl+IApmvx3NE+YWFcor2vPjkXPsNIqQq
k6KJjDrjj7+vg9HsQ5YgaoAZFbDdLUXRv1SJN2H8b8ZimbxzmheeFGObDJ+pCuYe
Wrp9yLzcuXRSJ9EWWk5PEE8UviLAeiuU54VrUcK9kU1PHi+PVGMgrGCiA4uUVSbo
5o4YVzCT54yrKQVDi3YJVVQkDvNI602J1IsH5AuOxWqjqfYULqLMsvE6auL97Xiq
ngR5343AAZM4bop76pkMRx3BLEV/ueLYXPA3Zk2XOTEjHtrOjBGTHk7JhrLPUXJG
eQxgoyc0+1dFVg/xeMd9hWHjPrfYCLHx9Rk/jqk7ha4iE6vKr8lFRomU4LMPjut6
UI/H3j+egAkmd3F0RF3C85kFmu/ksOzSHwurgZlkRxCQ17LUyG6z+FrI0fC8CacJ
FpromxYabrFrY2vfhxOX0dPwcpiDhwwFuYqrs/UGg7r7udoWF6IDfU5LiQkwwwoQ
lOP+NcRRXw3K9YWzVoILTJPZKDDu+NOsBEba1yBKwWDyRx29GDXbdtq5141lALel
dQWxWrx5KWHp5dxbTtmpwJAtQ9GJqa/+AfdlkmWZD7yzKnwB0KgqPLZJTD+gLKqM
C7QiqbE2HjJh0wm6lpGQS77GYWzo3YnrQdtJPp5uY0BT81bDglaWDu0MkIwhkaEy
soptmBZa4A6v0/vWeGvfwub58U+sqVwUXorIjO46cz8xKu5KaFfSgb+YVf3ea5BL
cdlsonaMnGwe+smrfD8ZPwxnyJz2U2FPJ/3Z5RAMnDd+UVivQi6pTX+I7oPx6peu
yQtw+1kDr/fv6un7yUUzyVghwwJVNhlZ9X5tAMsQnrn4O3klYzAgco+DY8+R9ggd
EwtacZrO4V8J7z0fIAy7up9xZk1NSiwVDIwlGzOLSvECHOWKJiXzD6VBhlmI/Dkp
mwbcASafne+UqEcfL315HR05rhbTV4s/mkLzwwWkZVIVtSHzE1BcJNTO5jAR245O
XvrFNZpyNS97cn4klxV869LlkTuH8hshmkRHrOXKysuS4UpePFNjz/fKZTYgFt/J
+BkIf6jDDyy/YL68jU6YlMFvtvXOi1pMqELHMf6INjDrcqxQKeNpclSDQDhrTMJC
ulxyEP3m85kC6J2cUQx0kqlYZS9RhQ+qWc5Vlfhj2HXDo2lwQqtulbmP4bWxTctc
Ztj5SMiXeNf6df9UiizGzweA8Hfo9nxKWi+zHxgfIbWI1vXTom6DkScUPdxy7Led
/HM3UJrJ28iMK/A77pqaQs3FHq3eBiPmenHSPl8/qQ8i1ugspkw8hgwJYCFrmNFY
WE41I25WNGUv3a8/uq6CEmTAD+VqdhxlkzYurpTsUsbDcIBYfh2o50CIQFBFiEFz
7QOUL+9OTcb5KndpAGZBd5UNN/M7ym5+X0Qx5KXoxCyCrAVSfpg15OtliwYgdyyY
suuPGNCSyUeToAtdK0oivxHm6O1e0qcHz4Wv6y5wnE57ZoAIUuoAK8mbdKIVX9e2
Mm+AbPUG29IxrZCZpfJk27vI9GNAuyxat0N77G67tHlu9mIT2K7HwgF1t08GV1My
Hdvq/6tv8j9MedtUdBu7bMZcL9rlhvl/aEHhkx86UGBOraXd+XuEvTSsNtNSv7rH
40YqKl3UF9UBLSQnrv0DZm/ldW3slYnbnngFhVTaTTxEIThzSeiHA9o4lr22C+aV
0ejE3QXPqeG7q2kxgONF3EW2t9qUrnb5DSPd9yg7ZSem1su1RudXLwmd6lWgrv9F
vHnlJQpmx3yB6hc4H4yE4hrV7CekMj8UAXCbjidbKtcFS2ilWwMhdjVS9mKG6+aa
O6HA1OjOCxPm+14vV5a0ohrCvDltzTqFxprlHN/1VFIizjKaazIRI1o+P7FDPQUj
qOa3ixAX7eUyQqN07h4p253iHsgyY6XES42PsI98eeBwprKcAZ6FbGe6JTTJXfmR
nJftRN5AL5t2hYSyhzTjeJr5eo9iAu94dJL4MC375fYI6F/86ul5Gdcz2JN6166N
LnGpMeV8gJczhuwpZylMgvXJWggHWK+rmCWWELLi4/fLMmscmVtVo5gJGx0P8TYG
TTyTuNg8ZOWoiyJvlTMUD35ZAqPX+gralHKTLA/tb6h1hzcUPGOwCWO2oTN3GK2J
izT8phqjGA/WLMNjXZes/m8wMC6tYrZpnserjcd99l5L3BQ6kxO52y+llq4etfps
LX6/XfMb28+tlXoTrxCPOoSr0R1fC6O1Oy5ggrgGsLMetiCf7lP0EuczGkh86vgH
d7bxl/EFxh1rXlR8j6eoD6Pc61epTAVq7aby1luBV82/qIOYASCSQLvvz7u2ZW24
koYYTl874v0jOZKgQE/TTbTalc0KRFMNUe2Q5XPgYroqn7kUZBNNlFWKQr/jCU0y
P6htwF7R+s1oSpawZidW2a9dNqHARJ5qIkAcErODDTNgNHV19AwCrjoxY4NhW2qM
nvbqTDmlv8ZwfyVBLdgKXwoVF8tqwKtywppFAQB1QgY4mFxE3cYn3lpeKhn4Jnmw
R0INB5ZzMYXrI9Q/ktzFJcFCwQJ4cmV1Mo5Fi1ZKedSAv1Sb1QEyfu32hvkWKvzO
UUOOcsSHO4azEVIa9s7UUqQWHjtk1TuecbMJ0W/vUs4KfLdI9i2tUbulQTu/2kCk
VuV1tInJBsnsKtqqDurdlUCfwHPyIRi9g/xDPQ8UDGmwDPiwZ/j3NUEuiBD9+Scw
JCKB5qkXlM6uEaBbr+JrYehDhCw339wsvNPxRXprCvkaoOO2tOm+hhZLTxJPoP5m
pQrHzdGIOaKrzx15npLu8M/aS/QaEtf6px+iyhGlLa+EwfVT/FERIVuibB00sRlu
oPhwYj8TVQEGfvpKlDHqT7I0SJwzJslvBNJiXHHxEVmoge0PIOKfzCdAAMalkDh6
dEmxK960/twkGXoupSOHqiVuIf0YqlPOXZgDFhq6Tcd5v24CcgVQWcR9dAH9mIpj
tStUCbNvJhlSb5lZKky7zHCGwCmAcJlosK/zDUYWK8wY1zolPjhXGe73s7KGpTi7
bvrreOm5US+XFS37pUP1gVRA0LeHRMk1zuowtECEd7f3oNGcBcG8HVQHJsmqOvjg
zsMvakQdpF9ATUpYwDH4pOLNfW3gej8oGAYSt7nKE7VnKf86x5VKtF1A/pFnhY9+
UqzLsKiYvwd/uEHT+L/kLTTMG+JDs+MjNrMjj5YkjMQAeUMQ7Edo6NUZRKPAThXi
qCcrHw/havMDnBzW2fTZYfYH1/ZoOSMIp8zX8oMhoqUu2if4z+cKJGXsgqHc7VpO
6Zs8nPJDCSaT+xnuOGJfObClSyyr81onPv422u7eRM3URc7HjwHAVsNYrjDkkuJs
DxW0WE8xbrS6H5uOyXkZCOm6s9SxPGbfH+WzGz1AszkA8angRqc3KVvazqaTfO0E
pAJ96JRD3Ycnc4B0/fPqeABzfAbtcHYDKRHoYIIePVOaiHPQHJi77KV35qdQ8M1T
+QF03Egi+pTk9L2l8VuO+09B/qj/HSjjBmsBzn8hJNa1jHbIXrsypZRf4dLPlaWG
GW6EZZBvDC51nXR4Xm1QIz/hIrKkbe6QAOSmWYSZblP1YfRyZ4piTe56nM0nTK4S
7Mk784znrAspGunY0Lijb2OkCjCCudTKd4xW43eKZRlv/OvIAIqtoasgKH3/jqk1
hKk/3oZYJzP3Tp66OOrMlvdhIcND4p6+nMBVDQawDIT7I6/quTn8G8ewfSwckAsC
Um9E0lWgrMH4uTTW4Zd5JQHcZOUzOWCS0XGldnMn2at5KLFSMFLpLGs93uGhE/JP
7fPNpnfkKIxpxf6uQIe0AbrOoLwSpms4lNJKKK0lYItjst6JRsNQboFfYYzs2BkY
fxYeKf1OYW40z85OLs8rJw72EEnB0mLq2/i4aWLrVpsUpPaYzgn0BDeq34vH0JeE
JA2ydMEHx5v2zxc1GwrQDuIffhUB3AqCmAZpwKk3fOPEBb4kZVggCdFFj/iY6PFN
P95QqhWO+Mu9RFq7HA9kSUDLZcZZXsndyNppcB5isz4q8r+NwSLRKelWbkgtW5VV
BqL2wW4hBHKgqIs9qGGKjQ+StvPlzkNWgq2no2ZmQj/eFXjkY28c9bM0+MuNF2Hu
usWJfboxmZcbnZucQkbv/dNiEEBALXNPApXyb80gMrIcUt+/+UqrLd7amIG7plFQ
TEYbGAOkkBiiIBlFsxT9i8gLEOJpWpOuEgbanok30wb7ZKHn4ayfllrfaQRPpB0E
mH4la2//0bzPDhedrS3Tvj4fIaOjZwgHjZ0cEgROq/ak2CjoKuRVpko+vjn8joAV
VgEOQYQ4PsvJTW7d7pHhf+9GziRyNwuKnaSrwMAnprrx45JNllzQOKxyYmC/Cum/
HtTnd9s7Gqp7aQ4uetF0KvYdqzIYAkgGwxlSigw2OlN8rld4pkdYU/DQy8kKu75p
Gk/IwSc2ZgZC4hQBzNdTvlVrsZ2HiUK/qXR5b23nHKdW7TRoCkkkbGlySUb8tOm8
IXGOHh6yB8mjNZE91n9CVDXR9OhInjNNCumQCl88gKYFcqNwCATWOTp0i7UqK5Ys
nRQ8Xsx7KlhYWKqdHvZjA7D9avvemrlTQ4W3cC4wmDTJkD56kW2wTtSupsx4JhdQ
WfzpeITDEI16hVPfsuvf+FyLEXmvwXCaC2unCV3kfl0qaboPDIw69RfzDsCEtXbA
HIvaxe1LleF//35KJvZd+e95SGYJmRWa6fNFBCJ0Y2HPaszdDqhI57uvuCsMJWfq
p96PEYoL9aaCGSrN3ilyMSFpQAqsAtqC5iTY/1HQ85ppZwpkSqQgflhWR9rlKmsL
9QE2cc8UO5K0K6lum285FqyemUQxI7BiTUYi/Tg7wIuf7px2Lu07wFt/JUKnrdXW
dZET6HXliq75Ty2MOVxnKj2+SRoqiXbj28htK97iV6BzR9RuIM8O8xGVTddjn7wn
x94LQt+AAyJ71h/W7grnGDys8EqsnixuAvusC0N/8vGo5Vvc6BbKFJTOPOYTZcbK
/Mee2CV6EVzRxofbVtJw5t+hy4h3k3Xrdpk914jGhbSeX9PFX36iWqezzjxT3fSP
9agcfRSN2kzCorprsTxPLYdz85G17t8c0QU2omB6sKHdNNbUHZIOmlDW3/GomvEf
RTguMXYQ5HESnQb8cqqahnhwB6RBEist8Q3NX1VoMnFXNJfdkP0/AIxGZU274I4g
2tjftKWVUIBT8Uhgzy19q26aGf635oQOIEB3jaV8xoMi5efNZW1A00fk1MRwuKg9
+5l1IawdpOJFrutNbP/5K4/ohDQk0LoBm+bW64kQDmZO9IXGNbZNDKoOnEVFkx4k
KdBxcGF+MPUieax22me1KrtbyIn614ZBNepRq5Fz1i23fgBKusEAUWhGZtIwKlYn
wMc7BPN777CJJ7tcTEarUcrU94FyP8mEYbrpqeJOHzYEFoa6xLzcbCWFl4VHeV2h
oXxNTb4q9T6LyPzbCJV8RQTu2s0AzEXI80PxMu8jse5xOmXOI7y/VulY7YPxz7/r
dsTt29urFVbz9pLRUySIfz6t1oFPOJ6OzawIZ7FKqLtEIeFpqnKJa7PgRQV0v0u5
gg4HTs1drAd2HZ9fE1S5XLQLUfoMMuIMo0xv/u9IDGUsjrQhaQE38r8nguaHMtfg
1Q7zRTzkuFIfXUt3G0VRONBSEJMpFh4L8X9tfya10s1xsG77trw/vlLfyz15icwW
WniM5hw1PJ0zJRHViyzEYb+altPiVOr1J/Q0MKG8E0PKSMTyY/QQLybiWd4b7hsn
qMjTO0/ggghxZ4+r0P7Shs9m+3VIv7ItaRq+GX91Z1emj+Mi1XRuL6wQ581kK+C8
mPTC6Ieba/Smt8+JIm5x6N7aNsMwc5izTQeUvw+env1HvQJTguCMJu8ALl3cniTr
VH0JtYvtzxOg3ir3oTs5QuJ6WK3r6xleARHXhmt0a7DtMuAfd7mAH359s3N9h6LN
nIM33iv6iLelHph7lVcl9P+fUWU73fQ9rIGxT+5Uzp+jXgI+LDAzkz/ylfB9yxjB
WluH4Lf6+/phBbsEVhson+Bj2FybFwaG1frLPMoDfdshdUwzob2XRBRO8eDfmqpS
tYkcUC3M3MaKNVjeJjRSaMfuyB+LgSbaUIV7IoZrm1qhBnZeD5BhrBl1T6a/846w
mW7u5GrqEtyajiKmbWN6pRFB1YkEYtFiq5t9FRIAX1cfVqGZzBbmU7n2q22L7ykW
8aV4BYcWhlIea9pgCM008S8EanFOq4Rbyf/MlBYC7ToYkCptCZLqgSqw6vfR+Epi
XJ7HuV5ObUkDkwLp8Z/ZWQW+ul3Hi/PkUGnLs0KxoFd+4iZUHn9JGAVxS47NfFKc
GLUORF6lJ8wSvs6bOR2ho+E/qnIIT1V4BCk6wLApa67uJonhpuyVn6cm5fk+jCyb
R7X55eAlveYDT9CucZ159sR+5XmFNXO3cUYd0KqnZMjkBgNv2ff05/sCs9vvsmuq
6u9FM7X8ppTCI2vSw/cP75myvpkJM6+VTIuTXDcJ4gAKYZ6YEzKw1GOTaMKpuzge
C+0k0JPp2LMcwu//x4xtZP+0lU+E4w8wa9P2GycO9ARLp2cevL2qwwZcH/0I2zGe
/AWTPCIIPpnZHhw8wV77EvqX/2+JXPWgniv2xW1gMMOqxEp9N7zStE0ES2ZPt/7X
mcJAjPPEtm+wVe7/3JC2zafOaVkoo2mVSV0nAevonkbhrePCMsO4ZRDThkghmFnh
YgajQFrkThJFWQZkuNR29fxDcufkz8b8gHY1v9BxKYKNPz3VRj5+9j/lPU884rK0
RxPa5I6n/cxLkCTPELlqJktokJc3uQc6NES2YdPd2hpQo1Y86y3qVy7y8nifzRri
PfcuKHTiQJQfl8BiqN+cPZZTRwVV0BVh5AFdoGSABtmmU6gZrGuERC24i/4dWCOW
ch//J5U4uSGd6nqm4uhtBS/9RpHA0faD6xd9V3e6G/DStAtY6RscA0Em5CX+y168
/mlk03Q920Ed5DuUPse6xqa96NfZvnYpdk8p5Gh0yOVZYfn6EIT+HR3H5AvLslFh
RqoCaItHjKjXT2QqRQuHU6HcqZujpegS05rWMCniF5lCgz08Uh0WjGem4KJ9zwjM
jkw+ooSMAkiYHHrFuMMn2M/gfCcbSySqyebrxsV+OdsNByJiAtXyZj/3E+jGOsQS
0DIapkzCOWhbJyZAbxUZMrrE0RHjCWKfZUphzLG1d/cRPt9c3whziyjLyNHaQ+1P
Q9LU28FFi0f5Wlrrw8F1iHDQ2Kt1VQ2mL77t5U8xJMMQ8qq3WOv0qhH//Wjjsdnm
YdEUEhrZkPynDkkFd5bY2CDfT22D+oQBkO2iL3IvoPvEFlupJZA5ZxDySTKEDe+w
S+g0ODLkLRwHRRG5BMlWsZmzqRnsTbbW+eaPhVG0eENFEbM2p0GZJwkoi9TW+0kA
Nzie2Bp/bBn3EwalREhJVYgJTjE1Q81s2m60o5snaioeY7MyTFoFHiy17A5z4/eI
qeuBTfg8V4xDgF+uz6n1XcOVcO2EfT3Kml16R6ysyM0ORdAlRGTekSVyJl9t7GJj
l6OQ99hXAYxjkWwV7+c+fwqRq2TRuAsRTBZSfMS0MfiT2VayaodxiBByjAuvEjg9
Z3g3tRx2D1fxdO5youVc+Cdfud2SoRkwJImpobvqneh6Nbm68pZxipGgbl6gK/LJ
x9TaKAeBlzLnzoglQBkBSfwlzElBkls/6BAjHqY5rb3i4U94PEjwL2BWUxEL+FfS
PN8RggTr310kAUlWtDljeI3R6og1duSLzYooXyzhNhOiC25s54L10GPBQFKDugu9
TgtBr6t/X5NwUoM7K8YRaf8ZrolsnPW2U83g/lU+/bPUknYcA6Sl2D/nSQSfpZxV
sGsC58u3s6MxcnEselkcuXGWJIUNaAgurLMlJ2zzAAyyBTTuTHFUInJyo/InnxKh
AchkUO2Od+2JtgXAS7YijTE+WD4XNXX4jWhOXzyqKjsuMgOqp956syK8OEH0ams9
j9l4W8aOX5oVQDu7c3n5Kf93q54awJdni1o2iQLs+5ZRGlFHIq3ArHm7TKuKqsy/
Qp8r2XjVEObjWTkb3DcWsjbDtQD/XU/t/ktXsYWmytv42JqXEkzQVuNX0W0Wyflt
zcQOdT38d1BaFlZ2cKgoP8AgZnZkkFK/MtgBseycYHCyCxDGEziHp+oRDXyTKoTU
A/9RgXr5D35/8XiIqXBX8lWklXlebpf6hCmcqpi5o3fYeGIizYl5POoOTpena1GS
P1hDcTumkT02E5A2WQv9iV0JBKvIX9VjEaHghO7mIv+GBgC8uQHsxh///unH0L3p
NtxlmfTTeiCBAB4ioa1FB4X988JixmDz1UXKuns/RShS81no72rDlvI0fONIrVg/
/TctRunh/Z4G+x8VJJcdHimUu1+wwluyZ0NfBFFVC4S92BEKYUaoe/YwUG0MgRDv
ydaXbL0JaSjjsRC41B5KOIGUnb4h+ldKITixbBKwni3nxhII6XBTniaEx9DlPkSu
Ynkqz3CiYVbV23YWS1v5NoJWbtZryPOMwhbOCKgu5Fu+nwIgseAV758Jd2T7a1Kf
tDrJIfnpV9RcWzthVikGzX2rtZwBhBwvi71oJpqIed2eIVQtYY6OCRB76PUn9h4E
PPEXTqX8aXSKGcFztVV9B+3SclClFrcJYUljgGRzTgJtW2ctTqiabtiws5chiDDv
JxeET/s56hJxCuNMlfOoGptC2EdSGT5a2i51JaFaMxxfwh8kcRTHLPgdbgE2mOQf
iYWjYpRSOvPQwILWEztOyPtbo/PQdAeAs9hhKC2kYuc34A4zHcdN42LAd7Ymktbv
AMu4CtUl5R4epauwD60vOBh2m4R36tOS5LezcA0MzGC+gJjsDPx6UBzzETsm6rtf
dQpFS6GD+i7N7lB14kAxVpon3GwBIGK+8yffhJSYWQJczZs+XlRf7TGPOmgxJEMo
zq2Kn8walfYmDfhJ/3t5JFG0cXMNFGmi7/UY+uqvtw+dO5ht7j99QjRuWVp9Hoz6
6Ai4p19DKGru4cH8mDI2Ztfq5hakfvx+PT+zXwHwglADa41lASDeQtD8YrWxjgYk
TFEwF1yuspVCCAIg4A+ItfarEFC1mZe4mJbuASvQK1hZkjmmjgn2Rfc9Ar++tu7z
MuPzvBpnliCZvydqsnG3yHHWd5z2WXi4InWv+Z91jmXT6O4ig8PvogQhFufdPTa3
EKDDrYz9SSz7sjDJtUhq9kS8Q1XFbZo9SOdAyxuTPwTQSexxB0Yd68oWc5QCZ0O6
upwLURHmv94l6VY0022KJeciNJPOG8BSB0FvArebNtvf9b5UOhDgBg6Mx3AzWIxL
GPFThCJ6UMKFoiC0i754kUoG6iaTK7Kjo/oOEbyHioKfDSbvyNIvhxlWdFfDyjIi
ebgFO4Zp3ri4Yr6LruB/heyD1StVOeHotnQZeUTOIyLd2giRAjBllxCCipl0QS3a
Y899fvwqvJOJd3+TVpUQ2zTRn30GU7Wz3lBVRk0EHEI8O7V+JIGBpFV6tj1hGDfX
PSnKy0l+vGr+mDVEi96AHzgDFK06/bL5XrMZl1oQFiM/k6Ygc+lPp6cklXCgEmdw
xAQ0J0gtuzwEne75DKrYmBacnu+ABe2pmrriJcSuJQLIq+38Ut8DBoltQiAs8JRi
5/z8v+xYKjAn/tvq2DDJJQVOqwRSxxPplX2ljgo2RxknciU0IQVsKnVkpU6AZy8a
nlQlnc8b6WcSdbz/0koO4gWJGWD2GyVsV8mnOnx/0pNFXY/2ppysdEH8OBCQr9Ts
VhQl1rp7+qtGLC9hTVtFJgC8Uthd44JD3B9eqzzMW2KsOU33Dtc5TvxsauCH+IxZ
wXP0ucCOdFMKe/qUYuQlGBS4jM5FsP1q6xGOxzt4lQc6/wDWUEXMl+mTiMJg5l2r
n4sXv/9FGA5iP19cExqnwFN9p9OrWmi0pQTH460Btu9BZaVeuQbumnjw2TCK7DII
cJ4ascNltPV+RQYIpxWhuVIpd8QEp6mPEtrtMVbBZa6eOGjJuI72xCb1Gs4EDXJB
T8MpHXRVHcDE9RKjWomFg61l7QvSeJu3e6QmZJ4HKYHVqshmZ8F6+v8sYg3nOkVl
IkTqVrcSKoFFmWKQ6+ZMyK6ObJW0B0QvMzWOtG+K+SJ4hRaC6rP9B/crgb0jsESL
UX3UvB3o3+BnZZHrv+pCPJrO93H4CxrPOUx0wAuHUDNtjQ7da16JF27NrczoqhVu
yxEEV/u0vag4+kfYJxMF74tIkpjdN1Sl54suSwVn0kc1reVfaVQ0kBtVPdTZ0OH5
dzwYufd9GKKrj2CgqVYvyYysPWQ9ljyFbD3SYmaDZJEj2dJWgTayt7dcCffFSuV6
gD4acAgC1FA5y66QUd6K21OFYWEPCH8MBjJJNGjj9Wud2zGxbG8jktKRLyzzulra
BeQb7vh/VAgbhWu72yEtPuiNfqbCv5msf9aG/2YYMv40nCCRh+bcy5pG6XwsR01F
OGGgbskdbW4Z+evWqRtKi5olhrfvqZF108/LWvFvWAD9iRHO9nBZrtIg9D2RaJ/G
TI+4MOOFCXR5OAQnsijYm8z+zS7siuXzOa1G61fnpaKX/HpZpsykuI2caHRworOx
v55z+/SQtMqe9tDjV5HXMsQ5VPNVFJSudSN7Xy2PBHItf6RYwuuWhvPUn/4EWH85
s3IUC5fhiSg6twzE/wmLZPxFe8W3LaVvssM75Ok6yYed9RZRQbV+MyL94YqUW1Ps
u7fC4fD2g4unCpL9ck0Flzmhoy/UjR2Gm+M3Tz4iyJazRJLR26/oYwiPbozQ00F3
iv5h58zG6m6FGbkJeY41uSqXZiKG81BOus6DHdizfwVw/M3UXhjXpF//6IQyXJqH
WXtApIkFLyVKd8XexPxW6heVCpWADu8H58gmgceGBLufjX3yQ9U3WcfmYWepYHjX
tXDorYtq3QNwYX4y9YKo/zZ6CmkBGu9/ONhnaVyKE9zyj+MwRsIRRDrVCD0ngww+
a4bP7pPCn7J+KrJwbjuL0mQTSkvbBol0mPUr7HYDSgVPpPiHGIua0NlR4n+KdE7m
U8+RDTB4QWO5JsZmQMIYiW6DdzwPLZgi3ZY9eRQLdEe35DqcvFSTMs7NiGDKJmYN
ztSEUo4usRuBw7QUnPfSPuW2Ym323ySZUPhTXwLzqjZlQMN6wYoFGlZmVK41vl+F
l3y5bODA1FVg2/6s97XwCIfJz23HQKbEeQmoB42gtXzOwV2kFxIcQcBhf99DlW2x
RlTFw46+hVKDrHBn1u1JfFr0AiUSI1rk71Tb2kEBBgXD6/cq1vCR7nl1HjW19Ae2
ospoDVX/luPAzfK8svOBOKWkCc9+IVXNOxlGd6EYbIijits1bOeeczIaKGaRWkEH
04Ct4cTOkRe/OPpve3xuHJWzHKfpUQAaFBaFp9sKJIJ60b1CZ59hBub2WoKk70Gl
8EENEkHqIvBilr+39crSjbB/azmSEMbxJK07aAcRpJTvcR3LZV/5bGVnNQwzk7F9
SLLi4L7iUxLsjHPG+m496iowhYHqpkA6zwJJgJII3EY6t8y4vjaWgNs7OPR16ccb
9Lam9uBVNaalNoM04xB8ro5d7c+nQtI3SynW7Is2kF0obihpebdw8BOPpfSlEieA
b8j8IDYFXUQxW7kgW0MhKNeJ/VPAYU5oSGHMcoRdV3YiBvZGDVU8dJ2vmkHmPPHD
gwTsSFaYmiD3wOgho8fsNKYFcUiiagj2sBen+5G14q3eLFnVipgLgiAsuhdkf4ph
paGqe5i8dLqoeQNiSZsKsWtvjQennv6tFYZR5heWDLworw06DlzzpuXPWgFQw9Ob
P+R8I/TMEEYK7Y48DS7Qb14A85br1ZvwVJxoE7qJw3pb46Te5Ydwz9D2wY3pn0bs
QVShVejV4xWhMM4nL1CQ32imewvNAa2HCs72dbHUEyVYHclUxui8sAON5dx0e+Lt
vKWjERhh2IiYdlqBjvL71MAZ199R9Nc60PDmI2XC77qlmtz2H7w0OL3SdSZBOv/r
CA612oLXgylKciAhG7AcP4ga8aHF50zkUn+Z8XpAYfJGIVeCXkl98ZwXQcKl/H2x
CYqyxrvWsWevG8APhgItde6692gWXCOR0nl6zg6fNQb8fbtHPzATTEkw08nLIcCd
z0RNB2MTGKASmINMxP4uWoPsI+HTuNDQn+5LWrTCZRoTTvT77CjYaHWNwyl4Be6b
qN1unafWIpdxY1Zi7oze+sANnXooA8xdesKYIghs7twzuVeRFToiVkyxy+jvWdrE
SF94xhKc4rI/UvNNv3sy9SX/z4De3OTMJvvo2ZrbOCjuXH32l33hpt6KEKU+3Bbl
bSoDGEoERaZ82h+L2WlIovrlwtEKuWut/X0ou7rznH8vGyRxpIR6HF5V+AsumtIY
rgurasSFhYA0FsCzkWMAyeYPzi0Rumfr/z3GQtLilupXb4FtNEGny4GgtwxGa0Bd
AgWm9iLpSH89ci30Lu4JfYfVdF4OtDh7Xuc0j0X/gDJFBtyFhRJS1yY+8YOplJfO
33Wz6ZzsC2WOWABtx9hIKq6R+4wlXgUMC31BjfjD8nnkqB/dRcpR94yPKx4V5Str
3lBDzcmtrlONWbYu1IvdXvJL9nZMI1M22kchqI2b8UIYsNmrmTpu8rm/hp3gNts7
NfZU+Q/msp+qh5FgopFs3ZGxozm6uzuS0pk8vGr17zm20BducPnPvvbKxaPQe2rx
ITgv+e1aDNyVx+pfBTxb0SzIq8W6CNMg2vFurDMo4YhUMhroQytAjXDLWC5Lc0In
V2sl8Tls+zDCWwiyyWGC2jw3eexMnCNXvlT2U7J8LLXDtomVVSKCfrEVfB2lo/ib
rvLl1PNYI80UnzXGbPGHhAnoI178RxtU3Moix1XpBoPxLjLmduGgYNfbVKMyD0gj
E6gkRMFVOKOthazp51OVW9CUfWIBuhafE1rVb0vw7AkwQ3Ie//2wb4qxdKONbxTv
pca2+MrcMoEoLicUxHXtQMLE/QYGECYkm40YM1OCuyZWQmn+/4Uasg9626WtkSAL
wOuPoE4pfMoolbb6I7DCvAKjjsqaMflz7rs08i0+LU+oBpkkGEpzHSaJD58jr6tF
Ob0e2OcMorN1t3lD0ar1g8e3E+qV27b/oL20jPvB8EoVmxlE1SHsblfGyt8xwsBS
hOLZh8sbhyxcvdqlxsuHqk5LBRfp2jnFNtvQ2Sc+NitskAy/oEI+I1zPpGCsRfAu
P16UGiRsq+xUK1l/4ysmp7C/qYb/PcYFiAXJkjyJkRF19PCtdEVUdStBHLy6ZoLq
98M1/EejJ3z3TngRuurIHAxQM072iBFrs1ONut5HaAvybbzdB9WwBOjMmOcsoBhF
c7BdM6epsIScvuWQB2bteIfN/tXraye4MT8wx/WX0hLvsEy5udaAIlFVNp+tWBI+
oi1OR5Dnf/mljKKCDe2nwyAuiuAoSrzk7BzMW6ynQNsKguQ9DGok5pNlg2Zl2y5R
nNAQHuHs6V2DaT5NZ9AqZctC5sINr/uCeDIcbbggSTzQ3gjfVcQrZ00lHZqX945n
2dH6t+CLvRY66x4VIWu9lKWT2eheaY0I9C5nLHDTITcQ/Wjqw44kifdaayXVpIJn
uHppiCCGX23jStmOWrW5ho0BuZbPZ2jjQP6V3HaVozfZZJcDRngwPwJ/nHD+weMv
mML+KXQ+oJsNEHZ2K05xbvCcK79qwNY/4TyP3HMUzs8TPQ9F/1yTPs4Zjg5tAG7L
p6Zb9iWX1pfsZeIH5ylFFv4zAdaOqo7KXpCHjz6oeK+ug40/ApTh7b5wh8uIk6s7
ZTfKxOu7EhnEyebF3kv5uvUVPvUAa2zF71Rgo+Vd2YxtnMfVZ/kijPcskVBI3R7G
2o/Lb0Lg2MlVSmwZJhrdbrYHP1TbPwMJJnDiIowwEXShRo7P0ocI47iCenUY6l5t
JtswD37Q/aT9W41R3s3nSR861aQzcbIc0ajCMAJLjI5j6YF5mTYXnav5eZry3ORz
YWczlFDELwOkZz1DWQDjhN/2IoInri9bwvpHpoSYcSclY8BjMe1dqvPJjk2OT12R
yTdr+3oQ91Sm+Ol61KkETZB2tnaZsJk7HDSmBL8jhrJOGwp0vNaj2yDs2zsfpu5m
ivoM9B0pUDnbFSX/NNoRSoH3tNhlPeNQMAegCEojE45OuG5UgYO6x+6MU3mPor38
xc0E89VYLitiWrpECGtk50oUMbHStpiYvQZsautr7NHwu9YInkyuT7OVheIhtB7i
ixMbQVnJODtKLMxtFMc6DqUTNvwL1vip8WRhrrtSAGg+7qw/lcnS1c6gz4jKuw8b
QMwnsf78g4WUqm2jcPhCbcmGEVNtvJWT5RbzVtxcDh+VfTlAD+LMD6pYTWtlZ8ga
5TBOJMm5Zxi1Nmn2c8aPidgZVSJ0Yv58j6WCEIvJscy7vqRIZXRMAxF9/69DVfXY
AMOywMD52bXxmFHgoLis9bi7VHcRbmETysH3lBVecK5khfjXVIBFzjX9wfqQLcO9
yFc0947PA7Zvy8ZSEVcOzPf2OGzuCj/tDpbUPaocX7DkTcCVPrKgQhKZrzAXcs0p
4bi2l+MHHiG8qGn28/a67Cb0Ex4DLR7sbEk5fY5UQ93KOsj04e2F3NGOB+pRpojd
eB0kLhGyjBDsfdEFDbdKfLd+0rYvGgcTy03Nl5j5dWlTA929oLQiq2UiUr+KAcFh
UPmu2Mm61YdwiHY7GtK422yen1XzSk3GsaS5jUUiPXJ2lId6ulLvpHKzs/z0fUzt
aS41p6JdUI4jJS/HH1cowtiHnVQ5YyC3NhqFlq+nhCeCd7YN6FqgvQVIcRSbvoT2
uQmLZfnOnDoEBgHf/zsUWYyaRYqc2LOXti2NJ9p75KIQ4sLOUeCD9RBDd0KS7gUw
oNbYyFS89qgu7PZSxAkpwmFccIAcg5WlwtrIPTdmU+h8teSL1MLncX9NltOZFSkJ
SZL9454agarohJfIEspEKmN1qTfSjg3e3odNrMDhg+zfOz/lYJFF9KgzNRbJCFbw
mTG47kkAL+r3me7yra/j4S/t0gA2EcWYjsFlnI6ptdRKxE9sUpptBwFf5J+A64ZP
XPvkIyqo3eqLus33IbDNPePiIOCIeU0WxaQU5t8u5rWLYaqtK4xOpc7vImC6NmmN
uMskvFAY16/+OHN72sHpo5ddk8V88a9My2fbdYOY1MKcOZs1l/5rUOTBQs4uFYGI
0tMZlc2qJAYL5LJQ5iWUtv/ljA5B9DX9jBEH+UlvEMBqTQg/iNWNPE/x6BQwfnXO
0Co/z8uElnk/jzFrdUp5/VMiYIFtmbvmd6seYDBXneoBdR/b9Z4Hlo3htiopl/IA
D8ENnGSFyHYmao3U2ST1H0WxvJonj5F5NJqwHkgtxZfNI0Orrp2R+bnN2QivRfTB
474Ly+cqvcgrQS7Qj5xtiOcxrqWOq1ocC/jsdPMFVuRw+M88YxwYnknP5hNiE8z4
CPf9esSh9ncq7B7cQuvcrtDxmcSgUjR95zlSEHVC+sV0a2Wj56Q0BQVzYiK7m1Tm
odMyxEzTkyrbtvYsSdfv/VxOv5Vw/C27zS6fRDPQ+0iZbPQPpUV9yRMAUu1+EXGo
iIkQrR85a0Y8snq1c4INO+mhnPSx4oBWjXEkTEnYHPvdrFISRaqWK58HGSBY84mJ
VAjYgSGI8U23DhtIRUmtdIVK0+TvCZouXU+ny6MpeuV8J0K6dcgu5f1i/LyUExZ+
+2my/Cbj3ujYVT3+hqGonCGiSSLh4CRxofwKaKFqM2vgXWDsRsGnMYO/noZZfWsS
2z80ZBfm6T1LV3U1ApVRtJF+PfwpZm0/wKz9NSKhX6WgX4v1h1FMdxqwLEBorpIp
tPnbVDPQN3PrZ1TKk9+OJTpTVBTpQ9F9ZbUtGO26H8yq5uHE9uWyp/E+MryAq7kT
9JM+zgLDpBGRQ/Nr1fOdBpC13qPXmGEivMQE2XAxlUznSI2WidY539WPd5FYqsum
7NGpmUobky12vJQ+Q6yT7BAkkMjop208dHevkfxibu8iqyLEdPHLkPd2lUM3/RI5
HfQofXxQRtRvxPzhoFfjjtpsmj9lHDDl7PFW5m8NNe++i1lnoJ7c5yrtqNvbt0uc
nt4nkkoe1/1g4uIpt9XZzWHI76tDOp508OGzmwZt6getmoA/cK56W4vIJK5cjwnS
7DlmCMsh4bxx1IpAfaD75Fm+QnASEKSjBWggewZ7FBLmKIfb0uNq9Ddr8rYF2QXC
efev/035TVHB1yFO/NRXSiGAVAB3wZwKB/ZlTlWvEevcE0ugaqy10yNrCIuCrc5P
OCtpr38cnsHEivFH0kg3K/wP5l5Q4x0EroyURNbdPHnHRxXMGLJ72hV/PHfbgfgq
UyDvZUamhru1bPFteCObM+AAZYfLHlHWEAxqhgynYyupadhfI7JI6gSIpHDL6SrH
ty21nLOeXS0hxrBcIxHfxAZIBMbDAqT8402leg373XQZ2LvxI240GZ74xDSLASVV
elqgfbP9NNMwe4eDKJ7OI9H8vXZzHnJ2eiBnqYlf3Gds6J8ruVjQ6g70kw7K8C8K
zzrwm4Tc8LiE/gu4xTUHFcjs0dWCnE47Z2WsaHrZmSqY0cWDoo8oHnuB+dgT77YH
cKeGJxC2xbnaVqHpm7AaeFQcN8+69H8vy5K9RIsXL6ScbsxhZymxH2OsEIfhpYr3
JmXibTw/85TZkryf7KwT7C+tBjEhxUQ4gGxR6wYfH0l+VOZOXtypcFhOjAR+lOdx
uTKg0iJMg3P5um+H/t0wqftREYn06BxQMW06qoeqxzx/KV6slA+VnKrmwJnU/1sn
ZiAVw6RAiBGK5kTAVxcRLQuqBAc70fr+XgHzYJlYsaz829kirlsPG/9bzq2ErJpp
IcgaZwr7eCu38Gz30bGxd4E1v7hXvviBMG6Bypv9FAG8Wda4t/vCeJGvVzJOXWor
aa3chDLkMoBNp5GxyVmb0/xplrpIdyC6llG2pnohm8/4Cqlk+2/IHyFQGq8z5OJT
DmCNecu1QrOdinl3SS2GlObd6qWnH+BNAATughkqp1N53QGZ3Mg0q5lZ5zJO2IAf
OzufDEBH3fo5ydGN23YT7Fpl+QpwynWwCZiQNyue47fY1wuXzwU7KuedqpCyGv1i
3bn7yF6mYzqNDW2Z2qnXxgUbnDal0+F3bC+XG7gFItCg6eht5agschVum9dqxISk
lGFv4Uzk8qBUChL82DCdlsY9FG2CQweKK42smmed+gE3StdLIZMXmLu8M7HxUjGf
tqRDsDT6oZcEzVL00/z/8GNG/fb5Bofd4C4oMQL4ixPA7hg1NZEFgBA0Jlxg9g6N
kJcZy+Tl+0u3Lj/T/j4dEDlfnc8Gai4MInEQdnZtJZh3v7JGlmWrR9w+zhwX9Fmb
94iWPUGKi4hfxbhMSp9pq1pEOf8ygAvIqUjMRA1k120JhMzaO+bpXWFbMydZpzcV
d3yzE/ScYwqjGGGHKOBMN0m5a6l4oMReOcGpyGHgPbwK/Xmfe8vPttL1BvnxcSg6
a0nMDPXw6C3RZt7hMsTob1lxiKnmOEMugAc7WRBkJD4RR8OE36eKcdx30ho5YSj1
rrFOl+KTanBBmc2UUNFqsz6dIsjK+aMezfxgiL/tT/v/KHGj6pAd7Gt0BHbZZ7FB
brc36gXIHBSp9Olz4hkgL/4KPu5Gpq/deqIpWgSyRr/YChqTYDGHlEinzlL2ESlK
cgb+jwALQ5Ij3sbK3wdbuZnCAVG5SL+e158hbIpdHGajsMtainOpum0mgflMVneO
gmEt8Kgx6vtzVJDfWLX/UiP5Qki1mk8avxwX/t+/eUgkd+xSmYF21Ax4AD7Jhgzl
xeOb2zqAKbYqvUT1YhX6TPrBhQpEc30gkprMBAt5e6CgXXGhFdNIjZlRcUq6Ehd1
4EjAKCwD9OyhLMSX/uJ8XlCK7+mj3VJVU45Wm2CFwzc3JIgdVqcKdmwjZfR/l+Nk
AYU6++cx7LlpkTkuWME16wIPNU4awZbbUO99QSQHY8pKYgJtWp5OJZJcT4qZ/mdk
oEVn8nXXSIDZqcOIFARMUElma1Vw5FLWJrWx5QAwOUFlI1UDin1pDL59/XxEnn1A
YVbMIimHscCAE7WwkUPrEZnxLkXuBAy2Xd3bQj8BIhZo9jLg72da7ilVpU105LOn
9xTDmFWZ4NU6X++J9P4pcWSlyEJCwkY5Kc8LCEiQeHAJ+cNkg8AzC55pPAHnMULk
0IIhj1SyCrUBrhm6d2tAjA0uDOwx9sRD89zMv/2U5yni/5ZvIXYzm2qJXWqmqaOE
sdvxD61Z6uSeKWKd7/h8MQljvOYtA8h5NYyhBP6hqih4hYWRpQWjq/UvNuQbMni+
HIF23QhxtoOH/NCjwFVz2SAYDKkY00wm55Veo1K3YmFMVt0sNbn3QSTNVwqHBiIV
wvtk12Y9YdaTjadw4InkTvFlBMlw/7QBINCONc/0deQTVAFhOnSySA++AQj2xeEp
N7uMfaYXZ/4ve8hFg8LDxvxi46fU8uTYRd+KBnQe7C+I0T7eVd0TqXp8gU9p84vq
WwUuylVkCevTJwbljw6C0w6IrdIhM0UA5rtxaj/B4H2di7kwPkNLpQqaDY5xOfMq
PweRmzGYGYnSb752objq8nhSMMqqCwWpLyCqRFNm86ZR+Sq64gZFl/wXaD0Uq3K8
Zh7XNhqLI3pXN5WjXkl/eDDeTgUCHlgUFlghPF7ayHByZIGc+rIdR6GY1wuJXJvo
2/nXPbLt2VIUsaJaGHz2JdhIw1xjjiz6hz4GX6mkKvwNrRfI62npgedsmD39QCwS
gg0kOBHYNrJTUMFCH6nnkmRWCSAinI+ZKEK7A6VsCRjeAQD1iyAZS8oKQ+nw/3UO
DmOi3AxSRVrYE10jJT2nv+9kFFTnJCan9y9R1DfYh3ndvqNt35dabvjWhejdh+V8
4IvaohN/0JFkVonlw+3diU9aeRai5K8v/cPMws+XmLE4vySyw1U1Kigp4vrgbHVN
QESXrlaFk/Tw5wcghQHnZCEZs8h5q/DILIzvDFFcr7c3yg6UKvL7k958FyUV9y6J
y5wl9ya1qP1vDRI/irqf7BYZuoq+jbZLD5WgUEMOG2QDTmzMYKrrbQl6rGLZq8H4
53sl/GdWJwtRXosl/vyNw7aViTF3EV8YGxO+pB+3P9CK6Lv7ELUf5OjYW0v19cBm
PmPcyzXlvux/A65hvRcJ1ognRHTHgOJpokir5hf5NtybjbVZTupovJkjjEAXsdNt
KGuEu4PMGM+wbUBXVG/h+Z+VjR9Zn61SqZfdv7SS0m6QoMJQD0s3r6cV/bhLP0/w
QyaEYlXuOygl6ycEeuJmau0OjQCXz3Q782/uy9YrAKYLGAYW5jAL8M8YG1VteBz/
SYiso67ppuVh3i8sl5C+27huAkW1noZ1Q7OOJ0nzKdUSLsOpBWRwRNrfS4YLNQFx
h/vSEh8s68axJS3QtorQ4AI3UAoSw8KUuPDUUyYecl9XBnkbNMlOz6YRGxo+oWQT
Zxv0V7/NCunnsTAjNk6UPggu+AmX9lfoAIzG/mOKa+TogrUW15mXWCRy/oVHI8lo
lsDIP6YGeLMjYszTioXoAWNIqt8arBphy80uptu3zho6eImLqL3y7A7Ms2b2CNIr
`protect end_protected