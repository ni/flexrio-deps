`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10128 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRvp3o8+RItkxKTewZIo7szZvdGo/iNhFVQmsqdn5BB31
cLW9sNftAlHSmSNstmtMZziDkGpEWj/qbYc+f9wig4uq9EXrBfNEyUvvMTUgJmlu
wq0dHooBeVzee+K/lnMtmvNJRU3O75miwXyRtJpvji7+wjy9MOpHSJiATyw+Uyy+
fvdx/fQ382uqT4uwFMNksJ8R+8CdjYkfbcBivo/eALRWAXp0xWuaF7OJS3uaOgjv
Ozjkmgp4O83XxuRZ66lgINh1fi8UMpiBkPSlDer5P4LoZE2UVKo3z25InU8Rclq9
9A1whhdhi0cBraRnnaG6bXIGfIAr5+DXhk++rIRAVxcrFQzaeJG2Et0U2SE9M8Ku
kfFEx63+mSJ64H09Xs+ZJKIdJYfpzyIcSPz0p2eg+5xJd2mUk+xNvXuzO6akeZ6h
S0Qq8VFgRT6gpuA5NQnMPUAUIGx0VXFP2kE6uxMj2rZyeHXzbWbWf6OhVQ/K9m9Y
KmbUAfslmwi+uULBp2ZRZDT0rq0CoetubIrIBy90VMnlWnwnZefo21laStIdczXJ
FqrMGsP2koiQHv9INxIzNZxk+1ImoVgdc7lncb0LxlDtM6HYL/UUqVzOOINwdle2
7ssuZ48s/HIl6ZJbvwttPWBJYY2k7JtAgjas+nTvDfBMim+c2G0mbW9hPPmbNUq2
tUHJRRXgHp7GnOm7I2hu2h9WndRQDlLcXNSJVcKsLM67e1LuFDf8soL1eHy8alnW
MjWjAbZ5Ve/0aS+lBnWoDrF68Q/i1RfKCAeo0FDx+j+vr+rP50rsBgoYYc6K7qiI
CJ0k2WlgIsyxwVlfpp6+jWL8HtiXD5BHQWC35ffGmTjmjYPCBQOxFaVzLFmNii96
hqu52jEyHILc/5zbc6n2ls107pGdtpNTyC2clBKDSbaoFgd4Lb9g9Gj8G2C2Fd5Y
KqbYIbrXorTSWq7rl0ZZTim/vMJPgMTEu57etXZND0h/VfnxvL/9ifpZm3hs5ipE
6uIupx72vrOistARKqSzRAbu71Dxhn2XTAPAEgQSrHrS2f8FJRu5xDXteYPJwlz/
WXC/Df765gxJ2bO+XY0oCxeS4Oi+iCbvMW/znKP2si4FKHp1ZtlNYRxuPMClBJC7
DAQRWJ+i9gah7R7aP+uI9ihHMwnDOKrgRR3jHej7DEoV1ZaeQgRUa5IbO4pggs/l
dgeXYWz9E6lk3re6Z2WecpCpr1KXqFxXds3FxGRVgr47gH0QUj2Qswu/SPRszK+z
7fx96fM2dmUBfN8N1LdCbrPE03DY8V7lJ+6FFbcpYh+gsyuM49ff/2WzKmpy5pO8
B2qJ3bfYvQyxWiYw/dExnXxJatzMsUBUKCvJorFVsKQ3hy8OlfTFDRnH/1clVmil
JOhLyGEsgfm20mJR8FVWR35IHzVoxuX/34FewpZehdmYNRHt7vpIHx6YXm2wDpDC
WvrV09sblAW9iDEffYucN1yMVTIYugiHTAWU6giXf9qz+6Sm7kXLq03M/HOusm5h
xr9rJuOeoGIW3U473JI4yoKSQ38aCPGj/cly0vrsQzt2U1MYQF0cwmLgwJjKZSbT
n1hH3VzslqzkWzy3Yujr36sp64/mTL0yRiNnMdfb1ZWkorvz2MMaaSH68dl891Ah
aDJv3+/Q0azoR1KFKd0pN2ANhFKfQh4dZLw+I/wubA2DHaGifLr10tnoP2tWXDkw
qVMiXDyUE4NAqayyz77VaVUs15K4+Tb3ZnXJE6eFClNF5kzumVWvgya35fV2ZJrP
rcD8TWM1N9tTARWBUVKLY7ejFKDDOsDTCpp3MWLPsa738XNkeqPSe4xu+SFhjLGg
NqCqzZmMoEIobnMh3U9o7FP5g/9MdmJNDKxF2HNk5ha93kBIAUnKRdX0VH8qDJLa
wUmhc1uSsI3n7JILaRrFcP3aE8xmNu9gQae2QCHOTn0Kue2QTubYbZFFVbtqBvP3
yDdb7YsaHUNj4QZbBN3GmxC6BH/qeYueZsQXmyoU5GXg+bXCnpjywSx8Mf/Dixrd
BF+A7uNKUjBu5rQ2sUXQRdY5AK6WKHE+AzMhEmoTvghYU9sEqOPj1UTNbTTbTVGJ
WA54DiDF6yYoGIGSmxWlfapJv4klHPaEEJo2yJcgJCpPycpxBIFS6vBx3+0iO4E8
3ZODQ/eYFYfwa3g288fTIfwODphNtKT3FJTgpSUv+M8T6ifw4YegwbYGsoEr5dvH
SK7+fHmlxivSOrAIbekD+3yIbdPYytWn258Xd/jYma3X1je2YYg6JrNNqztCV3/L
6h7AsS28aQ8OMOiZPzI7ONCyNKwsaTn1rj1WFNQ6WPU1g7miemkc0WZq0Q8DBSQh
1EuZtUEAoOKPuSgV83hYOBicrMTCf9fzgNtFZjIz2qQnePnjuWVCRH/byk8psrau
1kIlgG7Zw9s3FyZavUUHsxspL++08OP3YSE32EDdcMx/jY6vQkUY5SiFmYkVXu4q
GuF0wPF9FItrwJcZjVxsSZyPY3mRI25eTTbiBtzAIO7c4OLq6raitV6Idm7oipav
O2kOEpZ8fw7allwkPpxO5lrHRJlyQ0HDvfqtnhtbsz3l3jMlXKgi5q2z7/gWPgyR
GGESICC1wUxEkvK67c314au3jedTVPOd+CZu9515rfzT8U3o4VamB62eD2IQYNhB
xYGEv81HzkS7Mq+74EkxU6ciReUab5+j33Eg7QDdBLSfKR7XCYYDTSakQ7gVHhv8
PJuOr5BocLLXrW0TcaJo6MIbioXflKN/vuLrYcCUpICHkZ2ixhF45Y6pCeArUEXS
Atd3aq6KplV77B3BPHpSLXjxME4phLAtGJlKTVJlTJRBbpj8MKNIxAN7dKuXYr1o
t6WCgFvbWq/673IJLLXJSUVXKXjPu2EjvllqZaPcCzt9RQG09vOqyXf3dNzlrY3F
lSuLPj1wgTYGyVwwmgAZP6MFsezly8ZYc8p7A89xYSnxNqNu8dOL+4vx4Gx+jMfd
uAnEenRsUd/Fp86MAlJehc4dN4w9HH5nzdwgFn4KvY5UEBZkhXHlVB8nCevIsdL8
fIUwareSqK0x0pGVkzKwn9owpPCNNs84CEuriLu31JtoXtEe47RPTklFk/vd214C
TLuiL2hDK7VFqqwm9KjWXeocIGQAjLEdLkXIH0Nb8eB7LHqYr55e1LSyk4EbaDsE
aOPcDYav38FBJd1qDa1E5a5BSFgECRZstMQVqsg+jLogleEIB6sji6gMIKMQ79IH
ct0/KuaXwFTvZKpMTJX7grCCzHMmvl/b18vjNvRgP8tM86DwqBRWKk1J3DsGr37y
1dqE5OPaU25I2zQMHSdKwgCdXK1Q5cia3gOqQAnWl9dj8KUkEiMdRnlbgeB0sQax
YqmP5iqRqA+UMPu4/NBixEsY8rLut3ArmMc/YCoF/yccF/0jaJen8zp5izU5F0mm
O8bWN8paR57gztaaNPuo0L9MOmMNfnF22lUar4wYlMbeKosP4Pnv1h35v8Dc/fTn
U9ULG2YBdVBZAQVWB4Tp6/nQGsM3Xjg2aqYBpY5L1mLR6xyNslAcNe5XsZ7V7Mh0
fhLaxp/76ndZsKo1v7JJOYy+i/S/uXnf6quq6XG7/8nKaoaijj5O1WwpLBdckGWV
O5l05GIe7V+rqzSo3vJXQeKmG9+LfaN8xyUNWY0MfvaFubzXSOA42T3GCMe60pnG
qyKqa4S8tCtpzOGOpysPWdQPogjAfu1yQ2RkbXeCjUJ9WGmdeKobo3AjZKP02y8n
9ajPfI/3p47GRFTOkTAbmkuGVFQPE0wvsOPdlz1DplvGcC7ppdNq+LfVW5A6bYpb
8MIOLnpAu/9c2RNoqCLkqlkUMcEpxFvwWK8GO6k7Il3l3XOriyck5mL5qQYqt6rH
xs1sUhqLQoR38f/9P0gGNGve8THncmoNZDHi2V1R8Pg2zqKG5512RPWzQRWHwY1X
atjDUsC1zyEMmvzHA4GilVe0Q118qTk9d0Csq7VEBbH8LVqZYcJHTJhFQzg7oL0B
DYb0RtX9OTfkjjkKu0yZFASCNBljYZB1wHF8gaBKmeooEkiMVPCZSyi8Crz+vAa1
K1Hr3tqRVcquGGovI1cIQZXMhV+VCKWO7ePzLGXsn0LiOM7gl0lFyES8hmMzxsUn
BgjtzVS42ZE+I16SHLyROu93uTBmRxZgyqHs4csdgoUk5ZOMC+XE1h65qp/TPlvD
ZX5H7pz1ad0HBIDqOYYM/sLxj8pPJ9xeuJ0hkKGXJVIXewyvgW7zCeOCCb3L+MsP
AvrtrXpkziGxCdMJLlTua12O5AMyp22RTGsmlpEtNHNrmCHbKcGKqttiBGXfpCwZ
7FBc6R3eM0i/eiOAOSW1ztlQIinxfELJHtV6FDvCVrIasAvWbocNTGovAmNfBP/z
VENyGbXexPBCdrOw6bz4zVElesibr9zN7LP73efk+z7MMKN8kDHqOEmAJsyqRGY5
NJNspuyCOB2TPgqIzIiC1H7cLfYq/C5/VkGVDNGVPwrrrvrNRSQkMoL6/AVxLqWX
LJ3AEmf6yhDi155+r5gUorHXnIHHbumd945hgkUYE/89K2rW8Zwk9NoPGGlSVOd8
5DtBBe7BDuTaRJczTvL1x9DLND0gwo/JNTGxYdqlW847LUCzuhfhQaAXF/OmJ2DA
dq6skUySqioEsIPCC6XWQfrnkmCGRJHp+sEFg7EAGHW1EkqWMg19j51VsI4Ow1wa
04E20DqCgSWbSCMgArvWDrh8OGYObcIh6p4b4jR2KKln69bf26/NOI1zpDbZbO1Z
CHAFNHkYUtCM6mPhT+Lfn21DSZPA9lQ2CRKYePVS6dhURJBMXdsLtfNbBl0AxEsx
s9PHGp8MREF8+uPrvKToV+a88nqQHIeEgOoSXDzvbnaR0i3Q95FgSlUyXKp7umOi
gkSOQD44ltdd+YiMLyGjKjdPc9UNrZ4V8uIJrMgv0wlZB393sv8udEi4MmYLK/d8
c6gP9zvgLNso8KZhMg0M1F0FCypP43h+fd8sDM1Quzi2NEwDHKT1MLGS4wWzKPFT
Qy5eJqLG5wn8lj0/uuiRhvG4mHPL0C+P2aU4r4tV3ja+Wo7zBoYrcacIlddf7wIu
ECIZGYXY9Egx0k9AwCn4UhpRHmyBU8sUxjJGT5VcKd2TJRsOgiOqzTH5GBU91xSB
MrZofO0wODkAuJzkFV1x0/4Yxc2aQcOlsqLpwj4/zcRkTiRW0OJu+i+/1vl0RdMG
j+uh3m0o8l5zsYFj3n8CHb5oJEAAMRad+PnqTOO5RjnQ5I8aZbRjp9U9hhwzTK3e
ZSn7rJHt/o9DyEgiNmM9Dxa6jMcrSaxl/qenTS1PoJMGOhSLJm9R5fB8HrUCRWDb
XBKWvpMk8p25PG271E7+giIYN8OHEnLikt/zCxJkAtjIeTfu51cQ0N5G9rVosKww
cktqL8W0yJ5L0Al+5RnrMfepgBcO4cgMdKGf/YvZnlNQ7+rsnEJiL8kX4YDHD/wx
oUJ2Lk//4GwrTeS1dbf6vBuuhFaYJpuPlDf/QGKIr0XQJMevp1Z+RTV74/m/d8jD
c5jYrbqbRhv0wQ2RlrtODNEwDjeikzSyGTUwnaB6Y5jAILk+BQLElsosGMOiUgZb
ofOGglRwQwrlNYAYkp6x/LJVlOnwd6BY/Ijd0OK5wZMQw6OeMH/XWrIyVdgfIknz
0CGbsu8GPf0ZV3+ihmcOQ9aLuzIjLV6Cs8NhizD32gzvx7aJfnRGpUz6RN/J5KKL
Avs5T7b5sP1dZ4Negt3LI+yRSuon/VcnfKbkbhPd2YXUTzpfKemOtJCs4bAdtW8d
Zl5PeoRbBn0/ARcAvQCx40YmOPl/mgT933QmUdu/Q29N/UZv6ZzbyFu9FJ+aIZJ1
fwtSS0LfKHTYuodYBBXWDgnwAw1PDetdiknDhdUDF48Z2kLUrQe9zJLqka30lDFR
EnraBdLtC37cXDrkaFA9zSLG7bE+cfM8qGoXMSoHtFHDui8pnqPHPdMpK3SWbkRM
bbXLnh1Bn9dVm7EbgJ2gfHr6UfwQNHcrmohC/IX9b1CO0udTe47eC8uWIsUwabFt
nVQI8/BGkDsnvmgVma/AHfa2RmIvWkbXSd5fwkCqfcFSUERQtuZ+LlHBilj9/dll
AAAdkCNRTUJ7q3nSX7YmD0+EL0tY/9dsSWmFfM/zUI3WV+6ewstpJQqgzq0GyLzC
jVnpHkpBvFb8iGpxX4d5nSWCSJFSJXVC0QLcGfJBVbGKpgz2GG3RKRB1UdD4nhkO
qKvL73C0Ya0WVV6z8GuJchtXlvOArtFqexrlJfajDFtIXuZgIlRYb97Mma3ON6Db
njGNtqiY7Bh6ggdx/qTv6LsLCRk+SWnVMaczJAEs8ObtvRzDNmdk70q2ED2LY2Jh
YwnPlVhzGq87P2It4mwX8mn7ICO1obkn1O6uBCgmqSqu9sPPQ7qFMWTNdK02GD2u
T+jopzE88YI7wq9oON4qdv0j3eF0GG2cwbP443XDqj4HAUSsNSD6K5F8O2vrYj8U
QvF5zwRwgcKJ/WQKBz9LkaNrhWMmaGYM97ewLAmfEXo/4p6HWWr0hORaYZ5fNotz
dJSkiX1c+jZcXp1PalxO57x3Yw2+M0cRKSjUTwr13zLFnj+49q89ATLnuGxxKZ3a
rAQCYtuUEMXYvzweVZN+lox/C1TU9SJUBUGdQOCXV6z0fjZHO73Q8iTRLVWzwZ90
yvCOKQqOs5rBZ3Rh+0q52neVBN1KBA8br245eoHHVcnAJd7wRMQRN3Row954CgEE
NO7iwBjr1nxQ1KsaHhHsNS0vvPQaR3TOVBz3upTzVMfa9ITHvTzf14J7baOnTk1a
GnvesDOXVTYl3NuicSTleCtv2NxFxrR7l/+VDse2qoZNbEeBEvDXFbDCsKnRP0VQ
n2/OFSbZmcMNhPQoTEb8r6gCXw+Xc1pEVWAgclPNHAbAUgmNPCvlUFEdFAfjWDTR
P07jTdK/wu5AgCPATADP5iWLYBSLb1Jmunyci8mcTSGPX0G59AHzbN8azBQZztLb
S8SP0uA34ghV2QCvROF8mQco3geEdgfxlhgfSGpLv9paaBz5J4cUs+xSCqJGebO0
azlk0L71MffFRyG/GdbVIQGAHm5yIXNbv7qrsheH316Bfy2/miSjpWPy5sbZAyOu
t1koOo60G3fldV7N0mYO9t8guo5sf6puxHOyeLR7qj2yWLZ1WxVI/HP9RUlLMW96
w/xxb5QPtyuyf5r1WCKuR4DuINfFsWw3U+yp+vBouMKuVnSEBz0USmPPLSn0m1FZ
l5IilA2bKvBO4d2XVlfp1vKOdhlGSttkKgc0AJOvvFGjlmGdwohP18FLkBSjGa6Z
QcGl4OwKiyoUz04oDS0XT4e3op1j1Zk719N5d6gYVByodH/EaYSFpuidU5N4oH0C
yPQRv9S+KLeQD6UtPig2Ahb8Wgd1K486Yxw9V3iV4mXY95TNVvk2KGn9V+KXK/J0
9JVM08Izo4v7QIoNcdQqZ99tIQHEaSUOfV9ZT2PlxIgfxHE86bCJn8FN7oikuVeb
iHTtR8Xv/gol8Kjr20wgCl+VzaGGkiKzHS1bXVLoX+RJ7xWYLcuJ2T/PtWiFw96v
jzQI9zw4cAM6irKrB+c00qbd3/NYzSfIGKaH+HUpPH/8vdVr/dEWL7PblSZycQG4
28Bba4j4KbyfuuO/dlcD9Eurln71XrFtYTPF4vMwqCFfUFt2KyPi2cb6SwMjsn+d
3Rk9gsq96umHYT1LVCBLlpvLJ8DWPb9tZnYVbu1PVAC1ogxOxFxt8PwdVoooFMf9
sDzhxnRy64UjSO3O2Nv3ka6fA/wTg3V+J1RMqhU0mIBgsyBfDkcFNwZIjeQk0avr
Wyfr7a+/HySjjyUhmoZDFvrpyxkgfqdtL6hK4CRFGUZt76KFX9NXIYq7z8DUliZ8
K/tMawYd8bMMYh6nmVt/HI9Fiat0M631XxTmMK3MObdY6LpxxOgloGs61dKVsAhZ
U5fpjci/6+dTleQn07xIeS0SjX0k5dAJSBoVnfq0RVunQrU6bxDIfxWMyVMwE82O
sgsHWqYCOGlYxjfzqoD0Un6eLoLwUPeYv3xtlnOpM/VBuxiqer/4IWZJ4VlzlMml
gnBntauj2b2auj7INQomVSJ5B8HvKjV6RtCHZa7M0JucJYJpIQ1/hQZUd/2QKOvE
VR+52KEDsQMT3F0HYi2ERiUX/rFPZ81WOFoIvu5t0ZGhT82k1h1pPNKzwRjCe+4L
PoIHFrq4VcGRbDE7+np4rYpZ5zWlLQFpPC5v4V3AY5t5ANv1a49evnA1scL04GRL
id1StBkA91iSvXGE8mEfHSTzmpjRK1L8D2V8wfoV4d77H4pUFEgiXnEtxrSfm7n4
ioB6fCRol0sd6c8Y/yoE1M5azmX2tmBRvhkxPrp534ikV4LCHA8yohPG41W3ljVT
taHNsYVYp/ro8uKpphSXLhWMAfArokMOIfboCnUhduw80LzkBM9oLNo7a77izYn8
sxYG9mPIZTGijg4rFJ5hTXAmq+xCv80z3PKLEA/5+Q6ogozYqyT6dl4RUnqb/f3o
79EOGj7r21SL2TFbDHEbbAWNHmicWBV+Wiwspng3bpN8S9KYuVCESm6ejxtD7mGe
GqvbNUkS/21c5Fi6nOvAyhCyecgoBelVTWRrt9RtCjFnmW3WIrTsbvSVfSvTotHP
XmBPtQ/0jKQHkLh/aOqfo0zNTUbdnySGf4b2+VsJwQ8dZPAQIDqQeJ+4nLGzDZf+
q7ni4OEpgoaJ1jZVs5WslIsPbljKWyGbOW7ycD0/9UP9Vo8FMAu2EL6x4Y+F8wzk
T8DngwwGUssC4KPrG7GoBxOevdhLRwt0RY0PPTvoYJnnQK7EVGAuF3iVoPAkL3Zk
WwxiDxg5rTvX+875E0ylD+hD1e9p11X400/Ibs2a/qQ+EdH9p3WFy5+SHXGJne8e
fwwNM3FLJs+9MXXk++R9qVLolL1sawC4CbcTx4YsnlysrAKYNSscbsQCAEtHN6Xs
nSmfuO8YYtdsjJQ5zaTM/oMyWmF01pFzwQeF8ivQ/Nc4Od15b242byFOm1o8X+Xh
9kUU/luIbYaZQY+ia7xxSGzt7Rv+JHIQ7rJjCWGRrTUXmEPzucFP3EVg8CxrektI
hdRxON26BC3DRjs8AoDJy/KXuhrCoJsfQbVacY9Us0gmYHDXrSHf+K/53TgkONFk
lNRQFLvormcWY+NO47WS8DyWSKAvO4M1m/XIu1Oy1f96wbymQQzPd2moESoW+KVO
yvQEbZ8wWeMta9FVCk83jhK8o4Aum8b8l9uKu2P0a68QzLtYR9LAWI7gg/5T0Uws
TtPW3GIVaS13d6Z4NRr35wL8C39Zsjp2BYrdIvSaPmv1mm8uqctWJIb0zpflVCax
HI7Obvn7WQ1QW1YREpL9BlGCymzFqV6UGC7qZP8l0IoCFTT2WBQZJMwSprR9w+9r
I9Mdn/M1xlswEgniS1zzjunAT2RnstSXoys5qsC2wmoIy5AzZc2OispSWYnhgZ2H
OQdpF8EnmEvpon1AygDKBsmCzClZmX16i/TBOXx3RbsJ3ifAAIjG9JKtatdeXKDc
r22lytE5dUoPCi+gl3ddBSVRY5TKTNV+05tSpFdriuhiM82pkjnhl8V+USLvq1L8
+8rq/Op1jrYdylSBUxML8L24wxuVGfbvK3fIde1pqT8wGuFGoj5Xod/BSMyK9Jly
sKwHYUbXT+qIWJVBqt1lISSLL20VqoQ+0/qdUayjSAcpNEJxgTEDWmZORcvhXPRN
ju9yZ1EUx3rH8yMvjGkRftILC1i0HqrsLQg2WuUHdPP6mCHR/FOCMwU652KSWfs/
dGH/9A+Zz94vnCFJGv6pFFAh0Ui6EZpLPRdlLS1U0HlAQCyhwxE65BT0Jbs+xiO+
5oXtLj3dHrh9Y6fA+Mf33y96psjqrH7xTEK+orjYjTQ/BGO8Bi609fh3Ztb2jJin
2D/MyoZZnasSHFLw2KIc3F5TJTtxHO67l/GWDEhlGr0GPaYrnlp7PimGSui7nkqs
EXO66fZxW4GI8koXfOwo/Ng2FUiKtvZLd8Xi0jJgjOduZ0ZMBQTzodIIvfsQpXQL
omt2n7bNpRRHT+kMI81DknOawuQPMGM106mqoceGzEx+9sFBg/fLrBekT7gv2iIV
wCQeu7+j4IfNpX50sIuxzF24MGluV7Kf8iqlOHQ8S1InArrz8V4EaeIX/Sdz7ED7
Z57GwEGUgEoYXXoZeem8Df/OoC5HZGrJMo4na4dwmSeKImXOdSHzt0OpLvQhf9rx
OKXGApE0vcQQxWDtZtnyg1WQNHLw5CUOTyDEtyhmh1604MT5FdFzjTEfJCtG1igB
keZoVgeinccjYX/WiNqzBOWVy6+wL8qyacVzYJMj81qOJtFaZ+I5P8D8znJ0dIAl
XwTQHcI4HbE81sObKDC9urmCmbpo9C/zGKrI09Cp+Kik9OjUzuG2pXxtBbGOJZmR
/tTXJ06RgebL8nvrWD5mV9dhIupH6noIPIYA9MNbRAKObSae4NYMgwuo4Uz53XCR
BH3gGETvk7N76VsodPmHCEhDsiqyW1kf6B5YWXPzuADCnhGg8mMkm/OEFtcydNk7
EIwcnXTGk0Gh9NKijx97+ETQy+isBBQvOTjDi7+B7yhTpTPCRIQStUUlAaxfCTSv
eY20om08DU6nDQhBo5p1bb8mIH83KsND/K5Q2YIc79e0LN8NUPOtX1UJ0Hym6gs5
Rv4XEqMerBq+vi4o944ycYi7JFPFgHdhJYH0BCT24Ft9snsEpUs4j5v0oIxQNL3L
XDP5NkJQ3ueOf1jaDfHKDVCBWzeNSTHefmjKzD9bz7bsR92wfH4GAz4LoSyrhB6E
YGyy9CDeR4Bhd1O1IxEMobsG8/Ee5S8hNZPuDt1/ssB0xeljKfKJF0WkYFYIAKhv
+sUFCc0u6G3gtO2fd/FkFAJpW4eLRGnvyZwtO4nk9lhjyypBboJx1zKKK2x1xQa+
MNsYqZIdx82R9O1EMNxmfKlxuhK2aLVgGumXL/O8BbuAzzSG68KtJS+4P+KmVD1s
lm0eRX6nABNHsMI9j/EhcYbzEXF9qgPRtSg0wyurxCPcVdzb/t8JTA9dhx0Tnj0e
i68n6FrA15UrbdsMKaFO2FB29tfMs7k0liWXCAjou/nH+nyJxotg2wPBQO07EGQN
n0NPJnTdn1ERgHtkxmmzDVTwYp1QMY4JVf9FZQ3/shrKv7VCzCJJVqibsqRfV8cV
k7Y7igqRf3Nn3LQPoFMR3NhFtnxA8DYaOGz8mDUhWxNGRWqtCUjjc92mFzi7huJC
qRS59IzK4DA/+2JGj7XyV/lEzgzDSq5JALEnl991XWk8HZcsVHophyJK0qXkaSu8
Nkh+BQbtxjG8BzstAM9Vasohi7DABZob7e1W7gGp6enCpbe6s5fJNeVPWp2mlr5V
9cxr3UDwGvo5WciymTlKXfpNTOnGa7Y3e8I2NvvQrsfJUsGnL+IeJlAY6OZz/KH1
GiQpJwjS+ad23O/+xx2Ayl3/YaecMaz3mFKvDZtUv0oJwdwB+TrnUZ+lq/EN7m+W
lMRFou7jpxpNAvT/qz3jE0Pc9IvZF+QCq7Idv1MLtHCtLNXtKbSasun6x8PhDplb
1YhTRN2FNvpRqhLTIKWcFiBCbJO0xDtLnWS78fm/SbQQ9A0sswWytz95Rc5cdvXh
9koeFZB9SAWcnb0ASWdD5YTle7CrgN4NelqBe5q6vhI6n5bxpKp4a9j0wEiTgh4x
EE3HU4/3LzUpjNFznL4Z+6J4kt4GzB66BgXXSUbvmP2zSqb+i3Cfa1YGDC6Om0lk
p3uNGRp3DCbzquwMcKboYGM4haWKiX6ZgmJIzQaJZp9weF4NcVG9zmG28PaLCfbV
jw3HqjUiqO3bLFxglXlRZVOd+1EJ2iWjAykuKJnml5hvYgLO1DDO1J/aj0Cwn+WS
Lxhz0eEKJOz5p8RbPhYY2Jyk7MnaUGMMYdEW2PYxEg4R9zH/D9Vyeryo4i9lq+yw
3U7vCR4VY4tTKY+GFageJioozK+jZb1Qj8Eftt/+Z9LnJhOG/G5GMS+dh+qp69X4
EDMasnVmh8Qbfz0mDHBshoysBzsccyOVpWuCwIeD8GNcnVQ75PkCPZYrFVT0JE/k
MgmRQ4fGSMv8lix5ZQTDNcRH24q8PBJeg1ca82hYUkBDOUSWyXnaxxgYSrTlYi2H
HGh9CuunTcvsV9zMLWcvD/pifIFeLjA7pPh1Ny9F20k3jY+SCL8UuRu6CNjlTnvU
4v2VB3clxclyr07sZm07dFZFBI+Q7YWTLZHdVX9bXPNLt53+CFpaFjXxv7dnJYrM
HDsssfbwp+VGDTS9sL/AgHbFQGhvzv90FeDJxz9a2+iq91goIObe8qJ4VBDwDLxI
ywVHmd6h2Ij4V0dCyO5MZEjyUEuiJqNO7TlXuTlyEtqeQ8xvKaqTazIODV5lgfyX
184oO6cdwaRKvuvQ20OK6AlhYwgfX9cJkBk50PcwuNuJW4ttBv9A7xKEQko4qoZ4
DRVYbkUqlwbdnBkgmNk6fzjOyw4WXl5GBm6WufWvrlf40Z+hP5hX1USHOZmhv2Ys
MqeTl3nGjGe4cYyPwT0a4vdGm3KHdOmUPkVyP3SSdpVoGv32Y/WyXIThV728DkpM
zQU33YmBCTFAxsQk3mOY+V6VqrCzRIzc/fUcZpopB+3326AFVdzVvQ+j+BSerNT2
SufM419C2cCkjFLKvXlJ8aUucWNt5pXxMOLjYV8N0Ajs7ZWMfr7zgd5Kci32gMvM
+WBqcE0PDKEI5yOx9MOrx/5A8nqyPusGCRAluApefB8cra5c8F+X+pxcx4UzVBFq
yyD9gkAUcHLlsSL4lAsQe+TEXkm6xd399IrM6f6EQxPdVmhBsgIDOfYR4yUgMoPT
7YiQbHk30MoWJGO2XPi2igPwhFyXRiCPibQnU7iGReAUNby/Tgt/A0JXjoFeM7Rb
sBKiwWrH2MXTn5cvzVjkFUNwFxYHMAJ4i9ZOJOOiGUF169xp6C5c9Ws5Gikpy6sa
lhAbLltsVZtCE9Em8JxBvgvvHU288FDgCHl84oORJ0vtife1IwjTze0tYB7EI4DF
rHL5Z40W19nt1UZ2NLefOGZDU//PSObdr0dfYMguDbVbOQ3Ewneql+6jxYlgHq92
qZDYnZPcPEdogUI0HdKcPVgGYzJ1+IiZxttD+ED0Cb7+/oIfUJfYWHsHqpvUjSWp
GpJd9xfsx9AxEQjbcL9F2DvhHjLK12ubBHWrXbyRybVn+z9snzCPbCz85XqVErbg
GYrGXaLe9MDIu160suCAtdtCDT9tbN+u0GELj94QWQ6ezlsl0OUFvHfCEXkIGOG2
`protect end_protected