`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11328 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmWdo24EC1SLhDeUV9o12ewQ
ulXp2xSZ5P2RSggIKJUy/Zx35vo9seYTXEAAP2nVUE5utAXOAtbviXy2bFvQWUo9
447w96UgZgt5E/OYwYmAjmbUN5ANvR4cKZthyHhHhOdS2vKGeOGvjPeY4fYQI8D/
EqG0RJ2+fR/6RHLZP/B3vVHFYPLkvFij27FmHP/sIEXJW1ibqGxVggewlwSXUOyz
P9if5FpEtE4nBTA0MO1m4oMxLeTTFz9PHWMQv3nLOawbxrGDKWD7sixDJ29g4+M3
SzhVj4yqet6eeRg3oWRFa7yJl20q4kHrGw915IwjhXqLiwnndb9PyAyjv64Dou3z
SEPfzF04lNnhZx/ZxM+ZZYSh4iLeTkYCUmjrY0ri3BBlpUvafe/n5k6Nn49l74B9
GQqTkUkniSz00ytWNVMWfs6HMWeRwJm5aFGfw2hzD9NOACS12IWCbORQFMtZf7I+
m7h20FutHMzpLzBYoxOCaogScAH8hO63IBCaewCTwS3BpQlYIj85mvDoKpTVtG0M
60ZD0JcHgncz8uhfX8Rs65VXrH6vIOJ51xFU+y4PVOsZMB8g0sJ9TCCVqngr8CyG
fz1QJG6J4/1lZZlH/efcV70MhZ/p+m34KcuLbiSS05WntXvfVHNgRW8quC/11U/A
4t+W3D11HE9s6Jv+Vp+ecDcpYCU9rRrp8HwvtJcTXRhQlXF6spHwf9SbptVX7KfX
DrNCX+6jzq/LezO9l9UcTcvmTdDjsTo+ubdoSK+A7pvx6OwuH3b0XhIBy39pYlLa
uCrAOGQCYbSX5ICRCFANoDs466STN3TNJtoimFi9UUw08LfOS4tsXpP3acdg5pJJ
fW/avcUDDyq6OU06CKFnaNuE5jarIcUS0fwvFANovj7wWIuKPA1H+t7ZEYLT9yfB
hdXifhOcSLHzTA52bE9TFDLBPutz4S8cUpoDBlrHrp7htw3au6SUYAgSi26r6uaA
Y5qcaLstkGLdY8dIy5IGnRcT9H12vfER9dL7PFNZL4XIb6Y4YQax7wW1KTWCs5Cg
WpcxN0bZhUAnMClNToc+f37YnCSm9IqIuBoQayua9Hb10wBFm8iFwEtcgXydNCXx
f7HtA3xIyrjfFdRBK1nlRdcjVWFnR4MTc9AqMqqXkfD7kWmNuFUfmq/uExoP9cT3
oMDzPPgQR71uFKZcLJqoLmrxB2kyeSeiijm3bw+B+c+3ox9E9StJptKv+yg0jstZ
yNq1+lMnfDhiobE+cneEXW74hvKVz4fYetamQkx9m8WV3pgOqmAbWIUbbyhTH17c
4AuGJKg5YioJnqWH1EDernaOr7B0eC803W1c4DVzzB6VL7j9eVY/2T2Gry59uQT0
9LqFwnBrtZxm5Ie8eRVcS4YYRBlJhPzgUOPu9cQK4+isSrg8B8Ywig/Vy5ynUWQO
z1QbjBn5m3BwrSaFhmILbHfY6JGAmKNcptGgahtZEG7A/0pQVnMCTIaE6On3Ryio
C2+MSXxs5Z9IlDW+U5b1L/LFpRDdlY8dR7AIuaCKSp3/DpCHQlHiJ1PXD83y/NFF
mL3+kFeSUwy/quhSB3rCg8MwKgZV96hhlaAUQKsk6F3fTl2K3dsQ3k4CU0iINIvd
M9Q/oOH4sXQBiiWebSVFm88iqjcNO3GciAr0GloxD6I5C53Y2oYfUlcB1ObByxlE
7rtEutxUL4D12wHyTtxw5YH59mcT7KrKrmkgULIU/ZrzkBsmOUCIzzqgHe0o9i8l
ZmWFaSOV3+ysFtgWxyOfC0vaTIY6LrrginwwznEBi9p9Iq+SHb2K77qvWtBclEBx
h0jv+zm8F3ioeHhqiO4ujW+GEJSZBmjZ159nR4XL6cZdoUpTgHSuE72Qe8kMqY2x
aCVqxJSinFZn6S0LfuTf99mHbUahCtDLmHtCiru9Xf22xP8OJeY/BHecBzZ8AoXt
es2I9XHQA2MFsunD1v2WFn4K2Fq3F5B2QiImxdSEFHjJMMDyLCBTYk7hp/Pg1nRY
lALxMcWAcEnmXz3++Et26AZZ3xxTtBJgnwJC4dfhyq21qs5yxxBk2W7ME7PtudvP
Y8SnAPopgtbaOIRXO8j+YXr/QLBqBiHtAaqND9VTSUcH6z2JAUDTAwIJtudm+Zrt
adc6FkJfj+UkxDsUoOECP0fHDvojHjZGRlKGN/QQOK+eajZVbvO3Lw5Yp5kalCKF
cpE0thoCV5ASSiHjNRhICk7f1dEu2wQ9DIcAhRx0xkwnEksu7gLUKcL9AQb7svI4
o/DgtJkYMgVYVrea3Qc3fkO0QzPPRU85rY9WX/LR8JZLRL6Jig7J1OIJt67skQJ8
eTQzMklbhkDTOV2uOzv7JOLSD6buUqoh7IL1l25iynIAewO58WFaxQYW2zzqfmZo
rspWf2cL0b9FJ+QkW4Z9voboFV5bnuqD+lJ62rHg7quXb/bg2H52dyEXYLzHN0w1
GqQfM85boMRC2QzwQocNlQ27iWekV+Xr1hVkDybKY54/NEe3+pxRiNUd4EFdC7ZA
J2zTbm6vehSC2waAM5agt/tqE8d5m+LJW6gs9+lomFvvMLDbVpiwPxcGz2b/A5ck
foQTiouise5cTGBq5XGsVca0d3vLHnKDWCCL7avFzfJPdDsDm+81rNeWgU+9lFsV
4O/5/8+JOZwOlGJUE8OZhj75sBYMjT1XpFhX4BeWi2Df11IA8xf4AVJZChfvEl6B
m/ruSUWChLRqO2Nm8NvJ3/mwE7/DyqCM1uCSIVPcC1gljW8s1eUVprKXrt2pFonz
XYQcMtbuHITeFWtWOovxEStkqaypY9dnh5ALUkr/TiBNE+Q2D/sd5D/BEkXRr8/G
gR4RyTZ8HDJWxDKww7YbSVlYLtk+qCGl2LZLFj/zFRIeNPv6FkN0iMtTzOCNPOD4
NrQ0hV5sJYS1IgzMvFLlN40yfKrOPQrO6Jhg+a12mQZUn2HnUmCXPv7WuO5jpMsU
np4pCRXWIkqXWaymkcFBe0nYQzgtl+hjlPcqrx7w3fHckrBQjhsXILdSxVBE6kIT
EUbjCqnpeHleJiFEO9fMYWRjTxUU6O7qkZvnyWUonJugoPKob+e7GNCkd6KrIpST
M6GCe/lQDXwBe+KiMXctoqlD0r1KqKGSqt25FEQ2aW6F86YtziYEIlGCnqMH1VJ0
+DHaJ2kJGZla3bnnvxSCouEeCVWPskOI65PW5nEfaE5pdKRRXG52pmG/BbrL3XUr
ttKWPW+5NSayBQOFvxs0+ZY34aIipa2JNbPPzLdRArHDOmElK/560QVt/HNCgvQu
+ukQvDYTXqnQ+JU67KKWBXSFJHPs6/hyQIxz6BSOJe6IFtpfc79WMK9OT990FZ+i
PSX8iZg3UtNrM8E1sCuuVLVuPrrKwNX5fZk3eaeiYaYAeI0DOgFWa2ntrPmpufiX
oNSMHmb6p+Ph1nVQRmsBaglCsonqVo5JN15X46dBzXNr1GSDvJIjlwk8Wrp8BCuj
ZHu2coDa3MvmuaoW3jChiLdzYwnMKeajS8GGtrsRVrGCGasLJF9VTI3pM8wfETks
IXEhEjnz35EkKWyjBST8Ip1cNfnT9EQ0OOqaBy2jZQs8zJN6BL2jYW6IHY1hJqjJ
EPIFnoY4D4F0v2vJWpNAlOfwFaYWtNU74GJd02pYEIaewyFiQzmUJW2GGEW8AIuI
kBBZy3CwVatAdKtkCdxNSGtRNJ5QKoLSIoPEsp0kPM5lrwEdyEVI8+IqxJ33M4ck
/39dT1IT1RZxxGIeYKx50W6Nh5HvqGF5AEDeR0iWJwLmJ9UgJYsuvdGCKPYaquWW
K8wevA7MmlBRHiqmDHcmO4zW62RDddRMPb9PUUnyJEB24LUlcrwokw3VbRBRYvzh
qVoFEyXtmWhh5nFjQZ5K9yZ1qmcV8HC3pucITY9HxodMcWzfBCe0+UTs2cPC+x2t
s/SBq028E27ulWUz8UmFuIdjlXAAWf+aWGizMcpZc6jNs6MohzFeH6UrWs724A1j
zGutbXE1aAJYOgyKu2FPr/wMicdFbd5xDQW499sXjyqOiHjZhnJobPksvzv6P9eZ
4YnOaSWrAF86r7Kjwc1hzXJBc9hA+6xWJPV9SuyZD7Nz/9BEp6zCOYR3EVs44SN5
301Ila6OL18P8cC+jUE4FXms7gE7da8kGoWFZNdnBguN21IGEVrD5n6+EW9dkUac
SrkOvrZ3OMcUqCmpOLtHbdAn9jm423QpLYfZiCGpQpQPw7au0BD/4XhE8/+W5i3Z
aYFfhgoOJk1YCcqJyuaORBr5zfk8mqdTuyWxOgxt//K57k1EUYbCZKaLJUMhShld
HmZPFtmWEMInuL9iY4ZDgXd8sGHrgn5Bg+QtH4mC6FiqOKwBiFBk9VVO6Ztu410T
S+neYqB0Db9yf2m/q36EeMiW8EDTB4bojsZQvS888Rzk7UGKyjKxtyFfXve56awf
maJWHVYwYPwPYFXPv5y6MhmJqBdpHm8MI9d+555vsipqGynLuNKBuwn7VMwVfCC/
CKotizoJEdG08zpWFMzhD/4deh7CMUupus4sGkZIerR4BlddWLHcrCmZtaksMmGn
aPbokPQf9Vq4YctaNyZGA1Lb/La2AsgJyXDNIqxH7/lmXgQOUFkzs8iivAA+j2GU
1bUvMDTyOIhd0skEeFWxPaQ2YyN/q+yFs5BmcmqC9MP3cPGA/wfC8xnQ/HZVvrEg
07KKHnkv9PFBBDyTnhz/qVwSeIWMMBiaLRKYsR3P7ZxXvkQwXOg2aQouBzk/6g6M
y3gxFtWoEfj8cqPuX9WcDS40tL88arhWZk9hRoD5g5A5eOIreBBuTKSRr2z3kT1J
LdOHvIqIsCCTqxDrVJbBhVq7b3kyTlH6IXhkwZT/gqkXb3ztOzaBrH7SMpA+XS22
K8Ql8jGAqVhn1Yqd4ocpdfu4dJKPcdqbMRGKbTDcxgUYPc77A0HK3RbEnDRCkGd6
7A+lJLYtBEHJZXqXc37EBMIK7dp/Vr6U+p8PNOYD7s6DfemWtUZWwbDQxxRrjmBx
zyM4CUNVcVdIu3NwRi/J+wekHUpUwF1uNuXU+GTZB4Ts0IXq5SYBmPCgoxBq36HR
ntdLRbEeOvBqie+mL6QxnVoav7njXdC2/FWikoGnrpMVffVLvH0BEU26mueHkKzr
63T21zCcpV3QDbBG6CQjgN8EKcply3JOLnBcW6qEphD1gAXovWQYgWr05Oowux4s
+1IiWfCcvHyzvq7uU2X1+5NU6A09xldkncIn7R2SEGatN+v1VZuJJ0L9nM20j9V6
Dlta2/U8Um9G/EDlJzFJMa4UYq67VUJUNVsqnheAF+MeMtEdE24dlKCSyb86VAZN
lQyNdTlV8g1T3ShHZjf1DwngltsMR/c+UOLi8HG0n0BzaLn3E2MkLxn/mkljPQVT
7TcTKSZt1C9MhFtjeISV5Dy+AQiyLr+Hx9hM7PlGX1yno+sXbepyOTiTVtFn4j2y
4afddlQmWl2ze2/YUF2k4StlL4E+9+NYOlj43DYj56TuBffV2imWyL7H6k0oNk16
mXegMcef09KyTy+fyPC58fj26Tg+8ufb21WyROIspwNp1+CYQv2EV+2AV+miZknd
91KMKMFD7ydsMcudPP7NIoLF1jG32gyOTxaC/n7v26tVkvoeyVR3lAPzxM40gV2V
nmgXFTjj1dIcGZgDDxLXtRUspjp71Bd6SgKo/GJz+DSs86e/2NZPT1192sKtM9TA
jwCoEw17qRNZiVyhMVmRZX2wkn11inBjca+gIT/sTgr/W+lcvM7t6vxPyBgx0DwE
ijMKJXX3itqqvaB3j5fu974+Ecn+g7FshR3/PQA01RFHGIWNbES8Lei83C1alfoD
czYbDSAsaWolYZ6cmi2sbrCPpjdHyP7WooI3TP+tEFRN7LXNSMMa+PCa+eU41m5h
7Fq7Q6SA4Hr93RLq2wjcecaHv5VIp/sVCU2Ey/AqgQpuoYgecewmvT0l/qNZF057
JkuSIfMh5LKUqzUnnwLBMeRFJOoH1PYFexG+kpS+fD9vGvFFn7J3UHCJyzJKpjUX
Nz+hwGFH8YfKxKrIcu7mhBljDMa462s3VB37UMJcFUwgz8eSnl5Cif3s7fjGnIU+
deyrAipnH8sNh4w9miXyp5l+D7RJA1GOeJHroAfbaOL/r5SB8WtqJXEnxvBDMs7d
VhbsYo5vZ2NF28HxbIQCbUwQorMs0EoQ0qS36jyZfdNffejyC/c0R4v7uzzVVpnH
NyElnCjAojcE0Q9NgETVnncWBLGY8M+x4vAM7AldfO5QI22I1CP/qDjc5s1U82r4
wzw8j8n6U6krMOiLg2WozG8cUbHr+FLSpVVg75cYIeq8Og7vM6+SzsLVoHEEyBop
Mc+yrKVqCH331uAlXxKUO0r5LnJEfukNvww6zI4SV6j19tg6TjWKj6dqeGI5GPnR
o1CeSjBr3CjaiT27olXdyo6pjkgNpl1vZDe7RRKJg+EN6G529NakS8NpmsXAlS9/
HuEsDHuTUBOPRkPHEdhkqY4HjamVDWt/+hTmitz5mSAfg5FWq1f03lGqJEFIoPK8
ibDuEsaDDL+5qUjizIZkGDr2cXvGtlDApZpTSSpWa1WvJ2mZGfy8NoArDpNexdUQ
Svbzgs8PRCeIvzRe2ZLALYNX/NNY/hAA2uYabB8Drt9UtVyq9UPFJscKhA5ox5OQ
9xqqN1gw/mAMNEHcHx8zwbg4Vq/ZghIbHChwLyg2XauLc/qeJlAwed+bzr21aFg9
vMdqcTMo1MEEUmxFPBoCp6Z5PCeP6vlVE3f9HK/wL/xaECEsSFrCq1ueQ4PAVo0t
RdqoY468m7wJxQM8NiiUOGz/mXE1OKbRznmQ2q75+Fgo47vOBKoUj88IgA7PtRwG
7iV0aCa5fjWDCq396NUAYlwRv/IdyaURYmDy7qVJzVFXY+9eOJD7rpZFoPHywtuE
sE/N2JexMCLmz+V+sJhCWqU5e2Bc9z3B4hIRLUITEkN76mMTw6xqFxAfNLWnmdPj
V3b89YgIeG5rEXlW6F2gBYDejp4b1+uZc8Du4FfSw+uE4Yt10Oamr8zBAEaDncxp
+pL8ubKu72PRsCY71TsiqlUWBIDSRkTJBwrk0Egn4y4UCap5r4IKMk3ea5mLoer0
iICpYWcdqQ0tyW2uoLt7Ps7YNNWmNYmnAKAo7x3AiWgxgga4IRWf/hGltSTEfwYj
45j9cW49HSqm5hf8H4cN+n5O5ao2Blz25RCIqV9vbDfSm93o25akQWQT8aaHeN8b
bGhE2CAcc34edsHiMSAV3DPvUIL3E7PYce99ptuaOy7M3qCGC46CuQ3FXjx03CWn
GDIJ0jGHswE08KZCgxTw9x9RAG0NSMCcQj252hixOSDUAhpniIEpivZ+SikYHnTL
wI+p54FhwwaAZ/JeqU9SsmMRyCJRbPhs8t2kISA0xDQrkdOQt6gOTxW1mjIeITAS
DaQuFhTov/Ko5M8sUpLuDx34nYR0m5Ab1D13xbGR8gvBZHXRdXHZNwPDev1xQ0MZ
5B6bkMsX8WsyXFIJFZxEmQIM3Egey3TDePGpONJWfRuTBLreXzX2pXcsc22ZnoXx
5hFtAQXEGBWRDVeSpEPWyqzNugQfJFT6UJCz8GsVvFJe8WrxZkbrYHf/b0Gxrx3K
+CMxbPkWh2eitpgHzdDtRzsnOJELqwe8HWkvsfhgXPTsHMFnWbWBpXWVY9+Pm2Kd
gdeKzpcd/sFjy7xFfyXl1a/RRb+esyPMK+uydYBdcGiMpOKjU7jH8AT5BuH/XVEY
96wT9dlzeKl1borJNSs5S8Tp98z+rBMXKvNnvBkPw+LiGsB89HBnGlS77JJyUWlW
JE+jmu9C7hjZcPYf9hi/B0r5mmm8wBV5Qod1aRf6gfpEl6Bs3YqjBbWs/3ksTb/s
g+RssfPpftlWL8+E4q02i/VvyEJJlxDdPDRg6r2RWPRe6O/zusJBAJe1FbvwoHe2
2nGJUv7prYXufRgFgstcdMU8rZ6w+84ySJhKTBv2vOSesAk2cHBme+Dkw55+pPpz
4OMkngeV4WOFDuBw3kH2MzPGzwLyP0R1hXYK4G8ssso3jl61nvpNE9TFQjsK3kqK
oFSbLJXCsl3bFegPstllYpOH5R6bMgdPCNbot3lEk30QZCOHiXjK7CC3AgP5Ksk4
9jUQh9frQkbQLldmqqd5Cp0sMzdlqhaYt1AM1ZfDluvG4Is0O3dIq30fJr787rX8
SO5wBFo9h0ligZUaY1IwakBuMzRHnKLwlWY28E5iFYJy0bIdqlEpJhpnEXaQMCqD
z1udfn8MLcH4rkkVit+97VHlvGvbGq69FWkRtDnTRSwSUO8R2KDgPfMXFPR1z3FM
OnJxLrDr2HeazNYOBM2OXj3qTmTjSZnKxm2yClRBqf2FrQdqwyIaYSqCQtTihoDA
AWDNssYfTEOJseDRYgduV/c7KXuiQvGQMIjIe6KBk1ENwNznAtwZdQ6KX8A31mLf
ayXPYT09NrM0S8Bfr4REokWZ7U9YRrzpgQ5bD4m0pDhC4QvD72eE0FqvNHGqmR6X
G3NO0CfeATJzBCyIikobm41ITmvUzMLJhORfVOeEwjSseUS8qOpsUmnDyrcD8z6F
krQqUEy5jRzI/ANuASSBswXwTyZrLxzM1qKFkJmwPakRsNPEO78501YmfN8b6/kd
wXNLXXiv2XqUk89lOAlxWuS8n4c+jSvXwBHibJSGmQj9d1V4RnWRfa3z+S02hsjw
L1FSMYeYR41WiERrGvmYiE0Oax6REeKqm16Tsln537xdMnXQS23oTG6AkEERuKFn
bmrC5XbshUvpCkSEeXql/nbnL56TlXu0pFVaArDlhphsr3Y568H+nSO4gfpCqv7X
rVdSZQZ2LxzUaRaJl/M6rh/rmZGDyKeUP7xnMltm49Yj/fdob4ZrPi3p9kHc3O4W
xtIUrpwbtgLNcxg8VbI+k00+h5rWjsPNNgM18GrcfWl/hX8L7w/Ij6me++EmlgCq
IcqJLz9k5jv8T7sTpUamjEA2ZaUaYa5/kI4GhN5HV2EXTzO5TrfOZRmrezeJREuJ
s5z27AfFdJsEeyuErDbtM6MQ9LC6OtprtyjAbcVqwcUvoOSt3h7X6gaOBhNL46wW
lsg34lPZEdnC+TU72kI51Mc6yO5zzMTY27O19gObnjDmgomn/SJgfkWZu9lNBkPr
TrQtXp6Zvo8tayOgOhjOZqh3VmcwnbTBF4U1obOZ3Jjoz2a792+e7nACII4Xt6u0
qIZO5R1Fufgu6TKhcvtCh3wCzvn97e25x9wD2z+YAMeVFuqfHigqmGnwsyq/bVSj
pRLHreIbVVLwyPXZprmxRZjtfd+Wl658GoMaLvY4Oig3FCnX5LgJXTTQ9mcmqR5Q
zNPyiwR+J2twa+7dS6muIClsSk3VZyM60/W1+JzNJoqn4gRHcdtCh8HWouWrMyHS
b6mzcvoRVpgFcK4E7+nDEUD9rIQEM2hmutaL+nzshiGhXgZHL6ReZAwDDdn3R4sc
L1CxWcs0Ns9jdAVHNoI4F0HuN9wFZdWijnIemJn/8n2axnus+kmwJCPP68GvY87Q
nrAcH3wkSIA5y8ipZ8R+U9UzGLcOGLet7nMgAfyVHWo88KDqc2OldCD4g/zSVuDH
doZB0clzeDjMHN4tee44xo6DM3BOdA3S9K+2CTXQFS49c3e2RCscjYuFH/jqYghk
ZrxlV86M+s+QPHbYR5kK7gD0ijupj7hy4MSi7YmqmTvqeEKNHc4Nd23hyyLPKS4J
Cio89DVzynwjSjcFdhOhhLe03k7v8CC9aD8mZT4i8Hy92EDBJitod3mkM5IWq4DA
jwAxbnKepK/+/HQawe/aDjiRsUj1aJCHD6mQGe89m4tuGKcmu4ZRWMNqLwUkukuX
FW3pV2Jybf7SpptPEwFxYcTC26FOF0EuvOEPHq3ryw7NJ9SVfBk87zpcUGPcnIaC
D0Lknrap2ovV0Sm69E7qTsCRA5iXS3172bYcGxmvqydR/dTDZxxnxRCq5TGq1/Si
KOo4scNw684jQF8rEwAxTDrd9/w0i+J6e5ESVcONvQuoZQX2RaWKgXVHfMLrqe4G
Jz+5AktkE793N56TX5UPO9B0Ch83SU93AG9RXBQ8VZLy5Q4AW08rqFAOoI9GWXuA
erOifikZqkHyCh0G40VMQqV5C5mv4KxE63L5dnq+rvo+RUWgRVkTJBpLgzxRTgYW
xfx8N+b3+L41S+Dm2OnQnLZs00ZrlnRT49lsLD2I82UmFrp9xFDVzFxu98vlylty
F070BJCp8g8Jn4TtaTRy7OfQ7dWMLvihNiz3LqDlUWneEBfRu31zGGHq2ENlJ+Tz
8dssR75tSFk79vA/P1zr/N9iY//vE5bRkwx3/OUMpB27t02NIV+vpHNLN5s+11kl
RXUPxZaVK78AGrjoSl6TMQ5CGBOv0k2jGQxgjq02rf3CV59pYnZt7g/cgmdPvvhQ
qM4nIDHx8DQkEwbW5Yd2qLKj4t00u0Iw2kCxFu0eBKV500ReCuzJZWKmUokP1Pcu
nR2FkMReDdth5m+Fv81P6zPawJdMerZAGngUbJ+gzc9KuNncED6D+ecPwY180dhR
1/dH/Kn9W/8fnrFpfOm/PYUHgAJMWVdeoVIovoYj4+CGJjFUCNkf2YXrcL2Lg2GF
fClHDiMurwRZE9GTpGPEbVQQcc/KOatbF8ezP08/K49J6W5PS91Igs9wjPEmALeQ
PTTQcP5ueAmWf4ED1+pcLqlMo2U2OavTUcfJyDoKagB2DJPUPkYRcFXk/0sp3+iF
5n15xtlGblUOQ3+wUAGKoo5J5KBjxUhy5JwPDW0P1eBSw6TpPuYvmkLb45EkwH8L
UVSQjFqEGErTSFJBnA26ZOmlXRoGhXABLdGmf6fXSS9Fxjj5eVR2E1ibZOXG6PUA
YMt6eByEa/SNdur3bzsiedDoMp9VkRr4U9sNMC37s4TqtYk/IKbCU2em3pR/5jXU
3Rqa7Y4jh9fOB1PpsDYuxOKKtOdMHfJ8vm+ozUvsTH0TEbqkc76kw/76Zcutfegd
bEqwjWRj10Uh7PcHPiH9TE2OJFy2XOYxpOmowzR7HjDGRe1qZ+r+emn/zLyPEc+T
BdhO7pk+H5qH7hAf0TI9y7VY8gwdOEB8QiNN6C5mqAPFKay3HU73fXDPubmmpyfd
r0e907u4TNFnah635AGaj+8kvgoDz1M07/Xbshr6yKiDB5Nklj3kAkgshWxfvWL7
u7bt4IGKSqKgvwPl6m3kNrkKnqusG8soE3P2m9xfQVTcEb3h4AARsqqZpzlKY5ew
iy0la9HPbG3xgkbaykB1e8A8L9WcP9KJpiNvC3P9p5toGwwHg26mjqQ9siIj5wbi
MANDabOSm/RjwTe11+ABNS48kK5SPDVfeIsWuPKeQ/UUWzeYe0Kdh/IETq9ynE4I
p++C06cFTcWbvmXlufzD8Ns025MNLxDeZUIbDUUfyuRaovoe7SdYuKkkliue9ZZo
zAvwWaI9PQHPHn2y7/qSEXew9Az3yM5N6mQk9dVDg28dWxj1oGneZBPXakHSZz15
vbAnb/+eEND8zoQ/UN+co/yq0pEpodRpaa2Cnj/QM5NwrSpWHTilCbVMzevNWGpU
jYL0ndRCHXol9TFyNVT4yufQMlPpPJtf01EBWbeVPA3hdFRx8uaiABdynmOyQePM
od++iN48kH0sSuqc1ANxz/BkaTgNMdMWwURB4uJ5x3Ew3e+3PpTsrYIPXKhbiP49
hk38n1xVxX80ImbdlXFf1Uy5ByjJX5wpBOHbqAo4h0gzPczHqwPjeNhCgJtjtZYz
l2SWY6Mmb3aoJmGIOASWOb0v9+2gdaGxuk9fb5gV8Vkt22ETWUoVi3vavT3WFo0F
gw4ekH88tPqYzZ5UrooiYk7hORxw/fZqcGFP+otBwoJ9ImA0YtLkTKWSl1mIH+Gw
vIWEpyH2DH6yDs6t3Xcdyj06f5YxgirI7PoFW81lTSN1LBrBtZjiQkazozBwdsWo
wYP+3YQ4ksYWI9vqtOg62NyYFcgmkq1gu2XmunJZpdUSwVnNiuIF0b6LfGw2B1id
+HbYPhvQlcoNiCOyGtrkYbRGnJzTQb71fE9+ab4qajMx0f+PfgYH3Ux93CTAypix
AQmeIqxye+DEAPkjiqYqd82VFYlPyNxphkh2hbeVHyySdk18N2dP+e4q/MlUkzLP
Z7TIwqU/VQtxhacG01rptyWuQhbR5y1k7c+IJ32nPpJA3KX4KzqJ4dUb7LxZFC6I
7Qgp+jb1Jx43rRbYQnd+to24cwyL/DJo2kLBx6ZaieF2e9oMuDTo4mCQROooLEyQ
KLZEiuM1PSkeDYFIxwKUL9tVSFAakikwQ7lxBzQ7tdgyYjRwtbHoqKV/KUPFlW2X
QuQu6o70Jpx82x96jgasD45yvvStuGriWJ7hRsPx3CN38Ktut6RTao+Brvv+sPfJ
4GRsvauMuKXAOypdGSxwIijpdL3JgUmDfO//kOFySiI78pJC1jM6S256MZnlVhQR
6mHxTb8ms/vKAZoOQlfOXtCiG8xkxGLdP1yqk+4JOjSu8PeKE4WR3/bQxhsBxBgV
brNGKgVJ3m9PlmhBa4z0ZIEc3s7uH+EFXQjMhEJKVz2sRZLNIWp4ZnTBiVxi8PAj
p0e9w09rGHsxEUKavZEd0PV+Xngv/0m39OSQuwPUVJ6kDFiIMhheUOBnu4XBlFpg
eAMyw0kUrYG8TXxjt1m9yBhVhxNaV9kE4oDKbvyfUhMRIOnRfkMGsK1wpnjPodWD
F/t6lX6VUCKPT/zpZxMPbl9Hm8bWF/fsLk3Axh+SfYR8sA5P6DjGAfOD/OjQOR5y
fU/pvOXzrRvMGriYHW9ubBWnQS2EYCz7xVcBcR7Y3rsUurZvsCqv3ylZEfnip0JE
e1vr/KAndw5qh2p7B48evWNPAZI8BhFOgoyIMUBot4OhylDZqM64aA1jw8KQ1lR5
IfT4hKZmYIfEzxXD3maNMYUGsu3EKzYrVXOw8kBEuPbOhGGWaKKf/3274cSgRfOc
XU+1qd0U7CxbA6NJszPPgB3xKhTiPFJb6ttSOWHRa12T2j6dsiSpGvA93iaXeyRr
TsJPuvjNMyoVJwtnUaWGbc8kP3HaHtfHQh9Kq4OQe9AFQPoteAa31AyZL9Q6/N6P
gjAz6G/gQv3oGTutU2mk4p3iOXah/dDMC0V+RPmb235nLKjd8pZyCWQnYaqOmU3Q
t8fs31v9vP0NJsyZHof80CXRd+hWaQE9tplRyafyMEqLgwDF6w32d/pUt+MdLRUL
I7HJ2Qk+ZOuBL51kuPpd9bFW+aOU0kY49tDV4w8p9sMGs3qXcCu1iEo0m87kHYKM
9UyaquwcgOb8cyQF5/+kwpb3M7j0DGkFmjuGMjzdrNU2xBTOq4CshL5pP7fv6nip
LXBVUKOGLBHGPz7TZUdxtNOf8EVS1S6tAR7Mo/2I8fNmtTCTgDbCE2kD6Ou0cMvo
McAaqzkJSYlybU8aT1kwuR7cOl88Glpf4ZfOsfrHwP5vTMxb2oZx85MKRpG8DzxT
EQLjsfqF+MBkUOMhjeGeH6lTpXDuzrBmGIawKEDDhgPOOqhKnXFQ5yz4/iy1axRq
r5DHGDHc7gytdopXWiF1AJrZxVzsTFVLgl1ehnKPXwx408KwwGYXqHK2Phwwcvl/
BN+Et5huYFXUhmHuXk5/LHMdzt0ECYOCaWiasg/v8RZXZoPOfmtdZEQnyGuXZsAh
toaqZCNDCvg9W8FOWGOLTdkKTGo0gP+NWfIWAiSRFdvRnhCHd3uB9Qsw7Z+/Dcbz
EgWR5S/sOUG/7PVNxRLPGsRs7qJ9FTFNX0TtovZ+uvZ6O9qNWYyPyQy2V6u8aIvj
gOL9gCsOwHgcNqyIGv/xTmPbaHTaUgRcumrGI3Yfa1jzWguBgQAilP8XIyV2u/mh
p5EymKdOh8eLSERJeyH0Iw5E0qkaOEzjCkD4hIPziIDqvYHd0qt6JJVxPllAGHFs
/ZNgHiq+FsSLpjF6fLdnjXCMijUkvl4Zf18FtcTXuD3zRqMp+4A48u4bQU1YLdkX
7gKUBUhSQEoOMHJkqiGzA6/aPklgVmLml7f7LRQfl+V1AloVqlKqo51QWrTZK/tk
wWDnLKWu88E6NVlnBPDzze8AI2xjilmiK/ylk6C9CSKqlbnr3G1J0m19uRLBNfUq
Tv3LNoMQ8mOzWO76hq87ITeD0Eku1XCPY2HHm9l3NlD4ipRd7oJWWf0CmNzl4CIc
inc976qXIJqoiHQJXiHJnRfRk6QP1nr/WrwVOeGUnH/8R1hoHkVAvqWOcdXgBYuK
NOASAa1DWlfCxi3TccXNRON0crhVSyTQYXJVplEMQ8q7vP7zZX2SSuSlnyZ32qkz
NPbc8kaWOFT6ffszBgmtIp3aGKSwom3oCUN14RXHmb7U0cE0BKQLUApDNEkVpd24
34UOpYCGRVowmLSh98RTYQMEi7/t/LKFU1qDrgV99U4CmJQrqcTyESen/giY2wiI
dUuI//xwMFM6snIVjjP/0k9e8ypCQKxi81HB2+5z9c+Fv9xiS6SfvNB0s1WDLCUa
b/uT1zGrLW+iH+P6HiLQUgsjaA4zNDOoZ2e/fw+7szZ9JnbGbBGQ8LcIteRs+/JX
Jef19Beq201MId1WHT4D/0I4GatZJwkdThrnN34XCDEKn7FJxkJ+JnaSRUfng+kP
IgHehjTfYQhJe2pd7bK0kkh0JC1jN7VUtgta41brwodcDSTUKx3zQFCxBZLXrrMm
jVbdepUFg69uDLhsKZWZuf6u6vJgOf82HhVDaFbSp/+Z47AD89edKIG526L5tDvb
QtnZiJUQtC5U9FKPsGMRRibFEY3j2CAF3W5asGmP+OlZwwAW/oK5bhRl2tODwqQl
fuBq3t+Yxe6u18p9s9+C1NBpI22x/tO0DmKwOM9gd5Zz9auxrXUStWJYGZo1Un3u
5vEaL5b25jNOWvH+86g9BfcN1kbQEeAACMN/iZA8pGKPTc8IPa3+FYcwhvHcf30M
`protect end_protected