`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 61520 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRqFIMsr5emsPPVriiUzOHE6Mdmt4wM8IGdRVanZqj+XL
r0EgfexcE+aZ8r4Ir17I751pajoEHmULhHVJHIjRzavrAeMVnyM3r4dvpKfP3m1x
ENoxy12n+QUtcx58topsBXPt5RHtv0WUmSGlH14SEGD/TEib0dpH5IKqS2qEks0O
V9hK1PqqyWhmvRkEKWvvFGfHfWNRZueFJBg8HfFHnn3zY86TAiz+wy+ekboYk6la
Sb0vLFlDwR4cd5RdGY+GcLySVS+E7C8KTw8GNoRNKBacnVE2LSALZ1hDRp48Jy+X
LnOHqXg/tqF710TFD8kEQoZ5lElZUkD2zKUZkd6XBo9DTOxUaC9YhC3qfniwAxZ6
myOw2fsoWsKhlVk1TBAFkU8O9OU6bIQThkN6Xc5IBHjlGgIXpZ/WrFeK2RNb3plv
iOYKIB0bcdJCiooI7skBZ0vTjkOBQYispA7+FIPwyt9x14DgqjFqQMjuCgqZ/+ac
/ruIPO3/f0N8Cs01NwMEv4wT6BRKciQXt1eCZPMAZoH9KwjL1KVjT/KGaGBDZ1oU
SnPvSl6m5A0ZJ/MYkhXikNZc+uBXOWWH3mVXTJ14t5AqrvWgb0flLib8wX79r4Y6
BFjtYbzOoETqbuCLPBsmmJSjRhUvX95UqDK/8ailDESKIrEONuWWWTIgZWHPJRs4
7jz5imAva/R74hNpEFPdA1li8EhUoRDtBiudxyI656IuOevZuZgN6RmB5Sp6Gt2Z
qj/fKWgk9BJFDID/BBkl7CrOJD0GPofKKwxjt4kSeWHk2BB56iTE3T0eVtQHsrf0
nFI+5YLrK3+zqz0bJXSliPf5DWYF9O0mT8PxZWB7cyzQv1Plh4/eeBgPL4b6qbsk
eVLy5D0TyTuVV0/l1QGZHkyjmwCP+2M0rEsqaH3lhCxPtMh6FoFV3jHf7e14qVpH
hKePUOjZk7chn5CFYVLKMmG3uKoIJgY/Qk+0s0bIz3yUQACCvlwULjt0lSrpj4cg
z8ZOnOtAFsVUA6z8ik0TyRpc1zoDWHewooHJhIoyduUlP2sSEMe9ibQ2nEYiollK
iKTYNOUcIAr727BT8lPK8VNRg0kVFwhQFeYIROLqL4mbyIOHe3CpQhdFNaNya+nL
FPzijym3jQonFeZJIkfUkzz++QToZ8Lt0akxjwG5n5KR24BVvKhTsw+xkIo9jvwq
wgjeldw7S1ItOE1sHsqlBdxe1M+aSVgh+A6qC7vAY8c8TBh/mCdheFIx8stuo4Fh
RtDCfhPluVV158kAsV1RjEUCTHiGVKK8lLaeEsfqyxARGVaIK5OSi3bRYg4nOnjo
ImLRrh4CaLfrwPRzHfAdkvaydWKhuSKdcrAq9l8jCoswjlrwdKquoj67cMcFygfs
If+T2/hkeOm3LhF/qDKz5390SCGviBJe3QpbmjBKDzBrW6ENK4zxWDVDzx/3fiLY
UMFMphaZqx/0XAK/Ogm/R3T58tjoRZa+y9agb7Yxj90g1uZJ0mZvHxyDBpmz5YUO
xRriX9PLlO601t0W6THBq1VjwFAm2SBcVztwOYZuT8kun3SKuko2PWMcthBF7Q6T
jmz89vS3ZotMNFQ3gc16Xx+NCdzyHPww6q6gRPIxEnNY9fCqXTOkdzv/Nw+f955l
XSIoqMsUFR4vXmj+8IvAqkNtqfe+vOqNT5Zbo6ASs3da0k9OidC8lZ9qZmYYAj6r
PilTKz5tPIrSyYoxtrIpSBzmr42fm5DOhibMwjIXYX0QIAs7mr1q+VIVrkwe5kGL
s5v6nAyAHaB/XnppxfA5FJ31unnJbi9nNyFBPFdZL8o5T8pOAOuvf1dCB7ithr3M
ImyMeM5XbprNswRJFl8i7cyWVu3hGGSzJEhgp0iSvlxhaFxxgCnOm2ZVOcPVGQAE
RHP/Z2KuP/jKjReNIvKW1I132ukVMoiZr88Tq2vInkmSA6wN1JxdasVGUrvEVPUr
BfHD+ujOTOFLO4u7NTKuqG4HJFgXRfkFM6dhQ7wb1Qap5iphlYqpeExxn1znCSkn
l98irmWSgYY8LgCnJELm5ZNeAvJfPsajDFfPh702dUlLExjAMuc+SaYrZN8ZxKP7
LHqE087dUdB5DG4CtY9L+u2aXYRJEmVKEJt/juzwozn8wXU3yJv4e2ay4/xICJar
LdFpO0js6Id/e2dplalfOIAviSybiS1SyIe12qWLnc3R7zEeNkP0q0mkowQVCuFa
FW/qitQ78EC3ZO2CYCsbraKwWuXrla//HhD8eCm/JNpqI1xSDUW5O+/oVFB/ZTvG
+1UbtFCKbchrgepOBYoSy3dJ51f8n81SC3m4ZyqpDfH50UO5SP7bMTmLrcz5LazW
0PKS6okT54Ut7CBzLp9MW9ZjUzYsY4CQxnhaQcxO8QWRUuuvt4g/nYY0n0ZqVgae
yudAqc76vOs/3VgLIVb+0wmCXp6PY2OsgBGvyey+AvfPHlB980OlxqHUQ7n242k1
yWg9zJ2O7jloQSSJ/DHKWZgaDQAckZxG2QlmVr3ZbV3sgRtcqsgO1ndHTtkGdhYr
BBPdB9NnxUv3iXvyDctalGjWh/F1eo8MXmFzaBtPMpzfyvYeKliOF+JFBETT0D3B
4EbtjMFvRigSgtqBGTPvtoAWcqG8pF189FWAX7qQdMXNACmMFBHPQ95oMK/91mzG
VA/eln/Zel5wjZgsvRLXu5WsZHCf91ZTooQy/S1jg1lDdi1HwS7u3YM7J2hpxTJ1
4Ah6e5cvUgvJ3DuuxryKWMvUofdRFN8gzfC1cJDxWjgp5H4PyCEAcuaKaypS/cTK
gdH98MNh98ZM9tc1Ly045vrLdLwziumM5WzbO6N9n+HF5M80D/L5uqKu9Iw0bo++
yLQQ1xALc1wNMKQotzAGPud8zDChF7OTn6z6fzhWEWHi0X1HcVha2XeCMkEpl8uO
9t2UijRwNrz5YgJZjbtyD5F0v4ccTGChq70Uyk7HBMZOruWn6l27ZTPlM+Dzmmbd
1lRZk9CYwoIoPBmNcON3a0JAZisRV4FTw6Nu/7HDJ3hcsiakZf5x7nR/2KVovXxB
ETGU8IsAAznKjiV/3E/PqiIHfoDMZPgyLEqhfl6C4ZRvRC2XwF+cfi5rMiWtqBQW
mGLqgfODK6XPOQywSgqrNfrC3pp4KMraWC1fhdvxnDRswAoydn2n1Q/rukRxgf80
HkUzAM07/vZizkWsEEiYy49Y8Eo/2S9pX7WmuViHNX2I2Hksl9BMKF/eIGSp0PNE
/ekhYDaee0m/LHct8TtI3U0WRVgfAXhqZJGH0Ubk/U+tePruuRXrXGg3VOJ9qipz
ZUtYdhQVCGKJBKft2xI4dlxGg3aA413pGe8bC+xZHTqUASyl3EWVKsRnPuCVlixD
xex8Uh+buZih7Mh+wVnl5dP6GTRMyLL9p17uRBYm5B73SY26X/UTwWhprqgwB32C
hhM9aR//dGlbJBq+Hq+FxvnOrBDDof9PSZCcqJH3zPVVm9EFQDfVkdh/ane0Nh7C
YyphvFemLjfSEXRX4xMROcSB4lw4oc/uImovAEe7Gg5oMHh7l56+Cs3rWaS3lzLm
YZOZyUU6l7xz8qlK8kOONiXTp/LOxplZf9xCAerYA7iyZXhKjNI7W7AJ3vQXuKVq
OlpvZL4rThG5/bWtemLet0Rc5GpA2TIMzoX0huTWla7YcmCbQ83SxmlOHH5jIxdX
z8mYML4wKhoqf8DVLwISsWAkv3PVu/uv+O/3e6x+6Z/T17hzOpFfKI1As+gv7lIC
3DjhuGamE/up0IXdAGF/7FmaHkiusRAGWuFtdxbnpPF65cH0Itj0qg2g9sOZgi/6
pig+uv7vZoFNRi/IKEdkbg8sxLmVluEgt4qQDNH8ks7842U9affmkiDh5mDxCVnG
g9xikqG00O8d/NXjk+J/bc5nT31I4rX54GI+ssL0SjIl2MRwsO0ZfOkvLGzRevsS
stdYI3Vpz68/SFJNqa/kSGa/aUgF+JRLR3RW0BCGu3K6JBbqNKqjqcDfet2VD4dD
2h7tj1yCR8XqwZMN1+Tu+BExJ6Z7Jh1/dYqEk584MPavKvJX3PKvgTdNOUopuMB7
wjDCU6wA7heV1To4FRZO3pJe3/R2GA8JUvoRSJXSAGbK31i3oBBtWdZeu66RigkF
78p69rR3li2v6/tMBDFaqNnMdtswklEfb2tDK4sgZMrh+vpovrjMjaDwNaq+JPx4
c7OUxjrJ0pGgOtlQPJH3CnN2GNFvn1fo1OomrmY7wn5kASegkdUYS+rHkzd4b8y2
4dmNhWvb6AAVts/3fCq2rQJ0WSdU551K1Bfqjr9rKMxe7POm1yEckNfvd9RAVUHX
QirbPdpzp1reCu564mH/RfZHYzDGSVimekT20Qxk96LJERBedZEcN4JBEJ7RxGpN
IyMOCE4Fv+eUJ5n5v3KgidDrxh2I3tchXwz5+tDXt9imusuO/w3tuBALnWrvauu4
fuZqCGNLsFsDHYI5NvYronV9xmiw15zwOm84O5S+TyM0f5JWUdY8qy5yTgOPeQs7
k05kOm9mGBaEHeqcKJdoYYY7skIiXwA6j8jrCVv2HdSgK/VleTPJCPl0IWrNBdwX
xpFxVtPCbIvgUJIRsjukrobLhJwfoAEQ2cugfsBpbIcMdgmTQ2B4ugnMfxgQU9zT
+ITeVJ8C5Iq7dsI6hQh70SVEf65/jI4w7S0qQy7RV3VU+NjozTbbwGqS2P3Yk465
FpasqkuNnc25IsK/zqriC1C5h4uB6dF4EmMrHnGYHeSigvYGs4JTPH0szhhEgE3W
OAT46GySi6WUm2v5xn5Dz18cI2E8F0ZY2Xa8hrSrUQD8M8NN0ulQcJqK1LG5OBnv
uAb8sFrdEKuy+bhbabnJO9xKWoLtLBati2Bh7N7UBA0HLL/PTbskWSK1d51cEDaT
Ijz6RLQMEGR+y6gpYoOxTk96qdc7xd6/Oi8LgNHnlVdr2zSXjyE+dyfwGXmdKpMr
WBg9AedNIrP5qIjHHpV3sklq7fRk1T6tPLyxjHxsN+66qtMAJuNJmE7yqeVQukL3
oyKTLoF11F0bxJR9dGA05x13mFX4kQemQ1Rd6TBmsZNALrgmI10bdqorBkkMl+BM
VAkCzD3xPmJIvORiZD+7l9UmBFvu5Bs9YRpA14LiUo8/Ib9O6vKKvEDRTxQDNIcz
Gcwq3nhjfPYuwa5i2s7xjzR0QZUUPA8q2/VOnFowvNejFD1Yi0E2AlzdBl+JMgGw
sDaC7yGZa9RY30nIT0rBRM5UAiq1bHgLuAn+SswvsuMu/ciZlDHn0nRdeueb4BIM
uR9+8SdQjrOJMUSJZx+lm01whqzFHyPWto7Qw4+BJYVWVm5PoWJ5gGlODvLyHwwh
1r9a0v6Ze4YwyHRiP/THZk1pi141obPJ9C9jE7PLpapm1WliCDAj8gROiQVI44Ay
+kf5/7dW07+UiGsLRoeOs0SPnN5q1x85sOJyDVUzXhk2UhTzPxw7ev50O3FPSSE1
k7am9P0FDTIWM2Nfi2+hPXkvht5P9RRURZa317L8shPbVgmV8q4piEVHqacdO8mG
gMzVhwUX1DYtTI7Q8gqWZGn2k6pIUJFbReNCYzCjyvNki2T0jJgdbH/NmtTyDs9x
0bHAlYtmanyQfswgexxO8906ne4yc+dtiwu7DIqwuEjPXpEx8zIcnlalPT1QR58E
3lqZP1z6do3VAUydYXWYk2o/KqVABWXCYNASn7dc9vZcRQWbgxkGMaTX07AnOmEH
682uDibZ40e3JdGzp9U5s877D9r8VkpZpXBjirNvN/AFhHiVeFnNpwJdOJivzJgz
EX52JE6tNQlHxDW5gfoAao9j9gs5/srlJvEkwJaB0NykK3PXw4QwWfXcqEYjKc0X
EEn0JwgEWlQ47s5SD6On0EmsQsi0HUMfozlkvllSVacEDWt/fqB1XAyvEI8lU/gf
T1JwsssYtH7A40eoLGAeN9OqKXvASfXO5fRf6c4+pn8y39ZrplVnphItVPfTA+F3
5769WAPluxW/zLCmQUeTa+27ojTUxXzqS+HXotuin/QU1Nih644/ee2leKy7BoIY
rVfSayhZJTkMvQvTdGHDPmkiBhXKbLu92b8kYKbT/HiHPX4KjCBJZgYABp2Z0q1o
nKFpnjnDdD6dd/xy0VCybVGrR5i9AzPooTiEX0FIFry9KaUgF9ytO7dMA5/Ee9sx
mfLPpurGKyeKlOoxJ/91sNOfVWdt7wIPOUyLKnyUtap8f3weguH/rmyMvSCiPSq4
xsle71kAhtZi+k+vut+iCeoiDxRA97Qb8gF52+LT6+gIIVa7fM9Vuro7XIQFX632
8R0SktnagXPm0FoIX7+LtSiotVjZEqkbhf7Q025nNxEm5MIdUNLu8qktVBwc9TBP
0bcMIsKYzmf4HumoudbIPWzuQ+8YeLwBKPgQj7AalVdd8X0mtbY8cQp2K2biq9jf
bP4x8y8UH4S3TRXEsW1I0fjLFgiK4hcRLMSb00w5nkCVdwUxQQ0ewniGmMWgLlJx
NWXEs0PSZtUyr3OXLj1+WjENEEIRygVWF8gX2F+8S3JnDAr/GG1MwgUledK9In5l
tC7suDlXl1yp5gzYb7dQAqTzXpJqkNyFPtgz5EdfCtYnt5WAJ9MDktPQsGomlAMS
unYwhv5dWDmK7KO2G2pug4+ZeAzfe9Dzo2IAnSunDNzVq1OoHZiLKqOFZqUCN+R4
You0bQWm9QHE0JVuuBvQmgxVxD+bIUaFYv+te86GdGplRMnD0cXCqZKb5YJvWCRE
4sERSSNIaxHNc0oSDZUbWAhZ/m8voEMo5E9P1WDrVGYS+mErupRHTn0r8+DXe5PX
yvJKRlZ0Z7GMDp6wew1jZlauAFLQj5cp/uuAwSoLJlexdSnHSMdxMusecJCyROqY
0rcS0ehjq6sgx29bJr7Xsc3JLaxh9OuGxdi8Zu+5GjE5clVZVL25rmOyZuEaKPcM
NYJLXvvlYJq8uuger8VUe3zpmjg2mU02r1XhIiD6IT6WMWRz4S2wC8htZ5+UD1QH
RmNBs2WJTt5Dj1CzD+36HhBidprCtWHYWvTZsudSHewmUJ5OCSiQ8xCVxScJlBaU
kyaHEv76ZKaP/6V9+sj8R8QLQ9Q89JL+BzdwyXDbaxYV2YEMYCSKlybDg2Qdf/GI
DFLqzRU1pS7yzlBLWSTsowYFS1OxmbUaBwOHg7Plvtu75jQ+W3PMZegXC1a/TiOl
J8upQJL8WBreaoDuWcC5KnbSDuN6KmtOBADni1c/37nAc6mpw8GT0eSN3Z9ZRIYf
GzUlPvo8eOi4hcGS8wuGZyzhNXGOxJHRHzzteL/JNdjkExcc3B1BHohWyQH7wL4A
Nc1jh75KAZY/Ea+QbW8j3XsB1fniku8SN5wwCLq/Pc4CF3Meh6H7z7sCHYFiEVTK
WTsB3Dgt+9N99O7qj8t6Q0FshquEy0bglh0DC5oA8N14kmZ1bpdIUCISkwdGyDgJ
k7MGMBjsSjCSi4y7jI99eLhHmZdToxFcdxSzFGshe8gXCOh3xInfMw1zCkBPAk95
pymI/sD91pAqteWanByNVt7n9ww+txy7h8AJWhjepEr1xK3dccsJ/2t5M+//OQS5
gSjUYXQ4mQnyS9VO+Fky32J3BS7fFnzq/gd7PwiZ3JTuxFSiTGKMQSiO2bi+W7+D
RmTilBLCBkSGU01ZgZpbXRE0xqsZljz8X7Vfkm1R2Vm4/Jr6HoQs/etLGnU63a3t
O3WvBoeSQ+frJcmL535Co2wqXSK3e40ZaHfjpJzpKq/U32hnUAHVbSOEir6OVvEO
4f2FLf363EjGGre8AWMGk+o0XTh4Z8Sd4rLVyCNwca3A9LVkA8yTCwB3mYJCzt8X
O8BMtnD7b8ZAvL/cMIUWH1wBVIoRSDPqIn1UY91FIj8pgx085QI3z2+OxbSPAMd/
65R0Ev6cta1CywjtzkhGyVPC717n4oH6t9MHSe8cdw62aykyrTp86yKUUtvBMysF
no7UAdb2EAocXPJVsKxAUPuxqIL1gKA1mqnyyYLmD61r5zc6/mmwNT5w+XjNv2ZP
FefxKe23vsQTk40WqOAVfeT04qA1kRGokKxszgRs1GG+yIXkwzqdz85M1/PwNz4j
8b2s2X84jL2Q9yOdOX1y9DUH0P7r1ASqQIDO/ZBumGn2GzdJPvR0q4VnKAfsC3DD
k9BO62W4llf8lEpJZFyKPcIEcokJU1JNU8hVDwLu1tT9DsZ0yCRPqf9j1ficNR1O
F9IAgaSqCN9i7tPmg8UCS+/k8QkIdBiArcfsosAbLZXWJA6oRcFAH5CwtS3ThuRt
abyWE5Qx3OGBcY4Kzu9R2Fj4oRF19ZaBOrOF2YAmovF37b3G570uWLMJLhqo+2Vc
D/m74eP1BPEnp8dZmFvzHp5xEfWrEPshaGM/TthNa9ptg3Un8MphZWMTErj8QBUt
mDWWA5WxMbz2PmzWYVpBbWIb22C2bBBdCGQ/pCMBv1v38M2On08XwpKiD/AON1tg
sLbGhbCXb7Aclb7Pv1M1IveTasCld57As3gAGBfx/pd92F32aKEL/daE+LSJ/flT
3A5477/ZL9ugQ8X8r8EHSmg360lQ3aHvGX3Uv12caXWYiTopTm75xkuAaAFC+uHV
6Q9yjdctt6daWxPIpu7dzCO/PX/2gOh8J7SnbqzZpYu3dus9cvtEkAL+hzYcg4t8
2tTpcobg64jfC1OcymvMGVJV43ScTB3aEH+L9XIfO59DLIPhU1pdY8cegiw8MdRj
Vo9fa5WkhTJNCuXuNOMH0pbvpa0N7JKSNI773Px+tY9ojJiSMo9k5cePslzAwlp/
2lYM8VRybipI+71lbEjpjB8AnOPCs5lM6MkKdxGD1HmtwwKku0AVanEYFqCr8hbf
09wLnbEwWnJiYcVJznLkgaTIKS59WExKX5q4y1ulRBVYs/v7KvcKUV/U4YkUdqHS
4GV8wO2KJ2EJtVZqQXST2iBNJG2oCLipNu7Cr46+lRXziGsgRNXAkZU0QuSgB8Tg
NGS//MKB5OJCOoSGLQ2iKC4w5OaukLxk3hGN9Vn8a8X0NNhvHRsXTpKqnEhV35qW
Utrzg2QdVMThAwaetqSzkPo9B6DlilzDCJXDAMW9fO8LNvQGsWFRz5HXdllijjCQ
Ig2G99wqUczmhvCakXbRFYzvSM8ukcdoo2FKaM11yF8HR0jt5IXWhhLU1gKnlr/z
Z467t1hdvviOFgII0Rc2oZF0qk/c/0N/t3OfVa38VC0p6EvTC4sWj71lFBQcsGAC
ibP6BBb+JwNlef+VZeQfotkCYVwbz88DBbEi1Kid82ou9AdkwxJuFtZgFBodnpjz
Zw7ulcQebGkE3/2yr3XhT+2IYN0fst1YjIbDoLtxwYcC7qPx5m+XNhsOELgkvWKy
eUuQvh6pjnOtlxURpV3sZUVKTN5qYsMIO371a5TvMxWo5sby+MSoceHypz14WVVb
XzfhcnJV49UE+j+7H+JdzzB1F0+UTYV/4l1rbhOIQNGdp2I7XX4GdenIcjBD+byU
IfWGfsoMtwKNWg16q5h22VZcqXJyqEQ0B+fhXcWqWNRNd39AhciTWk820m+wEvzQ
4Y0vMTdHzyLGRR35JORcbLnEFgthdfPvexpeXOLi5ev+yxpWjf6WdcX9FFh+ixDk
tr52gYFZnytR+8g6MS4Q8RLtp9QEXXzKq4Q1Mmkr9PktgrYcge0aRI4TQkVY9zLF
QLDP7H6/CcSlcF8NPhWx7DocrVCweuDTCMDq5nCppW5Fo6fxa61plUctXBQAzaY8
+QyF5yaz2a+GqfQxleaOM04zwBsQme5Jgq9QIOnkgmbdCEF7NTemXZOtlmPtj2X1
jR7fRzzkXaRVuYHwC4L4kT/1XrnvpNPwmkWHY4Hm3TUyb7wl7cM8f2enxJ7AC1JB
ExXLiUkhOocwkJWufHV7ieMi2NXbCgnBZ23KJz7K/+dWf2+pAFDhk8YgwrZiz9Is
0dlnavFvRlhLeYnfZTF2lKCKfBYq7wbTYUBFJ3ct8tz8tlG9b0gP2zQR/sm5gazl
WU30uLYc80ZW532hGej/MqNBP0k870MiPGbvgGANocNtHZoWilcrghT5gOCczD4u
CjriB3NnseUPMAZq4eWw8wB0R0yXaCq1xujTiA9phXi27ajxl9y/S68IvmNXVlWV
Tl8cdctbYEQXguSZHCdrZkmkBAH6bNvaA+Si9Aq0LLfrgBMc7KjaRrjHlLBcoCv7
FAhwLvgiDZSeZGaMJaJvwUwOTxSyyCSiTUJoHexKvyn3Pp0RsBoPT1ovmLxjki7e
JTCaKDPmaaeVyPmPqRYG2Az7lrsbZE9Pb4mJ/q/VYxY5s/toSibJ/W4QVtkQKv11
sfexd1xOCc9gRgB0xUPOAP7845KxgaMF1cFxG/hxYh4vM8jXfg7NqfpLdxAS+38i
NslmLi2LvQwEM0CZtma+qb8FhCn6zR7WW0rdOxAGyXOxr5PQk9GAv4t/NCzRkWkh
E9xyJbZVnqpFcAjlcAoucQjRAtG2IYq86UhVZjL6LDHkYQvFtNhu8fCJNuSRuvyl
bCCEbxOX/mpCtf4bWVBdW9fqJPEDjgNbo0mS0xxZrRXj9fJxo70xAC1R6Vcpad5H
jYpt03+FNxQ7nqc1c50rnpHDr1kQRPvv1xcduVPyOxUkTDrR1BiwFpjt+x/ZpUIy
2OyfxWWXyfBxcOt88qIz9ea3Cr4WC+23Ye2lv65hW6Flskyt2Qx8CbLXXwcoqFW+
TcQD0z8WwVvBS+DHmnjHW4ao/visXFWwxgfwaoPjn28xEPa5cJ6nNp1vNPakjDSb
BdrIduCbkdQAwvqVdS+EGVZw9SdiU72P3066t4Pr9Do354qRAckNh3IkhM87a2JP
BUn/tq7JOyNp2H+e5bZKXSUkyO6L2TnFUhfLiQqDMDCyrs/LkOKUqYTD7leGtu2c
RptG5OF+771HjVyx6u2F5cIkdm5nOvvkSuMhHQrwE2P3WF4QdrrDenO6UKjUJgl4
7uFutbIXccXXt9OwMSRcmUh/fF5a/1c3cgRR3TWLiuwLkAeKWi/bJp3bEfZme0Cm
pCLJSgg8CM8/XartKeqVUz90pF6I/CxTMtzLwRZV+HHcTsUXkx65ooLt/Hyvp5BG
S2pf5lMjaMiuKTTC2VWefTQfFvxtZypjDcoNWfW9OvgedXZr90U9OcCtFh4x7o2W
Wbdr7gHL0cCJC/BoOQBpHwooByyo5QW+hvUw2J1NtisVvcwcmL40XcUcEpCmT18Z
vLN55MtxmzVekiNCQiHYXlNDpJwtCr2Be0CibG8YWCmz62bHUVE3Y6hncq9Oxxlc
ulN2NKGUtRPE3YUM/BslWiapSiKp70WPkfPKaLmRShYLFLUNG+kxwhUrTfdG7X3Q
4PXeCM/CUNIKNUAA4+ZZTZ2LzZcBtAOixNzsRAKzzZxvj5atkWAjphvR0TE7idKS
zJFphrmj3s1U/KmsA5YexqcvueiXo6i5YeYKMvhdfyI3J4cY6Z0afSuOvwDJ3zHT
R0cg0LbPtdM/YzT/x3EBRDtmekhtx6WNJtAdmdsjiwLaeJPC8QRiBVYo+9Jk6RPP
H1e1TvYjHN6478QUrhQBCrqoQtjoHBtKmUvL+6kvZ4RIsqsrvnBBl60Jq+m95y1k
wXlgY7vXcAJ4nsOPCWAScuyYTG4QfKX9kDxPFfrfjEoquPWE3+a6EBMdWbLVdBQJ
xR6SyL2Hog77PKZ2ou9J/cvOxFsF56n5JOyfAs+tTuns3qaKUShDT1hgvoa05I2l
h6HrODUPyg2mlZt8RCnXDAEnAAvlrKzeQ3x0OE+4HBCiUwVU2+hndePj3au7rgIX
UIdJvOPTsrrVPumxWbY5134buv7EtaXKP6AGP2YEM7B6Djozatj6URtqn8/3785e
uEvLPjJXaKTu1vSzp4Sz9RbP0yGCmAwhAP/YiHI8al3fzUaRRLahTQzfYb8eS4Mt
6oWLYHGfnXePTBasj0KuycZmXc1f09MHxc8eljs2slDnZ/KbvL/W74EbE8TAxq43
eeSHKmhNQTq3Uv5mJKFbC/WGWjvmeHphaOSLpHI5AVP6jLJEovonEb1F57zZCtNU
rVGWkNiBSA+3VZvUqWG/csswUrBa7ipQDSKdTeo/8X9tsIwJukcDNTPQbZi+O+ee
Qd2s9ODu5PDhHmsmLitWmAvlerA3kGaQnl+F3oBRTObY4yCFARvFxzqSFfPqfYiL
EUy0yAsXTo45wM3vsXvOmUhHgnWS07hcAYufdyobDOM+XgiFGntTwJOZ10ARCQ0b
ZUB/gVYorDkASq4VB09eNq67FGM9M0rwHuibjblvPR5Y5nAReRZs1VbomBURBT9i
LllTATi4F0PUKYU5ENY7eEBk9asWNg0IIfX1777bDfbO4vd2XIRZpxCgMLxa+Qpv
jNxWGpZvQXDcsSMxh5A3X4S3T47ITjnNzMzMp0p9nqfJUtcyg3Viz+7uTTVrBpIR
f6D8ecEnOg3VGKr7drGvMndTel9sAuQE0bQ89dSoh1Tz2R/36ldlfwwowXVkyHSd
4OKMOjMGAr1DYIt2y+EUP/0RHVU91xTJT2a3GKA5dypy4tyQyMrsUUzwYAnVG1w+
1vYevMUB83W7RTF4IzeirYdBA4jY2x9c71oA18rhHXtGp4CPK0I5b7zOq4T51nJk
lQipQ4MDXxJZNm0yaWsPWSJJwV42jTAePsAItPTbk+mpU6nbUuDCkESIcwwtOzue
VHqxJWz00KNJpkocIqITZhp8C2Li/XwEgqV6c8bOqRVWnH7s0rIhO3+NVxbY7ZDU
VOeQmz1X79dow6RcEqtBydzeqHGkkg01/8drrje15FlnRGdMegfZLLvpt48ooKE4
a4/okHr941V2/NF/vRH2vK2rdispJRbEVOlEKRFuTY7e4f1BZSrg6QLLMiXbDI4E
ZWwY9CRHuwZabt1dPGFcAjWBjuT/hoC7aW4qTUeo7r6+v5l0avRELOAB3sgvuTvt
RWMzS14GlHlTQgmqjLu4Mb/9IFWYbsciMr2779X4AwZSjkKnn9spCAh8H9A17z/7
3KS1w3WFMpjBcjxwE/QjnH1QIDZn6UOAEZZvMzIfA1OOLZGAI2AVVBIKNJjQMxSF
b3JZFBu6ozy1lae0/pxQ9AWivjVc7LBI4p+0LxXSNhi5z8oEK0Fi8U3RvhCROt89
HOXjMLVxB7i5zZczbhmyz/jn1BwOk6I45ELLedp2Oxx3NfEMDx1GcSQpKsohuYwK
a4KZe6yNAogEDQfY3vn2TGUYmvDIeJpM19p1k+KPITHhbL/4yMFOm6aL+invNKld
Wnmfo+CqaiAtDISpMyzb06QjbJq52mlKHZmkPA4D5ERQG7kSqP47QM/DOcIvd1/B
oZXfRjG6Tx5ZWnNAlbuzVQET/TUdopOMOq2wFGPlM7v1LYBc4UtfUYkjqy7p3cOx
Y9Lv+cdm9mqmevZMnN81xMRqvIM72aTUV+tcLmHWYsqNPFkCRhUAFbHk69r+4fKl
uDfnfbl9wfIAKub6CPayaLbjIlGvh0Q7w2H5QDjkKo9uoo+JWZfMBIhBHroau18Z
qxKyBvvVer/TAB5eL6cs65CPYD91TcQ4ZCyLiRjYlgBcJitFL3lhQaZ2koINwZWI
eJeV9AGaj6FLonCbPNi7FVlX54yL/JDTJ9DMIxHS4bkRDhz5SlMY1MsYp3/rUBsN
KiDGZoyx8cORkYtM20LsPXiAnBfRUqbKDCv/fT/l2e7TtHDAhw2NbaWh3RUKgdOC
Y6OqvgM82elZk0hNKTbQCQok8f2VWeKU9r/pm1uU1jBADqndSBQnC0ySqbpSzUsg
wDWGEq1ulv3J8ktmT5QxW4cILO1ZANgCCQq6xFfiEe6PPvUsS+CzILvyfijkd8jt
xj/WR4/bxji5Lneclk0gKzLSE1KY6Ua86QV30IXDzhe41c+z7ydcqWUjUqAxMDIf
7W+Ni7r25jpoBJewvPUcTFmOxs6RoZkLvil0//Ox6Al3mfqYuWT766oT3Np4fsSy
SS3g/6QOfTlarSgdie9HsnAjVNbaV3P82V/4IO7Q8hwFj2Sc6L+bWQh7NgBaXEKH
KdXqmOV3iqXJLGvdeZgL0YHMiVUnR0LirvcL1k6C2RmoggOauC0uSFsugwSrKESQ
l8UmTeGWleGgrYCEXlXHynpaUxQzNjAez0EbB05g5LldYO/+jQoF2bcCfTydFjE5
8/oMw8lVIMTPtB5DEQ4bPG3sTvxGlveMym3LlcjYpraYKRL2BD5kyNPW4ipA8Nyw
U0ZXH+DiwJn8SB8YZ3XbKXXL8ROloPDyQIvRDzETYAmHj9SKuI06l6Yas9CZJ49J
K6Fj6fw3k/O6wNEnIRA3fJDlnZT/2zNJk6Pr++j8gL++QQyNQWr413l7lECadGva
p6l9t//s0dk+yHfEw/3i4Sc7wLu9Oe8UtAUktLlEp33XWlf02CHCRnzOaS56+d/k
wAZk/Ed48ZD2OOwjqa3gsEcWusXMl038Disu3HXR5uupZ9av6hIZQRPCtkwUzLMz
bZYLnTV4fjWaE/ntboNmTvjRIlIK4rijBp+pkfjvyETL6+L2cHS/r3iemcklgiFF
v/4HCtu9/1A8Z1cg3JGeqoa9Rmvho7+6aFIJw6ld7RflbDsIbgJTSrgdHLPuuWRb
Y4qX9RMy6pr9Y+IOx6K4glNA2L7I5B4MK/Fyx8+bXir56rRfOVU+rnHobeX8myO4
yXox2XeaA9aKXVqdncTw58cQZK/kJo1y6s0igE+8Wd5j18w1SRwkEfBhqK1m3oFg
fAUpj0YaOIo1EUbYk4XR2wzmYujv8VLJLJp7zNa9Hld7YdFfKx8IyNXswyY9a5ht
ngskDNhABujaCecZpSoi0A5udmsrKuDRmChcJl2RbagZsWJ20rnl9wa2K2Z/Kib5
dXcKwRv7EqvzPDRUoOOSbOfD0ZhFGdL2ssaMl4K2xhsf1HndO8+YG74HAzz+E65j
oNSQPArHrDYQjanxF82SE2c7mQGI9o4Z2Un1xBZ3LJFyLW3+sP5USrjz6OXkNTqn
UHb8aKcvr4hwJDFwSHgL/8zbK1L7i/GcBKyjYAJenw7wcw2iY9kcXPlZJ/LRUWMB
1iUNwcbJOE2QDvlCFYo5jMbaSgbCS9xOf+pKzxVSgndevyKIzu/hqLVYCpX4za8x
pyd6IFsDVUevQ+afkw8LyXM/2cuQ2X9iRBembWT9CysawxCYWD9UMTMV1OasRqJJ
BHkWKDKxT4sFKyvzIg/4lT+yV3DvCMY010lTxwHjFqHNYHrKxGoxupv4c6sXj/Yv
37ZmvNfEKXU7NRHxKutoSX77VkBrZysz2BonD19wE9ydcF3KfAj6zQTF5pjdrgCm
Y0/VWDd0YY70SemDywos9sR4ZJ/q1yPIFp22bB4CYt+YFtFMWEe6lhPtzWgUlVR5
324RFdMlDrR8CeThasrxokcmrPUwu1KGmZ1LIJrQ4EQ6iFC/y/8Byip50om3QiG5
9+2n0inJhk+5TeNXH2DIgG8659kkXRYtIxuLyyphZmcVAgfmfykhHYXNCCZy2azv
WHajOKrW1FVc9RS7H32MGhc9ukgAQKRYgcRvwo8x37IXuNBGp0IM6dGCtKLLARDD
a7uVNghBl8T1PW+ga2AAJi6cI9U+P8wpKIePPSE5RZKgihQCXCP9vhRGlyJpQ7Oc
r9Fh7wvFjJXlvZjUHVnF9eiKWhaPW/SFItHcAdhQxLQxBBxHEuR/MR2482wI/dwM
RFz42KEeqxEhpNdYYWYgcAsIznk+ZOdFEJIbaC84WENQX/NdH4s0k5cWsLJxboC6
p0MdLGqAgVocFeCiRwlxdDFqyzS+twjjx2HxBdx6z+4nqYvUC+Mn+taJ33qsr6Hz
539M9gOrfJLEHaEm55UE38A7+cXSd4qtTmhWFI6s43q2xMtQVVbkT1AUawzKe/Hg
LEh0EexoDatDn8ExH27vZ3wFCirt6/tYXMYJKYT+ewutTuTVtweRMhUbbI+DvbuV
rtGDz4yyxQVBIj253ML/odNjLY2Scc5MPG7rQ5cv5rcTV+j8AOpf8LJEeTwB8kEl
v/AT08H7J+Fjg5FvPzF//3E8Y/umS6apyENYxt9BHx/ilo8zY6JiG0C43Kdnzfce
Qtr2+jtsvXA3VkX4AetFr3JDUzMIAHqKeSkr9DJZpLtzIJrqdPgLOXOKpx/KKpem
meySOolh+wydIQdJtRhd1DFy+4mkpuW8MpUOvnUZn56+ceOI9Rlb09WxsPc1ISkP
ZXWeqqCMbJjTaC2JK0B4Nx7Utq1zXmSTt9Mm/3YZ6cAOAx9OaebyBjM5TgkmRKS+
s4xBHlXrqK8OYARcwVZkMIRnUdt0I+DfALIl7G+aD1bK3oVG3ccF0jRtbI9tkUDl
svskhh4zLO6zS3pmTxDSKV7Zdo5ts1qbTBZNdHr+RH3J64xm/q2p8PhX2lmywAXo
MDcQAWLvWpueTfMRLNw2qEua5pi4hzqMCMKf1I6+ScLwrS0PFYoRtVUqBfEAD8yG
1tItV1FU0Jq45KK2MtyJO7sczPcTax0FIMuiMrewdYosWZwXWd11s1CBb4gAOkFA
TqE2Y7a2NXvraJj29HQMzQpMfYJbE5b1M8Fdhfez7O61vkgIi+XvKmaAe9Ym9vVl
SXCMmU/MP4GXEfNTkaNvCZ/8EEcbVr3LRsfAGd4yJCm3r4gmxtoBaBsVO2tc93Pb
vpI9wJ0NAkYPvk6kVJGdnvlYsdlIB8lapD16K+DVdBljTZF6hC/Vk2cwVmgxhBVJ
C/FU3syLLcO3JS9V+rMC5gV9p+CQSg7CkPEoXFWNkvTYxcYRO6EM6qog6fzI4qGW
FPvHuC+ZfmGJkhYzjJJORQoafFTucgp+xQnVfUkiovP/kKlX2q8Sdo/GbGUQTNxu
qR078qOgkhT3FeVYU4yKcQ0GWpzLzTGHbyctGDrPLEl4p2RF6VX0TGtnNuQCUj6e
r4VXpzTBO/s4wwbGCmO6FyfxiTuAImZZ08tOrDIxS3ATM7FC2vSgwp7XRzH4j1M6
eysIrfEAMB3XGzuniBGYqbksCMgxXPx1Q+y1j48mH6L0UFS4ko/0wXgDrRgTMWbz
VQ79D70MM+LIvf70aZZ7ufy3WWIgCFyJSLTsCLYH4ARwVEtYuo9bNjNZ1DA7Xfxa
2oCI00MT3j0Zqnj6gMOZjJqmWJ7/650i8o6B8J0+6IpDPdo2wffseWRH6I/quA3x
LLuMcmDWB4i8uInLLL8RTIiYKJurwXMnQ4NVeEH2yU8rGc2/sa8ZwM0MekJG7RQy
3W1GR4gcPU0+ot42PRxWcPIdayZekGl8l+nR/1VIc/kEsayl/mBqVBdS/lNIzYKa
SZNjQcnKpAdQpgz6EsXNF8R/vqxmNfs4HGsnV/tYvlvjzKJu7K8UhQq+MdhZScaw
Q3VZMsgiqRhcA9uisOveZ/1nUQCP/1eFtOrgEdK6P//E//6RxgXL/xjVPqJgZw+n
c5hZD7SHoVca/JGueZdUPArTFUqSqeCssEkoO/Yn0Qw0Kj/y0G2N66CCJMhQHnI7
+W9aVSjMhENZlOY2GY0wkHmfe+BNbxe0ueTnZoQ3YeRki4E0iFqOfAA29/ITva0G
8dqbpudAHaPN1OzxQb6ufbgS6T5zAc70fzT8InpmlHQMBHdqN7/LQHk4alhL6r1C
tJsyOej5DBS1+Q4WL1AhevwrDg/4Y3VGnNTA01X7FvCj2wqmYhv6YFAV7wVhMscw
Yv6HNSs/2gYLBTRDLTa1G3kJ1n/51cM9Htldh/lrnTd47wSZickNRS9XahC/94tR
H7Kw/pvdTJ9ZszlFCDywcU/adEtG07MreK/rGYD8LzruzRhIXHCWNB94z7N3KG6C
Gugxn2Fnbpx5PmqUlY3bU78PqmOjOyqM+u2N+XYZDs9Y1+y6FIWQKkZg1FeObkGs
F4SuYHPjWRqd0NQX2Lzljb2GMzf5XTJshWAWYMczyxSpTG9/3tFpBALKgHKUcsgf
at+xGt5/T0hJUSf/Ju0CuGsARCohRciQCAXsck8tT88V9zgTqXYhh1n1AKiKe/5/
5itGCnBnn3fWkKi+3c/7cWOfOwy/QSK7cgYntvDowawH4vlN2yrYo17imojryuXI
VCDXuwqEK5L0NvQJxrco2usrt7CFJzGMcn9GPkY9H/yIamySzsuCUeJaqPP7gWLv
czNrc4yjpAWi5myea0y/82dsP8KZyXZbn+nJcfCXa0l6JEb0PPKuTEmUD7iEQjlF
2CkZ2pnhEMAVyz9Dpx60gqB8bPaALa3RTc2na3rLPRZB6qvTgK2MbNnxWrWUG/T0
ZeEJH3jic2zlJxjo4cOkbmgWEkzpDEIaZOjDxXQBRtZ5U8vZjoTPzHPTLthSpizE
oL1qY5eWuur9OJz8K/qdSwMboZ7Zj5prFdxre+H8WSO8lvQZkcOmhmcy8pkPIbGx
QBSOMDTE+U7DhA8nAuChfl3pYo8YnFxHraPku5l0rKSr7V100tIAGw/+RzNXMrMk
4T4fFHMW5KlZId9/p/NmUq60rAc32m3hHTzU6sds44Y2YpEH1uxlITDUogrmwWV+
zw91LTMFCX13b+5LNVrM30Xi4r4kGB2Csi2mcg8O9sMMlVe/ifIaHlX5SmyD9SmH
bcEZfzx7VwrIFaxcmekYJgfwmbPgcs5dPCEyHXLx3+raH/85C3OT7FijUh9wCDIE
qOk/AyZInoHqXFlGsfn456za/4hcj5rEUbCtsyVQmx8EWIocYjzDsfFeACUHmMEH
rNK44MWobH0bgHk8h2L/hT6U4DH5zeAZ9DUruQO7tJv6FN9q8zB5soHH/oWCU05m
rwmk+kuX7VmjieXf7htH9gG1xg/C6Npr7rpZ0mPaMGndi+q7D2oK6Z41YUe8E5d1
c3ieWkSPXFLX0pWVIdgjBE7zaNoOAiYuQ0PEnlFwX7ECz3Vz3y9QZP3mG/U2KX8Z
PO6gBWjxTo7DcU8yInWkmmrQ7LWo1OmkaQv+tUTCKa29PPL5IE+nowkXkwYzHfbC
QouQqpHvnD+OWJhhKI5RJPGKfIkkwZg+QRdPUXHuuIgk1WvacsKOnyOYTgs5zlz0
+4CDbdd87lsQG0T+ckGDvbuPBW6JZabAWQlOecuRZiUpdD5fUbHaJzCFpZzb+5Zd
WdWvP4TiyU22l7f/3Si6bQFObJN/zlX8v2OVuwb43YyEUOqMQcyhwIbBgPzev8Tl
OyduTu6dJivwhA2dAqq2IYjxak53LD3R7b/iTZ+KmqkIEYxi/m8ZhQzvVrPDGy14
KR8irBMMH6/Dbit/X0zjSRI/+0q2SiEfTiDDHsVFBsyC5FdrOILY3JfxfTNYEJPd
eh3sYJXirUzA5fhw7Vox1xyfohRqc6TnuEyKznQqVBrGxJNgZUKN04SjOGrRRJzI
D4tLmLttjyukDhDA5H48tt+Q+aNDjQqryMythsb1a1sZdt8egbUwdmIuH+4fA+63
p2VvavqiCauXffZEjC0gt3mbcy40Xo30kuQzrG+kSvYKCTd9RVB42h5r1Hrw+wPb
BedNMFQp+51BSNHT4JXLpn1yxZZ0CO+x2LqnNTPR3LBxCe/08/a+NaD902X8d80b
LeVgBij4FyNiQeE/gF2ANx3CnXzBDyIJHcjgfY2nqmdZ0SSGOq2AgtJeOFq99KPK
BTEFAJw/LPLBw4MRBV2mRs53FJkXh45TU0hLsg7axDX5f7iiZKq0AkjJrn9R0Poj
t6GnN2ow3CBLb2lV0uf96PaRjHXZ7xJgAvQIEZJipFFwPDvWrwo8W+1NXOTvHr/Q
POHRM3gIwkVVtO+Se0+9diTSgxGat63Aa5ynmBdWtw35Zp8/00VY7nniW76rUt1v
LO0O4+HLZdBpsUpdgv1V10tLyBaVZtyOvowOvrBkjR3DS7+ktR9/eVC3N0CVxlJg
T3xr3pRy2bqVm//T0ouoQi5e1GlnQc9y4ZCcq218gEf1p8tEhUGgTYwjSeOaty+u
7Xfvj+CD89oTbAn1wfo6/ziZZZnWE8KZfRBXqIYmDKXacZ7lptstjoDM9+QCHonz
QKgSqDR8n6nJQLxCI4r0wKAylXTXULQQ0FV0bN013Zr9eAGbo5WbB1bD/p8/irra
iB+pEfaU9TXrrspWulFMcueIhIaGH4RVOkzXKiK6PyOG6sg2Oljxuast7m86XMaw
+U8RdZL8r46lQZQEf0UhgRA9zHn5k9TwZB6VAEeu3yDGziJcL7zUnngxaSyx8zpa
ttRNMr5Bn+Qq5H1sKHNgckXgC22BOJcx6Nsjy9UoaB9xc85YaE384xb+QG2Utj8D
KRy3e8lxsG3prmQqoisiEIyvdJXUjwRK9cdY1OA6aDpcZY5j18pl5De1sFcdmrEx
Ay61CWuSjaa0g7EWV+otp4hrhNpYbLwAu614eL+cff0e+br70jdsfaTm8sE5itgf
vASTU4TRzSRuprqtt+XJetu/BXxNHlxPFhhKkbhtD9D4f4tfQ9B778F4a7dGPnzh
SoMUYIZcwj6GQKsrb/g8Q+m0mD6L9Ri1h1S9ACTpdTn8jcI2Dj6tTpu0kzXTaKTg
Uvwd702JbOMPB6/CtMeR4pspk905KoRx2AQ6/0laTOoRR3flFbcHs4QUng8Q0RNj
InxwTX6qOOcwmiw25qAbzxyHDOk7g/HrgTGj/tUMNbrHOL8Gg3H5FCOI2/sbzzFu
34YCRFcuWd5Dc9z9gpC3taQy54h5tvn/olT9k7UnzLsoslCJ6WQhqD/JHf92EmNr
j5dGZ6ZYi4eQtbSQkIJVlLLMQzxfVeC/yvsxyBRy1t93k3TEbzJkJ6Ut7SDPIjHO
9WjGxIoVycrVL6xfTJhU25PozoifOyyPErVGNSbDY3nOBZal2bSltnhvGlqoA2CC
3QUm4urg5kRIOioZFevTaN+NOE1Lgk0CsiGxWkh+132DWeUinGGGgvGFiIhN/I1X
Tb0Zuv2/7sUe2D64mMdFEbL1JJy33beuYkBUnLsCgtf0g3vXFX4cczINx00GviuJ
PgcHkTBIouZyAtdpBVn/Z37gwzqYk9rDZiNMqnBEdmyLA6QHiqWcNukTp3KKwa4k
479Ccx4V+IRJZ69SxxzR/zOR3DeY0sO8ldiNhrRPzgc+c7Nk+qnR6Fts1mP4adyW
XZiGJDh3jsd9CgR5+7C9ykL0OIVR0h4t7+lkUnno1/5vEPyVYATqZ7exL+JgJgFK
ZIKDWhM6McaPlFRCFslXSAPANMBYsXgVHHX0Tu7LC/E5Smrtv0K+ZsIhsob3PtE/
Q29sNaeUUsRtC0q90eiJ1bjRatNcxUHq5zdIy+/XPKDlVnrt8EvnXvlIIPpHptiq
NJBDWiTF4cLBbjWht7bwFQnCJ9osppRk9H9sNWD7g97FbpexlOBFU69j1IOH8R5P
iCP3YDNM24nP/Omgjk5dH97WLhCjoBP5tqUfh7haErUyKb51/EIkI8uRttaLQOdD
NZD58kQ3b4yMg+dZmJ2NZ4XZr52M6Dqkr5auWu09Cqfv/1FR66aTDszq+6kl0h4+
68OUDIBZuNidtAjd5RGyAGsiDQTN9DOQWkYvIYlSecgq0a9Rm+76hzFhyZ3I6xhG
0hoc9aGeJB1nURgWHCRgadGa4QCgIbOaWtAyEiA6u5+4ZqUWhihFu1rrfN71FBb7
0hq1XUmzGs+OCSucrn23OlGwnvaQglUHfGIyzBhlare9+hpv34zDdGEpjAaJ0YrN
3xFZudS1S3Q5KFmkP9zBWwH7o1cJlO4ZYa76R1YOMerAaEkiCKexCuS2lkzK9wkc
zdL4KmhWi6K3c+aQGRSr77N/7uNPmYRRy61ugfVfOrBKnbN2R300QOgxheQG++Jb
W/6kwhl2IHi21PTCdx9813ugtit3On//OdkVFzzO+CKCtfM/f8FvET/wkQmTm0cA
3n02TPYEwum9UOfyiRRe30gRDUnrtaT1MLJPFHQqh4X7KjrMeHSemysBhpZS3vOn
Vacu5XmY5whzeClNxgJCAaGpNMcF0bkyBMPhfI61bHH8XIyFdnWzOHqYc+c9Quzh
5po4ZPbUHm3lG25vCqK/lmX4KTWWCmM4tQLPfMwN3L3MBj8+uM0dEwHIdtZu/pDv
2/3BVTOXK3XXLfvRGmGAvKTjV6RbVAprPCyQpl5rxwjDYp+B96ZEu8m1IjnmQi+w
p1GkzdTZmylCbwCV8bXiV9+yfVh5qW+qgobZA4TzSk9HW4vI7w7gqEt4nUX0LVqo
BtAtT6rnC/yL8rC3RumUDLqWmyuRof91EBaTwlORg72U77/HpV25kPSDEcwZ7Eqv
DX/Muyc8tLtg5lWkJF/QpMSbyWuVXT06A6Ud4bkOIHbOyLkysDlCqsMKIfu4+OpQ
nkeq36qIOPpxGlrDRSaRMjvIyjJVGl+eQv3iLKMX5p8ft41n9bKQzVSQ8p3UENmU
KmlJggdjL+Jve6PY3PUsk0Exqa+Ru2uEQFhZvpWnNIi2QgIAosZrNKON8Ao62b2J
dNFLcMh9rI7IyCCr9+my6ZVdMsG8VVOcC9ZpuvlSm9TdzDpREVChPYSalVx+3wWZ
y7pE2vpLAWPsXQvPtDzlx1lb5jLtzb/TW1WM1jTjrdRlVcFDRvEK7KimJi3C1rtv
Y1gE2dy+9gK3Hudsyb1/ZOm/W86UYbgyaXQ6nrbP/uFSzo/VpizGp7jEjpq0A+c2
dZi1eT8vWBfTZINReBl+EcHXJlLghPjI9gUeBxG7VdYpvtoYqvNzXrYw640uhOLR
Bl3IQMg42uMA6+I9zYLH16J3P0sCInwpRQtA0dB/7EWYYZrJ+Grw6AncpAEKHZy3
zBQoMWKkbgRE8OfxzhcKdEqCWEM8oa1bQNMXP7NJjQaD/33d4rVDFhHNS6FdUN1w
g6QVQVuhb5v9QlSCnqF8bTz2fMbgcV+SNtahc67hqEfRtYfl5RV4CpRsmyaufWk3
zvrHXHGT3MXt8QQJ1mxIrarXVkJyDDbdJV9nSferl4uQ9M37AjDlSPGDdwGTrVa2
6mdLCQEl6FO+XCcLH0zxlLRVRDO32lwpdI9v7+mb6YHB8gsTxr28dHE2efuWqn8G
CCC06JvumEJdeXvt0kjiF6CH8StA96V3U3z+kwKeQu2gmL2LxT8RxWxjnq6T1sjN
xSp8wEhiAnpNNhfDyseWdTxtWaQKz3T99K2l6Q7jMvJjQlBfORQ+dmjpw1LNxEbg
N0AZwmwJcU3h4Ln12gzn7pNcvP/CzheMEHhw/SyaEjVFX9euT5R9mw8leYppp7z6
9x0pOHrAk7HNuLnGFnAA7motz1MH7WrNc+PB3tpyLnOfNRP9pVXTOh3LVBvUo1tE
dohsdT4mr/lKc5UqLFHqjtUUxqk3nBjSAgTygqdyZYZU4CVO1u/NkVWwNPnuYHMO
6p6uGpNlDfWp28PQGze9sCit1tr6gLQUDun+FlJJ85iYQaMFwzy8HzBJ7ioqZxtf
t9P2melo43BDHgdnJDx+qC5qJId4nxNbXCipWZYankvsh2YLqw5PXkl4CwkTk9nl
qhrHRBiX7t/n73pyMa8Uq5QIKoLcseZuXqC2apd6tWbWpf3s0nBw1Ypo69P145gp
9x+LbYd2YjUDE+sS9iSTB2wbqTdR3NuT3cVNmZzHNMtuQcFIUdPyWHtVLKWWm7fS
gwphM5bmuwJwPIWvCEUuU6+7NIp9IgymqwwXqoDN9inlA4+3dbBpzW6aGogRngFg
AIy4vzwnqH+PXt6J1ic7IpiEyw3+Yc/O+MoCTaDO2BAyFfJWDfHY/jyn96SkgE0S
2H985R5uiHMFKsML7WqKuWqOcHsuuJPMLmzUGSf0zeevIhDx9nnbTPbRBig9sDy/
vRSjnPmMEK8IVyCRWf7FGsvkv0QH5AupNuNZ62WJK7P/KweMRvuWz4nzY+8cLsuM
Yjmbkq6X3JVp6EUrgxb+dEMc/6YhqbGiAiZcn/GKiH4q5dkrJhuAjiy2fZheVIk8
+3y6BV5L+dsoXh1Yp57rA+0R8hK12nwLFPKpoP3HlL4fiZOZsdFHpthcpu9dVL69
elKkzoeN/i9fgyyyOwMezP0zmUTkS96i2we2P7acp6dv8KDcUro6+ktIg750FWkP
2Q8j+GGsVqbqrTx/FYBnlmhml2dNtHqeor8cbRhXT43Ye/iU5F2aUNw8DpUzL2Vn
m8l40tkV2F5fb0dakKj2nEXEyhkQyi0ax2r9raQ+KXyIEPxLRvR/oV3Jn7HocHLM
1ufBiKei4YEhL86E9fshhOMHMS8kk5+4KAmmMtVDXdB5WXCuLIfi2ApI4v9florl
43cb98vXGCvWASqKo8ZhSLV9gx0t5NPkJyGdqaN2fvNXU1khH7lhVJYaEgDp8mm+
gICS98OkKA1TGLKsMmPUvIdWVJNAbeBhjMiyCmtFvl0qgx5SoDqfsoAtO4b+AEih
162w/xR7Eecz2YHU5lljePBxKBwKScpsRf3L8BNAdQU9TBra0PueXAbPrG8xPNN2
Gv6a8OORxEIHjQlsRityTfGYBSka5KWI7o2tIv2aVDCbwMHRUuUX5uLYpAUTNKDo
8W3IYEwfq9wjH4RnbeBoo8aMup2pbL+1CQl0rdIZ1U1aWYpM6RvjZIN/8/nJL12H
/AqobNDpPEY1jetqFrckUKlOgoBwhuoDccB1VvU/yjy/Owgt3YjXdSoJlsWOkOVt
ugP2p1EmVmpkEKfj12NKVa4HqvxXWxVq7hIP4SotvS48qW4HCLsSO/vd7emgSr5J
CfizzkMntm0kA3AF1Mh2SkajXk6hg83bH8IbE6YNJZtnpAIQzVcdYJL/QkzpGUxq
agObpcMlwVq0sNTg/1Mdu4z1ihi3Ruk5TDJC5mf6BwKzwX/mdhqzjsIt96uIu4gV
s1rC6nH5qL4Nl5rxLCi9JYpYfa8F0qvUx2KW5atiJymO0PZoHwv8QD2dmLWhORw8
aUUu3wDj/nU5iWXZIwOUXYY7udK7fpZYUqDJu22hZZWmNO4rMM00CGjgRJ5ASsa4
URh4sNoCfNIAkv4GUAFBuzB4Xhvy2DL7Xc1tZF2KHc2BtjjDy7/z4Q8rNAKU/vR2
QRB3Y9u4TL2IzYCYCyvAqG4GveqkP83+e+mQDi0JSCaqSGxl9azG7zYpf99oqcXC
BeXToEYorZPo6Nr1U2cjG7IexbeC4Ttyjph4S1F9HsPBUFq8f6jzhyutG3RFhFdZ
Gsug6U6IpqF339fUfI/OYqiX4S/f20q3zIj+0VggYhPgMgRvLyXZMpVOtfYrZs66
6vfwMXXW8k+dKUMT82GXQrtjnx1Uwqtr2880auoy+aO7dx4TILuQrnP45kyKk4Ty
Tpeqcl33Nn6Pf2vNQPK/xRA5KEyfOkLABJmr8cYsHfvntkIS0rCKbsiPeqq8t4E9
RUdTEWBO+Y7mhi+oUaz94bjwmxlUvtrqAtWv/ifM48b9hINOLazEGYZLpjbhkYsC
4z7Gd3cgZbwG7oRBb5lXc/+ABonGRyQ0vdqi8uDjFsYtGpPACf9RNhQ+Vhm2oCmX
IgbcWYz7YFvLaeCmCc1TCTQP6W11dgHHavA1EjNnFpBWdjkLuVB/hzyNY/UVpIbg
1ctUYXGFMFBfkYzmRcSCrzyf+Lx68ZwY91cC9G9RpHxD4BBl623oPJOmz4Cgx8Yr
85Qz6gdYOaYUXrgQxQ3+PzyIdLCxmJ3pC3NzPA3Fq8BMIbbyJ+Pb4Mw3ZtJ9Gk+t
U8R0Yu6DXq4XnDgDKHl9n4mMAnzM64S1i0g9TlbSssyVqpNAZOJ9ABPdPWj332Vh
xn4yimBsd0dn1CfFSn3lPo8mfId7uDPR+dM1Fh6i2Qov62opB9vKbwu2QND8bhhQ
LbhDyhvAq7hwnXXh/1BREvZDzsUfO7/RTqsGePVMAgfMkWsIb7/nIfJRQo4rhvCF
+4Jy33k5EOtr1HsFAI+gzsrJN/WOusYNdArpXBNZFClHnUJz4H4Dt5y0O+SlW8wN
G8g7P8NzSOiVs6Wj8DVNNKSwT8Qt3O2ZngrcB8V/Lz2FiotvBdyDEH3f5mESVRA3
CgXfp+6Fdy6E8mV4V0GIsGcLZJXYurTpGV6B9SxXA2iIFjXvfBxUim/VTXWhFDgx
XBkChuCEu7vls3CYsEBH5NMcKCYaLEKCq3OUAcgzdsmVKtVlGEYFp7xh4ZwoA0KF
zXR9O21ESi9qfPKBREJfAU9fFqDtoJ21toHWDxWsa4V8RPN+6uIepBD4hIkknUcm
PLX7Kqy0N2yi+oKb+9Ig9w/5hYzXT9gYHscqXzQiarwmvz5EAvB3HjEdEpaBTDDN
svL0vRT9k22hTpKC+0jWhKPY40CEwLHpr87TDuHze6hC49TYdWymuDE6CTCukgk6
M3gm9+qOZYMm4U/Q5HyaFDHvs9v8M6a+rpXfI5eKFXI91w7IBrTmUyrNz6/wXnVw
fPn5hExVDzXEW42Z3dILhfnXxiV8dk21z/o5YblKT3gxO3KN6udG96qc4p8Yd1GN
D7ZfTfM3+3jajlqhsFLr2Za5m71F8KFpOLbKvyvAS2fnGu1iY5y+LHrBLmwBXh7m
RTYBicuKnMdtPBSa4UV9KVQBQczj8eK1gTI5jT/atWDhHE0tVKZCT4VSBjZoT3Sb
uUOK2cHiinTpYk0xy5BdlpyFUBZlQBAPhGJ/s+xasCdV3pZ2xveM6p9ukrch6EBY
03pXswCR/VAlvZM3mMxcCBmbKD5b7kQGQqgxxr8muFHF7u+j0DjuMe5S+/Iq07bO
P2XfztcGO5tHpdzcHnZNFsnHtyiS6zilNxyLKhv6WB4by5INhSyCNfnjvjR6egR1
2ShQRHsE/rk1Uspq6bpSV+eug2wMuqdNGQY1f/iOcIBZOtLJf0vIdsbdb2SuRayo
DrlgMM/wYH+clq+tTMYc53wKJs2vKFXYfQLUWIlj7OnidPcz2jrhgFa5+E1Spjm3
h3nSK1fXnIuxQ2rSMKCNhy7nABjqm0CqmK1gUiXzh5PmUsATdH25Jl9StlpOMB4F
Nvc7VdnAF0CrkCh4zoO1VjlhVJa3GUVuyn3tHHJOB1BBM75eeOo/nXtEe1Ru03OO
8s3LNYDFVwVRTaNPfEZ8jRyEZQIRVkvHGb9J+oS/QHcpFuoXbtvLUPM+TM6KQ5G+
I8YpXavlfJO5OVH10i1ZZsbGdH+d0hS12Myt3tUt05JwipvxtPrx+Ac2MXqK96Q5
ef3G5ko1QyGL9SlP9oKyPJlpVWj+6c/pCjWEreS5WbQNr02VRK29moauD3Iib0RY
gAiIY0akfv+alXoxE9nybUw0lpCdxDAnnfpYPwvSm9+kGTeRDkHr+9ywo30bJgHA
wsgq9ZvALaKmPtT5NJXkuHJ1KGzU8V6j1gUiWIYkai0P/YtZN98lvwv8iXk7FO7s
jTDx66dj6CQl8YUYb9ta3WnOw4uHGdBNxvs+k+LMXy8x+oXUPszgXPI23puE2SrE
36FJ0hMV9uaRiZh3u9e9TA9ER+JFp1WKGHI9tuyX/IBIDbZwfw//JZYfIeLoTGX8
rlla3L/WP35FVBAdUGIhGCL2MX/LXJZP7fhzDZ+N+PG791J9guZpuQQE0POfAmK2
7zvE9LQFu2hkp4zW7PyXdV1QeAJYXs2+6tKT7dyROfJlqdZA65dT2zExn1a2xrWJ
baOxHKO+UPOsktj1wvmjp6jZc/RrYYT26F1OkpmBn1G7gTWVpi/d9RNQfeIVWdf0
f0ynlslDovP3b6xIo1t1xAv1KUzkTgUt6t90Lh80mUHPPKOCZyF6TiwJt+fXJ06B
KD4k3jmQ0eHLcL8Zh0ZXwXYYElM1Mr9BD1y3Pxx/T7JpxWIThtZj7dul37w8JNPE
Vv4Y/13m/5MCVOYkUIdLhluzLdwzgwu+wcl5hnY/Q4YH154mz3169fToXiIzGPzC
aH6gf5+7rO42fND26aVBrwyYNPrV6LEKGafxCQB2u8qSWhCvTT5VNFUKerKid1hm
kVlhAt3kiFngq4bnE8xKfV0vKgwMEcsA919t7vftg1+zFHP+SibBFO/DQKI9nSz7
xbCArdaVVYQgAU52OYD/JOPQqQBBf7D9asGKEYpKvyvhoQrrqPX8cnSku4j0klA3
ySYgyJBO3Pkm+QauFQ+wXEgVKFCXaHInwKRCI6Miu04JnIfKB8La4xcKbNXsjwoM
fASZ3Dg1a+266iGbSAAv2MY9+XLroYllm4j7n4wCNShGmey6UZ0b+BTdoEossRo+
cqZp9U6WbjStJd3JXhf6mkZBXZnWgHRoe4Qt/HKSFs9TRKwBJB6AS6EM+mdpnfei
oUfUll0UWMtaVSX0/WmVN+FmFQbeKJba+hbEl9vBgkLv7m6ieHj5Jt8uDEuNOnET
/JKGaJkvgKDqO7nHvODi1hNoUVoIe8CkeNsTIixtMEsU9CLtNhKtchxLArWowUoj
DyymniKAUlVxjZkZ8XSpPqxrVrZSSyZWhkdNhXBYXrkaFmrwTOYMPU6Zhtm3rR8B
8XrVprGbwj95fCTibR4asDaco0YPv3Mb+SrlfsLwjTdYpTepMNx2jysFpiMObMXf
sU/K5rcMLHuKbEpHBbnU2++Vy1dLh/acGf3YVTz6NI7KebjG5FuWgxkaiweSaAqn
W4MkX0zSXWG3Owiv9h3M6whTzjDrSxPQB2t3DFI/QGE+OqMVjKNaMbFQtI/QIAyG
POX+dbLh+ycIgPL6z5B1ujLmDedVw+qIsYGp0THZtwz+TXgq6ykdM7dXOrz3DEur
QhgofViZvMzH4rUuCxF6uBx+PeR4ujcQ3DCp6r0JXrshDd6r1CYJSQUyKJNJzdXh
BXcTBeo/BFNey0vtO/B9X10amw/geUJCE207E5Gh8+WlNZejivUBNmB1PTwYtBo1
MCPfjnRrZKIROwgRqmjoNJpeTtggbPG55scFZIctQEc59Ql8010rKwaTh8YG3PTn
3lzTjDqmsw1NzzGBXOY7i0yIa6+VTh3TzrC8uJXWAG6VMavyj6jRehKUOPyYqdQx
GvH2ibBjxHLITF7xzmvCgR9xG6Apj+u83ct1qW9E/UpMNsq5k7WbgpFhSfb5+XYh
07DF5+wOamzPJ4rj4UjH2cU4D0ZZh19mqUzYiKIWfzH0p5EU9BZ6WWD7YXPEVDAq
6Qgqhs79Zg0Aiyg4P427zXcgYeAUJjjL3zHGNxWU9IKUmsd+N/GjoiUjyN/pXOpw
CzRUVRxy5pvb9KjfLvqcmoUWRRrujEr5nxkJw4+SSNV/qUawuFMfpF5rcONrXBAT
Q3HDggg1aAAm6LXxwIptGrEyAo/CKZ5FiaK4ajOnrxSscJNIFDqIYq6DoyUZR3gi
QcDz1LIqZPQFZvZUI37fauXBc8PFizfjmRNeqaaDutkqXxEXJIjRuIHWQG02lIpz
xOBOpS3ZSFhqy3eHxUY2d1RfAay/vGLL10B9jI303QcZewYFeFFr4ecIGuuoTmJA
N5SouXy4F54FbRtYgDVqaTQHAYCUy1VjVcLeNh38z3fExHig9o+kMPsNFz3zqXCF
CRdy19fQyI28D/VMEYfA5q2DsntNTD/6uIwt8Yl4Pmo99c/0XdURrNP8IMlVNaRH
Re/nEY5IQIHAr+JDKBk37hBhulGDwmFA8ey8ClQp/cB7Gep0pDoyhPb42r3Bm3uk
c4iiCw/+zLPogjBpAQR4tUmoPdq1n65YN6+yMQGCcGPptuObWHw6HOcWVrTP6K+x
oqgY2mwWO08Spl5iDKAXuAkAmQNkko2rnftN/783di6Ob2ZcP4SbnrCALrLsD9Dp
FKdJGLWh7BW6uRFXsQg4El5yb8nWjfq4+sMOX5tJmC9VJsuWrLl9Ht44KVghScbw
2IpF3bxqvYma02rO+Wu1TDaoMJwU8v5o/ou1gNPnvel+5LzM4HD0Ja4MgObcMDcp
BxjJgWKtjLZjoKOQGNb84h7mIPUJXlJYhERjj6IJV7lQPr5Ox6fxS8Rh20CxEqTy
D7P68iMHXcztydBp+MUrMKyK8vz5Al9riIbFQQw3CKtIgJuOkK11GPc76dA57OS4
y1eHzvAd5Tms4NbKWam/ED5HuXx7JpNQzCCZQ8Km7jMC6rN3R/2+hXEjp5dP/0sl
ijebMg9za9AiurAF4awoBWQkprew9J/hopARa2k84b08GxkV/MWP0YuTk9r6R7rp
GhZ0gNhmcALpAAaLKpQScSA7D6WBuFeJMLOsDht3EuILYq+1IykuFf96nvzN/sG+
X2QKPTkjcJ+lOxWaQ3HuyxYL4X0quRwP1fRjKwU643fMmeFM3RsvwkB6KZrga2f0
rJFjBGe9CECtRA9MchdI8zUCLSObLJNRZrXqOqTfksSQtdtC9U3aeo3rz6MBFfME
5YZoYij0ZE67B5ITnwcUu7tsFdFfpmcJ6gVPVAWURPTgN4fu1qP7sUnsKk1Ceihf
8L1TQ6zo4KaxGynaGgeKOd/YEANojXK2m3/n7L0f0jsiz1LEKGMI6zubcxgZqGAf
fCCU53mwsxUxBj+TLG3O9n6pUAoR97WPbgLH3IqSiwuFBRBTCTejhGmtYGiL6UmZ
OSVYXpG5a51IP8L4tw0npd7DKdD87zcpTEWS/VnXlqwAexyif9+sfoFSMzlymOb+
/SpNOxfQUnpXBBDg1SxWt4cPx1x+f9k8j6qq/bBZxtZoH4TQeHvcLjhdRCqPpCl2
hf3xwMcX8IguOKfahrUwmSXPkkNmeJjJPxr2h+u41MVP5mhxAbTW8l0wRwSs0pAx
AVGvrH5doE+MJ/oooIRkQKYr76/Vt2KYars9vCZcgNBvVoTaLtOdR59Ytifn1z9J
ViSy5BSs/GDyaFPB6vU3WIWVkB0WlbgowTe2lK5Rn8wLCMYJdvMKyP1CKrB0ZOcE
XH8A0X2gbu8uAw8EsTVp1hzYF8pHd+M4Xtu5fgQWZ4uDQQz+JNXTmB2wzMVAW3/O
z6sPHV/d6aSOTGAnU3I85CCagAizplBVN8akWzXhk83bK+27mOQd+KVvO+wmiezt
y1Tq/VRRpFcGAXUhFTbbPjAakrTaA73NhCbC25YLyFLteyFDtrAHZg5MW0y5wQCH
VlqcL2z3F2GY8n9CbzzIUD1cTKlsI4xjN9U9KesnOiPDZRbBfKNdsDeVn91UQVz8
/R/3hPRwisjIkSUlHougrdrjXFIVDz834gmAt4aDtuS8UERgOqDSmdqEGTS2G/mH
hctleemz4NIbIpo6wATBYkIDVVhGevdkQ49czVgMaGpXmX5uYwBz7/f+0GlZT+Q4
fHwoGUFjEZdRbYxG9nTNiiPaIrXVGZ3IzRzwxDUeLxpAuJf30vLq0NSmm9F8i7Nt
ENSLnz0BOfWv18HlQEXWD3jUaOUk3yn9TtcS3KIXBnAx9jqEXcERmslUyCkO/0UQ
+GUKaTC2kCSRgVZ0NBOMShIVKA+JYeCzInkuwHOEQxJDwhcTDqJ5NhFhjL7T3vnk
Hg+JCIIoSgr5/LEoNmQehp7dHoS0JvBGmcyCzDNOKIu9JxgFijHOfBHzUpkSwbCZ
Hrr1uPDYtsFulOrP/8u7YuY7sTOn59tzGaH1Pb/p2hguy30hhSYzjOTLn1+pPKCh
kC+b9aXi81K7IRLdbmKkrlJSHcSz00K5ft/7+/CWNx3F5NIf3/XBdH1JFxnpWWBl
wQB2jkOYpGruDuaFwALPeRHcg/MNMnhxDEuCMQ8X5jtR+p8yeRuHHuOa/PBriLA+
FM46HsMlmOANg0Q+f4U7+d++CPOiYNTlpOmeX0tZv4AGgyHaIBhjYMEuU2KSIf/f
+oiw8/lDVnd+kG6OatL7zG5SjiJWlSIe+7ZbRM+CvRRM3sFh8dmP/kTnsQ51XaDt
LiTMqt2RU2pzkmn61YXVnthhk+pCLL9rgN0/N0evyzYy3PG5h9JP2HE47cPVgX+G
mppNfF/RnY2FQWmAJJJKgxLDngXl6xTzebO9RhfTGkx5ZPn/62E8Mnj42VUWMHOD
e9wo0q02IC0LFPfiqtjc4CvnYMMEBKm/vDdaHLQ5KqM9i+Ls4r+W+/Dldc6updIq
rFdu2HdxNMrs65ELAs74qIswdFCYM6a8Js2z0igzO05RKgSDT5KId7RUwGfnvsIn
5qaXRXXmf0iGOWI3/8iqyxe9Z8Sc/bWys0y+8JW7JmcVAMxmwt4CMGXiS/HlsoyF
Xhcte3tJyohF+QaRwX8/HbJpBvsaDaacueJUx0+9k8+D+70hbH3YUjCYoK9D7kce
MBivFCVRbZYWQ9/cOUk2om/NX3ImTQ8mAd3eWpmd3IU1Gk0e38Qb4BoYQHmW++kz
caxxXeW8/IaRSZmoeYFhD6tl7p5mh27cKa8Ec3X2GaDn7j7uIR49L4m5/jAbSHDl
xzq6nPdzsq5X/KWi8lziWBn2T1L7xtYtAx/goO0KmOVHHkPEKGrLaBjO2tocy6hI
pf7PFIumWW+ZURSlw928VA0cN2kb42LRuqpkhj0V3Y2P+GQxLywU6EZ7SN4hz9vF
MUoeD3ghzseA184kEmB6f1vKD83aqTfbSmlKefFKvVkAO/XGSgdgE6ZeESesztDo
wPyCJnIr9lsMOxfHiROqWw39LogxtnQhHoxnlEQbfllbQwIeIunVWW5stPtuGJKn
MFhl+Ve+9iHNJPPYwuoaW2Ju5RmCNSJ/wJoZvWwKoWMHOi3krqj5uO1lrVde5gaO
LLGsoioqiKErKPuwI3MNzyMOxsz/yu+hAFwoj9+hJAcxgRLszM7jWWrR1D53N9aI
mtOkxHXvAXYjiYO3UhSwOn1vJT8Px06vn13ngcr5q8Wz5XmbN0Mdmav9FJ5RJwW6
NyM0JLcVlJmPoX3nWSx2i09U20tbJZCs2bN1Fg2K+FPJI4jt4kYXLK9HcgYjbXN8
A0sE1fDgOxnGRjqQB8yYqp3G3a5UpBdv5eGGlWRjgZ/ykvfMC8fYTSA0T6PW3wOS
G+swf6kfumVqwY4TZtxhQOiJLqs+HAS/w92cYYEIVkQPbc9ZfOEXlZ+BjG8bNDjN
0/bfxLFCs7DHDUDFH4LDFvhv2XZHcmh7zmmCH9vwVu8mjCEQSH2tWzkwUXqV0H7k
n3l8xZnb/NceltWQAUjUAaMTb/eThfgt1k49he3f++87DF36Z6zOc9KRvdWxbh1X
saEphCtUbLFAa26Haohqz+OvHvtB5K62mZzmSrDUPnRbwmFMkm69ASaHydGbwQMG
Edf+Az9FNKG4yjbYM0ZXSMDtdTy0QIDgPNCBpYnOJmxuvpXWUrAvOkboEsF/caVR
/wiih9cqQmJ09WG+Irofi52x9ChCjPQ3ZrHztHQ05fvuQ1cpBJEiSJgk1LsUZhlb
0mbob6faob/BIP8xG/RgFtUpZsJIdK6qJ5oviPXl7hd9pSQMaN0/uD8xbadcAo0h
rMEZfVHfPFQIAQF34+LVB/+8YWJOP42a+6au2tnHtCR2wgPNA0H9jmgHLEf1fKVb
9dXlj/w7k3hFfvWy7/u5/Tqs67xwjDgPbnbwZddRiBUxXS/xExKyi4ivMXjzbFxj
aHNWIYMfl8bv+xG4kFiLUNd651cNewtxEfTz5GZb4Cm9kTdyaOXWZpGViKOs1wwD
a3wNitUB/uiqXAONaPee9+bT/Qb9xuX9Aj7fuP+f6LlRi2fH1PFBFCGunDa/zDCu
Zwd2HBPbRgaW4OB8NKModDYeMMheGHNwLB8xSLiyCk/gfKczOHjPfFVJD/w7zFEV
MYdhOveBzQ8t3e/06y+9DFjzA9/nmdbmXtvdU6eJ2dwYFauJ4eULbaCuk9kSx2c+
VhndZJQ9tlMoXRrVVpgJxsBmSAMERnNXbI2P4wZ83jLXIO2yRMgdsEkLlANVnMq5
ppLN1f38pM/20t0mIP7XUtqdDgG6wdiQc8uTcUHHQhy8Mv2YitnwV82w6x8DCAuT
6RwHufxfklcnp7/7XppWH6emivSD0EvtrCABG2QaOOOzuWa3TB2YbH+yoMtRKMUS
nAF7oOvFACOwlI/7Xf6vBRfqFEEzrEDize/82XpyFJNQxwP40g0GDbjlzsn2/Lrc
zBbaarUfRGUz4J3NswQd/gCbcDdcP2Itf8/Ti+TdI0MwRF4KlDpJoRM0+M3UZVze
WSafMGMl+PqYAD3bTU0xIbhtGTgStbCwpWad8sMsjaIvq1OkFCSZvmfiEY95Yjht
CK/CK6QgYLVDcMt0QbzRDaJYxgvVLmHZP+PuWONAM7D09f40obcS6XcJzWEMCxnq
O24nohWF3iIyQeo2eeBHQ3TGpmUxQTl8d//POPGK5uSp8bvwH3U/G+XXaanIRO7b
FfPwQJEjg4nBNZJ3zAcoYm86GSqL00MFoU3/aFJ7IS6eSFfIuhLchj+m+O84pBNe
J7mc2NEa5EcvaAstYI1VYR2aGCDMtbMmBIr/d4gd3/yLcNYxFYQmJjKtJ4rsQR4s
7ebCuG6t7YqEvWFDK0t6Ank2j57wMaQ5A3W/6DLwMzt0OM/gv6nTgTwhC5mVdgFe
VfJzmxeTAUmQmZm1e3mRwv2rr5JaGD4an7Q+LCv142Uz97HINpsthrsZWyzQeZHi
r/pOnMH9kzGDiGk9RfyqzLjVtg7Ra1FIMdoQojl8budlpEmoS5tbGEJv6dQ446q8
Nr3zb+jniGaCTiMem8WhoqbCSmwo9txZxwUdr4tIcq9Fsa+lzqPflgZJokoBdTL/
uIly8fOEb7NccwzO29PqLOmYHk27gQb5rSPm95Jir4vXiLMrratOQc9tEZZ6LqXu
iF/s/uly9GwROa/jKIz81lHxYRXe+HPTodlMrFJ3crvDXJdjqO5SbOWBoF76hn5r
aZ8RIRWgq9BA+sqZRD9tJBb30o4XVBBUN7Yyu4CMmC6BaQBg3VSRi7VmH2vdvWyu
ShTwEJLtzj8XhoDRlk5S7ZYUvdwLVDWemwrg8fTRJ+Do+sT6I4pDzHATpr/TCzRe
3u6bSDllQUN0+/zbJbMZjpalfDOIV8anR3n8CWpMXGwH+vX5oAMAN7p9fFpeofq/
akEFTRAlcSiBNMH23eJM9XKMMCTNq/gjq+78byXL0JgGaG2D9C8vpiK9xmcJgkwL
bICueeG14krvHx4OjZYGPKPMl668/forSgoRi0oAtBRXEN3WDhpD+kioF4CpS6e4
23nDNn1819qerflnlIpWVyBsgG7c5njPqWo/92ArUWmZoAoB/oakK9BKX0z0iQS7
mMNXtlXM7Qp4gouV+PhSk5YoFGbbPcBRQxjbIrNC1r791cQGxnELEJEQzrsqBSGY
mTmRJAofg0s3aaHUtTKBYUYnJJpKXphGKa06q623tTfaSdFUga7w4MGzoKBZuaYO
JfC0aNR5XLxYEZcz0bq198ogN26wNjgeMoXkIRQ7oEMxJxSWCd9knb+WaJ3U4iGQ
2NzhT8dEBh6roPLOmw0UMKZ4J2zSvAOFjNjY3yYjIiXgzhZLwieHH6oDNW3Dw9vZ
gXUzWSP+R95RQ0OSyF4QPAXVrTi4GaVM65id2CMJjKYE8dk0jcND+1jDmonKtw1E
CBvFecyp8eyZF0WmKjYDCrqlkTt4NpqkMn+IwzJMz+UC4GK15O0akDG7uYlNDeS1
diAolJGQrPvA8X3irIL1FWT7UIDQad2NqCYykvYBX8xawGs/3qr4Kw1t6ViWooR/
l+sL1zNU+xGsNO32VZm+sdpeMfb1MHy8q7nh6XfKAYebSPjb6n1Z3LWdk26wKb/O
KyFicatYR45zdQ9jRftkjKK+jJIEfDrRcZAPp4YP5y8cRyanj7eQisUUJpdulUaf
50tcWybQx/y00qwDLq5v1XPAN3QTMbNWDtsId46a8DEL/jfUEa79yhBSk2a7gnJF
I9/afH0DyhrOfmaGqboFaBhp2tHUHabWJQNT6xUxjVVmSuVey9+Uo5qR+RD8dooA
uEpH4H6fYfGCYLKeUtikwOtmcraVBHXANbH03cJF1by9QaMqYdZDEnTbabpbqJdI
bUQdDthacjIogjoL3uGzKU05CCYvUNJjsLqYwoq4XzZ0M9rmGnAJ7022FObJfZYY
RNPa0kNAxXkZ89KwXoBvVl1NlrkjxWo4CybjuHJJnp3VYS7BCTjn8LGSCLR1/1dm
XXuOg7Bgu1kpOJOHfsuLyC2uH0QQIJt/yIQeY1YGInj+2KEkFTr8Ykf2ztjg8EhW
KtaIw3ZLr2l4CNvtQr5dBPZkRyVexdrFgWZSxDMcLA06393uToS/sjbAIwTXnqDG
InwzDmR4JL6L1R0NW8tsUClksKrLIoumxKzK6buoBQ4jRSxRNMLhH1s56FRBzY0u
bs6gqvs5W4+UK/DYe8bwV5kJHjFQYUMtig3Cd+7RbwL6+9N2FLtHGsc8iozwsTpS
zJlgsgrQ3sTbbVvSLFSg2j82inH0dYozN47CxbSxlI5rujuikieGnfqmm/aJgtFv
RPzgbrV6OyaSa/FkTfgrALQMLLRKrwmZ0Avjyc9yrjSCopHJLANULimBQwGJhFuF
Q1tadgsATuhy2w5Q8LuhSY2AFmcnwZTwb1UVH0fzPX8/nqPi9agW/D9Rbs3PHMnk
1XfR6rdtxCEVNH5oAdQQAgeRgWXXBrcUIgAcOrqERnlJoEopvXer83lqTGTBAg19
8tKQqez0fKt7RhBA5wJ+WPHftN/w0Nfpz+OMjcmRPilpr+JK1xGr2tmu92ItpGCy
XZ5/bGphaqAwYVsvvD0Tdaw7SpKwjH6h2JlHNjyHZiRDS9LMALoXd8x4A+bBZBs9
LY09EX67Dfd9ih9rfJeho5TRUb6fxjtFYD/0ghOTXuOuZM9dSzN9UxEXD4YfBN1v
Ck7C29Ny53iG/VkaXLEbK5pij8xRpIDMRVkwU1j30A9xmVI//+kVDBmvLv5zmGmB
SfXy+8PKTNobrcrmesAHl25Dyg+4F2GoRRwxtiMPgSQElnxCFea2pLsl/LvnM1vn
+WJ3+Ba90LArnmz96FkVgsOEzMFJH2MfYzZHlcWCtuijcudIDHElhSt10OxcYkoS
ReyJ8twHIJwCVyD8MUqmNm4yALkRie1t0Bwl3N8CYQZMtxc/PekaKih+lq1J7Ks4
7SG4YdHVTC4Y2J+CSpa5i3+u4hBe8lO5joz+e1SVBkFNnGX9OLcmK0A6pezY5/Fz
pYuMiQDj6Pl5TVk1Nqn2wD8wiHPANIPlGvFh4jx0m898a0wyaoX5RlzMMmyG93IX
Y/6Eue7aj1QyBAMxPpqo4Bc2KtpHGpdVSa4YkhmVZVzpszMRMQ33KN0QoCPXUZ7W
VWVmusDcrxs4JawDvqxulZThGJeyDyTup7wqrVuNAGr1vhYUeFszzTU8t2Na3L2H
1M3P7VkjLxG1crGeDJEC+mGQhhEF0/uzzXPZlcort18+WYa8x97ZavaeeVJFotsZ
GM0Ld5aHHXVybro0gxjL47IBfVBSzlEz1J4NKRVohEEHk6PeXuquRKosaFctRlim
QK955eJOqistSobzO42ZezMiZzGUxPVCuVNC4aEg2uQo5GYKEcGjTsWutiZ2o/m8
8MOl2+gfybxiUmH5uifFjgF6DkrN5e0y73pKjEf+129EsnD+Bhi8xM7jVxRTPb3V
dGV+OwEi012QVGmxPrdPN/KOrHbhn31NWU/FL+b0IduMHj9NoDF5LdiQAsMH3dNQ
8EpGxG3qycsd4P+k2cdHvgRqdPQuSeF6SDaCcwtRxtTU+KaN4aBnNiLnXgoWX9p+
OJ0eU2ttDW1RqngfWictP9TRHDLQZKF6MKxrOkHf4mw4rFIFyp0jNNLq2eFC4vxy
ua46NiSw/Vd9Ur+l8ZQRmyBttpS+TWpm4LjIn8QcTA3iU9dFQ384qB4ZDHNuiceu
fX2S0TC4QHFkNBuFGAYEMRnOobuLLu5kRq/DiNVvx4ABrptmAZtz8AduKJRxosws
iz7PX08gpIt0AzlnCzW1CQUPy/AV1+pWUFWETCL+BbN8cp1RI7eiRDSPIHYpGmvC
DZhL15ZycP943pPvEB9sdXninY9vK+E/+hdw62lPNNpexjwgyQoNkjaVjVIMEqN8
0aiqtnHpSPW4VOD4+X0LLn/Xyvix4acyfeJL63jD0AILg1TV+XZ2BU8pv2ZXO5Mn
TAr6DV/jRKCyibJ4s0r0rMZa4rNBTaSKWCRiYP8kydQY812c0GqOwqRdikN43cEh
p0i5d3YbuucSL1/ofrVifv1tLTdweRoHvJOuCvF+94aZH+BohkOR43mQtBEq9iF0
cNy6hC6pmGK93ACfbg/siW3haGqCq08MNeAK+Y9Zhcb95ADfQFP4HX9nQtHIVq+e
DaxOs3WIt5+iScqwla+C7eK8GlPw2wyh5LUZs4yWQAdsEeND9RkRpvGa5vVPhpUW
ByoSmP2Au/WoWOXxcUTNQ3mVHx2psql5AVLqJVX1XHskC9V1tdLwz1JYMjtMfxXZ
ngmz5IjF6xvv/SXCujzOHOK238y9m35Ik4evIbQPLGEFl8EGDGgtIgzjHsQ8eKwI
bQcPrJvqDTyR/6Bc1xC/8dpS1x2MH7pdOL7+SFsTg5P+KKU+qoq7OAZ0uZSolx/F
aRZfKFD41eSkzCxnmUaJhUDN06X1mPaWLnFSqCdAj1qAOOZtiJaxNEE2vtI0fpUV
79o+o1tAXyAN2wg/yWLCahbXgUYsGtXGiNIOLPVIqlN0IeVRtpak2ws2jQQ+g9JU
b3pH+bQyP0+gy8nhrvEXBdemC6wIFOzNPvc1PsBZhHD8BoNohNrEGEjlt8Gp0lWJ
fWx2CbMS+j0MSUhylaHmEsUNPQtWtRNHwICNCDC0IPGikw+iyJD7EdISH0daH9kw
mI+jaEUGEehw7aLbQPauO4M3Trkwy2vlAXLQl7Hzni06iwk8FjADRgaElwoBxf3N
FEGyMhBfx/I9P2Ripapz4exZN0Ak5jjtHcdKFRaCUruXyk3fALeGX6kWtelhTJ4M
2oCRn4nvoG1RX8/cYM4yJXjmIE0rJUCGLx103CKRnP0ISxwTA4TowuM9Ht5RBl1Z
h0kI8BKcaCehg2vSoRLyzCqLkf4ZETgk+8K/Y3z3hZS0JUJ94JKdB5wnKqlLU57l
tLElHLvIDQeQa0FA/koJJAorJNs8veM31NHe6Lo43AyOgeytFTk3wSsyVMjSyMd1
GzTHQD059ZgfQk8vSZknxF8tkf4IFnB0gTgH87XV0ByzIswaDu9+MmYSVRvWozWt
ti55amdzvinvC+JmjME/AXbUWNkntFiMNZ73BNa28Wy0chuvWAThYhpidafQ9scN
n4R67Dzzdm8+ntvS0ohKkXNGcczPgMbNAdfxtCdrm+C7r0pTHuTEwPtGwmsNL+Hc
LxCo5+cmQvId9bmWqXsjsLYSnTH4png142uRfHo0/A779HZQT3QkKb4KLsbYGhTJ
W5T5/2UmXr1oiL1DUn5T8Dah7zomXlk4k5CxTlXw65l0j8LjMDtJLpzeYRFCE80s
x6zQiAthN62JPGmTDLyumTy3FcSsK2D+9+q1QthEqetL9X/THJMGGrNdKxVPblZu
iI1wT83VfaGEHFBTzExpS7VtRRcZObDfiDlfu9ZfHK4dx628Sn4kOjYF++0JfOOx
kHaNHXYcvuxnGjXueNPqdHl2oYIf9WQxf8QOu/u03swqdd4bKL/9vjwKMZRT4CYR
A3on914IScwaWMFZdhm5FzOiTROz22TR40qqZobveOqqGuawREuRarjgGZIEwfDe
7fJyARa0gK5U/bhy/61prHvtOrf/D2m6AmM/28d+q/IWYc/NYsJsxG77STA3XbqP
hoRChWI9OCxrry8ynr5zLhJieGJDVZRGCcscCMwBQgp3p+my0jFf+IpF/VN3QiWy
fCNrI69K6Vfm2RRncMeWMqBLyKZu0tUzqesI0zDmZjo/lvfmPMK6aPb16GZeNItG
YdBb3yFQZcLI9iAWJpWbl0UvpjCSbeHRXcsYjEqM+6SLJ2vnc5/F+SbvDZv8Gb4J
7svKwBzK3ndKKTeM6Vm5KgcCAnU14kJ1QBn9q4qjXu+xSsBTxfX+T7hRP1Vw8th+
TAcTKSrfsRc6NmW1GohcOdBqSEEoPrTG6XUCW0UybAqHoXxvylOaBIiPE+jXJD4b
JxC1DlsaXCo8tkFWAhCieHSjbYp5CzbLiRXR4lVj7tbEoUC3CyajwgpyZffRcIF0
TlfEIyYc7o55ggnE70Bxo9MhVjPWkeD0+iH5lgkwbJSuqc6TFMr0k5ggMLu/m7AT
f+y714B0DHf0eGuguVY6sY21mNjwtra7aHkuXKDeOf31keEr3k8PdnzMunkk0y6+
h6/NgFxRgd0kg9Ou9DCKPbrzfNbpqJQ0NBilwsUOMRhvp68CT03m3J9XBKFWoHUJ
Tt2AIjBKTkZ0UiXo0Uxs7+oalSo3Iv6kznj/K/NhA8wcrBAkh0g442NfsojME6qy
gBToHG4JHZLj5tB10eu7AHKn76kDV1Gqk7drrB+euoobI/EyYm7OyBdKwFNUjSLN
LTpgfYfV1buhDotrhPFg+HP0C13POaLIXsHnOmTAyDSPvvYfmw5N02RSHsXpisOa
0wKM34gRUTDcA8F75460RZxGxD61JyzNNakQrmtbO4bj7gcbT0NSpRWZncgLHgdI
Y/mwcCN9ZrvFGtV8zkfz/W5RUdu5vacKy1B2nPeeavAaaN8IYZT6PY2pO5WR68Ys
Z0a0cGsgOx4td5K+lQqIRyMC0387VNL2GrKRI/W/Uavrk5WXdk6qqKdCIrr+tt1s
fR2ysoJl1RjAuhj1ThH78w1gol3Yk2QuoNwt6QsgYCFoOHLWFIKAylF9neSFHDIX
CuKF3LwE12il0yV92lf6YC5kyUpCOtqmKACSSP+cReVF7Ss+0XFi6GNNONZf7SLj
bSQe6IEBHvpSx8BdQH5eAlr2Iq3Vto281HLhz9m/V3KfdMyxWMvYbiBAgy10Tmqa
+PNTSQXK/S3pWC6LfeRIrWu2eXQrIe5op60bfM/+b7+1iBeJ7pOzd5fabyVibw1N
jFqJjsV9lDfmHSn8jF2ZgIS+Dq3+kBWw6HCYnfQHrNBfNgphptgWtjzEZy6+5jss
zpaFf6YgjOUiaVHzjzZRlBZFVA1RGKEf2ZCw9RXQ+jqGVdVHGWcRM8I+WCwdZGP5
SGNmD5g1RBM4laDIP41+c09rwBDniKLtTeuZFnLlAZ00utGdN3N6ZEz8+DueKfDa
jOP5RWlMlsbcTGRAU7Mp+tiHsn8w6z08d7f6c4mdUlpjnwW+UzFrJNM+tzMTt4BU
zMJxYroBi6H3FwaStIY+HQP2oBc+heU//ocfTnM1G5bY/gRBbLCFYBX5qfSygfkd
n7tdRaNQIMnBCZuD7cfiP7jKeuX43zdwsddL2aSSsstF0Gcx1L6X+stb21u6PR7d
0EMjUPcoPqZiA8+IR0dKMVtlyJya3N7VQjPL9CPNAtZW+JdwHBAIknocXBgK5g3T
Tr33GP9SenqLuZTEB2q44WFOmZtE1c/yFCsj9oyGYweDnVpPTrj+vCarwTseaaIa
L2tOZmLYfuANMBJSuLqJl4gVrobipaICoyll5T9l9usqdARYHl7beiqIEK8ISvrj
1vKyMUJwZGfxAqp2Rou/bZ8gb1RpMHtq/vvFE/+l+lfy/qUWPN5AYTcj2Jb13cjn
rybK+cxTLLEDXk36Ialb2DdjISVi4WE1XMwOv96yKRnLSKYE5XiyXQqMHvS9krhJ
YT0zXa7fwD4D5FMpZZSKTFc5FHE4fvFT50uKRV8ib1K47xGI2YrP8k+rosXiZTid
h+auQ/Y/0QdKUs2lDM+PTAPKBX3G9bBHJX/eeZl/Hb9f4kWiz6Equ8ohBYDE2Rc3
+phaG/T1mtBNWbbKt0Aa6Qt7/LQnxNCAXexeRZw8+x5iE5NSHyfcF0QTPBGEJQ7r
9fzE0uoz4VRgv2eY9Y/y5L7a3XbspInVMUQ/MfLlhOIb682VcXVeliqXqu4i/gzC
ebD178bFC7PsoSQCSJmvPJ8DqqVK3Fsp9eLNaWmo2eXoKTRrzqL3QUpeg/rhEhqm
d+5gPngw7GtCRT4pYV9JkAOneXlEDbvKrLbRzE6FHCFFdOMoU5jnLl+bwoHNifpi
vFwB8rmMhF7DqSc6ZwCvS+PIiBhwVa3CpeYM77P2kHxhfyu7CXOP5IyLOOLaTZCu
jIVy3A6r/KtLE52M/5L6XgUsPZLyrqJyDBbsiA/9nd1KJA5jGxuIk0ibixU/KQNY
+0AAyDKE4XuZgCzeZd2kboiTcCuI8AT+8Rg74dieWDVtXkonuuOZzcxDqceYSsNg
ZZtFVJeIc/6n7WtMXHVGCfhYGL1396SuDpHScsj2bMV4PNrsvvUALHYRZ6uRT54Q
/ev4rhoTlFw9bITHVMcAu9zvv2bqW5qHHNiIrnWb+TT+8ZP/YUwAKnCssp5VMYhH
k/Ekjgy4MppfZZXWqdwT/Zissx5IqTm7RFIKvzNsS79jkLXfHxRbbl6lIduwayb3
DbgPjf2Qh0S+m6HV7ytJjgRFjFc6i1qDXfejtxxLDrAoVfJYyb6FQ3ky3rO3Cdbh
8sqY2wNnkvsrI1z/Lqjypp3WbhKOEy4TkuJd6ZsEUAasfDiT5v1EUgyraEJO9A9G
drnxs1X8H1mv9wSwFiXTZ5MeCXorxRpnZTH8p/8f7lrM24/7AJzumcZsGE7FAVhn
FusDOktYyhelWWDuwdBAXhzSL2DdD4KQuVGSwyVPQ2U5NlS28j79yJNOCoERgsoz
1FdTfCarXDhHDZAAqZoa4xLFSvl8X/ipq/a+HQ1obeHC6/tXjawRjX2mlTKlR/Ej
3VYGI/a4rT4YBbGPtT0es8cvfAQfHiktbl/DjapXajNKb/apA8422TUcQTjN2fSy
Z7BuANebk9Dzl/oVB1hK5AtSoOM+xGe14b67J3WJg+A+VwSIuZ3UZr0fWs2U16Ag
F94Wdg86693orlXytnjO956nO5gb5yqVF7ZHz6Moxh45U+B6gnTds4lXdXRek3GM
ttfLowL8iSihRjUpXRsZ1ysUYptPUiq0C7h6vlwQyIpMVJAuv0rI6uMkh/NYNByW
qEMbR/1iFbolDAVSbR3NnVJulV7UhW8io7jkiAsG2NS9ozvgnNF5opTMOHmQNLfH
4D7hxQRMass9tIfcdxlXft6fFBCC73T50giySaBVgKkVKdbBIDQHjvLIMeDzTmSD
HMyf4lCFHqOllIXrDj/v7U2PueSNI66ckq4xLBRH1qa4KiICSUibf0YJdJPWY4g0
fRAkZLuI2PxgsAJKNnb17FWCDxdBkT4mPFIhYMJOW98AMc6kULCCL80X532NHxBy
fR8ftenhXe5tEA3kDuqo1qaU+byNbSrmnJklS/whIhmeEukgWywdZoci6VzkY1AB
aFt4zHjb9dlHvhX2TozuCgRmX6kLGH5JqaW9IDyYY8cCTiTKHObMA3kouK/eSbde
++Dx0Oh7tt5JcYLqEx9+X0FrD486MoSChP2xofrv51+yNiI914zfiI7rMzheuVuc
XMzSqzN2D0Ek3YzZZefHungbmFFfF7o+8az3Mh2uwNHuOOgprm8An1qxpqUNWg1d
nrOITIB4vz8tQk29COe8ymEDCMtUuMxPzShcs64p5YEJcjCqhmAviHtfuJqgCZNW
8H+vo09v3RN3j1Gnz544vv82V/NEn7TTgXgdaQCnmWdgNjuJKvtLb9h+gBRgkMDw
AS85cd3aK9ritJFimK5KTSZeMTsR5wAGH8GV5ixglmK1hRyZDit3bD1bGOliytUe
a/PMNsesABkkCKhnedzd6vLrdHPt41veW1NcRXLOeQVRdCu3rF9JYXfODH/ONRS0
+dCNki62d6NFY9/OUBfvunztNxxLadDUaUI74gOlvSVAQvXpgldxur4oW0ceGVL6
0Igortc5rgGo7ALtWaubdKmS/Ajg5a30Nzc/XL4EGRDJCa/b2JpAG4T4JU2myQkF
j9nAL4qylZLDf05x67frZSd3EtLjjufov2wwb608u43dS8x82hAGpSUPV1JtPKXz
lJbjxxfWZiyrRzLPUMUKmzhu7hNYxb+2Cdj+KTPsufp8+Ed4RVh4a3wsfPSuK4Jy
FfJ0DTnrKX4j2WEosCtyZTLfxOm4WpzZpw4AktNhc9JQzwNVck6utxkDgkf2Z+2c
XrPusOXYDbr5Zafbc/PtLukInBWiW/DbI4i1TbdxED3mK1LPG2EQthvqljkIK+m2
8GRgiUCZLN/xDfI1xoxPgLdrjiix7s8fUFVrV84UmTC/Y/LiK3YF1mwxpmwzLynq
3TM0WXDmx/MELH9etiKRSIabqbZcHI4Y8J3TEI6hqc4p4TTKoMWsIRXoj/IlUfCT
xZMgHwfQZ5oR1Q3jy999zwIaEziRMlVEdaOcd5OZRrd/SxLbOSYpkNqIjhdshGOE
4FzgKShbmBpcmz3qTlNjSw/Yt9SRkBL9JuFlpHmhFK80IZ0EOXvDAIKMt6EpS1NQ
+Sa3Hbfspu2XKI2O5tTNw2LJslOp/dR0IdgsNKI0LbW3mFcbODKycaW+zUw4gBkx
P6ANBQr390SglHRowNU4ShcGmYERNA+b0Cwg2SYOe5VT5ftFWLP0tKRQwGAKKLoH
LshjI4OmHGPbOBmFou3JbqK8w4XMta//o2hjVGKxrSVXEqVlQSnTWxM1dp5y+JIH
9E/IYdyD5pRcgMNzcQpLim7dvKMUAtSWQx5oCB7cyHrPam8CxTH05atTpS10nwp0
U1fCZviujURtqkd/KYxgB63quBk4T5a6axNSGsmWyb2QWlSykjdLGsNjdxJ4J5l+
P2JNaw3v071t5lJ2wmGJeRYY6NjG4wZDDRllAvOlePhFQF7RPhhfpg2hCdBTR4Pl
Ri28xxq8nYrc2JBHTO5wYAXLhsx9t5ODp2pYLijCnVdkqZ1WJHjGV2nEwDHu8roO
UCHPljEXen0e6bkDSTmPhVKd+063hEVJa903jIbG7dDVscYa12/mLf0PIkiYrVsP
idi2fVr8kiRkr498C2lUbFyHmWYYrN5Y8xEZxq03FbVJuwXpdiA6XaRyz9CsBnEL
0J93OZjtph4YNxgwfCSCwWkibvuPDV2M0GPsdreBsbEU27JxWNK6kl1kxOuVxhUr
TA3jOe+9I8UW+ZXYKk7Fynj5iHORex5saMNJs+cjMcGeRlbYKbFm69Y8ldcMVWCh
vv8u4SWAhaQu3NHkU8G0PnfHseCbre2BfmRHHi4jWRxNM2r7oJmesI2X04es3eD6
r97ZfSug4edrRESmo3pReCVe/qrBDQV8Kv41J+/5SCES5FuIJWoKkMkzV0EapCVE
Z9WztsoN9e+nbSLi7NEFD3T7uhWJtAFftyenvlrEV5Jhh6IL4IL8ZJ4r/mdeo6uR
O6cfHfTMi5D+oxlHjN3DF0sDnTUVjLmw9cTbVyICOPwmGGeBa+AInDiM74yQLe06
UtaKnYQZLUGvFhoS20k2k+JrypU2v3H+g0wF89oy7sD7TtQYftOGBk0gNE+XKKin
UtJrIDIAbd8Q39MLQ2Ns7KBQiP4BKKxTBF1HvZt47QituqtfzjXxtaAMBIv95m95
b4JToacSDOrLvNtZJWPsWcf54Ezj/SCGPLt6DmptPSy+GOlr2jbI7nV86wQdJY53
to5NfH/S1wEdrSAQugI9AzXveC97G9cfIMYwEnvBVl856Fqeg+QOEFwzpuxONfW8
5QNiWin2XQGEJtDei0DTFLtF9R8VM31jf/Mr7CKw4bUMRaaQ6mFBgc9fDATyGKv0
6pfoU41BvkYA+09B+IcijuqzWxxn40K0hCY80qBcOq+ysXvsfHQG88dC77makOR/
VWvxrfyK0aiXrlW4+71Dd46uuB9i2IBJyGlwSZWjeFOPFr/IFDQcRny8JPYQIcY1
JS/FgEVPR9zzM2hB3UQOTXz655444O5eci1zn4MHg/IRZ/dpd5Fy8ewrsiMCCqhd
VUMf3J1xHuKFbh8QyXdMsN7IIc2lBXMxLF6l45wZZsAkj7r1160gNltIDaDkUEj5
J1YCrhnOosXLssMw17l3uEluDwycBob6CdOAeN9RDHIa9y8VvNdVReoTJLUurWLQ
a31QH4KyuMytPWtp+yPyvaEi0fG/cZE0IVtXsy3cYeUVNR3xGR5DtN5lZVy9A3X0
AfZmaaElUFfiCm6+jngdsppwC/P9v85+6naEAl8Afg02z7Qmaa5afVEN7HfIozCb
w8QJ+mMId1nbvSxKlRLanILg57bUzR6qqQJd0LCG3q/RwQSWIrSbS44e2/gDHmof
ILtPz5QvkNuRmjG9h1AG+gjtn339VqwyCqtC+5OfLhNpzRNrIGXGKDQ17kjy0l+G
V5nQVEnO4IcDBNZGtN0Sz7XM3NMYk9R1ef4F0d6XSdtL/i9ZV6JbBxrS/7TCbm4j
FajjPg4upRMObbuuVGoEEyZhfkafMoQzGRZwwe0NIbhy9pxQBgfaQbg7RaCwDFht
FhUPfECn9+D3Z+7x5hsEotr08JqiFZIPoSuDBwdNrlHDV72TS8ZqJpvL9Kx6mT2G
0bfWu9Zzqcse5itJyGgK8oNNRoBCs7+eOO9uJsSTefWprHQJA31t8Z8rVi8eNUjy
epVj4PvCqkTYV2ie+1MwkX5cBV7PgwHFaav7XCuB+XdPLwgG4wKa4GCS3PKS0dWj
1rUTLO0YdNh2D+8sWjzhSepQvY36GCkio4uE64tjZifV6Bm03SmDxxsX9r8EPBE2
fpl4s7ARR4KNGn1kdA7O5Uu5notYgQJTSEgyKM1dAThXC1QIQD57i02neLlgQYq/
0MpZNGo9aUuI/HNKBmbMFeEsdJ6ZQEfZ00fyzch+uE+8fblrCRsTmX06ml0iST8C
Euzn/GToNiG1rHARcNdELfcIRtS22ShI0clB5SiqASLkBIP2HOc4g74owxsXkXUg
6jeryDngH+F6wCsfGAlK3ryTle0HaYEKE+Vb1/DRNJzLjeuk6X+Sc5RdhBmdwPPr
LscDLsTjpjCqIGYIbKF4NtfKOYPxWb1VwrvOgPLGb8IYaJz43K1Wtcm/rp/vwhSi
y1K7THXKS74JAyWx/8nl9m8p3ti2r6smQaDD3LiKVILMhRqVMgX3GSy9kOatQ83s
IXSw/rBEUcMlVn24HJmXd42uZ1LssNAjlteCyyFp4II5LkQ6KSeJwDNEIzPHllY5
i99X4cQh1sWT01jTt6vEJr+GcTEtWWUuuF9BJWse6MsIqoUFIyVIdDa/apQUYKtI
EZiH29SWmWK4nADxHq4wqa2PapAIcbfp2RGmvW5NaQy5AKaKMYJvqtaWtxrTC64I
Nar1b0xWrXR6McPrrv7qU4H6T2Oiuc586PfKOHRfX4JvAc+xkr8VAjUej6/0NED4
kHJqnZvg37KYSXLeR1eRsH3kRrvI9yqFVRex5nZoJ23cV7zdnuhJwl2uEBGAUDNA
lA6PyuBDdJJDwDaiEl5oNJDCJNA58jzaNi/Grp4lRGYRmHzLILY8ZgJ4y/R3ylU4
BRRIbm1+jV9IzQDJROUeG5lkbCeSatT6hysi3S/XN3fwweW6cBTlWYovMdFV0IVL
jVwhQaRVExwunRLffWJKNZ9VcElLlpwUgV79hgIxK19PLuDNdVuCaiQAhEtJtP3r
5clFxk7CCstg1p7P5oIx00DM30LB3sJLm0Jnc8Er8jCSD7Te1MmcrHSkkqZUHqir
CNaplxjifTwXqn88Mt3//v4JrWPUwZb1Q9SPnr5gp8Pb8aP9vqvEsTvxms/shHYM
wCFQvuptHyjc1TNr/2VDvTC24YPPsUmxQ5DkuLzVOgENIRB0Xyd18+UYqZyuseN/
ZmDOxyxdBg+OK52lp7r88NkMaVy+MLhUIW3/y/GHrh2bD9aos77eIi+dMZfDHW4X
aDH20AAqenGV0Dw3NVZM9TALGlQW9IpVjHY40bRTaZticNjoO9aNNp+Vi88T0zgs
Jb+eRj08CLTenlwvXJ4ZpdmmybwRiGqUkWAOWXf3aJc6a1FaWp7LpyZrTHb6P5rv
T7elU3ryTw9f9EH/NTS5YyVfRzSFgiyZi2tjAcArzC+le+4bIXtoEHLNUkkwAUHo
F1/Ma28DMEbwBqtZLiHL4CY6ybAjUBG6/H7rke+6A7kGps6dXnJL6uZOcnQzcWRb
oQV/QCegUOUeuWlJXkQ0y/io4RWokBYSV1sVVkQeYIGMIctMX6neI9Tuctqgjejz
5kX+IN0qj1vozfpWhFqxeQ7Z9ph87wrj2aIC5OB267KJttuWnnSOqyawLsEQ+XyB
9Ly0ezr+TqT1/mnoGN/H5/0XHoMLuKvftm7/4Eset66JNY/R3blMse1ePlcHIV6Z
/hdN44TfVI+IxAqXyr59cRvsgzT0NcJ8kM1yopCCeqZcTNhYVzO/XQhV7V9wywj7
lxA5jF8Nrtma1fg/S4Z/4PGNW01xZwapWmqeb0JxyjoKYFAXJ/59vM2fGzcpiHlF
+Caowy634WYzS0vh4LgUWsMwD+8eolxotvf6ShlJhdrPtwmFClR7b/duVYitCEXZ
BO6l6Ka8uLnU6drAmvR7Pi3jMItgoFHUu2V6DkQMzYAovnSU9SrRZKygPDLNBiyg
p4x/I7cayOaqEBS25X9VjjL/kzFFtP5xArruOEUQtvo4nwre/lTn6wTc3Fux77t0
wcHtY2TiuS9AjcjTg1v7bM3UvsqZxO2u9N4ZmPQjM4muW3R9K4ZdBOO8jqA3HG+9
xBVmW2t+DkLQU9iGdnk8CS9aRMikXIya1z0ujx9mKsudDw2zDATog7PYtdR/cF2S
T50IrGWkkmkL+MnOApSr1738J4Jcyn/jVWjx6t5Y4JJKTiBfejY/ZDpUg28lKfAu
fNgtAqRRkU1hOogPiT1tyg+pAv7xxXaxkeGZWqcPnIGyD1KofMPAaOE4rYZ3/zAz
6DYz/5Ye9EdeNCfu2vDZZ48xnhUGD3hzgIc07cMFr8yiQEnfJ+/so6N5cfsYzLF2
3oky5brO9ygcdC72zmv5ZFtr2A3OyxD830WSNe4VZn01a/EmEUrpawTfodZlTi2X
fbj5deRZu+pLHw22ICpLtIgiSyZAwffZqWuRCq0xbbz7mJ4TCvGXbeoNVmeGHqJG
s9uqVaI6+Elx+4QFHhHLu6lEaB7PiZipyzswgCaaNS+PdaXTeX77w9fMO37Vi3dY
ALkOfpVUaipGPMExR7iSEoF2Su1+7RiofEAc/mcvcDVFCYU07M+IQTpahBvLSxAh
0EMd4E7NFIf5bJ6yMbam73lz7XTbFhrRatm1sIHVgQ67QD5DTfFE/sTp26JCmPaZ
ruQE6zD8gNT12mJuZlQgNUggogqLFkgDeeHa4EV67KyNvVqYGAwrW31sbrKcDkss
G7MawWMhadaLJO2sZG90eXii2gU609hyHYOycAfVdxHMJQnjz0jq7BfpPYi/xib1
GoSJlBy0PQPowVo5p8crZ4SaTCTeiQedRj+ehVTo5S1+yeevN23QL0yFYJxdsGgk
CJ70d4g5k8XU4+BAG/S/DF050eTN8XknTsTTUWTGr1gh+mc7jQLQUUgoyrZtjrBU
/U8g27M6BeX2AbKJbC0AzVtIslGHpOE5tBx4uVxAvdTa5Yh7M1E4iAUlLW9HdPUt
C5wfVsqTqilUGlZPfAlAzagMV92FnVOmF+NFgMWGTf5R4fRNLBm3JSusckx8nD84
UyKvdaEQhEA1qx2QgA48PxKmK+uq1e9QeF2Ha7O5urFH2LMvJ19fmJfH1Pwfsoju
4vOpEu+hs9BKdHvIM8dHeBFJVCGVRlx0OVP7Al/g6onkhXY4pPpf7e6psIcFbYAz
d6D0GSHdsfEG4EMkbDOU6y+Unnz8yOkf5tgr2pd2QLgOeWr14bDVnK6cY7jGUpiR
u+PXjanFyx/1O6gMXtxQ5gH24pBNnm4RvybNxOgOA/GcnZNrMDXpOZ4krj8l6mvc
DPVuaT82M2ZcGT5C3mKgcv+0f7OUBdHvnF24MY6nX9QklVcxWvLKgO1CJo41Nou8
bdSsZKnrnIIzlaVnbkdlOr84r31sEWpJVBFNH8hJ7zRBBEGgFpVIS6AS7l91QkGO
3O9/9i3D5sO/epRNH9gTrr2ulOvhkcQdq/sFAIe2cTad52cABmPZxK1G4UiuklZ4
LZSsbkB6nw4TJ5tIr/awxzvXTMwvpRSCpEq3am0LF0ssRQqNHt9lEU6bBdjgTa+u
n/1yTb9WBHHk70dWsAxMetknMmYpjkzIkQTdDouLt8tHK0+cEyTd1t/P7EP7YywL
hu2kYGADV5MI1C96ofHVsZk1ItVEo0dDHW3gEGeaOVfGQe3Dilkb7tHAmeolIWbQ
Km0Utx8Ckp+Y/VHRBh+Ww6Xzz84w5K3R+/pkUkdCJ3rnbbMc51kAj2Zb5D80QA8p
bDt9wxVx4DIwIn07fczzj1ptn18t7C2ILRySvQ3u+YOcJc3VoKGgUApTaQW0GCv7
SBm6DmWsdcm4V7Y8QkTZOjZZVso+frXFJOi7SZbhSMEpBh5fZj7Hm6IvEO35g/Lp
gc5OH13Z2Hcf3LW88T9NuE4lwvksW/i7GzOt2kj3kwHaMUVwFZtf3APDzjfS7wt8
+hUp4CtbLExdTHBahiU/0RVMpXJF2bNzIZ9JUr/CqWFxW6NVvU7QqX25NV4Pxd5z
xISk/DlvI1BVIu+9Q5lgj0akPxMiirxAlZjs3ZjrNuL/qVEd/+sT5CpbfArxy4XB
MTjhg4EwXg3FDjpB/pyDE+Oga7LBqryIWTLnHM9WRPzi4zW4fLo/mkwpsIMuLYA2
+r9+PzjhqCm9jEMNnU8D7MUQeRZ9L08d+hfHSiWHq9PQVqQxGpNT1rUVh9EgcvbM
Tk7JZz3u5FbkvP3Tzn/TdPPGD4BjvCn41THuHxuKtE5KBYOjrRNF1qc1ydjBkb80
Mrjsu9rvQyepxqkIl09QhQoIVpHZxOD701mXClIJg7LVgWOStQ6zp4M14DvMJlmi
g+OHmYsuybeWGKaDr6s/hiMm9WI1zWVWzq7OewTuo1G6KtCcN8dE2QqtbNejpqBt
Xas8EgCvNHOTZrS11WlKvO9ntQ6zQpMDT4NSlrIvsDvUBOf3jRpbS//BEthiYqc6
iSJEnb14idXHiGFvxxsHoCQn+M7OM6cMlQ2cDfeCqVHE0ov5z01ca7va1qW8rvHL
tGYGaA9V74V+z4pBBqMC+84Ka8PM7jaszwZyy9pkFXjFIsosVK5bzwJhDACnn3Kj
y0foayGwDaTZba4gGtdLcZnZhSLIm4EE8T7YjbHp2jlRJTK1d3eoUTEZ5e2YN3X9
RqX7NwyC0KOV7erJwLNi4mymD7PyyvGJxQUoGU6fVhyuqq0KRax4iqFrFpQXK7Zn
h0grgwd51AL9SCpoOz/UEdDiW0h6eEztiHkEAmIJaLXX/9X3xs2lYBnjqhQdf97s
8YtJ81Brt4a98AyF/dJHHTHOJWOy9kYDgw7Cn8MT0nv6nxE6o+E/bNS20ZX0evKw
YrQTUhDvfCgSwHwzAhhrSjeXo7vH6bu9Dyo4QrdHXORbQ7/kes8g+8vqPE5GEvSB
wRLkZg3hdSd/VOx/XktOxQbVXTKErto+kbKR6vdZi56zm3h7Yw2pxVxconY0SzVU
cjYnGoQ5yEsICX3mfw02CfUOgsbbRx8Nl0P8pkNqO3Sy4wvz8fDRsGOb2twSALFG
c9XmQkGSPOlaCUwknB+HQsdV4F4t1uSl7OK4zGhaSc+8zkPkTwlV9TY1Zwewgqoc
rk9tf16uK3wX5GqLDBUTXykxgfDLFU13T78HTpb4UccjfdlEsOwevwz4qjc8JMgf
xaZ8qaOo32EELsDQkNZKEDJbrM+2XNllCAjRGgqlhik6B4ue5FbXZWaXqaiCCljs
EcUAaAc/+iigQ1ASKw+czzHsUp0BxQpwsqTzV9UVeZj/UV3kcDWWVcVLUdYPm1VW
+8c34Tfxa6Dl5LzAIrXIOXyXUtPTGYtRParqoQ4ef6c6dah34addIUVNuIB4X15u
cXqCSGDSALyxyKc+U5VhmT+uafPVqrsKX0SxZiT0g5MRmdq0vUcrq4mSCvCfTleu
UjpKExZmTfU9s150FuvMavwCDbgqcpMY4Ry4NBpzE0GowfZAJaMSw3YREMX/JKfC
7oz8DeLq7KWCqkW7ZRzeEMnH++uELPXts3Nt7bykcPw5VomdwUa9N0fMGrCZIvX4
kV+uxiuRkE6oTFXuTp2SN03cpiCvOagpu4XQ+DJJRLs8ZriJv8wXaD8lo7PiRZ+/
DUif/r3jJ+WgeVgeTJ08ZGualikYXV1UqDgDaeAZoZc9gTnE/vOTS1YLhp0NfTq4
g0RzuUrRXLRo5124NRP3uEUvNglPmrKkd0LIGKxMaFc6A05jhGfTSgKxfR0F/AUr
PVpoMqJ+TM4qHfBRzEQEel/QwlBnfvM9Q13UyuQpyl4QPnuVITuV4tvZmzSqI3+F
bMLPZoWz1vH71+ry2pM6RwfzuoiYg3+DM+CY0S2cKrC83UWJ2al5a0dY5mkObIOI
zxd1ilxkZzYSut5U/ffyp4Sdi4mdVZcQGfTNmwqmEBUC1f+kOXbu3oMknTECDpGL
gYou35xFnEE7PNOQsvhvTtE8sdUdc7HUjW/A+1aH/i+9VH0YMnWd4TbVwSU5b207
MPotImHDvlv/NLJTSr3cSuLzpTIhqo1v3EhHQkZZYWD2WEMskNAIHHTNAsj4tTRS
moxNITROv85lpo6S0HAQPTDtnh2c6BO5IDyRcW1DzkbrcrpTeOGofI8xsXF2GZTc
J7EvAyj2Nzc738CAiHyEA3v01yHKSSw8yCXx0ZmzdDS4MUzvJWeW6G24gaW8zP5p
Goo8y8fXqjgAJnC4osi8HBaPE2A+xl5BSma4k8LgTOQzE+3Vv/VJWOli6n0uzRZG
pwGTBU1++ZJjbc4b0Nx3pP+r5jXutR8zJsXGsgE1vTD4deQqXcwvlwKOQlOlMjax
BUBdDb8MXU2ZNH3wcO8RIVyikic4VhhshXby+lwS3CsOq4ytcrcgQFg6drYzHImW
B/L92worEHMkYh06zXYf6XVTvmzM0xhREBaIlkay051NM7DzXNWnNp8SVmrz0uwu
gxWKja+pm4Q6BR4KMkLapSje9LfHYvqqFGPKrEDihEqQY5oqJorKKcvbC9WWsa05
Mz/CynKq2mic2JzEevoUlGoDM0u4pPMHQEAvxd9G5qeZIyCWUgjCZXSAF+GXfQZn
zzS2efiydfJp3p3gsVh05N/6mzN6m1hmmFI1NdpAckzx4YsduoFUY1JQaPkTb1DE
T4IyD6+hfUk1Cnx+4pGnSPcvhQrOh2xTXP6tWTvZy6GPmUZheXCu5j5N8vfH8u69
uxzFYZ5qwynJjzv1OWstWFNh911Ksf+uvmU9vhAJv59CFPjcpBTqOA1k/DKiDPug
ho+iDPLuakCW3xDHoy/SpodHE9ahWrE7EW5viIapIChKYlJn/x2/oqDAVqT78tA5
AwRidU5Kq3xiYdj5B+NDn/T2iv8EKDXOCDxt1uQVDowSlzZnDETd2Ecq1KWv1M0Q
292WN86zYNH/7pT/asNYAQy/sUZihhRBq9tLSppw9t3Mup+RcqWlu3fifv0M1iGw
1WfG/NplFqwkpcD4mM98vyBL0Yam7e+cmc8FrRagVWqVkPqLflL4P2lxpOcEmq36
1dGaG9P2fiw9YSMRjwKgS+IbsGuk03DcnOwIrlM3Qp8pgx6mPkrcKaP6hEG2mfaC
oOibiPwOYBg/B6VvPRqWgxXTIRfU1Y+OT211HkReUUjRZagsl4XewzYDcOHpCZ7l
aHnU8VOEzYpp7hj4dwdsagJETW/T2PPJk8OeWfBDuUDznaMwFx1p/t4VfotWq3zc
Uzv1qUbUiDZf6JMHU42UVc2yf/gjQ+shX3T8Vp6Ebk2JjP0VnHIG4MQrr8gYqwIx
hjqBiTD6uVYVYwQ7KuxHRuNAiKIW7DOQWsj5TW70KuWrJtwJsbeIjY4DwQ5usihG
qmPuBE7VbU4j2C6HhhPNAIFvT0YFQdwwcTxNqhz6V8uvl2lCHUgHwUMfjE1HWTgH
Zht1NT5A1M9kqYreQyr0qsXoFWpibb/Pt9RGkV0rGrqyb0DeWs7brWAXwfB9dMOl
b8LbrcGXN7C9I35xIzCSwrN257Rgtovkvhryg0lxRMWM1VldT2t0Qb/X1ljinEfT
1dlMn8HKGffE2OwJ/XxRoyAbBF1urz89Cy54U+DchoNQmsmXl/aURD/o53xc3kq0
aMkIcmiDsb98HWB+UURHRDjioQNuEzUVsWEbVRBq9N+OCC71/ofPUrk/6Py1h7hO
VlBDUj87JMZjfqhItZXlubnSjBl7ppgw45whxJptNMOjHGdQ/wv/506W/jiEOVZx
Vyog2WpVt4A3ESRsEnOhYAPG4ropZylDSsx1aysU06rJMHkTsQ4z1P51eNV0ae3Z
wKFnVmDNvD6gv79PfytQRcoOuFAhosD0bsOYTjChF3oZL/6IlpNzkjhlAXe9FfO3
kwx0ZSh8ic8Z2/N9f+qfvFgi5gwtv9nWiFdQu3eBxes/QkXDmgJoQDwbAL5Sqm5n
eqToK6DC0NmVs3QdnKfvg+7QPJ9hGyhbgJRrER2dxvUX76lga4/wx9xQ4A0drRGr
Al7BezWWJv+zzGMz4qsylawJ7LXlAO6OL/Omk3JmuvAw12TZlhs9v6S7qXZ31/gt
qoYVdyAjz3RL8AyCS9ExIABvwyODqumjN1U0ghvRSndL+AlAzEf2l1DSekyANC7T
LkWM5jD8iMHnXeNBwcVt7pnla6mBolxtMR1cMRuI2Lai/FOqMvCzIHw3/TOozyW3
lXDr5rqWPU+I/uMrOsFiDmW3OvckK69RLzwtBSxs1wKaaLGtLlc6WV/U7DSz2OQm
t/WuKxeHjwzSPTxg2/xNDDlR0OpzM3+mvc9kAwnumVB9waECLmgKFlFhoJaZyO9K
+eMyR53rQXVJZBJxrMZrmr7ILNrwWOFD95rdEjd1i1tqMDbs9SOmfzGKd6v+N4TF
KdZM6xcaFSmFkXajIqkb0e59yS99lYmSu7T2z+EeBjLOWsIbyLtxvAv91FLpfo3B
txJwoVSDGw2XryNJ6sX8Fw167qDuFN8/e+FY8p/Ib+xZTq98J4MShTdhPSQ366nk
tjsqwAy5f+IBitoCB7ylrr7HANk3yxUMY4FJCauG/oLqbPyzrld/QfRm37keVwvB
sATT5dCdwwfjYIr5LuJPKqKcZa9B5i6Y9kDKeZZr3xuv0+lpSp0X2zOL6fvSLkc+
wifACUF7i2CjCukmerbgvNywSQ2qBSegEdKvZ5qPifQ/yaDfzfaUoxTsziYFvLOx
Zkr1s3xBwlqOKBA2fZJrn05RnJL+88bPJ4AZsFDUI1IIGBZAguK3k0gxRTrh5COY
o4a1qw5k7OUT5hyCsv7px8b0evYpYMSXQIT3MAXp8daJtOQYyLElJYuANRkxvACt
X5HMzWkLsXZ5somMRS+JXxTWkgSTJ2HVtslrnEA2lDqWPBKlICwgw/eR0AtCqULE
xBQ0u0SLtc8XNZWDtI9nGKQb1V14bgRDpogpGdyhv1qdaEjrnET+VaDItCpPa8bX
O3iCNjnHVTDF2au7vUi29fBln2GnIFWfpVa4p5dwZ/3r/gh9m4Gqh02KEAzeC0lO
j/1PGk49fzHVhL10ra2ml0SfJZfJ43El6mibNs5SZXYsU+yw3jAk8vCjwH2TSwrZ
YwBdwFbNTK6v7rXEodk0l4ODaDO+UZgAczS3iyhQSUpXN5ZRabGqslyaZEI83A2j
Jhq6quPnU2G1pj2WZHDZ0EUWjOFnX5SvkGZXFV1+55GEOOSUjYV2dcg+doB4sN3T
mAfemJfP1/y3cHcXB4G4GNCinteqquBhXQ2DK2Qmbvi9x1xRDOQuuhPXMPOcr+GY
o+GGzmF4w/KUKhsVTjKqJUbRPCgEmTPforAXZk1wttulsM+mf7GDbbwblFPh04BO
058CnfmqcT583fFjbbalLNx6pgAsY4IO3RW8YZctDjDVBb7TeTVrK4gSf+CI7gXN
+3hovrySQzbWaHhNxw6MMJFbuukzMNU4eZkjphZRgo2mMlsB/a/zbd9nBiliXNG7
XlI+4gfrpXyBBlkVKJwKohC/RPyHY0cg/i8inGnz+u3e1vHlwx2tLUJZrbzM0vVj
LdYaIjoHyMmjI21fMEjiXlwsKJc44huPFkcKSnxpLInGletrW2D6r0Que5NmUS8y
iHrvaNUqh2/cO0NPq4QJfN+74FMtcTWC2gefA1qgUGqmDVbGrY3l0l5Rtki2fjV/
PHxlT5H1LqhFsfMvCccY3BCFqRpLV7K1Tw7acyPHd0om69GzF/KaYsgg5GYhpEvW
GJeZqfdv6n+daQZyqoEGo6Vol/E97g6FcI+ObV8YjBMX28AqI2qNVZIKl9xMalvW
s7N8erauUGE0sQNp8vtbMKHfMT8gkr9eKPiu886Ubr1MrfnR4sW+ex1XQ0Xklaol
KdcAUqCdY7TmjNQdQiyabfpY9PsIqyBZ09hLCfotetNgHhG0MDXNKuiuiYnpIi2t
S5VgjgIpVwqfSDAPubfXJGV0mYS4v9kRlyPit9/tqxkJkCmXGM1bjt4rLBWzDevD
RqUIjfS9BYhsS7PjqrrEWAGO+XTjhHkDtpjt3b5mILbmyI3fgUZQUKvYP3Nej3Ol
EXBsBc4E4aw4nrQqhMRleRPOsrHg+nK4Pmp767952MEGJeSyi2PQXyA069reWEG9
YkfK+aiYf4whkPl8GbQTp7zFAUz9KTsOFXWA/8tLn3TNNS6gx+FxWTeufbQVeWjj
mjWTERhXayGVjLd8M6zjrzaHPZhXG01V0F5sMndOOeqTRGozZJss2ahtZLm0czLZ
bKvQ5aNFllir8BqV1z+yGSGKxVYXpbzeI/Slg0/+jboQHODFkQsfyh8HRjiNX1vO
dKjRSRm7IJXKnahQwu13jSbtoS9OMZTi7Ca+zTg9WVGrn5UNqiLFb55/5PmYWSb8
zCuBBWg0crIv2bwRnoFOFsd2Sn9GtS5bRsm4DpEVQaEkH9k6v18E6Sl6S5GFWksy
Clz7EbBqeQTe3Kl5X4y8QPxCnkd2hC8eO9njDZ6OQEUmn7OblwhZESzsLC4KhbJJ
8WPGlKuPqDOFGtuktQXOKX7+ip0Ge8oCJ0kinenFJnng9fzZi4GffttE7HuZY508
J29LJQoMaVZ/+/s7r8UNFFPrdKoxUZZ243pXrcxuVlqTzpkFB6nM22bfFcVYm6NM
SHlIxuHmTd3jyBjHDBOcQSuF0TE8apvj1fODOiy7KxSx2bQ+62ZX8V++Pf7/B9VR
BnVfQum/lvUfwI9IATF7DlUptiESmun5Uuw4lP4SW9ONCQeOnBAx+JJpuwBAoTL2
teYqqLchE9WEsAdZP7dA4ZkFPZhdLW4gjKHP2Mnxs7Vfoa03Skkku4xtnddPboh0
KWFNYy+bpeejP9TOVB4YBzmQEc9X8mOC9cmj4SKQBax/D2a9Po5TL2i942JwpauN
lZvvD5rF6ekkPtuRmHuHkO7oX863wEReMcgj4ERJbJ/lVxKo8w2ue2d/mJ//fiyk
DTGCkpqRxFShAMXgPXj97D91silDQO0Z0gfTKekejmFVYq+nJMTrMBWDlnhB6o53
ODiVIwXKsylgAOrocurL0PYz1yCS2FzAgnE2DUn+R5lCOo+ertRIlS2PsfUHTpBK
cTb8ALckbiv+AEzdxfKKHwyxZ1CL5KtwfGQ5h8fgVZpmd6m6uB9oCq2WLam8HjiJ
VXtK+ml0WEHRKVArWjT3XWRDtjOg3DdkXg4wqq8nYS6PQEcrX1A9Bup8kKrkSUMj
Qb9KwnEAxvLbV+3iNuFrPT6PPU7Ds7hdBsUXvjUhJo42hWvffsXgSwgOEe7rJ5EK
AE1iVrcTMOx74LZK7MwEk0IGL4sejf9c8ZziPo8FjUb3fhe+FX7hvVNxs70dRl7u
AhsWpZUDKfNk5I81HH2O4ioJFrXsxXP2unIeuF0uU2ktJZNk4IpPT/uXC9zFTWmW
aFOilXnHy4RUQCcSrxkaMwUzq2eCj6ixQd+qid2opHfQR0fnsbpoLt/bU1cIb4xV
FEqk856xsPKKmYtOgUMjwYDzfxWrjFSin8M3ye0PA+CwhRdgZJEim8uHdxgju7lB
DYtj3fbchcSniEE9UFULMdJS4RiINrxai0fMEcm2QOhK2SzAob9IQEhY7wsizMgL
741iuV6tijgpquUjjLTgcJsDTz6pylMLjJxVoB4PSkJSGKyDxB6naUIBBzPXoTBp
XhR/ncL7MN5HsuGCZIOviosQxZWraSOBGNqRDaMbw4s+fvSaEYwBLk+Lh8xXD1fy
21pkw3JF2uk7kYr6u9xnKRBES1ytexALPpcyvAkmdiJoharmp4hL2n0G1ks5RO3I
GPMhB0arkUlrkjDlRFFm5W66QNJnFF13nbmN785gECvFg3uiDB0qIt0CV2LG40ah
XnIcUc5m2Hxh+wi8XVGJSfyrvUfJ2Lqr0lf51zyvUTzcxUNowwOzkZhXPyGzWlAA
EWoVJEZbq6kpjQxMRbgxaBgS/Qs0hUKSOGRKupmBN/T0Y8HvzAGHlzs1P5J9EVi9
DCFUHRmjdzykx3XLZyI5JpvirVWTRAnLvpudT/3NMLVtnAehz2jqDDAgGGeegQuQ
PXQXGgCPxEeNXSg0/vMJJj7eS+/EJyoHLcm4wVLG7WUwFyUfwLdaAREDR0IPbgAI
kHQRtfrwBwITQRKYS7Aybc9bsSvbUrDIOkfOvPWrhBniHit9uYhkxpTMEFJgqNlK
pouYnFCR9UTs+rlHAGpfWPc4Dn/i0rn1XKXJ91PybVwaeSlEpG0+f5U1U2aTuS57
p/X/EuHZCxVhDAtsAma26W6rfZDwXZ0yGJ5myPJceAgQY7Q4IcEvss/oy7egmvND
utfRsp2dMiqyOGIlL/psO0tE6r5k5AWQuFvEnlgLhYFQGWdK+Ackgi3u1zryR7O8
lodxUlzBnXb0uamvysaRxwTDWd7uhmWLLYUdZ8n2fvk6gfS7PEEZmeNx/UUI3GAc
cdwbgKsAsOXe7u+LM8MInZJMr5mr9Dm8G0PsrlVCpDE5PThDFKWlCHFKCgTa4eV3
3dB1+Fg/evYjZDIQfsxrL8HqULkniqsqmwPRwDcciJ/1kJ9bxPelJYJmSNtwXo2g
yx+I5R6lbw6QtTFswpC7pdwzmlxPaNX91v7r5Su8tlijUGK7urUKb6BiL4+QKpq/
74K3d/G6spks5qDYS8dacX7fDy6/9/Sns95nHeGY8BAOToMRjFkOfog1RLBS/s0R
YBs4n8jFmQu8owC9MicE4y8+fm4ZUb3mpvH8blbW9JaxpkfFnMeHT4QgAV5Rby8K
O3v/infC41F45Hm75TGmJfbXCj5VtJYAtPUx/wb8C4Z6bMOx+uTXtYjzJAHF7Xre
33QT7x7B2bKu7fNGRiadf3fxJytFcxOjK1w+daEgO+2GX1xOqITW5WDo1MV++OBu
2NNymO18awtUyndhpjjyY2z5EiDwvSbMZPAtSnEm1BiUJCpcus2o7LphV+JYfm97
IvyEGu7PjscbboUbsluPB82kUQ3Ee5JN0I1Rv7brewrsYLY6qRqutFB9kKUNYq+C
/ZfbTKXioIbyERUQizM1yZ+XuuG3Tn8T+iZSMnUhnX42xdM0fcxTQHFJtID4Eq8q
FSWxW8ne2EkRnmGg15zocR9ZeIqUzQMtUofREdXECpqPHeyui5aMezKuusPj2NT6
t4IQEbd8FMASFHTpUinQhFhrX+1jrTJRWpQnugGPMOUImQ9hafw2QIhEENKoEQJH
OS6M0Iczuui5pSIbscRP/f//Z14RVL+GPVuzsdnw7+XH8ASfIPGgfGSgpTnt04U2
ricz8FgYwnaD1imU1C5JyvO5DdAC2stScT2cwnZ1dUl+QxBQLcJD/apx/NR1u111
69HJmzRqm7UrTqez3KffYCTZDADOIHPiP/DbC6W/QOXyuX5kPlFtJT/9lavA25Ft
IOJGZRhSYycAAgb1/fgE6MWFLLdvXzsow/Tumled9ABDvE3kmoQhGs4docPsT+yS
osCSufmpBjnF5Lq/vUJo64plyXbrxFNdhRFxw4D/w2wg3uH9MrOe5TLYJunUyT+A
1OsTwbYd2i1+ebKyP/fnc/3PfubiKYEwUe5A2yxmCCNY4WJ87baLYekSAvN3c5LW
QdRKCfWmyZZoQ1iUuepodFzTEL9gf4/Rs1Z5e6C2jUzVIQe0mKPfGnlVp0sTiSEm
+oAND1PmLRMWrAEAVJsgSXX3mRM9SPgDdiU6uxmMVlr48nhN3VFuvZhk7DHFmf/h
2q56esAJE/XuRYHD7cHZKHQYU2eLA1w7IlOLXjoLr2sgbUxGsTNOJM7a6XzBhRNp
0wgPeN59t0jwUpTgdAaAw5NVAMWxHBGqD3wwhJM9NEpDEm36Q3idgM8zDRBz2m3G
OwPfhPJNF9aYwcJKraTKqzCS5lRCcuK1KB+bnxLp2COQvaFxUe2Lba62Mn9qgFhL
PlWgrdY0Md3gjQyenESHwhS6BMWNpuRuFRUFqS4zwg2o+VkLkrw9/7W60bJ15pJB
nQCOH/ShBvC5ts54FStjWbdorObN/Eb8rQ1LzMO32BO/sb4v0PN5nXhusr4tRPq4
n9oKz2l5Sr4j1Jhoou4I8ZElkiy1AlhTGMl2kp4lPEADjILyhy0f8cLUssKygceN
uVmH64tFK+HyJpa1t8/S3vilr5NMx7OseIAS01fvP86qwQ7rL+SimZdG8xaZC4ui
+JOt+p+1T/Do00lBWzKtCL8KagTudhXgZXSujk69KqOOPrZ3JlrPWErSsb/OvltO
Ata7ZyfXFatD+iXCwt561OD5EDbSc6rNoi3onwxj5XONiQVKUxsDwVMQN4TA+DbB
ae1Mcvubr46rFkEYcdBg3ZUnj/ewuj7aUeyy8UmmbgtBQG7MSQJ5UHWkD6G3XMW3
8tufnxINLixvkTloEaJk5ekH3Rh8p5qnJErdjVBP2gX5ZDJhWT1kdGUQ7m/70B69
BDE/Z1nj/jRXzvXJhQBFnj36tsWXGdLzGOYd1XLmiVItR1G+ynlfrphVYp8uB6su
7wD6SDZ1ZXzdoOOrbLRrrblSj5Wgh+Xt1+gKKeKBqSHGNYkuVangGwzg9JEamy7o
OkBuVRn709rd5ioiVgUBV/++OJtGldK/BEB7/H3ERjlpFJMx5tfTm46CCJ4K1QXX
Z89Nc1eHqkOdWzi8/ONGiHeWcIFb2lyCkUDJVX4QD4Zb8enLQf2jfGX7amN3m0N+
o+lxJsM+Q/A/U4RjytEgBv60pYVqbmcyD/a4MQMZ7ynFAp+NjV3ngi9r1dLIt4Aw
XTlhWlihbbiIDy8y/HkO7t3UbFqz0+zGSxCzq3pK7aVVfpkyB1tZKXC3AW+tiwdz
hNyfLOjSLGOEI0X8fqk+x1SveSC2UlOxIrj8lubAKokCUfndCLfS+m3T1mjvUThG
CpZ/sfZd2DofV5iCJDpZ5Y65lWDoXZdu21MChb6AaLUkmXxEksgPCZNy6IldFI6a
gnUw+3lKhGaRp/iv6XIkL2SfWsWUa0jk0vIyWNV3UMcNcuiQB5T3N/FcKcM5iaVK
VEnHYOkfKJdTZl2O2CYnlQcLsB8+WSFgPOkiepM2bsPz5FztpJevxX/oyvEwCk1P
aR+Ijwg8P3G/OQ9BFQGRB4njE8r6Et7QGJqIGBmz+0PnDP3Ixn7RRiXM6I0Llqo0
/DlS392wOWMoJr82V+KDKcGOdPeUSLLcwx/jlg5tQGunTADkWwDwt7wPiqabSfQ/
pk8hpC39E+W3wM6iQP6uOj3dTnSMN9kRZyLmghxghhbexbX5Vv8TNFRJEML18vJJ
OYdwAg5xL2R8woRt4jyhnSaxP5EBTOuajs65q7m+BtwyxQXU2LsqtYC9AHTlr/8V
GXZu6ziarBNpG4327Z0wCxLCpFWwjAwIE3PAvaul2q7zmxdzp9ZeVqY9GGtnmXA1
9GiOgpszPKzlfj/+GUpYwq2YSiDIuy1IZmpjGVAMQSeTnDXJ6UmrygHilX7WkTBy
MhMvx+OUmyQ81mY2OnUEc4Td4AtIpHQ2RfvSea0bZ9nzkL6Wti9X1YAe2aUWXKin
fCzO1sGJDIYAD0dTJ/7JL1gOoSstj0qp/af2yAbS5JAPerucdE4+sDiEzeAcJGSK
dqKEGapTsuu7mhTV+zsjz2asH3TPhg1OOswdih+OT8zB/zitVJMhOoT9NSXKRO2S
dIn6jh5JeKsPPDGowA4cyV4qSZwtPfl/zn/5mTur+m8fcEzwrqEsJn9bha4ssGa1
8EPW/fBxYAadVq64Pxu4sqsoGAmu74jfzWujS7XWXH8vTtB1bLiO2g4/iCUWA1O1
aA/JE12nHMN5BT/MZlJ6hkn828LoiNgJkzBT4fy2aXzORaFxTmv/MDwHCytLao2Z
Cg6DgFo59nE4+Kkef2HGo6QQmEe9BdvOdgQt0+1vrr+Clu//E299CiURavok7nEX
CVvQ3WEtHJtjh/6AynWfs+Cxoi5m57VTCRQ1BEJeLYG5K3xzZMmjbijXJqoj8je7
np541OzvTNDLzRy/xIz+45w55ml5Zg66GXnrR+x/qmWre93ZyXEXby5GB2nC2JAH
9+LaBi5ckSp8HzdZqfaOKj/3T0V6R48HovQQsW/Hg37SyWV8xUXmvF++NwzdABfV
LY/U6z/8m44bkVnBWRcocOSME/eQ7V1y9DQVSAasfvAWCr0iRs2WyWlunB3razxS
Qsm8/OYre+ZwavG8QVfUw9ltpjtDtNJ8PXlYssngsllZNrIuIe+JYqmwKFX2uDLo
zcvKT4GaVy4+bST+Z4z1Jux9kiLVBmtizL7J4MI4au75fs+x4qV2E/OaB3OOtUlJ
uVxA6zAO2SjCr8vMvMNXKXDzio3MnKBqFm4gBiPUvOtL9oSRdN1/CsQXqxHVHsTt
Mayrs9Xth2NSd0I88mPNihgZbsYTjfYABHung9QdPOmZZ2aYVCkEjaWRInyE0DDx
Fi8bGP3rr42at14zG99iCUtI8VpkwWW2FcnatE53TwOKVLj+X7UmaAgZqSLh5QbV
x2CEsfteH1fHcNPd/2te7hNC42tfpmLdvHDF341uRRYLXLWvedi309jrPWvz5UUe
FFNclroL31lsyHycuOgRkdaBT4XGy1tLbNzhIZyjzn7zUTdFp6dRazWzdcYm1IRZ
Y4shyR2RSut73kfF4L/AnjOXTsCeSzvv2t6053n/xsuIFOac6SP2Jv0U50vZ3S/J
brsya3YTpt/lwxbbClkF5++YDhuU79ak2hGgQFuDP/xeENHCRqj+UVvObz1vnPFy
H7QSVMRNBjRJ2G31ZPS4r83GauOgGqO7hFQxeY9Oeq+WYgdN9y+JYvpXSm9e6BMm
giwRn7Znl8IBd3oKIEq8DSgmO3sX0UdrhS0v/275O93a6IzXDFcYRF2b7vYVC2rm
nuFBFDy5R4yvzE2e8ZN3Zz6Hq2COFQc6oA5BiNarc9dIQCq8YbS3Yb49peWxOVyy
UyBahZq5GBz372HrGPFP+bgbj4/6lpYkmIyslha5yboIBEF3Nhbmh3jlBvQNoyJX
GKUSmOSQsLr233rK4wlqAL8VxAbEwpRbr7oxLMxsYbMxdKym3oqwvESIxhS/BpQ2
gE6oJqK02naV0E3gLHegbzXjMTdMc+43/+crLN8H7+57cKDq6rQuQ5TL4CORqQ1L
kZpEGRdQCGX99GPU5P6cgMKZRKdilLVCZOEL9Kx/djYkBfz7+/pdaOB2sVieUles
0NCDCfOYGZX2qVXtAFYKA0OyKiHGFYgg/05UBurr6qmS9zwkQeCkSDtYS6RWVDu5
xd0qPvk3KkSDhGbBOL6m0VstA5NzG0AP5EVwAy0VzqNA1w30iCeEGaM8/G8RFmnY
bGw7M99H/hcaaplqNlKH56plyfmWWTU6EYDDu2X9BkinoX9HjMwR9uLoPqE7pzQM
PWD6aPeT80i8eJwhOzf214iheBswy6UVMrgBWftPws8aFQKJUidrPVuOTbF+NaZH
EJQNdgitOL6wfqZOqnSglmVd1kmIz5ehV60ilg51vH+FcZGVPd1Dd2erETPrkb6W
tOcH1k5aFai6LUdsshm5PK2D026DcjILWV/2TFCIt7AQH0HoBhtEnzHC9giynyiT
GtyyQ3S0ECyHDrlgJY/v8sdFFJORyZqFLgR39e15usbPSXN9eBxdvYtF1v3nflwC
nc8sOK166faI/wCJZSnmg//2jDZPfnD+xWp3BywlbGOcrK2lVw2w7rkq2b0UMz3v
8XIR363BO0k8/JcPHMdCJIAVp9lXIe4oE57IO4R/0fHb141dg9jiqJkLsWVptFcV
YmHvE9E2/vEUTWyHf0X03X/qVOgJuQUht+ZB2vRGdVWdTuCNqkFmY2YU8/KtaaoI
QHUrHcCsIGafjJrpQQBjP9Aga6/sfjOruxWRtlBiLAzPs4w8lFW/rwW7AwqMf0OJ
DZUsCKyl+G5lVQ2v11xAiAGUzB0rXhnsD7x+KiCNblmdqD40NboTqMsDSRSPMwBn
xXDCqSvq7SZ9m+zSAufbSIwREAxS5ZhlQCO8f+cQtyPuAymKJyFNZ7Z8wjnvybb/
4ySRg7aJDlapBYqYdUgMxORXgLYuzlHw6Iv/7tB5WXR3QG0td6B7WYJqOfXFHdBZ
OYScF/FLIaDQrTzlt1CZ8GrZSKOcaIkcw1HlSuRvFG6abCj13/pk3++5YHEquv9K
r4qp1XaIA351juOnERLGAFSuLsB7TyfgvhJTZQ8ZAFtnkQ25fA+SPtBSzggxQcHJ
tl5epqAl5MXBZZyS5DPhXqzsA7QvdykRyeiD8fKsp+rvERYKz0/Fpx92ECgWiDh/
jSSF7QPuYJ1Wlx632dTjeeedjf6tOYmiompoMfY46I7fkEgOf+dMLM36LQQm3pVh
Fp3LvGS1jDcHfUP/qptrL6VxR/nPa6XTWZugPtl4PIy8g+Lv7XAB/AAO5pcMVx4Q
t3kBB8050I4WGAazwZLWHYCnLFUkI9FKcibzBvP+UcWLNVwkhoP7phu4ITtB2i6p
7sLzRCJ5RicbfjYZ5MrKhc1X+q9NoGbIc6wLY7Jk/p8RMFERlhjpDdWCq6y3Cogw
9WTjJGxlpU2bz4fFdJ6f+cttxQSQnbgjkD6oXnQvAVEUOXdQpn0bDlATploJx9qx
087NsA4t+BZGrzN8PddjTfIgBvoVK5N32zHHZjD0weKvVCDjv9vWe7FAVKoQvEdO
hFHnt9/qY6nYZcF6oR0VyP17T5bxLYFaO4ddmhEK/6ZbrVfZEVowc2xIaaKSYiuK
Sm64wxhl3LnC8++HucXGux9br6Gp7esNiSTnH4LYzQ+ezq6On/tTG6wiPW05e09a
4LYIIV+RyMstd9t/pgqBKeU1GQE2lEIyIlWXr0XAShFxWLnSBpf7utaOYlxlGXJ6
OSJyfyVc9BfjxmzF4h62+WoP3RujHA2Kqa6U/TOzGOrIDEDUrDLXoucwUEL8elQS
b4n9yskkXKNbLuKDtGmSO4PJXz8oFbu5sFv9in0ZisOacohyyF5agya0o5xiEX8I
Cv0NpP2dPoPWd/LT7dCU2yVUFyp2lIF2ezjvzQImvbWL3yXlKfA/JbLzjZHXhIJk
IEL+iYV8+NOplY+yzoU042/dOnFbi1+c/N+jpeewUsbhHclM+7JHpFS+6aidWfuM
JrIFY0oc0m9vOaQG79P5hAqnSjivgODM4qLAhLS0NhQMonqilTbYsNgKke+AN4S8
wp5FGKxqPMRitMO2TFhPiBy1s1mQdheBTK9NgybL8ciGYzeNUbYJilDbvDcPwoHq
Wz36T4UQeXHVY3i0bVT1Rq1lizK9f2oAgcuyslxW+fHYYYcD1qUBvAvahwcjHjW2
8IDniHEniim74ye0nQbx+1l4K2+jdpYPZ+99bPdAkILzBGm+V1BNve/VwGzROqBa
V89f9tvk+dSI890ErOCPsNZKTCRdvwerne7/RKubAncW8TWoMJYB6ZZPYgOY+2Ig
uMkdklANPGkBn0mUpYtgT89hTQOTbLrJkjDYCYgmyG+T6NrLZFQnJtiAcwL4m0HR
JORnws17Y2LACyakINLivO+ait88C7p1sPUl77yXzlPKeCC3BZlq9Ef/yy4QwLd3
bgsVRcoR05HQJN4mgMhIg9N1GMovufuQaiHnlKYL3Hk89xITGvLnq1H8DzOySum0
dyT/obbegcET84YZ4Tsc3h1vMzHG/aobkwy3+zVgaYCG7lsT6EnuQtMFEXFmaT05
qS10WsfQT2bsz6MVqHOwuCNgy3diEIAXqAsaWRjdmNY7cfVAz4uCiqb9d9KfmO9h
GytXMpvc1HQfNJV6PUzK2bErVOqiLfjpj+tvTeQOzMk3H1altcGDl1hnc6e6ZVjk
0b/ACIJuSn1hHFm7Hv58qt2a7SiNZh9ftrHGfukrcanhk/btUCW/Ux+ptpXRnxwB
Nwsgd7W/VkcTn6S+0fv3YC6AnhADBW1eMHiFkZwXMDPr/k3q1lr4J0SFFYWFIox0
b1M/91TQxkOtfI4SyVQ5r+yoImi8Qe7kkALKsnFNtcEu5/GPEbF29uShtKj0UASn
VH8Wq1X1z0sRFH1QqTsqikiLBfknvWEkTgpLyaFwSIV3As3jpEWZhsZkJJr4aa8m
6GEu48r0iroNpNO0vuE1dTfzRy+QevVOEOf/sUGLKpSo5XOYhQcL3H/KtTlV0wN3
g9nnBX/uWl1RdN/7/Ba4ZhqK1ZT400v4DcSTaDO/MOIt+0lWnLpjMvEPPOIJWVqn
+Hjc7GkJKZkgF6iRhWGMrpgzsRxAjEryd2cdEGWEQqcSQyk/Bj9PxWP5xVMZZI3H
tdOkfEtGhxaDZe+e1aWgD5Sef29OtIJ3GIeEwIKXxgK9nBezpZf/9ECsx2e944Y/
J22+V69MaNXXqEcO4DcFpGFYJB5rm78GXztvw7+qVbisFsZi2v9QLIFQwAhp+Sv4
x0l/u+hwin/b95nb+fVOxRqTUkW69ZKBHI+1DMhO5emECBA2HBDtlWp5uPr6lH+l
7ue6bdS3bi5Pi0NC74NduTFcApMnpi0F1DHq3fmUpanHexWEJHz8CICahv/Lp26u
XsYnzMg0QiDS++mXowdyZ/eF7xyjw834WAAyZRUODmprmj29XbdoeRDwhOcWy69n
b063y+aws+iA84AUOF7AZy5HHdMJmJi/G1MCFTYwYNC0atE6j9/JiBgMwovIoiMM
Sxp/zV+b3qu4ltF0d6s3P5rZMfz1IPZLjo7IfGzsBprrQT/xSKB9XTURITOo+q6A
Shwm2NsQozLft5ujvB2Dr/wtSWC3evHTi8XZqOpVlKqM0oRau1nUPpWWCUyVzSpW
PIXX2Jx/B+UI5oPmYoLR0mNGKDttZ4KetR2PJfdenY935IdsLxZcPr17ua5KJLtA
IBrEQ8a01VP3oD6mm1477YD0d0tC9isEPsUwwxupy1L+T2mqLZX4UBYeck/+kEqm
YKuKa05VhtdtKY2q06vrjO0GQCBgikA7Z96XHcWnvNxR2obFXs2ccEFfKuzN43A5
fA1Jt4TfELmQoyEjv5SLLOLc+9qnZ+kmlGJUt090TzSjcQrUZG5b4x1+p/Z0KES7
W9QSyHOP/APB243QTCgp7/6wmiE2AJR7P9o3c0EhfaWuVESVUvt6XXxRvKj6yKUv
0Fj2esDamYQCPzu37gc0miXjMHUF85N3/oEf1FLvvlKwQZIMApZYc5kT/wZegYLd
Vj+8Fagwpr3Pd+0LG1J1piYVP0LnlVzyxNosTwXXVH+/KTKCa8P5IgIfwStkVC61
U2VTrlCcibq/lCi8cOhyKF1jeGwyj0uCR+ia4W7suUIPLvAxjc2ehJh9VYLY5qJO
iUuaoPZkHgUw9tqrdIgIbpLTUdnt6klGi8OC80x9AHZ49ySTSPD/6fd6o6s7b2i3
1PFR2BXHyJvl/EYdaOSjbbPck+auE6ovOeUxaI7zTGGbA21a2Tyc6IRVQDmd0+0j
yxv4wJUFqQwWAOeUEj7CjuHJRFobouW2wbwBShmjpohqKOwIFPcpeEzKicq6EFdy
NV+fxSHPwFSucBeUutXsT2WbBoOhoOl0TQHwN3s9bfZM2etbRRAMm3hz7siVYWHG
AKE8mbHwMcEIbo/dt2SArgJvFjCRdGdWRBaeP7IZC0IZ6Wjum7ZKDRT/K7YpsTdH
UCPXhcCf6yluyf12yowqcyrtxmW/oJhehAf1HPv/L4CBXUXgGYfaFX9tPxYB0Tia
UTn3wfLzobkxthZgOfs9hQwFYGmR98kHp+oRRe3rQcXPL8Gnja7YM8btB8uJhCHW
XZBtPt4XpRD/bXw6M7HGps4lTKL8taC48P5FD006zb5LjRuYk4aT3xKg1bZLkrA/
gD9jDSOcZ8/ZZxNw0/cM1cPEmv0ik/SGGSHkihXteh+gdeHi2F0O81D5UHZuAz1f
Lh0UpAzXviTgXFo6geH5SWf1a/+3JpktHpwnjmhYEb0ov/odTliehtiPLTJqel+L
igR8M2Ud2sEC6994ZvfIQ31ylTdLkxbD9s7hvOgSN5RHJOJ6REFarnrBZZ5BHZHZ
ZfbA3YS5G0ADmu30IvU3+Tr3BM2HtWUwRsD8b22U6j7yiuVPpnWEPhbUaIOClay0
wFmEkpQvOwo8kZToroioH0wJ4Y2MgUUokZTWHYl8bG6Bj2b5oTNMlkMZaElAOEGo
yyKLEn4Ajq6ld80YltjXmdpk1IUUjRPmnftsS87JGqgHBj1DBfhIm0gFp9LrYbYX
8SQz6WE7IE7Vgm3lXGjbLvIsM4CfkayeN/Vjhu0ZEBsmGJhpNYL3j1IHhZPeZhWu
/z+wPSIxCgvksyDllyiDTCSbyOqz6g+0tkq9TSoL3WLkD7toxO5Z5b65w6NGaLBQ
Ly3P+nEbT4K7yprtDUyQv461c1QjruzFTVYh8cTyBsC9ijmFRcVhxfC/Y5GS3Itf
qEV25GIqDcz+iEYVluxDmqswdiy1MTY7qtFood7fxOAYLNrb6Rez/Tmesqf8Hd9B
thpq+xmJKeuSP5SyJwwh2kBcILhdwc9F3cyVZhXdgo0lSSmpWLMw+SzYe82+Fz3T
iKoXl9Y4vQvI2vkh0ccVR38WHWUXzNpvei79z2ck0/WFOSAk+RyjhP12npJGicCB
XDYCIrSoHNA/Rgp+IMcn9OYb6NmUGIJjkurTpsZe9AVN8L6Dq4LN655xL62HSic8
m72WrLBKRmfPWBtlEuAMkoawcKquGUMh3vOa9TLnDW6eXWKAiUDEtxG+BCdrtHcm
tCT8iVjJwj/+rMbx/wODR9CNsuwqPm6FZjMRWtbkz8MHxKzBKMRUDIiuhosCVLDB
8VuHD87nZcBgDNHB3VbCjwDon15uAvT2dT+lwv69G/2BiASEMmnTm2ZCJeziAr0s
DSYuMUQ6+GK0QlJ3NIG2VtgnV7pwRT9zSIrR52wfQykWq+3m2jnjDzNIemMg3Vnx
bjAJuNJKnb388v9KOKGGATvMo4TLf1bvj1FGHhmWPZg1FaGRdFc8S+JEcw6XIdUS
4RLk38DP6DazxWLH+wD2FNEMc165R1g7GnoGgU/5Xs92YUCdbX24U2aSeJGIOFAA
JCGX8VEtkFCko9cSEiKGoi3MWJZ18qYp+ZNoutNWlu3jX4ucSNw4/C1bxN7smsYY
ptJsNWFWOXs/2Q/HDw7NOuqiuQKanBeQVFeUoh4vxTugWMOa3GrcGed+y6ZVTDUw
s9v1RvA5TCT9J8TLr3DHsoyHRDWLzDGhJA3QJZAYXxubCJScpjqj1XsMzGyUxPDz
eRFJHUqn1+SwbmOweMfXJKQB0egicHXeCN6eXG00IcnoxFTRS64Qzbo4HXyI7Exf
mq6eHEuECn8bfZeYX+4D/M/rWsHrDjQOlEFSyWi5vxlkXzu1mP9kmVjL3cEbvw2G
ZV1jvBa8ptR8PcQdG9pxujC3DVXxpV+JLeUO8K2aGn+nh93cfQe2Phaj42N25pW8
XKwZY5pYXYuVHXw/ygfD05b4Oe5XsWQmbsn4hQpojQKqpruBDw6H9M0ScumDf++0
a6FXnYnEyu3juyesrGD0CC00hag24cqi5lUK4kicHHeagfvXaUasfG2D4Ae3PvZW
BvE+nbgWYHKx18pNrqLiaIFLcNd9AJSTAu6orOMVfuZ+SAK0QrEt6GquO/orWbFz
gKnqsXU7SVQJfVx3zS16HopIJ2Aaotqw4sdXsFzmO8ev7wq0zaKmHW61FxEtStCi
HzNkX6/B0qhD5R1q9shRcP27Hhaksw9cYk+EO4R6FbjDXIHxMYQetT+4IemAJQrR
NDqSO9gyGh1uiP7oFynd6RidZBpH8aCU9um1A51BQkz4qmnbpLoS5apiiFRHFdNn
VGUCW6fLkSfK8Ta0mmleRQSsmM8LsLgH2kEFojDv65HVjK22ctir2RWwG5NNKiho
jMlovbXUlf1HZQM4sE6m59mRD9OPLGDa+awLAYaclf68Zdd5Uz78gXZDYGuxtQ7g
xLbQu98Gy1UEeK7Bfd3TIzMSunRBt/h1VMsYt7s6keahgF7455nU/v2oVJK+VJyf
P0htadXLUvina8FY6p2ILq6DIDV/N0voJVp4F0XAd1+PYfyPX65Zqu4WGl9+pGtA
HlR2xJo33mfco2ghkR20x963hsjrB/dZAKUWi+iOs5VPQ5UoTHn5B+arewX9PLO0
Dm59ztw+HvXziAn5VgzWEntwPfQRnyEQXfmF7tKmGRfdBKzKUC469HH1uXC04fdN
qBtFWlwc81qeRzb02+qNXfaj3Hg9FoAo4akRt9NARLy5Hqf8iQeeH56RHqOtjl4J
MPPQ7lnL6Pwd/UXBDzN5OU6eURAWuypkJMczDZI+STbWAdBUk2vHy50B59V3wx2w
eP0rEISiUuzKcypjUHwPg9UGNTCkHF4WaHVdh0Fq/mGIMEoac+e965oYd4kG56Ph
qpCyBnuBqh4GfmoBhDBvzOAWgrHwpXudY1rdPAyVaGxhj4tbYuQd3gl8WfORQIb4
r7yQG1bp9610sJzFKkztFUntGIrQVOGgw1rR+i/Hzx2brFTMRxRfsfWsSIqcFtxc
OdeXxVUZV6ttnkPE9CZDrpgj4O2dEac6wnjX1zdw5DGdRKKsKvReejrCKGBGNzEx
JTKQIiVng/5NC6aTCzrpUgnIliNPfjSt25JCeCA7vXRh0A2KLNdHu0fjs7WXkyv+
1LccCXGkJuKDOHvMImwWHfVLx7yykYv2ncEvhqfKo5j1toVecnJi/7leOVlYraTp
dMvqqdj3/67SmjQh2IkOPt3zcrAEgnKbMjxiuQkGmUnotzJh/6x2FjQS2iR3pNiw
5JgoGQrqNhjnms34hYd/Ana5Z91+daoSTiTQAd5J4yADE4AhXLwTwZKnQ/ZIqxeG
Lu9UYBlquEVX81YHYux85lDn6sxcWkUnB3HBh7oNN4RuZ5WHDR5qfSxZy7iGchrW
MOmG6xzYwlq0Tyg/WJ/T1RmgsYmxfNSFKlog2cxSXIb0KD6F5v1ZBU/5Yw9f3JTM
4FWmNXelnwRrchOM8zFjAqmGuqOEz84eqMjB2ped7IRX22tmYeZi8vxlG7o3Rr3Q
NCAnDmrf1wEY9oIgUY47caNokpvtht893xaLtOeZSaGYkFird4ovMMpST/jBmSym
tA9LiDeepwayvcbiJkBUFtBKrp9nM8NcDMjL6vM9weuTI4Buq6RlkZnT8t0Wut45
biCus6i3DCM1eOb5PdDCrjZbZdaTJSqLBzT/yTEofi+fOv/GteAbePDDoazdsbIf
Z1OkyR+e2svMPyZpHN363Dan38mZphminROURAkyROOpr673OIq6wMi5A7r9XIYn
AdU2la3DwxFhG6pYF8sFRyMRECTZf4EV1NMing/8R/qLO7c59dEcBsl3gnrijFyd
nHiciMIJ/j0o3D9KU1dL5EmmciIrHZ5aB55vu/ibEik2pY/i/+xSRE4oir8+RSim
TsVCJpv/HCgo5yNVHqLxAOo5cVcroN4p1v0H7VXaif67pemdyOsgksGipYgHEVTq
tUFoYyxPef76t+22BM6pM0b5XOGBT7zN+7JtjRmaun71eKxaeOfHC0oJjAdGAlU5
61HI3c5gltf7docpgzL7yueDZ9/+M6ej5CAKwfAd1WpYY9vtmwxNRlOTBujv++nk
FP3eTL40sHPNKI78jldNi5YveA8lcidWSvCGNqbM52T1N8EhVoTuJ55F429CTWX5
MyHOo79viBTK3e2+mxhMVZsovEzqM6KQyUoJTNvtSjxEadKvJmXiiMcmY/YKRR6I
iPyxug/2XOyci+YldQNs0CNl9rNYXEnvJIVYNgkoe/oGLTqOCzUvtF8lsopzPXpE
eb3vutOClI+mp4Jb+LW4LFwS8J2iHbBqP97P3Fdez42UhKudQiGHL9joymL3oQeu
Qdtcrg05gc9znr/Dh2xhO3O5Kxu8OfTJxLzUVnKI1A9G1Ccmwb+WM6MeG4LdEgAK
gbevhdokICsEHY2Wt3cUVQP9YNguEc1tvk7mpt1XCfnoejyv89HnH6t1CAMD2OoT
If7WDccp8mEdytkvmKSDKRVftIxHaB/yudf0GVUZFcHL+2tXsNO0ricNfjvNSCaT
2IFYXiEs3UoBMNL6oGqzwLtDz2YgXQUEXDunCCeT4QN4m5VSCFdtbEbzFPO3xVUD
fLi1BrwaiReEWOeroGU54+S9IEB81LRyV32xMuUdvPWV0tLY6fCjzREqF90BZhVp
BHCYQSjOAP3YEHEBdBkQbRkAS/Mqt5lJvAaq0EBEas2E1+3zR4KfwEwXByv9T9zb
QtcxhzoU2sotVgNbehziaGLvFDQ9d1YAKOYxpwiW/4guf0qFIR/kw6DM+/uioblj
b6g68CFBMsQF/iNTxqLtVVRepu1AHmpcfPY22SSJxiMI7lI0Q76o+rJ5HLYEPkko
4Sw5HwmJr/nEt2eFWDC1fDrEoWZ7RmVHWjwLrwJ9GXJjqAEDpqwmCWDisxb3YV3P
uD+Q/4fzgI1IeyG2DlR7Paa+57bQTNBNNUhrzyXiArQI5zQAYDN8Grud6knXtQ3J
6h6AKeyCZ9iJgzGSIszmt+kRxQdHIsJAnsX/wFmRvTvWKDGHvsc01Wyt823q8pf2
L3Ym/98juxdH5rxRge+p4Uynsra7oQvevMFDVvBhu0362KL2ZLfpoZ/C1izr06h5
GJC9M4RpLjT25bhs6SSqfMCp1IXt/hSGzxtBx3Ghtv8Y/lMRml5RfUsdX1c7IYz9
TUuzdNHjDRqnF09ZGOQtaxC2ND50zIFXTGqxsWNYRpaM7LrREIxzNcIDNd/tGEJQ
H57mglSbgMAKRjgYmBFTwyJG4RiXTqwtOyj7kpQj2Up69XWxYe1CxRtwAOgaLpQv
qYr9ubgOIsE8XaHGu3IrkHLuE5Q+oJwZgPoGGNoxZyc21WnVRoq4/tQdDgiTNUhQ
6W5KFurnvL9GcZzAQpj16VYMl2eJiwLnOqQrU7qLiqCcIPp7iMDwtE2sOWLfF4y+
00ocizp5A4byBL/41R5LHgch0x6OXwDbL2ChXNXjPggG5Z5Myzc0dnP5bCDD21lS
mqUNNRk9g6djLf4GEgKhUo8rboIqnksg4J3nJPMsegGMEHJzd9FIGAiDOZ76MeqM
zRd3K9L54V2SgcMTMyHQauiiUZfAsfRMXmkX6bcDkVINoFSFb5OdNE45O6z/x2vZ
u1v2U/SSZThGajKNUIRuXLjxAYtOq1J1mXZUOY6JcRNTVwekloCMtruRoCOXGZ7E
qo7GW9nHCBurHZP30tewvCySx2eomLM0hnMEPlOXwTmTmck/cHjFCUYc0WbyNF7z
Xj8RuyP3z1fZZ75RSg8AtQDa9VPHS0bcW4tS86s5N+2wGlLLHjEcz9CdO8NWwvg1
SNSDnCVvYKFbUnbgCbF3pSEIpKdMxN2ltUJvorrs2qB2AIN7KgssQUpyFGxVhI1N
ydsPVURiEswhfLsIcTeZagz8JkQE13TgFY7WF+LVN/nYv7nbyHMcIsEJxzNBbxCS
TWxrDqxv7X7L/2NnIJuDNMyleB+8iO+4XbgHbQydsCrg4abC4/QN05LqtjSJMmEz
0Pg/kQJ0FO0dIvSX7uhSI5MBENPNgi9WQnh/ph3JkaybEl3YWgQ5yE3L2aI1XCRu
9Fx/ZAUXlSqlrWCzq9c5MQAzzJ6/28JnFG9Z81KhqDJixXSvt/H/hp1Zc+1SavkZ
GAE/+0eGS955bXO2a92ReOUj4SH39cn63i9WN4L4P9adsSPafVpAwZYaZiRJ5LDc
An34CW9E4WmwpFTZkg09cNZX92faaBqNrLgu2ELBKzcwIUkoC1Y4jepkVqN3N0Pp
FjerBjXXFsXFmtdvj/W9hN7NNGVO1IMeX0L2T6G7yatCEpXLCkCXc9iRofCvD601
jXbgVNlD6VKwYjuHXTOFe4Jw244mqHpFg6RDA8zhFbuJUs5oAqfq4nQ7PPLXuXDm
Hn1C2rSl+QoSuRstS1wvsjNsjIMo1VB9X2VmOVAyRU09iesHEWu2Tz9HqEsUIgCM
zl1NHRAowdA0Y3L0lzivo+nnxB2SC0O1hSFOcL0gqa/8HSv/CNeH3i9iMwxl+28f
eGH3em/5DEylcRfPcxA/q3re+i+PgJNzddo/9rsF1cyDWZr5Eo70Mg4PfzcEQTCB
5IfTjM7YCy1HXhCBvMVlFTav5MQpQzU/+L6FetznR/Wxjht65XsKAwV+7uz777Ud
rG6+9g9ehcQ2wJ6up1MxA7Q6voyzvCJKYzrq9F4qY7amZnlxKYYRvBY63st3j1Xf
h0OhylRC1lIepU5ruXkEKcuSR20OPxAKq1MeTkilqF1OTeIbw2lZHA2Lw8vipZUf
qBUDNZ39tDKeVrVtj1ykCHY+A6lZJn1A9wDbVXy15K4tmg4exo1oM1pblZQOfjgj
KMlYngwhgZYCVMcmpsaMTZTvB5PzTgSewDoK24oJR6tADjgAYNrlK5TOfE5/Dwxl
/lnjshK16V3AVC4IX0jHUt2ZfADGKPjS3aMY5GRknZ+SvK6ssK1pPg/wF46cD83e
pZgm4uETsHZRwdmmupljFnZFW9QH6dB4WgYubOBsAbjTWTHvCNIDxLMqxCGxgfZI
v0F1xK0pTRsspqhjnKuhB6fDuuCMzlHaIfWMSHeNLfLmE6Q3G0nhy3eAVRjlwyFH
Bokd5R/dzo7AqucsctVOeJJh1pEZGdETTzOm9x7fL90UIt7BQrcsCdxFB6PrhI31
ocCfFJg0lIjX2Qg21nqUz4dLqi+OhqoxVGxD8jbsfSut+IYVTY3NLxo2mVEof9G2
Qd8Lx1SckeDu5KezF6ZFVNSMp7ZQVZDfxMUztl1a+30tTb+7av2fODZM4iTF98GZ
LzZmGM8Ct4FoLwCkbQNtAmkUkctZ3qUq7zGq/p8849gBhd7NCqGCb30WWNqDKEue
9p+k3XduVFGyMJCrbQ2v7/lY76f8zPT8WDWfp9kQalp81iobIzEP5yMoFnoTaIbj
lOLp8oQC+CLa8H6MyE/7UakXg8rthwjb3WCNeC8wikRSyXF5x4MggQdYMxhEwefb
k3Cz1VGRFzVUZOnQAt51TIb6o+aEWGRFU/v/V98gZwcfIXdY61Z2+9wBLJaceSZN
Rwh25nG4YIV1AXrdf1bMh/9fp91IAZEGCMrZRia9nhhed+0ESxVoVswgppduuGhB
3evvHaKloyYyUBeHVIN5rf9kM1NZrnV9n9582CLr+wXgZTpUH60BLQnb9eY6SYMR
7nhCKTe7KM6jtkN+KM8Z4dG2/VBdcvQhVLXwYl5N8EnwkmuTDY3FSb2AQNMKeY0x
CWKyAOVZHUeIxRVKVtvbf5ZY0kuKubhezEfV5cjsA8WqdRL9kwlEcdthAxySk4Ep
S32Kktdtuyh61ih91/QTA1gi8owQf9Brfr/PcuK0qbVANBtG+BwDwRIBIvCMpLkW
dKFwlcCUYKx322iEZOCvOBwVENFalJqHuiEeqkezxVaFUmaJpXqP7k341k5aUO6/
Zllj3UYQmhWs3M0xqYC3OaaTXCe+3w8J15xf4ucGGDjHTcYsSQ5qNYpz7asLhAzg
J1AIUARacqD5kciCeXKnwOi4gK0UVJAzNxbn93HCl1eXTv+j8SdW/fFCrsqAGvVV
E7+y83cdna9mDc9frb0ljJisNOEQDVLpINFH3owxFEV5nmjb0U4Ca+m5pQJ7EuMI
JIl3Trbf9bdNCh9TRq7r8/i5Dr8r7elt5CoesIAPERw3JqKeJ7ea6kyd6isfsofb
frviTNkaATmPRcFXDcL8HxyJWCu4wEJSE2x4/Z6PpyC9j8aYI7IdpUiWjc5BoUEb
6m6BNqY3Wv0CuypsAR8zL62NoIWD2f8S3pC+TvTNzUO4urLUc1eeNpEtsOQ0nWpI
CYYTUrhYEjnFDLsjFfq3cXhNXbyQ+Aq/fooDB0y00Lu56achZy1pxoHCoBVt9QX/
oGxEN+JPpbdhMCxqtHGLMiByunY2aVRsJdOw/lx1142MgyEtSEJaw90Ya3Gv8oQ1
JadT/6No0VqqIpUSi66OkD6unf3Vrgwn4cl+yZZ5xXRKGFjYb1HkZn5+cXebFCmm
gD7lcCcFjti9Mw0Qarc8PAG4a9k1WAygpXDZRINb2lFvLiRBMZ9H0SbfBDiMisZk
39ht9VQaIuQDF/yTAi1xy6BaAmONI2nLQFkziGRCUrwclMQ4rZtW/Mx6XZzWhche
CWn8dJj7iAa0Fh/hbM5xxG0bPg92Dg/DUGpdc5L9DuCpfXFmETEZ81J0zlOZGY0Y
qBAwTCuDCmbrf5+GosNCSfu5dty+U2mB7RNHBMwht5zceNAVr/VysSxjXuuTAfgx
FStrjwG/0RgBa1Bc8AFC93qvMxTlRyEcB0Q5ss8vyAKCDJHhWpfxaWXwmiW8OwHG
WdtVgLVtkANl+4oDUzFfUVjg0NIixxtkCp0oj7/zgu+o8HeuNHrSKH/bYahU2g9R
UnTJQz9UEpYGpt7FLWfB7ef3K25oQu7J2KUWA7pmSx0CLOZtt4VUd7zlEUhVc5gr
gHYbLkZlG9PNjXFI+dKm8WW3MIMLgEFTS8/zRbX6ainZ4LRr+y4HOl28/VlAkEkl
XUhi3JOi9OiHdDGRnNcl8mX2jAydSfZi3zXCAmxRC9z2vXNDHOePuWKu1s2ucutk
hU+WhLdnOIrAVDo8GCalSXBxCIxh+/d18qGm90Y5+9WyzvsBBtCNaz50tcEi89xx
OrMqw35hLCVxcTyhndYNEQV+h0pbv5b8HPePXH5mtZiaxQ29uP3Lg8UZL1lC0xLz
LdjV+Xf92b/c4IyKeRdp4hhQifBedIkuNwcMBZgWGtEj9t8rrUPuPopQUDKR9Ysy
R23BbC54b29wb1Ctkie255WRtv+hysu9mjWHovZvL0AFoFdbhGuW8rqm7+/YmGZ8
ERLwlaObwXX6NECqiB1NaKVy0A2Y+EuHG5Q89RisClTa3acCHMl4V2WNIEw+eZX3
TmIms0Cmtj/4SNwzZwDuSjY65Xqpc4CMzAo6/qG8i0vfhk2P/RobOob933u7ozwV
av1Hu+epEs5ixXd7BvVpzptAwrupEV0bFrtN5IHBwS98IeaQkk2vtn5/fRUXJ+In
wLJ62MBVYtuDc+hmE3TKv/D2vcg5ewnrcVsj2KO5MiQa/6auiAOPU3ekcI47LU4l
QlLrb0Ch8eqGHCYcEvieJfzgVVdKSw1QzNbOJAIiLakofg+hx3/r2E2CFqUt1kIF
CGFxW2lGqM6q3A81EkbZ9c2coYVNrhIwreyCBZFP7JkxSDXKWRwS87PZt9Ubr25n
ecl+qVAK9AUOUC98gDtZ2OfVjoGN6sMo5PmE3Yvfq9/e6ILHzWElEaCw3Kk/bV/U
CwqYiHINU7+HYo26pufRaI74+y/ae/ud/sG7v1wv7QtquKc6cE2WXX3ax/NKERpk
aqp6JOZUKqawxM5ALz/jj9SXUILGv+6fjroBiyJdQ6QuxEkpmrAUYX1TC9HwnI3D
L+jLt2HSIqm/bV8v/FpmqPNV2wfzHqIEpHyQVqSJmo0xYsbw2wC2DhlaEyZkwbJh
OvBlOEWvISvJ2TUyHMvKFe1gFAo3c4N6VXFVVGCCgtmCFRC7WQoiu3CSas1K0t1j
9Md3r/TgHuLiId7aK3Fdnu4zsF3z5XJ93LVxQQw4KncfeCPM89prl9JtwFywnMXZ
kqUscYTpUIxYrr9rRczmIHGtsjgpFEqJ04Ji93xI4pkvf+CxovkMKwkLU/ayFc9o
tpsW1k2+g/uDm0CTv/diJgbRertWphaiwjHbiyEc0sINLCWDdyDFSiJeY9BN0x4x
xDOiX/rgqR0OFUKqLGrkXznH4jGYxQhO/73QLRfrkVzR3E5aosATmAgS0JhQX45Q
ORtgqYzz7EoHsPL+U6wZtR2UWTFi0EkmTD2wpngLHD5XdBMv7OJ4ewVsbHZ2tank
bxF19KwH6ZLBbwcGaHWdMf1DAI5kuXSJ5FQQgEgHkUhvzTHlRThlFgCVsPB2Ogjs
ZagpYEkYb0/0DIEi5Pn7n0rlXr1Npgkn/E45nAXmrOJdFS50R+VAZJ1KYtCxWvAI
YbDozRZjoPpNlBT+MDK528vxf53Ue9wFE2HfbUpqzzkv0aw+/+nStSB7wukB/RXT
2YGNCyCP1pDEFWXXAngyg9iqxig7ox99RwqYSIvysoctM11YVLNWOUsaFBJbIADU
+Xb73vDEC2MYNOUKsEGOtlSmoFBinx8ppIZYCYer64HZWks2W8gRIaCsqBvqIRRc
QBp086nHQBRgRJzPbjCn/s6F2uAIywUqlqUgu8sXz1+fi5ealtgxtOGHpmjLMSEY
agYUprxKWSSvrl6xcoQEeSy8fTeJm2lNAiFbiPI38nuQ4R/WeMHWMVMNwKWCIK5s
LT3TrRKCueTMXbKP+EOVxrbBiUadkuj7ykqeIk5B+SxXq/uk2Ksc2dKi+mF2J7jP
qPN4L15ejpCQI71ET/yjKPERKMBOD7RO/BOdOzddFu+DcBHcVkFZnJDQuNF6IGzw
KUprnZkakJoBvwfDbP5thOD51oUS2TKdDfTYVqw+FKG10OhUmU1AbdoSr+1cw7Vg
8lRfXrGuTOtUYpiFtXLAyy90Y01TI1s0styuVtHnSB8ye8hZrPIsFG6DeYoAfwWb
YlTZYxfhMk5D2Sop9mNOPceCGdMO+Rp+Yu1FSzmf4B/MJ3QIjRx9wlMtxcexJ3cu
KuVbdor3aw/+eQWt+L1uNt91kfft/A+Q2V0a1+Qs9MkGNTPsPGhQ0yFT5jYJrzZk
hQyz478q+78kMi0Yccd3Dctp+spKnkXLXDvJHa6/iPDO0AWq8EBxZAscJzyLf5Z5
AfNTDfBsbhg41rtYI7aNkTjgyvN0wrtVpfTULTgttTekFAppHaWsnCZKmcpvhDgs
gPyE9T4wqmkwkdFn4lkXlM7rrIahcTxuILgKsqJzVWYMmKtow8xy/D7WNu4f1fzV
7+3ZWY1DuGMspGeJOLfjM8xcyXrxehSpq+LQcgCOtPGpoci5Y7HsZ/JXxmdZhnXR
yQWnldwLau0ghEEEKiQ7SIaeLz2LUF/W34j3yNehjW2+UpWf1vceLMm5hHQtYz/2
TK0ijDjfk6pYlTAI+i5nUEbHHQE4uq/z5voHYk2uDhDYSMWM0bsv5tkwIyDi5zO8
nEqcE5kyGoHpJGiatywGthff3g+a7sHFWGGVIsNx5JKVFbE2HPlRIH48FYGCDgSh
FZHDI7YzT2t4bYjaUPHG0kdgb7hctQJ9vGMg4JYo7M9ltQN9E6Qa0fmWa7yUeuEh
WTYHmVyxDAV0sJzkzjCvxdx09dm4zKQ+PR4D2/AJ5lm9Q1jC+F1gWLJgZx2PrRZB
janng6IVL8QMjHKMo8Z3ukJcsrT98gFu8d+eUiv+AsvbEZpoPOkNrgNwY2hkpWs4
Vgoo1+QFbUdJ4dxmxXcRPQCwvod1nbKoV+/eItFZGPAUZCB6TLlCdQD1b92i9p+0
LoZVhE57sV7J3w49Ket4r7P2mM9h9hEY0k9LYCA2vDfQzNgNTkbvqwvTo8IiU6Zm
5d7p+J87EMLKfGA6cf8vAec6hWL5NyPKF9uBSkaBIbVY5SGYpYDR/adIYdzqYY1a
lJCm0mqRwSXORv+MIM/OoDoDkqBZWeK1ZkvYB5BcTbwdjNd7PHLXbj5j8AfB86BV
P/uVcZGoptr5G/23Zjxhd5S/rjFT8nztkRRE1hihbUsb2unX7VUBmfsl3PNrxY2c
I2rr78y1TIQkgN8KChDaa3S2FkWJQAIlH09qv3cCXIG9DbScqGRezg7cyejTBg2X
Iy4QR1WNWUDrjVoMMv3RWbm9JvUdkfGDlzZqD4NXmW5KqTI7JAyW4ly4i0KFZt9W
1IPkmYpROkZ2N+ewFJI1E4BvuQgl5MgAafgs5rEZBA6EPGeoisQl2wdTwZ9QKY05
gy0LnXANj5UZGT1ShS5i8VELY1q4wOksWWOGOcr44CgutsDLdoaYRJB5XpHA9kQR
YUIN8PJM7FS49uCRG23WvQk9Igzg2j//0FmKFbw18p+NcwhsrgjKVDdZSAbg/ZjU
gshpmQQwVYwg7JJ9AobPiQDXufmzEJz2kcynpkbBgYrutE+lC2JQzK2ZzIEZ1zSU
o/wwSOCZBn51vq+A6WhWsCbdsf/QNTLIvhCjemLz09H14tzCXzFmCUW7UGU8Boqb
dyg2ksnsJro0CeRFATfmku6Pu4CseCOL5t4sslTCV+e4fIo/A/xwqJssFkRhGIrg
fF/JDAb9GAsIa9jt4/rAmrWA+yS7k2TqXA4rT/70D80WRNplN3fG1oVYu49GL65J
D7s+ovCWYRaON3q9ew3Q8ZVHU4g9iIQvCaIAh6pv2RxgMYI7mpDmZchA67N1vECy
yo5aRuptBjWLTo4Mzu3BUrC/P/tXpw58SvF0ARJx2Y7DqwvZjeC6sHrN3lo/SdZx
PCN6OCNqEG09SmY1cfMu0naCGBws0o2A4pLlfpmoF5flinOSnQ8rI2t5E1Jg2VQ+
n/GZQqJ4aRP6gVd5HJbIwDcooH3tMK7Ynhm10G6NCINIR+47LcnoRbJ6LBC40Dp1
NoyhGOn3jHAslaPt89Z8Nb8BR8wXG5qNc94oIVVwZA7GerWRbvLZ9462G42Dg+No
EokzJuwHPNZ8MtV9VFDgVQTHC1FqyEWgWXJnMr+cntM5VervO1EEscfeLZ+u751L
foy3B4O+7hkh3mOGxXwttqGTYtc4L0RqdaB84xagXeirVKtFqPG3G7oeQlLqu4cc
HNH8on1aRHMZZqNXI47LFgTqjl8S06rrkLFm/lvPH+2Y2bk2ldHz+L3+kqQT1CcY
uLGaIcpt7UAVhegcfrPcyVEYQaGWGMvwwru6Fw9Ll5xY/Uhh9DlqplJGlVW2WjFu
niS1wSuFvuwMhgWa2Xdry2+SZs5xCyLWSiRRnDaaYoDNjrePhlFbS0EDrM6QFvOQ
2pWfY1LsnyDOxyQn68GTeNSb0DCAyGKzAHoIAIsYbXfiJKpH7dG4MOkBk7lI054V
Ba6aJRHUYgXqPsjWmUoTFGSn2BSAalweqJyE4T8MjFRDj5JHP77nqMYK6VB1I4Va
lHmyyMYGMO94P16HWSwJq+x4QJFqlip5Gl8scmvKUVOLD8IHQipRxOLrhdriMUEC
RlsUYd9HUfKJgH6PmFY2frqX4vf1XFSq6Ac7Ts8AzqoneE5BMHd4N4CS0Ro+xl8C
HmsqJIb+NmbllkMr+wt57R7luKqild3wW7eqeBbhS+xZi2DlmuvQZAb9tm+tbXKh
whdspXoZvkuDYB+5r8TIsff52ueFfNaDWwlp8f+yKeqIHJWH0WFa2oYjJAl/hwZo
pF5vdZNJOfbfz0Omx3JeqP9ZaeH2+NkOIpVqjQ+lQKvIUFqNcR5Ib+8FGZygSgZ5
Kc+VFvDgb19bUyx7IrkGMu2g6WUJZu/E0Yk0wRsCvZZSG1DqzWZZG35zye85fFP9
gNjEGTGy6VfJFh+V1aQ/YcSDc+cHKjMh1wrZi9xF6xf2hHF8FZ6DR/JJpQKe/5iY
V2Es2blIZX5sXM8sxt4GB4UXn76bax/t1NMt+H40KwgcYIrMr236JcD1NhwSZ/X+
U4wserIvPdiTH4jNyAuILzTtYaqYM1FBoKITiCe0usg=
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 61520 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
/GMbQK29Y+AAYqzOrLs1aWsyBiY+5Tf4mvOc0qXiNaAYrAvkyEOgA9/WXj7hGVA4
XgQg50hTlJetcOlZCZWNDRjNFHQiQelNqVHyjByhEJ9YIjXrbpEWf8HHGIBXbwyg
wpV/UxWKb935aoE/EZyDavfc3QQQp9p+nh0+na4HLstR7r9g9lJ9YNRW0Z67n0Tb
IhHpj2HkyENA9YTRFaSElRkliaJCOScfdHfVPctdn1A7GEjRzIU5xAiucWtGNm5b
vATgiihnHHHqvFhPBjVHwE9yquprvzFtOrJ0whmXuO3Bzfpg0cSyHYlzocR1MbMe
4hhSF6MIl5cQn2roV3tnaJJGvcbaNb6n154f5EKVa6Fz+r1RWpzgOUzApvAFDn6g
lWoCWv9w3e5D0F0WLheT5G8lRPb07UU5aHc8PBzpoLleTgsCJEbNJM1Mh6GCedyO
R02JyjMZqrvrohCAzsItnm45Qcq5o4jnhm/YAQuRuaHTcdgMkKoLJ3YE9veQkacT
tc3qeUoCIh1zS/hlrDhQZ6gZs2oF3LYX96kOmtW9m8LHU3pgiysxYon38s/QqOVj
pF1+5d02NJzGK9KnwJxd65LgYuOqX4SUslh57f6AbXXwcezR3noWyumVO4pB5Nib
uvoEhlKMTPp8exAqX93tIAyEd2tNUcfNp4G71wJogig3natj3zgdOx3C9rcsbzlF
hqpaouYw1wmjLy4PTOSOYzjLy8ELnUB5e4Ap2kpz5huCk0mn2Jvn84r2S1zCGTl3
7Yzs9Wf5/Z+tohv8p3ZXMn7a8Is/ORnmr88JiFbUBu9lTIR6DWtnIcRtTBeYBeLU
1J2CumflXgNgwSt+tf/pBaD4o2G6KVT2pWoJchEYnyYGiDBJ9f3hHsrij5UK7B+f
1gEEeGHwfBugVRYaR8+GofEsU8j0d1gZZIdZ7nq74601SO6nvjeyL0pVQ0QAdcQz
wY00w7tpdgAkZNiVkpTlwiUze23DkpJe0TnPrUkEGWS790NBr03Zt7IeelifKQ61
AJZ+L9DW+Nku0Jh0ZZPOKiuWLuye2r6XMwjdsvoMpcMhrCVq3UC5nVbjqyuWXygz
7QpZ7McNhjz7xOHADjHEr6CsWQmCx2pgqJTq2jvmyWBk9ZOkYFEOiExLIynbdXFe
yl2KP5uwTsUL3LLLVEHikcq6JZeg1aMPtTqBejnHkAJNTc/BJ5E/joQavUFl0/3t
I6ouyI9xuzoLfzc/c/Ttsr/SzywjjZbnTM+aATJ895bRlZ3F/oJIcuUBzWyEOQsO
8ZIvqFXEEf6jBwNNKggqfk8qryyFSV+SzlXQi0aLh8R3L9a4+ArKHP4Gs9nsJrUe
UL+EkTIZih2DDLxW5Ud9rKkewxDp6fn4wforckueSjbcPAoYfTzXgLgJXWx+LX0Y
f9wvYf4qvK2SM4ZEcP3WkdfpUvlM/2GBJTQu3HlRUqPxghGjTsXOjR9gp5YDn7yt
NslT+sqSAbGN99rRWHqZqgz1nBlEVRhGIIPyIEXCAjbUlOGNnK1Wqt4RBgEqFooL
Nk0FyocAW8p94WE6SF0vNhx185y/YRyudY1W9YDSRXk+1qaTnH6W2pue6iACqO26
E38X/GMt8C6vNJgsgSdtUimdzlrZjGIwX7Y+8i7w+YUsFAAXqgRbR/9/siT9cbCW
9dzpJe5yCwNATwSj1zk9gq2okzJzLL1MyUmsjEFB+Y98kG1n3b2BKIbQXygWtmNr
aBMIwQdMZJw3RWMOy3+quIxSOu+07xGxLLclnls2VXPTlCM43SvM77snkSlMcD2p
lRBSvxoLylLLT03BdDybWiVcJf0/jyj6oqrdscWbTAQiOlXWExz/V+yJFZkTe70T
QOspofDFVMtAr6kL9o1lXGLazQCSUBuYwknrSW/pGqlxKyh4uOrelzBF8e4TSuu5
d+NDnhyhT9UCXRJyrPINqulPhTUfgn/LTR7jgru3F2B7ugnqrkd/jDYEu5cSvfpv
T2JgKBlgJC896ciqOwASVy8bJhIMwumaZDpJZ4+Tbbk0vrdjc0HoxrKHbSVQr3Sk
Zj8PDCrTyVD9Q0WanNOz57FQImsB3rGWuwiR2fUnfd/rqqP5VVnrzrtwqosDee3s
vplGladBx0IPqDenOTEmCTAUfXTMBocH1gb9e7YoVNt5mfuZq1AOPj1Rl2grmN/1
Uv54jhQr+mPjtVM8OZ6q/K43HduM8hHln2whNP2PeldEOcoZWFDi98n/PuIfbcmX
/rmabG7K9WmI4aOnTfkrcu5RmynMf0DnWm7opf2s9mcL5opPYA40fa0XQXh06Lf9
UJrz2NHAaYNMRsE3fWFidCmg5R7wF2ZExjk/EDr9Nfd7SiIafQAMC84GCYusdYlz
fKt2N1vXGBsTOUuqZ++YzeoQi2BezWol/3sK+r6qoAIXXk4PCuinvzXJvyHKgloS
+ixbERntv1oNHoM/q/FT/CVPZJje4IXUPmM5CIQJbszOVpdpxBViWkWSdcK7yAsa
5riv2g2FtazzaCqvS9fE4HUEv2T0AzjRJBDroz5pIqEtBd3o+R/BvqtECReDKIYx
XZrIxqXKVsu5xEDiv/dJQSgF4ZbdBVeVwc3zjna8lZjVwrgXbKazsw3bERZGSTzY
KZ2+sBup9WwKwY1cPzM2En/bu0JfDDZLZr79aEfuRX8r5IKNVKCD4Mk2ieFbFETh
Djiet7G8ZZWoTlYaczo2E9rOwXV+k9hvBhJqIBWy5EB9PNnWrQ0HYAuPzWP8VXVk
VvTLE44CP+oqy2kSjqE7tDmn/ygkoyLQp0Sr9OVye1jVNrzaYtXPWpJqskU3/5if
rKln3gRZTBXFw6DRMxyTYCsjD5WXhcT++qzVhW36FVNCWKXNDcGkvbjJ+chW9HQf
oQK/RAWK6O9tzC8KcmdhiBpmco3UmOjbgvwqp7AL26ufXSe1kFCAdjg9CrbEpL9w
8wRkrKUY15OR+CSaBXmm0x9prAmbGtNUSdYDnrHJOE+fc8lvvUcGiC5A85H7e3Cp
1OP0jLuovx7XTCJdD4EXIwgyFzpNSUriPXiYVhjOB7ySHrEjf24gt3KrdxWtQBx4
5+/WT4Xcgb0tKbQr1wlf+FZ4r8KHdG2nOqifnUECgSmkK+JfQGGk3vW+nI9e3wNf
S13eFFGdJXLVHehmA/C62gRIItXYq3TdIOEeyZBiCvfyUQwZc1qXs3OhE8weHh2/
F4sTkKLMpbON+UA9GYLl/rherynl7aKeZLTRGFnYBCG5mk2oxC9k1XwD120d8GJR
rU3Y/ZjbW5GZmAG612dNY2kC/pkwOWzZnq8ZE3HtS9sngcVPS/vRYywILp6BA9ty
/SAQg63aFN9PRyWnTx7FBCKIHr0dXsUseB2aVxRjwArZ6ZFiUeIVmFNy+F2vdZHW
wn/0x/TX4lC9eCnw3a7O8V6OkKpxrq4tgCJ0iQFT+CZ4rV3eITmW9GRKSS1tthQu
wi3rJP0cUwbSGsOYYlTt2MEORWbrmXY++Y2HRQhKWdmzrxg5JbV1zKfM6fr96loD
JMtzifBGRWLe9UoZTPN/4KsN5hZl4SAVkDzdP4XLnKGz5d0d67cJkwPy1nBpjjlt
kcyTOjUxdNTn+Z4BGliWZ+4dsqiS16O45YyHhqerjuuXrvnTyhI2uTMGjKrsXIm1
OBjv2MJpDt0uiaK8zunmGdVcfrGnDW7TBbCJ16hUliw/tXzqykbDZrRNcRYOPe1p
olj8DeSWIhgSBUG+q8RFtrtHgUe9xUsXTydVcAwb7LWF/WmbMC1BLvazsxnuQsCu
Df6pH52JALGGaJxtZvRj5BgUhWN90FdY0wwyRZ1G5y21JOd6zEBjmSjWD3ApUgOo
9GqTykj+BNL0zXjf6a8/mLhsMLFsiyipnF5JjopyoCTXTDy7N8UtjTSBNMZkmZDX
QqiuSqimo8GeVweL+Nqak2X0GOknuUibVkkjvqElKYTfDXPmN0DzyqNmR/vip9+p
A0tW/H2quiUPbzhYAneuu1vUEpStWA0D9PR5whMNiWr7VDmYC4kTpirkw4SH7Btw
NZN7K8NYQRICcfmYDTFU8Cx0eu9ZXYXMP0UF4rfiI4h6hjPIxH+8xR3f0ljUyxng
VuTLiwpxcBdzVXbDZYSjQD+BicIwAg+ZyjjrXciCoBdSsQJxIdA0htoAX2kPmf/h
A3kZcoNapNpT/6Fscgb4RbESGGcryeA3eNNYpb0sl7cZ2kdfXYv0HQDRtbEgwpdT
L/D2RxvVH270oTjoVdOe4VnGDDrJuyCgr79SE6wz07C+SjfAaX1rpGakbs97DIMp
EeAOmlVPwdIfT14nREcZOow3dp6MdZrI6wbe7TuhmBPBkjSa1ZOM9wpVy90fizYZ
xJOULT+CypBOtvo2eX2bx9PBAAHY4IJ7JlYcokTaJ04cx4Mfz08DLzOzCd/TaKTL
Io+TU+QH0hUGH7Rbl61NO2pH+oi6KP194Sr4h7dox/tsVuC8/a/CJ4El0iJE62nG
GDFEAqqwAJJC3FLJU3rTF41ZKUw/M4eSrp2uTNnengB12BjXAjtxO080zJLGsHqz
7QOu5RPJCoG5dJOM1SxnJqC/GdUNCsuvpB5b874CSClOYxwJOPT45XuWLl7it9Eh
dteNsvJIJMPs+LJbQJijEqJ0EXEJNf43tXPkXWHkcurl9sLF9pYNoD2CcipyhHXJ
NuT1WimBt7jbiZeF1dylCSWrLuSrco8d2XIAyO7jl7BN93noh7nXh8GBuDJG13e9
B8GwX15lJnT/cpqqT8wSbpDzGZeDoh4U03PCwJFSy37vHaL3Y9IZZZTI4Zo6KJDU
+Zd9Idxy4LU2p3S5wMWNilgH+ke/ndNGFJVidPpb+TrDTSz6tgNPkAovHjtAnob7
pmsQ7Vl1EAKg2NwDmB3VenKlSN+Ku4G4cO5kpGy5hfDUWbpq9UsXcHLW6lplkS3G
6rnEbVqKs5XzkbUYl7tamHBm4HloYW8E7fgdKktu21sgMXwR2lC6TiEJ3tAbFZow
5rSPR0+IjjBAIzXoRB8ZFOHVLiKLMoC3UH21Ba1iv6xBM5px6/8nnyTJzrLOa6yn
5vsRwFpt/Atd6EHIsNMLhEHnoCagK7uMiqpcczv000vFmE/UYzxZ7fMePxfHuhbk
vOaO+A7DBjjcN2mw3WOQgYQ0C4ZJ2XOH0aEklaJX0+OUpqCn4htCAlKsTvK2TdG/
MkdHBDtmn47GeRNXReEzBmV+/4rg6c8NxOqaHEnPfoHTB1o6sp41ICT0zgJ+vBXc
hfuCmLzNZs6tHcJ0wYJAllJslbgwCV4JhJTx9vAvbEcMmJejYOD72zJe0UU3ulvZ
COsMRWw2vRjjCLkL/rt+9m/7ZD59fXrszwqOszx4MDlazVwxnSvmhBJpFtow6k82
cdKRip5Dj1uRj9h81VVVjZcVrwRBKV37subqQY7QP14Ywtbd5HGFjNf3NnmOXU5g
Lb2IuysZu+6Nzqv5g23nKtO6+F1Tityx/eEoscgxnfeCmcGvuE8tImOoRvVbcNUc
QvsqegVFLOj6uWNbyXsV1ZGxKJK4X1Xo8zkDJfyaPnegf4j36uW7Qg5ifNIqlW3a
JaJd9pcBAcXJSDP2RZG5MShD85qrOqT9PO8G5n7wgeHqIjs0NxQ3brmriMjGMYwD
oZS3Z/WlF6guzxKMene4UYZPJi2bltXpD3qLNiMDQhAkpuKMR2Ja9KMNd7KbnZ0G
riMWsZFLTd7rn+GE3xHoJkx8By9Zj3DdQpybpgs9c4r234Nr/EgyedFv1rQxnzoR
aqxQ+2kSwtoDC/jvBALqpVAs6FjvNYdRk8l/GaYnRiduhn8d2pV2wq9+Cq39ZEzQ
LIdviRSULsgZ8bkbbcypLuI40iL0ysK0ikTvcrmtT6Z3NtukYSSHvr41aWZvsH3s
pWjyW5num7hXG3gtHrJFcX1ImSx5sZPtgt+TxUCM3PmshWhuAWA8+x8bbKa6Akej
dNJtRGcc3vydEYMzen4K/f4Akcf+sspm+S52zFImSmZW4fJ/D3/VymnjsdpSajP5
hMnBReTknXN3KwHQxd3J1KsI+RmnGK+aMqTqUaknTSiOGEvwo+rFElK3AIckGKVw
QPxs6KmMV+iufpim2qAgDSB9QPUFW+tCg5dqDDIQu4waLgjgga7j/ZVsPvWzaqr+
LVTM11hUYUbEGI25nwg3e/mQCTsRoY06FiJ4ssJJX4HGuRgl1sKyVOTlwpjYVTya
Ddk1dblTEi7ofkU/cjR+luYVhkPqZRm39WxMhVPlNNhPZuB4QwbT7+4bLsdL3ee6
0iUGkYxXmtP3kbGmQ5G8aqozYHAP6rv/wHY6QKSxvyWbcaWq6LpJw4LF39RzVHe+
7tzve4SXpLyIx8bYKZb9kXh0fiXfQY1X8nq9kLVzbB/fakVad+ZJOc3XCAwYaR2a
u3B8/oqQlUzBQ48AhJS1I3z4BAtwgLk9mwvTu0Rxn4NLnaqEM+CQcPKXpkZyN2R0
AiA4b8gJu9HxlwZYZ5U/ko5D5+iZQZmFEL+NF2LMTrGtQ6M3Q3dJK3OX57bVFp/C
97H6TK3MJlLZEYYmNeuutebCWIDAIyzb/OMve4zQb3PBje9S1qKW1vJpzlaa3L6t
gVkwZaqS7z+0dE4wIPPVVIXoKVPxYO3+5xcrG865pmhT4d+Ck4YsdvXYXbPLGCN6
Im2OcBB0c9uhLnDdHXyccnd/dKHSO60JD8qNYQbGtEej/tMt0QqyPHBBh/XCanWF
3jWmjcdjMJJfRLytDApxeee/eCkbba8Uol+M8MX6hd8VsTC0yB2U3KygnioZ0GyB
rGNBtNxnLfYUnFoRoitZ9HluR/BkDTLu+FwmUeGIJF/Sp+8zmm049Bp8XS9XtT9w
0osEnv/vuBQ4Px7zD2xQVsY4J/2OLtrIZY1aBhmghekLinqMOIkfTnWMmZ/ognMG
gLiUYr/9/nRUVZ25bTxi2BHvzhoTW6SpR9XB9KVS0X67ch7v5PcCX39/qozckBuH
2XQMyg7r+XPvGZXox6eZx+ft8pefnNqx99Z2N0TvIp70NMei3VIY0UPXKFGln240
gZd8hLaN0+zDHw5pyDLPHqnDzx0HRqKXC2bVKf0KREH46QHjfnvS7lBH/8I5tP+W
xD020iLr8P0hn25e+zpSAM6KuFJ/ylqfEmnjznEHdvGF+x7YIHSOb0WNsHjnJzlK
PJX0M4rgEFkeAFtvs/JX0XaVfNXkbq/A1hr7DHwL2FuiwUFVemDM1Do+Bmy6VkA6
tETDVQxBgMLNdVEwNwta0SM4nYfTvfGhOZdpqv2yo6Qiru6wFczVjunKlk8Y2ckK
SsjMGECFwzGNEf6PLJhtCiJTbx6iCDv6sqdXhUqmBJj/TASHO6xjcE6CzL+JeYCe
vWRJtBc9V2EuN9O5roTAItuhK50uqIdXHYWFaEhC/yM0vS4UPExPToZgRmjTTb+M
/agJ/M+Jk6jZQLnu5XJ+hZV4D+msSQnvyK7FelA6ScgcI/IeIGiqrOUS8ukd5dTA
ADEISdlbgH5VUdqBPVsqLq4JtzmCEksxBr3uGScvfkRmdw0u0b5rtXz1b3khK11a
MQEVX82Z3UDaictGada2ghh85Ap+GRDD3w+OjmLqci1LzAsProV/KA3Bfu2KsG6G
9usgLhx78vIesUkiJOkF8APHKvmbD5nHVuyU/kF6SKgMPfpBXyhOsDVCZQDCIYoq
/tG1iixuct+cPveXfGGFhuPAMaWjHEk7S0NjE74mR25M6sen/rh0UOmpopLwGP4g
2vdZEDhOrMFK6cZvI8DnlApV2sYfGvLbtdFBg2RR29UZlrkbmUpnF5jQ+qyQXS0L
r/BDmHd44oneCQ2cwu7siDMr3gH89ahyokQ+aSi72KJ9Wduy8uYz1hVkwgkwDZc7
Ydnq+w33hn93RIVRMsuQTS5VlR3Gw5/4xbwUM530KCMTU8FuUrzLs1MFNTYkwGqV
6+4E+MK8nFhk2MeqJWGaSAuVR+nMt3ug+FhIN8qPWNf/sdDobpFhfSMZfCVwU1Ow
JFa5zecLRz4miD/V+MkrfsXFy+1aTDeXnZ5Q8TEs8N9WMBXDbedsF3mZ8xlrxzSx
NSKtBHonmYzux9baeGKPeXdUmV0wHIDiJB8fgRqnzhIFjrIDJetFra6Rcg2mGN1F
gRDA74Fd9fGmoNJqm4vlkIahWFFbD+UAl2TxZP8pBm3olhrteOVUnyK7gHiwWsNJ
wFypFz4dgnMm8q52vekdFeOnpxBx4z+DgsQSmRaLFTObrfS93Zqwl0nKMMhVPixy
isLVUtt6uV6u2TGttZonykurOMd+2TASrdXuasIlhgrXY5u79uJ1Ax0Jy7SvpQ3b
KQ92wGKgwPGWC911jCGjN7c+DH69MsaKNobjXEJAhOOZP70p9J8sMdUnBMWDnOfg
MfpoG/ccoKzAZdUmRrwiDiU6/eV1Om9rTVW8OWZqLSOH7n3OhR5T5LZQdivWywdK
aw8lARObn7Qez+44omKGFLcugOxCztmUJofV+/iSbBo2SZDN2aVkrIK7W6ZhpLx6
6ovfJePNkAv//jcM7t5zJ7vIe1mbqm0+9/iiMglv1njhRHDeXZrGWMm9xHn6umQF
F4EuoS2DWIXnlaCcCYxA6awThEVydxueGhKtFED4obeozMh5EEf9MUyCsikKu24A
GdLPh3YRIOM5rDGEalja4yoCzHyaW34S4BN1lp6+8YwUyAbW+9fAh5fTJSl4mN6l
JERNrNNJQGiPlpuPMVjuSG6Ljv4qx7rrsTMEhIdmS4L4YZXcOH3/B4KYbLDEx/Sf
VUaupgWRiy2GAQbmEuzbawLu0NdZhTD0xglDMc8Uh0jsd4evEySF+xT6YTSut9B+
3AgnTMyTafdORjqoF66nbhgcctcwJrvbadQdFps4nlGq02G4zZHEC3eRkAFRUXnb
Djhk/BqCGGq8CCale57+3eeJg/Kfcb6Ob2k0Mt+9+D9LMAjdap9UrEZTShcu8NU3
5Rqb4gIAYC5mkYX6Z4ZeImYfLq+sSLSk1PxEoeWEQQy2MH19oeEvnF0VMbUd11bT
eC6c2YwKiH95xL0QB18UBBJxR6xxyeQe8ajqxUB0Z/1gR7J0iFrMrVnHQM1Jka7f
EJxB67ESxoq8/XfNxTx1OJQ2RFtQ8X+1xWXKasoFd8ubnL34XbF8p8OlahFAR+ix
AhWWTW5R99u1+7ROYeGmST63OZagg0to2qgP72Yq5CY8i1+7NEG2jUGJuDctICK+
1DtyxeuCxqvbeg7XFeaJaI3rsuX8OCZQ6HXZ7p8/VrWitvuwc3NIn8DmcS4XqYWp
fA6m7ZeEpV0DeyrRAR5dsSP3uAraPtVfQ+rkMsk2oy5HCMRfwRS3u4YdQDxReopc
bqD9fU8j6SMQoDwvQ1wSZ0L4FvVegDHFv5owImN0c6cTS6HMGMd5h86PA3EVbaZL
z7V1fuQS0k7kdchE4tmiwtfVs8QVA54pBDL5A6dwR9zSs//MOSHjUGvWvutIBQXP
AzQl8m+1gysDeGsqGkGFaKQhPDpYRbW8B1fhBFQ8SSovgOxz/qbbgx/CeHC5qcnp
8dHP4dB2kUj3LBa9zNtMtuntXofz+mDcAruiMSyZ3hGb24j28fiii8IWBYf89Q0O
IbHIJL4eQgT1dsEklGj/9GmmxpAIk3t/ktTl5GwSrJgvd2sVvrWHJKu90Yuutq53
D0JMO91OQSmLgMHRE6zohqb8B/CBMl33EO8UTadFAXg+abaTDcLb+4AJWXKgODlP
Lxxw944XEuAF7ue3fIA5eAYJtJVX0yqiOjlblaWTI4RRMDEEZSQXrtO2JucTnlHa
8edAhgHRbM1VSnVaDcIOF+2wJaHF3Dg3hp7nE4FNWaDj4i8FRR/9RlL9xDaOpiiQ
3c3WCyTXlF48ly0OmRSeSCMdYOO9FpAxvzRZMadSgIlrjAMksQ4tfOPHYPUdDBze
Jqc9WaC5UfvI5tGgwN24rRHHYtEJQwEBt+QOvNUL8bTuagbJ4JQMbRjs93MstKxX
4QP96gF6aRGediLvPDmvsX7tRUD6T1PTfsMpNop/hIz/gVs6G99yLf4/t0j5Sh7o
kESii3JlcDgVidF/xquMvYg6fptLSE8cJAZ/KHKHzG8pUWLVYELd5DlzWcdrVfGV
+zRDJsVAD3ajt+x9MU9rSEdG+UxFvyX7koO0rIQvXyk3Ytt0KRtVuSSJ+E1pBi84
7uPl4R+sCaptZVcABd/XC3G4M3J0WdcQCHlfK9NCBJE04qMvMv/YPjW5BFd8br5h
ECLCxnKfjV9QkvVkmrWOwYUD0hMFsbmETO541VmkJVPCpfZt/kKLYKKEcEH1/03A
Sbx5vS1Xup5IKl586/yIT+GMUpeZPPOfBWeQbv2z3mdIwliENKCuGckLySye19k4
CgNYGDcYRoKqZQB34Kk+X08rMU7bBoTGEAipKQxJUwA9PvSGWmPojOM/phOceKCS
KxNst8Ns0f/Z338hUwu9FV1cOW1Jctd6hbprpik2SejKuQYgG0SDrHhOqL7pRLLS
ozf2nyBNK+xl9K5AdlxBZosm/KYsqXsvQeIdMQ8IiA4edk0pj9ccjac3ZKk9UKjd
+gTy60n2Uf3f8jtoxiReoeGZzUorM8C2syM/jt5cf4d17BR8dt5IzVnz7bVpbvdG
sS8lj8jFUrxL0NAJ7YdLBfFbDIY+LvRueVGHvlJv4mn66iszeKOI+EG5kRT8ko7N
24iF5BpCD3B2Q2PjQ1QH8RCYFCemxPZA/f0ExDRu8TMaUvfslVHBPckdPD+IKXbK
YxsCnOxNL9xs90zA7os04TQim1JwHgwJlrPF8pvoFvk3oDJzxvosip2Pms9b+duN
qXygX414fKkLJ/kjMk3vlosFjTuLKAiTtxZyEvQfOVIrV0xoQbKxksjHdumj6OPJ
wGAwKAHqNZm7Elu1yoyJeNcQ+ocooGfegL3UVBPqSlnxDUo7jQ5YTLNT1GYCNois
Bb2btteoT0IEPZM9FuCPM/6XToVpoJ04/1pgOvO5h3kO0lta7PoZZSYH21OhlbkJ
7M2IyR6UJEU9fNwlaSAxrHBsuEtek24S9hNquyp24P+jVJKibszOgGdgEYcijTGw
Lqn+mJLoJXtfwL9HZGg0XGDAcwwzy7h7EzhAMfv0RXKTZzS2T5xnhxt//ubDQe4e
k10EhmWoYL4sHDSHgG4zvFNnEv6eGr3MUvlozv5FdvGBeYSMC12ANkmYs7USHUy9
rUldfEc+q3K2IS/J9o6y9YpVL74lXIco4a1Xf3HabuOWXCalA12pFi1WBTy0CQDr
+vZl6OJjbHrL0phC1EQf19a+3k51JkYQqilz/gAU/9PSqDI2zJnc6lUFKqVEbElZ
DZNnIRb3cc25klAoNCTZFDUxWUgFMyQUrEiDeOr0qWGiV8yBMpM9JmQKjKIAXJXl
r+yLFbgiPB2GlN1KvYQVbgFggYI7vCBowYa4D+IRMW2fpkNJYKRkZdt4eYxBW6d4
Q+irx8dCRccnORSPMM8pN21/3izDKFXCbqsbxv2rWaBDiTMMD6tXk+bb/oC9DzBZ
8GGmm/6imztrB35zy+PVywGTSG+Fl6EllNMWsQOLodCsxNaMU2aV7VAnryG3C9hV
qoxrSnu1BS0++wQpib18MSGfDuZSAs1Gihg0kKoXeT+zEKzPdsglVowamgA+hpUO
iD0AmrFVHa1uel7XP2PeaKU72RDnMfLAk3FkDewwo+DW7jbih9TLUgJS6ovlwhPk
Qze6ZCHaysR2EA6Cnj6kRd+BWkpTzUeU9yl/a7PGnPX/onNLRwbtmKZLNb5UD8eT
K2J1X2qeeZUHxydnE4VKGY3mOgQUXn+PfmVCsVKourguU/+D+H1Cgj8BtXGcyiXK
+e88HVEXaFlz6BXmwestJAaPZ2nPSXDqdHSOt58KiHS08rNyrUftVrT3XrkLmaqn
KivjXx4cVO0gihwZ05QXF+Ynt5y01y2/ZAk8BzYyVrSsgEdamdIQOYbWmJ5y+kHF
BigaEmjSvcjPxlD/mr9pwaWIT3qYqAN5saFCo2Y6khqco1C7q38ks36fG1/302kt
OuiE0bRM013yCvwQuD7PnI1lewkqCZ4T4SbkIGW/IIs+XWIM26ehtjqadv/7t0Bw
hUK6kaX8QBFch17CNFCqg7FYCdFJySt/71z/g0uKV+esR0b+Dj8DNs7HdswabcMA
z062TNAXOI5JZe8aV9DLg1F60okx84DG3vqd7o0fefiyfOB47iPBnnvGrTZC7zem
ZomAf+uGI2vSI78sr3voUvBs0GZhQrKYgsor+vZaEONjQQlDg9GTENILSYz0nwFY
SdT2TTnFWkB3KqGeSmeRPnHOqcejLABwBNwCsvWDbPPfAOJPM8dwdCLcb0S1Q9uV
24chk/cedfGOL1xXnfkqUhfBLnPcbzeeZt2WOIyB99WYBL5tEIKWcN9RQ94ZOrIP
LhGS0Pg3jJ0nelQKA+wjbP8yGfBzvRjQC1VC6xz13M74K7eqguo4UdP4URYVeIo7
guZz+pvNaKcZTnNj7auSWtd/1eg2gA6NS7J6ddqG1w1iVJpBvHlxkLVupaQQnQwr
hfvPSJz/fiMiaXcY7YJiqEy9xUM0IftTD+GBX4lPby8mXEpZ3qb/VVeG8ZByK+uf
eEovzc0aj0dwPw7LksJ4w9Kn5BcPk995xrSyhJfmpr+rIWj2Jz33xC1o7ubJz01G
l0/SchGTIMAsjKdJ5m1pkwfCTHNdx0q4LeZAi2IWV6Z8QEdlwqP81TUBK3CmYTow
Ubbd+SuR0rPdx94nO1Owc91qUzcnHu8LdXTzCX/XOVygAluakj7Nb1UIysymIqX1
Cj/Wyy56cLR31mwUHNumQB50bRAM01u117/C4GnZZeXNSZZ5+HNibKtptikh/4FO
58f8K3tFuXZIBNDZmxz41mx/kMLZglzftVccypaEND4N6AQTMd1/ECfqgSrHaoxS
lkDubPi+cl76litnJdqQsBSFB7dRbX41vxaOH7lnuIjyF6BDGJepLpQfob6wFJ8D
D0ohTCN7inVnJHo51BKKrWy5QEHRZYhIb/VCoB7wh0rshopmtgOCF17Z9A/oZIEW
ZTc8UAPi0iL1SLdvUHQiVMWldiQcswIn3fnxkEGE3rXAXq4LewcsPr/P1wy2R1Wf
N6zZUAh8vgtjt2le/5RO3XLFUsr5b753QN6yN9QDaq2DywFZg2kmD9pkCsJiiEx6
Dqgt5U/6VY/oNDgIZ2k5kHDiSr+T0olnNxyomkQxwOXq+kUNhymfg0rnqMiNzpRP
dtJTilSaB14wLpDiCMQHspAPdu6316bAiNopq0GVM/zYGog2GeL1xbNA0slqJ6IM
iqZReTLv/thz/aQoXG51AttrH/85lIqPvp2ex1ASAFeaFXo4nJ/xHcw9RiO+mT3l
+tld9DOTVk2+N83OTHiPgt1p0kzY3ZzBLdjd0h7NXTwHTIvaG7wsIxKwY9W/4707
FyHweMaY960FTgNSs+ZdBdaK+c5/xtECdJ0hMs2tIFYqa3WTgOvPz2SBEdYqN3Un
tNfgbpaMUZuN0O6W7IR7udaF9n9ZpgL9NnlmrRD+T/MWEcEQsKUt0VRi565/LMgV
btPorhgFdgyOo3KlCcUBE75b3ev8nKYxdQuuzqODJhGBgR/nxwoM0rZB95BEjbjR
4Smm+02v1F7sqokfayIfDAyKByIi0L1bDd01AJnTqTs3sUgG5fr+MeKjPUOLNXr5
XUgOJpqj9tjUZiRyQiVrmLeMN61IMtaWbTdrR/intvZgFo44JFSRZHUY36sOxBXB
/62LzYhdf54HQs+3HKMQcNIE74AKaalAsM0Sw+vSpLripedy62tOhZzjjN13fBKP
l5IFvtV1p6lPfrcJ2O+ucix8KYMwlljz4gfaaVYaVm8rEzeXcJGMGpi02UrJWkhL
LW20ZKriGZUEvzL8gUruMAxzASRiiOBTirqpQ4ys+6Ra5547sKOsQtjpeQ86ulgd
Hh7Y6Rqt56PMVzBu9FGU0tLNkJCav1HSnGgpBJNUlAwRJVbPU2T0hb8FC2KiUGP0
Bj25QCINJggQFXuiiGAgDzODYPCXY+HkhsqREiPW5Mh1L9f29s0rSHrLvxt5DORR
/H4a1vBoe9BqwjdH9ASu7cmfxjt9c28K4rIRji36yjafIRSllpxMxfM9c7szRpaJ
b35k2f9LryS43B1+RdyLrjEu79mBIm9mgwFVquiHh7Txf3TXkWdqUqFrN8DH3ExS
QLUSnTCAl/WzoQjNiDgK9b3+0FsfanTYuiDsZY2LXdbDbOa49qF1yV+4BQNNS+zK
6qxlE3idoyKh5F+d9b0g4cvFeuY02Lw9SUNT8uK1t3wKCz50tP38r8MrbeQW/RRi
Agtu2/ys+bGO70OhAyWd1pNrWoGOu6Bf2B5NR4ZZYiQmssXhehMgEUbD/cY2F9i/
DbMtE2bVmQ7qD8tEm1b2xQw7dJhhEYHrDxFHgvbWQpLg9GUprK+dVn8DlrNIFWx6
uk5tDpKUepX0TcDhG/YAq07DXPy3az8dsf6WfzhPZfe4/swz3vXO44wVIS4wcJpD
z6gGThAzHtSRMWkEd/mt1ecgPd49d4EER0JRe3Gu/l1myZlnHfb5MgTxsj82+tkg
bgBTzNOy2TikSFBCrlxoUfLkjSYx8WMHKyichIkp4xqvDv6izN6Ytbj9efz2FqSV
LisD2w2fNr0zzaN2g2GmoBpaGMJVo1zHuWDoThRC0vQv1SothiQT+/fV6CxPRpl4
Xf60har5GG9/DRIh5G0kVZuBUYyZzA3yKbYYY9ryHTMoClekzhxUJuhqdIrVUdz4
ztVtjNOwFg1HMAK2i57f23Rkr3tH3fZj0AbzlDpuOislNji8L4j93wNIjf/qrRGS
PpQo5x+4uaA5tquad8lKFZE0/TDr0hxtTfdJC1fadJwxkT5obx/GhuQxnr2DIuRN
+4/XP2r9cu4D9IcJU05DmZ3JrUjiOZ5mN/tzy7EW7/vgAUN5Ckhadnz30+ORVMml
3KMzlE30Qkv9Gy0vMtxbpBfHs3/wBhYmTpVarp2fEO9wvAt8Xla/BV8YHp73cTts
AwyBQ0xEtDo2tPd0gVEFiUjsfGvnjDuqt0k4aYOL2BbbzBZSDpdrbVXDVyJuDpNp
V4P8s6z73Iyexl1CvvJ1IiYAIJFEqZoeVxBNOLRU6PFdkQERI7Ct1fJZPIQCqP3c
wAfFCG6V9J7eQQ3kL7sv8YAz0JUfWvJ0xgoKaKRK4uPcVIWoLZfwTIplBza0B9QE
dohZErwwIE0SqhwLzv84ThwHv35KJXPEoceD+arJPhC2llYwEuMfDibhNneZ49Rx
aIaPvT5xQ8Ozg4Lvrx/s+Ph4XUCBDrKZt2PKZz2xpm7JmwsYlwFC4tqDhPnuJ07R
ze7TdFZVlA+MAm57oXjkIvtoMKBao6HKF4yKkUjBNmVd66E3/fFRCujBTcz4SBYo
pqDuMDKjY5Qwvy4mhsyZLH2Y2KQv1g1jzmTTRZQQxoWDTThdx+sinYD/lOoL1u02
0k9wS6EmK0UY254DHrgmTRbyDwMIkKvq2bKL0IAWX3cpFA/f5Wu8uY8QzjCb0fxf
Ezl4doy68c7ZRQuQMSzjoLCmP76Y3EN51vPck5liqHAdUarfRceJAXiQ2p88sJs3
IN4vquFFkctBAqEsFAXMs0Rsd74hvW9igoUpStQdnDvS5rKNH8zxNdOA4alObixC
+FOhNj7Y1eY3mLpUu7vDCQoGq6LftomtvqRoG3gR9HVCiE6CxEeV39kwUt2440en
RSXgUGKuIQdzv0okXd98cyqfHrzg6OWNhbZdLf0OxVtFuNeda9QBZhhxxM63jJeu
KW7QDiUbJ1h8zFJgBWwKzuAPkhBAZdY/7SFrR/3QmaktyjyPKKOb+UB7W5grkqk9
paY2aToVEiYykhaPXnEG3ZLDGPP0Cra2lVZrGfqU+h6IBzghq9gxCAT02u1MClbH
pIwW4pczGH4F6Y3yKwh/+fFcQbOJDbRH7e6OrJ1rH35J4iS4lm+XsiqEf4648GNI
EiGkV8wuEI423WdwH8luBPfe1i0pwvIDcB8T+sxd3Dorh3WobIKswDEzHFi3Rrsw
Dg9kyC/dFYbRXszZzgANnH05Gyxx0gTfBKnIOzFWNhkTS+mtV7E1OfJmTpept3l6
0EicMsregj7aKX0SPzwQrjwpOnJX3wbR1nDOvYBu/Lx5/mtnOW9SQwTUrPql704D
aEOxW9wNPWJgVuZUiQlQcSkEI/0OJtZn+FkxSLDdXhu5Yy4kUvkZyGI2RYF1s1FO
XPD3ubZVtO/jZ4zxDJ8w0OJcYedOFkeC1bJlbnkmadSrNBUh1vsLYvckhjeqJGKk
xI/XSEBDs22L25uv7e1Ka5IZPeW/JSi30cFUCaaSgqpGZXV1Sgcxm101mS4rc2ci
N4t5VBDGnc8TN5SfAgZ1lJDaO7tbARqwgvZngESO3+rOekR2uwZ6AwJmPK41ApQz
BEUjgOLBT7yUxP0N6nUDubvFVbHGdKDA3lvdnb2LICZmpaXG08tpXJq7GBNo9K1s
ihlIxtIpd7OzkcfDxzcvFJd0u+anCywQEDijflaExdJ8JRH3ussjDDt89yyu+br9
cnNfL/JbDSfh1bTlpPK+3+SdHGcznrgoekGwsHTbm/bfdHxEXBjnAT8WQWQkfW4H
SvKBrIsl0/zsDk5bAZNW0rzUcVZi/+SikzOUYMtGyj3gybWorXlolqkE00FjQyRG
xZ6p7W500NYvfkW7prPGFYZ8pOJOrV6Qf8cdHfqb+MGCXt0Qy5jOCpj3zKLQvYVA
sRqCNE+U2ZEqcBoDzvQyva0QHwfexf5ySwiehhv99qyqxIqVa1tJNaZiYsMfyFim
6WC1X+8qzqgTe6OGTVS+8ugyy3jrij2R+G7LShSsu2hptkXbVGnRT12H8Wurm2iR
Go37DqcA65RmduH92XbltV8g98faClIK8yhdXUlTCkBf17BLVrY/Lu+dfDFIKmuW
vGwvBtCFrbdgHGFXwVZ84uq78vTgZf7hN7+epIEfAjyRWp8kbpaojCEfr+UzUezT
o1/ej6i+0D5850gDwozMyv018x6KCshFPGxYc1lbK9gOTbx4/fsq99iEl4Sxgp75
sXktXwhnhOoyUCbS2J6+C8snY1ItTkk32zwnilzFqy6VymoQsp+EcVCcCtFjsc1L
UuKrKwjnUhiu5KXoZ/l/pZr5uuHarTLpXS3Aq+WepqtHPPIz8qxBgbB/z+mH6s3h
ZRykaEYG7jMtYEf4w+rpzIKRLhcurcdiEBuvnvmICxr3jeDqmWyQQHxND0dz9CrK
GALb/ULSGhJRdcjq7lkst3VNUmmzpDycyyykrRrTtJ9nV4DZoz4Yjv/296FPoaLR
P0xwdAhq5sdHCul3BQHFYl6Wrh1AIAXiMHFJMWpFTjUECVgjSHJlC8oeZP2q2kYh
Zp3FRHTIJnJlwpMlTTCcClIluNgGsKbpQ3dXCzNfVWLxx8dpYHswk2yznSyuVDb+
R0/akG0HZOursMqbSgvlkuiwBdScBt2qfgaLcAMwz69c4MChHO3s6GRGSFH8vjx/
uzA8O36fmovQMuPFPiyA10aJOT/cgGOhkAcH9Yw4LlQbqPMDxWD1H7VwRpL1bTq7
jnkjOImp4qH+X9iO+CBFgX2nBVJyJ2kzsLCN5ic61UHMfvjrY0OJtKZQYM2R90we
pWDp8fibzvnIqHCzq8uiK5HgzOItiqyRicIEWhKLS90uIX1PGOoL/3ODPdKxRh6i
KJJr7Dmsj2u09bqB2LSiu+TLRHpG5myGe+jfVg7rgvnxLgbSb9p0ElQ2XWFxdDHZ
8D1gRm5b2lVHndiABMf2tAzI9EpwRYBxcRYUw9Yi6159SLKI59aIUIQXXrVTXhI/
jqFOmkVk7JG8EGPN6vyHiuytM8vpup1fD7tc0TU8J15cmcxAFrcsBu7JTK51YdiS
TEIJQZl/UqJKpMXCMh82+ad+pJbflpgo25Az48Hu+PaGwFR2xS7MH0MBjZjA1Fvp
HdbyeiXXFus9AnYPZy8Yc0EYHQwmzunblVTJ70GK01iKcqxJc9Kl5dFC3Y5Fz84+
s8suH7ZZyC0ueX99zzD+2y3WdGrEMZKEKv/Dvq8SUoA2Zoa8eCCGTPIEDLfm8XBT
Xmk/iKU40x/YeNjvRIrEsIINQgLFaGHEgKaw05U3XtcDBOw+kGyEOYTrbAIXN2ZD
HZEFh9yWJ8FlaoztwbjMbJcm1uWaxucSn7E8T1leKb8OizBj+k4WYDXXDqBYLrOU
kGdohzrjJ9frAc1IL0J8GPpH72sFCMqRWtZrImhIhxEoO7KbmVK1MDl7y/wSDqYl
N4tW6bL688CXpTxH/0z+2hrvJebhE6D3JAsrtZUCdPad0WE5Sfh+x6fGmBejGdM7
2I8sm+dI3mYL0eC7jm8wvBf7sk04yvi3JIIUT5cFVwX1QHkl7LBxFDaC3geu+W8q
CDHrm7l+FsYptvi4UuCUzEmk7rfEaefiAIPVChU4258DlAXoJ96uTaLOafUI1n89
q2QkdBLFVqmLsewFC5UjlZzZYqWFOb8djQ6ZdfBTfE95fHIn3sXV4KDkhJOdYXUR
nKzk50YXDMr/IVv26IvjUNFaGLnmpQ3uSZ+n751yhIad/RJyNnTY2OJ7SEizcxMl
8G5AfnYwsqfOHlXl86JDoW4h16kllXRJbMUrN94p2f1e9e2JutGMCThu+hXYrfU5
dtL7TyktsS7NlEc6QOTnBvoXh2dYth9njU8X4lr6Yjd1UC/pGKAJd8SHxZGYT9LN
9TcGxmf65EkmJPZDfPOWm47XeNKtseK+US9Dt3LR/+/NzNPFM35EhsQa6fcKf43q
PqZ1pcIIGk8ye1d1oSaq3Cp01YXlEyq7KSXyzqAC4mPe6aON4Ijeb/07CeIsiPwL
sa6F2AqM3dFul0CCF63eVztrl4+Rm92K54q6rvtyghEKvvL+a69TxnUF4m0aB/l9
O3etY9HG5gTgoUQXs+ySKdnYe/8KeGZ241UTj+bPFH9OzXHO/HtCVPuzoOx+Miyc
D/zi2FwoydhClahaQnRl6VDcrRvu3l99nzI3I3KNiI2/Bmzd7OPLA67q7yCiWzdu
RZaKh8XSRoRayX5mu5EsnjqodNMxAA9Se8pvw5EJ5VMrAz4SiEAhP9PyfPGzfWaB
ZvGqwiJbafIV6z2Acj5yA5iWICeV2/PLg7LnSU9z3QDQPy8TDwZH73cGqvBnOpPq
PXCPxjYFaha6PoEG04zNeVESa2ztgnz8ca7hHMOba39A/ltSjTWvERhHkB60cx2l
o+HzjC5DhUepq6OXBmDvV4bWI7+8V9+0CSpjABC9g6cKhQv3P3TXLc05ybmT5e0c
e0xlwpaa5NMobap3eTnq3AdpPXJfzWf+7w2RnBDNWGKSCTC12b+366FFuqj8Z2S5
Oj32WVolN75HGpIuuwa3AZMItQB2RtlaT+JMSwPbCxdO+nmWr+m9B5lWlCf61k3C
6vbQS+79klTO4wJHgkStksXHussC09hphfnz8D5UYsQ4jUPyRCpj6HhVJB4cb3RV
k7mNPdXhgZWc5e4hTHgnz0uMRQqIdvgvI6e8O1YF5puYa2dz2wJRxZ727rBLAjeh
Q0ExSfC65BiYR1tUg3C29lWw/7mOHc9KDOR4mrv8z1Ih6kg/0m3yHLPpznMPyFVF
nhUQYM9XOPmPTFGyq2S1nh/4uww5YrQg9MFI/+s6I3+C9aIiryllcsMXQ0/rLuMl
fuH5n9gVzXMqDHprzJ/nmn/Rjox7h9MTvHDv/J+0nGz1rtqpAroaVDDiy8BF+mMU
NWERZ510duaO2crDBwy4nC4qPnkuJgtj7rqj9NQmPXQ8/1jnJrekCy2FjUgn0/Of
wl7QW2isdzGYemZu+6TGOom9X6hWsOhnqs+ZQ/nACl7SUDAn/DfXbqsgt82Qum/Q
HCpj0VltYNxvzQFGjDvtcSrqXA6L/kEIqKESystLFo95FJBxYKTWGJiFpTT+PouG
mRBSGQOO+qc+4uzURyzGBV89rwLt0YWs7ISn1YUDzFitEIjy6xGQUxld8ILE1BO1
jHmlRBF/fg3PkIHhJ30kC7NO3i/g7p1o2R2htneRoSZI/8Pvct9jv6JknOzt3eif
NLWTML+zGCYaHXuAkQG3JYeZolJ+fZRFBFM1EURmaQcahmBl7cbSGt6K73943GH9
arQlMzBwOd032j9IzJKV2q+THiSPIUg85Ur3Uzx/ZX7r8YtwIVcmfKSf2dHi97py
Xvu6ua42LvLfsm6H5COg3pk0s3jjHe41NCrtuyLgbGtkykHHEzGQQrA8YCQ1k76U
6bI1ND8/W+mtZCJQxJ2CdTomy1379bZjBaTEBdtL5KOvAi0nEUsRs5a8tkI3JaC1
Wuqp0YCtjo1B/kTmz/I4SRFDcoUciTswWexYVMl6Z42Ao+hrh+RLhJJU0t3hJXxj
T/YfkG/Mo4AfpF3/Xu0jXj2cIX3CMYNUzde8opR8fV+ojT+QoiE30cwOoOTuCzCW
ZVzMivwP/Vr6k59WoPyS0rBhKXerWoHc2HcDe2xwQWoyl++Hg3qvFLDCNRSEkEGV
5JAWC1YCH6lPnqkyek3nq5xtzvrBhopJXidM6kujk/dEYRU6hZ6drpTC+fYTV1TW
CBPoAIfjJJKgrFMPUQqeADog5hyCqpSNKE8XkU/KCWxfSo9uNFd23bx7fo8VY+Q8
F6Dysbfd6cmzBHz5HWBXyMzybgVgsZptppofoSyOwSzOFLwCoggtzciWYrpKpyxG
KZqwodVxw5HppH2hy76R4U9ZTbAaXakau3LnXssAOvPUCa3zuyJNJJhDw9Z0xTWW
gLiEqIc4TA75dSmQFqPCan9acgqvPNJs6HQBUdAZtRCzaS3dihS58Oo5Hkmxa9so
sd7Bs7cLrRCSu3/VBE8tAfUpxCoBSojwt4hrILGFAF+RNeH8jdC+Bi3O025A5ROt
OKC819bm4g41cXVdXG8lK3z7vquECqrMoHyENr5TszJDnIXrohECoMq/JSYaSSux
rRtHFfAT2FK3ZJw1eGkf0D9afHGJmhPCGFZoQEAfIwH1zydezJvaFLyJ0prfTwv0
WasxofyvfGPdrrm4eZ7kvhHCePIwFNdDGSvH/LgM5txV25Zia2Dj9lSsckhRLZj9
4WeO1P9+5Hlx3iwGCamuEBPdABCeCbu2MwBkW3eamuh/BGqIYwMYyBlP+UrBG4gM
4kmpdbWUNFwUgApPjFONUinYJNhn3BjvqcEcZzUlUT4ZpzOjVkeghE3+hFVCf/Ni
aTNfA3arV6aRQojY0wInGQIiZ1fo1sKO40LFFB2AD425uXDrxD0NEBQ1S1SRfQAF
rp/H+2Sjfdp+hSRLShJEqPLSg8GOR61UoANY4VlCl+F+q922wk60q/ZJFdiY+F7W
PFS3Tp1Py4czeUUMFAibLoAhvRXHt6Y0I452dpmpO+v1Ns9DA+HVvHW0PSsbWoVN
cvHtyyrmJzfCPPCm4zykcEpJfFKcTvF0+F/6k+eI3e0j5d1fnTHPBhKRWyhxBde0
W9HyXinGKXX6hPiFru4z+m+o1lZn3N8DJ72PwQ2qrpdvBnPvT6fWqG1lXyL+4+AM
EyztUyRTMsPB3y8F7pVgZFJX+Br+wWzB0qRjSOU7duihEx4LI2fci1MAYd1vpJGp
KFriQYu2YRxQWTeZYG/Skj4zzrmCf0x3nYVC6plQ6TY2lr/qsZ9yx3f3mky/D5+Y
fARqqAJAum/JgSlzcMj8YTPVnXI0Q9OjAAvLTdURUBg/VUx9IfjbfnxHO4dBsJLi
y+nkz9mUh635PtrqIDNKe77ZOuCYycwnU8snlAFCS/wN3AluXbTJDHfPLrv7sfyo
09/6VgFaxJOS9K3Q+siYakToWc/D862uFZqXWbfG0UwwZqaLTjtjhVTIl4gj6Lp6
IcOgEitaxczikvcIlXm7+LVMuUakapoTVpAwDOLWU03+bl3nybuEwQASM/n9sAGU
827gtn8FA7OcJKTLaeR2ToPScm6CdF3EDYI1ufT1n7BaQPCs6kWk/77WSl0a403s
q83sac0+Shb1roipIWpmG1AxkH6X60dumdd3PWxzzN1DK+aPhNv8TuGtwotmKE9k
0K0U3uOeB8i1qdQ/z9rrFRLFVLTAU5WPZldWBtmZ5TOpGIlvlmrIrtoRYdOSiPIZ
vRwXvMeY1yioRHCM9vODYOMmZVxcnTOjGvbklj0ayDLvSMl0fayRWpF1Z2HKBBIA
ZJZSaI9hIWk/7yq3+y3z6lNnXVtZDmfjnihHeRQhWONbPJKAYMmx6tCaYA/pjR1q
ymq62R2xzWAv/mDBYWPrvv8FO/iVtAufOPhorqeEyWRDio9IM8c2EkR9YSDDymla
EZAZr/DjwwLUQPwbe5SwvJqtcy4iXoRfkZ4zk/e1m/TeARCgZEuK5xKf+wseignM
ZilunTqU7XPrhIZlcJXvoVmEeJJk5ZhC8ASm/7SMrmbhx7AEnuYWu2sDRZ4gdn4z
nuRqG+l/BiuxJMKiQZoZT8HV0HUolPNh03iqRoS56zDUkxs4UXAn0Kgx4mQUf6f+
feb277ZjnJaJTPxWPUmZLyOdml3mtLO5k/Nut1N7AiJhJs5n1x3tLtBcb2Cgws8q
dKcb8ljdkRSwyKluEEbL+Tz7+v89qgUU+9vjdXL3kyQ8EfdZYENhFCIBFw2NWOgX
jwK541ke66c7vTTnHSKxQVwtkkERcwEpfO1Ac4S8+840rIpwwPf9CgBGT8s5BWiu
2eLoPFb34zhgDMI0XfvCJuYPgsToXQdFqMhJ1Ddjqx6JFhiuT0a537oUYvD0nra4
nI2is7VgeWU29Z6D7qszTl1Mtojm21mViYOYMu01JvQm1htSuCZ95W1wP5vCMdwL
H1n2EDdF9o5vWFvKjgeYgaaM8PGMd2gtbfoEEDkY8yT5pI+TPkPAZ0yRi37VSPQ1
0S2uCc3KAO+gGvQQUbKAfge8s8gcAAsWCsikFsp1rnnkr8rX6yXxC7wWK0P+z5vV
HoF3PS9jR/6E2Vvivl9kH9eo8Y78xUwrljEkZv0O8vD+Madk2zPUDfAne/MyISPx
nCU+oeSzWPXEsOJlgQmrK4Xj5exCJim3y/Vwy6r9gddv8CRaX4mxHW/DDl04/dok
CXUmr9i8M95rSvoupGgHg2yQ44YTlegA2ZNcuNKItIhF17aCCtfP+tBDFudMk1Tt
rPtCR+Br95yLRMJ19ea43lYgtLBwF5q5ph0mwHWIjHM7yp/PaqNW5wCIYRvH9bgi
ce8cXD92IO/+p0Sdm+RlMl00nSwhokgtYK7VAXbQY0/A8wJgTOhpAU0b2+QFP37B
FNQDeUaQsc04LYpJ1T3FCWmZaZz3P1LcEL3urczFPJo0YGYa53IQiTfpG1nMLxha
4wsZHdkek/n5bpnHsNhMiwjL8FzjmcF9RnA3i4O8/7NSfUkKA76xoA8HpsJKfO5P
R/iewL/ge5NKZWp1qGCgKJpDaNT2hw5wme87o0i39GOKxjjA3hv6R2cHX9kzhkJ0
2x76bQ3WqI9Zq2uHrTqkiM0gXR2zWwlAwnY69WigiEHO1HV7OBKjro3zAytyGuIq
TdiVJ8zFiWPIKB9hqBFiJ2NegtpJp5ZaxVt2UhXTck2RWiRzl3h+v/fcPXNhElB8
om7EMnj4bxcqqj2kfNOobMjL0qpgzmPTHkV4k1QLeEZGocoYIyWaG2V+1bXIWwq2
p62D+uzmc4owcvGEX/efX6kGjXbYq0tiskSBg0g3wWC8k8B7CppQHWRwOWy1ZUiu
p2mXTBhGVmpegfN7gpk7Fl2MVXrYSxBvi/Q8u/GiQXpJkuod1bFnZC2Jz+AhFPEe
RCSwHGVqP0qWnUHhIquLdPUf7/NHU+agfh4xDTk2avHDSRgCC1ab50G9HXwRZRt0
UOTXfGOu7l3QshYBRWxea4E/MC0mIR9f+vAT5gdjhqc23SjIATPEh1g1QYN+wL3v
xjO+KzfuX/VMHIUu5O+zaGKD8AVS2chys8O51nHFKPXA6jIVfWhJFGvIvDwlS9yn
PN62PRtS+sE95J1Q0OocX+hjZEAoQuGgHCKhoNPAjyTXENMj5oMTD3S6dnHY7if4
lVWkGOunig6ksi/SNDVOEDurXyv4XHtfszEs0wCFUFsWpHNrW2K5HqJNX9EA1fzH
L7rvld/+oTbOO9WGKhstj9INPXMZwBaJlcppdOHcfVo2ttpzkdmasPI+/a3NpWgD
QSH3zZABjSJ/HmnRz4J5AXTj1Xc2h0HrP2XpA90dqXJhl1PkroyqhLkwXFCytCCl
JElElVNis249ojGFdKlBvUGtQN2oUCWy6XCR97tacXbYGW9V0XP/Bjw7taBQowsE
+xfHNBevhRIgJEyvEAxWlEXa/EISslKdANhhbxbEqPoTD8E2cI+5lZqiEcAEyg2V
3u8FfdWSj+qhCW3ySTcFqXqQHuP+MBRrmxKGLOx8e3FTkRXgiFJcJUo5dsNpiIjC
KMwm/IHpPjmRmgC+Elpn5aerw23Z5mDay+YJhHTYmtsCrHDXbXykbxJhsbyZW6Ib
XylM8JTvcrEkPEtDX/5TmvQoTvez/T3Q3BnXCDk4ZUVx4EF2OgxAW6fa4XmF/HZC
tMYmDp/SmOw5k7shZN663a9MEaE32M/vum9qmti122v90hNnDUYcPn/9UjZ//UEk
XA/U4POPsrUjBRYpCNFd+1MwJQjDGTBaZjFAVg7VumlPtk7HVFIO0J1dCj8n1MVL
qtaVIVwogDVEdl/c2FmOsaaUNBzV8UraezmI1klRljpJdGZNmXqw2sR8WE4MchwP
igAaHW0nNT82e9rW/pOY7VKAvdOaIhy9fIjKG5WcrpU4O+4UdN0d/SHKVvE7XIVM
4KvehDnMc9zvBjNZGaX/C2HS8thAAb2GpNIEuv6xZZciFF1tjVDz7VO+m296SmGM
RC8W6NED9u3pjQkioH4Kv0/bMuhaXnbwiBQxBPjdbKHKDs2Oe1hYm28kKJnZUfd8
Y+WPmOf7OgaD0jhHM2bgdfZUc77OrF4o2QGrPkmgO+3wGeb0wNoI5BMOUULnouKL
5f038Qz08CBzakWlbzH5n5oY4mQApPJ8iMjuv/Fa4UV0s5Vf8Kjcrsro607Wcj+T
Y5eLdW/PCf807bMTkTEA7nDJzbk7M8Yrumsx8mqoy6u5mdebRyt7/MiH9F6O+cLS
JtJBglyx+wXFER+6kHgT6BWD4yvKCh0UG7P4LUZKjxfqAyfWptPQxf+vD7O4+UX/
0Ck5PqhhZD/s+B129u1du1w8X8kqh83ujgmnPInOLF4KpQlN9FaBREEMUS8aBg3r
j17H0g3KkalaKJH0cN5X2C0H2RcD4xWKg6dk/CgzR4KALUSULiZg/PY8/ucdh/mw
YrBGd6ZJ+1jdDPK/qIv+ViEamPzT820TNj6I402xMdTLKiCm2+Jzq0dketz5prr4
QhH1j0kIc70VKRCV5ZonSS3LROkn0nP2a8gW3MNVQPVl4v2/ptqmJRgTzPFcOvKT
pJPPHiCnp2fIVvXhssGds62C95TBgjEkCEp4tWumVSPHKpFynSMYw0QyLVXhxezC
9EVDnz1l9mpzAxcFdh/OyLrX60UZYu7l+AxOQydwcyjMDy/o5VMibfuUnQ/Oi0or
8d76kLIbzafTx7afw9kFpH9gD/8skuxi/sty35fXrGMwo2Ux3d3nuPuzp6i2PLX8
1y9aAoBmZ/49i5hUhiitAeWCoGgwApi3h2X6rnvL3qrJoiWtjWNNNQYFW2kVJfI+
I8o5ERMEKWEpzLBskawC4JyxBU8LF4FtI6YzNk6Gn80AMP38pRSxmiOrgLUhDF0b
42N5xOvwc0XbCMk+VVqvI/lCp0B0e66TII08MTp/CPqyisghlLcXft0Ga89yBng7
VmOEaCXZAe11GaREDCMoXaZeIwzp7pPGthO/zSK4sPrNcTJNYvbmJ17oXbUcpyt9
1uZZtHGXXKty0d1PlV6TSLikx4ffbzdp5b8ojewhId+HPrPkpbvKbWRJsbf0J1zD
CvnNAIzHcWkOhP28K0TxCKIVlYltNXUZY0UC+ifwc+ITcuaC9MmjhS2/bm4kFqI0
EkSbXOdcu3rfyrd7s7zthcpyfdmATJM+XE4hfs0rsTFQERAeYh5+aTYVuO1BXnLu
hVe2251Hot8/zO5pksPEklVJECWoMv5DShB9iqVocV2SI5OnyJIJHShk8+JZ2U+Z
PkjSGhnXNo9ElnmsAF9p9Dc2fWxIgsingY5G+ifXGqRmD9xY/wt2qBDtbFPusg4P
x5/mNe35WfOyiwEwd3NP36FBcpoSIMje8CsaMaaUuuOEACsD7mmWEQob+H1fHJwk
89LxDDCdTCR01ludWdod+IEfaNLm7D+XRDtYjDeq/R392ZVqDzUS0OGhjInMvjGa
RbMSWH9kmWcYZ/W+X6v3hQ3QzfchHgYgLw1qHgIUdiclExapgESArwsWyNZD+QqK
iPNJqStABurC3GSFe3XJ3UwQAfeN8CiAEHBctAmhNfXaD0TpwYXvGrUtqYonvCs9
uLSiezxaFOPI9rMf14/M43nXLAy3j9O3COxw7yca1/nWjvEhOaLlhoOj/P/QNbNx
j4ioWyomm3amQSJ2FZsh7NS9mQnNB6QPzXt240Dpg2N4FV38mj19hyOET/hScIG4
AC1ZY+fxUB23W0+V6KQWzHiNTApyOqhuoJBH2sy8sk76vsYMNzN17RhZbZP494b6
vW1FMrPwV3yrLnK68vk0m21CqSWfOkYjHAy5l/ceU5m1oae5TwmmKgnxTX5bFG6D
eTNXxq8poOyswyd3RjYzhJIImCxzTLKC6sbMebXmHA6IhhdOYNUxA11/ucLxc6E3
gX0/fTbsiTvWWo4JGlD/1esqvapoi3b/ffooFljJHbvo71m50lpzHP74LZMXyHz6
/Pjj0O9vUDC6fG3OcQg7GsoOm8j9sUG94O8LuTPJxohtUpqY6bvQWFS4QkYFWgho
GF7EkebtQAYZynVjpza25wcl0a1CcVdSfiXZZ6pgzl/+tfGUPvK8ZZ6c/mrButDs
BqGFWlQcNQ0/EhJo8x8Vk5tdmPXr6YEcDmOswP7ahBttRX+D9J+K283a8XUY+y/w
hUhA1oO9UGlEL/89iA/YL7JjapsAdZWh7HdVLw8+ArMVTPweWkQMKko8Z18VCUuI
D3XomxzsP/xvngWhU6II+06fxwNUhk71WECLAz0FM0g6I6jLJTR1n0ZjHdBHWs5d
+8IjXQLQndG/c55/fH70/Ux1DsSsiwcEpLc6WNJz4PoyCSbfdXQez1DJz0OZ/qAm
IZvQ3jxY2YOxdFv4N+BG9PU657dVFRG4G+ouObdYbuCTXKjIDYJevsE9eHt9FnDg
ExQDeKfLeXilVmKuTnmw+M4v4e4fJ5+YkU59m8lOaJF9yrb2ePYPQrTJX9lTAIwD
Jk6USOupoaqXqDRkPlSWT/cVSgFrqLFtQ6dkphRrQwZHSd+Ls7jE0LfUSa+qN+du
rQVr4WncyU3noKOXDSJb3vFuJ/xehWtOdkrKz//xPN6SXy8dIjaWhp/mXMCAkr4u
RhsL5ki6w1sYpdVyESva9DPKlYWMZ486Zzy0geZbz49lUcvCpiEnLyTRYxnpxymz
8t+LAWr5S7FZInwPHca9+FRKOvyeD84jIYAIDPjK6764nohNFJnABy6v9mm/NelL
Dfsrt72r/eCIIEboL53oyKlQN1y3X8+lxRGGb++KxUpr8lBE8VCHX5Azoxt4L0Ft
7AUbSmrIxKyxMxCi43TBid9sjsiaZdt81CKVOhZgy6g5Mn/C1yFrdGnEXInT3TY4
En4K3/grVVRLYOsq3NR9v7XgWsMj9l99+k1IN+R099DzEl7zEbeD9FzVnz8CWno0
scfYEfjEDVUszrMoWHKv4uBwR4aEGFglFZZ3zVMpdEcqazD7uq5uiPQuRGDhtjG3
IbHDzt9PZhX2Fzlc2kyU3hl/rm4951H+YM+tTlYmAutWF2I6D4WM8W6I1Lt18XLZ
+dVeBh+hwV8MwSmVLKkEKVbUnKlzDhDe3OyKsvdqkgQQ7m9NMP6mFNeL7ynnvEBo
SbT2ddWj5QqOOWsJu1M0ny0JIxd4ppRl2yA9TzXf4x8bRqdhXabueYAv9/N5wxZN
PC+RirHHwxxg82M4347yZPjE0iXtLLoYILeXw75DJDS1TMaHe1KZjX+fefc1ifMC
p71EH00f5pSRqaEwNhsHkR0yR8fmdTZkYFV8GAlH819AftbO/wpJag/daYQFe12B
xmnz3ALy8q4BDzd9XW4vhkIpu5I2HOmXZKpaKpUjxpmcxXdCdXx/sDWqi6p0R/s3
GbU7DWrr1sOzyvGmfdBUwaVUk/VAsjfCGpsrUG2x5DAk5SSEj7qemzLSRrrkgC51
sX9t6wWTPN0foduueMQQGobTYDuRXfu9PhZaNybWxgAi+s5JYXrRGHZCkOAr4nr/
7U2wyatzkVpUPhWXUXzeH5Z0G59a//w1QvXgB2tQHQtfuXgepGz35hqfVEQwwEkU
djaf7XrdVM6G1FTJU8GDrTna/qssfbUAY9kjTSnfqIaKPQLZKwlcjZuldstCYT2H
E6W34ahk7iWr8K6OyhT0PUEj5DTjzUugGk3Ny+vQhHoWluoBN8JlDZZmS0vlDy0V
K0OOaTqKzxNTOQKXSFykK1V5xgFL5qH+CUt2pHluG+kn9BLEJJiqKd696vhXteOd
792/GUIQhnWKUcCRcEEQeJruPAalMUltCAKNG+P1vgvmnliX+D/9zrULTeCpuo1S
XmCmYB3Qft2kreCLpRj+BzHAy5t54WCI+qWMJbz5osnTodDLg6oUCFXYjqsIMwzD
mtbSVqEkquUt6CU15QV3QO1HCAL5/8Ve8HCa6zd4Wo/d46M1Idm5qbAHqex4U+SC
e0ZFWKBnT7JlBuk0110uPPd49D+RaTDUb4PPtTBhTHkf/nT/WJiTDh2NNNzPn7hE
keKwwMvO+OvOUVVMANST4sZIYT/Ho9TyqE+e+blMFX267BSpR3nMr6mvUV0Swd7h
JTjdFfrcenpZ4lmmqcz6HjLcPriiVwJXSYemIopEZ0KFPt+BpWk+tkfxX4KC78PI
lIpw+xnBOUTxaZfoGaNoxtNdLNMuRwBLGyxj4EFhr0pRG4tPN8aHcfmCmOpyXVpa
zejqAisCs9RoFv9pY0KYt3pSi5jVCDU7WEiCGNRAeULCyEmYixCqlDuTlrW2tggW
DUEM6Wsqc9LtzhaEjj83jYHcins+211QReyGqy1BVy44AjQqq/Vjqw/W78+3vwiq
OdDqyU2HTB5D75/KPWkcFZFyowyzhXSpVVYYN4JUr0xV8w+UK4MYISHVd7D9KjL+
1heyynHx24DTdXm6U1euRy30TKIPxozBzWpw8npbrntxr0FU5gEdoySsdwEnjHKS
c6FMAjmOfQ55yoQitWch9/c1rR8Dx84LgHfKucAp/TL49pSVsiTK8Vnpr6t20WHh
V/N5otHN0FhNEEwHFPs6IhhP40aWcx4WBi/M4aM/C3DflhDgTqTVvBcEi+XSVocM
5mcOiiz+tn+/yj8Zs/GNpTZqC9ezJdxFVcvwOZy9Bwjwcg045ToWzEb3l23eDYUK
7aZM+Axj74PkuILhzWtZwFW5ewhe/QXN3+VVUEDZdit3aa/ei56QDgDHPxESYDKQ
uzvZwF7chGK1k957kgzseL9TN17+uLjjFDAZXxJTut5gJ8oBYY+dv69b3mYxljrC
znViTVDGMAmhcFvt4QqjSd1MPb//Q1uMZlkQgDMlyFKYyoC+lOp0NoMberP2b5lC
stpqa7Qg47o23kAXuVOwMjcFt6QOPdJ4PUlkkTDBGlmjjuzDdNmZ4aj4JxLa9PSQ
BID2F9uc3N6Qvf7tD3DacOpeCuD0webRIx1pJjaFfhBZ4QCDrDDFbkr36azeWl4k
6poLmj1Phlt4LyDGydaYvREr4nJDjTAxoQ597fapohSSmo5fVRtut+9quDsduG24
UVFDYB58h7c+G6qiQAxZDEOTD5xAhe/sFC0sCvKxTXPFEdy0LXkbzJxsax7GJ02a
SudAEL9HOFFIh8C8OCiysgDHKCzkDroU/vz/XWuDnoZOdf6MvPXvN0o4mNbWq0pq
Hz+uHo41lO6qGfnSlSuBZ8e5Ps2B78Hn4wBTHjyOqK6F5riUY0+e892kdBJeUHYJ
511XduSHj1VNFwjQSkOzxo6Wb2fSpJ8lSQ1VPYX//2ppjqbKor7IJ4n+tN+LejlT
wBhTSEsE/nsF1k/zDQ5i7doCc71WSGSNewQu8LC/MDpAvC7rhsLLcWiQqhBy0M9r
yfLq/ZeWg5nxbJ+r6UMTa0zajyW+99bFb2h/hZLk99msTFx+pNPRzOkEK5ELH70j
yxADl1KmFAQX9Ucsejp4GEKZASrSbLTJZfk1/C6KDPfLG4MWa65hdXRCCbN6bmDN
q2N0F4BwZj8C7SvTwlZO0663KsHt+5gKQJCJkIw9NCK8mDm6Ot4KRkgjUReRgYHs
RfQEjAlDdj2W6HEKx6xNoFjN6/lAJEUTCq2YTj1xSmjXib70B7yUYW1mfbF0r7L3
T/zI0TPbDha48NtbfyTuxLwaqJcCu5/5Ah/rdYTSUQ+TS9jcgEfzitPz5Cm115fH
vicd+2NHiWcRdPEgnp14WqLIRiC7uUz+WmRemYKvXaJ+wC+jPFTxqSkHe5cYdED5
og3wk9Bj1I0QiSWyuC2KqoSgzzAVRUoHmlctmKtkRgTryb+pT/8UEcMONE9G2oMi
7FT9RFc2hgi16KbeuiTEVEs9qAAPqZ44UnGl5YLvYkQBpkqxxQkgzHjngH+ZGVFq
fzCJlWpHcUmD7gY5gsD4kuKdZaEoYMrZHrW3r2k++khGBuuB2LC0vfMCsIWtBGmz
bC0ht9ZuU5sfHnetYL9VMnTTmgKenAXZggnDuDniyUvYKCj4kX4kOP8dMhKWKhZt
lIleVgX5EoptBkJPxHosDsVdll4VPdTIruX1HkVySM4ayTXyzk3ohGiP5PbuGToo
uN9gKUO5Vf2GvwJV+DGoabgnIA2SHFj9E4X8PsPskGgOh8mKu/w+gvcZHPXTw0dI
fc7i9AZFYOb2re73Y/3Us0CRODRmisbF95rQlKWYZW/djunVHvlCoONEegB6TniR
ccOrcCNpfIgl3KZyle/6gd7Ng7LvR1xlgWPK6DOIxDwTT3zvNp4peElCGHsxiNVg
3lRlMDoQNFDQW+bhPy7IcFrsqv6swzqcb0PN90kM6pDzxfPAuRnfl4ZddBwp7I7k
a1nZWkJv8cb8ukxzwUn/hucGS8WbOuQJD4hEbvdlSP59qnBvWhy42Kpmf6B4bYWP
lMDsIe4zcuM/qQe+LLO1trVY0RWrV5PTYVSKHWH5GBGqUfiIepwSV91m2PlWhV+8
4f/lUyPDa6q9xw4gUlpGn3hMjTGdmzk+lZ93LAwxCrz36BRV3q2uHIDmjZPQzC/E
XEO7LE3sZ2aOMzRZpZidE0+81h2cVliCQhc1KrQV4UcdpgXdnKofvEWAKSHIWPoh
gnyCvyqw5WYtFI8M+MASQDYJ1SwpWMCIEckZ8eRjcd7TAqvQnaH2Wj5YjQW1Wlhz
LylRhTSMIiPEvaG8kSerCVVWqOksNlUEHquaBEN+hoM1QjkJH2RDfBhIJv+IkccF
o7WyjbAH/fYToui2Yy4wVhvhQ4T1FZ4bOhelEli/di7TvA6G8vKCf3Z7H5X/Fana
59NWBLeOB7KLBcQBBg+aFHqHuZ1dFJwOUKTRMn462YlqvnZZRlzgPQSOs7c3eK+q
p1yYbAWso+51uNfIuKcJRJXPwAnBLIgJLqaicgyoZfYReuJDYKWUa+sXcFD2RaPP
qgZQqAmEzluimhOp4utpq+mbhJET7ztugVaH0mGEr0umox2GBjHo+NYc1ILZcVT0
b4iZS35FbCoWzKfLCfqUSaKE09mthn/+HWu45519XyK5OhTPavQBOjVNF17BZO/9
9EI7jcThAiBk6+LuJGkoAL8wp2SmeLhl/UJdojRAHF4VobnK3XTIxcvU54ABiTXL
DLlfEV6VsclmGmLTPZAotP0ZbhZDa64HG0XM1+DEh84pVXq/zrgVfmvBl+NZsYlw
9uuouyQ+7WEsAUxMxlv0LdfBwo3rr1FPSuAsB4XyW9zTBtZaJtSWgpBleMEGfJYm
p7A4DH9/3X13CJR1HeumCMtfJgCY/583tVG2ayATFwA793v7DSno23jqWLO46c6E
nFHO/z/D5HFpKJ+F7CWz8Q0ePDBYje20jcTUtuIkoTRfq/CpM1kkFMAent5UcueZ
iPVQAwtcm2ECN/M2AEuhcpg2h4i7XQ8PLwOoZ7Tb2eGuBuJcdlTrvpTNGunkSQ4T
1dz2EmSdV2wSCNzqINIUu8pI5y8eUmDJ9u1AE90CgXpvx8zcRTQN/MRNKLn7aSTj
5FPZTCDJodwrdVZ1P50ROcgqb5Q1ussLr32pxUKQQE96nKEZD1CdFLIQMxOD7xB5
3N1MXWl0h18fLn68D2EtUVnCt1KyOcYWFQLp0M1e2Zf842vyZ3jsLqHWMWQ9DGVy
LzFCY2wheIxG2gYGVcUkq4D0APJMheLfoUVVeYfTmgxMxV7SA1vzQZGnWBgoSQEd
eINS3DXzjYa+ZmAYIb7rULvm7fnWo5TRZf/qtJp6mXC8PvvH70Rbb6cq56D7thH+
IxkhJ/EdJeBKdOzZi3D9qbfHdCTcUqy84fVsgkud8UfYxQBL5A3VqRUfEiKjwOkl
78dUe3ePM7bRJMqB6QOzAfDvjURfiu/XgjIXtVjp4yv0w7TrsDKJHywPJcJD3prM
wanIAvElwi8CjvNoJWIlPMakvmjDxAABh8KpEvcXv7zMZgQQf1aSEPx6GFE/WOmI
yTKcIlwK/QwtLGcSATtnbvrAcAzPXDBSNOyyZnYKBx4yO0ykybztc9f87UiGIMhn
Tj3mEl7VT6VcDPeLqav7Y9mvdcUdw7Uj7kxq15YjIw6tT0UMCffa4O/4jI5EOhLI
cFSLFqrRz1P3+w0+M6J3wCnMugP4Euf5y+Fc7wiR57HQVr139Dj7BuDCa0sA6vck
xOhctW7ubgsfkhFW+YH3JDqmQbTEblTE7aG2FO5HAl1h4hP+QChMOghXeW0iHU9+
9/Bbjx8XtDsfzHvm2EfrmwEvkJDs2dpGDp8bdzIomD223yvkqjYKrUxKyoNHb4CA
3yF7vXT/OouJG6tqrSXcgtysfxeXyL1IRIl7Ue8zZUj69enSL0mmIh4yYGwBPIdB
NlyAAbX8p24g2YHf2gocUqKvL07JFgZ0XRTeRT1+4gqU3A6RJsnUYDM6U3UsemyY
4jFbd8QCWtobR4PwZ3PBUcCQgWDLvzteH2DIiDAZeTFimQy3CRdUO4Ty/4SUOGfr
VR5kOPsK49ToiVkpsSlsxrv2txwuZleNgvyXmrW/qyzhMVEwOEKCJIyf1u7CN6bj
VaW8wyzxp1MNcrNkzZksjQnA9T9tkfZ7l9AOsIbNWUomNLc/ZSj+dlEody3BbXt7
w3i7jyzTnPHLE7WFuJlrtK5ZaY/6P9++POoxKca8V7wi7LNbyrFY+pRTrHNTJiSf
tIZRwsWvZfVXhABqii3u0xNybMXd+Iex+skcrLa9koYWh/Gdzj3t8lIMyHkdYKFy
5WLa5TOEWNBP0p4MZBiF3LVH49DY/3DYQesifQpTWxVO2TRTW9ZUg3V7i2iLEUOy
l7bQAgFh5R6Cog6fhLuNl+ddEEPB191PQIRuFKEwXtfe84C1Yi8TBv1At+SrJ/Qd
MIM8+70Pq5RdfRVL1Vsmf6H04UAZlNaLnxSAwtKnbZPECWg/DAIEApMQl8C/g4WM
mcPejx6+QFQOTjCIbNYLDFq2OW0ikT+eMdgWAH6RKYEGfp6Sxjht3gjXYhpUtLQY
MmGd4okh9c+NYG+b0mCG6MJ4eTu3ihq6CzTpV1Q9W/x4zwp5hkKv80vjhZi816QH
YaP9ABFx1XTYB+n8g9fVhi7hpV1yoSQyZMRLNwzbpbfK25X1jIampd8ttWc5UXBR
+kpvMjTqo71U8QXkID/SvL3hKVxl+WTmqKeceq678qcHhkHFJCaZhMINQnywZKSn
SC4xeJUUcuhIEKjvHB3il/nIGeIbyc0c6GRbs2azpDQ15/IxLNu7UkmOXEa0se9L
pAaBb7IqGjbG1p6IriK80cEX7wFjEYfc6fYS3Xgf6UjHy+MvX6YlXoHzVxWj1QbF
Bq7SdK83l7N0NuqRJv1Ue0wx/6rNZfGkvP1ykn87vt3FqTnTVk/UseG9KwqNF2Fm
kDutyCn/MujNLYkK1bvLPX3wfyiVLurmBg0K2l+kBlPGpyKOSrhv8riwJmkH5sL7
a0BJDO+0ohm+Q60wRXHZj6hEh7eF1K+1ES3TagYy9rGLZNtdcEZ8w5TgWOIuAsnT
e3JFq6mONFa5/PZha3YQMlgJddYOoxTo2x7Nh5UBbBFu8FGlOy3gY8Iy5LHmNMjv
Z/yHTOxB4F/WcAIdX+/2foLK0Ae93S2bnG9M+gESFgQ2XTIeko+gfT4Xe7WPD2Uc
3WJJKJZWSZfTntuZ+kgMtVbUwDdk7tae8KlBQAHGm05Zt1Zy/YVR7Gzl/Xv53W67
BSPgpKohgNOqCgsBEZDFa4VPRLZ6Goz9UkQHjM65xNTlaJ5jBS9yDEbJBauvEQ7W
I6EGxu8uoDAumjjAgAw5Rlxy+BUuCx4tvDZV+xdLmnKNDTLonq9/PrZp0tn8TdbG
2T96IXxOwFFn4RZHEFLI7k+Ee+ZRbW1MpUuSPYHnOEsOPxDhIpizsHrsiajlhxjs
ejX93Qfj9L+9CaMjW30VG5elQYKIVS6kboxJXNxxPsqDMXF07Yw0ogi0K9rRSoGY
g+OJluH//+tsMiGzCO1cAh5EqB4W9m5KwGBtb5bEEr42UiTkwqPG5wJn+EMDTZfA
awzIqonwgR74+H/xSUl4IJ1ZvAYU4Te8t2gEMAigWUPpEyfAyeEDaNEJi4+IFZC3
tQO+z287NoNSavhZTlaRQHpkBw7Y4dFqA+ilNabG9aI8aAnVIq9hA6sUQBAsmOpy
P/wPUtwcKzrG+036bKHje9v9/CQTnJ8HHCKrQ1DSaG+1dxBfaikmAGZWWYqIs2Al
LpQevL58RrZx1yLdngKZsPGJWG2m8oYWwWRKXv6wIowCg4+xMC1Kj1D7Q69j434D
jlI9F1XAIkj7LDAJCeiZZx12xA2pU13wKWp+JPyvFlFwIsdT7FNOQkYeehDmsJXE
XCbFyMeuG1lgEKYW2uKzEJXZtm0GgaUZuyfDSGpXbv96o3FLSSP5z0s9QyRvZWkt
AHH+auuEaLWf41Fwrf/6tKys22LpuKw4vLgGRTbfm2gv29ax0FvjRKDWm5ZfA/k2
pQLTvAv034L/SvVZiZYeXuCvSicYEyh9hvNhXWbjgEHFqKOfvsyNYsXtkYqt0c+6
uZnfabHa/oiAnEjEpRjFa8HbiggyY92lYNVW4IN2lqHHxwexm6WVzT99QpNpi39A
+8JuEgfJBIaKM6fdokoHPaxL1O/c3rjxdgZ79at99HgbadbkiQ7Ggz63orPx/7t4
Ze5378wSHdLmHboiwabMaSUk47Jp2idMzyXdxRxXtw1ANlEZVPPRpXzk/zuOXN7I
gayJhnSI+jBcyrkTIn0W2E/OcVkvubrCAnOhNRBL9O4B1TaPW8UuZwqQuSnkhgvI
x09Wwa5GSojJgmstToZE9uinBZaJ2cZEBiqTAFTzVb62kVrUueTQGIEoL0AGiaKn
EXPodQUeSMByHe8PS9DbNRGyrPkBAqTwcjEIU0N0tskYJr97/8Ub6z1VVWtkQEGM
0v66t5g3jQZL1XiSzDPi9Gaa1seYnaI15BeSdRLLd8OllBi3eniYErnf1H0LXunz
aj0DzPjx/7tkhg1SflhAoUnqmSd+gwffZlkS7bg/xcPuOQji+WpVlxUouHmtRNeI
VPvwbI4JwtvPq6ymnWqe8eTXXcKXO/OXA/JnmFctox/b+0cM1VHXjo7HqNsqk1+j
EPGwJ65co7VYyyZ4GhmxBHwpmUIRMAnFYBNsgeXiU1ziUbgn7lfAX0BM6XZB6MkG
x+FQWHFhEfwYnuunrFkp5MSwEA7xa/o0Lszg6q2SYcnk6yF3PsHdgkjXjk3tWauk
od0/3FFO3GVXC30M/FEKryGz71evKCPC6z/EbfaAPCujJ335ZMOipgXppv2po9RG
xzkYmyZ3pmT/8sPgYF3jOSe+mb8VGARbJg7OvUZeZrqfZryHo4UIBQ0Mb26UaIBg
Kala3TT6QrwGgsgTuHpNgPYI9xfq7RXV31smoryHGfQaMY1sMg8CC15iontdsJgJ
p+TIMDuB7OQtheIpYcdzDsYAN4jRYvKfVJiLzYQ6a4GqvcTaX/S23sYvO8JYPjBm
aONPAdbecUeN1aYCqC3Dkup+vmv/cRXWZ++7RoKGfVsba1JCibRUsY55fBxIB1tY
H0puoW268QubOzLmbr00gFt+O0WXwY5GrmHD2prtNbpOtaSu4h6D4T32ipOHq11l
BLc9BfFmVlMKq0iYp6ECr3Cy3C0+bHVu4u6xV7V57QnkkdWeG+XK/b8QbUkIWF1J
vnclUQiT+r0zA30KHoepTI5/+lITfpqRVD0T6YtvWnivyWCKTvSL1wO47OKxJHN7
znsKzu3QpqI4io50H654ik2N383dnfrPISXMXp+cSykzpUR2wJH9dSu0MLsWOqPd
X72QxDB0QL7+0L2oVjjkIzeVArJrAhnyrWnLlz68jVsmv9Xd/Ldb+kOpEsz6OCXP
1ppoQQQQW0JWK+vuQHTTzOmZah4v9vhEKgP9+JUe+L9w40ZEtO7038gefi5qGBNg
uZc/JP7V1F3b7B2DKKIcX18hN28spVnCu1WtWcVxV86qrVxD/QQ9Td2tyG7Ef+Oz
LVeEyX/KuccpSNXMwxzoyqzUVM/Gaep6Ta3QliPdav6PPFZWeE8Xz70xsk6LKKYQ
Hjbo/mTy+/gOXMlAFUJP2HJXOsLMD7Ai7zsPQN8DEYXkOY9FCJFfWNhJf9fAH5ml
ZZTFzm8Dz6J6c9Dklr7E5DjtFk7mism6mZi/q24o7p3KobfNSU/vfr7naRCm087E
aprvUxFB6HndVlFL5GYek+p2M+N3Vfa5JG/u81gwogduOwQo5xCyhfzMtCQb9ifb
qZsDC0uX+ihYg1YCvx0EomO9G1fO0+wpqZ9yDFhNzy49iB/ELZKZPLEtbhpYhsLP
j7Hi3js+MnT39jfUHwajnvNGRj3t1Nj28zK77iQrCmiymQ91t933K4MFVIuDU+4o
sXKbMB8aVMvV7VAXUKIyy9gymcDhFIYNymn4A2x1Ct0kg2YZ8phCiNArwppXVr+B
AZl9kJ9GdhS5hxvrNrcW/gNrnemITD/h/3LFymKZ/27Egr/chQzHbhXN1vBWVdxa
HKYShppuAYt008oKD3Z/rvENYPSRZ9LimJlI2qXnURwkO/Ra2Epo15kSfxHUedF7
BMsWxWn62ShZ/+5lMWiZh3CZHaR8+3R5qcjvWJ92rucq2FALpKTfes8JHE0Z3nRA
2a5uKxauSSrMwdyBiQ/QYUON1n5612K7FM0FSBAIW1ldLn21LzaHv3UF1iOuHhZ4
hC2/DQqTZ3FibTHRRmpdpuapwn08dsOeaf/8O2UFJ9YIkitFgnjfbvimSfSj17Ht
4zpbNtHLM8+LIQ39Ls/cUTyvQHyNdSRwHgImc1I1O+ZweVacWgcNy2i7L8RD9jct
19tvZwFtDdAV7lZnBtUmV2GgIONOP+KjiCJPd1dv2/POBTOTJ8Xh8LF94xg7Ngnl
UVJPrl76IbAgnH8UgQZmYZFhapD1PKC6K2lE80B6OtqhVeGo670HzFboQjRJRncH
4Zo040w0a/mQdnnZjcBDE8z7nl+B5Okdc0KEhSgmmQT8oM7LfZtmi72UFZzRtCgl
ELMMubjmw9YWGjNmuQNCRFD8qmh4orIG+AoerGt1NG0qyWQ1EPQlx7gMZYP0m5fb
A57EQFXxUb2WeAmHy38wVDT2mwW1gtrvJ+ukZ89gBfkpk5Lza8DM5cJS9om38AKt
V/Vto2zrUILLGfYN9kCl0bO40ZGhDhf01ivSiVWhaorZoimdI3cbVso5Wc6SFv6v
M8ka4R/wvMsPYyklTWkNdUU6FOJKK3L5EkZxn90p3rCF8VgCxpc6iZmRNjgpgM3n
suv5+nqq7mbBNiE0XFD6tE71syWeztN1khXjn5q+ucsfmul+zVfrWRwI7KqLw8rD
hZQn5NOPx+bxmusyWRcLqvIqcBtEZGLAKlSkohoI2lMpUVRhCKuxLnapFFp4eStL
M/pq3ziiLEotaVaPZL4cbDldpiWc2jRrH6333IRMHteTKKNLYYWwXTM9sIZ1uKF2
/PJdZVWgqcbkllXnyuoZeU2R3jJJuxf4VE2l3jUg+RkU9OJUwC5ZIuU6meSr4Vif
O450KXVSGs0c0ckihgTPVdJ8jpkTsRiVx91lBG6xRrNH59+hNcfO55PWMD7lM9jc
obaa3NVEYDPX1INw0liG0UL3YOkyrACyyoC2v2yPtZd2CkJVuAiuMj3/kH3KKhOw
qhvhy63/qaKsDKxVcMiWZVPUlWEXmRvDIgQEzYkFnnIKT3M4SYKtFr9/8tY65Nox
GxDTUDRuGI3tRtEejxVU54kOHqanYaORSQQedvEKJGlzSpO69APoebaa7E02pOYF
pwrVgIhp9GVJaTZI3HrJ3gsMIYWPxgx1oZQ6WiNQeoUPyV95Y/fwiX3w7zPWcgnf
cwvQQD5nrptLLp1F9Yk/1JO6Ylf+lzOPcVZzHw5YkCtqL9/ot2BeABaCL0sctqeL
m4alhtBrcDOXL8wPzO0V2RmLSbaNO67I3u1Jo8PBCgMHzgxUOd03MCOQACednkHm
6HspTQsQ5d+QaP/g5VSHDRR2CIV4H/2eNTEkFez/Sqbpq6TKgGN+DvdiK73SIEMb
sIYx5hyASfzHHKv5hrus36x0ndwhHqnzOo23WkIaV0rQzV6C8hLq0OdgmIxQvs24
WOohRhBRLZy8DINbJ37hwPcRixcuENytOCX4HzIZiPo9QexCwCI5TZ/RMBLDUDVi
lwJurSFoEY/tPuSn5b9gB2UR71J+HubSNhXsYKr1T3AC4wqtQywcSlkb1A+i9QJR
ngLzGefFL1C1pYeAuE0k3ZVFO69/QXPLeetH+EvjXq+MT5YE0GjvTeKvrajK+Jp5
gNB5wxBRoevpVNFMilRiJAs3F1UItmfbrvSozVsqRo8k0KKl4D8SLeMs01vyMR09
JsjZediMhZpq2oNVRxlqr/PINK33wWpuj3NwFfwSgkq52aiL5ybleF95+byGLMgI
DijbWWv/gtok10xsaQvIp5SJe8RQC2RgAeWxWBCelUw7ZuGXS7CzLJM5kVO9YXIH
mt6eNnwFwuN4lzFR1yqYR9uy0MysCIu5+IqTiw3oVmyOdiihky5YO2cvqzM/u4zr
3HC1WmAQLA3sF5/gyoL9TA6SC/8EWYxtDxDWvsZhVbIyRBozouqJxTqn92BtJG1L
gmZUhoWKSVLlFhigXfcdDO5YRrQyoggBazHY8nBassp9DT6/oZVAy6IiodZ+HQ4I
eH+WAmNoVKFVfoYL3hnHriQXHtSSOxYOzw9Kl4axN04lgeS/H7gCj2kH5J/looai
oB41YiLxYzCKyy/wiohpGHKHY+yCsjR56eMOZMQLjojGGyjSbYlIv8ltRL3cnTW4
VZUh7WJr9KoiUtkxVqd4nZ/9DGWkH4b76k75PSs2YgyyyqyYdf/aoi9wZFS4pmMh
E1grkMqQ+r/6f9uZcZ20NJ6tjOu0yYsxSof+bdNSMXo4NMZnnETC9VCV2OweGDsA
5RQLAZHDia16qJSyLeUC5aN28nNg60D5KM9StxxnNVUsBuXrrSWfbN911rxT38nX
9QzhX2X0kJKABxF3xIpIj9zOn1IdQuhlA2FcioiZ+QLpV3fAwSVOsZaOecr274Q7
JUuIy+IszTAYGuM3lzIh4EGUD3yUqE0R5IPJ+LMzyE96iivOWEn0jScb9tCWJR4F
gt7rNGKRYeAVRR/9/hlTKBj6xGP9Do94VMCnBPo5Q/g0nLgGTg4kXDwHk5/nDlD2
Qo1YmEjoFlIhF8AMz8iGTvrQASpReoJ5Z7kI4iTlGrAjPU7EOLh+5+zzyovZlg4d
tuZc/KS16ViGgBeLRZvlb3Yl7v+Nca72CL+Nz2RHkoJsSX7owg93snbzZvwsfBqB
XFE91W6cBM+yhjd1m11S/O9btnRf9NedRp4utVUo4ABZUlrnxXdEpwnM6j96FINM
nvFhNnVLCKkaDuL1uOZKhw4UucKBKTrrXoK2fVy7Iqz7lfKiCmQiQl58E2ov1myq
0BYxd4OVrAA/ZpRL1+P8XvdJxw41R6O5KrFU/d/m+k56f0yvaBYIBdQSAnu4ADvL
B43RQ8L6lv7QvMMK6kkjnpYUZGclRk+j6UJRt7KFdmaKMh895Qg4ACLHAiHrLvbW
TqpXbcwKCoj2MGMPJRmkBq1PIG1lHBPA91AtUy9U3TwoK6l2xvpB7JzG3gxXcms+
dU5VF8Xhgnbrjs2lnY+N8r3UEYCqqWshKFDnPrK5SMQwW2ye5UWCkgEz7JnvSozS
x+KCmhp9Aldrsq6I1aR3arzPC9BYthI8DOGUzzS3OGM5bqIEreBm9+Bks7ibarh7
8PR7eI4HWWiCE3FttFbtp+twesfp8+EBYpJo9V0bwf2sbRFMqMN5juwPWEeuyHD1
J6QJMblqeYtYYEb9vU7VjTh7fbo7A+L8OTJQgeWX7TI0cjSWUUGh5Xv6eyR/1PoQ
vBbNS1LsvehAxC1yBEfYtEyFpwWZ5TGU8jhfSyizYa31ruOxpBhMUjydy+M5P2nL
w6s4ggaKg4JM00nZ7lgTw/zHtk9OOvTv6ZCTge9oltHhytML/QrvMiroTMVBgU5W
lCXbOX1lxvA+qqvcb9rZGLwX5RZczZ30YYDok8s7TwvoJio0rNxn162hFyeH/ApK
KAC6+fRv/PzYkTS5Z9gj4dpiIFI05JdXDlGUwOAl7xVtcROTdZitBSl6obl2R3lH
mXrBOa21AgER8ywlJqb+Qg0iW1bSHfRqj2K8CY1OZmRXl5X8hPd7zPPvgwtotU3J
N6PBCzwkezanZjjDjC7xjk8GKi6Yd9MOSu+EqD8Jdj7PeLP06VaU9VF20BbU9pl0
fDht5/4depoSpayLsJaC3tcWnmT8j/5xDmz/KlgmlGQF5+AcVIqZhFwoqd2WtNzJ
dCVIAv7L9M1SI3TTcj1wZFHN4BBtVgVqmbYygrZfvhQ6pRT/fk47Kknp/MUe6BSH
mXn9C04j102eSkew+8f+U0tyRS5TL3/q3BDg9M4sqMojUOgao9dLomOPJ2is4GA8
oS9TVS3DEI4eB/fh+0UCFkbFdxHKpx/+wntT8pG9axaF4YM63jUeHrQB8WMKj6Aq
74MAjwxKA128CeAuGyNZfYLSXOfaKmH6h09c6tXWMogY6RJ6H8lEgEdZ00qqi7g+
3POmRNI/PUOuIWPxwwI9XhW/LbsEmhu7K+eotibHzIBy3V9JCxMEVytsfZJduRDz
HGNhse2kB7+udILDYLL8yAzRKQ/uH34OQGJN/LL7jtWDr2kb1EY95moFoaTCnSz8
lzOsRNLWBY5USAynYXcQK2WwFgumrkdhrFoIAFfwQx+I1uzymm7OTUNHEnjfzv5P
jGB9aQdYM1j7qlrAn3xqcFOlqXKz9xCLtNGbny8h1rxzCLDskuOnGs1bmVwRSaey
W04pRa9XWJXjvaPuPnt7oK1RVRQNayGEv6byUMns0P4cB+FOJroJbGRAdQcpHOd3
7WazgmKFRgW8IE6d/dMlmDWCZCuT4+4L526liGIjHgEyvsIn8NOrZ0IA4n6+Nc4M
H5wWrF5T3QZk2UoanjB04w0/qD+EmPeBHfK4oLojvjXqU0RXBG+O7uVcvnmBV6vs
KBDqVV4zlr6U3L3JE2fJej5narIH6WYVAEj7Z2NZmI95x/m/leTsKo0DDBr3hcrL
xWaVwCOsxiDaaewC7nwHXwu4Gb7sTXrrmsAxR0wxskJaefR8ulT28DZ5Cr/4W2kY
Ww63vSiZ/R2yNOnQUfP+3oCCjSVAf20Q0n8d9qDFMOsvJ9ygKAF59WraQ6XuTePh
gTtBT7zSaEhW9yeceW8PUDNO1sT4W4WZOF2xTMzobZ84/i5WwW94hm4ScCPNk0YS
hviUXUDXgqxZgBfHN0zjky/d9DrF9nReaJURM7zEV+kt+Rk5sd+eaIK8bFnhLGvh
nBuq9VmaFJGyfmviTXYMvH09x3VgVsfTmbcXXBadPnFqpx01tsLU8CESTI0U2JPU
dpPKIthjccpsPm1omHrG5itgv0X60SqM8eCe9+rk6beTul6HpUSjzoXhVQVFLPlG
O0QNLPJ03wA4VVBr2P6OK0fTkt7kcGkg1juaYwbh4i4i/t+fBxSDWJjLaVaYX3sc
/3/E2k8KwbifbSsTgvs+P9RueTuhIdE6ujGXGwfmwiIsge6IxJJYj3MT8Loca1rN
x9mu6fg4L4+fhFwYflKuxiLqhHp9dvJDkMwebccmM+BV627Nwd4yXXRRFz35Wi0G
fv/IEg5R1A/xXKOCP/0HIPMclMDdTBGDrrv64NzWAXnbkK9/zIql24B7HJ2j3x6n
IGojE9a9KKkjpPCw1MawPKtHEtAL2Lx8yeiw6wDvHAWYnnW75jJvxOJ/7U+1j0OP
YyZiCtIbubHPkh+iEhlXnAGMskc7eNYM8oEwp5jNVEtYRvQrraz/DoBt2OBdNY4w
aLfQZETKecwK6/EQ8YecOtfoS1rrAEi6iKEhxyldxPLVHbFTgPhfo9Rq+3qTVRAz
tW0C6r/Mk+8+CqqeLFo7nlv+sK5JX/DrZ4SfzCG2YXS6oWhWtPVgE+Cx4SORE4bS
S8wVpwPmTQbV39AKAo9UaBh5jfpaosz/HVXT6LB/Slu2MxXbqrv3Rxg6ZuTkhbZJ
GhQX2eVTkpwwxzCVU8Bsran9E2wpYMHRbvcjXbG/rhROxMto0AOd7hnDJm40clpM
HTJKJ54vnbNuPZZfHr0WM6Nq+udjbZwMv+qVYuGWfdgmRMkGWDite+ZDA+EjBwSl
DBVVA/DM5b5qRavJEB4mbQ1Q2GqqMj+PpmNGeXEOxZx5cZdIMqpykEJOBU6lchok
nz5keASrgODzxA8prMjqU+5EQrD5ec/xPMf2mTHkR8gDDgSaQfMd3u3yRUuLw8YD
+FFAfm7GO2hvasDtD4lFS0SEMKaJAoZTXdxFJtcvMSBpo1IY2xtjg48s1MEd0nig
6yN+lx305+ntrKN4ejJ271+k3qtJJvjqCsU8VvZ2oakns6zoAJFT93RmhCYfjjAc
JKGVhUCTa+gjs5QZmFpKdKfpBeqvvVtqxprhhUPcwoUCrQJiWP0he44z2RBFOuFX
QSMBIY32G1m3qBh7H+dwdjyLfodxnRTbZXz4SJaZnr3hs7BnMnCn3x1uzLu80bPN
Nvg3aJDU5+C2a2Bl3/lc882wa5QoFKZ2m1KNgL9N7D3ODzTOLHiMJdnuGBUuEONO
rQ5iBTjxN4tL8NTXFwMqbKTihvONp/EULiaOt7Q9IxEZ17HdLGgF21X7W2VzGJqO
lFW8YlrKP7rBeIs4KcT52edYh6xJhHm2co9JWL/PjgEfm42F582FOrdupXLFvNEJ
CVyxwMKG+CGt90Uk18LK7DFIpGbyjjx/NmiJrLM9XOVgL1yWbFw1HeLz5Z/iT6Qu
//4WkZnJXYJVIhm96aqEtU8i9ewTWGdVT9iSDFv/SWO4FfhjWYkclvTZYHv5M0JH
BccoczUqVJ580L0r+6D1UlxjltgHu1Eb+FRszzraNF4Uri78MnpIJqPQipEaYXvR
IT2XM+NVpw1WtoDbtUYOx3Td3otjh/NhLyUPErNypSvFhdtvQOu+HwCCnrOQvMiW
155ofL1le/4FbhwEQU19Skik1qKxZDXWJjk6vb/SO8dOEbEUtB9eDvxgLWGFcgCV
1wcLwvs+Nn4gpxnIsxexMLZPttG+bZf6Rv6pOigVDOS7KCNhxm+RtA31YeuqSA6X
tKBfjWGuYxJWzshxKh57CGEmICn7DINu+D5Tg8fNDONvspFMOQ/ranmEjJEkQ6Ki
ouKc0yaBRDDOK26Ujhg97FioKFwAuhchCeETw6nCEgiKgbU8ydayzPk2+cpWZLfw
TNxfgbNR/kAGaxUs2WL/9w6x//BQ98bM8qB2h0iEB9WJHXtpSRMD5rs+m29GM2+6
bvUhuyoedleq6WrpXplREFvr15ZBBjceqxzT50HvuFHCYgjLfLCrNQSzdisQOeF+
mPePPSx2FKLRu0D/48UPfb9+x9cllm0UGZ4S3U/0qdILj/YWa3a+GJK40EgUp6L5
wOAS120FjNoLKRibMxiLgQjdWkLrCJiR/5G6qV/AqObIG7embQSXLxMQgVz/Yp5i
XnhyZtgFMxtvEvxSGgZme+eGzPqcUcFgn3fd7DjEGV6ZLqWG2QdrCWvGR+lSs1hr
YAGfroyfY1UZnqdSq+h62B5eOjWIOCFB4PwbiKpzGSNZno6DvuaMB4IWq5vMpr6F
lG3fUoR0clezRH/IAVE7Znk730JiExP6fCvo/05nT0FomMdkd/7U76xFze7QymK3
uBjZ48jsGhuRHeKMdG9TQ5Z/XJkVcNn2VaEUhESqVsNfgVb8Hidy29lhjF3O3v5l
8JvSlVerU8cw7385eltVGe3pKa+6rkJBscduvb0cAa8sk25Gk4l4K4OmQo95fGMy
+45wse1oEtMz5/Cj2A9Sf63z4k5OoEtNTRHser2YxttFIN3Wc8HTKpIwR6Tigzk8
hcW3C/2GJ1G+Lvy/Fe9ZitYB4vWsSHL5mxFR6McdMIZp7S/glFiTLV86s56vHTV4
0UbkikB4ei/7Pe2kPMRB/6hpWl1f2YaF4y9fnj/f6XkReHadDVDT/7b+MwgkxM2Y
FGQxVwgK1QrVXZmDoDOGKQG+l6tVJC8os9ZWR9CpCv2d6l/r93ZEfhdbguzyaCxH
p63knYCtf/dEUFHQl3EYaW6pks/p8ZOhx5SIDsv7c7rV2nrNAlUUFmIk2UCpEzH8
M70M0knvvsisxHddXdQKoowiuja9bTK/uakPqUig15TVEIEGVjZG+YocpfmLk749
NPKMp2CqVR60HHoT8dlOtqLMyCOBeN9m3SViKFB6S/xfkn6n94E2bh1VbtRHEK3N
U3yHthfNnB5nY9+K9nHinqxCrXUpl6Vh1KZuMfebgRHBywgvlM4DPZtNvQJIy2Yv
sqj7MxS9uHGguoiV1d0/ffxDjOTIIQTeyUUfR2R2afW1vJouFy0e+xxm9d0j0VBj
5V6sfreJ+pN1y/OtGCegUAOtPZkAQCUQbqRpb1AM1dmasB19xLYSzaG23gLzNBuS
BSqZrewxW/ziy+klQxjNQ7lfo+lp/3PT73Ca5NHCY4fmL9VP6FHMb+woXIBzzb7i
5g12YDsWFPRbctVnVZJ8Ygs8HnXbC9BniD+IdphVQXFu/U5wCtZL7Xs2Ez0LRFz8
L+CpW/vdTyMVhUDGIfnp6gOhdHrx0SPmnpeYxJg77IquF6YbArNAfG8VebVwmeJr
dnanQ13pTarDnXeeiETck20KMPoHlak/TmgSR0JNKWH1t2phPPGsGYL/avj7dz3q
4gAISayvM/vndXzg6euee/euC6GiJDSy8+06iVXjSYZVshJg3zbJ4TOrcuCmyYhQ
5X165NQhbOX3R6rnLJh4FXGjKMkDPrcIQBvng2y5fe5j/qTHx1NJHVnr85qOl0Z3
kqj3Eu37lFuLDpA4l+NRGKKZeS2NmMZdd1VFRH+B3XUw7/YXCbwwJszxeLqP5hgX
RWVOY0DrC8/uO0WdnsKrji7waADHUAAjK69iG06N2722DHuXLGiAWZup0eBNxRMG
E7lbEzPKqDOOPfMvQ4tEhfbFvgwODkIx/8UmcyhwZ2An9JpyBkar/1DooKaa3eps
LMWnMYOWrXQwll1Dq4ZvgQ1f7Ozd26dnoX7iAndH6MERhDkMkUIugVMQC+gP5fla
l5E814FCHCpfglNCioW/BAdmvEIl4YHYER44SQZ1tfdgKSyYCVekQd9hGTROOxDp
SweCr+zHu5frVPC7nJzs2x+SgE7+jkDd3F3JC4BBa8uKScfgkLSaEstkbRZkfMjw
nAMVEn/PLLyPeu380RcQuFu2yaEv5rIf00vuUz7AJwoxgkw63k1LlUuqq9CZHIEO
U2JbPy4VaJu0U3dyYIeEa9DimvZ7SBwmJZ+VdqVRX/6n0sS9YyMwdB15SfhWcoau
crq3aj2Wz+fKFw46j64fXQfnV2Up6twJnGupL9KLHeOKua71fOzx8240088qsp6X
9sgZlj5tp8A6Z729qWkR0/P40RhZWbJai2ZgZTW2x41BgusxOuqmEiph98O94hUK
XTmUTrgxNTVAtHgYkGF6B2POSVOulaq7bzuZnBdSf41Eeti52KIIINNLpmr0O09Y
nMysAuBREQjvgX4jJI3bA1p0FoeF7yP9H3QnNASiS7hJfuMCa6Z2UHL1V1Epz++2
2mT8M4p6t3+wzuqmSPiLl1bqiyDQJcHiceORLrmv7weQ/XNwtgvf541dNMiXcTqG
1ArAh5kCWcusFYr5I9Hk8MDtl7aIjKqiKLYasMDqQpUhEeqWCZ+5xtK33B58k5n6
hnH1Wk7c0CguM6dKbpPackpGfOSKFtUfouNhpE2ZFYBAafqkbRWoVw86y93fjVt/
tfsTS8Q6mdlV9j4PWMneRLf3+WlUzcdahj587c8IttHRIp10sCOMVeXXY9bxUB5l
9Kyej6WezNXp12U56kmWlnaUxFzHrxdgQ4gYXLLqQ0izv804l0Jaiq8qCdetsu3A
oiyJxr8nrKX1dOMgYmWW1Kru1x/cG0YR9QRX5F7rBkS63URPaWbN3X5dwGNxLPsM
TUu4/Ydmpvnc8moBGxgdv7HtwpGGEPjwgw41d649PoZUXmD8eHjNYPAKL09xqG72
TG0lf8NykY+aFHLJN5NBOO0qvYkoona++T2GSxlCz5soB15FG4sbeUTdmu7y33W4
L2xcgHvLX7UvYMFDY9xhqhmaTUA73YS5nr9NJyRQOImxqoL5leGRD8APnGZUGqC6
MWvAjZCbfy30D7hL+EHKPHn8BxLGdsVgI93sB7gNixBF1rnNPAPWmIo6gBAwjzTh
D+atpQqBTs7E4lSLVZzU/c7qIYbSLJB/zv6DcIpDtduQnXQ6snzk8hwV1wy9b2FS
gAeMZhSDf72Rh3SuGbH28v7jzPVck+V6wTawnpBXDLd6avgqXja4qQPFSLuTmLuf
JhYa4tnHwqwVyXOkZjMHIYrq332pDtjxFNOTTYECBeNEd68xGGXC1gr+nbQa5R/B
/JCSiIhVYldiqWKvXxsJO109ZXRzcNh6gwkBnAZ0TFqclYNZWM+NAg+LMlFcv4BB
VA5svtPNGQJqao5ZSCy6qA5TstaiG7I98MDRS2DxbAucLz5OiVYy2UD1GCOIqEYR
RrCWwBx7hn31oCPq5o6C1WkrjHzqVXOE1S7Rh0EqHbwqqzfHP0Sm7+2ACRh9BTY5
sVbsQilOYsjmHlpG8/xRzX86V3RjId4dgUgPyoF4ZqP6QzOG8xBXZbjiHALsfhBA
GyClxJAKOaMwyMZI4hNddPbngA1IO6XsIiO4FfE8Rr7Klzfu72sdM2W6gkJ3xY0N
a//hdlSrjZ2+xgbrKJRE6yzSEtTeQNzT2DDPHilQlscc9tBrHxHJhZEKyg1byvjj
JrXhTM4fZ3bBkUCt/TPJIlokd6HqxwaIUYg0ltd8XeT82BFC89xraUshB39Kh6m8
ehGmt7HFtBkEhjJY73W2DpKUfx5M53zMC4/xdO6bENMTPPiPe21RoJmDCdry3xFX
wMZ7jGvkxjH+Z2FaQCQxuMwpVyCMjowqNrRsVEnyY9U2m2DTFrdBSeZvu5ytbaty
jwPRJbHl7umXsaETyvbMt8X1CARwkg484wrD9Gdal3zhwLw/q1yKT+gxf3cMWyzT
Q2d7XmH/tLbXrekoHRs9yLvvvJvB/rXjfMqwNawrYYfkVPLsZO5DMHDtmOK3Dbio
L8JzArw1p5LxI8I/CGQT9f7IJk1ZfHCY/WCdmQEGOUOBSbUROh3Ot5jbt9FkaygG
UhjE0Hoj+uSmXjoescCa2JzZS5GGCwZxgFrPl4LaWDZ/IOLRm7G8vxOcV0by9x+b
883sYGACyIwfh6jqEGXVmSDSh9BMdpM2xGu7PBHW0j5zBBIGc+/I4Hyv+6KHVj95
tNdvpBARV8Uv1nGBl8oqyYE5dhCsWu6Ir/x1UsQHxefscXaSuYTFMUKmb2+hdnpJ
gFHpOe8+4SmHUCiZu+CDLgiuLd0TViZf3GOmGtGp5budHfZusTmvFw9JpaNL80FK
L4fRFO1Wys2zFANXHLpEIrr9zg0u0mjLsoJ3RcIyXzctts2LXj/nS5218qUlAF3Q
hzJAvmVaPNmAasE3duN7HThUl+jBHzYNT98GL/kO+upXMvmLjLUU+R6D4qF+RX/j
Wm4/jFr4O+dIuqBhkEJAwzTNxgE6E8++GjWlhfouYW1Rsn808IPKvrSiaFEumKPg
hP6D7k3AArS8c0TxTldBp5P63OlsglgPe5xQI7olsjbh9NS/ADGony/C2N8Ps43K
t0KDg5EUZ7sp//wd4ucDJOux0qcVyTR1bJ9ziaBon9KX9GjRbXaiZ84YoEmAqPTI
K8qctAsj5nzEGP3SPQmAOAoEqzDJQzyWkxLMaj6FvIScydbEUFTwgDIO5k2ugGY3
76tToxYZCNNfnwDrFCOayuNdt2LsU/uZ8/aFvtskVgRHn9U63bl2MuVCHK+MzaLv
Q9wzL4nM2GcAar37jDyl7MsVjtKp6P9wZ/2VXHs8skvdQnsQmaUTiWmaGMe6niUP
aBC3P3wHHhuwO7LRsms2JQYWgT0V50xNKIvgfQS1wEklYp4VgEi+9y/Elf/ako4+
6TwyIwAGYUMEoEpH+7xEdOwRpVryHOPYEotQdWxTFVgmNFSDdppErU/Y3qwZz2p6
pTOCoVf45Ixm4DessHp9z5bhkPFNzQwFN2JaZqo4a1VJxW4gv1Gq1QgDfWMbhenI
15qKhqJqq2qCoE0m2ZbquEQgL64yfR9KTNGjzbUwiCWxNa0RJu57wWOJ7Iyo55vZ
lUGby4k+qKEvoXbEwgetMziZsv5Cc1F16Jom7qU2tBoo90J8AeGEgcb/DeovDOXg
FV+y++5761nB4NhmHpHsUx1IxzhhY7ev113xZLNlG2jUnbtNiiC6kLH7UNoF6Rgy
SPuiiWstu0ubA+WVcSVrY3+2DY7x0mAzRIEKoX9ZLSDwzGuinUGL/o8RjfNVA3bm
EKKIU6BoyI6C9QTM0llREZfs6SVuBgS1Oukf+TfLo+vxJlrrYuWOAHi52npUmmnn
bARL/lT6lNUA0WUFIw0Y3yoxeThQXy9IPDKChRzpudSgJixODNhDcZxqD6saiJbB
S04l3brUWGF8hcoaxDBO8xQ8GLKVgIwoy2HVu1ch0k9VMaNTEniqB9W6lpOfv3J8
Zq+UAd/QyjwfN9Abb7x2JGvI1KTHe/5UbV4jvyTv2rkh2v9FU4KO/74on02hWigM
j8rnTM5PzP646/I22gJ8eQyQw4hMSs/WR6aot8TNMSWheaNa9072hzTZdzqJ0+W3
mLgjvfhFMawTMKkO/wA+87akOcAhyi4WVUoMdP9GeDiXzQF+Cm/5aDS2TKrpIZi/
4T7iW0UvAujP0WvYYS2hyWTaccByU4w0Lj+MZNAsOpqz6LMR7/MLHRBcl8nIJDmp
y1T+iCK7r3TykNC4WlXyXk3/ixYsOJWD5E5Jh8La31XhO2Npd0MEHo9I+ef/OTyG
IBoNZEeudk/6zhUm0K4C+r7JCfAqtHfrDVEWyyHPuISQDxXDmogtM8cxRbfQfF37
TMgoyfEj++4kW7BV9jbwOk1+666ZGqbDSjbDHVhx4l1w7dgYzekro1R4CRLQNcL2
QyVvxnuPY6njm18EtRqV0ywKSFDtNw837Alp+cxryerooJ4Wpi/v3Iwt62joCiUf
38qp6pvXZT8fGJQB4ZhBiTh7y8WYkpGGgkr42Kzx8RH0qPLnoSTFIhINpsePnnBM
CVhVzR7nj6v3dR4RfwEbis87O6Pae77d8h+BLKworFVF23wBcwDTaXgORXzUiyh0
QBMWDhs8ec+nFRcmxsh0YZ5ewR2ZRzbDU1SEEK1u7m44A7DGq2hIs2RKioABLifb
aE7V3FuHBpzN4jhtF2k2b1QLplb5GWj+iyBnnaw5OARDAmpdTvRyrrEZSpED7YBi
T3ZBGG49Qcp7rwQascQM0hvHN34HbV7SP6d7XV7K/pxROfOzQVXiH9DtiLmFRhPl
xK2N7x+qOvF9jJ9KAc9xDB7K0KhCO/N1u9G/tb4MCg4rIP2vdMJJMuL1bDcSockq
I3cmQJN/8FBy4Z0TtXtQvGdv0UuFEHboXwFvR0FbFFT3OWFNzyy5cOdWu2pi8s7E
WCorg/VCioti0+q/chB5uSEVMBGoyrl43l54N/mYoH6GF8ueRj/b8sY9ikiC1Mud
unzA5z92P57zDigrvPo9qMZ0EGNbKrXTS5n5kqxVl8tb4qhOgbZliScHahVDbszs
ESIxSy8l+3CrKvng+fAk0Sdp3xStQqPJAbgtmVldOSKDN2sNyroN82t/0VyjSUzF
V5xUrMMA1sZd1TKVMJPgTgqEbGF8lMDQ6hbyuxujvPrgXAcyypwzctGyYTfDHtD8
MBMfyqktQGEREqucQsoOPXLCkJBsomOv8Afdqu1SrC5g8PdCp29nYSVjblbgLuVa
g8Wz4HZkZfYSt144e2SYFi7iigOXiK+vQLCqpQXpmjXKPdgmVIJRup4qUHvFQ2Bg
zl5y+iyDNF8WaOEwP24fkWmJ2PWymHb23VxxglBF2dsSZu4hf9ENpIPXf/fMLqw7
Dav8Tzw6mKMdtNC+3R5zFuIzPHddFs1HvNESx8jmK8Gh0G21HYmfXj9enuy+stoM
nh6/jVg+V9zID0PJjhKawapiEU9FOGlP5CamHQ+PEJH95/hw0Dhk3OnzD64E1VNV
DW3UM+0IGKqteXa0sCQifgKJCyTgP6JJ7QlYNO2nhQUkeHjylfkizaHY8sJLG6/H
k08Y9O1wjYAULY7n8SZRfdTojQbVqhP+1XKqHJiiod3jl+q/2eS35TME4dpxApES
tGpL+kry/nzNnq+QlrrNA1Bj7TkbKt0TQgEQM4/zwMBpM+on+/dlpFb2jLQYLZBx
IaMQvKn1oSYcgybpwenMoY//f3cEXda95yGSORdXz33KwyzH+WACPDQFXvZRPvJ3
XTM5X75mSwqqMF9yjp9vH8N3lwu7RzYA2+P0hjvi7AcuRIRo9r9CgvlLvRkc39da
BjzgF1S9DC+FD0+2RjsRMpSNm0TROU1ocmspnGeAGUz26tr9g30+i9dtmOG6hFqm
PFHgdVgw01ae/ydt1gpgKURA8WBR2CYrIsH/CPt1VppdXQjO3QYuUZgyPdwz4hww
RkCmlIpnC596lO1H35GoTDen6GCk2iaPl5Jx/rZhXbKV3nU3pfC+MkyM6kTVYiLi
t0Re2mMGqjLHjyBZK5TohnBK8FVog2t8W1v+oq1W4es087Ia52s6s8w2BKwa4Mcw
cGP+LZ7I87gEu/M6/sn8QhnsU6KyjfF1CpaR4D1WRE40ShV+02RrpLvFivksSEv5
g/CTOXZxDqz6NLSN9nQdNoGWLc3vfMOso0F3L0W6UM/wwIAMOyjd8ecQXy15SfkZ
EeU+v3dEYtp/UhmDqMjMBO+OEhugSVWWpciyGKeZhDpJe/mR0nN8jfWL/eWYxqSP
cd6XH764C2xCDcGWoUgWQbnTwLJDjGZkSgKjj3+Le1kpfCw24/g+RwvJfiw6vNlR
qYg7o5/AbYsfgNytW6LU7AVkZHnVnM+Kq/6w4ntrq7j6qb2WaFHtJs6MWa10U8sw
QOMfBPOWS7maHwXOgPikHBdHI49i9LHCDyjtw5Yd2cRXEJllH4jjb+W6HliJETYO
4KEGGPddYTbVIoFbYKiVbXABz8CS8UpeUMHn5fk6DtIRneanBTttKb/bOJTIeUSN
K0W/Ft8vfgtSE71NhSv3RdGpfz9mdKq4JK+BVq8eIecZsUVGImGK8BNV5ocES9+u
Zzlt/w5zWZ37dyl53m+2gY6RoGb4C6DlU8T446X1eiZd+uic9uFTjK7fFFb84XCr
R2vfbffJ3RfUsMAi7Dse5Szp+ovbD4RN/d+lhrTf8UNl8lS0saTfSHE6FEilDcr3
EipwDQ6QM15q5CVnyrdJLfmrPJyqh6SJ5V01ABBi+qaNGH+QfWHIW9Em4UBY/pg8
HR8rsul6J9kemq81Arnqifn4wtIu301wdCESMkLzhgG+mamVQfbPSDitryoCiPjL
pg2BeqRIoUgYInSfBxmRrbyVAK72mzONB+i24cHYLVWv3hGCGcYaqoyUYY9hGTGW
WAAjymtag45evhj44bJvH0Qn4tgFNqPzDUzFVyQVu+F83sOf54CdT8OexGKewcs+
lxlZ1qydXqmdOdLVWAlHymTtV89wBiJDZOufdOUIpXgA1kVrhHknocnt2kkZzJaV
gZY77wGaaCiv96wEY+pYi8sZO8YVmM/IIyyVxC2D6VuJws4ntTE5ndIKnknHyOtW
9AmBXsNc77tb5uF6DZLu+mW9CC+vqvt19ptqqemFmChZ2lBmwpv7IqpoYSoPgqdK
hpg9va2lFtuNDGZ4fjcVTgijhKam+Es7r6q4bU+dJQCWKsM69C49o+bxUhywtmds
CuvHgX1doEVnN1MinEZ/6em3ZpUFyAXTO02biKva4f7wKJN4cU2q6SfkwYOqehcH
09LtNpmQBlZvWe5+Yx8QyB7JxwCFyfgAYbLVzs7kl/AMEn+otz0KW478diFLg0fu
L+kVByqkwVHfRsLyBUcGZHQrAA3joIkDFiB11AF1jgDMuoyaQwR/9Ki373rr//gp
aN5NR4FsB3TDF45nto+Z6rga6Ldcc51aQfBWpZETyA70zcDuPffS0QHxou1Kr4PI
EpUYO3enhb0WohbHdA+AP0lrzAB16FoFKabRg/3SaBFs11BaKj77iHsmHdg70it+
RaKzSLYmBt3WoucI13fbCAUEPr7UFc0IpVhRvXy8Hp3Af2SJVF3DskQBrUrhGXS0
oF4Vzow6n+9blzrNZSsRejRntT79C4wZKEDRHOBpc7E7rFFcTlfXLiNo2PmLkVPR
zBJDBxYcU9+YA8CC+gvpOwCGKZ3bo+x8tOce1LmxCFVdjgkiXW6tqB+/takS5Cjd
iN+aU8fahktIKRPJMPyE6csAN7sSXwiOII1QB4YhH+C158QcnhN1bTgStHpCw3me
kzqx3yb50x87+9aloxHSLQWLxdO67XsNX0NHfdmniqwqdsJHaTQFaT8sU09Rzels
JeNTqoGd85C2GyiXK6+525LH+AuYuMM9CNpAEcFYHQXITzw7xLBvFbjLIGKzZRt0
bNA5/wHu02p2v/wIYvcPGr3Gf0CM2M4ZfAPmdoAXyTBFOsJWnICFkmZCr+lR8ldY
fd8GuY9MwrrxaZ2gQ9taEXtV+0o25NsRcq+/LDdfA1xZYljNE7aBf7GU1njW+qzF
izLjnVP47fSxQNwvuM0Ls8sSe1W22KwOpyNfQm6oLWmEvfrsoMHeDrPaxJvIiZGh
StnkoP5Sw7OJzig5UhHcMqtP9RapOImK6jBQb/+/qkxGP7pSYmsPVsjGftxMC6Xs
EGph/vNTZ82jh1tVNykTKCMxeyNJI1d/WHrLjl5ixK/ZV77tNBksWmDZSqR7LpsV
0x0WtDe8VX6JNGyBoglQVvIPx3LBB8eT6NSF7eLhSE9sc2plrJ/gAmUYjCUqzerw
ToWbIpPuO/MA9loBEenlmFRjivFoOt+X3qydpVc5Ok2L6v/vKh+qbZ72Q6A08Ah+
8ZaHOG9pPSBp3jJnh9UiAql3pNmka1tQkjmuEWI4QQagpXx4heWygc3YZKkRUQDZ
ysdmwlXCfynXFgZVxn9310HqoJ6htjYUYjB8monmIru8WT7oWreWwZtQT8EqOiFB
bvfRQgSVUW1W8Iovc7nVNoNXZfQuJgwqZ2xHBY24ra2w/p6L/6kkibQhpX+rmxh3
1mktAOX8dnvLOIOx2Bmdqhd3fSTzVO7FJZxcJJbV72tG14tL166U746bHUy6sabY
hOl5lOiiFR3xWuE2msuGRQcsztMOZMZt5XXxre6qlX/L6nARJjrpPDZMKvIPJ/tR
z6vVJbDWTB8hSZTRG5y6sI7XRwbOysEpTRklB7ZGGarb6OzWnJZWBBc+UFkiRw7O
Psn/b3ulrsdLR+BtQF5XMVedRk5pBc1i2u3Gk+YXx6Ivo6aetQp4+Um9bPnc1WSw
gA3AEJw3ftMK1haTr71AfuiK6QjOmzoDr2dULpFXeUr7sk3/zDpkKmfs0NbgjnsK
swipuc1JMxx6KaUrKYxGxm63/k2WyzpPp6ScW1+bCmk/SkXDTJq7WMbaOUs9O0bC
XDuNlzrBLcXuoTWnuFIjnEiDFKiwKYb+LEmYvaNVyGXd52lyNFoH+NiebfjLHbWH
RxjCNWIQi7q7XenEygLIOKlVALP6Jr34oHxUYQ8Oe6HSgneF6vIbREmxNTBCgko4
UKi+Mbbv2sDZ9CNrWlDeKQNsgf7pmKZhD46ak8JQWSDwpfR6tmZbv/QOX8rJcR9Y
KtZCNgywoZj7PQ2zOdrMj1wC6KsajgEqsS/o9f3SKC/VcJJHvZVBatIXaGCCSQHM
0Fu6qGHvSyfEg1BJWcTUpiV5TnUpzBpS7cv2cleztlnsf2FC6cgiZXqrFnhWc2Z4
fdek4YIZn74BsEAHH/slUX71tAG6qqhj2N1+SVue48PzfEbebfvdNbR2/dim+a/l
v4cQMSKq0cbdyGBS/ANw4UOoFvt3j8v43zkDDHOI/WEZTaq0tOv1l5dSK+pnxLGD
1DoTCWZoLK8iWSQK1B+tDENfB99HR5SancPDrfv2dXyC9lQu9Uh/Ycv31A4JkQz7
RB6gwpEMODY3NqLAbuLjLqB21kfSGwjAUdrNCIf2mhoiTDFH0RcR8r1EqVQXsfZK
IrpLbsD5EMoi6/KmCFykrTcep/mx1Qgg+ZosXhuMPqbEV+j79pldS61bcBKyCxfp
p5wpb2VMN1MRtL46JQIErFvvTUzIh7etGjVnLcU8hMq0yJIosy4wpZsIKBITIgc+
qH64hJOEdHM9KQ7+9hkEPULlkw9GHCH1VMZQHjJX2AATdCpU8vZcjh+u+/8XunXi
rDEpjMQIM4l9J/B94NPkvlNByqKxPXiEoeCgnnaHohaLgtUUMCBG2ts03XgPrZ/s
RCUjZGK75Sn4E+6WXXEpbifWg4ObonWNu7lZaYb1C+hW8pc6vURJTJMJnpE+FGUM
iv1ZCTs2zDQI4ACa4IVc/+MIw0xqGzxeZUbd4WapR3PExOulGup+EVaAYANvzPZT
QFnhSyFtUa7GWZ1sUbyZoZBLbhE0KVpKz2VNYHZgrXK2dhm/u9V3eEZnhsp6OvnV
c2XLM+5Uq/Mw6nt4QdvZBi4P5weIa3zkHFSuGajv5WbwLBE5x2kEkYxUuipS3RlT
hRWn40mFQp2NbEHjB61eYKIpny40HrA2aKMGAXUqKKBLdI91RKRCUbupOdpQk6SI
FGd8/7Zj54K6TBhaM+R21gi4xYmuJWseqXJVMRvgq4nU3fovYsAr5uRGGIiF8Oay
dn4GqQ9GwFs0KSuvoiuzFrnQnQDOc/8NrtXnZAGVpex0yEGparnT+pm2Vgob0tTJ
WbN7+293XXt0hSM6uh20DDZTpw2mV8Dt2WjZ/XMlAFlCZPTkTAdzn8YVVurd1Qb0
BIJqMQ9hyhkgzLIMNmIwc2h8bJiTzn5jYA/5zPYqje25BYdVzQxKtBOyarhSJtu/
9uvwR05h2eYUmaLHHKOh2HDFUq0kk7gOZ1qjD/H17zf1rEY558nQYVxicDE4P3Vg
OO9b3bQhKN+34WHDN5i/fytR/ser+tvPlBhh0ghE2tUjPTfRp0dKPOW+OhAdMyH1
ln4a9QsrnwQCM6D2EgfUuX1yGcX+I91FgIOe8y8XHShjPTjEaQFDn186iwY9ThRt
8WaE8wcIG9KlAB79ihfVauuC4FOcEN/wQyBteifGu1L+xyOmZxwgxSqd+z95ZD8+
lQHc+e2xgtc7Guit9j+cK7hnoK0JCZ6lf8yiAf3nk39jwSLHn5RX9iZgOiq4XLUj
qqLbUKudjnGuzrDKL5+WALLHBOwzYm/UQdv7meyixb/1l9MMw3ds72PlTdskIR0d
3pm6erUSbG2gsMa9D9pq9jl2GfMjaiaQFxVqf4lTqh50XYjZOAkXr32kcdink0pn
aB2puDKaifQNBnm6S5i+3ieNRmg5vJtiHBGBHmUhlt+yYqmoH8AoZS6Xa8Qb+wTs
/aG29X+sEiVr+pIZ0HJ5Uir5YBQDR/ni3TODQ50hCqDYmuqnMWO8/7qUlGcPi+tr
j8L1gQ7U/oBdg3587VJ9dkJ+qDgmiPIDb4l950gy+++GxII3z6y8FWsqYUBvJV36
+98DLLS1yrfC2NuGGR6ChMANTuq1m9rt5iuroTR9APGf9BVfW67iQeGNrkWghPwT
P86HQ75s+aWJkjjleN4M6kmexXks3Jfby6eNL/amUSs+unGYqpWwudQQCsHb6D7L
B1PXWVGzOkHr+JNZG4G61rk4S8ahEZ5HrbCjDZytYnIdTKbQGiuXZVdZyxIE6yvh
WYwpnkUf+v3XyjHrakWL5RL5zLXirsPNA9NkxhoKD2NjJU8O2jA4atKf3sga7FBp
IJXq1T9/pjSiaycTGc3nHhF3k67rPwOq2Embbb3d6FJLXR34xvJc8J3SmpSvkQX2
5IK2JAr0cZ/TdWd/nYKie0PdEnZ6+36zOj43GhtnKPrN10lODnGpquW+fyTbINjR
PceJ9LcR/5rV1LJb7tvsDvBcHdIgtndqXXXie5/+LaUJijFpWbe7s6wSBHg9NX9p
qodQ4bXMt6gMf5p/nYae5cX3RhIpLnqP9wLnDTYEmiG6KBG+DOS+z2w2V4u7k04w
Y375gIutrvgmeMkAyMBXwOGbVmIIiuLTZju8io40Jz4wRa31vuAMBBxuuVlOxSXZ
SmnyAwl9MfeWkx0EBHRxthS/qiYvdgAtjMGOYQNgD3WtFS7BLUueQCCZS6+rfVbk
EkGqATNN9H9FbvMclUDSpcxrgD4K5jE5c79Su2u9rcqR12eLLHrMpdqxf0VjeU7R
7VZadW+wfllIgwrnJ7Vx4V0OW3W42eDTLupza8Donv0lvUCgPC7MhkIqhJU/FGOl
pRANTK3mFFz0JjkHQo+VaZFky9T+v5Z8J9Fmocs7qokDV4DdSdSOFDuetE/s7Dzr
KaNxLGP5DUTTU49mfDO1WS0EQEy8HSF76ErkFSGOjJYJx0xXl4MrZRaphlZHyKsF
pzZoaGrxt+dp7x1v1//BgVopCfABCqzqoeM2gJ5bUstkpx8SHQSZiYxC2Jp9CEnm
xZtexUFL1Oo7zZHPd+LwNM2i50aKRuqxFxW1zDgof7FU1OzyQ0nTN8Fk2lsOTRAM
OBOM4UiRkbqTbugxZtcQ7TX7J7KiltiA+Mi3wZfAKy9YZv4O2WPd6Rok/vAr3a8L
kC8mkTsAivxJTIYY/TR+7cIreEfcMJzEqhqd5Ax35w6K5YfsXlaMp6c7F7484qeC
s1Qh7Fl0qbw/rckRl8GkDg5DoOyyDkBoP4U/sMrw6MDGxa0Pdw+ZnoAp1tRzBbGt
1Ieuj8lfAFLGaOdHSe2q1B43vxRXRJ+WfXhR5Gy0CxXp15ywhQwDKre9tuQE0NQ7
IvVF94X/ibmCaAfQaObULJ/2LN8sWktoKEhMCz3neqwrto8f0+pyrV0jyzjTGSe3
tBqEWDrmoxfWGsWd+pHvhMNpBkajR0jZpBpV1g1HPbBAwUNEi4Oulq1/Uizf7fNP
9kA/ZiUGmE+zEtAnmfk0oGAmpfkYn+3RjBBWE/cmGC43M015JrJEninXrwoQMBSt
S1uFkJsB6PoXig/VAtRklOqwvRv+N1NxGdsF1pz9cHUzGPi/O6eFJ8qNEXMy3miK
pTgO0NZ4vs9Cyi0febJCI0zyhDcItY4YfAYU8IVqs72aW+ufO/YXOw0ud7ZHuNpO
FNtIlCPKNLqlA6mPuyG6EQZo7BtCTUSHaHNRuOwbbiup3/dPbA6DZTOGGYMiNaGF
SIKPHbvKk1Ty5VntRV2jVH7+S1oZMn8PDDUEdN+xlHdI2EdQOJiLzQy6j+DXk6vK
UWr3ZFCffIXndV0H+CTZSoXSfM4D7znAdpAZRaSKoLjZgaaBq2GNDHV/JoS2NKe4
mXiHCqJNfvGCzQQdK3NXJ0TLodmdRk1Vnvm4yF263MY9AGrm/Sw6slmjmjVl2U1Z
yZr8aj3mzYrp4c96e65d7NqpEohbBf7cFExsZUW7hN7HReSh3m8j3J/VNrQ7TiXY
eytJttZJxMwjcLAjpIrIwZmFVwo7QlYKa/MxUjme2Ms9IQqqTxxmXPYKESx8ZtVm
DzVwTwpmglPvYmim4hZ+c1wXT2U/GmpdckWyNVDi8XjOhaZc0qZVPF7zgikU+SeE
wGC+YZr6TVPmKgL7aHw3gFO49R6hXmL9Xed5JLbgRtSUrtya5pyEgrMcvwrHAXn3
n2ttl/cBuuYPoTgOjHi7c1tRABjwkVNRd1GKKHt6MEb57tSDG7CqAAys5ait6Yzd
oFaKKkfgqx+UT3xpvP8zs1MeQgwn2bv3kHDH6y4qObM6/vSbIoUjQBej0Y6n8qTr
pnyzzY7wxZ+QCVDa3qGLq1uyvy5pAwo6eUnkByFEE7MCnqfyKmM3hi2QyqtEkxRL
fJD2KbN1vaczjlZ0IbPvtIpr1wSQ94yglK6a5TjycVA5LH9gYlQ27IB9xY/MUbSe
gsiynIBt5clEgmJgP9idQJyrcI1rPHoxH47OI3ZUbXlRJ0QROtqZ5a2Hj4Dxb9Nh
OtlG3bh8IQTIMrWVDsWhwGe8mKoTsGf2DB19/70bKHM+mfLpnHupGnSUELNYi63s
SZnFj3U5UM3vVN/FGRlqXs9Ee2WlYStNZpk6ZskVI9i4+FnoSRomk4QD6GyIfJyX
zrij1MvR96ord+v5IE4lag1PJ7aZI8191Cok6aZu00rsyeIgNAEnuLD8BWdQo4iv
5MGOszAPGlGiqt/6E08UoYmvYF1x1zWSB3k8f0YlTwUXrGYpo+FHRzMHy1zon5/J
rd1Ga79BxXo6Z01KHfJTAhXFt5jfhZHVJDL3XLvX/Zp3S/SHEMR2H8q981CsXtQ3
iab7fLMIhiFr2YMLoLgAe0GAp0FTq6Ab0J/VCN5aIsHJFvNfO9QUoXbWetz4MwI1
J9sMvtKL8p1aVJ3mJXEgAsTC5vIziTHqBlccPxUkv10elSnc5PV9LPhwshYeuptq
k2hngk0dB8Mt6crVmOWltu3t1sogCYliDteUy6h95qsU0H8S0mdHsRml1TK2u5P/
AIyi/s5YhIGbH8Z6clW99tf8raoHoCjoHBJEOK9AWU5J30tVUBjRfr+CtA6/4rcP
4FJ0UPSuMEOpWOMGRwvLULTtNelxXaoUrZOWU/cDJ7x13Jl8BjVfI5WAMtaXEFbG
EdWkunjG+t611qAGGDnCXtdiLL3+eSTVtYcZHxbpWq2x7ZlZ32Uxc2j+GbSkgYzt
JkYKGIzwLaU3LeZXcz4Q/mdNkZU8mSxeNcou9J+iPV1PwxrG6uVxuyw3wZ/dWSI5
v3fmE3UkGPxdym1JprVlOhGStpxkGFtKDpCJJUsR6zU2Mj24oS784dd6gLdPCmsg
nGNj/Hq9Uz461iPW4XBOLj6WkeLKXgNvHOEe1yxgA+JXml9jRfsbntNM8O7MtKz2
Qt5XeaMkY0wx8adI/iHOw6qb9Vdr18drpNvm/H++URc9y/8ttI9BywLW2H6XnlsV
4mrlRfwP6FyPZB+C9kTuTTbTgxs8tuSl+xZBMkop5Q9JvF48i95W7kX9czE73T0D
8dVlxF50g00AlgGs9rgH2uYfXDTyypkOOn2rv0WToFFWRm664Cwkw/3P0G1+Sk9t
OVpu3N5xlHC1sLjJXT2G8n+K02N9Ecbrjqarf10gy/mYwMTPS8V1hXzZ+W4psx0D
sbvrI2twwwq9ees4leyveaxT/CgqAOR/YlOSIlIyDgK7m7NR4iFxCqq/LZO9M3V7
peyibuHx3dJQGX0Yvg/TGyid/Oabm1Bu8naaHe98468jkbDoKeNiwZrTgN0nPdbw
gteb64HRvmQCCuyeMuwN2TEUTW/mmhkbnpZ2kw8+3v3kAW3LW2Ar3wACYMETXo6t
Z/aBEoo2tSFpCNG3yB81aj5ENozhff3VYeI9Cut1pEiD9GhgXPC+s2cHRpMjJsXX
/14jKJxkJ1uEoFgZRSkIoOcZu0QPD9hvzJKOXzesVKMAMdmNl+fVKcBU5N+CXQ3h
7ytCrkcLjTj+RrSmueOU1AKAUr+hiodgc7qEMSu37z9xSO0Wl6iz1Ys3Ir2CMzEg
8XXGioQn8ofh4o920KCQBvQKyYqiQFIMV6gjYx8ehjkqil+eZevXe2LDwd4rK4zw
Lpo61eV4+roCZrl+jp5+VDTvT19BTbihPD9lFJ2ILS4CfK+/Cw4GSt8IqeV7m44l
klb9rgBCo/1Be4RuBpS1g1cl/84caCiai9hMa6JVlaMn80Mz0UgBG4nj9nCwyg9C
wNOqWB4OI/wY0UU60Z/N9IG++ToSEQ6RLThMOU0FYV5y6P7u0iUF1YriNzmE6kWj
ICCf+GHEJLO8vN+tdR9X3e8DCKbXLt9xv/5nxdo3ipuUGlJaD0zTmZtV54+KkNOB
1zNuxjGxsayCYqeSczzJ2TbAnGnkmJ+8KCB+jeDWmbJgn5RA1o1vBoIqwkTLoSai
4RBNHyClc3IjkFBG3lLbP+J/9my2Pr3SuD5Mps/M+8yztR0FG/s4o8ennaOEErIL
jWpPbp/CS3VTNCnk4HhJ/PELVMhMZL5SRP+DshoOZ+ZtwbH3jXTrXIlODIJ2+Uxp
sawY1yj2uCfCyF5rIIpIuYK94S5sQq4Bo+nSgCjQBep3quUG0kwZokMMT3cwplcd
usVNkry0Bjdv3L0Ca28eiUYYs+t7C3hQFvnJK+SPgYo1lHMxQLhf4JBiqzWA/YpC
M9DJjqwrflwLzJai+Ov6o9LBVA8RDEkNgKJo5ODIohnWCi5xjwv0xhmV1arFhczM
0fbwfsPG2PSTikt/x8M22Ce5ydZARH+qZsp0+Gm/QppIaMDQKizOfy8uqB12RN/C
HFuIzXGGx/3ekqzg2jKAsz14iNf5xHHTjXu7X5M/iTU1x/Ebf/sUDzSPU+G8TT+L
xjFaXvKk9HS8wxjYlWMzRb5eryccUpjYCwwoNkokCG9wth8tubO1iWVDWG6r6ggN
h/b2MH/FAaJNVapMlwnW28Y6iCZzvtrqnGdIdpsec9aVVe9kc2ARub4RKwVxZjnV
iP2nodlRb5l3Wo1w6IpygCAdprpeZzWAzsHoT9JWgbGaicO+QsPqyiFZCeSnyhLE
Q8POzNjbNOnF6Ea5ipfPfb7wDZLaveJq/qOIzj/gI7iiKPYPlcIdqyN+d/usCNRr
3vrlUYI4mLwVkdPCbcbV76TYYdJKd0YxLRZkAVlRH9r87v3JTu0xFCR+fEzrEZRY
0R2vbXo+BEtjY3XMLNRZOamRcg6Stjnn5BxAV14i5a/U61P8BAgS/Ut29pUa6RFc
eQ+zl8yHujC0bfxjHvJW1B3tKqkYxq21WtnFhN98kzUwtjHVAIvY321lyx8v0zio
eQoc3oQJ/MX17PqD9wW97aX2y3wSx88XcLl59Hd3zes8t0iLR0+efSfkiNnt/B+q
zSgQyg3mHL0QOB4CkT8cgA/PDGwUNCCsTLaqONiZ5k3O71D6u09A3VTzKYkJCUmx
Pry/b3VpwrKDErWNFIGl9bB+jJnaNwncp7tko0wTLaAvyFuqFFOUv7S3qhABDmYW
3sYq+UOHPelwbytHqEmogXBJHkxbn/6FPft+TSpuFlNzoCKMra3ucxmQz7tBmr0l
2my/b692rcHI32mZnTfBCVoQgxmqAcnPwYU612BvU3IEI1Fc6YLKw3lxhGolXhYb
DBXubky8qMb1JfbeiMJkh9vpK/7YYwKp5QSyJsN7lxfDIY49Byq3XKxXjTih97oR
YPd0gBa7yCNCESmeTXvOIff5XUKs7CuzMDwnTgcFwi7cLyiYqjxuV3Tl7P4kyz16
HX8YaSikEtF4f6hf1mIPxZwcLeYbEgR7L+bi99xrrK2AEWSj/Emh5n4g7B6fPonf
BQW40MnM9XGSXybpOhBB+3o0BDyEqLtB7No7Et3BcmBmXySrIyUGlSsIojcF31Hx
W+/diy93wxSP4E1H0oQN41v0Uzp/+z0ae2UBdE5sU0kPUsM7R++OXl0LaU4dd4dX
ohPjI9YSKa0aklfvnlT5+iF5MBZUwuhV4Z8RCaOLsxqHCxXqMGQc0LAChPNKXnLS
ryaKpZdfWK8DNwsp2nxQ4gaXCZ1vs/NH7qwkpexJhkWaksyRK3eOCFD1TvK/yBKK
DlNJAbRgFp1/Dj0uPDlFUsEschJ3LZVH3Nxkhe5QRrk3HAGF3dOgbzzfVWnhI0BV
QwCdHMlgQ3D6/JKHICUjnBKgYzUHNWt7DR0sOBtxq6IxIextezFlUKr0h/8xY7iN
+OuCq1IAszJt7NrCkT5xwdbvMKjQ2xMuLF25TDGFRiuIg8zk99/XJiyLWeJmwwq3
95pl0UNhlTFaogMXre8VpMt/69PGDRwWFTOHV7jUGVj0ZzmqfsC1W+PHcYit4yBc
nRNZrWVWyLbKKF+R0962JGphcbecdG1O6SurJrH4D8DGLGnd81aX+0eI2ONxNNGf
qRU4jvDHZ6s/ZELSaVG7MOpVb48cDN5PhAlPO6DpaAnYkXcugCirU1ayW684cGeP
dQQo55ZvnAMj+viedmJNyHFchtxR/0LrP9vqTVFF94T2jNygRrPJfYVLfo70s/zc
PBPWAro/3+aUDNCpu56Pb1bTDOEbUSL07W6tJsbYnQydx/TifY9buUZ489JJNmqM
S/wrxeiyfhoz7tkO8+2o/1mSSm3RDroOET3Rxr8Gvwpp7uAnhFsRsdosu9g+voLl
XFGB+JvXgXss98VE6tmYsJBoYyVjhzHY2pJSpKuxKpkh9MMFmagkOvbxEa8N3Q1y
kEfzqaiNWgn4EIur8l0deRcEIwfJ8TUEokUEIBw1yX2s4w4KX0BItBJNXf9zTKre
doV6Ux63uNan8fVqao01llR2rGjKCYM0F3JhwUTHFhzoMqH516BGrR1/1OToGoXO
mcAoDFBL1z2/SlYDI1jektCqyD0TpoEz4ZRAN6ZY/VMhhUzJ1NMprBToKq4zTU/l
bIfm35YeOjKw5aADRb2xZFFQhdWZgSM10Sm5z68LfRRwABcgD18EWmc3msYYZTIT
ge/4KWLu0DrCEOvEGSpKBEcsOLyy0N92B7khJp8MieLRf7sMTJWC4Nbk56jL5Km7
RyjT9XTFJ/LjrV1Mgdcq5KSq9dPMIFpevswTYphOMMnHAL9KFMFV/xWtrZnZ8Ww2
CYMMKCGapC70PpDSYLCliu9x9s7+3IVBrwg2vjal8EhTDFY+tKNIj4fp8ZFC/OBE
y6qU36m3YTNrOTKnR+weNqmwPuO2PHRDqO2pguoWEYnSXgavMmjgmK1XI3vLXQ7H
TivKznd9rfQw9mJLINreT9NTTjv0yflNqXOn9VxID86al+B2pawZrso6cNVr7o8A
TNHuhC1KOriMoNiwcXCsohGm8W9rLrTUZHuS9u4ZqVa6tKa5pJ4Ecbs4g+0MWm6w
WEiFbektemmivu9UNLhGD/BCq4lpJYXjagY+A5P8Gxi0hpRyGcqjfjX0qPopn03p
8CmsITa75AucfO6AQkIrQwMEiz8FAMFGo3PYoX+kg1IRy6uSdOxydL1dGtcXMFek
7gkiC0hsKZJIW/WRnIQYYYsL6H/w1mt/p/xLQgbSnVeoe6JhQAjQAe2eEGPCakvR
8595QeqkVOy4Zfza30sxMlReXL0LzE+YU/tALSWp0D4B8vOH5aUJGeDvcg6mVUh5
wh1nnMZtTtvDi+6cdsfbW9DDF+9hMQX1ArUWowDjbIYnnIDdOuKYwBM+thCMn2Xc
RybTMKC48TqnQE9J65czUSpqzFa4gfktnF+8yfuOIG6TlG8NW9+z1Orz/wdS0K3m
zDB1Vmrg/D6OH5C1w90M382hMC9ACgc2IEn/BY/IILctPW7eWvMiDEH3Nx1K4zyt
GIec3XzJRdCn3qpKafwsE/yK+jo8299AbQ9ZcpSYoMGhyO+qcmsUMacHiSlfHSDH
5yD+blvnHk95uH23MhcADsRUOLGAXIpbtfAaHmt5xYxC1rCo8vHoS3H/Mr2ghgUP
vf3K9JAnmsMYht6KZKJUE/SXsAg7ut/uPK7qIFkFUfySRdzDpxG+Z5sOx0veVlJX
bY8v9JeE/ZLXXFycg9iQwD87kWBkCACXpaCtBg5maTLpvP44SL9YCyyi5CffnG8m
0BO0xPFoLWzHLHsxe4tW8FteobEOGoE9U65wTtJ0ix1N5CUriZilRGUXyM90mUIV
Oe+RmZbxDqonGbTsPTUL0hj2O3qWTrJI29RpQCW7FVmAJKSyPMOLEvQvbu2UBg+P
11GT8Y9+/Hh6HnvsqXHYlZgGr29xrRuuJCY0MhjNkgG8x4HH+9TikIhfm9bUrbAE
cBxyU+aYjIWK2YYWK/SkYNHjpWxaSSBzKVTXfjp5eBAXYjDVMA8rYrvntv/iYw6B
FlTMwPWHJKnWtetGlWq87BbIYtkzzDLgqfnV4JaTV2iCcdbA+H/TejUT2YnW968o
RVBm1TSiLDYYZGLvgkpM3JveCGMYRaZ1VQoeZ7aVMx+0SfUVutHVJtUIjUQ8fj2M
MkEpOyBeMY7piFfizBjmn5MnFKOTJ2UEayP+9DdbB2v4bytsaSKrlqlJjUVqBiYP
zoUxIPO/XZD/tQQDgX3HB6wW85cAQ2AFjvZOTjimK/zwziLvJfkVMu5VpaSCnyTz
OA1/6QctTsQ+VnruinHuAxrV2AzZjLdwsPK1cXJvR7TKfbu/jbCcEHEsp3miaBTT
2BM4Px3Z8kVFBWQ6WTJ3N7GzeQYBfCFk9WG5rH68zD2FaqemOk2HnzdtvoJTg6TH
7ELEdz2EmpMGfXqX4oBL8ZaK8MOlMBjk/Le7DatcWI4crQi+u9y/1f0qdGoh0X+B
3C/fNIDQ/U/xsgHPLViWGV3y9KVPlUc3G7XZeO9BkaPVdciVGcyGbMXYT7pPfE++
rnBKKrOfh3LBjPyYOjg7emwc0Oh/S+bSqe2K5nU/vVvGvPOIr2hWk/bQM4ZQzOTR
t3ZU4Ffr/hmkxGgShDI1G1QaJ0cWpbV/b8NQut7I284IpMNRY36nuYyVsCplFnOA
BHHqPUO0/ATIfoTGNwjNian/wtXVl75MpGcYsmmgqlMpzVrHAfCTCUs0E0ycbQKz
lLRQxzp6mI5MD1y95EG4HinWmQPq1RIm764ud4mfjKX1loLR9hl81nXiVYpDKHed
7xrSRq/Ah4xXbQc31ipoLTytd5ygpcObT9m1sJlAYOETYTvU3rhsfUgb6t7o+Rye
lw4ERtpQEabvJ6h3bSutyzh8uSrpi7ZwHpM3z9+nijoID65f5H/ymNCQymEjajW2
Y867J58VlzToohTPUDd5Q46oVpTFyNgGql/pmpNwgxOvCwCxjjh8Om26zw9WRTUf
Dky64IzEUrOZoEt1AesVVlcNk3ph89G8avVz78jnp3vzJxbAtxxO9ff5Mw8FMNPT
I1hNsJh//HXjWn64ApIJf6oDUGalW6OOY9x3hMM+KofpIGx+aGh0flHymAgDTGqO
5QiY5IrClZKOEA1IZIwBU7fQqv/Gn6PJwBbwM1L0mq6nSEfPBG+oDMI8WRZaGp+Y
1Zdy2ucZugSvK3JQnjZ4w63JZDURtm+XN3WlJk/0rNzRg5PYpZChXPtkPxWvTVfy
gn0DrNralAyYjaG/dipVxjwjtX2YNqAVBHG1HvbM+aEpbcMbl044RgO0y3mhJLiI
3v7MVZBDK7nvr+vwHjnFU0e3ZcHxduQfaaHwVgvyXwvlvjmdlmuiOzYlOI1A/p+L
5QYGDx9FB64anRvm7rIbJO1xEiSC/EvGMC05OKiXLPIIAKxONWfESyqRbIHwm9Lf
kx+8UJdukEiCI3e994Q9/6nzy8IewrYnTT9ooebLb/Xy6SFAlpv6vFWFfz3seTDa
uDTX2Dk8+0ObsCVza/oJIUAMtwQNqcQb5QgOXLbkVrRRYm0SA1JQM1L3RDg2fvk/
gLDJfj/tmk5w+1HmbUsEQfsKScrOFGtSL2BRzTzxbhr0V7dsuC3ObIgtkBm9ptmk
uYL7Lbd5FmEOsOE+0vNFgiK5aF828Zg1qQRtCHd4mEUQAHGDJGBsVRcALZUkNQFK
viqnUPFLNFPq8Xqal543N/7/x6aJ7hnSxbGueM3luoXSIu9dXaB4AkPT8iCgyH89
PeXq51ZwYtkMXnuTLM1WPZcXDKSglDdYpMVyGXxbQYL/AYhUkl9wTWyccLuQ6QVX
t2s9LCYEUvax2hEH6OgbFm+TdF86R456Uo0AYAtR2se9ZhvnPYdStBZrvh65f6Vi
6Dis4lvMvaC3sZjf4Jnp1lhuiOKDMoYBwJOP0UrL/Rzm3tIUwezns8tLiruaihSx
2skvEwPKVG4WE7T8Knsq8SbMX8wFIacjpJ70v9o3t5lzHViOAyepzlKv64S9PQXM
+DtxPdaOGr7Y5rKsjLcoJc3ta+dZZtIBKLsUP/tn5lK4hFq8rkRdrNzgqVpFzAZo
hWQtTzZmUEPWW+riFTugE3digyjoMX+ku8ZhXJfqdhginbfiOxaOMWX7NYwXuOkb
rLYjAESvLPmRoKgGcTpPhSN8NKxfvAkYZb6kDkjvTvm/EWkDzWsd51Nvp45ogM7L
AJ4XDovjHDHVUa65R9WUG0td4qRaDQ/mRsIABb7QJxUTn2FMbDmMh2WX2jkzrjSo
YtprQbO2qi8GjuOOmm+tjzDKtZxlAH4Jysr+BKclPatrzKy/4Q0wvmHDJGPN98zE
hkX6nAROc3GHHS7BjDeNhHWIEJZNeYPQRAgGUKOXeRCYKdhW5ImVWgBqLfku4bJS
NpQXwbn2g5HMjyYYO4i9r0z6nSA5Ne8/HJZBCk+We7RXczg/NZSTYwLatsuU6n90
Gw2/Zda4W5Yo42YfkbZFNKSlQZTiysHano2XpXzZFs1lG+lxPWkY1qAq3JvgALSt
075e4SF1LztyFgPhxWzyoHVtvxoR4JvyPMntBIHw7PnanzGjmYTCtJXkgwaFC6cP
Sue1/1YuVv4niqF2V+gS5OpFJktwg9snzfwUeLHEl4my0OyDSro4FArNp1AnJ2ff
JSbW6tDuZzx4QBadpnLpedTCTD5zbpz0k2JBvBbmkOdn7zqeSP/uqWRSOsE0vN1x
ap7ART4ch7Rrs8cpPu4oSNV51ino2GRrpujqwMuzxm06sZIfyFNsULnWvsDCvmM3
GW2JrgWYcy19JJXLYzFuLBlxomVqpu4+l1H5SHK4g6p5AhmHJc253mqyd0OpE506
qmgsWuCkvDRz4PoLap55+hCqHCDJGWc8oFzM3GIXE+tdABKVz7vXF9JKoYGCaL3x
NrSco7gOw/ITiCbY4KM6W/Bm8ritH+9ELb467HKttHwAEs7NMAHVYq+VYFstVcLZ
XP8LalvDTeVq339qzCRNfXJPT8Tmp2dfGC6IuxglJrxaNWAzMO37cZ2sCgcNgphe
M7Mf7YNObXao37yXj81NR77NdLvnqSv8nvrKKXYiN+lrvSVeOM00xjVZ20nEvSVK
twd5POoYp0mOr6vZO2DiJqdp+f1oxJaZc35JeJbf7J07ooz9IT4JrNhQEh89CyKe
M0OJRaJVwL0MceUs5yO827dJVTZgTYAHZOb8BP2Dnakf+6hjHjHObLZK76EQAmlY
bojYVJ/QD7sg43Pq60PtLKl8B2S2dvqilrHZeYUTsDy8NVZxcrB4Jt0gRC6XD9Ap
cOJgq39CHTOPrf6xX7ZKqGALMqQsEcjcCHR2nHKONO2YBwIBdwZsyKOA+htd3u5o
9VDuZ5Iwe+5YGYslsFWHXYSa2lu2B+ygIJhjuFQisMta2F9Cer/LXPjO6bnW9AIp
zBGHZT+ZJlUq06bVl2CKDRbrlAf746bA9E7B13PlhxgOQriVBCsMhFHfoQRfdfCW
H4aiveaRMw386izW08yAg6+O8bx5ZjyxqJRA+JhNEyxRwagEIqbSSMSY16CZPWh+
n3cJUoI+FySG1mfdGOwXUzOhLh4SdIzBTlicOCFqXRWSMF2aPX37gdQ8p+raes1L
dIugvW+Z30q9wGgyt3yey9q5nnyL1qg8TztW0QSQ1r5AbTMr4lcABxoWsrJXMX2j
aMLmb7/O8R7C16AxcaA//tAhwco6GA1oP3HZX+J/d9CR0nrZ9hUaE8kV7PRWn06f
J24Om9U5lhggcKJfwOpJaIhwyF0CQvx2nNBZY57QODz/+4V/QvvrQTOQctwcR9v7
xLM2hJrbDzU/vvE3IvSTsDrixTCA5R821Q6pXKZlL0SjK/x2Yu7urYvpWUzIOpjU
E62XS/iqEKcmU9OUWSwHnu1tyxwRx9d69deZdaAr4KyfaTKJLbXbb6Yo8ykJbpMK
HUuC1JoJOMgeWrHSIz2f4iw9J4Htmd4v37r+pzkFYgrVtX98tWv4uZgUqiPFg+He
6yDBqW2+FCVupNJICzecO1cJ5zFfivGMEgS6oMP1yz4I3NIktdkKgpTLihXfVZTa
XluRjJVupZkiLhaRW4Vq5wLu3QSyAsBPryULuSzRyR6FfiNfIn5G73VAHNCzoio+
IR/LJQaaLr8EziplbzAzAAkLw07W78asmABF4+3oekWJIMxSFiKRx1W3jiWUhLqI
J9f0wMakfCmJtF2nqjo+K1Wm3ZWkL6BJNb7lUmsUW4PqwjEB8z/kCSx6bFMJTsMQ
zmuY0SqxzkRJSpS2mMzv9wM/PRHMeZndp4ubOJlaz45ms0N967Me4gzUO1FunAfx
6GSRU7H4G61rngvVv6wcbq4XSjK/PVUyqoBSNcu+mcKb7OAG1iYIkk51qupufqV6
RA2dEDLiVT6persF42tm7KHV7NYxxGQTIYsixpVnR7omTsOl8qMs9Gw+4zEV5rVK
pAi6nm+0hXsDhu7xcrDy3nt1PSWuq+VJJLQwSEAwG7wyvAEjDT0qEf+68QV2iWxn
35C/ScNAYbj5meiiNQbMh9gUfLdieTN7Fr8cW7Z7aQ7QbMLP7U0TZ4YHSW7TiTZl
U3dmU4fe9tOKhBJM6Gty4RkGZ/+iEIFdszNeyH6Q5+Ue7MmXw+okmCzVOQkaSOXr
qoUhMWtiYsW+sSvyFjiXO0RoO+SPQYFwmrQkabxcNZxX34S0LeuJlccy2cOtc79t
TnoI8uEbuMnm4DTy+qLJbltxiZX1Pp5vbqP74Por7sUjqaCp0UU/WmVemqRpaiJP
Q0Btf42X8ZoqK1QI3uHOujZxx+ne56rtQcgA2ZeLpnN2FaV2aMz0SxHkd7+Vrk2u
0F62eJV2xmuGOTzfOsZJU2kqV8UkWeEsOsaj8spmGTjROcUK5whR3//iuJ9wfbLy
bccVPdswjFoRjzj0RaFeI9/qeiLdfIu63dTnVK9UOl1+g8pfpLjDZBj06+mZWqZ2
6LBX5RopDw5a1ifVg3JLYxfgX1PZ5eYwM8BNDEEgQZQNyP0w4OSvSSwKuTTs4Ymc
ALz2ZT3dxpH6Frh8PW+hydbb9DH+KT7FO5ln3mipOtCQxS78XxHzT+OVXb9KH1vW
XZZaknBcDmWj3cdg+Q2F+BCB05Lfem6isXZg6gNOf+H6TbADZc14F3mPEf8YYR0S
x3b49vFLLdjEJXVDdyr0cCIp5/vGl432cyDlZymOhBcyLidUy/EUNbGqVF0usxaT
deeD/Q/c8y7qHMdGZa1U82kK7lM96FiVxonXgQN7GV2h8aZ8Pb/gkkAONba1xotf
b2RQmv/TwMgMmPYOck3bwByPQb6hC6YodA2RNm5OztvdyFVZh/j4qHpcwyOo9EJT
71IJvonxkmTeN51M2lvCxrZrR2Skaa/ETkDgXODaHenmEF+1EN0vBzPrNDbYHbGN
okivxXNldnr19+bw0yh376TAcuayr55W6IkiCBFXREUetZPzKTvC/n7eP3fsgkN/
pvUe1VfohNB3fvPX6XuWrw4+ljQ8dXXmp+QZSt917OG3ls9j7hwCKkZZrswxOrUG
hC65ySJ71gf08dr+OP0EY+7ZUnrBHsTu6ADxG3TB+BlCGV0llbaiRoOn0nQ+6Sk9
w3l4NKuIAT5KgSjCgjeArDRs6MGzINkPgkWjya46YursEySu8UVMZ5fZhzuw1QMF
otEFiv+1cQeh9pxYEd9imgaOpLROvxP0KosAUqKeJeOjPtGTRRS4CjAaYfiEChNC
KwFsqO3q9ozsZ6+bYhuwGCGdx1PcZV+1ouKIjQ8FiJ1C2E31F4FhaJZpzbp4i85V
/REyhC0eLuJ9+gIPi3dTyRCho4NoxzsT4rZxqg5//VsZZsP1/REunFB6uSH+biad
wgLObEpFjRK9m6K9K6ORn/BTMR0vT6cx64iaVcM2I5cMlbnx6zI/O8M6hwlvm8NV
E49wLs6oUWSUJrXh4xJa/T2MlrQEae0kwVGKiLL/tuB06pHaQQ7iXOWWm0KaJBUb
pW9myX4QSEH588uolA1CIM28ddRxvEkk8kVV1EHQ/0PypmHkB3eG6XLJCpWljOyu
OOJ2d0y1Wd34TC8I/d5hxavm9gwL0eZzsmO9x1hfDYJJ7WkipWmHYmv0XZ2S9rkf
2r6MsaoT+FFz08QZekmNor80Fni8YEMm+MEXM48MAxtvk7Y/UxVPoQ/upxItmSpL
OP9a+iz8lMa9KwekI9KsUmE3neerXm7uq3YZEbxTn70x+lxtBg8dECjCmomC4xHc
EubcbRpiSkijhIlxGH3utGyidrRL8KABdbWmSadiHjy5TaJKody6njGvlXMhDI7Q
yxn/Tf2sEfn+hWBiOJ0eFeeXk5bY+h1prnm9ieFjxBReQwDYRivqMnHezbahKIuF
++0JsvbBZiacS1YhO9KfDQfVKwKFZFZPzk9ntYLOHxwUIr0nIsPxEebVgMakg5vn
nFbx3T/WZvdSjhmGwV109uj2z/xsr8xzDqKz+3xF16OAbPjSgR2DAeM9JIg5YOir
R0TDPLJa3V/IEjbrKL+1zuAkls8tsNOslrp233zfm8rQNOn4Bg96HzwH+XuDLxBu
WElofN6oUynPSp1vQkm8UqXenqzpb7t3v8hlJEHvdiBJmmGXRm9OF4mSr+Tkirux
6Ac8+aUXdmuhgxp7eo6uxTSG/7eNegNIkTCVzJ7uM5NSe6+bTjQIOjh7xqSk1ECu
7GceaJUM7nsCFPRX36BLY4/N8O4x8tQ7uWM/sTebHS6tjKCcvo1FRiFviUoWkxfN
dbMseMsFepfrxKBkmfyOWIa/D4R8eJmKtD25g2bGAQhiqtgswKB5jPWKNBV33HYG
k8YtNFNiaV4VL/PUDPGKIfa+BQPAEITZQYJ9tgfOybjhOMPq/9S5olXKyxzL0/qC
Ke2C/k3DeruHt4dMfDdBZpYtVEP7dvTvOoLWlPGsRUq9IecLc+4Gnp72qKZmijHu
7dBcm0AUmpp/QycQqzf4RpvBVq1xP4J1BHzpc4zvUtt/r51dSqdoD1h4TcTZyNaZ
FBp9Ndgh05U/RLbpdjy/L2msha53xbtxqDU0qoP9RCn3apCiUA2r0VygavskrHWT
Zho5wOdlzWI9yrYnUZIa3b43w2sqW263jiD8DDJ96Ql7lG/4yILyxLpO4jqEv7Rr
HZAXOFF058sArdO30eF91pby7f8JevAZ3DxY6MrKFBikwwvgJoUCSIp3lbSyJ2bL
z1dntxK/5ZpYBEW3e5H/SY+nGX23cPi7Y8hiBOjNYTu55RXO+g+9FERNfpafnu1n
s/n+pVs2cIe0HNUSfxjq9zQ88me8xrG/O8NVxvBa7qUUyRu+gXqvOi5OASNz8Ynb
10PFqJEF+25s0liAm++JOCF2wxo9qq4pE1/hqY14oVkmteWrYPnixZF4UVjqEIjh
bIIFQSngJH0eQ04lksiYQJW3rD/y6QeoaJpz1qp1maaEMVjwhQmVpZlEy0Ll6E7k
jypd7MmuhqIcDyjWAtrzvnI1xVSHKtNJ50KezA5EDjqWROdRsH+ZbZRkC+ITupY4
GPD52viVZpx//5aDUa7L83cB6dRHL+eQHpj5ao8QZ0hoLywFvc9BDOyEJEnUAf9o
A2+jcz6QBzwnsFISRJfBYLoBZIyNJofUbHePuwwjQmRDjoIxsoVrjB5etxWOBCcl
ZyvGgNbNdNYf9Q63u4d7oCvSz24lfpIUKGWUv5b6kAPKE99C5vZwQkhZlSXEGjPM
wC4uAMs7NZ5Hz3/gFUz4xCJz1XuZi7V4DcS4pV27HYKgj5w+d0FzQDUwto5DgLu8
pBp8LJYAU+tHBwH85UYvEi5iNwVaIDllv2YYWVHpvuyBSPmO2/wtlGnAzDA5t34d
njmI4Qi2US+BrZYhm+/OiXL0vn2xy+6mqrP6UTiZqzzEkoWTYXoRRI0radfEMVBu
RqH8eJyVAwCppyE2xvKarCc+OkYnETMmoNSg5qUrafOhSOKE+D2G6LAJuzf+MVJf
wi+Q+K9Ku6t81HUxEOXrOTowbj+Q+TVyndME39G2s2v15H99ngAzpGIjKTaUOXRV
rIH8dc3sERyAxphPo1/zaYPOZBQygCle8ALFnSTekv3M7av6HeZt2Kav8pl7pD81
6ZH4jJMTCVp783Sncu9Gvas2Pja/KyDU9iDkmrx3jB4ltAgobSc6WEb5doiwx81h
kyFmeAdLfO05akhGL/CyxDmNXq7zwjtDHrRsL/V3ffy0mVE+W7JnJckFdmoQCpKu
1Oks15A4pN2I43TnkPjQhZY4p1J/pjL22YQ9FMIqCo8MA8Vfl2rG7G5GiVF6v27A
r56YSPl77VA+yCjgsPY3+TpSbCSzavxdeITt7DvSLjv0sEE6qhhOFRuMAypxCYBq
d1A0auJ6SNV6CilTDQjTGlvxQs7vlzZ0dB5ZTm/G4uq2r6aTHZNL+ppqGPhD1Ypi
JXagkgAnjKkrpqomccGW0I0eFe161u6Vr1yzi1dsVotUfsbt8y8J+DwdbeWcpZj8
/18an00UilBnKENTfPqtX+gl6e0SgG2wHzeNiPCj320NomrDgm+tAba/6kiW3O+Z
2CEIE+BcejP0HnYhyAKBTcqAB31qS/wOGCZXX2nlWBIh+1QGWqqAajbl4pKm5Qm5
fOoNOYV5UGjUISmUGmm7L8mvQ0PyQJ0Y1FXm96OUy0om9XnhLaC+/k/IO7Wa6u6Y
aEzWxJLGe1LcQhOMpetV6FsZ4i/5g+vUzy01dAZlrF29f8sLc1XdrqHKG1JDPkCY
YDVQkVpSYs7KhKmNln88vDA/CjtzhsnESdrMCsltsQOfkut7PzjKt7N0CA2NLFwW
+0Zvga2lVVSAirOyXURFXM/mBHEm/PCZo/Nke+4YM7pEhkKgfVyiFeB2eArJctSC
y8wtoJ6hKQdaMoSet0vxwox+jJD0Q6qcvJtWE4+eTSPyaMAfS1feD+1PJtmL9+h9
+uZGlKgqGOrQWFpKfwwCpNGLhRrZbea2Jjl4I6AwnCWcfPKDrCugWSvfsVct7gBp
n+99ncAspj2T9ZkdeeqI/Tn/pxY9+CD2Q92psrp1eD9q2fZj+6RwtZkL9r3V2qF2
Uu5urz8UV8ShJjnFlNkxYXZwZsLhG/K7VumJFWjJ5hQTRq35PHYIWDeRQeNXHhCS
rRsCKmGer7RFOhZcDssQMw/J7DTeCAroNJBphAo0dmDmniMyJ1qfiUj41AEzjlrI
P6Bx9+kKqHeL2ZatEG4qcVwetsVmrs4lSFqo0rr4gCz3pliX+up89TUGfVBLbM7f
tZVVOGuK5Ekecyn7dX0P9ZUceiNH2h+qj4uALVgQN0mEwGYAoXJ8oIf3UOMtEwZp
Qgle4oO2PkYGQlmR5qAsyqQBzfQWalbNSrFJtgM7kTqfts8ZTgZwrFVrsTgTMwEx
KzO1hO7fxSX2XB7NC8Lu8vrYfPv97orDxd6Tv9KCVlQR//CFLpmlKQxBXNCKuBoE
4foOC2Iunzad7WJUsliEkPeDZngKRWXhWJe2Y2KG+8RPat2G3iY2+7DWPoq0LNbY
cNmOrjdFc/kycObDPcFnWrGKPrAJnu9NxIz3KcBd+mhcobLcqo5U4nJ0/UizoaZa
atATmSGE8VPIiH53exkB6QGMg+px9AuSjGZV9QD5PqK0ZystFhTIaRQZmR7krl5g
sE+PrU4Mo65QwkXJYajSNmtdxGKnD9Hon4DFRD6gcvJFt2TI+DCacC0/E8PhtfAU
s+kHsbmwNfkGts46cCI1IllvWYpal7B2AAfkXBZphGA9ZeRZjxXQecZdCzVvx4ex
wOBLEjIbNSuMGHWhei8IlEdcMimpSbzuf+9iiqV9G0ss02nsWhB09rt+Fycmhfe3
EKgpRLRxaGVCb+IpFu0u9t1Jb8CPtjPF3lirsra+ZtXOSsz0YuqHEj1LqXPGGW22
NLTgqGN9OtQqVT8xUmOz6y7/wVQHnJdlcWFmAQ52vYq361C7/OXS65HZiWCtd7Vf
dC5FpKPSc9/ipIORgNJ6V2eA+V/jc4Q53A8SKLjAvzosEBqmjFss877xqRMWZAPy
/Qx4KjANdtYggW7jtDz2hkSkh72eSaLS6lRj3QmDwGl9/T6heOKg6YJyS9EqFKG8
ZrwmHxN2ILV8/m/qmLPopPcKcEY3lIzI3jLrY6YbvafHhN1D1PaJVOC9FQl/0ILJ
J3uhmfzTBe66wgV/k+jZZHX8WQyema3uhYolB0sxd15I9mQXifxRLks+4HMoLLwz
KAH2L5Y6rWuMv68t12o9Rc/uz7QegsWHHIdoMyOGCzdfBmY4/Sje17owNhRCTvVL
NhSNl/v2hC7s8r/2BfIDPRAsJGd5R+ViFKOB1lOW4lrtLZYIT9xBMnBj9pIcjW0Y
PfTbK3c6iyoEzZUmKR3YtrpXYQCYZownS7rPxmk8JSq+iVC6uUgPgd1qtRwyQTiO
4c8jgmm4D2mr2xTqtCbCTSYzciQE8Wj8k5TlrGifS9tvoRSNrOpshRYJXIp6XT/H
CxzoS6i8Bu2HywVDn4zKN6fjdn5aFFO1saJnRBXh8Y+uUXtwfdzFYktHnAC2Dzyb
0IOIM28Hh1xbhmWE5mgxGHJz+fQfOdaPLbaQpds6TAKg8+rmBbyIK0Cj9eEP2X7G
OuyeFfwKIJG/3Z5DSzVWF3qZW5HS2EhJPihgRZ5WcvIpys1o6QWmforHt5a06qBq
zEFMyISepDUteumVg7GtFwCMjF0fVfGtyGdsTcuPMOkGiC3EKPy+lVxM9b8/P0fO
aTccyoPH9t3j4jTTQie9z6mhsPsQUVsQzLllxC6eY7uLJwjTHw90PLmFSNekzdiR
eadiLSAVkG28nlWZsuyVEPAIBkHy3HCYDiBt69+jJQKEaHuUF53Q/R8XuYv9RNWD
ijDAjnZEudbUwN2Y06mehiVnnQxaUQRB3GoplOHpyPN3W4t/xv2xib/klZya+5V1
tRVNam1U79oIrKcAxgptx84zqnPeRo/vXjXPJzoNm6FS9jug4nFz0SGnKPnHICkt
jTNVvgJ6UYER6ad2cqIJBW5BwQMEJ+tWoETgubwwmrR9330XDDK4DRhgEgweyPz2
YCkdxWksZmHAa9Y7mBYYlHZcnVaT01m8MEH3d4U5r+rTLfzie9AD+jLh4mcPu2lQ
bkIwP1l/hCfayJhoM2cT4jt4yTXHX1bDnj90ecB3tPRK95kYFvOaXpinaURQchzo
6LOa+C9Su8WobHS+kUZldRUQMinJLyfdzj5ZSesstbJVzdNlMhFDb4ZwB2nu9/uI
XJDKIDUBUyOjoYuboV6dMnrI4ebGthPycE0jL11ajIV3yRFN1a8bhOKybklP0y03
Ygd23u2v4FZkCvhKv5OOrSwR6TUee83UKhEfEHH79tI+qExit0fK8kVUG3FuQkI2
xdFWSERfhId+zU4hUhRYpPMin1BC5BCnQ/BMgrP3emO/cHFcSSUQo3nLF7HvHgkY
tm4IVUBRZ9Vhc08rVKqzVtI2AQeD/NiEPRZhZ3pv5PwT7KC4M1+ZlUHR5dKRtOTb
djskK34tLv/PUv68hJsr+Pm24+uXuOGxLaaKPhrcQjz7Tzi1eereRrXDbusrTdGR
XeFA50D8JdbsE2+XKZzMljz3EH10krs2qVUAtZHY+G+ONrfNctQlql2bEorP0iwr
fyPP3Z47LMZgDGDVpvgtlWbhhbj1eG0kKYWvmjMu+LZnUBDjtddTKGm9TbLBax/B
KI0VqnQk+cHpB98oi4QFuE98HFin2DlGjwT/xX075wAEfX1sL0r8majbXIwVHuw4
BMHpY2fQKHe6E4zIc5OOG1gW4uvxhqau8VJsRhKzuSMY752lVixD7PMFbaYgC/wr
W/vF6gZQuuuYEyF92WVPRCSJqhDabxWUrk7hcQ0Dg6V5H0RcXOKryxM9tVnw4L93
9cJW9QTU6aIo1lBfz7aqcTFyvQ+vCCnncWUXnM7cmB0Tu83t6F8wH7ZOK2mbZ76y
5AFUq1O+is54EvCFvbvZevtL0BRPC1YPiQHmmPJveAX6Zy49kcIKsdIEuB932I2r
7OC4ClvRV64nARzbUNymD2xNab5OLty3cAdH2rG4lFm/xA1smoV6ThhvcRE6jrNj
ELgSLvB/O1XttyYonrGEkWw5JN/oEvT02Snc3WbGbKbO3zLa6iqJ4+ODudi8yCdl
8DwGvFrst23scpV4RkjsoJ5YTs0SNrz+RheZm0UxKtucc3p27SX3UC3FaDsOrOGs
U0kWuS3BVoCgwJwXck3yQW8zfKVihXG29N8hs4JKqW96Fh1hhhCMVl411JlS5E1l
kVuqgOcExFqADO8PojyaAuho8lug9dzWcELEg0qIZvHSVeyLCiE9ztX2VLt8Y+Yx
+LKGFEk11L3+PGb+I3ZXh1SBTyM3vHLPh76PDOXlMsyeLYoRL7QlLJlLD8Ab+0ZG
ubY/T5mZ5lweIgWu+8YWfRO8q5jpsDboUqGeahEhjHmS2uA1ku1+HHH/mIo8FEzq
UZlRBfHqCVwk0egzoRLLb9lVihjhhRiPMZqBBJIxFcXDBme4O30szvQ8+fmvAeOQ
LjLfnOoxUn7Bw6VXBgYZghFyDNYNIgsBSy06STMuj/kmsiPmom7ONLDHmMcsfgXq
XMc3Uv4IyYmwKy/wYDkoxdC9tQYFbkmtWva+ZvlCxRZmfOVEFQmC3P8nwxTkJ0MM
WHm0bFCZMEF7ETqAH7LM2gjtKjOih7K/jdgo/ueRK4Di7QI9Jm9RYYZ7ofOsbsOY
o08dfmRsXSrZW+mliLJSmZ8L7tNjPWxkRfdDAq1qZzP9r3FTetmTjDyXdFw8rF8r
2DOFwUqAFYkS39Uc4vPH5zrefaYyR010ko/FHmHbKkxUFwLlcpS9+Qbkcg0ljgta
jq+m4oHTyeQtUMyXhDT6QsKc7yWJjPTms12DF/vnHerSKltoZh6ysZT0qwjgj6KY
e9aThXt5pcalv6jlxr0K2DKu7rBBENUBFD2IOv4QfsP/5e5LTdBGifA9cGnP73lV
MiQPPt7DtU0T/uwY+NhcfbU5SPDaG+DD7fifAIKbGDCxRukphfIs2+rP4vtMhsdi
Al382+Zk/Kr/VDt81elRChXrGD5HWvzvm2o7Tf+DghIlJnI0Adz6ku6OdYwgdCJ8
mx+QCCvToYJQzIipqkqT+fJLawtHP6yvoPWKZSp54xgPNXLKODagdnNIIk8cVxtS
iQ5cCafFgDDLQBwa/XsRQmY2+Uo/5Wjxr/hneE3lZVriaQqst64Cm3tYpUR/L08A
Kn5HKdTcBmVB+EBYKQ9zSaTAM9HrS5Q03cf/vuz4k1X6siPNeqWBOYVcJjejTeNK
zjmv+s2QqxfIXUFofoVfZc11FEleScaFWQZp3tMHzpyef5kdmnkuivYL5pj1Jgc0
GV5KA9oIN7aJCw0ebbGoeClOn2p/zZZ8fX7mVywSGzfG8s4ZFndDmQxJg8FmdA74
a6btxUmWNgQnG9q+ms7Jsn5KijcEQL023/GZTvsY4QVAazn8HNKj/bIqWGg+cugA
LE/Sa5+xc7bM1yCUOjVnBpXjbqWxVOjVg6Jla2faQy6ZGEVo7qfLjEnKFY5dEBtl
gkq5QjwM3fDJkdZEmcfLLH9em4EJf4hgaRE7Z9z+lREXVjqCprOB3C50KzO7/GCk
201SbE/cQMRkoVhUB8TVJuPVxwv0m256QUZCCfrNXMEg4ebyxBJ4m2dXcVhA8mDJ
UlaoyzfbWNwpg2Lz62K3gxes8gcjwil7vi1aEcAKgZT72KWwLZjpxfvEepzKagwS
KGsSNj7mqOTto34tjRWlBLsjQUDyPwep2MemEOsV0FTRnXndWQUPyiZUZid6rssm
5TTj//x1ZfhPszNtQEaRjwJB7Zr2mHIoGXl4vYPA6M4GWUkY9DjrW+/BXxmeyMCS
FN2r12SPbQWSsck/Wr+8hx2fX1KQCitO0/lNznHc/vIcq1/RO3LW5CzZrQR617jP
buZ4gli87gxEURBXKkLQgQ6gcholPBA6wOg8XkrokJIElHBSSUkctz3RsxUwAgin
nL9m3s6guS8WPfAncuQdx1d6CUQzYOChnh3yNS2sb5wKG2auCS1WwlXc6sdmrKXC
n+RsSmEQsVr8rkNWyMuSP7xHUxAwqb862obJBhdKlXSNBYyP/zw1JQ81KKS2Wlt/
p1qDJHLcj1hO08e9IIfrI9uAhvtnh+LvfbQqSYYjcb/zdgzCteTZqkCR7q8Hikp6
kWGdI7hJrvEiwOr9UFelahtOWvTigOH5p7Qmt71u9RGmKyPBGLCrqUwnk9Glx0Cr
Zm/AL21AQUg1fw89/KsOzbBQ2ktqYBJqb8+xKea7Q8YlL8CS7ha2MVmKpIotlpMW
XZeSrJp+bFy9ftmlqhnwR74krJepN0wTUa4o8Zva2mw6VQbS9mzeg5Q3Kdu0WHg4
U5TlRbRy+NI5BFEEi+TSNIRCEri9mONIrfP5IlCKMNG0XBKNrBaXCBjdYCjFHFec
i5HbHIpSfpEGJQq8tvxFnDavZfkXLMbYAwfu1Uws1uUVhl+WQNN60cFvKs78SmJh
H5hqhEp+nZZl/ufTSaQvg5Q1Ww2z0tgTJH9O+rtWVFgVhpOJiBFbsZw3TmOWdZGS
n5+w+5blcKzMCR5NvQeYp8rVBHwdSBTY5B/CcpmaXAb4ZXXNllRyc9eKjH06vwdo
c50MKGsKxSuqiiaVTsRdt/VDxLRhZNU2Q6LMZZhuyDDfD8WyEsnslfkhJ+gL9qUz
5DObcHhdV7knq60oOvJzuBqqiH41OQUyu6F+gyf8ffWgteObzN96gGddht7E9oQb
gLNsd2U74aXyGFZF1CYhWrYhT4ZrJGBRH35BHcQphGJAjkUeSXjeB56/T2IdPrRv
A4ctyYHTr/30jSEG3F98cfaf0FL1/CibLef8V4VAA1iwLRxfE4mqZ/RiWeioOhGJ
IBUSGWOKbAZ1BSvNoSE0x0vnkmKeTZmHCfMV9kWPSb4XEHmkEIS0DzBnmd8jfZ/L
XzlJgIUg6+vpvwlyMn6R2jrK9MnIsb3bI1mrjUKWVKvHEavzfk+SV7RI9I2Q4Fya
qBTz1OCHnVIQprHoBIeBBWmoMwiotYn/Bi/tn1EMHymXEsJDcnLzsA222zBqeYra
OHUTGbMS6lTB9TwfCDYJQfvd7feuq7GRJ0HHpzcIY3xFdXRHp2XvUeenh+WZpXcE
QlgN/20hxqcEWE4c/mkNEWSGFtF6+NXc6Yf+tjeK+w5O8nd0EcsTtVGdEPoUuzya
NzwLuzkqcrd/7Cj2B6c4sFnakzYXtFxwc/nYniRmCgM4Vbt7AzAH3fvnVxQe8sdN
TXXYQiPAndmKtcQIkVgmH7nXyLQY0qPtpY5pSiHLkb2GAcTmI8Umg7Wt4HesxHh4
h3Emr2VQ6iKs/TfQuOaCYc6e8rtYpvNovAcR+vMmi4kdnZnPm/OzKbbV5ydGYjP6
7Pu7f1NBrMydFC2yxdfWIePdRHFoBZLDE2fNZsBkWpLs+fINvDqwuXG/NiavMpDe
blF/SxNaPqCriASmeppC8VU1RqH4tQMXWHxZwlM+BB5IXTA7JeqMlq7sUShU4+5L
wuVlYGZoCxyNiAEXRuw6L5ukUpUdeXZ7+reLZIUzs7rYAPYH67tlun10uSWZ1LOF
vc+ZLEc2NlKpxkubzY2LybA4aTg1QnRG2Fdup2p5pYszm++DSP4pvLcZ3VceKgBk
U1Fxz2wmBWmKVUrCHe+GKPewcrHfDc6wjKFl2VsW2IUCPDw/rzLywyIQYOi7jpu8
5I4Hh+YdJQBYxJ30dbtE6t6HZzcxcetWevQMkcpuMxa2eFYQyTMOdCQJngAWH+oO
z56Ds9LvuAUT4tYcokxfUsj1IyGJOqgw+6ytAcJsDjnx0uA3IRGv0eeAN/cm9P6l
VNoxrngzXFC5nQDWPY84pgPRs2yUGhxVJypVarRkpg1xht31xqK8E9sBzgb31Rcv
EJMjPUUvFCgpOx5X/mpmgGld3vS9k8HauLRQUme3ialvzirnuwNIxEl7Q+QkW5YE
ppiufdRW3B0VbagMSVCZrabvt1LbqIWgnDPhlaUvQE+hGPu0RgaQapZVCgiEVkQY
If6JD9Ij9TT9YUwCLdvPkk5F5uV40SJF9zuTuIdg9eDtnXFMH32cCTu/h9zTWzA7
RMhpLheDeH3uWLAzlv5cGxpoe0O9qgJCc6uCCZACgvcRobMcFI6WuXZL7cMa+uds
CqlVVzmLT2SLKDVigA5j81ZiHXGPRtSdZuPaveKFVqvlczU4Dj4JvNbMTZC3CRXW
oEYcVr6Glj6CURwMSHZWrKQ9grkK+Fu0PRSLT+ZVxsysOKBhQXuHocv+wqPBHMio
N6gMjwLeUbc86xKIuAb0NYvnAG4x2fvhrWJjVGYAfP1984i0G3uSOr78cDhQKf29
51FOXbh0uOugGs0izwrBiZDe3aQk6b3GRKWPL85CBVicJvZ7R+JolWgjv9/g6FUs
lRFRxTnDzkPdximYyPy+dMzsHVz5l+TRAgVR4yqwuF3XipHYR1hp3J/hjlAGzYQQ
uEeCYXQxGw+7xrXnEZI3bbGKM9wYUG4aY16rQjE43yvaD6aG0D8cA+RiXbKl1n+c
+m2vEyEwlPx6hRbi0Y877XOEq3qRXmtJYfsr+ns7vJPgs1FjkhjWbi3gRDcE3f6W
snrpvhp3bZekmnXc7f59/I93iorch4LO4cOw6MuVfkNvjBQcqr93NwLhz4QCcVir
U0p6QFMMOnAoJATAF3zENkgwKRY/Am3dKbnmisG9c/uTFdyesg7wzq5RMoGM+mqk
Avz38lFlXk3/VZoGP/71/+qQ8XQpNY7zZ0r/g+xrRYkmgtQUg7AQ+PAcfiYSb/PF
tHIoZeol5BhEwUmSlhqg+iBUOyX19G51xUp/PPU77tI3uUUA/tHFhSJYM05RfSL4
32N7ptEMxQIQUR/4zoUsT8mzZ+hXII+XmkXMHx6Wk7KQ9Uy47Y2hGh6NyR2gWT18
4oEKov0qejykb81c1pM6ZO42Ofhh0Gq9OgSg1Bdd8Ul0m0dBwnGtlGAu3rXSe+39
2YSp73T5oSO/vSZDV2fTM/Pe/1eCvPmxo06PBQ5BuK6jpO+Z4BFgNroePuiUGPBU
GC4XD9yNlWcWdLEOGxtFRC0ovtlSFO1QjvmNUoayouw=
>>>>>>> main
`protect end_protected