`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5408 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
jsJpSUcQTu7cBpkLybExAtJEIMHmXW7BEA+cLQU5rcFX0mDCHG04tueEyDbdt9Di
hRrb4cIi4VeFuA8K74AdPTk0oPmRdfclmgVB6r7PLvHqO84ssep89ooUv5EMA4pj
6GsOnHiIK1fvor9tw2atHoYnO2A57XD+tIZg4mbG4a5Btb6WYU7refO3SGnwIIQP
Ur+VwPrrE6HqJ6enCW5K2P7SRZFVBSDzTUeKkomyGzU+0iPqRkUF3ye9+PgXK/oi
1gGbkVUq8+v6o0piBIU1e8+BNRWArovvqQmbz/FWtnMJOjqdnh7d0ltqZpDp7aoP
wOh4Hu5JHubPWnHdBYWzMPC5ads+cOqIK7rF54rjkis5f1q1MfxZn3O+4SPiZUc6
KCftNjevgeOHTHVSaApQJt3nEDtuK0KiHY7/JsuOOE73T9yDe78eSd8z0PeoS9Sz
2zvvc8o0HVrWGC8psGYCZqYQU/BYAhcwRKv/mgjIbp72U/y9E9faCOcsglSqtWQF
TDQ61/bghEGb8ly4TkK5h7sNX8RJmZ7pkxa/RWdYwZEZt42aDnRDTJfI2WiPkSnQ
0NtfJ2urY58/Lf0RftPtv+g4iBPTx9Hrx34k0nrvA/3fjcELl67uXqbCbJE/6D4d
QCxiLOE7o9cwRywgHB+s65fA+d/6HpZLRjQczSyPftm/hobgMLvHQ0YG7Pm8qRog
/wL9KSq3zfp+p+zMd5+iUV8Fpf35kwOCcZpDPd9FJQmJmL62TlIX1sh3fv3DQXCM
2vtXpgqX2j3iKX++4/SoA+67PAeKh1VjaoGaegKFGBBOHrWkBi86i1wxfGOjWIHp
KPu034g6QSUythuNOg5P8q/rlNohIgq8CS+F5VN+Bm1cJUCU5w2ParKsr85SrBVe
yI4Bwrp0dLW6MZ6Va7q2sU6e3e1N7kl8PJ18yrHicefh2SQJFgXDFNknF4dIT+PT
AHB9EfVN7CBpS10xtCgJxYViudFDiBIOvbdQeaAFE8djfhdmLGRlNomhZYseMSYP
3YIVsEeDsAYUpJ2TOXyQ17YfE2w3Gz/S1aXQsunbOVPeUpfUfS0P7t4LeDoZHOBh
d4Qrf/BE9Yu8MZ5NnwgXvdsUzzCiAf1YwmQWQG0PQwjBVpMI9sRuQg0g/VzZ2fNt
u+5Nr+PX9O/Py+TNIxyMNDUcA+atjQc54FTHNUmeTTF/1YVE22vqlHAOlPHVd8Ys
JeoCygUDxeU6S5GxaixnYNwl8ek3nJh3v7zAikgsI8LPQ8CIJ8RslTdKCQxlTogv
9c0NEwIhPZlJRYwkRAD3Oj4cdp9N62KSJDWoW+JAXXqwZ7vonw9BPA+yurvfW6Sr
kUVPxl3/vQMQK38pzz9hgFMOqY4dJquDVb2HjTlLglWkxlWpcYF4mdiHykuacED/
ivFDslIcP6tHGpti2XCLIIDZO3d7VFt47mEUoCzHrUDGAjgAX4z4Fx6i5Iid082C
hjzDv23Hg+tFS1uCaWPTyZg7zsOgMu8Eynur2ISp7LrcpZrqjINWY++4k5oOXOx+
ByHrDuW8m1db/lq+/6MAJ6Mjp2ARicMDqD3n6Izbx9rBZriLfN9sO0baQJlfSOeP
4fKEtRoAOCekhyAMifZO7VoMIGMLPaVQfxd68Yd0ZpRtqB8UKGMeFnOoD1ab8Nwv
3WvJrlriuqvHmzmb2Rc4mXwzceddg1b4/NqKTHhvfKV8uMh/3u0pB75lPPPzxi56
b86IZpKG3MqqAxbTSJYqPI34tD8sj041XkvQu9/74PKOaJkCRcv+iDSV/06J7WSw
XxQJSYzLqnh4KmSP4U6em/b8Ri7a7BkCWfQ00xeTa7+S9o65bWEywRu1aYmRCJ43
KVSuhhvUKVap7wHxFkDuT9qqAHuVZ03UXv76Ax0MKOF7o7bvQTzTcagwedY5pVaO
C3TkohE9lcsWX9+eGOJq4LfTp7FMUXGgxUD7V3vty4pwxB2iRRMDJj4pLno84iBs
8FYpKBI1pZNARd3MXaDxrTUME79W9qSiggTkW+HX8cPRW230ZN0wHX1rj8P/Z6WX
1zFgAt6Wj26lL8FvUTf46DWCCvGSotqvyTmtv+mE/NkfZ+iC50ED62mEKF1ci67l
S1X8z7BlChNb/HuGjxe6CLJMIoDNHt2EzGf2r3MIg+kReT/ThX0sekzxzkNg044U
FQV3kn5a8xcXFxUIjFiZCJaZYkdIDBvvy4V83vzRFLovz6blp+W9G2iS3TCtlFWW
ENmeebq31Gl6bOHorGXfbQgCOuAMpm4Pi2VF8rUzwm8qSHyKtsu15vopCUw4pwat
xKH0xF1AZQetAVIUQAQvz+2trQKXLdoq8mvGi+gsfvUcptkXwf4trsAdSN9+qFrV
nBbtlGzhKpevDj+JdEP3bZrhU/mVasoVDCIcmIlto7E/lW35ln++ueZT1W8CM0KI
ipJZT6PWQv0clTO/S6nKWcsvl6qxqdLXspHUhQ5fOKXmFHBE2LsutmjGU7MuVv5h
/EhnMi2yt1KqhVmDQC4b+MyWV9JBeQCSeZ5Y5D8gsS0xpAAGzsr2YdbI1RbM2voh
kG2z20ALtzvWdaFF6fAuQl8z3ps/hcjFFMcMvSxuY6GGQ2M1iykAP4Uspm7ud+Z6
pQ6HuFRPuTEEeroPHKT+/RFxKyr+BQVb/8wOeE6c6c2W2UeBooeaM4NXHmtApsUi
CdHVf9ARY9kyYOQSnCMOZQ9EKXYW2Cd0382NypxGD8kDnToBC3If5eoFXr4DIxxQ
bHW8F4F7dHTfCVOd/Z6SLxvasJAxM093AmXxiUkkpiiVmVq7rJE2HufZcKhjTZWu
mdpf2e3jt8EdpfdHNttXAmwbMwFwq4VUTrVmGA2ha6KOkf5eURqXLRAycj9lktan
lVuSU08xP5d5F+ZItgjKgzPSaZUZ5B15wngcEdgHC0bH/bZY/ftPD49TEtilQY9b
k/ShH5Dsa2vma14dNKuSPWob2m6qDQllagP4Kt2aTf7zFfugF/S7/Ka6gfg1Kt/7
y3oSHNtXsF2xFBO35//vwiIwLeZXANppnZH3ElCi7EKesyjXzm1GFMcmVrwC+QUk
nclA+iQGfEZZ4hs8AX9IZRI06RwzbWRrneQCK1/N2yy6Pd3MJ5Uas44a9rc2Rg08
2pTd167Nn3rhRa8YBa9czWy8XCwHHTfGm9axDif4js1YYHBQ2qXy+GZ38sQI92Er
MM+iH0xLZcSiXVtIg/vPN8iWvKTL+cIxXBtM57eLOtJ54u+zHK7G1349g6mzGjsp
DuLTyvox5/iWQRiN2QcdStLezg7yZizuKJlvNuOCHxBsHomPcSEKxoicxVetgXBt
1MISawNq/EklEDdimxuzebcoVquSufB23MggOtJN2CFrIEi0Xq0rWFVvQWZlrCv5
zluipQJX6cROvkX7yzMlDD0/5ZgW3EffXbGWDJHH4kx2QgiFR8TwS1PasIha3bmF
314DlFyX4sUH9sprv9pgELHdao1zXKVZVeK2HCkZZHmOpHW9FwCTUjyelwwjFXvo
x9Y1y8qIy0kLCXdd8j+mX4bgBovByK8OZWgIhcOfUKo5kJWDISAmUF+ynRvFilhM
m7+7ICHFOV6VLoj73SqlpBpaxQPlKMeMkofK/qEpJcmCIf9iDdfUmpnVyuLFHdti
RnMqF3nz75hrLkn8OfaDZF2hUhOK+LTVZZX7mUd0MNLiGYqGE4wAw/VDVW3cbXGP
n4Xc/jo48aDSAsy7Ih1HsMqOYpjx0cVwDU/mNxFnITcGtajGINrgRaSP7/gQtwiA
duXIadUHnkgVvPm31XkP3hTUdvVqee0UIiX1VqxC75+RxroU5b7j6j0t8rJc+XFs
F+LhBlmBmqD2zN9A7Llsxuj9DS+6Jb2dpa3AgqdVh9AAcnazGfYrqGE/QT/MJ2zX
y6QJxX3fqybL5o2z7zKgPEE0DrQ/zexjTHi1/NIyBDjvwE+EJFNSYK/gfl99L9aK
IUFDVuhKfTYPo2T6m+HdNNQJCWFNTxp+pT/o1S6fnctFL3Jlw+NELZxsq4gjFZ1d
DWvoUzJJBBAl8cdy02HHTA5Igu1an4Qvg4tGQafdNINQY/d2fb84KawRZM3SPgdZ
B0MJ5dEsXRTqbbGQsfmoTiR3eOabBCFt+6npJ7btha/OeXU4u+SA2sjAlxpuIZ1T
za6dhfjkEY9ryrneS7HmvRxamFq2g7/YRWddF0voBzResA4ff7J7TYYHFCPf/nQr
Rd5uVNB8rJr1pMyb0IOIpKJhxRcR7ERwMha8FePXirtFI6RdCfyWdd4COUJfpk3B
7m9eZX8Fug4KI0U/QdxJ20FVw/tZRJGVFNABzAWe8iPtPsUFCgqY3q1TiRDDzOjz
uPNT+VJGxqm/m+YRQV5zoclhPbsrZgQNwIZBFa9H5Ir92jFn67U+RThEYvzFqBRM
pRSzCCTbQ8XQLzYGQpto2KCxT2u+pNmgnbSiZFHjWHIEabsAN7j9wp5MbXNjxTFc
8oPv13HXlei06qFw4/ptzJO7YvlO9G1J3G6ggqW61vy1X68lzDiv7032ZXipZwMz
/Fg1HOP2+96d9eAR++8FvoyfFH7419qjqtCrli23RVyG/m+rjWm9aQEkgmjKYNQs
2UE7tnc0ZOEm6lpd25TsNe8QPJhZB7TMCJsmnUsYbKz8oMyJOC416auWulMc4EzM
vF+9L9gyYC6WcDBPGAR1HZCa2TNkzSSt0c+kekIgI5tOKOMyBsoYTSX3Q0q6jMAk
Dedt4sCcqgUICIqPMuWsrtBUwVyNhIfKl2iRQJftggFn6ilDXNun+pObFkrB2CZ9
UehIYvcey8K9HeDk2E9+zb+qc2ngtXix8arVrpuhT0CG9SiHzFfW3/y3RjxZulsT
TRGBaHvqGwiXJQYWcTUXHzmSrUU94nulUFhPPlw/SCHmQZnhp19/S/qW9K3g6pbl
bsqeDH93lhxacJIESuFqZy2gOzfY7xshvS6M/o2xRhilCUzpgAVWJql7GSt7wO0a
Aon5Ic6IbKyzKnd87u2CB7eLfGGvXjKOWuMxak/Lb6ZEKp1WIf7Hn2MfKINZoyfA
NYNYC0yo0MC2+lxPAenKog19ECD+U934Sw5yIcKHzjdQxsiawmn/KgwiwnnoA277
UqA2Oq88PVfdQDdwB7xf3hg4Zf9k/AavUzrLnpQE+6Zl6ARoKtqQVyENKIrSjrBj
Nt8f+5PsI0ySJyWC7h9a+qT/xOrVhs/qhf3zazqu4l/EY6TA+KmATCw6ap3kPm+D
idRSMk8LlJBDUVqE3yiqBd6Puyap9iJTqjMp+57mT17oDaFlq7Mtambvud2wirbM
gRoIfgbqCYQtf3OE81o7DIxb2aJ/4Qj6iOldW57mqW7oj4SYTR/2oNqfxJ5aVLqb
ij6YsYviqSfJxrwVNE3CTgBJzQId6fXJar/OIr+YaEX+6c2y5l9MMTx9gbMm5BPO
9lDDN1LjqyiY/LO/La9Lz7Phv5V6Bvl8jE5udfmOnFbxwOS+BCepiNnYuBNUw0cK
Th5JSxPradsG9TlXZqRnhUDJ+dJcoxItDI08GZrvWIk9pE7yhvQ3TiM63m1DsebO
5IIxgrm7JL9glLAy/UvMgN9/lbGnXT/YBio0iSyMF6IRRC8Vyg6bZ34EMK4XZdOG
OTfTK9VpPjT4itkT7s3VhlqL+ISYYjQf+d/UaKDIgfCEFQEz1lsBbfkptYd/pBSA
mrnqNIKCfErrkdnsE6zLUle1qgCI5XkOPfB6Cr0v6eU6Mjk4wQFSL/OjJD1JkARy
wvUV6hK8pcnoF8hs7XOcLw72XRwNFsU1eKC/396filc4b4S7mepHr+/RvfCtJhVV
BDruR6I7UxHk91SkRHpLUIe7gy4jR3C89dRzIwxM3M5xwXoQDn1EzNa7+B7TPFnJ
pmK/u0597iCzqa4ow0ddfWszFu6erNHCm/yQmq9NdWGnVZuxxnNRsbp7PNxIqTdn
b5/QhxOS6qyikALDE7DKpJ/kEpL39yyweuuWES9w0DIywkjr9RsS9ibAC+Wft4Lf
IHgMScE9dcw9ZSJaESeFXWTO1X7TvqSa8Y4Ywx2RDQ/nqhqKRPkwEEX8UxZT1OGF
3Us8e7F/NkizlAFAH4Jlxdkhl61zjuPKa/sD+tX2/Amx0k1HRlFIoLmR1GsOjUMz
+rOpiZVa3JOGigSwWeIjgoLMukpJ+I8oS5UKxB8pI2SKY8Ix34Ob0M5W2k+Vk6zx
jIYIfXnlkTZJpZIxUBcWVZbWgFWFYpgTn9kHM7gh/g4m+jqFrPmsUdYjV1z9+7ex
aAST0zz++hzU3v4iznm59AxNh+YJDkTxa/9l/Rt/n+JX3Mi347oJZInwUIBoOLkN
kO68SgUpNX/77xQMVbmcDttNP7Ba9kh8+RNuiyt3u8gLmrIWp7flyH47UKN4wJIe
bdlUkr/PL2dhMgK6nqGQoInwTaZ7xCmvUzFl2N9O6MGAQUZmbgLIukHT+XBqdVlh
OT75iBFlBu/z581qRbK0IG7SrCQzlGvtimemJV5wTXCf/S+cpexJwoW59RpPcLy+
Qa4o4VcoEuGWHL556jf9JfHqfcEv0A3eDB8xWWCQKxRcuPbeHFZ3irHeBbS4wAs4
KpkEA5SQXhjSAQfNaAW0OiWgaJyG4T4wXU1RYF3Ry2+yzb6joubBqNErHTySCvB1
kGl7POYlPUGO/zEr2Q5IFcvkG2YTs1TcZynEJFn6dl4HVF1Yn2zI9pzy1QNj3muk
JzwneWBXLzq1svAQFD8GfnPbCGDzrdDplpHeKMOWo57JFgrEOwoZYfy57uIacV+r
IV4Kn1AuaSdiDURyCHIdSH4EQnlqRbAZ/K1JPP5VMmliUvj/fMoKiXAnAafnBgWU
O7Ja6h86HTl5kC0KDjDFWzp6wVG28r13MtKrtxokltCsMFXj18LJZ+vYA2sYk0f8
TkTNTWHgKX5Mz2QlSl8L1jk/EjjzqW8yzIxPdz3ad2sTK6dzNqyqn9CEGLnjCl2j
FizoFOv28xzFkFDNKR8+J4mJ9/u5gHI8i2ZFH+7wVzSzz3+uOf3G2yb1qV7JnX+t
iY9WEB99e8Q4o0fLceYnxMtW/9CNwusSoEf8um4IVBA=
`protect end_protected