`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5744 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
/vEkqJfyK/81z5lf9X8oFbGaSsKBcqQlFpb6lXHjj8ppPCJE86oRKU7TMNQDujgy
8bEm5MNfXj+fb2jBTIBwdw+roqbOMwb3aJ/hrhwHdGZt5aFXEhIcV9jaPTJh9xCP
Nf02RY+t02OUJuqWK/QEbXXt47TABpyWNzzioOAwWrcx1fDr5iUvO/IllzcDvG7k
dHOnQR6PpAT5FuTKpGF7DEiLcGz52o0mgfI6UlTdsvkZFzVbmJD1O5DbRd3+fJWZ
IbAbA88KCLebuGzZxvmC1rBnSrYrZzuNya1jiJdrQGOD6erI8NCxnXN+1oDcgQVh
owC/+L3nYf0HOGQp6B9bsjhEShNJ6UUigGQvjyZnPgiiWlsuxryL0TlIiWRc5oAn
AXR4JAI/Yt626b1LBY6z4hMjDiNv69CDFHthpdvOBTVRMwLAY3J7wJIoeNDNU3X4
nc6CJ8BbvXMlaSz90QSzuJFYAqyc9oLsvVQxn8UwHRnkTlyPXjevRUJ+tO+rsGo8
SiOQbDqw7QBRz/FxHFwP8rf1qW/czHau+QMpxgBYJlGnMTky7W/TjIIkArbfooH+
4DtrzhpxjXu+iqvAHKlzE4v+5ZmZSaoubeVtP/C5x/mRtOCm7vFDORbl42LQGpmZ
+8pCmWKyISEJzMHvUqsUDJ778gSuajh3WNH2t8miQIV508BTyHq25UJjhG5QgXJ9
58pb1/IeFoa1RQWhQFZT1DywXBuml0llWc/Od8mifV/P0ZKsY65WAmHk9+h1jwfU
lIj4zM/hcg2c+/Qp03B9prDVeVg5/IChewQxQrTZiGkWkHFvHi7wxENqa0ePaZvB
13x8MaTwCHwjeyPXaUAfL8pMcqFkxZtCr6Q7dh3ZwNxU3U3/AZxA5tJCo6f8m91b
kDTyzUK8SnPvO8Y+oUSQc0kuvDqKOHWEYrpLsKJF2JNVjf5hpqywfLQa+Bcj/rZu
pXzrahmcPMB1gu8tpm+Bsz8URVqQBuQQLn5Zr7tkz7yM/ZpevxKQmShoT06qMpig
pZs2Tri8UfHlb2hV9ekSS/PUEEcmLNc7bl1q1w/4eI+I7FH93YvH+mwDox3UcyVT
fSW6T8o/MnS2cdwsRjrXN64Fnn4bqJ3RdTjVziuUPK5y80aPEDZ3DRkbpVml2Raz
Vh3uQvgEEeJOlabsd0pknUej9wZ9c4xzUNps8o5VzNThsn78QhEO836PVLYNQKtr
8NRohap8ZUL29BzVKBPDbNR7+9QJjUonDEV0ZAAHoATFijp5MHk1cTsZKDbcldj4
9PF8AW+wSnj+U1DKy66+LqG2VjRGd4GORJrn7Gg4xhuaDiwjZ0vRZAJ1eCyjl7Ze
ZDwTbEokeDJakBQG2IOSm6Ut24Gb7C+XbRkl1+5UNACUDvzBaORvklFrypQEaJAq
an+KwojDyt64ei8+KYkxkJGDEcZAFSPzb1j4RggFTJdIqKofXfq2W4Okoy42wn1W
hVd+l3bQH9EBk0MK0wPOu/QWDpb/BIfrZS3ciYPpnXLYhK+sQ40jBky8Gq/lDjkc
4ONzvhweVoUsPAt18p0ZcUbs7h9H55iWGKl1LeUA8xNOsfi74IM2wD0nb5SMThRq
8Zs2miHxrQNbMWWfyQnqIyhXO0es6tlgGpp2UdJ2bMfQZr0eZBm3KDiTv4VglX5T
Snqu8mx6XhiILbk+TZfI/jm0e4SKpjp7cDK0XSnIpH88T8BIvYjQz0RTCPl1sQCi
zznjBbceN/RT0icHga0t4QxHNGAEyIQRSzTSO960JqhhlhZmhkXavcyhIWNzwT4s
1rjvfVOIQX6R6aJvFIS4LPioc/EaBgsFsh2A7hy/7xkxjHICwqvujM6N0bEb3oc5
mtCTbk9NPCejhZFrDtpunBiKK8LPUK7a1VhoZzS/C2cIfHfA9HoD8+/DN7fxP1D4
DxIwogAB7hzxt4C7Oma4Yn8MNL+n5umkpukdfuiZl/SKh7qHdYK/3akczIDQvzwS
V/c905Fnuyy8ypbvv83Iim4XeSzRlBYG4OUpCAee15R9SQS0txsKFdkZDNNar201
VDWit6U+xTGKdGtbTiHHVAxZpdPtXt4MUcju1JTgNxLvReoMvdFTtnpU0iyZwuyh
xVr72wMxaGS2NcSaL2x0tjPyoKGDS26k3PKkNi54PrPu2V00gcVSOW5KloNO0Iv9
5t/dm0mtT3MBggWXipzELTbUsyoGE5tixw/uBwEHz8JrtFxLAX8XtZjf3WTEqNjW
Jrs15L97pen/2A0xPurpWTWrqU+S8OajFX3llQjNrFd+GXZIGozUhAEr+y3jdnDF
svkqcIBaMmh/mxLf9p6gzzVLz3YiM9eVBn2M9s0zf1pN5ROmUAwQtGqqhtj0I5Xh
4mpGdVJndKdGO9t5Z636bF9W5y1O7KZQYgcKGe320/WFn7sDZBrfRvgUP2EzSOsD
Lxwpm5k2P4pZEnmyb7/2NjarJqLg0C4X81HcRNVIiJX2PUx+JanFJK0y+FrqWAgR
grdbsdXsFvOCrr3TNEyWty0Wt0DOVBmnS+O8BfOyFxhQDRDXck8J4eYy8bYEAxlk
FtZ0WfXX1grRGtRcRqEkMRfv0JTVRZctRpaPlmiAlva6lAXrMWorQ2PwZGT+a6+Y
7AnFw6k2PvYiBxv5xQY7pg27vornvtj4sVeKu5WmjM+BxF6/9+VB8iRhGc9RFzi0
ZRioxSm+Su/XzaNQVIf93oRhmphkrHVJANlf1bAFxrzNuJrtYFCRDH/JNq0mlz3v
S0nrCs+0k4GM7yca/t1TcOOOgT9KEoBqVjpn6D7763PaZR3vaZPdHlwONcEUCv9S
8YcQH6ZZqJ7Oixch0zqExJ++tCDCR6RpjAm3VaC10OxnlQgmkNvtHDoXYTy1QqNM
17OoM0gMv/uJFUJtBze1+iHDeLE4BFVL1meQOA25gcNXDLMgHXGlRl6Uih8AgDZX
i0zG+ZICaa3vAJ9D3EXJ33PoQNA2WxBAqmlSbO/kNE2xPVVOJ4loXb5J1Cp6rElE
WsMyJZrO9QMlyBwY8NvKQZfi8nNe19CqQStR1wCDxg+Jj12bWtQcBy143o5p5818
qhvVbmlkodYT6WJ/zZjlajNn1OhXvrS5LDWdbvPxYTjzUyVnkrqTpVD47ennFaxZ
T29Bhee4UuIzPOKPvGUddraqHFFd2h4GOyu/Ty46tfULCJNmJJEcmGIOb6nm+/TD
x4XzG8RjTKcxzBuNv0aPxFsWUvdm8OTEF6qzOZ8/EQfQjmaE8nXgIk0Vr6GEP1p2
/rHyinxlh3VrpjxfMHx7xBjorz4nE/lhmlSTOkft6y1mlc14OvRzWOdHnJTMCCKD
nVf7tizBCyMIwrxV2VisDxhdUhJQw2qgeDjNarfXhzu3brDuzXgc3YT99f9LW6q8
dgfqoKYUrF10csPp3Xw5ELRmR2aaXvhxkoKMgWOLE9Q0DwhEfPGnncTs3kLGczrE
+6pr9FnZ346Z6qYdV6hO0EGsVqQNuG5rO9rdM8INiWVnNnT9MnGG/Ge7gNPF/HAs
+qn/Hj4jQryERJMWjXPg7pkulFgkaonGmQQyhamy9WasOuhDXRdm+nHtYviu2aQB
YksIcXZrnnCWAw4kbRVFIIgy+teFnTAULju+YTyUlmUeomlIlyjFJGuMLtn5s05Z
kUEpcrWARu7CmcLtJo9oTRZZjST0McTxe13GUK6qwmLHhgoYegZywjoFR56X+eQ1
xT/X2DqepX+DqlHwiAubpNc0GWBJGqM5l891+DoEju15INtZyLxawmFSA+f8hFoI
4ZoyIu/19Io+jTl2f7fo+zWi2kmlutrM+YeJpgTPYzY6DOMrlU/4M3Amlc8/YgMZ
NUlRkobdGTgx1o3XHYOUAN2HcEh2vrTZ0rpaKydOEvgYZtoDUyNIdYNISLHY9/S8
aLlmmyVPnRJb0KDPIpNAoe2CNovgRsVHnUb/spoM6Cz5Ue75r+fg6W/crbnMPqxN
cN7UaYa3d80Tm4ZulARnLg83srMZ6ONtqDGwftpmF8feZ1J3c4YbxegAjMM/XxmF
mFR55Z8vCvOM5vNmSddVB03UW1vVUQwHAXlHIjNZDIaBdA3lGiqIcVHm3QtNNQYo
/dJydKqk2xT8QbQ+//n20MJDoUkpwQpRFf7fLFTJNxwdgE8trAMJXG8KNYPPyXxh
w7hNyknb6cQrAIxobo/9wkfg9p+OCuPkz1yR85j7uyZUmZgk9f0MetVMTzACjqVG
D6bJHXTkmtKSu2Ho1CGZNhFla5E6h/zYlHwPXBb4QV724SlQ+ctTh6PS2LULKzcY
kKgGvXm7dioDCz7smqUiS0RdJgFjXEGPoJdAW3hwjBS9Q4Vm0Qx99/EbYgkAVJIl
DiwgZ2EhgC71w4a7AdUQVgBGztK7pJQbgzfNq6/2QNt817fjE8fdoM9Vwq+dXYa5
W2p9bl/dzGhcwUXxdd+5Nx6j4Bpi+xuLymVmpRM3Kovt/snnGrBqDHD3keERNrAY
uKcBKw+2t1rXmUlhxOJ5/60M8/1bZMDqOEvo0u5b7udveB+LKK5vYBEbJad5r0LX
GHeg5EuHsR5ZM65x6G00B9W9nEQY5tWsu0JSk+lWhDpioXg9qIfny3WzVAwywLAP
iH6/2hEW6YTp3m2MZtYBTlgDH9/0LocVuhttkY9XITwY0XcfziPNVPiD/vhFJR3t
F8bo5oiGBP69Zo7pHG0nAvrIKlyNXbL85X4bshIkpI7UImEdTcqCiClo45Zr8XsB
xuu8tScjZipex5CGRJjO0LPhuU7YOFZfxIZCkJdbQ23zY7HPrtmdwrZwEyICX17F
aRisD8wfZ6lS7m/Oibez+ew6YmQR+8Q3LZHej8qjGzzpZsBVxIn2ODmg23aKy8nh
6dGeQhMj/Xijsg+QEVehjLnJ2phLCdXdezuA6IA8r54xRqiy4/gHRgqU3Kwhc5H8
Nj2fEFGWsxl1evnbIasEN/ycC7D/GneMT5vBb5hQVCw9M59+VndCeeb8/DnDQFKG
qos5RSiNSRPP4qYUzUnS/0IdUANErAIRRh2wT2TOlzliD3DXYu9xpHXl59qkdu7O
/sXZyL+qpLHxM+nMq1+XJI1mMdgA2ZGmUeJ/0SQebz0u37UCkjt1ttzz5rAOr+u5
mi5bkkCUKPvS644tEGNPF4ulePsGq7WVBKK35j0Y8jFMYSlUE4yiiVV1Nn3xtPw+
Iu1JgD1amG41RmkmH4vlfwjmgo2X3IEmggbdexYLjfbIhEHSN92AQczdvDicxXvf
pG5KyPMmQExyWMSjtvnoTfk9rP1LLOZmjeiMbnsMGg1WSIQhrW6IJW1IM4xs+lwI
WegwO9WbVEPyhDWu+lzzhfy8VrIh5qxrovQR/z2jpC23ZNKeaC6sptW3WA4EIMR7
MvtZDprzXUy7hqF0Dlq9/wwc3ZhZD/99j0KNfGOKNWsAyJOUqy64jDyRUuzhYOkW
FnxYmpA/teJMX63191obtSoNCHq1q0Po6z32wsP2vfCHMCcJ3Qki9POnic2nF8F1
Peb2VRAONW0vLFrMZ1SyCZqTj1dgwDhMzyeIAkyIZ1fotFh6o6g5eWqWXoIprIWj
5NA3/YNlVCCfn4uDsS80F0RL9fdUKo9ychGY1K6EIDeV8rP9Yetq2/Yshp+WqNXk
YAU4AjAOKNTRZVqQHAEw3AjKZ700wzNytlXYyvpESl5HIA8d0pn6f/+V4OaXysDw
B0MaTdQaT1iIUdlQmyyEFd4IuYJqEULRbt9Tz0r4BxThKz5Emdmk/UjKid7e5EfA
n764kSv86ikh3i/6lZx5QeIl9f08P24HqrNwewrD+Axi7rl+dPyL5HejCIUMhDDv
I//RNDetdghcAKoCovg3MYLKYe5bPEZBhGE4uy/kR+CzFxM/+D/ob8JYEteX3vmc
w4J+9Aj/2+krVCKcG2MmmXjwmzZ6un8DGV7/Pjis261qbHCR2JYCUp3fhod+FpgB
QftTrL2rb25nMt8/jyMj8uNrZICFNK1CwdD3z6bzp9NTyJjT9JocmhQlMWfjRSQt
aqouPX1OzbMRfBvmvWCwXLUihBALkEXNzl7+H15T+2pGicpmNolBShMDYwbcREgs
gmhAV5jjBd+Kgnnh07M6cknJ2BDbwGHQsPhgehT7uFiELIxYqo4KsXdomO7Fn/eo
QnkfwYtMdOZrNNWCSxSfVAx/P3V4LMjS0vE243teOKF3jJ2/B1xoGty+cOBsYxx6
sCEJiQRpQRZWOHMyc0Z13VK/ZvXvE+4K6MIKJMMgvcOcHwnB32Do/Mdy8E1ZMCIX
GzlPZevve1HlxhY6F/YGGL7etPExt3jPXjLnLdjShBhftvnWeKErUIMS+fkS/SH3
iz1Aihl/9RSxLT4dPKE6E15nzpBghO5KwjvkBSC7oAOt8YAej7gEIXCpxPWE0e0q
u9h3UlEkOO/2skqBRO8rXK3nJqEoCPJvpHVUOQjE5lO4UgRwWFSd2oPXlYcn3oh4
hBPvz4ZicT9MiZ0gS83sZSxNIi1Zqo2WQfRBnQ/1dOBtmpoKLPLZ0CdyRn3/u0nv
+qvoN5RoM7xVvten6NFS982zAmB2cep7Nh8PE0kf04MPVkHE2hXzls3EX3jnAHM/
Yhk44p7L0IC0Bp6mNv+6Qb6rNO0M7pnyhUzK9Q6g0aWKQ7hbUhA+afPqKNuWJTUe
SlWmDyyC9f4msgVd7s9Cfx/BxCkVwmCRIiO9++DiUuL+PQ83Ob1+gwvmk4nB6lLo
4Piez6tYFofb781askh5j6kIbIo9mmxBkbaaCrKv+S/LyWVzSLQPFw9jVwg2ZX5i
7vdfidGXSrSe14hI7rbNr7mshBOctbc7pP/2St/bziDIHOjs+YHSxssbWZa8rho7
v/zWfGHerT48otKaEoWSbMY42AsZhEHtoXFDNwC6rnHoyUWE7Fbq/3GHgCWc1vHz
ovssOa2MpTksWnC4gxlbVBeC1cFRtaz3ozf21crT/+F2SjE5WIDvP51AJdJBqkzH
Y7fl1htpzUHiPiHZFGDFOj3MnVAexxbuMvtEOMNWdSNEvB4QrALPYWasowNsk+St
hk4kx0fOUHEfgSloZHA9nbG1Lyw91MtdIOMSN4I3IzDijI3uIamQ3ajWOz+46gFt
dX+LT6SJzESeKqIXM/uT6rNZFJzsv71JyB0GsiE9Ni04CGim9ZBTZ4aLgf0akbhA
bBMouFrJMblXdAwpA2OMZAi6XTadOghsQMHo1NtpDgcs/VnwUhFhpvliiXYOZv8u
bYK5fvQCO+i7Zj3KsMaC8EFQEAUig/2o3Zi76KBZA3xwnD/x/R53YxNXnDDR7k3I
t9oACzkcjd3gcbzREGNq16B3U3YVjGun/5m4tkl5a3hkK50Jy68U802r0cVGS+HQ
uE9U3qQW2Hsn/U6b5++gJsPDjH1RKg/g16rJIUei64EJpr/C/o/dHYbqEYe6SHcj
3VqnHmCw6uPAF6YoYmw/uIDIGgoG748ydI8utk5GfJ7vJdY70o5suJXn4rVc+eUp
DZAQVHozxr07i++UyrGBOqLS30ULUvqW8PsKO0kBePY=
`protect end_protected