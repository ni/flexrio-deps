`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10080 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0gkD44Df5ZOq7aSVZjrWjnJ
/WXLKlHeZqe6U6WSOPkhl2d/np1YmjmePz9xy+xt71sag5Oy2k3vJKq+JYzWDb5m
QlrOE9BJuezC9xSDnOjjkFdC4kFtyTfmYcCvQDHZ2rC0/uBJskULCCgCAQtw9mf4
JZR5M7LpVDywGD3JNsupF1UvfBGoIboohx1Cp8qpKlacUH7/MX7uzevow96rlkfS
ElyHnoQ/1NwLgtcBuj+yqbOkRF1Yk3HXnvbeZXiDNvmuldWxsTmLTTfsAoOHK457
S+mZrs1xVMYJwaVp/JtMi+znuH9/cxvsIP+hJMLNRoEXZATTbGFayX96TNRPOpCW
2mAx033rn1QfA8/aM59z72hN/RyicQXvbOVMrh0FvzZowXl/4YnFlJNIaWygNnK6
YP9i93BffCyu28PvK4zvmRq3pJSxLi5v4SewafuxJWUiV1Vr3hCKb2C3H5b8aCd0
rz2Nx3SwomWohOZKxV09qGKqPBrxRtcdP5/vXPiKH6J0/oLtWE9XJmVgDr6pf2qA
/NZfS2G19M6wDm4p2P20tF82ZjRElW/pJM7nIDWI0Hn0JTy8nPy+ECaFfuAW5cLD
VFZBkmphy6tSTkwLx8GkcxZ5/6KYdN5vt2QCHTU/Do+zkk51+UMzlDHBhbE7chLG
Zl1MwmjqhEJAnUdEjbvIXcvfcSlZVwO7Mmc+apuwoXGvDCpwZEE+4CmQlG++c9Ir
3HkXbydcNRn9eFzxQEkAq18jcHSRX45WZ+tA4HNqkshdeDQHucZTkYnB6wbvt1ny
Gfnr5nEn7zKRe5Mci8C7UQ1iopchOLARy1mdJYlWn4zZ+RFQjVhQzr4AT6qqqdjJ
E81XjlST4yw6qFk0n5RdEjHflNMkhVPboKg3jtzdTFXjCQ8aF5VHSHD4RXSZdTt9
GwhQ6oFCCTVdPLuFBevxbnwBhL8XUOt2hPwhs02G3PLqytRaeVNTJyjMjkovo3og
I+K0+3wuJPALshjSrM7X/lquh/uwSnVvBWlEUqt/8YpGblzNsSZE/P42Kd83Z1aZ
MJDiYxlX1MlTHXnHnWFRStxBB65mBZJ7xzDZIb11I0iy21YkR0LHPAzLlXFaNvg6
WXNl1CYUDfg/jgWMCHXY/ti5MGOLA0874ewONpKqwHkVuQBoUntNbfT73DiJj1AH
5fTRGBST3yLmEZAtIWV+5iR7LiB5FrzkaJLOz7iLxAV854zctWVV8oczc2HmRoKP
eO8Oz+7ks/JwlyUgEzwhcUahF30OSwYG/gQI4igT2MTN025BWMl6W+X94bKLdyYv
aR70/JWuQxY/0wEFVg3o2ul1W4yPp8AKQ7m6NvpJXD8Fai6d4kOVFyB5she4heZB
SAYruFcxwWRxGn2EHY7NKRYVKmMfOIU04SC+xYV9iF4KCj/KnZHmuf8DPZSOOrtQ
rb2Fa8CoUh9QkeYZNqaE7i321TTvp85MJ/dA8k3effcRWjvaz9VImq9DFSNZjiRO
FfvnlZAkoptOsjYmXzSKEN0fkId3Ud6AinOOFQkvvCYtb5u275rZ2te6nwnKp3zx
gvWPLII5KmYn7gmvKX4MdrA2Xcsxxvtf799ODXrjNGpazXfUCf0jPhg+zzIo8Uf3
ieY+dZIXndU0R5IFhmLZOZvd2bKLSYwbiINw7CR4KZvQo6nlsH6KTjB4xrkJCUbN
zOvLJcrqoXObRIt/nCqc4M9MyhMcJwprJh5kgenQ4/WPZ7zwmO7a8Pb6n/wz/NbI
QCZhqrj+hiatoXeJyxT3VFdZ2g9wmgpRgnBgV6d91kMpo9lJWLKffUg86SFQ+Tot
cJNiS/EJlBF4aI0XIpIQvZ/fnkgmvj7aGjzDAzwka976TNB3cRw9XkYxDG35zIru
lQV4Uek78YHypprMWJ/4uvfOESDH33i+WovDNDBe+iOEZRoJuh7Kvr0X7TmzD6sl
Eg/tWQONYPX0e+1qyKtXWtLX6hsym6OSDFEVi7+r/4vU5EHtOR+IUTdiIpbDdFSt
P996MgxMVvrvaPW0Hhao0CDeR0LckNw2xBW2Me4NvIhHEX9SXB1M5SSq6gM/ED6I
6jHapCyU5GYzc1nyXH3vEO9FQ0p7SISl413BxcMbL+Y9Z7sz4SNsMy6M3g2kdh6F
2Hl4JR3oC89N/lldD1Z+sNiHzi7OQDqFnL70rdMeamNhC0VahRYJn1PSVTFi0oKv
8kdp/JXDwTBl5o0ZUlH8fM0rpOCKUeMnoj1gcS18Q46NuS7titYRvtBbgnIHSr5T
Wrrns8gK3C4BH75a7o8K7VG9ftq6JxnXFkh0a6Tg857F43iWk0vvX4pyBO4kKZVf
SBu4KGLzjQpdeGT4+Jy7oA2p+Rfh4JkIbtF4qbjvt16EW82I2TwB/+puXgog5yHv
poUQ2YqWlw2/6O6MBSXR6MYn/gGo+woJxRm0PoyF8QLFdO3uD4lDgRvu6918tFSR
Ocj+AtTORPBVZwtm1/OF+2YS/kpIHbes2jGG25aUzfAJFSDk6XXdDbZupuTwIK7w
7ywIkjICtqOGe+r2bjfplJER0cAgibxMtnIBGMl9W8GdJUwH03KHNaFN83XYzvFj
WoKPpKxHtoPwSx121ODqVlykYU0PfnSDkPIlC5YqQmqMuT50i//qZbbX3ErX0rav
SZdyHtJ0dcmNy59fNLMp/G9sFXV7Lw+UxgHfcbzIMYjybWYpWqgH960b7MyR7d4q
2cr581KpF8VJ/2rnkzystCO0QbQfJERg4aATbYSr8djtFx/CgGnRCPSCIM7DbAbL
0P8b5Tnvm0ZTAbyyBCppH+voNHUB5ELLtxMfcckjO2x5kJN/qGOW0AsqOOGfHCr0
uUjfBURlulNC4ewPg2QIRaNH1dhNC6ib6aUHvDjjwsOQwn4ENy1fV2ftwGom7qMM
IhRK0OA+KyAOQ9B+UBCtL2XXwTXWGITtExbPqj8Xy/XhjS8p6qI2mFUbP5FsT8Vk
Kr5tfEn70mYYQCzxYhchsUQCvj66HVsZwiRyv4cLwAipQxaFA9hQ+s82rAW9YikU
gLtCL9sAwwDKrMNXtCH+2LFoKwtkX+/czycVKsbUphEbQm/On8Bis/9PvITHJzdy
yNxOXTfRAze1WeES4sHJztKbSRMi7LyLMycUomQxNd7j0rs9dvMwrNzzNakMfoin
9/YM4VSvu9SXyJMzgGFCeqjtKmnMhe31AqtWdQglArLC8eBzjoU75mv+IfVL9Mm9
gqP+nf3HIhTtgMjH2fBkPs31o0/yTGG9k0V2fEzl5p/5xkyuvnXntppzN5U8QM5X
X32z8sIxGg7PB8JNqRdjL/MjhGziikR5t3dXRWiUFn4pjVMGQHchEQ0Sixj0ElXB
q4EOi0HJukLpmzGv+tPbaXMMlv7aFGy1S41C/LHsCwH8I/2lisV3J6wlupnZ0oPg
sH2RJiy8Q9xCgChoyiO/GzH0VQKY3+V4+wCYqd03D7mvuQGd+/ZRWFJrf8C8R2mK
E0HcBaUSYk/6EdvEIWf89/3GwxT7//z/Wn50yu5hoNLQC7ig/3wBtINlF8XAxYLT
/kHefG5wVVYBEV2VefXR5wasuzQXPCoEcTPkbmR1P9j+MRW5+//O2EIGOL32KUu+
7iUunR9sg6Shg+deKkWECC5q4UwK2oZJW0Z8OqIrk25fZZZDMN/EkouQawTM4p2L
qCMVC9T0nainKMrbW91hGZtXQnY88BLxzV5gkzyQD86YWRNvEgWF07A7IHFkhO/1
F0HhX9eA9W1Bp4iVXmjCeVmOOSJvY6PbNJeTCGt/bUKnWP7m2sZLm60SfF7nCkYG
OMgqQxkrJpfXBOMrDcXEubczhgkP3olvShfWG9uMfLckFEFNcDCWDWGYQpQh09V9
ITY0/TPCAps2GtDoph9MqlGawcpUHP568QXSuPqaeIRZi3SpLNxUJmPcdhuv0Id9
QAk7OxqvyAH31s6BuvIgtHwUoUpZlmVQ5E2vLZl7qIsI1bCoIZSM1NzJf01sV4iv
bDMtJsMZeejQLctCV14x/tYP3jqvVDZXwNgUUmMs89mPhN1c3hy5NE5hxjahiqtA
O8DHXWrF59POJBXKksM1Dbxm0um4oWGdzgTkJsWIFPxI1zKFn4UPPPTscgIsQ/aS
bMnS7ytfhCd/eMrfZ0ZScRKkyMbRRgFuZvjtOtsRnVGj/UaIM7b5AAZXbbM0Sd3n
oogTPAJ48ZJ63n7MH5SB8qRw//gUXI787O9PNG/awEGEetXZOan91XPGQup2a3wz
jWig6eyEb7q5zVbnCgU1zCoyHkzuPzr8vVfvYYx1zgn1NsFKr2qVAi+3xBxyFdey
DTRK82TjpVtzSNFNFVGZUeuCCMp2sA3PRWvUBbTJGE4PKOfK9l6fjAOe2ovr4BUV
aiR//5/FGaH+7zAHzV0NyWrR7VDang5Z7uh4TCKTxkFeN4B31Rqa4/tGMldA/rGs
hgLA/KiYaP2JeD5wcX6mMEAEY7Yrex2p8yl12Cu1Ugoe6rUz/uowa7i5Dp3mc9nZ
dTsr6mf4WznzbR3JXrkWBxc8KHkH8DaY2mNVHok82o5Jwu8L7vtH44NdiZ88wQyF
N0YkkWxaxSUncMWsYNsQBu5zkr0JXAKNbN98qKnRz4MDh7uQbQcKQ8Anl0IVqIkp
lv1cOh6SxZeHm8Z1ZTCzOdXV//ppc0RrCMCDDQbSyBS4qOWs5o4RKeS+yFxJkDyz
R5gCoDSgaGfwzvwR2qyCRMtES89gywan+oTZCkC1JB2ehi3hvPoVXjXG7Lml9S0w
rxyRMdiv17rOi++w0bj1IKXU6BbwU9bTd/bXrz01Up7qIbnCk8Rho+lXj/HdFq0F
tGW8Lcps/cil0beA3r5hx+HpD1P+XNc/YWjByzt1HxFS887p36LVQMmjjjpUbXqM
owHCzniyFu+OKEJjXtgjoC9nOx/qF4A10chd1/5aARXl+SNj+e2SVayoY0iAKlj1
8KQ/obOIcNfA3ChIJ7OAZL8HjxeTO3Rd6iNBHbUvpdp50Tx3gjAWnzQD4hyCRcSP
+UKe31GncziJAy9rdlL3y1v1AtRyVO7oyU+h6p1bRfKk6ZHlHZUnc3VkvZmuKKoC
6jf+3S/3ZLV6A/7Ma6A/P99QUrIUCuZYn3YuQLwnG/hUVQgDoS5sLywN0ZOf2qf+
rxXCjzJ2jJiv2FXaqUM1nnX/JZymJ30rN3NcoFppW47+yk1aBSPamWlpZs2AyzUi
Llk7xuFaomTFMp7mgUL0N+ohobMVMgc66zxXbxpNT3uq7YNOVho87mFujn+SFtmE
ER6tyPCflW32yt7KoB4JZiBgurslQnudfBJRgsg2CYiSw1qCEqtUwkf+VZgk1SZp
99qecw2CtR/5tGXBFHUXSXR+s/Ondnts+kdKhxUH9jNpB+L+ee7kHC1TiQ/Zi7nQ
m2OFS8WryemDSZ3XrRNwuKlfjUSOCYWfkC2N59AeiPzSQ07lg/NWiq501zEGSAvr
YvrUJTZaIf+HYRMVK1Ow4LeyoGEx1zUukri0UBpH6iRCSl5fFDWEVKjpEp0X4oOi
B24/Z5yFEuINQYJLLc3URZe6ED8l3anbNeJu4TCOy7l9FH3Ecq4p1frL/JNR4mIN
b3ebh/nLegQtY7+pXVLyYIsoUgbFxypVBgNVJ1vShqSaO7CbnzvedXkCSQEquqoj
SI3t1ixGnE+HfiEajA30FY1ieVVi8u8O1QF2T7wvIzxxR0gO6iQj3KA9rdteQ+if
m1S2fi5Z19mNZho318KdedE8qFnoNp8EP8rWeuSuc3TU8mo0ow4nghvcTkM9ibMA
Z3GzqZ3ZZPhEW3/D1yxvsQcpSHhNBopinASmDTuwLLskavQMuMyssHaqE2WxkDF6
VnjvGww4IrVdbIeQEBk7ReUzQIZA4xHUZViUexcfZPzTYJuB6D9IUL/q+iYABb37
0pVDhYq1SavT5UY5xuRC3oOVqxXEH1ruCp7ZrmiSX5pZi5ZfzLDsDb3dW0Sxq4EE
Q/hJnzsiRXbmNXJwQqWATAgkWBYRasbfE4MYyJKPFchfW0mac/gmggygtov9Ogac
wTVj2AHO2Tdip1Gv7+RKX5neUCkltdNCSBfZ1ASZLwcA9ZvOi8Ge6RU6eDFXsXsS
Ox/4TFGlku5l9VjPd/3x9N4J/OkT6gCNbh+4pHDIOK94d9cThermBQZ2mXY2mQeu
uBo3yzNrCBzPO2UQqeWa2tbMs5cWe5TLKPO+aBUpQ3RhV05fknj9Cz+XCCsv0Gdb
TaBVVPL9NUyeC+GnAiz8KaqoZqGPugJqGVk5mqCH/MamjwXdsALlND/hmrAorNxp
7ELEG/1U5+BEvY6rvnspLrr6MZ8JhDpx5EBBAkfnWejwf7/SEPrxlT39ulnE1UYX
LIyXW6//sVp1GPgCesJ3OxT6C91O8EytkaKkpnraq1AjKYpC6Qo/RIT50F7B1VKq
l6RbYYT9KDusgvphVI4fEF/CN+fCBphpI1OKl1YKrZ7L5Jnl5Pm3qZCudClhRKDK
7ztSN5UxqkdT60v2DxZXDGVd17zc+oFt8DFhiBH1adySkCJkG9DzAyDwkILtQLGF
AGbhckaT1wmviHwcedu0R5ESaf/VOnWY0RFXFG7FC5M2cvFN3GB+sOoHu7HGSPDs
aRpP94abJWYA9U1UUr4ULJQbnpesYs2Y6MKfhDbjcTzkqlGM0+CciDrK5kOAk2Sa
y0/BiUPDiqLim2TCw8LDr7CS8J4UQv7KkRk2hfVgI9AF3dd3+sQNncdT9SHBSGa4
s0ZCyoo52CDTVbIyqsLd16XoFvFgnDsREyqTNbmq9WLSHjjaZyPOLOeMReOvw/Jo
CTrN7kQlVFEWWtU/SsyXqk+ggTimGJRthAHrh/nwE+YJVYR8Q41YilunR20WTYWR
OQplFOWLh/wD/wNdrHmVEYdJYNUi3vVv5tlvECN9S/KPvnEUK9ezoDI1+X06nVT4
t1PJ+eeHk6IOQtyHRGj3k7xWVzd4cqNwqk5TGQUWCkgWxk8ACBV2l/YXUV4XjxcI
8fxDx4X45isi/LNDjXu9apWomgQcu0iQj1t4DsdnMPpDUzgzy3Euv4qCIuZ2rs2B
I1F2TPJDFMQwCdBfnOiBfvqXoaW+eSkDJTW1ydhGldGuFo3s38PRqLnRUB4bzEpe
8bYXD37txtCvH05Pii0H32IXBvpl7JiK0L3/Rf0y0/yQlo2ELSxl3gIpKc2kMi/N
BNURCWdUvNj5fi55SBNPA2nvWu74Kg1SN/42y4PUm8oceic5SRvLzXkEQJQWiCBQ
y1Iah9Uc/rIevf7+pNxNu0qOiHdMdf9ue5NBuRePAyXmUxBIVj0vYn9ZyvanAaBQ
qZDQX/Ch692mHbyUPU1g6OuWBu/1WQwoRfB8kKOh7TSlSbmPyJFteD3gAC6+0qX9
J45cf7O5oKe46lxu3By5b94LC/TZjeADzFQNBYJIZmVJLlYIWG/gVglT1ZPXhGCW
4R7+K9geZszGjPYVs7dNCxVWRnP56ZmqsokBwrGvl9JSgWyEo7iPGtKCds4HDuxd
5N7GwD9HZuhGkV9gDO62IJg06vtgndwcKLH7DFl3ALMC5VW5ZqsqDPlKLZkuGBpc
EWMOpVKVXtNHXgoszdxZz/oYszVs51izmQKgzEsSqGG+xeQbQTzuzBpsq4ehz+jU
S2MqYWkA739m8gVyY6Rbn5TPwN3PZU+U8m0OMs3Qk91vws+2l8RZICqxqbjQNnK4
/uOS+KAuCQ8ci0LfrzJ1E0UPmh6w+L4ZLTVPu0ewkkpqvK7MG+E/hV80AxaAPiNf
6ELcVeiR1y8Gt11BGcBpaw4dzDrsRrfQkt+2I2gtZxjFJ8jt2MmcOsLWBMULIK5p
Cdcy4CCnZ10zWrS0gz85D9WMwSrskELdmObKv/Sf9tvMJtdsWnaRjF042sgaRye2
yr4N8bgaolW3jzX2g6pLc5LUTHwEdjK/6zw5usK9q1BDmVYBhqNhhxtTDSQnoC1P
EI4qWFJOkREvgaIjsQAgtdLRBl9kN5LInUWKKsCpgycAfn2VFSBdg1WIwS5oAFIX
c9eSCkuHPVa5glz29/U9N0w1t2iaiCoehIJiyPUX9hsn98t2VuF14rfjecmsV9Kh
mRpns3aeygYnbFoZlg7X7BmY41I+Wz6ruNpv4NGb4plgrPZtDrscyc6une1LOJIj
FyPLDUELj/xDNSC3O6/F3mHyxIHgFjII9dstFuyZKEmpVF1CGRYyZrPJahfEYHwM
9rrdpegxu0dQO7J5+YZyYOf4GrA5IGBQics1ppMCZwtApduu2sr6x6tx7YAftC2p
pHb5tuBVxIeflO/a3DS/SuL3fzABtF8dWVcIN6qhr3pn43hVNkIXQdgkwhnn7H7N
ZdvZy3vl058b7GpOted3CyXSTnM7cE28SXf7J0cFTkchPCNgbRKv236HzKZdcmHX
Vww8wzURJb4SA4TRNqUeOt2mWY7/bwfQxB1qe80y5ymd3VtIf7VzAo3xU/5645hX
IN1TG1+Wosz5huX0c3HQnF6wdxm0y0JYQSsJ3WmUF4wX8pVp8yP/1aMqV8//OFRX
b9jdV9aIv6AMd7PRgZT81bwC7FGebSVMTbaCQrZAzZ8fl8grkocz2fPsM4IADiBn
Aj8h6QBMhB9hXbI5sFDIhaVEBwjE2JmNjMuX8lBS+6J+7NquhFFnFV14se0iQcsx
f7UKq+i/ZlHsWPQ8tpiWXtIJiNc9YgjO9pzzWzTJwlGeMdLTXNvFx8yzuLCLqq57
i1YTPb6Gb9I20bOr4raEZnsU8mFrz3Yzvx0/DMQSgWaznNs3UsVnGDjUSMmel61i
J+dibtig1J8Y29jRiJjrP6fuzJJSLcBHknKuKgJx9cWE6bRH5XuwBQB4bPPqGUX7
O4Nbt0xu0K8lyqo+S+xXsh/4AvXvqUsWRkkHNvDtS65kep0KLKhtoc0pcnBrK88V
giDNVMkc7MKP9DCY1VvDWREh7RvlZJsGYKDrSRv+jBmayQH7A21yAIXmg84267pV
0kNm6gVc5fBkKol+NOUJvWRw5aAl+CrfTSk2ymJCpmc1T63MkzZhSn6krLGTHSq2
FQhuYXqrLUT7nh/0O7qniQFK26hlBgoPOzetdhm8z5/pM420F61y0ZY01njb2PmA
5vzWkLyRE9WIuLk1hBg4tSYe//4psE2IjWZ5oXQiFxlCVhrG1Y7Xt7yJdeIftEXA
KCyHxEvDMLnFI/WnMAGqeFvGjXBF6HHywsiJh7OmNyx+tH8ttXKZD05sXz7aefbp
Mp+EbgDdj/yTxR2ztjYlNUTLe9Unjkae8iqL+qaba1K9UiGX0afQ2tLBGTZuenjC
/zaM3PGpbMklA3UMpor51b5NR1l62ymRueLGlphithb9e+P2G6HABnemr8htxoPc
q8vsZ/981t4A7LwlK4FKWPNUB9IDNIKjb/5lp1Q9hZmcaQXI+ni0eXy6EeHJG0DO
5nOkuo5yiFgayXNF6LMlHTWrJUeUTjT46cwjH2m5BHQBqy8+MXNZIxHVGKThlli9
PKeew/zimc3DuonNP/5Xl8XEtwPSFREBOF6wUiPXNC6XLXmbMmihEMttfYy341IN
vX8jezkqiqfHdX69Qfb8teQnyGh85a9fg0S3ds1nzeqrM2qlp3Ll+qcj+lLdx9aV
aFVUZxgTSpHC+TDfmLEJnOXtP+Q4POKGU1vVcDgzUBQtj/RKH2oub0VGt3ZvBZRA
e3snLjwFa+Sb7Z3w6x+TIpx7ZE3CrnZuz6jUqcwoc1eStIiXcu6lYpvbWPpxFxYv
4JeEy5bGNgzt0ePkBxelfNDMleYLDWwDvZiFJg1ocz7rpJ4HjZ3xxgBI5FrKll8q
thpLGGqyktNbGqIHx0+LQk5CzzGgVHFf4gjXJRSl0YvIEfcHXXNHNp4IO/U+3s04
9hxwiLo1ACoixwKGIPc86d1RUEG236UG51c+Uf3egbr0RTr2uTf3A82HAS59gmbv
npvSftW/I/ck99ah6cm7pQYS/dIVvpnR4tigNsP0skDSfg9RtUCLZJfF5JJjPsgA
qFTovAmx+UIf6u7QCgmXEs9uVuAihIVx6bT9P7MxmHBGrZCHaTOaE+c9013UToxA
Y1OgALiE51Nx+bZs6GHSdbq2pZUSMPlNWKU/rLrYZebv17S9tClIAwH9RsoAjuLF
Dx7x9fp2hIkd36croSaY4axIXV1Um95v0T3xb5oEjmzClU9570uobyXjux0utM+r
nNQM4LlO5OKwX4y4cK5V86W9/wnzZ0X2V6YLBt4dDlUS/2Zew0Z9aA1ovVESwP5y
jtnhEl/Bd/zBgW+APwRU/Bx0Qwi8hxGYYHAhF6NHNnEMGhUZsdOM1Rll0ROx73Fs
XZLKN5SkbGvrrhKNbuYfAL8jWgigGXIDlD6kG2ube48iD6uFyzvnvupk6nYNKaTZ
SA8dxugvr92k2WDpD+Y+J+J5dH4PUK8+bMMUWznXlP6krg6kGibW3MRPow98RDZh
n5OlFlhzphjFkGiabt1ZSo/fUZRZc4/Yu7ieOSpRvyZL0h0soOHiExot+Xosnp+L
ixFKJv5gMg5X3YNeu21yG2nvZMi5ngb1iueTqBgHSqhYqz6eni6Dox1H0hsO5/6i
mInQa5rJEMpuelfZfQZ+F1u4qMd6z+qDTiUcWM4PSrHLqQiVSB9TcyPjqk4BqAIE
Vg4wSuPVR9jXse6AoTQnaBs/ayBAPZMAvjuggu8W1wMGmUHEn6Bmv+EmugrZmKyM
c+Uudz1ubB1zXgGnHc7XceU6wiWGdLK4GYdieETfHsPZ8lWqC8nyMO6UXkzv3PtT
VCHCDwy52qnWb6Tdoj566/M7tpRrQeKtU/77CFwxB/o7fTzFtykAk7QbaSmu7Ghh
9SWgo480S8nt5MTDkAOpoH/e307stQe9ge5c8OU3i1OTbTg7V5UI/8rSi/fX1Prz
m/4SOWzkzDhoJn3REzs8rz4z0RMW70ySnuj4MQOtYkGDwN7llDunggJ4lHg2UxIY
GCp1MznQ6Sqfl/7hF6CJnfkd7/Mlygc4mAmcp3YemCbMOwKT9mDBB0JdPF0/NeDZ
izdndBYXcKjm0pVNvS4zf3KY40gfiST8RN4bqm6nk0vxJG1anYMZQMhSp0ZBG3Fm
4bvVd1y56lChe41KLFwMJXZvsHWl0jS9AS83eQ+JttbQMf3PyUELXM5or34oD1ZU
79BZPvwxwdaejXj9/am6fUJtBtJWkzEpBXgqkyxNNmPYk6UZRe+YeyNNUeK6fK2c
VU0nq3DbC4yx0XXj0+3a1n8NmFju2UyGIvvl8movZwXz+2eSs0ZaUvSrYwyu/doK
Aa97ahOGpoltuPHUFMhyLXNTwg44VI3DOZjuu/grYU2PKO2eueS0tShC5mzWKveY
UQuUTqj26ixqNUwkpqkkWYG2JimJnrN0zjJnq5+6iSTtJJM4Iwpik38diSRpa9ms
xYJ2r+xPwy0M0HiY0Jr7Qitx/ZwzprvQf2CF89cR31YodVbt0aFI3pF7UxNVvx1D
mb1tQm7gXYYDFQ8dv61gHprFvXTawQNUxYFb6r4c22Qtquxd4TjVM7QCr2/Wq+ud
xk7NgdqmJbJLfgwy1QQY3gLYBI82+IlVoyBnFnwKTaVCmyftRMcuLl0WDPSBhJ0k
zVzFk0agYjTsvm5SpK2t7CMmYJzBiSAXP2KicHNvDjTIGKtXPfcjDfl6UynTFl5a
YkiPLoh3LUD475Qr+FpIT0jK0ZUd67zSjMfnCh6Tl1ks9798S0RNo8UvH8qqqpGL
opA1TDqPNmkw4psz/Tms4XtaqRfcPGFOEhpIOrJH0Fnj6As1Rj4nqmQbUdpuSDmy
Hg357Wj3LBQKCXPbBX/MZAuyx0DtMtECTaRLvzBrKvMIpz2Z3G9DDuMhgqVTXV9/
OIZ8CFbAxAYeb/yG589d5FTJWvnmzikBEdRVsTsosBuyokRDJpGzpUlOYfsf8/gT
6dgm+0tG7BldQjiPl7pbL6PhL5Ysh1YNTX0L6yHXyUEArG6NVYDSMynBvIRdowGZ
Td+la9woEnL/dFAERtMzgUzHlx4d606snM+jexm7zKqf0V2rD9SvJWSkgOa3e6Ls
VncME31yl0iD8oFcx/k2mcURaqdwT7o3lItkdNuD/TaDcWN3Pv/0IAIlTXOKvrta
Iv6nV+jAnQiW0kTMCIzBaETp1tt/px96fdy/mPc3dnkL7atM6DQ5qkmt5O6cPMjZ
BhfG8qM2aEN6mfFTaHUjxtdgtX/j1+bfrlRnhzgH/fEM6MDHl+T/tOX5rw/tv0mL
oLQTqSBT/prepzv6BVvKQ28SWYELPc1DtI8wta5A797j7Ln/KsGF+gbVSQdhZ4xq
RN+xo407Pvw7ml9KtvxCL7pHNUUBhPWeS2pzlKRgKZmpq6GEU0agH0M0oqGxfmfF
lIdNdH5qcVS358wvytuGixN9b/SRA/i7zW7r8m3R6MAH30UV0HqDOswdFYg/5JYW
NqAtb1wfWVwhvk7MuhZJtMVApVRUHdhALlKV5eVVraMssuKWdGZes1U8U5iCOtdj
ZdhSeeyorVgnQiHtABI3vn72YJo7GizBuiNCLCuuO1B7kzIkA7o1yJYYHd5+/fyt
SO5YP+g9xDKDKylCRb4JSqKV9wsEneXaCEsorDo10N5r7SAPbSG31u6hOPBmQaPH
93qf/ez7qfQidD8dlEKDS15qUOP3qF+AmQkqzynWXVwTzS2lLWtAdiM1oghH60Hr
eQ7YwzW5QmrABfgGOvHa01MYZ5cxKmYPmDjAqyel+rrjH505duoTFo4c+ppBxX05
cnIGpioVRmK8jqsTStHYYB/S7oD0LEWS6G/cg7ppbGqqRoLu00GDVWfLbBUyxPhT
fQuRAD5TjXufD4pe9y9XHWI/1aG4OR12aAYp61VbvK8bsWyHZh1MRdbj8xOXFtKE
1m2pz0FwPi+2CClPeNrsd9v2Gr7Q0eJynOwnv/OhS5E6jtuXY0xBoWuYyhANiljn
/SUyiTW+iBiIbZuNAZBwYinGkLpiO2TkuQ1h53nWcKipJvyDNrHGgqVfvGmi4cmu
lvmvUW+yvYxI2ufA+zbYhy1FAq7Hg6aRx/2lzuYhLzwDDu9aHcN3kHujTAaTi/q5
MLUH+pOJHxku4Ndo/zCMnYgB0q9kSeC8WkYPzjjHXU6ZiHa+j4zgF4bAJISlESta
tyJ3/FmGWDkamdNiBdmx3cuUYStzHpKqyyjZ5CM0os2ZS/ZKtYdS69I2Pqkx0SE7
7z2UZoVRrg1O9wkrW9II0WZO90aSKBf9pYRmFP15Yh9Wdcrw1NfQhvBcii0/KZ11
jT4E3KlAiwms3Kghd4LAhSbuqbgIgWmoat0r5xe9kP4xhZPBVr/m384TIwng+V1n
`protect end_protected