`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6288 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
yB5UT5oQgw999PzwDg9vEkb04KIzZjM+3WJO9pCKr55wuMHu/Sfwcvgxcmjpsn6r
iUDXA975DdowryPwtNpQbap7R3gtR7CMVCAfljL5XvQmz0dA86oIzKErLxryc3DJ
gdBiWeDXbyEL5ksapzJKH+D1HJ4H0P91IJ2zYDiazvrSWz89xLdpVsvpDVapeHB4
yZEFlYffhDra39AvLZCOWPEMai1WTJlrHSzVfQaUyO/Iqv8FgUkUm/Z/44TmPP2f
+7hZV7YyV2d0s1ad+sT0UJRs097s9r0OFwSf7/Cm03yIZkZda1sQsJzgYeiAl1KF
PBkPOvGDsT7dHK+K/WwShVNsU79CSYQIYx0Fvk36RwcGb7CkaCmKxnhKuSGroSw5
BJgvFZWhgSMv+5u2/madx/T5NpcOAd+a2kRLcScbavewIkUBY8tOaBcdgWHWzXOK
STQx5Edr+vTg1ekTeTg/BDT+5Ym3I6uCjkDN/xthYmcpbsuFRNd5qQU3Cw6FDJ21
TarOK0DL0gbMIk14ugIbT+5tqc5Aph7wjxeFNDk9rt7vmq1FI74y4YHpPFN6o4LI
8yATL1Wh4LHxv7eFcRXndckz1EtptQE3TPUhJZHkOOZ5Mx6wKkT4GwTXoH+NQnBv
kVJZ0sO5S1ox2IXFFp9ePIGK3L6irVosQ4f8FqDeEsmokUSl4lCJKijFP4xTlawg
ofMxgeDyapXTHH63b9Jfn0KYSvSNIdpfZ6sX2zcTAI6STMrK9ujjbVKWCjpQJykl
/F36A3dHPWTD4W1NoCkT93ZjCRMIZ3IZZ18L7aNYr6rhciRnRl44BUumI92VWAjs
q2SRkfqmNOt+osOsKwsfIBUD1Q8/ga9ie+mjC0eLyqXUNDpdF9NJ4KyHC8Ea82+N
BkKPho8zY9ScRxq3s3Osaxj8D4warQCqZ4YN7c5HBDlavI7N8sBK+QmypcQdgqeM
6UmJLBtHSqWuUhFL++b6ttPn6YsK417shWPQTWGo006yYKLmS99Sm3EWEk01wTo7
P6ePubvcYom1OtNEC/TUm0kp6OJa/mKEelEFK1GE++kL4SFHuVduSPW4qx6ZeMPy
sqYa/WIQM5NMVPTgv8vVQPwLLZczIWaFwm7jO5ITuAV8Sj16PPpT+dNxS+oiwGWT
9aEnpAASYO6TcOvvCG7Reg100yKV8Og8kNNfBu3j2TzkWYqaYag6uKwMM9F36Sgk
OLWA1NcxbMHKFgoOkGQ4uG25Vr+If278P04LhXCswjjsD6x05esQXsZjOKNejFha
xwLNODB/pT7oKDc1wMqi4IcXdWoYcqw0lBYLvBUlzn/pLZXL2pLHQLT10KLUqTIv
+r+rsBaoeJP6em10FzFueYLvJTnNxJIaEXnyUnk536XOaJFSZafTsWT8JpB2ItEo
bUzipQlHasaHA2wfTbgevM9CLQZxWOTmg3JQTIgBTmJ9xmB8k72KOJbPkFaphc5N
cFo/oFn0XLgP4B3R+wcmWEVknarjxKfzffn7wT33MHVr2vNGsjWLaTSc2BLIJ++T
Tyt+27NRs8KVXld8lWbIYJBHYdCNhQE4wS8U9hGdGfhsnmDp4d6XSX/dNpHGEFEs
P4koEGnB3CohQ1lgJFURXwhCtoBObDHpBBVR9F4xD/OqrVRua7XK3SkXNOmdKJwM
K+di2OhxIvfqYxRKZmB16PwLio5k+MhO5wYffXbMg+nmlg/O0qK5hKO8ru8APsS8
9Vo7+ua3x0EZiGiW0tHYXg4sxGrF22gaMW3F+mV244gE7rx8MGwsKAfBD0Gsi4lK
NY9VEWwZHzG31CXteAFOz4i73cYHPXFEz2vrDpzz2v6Lke643QYMiwHVqHnooTD+
aLNr/sB1ofhhKxPToF9cpuCw4aNGjuYI2xiec1N1MDvYKgEdNEUzdCvdrgAJeCBz
bb6tu0OdRgY8Ni6cXxtW3gce+P4sy5WNE3vAPbYUhzkf0PEZ29Xx/3YuR3WAAedl
Jh0OR5hFj2GnCTbI9KqhP5GDubeosmQpFs96vlQSiZtedM7Z3/Bq8Bobbb+eLz3s
E52biPvaopqoXwLGzBxwGaQMhz2naWuTHuhhV3jFmzJbFtRp9BUtNZvZIj5///vp
6XIGJCeTAfgpfG0i+9ox/mifuBt66rMINPqyA4QWku8C29PBY35YYndlFaE2HCqx
GXPoz068bJoJvtaFwU9b7JFCwL2QZnZ6fKA239oz98cjQIhLkW4s0qfmVhRd7GQD
Zsi6bL2IZRofEQj8BhA2ZEu59I7RpQFYV3ft4qHC0lqJ+tiprkspcsDopf0UjHND
Heex2vj5S9HCETM2YvO5S1QoyBlXy4IQyGd4udHPwKgbPiB30qRDr2X/5LWPYQN4
KcIADYzA+Bz0bn9WtJWSZSqYCDRTylQYzkYv9XGkbgG8BsVB7X0QthR9HiaVpryB
k8b4LxEQVk9fSbXVsIDTNkUkbxFparnWxf0ekt0WmH1QWZMMaIVxOvgv9EsJ3iH5
3FK/kfj1dopODzHctMqMWXR1XH8wb3bSCyGbXrHtd/Cm27cbsqD2ykF4CThg/L8v
t7OugSo4w08wLWuBOUBWKx4T7d7ohj4JDrHrYaGmtLF0jkLIM04rfhnO9Y2mWig0
mA0Dy2NpxJm6xy9BRKUug9nn1odBPAgMLnU817XQJ8fWZXpnd6r8x9X+xEPef6xl
/tTjwTrkUqjRhv93pqTGA3YwBvl1KtammuSrxvS8CUPmEDNvr4WzHYT8ActpBNoS
91a+ZxaooIru6WdkQ7wkP6rqjvAv6dpVhgOtUU1hwTXxjpGZb1TqQb9xJPNkl/Kx
UXi4Ath4C6n4QZB6DyjpLlYb0va7b1mFUR1c7Ay6w0TRDmuuVIHUkuojhj4sxGb3
LUezHuwfZYbL/DVtTWs2ooOvYS06zvNriy926DFclA/CPl8W8V5A9/E20IupzeKR
v67HhI0ku4360lgmXhAvgEomuXnWZjECGPNEs/sZIWZEwCOGhpfleZZKxgo3QFXL
NRSuUx7yVfd2BbKVaRQsyniJ/znvLyaYLcNFrCXmT5Lr3NXPZSKJrUv6huivaK89
9Y96nnODlU+U0P2D8myAghelw9Lx7CHC4mgLKFLisr/weiAuVPV5Cwn130Y2lW+v
I7V6S+Tu7k0KBjDPwNATrHGFU9injtAIObJ/89qK9z/gE3F6KiiSd1bhcokg0awN
axMIB6x8SiMyE4blo54r7fPs3hbOCSSvrIkBkCbGscJL99+TNeGct+Yq2nHeXVEV
/ev0uT36ffkjPDh8Nnzba+cmrpyfS8q2Namta+M+9O5DbgBDQ1VMGtTHtivsccsZ
zj1e0X3Z7e+8Ytp5c6/7t+CSrmWoz/SS3ORasDjI45X96TsQWKNYl5VeiYWVKJXb
9cgTNSfdbkuymXBTL7YaAWKF55fYm7KlkYfcC/IF7qbr/zDQP3YuaLm8f7WzoWRY
PDT/llYto6tS8pHn9F6bqKsty7ZCUeXXTmzim/DwzUHu/AnYeFrWXlZ+hbQdWeFM
vGLukCHHRvjNoN0cBykWShd2iUMrInuLr5MNiaRK/+dlgcJukCnOZ8F5fkgDHs//
LFGg6D1ZGYmL3rDfZrC558+0h+kcRsOhB5HtBt7oHse3U9sm83T+IEzQ8Rs1J6wz
e9lwrRZQOk5yeOr9a6733Rtd20iSjilZjwV5uFOTCGjo5Xl+fHc6krJQFF5vh8zB
ybi3eklc6FdHmIn6dcCSwU/f7ue1eHBq3x4S/wcRwnm4bYe+BT+rUn78C0f9ASAo
s/lEgu54+qNoqmFQ1e4jBoTsOTcoHnHTKB54DJH7/5UgN7x4fSK/PKvsjAESuTge
Zz0Ye1oewJfkYjo3vVu7sjOBQNEU84S1qt1smD+YpVoWI9AWeM9AZh0xlakvBNZw
DeYXO8BRML0sBr1EugCt1wfMIwAd0tJo2hgL5aNguBX3WpOUJBPwtsuIBHR799Se
Q0NL14uhMpnJ0z/dvGZ/dtQOaTssHNCxWXc5iWGGtbYnBjSZDG6gjna3abgGpp1Y
E5LSk6lmEZuJjhJSsm27nTIExlX0Wv7+kgBSaAM+UIH7G0+lwUbpWntegYCVtGR7
ugWpzyXOIPBe2BXsFk/kySzaXo9Hzs9X37ttkDERxPURa7viwmoqiwIdqIAHhCAY
Um3GRIrt3NDNPL5YBjdGkXi7RbtdmczvvzTUy0TRX1tsCYhDfjBtoNSSuPXcVb2y
o4Ik1sheDzCirk5Pl47yTq1jleIlVT8nnoMr+4KS6XRMMOsKVXKVnP79JJVYFztb
eWB3PWDWlG695b0eszSOi2Y3yj8V6mRqjJzzEJ19USO0Kxk5lAe9Nc9zryQX+bSj
AE4IZzsieIGN3z0M3KV2ITRI2aEXObeKnaQAK/rsrRBU9aeQPDpJmP71EcDCgmMm
tiu5AGPLzp2HYoxB1wsGslZWH/Ml3SWnxTlLKnsK1D5TlLIXKYrlh8v7UOoDDGOR
HJqoBj+Qhiq8mfKVc7KkYCDI+Tt0guX5MMee7uMCD2pQ7NtNyIXsfiPWUYX+2v2R
9ciUCKPBOHudZhbGqEDU1uKaCo1ZX0ZiuybjPIp+0StyVf17ecZIzYOQv9wksVzK
GpKCz6mwvcrEzd+nYqXvT55VbsHP2dsZlq5JkNWJrIBZPKTN99dJ5A3HYgh6vKQh
gfidMNHfsDCjvpd7lcsYzgNqnXksgB6PrvYm5IeMRZ6bWu7yyPV7D+t13tUgQKkB
QujU/x9eb7/MtsArwARbmlotgRA/bidqXal8GDJoQ2cybORraqu6FI6AsFl3KWVH
1Lwqg7qzHtJVT5zDIn2jJTrquyOW8Xe+Okhr9ZsTu8UYmcT2ZDKOZ5erBkK93urI
ZGlP07rD8vpy7/3z2cUiqX0puaTR6sEktE/V/Bq5yLnirO+jNXQWEGKX7SW1RRrP
dgS/MPwsbz3BkdfDUDcQaoNvirfPpCbZjHyoaglvRMh8Jqf9Dzfm1/RGBAQDgab6
a9HXfjXr96gldZB0e7FKTFlVyG9uDuBTXa/uDIU+DWzojCt/9d6SToCdXV2Q/FcT
vtmyUdVcakufS1iQgPoOyTzsY1Te8irEZgT3FEYYQEz0QX373UFIDw3PF78rpOgO
W8AaFnrOeQbgWw+SlQBM/GhnMEDk+wL2JuF5yU38Ty4i++1f5oNDSQm5jcbakpDk
i+2DFRJ4fvAOfWMkQqJhcyflHSnhpJAc3bNSAJNPB4xvHhJqdi3nTWhOuV1nzhxv
mAeH8tHfqVp7JLA9BV13ryOrkHfPQ8drzb8595NDZY4Vbi07HGJx08TBeNPKnHmV
u2X4dOVCqcaLjOj41swezd+o6D+3vo4h0C6N6lKFtYxlry2buaYdJMBirwXUxZtL
z1swMyVdIb755N2Pn5egmHAQSIESMJEL7Bfz90W3DfwF6bslqfD/qLnaAjxLM7GT
5orgiRGmeCAwvAPpEbUICq2tplTqqPBNh0ONWq8JcT3195eIiI+Lbw+Ea3X/KtZI
Oa0VG48DMSgLmkAGXRSm8fndaIrdwc+VPg4vkJ+uZiLccY0vqbrbSRSoDQGvmNdR
4pXsQ2VCdXYguxicsl+v+4sQgtQKaNvkJ6kmZU10yFrCc8cIeelyBYq3jVU/aoSg
1NaiwEm1+EgrQOuL2+xs0EAXVTIDuGTwCJx7R6vuXu27i1fRq+rFS+tMkpuBL3k3
px/g4ToR9Azrf5ekwE1fRRIycSbFSQee8jYFaOJAk+TIO3VZRaOs+E9NZZplCP7J
OvhiTjbexhURqp2g3gRfn28/0sa0ifPIo0m/O5QPXZ7z7s8/ss++mHxnnBitGPM3
Onf3POiC6aUoXsdLTtuIefVg9bP8NK5E7pPIMpPA1wez08O7a0HvWjQkOKZBGArz
XeDLnSrdVh+cM3ZARm7D/ad/8HN25mNv+cQZot2rMfiqOlLX9fT9MQYrCNYjyiRV
dPlJnPH50ynET16BZkv/FNappDkzgp7NYR2ZSEJVaCGbr4C/As0pTBsw5TzFS94H
1Sp4enBsijh/K1IKsPmuwpO/TE2ZIHFYHwqaANjJR4XFDhWSSErN6SKZ7K+l8e+G
Vx6w15j5GCLMy0HppGvX95j9sVHsUA2GEC30xyrliqhygCJNpX6ps1cExEGEml1p
wVtEsUTzyljQ2ZEpp6jGUwWSrfEf4aUutPCZs09jMhYhCYxg3fGN/92z4Hw41ERk
9EAG0AX8xM/xuzEWdg/0++xwu9JtfOVeq9KQLltwLskr9dTJCkF7IHHS72o7IddO
LGfUOXmwOZ+Hvj7sf3eBYAcoJZQ6fKSoYGbFePzFD5AN+uKgfjfvuxcVHhUtmFSK
tmj9TN/GNZh5dYOmUvr1YRl6/nooLyAxZ4gd8ViZgvrvjSlJ8dfkPIEubXd9nmlT
ro7y5wvi+khfjK3EeSJ4qV0tklS2TeV7fUZwzQMAOUw0MGPllo0A0autmCANp93Q
5mYPqwURNRwypjGHmwzaQ1caZzs6uYOyjV9D/lqT8rWMBXqCYFEXaxIdQVyHPPnS
w2Yb2xujsYbCIUv4A5WUCdBcdrIqWHZ/jP5vylr3fO8DUCaMQdpS/MZ3KBoxQwUn
ABvO4R8JXbN8EG/B67u1E+FSd3NjlzJlMT3C0C0nrWZmGE7TH779ObnmGMcquR+T
kcABg1SvzgKIJek3Cs+tKjrGSdYjS+FfMNxr7wXiB3iTlaBFk+xWGiJBSLl6NhS7
CaEOJwtT2nUcq3LMsoisY49CQ9p7b5iz65zLtp8zOrNqyUhK4/ioRQEMZoz90Kbg
coavrJVtSDf0F/BeY6xGFCpP42fFP4IYIJRnjYFiXEcL8Up31L3NkIYgfUVk15Ux
eHlcI0ZHpuKfU6BmRoYmSiOXucCrXkR9YbZI7OEKmVjtyhr1sS18QcBMyY7GYP7r
8NZ81pdmPTPec4J58CSf1cEoPV4XScxnjlhCqU0rXRLz5wF1dTk/XgIwt4KD9OI/
hDmuiR7diYBYJ9eFUqefuJIJNnd88exaMfQ1jC9NHFRWegMhD1CohIngD/8S15x9
xshmFciNEdQO0laPs+/3QYG5kqB7rc4dDl8etmrUuUKqWc3CWxZfAE2jh5GyUysu
6a/tPvbvbNo0lD1yU0WgmtlSuQL6Vt2j6y2aZ83fsS3wnQAufzxfvCfavKJHqBAI
HmxlGrn/+WO+GVW0d/TpXJNL3rP1nAqO4JSMK3vCnl30CKAlMGUFa1JaSWUNG94Z
wThwl5NzZ+WL8WqShdTlOfWvn4nIhJrC2JoZwzmjHHb9sQHv1m/vbKRH+cSnlwBR
sbZAEnB87j55XzXHWgKe4vcvKH7YRUtxHvRfXOCYUcXsAjjByrBojpiOUGV7xi8g
xLfAspNE5Fq+N2oQxz5U3FFf/shua9QF57nws4PWGLj5KapsiX+JND97Z60uOvKE
cTGvGR3N5pv642+HZdLXWGBjupit5+HRcz/deZbU4RRsJJZB7tne+XZFMf+0EzC3
X1xnaEowW8FlLEAqHHUJzQmEqyhiROqczaEjROBSNCNLqNfxITM4axVK1iCP4flM
2FoeZTq/eOQ/JJrPyQUK/2S8697jC7cxr0CvbHkA+LflAws6h/wIyUSyqhpPBhmg
B+fJwAGY2mtXvuJ5nOInpBa/Z1hmrLKcIQh7Q6XVB1ZgFsi9nk+TH51g2S03rXQX
CHZx9zoK048FUVGxPcEJ/JjKNdVz4LFEcdYDfsnmPYjQWnx57Quit/7I9k40Oj96
20SfMxmq60pCKFw4k1KJ+5qRX5NKfdUqC1aMQjuCHimRzewJ32y4vkeL/XA9t7zE
D83wOTCHKlw/W4Xe5eReNrudIL+DEaVlsSC/KhrLDz/hhTFF2kMZ35JyBe4Tw3h0
to1tsD/LTNKcCxstOwUaD+oKqlwDH9j1AjjrNNSLjxvxqhAhfFxVLF74ubEE8G0h
/Vi7Wm5suyMHeulFQX9hQlbF/lYQ3/Qtar1G7GLSFXCFs93MgSce3pSh3lY6VulA
ebMYK1a15AWgNpatymwZrCX4Hv2b8sKRQTpdKq2K0nh+XlhLnatn+lvIYa1l/Dkt
7fAUdDzfMy8RZkvH6xabFJLfPsmo2vgqFPYny/yV/4X1dtq70v2iAB7aNZCHfBTX
sYtvzxtL92cqxQlhj+SmRBUadR5iaDl4SIo6FyrOYn+ov/Bo+gTHlrku8iIiNGjA
BeCMUm/vCODkAO8H7GYqutQE+TTMOjOelGKTAnX7GatkJeQb5WSKIrFlW0OCKPGo
`protect end_protected