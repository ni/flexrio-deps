`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11328 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0gQgIG1mJzulW1XOK5NnZR8
C8XqDUtXW7uOWTnSVqbIbjyY3rtHDDuigL2b3nWaHShLOYCemKMIr1EALuwYJmXg
so+01xhJ5ZIEzMmuQwiOpkmAsHwM7BzVj+kM/JNDDwQOabRRSy+OLfNGpyYkuLIx
bDldEQ2tmkFyDFB9kXT9oy2+NvJhqMPL9/j0L2UrR9atze6SIgefTF6sltQO43aF
sdhSCwfNUkOR9H6/txrRiN87nomjLIVWJ2L+gLOHPMeR/HAGq9n1cEel6BNOEale
hNOJcyx/WvGlO9Trd+vMP4ztmZi7dpiXiLO6RIooe/gVqCXjl5OAogZpUFAi/FQS
ihdjAeTtGf30LffUdJQqYjydEM3WW44i2GuXd6Cc/MioD1v5ewARNjEwa4axiJpc
4eUZHk7sG371qrORlBTYK5EPM5IkbsbREb1MhkT3NPmbCEKxrDjw83QGdZuLxZEH
OQPn9EXL9O6JrLgpfia1ZNluoXXAl/3MKddedUWd2FYSRdTHylGUhe/ZLY+ulGba
DObbVFULSDM3K3uW8KqfXLglcuQKNNKuk/OeQ+YyhGvpPPtM4mYb/kDEgwHuKEJt
EVu3JGouSFOU0LJqA/88lFA8ZGSH2Uc6ajM0hpMxKYCcWRxwkoCE0CgNj8e31p/r
ZJHXILqgB1qfJX2eT42SHVcYOVHGtL+HFToL4TbeDxTKR7pjkdZHoavAnVY8FyuC
dxIikNnfjYgXIrPEfCCDVLPktI7MbKUVVcPaxVYLPrqIzGdhlGOzmRLiVfzPmfKf
PDoYNwZMOnN57fwGilHuSZfN0gbOIhOy1b+DyVzYbsX0kjbB0xkQL0D/Ff58O4Fd
JEMQ6Zg3yXNujKid5qQscbMGQgsi7TlUS9GAEByg2oNCo8w/3Icus5iJD5Fl1Lhg
BjXq07PMIgG1kRhLr99+JgIrNBLoAFIH0LFFW3jBDzvDimdOwOVD1diK9eFq2A77
W5FdbGck2CP5selfO/M4wn380fZXM/6p8oYfgvxfWimMO7xTiwvy/xZb2GjdfArr
CZTzKK8mZAq9qSD6CysnfEgBsJeqmPsZglK4/Rxsup/oHpcMD8Oy8cPUsU+Kocv0
yPf5MNUg/42lFI+iteDr+CFZqXapNBstjxRLYFY5ouQLsiIlY62AJACfOxI9QlA3
K8D2QBGen0lU1HwfoIVT0gMONSX0D3dMOm4oNKsZNzZPMtXv/IcuKgQQVAR52Vph
0LDsZ2OQ6tQ+2pgsKtTF0e/O0JeKwXMtiVAKeQCmD7nGYDOm1a1kJePocLHjC0mE
rkUgnhFjpO0v07iISes0/25jvfegLAwlAieXi7w+8icXUNBD6n40+pdmr+74d0OX
ibKvJPLDacCQeOMwB9QfWHbq8CSqNX1hU4Okl123hZ5lcPadH5Yo0URZoHAFZyPJ
nLdK9YmVwY+6moum8QUHx71xK06+T1+feWgQW1w9Wy1OOtD87AANuxW69MoQhsJu
nrg9WSBNXKLtPi3bdvM9bgV5xM13JmPduu3JPtrSvJO9kIamUnOrv8FhjmQHbCWJ
YTo8cLyzuXvUFG95giYalPWqjvVPl4Q1j7QnAT8b41GCyMNcZ6FzcrWt//mVLScx
AjsyynCF7Z1o/jb7nPefpXuzxaMSQ1ocslV5SsFH9PJVi78FqBtoULHcTT9tdFZk
8sRF5RHjBVnGH8uB8MK6S6YPwAYCUK5ucCK3jXaYY1mTtY1aioBwewFBsXW8sFLo
mM6AAsQgV84DmHWjo85bQhenvoUgHywyrG161FOmm5ei2R9xvZ8g+7anY2+Yx0D2
uND8xEu37zWBncA6KUjO90NWEZ7wgOkq4zNqIbwEOhDsQu3rYqq5JwcLRZ+WemU7
sPAvPPE8SKsVghtJrjilPDkqushLz/29rTcnKN0vP/PmgDpe4l4QtqF3J6feK+ab
JwtqjXdYhWlMubypCnWpoWLcVl4i7PrVFJ3QRVPxuZ+t9MI2EogaSh5Ecwt+YSYi
iD8an6mq8VV6Smhsi+asMXKoSnbcYq93luzBUsKbdmKbLx73vARYz5Qd76iddueq
RCGQagTwWtLK/XVWLOH/j6SwvYSX2If77MrwKkE1U6+QTLB5bspz/ceve2F5ujBy
QuRk28X287QbOgr+c9UAGrzp9EGHnD0oEC1L16bGun7S2iHg/5D3mzcI1KmqSoZC
Bk1URPXX2HRgMvEjN+JSwp+tHk6D7wMvINlq29hWN+tyENxeylecxZ1OKwgXQa3b
yrWE19ycBeWTVVO3HT/JeWmyun1n0W7lKA2SXIJ9m0ptZYmDQIz07Dfdvxv7gs+6
6x71uSBtal0usvQX6XahZhFlaw5Zi4JoZsjPx4OTBXDT5vdY+lfnHx0Lqekw89ZT
NlVUGdY4Hxy6MvTl9ZPPSmm56496kYwJgWD6eQbR6cjGxQze2Ea+evTTBq3JtqXr
EKhHwLYW8B1j/BTmgAhTtJ2aGENmblxDu9mFDDf9QV/9RjVvUGGl0afF6tGghAoi
a+b5dOu9qFgSaWht9GwsMb9VutqoxJQKHI/wQUyl1s0DRSoldoFokUvbglEmutTe
mdX4Nj1TQuHGg1qB0YWG1UrPD2yIUjPL3OG8zMTmY9+nzd5VehUK42wrOfEkmppx
88C2p2tw5asjVaRjIOB5+GaoqJ3JlzGwm3362RNtQzoe0eqQanvzRWSbT3ODAPIL
YaAJwocH5rAlh/GZY8C+x0z9ZIFpA1aGvoaGwO6pn3e1s6j+gkPx7NLHgWDL8oi0
i0jVsWOZcAMVpo6LnEJqMAns8mZehjP8IK2cBMx8E6Ndu43XEbpmUAr9ftilrWSm
Put/hlp8+E5ayTjCFUVpFiwIYYgH+S7nWNEE9K16CK5gdqZ3aguPT0F8cGcf+QN8
W3Tn7qVmtVzjj4k/RIi0+EE4Hmt+eEdmPoz2I+W2b2U1N2cJhOJsS0Bh/x6b82t9
8W3pfvdWCoOoDAjRfWIy9b81FDqZTWPPk99v7RY3ZBd8IDmOsr6pKr7TR8DypkaM
/B8aDMnYsaBAtqCxj+xzibUC0Mhs5iBvalxJ8fR5jOrY370BYUmJlE61oAq1xv27
Y1k/kVU66dKFlaBjtq9bWYkIfV5F+HwPzwUq4yLZPNE1KfbdYaemqdDLtuP7Lbuf
Y+MIjdE3AF11wcFYsb5XJVs3pwqQY6226fvgZRAHwanzCkEdXzlWIjJ1oZxm3BP4
Q71jQ660pcW5gSH9ggDaVTN35KKaewtCkHMOOENgMBcLMnDNoFQC4RFftivlz6/6
Mx3GwDXqf1GhO1WvLT8alh0yT5aLcBg0XT6NT254JOOmXUgXKM2QNlWbMeM/Dhd6
WI3PMXTEbGpQ5fusVMEV5Eq+6+u4ilpyACeqNDljbvLTvBwboE40l74egjw6YA7g
O84Cd+pT9eRZkXHT4E/k93IBqohF+Z/QHOIT1RtfchI7OtCYaQ2BxJJFBceA0/BF
Sp7vH5EWidwQGAEk59KA98X9hzZFpGD+3quQM1j4Dk8M5S0sc0EwD39DoU1wteo9
KkKM/glts2Z2RCXSFsAEs+92TON8A28pAAwoSKRw7H+MB4FGcqvMH5Vu588R/Lyr
HbDj0nL880qEPkvfBSXwi/DVgI7eknWe03AaIcog19HgqHXmrWDAFiclRZDjxzDZ
7xsnPeZdNmhZ40PNkUDVMocVkCm4Aigf2FSReM8z+d4VtTeLKZpaU3s9VOhFZjDF
Eu4iM2TpehE2KX7lvAbZ60XeFe3pJk3iGnZ5mVbhIMLIcX21AAihMqwVf1jhIaJH
SlZAE9JdMiJ7MWs25Bu8N+p0rUxPY0nvOZxw3H876TQbrnbMUK2A4IYuawEwsPaU
kWZDz21fJy8eYIXxeBxByge9dRVpkNFAaAoBbqHjWZWDafO0U1vPcXK/HTtQSwVs
uLisO7aKSyoAYWouJPrA9Auv/bBAKSykr+yKUkll1OO+1+e50WxmfL3ToREC6gj2
fgnmGRcTdsvNbPI/sGYWTwXPmpEWFANiTd9EFEFWBnX6iCxHREfJCxXU+ID1XHdf
/PCJ2DVP/fBdzf/9ZJefEDy/17NJ3ZlkpNA/YwHfobpky19fNF85MBl1TcBJk+zg
ZgNau+qyJFdf7KvJMPZ54aQtmdSwmaIejhrccFLsnfmmoKVlKO+g+tRi+sCMCspn
xinHIxES4D2z58+7FNbK43Tf+c1YWJrPYZuBD1q/0wsutMdGDJNa5j+NK41TKiTv
RgxNPwO+Y4UEiXLhl3QzJMMCdKMAPNzVydSgSJUSCfn89XxO9HYvbmQxbTc2lEew
EwUk3csJX9VbPYpeCfALK5QMzDtrFQE8JZglajedaBLAzi5xQqUoRDdbPJyhZJbK
qUU/DXp6zNR77b1JKj/vxIgIbjQOxwH2X4+vevVdHCOSHonYjfCztKLRVQJKgse7
Vxk0+cod7sbKnt2KaWtnhYaZBD6VH6vEuBbYtXqEARU+Z7kTEgsY1lpTCU910hro
ESbkGKwOOADWFDyk/JWfMAx3B0j7SlMGaOBchUK6Dv4PMZJhLsXoq+7LC04tjq7f
JwvhtramFf/QNEn0vkolotvrc4Ex34C9wr+eyq0JF5DqSQziB6tSYzizpPcUMV+F
EB1M4LmTo7y1ufep/BZGfIj9ruiSIQlH2W5JL9nGj7cFnujdWmoLpSIwZSBtFSPi
PaTHz+w7g8O8YwHrsqlvuIih3rk54FiS+o+T6Rz/GD2OYX1ZUG9UbgCnwhqxfiFi
3n+OYX917WXzFzofwFhn76t5r6/JX0oTrgtOytnJfXSDqPdFk6Ptfa0ZReAOh4S2
E543KjpskTTv/BBR4V2vop+rzoAXk7XzP/7RPXjfBfj6sTr174yIIP9KwpoomIhr
8qDXGiRx0gMIppecsB2zKBAZLaTmuu5/UJ7+oSGhQV/FCF9keuzgrR0BQRDDt6g6
dU/EAxT1xbBJmu2uJwHGI8/pP0Q/dXmdjaTDFbLDPC3wAd4qHZLNu6kvMUoPicOU
4orBSOrIJ6uuXd/Qwzl+atTxpxRdo8oXLBuLYIXNfdPwAz5ryuxB7o3+DZtyZ3iM
3qkmRIpuLBrARfZlZazeaVqclbsAoanTs7qfoV2vx/zKKnpj2HtWAAsLTb6yKr2x
LF9kRCcq8JNM8wVvMJp5VNKOssUq6344aQKfihH0tcuCjNpXJFRS3UJOtUzTHLM9
n1v+3+3BupHTF2s5M0VQd5ebUirEWpcboB8voH+D8ZQv5UV0tPaxOYMV6J5iBHdo
oV521G6zprrSydsrn+hvm1wz0NpC6PzSdcRYI63lKMhdm64BQM+Ilj9MC8jeAQ+q
RUuDVWAnIdcXysBbPfvLeTX2DhNy1U1Ky05ut+v35oIlagl2b/vPJcyCL7UCYjg3
sFafJM52BXvO2QYNF91OYs3uONyXVMT5McpB2TwkMNvpMm2vtOam+Em5XZ+WCS3p
zn577ov8UJo/M03wJJe1pSjUUUe5UDZTUDTYMhlrPgnamnM6/40Z7GkZLfUMH71P
hmjnk+g7viu7uOiKMA06nY8UwlooNIMTJwZjekH7n4cEXUB2kMbSmBp03BIQt6hB
sSqIzB2b4FLqzdvDX4IWFtCPUjiCNMeNgcKcAtdqzU63hm4gzFsVqWVQP+LVrllK
6ImVGEfuUTZXAFFniscgUiddBMVEq9uCOeHLx+GBek8QaY3CsHnvcRX34oBflavA
CQCkF4WJPUjdJUN2DFr7kptYu59+S9zrGxf2mTk6FqZe+pQVLM+NpTpEUtLi98ZM
YPyXXAx6b7mngl4S/0V/GonzszQ9KGpzZVWzWw/SxH+ttvywSnK/eJkH/GIZ+817
k5fBDO/6cC8KBN3odxNxFIRteAYKq08oeCuHWTDtAe4IFa/XZSr4jMNqmZ/tYb4e
Xrvwou4DEJwdAntLoaQivdWB+W8AX9hdyGvAfqF3Fme+bq5BAjd8NZIhIwyCx7nN
x3CV0yODgDhd862bX+JbWmIc72w2yFPdpCIsiM6bmDnblmSku4kAtNehuL1IRJUv
OO9M3zxhnjrBVVIgZTCM81kEqZyMVgZ/P3nfu55xWwspkd1vTl4nW8EsvTgk5/C6
hr8MYannxTy6Xm3KniQ+NvL4obxzSRZuA6cZhZB/AxIFBt80yDxkERnWLRU7Wg7K
FoTAK3vv0awmFiQR+G4d33rrU59fQhp+MPBEV43QsTafhUfJmHGh4ELSv+zuriLc
9VNVNUGwiEHnB4nQEWbzOoSYAl3x+Tsuc8/5Kbl/tdqVDYAc4PIi3Hch7NHTO9RA
CT+GgtTd7TW70NhCd70FtyPdvG1S59xF5vzSnh2C4k+vYiPD+LmZ6A6pJdwaaoaI
seH+PLqfQF63W2sVrfOi4IZXIsrevtmEmQFHr2qO1gkHplPrkYJx5EF/S6NMlioD
MkGICqKNmBuJt69kbg0XU8junRvQQwqVW1GJ5s6QHECKgwc0jYQasyxqNooEb0SZ
gQv4te9OruyOu/66Tx/ymGfbISIHkmihL+T/hWP+71IXq4Tsa3SJFKesHkJWdJxc
mJROq2IP8wSntTLzGUI/ZIgX/ozk0EWQNC95S2fsu8aYro00B+zNNcfxQgvKwTU8
g1/uQQDEdHc1qTlTzmvvG7EXaTLNh7BWUp3bojoPROPQwzNU9Wsxopk0z3up4y8a
rAmEcXv9FkixunVYmTmvazZDVxpP5T5uCJ6TrteYxTh3LHCmbmGkR7bA4suUU2ci
WyHKzR0qAyLKGN0/keEGhB8RCngXL2IB4H1xCwEo2WFvGIPkzqzu0MCeq7kvpheD
i3Xgdms7mKrLWc9BHon08i73ck7a34ocyOb9DNUAB3cfonJUMFiRuGxENrJPwvAf
KobNbNGAcv9Pl/KA5NIjZc+DoEDp9tw2V78H8iNPth2bUTlveyKVHex6gmAvj54J
1Q1k4Duc9K+64PP6wqxZqn10kMHbh565Jr2Wa0xnH2B06MWCFHjdfoQAanqINNI1
xO9jKtaNY8Pi5E7sdHLEW25GrIB5V+6M9APC+D5bDh3myRtYMc8NZGvx547tPcil
rxa5TFR0PEiMLJ/mRxhEsGligZHecF+puzw11hEI4HoKO65VIxI+M3zY9IUcDm3G
YmCYJrAJ/YXWWdSAhcjYWLID/nZY0q3QjXpbqZlE4tTF/6dWaDwc8Th/W8tHbY3W
U6dTssbIrwBy6PqOGJI26hlu6tspA+GyzSRwyZRbGSFHI+TlZCm1rjOabWb8jtzx
6RCpgS+3VDkIwDV7zvX94TMNOxp6qiFWYpohuwKoEybTFAW7QnbL4R4wZ1huN6F1
I/jueHN2NRx4yc9A2w+OJF9ckDcvlo6qJ2gnkweP8pf+DKRdpfu7+ZLCDCdZoYWc
IZU5EO5Nf4dSZTXrR8D2zTs/MPrDWm2ZCh6nS7CYcVnqESn478qyd6e0zBRQZS6P
sssmwkW1eHqeQRNLmFReyJdebgNbljaphZPBEnzm18qKvApJ/SloEHYCn91UfKos
SIdaJhvKT+rCXvcEDee5I3xycDbTlLRe80LnauBjTavuMdWnIvFG4RwobACxxMCU
V2MoqXc8zRquRAenp8x7oAiuOIbv4jxdwBzad9PeAfBvwLGEnBmJLKwm9KyTV6IC
TaUoZU//UgCO2lsUjtakFy22n5OyBDOV1jAllr25PsqzTkDVizvP9QoTzPbUGNjV
SDMDslwl+39MfSU9doTBgOevQzFqhkni4TEz1UJdpJqDfxUUnRnRj31494oy4A6S
V4eh6CkM1I+YUFVlRf12tFN2Y5TBJ1WtkmNw5M3DcUs1NHMEBH6jwvig5OCaLbJz
7mCuTEWF46I3Yu9LSJ/jzXGcwtaPDg01Xsw2ThkVs3eygiB8uoTfNW183doXiYR1
pDp1uw44NiHJv3MxeCYflSA8Y8A2uhJ6V9q4bDQXqWLC0Akp7kW+FgB72FjnkCBd
NYZNNTuKgm7A4UcW2e47PliHfNjnJAkkbiHOiPgZfws0l+XCEjBYGx5oxbfHTxax
jfXCAtj1mzJ7foVGcp4NPVEReRnXyCFTMsw9vAtHyvrTD1GVl+ZWJdJGxEhBOFM7
a8wwj0uz+P2Kcji4ggu0dMDZTKzWH7wCBzIGcyYjs6rsP3z+t8xrV5m0k+HxML9R
n9mu/4S1Q2UIm/7FNExg5oJ7nC9xp+3Jo8WJkuH7jddYcs9bUTotYrGRqxUaXPyU
4uZWlz8fdi0bJn7PPkvDL2ekofwguQsFEl+40F0qvy1+697BOYVhpKxyoZbLMC//
j/8HPsXFQtvBZko3QDnlwJOrPDBDAYeWNLyBCIo8x9T6bItkOyff4bznZcO44VmY
mrk7tWfZz6ZP60eWE7NevtYlxKIsFfpqXSV14SiFldENrMvmHs8rm0XnX75+lObD
FgHIfVHLJ+OoSX0sgYyrHqBeALdQ9VEiIvE5oFscDrd77OZgXBq9GYhA0y4TYn8s
GkOHSHuxgS2T5nRvhAuvj4LSmNi2X0bGex1r+1CaovF36dV7tFoH8duVw/n9ANyN
rRn3jrC3dicx2bWxeEqQfywSqoWE+qH7ucDvXvMqun50F0qCG5G1SB3TCjnW64UV
QLfvH9wDKjhGMuj9q28CNISQdaw8qbkSMpBcrDoVw6/1rejM3OtuFe7w+pt16p+q
Iap6JG2YQekypSuHwwv/aUI9EJNBGxfe0aXYLsY1OtFiwCP3aO3qQt0DrQoPCbMq
ru4je6IEzaQzmG8AIXtzY93tOwloZSltcpwSyzbCvsqQrncFiCLxa+CO9Z8lQYgV
3RtKXWus1YtKHwMbLHK5Rr97cOifBXRKy90Xjp60yAqCF3LoJ7fjxuEuOrXJ4hdb
JSGgHQWyoj9RMG5r10JXPNiMYoabVvMsklHubqZ3jDhXVFpdILfLFMgMlLoUvwae
BNgFtubepBAA/tPC1BRjNK1CL+ZAcATHmwqQSsyNtorGg3gLLyzzj98pa9RQOOFS
46cz5riDhiuw9o8egXTmWmsnC0qzWZ/a/XC1XYxLxB0rcQKl57TaOyJQEx1x/bB1
vfR52R4c3PHglQAh/h4TgFcHqgpE8Ji8UsZ/DBNEapLbrm7CIilCGVUcLh/QFyox
z8vwBE5MpOkh8rwRhqF2WsvhR2S0duj1Foa1CeCzBzg9wfhvLjAn0QzTL1EtKP3W
9aoYGwpyDbd5llZrNzAgxDetpg2MRzMGjIJspekmpxhUoK5wRQpZRyddbzjQUVMu
QZS7M+Y/mNtMQTScdDC65q5kSJqpNF9k1T7PJUB928UrRxRmsEZ5bctNR+eviZjM
WvpShXJMCEyY6eOqaB3kyLHHsUAtw1I/4U+0A/LRDkL332Ptn+LrcA/9chCV7/7T
72e77PKEYGfNBQZtH20SyRtjYNpjncrMPtlxLGxsDcvPIu1V1zKXOxYDkSpqPUuC
/AVDAFBfYSsSgHG2r33OPAUcFgUT3ry9ayAw7EtdBy9dcRgQzG04H4Qp7Y7PNyIh
Q4ioLBvuDc2D8P6TVbcOBySjVt62iUa2Sxp+7ken/uIHMbgkReAUrKHnlogIcqHH
sMTH7DVDPTp/CszCQnMKJm95H1g3Q/yg7AlyyMF6W9LVG+yottITC6V7R2cBgwsH
k34D6uW3LkstNaUUHP4T6Q/8qVVqoAmQHxLrLNbOw+8DXnzvKaTYP0IuZjcs7Dby
OyGsH5gBiashnHNbbKL+0CiJW0HduKzS8KwXbAF7ynScSeBRrh0xrPf1KhlXI+VI
gQ3F6A78WFMZpTqMPmmDPVsL/OQ9HrsdTlyrhsua6gjGbyvMzgxgR464T/9p7cVK
Yca6/O6dBMYC0+cy5zZ/moRxge1T0D23sstQ+uT3BMogOgqvAnNEmiL9d7L/7irx
jaQQCIfp5dmkCfJaIC+LsFUhxbbP0PTIXXhrGxHCzad4sX+aasSPsyGmUX5vD24S
Hil5guRny40kul/Dfk+6MwrSNSoED9FNn3Wv1+TnszbVfIVptBE94WKT58UKu/jn
o3DWyTDhS+wXggpPHnNdF77KzN24nI63u2aqQo9kDL3YNpJUjeFYrYHgbCpag111
JXwqJOtQuPT8X0FqVHoI4UdqNX4VoS4BTNFyfZjtkAx+++orXNUYHunPVmfgQQuG
PgVbG2KncZsOc7f8a8phK89LR+hqQzCLYEUMrvw4zZXaTyYjoul0c2kVRucGyC0K
u0v+50281/gzKqNBvyKbd8pY6knztFR/FyHHZRk1rcLgKN8rhYo9MQ8YIIDRyYcs
2W8Yjkknw2cveYkdiLNeGcMy4A8l6QUisSHjjAr3B+lZEeRoXIjGOihPp0q2B9/p
2eHL6kZCgRhA6El3V1EONydeMnu2jI/29BEtFbcLRdPu4r0Ck7QH18i6nGuSjnMQ
/uh2cdTunXoPr86faCJcRhlErlla0boO1btai2rYmXYQFmIq7tw6nAxhgFy6rHm5
D7Gk/OMJhp8xeQ8r2u+0FQ0DudgZYEBMe7hb/fPg7IyGhqDMnVAgvf1subKPbBHU
HrkSTABIHwqo544Er37RavAKTBKl2Ji03DaUYjhtpBvjOnudwNVdGz/1nBiRaU/Q
FtaXC9xBmeGKRp6GVOETeqVe4hF21l6DL0RToS0tf4ZySyFSvnhJZQiLDyZ29iDD
WjK7RsrPB3k5tSKJF5AVT0dDKTjHhXLNdspe77ghjLPChqTey7MX4oiyihMP25ya
C+b/COmcigDYEa5zGij8MAKuKH/FVfwDeOGG+a21yo4lr985oJ57LkX6uV1Kn0Cz
f4i924kb09smTJ1Cml7WFiGN4llb2EGOBCFm4cXQrXebUcIVqvNmahElQJf7o7UW
3WX/Kg7CUaetwCp4CacC4PwOLTnW7dOdwVD8xvMum+vhH70zvYyipoiFH5uiQswh
DdEeZmHrVvFf0uqDEQgmXFkza5+kBDiimsN0+r4uPUJUgI3mogsehfqTn1g1R8wo
r0FKIHgQItzU5wOOmdPn3cR1WH7FzLaiTJ+KR+tlUvF2bUb9Tiqfy2RsOc4V9rUY
4uTIAmlE8dFHB/CaYrBftHS8esaYTRikzm+0hZCguxJEH4Crgj6BKf/oyJs5hQLT
xfO8fffa+r8zMMXmrGDwVcah+r4/1kOjK3CAKSpoBzN9r7DzeH/7WRbAHDmRF5Ty
VqulRYUS53KyonQVfbgRiOtmntk1LipEon9YhP1PsVhsH7vTYP8/O5NdUF0OWhnN
RhHml40/igEVpUZvR1H9mqHi5d5MrYm9e49C8bYyrkTimmU+3VMZWTDisrCthf+w
JUFaSJGKi+duO1WNAD7GGl8r5w/XprajHk4ilWlfVpz4T6e33QS4tEENZenuo0iV
ySNtKGB99bAvaucpz0qnOBNxDSC1SFw8A6fd7GeBYk3PXqoQFEoZye2huurq5dOL
CyHONQY1T5GUxYZjF3dFvRE7s+2x9Jl4SN7ym48TaQdEjBwf1PZai8u7P9MvmvVh
p1tAQWAxXQyxaCygvrooxQ4wcvi6KQyapfBLTIxfxbaGI/Go2F+VR9mRa7R+Sfo2
8zgFsfdeZnnYmcnmpRZ7cuTay1jArxTn76iOUsGORokKL0X6jWSFZ/NzhudXtX/i
lmi1L1MnSj05vcf+Kv+CmyExIom/obrWaYcU3vzCEpC94txlkZoW0LaDGIIQTOXm
o0nDxprNZb9xOVjPi3nd0Iioh7Mx7BMzLG2itDTpqgmPT7ChVi0O9irnEvVN29Oa
2Vc4loPyWwI9uWmKhwJ9nTQX9/gonjzWJyMqm/Kx//8GrTH/UOLETGHMolAPwa/u
JlIBK+9xPg+eqSunxnDR+Fc/tHDiEd4MGpxW6y1PKCHZ1pLoDv2PwF0xa5wTOQEC
dKLeQifFZRqRijXOgq2QRWDntZo2D2pGGcot0dI/5T07eUSWA6KO687uzOFKtUz1
mr1A+EtoxJXtqUSNiDuqTlRiFT2ZTAiRIgVVd75gmgno+BXArBu5cQxkGRNHWBGJ
X/+YMhiIji1yuqvbBN4Rb+07v06mv95fdDmP3UcVvpDQT1gwa0vCz8F9aQyZR8eJ
42Jv8U/nm6zAYeqNxzbP/9M2BzFnQ+meyuiy48REWNhkw7Zx9jC996EeOVAFrYsf
D+SJEx4kDGReYZXOqh8wI37xCxLL1eilK+zhj4pPNi5TWmq7B22hwaJ9pTfLFgMi
XA7bfgKfB/pWxh0g8NCPyIwjbuCgZkHqoDxvlgbjOL0rkBmsAPdNpGMFQNt2CoHo
ZZzREn/LxxKpgUo0d7UjpAruWyBGx1dym9UXttMwkMTIMZKAW9hR16XW+kyjXkM7
TxvVSkVRLYumS/LbtLtsfFvVlO8n00AAgiP8NFmBGqDWfL//S+5ksFLtSX/ZQJyg
Amlezwj3ZTBwNt+YHD1/1gAmSLPgBF2RXtTIiCV7gJFx6hq0B+wHJyFVoX/xOYwS
f1shQRpsLwlyWT3XYGI5eP09BSy9fwSO2b/RWD4d6qm9B8nfIMTB/Jh8AdwJ6EW6
dqpI6bh9GC2qpc1p0Vjw1QYCNDpQEA/mDBUQNHubbPuDpgwtd0rkfiA6Vi6vbcyA
oJ68IWXcNeeborrcz01shH7XsA3Ee+jXcNuRJ7gZOkDZPSm5N8l4rrB8t7Tsb9Yt
E75+tXDCgXcGFXneNCfu7n28NoQUfissQPRrY0FgvBY6brY9kx0drrZn5kl6hLlx
iAtSw1mNRilKxmZISdlWlUM6hs+gR2Y19jxB6WYhvlfK5ROa3Xc6Ovzsc8D0xGQQ
Zglpgp13f2L6RhK8dm+F8zTWZbjzkAs13VxX87pwDQA7AJ3WGXt+93ZPKvxBrKoJ
eC/AON7EkxOR+Svll9pmFk3TN+JjbJ6uVQdHg+/e595DNWhxwWUlBQUVeBaD+CAc
HJ/MqXHtDQ9rbM9YWZ4xDUbCT+R4xWt5QYyW+sJGFNiNdcmRfLDBMu9u4oLMDCf9
4qLDjjoYYtNZWz9RsDDRGbuOD1YIIniRQj6QhriCeIH9qA2emYQAzCLOil8wV+dv
SQ5yEc6rPZOZaKh3kbaos3+NN+z60iJop6HN/G6DtDoyhkMps3OG49n5FlQBmXeF
AzkM5Hs1+aYoMJqtZ5wgPpwOR6dNIpyIHgOHSneG0kzPQOQj5ZFjXdeChMGicEfS
nP4nFjIbzRsQo5qgDoyjk4gyzZDqNR2fP3+sEa5kWK44e+RwHCZQ9x3Q06gw1iV6
n0tfyXtMK9lS+zBGHCqHv3LBqeZqU/qOkosO0oktbi9ecvFYXiMW1oYOK6NJvxSo
zb0jhRmPj0Hydid4gBkYtoPjA4dl9UTSF34LtAxLuL5hMCXacITaUT+HsD8iezY4
xA0TFHI3w9rv2L3ra4HB4cLk2owq7MAdBevMbwwxNhYOne2+e9XjRw0AQsDeL5S0
RzxY8feJ6LS8WLK32j1SB0jpXAvVAevHnLpBqzpr5F8FSodie8DcUM439ydxtRrx
YRedGpHi0YKQEu0K4GUASllfaDsiGKVPWWuzJyFGYVYX0GeljfzPG/0rwyjBMR6z
NRTV8nSFYbGCljc765rqL9HMppZcAgzspYSDd0+Q12ev/dhkhz1J+PqSBdlUN0+k
vdpeLVpz+YhyMwxm9IbnJfjL5p2mCZFgOXtotwESjyu9RAQCl72Kr4UzizwfRSnP
4r2ufyBalFA1f9CyAH9ojAB6+kyHxJgaHxnybV0lGSYNZRIh4GwPw+4LWbW13szP
DEDC6lT/fEb3+qa707+Knnxb5C5ruso+CTm3a5+OWw0lumLXjvm+BWf4hn90CLj2
qmFVeG60/lKkI3YZbBkBplMkSGKR2uK6I/dDNdv6tq+1dTwIuR5vWnRvfR+CSwsE
OJqSxPcg9ij6qcThJx6lY2wPvUTs9yoNCx+ho6SUHf8y/xSyVP96a7f8nC/r14sp
g1WmNtn9YFQfLcp++gnQKUwLJPCIKqknmSSMjZMv10DzT86+/VdZM1PbSlzPcZ3g
R4Mc7BNsjIY6eOZz3mPLHls7gzOLomSFVFP2ZMAUskD11ATpNY3gr/i8vKvo7mZp
x34TIoYbjQ4DmFtASVtJyT463c+0yeOsxMqk2eqgNu34uh9avp+pLQtU/WYG01el
WvEQ11QooXD3apOxttgrfeJ2ONgSgVPqfRGBkLLlrkjzUJADeRguJpCAWQMBjvGu
ce6Ho563v5X/KYo4AenydBlI6Uc9G7puKnkeuXSK1YtK1cwgdoEYTEKgi3POoS9v
C+7hF8kbtO5pQf+ykbmXvIsITlXWIMaGFW+WAq7xRnnmJp/YL6r37gloumZ4AnRg
EA94QxzmRG63aO+5OrxnMhteVaL6omklv9l5SHdS12ADodL17HnYWUUNqUL8R0VS
s8EO5vwWfY+bF8j4YYYf/8Wg0dPQoJxx0h5E2oxCAjL2xdrzlp4vuUFqMR6vIgmM
WV4elcxa+L+CRpIO/LMo/dTKbr9/PmY86IFrep+Oj72uR+CqCh0THeOYa+RCgmZe
OSfSqhsX9jLMWBGcZRE5Y7pe1a0PorQTY+/m7NQZ1l9r9SSlGQ/+fMfz0tqOUCIo
8E32b2L37eMdFRDU0ojn7K6pGcXtWSBPzthypZrn3ihtz9PfSKnp+I5RRnnJ7L8A
/euCL7qTgDGRuEHms/IYEhPyFUaDd3TqkfQ1echP9dhnea9GKzre+GVd7ErthYxy
7w4uydUOAnzbrmkGWHUpHWp0AM+8kUpa9Z2dZqchiDZYf4AYR6IF3YayjctlEdXb
QdzWeBuyndDo5iqB1tke6pb2MAH5uib8G6+bZuQa6kDZg7O9sz/LZULZFl8jLqXh
t3NuN+h/WdduzS4THKvHMRERlQRPsCilwknXg/szrdxhFsPe9ohTwGXrcaxj9hCZ
g0NBGHGwZypiHzWiSUUcBwDKpgu8035cSrduIIsHIzBtMQPVyeyOWBfg1EJqKlto
TElbfPlUoL4ZB6rsoXfRiwYPjOpaw+SkArYI1DdDcTQmLiP4zho0AipKFHj/fcZX
`protect end_protected