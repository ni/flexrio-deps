`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2016 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
xI6xg28eTBkT3MzzlHKeZBbTE+RvuiPmhR9IDCKuD7cfdBTF+1JKD1tO4fBWpKx2
t+jBSPExgRhFFHnhv15qM0YoPFwSn7xStoDX9Ax94409VcXahTo08eQ26Z35MKfl
her8MubweYvNd+0DkDrJjyBrGExyScErGF6K+KhQ0B8U9x8HyDAioW7OrrfaDh//
iwDLKK/LNuzIM6FJbjyWKzRftWkywipggN4MF6Z3u+ZcuddAnQahymUaZqaBfZMq
aNX4W4jtsJcscQxAsqBlSPPlgzDdpVUrdjy9AEfae7bPfb6Bm79Q6kWDlWoeWY6q
x1/hI4quCbUJQzT7KionUgBHpIbZ0YJebn2ATzBehrV92jtYxV4GzrSv95X6mOod
YbbcUcsrxetcxNgnUO3i6uqxVggHYgDdojKFfA8Zf6syJD8N13VYxxbVrwlFjTFV
v30/ai2oegvK3R8vYqVqycqH/9aaenyuaXGJCxxC27+XOtnRiXfQB7b82DIyTi20
Yt6jrkiWUJBZmb3nDisWckGiAtbrLAVDuthcTnNYTwjy60V6EA7kMD8MdZu5pmsD
mNI24AM87kSmSjm3K3rmQsn6kvFtPGxEd4PIDuedCHuqCqWhKcLvwjHJFXh63aE6
eTucamJitpUWSgJP1R2P2t82PZeJLQf9H2UKeyFvcTji9TT7VAVq7495WwGlvbIF
3nUMl/ZgBxbe4WQOWzNh96qOwujmZfTP8XEdvo1euUt7wz6q2Rd7IJvjlYqiCO8R
jVM1bK/6lTgkHgsSk3dQ1oH1WJ3DgSem7IaF5K3oECb/FNGA2RQbH12PzJH8kUNx
36LmFDw6LbCTNlvATYafJgDx/BNiQL883mHAKPh8F/T5CmftJ4BMzT5FF09IFbbd
Vk1buoB1B3oy3RCo8CMfqSGCaQ+VTK5gy9YyR+FndUPEGjdTbKfikv01iW910QPT
4ZpkRYpIQv/CAFWXCdt0bO4X5ecW44RGT4G1j6R71PwnddFH+HsXHPDrOU0VZdHt
xArzqdmrJq6W3RRXBcKyQTHlVZ1RJrZ9K5aerM7BwhQ/Cdg+3+YKVWeP1fglwSIx
dn1qmjP9KrHcVzwIpC/YSfnF90l0vL/aUb4N7PF2M5THO2oeAuJSsvFWbHiLEfI1
LYS1Wi7rnM/H0mhErjg3a3Av7Xq0FA3PkXRRtdSio8ficrqablhTx9W6AcEjH6O2
zkTvM63mDDjqBtS5rzWL4tzeBB6D5wGjv5sBKJO0JijCIfY2QchSkhu89G37Jf3A
IHALaGI9aLZrt9UpdFCQ4aNZnMPJmtDGFOKwEX4p2N8Ed4BKpsZZWwzrD7ZuN3qk
H6+dh3cSxUyGn1AQcug5zprznBNOiQHbaCX1j6PurFDLFmnk6rn4fQibrnOUSQaF
NSnBgkvN23MiZStDEsaffgcHGEVojoxmhBg0ru38KPGAoNA2J2u2cOI2ERKrG1Jr
EoqWaLyKIPY4MS8A87pVwN25yr4Q+rMMkXPmJY1uQTBkBF+FymAkEHPiqYYAiEY+
Xskj/tfssFcJYR75ukPdzE/fsqBoyNkXIQS2roorGelO9lzfgpL0zEAv6loR4gd5
dYHLVI0Akjo1gSZywKCxRULU/1cCcCkl12dNgjp2tR4rgvidyzQ46LqgmMKoLSgS
mGeWaEJVLufKf93mwrDj8up0OIZChocGVN0xZI8s37ReH953sour2lF5bmNCPYPb
2aI7ENkoSF7W0XUJFO4H0po3vV+go7SdXLR6HEYDyEKOIAkG7hVjpVGI9IZ8+Kju
vMSK4fZCyl61qiU9H5cpDODLb3pqGshSfy3mkpqMAkmPseOLlQg1/Biq+oqGTn4z
pW7koerLq8sPqedHcIJv6xvpbtdi/3yM/Xncd5Wdt0SU10BHw9tscDIvJi/m3LBM
vPJ4ZT3fpqwKnK3BTqNgQKxGTC7csSo8ysdHinz32nlLK8Fe8Paat1wh3vfR3UzB
b9FUfP1+TNI2CDCL0DoSFdN7rxW257tcixmvhPnACW0GIZdgwXYcjeDGXAHhJiBU
37e/OX1W84qVmB16DSxD5339D7xKdkeVxuzTKGGpmZWUNt27p+oyTnjF1UkiIMT6
317f95QoQH394LuW2LTXdoccJWDPqs/gzULWOljVYCjvPoFJP+iyIyZ1bbR7K1Ye
E7G0qA6RXSnLpFrnDkaFxzUUJmgra/FSX+D2bKe4lAkSwuwEJlTn3LahbxsKIqF7
JVf6op71QB+MiVYkSTThyz6TkVIcm0XJAKM+PFvvqSnhnZW9nl689wagTQIBvm9l
TT7J8GTqtnVHEUbVzfGasDFDqXS3CbRfomGSahK622we19iwFv530ANEbzWlY16D
7bK11HOAK9tdXB5TuDzwZdS+19TNaPE/Q07v9uqergr2QoFcIL2iTLYGE7jm2jty
Gk/lW5wBA7pN7lOaivSvModOOiYjdSnSYxOE+id3WeFvm9n/3dorsYIu6FyfEFAW
EdxvgcWvGemHSM2zv0Rcc07vxCDeQRSIqEigbXInCa9FAxoPy3DXoBrWgbcODdSW
`protect end_protected