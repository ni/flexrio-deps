`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 61520 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
FPPR7ws3fN+RQyk1V5tkgIKK3Jr4ORg9KG0SJn4inw8C27ZW743Jzh8LKS3mU7vp
fBmdxeEbkou1jf9+CLfeyVe1QC52NKDXDAKwa9ppBZpA8UeaRwk/r1+spFLVNhms
kAWdRisN3qzq3biPF2xk6EdEcXB3HwabFvPXJ642xCZBqZBR6Cs0xuDsAFdMaZfc
41rP7MAfOHFzOrt+Pyj4BrqMpIkFn9Y2HAOloxoBgAPm5R/yzqv8zpZ+y7SriaxT
bfOEsHq3lcQV1SDubLHXi4qVDRpt5dsDLDsT392R1gUXuLYjbC1vKIldN1FzFr00
k2c/hWkJTqQGTXLVVzbEsdhnshg56heeHmgCnkr+Ts6NEso4ITFF5pgNkg0CBZoN
XonA0ujQels2b4Dy7ipqR8FMpueXZt0rg4tptdpNXLdp5p8gBsSP4NZy2uUUCN8h
HIzjSvCPPaTB0ZSvDaZig6kfBDQaFVxWrtiyS1qr4c2ove3ci2qsMhFdKWUT+Fx0
QFzQlPlSl54YXgmx29yBKJP4eqe3KHRod4WjNjdl+PEKquIc4bwReUF1RNM+vZLD
trJsjAu95EXfMUyT1JeBzgobrR+aTjkAgxcB7mKtcQd7d/xE6aovOJZmRbDx0fyi
WpApUT9ClhUkoQ/NDFZspBUHeSgdQxd2qC6BMVQVmloN3GKHZsIjJ/UI/ZUGAXOB
fedazy+dOf08Mkhsdt7U1a8yKsSGjT3D5cXAlaD/bOA269b+CbO15zDw1FmYD1Gx
YaIEG5EVIdZH6KqJ1VAhtRDWwzvNQzn9bhcJULCpMxqjnNPuKdJxxO++/u534aMT
Kko0zMm7XY6ao25CtE0VJO4uB4RBGUYT9VzPnKUyePXR8QDoYOf/zV8leVrFUG3A
MvEj1HC//bgph6afdPnLsyJenxwtnxtizYFNqyUidHkNTQHonW81VTrsZGGvH86X
hJcbpu0RUvsE+5T6WPb2FQWjuYFn0UKfWWPqzSr2NTE/mBxCqDInmfZyjRXkUu1M
rV22nYGK+2xE+IKZ1YELawrjIEmBXFi84t9PGmOKPJY7+iIHb8upKe8lkkCh64aj
Fj3+JlSdk+BtdttS2HgA2FPe9xRPNoNVHI/O2ROFyoZQL603Um2FGlRzdwtjFwND
5TfWseIjvvCs4yEWXOMLsvH38Oun5AsCWvp5LX5R8970Fq3V3RLY2+Lfi0stfy4t
l9jRyyNfKxz+O2ulnXJ9oLRgg4AEY0/6kdWynX22gJ409gDwII6/Kl1a/Ui8xQBe
Efw49XPmSdSaiH/XBoxomgpmP3PMqPZmV2AH0XNc8Ck/FMYSNXA8wQhfUxxKmqSx
PZ4CU4yW2AAEpMpx87whIRWgDXK2eHOr+2PSNcpR1aVfIiA80cGq4TgQKB4G+sb6
JOEM+v2S6c9pSV1DhuKFh8EJ7TK86mf1ZzaH65yjb5jn68h5v5ihM3VJwl2852oX
keN0NYBq5XI6xEM74N6d0iB5leEmemoEjMyF2H/viK1MX2Ysn7tIOz9BigBIj+Wg
QSlV7Ck0ioyyKLAQJpaSCvwcn6+P0fDnw4EZ2wsR5hZmPxZFzLMsclrSvr0eK3zw
CKpb8PScV+1nndO4uFdGMka881bDZn/qeah5a1qbh34sIfRWvYVx21Ugk+Nq3aa5
JxzxzoL97Ibsc7As2OYoNLcxP6c578NPKMw834hKWhH0HCQbQXj7E5uiIle+LMGG
t82DExX0qvvccgW9ysDuy3Co7t7lIMcZVundHl5r/pRM+PI/n0U5J1Wdfh5qFUK1
JQCPr+BhH9L2nj3tsE6FpelMd6jifMFBfPDYInxBu7jineH62wjis50oM9UAErFw
dD6ndOdj1JmpwIjJIAmcskUxzkfSw6cJnNIkYH9cxUPxd5OXnnjVw3Me84mgAylF
a9iXQazsQG3jDIEVUzqVoDaybU5WqoKfK0B3eZIJZSlrxwCdD/UbXBc1WfYdQk8s
1JFYoEz3ynwM4Y1HVe7NaFAhazOZKu3+KtcrbDF7DBJybG99zJOfcccShTLB5H05
OP5gtQT4Df2XYq9I7ewSUJGTbKEcY9lGui1amv1+uKgRadcKg/ZkAHDCGOx3vlan
JYaJvmloC0Zi6MAHVZIkAIrkIhXslgXqsvR1ZxFZyFR/AGdFYMf1foclKwKk9rKF
vpxRyY7yYU7RrzmNZcV0RVR9RhzhhV3cKwVdxcFCHyPgTd84mQDYDvV4n6dAKm63
kHRng30vH4ZtRckzum38yScPLvhD1EV3lIeyQZECj8+GIkkDmzodlPfZmGFDxBZh
/R/5x9it+iRQAZVr0/MI3FzP8FIoFkXE36vVFXEdKcEXjHXGD9e4bR9DJCeSLN9/
8bSjKftjBXJd39XeDALyG/zOjKGRLEUNB1dlfAxJaLCQJ9yXesC93vIX38by/W7u
xZPkD2t2WUAGJ8oGWEOJMw2W5O3mkmG84zETQ6EMWN4rfEOhVcDR7RKWq5C376+X
KigJZDJu7vauraT5c3xdOQG1yzX3kJcP287mHZfVKkuqQX2PjIzPXeKe+OjU2Vxr
yy9+QzQyciWfYZKJvjEtdPvw9SPjCiThCEr/tm4HrmtvCdRKwcEMyCTdPdBo9d8E
SegTYQTcxwstMTqJi8J9906o9tisei8jkxcW+7zSCJJLE6t7MikDxPX73TZPgS6/
8PEef6jcxvmmvmI0ZZC19UI7LbwWXoOn1dKfmKtUfyQhZppF7n6mpLLpZlSOJolj
SqTs4upeE+gusCnxxpZEjIzmgPmWlMRuU/6LtiQl0M6T0PbsUubQG8p5KVyp+Ooz
d42TfKC8faXfW7y/JT+o6L+HW5ebcacgRD7DoBt4+hwVoifoMdq/zIl/oiBfCusy
j+ZGOCaHwPgfsyabAz7qjn75R3yZkBj1Ik7KD6I2xLVRDP0lEXSZ3myS49f6MQtp
k5aTe1WiwYdTDrjJl0B0WwX0TKvkQnp1I6ZqnEWYhDMZKeb1xOqYE3PdM1T1rEF4
68JecbD8SoSPizXqo3xaj04vQ5o3wRfzksmNIJfVIiFFUJKg74bnAHCvUBqLIgPN
/vjaCqdbM56NQtd2sBtvBVCnCEyOzjOK4LjSUoQzNlZ0GDSI1xu0Qtkd1NTztWED
yrBLHWZzWEbSqK+lhVmvVMibjLb8nt0uFYJ3LQ+SFoMb1XVA7hy3GjP+nvf0A3EJ
emMb+oUzRVQFW0A5o6seZm1e+wYQx9VZUs813q6nP8KZLisPQhKbpuWvjbn3fNeE
RFXcmeKMbrxz7Xxwfmius7+dFLhYzcs1si+e4pFVgoAGEmNyKQRURCszw3NTa7Kw
oY2UEghgFfrp7Nzh7hLs5I/7d3OajSos69hlk66+fixiAPiYCECpm2r1+drqZM4x
Gux5ibmkPkNhXTfSU48ozB18mVo0V2/znA/w+WHNzEM67IBA6rDFcrRSiRWOcYj4
vTYQgFFHCcjuh9Ox0aVMhY2SMkBtegYKl0mDeXxx/EZBUSRmqenOiJcdArFjJ+ya
4P+54C1j0nhVhD25qesWLSXRDFVi6jrKMiCcoUDHrfokeY24RKbVUQGRFvgnmouc
Fr83PDKa9oY0fkZVuuCfPqOcaFkUGcBOdDnr+OU67/k5kZKGMFHjAEpHWXeOvDbJ
oYZanKPsFjHsKYEngW+OvgsMU5+XRozr3jQYovL+Uubnyd+c0euDKjTrL7mKBPeh
xmipSLx7xeCDwkPd+0H6dOwZ21FOMJSszsbjwX+QmSdzaMNvGO0Siwvh3IXdk6PW
s6Fav2E/op7NpZrk2Fp26Uy7Xz3K9gRytBHVYBZuRnZt057VTmY1XDlbM7DsTQ+a
xuY64gBdrsOsnKt1jIrfb04fJC32q0zEuccU56z3vSmbrBRuo5vZwuSeREHdV99F
Cl+RZdqEHCM0kY1brkq/caohFQGa2wPrsm9h7XSzJVwLasdGXwayPDk5pKMdCniH
VrqhOQiIPTI85f02tTkCTZlhmw6mBI6eKTm0a5b3fZ19UcWMBMqoJm+dxi0GWaIV
BGj9hjNS5TtLITrt9O+jeT7yGaUqO4GWEMChzv9abB5aqN3Jl1b33velHnN/TTS6
IqLX74Km0fotdwYGARQ6y5O1fmM+WTfyhhLZeRvPk+uz68tP5C9FMKKbe4bgsYy4
s2NLg7wUubPMhPlQ3o+QuxwX3H4WnH/ugGeGSmQp/iXMWrt9Yh9YQDTUGB/wY5Qx
54gWGGEW7p+xE9L9cnT6NBwyEcE8SCOgC2pmtRQYl1Wlqe02fKPYCpjKrOAeNRJz
297FATZkSSBWUhxF7cOlvvQLIP4AnkFLw2+cVnGCr0TQcjO9i4GfO6NgjYBG8CLd
NOXvuQ7+180dW1hmSj6+6UnJk3uivjCORjV34WYRzK/N5uzvOykEwtUR3Nwi1a+k
F83K6CElHCcrB9poLKr647XPrCzIl75TMVlHPM4AEefGR9itCruWBg2VmiUtKNsL
xKBuhILbxBZp7VnLP9Q9Ppcvv7CUdevzbR6mqc1+hqznsf6vNXaQCzhE1VcBqc9a
dyAhHzIjTJSP1kPsLMpa/YGq2W4PnkLImpSa0XqU0QzgZe2S5bGyGLFKKKAQUaRW
9muQfkx2oyYzhU3QF03EVbzUtuSgmoexMp/0TWNUoB2ci/eIjHEx0o4fYEah3qNM
v9gqpDzL0gA2qpmfB4MXfhb9ttriEVHUlGEziiRgDeB7w0vEPRVIzeHytzg0DB/R
A/R6IojBjPxeI0ZlsX7YukwcUTbIchd/Yn7eRU1wPXtVKc6WQPIr3Wn7akoq97bN
tng9S69CdMAubUcUT958adk3k0RISU5nWiOJCIt8UeKfk1j8DiZXTcWTmdEs/Pr7
vk0vFmzcnRCnisy8uE0PfKqUHD4KhwjnLzVJqiKQxgp3Kd3MVqOCcjYKMNlolZyO
TbnfwbMEjQcumlbt0ozuQPHv7Iej+ZyMz+Rdvy1YO6/QSSFixcYU9Yj9LW8Jjc59
VyhnkypsSvob33smOc9Tq0SNBcpzx36aYlFQv3CCm3PWg+pA5jAZ2ZGBH5EDLhaD
6E1wkTF8YGKY7wz19YYTZoOuUmfiqNodnyHl+GK/S6PImst6VgveWbOtXc02LVxJ
kMNVWekBdX3gme2APPUpN5wFbpwQ/Yw/Bo0DsptjzLjQbrqs6aamjoVgmjglbWMC
wU1vTStlocf/UQZbWGV/GKWNryoabcaItEapGA7FGBN27ujQmPUDntuUKGJWnCgd
HlsHkmXSRxzUWQjZJDHqiMT2TjAAiuSYPFCe45sdhpG3dQgMxzJsj1rwL1E1VRWj
BHYH52T3xft4Mv+22WHyTP9iZQxK2hIhbE7Jc0pDPOUA/glAlTc5M+u0XHX1uKdZ
RQ7TLjnLZoVOHPW/5fJBbVocOEjsacaeC5N3ydaJGIhPPjB7fTSG16FLRrER7+Fv
82DXFARJZXzKPVrJYzbOMvw+01FA6xTG0O9ctRhcaOC+L7vHLxOoRMA4HFFV4r3v
js4rsScQAMXyJyHvKXvXzszW6qnah4tP/qadccGbwmhUk+O22SVnum1Wkm0YXwUA
xu9grbi64gFDp5mKjjpkQ2UmzpCrCK0bvBwHhrzuCZ03c7vvYo/5bdMI4JKdvdmV
3agdnKyXjRulgaWmk4AaaGoIlihoxoMu57BDdow8ZWwwpY7Ih53tSwoD3z1UjoHm
a3mvteJU+asN0GR2BNSJ5eYhOdFe1gphKBBBTB+GgLSsr7xvY08Fqe0qHsQJv1Gy
K3JaT4sQdWAhcOoH9GqUAxZme9Z90zfKRIXcaUx1mVaeysL18/QXVItWUbfVHzuQ
LooR8IYfBw5fYKhhUzE2j7JpoHSgD9ytkc/CJa4OIDmvnfKSZfQ1BUiQo7bpjddN
aHQLuOXudnYgM5vPislCm8Wh0nsFbWoDdbdGoaFhVu/hnUHwMovmboIfskAZZ+NJ
jeGiknEbVu4vkZPS9yDmVshxnlNyVwIXqC2zY61bXEIWWfw9pmdMK0OyECqupOVQ
jF9jNS4MrLqFrWfDHCUerJJ93xGTQGbMcN39g6I+Y5PXUhJ5CAP6e3ksSSGKdNL6
SflNSmTz+yD3b2849A7xGtnrEj4tt2FFq1/G+iuzqcmxx8bgOFmW217Q0xyupinE
I4j1ZJIkRYc8utJMzIgvat81Z/Les2GjWQwRdFHjhuodwmKLSCyZLog1FCwjPMnP
4iAfM+3E53GhYUIQ34DuiVQbkVVQlva0sWE3f1NK9W4W1eXp8oD6De4GeUgUcuNu
mCVaf/H7n9e3m2TNWjnEUErEQf8LnDtJSfwnaRpR/ojyjzLKdRh2umriUpAUx1vQ
fcja4I/yy8V6YccvyubNKN06IIaGTvViWyLPTcKgmTQGrMixvVyH4M+QJ+iL70u2
VF0qbocYm2HqUp7UOzgjWC+HD/9viO3Bp4JtGNWVZCgJ8Bmo2SGrYxJy444X1SaW
qFLytQh6tNe5Ggp/i/KcMTTi8xDOjuJBFO+qIF1Cu/7cVogNtHFzejgzug06zM+S
8dfshGx+ibnciuijlqwkA1Su0wbCDHO5wd6RvcwbesbiimTTlRKc9An6JYq3fjQV
cxeE96uSCBVbnk/vJZSPkZVDVdtkA5+dv+Vz2kJfcSgwJtVB7vH2UfLVglX1wtc9
bBMB7jh47zgbsy6/nhgqu7xEsp40GaeiDwMzMNr5uBIf3Kas3XCYfxCMCBkEe9K4
veO3KkcTNmiGiI42HUxGbxPuLcMvrgzeWuWka6yhyLL4WPJR0RI8h46Ke0AsFZLz
QXRxrmPfHm/jUJELlH2AQs+Y/SLymq7gzag2v1gteVldZclLKEzl4w9gOWK5X/HV
DkODGw2DvnwQcPGjbXtlxeelIMDwb1laxY7ZlrBAZW388tRIxzki3P/7ph47Rdo6
BxSOuPTNhDPZ94cW8HM6qanC6Q98AQN0WTge0uDLMC4aohFtK+DEeeFz7Gyqg67C
bXeycnp4NnuRQ3zn0LsUWB9wWsc9pgUlAqavsdN+x6luL0RQuuegW6gjCOFswv3H
HAaIJWgFGdxZPFHSDA5EBAuOd0N0SRNsGNIJ9V0CY4hyNDd35sNyAFYC3mRTf0C/
HLHAZvYcLtOyle99DpH+AtmdjjY/AxjpMxhnwYERxXFyjRzGzv4ZQQTJgpXoKeC1
a1DOJJJ4nYMRpKbKkYX5dtd14Q/5mWykS2LTvlAc27T8K1sguGde+SApy6CRjPL2
pI7+FpbzEtEcyAZi00moZxevb9XGiF5tVpahh/c/FUqnLmkNT5bkEKQjJCfzqjDU
pnaDm8sM2APKhS7+jeXDGO8LX7BHXC39b/8RjpYk3R8i52LsjcqDuYH29O66TdEl
X8tOrjgUVTjMVQk/aeUJvIQFcNgsof7CDLQPo/YeZQ03vjb+A96hc6fXo2T3ZOFs
b7Pj1LlL6/qO4WBAQI2Qt8yDU8K3aubxhEvIhVuKwhz9dNbm8WAHOjpYrcGN5rqi
hKYXL8DjcxV7xvUetRcD6RZSSxwhR6sXzSXxa1WOpdDnBNJEUw+OAfMl3hhWoiTl
r9KnDSxoM2df20LUxIsvz/O5oZwncNuJq7FGTr7PJ1wHmlMpqWQ3qzS3rSbXMp+E
KG5hd43KYRx+++udu0AMOOL6M8bPJ/Im/7bDoIaXSF9FKPQfqbWr0BLaMUbZm0uz
pjHj19prLNnd49+RYwovO1GEQaeEdl2PXX4qBNfJhmXeGWucjWqEDV/QkQ5IHDkG
SJjNgIo95CtW1w68lt1/OLui+OccjmNITbmy/HBmBMOThRWArA10T9XvcD/u6a2J
HlG3oD1hZeZMntnj2Dhq8HvD50+XYag01GliDXdL/ewc9rQOZ2WWzpofEISmuNKR
M/uGoe3MYgCv7EYeK150wNaTly0AjKqdDzoteYD+ldfJIhWXGp+KVCYPKOIJ/IFS
aYjL1DrxakC738Doa6LfoFSsucCi1qQqoCn7spt/LzNq6Gtz4db/eeZFFUxZACLq
Xq3lIQrMCJ+a63uDx/jrVFN56L+jNMl3OW225eZA3Sy6/DsM8hK4drsgO1L5/Fv0
Xhv0HHX9k5IZO3mFmM4tjRCnyRGa3kr1b2kkHIs88ehP2NIU6mkZvXhdQEj25XaE
EJ1jtg/9BRmAeHtliXmbbGdctgg5CnOIQWjmVS7Fe5Is83BYgD5o+7u7vpmftoRX
WWARY3UNcLNG/cUje98K4/DOkFxpw2rLgNwCsT4/4b/0xK4Jkg1pxyUlfLczb3WL
l+VQ+Ip+el4fDODJQ4TzVoUphNQbCw+HR3jOwZGispV+Zq/9MaBpXjRH+hSbfQB5
OU51U3FfFSWGkbwdPZVxhuHt2D5Oa7yHUZEk81bbWH8eDkMNmQQ8dFsTxbZqMP50
J2EQdLpEwYAxP/YVltappi+jgb4iQewt0svT169KY/mrlRVTsk7DtJ2UWACjZ0Wl
biWxG6fLYQZOtAot8YY1hKADShcUn3Bevt4Ay6UQFdqZ9gcyqbvzwijs71XI0zeL
5DS7BOvXf5SWKAKz7Au6pLvqt9NpEhlRBCkNa3253PaF+0TW/SUE4kSXr8BL6jd3
t3Gml6UFy+1ZMxkICuAR8xUnaZDwdS1KdRrHJ4bbNrHEjqpz0/9Rfl4TVN5Dz68p
Q3H0L5zEk3GYVlSRSGYOc1Lt5NltxyxCfojLdR1GL8+8eKvxNjwMDmhTWqsBQZRv
+lQHCGk0dzk5jzVoK3NWzAUVxZftncQe/4tlCo9a4s2wvSSetwD7JQwLnzq8ysIm
YjHlHmSrcDZGQl9h7GDPdMjLkiCjh3i1zQTFl+ghnlGP6413kcd6hpQjeRLm9SoJ
cJxRRXoeaRz/g+jMbSZJYp6hYpMYuP6j2wuA7yhAMp66KDcvTmfYY9vgxfZ3nWvx
adKumB9LmXlo59yKP+gqMuzpr+1y0nW9SGJ0ui7SYjrVqQfoTrrgF4YMBluZxaRp
dwZMH9g2MsTjxICf/xG17Pb+XOV0biqJi5b4o/WcIywejiI3XqfimNKM85ajz+Cq
mmesota6ewDnmPpdLcdTBoPDrqreCFKoaQIoQ6BuykxiS+W0fxGjNzXaRujH+ikD
jZPATHzN2Ik7bzG1qQopSA9rBm3zUmY7w/8mECp4d7G+w0pyOwuQ02ZyccVC74rL
BMgpryb6MjganPyQIlqZMbmn7NQV8jXUjjUmxLGMMhoYybmt+DAuln5VXZtCTQNW
sG4tKxGEtJ78xJF07Jt1n8ylNvjhB0IdwiNvNLDFYPCi7WAI6TMEoh3qq2CoQauP
C7Oc27OejZoT/xSUkeK4keNRa2MQz5BjfxFzWRdxOrwBMX8tbwtwXTo0A58XCRsM
tRnaFnWfWdx+Bbfg8slE1blg4UsPOsuIFKE2g4YJauX1dB9AFozeyvYlfnqleMJz
PEMEY9wmXBV+0DiTYC2MtizA05XXO5x824JtLCm5q6kfP0l0QupBjosdZ4uIdhAP
ZeqYEKQzOa29HNjVUgd08i+we9BRluf5u8Daw3SQSCTZyHHvusnzcDz6ObLjkKTi
rQy+D67rORZRon0genf+Y9eQN0She5YJgHNyIbSuon1COhCbOQoJqavBkeml9GlP
tHcm7g8tqU9PZQt9mSPobwqibLgNinM1Sz6V4e1NAaDVG3AGOoUaOg/SLRC4xcdK
Z8EhThjMnK+JwcA0I+0ImDQGjKwv4W2R/OZ+lsdX6OW2ntC3a/53IElBY8N5Ijoa
9rRhRLzJASSgLj2DTIEQlS4E0sAuuUOiBFHu4kxUg/kCm7AbFLGdQVBJcJY4iA5V
f/BQM5hJEKPH5aTKf6+ThAHShQkHMRNSqmZCDnY3OA7ftwBvFTkrOGZ8q08T3+vV
vieVZvitPbW4HcMrSRzBO+EDbh0LSvOiovktWYzOscoCLIpeFnjW+CGE9rQbkeXy
SKIvK70z/UQye7imExMsTDpaaRBiPt+TaJIK2NgBRrn6QqrpMKxMZNw+B8LJR7pd
6W5WPxZWK9uAYamRyFcZQ0ITai9zd1AHfhy2Pi53dDQpBKLsbSzeR097WJcRP9tP
hGwGB7J6F+k42R3qj0FqLWVY2r6bPK/RRFaUtDg/5QHi5DW848bwYQD6w75Kr4c3
dXOJR8l897+8QiXBUkjzAAwNG2cSpRxR3NrfNfewx+kps4/qdyDeYfe4862ovFx9
jqdqW0oAPdf8e2tndK5h3w5/v4f1IVXFFsTEYzpqbYZgFNyT5Tmio8oiJhnMQLEN
JGTal5WqoccfC9bcN4F5fYiDD+o43trWuNH7o/l0vp4ZWtQpqVaKudbXRQfIRiM8
BLzRvUD8rh+/TVJYLp7cJahZySK1LtCOG55zmtdkQgsr8Dl0UotMxf8vPqYQ3TPV
DGbmMirX6dJUjh4xjikRskyIp2a4i5FtIvhbeGcyVccHA8W84a/jd1NoPMPhXQWP
XRoIobCd7W5usv4d34x558+Q3ACS3XBXZ5kMusDn3OH4Mzi3RTgAiQBkrUsCVi97
FG38Vygz/Z0fv44CouymIh81KQmpdmkefR9yZDAreRFtFef9NpugM5F2NPuGyaEh
h/hiYJE4dnc7bd0cDEI/782Mxhge2duKIUG2LHaaeaqoRyfCuU+ncw8SeeOExTK1
wChJanbOlMIxkg7KeqlzfbnPyuivhCGcy6aGXBjTLiyKCHa8t7ko7g5kFyM5XJ1N
awGuSgdzRDfHKtxE6t7BDhO8jPxKK55lnhoAGQBPbweC5bpiF5AGNFNCxg9uYmmm
NdFWRZ9yN312Sh8W47EY/EKAk7bA2txVRtsHU/mJKRuZgjUdlfNu87xpmdNsDj1f
jW50JAjnVHMr3AwcYe9KiZYFPtNxYrDQ4fV+8IMgYJ9VS5xiRxbX3N2Zi3LfrIPy
uLaVGQCfiQioni/RcR3k3A1gYZPHFGA7boz0w3gQnP96B8itUpO5iMXiWBpRTeZ/
rJ9LwVEtHBujHbphoZNvqU8PmkEuDe63QphP0+97mNIRqGHLIk9SmVTKBQ29Odgn
sJ+u+wDqU/N5O/TYqoRFtRr1IQ2YrfqArGxEOuBRI3TwDeFnU4PVH0DgXOGMCGZR
CsgZCLQiPKPtRAnJbCv8zHV0rDRe2BXaMMsmWDCmn33QmTKJuq7aIEszTDAsus71
xcxbKzkfoHWTT9g1pdabYBOQtQDyfCGFYi5OHj5rFdUUnRucEwPEwJbeIeWSR9tB
XVvzwalO+HgoZeX7eLzFtaayvrg6RgReq9OnifpL57G4FCz4sA/6VK529fpZh6Mp
z1VKgaYe9mwGJJSIpHN6+h1CPwi1nTMHFU/UdamVTqUR9yIWVSTAf6U9Piso3Of8
K752+AtHYzKYbbujYVAaKgTKlSaTgvlW2MH/KNoKmLBK86U14SgEPRUupmAmrs6i
Oj5OS7Wr//EbIwCfLdao8Avu/UXKDmTtFzamAww851dd5vuB30sUWMf1Xg4Q34ha
sc/7RioTKGKozRw6i3/+T9sEDGdRoL9hnYnpXKdNTaJGQfjUWByNu2YAKIgIN8rr
N+e+vh6ptHEyNjoLzLeY04qUMTlIDqS2pZVQCSfVDf8FRwdGZXYCIZtXItD7a2Zo
nJIYt3BR4Ks/b6hLdU55pJWcLE3FkDOGxFj7JjkN0cGXaWfTzlx5sqwTxkRozDRz
hELVJfJeGdevM9PlnqFXzpyWYDOnnPAsh91oDfjmSybl1oGvIMsJJ24CI/sC9u/b
9pJfEGh5+9O2NufXuCawHRCVqVO/hsfeK47vdvhQEmJT7y5N6Va2JGix7fK1ez6/
/hwe4TPVCVSTacBUT5XjvxnLKBaqi4A7NShfJQBrNnVbXznwGmBX8uHyIDz7k9MC
XpnPkRolyTzdqIDObHkbEZaFjI8s8iSsKGNnGczrb8wKORMFVj9QnVT5Hc/DXxeH
POJoae/gYIibdbSGUHTjPuh6YisL2+sHQkpcyZXV86x/Wq7E0J4hcqRO3+fa7wk2
xQwcigcX0RQhAnO3CAZzULGbJeda7Q5aBW5kV1+cRIDdqExMZ0qSh05aHVZUUYKL
PPavqQYuoTMA+UL2no2gIn/Pgccq6/CRYxI6L7azZ5WQqZWCqa6xzow6URBHBNop
L5hNRoFej8tz0oBx7YR6vDd0xIq/lbfDhqr9mjALRSlrR83G6IgiRY+KZ69f7t1O
9ta2EwQYud+sybJCdrhHNJs8y34BcwzexXM2MaqY1Ihw/rpr+0rCT7pi9fbpqqVH
pLlwaM1EFMu/StOYCV1GGorp/a2D/4MSHeKI/y3OZ5Sfnx3ON7dFAT1sghD7Q5yR
GDQ0SRTwgu/aV83hESV0qgcRSWGXLz2YUVe8Km4ObkQp9RKkc/8ZqdIpV0wINvFe
x8nSZ5WwmmwG359/q9KbKoALVoU2O0lPeU5U6Cvx9A6JZhcigrtn8RV0+fGMsDFO
tCqtBSjPv/YSElkW2GCZV6gyLKTg840Hz/g/KSTZmWjH8CF4MTBLAezE40rkQLo9
hivEaKEYyeO9ku2WXOQTCuEv6M1elidRssScJ7i5shbimUvbZINNMZAvk+gJWqt6
A7fBKogvPA7RrCiWLLM1AFMardNFc37wfVhqICrJyyYWFL85qL5gJvaCiBFkjcOf
oAp2TFHZVkxzUNj4UH46M2awCHWmctCvYIUaDvWTXk4m/4mWQFfTjaUV3rG2Znr0
gY2csnc142tnjzDx0FW+IV7rEJ4KxDhQlARVYHV2oNA6FYs6XGKSdhFk/LhsDkk6
2U3xZwvlmb7Xs5ZtLRUq9OiV2VJHK9aRM6vjBzWe0aE4c9tWHly9tokHfYU+dtxK
+joUCk0RuvRmOCUQA4f7GuRLw2fb4IF3OI2+iXq3pgLRcTG94dMm5C6BZX1nrVuZ
FPPDB2NKSFyIEKzajvB1Te2e2XJtXogpSs60Ve8xrIwQV5saYiFB9bCxL+1ygp2/
UJIpwW+FpoZB9EWUpNL6LLXK/mkwz2FnQ39jPhSQIKfZHj15mL5RTV2H5O/U87pI
op/sQ1BOQPZjTLBjIDjMIKAYx5kI9pBmeyBbuv340bVwbG4PV6ZdVk4HK/8D8zzo
I6+Qd/Lf16xYtuVqd7Eb1++9X/oKUh3sg9p9S+EiYeuj9rtGhqVP878vCVV3Urdb
JXBHPADMpIMyLvwVkoT1uUy24TmZIAE0x555SNM/wxBZ4OxJ71IEVh14JnhcpQH+
Gpc0sqvK8opPAFXlxXwSKE5hnonWehZytZz8WCOoyiuFQK6+8C4ZuXnUHCmIQon9
MXltYZiawvGNAX+DwyTDBJK6mKbkQD7GFhyTBRsvA8I43avnoQsNq0EjBBjSeoHO
m7eOfTbWM7r3cEoHWasLyx0Cldz8JUqX7rSYsh+hApKOCLNP+L233NOB438gdY2p
wF0evBN6h/FL+Ih15Fg5vQu43uTfFXFXSJ2w/r1bbJEiX4UUf2uglUwuK7OVT1tA
kfeVby9dD5jKiaFI6JnaLmyMndruvaYchuHVCIK3jKiJyxfYEfWgKOPst+OQ+xrB
oN0luARXKX7+ptq3HG72CV87F5v7ui1o/dDL/eKxkF1POWZHmi5sjeZI3q4PKZdS
/omqKiTU98UgIk6YaYhmentD5n45radOuvsDjxNaOXihmHbTTl0FG0nlLn0EuUFi
/6H2axM1tWVM1qirjh1aEG+IJa7FgnLtpNepEiRHGpdsXK95bRhm2hdnziV6cwLM
4rAftD4j4ZYOppZOymnqH5h8zCeQvQt1342b82HPAunKFkm9n35kVTQyEMqHBMW2
LwDPbaJrysNr4+huErFEoZ6dSAj/eMCosn2pTEeVb2qdlpZ2xIRFDNjJPkhJWonp
TywhTJKOkk+1YInVDit1n0+agQYVwdqtdy8nBlLv5d5SHewW4qkPXBLp90anSsm5
QoljqGbwlaie6zRBR7l3zP3QCQoyhU7LDO91jKC0//RAaUtZFzT2yn0yuX2fvL6V
aln0SbxyaVH57kQdrf/Uj4A2wHwk2z6drcEoXTH2opnAGb3TjwBGEpTBYgygKA6x
hYCWuHurHEaSjd242OSkdlTCCeFo2zCm5JgoK/hTpZoOLSGIeYuuAmV15F4p/w2H
wMbReVaLVui+4vEw8/ikZuNLwJdi7fZA05dNsvdx45LgdjlLMGKXdfL09ruWrhkS
ffxXMyZujsUw7E7m+pWXxLhvH22v4N7KtGAcDi4OqkJET8OPQBF9NaFrSOL9KADf
2zmyRUBICVPilChSVe8ZrYfrH3+MJxxDD039DMfW6NCV1ztve6lQFB+d0W9ufnQN
UGa/h0XRenosRIuNIGPRnCAVCzsu0geGkBk7eSLjnrJLbvqyF2KOCn/CiQYXvjEW
WKMrf43DMx62ogATjH9yrmc7nuC+QLZspgfSjknK2liiHnm53mPnrELIK+xgIeps
TSBh8slwk1gyh+S3h4FiNoO8bJNpOp1ssbwkhU0PiDDZYe9GF1Yg6DUiJhuowMN1
OR07utER+wWL9ih/OUwv/h9L4V2x8jxEExB7gL81WMt9Ml/VRXPOOWKTjaox+cWb
g0NXuHx5JwOoX6VlNBgeeLeDJ1VTfcAtvspQaIBAVF/jYR2B1zNalUWzlpsFAmB0
WmJ5Xl3+r/1KE6aagMrY6f1PLk72fJx4QIDghFC4185mCzqpdqB3Yypm6vWRx0FH
fsgh+6chzt59MpvjF+v2sFN+G9Fq+EVvfYKxdu+yeZub+RCfLqws2dYMExzQb8gZ
hKDW3Gy6Et0xvLuCXkrNO3rOcRip/+ImZrVlllqQHckf9LOvUKe6NP55fN3V2Aif
qeOKliB+/E4NUEe4yYqlf9O8t/OODkYKt22VtsJQ8V/3muy91s5XzsPr9AqMdNmM
QQhbd9CtLiNiM+vtjC3rxiL+aCbwAugFd+3j+R88QsC+cXWQpc/nMEAf1ITemS62
Jx0wVI0stK7SQ9nCI+UAlDZzKhPmxqygn3NJ6cONOLBn0iwUorovJyav/BBoz2RJ
pnZ8Asb6ak1da4NvLhPu9xxxkyMjhv0ksgVntwJbEl36lW50ykZeCQf12VcnkJDG
swjxZ4yfp77JK8Po0Bp5AnrLTtE60ydtLuLjorbk692H5ngJpT6KZnBN3DEd+E/U
Xm+zvcS22qfE6wQ1bvGztQllgwCBXPUcyoTAn/iasM8JJUXan9WHCLF7kpEF2pST
jOFYZzCgJo4JgQlhW4lIKxW6VUW6naKOabwONYVpx7drgTT4i3wNYioETAOzH8iK
HjOJcAEjs/KbdVwrd57mSFAs2lkTdQmlvi71szLOGx7rueSwL0VXA9V4nQ/I5o/u
gRRaGgMOcf2nh6hMq9ycNx3GOS5WOz1cmX/oVze8kIbCMnNojd73PJRMIE94GnqH
fjuiEDVI0WBEBNQpS1OLN4EfnaualLeM8WGDNK2tBgAnTHURFkQwkVD5+tAA8Vis
8WuAK9rbzfTQxxICgC7PEOP5/Jhh+ZD9DrxTVOHwO0NNL7q5c5Sdw0aTPSXfZClZ
8qtcbQOKWUpkaaRgKWCh076cWYJOLVB2+TTYVOPluoGjdix5z4uHqr/jUpmVF3wC
RSpcXKYUUUn73K/oF2tVSz++JZdEWNd9sNZEt4lz669Py7EP6MLg5hh4S9bSxv18
DdEk9ge+OY2tEOmAXYm1HeqY7FtnOOFMPZaJ9k/C0dkHnHb5N6xElzMGLUeHeCIz
VzZW48Q8iAOdjGKT217eYr2fDnNzPs3PzrOdiwbEFADpDFmkJhkcgdu3DzWHSp1+
QDpf9ZVH4NhuVKw6waKlbQLeBQZCbjecX2fB9DjUFk0O4f5/OLizTiZ+k/8eIamL
x23pncsyY0zDITaL67ixpLhVrgVcZbSFhHkQudcq/5E77XQF9Zjwit23ybJETnl9
kvTpkdTKzMwQdClzsZ6yFSzBcP/lx76HR88qlYXaHga3PqQSh3jQ+rzLt/Mx+nR6
tOUBxhSlmunrkYYlk+IAEvDdi+4R6G2T/KjXmbNRvu1hZKvWy2eM2pG+qbqRTiDP
BtuzkppdW9DKVuknY7Dhk0iDjoTgTNCZUfB2kjWY5B4QsGT9LoglNeUXQc5KbFXL
5CyxxFD4qdeA5boGVD+a9iReZ5X1G7bwROSe4uKuCFPUyWRACb/mpnjEbH964Yp3
+nIjrpUzWUeyfe3s+IzjO04YKxC16rrqFGgXJdn4n1drOYnV6YYbyIopnkHM1h/h
68J6wW+h3SWucEFvD64LFXukL+xAGWIifhCqiSF7GBjvp3JzzTAiNxmjmRjVBmHE
qQyIsGFU1t1djwbFDKdWhQUXmvAJu9ZKiHUAaucPqSt1Cp8Uqt2iaQUNsXSWf4hG
CuY63+XxzeGfvwQmEPWui5WfcUZsl3cP6WkeU6QfgIdBDgblY+eS/dztel0ApV+H
RpBJ351BECZEM6J0gWWbfCnF0DnmpJ1Fke/bHETy/HkLQl4FVdAs7HxVUrbTRtdP
EmS9WERjXEbHZtkY7M2FF4sOWme8aghfD2+WP4DQzFD8r3JQgOuShXPoLdYIZQhx
k1euYcVRxnmXnsoQlJQin4MKwfobFY1Rmxy9UvboemK37VcfgbhBsufB64Mb8PEL
P4j6v+pyL2IaYfVacIJVKdmdTVUfvZHXrXCqXacbwsm1LBQjlZLdwHlMteB88/j2
Yt1X5VcolP0HhVfAuBGqvcEvmLDm/TD/yFatp8tlfydFPUJafaeM3U4vDIS3vVEG
Nh2WaxYI+NZo+9FJnrTd2WKSfX6luTQ5gGLMyq7OTFLt4gl6jyYvqxyySi2k3loO
49z8y5qDH4rmg8UzQXHa4hpJlZc90vksFMBSKm8SPwwqGKHLdmm8z6BXivrD2UJj
rVixAszRTA0mcl8C4xpdPMMHX61BL7n3aNhvDmailrT2O+EdcRCdMtn0BlF9fD30
+HT7AjnGLzwhKc1Nn6jMjRocENT0i6dUcYFtR36cCUrMhUiqKZW5X+I8Kt2il/lc
z+7RuZZc4XwXvEFMvYPt1BuWG70lxO0GwQQwDG+nGBLMvQv0ooeymklEgHnIjwav
f6tplP8lr8vLdOv5YDh3WyFU3QLxRyH5C2+5xmY4rmaJPCSFrarw1JcE2jqYbJnk
3KK7tmry4p9YeBwMPo9NT5IKD11bQTYGW0pH8MR97YOkqWJ1j0OT5YBviaQPom48
v0H8e2S5cZbQ/B0JhTvzvQhTSmJkI2geW4hi7W5bkLzGw/nG+Fl4JqKw7YGgt/Gh
xwCl+8ra5izODNo0EbFTUGpOXC+QCJEldofoJM0+Lqb+T/gqLMtOB70y0fIf3zmI
H28453EjW4YkNeFEvNjtlfQyXQH7NAZxFHPyD/EBfbdFDfM0jJjR9DLl4tQQerw1
t6X28O+y9XVX3ud093M/xEeJxpyswF+UaSlB4AXSmxIkkspYTn4KqOzNEInF3epm
4kpZWvzr0poVRlqGsKLnZzloCJ/KNkVyF86mxIvmYiWoqIi1QiuEh5afnk3MxGgL
Nz3MlqfIOQ3JR8GzO+DjBbA2RcYmWvT+J7lOG1OAon6oFcExe2W3IZFBF1eVjVz4
hbp4FTUPMf1G2oP6zlZ4Gxvl3GssUPcHIWVF1D7RfQjbDZX9Zx1akRGdttauJunZ
3SqYsFPe5kBbO2sQv9pLqt2r5gx9g47AIBIwxcNSIExouzBo+BUAW6vGyyzV+IxR
bv7vsgn/1zOIn7FF0gzzQBWoVkWl0g4bz+uMvTRgxEevUuQZQB3uQt9/F0qRIV6V
OFhHxl68qpk+Sb8ugInQRk0jWtGApGdcXCB72q40er+PMpEq63Je0t0bDzJLVesQ
ddwMde6zwR2Gbh8YCGLmKavGGpQ/lw5UQuRzR2kb5MUOyPUCqj7vyG1jIRaVK7Qz
EOKOXWHKd+wQqVULNiAYXKjo1wrdIwqnLbmTRKeLVIuAdbpSv7mTKa1ymreq8j1V
5cWRkwozf8vIrPkWxwPhd/SFQJsmu5JAp8xwHMiFrhP5zxU+B9EnlA3CwmnZnwac
pov++9TX0zUwmmLQfBrA8iJey/Ng5roKtNOrZpfytv7VSwl/LzRNi22bi3yZSBey
Mym5RvBZnae9dXhx8Bs0MCRP5Clldf2whEjhhh1ZBeI4YpxLnuUJ1La7l/f0wj4B
T0kX1iCQ9RCj/tO5oJd69/7c0LduMH/2ClWY7AUsrRDT/aFZIGT/YcW7DJqzlMn4
7CfSdiSRc4ggKje6je2DFOdMKRZbksGkMZBAntE/jp5W4kqna1ndU4bGg4fJb9t2
Vk/3cS8Ybp3I01ofQ7u48f7wv3omjUglERAk8ixS91vjsRVmS4rlYYnWO/fZKuIQ
t7o+OSzG3DUZmgRWc9cGF0ru/AQ0Ztc/FRP8TU+9xOxkYy/IBLhKI8pYF1a8AUpq
YSUpEC4bfHPsBEFiPOGpsMOEErisBNVIWSfWhsdevHne/aCzsFwF90mLksDNy/aM
0Yc3sgd2xwgPZJbXOGr6NHr9q/52ayCLjTh/7px7EDMzJdHnFffYYVwr6tts4wby
GNm0v6SxQpkIbiELAj4k88hDb8uK5fLIryOQ+36bkti8J8w1v+y1qhoNNN3/Rw2i
2yg8vTm9SxII0W215KbKEP9OkJ1gJFk9zBWhfWSIRYti8bKw5J5JMtRiySJorqbk
j9XHqlB8v+8lCNDoFgRUhTjL1tywzs9rfCuqNJL/n+f/L1icP7WTP11Ruh5Lj5B1
yRGK/ww0N+hnSEQnWfp2SMYoNT14SZOjavptr8vxIu+1Dk+SBYM7tkggjKc/VN9M
lleImSFXufipzk0wqA+VAW7/Hv5nvFf/DENlwMaw7IZFuf3WNQ4ulAr2LpX0PiXO
ICGSvOgfqFnBQVKWbQBnjGO0Q7RbRR79INLLbkNrThgLmmpbeG7UL9oxauLkaCYR
Dp9+t+mXz4OJaz6wbX/vYuZPXMCbkVtgl7Bahq38p21dgW+8He8jh5asf1P4OJkn
1EUH2Ren07M4ANTX72dRSE3aaCEZ7Vbka26b7O2fF8UXXHv8YI3s5iJnoS6yli4u
EvQlKGkUhm+4RaUXrEYyyuY1XZvtsQdiIY7ekKFd53V9b1DFBzshZ/0CIfwlUxar
o0WnaAYZ7mz9FxXpRmsFjOG1KaVAVBhITvAbHsNVIVQbLVPr1z1Byi3SlUd9hVsf
q7DceaoqSrcSoVOH1JKD5/89WpdDcH33kwG6QSLPJQJhmtDaP3n97ADMdgzA/Gin
1gYm5b1XfgzCynRus26PHRHoti41a68RmsN8mfsrqfTfdaFfOYTI3iTkdAgkZ6jP
j44aJOaSyrIBW3/SwiOGccjRBSIXuTAUydUbAauS65bPwBVYVXHFRc5CWjyj+TCV
+wEbIbE0DckO74bUPl2UubLhnfonaogWb3Q7NB+tyqg0p34j5fCa1QKbudq3luyl
23UBW2TtzGbWK/qheBdaVZFuD7SqMF0Ba2LTXGRTZHOo5C5XL7873K5I7fTngX5c
KEN4bWpPFb8eFzSaqUReucY4AIbdSkr+ilt3DfwGN2vLKwtPu0/9U7khQCr+xdLY
ENPq6bLaRqSAgMfPlFJFdzEzXXHt++6TTQPi2T0PVuMMw2pCyQ6PztPgyesUY8i2
STX5DCepHQusR0aiwqXLGjMAgv5y9OsTMyw2oAlsQ5AJXIAuKixjzO1j10SYv376
VkqaFJj/umQWrpOv42ill1FkYEyuRIVdrEJJRPOzUOGHoBPqt5FH+pBanHlnk3PU
5iO/R4DpAU7MXV9I0dQH46oT9XwPeQAfZTdkJ7bAt9ZWhJtpodI70wxYcP+DZcEl
O/8wNxqGM0aUgkO9teh5ieyUama3p2mbWU7zkzCEwYDPT3ddywUAkDxaTB+kTeJQ
TfkEO1AyQ5NIA9mz6RtCiO4qG33lE0JUN4OaoKvSGEcFOKy2WD4nz2CucICpe7fr
pAXvzFu07eir0k0zhCvu0rMLuqmIcKbwn/78MBidEQ/Wpm8//mq3Jce2gqtza9B6
iUVPWA3vzPCXQ01e4CcBp1O8MADI0w18LhGtlso7oNOvGeBzyePbaPYuCZoJylp4
MlJAlUgUcsQGftQCUoF6Drn1P25pNbhEOH3xtn3tSdzWCFU3MxiYekB8MH+XEEDI
xmsLIS/NPnOj+5FyS808/jIi0DQ3qTkbwM9qk5ijBmEZgx+Yfe/NArqefsfVhzPl
PUhrsR3qGWUjgI1IG4h7CDxYvIKFs2V6s9vbvlLDK5VXYEage5dBL2XM/m+qHPez
7uyGx7YG6vjXhEOesbyhGvYfpOXK8vR0eDzGG+G+mM5+/7newjalgMiTgOMige56
6X5LQfYq05gy/sIn+9UyNrzGVqkZM5tHdGk7H5ID9ruQZ+hbanha839zGwfIJu8q
B/pDB1QksmFFl6zcCXTO/M0Jm/8S0uv3FCvMxLahmjOFNehEkA/7cK186F+zq2mZ
uG25ZGU3JpGCRAwgCm34+e8SV/Tgnu19e+w9NSQ1miNh0Jrq8ike4v0+9DFMS9pi
5t5icp71BPinrgysepBn8+gRJVenJOhC7xzdvKDy+IQbwozB4PdEGpCdv8eNMZTh
bNbwHND5I/WbvB6xBlT7rewXSRkeTuLaBe/zgWDwlfxADzEi4eA1mAE/M7A6gfor
bCsaJ1bY4xG5AzyULlj+MSXphWSmqcbw2eVRHYFaWJ5hPHixrztJxBpNji1U8QFC
8h62GYYcYtmTqVViEpuP8LLcwIRs92Xhm1+hAHLnfcCEqBn9VjltTWFlgSwYFHW3
7IO2Kb/6+SkT2e5utq+lFtXX79N7yqoorNY/WVHo647qbNbvhnUNFrCEkxswGhJ3
ApI/fN3F/CshwblPLOyxttfo/n/TRO1NolYe3BKfUu1Tfnc4lIVOoGVOrFtB4UWR
OqO7CkAsKowlmPXj8FWsJDwv03CToCucHlOS9foisSHu1z7vd1JHYDNN492gxbxs
H4Q74QdlUwzYEnpkVwcCll34iLrt2SboD9LEUISR0OoZIagndGttqP3v9kSHrOPK
EWPZMh3BQXFSd17r+2G9qy26ANTeg11QdAPASSjfsQ3GiueXal1t4IydZcpgXsXO
SzkKgVUppmNSLgYNEzxFt+h9w4ISQAaJ9l19zvlcSOhGfPlezNHgUwBmQtJqxI8g
JqmPMi3eNS8j1vx2t39BgVd/zp0cZY/9F25X/8Do3JbhbykeMT+3LAjObiT4tSZq
b3zSeEowa1RTCYthI89auVZgY6gOjB9/sTO1rvQ1qJXC+6D14cv6ZsNztJ/8Kfyu
crS/vveqwzmcSfeKPae7Kpm51kCZKTQ5iPYjmqGLH6ZCo9qUEBUupk16mYf25hGU
Ep93uteENHsxB95FMZHNo+cqqNHyxQEsswHNxxFcLsnJYv5gORea6SeRewIfKIMn
pimNFvYzCz4m+kcmvmNt0BwhG9JlcDiNFTedSzRblWH2eJlM3iG6kWRYqrUWZY/j
uTvFQXCISkwoTdzn+cmgRG8FJVS4rvh1fxlHXk0QQ6hxN9qrvK9c3+Uj0wb3NkPu
590L3vJWoGYuqEPA8K915+BUFWx+z0RwngM0/+UMsDq+dNWGySjFsd7PudMQTO4L
mywLsKBo/FjJZsIGQCM0xSk5k1PXZ2N0VrHuaYc/4fg9WJK73UcKSvKuReNSz0fx
tBCiraLv+a6fZwQjw+Z9cTnpkP3KFkTn5LJB6zfUsvfk2Tztxq1hNV1UL2pTRblf
qJYcT4h2QWrlfA9YPfebLuMuzLpbE7y7JLBcmAv4PBpXzbkQwn09bZbjlPDqh92u
iegRmOVV7knTNIU5eRKRv4C+04f4EcPPa5TQ1fSAIQkoxN7VcH9jdePfWdfemPaB
V1wKf+r8FGNQE8ggCagEhCkJ/IE8B6KBMTlo0Dc8retR0UaPFWt0IpHd5V9xtV05
c1OLppBYWXZaZRTSNP99HnONcazxb0b91YnyiDO+r4LR6RmdgSEVBZRhkTOBNJry
mo2fAS0LR3roGxrNn2HFDTladXIkd9UPLKLYTUjy6lHYqkjF56GzmtgEbseS8VuN
ph21cOSd2KgXknNKFuZNyltnB2bjrAt4oZC5ui8NO7UYq2COjOJpkY6F3h5sFkCr
zNc4F1y/ZfEZAKB4zFK8CkloLhak1bxbloJTsiO2tEMIJhWiq9xwuun8o5gcCTne
X21IrYpDZvQ4azmLr8xOrM+MDSTW3bglzWpY6894SK1v7ODZvzvJEqNP+2g1cWEF
iAL57jHERFYyuq7WgDTg5PRADPiO/1EuDzGoOmoU9OWpeM/gJOAv/yzzD3chQfmw
0RZfm2MitBJoUBT8/+MoUqqorMbIQoI4po2FATNA2B30p3b/wpJrHvDyOIcDMM9p
X1pVCotsGaYT5j0rfQhyP7Zgc+Gidp8W64LgQwkZhtbBkmeTN0SHzYq4qFua3tUM
rpEum8NvhIX92MA3STd02yqYeA3jPG3GIhRQ9Y1GxwJWtH+FEWSxm1nwkpayRyOk
+tWQRIDc01fYOlqffoQbktZGckcxbjUrgxw+9sSjNGAuZIU5ZZbd1wc2KjonBV55
Ikugi1WJBzaVmEcCN5mOo1xzo3S9bhKokGjSYAAgcsNV6VyUxzK7liNNB/RX8fK6
F6L3m4xZj0jlDNq4VqlDgSWKPkheqOpvzqBwz1nplL9xsMwaGWILFjzcf5PJQfH1
DxiLUlJoi7yV33q5IADtUhHRF3wMfekdQjqI9J5zptPZwnwTVacTF3OGMyZ5sM5Q
mA6ZMlgZ55CQy1tGEH56oZGp4/uhXslt2/iuiUApV+F4XwShNV10wanjb8prBm6K
ScKdhVE8QTF+Pq1uha2VyPKleukcY9BNsGPMDJQ8PVCASQTHL5np4IQhgILxBXv1
Xv7iHkzzAESk6piIhzNgJcIN7pqtdwj6QbBq3l5moxD0nKdhPlVM4au5zP4kKSeT
bR3lC2n8ocJZH/k7ueUGn4qO12psN+sFwPkIj7j3LxMYyeX+zYRPVC56kJCBspq7
46rnGLrO4Ji+9YiruJq4c1WaCjvs+zXijorITLmn4/gw1tguuUocrsK67PfJkEYJ
galX7g8zfOkHKhViIK4j/aoEzrGxSHrrixX4aMbqOOpZUiboKaTqxnInOiF0ViLs
TtE+g8u4L6BTOh2XZic0tIU0WpTY9e5GfCYyeieyiOd6s6kEvKl+wCxiEltw19SF
TmnQAaCqaAwGglYPySOC0Oskdl1p5ytxpxqR3R/p6bUvXgnusY3grw0QnI/DCmnA
azDi9eG6dfz9Fx85+ptSX8De+OOCIyulMpnINcZhlnUo9KuG97KEignLNE1AdUDn
4obdxHZRjUtoPKDie96+cQpIlBkJKVyVYB/JBL2GiAdYI6B+RkRX6att5ETsK7DE
e5WQWkHeLyKDwjXY60AQFFf+UqZQyiZbbyrP9h0b3KP3L5NG4Egu0jkbst9koPeJ
lcbAtt0mvIDlrje/x5yd4qIfFjBQoCW22Oe4ng2LgSKmFluB4b3DZpmvlNkpmm0l
Y9JMTQPcVW7FekCcEdhELmqyDICxwN3eiVf1LenChxXQfwpU8KfTiAx5hy0ttVB8
6qJXGwzHCp2P/boa0gTRlb5jS6LRQqmOE4dZTjMcTvqBCk5iK6qAe875XLKhvrE1
Q0Mse0JHOzmT2a22PffdOeBPR0xMfoMY2o082uPdvrye6psg+9u0+qygRPDCu/hU
HyKpbDoqBYf/sNmqMBGFQPGaC+1VQ8cZ3c0FUGWBtCHwlsJ440bcrWs+GeqxG8ky
oM8RwxMuD8igms270bsB07NxdIavot5whm+auIgUYPaP84W49YBtzuCR9uexbOme
CGavR5MIQpOG0hJ0ejpjpWQKmI54nVmLIZynISbFjZJwHrfImsMWA43mGhQHdZyC
dgizULPh+asjy+Ys0EjTVe7I+3i2mRIOKSAPEmdrDYSXyK1AqUTcnkW1u65p0TPl
64JMHIRLfuJC5/z93GknN//QjL9ICUuk1zPDL7GnkflTvBJ98P+zdE51aUKqUQf5
dQx2V+T2T8Eu/P8pQ7J0ZFvaXPhWFwKEUDZjb5F8kzuDuqhOwLRtpbCAG/spHGiT
qDjeoaAYmbWn9BfA4KDGrfUR1fN5d2ZzOKdEx4OUIIBVQWd7yfhuDF37/k8ANSnB
9V6HM4ZFgGAScsXARtoW/VVYTtkrHQ5PJIkN53G+s/5Stc0UdR9WtF23O6qfaTw+
mB4DsA90xBWYWhdvXfOInXmxvc4JvGfAsZr8Ux+t0WC48qMoX2KeXukFB4s8EUAu
fD+07u13kMFcoPFoqdGL/0pTCeH29fR5kvilk+elaVDkJhMLwcM/1h8tOHS7GXxc
teqI6Q2ZswdoeakVo++1de7tkOMLO6MYJ4Wx/xgRAQZVlXO6o0bZ/0JMoGzlFtyn
n2Sy0U7/cYw/LJVdajTdxW34uMbOmmiZF1iump+w4f0GomCIG6bhsoSucv1gwN3a
vIa2lSnLjvdCqv4sQb1Rfv+S83dZRjOFn/vIEQhnyK1Mg4Yw67QMIpwLAYv5dBWr
QmsLgz31zHKM0vYEx4vsnp4p86UodlML7HX3fKubaHobuK2Cc7rTthnjBy4GULMg
7ojd4qieNiB/6s1d2+SpKVl4LBG3hM+vz8gyanhG5mtuE502XKCgzD13ROk8VG+z
TxAW9l8Uk1pFq+m0zwspXv6JngNlsWiOGZMiBilyXxryULY+cvuEIUTLaQcijktR
fa8gMndX4pdmpH2ItIDeeQQbNk60wr1CiOE9bD44J2cci77zYFv77ku4W6fAfI7F
tv6ypcbjRaWYzcNKQVDOYkixxVe36CHAZFsxprW+yiUuqW/k4VJ5rFG6Zq3W6JUa
4buemJJFR/FQl1OYIawd28i3Oqh9hZGUBhvDwQmFnAv8IZrILarVYMNZZ3s9Os3j
AXM+yVIrixO0LTwwgXncRg6llavzQq9EjBphU7LW/IbxZUBxpECACk+bT32kn9gR
ZLzq4sAEwi/oHFHhhdLVDGFwzKTwwIVm2IBA3WrkHsfw2261ThXdvMf0tAbneI3O
yjpOSBhQ2/zdIljR/1yk2Bspf0RT/+yR2e592Xt7G/i4Yp8EMD1TIPvDKTLXvFfu
v5rGd9XCRXlnRlGFdvk1te3rYg/9ggGejCSNZNUA7DfV7uiJbZwAIoG13Noz3Gpx
K0hjxWl08Ix6woZ9WOGtumP8y6j+v7SqHOGxbM181a+lcaRDWI3bLOkrVIQRj6xZ
gmtuVUMcqrLGXLkY/jP2IpLqMRQg/AzfokPAmHwGV1ZZ9S018M9mY8mbLSFlyY0v
xCyirigI9PNPBZJQtchTgLz295Mzf8D+xwPxh/cSSqKqfgbS5T1jVTXt1XzRfNaz
em9SYCceWkXTfso6z9xlAa0zOtImoZQrVrbUy0ckM5e86d9NrfdnTl7Lw1p1uxnD
jlWfW9X4SF8Mwj642ye7UFlumJa4uOu+N1a2o/Od5iSo1Pn6e/XPAVmO3QtTYvKn
PE1NEm3fHt9eYPcJyTPgv5zcrQsG8D0SY7B6oI1CPsBdUmiE/JhUE9Y9kOvRuw8R
005KT9ZKqmYyq+0XnjMtZmywooswGLgmDN1zCy0lai15cTPTY979sHcko0YgRsVg
7yAN3BBAbK1RaLyNoeHtzfahyzLGmRRK0TmxnCh9fbCvcTbWC6TCCy5AM7w1QePS
p5DUcrnmQZHs3nvqNkhNxNMbwD+7JZ/irspOw2pifOwCn/J9M3W048CDdnE8A/Pa
zKJCgo92WLxQs7I2uZElTjF1Q8Gasw/TeVc2Nt+ZM9cyPezSdPM053/m/iOtAh0D
MZkNTCsxWLtmS2TrUHtElYPU25BwD8LuOBjBmMC02kFvR5qmu64z6QLlBdbQHxgY
16BaZ0L/joNAqBPQtROsNQe20UnnsUMa+hQaOXO4wTbZaS8Ye6nR/tevvGXyf0WJ
cYF1Orfl9eMATwtxYv2GT7v2vr57bdSiaC9b7c7mI/r+kYW6DBsmdddGH17kGr1F
CoHfQiZWOSCumSPFbWrzGpvbmBZ1bZLfK4tQ4w3eU1w/V4i6LbAjdDU460afu70A
ktJiaM2eo7LlImAxIpKUKNl0iVmlcu7ZMN5ayaqFpZnSXq0E/0KBD+wxJQRthBN9
YLsTazD5tjhoHAwZtxev80FaaBJ2L4si8DTiF65CKxVilpwOTZ6+B86Uaqnkmted
vze1+Jy14oLiP4xAcr8Y9BpE8jkZhP+FSEtGkOs4jdus6Lvd0GoYrmPI8na/AEyu
tKhxnnNO7LLiWoJTZuEVAJuJhcvss11z+wE08CcuSRYoCFkfOVIB7KxCdxzbXH+Q
FBpgVbRTWSCbigo6vbi/MLTNZkfyjdeY1D8rbHPjP8BQGPxX/XrH6/e1wCrp10Eb
5aeIqQGpS3zPU2xhZlmsr3sRUFVP6rsR/hW5iQQRLpbMNzsG22wzCe8+rSKuJjol
ufjIKeSLgWrLI1UfXTEmYk7KTmtsU6QYNRsGPIgMiMh8SJrqdO7tLukuM8LDjHUc
yCuhuCsD6gN6whDgsbMAj5b5CFQzRdsDqMV4kYI8I9zjUx7H7tasGbM/WsnjUyKJ
XOl2OSeJ7Fe6VTCEZR7NjoP8SLm4XeZsd4qu2UzQ7xMlLoY1uUGMLP+sW7X5cK0G
bOdgMlDTnGtpXe4POqNy8ugGeD/FfKGaDm/J5ggynzbu48w38ah17E0NSsM8O6k7
nmyUJb2TAAx2RYdDRni/tOV6NJIS3LH/sUjtDlU7y+f3NonWTx3Dkndw6O2h4Daz
v/PYuwLcI0GoMnsVj6MmMxUgQNF5Sy/8uy6PueecdPagAKM+arFvTTrbyL0dRvBe
VewLnMv58ZCbsxnvFFfHZjCufK5OgGXKDXBkdlvO6pnq+L9odwlCYHW07LVTmmoi
Syw8vj9rzsB2x8bK4q3ssmo09Wztryry1uSSgmfjVO9sX6CZFIn+sw+lhjw8qlPq
zUuxEk8bZ6Tuar7CP9I8aydy6PdnUCnjCfCZjNEBIUd4aaaeTEWc08nvlNNin4mh
aK39yCp40YT5m1iB5CuUujyMcuA5FCE+Nec6B9z/CopCv86Mht/Q4vjAHXExvvDo
Oo4a0Zc0T2LYtwo4zp5FO2zbTyV3J38ur365l4VXMYWOA1D7CFMSUeJhaA9e7ccH
CH3ykGI0YWdjTDKnPteZkrTSI0jDgJh5L9WejVUWB5UhK7ZW7YQ4oYcq5kskDhlc
LhnkqwtSBrDubsO16nLirWpvMaS3lYV36GgpURh+Bakqm0lBNZsoSIlc/JMR/oV7
chKUF/KG9mzuJNOkMMFYNfGQpPA9awh7QYZvofmDY8fGETeQiikflbqdMztGRL4/
nAPAQaVb9/DeXEaYk0ggRcY7kVi5U92uIAwroY9/bT9ush/DXpmA8207f4pUbR7P
uzv/J7mdnUKoN1lVV7gwyffLeFl0VFn7mBmBHFGTwz1NvFqUtFxWo93bpfSrf30m
NFIGG5glg5PGSFf1d+L94CZNU5fLvi+5a4XZXWIEA31O0Wp84b3NmLVMaxw5WRS9
DKSISvcoub1sqotVSYDlppke1BS9JiK5Dl2dRk27x0m+WH9LTwiUlg6q2hTjuuF5
8BvqqVa455GgGa3bc/SwTgL9lkBWa2uru/TPOme3l14ICaxMSjekr3CxG+HsVbro
wVJlhYsU0d52gsiWgcA/z896S3CNhLFy0brRAjc/RY1xMLCskfjK21MQA1AqqsYH
5HdYsVy1+c8pGzcI/YodUlyiHl/6cO1+4wQnyeOInPy8AuY7R0/tkmBUKtqkasMd
xdBrDtNSjEn4Yq1w+dJBuFxABOVl7ZUKlV5/BI0S8LAlL35x2wfFIv2DTzYEYM66
734g0mUhp+K0426vMbRte+qdF1AuenMkwSIvPG/BrW5xgXPGoMwTqjq7M7ZpB1da
TZ54wQBzwLRZ4OE7QQnHripAOfZt3VQiuMzvMprl01bp5P6MqzY+Egu9KXy+ASAR
LYbqs58stZZcI118s53FJp4kWC9xwe9oC2WO292eouSyr72uP5cIC1ztCw8cuXww
/0cK+Oa3Wu4EGQPGXF8H6srl9u+ENhO9OKOdXOfd+bNNZm/vsY/S8+cPrL6KsBBp
HBFb268eOdYEGTi4Q4T9KeYT0mTROfmJGPFKI+M5RcxdYDWHjJjKId84h5Ie5YdU
E9ciqXNGVGWtRYTicOV5keza+NbCibAwX1q2xH6pkApaqOfMKoCdlTzxT6058Ef/
ZqPu/wfoEJt3HZy7CGBzw/jnKQK07Qr591gXIbW/edyj+xiG8O9MBfjqvb8UdLp0
T2Dtopro//ltXtzSzl7BY+N/vj5MrVet197sN//q61sTYshuoiCnbxjJaFu+FmDF
xZJ/fA+CSX8MG/xv8Ckde5gYlRBPBpGwpiQOeTZNq/ki0S3dTvbuYNkunRFRlpOp
ypsW2WxOXDOpsmtYNVeVgptzVlRtLFd8RmxgfhVA0SFRhWdh6opNdONH8JqzaWru
0CVJQ9St0792y7a3V4Cp3FLUY24SVYEJjdF/PFTSpgiJ2RweTJnFRxumpk3rlUu9
nWhlHUOWh03iIK+KT8n4RJn9tYBD+f5/UJXoPZK8ekWoWgsQK4i9na5jlwQWihWg
uj9uaR3dV22mxitUnhJipslE64ta7AImCKNBWlpfedZpk5cpdwaEkTs/x3zXlboM
wIv5xLGQ9cEb6w49yC1pVT/8bvvoWsR1M1JLP7d7KVycSnIf4F1GOwLSA3X+wq41
sPFYqf9lW+VNaKyS32LXrZrHGOUZD6iXUMYAY3WSDnOhOX71fQyPtT5Tqnw5c4ou
GjC3FXQ9IMEHbuyXe6Ow2CN7N6gMVyY1oMRja4/HtF/4fzJYQYBQ7f8xPW2HtgaB
EiqD/nIPtL7D2M5uulhU+rN7ZdsZTw61T+bM9CjmPErJubKa72ix29cFf0jvnYN+
WpKt5XhJHyNZmMvkTW7oxxLmbBb7tYOdzyoLDXU7KM6pDgFq6JlGXxKqcim1FZgK
dvhw8bWeL1Jt6t1H/zraxlChuUWAZyuQdbtrYjRcPW27/WkhNrIBH3iZL3z5C0Ck
UkE5EzLFyHQ2vA/AQ93bcq9XHpM5vaCKY+rJ5LWT205dvgJ0Kgq7QVexx2HRNHql
U2GqXUl0ljM5Yahg5l1oolFI2c0RH8rI5e+EWDQpB1A3rDdju3N1T9+saY4G+WKw
qHx1Ga76fB9KB0A09GZ97ljcUwc0YbtF8OobZqibb13Ssu+6FIWaDqtM1otqUgwh
sSoXlyuH91x/b6v44YdI8B8FjulLaFyFe2Ng2QUQfMq+xgFqZDXEQ/qoA5rcM3E2
Uc/b2Z+EA5RjwEYZcsktekktsL/aWz1zBSO9256wUf9/xJcUlosecm6pu8ATuWMH
WFUs8rkPfjNMvovRbeCGJGbB5HRimGrREPp5liBo29hPw3NFr5U8oetzeqDmY7gg
iWWYTWNFiUs70c8RHFpd9m68PuxQ2YRb5Gt0NiE50m7+dd+3xGncgZBsSgMA2ed/
BPMFmx02HebvIwRxoV3fu+ytJ9d7Smq2r0SkLJ5wJ4PkZugEUb9tCIf8tffmLo4G
MKWTQ2w2Pmrq+xjBYaT+QR7ShGXIl/sl8nENMf24KNe1F9FeSk9opaXUZEdXGTxg
uWDcR/BXXF1fwo1R076ac9ugGC6L3sGqaPdaLZVshbvBjllWbbMqPiAXEQsLst5n
GSj9nG6gjMSXTt46/BPqVn9EEd6Z8r7m8QdWw1qL6sfWTWRXX6ftRZmnGfjSNqKY
mQzs1Vpxo3nlMTrzQWcvBYHeXQTC+sAWWtXBqwl5VBm5i40BErVZK2A2yGwNrd+g
9G6XweYbxpqSdP+ldQMRDJlKSgs4opCfWLGro3b5lt7Y/SENT3G6IB6dkA3fnhxS
VU5lvlGPlIrInMisSu3YYVWQ5uqo41sFPaHsmi81mX/CP7js7kro2LfzTyYmxhWQ
1RR+TAOuP3p5zDEiynnaAWO1RBmfKtweElWmkfn/5uyIvOiWaN3yuuLqB0DaisSs
TTbYk49PZRjKcTWW6p7CA5GtX3PC2rvhUYPFqp6UJ1MP3dmbUZ/zSOyDvQPDGE0G
8tjYskyuk2rX8s6KKm2c+vQnvoG8OPu434+1tEXk+Zwet80GTv4yIcwIbpBBOqvE
Y0wnWMYQ67bERrq7DYCAW6t0hyL5MwoX8pHTXnNfmIL5gk/LIbolJIiaFFGSmfF3
5dRSoB7pzr1cHA7CXe3NDtQn4YYqpEAvTY37sMkQbmG/BGxo31FtRMiadjUlUgwG
Lsop7ZxWVjBRIdQKu3Ioj/jxj9iAp+N8/aIYFSuumA4tWI83w+jMvL84unUgLG0F
6xBfPrlRseL9JOHbul1wgjHOLkQT95fN88QVnQRyUbDRts+gjLgGSREb+49ceZ7Q
ST2Zzlsz7dJZ695AD0Mf7WiSE6073tFEZCpLclQAVZQKPr3ngSR6b7jlIZKdWIro
K7zyb5I7GhPi+mOlPKtAG8pj6rvCE38a7BGqGa4oEV270SUTjndnyXRvXE2Fhx0a
GZFHqJBtmBEuC4LVis7IvOkDIpS+VrDxypBtZUx1rsXS9wQ6jumlc8kz8x6gT8iy
RltDJhAkbOFs2TOtWmYegpNJ70HBaFgc+I2pzWYiAZbZUw8EE4MZZaaKIf2/t/2L
JyM/vwhl5ffmeujTDs+GXT8i794QKpwez28pDfviiOHjlzl0mQi1+dyh1qOGMSNN
0qDXaHf9TjOhPu9gnkAzvFFLQCj11Ek6f2hMhDN7frb3BJ7SGq7Dl64yRHoMwBw6
c/YJZ6EzDHE0cEfGyPLeNwTroJRAf9fOlmgGMF6tAaxatSeVP3L6/X/SoTpe6shJ
k67JjwD95xiUHm9xjXxW7GqHbR4K332O9CNKAA19t38029Q/Tb/v7cPVdEMeOss2
Io/tG2OD9IoqAF+ZrQJ0PeZOXVRgSCxfwFqTl1p0/bSYamu+HJnV+ZS9wAGKHd3g
q/lNrQz4Jaiy2uShHWe3dPlTp3BnjU3H4eT9HgvD9NgghSS6o66vzucD5Wgvyq21
AeN7rvO9DHXc7dpcP/8hD6tBxaJYaxNzd6VZ9AasWnfDXBHiITJWT/M/4JIrkC/j
9O66A0a+89n42RV9V4bWgQJbW0SjNawJC3Gr/jdG8XEDRvf+uH+8NRq7lYd12aGH
iLuaoUBuBtLH4XpxU47yaetoBwBAy5A2fX/mcvDimiTJsWRyhPA/vtroHG/hCiuQ
lISrrgqremWlnJWqVKZ4mP0Xvc7l8XminONc58a9UW2BuKCZu1y5TP1LUl017BFQ
ORmpwNSTUeKS8AxqWdyMQQMjQRsZCN88VA8oBWuJH5IiKK05KGl6dfl/Xny/ww35
mrVicNCleIlAZsnyiGY7ZaSLCotaSmsnMWf95uJpvAdaXC7aQa1kfWUp46tm5Ahy
KYVR90x3Z+3HSNZ09TLWP53lf3CZIdMMuo+m9H0UIEEDTZWzPI0tcagA7n6PoMWk
RFn+7wrxo+7dSUB+nET3FafLmNT7oJApWgHw5GEQlmDZ6Xz5nLLuc45bFlWN5ayR
Ft3znP4Of+pa7PScsJr1XsfFZO8Y5rCgL+CegPRG72LxZG+ctxzS+Gmxkm99cB7c
EJ67+VoKCM4c2j0Oef3rdmZ/xBHBPWhpWiHA3WdBHmLlap5x+lrv5qIkXO8XMS1e
PpFrKlhjX6IT/jDiFUiJ1MK6D/GsvWIYxNIvgvDLvdk7FeT8yiL7VwF+DlOUaPb6
xLSDa1S2bXIFQVwl1bbM3Zt3W8NnlfOEzOFlW6FIhZu7ifE39MWREGboLjRHJubY
NCB6SJiDekGu0KV6Fwxb1Oab9h+hD41FaWOM+ATXBJzZmiED+lh2zY0nzOSLMiQL
xOH/oVZlzR4zTap5KYUKc4r8SOT1bKpDPJBNziTDpR7D1Xr/+bc6OfHoSm42MDH6
9RVc+2kaKl4JCmJMGf08iGXwTEgWj6AKZISVY02IHvV3ebpgWzHdy/zohy2bwf6I
BBrVmEmF7rviAssFBkywIWIq7YTaciyzWm7DWL62J7ytGGbPDWiiBXCioEoGubVZ
DcdN8ztzozkrWHqKFIk/GdFOX38emQNZqKdMtrl5Z6Q7vSOwU//2/pjZuQwh5Xv0
0e4XFueZCp3Jh2AcUWayJn+rAOKJggHSAeQ+eNokCN3qxrd3d8I6T5rTNzINX63N
dTWwQDI5o+DsAWYN7ERI0UJkcq/3ElW+Vc9sAQsNltHetVhiZAa9lBihxUK75KSP
+MbmuIJGwNvTz+b/dVWYp93Ty/6jiMOH3PJODpTh4/4EWEJSWkR4MHLOC2TWybCS
jpEw7E8z0P5YY99rS/kAzhRnORkuuA/LAnRbwbKKraonA4i//l7m3/gjk0kzQjjy
ylwXJKSyRlMxKG0rzA3MBXgArLBuV5BvjLRaBz8qkRabtno2WbCsZYkEgXCRyj7u
j0O0Vi+bVvC0RwvF5lTZAyxiY7H6YbF8nZ4p2RhlEvMgpdP4vBibI8jBZassBn1O
U1wQ8nWBX8LfZ8XGs2aWQew5TFb95QHs+TcjJFZNGtZBLi5u+GNCLFEDBKAO2ix4
HrKGAGHHHw5Dg7pXfhsIMhRakaJxE0mbb28Q1W1FDM9cv+/UpVdhuvvXMND1rUoz
FdgeP2NbzH6KhuS2hEwYaHp8rylvaW7yIJZwiiyBV3iOsGXORq2aVT4qkAoCx5hL
4UIm6HBOw2ZpJnigodxSQJbVVpQgzc+E9vwdUOvrDRV2iPE9dAtip50yKpCHyOY+
NspmkQeykujy3BEUa01/H6vCgTKUu1NLgisOk+z302LjPjiLgvHD/kTchnmLLJd2
AEhY8Qm+Kal4EuleVJPDFxOlhF7Vk7LWcUBvpmhGedwmeg3sE079QgOX1Hg0792Q
f4i1OUPtPA0V8KAF0EVgu4P07/Kj2TwO9R+iU8zTpMvizOYjMxWf61g0gdt2Dbsm
PFbzuHmLjtlSiAp8a+RdTzWn60Y/PQkrwUqE8Y3D+rI2gX8tyQJtFDuJ4wDRtw45
MXSNmg82S86EUqACU8PxTO7L4lormWFlsS1pFZrl15OoesjT3F53DgHe+T01woLu
qw3IkkTbwTHOOk/J/xVaKWWCEj5ne23wXFONrRsWGV2vOR/ZMMokkt+PXk+EjOGE
2jiESyrRlFYIoq2kuLG5oUwgDrGXnpRWbMPAZzUuTIb3+6avpEwxXyKGSA5W3eeM
lZkzwWE7RfBpa9THGj2I5y34eCBv0QM2q6XNhVQHOu8nzL8ZmaXxyTZD0cQWr4b5
b6nCSL4+H2UN36iryNVN3c/+3d0kYve74XlIHhEdQxk97yqrIZWldpMU20klC5Ky
H+6rgWt54bmR2lGqvNLacMm3SlaaeGmWMaU8NIpcI7ON6V0aI/LEYZivNYUcPbpF
6nEnU1qmrR/v2TlwwOm8Psn/oQPY3TMF/MRuPfknyDev+kq++kLd6yLFBGT0DbJX
bsGLl6FWasHsISAh1NvakSI56x2sbWfjAtkg8HaVfbOl74YTaFkukFSBT65YCKVZ
A704GO9d9SoMo5T3gV0AOC8KwTn15Ho5aLlJ9pbD1jGZvX6WMsmFRd2mV9HcYB42
0+o8qQn7fU5NUT9URuzFEf81ULBr7vxH4yZ0zR0hkW9Gvs62xzCztpjNf77ug5ml
krsWK5VtVRPKVOGKmu/PWY+5q+2xF1cPR2JAVV3E3K0Fo9P8DqSdUpAFuTzgctJ/
kuNfIr5+4TIMadUsZhpcfE7mgNdXqNAum7Y80CG3aQ5qj4molB3zvI0mt24QOnhu
LWMszs5DY1ZC85+C1ZSluj4AYRI7clgsI3dHy4lFEfuZlZJ/PEnJjuLVvSQ3t1q6
yYMgLXTIS0CSoexy6Q3ObnyB+c2fgM5jVzAHoTycTXRV3S7MzK/WglbMeXVnw18/
CFkBogR9kIjRTRY3gOasCFZNSUbQZCXnAY8uc+kfsoVc1erTBtNhQtMK6QC2N1CD
2b4hPdvdFLcJCHkTAFDBPKnkTnE/ugFhYZ9dP5Lz3GFZB/5KC7n0FhFx3LehlTgE
4CJzvN9C7OCxwly8NTgGJndHJwKPng3zNn6U3T9ilptxfnKI0/vwvILPLsgGKMKe
ALXaBUFohL8f6e1O+EO/D6dneLGCMFIyss8IemySIF17dYJ8wN4cDv+2a1H6MKTZ
DWs7uF7fmLPeM7IEZqmfmRDgAck3C//0mD6FJZDif6ptXL9bx5rsXMLNBLJERTdh
7UUXAa+FnR8V4g+KbApbfjlrSvarkWUsSXlzgnofO9UcozlhpPGmewXRNwdK4fwm
hXgJ4Oexzt8iiw0kh47M85Qb9JVTgGWsSE32ZOj96tlsWNkhdETFwqbMUlI7haA7
aJPk0ISHYzIAy5PeZ0UsPu4p7BYClf++BWyMGf6Gp+T2x+g9Dj6GZqwgo2X+eEFz
XxoYl/C6gsVmkpSIL73dDnKZ6jMCRSMknBxPwa9N6pN/7cZ73sa7wJIi8z3Ri8b9
F/jbtWb29KPW9iulyUNipWLPaX6uugko/Gw/2m+pBjcKxpw+Fu3gPpu+3YlUiiwY
1lAAMmZkH8/SC/1RahQawduFOh2FyGfzhuCvAkLArtHSCmRT7P2qKWJVFa7EQW+j
94rt0+DxczeHjizS5bMo7dWasKxIY6mDvuBbRwTFGBlQajJZuIWOegYv4M0k7HnQ
sBgPgdnXLdpfsEDdlzk83gCJjT+OmS1+KIK4GSnSeYGC5r9wzzhZiLeuqt6VCH8X
e6qkMxPTo1VgS3d6cPq75rqSPhwE1EtnW7Qlbl98kWvrEduxjZsWcvhcp18JlClA
S3lQkAZ/hMX/kGgJBqfRy7au3sF6l7ULZVMNb/Mb1a16HqAQwby7PuH0t95AtQdj
7fp8YvIKZk9g4UjvxAD5LBOfpeaK/tluVFWV/J8KpNn+FU/4iH4y28IVMozwpRqe
aAG8a+Dt9eYo52N56/Pn76Yg3RtSC8TNwwKn/7Nfq7olXaU1aK0NRk2CY1/GqhGV
HsgOY0QR7EbK+tBrs5VxsDlmXUZnfbBm2Z7Vx8SHEB9KQhhaCEMXGQhHxmktbMP2
ki+zpClRyaUrxUFGd2lIsWJY5CQBuVFy6MS8AZKDvsQeDCZUQTlsR88Ac+/T4gKH
yP56XP4ZeFGe2fVwJew2RO+R7mAIa+nwrGVATJ84ij+e/l+8P26SagFhqFkaXa8H
odTR80o3MXJ/TTQAkSxEsthSQvZCDq4neC+Borte0Wx02UBtTGJKdXebV31mUGWC
D4qLs0C9qys+f9SaLXwoNpVKSKpRZ1dpqJp/Z9yOPDEqa6cVvZeYiUOwHNvNennG
vFD5woIyn7SH1w4XwSP4jqOKkmz7TUj6hR6geHQwNRxAFw8ndPOKc2RdEEvyd/WN
y72q+NFrLNpJmLUL1sV7Z78BoPzAsrqJFWEiskq9bTQgcuqRXx117pwkVtNEJ0y0
GFqRyX3skblmp7ciy4djAxIV0OpgcrcYILdChrI3/+tVjpMk7euvT1pQzbTY5g+0
yhXXAO+wzqDknCnx/F6C/16svIYnIdceQ7+gWgkoJgPWffi4LdC7FKfotI9jl+cy
Z5P7b9z5qbblO/xG0UCF72R0FvH5b9toPGIxc1CMoR+hndmeOtFFYQf61Rr3Qa+J
8TIgxKutg/qIFA2UR+5GGqtaCMTRiRrXrkjGXoqzTZ4ZwpHyJa5SWEAX0ySR4iUh
9UgSMsNK1gxSJCdMEO1qO2PI//Ncddt83HBN3wZWFqtkPxM2GePc3KnY7C3dZzhm
XYQ/fKB2xbtUc7jsq1TRVkeJhLBjp9GCXAM5J0NvK5p1mfrcWs3FwCvXT8SBNyOq
VKRrlWA+0sF8kjkY0puR9Or0aALNEpKal0q8GQtToZwa0vmf0N+CgcnE9tsz5hac
hIjrHHrZFVnX83OD9zg2rQTYwDYmtnsmhW4ymrXdfn5emHHLETsb+aAtY9OP+vEl
qvKB5vSOX6QvkCXUgHogiMyLJAj0BhXxra4aZQ4I7TWc27/G1i+bLlt6L+lK3ZQY
/p7ScqSMyG7hpQZQVhUbyFXz4fqcoQth9/jL98Eqt6zpMdwarCcbubCdHWlztGkY
U41pODrGySd/TpnnDLhEJQ2sWmcQD91xu+5rP8nBJbOj3ceOYQ4EoKfCWr6Tak5V
sWhZwEn6xeZRuVyH1NIiq4tC0s3QYADs94iGPPJUAY3brWiHy258TVBcBo2qpTz0
i2gUCDISPjuMVbsxFMCODn5tahZqWXsJbB9+HN3bkSa32xV7XJvh/58SSYnXH7xO
w06slMvMYcombOZ672BGo0oMcwuGVUrFf2mV92hrCGpkOjCVNiE7JS08Z7kKOny2
97IbRzuG7/2DHGlN01Ef5gmtOzql7NQhV2i05Qm+qUqIkt5nDfwzM0WIIcCP4y/S
dWWE04UWeB8WDU0CN7fP9SyF0dVNlAypDACjoyWgw7q+Iy2olEv6a0z2AP3eMoaa
7SrUuQF88eajnj9Hg+4p8MNRXK9OFHm2AQ+QcDBgiVPGkzGQc2if7YC0kTcxULX5
FogFNuLpg3C3lbzg6ds1V9p/HEEEZ9SnACQXNuKcHOXQiwB7SgZPN+WbhiDr3UYb
HBmMHH4YNeldtz4GkMDtDrowrp2uHalmvWS6Sk9f3JeNF5qm1KSrTRWYCNYH3kTx
5sY6k6NnWET+SOz40kBsCySWDm9Y+cZOOnOF9JILFLWHobG55vdGrFWnq0+pbzPL
itfTG70qggp3Sx3ccrMhlY/vYaSlh7W+KbhmJtDtc3draLfbCnaOyHdqwiZ4nDSJ
Ny294Kvsf/HUnhDeqwAugc30M7kzWPhD96NVFeaHGOgk+WGo5FxKBd4XiY4NRMFd
IywBvwjY4E/5OVEw+sZbVmeQtioHQtKQf5u/zGswC7ikC0wBrw57pRYXD3Cut0ml
XYnsEzW+DVs4EGLCynrjvoS4HONnmerMks+IPK1tgdlP+ANqNDQR7xyT5JYIdM8G
9s5yd2B6cgPhByL+ms2cQpLlVm3E2EC61xr9y7s9GoIwpP0lUrWutrehsrYG4+pY
Hf3zpkopxOQw9b8sei01ZSlxRd1aQDvbz/3M36VKLq21XgHEFp/CMjGVG0+khOWg
M4F8KSbt71XjE58zrSZNPBizrcDqmXw23sGgB8qMeFsBjvo017bf86KYJpgGU6Fu
1CqXLAGuCqxGpZlHwudt7Z+doZTmpQk9VqZVTM7t0sf1WT5f7aJ/HR8taSUC5SDM
gJcwV6L3pi8y+XydDAPA1lD3gSBaCI/bQhSjdQzikysTPBVwzM8SAtflVLRvTzrW
ae5YXfccbHRjVFGj3N7+6xJiIzTuMP4vH5J5y473rs216/FI3Ho+nqT4tkPniFQy
abbAZn4+OyYyaymvisFsxQ7DsYKOkAakZ+CotDsBf4nhFsdSuw1r4C8VYVLEHY65
pWPVGfmIfUQ6DkQJvPVtgdy93a+d7KZkCh66QkeI1gyrcStHQsh5Sku5dHDRk/n5
lLFIE3bHjfOIDrIXnc+RA5w/64DE1v78jzmwBMWkZc9h/QPhZCQrS0DGXuwl+0N3
F/czoEraycgp5rHMB5p/U/BKFX5j/4o3r4RnUEGb22wCTQFpbgVhueWGQWTPxhG1
0p1X5WV2v4ZapzEL2DwoWFdu8824k7Fif63FwyqNXx2NEVFOKokeVtSxyrsitKpg
Dkjw+AJtTPSYCjBAq9brcmlfJwrCPDjEgNIeqKqwaCk9PDhs7G0hXdXYG4brCp+l
as2FesrtpMSY0oCqEYSuYD2HM3YHuvFfxFH6FiVXbVkvBeXS1IL6ZscAd2EiYsDq
OmQcmqgcYtdJRirfVrmzICKtlqyRDZq5POiKkA1E+6Y81b7drQp/QUWVpHaCdi4S
KZXOa09JN13MhMAvC6IsSeEqz35qhnsV/OODzrMhxZ1Bp/HRTtXhZP76WU3duWGW
D3fKxkjEaxoX10UIgEmYKtMdcLFj8SOB7yp6KIL7ch0t87XsgBteYnllurSs17eE
i6joUQ0EkwkbOGcTNFcoIcEGHft9tpDcCRbS/31FHqf0athuLkDFxlW0oa50BP3g
pocQ1N2MXWxKrt6hXKgynXmzoZUXUqRN3VW3/vM0aV0Aqh8hz8J1/F1wTzn397sh
IlpoVfHAdCvTv+tSydDxQGcIjNvpZpZlcwCzhjA/8IswR9k18aZgkagSjvDL/PdV
QMZmDOFNEohZK69jzR7JuH3OiytNxyp7swa/iQPcuIS407FeRiMZ3UnAeJIHPP7S
jeTA8keSFdnH4O7bNeRAGDkM3pGQkdDoD+SYpmPqc0EgSw8dedAJZ8MhJ5+C1kt/
I7hBUg+y5msKi7AY6h5FLglPnb8s1eatXIOGJyw6Hal4B+7/OSp5p56NnVOGHtU8
EAofFSK1spPHn122mRBd/yHyHjkSgADxd6KHnGk+oiljuMvQFNgURoVcYDaqJJNY
bxL3nC5I0chKaGP7Va+mDMNhn5WUYDO753gveJGGGBnVkeLMw27fOw61q05qqp0L
/turK8ryQZ00VpOOUP5XN65ZAQPj7M/AxGfzulPLgOA7uG5XZXSD+edrX3wBbs31
H9tvytv0p1CPiKCydeYb8+lSFl4eZ7q07lPAd6Xp7g9uJUcsTuwkmJ/XJtkDEMGg
hfmKee4JTuIICJx4BIPquzabosPdR+fdAhJUEI9YqVH8m4d14ss1zFQS9wAwSjPg
cyVhXarL8KFxVrctDW2lNJHQcZ1ufMfHC7Mi7bSpGVqqM8kXAWyYrL/o8DdYamVg
y7Hh8ofGsl4ubTbRQxwewY3bFEHxprvFKYrUmrl/xPjlaV0t678hrlH+R808LJMh
bLmO/p3fjYAVBlEjhRWOW191fIb6Q9ek+iCgH2oV4HN2Leaq/cxEVmHG1paNxrdV
+3KwpN0QfbbApv9LkweNZ51WjznkGYCftMGr4XdmlcdFxfejRZzE3CaENiOWFU0I
WHiXBaO5z91V9dTAfYU5LONt6foWAp+0QC26I5Bjhbh84rcZWdLqM+bITiWH3QJI
VJjX+z3pafdkS/glOjh48HY9dz9hkN2RlZwImXtYSidQcSACaIKz7uv7WlJAYSRV
B6oWXtqdposXrSKGPSk2sECCI/tn2mIFq2cElW/KqBmq+9EwQ4/ees30G4FTY7wY
bwrYGOkirSSCKXqXtZ2YvPChk0higDEsJ5aE6nhkmHioRfoDW03bjqac1PM05ypZ
xNt9YlC7vn5BTdLPGi8wqlB2Qthk9IsTABUA7fN/8UGv9xUcIqx0zhq+r9e+82j+
g1N4lleB4+o007AF/7aRlzTyXjyxoVG1dPZzi/v1/Fai51QJ2Mn6z85u4LL53RRP
NcoGu1QRsE9yUOoMKJWJYGJc3L78IkC6n8fPsnAJ/uBtXQyn3TPQ88eFGMi7IkB/
Ywx3PL8UfKQf20DKTdNjXyGjLOUHyI6GqJhlYi2KOHwmoGHSnN7B9cER/s7nm3xq
n5zshBeUAWdGb1SjqMtHNkfLSKkhRiD05b0vUNklgMGvPPiWPAhLgNd4srZxRikp
idOmB/iLaBw5pulfzPW8StstsSLY61yOD3IDlmxJ44cVBASXgqfpP2U4hM+1eWaW
xDZVlWrMKYuxOdZYKl0txl1Qb3m86XJeqcni5+rNfXIiB3e/h7t5b5xjBTjlxyE2
TfGU60eeSLCYxTQnJ3Z+/IfLL4sbDc/U0K7i4lrBRIs7y+RB9fZTR400GlFAM9zs
GHL3ej10AJZglaWsodqOkgDWHHmLey5LOeIa0WKMtaZqWtpRTnGkMd47kRz+Nu2T
22XKzTeizc94bpLpoKiGtDgzF95WBRmXng/fpCJPYygvBkyGhh4QGJW77CHl2YnD
gQmEaeR8vqSpmlG/XW/AqBX5zRzvjDXBkA/f4land7QJ4hIPXD7U3x6Gd2FklLlp
ZLD+jtFI5oq7BJWM9qneyUCKczvlVWRyN/ahxdf0Iq9I9V9VFhCbAQcTMjZCz7DZ
CQ3NbmcAOT6g/PcrtAGMmT/VoBUzLaiQjDzmrFHDXzDKHA7ZqOteVou4IBZeu41q
Z1JRGVyW2f12ZAUbhnCkFQyTZakYvZ5+W9MZLr1N5yBQ4wzyo7eLXl3dccCKGxQM
OxcLLWupIS98FGnhozFuX/tzPBX+zWlT8qo3j8HRW8G+MId1UcGDZTRSR2QPB+Q+
QLhO2FIIkZh44XUw9oO6xmz31f4K3A4pruIMERDuaFIC4xUp8TwivLPsmT8I9Yvp
YYOoStxMWsJgz1w9rgq4V4DPro9el2XMXf/Fbb/cetoFvx8sHbQVjrzMkQu6XJhl
tpJPh0vKKgIyC3XRfrYUxZMIzGcoUlTsri5MBDu6MeZsDhoUy5B2owM/iWIUxYjT
g4YaBHoXaTt7iGy6BOd8TaTjrsY3q8yviPC30bHbuTZUkY7VfHVRinqbF2dR+/Fl
ChWEAgH4ZQMyyj0bVSYoxrFgwkZY93F4NEVZ4qtrqA4Gn35TokgLh/BKojz5uio6
rqswFAFt4dRMXSMRQ4yp3oszFo7/uDKGtREUZFLwACK8ygZ8UoE0oZqz31D2RovU
3lTwCWuFGYytjJDtK5U3lceQOYLNmzTD8hExRKAMwH+L+1rb5h1rTC31vef1LUkz
2UUrTu9y+vPiHEiS5QvwDDIvXQcmiaR26kZ/KygWUBmsgPYHCTgHJlCbgcISmnRE
+tYwmEYuetSeGQPoRLFbAW9llLen2s5Yr1SmmWQLs8UJxwZc6mmJeV/AKP1MHFcU
3fhRdtrzoFdaZdAlU61Y4As7mSCysG79Ec8ndQvoQXx8CPvjs1MGqWy2iiCE/NJS
LgGhJPODESNVlXEL77OSXPzwpO40u1Gq8QBeM3gC48GEfASl3GFFb2/hLIRASYNS
+qDvDEEWcpEDKySEmp0yEmeW6VPOOJwrUlYSvYsiX65ql0tx1bFFIT3nbZns4Q1l
/GW1zi1vFAwygC/cA7YngwLwfxn9g2H/8lWXLq9xt1qU59bEgtAjCSH0SPfV/sOn
tfousx2LJlvh8SsSTF7GSnhegSBT93Xdo4PSyuLuHzeTLNczm16M7FoeVa9mwdoM
fEvLK47I3gWchyWyloGW/J7tyTnoln+sGHGZXfDpGnZOhQQ1buXKOynOkyp+fQFa
0Gl0BbbGv/gu9nCQMAlbkTKRefZscWMGySnSGe45ha3GaFzN/qepa8Eo32F4qEVL
pDgkL1r1EdzULa10ztsJ/eXv9ssPGNB9eHMASlNUvcXyLIYIVqn56SGbR3KDwpHu
49BAYo2TOQLxbr24DXEBWwe/+aq/n4cBMYf+uXdRIIowI1FMK7jtry13IbYmBSs+
tv1Hb0pBS+632EcNRAsEIF/LDUsXoWbqgsfdMC4/VLEwcmoALscWZwOtY3elt0rF
M7nYEULNZhCvFkRk+IPtYBeXQKgz1XS1wfy9rx+diOMPoQWwTje33GjavDqSaPlP
FEz4xyWphjiERrhfng0PpJ4JMHWDYN5qhkZLUhCUII2Xf0KzWue2mewIxwvv+Zo9
E6yqOKGd7SET5O+wNkPc2IhyzemXCx3H4Wa5c+D2VnaJgIJ4R3WuNkG+trUycFYL
Pm8uCC3M6LYKTG/CZHve2U0zb8f15ljWYJgZ62jp7VvRN1xF4VQy41fIByqLT3z2
eKL/pBqGbaIcKl9G5Y9OO8a52mUi9y6cP3gGFasRj3ZOkhLAf02zZG4c/CnqaQrl
xqFdUOUfjMBdVR2rToSD0foxd56RgkjRbWNIKYmzt2sgqkgbifjMdQk7+pIqPE4U
R0GmENT7r9853kVn81Qt6awdtIiHiPQ6OzPH3bTG9cc9hfjjt17RlDut+SR/0NOf
d/LtWgbgj9L8P5g5VCkHZLg5A9Jm8cV1La/ZOay3UlSYhY2sTdvFspajTj5TiA3o
F88KrlzB2Tc9O2udFDt53fad6Bo5ZWfIbq1AHqxsOs/gsDa4wdBtoNdkSuv3naFX
076A1PrWEPJTt9RH5wkjl8dfTjiwAn0KnrgJpFtcXmiZ8NHWC2atJ/yCFQqTRdT+
ULr+O3IQ9r0Kbsg2a3zz8iwYlb53ZKX2chkGZqAwTaRzaYKHtFQjO9ofi27vK4ff
2A9+bMLFpazax2wHBEa0t97lljkmLG0DuRGL30IRa0Xr0pteqXyFqel5ie3kIFHf
974hMYoAoxrsGLLW6QhmU1WNRqGHLdPnlOHbPNwKzbfe6CC1HJtkiI3b8QYWxPv7
GZnEoGutvz8cEldqUbesU7uqX0VsliGlJK0afuQ5XnKuEaLr08/bubiaP4tDhmSs
Tq/CICm2Efn22gp1tkMG2DnFEYFuc1ZgIqdGDUCgUOsh9Wjl9Ly+QKf61PiaSC/t
noogq8a+XQfbik2fnSFEHqFFYTMTnoS0l8VI/6hMoIhJlTD9Qdvn8fXI/ZG4sxFD
oq37oI9yDgalle6BCrSk0pcn9pN0toEw7OtzPJB0Uco/p3R71U53h7dOjvxH7nUP
BaRY93B4/EB5e35YEjdxyHix3IoFoITsLanBXGMTJkJLKa3hDdszEHDsW02+Rfk5
xMRJM1Ra+KEEdEZRizvYQVU2J54lmBWHjNxLWXN67ItGEjsfN9zIYtIeOQ4l0rv7
AiRgof22joYuRlLf6i6leOferPRn1SjCfOHbyK2amvrnh+z+8q8KDhtYP3c75bcv
UJ8RCI8sFBPqzxH4lQwQdIlTlZDNbCLIqlw8SV5oiLRhgx6MnIiU0cNKHbeJTZP+
zZeq4MoWhwCmBI7YsgqCsZXmNNZRTqLc0tgx3DvbARWPqiisrO+4cYLDCJiHyXDI
8Pa+KobF0mM42V+DppDJkN8iYtVCr4dEDiee3zNlyga8C0AQphmFNkk0eKm3uz7C
/FH3HFIlZ5nEn50hSMCQ79Mdfg5bqlrgCXL/YlAvfRY9mVhCcIQTSMi97V9chGZj
NyFLDW8HBJDudPhAMy6PcX31ldIO+kjDwTO4uhHEPid+OMoIReeRaKF8R4G6pEi0
f38ulp0l57KIFlMV4Tuf2fQf9aTubvO7eKH1KWRygp35mUIcKZ/kQ/bltlroXUxX
IFbhFAmU63WR+5VJ7FKuKETr/q+873fsAJYFB2I7riopic2ejECUXAiG45bFI8qM
YLp+TtoObSDTOFRn6TnCTzRf8EQKxoIrtw5jBLlDtMdb+vzCy4MHNM5MEWeae069
+QxdZEA2zV69gaHMSnV0A175FJCHST+a5X89ZxCs8tW0bL3/TVhz7JbiHzzfZrSb
d5CtzVzq/9Dr0v5Up/rjnMBDlmMqC4LnrChASplKWoL7E+SkCELNlgOMcKfIEn7X
xsT+f60cAfvCxKk3gxKE1eXMdXr9JqERHCUcYkMhFfKVUAEMwFDRG2ojrBW8PDIk
ccfrT8dYqYJMJE3WQt6u+Q3wwcsh1T0beqt+LQv52z7w9Nnm1FhJnlkDyR1YcZcb
cum6OmTbbC2CJkwc5OWkvxb2Y4RHp/m+qhZDaveupinS/F3+8dAzme9WAZOg5zqN
Skwy4NqaMPs6DfdIrUrb/CvuuZ/bHipwQ4QTwqXFJnZwEbA16iWygEvuF5BMDWxS
hHlToilRpcknKJhUMf/PvaC+RaaPeVMuS8/Npp8zHos6swDyPGxXEN8mbLsTKZO+
dzx269OkvNIX0UQ6PYtgKY6OoLgW1kfN1JYfFm8hUM+oJgQKiqZhrhNxARGe42un
suSxof/jxexJzb0OMj28gZOvewvChl32U0XhKz3qemJVBnd4Iy+nnMPCAtz2/kFM
oPF6Elm4Ukm32WkGBK1eUlz3cGavrEci/BlB7CNcEN4vWMH/nIl9oNfH2Fqyhzy2
ky8f3ta/gyvO5XU1nWfQXsNT6ZZk4nqdqquPM/cP+nitE/gUZyRPiHb9gLW4qG9O
bTgvX4AQt5If2RdNuAd9fxMYxml8D75uDTjatH+UGwvVXN3eAvbO8QPuUCqJ1yLk
7VUB2JWompIThARc70QDsNyi4ogtl7tdDYec5/AXIWGiZ6LK1ACrTb4wM0DfGqDx
hn1kvwHIHVipqP67SdenzeOKKjkDuQWw4zHXBYNtioG7olm/ce24pQOdW5PSCPWt
HPTV1pakFV+U8oHaflzLnEtiq7otyqWQCJAS0mecO9NUu5nT5yByR/GwE0ospJBR
P00ylistuRiB5dWyDgktkR83T5YSEMOgYWk+UAbNT3J+iQm0YpBOa07reD1GAkJb
5pcCMPQ0cZVDodABA+1DMXj8u677+CcMrimmDz94iYhrPn4JLIy7JRfMneM9lCq/
Jf3qTqOBbR5D7ZUvW/50udhGJbZ9GODjS9TJMU8jR2V4FWWEpQkux5/npYJSbShm
cEvUPBm1h1Ol8uzsCWvcuiaCB/S1Hk86j+6o5J/RgVJ/6ofYxtwUsanEMFFvpNL5
q+xdtW/j/aP7HaoeYSPhPFxVdQXStG9T502irKtdGs554fcj9aRvvh9G8xR01yYG
SD/DiA/ms6Vb3qqc/ALjoef7BlL6bzRmCPt4uf5fUHMbfgm9e1TLPdD6SAFNb+oD
kBcVndv3fVOKW+6DHshk7vvej0/YH1Ui8EoKzVtoSJw0DZ3FaNxE49iznIuaSWUg
dijkzsFmtqw8jRXxzQOxwBQErchrL8zogSl573CeJEVfCf9oxQgaEVjV44JE+vlD
JLd0pnPrG3JSPOcvzjDD2d415lsv/nqmluY9z4fxnTZMsWSEUKHYzCLr2xon+/r1
QUfL96Jj87hpRHACw1NqAkci2Ne4tDyIo++ElJXvNe3oGKCeg+e8uESRjDW9ukWD
jmh3ZjPbVx+00ekFp1LYcoRshOHm5YmiNrgX2i0/svcECJvDhuJEFA5GnEHIGtZF
ta1w+Kobyi9Ax1S9mdLIR/hGpI9qa0P6tTAAPpza69vFNC+taogbj/Y0eT5+BelV
j2vS8tXpuTPvD5qqqCNixVv96DBpNg+sBHHU0tvTvFo1zBIIc9nPkiOMXOirCmzO
/OwSosD0nQ9pB2DdCcpw/FIH4AMnB9nI4VszW2Y+ITAq76eoKeCGjIx/Xv0oCaJA
49a2ZbS8GWONBK5DpU6IhLeOzQi2JW4fHUX/UtV7s8NvkVEPlJzV3+L5fShzdcGO
g2ayrDzvg+Om1rQlMmrWtg0vXhqzi2ytxku4Jo0evJVlWTyzEk7HcsOnSP2SAGIw
YLR3fpBKWLteIPrKfoKZy9xaBP6jS0UkGPAE4wmqxhklGCyG1/SIOYmOsDVG6nLm
IF0aAn7nXMnviob/NFm7Z61BJq3Ww8yIsi1R1S0QRKrM9PomYhl7YxIw9Y3C59Fw
B/sKsnGPG3Xw9v40FuBXreSI8ETFSanUXL2yuuBpAXpTseBe5z7fXIZosq5PHVDq
rb9wH/HiIcyT9mzn6h9DVqqrm8GS74pqMDX/1Z7JIRUpBKraSDfeX+bs10Fs+mVd
yKeeLHQNjvgbxduhkOOid/lNojnLFbgwedNZu6DaoJwsmnIHpOnfzg9zpSXX+QXG
kKlbv3EFm1M9w3bFcxP3EXFeAfy6Am6LnqgKVqIdlEzYAubK5vSTqgdhWFhf2H+W
d2mv3ALoa39t5gQm10ZPHyjej90r/WKAO6tRaCtkC4aQbPStQ7qkO3MSvc//EgT/
NWxNET4yhY1JsoMo3zF7SuPZRZ2/KgqrUOxHeUbgQdvFhOIQXQ1GiUUeuvMkxZWB
fo536H3ZZPzjJC5iHljAV6x4JtYs2x5gibC/QcyWQfoJoJn/rS7zN3T/SdisUaV/
o3UHT7Zqis3FNAVr/M0RCr+yNKEqpffheiFtvhnwsD6t4LVnLfRAjRQk7rdc3OPQ
Hbo+OWrt5iwUgtmN28exHEQEFYKFk7+TEuw8qmWJc+rvExMaK9nmKZi8j9n3S3vC
+V1aavEHAyeCb8VOcEQNDyE3bQuFarHN8XDTA2Zq6+k+xsLcBZ/NaT71FMjg2pW8
VL8rFmQmbU4awgvUjhbSo88Qdu5FoviNTa8nNXMmmJJGkyd1+mt3IYLJM1fa+ElW
DvmGMq7Kgdn6oz/GJHcSF71ubsfH3/yOIqLaw7t1O3Php99OD60GoYY3hLeSt+uB
C2e9tgJBy7CNckgeM84SWmP+6oiMYdKOjYI06B/EAtBbhX8fzTBe2jyUeDN1sCMA
a2FnSi6JfLtdvr7Vt83c8VtKskzxyXEaJZUfLG5xxbpgJxvNYutxOms3FMMxIkLY
4oZ9Xu5b3TyUr5CVBPx9W/BFauk0kaO+4I50rqaR3iK0NkybSV0qxj2M6BLk4nwB
gQ10Wkl3FuomRh3PDnECEW1AP69PTAmW3KhgPD+0WJXLMmwmNqXWXxpNcCCXsX6R
9cyZld/nYjTTztCnzyHnxocSHZ3UMHI/GCXl/dTRfHy3RPTGcDQBvCAnd0ulEdb8
pQvEjfbdHDBNQlHI2Dg6g8bn7JpQNCIEX0CK8/J9M/TZwHtPjUTfBDLGG3OPYsoo
MwSXcigyJqZZJd66kY+StuIZE8C/8f+C2t9cb/bWdXEdHDG4WmBuKPDkoDCjgaGT
m7NiEzYUIvqNDSSOSsYKnkTwy7xLN23apSjRru+Pv3YZHdOtnfCVCAZNwj/yDN2+
jzBzE1QRqvP+tJWpPpZKziqOQCyB87cMh+4lmgFp7iEO4JL2bDndJBSBVLusEJze
UNwRmfO7gHzWEtpIgrMpjwiPb9dAz+smck4GJMCybEHY3HtT0WlMlFuSyl1m1whD
8xmZIKefHs30n1XjHPWEYxZUuMVBW0L4l3Mz4RloZlAI09phU7R/d/KVsyZ5n5Ii
g5icsVRFLNujXWrzlwdaVLaryzzTw8vA2HgDQvAZEvAUd27LNMnWDQwM183LRZHC
9SWkWZYdVv5MSeDp1Fc8OLOLlIyeQ2gdswAhZRQK8smOoPxVL0/iG0Qn/qwUzQg/
8a1eUsWnj29dBlVoLJo3yO5pPnXLft3tQ428s0/zG62fspnphcvnVXmDr/kfwY4s
tv2ip42ulvKZowGI+sQmGuQPVkHaEwiu6EzRXoesO2OL/7xrM10ko5Jn84yKYj0d
wvZ+h65OFZ0r931rrPUY1KKM+gvVgvDfaep/U+2pYbPGephPBzGPrcUGclN1WElt
GmLtyg7qZrJ2G7melcjPVUK4seamAat7jf3CI9j3+gZM0f2/0v6Kkm0OQokN8YJ5
wPWQD5y8uxDTxoakgk/PufBM4zR68k8PqLhZU6Ymb/wroAHyYgRnaGmYffKCKAq9
JT2X9dBGoHBM4FLNOwWSPv/tCqNcqNW67Yw00UWnjOAIidlMgO6l82jtW3FRS3B/
PPlMoPkVsX/WIVT7RHi4iFohZDPi4XLstKK0mC8Qx6nQO57obJx7JsJ+ZfiKw7CJ
QtIKks+A8dNGjcFeRp69t7xVZ+7N5jh5rXgeM/1bx104tYm0LoFmYvAa2CB0jZrw
+2NWfmOkbTfhQ27hCLvhDBQyDtZGvgUQ9Qz2+h0AH7ztU3/KpFf1TwIF2UPnACBl
TCf3zy7nP959pF+ZNblaud5wlOvJMzr2SL1RLQpXGOePAdLjPeQiqYcrMZodtSUQ
CX2c1dicpJD84Ljm+xhB1mEF3wDbbLRvR68N4+JRtxvgadfUAtVZO3DRgtO3d7K0
td8SYy5XtsZgCVf5C5YkzqiDWe0zavRfJqpvuJPHNE9KejZw6mxgZDq45O6OdO73
5ujcn3D/5ZMVvAQmiZd44vJq5tPe+wxBKMFOMDAsnlF8WA+hFL3Zag4DJmrVALTD
3igwa2S8qWS+PobMr4D73ZIjMdnL/FacfchbixHR0BbfL3tkD+ks0C+/r6RqcfIr
TEUMWNjK1c4ZXrA1E+0ywz2LdrXxbZ2sXzpFHv2UlIjsBwzYJFXzkz1vJ8nmCprX
Fu/VgJtx8c4TOlvQUuTGymGmvw2H/1vEwTwxU7aRAonhc05+Xye0Dr2+lSktoxAj
XF3FrXlGqkU0gL2gDsxkRaXR8J2HS+L4ke3J4kLepJPwgFRGNwU0kr8KRBGQx5BC
CdFum7N6Wbytfa6een+7xe+KRerjKOT/uifD7Otw5nqIxhjGasc3ouBnjGx5oSVm
HhRZB9lseKqPHULudAo0fx+kul5VwM8lOBqj3OoyAP0dPddMhmYwh6hPeuojhQRk
yBswuiLhkBvSD4vc/342eICwGsxVJEqFOp195VHYCJ2bzhlt5qDxSLUwI2FwiBhf
xDN/Gh8FqypsODhWtlwGiU/eCiUNM9gDcv9EJQMxUT9wZG/TO4vCC5QRe4KPO7Cb
/sBCVYz72PyA5Qjd45P1ZjxSXQqUTB+oIwUf4hqLRM1rK3sNie3vCPwKgYomp5Ar
FIykx08+yyFmpvgofz4Kb/UBpCHSwQ/zfQuqZStr19XAHjo9LXbDu7ERkLjEW0XO
qLJ2Ak6jZ0dLHDk5w7rb1pJE9zCkkX7U1j0ZGTJ8sIogymBdUgCMhd3mS0CAS3gs
Y7a421pSAHS4T+Hp1mDpzGt/8Wg4P3jWxNnFSkgR0hBN0sGmUv2150EjoJsPc86y
PROmxJYNsK4LHzqqBW41fduJFx2sy5MrZ8C+0Av9XQxfwyDLJBPXprkVmjMZc9GN
K6MtF3txI/JGHFA3jBNvstPY+VaRpFDPBaQFKNgvkXPX1Fa7ceXYY5bgwxhjYME+
4WFElLg+5ltaiBJRXffb+StKh9NFxT1dxZ1m6IRYMgoo5jnT3GX2ZLxcXEmZUpqV
90YlWG1rb9RnjCa0INLNZOeMcELsjS7RkP5qx6JhFfrAO8bHu3pqycBEP2cRcYlu
2SaNDCMzviTTX/e3CR3e0ifLuiostM9086JduALkt3zgDa1WkyuMBNa2OiyNKscJ
yC4MIrv6ZbM7qcJcxx1JtcXL2fJwUqUug3gGbzQOCYv1IxROJUl/Ycs6ZPFIxUHE
W64NtjidDxOetA53ATCrKBSuTYyKkLfug65gVZdydGaq53xbLb0WyFpQqgmHGU3S
q1IweS+MxRST8VfOloLaso/I0gLha5RrH9w5qhcFqtv4rtYrCjtRcuoyUN6zxCG4
XFtWHLUQv5Xrw8NIm22c9XqzeVQJ/WKpwNlcW/lPJE8ESFWZkgajNhZYxHJziC6D
2dJXcRmQCwfBfbSacZtDLlQOjqWob0ubXc0XfiQEzneVomuj9tP8RtebOC5t29AV
MTr/uE3eJrCeR1da4gOqJwqPifp0tQyudO3w3WNNZ3ud3zVZwLQEuW3IekSHM2eN
Z7tBVAF7gqfxNWr3m+l69oKDTA0OiH2FQkNaMPs/Cr2pssRv8jelMS1fCjTPJgTJ
im8Dg2YOmV7Zpsbi0pNxGSPFtOsSViE0+8EGPi9IOU7R6YFtsA6fu8keweb9FPc6
q4bVfywSkA59ZEGd3AirV3uCNQeDh1aAxZNwW3tFoIW+UQ9ak6fEAF6eXxI7big7
YJpe18nSyHk1S9UQD1vlATP2WpKiwHCLvcoG83B986Iq76EzeNQ8PglvgJJhYgiQ
Do9cT+cVuuFWv5GZ5oyrV6Bre6rS2+rqiLZZ8N1BL5ORvQ7pRJqk/6bM7e629FfE
5ddHhY1YWjvhWhvMGZ0SyuZxHHgUnMA89JnUkS1iif5MK2iOIOq0lO+Ov4QHHnHa
TCwnNDGKv/IE9y22ykpnHSo0RmA5BmOgr8YJkSJQ80LIokCJSZEpPixIX+6mL79E
MB9eR0WsN1OxjXsALLRJg3QUcC4Tczn26OMbzjFNbMUY8HiH9OrimqwGcNXeijfN
KLwEyw4cvKccdfVdgVBbaZo8UGxF/khPAy1CQozEf7uR9ACUGJ/TXI+J9msyAZPj
nAfqwbweNOzw6qXu6aACE0fPgUgKrSw+HdOVcH9gK23SU4pnqfCyANDlSsvN1A2G
fOIRDJeRd44MDmnv8Zb6E5ErR7+JkQKsxn3/7zEjZpgHegl+bB/HyvlTNiQDQ/SY
H9nl1nGqF2+H9tuBP434Rxhw/j5Vr/cJF3LVfKdWanGuX6YsqiPvSg6192tQzFgo
cV8dRg7FWhHu/jQY/ReNjMAfVND63jgsesEXD4oZRjtNVYvWat82xsJDc0kDdcEG
FP5W2jLytrTdWInw6Fu3FKDU2UCj9tBO/A97pXTdnxf3coTZ0m+w/RiRJZE4E4H8
Ir6PAKuevmCr4yzzcx4AAP4fU9FdB+u0GGP99X9b7njREWpnyWmhCt0KYSyGpfp1
CJp9w8qTCB1jk2EoUbGJFCryPmXBR7rzbrOXkprh5g7x6ScRb2Z0hNLXv5mR0G/h
1tB5jl0Mrox4DMNeai90X0m8C5V3BXLpxQigcfb3SjBibQRmgb41ym0sB3ZenZpl
du56v1xa3pq1MzNZLTi10FLWhvsLLWeFqk6p8cF7pHhXJ6K5U58DVRPzllzSat+2
BAuPMNjShtg+gey3lGlUFqX9mx5R19QgkqnH8giXZicHReoXJwoa5QsTSQHcaaxo
5EMIaaY+a8n1AVgN1ANefQqXsTKTHyEtTYAEdXgvIfnPCfsfRBVxOfJST+PANeWg
/JBBpvkJZDgymIbLax/Ln0woWn31zPiV2aACho4ls4iCEjuHblI8cigiiARyrruH
4X6ek6c8sMFCmq4JI07/8yPVn0XmbJu7lVD7G9FbxyUpOKdfDLhTo1gvH1dOItiL
SdTeZ6etKe4es748Upt+13HMZNlAtBSMZf6gikKTpHAOV5RdREDx7HGNHnxpR/Ib
knekU1Z74No5yu3r0TCJcr05mmt6ZQlUQIGu0L+zQGydLXz7W7C8enZKAP0D7h+H
eqWxs0D1c1Eb5/eWCvQIKYuhUdFyjtjXqXPgF213BFl9Of7fmno7RPph8Gv+av95
AxlyAosv/I5+ay3dpk9Q8SlgbzYiUL8uJU7iQRu7KXzc/K2+ngP2Jff7ZWzLLTOw
HLGS0zdoKdOk1py7d456eB0YCsgLUv1lcSW5fsqwrnZ1G53ufF3ed47rGEH7Xgeb
rhzygA+uZOXVBRFr/7jskiyw4YH7DT1crFYbDoTkkrKYoivZkC2l5jmNEvHK0CR0
zzMJOOdka+yBxjiEFRDCCSAyrWRd1136EujwRTF1jLCxip39fG9mMOxNXuhDQcWK
YhhKHqsfxw2kk8eVJvqDghjmsLiLsdFqRsgBwWT8pSGG977S4nAk94KlqDMjSsD0
w/jKU4E8yDzzaZHoyh/Mz9K8mAFilD6m6/if9r/7HV30/wao8hQbJaUPIzycxnNk
AShIaTkBjjAflG+JmoJEhNJ+BB58i9MrPqVK8bmM3AsWbyzLWq39GRp83fM4vOey
7GAhmhUr5vz3CSMBaqNoQLegOnI2HlOESRfs6IY59Oeervlp7L8EqXwE+ei/G2ny
A+mC4N2otVAjNvvGbnea6UMvjU5NJs145Pf9fmdo/OKkLskNofuYddI3Erb+Fidz
sOfApoWtDP5BJfs9d52tjBYdDLYB7/HdRqZmRWaQ6/wm5RmoyyxKTOVZysAfRBSC
35EvQ7c/wR+3u/sqQiYffKZt6m3mGSPBpIvrZSXOZx7nojqWBykpraycsmADZB+C
ivyzKREP/z/CvYuEYcThp/LW03wGvmOJz6V+v6SnsKZ6W8CS3UPccNepHfDubBDz
lt8rtAzK459f17VxMZwZr3FvNb9/zGyDbfZVXKg4n8e7ggZ0RHdy217xI6Ce9d4d
tctyjxXGTyAeyX3SUtV8hs0fNhcJZ40GjpuGL9ClrQ2zKVojvo3KxVLgZ1BJfR0+
HqKTrGaRFVn3Q2C9BKgyf9+ur+3WNalalOfiju1F7Q2LyXddWOY25U4xC2QQwg1L
uf0FX/bM1nBVfZeNQBo1/fvGn1n66d2/FL8vsOuwCZC/3q6okFqrA32EfD8RDvP3
KREuS2mnTKsfd7yJPYWRNpkAEScYPQX2AOBWXjOEefcpJ8Rx6GEuEGbP31sOKojo
gaoNVTu2F871EKnCA27qESHg16yT+iUrvGeHJu7xKmhuqekawnij9TnPzsL65mue
pve4ujpru/LP0g1zrMFD+VPBUTptA+QKbViuGcRNHiTCxI40/Ml9TYb0l0RwWHcW
svwDeaHWfsquYD7W9fBl0jlON7JvFJLIExXJZSFXMv8Uph6Er1TrKrURBKjaRfd8
MifHQDI9iERAZ0MQsIL1H12G4BY5aqPtFGFCKcjKzu25+m52Lcsxb0Qws+rsCIN7
wsaCkppULuo5lQyJbuo21+3RLFX2T6HPhHVo4l9NR17ykKJVY/oOvnqQPjyfBmw7
HXt4Z8U0A9pIo52cnlH3xMIAMrl1pBhpJ1ck2PloOP0FtM0xKQs2umqd+QIcSBTs
+MqsnwD9OIL7I0j1ZwVlvs71PDwOKyTXneT+SKAdTKycj+ggi+P3yBGzwUuazMMn
gbe4FfEwzkKNM3qqBuU6tmru+a+Ye0rYgCHlovWRnp07Juz850VMvKxNhxbrekem
0tDGS0JgM/mvycDfWxBDnoYVwJxEUIg34Q2ar1fEwbsYuCZEyoMQid1ChbUskwmX
6ujPpFsw3fPU1kW4L0/OpWqtyiuzRbyjFTztAjL/0hCWbexWkGAqV6/ywYC+IWGb
xrmH/GAPBr45710LZgJwrc/wSK4qa1xTT5W0vlw5VBZxTEyuxXzknbhPjXfg7+cF
5YSJRkMxx84c77MnMC4aF1faD2TRNRPv6brjuxBxouAWo2kMDcTIHO5C7k69bXyG
dJm6+suIf79SbKpYuDaxihP4AZi2jQxk1AcgdLMs5ECPgqZvGxRib548vKs+kieB
bN8ODDIUjvNqsesG5UsDB66HIgWdU33Xc0vN7+Lp45FySkcTDhM8yGsJT5kRgDoZ
ZFcJljoB82+gPwJDw4t27kZuaI1ZKpnoujdJ4U1p/44R4JcgyWYgwrNg+qN63oHB
E2CyshofppIS+MYEnKgUr5psItIUioV8p9E1bUxh6eOsT5P6YDo8gl4o2gD23Nv6
DGrCGGaEJHwNmzhBefOL2zyIrX47rEuZwmE3Yrt21mobHmQfsvpajEi73/AH3r70
8tZa6BvSwYuibiv8SDu9yrccHRjUud75o6HkoGiga+brj6/m4abZ2DoFvI9bpntR
gXBZ/BU3bsgRIcxGl3Vz1aCvxFAtiD+j5/ZrepknOH7CMyI9nE1XHTk3Cw7pehZg
8GX9+3etk9Z48kbBPG1fXC6IS8tA/+at2L+oVms6Oy1jR/TBhHj1Kq7rBMebsu//
ranIvTdeIhzS+CV2JCWK46XNz58TYuQwSyN2zo/D2mfwWuiOH7zen6g3FYh0op5c
elrttowWjEa1QG1orPZkZU6X+E8+yMWYMRi5MMcoPPmVPS5YzrscMnQ+VPU2MXBZ
+vQzTVTL3akkKPStDKNo7r9uZCA2H8IN3xeJEqZEqGDzIyMcW/pDItZeFnU9V8+S
dgv06pE39Cz+B96CICzYj40Frcwr7hI8zs1qRJtbUgDdJQc2zR/N6i34a8m9qYPc
PXyqpG++1kbpSRniKTHfJrjg+RWQ0Ansn5SND8EvXJCnQAoaiD4EoWAsUyqVD68z
KIHveMOR5o3AH9IoJ6vL7Emt3Yl77HcDG+aFrpbEwNcwSJiP8F7Z57b6B2X67B1Q
ru/kMFG0M2CP8zW1htoxbZbo8OLz/2U4wQTgYapBQraukCZVq/DIRzE+C1P6Nm02
TS+4H/2oA1KJfh3fYbgO8td8odymtzzEbk6o6Ee/CiO+R7NRqKn9goiKUq+wCpk1
t2noSlSM0NOHASB0nGcmAAaeS6dIlePkFzIINLGPWBvxwXIcocgixi1YgcOXBFxt
c9gRMW8NqB73WoklhZsX7RfvtkR9bW6vLv4gPhiZgU3hRlWJrKwCkCKUOOwM+FCw
2O7jeogaEYbF55DrwziyJa2+Ze+dJDgGL5juVNbxz2v3CGNU+xAAVdM30L9F6EQQ
7XeHYsjrmiY6Q2M52h5oLcdXQpGYWgZcAFkBXcXDrz7yHPzdMv5P7cV2weNO9msO
Tljdx1C5SKlpFDLNy9BghEPYXNlGzBUQZQeuNPHHPn4gdrC08daiwYoFfFN++tjz
d3ZYnJSbUr5awXOlGz7wwLArCecM+/iF3wzeFRlSx8hfLBdXMSnWoN+NotZhuarA
Jx/fOc4Goizt/k7GuWtGFWc8Y1+WDfqgXOteI27jdayTWuL8tSU4mcUPl+1zu2YF
zNSdC2GAbTZ66kZBt7NxUqVDjzAOQkk7Iy3gOyKNyqq4ZeZDvaWb4PloArVtVZPl
LQbJXPsSqIsGKom4UKXTSDNvJNAV79whDKFyvBPgjrJYmByfKzG2OSfI/yFHuSlE
As/S+uVqmq3Avd1jypGTrPZnr+kcTEk2y5ugVXQlYrlTsncuJN0sbcoaDa2UzfPM
bCtuYrzrK8pejROw3udFagChd+zj3BpDhNgfhpy2LHP/KNX0IOP947XAAkeRUBAR
aPE1IIJzpw4uI4p4/IkDVoCxoaWdk+AOheJ9kcUgT6hx5F2Fhjn/6JKKKtWLu28X
u7zA7SB64bmlw9ySsTpPLi2fKshgl4kpW3HUsO7QkfS2YllkkO1nWRCrka5RzDJ9
vXP+CqmhtBLD3dn5VfoZ5rosil96H0w0RMJX8d9vK0d/qz57xG3lIDkx//cIonnO
cRvW+tvYyV0JPBsgV35AZ0ubLvdNOdPWVNpxHpSf1MZi7xKAWTuzEgbA5dTbe7uP
vrKzxEeNCFOANKduTrf+7xPyAWBHgRlXqVhS5Co/KedMDQ0Lo9TvELvnmJPN84mK
0Q4OeDZhES4GnWKXdfcrXHZX3C/bob1337D9rSQ88vcMzrILIXpS2qNp5hkhU48W
a5hIBCoGMIx6ze6Cn20oiwRqjahnT2VRD3eidQURvatuvpl4iPirGBYRKZ3q+M3G
u2R07agBCvbJ21DPweF6IE7TzhmxZZ47JldAcokNokk9l6vsgD3RuBeIOuGuMRk/
g/5fIbTRElcM0FQeIuodargON28/ly0cG+NUwBy1EpxmAeKJ5DsunesxNLtmE4PW
SN7mLL8WXNJBp3fSAd6Q3I9Ur8j1ZKmln5P5SNk/JwY8/31ATE2cZ5Ij2q8pJfSQ
XKdH8VZcX1Ys4WoflvWvtacSBqGacurlrnXsipZa3BgKgU36ojrKuZYPA4G6vSP7
Ti6yQiQ56u2WYGUiTJbaVzAGfIUi3gWsiefim4H+ASt3kSwhjLD0dzkKdp4Gl+fV
JTkKN6cHNG6+WHN+C1n97+N0NZullfK/mCYzu0aH3qzI8P9IP69O0JLobDxz4r1K
2S3Ix6PiblyZKUjT0Y3VwtJlqUcHdx+n76P9mt6H9XsvZ6ZVqDeNCwPRKlsX02Xz
iZNKBcjuX25M+IK0mYWjx4/slTCmONIoHfM3blEmbvVEkkSuL5iDN4xzCBET3flB
+Ydy/zeXV8tkk9SBFCsTiYSpuH1nw4m7eNgZvUqulILMp3iRVyi+QYnxzwHZP5f+
CTv2T/BNnaMYfKGWmkr99ILuaKONRwe58zKc46BS4Oyq6E8bLihzLq7nDeXVD2sB
6x6Oelb23KAjRVW+e/LxZsOgr0WXP7ag15ZedVX+uOBoViJs+zpbp73MZqp9Tvqn
+NHXuBaF8yAx1GeEhu3xpc3TnSKWhjb2tlZMYM0SmsHS0ePSeEAF18pxcgAsVX0a
b8rJ+3a+TV6qiLh7VPPIpbteKO0nin20kATio4ZpO/dbWSQpiO/0InYN6SOPVJJR
P4EStQmWQstu40/OZzsJBzbFaeIphhtqXQNAJ9YN/S0tDQJW0XijvJ31OnZseTL8
+1F0EcTs7rEMUsPyj+TfLYfv0oHwkTATmIHDSK1j2Jpg7dVnZkZTc0jvyfm5tGMD
v6F2X+eDr5CJuL1kIqoOwq2oUYlKFAZBkB8oEZK3Qd8U6Asfg6tq6bqW19HzVSbf
805q/ruG9pEC+bFFSTJUZgoEh4uaWwo/5LMkzM7cBShWegchRy8SwKrci8LRNBEs
+jGNK5DKhCU7XvY/PFvYLwEo6b+6n7TQ/O+ELT/ce+YccxFfuO/uOhWcmB+dxm68
LUgGVHq65U79DdF1izXcotBwelqxGkMa0cSU0Z6Z5ha4zXqUpSExxX1rrDw8RWSn
GPqoz/I+G8PFn1X5mefLxsy2Yhs/1LoVdLakreBuPiKD1XlETl3pVsSHggo9KUoT
StkAQZKHO3JDlcTRxpeLLyFWprennuZ1Fxl3w9FSBB6O58E8fBfxPxvU2W7wVwII
JkQ8IWA5yzCW0ZfURBXSPY0SCC+Nd1BoKl6MYdBk19FyNrMwGXYnJm4zORcuobWo
fEnAS2Hmkxb+kVHyEktc419czz8jcGWTq3CtMMnVTgGvvMtcmXPk+HkVELD4Wkoo
iBYBDnTHVv+AhX1OJL1z/OrABuwNxqKDT1Goj8IWqO8UOlVkiiynO6izZ0u0A/Ye
o0jVigtN1MUMzePDuRbfWtEBDy3lXGsw72N58kCII0us0Sx+6us6CaweRidMeU4W
C51AqQCjb8Th5DmI6l2Wy8pO7eONYfkia59v5N7zpq9yYMbuHfw8M3UwiqJX6NxS
kBo8u2YYtYPqDfwcob2RWcfm9ry3FL7MkwlepAIDPKB7+kAqWgXqSeV8qfjB4fDP
VgO1bsvAexzigDwhS57q7ZKi4gz4G9iMkTRj4Ck7gbLRqZrUn0ZkZpZx9EItD7nY
N9YvffiEaqhyyj42E2rCpMEt45wC/Ehn8NcUGsAi4yshUajXyiH/Pmr+K5Vzrpyd
83P2DU7a0c4fJ2uQJ0WilnunknCRTIp5PwbYBXe3xrceIsHBX5jDuEqfZ6/j4ZfZ
OL8ed7prwHrmUdNCKeI713yWuG1U8iaVG1nVaMNivGLMqQhuM4I9QmCXfTL01VRG
UPWpGsSbU7Ns31wwFSxIGEYjwZRO/VY8ScTFC3DULXjtJmgvQl+NQjy2r9MYEx0S
incb3iXMcMkubhDJuJ9zw1n7XCTo23xguFr/NLQ6x5v0NOtRbluNum4bUeOOMtKz
2gWtGrrQAkg2tle1ZXqCYJrd5VOwKB+cdHU8KIHS1DYyxwBP4iQbVTtj81FBzPvC
ltb5qHET32yxtNk5NN6Yf8BUrHHMQULZ0uVrYZKnrEyPmgoiLRomGvmJHcIFHO4m
PBkk4zA6n5+ZFyr4xrWr4g/ugG7VzX3nh6MgGr9xKFZF+UlkDLB8WREo5lTlvGTG
83CdQoQ5DFIPrUP3UBR1pJPEUQOFgqb5mg45Rp2s0SiYHDp2LRdTzrdtlZV3orKu
gnivn63z9Ev780yM1YTfIU0aY+cm0rKDiTunjzdkitTThmVtOVpeRuhoiTavwfni
4swGb8AEYmFLAJ66jFicBL1uwGu7bcv/3kx6wVdrRxPsmHCUCJJe53PRFq+NfQl9
dacJErxoGVdahSQf7xv4OiajHvQJWf5Y0zQtADENn2PVFcNRyvVewpGzIzwsOTiJ
JueNhf79XnwtYoCD4iMz8kt5P5nKcqwMCBQBADSItrpz/kZpcxanWlPZ3v+cJmkr
PfXxBUiGrLSb/X1hEd0DtC4rUoOerqZRH8kdYGbmCm1RKzfVAE3GrLi7Bv4AOiit
gCelq3egaMe6Fl+dpW/c1GHGvTFgTc4waeV7rWVExJjp0V9T1NyiYNJJQy4RgmGG
YoJ53y2tiPZKKHe5M2MnJexorVhsc0jvl49D6rDlXCt+3FHVI9Ca8EX8BBfE2oby
OMnRaH/+b+kYHvX7Xx8LF+iehdImykQChZEA/Dgt1JVsocLTgYhiwL+aE3UN0XVU
12eCRt8Az5d7giJRtBCnyNrHk/l7O+QZbKnHMXwpRZiM+FexivT7M+V6fX4FhdJp
N36zEPsqd3bYee+/8tnrer0CoqUjbZ15Ekd9/4H6G8i0z/TTTyhFjMGQXoS62Kfn
RFqKe38rO7LGpEDqzo6aY+5FifY2NasZteeG4vn4v1WO7kdQaTn7oUgkdMoN5A1i
cFePeDrIWE0Mf6sVVhqDlm0/BjnrGAFECZeV2BLQCbH6OHcfIpbdHxIOly3/y9mV
q7tKGW9H9tQHaVEFUMyxw/P2yLr6nNII9sD5wSwExv9Jc1eiLj0OYw/6Tn4SjIvY
ZVB6ZOJB3sS4804eTxTz9+AOY2EuaIe124SqAcmtbNhufn14p8xItNI/TRVwvREj
ReAR8+2vaF1UuSbU41ODiv1mbkc/y4eP+XDr3c59mp952uGsdzSxhoKC86CbFIny
jI1G0R6VISZG0zhC0u9/faIqPwbK2qFpgnVktvqxcJ5NSRBzszDb/tLvDEj9NEb/
6ppHfoE9b/7vymkHbhG/GV4l0lnFwDsaMuWc1LIESUinuBjuos/UrS5r0edIDgGy
TgHFVOXFUqRMnWfQ/0XmsGnygTsAxBNNX+tYYfwB/uxCv3Xh+L6XPUsm/plFsQ1R
fbf8LebQNMZBP9jK0xf0hCemiB4xV/G749TlbgodYpvJD+2ktFD+aTHxKThqaNw5
YVdBGhVdNLeAgdimVC4LumNbWCJ4xUIVB8k+QhUAGzNBFFSuAIZddgqGJKxUSTVE
FJWXuEeKedwGbUO/xrW15l1t3Y3BqBg3RnG1a4Z3XxxXHWNHB4jusNLhHLSCFQww
vVfi8Xo+RC41U3HYJ6PxBhwV0q25KxLe1MkTAfFGcry1XtHm+KlAIVnBUQRWOxpG
Ape0rxIqwIW8xgCPskHviIGSVFKys6S+2jzTNkqk5bQhr1dsbL5NmJTjfnVS9ayM
ajyhB8yMHOqVJe3bXHMscXHWfKNIKEAwBe4Tutc0KxvLRANUWfMBwHn0VIm3nKQA
C23UcBy8FlHbn2UsS60RK255n+7+BiT+Bfn7vXX75MCQ9Ozfi2ORYFpPW8C7BvZ8
bm0ePtpam5hsf2h/1yGZOqO5G2YmUg95p+dWBDsexX9mV18e3NG5hAJV+mQFu04l
jQruxmsVjgyVmDqrhK4EDBie6MYkgspiEFyYnqN6wgTjHMoatd2Ze4KOgPNr++Ri
+Le0jRaaN/9OVJEJ6w2KF16ITCtZXZmoMroSGCzmSrPcIrmtI8xq+gqZSl32E/w9
dDu/MduugOpL11W5X5XS2IR9y/AqH70ZSsJzA2bGQ7YBTXwaLQ5P/QOrpnw3gvXi
w9CI7/HGSfnvOmf+ca2RDoSzvPUGUwwZFZUMYNivpFf72HzXczohJ0SJXPDmPTwn
6vXu4WhHhCnHS9xjSS1Rt0vD0o3dR6Zw5wWCJTlTLQXm4iegfK3tv2avGqYjjj2r
a6JPj64HuC8MBSSwsBoC/O9LXkYSLLYNZb8W3jwZxfPQKToSU5Ch5yJbG7ZCGc1Y
nfP4R6ErABo8KpS/DyTsdRNG8p1znwRDKEbEykN4oMrWebbME34AXuo/tjN9Cb3g
B7DfEuHhYsc+jgAcrG95SM9GTmbwfogV6j1H+z/BuNjkSXYrlHHn/pa96qK0Nn2u
PUG537lPERNIvMFiW2c8gkUd3igYL2hXvHLV2oSsWyLlqTmGzSjRnGkPqBrYKO4c
5rNYR9mYD+k3Agmm5us9pLbRq20ZpSi+5amSueLOYKnSZo/4HP++oaVIU0f3wIxF
DMhZ3ZHM0S/rhsxEizicenaZ4yCg3bUJ4/5fN/rQSlfOw6CfxmJ/F/TVz5hm16Xx
Xnymp0rtNAeBANjWbLuPDxqxY7d83+EX6xa0C3UWzG7uCbigvvN2TiPuWLrq7p9X
QOCmdwK3Ll8lbcQ+PMULFV/NxcLcSvnEWstP1LVFZRveFrOb25nhBsc5zxHyR8Sx
N+s+4ViI8Pp6qNMJZFK4ecKtjJaawS5Ls9UzzFBOM0njazwBSqrTA46F0pDHz3Fw
6S3NiY/bTYsGHnhdkSWvtHQHmm13prM77c3KfzP2OyuP3Cu2c0yGcFPZHX3OfEH5
QJFwymzHyiUpr9AxsmvMXMkFdWi5cikdUkPjGWWy+jMXiZ2XXM75le+QWIY0J9P0
W0EhSjSw7oJYQskxnmviZaFzrn1FjKJ/SnJ0EITqicyk9GQNBor7T/Y7y6Wy+APb
2NGeg02nuwrci8YAFJhh/GKYHCF4AlcXtYGXUEAlUPPfLDz06GGA2ImvCAKbPexS
BfX4vVCps51QoJ0ReOxBW+l2n7bQMe5NWHl9rMXmeUHRTQEeakptYYDIbtPTmyyn
jQy17FrNtvwuBInVhOUX1X31Tis7cuQctf0+8W2aYa1sJZtnQIlnqOZ8CVu0GSrn
t6uEOespQ903CNAqaQpHACmbwrwMyELJtX25bRPq1UWIXP4mPiFxRv9BWjVwpc3i
p+RBMAi22nus6BjUoIuWbV60KF4+hkA+IHs+xxVmbVtmSroQtPxJaIyngf1wSi35
MeuBtZLUOteUroItWyAqIz/lem8k9PI5CU2NB6JXWXlSkSuxOsPraH9zcKnmhG/y
FYF1pQEShQZybyVUovMwpeYacDafxBSSHcjqg8NFHcvv3grzRiIgo8Bs70D0WxSQ
sclpi/LF1qLqqgc1dMKrOXuSD6hpYsYDNVlrZ84q8C1anqsrMJ4gPJd6uv5vuQPx
LC8GZqPY27nm+60cL92gqbszXyBS0Ja5GgJNC7JAafUIsU0ZTR2ZIQN0E8QA6Nsg
iX4hCD2HbrDqKfdyi1Y5KduGKjIWV1S91hIy20RV7D4q1QT2KrRqt5yh5i5pdYVO
onWKt2Rv/6BmWh8nq3N+uiMmBGEeRxo22xQ5mNR7uAokSZvLkDnolqDWLQvIGol6
HWP+B0GRp+bMnhZu222FpM2eTBRCGDT2nGj8e/HM+hCEF1PkCd9HyaHCYmslV477
yBP6fs6kf3ipbG307Zv22lOgAR8jvyDARt+cwucTxTmhlvh2l+EXcVEd5qAlGb2P
+XXyMaa57usombG8dcjGaZ9HOtpL+EVjIDe209G6kDEKIWYMsZeDrvudVG2GuSON
Ar/NxCRwml80T1hT7hqFwZ/Feds8gbOx/u0GK5Tw//l23FoRRQpFne0SgBHoGMa/
6zS+AZl9iXb6iCJKIni4Dl+WAjHnClWzgqtV28snxezqkbuq5KMGQf8RAVaWhMx0
l7NTg3XVG6tunfInkmso0L1gpsCFKvOpQQ45jrdz6TvNKcG4tsYtcCW0rrlAH+Na
gEQMvszj97PZRPV819qao2peCDyXrwLXjOXBe1sYudGDMwdTKKMv0UAglj11p1E1
1AYfVtLdxWoOaDbrDN6EUTQ5sFL52cRyfcAignrfK/k4MZIfc+cdl+itIVdlWczb
HjLkLnemf1YAQGRMtKPi3uQMpwX/LOuI5wAeVBG1FOSgKGjDU1shS5Tx1lIXb4G4
gDSUBAgu1tYyk/R6Abql4Gay8I4nAO2MaLUY8E7AqCv2Gb1vMm9haUE3+igWCSjA
AzrKK5UovEgnXTbFY2QqhnPn20PGebgoRfueSjJF/6bZD1UWY3+jovAhFVxw0s48
FJ95FF+qIsxn6JYxOxDgGLDwBzUUIB8+2o1KkoQqu71Gjdwr/CnXk4aBP4a+y8l+
09Q02VrXAmapxiYumq3qh+hwM+Vjfgflj8Mcn9s0iQsaRM4qzZn0S9SdZiUyC8v1
T+D2HkCOnZqM+R5wbBMbVTnY6W+l4HpklLOeD9snOB8bOm2S5Z50gnRAZxnwmdna
OrY7pgQBs5gU2bry1peO1JufLz5T1v4fG3KxArRb0CEO8/tFFcmRRmP/s2fjVogC
9/KUCYOosJk/y92fm4M1mACW3sHiwY0fOJgENeHdCg0rP3j5IY12WL2LnA+vnCYE
ccIqm3yh6Vsjwo3q5z6HIRDfvrkqexvGx5F3xjdvSmKPuTvSO6B73SHnNWGSvr7K
wIeRr0fIhnSYxME05dduDZwbYNHlaJLPcuD06NvJ3qIdyiaLn6wd61TnNPUEZYtv
zqH4sFd4WSLStkF3TdAl7+GqydBkX11wNe7C5t/AsWSK0uJlWarNDbTUaT2UeJtS
ycXUn4ItauFLF3N3FM7zYVXBp1zVH4wbpY1zKGGjWXPHyMAJSo2CZDhu66mv7ACR
k4dq9rkGu2uz2LPxSBKc0x/eOnKCNeOsI9fXOCOAMDHKa3F7vG3Sr7hRJ+XvqbHX
imUlhzl7PCA2ydPuEVXCjQW8IJWECg4R9xGB6ORmEGA2CkqSTuToyLVW2cykPzzK
fziIXAfWubkAZw6pAWCbXONDYCJaIWrZ4VwO68r9na0E3HNRb29ggBPZ4CTe3Gro
MqbxYloCdnbKDbzJvW2OqBFA41gPDYR/+7c8ypfXNKAGTsz6cJXk4h7lXVbMh4z8
38XIqGwX9MQP63OhMUE7e8pt9xNsboYLFQYXx5ZY4q9NrH3/TjkH2/spPgyYtZLk
aIZQ0PEmCI6R5bS5Z6ZC2WSrpcleFMg6dNwz4H9+mVl36JuFdKPNG1s+3bC5KpfO
1JM32beRQ25dC/RUbEanXT/W0VpdJnuIMGAkLB0AdZO04NRejy30NCCo0qaEZxAP
FKpuDy0CKwl9uxQKZP6Htgl9FHgwBvyvGrNUoN8F25gUAoz/XE7m5EUnoGcmFg0m
FhxtDChk7nW5EKtLJKSlqyTDycGC+Y/1W+GlxpSHa6jENJjYJ++cCfCvXezhld3V
2RUGmnHTJ+MhZzTlT7/xp9qggpA2h18KZOg1DM/woTqnKWjezz14LFLd3uJVKnwZ
z7WGClFEHu2o0FHRZ7VsKlYjP0y6a2Td8fEsPCcxcGeipzV3AbsANkoNAxjesu/i
dNJ8vgOqiK0PWWHcOgh23WlsymH3V9yh1R8ux/GTTDZ7CiyIAnDwEHDkHK1dDH4i
Bspc3QrAd3Vvd7bSyyfOFY3lxev4ocYUWW0wJ/7Es3cT2ixthJ6DF+XsIKPJfTus
lzRdMoROeppQAboWopnh6UbvNX0JO7/1xAmYFXtbx+Bu6YbkBqtIYjh1IjKRJcZn
JLJpWrVN+vlPHOi2Du2hH5CRP4Dakuc4RSYIbqY5DzcMeqtCvF0mctVFHZAnwMJ/
6wlfjgry6JqHOgJ5uNslkO7NcmITdAFmsCAPmMKfOzybZf0YALq1tvXpG7LD3iLD
udK0XB94jnoTxPUC/Eo+I7D06rt0zjyCwjCFjVR9ZhhwqUOcuLxCS4WOmjOONF74
DieJ8mAEkyCCTAws4m0eQZotEuGxYNn2Yx+3wEn2sRrpmlMYNbcbhm5D5ZhjW11S
asRjLuaw+KzVj0qKrXHrtKt/gRS6kmKf/7OmKqmXjRSQHBhxYSYs7PsseGoa1zlQ
q0wHnOmPubI1iPHddCkvi6Paahua9Y3WmXDIdxKvyXtAiTa8qlzxondBziVsjXzf
NbXCmzyhh52eFICuZWdZt4mUhU34eMrlmaPIgTuBGiWYEO6eJh4RLJ/4pqmQvR4J
7+bEsFH2njW73VhHrnHV5j6rs8sNRc0BFjyEsTc8t+XEJUsHgX/tHtjSyNFM3il5
mgfr/VpyILzX9/hXSbI5xNJIA+PN4nxJ6W7L9K5UE55Yg7HkWzA7Tpyg+KpPs6/l
fqyF7mUbfrxpPYp6HR5lifAe5ijTP+XKaqb835BeNBqLadsgz1xbhHsgtAGT0cOc
meuy69L3UI5nxc9/4lDe3BX9bhlYbUs1gfQZy1rGjlvs8GORr2nDd2O57aF4RXcx
QA9xmJHpeIToztW51qgrI03rX05570TG3P+PqLFxcKicJK8JM3FdEoTilAeKV+eJ
WRpSLjHL0JNnrxhHZmnAfc5fSRPoA2/MX+xcao4Fby3yIOskPRb0GKmAxl25HKjD
OiICJ7rkjJhpA+f86N2UedCD5dYIjcOoolfbCUyr4kjVgMyX1Roa5C/COWZOwPFn
PefqxtR4D9ocIK/CUJlXk+NoKEPlQ9RCAa7lEX6hZSvQkCC/SqeDcB29swVhV2xr
rr/SphXlhaJDlbDO3EdPrKu98TqMTpEfNOuVpR8ccZfKlHxC9KQKcKlVQGcGBCab
bBydSIkB42k14nGZV8CvFcZvnp9CktGDq2gWIsVr5bo3hWd+aH7qtmljLL9T/Ibc
hgzhvAzvGm9zHQsDlH5yvemeUKdQz4yFrss2XGuK+EkL/J6tjKvR2NhlJj+RpQaM
lULuDHOhjvJyG4/OR0ZFeJci+nqVTnsQgH+oIRi28T+3Gz6maJEP6nB49wS/CEUh
1wrRR/stdF3xyIFlQ+K23bJwViKxGL/yn/DyDVRQfy4q/xP2ff8Cm7sxf3g7TdMM
2AmMVoKa61iaAQFmZDPxkhswNloa4vy9Zf18vrjDiAlBn8gy0A24BKFI31ULZpYb
lrbxnsCxa/ysy3k3Y6Bcwl/DHGIs74AB44NNCpXvB8SJaTKYt4GdEeZZJb47Nyx8
P7p+J/Y/tkYq1eBO5ClS+JONmvCkf+3SRMFI0pvNyVQxwTPBrYjNYc5oYOFrNKJR
fo6idHs++yZIr6o7rlakteJ8v3S6ndOJwESHsD9G3chE8weDXa8GaRV4EtT2OMIC
QChR7tkq0Dr8GuVxhRmfyYPBbfCBsqpuJx0q+HVI7innoWXiCW0IpHQ55IiywPrg
bmc/8cw+XjfbJTWzPURIdm8Qw3RuWR/8NFEA/EjvQqmnavkLadJ9obkcj8jZBZ3v
SQ5wSP0aeI1xJgJdc9vpCtO/GQeeL9ps8of34pCQ5y3MTwc2ZQON9E+5bXzx17+N
4SJD4Eu9vi4PfgqX2oqXjBYX6cnkCQPrDmR3WKAHONmNz6wS7emuqqKegsaLQwdx
9L9lJ6JN15t7wTI2qa6tI/BypZG/v6pSa9nEGseI718xa5rGd9NuA8PPHRNFtIRp
EAtQxCZBuFWQBVQjj55vEgirtBiBcZg3/GO6YIrjx122xoMgQoSzfvCS50ZJpNdV
oZDR1Ck+c+8XYThVDTUzoEfrbUxjtP1VgBjnU380fXQgLIDt4DU6q0Ashqmz6Kot
6xRs6EvZJQCEjXP2yY2+0P3OHa8pPhtNX+RAh+KBloNXH2fbDkWXRr9rswC0PH8w
rd+k5Xjh3yLrnTdbIt4/dfkUd9IILEu/2WOEqKaXyUMmZJTrp12RNHzlWBBPAXRO
mp9LOIZXg+PVzfACBsThSTBnK/375IhT8Xy1BYhEPg4KgD7Z/56AWCqCpzYHxbDq
ZsU/nzDfRiTny2vTXtn7ajbQwJYTc2L9sbWr4RV8KbBnIV2mUa6TR1ODWlJO52e0
epDbEM6RgDQXxtokxERhskVHMUJ2sILj7tO8ujuAlpOqot7M6kDWRboi6Bt7tQkm
3LYgekXb4AE2Hj1EoDpCH0CyRxwSpTb9tiP376kDZMgF0k2NN7/nGdmSpl86yv9H
djMR58sEht+kppRupUNEzh9miStO483v1eHuNTX3kvs+R3VtUpR+oNL5y15tUbSQ
rDNuMoFeHWgB27lJYFZ4SLW22eSUcWnIt7VndyJpLDJBEB0jkpbbrVJMrqqAq66Z
74QjdniZXQVvH4eh7Oqw16j/qM28U4VLWGZLHFZ5NYHkS3ZwylSA5cUAt2Z6XL1L
c1MxzJiGckn/4KKmIASce3ru9RG6wFYg3aSimA8o2dL2WB4wyBEtlkCe1A8Mq2ga
mM1SqHKrXi+SMj4hc4k1KCx+LK8Znj413a7L2FUfjNDxUzHR+xk8nW3SJyNm38TY
Gx22I6mjT4is8mbO7Y1B6xve+CPiUVukl/Z5O/WlrtV69vxATTAVFe+NbYHsSxUd
4Y30dpBE6pjOao74/RM1yrxAjxlt8Qk06yBWIruZldcLoqxE1WXI1wVEN3/W0x38
IqsyVK1/0Up/GnMl2qYUBuPuNik0qZN6rp5SEE9nd9F/c14u18AXo++YXDgbERA9
58jUsAZxYYf9G/tn4RDYlseFNiDupHk7CV1a4hXRdACDUffjYuKhClxSs/FzMGVP
neAdKFM+eCDUzmKFEhLrD19KLw6qnQYFvGem35c+axJv+LHOlU41Tzb4oZV2ymWr
Ev5vwYgUsi07tJ3FRhcnyHIouSJTkLn/noZvF+B1czA4mgIVKNmwqHU2FpabBqKr
mVOE4QQrbfPLdxOrHBrMmYKuaUYpwmtw8fkvAeigT6YklFJhEx+vAw/itvlyOyu9
sEJTfrX4jz/sPAdil608zHPqgEKEB6JeRU/WYONSK7ax78LjkBOcJrp9R7wq82mv
XAx9lrWkB7kvoGdDtzIINXFSoUjQ7ntNEZXfGbsCB7EqZk6v0C9/FjVbATAfUtZ3
/2NUVwaU6omUI3PxAd45U0A48qN0MHSdzER4CibS1S2UWze5pw+1P1Zgc4Qp9yv7
K1cpI2zmL379LftV6891g63irUBFFMorhQTTd8Dt3CMO/aaME4De06QlUby0t+6K
fNHbw3pSEk4OWOPktKPwJ5rHRFoAs+BQdEpAR9Frx1owRaeJvScISdmtBpnK6FTK
OJLedLNEAdaD+nAveLfLoTlscdfwCDxtD3vwa8q0tLF8L76TLYOIp6H2gtE36ajw
YT0GV5qjHNrIha+1PzKMKyATqqZ1XzgjheWpqBsTp6oezEZNfyE8RyCst99i3XOy
iGjKO5KbfYnemICI8sDRXbv/bYci66EzygKo2DsmKnQnnhIuH7e6zlKEIu13NYTL
iw68J7g35Z29Sj3gEAu94dl99T1sjK9QSFynGoXIbJ/WIAn2JA0z0XhE8RJgbNCr
gthD7BU+SowjzgjAj4gE/nDn7VMGXlQLY7Ibj70ePWH0dJcw69XW1NvS+W1mZUwZ
By5tf/jRft18Gd3Nx5TJZr8B9Hsp/cUcQjCchEYN2YhGFDLU05wjFwiA042SV9EB
B+Dv1JVWx/0C5jY4A6LijZv/8lLQ9SA4sdyS2p+w/9aySI/0papqogfXvgITskNC
AE7yc9CK0rbBvvd6h9NA5gEglotaOuUkYkgzTNYlbxknwKhccoksViI8u2gUa5C8
+JB4hH3HypJ7obqP5gjq2OnXkxhFhjXd8/i4w/8ZzetCcTnKpGZr2iWaoL7TDUEE
rdj2D3B00/1aqss3Y7GgT12f625vzqZ5VtQj40XC3Frl5b9g6FSDt3R03zEmmGQ0
yMQZpFNRiJlx6dIq1Fm9YGIrejXF5hpUchOmr0S6K4MD2Mfgoln9dd6J5m3R6sGl
px1afEGPhJmDgBWwQr2KV9DzsNPM/oOwSrucV1DiS5PHAU757qaEBOu5GTndCDdM
vptv6dUDl3T/P5jkVbUq6S4A8z84TMhSPQc5Qsl6soNJIzK4W1TYVcUvIAcI+JmW
aU4k705y7cS9nrLY/RQj5UMMg5SU/KILY1r4ufJADo+AUFh8Qu2TXBF44yXLkN5C
OZf1lW+Uir9PJ+5V6t55TNMhUJ9eVfFOtMfHLBn9KzdLGAL17H8Zvt+o+cJTJcgo
FIgzLZkLLNjUhVWKHoAa2xMdeLNiKhffuaitfipvjK1xDRb1YDBPnrBd52BBkPvT
iNt7S+3UQfmFpj9+POH2Rm5LnW9se9zZ4nyogh9m8mZJhp62hngRmVM6X6yI+bhp
94jqr5/f9K7u4c3ymwmKj2CsHdA987uVEg5RlDP+LGMCWjTG9T/BR8gbsCWl+58T
GCZ0PTB+9/X6eiF3CAoHyxqoS4ZciVX3nbobNMEvYpqenoHe0HIiH2M+IAHpEw1k
N0ph8Jbuo96yQVPFakitfImOiUY2PI7k5kUQGlBRbMZ0Pt9sceOuEX4m9HPwL5aB
YXQNc9KlsdSOxDFGcn4r1Ez0GwDCDnlhh4kNXEtZUDY4tQPVjiYYR+c2SQsZIHgm
NqnKsSYTs+v859PN8ERUyQH9Nn5ehBqNm5v1weMiig7eFr4FGCNv92hDw7YyGsOq
g9a3NdCVbz1LblnlZ5pxyk8fqwTCqCohxcXR2lbgrWgjHfcYRFarGt1JLPEPEQza
4gF7ar7bgFrjvcBnkYmsbYsQR/DkdSxiEI2IsC9InxF/ufBT2UAs3nLXvuFJVxke
Yijq2dR1YLwXNTx1NENtOG0RcHPMQME0OehHin3zTBMnKkIby9iP49a+CKqftNfX
4op/l3tKTVzmLCbgi+vLvS8q1dJRCTX4mctzjGXRNRRvG5J0baKJyglPNGuC61QS
5NwQKWlok1JgFnvE+0apChExP7rj4qVQvZfCpA7U9lqVJHSqUV2Pwaq8yrpVODQg
mrlK927WfAjpjB5gqp5rUGqzRi7AvmcSCYDFDh8zPNBeUC2lpqQpyvwE4KYiaP3e
YhZRUMCHXNauxgqTEbJ/eNzYiWi/BlRlgylyl0qWO9ZHs0xjpkpc2ndLgbmXN97m
u+8iwssxgDUNQJQ/mTjdNXPL/Vml37h5YsNHCOzDpmCWcVJyVTs3gnFEpxHBV/rw
NTFrPrImVlIX34FFu9cl0MSRbiMute1Br0fMl4gVc5rnvvLbE1Gk29Q0dI6TouVl
qFmaTO0R3NGe+pAV4ummk77Z9gqGhvlg2PpLecWt/Atqq4GMkfd6zCTMIZMVtITj
0vv6/9PAyyJyqowQIq65rDUQoaWNcafQdihtsmzmHXoqXkvVvqfGG0sguZn8DYQd
EKT7ofGgvCxfL7MvAYYJp8bbIOKkbAmiq+g8BCfipUy/cPtYYwvkNvhXfyduAS0z
qvD0xzhtqL2zSJHqxjeScVSvWcRbqqxwhyAppHmu3uZDirOPBvCJPOMXe3YUzY2b
+oFYxSAb5xrkuh9z4IcC6rG2Wof6D7aXm1WRJzzKC/0SWpDZnXoVdTZYLb/VeUCx
TNimY52l0bor/IQJGK3ugrGptJ4JECHDhGtHIv5idk7dKzsI1cY0Tws2GUFzuwe3
6FZdCBa4Fwb/afdsK+jbdq8TeToLyAX2xO4WvevGs+HTEI5q3XCpBFcTScJ24doI
6kHqLSQ6qBFGhZAYeFr1vUPd/eWbbYmUcqIEiW7DwBXjDzQduUeCKSQlOxNSUYN3
vbYMKko9xtobeu/og/dO2x/AuLlrUtAP/QBi/ZXxS8p1JM+vbOFMbeEYuJL9Qe25
13Ja59abrkRUSd7eT108ZDXKqxW7tqEAgUAv7mWGSDSy1KFXLh1FMX+y505da8jn
7tmRaIUeYEkC6p8uz51ipA/EagaLEVEHqvk6SnTg5omip/UzppeoOiNl/KwX5l95
ldKmNGgivFuknZOzuthgu2uzjIexCl8nSry3DIJYGCPIFKT/6ZvnyJOODClAOCb7
LUYe6aVmZFa6viczVrUE3SKifRfJt3SL7aal9qXg//tqy6rpJ91uXdUKsIdNTS4X
FOOWcznVkaMwb6WJ/s50lZqDnmFddxjOsSqhZNeBkhuO19lT+GcAqaZ9rIdRQdZn
YSJBISCnAu1OkIERkTbNWDbaXK4wSfw6rTz/hmZ0x2N+SOPyf0/wjEqyW3RPvbFf
YZKaELODSiegKDpQrLvm+25QfR4JziLjeIhuMKYSQ9R/JhNvxgQ1VBX+XbMOsVRg
GargAT3t6aeAN1nsw6KX6AEMhNvgeAU35/znPzLo9C0F2/ntx4mgpnyBc3anPVQv
SDcpze0ne0IRyLrXDZ8LFGxRrF6AFglJwjWYo3cuOqxAwQF68ULFB4vJETlpGvCW
b2LVvGqmBi+KYwSC9ptPu+ftd0Hugr1JJzkKyZxga4b4gLAmqyHlGxrOPpKaTwfC
sewXPsC7i1JzZ8INzIRfiRqcY7juapDLaUErAozytF1E+6g0r0gn2kLeY11rU4E6
xRThkQBy2+726ML6eBqQWJM6OMxwci+LGlddCIxETBFShlys5tWiCGWmqAXJ5iPC
kK3vn1MTqRUa0QKg9M5YwIsyvw8/yndDt71TIjqrY1AxhoubyYJMC9DOu+sFDOg9
lCuf9uI4g7Re5W3bUbhncUhkqMNskDSQeW0LQhInGECo9URlshkVL69RMg0T7SeK
WwWAsYU91hLSHl5TJrPb9oRXfkSwKijaiEPBEKoo4b6MMPByJg6WdSLaDPD3+yPD
MGw+VlMAgGpadSjPatTpyNNyjuxd2DcHmE+LfQVMzODUo6D+p0aAGM1XuejVJYDE
s0COqyFl2O//7ym7e9l2V5xFEwMcgN8LN1hGrG3Iaku7cGWDLNrsQ8liZu/Rss9v
nJLmbnHgEO/j73LgVNiNUyPF5bieOC8+0p1hl6lxkrcSDnUGfv+8iQn4dWf1D7Dz
USpnxUAAHbxFsqwPe6jiL4mc0JFwGeGKsByVxxMjnK+ZP5QWUnyjSNn8bvGy6bBu
lku15Kscro485Gf2LWOUn6B2wqqZgevDQuPxxwNcwuZMtotYDcN1/KBnVa2ulL9U
t3avN8Ex/3vFk0MA6bQStX0fr9W9danrulvkvWiYUqTaUoy8JswGd++ZPFagaUQr
XoUQv+VTcbZ2NkTPtawYb3rUGyKFN32ukkNsUbf3WpD/XWC8MSN7UyzhEG2M6v+l
BzQMtnKadJRwpDM72GB1A4OOoDlFYgsQJawMgrh3IOm1ROu3y5OcNUPhQDV7qGRm
DyqtFY8/qjOVL/VxgwkcHD2uP1nQjYCQYGjX7Mf2psPgtd0W5OB/V9A7rAgsjtQ3
SFWPE9zonSvhlQKuA2c/zXe1w+pf3XWAk5bwsaVaaL5WmeV4Yi9znTBQe2zQCItj
DJFi8jXOl92zrcubR8ke6Lz9yk6rxfek1ljhFxqrmwrAADGgkBdhmxjDGv5Nzz6t
tGVGvMuROsDv47kSu3VcH3gaWLTpvOXfs9VOSHVjz7vc1i+sYkZPA5mEglGby3gq
T7PO7Ks1Vhz9eSFlYqTNXxWoiBdizUYYWi6lPLOzCqLx/D5+6YkMSxT+QBEuHqod
jPXMKr8qlNzQja00V7CB/Hz7cutDvfuKO05lEBExQTn14yoD0GKhjjVR6+YB78dH
5itq/ly7rEQx4DqPgMD7tugV1qSHniIwYyOXM0hSd1WRqFt2rqHM9mIW+1jEBq5l
TYSbyNxEQAGnfUqjOe9MVqiGk4RDadQqa3Fz7ePtHEK4vwd02UDV4rHnHu/sNWbP
usx419mKC0Mc/FLejs5zIP03iUrmh28GI03wDn62m0A4TWkqeoplI8PahP1eSDm+
b7c6h8py1z2KcedVilDPKSHxlM3+EBvHLKu+5xzKtVbrEO42h7K/9b5Wt9Gnczjb
WluiBsczjbrhO4QchyFPD97ZWzCuZqLz/Ljn45v0fxQjd+tVaaNV6z1CPyr98SQ/
EhXSCZar66vRQsHrYAQXXm0USyVj4RvjoWQZT9vsfP34gNK0XleBmzCZCOkqWoRI
Roeq6Kk0/jfWx1rXXCCSyRliPvOvE8nwLXqSwhz9OkJ5ADTaxFYxOn0ewWA8DKmw
i7HpALyAfeZY1t0GonJxaYHXC+CiDHHZviz6zE/W5wWWxcl6aI2qVf82cpjULHN5
3Om/w4XmsiXZKi5UTwDbGK59TL98ZacAo/tS/XkCnQvMSfxw6IYu0xD3HM3fBD0U
XlZOqZ7eBR0gByR9+eOzwQ1K2cemb244THghfYQclG0q/pNBb90kYR+hUhysf84j
YP7t2sTgKcTwKBR118TW5eoIptUL0rFZGbMywrRtSQV0oNjp9BvNDb6SWH1u3P8H
zJo+r3KvTBKMBQzur+EdKnxaEgQeHUDYGNAnHaO4rQLN9Vcv/vfdoAwlAVSOC9Kb
OwBStyoAJdkqmvq3B8qwMu/uJPiC/xeMvVE4AxKyVgNBkAcbc0RZWlZ/EoEkjFmA
icKSdrMSH7qwEyrv6eblr38E9kRCFL60+3jgGljl53j3sUco/BCqILPdxl2vfdsB
FVPF4FnYpNzh2cMPX3r0essiWacH0e2mwMcgZlTa00m+0jIMCKjmVDzbAg0qwVCp
i4Ib1ASWpoajTt+BWgvqHM3edNQfwzVNgBXCrfW6JYGU/peulQ+E+3rmby0gSXD+
jUD9uMXLptHVQ12V/ra5DIIHzW2GazzMod1yXrs7GqR28f4AvaKqvXW1jAk8JCNL
IjWHwcoXBSel6e6QwDm8dwIRQgBx0J5YMwe55pxdrFYuW3CPsq22BkBGtx8r7GIF
r7emXN3JbT40oBk9gjLFLnk9NeNOg7c98uutAwzY1owjcEy0+Xu0X+bgWBR+Q6hb
3hXWP0vXnqSKK2Cx3n09iaQlDB/BF6ADAgq8Ag3dwNKxB02fj87vig2k65A+eLbH
kYqxepMhnLY97Tk0isCGGtIlKRgcZtytKZ2f+194AKwb6M40Ox96uxrpm3yd9tf4
h+JMhTjby+XmHTHMWxxZl6cl2uQvUllwvgUaCg+H0hPMUXjil3Ik/LB+P3SR5FYE
2x5pflALo0VwCdGvP7nsptofxdOVZJreyU42cN4RgjPOwdJZ+wnIpfP3iEPtVK+z
h6px8JhR0H2slskz5UNG2Th6Xful+JQ0SKwi41HVC4aGS1j0RKcGHAtcAKaHjDVm
r0TEt/AA0AvkXcErSD8KumzEfa+T1lMtCWkgXDL7a9CQgdx6mDWUkfMkBsSySzvg
K8ruWvb/lHIQ/TaProb0VI8zI39OrEc1mj4T7CmMSF8lL1bmMncEl+7A1FJY+tJh
wOIR4Xf68s6edWzJn5N+oR+wS/ZDg+DnyON+Ispmi78aD2HodFWo34Qb3UiB+H4c
AVHGzfjBHJso6bIgXQ2p0zqXogVCCoED8QAzWv2F95LlXO1/cmEg6uuXbAWKAMuc
ho9b30KDimfZPe/HRkxLlisy1kv5tnW3VWUZQbnbENZ8rYPf7LAXUnIfG1FbDWXJ
VwAOjfHNvakkuO4dcJ6LpKgiTSgpsNMY5sFHOHYcu/mbm06fGuZTK5rw+vfxVU+o
mAkJNtPih+LhwZie8a03lIYrzW5wYFfBGExy0o6637jDvqPmDb/FD6rqLbuTgERi
JLMPU2SlKkpjiL3cQKXQCZrkTcu09fhiMvU5p46NMvncnrG6kR9RyYNkqDL80CIR
39B0aIc5Iw2Tky4bnmSqrnd9PQOVeAwzxCyQy5R1CoKmiAORxQyfO4/zFoLFpmTJ
HQQVZmdw3ISd7xYvWvzSho/XsHCFSYIkMfSKcouMn99UqjmaLAqL/txqnu5X1Wu9
24MtXHStrGG63MrCJWjTTRfEIYl4ucFz/veXaRAbd3b/ZlEIp984Fv+Rv/+gKoV9
XZ0WQ/uMf3+t5jrpM4PsjKgtcJI4e8LLLoIbnD32yHxGM4KUsU/I7jklrCWuDRap
zbcDqekWWOPViGUU3ZSMuqfWDsJgTrYpOlbFe5gaC7O4uDaHKIzUUJqPWQF0fe/U
Z6G2Rn88ooZI6BEpkfHoZKaqOXMCIYALixnAX0VmF0TZTSuuebqPR+MWXk8bEhw8
6YOVU3BGIhohOsdl+MzOlseBng0IR8g6QShd2JSoFRimYvc4w/AydVQU1wb88WVv
SIpOg4tVqTuzb5Pr50lE8kOL3rxuAkHytQA9tW89t0w8qmX9vpdAtMZEr9clK/zr
7+Bpvj+GmUhysXsyMqVC7Htgnd1+qDVR0SToIVlArmj14zmph8WxXcPvqDldb0M+
Dytv3bz+cxF74edKo3nPNCmqc3djHICwHBs9vEq8in7zO7X/G545tN34CDOap3lC
wTW69gRZKmmdIuWbyEdJncgeLAy4+Gu0GNFU+g9uYOzvZMYd6i7Wa3opmNZUGjFI
WTmpT+3XuKcEB0RX+pA53fXwlXjeHmD6/6jbSnddsjBvfz2nyGUZJ6PsuTc9eWRS
roDbXC2R40iRKqsafDuKkC9ARQl2dEP9LRncru4QYzxplo5orBCW3aeSXt8gKAoN
9xdzKSlkh5lIBmiFToi8Em92eEmR9KdIsq77M8L6g0ftaEXioL+ySfa3xEepsMle
CVmGHlv76iwNwdpF9p7LlkdHhW9JrAb+VIgQIZOFgoSSkP4FrLbjIVP6Fqqa+hCa
34x/7cNvKTMPqLJi5wcLKp2D2fal/WQe8NY07f9XOcjVf+IiH7gq2u9oq7pOij79
tBkw/MkHbosUJIxVEvxRedWQjAB+mlbcAwXRTIwoH8cTwE5QzTovWw9JNC/6JU5L
0gIw6pNEO1bnMcJsTouIn1MfzrUSXx0LPtEDNu7VACVbzvJbEPiS5sooIXafZUlC
00oeEbq7c+abUIwRKH+cP5LM2GRa3B0Hpmb2Af0deV3okwsyTB2MTntoQnfS5ghR
PC+zv6OBOHFKkQbUSig0Kpqjkpq4wDMZOLJxu1NXJ+tAEP/d3yeJOpdvMvhoGGof
phOOaf8cXJX4lCnuI8v6X+hppoTp0No7Ns1fSR/UcjKED5BTgA84n8uZuN8GFmT1
AD6/JTkwnQMJ4/2emaMJfZGKIwuZW+fIcdF6H1wrVJsR3HCoS3+Tkje6oLt8bon+
y8qOgK7JcIhnpGtULwPEkpgF3265V7DVAW72PAx3KpHmazSiDQVHE1IZ9E5VowTk
tnI6pUQgscdQP7gtdvbFqSGDufX9acV++gyp1gMXfYtaEGVUKSBZ9BNjEgO1rgXr
EH1xr6P/AGhOKI3vs3yViNorBhK4emDAyf39gEMLDs+rCv9xNLCZht2TEW9kLqYI
4affpVoM9tR0MZHyu7jA4nFJE8s1YdF82AueS59fidCKZ6Q1RF9i6aLmM0UrvZBt
k/6FLX2P741dOnb3WR1nDrKni+w3TY9PCNig5VRBM3lL0PbKSvzjmeS/BYs8WHSI
RYlcpI6Nk6BTR1E5cFzKL7b+4jUVWBN5qhIBStlne1WbxyR+9OwhxBVgWVJ/CpQV
q6Ys3AI6RejiZjEnKO18NySzb62ZiW9h6U7pFZ8hUqqt3QlWErtNUrCULD4JJLMw
uM01Ts7plzT/anfcCs3VlqJjJUVS9bPY2da1Iy9oOVL26uLoU03hLWK5BQhJhM1/
Wz5ZMoe6nLA5NYZMNKla1W5mHuIDBzY+XCqbNUtWMNiyU5pz0QUzFHcfhjhMHgAR
a+jo3yzWEfNRGU8XQN4aQJKgFKoCg5gPxf2Fn56W+lDXP9M/uLaeVrJ9YoE/eFXa
lJEv0nm3sKCKQsUidCMkh6kYGY3AdMqd2BCuCNKKO6dfxF6Mlh8l4zlz6fH4to4E
a0C8LdJbVPUufwUa3baDNUY3gw0gviZHkk+62YwCIr/Xx7vYCHUS3D+ijgN1LpQh
QYIlK3VEx4rI9/Mux9Xj0a7Jw6dPNtcVFpGgAOiuejSEdhzSZ9JwsAGjp3ayiGya
beB/mT7bzBSTrwoOz34d85lvps/javEjH6vFwKTvDdJiIN97xmqkLYvjz5RCzG1Z
SEfl/MLE0UalMvQp9sPUTU1V4BUK9WLWcl+8yc9ii/eG6JI/isz+gPuemjqrebqS
phwfqaVVXqz+A2ezY2ECQVZUySdd8FHNSiHlgveNOfzl3SFv+QybRccdbazCcvaT
ywRqEM/7DuUbwBwcCyIzf/VbEgsiZRw9nO6PL7yj4yGOcP7tQrkeaEpfYD8AUiez
WI+7HaZIytGXnNeFh7cWkaJirrzUSsVrS4iR550Ad3hOJlvETf5aZpe762Yftneh
PySCcbij5iE/6prkP4nBGr305L+LrThaIxpVRDikWpbwyudeB/vBNnpPouEIcYMV
f5P2v5BzIxSA2qyYUJ7zd15zPHIdj1QTgzkzXnFTJv1Ze3ye0Ti12eGeTpbTjyLR
CC1Cx3kb8z0h0pX/Pqpf8UqeySS9ypgXx42Y1gZ9SYlzTaXSWla3vX62PEiSe7ft
7JQrWZW/tXdJClmwZiXzuG25UzrjnpmmrAghwluAYCY+Q/q4jg+47Y9o7XaDSot7
9ojKWRqTdPPl+LxP6TnaadhU9OXk6ldQMBHkU9o3/Bkk4I9/gkglVDE5EedqKdP9
iYPmlL7OR3Mw5cDZc7GqyqgS5fNaAPnIhSlkKDeMStas3zVBxHkYdupbq6limkiT
h5UJa2hJxpX0fMOtYwRAOBFnD4ibv8WV9pOUfOOIjs0IwCVsfIDC7I5yeTGJ6gAP
lcmtmxegXgpe6q2Ecab0zdHnRPxLmXCZPU964pCXw3vECLGH8pSR6QhNUkJIZcAY
wZiBMlROA6YaA1NpC5s3E9C5JC5lRd5sbI0pBK/8x5gJdKxNukCLMQejd6iP22Zv
HcA1BF1TzmfjOwuz2QlGXXMiqtNYgO58JiGb4Y+WnIAHMdsSX7VPrcmdrjdd8VNH
/W93uHMR/L7UuhTgCUMJm4YZYxBGGAR6vFfPyCG3qScrMSmdL1uxmlkZ0ZzS7yIg
xqkyMrf3uxBhaZIM4pVBBtF9wCFVfbUICzIPFcNJxntgVLSjHTR117DQ0EWsWpAN
YGdXa1ksbznOr6IgW4N1k5UNwpt88gDzIQl0a7w/Nc6sHWaOMjA+Al6G2yZm+1kE
KkqfIZB99TvXLzRJCXvJ70tKOD/6KfojkUPTz6eVZj6GyS7Co1Jc/2uEJmyIO0bX
tRzzmgI/COpWC3IUjCw1DxSmDtif9Zl/sx0oqEkYcbM+cSDGhk02noGS79cdVmjZ
wASaPQ6kgxTxJfsBHak/tyKS38playhgYTmP6SPAX8ptuKBAyMiZ8liO1GrhfMAU
UhZgFyQykqjEJO0MjgmWYLE8J2ZQa2SEg0PvTzd758ER8ATAbcx0Ipw/+izXPv94
4WeWepkfj0L7uMD1KEjb6B1zndIu9OcqqMCmCvR5PGBm1wQ289+8cgiDTIx5lfF7
5fNQXgv6/9+dOjabyhVhqIyfcIQjsyJpcUZsog/qhyAl0BXYMqGKU0sH8z31vuxs
37vlEcsVddGQDIjFbns3iL9qRBGhLr1kCiXY06Uiy4EvLtgsZ8dCQehgFgzE++Ku
LpjL85FNLHG7iTkcJJxiKb4OWFJ7RGw5iXrupCsVQjCa6qCehSr5Py9UJbjGgL8s
TRanRXITdiq3XMbdb5qjO4E6tatqD/1b1MPZJRdH7sqrd5DYMeqrlTBEL+fPz3iD
ukdgUfXB9UO2uc0kifKypQ/8ytdP+O/hbxi9NjwJZSDD+GeHo/xklZeZkJnKSR0+
VqcTvWnQS7f5f7StmUw9ac9CGz3dBdc7y+qXs4Cgnq68dDqMlRlMWBHxder3fjDe
VYt+HcsvCXUvYCWjhJYb+0Eu8iNS+PdbcZhd+jcEQ+gI+IDk84/2tdHPTKO//jWR
o+CdkIW+4UOkFTMkPaXXGxSa4ck1kITb5tP8l573/ltlRh7MT5gTC1noxOtqJ4Rs
sRiC5hOLXPT7ELoG3SZljykzHG5wkHvXNgBwBUIOXEpTi9nrMG3ylDErzakKpGCY
LcFgIbvZkrKX8Cjz1N6kZ458+es8iGQmSbMxOikaf5KaZhxpdvuPANbSiJTl6YQ6
mxEwqSEOAW6zkrWu0qZwhmnKmZVBa01YLLErI79snfwDkcgbCYthhNbHw/kkTdLa
Hc3hMA+GpR1YnvQszZjn2gXpOwSok0sjrtDOwi8XEKY3FWibzCZhlTXVzZdh912T
01POmpQ3l1TYmBGKDVhFBdnUI8VY5QYrubQUu3hlYGGN95q/YqPdJeg6z+Ift/A/
hoQXVq/PBtfX144so9TdhrH2Rfpx9fOty/mGwOXdEmRXur44i7BEn0p9yrryBw4/
TQptMkl4QxVNGpyt9jlUVxjyByHWkCmK4CxdWIlFsXsaDX54zB0vIdGJp28NX/Yt
Wr7me6IqFo7Yx5QQea80Ig3+Q5IXcZqoOFdHksOOdm2P4nfWAGIY3HAxt8PRtDnk
GSuMLNUDVVbUwVpLmprsG0oz9L16lggzYqat45v6jdMXPITfdzyDX0amXzspoVNg
kNReX9JW8mcMGCP59f+YgmItnOykJ5azErELTEhbKKYq3N+lvKLSLWhyc65ZRTZt
8a3PRT3tU6jZFstUiM1Vsfz8rNE3O62rTyaSSNgrolYgR0TFdijmTm+JgG2hnvSG
8axbL3YE5wiu7MkHZVypjtDiGAIBjLNSIaDN/SOhAmI3xOIETsG4cpVddsYtWzxz
LsDMG+qilaBeaIh8P8mtp7p7PIRk3l8cQog335MiuHfWoycE/gBnxLKn1pTjUUer
/NbMDmeTzlFFRtx3rjTjme2Wrz/BIgZIJXbULgOAS6LfVtAho7f8Q13Piu9Bu65m
iLOStKJ/OaV5XFS3cyfQJJGQi9n13PrgC2ucwFjwAksGwcWvhipB1XXGn0o9faYW
v9sosuQQ54Ebqgw0wqQ5dtZ4lE2GWEfccpkQ/GhkmUs5T835foeN4dSsEphmIbIA
v93vP85FqfJW3aglVzD9i5MywJ1EW8dS9ENmYyzlCaLDSIG2qkvYP91yeRlLpwxr
bcj4A5I2hrFu7f7GRsJAAyPFcGJ0TWscvT9lps9tbxj9cnEGF4enInJKlw7O5yej
BIbXr5pLCHzdwyPyZatpC3MdZ+DtXLB9r5gZJSBNQT0ZjKCkVKmKLat2liYlgwGc
bFq1uLpbQhjTNoULKvTErEmP2DImyzBxKJMsGUojhQEvQtlwqKdjak3XyomXQBeV
3qqIFkZFPE2yIFJhwFNt/jEy4TRxZsLlNHsxgL+3UL02TMfMhof8/g4a85+TdyoG
YRGMcnZsGK01lBGDZ5ZlUby+mLahPD5n5pqE6rRmPwAgrprpqykaLSQhHGTCmtzX
237+yG+GyhRXOdgvhSakJH1Rg5HXQRU0zK0d4gmPSwey4Zr+YZdzP52+vEQtgJ2l
7exPF8/r41HlCr3YNaZdCZThg0Kq5bmQfy/h0QYjPGAlOgipxRzZZyciCA1a9sTE
GPjf42khTaqVQCbhLtRye1It50GZtdJQZ9j7IlOO6zpAFZNUsMzBfuJaozIit0Z1
scS+UtErHSQU714OnWThkUMwa2NqqkqmrEcp6uE55h0bzyLlF5kUwbl6D0w1iJ5E
Q0v4W8M/XFFkksbekS95Sq6ZiFGNESu97SBfC/M629KiNkuJdz2sAGTaCnjKcyFJ
SCPrGcvB+iNOVGq3RVg1F8oAD3t7D2cEqxcTqiA9WSIHObyKjSlCZuHZHgAZVwwt
c7w4CNstcv7O1WammSfbXLIhjaoyf9GBpl2mFzcZKxiTfy7urm/CEWnaM3eRnJq5
WUBozaytltORCp32+RtqEkkcC0RoNPNq+rSwGIUUNZUjaM6gdLH+k8GIsU+J8BHl
ccSE5uuk5D4Epp/s3gGySFsP926cvzU6MdjkD4DWBFIFCj2P9yPWxKm2UzKGAFhm
Ul6yWfbRM234kQKFj3nfUT18oNWE05IPfF8TVjG4pIIijj0I+A31CimK0nZyCde4
It76ncEUWMUyws0ehaaFPqRB84fuHszo1/EjZxmQBYkMqUO77ZsthNo0W14Cywiv
56LL487dUr/W/a7rpCjTUhfbomaO81J/vwzt0qVSAHv7GTZHm8P+tQ5a/mTqO/eO
2xN34pljChtb3QX5YdavRrt0cSTsYcWSZ7kYQ9mLJjS6p4s3varr8AthihvBj3rO
BOUb9y5adAZX8YUb+5booIZm5hr2roj/yxe3WXZAgdpgF35gkDTlPO4USrneM0pX
UEOSdiXZNBSyxIEEYAvhpA0g2nAXE2MNAnvP1EFhs0SQWDTEu18alK+a8pIcj381
NkorlZScIfKl4WeyQ9+oFbIblpguuEZgdlsQ2MwaJPtseovPnxq3yT1f0JPf/0MU
lhudS9q4YJ4sLOgijQVeyWmwBOtfINzFMZjOD6Qo0OkAbpS/2PuoHVAxFqJcyLwG
fpcVbhAhqgOSFHs9RUdU/iLWEWQMrqnHchYCP2R1H209dBCvNQTtLbyzRtW/Jkvv
6Mwu46muRscUO9qfAExeZrmkY1hwXxTwgh1qHaGiWFrUAY6U+GgwShxWLpolfYKH
cJqUH9ZjtmVJs6eMMqJcIPBbs1SfSV3u8+ZF6y83le3ojb8ccviq5UT2MRHd/dO/
Cfh3PHf8onQma6c3mIduppSB+NT01Z3DMKad7bRKHMfaOjX3992+EuDtAiNNgVFQ
/qhvb84B4pkA0omQ3XAXnuQwlU74FEdGxvSxKXrqMwMTzDk2Ugvu1hSkTyHxom3h
MzTVuJOyJRPcwbt7AIUfEfYkD6CALJHbMg94mDKlQ53FAimomfQMgDTXwggkTeH7
cXvo7F1QmB9cw9uYKWo0spwDaaM0j8Z9KNZfA2Vke9gJ1lbqrlMlpE6TgNG/d+NN
988WYSHTmcocoO5k4BcSO5H89DPr3+b5/vY+AGPKcy2wgNaBdNZecKJV/xKLA2Dl
HkB0BCj8kuGSaonh8IA+cdxNnzsKlJXgatL5ELXWPL1yfL5tPp0Wpa6BnaOXDwXO
4+bWtB9WOgCmCZsCX+l7TY5dwtvhKE2m/nOCrekZMO4mBlO427N5JjoeMCjD5VxA
JKt223/vkv1mq+TSi5FeE6GE+/VpbEWQvjWUBLHw7kznwG/4FFNOVOx6kwARopNX
Wu+bhmIQa5UL6jLS+YIRmzSHniKxov9CG3mn9bMbo55182ZPMRxtt67pRavYbjdG
piIqq4kohfZys9b7KhFB1kxbVcdqKCCM0qpHTSsAel3LtqfRWiwnGRxna/7llCf2
dRYf7su5kdwf1OoZr2DHyoSVK+5md9VpwrtvPXXbs1mQxt89kVlPbKQVj9QORvpb
URLxdsqO8oR9OczJyiSdKG119U4Hcr5GX/1RWIa+XEZCqzwkiwKDf8upDxC7pDOZ
ffvzp5NQfUaEnCPxOpVcCBLWOE/5K+lWZcXWc7RanfgcKlG/ON9drReC4vjKZ0do
XHgHhcldFsl6K6Zspcnu0QJlV1LEXayKNAWvHcWZOYHTM4uyVDeG2Zb0e59KHTkk
i5/uDfxi5D1Wohpp42SFgcE+ErQNeywX5FYJbFrx+PrDEU4dZGv7nlrvtx9YY4n9
Z8tLStf9V2OzOpaKILKv3z2Mp4eB6LpXMWGMnHfq4ww0Dvv4yGUSo4x9ErRevBVc
7I+M1BxQCtSc5fGfBFCODiosU+iNDsSnDXwj4h+XjG+Bxo9KwkqWQJKCYCdkDOFM
J+efZKyTJF4rCZEX4U36kEJf8egT22UvL4VY/rfGsNzytfyz4upy0u8BlAWmEiOh
vOq6DWcH/EEBN15KT8lmGZt/avp9PTE35id6pIuAusuF3K3NpLRMe39J8mxIuAvw
dW3iIXSP7QFZ3lOnlta4mx0YxpW6tl+o2ZZaE1WdpZcDjzmkvDTlL+Wczd45apkm
5BtLVfpZMnUyYezmr/W8rfCmQDIiyBj5EM4jyvU3izYGxkFel2V/l1IUcgj86trS
GIlDZjNeahDaSZUQcgUWBf2kPvf3wWW347ogj5YMmflYn6xPRxJZ2GQSKQpFfHPF
bVWfPUY4iNufifgOiLSTIuz0V98ZeQL27s7Qu4kNyzpoV7z+/44ASAqsWTsXsE0j
Z1wmZ4r++x4cZniYhWwa3oabpqTX+SNFDKRaWIv43FH2hLXvUvpeQWvYecPApo2V
AqPsNZBPVE8Owm4IdxHyjkfjEOie+7FFLkZs47eb11VF42xchkg+FHx5jOP7DYfD
oJl+7U7ujZhBVUr/T/Xxat0tEMvUxeP3AGXo8uw8pSNRuAoeeOiWCgmNmrUtYfT3
OuqkvRZIGCN+HuLYdhevD1+0XWwzvtr+MQVhWpl+gERqzDtL2v3dot2DJu56uWUq
zsKwF+iZlrQX0auv0JO6xaAqcl7tJ3UYLA/OXJwH3JLH/MEnOkBCBpRLxRAftknb
uxdGgV2won3Wyy5bx/YnEyultB/zcJ+9lsGqTqgwfGBpSXfqE/W3B5JRx4quPRIt
1Wf7u/8XmdK7AFeggL8ZGyBrE/d6d8KZgqrO+36yk4bqYoEW3kWWsCLmFCGuxl9K
07fnXFTj8YyTMKHdH+OIMeZFttfpHnBP6r3gImF2b5g5XRK6AFLDz49Ppq/O2gg7
elkQb2XVFUyzNeF0CCzhvCPZkk9ADiUprRrM5vkg0bCpDDNclK5VYTkzOmCNit4n
7A14yS7/e3Bdpa2JYwi49i0G/PTehlK5cwVxr68S7iV4+xZ/w32ZJY7XJyqXqK/A
A26RPNPxHpa71SMMNS5b0QQEEFX6UTKH9kREixpLdvD9A1089RAAwHjK7Gd4FgRT
YAR/aDthlMc/TP6YRs9gkmKmB1uodpFVxb++1VU6q3I=
`protect end_protected