`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2048 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
XDmUU01KuyTGZ0KfD/yCU7ha5+nWkhQVGOk5EJ97rMJAluHRkwqgIjHxd/A5klQd
B4ldztEV4yIsWOeL6Oh4XZcEYZ3CMEdYYIkfvu7qoapJndy4Ag7PvbG3chbnvDV/
X7CyqCflpwRJkecAU10HVjHWFpGaoMzrzXk3n4e7NAi4uN6/woWiFXUa4gs1Rota
RYzH/jO/Xb9KyZKdYY00adLVUrlUAO5DpVjZLfH7P7YxpnvdMPf818H2XNnUlF3z
jyP6eCoJABtYq/PixS0aOcGMoKfTWIkKKbB09bOU57wF++Lg7/xKDexrodBDkqwr
QFaC1xWGbJSj2aTzm1y1FP6N7/kzeqEeiV7oUgdihb3ldA3koH5v/6VhV8em4Ocm
rceQD/tu6QMuU4w4BP6C31lijZJ1YQ1GYAV/TyqGT7ZNbqU3Pm2tUgwLODLInOop
egTSMvmeliJoH6jSp+IGLdtu9A3coq8Axz4/EBvEgogWyv3cJjmnAeSVUtE2HKdZ
6dg3WHwdv2jBIDKz9w+vJ4BVh2L115nrz8ul/Pm3+eGVWu+IW+6i+DJSoSUY5i42
Pp/0AVjX0Ptokkaeeo1yy1bGrAke5gm7Y1fH5xi+ZH5rcyP4dSio+xYKg7qInIM4
XfTiSSSuL5sAh2psawfdbogm7a0oAh+01mCNd5Xk1kza9Tz9jR4l5YUOH4uyjaE5
R6i8EA7FIkA1IYIPVfazVnnbQzyjK/dM0Qt85ua62mPpnUKT5vnytGy37D37WY0Y
g7TmRNANNJHm4ifA6+2+cbK8n/BXiVGttwzApsMod4Uj1A9X9hkpVwKGI+qxC0He
2Oh3kQk4JA3cAHSWokIK8zTDXi3EvgBPBGlvxHaZocbkw32w0BGeVXBr/tuqVxmy
eTaR8mCqKQMQNu+hAzS9/0R1+E3iUVBTf8Mq+I12SGRx2xCfZ0wwLd/xc9YxGcqa
8+RDtpNX1F4GHtp36WhHF4BAMN9lPmme/IAbqfzDuPj1eE6S24YjyZKEHGaee3Tw
c6biTosvNQfE1A7CbakzVeJEn4S0haGvevcOr6AIuuPcYS+Do3yZe0C0FVeqo1r3
ljubZ/83j+h9bNNi/sx8D4AyYaz6zOHZ+Q5uyMfv1bRNwUC15KYAKRCER+f0ysrw
yCzFc5P/40/JUzlPlwJYIQaQlPB59+1zSvJ8o6DE9aZUwhKEJX03SaVJQrN7B2Ri
1S1TGmKl02g03Q+aEBQvwQOCEmqsutmOFupT02P9znnxW2MipVna5AdOUFUeIqPf
lHeMwVk4BzfTGuHPaVOaK5lEdQUyWo0t+Mno0yzpAw5q1RFPuTd8Jq0MFJosJBw6
ElriLWdt38FbgdlRVMNNU+XvgmwixoQZ5d1NWO1JMS1FYaXjhn3xn+Pjy4DcfPOq
d7AZ5toNaQC3llJYd9PiDzjwfUIvcE7123uESqX6iIlmMcqXP/2q54A+J3I7tIVy
RxOPXcv1e3i4AVK5/i1+Qf/R0ksCY8hr1YQwVXw+Kf6GsPDYNFuTtm3eyzOxlEaU
zxVLCcbuY6pMUhQryB1UBioonSOcOgCpxLQLHMhLonmstwCfm6f0NZ4VMdN/OnV8
lO5APTcdRhBII1WNQXtw0dC0oahX5VfyYcSV7TUxhsenyhIUqsVPxWWfPqYqxVeW
s/rmpKWwRBFzxQGE4BqkhEpIo7vgFha9pfecOjnpoN5bJ1DfpbObJRoQtLc3P9G2
85zdILPxGBDus+HxtGXFOVkakcVgRWIep6VDdnJpHghs7lX2D7uwzdqfnJSfhFkZ
UYwTxNi0Tvxy5m+lGQbegkyOogINNxI5soFyo1p/bsLLfB4OigSTKgBAj9p95udB
3siY63BoL2oUd4sr6AsGUf4ZP1GtH4k1593wPerPsn9n78jRTZSFILUPsZSTDL8H
M/qI74GrSk0B/HVZQqChR7Val2MimnmR3nLz4Sq+ooJaj2My1AYTomzvIl9q3g+9
wJOj29uv4xmjJj06shqYwkLsK/p6SI9tYJpEPSR1x+NFirvAV8gGGrdkPsNrj9Y7
58za0TUx9MCKDTihEkdUknUNp52L0QDirjlO9Lu7S8wbJf2/L3vx779i2rwfbfRY
MMHn3IprmXg+uEBowgfr9wuyPdCD6wvUiJN8yVIR3zjv/DQKGCFyByGzPhf/0Hv2
ZJ2rE6L0qVjAHYoDXK072AxYZ8xpDbGcJtF+WUt1uhzoAUlzCcZmFc1QNLSLq5Ad
jqRhD3UfxMTq01tfJN8DuzuqGHIjpFI3Hpq89YUfx7QZ7YvyVNv3UYolHwPOb3dM
MWePAGSjCw9D1NL89xddJaII7NJ8ZHO3/7gYpZCfkEsp/oPc7UnbTKvTJP1P17Go
UVbyf51O8ICbE/0kyhrGFWThC68h5xwHUObj526Pg1H6JqvDJ5FeIGa+spjpj1Mt
UGXQ3/Ea/Qw8Za85ZNOqtKfuLt3dj14cybv15iYf1zv9On1c3YBikeqTFqQfqFUr
QklObPlKeAe05Q8jyMRk7kVZ6oOC4mC/JcngPcE+91IWGoTbPi2UEQb3Hi4v7Hk/
mwFTngRZuGkzdBop0gtdXS9L7nbUZGH2ekovk8jht1Y=
`protect end_protected