`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
YATj3kULTF7Ty4ORuRfFpnT6YIk4rUPRrM74bVTnc4GjdV8oSnW5PtQkMCLOi558
1V+/wvDfc3y0Z8//ksX8sZm3JZWtrxUppw8c14g9Y7owiwp+JumRtO1zuk5xFbe3
0MMnIxxoTKLhyRJtAxElG8sbx8N21OWDGiOk0Xyd5CqAmk9dcOIbxzMjW/wndBXi
maijUdqS+5KiRCM9+Gsp6k/iEAa2LnYTt4WtjkmDD1P5jZKsiMgFck8WOqLymplZ
ml3TTfn1UlLNm/+zD3SFGP0kABAiUT8NK2xBPQ5UzQ6sMFPd/np8iUZ5u4QLTWOZ
hTrU9OSX7lOvRUo8pJ9vPg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="BzW6NOo8eyBw+CxsNNo4wIDxODIsVe0ft0K5tGuSUZw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
DhjJh9S2BY18dG77XPz3hsiSQ73+w0XqfJhD+f+lIDHHVjOB7CfC8ieNRTexgzn1
5W+qoqOEwenoVQtit9u3XViXJSRJ0wfUC5a9axblRNyD2mUbyfH9+f59nWqGkVOh
ieHxkA/DPprM70F3APxk51m7/gNSLICSvbONgLGndWc=
`protect rights_digest_method = "sha256"
`protect end_toolblock="L7NTNW/5Dqy+2kJZXKczEa3js87UJ8H00YWI+92sDHA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 34752 )
`protect data_block
6eHODtGLmq6ccbB074dgNWpdzW45i5jL0Nzx5wwM+RA0eeOHXxEV143NNyQGmZjT
bzHAi/6AyRCB4X9z0c4MjyrZE8GF4crbMH4T59xFHqVrQ4zXCea5w0kG5yvHgpKo
2Lp2o1suKM6LQKudLJWunzaBH/GeJq1TUjUqUflVU08tJsc8e8lBC3O7Hrp7HnUO
9AHxgLS0cu+JXiiCSbJSuT34JDHAOc6W1URjcNP9wocDzWYt1hd+nrZjdSqpuWw6
MZN+QHKPg6JVZFqDXNVCPgT0DzaxbnhmXqN0mB76p+TxbmGZVco4V3p8ZX/8zHtA
Bcyy2zZexo4MqJ+chJh0Rak0hFyYWo0CqK3frZOQE9fRIkfWp7KitzS7tamSAwGQ
cicPU40OZxEDVdJC1vFYmn5XlBYxr7SX3zuod9PFnM45VFLvBmKpss5Q6MPAN0Sr
aQpnSk4XMMWB6RV+Qvoxs2Fk5DBViWGaMynHAjn+vi9nvfBiMqAyJirsDCEmGzhK
LVnh0v5lEYKfVWX+cO2+XkhTgeHJy7JeMv/g2S2FNGicgkW+TLOH54srPusD0Enm
OMcxr4LZHBFpGSxIWLNE/FhRhcpGISd0Dro5zwBevaLWEagZ5npos5FSGkrfY+dI
CsmZdwgRfVFLoIvVy2sWKEqzYlqNqoOiM7cUjUVNZ24ImHkcIYwt8f01ITEDYCGx
aEFIH9U2sg4H6Ktx5qYBsSiuaUA3jOTmCMzXVF1V0h3hErU87ORA3YnUqkybO8vx
r3aBZIuf+QUHrkia7LVot9O8YHQl7QsGEo1nOVgwfKNrIdlZJxwKj1l+GWOXVPuR
K/YGM/sIOS4V6MiLI18FR09Vb4OCKWbptT4VqBiKnyCTIueRqiSXaozNB4Cy7RDv
mCHKN5owsx8Qu5qEANc+xSLcBf2JC974N4jw5ItVo2P8PUGjZJ+xBmvWW0CpBB+E
xOci8qdDkUSsFqZP5oeljp2cHWEs6Y97r0VKL9UpLqt3/k1X1wc46mH9aGyatoBE
MnK/liL10zxn/bT1k8Ye5iPLSL3NK+mAwbPKBATeWGT4enccPUG8nJB8tGATz357
/BrF6afWsuILxOaiXL+vHme+SMSF/wQc2S2cvtipHyE4FzS+kOZm0L756Jgfl6pS
GVoan2DGaur3A0pu5xalIwMMVIaxcV0E38zKFuaXTAA6COOvuI7GJzrMW72ppO1U
qZODdLoboH8JVLWSpqKpCOFDX4JG3ZKxsjAnZ6WwvCXx9JmUFOhYuw47YY+SjZrI
5lJrle7gDZNwl/pEPgSQBTBnMU+M9WnmmTYdc0+SZZ8T7Ezg13KF4RyUQm5FdAop
PWubwjCIKhAv0HtES5V4armUr/dlPQ52UH8S2yOirmYqhNx1vHKKYMwAC7KXBqIo
TxdqOoE83uyyFKGLf9zOGa79kTJ9jzPZgvEhgsDFoMEAvcoqd+ecoQRNM89JDJgS
znqSwLVMa2JxUyUIYuntvkIO+7b3bA87E42r+icy7obc3W+CNUqEhoyqapFQnXIX
GjZL9qgsUDMpE5I7n0pd8FbmfYr0Oar2OosXv5eU/foexbxXPFPOLk6StrUwDHdw
L8fztnUtdcebH+MkYMaZTuZq4dIo8JvDSw2AVOvnPUK0EqkpoqUmqrt5JKYoXMKl
KRyBBJ7zxTBOrw460TXug0HoIGfxLA9bJ0bYJCCnt+huGUczElAVFyOntZocWYjS
rmpMVN9G8tIhvvKwIMSIUpoL1fjJoaN9u+72XZteOZacNEbcsDjBsEBCsby7YAo4
+BTqTgyax3+HZILzH5wTJ20YQ0yAzcFwcReW30qo4e2cowbTZBR1Bx33SjF9ZqsG
7BElV8g7TZGuAma/zsBF5JNZtMELptjjHmytB0deYO0DleAgwWcVhJduwVETcicM
NPAkxI5ySxDD0ThIQO7fTKc7+vVEYyvF1r64+zZrcJUaInxoQhdknZWJHm0WF6Hw
hBPhBHNIvmvMTQuuAuD0EulPS72d6hVyQJpv1tNmEeg/SyO52cIcTnchtb+3/57X
I/z8PIzjEhyI13wwV1+7mtcv/zGPu9A+lKLjrSw+LtI+ZQPcO8q18vNYLo0dQfs8
rJ39r+f4MkQqrvfYl13rvvvTq+b+F6yca1SmfkZ9rS3A8q2S0r8Zx5ftzY+dn3EI
jij4OZEGKtRWXTNntg5H1MByvZCOa0oXp7nQZnAsriHaNLZyRTPeWty5VyrSTPgc
Dnc5eVNxdPTRLv/ftcauFl/jEGWN2KfOBWzHBXUlpGMXpB7VtLBclschqecZXqIr
J971eInfpUNFzVoBdIeeOqqqXBm3p7sykDVftwlIZmiaVrJHIAoYY9QIN5pu1/BR
t+M3Sl+2zt/ctn44cBgDCMchOeTYPqboaidlmKCWbOZARt+vUTwsZgsKI4ae9YzZ
QXw1w9FH8mfVR2qznOnnOdntvjlu0EX1U4EYxglxMW0D+PPRBnrcRubipM0FGrOW
TGhFi6csJnIe7miM/+ekbrhH7e5vzYRtfPUI7+Tf80e4TaRrvhO1agcQiuR7sMY3
XH0t4EOORO/8LwUV+SGSHB06EawEsiKcjOWsN8zE17UF5duhW7J1vpXV1f6ku1fw
Ry2Bk8gGVDgQWUpjivvIlMvqGuE0PgvCDBUyYiCfgaKx7tmuEq2CLbMMeXDghRfJ
Bi6eatjyqqYe8HtOElqpMuuUc4SEqhlkmPQpWtSrI3QVSj+zT7DXcBYyR0a9heSP
yeqpOBRv4fzDJ3jMGfHHdyQa/0OUz4zA3jHUvzSt0lhfp4sVodLOh+RoREEC0KXp
PmmcGXp7QswW8caNazC4ooUQ8bNhq1uNmDV9R5GFuiKZdpsIH9RBOWD63d4S3s+d
fCh40dAuHXvicg9ocl0Zh1HUqErvxKh2uCSW2QY15sz6+8k5VL3YbJwXRAcWk3db
o+XcNHzjZGXrFe/IUc+mKmJbJdVI0POlp5284RcIT3jzEDjHoooMV5EcxX2d3raA
m8BH1qMUYHDNeZlbnJ7K7u9h0QfzNC0WqNfIf2s0wjPhaYHf57sojpOHPqBs/An5
ZEc7X1WjXYpu85aXyHHUB+Blfb8PvlbYS6XrOc6oWPSlmK8LSXJPzIgE4adGwrZQ
TRCSa6I02iQwgbV1QLawRwGC/MiFJhM949EiXCcD4zB6/nK4mNbMfYbh7lntqJFh
zVq9Kn32xQB+xAWHuHnrxHgQ430ANNL9UK8HEHijXDjJn0R0G+GDmbQTB4bU9sut
BYnaSEWQUQC8GTUcoytcTrZgUuK0YV4rcOV6GXzzG0OOiKVrZ1RXtMeGUL1y517X
TUAQQu4V5mfBxB6ET+Vy3d7JI4Kf6nZLeR2Amit4L90N5o7Iz5soC+aWr8QwMX2w
VWbrIPHl9KQWj3C/e56Qf1Bs6h/ZmYwKR9bNUs+okxVeLa/eCjzMmDtq7MQpsQ3K
Zg/nI+yLFw6wwDb9o2wja3e7+gfG5W1YGEt3GBY23H6iZ2Iv3Z+ef3mpgSvLBZvZ
PsgjVW9D0v7Bkye5ENlL9KaDZxd3aLWwZGSwyb17asal7jgqomqsL8OcSpWltLmF
nl6oKetV8S2vnYuCj32S8hKKggt1WM1DkRHSeMgiPBtEax6jjQf6tcB0SeZGQYaB
A2Zb8nvBv+3HtimriFBIMXAov1oD+p1sVFTq4OD0Grsks9NCwS+5mNxIMkOoTVT+
NiOTt5xtIoqiTAgRw9vl0pdHsytRzReYoc9EiXWQOcPy2kQeef914tNpo3qy5xxt
ThFJS1/ghGWhbZspCTZvmvkN6KjYal+JokHlNQ8qUFWI47YzYeVU3W400sMCuUCQ
thTUd08jyGr2LC2ohgNc49+l1TqO9qmI0aiNbG1gaUel7jod460l9bJ8sNKKGvOe
jKyAqbxgbtiAQ5R1GnTHYV320u2xDFqtkREJUA9HFfoH7AvDTOPv4NwEpg++BSvK
gFqedWFxekAHDp4afpXcmJmgnXgjQkkEFMMN55eDmlq7ANwT+v13wdy8qDctYxLf
e94Al6qoxNYT7j3clMCY4w7rKrG5ikv1dxX5ctc8Usnjve2GmGwGrHTXB0+nNrlm
KhZ6OncxR6RoC3xJu7cx8BUTBuo6/lzFod2gLdzANKW5ohSUrrwPvKn87HngYti9
xT20REGnApGQuHiUap2nV6KRcSN309mWXCb8Syhs9+70JKf5caDlYqwoxXfc+ucO
Pmawp+MfGWvr84WUWIgRwJ+5DcO08IM5JOI4cAev+6g18FKT52oUALojCxmvxZo/
5OqWGGmUPHjA6ToN/llXmvBTKtC6BxF8hdhH1gt1HnaHkwEl7hCUo1+Q6tRiIPXf
84PZ5DfL0znyzjuqx74l9OkSagzbs21H0tOQBUP29MzcohQUSChEHhKkuIO6lilT
1C14rxs1Kep1EUqvtoIONt6zpj6mH25mS8579IB2PyygzpF+cx6lEZdIRfiI19Ir
mOPrprZ3M+J47FZhWFAeXJZNRjJmPDfySTPrxc0yI3Fwpo0WYHOnXpmCdp+Eit+o
CmDGNXDsKCYfWepyjCJY9V2oWhR1C4w8r1P8CN7FG4HMfqG+S24ASizQGXaajzC5
aKwNdRsta95HYhnE6Q60K8PevB2f2C73j8myawGnyLWTn06b4MA28oyRQSBycIo8
3lrs43Ngm2QmhiDdtQiHKpsGPsaEVyNU2Ffojkyvl8jb1i/9N+AVJD2RJPIrjdjG
M1ABqb/48uB2mGbHVKhSfMiXRgJwvLr4yoO1Bqh2D7R95hVXucZP7/VNtJ9y9PgQ
bhjBanUlDF1DaiJxLm2lae2vkcVRGATUDPmE8i9a2TTryXXfDZnjQuGgPFJYWL0n
Jgv6uX/2lLN8psMq0KvXgQ8bt7+CePzYesmiN3hhaKwKPNsaDjRkSk92zz8Ct4y/
DHjt/i9zRN5HII1vNrodIVfkIFeeS1luNuZKkkJaXlV8KZ5jQGFPEQLDN0j4dEJT
RPSeq1/b/ky9KpNdgsQ9YGGt1ld3zZtWQ1Ezf6JNBe1rYaq4Nzaz4cUWDpGXIboE
Zyd/RU82GzlZSfsCmG5EE3FCAW90da9IhqKtmTkBj14DmvT4qJcQBU5ERcPXnRMg
ZCAjdxard2loSq/RDBqZ69Bo5SzLPdnHzMenvtOeoY4wnzVBc7x3SZUOAo1NJtHe
1+CieYNEnXjWiaFdWW6RNc1BxwRRBzCr6MU7kB7EIiabCvJn3qQuzmROGpvgFITh
Q5kpITldOwLzrJTHLDuKdVBEL5JD1EW29CVkBQsHwSpteJjPfXxaiHERattgZNfc
OXl9u3uV2fOdmkh4n75rqJkWZ/tUahf7lfmrnXFw5/y66jnf/IU+cRkEAcnV2/ix
nUxLnBIMIsB7hHWJzAhTgXqGHu0NUyoAifUh7vjuEX8E0yHejQGcND07oh+0cHOg
eyWtBJ8HJcjvXTfSs6xPdidJe5i+gy7K2WkMBgO2MCtHG9naXfWKv3my12+PMFtl
s26QVBQinrZtthqOBdp8N6OdlUfus26p7EEnP5+tjPlFG7F2yn3uHCpmTuup0fkB
6YWlUP7vN7c3jkvC3Cc+9pK1YbHD8EUVtL84jv8yU1zQ+wHtvQAO6xHX4CYD2mzj
50BT0XW6Omw3AC7rrB46H9qG49yVtiO6GHlG4kZv6chXABo+H3kIYvXD7SvMEYbN
TOoHmzsPapQce5Cn/Hwia6sZInx7+Oj5UsPUIQ4zjpfJiQx8PQfReLr5v8rDt69c
jqATGwq8zhlr2mMur4vumO6Cwu4dmE4gDYHGdazQndXSo7Vf258nhmc5Wgl7d4Qp
KTZpVgsXAiLQMvlojEp83w93lj7vbkflWWgaPakOPMqDtFvh7ndHttfxftSjvbzp
kh0Np8AMezobzHLKi5zKkvIlCT4eFPgpBOgd+KC852lKxPwO10ULnmCR+fG1vofM
iq6j7j2zY/UWJyIplYfIisISDXs1JBZaxjsCCbwVm214gWbBfByz0m9y7K9UMZix
sSpf6BvOscdDpjK1vRq4GCcNHD4DxJfiCljPyhGNzO3R4RMo2IzJi3mKekOx5WvV
y4NkBBPeFenWtwMocDV5a8WLZCEOG2f/cicfyW21/ecLIMbM2kAKLHilwu3lUKz/
y8q5jzV6MmmQMAzGPIRJ81N9SiuwghYWA19zMpZs1MgPdCF+diz0wW32DblXDIvH
ZAz/ryIKTgvZSzoNcjzsag0KLUTPIIt9hDDBKfuM8YPVzwemZ4vhIjzItWFkqXT8
a+1FSS49lylz14gWshicccU0GKwNfC7SJOXFmYTgslUuhLLcHilmRYFKEUl6NU4x
/mHBp+P1NCc0GGeo9IBJ8+pyWHIjeDBZaCGzyXNzVirCwty2M8YuAa9TJqsf1OC0
Y7Cr1Y4TtAZJk4nQrPmLN+MjyYxCElTQiOCVzWVUzJhnGlikDSQqihj91SayHTpS
sanUbEbPYRUpQQXaE4AqkoU91p4C+7AocpW6GWf7hFez3Tp8emONTAd0F2uIYybi
8IWb0PQPGp8e9Fs0Fp3xJ4euNEczkVuyZDpPCFkYFWQy7UKl9dJE5dv0ZPkyPKME
Ucn6YQif9b2ohR9Ia8psYz5GvtqcHiwc1oGI3xrnTvg2ouRfHgUOA5wTKxNiC7y3
lvp1sH7FcZ436aWRKzSrKTH5/W72BIiyg4WA9IgXh8at/fOBzCnyIe3YqO5zMvQU
kinJ0S6TaC2ENkYRKjbv4bjsJphwMuPgcAHyT/I3Pu3ZyadDAMiFN8SCzW7HyPrM
fpVaZPeECOrvjDylWcm6TQXii2tDkBPDNeGm/mEchhhJbYAAaKoKp1nAtGnv2KnB
yMeS7EGwoW+22+9cM+6QSb+2057wVHT9cRX9LdeDPmTEojqu0dOBb5v1Pv6RAtCP
tMN+IQsXDnHn5dEb2nyiHgmJtwYxzinEN+l740wVe/03pOnVaLhrDGrLhe9H9qrw
8Ul+lzt3bo+iYXmznk4K/1sh134GNnFXynP+8CKV+YqcQFa6+tYHdXyv9Z+ohhSC
18Hxhcx0YVmFA4bkmTvQDq2bWZJBwU+GW+O4c5MmsbANS+NA/Jsq9e8+PyTZ+XOP
wvWnM5ugPtqPGlK/hIN1kji6dt8z6dsty/tqp0ZAYdoSuyt9zDeB+qmz8r1QIcCO
kKY8dVloxY4p9luPM5lFTEX8bzCnVKMxPiTdMhmHon9EFMUlNA7H9+PmhujLfg/a
0ydSOoqFOLzSTA9GcEUGX4UtKhxaocLaENfpj5AqkV4o3LpkDfjYVTbkNGFMFlwz
8+oLStpD86o5VrWnZ5NryiGuA3OISMxKDAewYk3J4UDgh8UgN4CMpg+1a3nwRK8n
rglFhc66T2NpFyK3FGelGiUX4zQrh3hB8LMWwb6rQPwY5m73U6mEOmwtL733Xc8U
/r6sqGn5S8unv9bnBJFTj91eLS3BSEVGouKSmEsvhbjRqNPsVWWH1lY673SuLQM4
bxqJYRlJ3MyDJFFHuQ36wxJ1VbA8YgmUEYo0SWjd645ksGC6kQzOSBirsMFSMoGa
Ng6j0wrBQLf9nSMnwaI/AjpdFTekFdZgfaHz5ylvlM5csTFeDnTBUkk4TW1QoN7n
UEoBI4N85EgrpQmYJz07wz3e8SvGoX2wB6ExkGyCKbHuGF1rPsGFmC5fTkAgspBa
KNc0ao+kIT6OpLhZz87cu3ii8yrsFcrvScRzEUz8orB2LHjnVUWCfo0coxrj9o1x
F4WgaF11CiA2BljZwGipnxDaofLGgND4AWQr8dXrO//SIKA8FmJ5DWeOgTtSctm6
Jqoyf7smh1YVMt4A0pjvvgwLBr/IKWdPd/c1WJFVWF3DIW7C5AZaim3lNpgJ4Rfx
crU+1VVTp+fFNXahD/uz4inu7Dr9dSHqI4qbj4998CH4SJ7BVg10gYSY5Wyc6R5h
hRE547zsVbnDzAkR248t2ZKdTX5ZBqUxLTVL/2NoCp4JNBGefXfQQOegvxM2U+lq
GPXH1yrZuJzuYxOVdYDgBexkR+mdoU9HKhVVrkl3TcOYif9cA7d929wrE5QX8ddk
ICEuxE71v8eEqJz0sZMObpEfXPtLlImXZ9wUSGmG2g4/Y1fyk4I/F7T4kCZkfAx6
fkX5p5staaDlFXJCsvHGFBO3kYg2XHrD+bTZLVcLVmxN2u1CBxEgE4YNCxd0PuD7
WPPZC7RTzLx6rTD+wZhvqQabGwb6r0+D2nWUTfpPciu7BjVdHBULXyefOkWGvBtq
5fDIpV5yBFSRazrYI1m2bscsqt57vBKEua1lHF2K0IsHH19BDqB0eRXFjMMiVDtw
pu3oaHwOYCXXdBKhe3XyBIO0qtE79fJYzt856GSThEWUVnOaMAYWDfCvd+x5PLR9
8mVWNa9CDck2dkmvZY6DzEHocacMwJD1CKuEOmC6BiEbe3t7RcA1cpbjG9nsiEjz
koCKDOn0a+d3IJMJ3SheERp/c8PJMQ80eKo1eqbHstlkd23GV6C1QZpso6m73tIH
tO++51RHrx94ViRTxrYiODgAu9ISbhzgaQ30CFPtmhla1cV/NWfYk35MPq8xxoX0
GOmJxhUraQMU+SvdTRE3bSPU4TWw42g0pX6AUCH9jdhGFrZM/04WE/x9FrKKiT3h
Xg0jP/mr122rJpZ5abCaJdZZ5qtFg8AukPcMaa/Se0pnqsjMx+0XSO7tsEJ5NZdC
PO4HVVMM6qkNJ8n5ay353b5g2S7aVXVZ0vP+GTbqwl3j9FjBT9OJU6TNrWyMuQF+
KC/HRCzpeAO6MUbRjNGtr9HsVPx7tlm899xACv8AVgWYcuQqFn8Ama95+jDl3XAF
gC4qCRL3dPVf5XG0xuyTsRn7dwwnE22VxZANj5hrnVO5jLVqLOykxyJS+ghF1ul/
EKvpCG8UreYovqQZ+AN8pJmXby4XGPYy7FfV25HsfVHkYh9oIcFWKGvykRBzAo24
DUdI8baYCtRBQgBcjL1UqyQCLcBSZKh+IZagVHA0iOf9hvKNGl/B7dvltzBkYx+I
+TTX99gNmEiEZaaHJ4/NquhoJ49/YR8aw/pf9lA6K3KpDdredKDILWqzr2M6MSq8
B7i89dMxx2soKIk8MlTQbro4KYA2sft27Fz7t/2QZYpDltaHefABRv5CxCxqE6VX
BWE2Zc0DP+gr5q19XRVKpYLn01wL+0lGXf/zxXdVBdRhcV+rye2rytdqg1txRpgC
Tllp+wU6sDelIte8bMfCZ2MzHsXdrktJHVGtx+vtiUEmRwsO1df9TUwpyCqcqtTh
8x1+HvVtInMeO/dmKZoiPx5CTKapj8QFhoTSk5BxawGk5Vry1ZVTFmTGLusVJ3gh
n6rkjkI6AIKUtb3Eqv3UqgDbs+ZKPoPjrWlSZfZZNMIxNIZPZC2ETTNXlYrD2jOK
CK6bKqGeGVz13bbzB7wWt9VbWdnq4eVydRzoX2+NZwrNTTjK7tlSKtBtHmtNZyOO
h3jznNc0m3/gBhZaAmAovP9ybniNlrCT5qGwZpyQW9SR7KKp9k97JD5b1obkatZv
p1kMxJSdlCBiwUgY2/Z/6ZAb8SNQjPRuhMKZ/hpHARtMhq2yysD1GXhHyhk2d9ro
s0Fp2i3n4wqu+gQg3Cbe+2XfjIG6Yws5JYTVaPPQeFSzbY0sVH389dPvQvACqAz9
4ociFU51E9NqfeSrKhh88hu05nb4RjzANvJfQUbFImLU1g3CnRmeUp3IUyEbkwvW
Se4Ep0B5KWzlBMzS/N6OhbzPDosc0MYVsIN/WhgxCYU3MMZhJbY2zv2RnpeyKqaA
8kz+5AKw37TCraZ+4MtKaD+ZVdkj2RQL2HSgSQRYgv3qJvimGtCzs6NmT9n/iFU9
AF7CiwzcMjO4qnVy48Q5EPNnW2oO4mDR9xBeHitZzd/ZjskYesCpRmMeZlm0JnxR
8U7jaOzn/ZH0zvTqi05AasbA4fsLMFFOYDiDkOTpjT/ULCUCjEjx1PXnU7Xo4DzD
hxGq8qCr79nkJiQi6eQYqZ7v/DFqgaWkUmd3EO5Tp4xbZiGuUr6DEC7l4Upxe6aO
X4R8weXIaeW9j9WIRn0UDJn/lYMFX0g4Zamh6DdtSMDwx/EeqCtmbYrwEERHxGUU
Rc4XrKLrLlZ7Uhw331zxgKDbG13aXSTDDBV23UjxFPuBp2NDUqhrffncQqLCmRCx
mN3DWfF1Qs/lJiUP//6wA035CNS9SM6eGxpKvuPOW9H3/ovBmOjiyoDaumqs/oHi
VDaKdXagOWeQctI0/1qaEVu871PJUY/kamqh+K7j78p95qP6fk97QvIwlBMxS/Bi
y/rVs5h7UmxfRAbVL4F7mZGfOyoNhJEjfFxYTkxc4SdN72bGh+HcT/opzEO6Ich5
P0GfgbL1bcXFuJbfu6GiAwgLYc2zYfVARsAJtuTzorqct64LRg5F0OwEVLSxFDxs
nwvgDE9yOTvWUTZzWolarW2AsbleeyrFP3Gs0EZyESo4whE5ZZZRzgM9TI6oXv4D
MwNicnS677XNMas8m99SdnDzrpAYIoq/AfViQozZBtfiaMFgR1rEWKcRJcRMlavP
luNYuyMutfi4H06ReXWn74fbdHIwOtaNjlQpvhEIfBg4dbWiBSWNAucNF4JRXJT9
8+venUhmHPfc/T40kGqjQH/3c2TeD5gTFudpSkUB8AFXy9ZgwTdwca8dpYIDY3WA
KEmR9Hs+qpMIWY5g6OcRo91vHSQ1BJIlzRku4gqEAY/kGHNKW3f5ICbNewdgD4Bo
ga0/XOgVl2Sh79BezozCxLmguOtFKaevKuigRS20N8Bnl2zQE4T3AhGjPdkoFJMW
gTv0IXy9kgVp1lSKGOIAwwVWkXWyvCjuvZtiOlzUBT4iXKxL4SyEoHV452+IRFu6
uSsbGWsftRgMzKFT7pchKn7JhN7dDjedsUMNIwxoH50syjY/m09HLbauDDcMP+u2
gvLYonLtQeASpbnZgjTTfVXCUXCSJT/qGr9rDM4Q6EGyRmsx2Pbi5/Tw1dWZlY0e
qPtCyiiT4C1NJ/SEN5nRZ2uYouTgknDY7wr8A0Hmd6Jd5n+T1QP5nChgWpQfpdVo
nSnuB4lQhovS9GEqwH28xSkoKkwfwGtLNb06rK2LBwrqhuWX3oMTJQO15gWr5wU5
V4JFagwah2Kj/6/qDpXUCA+A0auwIsT/BIE6tIKzPYIA4ki2cCu1HAviWxZmAou2
nGNG6q7bkLIi4+U35BtOVJmkjArqsZfWH+ZItfHJyuBm/YWhs4kJT0KAQ2AU0uQU
eVE5BU7ywnzomcycyCpDuHwM6nAhf+e7AlcrLUyj0euwQucOmfVtUKuC0pO2HoO+
bpZiCEkgzhktffq/LHrwak5NDR0G5KE9Dr1+07kbrsEVbdrh43Uo3PuupAwLD5UX
ylMwsg8HlleRVomq3zP9w8A5MTlHyK481ZV79nBf2E0uLHkISqc1e4/Ifsccc5eB
a+6IBjyPm0MEVha9lEHmc8S+SmtVR5JvefTXD41ygQo7S2/9GaFTkD0ALuGCzinL
QmCji06//tFldjMLCVzv5asKq70YqWYhaizeVuUPkg1t1xZr/Q0Oce6/JQgYFcBI
Nyo8ac315YPcZmWCPltUaIWSx+paeSkL7ZKdaJjQVyyUiOl9aNXozZzWfIrechFH
9JJ2HL1GIbMBh7D6Hpj58/6DXP1NiJg7wYLeatm0uu3WxS4O34BgGy+Q/A0z7eEs
I4kar54jZA2P+7NH0TxbT/1CkdqHhBtMfqs4TysLF1YIpz/pq2npcuYR8gak7k+w
b5tP8KR2y6zMB1EBxi2DcJ7sbeWxFN5aBFx35iGt8EpGB1fE3xMuozpYK/IekuK8
tyLf/ZEAkvZry/pYk6XxTwi829um7W94DdEfyfkNZwpxaYighljZJtDzk0sJVilR
4wVMC5F3rf/7v9hWPlqg9K1+DftFrqEw5EH8D1vZGqCYDToJsl9/JAQKITFZW419
1MakknQOiSzQY+90+2GZ/+onDBDnyibysyV2fHnc9yirCr83bng2XfeTga1voh6I
vAbQZ7ypX1iMhx2xirkh0MT5ibcxF8zQECqE+aPLK1FiYhR8O3IJXu8POLIqsPt+
LXdup3Hd1p25tjAE6Ge8lHSZB6AAr6omGCgxQ3lQ1E4gZ4lYQodB1+cqR1XgPxCe
Is+hjqMtt/7cMXLsqaUX0rSLSYqifnQeTndFg1/7eOCBfU6Rx+1Zb0l8YqbL/pA3
iU9t+F4AAtZ5RzRl5+X21zoje7w/3s70u8zNc9vRe7B9J0+EL+5oHZTOosLcW2hg
yVzj7RlFvRm1OTM8SOe8Y1uDLZOom8GWyw5GXuZBfoyJME5Oahmx4sUjtTsEIu48
saYIapIO4sdcKmP3A4GXIWjPyd+Pu48rKR/mzaKULvn2AbLtSqtxLqzsvcYF9XHU
UnYx5Gjz6SaTGq+oXQiAGTsp34IZIVz4RMgAzzA4zpoYmiFu1qF8YaxbCICEWJT6
RCWWwZyanChdorCvc3BFdENJmy2sbujCm/EBF5lUp0xOR6pBITbLNA73g0qN9bdb
yDFx1hNPlrz+/IJg2EcumVSffLk7PG62MR0WEqa+TV7EWUmmkKIA99kUFe10rZoG
yxTIstOEnx6wF4umnnw07p3+QR14Nu336puEAEJBFmKgsS1GS2gqrxn5HJc5sGOo
guqUaaboxfsVaVuKAYGHOafILyAqE3PyjnjiOGLTTp3UMss9nZ+/bEsN6offsd5P
T1q7Ltf1pFkNFU2cV9ftmdLS0+WhWOI54lmnSwY6dZg7NQTVHIRSkIvHc1p09UBY
3a6826LLZk0wUMtmOtk6nqEbkXxOFHv7vkqaRUsorLR6nRJHa53d2Tb7cPREWnfC
sS6bMXt84YRmwJnvXlwdLvXSxtEGKm5nwRCajXlOkZyZyOqCqHj1DR1xchiTkAFi
exHc+hwEZAjzcY3uBaaryU485ZSH2eUMpROELlpDtxF3u8T1YZbKWt7WO+XEpynb
b++q5Z7uSL9AGUTIyRvqDoyBwdEFD3sMKxZYLmXtWQcsWNxv884ZACLv25841NIo
KEKjNE82X8gfyyTfUmpt1C7JigqqO7zD53Ht8HGNqFSv8LTCG8ykR/nkhtPKxCoF
IfFkYgdTba5DB5D1WfEnYZ22hQj0v1ajE5pzCJ0jQG1lSTXgQuao5o8U866iVDM0
dt5RTS3iMz/PPUmF48doIE1kh3YH0J3VNUmOOlSoiCkM0beezN1ItLxD9T0Xddx1
JX7YdZOy4pz3EujAHeHcCEQHWhnLsq1D9SbFalciZx4tgXXmjiQoEtlQRf3w2Vdi
KCrbZ2tD7Pz8SkMhEEWuCb3kKB5du18viN/jXoR8uLLRrdX0a3OeD5wNbBWDlkA1
+Qwl7o435xJXnYSWZMAdxntg5ReSVM5hqm6cMJKOP0dQY6Ff+W7AKzYe+5ghS/G2
P2+WrH+fP4HFeEngdBJ7xbh0ka10EFRmB0llV8LThQ4/9lSOfnd2JbgLsWkjsoa9
nB42HoicIkdTItwsbDGNpfHqdSXlG2T0eKCZusuJWGYn/h4IW7keXPvcozuTHRAQ
lsXU964gjX21nl6CD8BUo7ODY1U3d1byjDE5/TBAauX7rSDSzBWLWDWFziXIaq4U
TE3KD+pMl4s2ZAGKcoxwF+loRtMKVvFXEgF96qnIvmC5zji2Do9vf0MBgfPrnf6j
loX544rCtL+eJcGRDhir4cc/dMFiT3lixThSVnrdIO8IOIzy8JOwlvFi4m1ntzeP
YJWMeMJG6Qp4206V/rqfxkItM7dNQIMZHTukaF6m+of9fKnnfWxDTe97a6PAxiXh
y/7pd6oj66tPJ6cRSEsNmiYxf2/X8Cx5po0W+sWdJ992aaH9Bn4QOFUuJItsjcA/
Or0bl0Y71u53ZG4vv5XxHIYNUfG1KsBifvTvXj22SU9V+94XHSVJI61pa8GkFaE6
Is/D+oF/3HCZ0Enx0zjU1HL4+oPa+hVAM3BdWbKqQpHWhS0O/Fy5r2AQJI20Ve5+
8v0+B0ulUr2czXJwsiT/XCbkHUcJCEhGcaWtsLMNjaGbTYYDAvFC0V/B9rtzh6qY
9qnKD5Ys4AL4Cifn0KcZLxyc7U4zGjOnxUdtks32fXiaDyq6yVGtALGWQWCg5Pg9
1kgGvO8YOUeh90iltjL3UluDLfCiQ1QzdRoHXdm9z2KaUBCZxsj/GOpa0lL2LErD
+uiP4iNcm0/XQ+y4KY5hhoK3Xp+cO2RpObm3Lv4DA6DMSkxsiyAYh6UuAY6ccydp
/H2WoakpuYKZNE+uMntZxeeqSnt9u+oZCB0pafwutGws3OUiDFp6dMN+7j7I2JST
XQ6qBsrprWtJw3oScxVHppCADpRCR+DStgXkLhUzDq6b/vgHXgm9ANuzHmTj+X4R
MKmQqGAbeEdVyySOtj9i4B7FWxe06KcoQ9fOrsTC0tUSL8MWZab/5s3aIa/azIlJ
6xF4GxShAcI8rUCErGsjK/BHrIUoIVqG8r6gWRQpoxxyNcE0TmehHapIpTBNj0Zv
2HSE6WeRLcGJjZRS6DdGhp71BTHywtTtT6McK0L8cA4t1IjjiYyQZ1K8HKqFZos/
lkxpMyWBFxLHQMHrqGjw2xa8WydMP8IJ0uk8KDa2t/jfuW8GV8wTa1iQ6Lr2W4uV
Z7e4jG5b5MrkFneZKTXs/htfyJCKNHTwAOgWhpR5N+oOCRMaWj6QlqJ/7jN+5Xxo
hz/oVYedH3QVL++l225EZwasagOtP/987cq5fBNdAPgs2AHcCcoqygu0mlHDz1p1
yYWoQZUWGYbDsnn/3ZkVtSBL/K3LqSEW0nxs8cBP1XXDh/45Y5p+twYC9PXgiDKE
g3XAI46y3JJ6pxaj0EgR5pDzo7CCoTxUckn/My/mFUeVZrMmYSwCXE6XseWfUnom
MnerZuc8WV/V2+MsZJF0G+yXNRuLsBWOF7mkW4QGiQNPNoGZrvr+KWuwRx2JOzGd
v8xdQJFGFAf7+O3ubfUN5wx78htouHoDAT9JqdgosYApbUG3BO6HTsWp3cgDSxu+
cMLJOceGcCaNl3lQZPyqxy+iBYUwegEZU+Dp7Ubb9jBhtIE6yMCmp5QDdx5TNIuU
U4IqOZX4T+/5+Ze6C74zAQL3FMeldLxuJs+r1WF4DiyJSzK/rYmnlD97AAPj6cWV
g2s1wjjxyUdNGXIXKyi2kxGN2lhc6xKjN/hhkEN+J7tJAhc18WSF1UgQYTaXMq6K
ShnUcFZx9p7ezqnhq31Fyj/h5fEnnkTEleyEdOJK6F6npSVj6B3AOmg5wCwVaGV8
eaO/wtY/aTii9B+bhb96av7NqMnuiT9m1dfXvDD1vPes+SmNIdYMTT9d84W0ql5h
WGlfIhBo/mYz+AwCR6rSLhbAFXlRQoSnrali/7FsyPYt3TVjSahJI+ZkpSdUq+u9
y2YkVqEq2Kg8MbfZ7TIzuaeEgcYy8W4r5Eoo0ZMrYa2H7QE6Bb4+A1R+vXz2NodG
DowJ7c27uo3GQt22VkPPV8fE1lBKIikPShDPthUZWY4SpxbuDpy4n17Es5G6xrA8
s+enFVCNNMTN1UcaaKruvnF6bmV8NHcol7uMnkSdMY8j2vBqVCg8G47aHYYEN+IM
/5+/Ln86dQXJd86KRutH7Xciua4o6nAK5zQUP/hsmURn6Zn06dt24ZAlqasmSy9A
0qBVZ+h9aK3ljyGYT07Uzpkf+zYHAOzapwJ58QGmWcHgzH9DqcmAMMSXwJ0DVJet
M4qV5/ON5DERZAAKKC71nZuuHN80nh3Bi57rOE9ncYMlcC6MatjnQ1Z5SYPre+Dv
e+NkQiogTcztNFF2a7lULHpDUtcDDwuP5qGvnNt7dckQLFuHOmUkAPTov+84zGiB
2c12aq+6u9dL1dV/vs4j2bEKJs+zxwyz43mWvho0muu5MS3Y2OSViRC7CHhvTgyM
dnaaKsXDgpurjGmfpQ39+mpz2iuW2vi4ZuiFm6FOUFpd8XhszqHjhJNt9T7m9DSw
lAUP2U7GO7/qIXqB9+VS6Wy27QZr0Wf3btmDOKaqv7RHvwKwpjpsQEq2A7Jmu1gf
GHeC181TsSuJLkrj0b+MM2yvKsNJ+hqLQHuEFOxFtDZq0P6xfGr3zPTBgUXS9gRk
R+qRqbRFJ6xE9xz3ywvp0em36cLQI6F0lCCM2xNwn3SBIhy9wSWel//gqR8bdbsU
7XOUl6SWLOy6KU6/Yz0/TCbxO714MG1IMBkEr6sdeeV6GruSbL9zE68Fd02JlRCq
Kaj2WnuzL8dHyqiB9Bhbj607n2otk7OGMmcc/ZDJsRAy9c8mU4TmT1O+H8nRlBkA
u4kRqfYElkDfLYeW33FDL83DboEP7Cnp3vmDS1dtU9DpdLJcBGu/oGZVbzC0Ykz1
/HwQztyDMoWMG6ybT4ZlUFZC9GIwsSMPW/S3AyfnmUQULshnGd84PG02JivLD5y6
0AhTS2vY6+URsexZbDBsWrN0xXznxlp0egVvbJYXN5gge24l10FfpZUTs68V61K0
Mf3VUaU4YYoSCIXvl8CwUlZgZRUQLwIrQzwgYOhy2ow86AfbmESOvLfKUMe0enUz
LN3wqpz9Q9UMGt8ItubQarrH2YKMR59u3NcnNfoJdll1PZDLfT5dPZFbiaeuM6eR
N+PhAbhUHIilYZtIi2CPnCMQUa/fk0SExukXUO5j3QvMfXXf0DgXYVd6KVj0qQdm
HJjqEKYAs8U/IyHzMAvN5pNBv/LHTF1CNdFcHaiM2S4ZKNy05MAIRKxyBxFXI+Ph
6tmXRVHn3JbMA4NiEe6zN43Pev8b9nIFYIvvCFvhc0txmz6TkKfFMdX5KIPB9Xcg
Dnbz06OUIAkKb+ra2dIDyAj3jgmF2YU06UQVdEhqU0sGrbsb805yKC94zxw5UcON
sOWFN0DQ28RwB5FxcFJjcl5C2GmOdDUl4pPudKbK5w60y33yu7qj/l0h5IE161Qi
Fx4E7/CZrUAP478xjdxDrrZmT88vFapyIVHcYrsxu2YCySfOXFXJ3RjTRoejLV/w
/RJ2h64L/nG8C2mf00WXWit47JjJQzMXAyoNFq7Cg177RosNuuXYdYsUyU1Fj6vO
GzwkGcpmCycPXbU1pdIrAjrTAgLcZrDTAEvU1it/TeKr4jFQVM+bsSRiS13540ke
PJrkvSYjIx0aTtHLXuGMPKs84hC2p7Sj/q0CSBo5e+dfHR9pOsWKguOt8Z2bzVTz
XRcLvVAS9xbQwP00f1JhTIz0EGKHEHTCt+8loU6c9YMrYliN4g6ELraH9YLWxHVJ
CaxPColrMP1vonUB+xKT+ny+DKnBZGem2bs7syoxF4qKiHFbbvmyseM1RJBvbPFu
rwDU9chsyhazKEjkth+hD4rBSXBm0zB9rDFcVlz7qu2VqVjCtqxGVrlk6cMIBnBu
ZLqyB3xfIWyNV/CPrLigc4630stq+GXR7oqDLG4agBbDurmb4tV5cgivJJX7P4iu
J3Ic0hbrQS/CE7gDL3hxKJZ4HO4CcQKxStEWXpWal3/p3Rlh2FgDwHRQ5pnjhUm8
Fa4WaZStLUa8qSxtiEkvHRBEikZtVqY3JCzIez6pTyID8ErM23Gc8ClGRKVqaRR9
7DPPFYvjztUrzPnVTHZuCCinICPYgxAb2kTrMMroZmMm6XIoQxyHN00hpLqL1vsz
5UWjqh1R8q9jXfob17REH0YimbDECTn6KGXYWpMELatrMSeDE/sQqFmCl7cp93T9
vRxT73vJGr3i8IC8EFU3txMZtabhpGxceF3kiD1Z85m0Qa90IrL+3HQ1j3YRHBwf
PnhbQoC+hxQrQoKqifLCEu3IDup4wgOM8/70A5/iaygmzgW2vXKM8cQ9ooQTBuvx
6b8dp46TikKxHEd3Rlz0D51kdZWBuyt8mTEKluWqU/Ztm49d1/9TSnXNUow6VcYE
Y9Kno3d+qHPlQ8rj1bS7VRFlm/NjPwcdqwG4oQ/8YE+AKAbKQk/FFthVZKvH+s1w
hcaoq/OkquvdPil8uKVuYDAR+q9uo9WuWhiGduXpap/gOujsbXLvdozhHKatpKQg
bHVSiozIkvwM+tlYVMo3vt/vd1nNCpp0QTwPFRGLtUC96jqfoVojWWIcXwFN+d3Y
EwkvWgL/MtaxWuICAZhth+3fLvulzWS2oYbrh7OVekj6U7isRQzwS8WOAYz9Sh1R
RwhcVaQuHWMi+y446ko7T2YMhrvPvPSk20ByXrAelJfRoqc4k25jch0EFZ9G8Aph
Gl9+BOX5xGJUf0VkCqk9hEVUzRuAwpj8KF8f4aCxOnifiHo3IxRYrzV5jvU5APDE
3DGuMI5ZhdLlQCMm1V3SnMWOrOfq4WiTnyEvxtiNsu+aSgyiDtVC/18iaFnRmi7a
rY+jEINbz+AgjfYur3LFJGS7sreNJkkmRoAwjhx3NCS9rfr8EGN/o4IOFrQJ7EHu
+62oWHMMHE9U4QMxtiAPWYKttWeny9O5+Z+cEGV7skKrD/keKXPtkFxgo3HMHz4x
XgmXv1aJTuace/SxTIDgMMldCUW+FI3U2YO2r114FRAU/vvKZz3nvgbUwltx9UEl
36F4GdYveuaBjkPd6cgq50Wh6tQTvk2QRwc8qNebB9LC3G7Xbf1ihJEEWzXV0MmB
cJB7ofQnBaPjdp89Ci9rGhTC5+C1gHr1vqnuCdnXO31AOLhf19016BEXiaxVSCkZ
vuO7kIuXZrPdHa/7nEqyYRSPtPnN/t5lYwrFG/sfav/Rz/UI0qvtsZDAvGjvfuYq
IYt4wenbKxlyiRiYaxcwsQQjD+IsbSs1rqlrQ+edIZCHXizzUSkHNhfU3rVKNhsL
5YkUNj/Wzv5vP6l6KbA+rXRp73TbBD33m//w3UetXWWCioui/ZWZXezajXgE43QZ
u51uXMt9LcDDHwD7zIpgBcYXaufRecDxLepQBvZ2lhIXzT0XinUsENS0/1YpceYE
FFnZwhY93tRCDVoHPT3ewcGqoUoyn8RlizuxHzuqKmWvLm0IiaCgAb+koLU9RlCe
n9ERdbFOHO3VnzlFtUjh34ORXW2m3rbMqmlL8BZ7SKKK375qcdRjT+TOl0z1Ld7x
e4qW8anDzA6ug669K/+6Pbbsi62UIRrwYrhOUDT5YIUz0fW74fMuqFPja1FytHq5
dCRMOLBI+tJIHa1zJ5OYTIkGPxUNbgajDCuq8/g7aQYiakM8OAKmhaYeegb7ucg8
EYjmdVonNqKQCHGOUSDUoJxsYXZA/JZqZWb8H5hy++IZjTpfXaB8DfsSYxNYmRpg
XZ1pes6r6+D5MbN0GjgLGZZO8U+6K0HNpC/OPhpXtCkKss9qsdKBhwEAavmkb5fb
musaojPKwuvSnVUb7mP0Y+heJrTkL1R6kXg21ecuZbh/xbr3FNhhRD2VcV4yzmR8
MUrpioy2J+fwTdh24IyXXliOk34ZJOOov9D3Jui61PAuEwbDfadQ49OM+tD3oX3H
VWKV6HpLvrfQJAvpGfVp08pLyDBfMJKtlZyKqWXNA+kARIrgVcIQfoRcT6wyGDix
uPvVaGtlqQPyo0jEKSXtRO/GdlE+nrHKk12G1jrh0xmstLkj9hcnOdoqrxc/0KQd
+IKFFa/Aj0RlJXKNww7yvyOyTI1WOwrWf3cw3TjcObEKFpxPXc62x0kmQmCL1FDb
6YUz2qOGpAvc2oPxQXoZARtvyH1KUUoiRhPgkXofN/ZqFLAxLaJKbFPPVei/oYEb
Gc+rnyruOJ/lA3i4OOessKpjHR+sylyiZ6efo81iiHJcksFuejAIskr6Hh72TFAX
/WPjxdBPlHBThBM9WCqArjswU8GteyRm2/YVGKjkhlSq2s8sbt1PvdKv5rOgtxGr
dpsGoBI6EwCu2ewO+1Rz1j+OQY9MAHLYkMYSm3D2tkqAIMY7LCa8TpXN5DfRf0hl
jASGCREb0KHkro7kyGbQwoK0YCTOg9yhYbVqZSdpElR83LWrXwU6VGXWdHAuTft/
ff4yXWDfSOqqIQTToY96AJAvpL/VO5JcRIPsYSGsNK7XsZfsLPi3Ko5UYyN0Vti2
3BD61/H9DO2AZ3gfDSx5YYry+K1JujJ78Fa9ZyGjhLLymPGd8KVZCZkueWiThuBu
IjsggA1MgrNFcIlD6ddbS7DTWYXAKp1ZBZug3W9Vv+fHno/ZRjYNlTJO5PV2J4F1
4PDXDY7gQc8/PQcVGLCFM9NTxqdPgsrtvqoioViNkX5zQJXb37CfBKNiWlr7J+Cy
N3tj1fJPB5/nrp1CrK7x2ai21dw+6KbNdC9Vg0UQijKyabCInYpOmtOP9FoaraB+
cAWa2Mu8IOxfRfH5EsxckrjOyOP2rmvQPm1Da4HgYLU4Wig1xNbDA/nAwBIaphAZ
JxILl5rNcfUq7pJ6NjK/0KGK9TGxUewT7jIXTPjjTf6q5vtf5IPvkJJDHFvZUKL9
p6MKEh1srsatcFwK9ut4ND5SlX/WTHF1xU172IBjzRu89G8ZmTTfLcAgb4X2I/J0
31pIbDaJTl+s15YHNTYLJJ2+YKGp3Y4SMUPwVR9rwDE98dfrsKAjCzPOABiJULMQ
6+XUo5MNEWdl2MUxvJ4ZX3W06Ii4JPxyio/DQZselTc8dNcSznIoXF36H6f6TD8i
Bo1ybJvzMUD0p0gOYjXebgKDx6tfKZatgXUOkokKyBNhy5myafL8iwNpagXB57kC
rjcS2ZSJ769Bp7uLiLC82EjxA/ao5hqiZB8GYy4lWWRrYRjHFNvuRZNDnd8d5hZe
uQk5xxepaRtO3WGOs0Ns/LQVbNh2AvR6/ZnHZTd4t/jV2aQHhifnFuawBxhdHnpn
Gs+4DxwQEA21AiMlb8hGuGXwoJVtm8Q7TdJsFQ3/uwF0dXKLOeieJY0ru9XrAZKB
U8DdsxjGrXqowfFLNmcJT2WbsQCXmla5ZeDeYeBMqtjtX+V66ikyW+q1clgCr/aT
e+cuw+jf3Lz51wTEZn5t2ACsoVFP1wsDxUgYR3eXphNQ2j8zODUgLHKKqKldLDsY
KKauXwYpsZv7VEUKfChVE1vOYjqLw0w8NCUDuN1d5J5sTEWBxbN40up9bFnukWys
s57yH7pue8wr9AhyIBe8SVNlFp2mV2PYof1+TAYYaexWn14bGEpy2s8df5tA7TEF
ElQOhiZ5fgovbW1bmlhTaMtlLtODFh39XB246R8EC97HsNAgN717pKsQ6oJVo+UM
2IhbwhkUZWrDUznHG/Q8DUEGnUxC1vwt7FWw/1CMqsIRLvOzJIWGUC9VgAfJyQek
JjFOfCA8Q4n1XqYr2tn7cbMdRza9k+8bjhhOjoEOEMzG/RWeZ0I/DilSqWKKNO6L
7eVFum5Yk8ZCfwLQVSGxyr00Nf4z8bbbCq9kPRj/aWfxIgsVNI3QRNdzqZjwThhK
gUTY0e+ZeUbjUlELDg5qLdEePWC9LumI3IuYA1704JCw/qB0OK6T6058sj77qRby
Tj0UW7UjreEVBQ+e8fqaPgyp2Q6OAtBU26bhOj1ElE6Dx/X453Mx/ilT5v542Ik2
onioMozy4qDY0+zfDRmLu+yJ85PkX62MAkXMu96iIB9mg4N74j7osu3zXF7iatLT
BUvq3JaHj9jDK/vAl71ZJ6Tf6y6b8S3x173s3efpAgRKmbpVO/SOfxIssrAcewZU
J85awlBP0GQrDH+kvu4aPi7u6UqnUzMLK2iAklhyBEYEIdUN1Ur5vB5punOkBKjd
VvtvpzKLMD4oyCGhiMOKe+lSV5udPK/6QHUaIsZW1oMb6I+ZQxCyy0RPYT/dtDlR
0nkNEFZE261b67T+bf9taaDbZi/X3buVH442XyY5KodPuu5DtsZ12Sj+0ILHKIKJ
BJ0gSe6OW8+/awBMEImmsN+XbKexBmos3y44JBt13vENRLqzbmn4ofFDmUyJ/yny
r++U7laN26IlmLTOerl2MpCgbq5DpwzuzhAGs94UbdADZD6sHNfLpSmITNGy5B8n
2wyDbxfl9RSsLavgvuJWgQuvbbwXhnRpFy4pW+LMZREFLSjSFlve7aQzdgfiSqGg
3Dmb3/vZ3jqg1342kK72+augTGfuE3Kq0Qk+tMoUFDuVSg6lpKm3KCsl4wFN8cxi
Vc7B44zy/rPGf6G+pRH/n9SpcTxflT2BP7Z6syGRpFrA5ofmnfL4kZp3tgb08lWa
Y69CUgkgVEOMSjjGvkC5IdYF0ItLIrAQeHTHxVCmufQs2xB38TDjlZl14WhifcWM
LiMJJC0aImoRn6hkvjVjJ3QdwXEfuK8BamiJKIBB8bxCcm/93AvjsU3R9rEyNu1d
m5v4HGp7ehPyEk/sbIluY6hMurK9EjT2arw9B6Ne4ELBwkh+v2mIiklNAnnwyAOv
KAErzhfcl8GlPTubkWAS51e1fDUpmrOvusK5J3LFHOLw0D9oObDZYVYKpW6y1xYW
cyko3xxTVXkSAabedaGTthdnK1OtJLhMKL4NeAoPCha9dykWv8sCQVS849NjIrCb
FYE5y75JqCAHzp1acrVH92PA6oVOYPE28t3jCy8sT2ouSLZAIL68IW44DgKt3Ig6
IgnV9Lu0RzrHbhSEPpz+G0bG1/mfBR+0/hNm/IJUqykXtM07q0RJQHboMF4CW/Ft
5jxNUdUryIz5FQYGTtLJtb33Nof1+Dg6/K5cGMxabHcPVGcFh75xwCCHnlaWhSmP
LGRj/F70/Qm3DmwpoOz9C30luFVOu97p1jc9z7zZhTB+qDCrOh7aP9OBYf55hAz+
gRV4pJlvjuIA096jwi8fJKQ/VULfszfxlH94FD1+hqxXIGId1B1fccKTZCRWlSQw
KWazVBC8ViPc2g8aEiR/bL6EKuBiD6f0AiZufOAPNEFq4QIRu3h8E7GxG7Gm5q7c
Lk4GHx7ESBmhFZJMloi3scG6vya7irwEhcldj7RhauB1THO+auKCO3S2KoCz99wH
f+y+fOx83rgMHx522XCnkVHSE8wZeQYeZJ9tgoHt6xaXOWSVCfo/l5LQzJX7d1eZ
Gl3nm+Wq/zodF76+9PC+LY2RCLR27vwtlniEaXOUv7EPqMhpD+7GCIfZb9ZE8oNP
ArfZ1F7HeiMAnsaEsuu7qpPqmXfyoNWVk8ZdfTVz2gFZrNgaQWw7pDZmbkGso3B8
Chtl8nURbawoT9EgvxBVybvLBsLdJJg12MXCl1FAsOx9aCVyt/bD/B7ziRNaTH8Z
djC2hwtvZi0nQbWgHcQbx3fciB1G2Sa1JZibiaT1PjGCuYFeVxyDK+D3YLGuTBAX
wCAs+3UQHuDdrt0C6OSEpW/AETjRgsECMRQZqVwhldD5h7kKp3XMasrL3BjbghQP
NE1qoeLKwK/Di9J4FuvhtwPJ7elPHr8kKnP1tScT9Kbb1ibp9EUQZXnO9QoKyMKb
c+9Z7wr1MblLnaMSbK/VJ+d3ugs9guZ4vYLeb0mtkNgQF4pDAV16KzJcVa/FltvG
41rcaAmmSf4UpGXL+xSWw2bf80eCGq4Q2hvBTHRkUSvaeIk3aNJGy2KxIFk+AZLy
+1TymFGiZWDom3VGXmmoGtlN0zQoFMgq8iAEcxBVeSvvX4WfwC+tjYbLgFo8Zhyv
GQ/vpLngq/VPmon+1TxRHU48DyG3l5LqTr2Mzbmy96sWEG4oakSfQpQJMC86AZMN
SHxNYanJJjYYLm9m7SmezcTTxtnYysrcBrono+vt9pEXFx6ZOKIYohVst0s0uUYl
mq37IA6fkw9Oo0U9B9gqR2pxHOO2/W+RGFUXTP89IjfmOKLVJfydZ3+8boFAK32M
5KFTuZcWYW+QqQsQMUSnNuxMHoXIMLA8ny0YbLHjZm97MEEwZNN9qzR6xfJ12YsS
vPNnUJlKs+oDZpb2YQs7LOwOQddW0VocSqx5ULx3dLqz8LNc4fwDrjNUyQD4UpXv
k5ZFg5H6U00tYyLgIxyB+P2Cni/LO1YJniaqlviL/YGu+9SDUP6Kmqv5YEINWKDj
5v0TFL9Vf88ZdfdiOpin8N29XSJfph+KSb3++YJIKo1gPsCxSF3Ihm82jBF5Llsd
BfNRrZwnFplEMxGX/g7jaP9CvrQXVxHjdknjx1tlsOcUpYA/aAkDNu4SLbSQeDxS
mDSap45Z0+zajpkRC36W2RSXzmtVwCcAjYHBzMZ6r5cWGyfusg5lal9Fcqjyxl3U
g+dq77V0z7Y7dwnyPN0ItZnjh1qnQzJzpGooZ6nnvTtE7CmqjrOufdp5b9ccagw0
n5weT91wqw8yvsen5ijVYOw7RKVeSK2rGqtHgeGeVWDmCoAmRCcCZGNnHKwrQVuF
+IWS8FMptys3fsxv0Ent8TWY5ncoUGzwj3zBhxGag0WTPvoYkqTLRnx8r7kLbfev
zahoziuKjSxF6yXsPU6xHPUUn9IAqKEqmbYujkTYHpTjZOi8uHwFwBA6wBl+benh
EpaBWtbQOCb79LonmQyZW4ZgMpvD+yhwzA45fw1nv64DZ1fwef5QbVafluGPunzb
eTQ1qlQj1mFoYxUxYhhu3fGkS78Ck6I9xZg/YzTGJSlz+HLJXtWqd5vXmdEAcVSe
oQHJzUjIpRy66V3bkOdgB51PoBZ8lC4uMUQm+tCT2LspHvPvO8kTN8xampnAQ/hW
zqU2cOyKB9twZT1KNqUVIf5DsyaYvaqE0HNmr7BMoYtUZ1A6f98t6RMHThWG0Dzf
CgWW8zUrIykMGK3/xIerJxmWIy8Woar8RGhe9PNM7Wehew30aH/fdz7fh8F90DGN
a6CrxpVoA8yEHpXUvjFXlz7+kzeSPjdmGMHHzXRJSlrI4EOAm5ZGx2/BlqNqaT5y
iinENTF3c3XdRGY+K7MoPrIlbU++x8rv6Y/60hdSLFRVvmi2t54VeT8x0dOOat5P
EqoD7y6aYj6sqVWgFiS5aqvbfujIB6Z0l+/wvXsYJylxB0w4P/Vawj5aqRb4mzLy
61VvmR8Bz0nCHNMBBMmgyW5HKfzGJKT1cGDu24w/qwJwzEHZ4BWBj7MYrIoNU8Hp
t+JpP4kjbja+u6+heQsykHLo+SkNyjwNmGyoEpZ3XiXxqzkl52X5Y2RDMdShNHnJ
oKNacAaSGr6ENu5MUsB0EWjrYRvn3YIdSEYEWSxjXedtp83MkZUnnVagoVmf0r32
xPsscsOf3I+x9A3/O6ap1+z0TAVTX6nlf9T0jqLo+UeCURVWZ6KBF7BhXFlEc5i3
oLJKzhLaZ0FMkX7RRTyQyGAuarp/tL7ZdB6SnI4M4nshMJs4svqHCqtua93FQQTT
8frQOPaOcdVOzBIwOiBpjKyTUTNS2IV5IBy/fvFg2/5Ay8ZlXP8YSX75cPRLQa6+
/DOSMc3X/WtdAVfl/SYwmNm0fo0epY/NQeJad/k73EFRIC1kkwFaRl8DEPsVUFB6
Fuyzu2MKFw3dr7UHKp4o3yI264u7pGPrOlfSNZu6AktvamLp8LTf+435UbZve9Iz
9c9fCvqa30FR0nK2vsftR8vF4qZm8JdG9TtPXZbRdx5tqx63bDjpkTz5XG1I74yy
wV2Zpkp9ktvcoCuNQZyottsl+YSdel/l4Ddohnx5wfFQnF6OUWXiBlRjRAhAooXi
i8vwTqXxxDO6wVthZiQQN6L8TKttT+tP0iSKw9LOKpPgxNex/eQIVqvqr306pBMh
SKA41fCJWjOxC6BYabpV7n5gI0GCivp+u87M8yCM7+NSMhWqCB5DOMVvFV8mRsm9
YRzgSxbniEJziqjpxmnMKeHZhqDFOipURd8wNioDfH+b9sWeQZiD+wcpiRRdt963
FhLEL2N3bLCE+U20lsAz4nioRslFMn9uFlQ/HShoAV5Qb7PvZklKTWeydbawZtfs
v47sB8deCn86+MT3vz1pr/XsYpKMI5MlHV7Nb5Zk6pNruG+Bd3GNKkRH4Su75fwB
hz+deCMfK4V724DAaqNt9Y4Jtu3jSpblLeqePYQgq8qiI35gtATtsmETalTnBaX7
HLj6noSfhAGYMh0egb4MWbr7liRLGtNgFeCzOFcZa8nI9M4h2zMsFAYkZKzdpn2V
Y+yC/EybcU5EBB/cEJbx9l9FoI2Y3MsncAMcGET0p7GLILEJvgwSGV6stQ2fzs0S
y84CalKK0kB0BISAVNh3ry2VmzjTeWD9pXHUn4OCU+TPUMpy7SFWIt9d3aQ6rEKy
sHRapxsHHXe/+3TwRLtOeIKlt2o2w8wRm0uVBJRuE/eGTKI+70BBUWj6gmKLANc3
PgNBbljLZl8JGWVlqYgmQiP2xFEkYg5i8ORhq4Xu0lGNyC09RUnv5rDniQP/vq6E
pcxbYQoZyjZBu1OSCQnctMoD+JjMBT+Z+isBWCueACva+eariS4MqlMTzn6CWFZW
q09v5xPTrCoa0RyqL/vuVoUIZPYOctiDVeISk+rvWoqvnkrZ5nwnnxszW/xm8dRR
kFxQuJDoBZl4nqMIneX0i+zlpzApCckosyKbcdoByEnB03hOCpqqgT2KceqqCLxp
/gxJtGjQc5XTIISCQjCgnLrsbAxGIfiAb2eIdO8JMVKtFEj8RUPjZelZIDsicXkv
gaSUrNYM921pwye8U3O5YM7lGvi6PY/50BAs//vEVO8yqUg6SaEFANdnufKM9OHh
oX8VKuanseUR13jMirrZbQ5zKS5si5FjWIQVrzZQfKRWQalcP92L8FeUeFnOrQCU
6A2cihbJ74NG0WnRWBxB7isvxFJ6CZvHFcXVS6llXhPjlOXN/4CfQ62dpv8PsQUY
DIZIn6SyrQ0n2/pgW322vb+wLaQ2mgiqP3OBeOVLju+cuzDALAjchQF/MzAG7tYh
Er/UWM/txeARFGtTQk84F6IH7keMtbs+tcUmLT6kdhESXXjrglbOGZNThfrm9BiR
aMbT3KFRpySpR1annMFlAzY57h7+Lv5qYqjirS0qaDhGqxFfZgjgFkuFZhcEKDyK
tHizPE403g8krDg1/mEA8tXCP96HomOI+9K6ApJurD6f5Ui31LHZPQdGWOHWeuI/
BD5FZoKu+plmG70OhxFp5BoSL9pcT4LeeFdpFFLJ2CoJHhFHJCZSqCEF4lZKjfkn
boV69OYc6D2Oh4GRgym13Ez5m8MWCpgaSBatfG2qYln7NIbrGZqrt+ERRFz7a0k2
H+wCne/8IvhaojvkH2FoRbhb29IhNcZ7jDabClSKGLzAPN3Q0DaHVGypZJWJUAsI
NJ1RWU39Rza9pWRxqSzTVUAxsZe5+Ha3c/Z1GO46MINjhHiJAeBPkVQqm3VtlEPF
YrnIWrsf5wuqKlwwH+3xQpWbYODX23gUYfoRH3hmggDnzNMoeuLNBT5IF/xKl0Ki
gDCwYLZv/QHo+Tbqg7o6nbB3qTHmE4bSCiw6UCzCWYDjHUSmYwzLQrxuoWfXLM9k
xrXW6J1IduLMlEBUek6q37rAt8z/SytUQXhxVSqFCDcdFDiO4QVGBG/4ufpewiad
7BUdXD6saUL3oTX/W+jVpK0x6kT2/vt8yeQ3D5Pcfv1fuQ84qZTPeWGHWPEkp+54
4Y8CP2pw7GrvX9GCnrOgEJnUCV36IWgp0VtGebMeRZ0xtFP/TY1DHztylpN8TlF2
LxruA3QzZGWP8ebMQgJEikiCyNuaRnKBFMcaLkziKwCU5PTg3iUQGwQcEqTTi60U
R6pucaua9xVB8mLy6W0NSVv4X5PeasZ9yEqzI1NBuFl6b9D80FtRrJ1mfxPvbiYD
kxzuwCV9mq+hKWKuPD1FhN4A4apgopxsdtyM4gzOe56EtdyorwmJT7sOZrn7Rtku
kmnpWRFZP9KvtuFh+Xu/3pqw7xT+OGfFD8URe6k4BNuHzb0FgBwy0jt9BRpht+TZ
nNQP9DCuOSpRBnruRvbPS3yHc7ISvNHrqmvqr5sZHhOIMsAZais4WyxdGMS7vQFH
ob+XL0h6SOQTzSkz4y59gTLTL6H/D6IP20179W/Nb896QZ+sA9XOcH7WDEdrnC+u
JVdV+8CsS7aQb1bZH/qADwqrUVLckq9tPfNXcuQC0wFLEnZPjhrzW6tjcp2+elFT
VxmczWs8MlPrjVtdgbEo9BYu4k3lg8VYMOrBPPpHK94tw52p7ffsp0RQjsyOMkZ7
2E//YwcgdOmk1+JdxTm0Y2pafdEGGhIwMCq5ix+EcW2BAQLCaID3+yV3jxDO9RwT
OqmDdNpI2XvaZEPDCJMmNFWd6nBaKLON+Dn/lrSlyDbBjp1K+CgZ5EM9708W1pU2
SY6TcFglQKLTuWRMs7q71MvwlyFoZnKPOKra0cqY4GmBuBeil4u30eJGQZRe69Hh
6uUTsxXoIlMjiBn2SvIlacCY0YQk7kMQ3oeGoe0qF+b8lg5qo1rn2ekTqmAxxfHO
S2MAw1mpo7795i0QG5l3Z6GmZOyATIdNlL7Q68qJ8PUHh1pRjuxJi0DccI7vqTXZ
WJUXn37nbGNVaoEF0/oQUc2CVx9CZkZboLqxlWydvDsFowYUS+vtrKhvDSSPXZ07
/jBElHqUofE4F5jkXGhMTynQNrsQDFx0pwTH3LFZq/x58EQq6X7ssqV3rV3JeUys
osuftzd38fV1uGDF8ybyl1M7vkhw/B+gZNpLP148wvBRt/AJbOFJN1AbJVl4Lv0s
lsMlsVYC99efCTavv6dy2Ht4HVj+PJnuLv+VGg4XYhcdPwMXgBvRBlISqc5pTjkb
UpAnxUPQiDUm/abkjIepgAbODwXf9DQg4JfwRjEWuhV8Jg3IZ+WWpIMiZGh5DSko
vfxcTvVd66RiWTlnfnYAhlGZG9+k4eo5FBd61bj7dbsfBLRQyA3tIDAVFwuThR4E
LZJhcWBMdgF0dkLu4qxeGn7YECtHlI3ESrhPf7ddB4VfTGAVwTbQvxMzwY1JSSFp
V8ca3ZAYrFRMtB/nmP5UVOtWc3GEUaCjPWYwP2G6rlDgpcZHdXtHlflpU4U/uaIc
kAEG+QeN4t2TQvYEu84WiBzEyXb9an+wwf3fH3Bgm6cO3eHfzJtPn0HcOrOcNw/n
1LhShTfsqGVTIumu9rNgHELY1jOt635F3YHhtTLDuEdH7XMyK4Pi6YJ08DiJn8KC
Ex2Vm+bPUBVFxnKDIUQsNlSSB7wB0VDFnbrRrJOpYz8e2iVyxJ654Q7wJM6FS0Tv
ey//36ZqityWfzWYr9I7oGBumeHao9l0r6GWJcipz7aOCoeHKlt3j+SDAAEkhm+6
D5zmQDnk7/NlUtX7DzqWP/dmLxIC/bYhStHVcMpnecfc6cz5L1HYIL2ZdHj0XhsV
0ItqJm/6B3g3ycvXEckuvaesd8p63020HVLT5hzeI2iloJV8HyIS6GxzzCkINZAr
Vn5jM3xStBVvp69y3tgd6xRPp32By44MCGJH0ZuJRDWDtE9d3XtwOyHfEASVTfvv
1ro/Q6GCBwnJpxP3fs4e/WmReWXd5JvPLy/4NtuKNhtQDbSho+W7SeXAjlbyjQL7
1AEpQOg4Gt0aFSTMJLkjLRJtwGLzeqo40qwjxMkHHKiC1UxfzROpfmM9e9UJD5OE
CBUlDl4pSJLLb/L4KO5UVkAdd6lumLtSBEbITS44WhWwu+iaQ7jYwqN8e3L+Fca9
/0f5l+Z35dfPteIFbEVLsmKFcSVOhpi6Lmg6q6I366YyLX9rTCF9dY7C2FLkD/xi
6VwYd4rq/GRp0y19Vy8qress0AL9Gt4vTaRoZZFu3aR3JNpG8Wqp5W6IGTB6zIsC
bj661lzokP4NLoG+xAyrXSIAVeTsswe/L/G4UvSaBIT3YWZu8C3DfTNla0eJ9Znv
xzNwr3ozuCL5BgSj7GbOPFcBSg+TQMC1Q/HVEmk5ngdmZW/92uLShdakm+w/eCxf
EGKdcoBT9xab2yjssL+xROlOgbACmqlBIaehP7v8qsLV9zglgS7C3YJDchfGc9Ja
YpOFlvUrKyweFiwc0XmH8aGd6lRPmfozkuYSzdfq8GAfIOYVzt+IDvOK5lcxBout
WrBZY57k8XOsUtIFLWrRiy73n9/2zIusSIItyLaulSU7hbHgd98KMau4S8Vonu4T
6UeXyJH44xkNBLLrff2kCrcWRf6pEMje/7zODOLmVijoaWv2EaNKKwEjheUGMW8o
T37rGoXUUnpjc5vxeRIo2f1K0UNO5kQJXmDyv9vtW9WhVR7FCmiyLZ6rvMMpohEP
ncjj331CqbIrq0UxgajZoxS7HYfbMUmYmyns2gwVDhH+8zlU1/Hg2zgnAWadYTyt
HXfjV6T73in4+cFNDw2obTx8I7/9GWf5iP4S0JFmrlcnMNoEEfyhNwJMysVe7gq5
oT31vWLb95Tdl1gfIIU4BoX+XgfRZg7f4VpOTVo1gVMRTlu1qmJh1cAltuHfiLAz
+Ugbt7RLOBp8KhJCvf5KtftvLWY9UIHeqj/n/36Irym7mAJCVgU0SBZ9XsMrAASp
EDN2PyXK9g/ypVRPeQSiXwA/RI0+asmeHgfkruIJpqofSGmADKE7jvOZZ6Wg5+oe
tRKyVZrvVAX3BpBLwt/f/3UbkXTsECPpHMXrT21U3GnQLul3mpwWWjKDeERL9O58
p+hXDlbi0k0MxV+qToIhTkiWpWD72hoJcyp3KJUZty4JAHhOQB2SKKcynsilWkoU
ctwDBkf7Tpk/44roMim+Ouwk49RpCBav2PRxkw6Lgolyq6DIOIwfUnbseHvRrsnc
6KsDdY8GBDoP08jt6A/PdCWpYCsc4itzuDCMmyzE4mLYR8R/1zcQl+pUvA7zQy2h
BRF9iL+7JBQXSUjzwxcQARM6Ll9b7sgzKGn/r0H/plhmWbcffdJphHFmMD4UR+XI
v6dFPD8Yn2Iv/GB2FCyrLTXRCN9qL9vlPPXTe77m+673WrpcABNaTxK+aediTId/
sNVMDp7+3HYsNpoXwGXGO13Q36TDMgpsI8w31SLYG39VSmWT0VNkJZkvOMIteY74
Z8et8GOounITFOdADJVvjNixdVVGZE7O58ukSfI82uD1L6zlD7i47KJMkfSnQW6q
R+VmS9OAFJRSX54qywWLOsXuwFJ4ci81aM6LCmZBMMC3Y+O/HfinIWqXYJCnb6B/
dd5g3aA+vi/aeiedYukFnTw/SUmdonMOElpJ4KXzxtu+vzSaxT+bCfs5VDJAN5Ps
OK+vBNmyEoD5zfJYw3WfIJ4ubkBwI8Dl3CBcYfA281sw4gZy4UsgqfrwAkeoEvIO
URXOcFByyjUZC9OspQmQpx5VL63ZgdPDL9UzvwwMiaSAYCfx35viqIyz6n2Mp4T3
bIfydR4WbF2avI65be/FMwcZCzsFMtmS7mHxT7+8sEQOy0CLbFz5XtRMm1Qh2Sbx
fXCpVtmnmlo89hHRt6zlhHOvnaoN/AWkd1aD3DlNQgekrZjHe3n0fQKIkOsoAmbl
BkhDYYmntVqzy/r/8Ng8FI59+DAlpDnsppauOFR22/I+40Qlz9bKUk6TPYbBKjdn
Cl9nE068cYh44LmmE3HA6H4LzHcV8EynUzvrCVWwYnZrwb89cbuOMx3NZH2bKLRA
UGcV2pssoA6zRCGev5I6X4GD3c3Uh14VchT9k7Q9OkagQ4PLLDQb7CvGwau8nTHN
ZveTS2YWt+PJl41sxdebvtibIg4/BuuaolmVWp6slxySHk7ES+9O1NGwANIxIBVb
yIdFmA3sC2/z40GIuTefBlTvB7J+4O8qaCy56Pz/bVZxjfPeN4wpW8p5Ar1ZHVMU
ulnwlAybldCHCVva+z+GcvECwS8maNn7PhV5ryE8zYM8HUV6csYQtMMLzy678SNT
IIsfo/TOVBchSkaoAM/IRiiM2YcK2CuACXvkhWl8CiaU0YeNN+jye3YUZyVni77P
r2T7CnSTz9YBn5J1ygfrnmEyhC8FvmgY5km0UUnVSxa6lSLCZevLwaaYO0pI0Uo2
jIFylFaF4b4UjKzCCd+nQs4S+r6ROnkrhGcBbbhnmhSq9xx403Z0dr1Z0wfHotCY
CsLCI1k3sGOqzyt8FfhlTpeIj9GTDY4jbqAOxq8oY/QpVZ/w6r34dSKhACyPVQtJ
hULq4xIiQDWHBhiplU06Ghv0/zdmQ4xikMjT/k94S9FHWs8qlgLb6xvnK/5kQPjI
5Me7NQpZOBwxQSQZH8j8yfi7csyVPonWb6O7wTDpoJt+YxBjfCgKquj9IvmJJc4U
s88D0HdgPKppsdEtVPBJ13lQSdpZUQ4m8eHRk6Vd/ut3+khmwhI6QUSAkYmsx+Id
MI9W6h1sn56FLnUD+1Ck3nIPRgtK30C4cmoCxbQnnu+HbZxFyW28FvlGjVmGhMY8
Vbk90k/FnT5HWYdujuRCXFHf/jAHEzWdydlyu9YC1d9cPpZWGMAi6nNZS5DPrro0
oGlMuX8VW57JBuxVg3aGII593Lk0F1o2cbzvXVzVT7P6tiSezuJghO+8ecPS6xku
4vETBLaGg3vuC2w8pqT9D62iVr7SkkcLIwt7CV8s+Tv94UHkP3RVI+Nc/T4Izhej
VmCx/uHafNbezQvj450hbHEqxEfLjNNYOv27C28j/mDNUIFYTonCwb1nPweoxD01
e63gwtJP1tj1lGq/7I4H3S3W5iHkCow5ZE23rbrz15xm3dnW7o0D1hH/UovY4Vf0
lzbX6pkqagSLMAE9Hu5aJeeY+cUcBhaPjmFA+gxrCvsYqd8M0Ig+Dfvbxj92bskS
2KgLnAEg4HJG/WT9W5AA+hfvq3uz6Ut1pZjPP7ZHXi7gHnRNZJPqSFy+0/1w2JJc
Vp7WXeIbB7co5t+wEmT73O2Xy2pybEl1estyYPhntMhszaVcF4TWZuUDujzTOoYG
zGeduUwbvK0QtP74/dCKykbFhbRL8sqt+rwjO+51jYtSbuloZs6oZ/VytEJsWAu1
FIWfTQDiLBWvRCKX1DIycpOLf8iCxklwifs/aQ4Qj0wfL7cYiptpNxox14nC11uw
syd82kd4JwlHjspC6QKpFo69LZLC4xXN1slP+QIXRFOZB3ekzrFQxXkZGp9efZ30
66Y1qe19LQk0AXltaz7kGGQx7a6mlK8kzoQRNEcXa1HffsD8lDURxD3Un2PD1ar0
d2UDTyjKSv1Fsjq/87YqZ2EL96cmDcDzO6MnqSOq+NRGyuNtJ65r6wUPZs8Q0KSq
1IvDp+V2+9a7JGNIW//mJIjlcPuqYg7vHoNeDkETnwZl5+5xOL/MHMMHg3WNMf0d
ce+Cib0gHhWJxmupFX7OCsu/5H9psw59BAYcOqGl45JiF9nOa79IKMCzwTPLASvl
vjf1/dzbQoo/7z7cCdFDEentiygeV12RqYg5MV9mIYQ6yw4xKVXRtz+qvrWMduu9
RNfVFm8q8mM/8H7/aBRwdWurQuTfRKYdfZ8qgVjY+yvSGtC2Ery5cl1DBCywYZB4
mXxVbjOJKNVc9S/AtQkryAcb40FXq2ESERq7yN0kef3S+z4e+kbUVGDm0lu0fyE8
h7vbrpnDB88ypdt+ll9VaSyNnLocm1bPvE2xVjWEKwIO4Mb1MyNtgwUMHjttk4At
R2zGekqm6KCaJ5p+PRZBianlyIViBMwy1p09/K0S3+3aCA7UBKjdcPxqNrmvu8ER
PdvQVZBCh4kXjXW7RJc1lwRgGVqvSJYnWwpG2HwlWBieudzjnqr23Lf6Vxix5JO9
mjjWQ0suRFZQVY+XgtugGivr7+HULTbScTYd9uP9+A7k3IvS1B7MrZV+2UaVTJ5F
e0u/c+gV84AvuPccJxqigVd4EApPbczr5G9LGUAzWOWHG1N7UUdLTYu4NUibwoZv
ieydW0AjxAzxtQirdOG7NjyELdBn7OgBziX5T2qSvyIk53NKkfndBpK/Ny1cON23
AgRQa8hT70B6BY/4w/ToQF+izHnU/jO+O056kRcSppGQvzspOWKsQRkG/eVtNKqb
00ozxZSO7FEua/XxmBbqYxw63P428CQa7uPuNXHGMjRtipln3nJmm+8mLHsQEB+4
z6OdLlQwTYK0Uf2fjbdIl1VhRudCT4Nh1F5r4KEt+Vf3ywDOzBB8zZrIEhwGgInF
01a4n1tFNWmgUM8JOrcmI2jhSsNOvwNnbOz1r3wnA11oVPNYVh9Azqk2O5LGl6B4
Lzg2/V1KLS+dgktN4ZfJdY/DxSWlHyzBL620tXk72T+NIKXX6LH2w5lZJA6ek4Cn
R1tLX7RTifVU0pHczyQ0Al+s/d+mj26IwnFNZhfoiRpkj+xfhSXmONPCApHQxKpw
CEfXwQtoMitYo+WbvZHqS6jclRHMV6+VyvBHtLOGX4gR7Z4g2hkjnfbgLnGyCO3u
X8mvWcoIbxd7KSS4NTqkfdKh646ZpKK/4gtBKvyIA7TOzgcLRS6/4oCcOxMcj7v2
/B+Gq5OVR3l6H5AkLaOidx1nT9mwgnARA8P5u0eLOb9V+Ato5wjwBlLbaS8Rw9Cj
RScUoHOFr69iT3pTGQC5xKo4J1VQXKOm2+HmRt/XNvs0g5cjPqGPgIfQWdyc+gyk
8PJs8fQSI8/Y91aRjYt1n6lZMrbwEF6MGMJh21Fr0wiqFwHs2hQN6m7o0ls669GD
4bIJUwcxaiQmx1RGZuaBAGCsmCCaOQiUBf1W+EdyOXXTbWRoZCUpgRVeP10cXY0R
jhBwJE4o4T8XErfb3fDdhAGcAyzNSRuDHxq0jRVCfSje+0b2wHcSsQR5w9Ug9kXN
/TDkzh7WKQ1ZLvYh0EEWEtulCXGsGkRXiH6wIb2PgU3ydbgCpFhlpCfYNLy68wem
nRC78GC11vX1TvzlC8eLJKDN4oFOtPYEqVr3JwcBK++fAbhmRGCh9UqI8xIbk824
HQBvxXRRtVYyS3DV6KKXZKAIuBnMk62kPYJBTK+DGOP3y/hTLmCC22QVqJEcJAcI
RA57t48RUlxvhlta2kotveqV0t69w9RfdUBm3KYLpRBWEtqYEhb0fah1YErtuzyA
v/6V4D+lAECvdlaG+VYNseVsPC3tvmZBsAemZ6RZbx5MG3q/1AQSNEsVSHRzR1+F
8fakp0+ukpWfE6h3sIDGuDv3gTRk2nDYVxzvYTYFtyWsxkU5Mx4US427Nj2SRXTe
QNlTrNFPLSy3e294ZDrs2fh0Ge56I2PD5nR8kH0cyaFKooHesWrC7YN6imz76czV
zJfCav5syIalTdDyYmj3e6BYY2MZhsOB6KeqCRgePs0b0/BtydFQi2t4c9Lp8dF6
7xMNsr4uLRP3kn9K6ElgDZUTiLPI8E1fL8QYY4NX5+EGiYe+ebm1N93HSEaVTrgH
2lxJKx70AGuSS+/wNCNlppQrrdOItwzMiegi3EdswkTT5LxFzFNFM49CTe3u5Nio
KhWYr9oSZ9kcSKt/DxbOBFfJF7tNIYmImSRfbFE1wr/0aazCZeeThgctMmckOLNc
QoFbyJTG3Kg35kHt8X7dUnZ7Qkcae/usTtGKs9AqyCQ4mGnE94tFQN3quRsXTMfv
UcoNuDhvw4pOzzccS7g4UIdlJbNXR+3tkggbG5Juoh1qG7ofOb1OrChC3fTlhZmX
i2kducz5lMGvh+eSyj0nzsey2soFvWNWY2duuVad4+fUQttItN/rIaN7jvUVlPid
eejpaCWnMnhwsXjQmJUENkVxeJjikjDpDCjz3Q7UYTMKxGgqq7TL3G9VO2C2Aoi/
HlxUopGKSRzr0F3VHkzUMNzk66W2uMY0HMzojicfS8alJRbrRJ7LTyF8jaJHXuFv
/VkaNYhnCMZvloeISFyqKvcilJytDTS7g/o5QJLuGngvsVDCVRV+jXu2VM9eKToZ
8oXqWm8nEa3go4qNBGFbW/HxIY297UIn1+NO92jOnAKX1c1VE4Fv4uunTF1iTOc9
h3n3BkKnbMggCDtyHHQvDBsY5JSg6tQA1DqH5XjnQ12Fp/KfhnYmfpBFmH/VYaGt
1ekq6F4uDUxPoL/Hpo87bO/k22QKFxKSbQnJS4HO2SVys+tdvzT5TwuL4hwxaR37
pWFDSArpCEPOvVnbU1ZoPZRF/SEn+FzzLkgiG7cyY8r1/5Kx080RcVv2Jn0SnFmV
QN7fjg4rzfAGTwKF3tUrZ9FEMWl2GiO7SS6Ns433ClEaWs1UXbIyKQ8c3VDq0sJL
pr8IzGObFUtgbza4qtD6QqBv+80ecFpGGj/146JmZyC+zlGwpkHl+ixT5SB+LfKW
HrpOfRwokD6KmC0jib0gW2YolqeiBZ/SFNDZ/2MFbY8aHx4VJIUrLtuFWU/vp1Jg
6628W7W/i6CsEu7ipIgoTXAQR9BhZMu5IitnhQwqs29Y4/eFr4gvAlrE/WFVcS0F
bRUjHdPtiHfDdOom2s4SdupztXojQD15WoRKFw1TbArff3OTOO1UdPoBTw9YAmwh
UpN+37uaS7iAIfNKjYYmCZlJn9QisPzkMk9L651kPrEgl6Ewin3p2KzGFcM9dOFG
58+XxL24eNdJ9wu+QMpozTA8S1sT/KPqsSMpv++ybfnI6KlmQ2Ry5PWbGdxocqe4
UCmhcsdOBfIBqiKuXvV2V5+V/GMFC7Xf62Mn42iPoEXBZ4eot2M4tBjCk4eLrZar
C7rHoruXe1qHu2W9Plje/et2dbvAkTomRyHhpFwaSz4+obHLdH0VMwYuf+Elh14L
dGUQ2ovXV3c9r6y4VORTbb19xFkSEmm1sY1b4wtksWHBGVXa5SuPnSSGRUV2oQF4
ET4pzc83vpxXnkn9pZYBE648rsnXecxAa30k8nZGGyQ+Nx1OeSWDFn4Fa+fC99vq
fYVCPYy+7gbQ0jE8J+mdth17tNAPEuXLaHN/+C0QxbomfuySB7c3+NZOKJeuZJRR
6JfIVRcqocUu5txxiZFPBF4VNQbu3gS7Q0+5HWV7DBSOCJBiDkgmgSD/9/PeHNAx
GVX9nXKuaargy5YxA9S46giNRfKXwjcDNH083F3wkBbiV0Vqr2TzBlNLkx5nF2Tv
bZCUKgFDSNPDB981oIq1gwg+eh9zqj0lI8mb5molPWKd1zl1T6Nf8wXJlby08fDE
FGPG+NCD8oXAaLIvy8srjPl7Tl6eNGBFUfD6YlxmSk08W7ALieDjc0EnU88OlnwW
+o7kKm4AW0DpFIdrzXJXkVZ8phg7AQBEOnITXYNdfxEXQmucRdUwW0eqEJoLdJfm
mOekZPRBQJdNhyLTJTzZFyj0H664aBtNjD5qQ+Ws6mWijSQnFZH2ONSmlpE6wGGv
qm3FkZOGD1gKYm85zPVbHna8V1ew1qOTm9iFaZxPplQWlDm8nPKlGSmkGa8CluO8
RPjC6CWl2pv9hz17GhPnXnR5c/rTWsxxLUrgS3FAFJe9b0nt0L/3iNgkZF8DwU35
YZ5cqZN7ZS8QKwBYeUQKGMhJZ6WAnG/iXz1RTBW6GBkzYoNbMF6gilOaTWCHoeQz
K+rzloTo7uzlynd+ZPa29DcHA1jCNt4dnC4n3dFgtpU2iF9bFIK4dXM5DJuiVC8n
MyShfJ5KxM6OvA0YAjOUXM3x4pdQy7wIBPLTwPz187Vr5b3+zWVxib+B2lD+pGPh
H+vZbMLcQM8UP1WFGv/IZcgW/WjOnnU7QsQlZm+/XXXaNjWXdgsaaqgTSJppcuFc
+ivHJm6KIEtUtWTqtZoEH97IO5kIXeGOhXa1TUXsMCuOcyTaHIm1degxvLLHomRd
kMmwwl2qfQktIrkIyF+I5scQt1P/qSp4k+MN48I64i0D4HW76IMBFWfGmxzWfugc
df8AxsVLSUnEPVQa7uSeUrtx1In1PQcEZhe3db3GYRBvWXb9JpexnyVr74mUffF5
GywL89/hrGXTW7KX28t7H7vBOkl3dH4aaKPBX6Xoq/xePoUH6wJCZp7FkNOerhck
ve2ZIT6ZEwd/ATOsvrw++Sl4uSCLzITZbkYZ4Puh//+QI3ArL9uLUE8gh12cngUb
K7ugkTyQELmJ3FCu4jh4T5m0hDRbFwy67+y6LAnzg/fF39fIUVg748IxJea+1jgj
zRqCigwo+Skkh9C5HypvhnbB+oiBLNinNpOoUlbk/IXcyIscCGWSSMPCPLfqGA/w
524SrOTw3fmGP3mL44wxSJeTb/Y9KEe01hV2MaHdf+O7i0oKxA5IyrgOqFIf8ASc
MU1ifXaMxn4oyoCmZee4XkE/mtN74vM5/X1wWchf3F2uPsa9NuFlw8c57RCvjIlR
33vpcTJSW8BRakMCylWZABJdfUSpLUr7K6JUcArFQHJAt18rk4OR0ynWRBAnARG9
F3sP0dENG1XQU13JUZL/QfjiSlBBPCa6iVVhWEsYdYELZSFfleQiYWhlzyCV3I76
rOJA78yeaxkh6DYpqxKuQrC70RCRt3bEeN4jlMTDxb9U8Btm4sVmjKZVqESVgtog
bivdouBk34BSTYzRw3KWAuW2eRONAnNtOUpwRRj+ZrNQIjrcQ3mIcqQIeSyN6fqN
3uKHCxUkBnGd5IDJSB3SNEjmuPeZLSVg0pkM7dlvhHCSkra7BOkgK69RY9b65p2u
sIwBtAKMM2iVbOFYvfp24GzkmNhIlDXR9mtQ2u1f3i60tNKsGz1OVlCAgtkvPwp7
armiyVI9wTdHbUYl7SJshCRF7EKZhM1G9t/TFEe8HDCLG7k8P4b30IpS2YVdAR25
hsGQZAQxn7Ml532TU+pUxzaZejNhlneavD5jnVaxfJJc/SsKSkwsX1pgGu8otdO9
41nS4sVVX+dn2xgBRnGZdKsFdE6Ysi2wUa63PZtjzK+Ro7FXVWkNVOkoL9upwOnp
T5p9S5gLwOMGAh1YGHslro/582Wq09IEauFNSd3tPeND8gpDYRIRMARF4jgacbR3
x1eT4Dei0L/VmSfy/rfuH1WqunMo4GG+ZjN7vT22jHJ1Na74T1tQIC4UYS96Z6BD
cGJHyNo88Ps6wcD4i1L57zjkslauUS53K57OS0uzYrc+V9h8xoFtEkq7P3M9wk1r
wpK3oMBZ3O0i3EtaFBn5iilVvZahtTfqYAxfNzm4nzntmNPTSt6nMdE1BSqHM7o5
dGLiAsuJghgQdn3kXNvNWPyaT1Cf/7lw9iFpbUVi1CIGkD6wCpY0VtA4/rZW6MAz
OLK4t9bBujO8WGq3TkrlAmA5xq+l3dRWRUPy8P82CqfFlUqlZAETqCFW//Uqck/n
na0oDikoQzK5tsYUIEVFImT8kaPUz/oxdNoXJI74rZ+1Vh9zrjCVY3kaMyCmCTG+
yvopGpoZZ6lkH0hHTfKjLVKTF+wkmfaJmTUEM+XjjoUg9+6Wt41BofgfmDHArLN4
IPQUZ9xb49b1V6pRsfrKWaj4QYq86qix3meS0XC1t42k9oWbK2OrLNzQznAfUFMp
sKMN/1lWa4O6ep3FmXKhqcBu/ExkqcKMSbexpoctseA6JfeLk+a59G2crmfBQ/GM
iuodgqb1uHmm1PAv4Y1VuJ+nLfdqxvjdablnLuVTHxkdv6AlSf6qDWczqA79Dh3E
ODUhMltlv8B3zP4MzAaDhnG2A6e3sl+bnLsO3QBLOvkwKXjHxfb8Ztkj8wJtEqC8
uHZElctca5n4aiqHiWWhbOrlmZK/LvCBAA67oqK88v9oU13FUI2NtQQdHmFxYY5B
l7Ol+drMXC/0fxeBL7dAqnl3nFkdiHvIaoetOFXbASN8efsd+NwV1WwbyLLWq5g+
YiyJODPmob827BGJKMNiCPz8UKjZq+L+XAqsuPwpUow8O36eTmle8xj+GbB6s1fA
3niNztoAbHauWA431cI+ulDefLHBe4RoFC6QF+DPoyV/FN7y6OmOUdD83UJP4Mc0
LgBtuWP6pKMNe61QqJZf9XmgkOTsb8Fog13DeDIUhV3AGvy8DE5JFifzWJSiF+kM
aD1z7tjRWZrAKW1KjHxro1tH2N79DQclSQCUfHVDsJ+OVBhOz3jr7iztlKWIDRnp
cXghi47XoktMGjdGHdCfd7S8imRGUiFkaO7Xj2Z538X1fuUN3cmlXwv8Sv8WtGdz
jjPP1QfERelRibGpUWjoBJ3pjheklZfCNF/hQ1AyPk6IMIl6WbHhhhH99hsWXQy9
aMLYsHliysYYlWBq3FcCgVqiHAoqLDxVOyy5EaPtLp0lJEBf2sWc0NbtNyKW4yEz
JcjkmPJxvZ/wbMl0HCUQ++Lt/LfcA3lV0mh5C1LRc+yStUXVHqIEbE8EZEmBYevE
zUimjatSxqMNXrUEVecxBiCsw9nsiwQKjAzIfLuRsASmNnQkZflVtHg21IcoL5zE
rqnVnalBPHT7QtHJEipqXhrfYKxGCuLimBBR+n7D0QSzPtfkvyXzzGjjUQRNZGHf
a0O3ljCl7YHX6aEYXyrYtnUP5tZBquvPUDa81BOdIfVt3BxizUHkiJfwsgYHnGFF
GLcZUqUVGl3K1WdiiCxFvGKbfYp7Rx1AnMcb7PA523g0LwSPxouUapQ2Trop3/tK
x14W/22dXODqRG5FxPf9cNfTOXSXFIWEjR1/4NQxB6UWa4U51aCZ6asQxWkKXIuN
VtVZShkxcYAIuHsnQ3XVrW156rolZLWMeTHjKg9nYEAzcveN5czLgaDeF876Q5Os
FnbnvoxGqc/gT4AQOXB4HK40giOFz8rY/emKv/baYp5whiZTHBQKUSj0DsXnjfix
Dp69ShEJF3v38qLmHP38wwJg//O1MlI5dX4vTz3Js3F9uk374XsfQPDgo5aBkTd6
PAD/JfTN+PgATLHwliQk+o+Ev2VXnrM4onuZxWLfJS8mi9F8GTIDx/XIy08nKcYB
XzpwO25EEYoxo5Ks+2Vyi9mBEh0a7Csi7HLuzrtmEpTWA7dTnUnOCRsHwilYm1f4
SE49fsk+NdhT6eG0BETObCHtSE+A1Myh0tSAI1DTWQTnD4IUxu8yfqmEPgDxLszg
7OqKzwm8K5UtOBzMDuDcNL8xQ3KwZgCK8CtEPsW6dTp1WgWJoNNjdTXLI4CWXUfL
ecfBsqQgPFP1fFWOWLqcbQeM0rFPflJ2mm3HCfGwZ3XpWTrkn04Stvve753dAgj/
fysQeZXgrnSMCrSEklik4hGbsGhRWxo/XVy9vR0o4Jk+GHLe+WZGQ6l9VRsLszYI
8GI9fOVQEPb3b+4mJCH0/yQA4XH4ALNe1g/DTg2Af6L6HuqJz1oneSLG7Uuj/XEa
H9SVxuKHIyzRbbYEykrsOmiHwCQlYtn9W4Zp4iYNi1LThbYUO/Ttg3BwTYusEXn/
1N3BiibH26qb7D0zOSLcU5i5Ay3hKgiNvmf5Vulvn4wHweZUkmxoNpuraMlsvLiR
tePEf44VXYrrfqazr9mQLe9oYsEOIpLMh+unR76MuEKXOb4mQgpHpG6P2hfTiexS
KI2PMSFGuHHa9ZGkWDzqdGqLMviVTD10NabhUbvA8S/caHHCs7Jn4R3nl1E3O0tR
gpFFsodrpWPPtNCAcp1MQageXn0IabqjLy8TmYz/S9vklF6LWJwQfW3uvr3USCmM
fHsrU5m3LaQJDUyMqryaHDwDnee3YCPB15E/bnhw/FiWuKC313ozrouGx75Eqolk
80716ttghcfW6vuAowVSch2iAMWVAyyuZS2Rgap1NNIqfGpf7amySggdpojnqENK
a8O7L5oed0Z71gy/XHksbPvRYTbQfmGdhm0V8nTDqfjSGVkxUhERF8rCcemQVlY2
jP1AHByH5YX/loq4VUPoMkZ61NIK0b5iqhoI0+GzMClAInKJFaUefnL6lPufc7g+
/WgmbFjddgqCp781v4W/gBE9nzM4Vi08ddAI+04R3K/WtasUtxDkp+0sID4dt8ac
JLsX6K7Qi0kqn78vg6qa2yNFg6yplGaCsKVASD6/KTmWbe4M0BPuAt6VzqSE+Rkg
0m6CieW+psYfHtDPNmqA8UD9cQOgssXmjicCVl0Oe2uXp9hc2o2hibf6gaBHo5cO
jYtnZ0wf1ZyIr9s7cUfbDglj4mJiwqT8PmOxIffdKvnz30Ela9A3SLiHJAGiibow
YeGqOlhep03yK3XDgNlu8iHzKRo3BmSz97AZzSBgXzPO54IsvQN5KkHTqnbHQ60T
8GH8Y6tQrVl8q1FCTvVpFM/fiLh9Vfu124o5TRFXmfVGuryXVN335rW4qD4L7y8X
xDVAPaWiqNYWmqfgIeAvmEHkDYTru4XqxXl3IOK0kc52m84Bou2WGW/HwB5Q9z48
35FR9ES66fHoopmo5bXdgL9jMppP248Z8fpvQ5L36jbHZ+B09oXljOtBJtCyq5bM
8Oy86XXSCjrvbaG+V2RR73q55Tjw54yNltpvAgcM0xJislwyKkFVIms91QyeMpQH
ouUw+BWjduF+uyI0pBvzykzBAo33O2U9QjXIrAmrDoxEDvRRXjP2kv0uB+KPmbvD
cNoqtG+ZnjIVtEnnLcjwNqm+gVNHhmHdOSwLAx2MaDxfQpzZMD0MNbhMjCRVUEXW
+aGRp1TiwFUcKszPvHqUhZwsRhgGuzQ9fi+egfph6yNKnjmVpOZpkQctOkOGh6ol
X2ZZRx+doF4ej4dewExAxugqABVfOtY7No5Uu2t0cWtJVZwhNVX78NMvMspMA5lj
lmTOUw/9PO1kJdAtrEPK6HC0FmQtPABIfeMOklPIERLTab1w9spkgTKZILWMGT82
EvEhLBskKbv9kDDhUEbYKOcvymCKqBRRN2sRHSuKzJ6EZQ6HEpnM84PM/kw6zgjr
xnC5neMvF5ZWCKP6qzJoTj8fU0POS6XTXkuQnRF63PcHVH6MINNP39Oflz1vUSKp
OhyioERb4b6DqGviHBH03XJ7SJAoHVQ8h95BfMUCp6KTapsxigsuBV3NtCIOrGzC
2ZB1EsoPa6R7KAfphwczmkNZzecEEQnIfCJY+Vh2h7mTStB0kun0WlTBsaCLLdYR
71vphAoYja4D2oiwcIko0bbMPzHCZGj/xytMullv86eo3LajqBm2aXSKf3gavMwt
O3dMfSiW3eZyt0NiSHkFOw0IGqgsqwSSQj24cOKxSm2LwgVHotZFUnBaleAgH3ws
8bH2b1a3X2KoYqhfk5oSxX9DLAJAao9gtAn3A/tejzmLTfNXT3rlv+JveyJ7NThv
HrjFTaUfbUYSwzkDlhWJZY2CVryYpxdYwtnSnnP9N1V9pLcXn54RMr0F3FCuPm17
mmOSEFwDgkT7laTCX0vFS9rzoLMUsNbCQ06VMnuvfMg5prO/T/wgCmwScmor6zmB
2OXS6NDvFseQ4SohLcCLjg3EnhncB1dNkG5ohR5j+NpCpmesyR7n0UgccBp+/N/h
V9in7/fkj6M4lB65VaQG8lycOFLbZcebgr/ImEzOTJ4BZVQsrtlUDeksEx7wFCbO
cVghPfmKqKVVUhjV2hQzILTlSKYU12x3NZU9Q04X1mgv4wX6RygE7ccXnLJ3dGzD
fzIwBJhsbgsHorEZMaKM3ANnph3j/Vr1hmZJt0lYjeymKUC2sKzADl4THcPdoFbr
OGXsa1I8c/wfDYvpi5C22g8oTT9BVG2mxUAK7ozaUItsk/4rEytn8s+gAjcms6cB
vOhnFy8qGjZvzH/7EN3kj0NjJ2kaRwTgeYZ+PVpD2VSnwmWPeqVk+29cEHvrc5Nd
XrnTPW+XxB+t0lm6gGOOS8FdLUbaR43v/pNfUciATYVdEeJ138G1+fvecpSeYr5i
FetoIisg46QWBFN7iSgMtAe+8OsmjkXIgwew+1RXC2eh7ls1f6MuLddS2EQSESTr
5gwFpclkelJs6Ti3NrznqDjq6i4PqabWn0FP1ayJXlhXEFnCsZDljOwNIqoZBBsV
ADj2NH+aXxIfby30zK4uKiPi6KzpdjYq66IH1ch5wX6u/go53FByKeEVEJ7dS4YU
6QxIbVYG4yDTmlvKknsh6Wq6SbW6wjOWcQf8z8oFdPyPKxDHaBGAnkp2OlMq2UbU
7UhGQgLUEcemIKh+Re8AgsQz1iJLoeEZ1c5XndAekhEXCXsh09lFgYoQ56JHOy0f
I4wlFfG2N/yJdytuUpYpnRiQai9wv6Hp10DseielPr9hnzc+LRMjLvpAqgD7dyC0
XWAbgQBiHBfTvJDcw6zHl+9/E3OVNvYUpw8KJso24t4IfB+Og+6SdhNs2zV5PO+Y
9/3vxTlSHOmFoy//VBPGPq3uzHCU9ghRLiw4MWrzmL6NMLZHHbB8JMluTEoik3nJ
WHcwZCFsR/5ev0Fk5R9tcMffM5ZcSZcN0+1zNuLF0r8o0l3iS2ugtg7FUCQNXn01
CMEbYR74KL+Vc6AYe3tM3QjoEyOUgM+VbNXDr965rBotEiYsqGtjH4OY/D5fShgB
t+JI2tdr4RgrzLjH9WXXMwtNlJlRLrt7JE+VrTLJ7LdX4Wwrq6V66B3KbD1+8atT
Nmx2RHhdojXPzfPFnCJvfbPy+L0I3qshnwn0mISMyUxiqMqIARpRI8Ju5gf5Zy5A
yo/VgUWaAE/bHQtEWSwfjvfrGSEIW2GBiE7mC8+rBSMCh/OZERZhpVNpMe2zBwz7
OTW5pInRqmsnQT4lRLEqESdl6kvHdM2sFmn8EJyeL3AHGlND/JCWJRgi+6pwnsY2
BOwfaPMmIno2ciPWXs/eU42o63mrHp8beYwsaU1o3pDsT7RJOgF9/JWpfWq6aZB8
0SvrKY8kRy/EMVb3fPFp2VNJiFPFKszXWZ76IsLeDA0VFx+4o9nasvFylKo8Q60I
Jwyhbe0wwq2rZKO48mOXiGDmWlx0hWaDcP6OXAJWiTBsqbVmDv/CjPrJ/VK/EC/h
QDbrWn0thsFkN/Mf057OZ8O7jb5+swIGbV/yGeS/QWIwnAD6Ymebvl+OU6lRKGB1
TosxkL4NzlrW7rivU1PmRPePrdZesHzwPCWcHgej34XMDQ/KlxxwbNQvlVXEJiih
WNqP/gLJpZItrEup3iqO3+MJ73Z5mBhV3pnMxfVtbGNFJsj6Sf50+9YYU0O6Rkwm
wpsB6Ag0e5poYPvWLWqYHsxdds2ZAHtsfpR9/f51RGbkkCP5sk2iFGgteDnmafQB
SCIgK2pXVquVJIK3erkeKIwjDmnbJDuw88Bqi7vio6MujOl6BM5tE6OvCHWA2IXO
UobCZCBs62oQnF//wUeH2kimbCIrsfkSIhiaTeLiRMtxOjqh387oyuvEj/xiV5n1
hpWLjgqIkVpLgZz2bNi2czdabOIHmFYGalJJVJau++RJNNoSEeqnU7JBFYnAr1si
Hmy6v/8Qc3dVbacJl0wjPpGre548+G5d43cqQX22piCbaqB35ZqmzwKF9i1qU1sF
T6OtvJyJYTCs9OC1lRCKY/H17Bi0B2gdMJBzmjCKX1UNBZgf59z5B1O67kqpvK3D
kYu+6Z+ni282cP0KHZNl9tX9vP0EO9+rFk4cCOPZKymxXIahPjMEFRNaOFZ7HXQi
VgSj4OQMRsqOAw0zc+5jokujMPfD+sguh6wxAXCVJOgJI2wDJ7HDHf9C5QYGQKlP
mtX6C5mcPsloZVxdGo4lFpQiFtDk/MSKoi6MyMXKW9BdzQ+xZLk/WRk7HgYX2SKG
GVFiX0dy+XkVZWXScw8OOl9Suqkt1aqrwnqjL114FPJjnDiGi6iaZb8YwlUzRa0q
2DumSxKceMZDzvP0TqWpzdU7jEjkrVa7FH3xAbwfv9EOGgES9h13vUTBgjHfWdWa
U0bkaLkreP7u+Na/RyGNRv+Q2d5C9hskk6YY9+hdnXLTo81YzpZuZrGBXb+dhPhr
jgSJIz/BnB9DdMXKbbu9f6qJc8LnrD29ybQiNBDqUYy9qtV7FHcDOgqXkQlTUaIW
xndCTvLNvZApYCIXDlL1k4Y3t8XJ6sd2EkZUfCX13Uvd8rSAp9vNppIkNvhsjqVR
P+jFbmEP/2JMqLd0qtjXtsuWDQyUQD9rl5gnLpWVMXHCs9VGAOwLN8A2gcoz+OVn
6XBP42oaytZW62pDeR1sVeRcZ9xG3sYUPS996GuBbts+CSpXdxK/Z+iiRhhpW2Ux
9lBNii3v2XgN3oNgml45CZ9li10vcG5WhTNoDes/Z+nvqF30etBGN+x+KcjbYRyC
2UIC8Ewo/qHO/3PQLOOREMdQNnaM0HQKPhj2DxE7KMOX1WMkvSQWfPA3BuNXhS1k
r5UGKkIxgq4NhZDJ9JHAO5jK96xeAADfPlp6sJqVZWuaoOyqzmQXsuOKS6d10ITz
RwMs8Fm+DWPmuc19azeiR4edcid1FwX27flg14r5iOoQ9Jw6twtYGdZmcIR2IKvk
qZxatSCr/0yAWiSvYtd+bDqEZOMNDgyBM+/tnpHk6Q1+Jd6C6MrTT4BY03HaIfRk
XUFubW+tY1pogKePGq9qXeOkVxQojIEhxhNLrcZSQ1Vl43TKFZ/jf3v9AMPP13/0
DplRXHL3+Uw9Z4rV30tGy3zvF2sFGTggM20ae9Kfgw6/ucWJxnTNekvOY/2XPJNo
U/9I6C6MuuCEiVrDll/dXLXzlNyRiVn90dw9RKZQ81dEwuhXkceoVirYYd5x8Tg5
5wBQg72r7Ci20pO1ELDBCWH0uGRcMhMKecyxtUHmvf4in7SRCJjNOzlaNlfUSAXf
`protect end_protected