`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5040 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
rt/3AmmLaDBatPBsuoIl3n1A5YmUmuKll4vi2w+vCpZozxKl30rygdHgt/9bG6hK
mDQTFlhbTcBUtpvWTJ43jp4I5CzWFWZz0qp3aOg0u8/RbuFEVaPMWgA3i70jU1g2
MCwXe1zmXRkQ3BIaU4Z1z38fu26iQcm2ierZ1Gfn2jxjSXCVt12ZCaKoZ2PTDjlM
yE3jsMQC3e4lao6ayVwLleCU77FsCt00Y7XA8INFQRBSH4lPkWi/ibncGsFT4j6E
CTeSM4d/nybejB64E9rx+lriQBM7WhIH60aGSI5tEdcuN1kfTZlNT3rPMNGLh1sb
E5Fkmt3TFNiHRx1HuBrThAOG0LMJsYp5ux8z/jZDnU+xfgMgjYmwSFxFlHIble6t
gWGS1cStQUVViRb/tKtcjdUQtwqytQJzbwFsReLZekhLg/dW0j7AkdoDjL5h/tuE
C8TXZZ+HkWGQ7Q0lKydUM5ubiQp+2J8gSDVbNGnrrx19t444SD2d2yHD1igdU69y
pKLxW5fKUf7WpQ9qAwTJ3blh+Goe0phwhJPYiEIicZ8gGfnJiuxXLxs9uQ1ieF1Z
5+dDeMl0byam3c9IXeGIhvuKYd1eyhjpD3O1LOeCwdw7uELkH51O/tv5AJ+LrXrC
GiJqAIb2FTW4AP1z+R85H5AU9A+zDkwKNtLRaHsFtZvtgFgWeMAG5mTnHs0uAGsS
6JrVNGaEXKahnB2xf4Zhu2xQBSZcrsl0Iq1Q/UKXtI2FNt2DlkqxahMus87Hr/id
EZi01S0Z9lFE/7ar5XzCl+jxPcYXHjx8K9tp/xuzgeeNVWEveOUKWFpWyINpXiNR
Lf3r15iEopVx8pzgEr8RyETmFbUcAZZBEDmO+qXJzXyT6q0JtDbF4XxP8GuwgUWp
UhLdgKRETN0ulE2+vqfyJ4UW4R1ieQqtSTwS9CVgp6GB3fF4KIEABW60N4DXOR6C
BSnEkPYtZX6Z3KunyO+hRZg205lE8enjrcFVr4ckDC0CpeongiXrlZXkYi6g0XvM
yFO9beThrwpjpXE1ZjFYF5IfGMOHrPktR6TfVU9S3crSrmUbJBDlv482Ht6Qtyu/
8uz6GUpgLDGeJPfIRo7v8gp52x1V5T9WSSswaAxs/4ydOG10/DU1/rD1fZTINcC1
0UwMn1ctXay7onV/iSX6qcBvXEVVMQdMCHClvKZ70W8qNALBFQdhPAmSPFDRBbUg
TUWqFKcbXAIsfHk4yHdnyloh9c2s9/5OGPR/2FfIkpAPgx6l/3GlkvhRfKrqbp/r
8gLQEU1nR1ALQAMDx3qgFO/q6hA8URVwKiEOAB6syt/lDbqzhjR6wdW3qf5bUgn+
MZehxdXhkH1jazWIZeR5rwrR+GEqnduCv3PWy2wyiiDZEcDWk+PE4uNot85b50qh
NDsFUJ2etGiDZJb4hCMpylP4Tt0rArMXelnhzWVjpd6NGI2ylz1M0f9gLW5kDYxA
gecuf/k03bFfsP+Z/E6OnBWsSDtK9mrYMuecxJr+BxiuDsFBsYCqXReMnMvJXLdJ
ltE6TTOTdm71wcxpSnKUSxQ8QzBWP/huv6jEqEZZk7Wo/l3Zgllya/XRNwzq04mC
ZADLbD8edBpM4pX3hfzLW+dKd39qp3BfDn3xhggZnWbsGpPWe1P8gRUO2GqJap/q
4tq/K2n9GaUQEoyBWFCdVVqSZFeGegP4b3U20QxKPx+V3rPDqCsgE1O2S7POMpla
c8CBj31Gzk+CfPsTaUfaer4sqKUtScFzRFU9gRr4T3H/kicxRQOPNdtxm4pcjFx+
t476xG1fE9ghGm9nG7WUacthY8f0HtuMJX7yx/agKn5NbomkKWNhP/QCzKxqiAHx
qVmS0IkiX+xLWmR/DVV77FgLsscwyA8A6GynRqcBZd7rrzPlsv5bOKAspIcGKDHQ
C98LtdbcQYeZQPrcNpdFQ6hs/+Pld5cwW+py9NNLCphSVdhCZm+PW8m/lCj5SZBy
qqgxxOzUS5Qmqp34E1pOp8rvM1TY3CtjBnNHvtvwt4hJeKod8yzWEo/xstn/N1vl
Uh/wXXAhYj6LBPJZaj+79gRoDBmp1alweLzTJzaOGgsNMoY5jZwkMy8SJybnqh+4
Imzp40YHlJ7syFsbqOftcw75RS7FGOADSJDtKhp5OegW090tRQ/uVXafGa82lsJ+
tAOJ8WAPYwEUurloNuN8en4ikZKuz1sMcU1EF6kv5NRZNXDsHLuR0DBBcGLV6ulj
RV3f6qqLSHPXEgsSmRMIFX29DCai6K8wfOWzl+/oAVZtZzLNQhYV9bPZkw0hUudW
U++By8hARHAYzMiu2o4qaL07/s0fw23YEVfJLTW1FUDbSoGKoXaRQ0pTCfcXI1BH
SYxukUZEQxlyPhP95oZMsbaoXna4PsMG70dR4X9REpgtRBhDvsz3gpmsBavUA7a/
jbovYEHxOK0ceTY3mRZ33LCrOivGBsa4+uMF9GU1qL8ksCxeuQt2bbXyv9eFcusG
pcQb8LJhC8PXeLoeC5tA2lHG/S+9km9ZHp4Qx5H/ftsAqs5duzQ6khtSix1IDZa9
mvHNV32Sj1+G5NjEb8jm9j5uXC2HqlkiIFG65wPfBtif9xjAm7egfDnUPcE1AeLn
tHs6HUB9+4p+h2cURsAQrZ6oSNyzXD1+Z7IH0wYQDhnOekWYeyKGXzAHJ+UWBf1E
hlTSHrD6GVfdW+EJX4ADQIX7MLINxUZtr40ZRWhxg2Bw1WrtCGx8z6O0GVWMkoYN
+8cnJrluNnPPWNbeO+ladMdNalourbEHzxMhmFOrz/HqCTMefPjPbutgOtGeyhE1
kpa+QeeeZV7FXJYmHuM1AY20KOxaM5fZISVJjMHpSdJUtFc7Db4CJhuJKynuqw/f
T7ULovRfnvvif51phygdsQLTlkwAhnyEwFqSG4xXP3AWxtFZZlkuhWn56VjDAvCw
UURBPLg4zkPu4nocfIQkNtwQj5+hFTV0fPDKhC/BTGAn8gR2Ov7CKUEzLLfFcQTO
/4eSBL1hQkkbx9eqMsEzRvksBQc90ESvAEJ7hCeh7azlU+HlEkjJxN+gNyN2P5EO
VOpITKWkyOnXw4d7pxZERk70s1M5JhHss5Q/lYjEpDKtP1R3RLqKkVdpXG62cld1
quKA3Ep0t2JzgrF1Msbi0sSsd7f1tJyhI6RCfN9dSfRWPyJDJqQ/SnEb3xwNAtB9
jzhNu0FjYThQgoZNMsKnPJRuO4arwtIjR7vfXFKFZ7W+tJKR1yGE0IV8E/xZQ7Lo
wheZ5SS0kHz1v+F32YCxOA1JXWU9JlrnbcNlpSMfqQV/d5NhoA4ruZ6yUOqSY2j1
kxlU0pf4T6qib8eM+uv1qvgv5vlzyqIgWmyHmjmK1/5tuqImWXxtdt+ARbiSKgI9
QV3HcKtnYmzb6mAzYm452oZxRwW/eKortb6EdiVsy34LXWwOPtNnKnJtcfjvoHF4
ynzJldsFqXsyBDEwv5twj+0iJtdIGjONWEk6EVYqFPigq6WwR4disqiLvfzMpK01
435vAtyFRKW5fO2rJxiEYq9TJNnhwCehbRuo1RPMhDhmQrSP/w5SJlr481c3raxA
61/CfzSq4vGXF/iYj/zn0zZ/iNqUA5lOMWV3Of3VMGyDSPkMOx9HUcru15c8h81c
t8f4tUsueo0T4YSG93iMg0RPaXWxhaAWW7QNn0528i2/3Nd8Ak7z57xpy0zj6A2M
C8mpdd2jL92kiGSXj7FEofJlcO6JLmqlue0YH1yViPYDFlwlA+IrZvXMjiaBQomL
5Y6g1CDRLGYuJHkHPiF3fX+8XJd76G6xRBmXLxVFHkgmQjqvxtDrtZ+5SZOM2ZjO
mqWAaq2QMAHNHfI5aUVC/ZHOYY0e1/Tu2Ox907I+bpfxwKuDfccF1j1hec3HK+Ej
DaGWCKsv19cjeNFwroBusFbCi1ruuDpygRydCGr1+0YpeaNpHDhOrxMIk8XKBf/h
9geT1Q7lsj8dyo56dqdgpeiEQqbAUtIfnI8bfm5WFGU3O+47lV02hynp5e/9Txv3
DvHdDCI7doI1nyQBYdOULqHQqgHeEYhc0jn3mQPGlssgggEx8KHjRGXA4hPPCpm/
0SzRTQPiuIhR6XSW9QU0wLAjmuZH/eZZ0cn2XkgBfGPaNHD+reiqXKjRzljhRsX+
5ECsG0WchwZQdNPM8Ppl3vGmMOkMrd3EKTs0mHxxDa9mIjCB+HQgsEKZ4bK+8GVt
kn0dhnx1HsN5iWDgeefq8JpvymBCZm0jAQ74YVRgQet97ICes4fQt/wXip3e+O0g
sAsTbe7AGZmeSH7UCHyEguejTfa3N53P7GcVeX6JahsnYOLtuD0VaCHbhDbwqDLH
iXXgM0AxzZlpJZbJwfKnlkJPQ/jmwA9Vb8UVfTifQE69RRiHCnTTY8qR18ElXPmx
RUlmjgCmKYClXQnckL+ijpCCQ2/WBM8b9kyg9MrWfA72w/UEZbCzj5j4O64POeJ3
78jTgUmBIemce6NWEbT0fQR8oA+PtyhZhicF/CsxR1w0dmJerxZyS5ZKxKziyUmm
j8XOI1A8kXAkEO+ZFYgmf0wZtM6UWkjPL4tah4B8jNZFUjTNJZWKxCE+7BFTkvqk
GlX2hyJ65FH2MuRlCQMrs8gUwdhp9bIa8h9w9B0JQc5FH3QMJxggRozLyt1CEkfV
U+czXXUeVKCE158O4U8UDZSrpIN0uqfq+b7+Z31g5VE09NnDc9Yka2uJiKokSDMm
o00rjh8i1YjIEyFR3Ks0tIib6s0GjVX5CZMgKdyxmZ+qFMHrRz8KeKH1+zSTSvWy
wE0yTVEpSm6d8yKNzR/1GF5dh+CQTKY+fU6QPBSDluR1QjBRZs/dEog5+FBH/rU3
SVzaMsUknH7W13rhiWQM+CeSt3Uw/4ThzrBizA2dOe2orzR+jXOkDMWWHcF6opqx
slUofPXXx7soZIc5LjBXYTWf9S0zHedBJVdFVnRmOrtTDfnYKfgsg4Ya5oaQqGOo
7kebXIOW0jkwkL6TOHm+rE0PVVhPKL/HavkYjD8jwnL4CQLEoAfDq+Pe4mcc7UHx
YCksmrFD8lL08TQmtQjqzKsJzEww15an3mUXa9nFhXRwC5ZnTXe/6UVCa+xniFO7
Zkr/6gRu6D4vRaXiWW+EcVE0Zc9Xv/vM8F04bWer0bJujYHPx/mrqGJ5eM70Y/k0
ymD6un88g2ByDLQjxA9JLZVrfEuHDOcfJRXQtQvmnpzWuipg6nLl21mpOXt75IP4
Y61XwmgyMH7Z2SmbxQGzdcgOklY6ijtuGihVxg16Q0dPTNYvqxoJPrfAxEUdplvo
bBy+U3KqBX3Dnq9e9Xfg8Gu2/45qDH2hWgn6Xgcney93oAYMuQ2wd1H1TMoWzxS2
rjVduQZH7QDwBoNnl4zy2dabw3KRCYb5xXlBo/Algtegf2P5Kmw5jy/5Es71V1dE
+ySlkFe5g9YoVX/rBcMjkVMUk92V9iF1lLP6QHYUmEiR/BDn89NQdE46QJ7JoErD
ZyGYoRwg4NmDAbCD0PapI5fdo5brdyzYwIhzPnaIX0DqSbP1R5LsSWkn343BscGZ
ojIaSx8e9Eywmk3EXHwbqC4LYflUmqnnwSNXJqogcZCXxcMYYVQOLc7BWbhxdDM0
bAsH80o/7qC11oV1WZIh3JK/fepxodTFYqoMg30z7DDa5pCOoD9GFYWtUpouj0EF
W30JZuSPhPs1UU0j3o5lLJbp7YtPqa9mq5bb99aWlDNvX/EnVJ9rH5NtyMNxhcbZ
A/ueHyUPtW82HLWC3aXvwB0zBgPko7OR/DGszWDE8C6Vm3GkwWBGsVkOU9Xrn/HA
Dm7UUFUa0ZpYhgEQEpxE22FCYZTEAiiwiGBKC6r7ZDBbY60nuQqq++vGJ7aYZ2MP
KtghbCNz9JRsVFKKnWE3Z+91gn9Z7sC9v7dRlMtXTOUTTdRj/ILzOUYxEG41oEU4
Wgjt1lxnsczVdUB1c2E0bU+HLPgvpP8iwR7/oR3U+EcIi4wG1mppPQx99mg1Ao2Y
YveJl+zDZ63J1IG2O1L263iAwoEEPz79HNlCFEytHRYHK/q5fb8IlPU/XESWUT6P
u5uzTseE86VensZe0xPzwjQ3AV/Dc6nNbhSjO1/xM7oSF3Zg1PBwRvUx+/nS6WP/
T6F3lHwRELdAhBRZIciy9bLOhLORYGJWOK49eS61tFM5yjDIvU4xzIGJ4F8DdXRY
pPfcb+LlfEprnbv1E92l2HMyPd5NybBp95lLiBFzP7GaQcC1NgmqosoiTQ3167Nd
sacnviJqsJ2U6l6sNLjaneDF+a3A1Cd2hhP5+Wy7ylL/augSxMpctQ9N/OFYFgsp
ORxLcpjB27g5icqVekmI0dktqkJ3q2aTXQiV8JEaxfV/tDqjvLnru06oMqR/1fSJ
5nta1qFeInhIh0NsDezGp5nA4QNmEVIhA+JYi4CA8Supi5ZnFLOK8BLDJ4gEPQ4z
OOnZyAyWgEFyOCMWQzWM+zV8Mxsn7HQYP1o/16jDx2pTEKdbKXdHdmpna5sFy+6Z
dGz+IkxbFTcVogw6823yawcOjxCCRgNBdxACkGrQHv/9q5dY89Id40e5Hwm8dftn
`protect end_protected