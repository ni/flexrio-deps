`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7184 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmWdo24EC1SLhDeUV9o12ewQ
ulXp2xSZ5P2RSggIKJUy/anaBVTumwtXp6e/AWaEdudCxCx4R2z2MbSSjkgxnkUf
8YekdUNzI6HumgLqjqzjb1/3CRW6P3W8NhdbMmesZwlz+yoaLCdkbDkutUiVsGNu
N18oHeoLeA3+LUFUOdqIPpGiG6VWgj944jRlBSD6gOUu0nBCT8q2mIE9oO5faAe4
4jYKxcc7zDnnldz5CPpp4fCn0+r59w4WaHqZTWKmqXn6oNZg53N/He0ZsQAvoRYj
7Mji4bmEw35lomqGNLWky8As+31DJghiPNHa7ZiRJfTNOypcPWqWP/axmDq1mEzg
tAtIwavpYFXRWLGqfEHPS8+2REflmGIpXP/FEngTZvMxvOCbPD4wV39J/enJmJ5I
f8IS48qFERLzVDxU1sfESEA82zfSvHiia0DgS0Pi0OpLlLCXRjk5p0Ktjovlo2lk
DBf1WyCCsQ4Kx+6xEMjOnpwAwstC4DEGsVxgaU9KDnk6gxkknMdJGNeh7TUA2r++
7wOSH+fJV+6Z8TC3R0QfOAQen12Kt+rQ0KWdkychx0oajFL4e5CX+qzqsJXeUxhR
SvoNROTOuospvIsppjSR/E/fCWw0ZOSATPDYQt1Ek8ANJonkzfxZ6uXabk1Eq9wC
Fceqz2k7sXKr18NWFJjwXPPFIX1pN1po6LyjDAW8Dte8pcwlg4iGxBRVjGIRfz7x
vn2PJTgIWujXDMVFgk4RlcGhcEUOmcWOrEJL8yxY5zUT3BdDNBkdCU8QuCtfQdza
0vllPKl4hh4pXX+PGb3sS+Hr+8iF7gC095z9mguYsWgd31ky17vwrrch8isL7wVt
A8NAWdcKogb2lYy/FMK0Yg5C9vSVU0zoj2F1vfiGFybh8fLCJLVzX/+4VduCfdhG
kBSxzHrfuqxnRcP5hK2DL88huGtZuvoW04vJOcnjrqj5VG23zeJ+zV2iBssiM1OM
gncUhCD+j2p9Bd9xrpjD/W3FiAP7rcDPZMlQPcdWBfFw7ruKOyeHy80qBzOHepyq
kwbI13aXRbYMYI01LMXFKBsxC1qA/2bKXy1owvH33VPAMWXOWblzQcOZU9Kd6ktc
FpWGhTY4zCBuEkGf4d8Bbxjvl6QUtbr8TMBeFKb21jmtqT5qMZzzw2nAWMORJhI3
AjSnrPgLtGUzIag86SPkUQ9tD9RISSZD0HH3FQnXjxYLBLvj6OAPIFb+BptrtnUq
+yQjZQ5YQXu+2vinH/J/HYMbtSi6Lx1hyOZVQ+Vnyl789ELJBlhcR1ln76l5fLbz
pLlbNH6osnvXvvQmAWZc2rex6J+1bA6BncrdHuSLkEGjCFaBR8ii5RtAEmA4gWvm
SGC7bkI8HTyhLjR1mZK/VEpxBQRMljDfJBYSpWdhOFUWSD3UCVaQGdqOpPKg/B6R
I/aXlXz9cWHGBSYogVh9JrZimT43ppExyJbKvHpmwCFJCdAnYtSGWjEPoWbB9pTk
+2Mg2+YW/VR7cR5AuFXQeL04O4FTmNyR/mvmR34L5UMvIQvHCqsttFp211OqcTFS
yazc/fo25PLpXweelcskEcHGa8If3xMSvUXARScqf4dWirimi14kZCZJXGmepJih
EXIZ8G/RFPaARu6hUT+Gp60oTR0sb1BJ50J8U+/IZqYG0lG+5q0ORbzRY5QL25Lh
HekxTQ3ktgklNvHf1ApfiRttyXcwvLIMQQznYgpktrCJ7GceXrTCXJQfTbMD6ufx
LobEve6LnhzTfnA5PBY4rbJzdZNdu6Z1HqZMicQKxudmiGRukHd3Xc2UcUnAdQ7u
6JNBv1aEb3RAER1hMi5H2LyjORHeRTeUzRe2zXMB7feRZa0tUlCTt/gdVcz0wK34
1y17HuWp6e2izLi7zCTTAJ7YhygbiI6ryTbdI6FDOwbm0yFIjkLgym5r+NcXZmjQ
pKhmEH3Fnm/R9KJORBC+EPXicXCQ5w4TMLBW8AO3nNQFOQs5Apn4asF8NG/WFCDq
H1XMQROBSElgD8Gw0QqCm4DNqbyGcaAeFIFu/C1ZIRiA2MC2hIYEFsgMCfII1epT
yfl7oexMvA673Jud14PFyKhOCy21pJEwxpmPQ77bDsCQjq+WLIhfjkmCvXV4qr7e
gjodwWDePU9Fhmm5oUn3APB18J9clgn+RODf17Mgsf5u2caRbswFEded/HpWuWXY
LtHYU7Tec5gJAun8BAk2Fg+w5Ell57oWXPdIPNK5q9CyQGw+VeixyE2QNP3zJiUN
Sbei3rfpISJSwhTOBVMFl/C8rrSGVY7clRT3agmecMbdkNDSC2lQ7v0RXSkbjyJ3
yAT1XGQ8SJpfeh702Uw4hDXMkzB0nQMiXztg7gW0ZBASAiApYh3wyNj+6sCelpMN
Hltc/71hqFv7zYHsAhHKws98ZVVmoU7aZLoSY7ntHFLB24fyhTqgD6/c8H2IZ7SJ
3kaBCX4rqKEe6irekYgqNljcU3iaOt43/0unaQ0e/17OsonpHny6sQH426ERvyc8
WlzK6lOGEl5/f3fEjjjk24MbYqVE7oibum4BnbUMOQ0NJr86ZTTWgobTMnRvV8Qm
/pFIe50HpUFv5AHScKLID4zMNDIf7ksnB2Bwp2xhG53fL150PEMrHPpfEK0mRG9v
vodnj4DpDsUE1tNYEbOazTdyzRmhi3AdnhHWy17SxmlixxpRIT6IQ0N4Z+B+bM4C
wGzGQK8cP1eJM+5uz1wpUQclX7H91VdwQ0rvNlFtDQczIOkEJ5aJIYoBD2JEG7qS
M5SEbp5JvF96zUW16wrBddKiYD04pQTFiZAsIPggH5kNRy6/VyvUliHbF4P6LwtX
xd5PpwBGn4/CsKvr+TjkDiMGlHsYba38ho8Q5xETtxLoEV7fPxvtbdZf3VHg3hKZ
lt/nVBQr+Y4OtqWDBlqVYRGZaCWta7xEjt9WinHPGLi8f9o+1/ZLYCAOkySRaoW0
H4A0mUwnTqU50/wKmrFGb0kZ4y14jpKAq+dEit+NDsdBVFX2qdc6SsLAiC2JrQhX
hfelUwwULfZU0AuETEiGnvz+UO8QJMc3Y38u6VXPyRqSPP7Fubn/FdhZpFzmzK/x
ziwKV/G6SFUckaPPxRT7STqWAfFR7f3mznn4BWx6Siyy7Df64/6LpeIYb1ayuaMs
S5e6q/bBhd2xnE6X2EHm4GkJc8dsC8P4IKe8RbHuf4ENDUxR84u704kBOzsoUQIF
v1cxLcX7azmVocXiA9yx6Whgb5aHxSSeokG8Kndzx4aZBz/YmgkACDihSgHNymsG
G6dmey7N+zFHRZQsoY3sUqhysZYy3gi7cW5Ki580JHzhyII1xLuiLOrz6vWh4vJu
FExNd1/3sXBrXqsowdPz7gYJoQQRXQwE+lYyKEDVfkiDSX2e48OTl/gk3Z1YKHzm
ViE1HUnPNl7pNOaAswz27wVxHaC/43TqCpfx52IMMIkf91ZZI+obIe/IiYH+QSS2
/O5LxoxiTqNOEHwqdAdRX0DOy4e4K/2rHS5vuJEKPM9c3ACSblhdClGU33i9bqDB
Rn55WFsfJGSAWtSqYotIVKKs3f1PEJcxH0zlQCJG9kwTfak8pY1+lhpPYAw06V+r
FImpXEA4ggGwsqCiCWrsbr+lht94qIhdsQDSBAe2X9p0T8eqqLG5z9+4QIGZvbX+
bdkxUozDtDjKUWjkhD5Q9sqsms7p8NBuw2jB4KayFtNsjOvE6dn/O5/gn7WVnqUo
/mTCOUu0uDMQFpekuIpg1lDSRsQTODJBSORbB4074FPzZPuolFsSnyyVNbIB/Y6N
2PX7BvDoPuDs+KgngUL9+Z9RlMILNiIxGAdlHjHvLwUZJKFU4/PdhILBpQTuQbLx
uawqF16ZpWkkYAN7jAeH154YZiUazSg7/02RA2SGUpMSDKWyhniaLuUkiEVKex4c
h3dm2D1aG0rK9Jri5wAuOAn2tdP2azLRw267CW74uOOc8HZiRLuFrcjwqiHJQCL9
z3T3iMH6TGMnhuX3SM73RLkUlKCOSiFs0yKLyfxqul8ZExgjsmHr1GqaEx0gGany
EQpC/5RRllilZY0mUilfLhRKguiKkZu84i1zA0AmllG4to/cGogg8UlWslDhL3lM
oDmwt6FEFWzgLox/rJ86qjuWbOJiCuNFVEaaD05DHCtDciL6inLNlrlTArB1V/XA
xx0xzVOiagsp7l3M1m4RBl5opZl53kkeCwH3/F4C9AIJRH8/1MuXapLc64N+/GhQ
bHPB8kbi5UT85tQqxdfeG1DFNoUd4jRYZG3OnLwkS470ygQlo3pv/qxzkkKTvBYS
fpJfnx/Qwb1cUEXhKVN9tYns/hKWEnJnw3pFJTfnun43YozEFszXC619H/Q6un0P
3w9Yvh8BR5MG/UL9QweRTMwe0YisT3EVHT9hMdeM6oDoHbkToqWYPlrBsfh3LAOS
/MfqnDuTAbRL37sr9xYMNjYb/7jupI4WtF1DduSVgkFZ3QhdY3yJGk2BhhJdfiCN
uGkZu/PFGdekEtCXChJOvXJizGr6squWCeaWq96ool2INm7/wG1wzMH2ERK9dCUv
jPc+lZvlffeprdbe5v2/VkVY9q6boza/BB3tyHtIACTpqCdnbhOSHLYkcX1qYn5y
SWIXFYuR8tsN+DlazSkD2ai/NlpfLPMRCs0wCXjNUDr/Zm7o/Rtib8M9LGVLbIQW
mELBwpbYmunYh3l6QzK9MSisq9+DlqsqtjI/v6sdaxWOXApW4sqthFOZc4Dg4ncj
D9oc4ClhvzEgIzUw2Y8ORuuooqjfJ1LHEG2GBgJ4J+VP6ytkB2ieDIphQJLittJc
dGxxtgvEL8rc3D72I4JIpB9diQyiTL3oaDSixPxPXYYzA2r0R4pAFKalLUSwVUpP
BP1WBw6Nv0g63rJZ3N5wolTeA/h/L/DKcfHmyQrRS3rlYtmLv1CzJNIS4KprHcP7
LUmxCmvqbnRhQSrsKfrCtcHS2Hoh2G3Za4y7gFBWWDJAsuytYMrV+HIA/Ld+0Dcp
LzldjVEaiFrw+moPPQoWXVzP+agb4OTh8nL3cYHS+Oo+IPd5thdK2nURAye+iVCW
CsMiQW1dCqxkjp3BumWLvAtxCOmglj7QvG3mpak8nZSkpq+niNhAN/3IERs+o8ry
G/gnUGWMC6vbxPv6Xn8AgPyfuTLKiHdjFgfz2PS6t1ZFYCamdO/ClZk5IJKiYSOf
Twgw1q8i6D0X5wbEw/Eb8tu/80i6a2JHwsD6ca4QilRKoMSEayxyZU7sMdBVJ/h1
PtWp0quD4f66rJ1TvQk2NHByPdcaxNyibHKNLXbJIPsYtoa3EkQIgvG7mYuDUUla
/mwYo4ZJmnREY7zsk4+F85jP9sLCg/lTRttxK5zCtbbN/mra+peNGjl4GG6t4fxX
+MqjehUEFTfoBQtUoOq7FIhoK2JFMEmQklLp5dcPhpALCEt0Ok63iGwe7jHp0u6V
8iBSid4AQz7myYLvTN6LdK2nswpc7Rqd0qV43qiu3VlVQgkpLQNJ1oTL0dDHrnBN
nXCrHNSluROYHrAyQmMDmqNyHaTA7u6oXr3ki9I8Kwf6+vNm04BszaDBx88skVYd
wZGQ9yuw/UcF6DezD1dCbl3QpYXgpwiv+lJlUbIPYkMO+MyqskUDW0owi0Z0nMZG
40jjzlbjMd4KXFhzOos6A1Bgb34D3oVrsIu+C2RBldV49krXh30V/1JBNRrfEqCT
tkm63jWd1+I/eHAH8U4AHIAO1az0QTqDJQemqAVYTIuX44g2nn6bh01a4N3F1lz9
c70D/TpwgCyYE0UKMK36BLq/CuPSO2Az9BAENlCsml/QmeCvXSe1Bmv7iqqSxwrb
ngV9QgfPUEeBosWxGLlyEcZkyT04eWGmak02CPL5i/a8wod1/bJZdifvSiYfYCRu
tAN0U3tm7W7uDzQ+kRG1F9AcWynnq6FwtEq5L3WTDoa9Jxuga+VDECe/tAtmeacq
4/YkqkG3e9XH5IqExj+H97J6kB1+RSxQkqRCs8kWZu1HOoF38okyP24J71VZsw4g
2+BGGMV9qnZTmDZlU13TtYLLlVBpiTbxc/cPZ8PsP3R1u7Lx87rIUeDSQZrZFS4U
QsTA67G0gcRBiQySlAh8i1jQrXb328gdVC4c1wljFqLjANgKQO78LrB0u2A57cwh
2ob/wKTs8xLZEPR8VvrI32sX9gQKC2ddBJAPPS4Y5ehc3JnRhiU6i5oPM55nUkJL
SoYjfx1UYK/8Z/d1FA0zVXQsm5dBYx0MngEJZGD2q/gbD/T/B0MB4UJ8B0FoUCwi
fvJuo6iyLvEuuBes0k5RzVQCzSoYFemBiSgv640l/UwnOC84iyOk7DRCYx9H7aGV
SIHt+h7WwgwNqA+xDlXNlVwm2vZO18D7GOVA+wx9sZAl+OkhfDQaArRAtKSDS1t0
0EGWh1tUP8/9DrTqSNnjukU6kKprfw3A185mjN3+6F0ObUn+P3oDaF0MPsoMetkz
gUbgpdMol905UtthHglCWKHxhcbxr22dboj9jbTa/xBFr6uhKXjg3UO3FkAGSgzy
lTRcN5dYL3HNpp1yzZWjopRNMEsOIQZueLEB2EzrsXBn/IRiN0khX/xrk2H9JuIS
spOLoyiMcNmb4eQCVcyOlCb9hIq/bqy8IBAHx4+14XlCnjhBqb6tzOra01ku6U5K
0wj6LW5QYyV05NUOf27ARIP8r9rD5ZHWzBpJyD8vBoPPVZO5nPcn1iqzEC8OYdk2
oiGr0xVsk1AU3qFFI8boUVZjdim0jM2a6V/YYY82suiBJqWXJAzYFZTM6uwsklOk
PgJ2K70VUmDYLABFlDCcuWEXXrciziZfgcsD+sJ2QHj30e9Sc5J3WrctF5rhB9i8
i+KmvoO+q1ICqTk7HY1FmXUnXLvetsXA2oPdL9tcJNxfjLuc+M6QHy3L4EhWdnDS
3drgBWpwm7/1+tmw3u0reLzhqdWTgcdcAMh45bQ1mfa229/HtHpguafk4LByNkiT
4PxTvH9xM8NqQS/fdJhfBnoACx4vMeKk+6Bdwnk5VO0n6CLEktIGxN++vIUAYjkB
ncnKoOSQWxQkJ8WsFXtioeIp5aEAffdXrKIjDOftPuOmZzskI4i2Nsp8H/UgrjVb
XTI8FcSO18Pmxb0t356WckxwwQKYBvU7UbAhgFsrm8W+ude3LSEGhoFU6hdYEDqT
VAebexis6H5LzUTRxlQN9YhWi7S6G/2lwxwD24oG01m/ynldwX4fO/iYfxBM98Sk
vXIHikZld77Aqeltll7gByXc78o1pmy/sN4mwBkyGomWcklDVZJ6uPzT2KvGhW6U
6Njlx/8sz0laph3px4JRk3Y6FXLQ+PRbVoSeroPHXByGpIeGSJ5ErgvGXwRU2prB
CJlQak+Mj5Ni5sAVxIa1YZCeln+z9Plc5brIJPaNqhDsLGU4b3uiSfYflb+rDtb4
/PcHR8Xq1fdv3dMh56IdASslltrjbZ4fxSUF+uuwmg8/4Ao5D+g1BVd4jDLKZLtO
25JSK+a5/UKgevIpiOqSrMPt8rXTNUbzC1CaRx0CYG2zAHMBZDXoDAceXPC7+Y8f
g/VG0tC/v5mR0W/JVfpsui5houL92eZwfdMzywpDuysASYmWuVOkgdHAfemET8Mo
RBVtln/olawoi+X0Hw4DmFck8lCHWUuSo6gJtmv0x7TLUMFVxjR9MGx4n6KEY4TC
TcMrJyXmWt2qho8WuL8Tm7qzOm0ocrSqQxFyUq5NiImMrnD14htkeO93zUm6zZQc
TsvnZ4ShARsbYiHA4gSOCh9CLrJVf4GNrLE3h5wC8yFb2gOgfAm5rKpnJKqNn5uj
A2sZdkeUByfUqPgCu0vAzrxZ21KeVfjzCkbn8ij5bDVO2jANEJfIuDGQewirOt+w
6wgFn9eMpI/ON1mHfI7AAFEWrlSUejf5Ua++S/6TQjaTZIIYEclHu6aAmx6lfuH0
rjDi6T5ARV34AoXkvG4RLHl3g3L4Ks+iaNPwqibSYBF2My1jr/7NwstWjbvukfk5
C4jzpAzX9GfkbsplSoxWwWBTsNFjdB2osB4St0C5vysnM1Vy1Vlas4Cnnhmw4/+x
gRsG1VOAZXzwZhxLZ4vF7ngG7U7VqoXOBCM9pKH/78kc+jRaG/AnEuau7iukQs1e
DFGzndGFyYHc1VAM+fIOF037sFVrglsgUS9LzuFSQ87qqCkMkvcC4MNxPCHGpnST
T5pRVw0E02ahQiOeaaDCiDrosMAinP27mYBA6ANpolodKp2JtlIdFyvye1b7AY0Q
ksvQNTsGaKsyyPI4FYkOYoUP4gcnTEFwS/FS4yjsSmDb5XZfqS44zzavsjy99oa8
1iYXsxpqZx6fdlIVvI2bQPmp29H8kOPP0MXWO4EZJ2u3EFO+Corv8qTEJENBw6Dy
7pYqi8bvcBWm7yo3n2kIdmzpKua01SOPPBA/dkbL5SrjK1mpBOpL/WXUu/oSehhi
9XlfzAitqp1xUDnib8CyiM1RAWiatZmcKg3zyhTOKr0oMzKQUhefneyn+Jhh7GfJ
bVFDKnVj8TqzdZz2nvvyjVUzvVKWYwe9cyf8thuSOn8Dt/ZjrRRgEIY5yVF/88lh
Hq1mOv2TuvNjez58XYVVs5o140x/t+iDEWdErUSt+Q65mH5Ogn4QTHe2BAU1xV5U
VNxcDpUvhNdCgrdYtoErgvZl6JfV35oqtSJfRaC5aX6i4J0bootHKRESrsjQ9Pjy
6yiw2RBZiboXyO+aMEN8EB+MHdlMcAy6mNkNtKR2DePm1JncdTYesQIPbxONCfiI
z2hMEZ11tLAyyERPeEmfamI0hOjp+opSR2SUJG8rtWItLlR5/mbyuUKPKVEXnTC9
S5Fehgha/sKIZ/5KeAl/GqCJwQvEQB2AgQZzYt4E13/vC5PRSXXq6OqipXrQCVe3
/dYyIrvV0sOO43diiUNomwgjeVfCFENj1NQY3LOhycCt7MteMdyrvyFi9+vuw/CL
8zSWIKs3C0dB3eAfk2760Wgtnc4j0NdKNyjYjnaBYTLnrtY8O/bLPKcSAl8sNKTq
HmZsGPZpdmxgyii+YOiip8PobuvnyXqGYhljw8c56ilmlQG5hH23jPOEW4bw2H2h
yRUg4Thq+Ilr1FMnCcJMEd8OZrqwTL5HROYDvnFaOq5Yai6Y0cT6UXM9g+mo5CsO
YEvgHpkIm69C0RrR5NZO2UAWh4vJWpb/NSVPUYPA24wqIfjTjPvFu8Nl9QMdbKDm
SD3AhPUdQ4y29+VFpZOrus+1c8q6PnGCs9ql+dYDgDpL4jyQ7nIFBSClRHCX2+xH
mmdioZxMo0R51bGCNNbl+xJXdTAqHOwQCjkjBT2aFmnXiOZ5naiDBMy8NST25cFo
p8zSbVcbWVoXDSBlvDx+y7G0ikdgrf8sdfuOtmtMuWRtObqdatchaIK60iS8KAf3
5/0+H3/QzVnlg/lkkEBIzjeAW6ypEeiMmSIJhm7H6qY=
`protect end_protected