`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9776 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
DBGZtUPdvgnvgIFp6VMrQTmwpP23Dpd/8GUbBvKuYSfoODhtzR7MFjir4+eFmcFp
2/qtMmrVkD7Eve0two4Ol6+4GbSWjFWWGlUFcWtIAczpQKEaJ4jBjvoatK4FSyUj
wjl8KmAdZTl72tgkmhFw+PSnFs+XLgSK+5IYZxplx7OLsjiSB9V3QVhSo9txalLg
JpMhyuiC4cCevu8Nq24UBmWmyMu+3KlyHD1uodJnpydGhMXAos8rVyGMo8w19ZTS
2sP+mYlbeqO6bSQdNPGJrVEmljJ3qalzzp/zmmwyfCsSL/squyULauLrKJ7qjZw6
BC2anGMvWY539vccuOvUAbZ74kOP6Cj9zya2HTcEdv3qpDaAhUzIdCz6bUfjI1h9
h7WegKTHWDUlwZAfTig6pPQHAqdhcx2LEhtGRdgl1MJ99L3HMTA93Q+UlUILZx1y
PBWl6h4+jvQtnDJez8AtGBi5vLDwvVRy0uY5U/D13ZLmJIWEhH+ppfqp2Wrfno14
fM1SnqJUye1It8/J+GfdgYWTk4xlfH0E5sMF7+0b/aCqx++HJqMad4ruAFfrjpld
lZkqQNn9/J3R6L6KYgAxcdsBEoMrIGocUmmqELOhF89LtGW/+tCQ607dFCeSLhuq
GgUoAODe2HN52QaXO//zMZQjhHq7Vv1Vr8jUmSTl3Nxk3DRZgqN3W8K3UX9hyrkC
dEr4Dhs1KAmQAhx22C70qh937UM0SLQeOquRzJy5DumJPG662aOyjxsEIYHi9GS2
FAiPrf+JyI+qR+UZT8IEzLEspIiEM0h5xCRwqvex9OdRb/5JzE/wJdfu0jp9N/sD
5f7rJy3h/+BALOsd3Bhl5rM8LSuNGclufOvqYltkmkyrKbraySI/mLf8u1bdXL/E
wcMs4WAO+6GiSL00bpfUMZiJTxdoAN4DDXg6oG9uV2B7aMvUMt16mQHnCQ1dn/ZG
ZHKCbDW4o7pf7Hj+n/oiXkQS/9n9wWS8oN9usZcbmnT5PWM+34XyhRu4z11lPrhL
pbp48tCHKlEpmMneiGs43ced0lBzwnsQB+TgBrUNSQqJcbKx+g/cGZKtYUEQWZK5
scw5Z9ha50pMMu74J1+d13sWi2pLsJ+TEdylwD7DP1pLCahX0tFFLZ9b/RFQe/zd
5KGlaqJyz8Slp6en2M/WWbJYdV1qCWD8ZNHSZGBiaY3SECQjzwsRoBKRcoPo8xm8
DkyaIdvS32LObR5Y+vK5y6YS1Ed6v66XmxdHBvqcmk9SWUGYuoAACq965ND4gI5t
2DlFUwadq7Dt5O3ilQorhTaKqPQpbQo+wzgsS3robYaqelM3Uu9NN3TWt/8fSkIq
gpI0JuS1Qdd7eTK+19J/zBLi0taO+Kn20JspmL1TFXyIyqLPJytLSqrUp6XAhXwf
JlkBI2VQRM1phS4WY14IbxiFgCLMAm6QwzZhnKIhoGqyLgMAIAZX6P1ENYD8ElwU
odCSIN1UuCnnEr7BKKOKI8QItKTsIOjj6iVH0gutWEz6+LT7KxUpHib+Crgghhft
Vp+NM4G2L/lYCy+o/KWnpgFB3gQy0+m0Os27Cm1TlkcY4vVmfhG+wFBSTNN/Lw8r
2cjMHUffNfkBXULVrKxEOEvVnk7B/WCgaYk+UgXtMs+DaCNRG52SAGUBnAiMpfK/
iV7YblA9E8ZgrQlAy19jjnylQ4t9x7b1OG28TSyrJ7U+64QHtmvWeCD02xjo2ouC
YfyF4wLtBwICX1HZCOcw8WntPjG3Lf/pQqAYaBGIk9IBIAO+Mao5ZVDF8rxlxW8X
rYy5eUmxZLXy5yEHC/WcmafjIHVuZHM+phLtyk7aBKhfcCcggIin0x81qKJbz3Bh
AkQpv8m2BOrCaqSSdDhfeeywrZlxaDJwRpdViAh+IKVlF/PRda6kD+72h6Tz8GWL
WGRZ0GIcpBrG+qLpC/FaolSh8khdNDlqJ6f9RUxOVjOmuJZGjCi+cxor1AkdQBXE
4pECWeG+mPAL0nlcDGjJsCnzJBHktlFG2wznNWl4C8vZm7OWq499iEwYJ6dTBxd6
Jhed5YAxLpZs/NsgGFGf25IHTJcbpRI66ZceFdqASXO5XbTV2mq4JrITedwqpnPM
D5N9ca/CNu9Xd2Sd+ZtcHnw1NtCR+ix9xlI+NhqG/5YL0VTqqLsdwgAfcfbIxvw+
YN57x5v15M7XWl+AXafmxUdOkYF/45MdJNLx46S0xbcZa05U+xDeJH4ti7cDMVaW
0/wghs9KVcEtHqIoVXkxzW57kqPMVeXPo9yg4DEVsoD8EbkXb/yo9fMmwd9rmFyu
7wpYXW8G0suMGTSGfX0FzuLqCtWXd8HtBfnWIoGiNNyntc+y2FjTkNDjHHj1ByH3
CtQtb3AJXfLqO5B8gGG9hegemX4DdD2ROslGhfVGNJOHP1PPp+L9B3Rcin1+vXgR
rwDYUPBeogFrhoru4H0fyL6Ln09QyRyHWw5Dg9leI3tas2JedQ3FrBTFxpgxpQtH
+vX+GVYOD9zZR7lDOuEniouU0HR9fTLhqMEUgtcAMuMmqj8F4iXKQlWa8trYC0+R
WYiGxtJ5l1a1ZDWnhg6YlAOfNLbtwOPpSkyYLkWIvb6Qgg2hA/M0iqYoRBEdyGL5
bzf4qKcmn2Qs7aQnOczcHVZgfzB1bTODNn7MdcenJFXztfz3yPEGN08N5kOpiM1S
Aaxd+Wl1e6ET6kiEnw2RE4CFQkNOYFuSAVaofAjweRO3WBDCk7f4aQY1SsWjVDhe
C86Q0O9A1HCEXPYMaceBBheF303qlILJLsRgEEAPofWLCkppl6P54eletLcU7PLA
EZVK/c3CSmR0vZAKcyYPVHNPR4D4r/eDBYkROChRQvy9ubxc9mfyyWaYG7SxjeGY
eDKoFAqIL8Q/b7WiRSUw8m1H825exbrag6ZLKCTdJESB9Hf3CQnogg30+XNJBLYA
kKo2IdVcT5ygthAnpIA/MC63VQcH7LZUXLiPTlDiNiWDXSh4y/2woDfmoEovgz7X
GHqtUz3ueEhKR+UckC+teIgG3rtVRLB+jp6QBsGxdjy2jHJ/Ztj7T06UQhMSjIaA
e9wmkc9RDQdhDRpqrCJhH/o+8D724XqGiJktxka11TveDEzCJrLQGdyjkMeAZ+Wa
MxrWOTV7nRJ5ZF+co2nmhrF5lAth0cY+9wYl2pyCfmUNIf5XkLZQ5FR1UNtwGrlU
7UGs7V1NHxYX3jJ/1UgmZzIlegWRDgyzO7Sx5oks69Ufy5L9acOaxoZhYKaFlGe6
/srRDrz0oGSbY49DauUOAW+a+eDFWYo6aQznUOPGpkn0rRVFfveP/iS14KXrB8Mn
7SKy7f1hPIWVhYokEbA7DmBAgg3TLhhkkSITnYYDZgkRMZjBFcJdeo+wPEhd2LHH
RjgqTbe1Sn9sY1cHn3MWL9Xh9i5N/FB0n2HbjGQmyYMGvt1pubNeseUr1pCU8dWz
Wv3jsZUFm6T1p/8gwHNIh9Yikh6Ar8H3cSdKJ9X7DofVmE1/2uf+yurorgOpg42N
eY3DHd+ogioFqj5jZdh1YN27edAKjhRTYESNSpbWjhvqstGFMZfhdhKAJ8whuPCJ
I2SnKYkdghEVSnF2WZjC5tIaSWvMHDA0Slx532uFaSY1i6ZWgOPpBbKKwA5syrCW
qrOnABOF7C0FQFNQyQgtQI/d+MV8b6FQqNwBwDtjJVDTh54CP0I7l3a0HHuI29s/
MY1V/ijaO2SM+t3i54S7IdVlSPSUhYOJ9BfUuxu/ctsfSeOG1C2bQwj9PfLDlATc
bZlBKrveatNUV9xxxVClUaxKxduX7H8FqbZtW040Jz6Us8kQjCx3V7xNlibUSPQd
mZHDnQ/w5CrJ7+ChYaEVa0DP7XDAdimH5k46aHBMo8HGPalu/3PWjT/u3pnB4+gJ
sxpNDT3JrfU9YKJcMGMWtHSbi1vNhM21oyFtIo8q4Z3PGimOu0H/Q5Lmh8SytsZV
fqNsO9rHR8YTX9qSzXx7xjQYKDvBsQ9UnmbC+bTDZFS5vpJNL8LCl5U40MCjCB35
ZHP1oGF3T8yhZffMNE0UXQmCWz+fiKMbCf4Za37teqAkZYXF5XpsuqK4cz9JiTom
WN8MGgKXZTMUBc1QmQBt8gCzqrki+GhWFpypVWIAu9HWbMytjzkWEc7r88Bu7sTg
WGdgN5LmW+3B2+09jRq3Gol7Z4I0zQi8qaDBuotS/zSO96G0KyZJch/1UqVJn4L/
4LX3dWWR9Fm5vFEHSa+q9e/mMK1e2R0ZyL0LQoECUNboeqPVxb+wYhbfYtZy2K7M
yGh2YdPQYowcHjmJ4vshO4lHUpokBDd+7i1KKVUtodopNPJjxmYdEIa+QRZY16r/
MWnR29EujrwRwx9WB75dOOzvgDeccozJeog33XF5TuIcusozWTqNxOxdvG4L6eD9
bj6wsScojZI42nur7ghKmm4Vz6rzPcPsyuXVHZgfu0iUs/VBPE+uglvmAsAVRM3a
JNIz9ewBfW6VQ8CnOexEZXkaZnIXKdbnpRSuc+AfZXn9DOTYiquVtZA0KpH53MVW
wYxZV44F39L5T+Wg0QkJ9mEEOdF4jqOze+SuwIjPOMtb2vPgJwdVZDtQFYVAeRBS
tBIUjfRjb8BD4/G93bcVLS0oflngvqEXVtOOMtU2LUZVWkSWLywjpnKmIFU48Iv9
lA/JK+ROkfyPEfaOepFlfCE9j8+eVLxlzBSRPAQzSPyfRppk/s0119+7FEGF3D7I
ByO5Urn4hJzUylGJHp0apUmT1XOk1EoqhSvXZbFtd9Vu9FdVBohnBdNwRCUxEtn6
W7WYqCxEr/WbgA/vHJOd08COPno1d6WyCAps3ZlnE14KFFHs0uhZOiyr+Yy7wHST
F5jC02RCOYH/qo68WeDfNibT3VeTtL8gXAD2onVm4duuFAmtX9Sj9ZVTEoYEmAac
WJ6kNbzBgt95G1aHDyK7P3GNNQ3Z5hxTdyXElRqgL7P0FKsHl8xexgUseGBH+1jv
5gnop4QxxTO2Ok5bSZCxOCZeuhPGsLfolZLZbLRFIxylWZYedodI5wur7lzChLaz
b7ArZ07cK+wKJPsMgyTrksV7Q3SiLLPWSoS7nIKViPAIJAolEHmZsLJcab2MpDtR
wekiB3eTcpabfNSmj7MReSvhJiDp30kRGVJCQFfHU/bY8YWnQEjbE3ei82TN5DrJ
mP+HHU1dB/0fvAEj5+lG/av8/fryRtbngzopofkf/sFP1fOB9RHTL4fB9tQJ3PqT
jFVZEhUUFN5jYd0RrhD4d2/Ak1P240qYq9K5BsC6mjd5RBvppIpm7Wxg4rhGZ0PW
2xrDQvFp3a1Xq780XF1zN9CZrzMuZkP2JH71C4qHqMqw5UDwVbsWZPoWRwZLAdZz
5HtQmS4zsgEk7XUd9Oqp+qTd1jvQGMUwLT5bHXvATJV6mXOHAp80RY97GjLrPlLn
m1EaJz+iDiNW2ps2KcrKHcu1I3N1vj49rP+3ISSJ1ozPbRxmOvHOAFPYDBGU+jik
1E6sSdjQAuHzLZpuM49G49CdUPBDEWFyJWEcDaBDeN1C3ouJfUvFdU1CFu8NcgQJ
Ppr3RcdD8ASmL3YBDzIrdvfWCGjnuU7dKXGfgPAOD4ntqoBSca//tCgnp4nlECoO
Hv58s2BelWVLA66NsR5S7oEtYgYK25lBcugl757X/DIAoBxU7t9ERc+SGMGuY8Y7
nmx+U6iQ6t/mllwBlejGvsx5XP7CBq4PkHQzmLa4ta7FPhSadUFPKW2G0rAZr3Xp
AbVSzmaSDiuHs3fZb9UhUl9l7YrJoagE916GpBctNc+EF3O05LWDyVOQA9GslKbA
IzLzc6Bu23JEDNw3C2uJ3OxN0HopqCWPYTrQiTxfJCpgKy+Vu++9KSlrF/eI35RA
aYtL45ObZxYABiDNuhFnnX5CX4Xn9Vyv2tx9DZssOIpXnQgyFp1+hmrY3pQxU9IX
FZYlFTwIt3Qt4WAbfpipeNqTVUbJSW7tusFrl6QFNQ6cY9Pty0KoVOuVQbeeZ978
0SvY4RDMsVSRn9r8ISWCPRGBr6Ta8TrrFdnl8GSz31JAHJBOu0QUzZecrm4OE14g
MgEfWzw90NfP79di+rMVDRTizbTL1SqHbYGtc/DBaNU/j3Zo8jy9wPV5Isruacjf
uQKqPuoYRFnaZC3J1eVgYK1pNqQ4QwMtdv28v/amVQuxWwAqh9Sb4szMt70KdKYf
+2yTLpn7o9rd9N10LQaVx1zPylTj07R9TYr0v5Kx9ldzJRaUKvEidYnWKqXYr46b
gy87Fz5z/HRCGg1xsZgmvQ3aLmx4RyycfoJ3qjAbewO+lbnG3/JDXz4bwLxaahdl
cYz/7eESefh0a6b26DuZlaQbblsMP00OuqzDddPbfku5WfOmH9A+Yaz+rFPIDdF0
GYORy9k8ihaWcCu9yRrEYuAGwbXLAGBUcxVoyPIdj38AnACxkvANtLFX9OXYidHI
f6XvxeEGn7glKTw4kNdTQm/CxAjlZ9TeFIn4HHSd9z3wq4R+ZnSj22UKoHAn6EFb
ZyESVNMizdpXWHeaJ85RbM5hoFqB8lsn6UHEO4fTDtg9QOV0re3aBje8bioNPZfj
DxHDWEEa4n3PM98S/4kdCADAYCgPdeoLMV2apmwxuRjKM0+gs2xB001EsxHXVAvS
eGrkcQGa4tFm/8P+iSkwPKTGZQyVgGWv9KJuxRxY9BjDOb0+ZafYeFWupAW45OFt
hZwb+jpR7diKHcVEmpUFK6x7FX6HSIUo0WyREdqw4KIJmtZIObMpMDQcK4VwAxVx
fDJztj7TkTF9xATNqTpGgxqIyMV1MSL9juizwywYe0LobQfEF/qm9qQ0laAsiW3E
FG163Q4rqP5Luqq3ao5COtnJoFqGDGA+VojXlzuWQswN46SlM7FR3WxOfK1jnGwk
Y+t4RPXN639Lf2kkK3jeQekFprvFXTVZiEZjcKEw32rU8POsbN1mj+m1NFcaudyT
tp9ZOuuczSPPfjcNFKDGJf9U36hYO40p6qbfCR8gNAZmVPo/iSmozegXBTKJ+ngJ
q6zuiGvCoRjpZREV9PJ2cNjKSGwnqKBcC5YeoxbEeHIyf2h/yqIG9NFZt2YlqQY0
C0ctBoj5MCyjJk4LzapFx/C2xwtIJE6/mv8isQ0FE11YDExRjs/YisOT+G9gOO1H
kFQ8wWVk0Xn0eIHuUIhvMxtb/VyOnOP4iZPOKGtAF+og9Arhi5c8QHBqbPXUB3eS
lLlPGZdKRlan/8mprcUQWVMqttKcERugOX/Ar/6C/nlACam8ROUGWQWY+UNGT9p+
aHuGmajqHGPXOn1vLU/4tx8IMvRSgx+F1sz7vvbZiSJsiubo1Zm182QFjJSoXIrd
ZkLdYFmupcVTRaBKRsAvztsY0qtI/DE8bkaTMKo6iXP93yu1LRKnZ62jhJ7LuWwG
6DqpIAxD430bFzUeU+L33uX3v0f6jOB+69UcLgdzMuh3wkGp/3KDK6E3TZGXih21
JDX2iEyBgebqFXNTXHkT9l81rtb4wkdHf0xMjedcw5UEcQFQuWtB1y2NJ8fxaVW4
VgCKjoYZ84ogXwrBzPg4a/MR0CIDKwuQg9Km+DQhXKnxNVa9FZYHDoz8iML5hvBf
aGUb/U3lyd+zEVPWc5uRrydOwU7kA540k6L7Ba30a+mLrOpAem6WEKh7eXCQM1HG
gdU9u59CKQ2kFtNXcaLCQ5kwaw2bdjajdt3yZIYbFfx/eMM0us8fgmxGSNatEPd7
1WQd8EvmMI3qRuUZm6PR+lcV+QHDhLrZXiCpBv5CLTUVQdr4Tl7ndWj1lSCenY1P
iyhOhS5p5KUB+Jl7uIOYb8sF2KsXmLg2F/+7vLqebCRJedE/jpNSYPnhhnuGw1vP
IQLgZY79K2QcNgQZrN1mpCqRqEegPpAyj7Vl4A2duGQohdhoY3nGYGS0w1bmBG0f
p036g0S9LvVbeEkQk/uH/XyHaTUii7AZtYUZLbSfrcQLnFdXchKJZU7uTGQ7XdGB
KBv5nxL4M5j0YyP6LlhhT1gDYgFWn6nf1Jup9YyIGh3Dvxs4OxgqkK9ecRmIDnAt
va0ys25l8rcNHzmilL7Jhh9TX9/JNi11+/Ad9C4/hMdL/YKxmULToWLhmSC0wzth
mzcb0Tqn2EobFIZAa09TMameqyypZ4XoV7tEG8fPxzglFzfuPVmcF4NnLAYnWMso
2NSoXxaV6zbbKfN6h9M7cWwoQfbcPlR3POsSuyPp2Nyo30DZ9skGn8/E9dzZ4ozw
bHVam7VAkkCCze6qFknpAaxAfRHgfMXGHkDR5x1II460SOvUo/wb1UEzOkB5P5Sb
1V4JxFOR6l3m0y9GjmX2gTxLIX7ooDvqhFW4sqQtpUlpa4dp2IKEZdzdauSSnI19
daDv8U6GPk9gA8TLb3CHkYrRXf89HKfL6NrdSr3rjEMdi654gKgsZiz3f4EQHX3v
SvoHxbenhY+csKjIGqH5G398/onp/GQlddZhyiNysq0L4dCdhqqXNbJ9daWXKSjr
dOx9EJJ0pwDvNwY3DagQWiJRxNEQUjVLIWV37+EfsQf2+YtB3p2wDIr8YUIxx1Kz
DWXJECywZRlsNLIC5X4DN4pR+k7pirnvab+elENcVCCg+mVbAbx+lJiWOlI+ZUyP
cJSGKsYNd7i69tBgXfpS3J2Qn4npkaSoYBQ/37wTVVZAXgSxpdh4WDPcAOuIeQ7j
sEKsKTFVUXkt7R8PRNWSdVz1rkxBIw1KtHHof7Ca7mVjTX/JIKY3KMh87V/9JMY1
eCJnQgsb4SPHdjJRmv7hWPltt1/8WWb3D/sWEEAT3JZgO8rzGarEDe+Mj4LUX9HF
r8rJjMvJYbHXWlaMyaDqWtC8l05H9n9rGnDixa0VDwAvYHbuzfpH1p392IH7hkqg
wNBLDczdgB86GBfX98o9661qXoqyC5fMknKAxNP5co8Y0jnQ+ndOIUCLoFtSE6j0
O1mPAl2MTc9VOnkF4hhCGjIv5fPEbPcx/P1gfKTnGHlu5jByynQtHeOm5+80Ll6l
1ng9qZQo+zp+1hDzobfdilLuUeE/hUuUzUnxhahoSZDRngF2nZBPCKmuM4X0Pj9A
KA7528+Wp/q/Np1ClHUsuawFo8+b7Lt9DQ19eHIk4SQbZWNaVxB4KhgKXV/HITGu
+1RW3fohqmexniiX/KJqImMrXEY4cMrWYTPOct6QZZVOshLZA/2u/oMd6rw8Qhqg
B2ugkFhkHMRqo8fTODvoqpyE42qJFvRNd8+syEn1zkDHDbWJGOTZzCSimRWoU7iH
GtDE7H30Tm5vzbYgm+4SPRKvD+/yFMccuei573lcbbqtPI24MJghJfUqAZYC8OdL
4p66K0T5Ea/q548IhcYNGBLEMXG42E3KNZHzcKJI+ggVA2R4gvLv6L7TZxDv77WM
Jp5ksgwVlPw9U09pi1sYWP5bkSM+K0rDyfZ5W6Gm9I4i97p8GoKyLkuG4LpaZzgW
KudkaqrP5HkgRodceKPAcYvcz6v7RMsON/WfZlzH+EsTBft3ey5nOsZbrYXBFNYC
Rrg2eeaUyiQ/Ho/Mwr10tenhLvGGeQX+i0kAE2uzZCpZUeN4H2JnZgSC5EQqgmXw
mIYIYSzvdFYsV6CHQsLJcq9jPehgFiXvNHYlC0Hi6y3AazrwLUyQZgOsFPVuFm7U
1pvCWu8Il+m4WrQ2BIgrTYHNc1ucK0XItXsE0WNimKXiSsnFCHrIEn57zz17y0Et
sTnD6mhNNA27pkGq+NZw6cSlOwCA1OUZQFx2NWjh4YTkM2ilfoDQFCKlGRFTV2iQ
i+PijerlZXfbuIxbGHwxXhr/WiKKvnJ19cOUe+W+YmodWshy1IhxMZg/JGdUyj6q
y2yu7RPh31B04EZ3BF/hs4fEz98gVgHMRACks5Xt/3Z1yU/Zu782TqZtLWvU8XNY
Pyvps6Im2g/dAXuIZ8XkMA8llBYKK93sAP8WRCOJQ0XcLdpQgqBcpKTcSMU0hkr3
quv69wrD6X4oqnZwhEYn+MezqG7ug4U9lh6zR0AbI0WxEJzS0ORxbURyikzMuGAW
WGRz0uSqxu4C4MEuJyuT6mgmIsHIRU56ltSVLzW+yfbMIhUi9rvaoweuHy6CaDU5
J58rZkdzubaDNM+gfYdylEQZFi15BDhi0LKAhPcm4NCJ5uJGAhe0RQnzqmvAgb8z
evYt++S16RY7vdjaNDKJaaqOF2Ym5egdXh7sHZF+Czpv85vEkDk32FbAobOd39ZZ
oyDrhGeJu0JUHb5tW6dJUP/jZeTuCSGZG8ATp4cE5CFFFCUshORnpemfTsSw0yYu
LI5EtyaB3H7TokAAUgYYJUvdws1IKojpUfvypb+hhrds7dLHW5jE9Sn/jacEUTC6
B0FwN2E/RqY7FeA9wTRs2fbjczLDQa3V2aHqdLZ/XgndiGhw96b+UqciGjX/n635
eAUsNwH0w3CmkZJWACs5oIdXipb1CDRfmHhi+z2KTsE+61oVgoN2KFR1z91Lbrkz
hwAusHhEm5ArqhcJFfeW/bBzWFUtujIvnMU2kFLF8NwmRtAIMcu9xX+/MLrW3h3M
gTNeqrVZtw71rysNnIDXPy6EqY8bKP7JRNEvXtizVLvsmfTkOf+QCfgBLYHH1IC6
UMdlDX3ZjdJIxZvmyFru8u5cTqlflpo2tzjYjqBFgMhqbtZrkZzhQzk8VbhDPyEG
C8NZ8pe1WPsG6MkprxQx6yLZNeeNyxN3o5yihG5s8ja1Ss+DWEzA5SC+XJKoNe9u
mMfWK3gmoJNUgk5p+tzmQRzPYVWibUHFMOQAjgrh75KGGecpDV/eC4CfBVZLa4kJ
6VSXqwP31NYeVr5uv2sqPgjyqbuGNm4W/WcfN5TU7ScAWwywijwN/pj7S7SrWLNp
hYKFC6dWrn6sun8WNDl1zMarTgyYl3Kt5r3Pb8khWvV1WuuQvsZlgzAosz4NUS14
pRnX5DPGVuMlfZqMCMo+sSyzcoEHu8nDkbsbxfHaR7EFapP5+SS4CtlbNlKJGW04
AQNIpWPKcC4AzMrbikvyJw6RtBIoNEaMJJ6n/2tJvO7k+Idf9a9hFEr2+SqTKirP
zbJ9Gvd5WrKgBEqXfrl1F4LH6Tw5D4HjWRglneOzH4SO1tvs9TlWUIE/ZF9jUb8t
B75PCJCiewr6A2l7JOru1UVSWJsD7KiW/JvCH78j+7onX9wqwFGlyvBpPdQL0buc
HZsmuxZKa8SFWH5Yv5NnrpriVqGYue+HoQIgw4d14v5NN1aDFRBpnKNg36JODVPg
ixvhey/7rp3rMXhQtYOSSMPqorjKeZLOwNs905zJAULydm7L3KexSkyztEcn/q70
hO/2f7JqDUjYSjNialYI2OhHnnIzQmifCUb2VG5gl+gMMYn+7/Xo9r+9md9cmblN
FOxS5AYziHHAxvYiLDTKK0Zg4F/IfNA1RxRjASTn7PKpur/d5kSa6y00VZuWNela
CQIEKa01hz9+CjvRaVl13ZxTpCWFnpqKmSw41+YwH4N32fK4oFLIXnaVJ/4LBc9Z
3BiOwDAiNOY8nJmbNWEJzyxnUvoJFhAMW59VqZjnvJ2EaOGggxMVql2TVZVJoLDZ
Zmi587vx6+3gF7oSBbFEP/y6oHtUR+eYOa6VkOSP388QWPj6KKubL+VzZaSt75+d
v2XxdLN0u0naoU/4N8axXm211/0+6Hqq6FLjVSOzEuo71+GpV92BRcCZK+OnHYmH
G2xpXU0c+M5ztOBWHSsopWm0BIapmCVAb9p+UccHKsgWfzUhpXpmoAQW6Ot6OLzU
quwJ0VxvkD/dqTc5Huh23gGSOzX2lrU+0sjkdI2Rb9CWl0o8EucI9MXL90dJyzDd
xsPsVd0/q2Xqc4+hL7kyF4OkTNS1/+BTXFKv5qhACN/VDuwzq4Nx2HJa52PETpIg
0qeCb6AcDMr3sLFT6ygf29GXxnhoParmYphR+rXt3w/6siLTT1dkVsQnQq35vn3r
lY4nlAKunPtQ8tNHtibQI/4b63tqPTtn2tLPJnrlwTIgl1VJGMul0bGNQT7p1xfo
jPE94s5uiLEXbjqqImeIIo7PKM8fg4mUHhe1UGDbK4f1rGEGseJqRCeohDbJWWzU
I8JWv4/p150Rq1qzkqV7hbtvKoGGI678YcBab7es+pb4nSQEAkXx00J867xTuBt4
ewYlIRKL2mfiDfadambOyHEsvSDUwWm7mY1+ydc3idRceFHB0fRqBmeO3YvDtup7
zTEMSmNYCXlOhr28zYnUxxJbC8vuaGv7hXn0pio+n4NM+ydR2J4iNfC9zVUqVnPt
Mk5A43gPyIr2R/Obi0buFZOM7NgXAV64Zvu/TG5WyoXUaOcteUhZuJ7pt9SpNTaF
LWGp97Fsvpw4hdeX9DmSzBTCgjobV5FMSi3efLBc3hZC7Cz9pqa0G0yk1HuOib5y
hNn9MfdJpmHvK7DbR+ig4K/EGu0yqe1OqlNPJnNo6gQQEpc7B1jAjnu+qg2lupRH
2RLgeC5vR1TS9oDJ6zNFBALYaX1LQMVfFYvnBiyCgTtMW7LnblRnrrTdgxCW+qxq
gawImZmRAbB250J2QexvS8kKJp4DCpbD4olmOk01AeIhCB+FgUr6i4dO0IfRSZNy
lKYLchqu+lA5GQJvhQpkMDd1sYCXkE9FEiUQg9V0bs5XuBJO1uoYmclrc0ALH1mh
umoB5WOrTTV3HuppbrYblO9/Ae/0zCX6QIy1S4wn8/GdGRzM2P5lgMjkqNZy+yO4
xpGAp9w9Tnpd9G3/RHDNtOzz2do4d1bn34+pbBudBcFDFvOLBNKrgGjY0q/IBp9M
JGR+wcEucBWDcKIA0xZvodHvCqnnhpYKjz7YWsLze/Z/NQT1lR3fS6gacleXv//R
FuTnULhRkvfKiSlJjXL3ikaj+FAQXlwIrD4oDMp+wg0=
`protect end_protected