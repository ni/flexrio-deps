`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5408 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
K21MooLiMCXVPibvGUiGAbbetOgCWNgyOx/O8Ots+fGxt1suzWi6MSBpRA2atToe
iTBp6ZKb2YZ8jble5ljz/sW+Df+iP0D3MyIK8ELB9gdxjEoTutfgzWIBDmCZIauj
eNo0abMl4dPVVGDPJ3Lo7SllECAKQOt5QFBepGrKpoO1jgoqZs4m5WiWP3W+Cjwc
bSYjIgRGpESpt5ZxyzX3PhcVmwyuElhMAYjUTEqgya9/hWatQHkHSxbiaCbuv9Ye
VwFb8K2S+k1gUvRlGhix0qflsroYhXXpS7JbnZFMU8Ea8BWsg1EGB2VXjFUKWEsq
jVYgO73UjqCsHd1bdJdgYkCLK5wx07bf+5bBFDgMHz6Q6D+DIn7AAW8d6JLRfgZt
9oeojCB+lbqMGrpvWAgiWJrwPFSA+nJIxIOfZVDaGjydWAgnk9/BIiQOQNRzIYxh
l+noCkKHqm6qVztYskFyXa5pPA9vXB6abX6l85LYkFoxG8Q7A6G1yjkFnomQMeLi
qBk1lIKb7Q2ork5Zk+n6WrtsdclhRfu1te3i6fEgCDlXvWtq64jqCERY8t3cDGKL
bMX2fkSENYrcKWdSZf6KWpZXQTT1SrafAfx/5nskeWl4GYSqiWuPXI2I/D+01b2h
kowsfCj5vb/32Jm+ewdayA9fvoEdf3YGQtl3AmO0DxhDXHbkMyZZFMeri/nxiQAI
ezOFyV7mp7cWDmVVVb/3xPtbIZxKXHqMXSq6Tyo11/EFLaWxNxSGX7a6BOjaZFgb
LkLFNkeWQsqkrH3T3MrHUaYnakOorw5pHQc6RWGw7nlm2XbxJ7Jl0EtlhPbskETK
nCiIhZPJWGawLYOLSJHDTqZPCUimpJw4+EQycnK6j1HQWLkCZ2Lxn6/Sb4+2X5Xo
0pmlV7M9m/PbqNuNS+DuUzk4wQZYjz/gU/nBMzIFlGh6aJCCz35VXgY83qk6b1v7
dBL4ZRK5V2KSWS9z8bNzDlpSHlBD+MPsVnClqS1GvQIu5rh4RtUeXNaktVPOqIFJ
p1pWSnN0XDIxXw9rpjw9T39tO6WgmT4YOdOYms1sNcritaVGcyYMyK2k1W6jDS6p
TsZPmTjs6fGnX3vnwxmlowFsci16Z4f+MDt4w/qLbZpy7JGg+Sc03CLC4+Ipl1T1
bsIgJ1e4YfZ1KogPJuS5HkKYD+cLYuiehgHfZepkGZ8jJy/g58WW3atU8ylx51YY
oo9yQ1YF1qoSIRhfkq+JoCFIdUCcmdPTvVgQcsG0ooArz8VH4xxaAizs5vWkcQPn
IM2gRzK12gbW+QM2GkEDdXCaHb3sixjgoKrrSJzsh1hr9dsz/p/zUmY1hNV40sYv
ztOcuCEwvnNmDZ9eoRE2DJDVqCJppOAzI++8yLF6fKEOxFElSgpc7CsbEzlatvPP
6zTJW8UXK20HoYQqE8MeSXNaxel0z6aBrU1rzjpWNxt9OgiHbR4yO4Foz4/Crz+2
UdKZn/Y+qfSqoodMJInDecbJtjs3qb9txasym9MJuzrSZDZrzWxMt5OHzDjF4ZS8
aVFvurMEaD2AiIk1ld3GmBJJ4yTlckfR/Spx0yG8z7oGUDYDvSFwNGB9j0OglJaA
uDBsvFXet/Kn4GJ5tNId2PL9OFVtJDR6L9pDX3uH+0dKGT04Z1/iBQPPbfYyNZIK
JTI+Q9dEtAgzAiVoMi0ODu5lu8HdIp/UBKna0wcnZ3/naIT66DYs3+Q9Mr+mFbd7
LCUG5pFJkxfn0BoFM5k8pqhDI0MGP/F9fqRHoVCksYNXPvWkTfHDjGPOU/5Eaiec
NneiryKPrS9sFkweVn3BIcbWWkfvu5SivGy5ASqvI1CwLZaagEdPe/7AWUvw7Aih
JZ9m57eUezLc4Iuwy88rIvtS7GauqoU6HLfxV0riMHHD9WIqHBE/u+W+j+O4QmsC
rjkotdc71KLtqRd+OR+bq87kpR4ln1IkNRt036NUbzHpxAK4a1vlEcADFIyMh+LZ
K6D+mw3sxkrP33wfAtvG+25fCrzg2Cf+1ZiOgurHuXjPl6vVZz/srXq6X0DlP82k
7lRmx+df3/jmv1siTCXIeQJJuV3RtX+CqqqylBXCP6ac85JpTYwHnT8+FKD9A560
7OYx/r+OnsmwlxbR6Y2u3gVRtERBqQWMDZyq9UYU3yYewgA2yjynyvr1OvB8gvJ5
4f1R5XNij7EqeqC6tefH2X2sygldYYq0uYzs0GdyJVnHNboX+xwEaF1cCXvkMTYz
HmIpk0ngTkmHX88GZpinzLEngIx8aU69xEi+KlxfBmY+3M6qxfueEyPehTJeXaZn
Y2/ltMVBXyKpBsXOK10m+3bdvVm/wLT+YZTys9fr111TE26wmGtD+Mjg4IHuPzEa
N5ZOSD8tdPVCGjE3aXYJVbi1lxQqjYjG8tOChQ6GHRchdu5IarJN8blm4C7bc825
1xyP0zTO/gNgXKV/tXEFScFe58hgqbViSTL+cmWOpTofyDwyaJAXWGGCvhXgf5ND
Fe9HOfKjI9kqcOYz9U8/LwQ2FPMUYNv6JaQvxiXB9f7qAL2DdV85k9T6jkZhiHEo
4/ZP0hr10BDZaezppQYCNSzfxKuG1NyOngKC4MFqAZZEcAEtWpJ/orFU40us4GT0
CmT0S6dh1LbUQsFFB7nbLEBInG38ABsT2IGc0tWEb5qOpqL2mgR9rZ3+heMRlcer
QC1u/lZ6Uh+FRa4zIPzC0PPNtX1FPQh12kTfOSlfRtYZbMxrlGv1woWLiTOk0RYL
qkrqkqSHRJO+pKG26/ttXb21S69FhfBTl+02XzSQNF8vtReQ57vncyBt54t15K1a
g/V+Npqs55fz/U4Q/W5aCl9krwSWWg/vW9QumCJNwzUiLoM4KxwpZFsO1vwhlVfr
I/oA9eumy2OZpqqzEf3T4b4fkjhQt2oXNz02nmVyqxNbNjaXzZOHZzSR7b8xUZ9b
drCpaAUswx4qGQQRgUF6/+Ul6U6Ag0I0qt36Ce7/viXi+Py1erC7AFfScabl57I1
ae7dF048ySut3HjaEE8/uSHhTc+RGA93E2cwtDFGhw/hMED+mEiMLacyMMV/U49y
OLI2x9LyJadJzRonZWPXO4azYmmq53EWAQMeubnYkoRjTqki6abu5xGfuj8Tuy2r
NBY1nJH+vjloRHqQneLecj9U5y0TTG78pAVc0ja1j9qCHw/6GcDHTxhEp2Vt5jgE
A3O01Bv/N5wLVjTgSdbYlotelg65fDNwV/j7QB+jSsxRMk1JA66yNUItS2tzzjC4
lNWnlHiNcFuV6t7JDXpqMbUK+90YMwbIj+PWgT/eOoKYEEqCvc+pHUDtv//pRWL5
/+uv+umo1OCFrY6qd4YvnPxv/uPOaIV1209W+qZ6m37U+9n7ADjF03exJB5qyhYj
6Qk8ET8K9EZGlN8Hot42u4FMVFqe+SmLWppl92DqIxx0HJ8IrrhPCvb3T8bUF8pn
G1My/7VpK9XRTx4xNCTaBJJEBDc/mugV+WNHqjWdetrnXGl7Om/ykDetkME+qaVC
CmtzSKoLDx+FfV34sVBD6B1pl9r2JcCJJw95CUEO3zmHbwHs/oyuhFJ4m6dd7BZe
6xJ2o50UDpp4t6X8uDEmYyhxCxUIzmQD1FiMPYXeIjdtOAOqRMwJQr+fVvvSo9eU
9dBFvGP9TQZrj5P6L9TwoEd6V0pU0QE7H5P/cNr7pc2CFu3EEjAdkeC7LWil8wlt
JDeK3/Gv08GwjXtpxI/4tCktCW8bLUV+HpIpF3Zbt+igtG0NWSpf9dLhfgerBqB+
vTG/882bXBpB82s/FfvNGfD9g5S8Z3O+HOCNIRLo/YgGJuUvRfGT34ViHDfuUr6c
ZQ84TzCFJysL/0lwWNcr6BFgG2MI3MvrqS7y69ZFUhArQDv6xZK6X/2N3ek6+Vjv
UZpgc1pe9xFN/uwh5t7VtE6siBu3jY77qm5Ue+ejfY8t5cJRzFpUwil7fe7PTPk+
34oDMkSNAwvguGweR6Xo1FDR/iaDC4h4160YqOAVYbBufGm5MBEEuolmcWOh5pTg
+G7q2E+3WF6lpXvg26wU0S8oIF+N0JaHSgJuFRZepx9Oswrokiz5CZ8IjyDhx1FD
DtpB2Dtlb9GJFPUwq7s05465bvN2CBej+b9FpgU0l2I9LFHBvPhr0iOKK/sUEiEd
ftR9BuwxiYLOqe6MP0YToe/tQNbsIDD9VEr229PjhbTT4HnF+RlRByoh48BIBmuE
ejaI7xvGuxqIEywEV+7e6KUimhtFO22NGaKFFm16mc3/rIYYRkimo56+MmTGf/Xr
JaMGsyoZlkwUAr31wzbNgKwocZ1YCTfWhVccb/khpzJVRP62QcX3QFgGwjBeFgni
OjEYpA+6pfh6cPWQ7VYneLNJC8dtfJoQA4Fq2+U84ilC0uH2bti6ACmVfa3ziyaC
+0J/lqR4xNRT9NA7s6WosZl2blXzGXw+exPjfjz/jb+gpVcom3wsz4uPCzNC36Au
WNDqjmp1w+RAZahCVAOwMnZD/aJW7Rk/BZ+aLmwJMyZGx1e6rdeRa727upKbHUm/
Jfkrf1RpQ8RbG5k73rJ4KuHX+Tvm0B/YfGjpQx82liw02PhRIO1TluO5QshYCmui
bF19HnWFOiprgTcEGJHuE21BZNKVQSTugGYhtS5U+jlMrWyX8KRgclO694Xc5TC8
mu1HuPRerM+B26LR09Rw2esGae0C7mae/RenFxP1rPGSlrtT3xIk/e00h+AA7vHg
YIORxXxFeJzvXltJQUhyRjV6o9XFuElFxyvfseg5GGmcfNrRGz27opq6eohVMcPi
Gmi7lf/0E69SgLd2MG6PA2MKtySnq0+eZbGbYixjKyylpcDJLoWLcTHzCy4XTeY8
IKfoGMussnf2pUAm4uuru2dykpDnSmzoHDl/isiulUMj0vEgJiiDR8OKYNMjuyIw
q8gR0wW9bFUBtJ+HMRyVfyue0MVAifbvSq5wdzS3oRR39sKZ2qi09c4Zin0zPbye
z2a1rDOYAh/NBHPoOM2UOiBeH7/KGn8BXN4KNNOms/aaAgZMR35qSgegzJNbWKJT
l+TkoDKnZsrXXYeaDcw0s4fHNzcfw2lBJA0dYGlcGFWU8KYmW6odsSyBnEPEu1rt
pzPzPxb/PWObkfxNdwqPelLG3rk/PsVZ0g731noB1yGZDSVJDqlljcPeNLM7B/Nj
MiCngTpV+sxjtn4bMRwtbOvJQ/YcLWWbevMhPv8lXZhe2EeCPEKTCLIV+jrArzyI
J5hTfU8Lcp4CmF+7Qw++6l1tpsfwTq66mvYgTS8FhoeaKBg7dikoOHWoGBtNAzjf
iPyCNr4v3HjXzbivisI89+Vg0zHRwy9AbF90kenKwud7szB0d4E6ZvjwYeFqkEMD
GoeWIWWEKpGZC2LZlbIGOZNWikRNFHY+vFldGdesM4hBcAP9BTBpsV+D1Z6Sv8ec
OxhZPjQYKEwzWOwzG9YWzO42C7ZiFM97HwkLQEOLdRZxV0S1VTIuN3rUZskPauR/
d8T0IoR+mm+iz2AP2yyMT9LLYWQ3q9l1HpsGfHcbQXWq2lQK3TqcbHp5qjTb0hZZ
MVSxVjcrIn4TbKZyHcQQqvlQiYeRC2qgra+QtGcv4UVX3kGqRpfi6Dhb15vtux8c
KcmY4qJnUrVTUsiDcHhcUjn0WPFUQ9By1QbRlUvgSCWYF9XoTN5xHECiYzxm0Iku
Lvn4fLM5JX0dDh/eG9HopHsByoflfp3tcy5aBhjZvEd0KfulExFh1yzLtR076hR8
lBY1QA9fI6Wb3EXcvzxIOnj6v2BYbz4GDZY3Ox9p5siVfdm4B8fLiv0FhYqC0t+a
pqJ24JEPr1vCSKLQJY76GuyEl5Amu6KvClSnJP+XyJJUmPzm6RUSlEkGgzcor3go
IF/J8J6FxQ/PaKwrUX4WUkvt0fEQifVTJdVItBeHAoWnnLCLNWvdQqoqD+n+ZXnS
wKMntbgtpDj91fMzIz6daPa3KhUaKxqJ846hft1pItjD+CBZGg9BWKjITvIbMghO
6X1EndQExR2/bieAn4zj5XVSSXtfGo3pga8XqIicSr0mfikiaBbl/S7OiFlaHruL
pCgJqElBMb1KqReN/NVv3RWalixiGmg2Wx9eEmDiIoxF4AYzomdesL43TF8gcooq
Nkjih6qxqYfE2MVobdviiWwRV8mEoxxZVRofGwc0vo9R0XKFr04hS45iiQnXJGXY
F/aPVAb/t1PpqsIvBb2Ak4TuskiXPnNy2SNTcPKYCHHDc7p/HNRlegGHH31wG+pY
kiFO/HTSEzIGpF78qMdTL7L4lb5vSp8FwHHHXfj/+vEto5ImSOTxeBNfGrbcJMxw
paNQ9pGM1fh5ThFBsq7m6cH/FzpO+ZjO/Hi9a8TBeyF4PxZCXeJqPptpQtjmP0EG
1xCuNo5CEbutvCYuJXnk81GhYGUNa/9xT4BpUKfg0BKvjlR1jKtYD5Rs1zin5buz
J6PXvo8IfXd+jJYQ4Au4XvGIDgJmOv0Zc4cLTIzgO0Yr7+HO9bRqZZl0Vpbk1mxI
7NoCJs/7BSF8SxLRvdoBaL6JkOhnDHMGgSYPXCGw21WAgHWQ30Q/T/WnU1GnscEN
lvcE8ch9flchvGI/4xB5bWupJWVbKfuRP42+ccMAl6MOm6CVdTdjTMaPPqNyUfH4
TwYWPucppPc9YeUQCkBmdlcivjDj8k+s4DaI3EPlTC4fBChntWdOGhs1NX+WZ/32
vRxoD+deBqhzPUQlMKOxDKT53APUHC2vyQzVxfo06F6uR+YZjnrd2zkNM8r6zbni
vvHyUx/3EkHfZDaVFNFYae42Rju9xTZcBr+YxzfJGmoRqIKuCO0HHqHmu1HzUGBu
R2HmHVflcxzmWk+FHzUlw3vRRvcKJ5RIxdvZTAbklwjCokh2jGhYc1+evRml4Kwc
PoT0km7oSZieDe3OD4qJ3EmXEFhYK8pKr7SUFL7B5zH65DE3WG80RhZxO+vGVhVs
0ISKFuD5e4on+gjLPYU35S+0FEoW0Z4FluDrMa6JzpxHKGaX+KNEbdfI7r8HH3j2
QDczbJq63LMQiTyuVzQgtecXSbyeQD2HbvwevLnmpxY=
`protect end_protected