`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1872 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMWORzZC7bo0toZS2Zods6Xs
yljw+BvqICQb54hGe2JGpD/BBOH9keO0cgJ+2MpX11ga1+05lQLXp1uDGjAwjddY
U3KOGcFI9Xpuy2ePJYb4gmOy6OLAHrp+Huasvvp5/2QgPnb/tWkzKPlgAtD4TBt+
liSVJQUd9QGc9oMS5dzentTkPz3gHvMSfgD3k4/wAxZ7vfYmUtxIdfUQbOYomogo
ehUPLuvj/Ma5zu8G5rmCIUqg3vJgB6+v8STJkUxlZMOwBGjlBgX2ePWKf3rxGRXq
OpwN7kbYsa+iwakO8gpJaFrZVIowB3YdMLoL1lsQ1PJv/C6rmykLtYSBTmfTngQ3
zAsDR1MQQ+FwllwHRBzbl+WW9TS5x8TrOb3DJsEi+YB3ctgAvfqpkHq6+h5COCrr
VYHSg0k1Fj48RcSxzD7M2XH4gQiGRA5j6/Bv5wdpUtYmBxSsPRX/9u5PCyJCKE/e
CD4IMsUDH62gCiYAdcorDM9dmmYh8UAF3X1W/pB6Oi9AQGfKZzjYhwe6wrjTvp20
s9JAo8SXYNgD3eZKIKG+AiHwZ1NelLZOdrrns5xP+umZCtopA8UPLHqT2TxB9xkA
qvPemZmK8FGcfhPZmlUBvh4s4UBqmjXH9/TS8vY5H0Se4liJnqG5QfUhdJLfenjz
wNGWNqUOcedhmm6z0duSquvVvh+C8tINvLHu27WA4sTLcVamUxowR+MtyCtwsg96
HYg2WXMxXj4B4S/aoz41z8dkD4XRG8C200cNIkYYoNX/WXINbwIub8Lkh8JIyngz
+eiZIZc4av87UVjLdCjOn11BFxyf/PAOVfKPFahfAELK7r1SqBmi68GOxrMdbVvI
fKkv97fAU1PX8/y7WPbqcTbb0R1tJhRjiLnfywjRYp07AnHOi/yKGCqTqIcJMUgt
8wgaE8FsTRZk7rFGaBNPK8M4rblMkJVNcRVcYt83B8JB+dT7fSFap1on4TsBTu8+
PdqUFriIlJbfJHYSW+BAqJAT2V9W61+gl1UvavFzPnZIYPtx5opA9yUiANqxi0Y6
MefPjRdPOg0n8Am+RzQ/qcu7SKDugDnNNAmPCg5Dr0G+pglQnUt+cnvlslN0TNs4
DAB6kahoJEhvNww4TPvtAUa+SelLOzc4xV6Kkhpopad6PWCNHB9R/WxxD2ACHWxm
0p1V+bpPJ6V8f7zAzXr9twOP2xXwbk4GkaQu2a7tIbMWSfIJHAIjSb5shzL3kFp8
aKKqUFm1amVmtNl1WAXOBjcEVzGJ5VoM/be1iBdSqFDNyxlwi8C9ZyC+RS+WPK1e
4X+L54N54AB12XORXKsZDHWGYH3fGaBxw4klInpVPpdqUS73PWzi4Ezad7in6GYk
xqpYE0qVjrTc5LX8uAYvdge4A+juTwN1CpZS3J8aXeJkW3PnLlw0yMioCu7na+F1
YJOXeikm/pY2r6Qav8xWdEqjLi2+pnnnXk1tSbEI/+Y/4R7tjPY/96s6FSWnAIVa
WhKcaxpcmu5xs7n4O0FRWnDCHXY5HI3aEqTYOw+6VOcq+YVldqh3mSlTLnCZdNAf
Er3GMr2xTAZsvIHMWEq1k+zIPjTcHzhtt0NNfRx/VAj1argbdE+7i78SoVaTHBXo
nDy+DjUXjOGeA4bcbA/vxC8Nkxdhnut1H7875bou7EC/AbL5pUyybQyhIB9+ccTC
m+w5NwnE9SgsBdw3wFgU1PWQlSeuX/46ry+oMQjdmCYuHur4kr1nB7yhjC0afXzi
AfrOnpEfDv/qaLoP5QHYZuGdecls7x9dU9rAdIUQp2RmKUJqWsG0fyptkpUlQuMi
29FtY9eOtU0LvMI2RW4tvnUfLL1jySICefnmxGSLWgejCDxP57xseq0kLK6tVCqR
wH0ZpeJ82JG2oO9AIGUjdHVMLIyD2rryhKjXQ8c32Asnef4Oti/bgLi9giqjoo4E
oxO0EAIqqWeJ6GkBZHn6+qW2gYMNOroK1FEyOqMqXJVK8/NKb04rN76QDpJec+lM
lhW10V8mBa9G7oeIDqUoYFJB3owsCLXRM330PN9r6COCUloIrJhjsqZtFeCWKJ6R
+fXmw9r3PVK4uuJrV2YeQCxqcAsMtUv+0NnEUt2lGYJg1P70ZagG4Bs0DdOa8RFQ
5Sts5US0juyGdLdnpSSt9ppLNzdfIJY+1f10UTFSj5dKNSk8elWaB9OYjZDLaO43
+Kj3Lb2nYp2QBrVSkAl4O96YPPH80jeo7OvNaH7SO+UGSBqLI01xr/1YxzZs97vV
zo/cYB/QDAe55bu0502PjOLKSj9jF07k6+Ajqr9BLDX/fRUDkn2+YdwM70dEabs4
WaVSK+8zVHro62JO/wsNY+6oi5Msr/hGMWAGV8w8FbF4wLBx3WO9ARF06eiMe9Gg
`protect end_protected