`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8672 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRukXvXlqy9wFYzVV/1M8ArffFuNpvgl6KWmwBcbuLKhf
35GgFfI0WxEEeEcYUwXxYj7zS/Le6lZe5ndeWPjljqXH4/2EsILj35W5iMx1TLCj
WyuL0AypK/xiaIi7Z8NywL63Lik6T2mtDB5jVyKjOCMM2GPrkin4HJ8mx/zJvvMh
mOaTdblxEyF1Rdpa9ggnnbdr856e61bWJ2cEv75U95B98sLotHxDEhDJpHyHMtyT
QATW8ylJV4NwfrD7F7LfDugwAjvd6dXowMQp1vKotpOwiRzljl/OGJUblJQd5KCB
jhtVBqQW/1+/5LHEhNY2n98dnEp/k1g2RK8/zYnmvZqIWB9+HZfnM4W+PqnYuZBw
OKs6WAIJy82uShaLtRr/unlSH6zDNBbaMPMQyVzA+e2HlVw9Z9YSYcaL8sQFTFyX
l3fSmv6j092wcZqREHlJ3Wu1lOfFh5Mr9pfCQW2M6WbIO4I3EB9/Z6FvsUm5ai5I
KhVurH/ohc05sF9AKbPzob25nDtbbVVUU/klYn3ZYE6CZTQ94f9Pxhm+9+GNqBfR
jDQjYe0Cj9vyi3k3ZIdIFGBL3AkZoKDBub0Y1jcA99MQ5IdHRCJrl25pZD0/HerQ
UYmpQwcvBqxf5EM+8MmSxFORMDG41yMPL4kx+0PhuXRxzGVCm1ltHVbpXS5kauPd
1QiBh6QG2/UZ4mW31MwS/szYazUNo0pAFnnyQptm2d2+m7dgv7V+695bZbV71FU9
9hr4XWxUaRJmx4w8Ik4ym7iDGmLoI4KF8/Fs3RTWS9jQYfdvIzOh+xmhplE7+Wbn
5PoR8M5wH7t0K4GQYd5JSRGKH+vaRsxqsvV4kJ2plF9pF9CWscI7JTto4nZqrZ0+
yXbO+6WyUBqfuxhrnBbl05Fn1oHgYEcqnBeVxymYya9lSiSeSBxpSmqNdx68/2dj
3GwiOl3ZPFoPoo+gfzPoAZeuHW3UcefYhTo4lI5nMDJHIc1U+oDUrDqUkj0/SlES
d7bDtODY1foIsADzw33I/Z9M1LqBZiBVqY2TJyf8SHaj4hD/qwbn+a7uuuYKcv3z
rYK3wj0JXKz75bSHLqoZUfIQNjtpjRE3cNJuKHfg5hci86BD3Pnsc2LJ9CUtruOT
DFCugcxRWCTiUnIoJBsNtEQCzjFSJHK5qKo9G9T37NRZLHCWJEtJzFoqDNSml6eo
eyHnK2XsqCpBkQvnzQGReiXW1Kyna7/fwq4xuoOYEqMC5VKpjF1dMWvwtCVyutNo
bIzMI2TNWuuFnHKd7ShftclAzs5UckfI7IqWvdaKmCE0VJzATykgXkdkjN4MOwcI
v2zXjP0cuDlGJbXnSwgmByLfd+vlujLa/jwkMiMmuKkF6xNGJjkWnTXrNLJx10hj
Oj7gco/DpFdDxfNolHtDgIa/4tbtoVwbkhSQBnm8gbYihdRqRw9/6cakesoEDOHe
KVwZBxbQwKAYsH04RY+b1QOglA0Z+AuOd5Q0OhqH4uoL7E8SiuvSFRkkGQ1XRPlV
EsNbZwK0xfzzPVc6UmnB6/dtvyd2+0hXwYo29ReS1JHPP8dhqXMrz0ovsKLHaAK+
Tf++gtEWJ85N8Eya9caPzyW/khxmxzgIuj5L6fF0FCMLC8yDHtooKVlFJlM3XNRW
2NJq3wZIWMTVRP5Jajz1teVhECQ3+odnWTSnihFOBd9EoxOTdWGBF+LlNX7nhvli
9v4qP0gwsKAmAsizFZuJh5DsCZIb4YcC06lX9Smj69Ro8uqo9JdB40749T6J3tBQ
aCub/K0uhH7qAbdsgb02A1IqCw2Hdnn5qRzUpfKOIFvsoottYtIdbaWaQdwKNaxC
ARBVgzO0XXB0zbd6TerE7BjwUlkYBvZJ9/NAVGEMpJfZIBeruZ29IhW0ONUePblE
ERy9E2PVrBFX7WfyMrd0XNup4AJUMP09hwAWwg7VmN0wXMpKBMRpn9eQZNz1yMlG
HbBYyMK+e9bHvGXw7zQZh5+tjRtt3lLETxJkxRxJUscNK0QN2c4I/XZF2et0x/uL
/JqbHzz137K8EvusccFV22KOF0cCJtgPCIpMmh4HnzWazfUJAYeuKtvZXnIGbwKd
DOjijHsvaos0duW5lf7FtaOaM88l3k5749vN4gFC8c1Q6JAOVnfu6LITnn6vYQIW
AYDHd/c8EuFYwfQohSMRNWLE10UK1Ta4zNCF/rRpcFtSU4Gfqdch1TcU++7lZJ9D
1+rtOL9Mg9syzwm4V6Ek83jn1fvCSt2lSpNqfqpHZCR6LqR27IFBiKjl8UKt6b+l
KmzzcDYT64xqPgzfURUJe9VKyuRwjj4TGWd6XQ+j0wGKYVc5YavoF5CtKcGcGA7M
9tHF2flqCmG67HM1V3LX+4Lu9t43CPLfZwfrk9z/a8fvSPn0y/pmvMp/mwIRvZcP
QVqYUqQG4FmW/X12kt58WBNjMgbF4S07aXdbXz5yHeZrlcfS2S5ku5h6VK2hyWIF
7LGxLhHgdjdhnAwNDFJ2ld2k9WjBHK6BON43HJl5Q4Ji5Ulf9BvSv0gcEm5yq7Kv
NLQChk+B1PUAxjjBQ78ippiwPBkM1HpkeeU97xYQxgs7AM5nZU9h657M2jME2+Xo
lMxOozvy4wkStzmTgui+1W41f1e6oHy2/1cjkMB3XDVlueEzfCMhHfz8uSgPTkNK
aNN4fSFez5/lU34xG614fQw/NukVFUEnPuhaJwopbJcKF8yMN4LVXiNbngAPvXPY
F2H5E89SCbyewteC+U8NS95buSRdLqClrFRsDmEpiy1bgqB+ZGiyTU1PhH7rOa28
bknsev0InEko2YCLW3tMofoaK9ayqIuKL/Wy0tzG7cZVGiSByzB8jFc+KBJiIQ2y
d9rgrp/2MO/qWDXmYXQnRqqIeXL6XT/o4zIMsAip2intYNGO2lpuk6ItBbXa6vP1
clljN2NCfDMDBh/NdTsJs3zvzO0ErXQUsAZi2iy53NVhE7yV5kqKS0FAwNpl2J86
412RUCECsZRkA4rz98RRD/YYpY0bjRl1XsckK9tmVMlc1qBW/gpQWNJaozx2nGS2
BgCKp5zMKiUQ2OmdAkDisnO8alwXeqoZ1o6v25A/Y1w2ifR1Z1YDLCe2RqLZ8u4A
vQgetB+joYoJgt4bVCoVxO/lOXzQEsk6H4ptlbjulm6XiDc8owEAGU31wP6EIC7k
d1O4UtwDK89dTLyZg6KLgDSsZgNV7AQmnl+d/2U0cxWpM6Zv8xaUcIVJ84frTNya
Ef/BFk9PzLTBx2EjxRdU7IQ3sk/sFKxfITP9gtPvpkp2i9777h6TGE6wBZc3dHVT
BpsUPyreVfWmTLmAiXA28xWUpPkOghNOg53+IwlJP8o+LOQQDLH0TDNqxxDmjg5X
SOjczRXBojowGCWOemdt73FkdMRcPZtxABV2KDGMQ6oaPli4L7PvrF+bFszU9vXI
zqLSSbudM1/C+EBcB2EMhrrgAzPrL/MmtsJrGXiZHsldTcfTzYf6plyj5NBBn/cA
e5NI7UNHlmsAY/Fp3AekEBtggwzTObRlQsSTa7wvIQt9n4XEkgDDi3rmZDzHKG4I
2sBHNDMi6jNu4/Rgo80OYS7+aKCSqsFFhG2B4O76h/4xnMQEvVkAVatEdq0lg1rd
daSfzknr3XUEcpHJd0Hn+/H9QanlLIDjpNyPs1HYU9lzeK8gvr0+ehc8SA8YVv5o
Il/JgLj/aojhI1LksNol9u5miEzLHtGF+GyYOhjRMYMtoPYJTBzB3ER6WGf1HiwC
E5HUdy8phntAtgPldLebLGeeq6H6jvqzoN932w4XHgfdkLsSEpG40NBVMx4fMyj2
e8kFnRL3RBNOHYxi45kc86b2P/tWTlDU41wk2f3VgYCiNi72QHsxLF0aYNRwN7Zu
G3mJny9LwiHbN01PbEI4LU8gy1hE8xiFKlW/M//jFHH74tV4gUwTWrBVB8OQzvym
rjDFwiXKJdW+X/hxEE096gMrLe76QrzcP21a8BYkTel9+48lQAo9bOtPWSTdtfrg
mb6sxzaduy31ZLGnsUh+VCpw2AeXExmeqALKceZbqY/8ZoymxYT6lVxswVXac5iN
1/6C73cU70wiHeQRtdhQv52jNMBnhaILCJRH4JQLDQatiyz7QHqY4+LfB3DWwX2l
JDYmtNF0Xcg9/jWNWejDN1suyLh74JuBgQLIsZ2qYdES1MCOb/9OkaTA6gMW51MV
In8YMfLJotlsNVObVGFXRD7TIR/E68vJm1z7OqhPMzgmy7g4/oy70kNYDrd0ixoM
ZpWZoRLBpJFgftyggWu2cvsPKOySQkto/RfmMoC2Bp/taVaaVKjlUVjG8CDAgyMt
PJvoXZV4LWk3txmFmfNMKrjLdJ3LEOePeDnP0OorGy6oTgHIXwBqETp2HOOcG0af
4xAMbK3M7+C4N6aklxNwoJF8UUfe0hiEQSPtYrmLepd960+hZNvwZeZJl0fG9zMF
XocTUY4B1oCZJxani1JzUFeKp7iMQmHzy89SvvUIXORPKXkxeiKQH18ABqWmDiIO
2Wd9ZRqmwd6wOJqTCoNHriwYpDzcu1YLkIYUUQM4KeT5ybkD2lefaIwi51xuPpNb
EBTK/baupZIxCbUi37dVAy9zVBlTZ2Z8RZTVrZDVksIo8YFR/3yC/qR8x3X9ewOH
Ks4/N38SBszM60ptgiCuwxfKmDgTWEv28LhasuLza+uf1+3FoOPxj4UQgIK61QxR
1pnwCn971ZnFLJG/H0+X3Uwlnbv+vnxRuxDpmKlrS7/5XocoltqDTqpX1mCoX6GJ
xHGHlIvHkoyv/bAsOxQIjTfls8Zs2IKTtUT4QSYTJrJwKpNto62nxA7GkKEgyQgG
MK6J4e5o1Y2ar5twLnihBI45IzSXuxu3bFY86JGRcZ1bpYrPWsgQudex8htl4J0r
fFn1mIXmjwB5qWyzSRwNKUtwbJMaOZxc1sXD0pt+nXRgrYenbNy3NpLbaWt46Dyy
SBW2nqSCc9dzrscQnh28DDK9ddCOri5+7dlYgHgbNigWo1nBgmGR1HU/BCDkVJf1
frdImXnflbE1E/e/VJAnNoktaxbJuKnio/rPZmEZNUkPwcyBsPvZNdqZdezxXjXn
fnbiRfQu+EHoZTx1pWgW1uH1klB2GMU5F7DT/bcnHYfxI2NZp8xJzOwcNhQFybmv
My8OZtobjxqoFuNZqqEehAlcfhH8FnvHB+mDtnDygjPkKLFCopOibbu4LoYqDFXF
/GK//AB9vvXd4fUNTAMASviZfoFR4ZA4ATm4jb02+/PEIdUOS40YGaVbyMCP5s/e
/fs9DfSobTRq4uvl/4Et5BPuNAj3vhP1ry4VHH7jcDK4fAPDcAlLV4uM/VM1hGo6
3U6eAgY9y4s/SMQ96ITcve2RP+B/ZiZ3TXmWvzf6H69CRRL/i7YhIhQuXxRRgC0q
kvEoCd6O9LUpzS55eiCmgiHmMwKuI8Cqxl7mqOEa3XiKubhF15JZCR1WMifKtAb1
pzgCwPBzMP8b4oKruXXVszdCEAK5iOV9+2uJkeDKZD0TTX+yPZEAFQ6uw+6T2Qru
wKQT8ONDkveD9dvOnri9p0dyXsj+KgC50xcSFuaTYG9ElsP2NBHyw+l2tlzot1JP
18OzlmGmV+n5vLIsPO5ULwOOPv9z3mE6A7vhBlmL9nGKhv7ct2sm3CBk2gkbEqIz
W564OGp3xreK0UZIbFOybzBIxufxPt/K8fIfcJqtRMzZwdZ5D2NeHUHVpWVsZXrD
pUe0m3yyZcyCH3tMhBUgNwiW1uCwQfJ7bJcjQfwprVG9WTLgGqYQe+wYR+kuPC5I
wVpqoFo9vipHEqNSotCoRlX6Zgdkzskp8xJYNVG2xwXVj5uGLMKjtj3KxvPhZzXu
Ip3O965y7rlQqpKZBwgnKlwmj58pPArSMabSEI+ZlImnWTWfr2AyJMPcA0YLvReg
bL+jWVUva6HryCKlBh4Yy9R1TArpNQJevAyfywHz4wL85fy61A/WzmyiQKjuiMwc
JTKtmd9sDAygS/Q3HRN6r0/GFNVD/uEVGYlpXabUOYCaM2bvI3VtK93aYRkS7d28
bhp3GooTefTRg/ee49ApwBbWTdVpLaRmrf93ALxaeV1nbKo+Zs84OP6PcEvIIElJ
s1Zx3zaKT0VYbKOB31gKCBmwsNELBLqrq3XWzlPpDfVeDBkGUXu3EH1xPNaGXnho
6TLFx8Xcl2KfmWDW/SPZ/Z4jDBLJzDZBZYkFm1mepV+JgY40zBdkJf/POyUphlMa
uqOQaSc2nyrpUY13Qjv9Tqcy4yNymYPpC+k5KoEMl+P+usdvPpRaBFKAJovrt5kX
TftoVJNRYTdJdz/dZib78/y3lsD2hvzwK2JXDgeW7auijwn4uebSxAwY+eKXF2aI
VdzPHbTna6TXnjxvcN+nCtlLW1GpErTI/O+uyuTZCOX9oWcYXgBK7DH0M6BqK7Fh
qcjB9MYfHBUqpCqY9nvpIOy0bPeE62N3Zq1XTMYOL1hgAVAvKgUF0hEpF1Sz0VO4
/fwyqNSKEiOU1HlBD++2F5sg8Xn11bvkrcQ7oh4g761wUqkqOxyBYfMVn0Ou5Sjd
SPkzjfa1dTycuyLRa31nX1j6knfeffiD/NXaHM5gn7hPvLCrIadXEY4KQHhDJF7k
tDzwUZyhLe3RADqRNhkAzCopOA2nHNaO9Jye+09ExkoV/MlN7VeKXgYdW25L4DfO
s0G2fHvYKxX/jso9G73GuwjJUzJGZPRAn06bdw2D8NRrNqVgOy+j3W7jm0Z6tfpV
UHf7xKsrGXPIbmbqKuae2N4aXo9lX8/JD9FnDCfI4yhdI200s2zSEKrW3CMYQHnm
pQ/dzhaFagctE122v+GMBiTMCn6++CLyUqKNFfDHMyJx4/QPxsFFDRywVBWq+l1X
y2To8MB5FcTSu73V9BztPmrVrw9/rMfn+d/JXYtqBrfPvfjssWQZqgxyKo9dNmgc
OInoogp+jfWsFfyxoZOCAsVoWfsuLnC70c4qdKDSctmXLXX4TZ71hxJpv3Mh1hXh
DeMw+YreupVNGbRarMOAEnxc0ELaCTJevGt3hMspSm9LygD7TFxj5DSHjcXl+kUM
rq5BVn1SgSjEGMjVeXY0r4KExPOlaRvnCAMFWLIsTj3JCcyw8MYzggovIW6cZrDz
8Ybb4nzRHnuHUwn24b086J4Gt+P2w7Rc8yDdOJsV7SnaWvzlZoObnh78XzvWTLHK
v1k2PUImmNndGXCA8jTx8D779I+7Que2YHTHm45A6kiSyKLvma9bWV7fPT/mlZHq
52SDfJ5vs8FYVDiUVplripnGFw/dn06LhZ1ig98xzPQEk/pXjCnA0p8MgmFhMrg6
5CO5fDr/Kmk6w+vfs/Ht7f1srL0NklaVVoWe0J2RVIf+N/En2cA2XH+k96u8QRO1
SRqWRoP11JXvPMem3xRDUGs2OsWsMZomWZ6/cEy3i9jjpATnqW6zj3iuiN7IUkxx
KiUEOslcqynDU972ThtVLVIppyII1CZpzMuU+haNgDTNkpeevLAatdkECOAlRvbu
3klsY+LJvvU+nQihSuFIBxi7UirfeVvzbOn+nYyM8I6lGqfDuDlwqyNxzdAkFIgf
adVvqZRHzIo6lLTDfspJsi4K2eyX/VBERIiiIO6+5hmLlfKhN5R8lAmj1AptQU2G
4XGIb5xBPd4oYPrI++AZQP9pnPs63r//h/F/OsUEc7X7GUv+w9Jflrox8KeYcY+r
kz2CHtWHAGssivSonr6RvxUDGCA89WMxu8BdzzsmxyYRj9bjZ+NoYBesbUqasGvQ
wWSmZT82yWDzDPArtdq5G8juo1hZZBorkjAdI6mf+mGvnD08uBuWZO7V5u4vbDLY
55KOnQ0k1Hrb213m9onmRDQZAa/M1Bk9hHUKPtT1H1G/cQ7rkyOJNJcFPsCkklYS
FdctreRCHOZdh10FGQh5AQgLKBYsuWcIdQgkoxYb8FWG8kpoHbOo0vPZ/PYTLp6a
JmO4eSl5LWKRly/GvtsQi/ovnkUkBoj2NVaAs96ZKr3cB94sHFdJAfQfix0x30pt
Udi0OEt0uufsZ9kNbIRbEQqF5Vr+B+hTeNK1TjAWAWwzvKQkiLbXIkwnHjD//zcu
p2HENO8nWf1F+zO4tXVZnAOgBUQWEJ13Us97PkbPtewgcB99XEniNsDIBPmsBgBF
u9jRr32cwDlSHjMl4wE0HekrTgc+SLHsESAWrp3Q59EwiAfvgd1/7KJ4rY1545nR
OBE/efh9NxTuBhYsfmHl0PcHgnHjZQncKL8XSSEbgeFooEkxMgJtjDhupP6pHW9O
W77m2USdEAb3h90Y5WcA1bRv1TfXcK/vTxAfAbVFfXb/9/uaRrujJT90r8XutOeC
TIxSCkaV2RorkAldSVANkFsw7WZzNIpFp2Av5jJUM9E0EcTASORK209J5UvBXAgk
njc8Pvv0NsA7QmeSXzCrc6W+wDeN0MYDoWf9tgoR6xzkrc37N5bE6jMDkAAFROl+
m2Xt92q5bh5IIaFR3Rwv/iBMBGYCsin+oUrtYAnfqIJ16HT20H0KfrNRrkAPOuDw
/dIfHehTReYKLh+YWkuEomcrr+HS/3etuIWRrovaleSDGtches220yM+UsNRe304
kkTDHyEXPNMfsbfWXHudrPUx61eJDHU1ADTjs2sV/24hUsvaPHhFxdeVYhq25rM6
T04g/28HcqRl5CPXwp4gu38SdyKjhCP00ULzePtsAf5hJsPqWGBEXzx/UME7efyw
L6BqTKIrLL2dQ0Ipqumw5NoYNR4luN5TdD8ecD74PXRtIEW/e4XmcimMJ3e0d85C
7dT+GX8CR6Q4S4VBT/YbSLdbjWlrXaWz3NxSUWqUVz9iHlQAMrioqHHpztbFXtRa
+ksWMMGwgjDFFPLGOuACkYSkkPl4n/ppoGf/LJNpUtBd1EP6RXVKLTJlJHualIB7
sFn4d9KuIhCkmOqppAGxlsVDFtHfBe/u7q/x5fVMR5YLGY+k9HU1fGc0LRQ1pvx6
jRK5Xem6kd3iusxCweVnyI3sWrKRTuOBoimz25OoYYrJxnBeWaJgf02Cv/wQklsu
48a3x4FD7YlxVACbFQtpU1Q8MbZtQEx46R9MLb4Sr5hqv0VRXFVjzB9EDxU+Mm7T
e2sdaUI1JfC27okC9Qp651KvDxsqxm0V6d6g3flT6GWZUpjAf1ZoxBBTxAHuBOxE
IXs5ofE0XV02GwaYfRNP+fGrKxQiTP9jmlipd3uJHvpfOEjvhQgBQSls/DANysMg
ZgBATtR+t925KK/Fv5VC4SdUZuFhXznTkJB3FgztlDhlIoao8duzOjSh5IF8sxJ+
QzPvTg9MfZDBqMQNm1faIia7oyA/b2Z/kDQ4y3zVoTPGRMamezdptT70XP1FAqF3
4Ud/z7aGvWF/KK+IObWR0S+YHjmJaVW68CrCRFWso7c+ipU5ZLA0kisJ9QDBCJij
KgSOiINNMaHXOu9cARCiLW+buwkANr3K3+b/IQxJlOFcbFL60BABeFoL/g3nh3zP
f8wnx8ZOi8sn1BKOdNVzjaTPJxEWLoI/1LUBG4Ue/NvH1Io1AI5L53j8uPOAq4zY
Dmv+BczPh6DcEGU34CLu/4og8PxZM+ZLsqzvgeX8whmdvlSclYmfADAfOa0M67eo
1NNOl9JwveOvx6v3GdZnQLUrC9/4mCGcxmZ4TwX7872pUDmmE4+O3CYfSSr9QqGV
EHBKkTT+iaOXEoxucozNVfOj7YGF22J3yfIh6iFyHOqKw8sBsjGaxrzWK6SKYhvp
u/CL5qLXNIcK4JIgfH91S0lGAJ1Yys+L/a49LsBTX1KPYjrtKyMZoV4KklJ6ELhI
8d349R4hO4b0mSXWlnvA3JFcjjya3ExDuyQUO6m5ZWEKEklfTH3Zi9Fa3sHkEUp3
E2MUYvm1bTps4oIdpvZgcMnBUa12ncqICvW7yA3euvrcenJDKpJ0xfLKq155nxRv
eLONgxVqc6yvOBUvs4JkqOADL7GESUhZgX8uZ7FFAhLwGUcy3ohhoTd7cBbO/Lhp
X6QIv1TjQZ47C6JhUJistecffJ2v7F7pqqSFEnMgXqeUt+YWDyLz2oVEAd25NaW9
hcW+7e598I4t992kImWcYPj74GMTIRXjP5Dr9gHdsIhrfR9VPzFAoUGvGLDNwCMF
1YmqSUuy5TZT/NQT8EyHvkpbS+hb7H//kY12b7rghYkIMAtmvQehs3WEqgq9rGqG
e9Op6LBraJbiRFcfm6LDXVlT8IutiNZQ23Ek8RGoZX96cLJHFdbyorSEZcgdoRPr
GKi+7wmnkEjIlNN2kiMOhpA27hhtBJ3jjHZ3/x/O1nEHNV1jBr3ghOdGQkvgK4AI
o4BQ884zAeScYn9ryUG3f4aDipXbOxsBHcMF1ybIzmQdHyCDTkf3m9H8lzleJ5mO
lBxVFKs4NbCM64yjI/8V/S5/8vJq2I9oLrkovTu5E22f/YMYLEFjbV2Cx3xJHy6K
d4hcRpOfwaQeB8Sx/De2yGdvD0j+cxvZG3aBzhuk7a7iicKPkIWEn6RYfE/4C1q9
Mqxs0ESmJd34dWumbaKwxuAWQF4BBL1JSCFLI2aU0Aev1yRqk5cRAkaO/Qxbm5o1
0ayCXYyJykxt8U5uf3buh91fjf7sCzJXV4oIqqWfevKDnggwqlppF4wDOuQcBoFk
ih7RNgkSuXt+/cwwW5uird0tqUwrVJHCUNTCnPE28VVoDGJP4H3lH2uqpNNVujq9
byU79RRZQAoH0tu2Egw8Iok3s+jcQwdjYsGk5pydaBV/Tg2v85fDqvlhEarxHToN
rN+kWPMoQchW8TswcD6nF+EBW2yQUIJzymRznmlJMEVt8ugCWp/K5ObMjfUtM5gm
x6OYg3ACQ1tsZjZt/DrIbHlQu+L5+miWvVOaHWUfixm8EdLx92kqgTZYJAyNVJio
NHSzD4rmihgSVB9nAHdeQ+GxAKFm3E4++DeAIkjW/3ilcMGFlpf1HANRYNep42NJ
kjQLa5EEpgkpgIooUs/VS7IMsIeopCmUjGy0lBi4IbwmVDE9I9cQXlKsvVQ+ctl/
Wflvt++qXzXv0IrlKquTBWge3O6clO+1tZwquqE6dKB8ENy8uJI5x+Pw0f3h1Hez
w9Gm4DPGNCbsjgqIzHYUNLBxTceDAlcU27UwtQTPkmQNc0cXhto/y0NLgwsfTXTl
zZpfQ3+1Rn1P2mI0EjXnj5rZCUPQ/Mpz2xto554iiON4uSSutT9AG1Rxy+IRbAMb
vZ7pPs5jIMPG1dtn08ZRXX8DPuYfwaySIjY0BadsDblxDYhi0sZ28CrdQRIeK1UR
jGucZnRfQCxKneLMzHs8Jf+5yNqxDV8hUoP5sVBJx6KblDRAzTutG4thcgdRclFq
/grbDR6rvDApWheP4/FlRzRmyNkXmkn8fPLd0Gd8ac4=
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8672 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
/GMbQK29Y+AAYqzOrLs1aeX9seC9V7j98AHI2NaHVkyQ1n9y8bgh0Zm4AI2U9pG2
VYFuv//lNIjVvWyOfI5LCMXMJJ3JxC5s9hV0cXHsHbHgKagdCPg1rGpDH5MTJKFq
VXSUCMQmvt5rvrcZHzWI4JFY6V+l+w+mynKPUWHbFq6ogT34YGwoaBcrMh5ykSQG
G/ufrWzDzRFYoWvG0cOFg+pIRuimngoxEMzWh2BLKwn8hJ68KbLSstvO+MGE3GmL
0WhyfSMu+H6JPfA8eaexp8IxvCkVRCl4ZIkpwldRA2UDY6l0xyDJmPFep19s6xLr
zov3HhoooP/XqSncMKl1aFTV05Z+YnDRkL+dKzjVFaIkPlezsnktZ93mCIx2Ct68
I/iz56afYUdRq4liPNY3aj7qD61luG4AsN11x7GSrWXUvcrJdBNI4mbCYKs8U5ok
tNS3YE8aQiWybfic2QBQBe1trlsf1/eeS8NGWyDB1F98Xb0j+yIbqUF9RPuW3HUx
Jc0CcHYdxH3JBBwBz1KLlpvd63tnX81UYbRB/0BoYWb3YFEMsnyLbkFBct9p3yrv
+LZCY1/ljc/BXLEMOp+Xvmc4piF74Rh98SguyEgr/rm+KQIGf3HxCIjy5qvyM0Zz
q+nCJ6SsJM+0oVpEerfBKwWWPzWddq0EFBDx1R1AXXmfPhYF55TzBjNJzGmrtmA3
SZh9MlUwI6zwqwRC2q4Tf9jvPAb3pkQy9qmRZCaZB0nJCLYs73vOXa+TBdUklFXu
euq8RH4Lzg+L1ZpPQvdz/8GOaK8HDw34fuuycaKgl99vdaMb2IHghuPhjJi97o5D
mnRwDSXFW8v1Mfv9j++q1VhYFR1xu3P3IuhM/+e3LEfKu4Xttbb+J1EhTM258HDp
9txT2BqhhSfMRKzYRwc6hZ7UnL1bkF+ApQFXsl7S83L8zwvFGT0FdAUwpL3OI6Fy
h4t15eoeSqmTrOj86PwohV1i+bO8VeaYAGaqDMrKu04jDO3a4sQxPvjqHNZiIsVe
mIVwB2uY+ObAoWqOxN8UDbWuB/vws+7tEvqBO4xtETz9DIj0g5XwKv+rxX+ng3q0
nIgW4jl5uCF5Tusz5bWgTevZKQV/3qftfZfAB5QnDXk2mV9d42o9rwYQMBMEzMYa
QNq0gyGBkmB4N5UUc99hX86Gxks8sCCLd9AALGoIEP3nrQIPYHsY6/iXfKLqMnBh
y52JVdGDuEzHsVHwQBRhTaYqqHgMuVLAilBaEp/nyhH+LlpZb6NqAfTVIfIgQvhh
B0KefoOkBiVArwHvVIaA8x/4z/rkGfaG7K1DnpK2VG8vraQvNHR/EGk1EKjzcx4l
q1K69zpjd82QAu7imMw8UFvJtWHyew1E0DVi7dapCTGi0ly/dJkNcAQM6l/K6llF
B/NPK9bPHzxQwc3MMZitePIta6sBNyzqhjCtQqHl7TmuTce8YpwkTEahKv4EamEZ
LvAwaH2supzQ85j95bU2QRmq9LFYC7NefiHZMRH/DL6K3Ty9RmmDsnF9tTc444C5
wi2iXIXbhgztef+z6g+decjTeEtDpZ2oBqYyT/hpNxgCPk4yCVw5J7A1L40PK8tx
Vj2FFZvfic82pi42oggqgVl7nqOuj1fTNSbydFlYVFiL8CboKQTAb9yilCAbH8QW
NqJcDEQy/kRCN/weyCoiYxDXGnnhJPn0y4dmFBDUW+rMTInJ4YcmVMb4vuVWclFP
VUGg8caPtuLN8neE6zVT6OFYsBAKwc/Ar25sKE1gR8xHBLzfx12KrVjKV3KfonZ1
3OLMIr4IQOOMPgRfrCDTtyZF8XwD2fk++zsO6H+KbmrE3GSfl2jDBSZZGCc8Z32w
yks72BzKifJRe1SWB1LLL8Ec9IRzariCu0jXVs/G1odNQh9/DaAOmsw9FOUraey7
v2/0wKylKnZgRozaEDK98g/tEKXDqgCJhdDOyrv4ZxkX5KaqS+0YoddoGSpPi3uP
lt2FS8xpZGgw3zNUK+SZG/0NOIib9P4h/OmiMKuevqXsaEYp0TTy1IWMAJ/OWflz
VW/6FPZ/h3PeXYNSRw8pi7QAdoIYZmNAXKSrP7L/Oh8juHCU3SI+c+IM1/NVZr3+
0bPzSvkd/8jPUDeeREZO28JceiIs5NKjbKUthFhf5eZGTNhDOB7NZlswiYhGMsn/
relIbziZSMmYCzpqIe9tdPAH11aJcC1m4gbHuSc9dVYqouFIcDAvpxLHtx37aUJm
V1yYAHj0qfTBSmCEIWH/j+FjSpxJ8vey6C2+Jgh/Pxnm3/m3AR6HoevcEwqYOZaD
wvP4UpGE6TjPB1T4puMtuAsvGBHbVqQ1SqE5wNKyG5bdZUexBEKtXS74HRwWV+bA
bg2GEN+/qsUQ6QfBmqPvGTIcAa6vepKLUCghy+ns7XS9e8reTEPChsLMt+WGDpb6
Z24Rou+FGyvHmv/8jhsKI4Dq2FXY33nM/4ThGAAbVFwaJC1Qjjt9c6Qbd9tdcPTh
SzNvnrfFAF2xXwC1cTiXkyTUBxseXzGjQIPKUVR+p6ADShWlwKBtfFeA2Fs4wXIn
MR7AiR1T/oFkyy7uWgssHpvV90mCbCoW+5XKprfPkMs2gDukKhwWbU9+wZmiYFl7
T9ySro3DRU6uGQSDl7dzq1Vl5QFyTjvzQ+FyMrRBeCkytq8JsMHUNV+XFXdFNcdm
tTipZ+hjDxId2v3myXVnHvCjvs/sol3ae5qVmwcCKLo35qZnodBbv/lbK0gMNOSR
P6ce5qbqabtmBR/W+VAVYPGbBUzu90+w2YCePnElkDA5J3Y8R67j7jkheLVctnC8
oV8wNwYrCTmmN49RS4jD3A61aAnhzwMSATV5cDE1Huv1mdu8mrzt7hpObo4aP1s1
015rK1MI9PQJh36ScJlcKAC6lN2J1JwcQR8mWjFu9hhlMofaPCpl+ecdIii+rMfA
GskDoe+2vKA3KHx2XRGcraWSw4u3q5wkSlBKjoqja679cCaVQ63zKmoqfZfyhWAu
wfLoKi/hFnXbFMUBdkzGyleRAscp5lxbYSg1DGX4cxobvZCDu4sQ3fVsoi1MOgUN
9/MhyyhBjS0qxBKIkj8HAwv5dbXZAhXSzrnsIcMCM+LYtDcgf3lmMHBFmw/RR5GF
Icd3XeQvkcCX7Q2lQsSpIj5zxGN7BTUJn6XIwtyZnkQLpkutPhNuj3y7NNFkzBYr
cDM7qwm0c7e6bFyDadJ4okWsVPh6m0C6ie1AeyC3CmFLLNsKwAXSFHxc1iCdOi75
YapLIGQP3kUsyLshCG9UfpKKzMGPPSWf/ULeCC2wCFVmFwsA2dHGTbestOIBMu9v
v8NZG2l9hxK0j0+y2P//mcJCNjq7o3xlJapFRac6JYxyYmlbAaKzJJmkiYj0z0Zv
4BleJ8NqUm6tYiI0jym/uR9gdogrp9JSlTq3PNn3ynRx068VUjhGLIsZjj9pCdcR
MdYKdkGH2MpPWFPnFdcYUjx9l/R6al8kddH146fvSe0MYdEhHO2B4eurj3W/JnqS
yTvDXvkq0U3zbA1KhBJTpbrdIabmL0d+7y0RrLY2bG6hCCpn5w67Z0RcUuKWC1FL
9bg8UXKWoAW8pCZS2zsI3kFxf2Y5hkAQx/2/s8LZ/ahCygmTsK+XiAOu6wTgfi+G
pQs3hQQ5GwhxcKOsDwrEsuJ+3kiFxKiIYhZOgORTb0HMgGKNhn/TUKwyHSdZQHd7
GXWdiDjSI9gnMUz0R5VQ/QYaqp903R17mr7NC0vza1fzNOpX7tCtDtflp6h5IvX3
wxqFRBtfOzV98GyTw2q8m1AiofRMDvnwqDIW0GJ7OSdjYpS0JK2bDMjNEKHA8Oiq
IDccaofsPm1grlJwd5q+HW5nwZtXm0opi0kjDpp8tPL4Q6SRvrDGv5IiO0jWYdr7
2C5ecXeD1ZZRZkJ1oZYB9N3Xv/HRPAYL1TQzBcSe/NEfYy6cgc3TnovFCr7qZv6n
z5+E85NF9LQTGPqfzn95hF/jsXQ5UHOHS4RttC0+CeWZVdqfoAjajMC5r2hwR8EX
lK5vmwbm+vFB6IwjF+2JbD4SbuBN/JjiFVhGYPRLjHviX440t7mgrScTZWeUBeKc
fmLOMxEUt5n8RGqfRqBl2n/4zrpF+yI/YZjcYJX91jDh5tw1Y6cKcl/Anzu2t+eN
AGgjd08krflsWciMbzfRkmlUmfak9aZ4RdbPaoGunMcq4rcGa+0659tdegRoPKDG
XUsoSnSj5Wl45as9zSGJViHCILV/fqVUNEUTeXfNQoF3Dk6GLSNHRTZ5MCjZONFX
pXihgIQ7LSfuHPSsG5JxghWcSyTlFI9a9CbYPFw73C/pOXcR/uo/6+N52ZyZ6bs6
s4YLuqlFi2PbJo1RC61RqcdnBjk8mreU53GFqP6FuDdLWSvE1H+lJJgov+DDxElO
HRSG7EEHGVuPkRatnI46Z8aL3bJ9M/b+uX1jWka1NZXkmlxbTRVlBVuOyq3Bcfri
bcI4RXrG7V5L0fJvm2JUtHLYSmfEOMBSMuyu0KN4pcnOwb+Kip57lic28SsmYUv/
4epqxMlKf1hmMBmyiO/U5w/xKEpLZDj28lImQC4mi5R3wD7rboeL3pqYGPUkEXn6
T0bmcWpz0kaxNNXWFXeeYJEEC+d6rC2fhhvv8RbXNX0YFnjBtKLM4RnD3zQwWePp
Ls+mfoSX8AGVMBma4kEqRwfBmZXq60s4BDP2o3QkihJZxTbtYjSKZrTEf5vlPo7c
t0TEIl2UAoMgMy06ql2BJ0Rt1E1IgwWdW1eoJ6i+W47ALFRRrOCAuWqvZvZjNaS3
F4E0+dmOHaFz8KJZ+5keoPzqvt5+dzlJ49JJ86xmfX8evWzemE13jy3uIlueXcHY
ZKFjDlj9xG2zFKesDLk7Pm1F1u52nrBFb3Pe42XUxbEP+nUXpK0GYOBLjIvmFOAY
LSNbQAfiZ/Bm982OkUXkRYpxF+S/+o89ab0PqnlgOtg2NipQU4ocfhsjf1tl0OxH
Toe2LfdqocVW7wGuAx1C62y9ZbvDIxGAMoy0sNF5jcwhiSHt2KsuWAKyFtuAUkGb
drntBfV7QadMV3exLXO9fiRbR14dZgWj/0c0KkfiUtqvdLGjHAk4tACszMsKDKhE
JEcYOrKOHzIdeLJGxGyUvo8KbN3Ryeg1WtpeNIVLgnxQTqnUJM1FwlFlFaAh9PPo
et7/IB45atvCVH8z+HnNEmk9atF42GUfuzAxKjp812f1ZARUe3SBGRv/DEm+CPQO
j2IF2T/OcagWAwbrLv7OFOQXcE6eYrmAcOr3MRKSlm4d308L+mgExY5HlzU0mOfO
Mfj0dtrU7aXP8enPvXTFtZf3eTBHaWnhBYZy71rtVlMN+7fWc6BzpkFzUARTdrck
Nm7q78S8wxQk7cMmCuSqqT2VAqT1E3c75GyKnrVDVZk9iWBfmY7FFcCiLGVAeJdC
sems6ZG1IsLRwJegFNkIzKXXltJyJ3ar8W33qJLIwL//bBhP1bO0MwmUhHeLhiDv
Y85M+l+609qRdxjfKz+3nd0Qs+NW9XXW2IKP7txSivrp52Lk4pBJFYucuwCf1MOL
g7mi5P+wxKaiPLOK1P6qJ01tPogzuQebow8D9UIzo+5JySfE5/xZnspHQ795hJPR
IePEC0HW7MY4UBWfHibiq9NliEiOI2Mxw8kPAX0GZLinALy8IyqFNxC6W2AB1Vtp
caYOyKX4NqdaLEA26k+2Ed4t360R9cBIpYKNjq4nR4OdwpULh6+DKv08eY6XoNIV
o/Ve6qnzuvrSI/sbM1kXkq1l7se6pr1k65NS9sfCH6Q1+vsJDM/Tz/LCfuYQ/zmF
PUXRJwRvB83uGU+cEGH01ZGxJ3f/9vtWL3kRMVweyzbTfMsEhklUINg9YXHYaK/P
qzCNsAd8IBhJB+JhlFXTJI+hjmzxdCJKFqZTbWN2501rsWYuaadkmyuRTAHbNbnh
91NdaFeIfq31h9foD3yR3DMb7GsCdITGSkEXYgmj+2OsmzsxESqCghztyV5HVQZD
Z6ZoiwDlqLwtfiAkP4DoqhoL55BtHh/eBppFi03PgksSRLvRexEi7mxP8kN4yt3g
Ha+iyGhr5qdU3h/br8LGZyGWC3wJgCE6BcwZoqWP2yKWwyOw18DfIjewCA+YVcjv
EMdMeT8pvTnJUxbg7jsVI4IOSdAZU2znEkC0v54RExezN4d+1krK4E8takaed1Oa
kkgB3QDskjC3lN2O7ZNDINmfk2nx7Qq2PfS9w9QUMvbccXc0QqwaZGZPgTP5DzXF
6OrUe4IaxlmjuXTwlyy8Fx53HRAwd2JjC44s55qYakrTkRO8Riq1VnuBaVbalZ5N
IqjLsaDQP68oscE54O0OKfaHw3+Cy6ZuTuZmOXUJ5N7YynDZqA2UQeZLDJmqAR1r
9j1lXhDCGLbpS1v4tr74Qh2jmg4dHet1q/Nl+cecbHmSnJvB75Scz4es4juE9HX9
6yA7f8ri5RYX6R+um/XCQeUkK9D+i9nrhX0kkV0+d+DYoedAPk2XOAuZ5j51098/
JelBXz2DzsXkLm/KH2GZNj3zUzg90edFZqelI7WNic6RRDaeoRvaKY5Bt+3IVEqD
9TmmoEJzk9ZiCvjxiZ+iY/+OlylQXnrzyDQW4zqlCpl/5zJgJk8ovfnQmzibzbj9
W5yRVSDT6SV2Z0LkmYob6YQ9yOPtGTafag20HjllCk9rliTLxDStz7rF0tzmoRcz
VMuNp6ixC2VPEj+gGbeNaOQXQCnxRrbRuns6jMtTIf766mmonhqI7B2DUl/3RDGA
jPDHJmcFevLn24dnf/T39xE2O8vw4GO3KwV+9ej6zI15ZYLSlgbhTDFmzz2H2m72
b0Z7ys0mRp6kIpf+S9WoQPvOCWd7MET1ixOaFiLCt9bPgHdqyfLpUIfWYBRPji96
Nv3d1YBIdi7eYPdQDb2QUtAESbpxZ6xbS/4H7ttWZU/agzUWDC2FBJSfNml9+llM
xPv3PsKaYbGEKLAg6+exem/sXGoAPfx5e+yatD/bkh9eQKc+OboCKBAcbBE7Euhr
KXcFbAfYSehMJ2/sd1J/2H5hvIzlrwN4ZK8//ndyKc4oeA3YJJrqiMfbSbyOJLP2
JwrwoJNozU9JbF3zwED5AToMZH4ESqnGF4/4G+zp/Ay9HWNoXBl+SA5/aSfE4VWz
p/91Ic/k0UogzsX6JawJI772PhZYmkg9pz3JKtHVMTgTC8s8H6UUeryfrq6q9AJp
UIRv027HbWEfc4sWqzrygwA3/345TXHmSpuDXzs4KNrdlmjNoOcQPI3W10zqNPJG
DryMbakw6IHGNWgcPDxwLd/4awn6SAWMmbb/zEFkP4wcTH7S7dOY8dAVOtdsenXt
BwAFeZhZcfj52xNsYAINBv98bnkjkd1baCnZ6F6rPGTET0hKEdWpdvvJojOFrsHs
2Q5uaX0FxK6J+0dVmcg7tNGDq1sQoRFNqB90Jcb7t5gy0cExGJYw8wv/rq2ywGEU
0iUnhtVs/8mliBJyYfBg9DEvUQk1MfHbX4gGEyNpqxIK3mLI8EehT8ABd9/U5BkB
8AiBP5Jgo7o3sWN4iys8Mmb+xcaD1tpuQNC9hd0sIiDQwZIYGmApsDME1hmBAjFQ
JvTjSkRGiUpES7Hcq+4T1UuvxOTrSubAHWf0v/WiICzMJ3ExrHcyR731JbdH1Dhu
4dZOIDXSkUFvoJc5gjNG0no7+HdBcBmerGK6MEzhCEW3g+i6mt5aYC1wntQfLmMS
25PYcwKZOBOyzv+HzlbFlYitVz8BShBYKlMWNWNXbYYvEWImhe4HWoU2kqhOk15r
N3mXbLUUkg6nHGzP5tb0iNw/reHiTtW70u80iHRO3jwq/ruT9nj0CuOuWljxzn/u
vnPiKNlqn49+ZdgNJ0H+Kt5qFMmcBmt542mIN3ar+uEd/9GmHM5C9IY24vWJ0Isl
Gia59Nf0cJ95ycwRUvw6NPXN4KQY5dEb/9r2YVi2TwFJpC4kcUf3QbuIS+uz3QlV
M3rkpLQMhY6L+jYNv2sMhWsBwQiKfmhz4D1CbaBltJ1tBBA2FNW4QnPk/8881+Gj
a8Li8HASWuPlK6V6lAl75k/EQXrrDQ/x5Hhvk7De2rmUhv7OzRK/H5YAvsqMvmc6
Elrc3tFeluBthwmudy1kIwyFcGvXX6XLznXOZZUPre4gZNAVzcgAM9cyesBaUaeW
nwoMe7/hsIGm0I9PcTJr0pJNfyF9sGN+7YGOCGGhuRGzXSEHpZ0bInTNtGYTgqmc
YNwe9RxnKVer4BvWBge5ZE3Nr5GrdiH3yAvuPXMGSKmXAWP3O3pEuk7RIapjVKkq
S9DWwIqMfqdKPxX8dSEBtwkYihI8q6Xhit2kRZ91zM1ohSwYf8z/GGs7Qt4D1pRK
eyfZcHBozb9G2/FaNERhVSOeBtR/tiL0cCow2vFiDu3CMkyKIO2laLJJ9n3/oupl
3Omr19HUVERaoXnkFYmap/MAy6o0WKGRCbGAf+QkN6WNTNtE+8MfZZpWIRD7vt+A
wWrbbLGR/lzVb6PpIoN/uizDHQAyXt5VavWtpcT33T3BeNpOd/e3iHYz1CjEOJ8N
RliNAW24CnQlA9f2VJ7/pJSZ+l9uHbvKEhyDfwQchXj5mGUBrQoSUNo82CZTYfui
oI1ovh3mebzWI7VeRpqLHZ3dEyLy2BEfcICMNVFkL2CLJmqD/kEEpi/yC4ltXmX9
8UoLzcOm8X5p+Oxf0fJTopJEx5/saGdxL0522bL8W2BtkDiWLi9i8e1a4FSLbZsY
fK8lvrMdlYTI0g2sCuLfKwDl3dLG13lu120hXSsUEK5fNLfwLg327OJ6cmxDyUkB
4kSVKK49j8Uq9OKXzwWrXsPK3JxVjv2/qikxSdULQ36iRjaYfv4pw1tz7qc2PupR
iwDCJnDLSXAIhnWdPl3ulLB3phx72sR9okqK0ElVhZ+X8yfCkHY/EJRF7IzdDLa4
EYUzZG71vOxh3xxQzwvPf27LbSobB4Se1egfZonDhucaoq3372Lx1wbH3shrpTEr
gHzuOgGfMtIzUu5xDFL8wzDoXZStbsbGCalTYysxtzwLCZPaTAYAfH2RUlX4PVMr
z1d6X7DtK2oboS6kewkk9zMYVhkLHa63n2OZogNRN10qiUTbeMmIYi/VfJERc9wY
6A5jI3/fK3FaP3w+bRqA8FowMsH7bvGhCOt5LrMN1AWzij2tx292VA/fv5yS/mDb
pFGtI38RHw4x3LC5iLVfQJtj1mrFtdqcarAo6GW5cZmLucb+nqAGU4nVdOFmYu3/
ECdFx3NpeGk1Xf9AccQVte0so4LNniaTKns7Wy1zBNRrxgBqa9tE+Yv8eFrE5Kzs
NtUmXLQKplI1248hbkDZK3MMNRPqpd8z+XAj3xzNY6hdg7wkulB0SpUkRkomVrcA
p/Fp791PdP/3MXM5xXA7puwmCD9/MxEwFK902yCQrqeBkp9PK8EIwhroWy30ko9z
apO1TY5Sgx006uULbqYyIxe2bfGHcVdNScQaRIXgq/Uq9hYhm7o7JFcBEkXgd5Bw
VNhVsZioN92U0QrZL+tr4aGY8wijTMMH4qWLTj+98NZQQj+nsCZfmcq/F0mUZqp0
proIpkY/oITFi4ofjUf8MJN6SuyH/6L04GaOZsflwRWpxNI6llK6tufDIXpvQb26
FAIIWwFi8RFIHcttZV1TH4sRsreMAvfcM85G+O5K84It3omqEUbzYr/KI9u+fBnN
IytYfn9wmXoBZE1m0lT8OOQ141IbpraSJZLp2E48AmITvh2hWRNJdt0em0zCSmvi
cJ+YSW4YPF5F9sQSwmA90NiL47jfFIIzA9f9fuVit7Os3idEc0m/SXGspWIoIGKM
BVgtu/yrDqa7zXUFTxLOCu3qiVpLX5HHuCX1/T1d39vlrYZWKyLic+QpYBdskqhM
s5hatL5bsrQ5w2paY7VcqesHHZwKoZE/mpRNSHyeB4KyUxwby4Z4kv8aFg/JzCLo
dJQvjqVvKchbgCLS4oL9DXKSXcgtj7qx7ltBqCF2+uLeZv+6mTTf9xU8msEse0nk
Ke/aH609IBwiZxJLPjYJYx9OgahVBHY0w8DCGE32ENx96+me4SHbconpUUSPgTKK
FqMhc7blgaN40n+3NkQ9Q6/HRhEUSS1j4zPm+EgpSKaCVew6JZpc/FYDf919mz6C
EgEQKOMGK5VAvpV1DqFj7CU+4z3JM/dtPbm1ib0hiCWin5Jfjnt4xj4UPLJ9YdcC
LYlVMRYUJDXOxMUxYe1JlOc5FTw5TVSBSFza/FuB8Juowg/kAC5RcIKeRDowF5d0
D+qA2W8nds6E8QMfU6/JxZ6pOeS4dtfN0Qti6iMF0KBuypzFsjg208RhUIZKbFAE
Gc1Mz0BgkFSQIm6+GLPq+XLoQ6CMMJ/IXwZqaPb+d3nGrrN7bi0ajYNgG1xfg+tL
649SpxexMerYjE3DZzDmqtIGZ306kUqvxnHEcPzTs2RN+x/zOiBEflFwNMCIQie4
Qslzm/0VwK6NNXJkA4vYoIqyaGnINVLRORwQgruNB3f7yU+46QNJicH+YrfD2mhm
jLMbxNBiqjyGaWRoKdECRWnfwKzVSeRqf8bCoCjmtPSIzH5aE/Kchd6VSyy1xzO0
CulvIMPkK0zHrs/6USluJvTSqP6vptHteuQ4MsA9IbG8y3Rv/EGGnkAhVFXX/+dI
HQc+K7ZMUjZUmpp1fO11CQtS9ZknarEvo0avbGJOf63eTAU1OwDKGEDsfuZ+BSTr
A5N8WDZmIEQmmUptqmGL1Dh4+23ae6ZhjohqfKQuP2oIXuuH0qRHRVmyCCDU61E9
FQJaLpZ8ItvnuejoFdighATYs/5FmCN1GmFgHzYG/qAAhqrp8c3AlHwnxE2KYTql
FW5GV5+fP6qoJT/QnU3wXgsRlgp+ml9HPf3Xb9z6/tjzhot/aAjLtHbKs9cv8TQC
KNIBnYgGeojQrnxV2B5mybCgXi/p7rvYT2YN+Mcc6Q06MpQvRMBzKpWZL46iDNJh
QNPD7v5dvi1EKc8XdS263Mp6/xlDfkFNVMECC+N+ZV+06+guMRc5Co26uUYykY/8
HTpoa23hhMI/ZZwp8Lz/dghufeuSo3I2++bFuxXwYSZXOoAJdLQQKzBtMmp0Wsb2
Bx5298rZ091FIzj2KrRWKtABq6KuOILhHpY0lPNEk9TEV9NvqQqFdK0z7LiggTHx
bfhf8TQEdjig8wX4wEd6FBXjJiuml3e2SuWMGpXqBg/Bs+AFGR4a590sr+o3BKiq
/uE/8PR7Se5eXPKwgL0GKtgBTpxp5ZLW9MURw15pYTba4+lGKSIaJaVFboNLETVj
NqNgdbS9pvhRnv1IdEiXpIs32hghnC/IP8IMNswZ/D/yf+RrP+mRpdu4vUCNw0zq
jYHVLExLCeHvylJS62IimdrgOvsA45Q+gCu72JnI5Gc=
>>>>>>> main
`protect end_protected