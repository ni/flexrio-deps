`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6848 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
akBpHK9XojjdOyFTP3pOwlSQok4cVoDSkx2RsgHkU203RowL9Jl/PU8YXhReG1JF
xb9w26tJ5hamc0ujJO4YKpfR/atqDHISQE/cfwhexSpCjmXkJr3WMcJJZMAysFbv
FMO5/X5q6gkKdUkHTHwX65lwjbZqDtHQXk9ZjMSDGmVZLLaQiLycTUnIB30DQIQ7
CXzy2GDl1RqRJT46dTzghHxL5zQMWZDfW//PkC8AOtSLXiah4WhxORgsWuxlJ06n
LPUTmuQGihApUIGjWmaTizHVAW4elcThCd5RGglfPa4hLAkvwBThCh1F7AOk06p0
ALcAh6JX+Umwtqa6/MX0ty8a1Q82pKDam8CWq7/qO8iW8k+VUd7Or42+6NRcG3Bx
uX/oH1B2NIVfsuj+yr0U04bwWQZTqKxshnAYeZRYCTLFBKOsCK+YJ44modDAw7I0
cWc7ZzW/jTtASL16pphnSQUgFXkI0WYfE1vaBYxI2sPhT762EqlLfoDwh6j+nuKg
xOysfoZYU4wQgVK2RZLmUTgXv1vXB0Kb4ORt1kCqbuaAZlaRalEzZKyr40LcYEcQ
PovGjv6y0AgFrdzZhSnoi5tD+m8t/GSGaQFPAihkZxBp9pXxm/upIYXjHMaKCses
d4EwNJ+Zo27CmHAWRCHgnCH4wTZu+GBIGvRm60DQhjHhkApf7lsZxgM+9IrdcYgw
P99JPuH6NqIbVbYOHnFRoXY+FQbB9rfXwRXIq3B6pvpSVl11Dmhb39nBUki8FUr5
QjLrqaoT/7A1LCvrJXb1u6C7tb/O7QvBGiMo8K0IBXKSLBkVfvDmy/RCmG53nNHP
zlZk8C7NI++QfuYQYGKF5cozoNq64KMa04J6JoanpeRo09hGBA2KQwmSp44MPlcx
00Tb3Q11lGPdTXLS4ucjh5NkXatpgB7RSAGH+84P4Qxfb8hTxWCGEbRX6kLI5PkC
/Qek9aIodecury0oHTbnAcDBXiBX9TxYjatCzeJMoyhjErw6d0UmGdrmu0TS2aFY
7/lMLqaEgy19T6dajrSuicxXscUyXJ8DMDgh+GCnG75rSyzamS/cpgy7fcnMsWdw
9iF2hC7Z8y67ClYJCyYxs4gBMkb1wc4oWMmBIGe8XauNNgvIHO3chVaJwG/nRRzq
T5ly9ErAdLyz+ktyyt2iiOvtTa5kTKUVFXeBMuKgtD3nADymWwbjtJINionBLciQ
htHgZevoyYBEz/sx+a67yA8mad/DAlWxsHS+DFBopNyrl4fR9RUdzdL3/sRfghgs
X1zd4PQFCKBGzzBUCdslnzlpwYa8vjnaN2k+TNTkoUf1/Qd5nTQPh5BCyWxpaKZG
R2D7WU158iAgV3fbUaw1N5Po9gy4hwSLaTH4DgsNcurXcZXKOAJkOQFn6Eemc1x7
DRloAhLRf4PTpfmCyQasZDR4M9zpq8H4Op1Qm6KXUwYZkfnDPnLv5/kVm+lvGOX0
y5GOoPLWu3UsE0CGjFZcnNolGdzdY3N0i7mj1kPuHjM4x0wk/tnQ8UeVmvzm5S2A
Zg7Dux4ZQVpplifIWCGrJuPtdg1CEwGyXGIpDgMaKOdEr4MxRz2uZKivKWTWon6C
U7Tqx8y7krJ1thWyY4x8JBSvuc2ORY4VkWWUVCCeLK/+yVfJRiKyChSVdMsrA9Ar
nIhQg6tS+Wuum4BGPFiSAtoSk++gRnyUPgXyfbc/QEoedmr0c1KK9kw7FUZLnayB
pqzejscKQRVzGwQ0JMhVYboHNjSh8B+5H9qMUBJ9/CKNTdz5MqNl68V87+QcRwUb
kmJX35GZ5rDSuYNHsuAx6Oi9AC4M2CXGN186n/Zusjt9KeVI6CyJ8vvVV2iVlkGe
k4iLpZj0SVE5BHLJFALrIk7wbDyFEH61r0pdBbSNPfYTjn2zzf7U0my+rdQIhM7X
aT3UM2oOCSfc7ojHkjlb9LGUhf7LcHzdkJQmkVbPiZhxVyk9hBWIvg1ra/fMx/vT
ymGQ+boer73865H4yQkvYTlJI6aUMOlUqUWgz40UNldr0mJ8wsSbjtC7oxyJc7y8
MojMfz2bkDGXxEggINVBldqM/rm7JngYMCW/gIoOvBHIvgDz398Ii6npTSsh8Mhn
Trh2UZXadnLvSkU5fe6orOz0rAndOTrgR9EM84qNcmcnuNuVEkfx+C+/M5WN6Suj
CBRBHiEoY1/9g/RhXnglbU2e2jfznyESPl77d2cRr3FZdN8UN+hc4hL7w1aCSfo1
DiNZoSetmjVrUutePites7YpBGJmwWx4WL7PFxJrc/Hjm61njraQu9NYJjc3JQkA
G2aEStbOhVnDJsLiPfh268tlN2ZU8TP0o+EynHbtS3Jiu80d36AiOj2ycVxElyuz
oMkD9Ym2wkuBH5+uIaAWAUdZgX7snSqs14XIUYSZayKJFPfRUAUBil5POHbFbV3b
xKUJMQkiJ1m5ab6F59olm+xcn7+StQFvduHMdyP+LROZN/YfmO8KjusAdQt0etQn
83EN8udbZ4xhtiSyqRYQIAo7oSG/utZs2aPGuqNlHhxgay8p9l+71wT9SShcagxy
YEJdWRypfuHUmQ4zetlJ1V02O+nNHVgLuMkpGSnQQ5YEQBgl/5KtdpUgCyn/n/iZ
rzM5ZC5aJbyC3wzphJPE96Qo2a1oSdUsoRAoBpZRxmvloDml5m4tbwEqOhXu2hB9
Ui3q7aom670ySM1JHn2Ws/l0eVinbbArjrl3ZlZ/+s8Gl/hky4oDHNL6+cS+lqhu
30g5ip3O3/HG7447+clCI+mDbJXNektxZKm4bEqBWkV+b06YzR82QnWwJUjn3XAm
zRM9jxkeBGdfCrL5sO4VMnGfz0hgzWj7fdJX1F6pJJ3ZrDTjGY9/CmDatOo4c6h1
nlZBPl2xYBnGR4woRcY5nNJ5w00+7sySyjIC3CNqnSWwzz5NHoBRz1tH+R0c4hfP
jxnyrqt97Eo9AwE7Kvn9TCTtbSECZ/2ORApqTk0a6y/HeJrZgJeoYY2OvkzCliFt
U+r+zsVijXduU6+MM5rijPO1aEPDZ4Q3zXndZ8aK0rYy5MvFC9PPytD2ZvLxm5P+
8BNYNMA8DahVpHvxW1L/u4m8xj2wM+xQax1/LWrh8pVQlhUNPxiub97wMWHMpQzF
pjekOLQEfi33IlxFre1H0kKILLDRyR+S+q5Nz2Yr4eJCaECP7EPaooBlb869I6J3
zFCcx4lIE2L9SrlIG5bgK/kBHEQtc1DVKC23BK/3GibQVfWmsS9+xEhESbgcRwbQ
NAHw73MnYcnsreEAInhGs0SU9fBDJSq2XQ1uHyGyn7qrckQvTwjyimZb0lMI71Ie
Vh/di/PZxGz9APYpp2G3Oj35p03koiIlcPARGnz/KlFYR94MqM4RjsSghAJRfaff
vXb6+20fL/rpsJ5o7/PoLYCQQj/9QBnN9u28cgsQOqZZvnjliXWQOoAHRwdDESXC
ebNWsjNkl2wXvgN927upSasOfho2x2u9bqQzqg+gHZZ3H81tlydUgoSPXniluSr0
AcZh3kX8IJnj4sye/l0beHU5C6lUC3t4FeYtxWrwjB256tRro6PSW8gElZWvCFhE
MXMj7pALLykBsJP5Ng6yKN+GT5pPhEKzgenD8zRxiBS+AVKc5tIdIhg6T9H8BEb1
Y6RxFuRG5VwzcAh5fmhlwDHOYnZ/0Asxwto+PV0S9lD4QZafy1BHOD6vixzWbhBM
uj6Q4blcgKyFIwA5ybRX4G1zuhZKYGmyuMbLGbfl8UHG/9ynJmacVT+sWlMclTZs
pI5Rq+kx8gFSoo7LnXzOG9gpHaru8H7Us7370+vv/V3/J8OwlLAuwXSc+Jhmk19U
5bJiJRmfnZUYvaWYBfjPGsvtPX6AOiaV+Ny7/1mpnZ2iK2ycFWxqDCn4xHmKivdt
BnLxRpDnuP0oDp5Zpurt65HzbVSSYwq9+pLawyufNqJGwTH/AOF4w9VDvChRPsbs
bDqtjksYDZBy5zJV0cZAe3IcDhrIgB6geqT4l6BaTXLfQALAm3hapO+aK7OQCRah
8/zOOXovTB7kLZ5maLQoCHtMEiP2XcXkLNBhixf1ePNq7OBapguENRvOjHmMJEwW
tTjAzXWXMwO6SXxVhe1Mmem4ZTWlGMSu3fR3t7vZWb2XclnUNUtFKKW25JBQagV7
PB5jQTRy6A4C2j13+F8wEPpLN9BXWijjjvQfl26FWR49X04hoSckt7HBjfTFzTgY
2Xf4SAH5Xm96GbuLlk9pxutXgN5vTwn3/X6X37WhLgj3mhU3/nWL8Jz3W2j2iVCJ
5cqqXPiqhaSBvcDPGXVVDTt5J5rNE/0HDH3UhpkoLKAn0xDsO0550+58/cIIJFHs
N9AaWgor6QschmTz2xVyRCu0lR7gPXR1IxjEwk5W79HCkOJOk3N4bXRJfA43qeLl
OBIV5sjZ3to/pGKbQ9tiy2NfHetZkhhCF3uyRUZl6SbKwhsr0rpZTbaGBgjM/CcT
WApBHf6/eaJx34pFU8m3AmiDQwbVdaoeUrgvH2xOY+JftsuYiiFjjtstSSCbKQwi
YuuMnmZAIcppvC9QnjIU85QRYBJTYVXT9sKKRmhxuyzN7YAZXXWEJdF5oJvlRp6x
+4yRp6ouwH1vWv7bBBgVkawXeFmTD8MnKgh8m32MB7HvNiCClQqe0DqemnKrTPne
+tzkyHNULj4fqPvW53lMQpAEV1ScDr9uIcwjTawHe/Bmk6Jk0PzbDsHZ5p/jTMNP
lX8uzO3X0HuzcpKNKmtcHFzn85C7r59CFIqKz0KhRJdZ9+i+SUX3M1rkvNllwYqn
9nO5tyUbtgflnm3BZ3YpASBcn/dE3qhjUTubhNdwlCDzpUo6BXoNv3LytWf8cazd
bEWSO8hEJdQE9gp7dIuHakf1QullZOwig0SlIhInd1rzsr6XjHTMGNjiwrmCPsUU
17j9I3ASeQI5iLZk7SJA6FchwuY2f8x1O1RalkwPDJtasfUVBxTt9xvb0uzpIkNp
xZScDgJvor8CZCtKzZZe0s7qc5iRjiQHQxgbZG6vFMkD7XuGpmLqWCXUFn/dIuQI
667LPfUIKz89UpbUg7haoO3IlfUyPHHlzFVXWL0J/Q2htfIlU9Zu9BctK4I/RNBH
G9zMH/T9nLwiX+0+DhTiihJZCYDxoBWI/4zU1kkazq3PIWQQOf0yT+JmBFSkd+Pb
NP5zaKUDD5CnWrTcGPISEzxiIQ+EhJxwsLw2zx2aFFAVSh5NunOOTyKBp1dZFLF+
6cdFeAyUnvfzmwG3gWwlztJ5fO+A3rvo/38SyydNT+AyOne9qj6V9xHT3kO5QA9t
/EjHEtUhROxhAFepxQcNo+wGH34dSiljr3TiBM7yIOJxLZaFdgw0njK3u/fvd5dK
qt2S3nsANuqBi8NiAaO6AvsPY6VjX2YFP8CBjQyRudbr+eR92UjssngjeMlkss0B
ZREmrLR/fi0fz2OqOX6E7kMmNRdtuP/yeJz0ylmw7f4a6E6gj50yPTCczOuimFrA
xpFblSa+vmUqCD7sdQfSRngy/q9rj6X+pVYkYacmx2xVBKNpoNuw15MhZsJ337b+
dDMUr3hRbuSWWg4S7fm4yKiGbyzFpoAfTYwk+4JfFumMZAEqAR85e6YADP9VYbj5
lVCtePGUlsY+CJBiRryTPsYKLIZ/Myy7QwTL6MTKJ/Gjmkcs7orqRon1ViHa+soS
sZHnLBAY5AGi30QXwYgLCxNH080FJVk4wRbrWRX0bFRnPr78Sfo3k13GbhoLiBC/
bwfM17mtdcS4oLpR/lLVxr+cwKO+dve7yMLEb90lfpw164oYopcrLCNWD0DsvT/j
krsjLSwkMElLj1xuwLFnGBtxHYD9OLMpPam6olBj3RicTStWRHmiuAjfGvNN75wN
V1qeXjMB1tPgNMKlGF19pZuAUM8mQEPNNanZRi6GghBE0yc9FdC9LUFEu4HjZH6d
ifrLDa3clzloBvXcOIF66Dt5P1pGjUnY7zEgpaey9ITEkaysWsk8VUect/RhFZNY
uIpklhrOSWkyS/G78sQJRealB0lfaZP5T+d9C+Ui9ds1JBRmCsJJPUHd99m6UX9/
pomwzN5CnIZlkwhbzIDOSB9tuBSEpGMFTyAicycWRKHWyQnZvTP7+gvGO3ASOhmP
Ie4ezecSl6LWTjCCOKlpuIxdtHsuonsvhlbnz0HLic4msaFyIq8scHOjP7qam2KL
UmkJgMywirRbPP4zEh+An73dT+Hox5D6SZaUL8zjk9PR1thMjmYhCM9xjwlUAikI
ofWeY0eZS0WEQmxXNe+ylyG+AsQMFPXLtwqt4UQb4626T6SvKel5laIni1CDHPAQ
cBM4iYvi+FWapOs6u0Ox5pM0lFN2GhvXHTbdcoSYCq01EVmHw85uhLgedOgY/AJo
xL5HJM3I84ZsXDNC09EjCjJKV4nVjAxKl346iSEz9b0VGBJt+YvlqeXBtdSZgM+k
B96QvMUeI5/GGP8ymmGcQ5HQKmKTveJsrUQYPq7X7v82mEoOsfOxWJAcYpQq1iL9
m+ngfq33oicmDrYDkOsINp+c4Zaqwi0DyJXmEvNYCEOrEZYowPKdtKf4NRz/v8gf
txoNVzdGCJDsvDGSkNzc91MLUxQr/IOsX9w0UEBeUKKB/QexXwxYOaqL58iKXrtu
67If6llgVPKXFakfmSAbv3HZmHM5vCGrt23ZGAIU2rAt3IfE/TuLScStrPMpDjuo
tvACrEFp0uIoyygkGlzTtUIoFOT95asqLcieh+ezM2KS/Vp7tAOSMqubL5Gq4S1A
Z4nq9NGACqm1P5vgB4tmprQWhXCGu60nXduVmUgFmLPbtTJPbEWLcqxe5FZaGyxP
1A3E3F8D3+aK5k3QNYW4a6fTe5RabiVoJ+mqI00j0OaZ6+nGlHKy9DfXX/wel+ub
K/alZ7a0Y+dWwAx80KAU+VnYeLR0CZXydk3R3YPdihoJDBUx8gz91TTB/XW9e4um
jrDLQJezs3mQXWUehQIY1+73rmfTzZhIhYOZ0Bj/6uxaZimDDd38P/B1qxx0kgxO
X06IeeqLx/1gaqe7bHUqzMOh/uKX25wkMDvwjRkYJGGhI2n54aL1oucComKIFYV2
Dw9bOYENddcGubId8fhOT0W4uFzO16zctUdTDfeSXHnNptH2EO+WDgQPk4e+SC6C
tKDBIicDz0sq3BXfx9FxoPHGy71iJW0CmbiKVUYYFYEby3o7tZZKzSc49vCyiyft
CS1dpxg+tqBWBDHLSm8/R7WHJPnJul4HiU0cGXSBi3U2gDvpENFDCLfRIS9iqcLD
R+UF+cqKUavKD2hrjoDLNrqFLsLT2Rcgpms7pVQOAbejcVU3X+lU0OYiRMWnQvRL
WADarzA5SiCYqFs7VWcR/LhNJYVtc9N5oPoBwma3v8qyG/2EehNKgibRizMU+C7k
jDdUyNsENn3d2+ZiWipsf1Ld9CvzMaKEAk/PYHuTCY3mUsTr181ycdTdiWPAP28M
WH9niZIMYWIvrYKV1Iz3EKKSLiUS3/8jYm4hqTnSBVUa1xZbAO2mcQ6nR+tl/NdH
brWW9tD/YFRuob//gLhjmIdgMK8ulify03aonp1Pts9kSOs0DG5nDsURhi3FSvAr
E5fGtQotkTeUyU/ZXtRGeVQRGgVqBYK8MdfKZoKiP6FGmXi7/sBXZd7ioH4eLvHy
uItnBNQ9ja8woauI+1nUMZqqr6OekWtaOkOXVtic4sY4R39zeTlUJnBzTZONIZSw
BxuM83qI8Lo8hOKBXIGR914y1vdPsImFj/t8/4aMWfAUPyGILwpi3JlKUWKPnz2/
GEkh3H5wZLW/zB/opEMtFHkg7BSANY11ITolxt2I6Wq0S5ySmrJSL/Zga6z6Gnj6
1/Sd0BQeoV+K5nz0ha9NzgAdPv2GEuCoSZVn6mb7Eoj7zPXQJdQF87LPNQb0M1FE
+QM8CJiulbpCKcNwlPFj3AuJPX9cGpMdzTPNJwzRLQl++xhlnSdiJ90mqBvuri3k
w+y8SCIrvOHsjLWl9OAdpYkRf2OIIQxdYQGMOlXVpkw2k6xlhh8R1vDq6cRc8Zos
C80+lxGWMpMFWB6Kz+HzPaqUVBvm8lcnLO4JLefCmqz+zp355WGVDqmRIfLFTGUd
EPmvxjsuJSYg8D2NrwYhnfH/MxoLMWC7dJKBicle5zIDoq72yQEmOPaZbVqGtO/5
rFQjk5uSqoufzIEgVGPvzMwe7+bW71qipFaQd0ObfMnNKsNJFXzc03uj05i/9VjK
nF2Gm0zHz6ENGSEBz7Ffdm9fiivWmZFeRQaihxQRcC91dVRfyNadI8cJKSZhVBG4
Vj/z/GZuy6PvgYvt/FdniU93geHalk/KPXzPE3l/cdEPYVndmM9T4WIoEYr9M9JX
Ct5150FJPSssRc7Uk95pn90IBztLviWL6P9dXwQEXkLBpWsgFCR9kLe+1qKpX4Q4
0rE+2sjboZA64Wt0TlGRM+stX6SovwQI0Xc4h5TrYPvLPCVCPoEHKASD+O7Rjyzf
7vrH6917nSUU8uu1ztZB35Bkp02c5qYjt90VGm+aST/Dh2C/fkvsxju7s8uxV/bJ
0PekA0C20TzSmgfAJ0GFjSlN1gGCPGVATVHWtgc7UjJVBzHiCPZv4n09BxjbHfAH
0YZRLexS5QsZCrUdwn1Q3B5EGXXd5ZFvw5sDa8Wdvkc5dlm8PW/iMv5cDfxKBYxc
mxHgqdcd8qjhOIii0euHZKHJRdSrywEumxAFDTsaFZQNGGS05hQmNuj9+peA+h4W
8XsdmOz1Va6ngZ+wKgiJwBj66VjzP7RbcS8kXfOtqvsyhYnQMcL7LQd0BSEGVdmV
F+LpG4R69zxxcxJxo2mdtiZPE4xh5WUoeoo03BcSnpcsZaMQV1kqy56qitK3LBMf
oBMIX4eQZugVTylMw9TM84aeDe+8en/ippm5Fz0moY/hZXP83yup4NS18+dEAXbr
9i/q5nyFZyTAa02mZ0EzZrqj2XfXLkuPEU91E5UvYfE=
`protect end_protected