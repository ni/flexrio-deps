`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 33072 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
rC6KPz1bEhpOMfeLdNDaqGez57ZdAnh6/STrMHN8m4d0k4pgnoDvtveoWYivBJf7
tUtQ7H4WsSDJWnpyYtwfVcYWE+UMW4TyWjvJz62z3QeAsUvOlTBX7aXLT+vsGKww
kS5Y5VwGG5cftZ0cwKTMYY4ZvNQaTaBYXD2CNc0Qji3foEOQL08XuTbbHquMh02J
ju8ttVS6hUPgrGZFx18l2WGrVNmYWdU2m/XncCBzGrEoLtkaer74FDFpkwzj9ZyL
CavMjSg6mSRseFnWSgUM9WMemZqG1LfvlTaLCpw46snaGBKWGgxGmuxLwV+A2sHe
ZBbmyqYGIPEWpAnAg6rEHVbvTsWwDrkKBrkD88/Domw8VafSTa9YFGryMgASmCiz
esKRGkKusf85Mb/SUaxIiDvAxShMyk5RXE1eFoURegYqJjPjGQoy4DLkSbaDPYfq
H7b7Jrc2eLFwNzz1aAJleu15z2buNUOzDA16fZWxX1mQk11MBumcI+5NyHI/whhG
BsnVsrkn4E/sra6vH+EPxKdxLdfBK5mJI5KVGd8NTkNzb15qR4YUzFfWz/eXg0kw
fDwZM/CeWkY8KNP5iqNtRjOGqvLr+XS3jeZh069EtzkZRgdlCP6GIjN8rBJozmsy
POZt8boAGT2mF8aOffWEZFkqRFL5wz9g35rbYfPPVA7em4u2bEYgQnTXplUEArI4
BmEmpfNVynHjogKkk5ysxM32MC2BhN13FJyjkEX+sNZpgLSzHyBQWS3C37eSo8Jr
GjrrNeQMRZoAzZihGLJw5mXy27/GGVVZiWQ04Ytcli+EOkKt8RQ+jZT9PMSZ7jZM
llc+I5eDLFTnnT4j/NyUBa0U5oiv0AG+DEw8vhPeDXhkIjh67vTJHEFLNPcOFU9Y
9jr1P++WIxCIsUgHhegiicRecuBEMnP8Q2lHKrd6FbfjF1z6AE0ebhSuQITjShxE
2am4oH4F0i1cOpeKWVvJ6z4zO78/r6p7m7qkrucFIWscPmC5FfXr1Z3NksT8uVNn
gQSABgtchDHIldszQEyHn7k0bWvGrzxVLzJAAVNeNKJoCf2OhRrBq1JvpZPsRWdt
ydQ/nKTJodSGHP5sqJkrubpojt28lZWUcA3e3u49MRnPh8hVMZb+ky9bi4rCwkFv
Ouq6K0k0Bi6HdXEU2BfJU30YJ7C4cjCo2R/2bjlY4MKkWEZRKHsSv455N0MkiP6z
VHq3TUUKqCqoU/AhDg6s7JPEGQBlIC6iFzQniILqU1wIXA6Z+k7btp/fjBMiPCEq
W1M3oq3tnmzNdUbmW7JIlqg/DZblJeZ2LkTRqihhCmaQkV5pafkfpQe9JkrSYpEv
ifE/HwPxkLqmytoHatNbyh3KWgMicNzTbpog5iG/ycf5ZyOhX3y/Mav2WW3SoDyW
42HlvskQpf0FTMmKPb2brM2e76AdvIaW2P123JPEBS334Mcw6kJMRHhoTcjz6lKb
4K0MVgFrIvK+3gDJGx23YGcre/veHCsw/2nzwW3JLWwbpxTWcxD18H9Uq426Da7c
EikM5h/DFw1vuQAA1UiJh4LB3Cqd7oEIYBF6QIprcSg5TwrJzLxIZKKVf9nPGOjk
dk9K1P2fG2PvGXGtezfU5r9W94QlYsGaiuHvIVmG3F8Yai41idFFkwVa6Tt0JkQG
PnemAwVO8zExfsz4HiulgwpjBMGJ/eek4xdu7lWXXWOKA6TGq40tYo6G+x1GVXAa
N1adVEEzTq/86t48WvfdkBurCjZbYAeMw1a76z5aU7N+wgXVqSQPEGgXQQhIvzU7
8iDjUAFlfQFs9swSnaPAjD4ne+NgB50pbP02KFM9PXNFOzR15OSfNk5xFRbr5Wwh
uZ6NyuMZMW9GAuVFpiGjwRvMLLdpGs+XhMvX03U8S4LLYrhubqJuBzZOsKmavxtX
UVaIDZ67f7vcqIwWWSsQe70NOpqeau3gebM0Lgmhh9TTIfq1+d9JKgDjVsef4isH
B+dP8jVbUw0EuVPC/KluZi9ncicOjgfztl1+eFPvB7r/zknM5vCi2Dei28lfQUyj
Atx42wgYB7do7cT8lE0chL7Zyav5fjb7jn3l+w/OkHX5KH/uRFd+Db6qVd1k9Tmi
gjG3JPSgtNNmtQNCfw3GGwahgJ96qFrXoEboJAGk3XnCd08vFBlvonYAIJg8ZEcs
S6xUiLQeJ445ODw4jZcB7tC/iKDR5sYk2Qt6cK+82ieatERlqP823iJ0Z6tLLUHB
7tFihR/qviW6hYg1G0BFWMUGFqKBxia45sd9BY4yfhvrpTZtJR8RX4oHFkjIz+aJ
lnBKQhSS1XHnM1spene2ErlPpMRMyRf0Y9rQ6ZoWdDC4snrBf7MMM8KFrmzJj1Ix
m7SyKs75AaHOELxqMWJN/8Ld0QN/XgbqjBUrsvPCm9g/avJexqO9PVvvxFJA3XXa
dLyiUHm1N4Y6Cw98f5WR8pT24u2VhTHxkCtGcIfQ402NsnTefU3ceIU5TuUdzux9
j5n2lnYzVcW35hwr6rJ1KjTAL6zkad9ckPilzKw4+gHNjfgeoPo93rEwmFtkFyWD
hnJs/sdnOM8ZKQYke5dXGXgNRCM/Th/aD2DH7CyzHt3aWDD2pDIuHHypQDcw6t+h
JJOytiCKdStrjhLwaE6amzwMSpaikfds01dPG1lYlXzDxea5SWiKtqOPdn3dr3WD
H9FNMAiDLymeyVFVyx0aAHW5JboJ0mVbV7J9FvVu4MebRPN7e3vIJb0cBTtTExFW
g0iF2BAGZzpwF3W/WmQ6N2rDaovjCVidNysgwQ16AWRTszkm7oGU4WSGAkvqR4l/
EtNXwDptMvw+c1nn9brMasfT1UW6REZNfRDJUvJa6jK9AopvWNMi+tducM/RWd6U
cXTR1am6BpYsHQ4fe6/FtaZ76eaYF4KGXVMOA2EjL2+LFeXMKn721gX+usCSyrFc
balSWL4OkXsC5qtd9vK3qP+aaV44EM8j9E8J13SGnyQy9K7VSWS5GulDnTayDwz+
PN50nY/+SsbT9jR6rgFlpZSGRde4YFrH97Mg9saRg6JXUxdgPF7Fygl835jLTmPH
MaiY+h5O454jsqsx9ZqK3Ir1ppIffmLEIghJDBy/8qGvLL6D6CXb9WIDi8UWit9W
xfzTx33az5I4RgFOr0A+x2at2JliliVQs9e+ohabipADqN9ZkVfBIBwb8FPqa2Zc
aHCaG1epVWa8ND/OUpcpTu94Ny70Kbr76qrwMEQWDvEdmJfPsmBwTFBUoGb8kSbr
vMcGKIm2x/bBLc/DqPOPX1V3yN7rm1Y05SG84QmHRqng1+Z/wwleyL7+QIC2JTX4
pePHh/HN6QlhookWPL0/xP61e+O42biIbsE4sx5YZWGoOvVZ92UhuiI1Ccn9RiTV
1/Y8JvJHaPD7n9AQQLVqIpYfzdmZfI1BoVOCxCUb07baAJU2BNFyHeHhr3Z/giNt
/CBedfm1lRXa/NSS1qujPM3gTQNc7CkKOTqRJ7Q3qLRq+CIN1Yh2nrVTmqxRvvMz
rFKf0wrx2ljVJy9jW6R9poCAIdhr5qSEGqVzRCIpKityTJHKmWIVpjoEWgnDyD8P
SwfkRk85RoprYZUCuj3vMPtfol/w5p5vWbKq0whU8MHH4tvUd487lfcZBrn1FuJl
CanDhO+bBrdpxlyVZcEy9uEXEtTejnOadSN0qXibYehbFtJX0vkFT/qAe8Oav8WJ
/D6AP/NrzpO5xlKg7b6svacyOtvchlq1K0Xo9l8EajfUUgvx8wQoVqTyOYg2KF2h
YWbGXLvevzZhJWZao4svjD3Ozxzafyu5dm0YKRVSy/8aGXLqLCJ6nv1adyQSgWMJ
81mlrzcU7wZBIqYBR8cNZhT9qBdbgVUy1mfJBaF7WIZ+c6AO9c3c87LfssNhes7p
SyD+/0v60gwK8vxsho61naO/86QtZHtE4pjkdPOvQjSLlZoiFSFY7JJkqAP8rSBC
amyNC/D7VX8xFegK8HWjI5k0DSsR/FOFeyV0cO37ww/UjNxexo7L75ZrpF5pl5G/
rPvgK8qFWwBqAWIrMrDmCwzSM7sCnKuuhYkhN61+KF2zuZL2IPQJl1rUxdb3Ga29
Li9VjeAXzkcdKp4Fa3eXBJSCx27JJDEzZt3ogE/tNC/R41G9Fctkby3H2dY60w3C
1jZ6DWH4xrnhIuZzgIXItklYRZ/AaFkheClCPiB3DcL5WmF5QKenqGMi60W28RXo
+lkHPHQpEVZU54Hn0cU5/bP3XW6vGH6EjA3RTLGf6tNSItjwodyeUTphCobZdw0Y
dnPuFHf5SVLRDA0E2yrz8PpJL0Uj/Ir7AGVbknBUIWaST9fjtOjnnJYa0MqVkVo1
0BZjStDs9um9r0guMWm5y9D3cWLM41aOZaPbWj3+krM5dFxJ7QRdSczzGEnTySxK
d8VGN6uY8JfAAlIJ1RiTXClboPYgAJOhGtbkrs828e1MwJOCZtsm2sF5F5p8ZoJh
NaKx9e/rjZzz++Hye3XWRxJaNOhCNpxjr8i46bV+1ysCyMcMK1JFAlzycTLSG4BO
n9wIvECDeI4bKJTuBCw6u47nAVEVpnQwrmHwa7j76aJeipDTRn3HitZzouaC1Kgs
HkDeFGgEQwHDRJaBv28D4oGgYdeTr6fztpiNL7+qJtdeLpim519aS12vPxorq5nN
TeX2Yd2B4+Mcj7qdlnfdC9l6ytHsQNy+P2RfD79EtFEKdRPui1IDmWQ11b8d1A4R
Rtk28SsuObgxu+tq51BvNj5LlS0HGEEcD8ZEBdekAjYXhXuNtYZ/O5uRXBWlfUBa
LQTe8DdsWp6HZKUI2xbIjngKMdU3HNRW3lE1w5xFg//0zxN61Sbz2khqlj4aBIKp
ad2y9fxuys+Yiv66XjMHke5UkFkCSYF0zo7OGt6yC2uGIMSwFYaEQ7uVeA2X20/E
LTY0T1JSrVgpLduSdwjSW4MQmOWBhTaLoFHEg1cVpGTgIKzbXUnQzSjkAzv/RpHr
B04ShISu2VdLagdgNO1kICfppRf7tR9zwTRXEoUc2YhMipquaTYy1wUuv3qRoRAD
xNmytcrsx+wEnVEweGGm+jzQM/ahZ2wRkqqh7HV8JopT5Wz+h/uCxsyuwPamNLJ6
MWCiNU/Tdp8WVtbpPZqpyf0mQU5QP7UEKdpmhU8Ez4khrJY9BFrb8vmE7cwi1Rnh
6icZvFAs+b7E7CBmw7Kpk/uPS7yUzz7Ke4quESyPEca5/mbxbn1YrL7/07cV22WW
yYgA5YmnA2MNydCRTxZStdyrimjZ+Qo7VFVLzn6Exp8EUurs8XK7Gnf+XRolzozb
KVBuWyRy9wHAl23BENYoCPaF8BjETWdanxsmjuBabz2CUlQltFOX2Rebd6TeaASw
i3Ie5/JkCcX9ooUeHpuNwxYnbMKesIw8rYhGFoCkDLpkvgG5XbjXDBXgvU1CE0DR
uNeVIktoUybo8txltQYFbwJ63ahi5m2Jes/u/gzztymUKMwfbMbWRSsF5DQPXiOG
Q3v0yDMV24tXLSrDmOgzaqfVOQID1/IXt6Mimn5Nlpk1RD45eDXywoVEA4cHTChs
neeijEkFaZcEEIdvTvdM4WTfTcclAJVhiD41YJTZTaLUjCKUtC0lTTCRtmWSm1uL
c1FUDCigtbjUprCmbkRknwDnGGEcfcgoziP7WTBGArp0WTG2zVyfd/kNUaYdfyJC
h6Kly/vBhIiWwPvUt6klra/9X5Tn1EMZbpJSaXM4OORFSJzIECekzu0fUr0b1xre
ojXsSyysnkLQwYiv3cEr0m+7qR+hVQMj4B9v5h6yALBPYUfavI4SfG7LVNXQqrbT
pEdRVDZ91iojKj5aq3l/bpLHrzK3xVp+4zExc//OX7Q2M3RcOXK5OH8oyp8eY+Sb
bju0sF/3TLwshkcOwfLdMaMK4VD20Ow6v2DMEtQx1Kqry48X8m5NT88qfDO3OLcN
MEvOu2xjA0bLOajJTODFkhVjcjSgxOk9hRBbWEyarHUauHXLKvg9DvzAlscp41Mp
PUX9fcbyeKHi7Ko8QaqYNtVyjuvAptlL9ICnnt7uezgkqkZjEjEj3Wx1vYR7pn2T
QxZl3Mya0wtBYcwjwlL531sbAKZxtniQ1cmjHmP930kUF5VU1E7fmV3OY0sTTcZd
dS6IFKOzmzKx+AvVSm+WEC/inBeO1t9w7LGgBwd3Xa8U+SqmcohisquR/OvlGDcj
nV5srsRtSf4BJ6haTlLv5bPgyWlfX1nE6cBSjpRRZK090DNvJ6rUtgkM2+Qw7ZdG
4Y8s+1wFSBEI5wocKF16RsyuIWS2xxamytzY37y9pUoIUlCbIyKdB2oVfddfcZFQ
xSmcQ5gzOHq3jEFs2xO9MPTRdrRxkcN1PRgDdp8Dmsdw3rrmavYMJm3/xXGqoMux
QsIME6fAahPkPo7Vcc2ptfjW0dOfAcxvmBx2JDPCfnRJfLwejvkiLk+qS8Ecw0Y8
fDbAjdZYXPpIWJRT4oVl55LLQMiRAjtwFuBYAzOYVTCsQnJhc38HysjIHuv6cGae
u974lqKwGcuHXuKwuKuEMMTagjYRjV5wJoHUx1z4DCtJxftMr/kUOSew1JU58dP5
Si2zr85xA418CS7TdzTH5snRBLb/Wa5SBwwh4sHImPXbbKHO9fMCJNX5dkoLnp0k
McFhC4n66x+oNO9McNnEiG6mxO1uQeumc3BNJSD1xJaSLkRhVwiunNvZKx+hsKlJ
Zuh0J4ulehcCkuk4dO5gM7tquYH/V78wz+3tGcUoc9RQ+23jYJSAL/97EtZFQWHQ
BE/xmYvCyR484OWbK4fyQvazICv/dAgeaDFubqG9Z3F10vITmVCM/FElOwLiEgai
1pZAgrh0ZcVO2gylggKl3Ay9CvXaceBK3eBBfeWxTZLZ86l++VD8XAL2c9k4uGi3
U4dVMJEQ8RKokCeb/YsrlsigPFiHatgf4Nuvkwzn+zcSUa3O0buGUs4w4TqNOTJb
3TYC6vWTaUUnEAV7I6GUW1NndIuBZT/rJ+6GAspMRHDJSCCBareDy2ESJFRQlZI5
sseZZB4tO7bhvRJjUGNAlAMquHWmSppWtDEPbeqiEGYM7WjmmJ0t0osw33oQYBiY
e5UBXKQxNRBNM+o+9j21jm4OqwphloVk/00neBypQhNJ4k1eTgZfzEFRJQ8EbcQS
5rz95hFlKekox6d6HuGmcwXuYgfnDYpsY0LNnAYS2+VCGGkeiga8Jbd7DB3qFBiT
zXVzOUWGygTU7moQKhlgH4b7q+BoOPvvaX2bsBxkncUnzO2eEYcle7EjnWbHpHtZ
OTXkP7db2lgZc3r4gIpjXvSk6yXKHHvwlwJdm80arajhHRQetmw3sxbjxidlMQzS
1baPcGOKaEELPx57TktK+v307KbdPZmOHf2FOSDxKnHycZUkc+FIxIJTsOj6bgMj
QNZWfC04TDZ+zvoXfL/BowBgW5x86hky3Uo4OgE0fe48xq6Cl4ayCA1fUuKD/UsV
lbS8LPMYd66YGnDBm2uPZmkHQ7cgoauwrrRRASf9GDAQB2laWiSCTVw8NiIrjLpC
H2GQp0tDd5vrSUgvbi68kDvnks6FhlMWL2k05wSTvUw8E9KG02cGIUnucfFvHO/W
S2qkJfb5BeC0tiwOvQglqKbmiSfYTa1TttoLrxy+JBpz/stEhEU9n18DfpoI6w7U
KdAG0Gq4fROI8q9s1uyqBz3WY+FRTBNPQ1WORbfCCOny6LASRh9SlKRWRBTdHT3M
t9bLwR7ye2G1IjGo/lFZLQr92GCOV3FvgxNmU1YMsYkvwI26BOmV23BTujScSeK3
PSFcFeX7Ca4ZKwzyDRwvarkNLVVlgY6UmnwGlSay/QEyDXsdVwTJxIVYggwFOrsQ
JDkqiOHxqxl/293COIKPaVDpgadd2upjn7GhDMMT7U6nVXWqs4PYMUfxM3Xoepei
KpKjKfa41CT/ayISlGKZ2irkMwexc6wUdKwlV7BZDrlUxxZzaPGGd1/DHY8Tr35p
0dhEXfkC4IuO/OD/HElBHC/5NwXKucH7m8XTQpVsz0DH4Hx0MqrD8XCxm1HizzNw
+wJvCqmLqxDji26NWFX+lvgyhDNLboGvZSjDG6gBKDvwMMCzjUyHV920d3PGR4no
hJTeqiDj9qtrwf9WlCCPQVHQFrg2UaFusgukUZ4yn0e4xApSdiM6nfwD3t5hAxCw
Hsyhn2jxeuJbmAuH4+n6q4VFWhfw1BfmNdhCi09RvenHNg8BrZSHR+coDAH+CmRG
4vkITc98UKVqNlvfzCXP1nqZF/a6PMPLEk9pfAxvu3OEH714Sia9i4U3OpeRek+A
LXwJik/TZBv++T5rctyhhd6O8umbc1iKgOT0DEEHePuxd5UuCnUPxXp3FMvBK4V/
Q9G1mCgF3XMd2AiUEmPJJ/9GVM4TK7HcCan0KR/eHGrNGkCxJ84MplvSQdtvk7OB
LjMgbymc6y6YQ1uhu6mIPjft2jUIbq+1YWKK4nvac4ds4SHKJQG2WerSQFmjKStO
1URkvAl1bujTpCQPORhzBdPV/oIrZ+jSahHyiwcAGuXvd/d11p84Q0S1+EMy+REJ
Pp3wYYUSOnJUrb2oSa/ihyl3K7cdLFw/2V2acWcJhvGrQeWaenIW6BI9hO+K+Old
bL2ARRVdB3W5X0VEyPz2nATezQjwKWfEMyqBahAVG0Y/eK5YIq8LR64aFCwrsFIh
sB/dlzDOSRLjWE3e9qHslO7FAQE9Hn7H5QYiZuC91yIfYDl2X/Wwt2/BXl+wn0v8
WuqN8IJAjPuHd6B+f82aP+Fk4GxjV11UBQn54y6gck8ifK86dbv3lvLB8++Qluxv
+D+9bB0uTfQ+g0e1ELWsX2cqmZt8xni1EjLjMmXSIzcZU4aPFhT55FKPN8vfBVDN
6Y87Y8/UhLlbjyTk/3dkHUGD0hsgpqprRTB6Q6+dWGE5iRxG3oPscUK5zxQdsiAQ
a3XZgf36UaqP9Cilgzmaca9E/90A6uRgelcjl8ZaPfO0QNQsEeOGBRBnTUuWc8pI
JoSvM/hFN7gIP5/ihe3ehLGuwqL9ouAex+6qdMDrnZkXZ75mT+bl2lPBEESN3vkZ
vnKbptyLojjLr8qCZQaD8sPv86geS/GIHt2h67RIEGxFNFUm1cKR/bvTiANgkkt0
BeoPbXgZL/gsD+lhTL/0h8eUv/1NTWS/QORzid8BDtkOIIF/+I8UP1hXePSh1ENK
eKa/4Ps2H2hJEPwwZixyHK05vxcSbJK1e8p9tpcQNVPyQyL5k36EYCaSC1uIUXps
RgVSUlrYcSFQIj1ubpc4Nvue4QPrgxkE+bBOidgDIXKpltBRptjBXfbN06lg8P9P
XiOk6SjlgoMKTKrn6dMn4iAewHetDzY0EeBc26FO7lAgQMEDB+U5gXDM0GX3jwd0
X4EbrUZnEA9ImcXdUynvmfK4kFADgNBZPg5RgEMwVlJ2heK792uHGbCLIvffHBuA
M/sdFsb46XFAD0/1bKI46G0Ri9F2J8J6A2f7b8L/QvHVMUHEtCHFfEx4FZSFn4km
QxpFk5RIem2QopXTNrSeohXDTGJjnQRlWpDxKs1n3uV2BG8PgpJ7b55ZnpYCY99r
gzFOP7+1lU/eyynn1kkSGN+rNtXE0Y6qQl0JBH2PEO6jpyKJA1BKRM25blQuOVjb
8HOceXgE+/K5kqcwUgIqC5AgXOA7DPFoMhBL9XKLwPtdyD++3ayftzWd91I/MNPj
gUtOuiBUlpb2ot+seGJ8LF/xCWM02sl2fxLa7Pz7hPy9yXSIODj6ueXOP5LS8Gen
czo4rWX8xvD2HytY++jFRoByPP+pxhftRQjLD213XKHntBUjc7zNjNYUXzPjih/w
OUr6mso1P7NCRZw37LvikjbPc+uI3D2V5Vp8rMQdBV0b1+dsGuFllKcRwMIuKWWa
zxfmKHcBeH+BJ2tVCBrNKOFwysF1UlOvB7tG1kZNGQd3pdDmSg73in8rTXaVIU/+
zXiXNTRnHhvNscAd5dBvXrb8YivRAeqe5p+iwunk3ycowYQ46zbAIhQGvkqXalIT
2+ZJ7ChVm0Ihu4V4TrZl5LLFPQQzZUp1ApF/hoOvwObzdamkJHJ1D26+cp6kafch
2BJqNAvAsYe4gvgWKNrMlQRiq6+dsRODkHwxtm5ky1SED1ULh/YddsV/Zuo5fDPE
HQ0KAmOKJT1aBb+jqS6fL8ZVcXYTtc7FgePHgE0GiGxpxcrnm/iUxgO/9D7M84u4
VRXLRjDf/MKx1P4gCbyMYw8cDuG0isITsfzm2LwFxWsRPm8s5ZDF78/6npVvinko
0nypgCbdHlm1fXN+gluNnpbcs2BkLHukxAfEo9Qtar6N7HKWK9Lr/PmZFYNJkVbK
pOt6vOaHcl3PYiDV/e+pYDULi8Bk5v7XP6GoIanXOdJoRF65J/iXW7/NR/FAQENI
j2N+aggm9YssQLpyn9aloiesKDhoEksSqcw9F26loVipIR1fxWhzupnbPuMfb6WI
uSBmk4GbzWT2HyTEjUgYKBpBdUUfEKFjVCzTMFCNXb7sPDZp6dRqxPMpjQFn7m5R
zHYhagIt4JhS9uAsgEtAw3+a1UuY6yVwCHrL2qsBPl8k9lwuxo5hvIiIZ31W74AU
nBmG/RaC/BmMMtGhVr3G6r5oYefg8jwAGrxma6QKiueRUsr/s6vK3PIonNJXT2rX
KylYNWpZ9ie2lzBGVLKmNYnDURyfFkX8pfBZKeZMVDWteSHAo3wzuiXPtVeeGdut
x9XGdbE5+pXoPNZbzPWgTujef7tMFY+5EwQ9DCZvPncsFpue04e3LFTHOC/JuNx4
qlaxEZJAfNMzHuyxjh5Vea8M2QfvVLFvCzCwbcFmEsps3RE7CMjTbuZPPJ0HvNMD
2oDqbjCiDOJ+a8TlKrtNOLup2WZ7lvH/wbXnMWragoCc26FDUjnk3mM2S36FTVYg
B8r2BYA4RbvnOZbUFe9dTQlSk3ALYlZt/eeaE+wEKXbdaz7HqnuQALIbzsh9qARo
QakmtlGINEHzxJV3lM6RqdJLiiRqNBWw/b1uPukoOhueRbxsOmu1pC+7FeGqNMBs
q6f2fhedIC/Eqhc0qnwKGNojHTZ7iJ71hFiNtdeD8c3fyNvaOqZxEgY/M/kn1s2I
/ViTiAMTdXvBfS+0fcQQo2AK70O+fE03ls6j9Tc2gFHUMvGFfe/HCs0Mvg20kOJR
bDPaC6f/o/FifTYTRmoApsbvc7tvvEFzO8X+TrC/mpaCgk3Jfejf+H+2PetIPGIC
UPhsOQ7aNZPJF8Sd3PFQWJpFEoAyP9z3Kbf0Qw5hTE7xq93096PEK9NrO8Wz8M+j
bXufP2o1xytJzpfYmIi9XpJgrvVVAogockvFusVaRmCjanxXZQPAGeKB5OptU4Bg
9sj8gz6So3t8NPruD9ySiGPN5ac4/Hsy78kEZiZOO8GpiNHWxo/C3L1yv/6iFJfm
5LDhVPceZQjz96Na4i8ZGKc79rwWcxDcK1JNOk1Tl7FrSn/wC4OI/WsnsRftKKKa
C5R+QeP4fvifsIP+zYHte20sl4bWFNQ0mrN5PmwF/klEHi9Sj7tMZva0qcgG8j9p
Yg1YLhB6D1INq6XYWPL2UVF05ohbKynTrGul1wPJ8I+0PDrQjnXiUwpkntfU3ci+
2aH8mLGtxU+LvEEdm8j5HQi215G5oKtC3P/B3td/t0AFQYCE9es9MAE0+i7Bbupv
Qaq2tXcZgqdE/jusMYQzuiJ1+Q1TBRrHC/I9Kk+kj44XvCSG30XrOeTdBIT0mQl0
VBvaWSxeQoze41Z2y3kE4kkM0NCderCizWbXwzTHNrIvnACfo/k9rf+Ow7UK7AVT
xyUeglXUIHsUPNqHRCDn23tKGPOHJ2qjXwaxMCyXlzQGxCcUmUCTy/rNnj+KAlmo
CnGyRgyBZGkkYNf0NMwnhuiPj3ejHrneSRmCSXs+lmH8FbsrXfiZPRfy0/Vyde0T
TOJ3BqaLF53V/cqCkvpK5vSn4M2F3w2nixYEUXRyAXilKVkvYPXIP+wgrQuJi12m
F940J5Ur7yn20taQBDbr+0tGGnuejJ5238KdLt1/ShqXURyUvWdC2xStLm7At3H1
s7mYthGUU+qM7d19Aibpc0Yni3Flabd8n0N1xMT6Fx6v4nNDSb0Y8g/dkwPpAx/q
262OZFcLj7LWl6PgOZTkyN0ADlg1szLtx2bAdJ3lnus+XskhpY+JVSkWWwZQvMrn
3NJI8ZMf2/IFfx9kyrfZwzQ/Bq7b3YaipSAe22nk6v2cNaYcBrWYJJbonxtr4Dat
cQOJsRq2GrXeFF1NheC87hbCZnIGfa0/OYdvyTzxYL1R+pm4/R0ddmdQK+vCjejw
vfIZaya2+n8xZGrmcOa0lesQaslgQwCi9YdbA8yjLe8PtHZ7PQicPeXo+TbABba5
5l7bBduRyJnGmY5A4EayvIkNfDUAzWg/AMxj6GYRRJcFXHXZhTpmhKp7Z70/WHt2
2dXoUJ1Xp9Gt43wJ/lToW1GQFK7FTU7RqXRH8KNtT1OUWHML6YwwUq4F0z3gfLD3
pylK3OI2PMhLCrYR452rwklij2l3bbeA51aeTDKD8Taa321tJjlGHTJRj4iUlyNm
KembMOgP9FOCqvTY4F6Ncma4knhsFPtEqgYEBTnEfQ2BHXeSdXudo7h8NCDoNgVR
8yrBFQ7u0S3ldK1nh6s4FX7UdP7GK1VCiyhPY9iWIFv7bXtqbA0CP+azKYtH5DFc
JFHvnCmMJGzl7sxTKbo4PbLy7nxwH7KQ6EcZ+0vPjc9ridpR1kobgvvkgBC3FyGM
v9Y4KXSLfMFrakuXhpSTfcDG7o1b1lU1S7sPghmFLkw8sWzCC3jwM4tCRroUji/t
BXgTm2J8xyyoXUOIM81zCmQkA00WntrHFH8fbbUwYOE1cH+Jdz69PIcU1HWW4LPs
zVh4hlHZOFsvP76i4fUKhOEW3vG3XQcfNkeWOdrTD9cbNQYl35fuzc66IuyxYQT4
KCC/ZCsO5BB3dAYBhx4ZjQ5T3sCqgjJ9K+a8Dmg0rdKIQRzZp4O4Ppy3k9RSy9Af
DA/3U3Ze1UjvzuFhdcEkbO9FWPBd7txvaceVzjIDRJPkV7WTVxudek+DTQ6SR/ba
6HKPq1rG8hT3BdMKExt2hDd9OMRl+Idqssh7JPv+1DZIfrJOAKIvHsGOBnaebfdj
2YTt6tgdwlBgvdip3ljVTclXNfA2RSPbYECMDDeDxuhhnA4EPc4QE8j4s71d0r6I
dnm557LhqFKfJCxUNzOKmIePiGkO3XyU3vCDGs7Wqouj9OaSYO5+G8TNMjJiHLmD
lD4Y9HDvYdks02gEHHGkTUFDTVdtO1/Rs5qvaLM/6RvIZJaMSy81mPpywfgtERRK
GY+eR8Cp6DF3kHsK7CJmbfBuRRiH8wVlhs2K2GDJFBfeG5HzfkbvoW/dmtM4KhWL
w2/v+AxzWvT0TooDYLk+UA3QJ/DY7cDHfxFQqaG9B7kTLmcgl/qSgr/IWSa8YD1o
KNjJiVFu7jj5pA14TlRm20Dkq/93hBnCri3CVqS1yTQHTbOhu4phUotq4pk6SBAz
wQK1yxOkbkNVtiTieJFjhnL0ZmN0I21zrnCWSBD/aE6roke9ZEaPSy+shtikoPHT
J3UTh5NgIU72h/TRmoXeWuqfhI1Am+7R1zneJ7LiCbCBpwJTJD926dyFfzn9sZL/
8S1DeOr20C6rtJwweey8hO9M4rfpgiT0rl6iKS6nV2jBOQzao5KweulFxNY61G97
DeaDKrb6vZ8gkUkLoJK/KXTKLSuRSsDKlE7q23opB/geEtOLEyPHmlkze83no45G
Tttw0uYiswu29FAvcIYa2TEODubck95jfq0r9KRY6AwIo7RkjX9UTBQvdK2O2IV/
8Cgsd3fgEtq51B8ePUNHZBUyDC70XVR0/Q0mTJTC5XXa0033DZqdVDuESXiR6LYJ
MPbAGUbltG4aQg6LFcMMuJjx62GMLKnyAbP7qtc8hw1C4uIeNk79JExrK2U35lak
mjASQVHv5khjL6UPe6FFnyRjJ1C/2YFpS3LPzLkqsugwqDt2nTobj8yBxtSp0emK
RXUXE2S10EX6l+1a3u7+RWqTg31QQhtQ3++o2dOR4NspwIp/TnTccMWgf1EramYs
hx+2bmBUg4/LA7W+ZnNQQTeF7JnQksGZ1Wr8R8LCfUD2d/MAOCWTnr/UG2Wg2LlE
LMbCLOTHRp3O4v3ATYzCEF0VB+q8BUWZvTXvKyn/uQE0S3L4HhornfFSUsRZv4t5
NAlzUY1nZuv/LzG+fG2NJJJaTSlzB1kkbYbdEvmgLrv7mc9WDv/vmKd6uP8Md2Pk
WQDxPNf5THXM6FOBM4IKwEk+vevU7MdXM4Zktaladt6XFwNNp+f7ykIEltU1GU1G
lKVQcSX9KIubGRdCH2mgyKIhL3+Apys7fdceaNpa64/PsZU0RaB9kWSblpMbFPHM
9F2/hEGl2bNYlpJbHtN6W/WsWFbfcpO7DYjKIWEAMWqOH5bLtEYMkQAiMNsqhXGd
vgMgZ57ESg/YZkqPy2SW3Rc2S9OBpk9bzHBFLT5LfcMG57byGx1UMyAUbJRp5673
x+k8gp6SoIuHZLz6hxolzUxKQXYFZismZMVhVRBug+8Znr4H6EMLFob3px+BhWBM
MAB/XRLbR+5LQbPI5afv4/M40klO9nRxTUoprmQHQxVsEaDCYhlYYu0pxMPrMlPe
q9mfLS9Vovo0c7KkHzej1jZBhFwjzHUCmaNBy/JYxm0S1WL3UHjfJtrJ5Rxz0Uq6
+P/xxGnOK2ssvZpWNxDOshEVJGxZ+zEO7PL/5nFtB8lfaHBxLKEFFwLUTEFtFpvK
P1uJ7FKXJWTDj+m3MMgFus+sYuHGLuD8R1EP8adHThI6TuGFu8qzWmTEz+aHx99n
Xs5i7PAkGWYJ3OayzW+QE4zkr4Nm1KQsn2MGuAwbLP0PLD76fGojIZRYF6XVj46D
yEZEbR80N9SRjSPA7I4cgvkoyycJFvnTb8gFfljEEahV2IuxFVaW/hUCNcHkP+se
tymuumIBYm2yrigvTwV5CmIKBzHo9pWdBoqo91MbQNW2WehYSRYR5Y2S5q+4QrzF
Lf+YPbAzzC49B0v1BBuNYD5QFSMuTghCI1+rPvNgNPH6R4kM8WDFCPojqKMkIq11
IAM0U/jAmQH+T1sBRAdC3241ATVg5qENhTR0yc9ufXTOOV3Kd/1Q1a+/u4gLj+Wz
Ga/DsMT5cOckzkZCYw3l3QDaKtx3f9twQj90XW6LLLO1ka2zeJbBfQcjwZjN+3+G
w/r7RuRswvbF1i9U6CYkCH+rCSOPMJhGq+wx36MYM7silf36umLN72BIveHT8UW8
2rRgbT5n/nGnyJ8P1YoPRQGA8U+ThT7HbCIqhHZ9oShiRr9D0EhcIn6EXV81Qe3F
jpRXvUOV/Rmeim1iyP1ytBGfrFWOnySPebki5qMk0vM+nHnCc2du+OoklmWkMpbL
nXNQZUDnchY5Xmuw9t/w7zZ9ct86H6wnTf3oqcBcb9Kl5J3pzzzFPVqMOTsQduQd
AuDQiJVS9tlFtoIBv5EcrhxF89hXqCkcoFYCBHCVTHEQhIKgtXTH14D4FOEtjhfR
0rUjaTucLsHqvHk0L+oOCXe0L8vjSuYIkDlJIZznYtKqRDTIpTfse+71dje6v+sn
l1mMY1N87Hc0mESWsZTHK43VEkYJMJ65ZfGNHRIVs+0XmhAopNoWYJEQP6ZxTOU4
DXLIpaKhBdnadFXyQni7TFSbVOgJyQUYV/J69BBZedbu66PWYJaHJ7d9rx5pY/Uj
hVQlyJw2zxcYAZDqF1RZ1UiLDpxqIqDqz8WnDi60SYwcr97D1vWWPBPXTmBcAzUV
xclzgDYSnyfkOb6Q8+pb7RNuoqOhCRQ9ccg73Tb8NVE+jDYejwohJywo+Oktyzlc
BXmOpFCVKTqSPruhwyzkIZIQttpsYGnnf+7F8wUk6IF8lIF754cPQbnN3x9v9nIJ
ip0A52pwCDR7Ibhf1r0wZcpwfTTK4XLEm26L64jUk/gK2wfvkm0eLwJ1XMAcsszY
ybGUKXemOplujVoUmlsnZ3hXDItU5Rk5syTHLbE6daSp9jVM3RE4qQM06gTGGAXB
YBtVbxaG8p4w1YJHVaof1ZHaio/nnlwX6OAwwMZxn1ERIvHbIbaAagUHKkSCccqd
WzYIWXnqnNdUjfuj0/qwApL3+IMPnWF64zir5TRVSIGGm5EsUomJWNLLuIzVdBeA
8ZB8MktiBcwqU6JYNKwt6VDOPyApo0JKEdWKXrI/zkWK2VNd0JjUgfo6DonWKF/k
CGh+rhIc6CdikcSQWqf50pDoj4U0z/ilkkBuha0PoAcz6GMc20QZGaDgEY2/MQNL
NBXyK1h/c1eUJQvAb2cNkUynfB8ZtQLzI9IqrKyYIhBKnaGeubpooNQ4D0Iz0cWD
kwosHje+YFufJ2I1dCF+DV+7oApxpPJAdy3D7UAMz02Nkz4cIYXituvtzMkualvg
2AJei5GGm5AbvXiK1PeMRZ2xFKxRV0RW3Byv//GZoTDsiJehsx5SDFh9b5208GqE
Cvm4MPA//KtQHlXh8rRBeD0i5jXnr4rFvmBQ7YlQyWtgoFCgHGfxqIx4L6GqB1TB
cqwFQzs2KPm5UdrrwohRfuI/cLInden071tApRmb6qC+EleSNs6p0LIS1BUbR5JM
6HHUjiHYEVja6znbg7KbNd2YyQ+ulcwFyQlAN0hrfo2zBnKsK0NGAyLM4U4QPUdH
r2sjWrYX+94LyF/o83rk97Wpf8nSrFym8SgNGS76eS0IG7u5J4gbmhIosefN38Og
y5qZoeV67ju5LydrDd/YsEXZY0P1jRbp9lFnmsC+uwLjvBGNGX1Qvao00EqINo2P
ETn8552pq8guH0gucxDMEqQDAmIIzdiKD5TqgXPI4gq335btWcAxmpviz7DKCnDO
TnPo8p1YJ/D0NYWgmfb57uYTWoXkOgyVDgTxYtTxC2QADszX7+G8nihcB6nS/0wk
fa4OaM4u3Po2sB8zXnK2Bm6Jlo5zXpNN6FWNrKUJWA9zuYxVfkebmVA3ZtTl9pXh
kRb3KXuZ/PoSwyQqPjJPU+eihFmdSX8r2iYbeoZFF6Jd1EPz3xf9QgAuNutXu5qU
1YiKXGn0uL7FnCpYXjI7j1Y/ID7k95JxvJP8ay36ArnrOF0LVdO0QsvWHQi08uGU
SmwJgE95ITqUh7PM344wHrh2dWf8nmYwLgtirUJIRXQ60r9tojlNP7Rjc29mYdWH
cF1WUnSwk7TLZC6ucBE+Zy17WnyCQlISlwKpdpXtUQUrbhtHe86gczliIGrm8Qrd
IwC3HpTTmM+tvvSz4IjIQ0l4jxeCoS2JRNeL5ODJTSjKfL27u1MdHlk1j6r3OxPx
hWk7EqB3evFKs1n5Yf2fMmcwYF00TIMe00LKNQwpmauSENFkVEsnh7+lAO94jbq/
2W23JdDw6zuAgoecLcG8CEwwzBcxt3s5+GiA3TeXKsfzNo+4Q1sWMNPG1cXP+/KX
CCaRlnQI2HVZGgLNy/UCPTj0BHJRfVY8OeVNT5KJ9uIy0GpDRVYs2KpshIjFqE5Q
CaNWVNHkLOd45eYCn4SsrnqJTwFSatPLHVklU83yqXVZvnax2H3eOnLkO31RhEvW
f7MqcvrJZV7IpPg5y43fO1DzULgVvZ6WE0/aKzJyTPrgKcXAfrIR72/7cMDCtoqY
/REjFK5QTHJRUgeb7De1/oqceb5HsICj74SMAO0+poofH+8fd5LnNkJWP9Vj+nSk
VItaw5pfgSVcRXvERy76Z1Hit55vY2x+CuCBr0bbAkt6J06cBkjtqFNIS8WeeFD/
+9EHSLC79dgtTZoUviTbqyK5M536Sa0UdC6cR+L1mTR2QLs2IGm4BXg1HamL4H7+
qOdJhcFKakvS/EdVICmpf/ZBXdJpGd9IWyUdWRfIOZysR+oCbpMow+HcUGm/on7h
m6BwJajyyQQJ/KFWz+YDrsyMRd7Omo71mPQDramuAJW/7cUeVbnfv07cIZ/5fB6P
UM/3eH/S2ixaN8PwRiSlYdQUrcgj2HNmSGM9YvwJ53VM0S/Sl2BIM6droCQuWWDL
9k3HU+ro2LIXg5wukCU97umZxQnxffwzFuiN7IbTQAMD2+Z88SFWUlYakiumrdFt
SRgbO5EDAE8/WcY/aha/hROW09Y05M+B52U67r2GB1JPp+oWKHXmXbSW5Vwr5k9F
mHduEj8e/yniR5vXCSCFt0kUQBs8jHk3ueXO6+ZB8B+q+XO1Hj0lyK1cce118Rpb
0v8cCCpzPsauYF4uS62neCqtam/lGCFl57V7MrOn4cA9I+x5B/5dVOkMj528e1F2
BHAlzgIR42YxAzZdhHQAAyhERxgNqEgM0u6Vs2qHYH4rc48Igtxj3RPhYzoPCrlY
57lyxcxvq97E0SeDF9VtjwaZFcSuNeb1AhD9E6YLMTLQHy6QaVXfLfyAMQzTM9S7
Kx9nl5Mwy8UpUISxLOjl7chZ0bMczIjrvm9wUmyZpj8HsTAY1/YJZ1Zr0/kw2EMk
PMhPdp95+78NTe21m73lp00BG4a2XwwKifB3oCqYe8JdNhxTxw/QQHfscckj6MHc
/o2q5/9/8yCjqhpSAC6EfH4bbVGKz+EbuCXMPzIrPPRlYzDo60vw5NPk8zBD3zlo
lF4w7jvA1vdvDfd0hPSfyFPPdm6yhuycsM+AsvwAGVSlJnWCzNMppEtnUkVslio3
6H/sx0QkLsp51orNJqmjyOg3KSIOKQxBENvlG1SReBUIBBrZirP+sfyWGsB7m2LK
apBxMYAiRSNCNKtsKRineulQjYXro2wKfgEk+NHZlKkrjpoeQTzmQSv9chMM/rji
KL51Jsj9Wx0c/lLlZy/e4E/yD34Lt8j0CTkXQVWydiCvsVm1ru2TZTyQPv/yjp0p
pKXqbB2RanrEWV8mO90UiryTHBJk2Tq5hbROG2cuimqN7exGjSwxqnC+ZeIrB9b/
wr07XVKn87XSVhIyGCFZ7KGQs3Pz18Uu6q5IRQyjpmDNdjcVHvG3TYQLqjtAjhIJ
hxgEuVDYums5cjnv2IfQlawSukLrWB43bop/Ix9Up0A1PTa91y8GUmRj/kBMKDRo
BAXfrtk+x9ajE2LCIYF4v5g4hBHRJO6MIXTpNQeyZudQ8zPKvCbK4korNf4HF8ZN
1I0/Uz+UySWUs5vwdSABjGAvMoP+w74mWipj0jOkMQqBZ9Rn5keg/nRSfjaKeuow
7CLYvUSmh22d5isKdZOvaYO4UUxKs0xGgn5uXHRvLr0fpo+PaiWVeLOwVWuoIFF/
zpmrLRH+tZs+tD0O1+M/zZpRTcmVSPQtS7jnL2nccizJDskTkJLrB5dA0BXY2I2w
BnaRJ/8HdzrtFn9nJcDowiAj23LmW0d/3ZA4pqka+4rgl+baaPoiMl68lh5EF0Dw
2STWzKL/0ZFmNFx3b5pSebJIFLBtvVGGadcdoc45q6aC8+FTK85a7HaPJzAxw3T2
NyAGjqgKRGKuFirkWmYkBF2ZqWSeT8eDDeCo9k8C0SGtuJIUEJeo9W8h1yOc0a+E
ZVE0KLiDl1vWcHdF2XaL66ZaEZGOwrN0WnQRH65PBod8oHTp3Gd9wkWKS58sABtu
SPyv+VJddf6Tp9o/g+iEKo+A4D4q6EYcGRBmORTOqZfdZJBzQFCKMDvj6rWtud4T
ypq0dgPBfcwEznf7vRHhTGbAGmM7jAU79QH8uwT2/CMEqv1KI6zEgkrspsqpnSB2
RhS0A2PvvrY7p5bBYlYpN6GiQSWIeq0SkO7lWfxLtPwi2NbchwONLOpsIe6abPLG
F40mL56eF8BjU/aMZHmWLA/HD0TIUPAeCHxNanLXWDxlcQMUBXETskmL+OQ7p67F
cuSLtsDk0WuvHDK+0vFRT34pWuG+tffDEdGfuU/tUpyS/qsvC7TlIWj1d3Xk8fiK
cseeM0g1umXIHKq0xQZjQFpZOlPNNW0OqouKJ8eAJSiAfOSCydFdTuHt14p29waQ
y6be5zEYuPEWXVLy22Jy7VCVXTNXfCjq+Rly9+tfGIkNi0BcZzv8s3I8veliMYK1
vulCXf7cbbgpFKldWDl8XBy5K5zeiolykgcWfv6iQ2uyxg4MQvUvZ+Toyn/DmQJ7
VrkImYqJqpNSFLkHcRODYgySAhaV/byKVsixygKeHll+3bDGJViq/OOg3kMirwdG
/lMRWB71OkYn3Th4AhRaLGj0Qg5XacIn5wYw3Tlix7/So3qf/DZN+HtZ0Wxnmp8R
rC1xSVpIwdH20oSsQZEdADeE9u/AgtmdsUbIW/pG/435EJq3PV8IxHDHAGvYCug6
zzHgTyQiBD5rMIzNI8wGWTG/ldwuI/bSlgGTZ0EnqSrWUsXNJU9K6JGYX4RpHsyJ
jk++ndvxhFO66a6svnKqRFP3MKJlUT+p8K3kcXoUT3eWwQtxHwX4W7Kdcqs3+vbv
X4wVDDJ82FwOqAFqXanQ5YjTKiQsALWqz4j+WV/LRIDd14o+61Wk67aorjLvTgYp
wcEYw7hlW6QGnjpEoT5HmmT6HOfXL/pkU93Rna0lLkfg2aGnguJMhCNbNJkGFznc
+VCeSJ5JXASbSPvF8h9rY9YRLPn8vRBsdjELnUfmGEy1LT3cfhxbAlaq0o0DWPq3
T4q5VEr5MlQUpjItqg008gOTmcCshhheLgv5MvAy1lpCAKC7TTiseW0LFW+QoeoU
QncIRazMjuqujIe2ZnCVMLpqk3LfRvEB2yWIQU3+vegX/fGSSkOC5+PawJYhhG6V
1tjUlGJTKJyIgNG9/8LXRtrwhNFyJKEn+pRQ+mC87Vjsxlyixr6Lt9ymZ6HpAz6l
uVKZGoAamb2Ci+zG6Ho9ULmD1QZmhzZ3NDLC/vWXFH9I2kuzSWXNwwAU8wo/fTf3
NsgHv0E4FyHb9UCJW0bIkQa/+9uKqy6I92AMNQC/+D5URZi4rYb6TDrmP4ubqahT
1u+uF0woQnPbv5pVDOUi4Gaq2drc6Cq86BZ3/dkaGeykn/kmvg0PihDXQeYExm9B
aZY+BMTfEtUUb9kEyn9leqAga0kPYAIKXP5/P2xKCk7ez2EZf6eaTGcEMbisXHdt
gXnjU2CcwS8tG637gjQKRCE33iPeHCEbp/8WpNqOGXB1PeDMmsoui2DIGMcYQoRk
za2/eX1V2P/po4/pEIzOWX0wx7QDG0rAWY0zh77aBacULzgU4i1QBykPuTMjkO+o
nbMNrnUU23JtEjkfIQbvznM1z63BIoZzDV8e4E/QQbMrOx0ciUARefuLgiCm5oGN
3d00DWn+3oh8amZ+sSaRLw0itTkmN7UikH8hQ7pmkn1UAJqZwbNjylkefgsNqbUi
fOsjI6R3lMHdrFx8xy8pl+hRz78FDRjW5AlxRBcxZbgx6QHfSN/DgMYy/0LmjkPo
Q56XoITSWL9WyiUYJNKEYcnwHDzxKH4no8tAM/CKNqRsJIVl0CIqb0IwDuqrJdrp
OslwWsmdJHMCZozT/5DCgyM+cz+sGK7eI0nBnZMOfX7gbv3enoKlYKUL0HCgYSYR
qeGfz8o2TaLkm35R0aeqy4cjA8u4EFQ4pfoVXmiHYWCwsd8J0p4gDtBESN76h99X
KPDc0KA6T44lZm/AYn1gmtRs42EhvAtvA60lRq1c20Ag8BLc15Fcfc2XQrDIoBnu
42V6uRc/FpdccYx087URciteloWdPoaB5TxwAFb+59X/tTzNMHPRNkVm6W4aTCiE
YRZbJEyarhZeg3z8X+wVo+3zacfF6YqC4ll1u1tmQ2vZk2TY9OSTbCLXYVACJgKm
Ez+HTcX5YMaDShF++eguDlMWwTJRZYo4RuMi5LC9LLrvBaddeGNsy93EMlk5V7Sb
FaIgrbqzlcLY63ZOYYfeHyr07uzR+VQVpGNMsCsdvN8g4G0NEXhvuYGn326tfB4L
GBAktc8fvF68touxU1cl1y1sPwAiKqDEq0wK7lf8bGZd2a5ywgFf8tjImlMWD1fk
f/ZHNCoxu/SFz1id26UiZYAYxhIJQq5k5O0RrqCDAgTcVVJM9x5jOkAXA7A0Lr2B
YSzgKY9J9FNFrqBKhgm1L1A7c3PZH+ZVme/Ngdw5xST9GTIJjCjnoeAmUyBOxB2e
Ae9/pnUBClpYs/REYJqT5IX2yDCZRlcl6opb6dUXGnOvasxGS+NQJNiqMy9rhY70
gX/JiCyoMAyKMTeab1Nvb80wZf9bgEhPaMM1dzL63rMwcFbd5B/Z0X2gF1XqR2Rb
afUokgjLtGWKTzsc2zus8jfXpw4Xww2KTYtN3u7Wu46/dcteD+fytQ69W8elt/9o
Lc3deglCMuKVJcpyIZQNNxZf4QtZsJJUWwmYyJpf4RKqQDx6J7IFlpxgLlr3chv7
8dzKucO31XIzTreRUcQgfrzfHUaJ0mcr4WBJhcuI8Ux0gsb1CdpXDzqwdYeMzPIr
Y2fa1cbY7DNKquZVozp1vfmS76zu23IRUulNLdAiXGzrDtZOG0E2WDtXmdqisx70
1jLWN+e+wgw2NkK5oSova85WXJhUUSLT2XrFD83euR/wStZ+cTumjWYXjd6oPVW1
y5YJxvSoJbiD5kM6VxDLJI3SnkNF9kQ3qRDbsgpVyr82BQgbm/G/uzxW6CkVqoTh
M+ZNaYde5cx/Drbp92sVU54m1twuY08o8W1IUgXTQsvKqexPZeQvo5qNXjV+Q3yF
JFzHNkXyW85aG+7MUwfsUzQbb+apfL98YjmbTcIcPl8V+g6AwwV+bwylUrkva90k
2Eey9x5nR5IDOOk/mtaV3wJzw+hZ/vp6PmW1mvgiwtEYlpfiiS6IM9lVWOBEji2e
jBfdpg36ZuQzz6a3WoMH3x5pEQz85Gkzhi9849BQwKLZjx9JNjWzUF4gBPUhMoaD
Fn9cG1gC/8nZBg4234UfAFq06mWJhKkCRvh7iJKgo0JGzoNIerhVs0JRoNrGipTi
+XRMtEQj3pdXQLwklczCeAuIFIS0ZJOc5L0a5VkvnJhvOtToIvXLwDNUkDRa0l+T
FvY4EfUVGvKLc/mt3neG57jjWCu+hbRTzsZKefgQQ6BV7xTfTsnDAOwaAtlwip7a
b6JW4UFIuJoEzWWbVvTaywEL+GtZBoQtHP+zcMn8dy/nrrdsuM7gs62xAaMqlm4j
l2SngAvnQ0kAQsi7pSxfNcw/b53ojDuc7mKmNXJt7gRXGrwj6qgV8C8RUT5xW7Jx
ZKSb37yCZWsh2x+3W5KfrqFk3WSyePJkxgZ/Y4mkNBYhC8H9EhVtPQyH7udNkSnG
rUkpxgWSVw/reS2bfXWKfhIzQW8RQ2gG42NRsNJ8NtZEx6nK4jQ5dJBxYmgtxr3z
R48VstdXVGFbvFR8/Cr887MPNcIxvlxhQY9zTdc3DSyMTcu62h2eGAPOAyPoVh2i
BwHVTBy/bw6rkZzohsnaxK/5EwvVJntczVFlKjMpvm2L6DorLhgSU8O3bvXbBGoh
EeNBOJ1nM/WRSSXKR1+8p+qIVryH1Wrr5N80wMOtHXzWF+Lr991eiy88O4r2qHwr
IFKjS5brTjs3UV/50vO4zgoG6XAY0iy7xxy+Bzyj4EOeayl4C6Gs24co8e2VBtuf
yS2hSO2/fAbRc2CpqZK86sgFzhfM3YvP/EAJ8RRdvPg+MlJDAKWW1eK2rUCQLWXv
y9SWJ5haxGBQheyDWzyCtYBTbDK7Rp+VpkuwNqEJLAJC5CFhCtfYP4mQl5zyi2+l
uLeGpDMaRdLM7pZG0qXy1rhWR5IVa1ewKvpWvulm/Hg5B/NJTBx/QdBSMfs8lG1F
m/uwq2RRTjAqOKyP9JHsQ3YhMwPYj/WgzXwiw3BI5hAKVcKfKPk9Zih5Kwkq9l+C
/xH7PTO6MdcgHfj/JN1SoFQ2//tamOm4JhnFUJb7ZZ/H9VE31i3zrjZKa5tXLN22
fyz3+5vCklACvPNEyxp5motR6kGNMc2cxDUpeJMxm26BUwzgHDXbN+fNfWapoKIS
s/Iw3av8NRmmOAtUJbh1hdyk3t3pMMV+dVJCTmj2gMuB06a2eyYtH2X/O8iYu1Qa
QeA/Kdps1MI559MNHFibkhIDgJdJeQg7aNXCuYs5C4/P9pDTNXjc6BjPS5jJ6w77
KsxD0qNOObY98BIvc9GxaLlXkVWC75bdndKpowhkULcCOzg/zRY2QXrMFBfJPtEy
gFNFFaFTBy7H0YuHzByM/QlpjP53vqtjakkM0U35JCZMNJ6/HyfOyWdEG7VRDILs
KcbRMXT2yva3iSUW94e4XAUNyQZmEd8JpyV546SRe9MmjSMG/Ha9xvXF26REY9kw
VDGE1qL6kzXxS8qC1TxrQ5NUrXKIAYQZHc3bqbId8ylvHbN/5JnWpk9EGDVVYnxl
38gJm+iZQ5gfxkGEv1eC3N0OXcZT4xRisp9qfcuZZ7FnZNSA1Goqr40c5GPA0dfV
2RQMIWsZTDxIYg9dRfhCk2hPz21pfGwGDFusxrAhXOT7J4xdA0YOp4MQPCe0v4rX
xGvrxf7r6ackSeu6cF79uYkLrl7+UgqUOWCHjKqTV5TAVDWQjadO0RIe1FXwf0Ks
719wXy8trXKb+E+rjgbml3DV8cWkc/WddoT3aWb9zVQj3wM5nuosB7rVPfd2bLaD
aTqjcMrB3MM6s9cSFaWMcfebNIxhX7TAsTyARXM58Tevtcho54UlMhcU47sYj6+z
k/hyCsYRnBNS+IK/hiasxdl6QbmW7DEcauWRh6LhN7IaS2zWAe0kh/0QBAP6QytH
I3t3a7IZ+aybJ9w8ECJxp4ATaaiOhhvTTQ1XiKMNSUDryTPwCMYrSQ0ZoLeNEyHk
5IeFg/DRGaTgrKk/1loud6M72lvtAlfjL2EezWM5P4yBtiqkbslWrRdFxpMW9ohA
lQwTj0COQnU4UZfXwKihpZrMTt8PhLB+aVLi7ME4ceD06x48fjYNCbA/QgC0zjkU
o4YyEfz1UUocxxr8GFNatChNPgHPncRmUqDqAbhDQmclg+iB/LpPgEmDOBIQJqon
c7BfSb1q3ITiKhpO32MLrgt2GFposuJLMLioNBVQ+RqbkoyhWHtjexCC3hzji35Y
dNNg3bJqmKCj7Uk4xtyzdwpxFQCMxLdRSkchMgcrFSwXIeajl0q+guu9lFS9xRp1
iXQrNH0j72GfxNcvMIF8zvXFqRQ6Bg/svxoUdPjt8fb2vIoXrZVhz6ic8e89oCV3
RPAo0RkP4Jm+ibWsgJRbZm5YXMtGvttGGylCPGO2Up/rW37XXC93v8EzfIfswGpa
GO/3265VcUdFIUt1mu9dNxVBVxxKwVx6TUleVUbhz4K7aAKtLjo8c+PxY7bCSs4L
Ecsacp4/IynbawMorRZPjNmgh7zcs7MKGHeBSoHYjir9ijGTV++YPfS53u1/b1k7
gSk1VV9c1rVN0mzuZFjVQUwKzsrwygQ76aucRfTCfO7vqO+Dy72dxNY6L0jrt5t+
d/i2CDiAzcwTCzAcFXxpy7T5eh9SjUJy0wOgyvYl0Vg7rUdsDX3dhWVCQB3Op6Yk
4WYxfAsrIBgT+ztTkNJq+0MZmh9Pcw8k7Eh7SRf0C0gdUPwvmM5ehu6ME1g0gcAY
h3YLWqFXbJvnyhVsUN+kSuyHsToERojcE/esZ5CSfCVwbh9QgnQbEPgOiw5tZxxN
qSiISP+6lo1A7R3Rf92lIM4jtDkhgeIzM6uFzT0Pnia4PFLyLueIPhGk+WcSCXom
KkLINjeDG3rbZlfvAZmb5qO0fKXyf324HzheOLiRZWC6S0l9givIDKteMLPeYgPT
RDo8zR3tr/AX0FU5hKdaVSFPuEyY8VSb4lSh00jcr5zzIuOJkTVq38Zk0U62Pqom
CfiaqudcjAkX8aJ8FaQUMCVghLjILSxGW4cC2XlGFJnLUdcsTaXKHZjiCFbS51nB
xVvwYuDcGP7yF4BKspawCCoZvKg4LUIBirQrNZrFKII0kQ8uGuZ8okFCQBHru11l
KcNNEgouD6Za7n0Mn4KPpN2e6YRFvoLM0AZTFUyln8gywImFKAo1m0A12P9lc8Qa
y6YtcL2zCodtPCYOaEs0oPhphyQFs207coyj0KVONeMZYoYqgnQ8fHvuJ23oaEQA
oC74JVnA0EfDr27Z2P6E+wgISoc99xastyvKDTOYdaRF3PSjdjFcJNmgrArQwOG0
UJwqOxthEyRUGPkqTQrwMf5iAyehR+6TvN23i0HLA0mlDssOQrkpRvc8hx0tHdzs
5vMc+M/lY8rRnyqJVLP5G944HUMjzZt5WSxnv+TgT+Vmv5gNfM+2EtQj2ZGFTF6E
TL9agSqXOyKEfOjg/5KUP5oNG5JXXRX0zvi2O4eZOoQzD18t/a8F5h0NceffIZ+/
nq8maAAWAoXef+fdHHOQvL0Vw3lJ9iVUkEplNE3EIuDqr6wrSmqKJcqpRAvYv9AV
kha9e43k5YBWrf/quklI+rZoNqnMbKos7qHcNpn9up73wzSGBQwCNijEOLD6hYej
knqOnuielhDm8IOoxXmyeuYD7NB38a7FJHAe8De7qUMcQjivna2pXXRm74oAnqB/
mg8Y9q0sfeGsFUh92Y3kYNz5dnegCXKrpsQbQBbUafBli2+8J2gbiOfLxSYQ1igD
dbiNJh1ob3q2/ltykodFJ2CNxe3fUytAoCp60PmegnujJ3gecES1GG6ACNn1xxU2
w12Px8ev8W/PWsa0CG7t+UlTx1Dw+JGUsyxTEsll374S5Lz6XgLj+G0CfDCOUKzH
/tphoyz0H5o3CexwMpTzSOne0VKuxjJ5pPHZL00w6QaUB/dy7++H+IKkshWYWcHk
5HIg27tqTBkNK1Q1VBI4s/vGqfHWTBncUnepEfEoZlxqnRsuVTdR0eORXaFg2Yka
scyHxHFPkB/gzcTbb3hoCoE8ZXIgP1SFOmnlW6F6dANYQ5FO/ZHoWmDtrOtQincQ
skc6iCMWtiwBsWunChnwaAkZzn/dfB/Li0j4NNhb/IX5XTpRCLqMuU/FC466K/6K
sliLVRvnqo6VS4XZJQGsomx3CBYQkRMaEyonBpceToGmdWMQa8RlTUlXqkNFZGHZ
3EQt21iyGkm+zNL/7k52wlZOHHTZrNC2rCFM/J9y83euWjwECXT4TRLPnerVwT64
F6ZP16xXxPaYuSQNeYx9mx9gdDTjAblaLo5bM7lFfndQ7eYHBT/QAngfbmyaogRD
XETum9mJoG+0t56T2QQxW/FVOZZLF2IrBe+qs7b19bBJILp6uctmVVnqkLwan1tx
7d0lG5ix2ZsXxo45mm1S6W/R3OZ+Z6EA/9C6OqYXgatBTdl7JHktt46AnAtEixUu
CerW9eW6609SSHwVoxNKzMmB7Ic2ufXALnVHo4LX0iXGOUXyeBXni9QR4VMh3HSw
y0FpVMiA+6ev0Pdqk3yby+03y7wvI6oopqbfPwtdeWKmaI7jhxOscfgMEJtq68tF
Swss/YFWxWoe5TQeIt6FMs19il/bs7fuvNFIoGY2zIeqg5q/oAyGUHUX2e5HjM0m
PuqvfmMheQzTSuLczOpCnyajw/ziVnLRknSk/mNgQn0R43NzJfy4tV4xd8Ommexj
KYH/TaXZ10uaIiV3A/hvi3j/ibMMeXKz6ugXwRqdzzdM7+2n/ZkmG4FoW+EzUtPg
zL9Z5bGKEcamXCJbodrAprv9397A3lqjZLXAlohyftnE+Md6NhWsplgDNOAeOzD+
adQrdMX4UUpqfGEG+lnQXUocnO7D0McGd0nmrnhyRf5oTLjweLfjfFcjtmHq6Ayl
Bv1+UpxJSJD6c1HujcvB5fVUyEhcR/bBbcl7gg9fsx7wQM3899ofpBdQfXieIA5/
xUOumN5Gyk4uExUl41QB9C7U9KhAfQHw09j2VB1ZIRFUfgkwpkUwQ2aP42k3Ic3u
vAGiCJ9sXsy4nCJ/iCfzyPT/o04FomYhjlTu/w5ZCkG8l/3ATb/OxIZeK6gWE2/v
zHrRbQ9OWOqCYCO19fvoMAr3fnVXhVE4mOOXe53CRlI9/uTtZEl96gkntwIk4wgU
tml3Z/eo4NLsrtq6kSwrYbbswB24ACN0OeMeDC85oVq7kenp036rijJ1FPUjTDyA
3wCfbv0f2gP2Puysbc3M8/PcPJnFpm2bTs1ECH9uwN4wcMW5LneIvNUYnrudBlhF
+SEOvj9oiL2wCviowtIltX3OUEfV2Uke7UjY9DcesQ2FLc5UKE/j4QWL9HkMf0v6
P/alm1KjndCUZPXCDyS+apwH1XkqRbRSQllgytLTbook+fpWJ/DG/vb+gwEaZLUa
Llr3vbBHhu7CSTjkFBMjk7jW/375WSWjPuSj/JUadO+Mca1Sh0EOcuv2Kts79OEq
8nyx3FoupsJoLdfmSIEqwY2d4RyqwNOxE6NKgKOzYPNipiIEdK5CN1nHIeScUSjE
fojKhkcEptJT4LPuVHhjyJr9+xpxWCOJ+ILz1+nb0pdKlPGMEM3ESB1Jrr2lIG2e
YggcmSjxHPnBbkkchF+92EKJv7VOc+ldoG5a2DAanLySEBRXIFQqWDIqKcf8Tqma
/NpxE4Nr6d0V3AcrQE4Gzx8WlK5zhmIRj2+lo2wYx9u2ujEy3su+Q2oZVT46HyPH
BNsqOT1yd5eujEI2Gd96BbXBnX567R1ZI0dDGtWWfQwn5JubDX5yFL0rnf/accjI
zpXaNcHuH2qFYGamMb+8WIOJJpqWkuz7Xnfjpn44HtWrBeeFbqKcP/6Hr1nu1i6k
OvqbUm5qJTI3oSg6C86m1X4t58vJ7Iv6EVpzVYhToxvMO+bymAeH2oJJIXWhpsY9
jFpZ2OdXicymWtBDxFw0i+ev4mDeJXygelYHZgMjd4WRR8CLHzQP4GYYpwgMJaVI
TLRkF8FsM4hZX43NMLzpVekcGctXK0h5tJpPzkVL2L2ITzhxdWrITssyjwN59HbW
n+Eh48nHrD9E9Sz7LjKU1Un37WQlbBxxF+xU8BQ54+aFeTtsPgABhfkBEzqGXy7T
Ra0O06wLKHyQ6HpWVjG5/LIO0Q1tIKXJJ/1jeFWc32MOp9ESyZLtYbfkitfEEYQT
dsuNxUeLCxwtocHNjRJYDyMCFHjQwzvf/E3bC0toQDdXuvWV88p5bHsflZRTPIj8
bUFsE+TGF+yVq8/msCfPdeEwqHn8s1iCZVaEuadjRe3aCReYFgu81+E6Fw4Vbzy6
HvRZwEr7PhGe5+F1OSfUoaTAMtjbL+kVD1fVC2NoxDh/ptJrJbC1nzv2UTWlG5sf
VGEFVgCN7TlYvuM2GNcegz8oCsJrUzrWscB7aY8KAcz7Mt+EDHgPQDJhONinUpzh
B2znmZubjNRvmBnB9xrDmY3Q28mu3ZicCWfoeLratfH1D5xQNIOdrg5KfZJV/7L4
B7/u9JlEGvSRXxKaAsxQYRVAPwqYXR33ChBegl1T8IoxBKNnUEHzPcNHbOlz4f2A
9NNp3w3SAl64hwkMYEYBCVUqgHBDAiN/dPhCqZS9/syARDMfVuxIRtfETw+i9I+e
u5aVjIzmv3IZl/UAJhc+cGzHShMjvHXNznXDhyB5i7to0Zx1+OuPYzwdw4ObflDZ
AftzLppq8yLWCrA0SSd+Tot96/YRPSVsswPO+q/zQWY2bFrddCdwn16Tfg+hzCcf
sNMexyJ396Q1ilYNZ+Inv9O4P8HNqLkCtz3sbvqwuiSLJUwDoT9M3MxPvRFXdIhT
2nOIF6I2wrMbplpZHvNR5wVmPpg7VXBlBQ9FblTf61GzAuVF9/rtwppcl7hcDMAU
l94VpyjtFbrYCS2wCRHWNtiURiqizAuscfPEX/eENmYP+pIaODuRoPvk8yKuRSKt
D4wjl90ybHOOUum1cVaU0N9c7/7+bZDcJB45aK59v18YIwnf05nhTkFvgrxBksIN
aL0mGJty2u7X6NIfZ3Qemh/J4Yr7fpcvxE5KsuLcnMogYBjPxaFGumDmv9MZksec
6R0NW2q3T6A9Txi7DjmPvspIAWGyElvp0nzijc2yNpN03UZ696ILzWqSqVhHuOk3
MAWMxxtSz0+z348Oh22Xytc0jklqUgIX8ZOpp9ECEUTtjfQQWkdRmsPxuIDTO3Nc
5eSlUgZszG+NDXU6ViuSR09oxElJ4DCmTfVeFdiSzwIOdo46RXg7nMtr1Z0Nl0nY
1Um+p8+5tZD22arSbuESx/AAG/z5YHvcoPqhzA96TbWH4UGceTImJZUc3ePPQ6RT
uWYsu2OlBVKGHbvyCVPnDCfiBXio2Pe+6HF8ziEdo3Yz+6Cv2rzdlsRkYKlO94l2
jd6oEuzxcA2RyDl6zHCVW4LUSVfxksivI9J2l7w7Wy0mZzZhyDyryQpDZAOsxo0n
V1ckJSZlsZPuFMHnU2r0vyeEIwkR46lHx9yACenhCl7rzfmCrUHJYqyKfOLZ0pL6
L2yXntx1kQFFHd4SLq1cAdmyJboeZ318dnzO5CX5qpq929r3WPwXd6qjPpANslUZ
9KRD9z3y/2ZnZA/RaxsECjiWJmPNKCCF0bRyuJSEEovnet6d35q/P04fnAkjwyAP
KftjWOLrZtHcMyKlePIYES/Dwiu8azvOW+qVm0F/JtDcpoKHOfZtg6B+SpsqKHgN
PruceEzsYG4+FHBwYu0tYonlVCDoVEyHUMtoyqth1NUTSi3IJndiepLs7zePp1jV
HLt5+w8Vt+AjLEXShpdZKL3bJL1QiNiYpQ0Lbf8LkU6sPGs1ZDwBeZ7BP/oYSoqh
xftIjDMEru0ZDePRQcxArGLdM/l5MfZ/1WSBGKEHiVTXxxKS5lht/11hc9gj3XT6
Ej9qbi2YW3HuC9IGZelb8WV8RhOqEwBE8lwz1rB4xKWWw7pc8CR4+kouqOLYK2zj
s1dTogD7YO216rnigq6lEyrvGCyxuPpDY5UcFGvGx8DwEAGJ1FBWxjt8RZUFI7jW
JgCceVfAAoX/z2ChaX4qWvbo1bB4OqPpCypfSJOBPUm6pwafhdcyJZetQCDKd6H9
pma5RpMjQCE5LGcgjGDtKT+D54WIc8TsTBYxVFd0lPuQABsZDVMs6WCoETCgAqy2
712iKaZ65osB/VWiO5tnEnkioOvQfwQSCJ1ei2xjPjCwqH0DQDqgTw3h5fC8+umb
dX14nMlJacJwZ6ZJ7YxP0UBuvnWKQoMwXyiioIYtMli0y/eNfhDoZOHNtsxKHBWJ
jElgURLgekE0QsO+VyFwWKrTSMWgJ5S69XqSYnj2z6AUnqKnPurh2mmtDGtJP5UD
CZe2EEfLzXnpKewAy3OjRwMihbII88oe10UxMi8jeMBC6w5nTGykFyR50NmIDpl9
NG55w0MMIXioB+Epj4mBUYKpe17ACJrSdJ4fp367V1paDBdUdquUhWZAPXQ2jvdp
DvL1xx2br+Yy+1v9OABREVtDBMdI03LwmBYGEe1ND8ky8Z+QyTWpkjtA1D491W08
IsgEHykrIporOBCSl2BeH54hPOdJPZxYn3HXqBGZ78Y8uRMV8Mguzvcf2d3uhNNf
sZ5O/InqmwZaBOJGuV+AWB42P0GjcfCHyTVi7l6vsnqhxqW4Nftmod1pYwyXzSty
K5er0J0xrQp0nO8WdlllhtWTysExyRL+iSshtX9pTtEOFUI6SgaEg7/Nffeks/Lq
iuOW02JHGv5ymXdnGhzidhH46Id6aPwFk3IrbbhmbP4hUG7vXKS0BJeR/0GAv566
VqJ8arDt2QaCOQh6BDjJRo2nCYZWMShykrdNfueeEmnMVU/mis7uwJ6oTIEjPXXn
5pArXknJiGUjsCQkjeSCdoTdZ7FWVcAVS+FNGKsLkzvLIag9xhZ2lzV3HjFtMmEy
HurS5578lRBSwENspWcA0Fyb3Ynt4VULWVW+X7m9fFf0sJ8W7KCBFa7nJVk7KRVR
tCMPbkuBcAiSs5HO/G8jJOP+6dXhgDxHtZbdnBgkO243wTrGD3r32+vUgpTlS/Xt
FIVj4SzcwNRKopFxuSj4TcKl4NsKFvPkU8umK6bX/rZ2zhp1r+XLyUyaHyuLjcUd
pqtYLkP51s3j5KZOplx8yFIdljv1+GV5DGVBVm/6eCgs1TLEqfJo36JqyN10lppB
kwPBZKdhST9hCBfqgTkwvzQg8LtdazHiJpytpT496Tb8O0fxHp/x2LpZT2nskoeF
qftWw4XBxfNHBGfNm6SlZgyi/I4tc2rbXlMwvuUZeeUMrMsmQtFEds6///TER0hv
Bd/l9U400v5c9gLSE3us3bAEzYeNqzg/NELeRpT0BHreQraT4cbRkY7caPf8CRrx
x5cfxLFfkECUvRlkKEud1kShqlG/RkAqVQLJWRB7fYAqhKO2+rJ2P8sCKtqLCupg
WzY/skoQF57lkWyXG+cHvD+N4zfjRtDqneebN9PLCSELIsa26QWSIk2501PrIWkH
squ9Dmmm9iGbzoPRRhAoH10Z8xB3b7D6mIgiAo7a8GI1966u5Erl2ks0h1BRuTtw
3GPmzLlgwtJD4BAuCOi+V54f2czOCgtt//HtdWb5gcuhIAXHECoffk82ZmRRdn+i
fpv6rQ4KQoZyzg/kR6pslyO6QtLtEpBu7vYH6mZ8E2PjZJMQat10b38C2JLZYTxG
2/IHO+TTNCEQHK0tdNtucw74fE8+5L/JNQIn1SNu7+y9369qmMBAeAvt3h8UtTk8
RTd+BMOwJlTBDUzzermS8DCatg2IUB/CqLnRPzaAEhfvNStGi3rttos6L4MjH8Tt
9chVdmL214T/QQFODJ6+UtSbqKihQZ0MkY1KHIhO1GLnGxn9fVX5jQO2JE31G6yV
Fjnica/pXbIYlXQ6s38sIs9OUtTydXegKAaebRHB7e7I+92JW5AmpXXMv8ZexIJD
HOQWVeOAsdwXzFRhHSYKbcFooPykNGnDxSHy+7e6bDgQP8XhC3b2R+vDRXy03Nhm
26tfzHUybxtHBqdqLNN3vTQ6LkbSlyifEGdhF6cNE9aWBA8N5WjhXZodt1SqTAy6
r8QRBgzu5EP/e7QKQeThqHw5DMJ81duEbOisw8JlmCJDJnWrE7WSc+3vaVfgt4Zy
w7YIS5PCNbQY4oTsjAL1uTcUe4zk0sUafqarNnPiYcsET4b2GJ4FibykAyr/PqDS
FNSL6tUQf+WVS3LEUCkQIX7Cbf6hFZiAAzZeFPyOeXviN0ibL+fk2dGzD+cGmqkW
lDfSh9XlxWdK8fJOg/w0daHUBZVTiLewimjhi0PoJ277V3w5goAo8UEg+0RsKmGC
7Wu4Bp18SwO16hc9zngws3mGnV0vt0mGkDP09c5J4x7HIcq1l9kA7IJlsMydx5UQ
XxFaizoHNpEiFe5OE1dOvreb4/yPLIiJGlFACDNrOsVAIYtvRLmNbMklWHMng9al
rLyezWYLqZ+wNmAXfrpM17JwH1tbkyUvU2cQTVhXC4AhfNQSADfbwPWAKjxY4NRj
Y1L5QG8DSJOic/w8XgqY0Rn41rXGKtYPq5Qj8Ez8Cf8jjiM0p911x8c/rFEqQUVE
iSzRP2zRcp0ceHPWP9YpKJ1MHcJAeAz/6TvUlEbqUIdUAh6OiDuaJuNr9x4V0Epb
uTBsxt5P7X9iyN29QazHF0ayoSatpvyj/4aDx7g/dcraRt9E4MPZzGcII0WwXAqz
xzLWbu6DwQumfrXh/rzv3n00qe/u1ReZZFC6KBTZPvDgXJrncvc2IKHjHLfUlE4S
3tvEfLbrDVA8+SX69egdmOHxvIkdCVDrQeXco8dg6cv/8pTbvRJuvWptA9op/cQI
Wks9oqdW7gS62faTebjrjPZi1UDChX2Yf2E/YTlpIrfvIn8cW/ejsJm7/DOM6Zru
2nIrBeDODHCPDEuXHb6xs9Xoi7CXArPCdM7BaZCtqD9ljZZtRAzRYCsAoxgRIVNt
k/C1Ox6T2CU3yMbZFNODnMAZXjsiGxxUlLeXhcrCL3awiivqgiwPxZ1h85QmXImO
0TWCb6i8ufZgnfsLGvXI4wsWETfflgrMpRUc0A3WHX0R1ut8eV+GDV6lIy8Dcn57
yhuls0W6BsKr3emA93E4/MFYtahFqhI+/RDbhtfCb0dhzdCJ+Qlw5Ar6X/2v9dFO
2f/IfDm7wA2LGltVQ8rviCmNr3Ko1y0OarDEnqnOhh4Ld94voEDerSL9nWU7yWMG
5/qpwnQmpBTOMg4WPCp1qKVr84wTpEE60SNA1WA5nV6xxa41Vi8JO4v6z/0B0bnV
mvBYqFQDRKn5/mr1k0qvxa27poFRtLpBhXE1m3JFLVj/f8p53OnaiGd+ac5PU6Ro
JvQD2P+4JRwwh3zuqlUWL9PCu6iMXDd/DdeeA+1y5/8i18++H1dAwTGQmpSBKQKP
LvZiXHbJL9u1252fBIJZjGvmQb14ePp25wNH++v1hEaHmhf3fPx5DuHrWX9ARHUd
PCSJ45k9b+CinPJYmepfuWauNJGIJyXWOaQwlBq9lyeS22nahhke491iFTgAnkod
5wblsqc0TFp5tKYpwC3a3K7N+DUU2tvseygJfS6TnUowJCoh/0VRuFL4B4EtRUVs
6B8I4U7dDJxOk7uxmbprFRa+uN9RjauN7L/H81EZa1T2RL6LD7ozNnL74Hr9hf2x
3z/FqVAENxm5BPaiWoXP9e9LWwCkrZfSBVIWUGEjCA1qPYSxW9hdR6fYF5xIx5E1
oLcDVl0Gm07qLhZ36gk3c8YoFqIwhSEZI8c3UucSbYICPbighEm+5Ru6HYmj77ua
iEI211qXYDpbnDPbbA5+m9S7FFRUAvoE1SnDJP6PdsPpsqAJTs4TTMY8HpRN3sTT
70NCmnTvc4V6LsiyCckbkyZOe2uBg4Ym+09YmV4dCY2XAuOlbpXeR8KoNj1DU+bD
/LTofx0OF+ZXnwKaoXSx913YPHmCKoXQBtavl5JSOIOnbxJ98hp9CMAeADHdKrqK
WtELYE8EFJCDGBMBxZgQY/kVztaKCLQPVp5Xp+5lkwHUQ2fttmUaS79f3iGtwLJJ
DnQyxxZ2BsfDlZDNAnf0AsCdACOQaakIZbgV/djBzScNkrJGIA3LeMDvNzdwcKJd
h/9yCGgLLmbsfpYxe6mUchSANPaZeDpDuvZBK7A3OhItjGVLBLLMGiUZDdjWRBfG
5LC8z0+Y+9E7tZzGpazLmjSEpwHUJvjlMTBciQna8kMAqb3y/JwUAxsUpubRiVSm
7BWToi3QhrEQBvNUI6TGTVDQnJqF94a3xC0N1nyLi+0KEFpO92k9Euy/EsRKhrig
XyQL2AR9M1jtTEIWy2O6wAdI/2EDNEfmAkWIQyGp0QPMNoOKwYJ8gxZDs6foMhKI
oWIyOij0LcfewarxTeMSYQUKvzeOPSlZyzn/aA4mqxB9UYoLtkEpfRMYZsTSS2Yy
nm4aZDx7sucQ6a9xFwQIlHrSPjPYIKFox0soOjmwXbmqPQIaKDDye2cpTuEU5LPF
fEl0DVb5SaRNxtqiO2JkysiGAS4WA30vbKD+zXm8zoq6V53yT37hwhZ+i0A9xqNy
k8leCXqgYEljxgwgeQZPAdhTQm08EjPKImUy5Jad2INIjxZcdpwsNE0oeKzgt07D
eqcSv3LrgeW/39y1PXT4+jqd303e8oZav/4+2AWhairuPBX3cosxJ+NHym2FdXdg
kuLrtZ3L6w/zb8uewbFzoO0NU75bOAZ6O6QZaHiIc6ZytShPDKdh4uFEH2LvxtV5
YJs85Z7T8oMvvii/W/mTxGXaAhf/zrOCBhOKoS6SpbmuymlOGxDd/oQ8dwlBZI0O
LIBIu4NQALzGCRjEsQPdWBFmEHEWeObiNT9hvLVWrfaWq4v4UPGd9RpTmMUO7F3F
I8YSsgRQpnGYRPkw9HdlPJmezyGi9hxUVUVyYaCrCkasj/jGBtLQMbNeppBvd8Sn
+8PWKJTJT15ym8PCFjMKxB+wuiSfT+etY/NL0WtWuRVjuueEJ/Li3yd7bIPjJiBj
Pic6zuMHrnvtlcnAXRVYmffhXhiZjMttxdS17myKuc6uQCR66vJH/6zuPkilhYi1
Hh3VtI9snUAxwlzplkJ/d23s39zXwmHgcOSf5W6sgypvU7keNhDPl2Zcg4PeedSk
1h4lF3Qs3M4xONnnOqeNG9I4YOAl0OTvnXDgn7Kieov05UDPjSYnKnzlUsyqcgQt
QLmjWuFJSLM0SqhQ1vlyjILypLmExUqCfAoh9Q5bENF37Jv2ZdpCUNo6Kw0cGTdT
Dg6/hUEVmXDw+5qkJh693Nol0Lln1qXHcg970L/SqCsN39Eby8uwkya9jcqhTK1Y
MKFtXOg+bQuL/6A7TzO/y0bLaCqSRAE2STGL5QOCYdoGs9Tk6CisQAYXBRoUs1lk
lQZfnqYrihrF0J8NhZDCQXrBBGtLw6p9aMvctbPF0qPufvflclExETE73QsDKp+M
1D8ij9QUEL7Q3/U2yb88T0acNZ8poAP48XxjBpUSxhUlNRItX/83NJPVY8OyIGNn
oGEixeTLD+1eDz6LUghlKIadFv6SdUhcIednh5FFTOWnsSfpQuIi3agHRW/cfmj/
B/n35FQmQxXoxrq990N4TWZ2x+qiUnDPTvMocKgw3prU4T4kU09HrXUlzuyQHqhZ
Y+x6U/RwO53X622NuOnKAn3R4yscPApb02KywGxsuvZ4wosg7vBji3P/K+r8+AfX
SoTjyL1xo8N/85B+TRVzkaRhhHXgVNpRkdPo9QtlIy2YMAa++THLsn2qEBOLbUcm
U2MIyJNkn7+wFXgivVZRwfhr9JyQGHKP+wFkUmPb+3ftmomyurEuu9+qXQ3I4fEo
w82qEy3q/U7EyCD0CSuxVv8sOw8QcoZ9cQJKl/lTq+I5LWHYhgy6OJFZp1NCcSPw
0cmjvOIbiUSTSC8/74PDIJuIBgewGvS1EQbA20/FSh+cXd3F6Nf82JBxg4Xgllwe
Y0TENf6wjH8kUeI3flTMwDIimojU1j7OH5g9FM2DPjw0H0mGauQb34VuVL6NOMP3
D85yUONgZG2M/gBV7JGXgsM1sCL7087CFYEos+TGpJ8fh/bXR1tTh6Vep6gf1KbY
8HnbENbIz6yc5q2WZiEnODxce8zEDvsG/f5TPmQpZm1DuVQn05lhkuCas62NpSvc
5bDQ5QrElA0H9mr6n389AZtfd2huntAEJNmTBG3illbeIzH9QkFDhiSS6hzH3Bxv
ZzJDfdIXazc4Jj5nVITuyxf9mRCZ8NlpDtFkQ/iNi9BZyvPZLOlLQ+IlOk1UT2RA
aTtKOf2L7hJizKvB+3k7rn+XQBZ5NSISJKE1txpkmpQEzEotZRzBOQEXXqyG5ZNB
VvBi9KZZoI3tgKfJmr6THpvJWGfgg8LbXes5v3Mz+8+pUR77EI1veKQnpMyiwY9M
0kwyPhDRfpVUJUxrQoodqRywCukzX613uI7FbobYA9Qubuiedjk2c/hOD5ucgw4M
lMtgTFh+ZK6v99vJWfI4TxtOrhXmukcPnLLkTc+jb3RIXsOpUDxqaaMRydNcaLi7
pa8vbxl20RQsnp//756aOPnAZ+eMBQYNp+6vD7mJKCD1oPhAOcU0bjtDN96n68hh
4l+GV4IIpoiE1C8NT7vSxF429A0+LlKge5Ac8FC6LyJRkEup1rF+x4EtLl11zqok
uO8KXx2m/3zULFyDLi5MQZAKZrOYUWhiOEiACX+4E0vqYanP2LBa3yHbxtybzBKq
V9xSxI4DPA+i/e2EfaESciqukzexyZ05I3WdIhqjNnfuiWK2k+qExDtu+leJUB+Q
Wz/pS6rU173Fi1ybGs67YNBoj2ipswoS0BVARlD4YnBtbBoLfstwla5hQSUZyAVw
yRmpClQwTiZeuDnp3iKC+glKtkQ5rsZRd9RrF2cvjjpr6ziMRcGAsbrf2/a01x2i
1mprI2+ppmHxlNIkbwjxxoj5cjeMPgk3ED8TCyoGfDCqG995sGGUSHvNSQ+YWB6M
hi0ZwTlKMO0dqykk6M5Cd+LgheLqg+Y2PPpKcqM9SAisxt47+mVQ5L1B7fH0ZU3P
Yio5sahS0yHit56O5t9zv6ccqEcDzPKdaEKNF/cpyVfzJtvmpnpeAGgMZr+F0Ksy
MXWhgd+3clVA+04PtYBQ6FoZ29JaX9l39sNE1rpyLSpEnT4H8mbPOI0L1IjWv7YT
FfWvqV7RHpX5Swh2CTdQYvH9Ynayr7iGiZOX8VHurWwYmgrGhnn2F5XEbdi9Koy6
0oihCfWqrCvc81L+BrXIfOT/rc+cmB4YZnkSgbaiRCPszakle+XWCrUnrr4cvq+M
MEpDx2/+Bn9jfr+LLRI3TG9o3K02ptQB24kWDFsH3clhCouohCwo2UBtlyQLXcxU
uo3Sy3ZXVZukGFmoTC2eLhw11q+qlsKOemlCyuleUcEVwECw4Am3HCFvXOmdBVvj
pAgbUrWxxpOIGEFZsBC8z1UVTKMlDseNi/z62VljKGV/8jvtJBUrXE347q+NUP/9
8PO7bGw84bMjPqb7fqWNMWADjlDxHAYLmJVsiXZW1t7h3VFheofQK9es7Pb3PBtV
6LpoBerStBzzRbjEjLeAAQu6xtoA1dM3bi2t7Y8fKJ4EDhHxt7IIu0J3M90F+FKH
yP4QontVM6mdPrDr/doTc7MAVagfAc48msBAbf2CI3/n/3eGIc7hOw2/1CDMHOnr
nR47ejHFE1OngA1p818fVEOitd81tGkXggtUhxUp2+LYVObwH4r/IutMrPXK1HHf
R/+os4IANQh+NVeV4xYJ4hvtTkTZ/rmMou/2azQ/zL5nt3pQ4+QB6H8CcwxDBcUx
SOkb+QFV7t3hNnnfSKJZ8xUVp4ua+Vaf5pE/WwtPHYVCI5Fr4MqCkNpkKQ0dPy1B
5qWMMUEaSlyLKV+YNch7paGos0+0hRDl09Jd46vo61ChAHKyJ5MLFNnlGPLRusd/
18sBlj2W7prP585pM7JkznSkBBCmWJf3KQFIt9YY5V5NuVpdsmDogwpA7VuMrTtH
jaPFiq0rVkDyQYfJlhsBfwEx5cyY5hRODiMUPThoUSI61GpV/9Uwe2cqbpwXj866
AnUHnHAchn3kaNQjXAJmwDKNgJgsGWjK903VwLyaUif84g+kOBG4nxoISOnfKYo4
i82Z1O7h7GUbhz8gMCww2bmTuFta3Hs80ZjlyU3cS2KBMic0rSV+YgA+Djc7SGk5
V3TlR0TvObbAelNa6DJx/bMaVIYe0DnbOZIYTxBMDVwy/MFkkFTEXAZNhr5dwPZs
AWJMK12z/3U7QfCzpTYRFxk2L8VvIGTeD9HjAhTGzTMwbI3kzOw/J0/N0igkNhJL
yR5UxjfkINyunyau2dRM2Aos99F/HS0A9bTbUAJXaFyaUk5Zp3BA72KwSw8SAe1e
aW+6ZBjGukWhiCBwXYkxD3oXJOgM5VGx64iV+wxFKknuk2wjp1fxW2a6JyDCZte7
aexuepv+lssjRVIKJT+1BBr0de98qk0Q3YZ5pszYmswNDdYEZn/bMeVt/1cP3tRY
Z4s+B/gy+BPi6TpXsCW+RNShaL26T1avwnlzwHXz9nOnPzWzsyASla2/nEhX2RDs
hsi8ry84PWLpVpyShaYZGVqQ+/LzzkPUrR5L8Be2z2CGut8dw2J1ed/5SaXlxvxX
j66tX78hTbxymkLvE134+bcYw51c9Abs2qyJoaWu+msfGLSnXTN/5oe0vO5UTQcM
Pmyr3mUvqriwB9q6B3ya8nEDGVwUbd9O9KukggbYD3NRYcfND4joH2fN4DEgnpNw
KBYlD0YaEpuR5Ofzqr8WXi3+etvyujcmXVUauIkTCcx2BrnFAV6uD57IzgWGzSNN
9QesOUHIS03wST1Ai1Hjzj5qByLlQZU12hquFPcl9LnBUMOXc/0BIL7/kcvaZjcK
oIf1Hs6HE5Nk3usx7JI8Ag2vleDyN+eKG0imEVhl0e7ImjqPRvOP0bHmnhD2lrI5
VmkC8UCU3vrlz2CTXI0npPB5jsCwSHVYQhEBw/HLgqJZ4DEEybf8bUBGFE8Rp4B0
GG/OS8AvDzIi/SG1UUh1w0r2iyWa4/nxRTPntU6dBhK0HoCsi/jPlWulh9W0ALhM
cHXZ66QVXlmCmT1N5VRAxq0zMsYqc7qTCOTYQUVKjxKPy5RjIHAkUbCNTQUPaLzH
wxwiRNNu2bpeNvasjbLRkql9ECBjYbsiWr7cPnLh7ygk1xKUJU77Awx8irm9t21c
SOyJeXQUv/byvTJyINgQQmYpGgYyvVAHXNM7Tg4hruP1oKmcu0+I15wdBukEFnq0
igbd5bW+aXOwg4g+bIwwaDP745sJux8jq9biurSf6E9Pbi5QfierSyKrSvogvMfY
RDZzX2ySxknP2NDn04NnfBp3MPjcdJkv9fTFuckLLBQ7hxnunphyLB/TNgolNsPh
kBEITIUUsj5WMXfGorAaOQ8LkDroro8iL3pIIUjgv6YGmBMjs8iMS0BLuwMZe8Gx
gcFj5yLeljwAJm0E0YynyHLN+NxqTOW4gKBP1x48r7mBuXaKt2/5712sXpUyQaHO
maNsF6J52eiQcU5EnDomyRTWHYZn7223b4Y5clChYJq/EGKBTMH6z/1UIx4tBaWp
Ps7T2kZxRI5PKeDkpgtEjBbxyyGt7oh+81EuDm+GX32ZPVoV6hsyuNokJxPIT6C9
qqvMIU8jG8gycmbohCEagjwBx3Zps4v5q+n1yzr3KZJrjttuYo0rNJZF7KBhQnEK
QLIHvLvo7cK20P9yqEcjeBBnpasEYHwe/kn90ybiTUt6fIRC9T/GpI70P7kXqsuc
leEItsyOCSzltaTLsI1+HKiu61VuXNmQ6ZXPLhx7tLY5JDdk7XwCv6I2Qf1fUQyz
P0CYVVwC+pqf/tx+oes/DwkQ3uDWxm/0jEx7fc0hjRnoCQun4tTxL9F0Ot5YV+9x
JsJMkFkOsgNalXIC424T+EFXpF/8jVf51QNiW6tUXkkZ75T18GswUsuJ0zsj8OXh
sI6v443D6vdIAfCieBwr7RpaRs8RhFayPJ6Xf8Qfg4O2nxgDGSbWL+cZseQwuC8k
okaMmFx/sl2ZbQ6+zAqTvTK+OWG8KPcAqaqhezRLIFYC/+ZpAg+ajndgZHVf0UWG
LukZj0N4X5Q0BVlCGcOqd6piUd9NY2XU16Oc7bfUGKZgq5On6tAxrnFuKsEaNA4g
prD9pdmtkSWHiEbRSC1eSSz/Q+Ercerz+WhRZnLK6EWNpstSJ7rJHxT1Oprrx6ZA
/7pziFKR65IIEMR7FVXdC6axzLJrHE4lYcLOXIH7VYXwL79jZPaJv7pzl74v1/Qt
ZTXPd7EicltcYN+lEeGBtDtSmRTHVXuCrXFxGeKBYCeejLaVnQvIbuObHsBC99r0
QW2VfjwCumVCplWts2pDe8MqMo+WA7QOE/w+O3nNieaC2LPk+o8Srk6ilYxCpZfO
ONJ1czzDhNtMGQLHmi9tjVY1+feYUkVGKg8K7xovXMbICYmz9RyTXYXezhopcYQS
+LqYwpf+9+XlIWQVKp9PFTMjH2Rka84cbK+Kgv6/r5PhK7ZnuZObFrecEe6jlYIX
lTY5b1B3GWRUCFptjze9wFlrTMA5kYPWixa3/1HpGlUiRYvEfnC5mkdcCKPNeAv3
tRgkB7IVIFaj2P9ChkHV4gBx6SV6HoJ1/LiG4yJwWMbUv7cwtVVg9xXE6cEPgkUS
10YnTwhPKJqjakjai1IUyBmcjqhMUYdCQel8twTWhDWA8SjsfJPoWByyIGfltkIx
rEPUjG7c4panlOTtvf8IVAh1DqAMVrZTdOcTVOrq0BX4GYCeCTL2yQF5dmVdZ4YX
/j7tovXdx4gQWavDgxVpiHj7J8QvksvchgpBmkqx3MKHsvGBXunvfwGNktVGg/YH
Gr6aXg3YBxN9iCn3ni+lHh0TQd5GXO6KNBJz2k40qhhCEt5JNT6x5PIjbJpjsIjW
7L0W2e02j+GgKNPWVakhr0otd0cOnB5EXD+Y9+mC2vzlLQuJj3S6/u1UoaxkvXjq
IiOBvgWPZeOa2jDfTd1Ebswvy74d9vc62iO4FIA4n8Vl/cxtl06QXoC5Sfj2+yGr
OdhmcOOPUXJcArisfN+zIKPRsYR8UJzEkYZNN6Vyj7k/v9Nx4iCLLLZIgTfkb3xP
/p4/fNeB8LbqPaTWgEGxic7PS88z8SkT+sxBqllqdxLEqD2Ne7d6P9Tk9lsSo+jF
BtSDo/BE1mGQgZ9wb/0OYoVvsV0WQIMeNex1siSIE6e/mKLb0hgtVvj3FL6mD7DE
1w4AAgYpPx9Wix+7XyjN8/sjp3YZ4gbBDEE0YXRqOCpORXO/l+fivL1L0KxMgiNE
XPV1/gRvD46IUp4cObLoTgHFiKyPTGTUpjnydCq3SatSD+G3SFZ1+dbPiirYAgbP
CsT3l+OeXVKaeeubnm6j7+cR5uzwSDTw9M1rjuaYRbhLC0S57Cyv38os+dIwADlP
2CSaqh35fH5kkXTXr+2fZIbH0YQTJVF3kYGgK8vGFjvsRgLTVOinakApTBK981Of
iw5lgDG+XrGjIb0kf3DjZrM3rYUU9aXb+MiZwfzaUq6i9PH7NaSBzXlHoeAE4gJ/
M0fI9OyuPuFsxsEYAdWL4ZnKLpe+HwWiOh+bYsip3s1aTjTJCtSSYyfr27xd3Ct+
0Qo1pbNDLSbNWN7RyTBi1aypqOjTOn8Atzbqj5OgzQIQJ3cEbddBodAJaAXp7rmv
HwVg5riZEhKx92SkiQ5ZyU27b5zkOpnuK/Rjxrjt2tc35qiD67uVAOaZ4TwHpRzK
ZsawkrI/gk9tukxUG37SFJIwji4AKLflDA0BOUgcYP/qZfWFaG27eBrYEq+8Gv10
8oPk56o2iyQfnxU/sEXOs3KZ6ajjYCqwIdF3sd/UAa/j4jj5D0PsR5f8xPJZVYhm
0lK3JFMFmY3cnctAv9/RaCKLPXh2Qzk7kvcI4ZFWswFueMA9tGGRxaqBKZUPIxjq
4XrQeZjCkDxZEk+ZdymBRqWOAY8iR2yDsN5G/47VM+g4XL2PpL6+p5wZgaiSjZCG
1XiqWhRMmlTY2E2RWGSMkgoxuaUZ4a9TZ+su9lijwbd52/lpqTfO10bh0AFVz1/D
Bom6N4aEk+fvaOHSjcD6rvvIIi28F6z4bAeJJ5UlpCgTTfdtzf3mrv5PkCffXzYT
4BCCjOpWg3x8EQpM/2TUJA9V+Ck13KEcrdlcDL9Ig+Rww1jdn7XYXUX/X5GIKNjz
QjEI2myTdV2OGJVHLEDZe4Iuin66MGIjsDkhBKMXwzPq7Bc0Pk3/AaQwmD/i/edD
U3wQ4GoavqWrIyrNrP4W7YLk/GnYefXtiDUd35WhuibajsQD+bkeYCRCtsUdD9s+
m2z0bx2unaEuUZJ6DVynE9CLMbDDI1s2TbgN2QfkOGvqtD2P8oQaTB8vPa+HrjXO
DiMpd3ZeQRTUcBDAKrXxTEcCK1NPLm74NXMy4TvHD3fpqYEpbqGTMbT/jLP0F+7N
IwLEKhgL4S23oT7rSJKGd03qQwoVaqgTxoCsCj5+hFlbEsV2x4OwZmRKFw4RD33T
qRCAtNG9fjrPBDpuhXlfDHNTmffAVY97Oeu1anrVFwXROTUFVBReyk3ZksjwKVpn
6iwxhE7T/YN3Pt8Tnq9Yd4bKGLsIDfx1CUXL+5LbW+f/qixNchZODtP0fjZEr3Mz
RiBI1/092UPhD/s4pesGAho8GJ+UMBgKpRJFjLK7vA9JMiw18laXg2Aay6X1VZnD
YXOSe0vpJEyJL5640GMB39J/ZPFuQ+Eb9thA9VX5ow42/0s1+xPAdNaLW9pefHWl
KK4XT2cMzDshWJl9Ea9IVo5BdmnATafZHLG30EiZ/VcWM/f0CCUgLFk4ehZBUANq
aCzNcTS2IBauTQp4WIKAdUFNxxKu3ungcawp4ivtKicikHxXns2yqqyl4Zu1iv27
lNxayeFJwtLMk7yh668pXhYeBhRXa8PX8tCJuOJJ/69ykgUbk9Qn2fc5wgc39yZV
niTNxtTBJ+k8c6BhmkxOjYNFs8LNzx/XGQmaO2st11eRhZnrx8xOMpeeHhI+viUz
`protect end_protected