`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1648 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
HdytKcppDjja7VfYQkCqvFU9qCX4kdJHjZV9u2qwYZiuPyuu7IfIKBnxcchOYMrZ
GjQw3e/y7I9BtBiD+rsJEyrJTx+jzuxXcIcEqnixavqKtGHIeYP9G1mLY1qnyZTU
RDkLRy32WUGg22ELd84+5FxjMx/AlO547lHIWaL1GxrzSCvui3E4ZjfBhc/SF1oG
rs7rNf1ZcdWZ4gVbYODlttyCqzX7K0Fyy4M2r/kYhqbAP8akP2W6K+HtV8UeLLee
xjZ69B/I3+nSP3SVG0ZcV0FYFz2CIeCR8dCu1161SZcrP3uiqZLBHtVTJSajWc2B
VeKTUW6VVw0kt60S/2g7I3K+GwyVhjkEDfhMagWDq4AmzHoVmuvggcjdKz2U0exI
sTN0vWWqJjM1h0L48Kc03mK447Q++OTYBTlnnH9qigOHH+HbbsnC2U0+v52Y7V6b
T0ZsnScHemNbsIi/h88M8MwQjTsxK8T9wPp177gf5HVj2XDVMaKMF9C0IxHpcFUU
ZFO41F0yk4Qp1DRAj5MTRwBbPJWpHzab2cvgERRRKY0FGra4b8ogozsIzENgs4+Y
sIv8PUUBPi28XIJlaSECKS7MdOYK/Z2FHhuqFWAXCE6InfBEHQbpIh8+xdP/UKZS
6fngyLmR3f/LNSq3eAjLLdrLzyxYcOfRih/gXWaAyTnBlpPLX2Ytmxz/avtDNFt9
Z+k+xnLw4QdBB3BC3d3QMm3loXp6x9Z8x3HJLUkhj6oxik5zJQjJTH/3FbUDaDpk
sQjI7q9oybvjk781NKkgnnBFF0r+45zcdv7cdQHuIc5c/YxF9qbf1+HNa+BdIRmY
hRukf+2/xi3rrA/pXPKYSa1hT0l8L87Z7uZxvBxCiJzbydWfns5GL7bPR0VtSQ5n
UPQJTzonLHCiGGGbkJchVIM69KC6p1AjoEAVoof5M5ZGrH57GmelvosPysFNUjF5
UdmMgvJjSEeVueM5drComza+d8248KmJw462pAs1S6yoSPGE9yT/3ps89cSZP5Jr
Yy7inOrRyYEkbZYgQB5ZeX8d+f4ubQ+43F7LjF+s5J1QvRp8NOEVIXBzKixUgN0h
SjC6Wjwh3lEp3yKK+KvStIGFJCe48lv9+2UQon4n3x3bySyAIivEI4H4l7f0rvgV
mlv+ibesiVX/9Z8EpaUYHg1r4F1m1JxjVFJEdmhOTC+FLwKQi9Qnd9pxaWyL+MEY
cVfq2WD3WDwiutksfZWldwgcqzRXwfRsQ2dPJb1+U1kpm0N8i9WBmw5nWVQGAHMO
MOHBVaIzSGjbeJyNYC1dJU+DN2quAuzaV0Yc36NhjJ3ccgVV8tBMdk2hzEXglAIE
CWTQMLxm4NLq9qRQzsAUtLZuP0YB/4A6rKoIkT0Lc4b1oxAeORzkYCEH4+3Xcb+H
A0X/4cezr8hek337anL24UnewZGzeVMS31VrIinOfwIQw/qL5HM/B4cxUsodnHvr
5PEQwcN6R4VVd19B6EhMw7iDK86rl7LAvQmseeodlBADcCebOxe4LwFE9Wp6nPAw
H0elWI2wSkN6xAV3VxCEehtrruQkwICbcvvlGl799ZbpH8rmokijo6qCs+2WdEdS
vpIofh0nPEMq3JvsNAWzsZqQarOOYbDQQRz6F/Lq1WWvSvuGeRtVZcOhpJfN8BCq
g9DGy2XfpBRU+yNk8TkP0m71eHruCn4Vwjh0czwJrGnmvwmtxnRuiqC0NL8lce93
YSjuqY5nDcl9AhO2wtl0gmJo6a8807ChYQjGBjNfLvdl3NK3sUZ0cGfhhJEzit2g
I6RT7Inr9u/bAvzToWom70AXhGiUeLn/qByiFGZ7n//VLloxPsR9/1Otw/I/RN0W
KGsiV2VDGmjn/5Rf7FgYj0IHXj5/IGN99/OnPG5pnWjm6Ybt7tkqdgvl50u1d+to
IRb0iZ1gvK/RlHqyZ5qJLxf+bhCmJ0X3Y/tmXh/psXBHgRuR+yik/zrtZe9s2Zu8
/CuN9bplwTBSHhxVDZkxeQ97vRtSoknJmYK8Kbv/IUxFqsAQH39bdDX0SIULALIi
BlQoTOK3QRUBnYU7dkJ1Sg==
`protect end_protected