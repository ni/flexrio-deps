`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 41760 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
sTHDbAcNdRVMi738hx0vztNGs0FQJUM8ivjVMxQ8/AQGgZBGH7HgV02DHDyu9Wnl
dzdNmSlB5K3kcF0CQTuJOuzaehWMpV13bOGepBhRkzpcD15X5R1myU02hKjJ0XBU
vCK4SbEuV6pHUl+WGs2Yi+ZkQh2klV2qpMofScUF981jaTAQDF0mH6dzerPXNfzU
mSRIg5gBecTvUGbXGFgYuTbDer3CLJykhaXpgrGSEPr+8c+nUr4fjKUrVZVINgjY
egvUMT+9pbt6vJhge8QygBBb41gIyHFBEzqaZXknbANGIZuq9yMvCWOl/RDbhrFR
TwO0y/DtWYhAQS4A6il7tLcdhR1d0QfQARpvAd1GowE/5krAnGy0exTCbBHWj42L
D4uOmOPbYJIMYlYGWoeUF5l5LmGSVMbhanP3EmJEBYCedERlXee/PSS3oz85JFbW
f7xSRhu7Kt5EFuzOF6dNIDC8NuogWFypFHpeah4ZsyqBPGxSSyfD0mtqd0UYpCpi
DeuMsuPug23uU80qvTiCuNXg8u1wF8FDLJQUjmsGeM3hv9rbLN2u1qB+1xrepsWb
Br8Ars8M9C8Zmtj5XgfQGSyfLTM5IptGbUFXkNXhiv/1S3xPhNdmAaGOAlsW2n1B
0K+CuM/r67kjl4j1VAMUakfuGlA7K6iQc8PIBy6v0Z/uSyJAxbNqD7eS4SF+UrMf
wpKqzjohaomNNTprL4U6ALrg+Q12P+7c6V5sa8Up5IGrHeIaaxyoOpa2RH0XHCa5
l9QTBXozL5TrXqx47sjnYwb5nCfTD3+a41RcXcdOoEXaKsEWHSCVLDPijVfsJIl+
3pq44/J9pzmNydGGgapLL6JrTuHUmBaZ6MAOyacXqtLPboqsvbBGDNcEdeiZExpo
RrV2m7xoprUyU4zzTZaX34CKDg2/3A/X8KzMr/rbxwGMZXLx6qdY+YENX8KURw+y
Of4CkgqAOdm0du0qWl0phwm9mOSeyY/PJMGf0GD6/HBg7hPyk+QOiNKB4C2YbFDW
ltoRBhsVMtUDX2bkaNJFtxeK62rKkjVr98IvNIWvGa5u/VT47GTzoY0qiGHmqt2/
4itgVd31JuGOeSE05X+7UJ5DHGlkWqXPNvMtscvgjVckEKbxIjuHEIPmiOQgxxZy
8RFqneAnGX330smGKLBijlVkEgpo5glK5QtMG/UxtzhdP6PEX6PIbeu0tkwz6E3Q
BZlMkvgj7bXy7u2Z9qblxMYPByoCJptHG2QROWPFu8G/uqhG2G9lA0LCy7HZQult
Bj6NYjhde7F0YOEmx0xrIlC/c+S/jamLfCHIqk1h88ZDZvH3m/+7XDKBGXn0Ieaa
h3SwjP9ym/+MyXDY4Ta+k24Haad65uAdHTA4sRuDhCXvYiKHo21UU1429SUSrTHc
wyCp/u1sAFXn8G+67vPZHqGtJ41V69g5mI2WW3r4QRJtEhF2HVYSoWkyfgwsFeZM
9QZO+QB9dpS/Gk35UXimM8msSKpqUjupscc2NMui/fmq6D2mJsW6z659xg32+rKC
qB2tq4anoQzqEUCX1zEK78NpuVdEAeqCX7zvFqOmWkJzl4yv0Kj8G8/l712SgFsn
bgmyU1YOnmgi5ZfxENb00FSGB92pt3wuJ8wh4niJ2R9Fxmrl8QaD7Malxcgo8iX5
z7rj+guunUBgnJjvHVK7qYFr/BOEkJNSDX+44yCvquGFaOJcunkzy7R/fkv77/+Q
2mXphogLcIcebfHys6GNTfTseAakbNhRlJLQm+BpZ5L3TwomafaPvmoXTPsmgX4A
ZWve7nQDzqJPjEhr24M+7phj+9+aUiADd8JS+FdG3BQlMKkHAJTlSDtOvEtBOWpF
hE7QHL5ouhUu5P3sKWnl9w5h6okHzhcv1CQc68hR6hp+BFX89lOpa9pZDpZaN87k
AsOj6QLT5dVPHuZAAkVlILINofY/nEbBMcKAugRX+OKsVAxIfceYqm08GK56oMeX
bS4EprmXizGsAOo6el/Nb0bg1Y2dB3LZ8eJ6bWsGSY2IxnhpZPcMEWs3Tr5pFu5F
rlxotolLRtvO3Dxtq08LirPbBf25C3C07uEtTT8R8wEWk7ME/B4vc93J9rGpLABu
d6pQTvm35pvWYsfGVFUbpOG/8UB88Z83gfjIa3gjp6DrFogA4wPew4I1ZTIiwGZY
9UUHJWUlM4aoTsVytJ7HwhNcc0EVatwNvEAwAM6UV3K8dktX3il+cn9+taSDFzOl
lQJe+Ep1TQENwHNfuHVdM+ssNWwL6+sBIVHycwq0NN9rSKrhBmpyCbUEzmyjb5zj
be/dZYP4Q8ux828KHsU0thQ5vctyDFfOwBSYqLTDLVYmXAS6H7zpZJWZe4ZuXDtZ
40lwP5sZH0kyKooSDNdxum7oACFPU15wLUxcyRixNvbbeJyaagr9eB98vH6VT33L
UqCGgfyWuQI6ojqpnvRTGMO56JoZdohdTsW4JYOK62WU/R66Qyod9Ynt0Wtzke/Z
xx8cU1AE27Kfhe2M2GQnxVuDsJFfQeFBKwfxl33579FkC9g8mjUim3jSPy6INMmk
4gxeG+vRPrHKOtDWMOr9mlxnoqXrKkF5zIxX73ikqKk+di5jcoPSj/1JDaMpMIYk
V9N5zyzr0T7XwiRJXb8dIAMVFHppCX2Z+AQX0FYdZcSAr0TbxlBu/lLPX007ukFC
x4/wmM9TcB9Vitclfc9N4Sh4jF0ShgWE3rIZJLWemAqGFErUiSpCNefalLIdCNtf
+tj+oZxEULJKMzxUFtfgwqKU9m/eEMREPcFwEY4p0GljPPbTu1VA+XphyDoQG7NX
GD8X7jXgTVVTHlZBnePIH6pUIViXAYTlDWrmrMg9i8CPIY0zcaNK3AvUPS6YfQBQ
puKXeg/6BrU65UtQww+SA7XZ5J214nw2QAk1+vHr6VsmH5vK5+Q5ILvyxMxlpPDa
t5shBxD/A1L+pghTtm0bP7mt/GQWb6s35k9ImviaM4jNg7EqePIGf0XNs9nzzSSA
rQo4V1QcJG/rxJni2Da8DsiOBEjHYOai/2LJ9ZaE8rJ7e49I//jZv1LYApiwg/D0
Hn0pnwgelmcvEeLY9X2yTCpQGsBXIvS7azBrCj9o+Wq1hzveUkdlwnuF/4+ZVVow
NFuPCHZOlHUBiEDkg8MvU5UyLeU8pduFHb+OgCvnEMZZNNf91fQ8bMGQs2DHSDhz
h6I3GnPQUW6vIdVvS3VCb+lm3vIiKYWXftNDPBhPSEaYJEkn63MwT19CVO8vgtr+
mUQttLO9qNrpvB/noKFc3SrunEDxJXJgR5MRZXgQQE1GTa0hM2YDXnz/qzsYxq96
DiXMfgffcrKIxiskHKqUO0jXux1aI6xFdgCUbtyCN6CD7Oje47ko0hbCmsMG7nln
W2Z4GDV/8pibaX/Bl081xB5jUQxzRjhiPwMvBgX0ZAhYJCOtw4IhUa2XbLGMVxNr
vop2c5mraEp+Rer7QNEAVMdOjh4SjguyMrBqjwn07uQc2ZZ3J9/9x6Md3+Ea57+H
M320hg5+2Ydu44NZkO00zmHW8KGC4xeYtDYqdAK/iNHhmGQuSAZAZ8o1FTT+OqIf
ZFMhpBImRasIHEMfSOyoWy+zvo4mkKqYY/owvWmV801HW8yA5pL7KMncnnyhlowE
Mde2kuUWxqAkWAOkQ3uhrmoCfZsD1FWVgzZIPK3nCpIWoU1u3VHO4T5VVofYmaVm
Z1TqxzRA5L5/UrjIngc0YNPDJlO2Ix5mKMh2Y/cG993GcZ090Gy2JeMb26GvtG9O
6qQNkm6hQgq2+3R7ZN+XCRaX4vCzBEUUrroVTkQrp/rkt7lypyNHIEX1oKGUA6UX
NuXxBHrf4f6SJbdD2pm3cBCeVZ6lBGVKA21hedeXB1Cwu9cY6yZmhJWCDZPReV7G
wSPSEwpCDJPRO8IqREx0btX5AvNMp5xB3IrYlfkDGkqt0WUrSJe0RiibWnrhvHrR
sQJPcIIMtClHDxTDc6QFs4Rr6dZocSsaEeStiLVhauqZ7SPIPxcdVuFuXFdBwdxm
t0/cb4ZWO6AQybROkFU5e+UOVIyTHBwtQnIO4hY1hKexL925HQWT6Bked5qmPauA
wmMYizk3CJNSWgZ/3yH+ddyWRyYRs0ygDsG7ZlErV29yUf/PCF5FXwrWLyhOe/br
Zzw+Q31FxELiFgN3uWZ71er0BIPVbcdbM+eS0qgoBTXaW+bmq4RHV/VswDAkSmUa
JK3NOvfcgAIlRMLPm+LUF5jIp+4GSuq+K+BdtqAMsu4LjF5EVSMTCAPrPvnFgGNP
RggZadL5P/7hujzNvey/GUEWuagnNuLk7bG0R3dZMoC1Qp8UdNgsHVd7FX9Zn8RR
7v9lHKCkIoNutjBRte3eXQpXD2nHWRoLnspZ8iSF7ZqFqnAU7OxkvWiVJIEYqwZR
4kLU7ONSBaOMsYjmDupnqt4ohmPG9VZXsImawkjzj1Ejo0oygk3FZuSKp8Y4bi7Z
Jytx/kggz2es7VKaRAzq1HhheHN8JbAyEU7n/42K4Vb3E28PZ6WmHkTjIGIrnbwv
H68PIcDBo1bGxtBhS7/DAvy/FMYRsfbWE1qfmMjVdE8PaVrueLQGp9FksY2JH+E3
WoiOMreZqfJM/OfHeWDldBH534VyUWr2+P8U5kw0UmYl0Pdl8nlUjrIc+rhgbaI8
S+Uygy4l1OEk58DPNxE7imbRLgvK0PtA8O0zzrTVIorl4b3u2Q5UXQMNv2gESvj0
AX0skbDUX7pMaN0NImex0+K7XEeLFhz9b019+1ZfCgZozlHWwqft4gSeE4genfQF
WSw+IWkfvE/YEYZ621R8wpVq7jPjOnjHc3HXgv2fEo6DELhYS5jX/JkFoCp3wyTq
AkARMRhAW4TZ8UX38gHsVd8u+nD5c6by4FA9ulK0SKBL7+mQFohb1riQ2U3sVjPY
jR/pG62xLWgiOOGi8+e24qkenjyaCl/aPAZuUOZ+1xj/9piNNWoEm1XSKI90UJ+0
meeYOmf/zm0vWOsek5Tup/4ToS/FfsEJWgVrWZl9QFJMOZlrXAG+QMuJ14s82cyq
VFuXNvVQ+1t6+CBccyS68K1HzsceQt9PGfRscMEDV2DDFQifqYu+YRCy12/PmQBZ
cCl2rqCjbD0RujyX6l6hKXrx4MuRaf/3htj0+DvnaeVKQLpkess01J83w1iChZnd
xHiIt43aKivKduU4cwnHCnZkR3sdvlOPea0/RRhXGuQICRfUCN+8h+tfigsukswn
kOBOVjLSeN2M62JtlEeHnErrgWkEvVV4tLtCoV5qpFEchq7t3rEI6DRbrVgvS/qR
CcIyshimTWiJDIfGulsj93utuQ2I+Z5ZJvQAdCn2pu/JSLVSL4qDV11a2WyapxX/
Fr0oclY7XQPndOMfe8yOXUEXJq0qUNdtjtw1tzfWuv1OH0xeUUbwBd1xrcFU1pPw
h5vrNgMoQZjX6QHwscAz8GTgCjvwZH81fnUemMhXIfi6QbiF9/IJ+k8zf9h6k8wC
cD2aKWs6vqeJNSOOmnV17dXFdNLPuu40G7U5k+VPiT/UneyJerVxSomreBhzZYDA
WDwaj94SVzlcLL8pgCoIbMDNh2PMFD/hTaCw1DicZJyNk5q26KV+dWLWeF5hOl2p
y7C1eVCWG364WRSbRQTwD8jSXoHh3wh1n1pAKJd2rOmTwJQ9ZsyFHFEkuN0/B6ju
vOOw/AUJwirnKB1D9+QUytNxRVheVjYxnTgdyvEfsw4EARn/BCNmDXfMmaMxWJh+
2jxzY+t/APSRO5O8d2rOdlTD+Txtei2DJUCBSEeroLhPE1/A5r9V1wxrK6GhL/BO
TkdtvBoESKS928mPhfw9MbNLiYpb5lTWpdmHWdV+CIoP1wvQFQWrwCbnMTyxGOHO
cGYYWNjxjaJG/d6CyVoYKqX0jLP+8Z40g/QGMM2p5jiDwXZGDpFplGiiEG1lB1p9
Oke4i8lNbcgjY+bcNOhxXAY7hNSGVpV6e+HHMm4FMofjApIcfL07BqwHu/tytzG2
Byfu01Ypl3e6PAr/fXUA1tPGnTs0rO6clUs1n8I3i9qxJTkJT2Fb1+R+Jzi6jhv/
6SGQsmvTSaPigsg8kyDTEWxn4XbSAgvjwHWTmIQm9g7iP+6+Yw6johck7yVlmK88
MOXWxzZP1IyaxQvmvA2/nkfsW5PryOOjC2cxTlK1V/J5B1WUq6ro9gKv4M6VzNoF
5sRhWQ3A4+XIJfomJq694EOdmS/SIaE9tdR9wHomzpyqpoo9ZUgX+o9bKAa5yL0H
uzTWl0lLcuq6oTovN9M/N0XkSHIBPkBu/nuVKJicTuylMr8kX8tcTG7kxue5aaSk
i4ytPma88Wv7ETmWIz61/LsMWjDxByusV8fKDitt44MT41toDEKTA+9NE53ZvmF3
dqbAZanhsxIqDTMngp58NHmxGMsjtKAZYx4m7zx3GPYBJapj6rSZKkyWrVBBD1BJ
TLWLMYT9wPSEi4YusJL9Zj+6REyIU/BsCGRssRfr1EHRx+VX0y8/YRL8pBqlKfik
11KRJ1BDqfdjJo7aHuHdr1qvDk2gYYI0WHEqp0ShzRCQCp7y1zvisSrvsclSd/tN
77QleTyR8LDK4xffw3O/Yh27QSBAa7j5fiqGvG1sQlYJjhbD/mqrFZAbGMkuLEwI
RI6sEqjl+8zOHXrvxpGHwdKdzU6bjkwQjIXq7+wlyWFYsrEzyHPq8PG8CpbV7tVL
GTlFMqO8puHIHhziEOPgHriLVaq6Q8iP/DzYs1fXn3kqlRET8xTW1Y/ZqOoTpem5
THCcovoLq1mggMOCY0vLCaBlp2haEpZK9jwgTg/gStL1zHjSB0ofLAyHYZ+jbJk7
h+yhHIybGbXCS+MBJDh0mgIDP/joXXqwRVKf5acfxkXTKxPFF/MoIf+LVdx7TuhS
fNFtSaxLEdjO+GZp1V8KVn/4jj5Mqda8MpcboFtnW91Jq2fQNkCam8//Glk/QrPB
IEAgf26oR1mDtLl2gMmdDlHaprq0PJjg83uwv+ndsBZ6mtgLosVws+86pcN/VvCM
hgZEmKdkTLwSsoPXGKC77V/+oMqoL9bVSDgiWdxkQDCm68iB5ATE3kgQy7A2Z5J8
awB7HvMLmD3D4AEbnoFEsSxJspE1U6sLDSTtjkrN9qcpGfk1sS/IeplO0DbozBV1
04majggx4nyfOFXmaTOxSu4gcZw00Df++cm2xVXKj+ITNBiS2Do1z16lBconDIHG
w/HlJq1uikFu9dA6TqRXwLhRlKlN8HZBvgENVQEE+WmFcLsVF64JjJO6Y3ar+CKH
U/ES+XZt2ctqK4fQlDFu1GvCL3MxzlTOjPfLwFHkCRwqFgerLyydt4ZjmHUubmXG
BlrYij7rwbDG43WDzgBVl7vYyGUPWstEQhnUC/BZM3FjSIsduJ9RQBzMIHnGM0k1
APWcuOuq+64iVT6dJ+W8WuFO42jcH7wqUwMbp7HpozOJhiaTc3CcpYIXs34zckMv
010pGraZqtAuplmOAISkrhEgCf14PM5RwSpVFAX+ACLlo5dTrMxpYKqF5H1PKKVa
utC1n1pnC6UumPo0lzkAkfhrNIsD/irOQKnmTmjHcETwMBgMOnhC7+FCFeujC18t
tbvPXgFGtJeZ8/jH+HPKwsPLapvf2v/GV5Cc3CXc6oisSbxwBi0Suge3nqzxi5nd
VowkygWAHU+KpSPpa6ceQxcWPdpGhXi1+nw6HHGFAGoHjcSAxbxCDMts9nJJIAi1
LoeFkaddaDjYeFaXocU70KW1Ve86B5SuRsjH6AA6vXAjrTMq5GscIyPaqrvk94jt
SkBP3Gu8UWiShf762k5WnYh2TCJNC6gad4R2LloJjD9x4ytwI9fJZO6795Huv4Sb
H/zgoTZ1RUcgr0Jzl1hdBNlKmF3GIh8g/WnYzaWHU3deI1E+ZXd9I9hipNpsJSO/
WF1moRxLQMRfSDb73rrBKglKZpw6Sk+avkmQ/KfgeKUrGQ2Y9xoJLpXsCWYetW0R
dmxA7p5ooThqxuOHl2j4e9jjjf7ee78qrl7VoHERBcOk0VibGkkrLWrG72hkQx3P
clQCbL1Cp1ZXawcM6enylRpWoaeFbaaamRxswWz3sT3fnPKTTGhY28WO02e9QM90
8T5Nq1GAUhvnKla13XLd4CoukPs4FbpxCE55ABRc0vbTxrVVT9oHJAnDkhVGpQgU
7C/cnzksDBuErmLADk7jAfvsUgrkjNQ/kvX9xkU3s83hCnetuqGSMs+IL7DvEzQt
sTXEH98ytHIvBukyJIbWgbno1N+ExH6IMBEMg6P0hYxTsT4d73hNHdW6aLMHmeYR
FEPKNl1UlMp/XR3h763OTwvJhNPKToJjXKZVRvNyxFA9SPlMQ+I0EYDgUOWog9z+
H7DEFaPu2qn1MCegxnJyk9XsAD+kCU2osWbA4aJSHxvWSFAmTABJ3lfcs9yAB4uL
VMAPck0OwMRfqrnhJ+z63ZJAecvybl7MgbFnwoBWuq5Es+5wJ9rs9zurrg0abcRz
W3mb3E4NQTxqIFLGrZErir/DGw5ZctGWs+L+YJcsHa3aWPaLib7NzcCIny3YFRBZ
n6cA+hibLU6jiX5XOpFdXIcSClaXr5+kresXLCNR/yx3KtBSQWTZAMTTTM89Ss6g
SdHkQtsfX4tB0a4mmDU10d8tB+ZVuHTu+Enf7gNQWpRAJx5bcWMx+1atGu5gtQ0F
3TjxBAw4GuSLVvRoQFojBtMOP9mnIGF8jrIVYf2/qUzCqKs3GKQTs9AW7lnZQMTB
QXlLZIAXt9+wiatZ8Uy0Njvk7NNEonp2vmbGyWeAEwrqfECLshmOSr24xf2RpHqa
xiYRXMtVgKISOz040rYDhAG8Ium9/4A8T4Otyfr4p8lYlkiyfBOlHnTu6Na9VbLJ
sM0SmfKuBLQev1+PNq7HyPtmg5e1mFSRBda3NoxyixHsN1Veto7goF2X0J5O+1de
XFmQ7ItcoDMqK6q4Tx2bg0Mj3W/MSKnpgh0TyzHQhKpsJxczIDNDcwG4D/T1Ea7j
VNruBfm3l55awmeKxyypnNIawUrEPEqaln7gYWBbhDll8gBqnGvLdLz9qNWtE62A
QBr6iyAjLXbanO5cIh0UmfzPk8TcqW7bqga3Kr88ZvzSqAREZHKTBF5lD+Q3jVQj
1r5Vsll2Xm9FICJvCOZaa19jDWTXbV3Hwb0qcNGZ3cop74VbJ+5qiv2Yy1CnWDT8
+EdlFvMmgYHG+XKPtlTtvFjAey0v+3YJ5SJOVuhN4qqHbG5WeM3jS8nfzY1zy16N
FnK+5sjFAJXaEgV/KuH6oqNH4X4y0P1OKwT4K9CUBma/RD7SqcAUols/NkzC3cAZ
1joBkblO8nHo0j2IkJmmzzoSfcGfFPHMMphvtLj1SI0zQ4//+hOH3QAS7MbHb8HT
qTPjCB2OP9vC0cPE9R8JxGpjk8+U3BP2UNNv0LfcaJxDS2XmzUXmsVCpCvYvw25g
R3EI0iSt/vtOgKWW7sOYRxkVNz12ptSzB883jN5wSxxO2h46BMP53jH0jtOPI2A3
bOY2kmIr+jzUm0d5WMJ2yGu/7r5fFiyvS4wRDZMAoe2WkEI5Gxq0WeWLcE2Ggj0y
PqOdYcp7fP0yHxY0RPO7k0R/j2+at24nH7PT76jUSMeNYEaFk5/D+C0xR3Se9AH3
xpO1v9Xg4sSdae3cnjqVFUfWUo6gszeiJZE3j3ijSUWiF1fPu7ae1UgrgvCyALD2
Fhcoj6RlVEBa+ZdiySu4bvGFqVZ9+RIxd0EN8b0btoboapNoU77R+A3OA5uJCraa
7YJsutJq6iYBT61r1Ybb3Z74kXvsrpIN9XM5p/e4P+fOccfnZl6AZos8IremUuYB
L2n4+aWwHunVPJfxqZE/Y06C2Ro5CXOly9IU6Ny41aBo4xnU8O+L1WNRG7Tk+yf6
hW9fOVcS2lbL6WurgvoKfA4Bd+j/MdGRRxScybJ5NwSULhSVDd8urAIgOJ8Xu+g/
AaiVfJzEkhJDAE57Qf4HNpVUV078673/+sGGNQ+fJnnu9X55v9zlxfgA88zpDjKz
TMceUYXJUmFRdEOg9tNUuVdk+WhMCQWLTUehJbAIq/tqO4ebfbdizhbZUgCc4YI/
V0Y7H0Djg1FXeL+zBhkj6uItx+V6zZEZDrZBpo/C91rtPstzgBOY/GnUfVfOzp9s
1EICoT2DCKlfjDkm+ycjg7mVGs8i+LKPEmhhmw5GzzKB3a3PRMn0Dy5+8Y843Y2a
wEL+iFTua0kNKt93v3iUOH3sGuYPnJe3sMYMp9dGkr3jion97gTiKCT7iHYWsNNt
8j+rq9Ld+t/ZAzFBDBlknw4VPx6aD2W4c4rBHZHkh9gZzZs7z+ugnEPxQiS6y929
J6wD9yhG9JeFmtLVrXoH4tC/vwx3RRQy022hJ9haRliVNIHqiLUFhK2NWB1YPwXO
Bbg/Unezu6sGBxIQ4s3tXqNR3mm9QSnN3TyjJZ2zSR7zljIqY/dS8vS1xmR9MAmO
PGp/ERPPFeaH1d9maSDWSTFX0Sy4xlBTfmzerANexbtg/2mnDkFR4ZqrLzb26caB
dMDYDdGFvyTH6xGbFUeNEP9jq0OrOJEv5dedL2EM4Tzdf+9UJiyz3xkaSoZ4p+UQ
R/29wDqEqXaFnXw5iKDJtGO/QUuM/a5/gWsVNRJ3elJzQMQHKqow3sni8XzFS3iD
RmLGehyVev17BOpXpXMMC8R9ktrf06LacBiUyARxgP0y+17Wg12zxVCx9i6/l+YX
ybHfshKK1G8aG3jFAxrsloTQzj8T7j0e09i9SoVFZlIUoc8ZfKU9fQKAQnX9YwW4
zbsnj/hK59W1AWpDsEdFXwIdRp3F9N/1ue6NCgTPj5etRBhLIDreAvdDOPWMJGdK
gSKLK+XFalA4H3mGY4o9DdIlXSjcYuGNfbB216qlutViNye9+3e7hZTMSgxGGCiM
exaOYgcP8C9BETnCKpXOlYYkco0A6YfXAE160LyDV9XycfZRt9DacygAY4leV66+
F20KeQSy1E8/mQARMfsh0rvctqAptx/L3ct42gnmkte4g4rUD16I+HVQt2EQQJVT
FC7bFn6S95DdqcczojYXeWIx4+XWb+2LEnay+Orm++IUreLQtcU4whN4NOhT70Ir
r2Yf6lqx7RF/ARma1l8LbqezRa8cbNIsrvv5Gbe6S042nqe92Neocu/263toSccL
AXVm8jGaW21FgaXO4dwFVnwX640V3amaoCjsf9n9UPkPA1SOkD0TXiAEwGCzvLK5
nXZY7801rZq5VYrSjTWc+dLhqP1Sq5rHi3K5PC5fdR7U6LvOD4Thy+8T0o0ba96i
6D9jEgiLLsVAaMa+mWOnuooTH7nvr0SSHr8IsQRGnbUo1ryGTKGO0Nj+eBTRWXqU
QVy7j6LEc/QwwK9gB9iiGHGife2HGoUNxof8Jhhc2EQ0jBgQx1dqosovdGMdp1s1
r/NjnLjxR9WgrKkv9Uc0LU7+BuTguk7u29bygbmjEtmFTSk8PUJhB4cQt+30KENH
N1+2LrD9M9fHY+4SytFos2JGYt/D4jwJg6wW2x3l++JE/gfzXFAW8rv/bokzvoZM
DUuypmJMX0lz8SsicXfq8xPhCczyBslwO3vr0ZuxMWSyZtt8/CA1COEMhngqxIwq
LjLHAVxuA2kLRK+RCiPtnRxAp1d/jO9sH30+Bd0AGT5p2ChmtXno3sRZDe0UI8jo
R0CyRZWghkusRVuopSMVSW5DrfYyYjU5+QuA9yIjboSiM0JxlzyK6LvhqeksLyn2
C1er7dJzhmHGHMd4CCpmU5Tpt9QfubtlFqsxIGlbxC8VbHTvKzbvfRV0sfq5+37s
mdFSCrX4bA/dEAB7MN2PlHdwLZrj4g6gw/jxjHOnze399tlBZiM9Pi+vl5euQL30
1R3RH+UTERhTgOBJvsdhrrHBx+djkIlJtnbGUCsTvTYMgTDClbOg5wD0HcSqXB4i
6btxwLwMg/m6BPatLOeUp1MYTaTPR5PiAPwV4wqjB/25Taz86gqx6HYBa9SU/0xB
ww4b2Hx871npbLnYrm2H5yoo+i1YSFroUqSqG8en33xLPVA3iOr4TFat5A7htuko
4GFgGaVD0Yp8wEVpwJAaUF3/o+//zzzVlLmrNJEVgMuvY8f9whpHl5tH+m1Lddcc
xxqRY+6oK5bcEutgVOG3d5bGDAKfeggNxdqphwxky33b6UGrVGgSnrYPh60FHepD
8an71oQb9QLUxtwjkKsW0v6ZpgsXfpoYsplbJIqojwh4eNKIuLEhKMUxVGk0jren
TfHmJIp9KJPluoOYnPdeb8NU2cWajgPFf1vJsHdd+tLi5o4tsbLUxc6JT8WLIZV+
VQUz5oSca0ukN4dasf4QaBmAUspyTdYiMcbIlPDReGgs2Mo7ZaPXXB/hU9B0K3Cy
s4C6QlFYcBrk7EmyqopX/VjduBzTGtJytZX9syj8eFR4VgrU5WIh9w18YB+Ssmv7
sCCsQDXDBBRj0wEmq7F79S8nIbNQtqwpwZE9+080MEd8Im8iXB6V8+4PHpGLn3HX
yerYSMW+5SorPgvL/Jx2N1b5glQi2ZFgIe0y+X/E2bmC2lM7tXkm47M3aWpM8aPC
r9JNx/mWfYLSI3ZBI2Xt4mPxGyrgHuKS6qQFQp3LW8auMXZceJ0dgix9g+sxKhtZ
0SCU5xlXpvuV9DZVAiZB0a1ZpJPl15Amio1o7toRSqDE4Nkizimoc8gtYumQMfWJ
WGheH5oh7u47P8D1LG3qlomEFPIZbJZP5hDABGAEwqt3H7eqmO1vtrvZ9tdosKB3
sM4ugimBkS7ggOFsC5KhOgmrgcuySKARLiy92IKYOG5VsK/IVF1kauHaCD5i0mYb
8GKr3rvVxQhdLsZLXt+qX/gIxT1v99XY67weo31SzXmhyQ6elzD3xF1p00ComNH9
w2AVJtH1FB0ZCHfvIfkW5sHXY51PO+853qsnFidAk6Vd9B0Zuibn2xi9z0S8t+44
PyJEXQ5TuUfM7JvXMaxSLmPl3Jg423wZJxLRmccH6Xw0DuM+oJX3OY86qALu+SV4
AvgI+DhNZEroVSD2nXpviMKmmJ+CjhyT561fchiVotQLmX75F4rGxWpuIEcrCohc
n8VDNL6HGjXC6lIAA65jeG/pU+5Btq19PFWDulDG8GUF3EOwudo9W3FHYEGPT1Ko
SG6cJZPbUCTNkzeksEj3uIdINtsd/S/flTmBIBwEtS6yiYr9jbLkei+eL2qGpzpv
TNwkXnk0qk68GnECbgnqmNj1w9wRFU4T6oXUlFGO8r7Iez2hpKUl1b4TX7fc1dDs
Aw+2M9E2OXH3yS99GiZSP5/wkj/3m3hXditmr8XrrS3orF5OCPjerxec0U0y6uQh
nxV7O6vgVTUjxJBR0zrVeKf4qcpVwSefEDgLG9dxTBEf15snkG3Z05sA/prYBtkW
/JRHihaGwm30da2qDltPxIPgochLu1FjIBkyBL7qzEBXenWr+FDBEJsGHp7/NzRn
QQ9h9UIQQcHi9Y7Kok5fEaXcGKUjVnY6gmBmxF39Dk6FPhoRsPKIwSUjUmKiEen5
7xvIZabjQGUc5SwPX7vauzGXTWHuCPjdjNTMLgJEDYzzuR8vzvDPfsomvDT/mqTz
B+/q457PlHsgDQ8cODIxcvkaKQayTCDW7xZDtMCKX8l9kDdKa2qbIECcWg4xM2aY
iBmcXQC+DiP7bwwqo+0PVxzgni5zeMDt+Tv2+8glu7eGvRIDqIGJGNE6yQlt8Hct
zM4wop5l6dHe+b+1CVHU55aCxbcVdNLKnylWZiO8mYrQ4m1d8UmW7B0v/vrcLyWT
bZgO3RbC2mfY/pGOB10PiE9avxLHlOZK0V5GrxsbjAzeER5mLzn6RbGNd+qikzEM
LmhVAPg7Rc6Q74Ftb7IMH8vf6Lja6PpPmdOMPyotUMZINNgY0hkgT490OzzpYzIM
Hsd39HMyq4bNqEw+81Tsh0TQAMeLDMd0zg6jx2fSu7PQWA/al/h53oSTb2b+WjQg
Fu6cUPfDyOKVfShcASPWTcyLHhMvGWyBhvmqNG+n1HVrcsHjcjFNFdrQZuap03UY
KcG+AkQnDAPXsiGe6229GLchvvnGyhT6fVPWa20c0gm/b6rAEhpUXHsFAD29PApu
/0g/7pJQMGQju9F0s/PZIaAUP4IWI8u15bcI2Y+VlgCQraqnkINT2MzB2h2ajBju
0zXihLRyJW+Voie6UF5/UJJAwjQurJ5UG9ulKjtoc25mn1qpPazaWIDnd2L5Kfhi
bon5jTtJWmLcJTNpJiOFfgtY3+H/3KIiGsv525zMvvKSqwLgsjwaEjd65oSpD6Am
xi3GsBZ9CIkOpqjQQeLPanGlQ7L0zE8h/SaJecf5O6P4Z6epCyj/CZSygQyUK16d
kXWxFLFueMR8qQvMJ1rEFNITs5hUBdmhYJ3Nj44shVyWaLvq+f/gtSXF/AVYxCAQ
ugmKsoJczmM2uFtxLzlWso06UmaKdC/l0y28VTppyF2j3X1WSEFEmz3R421yec02
kfT4q0qiooXUJDkErBkcO/3TJ/Tq2nAg3abow4BOd2YMyqOV4TmTDYmveuZ+MF4i
PZ2KlC4hS55H9hA/vE/edz8O3nqTNnA312iP1p4LbfOTCWSixsyVFNriWB8tf8FA
uVJ410kG29qB6nPWNECzoMPXXCxMwBx9V7rdaU5H+Jrk7ABVNZ/ySwyyOac0mv8V
ho8r4W6iC1UXK1Ay0gcJBRf7im6A6fbPYz5rZ5EDFFZNIducv7Ej/CWl6EzUQuZ5
3oQdOUlBfd5ZYxabH50EC6cdSEP1rDj+3wF6HhKW4MChzA1dM3WxQq5NQdAfS+x0
6BHRXWIXjFpuERvv7jUSMhIsMD4rYs5/fH2XF5jtFB7fh6UNJtMZrH+kAZFeIDDh
cAlJtQkj+QLjfJ8rNAZtrHe3X0t9xy2CbhopT73e6HYDY/h8+p984fVELEBr8qHO
I11mn+JVMCoNxyoU65TRvRHjmD7FlHHEXA1EcC7DZi8zHKQv1Lz4Qu64D17pnE6V
JAQ0lUIoeJ8+5wRqT227P4qTZBGZ0/F0W7tvFugKYTiwBYOvTIqwPSi13rnfgvKO
k7l2+++uk15JxbPIHt0WaAaIusShHiZMFDgvRcqQOcGVeRI2FDDMsVYF04RJdWdx
11XRhpAe0mNGr/EPpXW1nE06gatCnW9VZqgbweGsKoj4GGRHkmW/NBUELkjb704x
1WGF9GBdovebvic7bgTJbOTuhqQdw+CdEqOnFUr8AYiIT6N1A8DnS73IDAQsRwvq
vuAqRQNumVL4cC9BvxSRcSQzffph8HYbhPBZLmB7SvDjEjtc5xuv5mCZI20kbUyQ
X2yMhQAder9mLCjeseSg/Qt/XjxlUGkxve5JSDBzj99781iV4tNCqTEG9/AFq9e7
t6VGcSYdMi3XCO+c3b0YnVcmLyAPmCcg+QjM2GYm6GX2aIM3xpaP9vV6jwOHsBtR
uyef0jDg286iN4Hl6hUdZVIGXwRUfGwn2kttZhkyrRv7Uc/S7/t8BqiZdMpSuOiv
tduA1bu2ixiyQ1Mzv4h/S1j+WSJUu9ywoPXJjuqAsdYvNwmB8g1nx79CpSuhhUjb
Pnw3EjKQqEl0e/cE5oo+zk3zGid5yA5hEbAOkodCp02sdCH1nyphT1wuyW7x7E0d
buQND4bqMbbc/l9LucvjSMljryc7DSifxpuUqCjFDW6RRDx5MFJNPTHHZsqjk9SG
s2pNsnem53Di3fa3Q765aLkPhWwQPRDm6StQOFkoVPdaRTmWkMQz3cuiBQWAdcgU
4aVybKERQ/BH7r8/acpkJRBRC3fWXVsoPSA8+0kgIX5yamn5F4Nl1xijc2frK3Jr
Z8ZxfRpzqcTM5b+roqD1YIowh0t6D/6lRfYQmNGTMk86oWfnL9r0xOn+A2lWyhlO
1x0AziZwnT/gWJGwT7+lQBWTuqU1nwR6iPDZvVmqEXs1oT8zsaarPeVrBLrjAXh8
tDJeZUtUnTOytSN+AeiifgNr0mABNPTTOCvoKjaC4cA6V8NXUdN8aWfTSuNaAHAB
38wGnbtu2qkVY1eJspvUCvLMht5yO5XVtbCGxFGwyg9UXQ7mngH8Ns37rU/LxHHX
eS9rXEJ7aaqkQLrrxVYeiF6SYQKPTSqkMotXs3FJnhxYRQQ8Ax+g2DSQclsk5acJ
m/zwHvv+ljuSAJanEAhkAVHG/gCnQ90ANPxYHW/xq5wp/B5RHgX4/7QGkKqnOjAO
MYeL5aPghEWBoBnJ7ZaGNTGkT6pwNlVD1S2DRy1TEULyvxEjmM6C9u12eEcO35Io
BSS9nRXg7wshV/2s+1yqGsmi3anC74t0POQx/0FaslXHyZSi23UXlYA2W0lGPTXu
T+tB1L6KgDYkp327kH/ZagfMShVIdLQB271NI2X7+TQdiHSp+zJW8SsvCYcq8hFF
1r4JvTCRSrmJv3DIi1xLRXTx4Y7LgLb5/In46Zy1VwWTic/N2M4CC/z2rNEQkJZR
xlW+u9OfZQLCaXvHFCG9TX8TlptpiRg3FnbqmDY7oWGWUngKPsDKoei3s0p2ZTfW
lBhQU+6G51h3vNuPwOxUfAaZ+3HRRU6MuXrFyHRBz1++Anj+UyHL75ZH3WguXPO+
B7+zV16bkqFfTGxZTjCdYiS1DyhFFBP7yjahLDiB51fpxoLB5DwrYcAkQq8p1mlq
M0hx4KYsjrb56mppZKBfFdv6KYs+LxP1Gy0JfNe25+1CQgvo3JkowZKKzjG76S7J
fXnP/CGQiDLHvrt2196ALgMi4U4JCfktbP+a9eQBccJpehM7tB1hgtP9pmTi4qlx
/coFcuYML4pjNdbe0sFje14R98zzE2Y/JFTtRcAepmdX6R7Uj+aOk8/H9BGhtsE2
VZN2EidNc6uTjPVt4SZAMNmFJ0Icyq8xQpe/R+JM+r09HR5Zzu64nUTM8gyU4Q/4
sDP8KDT1/OdJoYYR4KHKUig9BI588nRV+41Q7OtptDX1d+03rKRpfW+6eBmWTyBX
8MmRflLIl7ZEAHTaMJuWLFNLZwdaQLt7b/SU5maFHE9grmQTL7KObGL4iwK0WKrN
YoUXf1y4DyzmjJvl+ELl1Pm9Zr3947T6aCSmjyd5R11pmTp5gI3TSmt7lioqI20F
hn4JOE3jCfVXj13egbmiNCj06qg7eWtxy2pMIvnFTtWrXX4Fv9qMnJIEihX2yJFy
EFXPi2IX17wkFrmmRX0BBxQ+9YpQiATgDO4BT5yoCktkufLaPKyhUhlqNs3CJjYa
2YYURyGFZDNJ9UC2Jf3XSn/5owfHQigzs7ZvrH33gznhY4maIbV3YgtneBnW+kf2
Hl6oaIMm2U2zuEgPE4P9Ypqes0HZlBFAShBvZmySfYFp31B4Gjs8+7pjMvbJWh17
E++CbXDWmpDRQcO1Be6NVWFKFmffXViVYHYlnDiHAU/v57Heq8R++oYCLDSboNBL
AD5JSHyGRbLcLy97R0HWvhNaYvX7ps4rUBbZAp/DB/AI6Md71fyYt0tAFb6pnqxM
OV2hfbBWSuZ+13yoVuf6GaX+z0h5Y3NE5mt7uzw8f41uY81/QDsyLPTyVdr9SL57
W+p/DPhYjtTVtkioNz9yVTq1hF7/Ig/SjM7Ebgbh1laK6DZweLZDeG3rm9Z3NC8t
9lP8a3tzPUMcPKDDUYKv+AW6Ah22lfl3uCiHQ3xmVDBiNHH5iU1N/R/Oqm/DW6F3
6MSqCghEOPYZiJft00xmN+TKoOAJWZGHd/ZUBq7rK86Dc0j89e/jD9qG4WLJAOV/
92+U3T2J9GF50Gf33kjDRRo8HBjs77kKONC4EYKgWrYpDJdxwqgdPR274/57xq7/
vfLzd8wyNR2DHsyxyiDYjQpXBjcDY41pqDjrHEKmU30/OLg1E/v5geZJ6RyJVoWi
cFlVKYn6tO3lumhs/GHikBi1BY5dY2iK3GNmkV6AkBYBewkSkf0hpgiljIb9wnCX
smZBuAXcG9fVKfQ9EWLi596/PT5ypKkQnKhoIPZDfVt3ZQhpu5IbhPQyOSiNTBOu
fzuUqRb31ycO5y/uDTLVl4msK0hyQf3p8ZEcDqoXkTCIfPawRRVzC3gD3Agdsd1B
WQcQrQ4seA3H65PH+9Gax5GeVukG7YX1N5cXF0GxhjNmfJ5DOWJWNKbu3WDCRfar
gs3xH++LdQfkmvQ+xZAzqrLRzAEf71qkQSXpHYukyGmueQoBQC4eU00J69GW+8eP
KqoEIyvwfWvj+aaygB2ROXw1/1NLEJC68tjISIb292A7kMMrTHTopv5F353T85zs
JHi/kP1SzZ68/QoyEwDKBb1YIi0Eqsrcy6DD/WCVkP/h3cFdGvQstfLFLqEz3lqC
BvYySdpuha7j7Rq1IA7WQvcq36TZ4Bu4bKqVh3P2O2y+qhNSWNe0jo3ZfkFFXBGG
TEP44xguGp49pi2vNW66znlUjD93n2+pvBQtXkofWjDvAW4SfD8qP27iwncvEMMZ
i+NqmThcbGp3oT4//tGlxuRV4R7zWmq9+7Uv2ALopWQmDrILCrS3hADUAhTHbK12
bw0EeMF+NfAiKwtCh3CINXRA5n4JSJlHfAl8whoxhwTyct1+ne4I54FfXuk0/Q9V
7/9YXR9mq+Oc84LzOjpI3sn/9bT4ybumLePeO/yuu76W/CRCBT7HMjGQZCmmRUXG
OnVFPpwJ8hg8noSPcntKpjpW4vAOr9FKfBxHuqZcNXFDuZ+YuF+WJLjdQPtDP1gB
pnZ5PTqX7rPvKbuimUAkgZQ6+usxFfNXduP4rkn7laYniky2+kRRHYGDa73L9f4h
mQ4kbpFBa0tF31Z1iRtOgXEsWSw7nAda02pTrH2YlyXdPYlsUDa4TjMASi+/decl
6AYtzrFSaj3Snzy34SDGGICtBSVxtQAr+R79WGakXIDvhRx1we+/A37JBB4GTbqz
Y0nla/jocWz7hArjl2JKp+CLGZ95XfS12a0QTI3tWi3srYDjenaqN2JHcTV3hb6v
kljW0yVzREo497q5tuxt+JNg8dkDFSjJkUIXjVaDyneufn/lvej9cP6gYnqUgXTk
KG7FkS1zUG4ugjZI8v2ygo0XgpgLQZkdu44VfghuvJbqeM3PRTElaxB7Nvjk9tPy
agtw6KXy5e0dTN+UCG+iQnmxgN983e7FlxlIbntg3XpECaJmblgpjhaZYTx3C+4v
Bxdxnl+eakY2EfTjxWiugJPRZjuiDYx3r+JXGrp4vlMYJAuFAgDgWR09YkfXX3wY
kL54rV0UIqQK8BbAx8lFnGtGmJWFTCTV1F6w6kpzXaKGgQRMJ37iGP8ojf+mTvuk
aMQGEKPnQP38T9VnHwhYfJZ+mhCDvbIv2yf6Ej4RYJUMGsW4ActXQvQccpN5u5Yv
K4fKFcamCQ3Pnqp6Np7+t+LqngUNBDZf7k+WJvYI74Ulw21QYJWmJBu+6PgCbTCU
QLm0KlYh0Eo6k8Lb4fyfuMVMqxEOcS2J9ozsEH6E/XoWrw+6QbeZ5BhL0CqzyHZg
27FR2lB2H2qHJEtIfPFWQZnaL5LUXH8K7IuMNQccVgiGC9mFaHHVHtUgQdmlCLmx
jUTBZiJkS/DBGPUD0HTc7XnWHbv6JDPUWhrrzC/DLDC4yze6VfAMmoLj8MmTbLNT
tdipH5o2ymAN579TPsvcz+lNY/dVHy6S2+So3ppDnz052E7/xYt8sloiZmGWxTwp
8wJCubDrSXfE5A3blQDOG4X8/Jsf7z2P5CAGdLIoCpCEasXybGwKwDFs5SAKlTYs
iMZmQjuSQNqypfFWkBNasMbyTQUKmW4d00hmrG0o+LKYE9nri4td+apbpADxO+MA
0lqmVjxpWZ+P7G1yGY8LzlM09168MUwrxp1zv5agnw5twnBBMc2vTYOLr+gcF5bV
kGV2+zwiQ3p/K9zO2AsjBgVhmdNS29rNJWNSo2NgsCtk0lenqz1ns04glFPFPe0Z
Y1hf5M3AfVKV9slsFOPT0XsoCL15SjxmnXUa0d22ZEPGIcZOQ7XFxX/kX4YC2Cg+
0MvsQc4wMhvkD+6TRQEePMjZ18OJIbsG+wNeY6vMYoxbBwlnhgd/9JhQ57yEAv30
A+l3WG7U7v2oJMbjjCzHLxqYD8xAZLFKksvbB7t5NUF/WboTCA2Cz3wkcNuVSRAh
gUYGfcTlnmXI1dd1Bpdb6SO4yj7yT7CSGA6MlAw35C2BjWE5P/Js3SAPT1A3omBq
HdMevOLolmPub7xk43QAmmtBeJGocLLXZ0ARp+/kQtQoUUgKHRQxcMjsCvBi6kZi
QGgIW6V2TqX03yr2fKNRNegKGBFOMZIerpyrO56cUydR9QBu21WCCeh4eBRqeatP
HC+KGv7wYea24XY2z0x9WWCYy4W8c17iRUE6WXqFn6a3FaB/o/9tcInfE/lwWMo/
K41qe0eUonBZjcjy+YzGbZA8SE7zB8aI2bWJcNX8GjctmWvlRHfkfj6zd5IxLwYu
/6luSGOOCCUu8OSQp05GkU0HQCwjj8qHRdN0lsvwWpP3Z5CATerPobwAtgcrf+IL
HKKQcOf8kIlvkpNAggrtVQWLBgrZaWXxiRFIbcBzarp+6oatQYpw28g2DRF/S5PV
a4gDGsboS3UlKgtshbVseFbWcgL9gG/1hKlve15fhzZbAUVA9Blo/7GryLSJCHGF
YigoLjxL1uAS6853kIAeEikEKd/Dx9d7Zi4gt5/C6ZKHc4gEGXGGtfWhKMnVYe7E
nzGicrZCZdBLqh7IoUl+NnOl89nttssKQnhiOoPi4WCh6gNxOkHLInfBkFXl31D8
czb/EBGGHuDufZoxdCsk1OgU3oMz3vaiErWgy69yJ6e332IzQSE1i44NEdy68puZ
ArzwPKaa8CQbwRfxFLreWaQBUnlel4l3fsX27vwmrFYHi/opyGHlyLTY1qsHLVbz
4hOnQp2OBrSMU7zM6QOheSd/807k6BABAgDbPh0/PThExcdLGPIjUmQcoz8MYggk
OsbTbKUnye/WG07PfR+qCZ2G5q8NFsgwLc6iWee9osoaCgVbyYRIaExDM7YQiGjl
2kPg4lk5tXBFZRyIPvk8yp097yX8jBDz6RtZKlOZnpW1CN0NVrAem7uiAsCfgaO4
zPa8AOoQSWG94CYSvLwFxx5k6Y7uIUr+CrAiA9Ay0pmtyb3eQwAsItWa6QUXfsSZ
tntcGt530My1bauLiPq0gnaJDUz22oow5ketN9ILIp3Hw8px2TaYSIN52Fc4/qme
sXgZNlLdquBpQxY4EB5skylz7PFeGvuohr/QnTXHzs+cSDuOzXVJcgdxWzzoXGO/
kb4rYVGXp2BxqefHv9T1n6ugUCMolfwRrrX6USykBF/73c3yMnIWuIQ23FzL6b0B
V1CaAFv0DnnYCyddsmUGp/v9T/QEoUd/VXCEJYaKPMqZB9DwpHEoc2n8mbnMqbLx
hd13ZGsMZL/uBEdg9U09Gh6ZD+xamlsL+hB6KlqPZtoNVzpos5QRdBYYOKFmHIs2
7kTdxhARyPZ2wIbKhLDsngZPBabYl1GeBbjxeGFFY0bER1wNW0Yb2ODp3FfBnUsI
L6w5R/zN8BLjUGj23iugcxGYZZzSBQC6kiX8vZY1jtepj4YyvQsm9DB26VRR+A0L
ugc9AkGeACz6rtuzNFOLzYdzhm94cy/5I+4Ymw6Uw5ffpQk2OEZe707/lfcCjRp/
YE/bnzAlIzCoKHaw/ldHU4gHe0Wwh2efxmZ8BUvspGsur3Gx2JIILxNA1eKZDjM1
JpwuOnIUkfraSrtzLIXjbmEsxlCEBRppiJN/b4soEjCWliuPe6lN1eUlXu+wBe2g
IOkXTtGkoREboRz0ca8HqRAv05xUDLMyJZZnYAi51TtD0pTxQ3gShhRNTAdJs4hk
o2RgjAglxS1goEciekQSD6W13p8JXy9nk75GErsYK9aq0wg3wK8meJ8gmaRlewly
yJisrVQZMYzNSYumh//0GV9Ck4ywFC8JcqqmkuD0DZtW+yCIVPPzPEy/K89A0yzT
oHgYkCVMfdc7ApQkcyx/iHbJ/VUiKIF1daDK5+VLi9I3kI7hLcrSZrxP/RqFFJ2S
HSeV8IIJ+J7t0f2KfZvdZRHwAucZHFQ+Y6leYFQh4uXyO0Z9drvyyBm0DN5K9Fhs
y8rHuluWyccgCRJ5ifsqvCiaNRQ8HRXvI7qHPYG9qan7LmAOyId+WtQV7qkxiPAc
Rn5zz6ts9TzuFkVpYS94X0G0AwsyhXiijwTc8sAWFMpP+IVIJZ1gEfdq6JNXhV0P
zEUPscWC9Pui3/hJ2tGNjczwyzYneWmetDJvMe5Sq5NH0qdfKflqcR1rGxlAFGbG
eMVY9RjT9kT+piqbFzq4qnQsi3dsXspqTGK+NZ6vYBeyJ4AHwSYKy+ryVjzYSxw5
OFVWfFqRzfsb3u8vXV5huMl++yo79VmeAyxjDZ3hYBLKHGsNwxDI+FUehggSojBj
aWBVnZBr4EqE7RE2fGhdFV4vyWYH4yfnSiZqhITlvf6WGSiaZWwxlnZfUkf9aKSQ
rp+nIAtmS8hVuro0Ufc4CWuEn/x03jcW+8MXVbMHch9pzRHw5uMkyC+t1pDzlfdq
9Su6z1f2cWpbV00lmr33iIfHpOvoijcN0EQ2REtTb4uzWoLInHjAE+W56olb5e3W
6gxlOTLXQAYgsmU5GoldPW6o6Wu7+S1neyycFNaAj8oDfVi5hFCmRQxAwjEN5uQc
8oSVyWEifF+eGJCGVnupXBxHfJ+D5rSIPDDeLl9co40kGX4XcZbb0YY5aRJ8rjBy
JkuOWdgY/f1KLH7Fbq9x+89fFCWPC/8IuqsptELEPn9NggkZiZ/C3Vbo55rnHSPD
8NO6AYhP9bKWJgqm2SGPV6+Eaar6Qx0ljwN6fQG29OOeSRvyFRbXNEjPACjzopvX
bn7DC9/aiq6iYTXsQechMOUvemFrHn+bVIIJDzh755n5c/eCh43m0hHW9Z33rkTh
8OJWOOzYLNrKTqyLDw6zZ+5NR9Y293JdXxujQzFMvS4fZz83iI+aMF3Su+e0XwUN
Uxfr4kRuGPlV2ExQDBPHZGY1yQvd+RSZEnuUh1e2tzLCYQoag4JkFFELoqelAXkb
IDVdae4xH93pmULJwVppYNHDCfH+1V74Ji9o23a7RuRZemoSvl4UKR52I3UuntlF
e1+miaI/64oRp+AfSp7OnsoFh9LMVDdNY7ks8Egurdh91XDoOo4sNgtCrUvQpVgh
pR4F+nV+Ll3ZwY4iHlviI7V8sAGEMx9Vjb8CFhpzVDD9wmFuuYPLxGAZqJozFSL8
paboFGleRYh2mZksRbfuPdXUPJ+yt6adqIRoO/M0VsWy0ZsGz9dawxJqR5YjmkXw
S2SvYdJIKQCZv43vEz25NUHqGNnnl+34fU5cUvKAL3bli1miFTv/uCorcJmEKFRn
9J8qcpatasH5VUmcItTwNNV6ZI87BlprYliEZT6UZy66sSzBzpE8nNbxdjH+dkqg
lbPsQ2Pxzkuq5Pv1p+bFP0/RPMmA2iMngwYySAG4ZZH6PNZj4X7AEkIIdN4SI6qB
Q9PWaLiFvOhNvuVCguADaejH6bSFRY0A+8jZucGk5yYTn6PSASpycRgchLzySO1R
VwX/scEqenMaZDOBQfcNLYXF2nM++3tQbhs6Hz1HoVRhw6YgCk0iva4fFuuEyta2
e0/5wkATXcRBBsWheRR1+5TyKycWouj9qBcMBbgPQJr/WdcZb1E7qdqZW5B7wive
lR4xbXY41+Hr32zUFnw5NM/ebZ+eGLZVE61DqWxPIwm/PIeTVk9upDbA8QAiAyRo
W1CHm1enUvnViZVH/iYmiUdME79xSKODxZwRamMoooYsYqkkkBWVZwvUL9COPttt
eLOhgN7tieqRPDOrs2+sns1JLCzn966U/+fWncIn4erAj1QyOma1kXFnWljHz0FT
TpHcwIxEq9YDveuYq7vo7RVZSPW4hUbVttH/jshH8P+eBXUf6LB3pJUCPqjHWubB
kGWW6E7sNPXlawqFk+jQLNE9aeGaoNKt/jICW7lXzAtREAMmPkUBED166JV20mD7
NHFMDGYCvmAebcCkF9HAHneGUJiLLR68U1EHQvx96G9vCQPYZrHbdqj2NteRvQlT
pa6uMsTQe+lAtJZowHeimBsoJ48fkHEDms4TTU1CFqnZEhvvQRNdEpZGQV+gHLzC
OGkGhQIO6Rw4K3SrdAc2WIj2/8BKuwsxn9kB8OesHTRdovI9JD4swccTsGh0S1GY
aHnLEXlUCQ9PkRnr0+qQ+BP87K+qxHjpIBlH9Z/XvBlBfvHrFxsGj+ZR1ycsHC6/
P7RwrBMsRj9em6RgHE4QzT/L4BtDHr2ZSNFT61rZIwv+bzBTzZKxlC7NQT/sCZwm
ejodOJzyV4rPR75O+YJ1ShlZymb0pnefLAiUFH8fXG2Xruril5Ho/Aqj9ycEisAa
7e/oMUlvebajp95+V9ojZmGlrbIjANPwZyrAYAYgh9GpuP7WxbnDJTDvBAUbc+s9
ZQ7CscQRxnK4Y01xs0I5ohWFlMi2WsDZWstv4R0Y+QxYIzrR9t/LZDw0xst5zx7y
OsPHVv8n7CCteQQVGaOsaKpZFLLMw44RiBv8qRhDcPt57KBcSLy7TlbTCCgwXA68
tddZ44CsL6Frvr6MBE+jJakbaY0wztyfbWEnqy47E8itjQT0p1Vn3S7QUkUvPUnM
kxrYsNVaHa/OjdYhBxOZVerMaWD5dgSFJvbm9NfqdHezMJwHalSoezs8lOP3DnS7
KBPl7npTRtk07FwCRQK7F9C8BWc1e/+SrQZeDBsQD7qSZyawmitW5ckC68FNVqMr
Bor0PpzVP7hKXdMlYD+2Q/hxvaJlIRoDDzlGy0W+SMf8nDh1GPudQiAUxK0LeYKF
5vWT1wEI4zncDBYN4YR1qsz8QKtorjh6cP9EytL1Nk1faEW6xaTVeV+uuFRAS8n3
P9dHMUUXFyFXu06yVrhTffvH6Kn6pHO6mmyJrsaPcrUwyPC/VXDPfg0vaugr/uK6
UDgxa7r2b+fT/ON5JPnO/PSywvepI5uzlo6H4qABME2vPy1YTxvq/s0UcaR8J5zl
vJ3zRaqW9mLnofrTKZ8Gv9lP/J/lDqw+/OmNYMeCBy+vAAGsRNYleSZumjHag+Aj
wqI4BtVfZhWaQsUaUGrTn9IsczkVexmpLCMrFWIQrkwxugD+yKKtOJSS5KWmuQjY
FrnbMxJCXNtMSZuiejp5XU2WTL0zAIvpfwfgUPildAJoh8igsrEoqJoZyL8j84D+
6PqiTCYWDk6CVAHDetLDEglLgGRv+3eeoKQ7+F/Z2zo//5TSZGxTJsA/m2WPUqHG
05NtMhRh5vRnwzGlK5TuLJUh2oGNGPZloZnkf+Hehcssf1/HvjsCR1SzsdEArIPu
BoVHElEGgH1MUfs1wV8+TO1js8atcpdqjBCDYpi3J2av2FbnKpMeMwnzaVLK9+BN
7kIJn4Hz47ODD0/Tm5uC8dJaSLckI6yGPFVUGHVEoko7uLkbDa83qTpkV03jWgxt
hvKs0Rn+hvG0loPG1vq8jM2gnG+jwvNahNNqbg7NQ68MHoDNhv1oXQmu2aSG/Gy7
lCrydK//QBUOFCPAC+765r68zmb93NZ1c5uX+LRP+023sdEvn93xmyR3PXLpAu1m
DR81Wgms7yrgXAUNfbt+pB23aDHFd2e3kOUH6aKLrHRR2rFhJbsPZ/7fKaH5h4+M
Kz163pt2YdiMZUikE0/MMH68hK9nkLWG9Z/9WOEQyIQzykw2pv8XVVX6UiZIQvIr
0AFcxQlOG1kqZo8vSMOxU8m5K+Lg77B7Sz5fmE+aQn9o0ZicAzXtooyysc9JRpRP
4ncnl7Uzier4jMY+ZJLU3noGX3TmNM8RXC6vr7Wtcr9omcgcI9BXZ5yuOb6q8UNa
RbzgFi7e/uCuRe9r/kaBQf7mkU1yAOXauGFCHF+2dWUdOFbp1tIM9Ywxzzh2d6Yj
F76gIkx73bOswTYxkqaDG/J7rRiMy72cbX41FBhrsQwR1a5ME5u9BNHLX7vkSprQ
CsJePHc5+hqr503WqB0dWO7pCphk90iDHXRQLqcbwmd24BnDwYwRNwa/z9/XA5AV
ppr1Yf64hkY3zSExeMk3Z0NFHyDOORlUabukOmt1DvPqUFklt28a80nmVS0T/Y5X
BWZytIrspGuWHm/d8kHxw9xT+d/y1IY+aauNsqdA9bKTLq+p6U9ByERHhS++YiqW
FovCuO+C8QRyA7eEqujj6X4x4AsrPvOvX6Ft9nKXbtKYwkduNbTroT3gaG5dS3vF
FbQ2BRZ03QHxwdmt6EpS6hzCCY99UmHXZsglBJ2PdIXWYdrCEEXeKKqEbi+R1uXO
Um/74YYEMS2x6f8+LZwQCjNy1ocPs61PRGUn+FIZPK5tpn2ddyGr+XvkNC+XwfQd
POUF7RcmJxekakJ10HbrxV8bqKaVJRBN6A2s0vR18gaYz1T1KugcDn8QdQq3+vM0
sbFVrBcKAH/J8oaRAGfZza+YRFLmRPAHhURw9IZSGUuJgYTfAoEYAXvwba5MkEie
83WbIbk/lIZGWX5K7fhXtpIEpuoRSkLDJxkwTZhC0+0i4OYjL823GNhqRndBAeS+
NIEdQ7dVennBTvuscT7TNGsT/1exMQgeAeJ//qaTRGmeTjZg47zrXcBCgXNQWe8m
MhTfDMJV/TVOAbiN3wzKk0sSlA50HfBmq3kG/YEGxviYLlYesinQS5izsTcCsqOw
9YPq7JMmJl8rVkRsOPo+2uJ6JF+9BfVhwA/Yro/8d8i8WOiwDy30DncP94+ATWrc
0y0ha1zQfuZZxG5uyB9FNwLTKbusdOKmJWsL6mwYYob+XZ9vfs84qHkrK1PprTHz
6ABT8497ztf7fEaJCZHMjEou0vBeXkrZThQpyzqf2NpV8AAqucHxpagvX1exJ4oM
fHRO/7cBIUNZR9uuxKQTvNk7fPav0qtCYOG0mdm3gVOg79SxpbWbO2/QZNaC9Ww7
Iv1TivJeK9M1a9zw2R+N8IiFVfIKnk8l/Nydk0yiG18DSFQQjVI0+WQRu/LBOmXN
bUqAM1l072W4LU0X8k9XtPbzlZwgpVeS7HIGQ60ccsmBJx/lhEwokToczOR7Ekyo
53v8tZnv2fax/AONBPw/Rg7OJAIQ84ADPu4qoX7TO1oXf8nRF84oxEaSfOKsgYyu
VFdmYfE7b1R+FzryEcumN+WZqwcXGHjGXymYxYOxgkJs3bnWTvY4aHVq6ShHsOC1
ChvEG8/WLD/wXGPkk4wxbIhDLp7AwEeoMf9iMrIDySNCZsmw2goGdF+TyRyxkYt6
CM+gYPyeYb4Y/I//kICzakz8fcKN19+oslN2qlCsjVYHJ2ciAv/7T7w/azj62U75
YcX/3BGHLxKy6rCKN8iNY+CxMRJCBKw8+fOpesL3srRRvEmny627146B05rOI5il
gyl3M8xTOZM4DkWefHrgg8mvMsHffN4ahYaEFIdpTyKQbjLYPMpvDUcliIuOXEbn
j2svE7dcyYi/c66PrX+UYFVzcaKfG+x4PzrsSr0Z/1vEXJHzJbNiQ8j+ZvlMmFfo
Yt75ZAHbs6VaY8M8Ymf5DgijgcKlp7D3Hu3iZOYwwdXC08m/F1IIQ3UOG8Ro11C4
XqYyIkFPuW0QGrw1gFIB2MZkLLT4VJEv9lTti4I5NQX2RSKWojcB7ijavAhz+jQy
bstvNbZZC91yOaJ0pWxNARU7UOtRKOXrc6Sh/Faek48sRf56A5UFId5EV+ODCuRT
kozZGsmQQ/vL1a9TLRy+ngWIPXGQVsj3aRL8VAPGET50zGqK4wGoYGnIBjWX0JZf
n9BV7ZHgseMaVwlssDZ2/+rOpVRCSqbQmpRe7t7z1wf29wZpN9pbPVFHpI+CA08R
SPrYIzGKzU/si14Vw2a482jdj0LGARL3lUGOaL7hRI77YNtD+qvoNGsoM+ane69x
EXYrhX8kDv+iuYN/wA5bFmW4gxCePht7JbAUVnn/wQNzJNculYUX+EBn7nHJWhqn
e9j+Ps9c11gt/DTsNcvaAw/xP/++lXBsoQGlvOZjSdW7kVR13eNaTBj7eFfyEhbY
yYsvdijOGoOVMlcE2Js0j7G22GTnoHpL6GmME91zR2iCVKIJNMHnaUUqxuxNSM78
OnSfwKt30ktNxQWoL/wAB2nvWjMkQZpkIGUHze0npvl+gL0SjdgyOaNAZqfW4Zno
4EfBd30ipRaOsQWRlJwoswSZQWJYmQgdi2oy3c7tLuz/nAMZUI8wka80kHqtmFQv
E8kXL38eSqmzkwR3ynWMTGq301s4Ztwuoytujqc9dBgXl6WPIStsqVtlMb2B8KmO
l7UAeX7Y7VFURV/HGF4i9DP4SPbW/S6kxp++GyPJyMDQTrUVlbI3h3CsqW2K8oD7
9WHHW+bP8ndvpAb6I+b+VtIDaItee/CnP/4AeQpkxiGuSvofxqZQwLCDp5zIR9Mw
9ugWpJG9VmP+WUQT2CC6dbjbEOaeOuhH9hB8Y1CTr4gbOwuKAHfnNjahuDnK3NxK
7JmzIZKcZa/62ghH8vdrT9Cc7iZY2558BebL9Q9FGj2JYKW0a0Azffm8ZgmF0sj4
xntSxPydp+mCdVVD6wnjt0D0jowOfLi1mlifhpo7PZLucOqkmQAIQvZv6A1/V5ZH
3NDZ2EMfjijYzSrQDdOnLDvkMD7eoxeOTkbqlHv18bUYLgdta12FcNXMiFQxfncR
7+WVMw2gnFDs5ynfL92wei7WiLZXs6dFn2nD7jpkWqbUgkcDh8b/AgdX8i2Xxpfn
YxqvWQfnCSeMGTmDK7OBdxfemNbe6WNP216gG4fNRNv7Y1R5TYHA1mPKWHRz2f3/
vuhOL1hLp2pNHDwclUJRzh7g84llGvq4wm/YCNVGqNJB2pFwNKWWGMLQd4Qv0Xs3
GouVIjWTvqisP+/k5sNuHdGW912kxcGneVU59XCMZjrycjuY/SWDZ3gWpmh/aAuL
j+LL5JkdTYKY1n6meBXttah8ncWyYYJezRznPEtMpeQVsCaImOoQ9HVxpHcERpep
cbXxTG6l6uCYkpxkwiex9RVcw6ulD1qdFBjJBu+jrmCd2G+dJlWiBd9xNQMHgHAR
FBegV1mEqYHwGNqK+mUVnWMjilZSCwmZ3HWk3gr646TDWe/nxRFIYjC+T0tlMjWZ
AwyeD8j2rDhW1jYT5VvgR3eFrvPmqH8QrlyzPC/1NcJ8iBtfxL4C9Hc2cIh8XxR4
gUXZiE4NXCLAx43xq1cT+JolWeJCo1PdJPo/hxN7ljBp5YwueMhf9euThcFXCqa8
B6KTsHm/eFaJYdVk/7YW3+BJz4pJa9RrjVffRJ88jcPwtZabpOyEif/1UJzfeG8t
haF5S6wrCDI18FQdnlu7QjBRXjppEKTi86LcG4Yt5w8eK0gu6PLDg9EsMELyihEo
552RGeefInXWT+Mk1y3argYvYmKiT0Tdka7rBE/UYaRBfTc9hlXYTKeYKq+fnTjv
K57pRVRUQgRl49qnfHuJU0JWuYp8fahNs4fu+8U1L0ahxXGCcgK9YyuqqcXhkyNy
DbiUl9UpPenZTLy9VlKHP2RDuKzzgCoIyekku7ciPTzJ8cSlfiLPh4fF1iv3HdT2
HyOjZG5tViQ5LkIMEqVm3HkjwYPHVSjTBOJSmHNhRMXe7D5nm6B6zI+uuJKjRfLH
pC5Jz/YC8+0jap4aJkm2qupP9dJvDK2MRVmNe0P5i7IHsY73ckT5xekZN179q8gd
5tS7cmRykNC2hBm6qdWZ9yl7IWxou7RMTR4KDVjFKibKw2puWsMn7Vl0WVTQ3DbR
iEM/XBBu5k/K/fxhfx2vUfOSpd78yf09wkRNY/yuBzo/wnWoWrvcD2g9+umsOpnp
2i+VSacqnn2RYcPQLu3bm1DQZIl1+1IWTwQzlVminQkxLOsHwDVOeOKdQxJhQFJc
De0h0hpUQ/NJ3k4sQWfTYK0SuZfwMTwH3GLkHQSnxth7HqK2OUQOs/LsDhBapFA3
x5DdzdQZzzzC4TJSMNKlJFv70ME/uI7HfsP4UUWrEW7mSVorz6JD0i4gAfZDYQML
GWsWg9R7bY+9hZ0JDchpUce9UQDpC9v1He8b++A8hKVgz1y+0LMciU8AooZLVlgE
S05aUzd4c+9Db4KH33OqWFM3Ml9jmsnDwv6DIwQnemxar6nN/8ozL/yc95oGPqF2
7Vt1+SA2t+jwe/XzjsCahuE9ALH0MCdVjaG8ajU/oOVkL0MHUX3+zgg3153d+ph8
aEByhpWJFTqeQmMFhxyUA8GuANQGC+S13pHs0kH7ufhbqpP+xICX85TrVbzNHd9v
FGf44ARpLqEndH+uU3AZztdR54B897CbCaiTfRDbduGc/ftBi/tIdXe1Dz77+MIc
NeUeFOgbuoxoPDNOZhfGGFF2lVoDRDWkrZCRDqEb6SosTB9LzZ039Wg+9+p/rntc
vLcuRr8hNu2+rliu180eAwAs6nQPcjL1mXD4/oIADYBZgnCPYxLf95SKWBnXU4Ux
3xNEdG0LI5Z6kq4DQwt8pRAyIofKzJzaUTKdMZQyoQHJJl426WofiuqVwNVKq4Gm
50OB0xw+/wkpVruBNTg0UZtrjJ6lE19ukKlSrak+hqWfpP2iDPffmkyw23CdOEXC
L9H5aVi7xTHG2mMnfkNvs7rTF14lJAlUB1msfzvwZGSQ8RJGRdn1MaPrMnBdEeO9
pDtsT5UO1wcPza0zY1r1Jkoq0gal8QKEmmbJuUKlwQpNs/au7CrLGFNxJhhEammM
fQLP1mTWnkWi5EAdD9H1ikWdiItWwRrmU0K1EPRyHZmBOQJBOl29/i+YmfWLL8Rn
JCYFI5iYcznZJQS3J5HyXTbUSLBv2hdeX4WEqhKSYZiCtZkZiXc9G8XRxY9qMmjS
kBMjnYqNJ4tX7+olTvBDtvph3+9Hun5NIOpCU7Ibr8lz8AOshRsOZcZPYaXkQdBX
oQDbUF4TtCZvgFqNkiOM+nqPzTv+kwgD/d4uvGH4guVwFmnN7Rf/ps9x9MLMTrkV
x76qpicF0khbXMd2rbkY1tG2oXmzuRB/yCkNOyJCqLdoH1te7wMi+AWL32ZVwpIr
1HWlqGb4yTWzfye2Ruy2aid0ucO6B0NGNh9+scgTF8WdRZtTi5P5ipX/hINxwMok
STt7rMkGXzCf9cHpm302axwYNEK4sAfPXDZfKDYHKMStYepsJwnapQI4xFY7m5bo
cTDrOvN+Z/2fbT8/uO2rUgvwyfKGTbIBxvDtJGpJYDuj8KRG+Dr7tmTE+rOEUlOI
mJPJLNYh3xAJDxrF6S+3/HTgnpM6tIBCiWVsm17mZHHGrxJmdZc+1hm9NKxfCDy6
ikfoXXX9EeKmEoNDLmBeurOTmtnQCvdriDMgT1H0ClD/+cZXqAbma8nqdDc5+0Js
I8PjwBDbl3SiccjaRjiIJe8o1ENtJmnt1G0oZ+AOdx837RhOfzfJoqiUGRBytqHv
IG1iwh3LylQGHcTiJBeVdGnWA7fchQA+eYHrPO4E5Ig/LNTsntilm5UBUJHkmm+f
4sjI4Hx+3Rduqu3M8b2Qqgal4VsLOX69FnzkKSROAb4Ii6CDIP3VtMm+T6HFWOMK
Bz9FhiOx/arGcf5EeFByoYTC28NjmimK3d6Kdu7MqVnhCK4ylNQoOTMwb4pfex88
QrsMLgsU+Rg96PV0B7/QvCHAN/CJ7n+uzw1qc4QRPp6dhlJvGstE5bpF71v5uYj8
Qp/hPGy3sU5ehaA6niHDtT7OZO488LtJifRcP4Q4BtcWyAd7lHaUmcKzEsn21TYh
RugTH4ZXs6X5wnoxaSDsmEDhladnNlke2mmYx+xtEK5fScujRI5VAAEKlq6BHDJi
nmy/rPAEHhVAN+YFI5TJWrbJeN5AVwzU1DfI2d1OKVp4A4OlECgrH1lQxeDycmd6
ntg7qt9a6drYAA5h3RnQY+nZKy8YkO/gn5yrrPffS81WVG/ZLsPCiGoNzLxUY11s
ZpaGeqB08bEY7mSfjjKloTa1ZwQ0lg/Lqrx3pp15IeMZmYJtzhVNZZbfIbiz/TfI
vFL+eYToOevk2ksseBEkZ8t3GpM9y7EEKrjtKrS1zG8owSlcyRuRN2H5GclT/75B
bC+lXe41rhQEgS6bjVqg4eaL1K3F0VUpT6oc/VtXY8RIG6TNiug8UdcXA076gS5G
5YlSl2zRmkvmjOEikBY/zh97HBK4c5lfuDddD2GiFRkm5IYJEHqtKFqJ8vT6jC+e
dGwiVBrfYR3kjOH45/39iZ5duuT/bVk9szqdAK9W0G0uR2VjxJ/kbYQZRAhYuwjT
g9dk5J13I1hvqh3PmmeRSjTUMxrfzyATXMYGRRWUwUUBo1S9OSth5/thD9BbBq4O
J5wnEiBRD0k8o9KSHB0nr7sBsonbbPfKGHuKXzQ/4+uKXwabBDwXDPqxnPIeIgzd
OaF3sRyEB5AMnqvfPLApIeK5d5TwvdKV6FoGTywtHNm304cYlCcF3ii00YHoJcA/
BaA75y7cL1eFXXo4UMCP7YgNWZ/8XSZ+arM+7QxTxfKMfT0DktEC0deWS3s2PuJ9
kfXdcdTnsmImSpc4zTLNHJ7MlptJfnIPq9cIjo76JQ6I4tifH6g5Q/1hngLgoGsJ
gP9U8E9qamQg73b51XncykaWIVz9C5kNECh5H3HwTv5TrEWn5yZ9oLkrlm54hL/R
awiYDclUKr6RncxJGUIhMmsf/QXn6sq5I2IWyf/SksYIbg+aIEutogjHNG5OjZwc
lSDnSre2e0Nfjr4+zqOhrONUKymerBXgIUlYciuDM/hT5ojXKAnBVwhAwAcpPYvR
owJniM56K6s0Yj1StrsDDjCUW50oZsZABq3SLHzQC2jGeuJAot+NhbZOeMDHh5sz
ybdVRIMFvF/ecdQI0fxKLqJToPNoVDIBXUs0MEyadpfi0u66m9lRqEHdyMfVbTNp
lIFPYbNY1OAx3XofL85RFGzl+KZ2ofd3T2I6wYZ3AFcMmuObjCf11GSUb3hQNeTj
GvO3ltSGIFWI+/DFX6UUk166vrkbUkeM3m2spCpHrUu/Z4CxMCKUyQFrV/RtC42j
+cMsNbWaTlnh1CUzrAdltFr4BO7WzJ19yxZPcd5SRyMlVVjqHWy0uRKuTqdmVUMO
AnbFwvAPSgo5hgXAhUFq6MdHUfYFE7uT1nDmyMkII/Wh1C/zkcaXm70Aztu2eiXD
+VZo2bqssf5xuj6PBsilXQwzUQg4Q9E6bRC5oVit4BcsMvpbeaTvFZU7PGgwL2kZ
KW2zR3930e/nz16LSdVEgIiLmbYD3tR+P9zQ3zyxmUITF+cS0GtFhgN72rytlbaN
JYw/qRNnQ+c+/8R7pCO2BUK+bL4+yGXNP7ep0MPji60mUBDTFuApLoaasWNjlHne
XlSOoVu7A/agCjnhG9TJJ0P5femm9Nwm9niEDdYO1b7MYqKVB07UgM34RwEkIL40
ftFgT31LWq4Uars/AYfILud4+u2+96SAXr+VXcuVMbrIdLAjr6obS0dI4VJq200D
qf2BTIF7gxdRBiulZxezvLYuSOyxE2q2M3rrPrYfn/sR5GA7bA2phTHsZJpRQYhp
bQTVMShsIEVAu6XySIRI3PpzuCdfnMKJwmJGXOhfvBvgUxEXRfvRuDRuJndQQ2D5
xmekE9uDe7FNvYO6rt2bcynnmwMgTYYAAV8jXPlX5VtBGMDr050k8PCeaIf+RIA9
87/eUH2bUjwlllsqizKsz1/xG+04A9/7mr3Nnood6iGHIbhHUMGmQRzakbY7wVIf
jSTs9o2pJSzBRRCwoZFlA3oOo0ci+tk9eKvKi5796DvLcVLCz9+nPyjnx37wsor5
w8QG7Fie/AsqUgsszhxoXgAe5HuibR6D6GwU42aLUClqWc96CIzjbD6QBw2JJVdS
CkkfQXgcFaFviCBLkNirw8IEf9N1dNVm5OYlUknB4IhuEUr/FQ2580/hDCTTMzlg
bPrd8Fnb4xpkZ4aMpCQ9oc8zaSxpTSFZ0xMZn01GT9R9YL9vsNMhuI8TmUo1h8bu
wr2H239R/MykFGEx1LDe+xi4FrnuvR+afx/+vxMxeyM78tU8a+jQuoRmbdfqltSC
QItbJJYWFIrZW69tfS5pHqHcFVP0Z1FfWKFEJO6f77EDhviGc6ETxa5ORl6nyd2y
caIEokgSGsPjvXoc7qdznZKsfSsnlD7yDhcRSN7BwKVtRBPz8xuZkuLV8WizZvh3
U8b/zddHia6bn991piUdGPMOET+xNKXf4DgN/itObEGOW0wa8BLJx+TESCJjsKoG
/lYYDis3HE3q68Pa3E6MdftLDU6j5/HFgPygDeUhOLo/OrdJqnJLNEw+0Gt0vqWV
DpG3sOcl7feG77C6sjMHdTChxp4DxhVHZFTjVMZdO9CsJ9i8YMi2L0/T86wj69li
agouiT8DC7bPzp/oHgJTJfbB6xZ73zoSuPEHg1kb0ibnkhMJgN7GMUXd7wnODs7H
1pGNA/wPLL9npu3RB1h1IGyHRspQYLkLXqfZ5Z9p8+YSw6HzgA0fQgsUg11fDBSc
jb82TeL2JMgd10+NgdWSHIyr/QpVGvN+gl3hdIfKd5cqWYKmQYE7cv91qu/r3ubz
/LGpzQJbb3FCwYMA623hqk1i7ctNQQgEsWMuOIKRusrFdE0NakScnMGy3btd4SXJ
Xg/j1XKgOW7LUGQUp1WPWb5+r55WQbeLwubjk8ySdOdFJSk6Wyi8xkH4prOLyQhv
7X3PeHQcm2hX8iSscG9E8bQVO5sBOJi6q4DvT41duiPrYBasHh1EDrLBtB+buL/G
zWdqDy292YA0ha8h16CNeBjCjeuWB/IVapFfTgfViR3Y3IEiqerHn94k3MFlUwdR
rvzF3r18Y9UD4GykigUvztwSuQDKuBPt/cHkjuVYhBt3J/H4sF7Xr4YFMM5zO58u
4+EPgYrHfSl7r5M78wk/bibSN3WS8FL+rfP0bPyIyoMPXxyemQ0QzwO40C4SaoLC
xAe+EBp3OrlsT3xVWFKlY9tFwNhn1VaHuloOj5qhdxaBAkqyCbMJHpBr5rnCitWL
89wWNPY5F8Mj4znqY3KL+mm/hiEvefSr6cpsvmpBmTGhWKDjxLGjWc7O+sYGUN94
KM8+a4WjcQh+l+7twJIQgAvWxgecPRpnLEuuViMGds7ihhvvm8L/2ZmSXt1ELVMf
71E0adgFwCj/trxdKCzNk9+1TCHYk4Pbp2ZUaYwGnfrllxNHmdbbfTGJGNZ7XCAM
LrEGxg+lFbkvIHjX/EvZqhyhGDtXAAwM4KYHoiU0X9DPHgVu98/p+3LuLi8elOb+
WUBuVNWMNQmr3RI+/Ix6Mp+AkLnUy8SDfsqqDITObnU9WwTs5uH5/gkFBZ+TqmnJ
Bz65Zjl25DRinNEVqQn8DsUwtWFdo7uQPWEMMR9k577b50Bs+R7Ub3WGAMaw6F/7
erXBdayP1XHh+2DsZmyJvPqDO//8iyf8gjDRF7qPVg/fh3I7OF4CkBw2dCccHAlC
hzXExEtWfyBTUP/uhcghRgZz6HmqHWx+JvNx+8jnagENHzJjs32CIRfmGpz4afML
TQccHaxNyz3drBQopp2VyWS1/CnaeSJN2+ZV1JBtCBtaWN7oGZGKLNyJBLDYmB3m
ZVqDNOMVzVe+sXRJUDCmuQP+A4hB9YmQnlzoa436M1mHvTdjuQqUZpTvP17gvw2c
l9m5qcBjRr7+dtqbZc++aw8E7Fp79IMnS/wZmCj3b3R717lt6HOC6Kfws747D1dn
X2aaQar4yUWzoJDT4NVw74PwaJ+EVA/gLgWSSJgsykykREsPV9FBZNdmekkzNdSo
POFmQBvYOyiNhc+46hS5+9JivzmqOSODtctQExy8g2qpBOxYaDe+lycL15lcpHeG
TnfAB5LV/dgPImtZkRUhNHKTjZU+rLxmLM/kK/WXDtouPLl+YAbbvp9WW47OgBph
Zt2D7GmfumVeCqFHFiQWwbYC4/fqfqsHqf4Usxb0datkhvfKTH3FlmRnHBnt7OW/
O4usQEqxpfzYj/L5dFesnPwulttKJDm0banbBGBEp2d2wgQuJajEqYDMSsvsGy6d
QRq2/7f25I9m8Z+r1SmgFzqh/hnRIV2VnjqGPjhCRW6x724KT3pWSy2B6f3AGtjq
CryDPZIsS7tFaPLOtOZgrJqNn15GceSUWjy/KtJ5mZ5rTMGt+/eRRM9zKGJ5ml7l
OeVAoCe24ED3fKP5B5phVs7qdyqo/OfwXjXUEXQdboTv8MvaQ8VnJCQ/nsgs+mee
dYASA86SPzclgeQ4mGBPqgLvMsvgtafDSr3UfZF/l5m47thXcob1FHUvsqDTE96J
lBniKZG2tU9anFqgE2m9lYkCa2Mwkmu3ea3npMRIr/FMYiA5iWr/l4lnHkq3JrXj
KKsp+FcWRO9oBPFqJS6IoyZZOLq0XvRFT0x8JeilIGizwwv06mYOhc5pUE1b1JAq
e7VDO9pihSkIgn/6V/gtWXMdkKB3T0f95ujBpYDs0V6pRQ50ptmxeq21gMxrd/WN
mAd7slyk87HWao9ffas9GUGwDmnapVrnV/tbIyD6/GJMdZ/BGEr+QQA0dryoCQbw
M5FACeKZX0rv8NsqBuUTLxVrHXmOZdl1ZMG035JEYsi5CGI9j5XWW0bdUtEhVnoC
ZMStNnTvDtrvmT8gBsrlNwDuW0kOc+edZtFz5XGZEyhhiC4BTXiZHoE+sTFVhdGc
577GGlPx4fkKtaAhviIE8VdtFD+27Sg0OvIn7xGVq3rfJkRdoNZjhANIUdjJUt9p
m9iEOf7GFbjbQO8FwHZN0wswJ+kcRuMskvfMtbbZocY372EmhoyZwzudyycZC9aK
Q2bc96IOVNyPaC4Aa5etIECxuAxjO+xxVrbrjG1/lMZRIZC6QfTsToqxM2oX5E1G
eoPH5CdaO0ckE+eW2L+ZJEsSow5Lh8z9VuFLtB/M+Wo9DPQofsP0hxhkbEpcP5lI
b4BjIq+9GvmEYD2HIaG2lFrLto+Puc+yVsUCUmVSmaS6AJvOoWmNMwev/1DJ5mWn
DZZ79UPYrWU+61kzBtCkdsaJ/uhR8GcYkW2gas6AHeG6OsSb29gw0z72lerEr3UB
cT9G0KkfgixYoRvsIByWzWFbZcHH9/xEXCkmNwxgNOEcTClhj8OFGVWm2frL/Sd3
0N2Gji1T8TErydESv8Kt5eqEOtuPjk3ktrW2bEDcTvefyrt9okFKroQHbCOM+3W8
ZF0+Cup66Sczd3J3Pa+tHYIEurjja4YJh6MZtmBb2kzXRc0nq2tSITWj/GR27eXA
FSux1EsVTTidp70VjByGDNUDGm/InsecqBbqUXkYy35xyqBWs6+uiM4W/WCa+2mV
VU0MPmgLQ3k2mg4+gvUGF6NO7XLyqydDYpaQDGIKsvdQOeV9qJumsVrW6ngr0M7A
L8qovh37GqhxWXpApo+q/dEBQqlNTSDBhmkjMutBpMOeSvPdCQ+qPWAhNkGmA6fR
mdXZNVo5e8FrknA2dLo6CWFMLpaZJ5Jv84JiSDsYnfTsftNQX6CKaWzYtNzFsbnw
8RBKYRLFAxQL8aUCEzdSnZz03amV4PXJM7IB82FjAfwGH435vwDrPZmi01+/3oWe
32PpQbdoWeDBzvfAexfqT5RMIjpwMRQd90XXX3OOZJ6bLPF5oBHzSuDGbQJ569rs
p0Xphyqim+84GbbAstwaPtwnxDuX3lqLPIS8uWrJDjIMHwOZcrHxPFs9QJbBSGgM
MFK27RXJSTziauJxrSYwd7uKA5fLjnxTKV/rdsfW6SlsWL87keLxCltYkpgEwKQY
Gmlt8xz2m9dBUwdHaf3htCMLk/G/G2Ecees4R3APluuYO8vQva8UzmevQPmrbrAE
TCsOaFgShrbQenY58T5BebqZYVPlvCNDhzUiS1xMYTveNnmiqs1+eVCpZjTuMlJu
cWhXkx2sVho9bkxd5ZbDV/CSsvcXlSQQPxay8J5UOZIDP7zQmj9yPjjxsxrTStWB
/C4hat1GwHNjL5S+tWRMSxJkd8pcfGTL1VdFcWbudzGNSYTle+7FK3dxxHfDRGXf
xLXR3N+fgsYlmJogZkOzNYHlQcb0UkTcbBq+W0S3wynID3tuyrIVGN0X98kDsxpo
3pKHaBQnU1m+N7uS4ODRA3pyv2IvTW1GYXgoO2dTz0RsRKXgA1gzuuDYgyF5UO7V
u0QUyHQWx6VZzAKQonEYE2DepH7R2CyVjIcb5zDnGW5TtXAOPRRlmBYxXYhlCRjd
w6msq8gweOaV4DGQ2JBHvz+FY4TmBGMEtOsw+XxgrMYUuVtT1LpeBNnk58RYpEIk
JOLHiTMnutaWh26IHKjMzjRquiTzvyWrftOiFup9Jzh5okSq5rr6I003SCC6WVDR
N5c04KL3XY398G1Ga6eL/q9mJpOY/6xjZOCFH3Ma3goGVCVPx2uu+mF8n3lGNdhj
OvS/ZC3uoxz4tK0g5IfIKF7+Hv7nyEmFvFDj5rzLsXuf40t2uk07qstzeAEU9KoK
FZn+g+MkvjiLIdKy/4+EayHsWhpaniNcg1YosmrKGyMxWAW0iymKHTKd67Z/tUYe
xKURKAmJBPjx5z+q5OmKSyzdsVFW4UNFXpY5F4E+U3mPybeZL/qwfdArwWfWkZwv
Gc7Kz/qj5ggHzdIgQKDZ131nmo+YjDnzQTz4wlJor8pKNYpubj12xOdemE32gyvd
tYxp+q9qdLMburoraAxVA7dXIsoXYwN5K57YXxUNjHGCh+R9ZXz/ThsuYCztGsIr
zxszF5JY0bRh+AWBXkxUqw4lu0z75XKtinZ3imq6ybeA/LkMKOSmD45yQuy3ysoA
2m7sHrJrTBl/nO/A/e6hfzr5BUNCpNFe3rIU8II1jJ+33Ulb/oUYwcbRUOgCgdcL
Wijhk/pjSMqg2q9l9FzrXcHxt9v5RVRzZ1rgGLJOvBDrhYQ3pAtim14mLe6rgDnU
0iPgJPWfIab290IjFqHihdc8cAA/05kF+qKF+buTq41BSIVw1pUnfsBfrf0zpXhu
264FLaCWqpOP55haVzYdFZ6Q0oyQQUCP2fUNYWFa2rfaoqCausSwHudPZxUW7POY
6S4+0sUdxZINEvPODZySJ5EoNrW6YwpJdXViNVK50fKFeJbS4b4OYfCv060XHID2
zOBCJyPXoW3gZNyRcQEYNfktl4cVcv58p57rms9UMHY+7dKo4ZGHnzxYD3uG6XTb
AsYb3HGBroxCLt70iL6nVDH04grrIzk1A+E8vJxLyoT9IwH7c3hgNYzRQdoGomWD
O8WDvmxK7Yf/WZ9GI80Y+tKfmGRjAsk+PGnKb5jqiVEqGM1vcRV3jJSRRV9bBSq8
AmM6X/01XwHajpGseGFLWDQZ1k/6vnebAV11wn6sK9ihaML+6HoGdkjRdv3ugTIF
wuAE+vm9YGLeznEDOCw7OoTtbBznIRVyUiulac8K8GmdiN8IcpZiwrGTx7aL2/Xq
ZoOiGvyfOIOJ308X5z2z9mUyEiQMxElKG5R7zLb8SN5pVPtAkWUbOK6P9E5LlgfH
bej2PXPF1w7ZV2/6R6+IlcgFM+V2kE/JI02CcBDmd34OnuPAutqETSBO2Dw6Bixr
FLKOc1jGiW1j1elblqVjjywao6cUcdnub8eMSYbbK/c6QLSugFzGdZ1B0QBnBNr/
/2YVCsrW3vFMTH+fiY2xJmQ+771xB2BbKI22pVeyUFhbKUSs11NfSwBMzJ8vAEZW
YsCjotbM/jWA+fKzhHL4AR9hz1d7KzXSg7n0nBIPbzsAvjZXhoyo64jtvcrT6TGQ
YVrju79Xghi+BAQd86mUQQztqzo6Lb7BZ0fx8MaBpjFYQMym5UF2XFmdFRb4X2rT
PBDvclACIUP6LUllzSC7fu8cB3EIVMfbTLCwPrvwwx1pCc2vjT6bU62/WC3dBH6v
/rPq2Cu+cTuGuXR9RHxMQioS/l505KlkI3e6cx5z2O0BRF5gsXwDQPa1b4B9sDLF
mFSzJ01dtGjUJ9OFclW3RZa5EZsO+pBXndA6Jy6G4PSUNSjvY4ooAQu2hRAVr42I
LLJbSMv64q5IrtBkEGL08f9weH48+qC4W1ZRHqgQ13c/17XJDtAAGvuRpgtgEm4O
nyxvFIbT6+RRpcmpGzd8NNNXkQTpIrw1zbuI+0CQcThTMK2tw6DsUAT9Wa5eWPgT
JhmRTeWwJfe1XjfTIRrNPI2OI3+8PSTy8rdmkQ0lhQQUMBmChbAwr9Nfs5W4VWqa
8NB6+hngdScVqbyFb3sBgpMD7aHUB0MJpw4WW5WyIljUnL2MoGuXztlRsFUilrHs
8GeUfbTj1VfyyNvPzHHlms7muoev+pbqXjCfXg7iBwNSCVnQgyCKEx9mZ39Yg/p4
ikCmX3R7cesPqTMNVGFyUB1yqkpTJug8Xu8JjmBrkYng0NrPhWAkMjz8/bLwNuUv
VQiqD5w7orjInc1etk+hgXxQPxBk0oWOVXp9NPJA5p9OqQ8DY2juti9X1kJCi840
XisKJlMPP8w2byaeH6VOWsz2AWoZ83ja6jcZMV+aLlM6qMqnLHdsQSeZqKZ8GhfL
1PqIGoY55NQ1bTsAy87PnVp7Kz/oxPP7LEpf976VOjPMDc2ME2r8RgWs4KjFBe4R
uNrsvGiupC1rR/86NrOlPlXCx0QWYyGVVdZrP/ZKQficlKD8Aurg9r15rXCTXOsg
3Bm35WpGfUAHgbYoQBHIW9sf+DhglYLBN8sN1EkdR8M6b3hwsMR6N/mS7V4e3TfU
A5VmEW/AAsEYLnE12uQcArvv/gt+pIzTEaJjQOhhz2/SScKijMWwwxSHVIvIl9kq
ncdjmNTYbY361ZgW3sowB4vcVH8eNTOMk1XbM/l8n6G/GYJkkTxkfMMZXRPhV1ZR
RdLYWDjpOMfVICSTFBVMdHJxGoqUhA61MurWsJ+zffRjU7ix/efUY7qyHSD8cHBV
1TFGFtchnWUzAt4rVcWdh9x+dZ38BzyNr6uBIbmB+YzgV6CMaCtt5loqTVEtzUrv
qDe4hewXLMEk/vop7/mhfsDcKfxkwwnLOFI51LOS6BOmBKwR19bNgvFrOLS0qOZG
qxKpSutigUCf3gm0nE8//YHSY2zmFUBqzbnzTq5VcGKc61qLpNPLVB7MvraA++Ys
qhQAcbJRmfyRuSB0XU5YJ5dzbhOik2++V+cx7Yt80LvSgbCD8k72rvXy/4TunfLD
fWmyWHCdQIvyEMW2AD90pmBlITQ8ThSGfORJwAPaXQrRNBtxaZvEaq8ATOJPGbWt
JgvbGRkO6u573acQ6pNhZHhG2PwCYwgIM7yIz92H+Dz5h8ZcYSULaOX7QIh9uTNP
pMM2ZYVP2s2D9jJ9hEx/TK8Ydz4yEKxWwQqf5sWCIckPal8hTl3TGSUXFUoYfZS+
b+KUU0RS7rQmVa44zwg0mC8TP0IjTm4iLGugN4eKaYs6SAURZmmsA5n6pVlHflyr
crJjjXp2RYlHgt5uFR45j3UShKGG0Y4Wm2zWM/fafoOJj2t6QKDf3t/z5A7bg7mA
LozvdcCgeYZiw8t2pja5GCJaKIVA9vFb8xUsTQWt5dbqywx2O8THSwCqgH5wLUyy
0BEc0Yjx76Tf702ybBPzDJ3yVhFNJcRr3s+CeabNgWhF4uQPN84A0JLpsNTlQIK/
akJj91DKp0V5WFrcrkvGZMX+iw9O38pAeY1EyLMV0PXgUsaQxgHkxRHqIlB8LH7x
i9T+8t9AZwB6bhmtwwmCmvUs6kzC67hcanq+UerZgNEnlfBnRyQzcjEmdsyIH+E9
RxcWAJpso0c8Y410HiY6i9fdoJShB6LveNGCqvLPa9awbAqUZu/r+po02UJB7/mU
fLNJVFvv/vCvMWqc2HCKWqw948KWgnU7OmNXKiiIAwbhRtxR9+m2FuwiistJWytc
u+ZICbq2g1RZjjKgY4PbhDO2mubHa5e/09PUtmLcd+y2xoyf4opj5zBGtos6eR7Z
klcjiY3F15az3vtRFxcuas40G9nxzz9Z1SbYBzy5P02pATBaOXbrXkzHK6ELPpve
OcyBybcJSKbdXZ6fnyurHbh3+BKDjQCUwpDMauyN7ABVY6x1/xOyq+iLPK7OMVDa
Lv/fnU+hWG63o5Z8KSMPUsdTfni2Xt9DAtMCTto0ifWg0dP3mfFeZBmDK+JQfCFt
00q0RIbCfNrqPiSo/4m4OHWT8VzF0ZTcmieWbn/Lh/5uQeM/cGEweQQE2OUB7jsR
WvwkxtkLhRER7t+1P3+Fodn4R5mXKyd+RIfadlgYOD7BSHsiu5q6aseW1co1tkVD
5Fm47EwPu4SdP/nRw4AS+oSaEPWPtcsPNNDMaWJb0Q/elxVNVD6bOp5H1cnIQT/A
XGMaPyvJzQDQ0ldESO8AQrhnicLxuKpIrXkMaW3wgKmfcT4q2emCn4qdYVmEueS6
uxAtzsjWCsx3sosLS+NVsjuPVIHBWV1iOocWv76Bu04jO01Jr8jT7/dics6XtFQ9
xBCs1Pry55YBm9kRhZ9SmdB1aCyPcjaKBXCPPcoHFqfBN3LBci93H2yFwaWhkmDI
7vLZhK4CssOaO/J8uHJ1zvOnK8PUDvI0w/2WOPDtWjX6ILdki3Z4XxVNavhlDFGI
u+OaXXJEgvEATSxzfIsJkm0L9MrGjCimzB26MnsG56KDC5WoKxfa+PAsjzehSRKX
th4DeYsco40LO6MkwQR/VfGlXRXQLTnYCNHjm/Or9RE7h9YPCSqhqcz55iFXa6qX
I35Ih2eGs7Qw0QeS1LIp0B8+iVy5+pojhXLGubDaAuhmtit3bk2z/UnveukgvRAL
aG67Eeq3wsPOcJqz35NPeOgrZFnD0IlY3yMFW8vJ0n5sZWD0fxjMER7fK0DfnWY9
ghsghHPzprQXVNpQ4cUQKUugPZnVBmuADDGL9DqKHjDGQJk8bQdatfJ3vYScgHjM
UB8EFY2YbZ1fDqrxGxEfar6OU2qcbpyNmmKCUndNqGlLwYAd6f6ilsiO6OXY5Tz3
+5087hdGfF+ljDjj1IT48072G7Znx4ZhlX+eRuXS/G7Rx2VCTJpER7DkJBmZK/8y
4lHpwWpFsbZgyDR4uVA8+/eyIdH0tAbTCGo1w2oOyU82S4WVEGAy4Y15OiUcUZEy
sOJEtHwxfcLSQCW7tDnHRbmia93gSsllwr2prt7KQVJ/E8Rgx1ChIYC5AS1O2J65
TTyBD0Oi6wgZeggejeX81E6y71DhQUvatP8TZ+gPDd1Ae47zQgWx+Uv6l9SOL8CN
CD4r6RWQDS4TObhF8ccUCl6q2/3+Fs+ykQ2OKGmxW9gwMtjLzWsE58kOUgbT+4n/
aM2UAeMLWiHtwJp8hsolPyGLCXKXQlBeL+bN1ulp4xNv8XcgDd/JOPVVRrMJTFTr
+7h6kf+1uYP7bFKschyQeN2TOrMtOCEg/PWTZrO7gfF6nZ+Wz/fM+KIWRAmQbk9I
MO3VWTEb75b2E4Iga7IcFUbzSgjTGFofgXEQ6xd4xMgrwiXiTPlto1+Nptadm0gg
FMDpbq0hb2QZZuJhZeigiIiM09zFlDBF76Brg66Ye+tePiUh3rNyJdMVkmjOi6XO
8kPcFEUm/neJ5oFGMilUXBE0hFMCI809tzlG7KsbN6P1XpWiyCgdE3q7gCPNH0Un
xKCz3AsRd4mFhbsNVrDukXXvmhL0Y/1veTl2ZpvoeMF8MZo80EHrp/8KEMpKSfp/
tsBTyc1ttLSOPe1Wsdn7BIy32ERpnEuCVybr1u3smagIOMvIt/8bld5zGHYZ6oLH
c0H8yY3+HUGxk/OXH9nhynoj69gxYDNoLJCFNSx0IHNFbyk6v6dx8of3WwxPK2nZ
/d4U8ZFaOyoOpgcuQXHzRwbsYSdGCPb/zuR92qTxlQrGNjWj9sRoejxo7KgI3YoX
QYPamh+KrxK/Wn2bu6y8f8s4eQrwzbosw1b0bTZSdXmbQQesFr+lXGS59MdlOK//
TWJH2l8lnpUz+7RJ07vwjK1SLCwlOj2USRcp3VDdocqVXhT1tFGuZQEtloG59qjJ
Ezdd9ry4Jt6qOu1e/f0ARwybNZXDvEbIhmAHfGQMIzlbrskutFbsy7217byWZ1/Y
EqUrBg7wTryNVXxxorQnHw1dMP4DJ33Ew1jNrSX5gLWqdxAsI6iUgkHy5LvHRAMJ
rq7dsc6d4GsLmwX47xOzZ2aTx6HdNFO9NLMP1Q4yfvoInQ9vci5ElqFfabp2s9o9
e2BGMWYJ64ME7NC2d1nBMoeKW1K3unhJFJNiNm3ANdOWzSlGgVOk0iq9qLME/SlS
J4dVEm6QwL+qdlRbMtbN4OPh+gC2VoQEgVYl8WPnUBQ7okqQpZ6fe7YRaBahSG1u
Vqxf2EHb0IAZiyBtIELQPV6qbqQapEGOjJr+lx+8Vfc1tIto9Azb4XWbTGZHkuCM
ewkkcYOFjf7KcCAiKkIlACH8JirrCwGdNY23pdCTDLyW/gMl3emThK1DhN9W+gdY
GoUABK3+g+CxmHDlIEeuM/dsnU+jsbbPHq0fgIclaPAQBS6VS+6XzZ9rSdYvsfJY
D9kXnj5XuasasMoIT7XYE2Y6oRGl9Ady9pMCeLyyyibbHrn3WndsX/DqPBH5GjT6
78z+0N1ox1iEhj/byK8tTtNKo/7C6V0zrOWJELCYaiqoMoqxrPbJCRK41tbrKSxD
HDjjCNXIvTfo/VTqWhlFi50nPWgLtv9eYeoBfWagkcdS5Zx8JH+Z7I9gw+tqe0c2
204iEzHcgw02sOr5b5VW3tcTDAQKXijUnRPKE2Skm85VhH6/OFDx3rJ1LgHM3BNM
9m1GIbdKg/0HzQ/PyUFdUmoBUkA3CO6xC//MCnO1LHDBOwnKNDBzfkALvm0Bmd8U
0+WRFMR8TQV1dX7ikx2h/gDtoFr72DH0zzMBwLljl5kYgtnNLc5tLBaW6gs+P1YA
0DdOc25xieJjBEx08xNojCMyM77b4xVjN5uAkDphSQUtuZS7qODD+vb1eOWaDiqs
jeO4HiQYZniWlgSUeoJygLOXyyxFKC08gc1rR4J27n7CJhfav0GAY8Pmpn3ooiSk
NKRWIB1TIlrJFhNqJbTAEnNejhLRudax1ot5uGpjBEQmBGrT6U/ttA//cHBdra0b
r3L+Xzlub1bSXdJu+M6jGzUbZhc0PEO9y5JMdsE+u60aXsdZWk3UAtTTZAvZih0f
Kry+TRqT+4TDR7gcE2d6zHZQc1twaeLQWIexPhDVRy7UJYlonceLFNga9cbUC+1x
cxUhKhLQEf/hEHwW1kczti7/CJKvFLtWc8xWTO/Jkv/JBprELAMTbXCliqAaj8Cw
JMned+TMkXmwqekjAogVww/XxTwiLaeNFlz1xOP7HB93GVtNq87d6jqBh1gypvLl
CQZMq5AuBgpWnyYQtuibq7GHKcftwoAzcbQIQTAwNhx6xE6cRnopPL15fysX2laZ
YXae73rk2Os6cxu5hitOiRaBHyFCsD2fGQlNNB99YnKxBehzV7ZU4lJF+CKvQdyM
PhPl58f4R6BuV7TESUr77cN1LT9zI33yzwZLWsTnjNqEHWlTDtHEoM2Kwfjm4wQ3
yMxPjb53CQlsxEGdudwjbAF44Ukca1MotgwooQ+nxYklMuKnIULdeva3r6zc/DOy
fZ/tH1woT6blrEA0NTmnmHfuzXK5ixCCreuRn9npLBPx8aozQm0d/YZoRfZ9S5hX
vw+X3Q0S6d7A6M4Q0iMqjCJOacyPW9EeKqFQ0ova25tht36rE7yCntUHyIkzLp5c
RJStL94wy+Hdzk7YKdOysZifuh2CUw7l/0lvYDKZBBV8+LOVNM4c6x/Hncanm0XR
JPW2o2ENn61PbUW0fTsljNoe+mz/Yk59ggOLrPY07soUvguP5VPeBA8kBzXDdvXe
rSd0om6RuWJIwIj4q7UcWUw/5eHGg7bCSP0xmNuykjYKXNrmgfUxl2uiV3KmopM3
ENF/IL6O7wqvpBNFtNLkn97zuxvrhuBGerzkvzfe40UF+EYCAWUT4PhjZteJjSZk
6r1CZLGZAnBCl7UMEc9chM5auHj82ScG7S9JQaKvXNxdjrfMlH6q3cuRWYL/UAIu
WlMnS4lluKlBhfAkMdjA+o+rf94CyJcCPxDo2vDojG7c6NUy+UN21J3ThPosNanG
9gl/14Lt1Bb7CE+Ly5B11XdbCN9UVs4lrEx3CakWnsT6OdyRQWeVMexWlL/BsAqG
YrNkoHvgspKUN45wqXXoVIlMm7HilxWENoUJNVsZHWhE9Ua1r2iHh6UT+BqP0Alq
FfIj1CvQUKQx2TnGkzANTznib2saWTGLwdSQaLZyniP+AvEu4CtS/nehRka4w6kd
Cy6ZXSW4OSi6ZOltsVazQ4eck1ickQWI+tP2F9E/xUtXEaxrMs+3DFrZIw/LaHHC
nXqpqmaXg7MhJNMYiMRqTvh1Z+928ViWzyjs/WH99rLBCsiKk0STvYZkU2/cGTQD
lnwK54JgxkTsa3t2DDcR9OCT3Gi7Nd0C7XA+eqC4itjcy+q1n3FME9X8IsZc3Wcm
zwuy1f5ea+eHn9QU2lJkvqL93eBx6xgy1w/oRgz1ozezXXj3V6n1QFWWUR5noA68
8fmI4qrZKkpT8b3Gx9X5h1txieEfTuQ5I9cqfPP4cEkMMh5mKHSAEGONtvfJNmQK
mt6wV4KG9EJfEP12GCAfL2e7KBjfjIMp+flDJ9GOKXqkF2GrS6u7Ure1g32MGfA4
vzSBfgWha/2GrZICFmFYhyFJxsL0XTv0Ijl5h4GFlqUBJS2w9UE10u0K8iNfxFUa
2KCuTjCfFvar8PgWbDnw9ldtPXfwlPWOgII7z+lmrttqG/CeFJEIFGOvmtQOiRUT
V8Fj+a5QySd+zZFZ1+FLAqUJ8NX62bAgeOGfMSU7E0gZckWM/L2IabckHEX5RfBY
e4WBg5duo1Y/r3GgotRMZZdCalPNndq5D99Dib/rzYfSrcZJBEFphQj8+5yIfK81
pKGGx97CN9YLpwbq2Z82mfakCuBnFUNgO/aFm/grmkhnrUkBoBNchulQJaNZ7wBt
RuribhcmXon+x16GWxW9LFLQCVNRYYPCVhrlGjEARvSf+9tGpaPsErvOyyuzOshQ
sIRz0XLxSwM5hJ1UYOX+plaVaOY/+W7fTfLtIplRsL44tON13JkrSBXWEeSGlMjw
wew4u/xFLdK6eK/csFpNUfJAIpn6LeQkn+851keYGJ5nUCKiwKdjuSUANLgKcvII
QhNiFrXBS6t6w6AcXs6zs4qpVOLVQaErL2FGoYygTiN7HsLiSYDsSFyStQzPDyz2
WMujkJC1rcJhj5joC4tv4Rk8aoEfyBmZP5R2SKXcueri0tqpbxXRSRBZAoQ0t3uf
YAR9RJRG5vVAKUlavL44K1G38JbXz7jp08V1bcNLirtIR3KFpvDBX351/spRkZGR
SdUevqiNOFNdOfMU6TG5EDmxfPytWsXlNzQorH21ToxvvjueIDEW+ubMDInRPT2p
UhfTdk4GOKR82IzrcrbGz2izBgpTXhtFukrcioolznL2N9gBKorVtiBN1ojyx8AY
CyHgQBbzVNAHUL8OpT/8gLO2PHp3jNr1VWM6bmQSqk6hM53GYGiN3+nlhOz8A/2C
AhkiBtkgiL1dK3GYzkvEh112MGAvAsOeXmqxZ8afqOp/a8JmAkKV/iHadXgzxz2e
Kg41LSYlZ/pIGBgxerbXj+JqPkbbMeLMYOnhYZt+g80MaPKaD0j8OCL063FZiw+y
+W7CO2M9mXMm9EfMHnAKV35Cj/GTcz5Usvn4qzGvr9Oz0v4h0v/m/uesWMzF2Pi7
V8VQNqLWGO0484Tiq7Se2EgdVAvhN9HHW1Bi/jFVdCOfeWJojQbgEI7xo/X80izw
22nU8s94abseaqCz5S14tA7tE6JgnGxSvthICDzcuZtQiYPU8vdUDczfGGnGy3FG
JQWiqpCMd4W61Q6quwR9hoqifzPlHoQL3pgPDJk8io9kxKgRFE6W2lj+NDrlVlfy
bzDdV2WF1oa5K80m+qU5b0hWNM5lGmNYdymFxH1ZXm4oxsci4W7NiZA7+miiZkMu
KXaKv/f+WTWlMZ9rh+yaPlqef/x3VuodCdL7HJzZUWU3UJBojatQmBLTJg4RZuA+
vfbFIf8L9zDwqmDVxxceSPd+MmYA81OkJZGgT9f7jRU5jDat+41RpOq/dwUWFpmN
yQTF/kRKZnG37flZZuigdFpRqh3ka+mZ5eGYlo96pHW5jWL3L4Xjq0C3xqiBG3II
QQTfzGLBvKljfVIz6Ah7Ecc2FFF3xGtpe7rBTU3AzhA6Anu3yDsxV2iMmSz8c2vw
IhtLh7FoCknNga4xJOzcCPPtZWcjLIb7TmQ/TFSD40RiuL6/C50HrTADbR9AOhON
tjyvPl0rvb4HIjJWg/7L31a7QF6OksRdJ5sSP+tBSvZFGMrT+9iIvQsntyrfCEj9
3jAgAsGWvB2NyOecoyQx1ES9SQPG1SMx/EW63bqQHz7tGHkimB95f0i3KLIkfvud
thISlFPItnIj2nFF276wiqKc4EUJel1DL7NjENOpJej0kb2KWOK5sa4wPDXGe8oj
eeYSnpYmyMFNggBZY3GCGAK+T1OlICyX/NEENs0CbIv0KvKGf7if+74V6Uz1mm3y
rEGBZu/ZIaoI8Kq5uL3glnQhDvcMaGHQTyiSmFkREfwqi0bxFIxMAnXdS+F/rCmy
oWMFDV72FWkv6OptRDqQHfQdRmyrsXV8juNFlzIUr4cERf8ji0B4fcnyOarzAy0h
lxy/dR/k5YbN93hYg+dM7eKA2k5DTXJh6Cmapn/CM5pAqyX9PigUkKWRRatoIVGu
syU6evdOxnuyEYd2n1yBA6kVnWQctwaxDuaAfVvtSof5h2/kEQ5VpztSvqUb5zEF
2HhF7V9suGCY8wJ0dcHtumwDDfq0yig6B9JD51H+Pj7/GG6mB8xUPv02CmurX/6B
hBS0aDJF2WADsLxN47aVRmgGIx4dg3KISSiQ5kFaMe9ntm37B41OlFrquSIj1kD8
1sKcyXgHhyPGwiqxO9sdUiixYTsdxSfey+FF4bI0kI2Xfthjn4tiGpVaQxkNo6/Y
4nxtn18TIjcplS758ooD/jnTcoWlAixa5y7on4g7DvNddy4hz9Ev2xOsn+I0XyW0
AibfEBKZpCqTLdN4cPuIJmgjH2Q+DlUEoX//rkvXGULQqVSMCgWZyesuPsLOx9oH
8uH9MOOaUXLbzq7MYHlcZGhmRoV3h8HPHB15WJV3ERHCTiZ09WcZVlv1NSU/adFl
OaLRVqsA3Jxkz8I674lfjbGYiX2ES03Tgz60/1FONPZmFya34loeC7SAHm1BiP6k
4RNpOM3UCOamGMv+CH4mEBfQhcWlftl03QZPaJNKhiMzYtCuZOgFyKTBs1FzcOGN
pP1cx9AWOB4k5SJu2u6bcrt1YHJtEtJwTDCAzkpz2BXgwgImQpG7ZEPDvYd0hk4w
maa41VLHub9YD9bKAB1OPM7MskOejArLbB70Wqk5b8yukCiULXgTNR2wqByIR8Pf
h3wPvTpDHYp5tsWOCLE3DPO2lvlm7tSY7JOhT5hcNGfoHOR/jz26x0kR9zJBJsbe
Roj2R2Gk/KKw0IhhGRhhI2ReSZN3KW9/2JFgRCDbg+7VdRqmmMfEDp0s9oNlCOYd
ZFcxKB4WdL5PD7jJGpVB+NdkLZaBgHouflXH4rC6rUVP6UxXP4LN8GN2fgK5Rd36
fAK2CFNRr0HN8iDfYIDqSFSnIhmwODZrXXvFGMMn6BlapSEoOF0tq40avpcpqCIT
OfDzotxYYwuQRoAn/gWFlXSo/j1/qgT0gWF5m4pr0EOgGk/jqOJ2HUBTEA7W6Jtm
Tpt7I5G/Ut2YddNR4MfXhfMyBwqoYpR8z1zJc7NvMV2PFD8rBV9BR32+TgoD08bw
FVTSXHXY7vtRrM1D8u5U5QkS3qB85/9hQIRs1DOBJ4Mp4bVPbtG8ONrj5+vVAwpA
mq2HGgMZ2wbv1Z41NLmYU2bHFspIE75k/Xrp0QCcPrZJOT7S6Cqtm6rZ5YfF2cFO
troGfXsLxD+oDZbYXqVbIiHMhvoa/vAsZ8MINvs/fNHUkQ8FTgA+bYjvYg3nmmtN
840hS0NceCM0egGdNL8V9ENaTCTDsWiRLgtjcOvZF0jGKz9R/PwL03W5TAzqx8DA
2TZtQPFUfPZ+Rx6iSOlCzd03gJMWIAAXWY33dg1TqAJjMNqMcUJ34Lsk8WPwLNBN
TyODRcUw6hVmi/+Wvb9NxGZLZehONNv0ajWAoU23i2gMo46aKe0nHvn7AvrBQWQs
333zUoZHQEDqD4ST6Dr32+h3gtZk+vae5HfRnJW4Nn2qpmU8O35Y+blfdLuvS/jO
4BmUvWWXsSu6POlT0zjV4kOmjXBWwZ2Yp1uEe/ss8pRr3ma3y5siq9mH17Bd/ZzW
n8YbqDoZVsIs0erGJ2od9fXKwu6gwvpBFeKNRoIyG5Nelqx1f/rAODxR7Fdwu9Wm
EcAG21TWa1kfRDuEOfz296LVV9zhr62nZIDrJYX55qmfMJnII3ewD1fMjaJ6Jy3o
nwNGNZW4LMPmNofQ1Y9scKV+Ionbi6zswiYCllMZCMB7ZSFUzHp1fkS+USrPcV5v
774Du17hoLwVRb9gHRcKMUXHR3UqpQcV0ILUg2jF3cjjvz4U7XlrPNYEVnS10wZo
8PEomC0bIASziBsuc20VgJktwZhqlUGaM4ib+DAa94WHjk3cNf8TZWvGS0XxqwyJ
dYd/HpkLWpLJ1Kzg3uG0KWj6YFHlKdOD7F6YFSIPs9H17hmV+T198EUoD8NAc7BT
UnSB29k9oiktcV8gSV2nyTJd3C8vbZp83ow995PqgojfGXuCGA5P9hdoV6uobhzp
JP2KyswmVaXu49N8Kz1zFjKswVA7UQObeKV0qLBIRwgAcaY25yvtkVZS+jNRPOze
0ZiNBh4AHGBooCsvG1skM+gP89cbOUDgV5nLxXP8xRzmBq4pgqHz6+jE1/8Jrh/d
/unSSuVrmY7IaESymqPO2uHQn30nUNsZt60Lp5hShOjM/TthhScv1mRXkr8bEk30
2L2A3UUrH3MoE4yWah+KyMP3lSGQZTsAyQm7t7QO3vpdAm54Wo0cXSTiRd0boWv4
n76thX0VgmFfHj0uyT6rFCYtjX1PXouJpyVJUjxXDAJM6dp2p2bA32jQuj4FPReG
O8EPo/PouVq0IywE70N1hcLvUt4PAOU/u3OqIFCcFISCn5kDlaUhFl1eXD7DOMy0
/TAm7jjtwWYZJzIwYBLTUidWgOEciDE1+4gEmEWoYkd1q4H5vGuTCpbbCzL4SXqP
yuIf4y7sctFTJjHKHaSgUA/WiZOmRTjDQxMcw5SnYErruCmPpvvH/egEVNBavf3e
DIGNvw6jHQUWvbKsuXj9B4tAUaR5+7K0qTRjgdbDMCBPLxu49JvfTS9ID71iBgUs
TRx4EY1GbWqiss8fOpPneLdqQL2H0tY/RH1dRf4Qku2lxAPIZJ8ecjzhC89jCiOn
GcWyG/75nXuxJfHsaR+IlpANe/Fo2qhfLXVWSt3Go9cH2n78hob3ZOEsZmlkDciF
k2onZUtRUcKhn5SPR/MJ5OIlSXE1s46oaW0At7WD6copmVQEWeg5grQzo9w9xYUz
2lepZBgUKfihSglxMBgxqQN7vb63ExI6jKoBZSoHs7CQ1CE6i0D2UhSwLdceCXI1
vcuGBt+OFrzBLx+d2rAEOySqsYDOJITFKrvjnXUwptVN1LUokP5xvnAxfCc/aZzK
3w/AzwOa9byWydAP3sFEHgJFAEGowhE/RRZ2AeFAZdZunRlAYed7ixFu+5XEwasQ
p7tafFAra3YC+yi1j7FBC/5YIZtV7pi+SJglHu6BIpk/MVNaeZLlPYfGurIZLCeZ
bP5jDKClQbf2L6fMdYRBNyoW3NIs47k1E29+lBGCZIsTjx26LdfolCj+0SfcpspK
M5SZ09S6oW7X84GTXLaPw1DYkHwsy2v18Uyuq3tzTGIbN0LkrwWCjw+oJziPRIVF
bvy2BaenjWpysJ22bbbpMpXNQkyuhQ59IGgVlF+ZdF/Q9VMu1laNDMeVu5NZK43J
maaXrT+FKoasC0peQs256Pay/tNWgV1T1w8Qsq+H8XGyKVC7Ul1k9uHKWtjk2EsM
5CtEmvnA1oXRN133mt1ha5xA/Z09FJz68uYPcf/5Lxlu9Cxty7h6HG36YsENEqD4
CzIMlHCxETj9uS7iGZN8TG7R6wmmqKjSOcUAwSI7DSdEMNc6pVaqmm4d3sq0mAE6
kjVjFCAsOLo8BZ/ToQPVPpYWODg4NpvB3LnVIgx0jBoTBKvmYf2eASx6QtZj3pzN
DV/Mq1mneYuSbshSffJhzYgtLUYMnZafRAS94RBN5fnh1g3wUq49qna/LNmKPd3Z
HOsMgAZ1MuiZ9cfoBI17pnMJFid+oCGGfdnSKEoDEPoo/ff6PRbSYIl2pFFgZ+sj
jDjVjHPPgm4+r5xlqiuj50B8vQVwZoAZW9BDoMKVx2n/9t0Q00bCswJI63N2KIjS
fCTibEDHD9/QZNmHGfKfE2+UX3NYOKeeY+p0iT8rvOjpRjPdSjh9s/MpHNoAOsxE
6q817XSjYSkcWCfefxG39Zn58ds+g4GRA7J7bgogGxkdnaTmB0Uzg69bMSUFydEh
2R7xR4fLEHs82qnsLRyU05ZKBQdBQ1If8yTmhzQ0SYCG/MlPiNpKGnIGWcctfloA
DE45v7YQKnt7+CbpU0Myn3WCuFY0PP07sidGF5QrXkYTJFApEYbcmt0kDmqXctmy
jeiooHruqhJa7++B9sBWPszp1ew2Spis1ldxe6Q9n6Lk0FhWlgHjjVECBPbY76pk
oceL/XIYqLSZwSzrSLLSFZ0+xM5sp2lYeyU0qIjzBGT/258c/S4vma4ud/gqLMV7
PL6QaLmoin3ZsmbK6jH0spGqazaf+h6+iY3Olorx99BA6sE9YaDAXNuYUYmh5K4M
ZrVjF9sAWdLpFDvzkx/i7lynU146GrTXC2UWyyOw2X3QqRBlZKzvwlT/jZWqLYUR
BETdjeeGrS8Zn0Nhavfteek6e6H+YT1Rwekf5UqLdC5j/4vs90aYkH55tFtVDFTl
818zW2M334ZK7gB6rwef+lyYeTQuR/JSND3IimnPnUO+NUSgk8GU4NWzTo9bbh4i
2e5tMGfVePm56ugNSkAG5QEYg6t2aliHQgjZeKr+PKXFDkp2INiqMn09+VtkJPNo
uw4F7rKXhBVMMRPnmhkSB+4hu6Wg1DzP25iCI2o5jYNcrJtnvKhHno5PZkfWoEsa
Pal5uihISLfY2lD5DQc3XJd0UmnhKPWCa7Ty/lvh57fawnKwICeUGpgEcQd9bvOF
5mS8h7MOthA4eGgZya/z4paaFan7lGNe/YGoeDOlO8qqHKYtjt0gMRwQSknNW3gf
reMSxQKDnbLQT1H+UADCIhI4yJ1EQBaKbysWvayTWLa4BCiJAr1XKt026ltfkT3o
EL22Ty2JZpAi4GtFx9BHeSIoJng8HNo8pUHlVMgimTP9Qn12z/iTRDYWuodTIQrb
P2lAxYSVDMpdo+FN7W12aFroGhV392O5eW7J/+xo4Qp2GaLx8t4cGJPq1HNsJyBv
d5stfkd0Z1zTf0XY7uL3FSsSBFj+U+JPYJ5026PjMOs7NOBimG/IDRkPCygynL2j
JNCAkB87Cxh0AVlzw4nG40sDMb2evT65rWY9oCc7cU1EijKDXNwzrS5Xt0DP+IvG
9lV0oGD/omCrRNUW/1iPF9Bn+qLFsy1BSr1sDJ7uuh79nol+VbMBeBvch8u7Nvrh
5pPhl4g66ocV5iLHMwj3YwIEe0qTQD5R2vK3FXzmd6dI27Mx5xf8IYilgT6DNjWy
oL1PkDD0w6eKKnMtKt1hlLy8XNhXgmWV946NoxzmQBsTgtrkWwnroLcQvCjb2wO8
5RuIGtv+yYshLMAKPMQ3M2OHnPwjJXLq6HIXN0V8ULmqHIGh9Yqcd0/yxSvv4hcu
6sdTeWgQiiRpm0IKOWP0MoFifbfSo5cxvS1XsxBwsdGsh6Q07xoQnHv0r6WoR/Wa
q5y9OwesZPoa+gVIDCEpx6TTwva/4dfivB2M7U0wkZmqGbqDt4Tgbwnc9JlTKg20
tZM0gESlbJ7fXRRDRURdDTB3Ylw00pE7vwmG6yj1p+AWo4TiUSSOi3ymFU5CC2Qr
566UEUVjZNblat63VllRmDT83tIuLeQOl0+IxU2MqPiIu0e0UhEnisjiV+NU4tNu
VZxx5NrBudOrwpZs/7Abjqgk7jcJBDIn1KTWbMVLFSHN86SDAmj40SuPKt1HXUAo
R6TPJhflTVrEgssIRJgX4gMnO6Iey8jukE5zlDuNVrQqoILhw2mxiMlyF+gjSWhl
IBObBA8Y4BO+WoPhVxX4GsEtNt3KNa61Ruh+u4JsgD+MCNNIzlDNCj3mcZmgVy9z
JYAJuTA15aoJ4LMFE8F/gUOcD5qaOUg4Em3D5JshQhrq6roMg9Yh6HSjvPoW/bQ6
bcuzWY3uH4jGnk0DG80u7t3WNV2fMqoSW+Ra8BnY8ChsQilJGRANPIbs1/hBWXmw
SH9TXxde4IMJ0R/RC59pBVkT+8V+r1Un+tgIaJBH6UbEb2/5+6Pfx80FywisfQrP
amduzQtHiAspKUBBE2yhRJh4pX/Uj3+A28pCpAF7/Eq1Ayu02hfMNEvhne26jxZf
cgyKm9kD8vEkNTJIeQCmz+7dNY0yZ4HzUjSq3ceBbwYak0ljXdvLy6CYUR8sWB0q
AQq9DLP5zbyOhKSJDl9pN1PUcJY3KTEy12yTURQR9+2ewEewU2QfvCk39twESN2A
cefXxRqqlJLaE4VSKSc06ZuCF+6E4KSaSFhPN1mjIwSY1aEbXkdYE/Hc/RtQ6HbX
6EXfGrV+ahurw9UzjMVf4TetLN/O6lDv4cYJ4C+07TkjVVIuTjoLYkJBDoGrpybF
BUvZuI6lzpsk4Ebxz7op0Hz078voG76HdCLcbcYLcYE6xOPjw3wvqSI5JyrNzGFr
6bufCqOM7+OgEUJPJPmMCDU7uh571NbZ+jqimN/v5DAfVafOhAfjLL9Ma/BWzcfc
m0Up0zCOiCp/HKcbz/WllfKpUTvoFyvGa9arMG7QINIxFsU0Stu56+ibN8SGpXEc
ryeWa6PwayQXRfRixDhIgGla4idWO28gXSSwQuqnpSDszem78e4NrD1ndPn3bSqv
sqSWi5Tbky6SJlBIFifQQNoXFbmSj/XoRWlz3N+/SoUhIwHrcVMB8oPpCZgvJSJL
VyaKp9p8vzrPmY4l3mDhWoijiSpgusf+ZDh/WTiEVYFk9xzZKzNiu0bSwPaGLjjK
7o0/8uFVgrAWqb66/e6686EzOsT7GAFoWbNqh0o7H9rKGhpRri9IFJufut1UobbP
wnip+BdWOStuVitqCUqS1rANhZgVvsNbpI1xHKkhRwpRSQIFZHTicoHih5wtgrSP
0aq58R0eRDchrWD4Scmt37oWcwNElFiRWuQCLAFkWzCCS223N6sCxP4vsnWhEJsC
`protect end_protected