`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 19632 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
FPPR7ws3fN+RQyk1V5tkgEsMooW6zJ8gNY8J24fm6AEeiUqtXBtyOmtDCYNUAIba
oKCRgYcQdMPFQdFDyl0Dljw/wHJlP1jgVLym9OYL+SQBAkXHpx5nfEyngwKDNJ0b
G85E9Cm6jOh+JTFW6po/oGr19y3egAQO25Ps5NfHp4iL74IyaL1++5fVKlus8tSX
CdVR3D4+4tRwQX/8bne+AT54i4JXYpG7GFPZXk/0YtNDLkM2oNrKcSoUUw7ie5Z8
DV5E9MAyro3dv6VLd0rIX84Rtb7LtazTwxsREKMaxRbED35elx/S7Wx+5N0Nm28J
KEHqvQjJGuOyCSHvBLlNGN/955ZaxIsbE2AvmXM7kKRhfbAFZoMvKDMUVELtcsyX
yRq/ZKLQSkoVhemoDNw2iXMucY/3B2FnoBJ2L+GyH5f4wyGir/RGVFWJ0CrQmp/y
5pvS4TfgB1AyJ77niXK+Kmq6LRbWUBg2DWcolWxWL4WgTZNwvaZWwd0h8vUMvQmB
hnt/UUW8okVw4Auom6EU9QlahLehoW+2oETmXNmunAgZLzwA0cLwzQ8Psiw8Huhx
g4L0FKAp38Pmd7OxnCNsopwM4aJv4VTxWbIv4SzYQrApkxQUyed4SLZc+M5CrXAr
KueS+2yMz51CSfFSNZcyMkx/Okh89GPD5tCe3vu9OUf/NPa2JV8BNWh8GvGs2t83
SfOwiUyZtPgvjNrB5UNhlS1QmtYZJrSC9HemveaKLxSaIrDzWLUrOxg+Bg9P88Hs
XrO+BPQ+iBQrW0ZG70asmHQXVXpARgu/nbczD5cRd+ezH6A8ZmKDn7rvgK5vv36a
mJOEdxI/fenNI7XxSMC1I6aHBCMjo54bYJv+vnrtJRkCKdvcYxQRGYNEIvhbsL/r
U5SkEbW069bXxbnYZwpLSTgqcOrJOJEQUk7+zDcleY32AHg6VVqGHkiYg2l61FvS
E9BEZTSaoDutv+RPpBFeEFvDwtg5NMElhT6v4dc2pW2xOupaX8S1mxhNeQAYGqjf
aEYDoMZxbE6A5n2WGVXTVWDfrz6iwAK2TOeD2nQqrQ/IQePEd6pI+RkLm/ViwUjb
DJzhYKIEL5GOd9uLNX6I1J/XWOSHWsftS6FtJMWfbwUZpxJz03b56JNdv9lg01d1
5f9roMxp8fp/VW5Lp2U1HYqCp+trA1Ju8bXl9x6P8BDT99AeXW3U05z0jdfUnhLP
IwnGUJ8NoOYuK7aFfkKEPmEQKsJtu/e8e8ZmMHQyYmhfr4Lv35Y/41nix+L3KqqS
8Scoar+/74opwEGCNld0YXxMSMeaSTsghbsjC6HjfWbYPpjgcMGKISHOSgeDD0A6
teSb+7PToh4QztQ7xvZS8kRbV+lDQqTKlda+0YvgZROcHkVBRG7yvnnvz9jj90Sn
S3oqNOvg1CT4LubUIyJCTC4Zzr9ty5Rul19kOJlw4RjOy0VjY5MggXATQZUlsQqh
gFtQvCRHVmmgMKKaJT8/cidHl8+FLImw+BZyhKkX+ngjUR/cadce6bd7j5hTEQMP
0fHy8ZjI6IAYAkf45AaKXfK3UXzW7J901JgcD0oyQd9wZvjvXlaQ5mBpwTakEbap
Y6wJtGZgVBiGpGvmY5uryqqX7nhUVPJ02NejDRH1DWf725b/kId+c5GtYRw6nDtm
VkodocupuQunlqZfeFU4FnMwHdryCBGDZlwwNDapWC73PP/R82X13WY6nIDx3czA
zJp6+fhm9j0MFAFSiFvydlQbOamaPCTCnBR6gJMswEykcvTpAnLbAD92AP2DQvlE
SzY1h4CALb57KPyFORBMSo0Wf93/e9ZrwpbGmSTwwgfpoYMB4Tr3ecXcR9QN76Yg
tugrJh86dR/uDL3c3y10uwSCBDCZM5Tf/5fyjHVnR9VkZSSjsJRVUtMLaxPvm0Ld
XsaaKY2RFp3ZNwiAnenkbgEeRMo4Vq9jh4KfSioL1l3C6GJQRDruVghcSiQxPmIv
TKQG2EfoeR4NCiQDdY111Hb41XbLMXIxa7uKfdw2nOmPqbguYj4glUf8UR/e+hUb
vPZJAANu61D8yOCNd0w/G7iXYMYzT2YKU7Rs/h3C9HvVHqjV3wfSnDvyRmaj+l3b
BawFxHDWWZzF6jpPQVfrh82NHhfsyJHDB7PaLPyEVe0amDN5elX00vkkC4LYJhJN
wnB6beSwO8Q6mvBo5/2pFNbJi/T6f7O7O4UDKS+YOV2cBVubhSnRCBwnTlXH+rT1
uqrF49j45Et657Er7g0wBFjVtOL4VylLsYMgYGFKpVk4jn9hnAfqlW6PcTXOATSt
0OhzzjKWZkDH2Z6ED5yZqAGus/F2vZwSm8WrtQj62/Y6XmuOpgZLTotRIHHakVIh
O5Xo1/JIOQNxjiUkcStRD/wrmZMPa53q1VJftyCrju904bV3QrWTcWLRtZq0JOyp
y9lbQaH3ILtq/VYbZyjlaANPrMVV2JqHxbe5PsEg9FDukRRedjsTKZSoqxgLfdZf
RqVHYWNx8EnREtFOQ+dF+ndGlmNp8MnYPOgtWVyv3GSBJqb57DpP8CZaQpYKe6HS
pF2w6rjwsUhPwDLb+RqhSVSggRZQAYX/XqLncaIs1Xjo95k8FcrGyzHXkMf87IAK
9VtKnfmB8qaVgDE2Om6hOFVDPAdS/oPhvuoNNGkJ+RRw0ndn9sD4g9nu5u7353wl
aa+4zmmt2Wuxy8/AR1Pc7+XuWm0tNAHtQCpzrcVsL8lZbLaMG25S1EBQpuXO89wx
ODdasKLNjAmwlfMgu+2F/MRbe1Dijs+C1zDe8Jb/27u6vDgEZVKU3bp3nMRcTaFC
ZGhtteCeCne8hwFvb+mwAXD8GyQ60zg9iHmo9OcQ8qZNyt+DlgN5XuCGhZhBHR02
xFQ/VmUMMZoQUrmMFA1dPAmBh+/w/QOnsM5mWZ5iM3WU1l5vZ+/PcIKLlKmzanzp
GrTtkP94++g+pXMLIWhYoQub1A44ja9vQbYcohDAsiGASpTS8Pdm8F0TTkOo4gm2
eMYdnTXGTpPSeeSmTpkYrGECNKxzRW0B3p816ytPS4oEKQqe18CY+rQZ+8ZGeAh0
5Zbw4ulqkpe6/3HeNLuksTTIQFp8fDwz1LOqv9gl9Lu5dOniBA0IQ9GHS1pHOhng
h8qoNu4YDlzGRnsPnYV2igSr0Q3HRqVSFbOcYUqcfS6butsKeaKtlN5R9UiwN7Ki
dvJnCIrcYRXYCLiF9ULp89yc2hlWFztKSfcdr5021IgdNpgUCtlNTH01UNqyIpiZ
BiVygts0n7m9n3nb3tri35EG4QN3qVsstMqZYI6Mk9n0cBUAsP4oXlZD699u0tj/
qT9QKMWtI16rqdDiZKWwp1JCuj5uB8nNs7dWXYbxQ/YFJv0DujnoWLjnE1n5HRKV
DHFWJll6fltrVmKpMZuGDx641M5o+UrwRxallank+M513I71B7QxNcDsVgoYarrC
4NGMCoYSkNOULMTcymtnw62MeLsjY5kk2xw1SwD3KqmF401fCJ4LykOT8nR5r9dG
oTJQ9G8jy3qLiYujLXzxwdGZJl7cKd61ybb2t33ilwxRPTdrh+wuTrTiJLiTPkFs
pTiY8y9jzK+9IXRKTIkAbqUhRZhgu2BLu3t5Mz4BW3ZFTNVce0L1h+J8asSAHdz+
3XT8lhQhUhUJRvHE4H4r/CHbrdSugPqc6topmFfTeHALyDROpAyEtP1pvTrSv2g2
/vg8s594U05Fmcb+X9yZDVbJr8pSAqAiWkYLGZTSYee97cltMecos2lNZGWXQukj
xRCSMacBjibUTanC+kY6AXaNj4IXXO3KKZftewreeSKuc7FTS3T1wBujvRH4fTct
RsF17L/mzn0fodBEeec6vMozNRtRtSmIwPkH655BKTKbPp5OOMotgAnEifK0OMY5
9mHgP8KI3rJHwB9RDXHH9H/Z0CredO0Ss+SqqlUNyHiNcwA2ULHhIukxzdQMYY3g
QBzqUJMHbMlcWMoRjLgSaR5eNM5EG6MFTvqP0LnRNj0j4H7gMX5gZ4aXdegSzvVY
126iw2XOFWDVWXHwlYTbeTUbiyINNUd9+BPWae2iH6pxI6TkeVPOdIRY+Y/xtEFX
JBIsr7nlpY/Vs2m7+cwzX+zg8sF9hf4ZSWH9H/81QI22vbMYpaGpuXe9BR4mOiYF
GlsMv183fvMP0AMhuQpVLKVI0u9eQ5q26OMR18tqUc/SXjUo53zPfcdBlZgpzTx7
bRewvvn13XwmAy7rFFSCtvU38XSmvEgAtkjxkd6zHHc2gQGsccdejTqPHYUPe1rJ
3ewWoC8qof8OcoLXw6fb+dqC5qI3flUvcIQiJUqI/t0bgRZ4wDkuaBJLJEHTBmyA
kVRKnMODx/mkazp0IFhHI0fUxPZtcjgr6lvuvQek+P0dtkQTCYubTjqgfX3pKB0c
zEHD4mmqDhIF4G++EnZpVTDv7V/PGEA4Pi8vvec0LIwb+PubwasS0LxGnFl5iPzF
6/nAoW4G1FWv7//BbOPBOxaj6yjxTglafdZjGylpOH3EfKt1PlMFqHNsk4PWYpKR
vNgwZj3euosJAh3r7iYJ5GVPiKfWpxytuwDiQG/6GpEpJRMfphwrHePMfcY6DYWn
QJ2iOEMKTCht/K5tL7ebRfcaKC2ogW2ztdJbUN9Ewc/RctTmM3HxcmJJq42eWOOX
8LU8Du2V7Ri6bqrr7Li1VjedVpZe2mI507YTUrQNp0oOuGxtZpNO2qIIuVu55lGK
7rJM4MqFBzqpy5EXktFtDy3fDN4YpKNWHjtVURU4Alm/z1vQUnBItWBuOvFXp5Ml
1hwExODHCgYX/3MuOY/GaI/Ail11i3wSLjBsw/J14z15xPK/Vzwb1lxu+YXqf/qc
bVSTmq6Ylkb2C3LD4CUuDetr/X03U7gLZzPyiNC0hd/b4h9P9VWF6m8K1nemzNix
GSE52dc97YVQXLtXRSY4cC6SPFgitrz/9y6Gn1tD9iVopsMuyE0oRRwTL2lNo8eW
KCoIhRRpkdaDSSI6Cq4mzy1Cso51Q1iEuBfli4k4lykDrFaoSeBKMLNEnMWuvHYk
aYZkptOQUikszL23X3X3xxfLHzOekWyAALE31NfUVN+7E/GMTr3O7gQetCU5G+PJ
uArixhYmJ3//u/KpEWdyVaQA1tKzDGznxaZbQov7YSTQRAqufSf9gsQB+h/EwJ6Q
lrKYPlVQvQQ2PicKtJ0W9BUlU/SKmFTohQsX6vH3RY6Tc/WGVFdyazHvx+8LmdMY
annQukV/9HHnAH1Y6h4bR+xEc8wn/Tin7djp/9qzF4S61HrWUJOAGZtObEcZBYhq
UT5Rnrf1Wgdrx/gfrkod0sSzF9KWhTQhg5jSz8am6f4ejrlI6xYEFp10D9q7xE5b
RoBYbc7RDteanhAYm83w6b5nAvNnLJIFR0pgm0brLCejA9gxPebIF3TtUrqSTpvR
ZoIAKGpc1XDLKfpxDhn68XMFiT8ZCQqJ2i+b4aZef66CtqbkKfL/A62v7KlpznbU
SGvulvNbOee4ds1022BZDIm9Mv3+eUePBi2O58/lUB02b3vDvRTfp8T+qlG+xPN4
IOr5kzQMfqfai1x12sAYG55ULxVYFcwobwwpVJJD/Vpk+rh6cQ/wBqXl0dnlY+h6
rUEC0TlS9M/LT8be1BOyJsdWQo6Z2lvka/pcTRBHTCkyL/y8PakrE48qIwS1i4iX
+nOeVdma5T94WVM5vbBz4k5U9Xz6/6zf0yk5yryEbCJBkPekwa3bHQ2Yve0WOX3q
C+wrAYE5WKaxzKWIdqe90TOdIvOwANas9fkFmPWNuK9TqulgybquboEUZUsnIBaF
4cNmcTnIVoeR6hZA3H/l1wtH8sNdBoeOSCbviQDsmXrzWpwG4Po5wW3kP1ydh9go
iCN8Nu/V26X+5vabOxJ2YcePm1udV6f9aFbi8yNU5dKfSzeYYq3pY2+KD8WPn4uK
o0a/G4BwwO6Z4TqFFnfpS4lbl/P6YYVNuxa77h/dhOU36vuWAcBMBeq3E3Sm/G1G
B9S1yeJ/AB4LSXvUnaFFnSIh4hPgwp3YXXbvhnmAMNiY6E32jPpEQhS4MrGCYF8K
snq2yOpGM+uwoSyQ5a7gnN0Yyu5Y7gt1QntucBt6ANeIwyxz8uBPYl0Ltlqf+nzH
2BRNl/O3IPlnDT3pqyWaJKsnccBgba0N8bCYvur/P1ydf8QrhS4+Fb+wKeGB14Ov
H/6jWw8KlBpSpQjPPziE0CcxAKqVTJewNa+jVLqgqnesbHKtsXgr1dCpgwKHIkvU
DNWaltklFg/4z52Ihx8Y46U7D9L4u5aQAia+D5eK/WIiNfQBXNW6ztVWCA+XBaal
xBBRUtz6j/UnaZ0uHVxgGU3anPlDFKRNwGV44tOfOoAzLR79VIdRK940wnumnjFY
T/ZO8Q8kv5Tqnmsuc/3TUr4wG0pvnJsgYm3H0qyGgDFI2OiUutfSVXpJVz4/PBOs
em6q6zfsNMwPZprZkb8583klOhVMLX3+gcOnBslrqTdQhBL/LfV33bQRJ32yFHWA
grtyZHMuQTskYxGFZll5dmW3ueab2GQEeiDm95nSPNsD/YT9/plgrtX4ppAVXWbF
/i6MHbiESvRiO5B/znQvWCdtiSHUpGeP1oV3kJCVKrBmMvNLNJratlv7rLz7S5JH
oopZ2S493IitAhNCJn6yq5egnmjLj7yEQW96KQsuBOkMncruzsTaYK/Qt4cG37JC
0GnoZCVbpuoGsv67aqdSXTMW2QOk8YXVlELFsJutmA63vFTdlfZigBlFXdL1nXxT
5GZz8VqZW7KIKYARChzY5bXVFG9x+b1tlz8gLuYP2dfCCYikKeUbwe09VWU/lWb0
5kunyBLO1CmA9yqejl4J3T/GaXC1Mq8iATAzvmD4NssprfA9+fDe+CLoKIyLtjhi
pf0uOyi6skhYVXADaWjccFKRfAbiiDNQI4mM2NTSCDpYp4gYKzHqV9yJR1L2zc4D
DF0dxl19HFXxONvs1eFsno6FtonHXHpzZBblqYGoV3kQhBQBdyUkCT1bjWLi4A+5
LAEX/C/y4SCluGMx7fMK/TLaDmNgBf90TShLK0paaAijKy2YBohL8eSu2/GPR0jH
OYawUTmfAI8Zr3QTVMs2SUEuCqsUkFMYKjCfRokD/TpgYLMmnW3dNG2jFM0u3Vrq
doO/XY0dllDzNrixBZWKV0jqEx9cGt6eQqglrbAF6VxmHFyigLeezuIEOQaMt9Rv
MxQx3CNqt4EsB1L9Ji1FQ6WDMnmBQIgTIKRGoc+pSnQ2OfPsz9PHilSxrH31M09b
Huuchqyot4N3PAzR3CDseT0LSCX7n2KI2yUTiPm0tdOOHhDsv42NkMB4kZKHwC3E
uLetRj1Z29nHSMz9G6wWYjFfgUc9IFMJGg8OLH9rMekL9+OizSBxnXYGd+enE0wQ
u7RxXcQKmAwqMe1ZL4RcJ9ufOMCo/zWZdQ3JYEN3mntdOIR6OPi+j2PpnywP08OM
bZXeFD2KLg77M8Jwmubar1mPRC5xUOIPmMD/eWqM3jInm0RhELdF4FZSghf/yQtZ
MG8Jiid/TXce3Er0BiLCuwMdYqzp0hJ7gRIkzup9FiSWSvYWv0VCvsubD1tCwZGR
gSoOggjzLQnp+GDC77/fOBfk/EsPqrBC2clfr3fbhp7iN3olc7mUbbtYCtoScQJU
j3lHVadFysdix4BxGojKNw7pKMN29MISreRkUdD5y0PoANOrKEc44C4GgzBCpXBS
+CaGveb9kot9wwwCWx+vzCioPLEISL21uzJQSldv4ggurr+1YjUM6lfmPAtAVpXz
5SMVPDhB915uejIWyfWk8vCXI54odyQ/ulJjEgpAWqZK2u4tMplfToM1nxt3PJ6F
lg5XoUheGMPOMQsnwJx3rKPWl/EIfDrba5Y035xjZZPBjbfXZ18SL/mVvVR5qgF8
bFQ3rQUWTiz+Keqv1AMn70PGwDLO0o2hHgpWIQP4eHhhRSCemExdaNbaHD7rVovd
UsTlsrv43F57AeR5UEQxw3yZSM5JVu/6Sa6Zp5nGBLV30lK5mRl6Ac/Yi6TENY/d
/vYq2CIB6abNUxSD6Ww1OUXi2ilLRvvQfknn8RqodFlsffAPHBx+X9rp35sI5I++
Avnr4mJkAHWz29XKi2LrdsWMJd1kekw4G6kKBcK07JIfBqbTwdIp7YmiBhhgGgAz
l7w6oTPxrqn4J1GqMbonYg5WM3Lks+/gegTTfc+wNGSJLsla8L4kzX61+D1uFPZH
Erj+uCnKDy586Qv6KLxQROHbNbs6no2aFfDaRKgkR6p0DmeD1Kg8U1v5F76pMiHj
mq+l2UW2dQ7efQIgNfw2ul9/RIJc7NrtW65qDuG5zqh0nR9qrbdefMhgCeiyZeZR
HwGgaotIYTC794+441La3oSAOCJ7+3KblwRzO/YGWdTO35BJC6YGdFaur91qQFKY
YxteU9OaxDVmr2PpUldc9veQ3cjZmZIgPIJu+aMql2FztLIqRSEsR/YMzmEl89wh
tvFneJwtTYXZK6M35U2SnY6z76Hf0GSHe2TEHSNawFjfVaF71r3QSfKoCI91XV6s
LUsOEUMeJvL9Zx2mdw0cVwBDjmfP/maX1Ckk1KZdalW/iCeJ3XgZiHeAVlfFRhXi
zhOgTa3UhXcWlhXg1FJD/MnqjiBSBLyVG4UkeKQNrRi4Y8fcnMREQs3ocH0nRfKc
jk9eRcCaZQhkolwKb1q69JAQLKdPpqt6qERI0SRj4ekT0wN2YKmFkCUNjuKRMu2N
OjwZWE9vzK+/6kVLYUK+uqUXy4AN9kqc9bQpHVmX7oIGFeMXdpLyqB0LG3two4dQ
5Mx7ArN9HN0l8JkPIvG8qUw6fnaj0/AyYewSIu6RkrM+poCiRQANii8RC48abkc4
LBIas5bXm9ivZ1VrpGvMdzmOdW2aUhGZnnNupQb0MIpQYM/siQqpLsVyVOw88VBj
5d1j8YK8L0ltAA3STSAnAT/CW2drl2NtjuLzJqUxbipPK7M73QcJ9qxgobVNLOrZ
fVv5qLflcxcDbLGFEZ1wRcvAF4xYW3ns/E6RdVjYHxhXMals1ebGLs4nmU2cQAnJ
bQ2qL82hd0ScLFtpKF86Sss7NKf7PO+ZPamHQ+aPwqn5DIXVDw1ij0m72nizsKEC
vBL4solWqcxV1BS5hRNZo6gL07ov0fa61JPoHIj2CcW+e6WxIMbZkl8zaM7SLask
qF66ZpX63p8FoqJV39TH4gEF0U/IJPpxMI7aun7A51iOQied/txjHFCMn56YJAR/
OIpHgBnKwW0pMLOc7Suvu7AU4TnskBj9VY+wFi00sGbKcMhfYQGnah0z1bssRy+I
6ygT19yQMEF6I+dG7q2MBDhnEgvkQqNh55SFb1UqILQgK8f0nJV2pZDSQMvlqzyf
eUElOI/yHNdVEEaK3cvPEVRWfIWP05/aSgBAo5HLZam4u1eDn2W9nzIpSwwGzeeB
6d0srVIlKzpGrA6tnNFf4lNtqyz9eyVn0jBTc3Ofghlbxg+2SUO7ozeYe545lerq
Xw64d5vA++1CJbpYEh+M4G9rtAEgy2/r5sCttjlTTxpCcGMOtul6vLpCTVozP0iN
AUfV2tLeFbzL+InLVYf24KY+avJqMksEPmGR4grLdH8rN42/VvMePYOcIV70RPNK
5o6v7zAasAbf07RhwlWyrCcKPwWh7bxcIgVK4WYfeOa39GvLsb8QDYidaleQ3KeN
mhf0TKG9cZta/1b2uXx7rI8E85fEwQHs2DTRsOSAX5LZVg2qsHTO1GMZz946TbGK
SvDKPrb7BNS4TagRG8dJxOOkl7teqxwxa8mP7md5uuRD6WLxGxr1vLw+Nmgeogy+
oUdZl3LMUumibk1P2Hen+sTRB6CDHKKih06lQF7P9rtLCC8poRCjIKFi59jRKbc4
YLEB+dQZB4lKjhqqRSG5Fsdek0jFSsqEkDIViNu8B1yM33DoMCI9SJSBgxkzj8El
qpQgkrU6ufhudbX9cICBanU1uDtM0ZA4IJ/1X2XHO6wnkmfTYQQWZqeP+TrHNpCb
+suvZYCyVMKNTZzPjk03oUWyzIYLePxkuC6BWiklkqBDaRHcP1A1o31l+gGxb/8H
GBZ32FSu4DN59037rkyQ/zO3hSlrZqYt3VesLXFko/Fqd2hImYDqDIty5JVWLbYJ
KVP0PYsM5Sq+s3s1ZL2Y2PGPyrPK/tScxQFrxbcv8vgKFV59gJNBKQDAln0mgzgT
YasEn4kMRk8IFwwQEpVeuT5amtibIYYTOCYzua8gE3hvKu2DWkjYu8GfKTIwrCnJ
MpsYoJQR9SS+Tew6o/0O3y8OgYusRoiFat1wU5XJdXpGY3iFB5kQj6hiAaRHz0R6
pU/0Itpr0Cw4ML75bhKUUxgLzwj09ue5jiGi8TdtDQ+2t5excVhNJqcZ7isT5JRf
leQmZYl3Z2CRHpB6oM8/o59Vbng4kvCQ20ZD6PHLWmxSVslIIvJACWQceXxkCZCs
TJYS51o3DxHtGDTq3I9lOwWpNjoqGkmobWf5M9bpuOeFzWpeJObJg+UzN/59fdpe
RNMuo6yPuWHwck6gchxzDj/mDheieto4MRoTOO1FeT4SN7PT92FZ3QM1PHl4lnKc
VxyD1qO4Tdp7jODJxs4ZIsY5k/cO+YGUlrUvUBn4fmTgSY1ZSszcaAydDUAd+/qb
Bk4fdIEOdBQQJVTmOniVAN0I1lBgOQ6qPFCnVhX4IZ+akQa4/TJaVOjii2ZqYcqr
RDUDhmmcHDFX5uYV8T6XbqI5yM3AEZNNUgPJpmbwt8cGQx+6t1Dt9S6M8KhWZuWU
TvfDdnMWDcPcFF4GA5k9E98OpXAgEltjl1lbcTsVgB0FEee0c68LRqO/zvbEYoxG
GF7QBFEEepOaigSzF0WAFmgL4ZH3pSJk2jwygKivTL0bqT3XogUZv3To/ucB7wdk
+cp64TP6xzsjYuWYYiSHxqXt61k9sPzZkkoiZwtne6gJhWj/eQPs3rfCWW/Ivmz7
dX1MXZM7sPzNRTIotFOjeFOshhue8BHe8lUnuIH54bwceKQwPSKdcS2nFdx8bza5
TmNoDWvdSbGmQxNXcKCPrKD2Q3yEROWMkk58JVHc++F9iXLAVqPwBq+2dA16Bk6U
lBoemuNTulEuDaUcznmjqVogrdkavtcazs6U1ROGAnkV5m+lMZCDkaSL9Wi7PZpP
86ArayBK74s5Vum/t1saP7bFmWzBAU+oAuoex44PoEKGINVFowOgg5Ry9t4vOnD7
T6/T3osZBdU6e9poEc6V5pgyp6wCiqk6fmI1ure5MZZNE4Se7QepkH2+ZoMSoNoI
ZKYFQrnbAf/quLeD3i0BBMrfCOY0HmVh2yqgwto2rLSNusgogjgBUN9v4DVfIUmA
nz5QpP7BqUZ0UuW3ptOSi7TlOek0JPmcp+HAehkSwpM/vhz5EQwa8opvbrRrneR9
yPu4+HnrbCs8iGvGbr1aHgZ4sTbnxusvrH8EVVUDfgPRn+xA/t8EO0Ro1FD7ZZRg
g8r90iwCDht4DQHAbnfTgE97Kd74F+Y6aGoa4DfWRXUudS/ZJ5WHM9YstBSk4x+s
IY3zUKpKUzFOjlbzIx7eq0qeuec0czcvTrqVH4TJRVecXfzFxUhiYyvly0KZULrf
633xoGueD59gVr4MSzcHnpP/5vlXKA2rywx5cfVEacT4mwCEZFviw1H5+hwJTVeL
vQnkY4g4+1dkvl/qRRiMU8+fwRjdaRv6l+titl6euAzcBd8Tlt1vZt3exojTY1mO
zQOJ+NDQm0yKtgSeFNQCVz8pP5kqRwiOXcPyqzVTol4nvJAOHu+iGDpe3EG10Vy7
NBc9/He6epTvYDTVBRUGYlKqmfEVkCufnh/zETszz6rist6t78N0jlJnXT6euMif
PxmJI0YGEo9MGlhvxIea2DgYqxaRS1o7UtGS5ewhnDpgZHDzakHnx4NOeyOExAHn
zssoWRhIOhBVpEI0HN+Y0MXOXUhB1H6OgUxv5EgzyUEVD6KNAKZKuMIBzQidiAS0
K/usxFU0HzE3kTWZ2o6++yE1tZobIIlxhlH2IKSF16M4Cv7sy+b9KeRpR9vskFEF
mVEGKBefwzFQ4tnPbNrNkXygOMZBH/0H0pK7Et/QfmSClLcZbSOggZh+oMMIP1YM
6vxOeCoVod93x1KwNFrOykBZwQopzdbFxfy5yvJj4H4deYktXVQfMDNg5aj5ocU0
Hy4iaK+DpsuWkgwCmhVwrZ3XBmb/CX3OZGPVF/mpU7mgspnBt0zWKEshHv+8zM/u
P22sbLRWmss9jct/NIwOMj5gnwdOR3CL8wDytC0CAUZEM38S3rhiphJ7cqBzXL3t
4NhGWEtOVTgYSTdYl7tCQsxjqan+OwpxUbd1o+WMOM+A/b+bbGtaTRgZh6aC2gR9
TZoLEaMRzb3XyvuTR+MyICmLp8AFyW8LJkfjfHRdksPDLNZOOIbFjXGxIRJrccQ9
kDj5WMWMF2E5dz8aZ6J9Jt9j5UAzyBbU7fFGF2VGDz8rQTvqvHCXzzgbC52fJCgF
5Ia7pym3/eN8ESWRtYASyJARHheqwq3DB1zgkWIOlPSuU4JzlwEk3wZnzMO4VeD4
2vis+Z9L8S6XBYHvaptuU/kdW/x1K18dfc60Kn7+qynNuAuIbqXnVX3wFPEv2Uf1
Tq7ICJRhF2UbT0xtyYJS5RcI5LHSLGnhgeGGqu9hEUmhLSX7Yd0xn4m53gvUx+Mf
o/hWad8Xu26zezIkmEPiYhNCY6pa+/Mwyt37xyWQoHGbdYPQk5bq8l9h6goWNs8r
dXmh3FTxd0Mkd/aUcc56nSdWOSOeej4SDDn1hc+q+GnR0bX/SLrT0vaxp6EvYVfV
svZpxUAkHdOkbzZwWhcSBdPecrdCnOv+CfOzP8BMdeLYGWRRGg4U9Ys215MfccGg
xjZOaJoIjuZ42IzK6IEzbXEjfKRD0WVVyPfSxX8Ry21zE61mj0ePO6d61zYeA1py
8ew5515+cRQOXxNde2vSGw1PiIeRAQCn/IA/prC/va5RMQL5KYaJnz+E6Xx1BB7M
W+hGiNTe8zn35i/VyEs7JfzeXsd3JmZBzt+QLa9sESCh0jtPm3f/RIZg4yvZVWBH
UcaU13CsClc3JHQl1bjoUfhipwKhTxz7wqTOyleg76ai7yHwyKkDgBCrsgHxGj5B
8mq4Xt31lzPmw9mT2Z4J23Wr//Ol7yyD/Qv2Xd9y2e6hvep0AHxKs9pdmuWFQIsg
UZBDmbwf00UeC0xMleBXspSM1hdDK3bThN6x5ad96P6AhN0XEzgpXJ9cB3ZQGkup
mxWq7flcKEVi7ViQiYbxnPPt8IDC50S8HUWOydsp33PwUK+og9imuK/pUI8ifIEf
sJgUEAFMx3dumWoSCql85oXzxxXQtV5UgtmbnjGEPQwDBnt0hEOTpLQ1FEJ8AmUr
AQFxFyfYW/F6sTwTnf7jokf0zfFqGMBO0FehVsul7HyNJtjzoZDJEQgtVl/6mmyr
2Kc3Br/W7vy8yWAq4hO6Lu61SNxyHM7fY+bVoapG0AMThT1Wy4G6XfGFWf9lRD6m
w0WltaCubk12GxJJ1qJFoQBhd7yiApxPvzeC24flzihJWHJSWuoY6q9LNSFsE/hG
DuPv270itw6cw0GzuJeRuBPWXrIUJB5KVRRt1Ga4xERan+T8zz2aXs9MBG5pAbLo
03Mg8356jjtva5lLaAypiQmhHQrHFKvtnWkYnPItY4dZsRYDRfy3hT1HDmaEn5TU
5iQtxtPPCVpYsfgXiYTC4c086yQI4PVl9IMvHJMqaxHURHJSAI6avmGRUGyncBiv
wsf9+S7zjFoyl3mwEhanH93yinUCF6QjUPZTz8h7/43eZksn0NOy6ZVuc+BtW/Dm
NdK400wniUMgYF27P+2BG9gomo0djXO88Xl19PLVePaaeHj4lz6Ivj2eEWqLmpqM
s9nVFN9Bo7RJ3/+ZsEvx6ReVXWJK9E4C8uL2yaZ0P91uIrU902CDzD6m8F/XrNhQ
0wizP8PZWflVGrwUpCWtXjQvDAbDcT3Do4fipHAOkeULpbG1CQnH6H8zVpGpYPHH
5Xxf+gygJnJNUSsSIPG46O5wG4VHNV1NNFsuzlXtFSoVpqHY0N1FLkUBeuWXOGUQ
46soOumJPZDyRra3xUUExphsCvcvD01p57RY+Lb2YD5oq8qiKLxevKqKKTvRPY4q
73WWly/LNl2mD3uJf+TXOP1Qv7u3GnE0lvk4or2plsbj3OmgH1WpG8X0OAvo4VSS
RdGZ5e0VzghdyEKxiWM8kE0rj++ZMEiAErS4mmj3AB05Qb9+RRlGw1rQVNoU708C
zJ+SYM7GVyLi9e5zqphvMuBdEA9MNYI1rNahlQCN4zsELKNmj7pxGxqrmITXbpz5
MEaij4L00ZEGbKThht1waX2xiz1jOwf80PjELMGPCYzEa6KRrnmRp+JVt/M6C7Gm
smd5ztcPhBdwAGzbYfWtFMODBX/6KtL4Bqu6FAJskE2Ar5iu+cfegk0veJZlf31s
fK0GVhc4wQdAtdYK/8JBD2fOvdn9SIytnECM3EbJZB9Tyrzftk2mnDSKfShgso47
Rmlef41zDf2VgFxfB799j9nI6FcQ0zqfPdZcRnF6XfPl+mxwWBLBNefIYEtqMvQD
GfKj8TAWVNRqsPpKB6LT0alx+KhtKiEgJNA3GU+Llcfo6+5957nY5hq97w7CwbNk
/12BjYnc7GLA81eG4FDvgyvm0YTRKrTtIVc5W6aAQyE854J36+ipgUMv2IA+oVy5
7jSn9woTheDows5NvcqpJX5PYGokRpEgxGnXQvgXFSSaJonbD3WWBk0wqjBotvSQ
G2Hfxdwqy/00Fq/IeOrRfnAzesK4ckt3tZJRc/MWrfIUUUq7YpI5pu0Pe+zdcraI
YKmcyMc5BGEkxG1GxJ4WJbZxkkr7yyCe2i+PHtbrVB6+oel3UNm0TRVmmsoCfZ79
2bq/d5HLIFGfb+uuI9n+vnd46K9vq4xEPneNe+ugaP1P9sJxTTIZJ4nLyc6h5mPr
mWABKyI3wq+AonZ8lgUkUld8xOFca9h1NsiS98rVmWzXMzXltk4wFlI3D9ynZ3tm
/qg3neCLC1+l2aCYlRd2gpN23mF3KrYHslmTGjw6VhqVlXybcUtaNyjkT/vebZXL
4q1DppdcEDDmPK9CFXKVwLgVpeZOExCbrB0QTTXdijQZ3uO6p/3KUcPzNmkQauC/
Cjb9UIR4+r6E91infFUN3Brt3qoSp43vmXCd6DlQZ2g50Z64uTeovw1n63qenQ0i
l4LeeQYVbSbNZIICl1ih1xi2K4YVMbGzqTCAMrKxEzHVu8Pdh65xuK68M0ir6iOO
l7ROi1TaFVMUgABNZZMYRUOl/6lW5efDoWEnTVoOwHObuH9xf6StTY8UWgKqWpM5
+5Ga+dpb9UuZdIkbVvJnQ2LUHpoBz26nIZENWqwPfh2/TP70To8nZBLTuf0gODI+
WA0KOEg2NT/SDuY/9gTnvlpm883oNvuIG2v5ZYANe9T7BH2NSepwt3XTWz6lu4OE
QSC3QnWB3lbOTZ/rma1XGY0DuINF79aA8ViUeOq5L0TkgWHnmPCL+V66vtTF1AzX
ODi6AE7vs9QKq5FGKSZVAUhJjqz6pi8x2sQQSgOe2qfTb/xflNsJ3bIbsDmssNCF
bu+b0YU9wzDVqJz+jcLEiZLfK0AYdoOTcBU2pjFsEWjB2J4JRWFxQzERJuNL8RD3
KA6Aim9/r7LGMhpnkQE7fJdUyM0QMb2SlSHGWY1h6F6xWA5FclNlCZfaB6XZH3sn
MUJ6R2LtB2gZj/XkGRaQHjcX4s34v4xN3wJVvCUAmJXHkPM/n4rCLcj/WEODSKP3
APM3r3HfetXRY3a21g6C8unbo8GInMbCrSAuncQvHadyGdEMPHOEiE1PCGmakJ/p
Wh5xj2RMlmfGalJbjzb2lbTdm/V5fovHP47Ac3BpFlry10AzM07GLbUqPn3WrpFj
WyoTC2fVRbJz59CawtjmCdOyuC++lzujsx1qTUDNOu6xl2DmHPkZOCYvjVOWte/w
b8AzYuJdAiHpuqexadkHEROc7YUsK3yzgYPA86CUL4MULteZqfIJ1isHn8HtvWMB
JGJnUbUH/lsTyRsQHXW3KEuN71Ku2W5ZX2c/NoTcI2AsvsZCaP0Iu/3vb4+IW6z9
fiFckukoIVfscgmKfAjuNUgVNh+frMdjYFQBN8vtmbhiWanZC0I1PyigJcGlcS7x
U3eaIbdKH5SCoNE1nR6LQKTkr1E0DT9N17zHQ+tqDpnciKghy89OSgM9vs3uk1uS
5+fzgOc3lC/kNpL+Q6pJm4QrbSSzfc65e1KzD3R6pZHt9z98SpfPV4SmT763gHft
2DKCN8QT3loqXaJyOb6PyVMdwlJkeGEbQ6Li3xb9UUR1IX9QwGxfKz8GKxVAEhla
1thTvoBrTwxjK231JUWnZYs1NCYMXplps73JIN5BAygy/CYMdeezP5F0B3Yz5ah3
6XXdEzuQTOziTuLvScdczGf2+w7D1hSsBtmNdp2CPi8hOqGwTxOKU2UGLbUsPV+7
NGrE2MTRy359/RGQC1u0iUq22BKNgumkk1gJJJ77hwxeaKz56akP8EfVq65iAAYb
7a0nbQ8VjCCn0yefGe99otUEBuxSPkSZsjs+qf6AYH2SLb/7vsFp4fGz95+EVJK2
65Uvnf7Kd1ukt0ytn1rAGCmVPtW2dZCVLPfEm656pc6pAc+WzVt7BB8fH8Jpf787
xlAUAS2Bc/0APuyjM46qhZIDgtel1WUthGpbkNT4BUovo1ifdE83m8dnIpwSfN8X
yJhZkgmLUoViUyza5m5q5LHYQJI8ToMF7G8WxsuD8c1FiSH54sBzqwJ0Krq1wraG
ByMw+S+QQpEi26SlDRI+5x+I+lpTGA32X6BknV7r/BuyWifRY+L+cVL2MLES4isK
NMqLTLEc8lqaJLaEmXXZ2CZbUhkgESnSxj+0Bu/8j4vd6wQufOeoHbM18k+mJ9HY
3q8wfFpWNBc/IV1u9G4S3J1cRJLm7LFzken7pdM+evTviN7n6Of1/TniQca7bKTo
E9/87O7mI0ScBKkmf9ITd0x6MiyIK+KRV0YeBVrfB3IzOkkeMoaENNudv9tzPHSa
ucLnoJSkPdyqOLQGObyBoG+L5fNEqxCz3ks8ENznR7BhEAjvC3CGQNkfugMYMB7Y
QTUBZV9YIV1Av4KiDyxRyABnPtaAKwXvjC2pJef4Pf3boepKdTDS3EIhPaY2KRk5
KTkrq30CtqzyYWsd3ISyg6dxwIS5s2SXv4vbmoWj0/OfOe1oqRW6QF7Z13Sz+ag1
W3MIuwgVv88+7/GW58AkfjL6lsGG9W3otp1RnzP0StRBZFZkFCgA2r/UifSxYTUR
/0yn/1cmn8gZAU418sFkdIMWj3o/ggBrbHyu5Zetaghxc5cuYkcXpqT9/suMEnFH
TEhYAtBWdyRHdYFTOgCJii9a9tg6tqm7Rg6Pw2UruccIzEt2nqo1HoQ85Zq4+zcS
sI9pf0cPrCR6NZ75fJQ4cr37zewdNHV2FdDEepn7kKZ3j1P/NvDIeKfm4JdYFLvn
TgMw4yZUrWsFVEBlc+t40/mMzWQrt4oOacomx4XCJLpJBSLpPDWe4HjdYOf76x6A
tWGFW231SyiJ1K/1poerFO4MV6sObrjRTooOxWQGIsE+ShP1V9jDEOSs+2/e+KAN
rq7iCr+LaizLD+RI54zGD0VSzMs6A5pK6isNxPh4bdrGLHDZBFWu2DfWSIIsYVLf
XZQMeByYWob9MFCYqTGeGx9WqTqJJjT2bg+e60kVn74XpfnqvgmNZ9zKBpWFZyIM
z48BEIvgS4wDPT1R4VzrLKQ/UDhCpncqbc4n0zG2jh4AQuUsNolQgrBt1dJROoY2
T6EHAqqosUED60FUtshpynPVx6rzdBZCxnwMCs2Lrhq+arxVaSsmZy2/tHf/OV3R
5Q5CvPD/Dh11ayWBPWYyUWrCp1WLHkCFv0PBnELoIjVERT7g9FDcGX03RZE/OMG2
rRtK+NnsXpibtMcP8zk+idqRxsCFJnznN6/EytwwfQ1+oC3DE3WaRMH9kHaFsJvq
/Iv3Ba3Zua6tzdC87mjVuvx0hm1TbN0atZtUoIkXxtiHOaSGZL/djBFnrY/covMv
BvnX8etnqVaFijIaf0wd2IUgz7LTlyi2O7HVHe7K9tcgpkaoLkY+aU0UkxtuiTCz
xUWrSihGXNTIcqfasuYfVKAMOHl4i/kczcX/Akh+57YLNhwLbvc50yft4Okt3T/9
UVtcs3Pn5qfmwc1L3u0dJXu90GNUxNuwbGpk010sf6mnYWNfPuRmuuTmd5Tue2gB
//RTKB/RT8us/mpicRSgJX8u1Hya04fyxOv1NWlQTUffWzyfeCn4gEGwIIe0VOpP
2ttMfwEHzhz/bQUgJK+MNF0BVsm3R/4lJvwYX8f3tGDlXi1OWJugNVd5XQzEl3pY
tsFBh0+NpWQYgEcnM8RjXmU94Kj7giwLGeECpKgsEISEusPpjHQa0TI35HEAz0ii
KYL7xUO8c+pYNXj42Rz/n+kG8APKcxSacWa9hXO6u7iJy9R8QkGQ1prJHxKuRANl
4Bw2RBN140rWJesxOHVxYZoXP+TAWFItr7hl23CRYTkMtKB7dbfZHmJ5pAqvJNkN
qD0IglRFLzr9558uVgSWmpOeZW4VH4cplkq85cJJZt/7qJRc9qhLt7HriY/gCTbI
By8Aq02iNui9DL0i1w+P8KoV5B8Q61NQB/iXu114eIumqhsVarPoJWBoyTEGHii3
HA/ccdZKyJThbATT/vM0T7tQrsG1CKf0oQ/10i1S/uhoIaJJxpjuyjMLP45qoBNC
xXwscxjNodUSxRo5N+HLJ5sYFw8X6qmP8f5PjI+b6H5arDnyNjVhM0kXnAc5Waaw
Zt0bbVYlVk0ErvjiQA2OMe4yzFbZoRK1kpXF7+Xme+riEF9VUFl97h2sHM98ar4V
GOnNvkLoCk/1eP4Vd1JXD88toywpzGnRePfCwk8/BcEGNMHTLpjQIgQyw2GNp1qT
iTHk2dx3zO6B1imC5T2EXBt72//3AAe3MXLV3QB3M73HPuX7rDGfLaTzBZqabF2v
FAmDCxZP8VC9iZR78Ay6stSKKDqismUrkNvjY/XHZeuTIZUuRQD7amZJNOgruoKH
Z+5xeFlbMY/9SmfJEL35C0rlLlWi5kB1VxR+pwLeoa8iM2SiLhzxTwqOXOitf0Wz
71N9YraBZx1fFgHER+PWaEDOx9ruBxMlj1HGEeTmumIoiu8NwsGqGvSn6+1b3DkY
4uKMlxOkfq6O3naZIdByklmd/RnKrlO7/U4lombauAj0MKxjqJPARxnT3pT4bkYB
eEnqoxYvJU8mzaUOKv82a5kuYiwnbYgysuQ4TPsf28HQPW+9c22tS6UJLEigsyPB
QmGcFbKfo+ItCH5WitOLPO07uL4nCfeD8dS0k6BwGFVRqxftRZwJAknpzNqmUkdI
bRIjbX0xPioQ+dl2K20rb9UkUK9dpl79kT5s2XCzxAwjlfnZwJHAnsCI4DWtRlka
iS0NYUSq/TP4I4NGQQfPRLVmJieT5eb1h7Y0cH2pwwAQT9jxQ/JydCJa6yrDaWHE
RT27zOLDo+Ua33uLsRi1woMJC8tw9bxQ9h2yvS20zcQGjPXbDEXGbzSoxrp+PZb8
m78NNnF+clKhnvNKh9LfffSq8gSAK3AhXnMFE7F8qf9POt9OiYGyDzuVhuUXnHGW
dXeHcFyFYAy/+hdBeUgw4a3j1gL5lTuJpFvSxpGKluPX5qplXsEbj5zPgtZcYxO0
DZg5SD/L7I/Ege95gyNqZ5eIPe+v7J9qlvRtZdk0eVN4Q4N5K+MFuzHCC249qpBD
uurxd8Ez7XNjl4deVexvnBHWFM2NG7G/olKXdR0UJZ1mZfziECGlr58eyX4Kabsj
M7VHzLNI6Qho+TaW9sn2fZ2ksQ/EgCDRdLt+TgrpjybO5C8GErpBUHOSo5WHYfdn
QCnbtz9KGI5iLpKXS6qEPYsHaryHkhP53NB7xES/DtNFyJ6/H2j0DkHdeHz2i2Hf
OpRF5FDeIz5FI/HHYSvRYFPWvTchHooG8CY6yn7RCkGxsOdyHhu48WY7totvMcYW
5HF3GSMu45VwBuDF0YlOVinZe6+aEp1YrRm1IvyedcOSixmwjuyqzrUbeQ+d+yku
uSoLESDBegENPc0ghOvNUqcNy3cc1Rte96MUQhnHF08Dcp1BUR/zrUX41WSdRyRj
gnPE+kCTIuhGOEchIVHAWW/HXniUwmWZGkGvdF9RdSmu3Um8xyCnzZmS9B5Two+F
QOZcmWmiuRADeHpMhvznMUBpvMQf83TtjHJbGZPdupzTlBkdUpdo1uRCNktAW5RH
eTAOljHaJaRpwlZi3FRb2uvLh2o+NBRTNBY7ncgQei27a1PmcyD8Ba/Q5b2AkLnb
EtN9mML7TfN5tXPH9kbVV1KzzX5VNqaYyeT1rix0blHtaL2miZSKIRtKi8Iav4RP
xevkvDe6mqtPo3wMsS4p7klSzuMbHgibBdICvvFOaEqWr8nyissTK80AEZBitFah
NNDe5OvSZP6WSti9o+eOjprv3fsvS85T/57PJ1AJO4qGY8QV35M+Pe/T1/yIKLIr
HDAEA1LZloEcbs/qzzN3tyPA9tyAAcz70O30lNxpFqIHJ930+RkUTkS9a2WH9kGW
oYo9/g8NzRqDf7o9K8Z31PU2j9XlEpla7AsdiGv1YyBU4HNXCygbqPh3LYr5B4f5
VkhinNGHDJH2rUpqsdGSkFtRtcyOmq7xdaNa0od6X62fwEav+PQb4wPF0yaAPjft
4MX0me7i9BMkDorgYHBHG9IQlqVc18KXYTUeOyWExxRvRioJzpHDUGRUiTZHUk6B
+GvAUuS8Hod6NBROyFy+4s7xBbMPcjHMO2zTC6BTQbbl/UuaHq6eZV/V0vJStnvd
JeVIzP/JJ9/s7MGqKVnaXnD9I2Iy87WxdEG3ZOKI7UJm4PMY+zOI1ZDtK8jEK+I4
Q6nUFf5VkWWyO+ADxwExIqutvTr5fFR5kv7sQ3cqUxm1pZx4H9sdeViAHB28ENJO
aY2WbRu1ujpigXUX2WC67OA6gnajzLkFLa/sTVwfix+4g7ktxjjkbNa2oS9sqB6m
Tvw/GMGwz3qM2o1OXOKjHB6a3vzBGBmTC1HkqRUGhqDubT21COPampAzBadFyCgW
mhCQQShCXSN1CJquvCU4eeEMcAfF96fhO1oqWT7QntUhbc9kcayPFUVG+fz40UAP
cVs0UXlOj8VtLLJj3MHuJpY0siDa4mOMzx8vP5DCWqybswp89Xq1aPqdZySx8rco
FAGwSU3FiTkVpJjgXFTQ8TaY8/rqGD7wvdeOfUeZExSmKM+8iqAbVM/PGlt2Dqr/
P+xDQ1sSJszhdKjyP2xexA5hXfU8qBzNA2L1Kj7jo9t3GyegGArcRaC5SrR5l42I
XPlN1P4scDHxBXNvg0hXjzDuLfT6BKlxAUO4Ovms3AJ1LkUxrYVvFKR7HN7RNcb0
bSV3aKLb2q/MylmFIXK4SUd2pBodJV3wWKmZOQ2tuFdENf1KCYv0kzaZgF/89DYz
hcQt+wSjSjKk8DE/f7GvKv3z1QdRys1aYBEB1gbhHWPeYEy1tZNL5Nkv6ABKwO9v
qlAzky9V9DV12AdSMWebqYl0T4jKZ4Phf3YaJG70+O7P55+0OyXSRRfmtlHAG7Yy
PfoJ/Cs7zt5Alz7dgU3INU23PLRiu7GmjwZC9+Wdp2jIm3fe18m4LfNp5CL/CWii
LDhfNqVnhtTUQmvNRSlvaE0rH7VHrZXh0m5AMkpyQUnwJuqDjbsfMMJbnzgvPs6t
0Z+cnxn+xpoYP1nOwxNdW0Q0938bCoscg45pBJGtAt2nxxjF7Mfz6UR7wAVyiHt+
nMhBCKQVIhDN/R0h4JtNrHfe6M5tT/2nJdiITJlRnYy0bmisr6be9BPcxAfAd4ET
nhyi2JdfmBIFxs+2LfWixDOP2u/eHy+wPf9EXnO++iBgMH6hynnfY9soYdUbVeh5
icUsJVryh5xZXCCK2N5zqDe8Q6e0o6c7saFGID1ALgSlHSlRJdirRSNOpcYpodeB
mbitgQ6qog5/b0QIgmBrM1Cn/pe6F6AUt7X5yAkW0ltPq2pVEnPoJJaPUWk8ig2d
CfYvVgR4E8SJTCIVkXA9n0ySdgJ9QtrLFyXUtaUO0ERQf24e9C/QWjMpw5Il4iIY
QAT6i/yUwNzPGZfoiYte4K15z619PVxf8bF/8v7x8tlarnFCxz03QHK4k2TW7+mm
Gykw/MAUpvG3OIjUCCNSWv8cQCi5H76TBzMz3b8bWlFz2BQPjgCMekl+D2owPkuF
6ulg9r23JWPJloFfXtLF1p/mUtO5yd2Q2GIfGXkNrIheL0LSyUZMLDy2n9f8ohnf
ZoeW4PLYdPyGKn+4WvEpnsCiAuemMErfGYq6fUog8BD1ux5Q/mBxMyFPVZT0bPE+
DMqjg6PnOh5flJ9UM8382+stEMEuHGwpbXp0IOc8v4hBF/wG4uKirr1/YOSo6dLO
QGZx3dYSDRTAifvGw1V7ptAf4EmQSUDJGCReDWWq6jPwE6gPfoT+HzuuZOc7LCee
mBQpTY1HPbdxdE5r2AMCTYaRzeN7X3AXrj4C0tMh4GJUA9W7Mj890KZuMTb3ct4M
lPz0TjENzlUYSYXfwvtFSHnHr2o7hjC/wWL6BAZSMuUlaI570JMR8woBpOnauZd9
Pn+JaHnKeXRarZqh/ZtTMzc0ckkLMMVl1WJeCEFA6k9l3tZEf71Ci7cTBn0dD5cr
9pl27dx8lLemW66feMEDvYSe104DLKV2Au9qi0F68H0Qqkj98UgUSK4mpYZl29Ks
0lFhS6zx2a3V66GhtyIGGjZ+FpNd0m75tt6JjgT0O3zdMIcArQ8F6QwDwTJM9g4A
dW6KXSGAPm+pZ6n17gW8LPlRhi4A54sB1He65suwqYfMi5BvOHd+kjGEf1ceG8Be
P/xKR61f2qfi7QRtnpmwJWgDuQ7D867EQgexKCtlkVBpGbffSrVZQFncWP3heUri
463hA8xa1b2vpdOR8OycSyErwS/tML44SKPEOct3FlvcZ5zea3d20L6gy4S77Oh6
w40fClhxxNQ+H7ZBQ3ZD/+BUdzGYOzTtrm5/ERefqVUzaFtDFAfDWAgwV5f/FPSB
dvfHBrJ+kE+63Yz+KoQ/iQa5ll5iminOrUnqeLWF/6h5CPSAoKgDkpgU9eht9NHa
GQ83edFoN0Fa0TyKsKBvdDhfyWgtxOIdY81pTZvpqhPQ5YnuSwA0DYk+IcVZokq9
IFnTK3qtTjpr08h+CTKjYawd6gmWtnxucKwaBhAvsn+HU/HbC2qeT0QgpHUMF/EG
bNmUajYafQBqJpHVoJXCGAP2HCXyxaOno3sV1fwfJ1scasUxVTXBw/TN/zqAE5+k
lPCkVGNcxSLePbkr64Rm7uC+qJzo0y31xhL4skpQpISofNldhQkOMWAySPt5loEu
8+DQuv4/7cj2d5e62XnVRyxLU+VzliHO6OOrTiFs9iezdVRChrj2SLwiTk3vTyCq
CSH56AHoy/eiBG6wGPTEX8QsarpKMQ5ALKSxfZhJ75ff/G/B1m0KAr47hmGkcCNz
dyxcduaZrn7TLt3gaWXgfqCkxhkasch6+M3SDbNwz2wkCOGdHX22glJUWXhZhDT7
FSlnqu7KI8a42kGzDiJwsZNnt0zl3im6N2FRmkaol97xeroMNFQcTIE1LznixbJD
UbLMCJ4OhJ0VQrcFpQD2695SUlwiq6CFoj5tg9GDnU1/ruedOwWw0ITdqU2dCU/r
60vGskV3Leq+NlFwRo11NGu5lUEvMO3HOhTOUL31B1/bm6TM7+hNWr0k5LcYfaIc
QS56RU1rhC4ZguoGoqFysnJ8v0BEay77BGtOvoJeqTMYQGznade25en4p+MpWU9F
XnFejMKguPXXXkPi1onCcgvHySUIHJc0ZPT0CZnwRT0CBvwospJYH8vDg5OfLj0C
s/zUng64WMoRYXpmcskIPpy+IWguunDxuFzbj/8cZFaV8UqmQU5XMZRCLpY1W24H
y0irwQrncuryXx8ltz2RH30kRYW/RDUo4HXitM02PazzyYTsBIoN9acssmISsyPp
44kYULDkPpZkdg9uv2NHSkT63RYj+bsQFR8uArt6OkOqiKU9HjQK1R46f1uyWrR8
HzeTDCzLgSX2FPObnvo7S5CWxxnNMCMnF0QALh29EKWBRHT5qwV2IjMDEFCnuwYA
CUgGMh/TtTCIvhyHnwExXuWUFBpWTdO12U3udM4MYRFV+ZhXEgrDG5utN62zlYPx
zzrvtGyVC8HFeXRcopYD5Wt75ombCBwxKAIZ7xb1L9XYOqMZfKqv6e/gAmnbbIYM
HfGPYkII+yfBrI7Itio+agx+VdhDK0Dx7/tMJDZNQ/6KbRPdsuNm5Xz8IDibkwvW
qxIOkoMttvy3Bbe7hPBjHAAxTI0Rg6C7cqFW9dc45ePLqGHbeRZpSiNkBPKcyWIQ
6dmSgsSYDuN6gvA6KFY4MiyvQuB/3Vuc0vvTqRktCqvlGrVMgGB3VAg0zOGtOhjk
VW5hvaz/G0Csn0NSESQqq0W5izppj8DXttDR4WHKSxl41OAxQl5DN7S34UJnIC4I
QhRRWCccs3fwkNGaW+qErWtkw/0WzvJti4uM8//L1rtxZ/q2c8q4AIT4i8OMDSM5
GaNTAyzs9z7kN3YfJ4pebeJdJT3aZZiaKqAOmQX1RoHzrvcxX4keSygSYAhXYXHP
WNAfI+hEd1S5IJXbF3+hFVAeKJmIeOQ7X83XRTMzHytfxYMjYO5YghPio6NpHc/7
Lf+QJZscpMU235Ylj/xnKKSuJBU/fk5Nqa37eErGv6SRpVRO5uWU2MwcdhETmrw/
P/XwCQEphqTBLoIxNfiSJv5GxSond+jz1V76dCOLRVqL5QXTyd+UiBASDtFhkh4S
dSnmIlnHWN/mtK0AoiyJxcOEtlfWvbg0zgxFtKsvpiGzA9ahrWnbM2X6QjqcQdAS
s+M7+vBEuO+gLdRiHrZwzICe5yO8tq9MScXrOFwU2DqE/XFCqbAbvModDSkEz6T5
L3vM+SmC5atxDLfAD3eEPFKBATS6/Zc9S3nIcXsqOzEFKUWDmH81HiYCEEdQNUdd
jgckxjoceo9PbaV+723MH0n3i7Z5hgXOAE8Fn6DqZjA6nHfiL9w8HTtcstYjX1pz
NRerNnzPXKs9n68sCN1KzJJgUaSioqG6G1WcePcJ9X+un5h8Ia7fiFRCwq0rHVK3
CwBY05j6n9DzasUhSIgt0HDXMDJZL+0Vo+u3rNvHD4gK6srypQdpEmuL4KEzFeQ7
TYxhHx6YH54PfntyRbDcBjsk0KoOPgRKuY3AiNdLRpwgr/9ANh7bNT69XAK52dj5
AqdoKTrqJveb6HBLpSoiL+urHUezbvHo5e/OA5w4sNIOxLspAcP7KxyBNfXfomGh
8zjKMnsPX5eKgAhvVltOWNXRrOdooMWsJ6m3rA0InoX+trl2qYDApEg2N2WiVLNp
uFNkAjLBsFVB6BpDLpj/ZNCdqdIzdPczAOAhBuOEkOc1rVnRIkJI3yhKi2Iy6npA
qx83aBTZ9Fy4Zb0SfJ7EAlTVymRh8hON2Xt46gUJ5CnykwahSppmazHwNwOLoHld
yPQP8yI8lCCsqIBcq85yXXk5McjTq8dDNl3Z5MwE9dxaIXbu/QrURMsVftz10TKY
IepMZMmqEu8s9alNm8hqaz4NWuIyRgUSBWTs38HNGCzc0DkkEgKqI6HkP7Nh3JmQ
RQKpFoTfgVN1Lh4KoV8EnQw8qUds0/Enntk7BrtSxqKfdNO1fTMZFeHoVlQsBsIP
fY73Pzy3PeJH5ce0sqE/H7WOhrbARDlqKyecOnlnBI3lybpqlynrQqBh8v4tDS8G
74zWBsEqvpa2rpOs5MB66a6HDpm+vgc+5gh+h7GMrFaDBxKqnb8UHK64pAoxAV6n
`protect end_protected