`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 29664 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
DBGZtUPdvgnvgIFp6VMrQY+w5n3/fykK7PLWV0u+wbjxrELga8fEt+JXenYOMVWM
THOEqMAlTXMaozuoWhN6LxXxB9S+hIdh3tL3HU1HXWboJERfyTARM50bLJPs5Zpv
EXWbM7opJBhrOSgHQaVKktv1W37cMiks93bQxYnJmAB+Yzk4rkdjFsJOM5ST9u01
GQqy9OdvgBjTQQXhCWcvIT6y+cy59DLFRLpxWkouetd+yiAWvXXGYMjv+aGEhTGd
0dD+YwcHdcr+APgpLKgSgFdH5sAWkio4Szp+PFFkwpudz8+CPzzf5ITXCCFq+itY
R3JRhtCCKHSltT4sRrKfrgOZ6YUykaXAIpg+HDnNEB0OkbkbyUD8lUKZQ0xjv+zY
aYGP8j0O4W7Ef7x1t7gPSArqrpgAwhn42Qhqj+LMJ/Hw4vG+FY9m57lpNJDIkIMx
sE3rHYtuq/5vvzHDRAVJi/Tzz62EYgEhINh2oWQQbJNmtZvTet3FV7OG/O+paY+7
j6PX0sXoOc99L2Tbu2WPZAHcWY8syxDdg7lt0h7m7U1FH/vnXv7Z5vx6XMGpbL4M
x6GGJxcUr8wx2s9MMe3aP3+fAO2l+olT+N1fczOt6N9JV//aMJiGolMc5qorAzx9
Tgplj12AdYWxHy01CmiC4KPY6kKYr/iLITGWlNogYW/uLvOM5EEVjqf8+SBg/ivM
VMzZsEL0t8RaZQchdbn7qWhpfu5dzOuUpfgTvtTpFVUDgpEGQJZqU2TTemrOFvWs
nqR7zLyqDK/uMvGIr142itUv30nNmnVjr8+Z5/ywWpWss31NHXSkylRTxc2My9cY
rstHi98Nh/oTcg5tvNgNlZYKnHS2ipBfJzK5RelRxLQdVme3oD2pTwHBEOpl5FWd
4FtJIoWhFwwnAK0mibLKOBZDO3XiVeoTR1Y/cUL0OE6tFqNqM897YZRWZichCJFy
PM5xLC6sFzcSRqSIouIDWz2GlAL9UR0SMomNQXMmBAdGiKlPDAGbZG2Mp5ptrh8f
nYvnIVSuoJc9afpz23PIesKcvR0KhSsDU1T/hZ61st1blU2T9ikIVqQsVg/9B69m
u98EC3Ui54+l8OniiS1ijxKozxI+wFgxE42ZNPxD2Pk7ZbOFrrR3Cnn0KizYwUDO
qHfQnHgK3B3sh3/U8COVfb9FSwBrZddmjm8Tx+LOAKywmjVorfzB68pv6orwJfz8
Q48Ug07QN/BcBcBW4KlnYvqoti6+Y4U8md9Q7Phy+EHnz/X2baBFhM37tHgFZF02
7i+a2JF5MNA6vue4e/wbEz7vfZ81ma3DUqK+8h5dcvgykNLBjil78DWOy5CS3wo1
ztDcewxQxStFiXV/WUPG4F1xiQFSnFsf1j5vhDW1YzJ46c4Nv1pjMfXHKzOtqBP6
AeUNno9BkMnurjXNSwXoA8a1IUm9n4Mvb0TlcsoMqnE15PUF1AIyeDc3HLDF60nT
O1nMv3LFbdk+bf+le5D/SKX7Y4U0UZjsP59hKP18vH5CeQyru6E45mBEJwMM9rw6
cOqs4K/jBAJt/xZEq3eUzQK93zPc56JHUbzLvsUvCrRsbtRWd/UFiuvh78H0nph+
IwkmgfO2Pw4o4Z/1kdXSwLGvXYVIo3utwlHExq9MkyTr+gRR9iGB/o6fxaCK5Dd7
e/PKcvptfyxyuhhF2xH9SlinefsJmi1OOqzlj+pGKUT9OzezZKhtTTG01njuCOIZ
iU9JVyuH6AHzXev1roNLPCjemy1c2RXOInGWdlcRtOahFa7mnJlvzWSTThv0nNmZ
sfY0/bF741rWrSzYfV6dm3DNi+afIBBXrJHSP5BtDm7KYy67cxvI8hHXUOmDxPni
UozaT0okXC+e9o1MdN0E2eLdAje1dqEBuYFRtYChCL2zW4zmfq3IEVMWgxNdFWa9
oPkSnJRCyhzBodd6hnrAJaQ3CfCEdv31/dtnY9pcAkAEQaI40G9clyRv7yaiv/Wf
W7zXAJq9ErIaIv3Ga0iPBmYedRFv8gKFzL2KULU0gMdkrIkKDlaqIOBxiIrVK4Fo
PZn6+2ohQy33/FvXWSkntXV3r8hA2nhwy+KzT+q7BUrLBnTqeLtbOq4F/1E8e12h
A5IEkt3Cghm2UyKFI3pj02V0NQtX59NHyJUe9X0FaLDqKET97CZUNZDvj1Ulh4ka
pmUBfvb7RcgDk+HAEH9DAr3tpSPpoPv73mYyIiU8vp9GZ8RZbHzt3lLaHdOsgbTW
I6V7GE6bgBUTI/Y9I34jmymwbLKoW7LUmW3Vu5eCIahuN4HE45/QEIa3h997rdpd
9zmcFtVqDWe9HroeC4QJhWVjXDzQE5jbex19yHeSIJyG+ZCxfoLfHoW2f0UrdNjV
9avUNIHkO4Vrhb/I/yXzGnsbd7d4VwgtJB+OeiwF6gvSsREfEBudGTFd68utZo7u
0JhW5+a/7FOBgrU0TKv2jScW4c94YWKU9KUDcKvuqFflsFgrcnXNFyHemonh3nOP
H8UFDOZ22bg5vrpert6RizmqjCPYzTTljS5S9xI+iYkLBt5nunaaYhhaAtmbrRMV
rloMdOlMdqshSR9qvMENl0xvAQaQtH4rRHCoC0zKSWKnldxDX9yGvgkuA2hDtPDH
ojDGzg0jI2vkSQDBujsfQDevnzaixPlQxrOe0d6+Vka7NKetvrmeSf6UXkyJh0nC
uL7ohsGr6/w6wOtVwIlZEXvwvCGxSeldyAgFAyzBmOwQtzi0uwXos5hfpofM872n
EKkILhyCx2Tk2Vi2A0NCojWaPB94Y3y4gA8DG9octbcwcNzjWX13E49eLe0O2aN1
korIqVen5JwfML8fIZf0tSywZlHCXmwQ/66sCVvYv1/A4PslhZgDPlLffsZ709Zs
EU9uQrHCAhw94M2IxSVIJhhrxgP4ohij93hOIpSnPToL2ZQ3JqCohkqDtt2NmDOt
qWU9qhNPWBVjkiQ1+ymKA3TrVboyNk7WZ15JSy1ck2fJ15nzwB185PI5WNKZP02B
CDLLLW4nyoc9SnwYEuh7gB1M7Y97ln/KxPkJz+I6TKI164Dp24GFpER0OFZkhvSv
aewDw9ONG2kCjMv4TQO9j4iEoEg3WymByXt1lU5Bd0SR/UAU4IzaJsjxXGnpf41N
n/6vUM1BzQP6Rmm/ssLJNPiokWtoxwfGF6DDXiit0yq03C/9vGqF8FxpolKasPVg
eeemkpYooMOkK5vp/Qo6q8l0hPZvL+cUmNPp61fFUIP9MKnNqwTgoXadaNJ3zeVW
6C1PTGOp8RBL0K652vgXh5+QAyOXy6T9ksP4DAt0ROuxjLgGlV2Fl7vFQk18zAdx
1hAkWPEnGwcKnrS+Dl1J0WefVNttmH0Ws8Jl1uVueouOHbW136M2nM9eTgINshkk
GMlhbM2t8++qctRMYC977WDw3mkdnDpl+wp88W5yIInYC2ooHpkcRnb6TcWTAYQe
9otTzcZDrQmeUAF/T8mrBj75evVNCwAvuKVroFAHfZaYc6TygDUT5SEAx2NqrMrQ
PfWRx+YMoQrf5QyDxiq3BfL0fMYcuJdUWd/HYgSkeF+qzlKGubqlWtd6Qrb2k5kt
YVufnytL3mSHB3hVqaE1RQl3HMddkIWfRLf/XWnhYy31+SnygrHKfiQdILozxC+9
cwgXQlg3IxubCEBOCkilzuts7+Fy4fJyPni9UYFb7MpmVDvLaM8X77OxPfqN+MDo
VDpp7BSR3nZGZrZusURkaBlzpICmbC0o8DRlqcoebP2b8/32A01QbBSyYkBbs9om
Ig8uaz3R58djGowFu3DNjVpnOTp27hivpAavAg1QbLjokk7QA2MfkdAJumUaX7L2
qao7m9cQPRenCSC+tWy6c8GhoRlg2EsTkXwzcYBKXlWfaNojO9vBaRQp4y4BNz49
RGk2HNVf7aeNZ3AZ5IaDYvklmhsZ0s1JgKTMuBIf/8QIIYrZIx3nbWiZ6E7tp4dI
MgkE9ZVabJrET4KArOYWycao5NBOg680SxF375DYWvVHA1VmYs34xnvwKBXSzocG
S3siyqTqUKeMEPFScD/q0VAMlS5KeewPabVFVrPc3lsZAbKfxnrQ+IJ+b2BhdXE+
wsAqMig7n/M6Oa3UsuysrWUZEroRpSHh0uy1/ci/nEk7EQpYzrG5qNJHQI0PKre1
67euG9xv9RReDnGUGK7nqMgPGBinQ0t6Ds4LZMNNF5RKhSl/xoBa3NPYbOn5zdCc
O+WKzGCXVPwHsfKxJm62n+ceWlPQKTXJv2aNtc0s/BWd5sjspKbtbtHYVkezz/VE
PKSpYb2AKebzGUHlLqsndUAqlHV4G6wrw9ud4HGJcqY7Ybi8Ht4qfEWdliwhhx4y
Ax8E6obWQqlP7k/hASK5qZ4ix9khKpFOf+ISbWene+lCc8MYuDpiUed5uTY/C91V
UDxj/sqwfu9kmeP+vUABJVBbsPi1m9vRvu0GQ0qnbREB3F9xmM4QHz/xJpor2Esi
z4RYIsE8kpa6xgMVbiSArbpDbUGUjgWHztA/8ONtWLN45AZjsS2H5qTCc0r4+thA
miltF4O4msbOcTJ4rTpgWj6WuvEOvcI7FCxRc2wRqS2bRgsSe4TNE9j2rL8D1Cpe
wKepc/cK1h2LI3jazSucji1T1XPsPmFkfbtj5f3pc15lHTo1WmQwUljdStHNYwDZ
vgMtUNFOiO7nrplFs/b4IXZKENPZH/skrYYjA5vWC3Wme1OnvneU0bkdqVnwAENw
1N0vCIb8LhDxUqDjDAIK2vr1J2YXkzLNWAtseY8mxh0Fd8OO7uS3C+Fmjtdgjt8Y
Q+ZMJXs17psATB5f5rhOdcsKJ1wu8uusHTAJX5RgEPvGDaXNzUShhZx9GwK+U9gK
TayoeeMTF2rnx+3Eo1GgRto5w3e/61G8zGDvhOdyzaupzgGKKJIe9/PKHOHW5Tvz
S3aK62QdpJ8SzqcU22Wy/IFi4/7gYslqyNVz1OT9izDr60Mh7Vw0QDd0KQy2uQr6
XoidhdaiKTl2fGu4tjtrUt5AO9BVbtlISUlI/rR+j+hTAQRG6qOCrhiaxeiEZ4Xq
CANtzj6ltyeeFyPVh+tHEFVzvToTyWvnHxQ0vgy5r0xSfQ16CTVrIksMQH+m15Jw
fz0H4xuI9EQ6Qu/Y1YdtsxjSrq+5KKspd6MaThwJ2TVPMKOiSh8UJnURo6Q04xar
xECA+PF7kGGEO/mxVo7sXo3q46SQ9qdmZuCfSO7iSE9vVLrsaiZmk3Ei1bw2kCMc
VWrl4k26wkqC0OGcfmkHv64oJ+PyZ25kx4N05ksIWsJ9YPAVVxkj9Cip3z8TLOKH
OV6rZobJOfx9BZD1QBvF9MsroE7AbN0Uu5vs38+pwnQf6qpnNlRIZKShKBRtcJPo
GgmFdxjGBMW+rLeZorB3Q7LrEOi4GBf8XKz/DgMBnDXw8xUW4CrnvcVRH4ennYFY
c7kjfxKo889B4bfuhcBV2+BP/JJvAK7arf9qhYez1wgVEYktqZti1HX49/OqnD7i
cyABydOHuTmdXPwaJ/si1lU5tzF+yO2xgiH9aznZIZ76R/jSqxyFyYZVaY7RjvR8
eAPqEdA+G8WiTMwxZi/ZwrhLxcNjG6OX4YN5LO754pz7EYED7H9iduxkomTZLVkX
vhyZvhsiF4qdvkx6TNfpcaTS0+OzxChAzLljvJTHE9Xg7wshsoP4tgGlXNrvr7NG
kavxyApG2VixqtPRAXKw3/yz4u1yPG6EJLRTc7/olx1yrVKSsCIQybxL5obNDBVo
6+Mwlp3/OxB8lJQUPSJ6DV+Ok4xEw/EvkdtYgG5kI6nQpG++IATrAXE9ros8ugSR
k/fXnzqUJziUlrGTL5CNX3e7JPkGxpozzulpZaM5YfJV84p3dXICF1LuoQ/GEDdD
mh2NcRH/NXEzND2oaEHBRLEsCrjrHXH6YW7oqN/FbEosnY3KYuNs5xnIMgHUkPW1
jfgMsWBr9fdUnGEn0zMdqjNDOj9bR6OkT1aYJvA0EokrdsgVYLAx0uHyZQAK4idX
qX1Hdu98A0jhTD25yLMm3sPUe+dYB6zwO2XceAME9qzCwwEh9+FACp9B+DlD51vM
t4KFeBlHV2Rrlx8AJGoDogAZoFl6opLHu76hncDwP71gDQY1NmBdtAeEffeXSn9H
n5rKyLMevD2ob03bTG9AeCymazA1udUsT/jyU6TFpgPaDCVv52nZMlNPoKCMpGsE
LYoc6VE5Hth97IQSwzyUyZc3gxs3JrJmEyRwKvO68P3CFHTjJWTrpkKvXOa6k4fF
NgQE5yEQqwW+yrD4BRFQ2A7nH+oY3+QGh1lG6A7WTALWfUFySeHnN+G0kVTvB/Wj
uUmaxg6vQW8osM4tITsdkvOCq7NBgSL9Uo4JddB9GBVCKnnxUk/XiWStHK7McHkk
gr7dbm9xamB0aqu4SkDR5Nq9IlACwNLv3bGuEkr9H1fcITuRZZA/VmYhTWodTuba
eFphLqxhxQVkbJMGin2aBjp439ei4uhRRq6NM8DRNg5rRmRe/uWB2eYtYiEZmccu
MhEcmnT4iOAJ+mMLUEOUBnxTrcm8unDY9nm2o+dOMD6A9ZNkIdqPOiwGGVuSRn77
uHhns6D/5NkhfgaJSmXDAAtth2UXBq6nlSg52CUDco38ckwTZimeZFlImLCJ1Gft
NMlQPYUd3ei0dK8maxcM77njG7wCDBr7FCqVDSDx1OMRSHi9vQH9DFSxQBO5Ay2a
BZXnbtHBJAReC6pTl5SMkf2mCJ/jlwFay8gI9jc8q8ZvOp3g/2BcH1754tKqfa/K
reiQZv/SsjJ00yrS3VZbGCqqRDammffXQOfeRWMFkV20vw7WegcCT2ZEKlLJxk3D
eWqtmX9OKqd7N5As6CRPpSCluMPiaGSShmBcJ4LYoSf4vHGYA9GH+aCNH0lbEDPh
dqS6q+QXa5ZPZ8+p3G7pPzvudauLb9ZboLebPTBA+D6pU3VebADXo1rFXHMwhjLk
JYD/3RGi9Q7lTA5aY3rpiMr7d0V3RvuNIBkZlIMg9wHM7wr9E4RQk8vx+0PMND3P
TijX/qjaHCJRsu3KNcfo4fwi3mTCv+OxxWtENVhh2ylruewIiyNsh1j5FKTYeNcl
ZmUfnqFp/u7aOLWlHUNXj6h2X2Idw/icIlaxL2YYObqQa0Y26UaY58nuYHTjnmZ0
hQ28kJOQU8wAH9F03XAsURONK8ll4yUjdfWiboxjMw2P23AK2TmGuRKbDDrM0h1R
Oap2wjnMi0gfT9lDKWGmPuFAa6JqqfJsD5NZH5TD/6ptue1ANQ2vpyuNOYrtykWD
Pw5dCXaGSNgdZGqa4Fh+z0ljpBZ+exC+GGU1vmdEVLT1YmItGcbhz9/YrJjCDIwB
OcYq4rwJJ74OUXgkEiuoWY48aNZtBlAOgNNTxDyQ2AqcjdNc4yDgVhoz/khy5JAK
7PSeP2bKt6pexrk5MI41GKVObdl9GQ20Rppz+EtOUHaGWjc9xbYXDMAJpQB8emuF
ANu+IR3rVmHizd9II2QPOne2iRHKeL2hLgOCpE+otiPcWI33tLPwVRib7vdsUyhv
KI0QvBS3gJR5fyLB69S5wRx6nCI0CCbdoORX8umsBJ6WPGJ8tCHBypAeGCsRxKHx
GdfA4l/utpmxVE+xIjYhEYeQGn+M4PpkUALVOqBrHkiHOMDMw0qH8g+B/n4ciFTX
5AUsdzdXF9g6fir1x5V3SYMBzEAY6BZdBUldispybCxtLLDXvNEg78oFrM9a6rLg
UhG+isNK4U/DhoE8XabOV6s/8mXI2MmBWEB5JqVG6KktkajkQhAZ5o64EzitRbLh
rlV7nPEZFByhL0kzE8lJi3vbIwDrb2Cb13TG2FVvpM0v0HIi4VMcTXxrW6vwFePe
XOWdf79vzoWRS0UUrMh9ntC1SnIL3Ck8DfuiIrxIBOPLCiyFzNT/zLbP0DWXsoJ4
6mfSbf1RwfGpDhckr87gJQzshix+NrcxfO/FakW9kMnRMs/oDNBmQ50W5i/fxAIP
5ztgU0655vmeT5hcMd6rnnmqgYCPrNE0ztpUsnQvATYzbpGh3O5RECkAlqhhjURS
kmIKIFK02WthW+aDqgVY/b4xtr6lbWx2iSB2GN6XfZ05j2+KMPJKY0QxgOnK+yXb
iBZNZW8+jX0TxYjxHyGBgzUMsNL26QH2PJlZSOO9vf8GmZC42QlkfzyBqw86xb4q
DX9SwJGNbjjPfqmMYEWqFblnwsUw1dzCxbF3O2224V9ueQWt8K0PMiA5zUB7JtKp
1kyuKynzYdNrGuqmKWeobfBTuZnvLsFh6a5VUak7PpQn+yXmXneuERnP1Zan2Ydn
dwaXTaZxDryCK9XRKz/aWnX38m1VGDRdNVjzHjM7Eo5z8A8L6KoIbTC1Or6g9K5d
tGhqKmQ0J5dnInaPRbnV/NPWOAZPskZqQ5TQfFl0bSW3+9DVHPGWF4Q/sw3zIa8Y
YZiRThX0EqVBDh6WUEixq7XTctSPT1TcFB8jdF11iC3APbOxGy1H3+oAe6k+jbHp
Lz8RPu6l/H1zj8WO19UHuseHyTNj1qawcCdro3wPMeOYqitORE+47ktrqDBAXXfl
TDt0TEWNR/eWs3E7jHw0ZuCZlIqzfOHI9LnM6p28edPFWE89ruBn8EHFWQRqCdiP
kQOJ74RhYxRjmtb1gsCh4XMGobeLRTORGmbszXPFNwQfm4ZLnByspD2jodUhRhLn
hIroS0x3aWWW2UdTm/Q/Bfxvx6coDj2BHDSUsjQUEyD9w4Q8D9nIjTrvLG3/sCKl
iu15paUwnk9Erd49HPX5AjWx2zbunyqJT1GmfN/FZt93ATJMvhSC1xs64mMhUIh8
kkN8s6oKC/JhKj6trtPL5sjyCUez3R3CWbwnSs9/qS4CGIwnOOUowMWeIdbfTa3s
EKxyidPIOVXJBGlawBCtath1jejryCFXeZosaPxG8sqQszBq22jtdJ4uqDkaI37a
HDBeqikO7v320CHo5i37qCe4mU3vk9DhLsan5KeLPPaP8K/sUq9I9KTmeBy58eL5
vZGrhHIbGxXhOOAbHYyfmPczkZ8q6rzHQt2sQBHOGnSlfDBW0JPEbvSZX5UKfM2K
EQKuFDfNb76Imid1BqYcY8RdvJknvQ8RE+K5/87vBVee8q2/hCSlyDGdt365s3Ea
6CHa+HV3TP1kymap8RLOHDa9Iv4G+1/tMGgvSJZ+O4hFpjqo/RRg6u48jOIr0hMp
Mm71Uq97DRa+VdyU7upM16ZM0TJng7R5NXjKmBKIj4hI7fQJt3dEyNYxlj64P82i
SJgm3bLOOD8kUaEZ9vgp4fi1SZbC6ETouB+OSKS2Tn3tYiS7/GTGN/U5ktNtGAJ5
9/Z2AB+TUgC5gOu+w82FhUrCKxAPgSLL6QMLAe8ZY2oh/xV1VNshzZ6BMg7CfnND
cCh+/ExVNhtyFAqgfUR17fac3Sbn0iwb0RpMfOGb7OZV2IIP4pSWRjHenOWSUdfR
1KwvzNOdfY5FTwztyfnsL4Wx+BPKAG3KHwSgh6aEdAXHlzFQsZ8H8/mclNX6V1ll
rWaFFnRofgCSMi5hZ688C4xmL94sz6u6gx90+TC5LxG99xDLNftAg6a0I7iINeQV
KO+uHmcEJRl0bcJMCaIT1I2OBy5C5IRddRNPls9KMtck853iqloL2OuRj7tuzTjH
npnKXd9cJcvqnIiqR3ABvROtyeI/nF2BpeeCv4FVQ4DKwUF9hXgp1yugPuWiK4wS
u67rT0Zdzt2M8DEu2jAFuQh2kjwcfEH1hRzJTtbEJlNVyQjadV2mwCsM3OvZ8VmF
deBx1sT7iH6sQSQ5xGShbOc8Pn1kJX1XZLgwUCdjKnQc8SsGBITt/1c/gOrZQVyI
lM0XBq2sNnjs1G6IZhd9aRYkkqwdQbVGpocZzHzyzfCahwfPe9yW1FgyzHlavFHM
k7PD1BgAIVJcw4hN/sljy7CeBcq0jJxsPT6p3icIqax46MJcs7x/AJarLFDKt1R+
wDFVkgPDWy0WoTWEetPfbMdmb0gBOo3nNHxrC00fdhg3NNPx2sfPOYwcBS+StqII
FMLU5jf1E7qm3amOoFkLYPXAU94+3h5LFwMJycHKicu5nTX5KPcPC2PKbVvXX9uH
qgnKAx6V/MXW3Sqg2ymYAKZa3Lj7HvAr30yFCiSUelDAatqmSnF4Cwb96ati/OyH
EKLzHCSsYAwzdxy4GC4NeE5KyvAQoZ2OUiQtdgaLP4VcA4lCh2/RthjaYDn6o75k
7XDc5DbapMOWQgG59oJeRTCl0zHqzoq7VW41a2Xp2FVUv+hutnk7e3hHszZG94hC
nXiEGKC93psEZ7lm4CbyuvJZBU3IyHe5/7lJxXHSpxq8pHkmKlJvETHQS4aSgFCv
DcVnes4JnweBmS395oDnM9sEiKo8c1HU+q8DWyx5GpgW3qttaoNZG4zzGqvOU2lB
QtBT+AF/ypXyXW96mXzyvljxwkWGbHrbR1qMYQmUfDt9LmwWyVZcdEPVOGwWHBk/
54U1a1KTZg6f3S4E2sxaAZrTQyX855tor1VDRi+v8khkTQavS3EwOJ2DkNwC7cNQ
Sj87H+TR8XmVySgA+36WU3VCmbO+Ip6UDGR9v6LFpZGDSEOeLXmVHBanJOybZDf7
1LoGdHOG5H7hWeM6cdo+MD2RxqXe6lg7+QC8Fa1IXh7YpojrIqtrA8ZAp/BRWzyL
xCCK2m3txAgqfUOq1DHCau3iqn2hBqbj1N5aV5IXk+u8fB06njr92Fm68Jn26kWy
U/Jxf3wu4OcAt1dNJqvjgcaF3fLLNr8PohGlEzfhLpYt+e3VRAb5fP+6ez+XZYHH
ZFK587FRoCi5PWUVZYnlrvwGWlm6auKKwIU2/qprTY4mBhxuzo6ZPHuNIhlPMN7c
IfVKOR8E+pmtomxmlnFn6Xwn2h8kp6k6/cZHhfhH5qrt+TdjDNHq1wMZubpndsVG
eoAgl6XsdBVNm/QY7XfaMe2caA9D58O+NlkiqmYtiX7cG2tV4oDT/b72BJiVyb0U
YCW5Gk/mKl73YMif/V+m7VnfZLpzULiQE3bTzNAEiBEJx0vNSa93uEpGp71dc0XK
MKPOVjHwlTNgLkpLuPcO+E8A4C2WV/098boPDd1bgndmqfqW6DjRZpstsmjE7vwu
dH0zlsbukuOK17fY6Pv+zgOtfpvEHTF01Tvlzg2ntWnwAoMVgaSBP47oa2j1Jm5N
X4+kPzhJOSNxY+RbUMzPlfR+RSnzugp0c+3plZet327eDeqq8sDA9mZ4V5HFQ2Gq
sz8clpNp93Rl/YLUp6QpOWm+QSCw/4smSQL+zBSOqvRdY7nhgnIGtBSDjcsu4Ahk
Hw1ZCCqS8hGN1cTG0dWNy7f+AsLBiJE4+iDdNerYpLhvMevMBs4yj/DHLulgMCCg
VjLZAxLETw/jRYDZWxDRPYW9UhTe3Cx4hphZiP5IrdwvvDY/D5ySxscb9VPUS/5f
+7ozAYiM2YiOzq+g9+P7tS5Zuyr4n18oJKnrM/FxkvKLDXpg7oWh9KYWukvyvIpQ
GVDt6f7gkdxLmSjfi8GfdWuHPz7mnMKFEwnEWGHhKhwCcpZgVgD7NRuC4kEq5u3S
wMOi9NFGFN8oZoAUZQg3pY/zByqDqF15q2cli5kOJlZdHqDd4DCN2Rr3v8G6sN/g
wLyAPL6THFjlXyz8xL2JQpmV+xNjxmSiDoT04lU2fezc7DKuWcAz1mOEk6udFRo0
e6ii8pzk8hH3dRXKJRUaeUr/EDcwltJETOSlA0J6v2/e8n+TMgDnY9safORIC9Gh
Wl1Ps9KkapP2yozD5NTq+B2hDu3LVDuvTlBLaXIsmolnaj9d/u+KZEa9ZkYeUjK6
4I+2BC0gf43I8i0vd+BYnxIH/mwGR1yru9WRf/YxOodm8F+XLz+X1fDv0fot11vk
Hf9b/8iKFQORQ3IGMgi5ILdKTnIol1h0oxcoqVH86HeO2X2lH0CE/zHUF7oxK7uc
XCU+NeUsD4N4MqOO0cIkiGODtoH0gQjvIc/A34xmglU8PJCWkzS1HS3E5HX6dy29
y2O7yQKWRG6F0xFif1hbf3LgQYGuMdvj6d1BI+Kz52HNRntBcv5/Wq94uJaUtDEf
uohGpAOmQZ679yp6fKMbY8/qNlIaz8JsgQbGdHCtjky6VHR6VL/uMBLb3r6CEO2R
72JM8TpBI6hy7whQfNsal01yL7g1Qzfop32jcfT0LOggsAqLTUa7jzZoidMZndA7
fVdmsnOcV9s7gf5dWjfMeXD57zYWXYbAjHGQ0gHt1cXtEPlNajqWK+ZChfQuxFyg
T+gXeJfLMzHcpMeItkpPzznc84afCfl44CKLZc8gQVY+f6n4EQnQERLioLUvtcPf
dMqAppWo3o+gUhbDduVPcHbm+Ur4IriNvbtwTRbL1Dkosqgp8nkmzqEoEDDd3hSm
zMQZouJxf90O1NQFUl8Ihmw04INduIqNOJIl4Q72TxJnZ1r2+Qg760pyZY720DDa
ccYjuGLQ8WHm7/7pU11XG3iu272tZo+CNj4ErQIIgPch9XN+5iHWQAYE3rl3zBa/
KxTvLDZtOKRPP3yXqkPeH5g/rBZdYpjMKJLs8B5ke9K6Sk3g1/8HheIJRe3g9JT6
uDzu6BYZIcSMN++6KZtaFQp8f0Gc7mckkQa6S6K6BU+bfl2G/+O5MAHiFrjdD33t
LldkPOBvdU+60U4aJ9wWZKP1GpGX2b2DWe0iB5n+iZNQejXKNLmJHj852n1gdR9e
KEvJgkQIZA7P+u0wsixg0+zxXvCq8t+fB0PmzcoI+eCsUEzBh6avpbu6jzp2Zbwn
oh9aH6TLEYnGBIG3k5Yz2f78jI+W4QGDWCYuRixiM3tRkoMedoRTe07dayv5rE8h
MCRAKQApgKLaaJexfF2wu2zxHCgMvoQNirQY5Q7Aeq9Eew1/YxKqXaTceFEz5P6s
W99vvjyXN6YYahASVkz9ppPBQskkLvC+wXzGW/zGhaNgN/m4kQ9JKPAtPJjhOAGJ
i+kxrU6sbtRSaCKXYhZYYjtLdRt4FdairPEcXGmBGRZHseCVSY7HYCaiTDToz/sH
zb4/vV9p9l0vPZ6D79yz8yRgZV45yvyXQ+tdSqBRG/XNjrnLR9zEviozC/wLkDW5
TQaAocYYv1BfvVGJ1nqZnTc7atY7rjJfjjE8j8bPML0p8W6WeEgAYvM6Ye5zyuYM
lgrQ7MlNMScwfqkj75Lauu6lIZSzmN3IzCMRiju3hWR6Py24ZfU00r+naWWDoOkd
q7hY3xEa79i5Gs1G0lN8RjFK2UkEP+Ek1f1+UdoOzT9wSM/215iIMw+8mxWlRBpH
tYgBD8wHA4KCpq9IUxpUIiHSgVmeKseZ4V6j/g9c24nvSfRUC8t//Wz4WcwTJMnB
k/ZUTyuG7BXPaZnWSIqsEncosxLMDgth2+EH7HWppcCIYUOZ5mNXWkmSR3Lo0cYC
d4pQwt7OfXveLsSHgwOeaiedwE8SC7WgJK5/0Q26GlOU1uNKz6AJptIAe7bNCdRM
MYRebkYLLc4SUk7FHTeXLzT+JPktlz4ZxOlUD1E8j5mhD7JRaLFtch4BTxkz/kA5
x00xyliOp6aAd6vMK9vyabizbYv+qknibbrApdEHqJm3QIQNcqUaUXK0IblyOQhu
Yv5i4skWchWS+eoYAzhr00poJnk2utXLEi7AfqIea3DN1wY2G1LPj7kMD3n4WqVA
/PoxeikfRTJDACw6blPu4A8mn/O66iFJFAJm6yPg9p1aGrvQMr5mGMv5ysTiMyED
9Ws8EOc8iG3rYgpmFQ+/z9CTCCFOQNhO8ahZfYBHjuKZsjxTSU7KKTs82sfzXWn/
MYfn3P9LmusLJHCQr86vwNZC988aCYOKzrPZovDFGQK//WiILaB9LzNXh3TUQdPG
+WPZKbNBxFMvGcTyQ8LMU2VkHhBJ+w5jE0rDBCOjgIGSH4ez37vPcwDjo1RiiDT7
kQt1wFqAj+RFZ/AdQgQv0CkEUVxSVMLqm7wVUFryLoNMGV+BmevUk0KMuIs5mHAA
M5xELoWLdoqTelN9waAgAxI25bf7XwSeZFaphKY8wpnvpQqIRQHC+Y1hdKgKI2Dl
p6g4KSna6TDjQMxLZfKm6QLyBsgN62rihQQghTRCZ2BmFM9S7upqGwoM4xrK12Yw
yWuS3YYMj2ciPGKyCaSMCIgfhXXKwdaD99N+IUYvxUPxvjj+zNbztAUis2REXVPs
qPwaEgB7fo93sTV0Q6l4KcaNxerQDdjAlaAgu7Y2KT+ecVEJ5w6tVU0z0tVla0+M
orUsXpBPxUVKE7b5wHd3nBTpQ4HL0gArq+gw7RTRb+NReaxOIB88cYoixZdOvoR7
FlQnEqoUU3dMk6H0X0PRreJq74R0UX9NBMSpZznJKCS5stb5FIrijKt83FPxjl3o
L2sYONIx2fHiHskRUhYl8itf+ZYQbog+QRwsOGuyNdOLGKAMPkFxW+HU6fLFr5yk
c8rRum/iuBVLQNib/mQ/7bcGSfoGBNcVAX49tAhBVCJjezSEia3YD5/+x4znheg3
l9g+hmV3duaZThyp9KonzLDI6cjtsVpKNx8SKGhYHDMyV98tCvp9j69nqfvnW7RG
bFvRQQj001bLVa02w7RwAd3Cs5eMYWe3ssReVQIf/Vaysd9JmDcaFTt73XsKFXPs
0k9hXycxpjeu5JQMv3nIAGjLzlGa56C0eiTinp+9GjVn9V8D4qauuCtE1QWAb467
gjcxy2ti7XZ3FvzcwGyuMf2C9ScC5VxScdO7TrNkLtpaTqVr5ca74fy/JBtGq4+4
skJwULQtRjmXuTZFqockPWiHKWt15uNwk1gIdrJUSHLUHDaA3kdfCf2SmGeaG9hr
HP/GEs1d291lWZgE8X/K600+0wCGa2i9h7QLH07gu6Uc3/fa3eQHhcASAgfcGMb8
Mi8mpEBcowpbkccgR1/oQIPJvT7fUe6uML9Ka+5YCaHy5T2xsBQUUEqf71kA5Xd/
66EZL2Nt+glsfNXW6fjZsQ38mT5wMXGOZNYxh7bwJXzSBY91RZGB5MP1uJyx/voY
MmwOFJjUkIpkT+kBPLlC33y9zCEK2PialnzxEQiU2FO6wKP4XGV5dewjhrwoVJYL
iJCk4RRXgCU3olclE6f/UWcxkXdIsrWfYpClVKhPsLcr8VYOx98QzV7nGpe/hUgk
tqBCaRa0JjGIaPT4JvXcHyIId6y6V99k1dWr9ATvSGlihpx+GYxUyribKywuT0d+
6q5BXlXuO31uYZoKvIePt8ta9PorVUjMfz/fRDNAF7hMnHoHqbVOSKSJ8DLr5hDD
wsmoV/lzGU7oiiihQvfdxHLaQUNxc4UBOumb38zeWUYvf8wWtO0z6a+bH3NafOEJ
E/G1vAJ8fphU0P0GebZkgyiswTFlz4SfAkQyt+ko9A1zEVtIEJ+5mLIL+JYzBb0K
p9Obvyo9apsrILXl4TiTD+M324t3yMejZRVLVC9sFPZFvshI7MUkY1wt4fAgA7Gt
X2N9F5rIIfhXDZtJENbZqpTuO4OzKKDs6gvHZIxU2HJ1hYr7/uYJ/TrGfuy7DEBd
MWFUQF0MMsMPKYT34jwl5vwwdF7eyeqaNibVVlJh132nXQfI8uyQColbPk3I8iAV
IJ8KdjByhFYXvCIyFwVXfs8EOIC5EKTiTzqrNL1H8QpD2Lov4FKEjCE40cSLgCT6
CxOJi5j0neBCt9bBl9WaFG450imJAQCRq6HKB1xQyNrnrD/HVtWw0LWxHsSMQ1iN
2hg2qb4dWGOs9X0Td5KB0kdEUdq3SUTkLcV+uYxrlo2SJvqKAVCvppFWik72OJOR
i0g9s6JFiiaEkJY2NVot6P3ybQFiGW4R78fSLIgEX592bETf3wiPPp2CtuMjOWR5
Gk6g54VSIXVgwc5p6/bEL/FtQunCvpgH93joX1axFz82gmBsfH/pGP7tri7G4eoj
74vi9CJ9SFb9X+PqeUGA3S4ux/JDy6p0tHUrOW6TJggcbf7aulh3+tMmKH4Z1i1K
Ghview0SGf2EorprcDUP4+mFEjj9XiW4pMhiWYHzjCEKCArTIsrBQH+vos6aTcfZ
1pt6XT1CoqwOaVtnsSmbiU+lejxR8rhWX2VCSgYddXpF0Mu271CfPYmhZ5zA556K
nxHjO43ZEagOzr2dq0l7l3OwpjwVmG/jH5zdDNtjeBI8ZQvT8DAgE1ZuKnOrbS05
ePmjRYlauEhHV6+MXHcGW2W+8owJ/w1K+JTwH8nyaT7UYl7bx8tqT3cISWm9nVGx
UWXn8WhF7spw6CpyLVAsCuX/UiN4UijBckbAY1nhBq+jJpsA9tiazlkC1VJ0G9fn
0kQ0ehiVJgxdkP/CdiMHLXikh488mv+15hqn/Hddxu0p5fp2uyYfLOE2DxiaK9Nq
p5P3zZ+Nvab9ZlFMV/vOMFgwHMZ7toeGf1muULZQUX2zLjtKh1fphorXzPafQeH7
cApiH0iwOXCtor9ur0s9i4PZwKNMl6yudklDx++UyoOEC7gF/uKTmmyhEWqwgmWo
eEvsUIrF4hMwmGsqgt7gMQWeY42qP3x5omW/iIQTJzc0cTJGylFC71rt22StxgEU
BX+e9B7OKEJc3pLutpeMns+xUYuW1nF6o0lxkIWx/yJ03eVoamDo+fKwA6Fc99dY
xCRciQPQ0Wnd6t5qXxbMtCVu4Bn/PrkIzx7MdpTLtt5TXrKVNVJgJaVS6mGFg7SN
PW2hLO5FBPWsXTGGb7f9vQqAOlAms2gRbXV/XVikwPCOcJoWjsNdYf/ECy70kduY
OvG+/IgM9C2MXigHi+TVPH0Ujo1m3pvS7GTZmtW0QqalgKvM41EpQeLMpDVuB+zF
d+4i8ImOJkuN0ATqEjUD0fw6+2p3Y56Bwmf3HTlIOOudFiXbNwzc7hnw0CZgjKcs
pg8DGf8Xcjx6l0E5Tujleh+R1WkQaaCdQO5tINgsk0UxUzQMwwRVQm51F74kEcGe
E+fKy3cMBy47SG8LUdipxwqAfDd0l3zdLkEBvBKy/svIRILf7pA5iaqfACQa+B6j
ycOJvoUY+RUneQn+nYTeGR4/poUuuHqSGzvo4U9/kWnQ2Ro1QDAfwSybazhKQl3G
UPJiIklL1AdtLRZj4bDSC3iK+JI/cFtcEHYiJkemW1W68PD/xIq3GPQXoJYwzTAQ
WxpTFtd5L9PoWrc7U4N/yOF1ZK1GDmf5FISf0/rH7bdtUIkY6iHVB6tTJ/1KQWrE
VK20EHOaIRoSdAcOcQWxOh9MvpVAIiJPjpv5LxG7JZY1RlERlFTh91ihX/VeW160
QffPMCFxHpS6neDMOLMN3IBj5nArchNzh4a0NFJH5F0SeedsEHUQs/ttizMlrksE
3HmQBduUwsDgBdUSs2fcSwKrbVpTodh1jWI8Y7k9K3tyBZ2771CGS56ztDrpZXla
dbH0yncMHIgPMVXcg3d/E8mND6bVNY3juAnFut+wWawRgodwrWu9kzdDSqPqzGXI
CPIVRJkM/4PMo7KpkEvymVVz/FWsdBR9mU2UwFzgffuMzpUvlKB7Tz8L6iwQy3Yv
iUEc6k7C5wfDZ2XGy+jsNoz3YDM+WOkyN7OrIOjkCDw1XY57RjOk8kkB/G9emUhv
6VhD9yihHFZbsBk8yvxWtYBR8Ug7tVdXrbYeMu0gGkrRNiISbNUeynbHVf0a7EBs
Uxpkj7b1gS8uDSeWnfmLGA5P3yRCSBF6AdhUo/AGZgArjz+HO6w1IcELYKhq5nxQ
cUdn2DUvwn81sI4TUThiOuJEBW6nGYqKjTcomsprPXJStTuZfNGHGnLUGiTGeZc0
l+CG7gvHUS4YZJ7vaax2cVTj9db3eoGJtpmiwH75e443F6J3Or3XVUy6vY2nLLGG
O8BgEJ4v0XA9y8j2uyQPX719Pmoil5LZYhfG/ZQVbOx4WGkQkaz2Bstf7k2NLWa0
38yb6A1+xq/mkGXyW0HXwfWWx89H0qp3dK9GXXAJWC6N3nuZyYK832M1VfO+wJNV
kEvvTMkF9T8GcYucPbfhKyLesdaG/pEf/Kh8VDAekuiBrujPWcrzQLL4cZ+1ATgw
LyGms9nYqXjVvMlqNWgrMDKzigZXsqr9r5sMAve5z6bvL48feyQJfQbvynE37gKV
v6K4Kvr/NuVLmrqiJwF5pvoLWETqS4yn7MywpwnGmFZiY5mHi4Uc/NNpg0gguSqm
DP2bscJbEgZtKB7lAmzOdFhLb89UCws4ycJH3u8uocLZ6rv2bjTugpSngmdcEdr2
G7xP0hcWcSOdfRAe+H7DcGZyCIWSNyLIsUUIVWHqf/WAagSaX8nKqnDZWHX60JU9
R/V4aQ7dRTof4uw4pJweRBjibMI/U2f/NppKUDz6UYluLSl+jGLUjS/4UDQBDuqQ
WavQ82+My+IviJPj9NyDzhY77FTPEtbksNvkF/TPs8Jw92mlMC7/xP40h9JfAGXb
NqhROUv8+s4lJ2cIMX9FpA19UtFWHbsigCP6SQgNgfrS+xm351ZOi4JtGxhSHZJQ
BpmsSrubdVBe9ta6NpehnvPFQhjMs7nPC7Nudf+TNcFFhLnXio+58/dj2Bi/5z3i
1opOH8Q0enMMUlYWNs3Je5e0/R+y+8QdWevyDNHxeFcOV1uG6Zol7CnR+RgpS6Rs
KOT14hWv0N3TgBEyLygolNg5G77zXF26iW9luYOH6VvnQqXdDP7yYX3hRTNfCJNp
dBWTLvBbuuIaSgpfGkO4kf6cNSjSocm/8+6kxJGXNZorB6KkkS5tX7H9wm4w6dki
Wc+yYtv9GElMmLQNlvd/9CxcNFgE6fB6txqRJzU2n19oHOUQefLs0ocAi2Q7QTbW
OMjkyBidrB+CvJLS1dmCaO4Zr45BWJnhA7G9ZLIkFp13fbiw7c+FlWPBugmvUDN6
xe8dLkLGqYYevaaKE/zVm15W4Vk6yAqx3ymxfa0xQhtWkdZX2TWcVcoD7UlxDMLV
afur8TwTUlt1gXvAra6e1H5STG4Ff2Y7vA34Zc3AdFBJNmbvzuB6fRUUddVCi2Jq
ny7hxDTLi0+l4pdUZNMfnv4kNRydTjNwMk/B1pr3tgWQlCqWhKX9DPznhc0bQy5j
5tY6GE5VLi/43cb8dJy+iZVHK18ef3yi+5l9b6ugfeJno5PqPMJ2ox3wJ9+tdg6c
rUNSo2X1zKT46NpjTQrluLtdGnsQMtciTlhwHwY6Ljps0qeLrbgtLpEeC0ffP8ZY
R+DuvB5zK40UDJVvYpo2GQoIfQ8veM1UnlLIpD5OI8bd6XntyLQYx+cFOus8Tk+7
fFHVYwC1BsM1sjIh/eQ3wZ2e9OTYpakjW0ySiW9fAkbApnq4QSOPZuLC4huyDw8w
HvU/gd32zTf0Mws5GXTCGf85LcQ7FiWfHGOjq3pcGiDut8GVHntuS8wze/wM0NuT
u2GNwKl2eWzwSnoSwu6LBseSZmk+JKmzYD/pYsnkfiaVvkLzMxpN4BXDfH6g0EY/
qZ3r+hZGfwt4lb4CRnnNPuXEbcBHiax1pxYIuMPY92cUzr0ZcisR2xviBWnKrcpl
qWddCxpm5TUlNbSsbmg6Tzns5Bn+HKPPTNtWLQwAtuHmdf2Zy3r1sK6v3u5l1azH
NB6npYhbs4KNR6gVgo4eBzGswjrs/RKcD5m+SqAGuPvG/2Wl/X7lRhAlWGBi6bN/
n3fHl/fj0Tlqt7e7zPz4SS/2KYgEkJed4kuTbFvCtb+ek7wmllDuQL2YlNJQTs+V
DtyaLKXjsrCj9fYcOdgVQT6IBNULvL4tmq1hjAB6MSAY0/yoEKy2x5uERYwT8I40
BjA/+6hlpIQHNwGcQAqQVVD4KeBEiAiHpmjfnqDyaRg/4pKOySSjWEvyytgjTh8k
6xEOteKvpi2JdVfa9QTNrvM8zJNC9fZ9dkAS7QwfpyMi100UAhTcQMYUDcOe2WDH
nBUKum2qwJ/mSkZsWh9dOfwP/zfJFwiEhDBY2FnfQtIwU1wNuapd/VhYnqCPXdJc
1OAiBkoVApiPjNThRGL93XwMGJk49IX23uEBaSWLgJpVd8xyX46bb27RAbnOe3US
K3GydUx+UrNY99NxjMnCi7ZAHyafuk2YR5BrbCnOD33UzSkI5Td3ZwwRY2mJUQPU
VsfOq+w+hZrsyacVoRqvtEOKSARm5oAiLOn/BJ3gbw27954DB35lQB9nHo9uz9kP
C+utp7UJDbBix+aXseOzBm6Ld/PDdCyr+44kZx+CjOtYUXuFIeGxOkraAkvaqsap
KEF/Ug09g9U4jYQaxrRF1lBNRKKHI83tb3sJ/aujtnTA8WukeE4v5/M5/VCpiKcJ
e/q32Q5EVIMwcBr7kcEQmLL6O3udqFBtiMQMlz0/bUkpEKCsRwECZwLuqh2EDQje
GQzZWOgLZjZbtrHPx3boH33Sxi+CS1OTMdpe70AHSKUofwgXlVVRt4ky8Kl+uYxN
w71ks3WsODrKkHRM1ahPy9UxJjNzrsOp6k3797zrxIburJkCcXsKRqT+0QiKx+G6
FMJq2QHokLJCM6dhWneQFUSFgrHxZvvTVyO86pNzwIwflQFwR8I46TgVmYpU3Eny
yFLxd0f35sDXqCq8Ylsvr7b4j4eYEydVOO3DpOwYRWoFCC5ONtoXTg7XeOWhpdJX
Lvhf5UAKSO3t//ogdsr0C9jbuyqx5cSbHV3S2zwROnSPeOe2LLe1aC7wE2NjFJS7
hjnn5FgeAMp3I9X3QF13UEPEVn8O2RUMp944VvWdKPrqeYwoUoAmOl2GCUbqnPeJ
fnbAL8MAQ3B82N3HH43DSsotimpDVLDZE9/o0T6p3NBW9I3n0Ub5Sf8oiz38bdKh
KbSPZdgRtpX6he4KntGvBHBuuhAweX+IeDgFXE1lwbeXGOFfpdcEt/UNheUPtiq2
LucxdVBvB9nrh2oWxHXyTpbMdIzKn+F+1QFgi0ePbQDxatNLyl9c0bnDptFSS+IQ
rYBCGO8CXqd2GpAQ0tLClZzL8Ongv/SQpOZ5B7njaE/qdNIEmLH32cHotMS/S2Hs
0P3uDrT+50EjxO4vKfUw2a8KPV+tt09InbYNxNC0DoqNLQFxxZRa9sfpeq2pdgKO
mdflgoEKhml/nvnGi/3JXG1FUDvlSgNlVB4RYzSuczoSDirDzSntssjvzm7Srfyf
iYOF5NIFYOLzfDsWz2g4H/zFqcvNXCrQfQg8XdZWbwZi00iV+0376C5M0UtA+szo
XXL5l+tbLzZrsiuVAWsv3sAg3kyo3g5jsSRgyytT3L5OzH+8kzMIHhnyYSM3t4NW
60CV/cK0cJL+aMdXXv3avaFC/zVMPIf3HRj0UedXWVK86LC3uLn3uSR4XVinkeOW
ipbJloo7ChUEmUD/7e5jd9TlEeiZVzDAJvJrnDV9n4fmWoTS61WD3xedYBs5chWU
HminyqHEEGpph4HJlP88ar0NEuFjFCTssybnBMFX3+uWcXe3SK5cYtmzoOYHvc5Q
/NY3ISV5dHHLO8vNUpJtALg5VQ96u/YKmP+rYjzJ4xKSFJ7htseInYZfeQ07kGmD
1lWClK7rOMo6Xas10QQ9Esk9g55tOR+WMdlGrV12bF3hnRZKj0cRrlEK9WdutP0d
2suDVufhy6HT+Wt2qMDxXO0i7KSGKllpjPU+4JrbEO3mnjEQ7MGCjyGS4U90Au0r
Y/bKNsntwg1DuFLMQn00AprhOHpUzP/5gXSTgvaj8uV+qj6OB8IpTDxg5BJphx/Q
HCnQ1Vuieu0AVdeY52JvEszhDfqcQ+DtF5aT5ATVieXkWO21bdi0xbB3zmUbOP6b
GiURWSGHZpbhPFx3JgFyayTurUb+hdKHOVnMGskQ4A0TOc7kWerd0W7CBcqmBCMU
loCVPWRxBM9hCXWKEAsLwZnBJB9XE59QN6nIQVubVeXHQ3fTGLou6ItASBqjq3X+
+vXvRNzZYGVTSl1SQ9l5bNSc6C7jaINBJ07ee6+WJVY1gTLNPQ+ab1uJrwjAW2fp
Roy+gIfqTDMlVdn9xqHTof1yR8BdZ3fOi+yM8LpOe4b78L3Yy5tk4qdZJ21PJIy6
m3YMXdzyTOmDHsgAXPhUQ6IGGmdvRi5xOQRDMhBvM5cF7iltDJymwcTdT4Pb3OGB
/qlrECTkOhLWBk3QwY0YVSfyXdWucO9StOwI5Kfj3tcUxEeh/GgZQmW+rS7TARoy
POBQrlZyRP2y0b3iIqK2dh3D0qTiMSLWrX4PFxftkZ8QVpC0VAf8q80VVBE/FIu8
VTrZnX0JBetVWtHcwoFciW1NxIWIPpCoq/AQlSjxSMRvEPpsyY8Sx/g5DausHAeK
NgSQ+hT7u3sSODzhehi2D1wqHPBEWpIsiJg+wluF9HNMRZQNaPplI2LCbMRNKDeR
uewmUll5RIzUvekRZZOJ0agQDH3pt12FAfC7Wha18lX7IbpJbC1wzTKYbvi3dwHt
h0addhQdYkB+E+ppiL0qV5pcvVrs00H8ECfBGNhSlegESRsz2Uisufkz5cZidbDI
rtC5LGmldF3AbixC04Jaqb7N/N+W8OwhJuK/sw0BYKLq4+5//9w/U717wO0URIcL
4+CbBReb6VWHUzrHRH1w6NtiUSM3Pe6tuDeJc3KltQiXDX6n9/OyDF4OEQCULIcr
G1Qas+54JqknC9rbcJNfzSwdRREWBkFEbNaAy5sBuaw8CVMhwNMTV+GJH1tuamFj
5fUk3uvje45FTv2QkdUfZ2CIFDvUPEaHFEZy468gcUBLg3m2YmdaXnVqubjr+61f
dqeVycOmHtmK8R3xAjJo+nj0B4S8IUv5/g2e8XK4zIJ69LVS/lIVtOyM/0DNcvN6
On/4df3qKV3UL7f6ZRGTFbNJPQip0Oyuk+tjuKN9M/ZcE/qEjzYtuIUYxeYoafwZ
+xSAiy3fGjVA7Gw1CdxmHuqO/gJSNXyLFknNRQqh5NvthkivCMb4gGPj7RGG+hxg
Z4qmm9kavPv/4srabG+c+Cuq0QqlYKmG4pr5z8QZz0DQbXeQgqaTxJkEcKjqJxJu
yYoC+KkhS3DCEIJ0WJnknAI8Nwf21pOewx0wHD3MnwnuQWrDb3Uc1VZwLf3HR+iK
30xiEv0k/lLpERG6kWqS/XvoLmsTn4TESv5+qPO5YXCOiWCikDj7iNNHbBUOBAiD
oFEI5LOQ3XB1sjS4N79CYlasmjgOZMq9A8pF2olHxobsQCGdsb7Eopz8rUVnhn7+
vEcmp12eJSzx8KsuuexGzMbmn06o7coa0mH5bkqhFhU2OT241S+jzmxfLKWQz0Os
B7PKQ+lySRU8jbPq5Tt24bJ3SHM7GGiFXu7sYHpNz/nhQKKtrVYjxWkn64B9wK/s
/2jwD7UqZa1QiHa7JBCdWpreXrT9vS2yuPBi76EQrAQ9FpfSMFMZyF84F8hzj1dH
bmDuhKDh7ABhP42Pl51MU2kdFL2NMRsqJeEkRXU/93WLNZ0iE/qRdiYce+3wiJLP
LFlrZlmu9jSUmr76MihUulUeezBl7h2GGMmkCSitCp7yOpiwsaWaheREbDHYgiLQ
dZNKepcS5Z1A7MFTHHVsaBoipRxFr0RQSjd8aZeqn0CVw6E6fwgiFZtM00CqoZD2
reIKM9WdVYK5YLWvTDWB8MqxK558fIBYLpXtUZ36Y3lZzuaQFWi1MYKTiSTTqUcs
/RcgFH+zMyP4jt/k0fuljpTgOh5SwdjR8UNUS00xnjQ1vrV2BhA7EBE8BnQhJIyo
XC1Cs+ixfpJr8vr7wzzE/Ant8LdcAjoNxv0p86lTcATpN2Mex0XZql7dhmnK3PbP
Wmx0TpbvzWNGBtvnSYvq6cJZGgPGYrVurEoMpm4rGnLPtBQgoWseaXa/PKSj+fxt
oFc8Y4nruL0EySE5XF77dcPoLhp3BYEL8HeoU1n6FrNr1ywlPotTA8ZjcLhyRFyH
5kvAgCMve3tgMniAgKTfUIlkorXQYvcYfn7Gohy2JnCsNeuxgfgOBWUrJpqtVU+O
qu4zyuDPuOJEFmNifPh0G6f50y43DeCCHcImFXZ3+ZFmlveN3qH9eTxQYoXXm2QK
IIlAPmXRzIS/cK2Zqtmlbq1WvQ+PM9ZBBdsDE2AXVtaTBe/hnkAy88bbc2QXDVdA
225pMWkZW7cxEK5RmMfQ+HK0Of5x2Xqdbumlmi2nVYn5eVJnEMNFYCbCOGWQmN/h
PeYS8UZ9szhsYXay4maDHdumkSf1qXxIMn0TOi5ZICATy2HRnsk7BAYe1ShZ4xSU
nLtHMpHQp49lCKeYJL6SH1mMKFK/9re9ki4nJXYLQKTO9/WKaXrTEVtnmodxAWNo
SeBm2kWoTMIhCq94MqAivef0N2EILXngzSBUIf6iMNrsfvyXlDEc1BUWdwvxoyI5
3HWOAZZ+vnIaxnXwje850qK+haHTF4DpMVrMCKmF52d8WP+oJgkUzLE80bSzzP+7
mAPN/A/eiM5w9odpxHdUAmr4BNJ6Le4tOmJoXZ2TnHHapzDvZsZEqA3al0VOl/9z
nKeBZzSPiz69v0swz7quamF0PcXv8Y///COqAJG6cN5Wj8tbcJkW0sCVmyALJPCB
YOcDHWgv7WyvwRQmo36s4whDVop8/IM//ytrXZ4C0Sd5hOa9pPwbkqBEpLsSH6JD
6uSwRBZRBeiVyITh2JAd7H4pyOWmcsIR+TJNyKpCoeeX/LUU/aI1CYGSwpV301MP
NLSBiR1yhRitNDXdoYQQfZTpW5sjXwBYSpYaGzWd/z34nQqHBEQ4ELAq/xm0XKha
NHv3gHwAQDJJU8BJ887Fpp4qBiEr0cLXi6wCxyV3d8ocgafq43rpWBdZRBJ92k8l
vrHl8QSNorv8LrSwzsIVfJJKVxJBJriE3dcjV0y9IX+1ldNFFfNvwzlJMbDtICof
o1XGy1r05X0zlrLjUIAEE3QuQlc4EmVP7YxlHpmj5MFcrCSeo458hSHz3x58vBiD
HlTT4dmwvwEsjgjyB50qKVf9R8kTXQiG2ViuPBKR2N/gxXy6FeQSKg2QAUI5oaWx
rXaB+A9o+xInMlXbY6cFhSfBAsqEEs4yeT9UxOnGMkwRFnlMRuZsAE9YyqxHPjkH
AZy7860cYO4WUp5JSL6MI8mgXAf71qZafzDEKBqiFQBxwUw9JSXuZnK+ABbUgPQf
MOzOWQNVkbDVFSUbxrZE9+sPIe1p79JzcWqt4+GumVj4G5u8nmERNXQpb4sGE54O
dvoZbFuTuN2EGCFO1RxhKgi5NPTKjLiRJ6KG9g14Y2tN+stEC2Hfc3NZykVQdK4C
JGEV+lUyIlCTJTkjGUf6MrS6sgrD2KlmSGQrp4O9Cm7sHgaM0IOcUMvV1usfLZsm
2wCFDHE/3T8zijc+2kEml7nFqE6qtweqq0rQulC4U4YAwlJCppGTTZPjav0Uf40n
209O7F+AksyFUtjixbONQPG9hJ1CdvXFkXH8dDe5mZEldtp8RRRYXhcqvmeVzJ9W
Nbqco8IeS+564MkgwCH7pckNpjORyPsmqT0RWrUWMgB5XBUvAMidST6zLTGPIjqF
8OIRnKvo3HE+aCR9hqb4k6JqUPfOnPcMGJfz0LmFQwVJhtFrmICjqcsyLTUGwiXO
PJpsewncbsz3ctZtPes8OJ/UWdxt7qGZzkWWwctfCXETCw2DtgTy9Z+JDiY6RQIJ
WeyjIq+q3pU9JbhVH2yKYVg9MLRChu+7WVRHKcl80S+B+eNesdQgoVKk/MISE0eo
LeYjp4cUEC7CltZVaMl+n5ArmV+TljSn6CtLaFD84PJpCsXUCu7xS2dPniMYxf0Z
YN1KmsLXiRQEn6+WAlJLrbeFdMR+LBknMl0smxvpiqniqJIQ7Ax20hYXO5/LdBKj
rsqWiZdDT69I90PiuFLM5dFw74dnZEZns/PSQnNxwQQX4lSNsqvO5zF3Mq/9uFX8
2+JU58Qz0pCduUyQGhh+xb/3t5tgZng0L4DipS4y1TR0TCGkzXfOBNuxxT0bwE2n
8DLtre++F0NAIZE8ur9z7o0z/LH0A586RO59rUBrYekjTzpYsclkYC1dNvyqJO93
DtZ2Rueyb75YtLAyHnGgQqz+W+00BFNabYFTSWzmHiuei9GSqAvTC7e89WZgg6wg
kpEcEA4cIaBeJfod2Q7Q+KdouHxJNyCOFZgwsyLPpvcvqenZBIER6uNK+DTndplC
+gNXi3b2hzPvV3Q3UmJ1N7HtJkklAk0gBwCfE8Uf83rqjGG0dKB4wvsROA83m0j1
Q6f9k1dzbtI0JFUzXWQei5Rjqur8h3wmw6KysL2jQ/pvr3VIU24KX1FH+4QYnoKb
XoQyZMap4FBx3A3/D4tRj1QbXK3oLXEfDRI9ZRiFGzacJ8nc0SCeJrNTk2zvLX1z
kEKhyF03fGFL7xo4ALSndMvo5cg5CYr0W2fUo2OqHVIpazuxPzYkcTbD+IydVR+n
u5lw9/XyKo2d1fm6wcQtQsCmoo85Ki61w+vLMOYkva5giZD01/Ggi1Fkd5uR+3j9
NMMTASSRME2SKIRgpp1YSYSE0VUlR6+wTXCdmVT7RJ4H38Jl9CBDv7z+AzPMivQs
iFTeIy1Bym8g6DoqCpjjT7+3r85HZt+Ig5/hbHja4HY4bD+NmvvHG4iuqVbNpdvU
ZaSV88f7jviRpCG8t3cVGeEpj9ge5LIv6pWQlAt8U/d0d9vU8QwqAN+3zt4DrsWW
P0EbrzOx4+FHZmsHonOdkKZFUpsUxOlVVu1k5EKGkABcTe1BqUAdtcGoboWFWVPL
PF0Z9aicGoD09o4zuiY69+Yw+LmVq1o//EVB6v13kuzK7d17y9NsKJiyKYaxSRIm
/u5IfNCSGiAjc148gyq9WoBWIZY7LCIYdzLwb8TDqBk6ucXNyDMyke+sL6yLcyJB
mhlsUeWOJ/MzyuN22cX1Vpmz0N3PobydV6geOaPbcj0q6OPjjJppLX2fjvxaTcDt
ONFghSd5M4DpmqiTCr8gyFpqPPR6My0WtfM/kVMdPzVwfqOyct/sDXXV1hypp5ua
kHY0EwnmzfWDPb3Aiu+Km+f+RAbB6wsZAsju/8li6TzT/P0H6IZQEWbGH+WiJQDu
pI6rZc6/3ui8bUASO0KHz/KIejoAlRBH570Rg7Hcj7JPrvS4g2T2TWm6qvycXaOg
/Fs4sCLwkL/CszF2uWlRRAiqgXAvo1Cfy94VD1v1n4SZpBjZ+AZLz6o27HdP7kzH
woBcJ63P+VTQkOEXQ8tsu0+lKvShRtNOvWpvQ6S6wXovO58osVsJjFBjeW2IOXT5
1glh/gqkYxYmGTBcyI+xGjJs/n92Fy/dm7MT3bRfGGwXS8U3DnMNKx2JXevH500e
IuQgynqoS5BJ5cfvBNeosPSqJs/Xab5LUdJCqN3TGZWslJ7SKJ6x4iG0UEmPxHcT
fhBCMumOCARU1c6q2WCe7IK78yeLNdbWwdRCu8WG5pbc9tMT+0/lx6kUz7HKX6D8
p19cof1j87JuvZ5Svn1jU2NT/0oJsLRO+H05rkEiirZd6ks/8CiMvGf4fZ2SdwO6
hfDjuWhoGeFJWHWKEe2YXtOuPOosNWfdmicfMjmWLo8XpICQpytGzpb8qjOCDMfS
ko7TcYb1nqdgMQpRZav/GuPcIA36RXGkrTTYOSKZPX0Q/VfXVpSa+En55DDdMK8c
qH9VTCoib7YZBJJLXl3Rt8e/bzCwy5VwFTUKiSzWPwiGv5X2IOP60eaYcI3V7OE/
wXxwEtghMlFzXfFFTdy3ER0stt0N5m3zt8z8Kk2UCLoaDTZE6Isr635Nhwq41IC3
C+e2E1d58dnJyCKLOfO3FOGN1QF4k9tsnwkCNeYaraWeZD2RyTHJQj8qQETnXv2h
I8ukTKJ6d4Ck2i9Izkf1O5zb+BDsQKI3EUGjPM2+uq1z6ujoHO94uVoVbIfo6Qvi
LAVqes2xMC3ir857iI3OlGCU2N/n7EwYjyok+h7ajQnu5br+y78Vq378p9iHBDW1
hFt4T1UTugNgv8PcmGmObshQpvijHOsVvCHUUZmzfo5M8/aJe/D0N0pq4kvW83B8
rb1GdVOj7Y8tppbm2Qg9gPxFJrZYc7OCDoNOomrVZJYn24M+bXDTl7mhAeO3YytY
oDIjvAY2c5ilkmCQYM9KuqEZbFVHDXnEjZIROKGyiUhsfApZ1aZfEy4nStGbULHG
1o/5ru2jJmIPuBxQh89F2fzX5GiF5Zf+suZBMC6iwEyX4Q4TkRE0pKne0bB7Walc
GpF70feYsa3Dvri4GidPi9D6uXKmTLCVf8r5Pfj9Plb2LhWtNh4N+LsL84V4p7Gd
YU4BaAkdo8KrMuQl4hns+6lhdisUMFngQPpCfAQZFdISR/UPtKRPxC9XaUS19qZ/
3ek00hdowQe9Iu5zFcdeOKiT5WGdCzJWuGRLeO0tLO/5c8Kn9V3PhrzrBjp+QVNY
8ooZUylCk/eNFOgerYGttKGZqXiztSrXPrcF2NrKwNR4dLTQBw4ygWgXIftz+edQ
pqEx5gyeEuhD1B80KsYnOE9eQS1CycNnMmk721DnHoI1tsalmgZrLwt5km9i5h8C
ibB44PURuOGkjCK5v3G5Of80HowsQstAzV3wmF23SgOpcnqt0KE7lN+F+GeYaTx+
tJRyry6ZB1s40tNdyeL3JWfdldyi95ckGYmkv7UVMbRmk+oRLYTKQQhaX+dqJq/Y
DoAut4UCOfEloA5DIk9HDS6jlCgvjFn/5w3lACPNovqCoiMJF5ZzPlnVrs7clI3y
V3csazmf0735dBzbAzkfVDNz74ADc8OwPc8xboC8gIFfoL4uduV84lfDLNR2lDPX
J7tU/5ubNqlBvpZ3BzpChKxziftTlUeDuTxveTSO2rgGkqo+q0aLU9yz+xneZ3I7
4V1wWMHCuL1yetwtNqim3NojyCXXN/dGFUF+Svd905jZL39EfE9J9i895kdT7bXU
zA9AipBCi0Az/h/QBInfVNXga+FSF/UYRNPVhMoQUUZXkkys7y+r1GZ7lZ4Bkdwu
fy8q8kW/D07NFTY2PHQhlPoiiBZVM4vvIbqMKbAWq2zOBN0M+L4nUS4JaVPqWc4E
AILa4xmoUSz1n3VXIeyOyPGLxtximP9hxtQFP06cllIdDbiinZXVxHmpyWuVYPIq
3yswKKTidF9aU3LdwXjNkjNDIVcMO/WFOea50b2GXD5ZWsHMwUOjQrCG8vGnl0c8
+4BEI2iAMMKwS0VS6gPKm/m4MCMv05g7MVfo6JMlXV5uM5tPzduD69ez/teArEjU
PkJoh2q4WATrTP8AfmJD8tQHWQ4m9ii66ZETQWsYLvKS9D6ADW6OGSomME7/7m9y
fN3aGqFtKprMrLKWVNlSkxPOgKaqq7QUl3C4srEyclExrmoCkjo3CMCcNwPSOwyg
/5SV+evf47xSH5G6fULS20yBLwNy1NiZ0XOWB/SKqM2PcCarphCrcSBzS/HTp52+
JD1U4XM4DB66MHyW4mqq2RH0y4g2LVrRI1xKFS8PVWqPEVth0fFIzpIZT3JgwS9r
6RcjhgLmMnhJHwJyQ7QJHxHt/HK0imp2cE4m31eeeIiAPqebibXXaz+Q5gnv5rba
ADuEFhx8E5+SPMfCUY1vbSlV/qJ8hCqOQlYEoD7ekGHAKDbIRJO0R+mEI2/rbtKm
7OOCSqyIpK/rNYJj6pahHQ9QBBQDFrJKHMTDzt5QYr77+IilobkhE+ZHQqt9g9GA
k4ZOCHxc58SFQ7A0whJp7IuUPXibc3Z5uH8zyvJlvvfW/QEMetboDNeBDA2t/V9L
9qXF1pJEkdnw7IYX2sHpKIIEioU4MD/JlDKrNb21h8PTIasil4X87GhYRB5tX9Ot
ovrX70263Kv4sY6t7kFNdmhpSmA4K1F/g3UidAQkZaNH/bFnDuJC9VI1u5i3SnRD
JJpnfctdJC1CHrMg/Ca8s0VltUdJ0JeOy1mUCC5SH1LVJ0r5tuqUk2fkv7AHCtyE
QKWquYvu+9polAjJpjgVY1aIDI6bZvchrGJTKN1jPtnsycRj/gZiEQaS0iI9f7y6
/bffB4+Y2PQLlvzVFzD31axWCDsH/kMPx4Ehfp0akgf+IjmkvZE4f/CvpOWRJu2k
nBktbqkce2ny5/tKB6UF7ko+Ex2EsIhRdvTlctqOhtnPuvorAJfQBZcXXSHQ7oMi
HWlQD5O5O8nEH/cnRUQbEq9SHxiQtdnd/aAmb0Rfc4qNoOSBKUS2+LXuohSdEkVA
l8afB+7v6XzaxqZYkRwzNDBoX44etYdjV9DngzAfJNf2Il2OqIlbMMW1fRCBy+W7
l72pvnbaom7Sm4kG+jOyJ/ZU6pEhjszdHkcMFq6y/in6F9Zlx1+kk4lcdo7+yP/7
BcW4T+4seP1r3DjHgdo3SaLbFjePW0yvRXIOnKEyNyt55XASAOXyZ0zG8UMVykVF
TB0DHzlgvJjpj23b8cOQZG7w2mmhMu+sN31n0eMfQTu9FP67/HFygZaDXF5i2eA/
9dyqIjcNd9JPsI2p4JPknYOcscBgwTtOfIJK6xXxHwZZZKW6xV7gHliHs5q2wpnB
envhIp/JBDEvHiyrgVXVfYjiutUpWKl7qaUEN7xJMQ4TVqcbA+ixWu3nbbKfEFfl
unZpIrzgu7bDyPs0sW85l8Xcy30ocA4GCRmajHKs6wa+BH5IQEsgJIb9KpSbgWjx
ZvnP7JOvd7ixeGypq+hPnHKndDf2WmkNOyvpke3ByCcEmSt30m8SQ1aU1JcMAo9i
I0nvfmdFd5RUUSvGGrABOlkiZZZivs1qWsqYeJJLPIiCKVdJruMpnmvp2WMnLcks
DFbkg/tmdzGlRPVzcrUI9+VAzfoXpHIl+zLyjmpklrvagl3gp2i+O3+XDBfmO3V8
N1AJ6db8VbVhhZWUBJWkMXOlWHL2/zt83pT4bMvAjOANw7TpF5SJcIYi4zDJ+BZ7
upVXLthrt2tvtaLxaLdc0KIaqGUqZbMUAFyiPDOwby0Q0As1DcNijRLZnXySx18l
WmWtfqYH6uU5Id/zd1jLiCtkb1mg61ZoZ93vuxwytMYQvQWRjrtWnWZ7EviaziHU
34BETsqNI3bmrmP0CswZOBqzjtUD80B/vsgwVVTIJbnopSkHxU9Dzrzw6EgZon00
7p4SZdR6Z0fYK8KPAEbevxRI9CCPbw+wU0qD2L3GZkzBbS0qDFP5n1zKasf7ahFs
mJEr4Euydznoyf7SQmZ4334GKiUzmuGwoa5JC+AYed6XLcJNlqAKWpTHrqHROwna
47FhHnOF1Utz3pQqxLPN/LcTFSl9s3/qg/Tw9yVxLKq0vyM4RLOa4LtgP9TevNhJ
u3Zg2pq4e3RdgZoj+7j17GbLovrFFystdnQN+B6hLDrLVuBjwbZbxSLnSBMjYAWX
mim66ccYa6Txrpb1Apryv1I+J/Lug+acftpV9KEQKtTJF+WjqbYHhxCwUbKjgZ9+
X7Dbsiy7EtMyIh0TTGh+Y7qPAujfsfyDpotFrK/uphhobwNcu4x6ZIPhGWzi/2lD
Q3V6wRdKCVOZ2fP496CqdM9qe4BASDuUXoYSF/461kcFi51Bw+RofUhkU0gGayqa
ftUqvMbgOBb3wmElCBoMMvVj4UN7Kq0GPeSjSAeb4knEiLR3zGXbPepWW0u1YRyA
A0Mt/QyYOeQbIit33K8MvD0RAh8SMA36pmRkNbFiXaq/wPW00vR4tYDVfFLKFhzw
YOn/kj1yxSPCQro8bvqC+StG45QhBxSF+b+XlOeINsiXz9Mk/bBRsoQ0DDNIUB/Q
AGoElpue8Rzjwxf+kdTidFhQpb8RJuHrrCo2VZdjCCVte0Q3Wc4YPqMvcrSzh3Pq
XCOf8rlIzICuPFG6XwEsPB+9XrWR9Kc+q3g2D70lkR6lfpLututWdDxOdgA2NBt7
rE6I4ieEeCbQljdrcAHsf3x7y8ozyNE+fNH1zdEwXSdYqHOohVqK1jqCkJDNfjcX
gUN2msp/mYM9y40SDGgP6c1jT6o1eh55UW/3Y1rqDvcgGQ2N7c+SsmZZCpqTnJ1P
aUzLftB7ac49+7NycTnr8a3xC3WzWNw6G7reVv2odTeUt/3kHgK10YSnycMRRVqS
QkhSXaxed1FasBGap7QZIju3GiM59mQtFO2RQ3ofzfBftuBivbK8HMpUxxbOti7R
bigQHLoduTvGG+HJutufez4FirI9S9o4WH66tgXph1ltd8Yk2+apF6KghhSl3zdu
8Gb19z2ryEMsnwW2oJ6+jFt9/WI3yLp4TOvzmaPN6pMHtDbfbdLND6pjWmgapjQ3
IMefLp0duRdpB6X1Rks3ELlZPNaEez/iWQy7dAc4TpP+xJfsDEdWKGxkEuhQdTpt
6+xyYvrDNT7VNoF7I2U/GbjESg84in9tCF9wkrYkm4/7ikOj0DoNGuUa10tGtiRp
SBrMGE9PyoCxdGRhzXE0I5gCCPgXo4GTLMqg84QPQP5pKJyxjI/OTLXYA6g1dKay
Y/vE0tgz6JebLur/bfXOwscaX75rYU2CzUeFAapEmJIdjCwJA/opzB92HobWzAys
WRjITcE+/PsxorkF/Il5h1+6tINkLId5Lbdsx/GZ1J9hiGeZDE5LNH8JlxhFLlWz
e6z+FLB5UdGsW05bULaNeONzPZ4YXo/oHpFUlKjcDXDQrZIT0QoQ2pQQm/7vGfgG
vgdMV2Rit28LJMz/bmkILdKLsQIMNJHUDaLZVuUkBLVN2inZ9/RkfEJUyRQm2C7X
qekKAYB+PM5jQptBJLvjuz9KeBsVEsE/0+D8c0QHMkO/g1Z8CI/RgKhALgjtQgw0
9IEHVWZImjECdE6ZGNmkeC1JfhEZkVICxKKwlFURbXF5yyukuzEvurSld4ExlDbU
hBMJa+zoMk7Y1e2KOfPFtBdyvEHis44xGOujQZ/yJlC3UnTOz0b/On5y3OzN1Nmv
eaS+zTz98/jlQwciIN1sSmwfb4RKYq+k0GysZSqjXfJWLlKGrVK4KeN7aa0+V5qp
97470ueYIgdWQvi/s/p/F65ejQs7d4lT6aXS/AQRka0Sszb4rHSyaB9TgYU7DDeD
W/EftSmYiJJwgd+oQgQ+sG1apFuVBJ2sy1Bf//mesMxIKIOLBltWdnt4+lDe3oEp
CFWdPKIONdAebFwfIzGiY/t1Rq6noG0vKxuEFTJr93PAmixxWWBfl6bw8lEW5RFR
+Q0fJKbHZ+9+oStubctUAIuYWyFC9449pg7nh0qEscxw0Vp4YLvf/oum7a98cOkm
QeqD83hl7qQS28d3y3oyi+PxmAalWGVsxOMTRjut8zaAxS3fqk5qILEZVEhkpmWD
3M/iBSeEbWwzRBrnVenLzTRYx+bEtVvL6RbhiKBp1xzeW0gFaPEV4Ajra6uzebCH
Yb29LlBYLKqzpxpf4X8vTNQBh9esPPvnOFXbAa5cuo3k7DRd+yCLVdxp7JFoKCbd
/TxD6uq1wHLqMAnhOqOvcJG/H8235ivAhzOiwgDpzcxjtz2ZIcag1SqzVAxsimkN
ZbH7vZKkn9gCaSV2NgNuBLnU1twUmgrn0SHq9zJ5uhYq67oSXvgpNJi08iPQTk9l
4Mo4ourS2t9zV0uVRMcPrlgyTN/D2mf+csudOlJb9Yi8+M+yYoKKUem9olv1yGEw
/wuKchELQbtD7UpZnIFMwPUPQW0dJPSkGFKxE42dWBvRfic0NZxC107Jquz/ZiPw
8pGMnNzwfRcdb3gvMQISyVvkPzcN1CXHqJQZS50r85BeDX/HwEAdwLTQZqQ4430t
nVTBbkMGrVjP47E4pplUbUIJ9pzG4A6Wrs2WKgZnYbIXo/MhFlnD/Kab19lIadlI
l48MvMqSnZBKcuylCdQbTkigvYheVEk3IkfKUWESoUbiXyixVeUJ1GrX5mMft9rd
v7Ph3H/iPsyVWw6bf1o6k1B6X3AirJkug+30sx328IIITt9PE0HUDuyMbakuC6WN
4K71x/xN0AWJ+CGbG1oeaBjDHhjtgSTtcu+SyXjxmB72v/XwZs0l3fji0haVd6Wq
RahDCkpopq7URDIEeAomVhQ1P+3FL0Ihvz2tHdnkYHvz7wwH8qZeZRc9tdb+3rzG
Zdq3LcZGV6wNLY38izlBioXpL+q5YIyH44ZbVwaNh+idS9vIguMvrbvAL6awydgO
rygGuroK+pXxV8WAZKvLvdCp/GNJWE1VxzLkx/0rLFQMk25GL544PpsicEaYyjTA
WUI8icc2yNtTLWV93s1Ns9XxP2ZddDfZG+yK2RgwxyANXWM0er3ltTOtGKVFlgXa
PEzcBTLDVTPIsCKAZut+SbLV4b4BmjTPDhjuZyvHUe/IBE8ZvN71kjfpLLbZgYNh
XcWJJO74PnraogAO9BRumAQzjbgUr7CHQsgW9b4ZP3UFp5v50F5NtsFMxwxg/h1y
EUtAHLzir73BjJzYEhG/eS1AKIFNKtbXJxDelZDECp1SjWXIAZ5T48iiVsHjAbHB
CBPtSKhQ359cyiW7sSmhw7hoNbmyzVlzxFrD7BKoGxNwUt2ejEJc6vztgnA2eU54
i5jbdUeIm22BMO58ab3Xy455vs1q92FhAO6hlKdWzwbblu0xJcz5T/4/taAYM6GL
8oiyXYxPZqHbgNstsqR+YprX/AtHpiRGecyly0B+pOZGtO8qVzWoJL1QFQMu/S/i
I+ZRPDmH0LadK0WTkjIxS3pxqWsRDLbvte7Acgowcd10tsZRv1NzCOAqg9WiUA1Z
ZZ2jEsl0l8g3XRv2Dw0twhqFuUZdUA+uC2rqU6+pp0D0uvt8/FNCYVw7PDaTg3Zp
wR9WK3PHGD83QGUV9o2TYPHo79gjmagQ+pLNjlUkkq2jV6ZV9txaz1dMRSpvnc84
juluK7Vv1zJcf+A6i8itGvF77ZWehAnwmut8hFcd9xua+IwZGSBw5QNZSu3+6li9
4IdmGoHjNgCaZEI87WtN66w+MKt7SXJhiMf/7pt8yKqkn9pblx4WCLL80elGc83v
rl8jIqX4xkd6vh64nTOxmqxRxWyrWJ+qB1Kkfvf0/Eg64XcdqVDeRBHORxQT6Vt+
2rqTvJX7U+teX5ILsNuXk8GF4mA2mQfAvrGTkBGRRhpvhCVyfQX/WXxSUID6JmLO
pyzqzO+39R4QMV3JhfJz86qns5CmBOoKslwtVO0GKNM90gZpR1Q29i3U9W+kVMVL
dkiu8pXBu/us82r11WYIswipdRc2T5xHufG4mauF/25aXmloX9c1+2ceZhMQ1Npx
v9w8p72sk1675WogcQa+BH4v3j9++g7knGUxFidUKznBs+nCSivr2MhzF6vyp858
JGW6nezWUK5Qn4VKp4IWOFtOiVvY3gJHivQqwhgtEJsDufpSQkyG5N6yJ46R/l06
36ob/uaMNf5BMLyOW7QqfKsR6qvLb63vrFKoXYxPl+Ea6/LYYFEj0Sp9xMO0m9Op
ce8r1TFo/02KIMciTx/gWwlXZ8hb6PXjWDgcWY1VT/61H1jiwiN0w3VxsLbU1U73
hhKLapNv/AlWxIDLowAw+ylOVyyWdm8GjwmtN/n9PiBIX1yRzMmnvE+WRYhpPFgz
mwRhgj6xiYglTa5C2z8oQd9iG/4dRTgNSXph8G0vz9eqj1m7iMIFOOQHV2MGnHkW
KftpKoznvzWMHTW+kX9Gi3YhQTs7Z8pnmziNhYe1/977+GjvWxm6hItDjSP0MUDE
jxxg+b5sW49y8MBw4AOEKQhKB5Ye6q2xheoLUJw69EAJazc/InOJUMYZMUeofCai
2il5T8/zQvaA79rAW0WTMbj9/mooLPbniVR5ntSTu5ToVjcD12Vo/JTQucJXbrft
xhZ7K+U31dcUE/uFFzhpngAz/w1KnC7nM8V+YPlOpYeuzUCg+1IoyQQXlXSmY/j/
M4yZfqCXHYOnOgog8XgHK1+CUi27LFw1Cb2X6T90wBJB/zWISp4PZONeLOmXc3id
DLWFhL5EWo2EXq63qQih6cMQbxrWK21mj2Bqw09X0G18vB8G9TTfqTV+ICCiJWsh
+7ShaKjZ4S9mhppEMh+4jNr2yuKLV8s5GKrP5ugx2e0acEl0opTmy7h7UuQfWwuS
UgylhfgFp7TcXkY7lXdZba2hd1mJJoXFc+pd69XFWSpAH3sXSjAPcgqSlzc+bFDe
QPLR3Gg6ZGfUaw6EVU8alaERcVHdDRQ6gnufBWGeCnqYGIJ0wSdSDtMpMmi/CRpD
EVGX/9f9braErKdXaJqWsF3mukCWkzcR0cznKDS0w+lvCOIHEDcqELpKWsZKJ8Ek
IbtwICluWwdLi7gBbrgiwlv12IwAu9nT7ZbxvflrhLvW6rMyUdt4McLmm8+ZGZZR
jmMuHeXCY4shUC1eT8fBRN4yaG6iloM6qbN3k3rVREzMfxJaFuk26WjNScUejoaD
BMX+9CKQmhEM4iywLPXR8Rk437Ar2X8kVDyB0mW6NR8AbQ8HRMA0QAddtvd49uLt
X1vTalX14KtJPGq93U+e2GUnp5psXxzOxpjxdV5v/HwUfrX+fSNDx/ATYPFmAhyQ
bnwh5JgTC2HwP2rO//RbqXT2CyenJyufrTzGNdJ7pZe6I9INE3SzWSDm48xlMsIC
9UK691B0+lh4RxX6WM4nkAmoci/XC+10R2KWobs8ABoFr+ty443J4f/SVbt2Pdby
5i8Y1hNXghaG3/5rKmBM7xtN4WSN4bvZutGppOIOuKjNZZDDwAvbUFu5A/TJ3CSK
oicX089UtOQhlQMcvIG4L4f4U3mL6d6qi5KJdEta2ZTPAVccc5/GzvU/ZEhB5X/5
xUKi+Idlvx/1F1gzLgBAWAImCC1zpm5dNKKf/MG54BcuEBYcP2JshUEafXS7OPhw
1M5gxj6wsVpNCB6kO2vEOCEUxpw92fAswjtoqUOrERdN2qjppcpD+c0pwOmvVAv/
r6pdDVuDKMd3Y1xgRUtfhxjEfSVjo2qLUVlZwvxgnuI8pLPQP2U5OBFtwjQPDiig
xNtY0ZZH2rGtwiKdlkpyhvwL504HT//sbTolib2oFH3tLghd6P5xWfc5YgHA7wKP
G6QRSxuMCoEYjfzEnD+bUftyFePsbUGj/N8bL0bDupLdVxjD1VSVmGbKD3nCWcFY
IPpCd0im80n+qcr8ovJW3WT0aLAtjtebKml3lEilwAGGM/gdDfr2JSCItEG44RjC
Lmtg89vSFFfoCLb7PjmskyRpXymBsUVnTP05WJu6wIvB4g1HcNmQp8J0UZTPCAO3
378tgaKTrGK2R10Td8oShHI2dSQ8txh+0FTpmd6UYwyFKShZE2fpk2u1oLGx6PZy
iS/a25wQkvmXr8ij1hqjGYO3mmSsLJWcW2C7v0NuR4Jk4fhuzy75gnKt6vhqLHrj
gaHOr8S8S/FDJKYcTn24JzTQiOtd4fwglNcde50xoiKpTh/dUncP2lRgHMTpyUPN
AYT1PqoZTousGIkOqHn5TWXqEkTXmcGhMnrlmqbuvc0ZU1rserFBdtqaO/G8zz6t
gog207AS9tlUHKFrVRw2q0DG3XgBZ00DDFIh2oTgZQ3pCh4ye3g+/ujwjb9Oc9Sd
zE5eaCpxH2JD1NM7XNAapARCyXyPRM1FStPyQXkmj0BdhzdYrrazHB2cOpG+ls3G
6GD5e59sV4XBlLAFvwx6Ss9xVf9+nXjPwbjxG4ftc7fuo/m+ZkPUki/GtzlQx+B3
h1qgCScpXZ7Sv0jTzVTnCgcxyRyGwLIdPxB1yfd2MpI+mYgZSFDPCHuvDKYFHNmQ
gpz0iXh8ByGUFPW9LZFkbGen4iQrGndnwcnRAa18N6yq2ZYKLcJ2Ql3KnwYjzlsa
h6GvzD9PBzeRvn3s3dRpfJ2iwm2w3TDvLFq8RpUyMyat/2kpkbClokUrFmD/gVxO
nr5TT5xJIwMuL9V4baTBFRPCgEo7Ot8LxiwPmCojyTFLE/3DnpwAldt3TC1snius
U7+c8bnCUryZFTlp23bJwNJIZDrhCOY9ig6KW5BEgoAh9Lh1okwZ6Ye0aw8lDSoC
g4uOmeANBfIQDLvzwu/bwTw4hxRjjGjAixZskiZz+gqXmKjjYiyCrmIyMMojOIew
twXSAY6P1csQBkNqf/aeO1MyFFgl9JDNpuuioDMsL2ukLOfhNMJEB0aOFAgn4V5a
xGKuIGNZxPPBt+TfGA72OHaPpQDpNuNX3o0yt3Atx3CIDDYLyCt1ybZnki2yAMwu
c/bpVgHgmEPGPVj2SS/kIOHRM8/Xj4lCjIcOj/iDtOi/jOesnNaquyrQs3ZO3ILH
yocNPn77PFGRxdVf9ONxTEWDdxEQ3ZxCkuovNPym32Q/cuwpwgmrMgMZrLNI/H/P
rsjxnEOeWi4Laj9UvO644M1aniqfdVaWiSFj1XW2x3ONxch7m0wJXkFRLOjglpIG
dHRfxw+hSeG+kJc7pBtusfJc3ANxFTVgftaqfyVK7oKOuI/3K5KTQAg5qO3oNC34
eIH9rqL6fl+LjjKDyxNBWBNLbdB5xRAQSLND99JHY/b+WCR7sKCIx+g9rlgz3yKT
4Zmi8OOsVu0zzXe0Tc8Okd+OwQPjpscB5yRAOEdVsUC6sbe84FQDapaNrIn4GGRK
8/Y1Wki/S9dn5l/jsVx4YBHsBTaqjl3iaxBz9aNPhpomcdeUwRpvF7josI3LFvY8
ijuN8WZz3cYkQgHA1S9ogUspfaF1yiH8JqY38tgfJDhb7Oara15t6KjBo8UgJSJ7
O5i4dEFAun3qqW6Cv1BptVjjJjHP8OrLOLeh1lork9P3zzGudKAIDBeYBYGhPr9q
dsW9u8leogWfsdsFLvDEBAnPBVBA0vmlec7nMFamR2RifecC5VQo9mGtqyI/vnab
wH8gYnbzvIt2PxGXpILrecnr0HKwXPlMia22hlkypSksvAjA9vO9qXgyM7FbTR2R
vZP5cKsKsg8HyIV7PskLexKpcYJ/fxagYhfpvC1r64jqy8n5gULNfGDzidEVJfNP
HL8jvxruL7aDLaOJCSlnKM1CrrXkf7WpT9m95RXif0dlg415LlpvB/LzR+FQCPze
18IMGXg17NEvSOpmMp1jYjF9xsHpoWD465RbzDebMU1OsqOKriYr0OvhBpuX6jKt
6PGenmcsKZMK5iNSeFGGe7RfGPP+uQdbpxkrkZoGCv8s6abOFCCqQcknbVka0mtv
j01gQfUvlz0s7SE6IFNZCABuqUgeBBvI5c/kLHuFvxndHuDRkAO65qmcjEHrf0KU
IiWh18FfL3asV9Vhgu6tp83g3P3jMkKFYJuxmhkHESIuJaf9NikBpMn6o1D1iF0l
Y7bpYg7R4+vPxQ5Mj2FbomeyjFaIDqsAUywq+mitC6Fx6063voOooEBn8uQP4yS/
1lYAfh4KZ7lCdC/k+YZHhveA68/qVYsg84JsfeeqS/PY10KpwhncYmF0rbZOlWMt
ZT+sJ0A7DOGZhqmvb+XCJ1tiG06lbTvIO+vRxyQgul3IjlsAK4PoIHrTx5X+uvCb
gPNPpag7nlsuorE3EeExKPSD7WWi+miA5Dy8F5jP6WZQcf9UGtUMV3jNdvZdRNF+
`protect end_protected