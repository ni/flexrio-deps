`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7184 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0gQgIG1mJzulW1XOK5NnZR8
C8XqDUtXW7uOWTnSVqbIblwOHrDC/GFb3kYl7b/cVSTt2SIQ7dTzgS/uSzsHBXGr
hyG/X7X4a3b0gDMNg315SZ07O822nXR6Ah+fVeuDLhaNdP2GsuIii25Mn/mMShEd
iwCzhYXbZARFyr1TGkLp785VNht2lQ6STKzbMps7RcK+xf+calOKlPpdNaj6DwbW
OSCIbHrxi3r0wPFEx/1LH4YcrkAZdRelkZkgPsz7TU5TH6hiW9zaqY9fT4GZOOf5
e3J/PqVkvxm6veIy3ENj0svTrkk6x9oDwvud9RsbfGFxGbWbRHYlQRhYpBq/FhdY
rRp2P7kNmEeCzxYgR3+4YU9nzui1PfJsNWv7mY0MLMqicwo9W+FSSThYIZlNMyiE
034GomDcOrqfiRDYlcGMl4ug0jCfDlr/pK9XZN2S1LzuqWCz8TRY/qShltZrgrL6
DT1IYO9fwZrehVgI1HWIKgugcOyMOLeOUFxd+zqMpIemmkLBrxjNVDw6aTH9q7Dd
e6iFOeu3uLk98CyHEAimIBEaokG780tdH3/wCrIjfXX3MbGFMz46Mbraejsp+cwp
qWxDwMEPibHR1Id49LWeLRGa59ffaYAqW1jJhO8KG9VGRKoVcGsJwxzMjR8IgVBt
8By/UyaHREA8KbXIa8dukGZC0PGXc+anO/p9ALyShoJIUqu7zkMPpxPhCz4vYjJN
gkEWyjcGje3O4Fx2nrUmeeNqE85A9rdRENzNubjTeyAADqOazMdECN0dng37cdfp
nkc5SfYL3rF05k7V+DSRxsMWbvMKJk+wx61ke2d4HieKm/SHQCBEW9Fe7t+aWDB0
tde2uoQzKYsqs70UnhHhkovW9TFwP6Le3ukmQNAbW0VKAT2CQFRnj7oiD8vcEqCD
iCVV2d2llESBwDY3fig1PHSlY8aiJNuU0IOt/w/qPAR3/P8hdZmLz9GX86rEOdzb
HMQzRSKgpnh1AXPCvtN8EltFWvNN3M2pYCtUnOQrTWX6UZ316RZzxpoaCJrWhstL
h8VmSCEqrPJ33JbD3oYp8vcLZjMww0w2ogihvLU2qMUeW7r6kYQ/bgPBKRaXeXJ3
orP79QAnbZHZnp6PGrce72MSc0dSe/17vKvwUT5c4g18ICt93KFSQLFDAjLD0PfE
7DSSmFcS9VB77tAY2+0tQeKtom0CK805vJyYlTe/z+Jm/lK8wcZvvX9dDD4UNxFh
xaRmG4GjfDZEXcAmIVtlTC7pLdi1+VMuLccsICo3E0J44fvXBZEgsqFQrKZMRTwb
W74QSbJzm7JgTuYEWbDSOGTNf8/fVruH7BJI5fSPtHiyIvo3wXH4MObhU3UnQzgx
jVnwdal2oeH3Tbs/BWNISf0R1/ka9GMj74wmG3ZYzTezUNwdZDF8C5f78vvtLCer
i+LcB78UUKG954nFX8NCjS01JJ8NKYaCC7vhA0sNWdVnbnPktJpq2heoOexX7OWW
wXoTkC+HCnFvyMdUjc3iYbaN23Pf5Az2TbxMGSCCEXBnSLR3xnxGVCHQm4vPTlaZ
oqZmKM1OsGWTCZG5AZM7bmCsLaQ6fd9nd6FPbTPL0meCBUdlygAPnrCTmMDCniCE
x/6AMUFZw3qsEyOj0rwyor+/ewxbIX9gwHd4LSuzscNX0P96clBy4SwB9H7zhFMK
lyl852ZJ79VCi7w6e/iEeu/2tvSd8upWIY0LlXEFdVWTKDHRwSyXc6FEVF/n+fGp
MGj/B9L1D+WTvw4WPrwd7QMyUanciB/7h51oKeaqq+tFIhkavW+RQiE0g5dy7DYK
mkWFcwpsja/slkhI+Q+AD4/iEltBAIx/nOxT/DeXv0oERAHW2agg0YrCh3yvkVMj
QJtheYs+hGxsvn5DOvzxAHLA3pYh97IM+F+pJ1XKj7OxYR2GnYLSOlR+3sS8SlES
iZuS7phEDfaEw0wMDMsaFi25vvK7F/YdQ2q3KGoNqVHlDbjL9R50D+wBS7Nuhgpk
rjX0Rpj/RF+DQgv571ZGQBj1ZpdQpg0MbWjoImE0chSpiCMe3m38mmv28dqKCqpo
e9+PhwOKX62IqJ0Cs3Qwnja3Snnf8SRE7gZ4rDAuFVu2NsoOW0UQqVlvo+hleV1s
jOYzJrKx08D95KqU0D7B+8teFVYvh5RvhUQNLtC59iHAM6ouETeHjQabjCu9kglv
VZAf/WXJBtaAITmQeOubnCbeY0wql5jZ7UpL3IJgGLUoii+P9V5DR1zD6ybEZDWn
LfNLWMfHAni/SFzLNb472xxaEHXLT5127z2fM+4SJtr6ea4OD3J8xPoMd7y516DX
f3x5Jpzf5+k0tgiUG1yxkqgbvFxSC3R/C+YVfOnOHYm8UunHNvGaoBDQPUYNFAzx
BxhEiCmlHuNqxS5xaHC28nHD7BpFo/gXr8W5G2xrAxO7I2VUUCIY5Vt7FF+0rXT0
ge8wgUqLccGk/9Qq1azlSs6kDnaHaBnG3ykabz5L3m3bYVp6mnxpM2Ok0AVkdtYg
rJUIgfDSHCN7QoV82xaFJDsXiRTZhPvBL20D6xEvylfCEBW4Uz58EF9wngm3Diil
/lZEikzMhDSeetEM3phmzqJVivipcNLXZtebbmLunhdrxLn0d3sQEzEcDjbckCV+
DtsXH8UF3NmJduzOWqnPewNNcWWtr9bvIhfhbbAYdqW53di6q5Xfxk8sCt8GOiBs
JyISBIDi6681NgiFgiw0ocKHHJOmrOAimb5y6qsavssg3ecEFo6tojpjSeoRpx9Y
1n4B8M5FkL+n7C2phP2rXJWEGzFrz/SxXdkwYTN3Jj/joIVN7YlN2r55qp6/pbw4
Li5gz5G0A8E8N7gDvm/reqqJUjDpNZQcecmtzVs36a8r/SyFMHsrWS7aqBv1ICzT
cj6k+IX1p0xmUvKIyNcHxxqRGSfjFz4Mkny14PisQfiM7n0B3IPW/2lwp8k/NQeV
vv2nfqh2VUxJY2jFeGA33QgxcrKzIwCC2QnovSUKJ9WwPucN0WG4f2e0WbFJYYUV
rsV21suAN7ny8IT2yF+GNi11TJesngE3fQcxSAO+gZGYoqp6pTxejqaileJ+svS7
VwSJUbTPHCrSEdulfLDtSND2g06qLEhzKrEkOY0/OZWJYRSHtpEL66OYr2VmGg5f
6kJWwKeuC2/0m11b1+YCdtAmSPIYpYWR0EvrXVuvXzB2HDrUx0J+ibK1O9h86FFp
5bA4VcXoV7hUrcFkGgDk9Fb6DnpuLdfdQS9tQPnhNu1ihOlD+ENoNjIYkbeCemst
Eq3qqMdn011x9aDykLRyY8poWudRI/r4tSb1H9+CohqZyk4elr/O5YwJ9xb8rTAE
9WOlk79xNHvo9eWmt7XGoI83yAiM54KuJXBhuPyXKG2ze4PVGlLz2p3bxOzxwtnQ
9QIIoySGFzV+Z9cOuZXLlrXLzit+foj5j1BcVodEQUPWbrPq2y3dHInR79WnfgdX
E6DDIkzUCZHyGrGxTTTtaLp9h9OXe1iOEngU111rNGLQxjzftuYkFn4/oy47EtrP
rFINvDg5RFbYOS4iavKiT+v4Ti1QMkt9HjvnZ/7sFJi9UwZoFItkN45Bfta5cDhR
PKwHsrgU3NhKG8+giSRM5JtgxoCjKLUndzheL8nyPeoLd4RXyhQ3TA4IzKWg2TlS
detB5nTMpeW+yAxV/xUmv3qPEeHxas0v+g09K3mTsTnUVKAmqmGhK0JaWHIyjaBq
jYdR4YtP4fxT965EPfdaqTi386v3f2wzgz2LaLdGRZbZLFXlOuTwp0X8+31zueRm
mG89R8hSHqxc8PktqiDG8nHvMnSlVpHeSgaoji+g1yVy+yrpsqZHBURuSD+DPaLN
UfR97ZXd25dqlqxG2uKE18FqAxIzOoqi++j9h7pal+Fr3jHceRjzOauoyyowpDud
8oXpc5o76BKma3d54Z7gxM1Z/6MHAJmVIKOyKJ66AQZFMOF6/YF1oigeZ/tKuUcJ
i36AKrl2IoVCBPlcs3KOQbeyLco/3wY5hp7Y55+kn1I5Hfe6vS0w05J9yPlhrT/F
AIuX3njVj1R7oNXAvLg8ila8OB4ESn7w4ZRJ82NTbNkiokIuPiyQP0nLA8s6r9qz
ZAExtpdFGZwa0G5gzWVmV0Z7rVCvUVanjIxjqE37oUH5U3ChbIdKF5Qq9Qn55Dlx
zoEb/uhwiVb+afVfaBZ/9iwNk0Vhtk3prVMrDVAX/z8ATAVB2s6g/DM9QuXGueNP
Lk6tln5QneB6VmOzwC/AyxWDoz9kqrfCKB22xLmGCMerDZEvkTM74E68grCVDBwu
XnboIoMubuzB2tAU1H8wuya8c6OnP0P/mT6yh8bQ/ADaUk6Bxs+nBe+xwEG0W78A
TGO43U8CHYN7WKafkY8oesvs0bEgM9ahlOy0yuT3NjM90k4Boyrr5MUnlwMxB0US
vyjv2RTjgf3KvUlbAPbO0cSrcS+Tu1VqT3GtsrLof1rQThgqEsoEZJvJDcAyf6ar
3OUzg5YykZzWzpwuG4LEk6jqIlLHWcNdA3ZT9pZtM6BcPas5XHufHRIOfXoCc/hN
qsukDq3WoEJfl1FB4pEihXd98ySUYogIFK88HYNihRej+tgadlGl4qotyljtRdCW
wgbhtdzZ9szvlrjypcTAE0Eyy1YNJWx7b0p+OXSjTMOwkYOHsWEyFqe2daLhQbc5
+JB43A943i3XSyao9MLhLn347HxEjFskHAT4GejkNpIVMmqLX1XysfJq1OdFxQOQ
uG1PBXSu8eYqxK2FZgZ62V8fBANi2NE2aMzaS9ZpkeFB/WVmxs+yinu3dE/rhqDb
r/EJOA0FjLVCaxyu1uePEylN5zEQ17D6/Xo5kv2u3X/+YJOp+7Jk5BBzXcF6H0gS
ezlYWnKwTAP9y+X+drDgcZkPGRJ63MEnYXFdA+UqAxUlcbFMrB3DXBmJvKCeesox
Ss+Ju88Y9UYgnPJrM6lwA9tabxg6I7Lk9VEesyiKWQQxA5ZAcazjGl7lAAD1lCUJ
UOq8GH2ir2tUTu2ow2nF+CkV1lNQM2KndVJMRsB43ePVuqNNAv3wjtG4V8U7dwWm
SIEsRzxQKO0dIqkk/+tVuJ82yVaS9Xz5ReiMvY48OWmSFAdshSLKsst5MjdRckRe
mi2JgzFesOUBAaMr7KJLVZb7rQ7rpLgWllzghaB7JS7F18a4ZhF7UZxBYajfuu24
XAkvHw3XKVL4gJQiyHAvdIJG7KT7z+/Z0lkjI6JiQS1a6yXtz2P/EqvbbQCl5TA2
pgFcKcplGk0p8+q2VdOxVb+5hK+j+juEvkpYlRTFMtrtavVnyc4gZ3PDqgmzJWpc
1kH9p1dY87RffqRQogETHm78O7wybCHcJisIwdKIsKgU7IheDioC06ZoQ8LXCtSP
4xV8K85sOAie+QntNIu+mumaDYlqmMArKyMkqubihHRNA1BkWSJ8YrosdYSYDsaX
UAsegVhg7K3A2OTRK/1zRNJXUqQ/P3Dry3SsWZNVcWWNPRW0Ae8tKyI9Hpivrf7+
de2jm5O3Q1mKw8bnQMcC177pCqLIR1LG0pRMdVz7gXq6pFVlBXnckD+u2hfZETqq
iCh2RmchGdu3cx/5sUefAh2s4ssPt6kXgf1jragkm0qeiE8M73ZeG6W+OEpcY76X
lCw4rjAYGNueGhyeawbaEw+y9B5xRBVcY7nPLRCRv2o7kVLaBmuQ5Byus5ZzcVO2
3KsAynJCN160PkO2UHJIInxEpSzbXvO4aXRFgIkwZRy7KzPnI2b0rLqniRWLrJ4F
2L4CbzazTSN+Un6/WDl2PFbVXWkP4g9UMeNbqsxp9jLWOx8gZtCKxm1p25TqBRXI
r6omIUYhHMtBF9acV4gxcMfwHJ7xA2uegWDFHYXcndidyxQdwu2dkkHkIyxr8lba
K8t++rL/5xy4+CLV6I5+adLslvp2yij0slGgoTHei8FuPh7rKqFs+q65eFyBQDFU
Cobhyrj9oTwcDILytdbW6RzF5RE8oULWWRDRKJ3PA0U27Bq2MbNH4o107GtMYUPS
7Z8yJ5tcBix31HCTWJhzWpK4HMxI2pRN8x75gVRsga6gdBKaZ/BoGQbzhaUGhq/a
6EwsEyo5WAnd7ocFYvAmdspoIxqj61BS3AKW/QFwh/zNYl4urXkDiXRYHY+e/hvW
S1imQgjnOMtoWtd7qVXBUbWMl2nFgFH8F2yUQPYt/RJ9IONzzh/gV3H+DGB/d2to
8xGBaCr5TcmLUqPy3red6FKK/R5Vh4QOpoVfCPrlPvPCKiSw8QYQsAhs5k8oxY2E
1XV9vdEMM85zokN274nPjxwckTP02AUYHSFQnVhlNs7O4I7asjqXJU0f102EVkNs
ekSJhbXuqAEfbwBef54jxygYZq3wVWAOSVTSD7+zB6qaVlLS8bK4FjyTr5UwKbx2
sbocNAgdlTI8FVvJJn07q+3fDPdIEwFNwoaAkUm67mHI6OkH2F3QtPDwUjjhpQap
QZRviSiNffCrg0qPvu5TVnhGuwIKImUi6Bom2juZPvKx2fZ6ExgeN4UfM4TUbywR
PpAVnCLqHv2y2r5HuXiMnw3wS2K9YIlR75AepGqcQC2mjOSA5tnb4JXoIxq9b/VF
KXxNw1dcnIglXhKbw+1KfqTran9b+EUeoIvZhSyu4Wc2sjhc4bceR4lerFFenuJu
nxbupzC1neGXgeXVBc8goFjtTsZV6PO/mPr/bjI2K+6A5ammLNwMsQyLUCWOnhGS
H45ze9c/abyJcNqceUDASYMUVHjB3YhM8DNg1eSkkukyysQd2EXECAt5zRli3lX+
G1TkoTXXFrm+MTkw5SMYgd89sxHGHK2klkxU2/I26RPdvhgCqYpOCxk7oibGOEiO
PWCGauhI5XDjCNE6ooqZzlVIfEFr4fUP9xx56i3QRLtMdYpI2WXZCMLujv3DDkl+
XUXSSsgcYeN2Gqtj9bf1VdjljnEyNLapYp+V6uzAPVoWSqx7w2jSxHkodh6oflYD
bzL3ryYOmcv88dzNb8ycS2h2T0hKwl+TrUa3wYFpn4WiGKqVzFcBwFdZKoJdZxUD
ySwZ9CzqDOUHn6a+ee8ONHkDRYpDTYHh6mKU6D6d6EvbYk8cN2p+TzRfWrCDz4Mc
YANP+jk3pw/a3bLs6szqJRpz/ShtGKwWrjFJVi50s0keLCoIT95gXizUMjwt86/A
EHLIHJD7bWn3XZcyK3BdEkGQfvBuzCSRV6bCoy8LTCWyZaudCpJ8jsRHgs5iAUDn
j/5JwlXTQzWhsXUWbWD47QO1DQiszuozWmtP1qb8c8ZAO0NYPULB8fqw5HlV3lTS
B9XlRmYPgFzs5OGmJN0YP5pO7c/X2x7M9i7QzDM5W3ye3YVsqv2paD/AdAhM1czf
mE8WXJSDRUiKx59j2RE+ZCt141OPy9MtSGXbTBAL0kEWAnymOrZsa+qIpkJtg3x+
A+zJ0+LOImb5yLJSeKtpRRuBjMvKoWPXQ4Kpu/Z26S8S2ASHveY7t0RDpWKMqt/Z
bg49Fm6dyG/40Ih/gPaDAghUcqgEiacXsuOQANDGKrzRHky/1usH1dJU7rQAS1KV
oDnbC/Hg2um6kY962g4EtW8JhKcDMsYkuPB5195l70cLL3baQ0Q1uHvHBtIaeXEA
LUxirbi9oOSUHMnbk8d4YpqpwE9e8yzg84akTdovEocWj4xYc9ViKSpMMA+IeE/e
X29xELrDp+zi3TwUWQPSPa74fbh6tV75BxNrOUbt6iJWGdl3Cu103MJoJDeOM4Ig
ZVHfth9rLpuzQzw9IIXR8CB+HHcWRAkdNGDmXN6stXbL36bad8xWR6yWnKBCk3y/
UO9oMWWXh/LGHVlOuWrRf0YiecpDRyAreUDFx+ZlBZPRHy03j0QyLH/yk9Jgz4CR
iTzuGNpI87POUS56BZjHcUT3qj8Ex1y6hB81jQmf669XD2TA+NqfTJvUkvY1FkY7
u391zvPY9WCp/pKtWX4nEcUwJa4J7cHoGAXQOXhOjstPiazNX7/q2bEhSZ1+ZJc+
6+N9BLXLJgPrveml7B/2j8RKfVjZvTGE//G1GaquAPiTmtuvF3nxyKGGyYy3QovJ
6MB+J5db9uByLOQOeRJYjxl9k+Xn38b+2BUi1ONlWHSNerSsDg4KoeTCKA66ogs+
c1tnoEeuhuxH7H0tUKLOXtd7N8GfQso3QKGwCvO/Y7EW14973a8Uo93Lk8kYjWae
aaHjz7ovjTeuaehJADp/1oNPOQGatmL4C54EZ6WnUdt4dgRCXnVR6Fwkiwj3cFlA
2FxesrHhz2INNPPcQZFmjM9+61K/Xibx3jHElipRMaDGNps5neh2mJpmyvvXlxVL
qA6Lh1NjRKGa2Fpysq8Du3wJRKQxxm+DCgXv4XkG0YjJ+tgRTNNy4X32qu8HXjGy
BJGBivdAmVA/dQFj4IDBiRrfAtatpJvqC76FqJ/HK2dwusldxNzE0nOvU839vzxr
brNDWp9qt5saAyMVwAm5O2HIHv/Q8n2V4Ae6Tz4Pr14PrcXP0/tEQLtQNPtpwI7h
lRfsI6TD9b2R2/pCRMDiC72JQ9lC2aFhDCA+kRIP8jCrGbzY1lPGhsUNeFI9pBXZ
MM/M0EPIaPlwUM2Jh3tKkSJqd3j50hfme50oHsdDte/YrEqhBy0Beyhm2r5dgEQ3
BUOot1ZrcyoXwAbQtmH2G+gj3WS1f1U2twUrsFPeufNZhtp//vpkaVAwclmvrSUz
Csc78sLizKzM8rYebVIfJ9WdLY15OfaeMkBbAcQvvSQ0WeMT1HeHhg4DCQq+69UE
/e7PyY5n0CQZL0vmo5WEPgJzxVEgUJQeAxeykyxi/JYa01EIrPUUghz6hLY86k4r
8hkSOFSZQp0vY9n0DlZ32ILh++WeENnFnsigu4YopUYnzgS5RGtdU0Neji2LRNgk
dvd2V9L9b6jqsfRDi8Xh/5EC1AxKCxuoNsv65vXhjyKFU2bqln6/5yFQusfDpfLJ
+SQNmOQWs0PFfYH5uKRb5/F9xe7mQxnp7mX3JPF4mIV4tXU+5wrO/oitoHHSy06g
N/N8EG1BJE9WKROTY3a/TU9PJIR+YW7Op77NmvIrn/WO/NBZIEJCeyfyOhIselnK
MvVKX8/tU+1p026/hMS8/WBZdOkHX/LXtUiZQq99ETA43GDRrl75L/tI2qEqCULh
Vxd0IYL9vIChpE4n5Y8Izx24kpQ/vi1x9Eu1pgkDQGK6HxYJxuCNdgy/sTFqjD9L
uOUQmX9Nh1QppzwIaIdWdk0/J0DVz28YTFoXqOz8VtKRgtE3mqdFOD6rBuIINcz9
6iG7vy8RDg70+wwQSvhB8JO3kOlbAFDWFz9TvuH3p3QY4EpjAY22kXIqTelT3bx9
GPeUCSbvgHBU+X+7CGJ1t3GTDrG3z367sjoikfBEl2SvF8Gl/oQ0mpiOhkuibNRK
RX7IUjqvfmMQOZf/aP2a4mTVrPJdeTDJ76eAqHHxpw4=
`protect end_protected