`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1952 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
2n+M/KhW/CoPvt8soGKLVmyhX3bcJyovdzcQhCHkqDYJUS8RE7L8oHQDtNJMWDcU
zmOnxinqurwFS3a5dSfKNxDrpi22w46b27RpnLkYR4OArQoim9wf4p0ODepK6tJz
TQx4Y88omxBEN0o+bN2YdojfjcO+hGHMUrhDpo86xwZyHjQyN9TtzawoaAxXzqCh
2/4cIocFmer77V/gAHBecDCitrQ3BbYyJqYxYma7AA8MgLuRysyj9g/JGZI2wPUk
FK+nEkhL0uhYhrFgsw+rbu+deIfrm57dyg5xpiwf6DqVolCkOWBEmxlIuKAbKZHV
BePVYOjEripxIPvaaX83J28KVXdOMZh8k/JcSLv+FgvS0qeGzLbEIKrZpTIpnR2+
b/LdawsmoB/hcIRtlKQKw3fQUijBhBx6Q2PUwvEEmg8ckER4zUKwsxH2UFQ/vIgt
F6DDfCkhIsfw8TrT8uNeyrvMChgVSdeClxG8rLmtLejcUHbzKy3JgrX8XqjG51Tx
Ls1+zxbCSfg8RMzhRsTl881HRr7YfSnEndqH+FqDfhUrblVTEnGz4AJ53xw42os9
o9OTl/BlAT685mf0EeF+BlI7i0ohHUCfelcEiozAhsf62RbpNvh7E54ro+gmwyBU
RfJVhIM2C0fpcuUG/BvNOXASFkCbib9hSu7oJgLTNw/iOfiQQ059ytPe5cOmR1Cu
eCqIKv7f5/b9gTFDIg0aJjhPtaHHggKMyCpdTAyihAfhFVfQpsjKj3C/OyRlyiJs
uqLHkOY0z6kbtuk29fPXLaM2DDWGOWJ3vMGTt/sXYyFq20eigVFgNpWgOlV+VTpj
CJwqa8QD4YQB3083R2UPDz1Op36OgsK8c42erWjl02p+iiu2Q7rULf6myzw9HOKk
CaQgV1OhPDeRSG+w8qQXVez6MFmGnw+TKWhPmQw2tfxEhsiJSim3SNS2Gw/7hCVh
W+TXJAigYAGxhnAU/h3xpqdKxleB4X6koxzqljkXk1swVGP/afg8r6aTYmDbb7vp
kuAmbNtYO6bREKfVBk2B+H87eIaM0zjK4nmgD68EPVVkK9lpmWmFMHIYvdcekXmC
7WojrmvkIHy9gGzN+TvEnjgQK8eTZinZgIH41rejJ1KleXe3UNkZtXMFdPZJ6XO4
tw1WHN3BCmM3aQFQvH6OB0gLAGOYGyD1kmHWA1wO0ifmBFzqfV7ZjtGv6seXtSEC
fxLHE4G1UOK6NLFm4jJcTe3K1z91uomNSZ8FWSUf3mOcyeRBUmHKhVpeHIu/6K9k
LEDipsWyneO26mLz7x/udx4Ux1qqerSJb4IBCsfFFDGqYhwirccvsETJ+B/nCFcE
9Ro8yovnrsO4ERg7f1p03DMXq5cDCX/vSWaWm9Iu+y6f6/Gxheh4nan2HA2k1VIF
nt/SlkALMRzT9BkAlgyv+uOVcuwUhBgdIVoh9Vb8geU+OnYv7HT5Rl078kHXbD1r
Nkp5EjEv5JUvoXjqD203/5MevP7vfrmU/aysaVhCVrvla2/jyz3NQ5AdUeaze8qk
5mBByeH4+GA58Coh0hSHDIfrjf9dtYFjVEe/U6h72ymUwFSvE9DcJejZiJTNt+Tn
Xj3wUzzFUAJDb9ky1gNjh2P+WN1holXEBZ2aFaemHcv8wgdY9GqOGDSALEPTvcKH
dbh/er/kkheQCxfVPqOcQSNgcBqEuwfTAGsBUKwby+To0BLWd6NwVxTEqOCOGAlN
KhwL9MofloClk1rbflpGx6j7B52ZAjMcu/NAwxgGeCh2SOR8hKpAx2zcTkWVS47X
qJvl0KARtsvPXVRVjtCd8Jsb3vf5NK2waDMonbFDixJTYJzfzrMF8KMpOgo8MqAG
zgWZGM2prroO2QxtzjoYsIkL0go8ERvUNNOmydT4eKkW9I29+ByuG9o30dWpZr47
IbBrinA4SyIvm25G0cqDXuNkdGJ7kfOUM/t7ImAtc5n5pwWzp8joIUnRxotXHeD+
qbyGvdAhdL3NwSBa4Env4vGCRWN5JR0MFK9NH2ORpI0P+yq8JNErwHQDvdmX1WgR
oS1S8qmKgVGc4g0MYGVyARtL8ZDs5NYsoKGZ9VZYYPoPPElc4ESY1wtl2J4is2xO
sld8XBjFcFKfLli2Kjpgrws12doJaFjwEq8vmlU9dO92lJKwmXmXz/1MjYrcw+06
8Hy8yx7NtPew1WfjjevZs+WuAzp/kkiQEAShPdj5u77Y6H5+bls70rW0JU6yFEW9
bxEkLuU7+KekfUp37wCb2z4cy3js50rxOKCrT2tCrrvWwHk3nbRiYpJYedqINK8U
MEA8+yNswIP3xrOpOCWE/JasmAfwSXOWAzMVf+R8xOlRTG5/MzZB33d/EfWSOSNb
DxaAyCFzgzUXS5zyCP4uAtsr8ufAybE2q/a7m/vcElsyJ9LgDxeX7lo6oBAaOGcP
raeCSq9d5Bl1ts+8+O+xAGUgX40/8VlTBQwRxoh13aA=
`protect end_protected