`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aMReDmrPskJscpWYThVKVItA5gecPPZO1R595p0GoIq1TSTG+UxXhmmUXc+VYHJ3
u/C3EW5qePLufxmXxmhmDnr9U8/cYC1zLfk44v/2OPb1TBrTsludEDQZdGNWeV9l
cPUMSIfZ0dHXN7L1M1E2XtgoTWQxf3VDHs7B7lU2y9Rdm/ibz0fWMow7op2nWdD8
gJ4QlNl3f9Oiotp1p8vz9RFzzZOF5gBBslZxcTF5+z4qO2W7+xLByngthWm+exIr
3Pzy8qyUo/m2DDwOz3VJSvSNm7RUq+0/yJNOOz3jr3j7ZyCj5OqT/jDAWjJSMH+i
2402Un+wDMOQxi21JLo3cA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="5R6K2aWI3OdbT2A+sz4o9+2XAInTqB1/cSw5W16RnA4="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
Gm/2BIZF5/H5qen8uQizPH9RftTuEE9mgEOF0SqeOKegtP64CfvEUnIxj/ahmIpA
6xUR2v2l7E5duaLZh39Mc1GYsfqE91NCPU5whLaBPg0UuX4cgTkO4cYbW/7yvcrd
4wavUfwXEp2VSiN7EVxL8RcZTSMSI0Jr/aojiilFqVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="TEmQtJ1Dsm7TOzpJk/CeTSSFx/zKExk04H6I8sT4Meg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1456 )
`protect data_block
nvPqn26PC4XWLLQG0Fq8XsMTlhB4evbpiwGjZroFFLgtNlE6bBjdtwWsB89WW4j7
jNfYbKN4sBv0hDeMH0AAR+8g+TCqoX7yLdIUd7aGwBUZJr6FdDs2wTUxRkXFYNTL
V2foUCw8RCp/PMc5/qua/o1cTs9+qVio/ObRRmBaBokR+0e55ezMye/AMpomTCcQ
rxpeKTtH4kAu/yb2TTaK+S8C2cwoxQvLnU8ELP3xJFqo/+rrxmR6lfPedEbbB3qv
2TW9U8TJwnUfsRUIinJiz8Dj6OkWDyb3iVxqOjXY22mKaby5maYsQswAMc1nPBcH
s/JR7iq7JeRBbj+pHKUeLFPmLKfQjZ1up1OUZUh4Pu6zlgXWdGJcwSTSvjg9bq5D
3EfLXYuO9f9e1LCrPTenmPj2gYYNH7sWNEwa1QDnHK4OwjSGoJ9EUI7DjCPXagDI
ajV5vVwLMCmu/upD/mo26FdF8CJ2Ydp0NBewG0J+iYFnoXh1CtikVxYOpDYonKvF
LeGA8j77mGuUtf7rshaMxC+x2zP29zk3hPPa+mVXb6RHHh5i74Z31wENXcpA5db1
/qIS3tqgUK0Cpc7ZyXGpbTmWuOxch7HuvPN5ahyaoaqBRGI4ShCjmvevX9r5/6Gl
AKotXNrwS3AEtX4k/6MYphZHZ2vcLwskNmo4X1qEi4DWCHVHUDy3+coaIsM1hBLk
RPt1l2GjS9vF/gL/SlO7D9pVQLGAx9XNuMQUpno3Vzc9gfR9TqALN57FkC6acsZ9
K6UsRIW+/Vh0h5nY1hbXbKKtFZ0CDl8j4IJa4TVGh/sD0hBc1N24mulYS6h3MnjZ
II9fRqxMtgNHrbAKZ09LobIZQnLEHqBlO9lWotiAB8Ja9tXPz7D0o4E+tzgrUfY0
DkNG0En61oNHcwg4MXPp1zVMfeeaXxf55/aMZN9nOO6ixJ2Wm1AEbyBX3lcr02Kq
7sotudzKuYabq9Ltue3vf1AKmltaLK/x4FPHlattYeXCIfqD5IRYM05riWK1nX/4
4/JXHzX3WS59yHxZl2EMp8BBiyqvlbqZl0sdQs2B9Y+g7AWuPRe8S9pke4ldDH9m
hLQFfKnIeM9/UACsg1Ta0SwiwKGqMISFLxYayqvn/JQMV9GmVfTGgMn/ydAYBYzi
6BZl3zgC6HcedY72qZI/T+B2ebn7pw5X584n+npEkT8Aai6+oPXazjSi8MQTAnhk
kONe/lBMtHCabm1kYI5fWi26hmRQgV8B33SYW7bgoA711eVfkmrf7bw3ghxffrPf
kb95jYuVC7tuwvbVCRc2Cq6dQXK1iv5XzwNulYPYoptHy+0s1DivTDynb5nY4Ih0
dYkjEbxyjqvhFdFHX9U3A9fBudtbjOxmygo6iC2EN0VoOKoms/EME5YcfcIR55z9
UZ1BYUw9FeNPnr91FmTL4T3MqTrhciazFLKCFeLbb5o3uSONKeHLY69uc5gL5S72
tns6h3w2nv7ku3/s8ayXs2V88hkKW9UY4004I6GNvbZ6PVUq9BlZu5LBT8iNeiBp
FqrVjobHsFvC+GxBNGbZGLO9ahBAJixhz4YfV3wmRZQSW2bpB1dYnCqw5rT26GY8
O7llIbBvMcRmdW4OPoT0pWFZjK3VqyIafK9eDAAxLu6sQxcN1zEbfzcLH71vzAQp
CyFTUgywx64nijRCM6EcNW2vMwpHd8T45KQgOuyGEKVf9XsOoKd7eIYw+mojTW0H
kywG1+jVk24j9y1NwG3/h1ITS6g3cYso3nsbiNN7Ho/JRnxBblbOHqB5Ft7zl6f3
8d3THS5+/HtFKeFuc7rLIuynQgcutn5SLrwou+GmS9roKuTSQLAmt6yxchmFGGBb
vTUOQlgP90YkOjRhsPejtWAbzs1SLhT1g/gNoPfWE8JeeM6cclp6wNdBtAfVJgDD
BNrAXZ7td8CbEO+jEY1ufQ==
`protect end_protected