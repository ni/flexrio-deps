`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4320 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
LfLaKOw3utJqtz02pVdKf6zy++vNSajXD5gU1PsmWgoaaUd8QUH0BnfIMIFOQcGD
STZydUWfVsyMNxxHa2ZB7bzyp/RRA+ns3yBE3oPCbBRfmQktNjqucfz30/aCh4LC
KIZA7fE2449HHS0rym8XHlw28LMxiJxruYexOKeNkBoSnufQPlsJyF0qj+iufSNJ
VT32BzKRe/Fg/3r8Z83XKDHyjRFU9AH48fmlQs/XWnPNagBs3aO7Q7B+CPwZgnSc
aud7+fyl7Uey9oVUiYhzVvIFyMsoqZV3esu3Yd0ThBBuGlAhNvt87Qqi07o4lPi6
hGJPsROCGSBmf6jrza5b3DLxkbU8ylxoEOgC3FjnPCjpQKX9pnqqEb5Pgo6Lm7rb
0tsAX8pubwraUlCwgdcLxmwOLfSXHohZYaff/2SEuxXChI8uM/H1zARgTqwcb2U2
EJZKbZteShrJsskuywl/mEcjGR+slOs3ZVKumtZZ/OpGxa1n3vexdnZ6tH5bwaZ8
G0DkQXQQccZM81bofPpqeztNICNw7tGiRT04U8wMZ3uUWBNOCEfbzZDJSW9h20dB
cmw8cIxQHp8TRvq5a7kxaU6/R9rB7xJL9aaMbbzkGYHm+HePkFvD3ZRUshkTnaPN
QMiu/8D0gC61NjPEwXK6FAyGYhp4ajoTEkUDYylIcI5FwGUKVSf9ikvlkc2YCaoz
GjXFgYRv2oGL9twtOSb8LjTOaktXDx3rkZIzMpJ6sja5rFV1dLD00++4pHcsI6AG
Xa55Pw2XKdZQBqfPjZDwvwEGf50VSbb/cWuXc3MxlRGiYJgDHJ8x71ptxxCGeSw+
1HaVmYuIkutE2m14ULC1BeYuIsLlwtnQWBcU7fAxvgjrIT0jANWX46T86/TzxbI2
wlpcxOFR92r1tWzRkBLh/87//ACUk5UAceLlBbIrKRU83EiR6FuPmobpCRuitYLo
1niRVfVhkjqR5IhcxMLb4gOXVbdkvkEavz2RCYudTWBWXHGs/aFgAX65wgKuAEYX
iLJsS4KIt1WjHVLTFA9YDjCslgJJfX1hWWQSHz3y+ep2+4JeS8QLwmLvZ1Z0ekeM
nXxUtLlrotxiqBOKgzw3d8xkMvUKWDhEnugHK90JVr5o//lC4hyHG0T5jtXRSqkB
GsQ11y0q2NCyKdWuE3KdII77odbF+4fTGUMKPkHA8EO2+rrK9nb8/RB4wqebyS7J
4o/pkILSrgvTRc6+DZ8mD5pGj4f6RG5/rI1z4RF/3I+sL1NUqDznkur0W6mhqqAW
DiL+5Ur/2fT6VDUylKMwQp5qByecPQCSpVh/jGdcGDiHamHmg8WPm8Fgtz2Ee0Tz
iq/1lELqvm+FH4WvYs0kdUTHhMdeSuouDR04tkbTRu5fJvCZOdPrWTEglD+3eDB+
ssPwaX4lVICDoSmGO+s/LLjTZ0yx4/tRwz3oTa9CMdOYcB0+pJI9D5KbrZntTHD4
IJ3DyR0lfOX+NpcNeiRTS87G0yvlnTDCl8vEiYVtYv/P7FLMpK7G4R4Z53PtCBQh
19ARTZ2hsQ2ggm5ZbyFjYzE03n09puCclIX8rwdF5laYv9TtzlGw0Ks/pxVzQzMc
VBTrgJBukblZOMkpKaOuqg9dDnRVeYevdnuHACMie2OSfA804EdPr4Jnk9gTRU6i
V5/8WIepsyFofK/Jhf/FBdfD0g7ciZEwaKOhnBmN78NHZcj3YGIXVa783wzjr/hW
1JzqWNgUIgiPnPYCx9uw08SutjpzLS4sL8eejmHObAH3A1WyyINAUEiRmSRy+5EW
wpzjSCoTBypDC6uZ+QBXqH6fv0r1ePggcsKGSDLBRcxSDA0VYj9r9xmyQqQ3S4SA
wnCXcU4R4CozanliiB5s17Vc6hgawk8+70Jl8Efsf/Musjv4dPHvrDWy5t+zzcX5
8Vw1mzzxnXB4HgfceN05BW+QVLHyKgAtleoSrAnVIQO+Dl3JwS6eHFkMrZOPEiDj
J2snL6y7XFmpjg/cJ7rpjl0Uag1564a2MixIb97gXk5Os9LInppJea748nueJY2e
hqrFTW7cOERX7Np5GAniXmgEU5lm510XtRN2CIdjvvXbF2W6A9HQEVb61RE6JAtO
zjVSD+rYyvK29LmPxin0hnb2eG4ny3/P8jhvhx9rYmlqy1lFd7cXWSw44H3w84b2
yujKxMUn4gWl3WOQYLFW5FdZvTrbx7TWmRqQrna9elINJbN7p3w3gwi6RkP0ZQXe
T9D7zyolqS0e9ZTeBhURIXdVnFmNAoViT3cWMay0aUMmJdsQMDBumZ3I/EuBKc/w
wY8Xnq4FaUBn8fshKfaCLdgsT3wVU093p8Srrk56LKJwCOLncuVDf9+Glo6IWGv4
a6529o/6Trv4kFHPti7dD9bJRln1u+bX8eOnEhZnftLK5TpPrZBzs1kux7/JS6xL
GUW7LfB0cGNWGkf9tUL6UM+RBkAPEINBTkzyEQXiuEE0YFOZc4aNYS1zGIMPKzqp
ZunZjoErn2Fasf+niFLA7RP/jPh0XUBFEdOXIJ2TeKuNeQ/lAPQMnrg51z/LgAy3
wEA385fMw7KWBI08fTIB1beNmc+yjG0Xhq6ySzDdHHUboijtgzXc7J1y7vCc6HSm
/L074DX604Y4YP6PVaMtBZ0Far+38NjOpeopxbe23qeUQJcx3rPZW18MJqxFRvr6
ikc8vlPB4AdfXuGyUbkNPxO9WP5/7hd+TAzotIqWJeyNeUzTsPP4cx0Qr5SsNYif
pZCePbmSuf+OEZ+Cso+ST71mory7O4PwEanJb0IZUIeK6ZmL0EZGMIBKr4qrH08k
CDugdVfyMZVPnHKLGAQqNsQiEXqeYzenkdz928n7cYiYketYPltdaUjaYKO3DW7n
xSq2xwevTWv8Et7x0rdEtmaPLeGegpu0rN5Ga4juZThKt+8cOaPRhtjJH1FzGFpL
oRIpTv/h+WvowzPqo0/qE3z9+l0r0OKPgDPHqQiaZE6df+B+RlBwPZtbSsEvm8BK
ITEpUosVHNx5IoKcA5QcwSoucn2SXOshT+d2Jkzmn6YBcs3rYSf1uW1YUeGPT4L4
PSSoowi2IdOAxS1W2WaLDHHmVAPlp7aXhwIK/LuvZ9ZLcRkYjlvq8eaU6pCkp92c
bfc2dP+lr+FlE2gqNxCgrO5gPP+wiOe8SHD8j5UwtHHb0dvXjT8D9Vng5cBlWBCU
0eqg2iksoXFwXkbfWLO8Ikd99qJ6UWBPv0Nl5jH0AdjitIxSqfSRjpxH70HsZ7Ek
DtpEnLDbtDcHHEL2/TuDsIlynyibwvh3AaSceypEhIVKWlfeAcn5v8QF4VFaoLm9
562hvKLuxbo/BrMu/X025K+DTqTFMQ1uKNwl1e3otDs0XUbKlC2voFO5+gqOrCa4
Gpnlv+Y8X2IGT59mglninQqC/GFiTWk0g8xtDL12Fr/y4QQs54VR2Bubs80LRHDl
wVYSDKwvV5YP34p8XTd58+akY4dAvCAOW0WRsvVTHNR2vvpylp4k8/z+F12LUxR8
CyblN1uzOKUpZ/EpLa/qdHWhAalvwm7q9JVacpHEhqLlF45t0dVe/AuD/sF42R/D
KlWTYIT1OcIGLsUWETqiTH/5Fh0spPdFxgzBQ9osdQ3OPBf4tOEefFbpuEGCHl9l
y0Bs7C7YyRlWSQLwf4HnWqzs1QW50s63ykAY6pu2SGTs5R0xV5kyuWizQCafe3FT
i06qwSk4/ld4RrsNAguHKLJ4alZQL3FZZ2Ls5bBpTgrVJ6mhipeNhsoIg/bNfqjN
u2Dkf8UI9422KNwUbQD++EwQ6KfCO8s+tT1z7IIqf33jv1liLwpcolwpHtpZHU8w
pkN0Ycsqho0X0wJVSIvP9j+S1E6BvEwNwB2TGqsJfvXOn0AewXbBfnNX6yPosSX0
m6UoNHQ0eeyfdLDHfIPrBswb3A9SXqzbjN4tPuuZ7pghWc2YiTJhHmcZewfefqPz
4xPvE3psOQDTykp0Xd5cCqv5bw3gw3VTB3wlx3yXfBQVKAeuLEm2fBWK2H17LF1T
PVr5MD3ehoE0b4TK3cVEaPhwb5WbiEnlEHpiKA8nVORKdUipV9NXB4vda82+s8St
Pn6PdeGGk2sJw/QLcfooEyhGdcT/Q2uIxhkW/GICCL2sMxkjEeE23+vQg4eWfBAe
DFruvw0NqL9czpoMjWj8qO919b4vX+MlPO+ou1FNONfbxrxkI56e7e5uuR2tSA2P
JRBDCsyeCf7bEbO6NZHLdNfhtwjJnoBsyD6hfCE5E6pAVsWMZNWSahtORhr1bgE+
xVFCQCbOtV/De6OiU/JnvEBF+u6u11JmZO29x+eCmcV38eIWmLl8iQNGH7Mc29M/
QVPzcznJOuMRVeUGHewlZ6W/alNxjnbuDKf1NERO1x/PXVwPgw+MpLlqDkHgKtb3
vNgUs1AZ8isy1zlhCaXBW9pwJffKKSMlEGOFm0eBXsiuXhFq0CPpK/sRlGgZ9F1c
rtO0Vxth4cpwN34qq5f7onZS5mVTgHcQf7+7lDU+UOIj4DAYFT24ugidc+LesqVd
Yx19TmsqkrkDpydIqDMO6jNCgmRhPwnSaUSJ2FKAgA+fl2qnd5NMGVrej4lU4Z0F
guVw8Q1JVHgwiAitVChgzosYCBn3h8FebyicF1RB7u9tyzXmBlj3w7VUQg3hRcRn
Ld8FZ15Dr9CEVixY20qTclj6P9JL+IQdGwYvUHl3on1+JTSB5Xi6RAIo3D+YH+ff
65Da3HNbOlvgbqp9pCN++DgUgkczbU/dYZGzUYQP7X9y5dMEh+pqoXIH/zfOjD+f
k4NwCIVbZbsxAnSSxkfzzDoVJkTpzKJ3n3QCGmTWz5p8YT6oVJ7mcd6KS42BLKeO
irfxueqwl52TWzTI6tDADJmkMLAZAwrpwZSKuz569+XGXAuOb/iRwDSScc+1nN+3
KwB0EdJt/97L5qH9fn1Z99X2NkYnj4BpmGEEzXvXe+LjI5BJu4LYQMeXhHhz9TzG
otnERhJdwOYOjvNtftNs9kfpvFJvIBtkCAOM9PBxvZbOUzJPCqAB21280JjzDIyy
6f+X1uxzmHoknlKrKpoO/qow2i5q5SsmH/4ZlKhIfbsuFRqOTH5VSGsZQBJAPC7H
y/+HaChK75ok3GdHQzrQYpTEYblAx4DaI/HVGu3p+uplR/N9z2eH5oq3lVBvKbBS
dAUabI1Ax3uqTHxyJ4BouZvHVQJP5SHCOzlApogJCGPS8C0TYmpIwzwo2GYGdwb/
0615gJ65aY8uaWgT1xlcaBRJiHiuyvz+3auyp4qaDwtCeHdZS411Atga8nSdUyGz
WDMQqaUTMOObsw935BjUUOrWGSAp8jZUvq9iU0uPhmK9apdpyYX33b5Aem6hjKkB
URS5+re1Uz17EQNergASQJCTgBEa/6GwuYRZ8MfsRbnr7LJcZql2Nyq5LmB5yFUQ
RW0hDo18dPSS+PhcUdzv4+Krgs/F3EDcAwjkZ+jLYAukAEtcSD5m8N1NxfEcBy2r
rpXo6Mv7xDVKvpJQ/3wyAILhpCvlzTtprsPLB094w85tSzurPlHAgKGdV5x2iRQR
xqdKEEj4cfl+s0zcIq/piiueJT/bMQxCJ0dMBr6fsgkPi5MsA7p8JBDenVs3YInp
`protect end_protected