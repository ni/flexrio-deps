`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
j9eMmSPGcKCWAR9PvkqZ1R001FU8QKTyJzFqNLn+qur6INyYDE1AI8LWcxAzfnTc
IpZG7ua3uuk5/kQKKQx8ZIPLfmv6H3t3eWjki8YIAtY/d5E7Gq8Z5mNxMYRzGGTg
TCMm6oOrOTVYlCXHE0X9AW696Z7UGfWirVibl8hs19hrFdeZKGiGht4r09vHR+Gl
FQQmSObM5aSK5wu5KOrK5ZUKGHyBhjnIQO5NnittDjOwxV/57nHVg0pdG6JUqyvm
tEgmCY36RCMRGWN7sekPtNHjqpZkmYrVX1T9QF3h73+8ZekZYd2xY2hpHHGYYeWA
t3+Fmb/6NUmoP8+Pt2hI6g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="wX+NBVcG/A5ruHK3pkDqG8ZVPdOz9TJPJ5saXZYSeQ4="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
j/hqWUoxjK88VtH4QmjIrexFOSwtsLKOZ/LCP4cmrqgzmR/e71apdtoL+o8nlfy6
eZxDZMmrZmJGoazz2oK6kz7xJU85UCwNc4cxAsVxNdCP19vZxph/nCYZQ9lUFkLH
uLBkOeFP15CD3jG5/dp945fHP13J9SzB/L9PWvDC/gY=
`protect rights_digest_method = "sha256"
`protect end_toolblock="sqDZkaglKf+bDjC7VKm3lOELrT2Jlynh4UhPg2J0Q70="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 33072 )
`protect data_block
f9kZDbPp4NLiAOFOgATj9W35i3s4a7wbt9jeHjHVcJxMoXY8rb8laqS5bNUhXGW/
MOc7UNc1VwolqhkS7G27SLamkGClZZtXSbRcN1N+5kZpEaBEj1343vVznnU2Dre/
1cevKNyx4kKswjhZbozAMgXelRE4KcDYkk45BZbafEIEjLpTUKemXJ3HGvQ594TV
8yEBVaQkrKKh8alrjLOwSAoKIJuMmuij2J6btOdoCp3XBn1V72i12K0a70cmyCUx
YheY4djALWsvV9bAZb9Ve8hzLwW0PoTbo2QrbQ5/D3p11AYi9k/pA9YPmyk1msoX
51WHL04DSSz2baPNrykuuZpW6Y7ozcM96gmvdDgPorRXtAeLeI13270b2CEHS+G9
mLQPp+0LFfo7v3x5ICW4wjQtwnrKAvaUFYzTyb+YsQl5uIdSDPuHINVkMk8YRseD
+x8yCHuPfWOcD0KzHF6gnD/mSoWnyXgmfS6/lO+Qc0Pe53P/lM89vqjiDO7pfd6M
BnafGBPwM+aqePkLEpfcFqvHMtV+apen9JdfZydGxxs0crKGb+rX0dG+WG0oIUj5
KzR0F/wElFeNn01MnOisvknFVkLM2VLkt48w4jX5ZFjcHG8SGea/db9ZLw5m8YK2
rBj6OZ+iLT3N02jkp3bBvY3VgEbHucX+rkyZzhUf+ZTmIeFmp/05aAX79KzOSxJl
zZHs6Quu8b7wufxeNNouP+fL1NHeHFGNF7aU/5Z6Gb9IE5zFM9Vx3Bqze106FX4e
I0hhQUK0sSf4Ly7wejxyO95SYxIW/MSvqexZE+96lf0n3DUJydPMETwIvGAFS+9c
bxHnswfEB2WrAZKCTx/ntzvMvGJXmYXXNpUvT3MwFmC+lwaoygSy4xPH5x/LXX3X
LGMLrC7YgqWAQJt3+v/j6QifV2tMIvViPzaa11rAh6ALFoIBjSTR69c2gPtHhkg0
xZ1GaCbOq07lty5vRjr1ZIdGJrUU4s5GHyvA/YtBq8HDFPUmH37wNYv/4dhataj4
Rvht+tHK46SqqoI6DZMwkMaeBtxsD9MJRtlZDKpVITn+TLP0gn3WssPuIh3HGeR5
HiY6vx+L0X98rVABIrBGmjUCfUZsM5kGecpDYDSE3Mo5Jxk8q3z+d1CxcweSmBlS
lI5CDiqvdP3ch2UOa7u0UbQ8VWJdJhZeEGgSMng+JgGJbh0W6ckx0n767OynE1X/
WCRwlCq6RPUqtJ2b+0HAyCkvdrdsJz0fbkuUMHn5b+FMdOgR0PFBn3cT36BHwzgs
xajlCux45Scg3aLbhO8zBgLYPQnbyuArjQt7G+SPx035gJVoCBQZdR3pCwU/yWAt
XnEsz1cImJk922RKMqAEO4WUjbCTjCAS9Iv3EpO5J7XgsWxKJeRf85/x6oz8OgbX
OCOYo/Jif8sCiQ1ELiWyj23ldiXrkRaObwEVj+YLGrAyQbbPjSWBuxc97fwM5ivZ
CowhKAmkVfSGUMpZnOhO1D76dbVLHdB6KopW4F+MQXMNk5U6LOn53CArc4mWKdKl
oJ7fDhm9RiFwOUyEcz0WeeZUeOJ8zxGgRF/Jrnbc5Fbq8rid2MoYLyZ/F0380cMB
xxMew+BCGfnwDHI6WxdHISwu/g2fYirvnjoQ7QPp2Jm1n7P472nUGW9GhzPFhq01
N/TA11pSSSmXnjLHEo4isxyXNDWPdMj2yWytbdJYuMId+M8/D8viTZ0QsM2j4kL/
2CZpXzFdBADd/yJAH38cc8yzG1cNRwet6jOPGJ2nH/T/b/7fypoF2uSXYZ1u0+Rr
1Irk3glbo98WnnGdXzADISBxwZidC/StdQBYQNynJ0kcwTUJGSggHcdhTNo8p+lk
RzuhbD47tdqH+Lb1bTkKrCzeZgyxMt1xNZ5cagSzqQGdIhXT5yKOcInqDsIrCyzi
ymNhwkYVRgInUAMxR1uxN7D6J8JW4r/b6pSeN5YgfzUZnjtpb3VoBk9mtyJghhqb
pqXKJDc2xCfgr7g3k3bDV+Pc2jSA7Xri5SDMb0Aum/Dna3Anu7DumhH2afE43inR
PPKb80tIv/wYJ0/DBy+OgUxV2lJeWgjFDJ1fIXkgSSmM9OEJl0vrtvh9nwcHoxb9
IIlEgUmkf4WyI/1bARPFfLnpWgijmU55agPoGtYvGBIClnhzTYaZkk9ilirRopXv
+yw8VnaoBeRR92x+zDPipWzT/HfM1VGYrz+H9GUqfB0whEsiwY5Na8z7lwCctHfN
pzAYXqjjMz7rJl5V1TF2G93BhMQzilwieBWqqXvvLIkQNtHyKvhIf94irLr6GyjD
YrIeor2diEAEEKEvwZl26C6geI0XdCcwh6yXT+uXQWXfu+RCyH4E2s26IPOEugVp
gAnaBVVkyOXVLL3WB/z/CBQZX5Y2Fsnfc/TANDwEoK9Ze7k8g+AIBL7y8YTV8Tp7
4m/95YmGb5Qt1A4F4pGu1D5qNu87WRvpiiSK9jhxUC63C6f9hi2r0foXAcZmFSjs
S2gphnuWAOllce9brXGDFo0fQiDRasUXmmD+RcZecWqjMK/qbops34pUXyZo3okn
qbIaFA3+l8swFVchSKsiA/pyzdqHFHreqJZiM3SP6GMl/q33S2Ng6S0BDy1ExMe0
45zhdL6H7DD0dBAx7QIVuy3N/QQdcAy75McgbU4JUGvCmqG1oLqRrAg3R7vTKPCa
BCy5O5guhR53R7lYLpTdTpVbXzxTp1XrPRFoRzj1u9sLuq8xNC0mHRc6f40KTPFw
r14qdSOyj8iKN7LtAspJqVsuUCLBaWxd5BjG1W5qDhpiE3adDXdTlE16ogh3wbFV
m3aoBbXusPbUvt35s/Yo4GVVqbet893bEduaUbKKlHuDqn7ud8eDjxCOzA2ZQjts
B884NPD/P+j29SDQBMlTn7WKqPXFhdbpT62V3R5SWJ/tbflKaKF2kWCXwT3AvC/t
bbmSk/0s8Jxy9dIR2zEEBQKGSv4CN1TULOhrocNw90FxHzUQPyfEhZjNt6wjJ2/A
yPXAIkOzNFxY/QWt6osAXQDARjb7OBgSCxChrvBYudijryNoSOb8AvnaF555PmCw
ctLK1PmHo8Y4dXQj5WNCLFuPLH2RZ9VcP7kxA5TmYU0SgMf9JBLq+dpGZ2thqdkn
ZL1OZcBs0tNdHVaWFCfDUudpS8NdOSv9HhwNmeKQFtwfsceDY9YRiUW8XmLTWkPz
hXB2YOnRiBy4O3hJaYlBUg5Z4PjR0Ks0qdbtKBQu64kCd3Or2WNR2z11eSc7ZZ1H
L1O6NQYq8OOrqPmZbw2ay+x6rnDw5mGFSd/ON/481F+59YMOg8MzdqOqwu1rIzQx
/qtVrrqDMcSD/6T7SJR6d8mMcgJCfwBw1605lY6LTOcIL/gv50IE7Cq5h2EnIbuK
xepwEbj/PUenrzvPeAszgxjZ0PY2yN9d8AP7OWyTSKVTQYzDXHQRwZirf5+j9a4P
+hL1DXq6PvJ/NzgV18su6w6nio6AYh98d1Gn9ZpIZCehsaCkSqjQ/DyPKn1EdazL
cfE9cjJyMrtZm4shyy4PaUT/Bfd9E+e0zqcU5xpIk33cP6aSBtliq/8HB/STJUv9
K5caY0LFnyGQBos5vJIEO2gplBCwxJNWYaqO90bxxUhpCnZ6VdwoQNIF3V2toOhg
VoReeLCX2odxpGHJ2vWwDuhLduPPYAZdsBG/LGQQwsxEJWcFSntGdwT40oxZtHhi
T40Nsb6HDObtC1S7TdB9ZhG3kfPCvOUg+Z9ylcxLZs1aw59F1QjxWa2kJyBDouu/
MSy7Flf+8S1zR7BcUlSzv9oZ80rSX4FM9UjLShewOIwO3lMw+WxyV3hs4WnzhtPL
RJ05IJYUPAVAmC4edKcri1Ye5/sceUmO9II1brgkICdt0Z1XyN0mjxxigyrZj20+
EpYf27ijHiW8oxf7pqWsgZNpynTqxl1Eu/T7ZexneCUsGG3DnshkAFt17z4+s/pJ
Dlt6iiFYYshTnrdGQd7VClIDau/3PWUoLivMnv4jp7D5pdIaM0dAUo1ylHQlZxNk
pyOmVYjeWjp9hpECeWqFuNlQNFkqCqrrBt62n6cT2Vki4qqUwoCyZYfKHZzEXH2H
NsSiWoRwouxMA8hnrZIN77fFDGeBh/y9mik+p2pdQ+L7U8z+bA+ZhzfeQxxQRzK4
H7tCcHsV6+BwXsIESKMKX+wd5o4IAZhxKvi96mXLyDkLnouaYtzJCyrbwFpK6r4j
vrvGC7zrEe3vCil9VctzQ11cvnR8utQcOwsvUO0XyMvROKaAkpEHQcB8+RC+LadB
t2t6lV9bwKBj9GUZso/boeg9+J5SJpeVmy5Hdo4GZUCAtpLMIH4MkCVQUInpttA8
RJFgThx3Gb5/03Y5gJLknY4615pj+gKo6MWIPBpgpwFVgd0Xp/wqysVj9GGOznNa
4LNoK16tXNl1CtHvSv2fFANHzYXI3EdmFRCIJ7idGWndeU1YndL4IRnBsvS5j+4g
QWlx/mU6k0MAirRwk8GqhfyNRQbUZllJEvHLpN4qjT6mY6qPmlRG6YZB2qnbVC7C
Z5WsIinx2UU9tB5bQZ7UoscBSzHdzxGdHeA7ieaCJGuAuTAhR7VVp4GMt8TpGyQw
Yz3Be/uFDzzrvW1F9uT5iiHKYn08klYr3CKj17QX2v474FV62aV4cEuh7xDWweY1
EYuKGAXplFWIVwedA3doeOzPqgpUletQiQr7EVsVSmAcdZ+16AAm6pJybK1RgI81
6sbblXdhcVcF6e88viMDB9Sq6Jy9RcIkyaUB7zOaN9hc3i6kkiipul6UK9iFDh2Q
jGBM+MtcnH8y0XkcqrC05xVEtnVejOWEtd6c+HIyq2JRP4hMxA9lS8i78vs8E0Xe
goPqyi3CKQLkLIXqvOw24maRPYGmYWWobYss8D9F5cTzkPrgNF7Wnn9MWpOqKgi1
OC2rhKyxMcEHbWU6wfPeU5P2K/C2rrIC33/aUMJKEoEQGusJjPigG8Wk0qNtWXB8
lBRMscIR3Bu1YzFkqXOtnenW1FUUghIolL8KBZHhMDjzV4zbPZ/Qa/aJthuuGJCR
ppfM+d0XwwrsPMBibPwDoqwmIh5GBhAd61sGQJCe3R5BkO71kkHgU9RGQNP2GlUJ
5hnmCB/JFx8C1ZvZMXYo1L6V7iS0g1laNYbFg7IZOVFzNkwEEqJibHyNGsbm7qtg
R4TmVjFOb/nNvUZ9bbysq9dZbSqiE6Wkt/mcKlADxAa4WxFREPAcdyI+OvrZqkBC
pfkTDKfskiLn6riOj+OWwwvINQ9OEiO8Ys/R5WeNiXdPKmPWYzfHtEfCK7syiCxS
Ml/9o3HssLmsuoHrje2epvrt6U9Y2P+Ppobl+Atg2R9/zCPsemwilo6xwF5LYW9p
CPfPf0BROpVU5PzUKdRnbGKaQRgH0A4U16pUjM3sZFfb9+QVmPAJKtCWpsfb6/hu
mfOfnTlQr653qeRc5W6OONX+o8dgqYsXvi7+fxqKZZQVZY6e8cLHzHIB4lBX7KaI
Zvi6OZ+RrvalUCU/LDM8Ms5Auf4DkfIOuZmZL5OhMmF1MeaM2ot0+ABebuUT/1bO
ayjS8Smx/1XbkLZx6upq9NJMf+o8YBblLLIBbOWwn9nUd4McmWz365H2WqYeHtYK
ll19tywwyQyjFnp6FrMD1s3+WsjPxJBnBJqcow6sGEU/uHhrnNzM7G85H+k8qx35
qTPEwLgOiq93cShmQNwL7SIWi+4fD0LZAB0DNnQylNJ4Im1pGLa1rqWXl6RJI0Bb
5eaDYLASpG0y6UBx4EUEJN9CLDYQq9d0i4wvlENcAC60cN2aqFdFrau5tmecl8Ff
ZGBsDgwwat7LDTuSt0vhf8/wBMoX+aFIOiLBlC5CEcwrI29BSJuFFqLaQ1agOWa7
t1JUDd6KrQM4LF+iTR5B9oA8ezTYg1nc9JkUKpo5u0VT/ncobPXaW+DPgZoBbMxQ
hSgqFaFztGfVH+4exVfBbf9BbSV1+5CJ5GeabQoI7vX1xoYBt3mDGKfblvp2LirJ
6BGtDueUShuamhsojuQQB/n4lt7stMDcGoAuJUQ2Ef0zjn1VeK0SPHB0/3uI7qCb
ejod6g7pMz4CmgEmSNXfRoTfRhdeEzbjmF2+JH/IWQze+PCsYPDZYyKWZV6aRoDY
/rozAPP2ArsJsgDcICjX3gg7scEt0KgvwOIGxkSgH7up8u+M1m3zeWWrqn4C2jmZ
HND03a9xzBv+EijOR3/C0ypnmd5t308C4HjKXVG3rUPqzklSqnCurUo6Axv6TWvu
kaNtGDCXiuBixcwfpicR7xyNqp/WO5gKNVSokfLHeWp1XT+aeq/jisOCjljlIXne
gD/RsimxFOp0qYdpLGzunpzSmN7UskUGW0k0jXGPf4I1yzhrwXkQqUbvqMwRcSWm
P7g6/lYFaSQ66rCWRnZsosrsL7Eev6+7UMZJTifGgrg51P3MOUSlt2GwgLp2MMpJ
poXo+Dzalak2lR/nfF4uDLo+M6AMihjDw4yEqaFSbWCWC6mSOGbXew4pGoEu37NP
QH7nIFKlXAsvVN/SReBR+QOisH+TQ3iRHfgBgkm0wURRYzL3wiX3Ns5ZuohWfH+L
x95dSlTB5DI7AlrIPviaN2JYv8xs0RaoTlLIoNvM9BUKsRd9hZqGclMmFmxbKfeQ
dZhttOlgeZZotcj7UTdaLqFq6u61ZSgPutuKyQ2cGDEzOnGyU9RkUEwfRJYNNWBT
4k76mYQJeID02Q+O0os3EXNv0yn2YBKcdi60jQbaOpMr0gqNsyy/GIy8EWDP+OLf
DTadvZTvaDToPgwqspMtuHhxCSFe1HoS5p2UEFImRst0VVn2UVFc0do3dnoxG8Uz
9bovOxU06ifNl0vT56KkcPxv40vB0vbafAd72191qKhGH/g+acuw2aqIrfd5jCcB
ysqmCbD9Hzt9HdBTNwu79je2+culh9EAZiik17U7D1ktj7sm+azJMAJqlzp6Wrsc
X0ol+sSff7E0FHztQy7H+s/Drcf7vXJK0swxCEAhd9+iZHxGjiLyNa5EpPfLSUqP
m7dBLQOWcgFdGO2rVCmgFjAr3zZDB8ryEMMj7IRVdpkrpbqHJd0okkBy5pjcwNyO
tfkll//WHWWb+MYiJwgBSiS+TU+OyOwjX+vRqVi7gwTbgI7IyQy3a4fMAjjz87fU
X+GiKAZ7C6Y1A5C9OUUA0Igyxh3/ezVzhiL7GsweRAdQdul8K7GR5Tpx7aXyC3CE
c2Isb53u0prS49tUm4VF99jfMnoa89FuP5R9ZrOs6TDVImFo9AZRMGFJ/1X9ywaH
n+Lyq1Mh/CCQT0Mltj+O3Ok6d/JJGU86SftM5Pj3vUnC37BOfKqrBJvR6II8EWvS
QKF7AOtDipIjGe3LxGGLNiJDTwPQA/e3EKMheHs4Cnd+hQTvP4EHYiq99FWqT7vu
oYxfV/L/jhUD9wzSWE6ObAA/+EP6hlsmcyLZqwT2qVQq9uqBrKLT05PXYsgMzG5x
0qItZRRNTawl9i/wDph+KjaNaK0tZCcpK3J1CIhH+lyzJ5QAW4yeHZoe97RJP1AV
bfe70JN189PdjA4ZlYSuC0+h0+ZYLD1Lx0c8wwkPZy45DkRepSjxiLGdz/vN3wAu
kJRXelxW5h7u/ZXRiL8py74Jcy/YNFcchwjFvov9pbTDb7nETkRajmLfyo8Mvwc1
l4K3oBbXBaXEi3VqvHqYvjKTI3aqbkn7z0uXB9cJ0uuRVdj8hAsbhqg7O6SlPWf3
+wXtccK2YGFVGRNOSKHrfHV6jSOmq7Dh/S0grVYvAyHH106j8Q7PrKgUrdmY+pgw
oVrCBXO6Nf0lADCdZJOHACtjAVM9KZwZx1q6l81NCteg/i01EoDbo+U1a97Hv2GA
6nA84UNceaCqrtTcArG1tDLpMRxel/10J4VE0tuhtsyOdHgYwm2NNu5SVW0TP5sJ
EQDMF21+0w1h+g0y31QjS3KRDpzxrEoMVbMdidokd2+eAki8lIJgNuw9y45ZzarC
3+rx1maNv2wUzPWXxv4J9U1WWnXxB5C+sUgV4TFeYq2ErK2BV5pkw8W21Y0oEjgw
4S82bbF+h8TOVw89Qc5OB87bQbd0pcSniLJBibSAlmwSAhMG/dmRAzPqfAtf9z4y
jnrwL0KP8r1XVDzyuEAhBPOHnEpahJbjkAI1nQnxWXfm1a0r3hZRlCxRKKHq8Jca
lr03TY1FlTDpB57TodJLHbt+hUrl2KQpX0x5r9nfqAnkx101WL9pru6BM3q1edPr
hqajBGxcXdJ/41sEL6pyUcuT0sbf2L5MgQCQ5dT4zb7eNxMyPdrDtjFthJUq2Xuk
E862bc8SoOExXy2OGyT4naUIfQVFxD+CCsOjzTNFZfxoFfDPFZAwUczJ9kHOXUe4
b6nvQh4W9P46kgYCE9PLNtls+NFBS6P/OxuJcn64GVT6heJ5Qf8+s1L/EOdMFFGA
CAh0iPMhds/ZpSa52+euARY0EeJswQqawEAnxT0OwRQNWW/vtLevuQRYbnqvpPpF
8d7hzrbGnOX34kEgrQ3L5jH/7AXabmmNRD/WAG5nkGPQ45hyu4GaYv+EebNYLaAW
aVpt2oEIKo405FGWgszzbmfG9ITV2hcbaaePv4yg3g9baZynE3BbVf8UHYNl9+YH
RsJ0EFEajg4tokoCMJBQRURJEYIb7VcugHp+oYXlTSzFOmMnECLxA3zT6B1eb3Ar
JO/QoGkn9wW5911Eq0ZnHRkZPu9TA9TE8KyePwV/QsLARL2j6oWRHw4TWhOyPooQ
059MaJPS4G3sG+vedkrhoKVffxN6LPc1TomBXb3WMAjahiKiTP8WyCPxuiPBmq/w
PwAo5oZXvwW53QlnbOC7oGkKdbfjdpWxPuz3h5MGSp3yIHkrAT4KTg4kE2STtKol
PwB/wI9Z+hyGDJ+DMlg06H4Yq0rNGMM9HtWRJ3PLOBk1rbOeBZ3okdTsHRCcKVJz
SneCCEbWyXpax1lF0zQlRUR9Q6xLDewNOpyPPfTxP2ERv/e1i0ljwZqnmeM/03XL
B2bgu3Gr6PXBL59ZZotB8CKLXfDBfJ0sOLf/F7MbchhEpqqpIyYvSlV2jkOerqD6
Nd68MoAdjD3F8dHBPOod/ybscNAt87O6ggoBDyvZPEvkleeN0WEYEquvbJiBOwNG
6w+qCdtVKhOMowd4Nlm/Iu8NCvb2f1P6rIOgjqB+Y851EnAxo27feRPAeb///k4E
C1xXnmBfnsCUSrWOeVGp4zaHsBvcLUBX1YAQvjrH8nbj5pFXoZ/Nt+mFGc9WqI4c
NP62tD9fBOWxfjt2wkkFgCVVRNG6aOHrjR5pR5qeML4y6HipF/BNuoWdNC+LRMVi
SG6luQW9TPk9g3rXsyHYIhT114hclzXzBlSj6DQgUg5SmyfP8gSs6rf3952npRXA
1lwcmLZLigJIto95/ZG2vnaNyBYX+PsvTCYJFGE9SZTEp0RKoRqJF/AUBPl9EhFS
Q8TUTW08RmCH6/lH7hh92hAJk4onbQLUmbR9zNpHxWj9cXtLdOD7iO+SeI+P/sIy
p8L+d0iUTUBqZvA1jrpSHY2DUiILQIeC+8imT/N8/ts5vxlWrdGtv1a/BJv31Ei4
zK9ay4r/AbV/aTXlyxHSwHNMvz1hxF5Y9c6z3mySDrHO+UmUn+47YP6HE5GMoUgP
v1nrBv322npiEJBvWExSA73bItcLpzj7yETHptBJrIjAMOdxxsFkraehUduqU1MN
19KyZCfSQAxX+Yuj0VUw4bWEsvrf/qFCGHsk28sCJlQ2XU0K0/ea5WZTFyarGh92
G+xvKVmuBS+Xhz6iDyudqPeH4Z3uSOyeI8Jm4in8AarzTIqX+HCVxfW3NzgUhgJu
hIlD5GIs1S7ej5/d+hSTUzIL4WsWF/SC2QGt6eKv5dB/osVyV7hUBMutWg+Xbd3S
P8s8/9DEY4/OJeW/5mm3aI7s+wXg1DjsfsIIZmtSeRyrbt/p2w7/KWMxifRxl2LZ
eYw3lN0m0HDPQnxxH7Wng5T90PYjVc5av6KdHAyvWNdx+xaO09WAF36dJmiuCM27
N76WEr50czY1PLXU2w3S/hHRCmBtY9hi74Q2LFN+HzKDDiZmuSkxBnqVcrsT+XSt
LKtRuf4DCzg+753rVjdEOv2GFlGG1az9DELs3gBITfxHJi2XRDAfWK9xFa4a/oFW
/rjJrYhjHylKUzAZd58p+uf+UJ0tV/6DNvg0ckmY4EvY+7ccZhFQloALzT83GUxq
HtsrHiwXO610mMHeG/QU1exNWjIG4HQeXNhLMSVIUQHRHuCt9EViASWF1vmI2Zx/
/6JMDll2PRd/Q9ACvzUrGkIfA9Jq8jdv2CfpW+g1j99PqRIVvQJTTjfrmpCeSGXb
GfJjoItKeHGqS59E9+mt47O5dJBsNOOWoG8nxdGkHgms7D8sl+3P/JuQshh53gTh
VAL0kHId/FtKUNBR17BfmL8AXbw3UQrl8FqHs2/WeG1k60Em5I1bKy5BkDNQEiIT
E/MOZ4vO/zHMYMt8gjBYZC4RBq13jfaWO2HA7ukqd2G0NGJ10Qvjn5m1yDaLGt8K
zzVGIkVf/5dipj5JYmzeNLIMQkB7i9saRSKcMHxVJtbvord+j8l1vb4z5pQNVHbe
qEJqgnq9+yHMLbER8pxZ6JwRZPwq6sa+l+/75LAWnwK395BPtKiEpdkFzwa29SiX
fHqTqvo1mP3Yf7Sqwh7Gx6Mb8MRKG7wTJ49DEi3fDG0cWnp49y+wKr0/1R/Xu8KP
A1B2DyBhagUTBUngvJgdhw4eYA94HeFm2wFL8E0LJydqioMFYvVTkSayGpa+Qh4t
DoQoby9iw97Hi5z+eevSshjW4H2961hvuhDR6AtSuBIusPdASECmprwYcmUxqVZk
+acGY4VOgLGLOhcfs4dvmYN0l+rFWW0xaTZMWRidNQLTJKRaqbx7Ssvxrik2dd9b
9FzsjAG5InZYdT5I5Ovqe0GfFEYeWPs6QHiUiUE9UfskejE0lW55GMTjURCIyE/I
tZ3JXH0L8H4Fa6k4k+BHc83tyQTrGn/0OYOlE2JfGliTs3aQ9WdT1GuBQxzD09Qe
YFbOS2e7ee7Lx1Y/9Ypvh3MhaVHFak+iPvmnN0QK+aFlIlM3+QTCfthW+5Rd+jrI
RGaRu4FNl2VoKwN5LVG/4RrjBu9MPe1KZlh5wsrc7A+QxQw3WMpS8vyYW9q6YyoY
h39SnHfBQqfkT7JwHWVNIv5bBVW9HPCPpHavIPXlzVyFM+SRbAgWKf2bcSOlwEgk
rdSqJKQhZDYYZG4AiN1W8wzSmyVBWzf0KEB1OIwtM/rINP73w/qB4sPJZZBUaVoi
lncLQtMkT9rBpygLX6nWMNEfMREZvrFquz9duXaXBig7wuxIc/uCvu+Y1z34cV7c
N8x2bxTr1qCQXgRzAZkYFThh1BFyGv5n2o0vxrSp8rDq6a9phqeIxWTj3bglabr2
wd6qplinPGOn0MgEUQWECIuqPVog6B+f/iht6cTJTT8GqtPwo1wnXJxauiV1t7dF
R8pE4Pfwx/YmnqSeOv6T/G/WL/JgIK5N7vS73/20WnFV1EWkXSOtwIohpVRbtcep
6krPJfAfwnoqT/0S4pdYEhqz0XXeojn7J+Z+25XAO8aljDXzNUu0s8vpc4inMNfH
L804dUIcR9ftmuHyhu7dmpNkultHqwTm6urjD4QZgag9vsJQbb8gVUZIFIOiac+5
LL+LVKQWFQyXZf7aqJHZ/79B9mLO2OmkF2oVo76ciQrCgp45fkoEOBir0E8eAVkr
Sg9mw9SVuVxO/e5JqeRCIW1sDQlbMfWVilsc5MpOCQMT9bBnBz4XYlySZy9jora/
lSiETirGzxI5CDO2e3iMyb9lXg40bppuLO+6HZ7k7uUicgQ24nJPDlNbad7QMxBD
Kp82oQujSAyvjr0U1JcUczpz8UIaoq4FpqpKkFaxmnPJTn7mQ01y7XpF0Bgw56Eq
+HckKOxeXCEFDiL2MBzon6rlGP4JjO5grqws7qmU6+p/nKt1FS2GRdFxflIWvOTR
mkbUDJ1fNbE30X0b1uKkLLUh5E1vAfn7CUqKnIiXpFvQKqaMhmPhg8Ap9C8pHuhv
9NOv+Z56iKFKBKrSwW2Kp/Ol3qtZPpwMJeolDLJPd1CrUoerFYPoSUZcX8LmuHGh
73uc3CBk9wheEwZTcH9IOM7dXW3ahFRDHWYPLDYWAOPo0IOfR/ZWa3v0juNNS8Jv
NLn0s3uQVFtxxUcXlalYxeHqTadkmiGOR0eZ9il9VRZpOHHlQDf0dwA/NtaayddZ
6zPxNvnSTmgzbpPQ98P9717aseXF4M7zt0JBrE1wbI3PF1/E8VUse6PspHW8RVST
IOqnGXALZI+yjihc6R6u0QnTah3r3rjcX9a4qdqL8YNFrKzdioEPnKXulokcdFYw
vJA2Mf7yTYKa2yZVqs4xswEu6m04k0XiVBKEOIarW/6geMSmSTSjOGbdQzHzgsHx
Ei039zICo2lDRnnJZeNllA9ev9dTZwcNCcLoJCI1iNHVLg50Ntp6hHFqElaOCOX8
7/g4Yw8aHb2hfBOA32zoF+hL13bO5RJqPGXD678cv5q1wH+rH4Uw4UD8sF6+++mO
xulhnG8kBWaJsO09HeJzn/Ny9dMA7Lu81dbDyBP10MZxg+apzRfJGKjj1fKadNYN
0FF4/tcmBGkg8VVgED2VWc2GJJ4JEcgE8oS46RsMWfx/6Cez9Ii+hpX9R/ad5rU8
46O3py9EsBt9JqcPQT+gKxR6aQbjMysKmbN8r/sX2e3sgvkAHVF5IbgRo4sOeP2U
pbZY/FmELLBMVXCJo+tP9wIYIjxzZNfLfYY6RupYmhVr7jiEoiMDXJn/xoaUkY3j
030XQzDYhCgnFstibwRiPBaSuBJjYhuk9vXeAGjBI+Kurjb22EHNOujJCbDZmYSY
/XJJtNQRcgZGdR7ekm8UXVKeIviWB+QEbaPRIEoW44EwbyZTJ11JAlSN0+W/XMXB
p145Dp/t785zw1MlbnenKWrbF9SM3YgW1l8H6IXiWd63jZc+upN/anEWyuokqBwz
nZQmZI5iYXfvnFFnhVWlDutw9k2A2YZR7MV4YYrMFt0Ncorztgrhdd49ZfS5xYvr
mKk+geFH3dJUdSC/5bC6tDKz1qQrlDdzysgTvl7fP2nrs8bz8+g4Lk1Ai9fO+Avf
Wub0CT5jwT2YmG/p+lVe4d1G6OajdmLnefj7IXFKXVtq1M8F4q9X0IY674/wB90K
sOJ5ixPpg5/pO/D2BPigGWjsFGtuB557FPb6Gp01ML9wxN3Afiv2hcOIhUPb8XFC
TtwF1ua0XSA1+oDFIABfHpjRWhDoWbnfKJs+nHYVb14rrIZ7+MFHcfTpxfwSmBIU
0bz2OAXUeC/RaBp/avHmz6/CM4YMYsiaLUXxr4rgOjNPYKOhNP2Jvn3apC4MdN8U
j+DvHI44M6Bv9q8Ps5VGxWINOzGoD1fGplp+vgTp1CS7SMhwPZEb8aVSrNfNRzLo
IfUBUOxwz92SpSGVtGLATW3Gm3uhEv1Wf4Jv2RZ2vbPlNlTuGKM434L456KL9e13
vaAKywk4a68g03IU/5hHAnF2WdGdp6QvvyXSLdqEiZIaI3WoIp+D5cJ5VCsY+zRv
vCB/wjVuSlfwcFlqkycRDvrOw+wbTfureXTp/KkrfHs5WekTXuKsprIh2pLI2lQQ
Gugd8Vz4xjnZF9jDBZzeq2l61MHqkD8TSOJCkHTf3uklqOnJdT8i084KNq12Nqsz
YXQohwK7+0FPMW4ou3bxiig6G/D7HRXrcyI1nBu05vse0lH/QNMi1XUOxEJ8jpBn
741+OP42g74r9VYwIc6WXNSwsE5AQ/0L96dti+59mPTXlS8DXEFLy5aUi3eZgdOz
j7U35043S0krDlwSHhmP886GyBeaF/nJtFXR9CH2wZzJDKeALQxCmPREPp01ZyqI
bFW/pBn94eWzHoupJCz20VJTkjtP182K+A9deSipTjFyrLaSr/lE+TDE5i0aeT6h
KjrAz0lYLyngyeVk8nfN7CMbfCxejnknbeNKHIqq7mzuFCAICR6gbuoMDMk0rvg/
MqT+4fBccPfTio9bOkadrS+W9fDvfO2zx6EoTvQEPsAAZRwk0C1UEQLfhEYQjPAm
CIVgbb8Q+pIGl8pdfTvRHqpNEgYQoSnDOOsvtzoryWWs4T4Uqi7NSfHyQCZZ2vU8
JA3A3f6DVoL7BQ47vhfiKaQy/2MFVtJS0MmGZQf3ObEBfZhfvgUr12Fh96yxLXIf
HVvmApnmnon2+O3SW8bhATxWYQJF9Ixi0lk+m0L98dDEChZ2ojyLq5tE1CGqqw9X
FhAcuxHQk0pqe/WYsfPC/1vfmsi46kELJyUy5tx0w+o/cbQg5Fk5JlMh2TNpgeJE
5KssfuHugv+apoe2//Cx5CziNBNwp84nizsYMdJGPRhPRZiKga7rdGXTJgFoWRaG
DwbsgkdoeH3a5/n6PsyWQDbiIa+07gi9NYRwFmRBNyFUX8vdSAIUvT9B5UCgramp
Aq8axabfTityhoMa5Hm5vW4m/wkOp0XfBzIT4++r/xLhkbTReYUx1MwhfxABjiFG
8q5EJ8iN+C+c9ekryMr0fvjPfYZQDO83VZGJp0g2+S6jom1QwEbFCI5ucUkG/vGR
LOlYzGFkr1hP4xa9fQgjDg6I/tJ4hxRTt2oK+Ld75DxtGNv6OHn5VcJB/tZXPdMw
xH06yUNz7tlAxh8nBYLqsbfy8/zrfwu5HtVUM+QLHOxxMXIftdR4ZKUc+sahekW1
NBO9NCLJfU8coc99fJFrAbQ3r7Y5/j+hvkgsSG77ZecUu0iOQDJSweCBHhPqqRsZ
Rt/z2tTEN7bJPt86+Aa82sf/yOnj5rcF+KdYi27+pVLtAueTieZGYdvb0F4sKWoH
WfDYIm9CvDYgxdhm/G+pbldrQc5KuJxQkjnKXnTCQLSZ3i3Cw06xMf5L8NcConeZ
J2s8sc+ALjMCVzeZRPI/caf0fG+XuXFlIi8ZNmyEI/NMqlSZmoctR1G8fOb4mSxH
GIBfcTt9QmIPEUkCTNX3G6UX1/7zzOsBMmjZP2wsAqyHBOpbelVTsY23nySPNARK
nigWppXglfomSx2gTZYKEWrHFzQut5EhVsqEukMr6gNHMmtJgPbYvljdk4QKHWYZ
pCxGvB8Q93xQ3JpddHbdq1clQCnCrf8r0dXu0cEyAb4wftYrxLsXnBSr8HyQlsOk
DJR158v4knbVDSK2U+yMhFOCQpXLWB4JkXqdhS4uBC3DKMtY+mU2pLWHLVi6Zjv6
TOwySS1hYalDIPaZU1uOhXMJDSld+7+UUeICp3hUTEQpWHxD1T1xNZXFJnT2nmnR
XY6NnEaBfIPTwCAmo8sIsT6bSBvVGpNuvwKAS0pO0MTi6UTag8PA+M+vdAZlTpN5
KlnFlTdLxtHdZ/2WscrFnEp5lAwDMvsJ70QGC+zh31kjnfG+BLt11gt/cFF49Ibk
jrIY4vao1VZeNmvmKIcMUoXju+d1entf1ZxxL9eSG8hX0lp0KCCg4a+G4VXCcwu2
9QOaGv06V+hYt79fY3hOtVWM//AgilRkhJtxXvcXgGrUq+SEWs4Sa0JwFXKpnPzW
KygWGF0zhknyHmYXx0vF56R6CFKmJTPj5wdUJTy+yaEWtebywdkgTkMrE4Bdn21G
CzThOEh3AtefEqIdt3FBihdHIBocunIVMrAJ1PggzYO4Mbs7FpT7LnFiJFmyHw1U
q8DzjwxfcJcsmqWFo8TE/kQfzac4bc8NgDXS7Yf/jcUgFNH8cMi+fkjR3V4c4FGv
pQVu7Zh1bVSmJpmHAb/D+j/UXRzxYFfWT66321glbNxBdfWMcygyFVQ1awD+2e84
cA0Fo2CTu5fvXjSWX+f7WiephDhpvgLcmn+Ul19Lf/CLfJVac0Iq690qnM5ZILrv
i/z620xVA7fSJMP2f+PHs0FTPZG+JrK82c21RLokFO4AVwaMN6K8R/7pPZlkCe31
jl2A6FsYhZA3E3/jlVyfACMmTxFbWeo4D86vdZSVEMNvI6Q7eyiNht5qgkQZw8eR
26Uu+93Pn5B2tQ6jQU3StwFzTU8vtuaztaIYeq21qdjetuWc2HhI+I0PagvZxUpv
U4V99Eny4yRhZoSymqy7BOKqX2sd9xmxTB61XZbevO+lSfXdHg3ZVfkqkDUJ5SU+
yovVBSm4+UFPzYjvWzgcKknFAmdCnLQEYO2DfyRhe8Sgjm5cvpXw+IrCAuDrX7NP
Po1pf6HmrJ0mAhLB4ZhCW8ajGP15K7tH/67bjQw/ESpd2WnpekpsXcENSSpApEzg
dFtt+5MF31Q3lJNyW2pF6zYKtbo4HQ4YcfBP98LNLaWZ6c+5r6XOdyPbf1aZG8AY
1qQt18x7BNFhndx2/5xb4i05JrIbm10rBq3GWRwC6MHuW0qzlkgAccHm99TRV2Pa
Iu+vqUAQvE5WQzZhtlp5zrRCQfa3K2G/DbWxY3pmp8EviVLfUwYs0nLcCgLTEnbv
iBBzhcphXDm1+27StTSaoLUj1fR3+AHWtgBxm2ljXTwfQXka8NEaxRnDoabFob6l
+F45hv3IuJJsprNW1BNero1TuJgjqe47uEty2GphV8hxDDLPtRA5b1cXUfFXeS53
ffERlC7EQqztRG/DuZnGIW3hWWPreL5wszWEGC2A7L6Pfww3MAELd+V7Idqh5263
kVjWj4zp2WydpCkBh6M1JNa7I7EYRcoPXUxu0enlIgpitsDbUXursQeNxynktYB8
2F+8IyUPxoFKxyCGvCMuAKHb18qA1MTTfQF4gPrqYVQpLHSbAX4RPGJKMPFFgNlP
X1k1g9tTrb3SWapWmRxhhbc9wlyyF1k9uWs05xg3oo9Tm8PChego1j9YzlNrOnQE
kJqWr4Tv3sc/TnmUx7fPVCaYQa29PlG3UkAEKSx6FVm9gKd5RFzTzhlURyv69tQB
bArBAY32QL6sJH/mkdudCERbxvCRG47DL786yDSl8XUK9dW6Z1RvCw2xPEjYMcL5
+Hzfok6k1CnmqjpCCUzzkCP362kDmSfLM44c+MWDOMmnimLvBGsTTb72HTrIo3N2
vzIaL7JzxVdsswoIrOxmPeg905jO3BtQnkEIFDhXJMNFTN61beXsbdfkUwzVUuOC
f/rPRV+G5SKllcn6vpXUVFQ5NZpdAu3yTVE9134XrDWn033WaUVli0Gtz/SAQcmP
Z2s++dfS+4EiD3MuOvcd/sblM9WJLwJ5uENGudLSi8y1Lh4Fg00UMtM3DmOWr27w
9of/C8h5NtSaVnp9giX8WhOu7/Mjv3h2iZwPDZmTEeUcfXrMgFK9zN+Uqef5vDnC
pnoMXNc0dCB2IltVhRJ6ZQX7LkZYJR0ptj4LUPv8krzPpA/V8iwkPCT2N4x82ABS
2BM8DaEt5WfgDz9ETbAmiwIK7Rw3Umbk/XyzrdhMwIzf2zptRaOS2q7OwsdAnFwi
iRGBpCjJMzIsL0XIZdgWviWcSjRz4m5esTuPfP6YXiP0YqueToQSQLwcYX4Bbf8y
qUTkhMDk+8YzSccG/eLAHaqOQ7XQgrcqgQN+/BuRsRFrleEAk9QIFaIH7257v+sB
ku7EmM/q5v9cymhB6WJ7/qJaLE0L40BnEBk2XSv/uylF3PtBNFY6Ni/HHL4Ak4TO
JBUlehMAvw0KQULRd8xoJeLlFjjWyCLR1gtgEvOBybKWIDjt5+wcHz1Ien8WHlD0
CUCXN3Nt6pxjjYR+n3hEaeJfOCWfhcJH90AeTIl4nx1nM3lnJZ07J2d5arGyz6Zs
rg3DxBcWOE9ywLvdgKb99475B5KNF19AFEK4qTQ0J2TryYGEdemBgIjF4mquuPk1
gbTEeqEYV960FkuphOhoiVkFBHS+WDTVDzNr1qb5DNWzQVikgy2zQbGdAKwVHDGL
H0LHHRTrkG1Bi9VUAR4s2GkGjSaeOB+a7KiWfHNVudgp32ZsAyLUAkOLA/4CuHOX
2hiOrrzlo6QXwzNFRnz90Yw9Wf7GvM1Mb/FoF0UlJ18jYm1UGqPI8FxPu8l7T6rz
hT29bOcjlHJPxpCq8GxqpsWj2JANUBMYwG6tF4my4JarAP1tMGT0gKCel6N4rdo9
HFukftU4RRk+6oWKwU5IdmnNm1F9Y24Ksrjc9WJ3X1NoEKZuTEIPXx79vMWjIgV9
lUhYexn4o/D5YtXxvYDGtwYxyHyUNKkV+g3caQFqxuoKWH9O9BK75/LkD3hiaW5n
eKOUzGGkngKIzUnvSVc1f0nIMMaM5vFtcX4K9FKozdrP8YWVBzJ1CiYhY6tc5xY7
bbAsc1zQGjBoF+hrFu7KFyKWb3k0oPhLNbfePj5nt5tRRK+b5U7ToCBZeanXg65o
rU3gDfNfTWckGgvBvRxzkzpwrYOZELZC+rvKj8IsJuc7yvNbwpn9Nu2VZ7H3f+Jq
OC3CPaC2mu8uuJ9zQpRqMvn+CbNtWvLxcX13D9w/RsjBQtL5btUGKwgZXqL5Epo8
ha+icGlEMfM0l5NPy5/6VWfLn5qRv4Ft5UgB7sUDBS6UdGBuc0e7FGv/nC/fxSW1
GMuQAcUz4AQ7bRTo6KlGzTX7j4IT2TU683BckboAfD4Dj5RO8Klw/PjbaGA+TAHa
K4TwhyuXLqNJq3Qq57DbzXo4V6+yu3ZFbBPTybfwFNeeB14kV5YwfCyvE61wS6bO
FLyPcmQl80kvAKWujFjqoYwRouonQVg31FQyqagBWAMckdQgpINM2bjhSut8P20h
gSt1T60OxrJzbguMHq3slpm3a7js21GjFNVIp0Pz0DL69cBXUYxQEafdXLwzrZlz
XcAyWlHdRHg7DcEaV/UPOc+LxCNHK8ylmgdIhmlfc/ZGpXfz30C17THDL4AxpweC
w6lDSEzyo38vr+O5wqzxj9NYsBgqzZloAOVx/er987H/hW8wp1vCxiN3ea1Na3wZ
MoaUW5WiYgQsI7Kp8WumDKMGO8dEcPR9E7dpBAyRFVwIFY0FCCTCJNyAfZ2qiK4s
YsxGxBcVTRDUQWG71kWWJk7yZEH+Ya90VnLBNkLWqi2F85lETSK1yx5GlNAoP+Tk
/SQFoQtaHD82th/hpjdT6L06080+pWC+o+mxGkrKCNMzzOPOJwg+N0t1QuVK1903
BWLYPMiFBz4ZlZt43LODlE9/JG8TO1KEbPW1xFL87SCCQP2hrrHbqZS1QAUWxNUy
u/8GNlhOkYcX6MzgrOvLmBpP+h1BDyeUTVofAm3/uofgh2SyxzNjFxJ7jNx5HDNi
n15/Fxo9WrhgbV9pi3n90lXuN7AoDwZABmzU7OXaEAaD5dfYbFN+VmEj6zSfautK
e88BCSV5A0mf+elTJoJ6UMYtJIcROz9LijbEyZgRu/EoUQxqKW2sx3wISaYE5SmR
hYGWwtqAEtD2h+OQ7Y9IGQXL1bAqKbAJ2XBC+D8jzZlc7940a9vclO7xsyGuMIDE
yFegTyh0puS7EarjTMDmNTQ0sQbmZBjagOnWJSyEuzvTg2vSf+otWQkJGf4j0Brw
E/Xy4vD1HC90e8dw+OTKVlrgejJKSDNLWtKQoc4i/8ajap6qnHU8n6STUPztnP/g
R7PX694pGq8+1t/IjpT0rHpWjECPsVtpFSPg6rGaThHMdQzVIpSWtAe6JZnHOjHU
+1GBvziTAz7dRcYlAm6sHQkpkrmUt6PSmUH0I0e5HkOYv8jeRRoVd88WHBmPpD4m
1xpMHKqIniA0qSfma0fJvma8hYgQ6D1EhF93x38Wa4bY6Q/iAFIW8IWzQYhbSN8W
KjDDZeIi5iDy+le8l8+38PR/Y2ukG+vI4aFr74vSr8e4cdSp5XI1OLGVE93cLXrZ
0q22wWFke7zbvVPcVX9BI30bxH50YihxXXn3bTBNegLt1tY5Al7Z9z8VTujiICjt
5cRSVym4mETdSmWr1E2CVfhVBtd4JZMLg4icgTaUz7haNUMCvVwQb1PpxQpB7XRV
Se6CdwM7wQ0/15WLbsa6S2FJ9Lh5JtmfFXFlks2VHFdY2RnReTbhPabCWbA9P/cU
/Wwv0NdAhpD2Znyx3+Mv0wYUWVBSzCb7Md6+TJ+7wluvJAwZVAaUWJ9mUVTNHtul
/QM91PdYULUn6gS51tpBIAwqKn0kEoSHesLBvjfJ4HXXTdtAJV9YtbQeATkAjQhW
Dzq8NxIN0fV4uBSIXwt6Kku6iRbZY6f7wu+xs2I8ITKU6C2wvjOw7dI+UTPYRfUq
NlyJkWlfDB63BjlQlO/MXqtVMOoE3aFSGd42R8yiwo+DiJxVTQS0GVSdPdsYcmlT
lQVUew2V/N74x9V32tHVyCagdub+FYtSjFegGHXuPHXmai6Edte10okUoRdlQlOt
+mz4pFVaNvevKoTPQUzxXCyVaODzzG8PDmo4WZJQKtobGbnnv1ABOxLYgHzYqHkG
buRaNpVUb9qRJSMVvI8g8XZ7+p8lMybnM595k7w3iHhc7+O2GztBa793ocAPBMbA
L77R0nCmEh6Gk96WOdcpAfjZUeBKaiJWi7qtAVTpynIELXE0QcxlYdcEeOnJBmLN
uiHGlFj3WpK0mDgr+WNsQTReq1f1gFdwPIW5whf5okz7oYTflIfuD3KPCTJy9gZG
FKc61PfzrSYqd7wd+VACuUWwN8N6+V67dfE4CnZcjiLfz0h+uPfGN035tCV41PTG
+Iu7lXJIz+Z0VhBL1vNlbOzNFL5gBBjbAONVsJZtnN7Kb5cp1N28p8gXWoQnkVIe
UwsOeIwlXUzcf93/UG8SUCWvHNBmJr+cV8yTiKZOigz9jpmyoQaA790G6QZzrfQj
n7fGWzUym4Qqvp3NVs1JhV0U31hycyNP6U8cZJ+Zh4cPU8DNvayevRBN8cUVtJ9i
+mPYLMmAX4rEfvzpM2wPmhzctRf+ELmsA+9on33+FjWazek41wWVxPnufNZ7MGZL
WCRgZIpuvGNF0W/tipcdOHq+FGzBBGPWYAAUq3aEVeXwFNSXW4fIsuzdS6uwwXf4
bZWYH++Ge2s/ZASQ6vE+6l99zAbtodEh0jIDPhW9zzfSmsT9U56SO2oOWbiMP5Ny
2x9lMoVzb6etgm0HHAkscXp+J7xGRWUiVo1+tRBqI5NDBmv8P5dKTcy2fq43TT+O
VIxC/kgzbkkYu8ZKrf2Dgvt9URn8IfSebTlqwP4Wt7nNzo3yXBr1EROiaAHZUKsB
pHdRxJhRV6AdqB8x48BB1VEV4aNS8uLp5D1oPsqEH2p2AwtrqFMulMieWgQB5c3x
yIkGPHbGGNn+Q47FbHvA5nYWawaNcs4d3OQ0OcP1KNfn3iLjotafQ1YYkU4Ag3Dh
X1vieoz8eKDm8XMTob5/dLu1H/5URrp/9TJkosTwsoYZ2Ilcz59aNjO8PC01G4Bu
qUkbJEbPZsIqvT1am6aVbjy0W/+TcKJS+lKwNnzT1rRWupt7603INYJseMwUTxsb
ASZOkwU2E+gFqWffPdFpKqAOoVIoMVE59BsI4/sEaIsC2fR6YDZ+vhZClzkb8CHE
U2ZnEy3aFZhhaWjv3a/rLwNahGQvxCb7swiVzkoMHiwKGH4VVAWllUbBpfOdZda6
gBwTxBbk94huHAJ0AqFxHjvdZXCWQiVyQLPVoXryU+6qZRr3EMGFLQn0ZovrYQk0
iU8xMmXHetKcAAVTE0NCqDaY7q0febxfuIrtERYTRlemv09I2GzBHMAK4v4l8INw
MMo5R8LJqopOJwgBwZQR4YPg3se/xxe2TmTxZor3Fd7/xWXWIaZMnXrjpvd44Rdg
oGpbZw+E6rWPUcfzs9NtGVP9eIlMuytQ2LbORQ6NEbyEq25GiMu3SkS+en+Z+N0C
beFXSaH/EWtIBQ0JTmrvFnjLbVF4XRSMRzELRT/4j65fKM0WEmrNDimI4TxSyhmb
LQtZr/5C+v7nyYIVg437cUVtRIyDf1x7gabPDMb0h2Es/kfEkB7XKArwURtq6JSW
RMGeyCTcXd8Ee52pmf9NxMVaGhqCQ55ZlWf5wFhbYxEZaL3iTWFIr2wZ4mEa4mvF
ZDV1vQ19ZpjOc9pxp40EcTmdobQcrwDw4HU5iPds8fmPkyeLoX//bCiYvuqfGT2C
lLzClXhp79O0MAtOFX0eBDFoFeErUjDdv7qPDTpeFqQNpT2Rq73RW33kNIcLJwQP
ea7yMW3n1ZaZWU1XuK2brM2ID77sqy46hhXhriDiSvHNYO4Hq+93iOzRfIyHjeM3
9m6Lut0C1GWGjFtrfTluw95paHFE/uSJfe6fegk+F+LolbkNDxyRZNf9jRgJYLIs
Eb9uqlhwGmh1p6fxMvO2olYWWAP1p3wxLthcESDC1DP6o+XXGCoZKbCkuxMLO21x
04n02qKoAFBdrtUElV4ulW9u+r+Vt2wm/luXE6WuGOc1PMPPm95+xen6cLE6wxNZ
wCokTOLwq0mhAVSq3CUChvXuXO9RiDfZZOZltbs9nzGkJfH/j9Q0qXv/v0wSdgnJ
/SHxtIyQdpr+swIsnCSektWI9eHJtCAypLPyAKs6DhQ/jguZE5nlc8kRBlG9+doZ
6mUo+gY59/LAgTEtSxy3aHyt+0EbIRaKSK1EWm9/ivj3FIwg/4Z1zjPJOGPIef0t
Q8vYAW0Ock4npH+gzKETjzeM8kkqZbmaLe77wNvnTdwp5eWjJR6UzxJTiedk+VPr
2kDvB9KonQP8VUunkGV6lyyGVMdIEDLw77BV0lsrsX8wMe6Ls4tHLMwwYCY1gESK
S6ZTGga+e5VRhWzp64qYlMI/c9qFbDva0aLR/d70JUeKMZFyU8F4jUFRYg7rXLkv
jOSDwTlDftoyMhjPGqcMgJYHPM6miCsmnL1Qm7zg8qqweJXZPJKvaJQl4I/Ey7rl
xJv0OXWQ2lxXqFAsw5tl/yTQojsm66SuRkRPls9JxbuYs6jwcpNmHHuudBuyT/wW
7GvV9Ik+2m6N/xOptkWHgBNV2EtOqporQLm9KbD+WPhR7f1c5yHlUed/ke1jnxNG
HxnYchV1qzJ5Zs+EUFnsWOz8Qfu78pfBeuUZ33yXAcuE8KwPrikeXgB3I4QDd6AW
Skb3pXnHuys/+s+X9tIiZiFjb8jQNH1BWEhV97Bb7/ZL6UdwCq9WUv22TqHzSVYI
nziwFW6k81UomRS0JmR5S8YpUIeMxAYnunTR0zrkeRCKyNaLE0CwXYG60tAlQxJg
tdNamP4UCNZPPRFYsDrqzqZXjlcUAWE+MPReA/93/wAqKbTfXfsARlfmXu4cEH+U
u7WWtKBONtcoBGZecWdQT+0iDlLHGml790p34AcuKnNHc/AO0BDYTm1fqJILw8ln
lIh4ZACLBLUsZwPh7F29dSLHgZ0YMUFWw67DsLo2YtmHqkaXylPyKk4xi5YavEC5
YvjllVVSyElRD8GOauBC4sPtd5hEKvtHyhAx4K68orZSAhTYT0Fb0WuqxbnKScUy
PDzsyKrI+LcCehLV8PE3ux0HUauDLKCD+AE8M2+LY2ICUqW/esvNvLYoAoA5hWyN
dUynZOlcDR2DunL+Nz9KOcihFJD/Lf3PgNvVmHPKArLPsksBRateCKxnHRLXwVi0
n9z/HlYRNV9QKt197rUYiPrPb8uYKokkqGspXkngASeTG+67sXcA/jvRae0pBYXP
Zoma06uPtFahWeWETbTyqeqWQtzX/Vw4YZDPcVJDcqxrdjV1G6FdqoRr9kMBhWvl
CJbjOSD8//2QKuKsWsnfnimmeUG0cHf4JMisQAseTn9AEQBn0cSD8L0zu+BG4uCS
rJFwt9XSdlueyc/LEiSxqbZkLE/xp3e8AP10R+8MVEs8ssuJNevrCCzW5cGve/xN
YcOqhGQVw7Qm/b7io0HJYg+lS3yVJmfaIGu5DfLCNtYwPw4lBo+5iX7q3zEA1s9J
uNY7s5wRNerBuuvtnCdStIcjPdHrwxxu6aZmJ3Hx5uQWBB8LKbOo3embVqdjeCzC
DTZc454YU3637aMOgf7HTYX1++LB0SXGsAC0GOQXw4qNoP99U39WSrAFw+XiWIaw
3xP+SK1q9Jf7SRp9eMHq5zC1bnfNjs+lvA9kNsUzHjDIpGuiQWIXEtcKLzzPh37B
f1WDKnILJlCxk+39Y6OCtG9IjfZN4bf/r2GIzRd6WJQoCVaCzl7z8gAyHmQPOgef
gseWijyQjm2HGqjpDcaaBvrC+zqPzA7pHSha+7jDLR/+ynlai4c6QckcTuKOyqcL
veIBkQ3/tXc5vBIiGE8YnlXB6nXyHLVRFGfrmMLJfq45Nsh/OvnF9i9nAZzIiqbw
23cDSsu1NKSlUQIzU5uSKfMJxKGN34svjfb0L82QWI3Kl+Peuvpv0JcJeg9z2tVo
+KEsMdsWfbIQuvMKRXLSqRY7CEqBnnzgyEZbWfj6/PIn8nL3muap1cUttPp6SaX7
kTdpSVFOaCauk85rtLImVei4zb21Jf/wb7xuKK3UVG6bYftz8avAbLZReM5ir5HE
Ym0iqROThxQPYscmIqwi/gtlTiK32vJA3NeJAvf/Vi10YJT1A4PvzWMINETmsbeg
IvTF5/FgSI0zK4VOfpqCpxanl5EQrUZ4ZZSd/iiS10a6Oed7TZclLCO5U8SL4UVN
IjK4vTJsAk5072jmhF6L3a9byAQRd6BtkOFGEKNcijPn77jg382lQ2mq1W1y5iVz
82VQgCyYq1BLxdgpzqIzd32/2xmSUI1y7E9OnXf6WbI76vFf52/u1VjSqEMpUJzh
Wheiyo+uXBImxrYp3H7kTV+Ni5Hpq2v9tABpDsbMr1LBy6PMs45gdRK0241zyAef
yOI+BKYo1t+qo8XcC7pQcGODfc3z0kp016SIs4ZSvY0orpSOATNmb41SxbMLlops
/SQFzP+wsVCfhbmu0+yf7USjRAyi7bxtYmCLWddE8h/0BMyxsc96k/lTDhKQNE1C
2/cNB29cyn2f+8/6pfT5WyfSmgWue7qxlzvirWv+NMSS3GhrZKP0wX0g7I2O86zQ
qmPJshXG0lN1KtJDvAYbYacBIlL0Qx/ySo4Jr1QQjcCfX3r4mmEbW1vOm+3I+43u
ZjtLyRrCKVAqz5HwROExpIiUeffhSDDgtuMhmnFcJsPpuznFar+TQ83bM5C0PIxE
AZKgNQc2CcJiludKfE9PYgaOSF7Z8ChTxZe/1U2QCr+MgUp4hV1LG7PcQbYVUlLO
SXG/TDvuGD1dmyzjQ8bl/MSHEVwHc8iAJWgqqysACmJKzkmAigAhyIsbgklddA+h
yYO/NybdATRbBtYh1bjADSndX79saILrxF9wNSnG9P3/LuUZEFLq9vV9YM1kMrNj
QAyEWaF1jxYFh17tcafuSB0gu3DyNo38p9owAuAq4DYncK8WR0umkcetPd2qSzFT
yodEwYxfR+LLNJklkvxA4/aLUuhoo0PgnJo+ApoPdakTs0ooESe8NMqPv0ZTlmPE
HE859xG61O4K5TGtbctNtekxLrmWNChm3dA9Njl+8IJ8472PNYLC87ow48+376/X
3lu4MNd/UH4EmKqvOBevGHL2VrvlEAUetrmcLjZCzdicVJ7Qs8jlJa4D6dT/Cda8
TWDjkISDomeQ2fJVinosIpGTZkN5PsA/7hhA5BSvmDs7eKV21Gw9+0apNR3AIOa2
PZuNpw5HLl85oXw/9AwiUSFOSclGZkA+YlNY+Cs9Faya2J0MOflCBbLw58wyNpHW
FHVt6R3C3nzmFxr/tZTS8mWE6MUzntO6P7YFbXVMmNC1C/rAlCBadejr+7FTLxkl
sDOQPIZEegsGMK0yikOIMB6AwWQvgGMS6aECW9fnW36sDzOfvbNKffbQWohCH09Y
S6tBMI80SSyLDapMvp1ntbPwEsznC8WEoQWZLlpt9JuD9xeNcq/wAi/P/z10Tyxh
IAwlHkeGItInBVKbTI1XOmxZTnDvHADZxBedCMJiXah0TBXOr7sDnZLM7VR/4Q6F
QEDX2f0A8abT5NhzriblmwxjOrk75lNt5Qlys0pLUV9xVXovKUGNF13/KkF0sUQ9
+F/+Po90qwFWX1K/dsa1fwO1fzZI/2WFLFoFp0/5VP2OfiaHIe0sIMRrtq9LNj56
IBqzL40ONRLzRKhUS1CyrVPrBr5rHWXWG5zd4aZcYv6OsIqiwK22hGwA0ROnLyT/
kF8ZimsQYUJkX0W3yHuint+AxO2E9XKQTjpKvfHfxC8NsM8Iwk5QfMDpuhbdGmaa
nkBZoVYnDvRRf5HjBNfQk4NnDn4KDdKu8j4Sj35V3uCWxlAt4lm08ywXtfyrDDw9
9mbjaQv4aL1+NCfRMsijz4+r8tpznV0lyS/w2HrvBLh0kfDOR15kyJvDDKVT2ttE
jIOhD3j8DkIs7lpmtgKcfzJBYLNOrnuRyVuc7noiULsJoMnkDI5+sTpq+tJgJMR6
h7IqBuo45GJkWaBvBFiAVPgs2SFC7VbP8USsoc0SIFP2VjQv4GU9MBe8ur/NE3D0
9dJ4q8y1XIQm5Gr3kV6/Svdaj82oL87kZnWNXgc+ReA1C/zDxPAcFEBBcKgkuPme
wPffKvbORUOEUGmSvd7kBMAWcGf4rKodfi4ohbvhCwsfpruR4j+E+b/3dqEqCqfY
CUAYrKXwbKvj+JwJBbXTrmDdgouJD+TRYZQYO6Wgj4tMYG51klOGseJs9e1+N52x
/qV+q1knxGu9Kw9yrdYfJnjduxVWLaL1w/+xXbfxjNEcknm057+v5fY1J2VEfAGX
sBXG3vEqOeiiitaHBiDHUZaSftCQkzo5immB4/uMbq3D7/THZD9yti5xjMIT6U54
QdeejId+7GHIb8cdPRF09KmX4hoWmpTE1DPd0FqQZPEKz6QqNK4X5eVb3CpmEW6/
IOaQflRiN9EKp9zIXLYaukvKp4HIT4Q0OQt7CTuZPTsHPxmaeXMaaqLcqiEAPUTm
mR/ZxxRE0GYevMRP0doAdQXl504D0r7WfWdzZFF8BTV7h8rXOcXCiWbd+5nD6TZQ
CEtszmEHMBaPMbGdX9qUiK/b7ErkDWiUKedAlNfbgaWRgtDOclR3iN0REDHWZTV8
j23SR9wDsWMgc3ddT+9we7TeuyJWd5/9HoPPiLPSV6sJc7oEkvRNWk9uU8XpfR8W
XUFnZAhqwoj8hu/Cp3c7l8JxeiQvMAbwaJMzt8tVECVgl+3RjJ2j9by0AG80l3Eu
fNrHsTpzwK98ZQDA/I6wIgMF0dfDn2pbQgqy/2PaXJJZhe1D9+YP+iizwhmXI80L
umkLnaj6xckeDoOl6xEp/Prlxv2YpMdJ6pdW+e4886zA49NMT/udqMYMCsECRevI
EO417PLd8zi3Iso3RDVRBAav0XLEAWZBWY658yf8KZ1Bh7/K9QwiHSNaoh6CQ586
3dVYB1+kZLJBY+zasVrzfpGbka4VvC4aOBDF8VUnip62eUh1lR9rpzAJWqOxgHXP
yBCafuTE9E/lJlvvfWfyztMftaP2k3raEvOaXa43uBjr83TBtc38RqGILUMU4Hjc
p06weHmWodGSMj6n4G/zAtRTOSZRjDwNSwy3bzEcUZ1m8AnEFvWeoCjR/BKXeDlZ
MtIy/kn/Q5riUv8xyaXO/8Erx/BQdzfQC/zmn32w4Wf0tKDBxwLQYSELwHcunOA4
D4lKhWAei/4jpHly1x8KW+lBfu4OR6Pg/ULu4/E6BpV+tawbhitw/Go8JxWWsRng
mc3TTMx7mxg4Axk31Y4Gtqpvnu7y7ssW0bsaAA8FFRVAdsFO02kH0mLGAjRAYEVH
2P0bLW/AETsJdmMJxQ3KObiwNjUEQWC+/G7/MUwY+OptRTcZY1Z5BeSW8UZtW8Ll
ouFBJWLQHolPQ1v+hLTLsiKyPXaF1azHoTXBhcgt8K7d3UO0D+VPVhlr5spUzL8i
7hCBa3E03JZBXF3guQojIibcbr6/I8FwznxDYYCmgvhs76xZER+VdX5k60mz26qG
9T2eYQOiKqYPG4IgC6BzLM8SYAJUcRLxQN0JQduiOJVH+8d8mNg4KBZLWDDW9MxH
o7Uz7Kn/dvCEx4LRazkgt9AdK2gowjndQ2B/jVoxj5GiT26iwfq0HHML9OQpFZTI
NanThiXs4ZVjhUgLCJof+lV/NwFyvauqYmzb6h3WuF/7VskF3M3ZwbhRorErPsae
U7R9zJEOJrD3J2QXe/l3YeEf8xnB1YbexNrfAX40EgkEPytRFHRJIKsMg4x9sn6c
ard4BTCuo4zBot4NFRWYixQALg/35FxE8wUmCrvstpY8z6O77dzAmafK5IzMg9G1
v8ZKz93kRAez2rTXYMpgGiFEbaStjSPDjTCAvHgzSO3FzFj0JSjPAvGpUj7srXXG
hPBp2uFBJv++1Lv58GUDxZ4m39bC23BxhZ0c2mhoxsWKXPZogn7NCdSwpb2eOxL8
PF8EeeXPSo46rNMbFv05Ea6HtS8oalEkWTH3vqDMbh55Z9kh4/ETPtyoK+vltnJQ
uesvFu+mt+OxP1LWVdj2DOBMbVc+ogPVibyNfEjjkYuQO7vZa23GJH2Nbtz/SszJ
vuUYvU50SSz6ssq8ZDRphBK2LI9CUX2sp5FNy32MplfOmOaJlewNiT1DgdCY+7d5
/ZYn+AqKpfYHyCMy5Qf2SbyPcVdpE2yYPatdDmDhlFeb+mmgbbvXkYCATrIviDMV
bUt11KykEhRGqvVKvrkVujHryNzzMv7WHdb94UJNYHz443Sx85rK9uxSLRCovJUv
I/4pYGbx08Ucysc4pGhj9OEswTaG9sIv85mFzyodDN9t9Ofxh/9iLa9UxGRUB0gT
Dlzim+Sk5TLxgfV6LI3zHbAXDwx3cfKcqzm5ImFF+Ve7ar7t2Vc+DH3clOLzXOI3
fHBjYeeNW3LjXdYTgyuUwEnkV/NjbEvCS0TM1Sn+WyiNIqLy4ZHjeSVwjyCGsjhH
aBHL1R9F9PzXLcsSLfBEjnPXm0TLrCXlOoX0A5/LuUfccrxuQcnMie4K+Hw+ugln
A77ZppDgwJ9Iv3oIy6Lfyftump3+pUaXbF7k3fouDZ8hrqL2F8EJNWuTzNYnzEUJ
g/y5QlpUbJ4z2mkVvD9VOa2BXz5c3QKD0lW0uuw+UZr3FztbppTLa0WbOKZv73gj
/Pv1W059d9oVWCqrbNJL8KVVsJiAgLzZlwHe79Kn7RHoShv+WmKjxP77JMVYoGE0
heKge6vjWoYXCLnlPg2CSdvTko8RxlLhez+hxW0SyM4F2tNyK19ROLd3E8Yu6Trs
4jT/AcRNgR55mR+UKQpJSBgaQoDYct59MOoSfGY7f+WCrHlt1dL29dS+4+3SFcho
EICXVMDOEL+GJxOIqZ0zVV+ckJ9fKGZ2jRx0L4u/5POsv0WtFvXFVeqqd3du1yh0
zRX8w14juXqQNR/d2bRe4A7wpyddyIR9QqUYPaxhadgBl6nHpiwebp5ocYCG2eKn
N6U6iMqCNgGSVgGWrtgxX/bSKy+XPX/e07gypiHDpKfB+rdVuJWEnmPgot+hUMFT
WNePx+hT2xG4UlSProuN39EIdqtrgd5rhAKyo/Zolqaf47kyR10YSe9gTH4Wjaod
TsJEkdUZY6R+pFqC9K6KopqUc3U2DRLIzKEvV0ueqEOft+t+98b/R1uyjaWksXIE
bqcJ6VZ8EJ1+iA/XGiZ2D8gP8UPY+3S/EGOFK++CZ0Y1fj1ZAqDhlmnTFj42AMTZ
rLEUjMIo+FYKGyGVXpVCjM8H2uldzJxZEidknuKjxFeANfk9es48MMu3URX26Otk
qABXBrLCVwk043AJgAjhgvTUAvlTKU59nYgNAu8L9GqQO6jIO5NXFEmfX9LhMcgA
6YDUeiqi0/FhYTbjhqeoPtuoTFpWq9J1SLTBh3d9E3GVoHAZiMd12e9CqrWGYTwZ
Ot/XZWq4jZANNDdJkjMZNlSjcliUWxQ0yol2Cyi5ubeuxJBy7i92W8mESLtePHLQ
1ZiBWPQAvsFP9E80/OxrD2sOowG2pqgVdnif0AM3XEyr+gkgTgg2hjmdX4exIcm1
PPihxsHh8UYcXL1dGBH8rXvwCS3b+FiMyn+uuosqueS8mgLd31roRtP82YUhlQmE
bTZIUlB3RYDWm53hm1PTleAwclGrTCrEY87mX7KHkAZ8fg3R7vmnyfXwMJg6tIYE
g1Q3/OgwI4Mx9H5S6VxzW0m9TfwMWlXZIYOb3fs/A4JEIHqB2DIFBRh5hO5wWauj
6EtdpX2QOLyLl/K44/7AQhzCnBJuTpskYhhVA6o6ZG2Kd3MHVbh3erqSX+1NcqU8
xxOolTtZqv1obqIPfU+LYlKGRASA/2irbpOZcHGxIAsT0rvBDpXXY7S4ZuGkhubt
8WW4MM3TGr04F2alR0RNYfMarLwvSYFr6iMNfBkaeGRabZ9pvzXXvfs+A/lElixj
BpK3AHYU0UrzLnBHE23ppzdzaPT19BIc5mY2MH9vpDzW/r5ODY2cl6IycMf6PBPM
es010VAX8ONCRQESnOhJL+dsEdV9JhqPHfOuVYXLyw0JwMpWwoX1oZbFH1DmhX/B
qiAS5HLpsUifPApFQJ48tO055OQ5XomWAqJm/nPM2a6xYJTOzOxUma2W/tMZT0Gu
3HkaBHFnORsIREKCggEMFAdbzQZhPHiKh8uweVKBDjVinXtrKxxWrKilxetlBchP
gqluZ3ZkyuuX9mDHsQlGlinRXhuTuErzNqFoEW+RqkuYVehhq9BECKXo72AJxn3a
lb/SkVysyRuDuHpA6UNIAJmkgwrg5GNAGyI48NBpNFx635aUfva99G8w2/7ZCSuO
2NP+/UcvjGhW9I1LwG/fi9eVTOVvJqual0o71cI8UX98BThnG3nIhdkxQ0FteZY/
yiTYtwr2Ab3JXBH6bDJOp4XWXHOpL8Qobs1iZpxD9lXmkRLh+vmVXY7rYdvTvMMz
IoBOP8/jNeADs6U3yUHbetPuWo6vByV0CRSkFuNiz4JaQpKCpO+uYeWAXmgFp9yQ
aA9Ijd1zdEaVRDOJDOZAjAmyqDx0E4SM4hN1AvOvppt25D/Wlly9ZhTwRFyYAGiE
kV64HRgTArxpkUWHnK8WgM9gfUJgFx6j5TV+xR1mxGQKzs9LqvSnQNVwm2FdODNv
zqWt/+OUhFFrR3yHp7IlYZuFXrw+6FNb/m7WpFdEFiPf6LqaZ7zpYerHCIt9E6t2
CjM83PEa62NB/Z4+HlLM8oxRoKqWAPH7oYg2PYlR7HbEhUPBsNPtv8PS3WOmA4fr
dCcLGUDL4tSBLJuwuBLJ7MBDNvtyDQjR8Jt4yyXtvMUrh38wKGuZe7u7ca+8T1LL
qovddG95ZUh41HC98Wf7zgrfWNgtHuMRsjrKeEiSq8dYoTgSbzEskxA/6pxQmIea
xuN80kUyOy2c7pWcohiVSfoQaafT2I6OdCqM5VpVsGmpiXfJF5PfEPRRDi0C1TBN
st3UC1u6449c+Kt5A/hwrd7pBse4jNsCqYO5PVdq9+ZwP6sv0e8U9M0V53YiqJ/e
K2PKzsyJ9bepVia00UDvDyYXoF4GmHeoKg26rqq/UJ7LIt7T67lKYXqFogIoKcpu
Fbpy3RGaWxVIQ6Em3v3J8PjT30N0huFmOD2Oj7vntN3DmPeENoWDzEQQUgXubWiP
myM23L8VS87ni+AXJ8iZblBBwGUeux5wY3Imj/sKi/iOnPMS0Oj7CbQJJfIr3SL7
QGqgXZy6/LTGWncNq0eN0GwjVsDPS1XbOzAVqIoaZQUZk+N/3Z8mCZwOODICF4VI
+QAv1/onzjAizAdrlJVcK2lUwYYGD5Roj4K4w/msWWRct3UWyMFH5X6rbHa31XpA
5BoNcDPnE43NcwNwdq7qNVlcAtuHUAKVruvwZ2YleeTKa/Ub23R/vmnTWgxkYVlW
gdB6gxKL8+33FaQeG2hC6I4cvky8rlow3o8EVsdI3kTGOnJALuF9n7h2wVEAPS4v
gTyNvLm0UkhPx04GwIOhGiUOSG0vagtRe+z4tFqrFRboIGER8Sq7t6B/ugjWArcd
aj7/BCCmfd+LwyH7LYz/nRjwFtHmaxgwjVPQOjgkszA2pRcACQP6AfXxv/mJ/+Eb
cIekPWOGnOPMIb4I0F0ZxhNu8pk6itMR3a0ac0c7yM712e3Bkt5SG2dFizqwles4
ykn6VC9GTGZN6580mudEjLMAuuR1CrkldrLaZ1CTN4mG/UfcHD2g77QOgGLXQPEF
PSygfc7w46i8O1Bbu/r9l/UNRBuSF0oX3LEWywpJ0GE8VR4j6uesFFyBoVMENr+0
DRoWl3l9A35I9nTqwA22yAwNKkjd3G+PZ1MFROe9IE545gfJcQjRCChnLmy25jXj
lATje5lkuhRHB2f3E6qtpebrFK6cu5FyTfRQ2MYxcUupQx6TjMoE5Y5Iwp94JaiA
pFEqOrsyKSn0UdirLgerlxTH9mzGDWr+qVuBYkJsneezIp7ZJDbkamUFeW11gURH
uWny8Bnexx6ttslGOPP3t+RnsPJs1ll1OnuomAlIfCMMxKgFBRH73+DafsZYSkfx
7h6/LzAPwv/8G8UTZddWHiBTi4aaCW7YQU0iKUzVDb9TmNgUwSspScmCDIFhHbzr
Yz3lJkQFU6YE397rLYBST2ChOf76Ba7Qnxa0fnBJP7AgAZYQaACzEVuekNnft5NW
Ds08BGEmw6GIEgP97Eh/mmhCIi1mOToNMg73OgNKEenxFf58KspK6+PPhlyvKoy9
n0HIIQ5KBZaehUdS57G/mipvViqsmD50VIDVJax34k5TNKwEZbUZoEU0lB2D4HKs
SkyXqmPP8k82hpCo5S6YH281Sdru8pjNIEDViszOkdrjtL54QiaeAThL3olntgPt
OOyLGqI7ICwI2//Ie+4WsyPPIbHU5P5L9/a+ZooxvEvMQrvn9BPBs9k7agk0bfZK
t94yDZlPFynZDeHQsP9ABO76zn/82CQAnBQgFN9siKtJ/5IY7ZUrnT2wUigZfop+
rAANhb0zmXnyH9uj+ukWGU5VuOmk+lpdXfaUxLd9tKKVcrGvM+9USFZMBirMiycI
B2yM0d9dhCbF2hYTunJKb+/x0MbIRf9Z8tsvsiK4WeBr+fLe/Y58I9MWvWdTX9Vd
d2ZdanZMWbj9/ND8hzinto01scXf8Q2hWQHUgjb5MMIq1I9j09SSs2Ex7CNUQpTf
IpYKP55TwNY0Brcehm9T/bnb8uo5eroUqCOOp9AMNulXgXlzVcvy27fSzgmR2496
xEn/qxlioOoAK2n9zSk8wuYAqoW/7QLc3gU1Li+jB49s4RM2Jfw5eLyFv5JXNXoE
G6G6uiu4iYL1iGken06erkqx9oy3ujz4rb0kqwYAYCHmR+6M0PGwyklGMi8AP/21
Sw3SEtueY4ZQpCmT3GoWWP4ObAn0onl0b3Qa4OmjdS361nwI/I/zRFEnoZCs5ijT
Qt0Wa3L7qejoyXvkoEdb5cS6HP8FM2mrjNKjjDbBL4P1PhKAkt0VDvlLybP2eLSU
465Q47vtPFIZVJZTKZlSerlZZ4f94zRaAjIWsEVWzGgW+1xDStTmEDA7skeZ+27L
KoBaHq9sQ++zEUCFdxjQ+4cg3iulll6xQlQV1ow0Gu2zHTIG692QSyQjvK67k7pC
Pq/LtihD1yIQGCZmExMlaAtRJQWizVCP+jXeinZJPPuxTsTbpJcpELDR/hA+P78l
7zQGdIV4nVgbpW21GCvilCqEM5s9ZNeEFQW2x8+VDF8yFqmNj/9ZutpiBemISJKB
Qx/i+fL3LRzQLIl5zIIxdNZRJBBuWA2RDA+XBE2TRo85nxLNxRZpAdkjcUwb+vjQ
sQuKty/9bdWRrS/Yg0dsi4FrFDhOsdWxGFwkleuSoEiWkw8kinWPFyAu2nsGwnu+
0PF2pZ2yF3ImVRMRRNaaj/5mGOlGkyytAWUP6XGGMfzr+1YDgSGQGwfMdzT5BtQf
Tg53h0+RrgcaBQ3qY/oxzuVIxtR+za5QJFvocVp3T8YqpPb9damIoe5tG1nDLZ11
NfKmNyQHj4yws5Nx52AZ6QcOocBv8C6z8oZimMoMLu1gIjz29tR60gI/cOzMMvIP
2HefsNI53VzZgqiCokK5Ik95nlgGL51X/PyBFQeYbuclFFsLEjKaFi/vjixi+aQb
qqltkA0bdAK6Ntc8ZQ0LS04X5cqOifjViRhd3+qWKg4hxzy1ViJK6K/q67DRySCv
5OkE/cpGH3OAwCdaOlYCNNzuXjmG4jiKwyWAXH1Ws1HV5qRU8yOuL0AZtnL2iC50
mr4eJZ3bauw26M8NIRsZIu7a+5HbghYrYobB4OKHfJwgZxphoKSLYiWwr/yRpdCN
ccskT1xP6n9lQAwo1Z82lCXz2HsfleOWOaY8RTds/mVGO9NIh3UDxoGjStIz+1BH
Ic5H8H+HxqhfHxD2GtFd0m3O5cbMxcxKDWAYxRxUwdA4folFltUtR+9F2LcpzRH/
pA7CXBkTp8ZkxfV9G1dhNcAW9cXiJyVDyL16WttUXzX1PI3kJomdYFtMq2mNqIxx
rX9sOSB1qJPxwZaQzQ5Rjk7hjtQCOQbcBf2Pz/f1sLPNQdEEDfZ/2Ytoi6QbJTde
v5615LRmfyfTjrlIZXQM4FzS+yGZx+BxRMZnnjjfXEEvE0247hj6zThH5Iy21uCw
mllbhy1NQlaa/1Q2yYUv5JRTxEk9TuHlM8i2N77c+8diYUiQ/D4B3Kd3eGtaY1tB
feD56DOuh34VMh5HFJbwNazLLgR6HPgd8VHkYkIB4SHVafNWT4jq259swOQqlnRd
MEu4BYXWI0lgTaET956vAWXOcVHiX3v1Nphs2a6d178kWdS4A32YpjRBQtBAqmcS
RPQC5/ad0cQEByyKnE0ITKd290XrlTKcKpu4n8qcff2ZAiZIcIuAz8GpzTnAUqiD
VyXV+oJMfV0VUc102HcV1Bdduip4+CuCPZ0Lc5BbsJOJaH+n4djASE6mvg4j5rzp
K3kPjoiwsXM6l3vgBNLWiwmYPQk6dJtl1d0wyzlYXpyVaMDSIaEUkBIyPqW7hLE+
45n4bI8OSGcQmnBB2jD60topwSpqY4e7dLbbBPrF5w3oNs/b9wwFtza+rLnbih2f
PCSejizxjPp42nsP8J3UrXUVknpyhrZaZ+quNyEfnVgHSMSiVgbo3ZP+Ev4v8CWL
6QBuSr1P9ZJuxCFFVlMWhrumnU/qnv2n/KgVdXMkqeBABTDFKj3QY6AD3K1Eg8QI
Be/O4J1xDdlrt/uYs0RB3RbJi0KVwljcJ6hfNMOy1/0pT9CZo2UEJuf1kqY0hBo4
H9PTrfAC9SPfENv8w3kOR48OZiI3+pHIg60bX7OS7L5V2uRrOyMi6m+cXR56gnpv
8ea+LKoVIjtu3oUjG7vPcazvqVcpBp0tLxqyAbzzJcRwKQRXSo6QufBYNoC52dRJ
q7kHs8A0VJ54lsM45tIV0wf/V7XkxAt555L5TUdoSe0uQ9EKYaVKFjppD+E/+uWH
EIMSHHokJDPzxmYhBUUvM1ua1W2WR0DndXQ+uLuVBWijLXUIHdf3xZ2ZuQ/lKZjJ
wo4V0qATGUrn5Cz0k4ZV3MBi4kJhPhZLfLX+jAajIrBVekFRUuUYpKRX1nHnkPhD
KQbrHN+eeJFaEmLOweQtosjVnk0m5yThHx+mdwVwh16nWcgN941jz6Fa3Jwxdi8k
4yr1QzaiBGdF42CKKJNA881T04NgTW+W787goVc92sPAVZ/G1zOAxhJm2KRWziRu
/3hkI5/EFGoSqfxbjNipev1NFwZJZMCAWiVnyoESDRusNY2o8rAwXdA03pKXu/0X
zFt2eMtISr80hs6plLEbWJ8xWysGQHbVuGYgaC7OBGs8IXtQAfkP+M/JWBmnMcyX
UUv5GbYwciUQ/sTjQDYV1DJRNyE9jvV0tSteDZDp6HaFFEYc7040ueobHQ6atLLI
7jOgY7VpFdDjYluUOnfHpWdsbJY35CDInZWHbJ1wuGyNMMOHioOtetA93wOrAB+3
ZY2M2N2tpA8JM+aD2jUsDflVDlSw3jF0kbZ8jqxbJN4ebes5a4Iwl5aOK92+zl7E
m/1eVd+rlIJPn1k4cppRZfB/YQb0fBod6kbjH1PHte4KQ5jv/YR42ZS7+jKVT3Bl
AQCuvkdVjMo4hc/ZKqzwNPK8lpOQGiGFRoMRDPRQ46ji98CjP4aCrfbS1fsdHbi9
JkPmtok+Bx+iUXkGyVIk99BZd692mM7j6N5reN2HWEbiQ2AS97n/YL2PJFZVf6Cq
aI1UvfcWVYqHx7S7l22yZBmpmxmpV9do5i4v/ojM5R6KxgqPXJOQKq6NLdGxPtUi
D8FXfWk7/itQvABx335YjLrx/XjSZtZD9HGPxSLwDKhVzkf/8RgWGn5TVkfwb+2p
Qs7mjWTaKXQBno5ih3ekRoBWME65wv6xzENGsI3akztECajNNstYru2ZoTjLz56B
PWzzClqbQiS5zNV4hwwC5HnMjqeXrhqmXUyuybmXnzMlzvMOFJNCOXeoMFlmwvwQ
YHlybyWuMt+9uCwH6cxSp8CxoFR4i9X/IvoHeVAxCMmgPraqouNAlLcNjH4AeyAy
KoK1xt1O3EqUXdQVRyroWKCER0IaMr6YiebX4vJl862vGT/d2SMsL5w7Widk72Rl
iIXTI/hndjvrSkSaJyZdBcC1Vfb4m02DIVIecbUdEk0BpZZOWMoh/0T3oogZlHol
5xPLRDAZr/I9mm1Wyt98xDpKhHPMwC/6/P1pR4mm3doPnfwCkaqfHp1W8qPPHJWo
x8xUoA/0VOjzkQ4cfiU/EyKZn0k6HYMVmRiTA/Au5Hy/K58qonYP6sm1MEo5Ak2V
PEwg9UQSRNCnffu+EtUJZn/1xj1oyWdWR3FggdBMpHACuRiE4wTpbZkVKlqyJFCu
6q6bTOdzF81KD43pPxsjFDKNb4jq4pwo8/5cEcPx16MhNL+mmXr/UywrQqiglEal
q/BvQmtUrdxTXPgt3wtN1GVXysyCpsC14h+PV/JUbmohlXD1AK1Wmt/RUNU+efr3
BnjwXxIVAEDYhnQAfMDtR2039rdxKjg7tq4GTXQ63pR/bbsy7xg9OVGGg/zkPcRw
HITEPVr8rpZwxKB1GETTwi8OvETLT+/4VQczgSGv8Jp3wWPe1rwQADqRl9l7VY1+
FfYFcF/Ojg+N4nN3daVnfC5LLee3ESw7xA5Ba14lZFnMPPETuu82Y6xK++MDkPQU
acmhXW/BUQmNZyw79uux8i/4XYR24o4t59PAFfVX2YWp7kmg63T6YmyR2rpo0MnG
evQazUoUV9ryfukZp5uusOkqT3CydmdPid9MF8Xp275xnCzfT0Tm1bVu2SdCxY6j
0jILIYhgJ8wcMkFhCPiia9r9ujOTx8T7lG6C9PJUTOZNVWZwMU/4NdWc4fqJBq2x
TeXF56LXi0bYQmOS8fWEbFQfXotFRXGJu5u7mcARloSjQyFRAkXgNP5t2bF//tz6
KU3f/eTL/YZGddEvHLB0HSljyTZO1pgQ2VPDIjYi1YMWf+luCHfkk9rTPBGjUfZM
A5fmx/bQt5N9M+mi5Uj31ABk5MrJEarrfHyvoBViY3+6zH0BXcZ92Kp2gENU2SxM
C62E2YKWj8YnzfnudSvxf9AY2aD+SQnRw17lUX0utJUzQijWhVopXL/JSKTLHg2z
CTFWhhoEUtxjTHRIGzje32yI8gUO/4RJWOQxi0pnh6R50M1m15U2LJx3CNTZfKQP
umP6mvyGBdVkl1C0KoWVAbJqXvwuLuyVgFL89KY1UlF1c3nuR4HzrEHQkHEnJQ+b
jzgGifEEkTnuyQWv+kxnEHgODc1PRf+wGkk4f8zwE7ip1Mwmhg38PfZeXGhZuZh5
x8g335devgB8b1ONF+966KbAZVKINHeMphgks+2yodnbS0WQ7vSRUL0JdoL8bb/r
LaXRCPs08FtE8zNufOXqI5pdF3DGxmzk1L6mKnlxj0T/3vVF17XGiJHDUxkMr72b
5ADcbCotcGGJgXjGDVIvaUFX4OI6Sy7AekMV08SQIh+xp8RzTjpvfzGFTC0/bXxw
f+RoLDj6vkuSrh88R0UbCSlWZ1n4LN8GmCU6sQMTTx306NZa3peBdN7qdhYex+JA
xjSXBm+s/gDv8guXZASGFH2nJCopi00SXwuaPz8+eqvePim/vBogwR8KL51WzFMT
gJq0QKcNfxelAog6zT6lO9eIBvV/F5Qb1+sn11iHO+ae8/hbd0goOwW4N0F4Scwr
rYnX/DDt1FqgI/pSOTy7nbLlHlpr7F7E4RWJrKUdzK4jl0l4A7IQKIo89Wff6OVM
3YbIk4THYAumKhmhMLxxdumW8KVoxassvpYpQ1MjcHfPPXwi0+Q9pGZKhUNK5k0y
ubNZWzAOtkgs0bEqlJrbTRCxpanQDWPDAVZBTLAiFc2GlQpQzu6DvgC34P0OAZVB
Q4EGw5YD6kocVtiYE6zPrRjfZIdVyn+wnRRexcB/t4maQ0Mr5LRo1YVanaCqq+Hm
gBJJ9cJ/XMENLNf75z97TrSLnCbCxi9cXPV0QXKTbm0hUP6ySMr3LazPKBKa4Z4w
nIWcwMk70DmIpSlMnnvaEis9hpeFxmw81MkHFBDQcFkoVDkK9qakxU2XWoFicNCh
0Wbf10L0bKSz0G9WyNJhFa/OUaxhSINKetJEM3OnAQPGjN+vEAxbJJScTf/u4ffv
KhBXAE1ytsrA456AkWJl6zou++WZ1YShyaOw93pSjX0DLGRzy+bjr9bkjS5KhMJ3
98OeNRz0y1NRJflkXYZn8tdDAkEIX3JqbgxIB1NvLzvCrAHtWNnjPw+TvqbvsM9E
14ebw8HWmuH18w5oAlx9xrz27SQLUjQQOJxUpFssZNPmu0VeqlIY/QN0c89kVmsH
Vn+7sM6f/sAPy9jtCaf7LcdEVISUx8l8LZxsyMlCthgNla/QOrPj60qSSDYvJiHf
h07V75lNj6A8e/96svJuBRdH6qUmZVsQEH+vUeiG0+YCocrDdQUPSQaWr+99OYCm
f1nacX259/gxFAUzSjekrUuX7ogdyrUahvpSQF/jelh0JEFwqQ+DJDfzr2+yPWGt
L1mUdalvHALXDKnbA5KaZRr4khYplGJD9w1NkbQEow4goF7XCmn5Uqe3c3sePK9g
zZINNezDdNl4xaETN8lmvBA3d0vikBtCQZ3+F/1DtplsMl9QrOgnmLqeBQ59YNYv
E5zne9mODvp9wKjTbQxQcrMd7Xxy+GbrXkUnk85/L9hGhw4wSjfu+7zeBYNOWxa8
WR8J+NZMQebHKrgi5/l9efqMXKbKFCHmvVkOIl+GAyFN8GDyLti1Tvm4PIn6076U
3kft1/BPHwFz/IeCNKQqSKJPoftahlnj1UU5xjPtiXstxV3c2SWio3R/ZVe3zHF0
1/uXVBf3aYq7PmYsEZdLcKDXosao0ZculkEFGJS1WyGXn8mF6thKE4TzBtODN7SP
FqSMKHQv51S1z+ARqtEKqSecJoD1riJzoMuhi7w7iLJaDZmow3I68QaKYVk9YMn+
psSVPQcbAwc8c5tCSS2TQS2JnKmipVopl7MP2Ou9ImEl+IxUKnYGMifo7mVe2fBO
NeWW7Z3wAQNnVzyu1gSz94x2fbqGJtqiW8sTjF/JVXuQbQQHwMvvQKfkg4kCNH45
X69Du+HNAFOqoV0p4Q2sC3Oi55Ji+W5/PN/Bf1S6KsbTsehZVC4iiYfePpQ/pztY
YHMdQkVmYXNHaYme6T/SDH2RASO4L3weTFRScPXik+buvJhozj6AVniZm1hkw2JE
SRLQG20vYiDn4DbYOAIvIZF78fA2w35ui0h2w7R/gycQS4Wt42JSFDhpkNuULs2+
4cuqBZe7W5T4XSof4lHEchbB4tX8Qh927IUGD9YVztdAGBZzfuFOzGZbUHH9/qsg
U3i+RzCeIIyjaCVfhIEu9lCR3K/JYdTzL9TI/D3Fw4IBnx5an2tiuWPsb10sE0p7
wx96QkH4+2k+YU+5yo39lpTLuyDHSJKWHT1zl9IZc0nP83HG9TPdi2zRtqwoEThk
9hIRt9vEghXsWv5k+09xYLC9IkkxwvcTrscLFzYeYLfmbhrfxpTwtJgIPXv8dt/Y
S3u992tZrrlzwmh+WRXBpOYKsNZgxARTCdIweyxpSBxA7LYzG/B9i+ul+SIxpoXe
J6jo/Gd1XxFka+oufZKNxi5G1UnvsZPyJz4e6LY7NA/14w4CZI9cIZfG1WJsDklp
pvmRzVXOInBFDTh9R1ZrVou63aeFXDR/JO7jucblXKYtMA3rI9n0yjmOmWJRTDfR
PbwFmWgYponk5DvL9OdDsaCyZn78qmYnDt7lcQoPFNDimO3aK5uIIlu3rH4RnLeJ
SHBFUlt9CQ6CLHDZNVJzu67nngJPzx1L6nz1uPZYodhg7XsrXeLcJbagpDnxH9qK
eMgzLhMwjJ033dU/Y7mvEp9OiTTs90zeo5BhErGP81fliklCLwkY+7Fpi+mHMlvQ
MhFquAJjBYCU3OOVLqJxkNHZHnRrUl/I4r6C+km2YvPsyCqiupf4q0fdTvJ/ZMnL
PelPS18EOUtCH/1TKFa0gy94jUcVykPa4obMxRA05g7Q4bMDdJBqeW3mb7E3IIDH
c4P8rCqR2bGyDQelTNr8C8F52qyw0KOb3UQbJgHwnMw+IKI8kKqes+X04vRQcz09
3x4NT+Sk9qhwXG4q57SjJWKvli3H7sJSSloBYSOGNdSjvKOvzajZ8vkaKlmMyQkH
HQmcPpDvmNfU7Vx1zp9JHvU3wj4U0D9muE7LUrAOmLhu11PLBKYCPCj6isCshX10
KuEf1UzbNO4+GLrLLUl5W+PM4O2kuN2xtRQcENcmpzLAtdiCziIEKKLvNKxBjhLX
aRCSSmcJHRVPIPF308jWkPsv+5Dzj08fFRtTkYanXRmqvZcViLUpQEZ6g+ywXWF0
FBQiy1FpU9nhGwbzPjBtPuSTVA4k4zGX2avZBJ/p/FkzRLkqRTNCq8oDO74HY+PP
3leNQ60abHiagpXnS9tz5rqJkfp1rEUzgStek5EN1B+9dQHlxddDvWkmH0VTrvJU
RKfREOUitv9M61K/cKtu7dUUJzH1ODMgZOuHP9KCcd30qY893AUheXcur27rn1M2
7ICRvtUScBQ10lSYS8kTpoALNhd4FOkLGZek3+AfgLdVAFSoS3MxwEtK46VZcMPn
Mr/OU0Wcc2Qjx0ORePwwc6L75gEjgOrwKJ3yZzsXTrMkea6WOF3W9Yz9gVw2TqJQ
Lj8LMMQgcWwkm8xuIhOTUmFcMIj56xcsjl03pahSAyqZaIFyMudgUEliUCWh4Hyc
lylpyD5f71EcaPTbuBk1+eqqRLlwcq0cs1bsQTbaJebIclQUEhS93nZjyjSOvTjv
EENDGiRGpQoVv3TYX/DVocHmX+8qTd20YB1szx+M/XIDlOzeXf5Zcq+cNh1bT9AD
BEFqLqMgpybgNnAknjeoi/jJ9v1HHWoe8+85LXLbiAUQCJPwJTulPZBgjDwoxhQ9
JT1ek8ofzHHm2M/HbTvmfsJQvYVi2L7ZLVBb0fdGXfCfIbaLXqxd9NVZ+Vc8cj4z
cI8DLOVmfN1z7c4TaLfZ5oTTqYF63WBBznCBcMSO/RrzJn/wePVxnkNooSTk0cXO
61Z5q2LM+K+cj4GlFYNsG58/+Rx2JFHp0oS1zdnzPoKHjqxfFs0RtPZjBgCBcp7Z
zWCyA0NxxrGzJo9BW7Xj41hIdFx6qvexFdOdhLGe9X85ETmHENf63nGsq8L7L/9X
ZzCI5oBtZpYogu5M4VcETZ1EX2GQeFA8XqnxAyFlLGPzZzV6oxFJYJEiH8GqNZYn
lmWnEgBy2n9XrP2Fl12IQWdUYbmVcacWYIu4a7ZDtZnB5Y3e9cn0nNKsnLBqWJxW
f65mxMJ6KvlgqiB8vz0t4/l0SbrNP/+k1++3l1daqwsJII22THTE7subAqMgl6km
n/DApF8cF1IUd/Gl4LGA9c4XWLE7zH8GrTqsTv79MCCDrQCOWyjiH2uO+6KM4EvD
Ut++uI+FdWNlWB8xlOPffZq0KiHW7PvjHaO87rrT5mHHRYolobJxm6VRNVUiqntY
RMFDB6xwl8/7Hn7ZehsSBl73ug7oItOTXO+hYmPM3yUnR/IqnLJwyly2phwuzs5R
02usB3C5HNjU1fUpYb8yBJwluaF5RHV5f8Pw7ZIgzpZNjYLKmRvQzVPcou5Ouecu
dXpsjlk3pDBeMSGfddky+UV65c8V373wGNpx8T9GOP5OWtP4XgcEf/dvWbMxkvdd
2nkOQ3lI0vLI8XO7m5zusjqTulkio3thJPinaatQvaXHVpRXYfqpdOit7YnusXRd
C4C/HV2KIpi5ZtnXqe0fKB4jVOJSdTUNs6ogi5+otol9wZQOxyKO3E4Lg0puuQSN
P5vFidN7jZ9Z0AZUQQDAel44FklggxuMfpQAC0V8wFlLEqNoTSUDv+b/9bXMbhkr
dq6hfzdY6WBO65WNjO80wlFfjRglhZik3iJZllFmL02Cqq1ESdM+BeOLf6U7FvZx
YHae4HWADnhV41kiUwYPqDamP+kb7h0qi6l2iYfWpO3kIWVGSzsG9Y8PR7KZbRzX
fpcI2KFoF7dlhXEQz3CkVgHjKdi68xEQtow6RpMfl356tEYL+ZLht6QRfTgh5ao2
BZQ7vDV8yCDwiMl35GzTGYSwHvITy4DbYLPqT9UaEOe3lveSJ31SHyU96LYU1tU5
PezNX6Vcb7hU3ga4CtbuUhpBHZJP70JGaIWy3ZPb34Bglr3gG/4j3AJd5uqlJlJc
olxErt7Vvg8E/0KeKWm0uy24gT+reDYeltghFm21krfH3yRHRYIP7SPs4eIrUZEd
EKLJdfiKr1ymySA2Z0WxBHFKKyWWqVHlGG2Op05bVlwfvNQi/klvL5oAjRag1AhP
3SHnIv+s4q1NdTWqK9W+y8JPqsq/iIfzsZGgXFR59DoRDEZ5AlOVYyYRBMAnTrAv
wj9wftF2BrIxLUINKfl4/yodET9e5d/7UBidUI7B/yD0zO5hW+EnOoHvDOHumpYJ
svRi3KGCr9NKasutWfjuitCpkoJO1ZEpdIjeyuZ50Dekyx8MopjQv78CAnObcgEB
D1WLmpqM0YnLsTinrXWfqG0l6/Wjjcv2bnnlLmMCaj0l6a2J/AGOUCm905PwbWCd
5XNLb27rHndsWTQEf0TPEH8X42B7JRbDa5NW/2AptdwWkP1HQZ43Yfet8U6+7iPS
JQigjsux8OVBawvgb+S82qUeGvidH3gYrRG1SPCgl+v8DxKBSxIDBMe4tSF2A2Kt
cq9bVWv1CEc21juSMQVcbs4O0zuPX9Cb5GWsTnHhDUaE0dOgqqBh5cgJ+fFr7IGp
FyL268KgEk7PU8qnP/xGbbnXvvnXwVUXPZIWF0s07eMM1QbTXHK8ZFYaEM18g5lm
H1JdE/R2rhVyods+S+fl8OUvSQFwcgWK1czpVoI9snbhycJW2KwoaqxqZzmbFaY8
Mq1WJ5G3qqJKoXRoVosV0yjt61PN8cb+994//yZ7TQvi6tVqYcGwh1nbCLAKju77
3gM5y1y5Cxh6JB0EDzcyU+lKAhijpRa8Q2yb1kU+ZCFh7F9kfoMsU1zOnbIL6ECU
sTdrvWNrVdpsqoF3idSo5gyEFGj+vWomYzRCuvPxs64tJbsxLzfcZ5pTcGo1IwEw
elCOwUt0fueTIPvOa/hXxbnz6mAQsaXHRMEPxO76YB+b+KPxDxd0OYbNGpvCkRI5
Br9TE1coEJ0hmeKj71xAmKmdoAfSwNGXM8Bn5rxSRFfv+jIqSpfmRnd4MWi8FiNz
o0B2umUGnMiLPCoH16j0Y+fFcq0541wFqOr7Ty+f/qg1Oyk3twfKc1xQQj0i9cKA
PBYjJT1gjVQfht/Cqd+JGjSll7ZtDkDHhPkAsthRMBwRmwLQCgZJ+0RrU2vyqPXo
sE+ZxosJcoq0rPurU5vCGIZMZlr2e3as3tE3aiRnP1YI2I2QgaDvTBQ2XnZbjrnX
wWQ2G0VOqx6nRg+a+2sKNncyUSAChNl4vuLdUmg3V2JU7RkPNe2qFNnPFmCZ98Kq
81d6WqnNZZG3uiVScljqJ2w7eXethSAmhYkFPiIcPmBVakN0FbOd9RKjQKsRwWIm
fFqLRB9S309iZMfloz++W6u2w6IGBW8qKIiVW6bZONeqgM4wuynm8jkGFj9hkBDX
`protect end_protected