`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 45040 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
DyUmSSJKy9uR92lovAin2vfMotMx20JpQzz2nkBLjlWyhIrVwxjoBveMgjkBmaAl
nVNdJb8FyvOopSioh7z9iaj2K1V8jPaMOZWDLAaE+ql+89bn4ictg/3nu9F4cCdy
hkTMiJz2PgwAO+wmfxZx3PzotswpMwYz0FbzRyHwbgLrpnH8oq2oQNzbCyMo4ka3
23vvLPfdTw/2k16vKlIHwkSN+YJ5PbIUhSLoEAeoEiuilt0hUlVZD+LtV9mFJCRg
4qJBUeHfzWKK4JRabuEtp4VuSTnKorz3TR3kqrL8zBKnIFEel/m5fci9oQYAkXxB
nuAcc3yZHcOs9zWJLg69e0zi48B/AAHPDtLFDEDsKo+hpWhsscc7faFb1yF5ZKlY
5+QW0HOw8ksv3m8h/gUni8mj6IuFNegmnHf5/GhH4R5/PXeb0SwMnV+6Ub3/HTs6
Ed+BySXDEq9mhVHt3bt2+E/Dwp08LOyXY56M8qZaidjInIe2ZkJRjzsYmNzysRYp
LrHJycFA2IOpvIIl1wFnTlTAGpWvYQfekO7eGA1blJQE4lfZUmusM6X094QMd0q0
weNwtJDvjM0VBYNJkNYbNdZ8Pps/q37UNI/mWwEgaqwTvUEDDYyj/LToTtgTfjFc
Zgf35u7EUE1TGRVkj9oT8G+acuHWNbzi/8cwjcFFbdyuEXBfpjkFCUBL+yaHD3Qb
SfOz05rcLMNqKzj/Xyd8XRbRo5hZFrEzZ+SYRwoBZGImGifM3rgWdhF8TPaAFLZd
8PcQc8XaWD+rOXM+p/j0EXFvf0tMDoKmLU/8YiHJ+CcgBxEsmuEoKNokGGhQ/qmM
9jfqVzZ8aPktZKxf+ftyGx+KyxQUc8sP+X4yZESgVr6aOPa8ZRL93Yyn3EMB0t7F
OJfOI1VvFEqyzO7N6+eymA6jGDoQV3cHr6aWrg1CghIlsxr/Sp6wuvPi4E7+zuFq
AqlD/IdIwxR8+tmaPIEqFBL2WojGQRKW2gSRNUZm+l8jAfjsao0oNMwZ5fotpEC1
25UKAhQPdIqdKLQABE47UK/PQBfKU2ohIyoywtl9yXDUO+hCxDwLk3hpFNkansuc
LNgbyfN/UExE038m/I88gbpgVI83K3kgrgPkz1I1rJ4H6yhKlIPrPfzWAkI6FNvy
JObO7SzNyC4xBJMIfYDLIz1wwMRjkuYJ4nwMVU9V2pp7PtkneNiP/LbW1+2p26qS
SVsu5J7QkXaq6+hbpDZmFPQ4GVknEhsqw63431SPtedaaa0tCNfY09fQg1cJ0b69
GLwriaR8uYHKdduHu2q3vKj9cnKeE/BenAZgAxLVhig9LTKhKtupK7te+83PVea+
LYDupWuJ2WFXrjzPb9Jgp2O7XvPigoHrmp53cOk6Gwe9on3nujGgz03syNX7RdXd
cKb9RTKzMQssnIdN1QoEPr4gZCuiFZZkFicsxkbv4hOxwFdlDfv5aGZeioaJ3N6F
JofXc2BLs9Un2C+0oi3abX/Jm0akIydaHQaoQFxHdDX5WK2apq+FgyxMVH2fBmhc
xQ2KJDmlfwzzRbDSwWqj2ZZvPafDuWg4ipZvByv96CzUvS8zjz8gLE/Zjdtc7947
k3s0gou11v8g23z0IslvxKe1kvGo4iY3u2ge7dObnMOsEi4BZoV/qiE9HW1GkUlj
avzCcE/MyCbSHbIVo8hL+Jem6Lv/BD16Do+eIzfOeQlob81VKLqZtYRL55Z3PQ98
jt04RTxabHSreyzY0GoDxY2XWnrAlYh9mp6a0IaM7o6SMyS8+oqFNn5+DS4+Ymv6
uE8hpeDi34tGJvZf8rUaPZxhI0WjIa0H0QE4Y1iuyTltURxeZ+LvozvYKb4R+RN4
Sb3w8RtG2r6owfMI0/rChMrzogZ/Tibm+iqphNS33nQsuAu9qIaFeDKyi9Vzevjl
D/WB91KJi7VuqqiS2jeVudoqPRIh6tXwPazE7SrZFXd78AxMvyXp+53zDfDQzX0R
gs0xKejetz7EmeIndTzhNhPGoTq1hEJQGiiOqHRCZCxYPwGq6c4lrdFQDlTrae+h
1tA7EeOxcpbpCALXE1JAJ1L7M7xmBV5uycfo11XZh7nEIoqlruU7CsPM3sPilzek
bGcKShfYtuv5RrK2WyivIwmikpe07HZdnNEOonncPj7SWsgZy64PcyGlE6TLe5/Y
D33YcIRbuZgxLwTxCnlvCxJ58cYFPpMPK6Ng6L9FwqRQl4o0FpUplauRII93qpxw
MUs1WoMD/QYznsoDcuXXXNcfUr6enKgIA3/ilPrpCRmWk4LQoQrsszQuuhr4XRqE
kAYQwe1LLmoPSuqhYUisamIGB/lRC+qxjCBNlC90fK7Y85PKwqDBOdoV2aQsxzJt
2Y/PXSclc2dZelrSf6V+FrQshp/ucjFUnef+jtm6376PSHxLLwcF3SQ4NJt1+zHy
6kEkj0VPlTcYmr/QVBuf14MPZlS7EvKPTFHeryrJ8L8rWOpKMPnZPzygZTXanrEO
oK3Cmax+nxNn6iIWQnFtcQYK7Ur6Ti0HbvfNlAjaNwllLyUXQI30Q9c6Kn37TUTN
TxR2hCQan/6c0pa+o63me9VA7oWQaHbirb+Sm1WmBG3g87gf5NBkElBwymBMq39w
WgkPTfui/Q7Scz14iQANO9PH8SvxTrQr93D6MwVaozgTudpoARA/jli8PZp9jV0y
Pj5tfSQOMPcQ4yYisC+t7tILELn9iIG7GVfY+NY/srtW5I2l0QufDkhL2jPgs1zb
BKWjmLujLtjomGBqMHpvALXG2R3fl51mh6IBRJc6powberIHaRYpDTVDw+EMzXZp
XNig/2Me2ndoJQ9AMQYMVXpwBhUhOQtgsRBXJ5RcpGd3K5n3XTWR4P5Ydd8lb7IG
Rxog+rZvoft4oD9n2krr/2ihZALIkhdBiMP/XaS5Os/1IO797OasH5BYeko7qo/9
o00OqQy+DyC+W5NiYEiRWusy/TBIV01atm7L3/YOGv+2QLU5I9Y98OK0sDQVUMZa
FfulgUYvtu8PDfZX8cleGeINGcpibCjw3Z4nSKCVC9pejdxDFqQFoakYEuQnsPkt
5ZZPV9ln7tweYsJGog81xlnXlPE+dY1VW6iBAUmJQyZ4YPT4YHxnBdev+Ns6H2kc
T8wI+vz/97o/b6tupaOlEcOkHQWLA0ttY83QN0M6f/wUzUbyTbaSKNnjC3Lup354
BbZbEfx6nto7zXl6oeJ0yYuE8BtAB9gvRTbGHep/qcEatN1IgACL+pYK3QzjNRZP
U7n/1MGECXONkmeX/Oyhz21wUt4mBf9baE1FIqFVN9pgtBnL5gC14F24J0ELxdDq
fnEau8reMUKUECA8dSSWFjNSR3Ii9Bed6+LrGXTBFNzbv0NoGM2PMAb1ijw2YpLA
470oIR5CHgYW33Nn6gLbkPM76QHY29/59RJ4Agihsr3PEC6Ou0j+jj50qxJhMEIY
C3djyCxOhFS9IQlvJSoMWT1sjUEY9A4U87Gz0L0KpKvEJ+9Wt4kLMawO0k9opuo1
Ed78PbIJnU3Map4ntWUrTZKQwrCWAKMS1cMLZ1j8CKB//RetxfOw9tRJ/kF8/6ta
3iRf8Xq9/kQlqQh3L77cZ4uOUDMzLNAIFFOWsxw3N6dpfxFrE0qQSBWrgxcHLQe7
rBVUnDLVP40cRQYzThqz+uUhsvTLHyBYAaUUwhmj2SBRmay3itB5pgVj0c/jKSxU
Ujw257n+EWn/LKR187+5b24HrLAeZGdEKLmR7t1hP7i4p+JWe8XYfb9EEwF7h0TO
qRhxMVKhnDE5DTiaNrG+deAcC8s9V0Ute2qT6W0nu4j6mkXdwwVTK69/cPia3tjL
ADIIfIrJF/0/bB1tOCZ9p/GXYvhwAVFMxmUqpXCks1eUybMHydnXmOMsXqA3sTIF
XGb0VBGCttrs0E3WweODzcaP7/NfNlYX0swy/x0rGAahu2GALOgffpxGu4LekYAg
U3pfOSHi5KUj4a2Bc4E2XBq5uYWc03la0u7QSWE+wLlxlIF0825Ee1/V9kI8L+GU
5P5hu+8j08tZNYqhUUsGWnNITiAQZFyfnq+2X+n+tEIxsn1MJKwr/ylaUEw8GFuv
YKtXuJCYxGZtk/ywwCh/l4SPEaKuozd1CPmj7pWm9wgS7oODrtCXGPS/lv/VOVXq
QQp3Yr7pWWa2kzbLH9IP0UNzypKADX0DM3H4butPTJyzE5QXFIpAzmJdGEqv5iyc
BqxOg2gU3246O81jmqk4qKmm+n5YQ7Zg7ILLdsx55wbfyjKKvrZlqd53OWoNZJCX
kuMwAR75M3EFul/QaoNbNG8yjmUcqV1YQJ/TbNGKi5BFT9ulJPrNz312+d9VigBl
QjwRx7xXMMI/njZFOgjlUe99qbvcRJrK0+OtxuBVM0lptlkrfcwIkfS3B1aVmdzV
XotQeJSgu7n0rfv3E0uSM3losW+7C3Ogo93rmVDCte9AGQcKXC9AonLVvC/+coJT
nB7YfucnEMwpvU+wtiPKTkmBWnfroEvN2Kohn9iX0qwHkyKpvXvsPRQM0oNws3RP
JN5EYKb8aNmCz+6kYIKbqT8Dwo74m8WehrSNb0t3Cg/EDUpPDYYBqlvzHzCDoIVP
wkcxDqNHlShdYGBtK/tXPtI8l2ZzfRHuNgGYWhRIB0vDelVMK2/C1F26f0kFSmct
Gqiq55bp3vrfL4nDN818mlUrLB9JMHaDXKaDsPHtZUGf4isR7obDivWMtUKwW/OO
clAX8pOSg0XGidakrzm2lk03i27x2vC06bs9BL4ZSF0oPlbF2rx/NowO1RVffWhH
NKT1MKGsbVFVHW0fIZpfRGCRZF8qmIsskGmOY6RTgDkKHdJG/hCaW6wxEBtKYlvE
E1R0KjIccqqnMgqXpbdxxHJi4f3BztDhslXhLFc2aWIZf9XHB+NFEvFAn2wOyEea
teS1ImYaTwMXqjlAO+kk2mjItBulgPjUCEggYdjLelnRg+uWgwdHANd0KfhI2zkS
nzeYE/VgyqzM+BolRl6yLsxgBDZV89BB7gTXZH8pKy2zdS/tFg0yatwTiKx35RQe
jSiwUa80KbG7KuNuWlIQLUKOHgCWi0cruLEBR3Msu6t/De3kAsbvJjk9JbgZFwWr
JxbHsr7DhNAlDj7K7enrOnWbDCNcZjTpaZujgthaqTVM67fwxehMjFt92BwxvKWs
evom8H+pe+7lYdBer9dO1TW48PHrVxRLsuYJweWlQFI+HrZmjBL1MaY4kK0e52V9
Gfqb0u60oOBtdAYCydqgXgwVyYUKrjOONWbWYCOmJ+K+HUPunua75HMQQTfzj+A6
kPgoQcLEZDshiABy4OuIyXIabBfeJd7r8g+H8NgENJWULH4awROIu/fNKtIxBneL
7f0CUMCg9ph1XcvtPygaMHsyKLA2n+JFYdrkNufP1T3k7RgckmEamxOuAf0ucRox
ApVEyl6GDbXr/LMs57/f5KEFXsC9QNf68HH9roM3qpJIZvyXOY+hqOSRIGhhvOQk
PVXiJH5rTahrNF8uQ5wkSK5eIfd0hGXgVJ64OdNCCBr4upEfdJzfRNFb7Zx8ov0j
Fh6uePWD3mrSr4A84F/98jkfvOqRoc1t9visZPCQv2N4OqNNSJF0rD0GPbNqLEUi
yCg7CfpZQ7/+HdR9Eh0RSkvoS0Br2XEUmRCGirarmIk1NtWBbakyjZQivTKhPCnd
Ui8/XI93BKawGzkRlo7JO9BbMIRpHqen7c2Qx7cqqJHiy/EhHNimhJ/MsQdYuPd+
1rO6mbJeju5hIOJSqTCa3y4exhVh9rOXGMmdvwpXccfEz8QIhwEd1pn57MKI65HI
ZipSt0bpKPTSaxy3XKkVlH4f6xrL2tDxV8w0aqgtiy0MYPgFVqPPl1cqYC8LIsX4
OVGsvoiMygKC0cogytwEKK5asnN2lGrp4RdomK9EtPtshU8sQ5fzZ24AfW259l+I
dhR3OL1vlYR2PrvqgKfDrebMn/kVS8kg0LzMg3jXhrzZtwUKz1NlZxpSIJsP7fjT
NJYyOFhcHNN8ZNydUC32qWj3TAs57CxhhFKNUd6EmQ06sTle3FWB0A4qzHM+PRDK
rdLTZIy/jAaNzb29YJh/XS0uER/Fs+Va9/lJAu4kqtBX97xar0nc7wsScS3CW2IK
orIyFOLh6OLfQDOyST/NHvIH7it+9pzoaZ3/zCDXVMc8Ydx/oqywEuYQIv+12VNP
IBV/IDAHJCXEu6d8Uzfts1SPh40dNWg/2hY7kZ19CBsjB8mKlmLwC442+pRshirh
EYhmNd6841hYxzwsbNYCd21hoqrZDJWgIbp+eFGzti8rgKaGK7FmGTL02vq/M9V4
if9PO2k73U5FmoABXv0dfAROSXyxFngkVUaqt1Mrg/W/tQ4XXoGZ5Y94jzhVepBt
2+z0fUpYLXWc04lVVM9XXW87r9Q5cQHohjO6o0NuWw9RuUAVjZg2eeLvtefTxpcd
jsM2/LJSIN+SWfN6V9qqIANpMDSywPCAewawb2Rnfnf2w2s4ClKcj1tFMY3wLm2E
N8N8UYZUvyh8Z74aKwXs6vF1UPNNeDBGFlA4R7tsKEtHKc5cptt2I1+kyffsQx7F
eMArwIPZFAYsZDc3gA7RZSohp/L8IYsj1kPcTb3oQqfNmw3h+EPmK3L1laQYCjyh
YAutGtRJf2v1B42T1ZEteOkmQ2FSjIosNzUwwuadW+gmQFjMAHfa0PhgedDwjTWL
nak3tJpJ5H1Xx7UuKDKii0d97SWxDQEymjkk2H+MZh3OyTwSPLfaxQS9VU7GeTht
Y3zHa7t6YATUI5y2nBXfo2bT9Bp2LBX9fpxsPqqUiJza4+PUVm7le8dkQGlld1Fv
1W+r1VD+EP0QuSUcypJVcBerq89Xhqm6HDWY3qWxQV6B1W24r4w8z5qDFhUAptix
71KhJ1LTF3O0/g7++STQ4bNsJJF1n1aWQauVXRBCchyLIcz3GO25l9679oRQ8dkv
XOdKACeXTVKaTR7TSaHWfzJmH6mwXIxgQjM1q/nk+qbAxwPjjqMQeYZn4hsbriaN
8X41BmHb3i/XwInH2ujGRgkP+MlLdSHputIm4+Lhic/Fxe4UZvH0l7bopxSDyKbC
pYZ2HYvppOybSQDzySgOrklzPRb7/lmx10sNfoIBmoTJp87302A61uJdeIfR9B+E
uwsql4CTdJOdQAsvgFdKYhHCsEG4VFGSYKPGmYyi9Y+sKtsI3ir/zIBCheSaMm8F
fifFOnZHwyL3WzLGvmqi7QfTaQYch9FnMeL1msVqsJNUCuARbBQwTjG2eF/GZ30E
onXj3X1baPRdxZyIXIvzDDzgSy/OBiVyvWGVc8PB7QTeJu4b8cnedWzUWONU0A2y
pmvy1HiAhBeX86scGaDHPScVNHFxvt7tCbQ3n80mZciK/8CYzn/WHzVg1Nwayuez
ZybdFAlygaq0eWs32h4yxGGiuplnn7kyyZgAs6RzdhXyKIGnJuvdusHXsAEzKCeh
8XvOIsVkxfEukpqECK5D+CVv2gfT9evoxRuL7Jjyz0CRSdxLZwrOrlh9y/qcquXY
pAzOhe4QIZw0eMhpCpw4bL6IO2vSDPPKg63Q2oXKKHacgmdAZ6PHHJYZy4e1mueH
gYZD8Ruo8wlGH8m++6oBwXIkznUjtfRhdV1uvKvn1Nt98XiXcumsTsdx0nrkuhHd
vAS1Vw5uGwXOx7k+RY5zb7HqK8VdKHFrukMc7CVZ9MAu1ik0rct4agNBDvqK/CxY
eOsPfS+n41nuSrihjPuiIY/XXFJPgmAUuvkaO872jlRELKhYjJXdCoKM8JvZKult
s+0dEqEuZ7lNgDhMbxgxxQwvw19mBCM6zefMzzYN+SDxV6dbgSvCQIDlZ2S5lJjl
mgEdRPJUuX2SNXZ002By6Vtkx46rmi+MuagRu6AnpgY6vb0Od+RanxIQKHPxDmsd
Bzt7sApTNaQp+F8zsjV+DRVn2Wtb/7Rz3pI4kS3rPGUIJedhSxwITm694wBd6x5Y
25yIu8rk9wF5VmcrZ/thv9Xy8Gf13J+GwC4Dej4Fz+YmVGXK9q43ZPPLpX/xGWPs
Plgui+Ib8H4etIwRji0yK9KUKRUUC2kYqUUWgyXgllvgBnMPad6gvF+24tvUsMw5
rn9ehihGULhJ1KzZu9j+TKf+x3F9uX/fqP15I8jzwggc2wjBxbnH/ECsNzkebwT/
R1r/KRSpdvteIdw/ttc//GK2G1TJVrG7Cn74WHfMIEBrsnmBzaadsMtk9g4b5Pr4
xhF8NHDT2VLNpQ/nG72o/O3iVB+gZnBXcvkhlRqKgGk9WRt9UUIlS+dbS2hEnMl7
bm+3hIo6TQjmdjzMPciyy2iK7PAnidqZl9okI0wxwREl79RYlTVMh82bkMy0wFjh
5vY+lOk7ZiR3Gh9VES5TRiu9SOM0pufiWXY9XMAvuiSv3wPh3FJUJ5oopxdtTx3e
GhktH/57D+7zp2YI2CAx4F574X/xJMH3tEpY7BbZPlK8o2tLIGN8DNeNWwtwiOuw
IsebsovZU2zSf/Pt10FzrSSulylJ+zIB2Rwss2c3tpN88I3YLlPnhIwsyenraZNl
+oHdoz2FbSq07q5OEEO2FC1JeKiJXSUNYbzbbltEJHtRePqV4pYOfhDYHD6nX4M/
9CGjp9HEcGHJSuYVBrzr8EpjeqJF5MaOxzkCyYlAui2TIhVwDxyflImXCWT1hsv/
P4/98VE5zWkjP9/8lZSgp5NLM1nTnJ4r5J3gmiZEur8NjuyLMKGMjwcvFOPlF7Wq
dlzTnbccPbAEbpJtPjTSJyk2U8fzEX++FZfsny7aAHCA576+WR/NEcDbVxNUF6Dz
O5NaHd3Np2Ey5fOpdCq4b2PmNsJhAETGG6RBql4a7sIskcSAEV79Y4AUuq20S3Nr
3vgeA9cNM6/kSTqj8LlXAGw0BUUaaZwHzU5g88XrOwGfAfWLRI5KA8aww4nUCoaB
2WXzflLucngLgJyxXQvf3NvX0IIEFD08HRcRCQFYrju+oc0ejyAUMQkAnPiwZxgO
I9iGyL0rt+2rIY1ZphHkrlQqlCLxoTsLWPBto/iQBoeoEg1KXh3DRmgxFGRp9zvC
ROGfBd7wb4K6O2JncftICuDlyxi1S0ZFkDwUry2/9HK9okvRdLz1jJVG1s4840Ey
aua6mBpS79hyKyp4//YFcVMqDUTfHcmemhZCL81pPkc8zWxiGlZE6N2OE2G7DKZr
2TWLya6i5GQFDb3lCkeDYrGNMW5RqfGEla7gAAOkiQFtz5bCaMri4+zbCYkoxEyd
OSMVEpI/0e30tEoj4l2Ns9sjTQd2IUCmcSbq8qg1wWXJfej6LWT7GtuMp49/2Eyb
uZq2q9NgINJE+Fn+K6z1054snufWVicJslcvivnYgjcvM+lVHq2QajSzT5uxWXjo
9Fto7fDcG+2P+A9w+4JwGhhJ7Y7sFupSeOBklQD3K3/hIgwDwG04gJOPtFKNNL8W
fYWe89CpOB2Qq9ulR9Yk6uciLdMxHqn3j9pSfwVNuLj3mzJxQegr0PBA2yEoP6vx
nkPwyTI6DtDTvhDeKVcGIj9/T4JAd4kWFc6uF6AswgRxOqZJ8ys4BS48BqhKMeTn
kIKD8VvApdFB2xLfWNp4dv0Wwzoh4EKpYuKk7KhwHkBV6b5glhQLe1kq5/a6owVx
b7AYAj0JYnNsjsPBbfQWeyl7Flcb4ee6nFN17KJ/L86KGqwRihMinIq9ZuAAGhXa
B7kvxc/7nJvfkzMPY4mH4JPMIO1YBJfQ59J03rZBxjU8n664XfLt1Hbf5antDtTm
D0YCNriehBCT6ZanFUzTu8BYl99+CBhG6CXop0cWcAPCBPgcUM48MmV1T1CXvU+P
JHwdBYMKhGJ7gV655NtSxUn83yJsiJTcPcw/eHdNyxmEqzBbQxerUcPAgoT3QgTI
Isxp7io+xLjVUNvRBMD1hkhomUdsVSK5doSfKC1oDNOezQn+4Xgvr+FnvwVwuPRr
ZSYh4tUCy39zL2PImTuv2EJkUOAWl7cJf/WjqYlb/8OEainLROponjNPba5F/hCQ
C6xS+x04IY+TYvbmtuZPwcMV9nZdwv2zZYE0n8enP9hc3HSzmbeNr/ml9/Qmk3bQ
6E8wpIFxpetBwyVMjYa0XUwqfOa0aM/OyawrbnyZl7Fvs2ijzCILmY4i2kKrWnbY
fb/k2MqYPndSODE4xbGyYQRJViHkLJYWl91W3vcL46bEtxdgvIYo0Vd8az/E6vaO
Q99tffhQz0s8jhAr6CpSm29nLW6PBuclYMO0s0izAT+ZIiB2Ktnp4+y4om4BHSxt
CVqqkueemdLo4wc1M0W5Qz74VW19bCVRIBEZ1wt08jMTq+oCp6OEmBqcGJe+X2yf
uQ7KMPu+7CeMQvZyu6JIsXgrno3BKfjUl8vm+Og2krku0vAlhX2xIPUEyxpBpwvP
VDbA6CHmXaUG4+QMBKtbCGBIOsgtV2S9k5iMkbQXvpYj5IpgGAgRLFaz1tB0Y0FJ
Y0+9MYEXUhSIOLry+WRDQTB4iMBtVk6LXJu54BjckfM/sGWnuDTQIKUGF795/Zjx
AwtMg91iQqcgBGrTqs2NqeGn/aH4zew3OlWRJFBBoQO9ZhhPKNNzTpuItG3U9umP
xIGL64LAMd4MO/yFxW5ywBHbdPBZwQKo36A9aoDdla0HFCGQbm7i5uJecZ5EEO8B
t2Si1Le81nt4aZy4u8xp+xftrIdm9KYwIsKWut3AE+wwhUAwPTxrCgZBjbiwUsM3
bfqfzh36UU40wGQWnyS9QQ8gPluEI6oAtFaK/gXWJW1JLFfOtkjw1Enlo6tfGpQJ
g+lepH1B5f3bt8Da5ehwLXStX5FY24buBsizjjxLPgw/ZoXjF4oh/g4PvUq1iX27
QBBw11V1QQ3uDGOAYvYDc9/BJvdlckEisJGLQy/j4ANYEL1h58KYnt617LLI87+O
RzoUKpzwM+onq3Kx2SsIfmNovsfihHk+RhBaMXDS0Meks5fcb9CaNudGxBjyBaif
S7KhlpLX3U1GQrrsPdhDA+vMf4iMdDFem8sbJmgIqWF1Of07z1nwOBYDPfs/YYAN
r0xMzhkjC05CTSqbn/qltK5unQVunFughP1KsaaFcgBv65o0+4dYbrBKWe4rJrZC
eOFvwcRYg79hHcPTkpfvl9uNKly/42+c08LYwTPR9z72SHi7NiaPOO9lgB7X2ES7
vbZWSqI7Yuo0QZu6SfjZQqQtmwsDHFshOI8bGmR5UNzLeXQciZj2hRGpedAKVvtq
n1yruymTgbXtJinBt5Oe1zzvHJj6QJ4RmGTfmhs4jRM7SuiOjewyrKzLlzzqKdX8
Cxf0Ew+eo1kcbTupdNkDotDiVCfdzeMER+b9UfiCRA7EGIAjgYBQ8glQ3dmSAAbP
oMMCaf0RtDUKEZyoa0x8o+TZ2k1amA7KivrM0yUsM4zXfXg5r+LNEEo5YCIDXonE
l8T+XlpdPHKPd1fBFU90telNM3DK16bT92eE0GqZbZur64uMHpVKHpY/kvWxU2jf
x9XDr+8CcFM14VKWTiUxuKJ/v8LfY9XpnrztX6hUt7vFBgbni/KLdB6iLxBcJvc5
SnUO0ChNCa+xtgEGZpfV6zN/bde5C6v8jAai5uCyCxmrj/lGoO959C/uWhsJD2qQ
IVS2cGqQGSvBM6ZwNCsESWulE0nZFGCS+FI04zxrDHg+zzmM8mgRyJ0saK3Xpurp
KZBdMBnlHJ1zgstBjvMWKdIxM9Z0xZqLb3/nshF4MgapX+YYJGZwZL9b+ypjZ7Yw
OBxLNwYcYclRvOQK3TXuM9nA8AROia6V5FLBnIWZ0UKKFI2klFhrfhUbkAa5mRGG
b9yoYwwUkEmsPyrW+jJNXttbAzUZEg00tVeVJaAUwtrnral7Bi6yelZ9FTRNnqts
pvyVoTW5CIsUIxMh4JG0Qr/nJbhjamoC+yhn8hf4V4JbsbaLE8kHLsMoWBYxG2ca
8Mkn+JPT9R0OoQUGOKxdllCRYn/XNAXKKBl/cu7uCdCviZyySvq5HXlmehcR4WFa
c5llR1bSaz57WcARyCV9xNi9QjcGNptUSHkN3rPogqQ8+WYy3sFL7lJHkAd8ohFW
0/R5zGYpwlHjkFuAXaaomV3vjmHpSK4VwCfVveAhegCuJg+c8ZBTHEBsXVyRSPD9
PyNX90hJ5Fd7r9pDIbsHQpW1upUe0B4Uufn6j5dnB0Mol78bkzRk+71KznQt6C6V
9RwyP4ooTjGokxlTC8DIxxNCRYleBLuFWmpZc0jDt1FzjCM0ESKRuVahVEPRfV7+
VrIW62AVrFYvMMwB1Tyfebx399+SDDAdBB2lJcLRz6I/y8AJwUkIzsTtpkGyCbb6
xy8OawoxLixAefxgWWZMc5B/BLsVPrSk85ZU9NNG2xSdg4ZQRON3+ONlceh5i1+X
ijvDq+E0Ja1tw1KeulgL7/wgnHbz603L1e7rh/6jA63SM6cfsQr06WZUqg45Kq+7
Va4UG45L+s03IoRVeyTweoPFemo0BIAa1UPME8dTgohqe/etzMh3uQILE5waT76j
g+nfkWVtR0sKSxFM4ym/GTEJqiIZvd4v0rvy7Xzc4vOSd2zoJv0KMtL7XEIdNy9O
tnpFMMx6wO7WWpkKLIBeAHAgetkPEDboQmch1TzefyUxfsk2EgChSUY3X0hOtoXm
/sDn+o0gjbmRL+A96jN+BUnUHoNVTPN7T3EzcYpzUUzpXp2cdhPzxbrc3j8iXWRG
sb1UGUtcqJ6ew1rYxWnoWyRnUChIkLYJaoGPCRpXtcmbxzs8rrbP86q/bNWDMkuG
f1qGWdJNFCINfa1Gy+4hS4EhHT7RYIdjQf2BLgSkotDrdNcIdZ3p7N+kmo+mGqAS
XYbJlYU7VKltDmjEprp5IgpMVbBWCgj+GgbXVBS4J/UMpP0TjdHuco1Zg4TTo7dk
5B0x94Pxm+Xgb5ROgN4zr1ryKcAQlzYN9CntPMsqwxB3LIfejaZ6tH6iQ9tAzRpw
hRI4A6cbM+Kk6fVn0CJssMPSezk9G1yiQTDfiJtpuKw2atLkSg7N8lJPn7/AxA+Y
kXkZt8XEzhJIj2N8r61hZZUu7mR+3SNyEtM6ejGN4uGR1gahemJ74t91uLYOiQ4r
cIvjAKTSB0XTLhYpocdkhsfk0NWQu7cWVfdaKiZ0lGDn5p0WHKjYwi2c0nhYEINE
NPcYHOCtFwt7i9QWbNeY8p60afwqHVYtchl8lqLPXNx7I/5oDYHtGk86OXBiLdid
LCWQvKbsiCwiO0Os0b8u8q2GF1gnIXPgBmA+mU26z+yQdl7QdLIV8o/cjwOJG0T+
j7sfcOdGshPRwCo9yxZ5aSW8piIUVh1uYjy7w2FiJ/2KjV/SUHOCZ7n0dQochSsC
vL/GjsXY6CnEVE2FNvN4v3tkR+ah7gu8psYnqaHaAqsAd7HvtvbwQjDtxTxvcn/h
6rtVodQoL/hmgfVN9OgqRs56lWyf5nEg3+SfpKqcvH/l2BnWsW4KUB7gmXefeJ1V
LRcv8IwRjj1XBUWMQwimfJATw1U8i6enMoRj0H8zCIDBLHE3oD0eJmYbrf3JnUoB
nQ83c105OlCkJ0TS0DWZI/yGQ41StdjPE++V3Tm22ZzMMXiPa9ry8o3RCFkQhhIi
gqgxBzClNrARnwai85fiOD26YJOOkr/JRVJutoN4LVlAkpMF1qjw7xlQd5rm9o3t
pEDMAbrRJc01fIFvJgYaoo/hLfY+bGSqDt279SV71VMm2Fwog9jaf/YAPH1JU1YC
yOdvgrv5nqql96zOZJtzbS+lJBUURj3emNnNFewKjus+8u1dwtBCKyV/cfdEBi5o
P1svcP2UGYxzuxEjuN6OBRdfHFY//uGIZCSCGj0fExN7wJFs340cEJsHK+xpY1QT
VgIyWDiarjEqSVsq68J7T9NjOE9VCSYXkayKAk9bsrZS4PYYF9YBxdlFl9WG8RJM
tWMgdiziHU2h1QcoEMMg7frt9cnUjqrl3FkcBnw0OTLjkqP1LXretfK1iDqiu1d4
MmEkm/fyhFucTX4Id23ZLhYCbnW2w6AvCJWNCmOi6LgZYMijYsn4bDsKU7oCNIO0
jZxpaDINDams9pkS4LLCIGcSzB41n26ba/hgx5wQVIc8NN7gPnGrOo3F4LFhV0V2
Oh2OuI+gEdCgo3unJGphMMQiIXQR2nWNxBo9T4QTx/AJiyjHVFOprXEji4yoMsur
XJW06R+jYCVG0d9pzJZMYsk5URcrbLCFA7N00uO+cs/knA6eSo0XXJxZLhOZTyPw
VWNZ4w/fpMeYBmQNIWiKZ24Hk+HDi2p5pcy9v0LTQEq2BqY+czaIyQDHpzoYDOgw
x5GW/v+M8m+ZJCNyDN4u0GLWDBK5cMyK5hLPimxlq/LfCZsxwrup4WSMp6xARYQl
AKdBL9ADaJpAEEpZwkQupmKgKPkOZw0mDt9QyyT64egHZEYzI9rZlC7fsRhadFSF
8q6v18HKXIspUFgGudoneNTAk5ogBpII7v+i69O61y226Kq3MKskMF3s7RdDxN8N
H/EqebXNFxX2+4P+wu9m99YKdgM1jgx5v2Au0dp1Z8TuUa9QWdNzqOASsyF0CIuR
qImriQ2/bSeKBmnNM6+O9XE9lQaALIoNwAhtvic5+SL9WWQpZIXnzV0BbTb0pCnf
GYdkq9emNRnYTSAiovTu9XdJnWTGLcSFBp9rxF/Zlwbl/s0KdnurHK5GnQkkrVfC
77XyBVFR/aHMn7d3owP1G3nYJRpQhuu6Q66TOH1tKOVWHE7jTLOHFrNmtl+e1cSL
9rq9k26qLFmgclen4aYoTkMB1NQNH9Z4mwWnKt6eZhKYpTNGnV9YCcBeK5gX8rAU
GYZjGROCYvKYxA6UUEkjiMP54svAXyYlrWSyVYYj1KRM5ckGhVB+FFHudl4Nxv2v
LIjybtAm9LB7kiDVmSWnwJPBab4HUzR342T/zNAlxb4QxG0Er9ZVTrs3dBbO4vEB
8EU6RVSdr4QpQ8k+G+zGqDN8U6YjjdL3BKTDEyvtv2U/sJVf+KZfhfoqDnMvwwdI
fzv+OLmxW8prA7gxVoDmaQchvAiFqebVqZgtDL+l5FbUPVdbUayTPVdgg2KSMVvJ
k/zizXxlao7pR/qgdkq1f6EYW7/Husf9UU4qOr/+ymUFIZj32tAMf/gBQi8GYpbT
rmn2t8WC3eZe7eGDrRMjAZ66suOdp2xqgEYP/79rpB77E6xBvXzEgyPVW2H4wMFh
idJSN+jTkYe5X6wYNvY/JBNqfuUSEjasy5SM+2ldKeSfWxi/3GlWtGXnrctCvXmV
zNO9IaKOOD7TvwhrQbdPqpsg+F0M/tByPOZQgk++Maf0JcXLiQaxw5N4gzW3QoQN
IpfLalOeKeDzrVLjlrudcDUacqnTGojRR5yXRvN4oQkkUSA23zHW08JNBARCMcRc
drbnzkNxcvNQ3N0Xs4nurzq5pq9/ZqeYnQe6hxjHe8255I2aA+KzaNw6kTdLfGjS
QjvAXAl237rlEsG0RTVDIDZlT+Mh5AJEscgPaTytLraTGovddq8Bd7vG050CS4wx
jHH+W954V/nirQdMASatrW7+YHSev/mP53RaZyW1GmvbqeypjGGD/ZShBWXqkuPv
ksV9rqHpuXbVbU0J6hQwEXvcEB2r+xXNxAR8xC84J0qrf53a/FvYm0VyXlq/LTsS
q51KD1OBswF4KTeMCVVYEP4wHtN9kBBoXE7dPHp3pFLP4dPtZMWWvjczjD3Er4NF
1BXwLLQi9knAJCfd9PgtRipaIxNvJFod3bN+v7B+4agjyB/Rwqnsg1DTGEPrAJ2C
xa4F0Bo9gWB2yewZEZrTejwkUZ5Iamsnhcgtj4ChExQE4Yfj98Jw16BEoZwQXl15
aErB7/8UVyAzym2n54hV1is78vwjhS9EB79cSs5015vh8Lg8z8/n9o5MYkHnfR8l
1OqEZr/4ZsphGk22iS3c2HBBBW/RGUTutAIg8jHDl6pCMggEmPkk7CoawEWwj/ki
urbsp4dtTAObpFh70J8aIGzIP3oWmd4FfOONQaIkpwnbS04UYrAu/XT2Upu9xz8b
ARuIh4AeGfIH+kVzNXg95LJihvWng8bXMPMlhNdXgcROeOJCPpqxZvX14qeq6nyL
AsDd2uR8kg9xpN24dwOnBpJEtbJnLvAH6pvq8RGB4x6Dqe6jYhOGcgeUaS05TYE4
ijkdx+CD0D/3P7sAjjJvVhcDXxlMVh6efHw7gB4T5mwQS58BjO87Rhc6SRuCA2oc
k3vVJonkokofLMY/CdJnLcsi4gjuwPOqWntr5d8nTpcGkfjwearba+ERDXQE3nEr
qSWa2CDgQ4dxQPAVv0PbmsT8vn2dxw+RFyLYKgJORbK1Oe7BsCe9F8YhhqN5FsXy
hrkvBDvQTJON9+tlJScwWQ9B4tD/Lg81JOmRwDyAaA4m4QJa0q6nMbxpLopZMNtB
dGpzOZSs8WRJKOKzRtbDPOrzu77GVnJVDmp70HBBvuYfSEw8xXoofoyPl0B7O17S
hFi33HA2ee3XxKNoGet8CDbRCNdF/z/kIweqWS4Im0y3Jf0LVRtnPrcwqrDOBO7T
czbHYVb70eSb2RjsQ2m4cU1ufn1ZcS3ZbhS0L3bXeVjxYc1zrtA28qpZOVOxNAlX
7fczxxW0tVWyqffFulQ2Y9unClD4kWONxSUp8zzv8ZkVBCzWwvjbyglnGDGWC6yb
1BcdKAtgPVrmrOP8sAsyZpfPEqviUwVkxpUmRbOhZEa4ooqJ6TG8DwXlESaSWLIx
DhQczhXw6eEzbM5gDBbW4i4YwIi1fPz4bHPrvBYBLgjlsLuqD4x+6L+8PAVayjTP
tWlwpPVxM979gV9xTp7ZIyOL2d4wVicHaw3b1GVhFtlm8/rgH56TpcFj3DLQ26jx
07//ZB1eV/YMVOVmSLfJtJI6qc+AytMc/rHSD5PfG0HfAF8jmE1vyC8q+bfCaGUP
m9eBI6mLbncF7xR/7IVGtqvDtBW2tSrBXR0rHOrIYqRKeOw+GgaJfdDr2sH1NMep
UIjN6wa1IjrH7zN3fAh7ZMcGJERx4ziPf+Ldp98ZKUwckIQFsOWbPQYMeloETCyw
91jl4T8F4o4FGetBtHSBUakDrh1MJ+y/MIOUQMVxEp5Lzckj4J2itUDyROtZ8m+n
GzyrZAeG3hHSVQ2HNLAII1f/OUAhxqV3k8J+ECH88lQc2z/CU4X1w3Db5TsN7fca
R2MzVosAvWLCkRWGSrG3uu1k+GUXZlUZYEEU9cxJITB5yYzpnC509uxZNPQrhvXZ
f7OaEXPahk7iTvYu/AqJ3KY5BHJIc6aU7zhxvTtrDPyNPjRAbbhTDcaNyT0k7SQU
mqj2pyws0mCURHBgll9eUzc26+sPqSNaC0JCGVkNDJCVxPCeHw8YoOusru5wO91o
UpVnqihH1E2jEOLJNA0h7Dnpz175y7ps0GLHF9K7pcjuEWclUz8zPnZk22bciaJ5
zufrwCiJ+4gPkuVVIwbI4C1SPWPM1QXSZWbwmo5KjBR+vIM//FEvVB1gynXnz9WV
FSJ3HNP7oLDsS6pCnklYexij0RlFpqLwu1HEDypuEevajseSBLQrlShbcLjER6/I
MLpDl0pqVKD0TZUQWUwBAAR+61WUHvhsBdeVreoIpSWXQT8zmagSi10CfMR2YoIg
F6dbQ+S0W9VD0nn+dIq9jAqPfbpf6Bu9BRuQc2tk5weTZI5f6fUCNziEH9gd7gR2
R0jflBqkukXKFK3DIAV0Z94TKW/J1869kddCgNkhrpgZ+apOgcu67lC5ZuGffyjF
QJyGhq9dhS6dAKqdeDTydI8os1t0AQLd8efoJlY8RR5/TBrNzeBDLoSs644DQXt8
ePBEoR8tjRiqbg3S3cmsyW7AGz4Cc9NYBTLZ6UokKnpwVzt0Tgvxxi5sJ91hsEAy
AVJdunHdyXJVvcQsCvkyFBdWyyerpq/j8R90r3+QoU68UTU9lpdkd3N+uxTuflUv
o4Jr/XggHz7IEBCxMTMzISb8C/w+P2Y5UhGqi3NXjby0ejtvsrqG7w8at6uWyHp8
6Mcs6JnRz80jNLgWvAh/tWyb/Hj2K5ToZTD5JgfpSrK0YTWlyGoXi5Y5Vpx6K2zI
EOy70X8ApX03J5EEQBoMUtqNY0POOcMf2g1I5D8QGh8aMA8oQxW4PKfDjfRUuYDR
T7hipe08KEuzivBh9zl+SOcbl3S0WkSCW2JUut0WOSV4GXblNB8dhCpuSHE3dp+o
7Gd0n0HWi6/0PjtknRmfQCmCjvTnZ9IQgw8RY8V93CEz6XplO0iaWTPwRoikbjl7
A//UlP/UKMoWm35eUDb1hK+4hMfAa+srDT4rKeGIbWkZq+UrYc3FWrQfAwkB17XH
axdflSU0IIGuzzmLwRFWslqfGuKIO6AbS6EHQcbBkEmBZzet0zeiDGW9Nek/uE8N
sN962uba38EZ+DzfprgZk8LBSJey4eePLBKamsV6xKcxBYnJRTQbdXv1S8bhINrt
gO4k0sOh9MbkYfxtV/NUp2s85zIC6lQhiK4khHFDEo0MILBhO/zokcGYI06JFWZ7
IiJGRVZUalvU6AorVCdCoXcilfI5QyfZgCl8n8R8YfGsx1Roh0yu4jfNRIDYhWsd
WB56pKQ2AzskQN1yclCk0b6KXpy+u/Gefz6UFKMOvUwT+siT2XX+f5qyzvRO/9Fj
WUK7O1dVIJOq6DAJmQ8jWXLuHfMjybbNB5UldLGEFsvLi32gXE/e5T3hjfFgcpPJ
f0KFEYdjNeeU3pX0TPAII9gDZYJpfx/oa+uH4a3vay9NflhhCFBklyCD828A3ba/
uFv5KzhgPP3fpTtycgGOL/nwmr3Tva4MnUxt+nWdrdeTq16V1SHSdGT1bfRaKYpK
Eze51gvHrrcb0M6lEPDNIpruMYy+DquTZU8tCAuej622k1EJ7Ct0NjT2HbCRWySM
FMg6uQzXRxeJshcFt3OO7mLwvVRAKRsyFHS2ywjgts9Kcxp1TuH8ra1djLa2FXcd
MIVIL9FngdIXcYIp4WKzgPCpNd90GZe6zFTW4qkZbKSDQrPZn+Isug+nto6+p8/e
jNB08Bb7QSScQuUxDnwB6jsH/HnHTDgeBmnDWXskkCsSV5sHKLqjYdKsC55v2Xaw
nXJSxMRNfbQVeuBDafCGDao7voVxRcjzf1UOHn9xk5f91L6TR+VwcbMqqWa8b0gV
1H4apGR2qHYjp86598PrdEWl+NIb9YjUvjHd/wQnbISMSK4oMn2tnaVxiDibSvZe
hKYkbV6hvST6eOA1Kvfv643HLpEyvMa/DKTCry2s2nsdCLn1P5reaAVjIQwY0Bvq
8+lbkGk7PQ18L73Eu93Q56UPrgoiLzdrAWoOxnKBCGFlVVjyBnnxPpHdDontX34I
cy/StV+stHIgSI7CyKHdfOWkpBKVUgahytnk8YsBHc95OeSEGsKjtnAmTRT2tVps
XePGgZdsRXqhlO5iHCuYJAXDuevxCq5mJ5psukrK0ElGyMovUzOqlbah6+63fOJ2
10X6LUl+eY3IDChjCkOp87ZapBh+fcm/1CB1nWauUkrInyqTHoKZftUIvsx1r+xV
BbgQXra4p7NwAGM8Q99xCkTRw5RVaEmwIykHIFhZxOhLOl+2MkMWrBJmZWIWp/0U
5tjfLdTUCxgo64hVloNvHkqqAt2uzeQCkNXlO8+2/0K8eWEpOGgG3Y8xy1pNHqUi
ViYyBoMWfVbhmxm+Bf2a7GPLQc7v6PvxpW1/Fj2UunzobMvo0bT/wGGvfaI/hn1o
703SgdfBjtkkUL4/9v+E0RWioq/p3nY3J044q4mUQe9jV7n2J8fbP1TpRyOIOs8w
8XWdG2sKBpvSOo93W5kINVC5MwKr9Ny7Ft87EqP8Sz9QN2+JxwmiZnRqXAuEjT1s
/Wgr008FjIyagV+KIrkO1k0uePSI52wbbZ9ubJLR8EEFHK9Lwmz5UWvJHU8Il2CK
nMlWJv0nSyvbXKqt0gIk9A0L2/qJn28bXFgZKOWufEpmE4O7sROC7bLNHc3KwWLQ
m8J8aGZkQbWMtnSrwv1Twf7WZ9SktVB/tlEsI1py0hPJ9h9ksPqFuD3Nn71i7nCK
VYLN9bUNVk9lUy2z2QMWVzjswOLR8FUwBvY/091tiLa/qrYrmZayB4Z0nQdSpvUG
yT4kyRu3dk0gKgKW+EPJqAiRWrua3ZlT1wfUyMPZ/UDnReSYAfSGRTP38BqdAdEw
K7god0uF9GLG5m9zGVV/5hMAotW+2r3x0X3qUt0tX8If1n4JptmTds05iJImtc20
aB7o9jPL6cCPxS+24tMKSLhr8qAvE2n6Q9h2l75aXYP78FbT07oZrooJf359la0C
aNUC2QQFDkn0VIYnLWBChSOtRC37I4heYVwCc8MVFLKDbcL2wdfpxMLJd/78wN8w
9g7DQf1H2uZNX3hGeCqwj7qmMa7fLXkbvsKT9OyCLYwe70sYJiSXDoLc5Nms3yse
/JB3bxtKuH6BsRZHmP360V1mFS36l+AH/Zznz9xHNbTbHRR2AbhkWZkJeTFkkBbj
AbLXjYN1x3KExj912+6CvaeyJqxjffP344B1NqgbeGfM12MMgf7KMki8tc6EQiKb
v4tzks4yoWZqmW7XkdU9+Kt08Rzko7v2aDQ3SCybJRl6opJcUASTG9UgoFhVOwQZ
+r4X75mVp4PmG9SOAfnkPleATHiQkra8GdeT2nPZFncwjlIc0yeVbHcwxvotgM6u
OPCO3ATQZwjkggDrnHD+/gV/N236GP47AYZwLQu9990LP4dtQh/iqulALEB5TW+A
49GY4QtUPHWd/VNmmCTo/d4ZNd2e2ahN5IaEQ2DZwSzpEtKaVOlxQCUdZr5VWnC4
p9XQl2Lu0MG9mN2DeKi9CpVkC/GXUI08kQiON1tOtyYrAI873qfHEd8HLouO4mbF
cJa6hMWjUHrs9qUq7E1XNw6ZXSOCpKxPno06OHkg7hhoGj3eEA5mfWB1z6xIijDY
/Bh7yLT6StRH8iuZnLijsl50Sc9/0BPTZ+/FDh50XkBWX5Eiv9NhdOoAMfVaKXQ7
b2rRM8bsjYEBgcNAskQuJKcrE5RXZNMp4rOfk3CsIBmM1KNzTRUDOm+jDVzqoIeb
CF9nCA+M3h5GxYGXHR4u/h1BF0QsWt3zsrCqthhGF40zQw7yOZdHO7ZpViPxolrR
XgzneZFM0VR714x5r0k4WlMTzT/4E1i14YR8s4Bp8TEGzYViasMGPBbIYA16h2Ld
YK1e5lSOhIejND7kGLS5bm51mnUAxudbZX/JVHeB7SlrwMOratHtt9Rzbsjmw4rO
eyx0nePQEsXz6V7zFpX75lHGar5zK08+oB80FYc6ZUilbl5fWk1q0YSQYn46IooF
ujzAMjN9IY80jYYi4Htc4c9+9VmqHir4cGcMQ72FlhWpCysKGIghk2iYT7FMrG4I
ifiV8upP5QAllETcUv79SOyS0dNWwpGlGiM4HFFNA7q0+o/ILkBEWgq+vE421q3o
tvRyxFUCG2qSKJTnoIbkv7B+xnR1VobKyqSEEWgCCb7Kxd5eL9fKWAZqRql+TsNH
ZXqOtFOQSX9VXOvEXJN7AzamlQDctsWiFOphg2sASjOBLBVtHmZd0xomqqtjKXHG
nYYSS5kqWz3a+oQ7xdGhQAh1TXqEblL/zez0nFpaatJTZIAjxKyVsCMjN0pnFjIc
GQinuaWnoPTnzdOGvW7HoaFSPRBXcs04MlA24a7HV5aWCycGkRr6njAvlgmzBqRq
mWnBJIfD9K8pdrdgi2YZafL3fpDltfD+tXkX+bzQXqQr1bCxnPTYAdYGsc+89yxp
L5S3DENIKHhx5hFq7kLXb7bWjttGn3RzgI7YA2Mb4KbyN43unkPbQebDBrWoIf/r
mbBXn7hUyogqzjUOpwjJfKuqvaoSWjMFsN67qT7Qa95HvKZeCQGU3KsRP6B1oCvz
eplUol4C3wvqgcsX0vHPZOshrjnXb0WiM2b/xYSxsMgH2WncSKqkrlg62+2TdZv7
Ekwb5bOgrOjhzmWiHWhbKrTezd9FqsfAIJTmTqmLidF9qeyn/uOzc57mbY1wUWh+
KST2ngZi+ygK9T1p5q7aKXDQ3eXzIaoX9RuQmbhUTmwQk2YGOP3P6+fEZmzSYXxX
nxACVpQP7whormmW3kVLydhUbDlMrPffAXr8Er6WBiNOTiGH8aNMt5un345BcqUo
RfER31VhsIu1EZDWvubnkwUjSS400XSRnlgmWwi+4vCDkCs/7rV2FymTH0IDvdRS
O0LIhPagABK5Jh9Cfrp3nRpVrV89czwKOyLqL/m7rd8r4qjFBiAxM5vDi/9KWaOy
mYiZ4f+uR+48pjjYWj02RdbcsrYSax/A596ytz9GvIwvSPyabvirvMwt+3HElFZl
QiB2fKQqG8NkkOnZRpJrtTlDprp+E7V4i8H1K5r6bJLaoekCevaE0/C9dQve1rKb
mwpPC9lsqdxjA2yh8EU5WD0i7F0GOavu8BP3PHN8MV/xgQ7PbiK2pVNaNwxk56Lb
br/VsS1vkQnLivQKh0o6fJ66Jn7VZXkJVhKjWGAjufa6kHJDlbu3MIEsQQsTpl42
NwCdlx1RMJWnPYzS+nZM4EAiF+pqoiId0MXlhHH4C/x6CJFMdTLFF+TQ5bapKGfj
Fkc5JR9toUVYuBtrl69qhj80+kGc8FEB2q8fbRN+z+4ibOzN6RTToVfGMoL+VvP+
kXZhrWSJ1bE0ynqfwtrgSvGE8RNSUMI6z66CILiKtAEXOBio7eClyTJDorcMt+Ew
S94BusysQYTtKll4/bxbin8Vg6j/3GHCi3egvZ9jeCBFS2Dff06J8IaQXqce3/+9
MkWW5h/cOXiTyhpoKWNNRbjcOVw1eZnpZ2A1YLM0iOFjIvmITZvEzpD7wFvTzwdK
K2+hWYsTQ1wOJ+EKjus1OtyLkkJe7OGe0ltXbBtqj86xF3NlbKSFIHsApBSEe0XM
EeEOJg6CDLYPEWwXZE0dHNWoi7Y4F2M6+RZxvNY4KJWckifL7VKbwhqg+AZ9OoJq
nYnKbK0/zRXizOG99ON8R63FW4PTWphBReV3VPBmy49YzyDYfjZNzDfkYu02sWEa
3NkDDDHQ8aqeLK+TY0gl5/+HGe0Nxk75BO+ZVRZd7RnM8JnclzqBWRZvA5LOpO3L
mv1gfRBSEhoPxAHB4U6gBMWL1jvY9+Gw4HY60IDsmXXznEXNeYrrHdWNzx+eM0mh
jkqSNGytv49QFOXNFQFBXYt/u69ajPQmhQEvRTA1n0fIpsd8ZnMrun6B4DRD0Jtv
RlgfcaIugVvnOjGHt6eCCmyYN4CslL9MH2+N5KcahESyMe8U5k6grUEynij3522s
+5oCKkCJWX5Ry4R5h/+wLdZifKi94+GUIs7zNLSQGQFB1MtqKsCp9qGNah4IoR/H
3zATyIStPn2wgfGhNinZ3xM2x85LDT7GNIhiY2YssdKoASA0RGBiKBYApuIGqatB
yYwyb96Z3PtQaXJVwM6AjRz2p26dgiesdDOC1OBFZBDvdITKUmCe/kafkWanfIYa
yNZcXjPjMKa5kUYZLt+0gmCTXXfeg/xQy14lRC7yGvOLi5WJndLGgUOh0kEgvR93
0lKy7hb8XE4Z2usgPsBwC3G0KLl2gqgrEbmuyu8WzHw7qGfdyhsVQVqqLNqjz4PA
wmkr6r2GMcTvnTPHaHM7f62fDvoFV/1o4gufQIoAn3E2SGBNLMGT9CmbW2LwzP3w
at6nGbZ5DNI6DgGTbdLYzbPncVXm/bVuqP7xF3DwKe0telqSJ6I//vy3/TM+WB+/
qsPkpmJTtot7SHn8r/+1hrBFMJh9e7VCoS0nBrs3kwcogy7gl2Vq7hR79t+rTJMa
MgVLXCL6JK17wiQzT9W7giROLYg9IrvpgVVFiu/jSTjxEQWsHLivuythdlutfx1S
tglZGiAEpJpjVHPumpX+34jEbkZipR+bu+S86r2vkRVvNhia6lqOkIo4HPa5aXIo
PVqpFAj/Ii0VbLkhs+dphSKjclLrqfkBKcJ3TrkK2wD1gIQ/qnGpMS6Fl0dVWjN8
JGAyPCpnKKc5CfCaboXwR7eU5q1OL9E3xz2Sy0fGqnfEZaG8vLAUMHLdrc7zrb0R
Co2tTGRSZc2bGvMKqWqIxmoSy0XEMhVYFat/6UKCiEK+tiOT5on7LKivTlDX3755
ipx/VrjDoU4afwirj/txH5hx+e0PQNGbTVzHnG7WyloN575I+E2EfJMMfcFC07WH
01lGZsWj37UhoFwvduKb67EWRDrItPvN3fr8KQnJmdUoiiD2MRU8hTR+8spDGB5/
YLtm+RuaBwvrCZojhkez/KH6EgSpGEiR5H2R4Bmy7VAsmpxLpZexzWtRd8PxShld
FzpRuFdROtxgsf0Q/ofNW6K6luiKCNQ2tra3alS/l+1Gwuwc8TEd3qdNNfFbYHST
8n/uLoUX5Y3CMdDPHyuL/iZJ0wHj3EjNRnQmKU6sJa3lVADZrM4+Qu0Kg9ygPIK7
VQSwKhAzavWrT2w45kZJRT3ErOEOO+Kv3HHw0Obn20FrDN+M4nOhAn9rxx0qZJXe
WAABtDtAzI0YPrZB17Ik+hwEzKXcVQ/ioTw8tSxlhlD9Mw15mTnWnuUt6qyk5p0a
qjX1Wb7wKWJCxPN9oVtsdMUnDyWjXYQ24OQVG3drZm00HwtntDH61HJ+FS6xzyNm
YDsUQbiU0w6hdaWzIsKY4BoRjhqYXHGj+VpMFlubRvx017MA9SgtS77hAc9LRMQX
tmQ+PBrsgC8EHjB5LB/wogEOefuBZlypou+BR47FS+PaaRhAa1JgpLBaJbiMjc8k
7b7nGiu/bYxmWBeOBtMU7DglVFIg1fAy8b2YWFLGTpKlnM+NfqnGW2J1ImmDpf7e
Hla6tUmIzKxZncHEImCIVODRpvfMg9sOQ7LaznoTxQpsj3hefC7JOOjS4DYuw80E
vuThwreJ03PAIRF+5vAL8HbhvJsoDuCNu2Gu4nrguk5JAiH+JuO/yVG5Y8/gHfNO
U11BEALq1Q9ZEuhQ0Y3t7Zg1oPna7TrEjb3yCqBFXC7suqfLi18L6mIJ+uwXllk4
oGRczIIYWKmACU2n03MPD0IB1dApJqoi+r4EaDbBGabSNIgXt+cz0UkpQnkh7lAI
hQ2J+zHti/nD/7dIgtbR+EMerxLE76Z/rh4DVRCl+udC/ApLI35aCnl0t9rQJ69B
UzBkiRBfw/TZ00DeqnI9LbxSp1o6/bABhnq60B1JWOCG1ARoFxey/ZwFHiyy66kp
OREBNcVHhCneBjfscRJm7GQjwx5CpMNaX7IQGijQ+JDzDB+uGBzDC6U1C73xEQtA
owYKm/z7Q0kQh+H+DwFYEWMsvbmKJbnRcLhY3uxYMZxGV/MJi79nkUpes45U12YS
6HrZLgMZD6BA9v4cjqhnARzQCS/Crn+7wCeieEy+zW/FTFFKqIohFtP7M5vQtOG/
MUKfmUnap1on6FoCgObA3mG9o8sD5aGqrDA6AllhxvKcGhtbw6Ri2HLsBKBHw7ZZ
jvTRMM6YbpB8GbL1FxDUNAMO+ioNy3OezH9ZpbvqGjIjmVWIbZ6nO4F5E8YJSlFF
gwuyN5yrXNYjg0nzBjU7btOeefNo2CncjQUIsqhZ2TMErBtU/LyHTXMffSBR60Jh
Glmb4qh5eJn1WYu7ZDzPft28n3qSXyrtZLjwcIf6dwV90X7Em/8blB6Bm6q4beLh
NyATEaBB7BWjBRwyymanGTHaQ8GREKFtacJT99IoQPGn5fEv2Sytq3O6tvafJqsh
eLmdpQ5pZ15RXKp9mNx5ZPVR2mB3si8WFU4rylAZUSgs8QZmqUZYjoEqkm0if0P9
vhQsAJslml4FUbGawfiCMX0pKAdEmxUaZ60940f5uaIKEm0hSKvklOWAaJ+M5/yx
8CFzyMxa1kUq8Fkdc0Tq0ziebwtm0J3MYCFK8Ce0n3P3+Qi4ldyvldPBSaPN/8/N
S0DUS0msKpw4cL4l7vej7RYcGJVaZod/6L1O54YT7MSZ6n1vuG5lZ32BU047Zmja
RrsP55AqrTX25egv7VE8P/x9esqYvQ086XwCg0tpQONoApb+nTdlVGpHAEs6xCqd
5vHJy4++pJmASfIAi7mbVjgnwWTOpaaCjxWlRw6dAZKMQnWoOjRNbmD4NrIOX2LD
MHbgst3pENFvQDIjsjCmmEUeC6j41i85OpVSU5DGv/yBFNz80f2uYPkOprZkp3hQ
ebJv1vonRcNfo0DqtMBj7K1vLtQZJ8dzkkmtU9rdYtZiXRn4bUeaCYjvk3rSvwZr
Ct7crv7FW67PcxhsO0qS8ma3/rbhlyJOcMCQPXO/+mvjXBRN9CSCgEa3ed0F1IUk
gFiLVJAeev0bQDBVHnhOWcrsmFxUr55/oq2nXX3+P1+W/uYrsXA6r3iZdCuLB/gt
UjKhTVD2PbbgsY8m1DQaXNxcfTleNILTPoyu3a3oC2lWj6k+qsCF5X3Z4bIzw5HI
/EV7WKRwNWK9zq/v/nNrfstcFAojAf4DSXpN1N7dMZRryIdPp0lAVIKPyE8n5Xzy
OmgMoDA4ListYLUv48W6fIJwHny8XOvxbfZvkugesKYZzXEOnOkJGS+cQhAvgfhX
mIcCcbSsDIzRJNhIEBfYibrTc82BB/ciE9Xj9v8tDXteuNuvsU3afR6GrLclnkf/
y3CY8tWspGyUJ1jVR9S9cnKTYntMAftzE4R0ExAwlFqNvAwQCwZsICifZA+bKsEy
rYFKtJaFRCn0X7In2tn3u3/sLXHJjAF7jaxJGAaTpC/z8Hb6F2gmX00CxSIOnPWj
vkT2EmAno303b/JXrJkDGtghNAr/x51+QM/rrys29rxlzokt6XD1tZNzQS70qn80
2b8JKjT/SOHT/wPzlbanXycp2e2scwh7TS2gzuU3KbFvur+N4I/Ead78vCSQVjNw
HpLincjWU9y1pUZCVRiQp4WIrqWGDWsQJPGIqfU+r161mEn5aVkQaGRSc7zN9E8o
E4t+TXdel2icmq7M4tDx19urCd4DSYV5CWZpZVeOk4fdn4HVr2oZN7My8bt37WDO
AuP+7bvgzdtTHOebawKS/qL7dnbmMYAfLeZR1+0WOowutwxtMdKmPXbHB5JEwLew
ETXr2DT5UqupzgJoORYnoFiZuCI06dzfDZGkTMajd6dnsIUZUPJO/8nXmT2mvYum
KZGBue1FKXdNvsKLPvpSxns0Iv67J7vxue9zhf6FdodF74HLh4zCA/hgoenXIiGW
xYh+29UEQfijBMpySXPLt358YeY98kt6AxEwk9j2SMmDALFrWlVuKcMHx6ETWmkJ
5tbKQgWxFAiHpo8Ebs+O6s7fRulw6DB+hG32VECHERUbcBAHt/1h5xjg84DvClSh
qnl1JrJEoI+/NBznWzx7mRBy6if81Nl7/J9FnSIm9kGhqKIid3OWLkmi4ub5+1pY
tAA4M1MpBVLdNoArVJ/QS9cJA4AGuVJ/P9r/vcXBkesLje+f4iTLurudAyHk97Ht
uasa3kNk4Ie6AyZVsxATSaASqnoUvr16/xw49s6yqLkXCcMrWLa3XnlxxBtK+bm4
0hxC/6llYEK9A00K1dNOhJoK+YiZMc+hW21D0KNO+3QvKE/Swi9mIJoqscGi5UY6
0PCQPsG30Ne7/cppXrH2kNhqR2F2J6gB9AfAq5VmYwrvvMNFreF6bBmAtHw3Sft6
UPpXNi40DQlAkfil3sgkeIF+MO/2G3BJvWlCPxtpCeMsd6L7uH5jDAs1oU0clmR0
pQSMNWoZtQmhZXYYQzrl42TOjP+Y8s2rLom8LFP10TzFeV/MUyDKd+bBPqzmZh8N
+31EO0iOHjTa618AHc/I8Sv22jR7sFx9/vMqueIe89T9RSPATQlHUIE2UUezcSoh
nSaKprIohVIYxOLC4RrHXHEKh/KibdQIgNzGHT0/oAfADQQQqckucR7LlzvEkts+
L9zo6ML25YpLULN+S5Vkqo1D0F9NqURzSRbzptC8EZUu9eIKCYDvZa+GS1B49UDf
P7s+WgWvWuGr0WKPNWdle7QNwfBeL5enBSxD0hB0N+mNYEFBm8mhMNjD9UaGx5D8
KVaEkoJ+2T4WinPeGihKmeA6hlcuk6ehOdlAp/O+zxHVw6fXr+gprGAyPkt5gBlT
RK0XSnYhAfnvx21Ao3kw97gZD9QGIx5qwgmsbafWIQjcwcxwPbuS7uVK6g5RKy5h
ZXDoEIbZLpGMQyl9oZpxp7+sfWmonM1mzKXQM7mVfek+b2cziyVT3m4C1xUzr2Po
Pn8vu9QdC/lTZ/ccLxaVB04afQjhQd1XC9eFhlcxIQmjyfvq3AzDex4xdfI5KBPA
mVe2lInLymW7dkD9PI71V6lrb83ihm9mNFdtlkRjw1sij78MZ+QxfruccLMUPCmx
ZBX8mBUUH1NhV/XvK1JBELOsUhzlqOH+Azkni71T5WU9Go4Qv88U508viYbOPv+q
aaxAOTodKUPXLXNSZK/6BMbE6SOm1jpTEogTCN+IcnYQrJC86FI6KvRQMavmZ6+Y
8zDA6T8eMIuBw0JucWS7AfcINuWuHUf8Usn3qJL/Iap0BN1TOgeXyhawImuj8vXT
87kEKSgQJLGzYT+XOxfikM7c7RAtBuvDLe64b7yPuKa4aOoxs0fa57BJqRTnyYQu
3Vxp7VGZZ+/aydFjePp1l3LT4vFW4BofU9UPr2pccs5uIITjuvJ5vgqQRqgYnXbY
v8b47n3727gMJ0RnHims/dOvMejfaT1GpOH1cZUwZQO2bT3uWsUmizXYzEdkAf5d
8nhbNpLiU9NeBnIkLU95Eac4jaK8lP3H4gPj3TvnxdbNVPDuAyLxVFOkViplmLZo
2SqXnacovu/Fajbv81McKowHHWk/VDXj0YuiemmkGySHiT3T50qqMfjtTVEHZb3W
ReC1dY5s+gMH84sHTqM8duUlx3MNqbmBVb1b8tR4E5LjBDo0w4/hANnMiG5qJ2rn
7YN1UOvLS/tvzd9OQDje/dErFtKjtHwv86JzqckXVxoPLvQisTNW94iX6WtHEu8l
TiMb1xQPrv9FwUQhCr/T4i6eN29Faid4OeJmdxK6s7e7i+RjaZSuAw4BwZVz4Evg
8KslhcGIoCw8+VB+dhiHQsCfN5y4xvm4E9F2QQBXUuUUmJuRwo/VEITnOhKmrNxg
YMqS0Ve4lZH9ZxxEW07u2ZkFkF8bYA8UH912mSO1HpJ/h0mYXzu2EykpY7NoaEJy
hMCLnAQsdMK5ra2mvsv+xiGGnFU4SGzhZSRDA6k+HlrhhhpKCznF2Woekre31g39
8i3yL+1/nq9PkP05lP+kj/Hf41Q1yBCaPcW94cIYBPBFXojymhOnV27FXysyAmvQ
GCsUC9gVNcr3LTJn4WOnPO0p+NMZOwtn+NJG7FmQ3s8qW5lMVAhp4Sy3vgS27cEJ
7Mn2JG4g6ogbt5TL0F6Myrcic9XhcUvIxuEzSLrsyYACjV4hjdbOm3CNk7coFt8p
1LxU2sykc0UJQKavZvAH/6E9yTD55GTeW+qutx04foZIR4Vn3wGSSvZStuxp/1ug
INjcm0WLpsv07LcAx+TCdeW/h1G2qFPl91FaQ1FqhPqL6w0rEit4lwYI0yXYl2AS
kEvS6wlAFTLFaks6J9YcaOA+rcqoOGV9bDuvx0FXjihs3dXDOp22/LhvuayD42XW
Nk7xDD1yidTCIqLbhJ1X0q1eJ7T7/pHih0ANT7eioNbX/yrUePnQJyAQWO+Uq+Vz
aRXneZqUf5bKA8JIM1FUuJVh4Tua8SaV400ceMlcGh8yOb1qO+dG3KnZxIISKD0P
JLsd1NrIcy2yP0j/nGvr/UZebuMLEOFAUIT8LGahUKJmS13nOQBi/moUcFhcFmc1
6npWKhHqPIeLo7d2c2nQD08PaFDRxCHECeGD+SVV3wEZHm7mFwaNcF8BONNZKhPf
/J7ZdAjGGYeFZNqVBeT/a0xayZV68+ov8/twcfDUl1WcBqvny9SLpDFJ27eK+slz
SSQqxBEo9nd91a5qUHLAojGdqY2iiEg+yjcjn7u3aTzpGsfm2wSO7hRmKrEn24FO
p9JkG9ZjqFIsg0/SX1Z4xPQcLmf8zojaBYO4TCZbFcSUry7TprM5UAvbtX1vKczw
NDIQLabLf8ygeOha6ibvvkPDwd/0ug59mHcU+n3gwnpwCOsu0qpATOk5dMlLaJLg
HI2ljitMJ72k2JAqniamjYvcuTsD/BLe9cKDd9mQrSX78BdRF6TrkSDPhxgmB+dl
q5a4/WYuxjwvz1ZaGvYdFMRMaGeBtqPff4wlzXUpKnX1xxzOW7yDt+fiMCNsYsQu
fhY4/mi6/E69SuZG3rBT20BBhQ4F8Vzs3EGyQK817i0SMGs1Ba7Ixh0+0mXbHheu
ohh+yv8JzQyxWdPUYtuYUVpaN5FlayQjSnH1xJGCDZx6MclWDV5+MlX5+laIqng9
hKXAlWtZhkjv7mjblNZs1LKPQl9TnQBPHjQ08wbPucWdOin2aaA8mllTuBblXyha
zX1UjMYGpHeu5lOXmte1jbptDX0cSCWw7niJ70sS/g4hqe1DMNKbk3D7Y0/h8/wD
MikRb5ayvLqMb9TRLnrYHAAGTcHWC5OtU2I45JTycfXvlNlnqvfCJlVh3HhdFxY3
44Ahxhfso5ufASbrD9Kgaux6EwReH9TatCTquhb6d7bNwJbqbD8C+dPj2x1Lzo7f
pHDPe5RT2aO5pVsDFrts8xblXfqb4X2bu7y2+md4aee3OdzOe4mnJTWk6RpBuBTp
N7c7ModQhFVwjRybuTEpakLEhtmaDsmsMdNelEOWjcVfO4XA6KgQ0IQ4ViQWzanZ
IX9q/TMwf23+QuLKVaJiomhBfGI1QuFrkz6HO+Y0ugKvNEDKr0OC7hfjHfsjKrr4
v2ptriJTyecFobwCaw2CXU3t9yGEwTx6S+MgZbjOsuq0arTRxraH+FSRDt8nL/wX
veZlisXBuQFLD8VwukhdMNegPOyN8WO35UAI8zX0NlP+h7o1cKVJQIcwdgH6XVnv
s1w//t5uZLh0Fy7yCpUhO6RbV5UiAkp0PySFtGsKyntnJ3QXZQURUVHadmKqr9ur
ou4tQb7Qk8/EaGCgj4H6e3RyRP4cy0BEIHBAmZB9TECinxXxetBvuOgwdf84Ka3e
EkbDWkDxjNjBcyQu5zVrCOcCr09lPpxyVSjpmOsIFMcL8+gbLRUVnUpfU+oG+7nP
mGuVNV5rh0mWgtjJJKF0BpcIKQCVsyGI7sJ1hXol7kuywRJY8xbQLH1qvt1o9CQb
/yKmlVnwQ7d3YDkKgkqrowhJvswsJpIjchQCODSjaENpVi4w7nUQoAz7I+k3rP8B
JDJTw1TxyM9k59R/cAcYj1Wo/FImwEqBRPBTCWtwUvhPy2TgRsR30EKxhdOYCe6D
uoYtaO6I/BHNffH0HJ/yjccCNuJg3aN3j1RhbGAnz2t1/AIhvB68fO4WOAnw+rPN
ar04DRZySKhcbM/zxTzMQUHBn0tgEjhmom0zUhuGcPNodI/fj5cgpNyY7/Ft5alu
FWGx3cNHlq9/RVegVoDE0BesXRusFo39/a7srKu00Oq6xHG9m5AnA5zazCsf8VHT
v7ZJ3Br9hCy3JGFezNb75aVtrpORAxI666Tg79xMLBZZlWEkH2IvdI4W9AUzYOCf
awbdFJy2Nfju8gmGOO432b+pCGLuWsxx5m1XHNJSLhbBzTxFHS7RspHsxV1GhEay
e4caIa3gc0HLvzTHKGEg9RJDFINOqv9P203Bn/ZciIq9lVmhCoIbdugL9NrtVuPP
3tHjsl+0CAQpBhiAYb1XlHDYipo8IXoW3A5GU1SrwdkBKYodH2XXICWhlj/Pncya
eqd3RtcNLBumw47bmlyu3mc6YfsfKSc1Fm31hYO27sq4vyunMnrb3+w1msWgLEui
u6jGILwgFBebtosCwJL4IWk4FeAm6h874KDsjoct0ytMB9Jl9Ep3OB+gpbjPcyQZ
mbpvqTBXP833JF0IYf5GPHN7UR4U/udAZaJuq3la343sOxn/rK+ABUDlJE/7QKbl
9+Fy3rHvwYU8M51rF+z4EOSHBQjui2xTVPYtirx143nUkm3RpAfyt7ZJOkcF53fa
Kko2xjJJ/U6Z210cZK9VQ38yQ57SCKWrjkeJktc+RRTd8yRaLMg7FZIJDbNQ8Z8a
+4dn96mHwqDsn07K5vFeFTkDC1xYeM8DM+U5s4IInhUD+T50MkuMnyV3kYMRGyPa
3zYLj75t5xLG5Xf5bo2W+UQ8SdLanUZPbTYgoUcU+4bbnGRDP+pmJRsQbfQrLtlz
DNlLN3xyj4a/DSfwKve43uamJBliGc+NvIFCn3yoNixVSGvhQZn65lHX/tYRPyTn
xES91CF/Pp0T3BrVXpua4/mpg7jph+tfB6HZ09OqAV7u3EJoCTIP7ATW/1aaRNZt
x6ZZSykL8Ay9CS7I4htt49vng2SWGlTl14eillgkW2W5PUa7RDW4OcaSB1jKhXDx
nnyjU69b+DfGl+0dD81asT0lClgwfLHRN7d91FAnrbf8gkPzm8fm7DENHb+CAnC2
m1CW3jfj74E6zvRxxzW4jkXiSthV5fMdaVgZEJOyLs2xKxxWGYftE5pbDSolxxX6
dUSkEOEBzofGxpQr2n9eFJLWc1VPxu4HC8fTWZySbzm2NbvWTpQCywydi1cXwxGV
Jndl9PyoD78e0xNdxIpmhj6X1RM5Ot3XNum9umuDY20eh2AIVeNVpzhHAHY5kOnD
hSRXgkiYOvS2NQUooM0pEg04jqdYzko3mtuv7pPOD3DmFjdGBwjiWjWB84w7TxR8
3rV3/deOSzFyJcj7Q7YMo3XYQqpH7SQc9OdbVbmfb+euLdkVjjZ9qCdUNhMv7XHV
jtcHWllSG0s6P5hMe/qsx9R3Ds4jlijGWJwQsi7OhGIQTNT+gAW9ltCBfhzlZzjk
WUAxaE2WAM/BT+fEz2Yx2ieZyfJL46U0LKHoObz5Y+u7aaqq6ssfgFJvlwfren7m
ybJfzxoSBqINR4BtAT60S5yzl1kAJpmJs2k+TLbn4/jcLu7xClic69lgsAtwQ9mV
zehfMMXcbyGk6h2hQ4y0i2Uc6C0dmMFDw+gvaYoGt5jWsKhNGer8i1OVZaqOEuhm
Z3uZrXSHEl+l5odaNwC9kYYNqXlQYH1lmJEzqxNuEuOHhFUIKrM6zHmFNR4iAAgo
TuaU22Ujp7djrY02Yhh7n0OAbzOOG9/MCJccVcTX9lvshD5GzjF8qaBWK2bFO0lt
XC+To5uu/+Y3wwI6G3CkWAUkHAf6eRRlmMA8X9GHMO8KbhUic0fgnMT7S3TRazvs
04LRmbT6Zbg9tQiYtQo0oKyQ0ulX1QU58dlrSUVmNqJwZ7+pzXATo0ie6k/Mjfpt
X74MlE4tB5vigusMfpOXEpE5zgtcKzodAFWua+i0KosVTxwZ0cm98/XF5vR+A08v
94j+KSset3A+IaUJCp5cwZ0b0fRAVvQlf+01uJI3IV+dBQcQJAmbkmuXGM3GfWD5
5LDlfkOvVDYC8Di32ab9KBZWniyNbhC5IlhkAJ1ZuObVsTMI6tl+gfVWxZ7Ut1iz
NzJVMQgcUkxTJNEnln0CBk0bKhfmrn8YeZ7pdpzkR3Xj3TELmjX89MYbsk1EqwMB
0AXQfDkNYowvgRocZ9ppq80jxKs6p3HrzKD6VQ79wrDjJEGyJGgHk97sVZUizee8
Bi9asrJe9y7a/h5hxlEwN8Ql0oBkW6hu7u99ot+x6gKZjalOFH8VyDyIRduDsItO
ud6fWZwEcQk/uJaEyYZHyW2Owy5N2InY/m8Eu5kZH7LvdDjLvJe/zZ/r+gsTZ4rJ
77hvX04pl9wTMQwnRtuamtvtBuyGPNRgFsZh/6nMh6v5Jldi5J5CsDjOjnJvTaXK
QmKSp+2fZ2qqtWYcmmVgjeJWVAwkdSFa70qqYhhNWapkq1P/AV0i9lv44vbVJbi2
THaJ8+VWRA49geMfi/rfDJCXXnFgdGCBFINgf6L+qq+yB25XfKKmJU1mTtCPsVoY
Rlb6p8BUl16ficE7A5p1nsVvfyBiglxozFKw2aJtu+85iUiWEHa4Kh5YOBxlBZ/X
LL4GFDgcgrlmn4AejeVhgRP2+uzw4molMDqSWQLxsCJaUS0MQ5OLZxSh+mJxkZEK
XBWBv2cX0+ObaydL/zW6ckvXzbBQeU/JbT7kYAZt4uQ9mm0Ng77HR43H9BcpyJYF
aMaptiFTnG2iAlvDxlB0c1EkBGm1cawZquV2rdU777VnXdXELUGiLlzwxn2LEdjJ
/v+G0gc05WsE++YpQ1MVk7k6e/HRDhhJGdFcv33+rKrni8RK5hbPai5JMehC7cDi
hzxhn4TnIKMGLCRHLrzUAiW3Xv4qsnChSRwBMWhmnaB2awUu9aXK6iMgpQOplR5B
H1c+A9E0RYZ+eL1nL+jMgQFX+0CAQyeqaR/Cs8e6NYOOsw8wWl/IdXYfI/w87LV+
ssoU9MLNKdpLo8l3wYAdPzvUCFdvXoEgBcqIuEY6O86hHHZeI6k3EZ374PtQe/2g
pqN1RCTu6WBafVT8E1Hui4onctg8MMIVjPz+77huKUbWENwOInTsd8bpWOSyU5IT
/uEGymqWeUtI0GbHSip1O5rpLDR+3gCytP9IFYVLMkUK83hwc5Fk41xntr8ji0BC
EU4c4vMcyM6Gducy7rpAxV3CWvEdkydgt2mrnHZf89KLyHYVceDZDvMj/1YAklEP
bVRSSCq/1DPX2iKbEWQRigr1tgJSG59og2GUiImWIi+SB6Xp/Gy9yO1zuoT3MRfo
u2UXvXJ87bmKNhCWEBtLcMlP4WznZJr2tXycDcRWq/SlM5rkHM5686ei4ZHZyOpH
MkStaFqDDOg3l2csnDeRBOUNRTxK4oaylcSPo6YdkwZBLy8YsqQc8THnRMz3+btN
tleuHGHANlWAQAFzYT9ai82l+O+QfUdDFLkx7CEJdk6xa5wBoMhfKzOIiEbjRMD1
GXKTk3cUJeb1SRRhIad0lO/JUcTD3ILpIBtpngSj0PSSyFYZ0GiWydoO5o8Xb5KW
bJsH9uH6C6SUSbzTj4ob2vtDhZv2vtCJVPv7L+Yr49uNIdAw0e6CGOzDHP2nJzBw
EOZtYbP3wygcIuL1oWpnXVu2vcd+tcsLzWsVoE5bjTTfAErlhSwDSciTFBSe3SqE
TzCmcfzWEVYO9Fr76374/yhLtm7i7PMYuwYLxRznhyDhLqctl3EywXdHE9f8l/QV
zjYyhi8/x4hL2W9dFcRfYB9VLzGnCLabdLepdLXYvtlX3shxk2PEIlK0rTdIk5cG
AG/wXUXilqeCNLOa5EOS/Gxco5Ts4Qf1XmBF6YgL2o5CyaGQ5YfYM7WxQiUUesJS
MrT7YYCxHV/C1Qx7zSASzqj8kHZuR98la744jXHsXc/sNXEDH43G3qiM1YXEZScx
sOfdRXsOhmUCMAXxjxydmw70rHfYjY8ih7OZpi67qvBO6dZoRbwypXn+KNvXv1A7
+0XH9vL4IwBdNOA3xf8DiuWr63sIJi0+NXv2TPUMaMZmHT7vJzJWYSLdRRU9Q0z9
OQCy7vdYeyNViNbP+U22usSZCtULNMs8ow1M1n2hE+iDJ4+0wXiLeMdoVPNc27Yk
k0HMjZX8ynJQg4g3vk3fx+ThfsBm8kNsHxgZNUHUVt3V6uDro3PyuGR5LPSo7RCX
p0z4txSWXPF6elYci030OLAuILWa+ht5wEc1aNKLt/vWUSQrSjSDVL4jdLScZ2n4
+8FfJJQuyMPoaf+vSLrslJXgSA/O5UK3iDUkdAOhDcWJHhJoZHC3Shsy+dJwyX9Y
GMZgboIfXkr+DtbVtKvuJZk4oirUN9tevc62QjQOIGGUoLjM85dfn7gcnbPouKQu
qgiAbsz6f4DfzTx1MGq/3SQvK1NvExhW+1efIjlZrGuSjdmB/+vKksFb+Q2aTCMb
SDvDa0hAijCA6evhGqMiTUNNvyurV/plm6O4T5Dne9zpI2D4KzM3NDg4twVQ7U7F
gjXx65Vx5GOlNPTvdyR5ikZdXbYd6dKHcXqY+ZBclaDk3mkoWW1U972I//oe4OtP
F9AU2Uo4naABTPAa1TdWdyl/hiItI0lKvzps5yxHKOU1cfW+ZAaIHOO2TTEK/C48
dOZgfWBSjb/vpGKUwaOeqKY13qL5/ObGKKbjgwC6cEs5CEZ+vyswQRaGlzMe8R7U
6nsnAXZuP2QHE4kkvoDyojUBOFrWI/3zHKcSdv9soyWpYSWbGtl9ZTNgDnzpy4Q3
Vu2PkcvYI/bb9OxM8VwRzQlGxITsvht7ILk/1pWQFIIKnoQ1DzH6SxoWL7TQnj/e
SQ1L26U2RQVJahzBpjOJsU8GVs4wQOfTj2uW8AvvsJ2wl59pfkIEvBISteK8k0NQ
DpBj8gUL6u8Lrop3qzvuNDhNZnbJgBe0CWqZCnZiortHf7XyouzGXooSMXG8IeY2
5lSPjQ1YtPycqX5l965basnQdTR+GxYYt7u9XS+AqALnQLAu0JHmZp++DGEVpeIR
0acOBCGRqsgUFxbS0FIE3VlCdoknySnXtbeuWuov3ulHS5DilF5HXzjLGTCF+2O/
hQWBvyoyup9fQ0ztoOw5pjTw7HvZ1oQChL1opXgZLrcvu5mXO2eiCQmqvo/Lg3ta
sqhgh4h0WDdixw8XMa/4xobROzGDsc2thhZ170qlGE8y+35t2c05+i3MftsYr1oC
Or+igEbWkEZ45glgytx6L98qJ3OSmJ0A51KVX7W+/jPzenFbagHVIdgAeFXikQXu
jNBHtQlrTWXJzMahVoH6kJ33/Uy72uKokeaW216ydy/vyw5JrS/2G8IkPGQRlGKr
/5wTiNC2CEDp46j9aAOJCg1CMhpqGwikYZvBUdI4wTKy5dr9CI8eXI5x5MzxX+dB
ZszUNZNfoDSMk9ydAW96IrcPczdmoJTT6bQvhnzslLkfu9M4EHM8/IFzzeVI3Msi
9lW8j6qNN9fBYTJziQQLrOPWCv+wFZCeyjLdYwkvTt2LHJ14EhhTt+wk7MNIOvTO
zFY/t0xUi+h69RD5vkfNxqUfcgUrrIriCfAN/7ZfMqYYkwCACgPERHx7k05cVI53
SvzVSQsFFW8rvN9Jxm+CH2iBtGMF/5bYM4pivawvxwNT+RoIUj+O5zVBvOW3OVMj
KLi93JS/BRbXYGFFv+9vhxMoyMtO4DsWMQiFvLayzxa25weoaBmPsEcuJSvhT/3a
Chj7ls2Anx/4YRvU9QfMYXzklV7cGf6ZS6GGOshXbiOM6C1Mfv4UlQ5eaYGdvmGf
8zxaewtWz1Pjqg6M8CMAzmNswiTzE+5wYtG8QU0zXryZ0FeLe9YzreB05htA2uS9
E1AHg9Y0B5v1TkLpmPNCq+shqpBDkTPwvE1vmGffAb2faRyd9uV7um3dfIBqFofJ
e1wo8e3T5BsHdFhhC3pUb/VnVxl3xP4BlIV+9aXvkT9FwmRYH3xp2JYqI/h5I8Sf
a8lNo50K3AYmk3qrzoTDNtEGy1HQulaNySW+0lT401tlmQfw9mUO1DUqWG1A+Imy
JkWipNoHOJQIW3RImxDoCtACKMcsFINURTI5xo0CLzEAATSHdggU7M+fC+WsFv6c
A42SVQBhmmS6xEyh+VKQ+MqNtYwQWHRCs/zXntmndggkhj/16/DGdKjq4M7qg/QZ
xCBIaz66ZBgbfgR4Bq2JVRgAIeWZ6n2vE/hBRbwo8saI/XN5NyI04ehyu+rqVnYG
YUCD0mtf5DOpzeXtDY17un+TMjaKbygp0rYj/KEJWZ4ocGUl3r2RdkfwwRqyjoMb
tHI1DOic7ugOEOd9n8+81zayWVUsk43FUxFbnpwM1jCamHmpGYFXQbr+svV2/CZv
S9A3lmPugouSW+ok4xUgVp6QQ/T1q91ujpRUfJ9BZDKp0o6H+qjiqdGDBAn9IpRI
uPuzhLUjyXG0Iizx93M4yvlhEy+hST9Q0Vsi6FeBf6Et1eLjAPw7Hp+6B+Mgdkiw
ZuQSK++C5wbaog6F0PwaiHJBTUbx92LhXYf4fBRdwRTvIMiZqv3dGWTn0GbjGLjS
TPEBRNlJpgtoL1fNjgUGK+a8c42cdERWpVLn7wI5AnZL+NCPedFteYdnREghLbU3
6qjlwgivTmraERu4n4OxdH+D7lRnDUdWNXHetw4s0MthzyblHLOrfS7Hm/GPhTWL
y94bCqc/QMjKLHxSdz46Qvt3nbV2ctspuMNk6d0C2tpVFapAFm1pmIhW7Rf/Q01v
ya6j9VJwmzk+DriHcBH47f0CAI1mwZqLqMwWYMqz8/tmWbyzH/32I1KKKbWN+DXX
3+iDRJNgFJbpGcq++ltAO/hmaf/BBqVA/HVPJpcP748OezO3KRB8nUCWjBdQdtrZ
ez0kpn2URUdDXah05lePhagQRpzqhrh4rJTyWt9UCVUa83Ti5mIOf5DBeFNCttJT
NjOqHPaQTKT/jZai8P1TPaXxc9ZtuuuMtMeZOzrgzNskblilqE1Z2X6QGygyvPaO
d6op6rDunPOkwm3kHV0MgiLo0CQirV2vM/ccqsz6tPmQgdYIU5cXXWpPrg1XOkrn
lBnAmpUemcdWEZfxSetOR5ZZmVp6iAjIi8poEucf5Q1ClUhbOHj1mCIarWC6UHgS
1qBbCWFz4yHjkDGhyVW/UYyR5xzM8fldTuoMuRrduQN7wqVwZ2M2VB7fLWvX9ObW
ZEur44dF/SlNf6CufJlCgTMjrJyca98ICm1TB98RBCaswSdRAmzZZpvRN2/gyRA8
PPolu/bqNCCT7XwwVPUn9XTNFbt3fvrkbIceQCRr70tY/j8acEG+dOHerHu+nmNB
bJD27EyVs3iIUTLQfmNdwQBAorB9ugC2So8Z4Bifn3Y20rLCJLXQL8qXa3LL8nZy
EDvCIJelwjgoR+FKM6G/jp9WzKBcVYhrNkhjpCQ+v1XxKAioSYzDA9VD9xnzBFo4
7pOWzk5Q25lMx6O6pXh++nZTOBaDn6TkMgaT6HWNv3eY99QhvGjUzMWBIpNaX7/v
+pxNKdwSWgCVk3jVA8VO7TOUcqekX0d67b8ml3jYteR/xj9aBQxN/gcrn+cVRC3I
mUcub+0QvR8Dg9syiieKAenGSaAS4tAliD7Hj6Kv9lw0pGmfmqhVx9l9QQwjXRS2
MOrgbMiguXYvCvLAO40xu6f5XLOFSsFij6YkyylcW0SX5mvdNLI2nDy/TVHdYB6q
ZU0c3qOZpXu+0c2tGEKcUNpXnmLWyzCWDBobkSiZOoD22pWsT4Q/ZdsUZxGCgJTY
AQeXBUjdoI2yep3uDTfY58QcGGJjfY0hdA20F0xzWRW9daPCm4pxkHzQSFBq6PKB
G2r2Ycpu+pPVbxxxYi29Iw6sCkCj6kgQaBiSIE90z+nJvHpi8GVKmVhdBuUZF952
czpJJl031falE/91w5niRU/fVBB4dKopKHYzReq6sVkmQmBm5vSYGIccMXO36k0R
tUjUwc2d4wq3dSRhm0Ht9k36OmFSdpTfhvjfooLdROGESrdnDc9qbffC1VGqUZvn
eX5eLDwkY5I63d5fpZWc2v6s7WujeJpWFNZ85AL57qafZI/D6/XBPJLPnED2W2WF
e/eplbfnoHo51fq7rGsCGiBUGybNdS7Jcc8ZiwbgXBEf6hDTMH5mC0Dm1Ggem1bA
RW6vxyadwf2i1c7qOuJgEDMwtJNC/y2vYJ0ENDXyOjdOmtDHNsGHJnOo7PxTPg0c
HFESwAmzMxmDYandpPtJNCWRslOI6VXG8Te5hWCOjjgfafmHuVc4I/lob8P7vV0K
V9MZ5ET71Tl7mITLj3Ypc9b6xMDox/kbvvlxBiCMlTKfJ8SWw/a0LrMnsxisqx1m
EAWTW7wYUz4UcAdJG1wbyR/3fw8q7pTVcfU1fw7YIgkFrKz9TtJYi3c4c8m8k496
iAMaSZ6zO3BFsXZ+8ASH7Eb9QYqGayeCtR8SgrLQX6765/YwdCYjFFBFoaYZv9K6
P5G7dUsFKm31v7u3gOboFd8vbty8jzSyqpnyerrHcdFcMiUUmRTHeUO3EAz02Ynd
YItoGB6KhcrxkDK1S+JGIB/WUCAv6PkR/9OVUD5/aWchIPci3bVQIPW5zLhRsMQM
FvbuZomQ833BWN2xoUvwdDEFgpKvwRLb8HC1r5qu2CECR7oR0r2PAntTnbA886ds
d1t8la6ao2fdvJDExcAFEykAUMPuJUB30ccuYOhCqRd84y7PP9fEx0sqXitt5MC+
QLMDnPfymWiAr0y4gm7qH+0BP0PoUlj5OuGPHAx9rzYHbnxrLXZFOy8kHzAIUl2l
fMSPyvcsPyGZ4W5ImGH9EKbE8qxIMO8hPZRM7VK8D5YVmKaTItXXoxuLghOxU2uO
ny6qwJhgiBAWlXYUvJwMajaSbxCixNLtT8dJuYHfCTM9ukrZqKuZXc2tZ6D0bidC
7hwE6wVi+sfcIH9ASbFmvdyA3n6/75CSfmkr5oFivBK8y5ofXxvbmJR1mnbmeiEX
lLq0dLeyxsx/Afe6KZqYxMqutVgXojns/dJyNBG/DDaVBdiKdUL4I6VT0AablUug
VWNYprREg89vOYKHhZx2w3/YnAxGqUAvSAcP/VqGAbur0eMm6PGe0hFSeYu1HWLF
7p67CYVMikkKIvOt8S1AbHStsZxe9XABR7CktrnLO/qUs7RKZrEsylwjCrq3Gm+G
W2Udlb4uqM/y8ICwwrAHMPfbDQdEwdCDDCkx/3ub+w21vIxjzjI/UsmDt8i7tnpy
0Rn3gvtaVxse0UeqXrMDj3GivNxUSCzT6PJ9xqGE0P4DWLqIhq5WAlnfgFRq473F
0g84jgNbMmfVrqAee0siJ/7xemOpng3iM8YBC8++j/ksUO9oXG+mMSZ2MyeO5D63
MuJL2j4BGa2gD72eIlD97K9xXhrIhqoZOirJybJIWSnr5/BMpmcZEsm4+65nc7EU
ZhOM5MLgY1NlkEifsodFtpKC1UYOSlTWQqA92+nUZz77JOG0kaqiec7iIHv0s7OK
9NaBhGWMH5VzgKrqYLll5l7W3mtTHT3sWyXN0dmvrhoMBrBoHU4RHAjCLLao6YLk
/9PykLkb8oHcmAMJmS4eOdu5uXN6KfCExH+GbLFSL2nQ0+lK5G//kiepNnjGZ/+G
+WK6lcL7b1FbLavGlJ7zsuh0btJMI3503lTuJDu1u1q49/mvOMnSHg4D4Ft4VpKp
er/mFM/a1T/T3QYdtHXTEizbdcoFCFRv/IB4ALppWsdrE+Go/kDqp/U73dfF0wvb
H9f4GmNmAwTu9sk5cZGrntNzh0aTrSWH/z+rgPch82sUY725gOzRPHV5Pwc0bb2g
ORGHDXuyNbU8ThHxNyOQt+RKugr47mspMy5/g6sz5U8kqkkjwUurEU7behkRFbpg
QS3GvQRhpjNYG5uh32jvvMe4eHS/sF7j2af/eTdbWNZjHXxgkPrJ1n08VSow5LjA
Ho0GL80kFGYcRQ587N2ZtwE4e65iBDxRZhlsWwj4fMnmvRdL6Z54/lEVLKuUWKQn
sHvYEjOtRWXejY+pT2aGE/9RnboKjhqbYlXEorXXTJvlCdL9rr6wWJT10yeGwzmV
Urw01eAhLIQNK+2sZyyl39bwcjAhH0gRPrW8P4ZxsqIYVi171Jj6qgBiK23RAWoU
m2uNFvhjJt+4lCMyjGu7nM8J1gPkIxKXLnz/DwY8qHZ2WFqVMX9Jlt3g3BmpqS6+
jr9J//T5FLyH++wSI7hiJYKRb05Qa70OU7EhbN2ArV4jpEIJpRP8Ak/J/z1sUrZx
gMzg8J+HcJRTfWReLwjJMl9DsxLokkoa+9xuKDehqdA86i0i1rG7MHSXClc6A0Nl
BN3EMybf5xyShr4bFSGUoqSXrcudQd4uq9llJ9cXDhMps6Ax6vwzYBEiW6+7ep4b
FHbGdPadxm5u2QXNBc2lsJ6eZcLANhvyAJuKpwIHkvt7JSO2rld/mVfHXD7PsmJw
0pwaAPXQ8AlDyXFQ06a7gu/7SSs7F9D2aiaEzCcsdCDUnAPaKlzsRdUUG9j3EgRS
SU/FndClcme67cdB6QSVZY59hJFz9Ot1Jka9hhuJ8wTKDoJWzuzUjhKADCM6SDdZ
XO2RTz7ebLNZTT9/0WyyXar4rAk9/x6rhBWtEvnMzC6skxlGjpsor+EbAlulQNoJ
aY7O5NYwjOK1UEKtD/mGJ+XYbAyHpY4YjDbP1zY/fmdM1aSupxzYrERQxG5HDGVt
RHVRRBr3PTjcZSh3cqLKaxZydV1C16uh2pzvqbq+gHuJoA6B+5bZkaA9wry10g/P
j8fwsvhGusNjgj5RuFXsZAzBftXFB96w1+PVUzsVMeI2hYy6QgJz7caf4nr0JusV
ysdqI8PzzMzxqFwNG0nOy5BC9J+fc/Yav9wJs863TWAvMXQBVKwhxNTYaf6wl32N
YQHAlPlJE75jcD1hZSNpRf9tsB3nA5h+F0LHLttL8MnKf/yVEUsg86D1GJCowzEX
odLkjYkhjeYTsdnwA7JGV5lqSgfayMJPd/HdgqZU0Qr6dJGpCz3Ao7wyv91jcwVk
D+fLv4UxgOL2O2cWce98RGnfxsfviyXrjTqh9/49P42eVRmQmnMLu1EXyYL9CACM
fKB7QcMvLw2yHYz10rztubpmtwK/Elr1aMN8b4JheCZp6TGPFh57SGRoiG5oah6H
FHJsOpqtYUZinE+3IBvfXbmqyssFErPc6W8F6AwOX5UH8ylKh/3jXtESuCAHIzFs
CsvZ1RAvL7EvC7juCMKdDTLup2WXpflOLWXhoojD/qFUw63ptyEoVTVDNtVXuDNC
ZzXTEJlKaDy2RZRV7McRqt9yvtbOELKGLWW2wHAReIM4OhkIiib35AgGrJGWw7oR
p09Aa853rv6mwHVdeFroQozjTKfmCi8ob61s03n5peuuLNZ09I9tFd1B8Rd+jjEp
+k+IO90GvsDeudNgubBxGALr+8meZyHWTfQj0ZizFrmX2p9P5z1mv0qYguwxjrEp
CXUC17NUeJQcaH4JVK05zfXjG1Sp6ntiONL19dUKPm8xz00Q1kuYSp4rZ9s9sYR+
N/WDAz53XyAMq9Pe4Jt9bxW0DImvnTZZeRT6Ct/in+jj7Rrewr1aSyLoDf2Db+wK
7BkTbINUNQw46feR160wvlXQkIVCd7WjMFVnhO+AYh898UATb+wnO5YnOlZEOUKR
VMcFaw8HmGRVhp5xFYLqrAwOF87mw88HiFxwGKK1p7oE6CssgpHV3ov1Y/b85S2R
pbn1ZF7Uew+1TwPHCPGeLKG1ojC0HZTt/KRiNo7ZmqrlK2055TT1uJAk7MySqrbM
fSk/6F+CxqiYDxgCYfiY8kWy8SOhpHGsO/pXX8Tz9I5dBY5kgtbaTsIlnngMIRMc
Dg3Ya0n5nQRz/9aS1cSUYYj3KXYCwkCzI41s2l9V2+voVV9V1UeYmtEHwRhn3ja9
DqGPZ6xT1BIWEh8+04ixAv0i2b0HZENXyTkTHrA4ZaSBfN/n65skaaeH0EVtXQib
gliyHVzM9C8/+4FsctXgF48uopghDJhT84KjwrH8+1hebw7P1LLTB+zxPuCgIPwF
xeTitpsk18wZ20nQPdpOacnpr8NIM1oYIyqUDiZ3NPYiYlTgXCK7kDm7dLBYML47
mIyIukFRRcNJcQfaWPK6cYivG9zLRfErA0i1XGaXj86mDsvaE9d+nxmjXvz1L8Iz
jnZKaeK25FlMNlYBwJG8xS1iu4TAnv7qJwXhr4eWuG+YfJuqd2LJ3vERIWSHwpOo
qcxAuk+wP7uF+qws/weW/6Ycvyj1D1cus2xVtANZpqk93M7ppRB/tls6hB0fwxdM
EQ/rXSjDT16+rJ4YhJ1eYlU50sQ/W9+H6gbR0p1YhXnoUImB+i4voduT0xVuPPsZ
You2Zk5MBMvJdLmJQJyy7Umy7Ga3OugzuZMMORxCFPl0d0n9/V8DeQEM3+a+Yw08
zjZnxEXUYB7jdY5c7JzfidC3P3+FcEt9Q6VQK77AMBIIRhO0ItFxtF1hvf8W7hQK
wi+MXTZZIBw+sZvSHR8tTYiDyZlht23/nGtSY0t15nOG1pEyvkKBpzYdF7MjxRcC
P0Bs3SrZU7mSBoKJJxbE37mdhX7Cx1G4GeG5K+6LYKnNBGE9TgwmnH7FFKiuD8ZZ
Fq3/7PgYoTbhSQwo0cyJ8sh3BUy1C9/pk8HGd01jMFZFKw3gWBw07tEkjW/arCGD
X6xIQ2tVTg1sQZ+uYMTV/9guLvHHnDuDM9UgcOcM/EYkGBQhHiEIAuXs8WF9pcvm
AbgKgW/kGoyVLR1oUfsjMubAyOjbmVqK7lgZ5zSyUo/RVVw+rjNwP2fSP6xLZ6Tx
ERJBOSIMXDkvYU991gGbjfCQy5dc0Dds26FIvuLgJyJza37D+nFO3VJUrqkOGKff
0D8eT0MKj21s1cfkeIGm097ZkmqYElI9J1ARbjj+ggPPO+g8RYIFzXtdUHMPhBqQ
UgPBe1ajbiB01gZCxfWTSpVR8jKiXeQyA3KcumrdNnyhlb5/W3fNpq8w8QWkxrcR
Xf5POHA/+JDagrgdxZ/7fWWNo6hRbNPTiB2AB2rS+Xw6u1O1B3ZRl74RnVMavhGr
lU2dTg+tM6/y/N3HzETpPI4PyeO8gDWtMBIqXaA5EXcyPMUuI+CdDu5Ijb1KEyOI
JCI5Fuo4WbyjOh7+Vp1a+/5gpw4Rbxt/U1mqmI5p0twY4RJLqra6uySbivEhJW7U
gasPDw66nkx6lWH0dUiHanCwtfRC6VVc0AsSjtgzgvTI5JG1qB/FtxYdQKT5lZqV
xrv75kmAsbGA73FHsOckwNnpZvcPH+1iI9RW+s1bv/IFUXg/1eFq+E4etTJo+iZK
JQq3Y7AdmtvuyTc9oDjndHplzvAlh2dVEhdRQmv53jzgTOizaa6DsorkrxmQ1QLt
UOZxWYxqdR0Z2rCRwpvzzuwKYWbt+hydzdvUGTl3i0dtMBin39FrxsAwJ1PF4GOB
ERnzKmfjBRt/rs+eh7oIjhwk4gTcESo0j/ZBVGK/p+j8vgyDn+HZMzuJalfuJnUy
VE6PB1kh/BERLwba8rI5fqAlZa8Y6/xorC1MhCZ+f97S7IoxY6kpvURgkO3uT7VR
W8efTuysmVpa/2aA/wJqztdUT0oTMYlGXUa20eFD756NoHmoHcUIG2X2yVIkEjd5
bUu9mvcJxijlA4ukwEqT09IU6QaXDGRbqXX0IAyp+JLOb2C32+P42Ek4gNrReHf/
9I+lEEOtpMrgIDJO6whcHWRMInblZqA3kPvcsSrzrAnnXoHAhwjin5mcqsZZB1y4
3znjkKvhnCuehEvY3ZEtC6NDt3bHlCXohmcahOOrZKzawi6tayhmOKvRCVWec/um
gvsIVFVlPljSeCr4cHaEBPViXFh7WPBkmPotX1aoKnTugrs62i8AIj5dMAY/j2os
dn6YL4OKgmSjdNmFU3CgCNpyHWV6IDdveMiDxEMcXGiiPoFZWP0ccnHy9BBVlx2k
0xXCVe6ohQFP0T+at+DFnx7VYxwZKQKZO9GESr5yAPBEUegm4NzW2NNC2jezohds
FxAWLaGZO68/gdI0qNRb3p2ovnZjcG2q4zC+u6Y7yU+gKp9O7mKbcVj9ylZNXN5M
EoPHk6znleHlo8rZ5S3tvL9HGnPuDNFUfJq7IZVpGaIXuEpr+MJOt+nCcvTJq2uH
FAq/kmSPTpFEkIyaCypR0iDLOXH2nO5nx/CHO7KblEcJXe9RprLbkxoymeur8KXi
SfvgNDa86X+1UrlMO/RPPZ98/LAC/SrYAxJnZxE9doQBjR6OnraNWfopFTRZA9VQ
bIrJIKmHvGEbRZd2vDbQgpKt32pmNd/zwttlcQLfdD9GJoetVw1eHzCuVo1e72KE
xe4LLTnTr+sBw7eDbYREh+gg4ujh8ZhrPR9ozvspsgoeM0PKL34/UHg64PgEptAY
a2MyuaIUDDEIs1EWR47EaPvyD/VF1kpz1TgmLBh6zhw6rJpFiBOu+wv4a5016G6e
fz4i3cf1pdUSyhXp4tXUQCyXXtOYzpfTEc42orQDhcDbaLBwSTIS5qABnTrmgp/E
lZymBL5TbHF/1Y7pI4KO9qd96aDD9dO5JnujEv8Eb33wQ7gEveaj8zloQL76L8jZ
2P8yiHpN/f4d8ANhdkwnb2Apdom4GZkU8RJEjGFbQHlyx+xlcOnKTMzZ1lV3PRl9
uSciftHVP+TYwEsB4WZ4ui+a0yFzE/vEjy+rc1oo4CxA1Kkdktw4epKM0GtqGMBC
EnoBSVyhID9+mfm8azjoIPYdUFnDVjyjOxf0uUx7Lm5536zdUEMymqDhYpLUj2NV
O6JN5safld35Fw7eXaXfZk1aYg63ZJrcqiEa9Zhy8U2aPpgIt3tKcz6hUjUZY6hX
O3XA2nzO4RRHEbQZVeN1ndiRcCLX6QAmKuwgOPp+k6B7vvxjH3iW3U/IQpuNezPC
rt1cLEqeI/jttLE6uO78vVDga83kOB/7wLVXodsFoDXtSS3WMmH7gIfNNjlpgU4/
FToVlqELO9T+xajL1MSTHrC3dprZAJQNl/L0aKsYEwTMaiNZZ6kd1yBEW1KYofNm
DL5Z3xHI9cYxiKSpg4qS+cTpOFVfACvFrMkWm93zFC09DsgRRXBCJ0Wd/J20lzgg
V9w3B6+wf3YcXG7kjz7sKp6xk+dbiBSKwc76P5f3Vu7nli04ZRtdwb8Y6JIGbddk
iJqHeVl5Si2bxk1EYbTwwTIbqGd4Z5DQajxD93kEZYAeZBuNdDs1CbBM/0h5k+QX
MlMcVWVnPXPecKl0tV1JiuieJJyPHx/s71UTSdG8RHH2rVZBUKI996BX9psUW7mh
xEs01bo4Z2UodtJmdEIz5AXyGyXdkxZlVyxxlcYXWwuEROCIV/w6P1OJbNbiorod
aspGMPRSm1SgZQanN7bkeDIkIEiENk8nnS90UKLCH/hfdt+OPWE4qIvzMMZa6XnS
VDXp8ACPWf7nXyJPt79KyFaAeS2FWbSO9yOc/RMmoVtbVdk8SjJKwrXskO84aLl+
jjxcr1PxCgxX5hX7kHMNzGsJjs+Ybv4tVGMDEPFkS6E16W8hbcyOn+mJMN3bseaO
CJyhHyfkaRiJ4za0ISQDg/s7Isl++gxV7FHsNF8RcuCvqBkaHL1oOTRHkm+XV0B/
zRQTZbruzjPo6XVp5NJo98zlLru5xo+0suYJKM1lcHqQwwYvt+qGca5NF+UVCMU6
UElr2R01hoPQ03GW9d4vZCz14JEo8v9hGs/kR7emSYozKroFMpEnepRlpKGuUUtL
YwxWgWIexlVBPXtJYsxWaThui08dUZ+OuM6kk2t7Puj+5/WJsluYs9wYRAZ290a/
Vsk/b92Ydp69FP+mR9kRD+tZuj6OiUWh7/hO6psj7w3GC7H6onjXJ8vVNFPTekzR
G/F0PEL/5w3HynBt/qNT++GpwCezYoxGfBG/LzPYAh7YSIPT6gvSZsJXJkkozQYo
qLUEZlK6E3UvYjelXg/LQattOhnYRo8JAHHHdkuI8qyg81gogR50TOpAWQPVgfWr
mv/WenB5tzqRaWLkLnSctUqvkigyj4Af05d1syzLBaIXN/oTC6OnMBUcORYljrR6
PA38r5fUDzWqxvQvl2YCxzdFveBpbQ405kTPgEwn2FX+L/9LJ6oaFa8S51sXOk22
XQh9gg0lfivox8WVuKkygqgu23xPJwvbSa/nRn+rdxLeNg77iBorTryjIoNLCIcZ
WPkE/GWiAIqna/VHhssw4VNJc8388Vh8/FYQufnVU3IfbHxkhdz/vgnbrbzidTHX
w79Q6s9kGV9358+RMBE89LWi9ELqD2ZP8vy2+y89sS6yNp6i8LRzvRo7q9sF3Zpv
nFYVxLXOAJRiXBIsIEhx1KHG3IFQwteksZEHKhsRKlroJeQubRpDnFckKJrpbpI1
gs80ZazsyBETYzRo7lpaP+4dGy4BgwEy0r+mh8M33Y53Z2uVVj4j7RnYhn0+gSLY
b/mNOqySCr57d2y2XY/tjXi2yerJ1Zy6IUGkllDjoqmwko+0ECsSOFfXgr2h5tQk
Y9rXC+EkMa0Hy7NkZ/0f+wdvtSXozJ0c1fwvm04fWMVP/mQUbdUxXQG4MAWjeu+M
4S9cvC5L00kh8i6ijKAECGxKFwe2bgqpOvduPBqsAXdyVHHV6naIYrCzafBPI39x
EaDaGlYNHj9rFKl6cDkmPwRQZgs02h047PM0rqmRAimZxMp/tlqpmRm6BNRinZaK
U2eBhzxUOzUtjq4C/Jr8jplrJzFl7xjDv8/ADqrPFu2Iz6fF7dvGYcymw8Cgl+oB
QhGaAidtoZFmNs8iYefIkwXkG1U/xjyaB0RbK5V1LZMRjizZwvF4QN5i3yfJOehQ
6s+L4fLgsI62EADUzVBEhFIkP3mX1mENmjVI4M8eaci6V02xEphvWjaOW/gXw5ZE
v9CqEs0r+M0mn6ANkLyJ1hv/3Q7k1Qls/fiy5kriUlJwe7EU7wkBN3Ix4TthLAXm
CFahbF8kzdcPbDlPCmjmf2kTYknThgE/OGgBNrycxg9IYfXaQr+shcM9YSTj5zIL
hSLB77sabnuy4IBmQge+tnp/LtIpK28YTDvxasic+snZKk215XHSkdn8dbN7Xgby
c7h68I23PyKdpAFk0s1CAqlh1BoeOMByMwVblEt+nU/7wXAOQPV7FRdKjGI5EJQb
ujubiTF2hSsigesmrjHhLq2X5fE0/YlqalDbRFHPgd/Pr+e+53lNVjrRWCclnFHB
vhXCApO9nSk2KSOnAHWImcWM6JAmRjuBAaoHf7HfZlRT1BQYRdLQtb3ntel73gog
wI1/VL/uHh5/L4XgEqBqvFHhWmBtpbVcYLivRlp4d7LkSjH/km+A3Agu0MKw3++q
FG+YqXSMD3vT5wKy9StPgdZw5ogDKY4R+h/ZRzgGpGEBnJMlT9WTO9Z+J/jsKffU
kuVet/lg+2/YMO5lBdj+Qs6HT8r7k/USrbRINViXx1TKbo84MJGD9nXehufBRGPw
X47Wrb5FXk5EsTmDE3ngBQXCPTeEaSaKsnNSwiz666bQ5FQJblKAQNC1vmb1XtJu
MSHNWhD3xf/kHjx0KyiT9kuC1XocVSAj04RwVNfSk9i8csSsF5OY7hxXGAEYPb99
zTM2Z+pUk8mZqzq2ziIjjFfNBJ5AjMzmRDA8YeGnrszPcizaNWzFHEBuwmfqxy4S
Yhu15C72ZGTR0eEXYKliFyin68ylJtP/FW/TPtdXw5tzpufz7IMoW8OgrkJE2Pio
af11NzQq6r2ad60SoqM5DRj5FdRmHRGYzY7coyRGTMn+oxJIBdObNadmvxCpA57T
uSxm881oK2Fgc8c9gpi9ff/KIZ/tEJAH653f1/7/PCYRc3mYk8FBC5AjnzbKX2NQ
G6UsuzWQSYUMZQO7Yba2QsZwGGlsDJW0BnhQ0m7WelOZgRTl0UXdzhHmSwly9IFf
wlauFAji3A63Oi5hcptBMd+61jic/3qF6OlA52mIss9iNuuV8U1IITtsjezimu7d
zTGpg9psKnITTFTnhcwoGtwcvODFW88FGSWVPV6WD/JMJyVKRqbG0lqe+cZxxzoN
LEREnvDN+I6vHIMa1os9Dp72GEPXDp0RN6KbRZw+9HXzPdJgF1cFbrqXCcAsy9lf
3OfRHIzsLLoua32B9UMXR6vUoijEs9xvVyI9pK21DWJRuryc8BcPN6LPla8UIk7s
qPPGNfwRVKMp4A+oGzmrVoSVMLdFVdLX69LcTCAPh51w5IltjeNyTi+Samf5PCRc
0BQbs2VZ3inWJHfJsRJ9pXEcvvd5BYkKJmQPCAH0Leg9AJekZgkyAgYPpuLFzNXy
6Y2Hq//HAh7vfTx90a+dvXuZ2Y1hC1Az3MTEPu4mapVGeUm3IA7UWZsMaObI3KwP
lvxeRsE5FrqaFXi8uwvvMtasxz8S3/JzbM1NDPbrDLGGElNOQNeiWeUIaS+/aGek
1Va0sEFlRvZ2AgI+pYo/O8unE8pIN1qlknYNI00uIKiuM6be2wC0dg3dMIo6rB3R
jK2h5jPSWO+UYiY3op2WxlkhSHDcitPWZ0XJvw3OgH69kuhNUnOy1fcoVrspr+1k
mVdEcl0LkSKnD/uNHb4nRHPy5XCk+y0MGOKPh4NxnBs52Xf3NWVCJGXKryyahpKy
PGA3l87Y3GajR8EQdrkBf40OK7j5uFVTXkleL6lsDv02NyTKcmzO48Zj/sbLL386
i748aDF+89ubI7AU6zpsrMKstJ/mZS1pegRiqXHq+b9m+7TSdcczHdG4elBc+0Em
iWlfNdcN0XBLgWWiPY/ydNFlq8S6Io2AqX7Qo39XhLuwB9VHDcP9BbVU0NUxc8du
N/n6ze09s0/bYUZ6JqPebBX6RGkFNxNzJwSkAOoSeQMW2B/eBSKgs61XcQQy7Zni
r+4OPDnpILHf0FfCT5l8SI8zIeiHf+GjSghiJf5NsbgUNVPY/x1Q13KBpfIUXwxH
JYyVJBSQVtwNQmH/dINTiCT1egNwB8xORJPB/33z3UCe5kev20Y+QfUZzJRhK9gO
528AiX7TwfrlfP1XxjO57ozHkqX45FJ5zZprTD5Q7W4kiih3BUdB0KDY2ofSRSh7
CFIqePoAS2AAA59tSeXgoUBdnFUgkJGcu8lJXNFhMC83ciFD+vTt9OxJPdh9bIc4
siUOLMj1Agisd1bULbHdZwQ7+igqQpnHMPaRSAwacBXUb7jxeLb8a+uQrljJnwjq
WEfbkgXPTDb35sWsIzVGkC1renYt1Qgs0JLEgb1scuEyU46lNcQRefCbTVmsMY/L
VoHAg7HnKOwK6SMZ+vE+MRP7kBpnMytWsOHhuuPOh+uaPKmzoWXTXin1IEMYd2Ai
mutwpXMn2XuEpejl7hruUoPaBKvd//5NfML+zIxanyvJC5p6+KwiEJiy7BsvLpYq
yEdW1YckdbP3VXSKDrYQpxXsiWiFSif3QqvkJUZkHQIByxb3CM7nSJi6UXOyrNn0
+j0OwLAL7Zt666WD99eWKf+zFHVmSahtBrU4vgRjrBhuKRjYgd45APNpA65ekGLZ
F0IWxKihrS4t3tq/JSf54DGD+hh2lmgioJ0Bgn/odYegZLCqG1YdByr82vHca203
ErCjkD5xWq/GMQIoON8X25rhWIriWSbP6S6tH77uV6s0M+ARYmUbSCgOpZO2xGuB
dYreIPeVOfytjznh/rdO4Uya4c4P/i8uhoSv2TWGlCoI2Y91MYHS8p+8ftSifTil
azsV+CrxJgoD0uynY95au2DtBEMkNW+Ls9WzihSCVltWvqDp9aJgM2UCIRaFvm+z
aqNnx25qosVvMyTYg5VXlCcHoyXv+RuCIlMqjammJw/V06R2AuxO3W/xdE6XzRHj
6RLAizv3JAMcvoRkqfOwxzV5GcbAJNUjmV4jnyz1bMnTT+22WkXTnWXhszVk9wP3
vmjYpp/KdojOJwSOmSPK3J+vVmCBG76nAQtU+Clw5mErsju8qA9IKJVoqtfn9Bdu
ptkoZV7w6EfsAEiy0uqbmkx09/kMG/joKXHvn5+x+LHtNm9tkV4sb5/uEwdzuUXf
5dfV71huuUOfY6IWYv1noJucL3QQczbquheE540xYgbbLKHpNmRT5ViP4LCv0/WI
RaAdjnqGDGJKfIGqjikpqVQhBMCKQOv178ilHL7ODI5PYcctLAP92n9heMOOeSkv
xmbjWXr5iR6XM/aC66OQCIvuGu57e5/y0tV9uJAtOd7PxcFFNSR0jP3aHp6LdCOx
9aQpTGd1pMxaBMtPfNN08bZSpZHVgZghKKgx1nmc66GQyshJ15Btmr4si+3+AQGk
+/LceyNpfljUjGehhdoqRcZz0ICkeu7XW0d8HIwQ+DgmskBEzlT3QCjRwsMN1zle
YOV60ZOSfvDRulgpI4zDUN6I192irMqkcFJujmCNNR0ANWdoBPUuyJwhnpoezOTc
JqgbSjWdQ0XRS44fbZxjVlG9KeyPi1UZmSlUrFsb6ti6ECUYuvZix33MNk66PTJB
n2pD7mrgh3VIke0Xgdy40z+Rts683UNL5fmfZMkw0TH+S2Qd1CX2CVX2GyEQed3G
W5xy8fd39O60hPba1cI3IZF37pxnGyt7BlFcfmq/rnp5NhYLfweaKtd30wwstFx4
R2dq5jbFsn7BiPER4pUY89cK2Yi98ErnPTY6wmLE2WcpQfsi9kfKF+nzbBpSHiaU
pp79T8K+tQjTCZQM067Fgkl5ysX6IaZ3Px5p86nWVKKWFeTIUsJpLFk3TFWwu7tr
T/Y736dq369vYeZCR8Xj4V5GDqVWS1MNmACw8GjRKwXBGEfUxHh8kysRTMcSsmpE
tvB84HBk74r99WSMOo0rrWdZZQovHVzY0TSgBGY/yt8ZEYST5o+ysXDy41VMeP4K
EmOB1Fyi+Erm6uL7nqEmyrLcfZVsXAvizFKMl1FKf/MhPp1uHIhWR+16ihEqcmXW
UKAKiAMsj8u8S064/tTagWbNmA86465EvTVQFELDlmYxkqTMZJpzI2UHdtqv0dft
sniaENlXmEervdnfJdgq+HoUMgYXlnkAokkzyDrHWbuGXZ+sGDrvRUYHqKmwhujJ
ChbO6cBmDb/iHr7FULfHryXNgek0sqwOECZn6WWR67aZxEUj+9b7GfxiLlIv3kUd
K/iI9rnnfWBx6n3taLvJPOKtpKCLBBplvVg1F8bwJTwAKa5agZQM2193O4SThRNI
2R3H18P75pGgeaiA9rT5kEW/OeqJFJDUp5uCXEWu8qKFnhaHUeVSCaXCOeUMsRr1
4zmlhqb3jd35+BWwi7j0pz/VIeuTrbFUlUtvC5n4S1u/LMxaovfLaGac20ZJRwmv
SAUJnGGSKe4fzm563zhic88xjxrOENbghzz6kr6ThvFUZc4iXkvH70iJiT1ExLWv
/aDr/t7DWZNkHwF8HPIElXbUrLrBXiiM3c+lAL0h80WnDpmqEmZM2wiVMBu1W6aW
PoFKFjf0Vp/T8OGBbQFmzJE3E7qfnbBikUmYDe455gRBaraesmbFne4QUQ/5+SPb
h816BIERyj23Qp4YgHBTOg5tXlAo0p1NcnqZh2oKih6N1ZsfTS5gi48uZCehQqMY
PBC3k1iSQH8t4Zmew63TGZ4seDx8PxV85XtTUmtZF0SK5AqS5+PYYD/78HbfGbtZ
ju/ldf+ZCJ/hGPN92liYCr4V6LZeRFCfFeyprPlU+UDy/BojYNqg3tGy0ejmKrbI
rqDoncFWlKkM68QPaPpzeXw7xkMIMn128npV4dKfEd5DkZORwweyTvY+VneQOGFB
zZQ8KBOEjmH5PXZ8ufvBN6ad2LfVPm1PgEYOLgVXdcrYNRdo8zfaNEaQMCs7UuNV
GscAG5srAC7vlWHHFzIkJlRmlAgiVezKeVvZBzzAqdGtAtV/TxjR5Qdk+jFDEAEo
u6ZDia0dseyF4pDIcIWn02l9wmRZnqprYkuGxUUnJ5/+UonQ+0h0kO1qKMNXfVz5
JAsOKMr/T/GSfNFs/bXb73Z9IRrsdWhRKqMT/eKQ4L8ngoqp8Dh63oSbbtqe0oiZ
zT2HdErlwELTMCqP95pIqjystpG4TfvtD/G1py/oGbdX81ioxDzm+GbNhp7vVTpu
TjdspO5Hy2hnN856ihN44wrSkL2OxkxPvUOG1skXd9ZGGavahIn/8RYXXRqBK/w5
xtxuMPJ7JJVW39qhsKgoAh/JN399zHEQmNvFLWFGWuZZl/3fpBPCtbW1rIHakrw4
FdI8Zh00HZNshPtRMkayOPfES06QGvQQbHBwN5MEbWKLd3E4anmOrNfZZVkDjtxS
i/3aDuaJeAqMNzfepO2UTlSKoW/fbdR7WFmHgUV2v1WZbksBHlp60eC8RQWurPMy
LgLBgj0xYPEqE1/M74PkIfvk69rOnkIZi9nKSO2qZXbHQKQ6vb6hHnrjHTJdxz+8
brdXFRt3mBz2Pv9Q7wGD4OGyc+EHq+jb0exNACgL3x1EV/9lkg02c9kASKfVvDjR
RCPte8IT3ugEOSBR7BqX6+eM6vuk8dOf//qyCxpBD6PipT12tLmT9qyY+8iKjxpy
qRn3ZM1ADEVDBXLyPdR2bKwly/NNGz+H3l4ZsV1j6AFUqMmGfyA+VgIPtBv4pifw
ddV+bBwXM4qaovlBU5TWFpno2THcytcvnx2v05cFnya0h5kLy0rckuweKONURK4X
OjMh5wwNVGvlNVxcLSXtroJAaDlEmQpMQvMYnAzkJbSw4Zwxtqm4c0KFT59mWlVK
oFrd4+H3P/8DNSKOoTH+c9lroLVdpBke+QVda1kSDbmODGKOFzDrZtZ2y84Iuryt
GfOsOa7nOb4Llx1LfvWIMsSj41a1U8/DWgvI+MDWFvqHjXIXVcLgs4gkfOmm4ujh
8VgFCvzrxpm9G9CTnAg7S8Z+DHMx3BJ/OZgAqyfpKGsCqPU/NlCFvmkhwig/ZvW8
YGB172e2rhE1Ki+o2cL4aMEZ/dOmiHK8V+1zRQ/0UbVFEfPzeT3IBpnvp3FSqZqX
0gzXKeZuPh4O+h7P4Kt5xhYKw1tGyhOi1QL8zU8u7beNYAsurFbUCgpwW5RLH924
NnSXsjI2fS6sIDwkhrQsqMWQcKi9YNrmcO75dHNJGvuLSiJKdg5GghVApf1v60nw
xGg+onHFQHWM/LMHvKJVlrFx94KEWCHXf6TKngbieWYKnyaAAMU8sjbs95UQb9mw
EfXbwoLRUZmZ/ymi9tieICCY6m6qDvZ0I8aNIUgJEQwvuYLnRio91zgZPwWvdRzu
L1zd2jGFNNwJxJRGfoQQCGOR0DMHRm3BKWh9KKI/ssyg6VExq5U5kiM8vjqUrWhv
KzCKC4Kme1KbT2Xze79QNQ6/Sm8DBoVDwpszWZQlTmgCS4FvB3pTP0+zgdIPU4DX
AKLZZL/0wOgk7CqYVPs9ppJ8jbjzr49LJOcqQPloUZqZ7b8cnO6XjduRxDOAWdSh
GCrqd8CeU0y9PzAbCJMDdMX73mOeCZYLNMBUDmJNzsOsDTrPcDXCYpBVYhfrLeFa
Wklc0FLrDpBDQLTcat22h9mQg22Izt2x43cJCSs8ixh+QxY+rjS8+E2z+YZUvWUA
jDzPsolbakb2F3Nnv8Bh8GGpZ8Ny79CuhVP/7Jjr5xVVPRDfDsBaPZ8YbcfSoCoV
MHwGpJaUcK/WxYGVzmpIBrd/b+YVbmBpToAZK2rwbrIqiKEWzpYDmWaLd4gWupjQ
Wu5HrMNsZCSOeaPH/z6sVa605TKH/TGettZTE9dx5P5TCxT9C+BsH7bJsdaYgBzm
AspNQ7GJ0dUaNr/wBIrOArZI9LD3A0vVB76L83WijDvy+AjOCGNEbFJxiQeLzSIy
TBkHe3lwkrqbTwrS+ppGg0TVAM5MIkExGJ3jyDrnYCeAsYns4K7OoahIBfvm5Zvz
fgOQGjEEsqtoIqvTeUHiuvxOBfxN7SJXoVn/WKS1UsTHOCVy7r+CLAT8uGasKxGM
po+mmdf5xv0GPUFQd/zqYcDzBj5GU7sQHi1c3sBZeKiVzJBEuP7AvIarUsRWxPj/
LTXMliwSPSYIi+ZonsB/e863WWLMpZMCI26/9wkmJZYukqeZaAjykr2cwHkgIbla
stmL5ohhTQwvqh0azbQnSW4x5rbvmIqGx75eB/5wgyj9Jlgy57G/Uy+tpPeA9Vf5
UfOPV6KYZzLyGBxxIrUhOF81KXEl6c9Df2iOtKsPw8kOwUJOcQdPG4AJm8ud1QVK
iebgfyWlOMCn8kLtfteVD5ZUVfzAdy1c2AG7irccMLjeusdla/DaEc3q7E/DzYy8
PnaYtffksrB9Bk8gi1RgQQ/38J8FD4RleqccGkfpECWKpmecDhve3P+KP8vVmvkG
d7ZFmO1SXXaUO0VlxUzLjuDY/FBqXz1gPwUoHy1ErVveg2Tlpb+qSeWkBBb5xWTV
NX4w4QPyqYaqjaCq0B0Bx28CO/FX/v7tyjGw27geM8f16vaGjpZGyK+E/we3MRwM
3d7SJpL6jJ2hAZHPvtZM1Z5MnR1gGc1aaVEMND6zqyJvJVlAYV18iYczNmEu1JBK
XJ2yp56hkTx4epn/ixnq5qmzVwbazaONU9Kh/9W+9Rtba8ZXMAtJnKfvGgph6sEi
yTXq8WwGT+FUYMFMxFVCNEpoucKFHIq5Xqj6eG1eyo5nrsBbmSVuJbEavn9OhDiQ
C9auQoWwnHOOWm6YCcAsR2anJErAcprhCp/tvtCsoH7RGHe9ipUJp5p6EZu6yD14
Br0BTrhwxrkY/R3cdoJJPAmEMtBYwz/i0IReHdes2fm21SUPk02W6F9FKPLD3gyu
9uSTSJsQoNKGYipOCHmc9w3PtxlqcaIWoQugTemvPelIvdeSO+CcOaPYgxPhlL+0
lL3m6CquLnc4oofebSOLcuqrS0063kdENYjveyAK+hZoWA9dAVcotfrygOj+dsX/
X0vJfWua+hVExD8NYQvJITSan7iucrIdbAnNPp/yUAUTmwXeQmR/OXd6pbM7+Kpo
P3zJP9mfKZNl2+wda7B6NkyG8wujDCGXI02aaZF7xA6xDxVddB+9ZJlmpSR4raWh
y4zX1a9XZIKP7z4htwDmlTC7/Rb0vl8AEbrvlZFdpWG8hn6Izrf9UvDbbrQbxdsH
EmoJqiZPHkwCMeCOfEG7rbMd0t/LWTgZ8NxAtasxEW9RoW/bdLJ2pdFGVlSN5xMH
7JXG1RlTdRlVL85c0QUlecHEKxn91BWHtLyjbIeG8FsgNhpaCe6HQEz4haHSXSw/
qpTukVJjuoianGhs1gAZJFsNfyXUP4Y/tRXvenNV1kfg15oHTiXwDgR6bNwFmpaD
aLl0CVqR/g6pjtekz9kfap2IWdTy9ke6X2euULOyJWSKNl6Meyxj0y0DJhxhqQOw
oEo8PkAcCb/iF4TYzNCuyFmsbJMabeE9MdWrUo5918UppksfKXhwUvE8xJL0XgU0
ajtT5JPlOJDztQANrsGIvOgGMhbfdtAKdsFnEYFSL8M4vVWKja0FXoKRScLFgA+Y
I83xYGd4pAYqxdGxTWzzfKVpnx150pdWEdPEeLzr0gkXzz+QVdK6kak98WkO0lNR
rr1tlz0YxRC6zgW3PTla83+E4OGaDPhJ1Zuu6bMxba+A8OxhC5/AhYhem9S9sCPe
tf3G2bws38xJnIv/58vI/7xlnfhsdA5fyENACiSWNdaBpFnywEEKw99Ga/DEyK2y
i7oSgVQrsDDb7r3e2d1a8NeBfV2Hf/CPRHny8omy9ogKExJGZCfPGpwfg8rWeEfn
yULNGqIUq3ISKkVUp2nR6T7tZAslqqi3rxOgrTErJwOitfaKiPtKEZMdyZPHVEOH
m3tx0OUUAShKBNwae8vK+eeWojSEKKlD7y9pfmezJ18G24RaPeI/irufgi/AzqQe
nZD8kvda6rMeXOKLzngjSKKJ8RTD+dl7zoJo+yMRBvImMGADGZjHWkGl+I7M51To
S5TBRTjPTuz2sBtDuUYmfqYMVUBgvFRIK0UDoZEiTOh5+tatM8D4TnpRXSNZZm7s
WYC0SAVXaNBstyjvmF1uxyu1dnJvHbMxt8bpE4VSuAN0Q/mtvZZ/OiSLdfHwvFmg
HH96Sip6sTYjtrukbKG7i4kuYqgV0bqvB9YW1KBiSW2DXxBq4Ty+REdgj+KIq1Ns
WDHc//giwlpefiF/qW4cQNbbPYC9W5AanToUZgCBacRcoaAehTqJTbbSNmz6XFJy
c9fJ2d8oKFoJOx2VNSni/SPe82Llo/bZBXqi78jcGkv3DT868nGf6Lgc7K54dsi7
9l3CztTBtQ5unVFRtxDuQcjfB0ENP2bHRayIXnY192BSl0DtpKnwV6RL7cTnbCIp
HV4DbOOC69ps6rGpLnW33PwaZwv9ruPG8YMjU2ABRAc+thYcx59jJyqejfoHxuV7
gEI0rrZDtAJnXqdATxzo6dqpAgfDuo1litrDvALBYgviOk68nHMOKhYhX1MsDacP
7x7Wikubmxr9LbVOM+BR/bX0XUAMVA2TO7BL6wpgSH51VfwddmKZWT0da1t1hShG
zTNNHJM/50JOIVlZ1T1lFRAJllZlC+HAnVJ7gvAAC8pvH2G7DhCHYQtHTWGrP8eB
5s34JohwGqMlGyWl/Ub6omMkY+AVw4sYfx3jslnm1ZPH5K6hRqBOGZnCmZdluciE
fAuZCgS58rKyHy6dxn+YlD106N2/g7GKZ5gFmtZriDSjIiHRag2asHV1uFr6x3CJ
fqINTCvGzo4O2ShK5dRvTDbkND6c338EYxLXbMriF6rJFn2EhvSDcd8fMI3119B2
GpGTHmJrXox6+qRKZTUnIyR2XYeY/b91WG7YsnH07GRwQJ62gYhXmYsf+AjyXvPJ
Kg478kp5gQRiuyURY09sZoEOjunLfVFMlfBcc4jCbDTwnAISD74HFCpX/vwbsmug
8UhTJBfIDmQbh25xJCz/+RGbLw6SXw5zH4YjE8r/sBW8IUjVn3ctzysVFjqFgoB3
mC8nDVyuCva0gOb4zFpNL59vn4+GNvtvw/TnqPKeymf4HTjRYCy9pNAREmbGy75S
EOZwzk6ChAx0az7GwrBF3d7G1C8qp1CmCWJfLXKRzDZSNPhveIvG7Nh0EpcRPt1f
cUAOSrvlA1WO7A0Glc9CpdWtDUHpuMpGtC/UUU5fByHHufupGLVKi41TQC7VZ/tD
EIQBErnICthChCMkU6K0WJ9GC7fXHvjeOYxBHuR/kt2YGaHpw9MxlByDtRL7efR9
7Mrv5Jm8owsvlcoQmZrw2r3kYtzB73OCumtNzYr6k4qn+iwsJDkjEqwgTwm/Xhu6
lPezjoszV3s0OCGYH6Moby5+PVqlLWjj8Pf9P4lbTPY4EZRKsjMZI7B22y90IY43
AkU556nZHo2T6BswG/pMpK+xE+5QeiuwpJ4O4MjMSDW7PXCcaIXpqU7SaOci349l
2Uzq9NaPlkELd2fL1cM0dnebNW3UiEtlpCNpTqYdRasH7tWNwFUSzijf/+Cw+1Of
CKFdwRwj7CmnG5gy6Ce2sJd/bOS9pMm2lVYx2UBC7GcZVTdiIRxORizKpLYFkJ81
5J6x8r4yDV+1nAPa6ONXx/Tun0soc00JqXaxo5joAq3wqgc4DkUDSU1Y2xKymj5J
cD5vaP6Yw4WYf/00aClEBlm6GhX01D6ms6uCQxXkMPki0VZTRdfg3+y2IcW9e6GI
+SwawLP1QTE/T/DFa5cs1VW/xNUSx7tUdOZZFOLLnbbhyA3Zm7B1XK7jJsnsimej
ypb+k6gEpeEDDiKIEhF3W3SXSX2qBS+xsjq5zHOVOmBvIIaZ2oWHg1P/X3hb2yqX
7rAcgZr9GwxyIlslqJUJ1qAx4fBaQQz7NP5jLrR62rqGea43LUJV7KAeAj3FbGZo
dd8O66lju9V4vgqPaDOJIUeIFEfPPjO7CD5P+gfMhxTgd3SPMOWKTbVq0mSkoGUN
AiUhaN9MAVRhZrkstJDotqpdOR8C8J60IsFMT4l5+Ur4Evwp18vNtzxfr7lEXhJP
GaHCW2s67VMiNYPv8xPdQ6d/hbv1m1CQiAalZHip/j2MFBuJ8UNDKxwXgHIsDgVH
qpRxpXeNi1G3K75gZpdhGqusLuAIzm+NGT/50doiX5HZuvTjSuSqhsdwOHoYI9gE
aGiaN5aZdTPVJny/5AVg8LZNktd2uf+7bbHXyWJeYwTuHdZHkXVShNxCfKa3CXPF
2DgEXQHxtjIiz12MX/B2NJd8BH3wpxj8PPJTOXR3n7MbTGyF6qVd/eXLPn7w4Azy
RvyZRx8avnSo+yQ0QPAa03XYpHTXwM3P+xUqa0fNzLeZ0IjRwZjLH8VGoO5JH1gs
yXKDCjRrWWdrHZUnlnrPxwRNuo3LDNizWsxK0FUz+TjP+48qZFAlYAuIjRm8T+av
jK456sG+He6eo2O7ji2yjA==
`protect end_protected