`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 43504 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
YvslINJcsdDabhUxdg24ayBYK1KuWlzBVj2WOVoyLNrNDydedPFFXXdeb/WQ/Cv5
Q+n5Yh0xyC/hkMlGLBGwCUsD6fxfrXZYQtpwqvPtWfmX8XveDFnIIvsrXN2gM/DU
t9xTCEo4kOhhNkfnXUOHpD8VauDTdBIBIzTt2KWtGVnXiPNVD3FluuC5KdQ4vmp+
AJztZVDFQcckL5bGUcBtOLAR1KoR74vRMG4hrGKfjt3csqcstyJjoI34wlEIXmpL
nhG/4QauTYR39YbwZorV41decWIB3wHDOGB1wnq8CmRaUCSGZhhaFdM39oeX1Bln
zasLzVqqv0wWzByMmb0ZzkQT1lQRieY9A8J48R7EICSC3X3/NTuBLkB793gCwYiJ
Bov9Us975Msjc+mSEX25Fz1ITczt62wf4OP0iN/V+081qJOLerHyTR6YcxMNWuDM
aTDsjtnnwcNWTdyayjXsya7KNJIcjvDZ/c8XpXHWqM0LOxd2cvnwijPn9MKQmsWt
OoT34qfuGnJu+Mlf6yVwIFyzC+FaETX72ZZHVYK2cnjO/Hmky4JpLj88qUwhvO3L
aPV4DO5aguK/QmOg7OAVrMc1aJH6K/LosVront07CLnQkmR9Na8EM6OK7ij+jgEq
0UJNa1W7T9YpsfMZAhDYihoXyOjmaHyMKtBc1wDELODh4xnif82HsYNGsPSZTqn2
eCT4S57uGgdfw4H85VjbCMemRIfhfvAe8+Og0mnXSFyPFS+44dshbMMqfZAXE4df
/Hld+eXnDT71x65prWQQehUD0RFLFD7eFHcNOf0iDyBnNi0O3IztV3t13JhF7Mdh
BVe2DKidRvhf+EbWl5UmzNb5MgFhnR7UJaN7YaXH1NygOSyibzWlY6WOtgpziWB3
+T8UfGLDG5F1EaGgh4vV28lywpSlv2Q2yGXpXUkN8yfZG5D2kSE20uyWRynz3c87
j67ZaHsD+y4JTWIs3RioHKHM75bgCEo+USh4/o7yYXacrxCsj4qmpnjxDoZr1dSv
klBceZYxg1ib98O8GLzUtazPC0CxisqbYybazotMQWGQ969C3eCNjKHmr7WpWqu2
d9xBlmeaX3TFFJ24zA1rNvxi0BUS4sS6889NwxawHvTUDMxF9HbAHkpOV85kd95Z
5EzprxbbR/3E/rnv+rcRGWFv2SDnnGDTrWJj1nyqPITpr1zFlRq7+qiaHBLmYWa7
3fl0SkeRWmFn9e7fsGVHWeSJfnLSNiNknxCvF5Uw4JtqNwm/HeGgEqN7lPO0r64a
r8eWZ5MEdW9kk8lJOGj/alYeGfX9xWc7+8IVUxizoPc4el9IAig+vz3lK0ktzmtf
HoF0cx0cxiu27uNP/RG4FdUyyWgI/ctVfoVlBOPUMd4oOcbNcAH9PdfOyc7khk7K
7g7znhSgJQ/XTMtdImEG/PYWRLCa98APLCfr+WX8Za+qPWGXTU7I8qWVOxjw+nWi
xZlcIYwiqPapNWxjJe4tByMaPV/e29bSYkUCNTxnFlD+nxwpLZb9/b6rtKgZpoSP
QCfdVfa8npPPmX1F03S6pc8SHNpDp34SppiYpi1VbIFPkla4ixqi61rNp3/zCAXH
Xl9LfyzNvQTDFeVMDcDR13/DfdP4QmCWSnZ17IRBzUYGk4cnbDsS8Yvob3hpCtUi
y5JB2BgQfWq1S/SMpifzosCG+R9YQWqNvSz3ScLeC7lVlXQ0vnXbGK8b6G5/P35u
3U3m7lJdXq7YJkWVSEKvFA5Nln3fwiKwaGrDaIRUPDjR5OPTO0dHdqk9SJBIdSlx
Nti4dNZcFqFvJDsTeYA0A1NVSqzOZdGLENemLnqP+BOzY8uOmRCZWvri7ZN9udz3
Mk5Hq53XqohOGGOzZKMnh9BYiLB5CvUy2YezauXQlwK27SNOiXFh8uzDJoaE5bEZ
Ns4Oe5oU1w6AYjFhU59CLFJkP8uwO2/xP8AnhQVPiQosmew/cbD4QeQ6bZu4hF2u
RXQXMMtV2tpzLi1FD1/siIR6mBwyK6gRwWkGHaSfOkG8/itddpBwYHJAiXP6Jkru
W0ZPzZCXcDKVXV9jKeb5y7FtKb6CyJv92JDVQKE+gb7h00do9vtqR/4/LYmE/SUU
7CXO8sWVHgGCwH47H+vHWROvXSGd5di9O0DuE9pjzMaIT2asCr6Z2EHeWH4cjsTe
hYClaZPNc1PNGUwbxmFVeoR9CQkQZ9zuAmXQO7Wf8dISZ4zTtcl/8wDHqR+KMXV/
KyKLqiAKhPsk7ctqW0F9+eVdCmjHdIemDMk/Me8hTgsHKqSDnSHJ/rLfieNUOWRB
F2LyaI0UHSEtZxkIYRaeOOrV9UFrYkf2pwM8RhofI9+BQOeE1Nv2B+0hnojFlKWY
LAUQ4FAx297XyPB8mgesh7bjK4S90g8Ibz69pZiwRN2JBd3eLtNaQSoEzBNMHscn
054rhb5/BTi88Ld+0D1Tlq0ccJ4Wd/9ja762u42aRAJht27rDTF1a4U40AaniIMI
M3o4lol1EGu8E1yDE934iCQdTX1k6rK1hcxVf2mrn5/w3B0JoQjfr5rEfjNhFzMZ
nWYUTI0l1XCtWHU/DdILTJQH1NGe8Cm1zDu+2krJ9Fy2OJc2cnDENVnq+7z5kSS7
LsjZnW5OSYRG4e+bIygGgns/+JcbRe1ibGhwPoBhFVkGXv9+TQDyvjFHBliQSEzQ
e4hPtkTsSBt65WJZKLXciXMiR3zynIgbwrANOeszBM3k1edZeY7KyTozM8ezNPAG
r88FwBWWrHGqi7yN00+aon2ueq0l7lIZvDbyQBZSla1g3YJRV8lfugBpjzJjnfeG
CF780H0mv92vo/oAmByZgFan9Gd9W5jEcLJww/A1LsY0P3XEAMUC5K9fvJK8DVQT
qC5S9j/VGyGKlanzaJkm2HqdWutQXVT498Y1veePKXHo6OKIWdqUoALWOvNeA2Fn
R405Ftd1dOvfgKslRMwcgAUcgn3D0eeFmhqRGcndOwRTXY0PkeqnxHqyQ/qqDMH7
nLRMTJ+NGGXt7uCThc/GuttJ6sVtp8Pw7AKOZ5cQBQQrBlyikYHbfjncL7dLmVgv
LASbF+dCuQaNNKh82nnG79ClJgZ9Xwec9HKHN7ON40e9wSH/PZfuo0WRxLC9zPja
z9YIs5lkmUGPerWmaxwwCvfoVVSKszo3SicRkAez4MNo1as8sNv1IJ0tZCSWH3Bt
dKwCfar8UTAxZoyZp6crIcc1ofyDfhFJAVXt2ylGlZOHOGbXh71VgRJ/GzGzlGlf
fLOmuN8HChgnkJ+aK0Y86YuWvoHEd15r8xSjm3XZ8YJMWE+QKBwScPLiej5ZflML
aNXHRp2LMr7E3yZUrvul/Yb69aqxB9h4HuiUNg6g/uhgUKZdJZBe59IxkEWjNdnr
QvyaEMfj3hKBi0FMW7yxg/6Q0N3h/0mpGHI8SXNZVNAmnA59Sqx5Yn5Y5LY9vYs3
mVYTjIaMrvmKIlYEI18O7q2+/pJEzZ56vvHULHUJDohUsjkTe6ceTBpEnm1+CIKg
gSaDDzTUmbY0BAZ3YrlxWOqprdOv20M3aiRMD6KfRoQzkvou9f6f1uMYWsbavmdJ
SuZTHrPCjuPS1Qs8tq6hOXiAUAfaUWPKho88QirObE57k5/cdLlyWkets6y8Yqww
OwIlIwjpVAx72WXstT8ze/pm0d/JuZk+wvGkC+y6T+NuUo2z1VfzNGnKqgTMAEwB
O6KuyI3zbdV/ApEweBDqNAQNXkC2if5WQ9ZACjrcZjCt6ZUydt9/Y9AqTUav+Ea7
HW+YvIFHTQOe6R0Vrkw5mw5T/lrHYcG3PqqcmOTQw87o/fnX5xdLeMfrKdfPtg1g
Ph3bVzDc4oA0RaHAiDfds5KdkDQymWaehrPut/Iq0L4lHb061Cz227oqTIs1/rBH
c9fcog8uB8z2JuyjplRymIbAqUs/DhIKRsesjCrjlx+hfZKl0KxwDTb7qN3HAbTp
w18/E0cp9TK35OEkRASFUhDytwWhmX8bpgelpP66afSShwSesNCtU8Nc/ZEoUswi
PNUXSyIb+2nb3yAl+AUWtH6w2vppZDWNueOiE52hAry0CLEhZOs1iNW9SwtPYNfd
sxG6qNW0xGBn/v05YIo8Z7MUsF2E/BkLuxMbEbQS5XQOx1HG/vs3Sw9QbI8eztHo
qMdi9EN44gl+Ggbjbub9vejIs++smKxxP+bykBH7mRuqJcDeXNyzyZVIYTU/yp01
VHh9EvhXicPcfOXdp3ui7lSR6UiOyicyYNAAXmWdk6bUa5a1fvQzMI6S78+Cq9hV
C9ae72MF8R9AmeilnqUdFzTwBcVd5G+X/YesdRc3MSz2NgbjQve1w7hc0GBQaMs2
jmk8SBX5kwUmlmt1NsFOJe4alAOHVQVDW8gjpTsV28R7Hq4mNpz9YNCzklbGb/C9
Q6mfaAwg1l/nWdEAapMED5zAmsvy8ncXB9/7uFve8KnfPixKdlLkpD7E4cXlwVms
05AZo3oDFI0E+IlcJENxlSvEy2YaPp+cyb0GzJsYKzKZdsMi9O+aicZ+Bkc2r5vN
q1AJhchgdabGXy2VwNkPNzPT5UqdIUDexoFU325XTtQnuMdDZo1c4Zf28ZdHXs3A
AGZW86J9WhV0xaThhrsABdA4lFhqqCMQtl7b+50iAqEfX4NEpZqzbw1QNJKnpClY
o/7yrNImiakDyArZMvIkwut/i4C7LIYYesrsvrS2Y3jLkcOqtCbwXx+yHRsfG9S1
UG1Xn03ifdwae+EdnXgqhbGlQI3/56LCuqVWNjU7PY7zq28E6H4X6TrMA/mcVYJA
Mekqlr9mgOz2xoW0M52CqiYteW/K8zC/g5UGUO6Vm21gEuvJTunST1CZOqM7GbWy
IeClQcqsVU63+vRrUvfrRFz7gRqkj9oOHgGv86AGTP0ZEG1EZCwLfXbpVqYyNocT
8cvQRRQ8iyaQRpnbfkWK3YmMO38G00DduhSl9bJ4MmaRPzrl6KsmBX51yuIvuCPv
nyDf02DxGy7Ab9jrQ6JXOXVzCPdlVlxOnrL0Fb81PogLnq1Ndoizq09ps5ccJOew
AQ6mhr1F0C0eU8RNGEghyHtMajrsvDxanyXp2yJSFW4boOTbcIVAtRqlZoEH6bVU
twRt1rtU09wCjEXK9jzcAq0xKrelvRg1h7WGUpOXb4+Sab29XngZyjaDFLvjADfF
IB4lc7bwisW6Csis21ePCCbecFVz95CzIkp8nyrCyf806Peeqk076xaDoa5JlPYr
k0EGZCB7+tgPkDkeTdUklcJq1jDV4uSO6CRE/REayRn9TOKkZD6jm4Up+QOmZszv
R6tV55QaTrklzawmId+hsivFvlarwqwMWVTQUtdHDd8yNHFbxcwVwWJlFpyUBtBr
Sy2CgwnvHHml/7svewcQQ51AL6Q4tkw7iyPfR6EsRcLrkKTYUiTYdo6CccjIFJO6
cQZaEHcyjjBLLz4GbtaXtFnCV8+9sZ5cL8twwpRyz9cxbSfVQM3OeAFDmJ593MuQ
KAXjuR/RdqG78dfbP6LFeP66IN8qAme57ouaRqBagR5Yf8uWTQsGYTUMyMsLM4kG
67ZIkIKFdoF0Ks+bDeeE/Ey3LNGlbMek3XuuvnPLOkQSyQ/iHEpjWnqcDj0fuPTQ
bAOf2JIZbWxJuYZZCI5HZhQkuuu3s1yrr8IlRigblZYptyTqvoF2E5tu4mYBN61S
acyuKGFQjjiM57YYoHUAb8TsQ6BVeHYUyxJfnMdfChv7Ytj273L5JY3g1FXOkG7k
eYiDiyuJtiocHKdkhI1hxHPQObgx4AxiBWnsfc/sehmIACoZRMC1v86MVxgJhyee
p6R5L0zUDV3ib1hAf4aSgkHWOznx4uyDYJSMYaSog8ZtDMNU/Dkfc183BCzwlqtc
r6M9Bat5a6w96sDudT7ih2u1C/b2fdevQFvTs5RN/EfzqgSF1qCovFs0Aujrcmqv
JLojukTy4EoUqxF5AJCLqvsDlPiHRTRJYoLzZkNw5TKVtoJDUABghS01HVwseZKA
8DN3eNNxgEX/8HEYIlUUKDNVEzMzbMYCX9gREUvm8GiyIhtJggpuMGu5gWQ2idjM
dI4/Utl7PqF2zypGMfBlZzXOLCMlUHIEMqk0vxyNnng2RjtqOgOUWEzCnIsxF+gY
2eieqpskiE0zScQrCQwL2r/8kdDZ+fJ1T81f1QgaoH4xow2l7EZxwEpSxA4AAjJK
kWKe8stwZEGFq/arcHvD8oCSCGf4UT49Vj4TdJEvKm3wr3Va3lDMqUwbF9c+DSSq
XOh7RLrzdDhJtPIPsDcyiZcBR/2MYZUIZzNDJv3kirMxy3jDbPqqktdxc/vtA432
CzMn6Ct1cbfuSKcULXttj1J03tGF8FGBzUAb32pLE5mqyzinTx99MHJUX78JDKG9
I5C+c7LZTsiLj54GkQ0RL/UtRdyjV+ZWgZ0W4/FboGYcc7XpaivdnEJB2HR2vkra
9WM1trD5TdsBijeLR2I3b30treKooyac9qxwFwz1vH4DLCRhMU4eZm0t9uDA9Ugj
vqFXnaQ41uUmD9ueedxAfqjKmhwpwWryZ+2AFY26ButdJDLkj5tPY89u3n3JI6m5
f56CfpAiM6OPKywSzSWu9vcMBkRhNW+F53flHWZgGe4sYC8TzqQHIrmZwUqf5FGG
Rs4U2FV/RLA+3mzGIe8ve99XU/fU0HmsplTFNxf8vHGQkJu+w2YcVXGVh9G+Giyw
pjqHGUQ6POY5QuFA6aWt7jFeAgcmHlMu4giEdl6UU2eZPMCjmtqs4ba39CpcEtay
y27KM6AsMPPoKh7ck7HVzLCM9Ky3taVTRghXjki9SJ7uqOc0MtI5s05eQnmwFZ0z
35MKxiL1QfRteLkqeLXfNTbT2+r4/7C0RWcMunwt2ZT790PhrVogWK2DTBjfrFvY
nbCq51CIzp2jN06bzhKpgLw7oFter2sM8RD+Eg5EKH5sZSyEVYrupFiItJYN460Z
Vto3evCBud8Y5QjR0gjiObvEs0/LKR3eecZhKbHR8N9HumPA8N3zSXiE1qVEtwbY
MVtF53Re+D145AkNDgrP8nPtfdWphsMVpKEWAHdhUspP852RC1YuEvKPOqXYpFRL
UcpDTkjWx27c8Oevo9oJpjlPNorW2HsYV+BiYpkCzKVHX6ng1rxJnb2P61QwCc1n
G3LxuZ33U+VYITLS0T6kA8RtaKoW6aUmexm3Ngg0gCVa4NbWaOKjo0sgvfHS2oAB
xG5G3uEcZBjoe6hAde2pFOQU9H0b+85iMzvHIK9kEZvLjtE+cDuOUQ1cF83tixMB
17d5Ozwwlai4crXxyE5xp6WBIE6fwTjAuFxcUGfOQ2ltOJqbT/ZIbSJXDSodi7yV
c4NTnpimg0AgK8O6zV5JxnjbEspmMUFANbWwesmap4QWTVWYugJOggDXrlH/T21b
Lz8ZmTTcYewP+noyEobARh8S3Lo577ZhuNTyLFBLOufOdefKZNdCTqPLu1AS50Jq
qJzjvt1Edm5aql9+DsdUyPjf7aPhgDXyMi3j9cZZRi/vZyY+5ivQKMX/H1qPhci8
M8VPZJgBwvn9T04UrTZP1krKwPrq2KdTUXsCT0D/c0GMakqgfY0pV05eeRzkiZJD
T3N5VQbAe7dWfW7tFPCeSS3082l6WaR4ynWlgxOa7JgZ1Y3NtKH4I9pqYMYoOWvB
GMnvnWiWBERLJcnuRfwGpjgFwnmsmX7qiEQJLofgptFRCrUpq/p0KcoR4GBhThKf
1gVrhRkCo1cCIOKLzDNRWl49aGYscBUNGQKLHkJO/pOLT4jMwifbKDAo6REjxD6w
PUTc/aF2fLELNxMOkKYX9xJNZOSisYZV+jFI30bRfX+Mvybtvgnlvh5ZLPTSLqC3
gFNmVgskZEwkFxcu+jNqq+iZdXeejqsu5r8NwnZkQa8ErrF86m34ZOKUEm7Xns5n
y4od3Ve/eOoDrSCo3H5GynAvwfIDOFAUAvy9qnGKzXwTYRjdOlJWB2Str1cXD4Oy
NSvpF+mG4cRnf8CbrTxsKWiq/+Wbiz0du2afe85Qj4WR9p2CKcoOQDX2b3jmZ6a/
8lMMxxKR2CfeZBHPJ7Q4im+83q5oMvF4IlNbLrWH3dc9YjhDkQf5WIOQpJ8ZYE9R
5BRD1h00QSWv/33lsJx90LDPCIS0U6H+VNzlT0moMS+9bJCPt4LsL771MSaAZ8Vl
+UKyAVZFYI29LJt/yKhPvG2KJJUL9psrTX/aW+2E/myYTtoQeQF5tuZNxA/Xai1o
YeRcKlkIk+fzvAeQzfvyqBgGp0bVbvxpi14Y+83e1YD6+SeFkhia7zqefXG/RKFq
yv7Rrpo80CRMM+DhK3TX6m8TRrYETdZWKFlZInTbd4yJr3NcjZElwzD14jzbqy+o
BsnvrEI9iUJww/jIsurC8x4bTCO+CE/zeRnOYGX3wcRmHADa8MutyTtScuYvce2i
HV+2dqTt2o8y/iPwoYcuBfGduya5LIyG6JiJ2NAc0/onVQPI8VsUoJBxEbePHI3Y
bYYnAaWnBSx5vAPGEnlacGAhdXB39wRlhc8a3vOqnpUBI6zmAy3XDedZKgTaNOXR
9FNc6ueWjd2KMRuPUvfG75CHXMK3EFnbtriK97pfLYQygIPu+LEjX2aftVmDfMvP
istr8kWuky5oKFMN0g8+LS9XW7T97DCAG8OXjHql9j76Oi8WW51NSQ7y4lgmJqPI
VjtcuPdY5TOJFIOyelw1JIsS5pxQ7V8Vkiq3r90xJ9a+ML8Hp6L/n0zmORMLvXe6
DIXc+14+iOcCPfoXodqUiJAwCipBVZWnuF6AjkY+MtNfv5VkYORTN9T2gRT2u0Br
mbPvZvUW6+PtCM+CiD+e1QBCAy+nnxorzzoUrlmgV05r4/0ofofrFm3YPsRGbSNp
eKU+kH6fOZ5iIcYh2CseVDafpSSOqwsbve1XUaiLiKdfCn6xr0tRGeMlOuIuxwlb
EKALTnaZ4eE7BhCKCQjhDYkDekwbOW2vXQktJaZZFIdxQBm4IYnlt/gqkXxL7FA+
M1VbGFgGAp/h4yE8mwlte/q9CyPWZw+/axF426mstI05Vt48u7KV+qbMPLrh/SAq
OGHIDWJv8kuc1MprJ9YzzIyPctK2UHEQy5HEm+OZr3TP/DvJMySmCZpRHLRiSnDN
ZHOKqfhtxWu3InqlvLVv3p7pPoI94mb5T1nI7BvvMCBPuqLo3d3wMiddxEEKlPDj
K7vy6kNW6GEgNOyShTgbKnB7X8u/a64kdSOxUaPpnoPCnary+div4c+9FhFEV+VS
n76Iv2MWGIdsyer4m9jSlRBoQzpKpZtghJUEhCVKUaTQllh4aQV+t7kqBEPGJJrQ
5PSTSWuFvxg+r2g+ADbUtS08Z+nTBbMOQYreVpT16zDSbcttwzbw1aY/rIyYz22l
5n5Ssekaj0g9xWDkyjmMW7uohWUQqcC6S9JuF4FNC7w7Ox6M6pcnfDY0oOBUWHQA
rlawMMkbarvf71FniwkmZBtupVpfdRqlt/53yNa+DhdEoTh0HJJj1D4GpzvVFGdK
dpw0eHGwuY7knxIEES76/lokPMRiv5RIlZDvsZS2rQmiyalF8Y7OB7AFZHYB/6Ua
0b43faeOaY8Qe6p+Hhv1HIDJq3fkp1JBenVUsSRZ+Y6HLl/U2Xx64lFOWCzp8oNW
r47bk110D4sWLHUT7QwuHrZadorLLMu0/oMF/vr4Lmh+m3IDVyn08OMwLCHccYhv
XHLWmNCVFy4Av86Yx5oe6C5Ku7ZPcFholCxEOCIhrWrHe7mvU9tbnG+AHo0zjg2G
8mzqivMDtQangzdzLaVSjP3R/pmA9Amy7+RqHJhVLMWEGA9Qlcr+EmboYh7zpKiU
WuXjJlgLtBitqbaopYq0sm679eoLBEC6KIccQvZVkCGIdO/VnffUarBKb40UlCqc
V2+zHjxnTiUFdERGvO0LDiFIvanYzRFYMAUxVLZzEQuz+GNHIukuw+LcpNVCF/S8
53oL0G6TGvD0WTk1ZpB0S65c+AdFyOUuw/rkrWVAqLpMEXNnrFDSMQElTaVbV8oK
/grW2/ESWVBrNQvCngzjSbNqSRNKMp1yfBH+SKJ+uH2BP7Z90d+N7K9qOky1ArQp
aJfxKCgAbx05yAN5W5oatF/o8aIJenuiYgh8omiWcIarKL+90kgACy1p45nN/SS6
7KUF69+f5Lph/faJ4c3OJkSpRMS5NM7BZJivJDwHBTNCWY/FIFWQI7wk3LwqtLEx
jvGAggPCyZdabHjUDmZiBehbLyv5EqlE29ltKGBUt9OwmX0mr2iZvmc3VQ892Xe3
WnJP/UVGZ5PzYyNPdPEWmRX+Xha8aPfT3CoiTitt/LB2Zrs0iJY3rHPIaqpzAPN1
pOIBMIHyEOGKIOs8b9eqgQtCZzG1fS0v9YBudOKVPLb3WKTytI6Oi4ft7iZKCl6C
xHkZsQnp2bF8EqPCaQF2XZXcQD0y1PJ+dkYNIeJJjH9rSqTjBklzVqmutd9mlZg8
eArpb8ZXjh9d5wavFTKYuwGbbnaURw7pX1eRlMe2t+pOYBBnf8mCjt9/G3j+p/6s
6T/UgWJXQNSkX3e5iywHJH2WrANdv5sxbRddwQyud0Nbww9qduF85/HV+rFSdZMI
mqAUuFdal0utX8ITCGnUI4lIh6gIki3SXZgXfBlAXhVr6NV7Tgq2JaVwuhERZAAi
hUY3oNnf/iJaeFm6TOif+uwOxXCCyoWoAmd2IGu8tnut1xWJbdwgatp+6MkfpwhV
wn7JHiB0w+Fc/LqSMyspis69UqUjx4XpuYEx5eojONgBX87U2pXzUizo9tjeyuYd
jTylC12rfXWF/slQ0+KIXT/54MezTTgYihU7WrLlNgvktej7tlemkTgIOnMHWeLo
YY+OqZMeRffVoVT3xQi5pjV1cZ1j7nEBW6SN/7gzyZGNberjBnonMm+c54OmbFGI
b9Nhs4qSR8MsmiceH6bR6PNcxFkmp3fwoIbRs8SWh7BslLvmS/4MLudneZE/fvXP
3Y22Jk9RoWqVqC/ZE/AY69MTbdFmXHoMSmhgu16F1HeB8fOPdsRaJRkeNUkljhS0
OgudILOwIOHd4/PaZnexILTloBjhvh0CeQKY5HvHyXSBhpbptnAVbjCSyhWhD6Dw
le+Uh1WnXCn1bvbzA/tSiX94ngIz4v4ghEFdjku0kQoXIqf6xDJm3Sn19cSeqRTi
xMB/PoaeaCxHHSZCAf1TTJUDyT+FgKInzs9lQ3w+UWTfMn5LjnMhrgm5M1Giobet
+P/RJarKA4EhdvgRvMl074ibb5grmVJ5Ny5svoVa6G7VpLDkI3XOzCh3rKmtscS7
7qitYBz5jjgUV6+p5ns/HodD0FgoPSZnxMaHQzk2UQjNPE6OeBztplUEB5uIqFOK
fvsDwVKKvkNR3MXz6wk55sv0szLKEbVYg6y4AFy6stDRJH9qxPXLjsZLu2BnbNvW
32RaYXHvFe2H3MlXo5actLVEzW2gjISaFXv+4B01ARu/Q7dgtE+4KAEKEmJc0NL1
nobmnRycYObstNwbd5/9OzH0ntnTA6kuJgDP3J6EzgKY+K8LayK+vdw2yD6BovhH
97snIpgDqj0JA9a8G7zTkXJ6jxPJLXX3F3qfseNloZV89MDSdCisR8Eddo3d1a2L
AxoanUN3zDRrV9KNvd5KNtpGtJ4xOEpqkdbcP74KncxGBQeOwIScducWzXfpL4yy
IW+ogYVY0kSBFVem34UTFR8m4KHmfG7xqvOIC2M9MUOqsPrV+UdejH4VC0wX3+6D
8TJdjvrN/nCOVUjGCJ7uLVojai/iu+U0JsckUVuU29pa6jgWt2BZFuDAICPQ2ou3
dr2+7NDlFYBMhEEsGT2Jt6V0UsAyvr+Qx3sTOIU31vj1p5gCqr9UcmSIMpzePeo4
PYvJQg1wzaERHYOrUvZWPx3PqtdtXGrpu8qNr5KDhaslC6pBnu07yXlVegFgKsIE
abygDN5Mp/3Ju2estv2JAhr9ckdGKzFY6YxlpNRIob/33OXZ8eQAJvZfgZVSteY1
MlrCNndUiwyinKKmE9NM/gBFlc38K7kNLlfZdbInf+NYhAw1DztOpywe6s2VnNcA
ELSF0A/iyXyWr+vBAriUMzHrWAoEEkLfvQN7SmKLJamvBn2pdmiEN9/TmMHhJ1zO
q5lVlH7SkSGl+pC+HNZ87ovQO6CyZSHLAK8TtSG1CtjkLYbdRToonLF4/7LQwBsM
o/6wMG1jDBkpKbJJfY4HBTZt3XNVQaWKab4T/1dMoTHiL8SqeVsQE6WPtRrwQdFI
eerMsNziDHLXxfkqp6F9CZHfg4sPa8wrGJ1lE1QM51oEazMZ6M3NHCS21sTYDCkn
mnGGaJRt6obCcIxckyZhgkEd4HgrdJ45d6gWE51lj5JJkZixp8Py9yihbY5NRV7p
SP+4ZxcpTDk35qIUg8SYW/ktf2TeNWANnsHeTKEqgP8jBsHvX7mrVI4yGxIUC3OH
o3wx0aImbZ6+ClvCQW7hiV1B5joQVjzSE7FAuyNZ+7rsJGNFHGUWGbm7O1MFAeup
KimIiQNzRjih4n/bg1SvsgDHEv7UDosYu0FOMSSwzikRseERapDIlJnqpm1cUSH9
jOh6POo61eXWyxpjvbEdoisAQsf51Kd9twpZuYxUjdVLyMCv/6u/n4eqdr5GsN9z
Me7ORN9qCd74wrxlO8nUzqNlC1Nt+D3RU5hrBoVKb0//5JIiTm6Txe+wViZEIBW3
wHJSa/nWTAThc8B+6PDK/ngF1sC6b2wdxRX2MaIJkj0le8sew04sDjlAvatZu7I0
xOaZigLeEpar0aUL9999ITD6HpP+E1VWkcMs+LIxyMnbY4d1VTu+YZ+OYhW0j3Tl
O50doQ0TAOdln9MX4k2aRguaJRH+euFmbW+2HfCM6/J221HuFn/z3oOCajP4xVIq
EtH3ngt10JsERRdVjJbQT4L01nJMkFCJKsNgln253XjVscez3yJMgOLyBUKbfChK
irWU+wgdpQ6C+T7r52WMX4e9ivJ723LTxcAx/zneuSeindaoXOXcfMQJZZNJiS7B
fn6OXiiwV21FGd1R6Z7jmFrkIWaX1CDJHGAcDrHWOcpkedUakxuVTliElPxOUc59
t7s2DUCo5g61OH2vWNS6Ntafb3CdQmiXHublqek0ooBy4E1J4KReQOmZBIbmbUfi
g6lp+nUTjKNPvhNlwpWyqcOMAhViQby5DzVZGp/2A00xk22MloXkpRH8oWoG7MrM
T81WKdAIQm/qrPp6Mdeu4CCfU9Nu1bowZ4QltFjphmmxsuhtYzAyi9+Drh3lhdXh
JA7OKojTThnMcwwAMRb2zNYGi6ze1OHxsOTnRMG0Sru84e43BHbJU/6wsDThv06W
NW95PTmNIXze0RLOd7BDVsfY2K+IidizvAQMAS8uMjMrFnlZAcPtFOGCZT5+/Wgb
KRm9VhMMlAWQphGyiXXZpLCf5fiAB7iCkq0RW29ik98ZZQZW+QJztRsdLyvi/Z6Y
PCKnWRWo7cgrIaquEU0HHAHzraDtKNuqhI2o7u/45TsIKtHmmJCPDcYH/t0yd0//
P/zSKHiG7wwh8AIJAr0c2ibJQLZrmrEfECwLL3wOn17VWjKXbIk/cuY293TR515M
a0XQNh8bwy63sX2vrG3sdEfJKOb2xa8HgFZkDJqv8P0kAy78bbY+jdMEiWYknWGg
DIaDzQhHf8Z3AWfyonx2J05gj4dnllk21PsOJNnh2FfGj46RI3Q0EFThhdqLsceX
IfZhnphlObpPmbEfKqKRBIoSCcFMO9Hiq1s26ojh8r9fXYaFoyprjc+9xSjAZS46
7M2DBw+svM1EJsatAy/5nB+gOh1SPTHbt6woU5xd6jRKyotwYGiSW2Dir68OSMRy
Hi5Qyrgm+2rUSOEbBvO8tpQW7OHF5rbzAC7ge5cUx22EiqGAjHAOt3GVt4S/xQ9T
77L9p+sAbbKCexxkZB5NSpKV3010izCC8k2dIus1wukN/jFIaOFOc2TuNEOXOzI0
8ubPolKnn5VdccWbMWGqCctz4Keu0sFe715bIqGivu1vDlZwz8HdibMKyaCy8rQw
IGcCK4XrwkfO7cqqgjT1iOup/E5cg7KHcndZuAkZ+8G8d/t5dgnyJNiJzPomWZgV
9kXu1umhB259UZx+SIEFLFZwA1kVR+o5Lnj20UFz6A/lYAhK4DqlqMXK7Hl9rZS0
ZoLcJFJHzQ2AY3ao2Jgo2Mm+q1N08Wv/6vJvzH+Wb8hmcl2orR1eon0i+g9a+RSv
T3g4iw8A0lKzd5lAgdavZmVmHiTUv7j7xFyZkw4uZGDyCw+PiW9Y79kbEWSb5D3A
6U/ZJL35fG3kmPzCnlRsPJFu22D0Mtl3HFmNOTSata+UjFSY5YFsz7JWZSnCCOge
vexxjkDAxsKeF9k9NJPou6+XpPANIxBQm7DbvrhxmCT8c11CKsPBwFh2OV1WqgCP
SVJtCqEOgNVHpTeAQNmdZr9CFeloWgpFRsiAILQEfGmEo82lR2+z+Y/WG5qWiO2K
TD2+w9AYyW64mmIQcu6AiLDMNhX6Ofpfqb7LsjAG8PrOBGZok+1dRqrXj7b8DeGS
mC4DTzFte6Srn62hHJdOhuAqqFRvPHRmU+RXF5i32LI4V0QEbv89WfDdbKtpuf75
99f/rI2AY2qGhZc95hso70mFBuRyKmVJXwGiswYKgh+WM/BmecEnrWsuUp1b//PS
P3tj0MskZUHwicP3pdIKF4qm0iqUL64yd5DWl71cW56dugRz+ruTqMD3ZJwTTgdL
mcR0F3Za7P7k/bnB59+l+6tgzf2vHxKxK2Kthp24sW09Es33bRItFW91cVX6xLX1
FOrREZai6xTXDzQZSbHBflG3XIKyNv9FcM3MfG8+Sbc9yYwnJVSLywx67FfV0sMT
PiaK/0lwaCnA5SLbS4M6uG1FnImDQwieLgLGVrGvwSzKYUooE9pFwC3nwKkZPSC+
hEwwmQU12FCG/l4fSi7h0iaPAD4LtvB89XiYBKjPUMo5Y8gPvQ8pf3JBMJugD5+X
Zbdo8Hb2fZ8WygQju63/yE4tcJDXSjwrK7fSLe9hdhG5QaQPz+ygOBPk2/O4+h3t
8A8RXc2sEks6EUOURPfbNHF/7u83H6r7YDnvJfhJIoUY88/7+xanqAqb2AcCqjks
TxcAo/VAX3ovOMKix5+LL3+rmgJdcwl6kF6FCizmnIb8ibGFHKi5JU7df1ahqPdJ
7R3TMQ+545SRYcgVo/PatxM1b2Si8GTp9IGis0/cqo/FN03C4uINfWLETipuPXBu
w49FmcWA2qZdb7GL8N9QPc8iWC2vtCOn2XzvPb2ps3vbccXJEqa39tzx+Zoa2yBW
fdHcfOSM0sh/LhA4eXBTGx19HGhTHzLbvpwYuiqkzzv+Hf0gXfVBMKRcID28rzUi
7pspZm+hcHCznDpCa0cEeRKyeUn3BUckNevvEfnm3pG30kA/Wk48Hqx2WztFjYfT
XP1HQX/sr0IJcxXI9SRj7FcbrhZ3KDIrF6Fr6qRA0IzdJiOlv0MdVwWddiDPIcHm
mOuxWM5C7O0+DXmnSk9y9pCI8MAiUYh/OxLZmgV4dPXKrTgyN5lzEGMv/qgbDFxT
Nyn+coF4N9Hw0l96kTD7JvGNVzOtlhq6t5PnE8NALxJyCB48shn+5CN4zMCLs4Ci
cwHN/hz5PnynHPrapFKqvQSNfvZJ5MdKbrxANgY3WFj+24UmmsXnYYL1A1VubkO4
liU2UpATvJ9q8hIcUe30cHzNyNHs7gxwef8rYNjIXWupHmHOP3nLZj8ruYAi1Khg
DBnUANuX4YZL7pJU6vReL3UtuAFBVnygNJZK+ws42P/oK8C/kmBXYcxXtPI4oHTE
+z/02eikWs1fB3PttvqGUYpxeeI/Nr4EiJVpuoIWF3NEW/J5OBF6vQhjLxJSVACw
Q8FbhBiC3Fzo4pkdZNwCDPbcKEXGhYk0OI5pDIvt9MazmkDCwQItcL7PXdADaIFE
2wS9Lzra0YxXCSKpNDvRRc0CrgxPZUFNsipcbxbv9SyoGql3bbPwyLsEvJ69t+q3
VYMElFPLxDovSyq36Gu2vSRNYq1KkjlFpwu9f01Ij0yT8zBgR5YqFwv3s4mtbsUl
clGJ7CwKo0ggsMm+qAY7Q6TcfwlGOlk+aW/JHbq5BH0maA/EKFf5GB0ze5EIApml
G89DAzAibKihBaXfzTkg48med8SIv7VzPf5gDaK8P2yrRpJKXoIBGa0YRUnU8iux
sES/f4bWpVo3xWd5lsBuilUsmlbQWcaP+Ybt6VobY9ZGk5YEsZ+I17B4yq87j6Ys
7+lzWWWHJPiODOGky8+UHREpkvp3wpZhD9pdECnPZKrT+HtnOmi2CD1UGiZYpabW
O3nzEaFQ4l/kAU3yUxudHW2PRG4GIp5V7roQMU1W4ZkekXg7L3EhOMoshjc5QmnY
Y0EtrMI+/msSL89Xw0IeV0LmrvsHCGAcn4jF05ncSqZOeoyAvWbXtg9CcC2Zgk9H
E4WVA+PWp6MTkQ32UI2klE700p/W+tyhdLqYlFMbuMFDNdxIondfZneSsemfREm9
d64S7kJjCgVUtgV/LYV8NTrI/kEHfINACITihPeB3zrB/zSLJKTAvT+sOg8FzoQz
flJDyuG4eHo5w44o98VBkP7echKEqLivMmTLVeBf8xjFq+b47FAESRUtSh/xzYr5
k4Xu7awxL0GoNCptnKx+QdSZysJIGOJLvSx5zcu62HKA7rnihz9TmlqpsUjN16mg
NIheI0cxg3OzQ8jab1rTnAKLxoYrszwzcq4gJPnhSUr40B2EWKUxdotxR+otzsta
xyTseYVTxDm8CmrxSanUpybib6BFbP6PIysrLh3SvU7SizIOWWlxjF+az2HPBxxi
NCF2ePjz1WHiNjb+nZDYB223fF7vUm3am7llQtKeI9o/I7kUxYqaJbZj7adG9gzR
wocGDyP1nDcNUsVVVNx8qQNbiyyPkf15DU+RaZBruEEuYEuvq0A9XYmbvnp626h9
7KZH4ZaVLk/uekl072wqavB4DAT0OSCQ5s4fWTBB23g3k3crSz/zQSN8fCdl7ItO
RJdneJoIE00fF0/lZ5PJd70+44FRLbnF1s1nv+f5riJiCaPwJLD/c+HGsLv0yt0S
LrIUXT8Rb8e2dRjAWFpg7FVlby3+dRqAlWLAB3cD79Q7A9s87CIXutA7mnOzPx4F
wzU9ewDyCZXFQ3c5fpM52KBIJKQ6a6GR7KuVQ3NVllisWiXWgNXwcdzm9tS8wAAX
Spdn66WtEEboPD3g1oL7Pk0jGquG0pUXkV1EIydmH4jtDo3a22cmBbIrv+M5UjWt
NkwS2R+kQI6CGwqqLY/TENk1hj0yWw7ivrWrE45cT31XGvfnWl5x2L/Lefm9ELSm
oDdkKTqwpyXLP15XqaVOP/nwJQVTYYOtqL1VfNP8bWO1jAv5TOLSaFlB8jedmVSw
m6YNtatFo7dJ7Cf57LjAM+1NtvFz4f+56g2JAFG+3yfrXRFF9b8SQ1n7geFEcyYO
2NWp/zszJa4nyIb0x2gv9Knrf5ZIGivLs/9RFicfRG2iSYByvaP7FHnqnRwmpZ/I
fOX8VLGWZDWZWx3CEAGx7JNLsnOmm+ota7iC8c+2LVHRdwH4nHlphcC4oRisbfCp
APlbUp6SjeCmWNXYzBTkBmyha0oy8PnOn8MO11S33sz3QQgMy+jS40PeC05hYtMH
Ch6noVxCPrx92JQHMVZ5eLf3QQCuDHc9N6+vuNvck7CZhj+WG60QqL69aXRfaJ0y
9TD3Ekj6EfozIV3g1y8rrvVq8UIoS1Be8LxpP75it9w1h92I4Jatb2fOHf5Y/bE4
xw0ZTp/D4FIOTHvMjJ61oOg3qUyC14Iwwcd9oddd6kSzH0gcgcIc5JizVtocSGyu
/kzqyQAhooP2Z55JYGg+Ijr0fDVGsCylLIqa1eUxUiCq35HVpp/XYcMhtO1wYVnf
vYJeXTMcgaBP9r6QHJpKPpGRooOI2XRUYTgQ9tg6CUIQ2zzjIGTGc1O5P4KeCllm
i9mI1PpUCyzLLlyW7o3FGlqt6F5ouoWG7vWAbO0uc39Q3zDJGcMYxOmaVaXS6FoN
yOQh9i0oxxaDYaSVC17RT1VpLZ3U4LSGCqPB0UWUVgMSf30wm7wFoxG4pxrMsLMi
w/s/EisqvNdwgXc8NZoKPE595d34nBZJGvs/SzStbVYmIl3tbwP9TUzC2h7J3R62
QCB0aBEWuKgRilhrNRoNLdSIqelJq0/ptgduRZNxXHWU+8mCbna0gLG0yjtUyGPB
rhDGY6g0VPy4d1R9os6L/vjawcXWU67s5UyAbLjO7VkcJ1IUo7VhXk3XwLAzKNia
6lCDK1Uec4EH/LQ1k+kBQ/J8TlQ2goOVXZkf75K9PHSpZ3IbcUEA+u0BYsQH2gw/
JDEhEfpcNgzFeq0HYYaqz4JEd5F5E2jfmHVFh/P4CgVeEQsYFXrZqVVaS+VJUHCh
3c6hKC+vRl7evRaE7407KAOOsuY3+D73EcvztwFIDFKPTVkLYxFPPxncZT0PHV23
jYlc3LCSCwGx2F348gBRSLlfSuT9XL4Nwi26AeyG6iy3E7WThhJDXBGsj6O2qb1H
cuN7gAfqqdINLOYLWRRjBepdvUY9XG+OkubWAtFMZbDf+TfBsv0M8EwMLe7d1l/A
5VMittMU5/IoYGsfFvEjHaRSJWH7icyH6z/sq657O9G+mRyr4PaSU7FI4WA1VSIQ
mYUDofxsCHgeN+2E07GMEx373ESju22I6fyyF14De7F+KoxXIFiFxxfZ1uwG4FEn
0oo7FyR/6Bb/9KxhGoWP3Hat4rmsjd6xcWrRmmqX7GxpzxIjtTay6Icw8tiJLQs+
/xTRzHhHY8l1mTZxSVBlJOlT0NWjCdGt9kas91BViDFu+UwRiBTXb8ui+O44bV5+
pG1YfvN/LwQ69GN8r/AwwGBC02gE/5+TlQGELAWw4SP6wWc6MVt+m4/j50eg+4bG
NuiNqqxwYAq9V90MdCEwKvIWBcUyZL/xUIpT1vNPmTw2sFKTDC1QDUSNhQzcqzG+
iqfan7mMitKFqoD65ZVXzCnQPVDjBpDgmjao5QTnSQGy5lsMw/rn8OxSmSCX//2G
DCVdPUPY6t/PA6CnfITHxDF/X7BrWvIvBmP6lx2v5xfijDE+97E+FNtA8K2ISZIa
Sb2q1oS27/7UbcVr2lNkgpVRhJImHmZSvZcwldUed/SWajU8YY5SVSesZ6ZVwsZB
peadKqvAyE/ofuc1j+Sll56oD4yiFpDvyH5eG3QvsAQsQihIxDWK7orksoMcXhHr
YYw0VZYPOjvkSWzZfL5YdxYW+Mjlppodhtbai9KeC0ef/YwXHAbMhOi96/O1+i2H
Asr7N8PsHszfozfMfJuARBgduPAVLqNSYYeQ3hdgRQ6pwkEUKGhQCtGU+woYDhTP
NPVHtLCWVoV/nBaC2kTr4Mlqc690aIPplylitycB9y51R7C9itpTMVVhux+Sm4YY
O2QZ4ib7IuZukk7cMpnY+oHP7SArzTi/HLBSvmtTVOhK/n/vxlriiv0lMHkfxhw6
vgb8aZy3Ic5cy5JVx9yxSiCwU+3eCc0cjs2rlrvRGVLCT6VYMycDbIYCPcAUe4ZA
VmdZ+kAP3lfxxwEKnAvDxCCiWdOMumutXfitw0liGQ2sRpFqG2ioLEY3ODwiuV6n
oGB2TAlewwQobMwq8+sZaQxoM+R0eTL6u6nPjojUq5SSwD3Jwvs+ZMfkq429R3nB
+3WDPLOBT7Jd24sTEVO58FKGM4odApahzPiR109DSXems3e2nWHdDBIS5C1AUMG7
g903iREmUV+E9HWZcdMpv6hzPcWWS6GjHSywq+N1NUkZ5hYabwfHHigMQEmr8hDo
S0I2ZeXQPeK4N4Nm14xY9sCryeQI+1r7zvuaBzIcQSo51LEBq4sua6qKoUkeah+j
fCFFMo/n7pb9KpzXfl6lPxvUpZiOQHQ5aTeGa5WxY5Xrz3vHELiQMQRDQUsxE757
OtDL1XLEFL2PKzi54lvKYxSfAl5zsByrrlE1Tlp4MFC8YLDqaiKWrbhSpA5xHwo7
ycPs1RYtOuK4SwnT/soViZy/LrHtpydhhXfyU0H3tPL/C5VxGDw7PnulTgDL9xs2
WLNhJTTelqd0+bFloZGRdBEAdyh+uHenEMVW7S0vsKiP7wUM8J3lAq4FDzUxa8FS
ny8/sAtt924jm5g5Vf9nZepWJAWo6HG+d4rXUjIOAi6W7HqZNLqbx0WFamOQThxD
tnLXjZT0LrDt+oj1x7a7A9uG/Kz4l9zwn9dD2xqmQ0nedKE/3F9JrbP6eBh99qZ1
ofoD8Cr4maLFFgECx76GL9PRdqKi9642maP1FDSc9KIwV1HCtydl20eFZJ8CUhQz
rclHBvt5V7zDOpDhulPh1qj6ruf80mD+O7A09bhIE1FJOBcZoyX918CigviJsBIF
pF3czsORkyaqx1vFZBqaPkCfdUIxFrlDzCz3rKn3FcYJ0IKThK+HrvgXRzxPiOsf
j7n+NS4JaKNGUGBwI6LTQSGkntWnJejAzXFH8rE6pWmMG8sW9q+kCNDm/mRPF477
/+jnrBdjRBrspD4poZzQZH9Z/xwUx45z89MXV4kLyCP88WVxR/CgbVjq1d/aJxXR
/WIpbPEXjvUWsT5drOSajEESCpoX9N3I4g+QBDr57ksExoA7GaGYDy6gh6RqiA9X
yojOe0v/adjD5KmrAIJB7ynLFpiQQgg87Tt8zo4xVbCh8CwhnpEhBYe2w10UEBgg
zvzerl1/grZ2EdsxQsklcDRLt/9rIeRiEed1t4/PzWHzLEfbjOEPLrhiXjFYVFWx
LzJ0RrZRQ7kzI8Lrsln+9v3f+AqB+2spiPdDIySbOevoC/IZW0+7rYiZ4Y3zgiIE
baJTzsOb+jif6d+HP0uNBjdmnvqht/FPharwQWxW511Zr+lkU9RjESHC969C3GqV
JPZmIG1SslYnnrEs7mrgBeagnA9l+3piTN5op3uN4C5CeBWU+urdN2YXhY1+oYpU
+skWr2jZadUM+0667cUyWOfHyAzZgQwcHJN4ax5kRXOzKMa7i/htoCyaE11I2iLt
FkpcX0WNF46PU7wFAZvqMZS86cVv55VTuaUgtl3m68lVBsEGp7A94XlhDRq96Kzs
oTOlLVOhIGMfpgkJTN9V2DR/c9i8sxMVrgfgrqPPD73tnNFqxVm2crswLuwyeuTm
hAP9Zb5ryXXwTsLPIsuEwjFRuZl1OZMNJ4mGuA576BuUEwD4eIQvwB9aQvxJ8zyK
Cl9BitEM2mTfoQV7kYuXH7Sed2l6ZdD1P33l73YfITnUD2JvEQcRuCZz+7e1//w3
ctV9QmfQs8X4lB1IOf3pIo+qTQwZtNm7Frn+M+xBcl30T8uW0x+RTRdfNl25jZG/
0RTBufzQs2xfArNPsHkFKL91WEyLgsob+dJZaS0q0ciL10HHYr677fYAo3LkpyQx
QRnS5L+qBiEq2XPpcmudmju3jpHEfchpKU2Lon1mW5d8PA4Uqly3/iMVX6chVI8Q
v7mGAFkd1jmkYHZihTq89X4HabWpFl2v9aIgXTfEEmZo5y/GtToc+swrRjWIJquK
TE44UVn/1lO7pLKpIg3PZM9WbUa/C4OHaDPNeN/xj7A6mSzf6qiFIbSYWcYrg44X
ifNLnJn4u2YQ4kq4/d0pZQvQlaiTnqutW2mmg9I/aZwe4HsoxmB1qwZrmebZm92y
olVfvOX8e2WTua2YF8jaPaux7okQNgt/TAfQfz2rAonjv9U/SueeRcER1AebZ6Oc
ADraidJ2ydqEsgvVxng5ERS5HodTVhNzQBkRSN/PAdi/Ww3lEczlDdJ9dpGR8zpX
riCdwk6mqGgWshJRmIfTWMHOLO9QGyxTSaGSQN1n1dGrVoMAKvHbjvexeXaICtlt
5fonUt2c31uM0mJ8t3e5NA0ZLkSmS5ccBTJmyFPAwe9okWhOxKWsv/HzrkYwYqHx
ZkPQvhkP7vty0nZ4frgTMw8hQ292Ytvl+BEz5Rw8788yhdprEpgSmvotnjvgxpel
fiEifEOuRTvEci60VzgiCJAHKD8lGOBcVPJMoDiimrLrABVQWAq0GLbtvjpagl1u
2OnGRpePn6a0F+p/A1Qyk7zI4dVq18qmp27XKRfqG1guXUWutFprJiFx2XPk8PMN
i8kApzQpTBVlOot0dtls0R+XrxWVOI3WRqkzFuVaOc1Rtb4sT1e/Olk3UDfF8+6u
karcRXolQWUKHLawrAjYt22qeBPGHwYuQ05yxohKM9tTiEdbHEpMiitUpHUggeMx
VlvyYo+xLCT9DE5f+Yk+t7zXYhXo3sByyZF1wpDZ7nVPurxnIYMym9CzDT+97W1t
Gvjo64qV8D4mgxa5qxdZU/Fqf8uVQKcXQI8dIN3FlE/C/n+UVQliIynj7a0hgsW1
2Lo6yQwM9Jc5M0KnryBdyjEEYDAOB3Pivom1HdznEeFav4sqtQZsTMX8F4K0bJSb
56KcnVwM1wP91OjgHiHr0w2x/8aVsjl1Hiv3DOIdblS5TUN+G6PVMYEvp1mcS3Ij
PNDPuFc2pIYij3iLJlk7dzGXOzsCmMmt3rO4gclqMkHsUwlBcc/tSmsKKgh26jKY
TNzA4hpmIK4xKwEhvRKQ3xh4mPBue6TZ0qZ9ZmoolX0du0YGgsIPcTLjmY7sngFo
Znal/INUlGslCAlaMeBMPCE5rupJf7JSkISvMQmaAIt3MfM+ux1WTSeQaXpgLus+
QGg0fjGRi21kTqkSIsq5xYws/qVXbDoo3PuOU7Dm4qDsgjKHq3hh8GHh/bJwr0Ki
CXrb7jlRtDI366Ejz6hF6yaeU65LoGOaFzwUYcyiv7FOy8bOKO7rjK0TVcAukY44
rdGVq6Yk1UQcgp/6//LEYrC3B5JlAvd/xxa5r1o/zjI2Jj7Ebwt4d/rRn67SnbEU
1uEOtME6qW3NYAjwSXnu2XpetpLZ27u+us/h2DiBSimvIVx0AdUOc4mO9KAsNpOu
o0nYOBZei+Ow2rAN/D+6BX6uZAzsnCrBBG8DYFidPSkdI/3lwxzKEEUkOmDzAkMl
2lHnRpSg6uCQXCc8N2Yq4oxd0Xktyg8BVWTKq7WHgH0QyOo+AJfM8rAUsisju5rD
Tgj7EiYMYquiOWMUcr8aRSNc1c/3UXWLraVseQb+h+gzL2QMCv8chck2/t+HXJkW
OMQf2To6uvIxRPb9oZvSn7DwRVrr7UKf7QPjCwuzJX/kGDAyMMAgnD05accFOli7
ZkjfQtiyx6CcKLdjUg63wWSNgPk2deJyNef97fetwxKQxyr9UvlcKzUexgS/RTIs
lYUXO6/XlP4BwATHheP2JDVv14LNgIaROG6/tD7t0H2e/Vhs/nJzmCyUv3h+L588
kkcSISJw+cg6aMdrZLtB7BxmbSSABBDTKCuLviU19vjxXgWcF41eccgx4IPsbEl8
qzjTi7Y7oeg2ZSso9NvScClg0om/ld+F5y5QqCKbYHc/P8I4+tdIg2NCSufWawgl
wHrMGWrpkzBy2pIk/XUxrVq2RK8XNXB+cSpgFHZi8JHvUdOPw0ObImtK5DV/ambs
T0IhNebUDW8/73xh3zRJZJmEDI0aW8TyrqPfLql4vBiqXHMcKotTz9RAA3GqaMLh
/ilPloRwc3WG5fb2mybMIyGiH/xVgA88jFv6KerlsEFJ2kAjoxhd/oI6gm+4yI5P
rm+MoMUncgYWd3jWA8zFHUMWmZY/b6/dkOCBsWbqS7uUP1kNJxPHqxbhQpm61xHC
v4p+noi+ZV6cl1qYCobyuBsfQZnUD9oLri/pW6F3SuZyWaqQjulNzU5fPT2F0Cnr
1vRSHtlOUuyGu+BRXs/rn7gU7y/f/AS5RIYHcH3f+SxDmY7z2pullQTt1iH9lLff
pb8VW9Nep7bW4rJ0oU8o80DcYIWjwRA7v1hn3xBHXHhFyPaxNWLVpU0AR2DOx6LY
0OwrpULgU9C4FvR4iYkeHvgEDKWBdwgA/RsoxmiOJglfQItz1Zp2551isyQ2yo9M
6hCE+TpK76PydfOkSAnYxov92xQp+QBl/RUR5OuNe1c1LYqQSFtfZ94JitRfvMGN
lhK9BR9EH2Il1kNiH/koAPlu9uGBBa3BTFYUtYr8BwJPOtpj0ZijG844icPr/S6D
N6d3KGX0FpyGepPzQwF6657+YjwsTDUVVvRIqVXPrS63UquBSlOXJ3zfB85G53Q1
5L6acmFdHgIy7HMxsdbM6qYVR2nd66crUzx0so+g587nBMkUI7zBSy5SCdAEb3y2
QL8uSOULVOnkw4we6XGMj8e+xevnOF6IWEtxRpyvkRD904hrDl0j9mh+RSGM1YJB
WMz3k6y73GQBomIjfbmVpytHMWy0xSXmDmR+R+OSptgyficrdY5ouaaYdMTmhvUd
5LGXRT6hQtpTEDmeyP5pjL/0Glm/gXCYKugPRRAmM1UIIH8LeluarPWmekBbgFVD
TKhj2Lo+EcuMVS/QvuJvyYSnMV0J9p4SXVnMyGW2Hy41dflGPxaGsi9g7jhF6Rjd
BKDshJnrSSNACQWbD5vCANpt41cwZzQJlT6YBt9cz5gGgnLBMJXeWVGagvT6kjWu
Qiqsuj9HSdyuwT+z+RleFvcJbFAu/RhNCywmAm9u9+ywU09g9BoxYyjlkhtDdAXl
aqNmf9xiQGJCd8iW/1eHlxgN455eS5aBJpQMnwTf9pdYNM2mU3lC1wFT6fFZogFw
D2xC9XAbOg6FUysBuk5kX1m0wS6DUZ5PASDgtX6bKya0sRK7VFRN/Kape3zHMZzh
6W1Rw8G+QUR6D9McZm0FA1J4o4rIaDahIERSUJ3MQsGggHFjdFldRHk5MKctzUyc
7G4wYLYCBBWjrHrAoT92v68rIoS/Sf88UrQJGGhjmwH0VTnAIEdeKpVD9Xb5/+wF
9Z/i4L06ejHJqPVgvGDrP1jHWpiICM1YFk3YIGIjinX8xad3E6j9PcHPSfsuebOi
CoSOI4g+w7EOiNwy+uVEgz7LBd0eFgUOY0AsQr4/pMrLYVlA4YjqAuIZCWJaNjmx
wqj2Xr3PW1fqhS7gg076h9PgHm9TQOr75AfymL2YZxy5wu4GXb5UeDXbM1VoPCc9
OHlKhUP94w9ulidkGd+z2vkNoP5xqFoZI0fO8grcJN1h+G9KUhTYKcpprI3XTWU0
wfskt/BU94zSoiJcjLgkMbEoXFamGPwOa8qSHQgbNOeWCHYr5u4BGhtbrYKv8qXN
XBFUgkgWwYfRAm+4HSnNue+rzcBIcWe4tGqB9lfx7ZCsS8Y94hZSFvZi/SUMLr0b
HicxX9FT5xn4N6XZ/LyZeFLbdNhO0npcI71UKQClKtzHf31LClYN5IOza+1UleSZ
LzwCPEntXln9XmINC79pXP+7224eaK0TT5CanWdQs1nYnBBSBe0sX24XAHc0uur2
qKFSoh+4r1Vide/Z6HIj9H9QJ49h9dpxvVn+LstJH0cmX+gOBhIfkQ2dCowywpeG
jNDKoGFcRGOoEouV6RJjEja5IRphF5bz6JlokvQwR8Jlp5jFNotvdsH0C+aVdOI3
lAPp/BSwOOsNX+IVvMogRPzhvEPexSDBUYHmhwDDy7mzI6E1ZsLEHZ1ooS3oKPCt
EwW4/J3BqWBqR9sIlFhd+74ZxA4ihpZWb4IYNQn3xdQsK/leuqfhLhhDB31TkVx5
qiF9wHfi7/gapkLtgQpDTXPRNj0JhFnxig8ClA+jJSu8r0cxIJTaKDlwtVoYAZqc
gNS+4gbj+Ej4P0TgeD/A7VrBnXoPzBf12NI7STSOwTrSGM67x6XzOEVEqf4cIwU3
Vxy6yZ+x3goHsntuMgt+f97UkjdT8BKYpIVb3eGyJiUh6sdboOOQoZvDgnyyFDQC
QN13fXy2EWEMmjYatPWVA5YSEY9mKfOzXbyceoh99Y8xNKOBwZjZs4EwQLJuuuS6
b3LyiwQvEFoa6UFMKrBnBCefJg8Rf+tUNSvNiCtKLa5e0hlmE4XBSvp3ZByxhptD
vT03n16603EQyia+eFGk4ii+9QCJCSZctORARAKNRxYyjz/NwElKmhR+93DwaOIY
13aOjI0xcvAB2uolJYQgSXuiZQgOOlQ+xDrStyqjPupXs1G2K2CoV4P4nwu3hON7
DOLlGhO1/tg6W+VTnTWfAAMMrD9WdHGklqp4m5/c7I3042Hu09ART0LkKrfVBNTE
foX1duRV/Rv+NTiKfV+xdHJLpMazzQgzZuuXpRwn/XJqpYxkvGBV/NWXDjQ1e6fr
6SV8R9cUJHrIYIPabcoXZQ9KKWNXcc8PBkL/2oumQuaYfLsV6ULoarFd34k4ergD
qK8qhdYKpVr4PKhppDXfLaUFy3VGCITBgzwJmAKNTqziqOmydTbBTrLZNrEdTA7V
cGi/AAch2G3/R7hLJQ6BxIhtITDPDtrf8TdgXf8PupJAiTK6jR52Q2mcExzlFrEK
BNe30JK/G5vNEUarj53Nr4a5yMdIm96Tp6AJYtcHLJbsaSoINB8aGqsZHa79NEOD
pZB0d3F/zsGVccBQa0KdKOE/kfThGFfvQO5L1d6gWNRXGJbr/fWu7PdcG2jbGxNt
+DUWAS+DLoZtpKB32ztRGeODXlK2j3cDC//XuoT71EE+WzH5KD8+m2BrjQSchhJj
GvUPxBpsE3UYki/hMQF5FV2xqX1GBE2VcRyB0yrvU4aWS4uDWMh5gfBBrZnDgPxH
24Mfnmx128T1dSmqwFg+pVYogADMm1YBEsjwVIagKh5myMDcChh1p/3vcsc3epyg
v/4PfFfse82XdbUSjcr4ReU9lfl3vL/cRbUJ2ErdfABfBoKDH0SozTLTPoIayqTO
OP3NIJYWI14eu5saKPdnIWuKymYU+YHNZxEjmYF6+05rolf5JJ+cY4zSoRkrbroW
L3WDuHux9cbh99ME73eIvfNXlKfYY842tZtxCAkq55xCoWkbzHr9fd6TxPdkBNoi
fTD14PWWvLZ/oTknDjSK8is3tNiyh+TFqVJxyxUg7sO8ABdI2UNQYKW6p9gPzpl4
JuNtyX5eh1m2ICq/COSGehqLFpjmd/RoE/vZ/xqRT0wqarDIXMlrGH8sT0+KPiRQ
Oo9IIE0sMqvVBpYRJVjhFX1xT+hSAbdP/n7ep+b0bK9j9g6WeoCeKS52Qv5ikBmG
Z/Gj75qEc76+fx0wVVaj5iRK5H4cA4Tz/Njcsrg6diRhQxzljIis5ljzCak2TzFw
i556FX06bn6yttjqDjXEFiAyfwlI8HzSBrK1st/0424CqU0c2G3EcCGqbYtHJcgj
cED15oMGJC3kAi2yl5DZhDvvOVAhkThT67vhOlzyxzLKqoQBFVAqPVdOeIQ4RZ17
8QbxCBBb8Nk6IEqlyvzmX5XF0q+ltaG3lEhDBLAM96bQS5j4scTSdcMhUNqfKtXF
juTZYodCNMAiBslwYc7RhkoLXhn/CMV9s5saXIyJyx7J8cudTocCcaVGCMDla1Fu
Avp5yhbNJjxGqliq/JpPDE5qCeQ57b13lULI52gDl76lmseTzHnyXxPz+JnjHqgS
sZj/n5XuEkPOEgzsFFe9QO+tPeh9OmGJswAKATYYEZmtAYlNqaLZnpMwQzMuQbrI
X9iTI1GSVxDgccrdAAkLVaR02M3JhOceKBAmKgyKviftEQ6gNx4F8StTKs6RUpQ7
hMLqLumqn+WeSKEPBKEWjxucb0z66Z94lRJ68xMImgMPj4tLNCAhRpWp/nYz8bce
KRDY8TFhOt3bXNfSBrIstqX+JX5NkXnfKvD0aeDPdwZa/Zdr5MojEhb0nqxDKVOW
J5IHuqsB5F1R/RSPSBppS76Z0hjzZwJLLIYn6l0EVTnPSYHmZQatfjjC2fGKGPxQ
KBJ5NoOxeKfauCkHw01HFNI8PmgImmzFYhU9ZJ0s6sSVa1IYqYw0J3V0t+1kyOyv
mppaZfJItS5e32GgU48v0kfUyjaU1HHrdbPh2Z+LRSYDvzuNioO5c75hxNLbNTGn
R/ulbXuwVn3lAYln38P8FLcUph6myJpkTMmi+NvKQO+Htrzf28A4/UAEt29Oz7Pb
BR58xAXIaYn++Agx+W2gYZpRwPWNoG6YbVEMQq1vF/tFaTCntSBt6xjRHeO4Dmb+
Q4kdZtvDSyD0KqkX+Dt+leHpYMxX3T4kv1MTxMI3YlqnAo0oqq+TnFwZj7iRiOtp
YVUw3WXWMH+H/Olllidm3mJDqoF9dAaME/K7MqQvnDQcpEqcR+LfEnIl7cmUstXJ
2nYN1rU8XZnsJ0orB4aT+cck7rtiQ2fvnp+6tIsdAVSS0N8w/g3UcIpTI6+L2Re8
KfAg8htIb3YHT9cpigxNJB0QUQNhf7n0lv2ELzian9SdgEXU5gU4K+NeLz/prJzL
G5j8RJN939uxWxc/UQZVnCsM1gvNN/EWWesmXDygOC/zAdtWxemmFtjbK5//TZt5
WkzNilhy54PWQaw2VQDr8LjD5RVDn1yIL0DxIFhLiJcVznuH6p2SOBQjotVsDbre
MFjObFLxKPi/x5OoqbP4M/S8bavEtmA3j5VT22utaM2tuKrtaj41tyzcQR5WQWs3
JZwXnnmV+3vpMUL6EssBv9OaBpQjRAy2iZCkUmWBBsyaFHbfP7eeWTzaIqZq4WSi
+ppnCThEoYsuCF+eVmAJUcy1bK0WABhsrd++7OPl2YLeq+Bat5NeRIAKOCrtb2O0
hBW4UNcEBr7hFfuXQ7/09M6uw+7DqSKLcFlSM94n2JkK6T8FIWpGqpxfm0Ns6MHT
7spmZ4QKAMayzDKvPLy/FnJsp32cP7RvR7iMcIQrHG2u3/J7WJsWfMDG1ui3I1Fq
XQEfUQ0u2DFWAp21LB3Zq1mhXtN7sfi+JMIPnONZdLGk9Aj0wb73ahEXRwg43lU7
u2ddL4nWleVvnJqo0t55hRrS0rudM3t50VpGjjQETf52EP0g3GXkybVPO4KC8o4k
WKgtI8BJyvcbmSfjOeFb9xqPlPZE9abkA+KcyLDxUH4HRF7u5a6mc99tGip3Q6RO
YK7MmRVf8qnVjFJDtqkp59fIBLVya5zKH+vgrT82EK0lQXTAIz5eBIIUqeCQFPkA
GfpGt9zC4GUjR7d8uG0cG7x+PbdGVzmJz1/g1lg6J397YXJOhaI+waujdS3iOFQo
9Cw0QyKQaVBxcNeIRGSOQiHX2dPApzNjAk0GdZ6iGfvVxgMOgdKsa81DF09Ew9iF
WNk1saZ1xgNe1KZrEm0/31QDfWRNmL0vrOKzhOunnm1nJLwTxa1Qf7CMbSFXhtuU
C/CTHUvHc0fj/OHOmUEkr4Xw/PHdM9wG+0m9xLvZWLGJ9vwARLujuTO0UD6BL2Mh
kJaBYduv7OX/v3/Suf1m5Q2qATr/o6paj8N2u1sGyXU1ud8a9dpZ/if7XpFgP9aY
ACRG8Yy6a+GMAzpMUP5wUfFH1vhtX8YmSL7oR/S9bj5SUAbuoUGMp+OUaDYkohW5
rPNmHrDYZVm8PE/KWopxHJnInidZK6LAVo3j1UcF86NjiJVGqDKri9jJPqiELlUr
nm/2v+4TyrfcMr2m8UPJ1O8ceLtLIZktue9rz6AAWMQgLpzSPaVDvtwMeFyqAshD
0dRKnYKboOC8t5zf8ijm2HGa7uDD5uzDDWeluy7fOreHkiAGhEDXr14f7MZesw8r
q2Dv9z+25kp8LWHbI54e1825FZ7Pk8N7An0JOquTPExFDvu+yxQQIArtAM8nxXrz
n3nGZ3W19H4dZOswY50fcP37iqo3yBFkAn1qSTyMRXLmpn7m03UOSdXeafdRuNZQ
Z0DnLrQAjxUgbLl+s45wz3a+rJJ/2yJDPGyGBQrSNYg9/pUGbqroAvRSC03qS5fx
DeSQHYzP9TbEj4tKQEH3PaJL/S4pqaXKasAwujpn5ezGtf1GElevSH/Lvdpzft7Z
xB6ee9AkGE27tIcg/6kfmeBu7jLd2Mgw3yP+Y6BznSSM51+u3ykspyF2sUTWWH9w
dm/UxK+b5hQ0tydlmM4Aug9KwS3ZzS//2/HHfgHv+MLS8BtfmS0bAH/So/AGIFY4
hgRLwxVbAB1kkR20n8kf/YIbrlbISsxns0I5GB7hggm7gOw4zjCsMa/iTOv+7KMa
Wc/mJoFjgi3HLVzjCsyNRSFOuCZI8DDXim6Qw7YDuJG3gpMrvozW9XdIyRQbTBnS
EJfpwFzdSYglBiNhxHDQwQeY6Podu/vE9VyfiTLnPB1qwEQBTSdT2gCxmkWDdxI9
xEYauCHwwYkAKmACTNCuRiWXBd62jzHh+Sa1tC+qhedE+v/wMyMJQtmH7UHdOpF1
S9SFQsba1Kazr0xcs65bV14zrprYaFpP/XwDg6PYq3rySQvNgHvL/Ec0oGlXWWx7
q1eeKupetd4lBh0fjQUrkv6NZ+q6mqtnmI4Yvsbdrcc+NDbXsnZajZD2vTRSWR3Q
9SHCbPq4/PhKBgZj1a4KFfthRnLODawnZz0L48TSROc3TPFZGexb5CBJ3IO3vLuZ
TFrv7IRMBvLv4aEDYEdL67/F9VhTDVptRCmg9ubtKoSz3Oo5D0V5pF8ADTcJK4g9
+lTKd1kse6Hluhtblw79jcgYW1E0IUMu3c5VKl0ckTl2iFeV5Q4nheqcDK9U+1YN
01A2zWEjxYbIHxWEgOa9n95fiCpYNfsOTXwgk2nrsvvN1c1CGMf8imAxauqnhs6P
Is0zyxtdeL+L3mtkx5GTWqF9LZGekgq4545jNGqtMrA5Zuuh58jkgkGOFECiUKt/
dXh2CmJyJl6kEcA6jJlO4Xk9ji/0AcJRDWJgshtw9XEfqEl3kEvBYMCb6n+RkbER
m2ZDgCmGznlqno3joIm/jaKcwmG+Ov1JUp6NLIFMfY9FjdWbvI+3nv0NtHPY3dJC
vDRKC75SGUEgGyA1zPwrbpue9CnqdS/kznBMpiYAUXvhdVVSAJ5h+4y4Y4xgRcO3
V6SFNRzRYXdvm3TYdZb/LwJ/uLbSxxfPYrMe3zX5j2cBO9EYebLQMYwjOMZurnjQ
ovIGbxaCTVDwi4XA+I5pf1fksE46kSBIpGAFZwG83fwgAbJpJNQu1OjuxCzttTNm
PmO1DzPMTUK8zFBk1h9fXc2MZTa5+OG8l0jfrARqDwCC3e7TB2Zaysc/dyIXsGGh
BDgbgEJNxwOdIKL4wHC/EB430JPWiaHJLCU5xOQUitWy5I8ijGezfIQHDX6Ds207
P+7ro8o/tLRbjtt1cVD+OCz/EpP3B1JoMmUhLHxarreUjIHT//vxH73CreMD3YcN
csJ9kJAmzVNGF+qZDGr/6/Moffz3tZO3dmqL9k3pjdCxmfPNt6uAMiQXsH2vea0A
Yj03WutQvjK9EsySJZ4qtUzk2ifFRvH4jG37RrYmyY4Erq24H0g5bEvFIUjVoMps
M8UzzKpbWQpXxv2sSmZ6+5emQcTu9YZZlBHzmI706VYl/fdxZz/K+UFME8QY9/pp
cHh5LGGuBRQiH1ykHpX/D0yh/bOgnYYHfuTASfmCoaJqL6VQmYXWRdGFYfWnOizO
GHKPqweDhFp26ki4Ph7iiGhOlTl8oW8yCcfzTMDZe9So7IPzV5NcdCs1g2CWgahm
ljcUHZxro1EDOGxRrVViy5IC/jCA9WyE1k15FmxatWcGHNm51cIpyYXd+vcYtHyh
mhvdjkjUbvvVgrTjzg4rt15u5PGc9BRn1b+qEMtO2TduGIgQ4t/lFknLlFoeLQKR
FXPDH8UkDihk0Jdi2Tx/esRSImXhUt3aDRiO3y24aZCXtLlkyGYpBU6BY0g3iLiE
0OJaehCyeltXqeyV2tn39LC37J+Tpr8rSeCnjM31HA49Ze8xA8InETdbzYkJwPXt
cD6XXYDeZjcvE4sb8dQTg50RtCAzq8oOZrumC/Yin9B3H+Kb/+4fH7Kmy/VbNax4
0NVrYKCc9ZMQmtNY3qLOBjXMfyDeaHuyRS9ib3ueMxtBdq5yksR4f6AzaCHc6Rk5
u8X6J2Nq8aof3R7qJ82PnMnYtOS/NAk+voxl7704CrNOira/1HDJ9XqEBden6YST
o/p/R501BcOLDeO3AkNAVOqv1H8UZVPCoWyN5yyki2rTwS0f12gfNfRVLGJPrsl0
q8SLeXN2PXypyeiGL42wSDDo9drgndoAYxAh6OqFKAt9+CDgmva0yHd2QIXd0ty+
SA6n7bO2eWlnBkdSGeDbuXdJijmqjvJokox5wDNPX3i7o3kll5rCm77e83PuHTQl
8GZ+ec3GQACLJz4PBA7z66R/KJu+9NW7+YajJKnWXxcAFoQS/+yYF66+ies5csie
uSqgw8fkhjJ3Z4R5fNboDy0ah1EvhflK2ArEaQka8RtM4DB/C6l1mYi1rSRdBJUG
7Nmd6BqiDXoxASMnVtujT1oCw7MZ2r7NmoPzhGRLp7k3cfRZkNpjd1Kdi3UbP3Pq
1DEC8peEQOpG0VqME7Jji7XdV/lKZIZo2eiP7QLprRJDj9KpsKXwMFTFhBsI3isQ
q2DOIKR8j+WliDdhwYqltIRAMMRy2MuVIvjd1sYua05P5lZH0N7DYBKQfqvowLXM
FONjTuzW35oVlkNTvJ5sbJgX8hIeKxtGf/sSJDHPkZ+jWFccisUuUehZ+nxnPcPG
3emaQbcSStSl0t2yX1sOt6bOmmoxsdIGdZQhX3i9O/J3ykqdlJc7JW1fmzXaHqMc
/xUIP4KgPqoC940O79ASTvazvJHL0vHScFTSPapIDpGcljVrmCbcPMFdi9Q84+lV
nQJSQJJ82BUfMHikYfDeawYTYntE9Hzd04lwsvV5GNd005LJ6mpCR03k0/3l+t1T
0LgaoeKNCJFXcAu5P8Rx7HfP/HvSKTf/oKzIK6zjp79PS83ssl+/2dAX3ItQJHLv
XA2IhaVdnwoO8k7BPt1Z+JS4Si2KnMC4bV9p1mJbEjDIWLkpR23kS56wRGZjAFLV
6T9ieJ7ib9aTF8GSJfx12towTy4+rTd6/yjS2fsMnDDVT6wcmXYbhyBx7GeudLpc
RyIWBgke8Bxnepq2ReCqhU84aJZIJuuDC1Pvy1YynBT4J+C/V4UyyJj4AulDsSSp
QQHpVUBkTOfUjd9WQoe6BYhryuvYbnWXeR3dssys59Xhfc6lftfToIhqRI+xH2k/
dLt+qI+D6i/zNf7+hAri8UYJdGE6nLGyGl4sVhsujyxO3YgzaekDhnwCA/df3f6w
bbJ9w58PSMl6Vy/2EWy2kFxxoWeFbn7LwSK5ezvYtFuioucCt6oogzPSF5m2McHS
F5HBGMqCf5M8o8yFz4lLE0M9qg0QofQN2dCqQDtARXY9/ivgkFMy4H3OkZw/k7Wr
P0URytWU+jUqQMX7BXXEi1wrQXD3FjV+nBZF7/8AJ9DRTSDPSIbBAZmPhhDftUxg
dFb6HOb3U6MuBitPk0lC6qj7iESS17wb6PqTf0sY4rXSPWOToVfezR5mWpexXEyC
jlXPRf6+dm1Kz14hiPGn4f/BAMwq8UJHq9xjroRfbjcC8cUKhGhrLUjeRXtpi81Y
J+U5ZjWk3sW2atY2X6E4y9seq2a4INphj/sGGN6sc3doq24UIM5m7dxDNnLVwLXf
lcmAIrU+RH+ilE3aZ1SGxzhJdM9yJFnzZU1O7VVfck8IFuSRdJlrgye02vkT9x9G
dQ4BEJqwE+6iKoNQwKUi0ix3gGudlTTDG3lGyHnKtmP6NFKewDfxzLTspedOzsSg
S0Y6a++wXZJXsFs/ZFsZofxX0yg1RK0GYkZ1GBDKPhBvSJvzJuBlVW1TiKpKXF0l
dINEf4wWGctMsg6Q+kRUG/86Qy3TlwK/2+9yBgXmnPkfy1M7Od3PhlaaXjknkQII
PNaiRsGAHu5qtuZ7r7tQLVgtWFimVS4nETmpYz4i210S3RyPOz6eXH2ICDLH1PQh
je+iaNdM1Zmath4P6vwXyVADs7/QmtZQgxbM3yUeohui8ha78QM4fOTV3lgTuW2l
GDOVshfMLz6t1wcE2he99hNh9fTJ9cgSPIXx3Cr+V6CAkavS0dqlLTWq4ydBUv0w
L4iHTnMkwfA9Pll3rAdWKNxBSWFkkWHE0HKtM5oHSp9+/+MQdjv2DpnpIIVPvko+
rLOI4v701uu/jIz2qbSResKQYYcBR4Qcg0JvQRUgBg9FLF6xjVq0EHr6/uRPd9bZ
nQ+mWIdMiUzr8Tp65Pa/pYCEyUwZzvqpvkkLLSACOkOiiUbNeUJqkuMRT0Pbo1Kd
BGQQH+3jKSzmS2c7xx1IYd8uSqId4R8cRq9GZTj/dRSjuEihp1wIA2pzuR1GiCTH
L67VR/bgwGlaKN057a2uWhNWT0bs9g6jPDR/eXSehObp7c8eZjX9kUodd2d4c0le
qquiHskjGFK+4/5oo4w+QBcpi0wd6eSg4GXzEju9Divaab6+YRuhL11eACu5Fep7
RIzGXGhG0ZSivkETn0u7ajaEeta18zBlQmARxFM1y3bBaHVtO9W/3HBY8LEGfbhm
WGRWZg/Khtfmj8pgcM+JS+8gDO9C0epYt94n4HtICbPgSQJotv87j16f4DoB960h
5ssfEv+exWL+NsIQ6ovkAAbZwKbM39Pf/Ko/PRBEYlUh/HtusEEGrMJtHNVbNz1p
RM3a8h4JQFCnQj3mL8dJtll6wIcryptObINYrYz3kEvX8kBzie0HiDx193M+2Bpn
gBK5ySJpEh4aRPrBZa8lM+ASeAm6oXr1y/WlfB7PcyGbvmhcRHrgaSey9KajYIA8
T0mg1QL9QLcgxTZqcL7zbafqjzcUVRNlPIEPr+ZYGR60qtHp5wiq4Jib/W+KK8sW
QMDHoZmaaRXGEBF1lXoyum6CRm3PqinpgWQtv12BXT78bNB0T399/lHkfTCdwxLL
cgqHXlmmKNV4CJxURBkVF6XInX0AUs4PuzEKYGV1vm6Mg+J5pVKeujXJHu48Nf6C
lEt9/U5xRaVYYSuKmGezPowCg5LMJMt3X10hnb4+iStWmAeXc3aYJ8sY8dmeqis3
BPkuYZ/Hvvv9MPsbyo5YRbDPOe1UG5nUD2iVbEpkJiFPtexLZulPXoIWqcBK/MHY
ynpG5LDtgmMQuIGpQL3ADSOFHHra2ZT8PLEa294+9kma2zQ5xQ9dniuORTBLlTUQ
XeItcojzqOzkoUrZybPf92SLYMoQ+fg5adgXuPiA6t2aYdwD3WZugbWlinJ/OiiI
2MY/8oB9GA9epRUnz5uf0+lZ6RvcQMxqG3i+9yPncTcc46163RGXuyCJXRgeQWi0
6gjhYssdrm5fwMRoDuCAdPvdwfF6D/ESzNGXHT0IWB+HZtUjqLDXxEAAkPBUeh//
8eBp3qv+mAJdjIXfqFIo0R4TljizBY+GiohblHKAKiK1ZpHUWP+qpOJG6j2JTVnR
9m6fnb+3xpR5avgC0BTMVAtHZlNsblH+tQCNDu0rJyfVodwP5UjU07TBiTLLAb9p
tUAi0EZPAYEv+EUBQ4w8+GC2xPwszMd7QLcmtE5Bc/y4qY4ARmD45ujFdtnA3orV
aMGbq1bb0GpcEa06Xgb9T26lvf0HcV/HayTViZV8cezIF2bLhhlciMpM3wkc3p+L
BJkkrU13gzblotfYO6QQaoHaCRVSydGKqhdCdz14zvh05C3fDQqYCYuSMsMLI8Ac
W0ljivquvf9cqcVqONwnDEuxWTjLYhV7rhbdA8VKbVZ50SpwJRLeY+QN9VL5VXq2
7ZRmYs1lfZEOhVcFGzuAEbgPmTZwU071P67t9g0NLDPNMR7JOsYiJWIgZnoB+l0u
jkwHY0kuiT9w6MznYaCBxIKo2Kty2mLAEJwULU2Av22uTht1ahp5miM+RWzBfL0p
obLWxFB+eX8KbbVeHPYsnhxe4HokdvReJr4BTHevHSdhshspLDWam05yR7geIX7G
FEkZjxcIaCBeR+0zGWjFASR/PboNFBdpKxSUo1NFIv5HtewmQCmJ10zxanYRK8kA
jGzUnb8wFuKuTDNlKuXosHKD+SA6rRSoJMp0tH2g9QxgFX7HdNvsCXR/i/baIkOV
5K62uTFAPAQ6tfPSV/AfaRr9KemgRkxr0VpiioBKnaGFjMJVdNd+puks3HhMD90i
OArajWEodor9wE7p1KOyFNTt5YH+xkLEMTAEvd3bZF+SRG0RpYi3NhOtXUNsLnJe
W1gEcBdBTvhKsfvxMMlvV7YbUk8tJCUvxUf/B7hNWrn25riZms8yelCk86nfOADa
KeYhnqJUZPG7rAQLVdngc+t3rYpYt24ZLlHlc+w0nRwywY7m2dt8Z2RcU0yxkDFd
Gu/yzI+nMTyulnvZOuMN77B13SUg4GRS5bpRdH46CGsiN+mlHdGGNSjynDjiznPC
nNolWRLzbOAPiIoTrrAvK9ZyTeSxikX387SdgRbnLJSOL2kpIiyM1B/L5vv7dDIx
vCA+Y71qPDH4twoN6JJBCL20Fgfu2MShQ1Y856bVlHxAGVZ/YJcMFShbcLRHoDNG
sitDSNaTtBZf2WoN6a+jidebg/xZYFoLz6HNk0BY3N1fHQnljKEnc7aZqG7w+c7G
p6DlvKmhGSjd8RP1mmLoXjhWlYXUjgUvnTo/PYETQMiPaKje4Rf+UsNityiYCXt1
qxcE3C3Z92vOSigUNb2PnlEPGbAq/9WN3HG2XlXBMbukK8f1hr+LaVMhQ1H6/n9U
b18IZtbKoluBUidb5sS8rWi+8Z3ZFULCP09pm9bd0ijt0J9m8DpPZXEE17Y14kVQ
gEloSWpNKzlsTlvym7keMqEiTCYosZaGfJk/nS/lrN6iZYuBf5aghQDY8BdStnV9
+98PFRue4IzePF2HNDALCixQ/99LHQWemXGVmONyDeEqhaaAdTAalIVOOGdYFniy
w1vmhl+3vx0+QOhGJ54WNCnh/IomFvNoQLax75WJ8WlgCG9IXYU0LoTHxqTXmazd
s+PhhCZymtq8xCgy12T4OK9ZL7TUkvAmZ/Sbzb0/QhGg5odNQWr6FnRZzIQZjJf6
CQroRXl6ULZ+ekwwy4lLb0CK/vjjr02FmutG5u5A/rf7G24JCe2isnNYkCVaCM91
4azCwdAfOH/gYYQ9IChdji9QjELxUzKvA6z3mVtVmRRhHHX+e4n55C1tinDPC/U6
LtQhyns4aqN9sS19VcSKY9jCWG4eZdqtPRxdIMIy2b4DM6vHUyz5EENUfZ54sseZ
kNQmZ31OTPHJB7C6n5v07oiOa1fZLYQS/auxIetP+kMZNv5iMHX+lCHMbs3AiWmZ
FRWSLzHjYRQl9oCKltrDFf/9lYcRrvBmcCGFXZh5c7xSutdTf9C9pNRiHdY39qAx
BjEy6D3JLifCSp4dB+0B+sqrouwZxojvMZPJ+xS5WFByH4WO1KwaNsqexM2TF/fM
rDAnmQgNPZ3yNtl6tMVSvdMlht2TMLs1G/wz5YeHi5IYozORAIc4mp6he3wkNmYi
SIUF5WjNPC3FPBapU/vuIr8fRPikboRjwvsBXD+VG3GCEcfkU41NaOgOENfgfDiV
bxRcRCWYumGk4k43Y29CWL7cOU6tCMF8vf0aj+a8ptjTmpZ4TAIdWN9MPGfyOnjT
WAz3w5RDXD6u4iRa2Xdla+UKdpLet+70U9xEHR9U2FJA9erVW+sgR07AoSXsjkKn
CzthOVHWGNhWBPbJ2NqGedsjVqyP+kVISmup3u36ylmAtoIgL633tdy39mJFcyk1
npakkjn+SEnp87UBjzF2uovXuDzQnlfVApg04H/N5JCrj4Y5kwuq2EYB0L98gK7C
vMOzS/G9i2rNY+STW3waJDYWcplp2SClcrryUmVkKA8USrEzzVmD/QEntS90LKaf
FhPgJDXjmbhqYS8sKqGCqQ5DZHPMVhSvLGhyLYAFcv0OUwF4JZcremhPtCQo3PXq
+j7D4LLIUbiPyEblXO4V3MnMtW2K6wPUhBdUlt3dTeinvMvIZSmKazsKc/WJPoeN
xKGipOSJ39SeRx5PI3yBYBCo0mcadL4M0X7LRwhn7MW0PFuT1lcNraG1wdXAiEv+
xWmLlLqSn0vljOBUVT82OtelOoeiTxOVanG0/2bRFYwL7qaB0WdgdESWjC0r+stz
qKY4JRmISw5G/MRO82IOIHCQAhwSDpGEYRcRYJ+laKqXc0ACBegLqbxLMqsRNsmu
lXoSEN8r5vzEi2I/c5uQ8aug4eLH7a5kuqP/R15PQeT/NibeEh3tgBOGxe2F1mE3
UZTPJPT7/Lbr1oiwmCk53kPPc9G5OOi9H/pt+ycodDqJd0hwZEmREty5U54iDlsN
pTYW0VUSD3nnkaV4hVYftxCzWKr564EEBUPr5a3eyeQXE4N6bCJy/RviUzR3Dp5e
XTaoheYcHLDB8Wq2duZxlSwQ9FiVrKsPIdfrbZy+Qofgpd47lW+Qq+y5NT7nyI9C
zp4zx3cQUASB2UfcbnXt8+uKSIwDpQRpaDEq1EvXXG5splI4mm0bRKEdyKWmJNAX
7ApAv5Ne/q74NXrCYYRUgZ0qwgdiKIoxkJ9YhDVBoNXyg6uqmoGOn+QUiouiwt+t
tn0chrLOVOJEUk6i1QC2yq3Nm1KVBxIk6lMe4AS16OWfDrhyHvHzymMhTZXhN9gL
+Wam52anC3hIRNN8b/ltzvGHj+/3lakXOE3NqDjpdHB8J1oZXIQUYFrcpeStQiDf
DnA/1+7RctIfPV10zeg4fRHcuJuLoFzL4TpdvnN4PyImh0pjcBHIlQ55BZm0th4C
hCedw5wosIIvGTBQl5SdZANY/TCTOyqXqi4TrX/Knv5HIF5DkjbXLcSoopKaziHV
mFXQOtAujwGRWKupehdQuz9QwI3OisqLY96MfCCv+Pz2lEt2fwp4YyRst2uuOQTp
PMZVocvzGt0AEaFSG40qAdNcUhe8sfZa4EUYZ2LLMUqi1RpraHjVUOuQAKHijUIE
UGtdcpeEwqD5biyvPaXXG720yjxwqrRTE3MJwZL5qByW/HpmuZySaRmYHRCwLZfi
p/WTQzuaVgO3HvFiH5qHoJVs+t7g+jHNUG7PnQKAghtyyXNE4GYgoWEBb+9Q46DR
ImjbnkIwYKkrqQcM14Z9NMq8eMANcnQTfMh8n9f1vbq4ETUEhEcWbi4OnjTqkoo/
FTy87O+Cg+S5cTAMlvggKYdwdnTcyLZYDbBIhGH5EZ4bitTSO0OKxk5Joha2+hD2
HANUDHG1UXPWLv9sm3JMOLBtPw2it5MnwQJD76SXFZOXN8lO9/Qwz1+vNHFyfcvH
kmWTAZ7fuF72K3kl36FQuEBHuEVRIZ8W6KPWgdcozfFtnbq351gjZQ3JDuZzdlnq
J1xxs2d+XqAMG5VhBgxohvSgy/8vG6FjWs0f7/Dbuikrzt2rHEhH294MaJumNHJQ
3ZYjKE/ShJVs5bbcgjHzAW50ac2a2sV+yC+VMeSQSmODx5AProu1YF6IDTLKg0rh
868aTc18nsNnfyvQ20h21tJsPNr0kCkQNUu87LgVRj2hKTu0/eDuHtVfcPmb+4TZ
8xhFBrD9KC2kmZuC0y22i6vvez8Ygo9ZAaeRv+3CrRUCkq68HX5fPEVSz9nA++CS
vVzhNzJwV7jUDZNqPizoHjgl01p27oO1DIo1FsmIBvfe6axkV9Z301kn8Pg5pKcl
ZuyX95dBILMrGNBSskQWnj+IZCt0tfp4q7qs6UMpg9tVgZMCoN8E/g7B7Qz/E9Ag
Gwom0FLFjtenkc49e2orHw+XryJ1gBdGNnlCZjP/ygLBvXcCtO61K7QrHv1CLRFZ
wRKOdD1AX/6bKxjXIsxi6uVrk+zztmfkIEwq5mKBpF6Ysz0I7+Gr97mgY5QH6W45
Q8hP205N5AIBRFD6Qkzd1qFKeeWhRKkmuFC6LzwY9Aadwqn8lVxy+PwSbSyVyMyE
cNyAF7X5JumO9I4StVWiGzERI9f2Jzv7Ga4SYuw9n6MsnFKE5MXhUbQLABuIhtLO
jgruSkHDMjK2cnTQOrZRzBHw1TVwUL74KWalISXKf6P9AxpcIct5b+LPwRasrOY3
IQTvbBXUxoXorZSyNUbS0wes8VbSuSIm14iftnNzr9FeFpih+H5t3h8UNtCyVuOm
MnW7pKTaquYuEAVX7zGXz0qnJJg2pVdYBRZI/FvZfw8nkHWLfFZpVYtFyCOT/F+h
y8G11RVbLTYZLmmyTnz42mzOeq8p91Fz0kB02PgrjdCfIpjDOZCYXqi+3WOmrejM
5d0Kzbqxuin81ty2dzvD4Z7Rmrz8qpCsXL45OY256+awVMDUicTvFiTGzeL68FPt
+QKHbTiSvJ0wb1di1T+L4SfTEyU/clerS8A16dyCGsJx0I7WBaUaSF3lKAYOKInO
epXGN9bYWXxciI9zG7kAKAcYC7bLgwgVhPEoij3KUJd8tjLDY57ajBswsEawxUeQ
A2B4ToXjQNItpwtO5QHJqB++RLbsLoG4GX70td4mdQO4U6j2FsY6lE+pPuyfi2XO
vqAB9isyCutpU2m7aj01KKQCFbALETKxiwlWRqmcWv62jEbuBy71POzPkgUuDRVW
bGxSKMVzPrbP9/92mvCS2MPlpvIzFrDNQ80BTIM/HcKaxiaI/gCfWyUwlxWkn9Gk
TDX2w1bxqqv6Zs4xy1NKHC0cek4FLTkktSNb/YqWYh/khmLs7CxJys6uYNuEJR3r
zvtLBWj/dznKDdxXYhsKHRt98PPQS+lcjpE9nmKejMpcU3SAr5+KtSDQWHVq32TI
ynjbotQoi5A4bq79sjEQl4Smb9FRL0EgwHp2syJgJIusJfwDMNaYd0/JG3bdc2JY
750eHGXQVOviwmEDpCofx98CdJklZqGXQ0iv+bVYrJ3dB8BUFVVzZTj2GJ3jrpmZ
edCRe2BvkeW+ClIDX4r63lVbaGbjboYWtrrCo/LIYjskznawm0Q0XmftlHaMQA09
M62QaAzdqhEpoum+6W2LAd8gYstvrMYX+LH1uxDifwtdU9hJR9Lj9bTGTnmTg6wO
BLf9ubtuTaNlq/G3yFIMOkkt3cul6rlo8Nk41Lp27NczkyM2vW5hgz4uHBiXa+Gw
v7Lo/9WS9jILv5H68zv0ExDKRoCDU3lDKHJWocHYTnNfGVw3lWskD2tWQ3vYC6Gy
wcxldx848c+HSpTSXFEGA4yOsv9AbASFuQkAvd/ATreLsf9jSYsB6TRrfpOzmEWv
WvmBSKrIJsxV6OPnIG1gbcx/cjWLSA01m/qvOg0mHS26rU35AG+t0ZSwyMAMIcK3
1/E6Ao4H47Gj68mNUt7Am3xRjzo01eOlP7eTX2rZY9TM1IJr5y77ReIu+ade4s+n
hQosDsCLg6DjgdVh/9CzFKQzKJDOBPwZDGDqTVgyU+Sa147+bzqApEAWig9kT5N5
ic1qaR/i/FLe0v3+cUiQow6ElfLkaIj29fTU7FdwDaEdN1ajcQh+33f5AoyRBGjh
2vOCe51yR9YC29gSCtmwY5qqNdXZij39qgRubG8zJ2oIsEOnTjnCxGVDHfpBT9yM
I+tlMlkOwRzr4DrYRzybDmvdi3mcOQZeInxgDzw0GeuG2mDXMLImi5lGh0FULCAa
jiTpwcZJjyZrkGMVYeSof3Ho+bD3nzg0Z2mmvgynNV5DZynf4t+BefnkpAw4zirV
FldwL5ofFTBvDkbWGIc2VLXugpDdzhDthzsvdMzvJKJRYYyLj4MD6pBRemMvDr1q
bcURI4x7tondzzcknKu3zEdA5Vbo659nCqL+XSujqIVkQyVL55j9yNJFDacz39a0
9liV9nZTGLAZVYxgyTYGlEndewP5vb7StyEXWV8rsIER6qPTYFJaa9SSQMc/Oh2t
ftMe6oQLIB4+u+2QR6oC+DULNp+jx9L9FmSH4WeINT2co+zvjRcD3C9Ij9qks1ci
2kEYfEN7EtpuL4YU8zYm8AMoF0TjQ5Xqqw359t/PFdJfljFpzzTewjjBNIQsJFIV
NAsA6mAqxoLYluX8anb3jUOAyvIvL3eA4IllszzKYPXWIpAeDoUPa6B8JEVUONmL
2MtmFlX4IcnZbpdPWcJXOTCe7szd9hq2zvbr0FyRfP7tMbVoihiUOQm6UREPQHMn
J1TOuNkhfr3bn40PNQx721xkDuvwgoNmN/JqH5Rn/dMFQXfZA+59xm+N2wwi5oIe
y62LslLZOhqgbs7YFgrFDmYIg2QK10zpl0HT7E+ypjDUxxTkmWlmNYaGu927WScK
XdO1lVDdndKaBDmx+RqaBcix91zY3nqCRSqFXj78DlEP0WIapqw37l04c5GPS/g1
DJEQNvtni7IlmlKKGKX/Jj9R0rMU58TcFYnKqouwimRZQrKcvWM6ONVnpmdX8Kwh
t8WygqROZLYWkX+gCDTLjve4f5BgAo6feNi7B5D4thx+Ekewgp3OJjNlc6ibNIkj
+ZmBjQyffqOd/sUcZ6n0jf8pZkmccL5iVZNXI34m9B7ER/l36MMqHvb/GiF9dGQ3
W9xqM/s7N/ylXe6Jo0Xsm2Rs/XRvZ5F5bZFTDMGxJVPcKzkOf8ino3DcH6ORld8A
1Qw0VRJQ1GwezSFJJb8YR6j94QML1+LrU8yihoPJAqnzovB3CV8MJCBAoUXgSc78
VQ9OLVR/ZhNo5qNwfcxX17SMB96fh/FObdJLVMy8kc3xBchCvG+MQLCU7WKhlWO7
ZsNrW0PR0ESUvEcz4uNr3bFNkljyrMIyhhsN2P4KyZpkkaXm3drXcqvXFRC9ONC0
J+rIzPoBIeptMPN/pft/tHOzV9Jg3FTkOlwqvcLsI5XngLq7JhuwhqOlilPFSw5Q
wiOve8uDRU0xUl32C830kSmQaanEc8rofJ1xi6d5mIQGQOAcoykdhWJEaqcm/7d7
NUk/fAOgMFjVtoVSr5fMDQDKcH4LpNlQIe6Oew8b7CytoOnnXx5iaLQj4ECsE4vJ
riE/3tPZKozLB3XzmK855GMYCqWKAct5EfCVSb0V9cIozm1cEYeHyvi13mMGPt/L
XtB8iNVbrDL+ECwAXsQ7LT6OsnjXjdB7y/TREJdFSA2J/fQAnpgHfuES19bu1ogx
VmVzHRZo+gtiu9McowzEcGK8J8DwoB13ARzhGXKtwL67tAz+7aNsmM3qW8SbMBez
eA29okicZhPDT0sjDRlTw+55qWhJsBmhgL6YVhXRozXqUs4MQHE2sGqru338FYcT
d+fGsopaotyzmrPKNwzHNizSWa2RfiYNghnSsne43T8IX18XjxKdn7D2P4hHLqzQ
KNyRd05SMolb2/DISjXrIRIucwVr8WKpaI/Wj1csjIv2cpJCUNTIaaQn+3tdn5ht
qMAv/oSgRzXQviuGaOzU9DLGZ3Bd2LIGfVv+hKaLGjAmB3/1aDizGhmbe1VIC1XB
GTXXST7dsU7qIehwod2xH4pdo/ii0Rctt/wpoCkDqTYQHdxLCb1lKgPoe5SGLV5W
Q4gpZ/nAZsKS5faBgHZmMm0xnHHeAa1jwrb5f0EXxtecZQfibmTuEI8h6238Pwm1
vN56A7oaycT1H/tRBw0UrgeQalq/7YmICZhrz2MufLba7GXUtsTq9VU2lWhGCyAx
yhJGmH0GKbaKBIo8pexHa/GVGFVxPcIFl4mXvT3k4YFWtGIhcRD0fovojKlfojwk
RvLrrpIRH495LQEuFvZpVL+7mZyteXf94rFLgMawr2d0J7BwQtgzHzWnShbid2bw
f9e4pYqT8w+2/GRM+IdqKJFsq1Z4kZXXdiW92bnj/EeVrv/27RRbOZWtSnBKQ8G6
kgcZiYjmuGqZ36q9hgIOlONsx5VzIdqX4OnQwxYJmJvCqkrUtotrIswH9Jl6gKPT
Sr5PRszjcmj08MPvKdeeoUCtIPxPpRQRNtDKtwVmxwNFMLwusMOkmzzwOsuQHdLh
8keHtL9k2ftM6iR03A1vl03ujH5tRGxAA0u9fYkJIhQBaz0LmlGUNZbBBYhgp3cY
3Jdzy6g9N2ffWmcmAHdi2a5ydxjrTvnIksqlt64tcaJI1rRblpS1gQb1ugSG7wkT
JAcuMyeVGogRLaSwJQJXCu7o6gfwmZUkXkzMEvTj3CDlag2BsnXOuIpeFRNTMAt9
PoL7bPTs3whUH/HbEoCt2mbkCpLHN7MO21/qPp3UTA+yazDLdVck0TNSy71NaXOU
i4LlCZbOoMUJfO+o7XoHAxYgcSUmB1N2h8pyyQYycS5/59a/sapUtk9YhIXUw9gM
IlfWk0a4h0+aPTAIpiei7nFzbHtXJFfH6NFyrJA93dYoqHJyCgyeH4jGwV/iF79E
O8fnwdGyejUE55RnCUNIDVFo/z1fDNS2NY7riMymfaFuhWF71gX7YnSUfrUgWxx5
MCKyX74Ssk5iIDmrYPe5bDQii8XECbH0ViLdtCnSFuV6nJo0WdMdGyOrepn2qx/0
ghhng6WWY/pf2CGgYhVednNqAXuWxB0+4uXhG7s2b4I+IzwmxZy03I5zD3tdZ6aN
Mc4o02xyvVxF4lI/XsSUOM+u7NYbubhuIVB0wUnhN8WddRz7VmClxa68v35aOFnb
sf1HmjONZs0O589wDbUByidWYBSm+vBogMxtEbCFTr82G8+/SI85R6j7wfN6GlQj
r4Ta64Gec7kNiH7J8zxbbSNMe/zFVhOYoUve0Wf9wGAZnVxkzY5b+dq1ftuPVrVP
ABE1HAPl4VMd5dQ8QxdSYzJDb2GavY1fvuZIF9AdK98st+/E8CoUiL2EUZXkneST
8ul1Kfs5ttrB7boRw4ICC1ssAKfEJ9FCkGTVk5lxJTIW51M19diAx4k7tHrgcmUi
g0NvAWZhGwbfyNE8X94IboT7joY2Ui24YsP33rbSAoi2jexXlbe5bLyxLw+k8pue
Bcg3Y7+uLk89CsUWL7an39c+v+JTr6pwucSKea3d80y8SNYyvcOX+J7MdYp9yJXv
aYVQ4pyv8fUCefueoD0PQJPGFb8XuaHywJQQ/HKtoedQYB23kLomaAWceJq/0QS9
1CemigUK22yfqluuWwclOMKs+wQhJigf/XJNj8PXK0NIHR994Y7c70xp/Lh+/NTr
YkDUSQYNkQ77uDh++KS2sw69XksmsenlrAjqW8O8dcvN2uWqwg3YIQfqkuSVmISH
hsPsxtsDcxU9KzWo+eSc1rixs/FIZMQAkke81JNH4tg/rt5vQ9KUOn5O74YV8OJT
Aa9V7bkDwKlasydBDP15FCLCEC7yifSAKJZL5pUldtCLl8hLl6rmeeOAYSa1ioA3
NLpkXluzk+RfxOIEV/i9DfzOfJE0bbXIjVZbaWgjqJisqrp2TKxxb8JSiQ/3TMQb
JYGYla17Xkjqx6a4hB3adF238Z1V1wnNpRlzAMgDbBgaQLRHD4onWKOQZLhvp4sn
4M/dWQNmBGjKkkQ2Xpx2Bm0BfxJ9jfXKEFkNx2y99P24agNsdLW0KV6AMtqB76YH
kYneUWRw0rhRVofPGuSbjXJJwYebd2YW6pmo9Mmtgfu2pVhJy+nunkEqvpH1ht/W
f8meE8pC/vDspCRHRPC9wvWyqYpgA6ocM2COoge90awVu99YvMt+O4xBaE7+eQ0Q
M+/fD487jbQMoR5bujvU4K1mNnz+aAPeK4xVNiF6g0Ywb6ZDW8iOMshpFsh/EHw4
USKL+hqwcur00ai3co7R5N17pVcbNX0XgOJ8tyk1L+oyOnvQl0ygbHaC6+lbR7Pv
P6MmcdaiM/VdEDBI692vmJWeIf6N9JCxL0CRYt8oCCFYwDbsyTybA+lPezTwhB3U
jmFFg+De87elUBXwrQz1RY0RmIbVgIeZScBOZZ6iB/juGq4g/b5MBogN8Itcf48C
/UwoPp+bg91gs+TbTVsGKp6L/fXGq8Lw1MeM4XK06jwFxcDZqJwAmQ1d5nHdRqRP
Sc+GsahTvwtMmnAopP4Obd4vqCanK6do6yEvY4BoszSI5pWld5kUz3M75dRLUjwZ
cOzpqYrQS4HV4QhfgCFtDZVbN5BwUjWfj/SpowehB/+4aLnQpeLROZpicrYx+CcC
sIo/JlAAvUwUb/TY9Gp9ldvPyQGZxc9WMmJsAqdHfpy6PyqSZCGM0d8iB1yBS+ob
rYIORL6xmiiyyPJ+SANgmCILrn3SAsZ0JTM2gKpSHOWnrJGYURIsVgu/995KK7qC
soZvBDtde/nZgdD7SMw35A7b0UOg3bmGhM3I/nyBeVDRh9P8kpjC91qyTwVDmpkS
LXcHfwCspQZxq7/lFqyYvtnt8VbtPuyVsUWyowg9fjQTdGOaJraZx6637TlRBV5t
v+ollvNzZgscAtFriQ0erpfc49RkTgQi3pLCrhzQKhGj0tTZnluvufPt1Ey1ngeO
la6xDuPqU8Sn4swB2c0L2Uw3jKlxsALCTWnjRaB/KOLhYkIu1AOk5LiG4kdkRZVA
oRbkmtoyHVB8Rf/UOd7ZIa4QA3uK0e/dEK2c+Xy5s9a/5bZBGUJHdtP6yAm7S1L5
PzCDchdTt5V2QaVs16Dfxbg88tPSGrRlAIqHCcX6ksHaO6lflp1XAqicSIrMkNib
N2Vm5daAk15ZBTvZQwdZ3LMYAsep0+MT9km8vVof/5lETpI83QRQfLcDekoJbdfq
h4ZlqqDIYNLLcf3C9Y0oOz2I0oRlK1Uc8x0Cv66JjzCTiKiOJSNy96Zm+xeLIU5c
uuDiLJM0x75OfLrivrIbkLoRA9FupElA8eywnMangJSefKDQZVJNbgSgxvUGHBwS
rfk7CKBeQH5XYYymYrxGXw4nJ8tiMo0KPlj+VGiQ35hXzurQA/KZkxs3E5hQoU+O
7WOI70PJzBWOwFitXY9SBpxkLbOeX8yHOeoqWJBc2NR9Iwcslp8IskvpsTWXsbKf
8V57wdBzJX2UgJNffKBKY7VvhT/Dzw7NPoCuozslZQ9T7UkrSAfZgAO8FB94XsxA
R9Nncirz6IUnVQl/q6iMRYKYTMQzW+By9oxzcqPVDLSgrmpsMT4FIZMj6T8GSWFk
YptMo5AOQbWCXSOozNQsRQiypwkKAzVxACrQAlyadN5FkdulSFiK2mN6alKtlUgt
i6Ym2WKtDAbjreKEKZp3yoHH1ClMnWt///gZchFEFxvEhT9LM+P7L08ZnTdi2OnW
NlKB5XancP61SBy05lwVpX9ncGmwBCZL3Sg1gzjypkXzUYiNeJ41kXty6vqIehMR
Ule19ghzIBpPGh52pDJErYd2JqHnqyqFDKTdlbzeP70+WeAkjlOa3SiyUJgWo1y2
1O3WV7AmVHTiKDgKvJpn+JQJXYjMEdBa09S7chOdF2v2pt97rO4BHmYTjasHNJZV
GHNuDAdh9rmB8g1fxuJuYfM0KhybEMomAXQ0M4ydScD7A7nf4vIgrjVjhp2tu7Wv
kmWoeRJqSYNivSJnwcn7aGWIocwgrLKzf6QRcY0yg/R7JpUINqmLZ1sXgMyA0wiz
9yqbrOz6To4kjGJcWfe80iUOQFtsIc2UHSHuP01ZVIp4w92v9JOHDVLIve3+EQNK
eAO9A/Nl1Uo5CwIlld16div3ChNz+TJAEpmzQn9WzPmuWLjgSgR1zhS2wLwqQmYK
59ihJNazWUQUu4QSt23bKtWWtTYqxIqHZzTAoligHqQyyHoeg8PT+rWfeAkcMEPd
3/9PcVuDY9Qn9AQ8pU9XzBuJ8WmrSBegDJpvPYQY/Ac5756xO21U4qJPGggsOWYU
XDq9xJoAoOBWuZj/qaDZErrcqtOvRdSDATTNfqxp6k+rjjYc+8L90Dtsz/exvmsg
ktJEBz0/B50Q0VNHA7kKY0dp3pgwt9lbQE3KsaZ46Skl07++vN4Zjdr8oVLev6zh
9e7LZMvpBSmat3Ji8v23MBLMFoqaEYS244AOOJo6QOFUjDozqFWXrTJYp8h/CgNm
WSncFlx0XmnJbHcTonjLHzsSjKWovp3+46szfmqTpA/XanbKPoRWThWhBOmazSUH
Mo7zjW5ngwvQXLog9pn3T/cg8xJuXTGIUMOo55mDSRXwr6L9Zud/k7CZe8WdeVu1
h0nARTauC7zkPmImkx1cROdqQFU6FIu6y8bE00nNEPKT73KfnX6mg9UCSRm8eANI
+i7yYmsBdyOS+9XR0pwUlPL67xjzQ+N0bfYH7woGdY9YduQJ2qqMxmggN9nkKuRr
NUlgZ4+ITFrDvxeTvqTMO/rwgDY6D4UG3N4j46Dedtl+KonEYxRm2Pm7wx0SUnpG
nbGtVmnWRgur5H1mlCV9i+qzZ9e3FpAd6BmDVVibp+ks7CP+g4D9voR3azCtae4T
LU/U0XfONI7licMOESccWUes1SKajxGwkjBGceAqxWXA8QgWK2dnf4ii/ENsbn2e
51mHiTbN7oXv+83va1vLg/MM8D0zkIie75tEVu/JGVKcApXDvyKZxpTSLMZC9wuX
WeBGAIBV+b+CjrJTHDAoTFjDSAsJOuCfJohfusQi9bbVGBwJDlRpf9C+AxFLJlJk
HqWl2Ye6enoNQ/X5RaFuHvlPtPxlHQcqfJ9rXLeAWIJGCU1a77iV5BIgVwQAza0m
teLDJ6cEQ8cnTw/b7gmN0wl60QWhQUmAxYUqDr7ltj0sO/NdBkib3+ICMOO7QTY3
v9lCmyXuMGrncbvEf3aD6sJjnLQXgCc+epLqfGqT2Y12zMEieXFfjd2FudX7lkAc
j6LPwI53OAG4i266AYd5FfVFy8FQhj9QSIDlaiLdPXA0mcBUItwRETur+ruAcR1w
6Gr4HOb+MY9O6gHh+WZLqHXZwbSwg4l3QIskmO+hYBEXoQda3spZ9h6rrsbYBMyj
S/8u9SuvMMV7pI1mAI6YHc5hbheGIWcAcfbU8RduzBXoJJtgzKls3xcbSftosob/
HrdTt0f2jGYjaKjOkToK82A/nxOvRQuMAC9zQ/iNmXOSq6IkxifJpwBJqNZIbH5Z
40DnYGYjKt3fffR0/YKZtW67n+tYfaWwai+Cm5HKudsgITHQ/pdB1UYMqHoORmFz
xNYTXEkd1nhzwg4Cl1m2/xa0WaFdttdtqQmzsbTc6fclDZd3ujCIKbBo0dHFl9lY
xpJry6kGRWaf5GUoWIYQHbtSuF7dOhMqgL0jaeV3RGCJg4EwcLPYATqwKeM7RoHW
ha10/4hgFx81c7npvdGCPSP0EU2f27/mJ0CXKDLi5/4VseVddpnGG8kYJlEfDm1s
C+DbIklwxvM7K12sGBOKhX6mtyhRBvJtYoZJA+tScbvZI9aq39Vt6w87VsR2D6Wo
owNbY8gmySVHgxm5bNtGNCq8f0DCk/cgDRiTFQcsvb+mhUVTBnfj+ml/miKH4Um0
zQ62BOa8WYJsfPEuH4tzHXopG/4bKm3Ga4lV9Drw4WYPmRk3OcTmT7263djZHVrQ
7uakvuT4YNlKOrimXsQmQ4ZUPw/ZrwBTpyU0bAE/PrOqpEHO5+s30YqYsXB9/yb/
ifGFQM0shy0sqtCuppKud6LPp2aY98rsgH4EAkFDN5WuRdmvP4PvSIny0HVxLjRa
+EY21orvYNcCiGbxeBrTUPrKqeDITGd2JRBILEPHdrKKZK1TdAjuNsdsdtBbD24X
xYGWuBSpRQW9mGYq3Z3M2I7CHyLMWsOaSYqcIcG6Uuap6aKqpZ82kNqm01nMwIiN
34MJ1hyc3W7g3fkiKTfllWpwicKbRl5Flz2cgoGRwzf9bJkJOlcBJUSDh1KCPITw
GJHz+8GK/0L/oZjqi2R/XnSjf7ydWPj5FKEfmSmb94H9QrOZzTWpC/Pt4t9Idk1l
T3qiuLUQuh9KUP5Z0oUKwH8G463NVnJOkPm4S7WIBrtgBBuq9YIT766iP7MYLzYm
IO7fOhUsTHh9UegBNrI5dXMJ+zYMMNumWtecLRrAVFkwLds6La8lXCCFloJwv4d8
E+wU4SZNPmTIezaYtra092FFp3xsHeQ8FksD6bHFCsi8pLWhs+UO129WZIf8sNpa
Ut7vpQMQhR54OASwJorecZkKG1sL15R8oN/4D1vSCXawGxVXb0okeXrElPtpjFz6
60nFX4cIUqKQZg7weUuSjnWdGwQyDQLtKzqrXUaYyWKf5iMTX6V2P3+k+HdVsk0h
jDkphz9VFoVHixi3mnfdeHYU+faR1l74mfwchDMeixDlWW37nMGTAUBCKITG74cc
GkU6litSyVMu67ppU5DI5s9+6+VsgTCVBm74/Q+lzTUi5PFlENAwg6Z809f4Y7Gi
BxQ3Rdptr0X5wE5VdrOSoEpqKhH4bDZobxRY1FdwCQFhSahnN/D/78QEghb86NgD
dq/IpxxeTVYDs9RRVCF6bZ8ovZOjdsNVJdEuh+tlEyxZzmSvfZDYSX1CmY0pCBMy
dp51BsFwfAhPVuwonHtjnQjn2WnutJ6iwosCpECqgVNFEpeykpcsHv+ybLBBZDtg
IOVWVwoNTH+NJKw1Zy/1izwfHNJjrb5T6V0eaS/36XY0Ts/Sb79+/vSmRnAHm+y5
XcjHQrZZZi64B+1PXwvnCUj/Rh/o02Bga7NUMG2cEjd0c+DKUMDHWQkio2Qb1tS0
Dbzz9QSxsrqtnvMDEc1w1mKB7rMpKBw7Ur1SXMCQ7qSFxbVNOkq31oc+rwWGMNR7
VsHyXL0sNvyPzO+OWXQ2nlWfLHYwUqqQvNY0abhLLGq29DpUcOYG6E+0A8w9sn99
/PNVcyzBmSD9UdBBt3VE4RsS/yHQcdzLzMGSTTrtXZM9rosUs7PiuIBapfmMcULn
7cttygO8LnpZUfdESGQWfrhZPPxnrXUdaLvM3kNC8whAXfthfnPwiIzGBXc2kmyI
a/fTQpK7pZDbNO4Xba1771XYHi/J69XpG1H1XtBn2+m5ufGt6NPNfUOI4MdzXEGa
PRxVGbDoby9UdN+gusQ3yBij+FdmbQpdiK2BHmxfc1bE2QCuX+++8C7ziXAx2wUv
BHEd+NZ2L/54K6eFMgK874Jhmb78gL85mmlL5g/hMxtDxaUSPZeeQNfYbAturMe/
BIksyTc9sglcY/6taav7DVP3FeHwuvFGS8FsfOYYD4p80fPDWjGPWLAUiXRzrv5R
qU/nfWWhJFtaZDJSyFQa1VZSgoFhTSLDM7AFRky5Bny8cQQycfn5+/Uy3aWx1dSm
MtY5s6rUFvFy4n51REk54vYi5o/FMZ90DL3IbA49Dn3a2HdvWJTcBvPK8hQUSRFC
mcS0Z+N2sH00WFwtqytRwPR3yiM4wk9CBQmk6NqlOmAg/T2zEoXQEawpMcukWnj5
eFgP6D9fkzvnQEAExs+46hVll3CzZPoa8SZjsnoTrbBWNBCzGeVavh2qmdhGAogY
RucPQCgSs/lEWthVcIaSxWa1y0jgBVxxJQB/hWV7d4s8S62gAHmDv3XVe78fPy6C
mdRaux0vl+QhX3VMORplNWLgAy0u2vscJdwYAF1rgDghvh9zvvU0UcPqdkR57h7Y
Kmd2S4CSmgY6waJ0ZB7DGMGj3av/UeERZJPJC2csU55TZr+1pwSjZxJ8c3//EwYP
bn72fLAhSgZhAX/XnPVfBNz0nTz7XgigPtaAgzAkXsioSDqQV3MohJpDrJEwtRrB
gGeUbVGjUdes6xgqnU88HbwmCEK7ZC34B/e8+rPtxSUismVep0vTzKabHJf8yQFh
Ha4xzMJsaQwzGVW24e32x2tlL40r2s+ZBCK5bL3Kr8y7sVYtqqOvQgfoOWwg37dK
7xxYKarWQ0YksUZLH7lsUrlsvUBTczcmzhMo2eQkJ1MkqgYz+XBEnJehikv7hbCe
1eW2QvWW9rXPhPrPQQTQN4FaH4/AI1y/wFv3UNLncJYYxKDU2wblM4yN6VvRiH81
1t9Pun0EYwpLyxGJNKK5iV/90rbtB/C0KnrM6xb51YBA2tdjRZBOuYjJi3p7J7CQ
cOaJvc140m08Lu/MN+nKlNwzuN2/iSUHXAFVecd0VCV2pAS22JRCBU5r+Is1TUgK
7zd7ByBY1cZlXUJX3SZPwG7gYSQh863sS6n7usTHzid9Nsd5GTnOxROj53B/KDAs
4K4Bt+9XEHsUy1rlIudA51v6miqEb5of8iUdwR4S5VZodkSfxT1uDJamCxxRiYZ2
wVYI45rRslP9A5m7Th1FVikzkhVWTi5Rijsff+xL/XvvEZGVr0T2Cx7Y+i7R9faP
aj7i5kc3wsdjSAEDY42pQtUPI9nPie9bBYOmho4mlr2yPB+E59JO+FBprGHBCJEz
WhazSmxG48+70hG7UaGk8bxxACJAc3bqehckOi+wGTkYZRo5tT3TmttIIRcLuMIj
9hTrQlG4nejDLCXFWHL+3bboOJVutDaO04+MHYpilxp+0FrSwbatirNVBE9ob5Gt
fmLWvAtfcBQd6bXgQoKnV/c04Q7uiwnlgoDFXbdYeprBl2LONRLinDjLIgU7yTdB
G1C0oz0wOI6owB97+Z7djobddzVBZbD7dXxYEjCAZLMDYOmbkjWbfjdJkuujkl0u
QHSD2epa8rdjraGjYDdkazjWtsj6Z/EzM8WAddAOPjvksVGOO2u6GH+jFkYd72my
WgN0KYN/0Yzo8JPThB31woC9eIklHUvtFIazaw5TETxrUsZPSictZS2c9/vayL42
dVahofru2XnFo8wSPxXKKs+WtxidoPB5XpnY0VST3r52MELw3EgBvux9vLcBN5GC
RzfoO9YQsRhideUQTDOsdvSzq0xh4m5zBTGJ+qFzIxVqN5IIQOm+E124bjriZISC
+g8QvsltvI+yUWyKriO+/6InrmxBrkkh/YssUJUQXGmCbFw9c4yYxGLCNd8luhAV
AvBkSeGNugGadKHowSZrE+KhkSKlGSxu6+1/SXMT+Fof0QAnSl8O9t1VUfXZ5sgx
4KSNF+hcgVy6KGFGwrhiJvfKtELiRVZqL1H2pu/a1tFyIY9qjhKVV+Siwo20HG9S
1Oqr7xu9sgnjZHqbuEbpw6yZibwcoVM1Fx/SWkFJxAf+vOEjJfvO8bCPRByja0At
flSqD+0YIrbV4Yke12BbGSOD84mVrPSiWf7+hZgqlPQiebjxtuCp7kmOx2eyr/W/
IgIx+adXmOzcFkN1KssxrsLy8ZEAltOFn5bcRY16HtXAFP219foCkc93ZapIWjdG
jY9mNNgvAGMSJf1PpuqYfeCE/s3zaq9ajq5wozGstbZj9xenc//XAvinYm1hSWa7
V+A7uoJH341TKVocjqhzWxBO8Td9Fc+PGuf/NWCZKfiDdWfmlXD6S+RNjyz432Vv
f4dopeTxoWbrVf+A3ir7OMH5i/0g13cmy239bzBNXyTdJIxqaAMysWfZFOpNmO7R
NxCsk0ckXNwnDCLG0vInd8CxE3GlUDZC2ZDrgTgsCBZ4438GAyGndaQLbV8KdWLA
9j2+UfpyrW+9/NKmxeeKmsvEHy4HfC7HOUgQ+4tt+0iQFQMVfQl3LsRR2n7E/cZd
5B+fSle1UJuOkQUVGl9nmM/CPJpdDEELObHcsrAxBCFsASijqh2XgUx9I1RTwJFX
y62dPa4C2HoKb8ETSfUvhXDYSuhkwJFHzRQ9YkODcHTf70uE8ohFM8pOdniis+1C
BGaNmdkmUCDZebB19kSZNhdqu5C2HybyNRO0MfkJCJB4oqelsx/f0C2PV/4Dqqol
um1nHdSRqzDGwoJ9j5xVbjjsGCEzDm8lWminpjIZndPi/TqhOgL/UhNnNBhWIRvP
++xgzQabpZfBeJyq9xRRX4h7OuEdLfJUP5tRU6UZ49Ufcwde1z/LGReCLJ4SKOcd
AoHBeLWfjy5tLHAaer3xCepp1whccWnUovhAUKU4TuaL4eRscnRPys+Q7l7zSJWH
96W+ZFHpKplEEyrv/3BOgDDIl0EQTX618SkGAgvUfEupJI/nVpUz09FilZ/Q+E9l
jVZye+V+GgN2jvgUrMB2oTZH2cjdXW+71TEjriXg9xvjrmjnGRcWNZDYlGZAlGPS
zsbZmkypLI0Lc5B29GJheg5H57lLfylHYTTHF9U9QL+LltyrOsiyd/fn49yRwv8R
S1uToYY27koZtXGyXcszNDPuSjyxCQxOQ9bc32X/ZNrDqnTjWTHyMr6LcywApkJ7
5cEVfqosJXrwBnDGS3xpc4TBpHUWnE+TgNAYHzL3bYLTMgr+sl4DSKWnCOLhPJM6
jgumkxZ5r6njrOjL0SiAwny67LP8eNcnzdRbVsxoyPkqQxiUIIxZayOqJsOW7s8B
nDEi/6n6H7Xj3WsxawcCG1dVuRgiO+ktQU43SL8/lBDSnapNTx0fZ4w3otRDdqyX
jmMXlC+k9xVv+r4Hzn+x7++Ptsb0WdkK94lwg4KnLKSOOpU+ULhd1IosQikCNFu/
Atv/liXae9kmdJMm+xzq1gCL5WZD0Dn3WeFlaFgQtAh+NFSDuTXQu4mhF8uA03l+
jqjmnkIb+YBDDYkJEXKipuHpvT9ZiE7jfPTXIti+oSlKWRtGtrLowFwXnufsyVVj
twQMSK4OSuBjpUGzlPy5yqXyDbBxa/4TsOeQtn4BxltNIXAYm4gkIAWd/lqBZraU
4/Xtg7lD/V0eVw3yYmrb/BLjRrcnl00en3ILtO+ydBpFVIIh3mxD07bp+Yn0AJ4U
5Q20E7rrDOuEVMvMmwwWlfAG6ShWwaEylR1fcZ50lsjLkZ3r9U8k1kO2ZtmoTqrg
kTTOVn5Kvv5UGHRm6hBECr67mIUljrrXfb1I9fFRNSxJzfYiai8f+u6ibJIzPoEo
CTztY0A+y9MSOtWDf+HepEsKVKwlWJgOMujMQcOO3r778PA0Rj1MRBOMuFlkOyAg
oeVampvW9gl4ltcvKFegFgqwG48ApTLmfnaC3uMj53LA4tYSpXgHWnf1kI/mzM59
XIhMhr6s37NpMe4CDWchWZvFFuZpVEYs3sWd8o6HoEJuXSh3FeA8GLaf/og4jpBt
1m4kJauks7lvvduNbao/Lflx9Ym2s1LifHERCXC7t2sBQpcTYJ2OsyBU9l5yCP4r
/I4rxwOZJMBlEG7YqeyuauDnV4Wm60aH/xr4lqnPy3Eemzz4pfJmzAyOOIOf/OfU
9f0rpgrju8aJFNQEq49CokNAVUgFQLzAxz9UCy24QmNjlVjQtoGqWX+EkSSokVta
m5ejniMd7F8u/EgEYzgKslE4ScXkxBH46DleJ3rY1+qP++7w7BFeRSJkM86JLwjW
TxGVhWgE5ZBjzzWHadFeEG5xVZO/X9LK1HuUZwyxqhu927pYgDO6LE8PQINCa49Y
SLL1JenwNTCo8cDYKwHnquegxkrqO1NM3edyXYe/0UuQjyloYj7W+AS56t/CSN9u
2lXnPeadhUq4/stxk1ktcVhAB5QthmXer/F0Xy+KCQU7NZ7qjrkBUEvcQTFRQAH6
snQpCH6pKeybhchwLQSrxxKs1+o37Hif1EfW6lFkrVBV1dJVBApuZJd8vATeTikN
dAzUOYOWvOZdR92U+kWK1Xy5DpaWqr49O7qJGIoVbywcwido0nWO1FeF4LswAbuS
gxGGXWeOcTKtSEhGOedivmpyFUe89pMiolbqrogyMzbCqM1Loni+nKx17VbKRWY6
yhCvKVxZruUk5XncrZW/wVFx/EQAvks8MCii5HNZKYFWub64qgn7izFC6+N43CIU
aATBaLDBTXI9DzB/dLeBH1Pheu/5Jwi2OnjO0cyVwITVnsLGyin2sCTFittj2oF0
3bAY4JqJC1lDhJzRoU3eOc+34iXHGdDlBneuUSfh0/FRqg5XnaNM2ZioxFa+IoBM
xKjW0eNIbJSxWVJDQmn/n04xP6FqE8wlYsIaivqbVxKlRotadwjpjr9JtYQH7jhi
LEc4IGMyB9+5UF7YubCtC9SS84LvyU4og5oAp9qY2OwpPd2EknOcKKmPGGrb57Nh
r4dMJUsKgLBVc5QoT8Epw/r8gfubAfXGzo+aaG6i4lIvsAGvWv0PdWJN9ZQ//1Gl
+cfvmuE1RCJGSjnRHgAJcxcHH7xFc6ZJxw32CdbfPzJjK0/FOTE4J3AtNGD8OXqN
f2vHobMYJYg8IMbPUyLpNGH+6x2o/sGzkfa/+NYcYhvSpVpADqZbvAGjY4ZOM8sI
P12ZLwr9HB1BhVMJ97m6FpUyW0ut82bxccNjNpoJ8nwZoqdCncPnyeGXs8xbhKRk
xYXDh759FQoLvC53U0FYAlki+wJXX8/Tf91k5U4CaY9DsgsbLbk7Kysoij3oM/AA
590g9/LnDMcWfC/cHMymMk2HZtKEliENUB7f0unW6WcIb4wp2iqoFgDhoIuGKnrn
/xiRF9hF6Hj8Rd2wC6+QkhIODQ05o4IRb1g34Gs+u5DUY/6/PM/hOsYNC1CL8rPI
9NjbUIk0UsvGtfaFz3QQ9KZtqbg0QAhA3OnvTDJkY7Fs8xewSjXtOzVhzAC/diE/
E9FsFblFhvoRGXldQexGck5SwAB9246duTDmsldKfs34+S3BujZHeDWLXqFyIrCK
oM2Hn83j1IeQW9sIWKOsLsy8lLoMpCE9hYLnBuBmtPVy2gSUPmmUrUe1tomqG0pR
JtfUdOsSgz0zaFqzBXlXfNfGtMGWT5OTOcbXdo7iMrgt4WLeKVzVtvyd+j90lWYT
WjmzXC0LVKadYFam7+FcIES6+D0DWTsDf+b/tEaPGFY0WhNVl5cv81qib0byXepq
pU6JXKsK+clkX4JdwFLk+bJmHJBcvdH6Nis5h4nU7bAJxPOk58PCTexfilLfi7zl
den3EnAEeg6xe4k9sRP3fRdgNGCrIfpKxOqYMknDwubedVQui0Iz6uanffKip7Rv
8zkawj/BEP6i6opLja6bCVj6iDwIFsT/XKEmBMZFmmqIx98zej+5+WSKfKe7vc4g
l66CyQ72d5MRaaMNRbZyt69f6buY49a2b5LWtUgt0yP38u5+cFoH58cGhQyclAmc
jAKbrbsyJo41QZ/ONh13/3ob6F4RqrtwwSIRhu3DPEFcAe3kxtK2Cni/GOBch8M0
mZZGzUgoEDcpBuQm1VjIvVULQ4Cy53VUnMBn/XPL8Hc+hh+jhHSouDulekaPdLKA
K0FMY71SQXwqNqz+6ucU1WZQdCzXdCHyrQTBw8n+K/dscVWpm/RmjqJ1Cpt/VAMl
sBKXaVcISkJvVzNw5iGVygS9bh6YtzmRqtVBXOXxh8m+U3bvQoa/h7qaZf2k8eqz
Xc9EbOUMwXuQWKgTXHm2ajC0QpHbOBOPiE54PXaMaVA9itKRXrCul7qFjVLZOKr0
Y8DEaXiCbM8aBErpwu8qm2o9BFHsJh1n9oQz8JlE/4bOy+Mi3CXhuyCLs9PyJZA3
WyuE80zyDiKKW1sCXAYV5xc318VMlRtzSPCEdQnhgfoy2bE8wNc82B435NmGjVRJ
nh6ja9eK1qj/TONZlDyG7tvNINkXGUJaJJH56tHhjDSVzjBdE2dY2KN5YIlS0IGH
69UDEbzY2haNGuXJLny/L2DxsZVBemZQ6AtYJHae3h2QqPsBFPRESnPRs+HVfSmj
Od6PMqorvF/oNWKzud68QmqM/vDo0o2wE/mc2oacudX0hJ3FqUa2owU6n9jUus5b
PlQpykuYUbNiazPnq1qAPcKRz4goERkHH0Kpv9hp5L6LlhzuSOlwN/ggXIZ0/AB0
PP8fPUJZnd7zSlDwQ456rLumt1xQVjKhC36Qt8zbJ2JA5QpAfFfrftprjkSNb5Cw
9hmzQoQIr1iH4S7olyYWa3AU3sm8p9weX4gYSF9LPDykSwru+A5y3/LouYjrwKNQ
4uco9oS9GZQkecKEEdfsRuPKMpxbzEomcugGPFtkGcAvpQldifkpMVNVQUjOiEQr
Xi0S0Aiur4ugWEZKnYO056G6+VCCG28D02A1QfGGHzEXBeIiKEoqQvxW+lEh3QuP
AwnPU565iN2q+KGlql/JoC4UjuOWtTuVg0+HqH/8/rm1l9IK8y3UBRtPPvZaCh6H
yrPzegGsACxU0hsrgKQW2vWG//2INY6ZMdV1qnznbcLX/KIFhnSMlnCrdTQ2r0En
L9ws54VIe9KBNph/l5U7Aw==
`protect end_protected