`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3328 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRo5n418HUi4GlaQEf4lAMgCmjPt0lNDT0WunfZoEyAYU
XQtGE2oF/Bv0uxmgfghm2Ob+VPSxb2zXQ4fbkgxZ9OqbjvL5I9wwF+iwicQdnwF2
IqwBV22n8nH0uQCuc7OEFduTzLDUHovlLf/oym+6BCiaBnyoClF8s03Wd6FWiQ7c
kVZvMsKH6SfgQpveTsUNpBUMz8H4oa+x5J7b/4/83mcPluPDetqKd5Dri6Pu1mbh
4zxwr1vJdunJN8FmsgZ/vXuIf14S3aURyyAVS1ekIbOSlS+pvEw29Gq7QlHuN3pU
XkR/Yu+CqbOeFCrnjOxr+f3b/6BYY/LlGFwjf1BYzQPRBGjzWOesGjR2iEa0nUV9
W1ZurIDqw/ofbfhGy4IVRBUmTztu95yu12EsDOPGYUN3JoRNFAyo1HemqY8AjNYT
6Mc2A/gE1fr+xtwVa6RIcHjA8r4C7LvDMYGKxqafYWmDi+hfoj0lj/QlQsLK8q68
cEdiiQZQADCJVxVovYOA3MrML8GsdDoOhG/sxBT0XfeXKAUeVB5+NxeN+D9LARpe
VsB8rzBqGKUDtixrBHvynwE4Z0SAPLekaZK561wp72PfWZpjd4qwZJgesZHBgWdr
fwwY/PTO0kPk8yIO3TflZw1Z6ilgR0oPyuOrBoGtS5UguzarFuM1stziQRSKBPqL
RSQuLb2WC2k5UfS+2Mre+zcjSCR3+YPUn4eiH9DPOpj7XrDLxrNiQE5yJ2VauYg5
/VANKVQWt2yEQVBYTGCm7aBHUWb8bysEaDzkaXBAfeJYgcr7XX0H3QCOK+TqP3zk
nQZRsK02Tt8iqGx0kNDmr4MM4RiXQyPntyGqWwNnsXTtodbKDwhAMEItJhEJ+PPf
4EGID6EAz0fBLCneCDJyEeOFBDVwXQ6OwYVSB1cj7kMXQR2dGurt4Z9kERxZPo9w
Uea3dAx1x5CdomFODorLuyAbt+SxN9DXtf/PY1T2NGqM5lNcHJJm7DfkSqIILSqt
t4TqjZjQTr9hU0wbe/1WNhFDGAzFQY770UeCWU6W2VWLYIw+B/dswjqlsQ2X8NdL
5vGc2GROwLd1ZUsZAaDpEP9LMFsKI/xRz+Bk8aTRPYCFpQyz29n8YX9xHOF0DSAP
SXhj+7U45hZJWk4MEckfBw4KjpiwahNaP4DbrXj2tjyEGt9sJNlNWB3wvPBivvq0
XAF3WO6O5FcOghti9Q9gQ29vY7LFoiEIDVd/BzpboybpncpE/WTJMlZpUkN/0zx5
Fug7s1RIRGY5unPsnOP1wMDoXsI5Xcu8kWcACD2hzwrxmnx5OKHaizMOwYP9DoOU
yqH6FDMSy6YDWwJk+Tmg64sHYuErP9yuQh48XkOtG1wddAKR5LHh2d/OlEzN/W5s
UbOG8CnV75QzzHoETT2fhQZvu24RyZW6Botoi2jtjSIGpTJZGxAYZ006bA9ry/6m
pJ+f91rEzfibzP08x2joL54P/r8jTK6IprKmW1FzggmAN5i08cxop5ePcX4rI2j4
Y4miseyVswuX12WINEh+xIFtOODCYAdiA6aAQxn8MEDnIVyVS6SPm0apZrqiSv8H
qbfLWPkjjfW0buFOgna0HlVveW8iStNDmN6GTsJkIwppb3fD3wp9ZM9DNv/xqAXu
FHniGa6X8+jEZS6esamJqIDpM4gzDTis6PFOjWTKsOBvzAC8H5N7AMxvVuo9n79F
MceGQZNMYXNeOfpT7CW8NCxMgho4/JExw0o7HU42ew2HFxRQCwNeY6oSwfEqX8FM
PxAG5VzTfHiLtvN1OZK28Y8gIuCOYUJOu8hPgcPu6lqjdocCk5xyJEN69Xg1ABNT
Nkd87lx86CmoCaYQmMLT84nGHzVCmv9QVprbDrwwqSMQbMb4QHiMWqb2oJCX7ylU
wDhLAmxh6Mo6lzBDXwfA3RWPhafRXCA3AHr0s4TLKMYxY84f8p5DQxSb7VAkGhP1
2DROljKCQAP3j22apNU+62CBY5ZmCiVtirhpO3H/OsMJ2QgcjwyThYgC9oMwzeUV
mUJ0cbm/QDuF75OYnKDTU9MXFdXOB/2QDWV23x1mrEmmnWwSAR2/OcwEwGAWUP+C
glBKQGsZazc/tkBzXdfXxtISBaD36n5r1dboFDMAxGfXcDn3CP1K2sZxbm5R+6Rf
4DdQruJOQNjY0RZduI+QsXXP0dXPEjBrlI10N/DOgumISNpAoDreNmVM6bn2ofO5
boAvcjIl6lIBzoXYIxQ22epfdilzetflNC8qjBVQmwRFE9mOXNKNxO09c4yixvOW
iyX98xk8LxYQkWWlEkdb8zZUnk/SwzRJEZ4G09CNWMagrETjUWJprB36I+FXSWgQ
qnHhLNU9APKuF36NzSLdBfQOGv18CPPhYCz8/0bgqeUjkVAYkVss3KR8rUq8pulc
WeNvT3wC3vPCkPvVNVeFqXH4y8hahuiL7gCICPtlRdxJu1Tby2LODMgeha/FZHsX
ZZuQYu4Bh10VhzjhGfdaLwLiZFFB4sYn7+CMr3Mw6GkyKVkXK2KVCRG0T/H99rTl
zYuhuVyt2+OaxtlwBx+plszlJMDw4tRfWj75OiDgt0wAxh0vJ4A44JPurvMUgMD5
pK9whxMW6sPo4m33M8gfvqKoS/0bjJNPl3Hmxubqs2LOZstvkCdoHWBBUj9/5hIA
2ELazf+09AtNQxs+WrWt64POL3NiyydoX+0s9RjBjSsOs8NcZu4ENrkQFhn4oT1/
f6Xi1JRNq1NXBa7+BRxqhISQ8C/sEAPrcN/4i8MiGj08NBigbK2m7cjOoKhHG/ye
b6Sl+5FA+ZL3u+9mspUf1kal2gNbHZZFzPW+Y0K4NS+zn336h4uZdIlRRTRKIcca
sXJfMLGnGKX/FAz7cPAesd5WO/yCXLW9p9hpKZlVDx7xYhfAyjemWIUNSpU1xvLo
FCmYdsG33/4kvES54R/NNbY0tw6V+EMvWNiR2JhZdftWzMwxkjf6XJPTnMp7FM7C
pvSFO48N8hxcxNV1BYOyTli/VR8XkZqs1aMa7g5Mgd9QcM6jCP8tjjDmjnziBMIk
OA362Ykc+2npu53EBmPNHPKuPguvMECBbDZHdzUJP4lYeFfPnXLWDOs2V3ecwnA4
02fu6PHmF+TugfrfYr0sF8u+H8vDtW6FLG8IwM8oq4CRZbWM1x+E8F2QnaTyeOUT
JcT3gsEG1GM7L0nxkNf87v5YjsV0FXqh8XkfN6QRSrGooWFk6y4c0xiijunYnFPB
vWcTq02kz5jH9juu9HdrXO92Wsq+xYjl/usNjGLItjxLmTEQYWpMfHghS1UNJb7f
xkupZs1lmTgy+mp0yBxgN1GX1HUk/FhvWaJcmy0AkPI0mvJ4RrpN2dZHckgazjwe
wgS9S5CsK+Q+pB3iJskpiCF4efr+MZVlqnMP7s5KNYvWcmWELaz0T45COvHdvT+H
AEOY0q/ok4dau11N+50olgBIuJxGCQ/dF4g2NPxYseIkqOozOu0Lco34kZW2Zjop
+HNZjhIRMsvwnIFW3PbhA//ZzKKd4OPj9FoQIoyJJ/K81j3c8uLAD5yDsvbEESXD
ujHQsvmkJXuTnDqGm+goCxEwMLlBr9IRSG+Eo7rvUqVP28tYCO49wzHe5TlIga2X
/GIgDl6LvEgGojtFMSyQlp24R74gv3C5CmpM8nC89aLy5hhtb/mWMnuQluh7ONt0
o+twe4z3MQmo43j7lN3ucaQPT5ra6+KMaX18eWVq4Jbu+/yhTEba1WfKC0n/5TIZ
dLFEZfKUc/6/abUoEoTr+IrgcpPpTD1kP9KZJuYKPciOZZM8+3ggHGhyxfiRi7KE
RQHy4lQi+KxYRJuhBEUGEKidZQeM/0qjvHBCRCA0x1mwB4R9HWDJOp3xwEmkSmuH
bqQ+X23jQWD5Mh6vlMPW3zfU30bjfXPSnEWGUOqHsWnTMHTa5hHGZcKE9clk+DuX
Rgx3eadRA8OmUftuw1Wowc0XFCSKrRxr+IojBXmAV4tmDdqO/defkHMuUoNAL5YC
Fmr/8rGhXFuEBEAes+r9D2xXQpIAWmgFXJ43Dof514KtYetqpH48eVB3956U1/cA
RObg0yW6CUJr2Do3RBRiW0pZFDhX7xQu3dM0BAwNCgfw0QqY2kVJrw9x/AXTA7YB
Ft/hxSx/2IBQgy5Ma2nAvYlIFU+2oTz4hPSr3Tqt3aZhokd1Uc8/6kr0rqDbYnux
R/78BI0wqZtXLeLzinQtern6ky/pjHk3mTsBroi5GF1Z2sWiUcz0AG5d49t5sgDQ
DCVHOfDjqqkfETn9QtfWJQ==
`protect end_protected