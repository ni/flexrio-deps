<<<<<<< HEAD:flexrio_deps/LinkStorageRamXilinx.vhd
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10080 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3Yu/9rPF3zgmGpaB5ZkBtHU
kEuSK6RotYmrmvJluUmPGT93qpfVkM6JkgelKbI/3JYb7h3uy9xW7Tb48n7A60sO
m4AvErxH65l6k6NFYW2C6aP5aC6JrY4ZlJXpXclFn7eQ8TPoFZDEFTPB1Wty8Vah
7occ2fqqRc8oP77XhG645UAV7b1dDI2vu5/OM7J2A6LNpRYuVUCneEOVrM5lQ+i/
0rMyCsgxRB0z7yKPYog5kdg0LzYuV86qYQ1cSzirKRlHYHLb1pYLRc3YZkL24+7z
yaX/lj+LFAC1vMaLuR3/Kojv43qrFVksqnbM7qqDISzGCfLrVk37Lh5hlr/3PJvu
e9KnzlbyDPsQJfjTXTYOHAiQDEdePw2mS8kE4m/NA17WjVFMF94z1OWu5Vf5AS1e
KuYXyLe6KtyfH6eXxHH8cqENP+FGlR1GB6MiaGeUrRixQto2e+bxvUwRLivcSTOE
0zFuW8DkQQPVM2OL7IN67Nw1nD6MYw+3o+0VYmaeLQVocq2dbQr9DFYpLWcvx93X
u5opQLXYNnk4ttrLOwZ4sgpGJLA7M93EC9kvhr6Gd0YJalPzG+X+7Gw44dTxem2G
2HyPSuOUOPXSzKzGZ02r9J2Dp/6r6Scm4sbB3GQEiAic028YxSxInRSX6pJ7RtPh
4Y3yPMzy2fMQLZK0SijqIUspyUJ53X13KR12sAcu3a/My1NIm9RbCu2ihLHDAvZO
IV7h5meagknDx8xWznIXCoR0rDbWjLWd21cmiM1S4T8PwBTzrNan8d8cr8BAzYWH
ByBJPdb/H+YTloT1WmrCp2UwuP4yyJGP/Bms0BoB0A2gZ0wagAODmK5PvLH501ah
Q/depIUqp+8RMBdgDk2et3q0euUMGWj5vLSA1hKAJrIY/xHaqO3TIksjp8WUY4vA
JtpLMDfvQPHA2Ojhs8tCffSJbrhBVdffc7yvfdSQwEi70SH+s48M7VXFksD49CeV
QSSCf/dYeWURRW9Hl7v8m4wfLUhZw6ALi6slxWLh0vPf57xWB9z+ARwepsa515rw
ZpofIiTzsuylPaJ2wHOiiMD+difCjH83FD0Q7nefDl4PYRkZy1fID37MgRIVPlBM
NzD/hO4a8xNaSoQ4TPaHZXkKMnKo6360HfKaPAoLF+uLlHlKB3kj5mAxopJAhLns
hAOJKMsPIL9jF7NKSoMOND0BwLn8QlDVuO1nbtgIF2/P3mOeNBga5W+CQu/VDMNU
TwoF8v6I0hpYKIowBitAVznmiwyUJ7tTsJZUuvQ/77B8hBPkXUmyAqZAYK8T2GHg
WMZZitXOlGueaBRbgHBthO+1lmddu7E6Nz+2WJIQlhwqFHLXc29DzMkvXeIirMwa
W05MFFPa+nEALi74fU6P6J8axAudty+5obKoS2v5r8yb3nx9NFLkg5P4zAV9rsrL
kEDssRBp8CkaSTIDpycKYx9dI1ny6F/yQe6gLhZ4+h2RERPa+F32Jcdkbb3Fs2PM
Jau1Gc87ZjJ3y1nmWQiqFM0Ki6azhcK0GdeQGlgTJBPkFVHPaaz9IZ8uUrjPfj82
WJEzcxsVyxVgH3r+2mL3uRwOpwSQjAMIDvXyr39Xz/bBz0QPf+82n1nrexFjpmvO
kKAGbhq2DNaxLbnI89EjcxBzG3Iroz7x6MS9J7WsD9uDCu9+1658Mzampid/nD9a
atdyGURgVmh3Zl818kb+u2HZxlNV0zPz/Wvc/i97BpwoLPFKw0jZTrIkR2kn2JeU
dfUUidM9hziViGWWXqj1xcWveBWpotRBB2isU98DalfHc5rHuiJWvH3vjwc773sm
qZCnCPS+9i79n2mHepRLZd42y++YZBFBvK5fddFMEFakjUHSWrr5eF80KhF5SPUJ
d8nzi/q3FFTLMNNUk2mLuykE5k3eKASEKFDRRwPUu6u575GE/f52W0u5Pf9wqUMm
u69AHLjK7ZmyCwbKHRwtEJYE+98MXCHsm5OMdC23Mtj6q6lW8X9SLXMD2PVMe0xp
oAh7aSqXf/Duj92N2Q+ZyCtoWuUiZca8iDsuXsWeKyocCR8IW1c8pB4FyZGqLOU0
V2mwZlOwfCkghAB+XZngzk9PodiPapgMg9iMyi2XC+5lPjDe0dgLlngFIOHc7Rif
FSJdZbsLTMxGEEC0EP79MAukJZiCpn+iVtnPciawIapAzGZEC0y688xFlLXXS7IC
6ywZ19kbvkn1qzypaR9L/mBMKttJ626XOfmgWYoj0ehhAJcPx2FSwc+gdlloZWn+
wj82+v5k6YPFPMDhJD6idMwTRwu1c/2N2x0NzCrm5dbzY7eWy8rwKAqSV8Nfbdvj
cySwOfJcYYcPOC0fyAAISOfFoNvyhSpbehCiaezX8lj0316AgQhFp4s+LBhHSxaZ
mq2Qh2U1Oy6EHnNQKUz4HwSH9XLjfAQdRHJL0eUjeTztUFxM4/m9hZUzGVbh3Y1h
nhR3MfdqzlFcyyaKSwj5JlhNTGHBgox7MYN8QouGY2GOoM9j/bg3/p+bV+NPqHCP
PCYFnGWLoU/F7CoIPmaOBrsVGCipmCv0tuINIn4tJcrZ3ZsKDgDXDZHZElduhNnf
FfyAXkJTmTZ8pgOvpk7Did/u+DjWo6IMQFCum3cBgC5vqWHTX3QkjHeetqye8BHt
r4c4NtxJGDy1TIMYVkxrFJ3pByjwsk5n0SwKDotUc9X6a43P+k9FWqZ2N46B9sTD
f4RosR8S38AGuxJsF+8Qorr4VIeZJPfcYAyHBT7xlhHeUGCNKlcqQiOu2Zw1km/S
6FVSSayb4CwBBYKA31Ngyjt3xzNLgb63v/ZMLEtseLKdqRXV5VJxCAZj76QZYy6q
kwSHhdUzMGmbzeuVMZVyuUBHv701bEiUGitqRz5Vgd2Vt6OEg2DaU2CRpbfcYyte
o6+hlAg5uMhoXdKYN+gKR6hgsgTsctkaRcyKVzfzq4oRqPSgo4fQ0jdn0G9sxD2p
2xh35m9kMBCsjDIHDcqPLiGTYX7jzLKmDsrumT2jVq+lXrjkjcpBGtLnIAKhxSQs
Mk+kFB0gcj+SiNWbz8FzIYgi7fzbhGnxNtUmtud80cCb5JI9k4N+sCqu8W4DfTgW
hypuEnwvOskGhvUrUJJKsKQ6iuNebDOdmbjLBymBotfwdyPJETPlr+cDXq70O412
guEp8Tq6WhxfnaweYw0ZfROLXnKBEtaJk5lqCAWyDQx6lqoz1u24amnI9zOLdQmT
MEnYENPu5McyeAiJfUFeUQ5/agbCsWdvHgRxPvD0IZNzfv0jrUfbq/QDJixIoKLz
KjDd7NThSUXp9Q+QbYgyf3cOZWQvn5Q6JwlczqlT3OdYdxAsB5SF/hoWf4crxu8p
/2U9ubftaM23MDehtUGBz4TkxoTlyMTnbp1zgPmk4LvlJm31/jYUKGm1oRoiILFz
aXC2HU7jzpazOWM0EFjJ3ql7Bo7LwbXsFcTWrDT7mxEzEunZ+pR9w0xiShJZf3pJ
YlXpn6ob9AFPZBVYrpaBuPo+gb/X0t+NCidIq4cxJ8RaBQeIB8oUBzchpffO8a2Y
f56rGe+UI64C8/7OpnV638Wt4A4CWbFpJxK1T9qO7/SNMwGn/XcC9j/fscVXfuM3
QP/IJk9K+ZzcheDI2Y7wg6I9jkYRFXwNvskrGajDKpvphMpWAvRc4BdR5M86Qb+W
pAA50XZ6ZD7KKCbWqAv8iNkYEmquRYncdyI//17ULYQmwOX2f3r9r7P9garOK86Q
DEDaH0ZS3yW5AeKdrylrXSzjGMOT45NaLySxyOYS+wncA/pkJjB/9ofhqi0/vLOq
6FFLupD6QqYHmA3XKpDdWvyVSJn4L7kXYmeQ7YRr5k6VBg+Nf1g+1ujw75dsx7j0
dX9tWUZx9dhxTaOyibMuRO+jbtAEjW3qA7ABRv0oU5uW1lF2llRFS5NaYcHd0TJf
n4WsT7VCwk5F8axohQB3kt5kf8zo6Mu4L/qRr8MbA48DN0cVviuenVpQoZZRoG8m
5frBAScBwYEdivMYnC70cLs0TW8YJ2QcK7FjMZM3ykApbCmo6z60KNlSyQn6jUh3
8A7ImBJHru0mZHtZFSQWfogkx3srsi4yh8qraSkG09escvIiK5FZcS4e98DL/Vqu
Rutvgmaf2es4CDK4i0oHfQZxpYdR+HvK+SOvXiunZyEhglBrMqVuGosNhNIC8w9A
G/u3S1hecBb71vfKnFdTBuMC6P4FpTUma/LVwp4qYqBD2LfUtB2t3LZei9GSKzGN
QWHVNqLFuWNlwRTSLiE/1x1JwUrVxQbTpabZLP+fCDvc3xnkFjf4xsm6nqp1Qr/m
gN2lwpoPubmXdZXrJ5GRZAZZikKGrvwshn9ON6T0uQNKWe6T8hmqvbT62i3wY3o/
r3XNWCIWUEvFaexOu8YxpLeEbHObGLwTdis+PUG+xAiQA35T86GawxtZp5C0H9L9
YWZbr2ygD8zjNglWOK2A4zsNNKNdLnevj1ELO7TSj5iTHg+EqNQFXsVmnDnxz0Ng
qHBC050CCnEuEJGB2ke4T12Gb2o/XKk+4/sRYlTYNZdnUlbMAmqIP4xN9FpiaBh1
zI5ep68M1KixDC0GNEwvoZ9yDC/HVwbyIWDlNh5d+Y1hXZVSDhGN/5pfrT/PoXWF
RHEaqvYWZV7u6PvgaLFFxNCzRrUM9HfNF+aYyTjj/bxG9Qi/Ww+vU8knDTREE8/+
OysyrYisdwxYWgnDATodw5D9L6Xhmr1fv+KKqWm4y/AWmqAJP/ldm141VI3f0HKu
aEkH37uuY/AhN6UgQf7edEvpMed50xuWypu/uXiRn99h43TQtL1VPD8fOn/rLGgR
DEK0pKfoWeH5CAlDzjL3hSlKhkY2+fhI2Vy5RNmv69PX8YmnjVRr/deLHkH42ZHp
ADKpDEgIGLh3lnr0/j95cT/+C3Oqmmiu5+Zx8i2C0qd2LaRq5bMMuuDikQfUHDM6
CPbadDdKXPC1+5rwGBOGOmDcpqA/Fpc5KV+Dl95UnaRoBA1uiDB4xvoccjDbVplN
ED5WNXBx4caCbitqkV5QFwUOiqI0V6pf20+XcGcSSzMTxZTBuGoaUYeC/Qo4TwqC
cR+psXPBm5TsLHsbaJzIOkqDL2ilg0Jen0gJdEk5Tq/F2otqsErgJgWuguU56rb2
pGBP1SuR+ocWLhD1BSrfDWn4/xmLbcNAkKyb46bH3rlvBMUTi+bycQwIRk84hTkm
/lr6/FoG7S/VoIFAXZtX11JEW3UrS9gcjmzGUca875PM7aUlCaDbOiJU/DHyx+gK
ssXwoo8vwp3nipDm3Jaxm3kF5Z3GV1PCkzA7riNnXlElMux+SXjrgha9SdKWa7Ur
RTXRJW/3dM4rveZ1nmmmpf2hhLn+V9oCxMQi425RzVQ++bCRMQ3LjXdDe89L/5P0
Y0JGqojLII8CsqrKr+x10EN5UtOoXrjZEjQxQ1SinlOOxHZyGPkYP1B2eqvj3MCs
Rs8LfBq2IaVIyPuNwg7Zzx2DtTbtDtGGkt7YMHIjGZSDCDRX42Bhq/ycvN+SM/TS
B9N0BhPZfmIoY8nzcfvfgSEpgoj+HS7TWuqEfvDsAzJHi69icVZ5/9pNgk9VoTFs
p/M6k6wpMSHJmqmHRO3ydxcNLBTUsIyYRGXknfi9zx3dvdZxLNT6U0fJ+9FCWgHz
6smarTxWNMHQrNYNoo7RkOxlAMRw/b0CDysc0z2Z/Xcd6QGlMjYKqoMp0OSsiC9Z
yvnYvrF1mvngvBZvn7HzxoqX905fj3eaxdzeW32yyNVCcMXRRQRvAbY4olWx9yCl
q8UXKQW6Hiti3+JnMYOxfSMnSQCi3rnjBDW/XDXxCZQk/To9ewfz65MqqVqyiN5f
LYb+36qxyDbdTMKNf14GLJJpMQvYTGTZZ+NRw0SYH2tar7af74hwMl5dBDC3vt3Q
MAKsifgdzvjJZ/Mo26IbP68PvA7CoCMXd5BWmRfSFYc4aQgbU9+4+iyWF/vrP0nd
jXZBeRg5s7eVpYOCjlq+fd+6kUlgzrYydQ8OR98qFzKuhKdtgJkDFNAYiX+zzGbp
+re89cMdpSxu7S0gqK4tBUVdDvZ8Jqj/3P9wOdUOUggaZBD1HR/5aQtbp38i7DiC
syOD818m9Jo9xcCH5IjXvxSVebRVsSye/X+h3++EzZ9R5WTk4g4ulzc+NTVoqt96
9yoTEfNOhIBLqVnNTYj9Tltzj07d6XdfdGROzblUrg7Pg4Mj3fX6+HEkS1UeVwSh
dOsUC/S2YQ7ljn5JClAxi+mrO/cvKLTYA2YiNcN2lRL0bcwpRiu/B6oBU8xKTE2U
8i6iYks4hYW+XLt13FpBVH7mnUt4r7RO1cMyW5nIVR9OBH890D5acdzxEUw0TqKt
/bQNmy2G07xgBGY1BFZ/kbO5z+FDdTZFGeEIR22mLZGNhOgKV9phaB1wvLgsBBya
Ss3hMX/gRYlyNiMP3w/m0tzoT4thJ1P5ZkDGEAJDzbov9JzSZN4KevZxMmBzSCOY
cIOk9exEaDkLl+bp7WEySvvemGxH75sKyCy8mgqduZEbHVXsDIIOAj69W8TjsN5F
pNkfnvoP1uSvuOx6lOby8MsDnqH8+b9RYPf9lOE8vms3d+yjMdwZqEEX4NN+KfnT
t5B6rEZq1hmk86DuuhytiD2CoQR4pZ9JFblgG1+W5R1RVmmowB0BgdmlTajF1um3
yscNcQiQprCBvAw87fcyRUy+icMPsTH014yP9uYA6Q5ZNEbTLYHoCKBz+vSfN5Vu
6XusYxSDkSAYW0v+hi/Y/6VMUOxI2QU4+P3+VKJmwDIGqbJ1dW+y/6fxkZP6tKvb
RyM+ehXKvOieBveJmZVNZ4yqNu5f0zPmjJhxCS274x2NgUWLbQL5epgjUkvBstmn
PS55ej+9SUqfQpN6Tj7g7wh7lY7euWhNLo453WrU1WGNh7j/XgQ/nmiDF05lGzEw
F5qVylCe+RzqGfhyzRSwe+n9b4sv5A7FkTRTEMPeTED8SFTuaXC4B8o3t1bIQ3Sq
kWrBSHYGBJ8Ibj80vD4TAAV+BDTs9AyKKKYmtFH9mqzOKk5p6o97W6NH6u2lC6OT
x2Ie4rU+PE0kZShLy+V1JZRUGIoKr9+j+8pPWxoXT4l9Rp8UR/M4Rei3DZyga+aO
5I+lYCYV8FkbEoaTLqV1s4HWtPWYp0i2tc1HnIAP8GEHjbTUohV/+wxW41nFmxLD
tyAq7Z/McYC5b9eQcs6wSDNId2Y40lXiiEtGWrACAzSrHOekB3p1zmJF27cU5dXR
Nvq5ASqbNEKVL4Y4r5Z9xHNny8zd/rA86MDWPal84AO6QOX8bV/TZYnmOkqCw1FP
D7UEI2f8qdeF1pD4K49W2wOAKOTbDAV+CKxso3JV3SPrGsswePIdXu4H2SgeJYVI
NLOa59MuXw2o8x7xOPMCV5GUqgVTpkMj0UAxRGKMTP6051c1nb9qWnJo2z76572j
HInvtffzZPjndVbGrOyFgESyjPfMaaG4RUFoYsPFKQk92/btX9kyuY6AAQhr+CEF
td/Fy5D97mJMx2R8Dhb8rMc8zX+0I1C8Ud+BRRGeEQiqMrL97pBLjChv9ys04PAq
7cTkGtYqnMkw91V4ubTePuHst6lWyoYB/xgZaimzsmswxuLA8e6dATaOoPbpUGgv
kZMwc+oNlWnnesTCi86xexiI4Q0kU96cYJpSGGhfCfJ8l+XAiiZDc/XyVU604wNU
qZHo7uBR+zxXqjkBk4VSNHey/fxK25IH8HMkBBH59NedPq9wtK1fufy9CdG5HZnh
ZL4tlTrBAEwBGDGUIf6rN6xG+10Sg4vCvRvXxB8XR1UPv5gySXIJ4CZE4BCBTNCp
sr+CMJ/ZqLVQlGhIuNJyJsKcabzssDbZA9q0pK+//bZCPzdmFwPPvaZlRYpIBTFs
yxxIVGe4URobYhpDRv12Z6dnshqXoT1fDsS2HN4WkTXnctDk8kth4Xi5PP++GQoA
IyiygjRabHNXV5s1DT9WF3LO7iZdFv9ynr/QuKWSelCoNVQ7N3mGJXTZi9bPkE2L
A6DUjyM/twgFEUEv5QZL83HsLdcJ8oEE123mCuN9AJ/SE01Koj5cqPIvtr+a5q+X
0/6awRZx0KYTEv6m2RmQwNrOa4vrUw850IodmT8RFkbv2domnST/S06L5CJZ+aO6
mr6larvmo2r2as8MD1JCk1HMg/Ju2CXtXuSmNOpwQAGix2UQ3MLYb+Ksyvk43B4M
4vn4bfDhfWV8xyL2CMXsaXtjTAT1L5EYCXX0AG9wSJxJtLrzu9Y/K37ia7UGTOYc
vGkNNZu71mh3bBWzB1vBS7t9mDL5YBijl77cjMDxfWcQgv+OMslc9vsoay7AC/RC
LUYgseNdryT0zL02iVeoHKwNQ9XSUNbpVpF7ooPzWuMZ5deXzxKu8JLzbCAr2s//
e0+RgI+tl+4JU119vGmLB7NwNt34IFbpYiSvu2/zraIhwGVI8L7kgx9H0tzsmudX
bn0OO6seZIIUo9rbbgbr1y43n/NmHPM6aeVkjZW8hsMan1c5ViGlDXtLG8Z1NJRh
6Dj0Eiv3f1JJnTasu49cVvac6O/X4JvOt1c47qCSag3CvQpfK7qkDldMH+qKRful
vp54TWO27e3Q44LKq7Fq5umD67mp1JswVKpWNtjb2rllapSuYV5rgAQHniRsKerZ
x17yzlncGI9H+QhbxRye8NlbQ6Mlte+/U52X+xePt5LX8KYgSHsvKkgnYKeyXxTU
9fTKj0z7QkuUV4rLjHDR6dxxjcIR+gNEEsXPPE7ptPV+zBrfxDAVXDXqzZiRmKyw
3n0YCBYErc8o+TND6+4FAtWlCmmm1WLBsTnLRNJ7jghpzFGwRIGcQU6hsJwx24Fz
8ye0ffOGuiLtYlImuv03L6n1pbOFwwWVeKrjXVUzKEwUD/XLWHDHEYIv9JysXuSa
38InENxiV4KAWv7/CX1gH8jnvytIki8cAfvVvdijQVbMZfNWwfWp4ITGcyRfSd4T
SnoksnQup9hoGQUWrTdoxmSOm+CQysoao9ZT6Yg26F7KYPbmZKw/8QrV7ox0h6At
JIC02HUQhnGxTC3ZDWzdlkq8TfsFAOXKbQR301qJzD2uLxDEbrTXIHc2oxE8ci9p
73vIcCYEjRtBfTu6Ivi1KrB1ELzjc4pi7MKNSN/6NPSOXnu/uyKS9LdS4OvTRU1W
W3ZVKhBFaHcYO2JMJmIM3IixP1E8yoAOcEyJY+g/C4Q4sKB53oue3YLBL7m3UrCq
XN2LhStYyT2YHRM2CSv+bd1xODKwDqzc/iUuv7k0+HR9NS7vFUE2jn6tMzUUzy7U
0cKGJJd4faIPquMxiV2b/F8RsxdEpjdrM+KbMVoCV2E+rrrajpvJ9x+SS/TDv5Fd
GvO1VHnk/BZAz2ICYCjjPJs4o+tQtthqukJW/iQE9eugVrE6Ff7c2ctyh8AkYSOm
WcBCBiXhqTyVcVHq2bNkFITJfi23TV+ZPLCUPOwmJZd3b2y4UUk+yW7A8tgN7g5I
Lf0GzIu1FyYBKIe7m278oC/jcJeS83rJPZASQacP+Sq5pU3u/pg13h1i7lBvvO+N
Y/Et3kSurXmdDvn79JnF9lAmWMPWwDKYeRu5yRAWFsuE4gQs0ehf/tt2tADGPjqp
1+bobyn20FImbX/HnWBVgNoBJSzCAtIxq/+obSf3p9L2xsTyuN0nPoLluWN1xgkt
7VkOR63XxzL19GuTPBOzLdhSs/mRB7dffDSPAjq0lAYzz4pw2tfTXTiGFORxw6hU
TwGCL9CrLocUDeLlXO8dKtdqbYVLoXLdFfnUE93vwcTC2AxfBMyjsa5jdICur9iZ
CjzXSIROFiV+B7FCFAByiCkEMQBTt0VsxUDqODmr22ozu8oyV9I6YZsV//kEdPXw
N/PXyWTyRXZdzsUgduRa+Ed6NusRZhTArQ1YDzRxajYsiexegcKdMOm/QdS0kEcD
2rbN2A0V2CsU+kyxrNYXaUh7RuSPZMzOaBVLSnqXhko2McFOydKGCeNk2n4loxDN
4se3Bw9OV8wKKzvF2xSwwu169H3VVgp90gfAg8WNKgYSn+5bqLnFja759whuVdSF
adGhoCQgDCnoS5nYYF1dRWMTvgK4tB70D9nYqidlMd9qMgsX+enJgXUqVCWnQvfX
LadYDu0bU0YXG6ydaOfxQ+NHoNcfTgqhEicujZDXuD8SozwOUh8Aj1e3RHDt8gaB
kLlUPxiITHaQngNnQrH2vZrchEMX68Av6ckQV+XqDvHdj7IfD0fYpMFcdj2oq2OV
oR8H18jiiJ0ohzggMonOeBRBECv8fu0n0TzXXpDlQpbwonkSWHHoD7xotoxbKavC
MBGDzV64oAR+SqXlP3LAe+Mshb9rlHiww7egDIE50tgjcgDgHdhoE5pGPZS7OuX5
gNv3Yh8QhM7Zw3J9ytSkCXQM3BI2yUtxGzd/+Bj2g+c6qumpdx07PP3D4RrXW7lT
F/JUzJxnbdUceVdpCdE/O5HSGrL9ckuFEGZyNZC6h/gtJ3FRqL9cioXwRrSzuXRb
7jqJWYOwyhdavjqCyH3bwAgG0Q5ZZV2QPWxgv3W2TqNbQQJr25z5lKnW7kLACo5p
Ky6auuCFTp9XxwGawpXNLkV2ZSa/UgHWoaxYh0jUgTWm0zJx2QK4CTClSieU+en/
UaK2iT40/WGtgF9rnOTIFV619m9J2oavgk2wIecECvOePiFN+PrFw+XGMOf6MXiK
UtNNvPvfR4KnyTwd0c28ZRhu4sg8erTE4AQS2LPC0l00kqBw8ZbB+S+EBa956tcg
JDfsXbzhjvzmBaoN9Q+25Itj6hMzc1sAHgdThTTk+J+SXCZIPitytUvVlqCkBIH/
qyNipnhkG4wTWcLquvNixRzAu20yg6lRivANWaz9GNpLmK6Vrz54vc2XxBw50Vto
ZFsg9N4fOxMYod/D3gT8JuDuqexRxF+JKXZc0a4WGKaVS8TpWm9qv7yCAsvQhiJ5
6w1Lb1sGVbwr2vaTGxkDv6TcvHzWqfk9Ab8FNUtloDRfQ6wektJgnP5MTbUTo0DD
kOsq0658zfcZJHBEkj1s08XMt9W2q5f/ouEAI1ZM8Phh87BilVgnQw70fGKuEqSy
BK5zSmXTd0fXAN0hxhQ3C/Qu+DR5Vxv8MEMjFCb48uFbaLfZm7zRvp1jdbcpbz9Y
6A2KxS45gTARK4liYfUN9gDIzAP8cji/M4q3Hb3rDMwAvPmSv4PxRYtVa6oVNxJV
1y076zvJ2P7ZFf9pUIz7CwlK8S6FUKwvUTKHLaJGfWJ9820ShovX9JqOTgGGA+yT
orp0ws5GPyAekpVFtg0pwmRQXsgzlOBNnK5/1u/X0rG3bZdg5BG9Xv4/xbsmH3C5
sW5tESpfFwF4I+xk51ah8ZeUwX1JVxznEwFqjfKuhdm60vfJfVy4/SGGvl6LRMbH
UK0nmSrneIteKWIOrdPmPI4hmPZEWWeEs4i4xzsF7tJT+nIkCgordLSlOSDoY9VI
89F0984FEuNwuf3q1JxAfZ8SVO6AG1GS8a6/i/0cSjGHC0tSFEJ6cDGPCvfwzeHi
NIgV0gWCEau8IElGqWlbqP+GupSErxgbdknkNAVO2SMnGJifihyxiUnHOIewGw/c
ZGAYHl8FUcoRkzUN/AwbvQlpcBRK623NgTT8yQVeLo6coKv4JPa452nxx918rC0n
+MNH01W1LdcgP4dc1WF2y6FvZHT0S4TU5SIJnQZwB+l7rQCUky20CfrZU8XnDtKK
nhxVxda4C5gIjHjrhQHZIdzLs/hiz0nh7hsObeF21XrawSAD0pMBgYG6sIVcpwTD
I1XT/5ebRVOAgaoG1RNqV6DvLdEcl0h5eulgnRwjWWOgDGbB0XhWK1dInAM1gD2m
YKPrLiNTHFzBBjiIEmKVLJ7TsuHBpj51/fZdsmNUBVcwWm1vNNDh++TRMLij24Je
sKUP7DA1EoT7w+9wRSfz8tHqZA/bMjwNHpuKNQZ9wVdMLnH461DqT5yrDXHDn+vQ
LmPCIjHs7EST8BXuxJGxDOsd9g8TpGS2uTLo8qkVc9Zx0b4HqMRjO1L99HivcXlM
PudYSCBodwRmgK7QIvizOtp5tpAvnXFOA1kA2J8Ht/0ZTyLMxxxfff00wDVHGF4D
t6sTeKXV2xSV7cEuSZqGeUu9n8SUu6E3x1J8eMWBqcUF/jSN2liiUOaL8Be+6TjX
Mk9PfGmCKoxYjs+fmnkwStCUXNi02jvprB207oUL1hl82k9BYzgbTHwD+RS6ju3o
Rq3LQoKqdIJdmOAQIRetdIWQ9YmBBuxTcRuNULaWCQMciv6Eplz1FP2Wba5bCu5K
0rwZxX2ifxe4N/jqZ6CqzMVj2DVVwVR11Bbaon+5zjgJ/bH+fiIXjcbreCweBglP
WEKdsEVZZcAUBZdhaccRSLkXRzLJPuoE2bD9VyRZIkUZNiK9n5i4cyCb0jlT0GHQ
SFKGbXuN5EHCGoM5Tua93x79CldDuWsOKtPTlbCFpK+h33ojp65z911+o4TNQXuw
gmnweR5BPqhK3uXdUNfS8+8gr0z922V1r7XOODZQToLhHtvnPKXDUIh4W/JoCJjI
xK789wKkqJ3aiXNzw7zRGDn9acLYNpllmQE6giLzPFpK/5//oGAV1da33htyauph
Np1MLsCSzTUu+mP6/F2o5vUFsWNBeYLEpX9zUeVaYLlQWKOPuOz3iLgvtmQjSTw8
vURQCoa+6rw8G5MZS9hY/i5zYR6C+1Nl7PtcwwpxP+CRvqffmt4P8N2TwP5KiLOL
HGK+47fsU11HrltuJejUJ+Cq0G6mtLVZIJbyGCe/eTGxTUD4xuczseq4Kw4G0zux
XVfgFAMpQYosjNFgMhwSvMFXlZReIL3tA/aJapo0HAN6RkilT/3idKRr2rZLx9Z9
hMhdkwBzpQwYCBvzsTSouC2u4tsIQUAYbeRq+IdGovdJxq6pmDDvsZ1L62XrQ7Ph
ruORGd4efuqlRx6xfcbEWESrSpOprHJ73nrI574kbBpOy0dTO02MyrDVBHliX7Lp
LTwyvoUXK6ihXUnBUgpx6XLom4w/NGkNCXI0OyT6KqsHcfmlEGEK75GsdiLRdnKO
EjzoKXxClCz4u7u2pVCKRd+6isxmKHK0O8SgMsZRTS8MM1k/VU0hxLWd+BhJPJ8E
qrzZ9wQH4hSFhHORpAT6MJKWbQvpHu9cUd775pT9aWpmmPIt6wVz58jj3qZw6YaI
+qF0TOyRodDLsXJglW3iEdojGJ4ZE2LF9YvXDKgDJfEH5Py1ZJJoKm6kKMxWXkSx
zzRzywSbAQp6kfN6Fm2bYg02WNZ2rru6sDElUshqVW9ApWJM7s49ZGihJGdQ5iHd
=======
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10080 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JWeJJ6Ze92g4+4wPuytvzVq
BUiIjW6BqLMgOdxnHw5DNWEQW/Ew2db/LEgoa101VlQcLbk7zrOOSuf7jO554NkK
LvIZzGhSCaoZNdRsHZRGRAaAr3dJqHoskhmWfwhLQa5CDYVyj6NoaA3VK54CQv1m
4lbpNoVgLNUOqrthe4uDHYBmQgikGIuCPGyij8/X3gXr3CO/EaUx7U+EAMohUAYy
VnC0VN/dioUoX89iYiaRGS0mnHSdpcLmW6s/mFKB+MTDaYpGThvqo/q6AzUiY/85
+CcMQINMEVGsOQ46l3Ly8uKIB4ZwQ0At7yatZ3Gst1WerI4nvaUJtb6TI5dUyQT1
Z5W4MvyMWEm4ePGyXsavkPfyjHU9Wn4DgsZBWp32gmr2Auf/6bRpBZ1sjduD2UIW
1p197gsIbvpyfW4r50agjE8I+S+aaSZdhM2oC9fX39aH2GuXhdoFB2U5x/IvwuJg
tYHM4W52EIp+1/lakcE0fSg7eaAaUX39Vg4cyRdDgcojsv+4rVF9EfMu0C9C+E5a
dupKyB82730J0xvCqHCxfTPynZKsBOa/n1ATDq7ymIXqv+T73ka4nUKE6eeTD00X
UZH8k+dMc9Vz4bq3D5ppSQwo5E+O5AC25y4AaDI0XUxDUNXyD0jmTwaUSDKB985K
/wFarIERcFNochNomsM+UqkSgRzT7S9xG/od1REFxjqz3e/PiZS7OfRnrQaKdFoi
VtRwdDx5XWcIHzX1NXkrwWF90/laTUpwTccIbdEQTBiVf+qoY1OI+z1p0ukAY8IM
4ejubMxHcYyrw1eGeZtQW+P6bx5tEmZ/Whpzyv3/xDB/4yjFv/JpHcPuHLUho0NG
wrLc9YoOm2GPzvPuODqGlLsk4GJwOpDny9bxOiskcYIXQoSZsrCWpd0wyZvsKDbJ
7BGJqQmtMXl4oiqYE3b5YwPhmfM4frX7ce1XceFwzGl3mhSCWq5LOwpoUTnP4xLT
VT4KcI1s+q5KGCfFCee53pISkEXhACQfTHlb4g/YagW+WmbeGjUL6L3MHqGuT/rU
evKf46vq5t3tN4+hOsJ75kkUDfb1CBSfdI6oS4Mw1tl4DaX3jkQVM3c5mn/cxNvN
GpaQeEF+xDJYTi53WsxmmcXAobQb972p8BE+XtATRO9Ylta0PDCFR7zD5qTbgdRs
oRtnrx0WfZrD4Ppt//wCR8t3TK1GDqPC3PZyOKxQMycSym89/+3YYdQSkqiw07sV
vfWYcQ7n/sJ2YkYaORyzmS+LUDaJpBf9EunQ619EwNhqtH+2JrLzNo5Kz70J0D0A
83Dg5701JsOPckLybF9mxrrlijSBeG46I+E7icBkg1KXeY8k0AJTZ0H+3zoVF7zA
KKQ8LzJ+4Qv9wYfUv0y9GboGL2fseViUutm8HOnSnh1OAnWB6Yty3oAXGKob/Won
tbJFsWPl+bxZQ2A8o+A7kXQba/hKYDOmQeKllFSZCk9jOj/a4BBD5tpYVdIQzFyC
xA9/V2RpTQeW8DC541ToNYiRc+XNul6TymeuZW8GLf7DAbvDGaI5XMTQbms9MeA/
y0iVNCcR4SiFPOrLHwJ85cwPPuLcsKgukbmr0eXN0C0VFLhb4Ya+rVcznIALz0bG
3VqnhLGKoF8I2Q8wdsNb5StK+Hxlsw3IaIkH/GRcvw1A4hmJkIcn+TcdSSY9xUhH
otzYnr74lI4xkG9Z23VYUrk1jUCG3gsvB7jntr3zVc6a0BjYXdmRStnpVoVLtgym
XDgd3I3sKZb8URuUJz0/UxUHMlobneJdrMi05vzomXCvEHwqwGhj5Q0czVGsSpWs
dZoSPumWJEtBGO3pu6d/Uomvg30YR74x6llRnfFdi57Bxr/GUiM0CkA9IZ0N8gU1
lQpfnMDLCQpQkArCFhyNnQcKT/8T3iWML3mcAgWFaggM7YAOcjQBpCriqnCmLw8A
u/u8fDfmHldZpaKfNsBiCMBKs25hkshPh7otlatxlj398iN0dAab0HfKYsgwhM/e
QsS5/60btmkMZRX2AFjH/oo3HSAm2Wn5s4QdzgIiZD0synKyl/Q+A6omxro/rv7B
h+h8BE1/N88C1pZeVmKsZW8cPGTZNrh4V2dmvjB9RLzCR4itk4s7dgvIZKd5zKQ1
GEdAvxqvoRjsCf+rhLDT7OfAy8F9G3ojnIAy76GJrysTUlAkE8Jp3Vi3nou1ofci
A4PS/C3bDZjDFyGkbFmOuNvvNvZHyGIA66qy7fUckZXpjtSZ9ciurZZRfN+Oykbe
U4oc4XLBbF8jXPbQCqR7UzeTxiPDKj/IY2VTss6wVAsmfnzGZs6IMOuebvPYb0yF
XFI0oIweZIhR1YmY9Yu6504+UiNU2NbGlyFlBRTBqSYGweiPrGinh6T4Wf/0lA05
rQZjouu0fpP7RlRC3xZFrnKK1/qtD8lSBXD9HMEuTEAOT98mNoS4KdJcQ9syiF7V
Eki9M+78kcvBvGi9ATHZPwfzaCOc1OWb2wvnBzgD4fQoPXzg+tHBLwAQ5JYu701j
3jdRB5cclU6HeV8T4C2UhpBErNuUwkdXukriszR+m/sv4/A8t9CYjA+ovHj5zVwm
fPP8u1TTIZynMh+Vv/KT62roa+9NtHGmQB5/cml6YTm4TZ9pvUmA49w7fUfaTzt3
JRzIBA1Y4FnXGSD3mBvBpwg/v+WganuHXt079s3EDhOf/hiNb1AeTVH0eufvLTv8
yuqRU/aArm7BQL6HPs8SVewWTpUYa0VD1q4U/SRhqxzvCk2gzc91QcNo4dSJM3vH
nvymp+o4l2ZSyVBiXGr3rsqCCr7TnGym2Z9POkE2EI4VIYmIxCtaYouhIZyXn2zw
PgzBzYIM66/GOS/Uu32SNkbmIhd/kHw7vawCXvtQpjCFz2c0IBvTkPQq6kAtSntY
9wX/yopHDaUN6U7Ae5y3EAzKr/JGh5yFgwVFw0pcm7IyHRusa8+MLr2MiatT+pOr
EQBEWXjnK2DlCpsg1R6Z25RDh50Ahqlqg8neLGrVb/B4xORgIv51x68VQ1rv0486
Zczs3WbbQujbmHhIbyzRJ+bLRGmJUSFUE8YiMPmhcxI4ZSx2WQOTeE2w3rJ2x52+
jG+a+mvbyTRAt2oMvDw5J3Fli5ws2jw36Cn/umOn5fMtiehvrt1FtjKuUTFs9YRo
FsBTbNnamGpnYPjDSofms0Ifusjr8Nsgb70xuxlSLpkA/dlD856XaBYOWgFZXO1x
XwtZI5z+tq7R/c2ymaBGYAypcxMXUeySmeZ8dv+cPZm946vmDtuYdFYAFlmPMqAa
Fu0fvK4EdxKgPHVZIz5KHJP89lmDz8MUH1rm0FQUcMmGoTHIVTJBRWJiKS6ahs62
T9r7AiOzVXWRVrr2KNsB3eOt6V2Wh6gsuBE+OfS2xZsOmB/0OCVYUy2NttPMUd2m
eek3bpE/mj3rQEcTi4kag/w/0MTPGQW0L/xpZMAKFdsD8FMyv8jHo436HhU87ygh
kbRZdiTuUg4Tv85WV6GQLHcs772nDHlS6ppJOrBfNfKAGp8GVti+/M6b9q6LPrbv
KPJApT9M/9oVL3gOm9erZ21gaIiB60kG6cKVK0ZOhpZ5jZHDihMcMCNWwRNYWvcy
KzrVArLdktp3O00mZmeEOrYBRZR15aEbLPyi6FPwi6Siyk4lPXfEV22SivXa4/fx
72xLkidedpTB7YD+v3LleNYCLvRtxzKouXwfXf8Ht9BVX3C/uPwvG4k6yLqStWxw
EMVtLNfswZdgO/vTbxJnNhdaSEv2Yff3dw+3xZldXZmgxmuNr8mo80qc2ECnT37p
jq8kSbHIuZolvL7ZT+4hrpJBaDl76ZlkHQOKG5lFFw7NIUUWDZDkkr1FcQsGmXy8
ZQ6I5Wwy/hbMg5xB4ynNIRMZr1gfwsVF7B//EtReSMC9LDLIRLkS6sgTe7MC/RTC
umM4BO19A4N7DvFQQTanIg7sFZapr8fChrAmQQ05dXeFBtIRuEbBnIk0o2/XMWxx
CY+VFMtGCLfTSBKiC30Dq8mdbHgxIFWi7n7+xLQcY26/b6D94Lmvf8w64ecNoh61
MFXGTJRd4916CZN4sUtf4pG8e4Zee5nc9wSvWO1LZNL4qxOLHKQ8GrwdMItRjRkG
aqps5S5k+9hD5urrnZjHRbrPe5c17PtXCsxj+McCoiCRvDxgbYHR/C35aUUJ7/sv
PaEjTiiS4dovqDujMe7+xYXKRntpH1uLNnwqoEkYMaU0VQcXzAvIXD2djLjjZIAR
QOPIrWUk6+N4uU9ZZmRXpKDMRaXBea2xCQvyc2YuNyKoqXoIF1MZINwad3S9txXU
HyqDfK9RYRBhWVzHJr1GQxibcQnGA0jhsaF2axDld0ykzukGfeF5605EDSWyp22p
rztHx1mrKvXEJ97OOAUyMcTtUkHDHcuPgEEAilXnP2IJcnq7G539bMUc0uIQzk6b
dEhGiN8LYEHvuxZtEvmBsCbAKhs+lyq8v5ibArbdE10PT3sEEgwz74Uuog50Qioa
OaJmPrNkdL5+X0sNf2ZZo+DgX2TzrwRnmKrOzbVam85QF9suSsmhSQgRShomVhUt
inE2GoebQ15PUyFqWVx5vFYF84O9Kq/nNu6AXLNQSytygReQKtdxHU32Cw2Vnkyv
0CbIoVeU3uQDdlKbs5wrtNq5D5Y6Gdl/QT35Yf5rabwYJobgZF9r+IPjldKfNuxz
xndhJTBWpkyoV/ZCpL9Scw0AjO+ZRxLgBqPzRxAfcgWoH5Iw4o1xomCX2eMzgyFq
46R/z2tsuklZwhr55Uj6f9kscnARXHMrvAG/tpyneTf9Mo9YsLeWKf7gRajLhioC
RnlU+Ab5+++MKR5FFF2Gj428+lGJn8uNxTS3LUI0irOQisNDFdeCoCdoq+SBvfRN
pwGNX8jEKG7aAbho7xTEdM+qqXJg0yFV7WSrvv/xWT2Mh3nFuqMJBTKvD19gZXh6
UYK1UaeojdzzvIBOaj/ifskNp0/o//j5mxVBsXgSnYITiR7LV88RWmbRJH2glnem
T9BjDlwjI2axZgjokjtrQsK9IsALDi23IkZEes9TiqheWaWWjkIF0F2gXari0Xn9
9wC4SIudeDhUFYDcvQpG1YALZdll4wfXcI8UcXg326KdrDczhTKDvLIXmDHi8Pqc
Qr3a1boqKUmT4UZ2kDpW9qDgXLrDm14cRGfSRjugeqLV9n8qdUO0VwAivZ/qv6+8
VEf/u/hyzFnC1Sq8Xw2AaN19+guyht6JC81C3mGBOCl15FN9ZaaHBXMsU3Pexaes
q/wLB2SJ1nFrHd5pF5ctV0cZY8YAFPHy5n2YACuvJvkRU5oMenTj4bXNLo5VUCey
qrg3jBXXccBstcixxRbhTRfgmqkm3zWmX6Uo3gqJe1N9ZiFcRdx+fgHV9Ki8szN3
cnmE1mPTmTG6QSkr9fMTppnrPW39YVscokPgy+ptaStKcuLXJHvAJwfL0a1A5iX+
s4yNMR4FI8+DC8BooElV8PibTvFf7gURMHRHpO/ueH704tMUzWMZ6S9FCTGwZCdJ
3jC4mwh0xmgpsBw2/KEOE12YKYNXHSD3PxBbMn5JpQ+6i3lqhiw3alwCguHwyCQ7
Bg58IZQfBHr7LpwW0WGJkmI+zCaTMpKXBz2RWQZyOlzjGgQtUxrdC26aylLtytMQ
zW/KDf2aHA9XOFPwVcJZkaWwfKzk9y4iUVz7fxzBYwygzT3aBGL7ylih8rEt98fT
5Z7bSj38vXMbmTl/3fKw7T5CRX0rPRYHOWqirfDehvFIq8KL9Y+4JGljGu4SRx2s
NYPlTg3YFcwAu+yP4Oj8dNv6Z/5b2jpeGZi0ucssriY9Nbq+LQOFzojaJphEhyzj
O9OOnSWHET2lM1Z5RvNkq9DdY8YQr+ruB3uRqyxkMKYDrvyyMBHIEVdBIteNOfFk
72ka3adxMM5xAg1Is2moGJeoNg1D7gcADPKXpFLVCSF2SQIys0L9T0Bd/wlbMW2w
1l1h+SeBzIlcSm9jrScUUf99VsvjEv3My6P6G0AzbGKe5IREoDcoZvnryldczSrl
zfDczSebtDDOtPHT/fHXaXasgdN2W28XuyGvpDn1612yFnpaDpKcnZrTV+qQcN/J
/+/1c7mb4inLdEDMY3ss6ywJ6yOyM+3TNgSni8MTNTx5mI9Se94k1Geo4bZ2Z1p4
f1aJvO6enEyVtdgUlhWklNvO08CJ20/5WUcUqmNje2h/yNu36r0olqasFGMDAWdD
dtdTKfg2xyO1GG3Il0t2qKLT9/9GJSeVSb1aFk02EugkQ91Z9eLO5M1Y2mLJdm8g
nuukx1gtbJspjCfBj/6cZQT/sNfUvmBewXikIqmbKFz4yUipPyK+25rSMETnS4GZ
DgM1Ee3dSr0Yk+kYIy4efa88QFS7qcmyRU+uVvvUiyIh+RyarmRLz9l/zuifMXlk
46oVHuLyhuyKHbrsOOn0KwsGB6AkCC2y7cV/3GTg7X8qTKdGlDoXidZu4Vtd1Iz8
6F8CW1e8KixnpjyrptvO4zwEnqArO0C8R3Ex3ZDzyS0aSkqkl2SkojdnR54wEmIR
iA6DhmzNP1R6UkASqARFSK6ejFLx+oaqjGo3yjx7gBtH7aEKP/AAO99UHgyAuV9M
XWpoSlECvQuBTLTUCvnqR+qjANWUlKls9KB7PC62o0wZajJ61vQDdi1ClGaQFbJX
odE4MFPSP4leCxJEu5ypt2O1sePKaTFtL+fR8HokU4ayb8o3GDPcIQRnxZSdOqSE
P/lmot8qOq6MJdF2pMq5tp+vTxLDSzzfSBOV6OTTeIS4Ub1hJwGUXKo1cjOwqHWr
XvPo7PRNvBc0hPWycMJb4KmgQGPcul5f5SOR5ZbX/LwxeXkrg/Aga4fy2XTdw7k9
bViuywe0+MBNJoEM9wHsnUOuppbpy67NWFC31fZ7lHA9eOt4Bu+TKZGjQmFdPPmx
3byR9blmO2yISADtxNEN5vYMvgzCqnyJWxgH7RM+HdVkVFO0q6wjku3LnpfvZnzi
XC6yCgKmKgrqWFzvKw1EQCI17B8jJwT9cGOwx4x2swltcmKLgf0PhtZkXnwDoxdp
UD3/wSzBY3d1+qvnGPfzcJ4LmFezOEOpiHU1UpwfuJjcYhor/+FyEB1SAXXexzfT
w80OWeCa33WOn68aD373RqSqgwgL7HR/JTQlgq2x+XHjyf3OUoVheVlSuFp+g9xR
41vPBHr90JU69IN3PXwWTUcQet8xAHEHBeKSAC2u+4yXY+CWabxxCzu2cOZW/NKm
dE2rHfTigI9yLtPyln/qOSjqqvg4HxaKwpyv6D8hypIMv44TIdJojxHZ5erVcky8
d+Fy1WNOCsjSKicpb/LgDgxsAJEn+JsDlXavWDvjdPw+qUDpceSiolUKyrRt4AFv
0yT6ekBHmmRSXRkvqKSdIfC0zWj1exhj58QQTIHC3TMu9taonZUndG7TACArGdDd
M6yOBzuoQbiGEdDg5DAOYhpmRIdEJ4ybAz3CIZPA2sYcavt2MHCRjLg9354zmLSc
IFJn2d3Nc6w3vsmX1E01gepB2lr0Wbgydct+D/wpGhRZcmH2kKTFucYh9rRNl59r
IoTTwXJ9pddwKrDJiJy7+nTSFyD9Kq1xBz75qD6NTMsvLb3rMb8NZIJ00WopcH2y
SVkJUfppDX1t9pPdtw3aCjDOkyWUb2HzO7KZyqq02fxijWun/VPLTQBcfOS3/zff
LeR8ZmQv6GaMN593+M8lJUu8pzHU1pnhnsdtq0jH+XMKuRTZS1ZYvKQd36wb/KeQ
NDnWtgNdXHsRYeAWUGPZuC3Y7cabRi0cfq432JT51fc0gmRs0oI+eszvmC78PIQS
B+SDy8JbZQAiPZe2SGDTfh/iuee0ZS41/GiKr+vrbxadY++e9msBP++/eV1B5MKw
EwsnpA8SWLQ4RRwpIEGB89DkG0QLQJTiGb9kOfpbVsp4lYTtpZo6uiRg1sPIqAwz
SzSkgzbBYzbNrbWBwmA+DJebJbtQTXR8pyumKIAxaV8tlDMyayJm9hQy/8i9goat
55UJ74nMqrl2tsd3/bHwehhQJdWDbSyG6hj7sAA4d2qm6GK4qMV2mMVQBClrSiPl
UDguvEzsslytpxxx7YoPaJzjrAz6EyAUrY/C1NHnFU7bP50LfiKDyz7g1W08QLRB
j3poL7nU3ngXrATm3tTur/E0xRu48VoohwxwWDS+WYIdWZyWkROd4gpoCmIlfRih
GTvD8an8XoVrz3pgwP+vBbL8tSTEdaVFoGzum8S3kDCbUDJeHLGHFnT+OTolhzW6
iuPtkQWMQE9qeFWF0gemXjxLGYtEwmWCsjpyeIpd5o+4+xrtvgQsk8JUCAFQm1I4
CWIEidIz7/18mnLmm4uibMMQhPoYLiiafkgOwJYjV0A+2YG1qtq0M33pnSFDPOjP
rsMGtpQI6Do23KRn/fu1xPwYgXAr2YJpuGgf4c6Q8XzW2ihnKZ5iLQoEl6n7r4He
6I93FNURuC/VLzlvKncCqLlvir6pfNEBhSTAHhb1Ek8mR5ZQdUuv34MCF76XC1Nr
NfnrM0EPs5Iw85si7yijlYCfJbohQFRNtc8vGO4ue0oOpPn51+1gOYTtyw4A1wr3
t3yrizusKcXhHmRryFw6PznofWBpEx2U20lPvGWpKx9RMZDhfG2+2lu8Nmezv9uU
Nk68ETGS+6mzTBw8RgqVPr3hu1nJgVaupCH1GkBBZIervlGXVdma5QU39br2Owe4
nTIBn8JROgMCqnhVZn9ZkVzfkfIxeR1mk5ZZ5ztTB+IJ8rdArrgVSHe+d2PB+vOV
25TVfGmCfn6ThtqRESJNseK4oPTr0EbBwN8Q/QY+f/iGtdKxgvUwd+xvOXyHFWBp
dKOqKJGbiJSqCbfLGv+1jq1+leQLIjZXJtEaAw3eUeGwfAp+ZNXTpoTyMa26ZR2L
5/8xIgII7l9QdfcaakdkANxtyJX17aZi4JTnw4RrMlwybKc3dbUF30rHLEwwIHQ8
2GuuhRMg27h0Xu+XcYcXK7KiVP9F25s08T//oXcKIvBgGWE9VtyVulrbgEeCS/SC
ow2WoeF11P92/2ccmCO+52nJzYTJymZzfuGZ58HQkOwQWydrHnpLgNHXIPIZCgzd
JcutLNk2nvUYBnZz+d45XJoN745O9kFGRBV3FctdH+gS10XZM8FWV2h7xF6b9kDY
pM1u5pzwoiQiKIc9lO4tGH0ncAGKdh6Bkb5rkIRV78T42MeipMn32ShKXEyNt1d7
Uzxwi/zfRxSHMxgdUgIskXPuCejoDWIJgyZRzvpijvYTupzCq9WZREy6wg0obo5w
dTqF95JVay3zh48p/PpzEVI/EOamoAtP1mMgXNtkZZ5mKzc2/Ki3bgT4ki6LICie
dogC1rtY0njImVJwWi8UANzeFzAeti9cfV/gqdN/hxnQdny21ScL6gKlCTBAaJnW
wkVADvpByKGQIwYfIKJ3sx35li1ZmN59N4tTWRIXL6ZinKU+/yNbH7mWXWGsMmbL
JvVXYW+htkia9QTW4l9pj7wiDcVgW+rXaATyHZG3niwp2DAfPQyqWOcQcrBAc9QK
F25iow42of6OXTiQFKTZz3rfco6DYae4NMBIit4GSLlma+K5Wnj7vU/p4uZq+WD4
Ecmb3YOIc4dYMTFly1seNion4eRMZ0/Y+Q4YS0qKOVjDGPBH50FS1zu3b3ET1KE6
lJoGnkXLpV1dj/jsIysc+TA+41wXKmlmQr8QcegFXZ0lwMv3YT4+ZVVlxknl3Yem
Hy/jtvG9vVYmdbbv9/jDofIR2AgJDd8ZiAL9H4BvW9UOoutI/b6w076IaaDSxKBa
pk9nWADlspZ34yP1TV6tpH5/J6gn8pS4njboKx7QetAaVVeulzNRdWngEizJcSQB
+9CRGJ3xEzLM7NPJo4edZMl/q3nKEkhPGijyPB8otCXBFZVaHMcoZaQOJsc3n060
dgXMi35EgtCvmx+dpKFbJjY2AMGiX60EQx1kwDK9n+hySmGI0x41IUC+PK7H9kFF
b6oI5wWV7O0THZh+CZIEQWvsLwS1i8kIeIkJ/81WElb0/euxb+W9H75ZrbObzWMv
gwso2uF7o4hdVmUFdgs1lj+HQM06tzJ57mPeJtbaMbBC1rGb3JodMukmNatl77DA
cScuqh9l7U+2zdf/DkdzH+MvCqSEAhRbTRJxCSlrvo/tPi22e4gP25TxLLUOvLWQ
mjy1zYN4W/h8CPQoFiL5ijuKJvyyWeyNiU3LElG7GZ0kR8BpfVVSyO6XhQHIsH5w
mF3QNo/8qaVzez1QnXKo1lIKO4ryLgVqy+mSRUP9ijfUUpJl05ozFMQmXJlxuItL
ofKrQDVkQyN4UpCkIZV0OoSSuEdvR9shrtBRwVH/dWWtU7agaO83hSwBr3v49pRd
rdQ4NKGeKf07F7WYoVYi/9KClTPQo2JqYF4zXT9vQuePBYRJlOsO3i1COzQCmb37
cBCNuc9Y1RvQauC8sVeYy/5Up1cOjTagkbBiWmrFofkJcAq4h48+tlAyVDOYPl8A
6dHqgBBnn3PF1u83waERV+Io37FWwxuIkqoSvyV+brkdEQd23Sdv4wSEqMDfCbXD
y+aDcoOMtiWBEnX0jjj9zH+KhfmQMwkWtg24XYFAzLoWrooghhioQdmJ3wc/b6KK
VpVtI2db/2hwdnd84BEYpOoKbXddFCHUovxcSFhjxK0BrsQNqBfPxLv+k3cI9vMV
cE8cqcojPvruExJmXlOkenWktE1AuQzjwd1jjkx4gz8kdlc0yERnMNndDHkUuvM/
Z1Wa09i4M5d+ae9KlIzRrhJxk7s3BEBQXswUWAROc7iog5Z7yKai0WktYxFpEVBL
1taoTuR4jQdldFfqCqRYoGoQyWGinR440SpIFVMUh2yw3j24M6h9NZF/Meberc1+
lPiS0bfiqAQjqD0l/g75f59RH/TF1v7O3uLsYJABk7bN1L4nRWK4FRgnvdv4EIby
JLZaJH47L9xIUa0jX7vNFF6nqGt2i9XFqeh3/dJuqkjk+i2a2Aig+Zc/7bYnY/le
r0rHqt91kR0XFHGQy9CS2YwCv92vXbwJVw8xQiyOhG7oo7f8g+xtxMo4U7bnPMD0
y523+Mj/B5LWh1+LkTXDLCeccvL9WFzI9O2/CCZ+Ngxx825yzDkUfjPYLcbtsjlw
RQQaIuKgWzFBmZiwWcbOflgzLxZPMYl65BNm4hR1z8b1lL4qGHPTiKHB9V7k8Eif
ZMpMEFzbeF1l2aJQ62ITpc6rHU50K0wSn3wUpXtJUnKaYUC5C7/PtreyWLubMM82
Fi5+rw8g7JZgGkFA5Jv7Vbgjqb5I0iQ0XLglrE4X8mcs9kCVA6sSKZbu7g8S8XGl
O5ZJ3bv8cpNCgYFME5Wdi0tEqkO1lwdRyuXRnvPK3gIIaxR46b5yJ+/7ZVxk/2z1
dy8/+/3E28AFuJ6aSNzyWoFE+eaUJXSDSja46Us/0oLXvG2uutpENy8oOcWqSQ2H
DyUNu5ZtbKQZPblH2MhV5ZUH1oomo86vEJHifYai9vpjkXBz0hDm3HZNjf+o7tsx
1k4eYhZ0JLcEgDAOY4it3uYWXVZiq9oe0BJOFloqdJkXPflMEx5nfltVhhv45YC6
RrLWbD20ROQ6zr2Hkz+ItxtS+qYJQ/eLzNlG1zQ1NH5rnu7y+1wLcMvgcKBBAmCA
/KR/LPxUCzc9i5alUdP222Ymdr4kHtggIm44Bod9JAMLOJjw16nGVzCmN8lvSnAR
EeUOPFQpsJnGYcHDp9xYqxyzHjU+UO/FrGayKnBvMKosc/6k7SenLfeefmZD814+
COPSmchLFDXYGjd+lZ4LLSQWGupyiPDKhKyyXJ77sgk1nGQWTxQIv+ja+Tp3Ce7W
AmcHG77UqTzBDZPU4veSv4lGRq2D47LGMjAKiDhvYyt6UwOKXPbhLhX09za2el5P
tEmBYoCDW0caLcYuHjAf6zz0jpqVDD+EI0sld0k+lkT+moLn5f3Bdy723IrpCru+
FQg/sO02P4NKSitSQiEQdLzVXuBkstU2mLgkWpBVQprRXVTWXYsxq+qj1BLeZbTu
+zYiFDAmXOUQ0QAO0VxDBBqwrIb6u+RSnIvjcWyzyaoV8TiGntV0MtQxuqoQ4LK2
Jjj7jLKbyCw31UiAooT1DNQ02Zd8mHxw11SbHmv7aKMiKJhAnNwI6mz+kVjvmyUD
6TGaYDFKJnTgTMkVYRChvSgRbJcDOuxxe00/HrlR3Gb/h2FgEssc7ipBjd8KwquT
i53LxsN2g4S20TSAlCXJYlJctRaLnMTTbmE17e0ALjdBF9KCPB59dxF6Qywh0Kco
hQESZa63VEGI8xuJAGaKdi9vgGm3GAvu5WCZiNcY2MVl6WofjmdwJAqvYoEXEBmT
hvEQ5yQ8pIqws0DhHlAimSlN6TEWliXirb17NsUiDjriZjqTgku7K1m0xlIc/v8J
RdX2FWsT0FfdKBODU8gzUjJWzryRZ2JcqP9fiUL/esvhed1CpFyyG2I8BCNKPlv9
bLupJ5GYrV7Ixr5yv9J81LQnT6mXyUwQzu12NWmlD93Vmzpdlqbi4/l7uj7dw1/d
QexGtNJHL0QU07Gbf9NNj+gvqWaKKSUd+lBvkwgt6GEUAaTi4H2jBbUDDaaDbCT6
KBOXm0ZAvyYJN1ouOVMTujmZ03o2U/LChpyx36srE8LEeNSh6gmuR9r6q56wA6Io
qOWtmawZe0HJy7tMpH38hyqV8n591sxSt3B7B8NQ6H2KXBEUE/IX3ywLPmEvWfKp
ihRY80CFeDCobQ070/i9LqVbhLYlDX9TTWgZTh7KFhOm5rTtnb7vp0OlQP9nQ/1K
/cL8OpLFu8+HGBMsbWMU+W3melAjc+MIpFrpEMp2vQns7pM6VMaEcMpLt9H2ZAMq
QZL1vz1uk97Gg2Smvvy3YkzRFboi04ErT9O2Ienz8kwfPfAICunsPD8EOnZEPAlu
bHgM9JaVSyNK8f0AT23fEuzSNnIQPY3Bhw3jfDb8gWEMzS4IDD+Z0kWCaoDWp3ai
t4O7oJivHVR7oFAYGYj2gpCOh6ELrpayDu0gmnjyosRmt8rziYbsDrPt8/o15d9w
7tMGrv1uyQ9ELbbJQhn/2NIy0H7K/ofUymidpucR0s8YYm0uvSxMjvli1VY57/fM
RtX6cbd62QD3TMlIFX1DJU776v13k/KMrJqvWE9khb17QBtW1v6KDHnrbMjGknk0
6l19bIBgsWUK9lYMJFBzid85Oa6EtyFLMqQ3L7FqIz/Ym0jGuBZKDgGeYxqtmioM
JrxFFj6Hcsdzxak/8x7akCVXeabQLIj8BH2u5QxVd1jfVLQgMKrP/Qk7DFJFUjXT
>>>>>>> 426889eb8ce467b9c9a9f74dd4af433c5046285c:deps/flexrio_deps/LinkStorageRamXilinx.vhd
`protect end_protected