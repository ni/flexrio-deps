`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14192 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
hRRAlfE1xLfeNfywbrz10PzJRff511XkZKpyIOZYaUWppSFfb85UVsa7AzF1qcyE
lhDv5Jar9pFjQ7xZSk9PKCYJuc9JZYdXz6rm68s3U8zVhtNPSma+9gp2rRvofIeF
KU4tJ2KGrz7d6DIdwBg5UDRPgvMKrJytIrDGGXTuvdtk8B0NxaPTtdHdyK5Yam1O
aWthZrMW+7TGcMrXfbwVxMg67+kDHA/79s5XuIbEtqykbIUKom03R9C4HcRoWg2d
152ktd63+F2EMXUgY+VwcI/Yzky8L99x5gjj3Ij5AilXdthgf5KAmxRpLYOCqHag
OOU7TeU5WMJ/PPqXkUOCfDmK+lOFUNWCBda19ERk9hUCWX2zHewUqWVJsN17d7c4
JLBZSz/dzvKo94GH75SFDoX4N9HnbO7J4M7L3cYPZffdB0896/aTBXvH1t5PDpxf
xoa9TgqnuXsXKbulNtJdv/NOu1r5+mIytEf7psfRYpUvd4wC+0JiyRenE8dn+4uP
Epd0Q5SoFFF/LbRwgulduJ2c/Rpe1/GQ9/gkEXGZ6vD/G7lkcyzyXz9PLn3rYvoD
ByaceDKC4N0zTvzi0b63OhYuwGtvMtgLgG0CAeTPiiIQUQ1bAEW0pjlnraM6/VvP
WY+H3C1yLioNVx8ppGwrKUb9zYu7GpEF1wjQvRgH2pmUkXLQ8c294fyDNUVZ8cgw
TV71rILThSY1aOA8uJiThIAZh/qrUYB+nrqRSgPjhoPOIASSYU4dlcxefW/QpunW
3voGnc3N2AoovBKhBhJh+/y/NctQfKB595COxLXtFhKleTs1JwdslwMccuR19GvL
gaOs2NHSaQfG+9sgAt/nLCq9qfBNiMij5h2y1D4eF4uTF34Fphv1OisoJt9APuV4
Hg2cMVDCoPGsCdXTj9k7zeUgSMfY7+b3Ud/oydlMCFGDq64ZRBpLjp5QsvF3dv6+
JaXpjfORhWGESykanIkkpx+yr3j7cZ36a32mMELrLDuc1BWKn3HjgT4w2ntk3R/w
Gc76wBaBy3BsjSlpSX8xdZhNiH5gAyU15aCfn5mJLJNUMWVatxOTpu1/q7yMCc/w
Ox1G9cHdjOG8Wf7M9/EXk3SE5BvxzjRdSpylUdY2VQA3bXYbgOWdaR+asLoF4/RH
Q8guRA68qAiQkCBBo0cZgTtX5boDAFZFx1dJy/HJ7WhAHczlCPXqd9fMq8tLNOx9
lBLhDjb+7ChACpFdoRoJ44fn4LDDNjiKIxVvZbwHvr5Z+AVl7iIBBK2Yd3ygIss5
SdEdOV+R0CFz1FmZgMVSPwbBcuBUa4R+jh04XVG1sMLIoUV71uK0j58LLeJfGwvl
xjlDWWiDPBvkpP5+l4VjDxlQQ9/POfZCq13Be5l9f6114ZytHEERPst9KyyZ89ip
bgKLqmxylWXqTOvPNAanYyFOgLDW8gxMu5/VgyTbPVYlrqQMXzmOEGfNcItiezyl
1BtcNbRZd7SCCJRgeO1iXKFKX8I2b/zo9Zv0lR3SodSzWH5+e4YGpDumrWVM9qzE
fYwUvA5a0QuC07nzPe6MVKMC83JY5Iotvjz+ZMOT/+OlPGaUbmJ3OCJrS/w0uBlo
8PbH+P5PPHGLrMhzY/YNh0pS4Xm3jz5aKqQhx9QFHDBfAcsUwuroIcZLXS7R2G4J
uJZ/19FjLOND9DiLRO8+ROKl+5OAEClujm2Pr/AQ64HjLEsiIWEgfnlQyVe1WL2I
O0W/U/VZU/v2rHXgcfqbHE6UjK2tTYIhF6tPZd+GXWDCYecb2tIffTnu3evYtD+y
UdmFmgigU5LDQ0SSgitlu/pa60S/gFIv0Nr6RMUwd/YCSQDMXKmv7/Vew8ZqQQRs
4WkxQkTJxibPdQrgRtzYw84bLdNaWPrNVpwJ9Eful8iTYhE6NT7NZ0lwM+gHvH03
rLjqPzi6DVWrG7NOnVT4olVNntYgo/h5tLbbvZ5nOZ/UCGOGMuISnPXpPxQ/pnO1
roBQBt2Wjqp68XAbWZk36TlSv7lRGBmWuwnjG0DnawyXDELUmgVGa5bD+jdIMTts
LZI8bUnlBTAcvtz4zncDFwJnOH3GmFDOldtyhTEqDcAho2nvKfTfyvKzMDRzDw7t
ezZf4HyCvBE02daDuex6sDqXTA4SAe5jO+ZShb4uLAqezrOQMvDrPrXsdZW75V0+
3Xt30uUoawqmOTOF/1N29WIUVILkeGkR2Ql/PHjhoA/GNGAUoDtsjRdrqzRrFPh9
qExrjJgbWam+4o59wcKV7B/6ps67MwBck85xI3JbrepToogp2C37H9RG27HFpmvR
d9jd9U/pOe9W75soyuTgTgESLxAIeWbsxllMFa9oO8+EYGS7jZ8Y4t1LbyL18G8j
GHgipBZCCiAveoljIESsLWzpAWYXrn0Sdl/yCwVGz5JXZkwSNEgYeXf9OOruMjZw
y9iJazeLmV1giigwQ1jK7GxIGAMgVAOaJ0bVYmFqXIKBnUBOU003xbBCHUec9PL4
OgLA8YXZzvufgfeo4L9SPMLZlwe6WYcbF8KIMbhcfQ7Wle4ZZYXpLYlB3TvFN/s/
zWpNnoN5psHyuPY55ljzDOBs9TvGcmzCPSBC96zrzx9Otb9IJU1ZVM76AhsKyjDG
RGfzOJGwoq/U3NYfe1TZYpmvDTyFqfd1rNqxSA3ExABIcjjA6JVNtkvWqZcmauD6
VUgR2gGO4Q6feE+DH3QFziwzT7ZO3NjdA/XoMoAXImhdYcNC3ykItfuyIiDyy7tj
1VrIJ0HXbyVK6Eai3P2aht59xU8CG75fp10iD3bUp64D1m+QRhdrYaw0NA2suGT/
YP/kIAzvtEA1Eh8+rEaoYY/V20QE7AgSrbKdz3sJWL19/f6ZicmCwYd3EhSHP1RK
u+Rzxeeb3AqQGAWNOrAZCIR2tPI+MBaeccCvhR2vCR+T3L1Z7TvskC+0qyz8OYV1
eko6R5pCANE2pdWHAql2r7Si0eErecBotJMUWyPZYNuXEjPMllEAoL5RmmwFeFez
Y608pniwK3HQ5CxaCm8N4aSdYAoj/fqt7ymYAcmrHWnty1qLcTUA50M/YgOTNo8P
VC6KI2PRJCDSMxgXbXbBBY1m3y7kDLrShmwHKSAvl+s6gzUIDkZ0YnSmgNBtKIFi
H3V0iyl5HsWrWtQTRyb4MgFo+RuRUxuQMx/5TJYmdBkFWWHYdn2bnIqWJVcZxe1F
aXiwzR5LBUu0qSFoQldTfw5zKtV2fU9as6GpQQQJDSi886txv/QuyjVh8RZM6vNN
N8uDff2COZ+TjoFytDYijcXStCI118xNqxpIZluxAGQ7LkK0fMNhpHPwqf9/94kJ
4taLpNH7tHIzrFMVscCN/GiPevx//PpwmZpl5nBec1FOMSBQDqFohELtx7KfuDKD
sOUiEf5lM8FuD4/bInVkt/pUepUfY7oxtqQSk+8sZtsu22gfNi53ToBnb50M9vwD
yViC/1LOlZI3ojH0Al0qfvykrfvAyBrGRDmRQcj4XmCzSiNot2wo/XBxAI+Meu9e
8u0pWfnw4XJFSza2r7b7oAHBX/UDKlTOoEHijzqUrF9qAUC3seitYyyKBM2Cap08
I5rSdGH5XS1XSIm3LNXABTTiJKYTsyAt5Un7C7x4JU3x2xdT6wHWWYl8tQnt0VcI
cStRhqEq4iWfaqbVMsuauzV8YQaNe7bKRLwvENysWdsviAUu2BploCbSdhy9GkX9
fnKrm4QPIVVw501pZQn2LM7xSnRWYwxqoRPjMFQtzRDEcYy3A+kTMl287fsKza+4
SBo1ibRAj53CbnGyGBhwCP7O1kmcnBOHHMVRxYxuyNfb6IJaImE9pYZDv2fwS8Wp
51gqJjTb86cZcYfr6LZzgn+vPb00RoJEQh63RSNVHynIXb34RdktYDUoBmfXP1ok
o96Cfc4VE0+Vddy2t+CkeaOrRSSncu61I8KRhtC+bafThm7lkcfUaPom1B+1ikgE
ATlERn4moHjpvQBg+SGwyT19ynQpK7MwUnJf4TnKx2C1qSatPiP3W/PiuevQ5aQP
9QTiZ8DgtXmPcv6+QTXzPxKHhHMIFwl1NTYQnqlaUUaF5lx/0HJF5jCY8oz/Ysbn
8lUlRQQAk9N1wHFGB17+NGbesJhj/6zsOJInpudOk6NOegRVSHLB9Eb35I6T9dwY
xSahDHstgvaJYJvIeS8+GHeN38RcKpkwEDAravRZm8GagvuLVIP8nLriJ+V/a/2/
hGntViwytnSA4HOrlW1lEuiymynzk+E8v4CzkYZ9+1sOhYQAqeZsDWeej+HtZ3/8
tzoTVTrbtuLXDP1frQiBGAPZEe3Sij6uN2atc5FnQJ59ZA2WNjXnIz5DZ98Hfxkk
Hng2AWg9uXwtoS/wwmFruirw71cnfPuDJdbYxr6SvFa26lwxW/GZOufCdv86WsNr
+RQnX6+j6q/5UO6GH90+hfquZvaeZdEcZpsqMdl+HqG+Xd6r+N0qacqLvFAxM8ib
4MGjiHkXL7syiOCWijnf6TB4Sw6cwfyEhs59Q2IrlTNJz//vZV4593i7EpMRomln
/vg5zF8XZ6GkX4mu01eNuEIZgzceqp6/KvTCZ3Kyrn7pP/Lx6iQt482U7C0YgCVq
GLPATVBU6wOtf27Zf4Ty7IAWv5GisPhKTed1VrvO6d18xdAJu9rL8SUitfL8vIH2
/sDyV7LtSiBpRO4STWDKfU1zvDxIe6UEXyUSSwvOrgxevCYU43tH9yfC6/naIeUc
OjUlV2s1sAgoxuiFWlNBxvY+XKI/zgPFLA8pyYwkxfzWQfPQdmVQ48WFiAhUA5SQ
aDYK4DZtq6pk6iFPuKgk0DX/0Gt+Q2br/bGowXyQf0Rlu+04umzqZjN9ETiYATlR
c+4Wzri7arAnuMwZPcNn5yX5bSZOF2RhzPRPvp5MJkYRdGVP9V+2E3vwCJzl0Fi3
e82MOj3xfZhDYAIjWykMpmfeysDhIJHzJvAP2PbyxAaPk53YzcZnorv8M8Kj4pKi
4rCzDyTOPW+JbbqPF4Ep6smqkG4kVdUddb1Dp8j/TuylAxbFToHMggFLuEAGFYak
tP+vPuuIRV4CE0mUlUHc42g6QKNuZiKSttC/CGJRq3YQjKJX1WT2S1aBSG+y8Ve0
TETtOnFHQTD6VDhJnyqOTEprdb9E304/IKSHFlv17KRL2l8qPBPx6tO9Zik/5NWo
RY/y/keax3ZskW4KUvRe/ZyAqaPYCkt2nIW7aswz764VJAZBct1i7Jf1m01H/BIg
BBEkIYlALrGjh8PVVJFS/zmjvyfzrVztuu1MmiK7JmP+685u8LNA+ERkxzqltaWh
XhIgREr5a5+gXvY4RjcnXMV5PQH1s91twvjquTT3xKuD6jKIP04+M3DbpGWQ169Z
nwY6pEIVLzRiYQsZ1PVtur4FxDZq4EQ4/AptJpHmlb9GagxPAS7dX6Bdqlc7cXSG
1jeaYw2zUDjVyBTFQ0sS86NByhtKWiGS0GdjHS8HD8SpSJ/s7zm+7mkvQ+yTOT+Z
fyFIDr0emV5ZzQ3iZtFwxuvW6L14cgef9b7Eq1tJ4La+vEeEFHqALUXUJ9MGHEVm
V2kqCyZdXvIKs4LyHk9za4zxx6mrVPfYzJDfprZpxj3jfPYJdJsKcCpzPCJx/ALg
oz7tP+rj1ajf2S+uGnAwUdyPcYgfRhOJodXFvrdnt828jISZqaQbAij+IuFZBZTB
pMS8WHYjP18CXWHexAz3oJXhrR8MV5aK7/FYHMnou4RzJxbLZajP8OOvxxA0nvWH
r+HxoriMS6l5XDWauP4sNd8XtnVgtIwzTJnvGwDXwgeawR5fun/YdHlNNgo03IyH
IgS8pRCb6kQFEAfzK4QLYAADuTgt1Qxazf97/lA7TyQQIdfKqQjoRchKOl4GTNeE
WkLNkGRfIG8TX4ZQ/iUmjtYRtZHI+9gs/5plkrUkDYyEcFbRT5GcO7vULYZpUEhQ
EUtjHXox/OBNzbsdlOAYYOsaVzeYf4CjPCLlX8BGKmUUioEMdYb28VRlMqud+1qV
qe0LjdW7+kZ18d3JWRhNNe3iZDBoX47Es0rio++3y1b6BS+G0D9QMv8WwhJG5Z+/
ZxmCUZRCPPPG+Z0eBSAc7yk5OC7XlimYRo82ik7MM4KWmfZhlhaHSsag6H/VtoJ4
xoNE3/rDxI9x1wI6A+pxC9eGU4/gNSLO9uk66Am0n9BAEispXbI9LBcQ1Pd8gAWV
XWYBBdmkL4YirY2FR/vs+VyBYktwoI6fgRtD4nwYP1Iumox4aT8pHL6XnK6U7HRB
LtxRZiwISQ0x1odvmYQnW/y+3R70yC2DDmtKcK5oTSe82tjOF0s/NCbES+FSyYRA
/8quMhNHsHYH7oNlE1MERhej/CNHmS1xNBgasa1Hb+lp/93zSAUdnEYQh2NBOx60
ZgYLOBXMPF4qQVSLfi2DOvhOmMcsD3de9xIkJIzDVytWXnZAq2uGPG/rM/WxYaYf
YRZPqfk7NEDcQ4tA2kH6aNjQLs5QzJx9EaV8FyC9XAGGLygew0wIhRzcx0oMkwP4
uPTg0PaOuUcgmHEGUzKte47StAgBLxNRSwytCsjN7i9p+ON+ijq4U5LlCpoja809
0hvor77RF0TlC62n3tgn0yTc4PtQOGoP60+p84bnkaDCZTBJZJ93w+aqmOGt0isD
cyYKlHyO3ZEc1CuWj2a2RrVVRqcqqvsXRvjWZktujafUV1sgl6nDRF8RInzYM2Yu
AMbu4v+nlExBkW9zVCtWypcdcBpyPnqTk30Xcd9MRFq3MuGxmbk9fLG4GJ3efV/f
37xu9Ie1TzCIf/TZxRQ1XI47XWyPVJQXG6zA7Ii7jXuOfK3c5by47zSp1/gCdtFr
QjDUzM7cyNKvcp+5TrsJEQNzMqwtHxZBWITA99VXMlgJfHr13JkXDSaP9bTw0Qac
uThXl4DVCwOuu+P2rqrh7nWBMCQm+7SypN7fvsceckfqzxJklmmu/Eqa8PcWtesT
53ZG76jbzZKAfNxHg9+M0QLHPdRSvIjwmsoLEs/GvZJ58oshs4puOtW4iO8xpBrl
18WFrdH9cjdRBiLTtyN57i7UHHniT4D3qNrbKvD9jA3bXXkmFeGG8Jiamc6H1waf
RUSaIUf2lJ6BZqD8SBHJIMnmUtiKas5g1ONtqjCcGnFcsaD4buX+oT5NTlO6/tvP
3MnrnJn09OeiMQtxUzVEg8SZIEwTDvm+hz9g6cIK4JNQK5OeEJdGXFSWb8ZPbmpK
dbMWUtQkva2FcpxtSo88t263i7ZgR3nIDD2u1DeBXopC9NcqQwM9dLLzA7USdRw0
an2uiw0vQYMA+FPPMuGZxlgT4F29xztRIWqbCBAk7XmbafNYl7ITj9s1Ya7hXXCt
G/vVLp52h4SHKjv2WYuUwzASofHM0wJf03jLtNpDmEalKK3FEkJoR0mLY3hBM3dO
E8xnVva0lUUkEQyg5PCb8kr/twrApoECYrVrzSjlo6Unaj7ujgEhR7sijs7INR/n
X6uvL11UEb57jPp9n8zvBPtExndH+yv65eyAmUeLWfjfDppdZO16XEMGVmrAoxo8
Qxcow/hlMq0loqH4/710PBBYEF9wMPl3k4Htv/dCIuBz923fIlsNg/wYGUK7jibe
K6opIMuKTYALDtr8WT3YuyznbSVD5TKcFbek0DJLWwkPoGhL2bTRXTlB1hAYbOzq
WEc/JDFgkdS5UPUcPjjP3lOZfudX9uoRugUoHL06gAch2y6FfOoL9lfyu2mXg0Vb
xkEGobpwsRqrngLSlrCiXOG1T8To6ZnMeP+y5e8fjjYowBYNuNjNm8rpYoLSqeTJ
OnH6NCilVJwLuXHiDhL+73w5gBi9iNT02PnwNL1Fw7IDCPzvLdNL8MKuLpbRk6U/
elRx+BihMGipcx1JzeNELMRKbJtpyzDzisjy6hcCO64/1enG7qE66duQfzCIjxnI
OS73iGJZQJjTN09CEHZVVqNUjxkIbAzUMzTt2ecoA0RfQb4Ux+wKpTvuznMGgxpy
uncD+tA8Dwyrjq0gR8qin4JBxNXIockuShex4xJSb7e/wC8+Pj7EleBDuUdq6S/y
gC5ilYigQt18XbyLxk2Qi9sNZCelWgXYFKpjAeqJGs+ikCxIMw4Ylr8udoyRvj2L
OSJpg2TFHlIXjZ3jbpRrLTvJJegCRw2hX3ZA25di9tkQRFY4Z9c3uzFTPBn4eVNL
JdPdUiEATb5/MjsOTPacFBo2XQgUHqTOT5SK2vdq8HO2FsVepjWU5XcptLRhgP4v
r7G7efvvyyW3sZGMXHSHIAZDyrHMFcQCMAfd0Wr1a6KHny25Pjl3q7YgmJEwMm/M
t9nCa0+3P8ohcQHkCXYhqPIVcSjEqqVS4n1Jk7sK5MfNsPNAj+72XiQU8f0i8bIg
yYakleZUCgJn+nMaKDQWVC8iFoGrCtWnfmhG+y+0Fy8g73Il+78R5XmffwTTgbk2
n656ZQTv3mn2uAcRE9/e6xpmSP3Znl0JBO2o6/Iglhkfh+RRCZq6Vktynskq0itM
Aye1InO+/25DSHDJzKHCFG4SBNeT0tURTAJi6F6W3UmUKrjRSyP4NvYOU9epWPd4
bpuxKf2GWQ4ga2BhkYzunwGT1SEs1l86E8IDjovc9/j4auu6DYgDdsFDXJ8Dp9fo
ksiRK+HQEKBrhYTc62tX8ero3Wfco+q9F1Z6OYdNDZexcQj3nXnuns0jSfDZfms+
ZjZiQWmSaRRjsxtMpnJ55q4MTCdtSgmkxuQVmWcuXndRAqDnNgnYyW12CmXeB11t
D4+YHUDMw//LsxKULcKp+LhKBcMGn15mz+yBFTvm2geCAgIY0FOaT1UPqcUTAc4y
FNpMuAa/s3vBwR2Gvmi/wPmHUywgwKqUAI8mZKKZE8vHg/kIQuHJ5+mYlkFfELIm
+5WqojWSYhkskci1bqwQR7SGKUQhu78MStq/kG/xhPIafFWwlq6kcCiRjSfR+ZEg
jGNjPgC5AU0RkT1DnB/dVUMZZY2CAtNpF1O+ASkYjBI9MjjBGJp1xPAL4ahK8sIg
pnQohAv+XxA4sizwfDKKN6FYLrbuZF7S8TXk9GFY0Udv8AaGi6kRdL+zV8CTVoai
rLqsoLB403U6BbGgCnCOtjiE4OAZ4eV/JrbJbP4mue9TOWQMplg530SYuGHmwKhj
7qObKm1UcIbRDKhoDgmD4z8/fSN9fL0U1AMpasPRH6A3dmASF2vX0K/tf19kGmQH
Rn4RGLSZadqgmGzM/qzD3l4/dKuxTgWRc6LOa8Y7jEQpf1IVQRJPVsD7+O9mmTRd
FTxTI1K+cCNY7SUCPfF7nuiII0wXwZ85gVTwZhiTVV/bZSFXR6Ay2mNVTYYd6AAV
EytvwPF2L3g7lOVJuKje/3xGioqvhD9TWIcpn1rnrLhJK7NH/xGygQX01zClitgA
FD85tkYzb7pit9YbvpSKorWJ6i1Ti2U5PfOHWXmG/EX+I4b6D17CPIWOlA1UNBrY
p1X+HiNbZW7iKSP+8N9AvOd1dsesR+rRj8Pzo8QSoVf7ookeueJ5EhK4aOzpPwEx
+v5jp4z4Maki3HhcUH6jUtm72WlYoKsif68hgFeUGWDVK1Tky17t1P/Leim/H98g
Br3RoqVYSpKB25WaEfZW/evAfILJf+nRnQaa6PEm9tu3fdaIOodi9x3F3Qk7nEat
xIaDqsnMBtFGqP8fAGsamWWxE0y0471SFgXJgsLo+5dEALry2VM5Jec1od+05t1/
8zv29l0Q65jaQZrkLEcroQzVmB2EAJazVij05Ve8YY7wmego6Kz78ChLiRnH+yPo
RVOHEbyMZ0JK6nGMdbEaWDv7Vx5NiRlWAwPQTXE8NOKSV10dpOW/vU6Cxq9PArQw
CBLkDE7jzGYfMlndGBve5EtqeUDKEhjIunHohPQpyrwUrhYbmUkzKlbsTPvMLiij
s31CsqcqbpkS5B0yoGUKT88GlEZ3TrU8E6TkAJ1lSzIl6QIGN2qu9L4pvSid2b28
bGvQTYqqIsyBJjDHRMYn5on2UnhSwC64y0zi98g3cTzrke7pAV/psbsuHxU0fZ1A
5dBMMRJkoeldEPWGWVg2cbLIO9iMB/4LpvB0zeLouUUkrqhxn+bDpfziwwwesmH2
pMrcLfJiuyCIrDg9q6QKLGPbAgNG9Ky3el89S3mqIf43CY4+jtCM7L2KGtoQCZrK
N5zn3GZchKQSnVAC5xGLMVKE83FPF27eJR+aoCGE6WMqxNv+EilhM4EST7LDnRud
ZAu1sDpcVc94/zuQsrRXnUJ3WIbE+P7JUUKXugV9VoEtrDM+BarpjX0CSQR1Gy7T
Qwrq2thQK/jrW5WS1LKJtPItKHckXqwLfeQ5EA5I6MTvfKzDGMprubhkfXTE9XCM
eOpnTL5aNK6vtHjIklGBsY1Js3LKv7AfOfP/sxa0x7e2xJbCy2aO8zlfHxpDnBFf
ghqPg2DHkLJ+M4ZLE+tqzJZ3udgA+iPfgGIEErk9pHWIxl67qYunWjCgjUqJ/bBK
2cYVx6Uvx6NMvCuMN+nBcR8y8KSqvVp53giW66FW9m65tKoUAhmGGQWTdkiR6G7c
H27MEX4a7yIMVzd2tv3eVRvLgJKFJkD0g7oHddMh+p+flZmiGEWDyVVJiSjoyEEO
MF4ZFUG1QP3GQvsdc2r/rt4IQrHE6dzs8Tdarj1cwbsX2OsC/lZz1ZA3qjOHlM2q
T499dBr0HOIrISoNJstyqogn6tblgiNFreUZ8Hno4XK3sjqSQqeeqL7SgwbH4Z7G
WyZAF4QebvnbXRpqefXLhaC+esrR72B6fnM8pUQeqOV5U3KwIksRSrtmsRx5oRZ4
CgdtBvbALfqK64dObHCEjkPVRo89MiY/63O6LcuW+rA8INw8ZrJZ4/cIda/+Y5Q5
Cl43S3ZoM/D9zGI9902IRqlNXg/19vJ7BfdZy0NJNPhG8GfrWz2xnGabiac5+81J
vGYn5SyZmYGE+PcLXtidCUnwy+ZOZfM4RFbvErGg/1rM8NYoIrAYaa0auojnAali
4yQy+XmKaw6FLbaJOHiAobfELYoOzgZici9RglKuTX0dR3MykifkVaT2/j87xnhA
7WEUaMDb4tkVk/IoIzMGf5rvomwtLGK694Xk99l5xR3GlbP31nkIZw73TinKPz3P
CtgiVgWNx2Xqipyxmu8ncxR6mDm9KqKkFwHIprcpvV0YEKO7RueRrQxuH6I7B/eB
2+xIuOOOWpd5bp+LxOnaQ+XnwbhLU9dg0PcNlvUh+nXP/2NMWARywpWZFUA2M5b3
TvJ9Bv7NZ1AKTKePp9oHa8eFUVLUYeCeQTq7Aib6YLeNBSDhKk4em4gYfS5EVpB5
htyupeEVbhm74XDLcxzhK4BKCCitbAxpisWis3KFrwtLdYz6l8toxKW+YyLTiTAU
z3LeZQgo0hWwuQD0VRmN+X3Dk57uCwyEq8srqngjj68FjdBGgj7pIn1LAqTArFIt
RlKx0pkf7bwH3YrfnQ92m9vQYitVNw5gTNPzLUDtEt3Sx5M0jwIQ47PXH/S4NdNq
Up2/hA3Dk12JnDakj/TCXqNcwBSkZP8Ls08zoKuW2yz3y1vzAh0bCP0rrgMbg91/
9B+WF2pluIKT8vTneT+S3LhrLGka+lIeJt6WEeFSXpschJXCv6QdrJ8SD6b83Lme
u4A28fJAd8oT0Sr6tkjZUEXMKKXhdGuvKo2BSSLnufUSmLm6mh5JjAiz6vePpD9d
CEZ1Z+vhA3c00/zMH616zL/N727p+7uslBGPgQLXtWUX3+A1t/QWK+1Bvjgm+s6G
7mJVSRZ5nN6T4fo8MMq50jQxbiv3t+Am9LseYovjSd1oCd4ZTLjcvwbXxEGuGITT
IikPNXEfBdTDrT4OUW6aXK8CdPFfs0hjgLLEUIe1dnqMf7GXt0ZxIhbx+pYuB6L+
LYAbByn/cwSH/YPHP/W9q9F9UzNrxICp+PERtMv29W+8y8sDg3qoQ2q9u+++XcuO
aMY/rqrAdlJb5X6X4Ky7HYXwx99B1J2cJbKBnOEmb2eLBUNl2B0r7QaSaabK1GcY
88k2sof95FCxgZ4tdmJgVX1dxWRe0d4/jGV8HpAzLm2iJcHORZva4pvM0sXix2Th
K/XOYm/uaMkXZTwwsN3TLAonbQgX/N5+9HSMFYxLvgoeizqlbs1Slvh8+ItxZ8ZO
9qt6WpuIXwJKUm/lcedvmJeCNJLVcAKnelSr/tC8kMc0biyqusIdJtWRdEWmUqHo
t+MqjnNsgsTymoCYRMqZ3pcjU031sPh9uiCC2mU5boqyPGVAuTAgmdlI9o/j/qn7
vvS23H9aPp3123XlcSIoA9lOCwTIWRC4pkrmVxI/opd+MDHZpnh4PRYy7HyHayUh
/DE5+6H6uLJEC+I3x7GeRSj3QfLIy4eBLEpBNI4bA4Dtlxku8Wq0YHZbEuqCX5x6
q7gsfRyJmbqcqanidxe/Nnkge3WTud4N88U1/khC1OTDz2p+gBO8MvOc23+kuwwH
XbAFHfYi6+mOaq3FzyQmCAf5a6aGPqJbLAhT6s/O1tIRhmT48A733jtj1m6bCCf7
y41BmLrTB9GE044knBkkzAeECN7Ol3x6ZQfVS47GBMiMKpSsQ2FO95XrZuDT+xmP
FRPRFT4LkKQxVNcemDRVVQSm3Bu+wFayBax62nIxc423QNPlUYujBd7SJ927eY62
/3nVw2ywQ9HqP/0ZmJRSNxWhJDbwE9aunyN42ZMPGQgzrGydiER01qpJbKA7RrFr
vM2T/oIh7pv7ijzLksQw+AfsjdHO6sGKt/zSfRjHWJxnjBh2xs1od4W1qeTAGpEb
E6es1QFBKxDPQwiZpbjj8ZZun2YaqhVNnK2aguBt+AVIHqCsEbCWpCSYMy1NffqJ
jmpogzlaMA3z7tNUngJaoTwLUc3sWQNYcQPaqemieNqDP6Z+JV9WkP696qNOLOOT
btNzBTtzel3jxq4wVZZbh8hvY6q2LvK19AEDMriOHFlIYsL16qyLubVC2JJPD4Eq
vg3OkSC5E+z/ej3uf5Ns9fGiVEtA1tp594YwLwd+HQD2JkdGgeN6UMYaM0NcL5vS
+L8cpevK6aXJKoVNp57g4Yxn8Ewlwv0KdfDkq8bqwFSmdSql0lbXT36R+NZ9lBAD
X/C8yvM7ujkCfGEjvJD69hH1xMSMnEBX0z5WlIyyM7BwzzXaN09jnJ26r6FDGBAq
Ylpoen3e214no9guU9gso8drFjQyU0orq9DnemNGaVhvlUeK1Pz5oerZ1x0XDN3b
sYm+bAwzr5HjZ1duQx9CNmmfU+c7n5Aafh+OhGOZ74F25wlANmd5BnVVzEPEW4IS
tzO2J6XMXIUY5g6Fx9Pqk3LRPKK9EXq97ZbVHctHJqzhzb47PoeMNp8bpwEpGlmb
KF0B7Ls/WY7igI6r5qw1MvoVEguyoJ0SrPVnhKEbwUwhJecyw/9cydN3VQTGS9uN
r9uWFtpj9vvOSqaQFKJl0qpCent3IDZBxRGVKffHYQt92xWrnk+mAkm/5D0aD9ke
0MZj+79Y44GExkd9ydMMz0u+l/gG0cPGTDmup70D8p4hRR7hmfVRuRlpmMRk1tYm
dZ73siCQkFUQf8d9Bo/DuQRxwvAHXE2X1kkuUXKXgaWvf1e2qUyGwoFWNYpGTv7J
zPKmxbIm4DoXVOHrr8gvfUhGM1GfUF6CDfCnpFnS9FVyuLb66qdbGNOvpRBn/LaO
+QjOrrnvuXTln9th3UbwPY0zJd6jAo5VKyiDKLdlHNgbgh6o7UFQfWq7XRq8zTpE
xfFzQqkX9xG/vI3Zu/o8VrKqFIYy8a6x9QjI5KA63+cl/qSAHbqUArPuQuWSozmi
JsD0+bCeZaXAFmeV+12OBkXzumyWjAMrk18g0k4SLa3YYKHjQAZfGUAiTG4YNblA
s7BRlxGBpKzrmUe9eWN/yjQ5gLLMsxxL5cQHvwT0umIkppLMQy/rd1ILg/ndXNtB
F0N/JGb6OBeldpXZGNbvgfW0nSYabiTPOR5fVJebN/B+yL0iU6bTXaeYF2smClEz
k21W/4Cp0YiFMKfwn5zsVxr/wMCUEXloTIVD3DPDsqfz8WBNpSasZdMCHBPeAI12
dx8S/xgxzzw2hz09K4AkvB5o+y3KBMMG82C7gAtDE+XajH7MN8LaR+wjqxU2EZMG
z1Qgcz+xEcrHNtAab4VvnSKDiP1zTbP1BNbmpKfcb6+Zy+RzOpRt9LmSQieF8cIR
MlK0dNgU9xr4pu25h4oAhwINfcRYYvicmomi0YqyMg6pCgC2/e+ga5HKam8LRREl
2kji4f2QDuqffRTjZnRSyBgaDLQ5W2ENht4A/mDZnWSSob3Nvn/rX+PXefooeid1
RJRKxOCnjkV/3MacerHjkQ9g32+p5whCGOeAUB8LljrxV4eisi+kQjFktBV7XCU+
wlPR4zI5aTmZvgAKsbEOPR+AZQoeNbnQ4+cygnkY/lSlKkpyZv/dw8SHzCMfuIm0
Smjjz3y/M9qFcYdtwd3yYjWIcWtRjAe1xzpro751HVG+q90EKUmS3X96t3b5ehAy
lnLvOjngWdo2eluLZ16wQDUdiwC1GPYqt+wbqmkpmeGbNxcb7ANt1CNXLEgIImtN
v/TuHjaQjcVwCUZSWozbeS6z9X4VLwldZcbnyzAGVsU4qYs3SoJ5ZlO8MLb9INCT
HApYtQz63x4s5NYqW5rTbxCiZB1sAhaq4XbDz1amx+JSHJzuDmbZYnMrh7m4e7hg
rY+5NDd/4uAvBql1QxBLb1LkbiU0xsuW8CkI2SephdH6JVPDbzn85JuqKsJW4GBX
CvuuslKdEqLVer7mnGtiCW2jkEz/l5sOK9Npu0+GoPc5en3U8dFeVf61Y+RdsdtI
mkMiXitmb9823kuLX/Mk4kNgM2jouL02N6b7kHVdSJdQtU70HIz7f21YwG20rN56
QXyQdleP+dSIhmBFUTq1nF8bz/LgCBbv/6NQr7rL4XRFugCv68bHWbowFBNvoFtU
SqIJF+pF4FLpbUt/41J3WpARxQxAuVbuPeI1mGvw8KT7Q3S1gLo3fYNS3xpYIuzU
2p/Szr1h9/jsGUYcrYEpiYpSKeXiabnvKBvH0MKFZs39LhakEhtYsXPrdbaXY8mo
IHGGvZG0dY53Hk28uKGJ1s0F0/keigBVbQGOxE69ZzzZ4f9u6dmBCiypY0h8RDvB
1dyXAl3o7+GrzksfjIpqtZrKsZnC+JBmgEaQTlN8etDCEwE4I4K+xkYThj/SlFM8
Vrvb7/xpwJ5B3fVWGWbXtBC1l1dnXHI8LAtJdsYgXL8FXA0U2EyBzKdq7fb89RBB
uKUsUisX4nbFErwKvlvHBmUT9ylzrExozzxaHjRgTE1a9g56MkUdGrjfKClAbibY
7Qc7TBZDhki45+iLhugplI213NDdbMwr5xsvWjnNeGlx+7MPKCjW0WjNR0BtT0Aj
qOPPncUcGKVrS7wVbgzNZDdgY6hOI62dAQ21ezdxwAsNtOHrl4TKS5/9sYH43Afe
CWZ/qLuM3VNdl5d8ezcwEDUiZAnF73qnp21Ik3wgz4fd3X14Eh253cKQEL5UckIa
jXhVkGm+uHsb2HP2CiojS2x5YdSAP9GxWdGRPX7B2AFhKAwcR3DOXp6SASSm107I
ZTzLIQZVHvT6LpspIkm/FWfYIywk951iCu/oSdJHec9iIbnL+sBRYPMQumcORlTk
eMB1E5Lp2aot7+aKHgEOFmPTcq55ridOSsggpfhPB6/k2QAsyYbFblkcK0KTZyb0
i99T3Jz9is0Z+x0VMxfXXRrXpQFxl6HWFq4//DSoTSRKRl4LPq7BLRepiFb/w8qk
ey3vPwhjvP9qUJA4z8iH0CAQLfMUjmkv4juGvWzlPIu1BcXmS7kh0abjhPPsomE2
PrlQlCLIwv56knaPWPghM3kJ7ymX6cDPs75NjLMzGbtTu5rpjhcRvJkQHy95Xf5k
ztNzvvDSdZWRyqU7pKpHNlt992ZtfIzJmQol352WDc+KSotkppS9i1ay+bFSDPQ9
5BeHcQY7DW4TiM3LZOkLwm+fL4mjExqUtx3JROkcH7UXyyE4B3suQP3N+LzDP7Gv
dOXm3p1Rcqq/ARp36UJPwrM+0lD99veam35n0dW3pwMrxKnYL84Y2oV+mWmVe4Jx
WWStYfxyCPuAJ2AQUanTj4X1yTerYBnXBOF3e8VXXjtwa0veuESJRlB3R6nZJ9+g
zQClvspaJkExmOKLPHkxfQVKHRUNwFFa0w33AzsK5URFp/WAF2TQlnXskrAgMoYq
1pi7FZf6DG96OyZOmBKQLGN2hBMcbgNHN0jvx5At5RVFDGhv1KrPIe6yFvFd0B97
BX7Zlh5bwouaXQb82VOkpINU8wn1FCmrUIPZ8t7knSb0fCZpVjJ/gxFdqlpnVpUZ
Pu8f5pjG1JpX9E7GKm/yvMmSbJc4RAaY7HTUaRGG6/j8jS6V1z7ilFvF4hbGzJ6u
2gmotW9RiMIhGQKePziWK1iy3QRKM2q8EjxKr9KcIgh1KEad/eGVgKl307+U0kTx
s2D3fJMO+tNqKzpsN+ZHRvj0eEeSUHvrHyVMs6WSPjKYxClcQrMFr1tM40VImWyJ
YfAELRR0dlyCymOH8ON8GI4PlQpNlZxwvo8Q1Wb6kumfcC+N/yYB1+RC1FeXYOV0
iPXJ5/6lfRjtJ2u/gomVVP3BbGedlJoe+OcuuW+uj1OouxC+yC5m2x5WSsEp6OEz
3zdgwM4u2SHTXCLrioCpelLEO3aTkciyqQow2T0t68YO3lEnv81edKtJpBo4kALy
Wd+Biq7Ap7hIZSbED+CRzPinQy6CUbz7m0IrgHoPiigWyHxnU19w4CAFTgPA+zU+
TArI59VNZG9qB+KT1nSQOW1hAKkcZwq5nWR/1MvJpYW0CdbtiHf/5bnlik9nW89A
xG8GtQuvoMwYpOHagpqoQdKNa+l2EBlhO6OLqJ+Nct+zlAbZq6LBJn0SFudoThQM
PY4mzxwH8HUJ4sHD5kTrNZsSb21uQ3efoiQgKFU5unXcRQdAtUrK2n+K8GB8BKto
Pgc1a5cUAkSNqZyRgRqZe+RhbkxQQHWqgLv5kCZqYfxKkgxk0SAtFo9iRIRQ3Jpq
cc+FXk8FLv9Nqw4sddCj9qXS1UUPXlml/wMH8/gt3mZuMCqhO9dkdqgO5YbQxhYa
mypznfGkFbF4tBvm/4yuqVZZ0+v3M2f7fb1u06NvGpjlo995JAGZRwXxvTPo7iH9
jg4GazNYQddhylpLJkf1No/RUO3YJ82BIRa3ywbR5/tSDcOolSuc8glDE4CQUDGI
h7zQh9eWJ3hXTmZnxkMhOuzzBC8n1hjUE9hn74bxA16Ko6uVZg+YXsAAV75ZBVfu
i7fNG51dt1U6BELuFgAZ4DAYAOdeYsLezvqW+p/LACEzU4PtUa9/LWyFFbrCR36/
SzswGL4srjOu2qbUa8WqJQHkrNSWrIlz3WpZvuNC5DvJ3iu7RCEDqTqENCFOANEe
kkTmKxVXraOAoFY5h0DjZAddmJYd0MoQQ7P1Ph62Ogwh3qaNR+JuS6iYcr9tVlx/
7lfT/pDRD0vBRPXr5vpw1ryHIYDtfQ3Dimune8Da2D2sDJaYxwLHCeaTy24LECkc
z+/PYDXuO7VA1UowqbqY3FYWL4JEU1lfHwH9HVnmzCrd0nQ9Iw1PDesEJeFY1nre
l1/3lTuplybq2ayjmsT/oqtMgK6W30PPZmTdPhLZJmQ8SwFDPwPd7XYJfR63OqFK
yjYYJ+AwwRwQX1+V2M4rVgi3KdJOdfNChqvSK7Z2tC8esSX2Wst6SjQr2WE/G7yD
UPwx9ATfRFz+QIZoupq3QSNrDhiDlYzRLQB/Gl99tXga7d+yS030ix/wnp6reNnv
UXL9DymycQNkY0MHiF6CHAmJk0mKoMYbSdFDNyxGtuUGQpCU2OF9aW/eagp/N1cZ
G92ZU8XXv8MrYJF9v9TQw5+l3sCoe7jKP3DxdjReCafi4k4CDIvPMNVkDUh72CVA
6806z7naES5FyKWDkqLAyq5eSJA82jPef0GiuofBV0E0uypGOCeZAtZPdKBWUxak
i2mJjhATjfHwYPITNgyIadYsoX+b2G5BKPaU5uVA1u29JXBLvXqzUPBOrPrN/Wat
LOltfDu74TnLtgsVOIv/lTnT+KHxGILZq/daDlKGf03IiDBUOOvbO2UIAgwCdl8o
m2Q3HOGahhRSupVw4Qci0JD7wnJjZq2UhorfemI3SKNsn0nqqzs+vtNZB1wBVTon
71CUjkPWZpat7iVk0uILfXL3FbkMfksuqcK2r6g4WydMhUS2NgixoLpv0Jj2ibRt
TfZ1bQUtWijNhLzx5CJyDDhJZVkpRcT7Fm7b0H1SqGUdIuhx1l0K94Ik/ycby5wl
CHfV6/QoGd/RHpjY1WwOaV2az/CGazXYNMWRbmXFfESUI/H3haiyze4hDlIHiuG1
NdhaQINUZLwC69On4nzR7mB94gp6z9JCO7Cas4PoQgebRmoymy7JLhqrUEAx8grz
colO6yZU1vG40UlgbrGJS8EfcgMOD/LFQu8v+lln9P9JuV1868zTFOfDsTTtg4bF
axvP5kqQsSl6clcmSfdMpTFs7t3tGfx17s24I0a/AByDMUaqwD/ST+flXXesXHlb
YLOfAcsnXHm7KEQi9jdwUBEtxujARseczFKNoquBe2C71Zvv2GjLfL8tS0Tf073c
DeJA2isjmjKLqRCPE5QqirL3ZaRzAT27i70zk9w2lTczJqrIaDoTI1jfZ1nbuznk
RaMiRbQyLAfpwjV6VlekOEo7pd05AO2rWUuG427SwNc=
`protect end_protected