<<<<<<< HEAD:flexrio_deps/PkgInstructionFifoConfig.vhd
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6272 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3b6eMZvf+eQ8z14wALfTJHs
q3E8aWgVMNpEXpVH8GIRPzD5NQ/qPB94fcGqRTdnakxj1sXO2YYjpb8aCfmCb2Qx
z18bSTHWigN0J4+6hnoySetgz3OTwLOCoQv8WP9FU2Ej9fhDo9w7qo6+iVmZdTRO
o7kuAyocy0dxFsXxzGljgB95lIwxKlJUkmWWgcsafd5RtRQvrIOiieVSq8lHoTky
e0I4c/ZIFVSTMkNVErO+47iPwYr/XqjlKB7k0KIdzsns6JfnRHgqceSzBTY8qmEi
KgquC2fiPo1wiVh1VSaL4MQFuIvKBSs+Kt6o3gHeh1+u6povvp3/dCmOWPuMVpe7
lt/k4XifoI6FGYsb0s2K/p0iVsLimgO90eEXR4Iz1rrJqmkt75z16n+KjXWmv/L/
7oael84LffnamizP8jYkwL6FqeM8vOq5x5n88n7d5uo+WxUzCCSjJ3azs09hhOlA
wZncuxi/6zo7q1vmh8hBejyeLgx6MSz2lPJHWl/i/dDF6VA5nMBgiajFKmczdRGO
AclDLoeYoRCyT5u9YXAnn9We/jk4M3UDUhtv9jF012b3efowbpFRkHp6GYJ/gGKn
06aokYye6Eiwa1grJTTQKsVrur1WB0W3oM+zqgb2TL+SbWgyvZDZ6Kgste3hv5e/
tudUsNVTKppBudQLXchkJb0kKv3xDi3bamI+8IV4oHHdu1KxephtEAjRce8KCEZG
Lq02htTyBQO5Dz8otyCuYPMenGqVMjpTGFjAzlPKQPtZwQJR0hqNnEIBRNRQU+hY
RC3cW/wGh2pcU6YiB8dQQ+RYDyzLy9faspxTd8amCoo2uRTrqf8tJZqx6QubESuq
y36V3XolgVJy184XlukKqY1CW/SLlWnZh9crde3ixAMD7WTZDfgSES2C5JYkroJu
J/tts9vWEIcjThya19bYSlsv1RSm8tNNtw16t+1IjaW7kTHhtHAUw6jf6J5/g4Qa
QmaxRsW3xzQx5YwUbqfyeqUR7lVIvB59o2LxTLahg5f4Z8mPihKRCFT9+w/NVTjn
XcShmskJrs6zgzXi7L6REfF6+k+2LmGxojRh31UQyUOIrIJ4jTfmEonf4ofwVAP/
1ZQk2G7qRFVXRWe/f06YXXlvQJGHXG/1R90xEnW2Kct9yyvpzPxl12dPZjQNw1Ij
06DIxgqTJrRDv5j+HdqIS5SkiLOnNttohXFOjLC8HfBlNRKXrondco4RLKedUP8o
jr35NKw1+B6Q/zPSJyQOm5rOHH9ZzeS5p1a0/1BzgIE/7R8lp6mrA2if/vNbZV+5
WPq9oaf+UEAPUFnD43WKO8VdhHh6uSpjbTZFUzRZUOOqY18VkNYJtDLkw/aXT0M8
MWQHU0hgGR5ZLWC4mGI+fb7TahcOXotzr6zc8eM+obl99ryD7PlVXyMGjWhsA2j2
FY6n9eYqV7xCgoHghevXspaM5ksMgmNfrzvwYABoxVq5AN9EZ5v1APWyi/MrNIzN
+kBoqwm9jw+rJzQ1IX7cdQYyiHjTAn837YGlHtigfbolweq80O/xOD9Nnqtc3Kna
pDKoEeK9Wyzg5qrEW24j3zuo4QNaZ6nhx3Z05XY+oI8n0qRm/4Narg9KvQSaeE8W
bs6khrnrPugekH1JuMv3zURrvVTjr6uD9VXjYf6BtU2qfx2aayqmvzj/7xu4y1ne
xnihJ8S+ck/2EdcVDW2V1dizjc3Sz5AC3a8aE3AnXhi0xlEWagWf8Ujrt2s8y+vp
3Um5OaT+SI+KYnagpFP+BwDjM98NJNVolk62YfOQAfQDqyL+RwkLrjIhADGVZq8j
yFPNr76kjGLK9zwgcurVQDE7vnr2HcYu1/NXqTRn9GVs12AZ7ZW9f5KUYAM/nBwE
xUffy7JPKoA1ASuqbYjI+C/oOFZxqCFfAfZsXPAH1cVvpprmXdaD0k8Vey5gK3vU
vLKOenaddIQrRP5hbD+3jSjBZV125KcBDjj4MlGRwJog4htmi3VTX+D8fnLVd19x
gDDY+QkbUsQDSfa7cSSiBFkX3DAWVHGD+aEEXNQipKD3MAQGw3X+k4hPrFYbG09L
iXCmvquSfBhXujo/irHMl1r9nCQ1VpztqR73CkV3bR9FNZN7SskdI13mqIQM6SHR
zHeWE1DwGlzbohCxoSiAqzndIhKd/ha+USdq2KazDCBR4VBGWaEBPSadz9436pYf
mJoURY5fgunwLP8TYZb1Ojq2NmKUYSN1X2AG8ynVePetpUvgjZ4dT5Gw8MRva/ts
DBk69s/POoBonadfHPEu1dWOq9s48+s0INEjQo4MOZJH20Cvm3B4YiuIYbFisjLZ
tU4QGZ0pG4PC6ouQbJRnKYF4EL/ywVCgWhPf4L7LfuDgM6Qu2g/AwevbSh3HERCL
tJci96TtJAp4Ur2/cK7D/n99fSqc09+iKUEnkBQib0CeM9aqTaeTQiXhBtvYUamn
YcTIgjkc0r4qajoy34NZoSgjph8hrrB6r73nKYPwrj/22E6JM7U/DBoq7a1o4uOT
cu0fSsZr2nozKQyPcewZgrDaEi7/Ydecqdq2di8gUXTdPudOGu68KN62+3uqmCEq
+4yWpIi5SvRNSkUaLysvQpwOsgizB+6p1Si4YesTe+OuJiCmXbx/Q+hUUdNJM0S5
hUtZfsI6XZbfx6YWpB+ZLWdih9U4ZXIwBBsbOuuiRbYZFQSfuSL0hLX3JUqjH1se
wXjeK1PG8k/uPfZ2zEffTKX43kBfe0VMoP2P0Ms/C6sfcX8LBgmRBoAgWMiLhtiG
tz9rMkXoCGsbiJ6UoxVBKZvv03+0n8RK7if8ZhyvIb5jBR11CMsfoLJzbpp87rzr
KWNaSnZ/++g+MkC8/sUQsEEPPlERzETS0I9xGGsBIQZDZEbAqwTFksxGPFJ3Mr8E
psApZMLQw8HQ+KBCBxexlJ53gssgee09NzFzGAI7wG/LjpQw5QpvgY0IOjo9F2ZL
c4TRS9tU8iqsFCw0f0kdZaYb7CfpKn58FXlOoVfxmfNeGho2+vPcJvLb585W7Nox
USE94VCUWmI418td7tR+iVh7wiVD43+H8opxmUIK1srawllSK0g6yWaOHR/hQdAw
O5Lasp0b5a0BFaZUHQ15VsUDKlO2r2CVYnU0pNUVlQf5H67yPQPIJfltEFGpoaKy
Sxdk1OPkPj68NyxqC5gwNfePSTv2H/bqNQ/XTFLKM56MspgKOFxDxCzSfC9/QvV5
7DYm1kcSJiLeJ07p2bIkgjsjW/2jrMVslcH7saK21rfJXvjww+Yu8j0e5vDo804O
2qAOc6nQLTs3FH/tSekUaIiDDeVoSTbzWypCJgL9oi2+BsjcXaCn1oJXiNdnEPgQ
JWWDkW/XsjjmJrJTFRV5Z1sXwh6uQCrHgV0H/zM3jSWHoChXxjGgRV7SmkUdoHAj
jr5KLpFXriq2dosOpsWwFHQcEJS7bjeOxa6bqk9zQPJuqEefnDScuj6I7IVBlWeO
jlVb54WGXiR2AA/wwGUoo0entFINLsw9EFh+oiAj+A+alCe5p3PrOdusEgSrmkYC
fbwxLXoTrpJWmxYekgs0DF+07OGVkmVOKVlqYRz08hnCUjpSdT6NUOVAsWtrpg9X
4D5EE85QHaFjHZAwlGLg5/xlAN3XP9Ziyr72Cr8w6AIiQWPZdVLsqE92snvoZF6J
XokwPZ3sme8dF79VA4wPryPCQLAZZsz4IGi574Bwc4uWeu6qJPTIkkpGGO5XOfS0
UhBTd/DYHnrTi9I3rG4ugaD6rpY9HT6ulk6RmzsvhKGT4tFYSi9uMp5rkqXhJkEP
zFF9thJ2GlMWoMhNwL5Blo3ZmN0b11DJhAHTf0y3x+Wvb4/EVDzftmEvql3/aWwI
Dvg4cRmPRghwYB6lUOx4nWi5QVBIrkXg3DhmQOmMkISz2/MpwHqPNgR/B5nEBsIK
u2AI9f8VJHlw7x595MtSkT4brrEHeC3Uopx1aosm88PhZ3+yeCj5uXM3qDWiQ66y
IyFawvXjK9A53fpoY3jmvOvuoRRNr3jCpCnXWKSxBfxD13hsgU69zou+o3ex5g7T
sp45xTpGR8eWwhsVuZL8tGbQva9BEYbi1m8SWrqpHl8eW4a8JtnmEFRa1TiW3qfz
eqp5FqwdrvvDyiyg85ma4oSp5NcvkpwLTmdtXFT5dG+OhxLcW1FPIjJzj3zRuozn
9ItGZSVqyuenDKh8/zLEhpY0ZEm01XLC3e94eSGA57T5aNGScM2zHbjrTQZtAv8T
/wVjzSGijrkP4UKpCdOLsOX7JV2X8KvbXSSWLrZ2VZBoXHOOqgVA0cbiAp6rlLdg
gQAVWHUjmOFhRhAPpWjYQkmrDp4jXBD41OdgSl2lIKL7f0hpRwFmvK4lVO00OiWQ
rEm/UwXhg31tQqJRLTRr6aIt68xf13xTaJ86pKxZPRZeOvFQVmag6uxezgzPKOor
UbOGCCQMgugFU3aVMKZS6qzpYtSBr5lri8ljTFHisV+J/yb6VmdVTWJL3acCtf0p
jZtmwLkkid6DV2E29pWi9ZVTK2rvAsKRs+Rqp61cr3HHCN69whGCqAbfGpTwWFR1
3Ciaihvb8ismdgUfVJ+CE7Xaq2rSYIwpclcGxOrqxO/BX1CQAToJzxCjDStC0gW8
qLd7Bg6nQZZjM+cOsz8yLKogGRyzP7Z/FtipC6CFVvgKNVRBNV9V5LLKTa0dTfaX
/Z4sG6efIGMX2gOdZXPrwxuJn4xOBsacy46oKkcVaPzUanUB+fuvn0x/gBCDOieR
6S31+EjmS5TgwAWw+yJOqzgVEdRnk2XhwjGeAybm6ZBZ7qYuM2Se64tS+h04cCoJ
QJCCGBKXAUPXP8QYQv5CwoCiHy4i4cOYiqjxgl+KsJxFL6qSnaKi8QIsWXtfnMip
17QLwhbJ5zrYFKVDFpyzZSj83OCvELvWhNMZXtTjc27nKRzuEFrPvObKTMeIvVvI
oXNw7xpHA33pOtMzAeaBkVrE24lb2bqQSQxQZ0Kj7xidY9Ryl4yXlxjm7BBXUS5R
13NWl3r0sMpGDUA6CFhxLYOqdiacKx9tFVNjvjYsycu8VCIOo9plv1DWaiyJ6lcf
LSKDNrcr26Y+CIuAaLZYkaVbml8u8BqkBe7MdqcgcyICgqDbVdwQlhl/SHWF6a28
3C69vOPPw0SVpEyiM0YnLY0MFhKVwOQGxOBc2Gz9KEmpZ12awp7q4NJh2kX0i1tc
9kMd2BcV09jK9diVOrkLUsGaHgGrTghsYGiM2ktB0r2jbY4hroQVBCjKageACcNP
SeZE+Fvu4OK1Ad3ThKZ45skd4hJYuUbDoVqskgMbamFnCyDJWtN5+50fCQEf/rd1
iHE8i4qZxqhFaJEkBnlNQJXGt2UKLDOTX9R+EMCk4kpCQOqoZWLrABye6AIgTt25
Vaws5Tgjrhujs7fvCYNBhgSfWjCO/g4dRuUl5EHiD8XcE35jW7AUWx7eF+MQwuX6
fCFdxqPiSWI1+fXMJTp/MM9oljyt9B0Hxg9J6h5NHSz0svJjfFyRhle2SDegpYH6
tde7k9FzfLd7S8bfV5FunLa7fmZH/QOCElxgFjef5QfGoix51f4llXMQFZC16JyB
Awv0SjTaMZLTLmDOgPRODqRv+JE82qu6djIZALH4fteJ7k9677O+ZX98g6neuL7A
C25DRCxnYMUmEq5M0QlUNVxIi4zNqmnxnLbSHgHeoT7iGCRMHLJ4pYWkZ4+xIhVM
0DzO/Bs1JKZocdnUoGXS/9uTc4pES5y/z+V8G6gGSd8Uu9+EajYq6PnTXm3aq0Wy
jYoejuMb4Ja60uQdkUoUCwWBnzxOn7/Zi/S6yI/+EC1S+wvEO08vOD1KufCVEqP2
67xr28HCOXR774L6kU703uoEw6XySlYJ2j5rXB3bZ8BRjJ3wXB6gi5vKYSa6/7N0
u3Cq/z4KMiWpStFZJ3ykaZ6V8mK3fvlisSlk+GdCwtaCGvi7AbhRHPY95x/Cjcse
iOG73fIjwBEVJSOf+JOvJRlx5T1NfKTWiXluVbbUji16fx1P3lqm07aYPjX2kvLB
NMQ3M2jl8XZBf0wv49xQlRExmeK6mcza2mNvomGk01cDEPjcjwh9aLfHYkol2M0K
w6rQ482Dj47zdVWWPfsMnveA4Q4OyXRwSShUCmR+XuFpD4NA9mQ/y0PGUxNY49Kh
DUTe9dB8E2orQ1g1CDYsd3SNTZcKO/8MTFRkDT7I0Xc5u+SSBp/gUbSSoXFO/baL
Gd+JREJmU10fCQwBUaGOK0YLVP0BIJpx6ttmd3m9+PnfOriKGvuLKaAn0dNW62TG
X8LmdRC+zxRIWZR2SS7ZTPobOoK/j6gM600UBFTtlf7HGHNDX1k+w/t0lSmp0yTU
1l/bpdxZuTnJGGJXjP5s9MwrP7Nu1LV/gjv0H3ZYkTUmjubJ+enN8LWcluij2crJ
YcjtxVT63Aa4+5yTTu1sJAqJoKRRq55Px4WlhEmsMdOplFMRHNYEgSy+WORgoIsZ
Ri7rIRXcVo5gF/6YgZ5zQfvDUFJ2Yf20Uyardsn/u378ACSR/XDJDhOYQ2GZVPUn
F5sAqOb7xe3RVhsd5s0TkpXbwsioZ349oaxdyukp+jVR4kB2siDhAJ7ByGJZ5lwR
o0iSIbmcKOmjvGbXffwU/VxJmqO2ZptReXRTLUQXWDsuAzuizLaVhB2jPHAEFjBp
iZ2Jkq+AFPrueX4BFVCaAjQAyg6UDh38OpT6fUkfOzNW7NGfLKmDF/9UA0TcQkUU
urAdlIC8kXAE+rggazmPa/FJYLQ7Y9TLka87pcikLwEJkJxjiNwRRxRlvQzfDsQl
jBWqel4M42UmLjc0EB2dJhSNcNZXW1xHov2nY2CwbKru3oDn6DSNjEn4r+fSRuND
PvxzaXhY+LH4luWiIJE2NTZ2dQBw7aTgnPir1Q75d0qJMFAdX81I+qSZmzQJRUoq
zQv3n+jiK4AYlFJuu18CpQPI6z+20Az3oi8+mlol8sFaeBUmOUiIeGXjRwbaXfR3
oTKuyYQLmAOPY+XUYAdML79rHnYOcAU6d/jb7x+jQ6u5qBiPsqNMe+qIEtdqZOyA
UHlhoJcxc9YHsTS77VfysZMAVU87a4J9BeZvVdJbg1PGUMSQIxOeRPpIUffQTHIQ
uSoa6MxIT6D82zd/SCm9n3wMUZxDIN4OwH4jDBXkUZghm2XS4wy07nM0szs1ypEx
5hInT84jXARv1RljmHqAsF6C37l3W09vm/DfKq3/h3cvrEspuXkeOmqA42IPmJPc
ARiaA8M9BTLL4+qloP2Jn/P3T9VTB2VgUkca4Rj+g7E9cJtsbrrIB55Vv7GjbSZ3
b6sMs3XgSzHLwXnRRNDLslszpiFtusLAz2K3LhXXoVGjrswSRczZQ/4c0DvlYJjt
mpN+phi+IQy+c6BDAE8B68QJy40pO+fsTPAoiYeY64Dme/STNi2NLEX3LCzA9A/l
+lqpGBVpG2C3dNXW7nTA1kNJ2GUIqvpgj4bE+D+N6utYjxqNkRipmvltP/v7nEwO
1gN0YUi5ebFf1SGgaR1PCbJEv9GiBZ81dFdOuLeNDezgaL3o45Z277brEbbH2os8
5oeHgAYThu10VpbPrRvZvdAU/D39qLyGxj6XY62cMwXWH1In7Ug7CL1xsMyIId1D
prNjJJBURco5x9AYG/mBjVCCApA2aRRXEwVr3egCn/Ay3PDxo6m9h2vkHizaeviX
Dbd2Cmna5BxS7Q3rsYk55Y2X4NG4W7U0lnI9gEqmoXnG0gmNDpx6lr4YESIhMrSl
SoE2Wqp+MWpInOK/M7ppRhmddmwOQbgmdy3vS9pB+YOOAN9NFsf1v7uhzl8sniaD
+A6HKma+Gn+pwC6OtdkbHjpaK4ekqMGcfeTpLNArqADPcQ4ZVlfAIzpDZgc5py5d
DCNIOHVi5Onzj33/v8ZMkvCKu3Of/tX7cYS2ZVtWFmkY3bfP9CGRMWpaJS+ReDUr
oWrm+0bjv/ECaGHpZFVKZHnZFE4jdMBP7msYx4OFcUrbAT1qvIyrOd25iwmJ7TUw
/1w5LFH/mGYi8EyXiCet2tnR6Qf88Bbf63KUbXroJY9vl2yA1pVLOWuH4VisiWq/
N8NhQrt6gg7E4WXgpVVuQwFmcjCAy0knfOyKGtfC91wBSPue1R6atsPpkGvVpzRi
CPqGrJBfLcbEUOUaa8cXWXtr90vch7nrQGjjENnP1L3mU79/UJcQEfwGD1YDyDOG
KJH32Afg+yWyzL66S4oNUowYM7YW5trtu2Yn+bh0VUk=
=======
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6272 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JXz1+zHgF4n2s6TEZD4KtuQ
ATkS0e5WlIVeyjNZ91Ns34mGmqHu6EGvs4XJ/VDUJsXeWBHwg8UKR1sksoBSJ+vb
8Wv9vudusuLMRLpQGEvrstqhD9ZpeK36d5KEDqk8Hy8KZjGY7QNRQI9ycmRPYFVW
JsQNsBWWuA+OeUixZeMPn/I7qCsD1jTDptAV+1fAbv4XoKCWE8x46l1AZrHCZi1J
n5LMoVjB8uPvF//4GS+gdVNX4dqPLWdZ9nK4sxRSpoRegkagvWHAjseimew1hSoW
+HvvHcXkCVf69F4fRPFvnU+tiN2Heyoeu/jHmxC10MaJWDUKbMtov9FfIvBDeGrH
AXlUBecASUw8rEVE72OsOoNn4grOGoFXWTC51LgZqoB0cIE/Y3bwTElT0IBy78f6
bFyiWr19rCvWVgUCgWEPXodO6ARP/A7bPb34XmfXqDuH5jgGytdXigCrcRebgDoe
wLeQLd4gkxgnOA7mRpwi8ehE+WlqtppqQMTQyV+++BHE9J8kdCy/uiWeOyjzWkKU
8QB4+nSD6yfC09kaePH3W+pZ/jKq/N4ZYeli5Ub8JPUIAN6XmBQOxd4wFBiF9twK
RqhcSf7SF7PUB6AdNek99rT0igrnUR13UF/AqXs/NeGUbdc1mwfCt3cDL9XXTTSD
3fNtfvrCxdRHQXPmBTXmqtNkI1YAJja/UEn+9IF4nDE2cCjFqdLC/pR8XF7/aFvZ
jDfNWqmywfel/0wvUoCYExpOGLvbytV/SM2N6ArM7bG89KRXWGFTQ4yiDPlqZWrR
Z62s7pNIbr/OIp8sLpJQCJX1NQC31ZMsxwf/qLy00F23da6OYuYnNMIrv027VHPV
RHLV+HaabBsOXbxnWrqacyNdHaYePWapoIXwkVlMht3CX+JSmm364O9fAwapO9pK
4v0BCSwoo0BB26A63psUVr0mhE9fedDne+cnRX5Vln5iyG2GbkU07CfB565Ba4RA
4Y0/lYOXPn0dKwCApJrqDJCKDnqQtprdgVL+EjOYsM/t7/DzlZrKaDEGdnoh2kBX
CfUDDRO64jbMcXmowx1o9BGlUJhv14kltef33OBLxGdCJ9nxmsRE3NafdinaIxTr
GjSQyhBWKFpe2oBmXguYRNgtKEaVyBc6ys9i8rLpo/vqJKVaNZlSzOL1Tc0RDV2d
zrwFPj5HkmxI3MnNaZSkQzy6QJaKv7auS2T7RYTiRRlYC8XaR5COpIKud7yHwkc7
UsrMtga7stbyzC+wDRQNB6AUo1Qp4ZSg0z2LvZIkZlTtGdM/BVTAAE8vg5E7cbc2
SS/BwZosgTQQBsHI48cI08zy41CRLe7mZpDlXf/99lVsRb1tEDdt9uOdbHCffwuS
VuF8slHpZL/M6ExHvMJy0x6+GgiCtrC7vxokQauFTj2Qb9iyR5MUUKuoEoUOLMsz
OYfYbZ3aIa80ELYq3ieYkGqNrC5oVdsTFvas1UD9PvkDRcfBeLwODYDNmQNTjEHS
qf0S2rnGYqRrEYANw64MxeUZiuHwqUCrBj5gOalu6J2O5a4Zaf33UTLEZyUBNFmH
shNqMN4M5rgOR73luIsWYMhWMdzhW1rqWIvaTuRHRCB0OZsq7XxXA+4DRnDsqEG3
2izGyJgKYLCiMYnyO9h7v/N0e52t6vMQdCC9imFHGcJIcLntsBaBeQcbwn+Urhrt
ULaUaW4npC0butc4juhJFFl5JtieijyBtwAnKlkcXeeQrbTRPT+x/ZkvMu0CpAdo
W0LyzykxKQBlXBYLc42jwvZ3GV++ihkn5fJY7ysQsmZqKgUVYVcwHhQi72tVS76f
wqGsxCu0LNiR5fgrTtlo4n7qKauuKH5TNCYgUloTF2AzI85QnwhNfCVRW/inGHGv
X56LSPzGWtbL9VyWbtDsdEYvNmqM4AgkTFh91w2Ihfw1xRZyVbYKn9gcHhB+RBOy
xj6mlXJQufrb5YYwVWhUv3QboA3HBogLPAIzdzP3sYYQcsPvzMdhakN6YAS0hvQH
kXDWFCkUsOkHpQzUor+A9DjtGom2B+d6PTe345Rf51WAwXh24/JkB/oUnWnRwaBs
hRKAJz7zRjYHjbRQ7x06+NqKFVUamqbBH8QlRYfOeOZZcEgyu/uTZPBnvTGou8ew
1zZO9xF7FU76NJTPsvcMn8jkhnXWZeJHTBO724pVNoZBMLzxWWAYQeJUOq92MWWP
LnoLFRkpLPaX9W1kkkblHDU2vlmmntbbIHIL8X29EA47Hmt2OgHozZ7v+dRbdgpJ
Es254kQKLUNMVCgH28yYBsvN9qzgBD0eW27pP40waLxaluHmgJJgRmATDj2Gb053
rpBvWtFksxnIUtC1f4YaDnyLOba7oRX8CU471lEmlrdp+cguPY70arIvStFk9KiP
HZ4S/db8eP1L9mllyeiJbmO3ztoIqVHTKQdQzSpy+fVuZbXdqKQgS+j3TtW+DLEg
dTyleffJYsgz8P6UMSTRWyuL+ZzZuiLgA5/s2I+WRXXjVj8pYDs+ekfJI7z87ENR
NOkTEBG8pRV0b/4IN/chuiSVQfdUGPQ8mLKG1BbNZcJAy/sJg/T1R6ujRf6sj3r7
VJocg3fDjdoSt3MWWjKd+bqYhhfl2UUeTOOi2ryLxhUsUqOL6DC/66jP0b2xQEQK
8luSERYrFvbYsVZj4/7ZCdBZQawJWs8MXLFHB2IQHQbttc6sJTB4rHY2Xv+C5rku
9tOBP5WXcpZ5fklGq38EN45GJP9UYcA2bZLtMEMGwcwQ88hHtDuhpaFnsGYuNOAi
KV+SYxXsQwtw/gMXlKUBLkClS2OPg3WdkMRu9w0PBwtcivG/Q/7pn8wTcHjH4iHL
42srPsCc8gqxInM7H7jDe5/8TU2OYzi1kzcyexVHr/L4JY1pOkEn5edoCUy7YzNK
2qpKswuk0GzlPzBQgm0VWDBvltWqJvjunPSEuTrluN9hw5GXjuWHvhTLSYhI8SNC
+K4KcfVlnWP7VH+MaOR18TDK+gutZbzGzLPyV3p2j2xvJ/DCDaQvM9jDfuWCR/bN
qcaXglUtWbw4SymVmGxPaAiDMiuv5kXxpuVJGVEj2IBoDOa500iYNFU1kRYj46zG
GoGteCnYT6G2gdzij6Pdv4vs4AZyKaTABekKZgBC0UINDkd29Bo9D0XKcW5Q07mH
DqvKl6OLkjJNLossCiJXhiZ5x7QiOgqwFHkCJ4i7cKsmX1q8roLbgpAHGGXW8Qlu
xxd3vjH70+xjjf8XaoqqvzbdIU+KoTV2ZtZ+ClL4+GLO0BbL5QtZSvCBZc2mQW1u
RpblkoksWZWSoV3Euh0zS8hh9BURik5vIXLtg39SeG5R/N7Th0Gykt5UUidTbkDI
+EROAReKStP7vzS3JI2RhFEiIGb0mZQHRQkJ9lSsRHwrbXWrT2YgaY2znTZtnOyp
t17n+9r3s+3O/FXrlETc1QtImbICSyQCBe3sXHKqKR1y057OJjhv24BDWzfxQ/RQ
IzG3mlx/Z5S7mB8qak9JOqPDV3Yqw5Ho2LO1v7bq8AR5BYUPknzH+VuscwBg6H0E
kachUNT0hiMBV0Xm9h2uHAXzfjlODWQ1VRKvPENnj8vHk+RgwV9zp+ThG05ygL60
CEooXj9N9jGVcTNOJuk9fDsl8XIgxyeo/rqsQ2eYCy2YM/QZXSQi7r8nYE1ZDhD8
tkF27o25PN8jHIkZHlu/+e9aKec2CFz6fwJgrqrKwaIRdTcYq4LpzpvDxgGRxkVI
Wj1pNHvGiolTc/UiWbGcdlPAqxhpGN5szLWJCgrGKzghdiJgANBj1h4MfT4r21/M
A8YZtVQ8CbNx1QQolP4yqcTflt1T1WIDpnVuwhmmr8StTs4P+riPDCVMQ/DD2+Fh
5T5q0dndey4AzhNDfRwwggzbQQy/auW7mCuB0dcJAhras8HOR8F0xYhAjgZTcfp+
j2sf7aNbDUTusUrg+tXJp1EnNNoWxeL9nnMgnPDUG4MbAU17hqSx6oGLmPfrEttl
bpp2RLhpX+OOBnNqnHPaHP84MFhgBbWwq/MNI5WDLP6tyFkoaIdTq++dqbmc+Ro8
1sEdfuySgutvpHKPBfgg+Y2JfcYvTx+1RF21V25IdaaQFv+d08pdvSXIYYl3VEZT
fKjtOOk7h25aWdtWWxPRrT2kdOSu6AwpR5sE3Blvqczt8FWYTRSe99z9R+rFn8vy
cQYlVwg6Z4VG4kCCN+7Jz0hr9poCed9Z81VX2BcsQFQvguIcGHj4/NY7QgTiXRrV
lspXSUAqMScBzio9l1fj6C1nXCDdO1jTvjXO+APjiOcY783uKVRkiwrFaD62zfwh
8/V4RlDXMMEcU1m5G19uUz4yHGWNXy60mAnauJamitHNbl9mDFRz5331IV85Yu8h
/PkDKk8bR+xvqEe1/L/iDY7FEuw6j/Fat2pxPh4JAWzw6qPbMZfhzUX7KVqRWdRh
0c2tbvVsX1/OTtJIMQ7Mrv0CRQENGo7WiK7gpRLMbb0oD/druWEeEO5ZXyz+2Ewt
0quZOJd+v870o0p7GJVr+NfKE0ur2d5G/c532By1l/nEy2/pva6OMcSWf/JEwCkH
eVv8cXDBqGWXW4HT60Rpv4U+IfDGWC7cS3TqmqC8Ci0nITjxxYlw0mbbfq9wCGMU
ODv5QmgAjOXvYxWqzgdtBqK7xLOGpJ6LwMrfigxl1kKH6MfPsI9XVAnRhnnfACYo
UHl90WnqiISEg2bCiXWJxW1sWssjKRCkdl9X/mWCL7lKmE6A3GczNjTn99bqeGZI
CyYmxSiHsuyD3B5/i8ceIaM6aHn7PMhUF5VCUuxvKnDCIOgvNYa//cvb24dnlCo1
MO0eCHVEWlNUGWPz/0mVlRfFLZoJuTvHW6j2VjhSSlFLsgQGfPYoeiQNT5eEZEO0
hV58vXxmzSRSe0HK9GeWkjt7/zlW/ut9Ix/QYxTHfoqucDXVKjD2vTS3Tw4DRy2D
ljMJ6EYT+wgaopxGdQ6oJy/7+KloAX61NirRP4kMr3thS8v3Hz9TWhDee3wjJP6K
07LXMTRkL4ulYTgwJum/TLRhWgj1QFuNL5L/cvJdX7MZac7H9JHqpBFOP/9V+Ybf
3wzP6/3X9fI9Uguxkx5Z3oZlizj+BCzD1HRLkyJfd4FERtcMecy91djMsOt5qSM4
z/TklxYoRgTTTvRkf9VaaT9A2toGXfmknCb5qTRv0c6r1lVaFI1iTueoCpxj9Md+
KVeQ05WIf1Vw2IGLya8/xv3JDO9Wu/+2XkfcZAtyD4ZbfqgLlcXx39HGR9XT96NE
SBENFvTCVp6LKyM8eUei7IbSsPKtOI0fGus9QKHzqAf8otKzblObqdmBTmbYX44r
L6eNdljoDDmkua3Xi9/l4gYrqEt3ddfb3EL8AaAeLaltE25h7Tp8QY9x8RxQoz0V
WsYD+mZLJF4Jz/UMHCTl0yxJk9ItKstOQLciAi2A1aoJhQYNtk5GbG+Ex6p+JUus
wFoXz2lLnbVtNVDV0p+RMEKmAWK8Th9MVr3i8ufCasEt3RE4a/lsawnhW0Bp6MN+
rOUoFJM+/rPoKlHEyMFuiiXcFzXOGDYQG9jy/hiL3oml9zPAjEUAZTilwrwrXBtv
VvJfeTjqaCpkOELIkTjXYkTuw6IpUB+DIXGDWTLGTGsN1cOXQtDT8McPiOaurIad
0Gw2+wddhbKQ70R4qmIVckp6vyT8Z5uSSmfxwvV1O8V9pqF0YaquiEbenrIYHswL
aZH1ZwJs02MPqzY60ZBpSYtryoL9+8ODKva6QrQ5cAxOl/2u02guoOW41hq2jwnJ
5GuDpc9OKxTOIW7xy9VG/kQtNP+/gNNWTbGcyBg7P9AuJRL+geIeNKz2ChSpB/yS
ZamGIcX0Mg+qHVxwAPmimDuXNjboZl9z64KS/B/lIhQJDzFkESauoiaJsm56lxyC
OmE7HKZTD0HyPiI0TN/g/ie6emRUwyjNYgUY4s0XFMn2RfXasXxigJLBl9xq37aI
+Tk0v/3kEXxjk/o1cRHRvbZ4Ai85R3FutNP2tgYOd2tW6ZiQcM5cvl7nFv14ljv7
A+NZWlgJg19iHj1iYDqIyg2wMgorATcNrYxZcUOXv9mC4ETPtI8iFkrYr0VWv6fj
aWFpU6MrX5+IeAwFxaezW7HYBpG75RtZfqS2RPrP2tV8qpTXUl1EBotHcpcc4d5e
X0wj3qFZtAsgFsJwRpSgvAtIEf6w561fT2qD4N9If/o6NbKgRalOe1HBrjHZBrzE
sdtFkVg54G4jmK683nXmb8mqPrmHZeTcSJ+LpbFtNKtBigJAelAsoj9Vy16Zwh8+
wX4MWvzFXMMDFa9ibqymo2M/Ztc4JKlvlwxR5fXXp1hj498CAxJZ6nwcxT5TrXAD
XaN7983I+TqdEtL4nQ0OJ+sBD6p/39nsAValr6zkoTS865Ou60SGA5/yiSTGiasM
IkDLiR0jo+FJTuBLiJ4lRFd2C+hU7YHKOfkSfYkdtzDS85oFEtojYYVs4KoLZOnA
6XPe2DgoHk0TDB175m3JbqznsXXDzxITPgZAea39K+wMqM+p8Ke7FfGg4haWhgqg
YXU0S4GMc9kcq6AR4VZUiUvMdJCavomzus4By33IK3A9VciBatOg5Ql6tdPDOBEH
b19yVtCBKu0uJ+uRHWQtJO+NaoPaiOhii8fdN0A9nb8BRUZp3owTTWQfLS3G3Uew
o2zbLA962pVOau5624xu4GbUYBF49j03Wghq4h1VABcYVeKdjkzGpFE2ZJt8H2/i
vAHYepSSdrrAwHIgt8ADCMXYCkv+XpO/wr2WuWiDPyjjUVXY+5lhdzOpAUNS8Zy6
v6oWMJoJ226uB5eAm9WhUOhwdY7M/vgqBJTUOUqPeSXeA7+Y1VkmXCPL98Q3hzUT
3H/rW1OnoG5zzQf4Vwl5LoSKyGMdY4zIpE+6+GPfoUaMdswTd8Ii4OGE9woN3/re
p8+M67uVqP6diBLb35cObAodA8Llh1X7HPOWHVA0O6b0J+UmD+IFmC1NSbS1CsA9
SET1/FECe2uTDMqd9OACCxjVGUYyA7SYE4KJEF1r0/pvf4wVsFbptN8kam3sGLkV
Fjv/sJs62WxaVT9Z8vhid8qwQ2Lm/Xs0KhxaTxbBhXt9DdwRSPW8a5Uoy5sSenVH
JDtMTMjHdErxK4NOjXRHDAxjVbzNYztGgrMVH9Yhuh5MWXsB2Jy7kmP8EAt4OFLQ
Hk//tfbqoWsAtLqIgTenW1v4QJOu+zpI6i4YU1tFgpiV1Mb/AK21hKGq8numy6vb
1kVR9o8mqA80Qt5RyMmiZdM33VSJar0swvEOTTf/0eQTU3EsJYt7HjoyrUDRSHyT
Y/vaOzAbVWtIyVJRqFcTWtkq2gn/YlIzcvCQ0vqqEU3j6UIiWGarmc6w+sV4ChAu
7nX0ooCK3umJJsDh+SnlMxh6qxXqVN1esaQnUxdXs+7hTO5zaQlD4/In/Ct1tMxn
4sbu9jbAocAg1FBwY4EcWFXVcOG5xmUIoJaOVGh6pr7OnZSkBKFHgCZODeKtUP/T
giPgQIdg705tHJnss4dLvdqIOiAuLja6Rm7ST+LnqF0fukTpQB3ptdjNwtihBUob
1opzZ9uKVhbbYHTr9VfuSUaaqBUbkN43kQBB19+hMsI4ozR+BvmP8YG4FLnFzhfW
EAmCtnnd8lrA/ziIVVUKsw7bg6xNqBpG9pAOvW2jdpvWBeyESD7U+jvMiuj68axO
FSHVQfdurJ0I8UySTzIUJ94RPthEyJYRb8M3ExUDaTnLVm5o1uHv4HgQehlheDPL
XK1sDZxoTMO073ZK9epVaplDt0x32iO8AQrluIgXLYknrlanAvBMRMhbJ2cjSJbM
UyCRvHGMH8CJmzTM8IYb5GAAr7iu5imbIOjRyTWFaoVNqNi++dPbnbvpeqezRQLw
ZKjf3CqYj3Q0ZgFoHghxgKpdds7cEXq5l215gzkOHuveUH25nrbIYuXpSjG/HrVN
vV9MjSnonPfhDY1KQpb2mymkdlZ2uMpwFfOZWJibyKtJN8XnqN69JOhb05D88m0v
id4CMqH2G0tPb1qMqwhB4sHl05+KdV7L8EyA+gPx5m8N4qnHu5Yclvf5FVV/flbj
O8vlLRb5hlJWdlaSpPQlWkgfeCymqGEeLr0JfFIHFMOzmfYIfqFJPsO8u26gKYZQ
4saeY0MognijV3B/lJraBRpne/hdPjN09yeSxaIYVhS5u4K1+xBSCvmrfqY+VToB
SFEiqkWrZZot6+x4dauFNYRGgEkaUp2/zVVs7sX1H6k=
>>>>>>> 426889eb8ce467b9c9a9f74dd4af433c5046285c:deps/flexrio_deps/PkgInstructionFifoConfig.vhd
`protect end_protected