`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4368 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
VKWNRQF+vfUNEEp7apOJOWTMCIpXUNmSX/EnicpWiYoGMPLjU0dbQ6WO6th6vqnP
AdICDJkMe5eMg3jpRrP238TcJyfWf02Y/LxSVYK1615EuaC/uGmTmTdgkGRuvAhP
HxKsnJIfnQ6FwnJwrZczr0iD/v2IxOFbWiZeO2xFHzZbA6rWlCasc6rUqxgJrqPL
FKQYawtUER1lvsck/xovTLHCfAHXoqZDPx23mn8AimKEHqErIx57chgMVKKucDqT
FMjKhlsKu1MFbtYQFxunD/Oo/eDLVDtCTb4OsFveYi3F88TLVtJdZetvSb2e1ZPu
Ii1NlNVx9s7S7PW3FFBc/jrik2eCCIrqUVFqGl+njT0/Hck2RVEba4nEQP4A42gn
EGEwV328MQOBtRLdL35bZmhAR4ECyUAbL296gkZrEW0k/ziGc23n8krMA7vVNNHP
OO/YJvo5yacrkPgAUVYORBVg3rr8xGHT3OXabl5ZbkHyTUs/X4JX/VjiWhMs5BY9
DtqRpWowWePS5XhDh5CSoKfdrhuqCOGPZakJZ7GY485JHq/i3Soo9oQYFlXC1rvG
mv9eslJayCyypFjrjRrlcIDEyAUgOWzfA0pvqQaTVh9hKS16tX2lvDIljwpR54pe
O16Af+fkHVHxIZq4lqBuUUWyQwSIpNEC5Exq13l8i72hD0bWJyHl/grmzsoOatyu
ZEgKEWi4snVB/T4jXxaZO3nL5vfzMQNT1MhRdTgvOdLERdzNTG3ge7+rG2sKxYwC
1d0BldppwX14vY0JiX6Ddb1/t6eHjYjaVhHul+A9ujNBOcYDoQrQWvYW4JLhrqf2
Ms0ZL63kv2gxPGBprfuAYJKhd3EZCZm+DQ1mdRf2jIBK2aCwlXDKb4exJogp78xs
9zMZR9FBWX2TvHjuOI8IBN4WnWEphwWXKAwm27w4CSOMv6hFLLGozFlU/K1BVIMZ
YT/7Me8KkY+EO1GHREZBn9tffOO/8b37yi8N0QBGDV8pGIzYQiJBvU0KsrzDsnGw
DY07Se0JgX1j1h3Mawqkt4U/dMa6T3ZM4l2YTIGGrBbT4d/xaHYLOxyEnsAojNDn
rQyifE1spJiz/0KdOWJNACCBcxKAAu9TLoiIcLnLUuIz1UhSLGayIKUsKEN0zXFZ
urCYZN/wxf1SI0orKFokUyHoGcBzJj0ZsTv6OrNoTvtccuXRTNTFzIeEjiBAO/hl
jzGs7pPxebEfNYmL0cFJBHnz2ilC5x0TnAM3o1ZuBIW7980nLmNUkrlw4F/yLw7h
CZompovIhpP0pKUn+0UgFj3aOAm+WvQ30NhBrDxV5e5mxoIntrL2slWIrRsuzHMc
t9KOPCDCD2V8Eo9zSoBkHIY4lNXUe5UFVVIRnbrcot2SRiJYDE7vnv9HGai3Ge3C
+xkkw1+qs/bqZiLLPX4gIMihkY8USqL0oTtDSmyfWImLB92R/jLrCDiQPGT3Zrek
5T0Lb4Xx6SwpLV4wQ3hwIQRGIC4SBafiCTpP1bmM4r4J7hNvp/Z/0hzCDSdzwo8T
7YxbrRYi07xs0G/Z9d8TeUZRLINkFPU96RqcKTtatvvOiAUm0Kpyk5K/q1+7JpfM
Vvd0aVZlOPLNFqF2Wyk8sEvFL+PrM1uX+MtY21cAC2oBQWBfB90DkzSJ4q9gYl1i
bnXW/O1HavD1Ng1Dxmyh1h2qP2WRhoNZQZhE35RNqd0NVdzC2qRz8q+R2GmWUAYR
uL96feSLWJtw9ZvoKakcVVgJyo61Cphu/e8Sct+mzWtJnv6I14DW1vxG3LRNQqmc
3zkJPlhQPHd3mmva79LTklVjZxHotibNCbxxua/C65TA/8tK0viCUfEhGBTgMvbG
sKjPgEEsEKfncMakyNbty+3crfzCVUN/sY6ffaNas3o4PHCzyMa5vg8L4KVnbmYT
+CYoWXS8ZnGQ42hBHVlKeqHjL37GssyTH4jpVG3P0W8JpjDewHJUmww9LI1j3qcV
a1qRVIo62OoQ5V2BU9NbWSzNuwZvpsk6/1aGzi+FQFBTJ6yk6hnno3PbQP/tCqRj
p6StU0lMNgyho5NnU7jR0QtQIR+Z8Vk+7fJh+yHlM02zDTuYywPVEVCVT5Ug1ZcH
QGJl71qWsPwiuPQFAyRftKOyjWpW4vpkTShQ0Adku4RhP4I2Z7YMmoA3KqlIw513
JgPoexI0RDDLGAj0S+C2luhtSQS7l6S4gvXh958M3qU9sp6BDTqSqu1oMT0FbLNR
7vj2MRdfPLqXHLb4+lckllPT09DJ8tSQPQwF0M8ldCjz1sjzEFXjEMYDMGFiVHnb
Z4A7U1+R7G8OwJ4rKwvLKDCln+d1gGBw7V1ogZyJ5xU0RQLPLO8VRp+pcW9AfGJq
L2BCOzmS0ZgajDIORxb9vGuGQl8Xm9Ft5JFxVujZMF1Lg2NA+00K7bh3Wk/wpgnI
RXbzf7Xe/qkLFWFzmxse5AJOB1MNb06NCELneqU7AJtWNQg7QM8gcIu8kJY230RZ
tcoculYgitHuh2ErsXkpD00QflIyQEboK03RpjMpBTjw1YOuJHoAaeNJ9G2NxSSv
cicRKlswkPuvpTGNoSsFtUUCtuX9fL+92FxLtd0k56bDXjtpPZT8cCY1o8YBD0Le
+GZgOI7EVdvblyzNSQtUZ5v4ViJYx25JbVp9Oo7/8xOxnrlI/S9jdL0OxYyBPud1
SF51dAiWSr2KTOSoaDExJR8oUNtc7yoHIPbcKco8GvMMhrB8Hr701znhf3bfHGTa
/K+TX1M3p4eOPcJ3TT48BnudAsAizy0/Qs88k9n/+C25VSazR1b/gAgoIh/aHeRu
ngjsc4IyJoQyeDWP9GR6X9EIjOcGM2jcHVeuqeVb8KQkboQNO4JlN7xczRhbYbkL
Iu00c2x6JCt7Xl5ErthDhzPSuF0vecgt0ERa9BGNTAl0hdDPmH43u7rSptETAb6C
WuhpLJ242RakqFqj8osVdQzG2FuF/A5v9eTtTdLqrR+nX4WPfXEQ8TMRt9zDNFeU
NjmUEHaMlRQHnujDYwzd6hgH9jRlkukqLiJU2zXL0ED8fskgM8mvof5p38zSAxdl
BCThxHeMVfjcmW9i8xGYDHdBgLcIp7ImzjrS1hStjpfS+jwpQStNDFWit76OJU5e
FuvRGhXh7pcZ7ZDOR21ub5mKVsJ8oMQvNOqoaQmhfY/sFaAIJdsBkG/8XiD9Cq5h
FcFYt9yAjwhM92u95FYctbfqUpp46xqO7HNGATZV9btLdgJ/Tj0Z2ws8ggkgdBFH
/kkZguCv7rsDF0XpGo2kiy6A0v+HQ4/MJf8z0IufDaKo4fLARdHvJzZDegZ51ywk
FBZZc1AVn2UpcXBzp+wDHvjmn9g1VbxheQfVi+1kS7spG4k4RtltU+zVqX0zrZ7S
BACABb55lwzDfCcI6K6+1smW5nEmvdKw5Ayv2YaagJHB3Gt91dtUcwSlRhFYrNp6
TBaUYEqSd7oElLc4Kaa0TxuiuOWJ9KO7hU9ZAapWC2b4+PWUquqkbHLwNSqcxViS
KSeyibu1dPJEPaGhRHXqXmbpwqNfbmB7dIl/kqFTZOEotXYMpJ39/UgqsWTmjDgV
K4E+RAcu+lftfAwe27289PMckCc4WG894wiBWmyi3xwYlt29BRyDexVkBao6Jvmh
nvdeDSWpy3bRtCXYOj1zZRElVDcgjlajxChtNiKovDFiRzZV2zkJcORmqzQdmhT5
a9U99DINO/L5Bq+1BNEIFxf/X+5YVXXFo5TsO5vm/CWp8DBCBILIKRARRxFZBG5G
oEIzEgzACYYQC2PBx0FOEXVuNHpy6vFtgFKc1ocy/XZWPgJ0UT/8z5dKZC4tUx2i
kFypt7zS6M7yZCMIXPqYBUKHg2yLc6ADHFExdDqkzBbT21Sos6Pa+qZIaapyt5gT
qbC0PCXCVgcB+zOJOrXLZRStc9og7uKUGwiUjGeWLckabOiE6s+PNZmwV1cAaXwr
fMZBU0+0Q+5njYxr+dDz3ajbItQ/WAaINSiH/0PMzYCDmf9UJ1hsMYEGuKScbJc9
+4txv/bSMZyYQ7T7bO8WgVzlJXVralqKKxteMZMLnJN/JS+mmtGGGNe+PUcenB7j
U3lbKNR9xVQ52A+xsSQsgeDSZlNgVBkS1Q7fTXGZm9agYDrI3eZ2V8yO4dnhBHP1
n9iL0pjwMFkQZAZPH/g1ILZ1emekl9CH9C0zLjP1tpKj3AdhlRKJxVaUrj7ibiko
bZZj7KkwUUIyiV768KmLEiBHCnUI0Zo9Z5tCasBdmn4xrli/Te0uThuBsj0fRnQd
TkTjER24dIY4V6HHwJnuOFyj5qbLRlEYqLr4I+qN1zWUjqG/QrPgMbY6jKIBKsxO
0RKoMT/ek/h6KHVx1WRHdL2HEt1dHgcEvqeFeQqXwI9jpZxJ/YztFrRj5uHmyKzJ
94+Ihg8I/InZzBP69IZ3H9wWvtdY3kvYQiD9JXC4ATFxBp6c/8pam1ihHADtWSml
cxfEXfgzzzTYejTTVxIYzueiLgHFtl2LxndoXT26qKcxOla/RKTyboQhTss+6lSH
8YFHzITGzqhhWLYZ3CQ8rD/tIg+Vpw+AJaA4oCCRWtNOodHx1ZRusFTuCuTNzY9f
AGctWIEhJweMhoO1oUFdGl4rSIpIPWKHv0Be/OjkSOaLSM+WEDmLNNl6HWGH1GkF
EG0wJ3ESZwa14QQF4hcJj2bu/cOS+yp9lOmMvaPXWKcPfCojRlpWWlT9ePs7pLai
GcFX9VCCWBWq4EaI+smso8LN0502W1lfi/+wq7558LZP89JBQhjiRUtd6b5GGKTO
Inb278XniTRYJf6OykYe1+EqPLxI9KNz/TKVmspcA8RS4WAjkLJex8hANzKL8ym3
w/6x4y+9VL9w4K2C39pdBfr/KTg6oVFWs9q0/nXsQmWKJyUZHDhHW9hl9AZGlT+g
ub6qg6l2ZREi0UhXpQrPwhJAZz+gVE+7EMp8lRvNSbQViFYttnFyjPERILLijeXJ
L/DIesWjSF6SoL+E96uSWsGWW6ItJUG16EBqfJDU4eOjuy2KzSre0DqyY7X1tXbq
FzBejbVm1qp8T2vkeo/N+mOCxEcQhILm+RD431Pc/dosKZ0zfPIkxzvO2Q14FS5u
TiXW3mUPGChzBaba5TyoQVvJ318a9e4k8rhQq+Aa9gLl7T3zWH/c/UFJao8sU2dA
2KqJuJQVLhnY0g49qpGeTEtnbU1QeZY/ALEpyprHJJQBLrzIujMiMFNzIzj9IYGL
hphnOVytOkq5R2aCYuBKTOwaZXErMUDscK3QvnDmKQ9lsngZQHa6vH9VXVbQSKIc
FIFW1XiIdHsk3f+3UT1jitKYCtXQg/JYFKRkNU3aJsKXmyyGxmjmaPLKtUEAS/rD
U1XPntTM5e5edGTpfVS3yf9g8wtO3f5bk2PsvKkoekK2klkKDILk4Fnm4Qsm7ySZ
w1PWUBiieMDoPYNNegJ0AC3k4eXVFjwCYEgbEP1KGxAP4/Rcl3fHHOI5xcbcLNf9
1sD7wmfbHLcxVcsOaTxcN82bT2J1LVV53FGcS8AWldDhUIhvowfjjVwodWS0nLog
0OKOLF5WTwIQo1+464AdxY/iBQdSsztF4hzWBiSlrrlbLTEICdGl6rFi3OgJB2sD
L5kLCw4s4p9OS6LvOzMMToxKUPM/n3kHJW4ph+h6vss4ahYT1OhbE/ycS2u1sCLW
`protect end_protected