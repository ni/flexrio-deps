`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2016 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
dqtlaMM6dsCHKxM+hr1+dhP1rs+emWhb/HWA+N+JVD6CxmK0nwMK3bJAsA1jnWwh
xePd8TdlzsTVKbu2el2msFMY4Kob1TVxjbdUov8mQw5JZDDNG5D1CZevIFpK+axP
3MgY+baKaXpbfRbS6lXlCVxOjwmDtPqR9oolnDFuN+dTeG4MuhYpZJJur+bbAJqL
xVnigdeGU4fiRPu/8JW3/Mt3SdJsEeiSudHzcNYS3DLJUsS/gfq2C+pXnRgMHKjl
YsUCopgGptnb2gMi8o110lZglmS/tncBGoCKOOL4YqRES6daubsI/psDT7onIOu/
N24hTD9Au7WsNVjSk7ZYyVhPx0hkANgUkKPSJ7JewD3GJYE5Al2xtGWvak0bVgvb
Ostw/BKV0lTFYbmKQc9bw9ElCSB9VtUhXWe4f/tPcMm6uN6iYrltnKqifGby7Sy0
MLVWfi44enDDn1UNrrMgTjh+OpfrAFXMMrt75ML+7TV7dNlfrgtQNlWgZMCvdlgB
NIxeXWuKn8a5MoZcWXNsJKOu9bTdn4lHor+2p2KTHUwHt1dkttV5/5aGeOi0fZGR
XTrvgydLIh0lrveb4VjJh/Mo0Pdis7b0En0wdd4OqWh9JJZHEnJxw1B5DsOCNoB4
nyiZEMW/ARr27IyyRNyugEi96WOUHBsVuGE4S7Fl0dcH22WOR/Zjnov6hwSaOkaG
rhknpvIZIYB1k1OKxho5cg4gWMzvNZqBDiz4jJ6yFyA7lcgFqEhgCJQ0Vrf2qP2S
5WImHaP6HLXDZPUoftHMGNkqwDRoAYEUT2bQhCoAz+zm3Sbf6U8rLiqF76e82JVl
hV/f99T6/xpTnFZi03gABzzTkbHjtpokXJeOQfalJFwhoCX0A90pNZPk6N0SANkK
C/zPvQGy8rd8XDxJj9/HD1kQHtDf7x5vns1eredzwfC6KC37eYKg+YMlFLSF/tVL
X1jjno6Xx5691Lyn+illYJuQzXFHSvv350L3P/s3SisMhBWv/7dxa45AjPO7xztP
PJ9sPavFgJYi1dZPCPW3kjGRXeTmhdhQ/u4tMzbcukg2m02vkHehuz1d2gGHqSk9
rIQZFDmbutXAzhPgdf81b6jwLKuflxQiZlp2PI4qM3GRb/EBavL95nXmoBV0tw77
6mIYTqjF5RXBiLme9bGznmpjhWnSpr3KVwIGZJRoMxv/fWbYP12Ru0jgf3K5YTwR
1JYScw8Sexqow5old9JEdpx5cLcPWRBprwDz/rC+x6A4x/Kmn/tGkw/nzbx66Uln
v5IeR26tsV67QQf78H3DuzVS1BHyMZcsb3PxHp7x5jHebjS5flGfJ0+V3ITur3Ic
4sPNiukM5QF4l4Nf48mh14ITdnbuwwGqwYMMXz7t6YUzsmM9KL3XEkZT+fmFOCQ/
55+eSwOs95r4HbFwGS9eosZdSKe4EiJ1M4DdBdQBZMS4NB8Vs4Sb5tnZKSDzyw4w
gexveeV1rboiq2dSg9IwvESvvI8HxmylMRKqScYkBmJGgydNXoniCvsVxboTirCW
W5QLtxjm3YvmugIsITSIlaYi2/y5rtbcSYn1MG3uGLVxo0LmzgxeTthI6xFAFmra
Rzeovd1B4RYTf8ARy35HKEtinTJpvwxZc1Dd/BcuUtGg5NUlAKoHYFAe832tVFO7
QEmIiMldHmIkImGh1REoJrhZ7VcEHYooPTUe7QYu+DbGdxQmte1UKbtEQqW7S/G5
EOqzn5Gtkm7WWWRYo120mpQPBbMxnEWuZSqfwwNEEr2TDnAVcJN7ZVxK3GI+/0EH
0CAPNLjoBHBBl+2waPQ8BBDZ7Z2KQ/l2Wun1wELtQdd4yMFIIwhsGF1+8ZCGFuG+
FQ6GNOE68fHrxNQzZaIwnm9fTH+WUy0i4rwa9NzsHpuGO/Azf8riLkuleXaeLg6Q
5Vdu+wOTNWRJeY9b1hY/+RTcQAMdxztyFHqQmrTtiEM4byNoJ6lDiijE2ryjqU9c
pwFyOZCTj+84lo//BDkY+rc7MueFwePUeZ82m+woZYjZk+9he/PWBizGSXtW+ues
Ug5RUBAp0M+c8BN8gfFOsGiyINNnwjxNl07Qo40Axt0rCAC3W9ixL9qHtlFWR+kn
AuOV2C9rKg5HSSCm2kL8pKwNKUmQnJVRejmJznCCPlK6wXhV9Ijmt3Op6NwFzgNJ
O7x52vPMiuxeSTvHfkzt9zNIHCUhulwSW0Q8GCLv47nNb9+zvQaTYNCdo9jK0hSr
ZtkN838kU+LxPp34l6VUbui5zvPau8UNJqvONQMOUnJjsAOMEZiiy8E92DtvOKoY
xBiGwJvtrK6JjGzitcgydSb8bBeJv/30CRseOro+3LW3K34zYITCRcQsJir/isvR
9NvvpLXZZbgCIiLorNkZb8XODeecoqMfvPZDmNw+MB4sp9uScJ2CDxDKbsxQrW1Q
DF/gntUHHteJbXoWuloAYpPXbMdTQGrdzjmqkKOrh8CntINao91XqARj3T+mBvyG
RfRHZgwkzQWK33bOswg4WArKMoh/a22uAsG4t5plapQSpaexLc5DATwrjq8W9oEo
`protect end_protected