`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6848 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
hRRAlfE1xLfeNfywbrz10Bx7C8kdkvT0n0Ec2jbQj30MAxIBUS7W3iVxxEQvOGep
NtxUJS/9lf6+SfpXKJTc0rkOA02qKgJAR61JK8Wja/HCuKnBa7b4rgIAmlmDL6dQ
01YHOzWyinbNtCzysuLF+zwTOOjCUdYuJYlqRBGjnvJHvGXJtaVoUH+Qw+8k/hfB
uSjvs7RqE/rOj5j7jEhDSwtjD3bkEWlOVrtaMjizI//9ElgqetRybktormgRCJsH
1DOHLfnxmNeqkXJSK5W0GOVqau32vbET1jhAVKhniADxOZY/0lEFkXSVtFp3Rg7R
0Q6b9f3SsmDSAhuooUiW2QOSKhkdwUTqMmCRA99b6IAbPkrjD1xF57kMoKMxR9c6
/z1rGAKtiIQTauQ8djItKkaSH/f9SxpNhRkDEQgtLw90UOBXqErbfC3n8Wdub5+x
duofuP5xKQACyDyOebPIuPSZOFEDmhJ1pBYfmHPd3YCWWzHYCp6qNvpylp5nSfVE
ZXfSAHhkiSMEI7qX4Ex3sXeu70/FHeXVw1w6I3mOT+Q+yGGvywLiaKd4hqP1eUpD
KwIcDg09yoNaUNYs+ut/43bsyoKPqqHx2A+/rMBXje/InYR3zWd8Qu5iZ+jxyb8T
9ztJwZh6rQe1zxHNy5m57YqBkRRwVg2mbSRCq3ucR5dNvcNJbt49k2hQ5kzlOAns
JG+rjE8wUKyQRnM0QUCVD/l8H2HDLov/TTLGG3j3GiVUATXzcP+yQImJ+aYSl2BU
8eA4gQjr7H44Vs/j7ZrB1l8SYpkUPd87Vh9ITtk45miEdzq7P0P2eW2IUGkmV6mo
kSKvUKLQC/Lb7C0EENtnEX2IdVzFyjYn5s2fJ51U4lnhu9KwOyb5/3K6qIpR0Mb5
V0/izW1v9ipU4M6TeyY/E/P+c4g3yFpEvbciYqggQSRskPEXXyED6h7Nq78S1KXY
ZXzmkoJqWhrdLY/5vC+G0IhMBPQB1ZZodJqRYcBxPT30NnbbROL+IOtwzzc5tSIh
GgT642A6yeg14s8hs8Hqp25hPwLqg4RBaIezJnyJ+eKr0pGFjuF2ru65Y45u8kk/
OcqDkkQHzVGLmYXUjLUfM+h3h+dAY9+r3bEcSez4ItaQeCyDdMXwNdK4lSdHAWvx
Y1tfJ007zf+PJmGfCEPKRlJWlOaoWI+V7lQ+BUm4dMCCRxSF/hKMGglPIUht1SUi
QOKeApA/cFEXRWC3zFk/7bUWkna972bzD74MMW4VTCX374Rx2gKw3Y32dSG9ORh3
JIgWTxJtl2siU46jRmoV2rF3qVW6c9wM3iXRU/Xv4GPUVW0fyHDQcqKFD/KoGs77
oJNoxs/OQwuX6TW1MiNHTF4FSArFWUDywZf+V/EsodQ58i/936pCQ8mEexrQ+Cjb
wWa3VgDpsxzy7/dUede//MQZsNI0Qw9tXEMEO/27B6OQ3FzbafBhSIQYbOMqazne
nzXa0ufrpcSB2x8KtfYrK1rdbx8JWOHsdq3TwlmUGC2CYRG34nUw3FOmEEQVzpkA
2LJ5Gu6J/Kaf1+5u7gXc87+sgaqISJHHxsLl094nTitnYYb1wjFnZPuOz3g2ZYZ3
VrBBEraMecMKXZmeTgTtT5VPRYhjGZHIcbpMB7VJKBSQSty3tF1ZXR5dz0jSLmM6
LefDQBLq9p3okLcAFj7eqtYocb6N8KunWlwXY8MvRSlpnijDXmRLDNIoR+niMJ8g
1hqBPP4W3X+/OOiuTbrOrxryZID/EEXl15UgawGpcDvGXx6qrOr4SsNKoqenPbLz
XTghBoicXLzuvTaVfOtB6KOsH5/GIQUPB8Ss01XmMxfuxLmfEHO29cjOI6Fi36lc
MfBF9EY2wAEbhWGurZxMl6P2EFUH//kyYw2+78CxlgwAlSm8h+tG/5b0ry9J5QV4
wFj1JPnE5b7K+jbWCIWMXjix44yxQaOssG4jPSH3MMXdgYwRxRX/zmt5JOuc9Xoi
PS78mkqQQEmqXQHZTDMLvE2R8/8YcnCkWm3BrnnkombLQyXzaaixVIdAsYFarUf6
PwDm7oFtHRKnrOn6KvlhABTNaesS3QRU4RkXWXiGnu6RqWZVbqhyDx2BFv9yZM6p
wwgmDRnIEf45URVRzZUd8vWB3V5cbOkdRQCxwUny5ZNIHHdZFf6qHTNCF9Os1kEA
VwIq1G1A4gTgrvN7383NMy8Lq2OHGa/6bQis/lUSEGSqb+lIqD53bp4o3ftTqJFf
DG543U+4GMFS9TKcUmZevqgdzw7ZPjzenchaT/GAFzMbCBCeuoUXAHIjS+RHfP20
/lFOeMs1yDqY8m8zPsbSvW5TKqgmAofnpd5cBtXd7H4HCNkQRUTyrYjQc8ovJo75
nX2Q2FNSk37OWuRaual0BTqR5dR8xmwc7dvVFcaQ8YsWzzUtQShO20Bg7P/TGJPz
6cHfafFm1SR21jFG9HJtGWve4ljFKJBYmZs0XDaYmMspAy80jFYe7EyHlFz89CUC
5RZ6qE67hbaF/YKHFvvUNa7mbwN27Id+0FBUVtA46Numz0mwRU4ue1m8kyBddpyI
TQ/7zk1h8cdzlAuVJwPz0uKMY8vjViEPSqieOl3s6IZ2BijDhQ03Uk3B0+kkmfwd
V0ciVbLkeGpN1/fw1K1i5v0Pqbr/pXcVXI3LyV78yrNXqvntjQjKYZDRhp1SlNBo
QzPXTryj3kC/3UQowhO+7IksqPmmRu+lm2e7SfPHIj4cGB16QUA7pKtNz7JMhJcy
i7jE1r7eTFSBBlvv4753lkTl2qws2MWeEv4CkjxpPKDHGq8ZcxRHXZM3qhrx+FJq
abDVLSvL8rQ0sW3rRUW3Rm1E9IiTjr4veKLAs0s5vYBDzosANoZ3UFrpcULgOAL8
kV76CbrpqDTR/EmAsSu6mlh5eACLN42fYk//e0kK/2R77Wgdfg0QuMhGbAj6VUuF
T22AO8Ly5cW6hswV1KQtROsdG11HO8nMWYQOg+xpgY7LKacqXvb+WyHHkpR/bt5G
/BrBrJ5MH7goP2kgGyHwm2usohxRVtAV2cj9V1Ye3IXi1PxNZzppADSZtNJ+sXFh
ZEg9wSqxnWyeTdce4lC185jX1Ux2hV6ciBMLaEhcPD5ic7YV4eMFCMA+4WkYAVgn
W1IaidZ7q2c9zaKF3Qn0+0lPO/1/1bJDSDENIpubmvM8xgzxfLVetfOcyVbzTVQu
BbQIPI4U7Vg/X+iuRK3npi2s0YO55khhxjlaMrA/WOQ7uhqccDT1Zc6o574qsONz
dgmgAsCkfZGAQPl4uPbJp1p3IK96ZGayCEqJt/A9Wg9Gg45LL8bVc5cRhl15reWC
+6kMSnnkJ9tzyXvqu4gDjSIdvzl4MsOACre7FxBy3LpES1qaCmZYpie+qUwR6OgD
2/QOQbzfHXjjyZsq5Z/4a21jrMoOFS+3OCQhTkcSbnoA1d2odiF/PFOQY300VWHM
4YQ7ZFmPIHlXyZw8CEGCMBIYcbaJYkzVnkR/DsHIoI9CUUd3yebOnNY8K/j6x4ZI
5xucc4WgKV/e8rSHxWmsmqIzryHdElhWuBWmN5hUVcxl1EL8Wy5Ffno/TI8WLTMI
eP6fzs4NGm0Vy9ouJLV2XTF0kTal6VT9IABKheNAW3eJ2mxMfAISWloIoucu+jYX
EImnoK3CH+QW/DoemF3Wo0FaIMPMlc4UYa+mei3BD6d7gRa2BJZzuDzCAYvYNvXb
wp5YHiNE096Du88r3SiVrXE5mTK8+s7Pq2NhFkxqw5sBeWev6/4ApOmqdQHvOGRP
AHIw+nB3vmqly06Xlx2Cqjk1L2kKqZYbEYf1VU8iE5bxelzfzx/whlgGL3iVOyel
/9PKNsGFo0eCImlcyQqF3JlRUIvSPy+zXcPmRWqSaOOr/VSDz0qbGa713/zHF2XW
IW3FTPUDYTptXdwca7j7OdfjVyhFsqU4RPIl9rGoUAJYhEJZc3Hck44vG3eIN+Ib
xwnOWj981vuLgncKIf/C1O/TCJZYiAkqsZoiecnTJSvDeH0PZywdjOCtuvjYf+Iu
GUBya6h952ki5NzLVnvdbU/qDNjbon5HUxm/8Foy5KI5JnsQk0OIX2MxKqHXnQMO
tyl3akFBDNt3IQsw38wX4bxnvZCBUlpJqIDIyoLCMqP5KbKkjYBa6kK0H9yL6xsb
d/9TwR21p3QdRuSbQKCJcy4HXNYFcUfT39zBrmzqPIeBQu329oGEzb56+rP5BPUf
JgSTYSfzpgG1qhFoMeSFbAwK4Bdp3kwrWEWnHIhGD0KmIb1YyzNNsS4UgYztWD3+
Rfp2dhhQrl6B03Ns5T0CaxGvv/eHOwwBGgCpCTwldWJusWrWG77iQfQwoDXtVU0R
w7r527Hzg3e2d5tAACcHxQBN5bRhcUhnzpgaNfjJgNgXw2Vk/b+u62qUgqMIXAab
MmS48X+7x78ddUsmuA1Z0cHZ3r7XUJiFrWKaPEF8S8dabkCdvG0QQtS6aEOWUpoH
PUflip4bciTCBzeUIFx8eZe2sOMYu7c0kIItnGYEw0Jc+EehrrkDGTxQzp/Afp7L
FDJ0wUlEoeSs01g7Tg3HZE4nEuc+gD6nyJfLh2t1a0W8i+ALB+PY0bqfnLQAp9h+
RcQK8V6PzE7s/xFvpoEHsHvzoZW6m8oCt5vHmLGjhY0Av+FpRZGq2qcQO/zu08ek
ycA+SniMo+NxeBZo4fMnvcmnF5LOFJzpV3/tM8gfCTqMFYCJCYEnUt4ShmOMn2l4
Qic1FGo5Etf8RRpq9Mh+2nUkTaHkvhR8GJjnHtRAprIvHYL4ws2bIoON8P7bB08C
B4aCY4Rf+Gj+4N8z7vcnfaxqBvAuyxcDz9r5cYSzZIN2m/qvjEiPWUYN7kY0QQUl
UQa/Oh8nJLJFZ30YWKUHVfcBn+MQqruLlDonxoiJmkaQHIhhwFfly4WhrIW7nwqp
N1/3Y8iifUfA4IG0nxPSKtf4ZV+39v86eWu4UJSxt9DNMH7PwFS0Z4aoITOgP0l+
tOdm+MLwwFWx9X16fBpQlnk+trAporPglYf1eegq7tw8zd57RBb+C/lDiIZZS8zs
L3CpJLQ5L8jyohx27JDD2aEk1wmcpzcvVq1jygp1szkrzCHBsbxA4X8IPTecJoc+
lzpY93w8fAvZFcUJFHkUgUPwBrRXxE+c4L9KE9opQQ84Q5Y5pa7o6TZoot5J2sRv
vvT0E+CdJXOO2wuAwn9QB8dwoTRf7eDcfQ9QrJY+gc9PChyk0DNey1Wu4eRn03yv
NhL9v0IG5BqxSQbSCrX0JJCQQgcPtROMuLfQDzg2AZon2FK1WjO+2BaIul+oz7NR
diAQwhdsVHdCOjBAQGkKV7gSgOiDAcTrnAUUC0UirW+vLMfgz7iUvwUwXs7IcbP/
3SvWNOr3US0zUbZOz9upXNovXuuHCS6N9s5pLA5pJlRiMiWzzdPil4tAHu0p/GWp
Cieeq/megnZHW7yvjIlPwWQ4INrUPj/Ngcz4+zi7wLpzx3cxjzrZH0YqfZWdeTRV
AtSMrqtV95tDCHL6UXxGWGS2IO6T2Wc1OogBpFdFCxAy6U++3Aead8xGKARNt6oX
Ui/MsfwtHYb5QjU8YMIBalRGlZ9a/oeHmgkjdOE1G30+KLRQ6AHMjxBCC0Y2Pgt7
Jwn89pi5IMs3S3cz7YHa6x2qBfGx5ivLKS9Z1duP9K6tnGN3wn7vmfVyP9yXGx7j
jD2vqb6eiuUBYgujhFjq0FeGOtWcrmPWQLx3moNaos6FNlIA+W+xwXXPNRmLM7ce
kXY+rRXsosIGMPn9bNP8fVAeR4nvcm+i5UJzeMqrW5iQ/K40ZyaUqByT71G3nnLz
q37JdCQ7QryR4fDImzM5zlERec7ky4lZ/qxaFIOUoycbjBZ3lRyaXmRJVj/Yp+GM
mwDzc0I8WFOYHTDzlLhgjOiNrTMKkkNY+hQ22Tqwm4Z5i2pzWOy/nC80SA4NybzW
tYy/vBq1nAfJAd1SI20dEg+ErfoYfW9bXDpMPfTyglzdn1sJYPVeQSVPkBGLN8Y0
c/GixKMw50wXdQkLcNtw2VrZWV3r3K3XDpa8AocQmCi6da9Ga97ME+kL28EoOdfe
w0uQf5bM3WXqZ2bzrfNw3VqI1zKJG0/VukhMu6PRdHJck89Zuv/yolo6p6f3uKh2
fxLJMYETyav83ih5NxF36pZmLYJInjOyWJutYG0JD1zIBKEst8kgRIxKA8MuAILB
t0QfmyVjTN7dWzT3MsP/oxIzF+V5iBREmaeGD9UB4eT4tntyrWKYFaNRHV7zwSKB
4kLQEKS3xygwqdy9CdlqQqviuYs0/xIBYQVYd5muOeTtQxdz+XY92OYjpUEXcqmT
oyKSmjwa38YsCa2iAw9Mw2h8Ak9onbTzXYrbliTjOhyUCcBU+rYxCuLao8Uy66M1
WTFtaXisskioGVQBV9l3Iz/SRk6/OjlZvVK5LvzG6LYuDjoAcS78voU6kLOpVFqy
elCNym/tTp1WEhyKEKU2ML7E59OaBoZK+YPYBMkXP4ATpSJl0YgFFrEcz0956dPU
+vMu9A1WAx+JFUtWsejW20A7thzsnfTBFAurO+qQWH0hj9wV84DIYUtDhJkQoTU2
9J7kv0S2tVzxDTSo3Pe6knbAowLNVjBUKuJJR/nrt3ghdfnG0OWG2BPSxDUWh6WP
rwmw6n9Mi2M5RzKIsDpw2whMSfAtEk8tV8otwGXu7nv9KgAlOzwcE+mOFt2+Cn9i
VI6kMeC/4HSYP2gJly6sl2Dd3pmkX8XFAWI+IceFCgdTXTU/jrFntrIyk223HYMw
ITzn4sA1zgGRoUAOiM6iYU1oWG5D0YQUJhLrY71+BHSTzc87CkDP9IImaTsWpwXS
dfZT3XziHx9EoqFivg8POwGoigeELPcf9zFF1mKgjEOcfBbJQMZQSTXaophZ3M26
VbWJjnPWpa3jbcSgilVhocow6owu2R/I/9L+RlITToocHi/SZc1eZAZ60wMOFMLk
G44B55CtMADiUJFUv7gDBhiAE03MydJFnfv6f2bynmoQ57v9syW/OVUBOZB77szI
J0AiiWE8yrLKt9Ju5iYY2jC5jPugG+JjlxFBT3SKfan+zqA6Pv1kU40UwypK/+s4
9udGDYky3a9616tDU/sPg1D0a/Vujb9CRllq+lueghYFocZP6DpXps9aqDT2ZKlq
LEz6lwymL6Ng83eU5ce13snX5WEXRqx6WRmhCpCP7mdddgRm0YHiB1ItqfVIaUs2
SLhbBayZDgB1cQZUqrXvRTMU4krlkVHDFwXt+PSjI2piJoES/uae4YjouAQCYSQp
nQj6VP+dEQTEFaRm+ApCcSQxP8K49NRZOOcNrnryt5CvfQJbT8Ywr1KLnpqqnXmz
7Vy8jo0VKh08IreAlGi4oIIUukX46mgggY5jkAuJsuc+JgFNh/1royRGyaxYPpfY
fLU8FQwhQ/g+TYx9I/vWu3n2+kRF98l5XBSJTiNov+u5e935NCruIiAT+amExoX2
jq1b9UR3X2tb0Ar4Bs6MuZq8wyjCb4iESU6Nepbmd1kV4ayslfUzuvJD8Zk7Gjc7
qrKUbWOF9R7I/rgTtF4PO9tH6HEpBiONP89y56bhBkY5G09maNbC4DS+/2yZNa6P
hWdSuvr2WwGG0B1BxMzi10PkuaSKdXQ8tf6ADJz5Guruk/WAJCTTmxS6Q8mAdONL
UfL4oQKy84Kpr5gRt95xe/gvDwQfKJxSWxsb0yq1bULEyl7WHjF8VM7pwOI3ZKgq
5g8M4oSKBTNyqP8A0G+K0038nkJh0msraRiUBdnfNwH22VMNHCo63I6ey35fHnWV
TWTD62NN/B4InoDCO10qnyKrIXHPJCosRbW6ZbpzOmrubJN39Uv/283AZFEP3fHj
uCZzP2ddMlHH24JEMTYlu31IuP95TQjTJndq8y6I3dwX5LS3Cx/tYT6fk4otM0i4
ARSuQCRT0s4wUIMlrmgN0C8Cpz/Fetml6ahD13ZF/I/VGYb/bUEB4I4TfuCyQ+W6
56tTkY+2XQ+4Uz+i5CTYAWpT2nYWZ9Mzx6raBugtYn28glYuZ8kqdcgdkpY2OTch
/zHoMdISNll17j87gwkU3yT2lgHfS+a1XNxgfVlz2se0PjZ1VJGq6OYZ6noswQ2Q
zwaqiKNLTU3aA6tXvifrajUYGCarAsqF47cVlVy6WVfxgq6R5ayjURZyunM5Wwd2
eCtsT8qNITVJLy+FNRbaq7y/6z6KQMfIwKSC0hwwvKRR+OVSByVUooXjzZUzBpXn
f8dFcuSHDXhwxt32SPVI7e9kv2DdJayVmlq2I+XC1VTDXZ8E2BQFFC2pT74/7dsI
g7HFGk+na6lW1iaghPCLuCQG6cjBcgpud9kM9dtTbmg/NIR1OjQOQA55xXqVn7H0
tW8J03h6jjGC0hQdYr4PPlcHDUTFAKfrv1AxD1xzSwXA9OV9cNzM7Be3O2woVNnR
7WYVcQotMk3tQYB2U0i4tSTs2p2zvvp46v3rxMtTr2mYgQbUzeFlfZXPmQEJgFSF
B1I5dN/cyV+TIQBoX4tkQ1wI27t1bfAqHZRRG92mq2D5OP1YNa4RNYOW8MDm4Ccd
aAre1EXrrEbSthqkA0FmjXtNMiNDItvQI6yykrIKq2tgayK43CtdO6Nv3BkL3pzR
e11uSlmLSHJ7Q1lMNNfN0QNLS9Eg5dHt0vUIGknvPBoX9JbBrNePz6ARfwrJEGVc
bhXFrMJ5bSLhwMDlnpUtzSp7xtJgDupzsA38Tgh98c/HRg4NM+MWyrME14a7dX6r
eCBIhzQlq4quIUyNkPev/U5WG9RNgEmg1zaJ2LZY/cBCB/HEIU56bk+85FKB2Yz4
AVjQTlTldOB9S/dQcUyOy02zQyFmge1pGTp0yWioVQL3WV3KkyaUpLlR3tYVfitI
/hCJeiYEjJRfrgcDfqKnReqnGGO6P+mC2b9m6tLn7oZ8iKlC0sMclvntl1NbwG69
pRzJQAJlwRfECGechBKWC9TnG2Cb0bg0u0ZuwBglGo0=
`protect end_protected