`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10080 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15np486+GJ6igjQvaUGiACBe
DPRiAto9cuyEin253BXF895AXpnZeuqN9YyVNl2kNbbZNQOeA5Qz52LJEFKc9yQ1
hgHliEz0YROnmvFofvUgcb5CpPl1tBKp4R4l3NqedZq6gDGFAEzp3R6hhWYbghOG
Et+u9BDeBHgjVNTsWFZk2B4W4NjmiQpEJSjw1DFotx9sjD+ZLA+U6bVJ7SZbOrEB
nOCy76pXYFV6DeqgYNaCjWw9tjVjGnFudPLhRf/s+6TaN2NaUiGxImkM2mzC3jxO
D/4+QhcB9lISA6iKXPRwX7lKO0UsL7xIRne6sJoQUZueFa0GaLjOSEzTu/uLKtvB
Mingxqqc1RVi/M4bR0bLPSFduNUpYzY7OTUpbxIYz3SiyjE4OOtRxjTfCA2AA++s
ATA1XmRuPNMdzh1Y8TnYqYPa+nM8XXx6cllW0aZ6n5YY2TbFdp9dYa0U09MSuANu
ngXm9Yn03Cas0Nqf4hfzX5cX5cup5wsDHoobQLo0KPPtqqEonTERdw9BjoXyH1wa
jrn0NKrBXFmBUHplzJ0urFBGAB3MVIpp0XMVrChXaz9XxjeI0I0WW6C/WN+7Oc9+
BLmp09y/uGMlxp1asEI4yQnOPeSOz2YkIhQbCpJWDZyRb2vnPOGCzuPvgncjt0kL
WLl4086egJm0VtyZHCLdxsXO4KX6PmUxWCcI7QJYW6BI7jHL/R9E4yV9z60Vtt5K
fAYBONUuN6aYki59V2i1yZePOnkmh2oU7PCtjEvBUKRtkyw9KN38Ry8VUnLrtKEb
fQLs3S/BH36wfolV4Hfn6GDwVNOB3d4V0VlWaBUr76xqoh7VEzZ21uZvtq/N/Fxq
F6VMvsTe3FEHs1PiX65ayRz0nkpPWmfVngAslbasPE0ra3dzFAMIYiHza5faLXqU
nGasmx/nhN75Yghs/+2E56do4hxyVjrLBpR3MVaA5+9qfbQDpoaA4F48gCgkyIj1
rrxjQNI2jE+pAsVacERPcA89lLlEBAtdZ8deG7Kv/+tRQM7zvwPuS+tTTrGAn6fG
QndnVI9ODSvDnTxxw99RvA0AY9sADa1WYX7Wzpy8xswqosyEZ0lnRRDNklKmOJFC
BAKxQPt/lKEqqjgrQD7nNCLDQl6rghrgMvT/CDQyO4WtSMGdi2bAdAxeMOKaVl6B
cwCFTgD7ObvBNkXv0+roZWHd0mqHFbPzT2nY5C5DUmp7iJnmvvHgHbPetTloVl8M
uOfCfoQxPZR9CQnJzlLESMl8+VO7Kr9cL26vVNpTlgXsVdO8FdwQDdASZMh4FoDu
5P6e6/9860rzf0MxX21GRMPe8q3hBAV3GFrM9FTOWEyw6cxkQGcMkDMTWLAIijH9
NKqls/mmBtaaLDUJha+2tRlOe40KY9Z34/znOVY/3N4l/O4Ts/KBV96HlawsEWb+
iItLQ2ZobnXbCgdYIlWdbhDszfwDr6h9OrM/MxRuGQySUzfZJBbp3JZN5dLiV08x
klaPrTPofgHF4GOEU5INA4Ewf1E+aKsBPHk4+/7vIPGILfbzIEGf2agyL1Un06UI
56N2Vo2ZIo+IT3vrBggkSDtdarPfLmmRXorUNnUvBXuACT2ZEA2DkGaYFrVZFyAa
xSXDwYfN7e9a2GsSZ5h5mAHD3W7AXa3FmposGU/K4n+Y7UZDio/4fmgvlOT4GodX
+Fp/pOe9xc7fRFP1yVE8lJVcgavPfXB6hPiNDQpXeusf/ke0onwHpFlYOmchsF/V
2SKfWo9RdXMY5wlyy3IN4P+Bw2cRt8BLrWMX4MvW5CPhYVru+bVSmJ1PQsp9JVcr
wJnq1aF8CZtMI9Dio5nKDY2JhHySap+0ftuC4Ae9FI7D97n2flkstrLYqBSwLScb
pqkjieIf6HDvXwSulN0RVlkF0rnWAI1ZLmHc954NLIBZHl4PcsQwK4eyTLcWA+vp
YP54DENO5U+56tOM+xRkejaNIjIjFIeodQVbNyTg/Q0Sd1nGhG55qymEtIzpGNWV
BA9Kr+GgRiU6nI4jOZ/jqKtbKqkxXaBafYSd09voxwcXSRR7R+q636BBIGwteSHN
gg8/jvB+0iVbMoekYiH6pt3hb2uIMe0Ccn8rWQUuYumMNEpUBAwwDWHVScFBmQ+L
h71JPuvqwenqUnCUjbGXid0QPmbSQ/hu5rBfkD+m1eI5J6cfI3bOYXo7O2VaSv9z
OwRvIeCXx62EpvIU+QIDO+endEp9mKvFRGfGB80agtHkoJrrvYLFcsfle71ILOUr
P46fUPA+NkdUfLRRX56DhQ8X++CEBzu2mkJSX0CWpeLsaDWU4DBfd4Dq01jB4RQ5
lQHweXiCZ5tVLHs17FIXOM7xy4sDkXSuQQC6PcgC6vwNNWicwXTIge1Pv8/iXyJE
D3EfeVFMVAXxfjMf07lEFvgtDoJbYkrCpRjtFUTPxYJLagH3fY7f4B8pTtT9oPhs
/hmd8JPj72XXJ3WXfaW/Aq6cznJnucHZpabc+LQ+xMM8uC623RFyCntDtzijD5XE
42Uuv4JSPPQvsuXJrzalJCbPNm9Iofw9jqIz7ymrh5KS3oZuQ4SjJ3rI0t9Rd8ar
wFUuYq8vtrMArKDYFYWZBkGq5UKB8p2wB2+8e1qsx8CnycUrspPSiwsLkA969ciE
WX7u7xBFaNGSo2Tmq5EfHDeEc7jMFclCkRIuFxcurZ73vrVtih+/Fe4pdIry+rRk
VwDr3/VrFRLEF21HLWeqCc+goSULCwWq5CtxKNLDVdm7sJK3er8yucF/hjgb/3/d
BcNGxps709werm7WfG29+6wt0VKqVaudMPGBYNFy94e8IUivqBT5cZKLQ8wzjuGj
+Dk7bXvkhXPTphY9/Zjom3KZ0/v7YWFwL0nzxw9j0a7419RSk/Y4vV4aU1h1P2IE
DwQn5LHGVIgp/K2Se9OoUR3lW1mNF8/Fnoim02IxEG4wCQIKtCVx9HfoSHyTmDpo
KDm4wiXgRoXgts+gzx9SpBrmhX3CjP8O4HKY8b8RumM41mxW1PdIIO9bzrnntQpj
lz/ynbf11X4fmgkBv+gCNxnXRZ27dC1B5GxAOAsjD0VdseRtiKbtxVMafM2BdCD4
Spmbuj/bp/XBd4NnO4JbIz51lU4WaNTQIH/79EhPCatuGagO18AMi6PwOxLaNu8m
BYJ4kJUUwGIrKgVPPU9ZwtEVsdy11NqNW5kGryfAzrXvA09nM7K0nRdbljyPBsFn
3pXVPiAUDGf2FIDsM0VChZMYahJulA6e2DCN4rF0H0CuOV1m+iCDR9RpQqiHaJ+j
C6q1HmKZ6xOebVT7GUnLX+QoEQyMsEglqkWrdZG4EoEDWDnEiS9Gs1x+KrPBkJQa
Gui+7bJjuPZoMygjp/f+s6Um4x+UPRCAh6EqkgmZIY+iIsFvUZn3BnOdzgSTl+Su
tAPpojsyzbQNLNJxpred0WmgRB/uZXJ/z0EZkPYPkJk1P3/fIt8kWgfc7hENs8b0
/ppw++tVu4mWP9WaKyM4MvIA6ApOx+cxJa2HQg/3AMp2ATKraaeJL4lgJvqUuST2
HRZZ09qJwqgnrp1VmHWTezTraChPEhIQYgq5L1O2/GWoyOXajgsD9BQa24mh7KSt
Jca1iD4Vf5rQ+UK7N7+9YFyOodVIDQd6UUK4Y+WE3fpPWSH9PQ77MGbkV3XsGYhl
i5/92HXEa6I+CNLejV2JouM5v2VZpGYEfvKvqyC2HYZ0c2BmjNdH286CalOK5Iq2
w4r+UoWy6AAzjTPOoBxdEOoBS3EQQrw8nSQKFKxdJEI2y0F0VLV4yt681TLFCnFi
EFHTGHWhT+40OMegOzq2ykrS1L2oiuGPGmCLrgf9xFbY2fgm8P3LOVmY2CtBCiaj
51cTcCDmJkhP4v0Vw0lfypSoYtNbuoTMKuUYNvHZBtEn4n0AvTkwwfH6ExkrFm7c
bIWLm9Y27QYqW+vU+xqAb9bR4/54ptnfpiIwrfDAxTc+2NMkIsR2SfgR4odkCHP1
Hfm69wEClayMKgUiLMi/+6q2dO1zM8p642hvdMprcMude5SejmRZ1+Gd585i5UdI
nLO/IXfQY7F6ArcvjalwSQE8P51kFCWNkqDws83eSWdO/Wv+5VgB1nhL1UAel2M9
LqJ4AO130q0F3f7si8I3pUfT/JGU4YgLSpsd7m9J4WMQks3aJJY8QD3R9+qdgFF6
0SeT7VGhwrlxzlJla4JMlAA5m9K0uwrP9hMM3dP4iLp36G/V00EgCL1XeDqFlPws
ciYaZSJLv6HevvEak4g+Vmv8YLzs+r1b7R/Z4nEND8BsSYArZ/ZMsoyY9SX5a1Ib
RDh706faBbLUukrfzix1epNX2W7z6c2dxq2Or7hT3NHZspvx5kMKPFjIlP0YO6Jv
Le7uzOiL+pSl9P2fpDza45iXqxfsIgZvzRIiiXiHAyObjYe7YymAZkaS3ONUUtNs
fpsGXDJNC7aUGxQ2HlFsV9SVMYVjFw8JO3WeBLQhOckNOz0yhKvEN97O8bFgT52U
thR7Mh+89492eGim3vSHaL07Z05+RdSE7O1kx6j1etDvOrRqpyFD3GzIqTjIMfCu
GA9DzE2BhywxKot3GbGbw1dGNQdlEAGP0SPcALZjUoBiSfbNBIwsF6Upw41VC6Do
yMSNBz7An6DnmjisrxeEsy+yABEC8KBTdURlJjUwcB2CGOUcnP70WiM0leViQyS7
clP6amVxvTQZ9JVDO9f67ZI4AqcMpmA0OruzzStQZZdI+04C8CVfckazGivBJ5EF
mWnBGF8ycLNjYtx0Xa1Mg/yhKIK+gdagbIr2Hv05dwwUixTUDy6udBWfprqUhusf
MKIr066b3NZQzjHUugr94G47wcw4W9TjRg28E9Aq1D7RkjKWz81v9z9+Zv1Z+hTz
gVdz0rBBCkS+h2M/sembYeQNMr6CqdhmrISSdMiqaIzhEKQsJ678y9RsoF5UJHQH
KhV6fOD79T/kJXYsc2BxgDraqT5ldRCyWMU27hzGpnIY67ggsGuaFsQTEoKSCfh1
e3zdz+iUa/G2SOD1TsIcejYiFyGSJ6UcGMuRoWnSwxqmFQ0tqHLaMphvhKhAgA3y
uZoAdbUqYLXpb/dsMOWzfV38qy4ezE37nouVcoOYDsxdnW0WY5+FozO+q4UKMQsX
9q+twWoZS5Chzh5uQ9O8RCLInlhP5UDivXdQtI7cqGpaDwv3qhfONzedt7HXkN/M
KdFBtd5cEx56Heufp0kW+D/w8DYCH8USXK/bdXJ/GmUyIj9rusoRBIswKv5zbWEb
vUzPzdt4xhEhOkFp6DCd5xKAyhsbx8IEyA5NkimsN9TykbSu5bd+2S+Yt3lw4lYx
dfOnF39xfQj/jyO5WqMtlxqmJorpZKwIrLGFQw/20nBF0//642U7wJego67sr1Hf
dmdaAMxfSe3VpoX//HiQEyW3PpWd6cEgIFMdfJXN/UljGwYEB2lksmrB8E6JjNmL
4efAimgj7tOb9PyyeDYECwqsFmA4qxZoVrddYa4cDTWt6B7TRTjJqZHV8IUIpU5U
8g/1Pw/pf+x58Jpj7rggtvgZHVcGEkQ2nCWQWMlyep2m0spaicnNjMFvgnF3tYqf
u+5VMtkx/t2M/ScvSum/qPtXv72u7F3IS6xZSWtdeVWmJbxqUAYTzYvL4nPHIH6p
LKC372xeT2Da1R9Ua1ZNEf5XgVPmfk0vYfcdOcFbeWvaXYiJ5B8V2WIhbLP+Hgbk
PpAIGcGHOXX4U5KpdfcMvvXg3+LfwhqCZWEcu6ClWflDFXkw0EoYPiSq8dwQOHY9
KOceJtnt9p/wRXShRsyY5gOCrgiD+pIZ3mFrhptA7ZxGzR2ZPh4kx2QpWDyDN+4Q
EjGrjQ4hgADtHFZPUdenzOqy0Xiyp7dYrWiYOIpbZWx8C2FqPN9dNZoZIoylzKYM
lvGrAdDsSWjKXBaC02VagkhLmQozNNuUAInSKSibDxlrFfZNmkUabBb/wXEx7ibk
Qp5URxwbr46/DH0OIgpTr4GP9X9UO5nH15jSkK/DGJtE7esYyeYyWdMFQwVa4O27
8OS1q5ExM0QkCUGdgGiYIFZlAwz859LqTMnvQH/rIWMGiZOFddNx06mUQ0cTresa
LwuO/f2NGbfnPHwHzNk0LFNU3DcfK4x68Y6qoTxN4vgdEUcslbGTywFY/kJVhTU5
NRHmfvIEQkc1MQ17SqZ0fe8f6nZiiPuBRMNH2UKpx+EICwcSmOFLEkcJtf/lJIh2
MUUOrLlTO2/S2Y+bnmqOwv5pUj0bJ+MHcBBZeeTAHuBeLz0ZzqVbVuk549Ww72kT
If82o0/eJX3h84G8x3jr/KQ7LxhmEikGK4ZHgcjoU+mTk4eZxarpk8f2xSWMkYYo
ucfpUOiFT38oAsl9SJP7UHc4++i7/EuWzQ/ORs826P9QC9mXA6qyCylcHhJk7Fsa
sc0VDQG7JXEiG1ZFRDQvrI0BY+0Za3DTAVSKP5qh1YAr5xBCWXNBNSQluR+EFnH1
bM2o9x0qqNvzJOH9Mtql1AjwJyWt4heENqC+m4DUZ0y4ksjmde2LKt/nnzUgYReu
ME+OOwYFQD6EZ60qvTkz+tmuF20hE49SLM0D/ofIQrDyDi/m+s2IJo1AgPnL2k3p
y/W4Tm9WakTQukbRMRKYjaaccW671+/MD6REgHk9ogLh5Taj2I4RzNSRRm7IM8qh
mmgqyISiDnnahNuVkNynpbp1wub3NH86AqvpElShQVchPUCUFuuCLbKk364YFP3o
JA4e52/5M2e28lg/g0z9ejKfV2KEicZDLFfYJIU6sPtPO1bnR9AGMifAktasKcnK
0endmh1ChCOhkAunLYev7pEkocVxdu/kJcpQDDkBXG8N7WNG/bqzv4FLs+UB4T15
hKao5Bz4kGGXlqifqq+7TbqvKHMJcZNB8/RQ3h5Zzc/Azq971GNe+bcVjmXwHI5V
rtjKsVwpc/el5ccT+dV90dz2dbwvU1mit63CFxdWDK8ll5JLRL3Qc9xwH4dfTN/E
n0Aeot+55KEe3K2n9z/XexF3I72x9GUnyGpQorX06GDuPzRsXj86GcTwZ0cgeR0T
JES95ew4SbuXdgmkJrIPzjxnhNq+Fc0E44M7vrFfEvb2PJlWW6Gpr+RvN1gaDq9U
a2UKtNXuvmR6NZEU9Sfo5RbT4ciVvwVQHcRtiBm0LSgBtU2o6YOMgcoPaFrxRj8S
50+vNRvDNlzC7hsOIdgIsS3ipx8Ncf5eCNaLXl7zIUnNLcX69rYSVjL599VPtujM
ivw5IcL5UkNIhUb/6DqshDAa1/Q54p7AxU0k6guXhPLdFR7ghgYvN+NaSmkekx5u
AdVqiyET92AXNSU2NmVfG1dmJODde5Uc8GDtFR+J+MJHeGjwZla/vtv6i7GD5h4+
1vEiPj/tKs+2OIDwScbAdaUaTjDJrebPE9P7PpWNpfBlaro2ezKkPbrypBT6zCg3
e/vm8NgZhKf1UWj3VYvo8/bSk2FhlM0UduS53V8wCjH6j4gDSK5DUK20hlH+2z5o
95h687WB2mskowVhHPY3nieq490wRqXm6KbxqO+I7Il2VCdzGeAbuOYuVwrUWBIb
dLm9xIwNgUoq2E9emWBbUoKsyoAeJ9p+bRH9T0jFG2XxoFOt4Zci/E882/RThuXc
gfAZA3D/UcLJ/deY8GkxxR24YpXq2SEkIKfmIcopOxdSL9+7B98WPnCx7+HM6gzU
JaxBNd8SvxzhVSO/g7AMUIOH9rKUwnJqIlgSn+2txlb+P4jIFClh1OGp52VY0OLN
+JlmzVKqhN1QbhGx6Q+rOy97nA07eV9ftMYebdXAEUKpQr/W+ISNDob5cUsGPmgr
aB5p8PXhii2VTjlsQBhGiftPmCDdMtmTUMDRcctUwZwf4lI8YRy2pAbgbfTwWq3s
JWFgcfhZ8bojJGP7RBEzxRB2Qj8cJm/4T6eA49PoBTqNFY11TuSFgr1FfpZVVOgx
+UY9I/Itk8Ah6hWPsdk6N0QwZMrxPwmvnBibWftXYuR6ptH6b5SGiv9m3LZN2/c8
z0YvtVuWljs2XGX5W2TBMQR7A/yEm+iSvOwH9okqR1dTQlXjjI5oTjeRObM+YnFi
xoijd8f86xsg9JuvTowfgVYvKSA3rKlECTdOPlA+QihjSA1lCNsRndi3tygRIU4q
zZ5khBQLU1Rs3rVHKteu7aDIxR3Z0luj1Z88mMSH7Rw0cvyAgNMOTVS0+6u3dbYV
1k97ESfN6oTiBKdfp5sl4pCXao+Ui9lA4d6mJ2ImmHrX0JFAAoym/2LYkRTCuYG0
LiR8Ep61ee+/tu4X2J16WbpI5N1WMCSKWBaKFb9JQEukkqRJA88AfwtNnGxUc2G2
gjHEtl+sS/F+SGSza0g4N7XYnIw6WJLMeKIrLBzLPK+5P4zBXE+HRmaa+xKSoogN
ZjBlyWt/N24oVzM0XW4X5RQbXYOCDhD6iCUMZ7BO8hIpwgQmX8wPuAYM0eYtO52Q
uYR2R91tUsqNdLaLGDm70S5NUluNP+Am9izUX2N8Q7JEzxlVUFD16y60eYXug+T7
gD/oul1Ia2/lUpRJf2rYsW7XG8cp63sVI0+tnbawkAX4bv3vi+UOIFE8SrDBrVe+
IiP9uBmw5c5AyZiZHv50rzqLnMmIOnwIygJfQRagt971ymDw8MLjTx7BQzq6EgeH
CfQ3Qo2Ml4YZhPkRouxi8kGEwD/bYxBP7EOxoyBUzKl0JEGQuhm8vHt9HV9R697p
ZCHdZDj9c5qlcs1TYcxc3O87YnOK0yJjW0IGPI5NIh/w/lR0rgkRWDHuoGogQo2r
W0/xFsEx/ykulK9aSf8EOM6U1psL/DX/Fyrdc39cKMGxcNkaaSAsixCqQlUpmeWO
z7Jukc24pJFXi3niz+J4QNn/WNOCAExQxe13/4ezLldxf/RQ9Ugp4Pr0hHceUhiO
BGninTlvClJC/NVDY5pfUj25RCbhx/rK2Izff+Lj5wD16oTB2Ypdvc1sj8QyqbGu
Qq5TOtXKCHHBowyORZktluO1MYXc/slLMPiGKOKaG6fRO1PcvBBRHOouGjzhT484
oSB44RgtROXrd5EVpUFHhIzqEVSr9xz3DmVC5gkgOkvE9hPkGwlYVeluRqNp4naM
TnLxKEWUIWlCpoWKcG8ULnd2wQVqBaK9GIcs9w6juZT9oTkmVbYNg0mgW/OyQoA+
IoKmmmgSLeVqL6ZNwoav/jZQPJFX7m2/Xlr5Dqn79Jvc3wGxFO7Rq2j22jlIIwZP
EDIS5QW22mnX0Rw7mQwuTj5kGXHQjIQczBSD0xJ/z/DpA0pTiPH7jhykU66n7qCA
ct15IEPw/W+WPd1hBXEIJRazviWZx4fwlIIMBOoHM9k9yt503EOUoXgOn3RbRShO
M6p3t9Vsl35OVcQVP2Q5pVOJcZDeY/RcaF9o148ozBj9ULSKSGIbMWrLfTAdU51l
NM4H82L92O+lvyLDM5owgObqwBAw2WMlUqAH/74s6+ttApIRGMFmwEt/d5r0OHQP
piTSKD74hxjp5yUEiS1Fu9MWmhb0i5NA5y+KZ2QRbJaXoPm4Z02W7MGc/i9aY2Wd
9s0wXRrpQVC+BG+4s7NdZhtm6dxcNiK7fQ/eVMleYO+/LcKg4skbH3uieR40Y6Z8
vUbVqzqzuyOtO1KKgIF3i40yzwO6dJjKulUowkT0rpX7aiAFQgyJxpS2cHTFFWFd
0v+R7tILe+0F2kUqbLw8ocEhVdFjQX2AORp8iqQlTba1XTlKb8gB3OJxoHmt9nXL
AfpNDV+vJeBJ0IavZ+2usqmtRK8hOd60ureXQJGE0W5ktgsGqW0vGzTIk9DxNTdH
4blIN98GiCfsZDBaawQZAZ/JKd/yLFi69s+yO/bpLoBvRHzscfeBAqHDLwywVptq
31nETYrvGl/vjBJcPVNe28bbohPiCBdL/LgGVCz/wD7iqhlKewDTK7+/BAqK+UAI
S2EZKHz0/woP2v4itlMzHkf8/QX5rNllXIKmT0pi5JcM/YO2EkF+MwSseV6bTSDZ
XW43to+63FYrUOcWy2z5Kd4DbR1VWlOS0t+1b0XKcRh7G6r9SNyoHIqiGvntMwQU
GThiFyw9SS/aK/oeHpKSC6xnHtxx7ICS+Y9mAZDMfm66kABW3XOE2uAwNVT/Twf+
Xz0I92CtjCRWtJ9OJMgtMoACZlbdhS/oDzM82qTYTuie79qUOCHOwILUdueuT5zs
cWwPVp5SPIreZryR60talwD+xAE5GFPS24H8WhHN/gmoPDUoHYhMd/JWZJZDlgh5
Fob6BZsjoGIHBzL1UocSnedmDfsF3gg8dMhsRsQwBMxHcUnU0XY378WE0T0KvGfI
6hkR2A9bY5l8aHPOUTnsBsA12ovWeZxBW/ky5pnK0EiefcFCwjCYzrHV3DdVwwFS
Rg75z2JXRxTjhanWRiE1m5Zi7dTeAw+hZaDwHjwGWwj9fIHjOumCOwM725pPzcbK
OiIn6tFhQ2HDfiUrLW4+vQwc1VyvQ98kUWMkkbOfkBGsFFTcPO9HgXP/shJsxtMI
TR7F+/YekogtPPrlxUbO7rzBpqEioo2kjPCX5v+48d85xZRMjM8+4fcc5i3rmYLF
jjn85An6gswRHIPE1akvQ6qiocceYc7SD/hA+sQh31cg7TVidlWuivPV3PFQmx5I
VcH1wU/hGOgOwTWg7GsU0d4uf1Gco4A1QwwiFFEXKz3wTOM80lWJvSrI1FdSi4YI
ZrCA01dc2E/ALlxbDSxePlnGajHLDga3UkUqwP09VjJDrlbQFzMW8iS/MMqwixTQ
wZx82t2rMoXzjOR9VLXNVbpD7SzfHYwNNKItltmjnHdmjVrR1KB6/PQOHGe0FCyi
/zWTLde9acr2Gel9rJB8/r36ESa1bnDrSpX+3AoEjscwtY4T9Ei+1o8ppXra/H4H
0Ttv628cmQL1jdige6xEXVkAdL/5F2LT9Wq0ZdiK9VpKfg2m3qtq09dz7OO4Lz2s
5xLy+NATZWeyceeYOeIjF2VPCYeBfLpNMDU0oZNSRxdly0Mz22e30TwKA2KfAeYR
Chd4Ihps7RlZQVhmeWdKl6EwUIx50Rps7UZiXEtmh0CAy79zK5M7xyGZNETEg40p
Tyz9tJqKu8sfrMAA+UMmWRqMmhH1I/CnZBIUy6Nf51WU9A+7ANMcUGSyce92bd6R
avQyDOGwcHe4x3P1qZx5csk8Itp3QNclUrIXHjCeYyrRH6m6W1DtTiN9u99NZeXz
O0g/9sxWdzVNI5em5x8OdYx7DBO/mMAScFyiS+uva4V3QI7LbX1Yl/hawzjIQHKS
6M/e06dCk9eFbKYvEN/iRYqCRAiYdpZ8ymCKGZz2m0RvtKsCrUpoZ3U/d3WFXK83
JSTefXunii0v2CWv0L87uuPpXSUGZYfAbSgCKAxTlhwmOl7nr4DsJcc3yUgk+bMx
PBuggub8c5+BJS+sg2S4/Bj1Zty7A05p6cnEuHEfXjicA93EBeCuKfeUByiTeYCA
SQeXAjj5dA9Azx1U8oUVa0G6X1/xX14v4Yb2dKyl9lb77Lo+Na8jYoCYL9dejnvD
j3oHPkZP78y7ardJeUMpgQ98fW0Fil1XSSBRiDdp/d/86M+IC1nB4BRwXjWyMwzP
dmqqn/iOeDw7o4etzDcHjSk3WkuB0pWKaUEDqVdDSGM9Pxa9E611Jhfr1DKbqanc
eAf3t8PFIWPl32VDjCChBN16CYubcg9mfiKLYcarJ94PklaMQo9nvZjRagfFhNj8
YmcW4Bz+damtmEZEReNz9i6OPP59XMl43tdZiFccj9e+YP9bkXMXArrQLFHN4yWh
WWR4ySmgBbdLhZ51m+jALsKu1LTCEI9DiR2dtN8gnL+wjtmyepsE1XWxn9ULmxT0
rmicsFlUgUFGmIt7XMYeisEz8lwFFBQLkgYYb0oaO7Jy8UbbB7xJ1LRq80NZXTmZ
6LtxK42/q0OmbUB5DXbi1tsgd5kUsMfR4VWECoymPGizKUirIlRQXnpVRm7OF/8J
LKsV1h9lZd5cRGA1InSwnD2IwlsG1TufHVglhjaepbqOK9NZkKic6tvQgcKsK6Wt
AnNP5L3SomH4cSQ+d66Ycg5h35LZMFXy1DBXPL7mpE7QaVf8Ol3cV0R4B8jqRFAu
Wsfhxzgyyk05mMS/mdiLBPS+egYIUCx8YFLBRV3ZvZyKS26f1bI6WxTSwWH6D7tK
v5bTMffDsYEbLIBk6BKgWzUEU47/oME/jdFmIrPFmlpcXZXYSvRMeztlEaOUAnhY
ULu4JYGF67vgDqA17Q6/d2NLSmqB68k+4xDBBDsb3R1O2POOUBIW1ofJht62DG7p
a6KrdDjCfr+Bf+TmjeXnO3yZiyjOnZ2MHx50ptIONJIY4ehXDdCSlNLG2gjEbKdL
ppfQsqb2H4vDfTUIGYqIxXLwg95vLnEQn1ojf1n1svAWMCFVTIcSkV21sAH+L/fT
45veJ7ARqWRoTQQX1kBEDRGX9rJc9pU+rPG1lkcejpHYlqlhTW00Em5zqemSfwII
n2eLEMKa5rfmYVn2sPZSe8lCgGhcEinPWUsu0MPTgpJizpmyseL6SO3QnSs1W7gs
qEbFimgwd15L5GY+EevKLBcrYoDfLZPl3DCcqphbUljlXob4SiRG8L46MGoacCCf
ZNtThUr/zBPHRMDJfua6POWaSk9uEDgG7jcIe92mOO0wSNsFYvCEfor/ja8IZqMf
HQLXa8ZCI+CNZS952fUDdlg+JTfKyFCtqYt6UB8+85GfwYe/j8s+xGDwsWcpjbNy
DuxugW1l8hqkbQnPwwTSUaYWdFMEb42BL6mKzayA8IuhJbm5Q9cGcPQ8uQ0R5Ri2
vLP03v/voRKc63f4wehHfN+aIYSQfNsR5dGzi7dWl1GK7+A+QvC5gCBfNYbP5x3m
CQaCjKLMKyTbDU818ZpqtuCLDN5fWtLcdgPE76/yTdBbqkqTwihqiMlLa2ira6j+
3Ch1riaeSLy7TLTQrlEPkKoQaVN+uzK/k/G0JjUcc7sa/ys0uw5NNNznYA7JNvGC
rYvGSFRweNkenxN/Jt4k0SLQXA/8iEfn3aPL/rxe6ZjKE4OcUaivnXWFmMzL8lGK
0wIfYXotBjE+yiOop3RgM46/Z5soyaL3i1eWrkasYJFZ+ae6Icf20tDZDlMMyuVs
qtV86LbgESYoUEWDqbb8m8DrguNB8EYZ+mRomBc6La+QLwo2V+kouo/umRDXHxzM
Sh9Zod7WkQCx3SD9J7O16t5fTb0FYAjQgjNFVn0ElFv4i160RtnbEIGQ1E0apkua
lzL/G4yUJfEORPzF8zYkGUNUQSYPDC3nShsAefp63O40TUBGz0cfRpYYs7WiAX6V
`protect end_protected