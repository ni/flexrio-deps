`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 20704 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
hRRAlfE1xLfeNfywbrz10OtvJixhnWeYVQCxik57Bc/aQN1QYywLuGBByMy37KIB
1/04XnD5N9Ae5pLg5AavmwexVzBj8mDypK0RDD6vAltL348XLy7eyOo1mfxyI3sS
bygSp5ha4PsMsg1yO2DNOsYnmOvtpnP9bH6o/tfKxCpwY+2wE8UTTfoscciDBbf/
IJczM/3+/KEJfgufIUJojk1fAcwSqGFyd/+9S2eYeJBzn91dJxXLx5EG9kQN3uDC
m6GV3+4P4lepo83hMOFDK/QTmFJiOBdTJ1Hz54TTi6a3YSL22VraJytfLSSv8QXO
hGvtgDdrS5WzAEPyhByiq/cMUP6soKptqhU/csUpCbWtvhyawwg4fBUKF2+76OAa
g11MtVJgzY0/t/qzH0B7DCjbSr+aryQ7Srk/ui0zS0lg0MwVXoo3qhpm+mGSdl37
wuRwmHDZiKaN9DuDtQ+vKaE7zRRIfk67xE9cA7URpOtK4hvBI++3rrg/K1V22mtu
DQhakfLmE3O1bBvWyjWzeqy1nYfY9lIejSlfXuIKxv0F9abDDfEL2DUVIzcZc98h
DVBIcpyU9rQabHQLAj/3GbGu+X/RIA7sr2gAn84Gn+1mvy/0uo5ScrEKR8VYpYoz
8WCfKYEtkv8y/TgVPMNF/DORg5a2/bkjrI8+qi9+LCPEuiYkvlZfDWEwXQ+ttGM5
Z/Z9gTE4be2sy3Yq1t+tOIEx9wyglDG8khhDANqKQdzeZOK5Urr9qUjVLWYQI6/r
QAOvhkliifzAinV4UAeAsxdQfFXNIBoYzcnX/22l1/GOgTtZMPGAEJDrMPlSR99j
vblVVRqo1MPH2DtF0rEiaAHyiXv/FvtnusKQFHyYi3CijuSyX5LJai8gSpLz80Va
4svHP8J5aUrL7B20s0gY/Cu+3UFZAOzfI6y0rtdDJiVds4qM6u9rONzQLVC0/PmO
edDkbZFIvZwnygA8TwPc8sj3yCemdbzH6KQFRz5kj5n3PAPo4LNDJMxIGPf56IVo
BUNKgleZeBhLWpN+2oo1mHFw7nVv/oVHk2EpfQj+ezWDVgktbYPbq527J1y9rOE2
vr/PdlcieNHsFhJXgv2cku+mKSQfkptzNqdG2eFw9LK8R7g4u49TnnYJuT3vddub
hcaufMfr3g5nZ5dig6b/uQFWQHOSRKhjtXX5APHm17Qhyrq1l7ZU06Cshz5gPI7u
+syHH9K2FjS4u0zvHTwoYMRTslu7Td2c6Em9dtOstbVbD/DdTOq1aHPgNT7nM+RO
QnFNvY+EKY4mf5ZJ2arcxe+fEpJdQ9ZeHQ0YAgxujLi/0PXozq6mdWuGb8ACq9pX
s0bYAdINMOtwqHF85jsAOHkCpj++DaLFfW8d/TiALcfv/wES/PbRpKPFNO+xLPoX
NqQ97JFuLBkUDw2kqFEPYXcRKAsjY88B3gQw62ODJbpwOPAcu9F6r3TzNEJ+zq6c
peyy8P26u5ybhC7pgYBlwulfjhojZei2u9pxrijqTVunRZtRzzif1RoCdemn8UuF
Q6oRXstK2bA1uWgm1N91VRq3LYKtwwTTlUfamwPxYivnFL1vsZFcEBfdaUOA24gJ
CoAYICRC8baXUMRxwPjK0v6ExjlbNhqyX6q0I6YyQ6vU0kDD5+wfa1ncCz5HiFnB
b7BQS35wkEtKD6MYe+Fep6VWzOqNPytgegkugBvFazG5U/Ba0Vvq7dQXOKL1G/4f
5oXwTegQyV1jq7GzLUWtFi6wS25r4xND76/v7R5whdsY0uDcFDRlpWFo1xiPn7PU
qEoHKH9YaOL/Cdbtcd1XzIbVKkB3UE5T6fSB2Jp9nqPKOBwJEh/W82N37B0zNgaG
AJCYWvX6osYuW4Dd6r8V2yHS5R/zy8YdsP72ja0hQNevb2FMMOCPlwLgvzgXnE6o
FLRsMyCDKVO61m3PKKRzBLru60Mxhurig+g0XsH7i9wRgTMk7FV+azrp2oEYZAcg
moOowEp0phb28fNQ0sUxxcEcg63f86wrOsq0kHKIVWZnbW6CYQAT/c1bGkzvCqyk
ZL1gFiRxLONdcEMb02WSH3tXiPbpQUNrhhS4n2Or3JK1XWAdb0ryaRt1c+GXwaIn
3I1MpPe19IrsEp8uRTtpDoe/b3ANqVSwNZjc7giC75EUGBjR5sKTKC3OAHfHgKs/
15ka3Z6s0kA8kWLBsJMVAxhN9Q6W6NbOQozEutgleMOK3FTbbDveaNkodSvrDK1X
MURutu3ahwABm+QzgzWxKMDpnVpRnGbI3uY92iP0QoK6QM7I4Aifc+VWdTG3G/hv
fQQ5P6/GK+TJTa8MH9NBaF4NXlmoeXAZxALy8bHyvpQJS9g6al4t0V+85sgkkzTz
CeK4bTVb1MrZc6UUTDEnnCUPuFNyXQvrTEzt6bmr0uW/zBJSTvqqMf4btlRCCW2i
pO3LyNen4IilYrm63b6MDmdaRx1whgm1CQtqop6+jlBVF+ZKseqL/tGfgmw5V9/f
sWQouvpM2I3cQ46Gw5C0M4r0HbFqdasM80rTgKKiTyXUE8WCnZu7Ag4yAvy9CW5y
HvbVAsOqYzy+FoaxvaWv9/HAjeo0uYNcjIPRwDa+BiwTUlufoQFzBjMMTjnL2Eu+
+ms8y6PGbQ0TEOJNtUWk9kqsPZhyWsLqvkjYeT7soNnsTjOJir+WFpQsUF2nnCox
sXyzCoPUlbT7/eothuR561ZFOWn4+KIO0EJGdnh6mB4ST5IOvUITD1pgTKNuS2SX
Jj/BXGbt0Xn4XNfQi56plcKGwc/UzOkoJn5LVpLbGXCkzdwtUiBT1PCmeLXx+I/1
NaBek1cs7tnWjGwPSivimaFxFnx4Gz9zc2JmKl1XhE4kcwc0E405bjGPzN8dkn+O
cCjrNkwfj8PXwOk09lzCbN3fuSMhR1bVGGddSIr9ETMMViL7LXlt8z5Llroh3Tku
tdJCuUZ9RK2+1dinlND8+3mmL/TeCqjQ0tBK1EH4Jb7hW+26uMkHKYw1FVoYuBj5
4vaBSMlq9iznjSf6vMgRXJiymi1KReqSjj/ojdeJZ+vq1oDzUSzlal3x8nf2p1sC
7xWw14vwOcA+zssir+Xt2hZ+Vr8G9BBq7zs6e37wO1frzbhvjc3n9e9d+C9MCatm
pLiXhmyDoCFhdVpX159a1v6xazgbG3z7nxcz1gSS+cPbvLQp+LSoRFpcLpLW5Y+V
OS6UPelcV1oSF/ZmIHQ7w54c/MFCnF5zi4+djjo9xnhdj6ucITpIJfsBgzzXA1VP
sQsm7LRFKeR0aAfKN08QA+q+IIFvGCIpnmpMHXUN8dUi9UMS7J1RX7aO8nmNtbP5
BFLDGyOGLts8qp5bThQ0xdBxcURpzLsi41N5ffyIih4P/AxOnDC1BKwabZUi5fAz
b1J4n5UFL8t9sp/BkxUP3f+gukQDhvIPKJ0d6B+j8KgV9NLBmIy+Cnztm8qdC5Y7
YcLCg3g4zRXoaqJ/n4pIZdoMQllSFXZ01ChoqaUzHRZIiYxgiQFSItOIPXeiVTAa
oeXTQDC4ZWvEbew9jyIE8DuaDZ0O1pkduBfNQnTagX1knV2YRusP8UzMOuUSlyzF
rJsKHE18fzOWyCGl2d3eDJXNgn/YMj1K8vpmvfPHQAQhf7tzPnRRgcySzSpbcTMx
qvjZlhEQ+y6jhdIs5DjE2CFckihJzMXMdshqK7+SFNEiNvbR6kfq3cuFPsVaCkQ6
/Qqz/abdINPzCxojKxpe9BMk3pMATBjKcfOJjya2lmZYFGyg6vop7q39YFkHNS/e
+FmxjPjWEwIS4gz5u/8VXuTZAHQFwG8IKmDlCt1qcJlcW4ywbRvp8LDVdDlj0gla
Earz2/HsfK24zgTaFqoP7h6QqHM/RpkJLNEqub57IpDsU7GdouYZEyb24gB73/66
CQeEfIYMUOdm2Dg6yOID5mV3tCiFQTm+plR6opR2uBleQPFFYhCrfuRj0SqmQUNs
LWLj9jvUQ5MrjbCJSlB6Pd5gm+id6v0UwiLt3nrgZyyRMQyrkGvsezrZYdrt2se9
xc6JfZkCRgMOghWjQw7+H3TTywTs+S2bVNs2QF4MC+mWcpYbKF7y60XciY7NhPlk
VVfcALABnULP2thymafR8fFYbN1Xg2qCR3zORqcZp0uogAwCwbSJJEnSAEtSJ/vb
OYZPXskevFPt7BlUZNV9+kZ8eoq5CLpZz33lazONA10bkJAoevP+iHB5+5gl+rCy
vv0m2n4uznfSQ73xOT2Le5elHIA7kMSVQDMYj580a3jzhlowvtpBwuWI0QL1fQqx
/VR5WYEwt9v814gkCUYyhjGf989Uul4E0D2mNONGfa5DG8diJmFQGJssNkEg8NMo
M3pludWGtLrgF8a1FMx36BHGijGnL1VjPACa6dvI/rJYXb8N5jXPwxbz6KSeH1qc
v+WrOa2V34SQR3ZnJ//ImY0cKT0vOE3CMNIrOahsq8AqHK6UujCm2lRI2qUQ4HN4
OG7NiVi6pjgFkmygEIXIHzhUYNbHI09Yze9QzHi3HGUQ0Kdxvzi2kFgNYHnSGrFU
FJeBAEDQwVU4I4oUefdT1zIwtab7W9kxypVo/kYyjHbf1SkSRXKryHVyzGTQT/Wb
ceeCdvHRYzqZLGrziYlUTIqL87yrJkxWNgbpON6H19cOW2kWjxUMSW6pxa1GNyPC
F43wM3CWCM05Wf/JOu9FK0oRINx85LVPwaPW1GDkk/5mBkj+qrzDhua6YGOm1vEA
f3T1LsCHS56XTlPkFfPY62nZtmvtPi6CwJNWoI+WZ4vV/ezdTo64fpROnXaYe1aT
20ZcY/8DUWwORCzL+3rcDeubdWFR+OnpyuXRLj+r/OlM/rhmLPJyeVBqy8GdBYTx
gcWrk6RidzJ74LAvbeMAdqVZRLDb2/JhEno34uhPvo+5SLPjSuQIX+9wQgHUGcC5
Wv2FJYhcNkSmi1f+HtY+2Y0msgHZlHxFQP4OPKmxs9/W7B+BF4OfkK/gOr00UDBK
rjIXc5ECibpkfKuCWW7eq2nq8d+M44DJNUK7SmlLHxaC277va7V5pCLWYuZa+7D6
gLdW1h3GuewxMXPSWBWlTVrl52uas8U5mbvnGqqlMeY+nMjqoU4RkkZwsccvaPIj
ZaXPEaAjIhHl6mfzuyucbT9alSyImfbSO23FOzCjMPhbLSCjOl8p6eW9rmp++OY8
pIvdG6c7F5nNCuiy9W5RpzzV8EpbmqQHuOvIhxOnLPWyAavhWuYIBUMXQBz05DHM
bN6Y2e6eD3VX9godBJcBQpMBwRa3z/zFqWFQzACz6Ac0vGP/YXlmpDVVX9vUPBYF
c6Z+na1wWqWNICKn756DbHQC8dWMbPa4xSenuV2tfVWmcT8qgYA4d9F5XgcgCsxI
kE40+ZKLt/HZ2bOj3fZH2OZYpEKWldXgkanhhHVEeuyb8jhTo2P3Ze2+wsBkecJm
gZ7gMyBcT1UgzEjqV+n1N1lt8WqQMd5y8snymD4trBU1O4W/WNx37noiLGsI/oCY
9g9jp5J9c3qfcwr+JXENDT3mRGe+IxVhF1soivluHeWKSK8ZJbw8eMItnu/Apd4E
TDmgdbX36DrE4oXiWOjN9xP2R+MieDl5yWvP1a5yk2X7cssw/1BWAoglZKpanu9R
vnKHesvI2IZmc919RaY6sqKcJeqTvrY9Is3OMXOfDnT9+Y/LREKFntZvBUL3UMBH
KVcw1oHeFw2A3zEv7QjZdnmy4Ixg91Midj/mc9nQPFnTYNeMdPgFBFLc7u8ci0CN
foYwHSRAoTSFhXgXF6Z5XVKWOxXLR4w5B2dLr5hQ8JT35khCnxyjnPGgUH4N351C
0oUhCwKVjPU4foyBGHI98cNcfHRHEK0jCy89x7wB2jt38PLXFZFnMJeoEoi4dEIP
MqyCf7CPJQyV80uCCLiQ/ftqpT53QchojpVMgLCuCdtAZ7FiFIw6LJDH2YAiLS4N
7fAi5rw/1BkFjdn2dyORvkNVMAzNsBVBX4ir0E31vOMCvO8Rh2UmTBSSu3O6XZa9
x1YutYd43ZiAubr3vKJtfQjSn5rhfxryvTUBGrwOh/nidvuHDjBzdpy2lrCzSbb8
CZ0vZSRWYYAsAkjpIv8q0B9/G6AJdqPAFFApztgQiXLey6t5mVKitbIMG+4g1J4B
Y9l44k0GCyqeYCKbwy+tO2+HqmV+vQpxzQhxGyXuenAChVTPtCKHYHwiEqAuK/Yi
Xbvo8x4aNd05i3gZ7U/VJxRLRsxJGvmku04d0XWOrLGDDbdbCOOp9CbO+qGstZrx
ZOEvnX/WC24gjoUoM5ruW364TV0DwkbNbulrtTiPvQz9O10n/r/pHoMnuyj8lfXF
4/N6pmXc9FozxMitW/Bo9ysvpVkv0U1slH2ZxJWA5s9ZNGizXsQ8p22WAgagPWGy
0BBUogkLHDXZLtu8NuEkxLV/GX0BJs1567UBH9wftY/HAJW+OKcA+amfyK56gKtt
b3XubcZ/TkrfZd7bxaUbK1GNYUmVD/l4Dr5NMtJYN7rJhGFapMzMa03f2HUlswyk
92Gufudh69MrA+FdClzUA2KSRBj0yzu5Q76Y9a1IJwp37plABv1aAko5VDiGVeFY
f0A+wg/zA5UwDJTaHorU4DTv9Wc9hYHwvF8CPANW4v6tYXhZipmAiyALuclD643Y
TpIQhdqAGv31bZPBX93W/g6xRLapundH43ZCal61PlGVw4txiGmDCaj1EYZ5U7+2
q0a/l5Wg7pu1h720hebTVzgkIa7TSfmtNvrD1Tzhwsks52XCtStRb07adr7FRjqD
yTuv/dabsLpMKiKDXuKj479p7EnS7MIu73D9EqGtzbiJB+J2ex0ATHdMNrCmVa/U
i8+PNC3wa60Y7q7D3cJ9QgFlzP1cOvyEw/FSSJ2l7uBYlmna1DoTnEbMEkGWikHa
Ahw3NHfe8/Gb/1d026AkUMdC3I/lGc39mG/WKF2cQmCMU830l3sLtOSp1p3Suklo
91ulYIY181HMw/6q/4MZA9W5HsuxhtwiG/vV+uo8LQOJ4IvwwHitUG877WAxcKE8
MgvgQLU2ig2DraM09trWNMekUA7LK0GPm0il7vHe1MkdaPwEiF7nbjomfbLL37PM
QgkxKHg1OCnuD4ZeNPtoFpsgDcppH79u7/vzDeyCb/n4CEMjAvlI1QLvVXPyITQ8
e/90HuSpj9cfdWVA3edpWw5nK+E8ez9D8MV2/CIT6MU4LqT3pTEJM4l7Qg8Ngu3c
5M52Sr5o7pCKTswoWl3jW6gGCnMv/opHtR/SJNQYK8PkmT+nvSHJOCbBiIotEVSJ
FDp53YRX7QkJ1/OSgGc7gMWttqauLPV/VGH4zvuUVyzkQm+HmcjlwvPdwqtk/KiP
B/SHoDqfKMUA62kP+duknbqJiPKqvDcRESCjflEwUjIlOOQotgZvj0ogVD2wNdDC
WlaiATbiSFvo5WBxWU5xJShfLm82kw1wz/8i/6aWa8EA2hCLbm6NMnCqInt/mwBz
cEnOwSIc1bah79wvpXnaozOxDKd5j+ucau7gJV6jjA7ya0Ew+Z/NJ8mKMg520a57
As39PnQTIKFcij8p1hCYBNJg26cUsUGUvtAg1f8oP+7mLtbOemsBdIKuLUhlbtaQ
ejYM17e/AM5tOgeR2LdqKEojhugrKTps31ZxpFaCO78ZDcXZH8RIxF7CJhFFzx1y
LrHCU3FcRmW8b0t1hcw1JH4ivqWeX+u9d/Wy/8blETHr1YfdZzinMdMZkgmTAWvh
e5f3laW+1vOkfNQC/I3t/gfH1UMRW4cCKGVMC4mWGLYeiL79F/lZAAtTbI3O+Yk+
rvq+A1CuW6nQlGXSnE7W9UvTLTEMjNgR6Fqu1RMeEtA7Al7Ts+cGt3kKOmgX6Y8t
lEG257MwwIoOXjJJAHOt3t36oNpUyckzka+ovfbpQF2lemUwoeJtX37VRtc+uN9H
Nv09324b46y4WRWCtmWrk+F7gvYjLtigdTJWYWtFTGuXXGRixR/q7nNv21ZMsCEs
9AzOe68KfN7PtIh5ZM+ePP6aoTmn1icQ1+HSOlVjBk2wUIo4kMthQ04xbMGQiXeQ
tHrFEvz2r8SsEv7lNdFQJwj1nR9thCh1ess41MUwA2NlTnGdIzDEPS5uv6vSHG3c
UgyRkSvf1+4QceRIZi6pMJpj9XXWtX7EI0YejJKn4Ff6E5eVXkDngHhznt91/aW8
msJL4Ibb0dkQxCanypDwxK3I/tu74dF8QlsKxEVw1qFzNDaedS4i9KSRm4MGqvWS
8DgiNSNzVqBydYgNWSsgV+6vhkEaj6FvUW9gRt7gYvmxr74R94/RVLbWRisvMz0Y
SPgedmfbS3Q9bfNXmnbhjDw5CTdUX5RvxjyARisoTiwGBemqkb/R2oYG9tk4xWfJ
AwVR/aaj+rH3MiWasIjXpQ+jIeyG83x3Z4T0Vz3fyXNlszC+OueUHg7KBtJ+8xEO
efnIP4tNeAXhFrcvJZKUT7x8AMPzGwtwE3j6IC6XnJRlNlZHuP2b+DgfVyDgvHsb
69/Z1hQatjJh+WOTweoPqhtEISLYNId4JBkqJJ4W1hKV8bv+vkmFzl9NsBzWI3lX
aFEMcb6DdSy62vE83Gz2fjXBGYrw28BHmFODcuCyu6vhdd7oGmWCJft+NQ9HsxG4
GvttzeSAcarqOUv1+FIay3tg87XLq2EY8EgI1/Bax80kBm7j1AlnWR7adCxISaxx
22ZAwPk9hKBu0qfBIiyr8Ots+ujylIbIoPu9JBtL+2mgoU42l+FL6F7PGCgc3I9U
pKKmWSsO+MJzm0N/sZeX1FjjF8K0tBjOOwZ26fvGxBDP+EOtIEgJj9EqmYRWYLRQ
gm31LrfdinPbJA+2+OUMykwAGz6icXw8l3jAv7aF+eSYsgCR222Ez7XyMrlg1C4E
5etGThCBl6K7chKMtmcfma3bb1/6VXuca7O2RQv45ZpfUx1SE5U3+7ambC3eU4VD
RAj9GTxuogAMVqp0vEWYVx12C79OMYPZ3ieSCcWoweBQ473r1S+gfaDJd8SatV3U
4chgekvBvt0ojT3CySoKpyzs2r86KL2N+8qJV15KZfJ2UrBfh6PB1nri3QXwcnSb
+8558uzYVVi7vUf7QJm3jUU/Vn1aoOW8kZwOF6CfeEpsYF0yAacI9sRcD2h5CMl2
h5DFMNrGk5KqZRr+QAhqFSyHGRB5s1MkLYZN24qygSrVybzWXqSISNRoJW7nfAyu
9Fl+PtQHMOCv6wYUZ8Me3qzCKSfwv+leNoZKMREhRymwnGU0FGb9Z2jpXYegwrZp
7LDjMWkMvVu9DX/lv+m1DH5eW7gaYdGeeBDTLhLbfj4Mo2QPI7fEo5PFWqhMv1n2
XbeG4JMoBlOimdIXoHvhfbBqUJRPqZ5YlMZkA12IL3l1zOW/d5IsfFLg3gkEOsX9
6qoQgVzu9EVhmjCTFEAiy/HYQQlKXM8iScYgqVVwZOeC+LIrMzW/V3ZSKFVNacRr
YWJDjCdXY9UYIKMwSBe5nvFsBP4cDRNDWB2zshAAb1UO8qpkZygFmwWB+ZEqb7f8
H5E/Xkkl6h4uyXAdQhiYafJ+dQBqndkKyvkF4DvGsGn39KDYYjZbz5k/eLMRIjdq
kIck/nJ+sGaBNiBzqM/Pn1zMVcF4Gpy+Sg9WxQE79DuTQyMsQNRbRn9JBuZnfwiq
fidhYTfOkX1geTgC3AVRvgMnwFUhhpueFqRE8G3X+/Psc1ER203VXOHZQD80Y1UB
GgMOc88CKyedPyhApT92pXedJu0zJ5BdCJ1Qkmm15KJS8tRMbLoVt0y8XwHckkL/
FhEkIopZxR1c0qAmWCeMZCqwjLNRG3IoGnXG0QqoqW/4HYwuDme8ZSj8J9PAnnxK
Hx2z8K/TwML5KmicdmljXb1rYu4fZmAjpkNVm1jOdedxi3sR/SlrmlS8wqbEDOCr
/2H8p6W2T1i0RnOK4tQJYJaJIfAwZAq7NHJj5/wL8YS5RFHfNupFKpZgcgFoEL+Q
gd0vgP3YAlcXoDbHuMYJrMM7UwupFVNDyvejj251jQXdw3n1ud03nNFX1MNf1lEN
DNjmkd4ymmlJGOx1+l/Ef2e67jWZroIGvksN7pjPLPaBDQI/H57sfE1AC5Y3EcBS
8AD7FOXqdks4j3ar5hX5YlsLEo5EdDZR0+PAxpFTQxVZ/2OMlikhszhT7M0pYVFW
eh3uwYJBFycvbdak54Vuq/0gv223+2R2vV8DXQV3/XdjZDsGlpeb8lxZVJtlZSP4
YzQkJxs77K0RWxKk/lvc28pX6PmCtZt/tLrxlhU/Jl8uPj3tMENZQQJ4cDtmgTH4
apYEj0shzPbMmMoy+Kq7BYsk2HMS+xYiAAUgCXYjS/MbFOvONx4PqOySLzdFcsVU
hk2/FWEyFjmmPXZdycWWK+SPrDrRKALKT8vlY56s8WevjQChLbRgnNp4dBb0r6uz
5kIpn93GlD0uCvAX0fwadIX2rHSYMoEJwuiALzigtg58g4oex+/3XTKlWgM+sAvi
k5FuWjKwFHibppBBVYpduoH8M+AWxSg1bORvQfFE04pzQg3/X8z17oUc9OesWlSo
+/5SSKOWiRjz8Jo8+DMmK4W9hg3+OBtc0mNeV/ABKrAZxQbJ3luPlYscbMnvV7XG
zmsKNU0VizFtbjTBL9AhoZQeR0njmqezEUl8T7qXO2cvcI9LUsYq9zKFRs8B17du
azAp7ram9vbzzEeDU8nMEqrQkV8zL4O0eYl0KHnJIy7rdP8bcnoS3ShXgqXssHo5
eN3nWW3xtuo+VTFwwAm7YViRvg6tvdKSepfu5EEZOykkNqnyNmZU0DZCNINBlMd6
GU4+6cWyH/RI2J+Br3StE5zu2rCgrr6BNGugnwSbXLW52l4q6pLfS4Ezpx+mCJ5m
HsIh4OrpLAsojdi1Fufktiuw/VklsLIp28VOd2OaMtsW4atlkd5eTXpKIBndj7Gi
I+W1tE9e1YiHMfxW4wSNRKzcDY73ezmeL39hDkR9AtHd3/5WxnNj+uGo6LtsL7gB
YoWO0gsaVUxQypNF2K56elp5feMP3hmU+SqLeb27KwpY1MzoMVsctt4PipgT2ewp
lSO1xrFB9GRHNmoN2AnNrQeAQT9+vxiS/nsXnnnv3w+yuPxNJW1ZF3k2K7cMu4bt
g5NRgmKv86AU5NYkEs+UVfGdQww9qpbP33XjeZWq8wMHcRNJR3fz08yvEcE9xkxz
6O1QRnqR0V473gV7d1UP9uS9xj/4CVcYvelBvdcyqS4MJNWh6EUc29IwxVnFxS/y
dkQF6Umh5OFi9x7afghmV2t/aD0WledfZ6IkfJXgCe+rXZqcFL/YwEpc83cQ6kW+
wz0hX6E3pqyf3RAsVf4gIVtAQvmKpYNFw139jBx9IBVAAJOwWOxFm0p0R48pj1y5
z0D5ZrOeI+D72M0wWW8xKFQeNFjIADvUjbFL5pGA/kgHAN6a1mVBvRDtZBC08Nup
p0xImamkOcUfch45ZTr/FWysf/mEAZw/PVGJltC6KKcQUAqgf8ksR51rC/CsiG17
FIGcKPFJSQgogqoqKff2Xu/IXaLPPGc19x0Rjm/QbZQDK2wl5Ef0SG1JdlWGWzb/
5fPA1mYYgC91lxRq1KsawMKM3x/AhZ0Y/Wrp6j9FvnjN44zlq4ai036l5oBpL7Vd
gYisrprd9585gHHve90MYmPG5J1CLaMXUkcCNFl5c0laiLJqhBcRVxxtgN8fTlP8
TtdhvXJ1EN8tvn7ruIiu3d8zlx53UqjeW7IFpbfw/fCN0tINeRlrYU9CoU7RoCjY
Mob9XkFHKMGSd5z3ZwSl6JBeiCVHCltlUYlrb9cit1DO21LWaXPO4TE5X6fNlcDb
ECUCGM1j4iBCNWQR3xN9ZS/L9JGquza0nG3mNsBlgJVzZD85fqDd42qrhLoCiTdM
Q9TNjSYcrtpwYnwzNqRCT4JYFWYfYJUGTbmHIqZk0pO5i4gHNjlUvZ+wVL3WTV2P
i4FejmFf39wLuKEA9kIkPmXixsdGffC0Ieb6RNnQNwu4gn1AjANFvaDn+sgC7sty
lnonA00bRl5NPkut8fTT68i0AKA1cOjPkD8rZz2MaTShA0f/H9erQg2C4Ar3kJ14
ZU1BKXzSLZe/xpIQ1kLJaZhpNCxMB7qWlJ3KwOY7TTUZezqIzChhTHUP5PJeMTWy
VZBK3cnxEkqgdYxUbIUUrfyiviXzmLtOrWg/xas3EnYwDmqSRLqy1RDk31EMe5MV
AxjXGRlrVQW6Po1B1OmhJ6DeIJcL4ideWrVyuSrWauX+EX6mLtcQlxuPLKCBhybm
pkvW7y/wFehahNxTWKEdnXGqvE8QRukdGWnV7RlupJVoLoreLSLSPQ3mR2dIbGFl
p0wf/0H9tCDBEgJNXugmANYJOWfITg4HHReXx76JJ3gcmBp1qwvRBVdQ5KSnzvik
MyYjZ1oGMLdHWeUGVLZwbisqXEyj7i+4buPIUf60e7yo3khFF7oH83pOF8E4JWT3
Nbmp8GiggFQoa+lpeefCuTiKALZFABe8dZioRYX8xliEj6oFWuCxz606mq1apzxw
efrXUHgF+GGDhIfvrB4B4L5w4dBJy4ffeO89tj+suaLpDXIll9Ns0k0VC9tF0LS+
/fKe/GyZ65Iri//aqeuhnawr84ZwzYKgUdSQYvy8GeetlRfBvNN6uFnjJ16So2FA
EGbooG3HklbqebmsxC18/D26rMio+GLfnskSAGhLowcpBRzRyqOWopB1GCVrFl7V
aBu6UdzL5MOspUvlNXgJW1IEWPf9QYCOgMzek0K+ibOP2LG1aHtfaL6da8uO2Hfe
KJfRklpa/yW654BxD2/KEpxeK7wn8RcrJIZ09WGziKlNQtbxbfw/FDTbW+3vSCyo
C+oZGfLtaTLuGEXpvBI48MrnfMw6iVsyFaS5b/4+qheur2Uq8C4Od2FlVik5XieE
DsyMzccUZKhJmsSS9TgLhti2lDcXjuSnyQpQqz1ye9gH3qV0RZ0zUrOx8NpBLaPD
185XT++AEC8yE7VtRTQrYWl6LQ0mO4HnkRuaVnP85VSvSywyLSGYdUobYfPjvK5n
wm3nInDVaZ9PuIxXgB881p0bspOb5+ZuH4JQuMBGeQMJclkTyEpuEivGk4jsZ9Un
JPRWEm9cl6Zvvit8U8bnF/WWNxTnd2l9o2tLGCKQ5ZNBYuRXR4aGE5Ut/rDpHufP
sxqBF9TunLZSvi58uU5OUhs7tj6/67iSE7bqrBKlyXY5s7DccJnFXrYOS9AheiQD
4BuDZC/x0M39kvUiA5jGmENjDZBpp4ZfsYNhy3r8ZYSqKKJ4Rpz7UxKcT0+gr83G
pxtNsUYDde+YlszUQ4ol4eHx9LMYIMqLzblLlLJjvyxCZchYP6CuGr/NZogZz0dO
+T1b0E8HPw5h9uxfwK9koQdYisSrPGILehSFcqWaDETueN9XFNFPLtR6Um/g830f
M7JptErrl9YE7keY3JBxc5fSuD2J3yMvwJvzhTJTcnHHEkDQjbq3lPBUFIyoR+Vf
BySkZXB479kBktBfPSEfsrt6kAjQ89lSEa80EFct6HyyDKCvmU9Ld+CeYhmHIUpR
TVnlVtSwlvVJSIdAgZ/LKMofXtABxNo7UlkLbpYesbdqvYvEM/pARpDjNOjsTCyz
G+SMDgZtu0WYSZU/3LGY1bFuf5l54YNN0Np6JYncrrfX5aw6Gcq27sUiFEIdG9PV
cbuNeYR1JklBlUseTY1UT6lnH9oMt1i3P8gSeonf4FmyaNEvRng56Jp14Jz291Qe
8++6+YeLZ/UyCf0F3caPDabGAXJ2ffEgu3tfqSWmUib/X9wu6C16Zh8gw5mRlkom
6AjvBwpmAY988DwDFp1/iGlKvDgzq11d7PjAUIoIyi0ZNqONkal5nPRRpX3V1Tu+
dUKV4fya6Omf2mSOrxHwPjV8XobGFPq5cG0+sYZRQmHtRo7mpi028eQb+XD7CcGJ
VfwVE85a95p/J2GIeFNGUPQaKStqZ5FJNkuq8AxwC4FbEG82UMzLy9wrGcmZWupX
MXeMdxd57ORHXWsTCAJxXAfQp81muLjPuGbIdvLvjoTFVsZZE0Ml2Kj8Ix3LW/68
KuCnl+Q6p+AI8TwqDlpm34LsuVFIT38t/jXHWaPHLhcFUEbKH4e8qDjWF5fOl0v6
pdTQGY0gz6XzC6DaQGYtCB3MNZRCwYvibUjFk3nz7oBWN8An2xVZNonNxe+me6Yy
WilrYKvBIH2A5w2H75rWN7ZO/sWFW6dr3llf7gqs4NNQrfiWWA2KSjaoQipZddqd
XN8cXeol+kFta4ow3xLz1O+X3m4MJVO/UKDeRO/mzrQMquOKNVw2QemyNZkDnIJc
jwvxrN5QBPdSpK8dLcC4lPZrJHKoTawvcnGWDf/5LkX4uNqjZDo3IAuzwyeQExkB
2vXCI9WUxEjLC+6jFKA+kAKT/1ynXReTOll2UbJoHgTJ76rBSicZFGQXkd2lOD+V
8Zq5B9cbc7GFWQiL3OYEEayjtXYyvb9tkmtmRgAFgWjyy4pXK6HbtXgZPvjfE37l
aDmGu7BYME8VhjuETAt/PuSe7+KMPIwtNKKGvFzrFLNuZHuUSd6KNhbZanouShru
Qr/XyoaK+IJGLIr6+bWMxrB2dX3j84ioh3c5DMfdqKsA++Uk0p/2j+8cm+3Wlt0Y
FC3qeweN+C2BjjtGrTXyhYFxbBcXRFW5yLC2W79nd1ai4NOcohBBQT++DdKQa1+0
5jvxgnsBTfbPYedJZxYgTj65Q27thuOgB8dZrQBmgP9GMg5buV6KHUnlsgykOY3Z
/CpDINOOhL9E32NG6CsPPUuCwOBTbr3z4nXNPX5DYhmFhI59MyuJzvT3UYPSoKZH
70ZVwNewwmdOajGN6qbgS9j7fUObIMk1AlBorYiIzt+bj2Adb+IPjK1083X1+6bQ
fQTOl7PGYqcCFdB3AbdVKMZEXuMn44DevtekfEjSmw7K6x7Kl4hf0ZLgDjO2DG+N
/Ii+8erjS3RGtyQO7j2w0kUcGmWja2nl0iR32H02iqEzORqXPYLApHyWKk+7IoTC
VvT0IVUBX5y8tgsY2r+y2iBgwDkPLyv3LewCwpx+yPKT1z6t2P7lw6IyIPtF2d62
ffXaCqY0JG0c7r3oUew/OfRj0GKSdLzCNLVngPIWaHQyi+ZVpNB3ZluMQlnEJrhy
4NTVqBORpXz9r5qzF1GLEXTO+zViNkXZhXtflIFK42ks507vKKqgiO5FLGi1dEvb
ZUG30m2CPh5HV1EG1ImdprDTWg2bDJ9JRv/ksxtyuy0vQoKeXTerXVLH7Ung8pQF
3VMuVZURVKT9beoCHqMIEaLF7anj48Z4RwRCzScKJaFwZY5q4cF44seOIKaq4WCj
l8Tj1sWO4Qgkk0BsO9Yi5Cl9Jeyq/j3kij5YViBUCbtxQCOx7fgbAgwpZKeA/hDP
WYwTfiMZBW42+qSS4aW+R1UIb+zqeWjX2ykWET8FkpnuM7Lx0F/gT6kx5IMQwsYL
vu+tcg86C9xvJHESb2tniMKSDQfc5UCd6W3bGo6gz70M6CA6GyUbaM8sIVsw0c/d
ZvhXBQkujg6yWg7JL5n2xCqFU3eOnnRH1JpyLF4Gtku+HsBeQf4SzLU+pmP1aOgI
VOKwZKtXGfcwBuprjdh9d4wSUN+7dxNc+QXpB23ERU6LVvqMUgbCp64+vEX0sW3s
nH0auhjAHn9VHnlDLV1hxYzQvKyZQUMYVf3QCqz6P2D2n7LwpoRqn80T2Qm/V0N4
HcDe+IlyZv1Ox7718A2pMCdAnDufG5ceLtFiUojKA/F90kQfGUqmZpPMqgG7PvBS
ysg2wSIw/amnjbjMWOpm6vVHi7VUQtLkPh2wp9Mb0+8WwseBv8EgxGWxBN6EIOLi
bKRkGr70tpxRXP+kXrRTmuoA/sxA9fwghuDYhh436uHk8X3vzpzk18sG1AR2G+ho
3BbttsdRv2Z82yveD4Vt1MDyZudenbzJlLu31+IRCuhPum0xEENIzkO4avhmWsXz
xydhatMCHUlLzJUwSpfRQ8ZpyHRefBge3hgYYsiNjWbo1PEZ1HKnJNvM83YU9lIs
HWydEd6hznqEVS9iyzuF1LupeBIxcFwDIz5oZCeaCAMCVytMoLqjgtaShZxA+Cvl
yz7wvk7sYnfnLIJIGZWvf4v/rglXCOqWu3KjetJS4/e6PN9repcZFEDAPpbv9PnG
ZrSEN/MBkic7Mo9g9fa8GcbwoHrNc7rE5LV39zSsXNDQH51xkfbvub/W0EW60gsS
PmZ0rf5Gp8S/jAVWGiQcMN2IK9eV308/Ao4bh2N4NEjxcVQe7BfjxVBtSSgzD/WV
14DvMOGmGsm5r0HBZP6Sm/25BaVXGxDrRIKDKUrenK6hsQfMfZb5xtCwXMKrjpYp
kany/BHJg4ShcRk/BebxNzMlK19CY8Bbnxez2o39Hy+C9Qka1TZquHQNAvB+AbPf
q70wjP/sxD4atyb1FwCpbdBAT2hh8Nc2MoS0wF28Knd5ssaNBydUg5BeVyY6iQqv
REeFDdabsTb7KX5+fde7h0U3Jqs8CMIz69cvUt0zs3cfYO3u0EGzsm93sH7l5b3N
NwA6a/YOS1M5IZqeoLM75oyWwg1uyk16FcbOov8Ynzp87G3KVKXC7AxBiDLaWnGB
eLrNhmd7sYbfqqG1JAy7vuNCD9f++s3CrbvKfXmWF5TmQjC37pCVUjqrtbccGNIR
IGAsvORKNrY8d2A9nb5miQIEag6Z3gZSux42wtDRatqWHR2bOe9wwdA+a2tPf3mk
sIrh9ZwicUaOssuz1cRiGDBNEAzuN4SisyZ67hu49JR5lj+LmS+/Ktf2rgXuLmyA
f3csr/B9Y0iFQtGPaDSMeiyn87f4zkXfa6P7QhizaQWJNPnVdtkeV1hiH/ZjgZY7
j6ucYpfyElHhUrJh4Y7zti12S5AGxiJABnNavWbAfRG1y2e0q5YJUbI6SQKETmgy
W3Wka8vXIhlhLJKOMHgczi+nKOgabJjE0Kl4EUk3zr4rv4ni2lvEmG1hCIw99RuE
NVB1UouX04jC9VTfOn29XHrWdAwH3Qwghl6OUJZ6es3l+URCxQyb3iH4nDvHZo07
7ddjN+GJjCXuWI/SZbLFHQqGi2dqfoP6OSnUhRs2H0fcn5j9ZV259O7QzfqW0ADr
HX1++M8HGNTRU7+l7TpA+75Mk2mMNVuiiFZd9TpWq6ZnvIDskKwys8GgJEf7aqSh
gj2sMyzg6sSI7YGzTBVZm0YPBZXbQMZt0IUMyNnFpkzBLvIK4dwxfkwYSHmUOPMW
ND4RjEU8VWkrJzDazJKcsh9URb/LNFUwGnjcToff6CAgidDJfSbWAwJCMPLF8hUB
jTpt8NbicdbwJrJaZtZ2lWM6aB9zqyxXd8TiVXG3gidLw3tLz6z8xx1t5DtAUmbL
IjNwRoEks3W21zzwMz/3VM8W76H1DOukJUXGnAzy+WTDy7ONjBnh339L0xr9KgrR
QdWVpm7UXHpaYF+NErCjYTHKhu+sdbWBRClC8wwjT10BByfF/72la9uh9cZlhd75
E2HRY75QayqGgPANWB+q3Kk6TfBFglzu5vGYs+rOShEm/1+SlbgMXJAlN1R1wDEM
v2gR5tIJV86m2kABa1WjXu1swkuOo2Z+VjoiLjGI8YaT5mTbJQ3iZ+z7SwCHP8Kb
nnHBpc45nVQBCZazoFO9opTG34PA/b/2je4ofYT/DQ+RSqa6ylfTSrQwFCCGO3I5
C7EqSKlaVwTWip/9QhV2ixyEKM/Sod3A3//R/+lwPLEMYUg/EffE40P5pBl47rZY
2L25H9yZvaIRYLQBhnBU0fzbzN1K/50yqJHeNCdsCH4Bgd7M0ivkxc0p9MMGXj4e
9N4IaauV0Rv4MZsrVXuH+5B4dgckvgSMLtrI1Q/wTAerF5qUtmUv+EsWFumrtlMu
8CIoU21E+h8VPvdaHma9APw/Ooyh2JBbLGqeylXKuooq6Wd4XqSESy10EBZNiSRy
8ZD0SrDPM7zEYK3MEpk2E+etrWmpz56MNXTM6n9rKHD+Up6nnujDyUN89AcijQpV
woMnCDafT0QVacJU46sqjAFmvNJiZzoFUIM0O0wsBlVR9V/T4M/Xpoibq5DTTUzG
dHBZe2ltMvzevBBj2Xt2DylrgZwcQIqMjPN80to5IgKQ726a31WCme/3Gpb4akR2
qb0huWT3YsBJfWLgFk1AGtOK1dX5ngd+3Vlc8qVud992zB+VTiYStLAWcluD/a8L
/0k6ujlhFy21RNMrF0hY9JtpoTo8663n1VLXI/efQsNnedzCRfV5uHjKunP8KS4W
adCe624tp1J9LXc6d9xe7QMu/olTctuTzN02hd00RfoCIDgs5KiQJqDjh2YpzzLd
NE0XtP/THMtaZls6W2JJLmmuGTiyxr0P+jf3O2zPWMrwLEACjKVykvs0vUcu4pt9
ZDdkKE7gINBBfPWZ9ER4a5lAW2Ohyax5E5BFZ+NfoSnd7GC+B4zJkvB40pdN5LeN
Q+jTWx9eOCD1BjLixTK7r+nqJ8FGT2ji+4h6Gc0xeGZoBdPNfX3JVwA4s9PJT5nc
s6v1kz9B8RZe2yrTKKkDYXc8zFW0f5tPVhJgBxtW/WXpyNFWqJ7TntULysZ8WVRy
XfGjN8dcq6p1ljZYdskkLaYJXMiDgMngKoTj9GrjHENIlrg9FgwfmyBZNcFDkig3
lPdaacgLZ8TZuSxguRhjhVRwBGnQxx4G9XeAPT5eFV53LR7hDHiRH5Fsgfq7DhDq
vJl36arHe1oTN/7RWbTRZ54cRf/lcADPfHRleIJBq3E+XAr3tUOVc1N9dmPlFQJu
et3QdtGbdrlUs+jZWaRC1gLKmNlAXUfswzcGszrVgoSInAdCxHAc/XUpDo5Q2Jmr
rhmmfp+Rfi+1H5MOJC1UIZSFql52Mw5v4vtyJD6BEvzh6S/R0q4S0+JLWiexEjAP
bO/smzFxQnkpKfalYBWYT8DyqJnXzPOsySdfCN6dWlukCnFKP0ukEwM1HLfYyq4i
05c66gfxK7BsDZRdYshuvv5kJirkiD7tHHBqWQBPPVGENE949276ybhwxiRdBbNC
aEezQnvd7yiGdo3+z/Jgn1TsEw8VOCy8XvqL5Gqs+VPErJL3dlBjpIBd3YbgYSsb
iTc2SAz56PmlMigauI4rNka6GBacig3EUkCMCxBWodcXwxTpvAkRIL3ccIYuUbKk
pyxhv346fT3ZbLMwTQX4guzUiCavQt+7f8f98cDM6noAbDia9OdiWojaZ8L0zsYG
ncEEkRMVpzfSGbZgeKED/thc9rib3bOqvEwOU0/GvlcFqZgeK2Wd6ePQoGumVQO8
8KHLLTeoIewPrfw7sKXBN9yp3itw05qxcRGx1jwI5pNGuZW9xN6klsrKOmZhi9ng
LQVDwE426AIGN9tLmnNsLF1rxEaLnBwGleh8wf/0J53f9SLYJxClHE/VQRq7vNMq
gFISjtAa6L9DKVrsdcTku5ePX9z43hfGN1GnbVu1Y0M+WyCj05La/hzylqkwI8br
FQG5G7xOCxgQHFcBVlL+8e7aFdsevB8GmxPklof8OxpM1dkhOne/Uw57YPeuUytv
809LbK+Uy1CgPbWyv4pSUk9dRyUW9cg+JkEmvWLZrwqg4AR+sKz6fzuLryl/9yaP
bKBUi0/7+PtuRvsxbCHsATTv7OHUNsCAKJrSu1LaDc6/CUomiiMBTKqTGbMsbdrf
YXtd15krWKr7B5lIQuhiXxNExvI2g+ssdmsA7CkkdwH6dPVs22I4MgnVcNLGlv4P
dVVkz+GwMH/+QCMp38Vq24IqHzYnlhHOCUWPe+7W0uF6eCX6pc8FUzWXf66n01Hd
ekvzd9nR9jB5UkE59NweGPZV1ENQy/HTYuMn+dQTM9EGgJNhVVcF1bdMae/GR29A
BRfHUzfwmOOO3HSd8GQ+y6Jc2PPM1Cy/KveMzYXpNautsP2teB/9k07181zGP6ji
WofY6zjoc64SKlLeNOLxXdFQ0fFEmgu1WiLtnPp4cLkAIi8Klo2cjncq72tuVOuq
LhPOaqvz3QtxCBNFOMzyrQ15yT8SUQSCyaBtZZiLDYNZGE0hZWF3eAvMowRe+F/u
ExeaNP7YPKKUgrxkOBr8G+tfFkNbBGe1riQ3588IJGrVaLK/t7NRPb+ieqG9BAdK
qLInO0Dd56thp3Gt8sC0yVhIYnGoKfOn/8ED7Zf4c9JvdLWsBMHyYpb0x9CRAIMR
SBxqbizkLx4egvWiRL2n1ZQPL7vTAPBgE4WF09i0b0yOIlnWxqHQFvjHsIhDOJMr
mrgeoY/Y0GD7+1b0hAvKvyreywhu28IJRr00BwGsiiDTq6ddjALEtJLlCQIJdPBp
r6JNQZZxktaBiBLNe1PGRD+kV/5BwY+a6uMd74GBWz5Zic8QfLa9LKTtxrYAF++P
3WeyjeReM8ZSEjGvA50T8xHRfPeFgcD96DhZc6yYvZtcBJZ0muw8mnw9uwHUP83O
+Zr/QXFX88UzNJ3wZeCCao9nSSCgMarBqtwisodWU2WIsfAh58Qw9unzmXzTGcjA
IjpDDKRVciYLsYrLn+2DEqfw51iLAQxhEnoYJM6Mdi8VrlzJNOobAEXHF2rOOMnF
c8jd0XhioqxyhnKtE8Oc1Ext8EkcLLR/3D2S/otuK7hF4Su7rGi3b6zSc9m0DEbi
OP9p+0GNviq67LFwWNxerjIj2rnfxcTof/FZvW259B7irzPEyIbtt1B5PI3DMp5a
t7nvhvgBntBOd7RNm/o2crGpbcOgz+UZYljOoeKUVDwKDrBJkdMWlL3mGtVnvHho
5FMp5u0f9Obyx9FREii4/4FDRHTV0/SXHJLrkNlkt1kD4OqQtPl/GYOw6qGOvhlG
TCe3cwV5zrEWVYNWv6ydKJusZBsf4y0eSYHQdsFArgJ4i4oAsbTSMl2tcUSy+PPn
fR+4p5IycdfePqAP0u4h9JfovWEoyGa3wBQPse1ykdwUb4pgEOIyk6faWrIt1fQ5
oXJCB5YCiGtNVxw2BfKCznLxh1U20iXEC46M8mKN9yIrpcpzz0Lfd+sJTgLxaQOu
KnKMCvZoPH4hLGn+d4WfJWSvdIo9OFzSKDD7bCSft2h0YrA+/XcKyr/BtedKIYcM
aPWA1kxBlREJIhZF2B/K+G4lAWCcpTvJrXJT7uuper0MDcDbndt8gHOPDxrgYMUG
uh3xuPfuSyr7GbHjqutlrxNCfy3GTdBbfMvMQxI/6rNcfh7dTX6NQSHXBcq89l3f
Nj9+m0QLOVZe1tn4q+zCvJTMjsMMLyQv5qLEafBfF5rQRKBhmQp7fsJ2O6VXudjs
4/M8WtRHS7te5t0zsSQyGevBVd6dSE4brWPyVqlVHeIlXo6BAuW+zRiAAGQu+IPg
WLZrh6x1ftmEDsDpb+CUx67ApPysSC+Z8wFIeY82RKrGfC1rXQDxk+TNH/RR1uzR
UCKSnjzIPJVIjqF3cqs48/Iz0XJy+sfYwITGFuj+K8Gd+vXjmjn4allsPtJbd4tC
TYq3OSZNNO9smSFQANuAWx7hLW2ivGG5qGxoSJBqN+37j19L8SIWnYpgs4pHPPPb
eK5jyYzUOK7NlC/O5zh57mZMJ9YsKgrVuA/gc92bFI9VcBzfbsBMUh5K0/JtBypZ
VwgxySnZYm0SjjDfesvbcfngzE+hRvZcdrK3QWpv1D7nnOyz4Y47ntcddYFBPHJJ
Kk7NTIVlp9PIulD4/UJjWJz3AUmO7+6d795pPgtm3Q0JCWHs3j1WrNOhmvNz/5/k
SkneQ7A1AfA7qbO58J5E0Lkz+ngaxVo7v/P1vG+wOEWzHqF0L3bBAyEmptfku5s3
qgfHte0qBXp8ODTOIZJo+HryK1MwKAXZnkeZ+TbDHPewczkbzxmEaUWgCxLk4vFn
5beBpX3vwanDewBCiGZZxhaXDZtcDl6Xmem4MalEIe+wB+r4ujgrDlT/zDf2NICD
FH0oxMxWHnrP1GLLCmkkf1d6Ulq8KfEFTl3+eXn62hQ+t4mKBNYoPPaBw7DmcY6N
eDnVMiEReM2aA5QTzXaDg0US0JpAQcISH5jX1jPpxo71mFMeAUb4gzRQEdGTrpDY
uIOKKHUg5vYJ4Z2DbE8YIp8jgoLd3FHtET1oKo6kBEiWFxhaT8t3LBdDzZJtF+VP
sqVab0wdrtSvrd2XYo+TRchDo3pgBxPmRp+oQIMQHIK7ko/ItsBnlrh1ZS9CPGlP
On2K5ol/4wPpcRso2EowNKMJc+ZJz13BpmZrxQe3QqaV5ETacl17DH5t/5mjmaTm
W0SXpWxlmPfejunzCVJtUmUxYwLMtVilSJ3H4pTZ7ccD9H2KAm9+qJ0mLSe8A8h0
+Z7jsdMEMNTaa64lrQgQWZh41B1XyO3LlGgXVH7cplzaQPyM+4qz4bAO24TCXDKl
3waD38qjj5MGopAtG2oIZSz/ZX068dfVfKSuSOJ0zTEQ/MWKjrcnbabqsujfPGcA
cIk0WMTZw/ye13E+pSDh4dE3DE7t0T7XKK9RPNgqJaAnzuCV4zAPtqXMaczLd8cP
f4Xu9DrOU3RUc/fZbPsJhcFr4krzwUVCDhWlMEJ1oUhI0z9HofAzbMQsqP4GAT3L
fR6w2ejvxvMVJEXGDAh8RUhMhEbPIXEra6lylWtN1dMkjr4WxBO58Rf43afqY3Hx
BXjsi2uvt41wcXl2LMlB11J7r29H+QZ0N6BVBUR+/R5qb9aMujeXQqIf7QllGB3W
QxlSwOb5/VZQC7rNsWjeM2R2YUeamZljZKF46VLygYHd3ltk/l4CtST8mw09qvWa
oQ3XkljvfeQEigb6mtA4C/VbPAqdbHvG20/9IrddJIK0PXJYc5Cp8A2ocRwHQuJu
HDcMaOHGVwfBgSqS/8BQRfQZ019U7mubrSdAyWlfG2/oehoZKrdIUJKr8e8fS1ha
NHAHX2uS3ihGM9hCe4hrrTe5yPFK/Nhd0iLNY7QYUuxwrdwvCv+S1PW30r+Lc0Rf
1YX1zRVFHQKWMdMbd9cbhKoeE0dEljUio2N94imJcpEDNsF4EZQAeeIbwlZwS6FB
MqiEjg/fUoDP69U11nFqNI5StX1iZ91DEFAYIsFHaJAZUx9mFJHjwipZbGsI2ac9
NQ2hGjrtlzvIXqXhFeMbmvyysj3Db+S6e5M/yyGw7LilEFE9oGk1BmBRU2Z1mNYr
X7xSbZn/bLdeQyy+tciBvkunawqbSv+0grWg8lGT156al51LG+UXY3PY9gzBI1qu
0lsTHeS3G5WVT2QPanvhfzAh96DUqe+ZePlEUtjW2y6Uf+COmf+NtizC+0SA+Qj8
TGlpOhxodaEmf2E/+QQL7ti75WSB5npo9dFovFEswsFn7Ywr83s0QHRrbfQ6w5MS
LEoHcPBYDBiOIuDRYgF2aMaGAsPf4N6+zwjYwuvzd1Otp/lfS3T+o5nHg4YDhNx9
SnonU6P/mjIWFejfjeMFwaXsdSNF2iQn227FWwGWArzL1N5PeGco0bP72hxJ3p44
IT1tEhlHLJ/AEPztA3UOqhvoeXYc0p0jEUwVbVywmbznVkC4iZXRMxfbK/UaqUHi
lbJd2fU9pQimLqKKG69/EyBLdy+ZrNYog0PZ1XQq7sIJjwPOPknc7hTEBKix3YL6
+KkOLy7vQqPLOcVddLmFIQRBgSfxkVIWCX+l+YgQ92T5HzNGgoCjROGoHW+zBl26
y/103klHYpcaf+XDPBtmDHgsQp+Voto51hyQgigXAbWn30zdLJOAeehJoYIu8lsN
6KXYIQTgjgKLwa5kz8AfjAcg5RuMAeHH74YwBpULZm+DZR/USP0Op59rxv033/gX
dOi5j9iWZAgdJd0ZTL/e7akgiJnX5rVk/n8nv5rtOHeYb0FALZ11K8dKrQY4luQm
555cUVf4IjONkrtaD8lXEyNjYsU47iFPODccC8ceu3Ac0CUQpO9vrM7r8PiwLRC+
FHNelKwqAeVoyDAmg8GsNv9JhwtT8TGXr0QUhr0bPJmNUzEBU28B6ycH8rCZm4ql
iySLXBGgktgycY/ZHJdwN4NJ0RFR6T3EmXb+P6wmV41Di4GneGsKH1XHZ1cNwKQk
B3yzSmYi+mQbgBRhduDGglLW2A9KGUsIu3oWYeMUaHySSohWnexr19Q2rHzdxEO8
A1DlTI4FTOAPdGABgFqL16rB1v0cJGfJZRurRGLGwQc9J3aNoCKk/QtFJTfoN6k2
j1ECbS1whUj3AxLvi0NXBptgQcEWNPsfBXmpr4aExOyUQ7s/XTjCjIQNkoS8BzRd
EVVHQL3VaZOvfisyfqUOtSAj9BS+jCjxHLATYH9Ic5tTgZLM5KzK9sHKyeZcNZ3d
HZ1N03m3J9oV9z4dCsBd0HwlLG15+co4dA9xgDR9uoqqcLGBc+ltISMfDhq355P8
ejDvlMlZv8nf8Dl48EhB9T1l0Usa8PZMvWjygWMtmwiiO/t/p6mbxDVyrnabjtUQ
MtrAQGPA5YifMonOntoClI2DYAWv1pR3XEBT9Bw/9fs+6y/qHFhUYhLh8SEXcVbU
B/lQtN74MnRydW3w+eX2FdaZV46XMq745jj7UF++mWACTvcBdWXd1cjTfWLbaRv+
pyc6zTkNwRC3zEIIx/Uw12PPzCfYtMJc9drJwXxmI4PDzHGeC02xCSQb1DlecgpY
v8H8GFmW40dtb51V8HdohwxPgYPKFTYRZjFXWjmBGWrxWHRNmsf5CFzw5MZFTA+o
4CwVyNoxyzrqQRH5m5h+SJXB9A1+K1pp5NqyZ8Q8cMgm675FbSMK5ImaCglhrGpB
TrO4nApluLnZrsmN4MYcZYPXbcyACsttmDDG9QTz9wikh4HwveEAPnPoHg1Or8Gh
dwtIrvsXxDhhJ3BTnOOKl8W+ip61cpm/cSqPdgJ2Tddy9vsqO8EhNdD08JbLQqCN
OTGls3AgyNm0MPc94PpHcUkKXw8WotSgEk7rShz7Wnvq0alUFOB+ale30F07GTTm
/mhMCZxdqkF0kiRs+zmwpO5SoZFDyCMKfNltfbYvHj2rB/bmqUIXPZKSLqzWSCOC
CZm5/BSGc/ivexYcjymUeTHLiybdBqAZSY51tbjvhskrY2bn7bzV3horI4F1VeIG
vX9XqGG0bbN+lbRbJWLOyTE0jvpHKwdF4VurPDa7hakg7xaFCuo+7Et80i4aJ2Wf
EG0c2Tdco79wBeYMnHj/0QDXkdPJf8jmDjm6ZR+p84rfcp3mQs5hy8oe40fpBgJc
flhdFwrD8VlNYU/tGd89Jf/dghhfDxAQIbexXdPxu++wJGauGcJHmChKUFApiiS3
3qIRbeEfUfY5bGDnmKmnyOTmE+b+hnKnZf7419vPT/6AS+mva4qFeLltYz2n5nPZ
+eJ6COB3VtTiNJa0lhOqPoQLRhrSwaG6VD/A6mXGbAPAu2Nn/wDv5EI8j2Vuroln
6gA0Haxs8J9YAjlr1YXQrDWlCQyUYJoEueaaevTQjQN/ILtR+j56BzLGX0Un2tPk
LPulRn5/RoLN9js/anwxvFt0J6AtkcuMdWBOD5SZ6hubs6DjKlYVcEjZ6GW5NvJQ
/y5CFENi8c6vCAzzG9XBnV22bnxOyPLrgUnRIDg6gJOugfHl+1Kp2kCe6CayF6Hj
3mwLbnLjsxBu58Yf+23Up8KeQBodJkfHeOaEog/gQ/6W9MhVkVJ686JUVHsQbrdZ
cw1V4KuIDm5n+jltrcp+rklxkXH6yUBl1PdiNbaDLX3OX8E6nTcAenJc2g6+Y/t1
4CMe+GGBsQBzbulhcG6XYcYg5V0m/wTOlzS10bexhHnvhEZZbTe7RxuYHozIHn4h
cAzxZ9rqmWsqojTtQ9P7YtQPZ9JRgQMOj6eM6ZL+n2acLH76n+HAhpPyAMduymah
bQ3oGyArBcjtmPM3z82quiOYHhqwGpiNfBv8OwExHqfsLcoXf/vFHcfL5FFyMghj
IbIxQSX4aHXfDuY3FcJWOtcJNlHw1fFEHEOQPV0zWlsjXBok9Yx+i393p9PgueNv
KixIljPxcCVMWi2jaafywrxPrV28IOo+aesHw+XFSYDHY4wedgv511rnyCURNYIi
Yc2TB23LBOcfbNOnE9J7cn1+UgFlA/Y/YeLZde1iK62RtMCX59AH4/5yG7e77SqC
kndsDKfcwKRJ0xHF/xgVPPAgjGf/u4cvAtt6A4QdUoWe6OSPP0UajyE98IstCYrO
VMwLXVCSoF1ysDW651bmBNLGHpmpJh7iNhN9NsyrPA7Wg0Z2Uv1bVUULgj+f87Bh
otZ9ikSGGl1HvIYQAoeTwFQbEoj6T+7h8DK4QYAbt9gXqp79aMhc2ySsBfjOTPDX
kQsFG0R0SJyoqVejxTV/tXhJdj1RcP2GjIMjMS5Ubj0QsYq1HXE3l1hrBz6A8n71
Ocqfva013urwbkLcL8IWC/Q78L5+AmHby7+6wYXjaNETaEI6ZZNz2bh33CXs6F+i
Fpw21w5KtAmInND7ddhq7TFSYccDAv86t2jGG70X6hzq/hYX0Wxe4+gnaUXlpZ8x
l3HG2bSnM/FOmL8O/NLo8C6kVfPmr+68C2nlOHIi2EhYrsGX9+Pn4oMIeD0M8+BO
iLlF0rb/Cwvs1GFmR2tgV+DyixsWDWaX4nvCzYVWM7qpqEMJ5LBhmyh69bPJhaiO
4ErCePhkEMkyN5D+cYx4ToRN86sb6tCCFjmTVABReZ5zpQbKXJZZS79h91H63mDX
/hsgrXooWOLhBDma4KwJ4rFz2ECIWhjPmyPF2jxhdHC7lImZa9bNVnt1cQFtaYUD
ATkV79HqsQpJKv9JeT8MyBlx+wSqqQIhzYQOX0bm47V21yOc23siE3VbeXIJhHQ3
Lk+5rljZjpDJBJJCLUf4B12cGP1lhkXyc1hOAmlNN7XwZc0V6PYASt1Na5u1k2i1
21v5XHduOknojD+TuFZJKKd5nwJVJLXeY90PiAbbJceDETtiBOQKfzbkWY2586BG
sABRLLzWwGEOLfjA8CuvVQ8O6b7Omtv1Y12inn8oQ5Q20ugTg/Wm9GX762k16YqO
2mFaiye3VKQQlRtzeUXgSfISc+QOTuCwkaBeMa0uj8xmaqYyyaiMBvZZVsAnlLeU
JSLE6OLDH6K09nu3zDKLuMQTsaplzBv4Y2L7+WZaBrV4RHv/d4BCIAEZMfk7eeiY
5mmQrygEGariglPkrPhc5CddRVENuyUTr8Vbj72oQurr0WpAvOwsd4jpDJfSDrIZ
uxWe50jkaxmNlnjAuDEEfnvo87aSWvlwT1mVLkKWnrHxffmg4XcuBhmk4IrPHY2e
04Nwo88ZL5ZcdF2ak9TgsiZ6W4kdURaCJ389khBS07jV0QX0F6wIP1uj21T8qBCG
CU6ugd5L70zi4f5WlMsXNvQTAAraqekpef2Mqj2Lef+mSFgs0ZmpkNKaif2GNO7G
NxZeL0YkS7SH3ylXCsT2S1qYZgY1SxP6gTcflHwjlyI4/mtAAiA1nxrlHzpniCqn
K0Y9ZIjXhFFudR4t1tARuQ==
`protect end_protected