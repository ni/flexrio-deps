`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
hVdJHWSfELCmA4ds+csnOQAALbB3ps7EiTSHEDd//nts1r+JQrRE4d3bDPRJpiX2
Sl8d+xAK9BIi4i+3ruAzYvB6kuD7r+gs02Jsvd/1kn7JYK4xBxCjtdDFjVHOTEl1
sSh1oNiYUwLuwR1yKfP+xBhqxD2Dv6pCKhH1NdGilpJQ6cvivGkSunAu0tzP76T0
4x1pB179E7uIeRplfHWX03KzEBF+eVtfgXVp2W1BGjfAe43y1pCvNYZOh1+TY62g
EgAFgbo7pAujZxZy/YSiZjUr2mGp7o83qMXyusx8+rQ41D3X6rxfuP0RiId2pOpC
6oq5Dfkx04a1dk4s8w8cVg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="Sm9DkM+kBxuxXCFA+l3fFkxuSWV4xqRc4Nn7Ji3ukao="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
m2emGBqRy4AuduN4dffN8194qYvc9UXRqiQc56IrQYMiIVQPyh59I8SYabcDdspI
7AFHnvKD5YaF6tQfxWm+mlcmMEk2Y//aUjxeiGGs+RkKgbHitJF/K7nqg1dmKvDg
a/GaBCq4Bqh0EehlN4ntP5HxM4qcvSfh5m/Coe3drc4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uG91daMWA1mGkhgP3oZKMYye3UAomMWgG80HuuXg2E0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1744 )
`protect data_block
c9NqBF2D1wSep1rW7utzHsk2j40aow1MnrccxUTvKej2Q1cyeDDbgAml4eTSXI8z
QYgCADtWi7S8BeChdv4B2VxKcS7CMq/DaQrOy1MKTfQzfAlK0iubmlTkljLy0Rwd
YnZUZ21GCfDuQpqHcw47V6oXFgyZi2iXFPLuL+oCfpc75jGfii2CznkSpcqCFxX5
sXsnFD8mvf0vYphsziTKty3UO+ZJZRotOFGsPdqU6ZOAPcAKKD2nyd6E2S/j13jR
7JKWoDYd5pkJUiEEp8Oj/us6nVuA9FD8EDe8Q+LOsWTmftHA7IlSpOlFX/ZNYK/M
t8129R1pbIxGKJKNEUKMDAC8RLpMBLznZNBVSNlgtmUkgzzjHkU886OEKELzeVwi
+Cq5dcfB+mskM6gIj+YlSpU3+07D5lzpahXmdH8o+4ceMRPw6Adkh/EA7669Ikw0
P/Cr/CbKJUD1mAW+y8Vlo0+m15ZjRte98ZccM54A3EHDvf6BOsRUapF5yKmNAJR9
MNkv4D/Zcxkja+ipr3lWPorBWha5+IBySXw64onHx2zppBV8ADY7mNNlbZZDhmre
RahuhBAL38+21ju235Bxg4eyt4HYHW8GAcX2WL52QIp8s+JI5NLzGiOmd+QMh9ax
a5lxLT16Xz30kZCXpI7Oqcit9A7yIH7LnpcSOex9ahLA+HejI1PzHGvWDaQNyS9v
jd5ERZsCoN8LD1sXLC7N32Z+nfCCoAtlwPJAgud4SqEmdk2T4DhFvCCSCdXTdB2R
GXvf3qCo9KTyZHRoGfPvdNpOvFRn0ekkknMUJG7VCnWjI8A0l9I2N0FZ/KhwVy9U
su3QvM0DRxIrYp0S6bE7qceleVcwZTXZRg3fNwGb+bxcDQ2phY1vNx7ewc6zuOuv
TNlwiuSLl87UYk8je2XpACnbSh4ZN5LFBvkumiZaOBS58t4BJ+EgC9E9vZpvnNcO
xR9wsXlBrkYkFLxXn3ZKkdS0vvVhOt9Xrb4Q+yAct7zXPMRoYEsWBENdwaSRR9t0
L97WfaQmHBiuBkBQ9LIwmB0crfhsuBMc4cLysa7Z/O8JfAEYT2Lz2AIAxEhQtpPN
rMXR8mkQhp8Hi/D7bmVP+RRap1Yvc8mPJi/+n2/gP28vm/ELwha1Yep90UyKsvFR
Nm89RnhmamFyWvwGgbrpbkdm71p8RkFRijN67fUGIjl6ZAsgHugF+d/JGx1zLbnn
eRo+HvjbLiUl5bgx0XBucnTP/XPxd24lItWgMu2LNJhNz38FUstC4i1Qt8O5VJ2D
KQ7i7EfX3eyoU0sc6whQXgEBWIIYbisdPrBXXMkfTHUphJSmz3xsuIciwEUaKeT5
Ig8VaMq5DrmPGa0xDeTPdb+Svm3VsSUh3pCTQScCq90OqS1IczdEBMF9UiMiVrWD
p7CRXsrlwFmhGQp+sYRx1OM6O9GVJXHszGwumU6/wdp2CWRrflHDgM9/88DlzA9H
Me3giULluOKrrOQhtnWSAKkuE+l3T1E3qAHt35K9wuHSCapA00aXPjEbbl3tBobd
+3Hx/XxLP8hlpTqXex2RBLkCWcUSdrhA7cIRtqB56EZYzuWJOLxU4UAv0R6EYaYL
gt4a1pP31bELs55bRO6sir+usW4un6d5Mr+esICgqAVf3Wlkd5P84rdNQxFuLcXe
4uoEkhZ5gskvIOYWTwPBn4UYxVUvtrd7EmR8gH7LmPNJM7vXBsXCGiE5KSpxskwL
YUQU7dPKECM6uVdAgybaojNchSCN+uSHqwQKgH9by/2FGVXOOFuUpUGNk9Zwi7jZ
aI791MvqozfWd9Npjkj1tTsGdghJGSGOj8RbTOAdAjuAqf++Qvxwc6ozRXqH+LYv
iaRO5iQHboURKIwdTmhzbmiGuo4N+lcdr7q1l3jNHRmuXuE6nspzn9bFUAQKdbPi
UIOw8KKLpY1iWAMooacgSwp5YVUrMbdywL07DFVjAfRBtTNcTHy8JA52b4dCXHka
edqZrJbnTj7fCXOOTlFsI1SvaiDORj+61bKfvYP1tYjBSU55Ig8A8z4Qa9lxOiMF
mOd0bCGgFH2fnYwOjshWDBBCLQbESqlZ1r6NztHZSYUqsTdjU0MkBSH+k0WaWE4m
huHs+sJ2n/XP2QVeu0IP9vySF4GT0J8syULdvUyoObDi0bEdHseJVpMvbsvfO7Gn
X5K9YtKRifGmtEHdiASo4qAEQQb+AWuWnjMmFbeUhUEiDaSsrz8F50k3QkzDq+Ev
//BHxToKeVs3ShihPsX8T6+W5jkFtJcGXGys2kiTA2481EEmj2KiEPU9GANsIrvl
PDz4cYk41FUMTuAvs6AvaQ==
`protect end_protected