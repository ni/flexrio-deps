`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aMReDmrPskJscpWYThVKVItA5gecPPZO1R595p0GoIq1TSTG+UxXhmmUXc+VYHJ3
u/C3EW5qePLufxmXxmhmDnr9U8/cYC1zLfk44v/2OPb1TBrTsludEDQZdGNWeV9l
cPUMSIfZ0dHXN7L1M1E2XtgoTWQxf3VDHs7B7lU2y9Rdm/ibz0fWMow7op2nWdD8
gJ4QlNl3f9Oiotp1p8vz9RFzzZOF5gBBslZxcTF5+z4qO2W7+xLByngthWm+exIr
3Pzy8qyUo/m2DDwOz3VJSvSNm7RUq+0/yJNOOz3jr3j7ZyCj5OqT/jDAWjJSMH+i
2402Un+wDMOQxi21JLo3cA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="5R6K2aWI3OdbT2A+sz4o9+2XAInTqB1/cSw5W16RnA4="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
Gm/2BIZF5/H5qen8uQizPH9RftTuEE9mgEOF0SqeOKegtP64CfvEUnIxj/ahmIpA
6xUR2v2l7E5duaLZh39Mc1GYsfqE91NCPU5whLaBPg0UuX4cgTkO4cYbW/7yvcrd
4wavUfwXEp2VSiN7EVxL8RcZTSMSI0Jr/aojiilFqVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="TEmQtJ1Dsm7TOzpJk/CeTSSFx/zKExk04H6I8sT4Meg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24224 )
`protect data_block
nvPqn26PC4XWLLQG0Fq8XsMTlhB4evbpiwGjZroFFLgtNlE6bBjdtwWsB89WW4j7
jNfYbKN4sBv0hDeMH0AAR+8g+TCqoX7yLdIUd7aGwBUZJr6FdDs2wTUxRkXFYNTL
pZPBKDWpw8SI9CeQ0UEeIdXqMzE1QqVpubV6QMzvXo8QpOUnpDqxDoyy3ASjEjDZ
5+OiZbPenKt80e6S3KBYdEmW7lqo+2Nh3IvoQGdK+qMv9fQA4pXtvKOMX2eGDlI2
Y9ucYU8Fj1pLnZj48geLW9V+tIx/nucdCc30xJ2bDjgJ+dwrILxLwEDLZa86eMD6
nLuxW/MxUhTIvZEIYE9Zjts4bKhSkvWK+t+1lSDX2afhSMnzQJm88fSUBY5RNaPg
FQvL0b5JGTMYoV8t+AMTvFp5Uzz9HwgPqptJgJYqKjehzvlsHw7SXZgfxD36REpx
KMPk9PNyl2gFNmSwSnUgUw8vYmA/3MyL8wAFGa0QjqnWuMmeWBp/42w6rcyv1yjs
je/Yptjehf3pF2ThEDjTCxClmSxDOh2CU20TsgaEjVUbCLR+05USGt0CM0Pd48Z0
WS1d5lYFHwbITSeqm2bJazoyZHZLpWyjRb9dZadQmM1D1ZVplFcQ+r9sedBuU/Jl
L7UmsXr/lBU6ZBPHb+3jVJron5KefRkmCthPrqtecAtLFHP+eb2gXoDevF5yiYA4
ce9DkFziwxJV/bMoI4lJWg1x3FNo+vpWWPi/I9lWFSANNeRkW1LJFGsJhz/Gg19i
mvpbksvzdzRzIqxvGH3lfIGQ0dcZSBVsI8TbJd045lubjwWE2FJyUJHOJE0vkIyA
Y2cJueCdkza6E6xKqp2mqWXu//0gg08qa/L55nHwYP4uLDwf/nT3HYtmaN3B7ek1
Z5rrHuKd6bTcWtqpJLG5zMWdbBLj74YSxdPoAWTP1Pai9jigK+F8DQuxr5B/j9Dl
J0wV17bD1YPgU13ZXighJpUg1JujgrSqTFsrP68e7rc75oyibF7mST4cjN+zquUK
vHKpV9uBKgNrjjlFmtmYOhS98JVaugyxB3rU7JY1EZN8o+8bQpXcjtNTvJcldKnc
NmIM7HEkGDuSs95r5TwFA0FBKbx4rJvoU+jpd3vad2pm6duu6/Dnxhgx1SDAKNtU
b7UD7FK2DTcrNwVJ6/gFPbWV8uZs61rRhBiKFsdb2/Jq60dWizMrfLTwRgLdLg3Y
U9BDDLoSWL7VhoC+L8Z1F3xeQFuTsK4XEWbqM3xA/O4oibBWeCIpUGeZCNc7z5oM
/h5ILwdHEDExLXYE/86Eybz4FqaGxLH/s7yIfEQyUu/1A42NMPWN4Th5RThPPa/C
CjjqV5vhDYr6k85QRlM3uMkqQarCIlN7YBPhMTCW3C3F1Xt+pFSaEzfZtuc5KjKo
thFqRHk39xvRG4lwelH0sL8FomrjMjRSL62/TL5kmiPqBSjGacAcqiL9OofNJ9vz
WEEj3nAPS1WiJNy9GCV9hQc65L9EhNFRB4949M5bZIu/T+Drlx86LCwjpvT/+7+3
qyhw5+94ZGm2uG2EnmoKmnwPV+w2WRgjmR68DLcco9tXz0loKFKV5q+MUOGP4VnN
3hD8MomJTYf/yRgv9nOSFa2n6c3wd9pTSQXkpVbLPEKFfNROeO6mAa8Y1GzJ51wZ
cWL+hu1muBE7jZfFIiPX7d3Nhtc+kXQ728JVidJ6s0XtB+Z7WQdGqYBnQutcyH2q
jiyruny7uDXWfVNE+BkNfYMUwpC2HDjrPdOcGQUgENsTM16uL9/KVDYbsAl3Lc1X
L4UPBvM1qv5IXqaImKhLF1bmvQbJmSTqyCdDGWIIU3qB10Eq7+YGkYMfOhcTB8M+
51jABX4YzT6EyBVGhM86AC8/UzLFhe3Mr8bdk2LVDZOovqWLqKpVaZx45o4iePYK
NLF7DE3/fLzLvAZ/UovTEosZaYEtfKifwRV4q6ajQ0cUIKiMpF2yudE3rOheynC8
vSLAMVQZv3N3xwZGDNlWd3cOMqKZaR5yzz+KzPiw2Ej5HKP4DeP4fi/kY4Dbl6NL
vYC2OLPHjpOVzBLKMHOL/1bBGnEIb5jSwPQDQFxkTb3YRTFyrKMHZqSiz4Hp7qa/
C4x4010TfXSDszQ9wYXOOFejU8iK871zIO5kjdrnz5N3M0brA5/K4w4tTMSAJhZD
edb7mZ2pwQoJP+f/lWIvb+cBZ3nyFbFS8BDA4u9k7eYDsY4CJfV8/rKCN65fAkrl
Q8/yT/bqSBFyVk0hThZ1Ra87wukLm2TvN1VnIrws5yXKZDyZIU4YMvyQBMaK8OPt
68OXKSxofRP5Gp85HgKG5+M8Hyf/u4uPwiUlzxqNSKzRj/rR6KgnrjI0hjhH/g8z
rY66RRCNjIkK7XQLqbBHzm8V0GRAAqijRtEySwUSBtnXaGQSTZR3fJk7rlYICT5a
j42h3oKRuvMYpAJGpK5F/4+W9ZR+vN0ivW/ovFTlH3a3jK30/cC4VMDE3XpZrMql
EjRfKuCQMOM/UQkUEz+Vcoapqt/0MP98lGxkoIjZUHorZpiqEBXl87HTgq5Z3ftA
NZ4FpdBjiDt366s+ck76HmrceL5xvKoUeV+jZiRd5RliJowOc9zRTXiqzQ6LYwHs
mE47Z5csyRHtS/b8Il7jJK5pp4+8mB4sQzSVAq4ZKZcQpmqTNq19zL2Sm0UFpL0m
jLu9x7572hqEXA1owOw+QONPByvm3Su0+es5ij9YD7P8oSZ8a8+TBnHHgxPJ12L4
KlYUqxKhlFVLb2ISGHelHCwVYYkEd5Q9tgf88UobNRExDsa3G1TW7Nz6n1CbJFkT
/MgeZxfruiOA5Lmn1AQKvxr5L1qBeEvGbkSL9E+8UDiBxKzVW/YQSz5Um/sV6WC/
EohRA1vUYzGwOkEv7EVmUMHkjR3/Gjg5VPH7kTSH4jF6Z5RK7mN5ILh5aX1rQB98
PP6CXeSGastcBoWw7n/yRMXa0ohFBBOPx7Ek90W03U7XEo3ibIkg0jlEX3UdPnUz
sBVdGSx7HDZNoajrsUJE965KPMqTj0wgRJUPThTCGoJP/1S5vH4xISEZMzOjtZKJ
Zhwej+Oq3vtu6NRPq/ngyeErwLpn4Y1TV0O9hxVczS+ZYtA9CNb/LR1TRU+7d/+e
6dFSU5qVpaSjrJytv6P3GoC19P7RotIA0bgPGLyWpsBuUyVWORPjRZiYW2EUo6zr
RM4qIzHNYi1deMLTgC7dXn56o7dDJE3u0vfvXzJ7sMqQ40LZrjkyGgagT7U/LaNa
UpLc8wO7GMC0u5ewmo608QH/AwwajgM1JpWSVHzRNr92aCw/gRt4QxGAU0NXoD28
NnZh2Hbyn/8GEzXzKnvI34b5MmHdHSF24sYh4ya9x8nssSnp5Xm8AG0gQI0A7Tx0
7cjAE6bIinltKh1DXdve7JXVlvekGXHespmWMS5MiU3J+dMy32vrkQur5rJeVq3u
MXt5k3eugo5U3Sshf4Nn44nz867M5ZJpftBybLnCnVdRsM4jPxNweIJq8rQoUgga
NEPNDhbmip1yeq3YuV/UjobWQADFxgGPq1p2bBR61Kp5Brs5TgZhdAjD4aoFSpis
02paHulqbbpPOnuMyQXj7LAxFIwGcWx1km4BEbToCLvymZnRb9e/5Bc20ACvBgEM
HQwzr3m/A05smokRE2p1x8FBZL1GPJdBd40j+fV93as+pnaan2lZkcGEij+iPY6X
A5J/+PSWEFpaJln+ug38Dp3otyzcxXLz5mTiVz6Xj4BpvhyNugpkxvGiKRFUpp5x
m9uzrsOfEXoXC4KRlQJuZpPo/qUA87QonhDg4k4arNMZW658/5sPRxsLiggUu4Nj
jeJKwGi4arrCGg1elhCzTxLBarYfsc3y6xYaVsFN3+OVjkspud5lUqmT9/77SvbC
mi5l1mgh+M1lfaaIH04j+cjrKVcPhgjLlCO9SgV2sh7ioexERa3w5nKa9/Oo8s1g
DtNcIhZ+O4X7hLZxGFDWsCZCGfbJTib/ssdTUXmAQ0KbJ+0mbPcMeTMokYZpiOqU
Sd6RRsmqJ3hl8x6EUG6xwaY6+a6t0ZiQ6cUYEFZ+tTeBPxGaaSjCYtPlKp4w8FBR
gbvdnYlFf8rJS/JPS1kWHF83zZvwNF/ASzK5R1MSbaMrDwk18rJgbak/OP/aR3pv
boiC7gwQAvaJiM+TNF8GZOAmmjiKaE9uFVLkz8MqQlZ5b0aEnsRwCevuwva1Yovn
2aiRFnAcT4GKF5uzOCrj+MsYA7jLVdjY8yYRf4g2EZewzRpghuOEmUWbdVQmMI9S
FSE9VY4auqip4nysCbfW2huYA/wJQ2v1IbZ8Ct3uXz7Goelhe+3cNYJJ/76ve+Q2
fP23GHWlqkm3rC3cXDBN+jXM43uB//3Wnptcs3VDTMUFPUyYspAvqPhWYzpzxK1q
mUmTB2PkLyDcda2TNxmmgt9ERR9qX9ZjyafxC9yOZ2TrLemsG/vHgT9oOhlyU2rT
QU/bhe8v/t1Es5YK10/VA6XfFGkRrlfM25XGqT5BrEPQW4xZGqbcZejbgRd3wDKI
hU6a3rt+kNIxSc0lzWpv+e/aMWZASJrtYMqxdzChA/lrIFoKz2qq6oNNHgSx77cE
oSWaVg38IdJpOB72/auNdS6Y88SVnJ9UKrnL+Crf7tHfqUsAHylTpcUmOKQdUWoy
NvucoRcqCehZMJuOO4ucRM02zbc2McI3lBdMKNPEqo9eAv4QxHRX2YtTfhDRDnu0
bAykhdEw4yj2IyYyhs3yK6a7xNvDHe4vXyPqn8Vm8ysHoHlKHewFcJ+4pehOdH8G
001kxUCi3o0P8ikrG7V6JmXgbk21jl9XMmqiLhZkrR3IPBl4aQXhGehj0rBD9d+V
1aRNOJFVbo2/pmi42t/abvLFKPlErvwLecIEFJoj4R/TEiZmMuP1wFhGPvG38h53
iSIiI6ZDFcBJzgeQw1p+NK5Gj4lG/ZmUdXh/cLr318Cgb05/wb5jo4GhcMnpFGE9
OkUz3XkOvB5xPN8OOUSnlxPvMnzFoU5FhRtWKiYlK+MPE7HrP/BWrhyrBhT/82++
yqErLbSI5xRyPZxExSC/z3FDTb8WIS8jowgwM6cPVl0oVlQ3yRVNwJ5xFNIr7ICO
4TO67fbnaeSiS55TLlc/jqZmaep0DgSos6N0W8+NkqLouBoY75IEW0GATzRPCzxx
qPzO1psFbDh0MXtsMCoLG2Dj6HbdifgcXA/B39dAufJibm7+1T6IjjxIaLxeI/Dp
6FCKRqrcxJs+oLRBTvmhU7LsgWmn+59yVfwFNrNPZjy6vvUXtQBsyjQGsfrDdU0A
CgdCrA1lLtzcsHmcIqobo1wGJM+4u0NammO1jyU0D/0iZ6VV/hKXHbquaIu8gCkJ
dxBNvxtxAdvVdjLVlqNMs11D69+zupgOyMefzubj13EbjX6LkQrWtxUdPSRZpkrt
gFQKOQW8tmMd0+s5uZV3trM6cxvy8wmN3GyaX7xDN28je4sgeG+dPbTNdt783yMq
/Rp65VUYnnyzF+c6EpI1PVjPPoKqOhWTxJYZa/1fIdck5pFDDR4ji6TrzbH8O7nd
XhYzFvRODFRDJfSp1vXNoyaBuS/6lpHMNuoZmEbNA1CAhZqpMqTZPRILf6Lk5xzk
JePvVNPK1pxu1P7Jt0tUMo8qe7fdppUSCSeRbHHOHlz8b7YvoQey8MsNqT/WV+L2
J9Q/HG8v71IvPQfs91L70GR/dqvAycl7mNuiWjBfgyfiPysCBbDQWoM2IQB4FKSC
qepaab16CCHhfkYmBrTt5ThEpwKm1wPa8wX0bcvGuU8C1aQpidWrTFDWnyXR9Txq
OEmzoa0AZLiDsY1RJMPjjlCJp99pHpnZqvPwEeMo1IGySn5Zs7h/tB2q8BhudfDu
V+xN+/cElY03jurkZLCmTPhxmiFau3gaz66grdyei45bim++U6FMVOgT8qLTEY8K
LAEURn8HhL1ppA+xrA0V4a2IpEyY8wxvUq/2k8WMo8vcYKGtaQeem0kjs6JNLgPI
dHEFEL+qw0y5jXWcJvWwhSSAgJUrrS4td2XaJ3HEsk1QgK4pyBJlv0AjhrzlV20X
O/3WxkUZ6m/QCMZ5dA1QqeOUFuS/wy0p0PmmlvYWF9cOj+9BJ1N50WFZcUQcYS2+
qt6fyaof3mc6Ott67RiCvpNdHFCMQ+DECmLSkNkXfCGtz6US5kmQHFwvGahA+wlL
NuNr4axA0ez6/MsaDxHIAkaGNTd4RG4O3LSmv1aA990eglTn567dCUKgzUoasTUb
9DtdRHvxVDq9htFTgcvcxXRr13PrVplxfaynSmUqH9TVbBNyLa6s8wsU4w13nDtu
uBrFFMakB3/tm3OOrAOR+AhUgubc0sApUYg4/9GIH0rx3xAn3JFnWKFxyeoqmB+m
HQjEUoO5UT+rYrp78kIpUYqT3seXqPwVMGB0Rd6Ec2FPYIhTNGrcRPaoAAoLtquT
r4zGRLT7DWoru0CPsRXCNpLGrcTl8S7b3BA1y4Yy4oxHTnqFY8F5bVgGmBFohWRN
Hc3+KQx2WDGZQYxlernFrDK+u49h/RaFg/wxiY+8ueCPqUy2IExnCunuZ+JL5jMC
3uiP5ftJiUSDz4t5JIhTRVZhikbEA+JCCSfNAXl2AxJ49TYhg0mPY6IZQ00y77TL
iKqJr9vSTF8M7heOv6U6MYaJrbCU4h6aeav5ouSky0jOdVnpSQ26CeWjCfXSQ6g5
yhTi9CUXNOwX0MEQrDkHwV0PdozXWPOpPJN6URcInieX5yDVnm2SthtkN06FXyH4
YsVPAr/PIjAt9pifR01XhXasZf7nYp+92dUh4KG7GF+gR6p3egRKtwxJz79Dr5iI
t2tuZROOMG7kY1qy4n89GZVMWJJn1iJNTN6cI7+P7OaVl46hktu4nQXkfbx1GTep
9Yh8vPG4AdUa2YQ6c/lT0XvaNSectHjrpAx5NoOiwXIyNqhFPrYJTB7z50eBOi0k
Tgqf0L2IfHb2f6puXbuhyPU453mO0Do2Xqg9f/GcR06hb+qRmmYjTt9Fs6vJ1d+8
bFtod3zz/XTCumOfMekPI5YeUR/mDLYEf6Ounq6pvWoE76UzdJkJgcu8To6pu/Oz
9COME4Q47BhzeA1W5D1qOQIpDzrqcecpdfkD/+7C1WwHxHCjJwcWiUJDuKcrNSA2
CDmzo8e1tuwqYXZbwu4vyK20NEL6sW06euj5l2KlhcL0nVzJl96lx6ENNzJ9S94r
uoGpAOphd3f0otPuUqmChJX+8Odyjkc5vJA2oEhbU9pNGp1etWnA0cFRgj/xuLsi
vQjyQ3x2C6LnEETIAQr2CoHfwu4WlaAIg2b1tDUGLEzKnowDfGFIiJyHMJCYDlvK
taNvowEYoo+cQ3ettBP/PLtVraoNtX7fTMBprSUdync6nfAicGXSyPETHHW4HfIO
YS8DozJuDXgCcC+M3O4SdMgptl0GwLiStsqoQTzdAtcUJ8aPVilcc4k+Xj/xN5Js
+vaN/LNh7sfvCb01kCzj4ZzNmDvpLun7mLveE8iqbaE0KQJUPYORVO7Wy4AT/Ydj
aiVGzjYyMz1ppfsqIQKmomicdSqpz4zEQGlAjAfftaoAPGXmFfaI9XJ2lySPan5Y
MGCdq49t75I2IRuA//hXA3wydifkIu48lkM77A9uMwdJICo+MkAZ52aWVb/NaUPF
vLA7Wo1MFbrRgnMxIjB6gmc//1g3qcMfRI+JdYTgdFGvPqNc+a8K9Owq3gj6LFto
1Irx0brMRXxN8i6XRXTOHRcLAOo2BqFN/xkyTkWC6+JAwAKk3gGgleaVtvSGyeEu
8uog/rL086MeetvVyYKanBdDDWgLQZ+PxO5kWbbZjEoIPIJyzaAF1EWT9sNDb9jq
0Rjg4tdVTTLO0X5Xe/J0zd2aIXkrY7l8CVjszxkvSq3NF987G9CxInHYYL9jmM5D
Ia4lx5BpclCNQ7K2chFlIOU0bjHhwfuPNhN/Hr/I1lpCps31RPP9yYHH84Ivtp7z
PEgc9SSA4tAtvV3IHmIJkPm7yPonugbZYNAQoYdTosBRf+WbugQ78ZCCjhgaCDm3
qKwDmfFl/vLZ+gH/Kp4ve4fVFCzkAHrmN7bQUhOKeVI2rM8f/tXe19J+wswTP60Y
nc6NvThRVTnEH7h01LLOJChuQz/E802WhEFxRfofM1dKLMaRVLT58l7QqBSh7Xib
Ao3Jy88Rd6VQHIqL1JWfQQgir4xj7DbnkUxRRN7ky73jMteSy+/vK+r0GwzsZ/8z
6AB7QHmu1gui3zu34dTfLYDYYlprEE587JzkbvGQIWLXPOwi9vkA0vCco6SEI6ry
WgDZoIaicKtvOOnTkrg0DvfxR0zKlozCMPurXzVTlM1ZPE0CP0Kwsfquzr85CZek
Tb0IphoXG8SRwVU2X1HV1YeCDABPmfLpnMV6Al99V/AeBjZjppvmuMha2fCt+mds
I1VFu+sO8jOXpTlRSfHZQnLHgx4lqjwgmZCBbwjaiL9peXrZZT2S0r0qhuJhf2L8
DCUDij27QN6ecfpPJnMbOkFWpvMymJYnif8yHpjvfu4rapLYpCLT3vyiKRUu+oO1
RA5TTAiwkrqdnqRecD7ykCVS54Gib9Vc3d4GxOgKW/gL0JX5BI+gLKiVn2LF8W0T
+r/3RQln8TrBn9/6gBkdeLbj+pGy55tzPMeojcYuB/0AwBKEFBhYHCJJFialjc68
sMZ+ebkNvXwiVlIJz+EFrShC7SeFnE1OBx0ADujlO1Lzht6b+V0bAtsOT0jePmbY
vDN39BYY1NveGr/7S+ZBY1cJarhjWzLdvF3m2aM5QvJNSMwOrI/Oc69XakRZtXnx
vFwf1i6YfgvFYJz4s7YJZ4+7mGC1oRvm2bv/4p542QXmDHEHe5qa6mO3pTd1/gqk
Zc+bcHxnB84oex3PrEpaOZzCil0yIoAlZsxYT33RQC6csQLPpuBZvbcSAlo4pEfx
g+Dcwinv7TGrTOzzq90ZK2NIKzEgaIWKIcLcjuKlLs0QYjsfp+Viw3xy5YpqpAUs
IHpzDsmqlX1nFcdp4YOCs2gzrAlxF2m7w9h4RA/AMwBjyN5A/23ALaTaup8CIAmU
fPCzs0n/Z9Bi4xcfpnuy9qMMzJagFptoTXZM0NbZ0J9tveoV3I98P2wp7eoaiJAW
lRjZlC2bEWQITNlTjApy6xlv3/y4k7WmLqojSpC+s8bI/gMcyqy7YLs31LxkrWBz
flyHNBiqN0M6H0ghoQARAZ96ZW6HKoHS7GkyX3bEMVhWMtDXCbMP6OpXs8b+yjxa
xzBlPJ+yxBhE9rGk3fci+DcLbEE3Z6cDfJTwXsRAxTtD8l59H/ovxNRwAgwSu8Af
MI44z1n28Pu+L5KmGb8E+DugesIP11WTWUC85AqsdUzw8FBz4hychE/P5ZO4ZE8h
iCzXpUgl5380HT7RLQwsmhWtXoVhPEZ/8682DS6jovFQv5b1U5isnYYTkh6Yv0Nj
YWNLC/A3fMhPj7rySbuon4N7dV7+gjXvunam4csdxTpoatUkzk11E7u6hSpNwtOs
S65T42gxM/bMgoLhh1EIyi2QXUuYV7aolBnKhhSQ8XVRKNQvHEXrhvamnJnL+vW9
PLz4bX8nGYMSZfIsvaNBaj4VhINpujfJHsg+xkRLKfyZ3xDJwiNQpxDjtEQmAQsz
VCiCQ+2suzQgg5YJCL20UAn0alAlYjZj0uz3HZT1Y4HnfZYzuZz2gASZjNbbmh63
enqMNlXjogtaXfy3fXwaBvbLpCgKVleymWDRPahwf3U7sBSDTdjIhX/x1DCdN/wL
BtgqFqg6KyHaJvrKn3thtYZHbKgv5EkYsklLG+XAsYCDEEiyX7d5peJIrXR3qlfK
SZKuS37TVMgWeXFgNQ+UeLgCKTFcOLCndTM8nh4aEOPR6MfXUOjAjw5WCHEGqR5K
j56fgE9ih+b5h4nQYgs7OfUTXi0NI357k9RsyadX3ewsz8urJXhUvfRoebVLt139
mQMnlhfADZx1XHWEFbTYbOD5E/PG0TNCn3U1gF9zgHvpcimMh0h/Mk2zuxZMOJzG
jZVboPMWWGadd0WLaocIN80G8URKTR/P7YQPfDXCPDFFxrvkb18CtZo3Xw8PplAS
BD2CcpkFqSFNkM+jn85XAV2sBZrZbqS/P30bp71n/NHgwQ/xOdQDbN5vXb4s5f1+
tSx6guhwWp0zJejcP2Hc8kE0oNDVwhLfnNAS4GgZwYS8NWsRKnIQ3qb3hUpsPaVX
hgn+AkwaFafCSan8Jl9CRnRLD5gP/x9fMuK+6GV/SoBa0/zt1ZN9tQqrE3TL3wLl
tLqWs1wvD+3FyEPjKdkW7z0sczIqPOU2/XA1JnSdW6dkJG+UKmixKb79VmnkHixD
X//LHuo3DRpr3uIzvMf8dh6Idc2D8zLZ4oMQI13Hcii9djGUTQ3lsMjn/zJAEs9f
68dSfMks37v3LBRZAT5Pbuf7i51kiweUc7/SEuBWbaThsgrud7xjC/HCxeFi/XZP
S5U51K3ODA0FENc7/tecOzO5UyK9FQmjiOb3ylEF45Uka9H6PG8K4GrG8/4x+24P
kYU6CF3BWDJgSlUi8wbincLfFqTqgR9GfYLKtkRfClZ/8N2XEry5L+eXFs38MAs5
UAf96ZdynYru+Wziw7zx0LEXQ7iyAWk7N1EAnwwWkIKYOEEI26M2qsSs8vwwgUgm
PeccLnUAT0K4WSpf1l9BEb21loDu6kxjq9SRfjYioEWuXltFiYs5+6GdTYGlFEYm
oBgb0xMsQ3CNY9xxvxRqhc6qg3Zj5RjOH6Y0G+Za3RbERObc32Djl8wuekywLkMa
JdpIQptyBQXCS0Xz9TRsgwV0QFxTcrmwtLkY0hDbjNzCOgJCI0guCH3nyLkdkeWc
tXhimy52mjJs0QzCWXTpxqaORKJ+0bGAtFeBS/F+cgXLvTtplh1Pm2g0WhUWkx7P
ulC6DPMiNApVJossAwjzQUWF88ipIWFEOAgI8VeSQNHHyra74rsMzPi+H/rhGOR3
ldvMD/GT1BEEt9GUm/QyxxAgitrUtbrAdEcdz79E+cCRN8Wr+FzFSQp/arMwBvki
O7N0svn6QU/NjHTKDD4CsLlOBXB0aeU3gg6UDbj6BOvVuHRLHOKwZ6cfB6jyq11f
d33pCKqa9Drcgn6aKaDUTLQkMCzqKtwAZJWF8JQjY6oTt5upvL6zxPfpjLivXl0Z
FciZlAC0pKk9EJ6N4tXI2F9iX4mKdcDNJfv2nv0flVGJ7vi+/67R9oRqgrFa5c6a
Np3y1Jt/P67Gu9duivqcnYuioAvBBsFMMP+W7S56ppVv3/IkV6fPIRfxqgMOKRVP
04d1H86bjF+QpTVW7g+ONd34cRWhhO79UMe5l/yWRXB7gtPb8OC1Pix9dGY4U5zs
ynyUSYEUBPBrXwQxd1YOgHL/Gde3dTkt5K7gK76Z/T0gHrEBTKt3HBWn8y6Yn32K
8pnFAHHprB9H/7W1ap1KLrWOZaFR2JHSR++YPfVgRyKk6fEPkA7YogQmj9/Gd61R
VwkzSmB2PAfkXOCJnicIR5wpOxL9HVxJpqN16o4V4nby1JozH8sbiSrJhHKphQ33
vdk7gnL3x44sgFgYhr90Eu8Z7GKVPEncpExCh7ULJEcE2AM+D/TruMbB7W+grsjh
p5UMu45cP9Ektz/v0CxbSLolCiNfqsg7A2fQtxpdJeZyyQe7Rw6kpX3WeZ7B6x/h
OEMNuyv2j7cuUDgwsg7aOL0wHHzPbLDmvx0OLmNjExCUX7oxeTvg3qQ2McTqymAy
gWMO39Y2gtqKNcUtBOB6Y0+0m1dsg7xUF9pl0DkCD2HGqxrGR9ZFjocPLdaq4H8v
qSifnq67ZEUWHqF4MNoU6Xl92sceiV8nN/Cr4QWzaT018FEPr1sGTREg+xV4ykJY
hz+cDRXUVSt9mG1w9zg3N+SvEJsQbIQYzC+vZS0pMr4RaLisg9v+mrdbgPoTuZCG
B5MTwr7gUEeSkqfYw9gRYgATbgpXiCn36tTT9IGTMln1/x0JQ9Y4FVP28sZqRX7x
NUi/yNV1tjtvqqhqMnEKqRQoZFoxMYZfNlaXBRf+eVDr4MxHF+264Yh2RGyOmrQe
x19bjFN+wMarg3YkmDV81bWOVL1gKZEltQugiFoQwI39+5kFx64jvBHiDCbYc/bV
hh/lmKGgem7Qb/w1qex67OfLvDrNH/psSMoYDnfbA/ulUNtqCTlLEaK2WWpARbQ2
Ttg4ZX7QZ8HmdkPB+MynovDCED+3hEt5Jk4sunLo2rveFlxOPHmBL2eapRSLCuUD
HT4cK/j2nbcP0JWAr1097JpgQO6D6fd3vlXSE9DEP40bMSRrRlzjxCZ/njc1c7sI
5/pS2pjJ3n+PGhxOko5vOyGJGWf3gqE1SlRgUN8kht6WGXvIQ1xveiXV7HiL/r6s
tHqGnAUgZLPot2/a/txfaKYyGu1YXC0RLelej4QewuuheL4j2ni+cjRabDl3P9pk
rdPz1LJvJVFsu2L+pT2AzPPOQH1cdJ1VnaN26gu8i7si6fIv9DPh6S1nzW4DWhSQ
qdf3T/RpFLg9a2+kTp1/0YFFOVtr07sRW1IHZ+4NzwVdjNpKHfnp4QM3i/XPXLQJ
wvYJjm7OUyIpfLCf6eZzi4NW4h+uZNHlILq4ByjLpuOkxbxKSfX25KAtuwnAG4ql
a2apPiun+nPTY4LwyUrNmiYmrswbvHjTmqIQJ8YyTKl8fH9VQBsx9tm98KwrY5ac
+6fo64NGN1KfGsfctkH2LJKDhQYlMcX/qOkPo6du2Uf6LpFFUtyhIyrSPN1Qlpo9
9eA0Nu0flK5GDEHEQi22AFdf/Zpxk6Alv/JksiWhxXSkZXlLyAIHB+2sgLfpj/WP
APWiDcfGpXWG6TuDrF0sHkFYKn8+Nvb6HduVpxtW5Kp/D15e51HZqYBO4XmfpTRy
/5cxZJq0+6uAewqFdvWMn+tPphXihfKp4TgfTpScpmXMusP90Zulh2sR5cPvB5Bd
7KdeuB4WAfJTJb9DtgwtHp59vXySzBAe0APqBiKmsLebeZnTv6L1fAn/PfO3shlZ
Trc3a6Jaw1FUsxtmAd2hNzPO4LuQwTzZaPxdUVK0m9oOveEtW9nnWBGbg73ToeDt
UOCxS+TVJXNW46yoaSpsFN7NK/tGZO4vBlbDMY/DRoAuxtNHCLnUHp6KQiRJlKcL
fqtJVBUBwjTJXCg4TyizQl5chqoL6Yy2iotx0YewweTsgmxeLtbP5IDJtlQY0rgX
u4vu6OxsxIzYULj9SslO3Yi8HMKeuQm8faycFpNOAbTn7h7/1GCnmqUwjPoL3ptu
DMfpTboqhs6FyXdNuISzuK5EWyEZ2gAgfgZcfjzoRXf20C9AL6RTDqN+SG9Il5zQ
czrNiMp3GmUMkEap1n3DJvTBo+j80KUsHglMK98KXwJjxyr6vbrqy45N7mpGYMh7
+fSiArsQmwH3munRkNJzGDVBhX2GKoRsW22C75h0sK54ShF1EWqs2+74C4iHA1f5
gZFBwiO9/dpmRBJQ2xyawcJUwvk+AWvhIsNx1Op4uUrraJxKXU5RtCC8MHOphIPE
0SoW8O9awAaFQydTZd+z6H/lsMdL8Q+aDEGOrBlZnMvAXI+ynHI5gnqDX1414W2C
GQKsbVbjlrZfWUriJc3/wVjImV28+S3j5Eabe9G4fMPAJMMmDb3Bd0H/XH4ZIgLb
hm9hcbN9JkJs++gE4DRrOaM//a/gTLlf3afs/uWdZplTz9T/9+EoQ38lqVPFQzkz
KyHojZLNS8u1VcLMQMIkChUELPcbf5Fc2WU6hlXxQ1ZK8FaBYqr9FpwrQvHz0QkR
2v3Z7vzm0h/ISaDrhh7i7POoSZMKMcgurM0GQn2vd4D8ZGEUunIdiJLFfKOtw/m2
cCgQUz6Bz4+ScL5tUewNuoe94qyGe3FPqbs5GHlWr61BRJuQy0ThITd32jr4Dj9Z
qCfSStfOgLKDhIinsWE4/0c0E65YdCItal4XMtG7O6Uk6tRP7bSQ2b7DOPl+Rul2
JzSVNpoO4q/rb3uOsiJ+RI3eZSxS3TA8XHnHlEwXOOdj52Ri+xVq9NB/iW1uCq+A
pj3wVs9vhBeerAPU5QMs0eqsyLbQTT3ruxi0F2h6wl19ViS/NILTeOTKFpK7toVn
nbgG4cVw3pWPLBUtv9YG+T1IwrIlHvJ4i9izM26+5aBC35YwhOqn1YQkkL1vkWSS
dq1JM5TBAOqj3P/xacaGntDuK1bKF9T3PpNzA+OR7/w/5w+u4RTaBh/K0r2FxUub
S5re37YVEnCb4OoEwlHTaLpleC9Fi8jBhgk57HSIKHqqAI7vmk8JTXWP0gUe8M0p
PNGRhRB1DoCpiJh6hG3ybjEcd6QubD/VttIl29uUXzWYL+uqzvua4GSvdojkAqO0
QNX86fzxEA8SAmSFp2lBuAYbA27A9Lk8gfmflkGNBK6T8+D1EWmxFwEEVvCm1Wps
1Ixkgs6BQzsz13c+wRUZigBX3HABkqIIuCdjwi7P5Dt4bYUCy6n6aWYDU2+h5PYo
QumJvZRp0f3XeW8xaVlR+l/d8bASIympEPB1IJyrCWeVle3QYbsMx745VQvaC9uJ
2HtWprWnv3lHQowEhUzKV3rv5eVQY8igLdSmQY2OBdKnwutNs1U0bkZlOKETGVLj
w5Y1QCmbID0UMrlIq7ppi6Npl/Eq+jucKdDD0pQ99+9kFzQDmE0Z3AmlkHRLX6Cf
tMmq5fxAC8kyAkpoIxjRMYaix57JDAA7GKeotd6/NedYE0CjCtQ7RU+1LRBwb0kZ
wC+1UyOX6bzeNwWpHW8+SrpiwKM7V/LJ4J265UaMHqzaW6W1+cJaFVzb6BypXRPV
cBbfN+FV1IiD7br63mcaY3VacSUox3c3MONWqkuMnkDCogpuZnEHt4HLBlwmFvKD
NGxzkeBI6m83EreoxRRoMI42t2NUzwM3umL1hctqZW7ULDLKEN/KdZx13GuxKgaa
N2Ri/GDMw78fJ6afr40oemfTOQgaHCNow1Q1qEfWy7xdl/4vFri+UCYhVcGk335V
QFo6tsL3hN1Tfsovi7fd/m1gpqnw6xsDbCgY/aRCqq26KvE/UY2ptEuEFkwh6Pxr
iCKpX/rsvOmWtNfMA2nTzM7cuFEDGsQaQ+RKY9iVSu6HdXhjAZnYHoW5R1JG5cu+
KKbD/dWMUuJ1SxSju5zgXp6ie2IYFNf3AAq0A0KBAkXht+xEfiRCX4/WpQ2+uys7
9JYP//d+4bRbadm/vLXuDapAomkwZkRyUK4pTPk70a8g5/wAYKWSB2BACTHoqZWR
5uY/8NgxwWBGOOJvQeLc6nna/WwD6/GFf1IjHHK9kG9nFVYzwHRuDHQP0ueUYBMX
LuZIQ9RkklSB7ltxN3b9ToJsi6CT2qjVwTq///Uzenkzqd4PT3xea144Glr3PPOo
P0JQISjEmMHI7dw65lzn4Fp+h7yoIpy1NS4PI9m6zXQDPKLplsLF7wqxxyJcJSOg
luPYe+0zN4XaIp2eWQ2aIX+HNdMCgGPGiXGwjjuChhiCVbDFyFDtGnL/PffYDTSi
USUJvMF2912mENW8XJK6G78NILHaNyKBr+1A42OdQw2rdJT/rvtq+Naty/hPc+WP
bGPBCXgoW5E72/eEvt1uz6vmDAqMmDUTCwWn1cjsiVWy1Hf1GwcMLWJIZ0Kldz28
PgTMYO8fw6TffJZSZKcgfl6HDaPevxT5GDOJlpMPNUI5PNn9rFV1vWPOcnQl9JIO
bKcButSX5O4bYQvP+Dp22tDQ9EftaoI9huqf13N5HzRJh7VOnEsivPoSDjkMCmDo
UiuCqCWmvkpfjP6k86q8LLf79JyBCzyBOh4geMwF9DknmRVA+30MaKzcruLpLVLg
RTKtUV/Zy3czF5flZwA3nITcUuw+0GAqqLAYM+QKUCvkGw3zoWehcVoVMABXO7mN
oR1AB9jBEzlg0f41snRW5kbyjEdqHDQTZF5HFLBbWXpgQLl0AM6ydFV9ebaW/56y
CUqlSoofav7b1ayE3ah0ryxW17H89/rKY7NGer8E4Ej4c1XpoZ/VYeKmfaZOCq/0
TcmWlYnL2Wr93O0/nh1ITXmmxOyKYji7MlRREppBkaT0fRqtt2889RjTGJj+c0cg
uxEYhg3FCD+v17tRrk8hHyz/7cczUmtC2xXrHIgIhEc7crlyH2ggOBSjt/Cq7dWb
nRpSv6blBOw4moaeHPa2vfo50stM81Dm/4Yd9onerg/EoRjRTf8FkQGY/ScBAIMd
fj6wN0/ZAnCNnWM0WwD3/bKGcxt+CyYNRUVP+3TwlGNx8+3YH9znaPcVtAQQIBZ9
/EjHb/vNMVp+d18T/U0b8Pb293Hfj4iw16cUMfXYs/o4SWu31sXRIfDFy2NHlJdb
xk+rgTR9t9u0PYSrwXZoTfLsOF1Sv669o6BMpeB/d2m5nBrv8q7Ah1+7TJUbRoqA
e0XqOTHnD71f2+x4a4FSp6yk/siVWALNqNzBAve6QBe5J2oAEgGdVA5W3IQme86y
Jevy/FSSwlIzYlhm4FglWCpE+LVgHUgXd1XS9pcT7gBYDeXh13jO3aWw7RfzVPhk
+HUvqgmZ7Lm0I6xv/Nl/cFZswxShANLRaB6c0cWPjxdw07oJUduWOd9VemzdoO5r
F8h5EUhEOteOncvQFu8vFFuE0I2o3FauVgQahdpl/Tb3biLcSYkmXNRww/ZS4ENP
mFpOxVZoZObA+d26QNgBKXaxM1cKkFNU2n1sYtSf60lJSDCkodsx6+dUYNWA7zY9
X/zolRT1uPaBIvipQPymov8CFYPNOr7XFTqH038PSeNnw8Z3sHJoMF+Onob0Htto
YfA3+bLJxtmfrVcveOayuIhlkxTdEG4hVyrAEpw5zsTOreiCYFMCPVGvgL6luKBv
NIB6sx1w2NlgdyBqPU2DVshhgWEf2ppXbPPguVpilg2mphy75ZdqhYRED7ww+lBm
qsNJ/wfvcRP+DeTKOo0MQO4r9nDDDLnVNm7e4R/LCK3woNDJIHWb92OrTeX5tRZ+
sa0ZYRcr4DMLWv3ya5cLLzb9am9AVSU8QRJzJoqTtjXEXgYgHjfXwuENehXChkJ7
RQ8SrKwDKMY25EfDFJwY8PExXbYODiBhSx9o2Bvga02h4N8SZ0/G5yOCZlgC9s++
gB340Y/EZMZ/8gcZLCIkeDzAp3S4G6OMSqKtvsnJAYeSTlJMV1fyKOcO9Fq5PTct
aBaA7q5lgMj2VBZLvgvskRCdFByP42OcXAuuSLKYfkRFw6X1G0oON2CW5AVI7jUW
wPrUnv0M+38RvVclFVDzY4sRtXuN9mwhorEvmEbGekV6E3w+z5Y3WdqMQEqdrvE7
qI2J778KVXgu6XbiIWhlOhgpC8P1akUhA9bk0wmVhvPH9LN9Vk8ZqcTZbFk3Qnne
oiyzJ4qeawwyPDX+SwJ/1Ba+cG/japmc4X9xOpAy5a7mHTBihgjMRcz0HhZ1pUwt
aEVz2roQrf6ARgDDwHKPhH2kmQjg7kYt/mfiOfBRV8i8nWCiCOhaNf9wuKrsdJ/A
kBYQ5zfAZ4NuBBMqB3Jz7hzBc1ihDWcPLcKNvpeU/qW2wUmuq3P4Clh+BdTokpFA
SXZioSOyeIpK+k+Wr4sNCn6JgOTd5PULHV3Fsxp26WkkEmwfm+fBHo1jF0NfFsyR
8oPIULdDd53VQtILxWeaj28xypGgglNm6+eKFnbm9V5VklC3i69dKrYL2MT337ck
kCPbjrCym6jwQ9rmrZFPb5lK96AGU53BbZXP+F11uRy11BLjJW+BKe85HvChNTfy
ER5u7rcQoJWhfqw8Zx6PtmePmssiIPxjsYni7Yp0ki7dVWU9uGtlN44g9GnDiR2w
3Z9fc2GvWHN2cxMAhSogqS/KexaMmBrovujr4Wyaf1dB8SNqcsutTO/Zrf6sMku4
tO0X2YZJoLfroA8Wc79AGRPNFUMBtAthdGi5Ck9RGL/jM52ELwQIcmDZ9ZAqaTJu
CspZrYNSoGnhNnkKI7ann9Rzme6dcQUe2Cn8iUcH23GKs9gQQHZKVY8291jyOb82
L6oCfJJSh8OLoPch/ctA0JcAJrl+24jCsObUbnqRDPMndKNFxKNE/PBfIveUwOkM
KXq6/Nyq/rvMi6ZYNUE/HZi+u+CapnxtmH5Je4Qwgd0aN529qGM4vcoJFYK34l/7
BkPj70zpWnXp9T/ojtq+r8GzOuwwJg1JHylpDbmbfFVN6YNLw1H0xxjj6TAunfmI
3lipDhUXP4T2RDYb0yfBJPsGyjRYrRENma/c2jvpFyunAy4sMOfLb8UIXvQXLb6d
ICOz1L5FQfhAAM7L3wTW6MguHHkDJHnu3K6Br9o80ZeaQAs0HOhRsSwg6IPWAjhu
QVishUKtbZlylhliPBTfsCb2fSXTORpIxPyKFbqmryq1r6qi2xi6dcJcEj3WxSnz
g8OXKeXre+kHexos4hglPSjicPrpwu1Hnl2pBHrxMpVeB5VzhjZNLuhsoL2UAK4G
wBFwZTakmKiQt3y420CIRruIVRoV9UDNjgjfohPxW7gAwuv6NX0PtcGqubxXXs1J
wwzz1/7J2gORE3hySS1hM0ibrMMeTYMxoknhW9NcZOwyepkYF5dDFHh16TpwDCcx
rxm2HugwC77kFtu9x2nUcpl4W0Gf/qFp/JcBaymkHLH9JXVuIDjHiA5aGG2o7d/Q
Kjpoq+F9HFOBE9iQfpb1ims9C6lc0ePeDg7fCPRa4tgZBzL6+rlp9tn/9R4iRIka
RcBBkFLqwJDWuSalosxraPu7XZaC7blK3e9y9nPLEExN/VuZf3Afs/4wTJM4Uhdi
1iWp21jgeJTe2lurHsw8s8P+Ag3Y0v4lfe4cgD2zePZxiTsrhlRfzVU7I4O82LK0
ipR+6uQavzhuP4JlkTYCKmHta+0rlqeHp26dkYhT9BRlewNiSC/CXNjE6960fYTa
1aNyRZ/iTWvYo7cCBZ555AiETPe71Qgruhj0k4NNYleVQAfeW4Cy4QfghwmI49u8
3JIt2U8ou8YNZjhc+A0aRFmgEfhE7kMksafEcOBW5tzBjZUM44MwT5sqWEJDTB6l
ffmepR2XO/JagcvaMmzw6+aIXW89SaS+NcZX/zBfkj4LN1eyXKu0pyPdtwEKMjZY
F5Ohf0zzblTvxxO5w/tiGmZ6HnpVQ+TKnWkqt0LUO3aj8PSb7BYw9yXCxMBg3cTt
obSkA62W5urragj/6YZRTvoZssQyjVxgk5uxCwvOBFn6doOn6/zmqtdBKuLuHHgo
tQ347+JNHU8F07RmFQXD6eCkn0WFMQzK/YInjF7+5uQsks5atnXAqf9MsvzHbL9l
i6XgGQJIGwmQFeCJrDja7xSbLDBV6OtzelC21vC+ISlB9zB5Tz4IQCooLfea5Jjq
T0U/b2+u3uG2ey+zSEtqqRSfGKj5mX+8j4kK85RJIC9d6qL/pmog0mZYYp403Iom
lGOnj3vzDUQ26/Y2i6u8vDutsI7rddhsENfzpBP3f9di8ytfOKVWu5h9y2PFF0ji
Etcy8PZinn8AT9+ZLTuobO3ADWHgBLVBBBmknoADJPwddqouyForAKSFY5WSjkQV
YzZeUYl/o/NevDxXHU84r3vHVITrL618gK0KstOkttwFWB+rCn0p6Pd24YfwX6RD
HUnFvwLHjnKQvVEJjtPU2fLx404IU/nCihszpR9u5z/MLeDzNqKqkqSw6t8b0IYQ
y2cOTIyp2htY/+7tbRv+zB07ttyGxcu6kJOCGZugyu3/IB/cTbYOaZ7kDsuqEaQi
Ghjejo2hs+fNX2R4gv1DviMDXkBoAtlhqzNkZg4YvkpOD/Eadv812O0zyD3TE2S8
tWWv9n4OSDQiWvLkwTzmFlOU/c061pCJQR8U14lIqlUXqa0tP0MoF16gzBIIbqo7
D50KC5HE+upZo7b6cRpyD+PU2btV3G7M63k46bQFzPGdVtwS574R2aGfZHzpQgpv
hKOs+oZwvOO9EE3TzcP0hVh97lPhM8LtSf+cvwXyaNV0lBKyqHxlG5CSWGg59XUY
R0Mh/GoA4y7g+pXTVDD6hMKWFrZptHoSvw8h2Buduxg55NV5mkVoyfc0GomPgqJi
vJ//QvFVHDLUy4ozgEavAC90WAnGy9k8UjoLXpzLsi+sBb7hy8lue3aPqsOkWZmj
W0kUMFAYFz7IgVXvuKwooHhHGNoNOYORJ61Ig74SjZ4+U54AogzZAEjWFF4fPS0u
ftyURQtItPsUOBYrdzcDjpWiXYSs0S4qg4mAXvhlbYpYdCM8IVQkc4J2IWB324XU
tvZh3MDk8K0kOGLMXP24HjN24rcxVt7D3rEDH1jFcN77FK/VV+NPV9IN0NXVYUp7
Qw6TRa86EWtkcYlJSeV6akMPUef+S0to6dXOMP8cXJ7pL0Rb3Ztz9L3FyJau/mMY
HTTFampQiU1DnCG/X6W2rhj7h2AZVX0Xu8WadqwPAXshcUVBvGUCen7vt6N9J0nG
+xi3JSn5R3jeZ/K9y+vgbaUfsOiTwo5KV4/z4vZPYDTKDgmKZvGAy+hcGqJvj0ke
cS6apcs9JaoGB6z5x2RNom+D/TdxhFb1zAGCCLRXqt/y7AYw17FTy91DEjK0+lOX
R2MAMBKHVdXygArNfsRc6iNS2cLy4UjOjjp6Wpiw9tDbqKZAmM8nEDWhvJ/DJWvb
5CTrURufWE+vbdy+2il1op4T6CpMSDEm7aFkIxDbYZJntcUiYUhOPE8ctDyaRcAn
jI9yIUn6pbYLjJSnOqBqivc9Hz0X45EZ5B+5T/cselzn79Xp40col8EwlfRJZjim
4kWMoe0o0EPNZAk/P2JgIFVXr2nGFZC02A+jcYX58S/WsFcYQXaUy1eQyyXBo97O
Nl0J+jF1xs+XpSUcsp1oFo5A0M6rMU2PhKmPu8m+nHmVwmwhb/0la/G9jmoSMGaP
AxfjZYQI3pWPjhWtnO1i3usJX9n99j7P7AN7DIEeaV68JrbyHbenwxTsa7wxegi+
m0yyK21Hkf7sm9KX1irRzG4lB8sEsWFHxXo+pcQqJ5Oi5TJSkv78+MzcLlHTo+1K
dNTvIvSr/PGu7pSqtWXIOIPsy9emfzwLTU9xxfnAcUTOYkKNKXyxfi+3pANCvXeu
T7l/qc2Ex5e3nOIq6CvSCIItRhoS4lCOF0gZ8roONNuRlZYc3j6ijUepuMuSj/AV
k1sV/hMQeAyQSPv9tKsvwvLVvBN0SUX9LgPteCgdv9hdrpjLWfrWTRFLNXX6mmMP
vhjDtT0jJv47r6DLbDvdjbX6sGpS+vFgLnBO06Lgo7/UT9d2Ey+ybFHXZlCpM0yW
bBUt9yrRuzvpRV9vREgLrk4m8tT66RtX/+It2VQttHbUe1tWmTG+3yJ+kJLX3HQt
9lnd36FThwzshselqYOKvukaDHzPOFnXm3iP9yWgWedxXv60VFRYC4oDWGLm7EUs
+hIRyV0cnoC8yjxxn0ZU+8mhYcH//qr4SW8FDZheBIJhGTvyLNiQ3P+9tvCl/Syn
rg0pF9C1kYsqMDROSt4CTtUXzDuxLjtpxHA7c8D2oHI6DrRMB3+q2bgn+QiU3Nlc
UiqAW5F9mn8mT3U0p639UqFAkUZF5TjU06fe56E6Fw5AVegVdVMrtWby6ft6drI5
UEX5udQA1Mu3vHByRDMSpJ5CiGUWEiM+z+FNwPUbEmz2+GW6KpEiID0UmYJ0FjtC
uZuON2Qe61BTpkQATNz8Xe+4nWq7+zcgHZi3fbxv/nDLk/pumTBmckDYkzdKu0cA
CDD1CO+8ufhP4B1yn58hijJiFUuavexuRu9QzfQ7BeCPMEP1ST0v6p4goukDPYYB
mOkQPw9snsJiiX/lTUFJGswAfrk4bE2vPXOdiy6qddrHtPcPbZMKych8TX9CxDSx
o1Nh6ltDcujEBuScvhRlssazAGLcmW4IR6lnwIJrsCOuDpS+a8S7ANvUMRCoGnYL
DXNfLQKJH90cKJLIwBk61k6mPDIBfIh/RrbTG4Srro9K/LtJJY2CzilTFzwsf9HN
OjWRYCtez47kx8lsvioJQz4Czx6UQO5Lo+TSJjPRperlKnFzwrtv+DeQg1IrGyYm
4DrmSPNqn5t8NVvxrI1dGO0WNJ22R4iZlrXWKC2hS858KM6Qt1whwEuqoZqEXuth
VtzsZklaDdWOJRNtVtrfRDSy+KL/K8locUXzlbfjYH+4nO/a6rqGnuxNHgZoO+zu
gTGEbwDCgc+iso8cJWlF0tCCBEIpN6abbtbp2C9MyZQ8Pu9gt28kVGy3x9KK3eeI
vViLDjWuHm+Ui0i8Ip9EX/CuCyuTlyky84E5n+41fauEvEKG8J8Ef0pYX5yJmPe+
O97N1FhPOgSI36/tsJE9ocrgVsYX8n58mklOwqlkwDvicomzfEFUSGl86z1uN/lJ
BbvteZ6Wh8mvj0wRnrG+vIsJbGWEnYvNxJe4wzKdTOOUpv2AXJpB/8pY2V1QZyuE
Pka0pnuLFmGDgvKF3kPyJOS0CntBAiPoXu7I3XQg0V4/h/nVKfgoSrw92z+hb428
hi8UWhIjZgIL9Ieo3+GEWw+TUSWDviR7SKvtRcTzN48SADQiFnNgGWGV0X6/yxBI
+Bm7pohEj+Mi91zADEUHzmDfYHMAkJfpchBXEE37oXyf01mjUH7Vava42XdIlyu9
6OSHBzf64tOTO1nxGmY74W6kYh46JMRndWfAu8As3PTry+0ClxwZirvwr5vNPrDw
WaF9awsOFsixMvsnM5eR9lZm8uXu4aLH8SaEYMPIPvQg4+eBZ+83gJzi4475Z2Je
YPQowtiUb9nlgOwUi+sG0TU5szhCdFq7cxLe6hZyuEMwIUKmHUd/z/XEdSg6oKmb
4fBAH0givICIUiKgTrYalJMksd6KbrQAZ5GzzWH3xZjTgkAvlcaSYq0KffbN5GrD
/SwUnfqOAjkrf5Zi7RwZIxidnoCYCbzko6APsZ923maEc73rz0tOIdOJw3jgNxn0
0aza4h8W4R1l6JBMkX2w91IL/vULChFfJMtSWTI4spSiEjSFTX8y+Ues6eXSDQpz
DFSYS/V+qG4o6YhJGm2uy7CrZg3WdcaZu731uN7lzmLBbCopLieqzaRSIw5E1yOf
0PiFlrIhELXwPvbrUetqzdKCkZ9XEfzwlKUobwIsW5Cyc8tVFWamJMgHHebp5Zsx
YEN423f5oj1UgKoyQs0gdDZQ5269fIdfgr9IeOjaFD1J3l5tMi4WVv5XGeTJQcQW
izfTdCXZ83RJomsB4wZilZtDcc4xup6GgUokp6Eq3B1LGoNt3x54BeOijTar2UT4
E2FVQQLh/ahUd2dWU68AMObjDrLxfN75xZ5oUnJqa0rGsGvFzXtAg1vbCu8sz0ZD
Pmjx6qjlNlnU8berEVaaE+Z2N7Bk3FzzvcQ3LVrRWBlwZHvEXamzqUTELM/uj8aR
pEw01tjDi92JHRgNQ/Qc5eltCmJqM6h/L54mEtum/1Fot3qIi0FFLFrMBUlB/DIG
N7XGN/mu+++3GuLyp6GtT2kYO79zxIDZjWQMPve2FCeEAJXK3PT/uoYMH7/cx2Ex
ba4B+DfXJf/fLDzVrmYJQJeQgls76Y+Agb1d2kIKB1EhCG/W/m93iG9xuPkGF+nh
idSXVQRuvPW7SqvFr+NbYW5Vu6N2WnXwdW+VR3G1HvgGgs0YUlvv8Hd8KgcvBUhA
+e+CJTYfIMNqF9kSTeRoPqeMjRZCfH9My8GrvLG20revj1JMpLJwszx2CPwbfg/T
WAcxGlnVXh7S9EGrKEDnBlUh88aOwPzcTXjSlHOWRS4ZF8gZEFCZ5qW9ZidZfThb
rfsz1VMG1iiktxv4j/Oo1DLXBkPSZGNJ7o2WiAQkchC1Aq2BKYhmZpA54Cbat6XE
FUX4tjuleYckZk+LU3JkgqBkvGGwZTLQEx3x2LPGG9AOon7+iIO6xIEtM+3iKZrf
sJeBsbbjglc6rR2gOuX9Lz8Lu4g7MAOVUR2+8We+ynIZjO9Ep/mIFyHvqrsLYv22
olxkJjU/dzySOCTG3+Z4p5MwfYJ+v1GkG5dm1okWI+O8hEu5gUOD1EqHqVydEN5O
sS+Bhq9FzP80LZPM8tp22Er2zJl+1WYpbzJID7DboTnzLPfbbJ2AIUkQdXu6stgH
lmrGFZGIlIG/YPGUnvkpEW8cCb/udxZRUaZNLd4RIx8fNGJz7lAJRcg4LUbVUdmh
E5vRdb6sYRAMIs31nxNnb1N43clsduZgDmUpNEUCQy8LyqEPAl8ddaA8gabZhlyr
ek9QnY8B+1RP8fNVGGbw6ScOk/V5z/qzu+2Y6onArc/KycigfnDJMTwmrarqV3jr
tuRTjoSNS/D4Y7cGG4YCXXNGbG7McMl5zk8I+5WztKlpXfigkIT1THhY5bL09Cns
eGgXr6XxLtGR2x8Nzu7tRVeqMLkqK/aURN3MfT8wDUL5xgvz/gIw+6hQoo6QbOoW
NOSNamGFgXHE7Sv4Rg9VB9ggQgBvdVP9etOSQopVxQsFNt8W5bBtfyuEA9iwI9bC
L3xbXyrOa+Jk+q/i4w0qkilVWJTYs9XZls05l6iyERWU9A3hykEKVd3L1TbIz96b
XUBEgxQLME2b6j5cFOTj4wJCONKGNqY2VMyLcRY3rjH2vte+/CbxmOZF6xkDElVc
gOoV/OW3qXran9OTLwL36KDUmcp15aP4l07TDRJa3rzjeG8I65hZBvFyUZxLkMbq
+Drr0RB+IB1TgZwUA4+bzJ7vWnXp9YjtyxMGnhSJW9hX7GFBf0fue7PBIS1zPOne
NuLD0J7oH25SB2jW2/wCs1NCZPoBD7x7rzHEFzCvWEZKhOI+fM32pKK5WV47RmAb
jCcP143b4u6kWRPYw7QAo1mSUDsgM3ggN1H9WjNThZxjfhPQ+z7I+nJ5DVLXpnWG
TLcTwutfcVsDeukNwaPsO9gIfKfyo1VKT4PAOIO2hLjzw3sujICeySlppYCl6ts1
GZ1YftifGari1uVuF00wiLmX+AOZE7OS8EJ/hw+tnsgaanRc0jI4F6CrqXgGxV8O
z5n0h7CpgUft5EtL0SqNNQDC/W+cvZt1a4W96tcnXOXedYNCXQh8gQsJCagfXfaF
EcEXRzuGW7YO8rW3l94uj1eEvt90YTiXStTDgiL7Kklwgm21HKpYO21o/6V6YQq8
xa6So0jZkEhAlwlXS1FSLs81fiQpCdnAgncIh0MtOLXyYXb8strFhyX8EFUEvBwO
taFH3pmkd8lsZPvS6/RD451NOSrrfPsbeGMnBygu6XHnySuxWv6qFmqy4ZgXZuwt
CgfGgcXSNPhBp1X47cvhnKuZppQSF5YxQq4OA/2inVeoZkkpAAry4oYeYEDIot3j
BVWm0jPwUtIibdA9hLbF6Ta0QjbuiAYF/e0OlYmIhh0MwfWCf2e4gaL0extMLcS8
t1zOJOjlyJHagtBc7QKrPRsacon9I7O0GbMSBOQqR65Mk+kq9rEdLUZfc1uUdrMO
Le4WTaeSb89sAw9bwqFHDXNBAcofEuqhREQteklXfnt8PqUe1K+kj/1HGDdAo7ov
YwPIAeE+g2i0EIwjdPkVrH4ghglqop6xiz38ZzPAjBMj/g6lERRMCWNa7yQsr77a
mhw6AMMXbww5OJyukp2NFA8xVXk2Iu/U3QMmOmJUhn/Kijf4KsXkuzH1LQXUfbyf
eUZYlZlUgxg9bOBmHRBEvJr7rfT90ncZYjguuis5ZpwYj1xqjjRcgnHXRBsqyO3W
jhyW9Ova18SgjbJvBj02nMd8/pT4GYpt6KF8zpqqIj4A11rbde1Ksc/SNtO0vITW
KqK5XSYMtH6GqKoq8kMq8opIH8KoniOAzmoGDwtBDpFgJREjx3d+Bnk1EMGUiMJi
JqYnc7IycmyftMsi2ykXOE6zPWrkrBHewBev3Q3Jz/GL9o35flezPsjtuDl59LHX
Ax6y4JXRp5hkn9YSLbbBNZ3NfBnnq308ChEPaCQh0PMz5mWQimmnsCnrj9jfH9HQ
WLytMoHXv2xLTpnYpjWzp/cz48IhZye8sZlcSRzoIPTyLlPr0xMnfxj2C4azXACM
3rBe6oaaYxxGcX6AZcVIlQoYoCXJTvUdJjt013eHA3zNu3V05P+qoKrHneD9J5F4
mkRuSQGKEgGEfCCFCvrs5LWoaHixMkCXHIMHZQdcN3mrDPZgyphELGGtbzGgN+Bv
zIj0OswltIssUmKHazvf7XCPyrBd7NFoDVIpEFIdAtP5HxQnxB4FgN49GGwmlWUy
WACy1HkAh2Mnu/dMwuVNC8lzjVBaHokzS8Wo7ChWTecbvxUZo30njOy/IQI/3WT0
5XKmqhhI4WiwUN65m/9qIVFK0OvFp/d8hhIv7CO0lpPfWxstWW7fzg4M67kLV8tK
IlNeju0D3H2nNxm9CynZbeQAXxbsO5v9QqjrkwTjDR3XFwUliQjHc86KwNPUApUD
KZs1guH2YDA8I+FoveZ7fIlROAwmDu3tgYFStw+xGqUqOMSnAZ/zra7pH7QtEf4Y
yypmPS9T3svTp6KEXYL3dJse65nkf0TnN7DLwXRiYwEVPC3b8Z8QZWDwVgkU3n9d
VakvB1u9ZXMExtukQHo1wv09rWXltTOWoBGAAGGNuFio2cPjtqy7MTQYt/XmHRym
hesdvo8yk05JOZx48sZpUykYnHKP6LOepK7dPezQgb3xpaqzBYd8a7kmfrdb12or
GffdvuYxdm4twyv+0+Nmph2/dFBtb2L4DNuvW4/gnSNVEXq6JlS1o12JLtn+aW4a
uiczvbNXll37csEKey6R1H2oPftCPGJOul8knmaV8pb8TYiuuUmsVREu6QQY1eWG
E5b8f2e8+5oE8sJ8HS1XMAtC7MJOkk2lxxfiLsGiuHaWPRKOfefk8Umk/z/0vKRO
tp73q4/j3LcJZDOG/0kw34vu7K1YLevZdVzmgUncEzp9LMZBiyuhIyzLlI06yh4k
+UdTEGHHaw+kZHMojszIS/GsxgdBGi8ePJk+D0w+KwSsNVDDe+LT4olyulyA+zlX
uhe/rhxHv+zd8MwFTfeUwYkL3WceMHKoreWd13rKpa4M7bOSrn8mjmZcVpnFyhru
cWQ1+M2Bu5nX9Lud/XdqQnEr0disCAaohR8JmPMkwlkuUuSVgwz5zKrFBjenm7Yr
BwKQaM+uTKCTMHYQ+QJ76Hq58pgOaYfPc1ip4Mu//lG1xNmthRG6Qb4TCv1AJea+
yjKdd9agDV4PcLUZt2qv3qntGdhX3Qv64eEgFQSdBR38EsG91lngZeBLsUSyC6bl
F9Z8N2KsvKQrRuUGORpaTNA1BGtVa+kYkPCnVt011mxh4HAoB4lo5k7ApBAh69VG
7XgMV1GrsgAkGCipDmC+Kf75NpMX9FI63iAE9wAiwAjU/GatXoqUoXXN+n431RCH
nmmDC8n5VQPiW8celZEacSlf9wJxuWRQZaaHfj8SofWru3t914u8R2Q94O3uHVs3
fq7q2XJYTLOX+lB9KXqHN0ZWYeLoKxwF/kPrnB8bhTUJm7hwP0y/gE8u60SVhtMa
PH9AixvdB0EIeQxrPfU8GH0PFtuLLe93H2GN+toR9WWaGEcSkkFYhg4KrV4B/UHJ
Swor0rhez3phUH9CMRJGPk3+PRXYLH2A7FeUMDDzdH41pLn2ISqDKnwL3n4t4Slb
AGgMMf1EKe5vyn83/BUfA2IIThpwky2qoZ2yxQ0zBOz3s1AEcTf2s71j/m7S81XJ
ntT16nEkcq6xq82WJ9nZzq8+uWOKFOAFDTNHXyR954kRAzxgGjENM3u+HcWZiQ3E
7lNHWdmhh6pMTS4cHc6PSleXZ+8KrWobr0/KLJH7m4MCr3KhA/p6i3ynrwuQt8JG
6L8j6E1mOQoD0nFb5IqD2EDB3ob71CiDdAY+sLvWaULsi2MTDKzFOyEv7edxffMi
hR7UEp6szGDj3YkEFdGTEbGu693tBhxDz99Fx65n2colGmuGigILxONMD/k0LWsR
/nMYi2Dss7MJSpETHE0qGvOddBJrP/HFG1jiIeEFtrBcd0lUZ6FyuQbEOmgcPG+N
lL8559Y/Gjq18XG/Wrz4IbVFiqk/qlmnWA7owzcKlnGXVBaawnt2tuYGALuAGETZ
O91TrZN2YszBIp/KSlo0Rpl+IZDGJhBsGuHf+IqdVxmhgz9/BIi7yeMUq999kHjb
8yJNCJmapgsJJFznsbedg1HECsR8AvpLgVHhfoj5eIRONsbKNz7dj4tq5vxsGm9l
p+jOq4sSfHwOYvdZYBnH4G/O4Z3PdoneWizQGA29CZMfhXxBN6SIrWDVNN1KDrJ3
IEpgqnaeU/YhmG49XDPHNaxR1L4cuNlDsdHHTHCtCN6YGAjpbWa774hRO+b8RLNj
eX1tOsKrsdF5VzH3Q7kSz6EMotaNamW7/+n+wDgKlj00ShnGphptvzBYeu84a+kc
G9DvowXBe++6OKgZUnqJ9x3W5/qZ+8VIUFsoFybdVUpewHejbcUsDDkvhcx3JSBX
CgNH3mRQLOpiUdBO7sRsDwavmc5peAyV2C/vFVQJp/x+gSXTyTFacmhHjrgnKQ1U
R0oDCfYgLLrkoILhYXrX2xlbMxaLKMBc+LaAjXwcSKUlZPxaLXoN6TI8DE8fpUTL
a7jSksnMj5Zt1krRHBR4vJLyraXz0BimzoUJ1rkDFbKxt12F0U8FVGfmTQkfDs7b
46YnKV14Sk9jEqm+q+TjpwTBqnP0KlnzUNShKrQM+JzRq8OU3tOtfdRsmohbpFAM
EE49LHFy3ni9KalPbusyj1mj0sAJdVfajTtA8kZdF05GZH9yW0WwNMqoMJtC4awN
rCTdvLpf27lNMSU/DS9biBluerheAYnrNGABRRdWQ5ii8BEoPHOY4RUkxbkQ8s+b
O/x0SVAC83MwsFMOxuG1krT/zAjrc4bloOh7sSqJUmdiWLTAxLuZCmZlRnxgPros
24E2F5g1tCuSeue6C+W5R6/68zMv4pzSw7Oj+B8tsWygQmffIUcJ5C9808AhRaK8
4ly+TJ1dJQC98/P3UfOJXHqLtZV6FrDWJQQmKhNI2hYgEAJ4FFrLwF9/gQ1xEh+K
Ho1Ro+7liZC6EkoZB4/8G1c305t3lm7kKdvK1wYd0y3ypwZZa1fjevNVoP6Hf5d7
AWUxKyTqJ/cqNpXJ9+chpbav2bip0MASqdGEHm1YN+SeNRkBMc9qVR8cpm0BObHS
kL+vfZfBPeZzAO5Wwg36eZRtd51PWW4KB2kgji8Xi+li1UdPPQy1fsYgbUEvGsOZ
kUFRbuhtI+VdHQ0tXvfk/9EwhzVEH+ciLjsd7qYzYfnj5psyp0tNax2OUgI4nD2w
WAp2VzVzD4ksOP5CaeS+K3R3x9fPaBgiZkz3Jiv4l+W5ei6jyK1lmBvMW3804JFQ
rKXPQ6Pg+kHiaXRS8G9ZuHP2eOZprwiYzUWhzi+JH144cSdfGIzrbwzwoXXnc38v
cNXLsloMBFksScfwvUCREopAOuSO80l8CjLfADeXQNm/u//jj5fLICZ5RyLR+a15
0UIr7iyfuI4Rxkx0sUfS2dn7zs+psEklv9yle2b+nXx3/mTVp8+ydJTxwn1iSrT/
B7WlWXeAchLdpyLiSChvgNhCRRX19gMUMTwmgOV8336pqj9gIHI/wsjdpFrqkVDL
mpwkj7ehR0B5YB4J0Sj3Pj02gQgDGBD0YntBXEBILjH9QXDGXODxuH/XdKKQ80WS
lB0rrDalmcNuc9q4mp92RyIoTWjQ0lbwGLz5fF+xQeTs8H+cxFP7ORa1aRpagtbD
YippV6FK7EscGL0CznBoq0akTT8ELGyWFUrNNp21QMWuxl8YgEHNQUwxQL95PhN0
31j6IrdkGAvJjf0RHFbw2SOMvIDZ4BhbLmM6KhqSXyEiEG9tWRgAlcwB54Co/zWM
gUGlDpzS8XRTdS69vWAiw4JgdvlN25ukv2nYxJAAyICSARK5IKeVzndRUKL4hk6C
9cRDg9faNDH2Nv+SZ0+eiKuOgkhr6e5vMO6+JBMYpXN4XH22lWwFN7TKPiwMGM71
RXFCytMNdu5wvgvGUilFaMRTaMUJ3ioZc3O0FVkNRYZclTYBM967GXQ3V/Mi4TBm
rYiiQijAQzRyaxnN2nmG3D930/PTgDvCXOhD6qZ5PqZcMtYg04mMUqW/xo2wbXkY
UQhd8wJpHqsIxuawQuCqb/07TpcS5OWaTB06JgWwsMlqbxthHHpTvodRYCtcpzqI
FFsORj5ZujPQLmDqKr2hw9k2to43kKSxWPmoBG6ijotMXL6w1BYHcNQ3RVOLimW/
hgRzBLcVOFQAcU7ggCKMuyGkeq+qwaS2rBePuP7Qltno7bdT4+EVM89oQYfJwVVZ
svSnqlV183/WugAeoSP6l3WBGbaL5k94Wi1L9y9nxmbxNMDbvU3H7gYykgd7wVE7
DyQRXtNBLOQcjRqfGMDZImTjJsAFCvezBXkrk8ltkSy6flFzbNC7NDeeE2T83REa
M73INF2siv4Ykchptx+0YIbnJnNq9GwaVP52eq53Y+/AXzbL9WydJepl8AUtnpvW
F8jbPGEADDzcoc6Guchk8TE9ofXq/9vo+Uwi/R77pI5ZkPQFzfxiMq7a4mPP90tP
1fWzvF8MlNHhGg0mXZZN4q4gOdrCxaOfO3mqHs1TB0SHeJBM86b3yft3j+3hoWYv
3u2TqxS+4BwUtxpiPBeC6uJQso4MvhN3beT02xNFK0mFXkeu0LsAIU9GTu58J6mD
W6LWHL2f8socPRMAqvaxZHfRnmSoZhd7Bdkd4qim/7bSFdgWXljZb2EEUarm1pbF
ZnZy9s0eb/Z90GFxpro/meTEzvGqvSOb/7Q9neCLEONdBk25jr42QrWMK4/2BeFE
3aFznYhx21/Josu1MHk6U2udkD94ncTWOEceIxlS5PcjX2zIkvnMvHZVMo7+LGeh
4VBjok68M6kz/R9mGyCHZEWLTIUnDBcVo59u7jpxqzWSVMG+l0I+VukjK2p783u8
jKBE305mVHeCmdUqRPcfnbGi8w9jg/BT1MamoacP2WD9yt1wUmk4yMgfizToRKKC
6o+5eOn3Z+tCsfQ8JT0OcwqMBTAXMbI3lheyB4nyH3qUIogZ4rFIRPaBbV/Y7JNU
1H1ZP2n6daAlHYIs6T8XnOVq/MRD08RU5hHoWidDvNaOB99KW0RkOU1oQaBaWGSF
XhPgubVddV/z+/EO/eeiVhXNZgQRSyvJVGdadNSkuUcIamTgT2wQk4+eLkeRW9/w
Nn6F6hrSOs41vd7EswGvHN8TQJZklf6beQLFLkS9sVrwqMvaCCWOxhgcU4n4F1E3
D9ARG8EYgDB+nTObhMP/clZsFdfqEnWoQoAjzsPrISnwba4rrUvqY2fUv+ig1i/o
NT87a1XhSRQczMoOdVXJivKUV43bjiBZpmhEuzm2nGrySoEiPse2FCLHqza/xmAV
vCj8FTkrkOinMoekelH0+KlOj6Zz68wXfAPHR+HsmGGM0sWMK46V6hQ+Bdd9/Ahs
LGNxL6DEkL9G4lDQw2t9JFVVHmw+Tzg+Yb3sjgQPF9KzDtSmsLY4D38Z1Lk/z3jn
xPH++C5H9kznVqEOcQWnkMvQk3zIlbkqWq321gdBcX5kEC/n8vOca0fJ0B+nF01D
5RQwyRfRjAUmcTsS9SWPS6kg7542T2GrpRx5GKOYOL9W7MwfHgSgLGxDLmNlTBVw
iL89PYuIyjuy3WVrh/Qc0cD086zJ8ritx9kLEIEGzjbDVdm4Ttgd41EIyWnlXeIe
wIPLrAWflY7od1Y9hWK26IDuO2092pLq31+2Yz0PfBsZS54/XUy0c2eB4zU4qW2U
NMcIxFljiXKWc8UoCrlZDDvAbDszwQKwrzGXp8A0Eh6+EI8T+haup+fEfpjFGLJ5
uk9AccCfLdbxmp/5hKLV4r4usRyls2lrkU//5rJ4jRPaepQgvXgZDOkdjH8AwECo
W2K77VEhYWmvajstUQCd457lWTn+No5teYI9lxPTpNOXqvq8pZbeSWEBJysGPy9d
7YnU+5eNOoVPUVlEPmMwpfgvxWoS6AAAwSb4JVIveM6CH6yDkRhSaXXmfhGH2GF1
8rJw602O9WxRDj/UPN4iWMRZagOGRT2EFAXmLyBUk1v/49UFUfOIzbe67XuEwa4z
RhDukaVIFdrvGerGnHb5kUfd/jXcfmzqWl4xRmmh6D3ECPLSoXJUuWGtbOmwqXPC
+7zsdtYp/lDhpdD7Aj2Sr5rC3tykwsg1BR43nZCb8IMBaZGiUY7E5pOgvb2ta67f
f/65Gmnf1oqybJE4kcx4Ots324ggcxOVEkZRQ6t+cl0=
`protect end_protected