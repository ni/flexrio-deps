`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1952 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
h3mPGhLvpV4xDnoJxCkEpOECxHFYuMzYlWUegCgnLdkIcmO+DLAn5Xkk3mH3G2ke
Qj5OxXjQd5+GrvdhX8EPk53XBjk1HNE3QL0KbIzVcP5qK2afZdiJcU7Ssab30pN0
4aHtMMruz20q+umlIBauPLE5N8ZSGulzs7CFL60SsrO9eGo4g1i2ROxpuoXvpfHC
zczs/FDpn5MspwOwt6Upq46RIvFSobFOqC/Bwk6h2yNlrkICBzYzbUroS6HXmGbL
IKlpiISwMrT0A7IxGt05550k5jatIcfVUzpLm3BffSVFN2oy34lU4yWFuTT/GZnK
5Z+W23zB56tYqhYnf2G3cdictmtWvOIxs8C/PJ4m5KOgT+8OIFNZT0oo7OQjDTBy
aIfNHbpeuVXlpakVaht+SqgdPJV2GykGd/D8wOO6c2zjgq+Fl+FwXcgopZwfJoPm
1FSnErd/RXo7gn1xX7nI/7HSxYCK0IHB7dOpu+uBSshEOqR5jGI/hXX6SjZC0q0M
s9hVgYPS9LQ5yBxHa3PTKyoBVv3z/HSlQw6+zdQBnwmkes10/HdnRU+d9d5ro0Hc
HSe2dUqY6caZG/Lg+cctSM/2NWviMApWoWjf9TNakDBfrWvgWQ7Kb6Pc5oiKfkdV
UpeLKqaMDoMLTEd8585EYkLlwevMk1IuCVHoDs34A77ppdWxEva1b5JLzxlZsMdq
2tC1cLEW2K4LVRHCW8oyNww7kIP+cCPdenZnUehNnewjQ+FmfoGL6hVHeb8H/Qrq
wszvYYiZhzOB74wP77N/05bKqKTx+3O45JFbggNUm7yqsHY9Iat+k1o1oiYtKmzp
99w+Xu3Z/ujBc/lD+zVemdfdhScYSiypt0Iip+N7wXhwi+XJT7Oc7em9OPqrLEgQ
HFuM/8q+3pFjmGi4RJAzu0LPbMJLfKMrRbvFz6K0TX1jp+f98WjsvyHblzdYqR1s
ON8XM3pSkrVXxjbVAVFGoeZAtwenrhjMMtiv2a4ky80OSZNQyKkKLkn8WE/bOHtp
84h8ZlF+rhtQ1lHLSLzgd+ok1Okb4XkAsnYk9jvkl1fIfsq4UmOUhT4uI+1L+8+1
WG3vkorC1p7zVca4PC5is2gxPBsYkpbg6YY0M1JAKlMUkdXhFp9jGaYjwnurMJGx
zYLEe+Gb0GLWf4T7jCI69E1ismpW24JX69F0OvELOpNngpjtxeX3V12PBwJLiCT2
rbk2c5e2SdL/CNJXFh04mHK16Zm3AnfPD279CJ+6GlHBOiNngrgZ5TcMiNt7RwnZ
a6RAug3EO/9jyS/9cbgxOpIZTmUF5gfZP9rmBNPClkSxi9YAK86K3i8H41IJazgc
rDEtWvPSIrqBDdzCd8wgGhFraEKea8QDiv3lUL+njd424uz36+hM+EYZ/MbQfRUd
n1u/dpEs0jfb6kzGPNATx2ulebtzpfq0dN6Y1bVOhlsSy6lsQDmdI1XUTXt6M4yf
S5mivG5N40Iibx0mG5gpj/XRXuaO6nW8FAT2p+JxSS4b8QuXoCKN46KMNIaEyh+P
nDG4V1EYAnfzYo+HE+USp2XiIx5czJpc+QcRBp4mqy66N3AF0Qqwki2JSjRCzIY4
Z9NmNB66zO+BbyHvOi0d5UwQue75BAcRalyaMBbTjcUiQxVYA3UbkxrtPbRNrQ6J
G6fuqFnH0y4IgevR1+h1LMAXDDLjoEYncn+kcTqpQ/B/T2XaVapNOddwC/kyuVoI
N+OhuH1BAT+zNMsDa5z6ZnU/w6REJ5ipFrZQRMHkiww9AGICc3cOD7kBUL0cFrPg
TkH2MRRQ9LGtZtbk+JCa4N+iPj7w233b7djW3QvlTFuKVInLnsfZvlpfrKjkr3UV
VSaa8XQSc4aAGvg1CsuMrBZbvnNA8SawYTbOo+vdfk8deb0i85U8Kbg29k5GnQBA
13vgbRCNOMs7Rgihq8XQUoV7df4E2eTjyX8noOnfr5sze03PggYPGqxmKozLizJl
r9pBYQBXi6BD++eOIAQNYpwKJ77F+Nu5vJ/PRLiUKqKtNB1knPYAU0tQEwr9TKtk
d2vxUZzRgngUFl5IPC8faDC3kXiLEjhw9j4rDTDbEOwl+hJbiu6vmZl7UFzt4M/o
pn4H/MQZy5FsTxj13/C3z+uX77tHabsuKuD+eM6fA8KxL+/dLaYGz6bCT2vrdvAy
rdcJWGP0S1MENTdhLdOFqgPVkHuK9G9w1R83C3BAKM1ejrh6Fx3l+lNPrb2rRYVx
QJymUe9s7VWk1BR5HD+A8NRwzxcSiqwItpM1pdXWvezRlJ0t7geLZIQ7y/SbxcBV
UiEFnsUeKBHO8ON6lxJ8O4MANaHEVNc2ZD4wJyDCU2kNrq/GBAj3V/wLMsCAgxVt
4EJtGdoqqTgLygieE2zWahjdXr2G7iFqEUqWbnYtDTiigDrc6pcxbKV6xRH35I6E
YojlmCeHC1+VjAMQgtFVHCb4NSMziuUX9Myp/iXst+Y=
`protect end_protected