`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6848 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRu5USVS7579wHpheYeWNqWFqZEm15wTQ436jZJWl2c+D
Htzd7ds2HQDtAIClM39VrZ4FrJekT3UVRl1wR9wXDTuNY7HvRIxNUV7LFZb6IPTU
qrusQW87J+XWxIXEeznL1TvBruHfhdftqTcw5bZS9JYdb9GzoxwiAlZ5dsPi9bvq
mBsF0lEAQsX/OETRpgxCxJB+fiDHJjK31qVXauGqgJRAVBEUqkMD3V8m31T246S2
129P0qCSOj71mmiDkYyKlQGn+OLeFm260OLgee2+Fr7eISD+TiRktjYXIAThqi9j
wvWByxng1v5pJf6I6R+qbPrxaxuiBsyjgP5pbiRBG+XjFXiLlCBwbPG/WGupl8Jb
dGiL92gYaHtSdcSoZ4CYoa/kiirplcccttZ3/qtdcNTgmWBCd6iLq/zFyVYPR3m5
AN0eePlZ9/416zQTQf6l0l1jC3zHWNHVx+rF7zycE71lxouk8GCejiWhYet/dlTY
eVksCaMi0KuuvmNRvpJdc9hM06O7RfIXWMhE7l2HaT/t9KWgyyJ3mGZJdzWqasGC
YQC4y51AX6U+QySqTubGzkacLDyv9dR0kEeJXK6+XMWj7ZqVzx+46Nh48PyTNUvR
+gq0dK5Oe9KPJt8Qdyowj5REZkG3Gasmzq5NKrYkNpbYsvpLWXOFZN4Bk55B/YXV
V/7Tw/m0812x1EnqSoBtlfNE6gi4M03DxE5pz/ootRNf1UFDvI91pGIcdZ+oddQK
vud4GKePzVmz1MM9ph+6QK4STVsC4SqOd2zIt61AMVmSmDP8lhTAxF3/hlDV3GrK
rkwHdOO0s1TkY7jrfW7j6lbV6qJ6bfzOV1Cd1cJkwYeL/qvbEZg+5GXMzi4Y9miq
n2jgDG1kCI8OtZ9qPbgGDmaUK8LEYwhY3oskPjDbr2N1fX9IoGOKQIZaRxRkVEhh
2kDWpfmksGxno9aKBHHbov5iugrF5QRqLsUqyxBRIHVWDZExu7vYfy7Nnk0uS5aI
iWw8iQ2uww++y+ZgHsVCffyirDXdLJGlx/3yaa/P1Ku1/78b7xtAsYksiB468J87
/Mgkl0EymY/omjdZxCBq/H73ZhjoBxvOEIOClTIdLZRcUvOPguMwuO80rgxreEIg
fJZISGkJZQZTY29kTWHY1z2iPg7YdlZNq0UemvL2SEIZ/eIWJxfwS46DWTmwivtj
da3RCazxfQ54o1yZcF8JKoPjllOUMunBu2wl8hfSS8Kz0uNYq810Z1l8PDRnI1AK
4JWwl+5KKxeo6Ae6pj6ebIQKTfx/qgM7Z6qbdlaibKIuQFM2H/o9hHAqdgvhVBvP
cHQf5tujWYj8tBwkemaWxi+iV1S+3Bi1W2EniR7w0wmq1C0f+wi6BQFcT+bNt7gF
TnFy65o3MWnwSfkY5bLNzA/0Z9k5HM/T59Qu06eU1zeVeEef2F8wif7k9A8hsSeI
JTGthveoOG1+9+H8ZeQzEliH3etik5GxeKUifLJAggtJPN1dVX7e1pFOZAnNJztF
lrMA5bkyh5lTXOfJg8mDZize+hbVzdnBUQWCaTVT/DiBLm6mWKI9hI28X030h7Tz
jKhvYab++7idfg6bGV4nRC3PYlhdbxeJczkUOEu0vgqe4cfDhW/ugo29HF4U8tZU
x5i9km3vbIyOXEvuO9DhHFr+HMCKLcDXwEqMNzSk3xW93fezkZbPEIaS+Nt3qntz
gCg53asq+mWtn7149ZN3MOgIJD/NpA8vzubtOEbEmAGfc9IfcThI+DcoODhxI4hP
6surcsnrff761fSH6cy22jccMGwi7MKRC/Vy293afxdWk971cFUpyIRU+itnHKpr
cXWHzbO74n1ZEVBKzcnW041ZkqUJGK3kRPh3V4jkY8NX+s63oQMcyXAkyetjYfx0
Dpmt2gct4/i1bdQCwqESssKk4jbnrRq1ZQtPHLb1LpuV4fXkfHmNMHtihiR2mjdi
qh9om2sFQge00J50vbbOekqP/udRGZI8nNm49cY1S1AZbINOmDF35p14jJcWVp/k
bQezf0xtuwSUx7j+KoJMiWBA7EkSBJJypldHiJRkwgeO9pdZZGsKOg8G7fNVzgCS
xQQtx7pfFNC3tV1nAMtYakboNlbuGLlFTwNTrJSAlzi5OAnRr3K1/9/1NV6UmfU1
cchLy8VgSmDPiF7gkTfFx26H15RuBso0QNkkUGexc2hxg7eqTQ8W/20ywOPfGssV
iERB+x/fM6E367m5tdap+OTYcpJJiBzSLCUICAtcJMrj1Ra3+LV8Co68q858bCaL
kvSOk46iT2Bh5GyYGWIluAITlAgGGaKcPynal2L/kaelcDx7gvoJ+2D1C/q1tqAi
TZMreH/dNZXZlJfS5s9iz5VfA2zwMPRcLge3M/KLDv1y3KIev+igiuuqZTMH76zl
Bad2IyLzKeEuiJnK6QcaRdlRqEhyOyRhbxsTT9eo+vclMKvNOqBMD96A/weusmNa
venIs6hu/GJ3pzz/2xsTxRA8a5crc9n174ITFvHyFtqyxGv4o9GwIU77oWFtJzjt
LhJzgzUgH9pjLcY6ocOBsVzPlQSmfKQnRAxLNn50T8me/2DRNhE0wdGHkav5TKBH
sSd/Cj7ohIu9URJ1+WIk1rQXfL6wNZEB+uU7m1lrU2hi9e9yghi7cetxqqGfN9+d
RsHAJoKXZFLlBp/NBEJqKeUaC6jjhJI4ckWTskzfA/K14BhY2RINcUzEweus03mc
vZfYUkJXVDFpDCdT6WyDnCl0rNynZrc0jYMu0SkSGHPdYmVJXSwAqXRVP9IVdhbm
dsO/hVY2/wBzLalugU0hjwRUATkmNjD5mUqw65Lq/b4LBEswMrBK0wzAc9e9+xxg
iBgUvNkIXFfzAjUXH7HraIAo1Vhi+8K5qIs1Eysg495XGx9197Az1CQ2v9Y3L59/
eXlqF22cxmkd663CrL9l8q/vdfs/mKR2AEJoOg5+fo3PDmLRBD6AqUsTE4kqlvFM
xlgiFsdnJsQY80xtIW9jRBxz+oMvhS2jypRnxJkJo5OgjTC4LLsNuL4/Fpw3P8Oi
MP5p4eEsgpv1r4Ft38z0x0B/MMnNmZWUonwDIn/3A4D0LuG51Oqm3C9ZTh4H52y+
8XQbg34WateU8RP9sBVe7ZY9jaiEbaxROYk7BqoBpwWGc6icPv5oflq1k6KD5tPD
FQt0zToUCv76iHbKftVS2IOHuic/6b1BqypJLVVsxD2IbcbJ++iAgEmFgXe5u4EF
U3dz8WvC/99xjlVSVTXmkXHMuuPoZDwPh3ClFJKdchN23iKZ0y2HqYZDtTb2QID+
LD98bMnybCEaN/3D1o5Nb9TQSWwGpE6GLVMxYGx7wyQvoncMEchSm2xE7TSU8DpB
AlbfSGeabCOtw0Oq8rJdPFfizyMwI28IvDqjVW/SfwWU5PF6yN8jvTG8KMnXO1np
2REvGt/yg2CRNRzYLQP9W7xzBQSrg52Ca94KusqhsMB5nl7PIqNNNPlqAQj0GYU9
pp6W3VPTC33R+065/joke090psn/6ePiJoUzcHUlelKxdu2/1pnUGTysaHFKPfd7
LluInVahcLp8j6jhuBIbgogjO0RH5XcD7E/xYnzis1AzWnJtbuvKA2R0g1O/VHwE
4G79n/oLvug+zRykdprGD4r5yg9hpRQXY59gLNwd+07iQkoQ02aV/gz+IGZKSs1u
gNgOC9Yi/sCPeNwOqSUd2SyeVKE8k8ccT5jjfh8pmGXq8MUqe0mx5vfNoEoI325c
1pu6og1DRWps/rQ+nuKeNb0/2UxZA9WA43g1pqztS7Fak5BvUe5R/kVZkpS9wZ7C
Wy6Wh2ncxETX56JaXGUKPuObZNvjHBANJdo2TKO3m5G9Jnj8qwn9B3h83btat940
jiUjPv/nJf5WZ37EpFtpt5RJ/n0vKq0po7/M6jXXpnzShdsz6NkURA5446GGkPZE
FFAYIGgCbjZg+GkjzMLFQmcAjVED9fg/3tYxdX6eFrnyOvNbp0j4v5fpDNuvua9V
tm415wjb+ZLr0c8S3FEAA0taDIgFFrAEqhMtAkvPveqpRG47zxtZhug8rnG01xcm
WeTNTYOk/Jbc3gCmmgEnGYF6IGlfND6mEM/CMBxevZ+k+LSw1MCvCBYehM1GFEgF
7WRTRsXFa8Ti/B1JWRKwyvn3ku/iAf2jSiPv6Gulrq2RevNkggor0XCQmrpEs+Si
NbFn6/iYBlsMXQwyd34YcpSs4r3lDOkqOAm3DQRshRLArUkxCB6FV7BC4SNTop1n
0EZ7FmQWkVK12geBHajqBOX0+XEL8ovzbOXV7tVjR4T8n9Rw7WIvL+mUK8G3zz/K
Uzr4OfhDuzzk0VtOHAGIsAoO4LV7fM7B0ABO81uEwIpHvHo4nKJJqgA043OLyBXK
21a7BIEQ0yYGZF8gFJw0CdKz6fAJHN+A5cBDY+I/kxIgmCItW3rGBhyI4+U8qxX/
R9LiGSDFSRDWbMQg94Y8JNH58kFpRRu9jYYWCInFTacd0f5y0uQF4u+r7NTGh9oI
WhqODKD/gOH8kOL0pU6POeUL+j40BY04RuX3eK51oUJ3GWWNsRpTm0tprf9ujMfx
0HdSpcdSfQeHRvro9LQnQKo/bJ65tPb4C6702wsZYo0R+Qch+wCaC4f/j+lRlx3w
56d2ufWbuxrmIPNDjDC8gzZXZZD2Vla1aB2lUCCJJp/cpCwMTSWKHp/Oh6ZZ863e
U11U/Cb9Kh9MfFZ1T1CxhzXg6gj+nXhxeE2OvZhmoNDYISIcsHkpDLSBFcRDpMMh
3su6QAMpqYVamFtnoADS1KTV4yZZdZK6eoO8QBDLd9Q/q2Rh+q/w5I0lj3WjuRwc
5ZuSAgvfGJCkOEeca3gAJJD0BQpO9cZFLyJD5BMQsDTG9mIqCNZCEUPLoAjiE4jX
GB5ngjCNqWE+4Pu62ajYWUR5R9uxx3ZXW0otkVB8fnlsyQtgRfGcz9OYweTSAWUK
GCZaWMu6wcMXBVLKLcd3Fau7gi6oKvjrdK5IVIwcOa3iF/wIRdQf2dh/Zj2DjhrG
VGeXUknWrtTHCRgJTMKfqENWFuag1AqYZYYY4J5+aEy8yapF6/FM1a6Suth+IcaH
qK2/LJaaLRIyJot1mZLTnWH0rAaWYJ6UFhF+eg2pZNOfozmymAqgt8WkJUoX+L2N
e+kG4Tkxxz6ADhgJrBgKbbKUfltyd5W9UoTyTdsU/OaCWx3zz87iPrcEFPUFFj6r
jfsA/xjGcraO+maz0EnYUqs5RLkJakZXJxOIabj1Gl7y5/Mw/ZT2DBINoKFMvup/
m56rkHqPxOjO/kTUtxvP6khkB2qgiDLql3EJN2iBtxB8AvfXGJH4PQ6UWPOM7P+s
3bMG4oB/mqQu74VmaCGnM8lQwg5vbbXCjE1usEwo8Qqr1T3l+e6TOXUjY+F26Jup
UPGfQdSjd+uWYXH1XFXpGqaQXeUXgDeJREITz50b7s8s7xhuT23/mNHFzZqebnL6
lJlHdOjYCQFoeccRoC61YJgY1m6+OiATwL3ZIG3t/vkSrwnCg7xXEh4Obxx2vTVW
q5ph/J0Voz+4tDk1vm9j2fYGQdYAme0qBXXgfrxWXbbDrghlRvfabUwpiNNXHMT7
ZlUcR/VcC8172gFb8IOfm8HZR5ZfOsn+htKiG0eZR43cpL0Iv5kcD1d0lYfgdCL+
tfT2MMOvoZLrtWpZj9GFyYRJr49yqz5CaZ9atlqY9/RDhXdecIgM2PUN3OF5AsWi
ss95SPPQB5WsyvB3taxfU+Mlw5NPnF8LhF/dS/KttQ6bQ5kPhpRx3LjZVb8cUQG6
Z3NZXf809Jz9lHexaOLhfp65lGLV4JuWdWyeFwlWp/GmMuErG9XqK1HVsqK7CWll
aV/Lr8UadNliGGNRYQJe30havezHJ6lWA2RULOJMumGb3+QSM4vCScWkOsAtw2Sj
ZF7vZAE9BduLI1lpWREgKF2DfKTCn35woox6/Y98MCFiRuXq1O+zhbgahyVP45q6
4ssEk2UM8D/lXW2K95exyGmfLWojEAM/szvsoDNFVbQYxqFt2+vwg9NvN9ECushp
4uTYgcla2pJGzpWrB0wJ6bXrd6SY5JhsHFlY89G+B7cbqDHo09fStUTkCW65ox+D
NPX2yaeC6am7gPboq0KGQjDXY1hgW7zMVadA8WzCpLKy9Ph9uzKWCBQB3G97+ur6
jSsTNshmvCjjGa6NovyJWGDgaLt4dWs6kXSVG14WIURicYny5lYgEt1Cyc5X58DV
0GVWWNyq2UnFLBG5uKPaq44A0dk+fcoW5B8Z+b7yAEsf1HhhqNuYUrHLvk3i5Zvl
FcJAQix4muN/IPqvPACqg8xjEWQIjWJkCscx+aa5/xLaJABbdZ/hje7WkmLl0yPB
IiwpNI5uFV5/JHIpeJNqCUXnkMB0Vaw6ZTRAGLX8ry7pO0hGSszgW09KvOywGug4
0sgfSdbscz0znGi4FeGXvk5dlYQY7bTYfvrAwhvEbAadrl2i+mqvt3L9a4qEeRD8
ZM1g18McN6xDuOmnrb+t0co7RUMDs8ZavYynAJcYhrHG1ns7yiB6crGDX7YBBA9g
pzJ02pXVHCsAAnpbaDGb/aLJr+JSm2k+SnpskgVvuXChxPVSAuR7Y00+yDFPaAQP
wr73H3Q3AYsy8mZgGsUmZdpPMmkXLkRckleQu0IeK72gRqnBR5z1URTeg9AZiDUh
OTFRI5i7Ux/AUNTNnq95CvgsPigivpkfh1VlSbFBqh4L07FEytl1StuIjeiBfOhb
7omDQODaefSIKSTVj5CLlxHs6SlNESJGsq05brUMd+7Uvfq9jY3xcrgW92ca3QkU
rrZ3f6BFpOV7mqAxyZhvG3CglSp52XKLP0MsdVnJExy8/ubulzFWj0ktL2joSL6S
JBJOHbe50e/S6cec+HTbaoGNRL7isUusGBHZNzyAiaMiQaXQ7QXPYY0PgNkGu5K7
zU4yj9VfqBRMLL9rDIx8NoxCMqvW1ZvMOX2xxmhAV20tqrY9U462wuT+5C9TUD/J
k7cRQsjknzX9Ho996nbDUszlNYOlGVkDyqkdO5DzEntM7yPwqCdEjsCb99X7B+mx
3p3A5DeoR3AWFgHiVHoBeNDYzOaJbflzUa5VNpYkWo6tfmZzcNjWdTYMIouovHtz
EIH/untWxwJt+zCNq2zdR2fLHp0sAPsgSvxZ0QeMpzUMjGtab1zkJhCQRK8EPt8/
rWJNNGVXjEt4jaFULVUhoh8tL0zvaVTqdnQ1TKnNn+sg0/3Lhfoph0M0SF9nfxf3
osMIfUzmuq1NX0J8JPq0PauAXDmvrmpEmjzElxiBZDb2m3JUvToNq5srCSXZZIaA
LlPuaysLN9YFK91sEyCqIXcjQeIZpEQulfR9PALfNlJNSMvg3aKqKfikQtK8g6/L
WEuQVyF+HSNaPeEup/7C6cIWqHg9vbD9n4GCJRk34kyP2TbuoguSHGkuOv92MKbh
VmA7eLdgncS7mi6wdGcCREQC4uZznP1nolIE0TMMbqRc3KZq6kGzc3TyXZqUa+mJ
Au3zQ+0g3+E8wxWiIwW1H7U0Ivrr/2g0KilMWQg+U7eyDSXpWvBsrNvDSGyBLMHd
AWz54c8SrK+pmHYIZOSqyuGOp1b4uyzFcy5HQjD1fYsfjg9MBXF8X4jAOuWbpNv8
7eXbcK5aBZLqkFGArSBNHI3Nu9T0xv3FkR9zFbsJdRmUn+VYCM8szg5VeHYbo+Ax
eUXgpaZJ8zCpSDpCbdLjYjHjwdDthWqBuY6LSrYq0i+4PSdrK3j9aetWObYTA0Wd
p42OQ9+KI5RyC3VjudonBygpCyMs1VumAjGYx5E3U8djUWa2E5/BKaq5eXVPGrq/
EVLAkQ4juhY0lR+q2od3gaff+rfjcUJTeLB/NCuAvS/yFS2CBd+nFrIKdi/c8SsG
RBqiESutrEn1kJIpb55MZ5uzLbv4NP4y7VLO6XIPp00Ko1MJ5P9Hj7rw/1OWvIMZ
KzRYUo0b8ojWSkx9de4XNB4KIucXEg1r9ug/liWGLEKvcmF5CCmZ4KQ3S0g7fG+4
FO71AZlyj0lbwgU1fpG2T4czqqneffQrSQe9p7S5m5vUqX3TpWwrlYLrc68Mi5b6
SvL1pWUY+dmemwgT2RJi2OEjpBlVvKNTD9jqGyqN8kOqcJhn5ffsYF6uZGZf68UN
py41rM45w51DThjTRlqdr6m8GhVf4/wMmBDxYZFoZzh64NdDbsA57phtOmtRDsP6
owK2bmUHxM8tmAXsanIj99JY82b7gjjlNvJscmreXwdkgsTT0m7jnrfutNsN8lSy
WVvRxrr3NaFG6Loh6INhP0RISfwO/gDs6u7ydrBOnCLfQM9th+eDbkDa68hrpTqF
QEZYY4akOqqLy/rKUa+a2n52yw3EUCmgWqiQ/fHTneamNokEjtrleuCNFG1hDomX
siFbSdx/vCkAJ5oGlPsM9MbUA7jONGXSgWf7cOHg3LwK/98m9+NGhGfY8tLr5BKc
6Qbr9diI/M00CsWBqV359XLZEFJBxRUm4xQoKNRiwv/gB7NoKqufAt65skJLhj27
9pnQUcdHHLLreTSH+xwCWmcw8ox+5juKNt3kL2FyzIAeBZbqu2s1IU/xMI1yL7b8
BABumseJm/pcuu8OXYaGUq6ctjBlH3wB559xVDRI7HHJHDdJQHSwfBlqlCv573kF
+v2TOUJWYS2ebuIqdklEZ9gfudyMAMHgns6NPwTiSCZvDJw7fhpqk5BLh+tagyxE
3DNcmGIo8oESFhGqamC1uXMPZYu3nuSs9HtuHSxAFqAds3Ara5vj487oFT3ssf/x
93a+MmFI9yXw7BZtJM3w74xZGF2XNRQTgb3bc6qpqgWAr3h2Uuu1Vu6gb+Nwq7rH
PxgDX2MG7eijCoD3Xv37VkdRiZu/I3xCcHyST3RGlP5Dl1iAgZUnJToRqwFIZqJL
ZK9Y/UJmkH5eAPJztnlKN/D8kTLl1crvvK6OvW1HVfI=
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6848 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
/GMbQK29Y+AAYqzOrLs1aQ2tVgDkcOAoodN49xcwNIjMAs5VdxPcPQQ0klWjGKJp
xMeHS6kzH5CZFMRJZbh3/ZYObn/zICA108TMFMpu71O6Z+6rqNe6SG7uGBDAvGMG
yOcFtC2tNtBueFY1R2HTQ5SAwgjwV1qXf9CSLlA3N2OI9fbCKqc3VguxtuRbNdUI
yMVNxMfuuoiqBecX2lPWjvxF42toDBqxcC8fArWSa3yVecYfB3CFzYlbZLyFYWuL
Mpj59rhvfCjmySyQjUbXMM4J/kbnrwi56Tt52HcfwGRmqqNJSfbwVsPbPYzSJV1O
v8Pu6A7etPmU1zBhYeMjj3mAHN+VG6s8573mjCDNhRp5m0VERbq2vLtHCQlXHPY6
xf16ftK+FGGM3lurqd4nDo/rLlyFfDbeo03R2mSkZIB6bcp2F3hWNJhoIxB2AZzu
wrGfNcdfVI6l0GK8KCU8FDXddYU9pTxTnE64cTyTIQYcvHM3QHcc+FBl6MFS5cUq
nJFgRVGGp6LJA8T8bl/HqyAja0GsKWeSI0RiPrJpcfC2HpWhEwI7sLMTq12lFj7m
U71jyIHsmrmHJRugvtd+iSQQzKGAglQszbfcY1gNGmRT8PtydGYp3vVC8CGy2VKx
jtwNx4QXAi5NtLzrCZtV+vdHJc9Hu/05JJoKV/nePhh3ntwEjuTSSNYXtQLfXVja
PXKQUU5BfY2+7nbCsUm4JCrHBCYueTX2tWW8yn40rlGE9inJhvFZMyV1NLDTOdwm
O1NVjGmO7MTOa799BGytrrjWdn2LOhZllRfr3gz0moZLTcwRXKbH1EbxCQb+eO9O
rvY3eQbM7UzWmQ2vDwjx/MmEsdkNUJ724z15KJ/Pk9uQiljvdJfNcUwq8CWV3wui
IE4tazKBiYo/GPZLEc2csfJo980ysaaIWWqyi5hG5kTBWVoJgV4ZfaLFm3Ruvpsl
uNoEI0SCKPXp8PjVOGk4lkqoJHYtb/5dmVs/aovHnrwtiB0F41tghwro9PqXFpLZ
HzaTvIj1vM88hTboP0nOlob/T/l6WydQ6B1TxW4ts9A012K/varIkI/ykrGicrrH
3XqBkBGFHW/pfDFwJdjstWMUfR5c6MoprIgcZl4aLX3gWLeAtrFVQBS3PuOxnkQ6
ekz9p+Ujt81yNWMARtOVcUKJqgQ5sS2iL1GoiaZpaaa4fwt9gxBC9y6crwYe+KIs
ajFZ6s4s11Opx7vHvKgxyr1HBZPmmJlR/pVh2REvjVk3YcscqtW1AOoy/8jw9ZF0
jFeG1muWm3HMXgDiwVbWsGdspnrYDjerAPbuVsm/GdwTd7hjTN9P00GocOU91yuG
WaLtcN1RXlmWb1ADwb2MC96wqfL8JIx2Kbioh2+0G0kkgSEtOI5rXag2C9uQKAJu
6CAxUuachiDVWWCGGOdYbqcr42kTTIyQdoPQohbtPZweygC5bRNQ6K/XOnpTgwdh
LfVl2S9UZtRiQ/jwhBOrnb8X27HY9kP5E1HIk0t/kUcXnwpXK4OAsGFo7s4pVBZ+
5n/VQT+vHXC0ayc94SagxNJUMdPaTDrbE5eDcVIajBuYpuhW7cuWTuBZr/2AHQoB
c4yHZJQQwYFSO4Gn3enzCCr3yaLYH/yWRpX4AuoXpoMI2e/GNEcLUHc+2zdf3IYt
i1MwD/IzBepnd2zEXvtHjGfn154DAdIUvViSMkpTlnL+odrL/idMbtkbbKZ6g/9B
pr0AW79kXvBbhT63zAbvqhMg3LVumDir4yndposbYlsPqKq3SdfbjT4hlEmLhofR
DjyJx0OvwM1XSr9ht9oMicpI/pC5cd1sbuLB8s0g+DwwOyRBUy8r8oj/96WY7WaN
EG8TqYafjSgeyALrflQb2/IdMGS6+yIbGvb6snj8jO5QHTD9z1CtiMIECM49jztX
5XqnD1EnXXBYAiASoXN+2LQDCvvtVgJTlNF07iQ2cwwjQtNcfCcbqdsY2/6EFBp/
gmVzc0ffwpmaUxEu/dHTT2ImB7dWppB8/h44uvH1t6WDUpU1ExQ/hat9WbCjd0p+
1ainl66uNmWhLDZe0jSh8tf57nBgN2mXFnfx/Lm8ZzoxmjdtxcnMb3Z3x0Sq4mKR
CmjMGTWeoQmKhcZmMfYwfEw0VX7K3x3yuXtw8EycLfO/KZiFkWKKb0htO7TNi6mV
ImpSv0o6TUUFvgxIpBqwDdcb1mn4WM2GHJOBd0qNRbfqrn7lybZ0z7BRIuycuoji
7DZCUk5qSpdWB2vg40Me9pkCK0WSNLOUwWYGeiVHCCqfUqJK5N5jA9+Ldg3TgUwS
V/0ejDQNEoHsT/KJa7Q0GNAuUKnDDyRqBAq5GOZb7Fj+jNQ1sTOSEQ1vLXXDakvQ
vi8QzQJuAMda8EFYQKudTLSsJLVdNM39WuXjyMAySdkGD28H9JD7PqRVEX3KnlBx
oWG0CUIQQcNRLnj0PR4S6zYt3F5HVO16m6d/vj4h5yB6CcPDvtcGox0e9XniVzuq
/Errf/Tq8oYJe9uIp6J9wDxoO+Xb+nsaEUf9nI/mQHfh7zSZ9lPzF0xU4oy41I+S
j+OnbXm4jozextq+MbgWb+lsHQvDarxyQXoyFDcK24HPGCReO5LTWSasfm73cgpK
apprnXxvUcUUn3Q6twJmXKJnhj/zT8e2rPmAjhZudyIDwf6SyE/fc2Uza4eKnGrx
ZRMjxaPCSO/ROT53lMPnrfRim2qZTo27pnkoXcL619+bW83Gi3lYvE4loxvT+FWV
OBeK9/lHJKEgicmKn/s9XBG8WjJC2kZP2QByHudS8KRZIaUKYCzOk+yJsVr3eqXP
Ttme5jv28qZEp7YJyzFLIHXg4kOwAqXMSjjo64HJ91sFmyseB4wfXjqGzTlCgfak
EqpES2xCRu5ki8DMDyMcBFuDZ+eeM05C2bzyaxq/xq4tXAhI5QRe2gtml/lfAGj8
AJc9AP7AAwEYqP1+h4HydDBCqkL7qQX/A6jToYDqgtX+AgjVw+5fYt/oGrwXiFz4
kmMBwdrd7nalHZwDL4ZrvuGAuRaJq//gZk/TFtxDQQzr/oEr5YH5E9raxs/vvrQ9
fCsPWC4lKEAYDgpU7OGJ3p2Ton555rryohE5Y5lKHy6KLFwk/Aa26RLWOuhnDPYG
zOXWoTo4n5feghS5MtdW2b8vW0bgZKx24rz2Ey7wKOK5SDnwg0Z6WYWXSz3jsAP5
Xuwe816asC7sM6uUT5APFoHQTgAPutDWetK0fM86LUBi+T71Y1QQj64NluhIOzi0
KmKbdnbZ1HxVKCQhZrQv7QMMvVgV3FBnoHubmLKX5kZ4DlngVf/HYurPtp5CAiFJ
2ShoW19N20VwQ3tLAPZssIdpQaaumGjwgSkkU3bVQrhlKIcHh5gtRqaVzQvY6PSB
VfMCs3ubGa7oXsNLFk99cvSm8l2FB/fKSCSWaZjcJ716H7klWNiIqGmQh4cn1a/g
yf2LIdwUPSkviR3oGVb0y7R6NyLuQEmHgW8HSr2ZBMe9q4ICNSanM28A5VTGdJBY
L2vC9phDvTlY3Zk7HU65pRUQ+LeYbtHUCnDa1tVhE/dGA7cSfhRrfBEUzJbPCYaG
gk58fNnHXC8vWn/ve/ifoQ9+FRB/5KLtjffkrFlwZq2FM0u6b9NcUhwPF89WREfy
IEYWgo2akHTwhkQ1t81/GnYCsoJKa7Fqs7ZB+WPeZi4B2TYu+TiGXNBYcB0UOyEu
TjHNQcDuj815ENvzefxNqP59scvYAtW+Qt3ZYdNW5XHVJnK9n+NjEOcBRNMHMig3
II1I+8xUEoCZ7NIW4S547iQk+Sa8Wcv3JVw6PqcFuzu+j6L5J/zFWd7AkIapFp+Q
Dts9xEKO+nuMXSPYCUq92eZO7N1nXI9ajDZjMHspifPWsOKiVW1bn72+xcmJX2fO
2/y2xYzawYfPC5rimAZ3VAtVzk1VpEn0QEfOtK/QXKhVH2OImrX+EQHlFgcrSVbj
ghHxqggl51ayTkQQiefyE7+lsB6xuZmaha/ALnCYdzOEIUFU1qBf0Um+M1s7+any
cG4wSjNxcIsY3DS+7pblykZexFiD58FNugpMsEhJ3BtLnlPxRIowyA0QSkGN7zmS
HLNYJWaJajoSjqiFBsc/oMR6mM48a4D4Uht2S8c2kxnHr0XkGgCDJOJ0kwXG2Asf
WK+CFQ4K206/RXT+W798e7EwsPO3Zpks53dkPElG7VW/qwYWzuN720bUpjlgpsq1
0vqVILa8ZyiNVHm6v5QJoAnTwGqZ3XI3LuD80Ht/cui2vvr5O4cV6JQq5ChvzUFn
ik3v4bjAnJlXOO2Lh8SCjIeB4or91f8XmAWPsy3MRTsqgKHAjzebZmyQPzls496I
5By5vuTpqQFdIibCU8jfXsC5T9n2MYyypJlneO8IA/axRP1qFQuLcXHWj2s5Ybne
V43AFSKYurLRFkFBkOn0ksEBGFQizNa90j9Ytg7u3yLLJYr/YeoJrwrUnrIbfeA2
K1i49lQowb5U+w6GqH2kUY8SrO13iRxdfyONrTrjng5V9PVfxeKl1TEC1CVKtCFI
86nVbCwCx01VpWjwY07xuzUGSnPuHChCVawDZgw23tfIO/sVRU26k0DIIohFXJlc
EfJK6Vitvd1pDm9Bjd5bLnBAb7lOsd/49g1MoO/LJI0gVPsEQ0qrYNlHxIlkeSV8
otiuKKjlPzZgCWsydhQL1CjXzU5QlkdzY+63oq8LA93qT8sPDmH73Mwv6eATuHBe
3iTzNxCcNkN/uITZUYG6roVsbFizNJJD8qF3FC2D5E8rJ6cP6eH5UZ0wiRUnDh8m
NctkycPYcDVqfjc1tmxaE4YzJjFzkmQLyUrYEQGhQ0L+/8k44csCI2IGBlDxEVBF
0W8WUeaz1yXcrCvNC/aaBH3qBoItpvA7LYCDQeUFFZ8/lV2dq6VKhGrZ2bA9n/xw
p/Xy6gZ+BEvjbG5Av9wicYIXsxdFQWluTA9lKpFnHz5jrcTcKGGciQUaAiORpZJq
jtuLhzk+7T3Nma+jzZ2xYHnvSZ3oohpG+R8FmE6j6wYQcC/uipUcqWSp7TcRyEb+
qI5JfSYgbULw4k9txKsXUofxbJ1/UxLCm5AVU5cUPFtKViGPHI7DLds3o9c0jvEN
ZVrFrTU9rt7Dxx+3dW/eRpUzqrBtCjRJKljeQ9Rr5MbQ3+SV5TqKqu73CnNLDa5z
B4eU94HkvGTe8QFoVErQxXvTZsjjZ3BH+n2CFijaJ+SRcbLJF23rjD3ljqJjHo6W
CAuCRs6I06udsLkTZFQk8O8ETyIScSGuEta+Yu83HpB2bOit+hnJ0V6nLaNFK7wo
77NkydwVhbtQmZZhzB6wI5aUG0wqvrcUkmZwE43yhJkIz6NO0EL6VxoxEOZXZo53
ZNzER0e19CGeEEvZDDR8DomAARw33YmFXsd39xVFUBzJup1e9ZOx4O9v6+4l03WZ
u8THVmhcaUzRM96lLk80k0AAyUMdk/vj+bzkIcWHg7rjbjufHiNz45R3KtfDn/mh
Btbm5gG8DLx4dYZClUKRPqS3ZewTM5fwcNYZhoIDpCFtfgskDzUSIOyoC0fvWMoe
g6EDMXz8StISYKtg2+bf+FvGuOiP+PHJucHXMieJuP+bathjUx8ZFhL277ALxlxk
/VdB1bdibt+EQ+eYV/0WgfxVD9a1jDKwKbf/kikpIIKBLg1gLaMjs+VzyNk3dC6e
poLxTjidLYw0/TnPePvt0E2xj7XyO3ZVr5dwht6dEE6kVNU6NlAwxFMtoFWC8JfZ
WTXAVVfArX8r2WKDUpaWsXcWBfh9EIbGXDmY80Gkj9z8wuYp1pUqDyvOZyoe2Wkd
hawB0A65pkFKrN2MdoGFQFT+AaFOn8R6eahGLxyW7tpbEIcXqqtsSXOsGTnMhKPK
tfbHE04kfmnhXiLxsGJgr2MmkcrurCmmvXJdjzmB+0HWLIveLT3DN5vvWNo2u7+/
LE+IYJhLdDetokPFx9LUJlNcYnJwB9tVkk930TEObQmC1H0/U+T9uTyGY8n+SKR7
tKJw22IgShrfhiBRB07EsIqxLt9iJniFJnw2C89/OTS6HomFRUvKyr/RAyPBEy5I
WEWBqE01bdE/GjKeko2sYRLxehjqNRpXmZmJC7FQNdm/3p2cTFDij61RBR4Rv4vt
LR4+tGRpfFrucxyrojj6Q55ajtvqZUq5QSvFvARwZxmDJqlaJllLJqjyqtNuyEy0
5k+LPXfdROjcHpiQ+/i3MvnUqhZo8J/5Eown0jH5w4gJ0EKKe3TZp0tAG3v86GQ+
uVfi6bRFI+SuTHOATFR59uuncHGHWG16RcV1PXFTf/zfEL5rHyI+YaY9D137FWGo
QqEL/mwPSCmtDKH2SRn5QirwjBma2iSLo5uZjs/pxjejBxg4mk1NNyagf0avGxI6
J3gvl2MomqySWZjetxiRmUgfdSexe3dxiftYauSDI3G/HsM+G6FvTqr5bl+r/qIv
uwCDSShSmUj1z7QZdJAbXNa6Ljj73shA6QGZAy9FIqHE+xRopoYU+fWVVLJKlEDI
qNmb+s/EK8sFM8Tdf3+v1r4Rrve3xhHZEViUmED75DB2BDM/jH7TalIBWeM6B4pp
sOVDhZlVVu8CBfpsmU77twycTZZZJLauGszaT15EKH3BaYblXgdRGA61lbVb1oW7
ZpE9rjLnJo1mpMifujKJj4KE42+5sKSnRWVWyStTwy0Luy3kTXKdlAFT2vaZO3c/
8GzuBlDRMHNh4fQIxjDyUpBZOpY/8NJTazeGVauF6Vw4YORciocBiUHaX58bmWVx
q4npVUClKwS61gOoHwfau7gSIRV1mtYd12NbRUVnKP8t4IMGPxc0vBIZleBnqP8w
f8G43GnnPw9rUye7lI7DC4T0xO42HmIMEY32ZccH6luE93My7ab6s+sySxncog0J
FH1RkCPomYJL4TCGGrtrp4A0tKmmhcuHd/pqkmnLyulVHccEVUzebME51LPS6cZh
1/3+osLf/4FRbCsduWO9dzbMFURqL+jiEX/5tCcs06MDhKDJfRdfQTxxxuzmS5jM
R8EAkFQPnpaXMRCTye7+1S50UVl59fPymP5qLrLfZ4XQ01zYM/sA0gQoYaSN81Dc
6+BVjpi9J6ZdNjCUbijV8AWk/AnBiytWV2zw9kxEn+OoOdfJ4+F+UlYPXBX1ssPu
ks1oNuVQh4bc/zAbA1Hzi5hmOUNyukAAHp7gdLDJiqUbBXltUDFYKGdWUQgRQsLW
s3SJRTAlOtyr7t/bWnhU9p3OntMtI0JQrFp9CLPy2J0XPi/BdIEcC5VjwE37fOr/
qzUTc4qjxjiHJdiLRBOXOtszSv5ZhDU3z3tLv2AmON9Me4TjBIFVBgSnhO3ODmhu
5+atwWU2sGSziG+6I0Wckz3h5elmZLViZdCUjG2rGU8n+flHyagtQk7tbHLqhunZ
wVbJNe5IPua7OGlkYKvdkGWr6blTr1Pej63hvr929R0tDfbp9OkvE6T9NR3V3Oyv
GJnqpfYqzYRARDlCWyS4tWSH4z59FC+VmPitVXMAB0Up92F7iofCXyJN0DHw9u2z
4yMlDVJ5T5J6Zkg418ZC1ujNeEDZeTTc2BSXLwSJjl6xak/2/7My6sy1f0S3LkTo
Vxo6cqjwJR9CVQUw3MmGzSjURaVrmwp594flqODnrwM6Ii8u0bl6X/ywY7T67PT6
tgIi5a0yzvJDAqtg0HHotbpROHlYXFgife9e/vBC2Nf//hq3a6QdzjtdrxqEGaBR
V4pOf8bkUHGToIrttVmD+HY9f2D/KQwzLya2CC8VwzHl5NW5a0qDfHGJD8xutwGG
P4xsd+qalnmXPxwvh187uo+/BAeNCXUu/DA80kdCQkb4LHys8JxPRW0spQvsYORh
YHHiqh6vXVD7YOYa/nvRnzsGyubU9pjdcbDNXX0Do2xFYFIidWNEsLW3b7L/q9N9
wzVuQ+9RrfsQdjRdRxTVV2UhAHNQuP5eLeFoIuRLuxWiwTVbW3eGGVpoUcDVGUeE
QzYp1haOh/DCSkmiKWGeMCvhB88hiQjP0CDXJhNUYzPOxjmK/d8mKMeW/9YX1+PE
IvDrcKiDJwdT/G/8WXsRy3SW/8G6OVNdawvzwqWxPdeTp+Plq8wty36fWeuJNjIC
0qTU/LS8N5+1Re0uP9QOJlHtfxPfSM61bSc0T7MrAa5ujefo6x9kEognzCSTQX5G
xS+aJJFNTeae9VX6jVt6gCFxb0WQQASIMtFUHdM6nN30VAuH1KNEGYqB7lh8zQ52
bUwhByYAI8GSjdpsH6NYkLVe2vQYXp1reBtfcpwyMcl5x07xEduS187F43Pad5KT
9sT67liy/LwXN/EDV1+APF0yFgDslSly4YS21WKZApxEv+eHN2m779RWNCfg5J0R
lTRH5ML0NUvCJMb+zOyyucmJDpoqsfYzjioLse5szH6roavrCTu2YmLqRJ5VdRHJ
mewuspnPc/qii5UT6Ys975+9ZlAW8/uM0PVM2MiEmbSaoUBu6zsPR+ktJIHCyC/p
c94KEIOhH3BdiMBHTvFnzeJphUvgvFXFexggdvvIY+aItIQm53NZsdur8j0LN2qq
JbtCDhhctb+uBh2t/X8DnGK0G47Mt47SNzz/oAhNpKzsteRvt7B0m6xVVK3ZIQNK
bNvOgXqeawN/SlImf7w5JfJkZkolAOeeQlcOBqFoKRFAMNrxQc+vsE1EMk690XbY
DqIAjbw9LxY9s2DeRCDIXZATEX1AMNts64rFJXMIczbyoY+3nt4NL+5cgEGbEWIG
k8rRfFJNu2znPIjJGb/D1zG+eBwyergUaRS3/fyWIQ2/BB2LZqzxIUM6Fv9ew2Ee
rATFx4KbUFcx8NS2jV7VPEpqAM+ylIp13vp+iCDrx12Ys7zKwBZvZ4Iwag44ZB9x
AOCULOlZNN5wkHMbTYwSwh3rSCaMStSEugFZTkX82/QsD1Gnbio7uxGLfr8liWvm
2R0IMiGe4q2eIElhNaYlmK+rJEvQdZDb7iMg6AAguAM=
>>>>>>> main
`protect end_protected