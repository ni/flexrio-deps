`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14192 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
sTHDbAcNdRVMi738hx0vzs8FhHEQ5k4Wl80hlbK9WdJWiCnClnXV/+X1vU882uzu
Ya2csqlX4JVWUwKA5SPATqHdfNfTmtILPw+Ixk71kJDC2t/gfWtrmcv26ISiacAT
ycOI9heBqRmCZKGzrZltHUTbma88r/9yz9xvN8W1RUsZyhWBttB3Mv3TXTvcQ4m0
0KBlrhjuJYuQLg+2vw0C+aNxIbLgziuvgJzqs+Ov+rdmt8cblgr7JK33ygb5wZEd
m/OgElbylLQ6oj6EvLpY+d3UekSmhO+N64yIj911RF4CD1PPpIiYNKJH1Z4jEnbK
NEqQMD+WqAxf4YS4hyxU/3nXFfKFaUW+4LLKNXZdwaXOcWb/fvcCYPm2iNwQDm0x
UntMozxYZtwkrg6fDxmhYHln9tdzqj6ZjYJSkOdbBWbEn9LoPs4ien3P1YXRqin2
f1zjwY+OjiOh6tooeAL9tVBu+dJwKZwuYn2IR/gR65cEvQiGQN35O0Vz5NPXy0Ww
NfunosxD02hkXuAfpo9YX+FtZMoCIWX9l4WYSnhALxsJPDkxY3O/PzSUloY4s3ee
PXczLQvbZFOq8xdp2G2wJaQoqu8xFXFiiK3gjF1P1vTmtbGW3SgvB+TByWcsE8gX
wDVcP1J7vgmoFB4+h1As+E37L7j1YCo72U1qFWVeMd3p+4YpABJE49Hfj9h8qqHl
532DmzFOrUesvYTi5w5PWJO63lu2G1B7V7GJuvZrNNYZ9njEBqHKH4MlMAdgRE0D
uXmmpuQlG4lL3IKxRmsJ0XKZJ+a4ZGRqz8yZEZ+ggi2CK9XkXQ+hjTqtcE6iYeTo
vfaf2THTbXfDACMPHm9nx8r4qnCaXiFGf+Al98rghLoAcRv+SnLSweJvSBeFZOQU
Z9VczGpYw70qMkrwWazmwSL5QGruVV8ZSdFd+U5DNIf0oq8WCCZ3ta40B6k9T4QD
SvHJZ+IjR7U2ot9JiaF6ALhEygLA76cU/lPEhSnXDaKhfo+3az/QcmOnnLSlyJfE
AxfLeSk3orA60qmSHjL+BdYhKSjYvfO3GyDJz+lHcrS+G9Yri3juA47TnWKgFDqE
Z1SFgxEWf06UO1KtskOOfcJxSzqT+55l7DVbbqQzwf0JZL/D/FsqppEmNTGxPSGQ
/ICfK7ps8b7XLPmr4GonpxNK16WtjzGho/iKNMBD8H4Hn51EDLBpMTokbbmhTsyU
jp4/RKh29rrpA3c3v+Vqzmtx5+lVJD2l9TwmxEf/MBeocQLzHkvQS5nxHDC1aS4X
/O9GB7iPG5Rm+hvHTvQgHwLskIrF8ZdzMcHxOgdw294SygwG3wM6sYO41uHLvRSt
3eb5EAU/TTMJi7S33RI1udcyWppqE4B0l1QmjxP4OYKcwVur5QZIpHVnePvRh+tB
QULUMtIPJeWQ7vibC5xez86+rl1cVGiZXg4toQV4hLo1bMp0frYDbdY3mkjEpAye
L9k9MxC1PagsEggZkE0H0uHBLizNLaKeH65qBWpfRTRtxBwcDlSKtNYL6GEIEW71
I5YI6EZJRgZSsRv0htaWW00JfgVY53H5OEkYkaKo1cFPLM6q7QBRB5WU7bMShhdJ
N4L8PyNP7XUWj/KKvStp3RejLbtodfbuAJ4o7Jb0d8xVLMYESQdKMWnoTLGtAQSw
K4P5vXIi4GRoA1vOX3XzKsZ0RcuT/GrR9LyoQJ4Vrzfn/9+dKaC6SJ0bpkA5tTUy
GmZTONP9mRYG5shsjHAAr/R5e8kcKdI6vdXVQmgp9CiW0AVDeLdUfmsXAiP7EvEB
h94T44ZhsSle6jGx14lOFp7GB8GKghDaHJ6GEFkGiYDdzdRQhybURLUemE/K4xuJ
dmywgjKGfuMBx+7HFCQ+Ka4Pjyif3TUKle2YyStAfIimwfdLiV3B2kyH+27zqHqD
DN6JRJEHSyTT2bke3P+sox2E7ko83IUHXTrKTJPt7IeNeo/f/gcG4WrDvb1T770W
R2W/F1wvC9V+01OSg9Vj/5C8Og8hvhF82dN4udr1KmlusbcXFv2w/5wMM4LpMdfT
AFFL6zK9diS9Xm7dMjsGQ/LV883ZXfFZPi7TtWmbUfFCHthC+b/TEI1Xx74Xdymp
L+CGfEQzgBdGCYTzBcUOA8aQmMIu5q7pvJUhnxzGeTRk/5rEEdbZ/yudINnTEmH3
4/I0E93j3qPbQKH6/SiVAL7FY4iD52BMRkanyJizlGc62kx10ftub2lRnrA4mpJE
ulISyiG1UGDRMTvtRBGqQQWu708I9Zi8ljTTzORE6XEEuK20aV45Sxvhn8KduDte
kAKuvIWgqGGv/YMsN6vTMuY4AjLY0yg/4Xqdl2GwZ2bw5kvtB1hqAeGghateyQ51
7nVW249OG43DtbFzkehy/DUyMRtjCQPeJ7ENYR8PddxFm4YAzzb5dYcj17jrF8nP
I42s2b+UF4w1psorBjFv2bYZAZppx8Vps4o1PSNPygTF65SWcU63k99nC3fUZHCE
LawIdxNGiaUlHUqQAurf5X/O9zhTaqIWebBrH5FpCNELjQnuqI+W/KuwBc/3aoN6
1ZPKTiH/oI5/V91Mha+O3XMnKsqC0MmbnUK/wvMv5UmeyCwBw3oXtj8KI+cW4HFS
YWKDCDKS81sgbeK5O5lPrJwlSyJCZkfxyJYoGowRHqilpSD9OJnDZvHZ9GfVS1Gg
+qhy75ydqLVUnZtVv/qJOWrw/64UxWvjmIqkzMrX7fOPFloMFFZdIYFe8xJvypsN
uNEDFI+7dN19PzYNrbCbzx8o16rtRgLsG7eAStad+Or3mUNIK5wt0jwlz+2vEZio
ASC2uei1QziohjEqsMj0J7xQosBQQznWWaKoVdrsFcnn05/BbEzJYd597YnbSVqT
cq7KpwCvIiDAbdQDVRNw34BYZ+0eNtT8L4Ru6OM90aEHiZ+jlrk5mfSbLT86F5l6
MKa3d93U2QF8fF6XlNiM4teqCkyLaFE7EkHx+xg6HZlKOFojcQM1kutIxBcprDuE
nmY3Eq+fqZhbxJKa2n/ykMGGX1Ivg1tlZnQP9qxABMCHQrRFDW3i8HXC6CDQYIEo
r6yLAbEf5THXHmUaa3tiacUPFybGCKiLaYv4njszwhRWLLENYYoV2tKohRYPnFE4
3vNmz1Uizv7UsXyAZdD6SY0dQkbVDebpJy6Z9HVnNUD8SKh8MuaxM8Dt5gy0etuP
RfC4NX2lREIzDOml/0IM7jiife567k+TQYjbMi/wwt5QnUAkTfVW6oqZ2qtEt4Vh
ZQ8+xIzr5v5EZAJsf+gaMFgVYBrZFSorje9O4F2Rh3jJede58YNDfWab3ocfcFYg
YvHAOswVgFTA0ESf4b5HO457pXUyGERmRsige0JB01le2p+EbiZ9k5TLSUBLj92A
4frQ8Hg194eO1as6T1rOrtlhfRutwqry2Ba/D/0O4oremjbPXz3zrXnTr9pv/cm6
HzHDbATiYfziB6P5bEvpd0L+f0dFhiAYtiOcYjjziD1wncoL6PV/9ybJu99aRoOS
+ePiGSLDuOyRvjYX+ort9AD59EU8P4aspILYv9N4l9WZsfhPn9gMCThsFJdCspDa
uusB7KSng+nKscLS3CSj38ddrud+Iimh70DCUhX90Y4Ok4LNZy9/hyDO655jH6Wl
M+nuHm/zZBYJB9ZjPk0HFqlERZ/iypfggKgUq/dixXCAG/s3aT9P0npFGxpp+63D
uXwojbzIG8bzulQG37pQi9VsDrNH4mMa3R2LwlJrAmMVrZDyYWWRjh4VBOE9UBwR
T3W8zKi4YQfasQhtsF86vTk8LkQls3fbzPa1alWnIoasXQwUd7FnPBuOUqCTooJ+
Ful3yGqWRkAmk8Mg5vzxy0f8XbYgz/Fy7JRjgDws4xH02znXqMYqvsVbZzGNRfNp
Q6WogTFsv1/x2uItqm7rLJiIk240+R988d/sNBjr1AG96L9qC7bgBSsUZieBkfHV
SzVRAf3+BL2tN74au6edtUxiey8ka9PQJNsQQF1R3kub0I76V5oXDp/NSSBLhqXl
pNtnwvPz+AdZmh2sSNkOakkFvM3kDjRy9W2uT7C7woCTQoBY4KANYLqFFj/bqMko
DlCYsBiOq2aw2CX0SunaBfS+YwNpQ4Xuhdbbb82nVcYo5VtLity6k8RzXKWygCtS
nyi3wnbVA1bw4N/F1EkzP1Y6vJ22LlL5ncWwv80G2fDeRD737nbFPDBvK+xCt1Mg
7Kt32EhXDV3HUWgKNNF+T+S7OgzIf60fnNQuvz+8zg64NoS6O9et9o5PL4I4xKPj
djPdocmQ+7tZZghERVRakKJ4kP0Ten04+6WNsiR9IBK0i06ZYTnZcZN7E5/x0khM
K+9fww5TdbxHQJhPGPJjliHtvb+7csDCGzh1uwK/yFyZmogJOWF7hONnPPzvnhMi
kSkdUeQgnqsgyxUOWRvw425Gh4lv0WC5pj4iDisZOyiLgVAydeuu63nkMG8bVLnC
NiNWEkMS32qrweU8iMK/XZOByTnmkOstpdisWonTXcM6JLMhL7lK/bc7fuibY0T3
xTpYPJ8nvtp9I+l+KUejQyv84LPsWHlY66EQhUL2FMUvaHTYTjjM8zTVFUx5Ya+I
FKPTt/7PYJPtTrZzphn6IQTAdRvt8oRqQgKPxWU1DY71+rwA/eK6A/C8Nu4uI84d
Wo6EpNbK/FFJsjNvmCBBSPCXoC2xQ/MI4m9y2jjeGqm3dsh9YtPRM+jmQI4K04yu
AmB+XUzaz9yHdFvkPmJkpY5NBupOf+qHHS6CAcbamTxeI7sRC4bw/wWOCnZe5tua
XtcLqFwKREZWJnX2nf8rjoxgPOfKHUPCcnluhYR38zZw8EOflO7Fm6x3sJc7XpeT
m/1k5qXdDnNhiRWZ6lbAa0291Kr1Nkpp0v8xBFnw3/NLLSqsJbucJ+ZtLzMBfmxR
jff+fwvBJCdawQWeyYMo+70xR4Gz8ZZ+yBy0YV5qrqMighY6XN10ZOLgxtoZGdRX
A4evF2yciXdZflJhy5Ri1jM0LsfURQIyY1LpJ6dBFWFx/TVDRv4ehaqVxSBh2ufU
EDiILohfGBJEoLFjsSy2evIye65wjokxJdTLgsn19PJQ926RTYBAxflqv5ZdV8gJ
wpGlXoVsaxPj007BPPTpThC+CqfDvL9s7SSI1I3aIZT8nflpTQaPjcTqJ8GSfdq7
KdImTz5QLNTG4amOcoyP0EPyVrUnlGvQWQOHukwaEXjda/i438AW2DPsEOyKxwwL
sRk6MzZyhlpo5q6mO6Ac1XUUIwkjCIDMyAmZmesz5yetvkVDtyVpnRLsIL1bXbV5
T/8nKUAQ3HYtCQqhWuv7S88wNR7QLlDzDuWWihC08uSHgnWKneXNytSeQtmPhKKc
PyJ4oNcKMTdeRl+knA1hU4WAmZmDVJ7f0Dq9SZX+sGizTx5Fn3GJNkBR/bJZCay5
eRYwKhZF+aQop4L4yvssESKHcaYeQQunivFa3VX0nboUfsn2HKgair+CeRd3U7js
WHeNEkl6NK3icnNKUgWtBr2LojNAbPoVH+N7TDXbJKcytIZAsqpSu1nj9l4wnkeL
sb2cPoD/qAKvdWzRDSvLaLD+dqUZwD2iDx+/G73E/KGxOS7DB58NiAna6m6G9snR
k2JoXVQGCX6xo/++g9X7yZrYnUtC29hu8LO52XkYRkeGV56hUFZyjXPL0GLfxrRd
bhDaJnZtGXdOI41M7YZdCz+zzmwBqSdVB3MxPzULTCZ8SIa7lY5Z4HxzyjXEh4kI
6nqkQKnrK6k54ekCQctDS/6HvKvRBBaJDCZVtFhpaPX+7nQoo5IBvjAQgO8jI0dx
Ece/KEn3xNLO9f6PdD83FLT1NEEjuAHHuMATNSxRCzRWpX5WUTNmU0Y+TNY57cKm
O8Ipkt9ElEZztQSxDj4jf7V4SzGBapxgmWfyWIS/7vN5PXzGk+w1A40K/Gg57b73
+cKGBYcYJaI47piabEyvUxjX8E/uHdd827aOzKagjeIN4UzQs9BLrJ6qvcK6ckO4
bCVM7BQYrjANPwj94V5BH4v01IXdMCLXJ2c/6kuR7Q0+4Ct4HiaSIuRM20Mj2jxC
nyGH5/k0+QNum1FkVLro6W/Ty1Tlr8Ya368EmZcogMY60e+pdDp2AW3qPCyfDZdC
VoLybO+Hr6nXYPzmWTQapzpmBTjbZJNWWvvFbUnjkegjAsjidEjDdEHl6F7toSNk
/fppgSo2SOhNbbVGdLWlJQF5KbzDzjr4JdCNwNBug3mwWwt6+6fbK0RA+SRqO1Cm
5EK05BK0VzE+skT0k/AyCioc9YPSiSLfrBl20RmUq6gggqpM3cJpV+BfWpt4H8Kn
YkGmF9YD6MFNYzoK1aSR/JJptA8LmKP0V3HM3peE8Jmtkzs+EG8jUIU4Qym6PpIt
QZuTaVOxyoDJE7majukXD5V/yRx8jfjZ0IpQGdGh0/JDPUF69WcaSwOIBHMW8N5a
dYsb1kE0hNtFzKFcpq9zk4BjtU5DUuq7DXT4IBsEoGeEg0BsVWn748q4pULAhtR6
92oDOZmZvhcEjiu/eMoVzPANcPm+N0DfCgAjFs5nTuYmFPIAuMIX5qqGU1+3TAF1
zyk7eIUequmBXl9HQpi5jLeQJnB4OuvayvoXO2tTKXzEa6z0xDTcIBE+XOw4B8hS
AEsSg0Gom5qiLJwmynlOnECsVMUa9BkRHthzpz+rnNTZIjdR2xo8xj6fS07gZMEq
FRdLx/lSriGhR/lJ0BtAsTQ+8VWzsT4V2mTI/5/Ma/ieWnqQTx7eQHlxKrk0cEwq
YGxMVxnLDWCmSmHHJBM30o67wm4HiHpr/yo/aRJqPyFFxnRvJIXGVJv3dtSJsfBK
T7tXn5BnozO4Xz1WIuSu6VMlSR1jXiE50QpzVq8RNkp6FVOhUvuaEX3UMdK5KO2v
P2gTLJ1GMQbLWdn2L0v26frMXqojvqTd4p5KsHEFEyjA9+W6csYfeAZG8u80QBYU
7+xQdqSl2pse8yiqlyfRp2hT5H0oXcmzK8Xoses0PcW48NuebPLDqVrvHWkpOY8J
42BGd1S0ODM3/9tG/XPzG5ZXHVUvgIzgva6rgnV+pDGWRdoUvbHhRIzKtqkkRxAy
CeSoskKF5vQAjcfn1+SZbD36hqxRfRPJw6YsukxiREEF6KfPlhwU4tde6JGcKNn4
AInxHdgDRUmPq2wrmiLfVfv+jIgqlU5PJiQ1OgcywkhM6dEqYF+Obl0IMMNvNBrr
Xx6XMg44iyZsfCRyAo9QRxLHhZTcMOT3oPAUY646KnPO0N1HRTTiWi5U2aTUDGgy
2dNgSy2ht/sa8kQDVkP8V0GGXKe26mxNAwm7EBBNhMFfPTY97Dlzr3sGs2ur16L+
UZYorCo5yNHKFaMGdIb27YnpYJQPbLCW5GN6hO1c+iHuKb7oW63zTUdUCZN0iu+R
tlbmt3cJLk54X3KVHWAhxFVPaOeavLSsmR5wTeGCdxd0uJjTAtigCkTctvgv++Nd
T825NKfcyP8VgKH+UvNHMsYqrrzKdEytkn/1NDBmcl6GpjxBLEMS4gMMH5nUHazq
VkxhGP5EsL9bOHCE4OpXmNgHhlKMoXKVn592pjIn5YEhzvbNLNBLeAyZvWUDWyC0
ECk0I0MUiSvKLXYGrIR7YMv89GOttavn+NqFZvs7JJUNGEAgROOngiHfZa6LxMtg
uq9QS0f6DRqgw7OfcDvlR+tq4Gzo2358iT9X/N4Su0hKdsp4xINzd30XwvDx2Oj6
68VTo3WlwAY6AtKICak9naooHl+qZmtkz4ccmQzrJVwRZJ0XwAQhXV8Ux4KoCm0K
s/U1kdMQ4D1UY8N7ULRoYUPuw8rBLWTp8cx/SFA81OROETpeXewrjMKsqkU8qN/j
nzW3wALjpw7p6YvaXBJ2oNrzehVm42IAgDFBIOP1vPEapznmJ1xyydIBkVinrDOw
Dt8dCo1g1g0KMkqd3SvaCOJxyAS8rsQK6+UVaoJpYusAC4XGlJnHyR/PUbsUmIJW
0u9akiwG5+syrlah7iEfKEHAsa6uho/eQ+pDpQ9Mbf7U8IWf13XDX3FkFmcLqFGx
M6l/SgPFHWGKCIvLf+RExoy9SEER0vGdqFLR+6wFSFhljrcOd1qdc6HWP0IfXJ3h
ECI7gRA+FD1FuLIOfs4FE85SryYXluiUWQLDVzjCOVfWiCEmNyDWC4NUVEWg0orw
O4gSpsDpL4DModXZ59amZvfqNs4DiqVJILlMqzJTa6j+xzy/2kFnnyjz3Ht6FTIb
UCsTLZxG3e/Wq3Nma6g8WgPLgKbFHqS/ORaU4ztf6YE3hq/LH4Z0Sgg7V+DJlq3S
paf3um+u5bzdWW4vGsAyYKhzOcC+BBaJlPRDWnFE7afdgvHK+bjEhFU3ouum9ItA
sYrmE4jvJfWW+K0pH/hGdmwwGvJN/d7mAc75uTsqEmqoxdMytu1IqS1IaH2Jj37K
LDjuU2p9qGDIyNdWsHko8oYP8/nVrd7MCg6owwJ7Q8hP3N64rkoE1bfMFAhZwNCt
xZ2evXT+Z2gPlQPre2Se4AJgHJgOGPBEXA2hHa6U43n0sRb4nM6aIVmHJG3RRPfT
06o0H8wwJ2hs9ToQZy2rvlwOWY90qbwU6dKlCZDd5sesGOWEbqE7LMjUOKN8cMY2
Z9WQLs5PJhob2eGS4Lh1+vg1WTndQsj4qluNnlZDuF6xaCpIYmmueZrsLvxKrzNK
tuaAZUXCTWbtZRhYvJcG3xRp1LIIq8VIg3bKtbTuJixz/aw7sdgJYjka0D6xRrGo
KrpmBca1a5Xssdj5xekqOr6XKTgqlPfF2V5gMeITuyBHIXoRWvBKhaD8RscUu7I7
tLIlHo3A510fToZXIWa7AzEr7wCiF/kgbBzQQzebLX5LqFyaHkJPe0MPiepOYtzf
uvzIQZ7KaRjULyoCy4tRMwjJCP5y0+4kzdpr+A4U+33Y9bFeu1BU1yLBQ+YetbNm
ti7rnM4ixRIWOG500eMFJK3sBTxsroNt0qZenAM6tMfTF8ayapszWqBA7GjUrbN4
FMb2bH07QFK6o6nXbMcf2ZSSS1E6k1BhgfJVulKPfnddA0UgCRzJrPlzzpefxvxb
FP+cLrxT7Vz5JfU29fRBwmUdvIqbQugxKHFTEG1rbPpN820/aqk0ZPP+TopzcRL6
VOaHhXA7dyQM55JPcbMNBOzH5L4nnBIEL4cH4YiSkNyPavzR+FI9EcfWr1Z1YAEv
q5oL4fWgQRjGwVIh5kaWRw/oScwIlCHjSdOo1Vt3ndu8pGL2dKp2B38sA38nEuqN
wrVUcWmKMfjzIIoh2S2UFabeGAP7Mjwo7D4yuXi3/dmxV+9cSTyMFl+j0MQiVX8E
6HjDCMvisSIzbn/bLxk9C4eklOWuB5hsLQmQ9F4PKooCOh5gqufNKc5QyBfeHXlM
G4TXWAYvlnMsshqGvW7+aFJvAvbiHZjdmPiM2Ttp/PhgDQdSMz61u45rwuXMQhnu
Axp2zlLn0oDXQGxBtS+YwKC6kIf7BN4Gfe1YDShunq1R9yv0PntSdTkssucE1kaG
IomhMj5gC8vLZdND5bP+lYbJx6vdlXS/ybwkhLVaIZ3GFwUkUWcjwpfNRCPy9axg
C4hCNGDZFAqlyayR8yhT6AXdNK4TVZVBDXO7W+qsCg0HKOhArHjzz/v6QuP+RYgn
RGAtlS4FnIyTTB2USN3Bn1lHrQt5qnWWrA+gd9E/fK6Glr2QgtUVEQSlP3ZlBSVw
pmRGEmM2qROJPje/dW7twpGqMgXSAO60Cf6uuIcR2UqpB60iOszX6KTTP6egRDuk
obfMQrMOH8CsnKX8GPZpFu/DwwoPgxXBB87t76L/EoPz6ZapjXsEL/GfA449XDY3
jQrgFMP7mUjYCNnCYYxzMWp30nUFC9Fbma5ra/JwvE7BgyK0Ri75m8jNiTlD8esf
JkNyJAb326UKG+hLklUakrKlg6j0guD/qFE++XBLJNAGF8hQvhojTLMb4odjSPpq
h0eltyfksQ7OoszIyQw4aZfymLY9lA2DY9AdhU2uW1yfQJGLoWYvMm0HxDQDXiOD
mSOPxN/OP4Gs029YAjsSZnjO040IrSU+X1uWITfeqmu22GS9MyFwptPxzzmxmeCp
E2PgtIjc5uP/Y0DAiSHh+ILYB5JF0nlKKzQe89WkLAn3M7ajy4+WH1Z3b0jkBmrU
AGiGFipaMBRAxCZ6/9SKqmP/2wJgDVaPTIsdFgMb1k26klHT6T+iOGe3mbJy0A2w
HNiT89oPVj8FdsPPF2fPk6YN2NeW7c5PDCk8PIcDc60TUAw1LHrizkvCwsEtDk4i
yA05vRIx4lbNZ85M9b5BKvS8zmiM9uZ9EfS8fRvmC9yPDuEuAfCfW2Rw+kifRIw3
EqinZXXsoxrLQtq3Eb+kgyfcnqx+GtJ4j0MnH+1dxEOELr1sHGguYFNpGf1iiIv5
1cxvyjRKldJ6ZD9ybRr348WEl8fIbFzEzOeHrq7ErOG5JJdtxShMOy8q6c75gXrl
4EAlLPWHHSSOlfFcNdqhkSUzqZn/NgGor1ZigwU9mn24vVkWg4qASnmFvFtJ+iW0
540yomLjqu7sKtZNAXw9EIJQjUjOtIiw0Lzrz0xvmJuDTqVc9cRB5RskUFR3pzNy
ldN0Eju0SU5bOCCeIFxJ8KrLZfvyavAkwkx1zEwbD0Wh5MqA2EU1XGdU1IXb8aLZ
Wbl/UsGmvlt0+eWX2s8zm7EYPBAeldc+N1ocC+ft8mlkrlZQrCLLnmq+JjX3mxTO
mvyE1+wJPz/aUZcgS+Xjfrhg6zsCRvJ0LC0k7L6ZmonM+jLQvQWCN99uOPk2Jx/j
ZAdXHdP+knRANmbmsfO1Kr47qmaVzqAeIUsqlnMysAtvUbF/lGUpzhedAUqswTP5
0oTEN2nZ4LH87to3nEI5KMfSsOQjJ9nIcWNB4cGlo+45bLqSzoBkpFh5RigVc0Ah
M1GEzWqldDKlTnWXTZb3uOYUDhVUx8y7XoU96yVmufskDeeSDtlsB7cYVWtPK0Wp
LzBeoMex0iRWA2mDeCURiaAkKdso4PbIw8GXKfECQRILSAwrAGizmj6hV952SpP5
KhCOYJUWUHu1KR9dWuceMvWWspL48W7avjn8iLUKwcaoY2l20FUR6yCTnMZFqlaS
u9ZNTNtWCntkle5xmWxHGj3gM4vX+P7Fce7h9MT8RMa7Ibmd5MY/OPZ2AuFLgynG
3kpOblkKHt/RN/tEYGuKmd5lkyhLgvPcjOkB6gGIIUL4q7ksbL5Mvr2k/Z054dAG
8hIyrtsj8+crNGm5zQ3CRyDoueoIbUNqVyEuuVicpc57d/spgjblrPgdkIesxIPw
k/LZen+Peil1nrmqjRfqqF5/Oce9L8G7Ew4SLbxtfPS+Bez1+F5XTNmZzjvWmVAr
NeyglH22Ta3JBbYZAlvc3TiYfB3XDc5ogO8dxlQsNK5owCYirZZPBpGNzbEKYyPz
h99lmOIm0TmyrLP/Qdld0RV8zGkbo/IDu4TR7t3V9uSvDxjGY5xBEHGVpsjbe+Af
PLWYO+CIF26qihLAAv9bOxAZH5N65VNNz2SHCpr0HoDdaUr9O1FFj2PQCKKpx+k0
SMrpO9ufLoOHlleYBlOVB3b4JHH4cqkg27tuPUlEWdlvd2IrAyKvS07JAZG6h+KA
DAGo+9ew0RNuxAoikSXH3ewIpko6UyINh0XmY72xs0wM1xUeS32DgUrJAoCSZrMe
SfvyCKQafC4AIhRMKIixRcePbCUqAdtC2jIik+1+rSpA0emRRzQgRmuxdWJX5I7j
SOH0TqB7mnsRvuJiCFk0F4T3zODJ9viKX5sZ13r6O0twBUj1k345HbPZBcWLTZAf
R9SXAuLGtbKyadtlRkn8fx0Of84iX9Mul1/ccG6lAH/Ds2NLuTGChK847N4/yws3
FBuEyN3xQ6bj0oXEkl76iBw5dipfjhxkldEUDaXLyWB2eQKan6mQet5JLC2Na2QX
t7Qm1WnFeee++TYOUdEarI1DEeT5fR/iAWqU8fbM0lMamm65v+ArMMO+fdAtfIiH
8QjmVqaCY79g4jGU7rhVNIiucvuSQ8ASfhfYm1CPFQj5M2+dYe+qutuFb914SSMY
W4lfnOuFEAAtNjHrQXbt7vMOkXZhWuJA4RWXUb22VQWWLqT6GWxT8aQ0lHYTpIn3
MBJbz1YXCgRPNqA1Sc0wianXc6Jb7sB+Az5bBLVKwVdXi7pjoyIIau/yG7VK4pLa
LcRQNMUu90J6FXuRdI8OJ9NXQja4z//NNtMj8LCQ+hSRieZeaZ5v8FaQCLS/dMkm
VlQQ8nPd7NyhIGRw7hS9amgpnKVeVUwrGKzR/WBzxTtEIshB88/Xgzo99RxZUULh
HPtD5MIop+IrWRkxfzykAxk32ZW7BoPxE4nH5dmRhUMN0tzp+783jpSsZLx8NcyI
OY6C1BP8fzp59sMaqHD763NlZ9coomXspfte9I/MpNaMQSRDxWEc+RNu5QlLY9zg
3w1c9/mYsc3rdG/buhI2F3341+qBCDhawr0t9gKII1FErsP7YwmC57vMdH+mA4wf
TlBG6sh7mAMBnmV0ctmpH8q7DTJNL7b8jAjEpZRx5zmK0JMS8IH/LfeI8V+dBrNG
VDXRH+el4NQqkMtdoDyKsvUY6hbYjIOvV8A+gBpQIuW9KBee9Lg8GHl3puNd1CfH
4vLyxWHVieRLfV6kf3lWYESFrT4ozjQTVezhXwpZfjassrHWunn/VEW2JOrVteEb
4zQnLwgDujJpw5Qlgg3TjX/yHQ6eBQMT3vBpWTEIb04vJdF59bKqDj6PyzpLQiL1
5T+SPGaYBQMtcAkYtt+Pk5l0qZwR2rCvZkM8a/gU8R6Q47JjCZYx9ywE5Xb5Y8Kv
ybz3sUCHb63smlAt9IfHp8GNagRPcaColiGwJ+kiqwXoYTtbXsDZ+gxptNl0KPZb
aj/VDspcPDMRdSknCHYtAUEYn0pL4iErMJ6ThLxhm3pw6muc5Rim7nMN/DmwpTBg
IiujhiXi/6nuwdlns6ac/3o1fX9gy7R5ptFN+TjcmqJ7B3cMb8VvR9xQVHiUHAh4
B9EWvOLq7fSpnZ00v3qp1EVn26XhIdznGx6K3bfJA+DGJOJ8wGbBedmI5AAm4dDz
SRLCHPAYN+HMETU4Jk+gCtKYRHzJqBr52UAq+bUDSAulUN7t5FFr8+vfc9Xpy3yb
VfwccJRq+U2jZ2Z1fu3bmbutnEAoYJjbiGHz5nUX86Rj2iWIymNRNsHFSO/Pl3G+
iU4YWdgp75Ijy82FsECOWZ8AVT5hcxpFbb0ifdFbaV8BxWU3RrrLZUmqFH6ECA0u
A+hGJLnK9vrU41qLfQxERylIbNLFMVQnLjioiJMfGjgv1gruYWKxgfQyUCIv4IS8
lAGNTafqJbyn9byv85Ax8GqWP9fDOD/0G0pZG4zE5wT47Io/hV6LrED/470o12Jd
y7o9G3u3CATNtTy9UARjjKvx8qWAfua89fiF4EZa/cqJmZ2We9nLMhQd1VOtHLf0
t44jKl+loWJqVMKeY0RzSFuz5MXbtmueFfn1ZHnLX6Icozfo6rWWgnHFCy/Gf+CF
BBugVUKQRQIABCqNlhveR1rrEde2AuvoKUAD6Y0gn5cU0xkwmtPq4HL17LkU0cte
p6AbaAKptedC4XgR+JEGF4wCJzl0/Gjik2pQFKm9NVzGmbs7LXDXWx66VnAmxJWR
kTQvqwf85fg9C37ld0p4jAVyyvv/1QO+wgCPjHNW/7iY/OSQHEbJMrt27DbUFiDb
iKFppqY7gPHFeB/qcvsdsEqab1eelqszWbJ/DpOcp02eUXYGmdhhCt+jI8WGD0qv
U3B3q03cAVk5bnGoC7WhUF+QVSf1BsX/k2a6rwecnRQoK6BNYZRJ2NlUU2iJkk70
zs1isEgWfhM0miql+AVlw7GrYax1l/Qj7KNJyoxaFjn9+Gh9BLt3s8zCUpwYpu02
lNlDwULMLPZ/nCaASXiBWmANcOlLQ2Ue6xufe1dcJKLFd1vkCg8730mByvExoBzU
wC+dE1n8U0TnyPsQB9kGL+YrUwq8Lkcwd7aN/HdJTcmGqNAakqsN1WUUmBmuZYG6
InCf1DdgRSY1oex7XHiKghAlULBhTjYNJxuEp19DgB90db0QiuYLKN6hZYsUFRo+
hP9niCkl/KM3ZNZVQ+utXCmYbCXLgXwuyDKttQ9lb/Mbl5qhpDONbvdaVRXoRNYC
bg20MkB885qUZEtOFAIHCagfcEBt5VdvBYmckIi/B9X8v9xNAg0aR/xOR02hNb0m
BR2827mM0UWErGuLK6Vw7caaWvZqzbrqywkmh7U78RVNs0LEy0H5e4DTzuM0QCV2
fLTPSCEUcRlq1la4AqKePlc94NUUDEHyXxVuKqhWjC9qxQ9/5pPLjpT6vZ55XOpf
X4XqziFQ0q6usADyuYSYuE64XZHBvT6zlfyaCTB+Dyqgmck2VF4rRgRn4H4qGlig
DjOnOthBpNoXod/lnqQ7ZsUCx3S6dDGxvVboZwQ77ATDl/HxxtMw94/6ysmmEC0p
o3Qs2JamVn6SzRO2rW0lYjRFSlZYE/uyOX8asunneMNXGvs5t1/LaRSLd14FuQQZ
ygL33gKDk7ySu/xQq7tdIVL0p0ltBndIALuLw/z943jQOeynEcNbjZehVdvDQChe
YmwJV5HCmKIgXXp8CPeInwWbfswxkgry/XZDlR/nabyxbqLu3s7+zFekXW83Rz8/
me4ysYiHjCgR0hFFaZpDFRR7hJUAXG3Ap18vIvhEnjPM7GwxVwuHwt8s61HcFGkN
REimztsSuE5+WFgUXHb2Pk1/xhIdC+93NyqFOS6gwhRi5lfGqFaJOdzsfWAotYL2
Vg0aHssesl0ww6QhXafJ/69xNO9sKZYLTPc0plrRRGk9muNvGqd/9FvFhb6satYH
qSLqD6GetuoaAd4+g0OhErLqm4vVEI8Vun7AWhyR/heMsN3vrmTM6/RTeLgfKGnH
JnJNXwlBVEtLvW8OlEDQQ0A/a3AcBHSzPDZnzL5Ecs99uuBE+c2/8qJj81+p13nP
dgp93+jGp5iYl3/car6q1GGrKuP/wQ0wdyibFqLuEVH/lk3SBbFMCyorb0F3hqwU
A9hivFgL5SchNh0/p2h6l90+4tOyFb0Ha/hIYzMMGR26KtwXqjFcGqWMqP9J7cdL
XljHI1LEkVMose5V/cKKLFSUg3+XEKn+90uwEIB0LjA4n2dX1vZOMo4RBND6F4hD
Qc6P8U2U+GY6NlgvRCBuyQn2NiO35+CMowh01vlai3V10LdbJYVYJCY+OP+kLMzI
SMvTKGwAPQ25y0EngChG1fB2ynJwKfIPkfHivcJDEZGhyExXY9W9vKOxX1MEHYD/
fi1TE7QZZIXk3QtrnjbOZLtj4OjW/KTcrH1mfcWhoCxR9P2Xcpt/BemtzJ3N7sWL
P/IxOsWJ9UkKsOyKep2GuvlOE82wFxrhs35/pvDJfS2GWlNvlEbcnOjHPKwwc3Nb
I4ZsFhKcTL/Nk7nopxW40fPQQw65dN43YnJR3HFROcMpBIk7/JBvVQ74EgRwFBb5
kYRfoRxpAlk+jJcJIYujVEDj8WJsZ2s5l1y1lhP+NUZe3/3GzlKbyeq/u58z8HkK
W9crJjJ5S3qT4TCya89LRBDQUsbkXH/iT5TU9Vs7dCPJ82cyAg/JtTlFerjjFThv
94jx3xeW6uPE2S1k/mS578eGwVbFf6l8ofpLUj5RbcvtNxE902KBTBiWPfDAtzHV
/AurgtRQVa+FA77z4cQz29tv5hnmS5UDt8QcnqrjYj0QXHwp4gKw2o5nmV9eKrOL
t/kQzFnf9eP5g5cJCXmRlPs9ztvNrvSvoQo9Ud9dWwrszMs/hq2MSjOakfy+aNZ/
2Ueoyw7QQkFCyRvJHinwZPSsb7M5ZfxHzt34YfrFDnIKe7ENBYM1+g3JHBcXojwL
eNU4xr6OrVA1w3jAGRwDr0gMLHUhuB5X9gbz1QL1O4vXA08uR5PSsVOX2yg1mhS3
/djR4BialANS7ei0qjDVzQ0TI3vkj6tbdjwWcbMdcLjKddFc1CXVDQyjDdLV034p
kaQW7fpFKEQCYrewSH0jkVMS7yFbCCit/cIeAWBe7OxdQh+2nXUJJ2NprmEsjKzz
E6hiGnZffCzoYBVI3Bkqz7vXt41WOgXsTJJqjWzRtUkm6eaA/+jv2imL0fp9tD+J
UjELa2VwGdIYCCq6msKCVkOmc9TbWhkaQZJJAMIFh8ElYff8xCKE9UYhgfU7C7ss
lTS/KC7bASUL7lwmB5HvkMDUePOuhjfeK0OzBdoKOIUvuMYkJ71dEsB8FgQt2esg
1l9A+Eiut0yYH2/R3fW3P7iJ0qBdvsFEbHycLKDtd1ml0XpE4qn0/sR/UqXPpKiP
BAoAsKQ3GSuMEibMJEEIz4JIq7V9dq/IbJiTVuD+0zq3uneGaQp3xc3JEsrJM8gv
qAZcCkp5vcJHZPh4AeDela8A8XqjwB3lDOKikZ6K1ETymHZW4VHRleaea1QrVhNN
YDW8ve+dJQHBjoHiHrzYIO6sLt6+emtE6RKuN5fLxcc/r2duydzCz+cpCzjPBKOm
UUCjgwAVSWJ+UEyIq4aRv2GX+RCus9GPz/2UAtMEWXRMKQrYn8K/Ds1P3f5qKYL/
kABmUJhM2U4nb33JOPAajuAA0I4OlpHmfqQlvcy3QmxdHWnxPJUrWMfLq0OB6tOW
D94m4QsGn0lR6xMFI2X6VRBnmI0t1oddYlZ4aZ6cWczQvttGBT7RmZ4flVOhZdyN
OVl+uIEtH7G29eA9NjAEx7Qk2kwPikfX+Q2qtyUGHsLsIGiRFPugzxjuwQL4HFs7
kdrmI/NSDYOBfWGp9un0wR6jJTy9P+6UdK4BrJo57psb2K3wb6M3bz2skEsNSx6f
7x+ykDMC7x/EsvSCTy8tRPRwcxonxNaA5erzNv3/Zv59UczxzQFaOnsY/+174EiL
NpaHnQEF0oLcdkaHGORL+zI4j1ZiwKz7MgX/cRZMSj01h4ioDGnsVU8gc+X7qQuB
2/p/GcV06ZNv44yOi0m9Fxw8gE46Q+RNU5BfXUSircLTaAl2Kvz+I93huhbu/V11
tlB8HBb40EsPQ0qJNBjtpF54a+Eum3zjydTDO2j+Eb99uaezdLY3g7FHlw/SJrtO
zQPkU3P2EM1L5TyZi63UZWW3RrywVQkYtwY4Dkbk6RRW0WeCTRA5jycQA9os9Dw9
yNMYJnz6N5qR+EiLmGPFjyVjzEfAI8kuurbcfvEusbq0eYz99v/Ums+CZe8fTQjf
MXcAMQMtGCYzUjXoPiV34sdBsObQnHemFccMmASb47/9abeZekM1UZP8vcLldRhU
g8zvK/GxUnkBWbszd1lInok++/DM/WtPBnWtelVeqv6klR7EBJhRScA8hEEJa00y
LLMAiQyFm5A/gvfQ5yEcBV+p0PZNDzWpQjIHkvj/UebUbwAsksvFC76NM6/qocpz
mYEW0c8qTGswc0i65QAcUdnrzO4aUjfIaZZDqm8uzHXtbF0sInYd03UIA02FXTI4
R0gEH7FnZwdXUStnQQOF3llZkpIdUEUvHJFUXusEdtv0Vx59Qan6KX6tcAyMBQJA
+Je86kWFKQJxfPPoVQq8iWQzYdygLAW7hd9Xmij8+zgBSICGh2RyNKg03Uu+9arn
6cuooBI4H0J0IBaPoe///0WB3MQ5Dk86xKOcyOdfGcPIUtnmBYpC2nLPo2ZFJv1t
w0vHZwnK5RUUTCDyMnDU+O1FauXJTYQpgyvzktNewQs197mwwC+mCW95ZtwE5DTZ
vHlyRi1BHqtfdME2T46jRX7htH3gm/TAL2851VmZgLy7WkdKRF1vyZwMMBLZK0XY
eo1QSiBHl5/JsdRi3BnpgfPm9ZFdUsI5svmouJ8wLuu5nrt1b1mk1i0fm3FXCnNm
jiQhIusOiusLghLeELG+qgXF6saRhY1T2lv82Q1aQLk/pAlnNhnPoGuizehwJr5C
J34p2k5DExdx99TVONYxM1CiuiIvwfoxD4kJVq25phoWVJG0Zqoab1YLkLvhPY9+
s5SINzcPbdl1dsZQuKnr+D07skSuPwLHcQkfrgJkd4AGN3VoVoGrln3slKDru/3E
VRqCPi13gN1yh0DgakBp2EbG8kAOoZX70v9SH5kZL3N558F4dOpxZmLa75wTyzKy
ANUlIA2uAEjSeHyQ1RX0+pm5V36fCtJZnD5IylmyZ4rVZyPzkDzpZq0+qQyQfXyT
OxHHKVMQq+x04Ztxpknz4t6O+pRr5F4ip7i9QmPj2Ywsx7FhU8+7ffOakkKH3MWS
q+xnzJr3VjB9Bdv8NgWZPnDWZUJn11J+G1Mlfy1bJqZ9Cw9WrkdjTwfKJcXvL1dg
yEJXGxlXK9UQSFJj+RozyZeP6/QC2gUMsnAIqwqAZ4TrbOQxlMJC6n7GA2mZOHsf
VuPFslphVKbJt976QXpg4phru4AZaFx69oir8yIiBv3dY6220Wzn6Ay0ws3T8yoR
t1nfgCKxy/oKWoBCRnlS7T9cxTMAPy8lieS3AoYoGi+wvFzCIKTZKDFObRk45+cR
sVcRV9oQ5BblDcKhCm0GYwKKWM+kVahhRMLyRN3YME/Nj8Oxz/PrKeO9u5L3rB3v
QwB7AHxOj9G2M8bJGWnspoG9uU6AZvgg7DdcZgzBxWlSnsS33xjAsD6D5EqjYfpR
Xc1Ik4vniT/izocdXH2CoNGISLKlIfqfbkySdjSwFIUhUhSKaIXnsu1z0YFJFnj8
dCOP5KA7p6Oj0GNm8osOk+X7gGaW09rxLpsTfKPrq1E=
`protect end_protected