`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6288 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
rODdjZZu2GxcKE+Z2A8Tbp9q3NcZgpi8avl3zyYPch+eG2Oy3riISwpVBmm9ckUc
TZpDv8vx9DtEYkteYAsRzb5qaoxV4rimIj1I2oh4pXt5r+bQfXS27CRxAOmOP2yB
4uBIB7dhwM9BOT5gOJsWABWiBu3KSE5013+P9E13D+5FsMGkS4LSfStNfIQegQa5
4v+JqSguQsvrcVWJJIDCQtyOlCkGKnEVEBlmueZ9x6/gmjBtwbliRZr1d8l2ZkmN
rbAgZW40/cVbuaWkH1S8tqmqtr91XU5BbrqyNNlE8CSDfnFWimZ05JeSNSHsq0dT
kK3vEXm828vl2SQdpeC3sFl6nnRiWPZFFcSCqfYGhnJT4dyh4GUEzzj6CV3E7d3K
x09i3muZTIJmSQb37u/k9bRjhwj2PiT/0xYKBuuYOoc9C7D5UiI/35blFdxMPAZ5
wuZ75GZ8Nw4Nr9kwAm8J2Oz4S0bYDSSxL06MFMVnOXkCAmqgJTS9RE42fgf3SJfp
hZnRWeQNOG/wIi130Ob/lrESsN4ffSh+aa+Xj8k22d+R65zrkqkGh4xL9UZgSnQI
933QZnoEHXXQMOVE1eI0yCJdoFvFpeK0j42CdL2GP4nI/5LbRHdLx0bB8AE9fnIM
89lp0mkuWvR4ZzyQfyVpqdgRLdLqkRHaw2rK7CjfE9/RkHFbl5zTdED1kdzI31Vf
sC0T6tYPGCJ613mkZcGx+tKU7gnxsSW3XpvSRrBWTJrW6wofBSQQ8gVeaDUVDKPs
ZA7r5jUZhEANgvq3ISwbK0NmejBscnRcwpJI5tnvYlRZSGGhHP8DH7cj3zz4MDnj
JzcB0SZnYJUXd3teBJEUfVzKGIFK/p7LvnjojiAcrwn0S+qwrs7FjBesFlR7ATqv
yr0Fmx3iMQe/fXv2lmgWO3fA4fDWLdYM0FLbRRkhP3dfIslSN5irUi9SdS1lvCpc
eLhliDs5HDxhaHrHO6sTJ09HINvAsEjYCKX5HGg/5fZ3Jd8FnMa7ws0WK8HeKrMt
7rfloEbNWMMiqsyiEoXAVS9cBw/lcMY/XOKst80pVXb7IECBqxA+SEtF6l/QCPk7
7qzGYpuXphcf74+L/+uqw49CYt6n0VeqxqVgNphE6fTn+BbQGnuQB5lhpMD4gn4X
xRxyRv67kn3rD7etQayhmwDgJzz9llKkn2I8wWy3iDvPE9IA3UPn7SBy0Lkot/Ji
bHXfpHLQP+z6qYt+DmQrfEky0xo02bdES3eXHIbdgctTewUx08MxlxYv/TilUJ44
C0UW+o4ZJa+P9O27bPoP5lgHZKce7MrUiych2E/EK2P3klX1JJyW21raSD1HxxSn
jRw8+yEvYVaXJrIb2TIqI/Z9/iMEyZwmeOETHhPfV+imC2PFHDcpS5jBW/oS+M39
4UayfE2ainreRKK2E/2fyG5UEn8cgjqaSZrO8St/QioSePtAx320HaXjGHxRNoOo
XuLDAIedYBUE2WIsRPGH3lbTsF8IYI5mk4+oaiw/53rzYtQBkUEchqw7TMz61EbF
J0P68fzblYIPL393tXGNc5n4ylH4CI5a9ClcBGsmu3UPBXr+wec8+BS55on+8SP9
MMcFWhyUgFTFr90/O+3CDW4fDzqpoAhXeB3rs9Ws5+u6B5ihWghOorojk67KFBye
AKkMMFgQVJ5VSfv0oaGY3l0u7LNaHdl1zST9WbqjOf54yC+CQ135AfFTANP3ZU2M
FqC1Ojwwy9iy5umLk+VE1RIKJoSRLLjDEXQmblbrFJh4eTThrEG584Hz7R4A9TH/
ylarcytC6VRatCQ6zfZrjyPRMlF3nQGh9n0IFET/NePeSfmk4KPepRCyJDg9Sgwb
LHz3kE7R4dcMC6BY2aL2oz5n2NxZZ8gaegjY/K1WkOY4GcV7hK24EMkfxBL1k+KM
VfmXAb1dS3afjKPsh9afcUa9ukbd4Ek7auSqj8l1duQjwafvQrUIpgwUDG7FAxx0
fiZgTXyW4WS42PWfZ0gpz/QCGVStQt+3XXIzuazpTNh0l423VvIvIm2JQ6i534O/
d135e0du2En1naMoV3fG/gjYVG/oq3OKspVVSk0NtLF//AlR6rpAsVLDokjnIrW5
5M3zcGh7Ir4MPj8X2Ago4EQouQ8W0t7stMyBzpq47l43KZrK0MNxYrm/ZgLHBmWl
BT5IuRm8k34XouEh4ojGPW6CipgSRnFr/aF6GqeGbZcmWNkjxQqatr2Fdw/n2iBB
mirQSMEB8Z2b7CRtYdJYJC25IB5cKV5od+/KrxKeTqK+QlV5+4RtFs+dFtS0ZRUv
5YD8Xz/IQtQpEtYgqiP8O2moQvgmeEBieLIVc2zRMpRaZdx0b7XaHeharXCQWVFM
33GuH9E1qDWp+Sbf4rXnt1iqT1elCGW4oyQrVIZEgK5cw8plrPUdoTXfF4kJlavo
TuLpYjWcqPQZ75qATZlTj32gD3sqt2vZTYGQfheEhoyxO/5TDNk2forE6C5Einqp
WDQxFg/dGaL+q1AJUYZlGfknpNzxNG3diY/dHwEtinkMGmwUxJ4UZsci5I+FwHsw
lQpbPFi44Vq/z7hAxWztg934RVUSEC3M0tXM2UKthJg0lX6uEP6b7JAAuXlLdOyd
3qjsyJfmeYv1BT6MgKF45v8IMiz36g9XOg1i1cyDvAChl8XTouPR5NIJHRGflVro
0nMPxH8kUB80TkpS29gPKJyBDOdwj4tavUI6DBOLe543sGlOsHS03ST5hMr96/yJ
i1uI8DJdq+9W53rSRxJ16k8T+QLu338+vKLeCPpq7XWkZR+mT7Kq9cRLcTVuc3AD
CRNBqOmq9INM+i3mGgTslXKFiAqPHRVzJNhXed7fjGUMek7r5U33DmWHQWb3OWPo
u1oCGt7VcUyMpnnOyevut47I9MIh/U8dz5daBKkVecMVpwjwkwIAbsGdjL3ux4V2
w1OWDa7MwBa+CeaFIGU6yyIxjONj6KztxxmgTjKMca1DQKXaj0nC3OiOBeZwFci2
IaisnyFsx5nhzYrxb/NhzRjxW9jJyfmkgxB9Yl9uMoG59EJsEuHztILrSJoJ4occ
isjlYwp1w+x5foTxK3rReB2zlapz25MeE4uaHYR54+XSfGnE4MYY1H0J95DhFxqh
ScMJXT2L/w4pkPSoz0Qu8e6xLGFbKNNbpdXpnPRXaUTCsxn82JNW48HVchO8FS7t
gXXqHK2zKRuPQko2/oaS4RuUI4kgqWoU1k4fSQ05nhY5eIRQ6EVCSdPQgz8AKLna
+Ths63v1onmg0ThkjaLzqN5yri2d7NPFFquqMDXJmIGGvx176T+w3DdfI7Zxbxgz
b8+GjZx1BdwSX8cnX9UdEzNXXCWAdBOLYlmx4K2AVfaMXe7xNKrbos3XsQT/5wyu
/POU4DOLWFJx4bKKyEVDIl3lUp6fGG3h9uiSq18MBovjniPgZ2rFgNgQmCIJMS+z
l9umyXs9IymNkfkIThFD7H99iMAPWAzrmHm1FQAsSJZIAHwY/00lkuI0dg6FOh7K
a/RdNsp8S4gxJ66MRBmsuJiM1Yu7BXbGaRhVpAQ7RQB7AOnGUiDUHj8L6I4rZoWq
Xq4RKVZiXn48DCHOvzIaoqcw/VKPKHYDNwxDuaJEwjRUiafrAO+OVzEDZix/K2qE
9KC0gbNNiWwbHwRKwq4viQaSDrFdSklBaKrHu7xS23xPi0+VJi2aGomb6FS4HcEM
xt+/FaP23aGKntpdMxr7qsqoPoVjLCg+YYslxg6hsdSfNlviOmzmhp4AmQ7AxkNc
guyZ/1iG+9ZtG+IHyzpu55RtQUpTA2Q+PsNpQe+rxAROrFC7pV2x+2fDLVr7qy0l
T7+yFXmRd5ZuyqQzlMp+LokOEoCrfDywIG8dAoj3DR4CqC/DF9xY6ZGtF3YxDCA7
RN5zj6iTwTjE+0gSZlGPCnEboglV26b9Ku190TWQIhSSyWHoQ2Hntfix1M83D3KV
zEWF+YGeyri9/yEHsKjD5kwtYa4UG3hr/HI7P3r0nzHe7twAOfWCplXQm0rXTuXI
WQVz3jjW73IlW54UNPKGRehHrqAuz7OznORNUvt8y8E3Ha9A9txQCLrHZO7C26er
CNIpFNaECGLZTcbiXKYlAoGBWpbAcL9ooAZQ5aJv7X0ahHuCZEs+AD5pzu5Godha
OUr+83QQxwSCJfAv+ZXLmq1Lz4Je1nmS+2ZQzszTD8ktcfp/yqaiB8mnilsmjfXl
/iU2ks98wvo1Wr3U6SShuvOpSDZETr7S89EzFVvkaZwbnUrZOvRU9yxWLBzaZwDo
1SN2Ck2AL+S7oXq9bvSZfNd507HYGDVp5vXqyowJv6zTd9PXwOjE7ZoLfhlrwtup
JPkkwqaipmERZuva35lS/RvMZMyuTgyXyqshErWaZGpZ+/wfb7hCRlSHn1a+rKTq
KcYeq8/2ABQGZqpavMgks/7p8WUgMvz9Z/dBV9RlyVKo3uA9kcvrOgHwdfKr2V97
M8/gfn08HhTAsmL4ANU+yb5B2VHURbu/aQu1HtVCIj0M6XLqOCPKekwDuTezH1M7
4P7qjfHp3G0ENXs6TcpV81+Me+TorTLM4SmVWmMGb1Fo2abBvIkqB9jDkCIho5p2
bszdsIbHazNK6juzVlzfwYDg+Dhbiy9UqjAnHfmcKtigOWJc2nPwzwmqzPsJEW1r
yZl1NxUx3EOmkAf+Qo6d+5hPUArP4Q6by6EYdc9lB5MvswNoUkszhPURYedh68Ra
g9iTo+IdhHoFhZbgVvYVwRrtpGKP+KNlNSy0OrGD3cv+YCHNGfTbDkWrqR/JtrXE
8Jo0Plp7GX3qA5gbLahXnlU1T9tHLnL8qn8xU5qs/YIrQWxuuLlKbEA4vL4StqmM
oBRfHjEoHs+dmJxeD8Wm+RYB3i91ixFDUfWtUZru9eV3QRe+BCr4PFuplZcuYSjt
dbi6sJLpInr5DB/SqRrHnSRp5GWsUD1gAHlpEzd5sH5nkAvW0pTBaQtATE+XJom7
1U7iBBBtd7fX8sF+GecyfSwGD4zB0urmApMRkUT9SzxlkeLz0tm6veaqeOwg/uXC
iW/SU+VIli0BA0oE4EE4MV84QSY/XvQNBEqlAngFWNM28iLt7j+hSapbe8MSqsl+
VMcsQ1BW6j0w3owf/R8u+xGQbksPKcahxjx+dtg4JlHloRXIPtAj+WZBu5AjpYa9
9mYsOFxm+XSfuuMEjM9ECy0O3uCcbtuyn2KtIAwIH3a7fB24BfudxhZhHcihuuhC
NAD/HTfPlmhJtN2evWvgrAgrRtGIPV2kue++rmnnILzCG3W/1T2fs3SZ1mVkLwq8
1wgC3DWMHf7G5YpA2ypB8+dr2xNNR/C7TPinaP9y83FeiJn1pyyjUu66l25mAXCq
fEJh9TFWE3e0BwhBaiYP+md8Z1BFmO8m14hNwBvYPTpj9Yg/8c8iNriDvFDXPreg
Ah4+jG+Etuuqottvr6eSbmx9jolGMjTXDEfqPcMjaBkThyqoQW+iM5+VbAnj2WQZ
VG/7SBEKOJ0rX0KFjGaDVE6PA4jBE6qdprGjn5EmfoupuWg8P/Ah5kV+MtsVlQtW
jBsL2pJCWVEwyCOiYtQf2+m4KdtHnhNDi88/lF1CCkFVjer2b8phBvjyp4897ciO
TiLJ/nsqosLd+cLuWFmvkjeBdHXQRbXyGZwt+om1oLQMztGjlHHgp5fse4qCFdim
n9UinfTffq0iTgABGkpF5+KEP3xgYxdcof7iWYQr5Um2vTPvz47FbC9s0BxQcOIV
V89DA5f3mn/IEgdUoshmpTg2WQ+ETt6V2HWrGGEKyId6mA1tdhBuGSvXGeNLxRvn
q1nEcwMmpyuhRSHwhbH4689g1JI7D27pKH6X3p6DFBO7Pzn0UMBIX8XoAI9Qt6ec
Szk1iMupWFT/5fRqTi8EVlft0BkuTXY6EyHwFpuPSX6qwoNL+dXj2vN1hu36WYp7
gBChnxewKIoGus+9yZ6pMW/vpU8/vEe6KJ+XIRAL0aKGfYp8z5XkuhhjiSlY9QsU
Bew/i9wFCjtjZ2CDhjvAomBwrC8eFxB9lQ9PiCrXP+uT+8wKUIGhEnG8kCWV8+WH
5UB4SMO8HHXCqIAV9746Lycxb5Yaz4xtFiknseaCv2LJL8RZu8ePMN/gzy5hg3/y
W/HnmwRvshiBmByU+ItqOOJiXBLOTnMnS1swan+pYFz6y8wJJNeo17QZbhI9dofO
iPYOHyuZ0twquz78tsf5M3GBcj2IQs0FFMb82iuPwYwDIBCP3wtAVmgjAtKNd+nr
ToLl+NohKedBE1YkD6ZsAadGJHbMNPxM/6/8ZXypW+9khPua87tAu54MjsLSwrVU
BXOEOUa/8vb6IHi7rO3epSE1LyTYc/GyRlrAyVi+jH1TkWMBIdXL6OfD8xkCghHf
O4xttj30LVCbXnfT2KvTl095JXqwEaT9RdfQNv8+gF0NieU8szs8JO8SsHySS7P5
PiHPDzdAqWrlTc1nPm5b/5yYy1OeHuNLhYwN4l1g39/sUOMp6djHESRsbduI5ZKU
CKkwJpUnBF1Qcw9UJYj6vlvmBmGYuQCUbDtLmzHYGx8xhkG3wLFpUXLEt4fDEvb2
BSmjsOIXJQpiLzPEpT4jRpQ8WfnbWvrSvlLC+oy53mxgmFR4kdcWgmIhi5AiMsDc
SZJ4fQhDzAVFtg3VeGxfMqZCvGhAkbiKhgO/6SduCfuQFGi5wg01iEPpHEFBL0R+
8wGF4czDTT+LIZ1upYUEcvWdM/cALNido7Oef2ib7T+4Kt9oEzNDWBNZOdICEEZw
YvUKuVNITqib3+vLNNaR2SwxzYLyc+Sx24jy6IMUZosKGWUHBDl1zpMNOoZ7lNwy
zUc+ylJjU5yIdK/QqZM/SmOJFr/QyBjyRAHaALrM3FTZ13AFWv0SW/f1+8WrnOI5
jzoH5U7E3t/hvOUeyunEO42sXUA2qDKjx6fad5P93XcTss8Vetp5d0OS3PUQyjNO
XfCp12YGdHJl9Wjki1zLZ9waG+NZd8HWVwdKC2dFB14LidxO64UjOzZ+ic++q5qX
nCJmLIoWMG4j3ubM/iJ0VxuUdZrUu564q2rAyeKT1L3d/ipC79n4XCdTqP3mRnz8
oC7rSRP38a+wNHfIQXFh9+1AMPUcwPMCQ7TZbJMs+JuWn4S1RaT3kVXKgs3/LkdP
eaWy9gZQ5TRL5cge4jh/rwFokLd60QnCw1+H1U+9HeC7Ix7LFdD+R5IeJrcNazoL
K63wh9HeiaEMCRMqJEhqQS0ELHkUBdFOFzCpLfaflNuBhj6fVupIn9PeLOm8B8xm
bxYaeF/z2dPLdkUiou9HuUA/wsTkvSkhgn/i3LYhFI7A4BE1XHMLA4a++WDIjIxm
F2L4iPp6Zn7j/m8lNg1hU+d5MTJamHGHgTolZ7dCN4WLEgfHcDP3/hu0GwgxTJFJ
a+VbHlRtaKEWjEnHWBKMedwQKEALHQd1vCKwsVJO799kQASZtpWr3jMKh0OZgHbt
+YQiEiuDVZeO8/f2TJOz3sq+rRXLTZesQVIZL6bNYPF0YUKCzl7hpFkET/BiIvyc
hmDH2qG31TtEX4Xk4Dq471n76Uf1694D62dqpzxgM3La6HH6yh9TKNCQPGJGSf+v
nknJnvYpgK4x4ZXHy2TTZKTVQtXnoyOUWDLTXMUPX9t1Yh02qexnPuCqYdTM2q1v
56MoHDmIa5FAqIM+syAiz4V4V77lRkRwhoYyMhlwZ8gF0S+IpzZLIucIznkAmqDt
v8cPNPrJTaSzoXERJ/ZrVwjNLPTw4IemzDL7/G9uWNsS+S5R+fYolyoqqmv6pczL
8jd6YN1k7sq3iIfKM12aof6trIYHhA9zVkOhRoeqClt9t8r9mlA31kVDPLASBHHz
jk6xAkugW/SA/k/6qyslqIVLQFfv0QNvs0wfJTw/oniNLvcqlNnb1pEEJzPIEWK/
Skg6RGLQdyNs3ikQirYddl64FS2/izh3UO5w1WP5rfZlxavR0Ds4S6BPFPJ0iqV3
dlieuPysAoIpkEfpJG6TBLfkgiGMpA3nuxoIIWIxO5M7biBsjpqeQEQuoWGl8WUE
uIvBemY6jiX3QBOPlN9GLJ0H0hzYdug5Y3XPqitZOBycVGO3h6dUrCxunpi1OUgn
XTUFM6Z5wwpes9mwvQ6sTnIOIhdAEAKhvMzeKiSDu0BSrM4uF2XkYFwNjkatQJgY
msnlKOfpjIpmLo1CSk989MQwggTTlodhruwpx4vZIznPHnjE3oxq7eHAsbr/umm7
`protect end_protected