`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 27696 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmWdo24EC1SLhDeUV9o12ewQ
ulXp2xSZ5P2RSggIKJUy/VAcWxVhQIj+Pc1Xl19u1zbOYUXDBYKKdO9WJgKoBALW
crqSVpHh95nCQHnMZsbfwq4MqPKbDR6GawQqz6sA/lAttsQRxFBZ0xdb3gYpVkIf
WZHQPFsaJ5FI7Rlgxwv3wjqM94cRIVum3zFQWsEJQpYmGrJLokTeNMW9e7BChUTt
s+10oqALWYtrk9wApkQ5rVdkvYEY/DXLIGZc1tr1iicKTc1/tZ1tzH1+DF5WzU2v
ugjoh1Br9nhlHYZMstE08IXnaNQJuBPxUYDfLFn9nPgbnpsUMcEAeUfiwQjrCuKG
SU/S6WcHT7fJ41c6YkwfQIUUvZm2EMhCVbvjIMQinsv7YpPYYoFt9C5yXx6WQNDP
qyvIG4anZbFGCv4r6g9eWMsG1yNRyF8FMvgUIoe1hBgllvIByLp3lcoS5+07zpkj
+68UWNDTQ5gGNat5RJ6baoKgczlDOrQLp8aS/1lRIWLEozJ9pX8uwMqCVjw7ICZJ
gt/2aLe3OkPPV3ZAfst+nQgX3gi6jKw6Z5Y4CTBEzfbI3fPWmXlt3Zghfg67xmH5
UNR4qsQH1NgEgNWqPOM+/bwtKNS0TKVEfWbuVX9CyzqDOmKVqL+CZ6WL1goxwIb/
KyPnWiLxDM3mUrmoHHr2VBl3ax4vIH0QXu3skZRwcuH9iCM5M1Ak0w+g4oEiWFGU
/hly6pPQPuTg7Rg0YVhmW8jSJsaoMd71FxtXui/49X47WfMQ7BBfBJFbGVA0sAO/
hqs/73iJW6d/zpw4S6Kp69JSbSZ4BssqC3pyUIfGF11+Nz7TAecM0oJtSaWtzA8k
QNhtaQcuVuEJVNTChvsVgMSDfRDo+M6Gfela1HMscJKLVuR8yC4anAPJayC42Y60
xntDVpzn9vhsysm8fPCrt6zFnUT1Aw0HEAN8bl1Dua9SkLm2+nrNpMEwfyxFSRWI
O3Ytf/Wbj/B6ICNd0a5k8ZqJzZ90TrC1MVZiEPDZvqyq63JDTRxk++hcvN/5779f
qdEmS/zA9lRKNs7xzQHdfF65XFcJ9IvZXII4TZR5H7OzSidPs1yF6ehHGafJ9iIE
hG92dsx6ZqBwu6wxpjGzoxaVjtgQL4jYI45jEfkaZUtWqSDRWvel9MH2rrt7H+mM
qAUgys7bdI5+QzHlGBaVKXTuxddHL/bM4ic/Rv4q9LDtbwYEsuqNQqIpJOrojtPC
lXQB1m4e6ODM6kWQ5eWXRuENWOCJwQuaR8ZeIQCStcn8vtBY9u3BOHUsr9xraTGF
42OwzLTbnPYzJElp5/YXeb7QEFhDx2MeuyOuIPXK0jVX79c0hh0i8018JOtWU66L
TfRnfKiJwGXFG4q9vWy27aPOZIHzBwgLdNnu0BN1mHV3rJ/V1eZhxdQbApP9OFKG
ax2s7ldH87o4Pjh9HKCAy8mm4ZbXK+O9ZxjLpHTW0g/D1d2jSkjB9Dy/SlmKjRxe
1mekSI+TGiiNXP3OpmOWZrGPx+D7ci8yCbEsFiK2kTGEh631g4GH3SRXb3uAj32M
apG7RjaYCPBGEwe5935kX7EwtAVkm633mLv7lEUwyAZ+zSGhCCDx9W+6wSz+FOv1
2YkbsDsGk1DV/0dv1wvEXEEsvQ6ravo90IGgRleiLTyCfSUEYhsOi8btYTijj/rS
5oBnMVaahmqqy5zx1qnKDDHgFcCGx96tlRgwDaz0MPpwkE0pbw5Jk1+mUnFX6RhD
XgutL5n7ATtixz+0BeXCD/AjsxZE9HJzLybJqaI51XpPm9MxBtFR+nuDTCU1/xpn
SfaAA3D/p3g5azGkaV+FQYuEWsKpyh5a4byx1lUiE2x09Iuoh+zqiLGJ+z6VtIPC
L5SI1X6jhdKX0F+CBxm2l4H/fucRG669iiT/uDUYrJQbokcP6HiapfFhGUnL3765
eM1e7jZHNXtlmlzLqZNM7C5mh0J4HuuWQZbxvDYuBE45ZZKbqMQv5tcRwOsBoiIn
Lv/XDAzbqfAZvfqqfjMOYadI77RgjChjM+b/c7MPsWO+lHx1Q1wGERyM8R7hmCzh
JyXMQPtUctp7WRPVjSFvdOIXVFSBzMrnrReVvIZWvISufXrgMCrVrEAJEYJvPlkw
6heCk3K8lB7viGqeMMMDOuZzjGhiypViCh4VXFAFr4qlXCS54HAntPuzaZCFFJQF
75skgT8j3VO/RDvLpAEDwDnQJd9as691qMn5EcXx4BCeljD052XNY0/XG5Y2s/hH
W+06Z+GQ0/8PEQEO9AOnfyDFQxjliODnQdLu7UjoCZuoXDZVmdWAEBnbbkIS4Bz1
nvxe7zGqNkspRT1ihK60tKZeq/rzLnbOGk0ZFmE4nLn2+vfzZCDs5MfPzrSEoHEA
vlW//xpPQm9qPL08Lb549q6PQ+Hwi/WuX1fuT+q/OEo14JplfGwkUtIm7o0xGClV
df5kA6PQpaKLLeGOloIyX1YxfdSoap6DfVevSSwTycRX4Q8ffFOTLwdYO+RRCQcY
Hbyl6is3BsUHdh6SeTt99Lp4n43TYJwX7Zqwobj01l6OzGPO/7/3RZ3Z6eV84GVb
l3ZjvHCIFXbAb3v7tIVqwXo7KIy96NkBZX41frwT776ZuQqlztWaGc3i4XVgZHUT
fD5QcwnISNQSGvguOY0qxBMMBXSix5sLs/IfpVyOQE6KxA3SFslFT+Hzje/v8uGl
s61HSb3Hi0I5/as/Y938vtRnn8xePqIL5vBgizOxhFV1PjM2K47wBkeyKm5AHE6v
wthhe1fz6JdXl/E8kAdZAD2CpN5ioRoyWAjAj4nifMWTg6AcqfmwdYaBSFWpi8Sn
DUs8G7fgJHRI29uRyssgrqpPI8tkelDZG930/nDQuczDSxqWGicNJzgfZhZyGMP2
s3q8RuyeBoWrQvVci/z/+zwvI55x6wqiLyAr0yiHS3NinxGKDwsWlHaBnhUKyjoI
ctkBuw4DA5vRClWTX+rgVlb4o39LlKtzSdY77XI+wq5R/y6cqbb2HhKrmADCPVIO
SOrLHsHsLCAoY8dtyLeJXqk1+xn48tzbY0P9DMPaD6JnMK7YMAhUWkjdeta/R1rf
bpWLoIK8yX4L4TU5hODW0vCZHMIR0VB4YYTydPNgOP/pGpCVlZeup/bOrFJJPULU
YXBoYDwQMOoncDDSHZKIMT1d8XlasVqYJWUKpNAz+QuhHKgqboiC9HknE8kUJPLb
lJ26Je3UCTWKe4Ao7I/HZ5CXJUW1gsc8N8QP8EK0ynwgILFeuOgQn5dXFINbPXus
rmGrKSRVxYoWukf0P5FbrRv/4VHiaiErpcjtxZEAQEuksV5lZ9FXbvjIblyLk7ve
hjNRmbYEQMVjGhB6ABIDyWUWLa9tjnr28IUbbIEe0S3T0NAUh2Y07zCBIGdIh3Tu
3GNtrUq3eRqNgtobjm3ODDc733op0h8QytxTaHSjXaDMIRhhCkQwF6e1E1fxL81Y
hMBNDLBJZ3k9Kg6psgfHfvPNviwRMdkLdpgAk2qu3Vr3+MlMaCjoMbLq+RomWRbD
2S+grmlOrxOT2P05T2V57nypDaCu8+xgIHmnvI96uIbWJvAEXLTAz8L0RAr2sAu9
z64dkus/VhkKTozLqVMpVlP6nVqp1H4cAbuYOeqNGw8GeMYftUBKRyC15FdvY2GT
PVNasDF+B3g8+pqZVnhTFiHhOitUN7qFjzauWKAbYcZuuNH/zVuT3miOT7tKjz1R
h+cRPRidYTpiQkP+wzaXvFhcS3jiOniqhZgBvkmoamZCPd9C5nFUOvN2nBZHMsjb
uXIn4mVNnC5EXpn414etpv3f4NO+1uqMAxMy44JuE8c208VphX5bdSTIiHtl+8OK
LOl08/s+W90zq7a/IoMl/ZxPVfpmI1aZPEHuIplzLH8nRQkF//fjc3CXkRzfvPF2
ouH273YWjKNkUBltomQI1u0SyUQWB2K0HXC75P6QL6tC9YmrgxPjbaYY7nbnMRDd
J1F29k8ufEQbamKyNXLxQhq+p3HS8fj2DEXfz9KncmNcNAlvrqRGKTb9vL43BVK1
gLhh4vlg++coXaMTk4l1VyIH/QX0aBq8iQ7C+k5W3ePicoDLGV3ERU/z+DtywzuY
BQSKMkFKaPCBQHTTZ/JjPcAZo/iKLJ8ybMNxdYdCXdFloArZR6i09ESNMYytvcSo
8nld5pEhSaYQFLtgRQ5KP43ALFykNlA7jtIT75dkKBJVl2RIPGENy17jdVghT6bO
ouHJE43tPU+dLWq4NaioVqoRFF2u4Nua2pB5Jwr/J36T8ABN2qCa4BHbbKAbAGJi
asaH4rzpLyPbelrnLGEtozWNd51DXgMCZA6oG3W/f9BFp0PKrlnOP4JQUotHvpSz
uq1i/PuCpe3WHupA36bLgFymjjpWHT+7JFYFc14D3Dkzy9eTe185+TH02/lQqZIh
IjIx/SpgODETw9DUtiuhkF8wMfvN8eg1yOm3iHUZPKZxfRSlIzDQw7GJEGCkNG2U
oHDt6DchecIk+fVp42isfy/gykM61czAlX0gcCRTuEybj4zqQlyCSYQIjbakrM1/
i5JfhnhL6ylib7bdN9hTFaMusSaMzvt0fYy2ayVtIB+KeNPtqlYMRep9ajTsu5yw
l5VKc5e5DkZjTiLFS5OI5EFsBfJy2OsukHE4JApAaOsK71/HUUTegVJA74S21LLU
wW3tzL39eY2/eeWYdrIgy3vNQ7bxeWI2gwbI11gAoFQ8FXOJ0zXrJft3K8JsETed
BQpheNA8fz/Y/KxK9DsYhSuaCzgzZQOlRO7bomeiDRC7lBfWTF/bMnNIaf1P8YbV
mOwufcpyXb5f3TB7pq8mbk+ALHK6tUrWZ6ENVI8DBBacxUmFn+CjJKwRoDVe6L8a
KM++ci2BFbbmx338X1r39Ez7VASq1i2PyH6uA/OxKsNADejlCjZxxql+OG59JEA/
ffei10N1+5jSmMLtHu/EKdwR6VzTpzv87l1AceR3+lQ4LJfllHgqHRU+knrelj+L
3EUvj7EPe/k4N2enw/iUWFL/INzYZ+XrGXXN93MnkD6TNEPGTobFxdOjCA6bTJFV
6vwmECwAzEnrIAKQiXuMVpICjvnDrXe4WUjaEuvA/LM/lH8shGCaHc4tLVLhvMzi
5x1kiGkQWGRxLwiUsZq6Hv/l5gzpiW58xyT7kMXYQzfGz4ia9O89buFZ4j2Vfe1p
i7z35N5GWPAmJVTUIedU3BpHxuF91y0/IfmywNWHSdKVqVyQhL/IrbGFX2pAQW2m
YIF0xKK/fbF5WHVkvS49CtjDJhnEeGOiDowUeo/2rOH8vneMhnthv65pJQI0AXjc
Zy2Xo/+R8EirTKygPNImddtKoQfOwcozNNO3ZlwmLkyFHDznywK8DaD+R2jWj6Lg
0THmQ33yztGhoNjCRoamXCjFex72eIwJgyWJW3+aMbipl3URWJ9zwrd5acQDrZjE
KvDIUaj0eTh5kcJInObDe+GrmMk1h4l6UKMInmCJ31lBHM2ZDpb49Z0OwKGFx0aq
hsQaAJnrkD6Z4hMEuBiBYXsubG24Tip7u8mS4LKakJ2By+AfllG8zctuRCBIgMRe
0ZMggadUyevDsqlmkxThZAlqtp7vp9JGdVsS8khr3iLefJbQrFzkBIUGys64KVjO
+zwoKXmyzRzmMTOdq50xR7Il7RP8fQBjdrJpnflaFZ0726cTGxABIyf6Kt2Pd50Q
NtOpaj5f74dYMHrI7eNepSf6iEcsU36EnYqpmBanOWeLuIQySMRUhTtXAbFxfLH5
Ao8zY1dO13wWBL6MI64mMo2iq+R5g1X7Y3WpsJxBk1OAa02l46mr2bWAM6Y6Xypf
h1OTIGfZXK01MZ83+yLA5FcIci68xCM5DqOsNZwfFT/y32Ag9CuRCoxG8MI5Xrm1
MbExNZxq2zsua17dLq3mUR+foM+xcx6hchKRfQtGfnUIpc+zxlQp/tAHFcfyxNsu
dsO8U62vLl+OqC0DB5cw4U74RX86E6V4tyIxC8RuwxxQfwMxocRRKRNcZs1Mtape
3D13NHLyAq4BKx282i83TvLCtoQs5v0hqORKtSzKxMlvakfDKqtYohebQ+QG2H8z
XxPbpf2oRPZfD9gUnk8ksXU39M9yQeCXmXk0o4BFusyTU/GI6bv4MX56Fxzj289N
N5ac307gSo3IMoETGXR877ixRJBgwRd6oqP+c6gAnWFziZNy0iUKhkzuqEarEZBJ
hGesGkbDLbNSARX5b/I2re6wzAbefH2ozddvNjsPvdsw6OpPUnfc0J/DSJJOujoc
y1mfJtyNGAi3iX0RBjAbvSf2AQpuNfaOizCWEphsGqUURsatT2dKKoAHRtUHuFME
HeSNRKi8R2SZhcZdj7iMuKuQ46UdVN6um/eqiDxk0gLxYOOehkgVJJiwIeJrUpSH
4Bp7uqMUXpWS9BQFIkI4BqA1rdlJCdL3hIZGRavydwl7YN4B8KjPRPRabh4wMlGy
wSE2qu+M5yNl1VE3ppcK0ed1tpKPre2ojL+GvI/MzxdtA9HBpPAdMoPOLnjlljuq
ABwXlrLzAabL/DmR3pSxtl2gna7bYqxqyffglxzNxkIkRK6omjaJg3cGqGRZBNi6
tY6zqeO+50gFlr45IHgoI00irQL8pQLe6fc49Zn/OvEFb/59lM6gU1vAxu0TFCnl
2K44lz+tRfe8vHA2fcbN3ZWwV7q8MCRyRgCdYXs302oKMam8QzMbpQdJ4Rf5IV2j
GreMkO7LQu0d8zjkkRLgayMHrbd9LfwMls/Tnvc7rY1JGbLXRxoGYypqlC4W6KLP
pHeDjQ6AjVM31/9ZhwmZniinm9aUFydYJR8jK7w1tdRKuWMwZBwcTLya1Zbq6aj9
YFaCLvEha3udiNjgoT6K2/CyH/Bqn+EaFypUU3gGFhfmJncaFslDwzHPcjjzgsgl
W2oE4YuzxnWpEz4pzxV6wu6/KfTOsEDiA6RT1oh4HUGKJLD/Cw7pMelnCvN782hc
LPuac8mZRsesCecyH295JB5HRbK2r0ki/wxiJQdv2UIiJOvM16fSwrJS5xf/G0ed
qGVc8isprzoVG4GarflZJuIav/z7yWK84GxvZ1GRb5g+KR7ToXZZc9eFeabwG5za
1B3TpYORbGhqkR2gs8FZlKjKuRDi/D1lneKFK4VOEm+7D6adOLHAIQPdP52OvBCf
BH4p/4IvIzqpNO9aVka0r+KKHvjJsz4BBf6qRsCNYmMdS538JbgXjW59q1KqXV+6
v4VG9W+78aB6B2srvN6eL8/SmY3xrHDQYvqoGGpOd+ERmevIT/Qc65FMdWmHhF9s
qLcVVDpFl2ZEB5v4QqZpcPgcGV+pF3T8T8p+E1wWBky+qUEy+f7BWRHw6T/FEbdD
gs/MOPvO6sdCWSa3ct2yyg+zB/Xfdd3+6k5hnSky9/77U9yG3q+bBpcanSvUqsWu
vMPnzySlTI6L6+LkPtdrPhNTTKEbZVJdsYWOzuwuowf8NRTzRTciICiXCZ3W3I4u
JZoBierC0n15rV6P7jbB/sOepGq1II+pyAPcwTVSrkq9rXWfFqoFPAyMS5QMjSnl
CklE4B1BfUDKGvhDlcchxm8Nr+Az9y4QDzk8kUGwvaKtWrf85cUm1DgADTuDMbpz
BL5gniRMMKbxkSKMhNHZzWNH1Fpl4pCSecsN4yK31rSW7GQW6i6v/LDYlxozthNl
0KApVitTpg7jdBUbg2SWlL9RrrzYdSBrCyXkCLQGk70MuGBpxETT1jyVzcgwkbEI
zOixfOgE18RD7Z6yJjc4R4SGRuIilm5GPH9E1HwL+r68u/THuhbcbt+9MPPddd2L
FLhKwj2/j40NFQ4uGByd/OC+c39BwW/c4CiOKjC5cGjp8r0tFUvyzBEnapiV66Ng
wpHP3aJV3kxtcQnguCm3papZVDmVqagYAyTFbGKlfD7PXD0A4ceLrfJxyH+I4UWh
3hKRU1QnSNekwi3uDH4X3Sl/XRw7iaCQaTRz/Rox+Q9W8C5DIB3fwaE/tZ8kIpJv
Bmcgkv8X+MjrlivmaVfdEwJ37JdbEKB60GglG2sHV1QMVQ0QIGCcponUl/IEZmLC
M+cmAicGdKrSP4kqkNRCz+XcV96BJ8OvDbO7nAwmgIrvjyCgkNAhVzSSmjLzqpex
yJsQ0X3tu2zxOkosVRAuvMjcEZNTzkx50ECWGfdO2WcS65Tm36wGyGJW0fqh6lWh
nFBpsZMdOJ+kS6v7GT8fBImuS5mOiAdX/raKPG/PezD+JhCJ9YZikY4AEGBh7jSg
Yu4UWMXA/k/7uyLRkeIvIYw1q4guf9txRQTrs3lVeTYT6HjoB78kpKQGA73uCER1
pj3CUyH6mjlplTiU+nzBR5hecq21XAQ1yTQMb16I/KiXTv30eJ2silCM8f0YbFKo
xiocNvXtWqaXUHEyVaJRvJoU8sMio+My+wAjRjbBYFSbkIPf01Y3Lftv8PF3vrMm
SCBVsCoWbddIWuyk4Zi7mprvuWkpg6QEq54plGoHmkS2+rERtRTB1lq+ypeZVVFY
6iMGseTYchpdfROgtjNbp3C93U1hPTg0t+Hb3HMSFcQVXNSgwOjF+uOHIJmPXcbu
8PospC0C2ODoW3sV2paIAvnmRHAb5kHFGJJtivDhnLXmujBo8WzeMKGyWRPmqgaH
04IM6atgLHusrU1t73+Yl4G1fUocNRUkyrWUGQJgdVeTgY828z+aLh0eR37Uib00
k9whSAHoFHZfD1mDMI/eolsK3ENGzMIlEYBfuhH7z6atrYNfiU1E8gz/Y8M/9unw
rXR7bkeVn4WZWcIGcvrWBsa/6q96xV6GDEwq+xUpIE2SpxbPU6inJsBAE81XWo8n
1BWgA7Z66LILe9QIVcNMkw80jynVO2wuhJg7AXcpxnKhvvFeat1J/ITVolJJxmw8
Ky8ZX8kcd0o56vIHACZTmHrUjUYT21iAS0xNRx6X4SeTsrtZiPeNvvB6ij2gjheh
DlAFyvi+qm7Vh/23sVCNH045u9nB+IomctiqnOEWcgQs1NZ3Qf2LFU/5aHX7ki8I
6uIU21APoWPQLn5PhkBsyiLMvHsKMmmziLeZwr4mG7RjdVXRQ5Cx/guGzhN9PcTl
qdobeG+849yQazarCdnvkZK2BfMnnNtufUHt10PRzH/F6aBQ9ftEmreDLAk7Ef9+
n3ekP9PgB40axUOi6QGfCv7QJxW0hruObN2QuD1pFvJTn/SCTYaFZrJlCxPkeyGw
JXLaaWmjaCqRBnOTFOZRb/VU446KMdL/GmPe//sI0hkKbs+p+WLKL0sZckyZoiEa
RnO9LEC4AE7m/AhOilGgx3rHqtWL6qevBYYougMYo4dwEfYHfA/47lm7Hhucv1Sn
XAdmtkeRwZcqnwoZpk+Bz/B5sicTSmF+68L0hHpR9HMUy24+LHJ5u9J50LE3OWJT
CIteJ2lebJxfTH77Xbu676T+w13rQxhAfY5TZZ6n8Co5NVhOkunRTv8w/kiONXb2
w93UeO2ANvF4A3VkVCytrHcKyp48ZM1Uf8D0lh+wf2c7YrjBF++SQZaV4hL1hu1C
5hCSTTXx9Od7m6b2KHWHFHSNJDFZ0CMsc/YY2TRSpuAvQJgMz0dI24AqObHOH1vm
Dc3dbnvEtqZY7hUD2Gtw8CnoNJ+JPohZA+gmQf320D5xK5WuhFxXzq8KzhSpmOkC
bZ7s5Qa2K8ALBKS2Rts+TzTNXmEs8tymGuRKQZB6Ju9d/79jnd+FFrBUeDXXf1Nw
xjCo0JlzQFlXWhgVYHt1jpqLS5Gkyr3pggEK6rTGXPZypqvsk7ln2EJJ6Jcf7w5Y
0Mmz7CCwKyndcZD94y9DSwd7zrUazeUXQpbKUDwy4WCyqC519j474C2iJoKMu+FK
QMe2ODc87FenB5izn94WnX4WhfzIo0pNUGs+/caWP02Ix6XuFv8AxOH+5ol4WQxw
QOVsE/ZOR5dS156dx+8ctkOhBde/hHWUn+bpwF5AWpmlfwZPTf8OMvWoflkrgOmh
tCp/MzoL0eptmC53uGYlp1D1cZ3Z9ZQNR4feggkHE/2IxLr5AnQ19BeV86F7ctdY
KMGGXGEkUQ41PkLv0KDOH+gLYX0UP5aa+9T+QAIgjhcujDVaDLPGm5hY3C61i1wl
lclw9EQG1PdnyVxrtWkoR2MJC7sDji4thO51zalir0F355cvIlpiFOwnFupO0tkr
HRg0Y4kFQVh8Yf+3evPVT2TedcK47Co1+CreTWOPk7+71iOSjPb5xsG6/grvC+X+
bCOMDPZNUZdl5aSQl0gga8e+FjEj1NI7Bk8gD8SIfBYoTFfxmxUBbBWVyyz+j3BB
qlO7pA5WA7p61fJV41jJq8pFdRa1Q0OEWqsvmJxBR3ejnZ3XyZyJpyr0HezyESNo
79g78BcQEZ/GHjsUtIWbtT7pEUBW6kyWySwpeqYRHPBHXMZoCWhJaQ0gl32a2h1q
023F40joZK1zs/AMIee5tySpVc4hhyghL/00Zzhp3qsDrLczDKqP6Kgk1LcqEGdb
TgcLncIv7aI45y1eXNWoZshQx4rW6LBigbeBa4TF+/2U0dEEWAhP2tUsD3y8hb4p
diZ8viKC3iEG3P3+ScId03dPMe1rxibnT4FB4rJUB0erkvvp/1ztNQszQoicxUTm
IqwlKYpYw7g+CzAoUPHSByjOM52LMrwHfkrO1NviPXjQcrQ+H6zPoBCteO2YGvL+
2O/DFOWSBMZhWZykjyIntTgzzm5368CX34vQQ96vixFXxrqJV1atwqd+ZZT7wiG0
6qh+lKRvI9SucwVhHG1oCM1pfmoSbK62SdI+aEzmquMP9936n57up1/mmfUzEimp
l9H48h4WhU/LDwh7U/UQqJ/tGenMcM9ctRMvxy0fpfOe51qmi8xWPx2AQpdGDIwU
ZwsvN6n/dGVM1RnqKog08Ed9VJWgXoU9WtHPoRntyN1nxjSBDCbChT9KRv8riPr1
bq5XH7JISIMhUweXcTMjLxvZIzj8YpYa5O8WLIeAB0OaM7AKxHbk8Zp4z57yTsRj
1OIMYSVHLe0GP43I3+tTRIWdsBkjsMkUH55RJYsCHPc7xVoPEuK4c3heV9yHq6BB
p6Vq/XkrybpVZ+h9QJn+6QnlyeyusUCqA65ChYdDgpIziPgPk3CGS9cNutQWSDyp
Rmg29W5YZ1JLwTwwI6GtCjoxmP4ffbFg76UO0N4dtatQoINJAoD4Q8Vn25kK1kT8
qvgts9rHhp0m/dQNM88rJin6QejCTg68A0+zzra1TKfgFaLlKyKXdmZ83iCjlUh6
40NFTIVdM3JGcPoq3vapj23X1NUnXTFOE6WKq+XcujRBaTpJ9UCKgKJCvZVS7nmA
GZykPDnBthMrxP2z/iYy4dKBiZEamyctrc8LFrvEQ+Rn5AOdkLYd65eEPX/ZkHiq
6vq44azhwc/Tpte+60uGmzp/9qkvXYRFgYfpI0OEEqevC5gX1ls1hllzUStfOFW5
YBWGhbUmk0VrSwxlbCt0xMjDelW7P9LhNjISxsv0YR+yxpVn+SIeas1pX+AJcEn1
Zy5Od1SMh5jVh5SYDnl2uN+bXHfBK5E2C3tpyjxQaBlEbTEeqewIO3M3S0Hib5II
4zfUHw+fRLQYbV1cVxd5KcAq0VOcl2MyBFB2abG2ZsysaZr5Ll4Fs8Zz11fW8+kZ
0j1sbwwCLhefbQlmIHvoisrsoYQsfHDZdbCcRCepZsc204oDm38Rux6LXxsMs4Ng
25/oM6u25dHtlPAj0uWL1mWnX7Q9zG0zGq/nQGbPC7FeDFCIr3w20BLBKKJg5vLS
qfNaRu1CAvb2XNVC7lNX8pKCdeFHD6KGO4GrTlz+er2PbUaVAijJGClDmq9USpIo
sKI45PzUvfNoglntXoIEkns0MvunnXO9MGE64m9pD+bC2s7sMM30mgfih+nWJDsG
8jqk7wJ4kTpGbBa41fHht3LxStzPW00euQq9kpLl1+TTsiF4bH4uOtU1c1GDg/kb
yY14pFYt46v38R03l3ADL+In6eVg1Uq9BgCr0hsXxAVOoi0J3UkCUiWilA00Otec
RgIdTTvBrhXbIFSGsVqZRjOS+/geMFOyE6a4565ql4d31n3mwKZjS6RjriK27F0E
RfBd2OVd5tH1gEO4zftC5S9k3tbSAjlrpSXrC5bd+tHUrumPQFqrXP1g87wiYp00
BAOabV+YbONSCWBPrNSuaaCXHgDjFE0BXVArMHtrbNIqcnfpCloKVaD5jL8l/lx9
zDC8Mt7FDOR0SYeLLpwt3uLRYcSRLx3oWfuQxEO0TLVoXv//gMrj/AfFybv1G7zt
W6pe0kdICtc5JKGFnboP77oXNjGF5QzZiz0lo2ziB0Lgf8/G0YDfBku5oSFrLyfp
Cg4VT+dC7sYwZGgyoRr04Ldpu23igZpailjFRbKnolt0E/ntD27+H07lfQtVQFPV
7UvSCwoMCL+PGcMj9ys3dN4WzJ8UV2K6J8Xlku//5pHoY10GAUKeZv5pl7kWvYQA
uZ4OKY3llyY153NPgMUsYzcWv/zWczZkM1U0tLbrLaV9T3ccczxYKqZozFV+SmCZ
ruBgUb8gz+8kW1/LsceVng3y9vwWF8ajwvjXfZ629pSvj2c6czLZt9amjO8LiMtf
r/MoMplVcxOuZb4zNbtUzLIdoH6kwhkZe2zAVUJsB72lqnrIm/ajQ6AnvDa1RvdF
86EXRc891S9LkZt2FHP/aDcMy/cfEiMTQnkVNVLlx0t34s5iu6YWNRkBAximOWIs
38LaujQdV5mFJAog5d7/F6TxBBmgZFCFUt0HRhEOLfWz5J3N613PFWg5EUbVhpxH
1LbFP+x5yOObm3qKVx0ktu1t1Xo8dSSghFJ5q8CUmv/x3ZAo0RI02i/5OcnS5ZVS
Lc299aD+ZfQU5TDCUN7ZC76CN7OzLLNL+E5KNhbjVkZ/JCKWuIskjHNLNPpKrt70
aco59IJR1iGwRPeHTiTtTWpUfVRyx5Xq6zCRbGrnt7YA5Jj2GycK/n7IWeoWeHBk
N6bAj2Co8vtP6p3gkIlzvcOH4iOrxHHN3z0R7geeO72NOSbfuvJdLUFngXln8sCQ
yj+xm/v6CS7LQIAOz+WMQV8HNQ9e5JRnfgnsx4Quf/9papKfXEyOqmRKptt+1R6D
QLOdD6EUeMlz4kcXDYrZ6oaBKD0aTOeHn+H4WLDjH8PQVEXeDAIf3bAvqLYR1ona
zX4Mpxv8sx4Mh1ZSqJN4x6GYuNIG/sNcQOUaZmOwW40nZ77TxRZrDdaFpQ+HVCkf
qZlBdNnCFHhGdrcbixSbDo5iLk1RIRDXexEtqzqg1I1C4zSjKztr6tzFxtKnFeqb
FCSpyhcSApDjJ2W/4Vpttb4s/q/M0XBSUhDvZ1Hc2RdGxNYBWN2lqJE07cqITGcd
G7rSddWpSU0v9aY7z6tsFQ/5SOYdGlqWo/izNRsas+6x+aVlunYe+RJ5HnRJCY7c
QK7RWPD0KeG63hrs/DM8w9wWYFHX0YIQyQH8etIfraabHxh3Rd959fPJlqx03ngy
5Xy00U42AaZRkf7e8Q7EHkD8nfgvbLMrhtxMrQo0qRYZnMK+Sl1twOO1R4LvkAlJ
vd0H/uAd+rx+v6sa+bhxu6VLi8ItoBFHjfkVqJ697g1leeL8IUIvgdEEwhSZa6tA
Zi4rJOgxWNIUPdpqlCIA4G5j79ajLsDby/iXbtlIx669luZqAmwHivvri4JVBFVV
Db913req1porgTKR7HZpOy11KK2L4VsDjaN4VrHTlCeG1Wuj3y0xCi9aRqmJFhBJ
w+0b8NKui1ZdzFtWQjFBEMrrl+2ttP1Sq/twVLzZFxVbCIkOeQJLZvtvbka3CWrk
1xdk0Koq97Ey0CnAehgYgQr50HA+cX8ImAVF3cSJGn6xbXZlBxRXqJjm5ZXR5CsI
fk5xsNes0nGcdE4ZwTw+IkjO6e+ORhn2VgNgLQPltKqfUU0Q2j672C9xxLmh1DCe
sLgytFS8m0wyPo5QdlRmXYe9P4lqYEuYq4wQBCqRlejGKEEbqUM493dcwlyns6yF
Uh09nMb1+jr8mOa6Is8PAAQKta2jVJ89UOY3t/zQ/p+LuZl/Vit22iRbII2pd+Oe
xaoZMc5aTiJ1sEx9KtpxoOjnsCBqm6uYoao+Wq0I7DsfCtAxnkTC3zC+K/aZFxTI
XmQwOyQj3o9PaWGGN57YA9OdklamBepNCxywxzV4vOYe9y0pduhmp26rV2YJVpta
xGniaLX2yZs+n/nQ2OoQa/1zCZ03b4EKBvuxSg6D0c9uA5CC5b5vEEGdtLRIP8QK
c8MqbpHv8IRIehhpJoPtnwmuDTh96Bh9laN6++PwhMSZRjYBqEI2fRsRI5T5TIPG
BWhXi26aZgHZQLJeXrBd72OyN6g1DJSMBhj//k4sZIOWfeYxY2h1WtXtHk+FYnmM
0d+ZOttP7uXexbzRfEcpZutjG2UeeguJhS0yxOcnvIhnWOGnXlIju+zhvDc7i/yX
f+wzGrRfkxVpAaNIpiWOdoJ5YsPTfze4jAtWxKgo0i3zPucJYcswcOZTSu+GvezV
wjwiGQfJovDRlu9vmj55F8Kq30u3z/VfH1SK61uIDJDYKRxwMaUC/DDN0U8hhV/i
jDB5TyprTG3kYj9j5jk/avHkR00NDR++Z+DGTtZhSdR7vVo3gmGIlfoc9AS5AxIS
J4OsFnDK5osMOcsTvYT1my+hZbgzVNt/qatlrnxvWmXWIGi6NTCnxitmitX7glfI
wGmfzoYX8Dk8Z4e/ziBrb7oCHXVqjs6EW0Ft/YlwnHGiGwTLB2KrnrIgXRx02tyJ
DxKomH+cfihUyKrFZJUEHM9iOERAOcfyjJ4s1bWgGBH0VpvZCWI7/lNOcRCvz6tR
CG42NGiLgqdAsnCNKubjNEt613EvbtlTll36EePs7KEG6SSKYb0IC2KzQQ7yEXh8
Eobnz6GVScOXeF25phTUbZ4/7WFa7i252bTtn87GelyNKpAk1sIgjGLVUdh2UzmW
XWlI6fOLb8ClKoqEqV3jmZiVlqbJ4Gw+pA4196lOFByssPaf8NRlRKkWll3uv8UH
VeqqN3weiloFOZDYIYk7RuCfWacEFA5UkD5mmYkCiTRi6JSMgsE2Nt+uDjWXCyYs
nz8kf6nim74HNz7TRS8w51HPOX+YNQDiUrcfqk9rj/Mlxaly4ORNkjncUG/4AhQ3
jd045SMx5wVwuP/ie+FQ7oACBik0nQLlAnNKd2YanpQa4HjBqoa8w4H6qxY+9XHz
/Foq1MN742IvzePoqcnDpRZ9XainDaMQtGa72D3UkOZjG3uw9nmpw5w5YUu+jmoo
MxH/BiuQswbWHmivg4KOFcxD8Smg16tBcVAvQLWrLxQ9DRPu/jYKLzwyobL8WIjx
myX2FbPQAJ6c7ziWYQhZfc+4Nrf60+Xtz65Apd6jHiYdFYn13lyeWgI0TfmjHrtN
u8plbLV9elgGqI+yLVJgsgt8sicFEKEPEENgSPmmutf+5Cfca+vd61L2os2kIZkx
vZLsyLJMQmoJHAPeo2xUYAIFeJ1I43Rr3vqv7LkA0ikNdEKKg8usPx1XLWv9UJt5
hhNeazx4t+2A7lyLSZbTyUKN4qqYzsvRZyrMfjakK7qpnrXMNT2VZIy7d7rmwjmz
te1Aomu+YJfFpx8TXoArlOhANVR+HQpqQEOhMYNHkZErhR07RqKDojUMGhWOw6d8
8ZS1n65BykPxLKFOpmCgWvM07B607+bLli06i5alRxmTf3SmRU6HhFEKpIWlQovd
25qwa98U0DxJb1ZB7nSTdUOb4Xku5G6gfhTu15XXjP/XbplvI6z5JdoEL+l2ueo3
wyb2zWRXWThFbgeRB5By/0qfQ9wphA/ZU+/pVoJ1MKyQLoDZWycDinmE8t3nM77M
1kMR9sQcgAg4HDnGzjbMwo1i1PX/O0lWiYYBtMxO+4xqb11p/IKJ932YM/oRkca+
DZ5xGNkLH87E9HVe90rLrWbMp0QqKZWkKQqB6ds4HYIWaoLuipULXauwVyLi2pYE
lYvvNYh4LGRqjjqJMFaN97hbp5XLeMCYa4nU9wEV/NqXFVpDC4ba+ZnRI+wX2Y4c
B1WzNhZqus+JmSTNOJB2/Puvief9SzC0KJo4f2imP1lSh0FJ6jie/TV527Ndec5s
vcUjx9+UdSswd/lBMwbYBbyouWdEXjrjUVEfPtTkwa5SuFQH0475eN+ZwlqzA0Hp
txOz52oSa8hh50AvNBdiI6D1NYt37mHiOoFT2oH7dYuvnrOGp0tBS2I0Hq/D+ltD
uPq+Mvn9MVrZvK71VJDKHljstvbMlUZp32QF/4OOWWigTkfCtZsxASzlQRnlm3kF
s2v9lL3VsysDEkRUZa16lWXaFaPzdNIH1K13Z7rh9CmK/gTzFBbqii+IiO8kjadE
jJ8Wy3Gbz7ntG4SDrebbzzRgbOAQGHe+DJ4RBd6Yz9sMIbus+vu+pIYbUm1JfUUC
PMFJnPbjHid24EKYSKO5wRe8BATlnA9fdLJQMxlTQDbIGte1+O9NdMv80e0EcB+s
y6zwTAoS5fN4jJgtW6enoNFuZkGRiwZQjc39uVWWfMO5ofWcDUb8kb/dmr0gobKP
Fy1AidYERVsGxKw/XkC11PBqvV7qfSNlm4C2IcnhRWRuQPNqq5im0d1a3wZSNkwd
AR0GorjK99jjdN5zuL9FOz+Yb25LUHgSg0dQDcGWwyCAyA74KVki8On9J/tzgtUt
eXbzeNDJC/zUmag+rH34zST1MJ+cgcLm0lAkjZvuHuInGVnsyr3ohlRFM1amPJLX
/ArN1TAJOdtP/hVChuUAWxv+Uv3nikKXnPXkSTB7G+LxoazPiLSCO9mGdeeA8klG
e7t1WRJU3+G3e0HipTI/++dQ+YK/oKxjJqBbAeW1gywoPLpNdrx9SqrGun4pd0u3
w4jEBy5VKXRS/H6jpfU8zXpDAaEvPLqVTK8XPIKxS2HoeMel4ksCkUssWdKxW5BV
rrS+YYpjqa+rK3YlWkvCc4cyehdnDKZGBrjoYXRCDdnoWXejs2Ea0+PP+9EfQTmG
dTYUyUCmTDl2RwnlKn5VAAcEpDE2Xhq/+lemDx5aEJcHWTtoTDDZMXNiyhf1R6zz
SYyDvTYp9OCSQu+aSl7VaY09xXyynX5+imyCqMrEocKs0q+hhA9+28XaXWKGsHQV
mh5I9aElZ3Oz4kkXHsKOEVybnRD2x539ifK+0sCrsaK54fx19uV0+q3JxH0KMSii
D/Ggdr9YTcERBp78Corv1r7M3q3mV08Dcc5lU87/rhEqsskuGT8gSld3n1x3fsWm
6IRIKLB/OJMiZAFrraizThhFJ2xrjZmOyisxkBoQH2Pf6pw3YpyN3KcrqjZiowG6
4BP7TTc5YGNMvcs2N9fHYDf77juCofhxmT9zbxcUucb0miteX0a57pqpa7qB/njH
VtrL2NC+Fkh4WhCdrcFb09ZJW6CfIDS7J+RFspGxgaNk33PPb32iSHgwqlqU8HsP
Ft9h4eAqG+ecb7Z3cqq5OkoFwHlitCdh4pW2Z4zGXPaxRR8OQiY3WQ4aHuHHkfMh
WVdqJTMdupFOKsrQIcEzxQFbIvwHqZpKuRssG50xkPbGHVNcSyZf2LZHM1xtBLy3
qNcACuVzJcpmPjTPul0NsvOL2Ldi5/ETuxy+ws+Vb2glyDlNOS6Tjf7iRCeVpznd
Zm5zUVj/ZpTSBHkK4f+NrqmbAAymC1tj1bmsVhpaEFLGqKaZ8yu2q7b8/YaMf1R0
6rDT/1XicayDSsQ5n1Pel5riTecrFQ6gqEfBxI0oRJsefstlEdw3sFbRge0tJz/y
ewsF42D5LdPxsbnNDhkjT2KnKUHUxpB4XVxu3GJ0MCg+QSXw46bSdXZZzQHORzyt
qUAVbLJWX0V6PWKs8B/CbUrgmbo85ez0OcAWUr+gUBkQsm9GensBwclxgKHo0Lxd
CG0/UHfGKqcPOd8pjllSBRMzd7kc2EdMyS1/d21rvfgss+rp8eg8chjaMmUPIDER
6Yyjr4DBD/a+8qfQaPwyYoHNaNY7W/ZLWzrUpAWipjcY3Q/8AmWcAMS5WJJb/fjx
215xsO34/+Di7ZIq0QPQGMv+E+DkgSoPiGEmfuP6l2NBsOHo5ArexLRxtcGazP7r
GPN0+0/IW++iK9S1UKtxrAG+oiwcBA33NEsJ8+XheDCl8FRphQbstR0x11MzWsMz
hhYWgwKRrxe0qSH3N/I3dCcn6BoIb7oVLHV82vwWoVV9e/J1dOomf8tEgfaS7eiK
KcbZZPI8IrZNcU7rXgxPLyS8VUlFO3W+fxpQW42jzBWM+3nqNEn77bD1tvSW0rTI
42Ld/NYMjE8pbgtFLCdkkLunQOMG7eqAVKUZoaNKp7xXR+VNQKQMhxswfjJbmfhD
no8d2BKChh9IoW70//J5Om/R77A1EaqQu5HYfZeO6dTGN4AIKPcunTMqvcXwU6DO
nd9ZYwHNBA5C1O4/egSY2aLpr3KAYkf5mNlz8GiyJRDXQcd4Fqz+yPiwvU6NvCR5
GDEKO3lk1qC/h+ZqtFPub4iXyx+AcIhUPS4p1hcY+mepSZ6hqy6uwA9fC5cISkVt
t0KtqVqbci8xArjVRJcPJ5MaIZBYJdrAu5qw3/x1uZLVPLOFQGCYqJ4OQg5hnTso
3cl54ECPTrEQSvhjQwy2jQv2+jKk4EWkMrhC4pCL7hB5JEFgS3nznQzWV8hMxzxv
S3A20RWkaxopW3eB2jCOwLua0bqJcmbCByzkWRB973GiEntB0YH9DauFm8mMXG22
/btXd0QmIfZpfnD8+nhn/n4Jbojzqto2tyI58EnUwxlHxTDRs5yGSdKNwCdfa679
QDKUQozScp3hjnba6P1VTkLrrm0V7W6sgMssLZbDed9OxmdIwgmCdOXbG0cmJd5F
6LjBXM/yDuwvbcqMCY7KDQgXGSUO0nxJLHXl54Z9YYUxAiDoh2pEoqPrpNnGec2X
TXmMQZZXz32GaJ3IfgX0Sjhww6bVKYWGEnOMcINtBF7+8a8ei774edYN5MBQ7ryA
t29sMMorSeaU/hPDV4g1iCN26TI316XEWZDPL2qe3YbJo9BVfU10sQz6YM0jtb1m
N1WWsszaS6+TnIrcnPiBT9/7G4wfNQv0rzfHJWRvIEKk/H3p2EAU3WVuTYXLTjVI
SMbCOML7FqxfhNSjTek+EVIdGR/V7hCoqmKZoAQdBUzaxISZwCN2PoqLb+g3kRkZ
p+WCMF/U7ehGIAqW9oHC4rQLlXPmNiAbnFdNIg3ZSAFXzlUOWsff0w1edGfyB5uY
jZ7D6bKypniur0MBulDmSnoKZWydOTcEmDw2dt1xnUzyqL7SvfXETTfo3FSqgCra
wJHXna+h21y0w6iNUtQ15daAQ3RE8M6tyvyFj/w+7RDRXolp0Jl/Iy0uzM2GT14M
YhUdLh42qwTqnQfJrlHxsYcgLIcHuwW4eWd1ahyys04cAwi16JYUgxHiosktmYFZ
68DZKO5AkEbRbtTXfTTrzhPGHckmDt4TclhCh+PKiltlXTBKDcav8D6dcz6KyrXX
OJGokwZU71Jga4opfj1+niPFleYVOxOEHNidgFVIL+zK5RnQVXjB/W80unr1pX36
Nutc1Md0lgyU878ArrP6WcsdC8H56xJowJ6DXgWmD9vDjjLyv5ktox42aEPrEiZR
SSwzkn+bdvQE2PUrE18hgRD/5jLKrYknCwCeaze+U+NeumyYlKXi6UfIcqB8XNoO
Mj8OizH2g6AdBUO/xXvI6+bvxBuNBiwVY6BeGo7jiKyM1est8KR+elfsqg4sRbtb
OasikWJUI4Xr60FLykM+xzirdxM4eHP456NZcshioLLOgSZZnQEmURfmKzilWp77
jayt8R90xYDegFoRXQ5YJCpSNk/JUxMHFnnccHiu7BWl94hmBd9wDdu3AtX4AOfe
39d93sJgv7PMJjHfRkjkrY1WpyV5Armzqx9R0T440F8r8lT6Yo5Lk8IDxQH9AN38
XfUJ0419kf/117mMCE4FzjlbZMf1UAW0xaLWLisrZgAqgwwGQR5SX8g7iqSOkcdO
3bzqFOt939Q01/B4vOCKaR3obOySBHJMiT9kjIcsCk1wZeT3ZBGTia+jE5QAqwyv
5kxKcNLBc32OOl+8XmhDXV3J+A+/KK4Pd5ZCxLw+KP8zkPP8IaGXw/3NkDD6qjYw
TE4fFmGg4CmT08nNGEoNjcSPIi71YAcUGlSYhy4q0GJWl+iDCwQ0ivzcZBW24nnk
Fd8afrLOf2BD6lGjWB0PJf7I0kPz5ndSr7PIv9cNcB4UfyCGkKMfa2A7JLk02pDO
KEX47h59DUQ5AagqSwOUS2e5wm0eApGG/jcRlb1ukStUaGg0e6mRJZrOGZXvjEVT
Sz7ReDi8iUKU64us4SLSsJ1ibyHlUa14y4suSeIzvgr3Y8ssLmgjIkjXEA90WbwD
9Fxe7dHaQ17mtKWpdS/gJzAMSBSOnupQZZcgWaxx0mnVlHO+5FhQLIWlcF+/4qcx
GH45ZOqwoIkyrzSe3lJ90tptk1Lcqboqiyf5gtmeajptlX6XfRkaf4F3fJSv0uO2
PwcKbFLHE8c+rGqXWOOEvAOemF8Nr/6jNdsCC/Lf9Zfl90TgC8V1OA1aubRY7KV3
eD6L+hSNk0YGfYLJkTfyzURvm1vqIzgy5RJgU3Or2vdmyLohTgFCKpC51tAQEudg
vW5cMTJpEE4jsSoFvEU6IBsmZs8+qTEcQb9XR7eayBXzOOkbRirJZk4wiJxv19p2
VJAjdBmSdp/Umt6PEZ4Kxsnw1kPWnwd/mOTbAQdI4Phw8aN3ExhA1vLlvVNVt/Om
GjHOQbNby+pf5v8mUGatTm7eEGRCsLBf+LVYjyEdtgqpxbu3i5ayuSlzdllOmZJG
H3OSSjCCsPErMkKCTtOj0jil/nfqU+VAi9ARpmL0mVeoRUS9TPaiXwnSk7s3nAhK
V3o/lNFMEatc4jApmURJtLaoL12QvjNH89wR7ZbhQCV2oTuB6BeB6KpZFXM2eZe/
bzyPvkC25zqfq1mHwXBMAo0dUOpr0kMlyQW8dzh1F9s0xsdhw4UJrFO1YA/4/Cbz
WHbB1W0eTBipsU80Yhjt6g/JpuxPrUWn5u7s69Z05y3nmquTSSEupqgaGc2jOAx1
zKskAK5fnlqVv5rYTEGXv4bI989Pg9J6dyLPkskT32uJTgeupwfCZsNy9OUJ1gVN
KjV05qDnzEH8Q6IX6fisGmF7iozQQ7MsHYkjTM21aokYoOw4yS+zHiPtMLIMVCIQ
v/8DjYr6K1tr25RcOaQmTV0wMd/oGQK7XAjdfWNJkWxNNVSyaotbByH3PfNZ0POZ
wvqkQEDdQMY+TNvF3yvUESmsEpYQfNBjSNaqbb0PtRa0oeEyJsUSQeC/P5t1TOXR
fBGjxHRL/Vq+tTjLY6+sxuN4pgkg+AoiBThLeBDo47gF8ZqFwrR1cctb105EF8zZ
psiOhz2f0kgqkTxQOAfTZuQlSeC2iMbj1zi7usGP6gzbbmhDvzI8tRxsRty7skWh
YGSNj22jhYCHdBi1wPc3ZhvBzJbi0XFn3ZA82PrumyyXobOaz+sEk9y46nOZan3X
TmDaaNwX96q5W2Kx74F2WHEzYmsdbe/s7pCLSKgxI/SyrqbUl3GT03YKn23TnTo1
8UVKgK0TTYomOR3pt3Iku+Xj7hmD1/kIydvhtbYpA16wxjdCtWYsWDi4GxoTt2aH
V2ZXeNwJyWDHPeE9wTMPuyo7Iqny9RZI1iFh4HyqcckLHLpRw02phJ7U9R+LSvpV
aLg3PyGtVrV7m1BMpC/8Uv/jSTCCKy5qizXWJ9hZ3EAGpNKjzVBYr/bw4o0Vhk2b
WOEk/utvX+rzK/4LK2VFzlsHNDaQkFa6MPMEwaIr0QkDiHczkoLugkH++TIye7JU
1sUz8IVCquSZJh9s+lhzGEEZXHRuQlQYffuhVNAarx+6l57/xCF+p+saZZEe0m2+
EcPu/vreDjihSPK0ir95/+b8LCI3L9EgJ6Ckhmwe4Iw8ubyxTjKD7ZwzY+OEWbWo
bI7BvHOQrnFskYzYanZYTTRYXImbc4rOsCztXK+1iTcsAKoJ4vdW6j/k3nNzkego
/nCz1poGOZ2U/rSVKhuPmDsLxlA2JWyk2XIB4k4tJ5BDee3yVlA6WcOdCTHQdoNV
/3NdPx/w3BnHj4nyePaX+eYFnx4T80iQD5xojEsoL5cJMxhuZbm9Y144PXPrjY5F
K8r0pYPOr2S0cBBmKnhjcK3PpTQu3KY8ylPJxfcc7at9wr42ekTCBSrqQ3+2FapE
TVXmckre3CodoooZhio8ZzguktYATfyLGWSxGYJ9TokQbZp0msJBuBM5Yscv9MVp
/ItvlokTx4OZrmlau01Jf0zG7hNK+GrHY2cSvkauxrHxoV5D7FWfrkWMZI55RDl7
c7QKqzp1BeWOpeBYxWVoLXohKQGC9wyad1LDs+DL92/RzLLcmMidOCQKYdiYmbdL
z7jokruV4PH6KNrR9fz82v3q7zsihHnvlpAV6BVNUMxLZXjQMv0r8OAGxumAQ7Bj
2obA2TiGPCx9KmtqdnWi+5RQi8QyWAyn8EAa58MeQDJKS6zzlK6T9NIogG/aR1hQ
HaGdGElbk2VIdC273gs6IghLmQ95/FBlNfWwo+vqYdSHB4WdM2+pBUAnqzCG9xfR
hRa0XacsIUY4EVBKMp7F9BUtt+3S4JkYj/3rm4EuojQ/I/DwJpef53Jbb0gJkJ4l
6G3VJffKKBXxdHwi5x+t+mZFADq1p2AFqnJsIvo1D28ebi0MPHSZaCGcd20l6ZmB
YKS1xAGZSvOFsEuicPH6xEupQ1zy/BkKKZ+cfGVZTHcZSpCL1ItdYEjfPnPJfq6Z
XOhvSmJGNng3xSk4AR/EiRd9hxsXEGlQDKXIhr1rOmJqwwUBWYUX3gIAYy4i6Zqk
52FX5FkOQtZa6gS64qK5pcHm4HTDB06A2PIh9rPYRMAbHNQncVAQGeBrnbK9BTqe
o2kz92pZ/rwl/diAgaFivL4AEM9AXziP+hJxyzZEyuTU1gKERkp4hz72LXnVPLYT
4KyLO9Hv7TuKSXg1pTwBfg/il04sCIwifJxFGgTRh/ys7G+tLdratEE9C5VdkndQ
jSq2zwp4btKhEB2oOohJ0Ltl+fIom+Zwoyqpcw9I9G7jk+I7RLWJQdIbBJefF5LG
ri7uLUC5oFO1NLTLbi4QCkB6umcDPADpoLxrBOIxNCAhqgygapKWEnXBAqgvHMNn
JwYl7cvExXydsFkECksT8eeWRBsyVzjI0UhZrDwXqZmoWgV8atpeqVidIGG8hLZn
s0wYQJ4yYPHVq+ywd0jP4gen0Ww9VmecGjB8d6cf1stg/9wHiLUBiTOjW+ABLcgF
fyK3LWfUrRap6i/vaPAM5WOjSwIB9a3Ef6fbyLFFbcs9C/7Ho9PcIDnBpyg9woRX
6oRFqQLzXA1EZb6wpTvFzQq1D9mxeUmKOH969abL9IxHrqPGURgFJ2AYIJ0fExYi
wlNv2RekNnzR+pkFSpqjpojhuveDEcRpm8a6+IVbUL7Nnm6i1gmm0YyDTpUImtgo
T4tz6ZRX3HmocnM8z74iEO6RDG7u3GJLCsVm3KDQg9Z2wIc4CoK3H45oVWgGBisX
E+Zdsr43VwEpksjvVo/x2+NhfMBZT0uyfbYJ7VOdXBODNDsclMrxoTe1sScwNqC7
5oU2l3Y3LS8Ka2BViU4oSNOPH250fKt3EBWUh589pSYHgX0g4x78CKzzCeaPDzTx
DX+a2+/FCKUbJIrGdT5J6KLxcHJWxTlPFIjcmsngjb2xJpIq8ziW8/qAn0Ys+JLR
0DBW1oNlFQky79yj6p3DbgSSc/FCrZt9gspte6YAYEfKt6B4ga3o1A73hWtTWNCZ
kQbpHRA1knYCq/gwebyfrZy07kx/J6zcXMI/sMOWhSpiHBNzQs5Bo6++98Ks2ErY
BNsBbNV7YCFS5GFlTJCEtbaDxgiQsJWsi6XzPaiWfo1ex+IM7hnbUI9cMuQFSPme
rzeL/3M0ni59fKigJcV8VgoA8ETsfKEYY/I3aPMvd7j0X/HdvUcuQx8U0Q5zITny
QtFure0weg4skEDxftHmqrRb0j4jzhpCHwErZyYXBgIhlOe5ZK3QcMQYVwaOx4yg
25WaZMrgFUrUxt4rHVev8lj4rGMRxt0CaNDmDbXY/1eS8Y44lJeETbM7OXQ3CKRv
QVjixn5Ga6suQ1/7mWvobtjNXoelt74H57xRPC9mMfqIY9AmFbo2gyicZ8Q72rBU
M1QPUVv5IJkVZKOCUlps0I81t8Uj/9ET3jcPFEgYp8MXbPt5W/BVv1ADMCQh5gn0
A8Wf2dF8p3vVe5VY4QwfRQPoNLM/7wNCplNU/cUHEs+kg5a5nEjex2/DyRVLyhGK
WVrvDa7f76NrgOkBbNzWmXSnPZySbOM4aklKDa4joTGR5+8mujFFaqm11QMhLpkh
6568I+CqD+7K/lS4O5hAb30UGYAwDpsCz3FnGvbVJ+3FMIOZFYsr2GjMYGCfvyUO
HxNCUUcK2FXoazWEEhsdnmChZcljdkS9rh01RsYDqVA81Y2yCxORWCtfbA4WkHwh
wYE4O1aRKn2Zh4LAJDGhIghr2Tu7Pcv1KUH0QqPp7ez84tyd4szw20sGpniFU3iW
gytNWHvKGZIObYFRa4YlWAr/zQOFP0wRJWoDiCTxUR6exAToujuotxD23O76+YwK
DJPuNDBPG2j3eR+Vw9Ji7rD4agTNWpsx9O1OajdwlcsrFqqk3ZUWluwZaPwhnjnh
KRO+OY/8UkmePEeJTCqbWB5Nd4xDBcYvsEvWAndmCh1u4CNWlE743Ph+WwhVOd0B
22AlaX9MAKLxpv0CgTZCgANRcCYCWA/sN8FXlYVvAqz1ph66T/wdvOLgO3il3fCD
cJKkr+QkQuyaIwCBDfo5OtTpRkMfm2orDVPHFJGYxCpHlsFqJx8GZ54rvCW0eJtH
boO4ETueosgIvbMqnaWNgrY3/BuUtklcWRJeIiU68ceW/8OY3fx2uTQevTIKWrng
CanvwbXsO3yOwHMOr3ieirRaNUp+V7DeB+j4Bj79sv0liBUG+oIOkbJBnjT480qK
izbaiokMRCjBaWc7gTinua5LTxA4T7WyzKEmsPVMTKa7IFMtK5S96xF43D6PVz1j
b52z2fU6rxecbSWJJItClkcgyIaI1wrlX6jroV0O/P3MCsdpglSRERrbYMpNoPHY
2X0Oob1bYv0QJW4nf+2W1a/5y6UIZc+pkMSCVeEUXmPDITAtC43Fp+Q9KHWxy5e/
ZWnkbTxHo2FW+jXAW7OZZ9SP6j2y8Iq+VC/v0iRWiUyDKtYKyPgxYP4y/eLDf6XT
28nY7ZvYamaLf2NqK9Q9OKoEe5pQ/pMml8h5HxPYw0WHL07vUAAJm2aKAckWxmnM
avM/O0wI/oE4C9Eh0wZcZjhuQZJLSQIOtdl6gaMbxptb6Bu1SAdCVxpsWpDmadi3
V5GJaAQhwALX1nw1CpiuKYcauTwnBL5haIzvk6SGaQdhm1JvAmTrbPWAL/pO2QZ3
4BYIUV19+KmjTNKayErThXPeT+xwMBGBgI7bHCUnvR9Z4cjdnJ2NxD+JCSD/Iuq1
qQZD19FcivYsgySaAKu1D9DXWyQfeTUiAxGkchoDttl53D5Y0Vrq6puIA1qP93OK
+/nELJJqOuYfejzE0kNENv/J3YolXxYCXB6eJeZ25Hc75E2rN2n7Z9vC3F/TA/NF
JZrhDGg2dRenSnKCex/MTQHmeC14CLEJlUGalwwvDayfiPC5ILczJc22Tk8Boave
MWg0aXcO9XU4KHBeGowuWI53hsJDCdkLvv3//hAxQSb5RKbe/5AV46zxc9imepq7
h/zAz408L43Oyytnn0Zz+GWAZH9+1sTIVqtP9xHLc1WUszAps1oepZiumYdxIKHI
0rSPRuyubsQ9YsaNAaxww+QQvicduafSmaoCIj+cCYkl+2GnICv4vo/Le0UEu61o
h3S8PR7SZ3QRVt/qJnRiW1FdkFSKcrKN30Xb/E8FfoVABQvxVFdEQv++J3szn0FF
xV+fVLBgO7p7FOFCUok8lHCIbvY7XSqiVcfjk7K6vvnIdH4/gCz/lw3GHmplyOy8
pFeXhdzSqeZGznAP/0evMAL2EuI4xofTS25U/dLDgu49O0XFcVFTjQzDvUEOOg9i
hXNMKJghKNxeVZNvrp/kTwVwC4veS9wDDOPzoixLk7q8AxwneS8D4xizX1QdSaJz
09eU89/cXrcaNQE/aXj4fS2oF0GdmJB9jcMPgvUiWToBoFA61DBcxyP2Mx22ABLr
o3Apy85/n8l9voT949Y6hlLe7coZn3I23n+Miq/DhSQRdcj3P73S56uMt55vwMYA
H/sIaRl+oq7gjrHD2kg8ekrndGUxy2ZbgZhsIzgX0mHvPzb0VfU8gRupg4u6K3XQ
d4tHb6bPEbCLJ7jhMbJhhTsgDZ+jt7ug8J4ceWoZxl7VBfMO9Tj7FIhuFVfgtp2g
XWQHYZantxmICjZ61rhLyh6gmclsYKS5BImkTZtZi0LD/Br4V+Jaa80JSe9RgxWf
F4vZsjbjWVK8k09SUiTtsoNVgFP907MUj8oiSmlMAWgR0+n721nyphWU7s/hPfWe
eQrXLIbH20jYhCLmcxL8rcTLU0AaSAdu/aJENcGJGOhF7GVA+nYMGcwmLEORTYBp
gRea/s6U9uQPu/9VnH1nU9uryM0ogLRwfCyjApf5S7hsEeOzg8kG37MF+pcP5xiE
lbAg+NQ4NpFNkY28TvkhetT+CzxQZJMLUbPsmjZESoVVnXMsWFdQPJ3WGmPAoNJ6
wEzKVT5rSTF9sBPive3owdnStEJLlb0pK7R3bMik11F50W/9kf01exGX0lEGTDWX
uA8OlV+qAngp5y9AmdSG7aefLOXxH13JYHwcBcWITiJ+9IaLVD+BOuTAxeWHyfDv
8ItFZNrm/NIvIZPSZZgNPPiYKvzkTVM7HPFTwZg+y45pBysf25ARUKgiJmDlnLAd
s9LojTJ/Yy91ZsDvZNr9r1Re9PfYS+srswNnvOUp4/NsxclQ4EB2LPlJ1I6mVVNm
Uby/Rq9B1e2xadCvToE+uUrqq1r2pU1uFBh78WnWheHciCDlccfPwBIE/+a0BrQy
5d/LY5NfwxWU4VYdOnm4wb9I4wSvZxHOGJAYWxNaTEy+WMIeUIPCC9dyfihELbUp
CEySj9SYnzs6wNVJx/gJJIrQsf++Py5aV3SMIxeQ5XZ00RXatyPN9SFDLyssuCDu
8xQ3DUj+S8byYz2nOLM0AZ8SZoDYWGXPSEfytRei6RwHBqksPMcoX90FIQtLtDSu
psOnQm/V8adRAje3RieIXzXuS8yK3Tv+sUQq/FIuHiChultDTD+FyBVb8vYR0fcB
MAqLT0tZvjs1SAXcTIuM18N0dMkmbCpgCo/bNiYWlnpNMZT35d9Fd9kqc8z4kTWI
VIAd8QkmaPR0Ur9RyxvYwuifpvE+QzFb7i74EY/uuQ1BCYspehFAwWp4wmO/iADN
z9eV0L5Z+9TFSu0Gj3Vsu9iG/z6hW6rMyWDj+EgjuVe2/czfxuaCFicOtK/r8NTJ
xseT+kwF82EdbN/RGYNdu5E0p41zCxtyc+Z3Qaery6miSs7WWr0O55JmVUjFKWlF
p6XGmouItvz/UaBZgdZFoMiAjfpk9jtugZeVOCopFuzqQ5H6puCH+gkskfZlraov
bAALOft1BLTxgaeNBvJKLbtot2RGAZmnfWysj90jHQiju60LOqHjIUxvv1PUgKSW
LOdOy3peGi0vt4EAgV8/kXl024GW+/V51vYuPCt2KHhD95c9rlgn8CqwmBhJP9dq
9rwBBNTztuEIMinEYArmy3dHJt1JSc6WY+Qc1n7gltOwgt8j+zAPa/XQ6U37Oewt
u17FsFLeDSeP8HEDUgylNldcfbvP2MrMkcoEIdoOTCiMmDqX8KNAviDaG+o9Nut9
E3FR3tJ2LXDKgUI1XU5omsHNPaQ/LFAa5a/b8CYwaVhrmkXN7aWYXRpjZ+9XzLcV
YYO4jN05+BBse7cn0Q4nTB+4+AA64ONdazTptNlvR9KukQ5eL7az+gOQPua8Am66
oBxN2ommbBwBREkk3mfDvLAUG5HCEZ5B6Ubq5YfmRun7VlM1cLB/l9gm0EPYNXus
JibCTeyj2YrDRwVV4I0ntkQ+VFXKive5O1KVtv6ZzdweLScpOG4NKj1Ay8Y6Y96I
zSshxxpM28MHJnOTQtDI2hovsB0wZXKsn/EcOUiuW0twrpSCMJI1Fc5eJxud6lZn
WpV96K8mhMATWPi+H6bTB/ht95lTh3zjhsIenFAMRsgxV9+oz7LWXKQWf3qmwpYP
nu41jafHR/nzVgkhAELCM3TZ9sk38LL+nt6SiQYDCpSac0jMwUTuxHdWSZxeN9ti
nTIlqzXCSzt5uOgTL1u74n62qlIXrDEJpmFs9n4RSSiOJ32xtO2TV9zWUH64bkwD
s4hjwZBaMLNGU9wT5GLXS0yTxrePLlM/IQYvRyxPhEU26znCFFRwI31voU5LBeii
5YPDLO9OF9jkqaGoWxvMUA45FqZXalf4baNkpEem8s0p24Wvju88uHDl38MGtyyu
l2BVcZbt64xyn5QsQIf/IwRMlkL7XKgFZ44mQSxyoecjfhdMUOoCNkWG3/bkIBwE
Wtk2ff2+tdicpuO+Xtm3PuHI/VrvNValj/GYmOjpryUe1NyF0WJwg9bbLwoKNKGz
rIDqaqDCLzEFpBFtnVbBToMqJrShHcgSbpXH9NC22IwtM+bxh3y9SyBVKBRCdYt4
P2Sx1lfeQBYh5d0T0I+xyHY9B+VlV8beR/sF8Y+9Y2VeGaISr6HsyO7WYz3LRY0f
WRDBQ1tH8zppLxU+V7DjGpEGsciYfxE4vS7lJw+jU5N7TluYsm3qPChSHSmHMYEc
tQoW3q3FZviKTKv4ftqhzgPaADnSMXBRbgyoA9EV5/BlTm39/NYfYQZDbO98hc5z
i8cMgHgao7obUIPPnJDgRbUc3awmOzFKaSVUV+Ee7CkhEkVUK4fiHDg+JuBTb5Fw
AecsZAmvUinG/ji6hbLBe1NdSty6k9D0KgU6BJS3BOYa7w8vH3tO4tKzY2nQKTEw
YpitDB2j7zOcGP1bIZMdys2JxvCjQ+Y+0mY5ZwL7Ga8w3QBcg7J3t1fspiimW1L3
K5a5CM55AgCT5xczAQFmZs387+R2Fxm8VP41KI0rXSUPVJLYfVQ/lkpT8d3E8H4e
JGEFItChrZVL0vYyKT1iWC8rdD2EE9uP4dX58zhTwhw+6zQn3RcuRZ4skicyn79t
Mi6tEj5oGHtOBugEgIFa1+w8wqiEJ+isTJWYraKr/zc0pcuXqeaDt8m4/jXuGYuL
qe1azB5PKQUYmN/5BTejExnS8x3JlFgjdGhH0acO50Pa3v3BriTLNdGjeGjvOURD
tnm60Z2L9Waey7lYCazxsQlPbOCwUjwP3b9PNlqkZbmTvrinnw/v9uRwiTLv7mVd
awBhHPyfO/k9LmisTDX3NgYewv/Y/t1sJ08jnSaW/JzDS0rC9EpB0iGW0wjZKLhE
Cz1A4nJ6AKWm7h83lwrc933LVV4+Dpm8gL89Lb3kOsDpBCxqKgo1TScrK0w2S/7k
Q2qfV4cE4hws4EnzSExeECh/N1+ay7rKMLnmJEMZsh+iM0sB2eInnhgdhOo5Stb8
+z3BhkY3Kg3jBaNERTR39dkdzm5MKqNRl23+Hph/gPP4ItdVtZU21X6Y24RRy1vM
gwr4gCdIR5jTAt0u+9RGxVD+fu8oiQ9JpGwWLnk8B1DKfkCXSnwY1ctNlAViJ3JF
ZM2pznSb3ZlbD/LZHAi+RSSSKGtOl4uPUPxwNQwOEUnm3tIDPIovXuB/LMFSZLnB
vlhgTZv5TCcSJf9pX2a4BindMS6g0BAnH1UitzSLJ3nIAhYu0Moibm2SPxvsQUtM
YyFS4okeZeMjjkyNiqgb2vKaLdwWsBe8KAPuACKCcLPbI/a/kdJefXwxSFh7X8DC
+Rls3TKjCeihGDrEsgfDIs5y1HLy3SAXdaBNtxFHVf4cs/nq/SXZkoyCt/QgNiVw
IjIR7n3eGskMCpDvUbm9WTXl94QL1ONb5JhyZMPQ7gjgB9QvsnF7G2zHbffNI+xy
DpCaI8bjY1S9jfiYxwa0v7T4WXbQZa5OaTObjPHpqPeJfbDjzKDHG7FZmKTy4T+i
tQ+cPyrZFSWgpSgmZHoL1kBHW3weWTQo8TWGnkFh2Xx+uvP2XhpigbXynU42cUqU
kgw8c2F05g9mZt7ktej9K8Z9J2QbkohdbufozRYaxEWuQusE3IOpZbcIWR2rarzE
4fPbkmHU2gW4A0iLr2AH4GFu1817ffkZk52JviHoz5XLal6utOVJuZOLy2s/ojPk
z0mj0Q8q0NAj6MmLl54r7U5U4WTwisHLmDB7eG1Fu2pcDuuEnReghpBktJUY2NQr
6HODUXmdrja06qmr/BXawRgkQ94UHGxkPvwLntyOme0EnLSHAbvCVon2VjfBuIlo
XsHf5SVr6xgLoZ1Yq8egEy+JdtXFINBbGfY/uqhRbFj7DkXDT9oCW5v9RoBvBnUc
pqRvc21UTgM2i1bS0A9sAr0u1lclGe2z+aNHKUVMfMEeWLc698JbGekNaNQiLMZQ
Gkmtuj+sF0Dw8ZJEx+RM3UcaL3lBBxtFKM0ssNbvwMaSMICDCCQrevcpz4S0bPrh
ov9lGZqupxBrqNKGicZ62WjHsqjd/Lmcx4bYGWztlx8OEl/m1FfvLXTrxw7qVnRV
pbaDCFU3G0bFOaP1Gxtmh9cncCQKVn1VeoOPxAhFaHA6lUSHmLpPX5ljaii7ay8a
u1yWYkQPGZjwYy9Tbhr253gdq6DuFW/knHBq6j4TiMzZq9utKEoW9a+rNIzCGBSU
Yi1PI1z9H8USOx1Yhmh+N6z/Y5QIrWYD/KF3GXeH+yifDLdkOPbWyyfll1H+pXZp
9ytyD+QmzIxp2HPc59CauJWc3AN+BpKYUwa/NwyJN8JpzL528fzD2mwPp2qfo0yK
5sKLx2qG45t3s/QXypWvaANbBadTGHR8W2JhRoN2HZbFUesnTB6A2XNI88tqaiHr
pz64CVdTLggWEP1NyMOpc0HJA7hnI6v6CKz7pZvcdkO0xSLmGFG/CAKOK+2Sa9UX
1+YgmToayJraaTzGNI1EuFMKFK4j+H5g+Pw7A4QmYb8tGQUbQKEI/V+cuQjurJ91
2F5uqT1ygmM9qi8g3+IVA52VhONRPx2T5eq1ZoIi1ZJIKqddF72LUChGH/y+bjJ9
SK16k00JTXCx4aFbK+IQ6UeCCX9zSwu2BpS4oq+064+Okc2BcIDq7BKOLtIPImiL
Z+FeQzANQiNNMeij5c6iYod40s3USoiY/h7dTrv4PuRs+/qmZ0imEcVf9MCHY+Wf
P0dPhg5OE7Fh2mrWFyI+vIQ6rBRluCyp/tSnulFRSOnTNsQ1wlmtfXQnNL2X6syJ
X8epiia84qkA2bJhP9AdfEM4tidG9VmmlBceqG03XMAujb99H6O9V9ffYnuQt88k
R1pqZ0XyY1pqgwPPXMH7jcqDcVhneRjbp6kueKWkbDw35wUqKkstRKBuEjoqlgrB
CnewA+0/mkF23LDZcj3RH5UzIrL+swqw8/vbsMccHbwUFBpOBMEuzAEY1eO+7VNL
KdqDX9kynLoRSZCeczCQusHJ9/c1lvGaGL8ikXWAW/Zyyr7b+MZ/mGXBjxNMedar
c3P40RzTB6fc3ZGwQEB/31X4vTqcaxosRMVvct36IIm7XoVHwcKQZQFEvmUevGOZ
MgjMzqgSJZsDn58RnaGO+KHzrbQzI/85SYVEZMsAcMwyOxaiRxAnFzoxTtDBOmBk
xKkW7s5x9IJJkbMjoPG91OYF5oNSLAKc/ASiaqvZP5LvgudAjnK/HlM8TNNX/ycD
dAuCLScUAoG+xHD7YCTT0xQLQabyt7AZtJ0oYfJOi6iS4jk+oS0iW7sYVb2rjmlC
FldWGIlEhq/8VPsiz9PPpXLz6VV9JtJvWC48ajXZ6Wij4EOfF9VsiblOaPHXIGSt
XNg7z0deGHNLo2xaAGNzsUiUvHYP4GCAjfdMoDqgQPnvNtxHy73s83ctJl7VLx9b
k2BgC+ntGOfnsCVIgc2xK8sAX5QnWRl3EujRE/CUXZCY7rtgtwOBpv5SFfMQkxjO
En6VVrR4IXPXEMKu4+6+uhQdoAEapOIUpA9do+GpjvqgjfE5BqYbJikCx091QKcB
SLMvmnaV6nLz/g+67dowmpJGHxwg68+jt7Nl/G2I62GNLTcTUGgm5Y8TkUz0tZ1t
UuyyvqIpTqpeQtK3GjU5qsMONcfMuo1ogFG4OxkLv3yIuG/Lzpn5amm6JJuaV0dT
UMpdQklNOlodlTXDmBnXwN0j/3VRXlaUzpbCIgQRUuhH1eQ1mn5HGv8G2g+fFb7f
v0j0d0BPpOYm+CdaKjOfPWo5f2cIs/RE4vwK8vjqPdxLZJeghqhUdxFusDhTxIoS
3CpQa48rEWW/M/gx8r8N+jJDcm2uMEkxnAEcIoOx12TAycvqcsJB1NLhK4riaO5t
KepfofdtXpL5eO+o9eLVKDaZLQOzn5dM+lGVSfm0gwvS29RuYf6mLF/ROsQmxgpO
ONK99IY9n9wPFIsHgeyp6/F+cldjKkwAhJf28Ow/L2NAuUtEGr+apkaUaa2erHfe
YUVLP1MWZW6GvlMZUJ2/I0JTzw8czApDuD4qjT+zDB2GrNxl5x+f7xn9R6+tA0WJ
zAGbWCZwk7kWrjZIz+H+qqls3XGWm00xoz4QU9Anfs8eHZalcmk44F+gvGjnXuQc
Tspvf4LD6VqosfSVGyrjOz7gkJ3Orojjp++ohX/cXuFoJ2zA5RXnO0stFlfZXkbY
TV6zvqxJurGjwlJA5fufZHJKADGytPRDOaZaNMbYq1cfHcv1w12V8fe2Qs+nCXkZ
n3b1z2eSFoioP08QdFeU5LpJeDszpTF9KszBR/TXFuL9xfHAjdoyJsq2VxlCU0VA
a9PXI0djqnVfTuap+029UaGrcd7kw6pz+Zw9vDli2DC8GNFta7+juAcsqMOBrySS
Tk9F0VV5ebGHg+OfU3sS97aLOuNr8qdVfP/cM7ZtOm0IpLwufamo7oWut/n/mNb8
tbSdR+CgPbhluu7JDT0JGAZaNe0qIz3AClmMNYoxH1KKEgLVKB7ikTDirpo7LU1/
y3D6tSb3QF4aEBy0nB4JDPv0zW4UnQ59u7vjobIQ37ywChCqqMCddyRVorpWNdXA
zcyJdKxzgqwdic/U5BE9HkLJBS0FIWVA4DbC0Scty2WF8gVfkFPBn0blTwokWdo1
lE2fo4+7lgRJ7cz/4f8v110AQG2Ar+cgThi4KtpdtZ7nGBHLsrRxxN7a9RvndTBg
ytkBswwWAi9E5sJZ8NjscIXpMr3jwajPLpOC57YNA918WBVT6rIkYtXDoPUuBm7o
bEZxcGdBNgwIdR5EcA3i988sOR2TucUSyYKafyHxeeBqcqq64x876vEEVzeVQumD
UDpnLnkyvOHByxt486dBcYsFyzE9xlzx32VKGupTJKtwvi86dVojHdjBXtA0QBN/
bnKt7JnxhKRxizV24yk6i8Zc7KwJ+ldf2RcGJGlWXkWARIqgPthC7gTAWB8g0emG
maGJi8pPXWv9NjagVqGc5elHKLzIhhkcDN8iHUg1zZG3+1Sv/a3CoH3vS580er7D
VwJqYq2GucnSDzaStwSAh/pQrWu4Y0MyILtZ2iQKhmhmh0V5hQv3BaQ7gITaJ0AZ
qrMUoU8crYXLkGQr32E1cQTLjLabGApQEa8qN7MKsbk8IQBmGy8mx+X0E3G/8dA8
deHXbRB8S1/6QhHguiHHmAUbNVbo69NsWznJtLMJzy7IGg0P7UbGNl8sdCoSr43O
EUHHAEL4HbQBh2tqRw/Bfw2YlnjjhglrY2RPfWOc/48v0RoCkjSLQ3nDGUCDBKL4
oUaIYRDaACjXzHw1EETGsiN99xSzzPamAG8DIAUvr2JuOWm3q0iRA0B6rAAPqssv
+V4TRsfEuC3Pb6qnxKbOFjC+tZ/jbxNM+PxgzhLKk73VeoslkhRg40edFii4/05N
9PSiNK5sBQHgmToX6+3xafAON+XavEwYVjL/LnJIOwg00lJItkLEWbtjyHfbhvQX
vLuYBewc5N5qDI8XtbRDh2MbvFB16aagH+OEr/klUJ75PubGW1FIOSNSaUEVzy2z
Ws+pr6bXZATlvZrXaEdl2c1Y5462Oi/OCAUTnEvB7uRv9lnH6TPmtVNmE273JO+G
0OkKZtGXJdgIEhLm+kSMSJGWwGNJ0nsGnhstc+NavNGazR4tX4hFMtwnS7886U7Z
n4SL2Zr7uPhWvu8gwJKMXKGTOEQtDYH0G3rJCfyfPkpx2u3w/SFuvHyLbysvRNZg
LhBay+iH/Pp29ClB89bPw9JCoClcTyabGMynTEAVpUNUDo6NmuGGM0CLzT3FKF1h
D+xbwj69UejZYVmooZ0+Wmrro0L/ag2qfCNPWMDxXO+nZS/5yELUVMRuysdmovnv
VD/fm3Y5AMrZvSmz7lKif74Au4KpEO2fA7cD3einQb1xi9kmL5iyntlsLBq70gyu
aZlI4ZkaOhS0oYJRuGz75pc+qYiSG7u/wxWitKf7dfC+Pnh0e6tybeS9ptrDD7um
rQBYaj0Js2wLhDIJCnqWKMW9Tb57lwxsymPSLIt0Afl9WZyDOJ+Pw5N0WVA0HP7N
B0d37BQis9L2npWVR/CdXLBvmhMs7bbBdfnYcqMoeCGAKL6KWfCJ8K4wR8hByvDA
uGmC8F0TXXmOYdC4tVD4RpeoDeb9n1oxd9AStsHsKmHIpUDjNIG/Sj24xIcaEgvF
lVpBOHNgrBfcPlolrvzMvISyt6nL0j0QcKH5fAIM/td85CyqVJRp+KyysQChq9WT
wWY9ZIGFQskpD8nQvWwHaL68y+wO0yW321n/n5RLBOUvmlPrteSjM3vlb/ga0SQE
H51cOVfhf8RvP73eV9Uvt9tCC+Z1bz6P+a2LeUTbGG7qItB2dt0e12iR+OTBvRnz
WHBCU1bUErHFseRkWLF/r62KOx9whwKobCQOWCtsTvSMF/rz+l9uC2uyfDgYJIRz
YIWlDoGbvR+MqXUbc+ezsxt38VPnvfLLWYm2NJ2lGvtEAEQ0ODUNbTL5USo+CQci
l4rWzz0LJQWqRXus5Zt5EOyY2fYASOIXpMLfwYSPoFB+upmptrehiyATdd3K9DhY
q9kgP4mLp5Qrsn6WdORiGplnXlZzK3mkpLb1OIk9QIhfw00vdeqjCO6epg8IW9ve
OVadi/y8X6k1wLGSYgaDrZnXRw4Uyx/uejzYUvM2PCSmLfXlymG/b+4nfqnf826T
zf4XSdxrAxV6SaXxx2bFuMbtWurpPiayMQOC6HsBmfqZ5AwKen1J1c6n9L7gRWmu
L8RURg/LtwHywCIsCIciUhfehQqMGNICUd7PdHvyg6t+KutNgWGgPlTrEH9wS3yR
DaNCtIeMTc3mzfwrMKCSrAoft/kaANew0JVGxt2NP7mMzTC/JtmJd6lTGsAaewyD
Og0bEmTalwgofip4dlPWp+ify0j8K7wu3DENGvxpNAo66DOowmGfi9vorUYHv2QV
b/4pbfnSLbUheRYn2u+L5lbPhtfo7DLq9lnghBUFFR609FmyTMfi0/o2b1iZGY5v
LocsvmTs3kFrfs3obx4hqv17nXTYDU/7gQ+pLSbAYPaTD1qjTsOAH65NCha3PADz
djGild3kRCll7cxfEl7F9iDBEYQ67HsY4yHCnTVnSUZebEYsnW4uRWKALOB8ZYD3
H/71bhPMQGJf29AWzhAvqv1e7rJAnCEKSrOCY6PhqhagqZ+URhui1Yjh/0jEP9tL
JAh9HEFrIlngSe6VzhFOl8fnK/5VPM7UxIBGU3IzrS2RVdNTPPlyPqUBwk6sawqz
KyCKEZWT+ge3K39Fr30afJrk52T+B75HMuZwLRmsmqVxQ6VyVNcMCE3EHTzwLvq9
xoRHZexFaFM4fhPUEL6I35j8m0l1BaOQyXSM0JPpKyBDqxUzG1aEB5pZgYPD+1ey
jIYbPZa4WU3tlqRZA7JGn+reXZsimTBQtI7oz35ltxSS7ialwKNMuyFloPlW/hxf
ec54LNK3AJpPdib2gLmuwgRA+LkEsJ7RvQWie7G1xsWetfunDP+rcYaYYqh/hqYO
fyjGJTOKuNeflc9h1pLKX8ayU96D9artYjLUSnEy9kZufBBDoUVwYMccXHxXpAiY
ywUH1VjI3FhJ0oJ9oWbiJd+obTVK0tfo1cscXZ27j1RJmquLe2m/uGwChwSYkFsT
WT8UmU64ht1W1HIFIAcQETEVGDM93KvzKvXajf/N31bgLuLvQYghsWo2mgp8Zat+
ZDgzQDeV8BStvkH8sCY8QBggeMlJrcI4BrHGkr5AGCdXpI9RlQqNNLXu9hbdz0te
8s157FsgV07kU+6mACFyOggxp9DORk8Gf+YK9wakPU7la1kTSdlIDmm3/o03cpnd
ClMonqZUoPdU3KAI+uV3ruC0azaqbDliYqVm7DfI5adbBiTvE35ypxJKoPr8RnnA
2kL7mf5QnEcVUAA9c0gs/5p11NouSioTrAOT07wK+emUWiX+JnZAB34w39LpdVuM
rLrG87L0/FunF72jE9FH/f3FQDKtN/1Cb7B7orhydRKjxGcLL0PWgWOL8e8pMUsS
WMnXX6f9VxbtPB0dGKVfxBOO9Oc43U3HPjM4WGeozEm27r+FJ1IDFi/A9NeoTHEs
`protect end_protected