`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8224 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMWORzZC7bo0toZS2Zods6Xs
yljw+BvqICQb54hGe2JGpCy7VfzPucQWBxxbAs+GRaiWI23+mMUGX6Bna1gCsp/i
YwjG0CfaztroJPi2R4MS315W3uWgAfx5FCQ0Gddu+p9zCrr/KMA8CJY+DeNFZrX/
b/1lo3CB6Son4R9udQGHXzWa2OBFTHvhOOdGHC5zCLjYATguyuptxKvNDnSqzN2I
YnP4aI0qah0gP4cOuxjCMIJTYIqov+ALK0g3ODo5AqvvTQfWlTCfiWa1G2EWRC/a
meaT7IwzUzsep+Esbyl5qFjOIEJ1gEfH88OdIVzqpvK77viejLE0IbM4qBMp3Yef
nSFdbXaYF1IAQGqIvs7Cs0cq/lqGja5p4i758uQ2jQOp9gAYoQ/5vZf4N1fzC9P+
GT78MMBwTMJZtbY3OklKfrVfx+LRukh/QWgIv6XsISx2mHEuEF6NUi3rzQpZXfNP
uNxOXmyE96dwUsEMUfIBXDyIEM8m2ZeCfl0VTtnpulP7+Ay8YAcloTd+0Dk2lYY7
VLYqS9hdFW5aK8XLDW2JU7QIG+YdwVtPLkPeX1fr53mJAizc/DSIlQfEmhmkashV
eUBoH4ahuZSfLtWrjNNRN3714wELr9GQ2Bvg3STvb9gp2VQKMlYGcfK/EvTvp4T4
cDUJXiQZfJjZgosLYWpljQP5KlruHDoetOK01/OFnHT/1BaPfdbIq1GNy0h0CaT2
V0IelQhC8GXXYgOmKYGzfLYNViwINpUkeEqEv0y5Xx6bauwC9UgUdHcWn0n83BsC
kSbLgS4utNwTpS0twxpEFj7LE0acCP4zkXokmMLU5mUMq0jtp3TcML6Em9tbQE4J
fcuD9bvjYd3k7l7+vKHtUhjNPwEiIYSeJPjHsJLCnfVVINBegErlNh0Eybmvq49g
fOIuWWnKddCG2TkEmWpVl8YD2acCOeaTmacE2N4oWL2Ok5gcgxlDW0Qfj3N6/UUg
999BJRaCitiPk/p4uOnenn4m+XeqmnjG2Xp72NWFupN6fBSCPKpwpJNY1dwFbctL
GEkGP+quTWqlEwN4iXbXUfa5obZuwvhju9+Miye60Ll2QG/9ZIYuShcogonKkNRm
CLE3vdCjtAgeZqNSUA8gHrmhIQX4C5H9Zw+zfQ7d1HiR6xsliWZ12xTm/hx35mfn
yQv2UhhCruqa3DesZirCKPmPyQSp93gL9nhzsYJmAfyIAY4rOk0gLng/U4/twpjL
qx2tvLXd1KcVHmpzRXsgZeIeRZyWARikMb8bBqEtmPkY5tzSD301sit+5rWE/4/k
YHu3E7SfhkDPEVlGJ1w8Ab19Q/4beweQFYRDRVsGg3tPptVFTT0saOJHrtyzAo2O
mKg6nhJrRXaxNubbad2xaPp4vZVRaVWv/D+YltWb5JBS2SKiECrcM/fzAPf0aX9J
2aIXXi9rnjxUd5OOaKwwswpxTDVbR8bMfTjd5+rnT7c2G/RiiXlCjbTGpZbPWQ8p
6X2utQwi31YZ2LbgxrwycVFQ6Yjsnuwi6S316KvFHXfiALxey4GjWqlUDe7Ou+BW
augLn21DYzBVkmrJWKqb/RhorFaF8fhCOZ0cWIFie6b+FLc30b1PLz4ZV3Wd3LPY
fFwOOD6A4pw1Gtee7gnGNuzAFm9f1GULFQeP60vq/3olyQnujBGQUJYp7Kaw65N6
/0MHiJ42zh/oyEztFic1QoDertBlHIy0maIzTrwWV6rEHjIwwtUsV9HyMZUap3Og
Df2ZKYM2wgn4uD0jRNcXmitbvvpMJei+9MaYA8VkWrJo0pQQWBsjNhn3l2SGzRdf
B43P1TFY8VkOnvNQ4Vp8g5DKQ7dKODhN6VEl8RVxTkziWOnLguCDQvVA6O6NpI0N
o5R9xi1he8x+0M5nJe7bOamFjGdfA3W/TnYipqo9GWvcD7+DR52C2dfB/qO+Qa3V
6Vy4PZRKJV6Em0otxtj4bqZ/5UCDoiJwhA/xZSQI+04c61y6zsOJdemdwGUxgc6O
XdQT+KMEzXmjNrkrGZM4HXKV4kIlbkEkdYV8zomp6zWKgg9A/EP1nUv8YRJ7hpIg
XTbqbKDdNI+XKupn8WgTqBzT0eDLzGTccuhYT2wiu/LJcNq335ApkqWezhfGC62m
2pU/pV7L0DIO5fKU4WBG42o2fOvVv+NovH6z8DjfIMzp56hCwlGCP4APg2YM6N0l
VDYwHBb/xH+nipwgG74TPzXkYKbdolhfwXLMXI432dwrVF+ictuINCQZTL9WPXgX
s4CdNRdso/9en50jHYQtDNA3Yv1WCV86ODdxMvSF4DbbK0xX+UBFzZOX2OTF6dm5
1iR8VpdRVzWmaIMSkELfv9yWwwiUzegPB8IGiHKT5LT3Z2Y0fdgJU7rCp1pQSxA2
wokp3hPebtSEfuOAefv4UJW8SxaVrhvuMRcBSRuFj31iK1ulY9EgSwiKauZrp3+t
xP1X5nQ+3tQdBVSbVmlIr5UvWOzvM1sm7HRqjBYUQ4X/aOEvbB1V9OqjvXxO84IK
1DbsURuHmopDXnfMp43HThGBuk257NsMkRgwJS0u8CqpApqyHmPTBixATO7917Ow
FfyA4NWzmqchYMonGrQhymEe0jj/J/wXkzLdnuybSA9v4Wnl9GRErRE4DIDI+pij
fs4XJGpkzo2JQlcE2u568/ZITXbyilrS1qhaYjQVYOJYm1fj2Q3jk8HBbsIy8gOW
L8FVNXvICbMI8151ysdVtKRQAtedqWuG1Z09u95CfSIrZntFcJGgwMDbbB3sjBGV
Xg9eVk7ZXdyKYmui3CFSxzssG9Ls4vQK+3QAeEh5NEZa27sfULnLzMlLbdQB8qlP
JlyTafhrA4z1XLOVWLyOyu1HK49kJIaeYIoAQoLEAr01lzt6+1ye1P1VWXw7xlhW
naYas2e8jZLtXCgEoUdgD8H7RZuIGRsArafID9PWhkGnhJhPLumrY4hJTQjomaYC
e3iSRWLCzwdYqmfdZGkroQMN6HttWhRaGejgOauzCZDciHkghKKAl27bn74lXQGl
djjVKVL3Ad46Lzav5hComM6iZosPqBgUYgg4Gt000wLunD7ovTevZ5wteTMEEB/4
s0nR5EDzKy4zew/QIr9KmhDHn23MwLcB2aRuyzRxgjP1GqddJutnIZsqydkSz1oH
CEVC+tdP7FtD3My3VhKScOgkuK9Fv5rTCCbWm9jZPB1sefG2IZYQk2bVf6JBDi+X
Bqvmk7a4EWqNt+Ac4GnTPyhrEQm3tKLWuhfnrITE2vYSl/0RdVQCBCEOlP7xDKXi
zkcMiQ5d6qElMgjFqqV2dopFxU1YafQxCJNXtfeQpsUxVUvOLQa3ZH7/XgKD9mKi
kSgksh3hF4BxkU9gO3tig+o6VL/zmhItc7bxYDUbmQoWcUd67lrDWUK/AY3hVS1+
OH9pPkHpNx0qr2aoXMCvI4Sf2ibEyPb7l1+n9Pcb9iYraJoRMrQkkiq11FWeVk7K
ww3nJAvDj3qI2+CukuNod3/PUVVEa62ZkViP0hrBrGoUkiO67bLTlaiBiPHCrlgy
kCqbEk3p1n/TqHLT11UBwUrqOt4u/wI3o7TDEsbH+fyuPSOx8x1/JRcHaUzEBma0
vC+78UySAhMtW4jDq97g1u/UPil5IIANpBFo99v7VKM2Gs5egnz1qF/SIwsEBll8
2+QXKjdlp02UAfh4UdcwrUhvsWfH0dG0WkUHawBJUqzql48Wd3OoMbyjnOcTCRPb
URb8+NqQbrBkZnrD5Wot7DDwdL7HwCkvU/v6y7rtgc/pSGDLN3kbGi0Uii2DpoYa
x2SjepvL4qwyPzhmq1ul3pzRvy0o3BtPKHSdx7ThC/N+ZGxT7h5E+KfK1niDrbIb
3cwc12yviEBRwpGOEVwsyj1bOGgwp1ljmij2MyPz95XkkVdMYCdhBUxFJ/r7QUe4
t67K1Epgze7e4utMXaykPDRz69mL9HemuPXDe2YdWvr3rrwhOcxsjIPCNRIF1Ee9
sjOOx8EHQwqK5HY/uZ2Xc0XsUNGn4ozBgnXMNyltvk0PlMPrOnS20POqbvRwcG+H
0J4xu6KfMD8Ni0fyE1dG4cAypTwMzbGcBtZ60QCxJqUS+tOjZ3n6C6RKRcHgPaMU
eo6EvIBQiFanMXKATvsiLLlO43CbqvRPzVDfveExWCMQ6Bh/PKLrg4/76ugFaG/o
UQEc5yeo5W9pDUpq3zUqK7QShX3lxx/SRfyIQqFq7ehbqdUYyqcqtKLoCj2a01+5
jFGkR+APdohQqod/Fcanxor93dSpiUWl2cQ6P33dn3VYvNyMr5QEavD3dI8+R65y
+kLJs5m5XIFos+y64hqR1T8b2+Pn4SOEaPnmE2Yi9t2ER2WYKPn4gRvS40uL776q
qrNkc7jz6Axk2LsISl5A/CSWSDzVLnqHu0zzltLo84f9E4bRcmRUI2KnS5+L2Q04
ZT8kQyEcZsBFVNeLXadjaECtlNeEJWAmmNOtK78fVE6D1rIjwadStGHwadx/s3em
pH7pp2BkbVaa5Uvph8iLyTjuBbDH2D4JW+2Hb6O0qkHr1rY3XIdJtWkRew3uFcAD
l7nLw2U/4rjloiKNRNZ+pFF0XQ7AQ1PfERjem3kSkFviCj+32polfkpKDnsIrQlI
cVP4aYewEguPGZGpQHs6lKWPVTMXy4B7wbQyRtWHZb9puH7GpdYHn/8hYs+ZLKn0
BpsYe942OghqRhYkOHNkwk6OH8lp7WmeLqataY6tZoHCAdQOgxWRsKRLxrXjHVKU
xH6zO3NXDbo92+8EuvLSIc9q+MTAa+LT5rMcMDvaQb1eIWN2Zt47oMStJS3mDifp
0rG+3Cep82Q5FNN0gdkp+jBpD6NXtK3vTl9Z2BHXJdpc1Amo+pYMrfVujqoxYsBo
r19hVEK4X7a4jvpJpbWfQvPPDwAc6GwsKD+yfDs/dzDLzJtGVTOxYxHNNiOi+bQG
q1DfIr3YCGIj7QaC+OmMf3EbWrx0BEYwQRnfm+XIXOWh5HHBELMdsnejjletXH2L
9QITDE9xwd5DItX0zUFwKsM2VZQREwiWestpN/5lMvddA3zMB6w7UG9DPAj1hJ5n
h9FdI8Tk9A2pf8cbAci1559mvPCm0L8pqjevioHXt9mUoRTRx0lWQ+OHF3nIJ5Xf
rHFek55kdpbw1Yt2TbguDyuFyBlldRpPhtJYlNppOpcXzyE4FZbGr2wxzVniJRfI
LcJJwl7YqBdh+wdkspoCoxpLY5vMHPmQ6BATjcWLE77hO/7XBHF//QkwwbnuSw/m
Bqbi0CRoWxpusf8/zHQX0nmTg9vVOsvfK37TRCNaHu03bnLAbRlaAqS7TKeG4vkf
q2sJ0Df/bvpBt5t1OJeubRrPV6n+0gjvB0nNzb9MbVusJN0zXPExrptvyCo7bBFv
QcFGAGAMqLOWHCfdE+HVZJIyGGGIQnKtaLcUTmqlm693UlcpGa1O/HV46SD1yj11
9dVW+mw8EvcjP4VvIlB3sIqx4Scq17Qqd7IbSqP27L1DYJYVfUoD/p1fU9E57Pvr
EBHxYASN1akU8kW4lFluocaYvHqnEQkTI3+aQ8n/VEioraiUJgVjYaMh0niKak0j
OkgQX+MoUwauhUWV+vgZaSkDU/YYC9mrhM4KYCZWUH3QWAWsfO9N78w8a96Cwi/q
dMKTK9CSbBtAxYnmh+MFVjhJEOaTHbudDcYG4jmF8bHjo0KbnMt/NwQUHCMa6Dsy
4u5jryE7o7J98k+QKUFSqa0jAEekGKPpe4jEASIcLJS/kuU6OFSzGDgZRUhVsTAJ
X9m07twYlwEcf8BeNlNbYg3j1kjsiBhIG8q000kDFF2yVzFeI18hhBp7Q+28NNyo
gbbQNoM2zITADRI2+PCn/GaybJVnj1cA1QvP5zbRwIv38386ZuSdnObGgKVBG6jd
ceMh0fFCru0G6/walyIpV+Tz7WyhWWA8rDNcACH+AO6ANh12fL0jFb0U7me1xaym
J52ejjQ2dDTHFTjOcpO7hg8gpSan2gxGVw/DqjO3WAcw8MDL2K6yt0OZ4ppeY7F7
Y1NgZz3bmY5jfHACpEk4+WYfP+WKlD3WFvOEh2OR+YstFI6UBD4406tmw0w/5udA
20PWPe0lG7/8bvRcoPTOxZdGWxPtb7+HQa8FBXDYTA0wnP7/hO+ePINKUqUWMoXb
MvedYq/TtaJtssnjqlDgX3J5h7786IgvlNIKufmyJvmlHcdxFAZvjUjY1CbeUNoE
DkQUOhGdzfTEnCsgiIGMIzFhcsBLmhlqyctWVCvbwJuYC4599waDksOSG5E1Nv+o
eNX8jbkboM5wJ9502zHveVVUob67Val414ItTmBbragCrSBqabz/LdbyagqBaukK
lY5yRGilPw/WjWSYpRCmlr6XQwSXpHe00ljtOCNhFn1tSftqHz3C9RK840Zq9cnG
86HsX5nqlH+1HgNLk+lavvn3LgN7+5ICZc4qXf65dhI17Lxol4QMv3oCFSGOrDj1
5yo9GFXKNXOoSBLJyFgmopAJX3mOcGNSKaBvjW7V4f6B71VcQIdM1kXKgBLthTf7
57qIaI8iR2ZU38HJxTQ+OdUNCq0bLNxGX3QcLzGLLye19Rex7ewLb1rq+lIVUK8h
BtQ3yvCSSrBXr/mSsDJOf7u3edrKxNTJmfJUCSEU7KS5lI8XzbskdMIc+y7yw9Is
ISygXGE166dPzz1KM6IDhLPzT6zZkOYwKRqdO+hgbuGOhvqUSvlHddv6ihW3LgO1
mbit22CQLjBpWqE+k7O9xCyyfsBspsLjkaZ/Ryulm6vMShKb99tYc8/wFhcAxfhE
leMXMaJ1YbMInJp+kq2sSNwucp2leFsYkG187KzSvb5QCLLSupDzXjCX/THWikf6
EITb2q7VzOls3I50ISRMaWc8XCvUshgmr+EVvf/nybelRKBM0C+HqBk6x+GG+yhX
kzTlEpUEG5LWjiFfHyVFhJgcUJ0UzZ8amwxp5rxR9dpDqVaMYuD8IAkzgzDNs41j
NUcmlgVbMX/7Tr0BbzoMU/yuBUWFjJfm3JxbGNteHFjS2Y97X4MnDZkh3hdIu3SZ
e/zjPpsZ3pClf8YlsyE2GmkaNLkGYkfBAcnpuq/O1dARy6XJvcZJFopQtXDHiIPF
KX0HspuEyiFn0gCMT82PxQl/B8DUBD22VE/j9A8iBSMga+GnWKD+Un1kMYpdMDGL
8HxUvtsQTr17HpuH0G9eCPUfErW+MiaQeg8KCiVu3Y/jlCXmiXIDoD33iWyWz/RO
L0mh4RYqArKzLpfAbBWYAVEzR3KP3vpV12pc4+Jhnqc3Ch41tU2lTx/jcV2dSKWD
yKImKPJYkHhrvc5IQjdCFAiuVbCKJqFK3Z4mUiPBD9qJ+xYQdJur+JcLwtDnwnKk
RiNFVHU7XsrszW5i0fyKI/53Hz+DdYN542A7PKKMMMekKZkLN+maMHK6bHZ9rJFi
1M3Nf1MwBeeUKUwilMTWX8Rb4Eq60MUsvU/bSPqDyN0gwkvinK3vyesKzFSUSWcO
omimaoJSMsvPpHO+KxQWEDDv5xgfZZVCZ/cAfS7u7lm3o+k/ANX9NoAL1cco/9uI
nuTsdI2Y6AzDa/rzJ+t8yVW/NdFdNWxHGcBa3FOageXedq05rlnpZJivC3f3Lkse
0hEKlebOIo1Mz/BMI3b2ZcYluCDtPLM0kvywLIHdqxGM/F6cJpV0r7OXtMSx43Dm
iEq1S2qBBM5AOdebmpQAEsklqXJuRs2rCXS22WsMKsdu/xiuUYWOjO94umjkJJK9
fsNxrXU8uDg/fEXBDPbcxian1g1QRwtCjyXrzcl4rx9HAXtgAQ4W94QPoR5OCwpo
mUZkSPRCS5/c8ml6Jk2dZiiV1CSRzcccH850Pr0d/mv7nbHKpzBvV6Shpxdb65xs
EecaPrzcVWQZ+fVr6LaVcud7L2w/pl8u3Z/MUbzX+BMdaqJGptJMRIFr+AWbLtPg
e2LX06tW/Oq5ksUnDf/rv0JX6D1Drm9YxOvWF1Ng45V/9rCdcwhEh090CUFlodVH
y2p/IqPKt22ewszvzYys8r5I/XKBeWZ5iklqY7UsRTc1xUzvaT9g+6eZmAr+L6JS
/VT6PsUX3f8t0krHdC1suf7NdkS2xyqME3ayJdUW+qu6k2qOS3klw2A/dmHKKNFb
0Ep7gfqPN25DD75ZlZ949JX4m9eO6rAVyW4HJ2Z+GJ49l3amN6a5zkynShRx2dXW
Ne2jSolX+q4zwkapMKCC5oIW3AMtJP8oRfX1YEteUZZCb05h5tfIXjy9Lqm4N+43
1bynpgjV2juIqIpZxJ5Mr7uPiBXKh2e8zOh64w3rXfehFmpX6lCC4PTUCZdR1/6y
j2G262m0bBMjM1XfOffs+iLaZY1Ntx8EDxiAmlzzzceFjzBvds3CBpMK1fapU34d
PeLb0771sG+hXWODAxeWXy30B1YV5gI3WrWt8e7sTEaeTXnOW9WLwaJ9XzdkyO99
HDquaezU5/8FJwZgASw5z2ut23yujfTUnaWHP6m1gSpaEUE3l6RpmRSpYJb0aSm9
MBautK+xB/cg6pgXyqrc6W/7ta59Lntw5hg0zexDhn5ExekxUk5JVaJqNyt/C/Ni
yu2ycZPV0sbBfzlOsWHMdH+9doONYzwBOFlBqBAk/JNMuVdSHBdTnnCf0P9wMPGD
UvZNjbNSJ9kDAjP38JppQ/ivadYD1CXTTuHoKEBKz9u7MiEI59xNThQZ2A9lcrHG
vN0JH1Ch7IT1+KqaCBMCYdwiOICncjOaf+ldSXCT6saJSeuuvPo/7XntQWDBYHPl
U9JNr34OEDcsfRH2buHuxBq90YTZ6K0x2cAXUStrLTMVvRYTszlsyp2l39pxt4qM
VP8iJXgpUBwi7OHdIEeJWZrMRj8qmbTds0Tj4+3ynFN9mcMxYDHlqcpOiGFKESoF
JDu4q65eiLfcocfeh+wHUS5aEh8Oid3zCqDIGDVQt67exE1hYJ+L1WTMcaygjZbX
S6tyO178Lg7eYwKGlABOb+qRWenCSBus9+yJgufvg5mTb39bpE1go+U2PmgAy6p6
smFbj8WCVHGM1nzGbBIUwsHi99P4Ow5Z5PA+cED3jZ7mhpcMN0SLcSgE1veqkkRs
Q8nOGuVi8u88xvSRr8fiu0dqwaipEFSKJhk1H8432VZzHC8mSvFnYxLCRd7mN2Wx
YG2zFjWiwM6PxKRohHPHqjcgLj2kvkXJ7U9RIqqXoUJLRWu9rwDDy90kOu6qF85E
Q9wbnlaa8+oI+5ZyxcqrfswA5mEbS5F/ojBPCU2W4fvOFuXCZY6bn+K1oJmrf4WZ
NDE4it6IGmNK4nIC2o6i5v/Gy08IkD99GDEsgqdR1TdEeJMNmeP/qBFMzbWzyY89
Ranp0d8uE4ouaAArTA0tyemRKLvtAKayWhT1Sxq2bn4UGV7Ik5TuiGOBKLaIyqz2
Sj12P9W48yjo2zw7YYIYtrbVmzmGAysMvy6cOrA9N7mcfXv9Yv06zS7pQy5nYwlW
S7TS8e3dHsMdXp9SlVd8paLIgYeQZCLKMEW/x9C1IKCTYFb791BUFa4SbD7yf3J8
Ao+mu+VOQw7n0vvloGqhB4bJI3FwxO9qJ2Y5QDYVy9OHZRqh0VE69DdAPGyYDt4C
aUOhDFbExfWsbqllyaXdX6K1xIL3Rw+lHcneeNBKRwmF4XVtz8NIkno2hzA18bTv
bzHRRAP+qSVspJa9j0po6TFzvASwTVCl5Ixjy98G+RG+N45TX+bu+cmATr0BCOdQ
PzCiZ+24sHTXRZE/DZZjauR+XKZva8iT+KIE+fmKLglExXO66xLU+/UpXpttNeEb
TxN4psVnR9DsM4XQp7FqOc4mvbWhx53oeRDQfYjjMKCq/Is8eIz1UI6OEHJP63G+
VIIxp/B8cGJig2ob50LjTHh1ZfRJGFZmOaJ2XCAim7oSLi43wS7Ec3WojYhlfq2C
/oznxdfNbjjMcl8enIMMcvhvGhbVQoAOnoRhlrxJdnvYPPj3tRH75IM5Ut8/3Vhs
UFY1QGCxXA8L3MmkB2+FLscwz4vKmznY3YmzzI5QxVxuv2o+TPyjBZRKL6yDdpzd
sVaHDGAwPmS2Qnvc0YhSfJ6JK6/PGRoKEPhzEDm7A9gDXwEr7SwXgQ/NjLIwOMm2
pXQhvRpnCuMNsuqjmIGPO8A0C91m1PpuJLOjVIQIeCQ2g1ldIdW0bcGdPMv3Vj/p
sNKuC1qwcRbLA0PCsBd1+EXKUzeGccnQch66F7MNyyS0FhcZMRgLXFSvzsOqn9kA
wh5PhbHAUHrIZlVRGU+sEAIEZ7aBwMCd/VjjW3lVyQyAzRVxp0XcU22c9C8jQ9TZ
JI9wasIy/sxtEtRWmNr0OfLWSMKLGwPyGlW0EDj2ZvPIQW6DL6WN32tOWBMe4ujZ
hvxSXpKjj1HwlqNbWgH4k8zVWG9v4gPUvfIJwUqB2hTEVBp8JMZytrCpxLMHnNh5
VYRawrbz+FexKe602gH07GEa/4arDboy3rRk5m7MHdJxJQGX7KzVK42PuJNLOtKN
mdWHWQ0LHuhWWser9EU7sV662wYn2QDog+dJyvcuP17VcZuRfWAgfzFOUQwhRwCr
i9vMwhTB8LnHsFYirpssEGt8VYlWsn7Y8DhlOOKZzpQ5C1gucb9A0ThDTk0Dh2zv
yB3AwVd+R25wvuw+BCzzVdZSspNONMDkzdJB1uEg0+eZ/vAXKz6KZipRyf+HUc7a
4DlnhmYbvzB1G0FPvyo0e2x0ZPbl3mQqRqOMzvJf/H2IIRWd8EzlCTl9KYVExda+
SF2TJqFjUewKiaDFPn8mrDUPn2Lh+MAq11srJChHfP1MgAXJoyDXqN8tcZE8H3ZJ
1BZJ0EREifFiqJx76mDUcw==
`protect end_protected