`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36768 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
iOS4T16637ogvUHHJHvO1N3lw5FMCE6mM7RNPK82KtiaR8Jhf6WXt4niI8BDJhkn
tWXudyCGUZRUGhvMBGy+xykhbkSKP1FSO+KaUcr+OdaF7dvHbCq69ouOaCSxEOm1
iDU83nYRuKl3WlqUTtSEwjCrBHm+PPGv3mddK3cdy5c7oSUlGK/XvyY2ymGl4G9r
7w0UcE5CTX/ZkaTT0ezunKdWu488Bw5PO4imTk/vPrrJY63RCk0YE75I4S8lhpHL
hladNFdd1cr5o1Qftqn9u8dR+vb+ulvQFhy8auZpwyhswifimDNElkc78ggfq5L1
u4rinSym0IMdpiff+nWk6knAekMUjVGHHnUGm7YtV4doWul+fbz5uIDJFVJGGHDK
Sr6XJzG4Ox+vhp2ECp0AFPkQ1R7iim21rFgPoVRV3BtBT6GX/8UJ6MN/d5WlkExe
Omm6Cj78Y5Osr9b0BsLwKyf0EZTqMmHGi+z+l8pbRzxV/LmvibwksH/IrN/PjTnv
/WGT2CtBv9STWyyMzpvpKWnRK6RCPPoMG952CibGeFr2CQUHmwjQfunmKjbDIOWT
3KinUuob3BG1+aZuI6gdvApIWw9rH9ts9VG3XZuwF5p37QY5JEsp9kBS+7oM2EZ1
P+P+R6yQ1foXh0i50hLcYFq7ngHngJ5+OXZ/wVIUwb/piyK1BvXkT5R8FWlaCG/Y
x9/T92CcepD1V3rZM96nLpNSD5ubIaKnjqCI/cvlPfbCehclDuK6IYIEEf7c+bJ4
x7i+a3K+rUM/+Vzc61R40iZRYhwIIFG8DJrw9pu3l/pRfTJv6quSZsIQWQf1w1mF
xdWckHihYR1pMBtzAscB2OD7CpwygxgVIWk3eMOYTZsue9GauvUPNL050KlxF12F
PI57OKN7YATgroGPIB0Im7Ilz+AQD+QiX3ywYb+FgERPBcvUeOPdG+fSOOqaaWmb
9Ai1ThX7P5Yw48rCN3FZ9Me1Py8FHruGzwMT3EZ6RDUxBl5sugqlbMpo4FTMC/ra
bjZvVnrnjUyJR+6mu9LRIlrLJNbcQkM/f/vYaZyP5DTcQF2BVvyHxpoH6+iZNRnk
NGJQe4IAJfCvkpsFaIfb5bUrZaz4XLM0O59fsbA6Ftn/rpi/hcfwiT0uW4Ea27TF
cv2hTjoaDmYZ6gRbCmrA22P5rprRlx0nkKOtuuin/XXai5W8/3CMQ/mUcHI8bG0d
Y1xqoYh873+e9eFHQ8J+wi26gxYhSlQpvtm1+cYkreBUYOOW3iedDkmfvtuHDIdM
oq8KHLmpvxa6DrFW2MFadnsnNSerobeAhHOM2Ozy8M0FNwV7VbwVgbOmp1NQIyY2
yh6hf8ytMM30G95rAqa+fhl4CANbpHMRljPVx7Jkwxw38fUQp5BttPD2263iHOJT
9ZaBqlsBMyZveq8E6LRV8Gzkg9g5VxTr83ggV7IJ0cKT5qO8TdlMd+kWTOaj7wqO
CYB4u/hHn2EihgCw08wluRC0ICIp4CDWwKBGpMMj8hPymXMdSsxX2FtyWxt5hE7Z
z2CYwqRU4XxMt2aArRJfB6bvORo0YfhmdOggjsBTCgkQG8i3J0Q/PAhIzd8UQsB0
P9qMlqrNZICc/bYDwh7NjI6SDWVt6GAau4uVld5wqz/lFzHBqWNaUO+o1VAe3SY6
hDhG7lDTpAKWLPRiPIHxRnCT2yNRDevZkq1lmdYnXk2IVL6KFnzG7/imfvDPguhd
Z5ppZdMtKhF+gMlYbzaja91zyu/uGZ+84onmZrS8UgsVyj7EGkpbUXao7IWnIQ1S
3eDJCTTn+DkuNWcYPa98vpwoDx8F+k4MxRns5LkPo9f4de7p/1DePoyg0Jq4d/7t
Wu0St1eABIFryOizD8F/3InhdmDef8yxW5ZYb//ad5Z6QZYLKa08q+pimGhkykNg
sKSiA1EtfNmTJvjzE/+c2A2QpZ7ej3yqZ3+qFLRvCtPip02IJZqvLHc4iP88tVQ+
m2H7ix2d3zQYHvYErcaW6cmk9MnjF5+JV5pcjJnU1hQrpLPH7efu4AHHl0iWloG1
K23rIcijEx8R+YKudVT5O9If2VGRb7DluxRJV0s293aEiwkIWEqj/EHumgMLk8H2
4DjDnH3ugAeAHA6h1lwYzma9ZFt4X44Ye21BpbKKIsRHUXM2Ka+kk5Na7zxhMQg8
2SSRXsKadJiCv9NtLgA6qVWyHkaPeGI1RUIbTvDKlvxLoFrBkuEjZsqGlZBEMnKI
lo01SSvQQXUuYPzKS6y7g5q2N/BeJrPUO3x4Buqydzzqcd8KAu9Kp3JxDERYCbQW
NHnlVvxL7/EygKOP+Hlrhjp52N22cK6yuxScNeX6QMqdWEWhccP6HhaGRRAwepO8
5RFlEiXxad5bYuj9Jqvyj2cO1hJ2/FInQi30Oq+MIDQI7cx+5UEdJ+si7foy+PcI
EQ8rEeWedaiaRhE+WMr/heQEVb99fmMBsYLUy+Ov6C6TMuSlIbmJFOVeF7GAFeDp
H38rfpOk4la6zPPh8wQ1rj3Nl4cGvVCSsp1Ksp+AVdqT/k9tn2Rt+eKbyeFMi9IL
zii6kakRBHFkiEzBHOble90D7pEJxrhENPEc+dOdT4cPg8ItzVlU5qf7NMpdGu4Q
ik7TyxAc/geGmtOqPsHYZeKUlauMr7rsFzn7AvDdMWgNbucWWz9B9jDO1cA8nZ8Y
90G5BTF9t3wABy9qaZ59dDCUmIytTpg5y6yILjIU0Ia4GOvICfoFYx+9xY7YLlQ4
LuD8JA3QYZLgkKgwnq32v0GeUR6xT8BP7yEDaWVTQkb/ixQ1ryYkVV5+cu/TZS9z
6UE8QVmhxQG0iu8LyeiVuOr84z2KP4gE6pi2meo01oOT3wPK+6EbEu6TS3cxv4ZJ
muiNUiDxU9OK4Mquo0xU7nb+v6/Ldo1Rfg/MGlW3gix7u99AyaA5mAuaY3gCEdw0
0q8lBPH+LP730SyXcb8ru/67oATN/dZ/Ex3ae0PUvN5uq1/l9Pk7f3S3swXgaTlo
bC1d7Sx4bskD8M8SZDEXjLv4fa3NfGNsvydE4Er4rXGGDqIe1FLXfUgqgmbpCccV
fekQ014itgt1FCt/Pu4h7WiEPCZiuFj6R9mFqDrhElDDxSLnxaDUT/CKO8AAsilm
DiaZILwSuDtzlAP5T08xXHQGvapq+3E5x6uTvEDrc9MUDQ6AH7qaKjec5dTogxNh
k6m80McvZrvH4vSqGh/Wnp9Vp6lGfNkC8lcvdd8wdJ60z4UiPI79axb0tashuWII
CYSvQYH0t5Kyl6+dDynY0OW4Wdp5iMeBBhmHjY/Pq4FqyM1/yb9HXTBA5CeTGfRe
XQDgzWFi1xM0eDU8TIERFhk4U1aao6RPdZQwZ8dO9MoX6DuuAzj5CFgAjETvZO/T
eil7KQxQuAm0g74BYgrs1gAAmltyqmpNPJB1vFBiiypkxYvoprfmj1wS8NmMQBz4
KAftOIhonr/fWlBaAmN2YHeaWxzraZO2yfeoMBTbu5SIg2BFGMGbzy51v3i9GOo4
AVi6fdHUzxrI8xFoI+zJhJ2CnwS5zVtF+mJqVQrkw6ouo6XjljRYPZDRmoGyxgk7
Atim2eztDSLyfISc5bYuHcbhhmbViuXPSlIE0ERfPAb2x9SXq747WvuL2bx2tSf/
9/O2mYjUUrcpSwLDM3PS22KzCAUcyQxIfXlQOTcZejX4ptmpXLFeR40sglAlDboG
5BX56qOTaXOdXoj0t632/lqGCZn1Bd7rxSEd6DxRClNflj6Ad5f5mHQiSmkZkRMu
MKgXnRnKRnaYy0Qcd/057H/re3/ZMtftO273s+TKzr3lzMgyOWK5gozeLSRtCx4H
y7QE/oBO9rTyVvwrZh6pIyulqrATJogEHVhAtuV/dt9if81FhRAizmzI3j5fQJDE
gqSsgFi782/youYDyzcEQu9vLjGadFWTnzlqMEoydlqa0IggMT6X0aM1d99e50FZ
Cb3jqPIaCJp9wsA3QRYBBLPfBeUdyFt8AXxfNq1QwNc1d7Sl9/FmpYSqG8WJtE9e
d8u73IY0iJNxs9oZ1c6y106QTu/MRonuSOJSOTK+oyuwT0a1OrzifmIEpPTTcJEq
0j6kGedfrwJtm+jCa+lrluEnAerA5sKpLTBTvP910P/TE/p82Me+q9llVGCkYk1a
hmqWS/QGhcIBjilxdXQJaoN+Cz3fnI6WOOJhGGsEyWU6wUT/OQ/8ZL1JjPEm9ybA
Gir96qLdQ8msWKvcTE08nZEYZtmCd2BNUWQbITUBFrN4FKobFi/ukDm8bFyCRynS
sFgoibsPNJmqxJ8rIGHS02Exa+gxycQAF6+B/CCFR7/MVy4GmO96URMZR5+5xHTf
frs79b8mh093qjxmt14sffifh4odMgBm+szC80AsYP/H0PEWiNWX7Z/WUjnH7afj
y+oCf89CFxvvf+eR3Rg4f8UgH463D0yoyBSOroM8BZMr8zc8PxMQIumDQ+L1r4GP
E7N/U/zaBrXBOozxN08iDg4MlCuTq+/3PkxKPEizLscWNch4DTyumEaRi6BuYlOu
gwgO9K6cTyvLb2gYHXSneVOZsiXNRdqws/SrqXdB7T1xOMWIjdl/UVUtAMAXKXWt
kLLTL+UpmIpNfuTbgtkbaCj8nhAGtrTKGR+YC+tZkTREzOrM7fC/V+QpIaSsZYzn
8HGTKMeEdm3UEaX8KTEQ2qfYNpOI7Yqmr6mCOrcym+yLcR9oFv3Xe7gtP2DP8bM9
DObwzAFpH7weQH1RL9wsNbcuIgydZT7NyaztdgieiM79AWzuy/6AR3XrnlJY5br3
7GFDoQtYwKVX5yl7H054N5tVbTJfgQL7wxq0zXG6bjmInk+B6wj4FUiT8FqpH96Q
R5VgCRm5gzkM4mLk/m02GcBKm2yfg9PNP66UikPQjcjgd7dHbxqEQILdv8lxCC9T
3xAfycuIcsXKBkKozAj5+l3jqUUSrNlLU4OQpDTJbLjmiGrx3ZqddKSz030zyAia
haiL3eo/MWLlCbpsSW7jGiM5Er8KLQnmYwFYc+LafmYHGtxEqbZhvRBh873f/j+w
zsQzLrdskENajlacdeGN1Tas7DxJTFiBJk7X3Ti5I7/AVX1KYGB7zjlUG7HgVDs2
MPBi25verJ6m4jkEWRzygNcpeamTyp3OhdwJlbGihR/SevHNukPA/YLD0wnhTxjE
zj6b5Js56bPDZnMJjfIEP/KZ+/D4inCBnDgwVM0d/A9+DJYNk3gbutPkxSbmGDzV
pqAgbXR293N4sBZMM/TkP9thjiQuzH8gQjZRLTJo3X21RiTOWWG9ncVWlvJgaqt9
MdKzJpBmR60tsPcpqR1xWjyBkHdSLbi1WEUTitv0pImlXYpyV3JTvcAxpgFjzuHz
iMuWWUqkEvHZ6XwxVkjOUsyWwuhuVwGG8/3V0kNdzXjImnqB1MQnICq7b0ft3JTP
wWcCZ67BFAvexI1oxVXgoc1gnZ5vFKHxioLA4yLNmpjlPTc/U48eHZfDaw2nv3eV
qiUIPEMyFcdi3nOZTULOI+tuQrEzTOcIxz21GqIpYpZkBwBXOCIKbXMzaNlhMoIf
IvzpNGvhwWzhDR/oxs2+6aLXtDzEcwMNt7tEQbj4BPz1EXMEidKtu1PkKtfqR1+G
LE/3BswOuu5mjM2uBkIVdAm5ilHQILpiedQhRZNlVyX8nK1+kv0NCVfWfrut8kzd
7HDfJGnKBcriKG1ZgfasBFjdelbzX93+aC/dB9FdIa/m6gPoGcriJEyb+pDgaPvS
uqEohlvqyYxgC1C0grqOS1o1ruSYhHbq6AhcXBgbpNbnm68g93GbVI/r/FndoR3k
KxKVEyrUDdQLxWFeKbzG90FpAYP0VmYw2heBMQOecuqEIZAUM6oGitJYTNub5GwJ
PNcQPyFCH1I5H/bh11WxkSh3PqWq/0wb2xJGEy0DKCwgkppZapSejVaK9UcZWLYy
h2UM7jiz36BGYrHh5v0hUy6tnG/VtdIh/R+jVqgpUcLDE3WNlqigLmVzdar+LBaj
RaLsp0exk/+F+XaXaf+N5NqGdyJAvSQM0c50wFf66oW1zuD4pVYzJbW0/vOKQLLb
zizAtCFkwzdP22dr7mZK2HCCvLMtleFYkonSNL4NlZ8tq8hiVsU4SMy/jvJ01ZEZ
WAbKdYD/HcUPFS2mauQL9cRMrGfL5OUtEt6vJNvk3JhcVNKf42WijojMqef/+aBw
jJLc+eygfVNZNEVkv1G6hk4DWH/4uva5RLgwKS4vZd5QQ775jUUcdXzA7tbldTDX
STbmt6rUFKfLfVRsST3ZwtJ0vC6oMxboZ7HlRKrPFFBsD8yszaqkXEKlA2kAa8WJ
coG05z/8QpLuSxNh1gbYFaPGpj6ZfdKK7rEC5+JTqWSEyLKdYYwKE1WNKS9qMhdu
LcEaQuPC+WQox2T8RjTj+ZMQvE40uErDLwV2ktmS8ItscAehCda1mLQ4qexh7tVv
tGfqZtCS/Sxp63GxDCDRk4GjUJ2mWOMgYXCAlqdjEo6oSOzkRZqkZi9mtjV0RTJb
aPVldUIsjZOkLyuRQFdXpj5hYYwbJSkCWlI1fIjVFWakiINfglw77LLhjqqCE5s4
vLyvw4mXCP8s3GM7zlDXOk2iDohXccxy5OUmnLk9mLVx/2hHAtedZDAUiUj50U7E
bh1jADXrF0OhK2IMJbrTGb7QKQfMrCr9XXPoud5+dSFKHJs4g1XwxhS3qGKt00SB
gFMFtoz+i1M+AwSU1NiZ2gFYXeFPNGn5aQcjMQ/SMCUjhzleL6mmprI7EK0w/ur8
1/VYyAga9GRlYA7tLyu6FJzQ/WSO+/acYGZtsqre/Kl+2rYZbbLNlKzPxHlKIrEa
7OzauGnVCKLWJRYbUzaAZhLxcvnp5t8i6B1yOShV09rYJcV4VoMpDMcL0tx32UGM
T/ej7bJF6vYcNS2Nq9S/suI8zeOr4FEPTKpaRA/OJYsVm+upUOUYXu/3XcrRWwKa
yjk6wSZ2LxR/6aMHF17QUtVpdJHt7cYJ+zxoyR10Qvzy/0ILrf5I66pAaDg+q1No
ulnOz5NmXb8b7t1pZptc2PO0G0MiJT/pgYn6DQ7uh6hYaTLS5ThR/stpz/h87Ho1
Zsx47DTz4+gvsB+tujSYayvQb34w2UIhUbQ1SOWSfCIVazWSVnx2SWRVJc2t5W2d
1WiLgl9puwElTYY4TieggAsFZL5I9Q4ZDt+G9hpW0+App2qY5G7POHaEkIVnJw4r
UjaOd+PlgWWQbnA0LGJc18v0VjBN8uRjX+AqrT9nP9OqbxhJTmJ0/9DUo5icl3yD
JuqIymEsCAZ8JLQmVamVnSE2cgSn2doZN8NkPB+OW8Xw9gjmDKvGINxWNmdwk2zq
PmGotZIm7HP+s3SUcQrzJO3gSAc9Jdy8xAwaWBGBKVqhCewy4WNG4C6YSatnFsRf
93Ad+OTv7GYO4kO2qeax2swDc8ExA0VRCgCQj3nltL24kyoaMbPcirxT2UxCYep/
y/A4rYXqrL5isHgqUHM+w0DBU44OZmFVhO52+Wu6bj5BwFjU+GxZCREZsXxhiJyc
FIrLdL+xjKJSTzYMpeYb2qJpGRWnf3isWSim2a72BnupTIycFeR0wYPXLdGqtJpu
b5h8OeL52m//bXvac6Eyi83QVbKbo2Ab++9He8apUfBaAmy9QO60fuNF3M8u70vM
mCdCpsQ86Hd/AkOU8uzrZAnTbmtMD8JS4j4GSMYb9uq10oxpGtkTz3bpn4AgZdpI
L++Z0evCXBIMos1YfAOIOHskW3BJQw4taEN3zSpY6Rtht/QLsWSKHVKSbMzEK/wc
FK0iXFWC/mNYkQq5IXlq14e2DMki0aH/zpukUGQ19AgL5jcjpkDLpcrlXo/cGJqJ
FbrrEa1coA/t951O6aYqjkFUHTrq7ee9pdpfR1sLISDm5Ohv4Z9L5pwKbzOddojy
MjUEUp+BCrhVc2QG4rEBOq7uEjUKNDrtQ32LtTSbVfzra0K67Br1gETVz0bF4AVi
eyPtvz4QSh90uVaZxAp5UZ7zAVgXnN23KTiVfXHEdrYRkQ6WdQBkaFzPZ5tAOhkn
+tg7oGV1J61BHk8Cg/eHssH7EDoaPkTaIn+GDKYHr1VUo6Q5Qa9SokXAzT9Zw5jp
mBEsNKR2kt0Rynnm8QtxNapBsVcjfnK0p6pIgB9qhsFvw5vsjmdRd3wRhPknEmo2
T3GQk36SidCUT1D9hBaFYlzZyNaUEhWT9P1QKKNsLP0HKISEb9+zvl8gyATmoXSv
g71FRrspcJHjXM/Z3wZBqjkKfzteAJ92bu2pEcpKcr6uFRoUVy3PbeslU7FgaNwm
9bOYoX7ITNjVsYkfhm8XL8u8oBouYdJZCyiPgiqF8x0wQwxbWYUoF+upSCoZkM86
rvcWzWSp6vzeCZT7tfHLlqnhJB5cUhwmZuC39F6zjI1GDlNaBJpyKDJ+/3YXtUFQ
9K7ev9S0eOPQzrBjOjpjwKGAAA12iw+2qvyZyFQidtH45jny5zRCJWy5RF/KtUrr
Le52AJOw5DPs7n54RqhJ+l31G12sgSY+2sBBcV2+DM0V5zg7gHAqfxpo7sPjx7va
yxiuvhDrmiUJwEsn20C3hTwCeqFSoI4zWNwtdafNt4dv/fHo1U6JirIhIkFTZ4td
rfLj2/EgTGCbeTvD5GUS2y2XUFPGcIfxtlHPpSPeV6ZEG1p6a3Ha5QjgrNi5U+BU
avNmZmXa8V3KTjUlsWDvoNYC/EDKYbqp/ny5zqna3WwlM84otHDhYzHFTI+3EQu4
oyn0zxy7ywdPtChHWe+izFTzSi35oNTOGaa22CjxopA///6UdSJUV5LDDuvFVrJa
X9HgiFg602gYaqB9T+sNxnP1jy8z+vBe7HQQ4IQc6tt8cipYy5G18hij5iIRJB5c
i04rHPwp0T4BV/4eNGOU8s1Au0hKsWkGftoGLGe6KhTwHmGyOAY4UhN1mmhAyGT3
xgMps+ddg4uQDTeZoLKmCSXFh7r+o6nuNbfXZvzyYSH7ecsGSRCGv+l8iUbdq9lR
wdDO4vPkYTonzWWNw3fnDpNicbHwCYu4+5iatnhrU1+Q2JENI6IMpBDYdRZxm49R
Tewikx6qvJSmc5z8v/t8qG0wY7TZA6hJFnfckjIIMGi1Ixmq3GEkXlnMPNdQFGO7
vr22tCcZiHrgr1v9zZNVZV1YOlrm9ZQd6r7Sb7xOSlTxb8wp+jv9Z+swCvbHFZWM
tvZTCrOIRw17wg+dW0Eja2uOmcuk+J9m+V8qLzJf+HH4QiJFUUsxmBQzVRcOWfDb
OKC5FSz1D1kSzsF53v183C1nEd811rIgTYa9H7eSG8Kdj4ziBK6OO/H5FTOz2EIb
chPBW1Ut/T/OyDJqiAnvz/IdqpXsz29HTfTB4iwq6DFw/Or4Dsif5lRgvfZ0UygM
9a+pvzwumVbm49nr4BdQkKPjCb7MTkqSKLP9UZJnRlB6jK9qwYWIVyqqLLuuN6Xb
G/Av2Nm9U6cjCMU4W0TBT1Hq8KW9HkfNata3SEBfMntH6V7EXhzE5VQUGr56lXBC
/pdIu8sCoFOx4XnXc4GgCeFwZ6V6+LOwRYAFxX/fXkF6QjLw6lCgPVvH5+pYqQMS
cbrx5wqLS8g7XBd/WpOn1I6MMHPcMV6d7YEeb1LC/Un7RKNIYYy+CNiNFyEKaVq6
MB+e+49qtGS5+4GkTRDj2UlZucYKQx50wQk4l6tlOS3NuVD+j1sEovPFFQPGPOhC
oQkPAlMI2RXa1znz9r7UQW8nPFfXcl2Vkrum/NKNkqLs/bperH/9IPK9zl04iRsp
vlkM5rpQlazG/xiSeC0LfJe1dTFu8kvgzpL5EyotorCIMzQoIy6s6m7LLZSNHi7r
EKboEu+Nw4ztWswcWEvm/2r8+Jwjj2BokWY/lwnnZSkcDWyWYRQv1r7ErCb2eT5o
8AQmh259K4qR/G1fMTzPWYVLqLbHWkgtjAl13RB+MsXN7tl7bufg95rpDHpQZM50
lpZPLcZtbn4aOSPo0pyAe1dHRMgmXBE7wdre/Ia54++5i04TIVV3wuUaPVjl471O
hIETviVPin/TA/z4OzwIzQ0QbDhf1A/WEZIUm1fVjf1vtpaTg7MNO56y8IbaEuWH
QrwpMT/3tfqRb7vbzi1SVAiCiwY/eWAZMLPhzLwpPVZCvb+b2ZKdWzqYyOhlyIbt
AiNs/K38yEV0Na+ehEop+tm8up2iUwEF9kPN9J6WN1QylSIZWa8+O0oYgWJaXc7B
hq3HtUeanjj43+s/cjkRtopkMAzmWAzQfGKyM2Wplw4InvxphshyCoPOk46kXcxw
QQIG/2gxSoPVS8KFEfdLawWgacIEEvwjMD++hePAYK6/q7c9eGX3RmOmTsh46sLP
nuMvYl7gcteB0Pr1luMz1VtaLEfMiByaqhCKvKrtatZiIKfdgkmxAbt/t3Lwy1AA
vWz1tnnyaN5/3BzQtmi6+BtTKZOHnpgqdpmDWYViLUZV208aoOB/+aPy/u/ARw2s
mDahcZWYBaez5i8/TtK2UdKrxfp5A4BKqTvn1rEKLUxRnIKMq9Tvivd5imC8gKN3
HWyW0/Fv0wzubu+lL6SCcKy/S44WI+b4ytSlgJPeauI+Ek6l2B7RG2o1gQ5tW5lo
D7Gqe5M5flRg9nwifaamBm28NNdMQFYB3j6mMxPkU9PlGSIJ72typgHA+dXQuDcb
zCg652/bRYFnB5FD5KDT2Xd1sy+DZG1kZ2gFwaJO/fFPiM3aXj+fazBDPtlNAu0j
CluXH770iUb1pOsGIEenYCm0PkMhZ1Z1YhvtCN59h+ofRw4LwsgsbunYcBG7WcFq
fVuvHLgOEM8ghIXqRaYZwI9Hc2weWcTn9q3whlWl5GGAUQt165F1RKWvU+qiCxyW
fzCNezUhOXDBfXxrVrOtI/6skKdddcbGeQ9aP5LRjqiyuoz2Vx1yiw2dL7W6yJQa
OJCu3FwNknZT6ARude7kEVWyQ3a9eN8w+UYPw2HdIYThUNowMZotLqCWWG8t8xWV
wuoWEXEyxHHHzUjQTgVhvz9rfkCb8habZz/dJvOd6il7d8ZYTXALt5T69O/0q/wJ
ag6X50O21tgu09Wj146V49GnbtAyumbK4K0lo9R/vVAircxx3I+XcmfVn8Q4IxeW
OB7wQfNBVaLohalo8ccPQQ7P3j6lquPRI9NL6UZLIQacQnqeCAjLKS2SaDXTsFsA
+kEGly590+J9wf8ESAfJaAp+ov9Ch7VSiExKPBtnkqg7/bK7+Gse4JN9pXBGrhse
4DE/mK68dECxANK+k98284kheMfgIj6nQs30KWhlRzb0Hi1/figoXg5GNCN7KNLD
x6SwgG+97KU0kqt+J/OzelEW8f11ThkAGKaucpm1mID1q3ue2PV89vSVKx4+6YwA
rV7l6q+rUKytuKiJM09o4rykpZplaMdxiHJ7Mgd7f9g9v+u5YaA1naofIrslaLo2
1P5/ujZRJTYikTWH1uyrHuDcKQE8BMCHvnRZnt5bKoCy8Kn1VAQ1Bl5s3ePqACHr
QIqOQtSqk1wFUHL4keIqim/lePzKbhoSxvbzN6oFoQ4dH4RC9dV0pEiclluvDCHI
fLirsJmIW1iBbISMj23WlHwk/lETowhiIEXj64EW5xio4qvKABMlnbPh++/+tLJo
DTXIYAVcQ3LflvF6zaMNYxCorbapjEdjV8evifbyzKL9l68zz28uFsO94Qgid8lJ
MzlpV047k4cI3onNxe8hGpYhsVPaB0GM69ehxVvOellbLpnnTThJAWw5QrMNxSIS
4cC6LVQUCyT2luc1DkZClDmthY9GAGd07TjwtAwsHRt5iZH/r/lVJrWZqZNaw3KG
A57xGofyGfbb76Sk3rQ0W1X82CvJmnnDaz21qrIkfl6y7wsrHeTHV+03hcxI1Y5J
YXCmg5R5oDPFDkERo/N2Wt0DUnHyhRzQ99HAGi1wYmIJlEnaXn7AiJObLOPhXkSg
JfSJs9aIjwWvLLeGSzD252Z265BTSAOCPKDEkLk+P7t+XQ4t/nj0wep8aZZkSTW/
P5OxIpty2Jre84GZcXPpiFkhNY+cDlv04Pizk5ndP+SvATFzbCDJAoueZmQXI8nP
rbt/c4/H/0aGCueiDUbqiFbMISUBpqehZ2lRfrD0JrNDyQrmUjI3rkRZVA6zSJcO
KNR6M0uTJE4zVt6kDD+I4OSnXdsCfAnip0jJGapKugjQBEceoDqLBbqGfL1/0239
DDg/1lJo0vF59upaJUixNrDLKtxZW2jye2K8EpQatagD0i7BFtn1D2Ur3z1+16LR
PSkGFZBVMq8jPsyL4ewTplyu2ouQGu92Pq0zd5enpC4lNdcfppiKM2IFXMB35flZ
slVY8yauWCApzfamV3wkM4G5avgWy61RXi69xa9BOb+9rWyhHeDDgPzcsSdUgTID
iX5tBIDjAMbSgTykqSIq9CZIcxf2wUQVZklIAb09wSD6Kq9X0K5Wz9+wSWN1qLVu
0z7NKsc4IV3Hg6V4JHhocZQnh/ItuGiPJEIdNiQE/01UsTYY58K1Ztw4a/idZ0xh
Z6wMzxEnJeJOIO90tNG6bTpvcTYvWxy8SfGtAVd66m7nrgszNMWgsTkc46w+F0bY
7Y9P0iamG10k6TxHZIykl81bLHiT2w7LcVZ3pv6BXSKRP2ppTvFA8h6iWGKQjHxb
2wge316Q3jSWZae5D4PC96KI9M4cg3FHHh3AslTYG/XdPC8wjkdwhK1FGBHXqfp4
/P6UPuMH/yA1sIdtEbCvujW91tPAnE8XtFcqf2H9yIQJ5tsdalBNMd1cAeWA0H+3
wEOHHm/WVp4DUjmV3XCeF6GDpVIuv+6pVNvW177JKLeM2ZMhMCr4AoVmKWeGKEKq
NIJNHwF0b4RHJDss0d9zvFlpHf1IE7SJdQZRrxoELEC6bWAqOg+Pt+g3XR7+ShPO
iq8cuS/kTSrGThll82lARb3NzDouVduLId4WBS+qoTXseDx5tKJoDcsEyeCOrjzR
KbODJrXwS5ikkofLV42RlfPVVQuQcjPz7IVWTBWXyblAkmhJibMqwojq9W1RQt9v
8yz0motrh8tIakgWUF+aMZyuDJHyfrKcZpmsyUa9iTyXE1mxJYv8Ar8cq5UbSikp
/OpFncDjb+y1tYHGknRKx9eBa5who/UaY13wH58Q0aOJ6h/H2L3FONAM3T/jm0XQ
8CdMN+WwOnS5LN0y05wg/IXZ16PvoJI63+H4hQ/LKL1UbhOno2CHLxNjjtbk5bxt
g3pH5IIGoLgfT+Rdbl9P0Yf0mcwm7ut3/OkJV1bFDdPMEBSlcBrbF3oU1VnBM4qk
5FjtjM4FdylbJW6fZ29PXBzjAxC+IcyXe9vVFFexYlnEiMv2vfx/CQukAue5aHaN
Nw0rYt6Ncf8XivK/zUCnbaprVt4zLoeAskS2a2yQVaUuF9/uuBUa+Ntlp4znBsqd
EdIvSR0cOTDIc43RsitwWkd6touz9BXqGD+8OGIZV0W/La2+eDC/PEFE4bPghOE+
4qtm99l4d9xq+2Xh8XJXswgGZ8sdFv9MpnCvp82KC3U3vQOvGkT2pExZZLiVLmgj
eRWHb0h5DHpCWNsJWQVW1HPfAq27TG7YedWqKbjlIyvsXHfGB6Z2cbaeDyV0zs1h
/YD90NQRJbyA+/OFmo6v6XKzQf7yHirKi51xFLrZ3cPvXSIf5jYcPkgHdCFkNhuk
ckzayz8zIAF2yDwaLvHfCQv4K25Slp6pDmlwTwCXAGAX61e192Bo2qyMoxWhdgfV
HncOrbmx5dJBLsfp0ut2BO4Mf2Wfn+VTfxzT9OF46owjwXB9T/nqIM65ZtNLjG0c
5HI2smH6JMylPXN3FT2krfL9rGL8B8inJyV4JkDoVVaAzmFL/JB/6bJTKYcfvLPd
FZwUtex8o/ww70OadYmMebKoGXGDasQ9EuyEvbX66TX7tUKhapjfG7xxttZ/hHwa
b/ICQw4wiESTq5I1dpyn2FuJyhhtSNT9shPwE+m0puyI0fghs/ObEg9tRjUwatP9
p66GN97Z5OjSIOQqYVvmyR4d3YMDdqIDfknfgemvkA5AOYS+X3QE4gs78Yn8yKaV
6QwgjcJF9wxCm4xw/66M/IX0i0hERvVhKAi1e5ibgt6tzCj8Lg1V76dQHn8Nyro6
e6P+a2vy0Lu56pGKVREX8WwKyXXjNjagaslwHGpvSYD1U7v979T7AeejLxK68Y/V
QRD8jV5iRcwmXlgi5i+grXPCDbtlEl811k768zXvYl/rV8togaHXnIQTb/TGMVCg
/u8TO2ffV+dPyDb2vXaQgwR3wA2uD8JL43lD9pR75RhRRsSKK7AQlIevl6IL+MH9
iMu3eC8o8oWKpMBLFwZdKfdZvSGhFh45q0+srwwxI6DumIqlXXZROtWGqPjZ/8NH
SpK7dGi/WOZ4PYbEEgOzMJYIOKQV8PRzuk1m0KnPrpnxB2DdJZ9XN9G7M81fZuYh
4aoDnc58Yyg5rK+WeOMd6ubGovu9S3vH7D1jFa47/9KkFQ3tycE1N8jeJI0NIxBf
8B1Kkb6apuTkgEtlyzlqXmD+BdzraypONM18wpIRwyD0tHsiCja6GnXC4O55n839
h/AdxmED3wlI+sOd0vAcf924A5Syr12zCtWWFN8MOBiV3VuXahLBoqrZ0CBEuRlz
iLwUwYvlgvK+ojfeIpBBl4JybA61YLWP1V6b5wCyZa5aXBJexsIbfp6cYv0STG0F
ojqEftDJHS4RT91kglxqz4Hy5c4Rj/SJvjEcFqYImpKwW325+lhBuUo96ciFjNje
qG6NAKJGXMgy9N2G6dSA9Jnl6GxqBt026fwhL+l+Egf+7mlVKIApQ25ujdPKBpZ0
YMh0pc2YWsNSUnO2QBsvNRmSEbfcn43EFz3K3qx0Lb33KGwi+0GRlSxgKhv6DcFL
LvcZrX1Zu66XYKbQvkkaEZPAbIHxeCSMvKs74AE6OQel9gYyvVb0SEDcMX8O8PLd
qFBevgThtkr6bjPbMajsb819FhSblN75pkMn/UVr79ar2jfCVb2ZQb9y0Fvw0DrA
WWogL1pBKTAN/DRMQfqWus67rnLDruOwtmWsA0pwLHqB7Pspt7M1gQgHE+iGtiCb
wZD6/4qpaGvh/XAiX8QlCkok0ccZF7/IT0t0hNfkUm7OKoU6q2IZLO/trMTwIFkb
gWg4Mmx2489v2e5a2yZaLdJktUzWWm/4aTJ9HkILBHhCAn6nvaEh4/oRt0sIFM36
UWsJrukKXs9gY29IH47WwJh/mo1F6lUYKUEk0VVdo87iHsn+0U8OEpDL3LGKzeP2
/HTk1jS2j+Eyf3S5EcogP0TU6ycxtYpn44rvuy+GtvuMzfwzG6GiawV5fHaYWghk
vPUtmQYOj8yzlCGWZUhhqIIAewY6hocVy7n6fAJha67AyMcxwGJOuI/HlJnxaq1z
7sB8jV4iClOSzv4bnkxx87WLUIlN0s6XWul6FSh8VIXspsiTyr3nzQy6BHy/WzNa
IKDdolco3xgYtS48YKBJlk8CJrnW8htJJ6lP86ySz5WsIJ+tlB7vgIhr2Y3jzhM+
NUvfQ+mDwDTHs+miHUGmTN6rFYLx+5oN6n6mMg5hbaHaELnoL5HWUCJsQbF+uZVT
S+hOitmAnDunbXRVEHWQit5wjGGw6QdiBiVJHKC3X25+iwIlFLF+jsRHTsMq6urz
V+t5lSD1yMWBni0hGt3RN9dOMAoQXc4ai7Y6G6gVhMo+2EiQxOqBxVzxdN6g9X56
m+JPgxa8BjNO0fZymNR8Yx14dnB3vk2lT1YoXgYVstegs6k0cosQXoLgagkx/xIn
vIUOurkVrn5HMfr2+V+i/vSrX4nsboF7yAsXBU+GxxzdUj+LPyhew8DyemG/Pw54
VI1feKldW8SK4nywOk0o2e7zqUMR+AMmTYScLcIdThEPGSuZ/k5RlmhvrVkYV+d/
Fj4SG35xE3RQZN60eDXZ1q9hAbUojNyRQrMCz3wlYGzg3RJxCT3vnz0WyN4KdwJ3
7F+nX8I8gOG0n2r1IRMtVaM03OITmb6KTn6FRmykpISJER97N5Yff3PPrxFH1+R8
myld1r/9iexHx0j8sAGVb+FkUzYjSGx/KSS2mm8FKeNDzErqpuYuHcspAZSwm1jA
sK4VUZxDQSzO1mNYz69NOUnl3w6ATXB458Awxj+FL/tOcHGVmhoS32C55nPU4B0F
F/mk7gmp7i31WTnW/DUu2K9pEkvBgHQuOzLDR0rLSIkt+cO8f42LJCpUGHL8rizA
ECQcJxCcj9MCtbF0hOC4lcpy13iW/hEZWbEJnZantZVUUBpMRuYTPo6MJoW3VS1l
Qk13C7ejVdwrR74VJ0c+DI7K0rBo0Y35peFSNcfr5pnScAc/cdL84oReR4xcdFqh
NWxTqdwn9C5g6LzfYnS8HUsgnt6tl4rK06JsrBx6E0SasckTd4ci2USVdubTO5u+
dlthcdMm5QyflFpQoY3k23gJ/+lVJeEfVN0W/z39pz2cZe44cSEq0kOA2QO7/epU
5urEvygxXIGSCAspfsdm4LZ3ftp/jZqZDLmE3Syg/dKc72+iu2ep+b1kA2anZY7v
QATGD8X4t6gAB0mACCcZ8tuJQJhgyBRf4x7wHQgYjs9gCtXSPGI+JndTeeId++53
0h8sb0vv6ret6+RzPQhO5Dmd5+pkJCyMnPJzqa1XmAytnfLg1u5s3AXVNkyvE3xk
UZf2TN/sQxBkXaajiBvmkvMenwmUAF9bEEJoj20jLXKatUFhKB8J2Ci92xotAI6P
64LX8eIpzJ2/cBU5f4cqEcmUhoG+/BXN/ECmzrN7bLDvz604AGdaU65Md4PliD9G
BX2beGfizWeOWsDEsS2JCfsZ3J4fMlibUUZIvV2VMsp1kawi+d67Mx02vWUzHrd3
ss1fz7Kk19D+LHqmg8o89r4ipwAOijP6COcy8APIq/pu94sLZk1fBnVhz7gSVGPt
Ij+OsNQyJpm0jxBtQ2I4kAzaK71WgzZhUMEvKoE5ro1/yh4V2cskCErznqUK3EJz
4Oo/3juCWjGsC3a8ysMw2GNWCjelt+ZMZgvpTwt+4qVCpqjLC7KEGrh4xGZR09rl
pD7OfPm1PwH412UtprTNWxWdW+gCu/e1zSGs2s5ppyOK6jePwNHocdtWuzUxhC5I
/IJGm73BptEWBOMv/s0JFLiQUr5L89HRmK+o4Wd0YYiYgCDy/rYvLPOmZHvGHbYC
75yEB44N1d3BN1EGv8AkdrxhfmhjvB2HUzw1sIliE5QcouQ1jdEny8kHhgiRvNYu
jGw51wh2Mzgip59JrLXOFluUsRzTTL7GsBHj2RKubMKQ46Hz2flGZSDcmd8Ui6/G
axp9w8FR2F6/3USYYk6CG6aLLweLnzXZ2OqgZqX58TIpZgZJHMELtikypaxSsILN
BcTFANpywh5915B/PbMqCDIu3eE04QfwhEwgsHi0xkz2YdGCLozdIkDeqNlbBq1q
bNuVxDq+Mkjej56kBPg/UkERLdx7wXJKSmVVjY/CamEKjNpmNW2+e3VC3hbQKbnU
E0KOWEGXxhxlf35rfbKfaWnl4z8u1gVTmlUBFnwpiXe+5hOmmjCySYp4s8ic/Kv/
OYZpjCpPAesV3+/jro7DWCWIwIl1KvF2s34O7F2GVBq1J/KQ3TlSO8Xom0ooDM6J
btKEYMfGxUiSF5VUENtE1yOKq7yP3y/KYbFWLtZw/xyXLI0vNJDeh45QYEelcc5e
xvUiwR3yQ1jCJYJIoGB9hrjvcgmkc3Vq9rw5T08j6LQYvc1fLsBrKuFbkGYh/X97
lcVmgaAQmh+5jd6Scw+Zce0iP1gHFAfGMdSksveasF0oQWyyIn9nej4ToNjjQp26
JQVtaxa031QfcynIVZIV5K5y7LA0BOhqfb95XVLxkxRG0l9gFLThjXxIbNEcG2fA
2X/QzjKExs8RXdbUt7nzFvzM5ngrjkF9eSLYkMpDdYrgsvzOmYeHZKA7eRkGzQFH
L2gF9PFcOLDtuapZ3/uFaUvgDP7LNmV5egdYSiVpZvxogPFTv+xC7LHvdpLyNUww
t7yrfaRnW8mNKUrCDzT1NPSWR4t0DlRNy0BpEetdlVWZJ2vymZtRkCubMqNfkr7D
dtE9Zn9+IXq1GiGBNH4BLBc68Yt4rOtNvHAidtfgtAg7Crm6QQOXeBjcCvhfTNmQ
0kDTcL3k4h52+yQQKqzSLnr4bpzV1uEMFQzqq0icIhOEz4nbkziOsnlt5Xcv+Q7B
G4Qg9xEEdeaHwnLqzt932J0oYO1MVjWM9U+iwFW4cVNnaMdB/rhneDo33ZWyiYr9
dBbKZcoZa36IOc0LeVhV4bxec3GLuVyxQ1I6YQA+ZJJWPR7B9ibny7rGSi0ms4oZ
Mepe+o/tu8vCXbtZM51TCxaaA2PT37kwfz9lLLsp/KHQ8nxo2wf/tlBCoy6NuwUy
BA7+lrNXAMcPmTZbB2Imh7r2SG66IUdFPzc6tJtAuvqiIML/ag5wMJ30MoUNSrXu
OMqGKUDDPDbo6r+jy3in5r4q9f+J/Ky586ARwFMbo7JNRNEzyEpBfVtKJvIPNhL7
YgOgzhKCywAFclZGsVrXh7BZbW/t1iq2L0KZVBC13ByyQq5DXAK+rwgc8jPDCIh6
/jWf84v9T+YTk3uZiA2d58A6t78UDVeIP28XF1Pp6o1z4vn1s95olfY05mRkY77j
gYEKJI+/5kYFs8akxpI2QSlVgwC4IZsYhQozTVSLD5pMLcaQ8u070MVExPfZuSrA
FJKqopvWb2bQVCRSyvnBkBIo2y6nIHMb9i4/NH4115+zr/5qrFq1Ren03xrYZ+uF
vNM2c/lhKQt6dAmB13PeHbXE2EDS2g3jcr6fvKNyZ4i9JuvhAVCc49ItFcavMUTZ
oz3p92BIbf/XzL7PbluVqrPIoSsg0ZyTFlWJwuhs8iBDtdq5JfYooMBlqPRaW3D6
fEb2P41je4LlfinUgsUcn96vwD1PepwUkFBsJc7XYhu/TQBSXKsto9eh6mJVtlM9
XM1Dsj5Rn+N6V8GovGezjTkAngCkIiwNY8mTjC/mxcPRLlIYEHnOrj1VJRKC5O5u
BZog75C8LrrS2pooOv1g/KqDGLHdGd6EGM92ugh2nKGUOiE79vY6FTYvshBg/8sA
sV05hAbIrs/0edUErtmivjb6dOjbpg7213RW3QHEkRy9XWIWGj9wG8bYBhpoy2lE
tKBD6COH+Hyue7gK0UwtWTVVjY6yR7TZQab8Xl+PdOfMNLgU3vjA13QurqXQXaoQ
pYZVm5wfof7bDZ7BXYDFEvBbIOTzuBCdgvEq59EjWStEl+knxo+BcZ6ElZgIHVr6
cpz8x9U3IWSWkgDYAVKRUvzwOVZB1GesZ6zbYuoX8w/nRbXuHGesHnVfKSRTq+oR
lVx6E/Z2w8REK8+jbqeSVOEgA4+AOMv7YfniQsAWPbCGa1hQJiO6BnFM5dHjV9vG
/Pg0bFl2tXvlHIP/GcOHsK7NXA1FTZ0iSoGa33vZzUb7wvdJ6mpiwX322CNWhLLN
l+uctBqH49EoyBGpsoEdGua9UgC290j859HlFrdA6Dfbwyq9SO1uQ/mMrs4uZrDa
aUv1bdufOu/UcUQ6/9UwcgOOr4QV1akOck7AY0BysJcnEuUwo7Be5DwfEKi7dxjm
hyGrU8s3ov1yTSNZbIvaKoteA5Kd0iAOk/Jn3Mpp4f7/jtnCNlQzcNeWVJ/EPo+K
Yo5ZODoQrgTr160KqpP9QaqlrcEsMzLBf5kiwqm8XO0ew8QmVpJTMzRoqXCRoWLg
Bq+E9huWJd/mEGuo5PS2eeE1TKdKht4xjvqaEu3Nl79OS+nIumY5Ah7q0aKFSXG0
KXRGk2eT3daZF3u6XY0Fx82Tql7XhsVnlErdVlw4gvS7Q6d2yDdeQJlndCZaA19Y
vZ7rTNDG2MGh9TS6G4Q6K0OVK2hQccDD82XcYbm6OKocKd7fr6w45p2dO9wLmLJe
UMHpLh9shwIthaaKDf/nkaNxD65rLMlbXYotM1xDeqNPH2kZwM+70yzdbTMx2m5A
TQs2TmHXBMhWc+gPdffqivu5D8V1FBocWlnkeNVvQKCbsQ/YoWQXVQOcXMTKkoba
Tv+UyZziVTx0g1mKbHui3XKLd2/U8MfMZ85AwzEUnMhPRptgtv7o0U9RliOFAJzr
B5NYdhJOvPLeDxIZnCjUVL/1WBWSatule/txGWW6QzQDkk/ZHirpJwDJFWeWdyY6
6pqiFTo0x0ojdaHwq85smvSdZCS0pSq8uWaafvhXWINE6nAwsZeEPb6TAGRxNghk
jwpayedfvjNT1B5BJNZGueMq9T++DjUa7EKiUfWYAlapGrZp9AWx5MOllN4qqR7g
2jeIM1bpSvd5xD8/0SMXAxej/hsPCyLSCilzbMh6Ogt3FhKDg7R9tyet5m4GsMJx
SKyILaTdT8dUIjz3xgNL/8dctXhanZR+dnfSACzPpHtNdiMC2akAbwEezWLLTE2A
cw4I7oIn18ZO1j0Elk6pbWONRsoGuhsk3RsNYBTM6W/0/hjd24w7E4sveqLurgrx
5D5uFBVbDvP4UzJcBOaIl3MilprbT3ITq056RFFz9/yrif9whVBMdVTN8fLLPHTo
x5b/omIaSTiALbsqyXkTzXDNr71rpRO9fD54f9QcOxrrgL8ar/2zZ1l36+mHXZcz
6q80Arewcq35l8uXMzVAsmMT7y6yU1k7jaTQRgb3WuiH5dFbqXVKPnPxTaIUFkKW
X69sVBlJDtWb9GjhInGYgMW8JRhqHhNs8jyRPtd7SAFy4jOEQ8AMuDX+D76SR3fW
qdGFsDGk/ia7m9HM20l2lwT53u7L8GooUV+YLCsdkJ8QptSSLGDbMEZFgRPYJNy3
AS+8aQ6EWiGvVgPf0Tru0p+2HpQ4QI0Lax9+Ed2oC1RYvGcPuh5r/EvXtLOKybNJ
YX4RwZA9tMSw/yPEDzIV3pqOkOb2HQe0rD5tSPLxGiRdx8KwaaYxjiaX2r+Uu/F6
xbHsnoUJ5n0HZPUqXGETCOocZQaQRhnsou+BeSvgUshypY+echgZ+IEuL9FJ06up
aXvpJbr0CGI8wO0QjYg+DXnkz5vu6cT/YErlY+wE1dtEdStjWJytk/WYETJMI5WG
SwkBL8xObAUvH0hDh0ZUZc6VsAaKuz9JmwdvAVyDp/sQRzuTQM3Ay13KmhnWxCyc
e41vabV9QzZPCHGmBagcRmqF+7Qwh5JzztQiOXfuZihbL5hSliU/1iAx6TURlal1
Ybf3XSfVbgO6zskm4EVNbdwr7UOpow/fR61R2YNnTVmj9ZgypvDv0mLbRINfcO7c
4LNMaGSO5PoFoh5hmjwkpetZAm6Nx6KZEiLKqw1U4Lz7Yc+liKTtcC4FuMnvHOo7
JoX/UdO1rjbXMiQbSt09B7+7PIJ1W+U3a/RTgVoyVUpXf1ATfMa3JFqHDG3CydkG
GXQRQ0PERY/lD8QD3adIoldMoN8aPLG6cBqEPEwRq4lKbuotJNPqTWNOrCNjqskC
0mRF+ETqM7UthQ50qd/ELw1SDeCqDqNTNCVUiAg/kHzLU+evuLAnZ7+ijXQ06NgB
Cnu6j4J7zkzVs7Kf7H9i0hz4Ql8jKpi30OIEpj5GZOu3LInXvsXUaES40WVgKspx
fcWBhN5vDUk/bFzTZKmRIld5mArD/RHyzwk+saTG12jU1Jem9bGNb5w9TdrcBgqv
0zPKToE5acuzIqU6fkzQfbDMCZGJZLABWz9cYb/AEFvVsGhIwCQGuXlLOFPUkeDV
IHrDwutkBfih7ERVJ/lHhvSJlITKdB/bOD0MSlg+P2Bg5ikmvQaT/yyYi13P3Ii1
yByS/dd/J/HchkWYKW+ThJGDjgWSdJFAVAeGm6qk3bk22Jm5GFdceQ/FdLpRv8NR
g+rxXCwiqMmD7MuBZoCmAziqqyFwN75Oc8F1hVOWh1LFAyBpsNkzZ/dMnChmcV6h
HiUl9X+Hw7KKwssB1o1W/J8lsI1AH0ENU2IbCiutrHoEU4f1cJM4q+eX8tRcpDwh
JBIGrDb1uwzM85AwkNshOksuCKNlgSYG72403ZoVTHM4rLGzUgmVTRQxsyv0BJ3Q
bBfdjA6ssnEssI4ILxcj+xAI98t1fa/Su8f4jWA/S6wHJbvFrZuYW839LIARtnqU
TCXr+gpjx0gNyxtRe0FjktgU8N0hw8ExZEYtl8yuzQtJwh0V28f9InNCHEorU6hP
ZfYFZcP5Ysf+nmrPuxqq2G9rEHDOF5knrCNA7t50metHvyG5yaUJ8VK1YB29e5wd
AZdmZi23xyE3J0xwEKMX2lsMN+eARg79wS09VpshW/rMpXM0XRWgrm8pB+05VlaP
sq3ExeCdiNQnH+hpOTKR/ubUGXvV1W05+pYsRRWPHOpVYQxElaCJL+jes6OuLJ7h
zxVJn4qbnBv3ou/++oTAC1XgjwoIjLkqcFhfmBsg/NtIgvJyn3miJOYJymyINptG
mQo/WoXzWz+Swfvx6rMMB6ojRFGM0yffELSHoRg/Tpb1Jh6vgyVHb2kYA56Z+7QQ
bkvSAzjVbOiW3kW7VxihaTCm+JD7GaRGxlFvKC2KFUDR2OnoxRrJe8/azq0y1IBM
6A6leS7zPSyTFX8jR6//ifZphd0ssOezNg/w+Mg5cpCv1+MI0Qo9rN2vfYSn00UD
iYQaGS4+K8mUbpz8FU/J4miwo+6FDcE/SdmHnyLvwQQKYDIkSC5SdN6r/VSwTJbr
YWM2ywdga8hPFquaBQxVzpIyELh+zEiA9Hl97i3PqAi5vmm2i7m7WdN6pCilsHxJ
PgmVbB0pCGqFZ+Bm4dzr8LzonkacYGlVwaw6zXFeRZMtM33yRvOf7I+jOOD80fQ1
s5jl1u40CsQORnDye6qNYXgo0dPDyGI+z+At0sXeT/JlHPzBX1PQSwvlRq/30++f
XvVZksULOYPqauppFcVfYSpTFR6DS4fXTpv8uBv3g+q+zvp/acTBPGjOgWA277Hx
LNAORoyN3Cll/+q2DrpmU/zCAjk5opA8a7f8xvc/zZMGcwgNjowxIQ5IYEgTe27y
abgyBZKkrhQhTP5U6fXUklByGcP87Kf3iEYhJI0V4BQFe7ebB8+FGHkTbPdc8SFs
XXJd1+ilHXkfLQ4cbEgwRAp42UtFUbhqqezL4xrBg50Q1k5aPDlTbdsP+TxgrC4x
aPX4x30TJUwD9YgEq60jgdCoFOYw1VqmqJPoZrb5SyJ2smlNT5/5HPHB+UTsujef
xw74XC2aLxgO5x/k5bQbrRscE5gZppFKe++qpCYSB3dXI/B4eL1LTcx9FKA0j6R7
3rnzoeru7Xv56boJfKytpo9VcSMh8hWXe3icygRMZu+4jbrjsFbyuJYfeM86eXx9
rTgua9O2Dp3QgPXnNYug4RVptOJ4vTvoqEJ0mdKG3pZgxQsoCoOlFuV/3CNYhUeU
7+YaMh3QucS4hxPzJ+7ViZWFwn8a8VwwvDXCuB7bILA6zSqqqZ/t5vShE2LJosTT
ocDdOEY1qqhEh/6tCxBsvaF1pFcGBTOPYY4+m2zF7aRRZTisHGLqbrzra3jv8P1X
JF0lyPhsoagdWB0Cs9Z11t3Ha/BGXdZtOerIw2NWB9HQEhRMC2N+Pg9NG8UEU9Cf
iMC4xGWK8yKfkIh86j24b3sgpDQ/w70rCzjwDp1jX1vhgee6HEFFdLZdQOwWBKsi
LJN7qBEBgpeIOKWP0/U4ixIoFdXVUniB3oApoutt6zes/d2gz5sxRUD661WTTnqI
nKv74baeeeiO67CdbEY60pxuSDyocNHvC3FZrhEmrKWVWrW7moX9eRRjYF7ceaQx
fiy6XYrxmLU6Vr+SPVaPJhGrnZtj8MaF5TBKpa3or6MA0FLpey1XGyVxfSAm9rnT
Ya9Rw0eq4+oz9mve5BIlR61ySxufdxuKgViUlKer54pHPkQuvRANLS/BGXoxkz2H
IP07etNzNRvsGURsIcaKEJWcG28P2sDeSNxj+Cd1hu/da0OBkJw3YQnjx1Xzdukp
9FN7Xls7+H9g36b2BTd7Izmb0DBw+I/bmYbztZ2VF+NTsWfQsqgLgnZIJ8qJ8hWt
VT3jTXh2cjKHlD81QdDbJ0B8FYa54Isj0HD+pI9XvqbVgXzk0AcTQl8Omql6QpPA
rZwNQrpqwMbyrX9uu3pHDo4G9ngOjUjo8a8niVhTZcoX07yFU0fgA+dj6IVbVMtJ
T6SyCpI/cbEx68dusXtuN0XDkvNkchQZTexFcuEzFB/1I/TEOXsCgqcBKggU97Kb
rl0zs73uxrvuBdpvfHj5Sf90v//gQsyGTuB7lstZpO/F+0A96lj6qnotrkBiHnEO
nZOMKmVciq8nd0NpaqCyKsVzJa8tWpeelSAQQTyDwAM2b18hrjt3Y9vlSH5vKd9S
f0dAkV2NlEg4zaAW6APLBu/kMxJNGqjWMjQODo6iAosZyPoXXMRf+DMb/XxqQbkM
PhIiWdoZ1oAZd6uJevh/b4QGj/WgBgWQBsZsgl/4hYBhMAMUmkQtGtNqY6bRtZ85
QV/Q91u15P4QQUtpu+c77RSjF4BcOVDNayjWZk9fJsYBlQIve4oDKk7Qw0eTrsJ4
twD4yjMX71xDqN+c6UmEJ/GCqAMNUpblxhoqe+Aq23MgfhIu/L4Qt3QclUulDnIv
w1nmrU4VEnAHY+DIWi9O/KzbjYORDD7uMXfwx7+9ckYsntarMb7L1ta6ud6Shgzv
41KYmlFUW6INzztSOeWc1fq8T3y2laevNJwaszab+da5ariQN7nBcVoXZQ3hREOo
/KMq/SjZbDRV6dY+S0/nQdyymVV5FbFbs1ivfM8xpsHsiYHzUgCL03TwlliTzT0I
IoPS/WnoBcJeqqGdT3PWJth2ClAfaQdFEDuUuKjmM/EZvipB+Zb3mawAaw6vroy5
iEoaonW/KRbTw9dRx36+XX5AtTHTtdhKGHnLv5HhX7ocXRAnJ1Et1J/s5gymha/9
jlQuKv3MCb5yCkWczeeN7fafLc2hSaaYQhJp4cP0Q3yKwYP4jkCyI7TkJdvF33fu
7P7RjZFOyHWWjxJD3bwBf+VvUCclO6ogVs64NH125+bemjeYFTmhMnYLTPSJ8bH/
6OU3tm3W7610mMWtaPviRKb2YBOjZ5NiSJrKlb3L98TAPQ8Vt2TNw+6GFIGmFcxI
R3FUbe4YCXiAW2zNL330qQQZL6VoOZaW+/A5CHqfMa30Ef874dC0BSr3kfAaNmYg
lmzMkcKFWlDFhcwGiujLrEyOC0UZAvz1y9VWqwcVl+x44/Wrb5Xs/djZSR7U9fgC
22lUs1nwGAtqRFd2cJlJPGRyL4bFPyGt0ityrtb7eAylLg8cQ/4nauHiO1S7yJ2H
Qx9vY1784fDN2DeQ7EfzgyKYA9iaL7toVA36OwnQuwxUF0qrDpL1YtkUk3I74nY4
ecj0IBB1+glziBZi1Chyfa18dxRCQU0PI/cSdaNbTDnui5U4QAOZBXHRyt5NhUm8
qBFlOjd8xIIPjlN+6nR/HuuwTdnwvCYxqf8jHqg/bkbOrnVIwTRjHsCU/OWODop3
D6hmuk9CEcHuDLk5o9E95oeyG5jHQ10rSdKdTK5BxYrmvnFmb2ygdqmy8kdljBqX
rXeZbu3bHlZ7SzPhiYu1SHnckluzI8MbV4CNzx4Rrzqrs5lOValkM3/wSQUeq/lK
rcB2B/gU/0E82vgocLSt1O4f5Zm4GvH74ddLTCM3Hgcf8mFWi+m5yJ6ftMujJRhk
/oFLoza45298rNp6Ulc71M/rrEPq4ZsyFga1yCjekF56qAGBdmegA+f6HFcpHsd5
a8uxO8GnQKEd1FS85TJclvXrewn0AYR5uSoCMsUcg00ioN7i9wagxLcUIyZAvV6b
oFJpMaL6WuepLkJnY7KQkzmX0EDspQkd3wG3FxzYdxQE0liCoOIplEJc2ziaFhs+
s+6I4eaa7eRlrWCPXwHjYzRKw5sUP+E2r5L7/Z0hNPKauUiYhqBARwtoMa6YVNYE
oeLdHBW/Xu6T3FAYQc1XfJDG+Ft7VYySmNg+vWVebNWRBHYUhdavCnyN/0OcKbB2
5PspaaUjci3lDh/MnJjRQGsFJs49IKaFW761q4PlppIv/sYey9fh2TyJ5DTrROkN
VFp/9qq54f0E4F3bNHvkKfJGLsOH9UbyMFSs8SGQu3vxHfBverrYzqL3jklU9wsF
Tzg/qVv473tAUJkku9JG4RXd+atPcVX8oFFNEHX4gT9UK/2CegPvjmkUPZ+SDXUs
qBSvlYgVaV3QimSwT/UxThmlrC0acG8Is88eqD5XTAMX+OtfohkIOaqf9IJNBu1H
q4++wDzXg4QOc+lCLYAmfTg+wrkZYaTEFDdqp0zJQSPVm/gqwnjJ4wuesTytbb7Z
btEXr+IA/uExbiAd1IEixEvoSdyUwcNwjIUxyVqEsUnX5vNhygRKGi6af+3jN4eS
PR2jf74fQ/45Bl8c9UAqaF/Q2G0wCWKHu02nYVF1HURoveuoAJZAL01M080UAaPy
2zdTkjcyekT955dhem7IFiwWGNZPQNFatJjhInHtYYSCKgc4s9Ck7S2/oNymgglv
/vOTAXnJXZVDgyLjPfOWVBoH1pXwIsarlDLDzuuQlX0HdZUy2pNx6d83Q50WFDRY
IHr8EpUOHIwLeJg6hs3QktxTGq8tzuFW9I6xEAt+yW4LGkiFE0BIeVduQKlejtOy
qyD4288IamIcP/tSw+BazO7KCdRI0IpFO/X40L7sgpGtsRHUtR3plghQ0jvhWII4
ORkQebJIj0WUCVmyc8D0wi4f0yJu2++eVBkiZgvoV/Z5hvuIJ+H0wnklUzVydOj3
z0e3FGfSZKJho8AtjH3FeygV9rnaFGsEa5I+wxuElXqriMf/Xp7NwZjrcTuN7/g0
JZVhgUYo9yLK4uY/vscyVfwV4VczO0bQ3IB9OlPkvilbN9iNNKb8Mj3OqdpEUDYa
H+H09wTD787uW/EAoy5B7zR0nDPg98a0B9nw1N1fqwa79oxxJIM7pSKdkx7j+pOs
zLRRX383deS+1ZEQ9K4U5k5tYfVpqvjOCC+W4ZA6udCJJp/P3AkiXPBeC/TxEeta
jv9tBNq4zVLvuim2o04RBoJCD0ZOQ491/r1v65NPFBUMb/kmUYSBoI6bsEpHtSSd
sRyb9pB7Ex/V91xX/7l7k/lllL2VdtYeppV8vv5BtCERfk7DESmtkPCEdHQZ/TS7
SNR+SLDemJT9/pCD33sReu2vUzNXHpWo6TrboY57zxUtMxxUc4Anmc/i9EObbuyi
PJIiSqKGRUcMa0Maa0tRtJFrEQxCzWdM+mgf7JyugVV7IvGik4O6wd6xXKTEP+Qk
9xqCPzTpWyXSusM5D7a1IRVRtjeMY3N05UzAXwAB1+e1D3/BgafjQs/Ky8Pc0Tax
rdqGrE/fg2XKTPVDWMIbrIvcCz5v8hcKopxqSBs3LzCOTX2iEeZEdFxUjCbeg/3+
tvYRNQgUzwPWeCL0GcDZFAdBCSxj8G4FI3Qej1/yX2DvpZ3QQ/DQvHn+ILvNpN4F
YIkJdjvzPmh4c3Kp3KRXK9UqeETQelIHOGCZVlnBkqmn6v4KIFdZKh+2f+Gl2Q9i
h16TpaBZTB8Wbo4xMNqQFMRMdxSrhtkYTbmiWJzvuTMUxGGa7rsNc7FKi5fbOKjH
Rmp6Jy1GXGbcGkOl1w/a7+4r0dMgsi0U0mPn+WWDUODPpY7sFnxinTyYJGv6Xqqc
HLHAFNs/pRCT61Z7KhgI8OouVEosnMsCy5Yz6AtWkUET6IBeSDU9Sf/VX9YNcD8b
zbgEBlLhNeA/kffbiz8V6ruo2TpmaE5iVGet5laYE3/pMyES9yiUad0q9OxG8ibx
d8hudWnoAeReBeQ83PMUjxkFEv2Z0x9AwfD3MjSF7z3GMdfb25EfbLtchRLj1Exd
pxhmlWMIpdzDrH8qI1XlSbY3msmQaTERsS5UP7PA8jS5EMweDE40PPLBpbF8MbWZ
jHZOhd5XDSI+qFaeA6/9gsAv2atE3Zo7w4sliB3uo5F1xL8eqOBhdUv900kdpidB
2F57TVEy+rIQOTelnc6uNzt608q3Vl/jvWEzl2EHCIO/E00lV0q7Krjzyan64SwV
jC4ivkMbOAlVxCFL/PTC4vsjx6zn6JMEHdYRMcgftRXpt2Zocm8mXdvb2fhS9+mk
kKqFyLVI87QaR9u7LTBp6g9tHa13U1gDWg9m8zwBZw60gN0mj613+divihDmH+rN
2si3quXvArNb/ySmTCEXojs9MUiDnehfdPLKLDgfOsW8fBwb4Vpo0TQtygJuBE+h
72d+eZF7tZGJVNMlP3fKfka4ApvShUrHQcIqAYttlZDEV4bFQMdK31NDeyMlBS4Z
uEg6pp5GW10xyNnPo4lfhMVXVCdBKi/Abw0rD1+UOQdCj3knZatCcaB9KoWh4sF1
h52bDRLdaYI2f69SuwapZf0KVZcF8AbeYa8RmJNvrQY9nW3iLUEtdVWGMZGShj1L
xAp53fcCjsVds3Rwmx+cH0fFAu79HN/6g4Fj1dZtQ2p/5CPDp4w0LZPHhL7CINOQ
/COp6g31IxFQLGuaPGkEizQeOOKSPOHP/uSesJN1sp0lNuPuRJ9tOdSIxtAu7uWV
n9rk7OGKY/WtqK+DShZhNNBDE0I+QWJFt/K1ZTX+TZ0Z5HOW4ozuZamEEoYbmEkR
nQx7Fvyz1TxDJkaeGpw2JUqtxi4uwj7UGN7JhhTwLBOL3Op3cyOHO4Pq5pysljwO
0KrCAUXXxGxCFequP9P8e+n7Ipb5E3w/lj7cTEdi/LxPuW1ACGDwIHUh7LXov+Jq
sL5YpZqF9WbpOdvzLcjMRcTOoQrfhZBdC1D2W8km29jQ4eCUs4lDujABGFV3a9E+
MCNH6KPV/rxYaqCwttdOwrOHOAc7F655fUpPN9CDAsR/K3HvNIoYbDLYpZ++pPll
0GxRwzirzHyNxMmjXcx4+HlA/PWV6xaZ3OyeiayTbr6mIubc8W5pFKkeBpmxqQga
jYKKqwEa70jKv+4LMG9Ch1HgWSTgZfJZQWBJu+cGBRMvOaLEsTobDoLaK7v96k+4
Tt0e0pWKoSWdGl3/rk2p8pkC8+HleIY5qgsF9TBGEUl5m3kqOzS5FLSFX/HK5X3f
NP3tV+a9Ml0lfN8J3y6ONLJmKyu9uVCxXxsQ680LgvN0KDDcmazi3qTuUN7Mhz9k
I/ObjD5IHc8Ehrjpokrxc+XVTEcwHNMN3LlK4pHUNOaLTDd1oXvGTVfMy+RxGvhh
njagGMwePmqIvOXhu0o32+IHpKRO6WX2DEMnbGTfWEXiRfFmVQOeUJzF9qPNoYPH
br0CKrPMCRlwCXfRJEvyWkfM8p4s/B0RUF/wcnGoZ8sxhofYlKrGDcdE69xJLzol
OHyMvVUxheeS17LRwGSyvLwp4O7oXss29OEbgxQXfwD5sGR1Zut4jZSCUqdZcx81
aBzUBpcq4SwB5GRiNDp969u/+scXV3N7Nu7hTehDsppG8hrzZEaz32HMe8QnSBpM
W/3wP5mje5wmvFsQ0iPY1Z2qFp7INjqluDNJh3ch93aDxb5quq53KQh+EKFcbtQy
PSg8V24Ni5rtJGtiNTTSkooqQQ1kjzh0ACgiuKpfk/3ew7EUUWZC5dIDSqroSV8U
/aoR7I1s+BmgkZ/JKzG3M5vRKyPCIblKupRX0G1Da4SgIMEFomL3fW68x6l7ymc7
SpZ8j46gnVSHMRiTquvxTuf7i/a9Hl+kDx3J4y1Cl9TurBtmAf59yTgkf6RNxslS
6Z3tPYFfWoAXsYi4iPLfkSog8WLVVeFUWt3WQdxHXFjjgY8KH9nHXsHUO4zKltNe
z6UixWNt836UFMNYbu7cNMe0/sApIaGfV0SPKR0UuZ4jalHwIkg8RnsYi7WPMiza
EdiKvgD2GmQwgrtFDgayoPQmZ3TsYQyg/fzH4RxYXpxuVl2bO0rNRfbH7IdQROHp
1UMbvF2BJhopxwy1d4D8A+CcflDk512TTq8aZJCF7nvgVabpQBCrFhsaNMRi7EAn
J2oIFxuUkhQIqB3c5UfFyfy6fq34hkCHjM++xWJX43ndMAHK8et2LIj0zSiz4oMJ
MDG5XHTU9ygWSvMweBjsj2HZYpwAoPuStwMoX8ZB5zNBMQH4jWncd1pWTsbdIgN/
mPCai71bZ0eK8Erb7HZVorFQDMuI4hkUUzk50HoYfT3aTjROal5GAWHQTt4zmdsk
vIXwQYMjEwu+HWiQFQjmHmIGqKSyQah/xS47/55tQlUj9ymqX1GB9MF+BFxNZEOO
X5LmmyX8GSEy3WP9LMNv09789J/tmAzgAlZWdpTi4Ow9Y2vQk7TyshTDMPVU084F
ee3LQEQypNAkIMVhVyJVI8wOIDTEPj8POYX/m6CdpezMsg1Isdb2LxTDYwJK9XGx
+QAH8AO6kJulPk3CHpj/UpVywcrZyb+O0pbGOpwXbRpKi4oTvq00PSidK2pbdwrm
6oQ07od23gK4rjjSc5nUfQDdpuMajsSQ/uvAu6WT6nZCHQlFrOYmy7IbXAjt074a
iS1+uswwp10LKha8APhNQ/dT6MFlKKTXWWkf1p3Jg9FCEZlP3NZ7C+x+A4KJXqw+
+xl4TjSdsNwoowK+uVMIBMrPzluzgp+7iIKYa+bzKnGXT36qR7E3Cvjq+55sIQDK
nd3ZOoPq5zg06KipapRg891jEbCVs/kfga33tvjeLEnQKydMgF5TjREvhY6I8FfY
jEHbVKU+5iDFF2PKpSgKePbWSru7hO3JWtBLiIVNLM0SlMt73RiXdOAK1dFldjuH
dVzhnw/DcWoeVxzqbpXesc1Ekmq3jSUt9zkT2ao6KgUqvQ0ScuDtB2lBFb1V7GGI
3u5vqixlylciJh8dcJatDP+RQxO+F3Sb4HG4ZqmAemhK89IGzkPb98rO6dBAh5Rr
jLlv2yEJog3z8ZyzF8XWQehL2MGcD7uvJItQ9qa1od6vZaTWJGivf/A0aSWKBHof
3ngaMCTvQs8knRSxeQysS8SU1J62NzqDPFhFzLfHjnO23OSIFulKuLSyzm3fCRTA
uOHB3B+7scnVp5OBPI3ej7OzRAmOdjKqRr4TQ/SdFkp1qJQWK1zDTVIiqtio1PJO
1sJ8iR4jgQ18NGVvKgjBtXuVH03CFv+qsT+swLoRfmfpgDPyOXB9/fobjvS+TJT7
2Xh0K87CpoUEki03FsMB3DSj3zj9TrqtQY1tr7/7EAGjnRm/6kFzBBI47IAob0QK
JW5s2B+Ku89ji1FZfxHsdIMMFJvJH0lOowBfucr3vfN7fYppXoJC81I9ZtTalWhy
q04K/EvVifLXzc9XFHSsWFbDgP+P1eT4k4x3p4GpPiuTfh9PrRs88oeXBnN+7OTv
noIuoXWssziiNY7cgRYWdcD64zJjxh45NRuw3PgSBRhsVX4oO/6puOFyLdv5avlk
Lj5ZHcVHhzAWncQYZql52Hc4UPIf7DKewiivuUTlxlUp/lmJ6ozoe9hccOsfjLw2
3AQxzIwveY3c66tj+r4Z/EWFGGst3L24gGJcyoc2HsepN0QgQS4bIH3WPPLqglmG
PbUBuoXHidf6shtcJz1II48i4L1Ni4+r0Qfcz58l/QbO/Bh4rn8kqZ6hzvi6OFAS
jhF5SElbOOHoXldW17vyWCLmP3nGK2g9FxWJb+CZGt7nV62xfg60PCs80ehKouWX
t3YMYmqWTJ/sUJXcQy0t3PWN5avKatx8Fdc61a0hEZwavKCFlYZbYPFG6JlMyIbl
tkAc99zuUTXuGJRYABXjN2iWLP/r0BetPiov1T53XDhn1uImJ06PfG6bf2Vy6pvJ
HO2QMyjaLW7pENPlGuXEyD7IUcYtihprbzHX6LD5jezNgboCw4THIcdgYeTMu36d
NR+gQJtc6QNakY6n1r9xUFs9cCGhOzFwNrRPO9SkAyZ8W9oVhr+EOLVq+xSKkzjx
9K23L9SOaRQiRSUBWFHZNg7hH7hs5u5MdwQ0QYaDRcqKOYEkEfkV10xPz6LvsLpE
IB3qRTye7xRyF88+cX+chIWiavhAUGI4vkoMbc65bLO9MFnXnK+TOy/BFDX0IZuy
WZC9flXRgoN0dTJ967FNnmR7lA7G/xtsqrBEWkQkoF4S3afqvw5kifNfIeYmuH+3
Yw1q94D1hkTGXWoT20aGE+Q8Wowfl9pEQlK/b9gCYsBYM11+6pIdlIQ2sZP5EeAo
m0950+mYcs6v1r4q1wlxlS1p/AvEMX8jHE8sNcvhubko2fUlofKa5slXN/3CkLWz
0k86Bj9qGwqqef+qT5as9J7HteYN1A8tIdObI+OFh3uhTwAZOLkIrG5zYKrVsnDg
7d67VMYRjqLUh+B8tzjRl+TfubIq/II966cFvDR5zRkYu35tlYRM5aiM0SJ2gcdG
0qFu3EEHtlzDipmu0KXsn4cSY00bH+bUBSHIFrq91y7YKOicCj6oylJOXEREOlq+
dCRXUk4xMlHoZ4+5EJ4VGF9mGTLfHxKUI0FUq3QiCelAQMSn+uzTDUC8aGJ8Zb+n
XJftvw/F9mI/WiBQ1Ka0BcdRfn4m8lGixi7ASMj43oab+D7IhIcD4wiSe3AZXDJ8
ugIpTjskdBpNcNfwovVy3NvOfLvY02jMd6I26+yl2LXM3PqsQ1YsXxrGBqS4mHxu
7a9S3+s0H3kB2Efg3veQL2c9Li6aX7/YFm1ZVfidxR3lSFtneuvReYrSkRCBi2ju
xEaJ8aSVEneqhDU1H1Fc8eZ83+S2ZObmdiiXS5ryBnShcE/ATQP7ojTkbaJQZKuy
HAYV5D8dJoNHdjhrjXSLetpqxvKhB2d0Oks8w3EIckcaN0E3Y5N5jScbwYiFiLjy
oBakVxmie1uwCiDJv8dtCTTv8YtxEJF3buGT+POJX4eriuz4hlbg8K37zYV44hCw
gC+k0l/MN0XJFL5DTc4KfNKm87aUxdmWMTpHCGHv0oR9py4Foq6gPO3Qp7DKsTvM
FKyyWkz9ouYWuWOtd7g/jTFCEHjgPDk1kng4kk/2mOALC+MwBz0gRh6c3MecvzsP
MCxg31bvBQ/FTUYyp21FlwkhYP0bU+mGQwSfaYmeQHhei13zH9cp22VhlsLrc/dv
NrszzzRD2c/JjSa31Clk68ldVrasZCD0uuE/G3yJ5JYG/1CIQ39FeVzLQi7mChn+
/SeNCSZy1o9jyUx9EfoCwGZXx0BwFxBvav/lVUx7DVG1Ype+JZALp7eIM2YJtK2V
oGy50sfoA0w7DQsKh601I87x0aTWrXQLZrNS9JmXZ+kCMJqcNZbqdwVyghXJFFg/
/toC55zPCqfKSwbkgEypaxKSvYwJduLF8TiAWK1sOI0H4isyHQ/WIF8IZjpHz3LK
kgJadrUO0WuEvLFtaF1R8+R6aL7DZmf3toi4SX+NvXp6UB9D4gaDGp5pd80Nst6I
zHkfZuyLBfZQdRprD/eLbVOPrBeERSN0kbNEoj8qQW1kt+jFxDbWqtpfOZfoAZjd
8PM2jbUXhhscbZYoA/n5zkMxTp3sCebSDc5T7qqXzi1FvozF1zUlyNwAMrjwf79W
8GySbupwe22S2MB3hoMCY7yoto9rXJZjBFPPKhs/hfDzBdagn9fyObdy1l0/Vl0i
/V8d5dSPHT9L/fSzfC9kuYT8xUn6VDkJY8z0CR5d6nG4M0vtqeOlONiVvc2qaLbh
q6DUr8qRIu1iUXklQtkl21tRPc43iuqgG4DdBpxAfYl4EgEqh27JOQWQNeQDbmVJ
ccMu1bWYUwEyUdXs/hFBOEfD9GvB8Aa8lLkZ7quD9ji+65a3s/B1Lizm0sKn6MYR
kT5b3LyJS0WYvquKwUt3wJv97whGQxu4GtWDLAtEmVvsFRU74KmTp50dg8689Phs
2b2Jne7NvDBejRHpG3S4fwB3zlEKA1YhgwXRHHnAMUg1VKYytp4ihOkfrb0Sdp6q
Z+MhdlOGnosHASg7Ra1DcNWscDQqpRs8IP6F/jJk6GhU8EuBxZfU4D1wLj5h68PM
Ma+fVBOI7qrWbP16KnW+0JFNtoOWmS5ivJnXFhcqtkGBeNl38jb6DJgG0t6ooly9
afLkNPU1Lp37NQROSuT4Fdwrsh/U/+LNBxh8Waa+YrYkKTpARB7YN/yuKIeo+Sa2
DRXAO+fC+vuMqrdZDg4WbrJhbnO11sKnYxx5Gcn+bwq0DZdUJE12PddNocfwkg3Z
sWtPDx9omEKYjoSaeoHYxhi0scrpuyNNNAwsl0YC3kCRQ92Bl8stvdACuIFDVtCF
fmhRaNaLUR7EfXT2a475Ek2diGdpLh90nM4ai9cPti7bI6LOAaif1ptlq0rk1bhO
BtDhXTTXqPs692yftNHppeTyy2uUSHszux9F/ZzLDnuV0hD7S1Oo2n1s4XoD4cK7
qMBFqLTXnyc7wtTiCB9hn2NkFzQ/GFD7uqE2KJYKNmiBCR93NdF1TuOS5OeFkq5w
/VwkeWp2FRQhTX9bm8JXQCBgdvEadKssfBE7Rne7xNgtAGCB+zaHygYe858M5jTm
WVS7H/UN2SPtssmryK3PoCrNwOzndwJxj/FlRYumuUQNCCz2uLAlfND+rKlAB2mK
uZQnQk8QcpnhdSPGoHXeCYnrwr3Gom8nmPM5JpGdFnD7K0EYaO+CiP1X7AdKPZyb
l/tTaicfjy0gRpSZpnOgbHbOaBTSVhpC8t2ziseOg5OLPy4Xa43rE+45teDxOpk0
AeCW8KZddoinkJlr2BrIDvfeTrHlcYXWTDWrf4tm2GYPg5BMEJWekJJGFC6yjE4k
SZzLkGwZx96kHnXrDW02VEacAvA8wPQ4sdcFzxx70JSVvAgl68Ezy2qfaUVcYxie
fJAxto71vJqPDRS4OZeVE50/FDSqVxYNlcaTM2qMA1ugLy0Igw9z752D6p+3Hf6v
LHzlbTqmbnC3J+0CfEg4EFTHr9cGm8Ff8NWhYKganWUKt5b8Qzl/VsWomlWPu0J5
N9MTw7LLMRcf5+yDAsdfBwrv8oaVm0S7ajtyAM5DJdrWly6VjFAGdI1O0k7A/KjP
XqTu64yXv4jqGmoQDJPeAuVys1Dn7iVV6WY48N0Du5wjOiKkOivBFMKcOt62WNEB
P0GguzXVrbophYe+JhzMfzH9SktlHr14WtQFvpInpY8Ha1M9iskdrLIy23BbkSFf
Oq3WYS8OGR8oiC96BMnNQCGCNg0b+JvM4ERp0VNor8/YkqMN4ZiZgujBqyqo/P+b
4dylH0qTxPCSnWFzI3V0+XPHrKxlEyfQp9RcWaQqA+aX5KuIk8Vbs8ZkabZQTRn3
awRbQLvO91C0G+D7kyID+nRzgr++mtpUT5snl3aAqxIiOWzwBjJv7xr/J1eAB22J
8uNtj1Wg0bkxkxGlOl15RPVa9xmfHMJT+uC3oHbCo9ZSlWqgjSZAjeH+kFxRmxBB
d0tqTVrY5WEVPCqpfyGrjO7EaoBb+oYPpoNjddktTv/PzRbqzas3HG9K75pjkmd4
lI9mi1yLJcIIpeK3QzgfoSLYAVxjyMZjkgzmrDHTbIWX1Ql1e0fLDbtAc7w2lyx4
u6vktF43PsNu3Es8VYJw0KD1X3YDXKmEA2kgzRZH4G3X+9ud42fQW+Ybf2OULaP2
BboMVgu1DLlHP5M+t6hK9WSe+MEutdQI4L3Puie5WcU8OrgZjBXGbpB4OfXhXGFR
NgF1qyXPPVVJ7ylL5chxseZPYM40aT0roVY6cPhNOG3UxlMfPaC1uTosIfv2yHeW
tKeZwopdaU0dQZ9p7L7zZbeOO6+IdfzDVBKLAGp4rScKg+CsihUGOCZMfAho2aFv
wVbJCInoiAR1+b09wOEk/GyX72Sq6JDXf5csvtKBLQz55lCSYWo+En3duqVPDIPm
2R+i9ILm/mcReBmlR2wR03cURu8V9aDQM7Ea1sowEKPyn6KqB7m8oKpyXLQjYzGi
E3HdCF0uJlc140sAPwa6AAg1CQoJOsRWzH5wX5ZGaqzClTUNDYwrwBxeq3w52uTJ
iZbtIue9aw0ZEpJOnj11Ytwu+xAaE+zGAtK6QBlk0lxxf30StRBUT0pMx1nKvFfc
SpjQc6oneGFgMQRaDc3Sh2LThsgYNec2meAxP7O1dYjT1mxwjejxnQrAH+hB7lgo
yK1zqhCSe0FhQDVXBZQpkWMsuzG4gX2tbdDnekwLjwsybu8MtPv5VBEb4rMZRfZF
FRrJXe6MXNRO2LXkjtV0gkrNFshLRAs+iFPoipW+nCit5iKTkUnL6bbejtkdbBfx
UsuktIWdGwa0cNroQqdKqMltP/EFNArHt6u9uYG7CipINo/HukmfhSsuEF547R8H
fB909cIDEzrHVmSd4Zuq56Jc5RB4MnDllrwRLa6TBoD5Lpj6Imw7eihrePwg4Mu/
BUqiuuFzYbFY4vEvvbpybm0f3fvMVY4gn4fAtebg1us0PvlYpipyz1yHzX8RzGhv
LX+bf9uOK2UFrsbCmfDsgHlcqgEfkIMpd4NtXtRoxPDq+paoeh5F4uMdlSZ57FsR
FRt06qQvji1EPtmmbSaFLkDrJK0n9VpDZlm4rMInNhjQZ2unKVTBUrFGbUMMdYyc
4rEPxuhdbGrKOeuIBh4SCfEY90bjocwieVk74nEaTFfbTRoegq0A6XylPsdFDX83
YXevAGswmqDB9g9bxBTPBUkqznFKbj5SgPgowHdo0NRVpU/CRPihiZadDs9g4weY
vjxeoxsnowlSgT+WWCoVtUKI/lEYaWPVEAXCXpePvyvoi5Sy1pq+ZXVf4x0WbrLu
p0HvNAzxstsXqKbi5i/kKSJGwUKUQ12TFVHmp00kck4mbOtWUiwFPfGmlIpQWOut
QbawAPXk2xqS9tKgC4Ke0MopzjngL4zAchQ+VmCRfDSa+EgrbtOXrs/O2pzyb5qx
LQgbqgS40XlKdD9xLeEEBHuDN7PUfA3ZPtk8g1SJba4D3Mb40A5rGWPytrIVMIoK
0efBF47SKL2MZysX4C8nygOzOeqjVmzzi6tTf1+nemycFAX6JhdVFR+q8RQziC3T
Undt9JTIbo+M8gImhTcbUwIF5Tk78mhC1ww8w8A/79fZPtHUL8HsbDzwHFdVrE3V
ZNrgY41Qanifq1NfEJ6Vb1d4xLGZo+OKad1lKLNb03Mkc+JIZcl82jdnGcIjI3SN
wBd1CsrWIcvInYjLblUJUtXFLKgoeaDUfp3Miixxb6LJefziAo1iaz76Z4MdrZoT
n0xqcTwoyhgADFqMYIJPwMc3yMu3O9W/ZOYo+kSzo3Oeh5dPJqbnGeQnxsQjXVoe
VdmBMlCrOUdNVine47HFQqZeSmh39qSAPOZWFaHzuom8Aextxwv2t5XKeQTODrIz
f2M7TxX8Xaszl+dk9o2cF4EmoQ5ysFpg8G5NbxYcg5v7/d3toJye8VPUd+RluAYQ
tQZ329mjGaLsIgwikqu09VH5QLvoxbSWeHvMYVtCYI5OMwkc6d5G1WRgO3w39IlS
0ksvEkw44Fqggm0cDnB0Ms5VDEShY1LGBiE8iViFt/4QuGSr4LFsL1SVamCIv29y
0lDeu1Gf+w4AeWcgCgRIANdvvCO1rhs15p7f2fM9nqjkA12RC/KBkvbFQou0lmZz
kUB62H5XPo677agGoAYlHytkZiUKZzFadjS8Q3FdD8w7EhyHDrAkzyZbPZ97rE6s
pVeAYALSYnFTM9FFSl24yZs2I3ZsltAwQjaP4GJpwxKj8puWWm+GYA/UOx6vdJa5
Ju90O9GWBSiaDi2ZYGFLW1xpBp9tOEF4P0P8QILSliS1NQGHfRf1I6EmmH7qCeeE
pLa9RmWM0zwjdvuk59Z15BNteWMxet58UT8tBOhvVkOnnLBTLuaIdJPRovAF0tvv
x4LyPuPeTy9fWG1r5AsOv37nACt8pxdzL6qe6lNg7S+z/GMfJ9XFWW8MM7qUlQeK
72HyUgqw3PdKWVLeI86FqWIsU9eXMxBabU6k8ZiOsS3G+9nkXC0hm7vN2n/tZuCi
XOAsUQYpQ51jNsyprqgcp888QCCRg/IznyxTglP4WNiBcnbfaElUMNaTo9cMA7Fb
HDEuK3S03D5a2FgCd/a8RS8CLwGSI4iGWqoftrwPNN5dUEnpubTEXPcJnh8NBK/m
S1hCyqWHkWenIduIZrpXDB22Y+mPWsd6xSK/ansvw68gDLm8Wk08H3CasT5XokDN
Bw4zaWOZTg73DoF53iIYGy1Bsahej8KMGHYQHKCtKCyHIo/L1AbADCTDDXtIGef5
HLM9V8QrADYFjc5f9xit2Nw0djtNYH1W+tABZndemVz9iuZITDQdv9LEdlZUbaqx
/OXFg3zEwdh//OJJJLxdNyC3/jOeuhBJAhpX0nLRSvKq2e2L8ET+uV4sIum52SCL
BkD8mgujg6K8nnRjV74j5ri5bR8gCYX9Rw0tWmOMKoykydZ9ZMEN5JVy3Koh5qCY
byWDqlCa9yn2Q/HGKqTH9pXGuFL6eFqoABqacrgn/jznUgQTu3eJmmUzMmRSQ7nu
6QGVXZg6kqHgK5hUEan7V30QSMHcHeghX7LG4fpkde2ACU3QVJSZXIl9SgKAD9px
KYTOqIkwHXzNG517zVhzYDYMXqcqXWvk0qJfDzMoLmgKsnoe1XpbmHHyWBkV7jn6
gHrM3lXs4s81DsSfO3ATicg8t31c7q7XmyZVSdc4c7zl6WN5eCrjOAGdW2Ul/hSC
NWt1ST1r5cw5nphqwxDNpPtuTktsUDsKcFlI4/dHMjwGRgnPYenAPagCbi9mr6+t
5sDzBMEYWNTgkk/NUC8FVBm88NgADyCj8NXX4oKhdFLdlXuINPsNc43Oq1Hf6G5z
eI0qdiRXJgX0bpZhteuzpS0Dw86GyRWgdlULEqHMkMk222Rw2/IHwAIuHoeiiXJP
y5kgkuiQ/RHV7Olqo/u2WlUsfHJiVTGMJHLb5MP2i47zQBowUsM2hgMvd31ZIOJ9
Mtn4+h6irXC/hlQEumbdSyO8feMmJeaqJN8OkXi93n+v644ZW1e+dG0hpLz4MswH
/otAjf437xpAuYiUjNvwp6IEcfCYP3pRheZ+AOWQjJ0LbNb1qjQjJByHnpRXdryV
7tfatjAYT0tatPwiCTNUeJuCPs7Uy8Xv4/hzoHy9y1Crkpmfobi//JG1cK2F7Gzj
y/RLLWdM3tlaREZGRzFX+AdDjnuAecO7llvM1IqfQfqsYs9U8t4F89WC+jNhts8b
vGqwqlu+mSpsT3q0tUKS4e9Wl8/cN7et4Q9Cv87MOFxABVBcM0nQE6YqtxSaue9C
9upM1Y2QZfxXKmzS3Ld5SPBrV9/EfSURiP3Cw35TA9kkWndvf7yVojMph1MeNJVN
n9GjzACLPjturx01T0INL0n1KU8niy0VaihCS4tdEjB3FbIGkkphw4SatoDd1Ymu
rXkG0Kkn4eFbyoGbAupO56Z2FSQPmpQqHtdGK4bJaM8sSljeT2jgVhlQzc92vha9
LUADTZcGVQmGUxq91k7aDHVdSAWWmnTJHJ/hWZnu1mo4o8K+cm5F5hB+0H5RFkB0
brZmIsQX6DMMnA/ZVeW6SLAsPvAenExWHn//evbkwAyoFGytpZ2mUosk3LjQ6eOb
u3+fiCW/7YUvIn0N+5AcD9ZPJNFVE9xLgxuQVh6ws0EV70e4/KeEd1znFhL/xMVd
MAVzCfjAR8K46ucXUW5SX583tRkvxivVgU+GXWdmwaeTmxWkZTA6WP+munH3WAI9
ZaoeWa4JO9TesvpXpqQ8T7GRlrPMZujwCeJTAw5NpMBH/qSNKov7xCrRDKBt0aSj
BY3wUB2TeE/+2LZLg0QydB87J1mFc8EBBvCAGEshsW3qhdozDXXahk6PWvEkvXgL
Upo2rt8h/olEzxNwBZ5L0jbl5Xj6HRUggJMmEye0lrZTvfKOAdMMW/SgoUIQkVo4
onWP2FgiuuodwEflAwXkmxP9uqS0Skhy0W4zz+b3VhHd3a/M5vzMkDZlW7ko7C1D
FHNyiHoTF5lCzoszuddklmmOlFNB9aQv8OvrG93PjjwoG/rXScMSRmemvYuVtXsb
QDQ0VeaNp1qLSDATKKULVtW6Eih/YLkmim5LGTs5qJ5P141Lg0FaVJ0Otg+cV8wx
WfrxcoGkUsQeGjUANWK950QplvDXD0cD9gf1cuJ201iqErEDGRGnQJgN3AcCpyEd
Ajhf1crfQP8f0J+MBdGArunno4/i/i6mKvvG5/JOREGZRGBJnlLdmB7Y+ubFODHI
NezIbZ7MLJk8InJBOR/AsRCKR/JG7064xtwp7YKUYG481FJ1Qzi4sY+jwEAkdHv3
Cy+BIZMHeP9lvVT3kfstZnQAEgQMEkE/2JdSbbelXrv3ow0beBI2Ke5QCQ5BZVkP
UdciBK5b9KzgkEUfkrTlihR0PF1MRD4FLfjmW/yGTip3trB029Otl+t5RWxMdlZ0
yk1P1c7wjH4HxezoET40y6qlL/mW1dW3PFW9yWJKHp8aHkPgK6eVuGZy6b+kiPSA
RZUtA14kbXfBF6R3SiYG4gHhHNozM9tSInKp5b0A8sDqyoBqXAmP6HUnEYbmrV9n
w+eq2yTzwwxgmuMzy/gPCnfFcINfvvpwDqS1Vxno8RFk8XVpzAuot7knkU4/dB8g
pas6cGu5vv/aRk7gvxYGZZT5JaF17bcvrMu9XaM4GuuaMFMu0+aa3dNbnVSnoCLU
LcsKucwZMm5XE31lT+H9dhtwT6/XxWWiwBxdRgIBs2GBHm86jgAZHuJERkz6UnKs
xgw9nQyiXBoF+uxzXO8ey1lrZUUvSat+6oqWEjv3ZpwnB5gJqDNFIJA2xeHWfOEC
s4Q8I+/YrT4rlJMlRzyju57XGbF4THeEJLtaGLBWuCniuJo3daOBe4G78jLEaQOV
Z2LqvsjA9OEdBQcqpsTs7cwyxo/zW7SapNjaRdZ+cfCoEXUAokqqDG/TvP+1xSRK
/aMR/JoSsm64osIHQkq0CHqhnD8npXbF4eb62ZF3QTjqAtaYh1q9ZtlROqlPFv5I
QFFVMhYPeSHGki0jaBkhE2CwA2RnxwWMqWhv5WWwGkZBsB3xL6BaVDxNXcm0SG7F
rsSzKaMNT8NHTcGGPyRTugOuQXXaAfaB7wUTGNHUXADDcReeybBsjUcHiFYn8XZj
OtVZwf6pCTvU5+ZmIWwDNFHOTuPt1G2mq+/aAQ4ejDTw8PKOioX+bD7vReQZ+9Bq
LGo3ZG+jNOBzsWPouM6rqoUy5zU/dwZKaQzKA0gKgLN+HRH8piU2JxDsRX/wpNWz
40ENEbpAyRI9o7rdd0Sm7H6g02++Clhl8vZpAOfwqxpo6M2TwxUBI8vHISsWEfKe
4FjqAgJ2YbwZF44/TfsPqU9Q621iLQe2V0pe4AyjKalTbwRJa5V714h26xIIAVvl
hpNtKj04qi9D/ivbEnZAzeP1EJqb24c9h4jfgGivXFushjBOOF7Sy9jsQ5/TsfbD
fLd84O3lp1j/Zn9jjwDCUxY4r3BUo6Y5JvtkOeKuuig1Pr77VKWBiENAoNy8rk61
a+gB5Txsl4IqAZQ4UvQjRDW+aD+BPVOkDrHr9zjulLvbKY8n1ihfu/qYIM57uytI
JWA5vEJriecOONiOYr18BlpkjTNvIsA0sbXSzQgpwxdtOfVeATDMAE8bVcbXuI/X
fW8N2g50Ayah2acVx9Jre08rMusEZuJMlui0+XbC8pKwBKf9am8LM4iA1+vbBLzV
gb7SwRNisRkpVqBC91HQlMRf3We6kdE2MrJKuYUOkOo71oWw96Crpx5tionZ5ksp
RwLGXg23DTk4kx8QI0F14Z9Gj2YOaGo9TojSjWaS6wGrbWI3TJHeVwHqWYwVUkjU
0hM+XoK/jV18Hozefh+6fAjlL66JYkKTBtLoaOOdHpEvEq+Va+excmqkM8RKQqhW
90r7Fga4Jy2jkO4P7OnJg5y+ft3zKZQZC6mfvRK+5g9V5skHSv9bw/queAwW6ulF
sOH5qm/bZwtyFhf2Wr59w6j9+lgB4IzzmIDx1LH8BIqaY69iBQYuIepJG8o1lDtF
pgv1yJO3dpTzkvuj4k15Q43zxdVDprKw1kal+zfuoUmzEo9zhw+D5OIXBmrCyeDF
+iN0GOUraIUDYqotbxpXrPEIu8Miu07Mxv5lHHVgcU4pcJzVYiKDH6j57HEYOhT9
48/eJlv2JGfA7Ycr+zNuzdkCUhzseJSIPS39D7ZCIFkAn0rp10VAC06ksGaOaiB4
DpPbjemOgEjHgdSeg+mwE55J2mYX562Q4olTBbb5unNj+zWc6czYUh+Wvh4FkKpB
9ruVQaPh9nrkhT/P42JzhFznhttpJo7t6yRRxG8SdxM0OstPdZSobYRxdOHpGi57
gZWP03nmR1QRwgj+gGOS9+CtkgaHzpXcX8i+DciOeFhJtiW8eWddha0NO7l8Len6
QPgod6/ijV+5zE1/UbiulyVEwFf6w70mzPEG6V5//GLQYyWrKoM/6Zn7czoWp4UO
/6qEe3hNK0ifZrrAclu80AIHFlWLrkPTvgC7SnOqu70wJX/qnI5v6lipEe00GHrM
mx/tiq24CVpiqNMcVgtgVMzMnnldsZajL1F6qeInZtQMNQssuaOOgEMBYUe+1FHX
hRP5VaSUPQrlRUHKR1dENu6IUtcbFC9nZFABM5iJx/rCxFBXKokMVc4OiLkwM1HN
rr7KlYsoRHK22r8mW/tctRScOqsLIm++u67NmmdzYVvYf4l9KaytZ4CWNLDMU4Km
vmffogO5QpI4xxNJyW7OOqFeQNFFFZYmHaZuIV/ugLD4pKriLA/Yk8/3HtFM6wb5
lvR75Z3Y2nXJZ9XVVLznf8nc8CdBWW9lxC2Hk8+grcHWPfYz+kTVjRGTHLI34o2P
g6O6hOBhz580dAcKPURd9iQtc5YYvtBzoTlDfQjhuuCDLUFQXCsvaZXjLt4Go+Lq
1ld8mvZz9X1QkEcbc+YPGCNPn9T9RjHISsGEJGUrNs0Sv7IZvtmvXCesme6KE0aV
vi8I8THvR5vXxDU0e0zuRl2XCmrzMXMlm2MlFioE7d6fk5olU7D3IoDGGWL2HB2i
VP5f74rfEiQ3CxCaMYcZZM0vU8oqRDnYNCxKFsgWc4c68owhWIN/PEbpssyYb+WS
577lPTDDpN3AUpmJwxAQG1FVZGB2cy/ehrFOQgBCVLgQ/blcdzgWBFyjfWlF8O40
/XAh4nOT8elsj/qlsUMsiGgziUs7Ud/VYVPwqoH5AdkcTsPjL1g+dTcWtHpT4jOU
rhRWpARN53MTQFRmkaAnKgiWOw+3Ufx9Y5cL+a65y8EfiWlSMuZstdqjVLDjsqFU
CYLOzpEMxT/GAeAYToXAbz2PyuWjDikClwAwuCC/NBsAqihjxRWNBlN2D5pWkXOl
Ae4YoWHdbw27EpvUbTnD+klZoGBJYoUatLzpeo01wuH/twY/mnUEYlYODTTaTpd7
f20kMlf3RffN7bC8fVt8F2EcAmUGUSADeaFFzcWWoB7JznR8xx7EBAyNEjS54Ndn
okRdcRRurcuFrG8OCuuqO96FTW7KWN4xIDmnW+aCyhEuPpROqk9WzFIxQ3lKeZ6q
y0d53ywTNaxLSx+xoZCO0w5h8A4lMBbYcUer5+IlQRPdLwzWYGjcu496gfyZ1smn
kYYTOsPUTQtd/w+q7ZwdvaS97JVV3gFbkVvbtRceRs2VmcLifsVFiywLpes3IIUA
i6O1Fhju7alIpYV57jbHV0GbjQAb9Aue2DlK4ItcxgOqA2lo71QpXSmscdzzBwaM
NIoyhfsSeT3XKokXLl1cIpNMB/OeqHp81QrryC8pgQ6abq+I/IY02pqrt/2pgohN
aTmV384zwLAOhZmfPFaw0S/fFZoe0iRBkyEW0hNH49jiDAQbWNJfSmEjA9C1Q39q
0QnL+jbKRQ494tEdausxtoQej1ZwM6lV8IQHDzbYfzjgreGeC6RCedb/jiF/pVEJ
TwoDAQQRbzTGsoh1OO6pkpG571f5qVexwCuakFLT2PNufl1/1MPDFU6FaCZBgTqO
04zTutG0LFAKDezXyEXD9hsSP47P9T9H/0cOzSQYKETXhXPE4M+xCq8owDtoxWon
XZU0lYWp5SU+/GISHyIX47A/YmJK3hdacPV/fl/2SkW6zIFAQNpHKdZv4mkALZ2L
i+S/lIZEd6NA22xHKUUdIrHph1ZymeU2J+EUIGDR9jhPBU7zaVMA3uxvTVq2487D
by+gEwwZL7a22NIGQeJ6AQ1gKm3BEV06bg8Y36t25ALvNTSwn4aGFxlNDP6jO2nd
2AjVHHj2uKoVeBEj+T7dRzzveDxEPNGvTsxdaq3S8tEusCfVnnzyx2dA//8I3OiV
23cMa0QftZFr+wASj6qeOaE0WMi5k8hRJAPi5qiDCifMSugxfyjfDRD88NiIZbUi
wa4rWABNo7nv2mhpaIZU/5/uStbUhIiewPqB11QPombQC6DTGPKiyPGfocQ39End
le0Cy/gWSe6TERGr5v3AyuSYDzrKzAB8OPjOZztdJg2sTAy0HUpwheYRjkbdJMkj
VyhH/bZaecSsqZKQav1/PWhPeGIe+2j5J9xf08uZHd1/skgZy/oVplvF+0+c14eG
KZ96CM6NAgcAQ9xeMEAj8sp34tQl/Gy850FZNjv7GnvxjxPWq6T3BLaTHiw6CUwz
arz5qohsJwwSSsMxr//NvO6DC0lrhwk/jOljFc+igdF7cyhHK7Z4HAeGILVhBIuJ
Yf2F12pQpOkuaqGAwh+tnY/bS4IPJnLIoqHM8fLQJQ+Wv0JK7SOBd+BcCIthP3+L
jrmhwIsOQGSeQITcEyzzTHpa9UiW56i7cSNlBHFlWxIwsomXtUn7zqtbKafwTMYB
IHIb5CwW+cs33ElWQN2YNxY9xx7mYZLjT6vYGXPriIIScCz++KRh1DGG6xpaQjN5
wchcWs1qmKhoA747ZTsm7/rxIsEmN2jc9+roPUxwzgFFzfCwopgXBkaWvMXkEa4w
dptDhWw8iWVe7k1v0cQx2Gt06xnYJLWfkplCGqy6yiA8Oil7XKd4jrymxmuakb1X
DCrpJknrGt0GGSqMW4g5Tke4XzGRlA/j2IJ+bE+kAVA4NYiQQsQYZ0z3tLhMBSDM
UQY+2CAPXzXxktgTANkwKvuhemVVrvoZ+3FnVMOXOBg15Db68WuzgPX0GG+UCSht
re+WP24miYPGvh+3B+tlDN4DgA65laEyD46/Oon+piqmMSjk5jxLws9IKgMz1A37
5/r9d4c8h7AOtrmcoLZq6LosLEfVdAoqyfbxYVcVLPAA3uL4bhniYKYX4yBNRSCU
LNx7ZwSz10D+WwBF8Oohh3ob4noyGogYWN+nE9LD5F1hen89VLrGLh3Fl3kpBcaC
aX6Z3TtysjMi+sl7Q/78G4P8isUcxGBlVXsyu/HcBsVsIEs15Ocr53MIG6FjxokI
pEKZ6mDK4lUqWYMgexbptS4LSLmD5oAHPQ88ijnPUFoX0b4cYg5FxO5BdiUsp2iA
3lv3lTML0/nq8suYgboJc9at+HH1sezN2U0dzh8bQQb7ePk0nGvnRLk+sTGw6fJG
/LhVV3R8bYOE2wNE4ygD5rY9CMZ5o3GL41OBOy/PiHQFUo18ZQBwWhjDzmVbtGGF
+ljMRGClCQEKXj9XQPHptxORu3zXhbSqA1Y0dxFRe9QdX6o79ChdYH/Zx/QsmtE5
i2BZQTRy3p7KYwDSDjAYBQLgOekaTvCOcYVXws5nAlh0a7O/0byLueO5ZmsV0BuQ
46Ef2PJP538aCvdQITVAlxnxrPBJeQqkCjfJ+ixRxfLuTUhSbrTwBptn0C0ZEvhO
hOVmRVye7bQzJWMMHMwab21REtJ3xSlm2dNwySFpeDHq98Y+w2riLsMlJuvDfok+
y2deLQCXwvKgeG0elk/4rxM6rQCbKPei61+rq0aUmJBakgsskmCAq5njM98wH6dJ
qUrjsqojzIqNXffLn3DWfJQVqhJnVQXYiNiDDUFKoI7K4OU06RrCFAztAhEhpTsV
to9yY+vz1IUhgrPkxzUDnTdOlgdsXnOxoSxhwHuvGjgE5ZCzdp/e4laExjop00Xr
ukjKGH0/u5TZlfd6N05FDwy6JLkZg5wj6DjktW9g2AqIiK6feWpLJejH8qpCC7Qo
aG0JQuDyIZG4XkImijE4LAanWnRuflfCne2KgVMAltrlvTlcsArEcjHyI+kWI5VY
lOYHSsSLzdiVWJAOoxR2wIVQYmNus0gCPKjR3Mr+zR6Du8jegRPvOBdwg4gsCcEw
EEEkLWNcHIucF1kKfkE33q6hW+wLBGswXXLGfCvhi9ViNQrGZnW83cIIvhtBL3ra
zbfUkXTTKGP4oLKt/uSljHNovMrdvIT2C01xlJvYpWDMZjiAWWBWU57uVC7EI2kW
pDQf9sXg11e46uDXzjcu9S19cqTF67CvYxuGFVMoINvgcLwKdhF4s43z2qn+KFGC
4SLwQ1i5m3QXa19xvmgXWvBJQQkeM45nIIriIWd+TFr8dgs1KsbOe7wT1kq65wA2
3+NCdFhfB2LM9KWH2wXCdBNZ46QESGeCgL7iPSWTBGoEZ2fsCvtXyVkfjq6RQWRV
2R3D6vq6iwi3n8JY0Dawvoi/QoCuFYiuvKJi0TOBFq4ygSVQBd8wiRrhtWiriT9m
I2wswc1THuLX5FJbQjD68DjpKGE/vOFRWewpNjWxnu4kz7SJQ8mOBTi22yTwNNM+
LxwkvV3B+hNjY/YTEgLemzrRi3cI0P2XU2e5eX8e2B1sfads3TE0bBRaw57E5EnF
ji3eK4wTfOD6vsImTN3XM0cV59u2W24TZkXT19D0Kas4eC6QQuq8sfpXwburw+Ab
m7CQlwssPQJJ/w6XuBHlBikFPtxZVdVxhrzNMlQ4oEaF47DHw+4Y+5A8MC8i4ByT
vZUtwHXoy08P4xZBZaB4rQaDLEVjzwBzB6NE/jgbAjIVOyyh5R2A8BOVUtBB/PuG
7NpjLgXNcLQ9rfDppeUfxOWU4Wck+F4hpOWUW7cGXqVmi7vzDoUd6VsVSFnNkEE/
FvOJ2qWDl9M2v9zkx9qwQCoCp0FW2IRo72YgGSOAI/dHHvv/+l9IRWQf6TcpwFgp
OlIpVonkqqB+/loG742dlwv3CFEnWCqu/FvtK0vVGZ+idRawpOwSYju5YfS8L7go
RCvDuGbww6/ew+sskkLNxLTUGjwcf1jYSANechffVpgCSRAOyX8qx0yXqqZmSJUR
JAcAaui8Z/ti+ynMNJ96zIWTAYeeBtmirUelgXIVIrbhorHKfT79Mv823GjnrTvS
OpyD7DVQxab6pCceOXm+sxUXmJY886abn+DTj1P+LVl1HNSgET8BTDlNkIL3zaPV
TEjWxNgM0WGdVWxBuz0XgMBWzUfuHHibQ56ZfWoqg+OiMrbfzfsbyzbp9FG3NY2n
UVO+d3wL15GEQRkfd97M4RzW4smYFw5gnzRPzNHEkdrKCB1E78BXCUtgl1rAORWd
+9CkNPxzCXOhtS/gOZBiXv86Rw9Wg8+7W2eOE5ODX1tIyfh9ZR7FEktdxwlMVGTS
StDSInifFLMLuiOhSHos1cctNH79WJ5iVS5r6rhgiYJaTHKbZwAwE1SZ62Jh7W19
Hi1BUxCS4wZdyYdqFMCGfKxhP6cZ6Lg/Zmtf21V3l61ZnO6w3cY8AngjXZwt67AB
QLuKm0mOZXZGHl/BmXRa0QCLljoctFKn+30rBJYpO+r5MDRJW0i5utddTCXE1Fsh
rRlISALDZcSScPKfpg6Yc20tREChQ3HJviHRnK5rP+bO1h+knT7h34T4akJ/FA3w
JQIV3RSt6Nb7HAE6BkGpoSYPjY2ocPf9Ak8LUhKDwOCIFWP5YLK7DDR9VwC1z+0y
eZx856L1Rpf7dNOcUBgO/K9iw8w7TSgAhTV2oOHyopkkfZ5LHaY5JD6yG1Q9+Sni
amrn/VvnJm70JgeQyQ2GGEr0xjGzwlhOI5nqXL8uYDaFMSCAPGrdQi9kVXYp5KIl
TH/m2AjcsYaWjUTJrZ1SjplvBIBC/bs7rRnjr+uwBI2CFduy1f56ZRQNRjrwT925
fLx5DgokgaiuTKtxziWJr/L4esxQ4lzfTsMGEWET2DgL2ZgNlXcSopWksvRrPoi+
bJdkG4B6YlILeWDmO4zkmOr3D6ToeHsIGEnUYwX7vlA7iNRSb4R5JyxObyWr+JVM
D4sNXfb7IS16VMj8Evde42lZ74HICuViKFFIeFl/ciimO9nC0M623QjYRZm71vcY
3oxj76SsP21shjMUXKBWuyZbVPKGq2IH8YIC1j/+pXiMhaQQrMicQZcqq9nChd1c
L68ORanfhD88zFGPkt77NbC9Suu5xwMk2VtRCHf7K7r74E3DsmQrfalWDxtm56sr
KiPv8ccGCI7NpVmpID9wNMNQWG/hweeUqFpbTFEUEALEosTkcFv7q/8qjw3STdfl
oyp4rumvxcgNunEM6nxWKmpf9DSxjTxUwmgo+F9nUlZPnvO+v3bxygcMKfYw9ZA9
aDul+r0A6bksPgGHMxwNPdnvEkdL0/S4S8HkwEjZy4Jyhf5u5cOMWAF+w53kiCTU
QGK/5XhWzUNmt2qkrSyAd/aW0LDVAzrh0qB9ymQciObBlWids5mWSzluOyILKEzH
/c9PGrOb2ZkdM01YDgUS1rD28vXafTaRdOnagPlwBo7HVEZrJX8FyqStUKkj8RYc
llWUYSaWLRYhwwc/OlaZpnTHMqyFR7hwdwLSywv58FoncRbAPKEZH8HQhnt5LXrS
ly3N3JbpUlvQb+A4B+RvT7O4UQAaJMk5/k8a3uVN7GWy9AroLEh2+JREdD+HlICI
xwMtMP2697s2dy3Uc428NyDYIjY3nY/sCGVuL7IvM6/jz2qUTBG1iZxvX+WlXDZ5
MTBB/Xy+ppQoZkTHgaf5wM+pXXHg8St/C5mFqc0WBY8+Ld3zIFjI/nt3imZnaxET
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36768 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
vWaiee8LnCgatAmbQJm76A/zGAebyhAD3IioT3Faw79BUTiCXpEnqRloS2SjZH1N
oZ45qhisfAZsnvtpRmNhd4qAFMlrHVezE8Jx9DpTulQiLuehDgBxJYx3BT35WKz3
kahxRaRau2oEmWbGOwXV+BeDZJCGelL54drjcM5xv4toVaUF1EQrETos5/bcBU1B
1jGhicgiKs4Lm30Dkly157AgST9A5HBTsW/qWft3+NI8wyvpnk80dSeyGAyN5lvv
o05dojjU1cnixf9VMDlHSPF6Lx/JS4rDG1T9MhgvYx1YnzXuQlfWWYGZ1xBKqZc0
6A6hv5rjNCzOOLasM95/TiSuFTQjiflIGXmT+2hHEBoUYfueDOtMrjqEf8mkpYTM
bQbGoAzBPYoZPoE5fuHkY/Nkan8ylSHX2Gnbh/LjIn/f6o1H06oy3W/bZ3CklPNO
SScINmtMafqENvUZdXVyZaKJSUhP8Ca5BaLvJG2UC10+qQnI5tKyIx+85N+UciGp
kPDIjoZFue8ICRSItTAad60JLm5uGr73eovgh5U495TQDfic7yyOQ2ry0q54ACjf
ZqlX3sMzUaWn8erKK4UkKiIoo64VXJ8gom2kP0slGpyQACYUkUAAbOngFFGSAoqt
biNjou3PPW7ec8tFrMBZDz/7AD/zyZ4dVmqxRypmIZ8xu+gC0OKArp5vJLv5EjqD
dd4NCqAWEpbJRHDFWVrFRdemEtyqupf6Yr3/SxUCPyferF4o/rzAWl7QzkVBbqsv
B2ul8NLIOMZyyUu7zP4D38wXCZXwElIfoPyVslNHtX9YsHIosTIH4p/PcqQd/ojl
4nOkMCP/tnK1QNuIw12mKwtCUnB/PKH03w//mrKKQxA+S0FbB1E/p5E1gRFhxU5t
cR3gUm+cOEDoIIkHP8Tghf4wWNG+/QsS3FUIDqV9s+z+gnwOLjMqYEurXlKd44PO
9vo54W9iaa66btmhTZsgDb+yHOxd5+3aV97dVM93sKiES/odGeeK4naYnZ1x0J6o
2bM/Q3n00bHR3EEjL9lVLd6xQycULUJrdfDlhJJbBwPPjwMbBT4ZAgDd8jh6sMGl
SGNhn95eCh0UASWwf/C/1lxKy2BhULwMpDo4jGzZHtAezJRtT50KXv1EbLmklYMf
FJHNo4SfPFSLJgYa7AkOgABqHDEsjfYgLwnIH9ZnedrkmtgV6EBITmrTfsTZgPcF
zUl8XL+Acin/AiHypjSUnf8Ng2V84X503qHW77iqRDzJIUlH5RzVM2Ri4RPi5euD
Trqk2JamdRgRa0XrxLGgej/hW17uTNSO4bQqXNdL/uS35+LW1+mP1aYkKYaxNC5e
KOf5qx/s7w0GVX8rke/OGDIEwkhNSnj/i5RS+xmzchHs1pUCt5Ng33QyPPQPinGh
4kIl6s+M0VPQD7Rm1yq4rch9tVoHDqBbOpzlEm7zDHWGg5qxJuWXHx87pW7Zpn6z
jqwzUadTTHZ1WqKfbws9BA8JlGKGZjK+++Wtl0Ucxq7FQlbmYy1OloeWIHudT9MD
8BF3pZJUaz6VOm+9zLwGraMNPCsA2HN6Z3qPJvIKS6QBcV4hFiHSEXsHMvpHg+g+
djb2+SyEev9EN7Gp57RMtcWMzRUwP+Xqv9doljV4mXiWHWFWTxSWfAH1DnZjXIHf
TU/84iNMVdm5HKHzwsi64iY7bUp/I6X7zAiHbTwPj7WTHnrrL55fKwmvqAA3RkZA
Xc+RGkHo0dDvtNN6hReeHaYjtdu0wIOntS0TcTQoRukyWmyFKs4Yr23d3XiX3zTW
5b5IqiKifH03rGdB5hqSkKwapo6x7cQPq/9X9eAx53XwbfwFyZyg+oD/tj2QN55T
MTLKZg7UqCfIM+G/QlYfbn9b6pYuiHcb+SdtieIHv2Y7YBPvAOTqHzbIlAfdP+4N
6jwH7hF4aXMArZTQC3VxKRLSAfXI+6gdH7aCuFFebpW/+mJBUP26b8Jf7zZNdjzD
zZGBrO4S4q0XwZpWzrYxXkckdoHhCOb81XMxqqwsBnTwUpdLNGKLBcLfYlRX+7c5
Jq/x2mw6Szu5ymnrCSXOQQDSI/ZhOhgkeUPR4Z5P5OFmbwvGlRvAIjwndbIQZvYR
Y0yQjbuS8sxMryjI4UIJPUwltJrDc+/DWwiYCHNOyP7ls+gXjGelUtBwjoZER5Hp
HMBscrbaiAkiTPHnZnic+rIj5EyZUITnZCQvZPwsnnMOMp791HweE18UiRiMoFxW
4g00wOOE9cAytCnOn4hWmkFKwyKQ1Eeg8MXuL/G61Hgd0Fnyan3LB3ZDsonF5Y/i
PUimhPzxUNUtTwuT/656uBoRjqp6wPzxn51ww8jT8qGClh/4GMEA9yBT3sektuJG
BmdFPdsbpm3nFTqkeNN5PNbMXN5Af8sNoCkzgah1TdYy1qsq/IAcKZo2UUVzT+nr
lwE0wEJnSTupA32PvO6JalMcaMYsBTBpgZ71AzE2uaBqxp6Ydn2RJWID9gIfa5wi
uohsBRWUhYAjPNS3/osQBg5dA66yqGx6k9pFfQZEaFjvKeaOtMOOL/8z1DnQ00HH
TrfXTFK2RpOdCh2meb4HWYXXV1thXb6schdMy6yY6bGSpgLA/K+gtR1oIt77/y4t
yjjle4gWMkBCYJRpe+UhYawhxxokA6LNI0V6VDmby599Kf1XlX6t5RldK+00XwMN
KY1VjN9a9EnzzXES6qoIs6ZmFtTjKV+YBUQhTep4FTBJgnzA2zZsTO/RiVCRhZ+6
i0DZc/LC+/9BteaYdwz7SU2K8mjEYEwDvwYfhKAiN83kATVM4mv4ho6OG/xJhTdE
jD1mas8+Z+oAWBhbjA2l5mv98rmAfSD1+rVzmxyNmA0s7iQ06R3A3JNyyDjOdIG3
8aFISdRNQ7PmRh6z6yga9I8nYQrrcGsY6+HJo4zltesfgqHQImyjMhrv3Qqzz9tf
+stp5u7hkeS+NHMyMDPFq0CsIO5meoX/ZuaO5CmV+37CqOdv+u953mpZY54yJigq
RX803qd9PEvOX/7Q9LXJ1iePme3wQt0SU6GbDl1QpCMBybViScZDKC8tOyKQCE+i
f7urfMPQnk+44MY92iedt5wgVXLc/irajsRA7lDItKrU8+rny3LJDdSoWvGomLEO
ZT4/hGftY2YQQmz0mXaS/h4fU0Gl+fd139YVgW7vB+V5gHp3EZnwE0qitDN7eKnE
MOOzI61y9kZBm78t4pSbC8jeNVdaUR/x+sV8GwUJWPvedkf3cr3tcTmm788PQssL
a4NmeQoappWyEZHkrKx62Yr/MvGd1ikckkZsR0ET6Q6zTriLmx/gpwz/kSx4+QpT
4cDihaYHHEBoCKDVhclIvD8FaaQKVHcXww+6IwxfDMCVmDAnRz+dzHwRiD8X5iWT
0eyDGMfx+VbWN2XDm7BQRZmQ3iIDbK7WFwsF3+2S56c6nKFLU+pu4w/lJ279NHsi
PaFoZA/BTxcUwBEea42/iM2kUq59sgnk1TbO9qRAEKAt5/HfS8+OR0OALcYkDguc
l0e/5oOhJ0aIR1Vs3R5CkGYyOWM7Z07IFDQdSDEidezxt45u9SCYdUolAnwvkjUq
s7MDiiKMHB99Nzn2QBDnk8FOA+ntht7wa7QN+scvDDcEWxGWZf2doL/BZSNTJDen
utNWvEQNsZ3BgyQRNC+SpmDEyP5lJhtZGUh9SNypliO4VODfx7PTE8eP47gKcJZG
9GCL4A1GAVL/UItRYZN9vvW6TXIinKN0VG6CymVypCdroFU17PdCCwhHNFT5DmNQ
/5Kwh15tEKKgWAGVr1vcf3IJytiPkgA2bFJOiIIS4z1wuEol/kdOhsD7z9fKecPG
eNCij2D9zb4a292SDlpd3zeJaDix8lDXc/kdjECftNphu3ZfFuVJGjPTXd2c7ILk
j46Rh37offJ72spgN3DPmkI+rmv+TKWgmOYtDX8Y4kwwEoE8EDSBRwlh82x6cjBb
4ZNfBqIrny0yNzkreMpHvvOMiFJD00nMaGFm07pf4yzVtVygLpjAAv3MhpSlCdmw
YcqeARxOYQ/ERuQxBi703PXeU+dBeR/Do/ngBx/QSwE4gsgvBL40MPkEu54QhSeH
XaT1Qb6ySpelAt0TmtOrpu9hnIClhriracJjsC4t3zcdLMCVLXwjXlMl3pf3reXT
SauvYy4rHEPxsWvQBpR326H4RhD0/f4N2tMXIOuzK8Ra+w+aKLxI3oRy6Zff9hlh
QHJLUYjX0D8Nd919JMd/FIZ+Wu9wgj0ACYSTzS/2tBs9NB1xDrgiSPVQpYJDD70b
Tz8Swh8vCQSzUbfctOtRx7yz4W43D9XhHDsmnuJXgvwTP4i4UKD0JCafBBxbjLdG
W5q6MZ2pZbhmsbKfYJmazdUxdLDPopodtRQMm3MTomMyGFq5aigAVM5d0kMvhPII
UUVzn8qy+d2VykKmT3Utf12e3n+QIdcmK6v3IyukotD7QOb3yZmaXp72O9QFJHIl
b1UHLvQ9db7YMBZPWdeTdtwGY9EhgvtyEfhxTB3n4ktFDAYphdVEV2aavgxl/8xz
eGV518TLcNH9AU9ws8DpJA93+HLW6qM9Wbp/VRIE9h/SxXHZe12DKlLFRfu6QFnS
btojIEW0K/YCpZd3Sd8E3rhxI29MTlMmylfz8htS8tfsvVb2Kt4eM5FAFtZYpj9b
b1P0Qnhq3NFN1k10+IPyGCVC3VwnEGk+LpDDrDPIfWD0oMVwSrGkfqA9J9dGYDgw
pCGRWHiLTbwAJQjUhWO6gdMnfPDr3Xt6jbiG0JHgDeH6P7ka/dWB4UjDb2whuJiB
+X1zumdgnKxxd6Het3n6un+amqIniv9cgzEYdtn61wu5UXOFYExYbi45lleCIaVh
merMzN9spwdiI+iQjfv63NP5USHuXqEyvGHMELzQAoyatSSMLITT2TyTBoNfj58O
NUsdeVc66S/yhCyGEyB6GmqH4/oHSlBkXik9+LT4IKRh0MMDVgkqGomkwiGyVBrA
70JpcnkAGnfs9EwJBUjgtNr0+qiePpACbbGVAOnR9rGs1MutdQITpA7CKMH8B9mc
09nTjz77mdvcJQGBdq/sa9ZfECwOwGLC1Fh3lIcMxc0scNRKjXt3O11rjpedMs1J
wGjJMdnxUzqMM7zGZ1AR8Kp7gAhskoniLtnRxkzRqv15IA0Am9oX3KbUFzuPLKtg
lxGq/5hbuzdn4bzx+cF8Xp40vRqjxaZXNlgoX+LE/GQMhJ2xQ2M7MuDB+qL04Re+
prhy3r4Da6UJ14fM8kRaFaYu/DviApWU9pIi68RMA3lfKw5GOZ5vrD6T2uG2MLwT
rY7rAsrvl4GXoKr+gUJiFhKRDBqW645ZfHWh4G1W4qwS9+IYxSkFgm7lSdN0Smck
/aerHoihEr8bIp8UWD8ST8NY0fsaYtzIyQm5gp5RAOXCNzqp1I97X9IMM8iEocCt
Sk0IGr8+/XX8wc/4XxVMKSVJ+UsEp8Q9aVSfUMePCC9JRYdFJ6R+tp1vqSWB76sV
PPi4R1xs2GXVrSPuexS/AJ0brK6lD/lAEPDj0n7V1DpqUPdA3G6ZslO7UNyPluDS
3seo2OhsnN5Fo4ulfPYr0h9Xaf1+ipfBRQgP9AE4bYoyh2QDMPx4HcsJawxKcgqD
fU/qIk6J/GFeehOEJl6gnhubTJAvKITUzoDeR8pLzHGbS2dvWWYo1pcT46HAtZGR
NfVKKDUH6tBQV+pVSnzWYFohLOu/68SUfnG2urE6AS1plvnFhFm3n/UMoQ1SFnCl
jKvyRoULxraW+ibA1gPQ9ZeyrI+u3GYxSmdGhBPkG5tkTq5vF7vPQg1Mph5D5pWJ
B2Et1S2alOU+LtKgfCjOVhj/3KMD8p4An7eIryVGFGkTTb2L0pgkyv6AuAoy4TPY
dMW2TfpEuR3WtfDiG28nyFPtqasO3tUuQc13gDU3SQ6TailNNYbgg90FeeWFsjjn
i6+TN2h92ez4RdHgYMkQlKSskxdfqtkhEmaN/BXJKFe+pSdT1IfQv0QUJYzcZ7DL
1jnVm4myrQqrgOAt7lqFtRyBl5Q46yDVjO0f53xXpY1MCMPTKauhMJVkiGnSJxWa
VEkb5Fs9r4rW/CXW17rZUu53wdIOOV2maxyjxb7Yi5OUcg8llnX0fIK/sCz7xUwH
M9r4Xpt/cfwaJf707XlO30tmrh8T8DO4fz6TjwsR6lCgpmELS1of56qGyIB0siG2
qSvo86O95Xpdb0pAoq3tr2dVm5utSxrqJcRi97COZF9s4LvPxd8JQpW0WXiIU70v
5ZCZ/q5XLSAooUM8TjrdXeMVXsZGHHxqUkNGTW7QpiGK2XBkZkq0fE8IZbgQJmQs
SR0scSo02dAvBISOt+MoS8RbfNv+wgfGgxanwSqkgHVPC819fKmXBb8o2yOL7y8u
t8gq3cbJxmuE7MTlC1qAxa0kt+OjyPNwrKK77cw4KXXXYx2PHGJDHxy8EP7gNZvL
7MLIfusYLb8v9v9Ndvgd0d2jieD0MkRA4IZvcqhLE6quGDVAKbR1sabCJx0KXMiS
OTTINujxEL0pZUJyOJaJBAQIaz5xrWwzyqEIdwvkY9xQydgiYBJTW5CW0vaJrwYc
XL8DTt0QPQy5lZSAWPuIIaDtPKvg0y56oZjewBSqZRQdg//igaYgFreR++lHZ0H2
7Tmd40FPtfFpneTUUM2ACGMhg0fopDkv0R6RxHkvEfme8zWGHjs8zR33pk3/+LMS
mM5pIHuv7IM82VhQKALfY5l3tWgnY+U13yvlmakLlZViA4LXpSjIPEhiFyVqBoIp
EDiYa6HgvWpw4TyEUJ98tHLcwVyFf+XXv4QOpZ/GTg5njiCVEXznLj1GQYPVZeRi
9LOLJgX5/3NSnmjrgHZRpymfz9dMAqsETOXUFRUxz57lMIuJzYAuuCK3b0JTJI90
nEKhXAc98yl9+huuGUo7T1BBf3SiR32wQPDEwT54NfLazzdbEW+WwlOBEh9P09De
T/+bPiVWA0Z6m/RFYdZvqVQszowiVGAcwDiauvpDy9NFxklhDqwtRgMGrC3drOg/
NAIPTIUvP+2BG332yIrvl8lPrOEBWZT3mdkpV1hMImNdUQIelBaBr+F99HwInETg
TcI8fu9vM2v7su5ODIUYK32rzbYULpN5gnoZ7UiqmulMJahySvP3lXWVhdQJSw5n
cGXO3628QKukm6DK/xIvB6LQ/q2f+TjQe4oKrp2lLd5/I7GcmigB4sNK8nRtA2Nh
GH2S+Jo1stCqsFEhK1h1/Xs8jL01mSbYbkAttWUsNwzLh3nyKlhksJTutTQqQlZT
xLvmKlYpqvXCoiUZdJ6b+O8STrxwuZEyo/RUS3p96hHB7CUaXz9InbVDZn2ogubo
XwlYfcJkSEnfImTxsExs/ooEn6m6bT12W3x+yW5aeZ1lmvlQL9mt4ly2/GamwhVo
LZgnU5y4SSKcfCHKpmt/6GhcI2/p8YzFe33hDN47i4k8XPwbBjvsvXH5K/s5ms6q
zK/7DrIblzlUmu4LvkZdQEbNiEAaryvNFBUse8Ls8A+66NaFgFf3HGMdH+87OHfs
8U9HsoWlkekdALXiM7+JXTBlqguehgeBwZg0yNa0h2eBH2oNAcnP+nEfbXAPNTtw
Yhd6IBDtCkF+wpvd3FrB7Ej2/OrOVqEt2GSbPvINCMi3KWHURhGoRslrhQvAm6cU
wnPm2RAoX7OGHmalT7TIuo7IoTwo/AmcpYMv/zIuIIPZCqVbw2DCscw1dA8QzpCP
/Edcue1xGbZ4m8XrhlatifNMJlS10rewWC4cXXgmenaAl5N4ocudsBPhH+NFLTZ9
y4U0Wgt+Ml3tv6pBNLdDqzx6bjcFlJ4cmjZURYFMSc+c/JjviGboUujIGt6be38F
ND4/FpjvepAXe28g7FMTbLzuDIda1ZR3B1Ez/pac3zsEUrIz8Se82KbmtopGnlVe
UJCeK/wLxPgpgeE+0Cbc1pb8xBfv8vxcSmQsEMpSLVmyNznLSWUbmHLZKMAQW8Ef
PY93bGa0fauwWSBLaLXN56DtMNMJm6zRKBb/pqxNm71CS/FdkqTlp7qjAV24dDbC
QjRNDdikr34tB0Z9WDhZkOrWARTtjd0o8LaUW5srRkb376dlFfkMJGycjjOix3TN
Fe3OKiOo0uuYaj6tmhckQ/AZ1d/5Fm8Q2k3AYYoI/8hVJGbkMOe2q7PPge5NYefj
xwvjibDScqn2OGxTBYclFknH18rsM+04mDRV0ytds2nh4HNh0vOCKzWAF5VIhLo5
PRW+wENdsYCgyDSjib7tpxPU747r8H0yBqV/kyHcqqN3BCmURCkCnKEo1GkR6SM7
95az9A2x2I4wYHB9c2TxU+5ic1oaGZmGViOgt9jHa0yzwAjVIR9xg3syC/4cwH/B
MrhN8ZXrIOozy51jitM1NuAC55vStzQNqDEOdCT8sT3h+17JBCwDuE/pFJE8TA+z
W3O4NILmfT8hGRQMLsN40xWplYuTxc8RoHKAAD6QGbEAWxI1KENuudEPbZXXFeo/
2Z8gbA7wOuN1HWeY45xd6thimXZz1dkwrxbsTvL78l9ybeQl67iz+wSzxQR0DpBu
QvrDZCTICqOPauyvHi/xGPxp0K1skKe/2NERkBVrgTD9fGUry4Yp6riHj6u9wiJI
Gj0bs/zWwFBz9Fa9JoZzioPoWNnRamV5k0G11VIgb6M5rxrSD/+YGu0rKp3V7hia
2XVOWyZwtD/FXfVurrhpMtN+5XHStR+5CHXPJoXaKRLeKEAl1hLGv4I9apxI5Mqt
wmJbqmeGnmEIlCYBXb4Q3tz6kAt57p8HIg1ZLco9ic1Ud5Cn/XGA7Mgq4FwPpcFT
6L5k9RU5Us7TaBgrUxvGr6W8uVNQ4AuoPuLeDesAXc0XRh6UdHYcYxU1bYjCI491
B9Y7+gzsSKz42kbmXSS5dpiGxGD6Cu+ybRju/NlMIWSIv7RzMdcdirv70y5rZkk7
ACGCZNixnCkugTGuK49lDSHcjTbtfMZbUdAoooTiMEWTEQNYySvJhNJkwA2zFyYH
Zd5UwByIi859IQV5Ov1v5cXCJj+bGAx52CAuHZXEs6LHipy6AbZjHuMO6//aA+uT
1qPVwArv75X760gQ4WsUbbz2kOZddWTuykrxQTHhHR9VHZOBdjpiVPQJoEWqZ8A7
sCPtmdpUkNLr/8VKRy0TS5PXZ5iz344aMyICeO+gxpiewriQlc9ulH40ndb0m+ZC
Pk3P++417srZ14DnKCtvk7MRNN5G5DrtjO6UHdFK8XaoLsAJmZTJL286qKTyeKYA
iDi3PDBx2wC5/1NEfEZK72WZPgcEAn2w6frsLL8hxzeT7ujQMrKf16XQ/S2YzllN
PwV92QZc43SUI8mG0MoVRc1mvxXsfqe/H6X0Llxy+NDZJAL9C3gfluEevWxaMBo2
YcdSHHURcOLYihwwtXdHnHMnmsiDznqGOt7tPU9JBzX31A9LSkKKv6ig1gfqhXxD
nMP9lGhHgLA+btpbrp12dokkfFro5UDFnCtin03Q8PHJMJ+VwJmiAip5eCy24tDt
y/UsZhqSEG5xbgABZ+xkvF4Q+rCPul8QvXClf2dR5ficM4264f2E4g2jNgC8hgRn
V+HVxrTyuQnUeSp6oa/LDv5UtUsv6mWap0Sx2xOCKpCaJVfGqXJxn9GJO62Fv5gd
uSfe2uCCYWnDzRWKAsUTDQ6CV9+wmsEQTXqsTeSR0msXfig5ytlLiYqqjENxGp98
PbC46iF319gOCiAwiAlZ/NyZFw/YMg5PQyGHF9Q5Evi+I7HpPa7amcw0Wni2y9xC
B+JDMx1T8D5vMRyQWExzSNsYTW12PRhW0PYxJXKQEcE9hohkLbCpKehXiYfhQSQF
hc6J/9vaoIk84KhhBLmHLWzPslv3zYICiMYZ6JuKO0r3rX5YkSJ5qpdj6PaoCeJA
MEyKCp9P1WOxJ08IampSUIc3cLnsqhzBNMX1RMokGH2jhDCJvvzr2yVo+R9mBUEO
YbyIbaFIw7igO3kZ1hd7JGLnbhMfSBWyDNwOFhq5bJW/JOXGsDbsgS2JBAN112Gf
1o3f/SeKqll6cqA3IsEN6zsuJxvLpSjk6HZLUDh47kwvIAUONJLh7bVLOyoZkYMU
ZyL9YBELbvjzY1Q8hqXNgGC3Y/EimjjPBLmbn6OZrhOXX9WSNJDsmHIkSAKSzCXx
BFMhXzWggQbrw6hdQ7Okfjq3ixZb9ukVhmera7DXOgfwOY4is/trw9vOsUXh9aTp
60hvNR64a+J8Xth9uOF5hoSHuOWl+I6NBkfy8FxPYph3pHzbowokbsSKa/V0DBTo
9W04E+ld8o8rQic9we9DBSnDDiZOBY5ry5L+JZJrhO2r99DRqhyHsLybwtckRnNV
GnJPVKwnIN7zBugthK0/1RZHCtyHZZQ94nCGmVd1e5niDJdVgb7dEy1wn7nEIXa/
pc0qQQHqwFfMV9kh4EJRZySxErtFFCuCs+s7SJkwft1rKy23aH7q1uWRIjOigapF
5CvAW5bxmrva/w+n9GZ21ODMMaaWXA1UPHakR2pzDmggldSufiEYvjkVfARXSGAv
VQdeYZC8gk/NT5TVBnTI1ZrWY3RX7bdxVfrDhvgfoN7xvF3D0yhhlU8P2cpi6knq
6cqbFNWU+YCOg4/YQCTErjxg18tmTGIVpcraCCd6NVLdZ72e8TbpfNWhUDMYZzdj
+LgqwLBm/JaLTMOEoqBkL4AAcjXjtT+i9/AQP56o1/YpaB+6woUrwrmTelLGOmPc
Aly9IXHOOi+U9Myc25g7e90OxdygdOVBxAt3OqnHsWu8/WhRCnliblXZ7M8DwX2P
bqMYgyoL5LyfFs/diFPQ8PCob9UlCNvzu94dY35rghg85TYwxsxpqT06+TyEb4Vw
VRj6G2Bk+OL3RyLRBNPeIlzc9w3Cc6DepRRY7AIbg0AsXGNXjpSc9N0CstLIkuEN
0yZinVx2axBBhjEfJk5+6l0p9qry80KH18fFK24/T1H9gHnq99Sgz2yBiI1GI1oc
OXlCwPSY6KBfTpm7JfMkPCXlSX03WtVwEEGjiTUqRup3be/TPGSzyrBI+QqG7vxc
At/cE9BVOmWQ3vOSYQtD7+f/2BDYDcUwQWIoxmFuOBCe7hb0DhzUuYayvNgxZr8J
GC3zMando6zt4t0UBiSlLiX9AoapN5PcF8/+WifkUdCTCmZTa5jyHHQWfxbAtC3K
1xeB6pxzL8y7kVOY2THLX1IVDJGhMB7cTmITQympIkomCvTO6LZsG24Vqwgje2T5
JCpsRROQJx0v9NqeAxgdh7KrH+dAOZfW6rUijbvOUlFrz8OLCV4b1ARyNjtJ12JN
PzpMtdi1JTj8wgmlvv95dVlr1NtvGVFvStgGg6qtucUdGIfkZFWEO0lXeQaIKJrG
jlyKjxxY8nKYLtrlJIMIHPKZ9TmczK/7zUb5AP4Fn2f40lUDVfgxXbGgpB9u5v5I
NA977s6/3zM/59G+7/S8AAianNnQFiDXFsGlZfXHd0d5QplkZof02lkkkrbeQSwO
Fpy1Gw0GzCgq87smqHABRXZHs2ql55D9lDXDDeK0xu/+nmsyvoGHOkKSN7HwR320
7Qc8CUot/UtiVNlj1R+ElBW6efdifDryI2NuKtHqWkpTHFSiSqXvEVhyIwHNllOB
AdBBFrKI6Zt82CsOLx41eLn7CWLowb8YqYMeSFmhkgH/0ZvRyM7clxsExFArMFIV
zUBYrB6Rew9eUjrrcMVjryF3ePrwsbafepI0MxCTvbhUdZWz4vOSw9hP+HaVXOOJ
6eWMdYUvNwuzzdZH2yAUwg1PfMBnmiHBclzZbysZ86RdRUjA+ZmzvgW6ACfTxh/F
nryGWXKdwfUGt/RxxhaxkGMdfHF+AdPnhxsMUE4YjrY1rozlBlPCm/ByJb75tOJ9
SkXbbtzJQBx2xpuE/TohR6hbiIglW34zwLM2yhfR6Mi/6w5linvb2bQGRTZi6HEW
vQVuUnzFl4JvUzVkLw/CcHCFEbxTxSSMewPPCRoKpoMemiEAUhMaQJ/Y47pN+0ir
g8AkCN9lRW7g3Ka0XVgSXOaV2opOUzR4MqygjPIC63Cb+ZcxsXvYbca1MRZWJZd9
BrELCjcT6eXQM0F7AcKVaDThCyyii7ElbK9GeR5Jv1qcqOryYheT3eJi1KhehJqO
4AtBOc0NG9IV3cl0cl9LPxNWgbiMeTpEvSNQ+vcZkGm7csL6cMQJcM8oK3F3dSV8
JTNDNUPQABzW4CgvKitxk1K2jNyMz9BZwjRrr+UEG0H4YCTRc1SsZvoN9h1gFpSQ
POQv+ta4CrBeLKGno722lhoXXP/hhJN552gPd6+FH+cPmZVO/qPRQqhS68SYgHTC
6mmgFWRH75q2J1eYnlsLt3UWTEgjzVh9NfgJ2czefMWXGGj9KocVH3PFNUG/wKbp
UdBT5DPNrRDRvhNHj+r4GNMbkTZPF3GPTms3rwhW3XqlY1Ii+QWv4iKZeVFNpMUy
hkZYcmv1pagFUc8Qpsau/YxjFAl2GK3EzE1zRimV/+rLUF96b6s+XRkWH61ZqgDU
C4EB+J4YQT7shjT195q1s61UecIpglwOctAzVvlUoSQa5F4TeO2o1UGJvySQ0Ltr
qFFVEtpOrqTL5RHVBKNVFq/8bo0qOVfNPVNC9SLM/R/UN/3RUaTj6vne0Vy0J30X
De+yBcORL4NV1AAKZYldsYd9wwTfbTWXUmm4CacmMwWnfjzl62MDTXhwMWMwoh9b
vTuQkEpXmYYiFGOe00Vr02cqPj93IlFMVaqEIHCnwlotnDscVUCocvP23BpSQa/Z
1yGqNnDy8ZmPZ8WLoZ4gThghpbIm8+6bM3GqejDSaZrl83uKUQtfYRjt6NoRx789
Cahf1QCRXLlVd45OxPCsw1I0WUnHJ4jDCpSfq1WJZQ3hFEJYuxy6O3t/5HTo6L6s
jwu0FQlr2C/2FpF6kFJH062u28rZ2q/LHmImhncaGQeBJzIpyqo7CQz1o3daRGA0
OlYkaqy0AjIeiF420BC6eR3Xv/gTWPfa+9SxehqzecJr/jXIklo38Ppw5RjPAY2B
gwcsHECHfdViS4Kmo2i0njskFmH3jHf1aLLhBvxlUAsfJmgo+ZNOhoyV+5FLhuAD
S7Pv362u89WdTxXA2kSPW2wfnaicdezXbaaG0jbTQhHpd0aQu1SiHyCwJkqbV/Ns
/g3R5bPrajdVLhXyfslOUCJKLci860Me3YBg1sUXDBCCfcUcCm0JZBtHijnuP0Es
CHJPm5N0U68v2hFcMJ28Bxrp+mEWAUjtbNwrYFCOsXgFvCXj56SYK0vW9OaNp+hF
GtNieYHQoxt06xLcZA1j/l4s31MXOF7/KLc6LmZ8sMvQ0S8AHCBtSddtZEgdoncD
Tcd/R2rWWeTulKcZt5zU3wEPGKtnzxMyyBLIAS6oXHFa6I43Wrb5j5eS+GmFZq2V
VVpov48c5Il9NWwLvH2H0TqHKETLSE6RHc+4LUIrrv+8zYCyoOvd/I5L9pNMRnId
Zl1MN1Yf6p3WgBvDxXB4z7sjAeYUYsk2FqhkJRB5ISNsbGurdf4BoMLqiTTDaRzG
1Zr9QZgjlixmjpCq7oo0Xa5uj6A3XQDmgYP26xtaOEIj6hXY50Rnas0jEfDfrHVT
DfMYZi0+Dx0T+zcBp+iEO7co/cJ8T3WC9+xaSM1UOjPQfzsmn5BqIP2tzuPFt/fy
pk5ma/aRYgUU973OGuHb+bZ33+0tbpW6LBNOxN/Y2mFmvi8x/JRgMGmvUPejjg7B
+Eb3BaVRvtZmNhhFTriV9lQtomDtZR6D7L/eEsBEXhoaf7De2RXdBqHEOHRGYFRe
AasZHVtEWBx5mL8Dioyu4v5mz7TXxOBoyk4EMYVZDnfM+c0F2jqZWT4Cy1iAlhcj
XzRPEM2MZ5e+KrLPGoifl2dWhmET8JtB5aWQw1KcbqnTqCuYJV8hNIVQy3n6fUus
xoP51Suj2u2dFvjxwFwU6KYXRvm6veX2u4wcA+5GdMZlSLEp7USfVo4tk9E/PzKB
wXgswnJljICwYCMoK2ZVMURJlSPZs1SXE63lJG6WG5sB/K115bQrgbe9Ox0TGnfj
0Z4LZvRbB0fjacbMy8MJX+Z0tekR8UUf74VL0yViMkKF7ZKv+f9MV4zQHd9g6GaF
YgmU9lOk2mFpQ+LSH7ILf/zVEX533/yOaQOK0W0BhBs2nWTeSp/6eoR6aWRU6P9n
YFldecmG4IDOLfHDn3FB0H679wg4XIvn9Q9pVzJHStBO3SV1RThg0i5egyp1ONYV
jfrYc13e5KpfKZrdTsATBs/U/EzZbcFmV+L/Xmn4eGWpRRSJGUsWg9RFLy0pHJb5
tFOMMeSN5kmffws70+wSA8zoAQ3FOJi5bSgjA9+vlUDyaJ5yJyuNhosARKogNZJP
gytY1mt/LZxAOCYW36mnPTSIWZIXa8ruvqvQWDSATr5EVVzCIFsoboooyvciYsw/
nQ/b3vvaTUUdXZD7nzt0i9O131O2ruixFUc0Iw2A3niO9jaa1ApfTehz6Mm+oemF
s2ifoTRYFqhmUndAXYINTuJpC6DIs/EYKJEGdHLu83ngh7wFXT8q3croAZl+OZj6
/94WjIJ0DW+0NzsNsPF/qyEfCz9b5lo4xMt1WG7eGQLjErUbw5YjtwF5JbPBhpnc
2Z5vhCSdBkE3BGtFS3IiUH4j/HV1O6wwoYidxfBDmXjPY70yP0QKUPmsWKjjkNAP
wXm04RsQNqn/fVxOj/ZhJQJAxShQBOaq8wMFtIwa2ja+byfGRaTngwUrqvG8tgWo
JWmYA18hOuboACVf0Fvi4iaNK/Afv8bFDvsGCpH98qFLIgynudR3N/zgJij464kz
WEtYvtcFVHAEwYKUuN54knZ9An3c+SsKtOQV4oHQqU7SimWZOclrjmujxUTfm83o
K5FZXUf9kk13D//Nm33AWRtDPqSsovqMn9OWuli6MjxLtYTUPfj6ADSfppw4j8hS
p7nGpICw2BF9lenUdS70Z/prYfxXrAQ29LTVQ5hzMNOxo+z2DVOg30p5WQuNDEFr
Q5iPBl4vHyqEW5i72GAsL3FI+b0AjPfB4DErNcAW2e2yL/CgrAs2K7beG9Eryg/5
9JHWQyn2IlfneMdmt1OkwN0V7YsAzoxg1GjohnPocPPZ3lekYRzhvqeJkMgKGa0n
as7mjUpQolGx09sGsz/MfuRZszXHa3YZLbCNLddoDtAVQ7L4ScwbhvHWLn7UpmjX
YiV17d8tTRA69TZY9Gd+2x0xRsqbkrEmpgk5aGSIFyFFHsWLYGA2bnExKwsVphCR
wkn4u+ZNssw73s0QhT1X6QyE15PIIZbgQK2ZGkfq8+gx1yCpWqZ+HDc6iGsg77/O
ba9QwgQjRWh+/AaDzH0vlSCzPmgo95aHJxi5Zh3kaH7qLRNjx/YZvgje0M9khXFG
5mtExK9fZ7YM5RoUEabtOxUsGtMWk+qoGMAd+wWBVaLnAq7iu0Ht5J1KU3/ZFOm0
5bTO4EbOWV8FjbAkSUa8l0O19ixPp6gZbO/Ze0kiQIaNN5gu0wY/poc3ki6JYJHr
9X2eM7FR29S8cQTo/tQbPmoJ0r0nhrgaP1IvhOnyHzwbroHEZFfQdG6WykPAiYsj
hTUAn9f/S4lgjLzf17bmWG2Y39WuIoKn8MAc9cP0LL17/MOWAzKVroFXBpGm2ZUk
aMabOfm3zRIqfHuRwaNcuj4oR6/g5mehf+zUOtspLXxDqRCBVUg1CPHNQpnEf6ej
87yo8gfsnUBjYsaF79dTqkVOIKKoQl2dN/Zd9ZSN+Uuw2HF8c+fgI10ZVotNjnzF
k9klwPw1tVVkUdPBIgUW6zivWIVKtw4xcqMwIX5y/g5ktVLk1Y9ZKhpXayB7yBdZ
7PGNsGFXCOHDE+N2PeI5mp9hXBH1m5cCd91Vqv2Ud3rQYOUOyCV9s11Ndx9mhdRR
P/Eh0o9fN9AkWfmU9iNGBkOzkI5Ax06oWUpN+ZoykpzPSXVHRuGN+PoFtxs/aEE3
D0MlR47ZLZ1h+QoRHzmVrVeoUu9nQf/YpsJaYj01m0G+yON4m3XbWhCNMj0giRW+
QEviOnBE+gKEhPEq3P1rJq+2CKFzMlqwYP4QcBMtLHpH4vuCMyQ7LVQFFFtMBfPr
d86LoY+C9KFqUTBA91YovxLlaAGTtMdPfIeXrwV8YXWuFqkCUQ2TBJZ7QRk9Znbp
d7u7lE1BNeoBiUTcEJebkQWfpYEEGpFZed/Ee/EiylcTUCcmbCRYhL5KeAqc5KJL
RHZcHqCdshRxNFeiIHcHgE3VvuX2j2eFWE+/60Q0pyfq+rafyT1J0ZkpCwp6dOB5
7WQr91HkAYJU1nvTFaMHNnmh0K6FCKT0jO2ZZceku8bgpkhP3nKHZe2fVMNfyNEw
8xthME4ueKB4CB1r71M3Vi9xfZea4BPgG+4DYjKAEUhwpGljieaObbPJwpfebz1g
POj7/uqxvIccRmVAf0bGOdTLdGfNBz6GckrXrBxkPZyNidTKQ2tmebPZNq2smxLu
La1c4tLwEeTpm5W6prN2DrGe0P9QKqMRW1ga4bUBUXU6KKLYZSBdnFS7XcmO+/om
q/m4K3S0BxBtGuGRRB/h/WtE2JJYtW3R9bxxTl3E7lBMQNkyPELD2dqcmV6KlZkt
xidl9+uR+Qti5f3+8bEZSHIyQ9K3zsb3OM+nqCfimYVh+/hjq0Z1clEMMTfprge8
8TxNagxqYVhym3LHkE0G366Dq36jckYyWGw7LGMxQn5oIIMQrvwLvDwwpiKy857c
mValEF3UgY087Mnk2kekRtiw7uoeYT52GAeQcpDUBffRENeILKcZWXcUcKjG2cO2
/ORAJiAWnIBaO+buL6HzEnmEfG8ZFggs5FMZCeEfqyT12zwc9XBW8rweXxm2hN/h
gmAfxxuOkYHOqnz1YcjUu0blktJejz1bHPCtzXEjG0HcRjyj589QhfMknP0YhA6a
4SEmRyWUH+Wg1tN0V5+GkPCKnLfoRbsEqt5+1V/wPilyls5wYx63aYLySSZsL0IQ
Ak8BSPP6feVZ0SQ2IGRhwMFP/v1MpdmpztsDhYBkt6KDAhP6hRi6q7xem4iAKttB
HWP9nBt7AO1JvDKz45/zpPw9svBK/8dcQPA7QOrXnG4YxHhXXk79wKO+irXUX4ij
VBRwdAUJcKsFEjM098vGG3lBMKapP/3/8CFhQerUr+YnRLdYhIgwWViuhLm2lLF+
8ow0w9vMLOF1soOI2qQI4yfpNvituxs3NottS9x1V/C3Ug2NBi4C0xl03uroWXqZ
rWaXqbJJyw0+fc2Np8njMZ3D7xhv2Cyb7izUn+NFfXkADA3JTeLx78Uv3b3Oa1aN
z2XvQzklNuhTbH1Phdsta5qke0+6rgfKxURAsN/5uA5+p34ugotZZBVPIKolCSsF
b1ohrEL7XRywX4RrScE6uGC2yRJ4L0MtbofaYkjJ6HaHBhHtmtXb5qVesAkiEMIH
PazzVEBBTzglOMiubnjUbABAadbXi1Me7akOy0u77HKMciqobddZ8sRWFw1wAR4G
5jw9V9hqAzbQzHcjOZhOx2/e/YuZ5yNMRtJLmkqZUBVb88L+hhYHx/a4hT8Qyfne
kqBuxwBjeYGHHSPf0WLbqHNbNehg4SCqTh3iz2EnWwDuJYmUo9RpZzLqXwEY4QCy
INzQ40dwICMrh3sSOCFCP/RO++Din6rVMqguCmKXFTtTk2tNtUYVtX2ZKbPefOja
dpokd6h29mxh/WZf12kSMYF8DsEzk61iO4tvZjMg88sA/Qbc+iyPgvddV1B40GG8
GbMzG2WIms0JACJQxNoNHYxgWE/tnxGEDeMTEKokPuibaeOwiHFNI+fk8x3SSwVX
Ma8f9V2XZDIVJkgcjaq/9FU7tcNJR2UuKHV7UyBnJpfI0NmHd+gBbVDT/OQSlNb2
o6R5Z6JxCC5CHibgLtgP81t0B2UIfptTOzVT22A2Vdh4h9n7eOo/uFUjFEnN7Fba
bjWr9frLgPj9+OY6oQVrx3SdbnZvARsvXsznutkZxaZCZVcGI68w6JEDGitAsn3N
cqlZBwy51lomgPrfjdsHmjryRtMl3Xb4ptyiacF3GQahHxvuok4/HA/bqvKEtg98
7WmyCQGFEdrXlA5Lve0K+qegqpoZw8L9Rw9pqi4afiGSdLTbKomc+6Ndz3hDBvFA
o8SyZrBZDpskNjg5X6C/pw0CRYmudUHaPo5GcL82bAT4nOX1y8M5/8cWgtrOGkug
ifzRgxUhlyvRQ4atLMU7KAgHz85bU16HNNv5El/PcGAOc49IaUhHUWbo/w5UipwV
IF5Xq7eKxUQBkZgKfFCrFajpHQoFP1ddpmKooiIEmFB91F+FvfQ4eIzL9kq83tHF
gu228OSpcGE/FLqqYvN/PT0rggajtzPgLAxU9u+DTt7RzqU0ZJrJ5Ttx5mXz2cY8
TmT6mKtE5jCz4tuDKnLn1u1fHzEejxRi5ohEPsR8YAYsQVZ0SV0MQhRWJywAdMrT
K+/eJiwabDuSi7er4PEN64pIeCk/YjvyOGdnYJUMuIp4GOwbGHFpJFJEPBCEndLy
76adlCM+jqR5IW9ngltQei4D3RCTsA5YH4oq2yVah+MfgiamzhfNl3g2ZphHO5kp
BVN2zvP7w0xcO+q9pDJNS26eVOd/dSiePhKsgJA/X3xZCNdOXHyrv9OcaSkUMytY
JgYCYS6Fo9PeeZeJdDDWLOkH0mo8JXR8kvgxAMxFOQbmjsCW8B8xpbCdfpq+qNyw
aVqO/+eS4nREaScSgCp3qqWXdJYY3uyPkuZ8mdbFdBStXV9eQMxd2maxMHAAMk9D
lI/nr0hY3LGNs46ie7W9scEJifpYE/p3A3qnJ7861gGc4w3ZUfhDiwUSzaUf1DAI
troinOKMZlm4D65ATQ41XcrbujGb/IDIGc/dUNEwKDfFMfJToMH+iY9MiyxV9Hnl
qyHgI+fJn3A4EfQGXXznpq2ZmMteTtHDk+BVyXWbuBMUfN8IKtgzcvjjaHjsMqAn
G/wsejrswH5nCDSAtGzAGM+ZrvstP6rX3sZnGb6ug2HuQpmX/O0SUtTYd3/bql2U
kcjW4ndkpOwt2MxrpkKEpDQNUyBO96gKXeLL88X6RGPe96gpQNmV/indm2EtV+Bl
yocDiTSOCuAygtZ7TEgq/IY/+ggjut248ytQ3J+wFMk88tSldK8ifvGe6jLpGIOu
m3OWjyn6VPN1CHXbjYf9qDIg1SAjBlJNhS/Mk2sk1H7F7U//YtmsWJGRUafGobHn
TTnaaB/T5xUPzNYMNIgRpSMkPz8scm+aJiqf/DlnPY6EolweFRtLGF6B3Fb7K9Aj
1fRvI2Acxmkqv4mKlmRIxDpqxAG3GYuLsQ4PfpHLrqK9pZfEpdQy4D0zdhCmzjFr
tEfHo+luDilu3MuALPK7KyNhHp0A/g5AZ+eiUemIOPKLosmYThTZ6eQy1pVkobK3
DjspnZDzYbidwPkaxDKBWx2CuGjBlGhnPLgA7fHOG+ORz841c71Qqk6RYo9NhdB5
RPF0OOoI1E5lYyiL/jUn9VqGVG49aeyR4/RkyKPk8Fy1UHIhgXgJF35u3/gACoGF
UKLC9ibfaQqH5C1uPbLhxSBV6TSDG6m2X1alepBEYdcWaGyOlgf93z5oMwLdCLso
tmAf4JrOtz8TiyKXXkXMQ0yqMpupuzCG9P3GTl7M4lKt/GcgDtKVvtRMYq15Iaxj
aMpzhn96ui8S4cbsy2vjDavYR+z1DS1UXIwtBSfwEEO7Wwka8mCybrAYq1xQ2RJP
bK+tOKsWCdb6IsHjpC6yEhf5KeJ4CEiQDPSxZzJ2C2G2mKBCki/sTf/eYNMfrQoG
GGEqgOFLEYlzwDlnMyCwE93nBltq6dJRnHYndPXS5JETvoK83uRxRBm0NgzKGWT5
bmJZvNDi71U0llF0NdhZI3Cb8c6bwuNqO/05H6UnTQahaki7Z6xY8pGV4jgvHF4G
JNzaNv7StK59jqcnAs8rvdKqyX+CiaYOWnizyOjED5gfxVzjMrWo/lQ5ujH+h2yV
a0G5kteeK1XPVE/8Q+aGRvXRzdjSgcRN6UO+9Nde10XMwHqi72jCM0dRewL7vQby
F57Ys8SfXuerSQwBk619rP8w4C6O7A3svPO5r8ZhehupSVr5s+bchR/odWDalXHq
Rj7YtgcBFOXuwGdKLs1tffb/piWkDJ/68tk/krEnq5edFcfOfv/KIr3d0znaON9h
uwtPnq/kgGC+x9U6Uq1r21YfC1leA2fEAmTRVZplZ0BEnVmBJy8ejATHb4i29aNN
7s9JUxYq0muC8kkTarhKWrqPemJ/+GT8KpXbKmNOI54TzV6OWgWQLIdG5L0XuHDC
asJzFANBtMTKBUgwaVC334tkmb9RTYsWfyjDAqTWUtsR4fk+J1WOA1vi9gYXlym/
jeIWbsVNR/06cBkVCj4uLvNPF994rQ2LrzzoVBFPB5VT6Vv+CwGD0CFKuOisOlu2
JwcxElEkSKk6A0Pd66/PBa27wOKkW0f1+vfCFczzn9n31PaS5kDyABVY30nOXBdw
6+7Me0SMVaZeSn7HysdsCKUJNGwP7yxrb97sd/qjE83z8Ivbdo9EjelQFtZAW9JB
bjTtDAxmSFPiLbOP5G0VYLWfXl2RPMpkzBK1s7efRMA0SAXOxaoLC3v3mWLwIvyB
VZrgjYuGJd0KIdlZlMhmoIR6iBIx4aklcAnRdgfQPTAvlITNqR2OJ6hSk+dvXW4l
zHc4WvroDf28CQJUipuQXlTmkgWOTSJ0RZnqVVOApfBWu0ejLQepV2tbYXpjSajj
SKakJb07Bg8OppCMXc3Vgjk6ED5I3U+xm19FZ5y1RExmNOkqniEeFMlANuJcYjxt
CU/3wBjcHW0jmI9ROMnb5fUDFWZCHBTY2s4ndbcbbDQj3Rmct1YplmUEAH/41gaj
0djwzjlsXORYv3NkynGgdOKWuNO5K7gDfUp2raOCzWGAcFFpc1Hxj+a2V6RDQnVa
DyZL415Fgmb+ys0/kFf03UfMfEAvWqkH4jhiMi+6oq81BEN9itndaqqTaU1lAejY
qCxV60FL+GbxToapXjUwTYmYkRgCbDIE4FeNGLDrDq7b83gy1NOtwmXup/LOdZ8n
6hblR7zLsvsHLrPC92ZTp5nltAR1shWGMegExo2mgiMDTz2ywuIJMKcIAO1/ksLE
dIHVGTeJ/k06qigbCU4ZB1uek3em7W/fdGL9BFGUJxKGb6DRGJ3AWLYqjSdxegap
dmRyU+tkSdY6TmuXrMO7NV1V6oTUPKoBh74yXNMzD0zG2l+yFVa+ykBDHgZZuL2P
rtfjLLyvkJG9H8YiiIeCrPTU+EA8bS2iFmzNB4DxG6kDjyVhAtk8yO0Bsx1FNmmJ
wD/AznGNj1g0joC1szPlRFdpEdHvvySIDmtbJ4OS9b9rzyKk5Fn15QgQcDODyvwR
6CFTN1dfnDonfTyIqBHL7EXfBny90XC32gOtyShdBoBptjLXfuizD71t74FiYiqB
C2LVXZdVZ0ahMnXX83w5XhdZ8mtWVspoPYlyEgBgKxXyr1ou20IbLYlLKzvVnh5p
xX4UKvq3YIre41J9PNMhfOKpZo+BKPgNduPrycjBsBtb7PG381ZNMG05FyYXqd3x
SpkT6bW6oqWkYzfpgThcUtuVAYu+FA0KkwXVZPYvc0LfOZl3PA3+nRUIL2pGdJnv
41aWBjYXIbw8FfdT8ju1gcEOcYXOtjlOz+u/iGJkOrH3S/qYZgi6BU4I/BQ8YJ9R
ynHyB7OFYgLOpsiY/ztUnIU1rK6OtZZTCyhUDX7VOkSt7v6nsdzPqEBjIO6uCeov
rZ80gvNP/wucJr6tmK5menUrHUfBNrHYM4/Z5TYmUo4Ncw9Wduu5nGM0mdkluZY9
c5AQWXUNUFx6ANB481SgGAoAKfxcCBzu3bUXLTihQxoQLIK42/RTxGO9FkA/1Xwz
fbxSuDEBN5IqHbcd4nlm9Qiipvls2F7IgyvzSmpPauIpyk26wx0iIJo5OqeAg7rg
7tqJHyxo5u+DjduDGKzAs68gfw2Z7L3dj5YlgpwtM1u220b5lVg8hStfq+IGGAES
g7vlA9Ehgs6lncV50/C+T+tG1XKfUpLxakrPSWCshcrt8/dceKeefUdWM85OMZmm
NEGavfh8xWyXt0xIrqAXl95Gi3lnP1qh38G1FeLbAGZKTRO3M/uDHgVPE3xkekfx
p3aRBnFirQGT4IUv31jQ3T/uu6DowREy2SKKhveQTIj4uyy2R0KtJOkacgZUFtiZ
2GYCKRtjUDwy+B707bMUdE6EecUlFFZEkSMlrUlZPYGTimVOLHKWJkyBH/ZVLEYZ
kpvV0UeQ8Rgr8CjZsprUAf62tEJSJIi2vEjLlrnByN6nzBVN73G5aT44OknGMtqb
G3dLqULe5c/daNRXRck5YigdcqUr5xaP9vphdAAy+qKCEkI/MyqIltgr0wYbcB4q
tuktu2m06wUa8nt6gKINU57PubXdENm9Hg8OIaKnM9v7vBBl+gXQOt3AtwV3c8ei
jxGw6qfBrNGM3H7mv6S6Y9CygfW5SIdULA1FHvrFUan5PaRMX5D3vNkizlOIy4QQ
GFWlH6avEJEAIZ1Aa4kgkKzMHFUEARuTTGm7YjDQx3HFGUZcG1fz5OP4PZpdRTKL
o+I16tLviTHeZwuxqTJlciYq0CShvk88NUHYEUUCT78YHNefyPGNjXfh76CfKczm
PlP2Y7JNZr++vqm+Ww2b0TM9x1mcZs3Tqu+L0hrmSpFzCu8XE80efHvFDpU89sNv
0a0mGMOvC8Vlm1vGzKicGIaL/ZYNGJjjVC1F5CIz2LYsNnw7gSCZjzLfOPpwzHUz
fsz4MI9BgV0aMeo5IbQtc8UmsEReKHj05T+idtQWehkj1NAiVdAb1mGdHgExNUK5
P8VA3ytjEz2lAKSXeg8S3rTsWujjotRa/1NvuQhbeCM9ANXw8OgTAS5vozZtewD6
ZTyqiVjbOgKcJfFNh+0QDkgFcTm4Cagy7aIKF1hTsHjfvKIIRc6qszvd6s1NtQVq
OFsfb+88C9t9tpjN/J+/e8kbyNYnwymaNwPqNEyCNWbqv85wwbpdzZA/iCQKbCxu
GQHRGRBUZyUuxypE9nsnNlDl2ncAYLYN+8ldA9hV0Bzdb/NPBZpLrUzznbeTmlv7
tU5v+PdJXhu3+eRyEaanHdE6NgMq/GUPtxU9YA4IcdQjzqpojD41agACpwOLtBPL
rv/5CQaJ6w6XFwpqd60PUKOd4mEgyCwplfHQ+aqC4bo6snO+hSMBrI8LrumVHetW
CWsLUyQDgFn+U64IzF6VxKgdCJFZ6Ir1k2QpbqB5wUvfmXcoXQ/gna5a03ly6TKj
5Wl6QGTFaTfcsqP9ZfQrh3Zj0YjZnrgD4YUMWgXK4fiQJf+SZlVhLpG113EQX1kh
67JAgTvBHAl6U+/mVujm6QZ44vAf7xI4iMyUcU6SCowpM4ARfgKhR25fWOurg859
dDVzCSlB0BF0ieh1Kv06pyCOh1rbKDkHqsekn5llFcehKOCKR4EWjIuOWGiBzoy6
MRZji75QVfCiqulEcPUKH4QGHWCN4C7jIUK8d9rTL9bEaqYrPl0rZb6xgFEEZLIM
zSs3EhOE/LD7k077zoiL8kkhMEXd+MF9VGjrrVUd8ovNvIuNnQIep85qkk5I2a6U
SuV9O3x+QCCPThaEFQ2zrp+QbAFxvHc1aN9isBOQbvOMW/QzVKCveY8vJOT4rkeY
2lGLXXmaoMm7RIWEj8IHsXCfl8SdxkyTbcAhV2eSMDAMLuf0kWnb74Cluja1f3K1
CUpebEk6lZ0pTkJ/I+TnxbMcfLS3Y4BteeB/q+tgKmYKRz9n2riEbQcG8PeRWuaj
M73lpwAV9Ey7dSFhr/tnU7g+ye8iJk96n7afuklaMU6Hlk9yKTuyAXiL/Sq5FV6E
mWjFb0Y5vbAyNoUoleZy2hS0jCLQ85DrcdSqhl+u9+S43W/M3mGdf0jFR7++Ml2C
j0v2F1ue2QG7O0oi5lYm+Ara/COm9yKt6IRLrcD8ekykNEPiQ+R8kT7gswpKlJg7
u60hDxMemi9Pd/vZ0c376jN1ZUTIz7rMPvWQzXSoYsMFmTRCh5xmby+OaDuU75b7
rfsAqgmNcjh7vp2BwYGMDuA+0BQe4abf6uaqNkuhXH7wFFYli/uXmMiaZUGjCL+8
PBrb1dgYWvJh4U9L2/InUK6JxWQOaKCxx8MKjqI8yaSDXFrgcAUjB0W5S0I7zDtp
zk+8IZJ85saV9MXyJcbNEMrx7eV2bQF/eQbWIRzGVfkmHpAywkXVgtGCN/vtt7R3
T1F8zDARXkBhsx17e/9JYcCxDwVPLyvjrMlK8js19LzVaYIZ3+GrtxFJbEGe8IRW
qhmQiFwSQdOZE8eu6SE4ZmAn93EjoXBgu8ptBa+hAITG+c5vSjbKop6AS2EHtCBd
w3o+1zlU138ZuLc6K1O4VhwSbZ3VrhrB+thn9SNswqrGNwjagAoPs812tHn1OipF
apRNVpegrdZ/llqfnwPu7sJ5dVZHmiNi2Lmj654lttQEI8Rbcqc0yoUoCKZP8kLt
zIu77d0vvd85dd7t1bzkLtWjBktJfXR7KGQiEU+1EX1GTCVBNiLlpBqEzN//jT/v
gL2YJoLoidcthjLrcz9cG3+sYu+LZ0g4r+880U0ho1jOUUdgV7Qz0WroQ9B2ScD3
BF7n3cPIYpj6piY4/js+mjPpwtcf7VFbZn0c0BgTSgNpaiCp0AkX92RN2hfvBQTn
K1AgQ962nFbqoJ+cajFRS4hO8bWwf6rTbhNo57VWAg99o8SYHgSsqB3O/3FLA+qb
mRm6XeJHpk1OEQDnJLNvwxRx8P6Nv0KKsQzuuxUIJ/TKMOTOkEF4zKHVC7qxddBt
LcTh7NrzNhcS8mZubHYy9CB89SPn7BZrv4uf0z6qEofuVRteMLQNVis7OVRORLSm
skv4gKW3WCIviBxxF3KJ1TZhOu7iEhd7yY5rQ1eJS0dvLqY0PThqwGtnF9k5hFP4
cQvKveaPLIBTTcXZXkZ5Kk4xCamJw5TRRJYb3gFKplr8kNLDHVYP5ht3FmQ8YOrM
nUKyA4LLGEatMqjZYSLeBWV892lpif6w7ICOYo8xOBeZYXShtahtEX3jOO3er4Ql
orjW6BHYpSzvvUUXZHPoqEAKZLXYDWO1wQnmlvR7E/CNrqGvwYWQwJ/vsxaAiLjV
SuRzT7kVM51agzOiXv0oWL6gw48f/itsEQVDTPXRYgL4MemIKkuEFyOq3A1H/zY2
XVTDgX4b3uOStbX1FLBmYGamSBGCnrh0yutB45YBnWoRNixZCGxe1sRjFpApOLLk
6LTnkNaIvGIBRQGzT+yyWuilNbEPANBqIHJJ4+g1s0cOybIfc/tYHayQqbTVUGqo
MbN3qZwkIPWDt5z3yH7KZWUkWY5KZxmcCr790hNaI2eBnN3Wr9DdCUXJSw5TX/hm
fELmytya/whLlM6lu9mJswr0EU2si3pcVfqOZgwHfYCoL1Kj/q+sdcJvrgADm3ZI
zQ7nnCNnfToyKe8PITber1FwNN/lBxlLVslu+ni7TH/UsAl4m13Z1OebGLc64xHw
QZVjE1hlu0GSki6mPzXAoJFB7uhN0JQLZ3IhCY403XotDwQNF33YmONfIVocld05
2Hfs/NKBHNs1Fb2K6lBpVG+OE+U4+6cvODodbAIJdKTrsbKcRE7PKVSXpIU7j3m5
XZHQePUaYqDVMgms1K1dfaEP+7QzUsmOQJty1zNzIeH/WTGTIoZGbEuinRD/N47/
Msjne1LIBARXA58+TlUp6F0WKbqZT2zp6c4ypjb34mjdG66rUSDm/VB7mNW7zE+J
kUvUy+KnUrbXxewlxpsh1XwD/ZMlzqPPXir2Dko4adrc4dIFcUDXBnZDIRBq6sTc
bFd6t4o8vB6SjuumI35bg1Bg6dX2QjyzhBOfJQr674yHIeZR+rFG4k9UGAVU/r+w
CK2x7YrMfcM4ohfymDnJNgoMK7Q1pvaNsDD3bjMcHbHqtqkzmEvRfJTuRs1RJiGr
4mtcnoSLPh3Pc0dz6M/6uo+rJIPX75Uspi/6mjLQMLCGPB55cpAw1ryVXjcq3N54
Usv/Afmiv3y21K4rsWIc18Ce0VhbZp5HvTcIvIYmib/NaACu5lNqyIROe9XEkr5f
qhrrcT93x7YKNCaDpwCzX8xEz2eRuhgClTURmVSnzFaWYtZ1H2BkUVyeOEIsNQwN
smB5vGrLxDGwKHmJwkjL/JgeKwf1/qxiivgMSundyXFQfZC89l7s4EAjpzOr1mU/
ggR+rwUkI7IlDQK823mARZHbuJBcD0sUci4qMqKe+sLzdzSblxgTJOpbZEPRbQjn
cCGOn3+Z4oXUlgF0/syoIRvsoUrHehduuMCs7lGHYJdB1+cdjharB1WC7p9VV6ME
Lubj+eGupdLGC8NCfV1fxA10+yAWnC6CLb56eADp+Oxpt7VC+ywk3ghkhsvootaO
1hrGlTocgnCBtAhS0Bs7Aw9aKpnvm9Zb8P/E0gRt1LEs33YjbWMNEC41/+DJgV0q
TwCnCwVLR5gL1f0J2CJl9bpyHfpcbX8Z1LVE4Bpe+L2Z82RVFhKlBUts3e73W/HD
k/dDqu9wdVY++30qdatE1Z7FwfFcSHBPNfJ+NzAR81KF37yT9yu/fsmO+v+V3NOM
yetOHmDjMKofJCXD01MKRLSXJ9fqK0lBNSusZ+fha90PheeobriD+qNKf6VKl4QF
qPGs0lTd4mvj5Ex4jRdju6yP4xBzSbFOCK5g8Gh8jEaF0GCHnfiuQK8/bQNiR1Z9
uQ7QIBYBAmLNEUI6ojddDD4/y6rIlcrwy9ThEa6mezcyJo/3VdL5DJKLrmFD8phM
GLDaXuQ+q6vt9ruEWV05z9tk6CqRDnQO4JEhwqi0jyCIpXPazXBEzWGN4eN5z2yB
urIgIBD4sLIF8PoocDr7QBm9kHG+4k7HBNfdCN21zlmcVf7mdMIRnrAvANiHbAm/
75fzapLOK8UBCXByrQbCohPrFAFggG1I0nWB8Pg7jY7rCUyJ9/as/nIQg2qJ4kp7
AalXycyzN4TdkPQDfpf+24gcqZuzKFl9f4nT3xaDaaL+/fWANGFKrj4aiG0B8ffn
T1u/FRZoCsSwP+GDqPoQMdHu6xe6yBrOuDVM3ce2+9k3x4dqFJm0jWo5tsrSoAkz
7IgS3EjtHKB2gXjMS7gNH1RHkeczW/1YvvKkDaGuX8luFf/oQrgl07ElRrZpws7O
ErxGK3eCHsTybnRcObm8KFD5rbSqrAcyypqT9uH5iPhlaN/vLtY9AxGadLfiTssC
RMyJL6WejoPYv191jEK5ZZkt6sXgtBq9yoRyz3RksMr5SLsN601n4knEwwrvF4qW
IQNsASA+uwG7hBpdyMoUNa0BCd4uTnkKyEltdUNV3eqFwvRVU5r2XqCwRyLZJDeC
MmualAsysPbkBk/WRW+QhglLMishdyxkCDBSqCU+XQS828/tuh9jEdHUMKqRiTXc
ewumtsSwdaHK7o7CtAG++EaaWOZKAp8CxRH9FkmQd3epFBDNVX+iCVV3g+iaLm6L
9hOH4YmU8jJB+bakOGy0WHruVgQ0dsCtjMdSoLNUVNCzh8iz9a29DQJa31qHHL1e
JSzJ08xlh4FMG41EJQvWSBbbKRCSO2SJuxZQRgzEWS2rwpYXDjpNTLmecbemAUZp
buCnYjzRmmCUzMEz4Iukj7R3UiXTS15TypuOw/XYyyMqIUWDNignGLHing3eCVh3
A2PCVIqrtTD0Kog55KLtr3haQcYNpy6xqRWAsCv2stxwl+aeogF2gEw+YWznF3o9
+KVkXBVOzLVhjoq24omSJNZivMirz6awYJTjTM16GL1CgeQeChCNCK2NP5cYq/qZ
vUskf4nknbfPkodRY8hrxazfhpQDNoR28Y0xJ83j0IjVktBtPDzIeWJU53kIbjYH
akkMV5ZsIzQjV97RqYmrRFRHeVMV17c3hN8lRSUdq8AnsNPlk8MxAA8TI36inU3S
6SL3zh7nJZoii91wJjM0zYoDM1U3LurLZs9sex6AlM7Olf2M1AI24yw+JDFoicgX
IIMSTtpm+zV0iU67FoYBCOYSNBP+OYX6jzspnSRTVxNdIjWcZWfucRhN7e3AXk/U
O4W6ksalYlt1uO8J/f5t8iyXLsB5WAm+Lina8P80TFn9LfV53sbw/FBvqIfxW5VP
6EPerQrking6DCJ8d8nFDjoc9eWszdOiX+3VJzgimhPsHoHAdtvwJtWNsexbider
J/BQCAbTUJG4vOVtcs/MAVfJNWQcOhcEUgajyDPhMAwQ0sSbd3cuRiKcUOF0mMWx
+zT7k9TZQZHOeiGfWwJ8YWuepyYYYOuwY2x4Fldyx3a6XR7u+UPIuJCVzu76tBmr
xoWvZLIoFXEqISXhSOvWtkrKjufwyZRwlLV4SL4ZiTe09s5eTA02hc/+WyyapYuC
3tNzTM4Ftptmkig0gia9AidSVzQjmBQ5vsfLZsB8jfc1Nll6FBGcar9gsS8xCSi9
YHipDLAhtgjFMb5nS8kr9n/8vhVjwNYy2v/Fs+Mf4m+utclWUr5xh8y75OkL4rI9
2J4yBxOyEd7DoVxrA09JkZ23FRPaqfeoaR3wGltQpWf99KQWYmMnUNKBh1JxkHQL
KEmTrfE134KRyzQ9MPjNviI9FZLZCJCcqzD1YvaBjl6XPQtRyZ1tfn90C7zhoqne
34P7vaXtoPPc1yZF/+Yd6QNKRqLUSaYxeQvbAIzwf9TPs65hKAYnhbHmhkPWiEXg
F5f/Bk0JSs+z2HC2nePgS9nHbk5+dAyUSlL0mihoRdiB1bEpWv8IkSGW/cR8zYIy
kN8rnN+X9PRUyoIqAGLbczrJYepobMH1hTtwdsqg8QDy5FcG+tei8wAEzbnQYCV/
7oQtGunrjgxln9bgWujaUCZmjHYmjoXhqprWJjXWJPt4CLvlqF17v86CVtwXBMka
ffzMD1iOb0BX529VvqKmEm+JNtRmYaASHhRHF2INHb2ZqsAritPVpop0S5j2hpTK
+JCC8Yor2H0VTuqK3t6UV/D7i96kpN0ur0ZaYFCGmsfupnsg/xmFmHUAllgd5D1S
lOLnZQVa07jTVkfECTDKVTK+6ShxI7BKhJEq2NqrZHxobA24gxL6WKGUqwRbxJ9Y
gxUvAZjxBJBNKRS5MIKm+spvT1cXaPH1xb64WbgZbiNfn0b3IAw5s35ahVqazHRI
y7rcU9GzNDu4LPANIHeeWEJKsjMrLeiaRdr4nEMGhM95SnlkwECe5iA2lm6yHT+g
fGnqzOBsFgRIKAjiUD/c8PMsn44QYO9SIO7m80wmPjLvY2qOowIF753QwgIYYPaN
BpmJxapz6ufL//VOJp60Z88hMjzhDkP6mi/qzT+KYQ8+LdMOZAignow5XCoUOrEP
QSpvGs7scFdGsG9AmvQBIvgRs2wi6YR2XF4PaOnpNBGvtHLMDDnmrx9yyOn3G4f7
Jub5kNRHpCu5+kAE1K+r2B5bHhVvIaabhuRiI5YUT/FSmet6nr599tcZxGBsB2kk
QlxQFacHJV7mTc97n20/0mPNutd5Nl+SP7Zpqcb39CvO4yxJrcpW/X1ns86s3W40
0zXxhZKQVDirg8+aUacXMOa6mGyoxeV2Jm+3xDqHi/aGP90KiBkH7NJRLNlRmck1
7lGl9fKZJRb3uWWacZ0bvkCFI3AIkiRCcPdCBYIckEtJZpJQpiHRnZFScf3iRoDc
ftaUdJKee92xrDQpnFDPoVqg5p7SVZRmYWyCJmx56WTll/6SQO3WDpBXch9MKl8p
MtQn5J/1AfTt5cJm3VjjFkrlY5U2tbC58Ddjutx4xwtaBzEqe2m/bAVOzpD6yVSW
febiU72qw62mExcZPoVbYo4ykJ95IYruRkVx1xMlh0VxL7IUXGCA3u3LwQxnCPYS
d+5ZctIKAdfMHsZMOCuhzcqUgorv9B+QCtNxw5r1aFLVX2bBquQj6zK9oxL217dP
IOp31URw85KJRGZBY1nthufa8f9Wn4H9X4lyV5HSc0Di+aP1/744n75egqkUIQ0c
lohX/8x38F6i7lr9Yu12Lqn9PTKouvlGVA1hv6IuabQTDi3v/GEJvteF6BnKTb5x
0zZl9RxWnaZGuXEbkyPnWSQEgzyEyviovPiTgK1yaJuYgBEIsIEWW5xcco6Lwl7k
OdhFHycbElNYP9NOILsRcg7z/9pZG4xoOT54Cmr5XE6ar3EYVOXUpETYTOu7KmRT
TQe90b6Vp24SLTR0z90Pqc77zs6ye9IHlvPZSwut+tQFoaG8XHQcSb1zNAAOQWk+
mTh+tO3wyXbj62kC5qT6+J04xhvpWLBR5kIZUOAZ3xUBon0Kiy26RLHmBHk9b37r
CQeHSGWplomgMi/wEasCT3tidhBzqt6srXhQfPAGqmWQx/2Wvdsx3Iiu396YtmKE
kkJDPgMem94Pbkc/tdOFjEjvObTpnRqO6aFieTWcv1qI6CWljKToPuMiGijQJrfa
m9mNJ6i+vHszedmIOJQR86q+PyqgaRfPlLu9emB3g+StJMtnQhC1UM51l8MOudio
tGaxK7hHIdFs87PCgmPgQbx3ibLqe/TANWBw7AZsFGhbHX7nPW2khSC4aEcbY3kW
J8OXZsqpLpdd6vpIvIXBD9hrSJ4+OsC9736i3BGzizF47daK4KHTgYlTz5cxH5ml
GgMHJ97wFAlAdbAg03Eah2kFLZNq8EDhQvEbbjh8uG1pEq7qc0qmuViDn1Pcl55c
/MEzmPKm3lxzFI8/bRl3jt24R2ZP+3HLS3PVjCS00UPsNfmk28WUwkMEKtpb3Wsu
ZgPyWlmj/vEZLTubkPJP7neDGSjoXppiVviEumDvQ2MKYu8JNSgrtiVqV4nwBT0q
1+EavLG5Jfo3nltfwBceVyqXzm/Kk1BtExE+6jamGfdOxRCxVnHLAh0a6zQbIzxm
J8qGM3u41phT0MgpZWYGcvOqLXVanbRXi15wKDvMvOwJ1cgW9fg/vniHCNhVrfMJ
kMlovYws80xKB+M9Wteli7/hVVbOV0V+6icpalvclh4UQ7FXekdVHWKI7NDy+DA0
n5EIK+eDANFJeuyJa6XG6WIpxHhvK5Kwxwu9JLWjWUR9Lp8Jvy09yL9zw53PI3qz
AhdF32pZRlviaUgykJJ3rBhQnUwxvEBF8DJkT5bn1yApW3YvtHi9xwfhYO/e05rX
lt7UR1bQzI5nL0GBPr0feaVRV1+JxX2KsTrARj59ElWQ++a6s8cJUXK7XSQoPyYl
eauZvxwpHKaS2w7oWSE3BVq333hEa0mI+HfWfidua1gJ0Q1W3l7CzEDmfV7FTsNP
ww/wb53Eycdw82WaypZ/y8sqJDIDfSVheQr25BAIDcgaRsS0gGu9WOSid0koarTA
6DK2Ya9U+V2fkPih/P5vQNqII3MtBgQm0UqBIHA3/6bKSLxR5+gfpUwqfY48fOAb
We8boSTq/zRlZMOGNXJXPrc7yx/thzTheuUNCk8xL3SBhmNfa+hJwFuuH3jthnI/
PD/FqR4bHh4tf/V2f7e/mDd1uLZJ6p/UZQscO/ZKnai2u1I8KWGgSAHqRLKH+F3j
mx7VwEUN1tr4R519XxMQGfbBFzEBjhmYUM3h/N0it9g/+UA82c7I54+bDmgXiL+r
hHwUhXSlJHnivF679mER3itXX+CFGTLpP8bhsKYF21oIHJU9ifwd3SUM6Yj1wd/J
T8DL6geS9ITmNPSEgNv+w+Bg1oRf90ceQxtR5RxgqyDaSuqp8ab4IxMlW9zWTP1d
kdYf3VMUsO9iE/FQgHYAQK2fvect6BraTwh1do86VWUxPYpGXxB6Dtwae5eKbrmv
d3MxeZOq6t+LRMh26Ip3Scz7cP2iLZm2mHg4BuR0Wmn4gSips009M9v4fuvjBe0G
tXb4LZ8oZH8HItyjZ8jstTFuA7Df/RRghpUEd0g70Wv5R0EUsYXGiCi696DZOfp9
CUGqKbz/oN6xZGXh7XnUVxp7floDZ3TgIg7aEg0MvWGD9a0hcjwsTEQEzy45JFCB
EeyjAd1ExWrXTCUtE2qB8LAaB1Xmf1YLjpwJG/85Z3M2fsZmPhfQC8YJ5yjBIhji
JYiob/HAfJ/KPfhfACLNu785lf8QhTI6XlYtBIGy3iq8YbE0FSkSRqFt+e2BxrhZ
q9/TgpjPQky0gCf+jhI8deAo8azI1caKFfQrtxtiqqIEBwaMFINnpnazk8SJpfJ5
AEw1YGVj6IYEPFBAUgY6RGBtKFw1UTZ5ahLqkjx81ujhTCGMws5XoLsJNO0ksy0r
O1QntMoQEUksSz98nll8j+TMiiHlPfeMJZWjLe2cNvTIYkGUtOy+AmV72Om2gadW
NrF6NhO8tXnWKaWNK3FmovR4Tf4/mnyVgS8JW5shk7RdnxbDqwRBH/XQTM00KNON
J9PLYfz/zoyOlHS5BWzr7GgDkyaogwMhe/0xQp3X6zlSOOBE8FJTK4Kq08wu+4vQ
QUsWx50jf6a4PNKEuemN6jeLk45ZEYE02jqUa/QzcdA39Bl9EfyBhv/YT05JlK7n
ROMaIaYf3szYTbEQTIPzaME7gZ2Cudu6QX53QHe80q/lvHevQ3irXSA34UDvdOBC
Gp41ihWDDlPmLQpDSyJVbOqKc8hBkcGsV/UCy9yi1gtJdK1BaU7EC+jItJwujWi7
dFKnIqXmc1j12qg0FPGslUO3KqsPMdyNV/QhUVwT3aIEgdI9n50eeKufnbEWxGGU
LYO1EBOb7wkrCIe0I0V+NAmUSuFbx4SUmMFOcNArVXIhHvLmHM890Zsd5HJpXlS6
jZN+mVj5FadNkHFpcBSXDlNx3Sqa9xCzQyWR0xf7o7lzeiXSbju8vGP1uLNb4mLf
h64rChcDqqKKlH+YylAKftIXK+8QJeJcKw/1w+oBHFAUY2irzhcOg43MQSbIQg3y
6R0dpuMzmtEQdXEzjzzWDVKzHsl2JFSRs+R6sf/F2DwYWxUMORgPgcy+2V0hrYIY
cNK38hNyYbK/Ibd5ZwWVbkiteaLFCk3/NJaKAxPQOfInzjf9coJ7ASgQoDZmt+k4
f/ZjtfNSvaaq13AIGZv0BEte99IhsBfGT5aUsRncpsP0nT8G/sQbQF8M5Q6iKetG
caMfm+9ZvLtCTcZ/9+066fHIV4A8jGorK/WNlLoFK9S73HEcRq9n/w2N0xUAKVy4
PDYBt1Ym20/RupDPrHtBoQCLQxnwwXeb38n53p/V0alOw0yGi70kkGnXIEnWC5OW
XH6FQpiMDId+5xs2HpKTxwm5S/kIq5QsuTVXDEAVW5rz/pA7CnTiCRKXDb5Xnp5G
GjGAw0AmeFb474/ugHewWuRGR8X6W+m16AS9q5bk95hOk/aokYzd5KCKL9c/s8/Q
dhDQtIFkaGiRMtPmR/n5/dyEmw9GoEay73Y0wKIOTkaALXzr5fwvn3EXRKBpUIFY
ff9TZ1WNJgj0d4kJ47VqO/YeHx5f6a4m8Gg/TQfPBPcKBCxt5ktIKAoH3fdz8y+z
VYKyXnM0jBfNMFRU4JvmOnHl8gPlR4UMVG6+RVWkg7UGjoaRJQO5IAnVkvN8O++F
jpUsmAOByPgEPLuS9Q91LFClrgQAJv2bqQPITRwe2us3jhOYZNCUdQwuyWp4EekJ
nvwL/9ooJXGXybo0TrFXgx3ANZbGTMM2xjGnXeC0amzTA1o4k1YZJbRb73cQ2DHO
pZz9OMdVF03gCHldvV26+SPJ1ofPIWlcYeg3XPP7OieSie7hUz/dN6umWlFoTlgV
NfgAnWCeAQmngZA9sVwWZvZ808mMvRy+BsKPZagwU8WHHTo7Pcu571Nga8GfKoG7
IrqwGl9vhJW3CIHxmweG2PV389DdicyAzvhpIZP8jKjKGmc+rEBblFb12nsEndcN
NBq0d4uX8IzENb67W1d2XPK5lLpo05cDcaJYETZHeexLuOvKVnd6ues7SVi31egv
qKWPjtDscVJytGQqe/vdE+AXmzGZDaUdVqsSFWouCLL2IoQJlIpiImWtJZa8D/Ln
FwPYEjGeF7UrNv+Uyj2dSJ6Iu3hsLoyLlR9GS0GdD2TwpihbhcW9eIsIiE5WDW/D
E9hVhflSAdM44ykK8r7RJq7l5vEHvXAT6fMMSXAvee8URxCppeADGVIrqFG74y5N
DCo33fSLYeUc5pZLRH9XimB02uamujkyFINX9wucAzg1qpbOWJ+vvxqNxiCR0P0T
KM7yrp4T/ambP6mw3Mt5fxhlfrR1sQhuWQw+kkrPzPMThzKBK9smncYK21660zfd
pH8B8vABxZiLF05sMomF1KvM4DcZTMu68iOdfc2njj53YBJQ0lx3172v9YCzLZzu
f5VgNJ9kKq/RMEks/s3KjoGIj9VL4Mb6rvdMtonpn9wTeIfyVU0XlswH0DFvq0qo
DqkkXtpP3PskObWAQFWY08tVC/Cu7enIL0kCjRYluPN54uLaiu8JL+Z/UqeRuMNL
KVXrZMvCvnE4I2qLV52aAsvSYaPclgjfz34Iu3bkaDi3pOTGHS/cvNDtf1iYBr23
FaEGeN6ae9iEWHY8dsrsMVshJwNyl+FDEe+tcXdvhIDllcgvJPyTo/FgyZ1LTbA4
udmnm+Cu2epPZwgP7CJfNqtOe2Y9Xbog4UEZadyrzTtsalsNMJr51yAJkNx+4AFx
djJWndOXq21i4LVW0jLMU0sdWwrZSPy4RdQbnuwMUf32ELGT1FvsENfTvgHeLtkd
ZF2brsGVVOMbYMF3e7Kzs6xRVEvH6Kq6fTmdtE26FylxqqblAI8gne7W1pZTjSyN
KWwJ1lujziEQFJXjYom9nKeUKdW1a/LHL+rCLudE04ncWLtjTqsQj3atBYR01IQB
r+GsdtbF6Dczo+39mwio50NrI8mzkHYuU4pWSO6sJ20uiVcUw0Ac97bQSOeCUCjI
obrMzw9l2SEB25xol5buh0yaoQQKqzAYIKJqwdds76OWx7+vBqSKbz6ZzTSLpdzg
WiwzwOOTa7hwp9O1xYMap3kALDbbR8h+R9Ghw00DnNG75RPFF/TwKUSNy07Pebiw
zeK09Y/2R6wxvvZw58dScfRypQ5vxFl0MDOjRjAsmRVwfGmQZiZJiRa8GtjMBvr/
vk8CVvf51zdB7qgOtZqtTwdPF//xfXJSTMNiM14Nh85NF2Zr2aNRhrlSZ/VM+rmt
PYVJoBO3LVma+rSrbpV4ZyN5z7RFmf5YWoYLvgfp9oC0dLWtLTQfgO/TtgPIq/so
7UNNEGK43LpTruh6aZjq5MJkTdXh1ii/FiG0LZdzOWKp2m3sGA6IcFZdjWD5dqNe
pHktgel2T3m2XXXl4APXaeDvcZjgXSZuynW8JXperbNJ5l6uLnTSjq3Hu19RUs+i
PwVfIAheejiUa14eIg7NBV7W4ySOGQgJ/XLQamvgLQx9VhoKSfzQ0pW6ErWO/OVf
3OSOUWh/kaiPoSH5bMabDykyrFk88kI9+tTxDYWUp3iPsbl6RL5VFgJuoyOcqxL7
buo0S2tScmdoTvVKQCRObVj2hTPJG3evzUe7QXBRdJFKhRTsGzlCuj2K9LovaznU
NHL0Hm4g/ydgy5qCD2yJJRu4k7gj3hZTkHQ8ZZTUpx+pgiMUtmKIrN2OfJhSCOYd
QOLLoIeF8sO8oyTUkL80w1Yqa2STTWiL8HjBPXLgW61jClrD6BdBfVUxFvvU8VWK
PZ4ElkoTpH1CD/7OLgqdT4yLFYb9fUPDfywsHqfQAU6Fy9sWPMk0slAWHihDjP2e
wr9pDxZwvuW2q8Kew6KFJPLeEQ05lecpM1+KKHF5fb01WbWq7cS1UpoRQqroMAJW
XgewioSjvF+tppORLspN/JCVsF0mu11qQK8TSrgzSYO5iRcIg34laVP1tADensEo
V7Scqzgb/0C+PQBXW3/DGnoZ+b1CoIdHhrBAgTmDRhKmB/xBREyR3D8spG1+S1Jk
oGe61BWW6KmvkiMw5AstOGiF70kodIlpYZ+H+KpzKsifkjjQJ/giktl+dtTI8sLS
u79kOV8aUk+0NHG1/Mx1aGRFiwvSIaza6iLgW9JgPK/xmyyA8bnDd15zdSYiQRa7
bVUZuc/BwtDK69Au6BXOS7GHioOYSj8jqdY6K9zVWh1n/++OaNu7fuiq1rOtvHe2
dmVsUqAa+kvC1e0ksryZN62sBLbcbFqVytlzJM7TVE8olkLh612IyPwuklqLH+xS
GbB5gFbp5Qs03I+NQdtPKhEBHApbLBY5rchd4KZ336qqtF4U0dmYxQgADgfuZoQF
AemIMXGaoQODOcE55NTi4/kJJh81rRfG2RrnfR1S1XMxlwJE/TSrisviHRkEY9ym
wZMW2iG4chCya9SeORMIPaRbsbR3ELhj6hOxKtajV7Y4Zmkm47ncMXEGk99AKtF9
roSVA8S9Ds8K8IwxPxDd0/u7YGwaez5oaW6j6OpeSpuR61rZC+/1VLW3ny1I9Gxx
+2VGNkLtlcnnhySjNhhevbnx3jJ+GKtm9fjd3t9lpFj8Rkim76DpkqG2BG6h/XG6
qa4iBpbR97lum4CG4eu+llHQgiJqaw7I9P2LMg75djjCss/WTpZJvpOqmjYdAlWl
AzNB/khEBlrqjoycmVdmfJfT6wOJxQ2uw+LExSQE7TJpzT2fEpOuCU17X5JFnIWT
M9sS29zM9oE4Mh1kwR2E4ai7tzrNpgTbcwEx9HbB5NjiIGP+t1/8KCJ1ecXZjoyh
U+d7QFD6ozk4GUqE/HcTYt1aM71mY6F233saWLi8TVzkYVG0Br/TEpBOr1cmI1yo
qyIaiYUw/z9Y91FB5J/N/KBH6xUzPWiDs272MKG0fTaAZ44Mc4ZycKDKArtw3nNa
3ruN9mGjcDoUbDf7Ho2AUyv1LvbPwTfX+s1/PVbCdEYrpd5l7tozH+ACb3egp3pj
YuqCHqoUf5mLZ/axLdmNir3wI7Sa3t3Q71bXNjUezIgpeTNyhYdpO5qyGT2L5P6O
MEUJrkx52XpDY3ZQEpl+NR5ZQokDwFHKUQ6zhdhrQOVrYET0JRw/y5yRzLMSw8bI
8Mt06RIgV1MozJPW+udLZvCsBaOGx3S0bU7iescjLT7EOvQcwsWebSo7Hs8o8try
z93C1cnHOu0NUAtWQQz3vBt6Bxd6yLIhUSPmdDgB1cobiTHDFkGloIousqC/DbB1
3HgOl4pBZkYT7ysgsKnXH/pH1FIeuqUWPrfCsYAeoAC09O3evUxJKY8EDC1Pgr6D
/pmcwvdzNk7y4ghW9MUwwCFm8PJuafgjZkH8WVyrbFdMk6zftgFa0kOI9XU+PjJX
qjrfYWDYNb4lcypk0aBjDtwfv2Og4Dk6cAW1gcN3fM12K9kTibVcTXBYZsNVoaIO
V8seI2DEYTVt4Iqt8ZH6igSQB7xR6L8qQ3e5W0Hl6L2YDo49/bxpBTFhympoesGQ
HENvYuGZbjz9ka0z5MGdpQ0FskG4LsCF9vz5ZrebjtZmYz3KtOoYKDPX3a5LbO/b
ht4ACDzQGVjVlhivViAixcyPn403YsA8IamSlpFcOr0pl2s9/apX0XrBhxPpMn5i
swT1//kqwvsApFYKzsVVI05WuWKW9N73b3o+7MU8Pb5/L4BggfEfT4wI+E4vUgI7
ayl877QAR6VU4QE0djsR3Oz8Nrg9FYEqxyJsuKTAUPFXz2x73EnLUhDuUkHWTiMu
Gdq4z6RwWXlnlNjy8b5f833Jfl8MscEjFYEf/GALAqL83y4vhSreRzIGE95mw/+z
D2TEiEVHdhr4khbqSaMTWpP6Bhg9EqY2bo50XQswzHFvJeV8jbe76g3zQijVl1c1
hVUCv3xfBZSppPRv14Nfz3o3Iy1r4zj6hvW6bomGHdWLUVQMkWoMso5yeu3oVosg
Br3DknZMqR3B+nKgyvZj5udTkIyZP7y02A6DJ3BoPgyTHOYNQjkIYCBktfvftrem
UBhdLljFyvsipBDSpr03ayU6ohtCMlTXVXCkzDzEy1vg641vp4xKxo8ZyAwqJN9D
za6C2Zn+mD52QlP0Mo5HFI34xHDyo/GIE5lZuXS3NG0H3052+UCpH4ODmy+f6R3B
WOaO3vbL3CLWZn9PGRXNEhc+Z5O3aOCT9SwcOikDrqEZmtMQaPm31dssHv3ths2F
EVoym0jRB5K/ycebAH4rEIt5w/F2mhwDoZKl+aN7SiCU5yNXOFIk8e0b6UvZIqoI
kLersvICy4HyNfrgnnlEzLWQdiI8dAnXJ36JGX3UxNSSQvoKOv1qjPbOTZXaihKu
QjMo2e8s2tvnXJJTudCo1wv0jiBPAlkW96JW/UJBnPzFLTt/LKhB/2DvlYiB/DDX
iHEIXkRCeD1xTFX8gOW+KCx2allMwP95PDQvHNdsT1L5IWOkLn3Jb0wllgtoA0ai
zAA7rqFmsSMeL/CQtfjDEgNQ5oFgjLMYNvb5MBlms4APfLnW1saqCoZCQTP5OLx4
DMUTlr/qdCz312V+AdQuq7/JwlVbMQgVL653wfoucptJbKJAF+W5BAk55f1pFoXm
CcQdEGZp2bpHaSt/8i/creYbzlRlDbA2sLt00oY/JkkAuvaqlDDZgNLYMSGZQs3t
3Y6WjJUR8lFxRdIK5Fn6HCh70MJTbEWKYnApUyZcSOguOMZtz2vzvN8NTSnM7tZO
jIKSD47boLu5dHLXxy7Mfg3P9TnsGRjdxnIqBEpbTE7F10DuxzUQGwva8Lww4KVD
kcdnj7Dw3ZGKM9VQo3BNIkGWwFGM7IcOHDASM8qFvVBp4puCPT1Semrw8T9jN5ny
nD52gSVo2URWe1WcssVWuKc1cinDDFQbbo58e/apOlY991vH+N+FiXUAF4nMOc/3
yRdtHAWl6YhTrCES/QRhuU+cOTyWsLN0yD8Af0mOmInNBopmC1K6Lm6oYwbFTR9v
2AGuXpXBqFnBxon3hHt7xfk907VVwufxvr9rJjIsOhzzLuf6EE3N8YLVjfb3s90M
r0SSwLQF1UJ9W9BLLwKi2FPeMj/rO3NfVmofS+8mr+yRzJG4TaBglu2uk5b3d0aJ
dEsrvjIa0kGyDpl7HgwfpC9++v6RHFgfzRPetMQuZXSFK6kD+ApnsWdaIggR+7ux
gKy9BXpjGvIeM7fAc/44XWdG5Y2J3azJdtufeNPMkIZJcYwqzB+o6/bkft3zoA+u
3sUBtmmI4pF1wX4Mg/JFDFjeLav6HvKepNesQU+g9k8eOVISz2oXkaQAYh/CjOyx
s1M4OjpVMFhUAs1UEmHMWOL6If6WJ1s/wub0tENwZql2XVJhrSK+wODkPsg1kYKs
uwJaxzGGGLRqffixeaSm3FBEy1kp7YsLu98mUewjh6l0GGgGF60R2mipvkVbg+K5
c344R6Lv10L9Jj3QDQOuy+i9Gp/nsN1C4bdtp83AjdxPe1b3ESuT/oEU5EEFSZAV
Pd1s05jZel573Osl4WHzde98mopELl67hf5kr3DgFY++kWbNF7T8cVtnyz8vx/Oc
qras9hjvqYnEBms4pyuT+zPjY+JhVnpbyzAXiNBX2XXSWvyPc6YPFyepwQiAcoOw
r+600DN4h0MBXUbao+DIIQk4USJNUkdTtxtY2E5CCjEowFmomguNmjxzOojiaKWi
ixH5G6yJB2Q6/8fQ2SXuGfrHd+9t2wzVZ81G9fGfalDiuSFDUVrpk0WwGN718f6T
nqcx9Awbqc616pU49Vzki65fLLJ7Z8h6vk1ZyBwHcj7oUwOrADxOOieE0P6gfOfP
w3rKbdttFMvGc7GThZvx5TJcQwUk6MUvtkRmcnzkVg2w/z5ItYGmnd0GbB+aSJD/
lY5ycJdHYtOn1jnCUNlKhgqwrSXxnqBJy8/PFSqL3xiwPy+1vdaTF5H0AxTrLmQu
beOOayfmfXpmgri2dDEaZFmzjUm121Hy9fwSdnR7MuS5BNu8MeZ/ujEw2yaS4MP+
GasKlHsIk9d3jJ42n7SRoU7+m7mJ2KIZE7WxPMZHec4DjO7Z9EbQTD0m4+y9mss8
KhRWbzQkWe4eGvS02PHJM5UaaN+OayNH61SmXyk2jpHPJNpXyiZnQXIP71Sydjfq
UpD1U0LpNk/mNvus3KZoMuyHfb5W+wTOL/UdLanfnxTw0OHObsBDGxrqyoRJOhEI
iJRLsTPJF35Xj1oLErUtN2ZW18PD2A1tWiMRO315yAvEDl1SajSzg+ctdncla/An
rJmN750QAndr+GxAjJtsCCQnXyu6NPzIQE+vlDAaz+lKB8yLGslwKrNZB/iR2UKR
S1CPMCkA1JTrmu+ZehhRg+3NgawCxcOvUaGlJglBwaqj7S6AP/WmSUNE94wc56c7
T8HLLjx7RA/nCuiVepW6C6vEc/IkTwbIvZoeyqFzn2xl/CeyTrkDSMk0amJU9xiy
yhfFidxXUZkmcAY56d9LyLEsITfDFn3riq8huo1w2zWxZgfaoQzSc7HXuDl9W6x7
xbFMgUoKvtodT4QER+29H9rW5g7hTUbiCozcIMrockFaYQaeLcj4ZOmzN021vfjk
Cj52QvganfOo/SuofF8tOU38+nKI+ghTLq2pTmdUS8RIhF5WyhCYWk1G5KP4lQYy
3EilG5HVUcSRFcBDtn9M2RXUZgYblL0f1goTJx7iL3+HMpuXnU50tn2H4asY0RjV
5TX66ISeL05XMNNmp1N6u1gsjAnlDKRiKHGaL7xpZpniKPgGjdhkWNwXnMJVlH34
fYV1MM3veZ1qvBcOL1y2GDZwSxIitaGBRluYtjw1GbComvUy6bXV4Cy0eM+bACVm
ZCUkvMQy9dGS5obw9uYoy330oRcrpP/+BoBatR2recP38ShPZbNiL6A6eOe9HL8E
g4+TpYF+NERGt6x1PxjJR93QdGwqV4YysPoCYqV9WwFnWEClfFMzFC4OyK8X3pOl
+wbjfeu47mPcFD7EV9B1lWoUx2/KnGyBNnh/g8E/Jbds0cd3R7NVEu5fd97BbwX+
ZKvRi/oPzze3G/Hm2LY8taHx35rvBm1XiWgPUMiz1Bc0F03Hr0Xl9EcrH2lB+1t6
pvjWONcDPLNS0kIBpUReSqm47JSZiul4FGoRYAZv+19iLIKjuxBIpCy8fzcr4b1c
SEwx0lNr40OVXZWtVdy0P7WIEaJfBRdeCLNA/RlM/92cLPJHhd/2XYi3RwsfZ14F
mXdPQi/f0ylNQ3RWmmusuU+YVQ+Gwp6gOksNxdv23K8yojPdZpWciGF3zUq97Eqf
OUiZADV5qE5AeSQxT27MvJrvhMblTAeVfVTxeYqCPlG8wSKnHvGXUmaHIqp0N08W
Fk/8yceOcOLziD3tE2QaLDjn3csU+nT8XrG89KwXnLaFg0cLXu++qAZ5QgA6Dx2J
MCCQOLpKya/8B3/OTLF+3TxHp1JkYtEIX9AjE0hg8JVxzv3dvDgdEC/hc1uaqFpS
ZVWfAjCxi/lAVPZYi7wjdK1PW1nXIuGLmaW0B7izW87eBdvxkjpjI2NDT7uuPDXc
K/+KrncNsVIeSQbTt4yCBRNazPcd2ypCJbykdJfC1fTlGFZYcBZihlsjydLn2H8A
V5xiyA2NK3K62Z2r4uC0yOSUYJXAum3FskhmGx3ZlEVW6fGIUv8sq6GE9KJrxuQZ
Rl9xOhV17YqT6Yp1xvORbG5AEn911VAyV2r2/NuJoYjrKvzKpG5LTp0E0bLW20mk
1eRulk7LDE9YEK4tgnEdKu4ptfwjxKw/XDWrWbZSibLlyWm6ewj2fVBxjfOFmrXN
Ojfo+uNgEj/jMNsoIkfHlyJQtOVstwSxGV/aGANyB0AEzOdSy37P32RWjyTiPiGZ
QuhCf2Ba8kWpQ+xLLyTNbqDrmDheKfPFzQsznpeBKKwwsyZC0IKgJoqgQPO0EKTl
1l5LrRwRthdryNvQwT+YD+74KkiY0PpipchDkxhCkVeAb3V9EuQoXKFrmTPlvY/j
T/y6jNk/W7+e9FbJRYqJpEAZx3Ib5Gc5P8zR2SW5WQhY+4LUl5YRDEeG7hdMZeqB
ckfn9B4UlqoO6lXd9+q39B2ZnAR+MEF6unWR1t21zH3JthMvRIoUzFihQcaenwtH
xTDjTGkFuvN0TNhBgC8XPsQyVzZjkJ7WJ28DFCnMuUVC6YcX2hZ+IFX/u6zwUgNS
IBIc8TKuS//D+WRnXDWfAi8UfkdrfTYA4RUlswcc40/HMO3rw9oTJEb4u3gPW4cL
+UK8RAxfUBZvmLvUsKfQcI1vO2NNbyPRCr1Gbyp6s7+1kddIVJhBtG8eYbk7+sEA
6efPdEnnR+YeqC9MX7hY4EngfIi9GUr1q84FOJZi5jvtviAzFB/BFK9ARa/1i/VE
Q+ZKwKNEIypF/OFyvCtrc+hdWhztUdVbX9r0sa6Wt7Af6xZ0SuoSagK3F/j2sDyb
k7NSY/S46uvOrJnRhs7u0MJxU5BKOMi/O+MtN66Xjcmidibmulqc/kZv8EpX2SdV
ie3bVTrr+4M32zHCMEUqkr9plr3T+yJ6k3ECPlX5mNA9Dy2IYTUFnSCwSmyDI35c
x1Yi6R5F1cCs2aSLspNGpneuQyDU7YiX5Vy/P7nIVlaGMNcJ72h1sCJiXwr2bU8u
FmIodDnGnPEIapoKlEOVsPxtOaNO3MPigQwweQoTahEvwio5m0ujftcRVbWWVAct
7MGM7+srrVQfOzNGJ5tVWRKk4HuPpMK74GQxTndXOsmR/XN3MtAHiJD4x2nn4sf1
69lQU/TVsA2cQwinwXzQt73x+51TuNwo+bRmvI1ecDJTt0ZPt+6Zqp2hqSlljFDL
h4TmB7dmL2YXxaBKkHKUAAikZFwEyKltDW2dYBXwLghEO9PORnigJ6mEnU5SJT4j
kKdVxqok2gHlmAfV+u3I4A8UlOa+z84i+Fc3WA/YgXNVN2rRUiEGfsWl+oz3S7BQ
IbedxYPaJhvx7lSuiBea28W40KuaUI/Tr/FwrLkY8NQ63I2p+3Pj8YH4L7YiYW9r
os7GWyyPHjp9N0b0E0B8H5SeRb9nCxUohUWu6CGciKBnb8fx/8bNopmzPltow6e3
pHh/Mwi8nfW5aDcPV7PwR+/xIPTLyLVgcliokyB//m8XF/mGmttQl6brRTlfZB9Y
q0TcYqZzxP/HeALI6CtAY+pQpYBbm9bgJ0v28R/YQp00NAUW/tY2GTwP7pDMeI18
Dgw5j6DHxHYeC7l310ne1VyGCuUQBzxdBV++Pv6fteyOzos9FODnzafEVckD7Oes
zjof4VqVLq/xRAamOyXeweoTJ5yKblmxrVBbnaYhRpRte7l2Mj2jf5acVWO9IJrt
kpLcHnWGPrD6gM38kJtrotol6V0Q5ynm9b+KMAWtaEkkrPL7IS235xP/x7n4GQA8
HOwAsWlyTdzEkw1I9238o5xvBQMY+s+oMAj2eh6/0UyQbQjURVOSdM/c71rhHckE
vwTIjGuyk6P5G1o3z/64QEdwDf9xMFM/KeVQ+Ogsq9c/YLLvwk4qZkpazQatgyP0
x8AcKmYKPS5iubuq1M3e9bmevUWjiIecisJOFyErm3npBFpBRE+LLvzUbGrQVzgU
TGB5DZuOPp5oTlgGL0Ngs1WyvyZ+1cK7na292TAsBWovueedE15wnkK3xnA1474Z
0esltOs4UiRyVgFKanM7f/mQmcYhF7Pdwzo3upIPvX9BkNpuvOwOTnoinSbwwHim
9FwKHmLZdwK4YC2mMtGjlCXFLix/7NADanlJPjyvRdq5CKKC9LSETNOkOuasouEj
mq7qsW7WL0TGrYcpdSD0DkSFyh22L2KsMeKrQSsNgS6M9f11dr/g3Q/UbCREEKFU
jIWDYqs8fOiTI9+5ULRgUaU3xwAgfHwoppQ1Ak8OJVAwRo9Bspt3cpiWjdXwtk6w
Un1D++pJeag1sYlne0xISsJ6ftONmLorTM42Bqs0QC4VyQHGZw5/7xoWU2U/EnQR
eawtzSDGa95VX+sCph7MfamlCMazMF1IPrwT93kJ+Y/tToQbe/GCPuT0Xj/+SBFP
h7GIhZ1FZvWpLL01hNPTU0qEHv2SpGx4dVmkPNnZQk8kOAulhio7xZe9JSacup+W
RY6J8HcAwNkg7TpJRKfcrZaPKYOZ+MLyqdykC8t3yNlDnvk1TeDsoYcS9leuOP74
w79cZzNl0r913c/iegOhdu/VgCPVCgvK0GZ4uZOyTjaQY/jZqdp4UVhqgzgwSehX
ixpJSN05qEYDVOZXrFrw6CSSeagbXh53nSPjTetladMa5pyr6bKSyicqoVcGM5ro
71jkWMp0TpkLQPk0H1BEKtkpfMDBs01TKYT28iQm9IZxNF3oiQJG4Dns7oBPTYH3
M5QiQsbwe/mJanPDYznkDrgRnrfsV6myWI8n5P05aH/ZfBImLyOwrXHUHp7nva2U
3nd+miDYGlVv+mXHo+G8y7kdeCzx7taPORVeJwABb0h9ewK7bE3X4TT04BT/Lusi
R1GEhqVmAkpD1KiGE0VX0Gq+wCKwuhh/NHRfdeVdM1WcRj1bB7Q50md0qF1/iJnS
RjUq5zzXYL0t6vjkxeMcpKWwv1eWuoglLPXlw81e1zLW0Ks48O0QlTp7me7xejLf
/as4k9KHi99+A8KbNIZUHSJ1LG1WU7t9ZC8HBATdyavAdnVSagBEuZbuCyvZtYxw
EV8z0KmFceV6cpX5+VUEk78qU3b9rIHLCVhiG/Yht/+fIm0kneJOxjatjthHOglt
OQp8ex7dF8RLUVF6FZDa80hl+q0FuM8g7XK7+6dHNBSo8j+iigpxjdWCZI6Ftaub
oyPwvVXPALJAOpslbWma7/LxdaEfec+HiI7rXDwnLjZ38kQ7OIdcd5rCJK3C4r0d
YyG5a7jV7NvrWBi8znvq60RqLdCH3moWf/iQuMguTr0Y/MUEl3Vq1A3IQHEdxB9J
QrH/ggItqywcLAmCICxTNfTRXdlGWUfREZDxqlrQFG3haxXL7DYdcW4jeJmyNkm9
Yz73rxAOPA3fIEvcsv0KfWHsYEU8Pi8nmwc4erbVuL4ymK9pCHLeLxOHXZ01VYcI
S2gion9szkXN6bRTf8oTM8pfypDt/kwDfc6eklP0b//pFq1FUYwigMn0NHswcR3e
KLLZdz+3KF4EM4Myq7+6EW/3RJcspuQ8xFHk9OMCN7SurLvgxH2QlV+ti2QxPlBk
n69PEZDlxnv2kpZCbyHKL6Xaj9+lEnhtsnhAQ7Tkkn8FHx0CZ2WKdF/6axlcUoIA
TueX2dFB17ePD/RgUaGEr5z5YcAqnpk3Y++OKLT5DP3hHzjbT714NxJWoIcf8N2m
vCBpPoBVTufxLK5EPZxh+pmF8wHxTT57ZvluWLguS2vhZW9toc8NupaIq5SGEWGT
AeEXfiNUFQCxYm1YI3knmhM0NHpJFyw2/xpj1MuG9/qID2ECUrB82ayfbKj9Enht
UwlFN93UpEreaCuG+PZkOBjNPmgPCQAI5G5EZU1jNwfWczHYriR4/XNW9DvnxeIm
a9FvTprV4fGioCT3EQWwL0qbC/FBrIVBUaSHhSo2TeQX21gypX0SKWJKLbq43s+b
/fDQeHv6Lze3gYkjpLiPbAJIkEJDM995dDC29W4/KM3gdlxcfFrmMClxEeJDZg8V
jBtvcyXPerlwZCxCXTx62hvY6fgKYb1onB1cF5KHNtPTzOQQZlVzWXNMUM/41QTs
biyTLmPJEpibZgwVamYroXO95PcA+5IvVqM6PGzXOXsPu/b1QJMuLy5kwPdOu+sQ
B2cP8XIBn2FuzFuVXXDss9G7g1rEqfUWUqlgjSlcOG9slCU++kHxQNGnclOcPOfi
2zmWMe8v4MchmsS3zkiYOyxJ9StN1BXrguy8AZUJqKCvElvsTszVSEmp34IBR1uK
2Xc7mx+Spubhy71MvckBjdA4uyXlC2q7vYkxNEUvr/6+F10V5CqehX1RQfZ726KJ
G9n6G+IY8s1SGEcNx5zzqml8QdyXB9MSDTBVd1cuxgArWfFCIm2N9oUh0X/VEbCl
X4NsZfk5uqvLWLevmA5ePxLtUEG+EULT3wzjJ1H+CMedHqjhYVeVw/NAKpze8ToX
w6CfwyT+D33GvE9CFgP1L8CrnsQPug+AMVuYuvdXS8QEMVlpccH0xHmgmvZm4m0Q
3KK9D8v1rKYbASK4of3RGjo2aux97Fj/DUJQhEwFBemGSiIFhLLegnDt7YJBD962
3V4Eh16zi1EbxnbXX0RoloWejHg8Azxu62gFO4eiu7Em+M3MundE03ExR56Tj6EL
c398PLOnVeOHJ49ZhkEjYWWUBrtHpCnIuoR4Dg9WzdWC2IwkTjSxgsua2zaZoshE
Zja7Rh5gIL+x8JlGRXdxZl/UJewo7twMbUTgAS/t0+zCrarzeduYg03QuLJldEsQ
gHn44N4aXtqhLCNn0eszEDOwd1146Vnz+w8MmTiFhJWwQMSQOeaAlOvsrnNGFp3e
BAhBwuCyALGzGx1lz5LgW0g0vyYucBkFm0a5KhkC20txE9Wh1FqDrCjuM+9t5/Fj
klsDSB2XCmnLk4cL2D9/R4XR674tGG4bf/SGNPC+B1FxVX4oDU/L2Zz8X52cHuEj
xhc1F67L3hS1q6jBjXzJBR/KQG2S8dIsOkHxYjvs2o70Ik+T8xfyJvrMJZHqR/KX
+M/vW3qXMQdgdoCNgrNG9QBwWXtE31MH80ogm2yFYTRnOsQ9QY1oYkoiXBtvKpd5
9ggT7TGhf5LS6vZ0upkgt4sVGtAz4FYfN8YLc9YxTOHJ6gUH7dXdQFMsMLQkq0I/
z5He0DFnsdoswQr1NGM/YG9tW7PcaalzqNDHUbSN2ntZBO6aVivweuJNXt5UvNJx
jyj7fdHbwdtIQhWe47Lygf5VuQu8x4s+cbhF2Fww8oBGeCjVtQIfUi5fiqv9LTe7
5AJFXad291QNly5LeZRz2ZrllnOFtIyY5f9Kr71e+FNYCemwzbBC/1KfMADVj8Gi
R58tMwAmXUmjtYKMjRD/5deQvTFlrfOg8BAjea6p4bPggl4fOxRAmdtTvPyUGdrR
v23HYXhPveKcMGi3Olyc/V+cAom+ih9hjtmMsIbP9gYthWnUIzrrbW/e8zxlkPyt
Qs8cYxFWiHMM9EK4CkECZ5WP2RyC0wBuLS4mPHsNJnG6SF/q1EVQVEOUhmBL/UF5
mjWSAfWqWbE8VTAhRfrwtVsUK+qSSuPo8Ady0ie/5kNuoB/prwt3mJBmC8+hcSl5
YL8HhqhwVxp1k6kMf5d16KiOFDYlu8gi3f4AmvYXXbvhld2sLfr3js/LA7vg1g+H
mlQKp0bgT45M8Wo0Gy9WsvaQdHWOjTxD6KOtHQPutpn5HjKXWrLCjuUDCCiXcR8U
Ym66N24+MY1nXP9A/HKJ02qy99J3jJG6l/7y75t32AQJjF1IDMObGMjuTep2rhTM
0fALyTfGliHbl6COpO5T250WrJxX+jnP2s4tQULzN8nAMpJHdVIlEiZmUUy38tna
n1LZdXNeAosPtTiBd2DkpUCM38B1GfTQgrbi2JtNvS4vxUD6a+s3aSUX+9a6U+2B
Sbz4kjf3caEI7pZgVWlmQnII8PGHZ3YBWSfJjyyH2ZA31bMYfQlLPySvdcPwrj/v
p33TtHjkWEPvb4Ayex3p4KrL/LM69ZESSB0tc1HaG2BWY2N+Mm45VBTu2g8Y43zw
tFfhIDeEPnARmGgjW3Mol3/RHMRN4EuZJ+MGCSm+qSlGVm3ine7V5TXZ8s21jVZm
XiVNhgmhQ96lr3ttyG0rygQrAG5BYYCFw6NMVoVd/C6bw5ZgG40UKCDgDyE3ehZj
mFy3a2oPJG2f4RWRFqDj2nUu2x55WTyM9G150AeK6HE/1dJvgXRZ5dnr1N8PA1Iy
kg1l9Y2gk+25CBTWjknaTxJzqmNiOWH8ttelCbi8ialt3A4Shivv5nNE3pQWxdrT
HNJuwSNkRg4PK0i6Frdj5VgOp2/cHghDCjb0vTSbayVNJMiYen3dLny7YAW/1gWe
QZ8nqA8FQfIoDB/00aLjhU8pD1uc+S6wFKG8eDoH5V9AxDap5ffjS25S1yO2WPZZ
oBVAHnKw7pAwqIEhaeEoqrF0FzCZGfpnYIAxI6mZjbMeR8gFZNxWyal0tp1kKKKZ
1k96jqJIfjdfIs2aeM3id36S1jFFxYNha1dfHty0+pQ1RJTpkCovqytf2Dcvea93
MEBzBn913v603lLt8lgEgoaNSLkW8OQsLyW1CIsYRXK1aym/xXq27JNzHBkfI41X
MO4RcDnKYnoLTaZpD9wuc6h67RqrUBwA/xwkFYLsUMS17LU979um596ZV0+FNugt
VcDZ+8q8C9HrLRadf31NnDfQS42ifmPDVvTKdgQTAiu/JvtSkk8vm+5DsEnKvX6f
G4SXA5VVmoj1QITxKqmllkoRNqSwJUtrzwjwGRYHPmzcQnKdgIPxNC2O6iztILrM
zamYYbUT7fPh8EFCADtpMmsQxUGTr6xRfnIz381RxA6yfYCvBLVDUbaWT22QI/au
nlCIGKXWbnaDE9rQVqtYzZk7nV1qvMeR1Bnr7UC8ylQEIqVMoLGW+mtDFLu9DBiC
22j4iXLGxpGG0DqA593RWtTztI1HgmYpbJxG70KOmcE96fHwOBBfrNwF6u2ohS5u
Hk2G3RMI6zyrZpK7JigcEaJ7YMN9MxScXRjKnc0xuKsQZfR9lyUQRuk+ZlxX2t1B
yi0zOm6k/v7UHYGJ5KVE+wu/Nvi8/T3RFGpWEH4rGB+YxuwDEAL+YPJrcSVPAoEH
2k/C4+C4XZP/j0L7kiameiadYU7Hsvm46lqUhyvr8H1sBw5dgfZXk46YkoGUacBG
AXQMhUYRpbOy0tKb/P0WsiIUNLGjj8mCmW5zhwTPZpktZbXLkdW8YErWDJjITiRv
BUYT5Y41T20iuKKYUniHULK4W1CISBEpGxvYQ3tq7fWrM0kVhdgc92jtFO1hTrLC
>>>>>>> main
`protect end_protected