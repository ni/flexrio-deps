`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 26864 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
ZIICkMu+S2rq/yOQyqhpulo5ukDc/tRQVITd5MlhjyIeKeQERvpJKDh2ouKOyT7f
kNvHJxU7pojY+iuCiCuWXZAhgu4Ygs30r+PVwhGFAkxKZKlJ57BGpb84OWBQ1ZNV
XeIuETrHu5+9zDW8VMbwiCbKCbO+wte0r3SmRHM7xTjRkrBMpE8zvYhFURy+p5k8
75/KCCV4wjXx+SFIWriBAEGAEyJuLBoBqXBaA4wGpbc57h7gUTSqKBMPKsXY/7I7
2x3WJpr+3Li6OVD0K3jt41ZcK1myfCFdAmztrZYnDJIL0JKNSXM6kQgnZmW3+fZf
ZJGOy+AFNCNWzL2Q+PDtbu4Z4Hggy9Q4hfjG5h7w0tqorzlZ/Xf7wNmasiBkgUx4
UjNz+gSgmx7XbKapBUeR29xjcRpC5/TR0gN4fq7ZCZ8PzdMR6eJVAl47T4T3yRdp
2tmOOERbmBdDXxHYXufx3mnbltzx6eVVEul92Qh5yuprHjBhFEzM/zlC6SDvDPa4
tsXIjIuSXtDrmZnNH4i5Oa9gta8Buz9YvOGXFRWhL+mr9pQ1Q2AnrA7idnCZsgBe
pd3wgR+1FgalqJpx7vwwuj6rmzwj+osDQRgkyBvx2NbLg7J3OLmXVcPFnoV1ikme
BDQBFD/JBrclp5dRuBA0dF/NMcJq5wffaLp1zvl6cc9nC6+IOtATSzwjL+vcXph/
gI/3RZyHI0F042uq8YmkFjfK8XgUsKI8gWJVt82VxvRJM4v/hrx9mTfzxVArvcmt
3kfDB2oYj1c/3gnzJczcSeIOJt+rIwbNpYjGX++RHh5Yl4VM98Jpu7eccSoRUI9V
wIFAPLJtuirMZLSSJIDoePSzXrV5MSMlr/YqBfl55B9fme0LqqsJH0zqVtNDzk7m
jv8NnK7bx28MNk0FBTrqVCgBKaMwm0baogfgzllRtvEw+e59haVTkm5r9KqP/AEI
ItMyKBcpxzwhHW86rmU7GCs9IY8dtQYIG5SCpHH/sTtY64ZymHV2+z7VdsHIgHSz
TkPtsBibLaePZl4IcaWkFW33sDHnGrX6tNQzArFYdhacLSJU35jHjoNQM09XgWMI
zvUYGv1IQD6XLae6rkFDXHtkPjv0wQ0grG01F7+VCd0b6pNY0KWhVQskEMNfXntY
5fdM29uxOfNsN2XaJOmTHSdeFR4+nGy9jPUNMJRZw3MqcKuoTrI4n+pLhqGGTPef
jPyeCU4A2WR8dJucUJqGPT3thdeXFzkInVhtKciHv7iimxwQrtNhKEhhz7ScJCbQ
b6ffQz59NHTEl1Xr8wN8NDTvUHZOFq4selU0iucS3PL0hEYK2CXFR7hwmh+k4kKC
T2eMMh78wQqQ3xU728/2JQp5i0PdCrf3wQUJKh9oSEn/AXyM0npxvklfbuV+kyNI
9C02ZonGUvbGYn3VjxUKYgsnfDfltidfbclRqlMiMdYCjByBu2dx1D550R02Qhef
6WiQdLBZUQ/4BxP7wD6yvgZxkZ3Ribc7P5EaB0705CdYntxfzr9l9t5mf/d1Vdzw
Wn6u87ZIgGfnW4HEUvTV5zTd1WIypzxqduSRoCs00O1M0ILkhqY0tZfvwl2Nw1t6
s35cmh7iagClre3pgTFDJ11uRsSFfuJm3PECcLxl6i4Rbn+gjQpUlkaTv9RljwBk
xcP5pX9EjCqr32huF3VDdzI2L5Ofx1627c5gcIn6cH9t18h4c/dnqsrLDD5JGAMh
SUUAIrKCpYbkMpnnAj+nt3+CzlfemDL4BauaDdJf6u+Kbb68BQ+yLvOcaOGuauj4
73Cc4YobxyQs4iwwxV8dha+KygCL4HdHgPj1RUsauEeVfRU8zNU94pwmmEjV90+l
oNNxX4DknwvjR64hc7hrkWNO3L/+5V12oWbrMQLgAZf/uksEE/wPbpYkU3vGwfPP
JWX2Z9Oftrcc80W9wYRWcRJ/MQf/a89Lbrd6oKGa8pkPmjLJVRXM149bfbwisytA
etGXzkdH8+ES8OBNHkUK4GPVbuhloGaB9indungCDcRa1FxCOl6e3v4rLnUDA72T
7yeQUq7fwL9pyjwqMeMpgW4SV5Q3KUyD8OztVhzfHgpyXmWM75qA6793vFkY1Rrb
bBSX5YQdS5RUZi1mKsJUk8jWwi2d6zXIiZ88hmL/smC8c1pFLiDs6M0lkiJSqa9r
6veCZlLstD5ACHNuzgXkLwbzR3s20EvkTlDVy/iE4ffBN/BiPjOHJtFqK3HKcbaN
CIMbCIBbfXsbW3JTKV+/7GS+MHmI9rqfqpL0WaCzJk4atUWFP1NekqPqkRt4HJrk
Epb62JBsmc0oxE2LpVd5D38wTPRw1602X3Z0TKfZ6igka9SWdoeQYa1Xu2p6zpiQ
/EId2DUFDuz/zWmqxVmBXtPLD4lylovPUvsFn/iuirGHKDRhbGPLCWBMC4DSPYKb
sTebIZfljyapEcbR+Pm5ixelaqF6jxFMnuBhECDWW41HMwoGoc1Ar1TM/XU7sWOb
warA0IVOemyQOdPcUwX3Eu9ak+wOJFIwSWuUz6lD2ZThecK1TU6iEJvP+WRX2S8A
QtvT/AFHi/OHA6UTI9QsymYQnpTy2lAeAMmnRlrStkuevrgV54rDuq2nT+twJ0yy
S6m+4W5Vc3KtF20Z7+FQgio7r+lIIK9J5TngPM4faya1btc4vRsmgyAUm6enPP1j
ANphy4oJ4FILvzJEpNjnAYLtE+qrtzuTPZPZWrsu4CmMEYXzpBjfiNCOoDIkjJy4
qBYGHtP6s/mJpPce6wXVe9HdlFG3jzBhMAu6+1E+RiOvEREJl6jWkDqv0Ak86+N6
+zFv9KTkVGzyN76izLXBjix+GZjT1EWBSS3SdVXfEsDZTa5WcFbT3hUJhCSXj99O
v2BU+XEi1A8GVRQRPpzVP0Ak9Ofa3a/GjcEVX1OxKF/GgxH+hsn0Cs16EjSooodY
aGm2LDfqZiLtpLFFjy+RPaunbHtbicX1aQEo9c8QpcPZqk/bIOYFKbTezzrZOiUB
YIkW2YJcJWsL8zECE5xJGB6axDpzD2R+tJ7nApGHcNK8FQ1W+H8DF+KDMdHSe+y7
nkVApZyu1vKF6EJAufi0rdfBPu7LBjkx3VLgjDwi/qlpWar/csJMju6nbim3PyEF
K16g1toNIPQF+C1GSa8oMvxpQKiF11MyduIw29YSv0A4l016bbrzTTKUbmON1kkf
eZYzagYNcaEM1ZwF5cyAj42U/3tlJYtFd03nO0I6YCkSQtWO0AFAaNK41jqOuroz
DtcG+Vt1bkCA8FV/HW4Y/dlkyFOjNxQlBFiBEonkpkv8Uy5GZzK3PZBFFcWykVUd
t+R4wWq9CiigQt+gd8yFHsbxIisqy+bKsw7/y6w+n4UXLBj4OC7mwv/SUKWHC6S3
7H2dp9L4kSenXdafDsJVGyygCqPP66ZqJpqDfn/yt6Oq36pGndOKzsKmcE2QyWBE
K1bX6V1d/gzq5JalLQf6f7q8K3N+fMlW/nHRM3ckSEinCsrJlQQ1mWhz12Cjr8wK
WUeJONx0n0xaHP4oIkzs2wmcAImdN5skn/X99w/TFtbzACAuVBUpf1eocJvPLrv+
FVMP+AdaFMA0h4nmJpvF9MA3Gna4NDHC/lAowpma0vX7lbC9kIs+7qF2O6pSQmeX
mOoZe0Uan6wb5YcJi2915A19ebJxx9whCj8e3f//gbNTeR/DTYgXpzG18vfJQ9Ni
83vN0qJbMSOeavRD8Xf09Mg8UVH6wtuEdbiVpNGwOwS68DI0p5HY+zW8uYAA13gH
uBlb8bD5rYAOLR7nNj3n4d9TGjeye4xc36HfYYLSmHFPBl5K81WDQAG4P7fPWv+N
wc7aLX+RCP7Ry0Lr9+Uu9DEX2bdmY1emUr8dVFkQv3soDw+mGHhPOOQlp27W1pxx
i1nA0qpv0nSOrrJ9YCgnXmmMDJ+KOlCOJYb+XhQR8lMmdPoAIPn4nqlFRp559ETC
so8m16VL7EBYDkzzp3raEex/GwqznrNl5fFWpH3kZ2+tQ8wv2kqhVcj+alhC1Dzn
SIaiETs257EiPK8xUJLZ25aQrkmVP6gZanM29MRPVqRx8RPMZeLdIFFjvf1J/hl6
JeIOI5T4eJkrr8OUw7QuXsx3KIPigexje9IDAhX0BKwaHfxTx+iJVfXuhLvwpAgD
oo+ShpeVTdK/NV9Jo70THmYu5w26c1GTZb9pt6cxvDWMhkFeE+AO5OFaumwBBsHI
Fgtq6/Q/us8bcRZLHppzlWrFl6Rpf24GtXaeH8VKG5EunoUqaUjMpdKu/YRa3QYk
LkqlR/NUP2wZEq7Zv9CpKTDPgld9y8/Bmz/cKhWd+wVm90IYgrVohq0PWAYpDaTV
n2zUzjcQS5h6Nuf/XhvuGujYSYju8RJ4gcxYAH/UVeBD2EGwDNARuVD/nELHzSnI
ijaD7EdHrtE9xahJwAJySY0FjGvuqwa89YtmgHQMyl17xbdFAIjRAUvpnPnNyZXx
XZCy2x0EZ4dNT7BNRTMjPUCPxms5u0POLfmXT8fqmp+YYMDNepoMybg0qxyd6Gl+
Skyh7awkYiBO+dy/osJhVhKpiTHBo2OPQZRcUnT7QtEUAqAdNTLfFKefUlyGEOtQ
9zF0I46Ps9FcY7c/f+f+1AostKzPOKprinhaBxV1CyxP7bOV6O4uxIdc4XFK6Raw
5+Xd+MYQKmyoR7QLEGCS3r3gY8UOmv8UX8wGQ8aOZnQ1ZnY4tjv7+GqIMeKOq8XB
CXQbMDR0ZCtOxL12rvuL280J2LStQJ6TItWNYxuLeKX4lIeOliME7lz/kd1uOuLY
Hm/mZbiM8XZb9idV7mU+1wsjUAhv141Y8MTSnNSmZEuDY/U0caxsUa9w+Vn0ANYv
+BOgpN8kwGNY/M6ZPr80acEuVimMGDM1DinbDk0XRgegfMumK2mBBwSZAawZIyNf
uH0zqP4A22pthCIHd5n6UygaUCQaRaN1wdJAG8sDoe5tZr8GmNPozqXjygVP+vZv
8XcH950T89qoczPVZbzqDyrGPS487UvAHsryq5SH44jOAMJmxhIZEAkRSKRa/b0T
TQNBhEDPXgzk3aYkKA2XqPAP1xUhHczwUjs12+rso4WPDo1H3s4Us1Md4turKzoI
Rp433LsnGVHy1kSREvj679X6CI9ZXV5W8r/sNWK7HiEMAX2FW6y7RX0qIs5qVlnd
k02qYbOEG/nZyxPxxa2MXOI+Hw0YeFmMRXG4DCGsOEFMZDQ4LmwanEXDkgbTmXDl
EB0++74Sz6b9QfIzzUPLEV0kFN3CWh0FHtgSdkXPR/dbYHwD30KwJkwEzjh5Xmzh
JlkYvBmvl4LlsBtSQSiJlggHh06W9hjoyazLAt5g7G8yD5dz++IChprwWh/F6x4z
r7OMQWtwck/ZTjwxz8S/BR1rSSiD9PR+xRy6Rt4BI8waoj+cK6kqgaaDMDOMtLn6
mctBD9AEwItWwNU7Q3lGil+1NpN6MUZQI1pKP1xRb07/HpLlGGB7tqJ6XFh/U5EV
V4BeGiJ9W9MOMuYwfuivQ89ZTdI82z3ggu2YrjOSTovoiOPqr9+pcPGyKcdj9R17
gqusvSVDEc6UngQpAciYoVa/58k8zltGprDzgXn9EqP8ZZ3wJdotSeOZUQT9RBXx
eu5lTnXJV+ogt1GQqEkZN8wpPwEX6GY4DT42Tehd/4NKFMcw/8Mb8MwHOn8veOZ3
IB3mbiW4l93eOnFZlvHMvBYXkpVjFCWjBf/FYJZwAlOGB3f4Nnt/GLiZGoaN1sLV
cem63oszomvoPV6cCenOU00Z6jjcjuNAq5JRP/gyMZNYQ+qP82ZX0132c74h4/Yj
uQZJIZ3PXAUsH36K1Q67itsQC9TJT8m9WCsO/70RyAkvmqn1YKtEXdMjrQPvlhb/
jsl0mxlnZHBSGAF9yvDopdaFeELKcc/xhELyFLZOa3rJMXOVl1i0C3xIB8k4AJfJ
Z7xAZBL/VlrQOMZZs9hTqlvty8++nFxT8Pp0+I8sOZEJvXunHF5IibcG0Oolpx9z
vnWOdEurtna4MBsuKE4OHG53lm8cRwmv/X2nJB24OApb4E/KKQ69p76vhPy8kSG5
+ygyMOef+TlDzFd/hB+n4Xs5JoF0XSOH1In9XKPeBCpSV6Edh5cPlY+NI/rbrAvK
OiLe9n8zttdx2gqcYJ8oAK20s3WZrrsBrw86sV7Yb6ff1DlC1AmrtAFdbVGgVJFD
VhQMRkInlAkwxlNndxtRo9NgbMl8Xo2lSwMzMKV658PGSq7v6HPAXIsgzkMOGvJx
h8D2zsNBNiD7gRBJbFW+3Q9S8XMg4rQ+7t5hrOdzYpq5iKPcQv4gpMpYk6V+o5s1
mv6JKF6UfFQnXwsfh+Yi4jLrv6kRIzF4erL3KhyEaItJbnxTTBvMNhF0syB2cZF/
gNlhMJLOvCqsfLaG9cUPUy3J23qruAE3gKpGYwDk7g7HzOdm0IORNhu+uHZXKu6O
r1bEer4NPg6jATw6gLjHCSVMhZkmES/yC/dHbXknhL109F6hsG5673FEchb8AmyF
HmqohZ9RfdrD9F9DqROCnCI0qRaX/KziUjCZy0jebdC/ZFhgJeN8CYkUh3Fnf0+m
6vBgZLTUnUD3TFkUBP/xSERZ/nGYDvnIRNcToYfsNBDak5wnE81gBMRqRus/kF97
Bmxe5HGLR3Jsirn3g/775L1fWpqWGotcJN/sQ2FVQrjgoCzj6b+svA0v0rpVe6On
kYNQS3v7W6beuMDDi42gci5t04IJNVWUVP9TDkStw9umr6/x2EexOBQKs5YQeLVm
fyvhIzy4p/3nOl7QQVZtU5yqxhEjau5AGz3d7GLMU67+jOmfsnZauaGaoOKKMUza
cbIxHzAbkPHwtPIC7YysXYq9CYZcQzmKwcMulEvV0vVgzCtu7PmfaCBX69vT4fJM
Ue2j9wTnGmQOUjX92Rhdg8w2rjs5mJiaL0xWhzWYYBj9MtSmMZHEg1+3iwWX3q7G
1jBy/aLA4vls+mmBMY324hIo4nxOhJpxo7DhZVafrGYEMDWoY/z1XnmYVLlIqmL+
iU5noSpJ9NaM+8GzXnU7jOW3OGyIb/9CLO/zYcPLx4EXybfy7XdkhvlLelHzOZiH
tRbw5a9Vzpc21TxY+va5POT1A0dowme9DguxY1OUuWiPmrGJ7uH+WzVJiSJFBz6G
JVo8Q+8WIr0cZ9rh+fLxanITYpijTeCQE60OxMi5qPRNWXQm+Mm2ddDOSbFnoOP0
duhN8dc22OWxFwq+dMwpDiicTspBtyk85S+9SWeggdw6MF4KZ3HAd6dzvID9KRRs
52nQ5F2F7IAZvgi5P+UGF3tNaHPtaxbP8l8TZARyMdowSa0CnqCSiafR01zM5+sx
ba9Bw1auFYZ/SoZnXYO7qUWI0IHcGANU61dQFKYehddTa6efN8xoKSVr0zYujBDy
ykUzrrgp8x1t/Sw1gGKeh7F+0anv68KNc752rjSycUbyAvtmrgbaTHBTiNJCSAkS
/LCzFPl2RUxtwVw/w284+hbTKUQWwFs6E/rnsa/aUO9Xs3IUURH+Pw+qMpQWwogi
MhKnEaPyj+eTyEs2OwMkZ5Yu7qacHkJYPoKKxkzNmsIwije1sJ9aGMDgS85imkwe
gNdxkzr3rax6BIMwSkhHC5cE0hoP+iBtjDjBX1d92mvM9tz5jjMYdj45XQ1eD6Kv
zL+uMBGep1j2iDlxuoUq90BTl09YnOGQOle7lFXFCFJr5vxHIEevA44/r7Uasqh4
N2ZuzqOsZRTkqO7YTh7rOMC66NfQVzqwsORUmL6KcLMfhf2lj0mND3ASmY9fx5YQ
d2Io0XYkcdVqGKEE2hFobN0SsafArPqLsSt5+Mh1L4Ag4EIVm8WKotwpU1oGJUeP
lMtWENA4z/5b61B6GLkrr0ujHSXHrrJ7GECM449g0f3CQKgrmm474dkpfmybzW3R
gxTNJaVCSMKrlCtGZFZpH2reLxG9q5tRmedmdSrr7xMeVSEpH/6jiTyRwLlHRxee
TCxuYbgKm9z1qieoRmEw4yy2daPZkrJHN0HEpvM8yPpmbGisbT51LfaK0o5akY/e
UDDtyYPxpZtL3Bd/e4a1Viu46Ce2lNZaXNHgu4K8JXY8wSLhRPuZXRS+rpIb6iR4
PcoVTo66VY9a9GeRiANFwZE7fOn1TTimqrkWPTrJU9ZL1ZpaniNIPbQs3pNNZkEC
KU/jKljsGpNcz9XnsDUU7+AIIlc25FCyD614FOe0rGS5BNKTDb4XC4zTo/vr28hv
2H16k/gcm5KYc1qW6kjllC5UydocoDOk+ZNK23T1weZj4eO6uFPqHhATr/tTPrkX
PHgzGfTtogsut2elDDFo4tgRaQxCl27zYdGJc/PCFG+SKMcwFIBDGaFROBOU1YBe
BmG/ThzfwCXxrIxOKPCc4XyGCvdbQzGZSmKWvq5koYTE9bPUgeZpA9/hh8Tejzx9
ol5JdbOlwTqxA+Gw/14ra59pkaEszRnYFVFcQn9DgHTZdtmeTMVk9wzenizYREGe
E1Svdm+uLuMGBfLb+TcqHZii8OXv8RoNdZRpum15ffj0X/oNUowkdOobcpfGeqwR
9awgThxO6CzbMx8gJLrB2AvOS8uuD2CoDOiIdptkUDnYEFKbYn8xTOKIo+mGgT4e
Joj/o0PRKJoityy8PqRAzB5nGlTcAh06EaygHqwkl9pfkr4UjYvuX3no2qklr59R
7w4QC/faAs7VyQ7A7IvO9qfYyPCLpqGOX4HF2zi9VtkG0LsqPBGUAczBjMfLNm9q
/TpVd/2SG20PZtfUaBlSMYN1QTTn7h2MlMIcjknV8ORdXoJayShCAa9JGnyGWXu1
edcjN89s7LYuByCXeQrsoRIC3fX8bTraN8QMq+mxiSLxfrVlgqVJfu2gvfp2DC6U
tOUX82WMxMdZl8V1HCy6TAOFGQTXtWi8XAp9SOwwMI4hwtpcKTh/U64xMMc+Gud9
v5sUmG8HpLyaiI/pN+hHrfQ18ihYcTIf/W3gw7/VKYUE9gdqUvQdCJzxF7sV5sKb
S36NDrd+ws/YJ9kV5Xokk6DLoE58Fnsn9zDeCBwNNT1Th0AOvnxZQ8bhP8I7dMao
E8+Rb9EOtwEHBqI8bjx+NgxLpQQJ47yXhYFCTIlB+IzEi+qSYu7k4obeEM7n+1rX
dYNwZhjm/LsPcOKcc68i3J4g8EEwm4PSIxSzvSBY1uKynYAcYPTqUEeIrbMqsBXC
jXBV+Q1WpdMfa/J2Bm9rVvBRSlcMpHYuC6YYROUuiXeCP2fjUT1MUPAhYPwETp/g
gz7Scf90p6IMZ5zxRkn6whblntnAULtQ1rbKi1b7dEKPwxmzymjICOJ448gUeD5U
m9Lkp2WBAVX6hqWBdxBe42RNw+RPR+01aMuTI+YXqlCvnF4Hpi75vshGr2DcsxxL
zTsMDhqYIP7W22hAQVLyrD8BMMoUvkDtbyR5hkgoBVY+mpq1EtvHl77IUYx7pm2o
Hx2Ltnl/8NpL10VA3xYHn2ZSWyzGYnceA6lWzFa7G+QGsaRBoiyrDbQFSTgbsII+
u2I6WWwkQkbDsACz0PVeNN2/53iMrpg5SxvqMl1fUYwkKQlurRiYRcu2bJ+8qF6v
MwDPyUUoENLd7iXQ/nRe9O77ehJVSpfyLqFdWxtF5bSUgyQ+wDrVZ0mV6QWFWimO
FUCt30tImtQXrP8vKfX6w1WVvQrhNic25wuxwPVtoCxFSr/48wHh9WQjuQHQcaXZ
jHXORKsiLwNZvgkWf9c6pVEgrl+k9RmndvRlgsZ+TMWxRR03a9PWM4RA/8fHVJJ1
x0aoQ780hJm4bKd0eci6cWnSRiqyiDu4ykFecXsHgiclor4rZwQ8MKbPkCutSVUw
fu+aWtW1+atWjqDedFPk3WsoQ6tq6BdNcF4DQcGeceITkz9dgVPvmXKCXLp/Wk4R
CGof9OJFAi5YY0HYnWh2HWyA36v+mbvXANRPzCIFaBfJJw5oZ0P0EjIPnE5usyz5
cUuio8qhX6lnFnW1oHXPD8X1DzsKnz87uEVD6K7b7qarVDcdvW5ueRfk8NJ61S2T
zjKBYtDn1If5SfpX1+l0qOCa8RBRKKmgERQp/GTV73dxlW85R//cEo2ri/eFqJnE
XqwFGoaXGPMumVJfeNCTxC8+r60a8dN81jplfuiF+6XxJ8Jy7kjdCnfV7b8Cifm5
JEznHQ4x30BKRzSSQKdFYgoSQ2xIxYESDRDDwZ4scBoPWP60aBbegImI5GSvu4j7
/VeYQxBYOUNi/1XOH2RtQVUBIA9DmHPa65R5/CstfIThbTqkV3OGtpd1mw2q1JKs
0+wePjSRvFCw+Q9tGaY3sq7T1LbUm26A/QGYYoQ2az1pPTWtLXJNaGdjBNa5IAD/
z0VfKvx1YKKmHsMDvnZO9dbrpyF12m2vdNyWoQF8Xwkkxfwpcamfr8NIuI//Qo/g
EgnYkh2D/e0hGPsKiH9vZyvBO6z6LoVIxTqna2ETrpY40pFU8JRnsmXQ/MemeXeE
i7meVSMHWyZFQOTjOLXtu8UqEQZ3Oz6+hWrzebY49qLNlLLQ7Haw2ug8zmKeoncy
x9QmeHxhAh+feyQWj9PuvMt+SqGQ+WxadxNjoYpDduP5pPYZqonbj7CrXRaVCSd+
ty6+I7tQNAZX8aygEgi9Db3mfoe1S9EwkKhpzVJ9pEK8E9XWJH58ZeBfG8fTI3PS
0XLs4lWuSp+ywHLrL3V1zXf18nWC7Sn6lFa/WPq7wWtYeV8HJQ8pWRS57aLs0Bok
M7gKyGhkBzKh0u2ri+CCl4OBSaBUhS4KWN0FdGb5m4aAMwfo79pzugS93yDPoAQM
pxGIZZ10y3nUMvlVgPJbXuQznyUgxfG9dTBo9+JZznuABmbRmgvlaPZ+ZvdEWX+I
UuUqRQDIidI1JIAz7Nt8Vkf7vzn4EvhwzOlQxdUUUmwMlbzrC598es+Q7ACuWRZ3
MmIjcyz/6OEDSvEDJPonLJXczSd7+4/3f4IkttWI2CmArWezuV8sWqUQr4xSBz0E
kJdVmvhSnqnMTccdfR6phFTc2AX+ss5/OFxygCkio4da+hNliqJDB0q1RNsm5Gra
L7ODOJSvYIS1GBXEfsJOcnTdjQIysUWMzr5oq5+RXlvR0s6tHaDH3AjgKjYigjNK
BvJsCOaNihDfcjVv+XEG8n6Mc4Pb1yP2KsF+QRri1c3zdWgOeZyOUyDwgkcwuw/3
HJkhxQQQex1kbqQ9nDgTenX1rxYRniBHsHxYaFmPr1jedaa9hyn99Qn7TuAmTe4+
n0JEq6lHK7ItX6yeM2LX9pxXWWbjTrt4BfRrqVNDQxTrv/atLkvC8rTtEaN27On5
KCbzMbiBVhoEmO0qYxMpD+PfpEpABuCIWrzWngZu37ulcVYgbEiYUvTysdmSG5Rm
C2sf94q9lxkkLQJl1hrh//kmJZeGckigetnUjXPrvJgTUhRi2ULmd/h2hF7rHyG2
OT0W58/TlnwWXhL/WAdu51W2IIdQP7dm7U2IPIZ2Aaq5f8bSioOg498IGbgy0Goi
kV+joIdr2oPrQIiCv3cO75q+9KZvyOCqFJaR5i3/fVWBvWPEeiFldcKgEA23PLhn
J2YDD8e2JfBQo2Nqanw3yk3I9MSaUhyr2HKobPLm/4FK6FIdyORnnzedGdqu1EnA
oln6Tx0FV4Tcj8JCESKBXyNdzK9xAY9mfWxlQVlT0GOXGrC96WyN0WgrVsb6N3zp
jRgJMHfp+ATRB1TiEh7EK6ucmO2X/lBNfrqTNgNvF+ndEPJJpO10RFRXkjZpm52M
+6YAevjNZNBvnX1Dalhw1seJjWV9kpow0UpCKjXUgyOovUAdkJ30nbKsc47fAvkp
skYqpBrNKbW1G26O9lIlohdTB+ACtNAjcH+HPUmuDmNX/H6DIB6dF1WRYbP2j1n1
83y5jxzPBO7rW95GcU28EDb/aPs+TV2ZKl/canNa1PE/weWmLzvbrbxXi+1WR9hl
hDP/tMwU1TdHNWvtturUKgtfRodbINtPNAd6IeiEyMN5yEz1/LB/KpINzatnyGwS
J5dCDnxjNTKr9dxcAWYUkWQCGIyhaxJniBpEpsLk3eKoZjN5vQlYFzydaQJPprFS
nqGu3FWxUD4J40XeeQGzcmX1wqObxtoUDwX1XbrjEtcNT57+/qi0nO9+S745MwzR
N6uG1U7d/8uqkbY7QGrEL6SH3fYI4fHUhYUhiIaIPdw+edWHsYUizc5Kgx6/cPjX
qi2S4VQlPN/9PyqBHcZmmTZnqnPcYmxkows3m6JthHV8gki/Fb0co4OuKn2HzD0g
jZgsjBCvXk3i1HGJYYx7feMVvgxPfJntGCSYpjwdfhKqruzEGrA4qBckURgWaYuZ
z8AvnMR5FcP4Myxa3dJDsHQjUcl768Si27uvx9Twz7oAXjkLuR+1CMQ2tQqQbpsL
tDUBtERJvuPZVUQM6VEodcPL4RaV1hMyOprqMjuqegIeHdHZnGL7tggw9wIvGt/g
IHbgRxLZ2mbvFH8CgKVg9kozu1gBSNwKHZBU+a+GXkGSsTu7bATUPx2GYDeESnYg
hDisGZN+B4Hqid3cKORuYZ/07cZMOtE/jMXjffPN8IlAeeRPhF480SBwJc7wrs7C
kmXZyOiycrUU3t5CVNnVanR7N/R7Aq+LY/z0BZR0mhwDMJGpRatJQLZu4c1SSx+Y
FrAG4G0iwEJgQQ2qu1BhVQCWHtbcAmE9AvsxVAEIA7C8OSaKJAktu0fZgtObWOwj
x5Jkd9AuM9HmVzNXl7FseoqmnemJMfC6osqlwIhyupnBY6kLqIxwh/hpqUYQbEQk
rC5FN7gy0lRgIOB/Ooxx6Dgovo5zF9+eEmD4hv107s5LOhiOySKE2nnZwpnCa04y
jEsZ27cD7xLkd06YmynvPyCpeEFEq7ngZUjq+GX4/D/2A+Mys2JqSjWuQ7MOuYJd
UH8JM0RxixnRu00RqkIavV7HUGW9SHL7geaHKO0eY15yKp2cCFmn9U2l+O+sO62X
lr7gAAf0BH7WtCcAUo1M5S+63xEpFUb37hgmLSs2tRhItck0YCKHZ9JoZcAKlrmN
WNraPSLV9YKQ1P6LGA6U0O6MlPbHsluC8iarhdWV7RxWLVRJQnTyV6IDaZVColJs
I2Ti9OKhqdfHzFdCprM5jHz1kh/n2ohnW4K3seUbZg+O52PxpQ2ekyv+/wTSQf3g
xtfeXZU4oibshWEOvj4uvv9clc4KLpcNLF9xjcoKLilYLpWKOz9mzEupRxoTAwF7
bkj78MWGOpT+1Cg5rO9v04hCShKvvZC/bl6TwQB2c1gaNIgHJQ2EXMDP64jq6NjP
n2BASW/k3vE8GbYpCovWs1D/OZhw2B/zaRoBpwNk5uqxHajG3YTs+Sj9qo6J8jvp
UEBXtTDLzq3OhZdCrKROJZdtznYo2sDtMRwbahspSPiHY3RH5jslWEBc7GjIYplL
VrEem5ax7dIwuoLTILcAXuO7Fid/hjlnLvecnSYC1AJx5eziWb58UpyQWw3ntDtF
AVAdynkB237+MALC7iiPfv1H5vxaNRZee5egecDHeu9qvODu2JGsuQto1bTVzY1L
ReDCRwIzGvUp2FSfmynZgK4RReWoALxZOnB2kw0wdpd6qahU8D1uJDaoiuGvH/r5
1kqnoPeZKUBjZHtvBeFnaMSlbho86pe6DgHQgrmMrxJtIL+XSOJ6ZHU1qZGX0634
/3C5DXrAKnvDY3UFjmxYZRcDG8iKY5pqm2elc14AmEk/7SQZGZbRsjtXpFDZARXA
Br4u6KaKNm4QtiCL0PlCPfh6INt9zsjgbR4uIUgDhlrUyH4v5wlCVPI+UJXFgjnQ
xbn+s24uEv9DwSY50ViaUzbud2zlXOgNn7YDbeLnSUkUy4HYvikl96mU2JusTVre
Y/nEgvkNiMDg97TNw6chrZOT/SKU3ydc+pwmSW5lkNMXkHXPQU4U2s9psN8fn3FH
CAeq5RolU96R/6q40gG6wUzwH+4csv3EpPIly2Nt8v3eEs2NRiRawnFBpSBnSDQt
b4QIs3K5PthC/eDV9q0ZCa/Ile42wNHYNTELv4pRkpWLWn2J0eLOdFlhWmOFom7M
vnQTapRybJz4cT5FjY/+TsN113PYoYnYDboie+ZGC5arEQCH3LlaVZKGGtw9pzwh
Yjp2nviGIP7n0XHr22EAgFKpUw7nZXh1gULjBvG7s1ifGesI9wtV9VGf0o9dtfoW
uicJTvJC2j+KSfF6Lqef9knIqnbCI7kL8/et+3+/V5qZEieQ1/8bFPHsWnu+XavZ
OtzziH8pTAlp+o3pOQtlIZ4WrANO7xgDlQoR/5UZ+OQFV/XawT1M97mb9DrCYF/6
HYp1ZnDyLULDjlfZTNeq31QeTEZ7BhOJDLWxztv9kTynvMw/anPJ6dkh/Ca4VihQ
4b1SwkJqGkGG0ajXaL1CuMfl9Fa7YqOBQBC8hAoAexMVmWaW2ZqIwZGwkqFrt42Y
seHpCtzGKJSwuMS4Dgu/GrOIVUMIkLN4S3W2ApBx7Tcf6RPK4JYv9GBU9StdqCWb
i/Mx9gUxHlequvbqw5jzDbzCUu4VnzFNilBbBWJvIzEvWmJUokJBJXA2HMfAtfmw
kTx0+lN3aYYGgz1q7TZZGcPA53DoM/imnPHk0bvNnh268isb1Wn/5q2dtPevkRiF
K1NBxhTB8Jwn8wq0Fp4Z4DsNjIVfCzOQxa8aGBOP9hEQ5D2uvwczHTqSYgwtg5hu
YZQWsYlVnRW2EDhYlgOqerJzSmJVNg4Xelzocl74YX7lvM9Rj1mKaXHL+q7G9H4f
8q+1lwXkeSUs86x5zHGDZyoO3AmAR5tPMh2Z5MAQwr9pG7ygy8M0E8tOpq1o9GWU
HzONn1Y6oZPa1Vdc8GPMx+OrQ7RvRuZ8mu7IKZmGMRLlvbFc7OwISslNbgxNIgIr
XzwHxHR3TjzR7WZnG9epBAQgAjk4Ji2ey8mKyoAbAGr/hi0uDKoensXMzUuyPXcj
jR/bSvxlvsq3JVGquGHp3kAqJcausoSWac0CFz4hDX/yB7Ysl2lI0eoETCPat4RU
oVFQ6zrKQ0KgqaixTmSHx5C3JPcXlw/AnCk7/kWQPf5PA8hiSeOp2vlCq5/pSBMm
S6it6cxT+2Zmesg7qBr1U31+i0AyjAAS5ssQ/vNv2ttEaJLDIkH+/zmjiYODKadE
30taS2ncL70ZykkAtQW8ih0PEwin4fC/VNwcFi4y/mFKin7czxVnIxUL65nfUnCS
OvL9oT71QNPx6f/iFnI1kIxMlIKvskBdO3dVg67ryB8huOtVXK3+i7X94IY5oMSK
5kSJfHoUwq+Y+3W5ojQDhCyR8MY1JdoBbjPr6WGpDVwe90K7qSSjiV1xZFi6c9EI
Fg69P35oOMpdBIczlis+yvxjtmHw/0rQHuE7JA21LDcliSu2jP06cpHlRa1Ez6Ec
iowKgzwolGJ9ootDaLpq0sRZeHWB0Vxv86y2oaqoy9u1hduUwmhIei7VMWD5AAyq
ls3eW4pUlZxsApIeS/ZGhk5gqV8vSC5IArzqaa4Spu+Rew51shILmJ2cqseb+DN1
0IDbKHk/5RFbgCKRcfpx1grN46RpFub4TWDsxPXiephgHqAt9Zpxn2h3/6Cs6zy6
3Aevr5uEOC4gzEy7avKjQFBFcYvYAEgp8ywEhBSnS1X4FPUnqqX5u6OdCr0y/wRu
opFye6lwaWz5siSs+3aQKb0YIeRx72x00xd3mnW+oh+MizaV7EBq+U1W/tGzAswN
LgyybOIO7nPv17ey/SBneQJj85zwfW70vU3TkN/H6C+Ro+vKn8bVQz5q6nio9HD0
uKqwUrSCZ6x8XyK1lTyMR1gzZlFPsIYEvQ1mmm4QUvodqxOoYkyZ6syNH//2nAzC
CUR2Lm37ZlYmcaSqnSZ2C0J3yX1KckbyDgQVpABavyenrlg0Fz+B/mlui0vMNYNp
q4CR+X5Od08/ZXmVK85x53+V+tFsXqL9DyG3Z+u/8bzyVGICwB0nR9pxvIr3TqVG
o5VhpcMjKoNJiuEwlkT12eW1XSC7M13n+f0tdZDdx8tJNtxe9cXgdtA3ZfSgza6F
rH20iVVvzfZIpLdBE37WD570bs4awLV4o9pztcfNAtMFthLTNErezdWrLRROztuL
6rS17rsLH62kk0XNalrTe2D+R/vK+FSVBCf6d0jQPLmUXzxNwduePfCvNGwepngY
ne5VAUpVEaf/lHBJB/CtjSFxL0Cgm0P2ilGL6hu6Xz81uQ1+yS7PY9SkIJxVELmD
DhkLWQ5iXfxe+Q35G6DsH1GkszOCRCooCcOs/kuT4HdUbj/ZqL/W6ev1+mC3XYDu
hD/i6DlZrPiZPhQ3Q7cnDISnsu2nJG3VU59SI7hTzbZPKoKSH3xuSrvO6fJhi0aa
xT9XMN3s+6v6ykBcHX+A5WVB+6KIlcufz/4ZJAGYod3/38kcybOMnvY062/m50/b
3MTcyruxVcHn3ku25SbmXmbmoXSKHgQAOBx5ixZaw6lGW0j5NENqRdW28tS1aX6J
9diE/5+n7mU2MA2qpyqZamqRvTu+WYeN/vdOrFu/YStWsXq2uGAa1jOqYBm1BM1I
4s8o+Wpw+z7coG+IOb8W4Q/i0gHTZkk0YK7pFJGWTDA8gCuifFfvTh5DUOUjbGYo
GLvDcpOweyt2D1Od8dq95W02TEyJN4Jg4nzVjrr6eS4gw7y9+I4n2vHnBILrmUha
T37lFC2YAobTTsvwh6NWlt1fqkpNAMhr0VOEIQEi+EacjSI2oUQBpAlhe7xaLych
3CoDNrzD3GDK0QXQMTcbDP4xaPwz/0AGOMOJnhk8iI9vlc9byn+AZVlUTEXWeENz
hqzvSDpQp9U9PjQT77UlgbnTiFnbeYeWkNl7O44xG5jqozwbmt/WPIRwOycIBfQG
72nOA9twJ25v5r/cXEjWc9tqzMrbUrZA4rCLyo3VVFTidnASOnNP6uZFo5NrKdSR
BaCnw44zIt6rXShxfWrKon+yOwzmvKu9U0Su2ZxVocoz+RrehIZbgy3U5NvTcdQx
xCu3IEOHwdUhULt26haBCzL8saGZoEdpjjWv4BuiDZ7zObxQYiSGscIrC4B8bXSn
TIEY9ltqNnHoKg43kI/wyqDaKb89S021SNX7r8iFjEGu6Vbag9HnGvaNKEb5lWa4
/jGUUgmiG+D9FLnxV9eP+4b705ogM2UDaoKnsPXHhoGyApsDLmui0p8TQTKl/Bgn
RPp3bp1WzlCulIkEf+QH2nLsaMansXYLPzfCzXcZOlubZteA/7Sj6w/i7mbmEqMc
uJr0+tOLCYoGh8j+Z1byrPtEHL50R5164M/LPrP7nswHghKeKb/CW39la6Cd9edP
Z6ULD5aMdLvZKTN+NnEuNO+XtPsTNbTQrR662wTeugIyhIWt7CksSA7G5Z8QdYmJ
yhzCJljOQiNfcM1hdpLxHEi+iVQVC27RXGdIxaHY2Wfsu2/qkX283IkrsfwUQB/z
ssILdq4TB0ipJrRHF7kv4myZhUkUx+gc8WYOEw9CuRlCH0AhDWYnH/UnWm9LBnkl
m2EHwpFiVxMdye+1k8ERYCpNhj5nlBvekhd+5cbmHa+gm6vaNiNdaxPq/NPxPoOv
ulbSxYfJozQw7lQnVXAbSVFje6sSgGFLhrD8x/V2xZCx3Miqa1PX59bnNa7AFMO6
Nj/pKUfwPZZak/s1uVH5lQIs0//5YYYoBaNi/OfUmRnBS9aREmuGz4ebKzZ4tyB1
Pv/mXCi8zDa8SHP3Xq/DjvJqKInXPHX1X4Eb9doek8eC2Dm7waJdep0SWOmRKtRJ
w0MhMIwvh2S36CrZuP0bmH/8yYIkrsq4bGJ3YI+NcW3E1G/bTaCNaBFTnMEndW+2
rHi8CCF/I/GI58TmMLB4ThyDKT0owoAHuNbSzJcr/sWcc+KqASMR5/GLGNhq/YzD
flQb9hMxCSYW9e0ot0q+QqLczGljtekn5cp0OYeEaB7oxfK0ZGhF6+qSQz3MYksb
Kdlmthrhsj16E8NzgyTh/9tcqcA1ruq5Wa9efP7vGAsorSINJ45LCcSfehr/iydP
FCqC7lZwP5jktSLUiuwIecggj4fxB5qi3F7KQ2OhfnliX5m1NbcUtShx9cP0hgY4
yDg+hvcbKYCrbfwrmuEtixJRaOCH0Ae+OKw4EjgmcKnwJIYjRWr3lGatwptJOh0r
FVv4uo3GpSoqVxhTvtXwD65a0TLPOOZETAK3n/OrGawvQezo4kU1gWY1aTOP1gXD
UsQpyjH5wPoAc3w56RChdNkL6iD9eQJ11aH6Q9W7ZcLgGpwchFNOt6cHd7XGdrCD
jSNV6zKs99+bJISXIE/sS7VdNJKHVszWJMbvJ2lo3/N4VzSmfwEkh5JZYMSKyGq4
FG5pep5oW4D/DYbuiumGG1YnIHpgwPZt6ISFJVj7dxPFslEiGim4RAFGuhl8tL2y
xV6fwVK/thm46U0Nm/6ffvMrj8RHlYJn/0FD5dNiHCHs4E0dH1QTbmCYvXxhfZVm
avbsaylsSbVQcQApFPT8qnYCMTqTyopDi3ar7Sq4sdKCl5eVZcLCEklVmjBXfmMY
D0KvPKmG6/p6fqkMmAtEVaMMGb9vZ/IvTZfMYsry9jZslLvUPy2Nm9w3QxETKc3y
Rhu0uo7Wu8BxEU5pTIMBbpsC7G4W34tKNxpCMe8EcJ4KMN9BSqIvVLO0crX621iK
2wBPDQM3eUQoqD2V1wlAu4jWQeDkE1dH838dJLB/uu0ZtGxcEoABI57wGs3fUywt
aChUowG8wY0rj6LJFKIr/U0sjBZegpEeERKNW9ynfSD5KsgpomBwB1XKvE7B2bvt
DHO4crCi41d3TfKSLD/lltPFwynMQVRIy7rgbrs9KMuAebbR2GjWUv5DouepcKHb
/5EX8BtUAImQ83YD5axUTeHyM50jvldLrLiaGStLcLLv3Okzl0Kpxe8nbQe/2DT3
aZtipmdedg4UINz68J6Y57uK6AQKRfEtAPEj6+TOCNhLBjzVLmBkUOubzqmy2CAr
odBi13KT5C/3L+ZeZOcub44u5PJvVLHZdsaxZnoe7Us+vGV4xe2AVWnX6n5GP98D
TuNGdS6nKe62FEEe1mzRQC3J1abneu4rgh02mgMS918+ZTT0EZ/Mb6xcNiaIDI8U
bVdlSaayTngNrS4nGHWe3wCMWWBF0ME3I8HRy8IGBDUYarZyyckmkm5bcz+mqAny
9sR+3kIuC5izBTfhOF09Saw1MrQhRCsmTeb9G3GjpJwDNl7RZv3GhhEH5maJe0Jz
XCnv2My4QwSmUo2JrjHhDrhDeG3iUrt5qzCCNqI6L0S/EQkJrV2r6ZmgtMkEreHk
gIfOxCZS25AKBAUOwp7JiAwFBqm5V8HrcXDbJQvQptbYijkXPZG3/phEMJiS8BGl
TmcnieECnCTT4fTrMuuS9ND69oaK5tQc3YkJy3IigOMeORS1cpU/p3kZJLZi3rrC
kk3FL6pHxo/1DLz0n4l5BBF0PWxCdhzeaz+6hsabOWZpWcrwWA7JOcRd5CU+7PPB
D6jxrAaKURiILrJBQdX4iLx4TiealfGFa2OVts1vY2K07g5PenE32pC/qUhgt6vy
YADxCZqpA1aAcQhtGpgqMlgk/xNMkmAXMsC6VjSg/asTcLjDIOfSWUhDZ1gLC4+L
zxFV6FdD6Vuz0Q1yKDGDHrfPzTgPQ6/d3VJQGF0eIBFv9GDRG44Jaz/Z4HtiMK1v
AyOM/BOe2f7ViCH4ODASdY0281fN+77bvjN2hvWMWqqL60g/hjpH0GSaBdYdgcDO
fR7i2a6EP4ezm2ZJ2aKJEqQ8XUygt0Dizga0YcozRkPHTpGRkSlQVfsqIuElkQxM
yeA4t2YWRySoS14zgMsYSVPQF4NFLcZX1oyVfUnGTHyIYHMu859A08ZERw65w8d+
fBCytwfATW96RxNN1pOtnuOUpBny3cHzJJTgqnw35cMRndZDI6t7edxF7XckdU0h
5rV4wgHNcuijDVTTwapBTBz2wkE8hUK2STAKf8cKfHbsVIvcMldzycS4AzeIp44x
QFioN4LPYpvAHLokjjmiL1AbZrj80p1/afPyXB02WO2IIyWvmMQLxfRFrYDFomCc
wVPlhFddEUxFEieIhj5J/50AqQqjnCJ87N1QekMRKwiSvvWD3Nj5bCtkE0/s9HlC
PaAunW0BHSQaB3mBe3YS6hge/VXpu3XMm48yX/6WDL4NWwlEdd8Ke3XYZ77p32kc
BR99hftbQjxziTdbdpPujk8ppvxcNiT4cbfJMApZvPqM0MY5fxuLqvjfrgxGj7fq
RFSDGe1ZwF7fB/eIUzqKzWFtfgBPA+vnIw5RBKMem3eWSATtRk0gWC2hjhCt9k9/
9IuYWVKbAGJ7x5kBxP2qEQztrM8CP0u38MTEjdi1HxymIAgR0hSaKhPnIe/XrfUy
lxXeSOqJQ9HFpmIMIn0dM5VwBP+B5Ph7kKPZ3twWaGwFBR1oUn30YsUqpooIoIIV
yL4an/k/FHnts9FTE0iyV7+PVRRLRHmfRUZ/XjQZCEltGFRopeT+5f0ksBmBi7+z
rbxOQdCuFfDEuxuFPamXI2NWbzQfVpjpKMh8zST0MoBsvwDnFZ39FglMg4cBSvi2
WS8IuBR6BHSyQeHeQjnalhzb1A+nCCGcTDZywuvMAZhvqaWeGU2+TjJDXNfr5yTM
N1ZBdrKYdwVmn5qKLQkgNeQVEvA3/k//M8O/Ui8y2m288Pim3enTpGwSXCgYkDK2
Nl8F+zFRJEGFZsvlya+y/aaqONWVAGiEigqoFHik3EmFmEDjN0s3DpGLzg6nvZmg
9OpUJnabvblidWXq96ZjV7Lr58LcFnfgmwxBPwzJxrvpCO5URiC4PDetUh4N36pU
+cy+SdFpvY07EWXqoQkO1/TCpLlr0iHvTpzNUlSfnwjglgf1egzP6Gnms7ETZpAr
tv6hMOQlWhzGuaF8O6K1v/0ftn9Idi3E+R3CTRYYlCkDYuGBwQeZpCBcm3AFQqOG
gxN1qgiUIdtMAvvpoiqjWvelDOnD0fkH9g9dQyEutzKEcMLuHC0gjFiz4rU0yXdO
cKQebALAhenPZgMmB8jgrjm3Qa8aN3E0rZZIQr8App/DGhm3QhRGzUipFzLqwnyY
rWnigtxFOpOxLeuDdlRHFvZ3WyvLzAxExQzs9/dCL77RYe+6fMyDrpZdbcQAi9mA
d6SWfmsw+7jORBl/VPMTUx3wp7ct7qCX5CMKIGWHwP35b+HDW02wnGmiIgvYukXY
iKs9YiIDPFYOQHzSUKdjjfe/61IC/6Ic4eNUQeZuGdlsUbuQgn78vTGWB6cu3Roc
o21GMkJnNC9l8U9U4voZQ/4DRZy5ctGLSJUFpotghVIf0TbFHqaeg4VGIbEWK1Mv
7JjWJXzHMTy/fi17rVpAXv4ms4CDlJcWZ1T9CAMF889XR/tGZXCMesUz/+OqaI4w
ljjNpHmyK73MRG/XvFt3jikHKXGKB8G+lm7exElitzKQiIVW62Xaw27f2jrj5H8Q
AjP70vXeX/FQ5LEOz0r8W7fYO+sOn/YyYt7C+LBgd6zRjAMzJuzb4VLmFU4lSNl1
bt5T7HLbigK7TX6ieaC76Yj/PfruN7sfPoUiXSD3nNOJ5Okxp2gtce1XEum1nYrQ
zDfciuKAe1SIRT/XvR6Nw79h7+BlGC1LjjOP77S34NYNdnpfNb7cxfg0e/0HrwZo
o2dFfJ0YnBkWrOBteiQYKqllHeOt2+ONYIdyuQXwgUEk4yvJi5f81l+WoCD8B9wN
Iiii2m3iGh9teJ+8m34eX6V0dIDmtn74tJ+7ClBxsw+MpGexjxhJy9rC4ehLMNRh
yHlCEir054rmLcaWa6i02KTh/HY9xij8tWnjEQImMerKoS21gRl8UuePuXrO6NNO
GkWQ7zQYMoNWIvbAAor04kZXHsqe5K7eBM2pLTJ+LfoTt6LPQeuZZE4ZOpzA9+PA
sKxsKRYDPOINGaUnykb+xCMR5CNiW88TAPZQlxZSapv2rNjTLMLW+J7DpLhjDWNk
Z7EI7YjyPznjYlDTLdSIDihVKtgCBP31slXO0Fe87b04/f+2wyiNJY5YG3TluWsq
f/FKQukYPwxyRXas8DTFWfXdFMESRbdB9jr90an7sZut1z8NystJdaOGisLiD0dE
WthxSFHGctnmpQU+Oo7KyavdAE20Y25gUEb6K0ULnEpRHxuSA1ptGGNkgw8R4rDa
pawkwJT/V1XdSZZGGd0gIISNO1+F9iAXjvTCibNSWWglH4YBiceJ1dHsVUHn1iTa
wabwEZw9ZlKwgKD+544MRBY/lMZ7R/wiyMFQHXotmoyXD+7lU5YiPpT1n09LTPW2
pQqnvjgrbw/Q+mR4pBiQh3sy2035+bAfMzanwFSG9kXv2wh2gFMaO7QnS9Hn9Y2M
lVrtbAMOQ3aSW1pbF0VTogFS60Wk/GRYEL8QaA4zKkVQZCi1WwgNLVbt3k1AZBAg
Jx4zScewFmACwEoluSpGFnq1VTkw1pXQVfSJjAyafKFvUADR3P6nosL07dwgOPrR
5M36lrsjL4SQxX+Ntb+JFhjh2N/MQR/zx8JYXnCiDpRSQwCRCs0jcVX/5kvufCmC
QQZtS50i5MxPMoXljTsxE3pfWLmpMYe0AvQkoveOOqYDOedePYxbURwq6ELt6Hqc
WSEd3NyCf+P3FVNZ+VCuCnJI/o23jt8XN22/HUhM0YJS32GUzuiWulfIOv62R9bL
13obFcYxIWtWm/mZ4rYSrq2ue0ag73dDziOMMLYDY8TtT9eRMJmKMUWj6IYV6TWc
72QmlXuIh9/bQQsE1LEPQQzC5pBmlIwyjc8wM8l8H4hhc8xqVKYizBFHEm/HDTKe
aLwUpyow/dRa9YF6e+SK3Hj6rNQg98pLg6uVxQGV7H/umr2dvbkg6iPXZg19PBKD
0/u+ZcagI7ULqLAEGsfCPF51AHvd/b/CDjuQaEYFy44H0YQ4Aqp5/UqKEAOdWwCM
D9NnczUZ1v/+XnNNG9CZXwqi710RCTx/kX0R6qVjT6gZjvOFoHEW1Uj8haHaKWdh
96oxnAn4uwnTEfSv1JpHhO0+Fa5q2vqVZiFZS6wiMKiu3Ct5RMW+MYHN5sX6KMvS
dIyg/9Heb1ibdtSz2CREALlLZtJgxxsmNr6ofYypXcQ5uvAIth6a1/WksvND2Xhx
QWXcc4CSbSbUMRGbLsUCNhu5El95mxJE9QfNSNLL+CpwDO1umY0vKqD5kBL+eFy6
C1jPQKAWsh9J+l3kkO/jHNjJyxs5dARMQL5o/A0dEvx2m499c+M8n7qAZWH4mhk+
0Y740k6QHsX96jVmV4ODgOCQdu+rAao5gYtqeCEWMpH3QObn7zm6cwviMTEuwavt
zh+yf21c9jbVY5IAH7w4NuVw/plD6ivnZNg3XnIr1RcQ06BegVAl9Yor1a7UxvTN
ZIj/cbZ5/jy/Foyn9DnWXVHeS1DrcOyLREwp7EdePlFpKoYmzDfHSKIqtGOJ/pYf
Vu7YXKbv3Mi/mLg741PRGtjN1VTnZp+9YHY3HHlOiBIfsFdG1WCic8zEMYL49vQm
+8zICQXqUYk26W7NgT6UWHT4bJM/plSnGUXmVyFUJ2QKI5Bd9V+WdWpbhkL1PiF5
9hfWFW3XTyk3Ezd6jdd+YHA5uYGvX9otlzVrnRkl+s6FO+g2pQxexq4zZCxQJamf
M+GCMh4D0QvANSkRrN0cy6h4hszW9VbhlO9cdrOgd/umiAgibJoXYsHWNNzg+2MN
lBjEkVdHktbrh9yUFoeOKiEasnem9Bg9wjXKjhTnQMMogLulqqiIG0zJJ3r9kBvD
JiBBq9GiDAN/lMQRVOnV1xGDK71bVVlgCfzZEfZjZuEmK5J07FwC/vAN1xUKGLVG
r9SMsLXQyrxuY/LZSs3qh3Q4V7GRfEV7mTAEWuniG8hMpkYv6k6vBgXcHUgi9RWU
K1TVEW/Mo6uzXrSVqoEsI1NmV/cvP9Rz2KZzDG9WJ+ET3wWPyWft7YU9BCMR8P8H
oiyczo3zNSymCIy8vw4SSy+ld4bHtZ0xF1a/dniRtJiE4TREDOXaAcyouAPhzQCv
WsUKDaoj7oJJ0Dv0TXT08hp+PQbayKM+OHx9vLKfE1wVhbS+4KiJ6gfQaUEXX2q4
02w3DxrQLdEzWZxfpcr8Tp8AtrzgoRM1FTy5JfIILNrQbkBZuFANA1oAPIZawAS8
9cACFCtjbACsarSfiZM26bRO/dSHP41PP5qgV5doOY3+M1Ld6HR8K3Q9d+MRSpjU
PDBUohYLuJYfuFPv18iCzxwTHTm3MskMomxzEYCdInpVV+wBu8bSn8uzBjQErGLg
0vYP0FBCvLKCmpc/PA9jx9z/8KLk1CHxZXxUAhzFkvt16dpt9zMv5qZgv5chKq5/
bYDBYQYSBk1vYU98hkfDPeZl4GHJUw1vHyjhMjdX6LSEP8QNpf3w5ikyYyqMlcCm
y23oBKJJO7TkA0/w76mkHpfwfeGMi+SlKkkqt+h/fevE7xr8Anxwa80jGB2vlcuc
P+xZYf/teGpNXRkW5G/cz2tCd3hDq9t9qWEF62bLSm8OclhC23FtCSEx3lhAV+0b
nqf45rDaHpy9C1skLK0WnTrSIzq4fPFeUiW3xi9KEdo+p2Xq7smHeXfaCvgx5rzw
INRJJVpmv5wR91ld5hshTCf1UC8Sjt+ibGQfRD+aPVp1DTxy+R03iLd2JliyS4+v
h1P61JdTrqANkjQ7ijqKTHH0S/YdpdESjy586yZBGtPdNrqmQ0EwNGZrd1tgRY5e
At3aDs9CPBLxVfkkJBUWSSBmdgdvlZyTF9uvGevsHHoJesXH+U7z/DQ3FJLTZ0Up
SmAEBfrXEahr9mrnVM0efx6/F+bKH/jPhYia6t9ksYKc3QVwZpHRhsw/M97zDS4p
+CjhFCGWb4wdGnZ9pMdgqkN8YntSrHVl/7MQZhs83Be33GaB9JyRdOuCQkIx7Mtq
h+pjDlqU/hE0TUvwf8MsqVjeWwKhgerwAujrrwt2xDbu6pzCwqMddB9zZAvUyA1c
P+QfnG3gHC6keWULft5pfAP5CMLwhomD6QJJz110zqcVH/Bf6C6HhAPpK362fg82
ZfcuK0A6nl2aoo6muBt7nNqsSltxMyxaj6oKo9G4delgvUSFj3R9tR+okKALSDtL
s3cwM+fxCuUTA2cJh/AYQgpDsCRpZKgGyd2KlxVhY4R8StQuZpdx0fXOQSq3eM6I
dftDAQE07LzB+cgJK1SgBOsadgOZqLW+PmBHgUIZUSwWyr7gzqwwwXyTSFOOoI1V
obpDab2dHbqZgMykqQ3wa4dmc5douKy6Hgh0TqvG3kcaObJyWSxeMfXIz/r6kO+2
PnusSIzs24y4Dh55fMPdT9jJDFvu7EPhGSsPeNdsuRQ+BLdfAIcFOGYMDyOQYCVo
t+BITB3BByNCwnqtcL6+LcrY+3K5ICtz3TDBSfZoVlcRb6LubzDA3czbs0HmHLj1
CVxHV/jh8TC+25pHGkQQqigSp0fM6AabvBade2qYHNG3XXRScyGGUBF36kz7T+uj
W6tx2chQUAA4JYmfRyzOb5VJttN4oS1ylARZV6IZW6KdlOTaO0QEOLevJZfGzlDX
9YjyI0ZrWw+x56Piu4bVM6FF7iiX+5d4V5oF5JIAT08Pz+ahdCAurj3enfzdiZMc
xfVB7gbqFlpPMLpvO4wf5TX4uUFZYg4Lo4w5N2wgJs7ZYrEtU8FfABXHk5Z/MDAx
W20pBY7s3EsS1CsUigkcFfNIu/zIeZN2NRP4JZ90ImYVibUH0F+ILJxdQ8t1A8ok
6nPUnZh/e2rN5CUnHB6tVGRh2pEXvErgoOJDKYvaLaA3WjP1C2FXm3B6FC+OGnar
04ePH+keZOB0RSbX6VKlLQ0LQCt8M8QlUg9go/Jq2B9yHTl6eREnidGEWLs2QZAm
m3KqXEDBdPA3KW7DwDC6Nl8im4PuHMW3b2NYLF+CA7M6EHFidETuYg536PhO2cgZ
AXTH/V2JvfvcgKPxwmr01BrEAtW1bvutw02FTnqJO5NMVg69PPvdGU8KbTYY4JH+
ug7opodUvnQWP4fRcm17J1srmpAYVFAT5qz9C9v1JoD6wnkou9bgCBxTzvGXiOSR
qveKaDHdwD5WQnkYmsPrM9RgL66V6u4pNzXyRC7ts1AAm6m9yezX6ziUp/qF7Lyt
JlzG+A3gheUvaL2zX4Q+NItDOWInx3KQiS+2PXcB74m/z9dqQpse68BCLEZwqVxp
8te/XEuCORGQ9ldAStvC9Xbl0ppSMmA+dSFAVrZCkPRdu2EKwyMVuRnQ/akCMyeb
JvO945Zh6efLBnJ9IWKvB2KQL/AkztuvtCn69+Tt+SNDM+7YbGqphUPyiwVa6NEq
4/aqEsZPdejvK11MJgYKsdOTcCBZ4aJflxRwCOBrOwShAWfIo+z9O/BxVws4a6J6
gQhcdWWaDQabGcLJablHGr8LVCNk2Vvqva+UlLvxU924Ey5LGD1qJumMK5Clyxtj
rPMHpFtPlhUhsUHLzqXx8Rh9E25se3kVKjyWEt/4Y0KFCsIUw6IaQOVvYgcjGSCL
uTNjGwwiIDDwbB6ruC3ZTZDbAUcVeE+FeeW2l+D/gBz3EU5BDl6nw6yXPFinM37u
lv3JAdN9mLzkCBnFfecbSsEgSdt/Guml+Mdj3gUexYfa+Hf/sNhK1bDh27fyIv+8
W9ZVDOT63ip8xOJYDQQ/Roj7AHXenqddaeGJOiTt8cHmcH7DZIuATKZHunNBqXXQ
A4sZuHpkpPi40M4o17nBEOdNZb5Dqlg4XC4rhQB8okg4scRzqilzDdaObEximT17
MO46zgX5UwtMVDY8zq4JHLnKcNtl6+JHg/xOYKwncJNOV7VKj8VQqSBi7EvJ7Qtl
E2qOFJu+iibQ3jqn8mvlWw+IUEev+6HSbiomABAcLdFAxyxrjFazmlAY425qBov7
K+qwW0BnZBY2YA3PzP1m1TI5rBfbnyriQ2+zYtyldZLP1cdiY4rjwWU4h54umJ1V
8hnCEFzcA+exCWxTrfG+6DGn8aWlnDU15EFZYY3fVg2nBMupFxUHb0JaJF0VvI4Q
ukPCn6o37Wwb9a4usHn1K3QWrtOuledhjm+4X3h1SJSYehhACG6WUZ7b20kSM7o3
ZCzHYoyJ4c61FiWKqCYFJZ7okWx7h8ECrcKm6R8/JxOpIHrSg/2u9YPlMh9FZqaI
FMPRtzpqFW+0XfDFAsOO5S7a/qJ6w3aVXZpQPitoEZAw8nNhwQ7a9ONo+2f3Agvs
5kOPBNZgMEpimFurUMvncv7TkhW0OH0FGzCR0n1SQijY9F+Xi5pToziOlZaSFFF9
ynW0zh90QtQIJBxw72DOvbTPESZltDdb7S19ovo7rYyMu8bB/H5gr8UY8uDi1ml3
pvWylBMcDHJiuqmpM1AyhI1ZXXHfjaDXfDf9WR2gbqZua43+WurZVhRZ85Pi3Q4m
Zhwats0313pH61rqFwhe/j5tiAgEm8oLh/VpwdQl4xDCfe4pjzY2iTmYdHw+rex+
rHqp55huKPoWgzTQCtpnqFhk7WkIIp9+z66/er46XmfhLhEKEbGGXKzFHFubLkXC
ZfJOS5UwIHWDWqeqoKvjLXGTjmifoyOqx3TifJ53VWK9fg5tWuMX9XvjfbTEAzQ0
YnMKxg1h1uyfQh0jmXNDadNCyK7WkJGiSTIYQ3flpBwWWyDE1/ZY7pce3eyteMD7
Vfaguio5L90++VuAJ16QqUUXE5k6+hkc/g8B6EiSU9wzCgIpKuHEj2QEbZlKyKMt
s5pagtX3pXWDfR69ktqq+6sr606nlDq0TgmqqD+FvwSSQbfUB2WGbvI4mgqt3S7b
SEtV3HzmJ6eDK6I1ToY4HXSthW1qVSOM5yNYQ+AVVTnUgo8hYpywVd3ppB1U7Wd7
TUCW54bwL+XqXGVQw4pJz9Z8FBh4lB6R0Vv1Erhs/b1U+/Z89Qp2Kg5Y6FqDD5Tf
u9sGnbeJ7KBt+G5Pmynhre9fc3uPs/LUZkikUacsQua9gluBbGMa1PMchuluBT+M
kLQkhQ3jTVH9WP5BGDJnHePTcO6iBDnIcBFVkp+XBqoUOCvrRXxgyeJyGccfw0qw
5wMUJqr95k/qGzrIBLAr58RwOP7ekT/JWQvqH+jM0DhkKdWn02wlAAGJsF1korWv
iUTP5w/0nsSe8QPvrTlZlrZXmX22emZ1k2NE3g1pbN5Fh60+AFDI31fSJeajCIsG
QOK2ApiLbeFjz6GVZraqai/ld6FRnSOCdS2CuKTEzVz3kOe4gqbYR+Wo+SOvobVv
poFTmlj+FRlhPFFL3iN7qrqbdtUrU8jGukhQsYIIh1hRuJLKEYvOfGCtyaPkzclQ
ty6R5/tWSEv2tTrmKIfSYFPT2n0P4yOeBMtQ9sDP1B5kbs/tL5z2fW1QwU/k4qCN
0tAMSRQNhUfLdTd405yUQXCQ/KOtX4Q58U+TYrF8RnvFX3F3BzfZWx3CaX+r7Y0R
R8Gl0SH6DIuUZXgUABHrU9uqg2XgxfZBhnLRtHjcyf0OVdO00KhmFF/qtiW5xaaz
eOuaNASwqNE2J2VNOZdi9/sp+GK7IgqqH/eoyXhP65q2WkVL0QN4sZyCECacZwJr
4XhSZP6jDqnqIweIr6VifILLqiJ4Kz4rheJx5bZUELmG/3q455ZdV/DSjBTjcqPR
P2HVs8dacP3GXBWdPA4a9l8c9AJKfnR7fQ+j5OLpjNTuYtigjT2anY7gmFmx0hRK
5YWcCSOOjT8bzP0JiO0C0Fb58hkLIq8nCuksP5f4wwF68bIPMBRyJyZvMsccdajt
8XpVlhDaKJ0cisjElqP6On2jdcZ5BCxV82ODA2m74mhz4a9QKAkTVy4h4RL+DajC
XXnP8oNkbbcBA7d0bKxElCM2VegD2swhgS84R3aVQnMlH+GbBgZXUDf6c8+F6UMI
3wD9a03cgi+9vFvBAXPa6SzQqJomtq1wT50KbgFJ2eccyRPdXxHX/LC4rdGHJY1Q
kULUeyytXFQywXF61KnpsXainiY2SLv0QQzE+5eyh+5f0eHpwamUjuXyFUNHd2uY
IvPyagwovrahEUIXkDUgF/8niAdcMuA7JXOoD5pDyBd9P++asG3DlZ02gwFoW8z+
Cb6n2c9B9Wq8oiHB1oGRG957p0k4x72vz9L9doS1V/bOm1NU6ONGz40qlzCy/e2j
ONgskVQBUVE0D1MBWRGyMBDi+m1OGwC4EDARjcQmw8U3Vv5mUD+m4pDmgD64jhqA
PqqKRHcwcKvsep0uIFys1ItyJFST6eqzlvou9dvGL+2+fbtfvQUFVhv+0bEzTjeK
pchFS4xZLgcp4xaIsJYgn41nlAdFP+8Q3ncaifLayfn6kdjyYedmI1U6ViGudR1M
I0xawCyUd+Zgce/NI4ql6evcA6clHJnOlEpIVd5DHN1w9kPgg2qelwJ4N2NqKQBL
GLqO6sIVcwZN3fj1YFKxv0657iCv2drmlmNcGbw6CovjXcIDALWCs1Jgx3fWmkJG
A9OIxnE+EXZWg0a3sqvlMm2LX6nZCaNris8eLpgQldr2pSThWCal/TZvfaZgNvGw
G9eI/ngBYg1Xckzdhj7lRdtXCBNw1/MxJ1g6uGq9d+H1T9vshcSl8m25tY+YpWia
yyTihgBLSF+RoWP2KWtB5XvA6ykizf0sTzN+RHbov2SNrNH8ZzE3ScHF2L3ENrQ8
zPP6TzIy+aOzWxWNgOLoSeg5nSAKoyvUA/O/nHZUxRXh2pgS0axOb2771QpzNuRB
ANDiwtiC4Zihk1OCsPmsrtT8zWNG2liNt/8I0B/pJQI/UdqY5bnkgJu2J2dcgfhX
Ij3fvYTKEVIHsVPnHEK4dUiZWtWVGs3gH83Cz0eDVUY01vpvPgpNK+4EkXx29XfK
oBOkOMw8V1Or/bPpV+dpPT4qMnGgA9BNHJFa0l1FQ5kMqBA3Hq3yKZbEGyhOS+Pz
qRhrtAkgEPX+WHC3wTYL5/UEhYiEeP2e3T1RR961SAHnSwVw+osbbdfnC/L6MNkI
oqA94an2yQOKToatzBgitckPS/Z8e9Z4Mk6HWKZqXaiXJMS24+PT+aqfn+Ozl1ee
8Mx/ZNFGIfH2iv2HwCV2abju5pyhyfilPNfh8cveD2pTiaR1ERzrhh1ABA41L8Ke
Bp65NA4JfIiYFvO9wcbFOb2I4iGrCvfmdT8PjmBVmVTBR2IhkCQaGu2SZflDMpr0
GKEQ4a3pmEQOMkT9CdC54Bfkbmwo+QT+bBXl8WF3/vEalmGbV07ChldOMy8JE9LE
z5yhc6bMeWfM+RbtUUxb7vxE5GEubNV0Uf3KYfGCOl2ZTXs7jMBTCEaEYto+2feE
LWqCCBG84Mb4brMGXmaYaJer49j6Panham/EaqwwG8mx2O2Dr41tF3dQQTm9BdUq
66MUa1Bc5/p2NfMdniMe7kFjQ1ubbFSMbf2diphhBxsgwuKbYy74sij6m7z3trYj
71CsqNjyWA2mdMhrSF7TU5AExbabsV9+gwMr28SMTzMFS49Nl+teqyC2rnQbCjBL
n24ggsy6f7oBaWcsmhQGZ2AbHX0SX7l4TwRsFLKzjXoOv00SAufLI/FK0cchm3zX
7ECg2TrNXfqzzL0T6XZkji0oKDuSOcPxXmYF9cXiie+izl8R3FuPXpl5zJuIbeKL
LUvNfijveGn1pqe7JFwv5RbxZ303ptuZ6K525tgJcJE0KciD4UOgo1datoxfaE1w
ceSQrKiOZCAoRTt3UxsObHcQqvcT3BtZJ0hd+1v8FWZXaT1tCMe2UqbDDa+0ssMA
jVUPGJGorkNMCXYThmx+szs28hgCj9M1rcLIuT8XlJTPe3OYV5wEyKcysLjrpbPE
GYooBKEQ5oyxG6GpEco2Yk1vp8yx29qKdUSmmMXccjYGjDb4Q3XqFVDuu5n2a8go
vWw3absS5mqF32ekrRLO/T1DjBxrjSaM1HBtI9SYGlVt+C9fXqNVXGCE8ENnlS1m
6GfgeSoxial4nXexRyRZFBBp8daQpvvvgK7FHtCQMbRg6tIlwbkDlpfsnECPnuji
Hy0avVPNO35wn/cn4JOTAYfQkJfRySzThEfU0wXFgjsU3u3JopPLDPn1pBx+qc7r
FNzV4e5492ZTiDJJINrIDNAU5gthjEulj68dx5LV53KQCgDFH5ANhGHOaqYvI3H3
gWEob7dT3nL0oMGoQ9/jOXxgifURlazGJj/RWLH9CdNEVjwz6dKgfzBrIcdB9pTf
i9KI8kEaihbvAbtEnGxlu87NdUxD1FxbHybd9qFqk4c+V3Yc+DhsUZp07w2NDq4k
NcNCnU7NvFy0QRY+08ygiCoCoPD8Mdepxx2ram0ehLvGTi3qt6Fp6RWYsvENq6vc
x9tSJtrF9qFj8k1Z4F8mYPGYzU2NyjC/IketZ3mLx0NaJImxfwqJQSM4o2qR5Bfm
wEgSCBmoG3GkLcBSNfVjf7rM1fRE+OQhuFj1P1sHH+dKxa5yywBOtchBYdJVxSTU
+/k3GM89+mh/okO0ZzHZkABGUSEmmyCsHWY3BxIDaQ/Xnlk//p9HQpkaJdt8Aooj
F10f+cm572CRn65nYepC1mjFqHBh6ii+qJuuPdPypM5txFMlnWjuYtEoK/DWIeok
YBJOaZX2nI/hEHzoLNVU2Q4CMQ/vDeErwitQJlRgaRt5FnP1KV3wNftyapW8p90P
oq6nGflaiFqAezaFkiNzlO1MuXdVjvygSyT+UGYsWHuGz6pgMYle7DVGBjD8bo64
bXhEQWKKkZqsTH0PkyhgLbbXco0ZqMlGG3I0O1PVsdHZP2dLFiT5wTQqaf4nmVAL
P/RdTUodAxRj7beDF78LD/uzGAx7MV6ymLIVzZQWKka563y1tLx0FpkmgjajsU9l
HaMRyC0W94g1n+heM99v0TGlZTEi5eVkTniR/BzFLFgrcx/mOoCJbgzd9dat+eFb
ho0xhu/LDrZRv5Wjxky6SikDyDAHhhY4aFA8wkDcjOchW3HGck9RUQ+STYGa60is
+CgkKiHlxDPpRPPDktF+AGUXqq8girqprpeCRcgwWf/k28EWX480LGavGawe3JFu
7NK84MNgQyamjV2C1iqcUgdEnFWCF2MMlQoVjEbQUIWjmUIggwXMLEl8uigx0EqF
+2GJ11sE2V1U+uSIEa3U/0CVK2KIwAcZh7mZY5PXbeUvGkfwVCkbo81i5iSl2eoc
/e0ZsKAwRkkN8SGZQPcCCD01B84YeJP03SoNZRvMpvC5EXeEGRZsHRpYIZjRbWrf
4F0RXdS/xQ7CskysllPjnn3u/DLe4XEyGf+GVnYu1g3NBOp4tSDuorWgRNLvr31Q
g/bIbqAZJ8nNB6dOdwpTS8fa3i1s7yDXuCsB8P3Ve4zs8L2xFR2nQ+WqJLBxSTQj
0gdgC0Djii4dPW6D4IaD/LC5/HJ6wkXrK6rmANBS+TqoL5lD7mhY+CXmP0CMVARC
SOzAHW3FTPBhb0K0LoXE77ziuUq4Qv3rgenhVcUvcWWCwY72z8fxFzx4xMrZ6sTy
LpiSoYROBDP5x8kmCUXBIOLjDDqd4g9RN6eBM7uB4x4yXmROCmLLlgtyYhtbcdLE
bUMz8u4qeGYKUc9uFr7JkiyLi2EG7ban9B4otyZa2WQzt0tYygDMEqcV0p8QAe4Z
XRD1s4LvFAYYYaqX9sceE0QZAfPmJpSqyCcTG/R/VM5YL3TBD9QpTiffzQqDjYrb
BWKIHVdYl2SoUrS8QmfdN++WmOFk3dpw3AIZdA7sTFkTFN6eutLqyy9wVyuD9H10
n2upP2wdps62qOXH0dKVsUB8520AzbEJU6a0TVDF3TwmwC+1I2x1GaKf6jEqiQf/
3/rgHVqHF8YbicjpfmO98EnbHzv5pfWSgWxjFg0jrMjYH/D8ZZZ1ROLwv34shLIa
/3KFsV1Gtltqj2E/oNONZm8cao9efPaRW5ir+Y5P5YixVgH3OJxlhTBycDOWPB/8
DwhCBOUVF1wlzy2pznBu140GEcHYkxxW8EUaVYmmx3gos5yDp+2JOX1fWe1x+t0P
ieG+oeHGNmlzZK0aXj4HvJHcTTDVCti0VgBprFLQjBAKSE8IohMLEOCL1kh2mUC2
KEQcSVoBUfI69VqDJbr+l8KjsEn06TGoNw5fcURQFhzrQhlExoVyYVc/3ckwkqmF
Q5aV1BZyNJCi7o0DvXDnj51xhcD2XmUatKWQFcD5oLHZhSWWeuomgEBufJB4dfyx
E5dMj7tYbib2smBFFSOCdIiytuCSzj/YigVocXAFEQp6ryc64LENMBZEXWeGTiZd
Ke4Q6nCRzg8ybX4e1yIWX7KV+RKSUNAyOtGwCAblXgzXqpTjB6cjfK9x2KU7zLlY
AE8PyVX7vfekaMVApejb0Dj7W5ypajGKuSViSfnklGVkzGMnytW+pQOC4gKlngcS
ptg/l2rPHeRqfMTimvGEQ3iBMvi8ar4QRXN+01yMLemM7l6+M6YrMVvHRym2K09b
RdUwlfxz35eAwGMlB0zgBDyfzEk4IrurCeP4Rnq9fwU714TCcCtqNUuvHRPnjK+b
F9ZCIG37Udm8ubgLAKHTDQWWSGxyDBPzjfWGEimoH8ZvxeNjXy+McsvgW5s+z1V0
XfU9yqpyDx0Bl2eMtO9FtqSDlQZ5tdOxIz4zvogX1iat8ElohcelhvjaEXR9IZs0
fyDTRiKvyVL0sG4k8Nip5cmra+PXhMk9ukaWZLeN/bo+RuStLBhMisj2FmC47t1V
5mDzxNY4K3Qrt8AwFVGWsL5HC2M171IPgp2k8z+otJcIj9OySUpMezrf+LkGRsP6
RhWIQnCWKy9sbHkH0Z3yb86W3bFqhfruFEhXBBClBtrtRgazHrTaVKVCn2gMz1MG
WC4WtF0U6w+Kb8ss3VsJMAkhaGjIKT5HDgxmrPcclf0dMfLjJf4pnsykbo5AFVVz
nbv4lK53A2TvRGDt6BvDdjsxlkF12DLwCdLsFNobyM/4Rol9c7MPc1GIUTpOgB13
noh6/lAlGmGc+Mh88dY2sCXJ21lN4vVdAK0A7f8RjRwofPJeQ9frtG+Bp1aXLZYx
W8SVSs2XqVUup53g4mNpHs7nqeZoknYQJnSMDJRQmpdT7oI3CfAAjL15PV1Eumb1
sdy1/uF22SYhbSlN/xdXfXCXl8QLVO4VZG+QtbGCNRahtGL/OVxmcts9asruLMQS
N4n/YjPVPFWDll6gxO6PQgySfJWk8klYi556XEbPCslQQkYNpO0vVDtW29E/BoeT
IVas/6nN3EF4glr9LZuARIfbUDRZtYv5FtcI/kVlsVacK3NtiVvpcifRVk+v1BcQ
o+v2pcPKP5he79hROxAoTWO23nCDnAKjIlgybGCTmt3PtGA8AYLP3g/xHa/tG0bg
9AN5zrpYFySEhJptVcY3zqz5EFGigrJmc6hKNfUXDctiYLn/pqm8eDFhP3k0tCSH
4gyFqFEkJZRVQHne4F5pWH9cSJIR4bUg5FrWc4y6mNsHmrIEbQ5JcJTnxDSiUkGA
Hci1D/LVrXtnEyuUKsCcich9uj7bthIxEGJ8ppisYpqwH2eqAJyb4Yn5F8OyjqZY
coQvXc51RbvTrme4l73vIkijptx/tGTAooFalZ/iA0sAvrxE+iZSrmS741FC0T4W
cuBPfHoGB8agAFKGzANjtS6ZAbu/beF0QP1RHIrBjjCQ1iQ88eN6KGkQWeF23i7C
pSXo9CR1YMICFdwstQmbrAwQFPl2xiriPJC3RvnMxI5jKNQocA20dWOgIYaVu/HB
uEsWgCcgeTjIyNXoqwzLczmIDcDPkJ1BLedmSTQ/VsmYGxiUR27aduOY6u5tKhPX
y7Btbz++hV2Z2aPyNbW1q5+59QCA79lJH5lvaQCJAzW8ReK+sHn217yYTDYTCWlx
VTExfjHfHIjQx3aBficmvsSh0tTu8v395rbFDyD6tVmRzOtfQmfxgv1MBG4d4CwB
bR0kVDCujBPXWMI0XUX8ziSiG+TdY6SSIv65w8uDwcIQZG2KU8Jx2fqWqIAlB8yl
aNDqIi0I+c86VPzIegxiYNQjAPeWU2+f7kQtySe1c2RkEAs+1QDimLZF7EFebo+F
Zekv6JDexVy5HY6QBwy/0Yz1cDVxO6WNIKWVfWVfczfWSYV87MFTjEwwhlENSo4i
zmRxOG/IbP1mTYRErHW3ZwySL87v6dIb53tZYsAWvKGPT7vCoDGZ1zGBhOhGXa4A
VEDYw27MBlT8ulloAzT7/8ddM+ZqYc5qscjuXVoPe9cRuujd08o/tQlpupYwnXub
t+M/LI/W9JGzEaFIpzhT+HxCwUc/KlgM0bd7zFp+Gpe2PYPSAkvnpanImpnsmVmN
6d/iX2hVOngn9IV1R7gHVb99kAWqWy5Ncp6uGgyld5fU3McoWyEPFX6NzsTkqMES
BKZgBxx+UF2dnwL6vbWSdYaIuEzaXzpjGjiah8j538+FRv02arHxQ8MVObWSYvbW
qgJ4uOl2Uua5T7M/BpVB5PoxAopwmhCDST8gsJ6U65k3s7ZisPBCjmHjIRJ927he
gVzRuYtk9jqZ6Q9ufGe47MUU2fZsCI76vmyxv4Ybq9dATsjaDi1HNM4Hp9kS4eOI
n7Wq1+n3/p3KWzFXRabPrbCeK8ZPhS9B2pWQ1j0tjom1ac1kn4OLmx+yaZUXtcr6
SCgean6JBuDxAOyqYHHW8V2g+8nc97b+cK6r7A9dVe8=
`protect end_protected