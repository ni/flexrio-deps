`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4320 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
GgG2UXwpbWAyDgGIJC8iiNXL3rFqsxcHhk+XUbcSe82b6qJjr1WVq9PsxlEuc/YB
h9UUj6C31qX47/0sXZMKJ0JRb5/NcGFvZ0kYNVeguCD9tUf/Yig5sdj1lUf2p+1z
7k0Htpfsr2z5O36wqXylCE2Wnkc4pSg9BkaJznP8uGltq4d0ASijzr3sUl3MuXqY
+WaSJFTm2Kri3tRhelND1j3NXxdGN/TQdxRWU40Z22X4vsusQmyCVjSbB+FdLaQl
dlclpnclPLjux27x6Xnd5BHEEpaC0KOYddFJXXEzMnN6FGNd4afnEAQ3KlEMu0dO
0VdQQQw/cWkd+Kj3Kl1kHsaPQNvXMtyV4nEyBqAmxuE1jByhcSi+s/OsObmup6XW
ozBRq9DBVfJ0Qw6gQB548Qxc/vDx07FHYRFYteTKCU8nDh40fjJIBH9plxROO1cz
+GZZZ/ZgSEuPGNk0cGR9fWSWetvrXroGYpHlE3ylHt4u0dKieBkQTWaDfyc4nI1P
Ikin/0UwxzYHTExQQEzX9nJXekb+2klXPZUNx0ZQvaUlcoLrw8CD33w0kC/K3VRd
/AJbuEJB9i3u7Bt8X+zZDuMNoAsVp6GN8nTIONZbJJWymz/uOjSUl42R1UM7ARik
VJ3NarqNh286odhE2M6w8entxIb2aIS2UYyOdm9O7dXq4nqkoIcEBiMZ8kmf3wpD
qpxjalc4krrKrsrdeaCiXPD5Jb+IpF6Ha++F4VUG+4MXGrmhvziS8433cUHwKhLs
Z8WrLpz0hXfAQPPr7wmsAKcogT//N04SIDGwdWzygx8DVCBHQL3mLXsKob+k2+xf
tLzI28JpW7LH6eKEjije/hVYZLkeoXqbOGIXknT6E7aELPclCi8HOlKNQQoqGBdn
mpE172RPxbdTsDqPQVhCgR4IPiIIdJMZgRf1kpaWkrxTMbozEVUAjE2dj2ufS+o/
BVvABKjYZuuyvwr//N91+LG4Nu3m65J0YpOkbeatGTJ8sQeT2mz/Lt0pJNBBCMWB
HW/7eCrR1pK/oDlmQ1rE1AOhf7C7VZDhM7iMOFueWjcGB9GlX4BIdvws/x+HReEC
PsXJdwMOL60g/RwjyYs0vmVT8tahIfd6XUIVawnrcJVWsJCBQMeJx9vLEwyiqyP9
UHbS/ptsdVEh3MRvEp2rOVHKbz+HKGJQO7aAGYoC/usDnfXDUa5G6b3pRtuRFG1x
liAAhJFrgvx3Jlb/RDlnqjiq8U55/Z3h4yH0cIwwYCw+ljds9XJbne16cBUbiiMb
neIOL92GTQ/tVcJ9VYopz6Eqhs4dZVJvTlvsok3D4VtqliKytD1FU8gVtDRKtqvh
M1ieref1KR2gooEYwbWGSbEjtluo236wDhb897UT5n0CZtXFz5Veh9DG2aHKOzWt
BKCBebPx7lTiUFkxK6d93h8HrWnljawCUW1teUNCugQY6x+0pX4oyR5ZBJHYSNGH
3EAh1NQ7o+LlfViaeaJiq+qRPV9Ic+RSsB3kMgyJTl8ylGBC3C3NFR/Vpa2kujmg
ILoHXNYLOEoIJxS5GLx7WO6N3062tnqqIFiX6wAhvpuaavXz8Z0kOWG6eIWDDQmH
a6PMolX36sBUYSkdc40JjtuzWyEubS6q++69Xhd7FAS/fvyA5vhFCiC+BfNAVk4w
0qn4oW7BwwxOneRtGPQWj00yqUEPknC0xs58iW2ScJS0YHkLjVh9Dt+Bb6UBz8EK
5sBp0PJA9PcWnIN15MmuBwsv59lrJl71HM0+hNg4fWlAno+XmuVgRRK0FmT4QOge
QZudfDNjYZxFtxXf2FC0j80TED4F2XK/MPqUycrMpwWgatGw8gEz4mTruMXIdMX/
ORosB91YQS15FGVUCNZdwUdv86KpcJAsvG/L+fxHKpyKxBXs1PVbC5jmwy21GUZj
mR/tpxqheL9G+yJX2jFLPt9koj9sPJVxqnJM9q9hmJwPmdYqCr8q3w91CayLW6F4
6pLshr0IDiMCnLMwU61GGrAbFCypyl3rh2EgJJ2WuxTt5Jx/88SMlC97f3Yp1JA4
FS+6V5gXa5CeJaAbSsyrCWEqYiUy/BzTdVDj28QRsjCDPU5xpcDGBASWfztv2QzX
9gENT+O26j+PhjNkTHCJQPmI5CS1FVxYo88A/PYoVtAOw9aRNDRATKFyNPIuD0Lg
jVHeesUC45Ko12tNLRmqPVdAlHmLdbqh0dsTmXuzkaQH7RIQa+S5e9XS5U8N4rlh
Ts0jxxqQvBqMgGSGorupo3HJmPGh6MzMZ4VU/AwPGBF67maEWS3ta1NNzF8t2XhQ
ljJ9r03mDFMY6AsS8B5QwV9hcCAHb4+mdA7PfqoZjsGkmidtidLdJDs0Ek5id6Zp
VL4dfReUwSfDTENM3+V61hj5qHkY5yns6U6OaPI3Nutsn+ircqff4qmOFOCPwiYt
WISqbu08j6E6Hi0JLu/IWzXOLPvdbrHaw6QJhfwjEUDs1RppUWkr422suO0OQ3QB
hqQfIDfAy1GPwWVMyWwo+XFyicD4IpuHSZ4hCqFd/lFG1YblDYq765lkkGntkbsV
szbCunr3PGGiblZtYQLzm1fd8PoW1UI/ogQTG+0iIM1CjYxE/LnzCxKWHrzHLx4Z
fo1Q+J2N4oWfqzAGui1vZkjmiWzIN7S5mCUXqGKUbaDrXYiXvBfd9kzVy8VJljyj
8TYO/hubAZdrm+jwffpqbv7DwoTvUef2y84pKMoeJCdtXnX4ECeSl0S57asHUUJr
o+ld6rlBZ4YHj8yjEC8ejMH9qGgNz1EhJ3Hx5IvCdBtrH2uYt9wViB8bVA9uLv/7
kC3P1V4bytThgxdf0Ceuvwa6+FT20Q/YxKUCK94oyT13iQ5NivfuFfJZiiigEIei
U+7809+vyto2e3PArwrFpyDS6HnsWLlGjNcM7AkLtXKF2eStrz9l7ff6fTeZ7kEy
ZXBkyxW6UfNBQhASoRsUasraMTBXRiEDa8KQQiM+htdVhHqEwLnxTIVN32x6DrRx
pksTI5QfOs/ILS46SmqF6LM+g4Dpi42OQqK9Jx4kFRpqLJHedjMgf4XpVa9bBfz8
TYhkvG8pIhHq6XQpY5Dog+nG8vIaC30xab5/rg0WewOcGd/CADrjxV0Ij+0VRhoR
I7C46UzDTtv0zv/1zPE5NbJ7DVoMfmf68xkCdIFM50VWPWjtk73k2kYPd0BFSLOg
aUcSPsCATKLSQGmg+gyA1D6vLoIboOXMlT6tKeWo6QnsKM0p24KwL/JnW2aCqSx8
WlLmhQrpZJqwXbxS+3cBrLOUfdD2N/Xr32bgLo4J2dbHowYmKOWzXMBl0/pFD1xm
4XobfBOqqryGjCVjfKeTEOw5Yf6cFyMky4MUhrNuzb3dLOO12PyYXcii0gTsBZS2
Y6RnC09d1Yq/eWSmnxjnPPLLyqcb/d+8LFteij1LfM9H+kNUP+dZ5P9BIDU4Jw1Z
qkOUI1dG1ZWSO08u6JP7Ymh0iuSe6ZTq/WpKiqgJP/HddfusP+p22Q9OJQh3JWsz
bZB3q5VUXUNWTnhUEd8KmU0xGEL77rc+VynzWzu8qNp3VurcajR3LwI15hb5K1Z4
vL2j7uxuMLNrpYaQN/2+LTaSghiFaNoLJe/wPeP5q6bInGx7+XPL4BahNwArqF2I
m+iCcUvyvyqhrNbMMSGoG/SN+StE/vpLu/D6vc7cx+K6tjF46PYhqPm6qK3kmzrf
WBSHUfQdsd4Hro6dSe1onF/0wD/YUG/UIxQf8yrdrP0kZpeDJ14DuaxR5tDeik7v
uhKUFEMQK5NHumSK1z4OVAha2dFT1Ux/UeFv7Z/WfbxlbcV+wqA1rH9CnKSSiWnQ
Gx+/DVZPqC3p5Z1zCiIGl+gVkxet4KneqP4WpyWn5KUINbk4brJk/1QTsxSe4Si0
k0Z06RZSftCMvL79JEPpyW4/4wpN4O4cVgh65rB4TZLjB0rOB/F3DXQ+S5qGbMDI
SL2y/MG0PZ2TX2VtY1fVctvp9IqoBzjYMuq9lYiz5VPcKD/9cQ1OtJdma1UT6Snq
4y2PQcKyYzbtz5EgcBf9FFRXMkzbd5cJJgiSkKVMAK8332pkjTJf0vtmWIxvraI3
S/MdtZI/Ba6ANc7HYh75ILnU5txJKdgSE2ZHBdh4GwtpnvVJEHByyZuSyqlj5pGe
4gFOKo2kn1R2UWZnDKnjDZUyt9EviiagUcvlEpiDhVEnnx5X0YGcLshU7azw2w58
R6/X1ZjrlEZf/w6mxlupBzzi1kH4Pd0jEJkD3yfUjKaUEAijUQ9GFnI1GM721JxC
4CaIeQfPzWVM/vgEfYaIaiSSpKGiykYMSkbLWGpPqnZYDVVjucKCXizJTxSKdy8n
E6xzS+8j1RCiVih1Z42tkRcQR8ur4JtRFVndtsKV1uoM2uZNBDajmkOqhfN9db7r
pXpPAgtUq695abxkGT6yAvVjpe5vDWiD4sNHsHFyllz9niRS9eWbtJ23o1KURkW1
6Ov3wHhK7CMNvPaY7kTTctKFkL7l0sa6xbJOlvTQiKM7GvnyXCchlL5cSw1AWwup
fdgYT2qdOMqRQswSqEBIzEC+yL7D1uSTkLlTPdZUD4b+zW6hUnjanaxv5rrpA8JT
4Sz3+DidngZrJQRjmvOkexDQDpInhocILzIqYxEz5PVPEbS26In7aCruE9U5DQXU
OiUJfXXcmCXwj8ud+4/dhGr1PVb0eO9Dhh7ZuhnjNz4F8/TftGJ8fkl7yQ3AQC/N
ihuEVxjB4jt4t1vunBMHYRrFkNUojX0i970JHN1BYW5hwOkwB/htk8SSB7GBqbA1
yZ/37iXlVwwPMmzZgx8xJvbQLdHqsFtbWVxTAdugHf1l6VsSAGSGY7GsafbiC0wo
RFbPFqqIXWlLWDvOpku0PaHd7LjxjhSwgE8nKIhBvI+ozgMDNasDLP120LLgpcT0
ykRVH5RufKkYIL5rnBjYpA7/eMZ/EqLcNhXhmgSqlRbKLXZ1qi8JIJSZi5DyxCLh
nbg5h8j1S6742ENy3t+mpQI6wiApirvgzZfzHhBA4HDTzoFiBht0nnc6IHMmOETS
kMEixYPJ3j8aBUZJDX3E6zIEESySETO4F3B0/1XnRWxLqLetzCkLt2I/PGvLUrVk
XLvyttjjENOLXIoarLLItrA/jm+rCsUBO6220XQY23RyZ5B9X9mF00TTOQR62Xbr
rMk0TLr92uNVORAVWbiRkEiGqZrX1IXvoxtugTKz1mULTILvkyEOtUBaN++9xffG
cWGDmUdZgVDyU3XArK+F8W6ld3pI67YF1r/bbzt8lDhxXcIB9nfvW1ReewVK4e+b
kayeexQ16tnSeuHMdr4IT4R3Wvt6FM11QqaJ/273GzzvjWFIJYnslaXnqs84QgiE
tXNLIRzdV1DV8qpwgVmD34cs5S5dcGXUEcVlxWpcD/1Bo0ykzJD5XCFL1d9fO5yI
dAKpppesiLBa49DIsIRPDr1/r8f91i6qcoZHnmTmVB29oq6Z7xHbgWOd1wSS3SvU
A/xuzaWJDLduhUfK6ILyfg2m08OtDmxVBz1aRn8WBHEkwJ1gLyiLtFv9lS9IKxAh
UDjVuxqRPmXY+sRbmtysUm2bYUIUkflR96reA81eF0lBOQJguLzbGogWaOOcJvLa
`protect end_protected