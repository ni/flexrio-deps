`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 45040 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
EmxAgecO7UDIr+OXKjjkXBjuGCy07FQY9JsUs1As/EGCZEI2H/GLSYvXTEhb82qG
/AgePsDLeMkFubBU+go7IJ2YSiv8YoYDp2I06k+Np7VBNlGklJ6wWqIunySw8dny
iSAhcn8qZV3mINT7xERlc8Ys/ZIgPpLlvP2jAF83IP7NypaYa1WFty2gnbfmvcW4
HrzEzRfNytKO+Xc1zv/Io0p84Q/9YfM0VIwUCV5jnSC/VL6KPr6DqJyEE3qtK2kM
+VvIBuKWQrQi0KGiifz0fQvOMxEja9HjZX7B3WrkmBcTHtrRlNzf9oEYLEkBUStU
M+dq/6T+Nbg4wF6xY7i+igSHYt6oGuytf9jQJVB4eBnn7d7RRVHdakfxccsnWvKk
yepNKDVcbyG+FtiThM98qbb9VXKXit63iqnmEbYi+Bx3KhyMZcrnlbCx5QlIWqsd
bGjLDVUBH1Vcyi7gqk4ZARR12WV98xL9fJieITmKF7FzukUCi4K9T70bKobQoLos
C5xSOjmfncco+egHkbngESrXajJZBHjtBqYhilbRpp63Q98xf2NYMtwuAeXdxmVB
Kx+w3tioOHOZUinP93KBnQTkUbWZOv1yrOfFA73LW+iEsyOXMnpkBuJD/PKJftr4
F42ggEboyUultkA88rKAHKwPLIpN6RDMCvOryqFwGoABbkhtmHv3kU65xBKunhQw
fQ1eh50VNW+AT1CukdRLBVdpw27kyyAfkOMBGOmU0lSOD5tMHnlnDkM5fG+Bij2s
J7SamduQ4GZlusMXZIRSk1g8szZI8EeOWniwx8RB3BE5ifLyzhVMeoXdfT5Q2txU
iB7gX5u733gnN9vnwSBVnETdsdRBZp20hSuALLmcDkOtvuNQKQSiMgsNjC5wvFXS
H5GWxOx8IKAUbYsjahm1iFssZOi/XNhiz4FUO79LqNAZg0RsLEJJ8dPK3MuPzcNJ
DGHbTutE0Up92kJ7UR95LNBQstrzIftHdlJZzwYaeX7Bqc5k0alDWU6IzJHYQuHO
VNuxAtxl3d/V4Hx7VY0ZVm9A1RB53E+ne0PODTUWdZv8daRkWjWprcZXAyATetXN
gnYqEZWZqRUFp9051DXzoDGzRnSKeEEOTIHR0L+GW2wqfcbldEY/4JlluZEAHxKx
L4t/JZ6fTU5YMcHSLK7Av39blMiw4Y000m5O9gKdBRtsha2Kj24lg4gxz2apqMv1
twmhPZFw25XzDdeOg/3yYeDkbq/GhHMskuY7YT2heua+qojQJrUesBk/K6/42Ft9
2POlye84bYAzhBbEmxK9rGZW/cfYR06Eb2iQEkoDiu5B7KY4f1o0xQ6NKlwLvXMo
IlLXrcPz4LS6euALdSXNslnKNkd5IstFj+eMzaJBbXYZ4L8YI9O7ih/AULPH25az
hLGSOV8EfzNB0mgnVW2EesQCKXjOQbqd2bJVxp6Fkxnl6p64OMYlEniFXKWAmTXp
kBEkdVrZDhCfaU4/z7q3jy5XBiYmE7n1IDtPE4DgE2S1RrYjafPzd/WW6uCdWigU
sQ16LJTG0OofV599YOvNTbdx0N6H/q7mpO2GX9PrZPfN4hfT4tkuqk+lV+odDgQF
dj/Hub02Xx+HMLhb0ZPdp+7BkLPCbglaLDurzZlFTBfhs/Ayf46RYjQNpSiv/OHN
YOB9Jl8a6RWyi2ghJFwk1mRUyUqR2T1/bd8s1GVeLcUipGmHB9Ka0JLsyQm6lLwX
POpJ92x3aY+j86w5Vln50pyy2ToQnz66x9I25w2Ugo6L/3tHtcKMFOtJou1rL5dt
Oh8TWEACeKiaHtdsxrq3RS0kB9UIQfhkhzIqdiX4SpxIEaZv6bViHDLZpJhmVtYU
epuBlOT1jSyZhdgrTnCx6IaBpGWVekzKusX/v/czs6bzdCiBAJaAzINng4IPluP6
+KE1rWa0n45S75HpSNyDxYKo/QSb9M/8yrX5ttitpxX9OOkQEF5aiW6iSm0pyAWQ
pClv6oSig/J5cqw1VwJtbS2UcxbXHo9/rdHtg8OASXYnL7OZOf2Pca2TPgppfXW4
ba4Hd/JzAgcOPP1hEjBLLY9Ucg2su3rkfkiSs32+VoHp4feY+fc20C2A/6rwA0NI
+ihjXvBUT8LOVlpebr59zTZBxNw3NN7q/L5pY2WrHGUSzo2owwMqOGY/F3BGQ/LX
jU22CC/z7O9aMl2FAC063eM27/jZgG/NqqxgaLPVW+D6pAKHR4Oks0lF61YkggC6
hWN6txknhMjir3QvHPhqK0LlQTgfRl56p/cNoGI8DD8otTViwesDJ/cJYBWYGLIl
OQwIJQ9WyUVDkFi/3hoV/lVC9UjpcJ7+eZW1oFzOeZXJUXBEpr1A9bWil0/86COd
D8k7tNMPmWUgpEZPF2P9hB29R/4lQ0FVxViTur2bNvYbOemQ59RDyPY4UQeAmE+O
Dt8g4Wqebj8m374C3zDZpnc+OV8RpDHxAT3P33WmGSY+LvlnfcZuNS/Il8yzzDvq
ZR406Ui0GVNLJKbrBV2wPEDUzeHZkL528ofMBh+6XYNkEeYTr7v91UAkGJcIc04n
3GBMCXw7dpozQtPW4IDZ4axH5esJhY9omISfUwDRu5FmCROSZzx/yGyp8GHKZqUC
aUwpkZszV91I49fBUAsbH3H3tgfhB7o1QlI/HEA0Y8LyTDCC8ectZEhfhGxgGGuC
9oxe8v6cH0cddISDFzIJaWx0DjAxxfLhUuE3pDOvy5eRwejIn7vB4Lh79fIU9bmt
c+na7LCURlWgn70g9o2X1GWt18N1JIl6MV5nYRFfCzwvs0ZhYlNhJl3RPOkSvzc/
P5n4/py+FJWZAMLDCfzZDUNuHaK4yhf24qQ++RjaMEypI18zj3D63+q6Ce+ClGoP
tX/RZzT2i+FAkX7A72/DOK5BWrvDupLTFVhP5zEIHUDegRXT0x5MxEek6BjxdP4a
ezGmBtsUuhyOeL0mnToF4UHFMa33Q6s76Q8e+dr0Ic61VkOy60P1pje/5gT/LORf
Fykd9KcIpFzTinZyWKgHjko+FLaoKpwfq2WnG0uTI6fgz32iisFckW+IiqclArga
Dttyv3Ujl7Zu9bi0watIhNZ9upUqxKu5xzJz6RtXUR9VjKYyXe4Yq+uTYL6qIx/d
y+343SOLalu7e6qkYxaI+u5wxLpn9GP4NqiArCQR9ZkvHiG1NQxmZxMCspEFisQt
ivJ1TSl2h6Jf3XvNKle3YUPEU1Apq7Pg7doWxm14et4wqzLWbiP3vz/wK+L+EH+e
/lVt5pjaC4hvM1cqq/npB8/UiWQy8RIMkmjPwv23OGNmq3qndT4pvmbyoQg343nI
Dfu/wd7TsYLPp2lYadz2HKZcYLyuaswSI4jWM7t6TQN6jG2ASMTypiWcQoYTS4cF
YDb6ZC8Jl8XzA+b0CjW7CDLYF64MTtNbfdG724TynFBMWE34gTK2zFJnimKkZkcv
TiG7ZAJKF9ayCJAVqOW3MV+N3wJazV50OshELk2sBizXfLCLqKKw9ihyABt3kwfo
RZnoqP/bp6wI0aRZn8HD2+rlbGYVwYBGCIi+f6u4q2UvijzFJur5C0X3Gg2fR1k4
LsILKZg9tIOjBYNhxHRVwj7ppXpvKk8+j9vWDt7KT4VPXaL22oglV8dyhde45otW
2x7D2xrjzSxQS/cKypyqCR4fO5LZbVkKOReAlqKwEfbi2y5gTTJNqI8nphFqQ5T4
Sa8oHYbbX2F25yBlFQkjhpcJAehA3lONPZf7PMe3iJ+xF0XBGzNB2LVo39Dl6aEq
1LNWbLMlMX5vq+aSaLhH8HSPS1eDvMx6bkfrFT1anIOQpD+soNDPr3SZeslGFZsa
uBbk1RfOecX0d+CxuX8ZuRt46F2kJXznNR+3kVU82Bvx7KGduCPKM6UfWgTw8H3j
htSXocLHaKXVtUapcSLmPMV83sNvc2ENutuKSZjy48HqDAIJ2Fam0mJDcIBFj1Ko
eLWm5D/UpbQ3sZc+f5nVqP+Edu2xT0x3kyRdUyy6w3dhYAAQa1EqwYjwsKlukGDY
zn62FkftYDs/2WqAt9kXD4XAImmKS/bVPVp1WjAneDNKDyHW+UEAFDennX83WvtV
LC+mHfNkbqM21IIpayydkhyJ/F+cauBpoNWsT27nyPM93Ov6h+eAcCIddPUNuav/
xO52JZqBXgMoQ9opRuovJKE0Y71zaqMXlmDvlvfLwVaE7t6dQooXedCFEZdRDLiv
XuhgGOtnhqeDT1TAxacuFfawKubxm/TfPCw/9g56T7VkzvIIHyhKABXyWU/F0T8U
fzoU7e39xr+aw6h2FB1t6l1hSWi1tEk6gVcfHK359MDGjN2Z1Of2MpYZuF9bzF3c
VpGZiCB+7BVaCwqX2ji7Olq+uPODGiGr8abXGyDXcSmy/oVcVioiHToFESvTH4sa
btwTCOumA8LH1SoN017lZYbbfjKRra3W4/jdlW4s7hqkbOIA+oryq2syNyAyffFW
elOI+cvz6K/oQdczQxB1LBnZOOnT9jLa8DnmsB2zAICkaqDXFYzt2Yq/MUmkmhEW
JxGOnRu+ku3IT4DXyl/PgDnbXtiBvTnM0405LJ9ZkDHsxmCioeq/f9RPU+5XSMIK
SeHl+7K7y7Yf6BkIliDqgDBb4t2rtKK4FMUyhe5psRe3EjGwDpURTU3HJdQf4c8X
svdmAuXw/FSqT3vnqqRpXWUjp60PtDYQb+U1+pUHtfjA84eQy9jS1ShDKRj//+fC
q4cSwdqPSARCLWmtnt1JfHk3JycyMpcSnj/PyqRCWOHNxQXz35rjdYEt91jWii7G
wunRwIiOC9sbkquoCTfKgXOtfzGCCXsEBjqXNrKAHF06L8wwdfMcjNR++IBK6Inw
bBt9BdAD033ZyZEImIUYtKP4geXb+mBnoA+wmKQmWEf1BxdLazfMAcrgtOG6s6de
ayUj6zxVcgBQDbAVo0ui9MXIJLgE9XggJ3MQ3eDl06szALeMDrOpcPe3nVlC8BE/
c0/Fm8dzsTw7MXQYKDaPl9rnUxE4iQsitH6h1vgytaI9ySm3Wk4B/JKPfwrFqUfJ
rsGqenRQMq9z303ojNudUeyb/uswbyFabq+In6k3REGolC3pHuH29+DPVT/Qeaot
uvVBooEYI2YRSTHmHRgeoZihpYroezCdFJ5RcnStD49L59p2C2O+9Ke9aAmPQTpy
dKUGSzn/W3QWAbgdMuAA9zThuA8GB4OUDee/hQCEzM4FtKyLel2cDAB9lVtWKW56
945PfRJQu6WCLh+8LIN3UFWlkfyO0bWfgrxL5zgoDI6WCySOoeDBdVWgflzp051Z
dtusIFnFpk/6qxwWhf161ee8X9FgBxi2bOZVU/3Q03joF5qcG9orxlepodB085Th
OgelqCWgNocJXUa+bAdjtRlDEVQ01c2Eeb8Tyd7g7YochpsFFWVV5+eYR6CSk8i3
We0WOqu6cUijk478R+30mhf5kZfiBHbKw8LLdIm+R2DkQYQ+mfrsP7Q0eIMeeeTv
zehOQLPyRwt3HHbW9T+h7vVvdt60gd3dXJhqbqk17HehQy5fVCHZolAjsZauItAK
UcPcJ+GIFidHcsLnwz8K6WSqP1JRvZS9zI9LpXDtyjsmkyV8ynRJvssTTPFW8BZJ
bOthqAFbfeSIIItWA6ZzVOo6rVzKviHp8tt8btusQnBbkH0UWGC7R6WUjHMkask6
0327/q6p23QzFhq2NdQvpwKjIxkMmuTf0uiNLjYg7iqqBBGSy0HAvfl+XXDFW4Cn
L0YuSavtBww/n8mb0F3b6PgV1fYjkTW/QnJIDfk4I0wKQI67UNfLs0DReZat3vZS
i4kgaLx2/l7cfZKm66X3sTrUavzWFX296R/iFe3fLQ31jEV3VbvdDzguVYaF4BOl
nFgBJuKXlUNjn/Afsm4qWE2fYhOAO2CGtHulbSN3vf30VwLrHkvYj/pBgNtj9Ev3
QkX1bzhzukUpcGaGWMH6ANaRLaeWo82CXVuesveO3gnWTqiDKPjljLMHMsRW/um5
TIm7P/WXPJ3eeSFe4dGipQs3s8OuPnUK50MFOCTFEj4k+waBVt0ClanKzdR0KjUY
cD/1ih9C8fUcGZEkOqD+bpAF/SG0B/0xxsyc6Wg7IkPvLLsF155Y/SG84dTQr1o8
1AmAr+LRmo77Gc6pJ/N5nTFMXx+GsaV3rS99QRyufW8a7DJIgdzFBGBxXecT8mf4
G9Tpl6UkhS8JEmT4VVS5NWRHha2p7V8JyyuMaxRy0ZL9RzDj/ExdFEoR04QsIFGD
LwfyiAxUAUieKGWrCwciybpl+qwAYkJ0On0ftCNuUoR9p4qDgY9QYQl55WkCkMXG
PQxI+w/Yjom6m7KIDoTcjAj9Z+0D3gOh1bUrTAtXEhVsEZAfM5PiZ2rchQ1cGwnL
WUKbyAd9LyuOyyqb1c3RuhWjNMPj2l6tT/IG7M1QOhbcXt552CHfr+QGVMu+TWVg
sGkpk+NzAhzr+R6bGg8ydbRCdOD6MPYO+snN79EE01SCzMM2OIEhSowiVEYt16Hm
sMbSmQFE1Z3LYt+lPcwSQ4kGaoGsOdHyxIgQsNpEpQmQVcFFD9atCTz2xvu57/j/
5Gfap+8YHRaSIN/9dzMMAK9OTjqqeBgDFUmkefSp6qyzObkgGlaOdeuDEiwdfuF2
HJ8ijbyPHWeCj++7OQiA4JF9tHDcjdGu/wTlXM/hfJNhUDFZzLbDloo0xFYh8lGh
FpsH3f6eqE5JD08jpBpWkjTxVrN4V2kfr/znReG1N6xKhpm7mUH617Vgb4IOIZYJ
oaDndNb9NE2wEd0YTm360epw0g7RYxBGccYLv8mvwVWU6Sv9W66w66rTOkp59g0J
dP8fWGDmqnhULvuVasXng3ASJgU8yw1Ewhf8VwOwSx/PTeyCLR9AclH5xtPCdpQd
o/FnemtTkjMgeB7LlTcBunoRUiW6u00Bdxmvcr18RJdxSDg2HKhSjWysKwwcLhk3
NtPMv1tJwAdJFDLKKr2FFu60HuyOR8XY378kOe9zaN4UzwKJIoCqXHUj1cSRQmZ3
WVO+F6fbCVph/i/hap8RoxcOhNqTh74H9ihFU3xt1DNol7A9A6yO3QMo3Y2aVAFT
/lwU9azp3LETK22Log8ZrS6Knj9UXWe9ogEBmq1g2p4SHcm+Pi4za1c/17XyS4iL
wGOz68Hh/JyTX4OOgctezbJbrr5r3k668CFRFwARBezIJobuMGSF7J6mX95690/0
E0LEeJ1moR4GrJ1VMiwCyCa9QyfSS70dHrkSui4x23tg2kqxz6ak7e/dfZ0RnMBr
yt2/kjjKd2eSUTQEEXb7DcXl34xXtmqZdj4ldOiV8gt0bG/igQvE+W6SokAGb5pR
5he00qYus3Qw1Y0O3R1i3HWlLvyWvJlX+QhELblKaPQsAt36zu2i1W9cmIQKaqv6
4npN5+AVF2RrA4uE4hVolzW/44OkvNac0aORewM5zQ7iC1rCH76qdWCC6RA8BmKH
navI/afGfKKGYCRsbcSQbeiUyvRWVbDvIjJY4BdfFt4wiAHsnL9gmhmC/2GCPYNP
8cvc19aVc6YG2iQmeV/fjaHCNsh2Te49j75VKYI/o0uMFQbLXcX76LMH7nVPjOXH
3n5N5j5FGeZDNnYdrDC+Ac8Tk2yWeIJq0Gglix4htsSxZnXsD/gVqk359yng6u9K
ftRZk86KBIuvxSQu1/bOvgzjJQixeIoSak2sNFC/E7zOfqmHzn63pvTZwWPT0gup
hIjHd6dtC5x+etG0eEm8Sr5wj+GtF6xxpeZAMH1PxMkwIQ7Ed3LvQG463l/fhfxt
3EbPsQK5JR+8ZOOuCEhDUjNBYIsHQd8esDnn1B/uTjYzWlY5u5ESC2SN8PTIrxHJ
SXqe0XRk7gHOPqSstkRUJv9fwu843EbPaKQ8Q+Bexu62B8B43OGfpcX87C/L2Hgg
BEzGvpr8w9lwzLS/NZxQKCjSntRsefU3o+WdahqBo3Y7zHXqu7OnAZjBnB+vX5+1
5Rf45oTMDjXv/meNfXQRQg+xEuDpL9XJVB5iCMXBf/a0QzWyhsQESeR7sCqUH/ym
oS1LllmsDczaq2EbMfbM363PhVxH+O81yKYTpUHrApSGs18J5/wqu5BNBLxrnHpA
nO+XyLFummbK5jTxX5aFWWNe4LhbFQdTqMHoNIGzTdFh8/vo2eYiT4KnGjC1yv03
s+q0+FcdEc0GNZa7xHyUnUNvlllCLeJajmHp28jTq3BUh+3vWea8NSiO7TbppQzM
THOHU3/yaW6tB6sVK5yqMhvXs7x9/qDXBRH+wEssIyDH3vpHzD3arCqmqT3IeTIO
Wf4YFL249Lzu2yKBgzZwhr73Po2RZ3aBDCwEflKJbkduTdKs/4nTrW5cK+HEbNTG
UMQ2uFNPt2/7LRUizXKzoSo7uQT9kE7OpxEh40Q9Gm0meJQh8vjp9vmgjZ4FBvfl
iKG/9QuhFPqvheaU+ngvYW90PsWXEBLzIkBF1YscVY0jcDIiR43rw0ZyqwqE2r8B
CUzeEo7j6nv2WPZ6S9MmjErgIHPN08N0gF/XIXqMByJH96Bt2und/lY9e1M0s3Ql
stfCnurSHPh/9YAeVg5xL9HEGT6ImZ3+FxON4fL5LCp5xVnKngS1RlI6a8gkhRWy
KCUwf3eNSMAYn04NNuAti13p0lwCYSvHdwvcg0eqKwmjKe14O+skZNqLB3Z6gCCI
my2ON15i1gj+gpnZnmHMfueTv4itvpB27HDQqVo+cQl6CJPao+PbeX6kDu1k86QC
jn5CLSqmWSdDrtDSny6kfkYVE3DeahOWhG9igPZVw2E2wopBzCZK9RbL7eAc8eGg
qKTTk5n6NgVpnxkdxacnX6G/sUUmkxMWZHENJXxl+xOidvicO5XpJHNUalFbDz2n
G1NrQC+9fbh0hiUBdgZBTzkbGGkfp3woZkEj5grqly3Hr8kFd4PsVBbakho7LjB6
Blr1TJMMLNJNj+yqhBU6cfK9JLmZzELwlSIlDoIAW63JY7J99bwsVJZgEt9EjQNO
u6z012HcgZ2qTuDlU20W5h2b60Kv5whcL5OCakBsRTu2NrHdNSm1En67Eltv11wD
3w6T6/D4+Slqy9inb06rAdwmqLICghcZF3khNQGcdYgT8J7WztG6laTDo26iHbsn
VrCtUwhez04HHy19jU+USZTirgAavfmGYLwY7Z/SJqnaHij9WosUblWnmo1T54BV
IBHfcZ9awVNVYYQJwTQAym3BADuuknZVc4fickkLBxB9YOAXhkOYjJ/JD8njEfDd
IlzjgSfVzXghKDH+EwYofxvsAHjzN0tweWrPhZK9qZ7arBF18HpQ+xJaDxIy0TO+
Gnn64bW6CJ6q4s0cg4Ob62QeH3Oa8LHRSEejfMMq5Xm5LFx3t9hrCae7qZicmpxa
3ucxG8l7BKCXYyW77WOZUhvRo77Bq3FGGvDeLZez6hO41Z73uMinXzx9kP+P5fWo
6F8kv03PXSHbdK7x3h6umYdh7IX1l+NAEV5R+Sc7oLzlM6fc6YmrIvIRdmGyYlrH
20YzPypI7IaZSRfYRykY712KmK1GvkQcfobghljr1J4uFr4qLo3jFi4V8vVZWwgY
h3ZCKjMVbbHlGumDddWkqMIMXork015CEiRzf0aeEZOX2Qra7Uw78Qm5PbG0VET9
ybv16Rq707gVy9aYM3mJn4owu0kCLfgBkgpGOAXMabJEqVr04lqw0pijUDMvWvL+
LNosXLlj0lPEiMYRkFHu3ljb/nBLzmpsNJpcgnMToPNM4dm2lcr/jBo5Ov7S+0q1
agIaQEo01gh67PfeqrOBTUhd9VcN4VvlOgTRo+NT7ohwKwADnRdljMhED8gfRQ1O
SoPHOrB2Ds8yTQl425sapxBJTru3QmYOLEj6JPunxrYeF+B5QEIHNVIjQWxBSdz3
jtmMrvBjBatfI+mCm/kkyPGDJZgQ6C2jvyp4tLrWQc296S91bf8mIK3kN/ccHWky
QdDcEUXt/yfrlgtxvXJaJmC68B3bTolwzGOtgpzQHj8XMAfOe7hpdljDh8mgfreY
x7itNOk1ENAM27P2vGUqk21wVp+4P6AqQAN1v7VHFl8O1RDifxHkRNTQbBDgko5r
AwTxvZXYDnfWXWGS5nWAkS1nf5VfTDM4A6AU8hNWdSE7UlUGJLTWuUZinx+QgG8f
QpB++1X7eUipenBUiSA7D3NDR3hK9k27cOSMZ9SN1kcXub/vIaiAqLfjru39V902
8iL6LWIcSmpxjafkUjOyDMvJ+fuPiIV1Bxl3qiUdXgW3REYlHNyltHLz0WkKcDH9
fpBt9S39fJC/t5mMANkgGBLZ6y5LyqP2lU/43QGV2lBTFZUsN7+oOjiRasfHH6H8
UgD6qYjGcud3kBL6EXDwQUOtWsGs5mEJHj5VuOm3TaTFZyurhp6tUpsqrZOVdyCE
Ldzettzpa+6RmdgGpX0Yu+REElTVQ6q74xyHOnPnX8rz+xkvrCTtS3FfZPPk87He
6KUAsm6hUpjqxHbzDcTVCMxT0EzxMfbdZw36pQspBDulUmQ3vE7vEbb2ubP6j4vY
YmHGm2VhLniHNsxdd7sfHFPFvSQbwZRLv5zWVK5dIvGUt67I+y5lfuTGGT27y/an
0qN60+dZfRoX3o79oCrwVreo2kv0gmpG3T75WkK8eD4DGbZ/jTcvJO5bER2aqVn2
jiJKTqN6uXPJ3Hlb2Mo4PFjOng9cOJ5ionVX9mJ+x6ePswo066wd/3/FsN2Go5Nf
HLjMW9ovDgGT6ty1r26TwPhe3yqof6xTp3UuxlAOiX+QOs/76bzJniUDm/lSqBmg
C+J5372HeCxojPejDYI6Tj14fCUxJ19JmfKLzyM7PNBudqfDIKVhFhvWzfTzj1yz
mbS6R4ExZKvd/SotcRZAnp0CU1GbZrKcRFqBo3Kyt7Lv6Adg0X5J4GPj6kGuv8Fs
uQ2ke+5eYWUBS4BYAkUZDzNb7MGaIQus5igI8q//sjmCBsKuUV1d6vba698c7d9L
Y61FfW0tw1qsBKYJZydyUOmAN3LFwtG6yBa0KJ1rPuWiR4Sf0VZLI4gYx9zJgVia
pkpxJGtpZHw4p3Dta9rOdcD8NiEnc4tYhLxHFrntJRaSs2yWhjLzpLYFY76e5yFZ
hBdtQIzjNsa8tym6FVcxjtA4q2j+s4xn9p/uSpudU9QDSVY3ev2ctg+Hu56QcYpK
lIEm6TuUlGZGUIoQ2fg8Nq72JzL6Bk3Nmvxl6NiP+v0n1Q9kMDTqT/cf1WZFhYHi
NtGVEj8dU4a/DUKPYOCxVJf/CMPMEzJ+tglUCfu3VBBtkL7vYSgpddbMPp649kKx
vEbMSX/xGZ43iTfOeOl88RePby7pqudYe63rIHiH1aGzVqRJZLo5pHDmnFy6sND1
AO/ihAu7nsjT/Pg+PNieQTMbmnmnJiEbMuZqzyKoXUAwr34Tssi/Y9H3yqzeRZXx
VCVkc2GQQo+uDb64K6L/Lg60o7yVix/rK0iHAc+ZwqQ24kfKifMEmc/vAwg2SgsU
z2XngWRQoXCWs3NfGmYXsgcHz+vhlfesiogPa0UFceQXUdzcY0URweJWPSihljCA
q8IQapR+ZG2EcNhF490hd4dMs58fzF0h/VH0vUjNc8ygu3yFjZBCbVlodPaUUzHU
yL/mLftjaBD0O7PGyTL/basJLoTV6LIjhizp+HQIEr7QNwAc6LToop94VwbqZmNS
mNnCQa3t86i4VBlJvSNe80AS5qqs96H8XLgr2ARYt4VAMj45VJG3KNcrhzT//4fe
sM+TvfVSU5K+qOM6iJRZ/c9E46m8VgPlA4Ha8//hMg/BAlUavLqNBeuDRY8JJSY8
REayUCUFHa09arS0P2pm3S9WlG8mtvx/+evjspnlaNgBVkVl6BQjdy3h+xsSiycC
+a9rFxyEZPE+eoR7Y7h1levQhZ2Kpy2rBpFbdhr594SB4O8KIgj8X3Yd8YvQkj89
A/nNVRcXRPcwIMT7ssTiMXx7Oxk/lXiKoLx99UuFAdATXWqqmx5q+8XlaP8faOSo
p8itWHV2nJkFUavuOosJrtc81KvB2K441e7jidIA2/YozxRxQG1m/fKJ3sIFYLhT
8V1eVQuY0lOSyIaeXAE/+snNU/Z9B5cpV3fecIg9Vn/MpOo/R1oHbYicvOtWaWds
gpHAVZOjej2JfPKyAMV8ALlTHjK2eJI0rVPTMPuHl1+gN8ztNQx9CHXyosecERDS
+OTGuYJRDV7UugmIffWRxXpxHPM7pj29l/76DUD6JiO5iFxfRMDIAM3IZGkS5L6I
r/h9Coz1GwIk+UQR9a7raHcnQtMvf8e0Pi+wuL1evn0aZLHm9lr6IlF6ea4VQTxa
ZvUhzLVe/2lqFXMMNxy03a9EE/7c9Y8ZWR71kUigJlUFn5u+4ZR1M+2TJJEOgaTh
C83rceGStAcQbTkoeP2XR2GVRESb9IFmIhfFaqM4AzHAV6qRv8e9DG773YciYCF3
SCzG0EF9z7LLLG/jWuEGHuxKNI5wRbCg21PNNdSkSuFT46JBLx1QPy6jf0gHTB+c
i5M+YsbQqlcVzlNCbW4rOPAYZR23bMIdrZX2ZafyudMkyMCdnDF2piJF7bDWqkcb
BjlzlAw0WdUqgJ/6giNor3nnOefalPVQ6BXOYLoK7ws4QTJ8s6Og8lfCzDpQNZ1M
/GITxCebEz0QCvdKI4B29nGwYWiLZu6EJOA+/NA+7qmleTa6KJUZ7l0CP8hYFD4e
mbNQROH9wJ81++Uk6nzMQC9V33YwcReXRZsoHk8HYZDV4nk275Aa2r7Hv9ZRiw7H
TSXR06iUig4/KSpTYTu5uz9m/nsxmTBoYvuMf+cQD9RRygFpSd1cfQfNCTg8ynIJ
djlXWSfE4K9nqQO5fVJXVI7TTEUoZ3mLIhpXZuRjMlJjT0KUig7XtGcQ/IqE4uMG
89MdZxgnS8PPqQgyPXXYuPUvD6RdlnQ5UNOUdhm+BzGcvmicGWrc6thoZFPJZ4Yj
gn2EOc/KK2BQMbVnUGIt4E4nXTXCuxo8rLuosZ6YlAPFhJGg3N8Vkgn0CVAqJvyt
10kuy4y9IOSyitP6kYu9PCgFKYVsW/qYSmIa+8XxKM9/umxQbW3izjxCB7EsenQ2
z+j3w7ks/BXaPwMS4NA5/wh4tYkv+bh68hDJfeHxJP+Av/uoe+VLMVZoEQeosoOo
rZXx28XdbGWkOTwZ7p2LrezmFI1sptwjDInePGpvLHI7gfQVwlQqYVdWFP3Y8Pzq
2aRCPmS4Dw7Ip56ZEGamWz5fvSAr1oG8FuVbNvxwihe2+I12wAz729PAuAUNqEzp
XQP2b2E9JrFEbBA4PZ7CCKuld9b5lbP2iX9VynXUavkLF4s3nlc+/Z3uWYDbdppn
kqbtvNs/Ux2Vt4tnICxv78IeOnZxe10sp0UV47zQPhomVUOV6n81r1eag7kByriw
lbshr0vB4fWIsaYL2r/PDu2XCeyX19ThQOwzoK/FA1px5XoXLieEVO9QbE1dpaGn
aA41uTVnKLKCKBt+KuZJrVzf5ZBnUMxECG2xQ8W1yvsyNcVkTqJuYMv+vIYRWnKm
Nu71X9d7YUetYzm2BH4vrtekcM5Lvn5IKGDvpXK6GprWQpHlCdPeWfzqYLnUp2zv
VS2w6pntZd5fbYFh3TjWSfN3CrpiyCS0c5siFskmZXp6Y0zWEQkmt5CX0RO5AlsI
3/6ivp59WZiK5PzRgsJObdbAqfbaCVC16nNisGsvV/ATej3cE4TZevu8bCzAyu6C
y5vmSkZHzwWkSWuofzJvY+nD/Bhy/D0ycBREPmfND0ej+Wp/eLFvVhpo1V0TBzT8
XFUziVJAj++4zbwjPT80IwWIBWVfPtW8ct/DTsobxza4A1m/BjGGUb5qczG3QQlz
+AIsvHrZT7ZGCkAfP0tQbbCYlN7Iu2Ba+tqz0cDxKwinp3J+REGRVomhmGt2twcb
Ga96FxEeVfytX506hSsY4PwoUE+pw209FhZs2rlswSqwps5U1Ve59iQaKkN2t+gD
MVo7lFQYEytfzgj74Bdc7fwDu2Q5Jg9Lls5aL9wA8Ixt/omC0qKepA6C1Knbnq33
Ct+HQouWXaubC7FAKjgHX2uyE3pSvxuQUbpEkXi1ZPxOXorWl9tWsiNfIkINkv1R
70AQaW4OgRp/XCJbHl0opHz0Bh+e+6hJahyIrovgQKhSAFLo02BYEMjs7OGq0VUD
LT7dcJmtY9QOnWkAkOeH32HA9sCLlZ6+s3hFFk/BorDWJW2rjT95LuKCPbHYRi9d
c89XM8ZFLmiH4AuD/Ky0mYn1RCVMHmhet1ztG/ZrC7KXLpV6Ub5KlYEq/P+P9zuv
HE/lIWB8pR/WHEjXgjC3HZ9nRUQZlkwAugRDJpgfNMUEp4DQq7AM9ZWoGzLCMUOn
5XfO3+fBksHv+OsW50b2xoQtRkaSvnR9EogyHkpqkq8gpM3XaX4RTXdoKL0Lv2/Y
meaQUloaIufgM9K39Z9u5OpXKtwrO4P4e0hD8cE5Fp2IlqilZWi56seFexmwittc
HNRAEs4ftNNgGmCqzGyoxQLvsQb9+Sq7NxccZvzLabFdVs/hikQMUGyJ3Jsdr/tS
zxK81z8C36qe6+zMLxQxekCu5e/X5P2fBs6NWXsCiXyGa4hVfEOwHPbhiyczZpIG
V8j+amYdHtfY1PiWITuDlci0uCqPZKIdqwwF4dMffckmgwCnFePld45LRFllcduf
4kvfu7d+8y1yuLUJbS557ya9ONLvxiEZTJZIv55hVNJsGuS1CBnv14XYYBvhTxXG
OD3R/tbUoNadU1CfPW+Y7XyJX9bBCRTmLZbLMLSJyhg+lUZZcYHEtNfKH1FmsVQT
H9anfQdr1dBF07w97ze3ZyFCDNUtH+RcLGHzZtvL3icB/b4SpE476fGYY73Xvm5f
uJDupu8CqqOZmWfvsucHd6r3veR00gjAcRgaZ17b8ZfNtGKIpKVnulbBu6Ntb7KM
s+kkkawuq0a4oxGM8taGxQ1LuzUkzc7sDi5FqviFBq9SeFJM9TzM3j7BxDy8ef2i
35xGbrq3uYeiljlPlJpNKL7PT/XPYx4gstz+9ET8phXQIZMCL2XGU5CGNbtO4tnq
WGH00DcbNHcwxfqimInCDhPJbZY9i5Vcj+nbYMptYcHHJMAjjqxH4mzpN80c938f
mK9+ybeXoFG8BoP4NQkcVg9C7lgCQ/MI10Di1RALvZwrbpY9caRQpoJHDlrTK7IE
86vVqUlM2jcucwiLosBoG84xXqFCUAVSfgxa4PDHCdNlvEMguJDEq8B0nVonQXwZ
VYOalQwZ3KmZbDmOf+9lxujr2DHIc3tCyCZJSohEyNXkS01xWZ564aQ0nIeW25+R
q55bw8BKro/EoHczN+chrxzpoLAvlpeQY5bNUu3PiaOzLBcoN6tNnXkG5EP+wkKS
cCp6KEH/io0PWohuFQNGVUrS/S9TokePBOJ6xjU093FmooX88DHDjkrkHqB/ZkXU
6fFNQqQO9gX+6m5QcT04D6BeqGGPWR483ZOO+mB0zI18qHf5QiHN4vFWxunjtBWb
E9nc6y3scqgXIWjfMNU8ISA+wFba53e7ltW51vce1CXIOxjjCuWIF/qIe4C6DnSz
PHkLRzwctmwdgyDu3ikF8KXv7pAbJcCZmabDURcUj/w/08AGahpKIi/zQ75FOwir
PDLU1ZAXgxjBbYr/tdqVs6VEPZ0Jg3kwI/WmYLr/IBXjrkb1tEHL/6mTHM2vYuQH
Fvp0eR2AKkLZ3Pboo0nnW6P+9Mn4xOb51DleraTBCPkAfz0v0+qKNZp7pSO6gKRl
az0NG368H4kEkZ5lSKZXbjMWi7oBBE6+qBiuPkBg/QKtsIE+8HUw00UXFk1QYuQc
PfAt3qdLwa7PCOK2IT1xuFQy1kIJLTN0SB8lxfgpyWP1BcsVv2pa6zyKEmVctDLl
g1PPXVmAJAX7gLnEDWVkTbV6W/NK7Zen1Z4vDbP65lpzVmJE3GSC1eCGOp6Yiplm
jzkLpPlivys0VnmuAkanpV90MxHoDdnnGdkjptzem/tDdCN0ff1XSLN5d0zcCh+T
HUZw7UpJ0y9D066g53xj18AfTQcls1r1gRHzlL6rnnXi70maknEJNvNyGA6GhHK8
XPQRJT0LRSLCyOiQ8w/g38bUjcVDfmBApD6Vkf4/IyPDZcihFW0GkPtCMUbAjXej
kIzB++JsEu17nlpHLOacR4SGR/V6wZrOj2VaQUvOdRsGL3zoSk3189u5t/aYqMEA
vvlc01L8G1JfK0HFiGvjTRTV4szQK6Fg57gBVpoZ+l9SpZo4ZFhvrXv6SA+mwAUC
tUxvLpf4m4nAdrcAceSzejVseQJ8jSghJ7jMHFAAN939c4ivdj99KmSj/H2Whzst
HJkjwgN8rlCNSYzckN1i/+cMARu1JJN9SrpksllRjGgU64SCPcvR+KKE8uHWGnIT
h9nXRv92GG+nWOGDvJj+soJuir2doH5m/FJao8KVbr/Ba4ZCFgOJ/dGug4Mbabnu
qRPsQAJYs8xpRF+e34imwlKx7+Y6SQ5scqGJzk7etGjwNJVB1sThcaBzDSoe4Ri9
93JegfkR+YyuoNpY6BKVm5tdc8l4+dinQ5PFobdYyACYaMerr6hGfsWOWQWcHLa9
1Q+W5vNSEqx3KtW+7KZ4KKfHVO5VSmLb4Mg4pX5AQItrKv/UUi7Joy9JBiu1sy4L
rMsNA5rx9uq6d4gintmD3kA2WCVYdN8JIqoOCPQhh9MZnXRQonBt4fefCEqZmop3
BD0mYEKywHs3+VaxDjP/PE9W7D9G1aemuX1mFCzGWn3ZZAuDJHfoeDYITslYzRkN
BlAYKtV85Bd2HFWa4MTNcxEQZeRl8cFPzgfAIxDPR4+LqyKpVrgipCcp/xFAWSqu
a5RS6x/EAa0P2zSmUnW7911lvHQzUgTp+Ml9uIh9GGIq+5Xic4VjJUCNBwpG1zUY
UzjKu5YfoyLY1Fvi2vs+kDfJvMTyCtJuAX9/3spdjDeGQhGJLPtfWZXK3tqI9flt
4SCoowxeHjV8Sqn3Nqkt+3HWgqCNsaNIgU0QRGVGz3tJb8iPysb0hb0I4RgOVUxr
UN9hbEW2VmPMgkiSLp8wE+jF9shAmjZAZzYQI9O/2LkgRzsiPZECY5WgyKi1p9D0
6AyJdPh9RgHn/ecWnSop9rSfXoWYwdgOSztGEkIJPV0splw9MsBbZym/gcpZHpwm
LmKVzdLg3zPdtYvOOdkXOJR5485y6ijX9H4OUPB4aLLYkzMYuhT+tjW//k4sBpb1
iNBCKMAjas508Wehtk/8q+4VQwm5GSxF1bsDXfd7F6d9JE8cfGuBa4jRQPX3tUHC
W12S84hyGOzAfSE/SrJVGsMlHp6+hVUaqcyz3BjNbDxpDcNDXTb6K0PPdn5iKr0x
SNaU2uP6oNv8RADCjJSoK2B2aO8m8Hrz2g0bnpBS2ZbnUFflO6M9lSmF+nVMtTUY
+g9hhBaRYDGznIA3bU+0JeLpy1bpZ9/PuvvoOKye5H2y90q+cbpEk+KPNoS4XzNf
NN9lwHmMo0Ncm5JdaMi28DkplMxF+QZY1liAeCJVW17O4677VoSSkRJwi0HDDxmI
1Mqou4Jv4kZXHkrai/rlghrDh0LZ6vaZ1EPkheUoDP7JcDcBouqPC8VjfZ/JKeLw
wXcD9AsLhcsGZer2aWyRmA0buuquuJGjbCzZdjVDbh86Jp68jbEx/rX6vN4Bo94c
ZxwWLXEhNfiIDfMVtDTY/xZWij4NmJV3No0E4rdu0FkSLP2056ANDFkmhIbnReAX
eln81kIXhXuRwUBtXHcnirurOh15icayAo4fBetRqVqaqhnzQ08BTdiun/vZpv6R
FZdhyC3MIyOIanXkLo1HXgTgxRTcF73ARZCaEvcojVFYMZOQjI5pS7m2iFOY65kJ
faPp/onouMp+aXsU9y3WW5Pvc2tSxAa1mGSKbdSBVwR+oues2+HyRaRT59DH5SbK
eeX5h+GwNILDfY2cK0mIAIKc2c598mDYJ1LqT20J04izMMiIUwLfVHH+HMdjMJfN
2wyPMo2WtZzANKNVMISgQ1Cm+lqWWt6GqHWoj9I9dByA+xdXKD9M+goG/LwYKTjZ
93WjxNkcvIyECCZNMPXyWFpc8DsJXU/VWTDEfuDBR8tO8VAURR5PRhhhmdCc58yk
uooOqPgycZCIQ8YVYPCCbwSiYS1LcXfRFpTIs9YCemF27+pKZxcl0QG7X1JmgiFD
0CFeBpW1dyF98wGwdr8fn4i0eRM/AEpgzULBqrF0JbCiJDveh/n0lC+KA9lLDJtp
e9b3l5//NNiWfHXqQHn2tJR9kqRhZqtefZMKBqNtuANAXZdd2a4vV2Yl5j99+aJP
BAR8dPXW1FvyysJfnED0UYyBovuPt/IxZ7ciwSQuVlvoQ59/Vo+A46CA12ptLXI+
q29pUtofHsPfjzhMqhl3w35gBUC0fc+D4rMzyPuEIdMSKWrsMr52GyNGNVlXpS49
ZbjuKHfKToX5qZN7svo+EA4e6t3gSYFElzanURAzIy2V19f+PNiSOyUiyYg+BtTP
ndmNmhU408+EI0OL/g+HH1j8UdBWxISJDrKRCFBL0OwIiKRos9IA0NN26F17Vcrn
inQ5aRwvp1yzZrmUEVyBbh29uzHw4JqVCZxzsLMncHcksMan0K5X4vbV9S6mCKOd
vc3DPkgqz2izzXkgN8PLIlxNe74xN0JGjPJa5Am+Tejf3eyDfsXK9BnPUwAKuW3t
y/VyDI4yIyAnCAl5Cv+b8mSdi1+2L7kxajkZY9ccGSBNes30YflULZbdQ4eAa2wb
HrqcSsBPRi3k2BY0v/JvCi2UVc6DwjrWzd2lAb4CjhqcTeD/HTKfl7v0o/HYW+jS
8gi1PNkUGD3jP6cflTkd7Jvz6f5d22i+fPJKpS+QUvVXSxOrX3q++S8eyEAl9V3K
78RmphHD3W9EQHUZZZYVFOTug7eLvpNyx9dJRSWX+/TWUt2mYJ2Vfufc9a1vXZhd
r3gpsSv3bRJK598wEDefakSWh6Nb5bEEMjjY0gmiT+7GWdcvMo/lDnQYB/IYIfiL
cGWGwi8QnVAEkkmFGgB9w+Zb5se3Kb+fH8VvGFGMhoMwVNeeku7mH0W6c8HUB87z
80jv1NAlkh2cOai1Lt9bVPH/JXYt36PvEJGGuwDqGE+l33xto3Sb3eP6QaHCeD2K
SJ3swJoK5ErBXU4FzryloUM0ns9jAC4vBpXTUQaW7AGF5vPPYZqBUZeMTKeQEHdc
t1pgfJMZA4bsQJHwA6ekGhr6yyoKwFwFuychpMRkryrV332vkGMi+Y7v9NYXUjJA
3ebMB+m2qSckAhH/vLPXF5CVgJ1y0l+utNjdrufiFhX/CXDitf+zXn2TULMXtC3e
CMvTWqIcVIDhy+6DrAfS1B5TGaCmFLvmEIfQMgJA6yHUJXCMPb4xHs7FCzNvG3s9
gsqqY9WkEeuz5rJ9xKTrKIDTn75LiQtBxynWCYtQO1Hl1R+AsRNecbzFM1jlTgd9
dd8Ya9u43nDMLcDQ6S57P3vGLwxmWKSNUoGYAJZI1WPqHvO9Po+kj5YBfmMvSHss
55+sjrmTVAHZeO4o6iXNkJWTdwFyOui2Famg5MJlizMeqxDxTD1QSOkgxkYSCtG8
5Wxx4tmOtt60Yksk+TEniiqhj2pMPUeDuYHaWrSDhj4D9S3/4v+F2AcHojt6ySSc
bduDhBy4WSFWVrDOBrLszalXHFNQ4N7mYwqNG7zHhdFKrwbRMwKm2B8/rnsVATAU
2d23ojMdc+sgcDar+doZE3nAYasbaT1HZRZ5yHwyNyNDyuRSTllvaEonetEw+E/x
eFIRLCx2UZrUHAyFbP6gBGYODwWDj0xbK3WZQG/6CVb+GDTQ2gbicCAd2uRJOXSY
azfsLmdY1qQpyG1eZy2PAzkt1xmLIOUs9hmMxXeXy+gj45YPr2zyyPb2DLVJzoPj
3mNBFMAOtuVJLKJgpLnAlcJbrsaiVVptm9QBnhj6lfTHm+DDU3nleK4VHg5Mky0a
C48hI45ZSvviT0pL4SNVUJu5+xrNiiGhDbJUYf4hMbfnJe2CZfTrmBulD7QEw7Pa
tGnl+e54/+CmwygGtTcxx66tquQCeS1RvsjlYjgpT+J/xzKGkQpYcxNq9W69qLiL
tG7s/JhLi8XN9FkwT0V184mhL7OZDE324iQnGoo2tV5dCMW54AVYK/kk+iBn/G0z
6HKD8QeCRBveufQX6kRuhuArozFWw4CPxsfh2MHSGvU8T9RXZauNVyXUt+rPMo+D
IAXvIdlSSKkrmSvwuO6xUT9MC+NLjnXaXrsSuiB0dl1yBoIDD8CsgcjzwgSqu1dt
pcJfEv4p1X2dT6mGmxp3vgUyA8rc+qN5EJhSuuun8Z3PY2yXX4YHsIEcIn9+NbFA
j7X8OKZGNq6czp++YCjFUeOxtbZM2I/TOl9lxfONL/STqlduWPtCGzeltQTx+B6s
WHG4tfEa4SYEfbMGB/frXPmGHHVe0fkCJN2KUMck9selfRbMiC3owjQiE1W6EDp7
nmi4kVhsTGS8GqcwUDhUMaOBnizulLtB0cXcnwBNpfGJbaIhTtP2JU+g5GagUrKQ
BngTWHy3cPPwfbQdUUh+xoCiPfdIgkglQMZTiCEXWZU5lVYjIwgSEKQ6GqodYBbF
4aVsHLY3gR91vBT5rbpyYk4Siyv8BvZxaEOXtkXcT+XekwW1t+LiLmgd1RIRjVWR
Py1atAQhG1JjQL9YSpaaotpklNgNO9N6ymkXPYl43sNd1AquNCV2LpVtqdLqJtMm
XAuk9kDUF9nR1DFj9Ku+qdykAx9VUtDQYo6X08fVfY42RUOkMNmrugY1X+4WtX4m
x8nkql4YcmD4biCytiPdYUtoFdHeZSzj7eb+PMZzX088Dfflduju5N/qxrwsAQhl
sKz4V2mmdHnT06fPHZvqmRUAk6mm+k49PzIkVD0+wF9WKcDnUjK5FEBRC53G07xt
xqItxcPe6i8HnF9gyp0sLnGml8Dmd+WwZh7chz6TPKEwUHJ+DkFyZr1ZJga70PSo
y1zxWVOOR3h/JcD/OAE5Kk0njLjHeiJYLsNbOpbd4p61k/RZ7xw9awJ2boq0KuMz
vprULxpo6nRCmj2dzvEY+uxnllelknequ7Z+dU0ojGMu7fwo9J7UMGu8gQnLkuoE
Yg4bv5FeBOibTbTZ2volJztqweC0Q7LbViXwy+1rCsE0acWx7/fcye+jrHzepXiI
Pw6bwYRkdWIBBYEvI6TW+Zf1gelwR3TNYmLjPdt7HyC2jO4xT8SMry3nmOdKkFEe
WHyk6g5cOnhXgYWF/UHbZVzSsBmni7SX8XH157B71QsL0hTll6AcgYwCQ7YyD0v0
yt+2vr/Cu3u8ZDS+ZHBa8Z+NBM+S5HhnMstLjhfrwayiqCQ90goB2Z0+uJYlNsPX
AJK3y04CrUJVQqnJ2d/Sw6/NvDr6T6cXWfODUqRb8qEZe7TUbeTIR9VaiPA9Jet7
/epYbR9gMlmGwL4GV+k3SRYKzrQiluIsSoNID8Gkfk44XLBsNMnL90sHsyss/NCN
gGg462s5Ht6LamNHWBzPXYFI58uDACT82zBy0rwyahQ9yfgRbkR83cIdjX5YRYlH
fvIuB475+WE11NsjCZR6bUDGvD6BPTqcSZ9EgLN9Lfm/DVcOBpxIlAyxJrCuu5U+
h3MrZzdinUBwSJ3/VwOlU5ex1+XKprVYVzGy5bMwChaDr8ZxcD8xy1iE3xlxhVsE
9AoxrTeO3jFMl2tU5Z7+AGtrsyLYzdkI1Ed0K/zqTMQrSxThGzCSs2fp8GC/E8KG
OkhxxXLtWU7HxaKjUU9gTstX9P4rfq+5JkAdNAm/IyvMISnhMsqLgacUJ/PXqBOx
qO/zRii/yj/hEILG1jeSph20hOLKCYMQHT4wEUqOr7A/g3TWM889ynDgcxQN5Z2R
kYhUEa7Cow1CuiQyLDY1fl4nO+7RG+Hfi0ipFUIQ3rTq3PmvESTui9R2Ld+ovWOi
6irrGTBDGr6U9PQC8C9IehtPxF/VLsUPPjncIJfcvp3w4F3I5paKXdVjlpOTEkfF
tiVP0PQmQx56K/ePVeGGlH5Xvq+7E0MLXp6hjyF0qfgdM23tFuuXc74xDQUKt8Ja
/nqU7U6ZNDnWQrddkBKW9C62QnD7IHAe2Qq0nfb6ZMy/SLe5xRoUNg3XesoFVNKx
BKEyWrqV/gnrNrkQtwxT5uGQ0Z4I11Eu6p/+8DW/pT8I77I0QT+sEOadH4iKr6EJ
VZ2ZUBF0lWyyhXl3bfKfrUs7atW3UnRSLsZ8jxRyJTbZ+qqcbg7VnmCBDH4N3+kP
EWwwLqPMMMBekz/tcirPGrQa75xci+hqOTX4IIjOjnXoyIXNXPs+VHxa7hv5E8B7
3MremJke24knxb9WiA0055gjfynZcYAFkzZxrxWd48dtHfMfTCpheGDr0hcrYIXb
4JaNr3LZrIvD3BQRi13q0uAjTVT1vrhDbE/EuinHmX2rVIiP6A95xXBS/FACq9at
1NqKXsg08enXE6we47FMpRqQ3xTWML81kpJfbV+sLbdLfb9bykYFdP6S+FNRZ8bh
0BFqGV+fm1TojxMQCUwmsDmtq9bXD/EjIEx+qycxuaPq2z7XEGb5I43JH8W5RTie
iHIIZI48CJFb/xFHosR2WPFfbBPKlY5SpzrJuC/9iqbBlFFTSh5z9AjvH0MO0SUg
lQ8Vm5psFbJEoZ0ql0+PSgmWDK78fMvOH2zhubg2luKKmAtw9/CNR+9Qnzo0+A1U
H5lhTe4v0Fzn6th+rJTUOZhKm5r/hngM2AcUdCwwf1fVCCymNBA+ZqtJroHhwhGU
dLBKtE1PaAIog0QobHvxR67bXA2V7YiSLRX1vxwMVCYxu+Oh0ZmTO0bDe7rcAG/4
/4taOxOL3jt2JYqJt/Mht9HqktYv8P9o7NWUH0oLhvqTsVuEYh8/SPeKGNvleI6b
vdyolhusyASH7KclvMPDVXMLmIjhBv5qDkB4kqRqZLgBZi+eP8vjEjFwWa9i58gP
X2SIeKWruBtsZ+HIZzgXircGzHQxJi4AgswFojr11LbHzJuBEFuaRXJH2ycIeVtr
O0XUPPcdNUG0ExMojmuLf7EyYXc44/nDdzZtiPuHeYwCSZe5wci0N0C4Gru7zgKz
u90gOu0HPaWiuez2kjwLBVdeoP4U6KxmdqYZxD1MN5gUk5q52y/4g+zgYihP9/Kz
7dTWuY3UIGpQ2Iatugc3DzyAIG/EJX1LRRblYnACoeOtU9rbU7IY+Jmh7lNYtohr
pvYDjhWYHO02HJluH1k0pBByrPcsuQrSeStOddxzLe5K73E7Fhc7XVMzuHSjE2+N
kYuN07OJsHanml6YeUKZ3lS3Jn9ciCo0CL88yzht+ZgBHapLhGvrH+RTVFiN3QOE
PB/czcvXrg/M4OGN62yZ5jY9RRjC40ICoAGjQCjkzvo7SPFc+8fHkaLReV9eXHmO
HTc0pa4qQUYEI85xnG1Q+tj/pC+1wmrEp3XQ2GvakXK9t5JgKPK145/KriEafvzK
NqlJHYWV3sRPGM9QokbbqnU2+/RmdRaC9L/I3rmjF1LQXEJhpFBXYmAJJvgQoMn6
drJQo22D7ir8VUruHZFN5PNQc85XrUCx/GVpcAy+DBj5P6hJAotomOABTAt27t8/
YCXJBBK/eU6ugfnWVx8A/2hvtE6uiFhlTo7Ylww0ckwsQX8Qx5FOTBz/7gQx7JdT
V6pdWv6tay13dz6R4gML/px2SFAVdtxXGrVs4ln0h2XGuTYZoh7kZKfLlwwpopcj
ecA3JE85wDn4i0FZ8Zd7KSCeY9/98S6YHWPTacQxpuMaQqDaDtLs4t1wco+jdjFW
1llSib0tR70OmD1pWHcwqtuQjXXnB4j+SY3i6mjORwVi3LaD5soSadXn5U4b3l9j
jspbyXUnaHqO74iU9MIxVuEL6dnQHO9LCv6qdczsImZ+y5lM7G+feS4fsjMA8Sph
du7LVpJSqxx5fwvq36OyT/KM0UUlyjfZ+Ch60EEKHtJCdAt0w4sO4qCAHFqNuCwY
QHez8NbriWbTcHjuB1XAfakQjUVxhLBlpGvEF2gz5M6k6/QbYE3amLZp8Cod78Vj
U60aLpHJzHs2i0RuyNqnbCO0RGYYrsdb20JnOt3cMPpdgPZ9LexqgKFXIq0U0tJ+
nxoec9xB7uUxlufy2K5sYMuQwiyA5NC2eptetmPKFuZLQiRZUOw4xPeySReqT4Ki
8g32nFEjH72ybCbhaB881K2cJvKXThtOcxvPyIy8P7c5PT0qNh5FexPWUJOr3F5j
wUe9J2AWxHCmJHwvUOuoCruXa/J7O+Mj/z6DmmcV4agTTgUSOsXsOID4egIOHT1R
KY6vpYJLg5gjMPtVlsXRWcMWxdQS3NKtuwAVc71Jt4HpNw8ju02gVmLS5ENFIASW
5j+bp1aeIjkyvzUat0NIicytpFqCQIXNCjVJGg1zE5FSAJsN5Gk0rtiGKOKsAVck
ezN7VfRxYDqGNsuFvRCfu6QbtISiYvYjDyCO5E2x3ZtG7Nw0qtlNdYKjrZaPTpWE
JbJNNoWZ+rleckvR+ADsrKe6VVb29P34gc6TU4hQCIINBEKastOY7eTX44Ev4Veh
DsUhfviXwESzozcYUUVL/wh1Pa1Z7vCO93qW/VennJPMk23ot2qD/w2eP21FyBdz
6e4f3Wb1tEot8JdqtklaCM0e84dsypX+EicFqPLq9vsQlp+4BKZ1dRWePzKoruxy
V2gr4QPSq+7WpRiUw4MdtYHxn3tTmA9DawaruR2eH7L46wMesG9CnXPBrCXFI0jZ
46KzqTTLjyU6qem0498oxSKJLNivJkfW0uEsfKKlgMMRWDZC3cveUD2dhynB4sW8
Xhs8wf4118peHPQ1VDiGVGRQ9bgZS1n1jJ1Urg6cioIuhmzQltGM7bvWzZISM8fv
Ex8F1mw8ePq9aoIsUBHy3EnQRwdeiogU64CCAC7StQyduRVz5Ay1qv4V41Lp/NfV
QKSydVkaHtGcDw4nvbT8t6xuEl0OK+VgSSqf2Is8pIeS3OGqT8t094vRMzdeFOq/
XqtS0x4IlQkIf0ZqDGxWBx9e0WXARUyrFv0Rr4YCalo8+JJSL8V6iHtOwzr0qbZk
BSAhrkYBXSEZSoG2ML4myLw0ToXLa13t5Djctv40kyvSQWvCx9m6wzTZ/ZZTBwUL
5rSClAN8Sf6DugJ/jiV+ujt2GhqEeORm8imO2yVMQ795XLl4LOR3qRp38mj0UBpm
9d5xNkg+5rvYnE56mmXh6eH8ZOJ/HWVLJsEHyxAvN5he6oOGC3ZIazOvgNoDdDN+
DeY/MDOxJ60TghjC+a+FoP5T4O0s5IRhK91e5Q5KBd3A1LTeApGNgwWgxVQAiDdN
dg936sZKt0/1kb6F7E2phyDfiE2PavTJwFOgxEH1XDSlnzqY9CarVf0htFWzvvIF
aql5ayy7Auw6ZVfs/1dMGExtjp4u0sQANe11wOzkf5dIeY28kSl/7NmcGnpnUKiK
7sVa0/gthUCJqvaecG1n61yHrkTnRm8OEuVsbXORmws52zMmO6tSzIhJQHCTYhQB
qln0kn7UNfw8AkIDraJfkyOV8TBRi4HMd0fzUBRVCNIDu5cMDuFr8t5re2eDJ6XN
s21WESDgDcVA7ycKVGu+7VfjpqTKWFiuHWZI5EPK7q4op0CJbeBDIxezyBXLK4A5
z+0TkDUE/ucwIsUUelinemlhmzCUzNhYsRy+1F2HeYqWQcedriQa8YrRRHSx+Kmr
qdovjNzf4O7EQK142FrWsZm4vCpovIlzhQMfRWmZYSwzzYJ5T8s3RSvivC/Qt6ZP
FYwQbDbD7k2r33Nya5YbqCBJo7O8Ca/vl502FH8y4K4YlvBgGtCbbXCXlPboixSx
VpHF/fqPyUAWopDv8v1ZMScqtDejLTQL4oMKD57ur2yXa/hCkDVdzef/ooyEd6Lx
OcFmh8QzB8rAhVf+z0bdG1EJwap5wR7t0nxzRSr1xSB0mt07W9lQFhZKpWtf4+Kj
QxZ9RK3omLzcw3pZ/y1EX+garfG8tHLgbY99Z1FB3aeltxqPzynkQQExpplGXljc
CYWRhZbtkDMrLdSrLZVpQovbQbEYaBTMKUDxJBPKm77IpS4i7uT3FBvkYEyd156Z
Cum5XjNtxNGRw8Cp91JaPsaXGJOfsMqkuKVwcmmbq+MWk5wAwA1YM302fqsBHs4r
XmAyPOdPt24cNLN3J0BZDSn2gfAQjusZO1tUKyZJuiQPDvmY3jZNWXoNziOPMm5B
7TIiPLzJPW+rVT42Zw1ZcsNlKyfAcMofMIKtA1tfrZCE9aRQEI4m+owVbnmR/oyu
tFIkIiHRzkOIRnakxvYRzWjS+pAagtoWbXg9suLDanSik5md4SV7IrBXNAM6u9B5
jUAK+pyD2YJOOYgKgto5ERVO+UIt7woEmaxQMhs7NgkdjC+CdlaUJb2QbXf+PVb9
0ov9bgppftBof6k6jBV/uuIjYN1gqoVi8tQPrZL2zfr9dav2slOypdMxnD/r2Wkq
e4pQBn6yJoETalcSXsSMCdEUtUMZtml9GJV4hY//GLzB8ewq15Wpe7Z0u9vJEoR8
n3Ja/sg/bYScYJBGzZRKNkHNaYROuHO2SAZOSwGxEXig98lpFaPrVF/jNYzxiU1T
/k2jXyP5PGB+kVhVhbrzegKcArJ3xLLvXwDrr7QR7AOEVs6xarjCwoID0TiVEA/F
3hO/TOs315SKrKY1QYwKMcShkY/wj6jndG/Xob8CQIOE8/R4AXoL1H2g4lHwz2h6
7kcw+Kqs4J2FKGNXv5upNw0laCfmE3jDnQwBoK7jflCevFq67fsW7y1cld2RsRbt
WUvygDqfA3+mAmAn+ojh5iVUvlN27glvwNiKVWZUS1j9QSr61HR9EOp8PQwhB2Gl
mGrQxyh8GYMzig/XvV+hxpY43QLstpIoIMrdR79xqcHAlCY4wJKciRzq7HzqJABc
eCQ8ubslLXjOb3GxdHpTWGSqT++fQ4nM9dKWqdUkMCNdy7LxmD3EiIztiEbC30K1
lAFaEmyTbH0a/5QMvZyFlBK2ktghu2Vdo12C/KJp0c9jQvgPgm1DuH1CY0AaH15n
C1Npc+SVnlDHHByLBgeYj7NfnX6F25pjn9rTNXpR07cEfXXbY8Dydmc58kPdTy4u
T559IiosktM8RBRi8ZGJsZw/gj4w9oC/51XuSDumsbb50p5Am8sSUHhoRcWxHMUt
erEUYUNry4w2hMBqok3w87YV+B9zvi8QT5omvsYLdrJ9V90LpszQWcu3RJZGiGIW
/Ks2BGDHSziDVCEL7Eb6tByDq3Hd6+99rgyHdQI21XpDGB1YBOq63j7/vSG5ynE2
fiSN6eKumvrxG9mqIcwgPmMyu0rnxAEeBk+lhlyuTUxVpELKN2SsHBYXhcWaDK5x
aM52CXcdn1C9Ue7RRWOboD18VE6TKkEUOmmCfrhHMWwkdNlu/Pnk9Bi3NljEpB9Q
GScpVWIYsF0NUhMRrndyWb6qW3ihHWw3t5zDOF1WYXlG5cDlFuaqRNAHSKjcP/0f
uS6NVil8zqhmmTRMUXpgrEBce9nkq52r7lb3/pTLgktaS9JnAjmUL3aEEAPFqQYX
jGrfm5haWIoWMOwDwNUAPJ+413SZI84BupNoUDr6t3uaSmH+pdeTwJmynBLY58J1
fPSTuORPY7P2s8S8Idc5HdPkSD4MgnKBNf+9XucNYbo7OhpzqtAiiS02ylKStAvd
qX07bov1FB080SL/Mx3s3ZJit4sYHUW6Mf5aXaZxICM8T9rjz0GkQtkp8jLJIpGS
FM18pf8l2tsRq2PFhvKCaoiiou3pR+6ykVAML/6g89r4SQqL3fGd8ybKJMA9G9gb
mJsuMCle3/H7PTULH2AORkhXBxx98Gpv/7VjKFfQa87ma7eg7U6VmmILVbc0dPSp
8bsgq8MGJWIQgcOq15MnlkUY708qjivl9CoyxGdw6n5uHB6uWAvkWRebIpybrHb1
ayJJoCvSrWZ6HXijm9ytkATnvWz4BJITH9PXM4svn6f1MFzPOwvH+qLK1dfbm0jW
kkEVn3hxDJmWbzoHueAYlWqFNDYFlWhLsR3BmBEB/UFTR4Vmb5GE1sHBsq8e6e8D
3e2YZCvXBgiX2PvN09p7hMYDZp6QruXzjWNfnv0f9OiPAWm7EOWoGRzDvI/WZYuj
ckilIEauevc7Oo6G7dYg+Za/uNJN+vSFb6q2RSxX5Z+sjfFt34BCNx5UdY4UQ8YZ
GGkLGUs/ChFPXSrhxOhlmUYnv7/gCxYgqBAlYOkf9Q4My2X+ThaV7IJ0OxEmZZSV
K9VXF62A7NIcz/T1GOafDgqley609uUCKXQsSJhx0unaAQQJ2y+scY3ovNOOJ0Nr
P5MaN0t/ggwYJ1B7zqjNvOwfZdaOOEHbxqaGG2yQ21isfLVzXDxTYQqSVA+5wQeR
0VlFv5N81RjmluusGfsJH1NG6ItVm3NVtuvgTt+nFRIEUhCXW8fd58oSp2Odi09G
gz8H+13w/BlLFE/xCoCer14y0Y/AkohB7/BfPVxu2GUi1EAdx5BfEJag0Xx4pXR5
HOZCdeuB1F/4xilAFaTdjVr5A4EvdmH1tctPeTjPF8GmqjP30N8gwJHqZ5R4FrGa
jkW6yJGpKak9zEsodfnMYp+K5Hqx9pUfRifv6oPTsgEkzo+jpFKLH3Z13ObD1d4o
GjvFq/HdKmY47fGRFASmk7dQKYrlRwF+IfZG0PPq4kI652+wJDzai4jk0sv2wjQR
Udr5q4QGmXMZtUbk6LD9Ks0C5xo7UH75VM8rVqw9PEJvcoMx/q+HqCZO4CU9gNrF
K8R40UKJgAQc8LyJUcWhOkQV92UZQUADggBmUJw4gtIFKTjHhLDTPTzd8v3ZTNSL
qnBgSUrbL9cODW12u3untW9wTizY0O4b5FYWdz0v1YqOYBefyXOkFxm7qUUnldGI
2ClhZCJ0fwK5odu0wYps3FqQurFAiOayKe6QHZ8onxvDmWXAwkbWUNdslfFVjXyU
2E7OeJN2c3CCav4vPsE84D73Kt1pqsULFvoNeSAc4y+y4VBW89P/bsJYfqkml4sf
vk42GpAzmUyuyaaL/2WjynayCYvS/dvrWMZxTmz/rXeVYOyzPvokiurmxFnhFvVJ
laUPig0YpLHVukXs1UDZIDn2UZD2s0mfq1Caa66z7ilZDgQ4+p9UH3oWWykZ3Rzj
p2Fgq64jxDP5t9m9VrWTMD9Vj4hxfWpVMflIgA+RLieWTn4JC5OwJTK/0zW2vC1d
HKFaAoIQ2YWmUhpRif5OeOeRKwLG3RTjq5xcP1JcByW9IXu3NMr3O5JtfLNAQni3
ysOUZl/cROn7d6sJinW/0LQCiq/etAP7h3clCVX/TXRJq+gV+kE4q6r5X+m+6RHM
EEFvHBxmjD5ibL87uEfifOcSz6M7VEzqw/WC1qDu424e5BQnOIh4i+ZdfofZXG8w
mL9NG6l2Z+QqcNnXNC6O1jhw+4BYwN+bJsJbe+n98a2UKWa09Xeo0hD34Wm5bP4J
9vk3a2pRXgjjz4UzuBhxH7fX1K8pA8YcWHeC4ISPvPIeiFci0H3HVjnVoE/S5WYg
3DwEwjUjk5UtsBDNBT5RtGbmV7XuU0Kq2uPco4d7K/NUA4RX5ag001iJW81h+QwT
8VuyPE1I+DkCXDP+GYdcTrUwzr214jhpi7AL6veXQ99/iXLdN3aSIgBNnPwfhHtA
VUzDTT3+Esrx7XnOp3+mLRWvEss/gi60C3MtFXylY9z2h8o9tmHVh05HCWZo4LdN
YOylL+/DoP+8UOiFdHrQqhvrHVPMEVfxeQAcuzuVsI5sAZP7CHfgH3BjtcBRQcNY
GGmKCy37vvsSr7zYh+osYRI6O6RchJsVXrH/LQTV5tHvjoQFvFG4fBZJwFk0BaJ7
kfjuL7iIxBo3tMEkkS/eK7iG2VxfHiVPdvR6sZKAKIRYmAohRoGADsr3gwiRQAk7
hc7ZD/Ktj4RCsDucLBrJiDyQPLMMPeccu1Py93JxAQiTqihl17QFSEaNwPr83eyT
CKpNESEKUvjTBh77iSgXNo8woJLx0YYGdKpqqVUgi58qHr+JyjzmbmUk2eS5TggM
fASqWGgMERmJmS2xtuwp/6i/jJM7VmZyjBI+iOqSgVSyVYorCmocR0WJ4pgQ7PH8
vDXpfSV8iapElqQum8RcvnB4WZQfYbtPgYynLoE/ECtr5Cl5RKw2fVZJQUXnr1Oe
a7xbA9GmVBzIJAKHZoxNV54xPMTMi0xhGZSm0wjDyKF4RTJuHxKyJ/Xvsv/IgNdm
rvoDmz91GPj6qDdJ/EyYjPtbhMIG5UTM0ZuRySA4blR8jxQVKygv5+8r0nz2En6y
zPI6T3CZN88uozEw2kz5WnclL41Nrqcgg67D37fybcFDXjFBsF+JEnY7WkDwRlNE
wtTnl5p+JVsCZwlxvcvPJg1xDv2Z/FtOHqkqow0jxqfy0cg9IqBuIbHIpemuW9yi
xdCDgxOw0W2UHOv55a8DvalrRyOv3gKjWq8uju1w6rK0LbLRfIWurbtj0R3ItMv/
LA7eHyGFEsGn8UDR14bfpKhsx2ho7DsnqcAjqTcVrp1+s1odupkJ/3eENHbmF737
tFW7pBQKjLPxtyhdXi1AoGU2TR6mzh/NX+MtSFnPxTfzlszGAxUxUYHOypJTom0b
mmQak3L7H4q1XGKQmWU19bEJLc373930IAoyWS+LbYr28KPeMT+8wLcjaOw2pIhO
MF68Wp5//yFbKPlPGIIhXgHVVyom3XYtB3rh19TxkUwJYgz7xgsSBs5P81EL00LO
knD3kY3rUfcm0Rv09mirpexUcDoFjaBXyi2AaYXzgM4sO+ftFaqas7N46aEz/qFw
SI4+5EsTx8yR2rczF4df6irniLTp/eTtF2YCniAp2zQrvMno5vNdL9vNpMkAlOPu
lzLFxHiXhKgpqnKbkHlmHtPg2T/u6eS3GkHOLMuxOJeLsZfKmdPFVgj/DsOc0n92
/v127ynsXD9avxEHsw0pNuwUVHPS9GB9DlCMcGwc/YpE2CXcW0hLKiIHjqOMw0DS
MVUdQUnBcqWdVuvMiUZtn2kS+FbStqifydKurtpqEybMiTsYiUyICXugpBx8agwd
GsBVUGhtPIY0I6Jk+++fYpuklAOT55eTlgzhA/Omj+7HA8f42OJQiPi4s3b0nPNU
Qehwi7bT3IlJJWp4w78PTBKV5mg+YUJkGISVdofHznMUnO4w/ep2wsbotZGgjApr
a307lFpKa2c0f8QkZJeUTlzzqfJM3MsEe1M7frmOCeVS886nHjMdEENH7nIEh1T+
lebrcffktfKUaCbBd1WGzsVYpCnMejpBaeMBhA8f1iULaab3uNkPgiCA0UHtw4+T
yVSEBz29nNHUbXs79Pevx9kmbLMhglgO+Tx7jHh+uT0Kv5+iu0tGyFQEu1t4mcx/
78ZBVrXz6qIp1stGCVEo674vB4+iEzNA+iD7Gv7XPet1yZHEjuRCmEEwuoXp/Z7/
aMWuj4Pll+xuU9KGE1WkrWQTRit+tJoepaYsaqR/ita3/9oNBd+Bh4OduatExKYx
pdhr3UeP7X29GYK96W+8mzzWmmHPEpIrVwIU/MvnDWwqzeaLvFF8prbiLr/QD1qa
EhkrEyWuxYw4bDdIm3esskvhHyuSW0osB4LL2QqJzLVIajb1UBL+7jJGTFqCKemO
f3SmQbRTLAioTrfaTibnD36bQoCUt4VhyV0dFHzhGaYbfrXj3yqDgvz+iOt/l/qQ
/SnTAjxlLLf4jrPXJwIGmKYctuRl/YAFGssvYo5BqD+SncpCKGw32Vo5bMn1Zdt6
SmgZFRG2M929qNlr+kGRQHHh9sBGxvb+UFlpL2MuGgqd0Lvhb2x5UngMBO9sBG4m
Tx0UcArUzCZ9f+VnFSZf3hUrWLHurPNOIsUdWRvjH8thSfIZDAYVtsCqwDaiGjPO
LxYG7evAu2RtbRwqSssj1s3VQRM/0470NTDbzN6TqgRgW6DsSvpRJt9eQfxZ7rzD
nT+mL6YzMjyHMtqOLMI9kpSSp7sJ9fY6iDtSixjBvsr9lJ41c0981cqt24leObbN
fze1l4HTf7ecPUCSYRe6+3XNMcz5DWfuiS6jMRrQ6/btz08Dszu9vWN0pyQmUPYj
4Qw3m5VZ8lKWaJVL2s8S0C23GXIVjC9GJ/CSNzw5HMsWzhMRmMIdJsl7E8w9adn9
2Vp2L2CLqQPatiiqmBIcR3hAu04OLidX4Kvs0gmqP6l2GQDaK1OYmZa9KrE8rCBb
3I9uYet+W0PLFsrzmoW6QiNVZVY/+NJmlOrdGQPGqjGU7Rnqeic1cXuJ39r/azH1
z26PnP+ThNo0aOV7f4w5JxHE+1DuZaMCdOjG8Us59xj9JKqeEl1THfp4oJJx1w0A
a09UPVE645UH+mjr/hR+0dEmyqTqTOmLsShW7Bxj9L5RYs0nXrhHw947UagQr05m
40mGS7vE27V7lLTyADA8GX2ABW8D8g7jjdP2KkbHW0AV+irfvoe9vRA+hAbwaipR
3e4iQNOJD/SrSIuIy0SpOfnx7vXvepjYYp6PQ74t/MckoFe1uYFnasAcwVB7rBlv
Ky7TxGiNTs36ziM/gnRuNHWKLy/fpAN+2ml7xk6m+qvIIuxf+yQxF0BdfgxbYV3S
v5Kw/hf4PE23e/JTlHEGgBEqi+RN0pysuw7dxvNbl8j+Y9zYejEG4Q61Ff/yFyxB
F3vvW9SjfJt+DOx9u3S8goHY3RoTKHBRKKdqDZ3IpdzlTGKUZCNLaiXJXq7oIsLq
mQbu8lKcRVsSBy+pQkp6jlRoP4WoLBCYcMTkbYm0uM7D9mlu0hwSfqGuJ1vvR2wE
O+LF/wRkFLYNRbjknjRvytWIocNpRkPHNfXwH/n2gcJ0sHsJjBfbHFg8i8+bsUGG
QZQIujcOish6BVmoXBbNZzOITK/XdF9Qen+/2NKu1EaOBrTQp/VmuuXS4ugDJLVw
XOQNekLzvUOHudPBhTQK9jPtUPmaccN4x37pQ451ZstGcfpmtLJ/tf2w8gbCqfOk
GQiJxDXKkkBgFeufWAR0Huv9MdzRXTtU6osfuO8OIgogmo1oQZn/PyWnkXo7aTxu
/6Ff2XnXZFgJuPW6rUUl7ak0axnZr71Iz+NrWdBL+VZk8VHcP/3EzQPa+Moo8QTX
SfbiCiM2SS7ilYFUVxW6Q7orL08ZwUz9w+rTpKPkV9JPNOFsmFtVGgHgZUsDfdQo
u8CHOwftV+Tq6tFMkujBtl5AikfUTD1/k/ejou3i17OSK/+OgfkdIFYMSPHcFvqd
FMokLrzdZlGlp1GQcMMCRJQHhpHEQIhJ6VL9g+mgndlWrpON8Gy9+pQdpRVJvHJ0
PNYEZMA0efbuAEJ31R18EEQPwqVS7hzLJLI1BeXoioAJzmdGtiitmMpEKwMS97Z3
CbW35GMAUwBFpJOp2t/p++R37//ghkYwcruWkgVhpo2LrxY/Y8Jm+R4malIH9ZPz
MjIcV7tYn2af/DzRlYai8ygPXTWclyMBEXoTEHUvLiRaxz/+8IjakZVZ3Bg7JWcv
JDcmRHEWx6JpyPmQZ1PxceimC9xrPfGHnEf7j0tddpgtmg5/frhYQK2Q/8gpxGTI
X8T5sT9UaSKNRIbKWNPdLC6zaerZkZbVo6bXvRNO7/BVnEGxTchPS1zm7YRsHpNe
YE8pXZujnah9mBQLFOzEZDimR1s/qdj5tjT2zqHzg1tjhJw6+k86Hf+9COhaSKti
2xlx5BKbrvc/UqIkxzIk/uH+5LmrZbJ2lQg4KpIoVPgFbSW2S4dWVFO/aRRKw/JS
g5axUvzMY/HzsNoVqEaD7JuLGvm7GU/Ud4vBDmkLpKzHK28182AAb1qLqiWfaRcu
XLRI2HEhoTurWoZU1tr2nxxhqUMe/VRY91Fo2TzrgXSpQrfXFDgofNEn+jvs7x/y
dRmFW674d1FOBihKtH/tIfDHNvh2MbUM3L0X/V9K0yCnxKcHoDBhsxswomC1tUJw
y/h6R5tZUDO3ipDPWE9/uXFNCqgRxvAFcL/yVOHy4D5qOO8I/rc3FfAKYdwcdcDx
yF+k+4wa1ND4LLorK4BNwSxz1amVy9FvM3e7asnUUaCk8h+WqPR7oL1Vyg/NgCHx
I1T175UAzHDKDnUq2yChuBOzpg2RZVliDcsTHt8vpgyM4qdoqFFX0I/hHZDD0oRV
8d51irK7bjKY63WryolI9AaRGHBDyC6X38Po+gfYSRlqaqyfutsSx3v7UfVT/e1r
RDyzaRyBvAuYEiqk/zjjxuf6B5sZqFAtjQfYTJviZ8Ql4UctutDKHMkJdYsPKFUb
bJZDKeSeR5CIUbcaUIWGt746JAto8XzPqq3R1Jm0Z1KCm6HrDezr9UOTzNnnROqM
BJsZ/YAPHorsbcYBnjRTqPIvJpM5ZEoLkjWpH9hS+xlf6oEJqPDfYK2omqW1/+kx
eM6tVLvFttc2L0D6eeiYtM0bi6+eR16cQzrM38Uw2EdYt5gddsFXB6Ujx8kWSsaT
XuMuMg7j9WzfveXfLXwdJ2/WHERGNUXz79R15GsUfKZ4Z+QV96jAh6Ttxid54pvC
NlJonjmn4stElwKLKBtDZYzJO7EFPhX0ia0HiIqSnxUQRQz4qpRXKydlrSG0KDso
mk0i8lkSameBMMx3SMFfsJ3yjFANGWolLSoe01RkHW5xrwNXlFZxGNi4UkWtaF8d
pJiFBDr4XYbg9Ooa5EMMnG0EcK9dioohJH5ObmBOVt8bTjAqfQfzpLvemOuA/dch
D8vvNBcE6x7a5cFFFdjN6VIe3+G6Oa9SZbH1np1y3NzkuRTA3jX9kaKnKZuI1NIy
JN8Az+2am2dXu7Jp6sUTvY7QgBth5Xyu11pWU9A0Lz+iop0i7InjIk4x6coXMdwX
XhLd3jXJA/sioL5rjy544wZeHIdNQ6d1hSgzyxxNy2UtnwhvYM1LwzEYxEVXwDEF
MfqPABuz7dl+XpgUR8yn6IDxboYp5JMIRo1t8QRayiPSrTIvgMXfF2iZ1CNg65wM
VbOObD5rUb82BGC36rxrxeFl5aAX5uKnEuISQVMZqk3jNSh+Vjsfo4XhbvE4mGza
BlLcn0D6/PShgU4PCSralLwxVpvcDkfspBVtTLCOLIgf8zB9MlG2vpk54HNCEvqO
xewHDypxceXaXllSCegFeVax5+woOH147Dx98MzszTM2qMOqKCJfMwFGeUKSsYw4
p17kbIS5sSmio8KMYg98D2/yquuiEwN9PmzpP6hr5DeuDYfpuFtVRMX7lNbd+ZUz
TVKyyf10K6lVxS7qg3sYbabMxynykEa+DjjqFZmaDdDtlSg7NGE8Gbt0gabrX2Ji
QoWFpRaDhnyUWol2BEAwfOwtgC54pey65JvGx0CmlN5oXU/89A6EEk/rugnI2bDf
sEkRsx8fsp1OQ0Dj76v6hQ06aWO8uzWp2it2V0bfcsLo+aw7u715+k3s8uVYcaXn
U2NNOKGwTckOM5dR7zOubzovimC/bbAQiIHMWQMcbiBUzREZyY5RyQyTrHXlKqgk
/e859O2v2AFtXse4zen6F1AJOuXzKi7odrWSMQMKmcp95Fd+r4MS1kziyMoFAkgW
DjCceDhqy9zRxZRcSN5SzcE4OvEcyBkPeeWo4ZH0ziUen8WGzSckof4qMUj/wVpT
NqKyIiVBO/ms0D4o5bU02jetUEG2Bt97V81xuNlH3EmjXonMWfA/vPTCsQSw3kaV
wODLWQmy3vUPxvDmgEEPpuRdLkP0NS7+KdLoHWOiuZIlvFrBjFMXF5CAXEz3yPUF
0StXLw7TLDwBuRX4bUapjTkY8/2X+AqWcvDglstoUkxCqL4nvzJ7xPwHBOd9qttT
Zuz3b3nhads3yxQs/RmT/GMRQ4eUiHUOLkAUpxW6kLmA6/+GFzcWf4tYSmDDPhfE
K08329tu0m+vtDzq4+Ozvjehp3L28fnXFABTPeldU5J7tb7ZbVWrsZy+5qtg1xYs
SglHAJNmVjPceL0QdSqmK2GZt+Q3jvhXPurwHNai/zTuA7LhFq5a2tRS86V2/LyG
5HWNeqNtg+dGya8sYHT/QTrTkVZ/x+K1CIiueTSAt+OCjj1SagW0tre0Ucxld7PF
bLZJGgoU9YcZYo48QBucCpEgbkCxUNeqmlJqeEA9ZlhWRcZfkNuxs7BUIi6IjLRU
LyRNYLA6Es3LnQu05AT2TOLntuLuIXUxSJsmQLMqs9HKrqOThFOffjgBLHy6M0RO
RCcx5DLkDFsmA8sC1I6UX8YQSyCSpZBg+kxGjlXTJ8GTOCN/Rg3V8FaE9NSyi2Ia
7c7/drNvrSo66/xnOjrbQIqFdxAf6SiQUwMlUluyRyjPMVh4FZ2F6io8wGc7sMoJ
NcY9DLoLQ3xDilLyraMAujiLDSuFISH5HXpE/GsRdE0X8hkg4sqsxZyuYxY66mnL
s0wUPzzlY1yy+ZwjLD6fFWCF3YvqzjbesENPA3gAU7CLDczSy7JX3YsCjiuHXLcn
94/wag6vSgek4zhNqeyTS92474YizbRqyzlzOQzdsXGGKSPiV3ZuBkA+7GrCKA5M
+hYtQU7dHhdYaHJWxWDw5y5YFCJcPY71fy59LXVA+5t59TRPY+Qow6lgvtTBaRca
LdrwAum/d6CEIRmvZa6UgfI6GOzn/LIwvMKG0kdXzZxH/97s+e6fhb9VQWYuwH7w
J/cMXHH8zZk75it1CSk6yFJ1hnWPYRD8yraFH5Ylqgpcq6hXybzMOtIorR1O0oET
yidZAEzSWvJ4b0g+DD2OFLif8JyZeXyV6wYU9lkKJToGoxxqLvrqXly4ASRNZm3f
c96lpOlWbPlYO6tZimm6GdyBNTw92S5XPzj1BlxMp994IXcleJFFsEMR0alpbAjG
j3gnGZpcCVk9e9wMpyn7U5iS6FKaxMc56+NEP3aDpsdXrauiy4uiRXUpvjdDG7sg
rXd4iAKYnJCZCWb9/D1CLBMt4SU/CZzLY9aKlZiONZhuDOCA5egCLzFfJCi2gPED
SnIMo2QtZoxH7AYeoOb5shu/2aqsu3K276Gy0QApLeNYGxkiuEuRw5oMM5AsqOsD
3N1rEPjk0QRTILC2L1WONloLN9fUlbfXW0n4xdelOYXfpFn3DaNDJkHg39DpXzg7
xti6S6pkMO99+SRbjFdz2OmgS/PmA6IeBx/XJRqvixmovogB1EDO9S7oHNTHrlwX
HWQe2dT0K4bQ4AYXfVhwvoMajWTW1QC3S1uCxtS//GNgKng23sRydk8fFMUVGbOH
NiJN3vdQ0KaBT+Zyy8q+pPHOWhAWzBmHxlnJfREd78qi8Q3JrSVCZwvQV9pAWKHb
yAL/LfpytLAJ+zf5WhiOijVUY/iVAC9EMn/uLIhc5aV2U2J9/VrUSw02P6/nXkub
+89an0QlP1XZEuiUG69IVr7lWSHVlLwZzRWcb5ogibWKnippdymqkA9nBKEllnR4
Kwvk7JMIqrLFY5rF4WJqeOf5nrUsf/lxvZWNg6T2T1dI5HTWapEhNUqn1pR6nZ7b
GwIFG5mO7j7IHeQ8cWYIm6BwZXq/4VOXoXv6eVf0Ko923WRe5FpTyhMob8T3Abto
JXkyN3Pa5wQd5ItAvZlAdIC2tvQcMHlhBNv0QNdnURTI/SuL3CigJggP1gn0A1LG
fISSaTKa2FD8LxNWrR8hPs8VnrUg1agvbUySqO/VJOthokjSX8A29lKdjteYBb9N
PUkrWoLqwLWpJivhr/ZXUNoaVC9WToxRoY1MSwAkVYx2LvZGEqsIiKlZQnjrR+eB
7FqNhqoGvvs4mSD1fjAUgZiJq48zbybJPn2Sog3Z9qC5wODsDyp+7SxUDvMzj4l9
yP1BXQXcAaGRazR/hivpzCz/Ytto+XdceFZRA6F80dyefVHUXUIa1YY6xc1zWKXI
AsMtFB2WfWjM8q7bV9MleodbSympa6oGZIQXMx8RSKJG92FK+k4w0x1d0cv7fsZZ
A5kgd/1r32B2eOqK2h8qUcX3Revr6J861YMfzPtwtngc/qWyXZVuYs85J9PRCZhF
XqkWm4sKeggPmZjntrSTmBHTYQYUoNZoRxId1ClcGRGYLNhWtnueY3Hg4Lmh51FD
Z6f+QoPn2uqoq5RJUKdHVOGdjL9KQXlmQRFs+ZEZxcch69eTiEketMxISsHT98vN
IA4MseDby9w4XYBFKfQB0LXUNiTdjUEbKLzj7yPTatsMNO4PX5L6e2gx2FEcw7lf
9307L37dDMaw/oUnASbhaZKszPTc20bvcVn8hwMrUb0ps1e4HV8ZYmxm55slnMWw
XkA2oYXmy7XdrFThuiIaLQyzqdai/sqRkznbRtF7sUXPEUeLNOiFO7YfFxmBin6q
sCa1lefVD0Rdo+dRcTJRaLEUtGIZ5tXPc5t0rfHItpH8o9ZFOMF4qzYLmm1EuQ+O
4P2P6SLzr2qN98TTYhOCVI4BtD0RdLYZbgnxrj2OhAN/NW5+Cv04ieaPJR/b4aC9
f9QyTHfnsYasbVyd4F8/GkMiuX9AmAmnRXO8cNAh6FYB9pyEPuDup+4kwyuIhci3
7uM7muLS592OsB//TcsGsRnJ5/W5eQnP4qxhUGYbmsiV2NzuQQMnf2Khe7CTCOPV
tLr1E+ZYeMIlE4FWl9E4x2bs4GhPXYyFroUVC3vxVMx54fI9UaoxyW96ItuszLCk
azl4jc8UZq+r6a5ZNMLXCg9hi4UNCh+/HWZ9Ex8wEnrFkmEcYqA+bHlp4oiQ/h63
DGdw2QXBaDGnxVas9dYH5tbYCI0ZsBkPxohhVdPUujCGEmqvZku2ChhjHP9ybvfb
uFdlpGmAwIsk1c4O43euDn1KL3krVRJq42Eu/6UEAGdUY5dJf+qavQtI/d+sjluI
I/ZdQrYOeqJkvLCLEiT+DhwX+Gdsx2q3F9EKhR3AukSUAwk6kD7N6x/H5e6sdtkr
VJd73OJ0+ojT5/qpvcYoS/wvNHDh1nxEyDOTUeLLQxJEqnEWGxZp45xHEl+pNvER
PCXo2uMVslKAO5mSdK3etCUuqIK8q97adFRqGzBp81PpqS3xTjKsV4X6xyawdU2P
BEmF8Jx26PnmH3eBvLThZN9mSTpTOgNIFYGFSjrNbvxG7FCztkECSuSML6XXrz5Z
NK09TvH6bOH1K3xr0QaUP1mBSemspzSjEBO0GwlXUVzEuRWWB9z83Opc3UlrFzau
m7jI2KLrDeKu1hIjJHuJCMfovaS4bDd1SiDpVyfR6BecEmtG9b+oZpd84+OhQGuD
W9VxnA2DQdWE0Aj9S2walEEE9FwMMC77Nj4e9i8Byytroke3u9txmsjB09lUR0uM
H55pZuVuebNgGfLW+vM4gw0Ev5mInYvdco6b65dFOpokcShUe51uZVxhbuV23p/s
dn9mEbiK+0Dv9M/aYmqjMJjR1fSfDoiZywnhkEM1DI+k6TQiRBX7Wxu7Fj0fZTly
b3g6Xt9nz00pZ4veeH16fRBbEfRSoG5Zpy/Ni898lumR1IXViVBaIyOXFIPNGA3o
COwbcpoYwXlsWy+hYKq+dOxtswr35ubX4d1GSp/C1oIPYG2xPQ8IezQs548c1zrM
SPvoWScc4KcVYSwOsgvZ44Wc1v66yTGhMvdiUSgnFacoSUWcs+pRPSBEzk6tPbAg
c4TPbiR4YIhTLAPYqy82qsvdzd+cpT8TYEjg3ycrHgjjvry/4UQG1x1OFAyA9xX4
IC3JpXCJgJzpb394EI9lDM0wyrzJRFUUES3Lauhm4Jc7LUuY3Q5dvNPp9WXsCO2K
wcv0eVWXFl+1N8VanRek7zJiWdvLF34lBTFsn5NzJ3OYAhoaUhxVYcujTPdodAaC
tCQRZCz0g2JUAGp+IQTOA1GMK5ZhKCD7vFrdpjF2Vz/PsR2sSTPiMGBfNO9peImy
dWnTLOey4IUlKHjYWVwSPdiD1XsQpQVBomamsdDq6uTV/418JTqd/ryrhqyC92ZL
k8ShVJQZXltpwLo8gREPFsaiYYebR5EXZRsdu93yiyM6uaQJnYsbWZta6ZtiWszP
VrQl2IhgZ9nNOKPUixSby63rq42VsJCnu50tazVhpJsI3szv65Ec0Fo+/0fks9vD
iE2Dd8gKwqnBT1kMmLmkubAPevQ6bQW8OqR+DundEjbhsXQWkM9NveFBFNYvKgPK
x/JP563kfhf+u/IYIcsvQSoqvNPxX7uG6T//HE9xfxLlKI4qA16cOhpqNc+hc/RV
36UtOeOSvEPZ18GfcPvPn5lOSigjFQmLT98m3UDsfoC7AEbym7lFruvqECpLGN2T
jcGa2iTzeex/99J2yWFecBRgyymY2GOmMAjQXH4LOkShUHnoqKEL93hYenrG5lC0
s8ADzlogNY2tVAC9wFSPgjZqSCBvHWMInrLRTBqJ+531NlEcar90s7kt5zPLz7aq
/231wnpkAs4hw+tkN9Hyn/SAx3jKpvcJtiNyxRfq6ENaMDjj95fwKaQEMTw7Pc+S
DAsXDe8oZPOZLaM/ykvKVIBMNWh/V7AnPfKSkejLiLWuzROmh276OdlvalBuTkKi
UIjkBDkLn47aP3XAeFHCs0mib1/vOZQcETN4qG34jesOhPwDwXhi0ZibhbhTBnvu
8g3in+xhlucqxTwhVHVVHuM6b15icsk33EubgfyfxO5yEt1uU0BtQgYwBaJK06yH
d45zXwg1S5R7phSa4sHWDSs5S6hNOYDGKwr6pN/Fh2nrJ5+57jeolADcGcK2K1vB
yWWB4cBwRHgqwh2p+0KrIkZNpNNOtGVbUUs07dAoJATSFZySWNhMNH+hpHAtSAVw
Hw/yBlWYbptcWOm8alTayugkoRI9WXb5tHDDLWZsQRFMC2OPbzUekY0VGTCo0z7Q
dyccWlcrVyXLLy6+mgSF1fb3FLDxV/por6356GoLEnijJ/qZTO6BHaU21WKRCsQb
3qpJGbizmLgthEEvhd0ng6YGXNdLfsG0Tg7QuoiU6MqxaVyf1AQKbU26pAxAZSbj
oqZx42hIQAQivIy5evNiKHbpoIcvBjFJ6T/5nj+aPAGhQYORTIGyllkKW1FEVFYU
wWloFDpaOVyAov8vLAvv0hIjAtOSJ1ejqcnpZp0gD40yZCwpO0Gqkz7UPN6X1cOF
gWfWE0Rwnu3LxiPlBZ5uppCdEUdUL2K6Oe+f1hvqaf5GCF3gUadnwKv/jdY8WESk
woPyug2v7vBacbW9tGmHSqQs0sCR9F/ctq079M4+qph0rC+/BPNqHwznIVs/4GjQ
w35FjwXH8zBAjFapihxTpuuBtxaZvDJwMlFArC21ilEfF8vJnSeF1lrj+s6NPvbg
dnNImNF7I8eNz1r34NSVB3+XjxcqOwcSA1ftunaCJj8MF9+LK+KWC/AWHldEbfW3
/RRP1259CpJp+MM89u0DAjwDMxXAeiB4GsN2BI/gCXdBWMlvWI5YAof1lpLIiGpZ
IGU8I6oVZr0vq6E1uzqo+imDDnwiesNq1ZovHSHc9ScVtPsNMskX9YBDpykwbTJ8
gSJb/rLQNwvXdAWW4w9qGgRxWqJ4clVftRiqOovo7j58zTqGm/H+CRPf5Jwq99Wo
yWib8QurVj7QjOlOY7/gzdDd5c8nBCqFHkXTOR2X0xBewXBTkac6nHsExKAH4iOJ
SBM5Vwm3M9bDstv2lJ70op8lI7OJe9cg0J1qVGIMavIa1Os5YMrK0UnsFqx6qYAB
CJcBvmJ+ydh8ESR6mtqTYOaY0fvaKAbnxVwwQyC9E4jKUQLsnvilXa+9RzUkcaKW
E5J1RbZ/PdluceGkJZE1e4yMORzjOvE1sSMY3r53lbPAOY/1nY/s2qi/I5r1pfRp
rUYUprQTEnQNUPpcdlHdKrn40403NveaE+GG6H20/CqYZ2wA2PoOng/SmlhlTbsT
CeiUkpd8T6zv4DWErhQG0mzoUGUHGpV4fPPbN/Ss0oeaIXntJyq+K6jgCVbFr5qM
nEB0SnXi6DG2hL0dZySh6+vfSda97koaSDJnriqgTL5OKCLxhvVZM3KWxb/CvNrA
vm5RK6Ke3MyDBxMSA8fDmAw9NGlzEnySCDoZu3OjO+KK1PapmZuc7a6SiBEJdwBw
ZSgTYIYLHrx/v7GeXptNkszPRaSaFShD2jrTjIrldRF9A0kNcTtGaPIjkhLrJjUn
Qf2rT/38zc7+wq8d0aD4fLUIKhETvZCYJ6H8NN5EP9o7pbpme7j2iRSvQiow/9Pq
dPBTPy4wclRNIoaIonG24Nc97iUEKMneRXdGbJE/QH+/1RiPTHWU9vXWUhHl4BD/
SwHAU1vFJ9DdAz870J2vvjFOgG3CJ1tN3p/viCJkniC+8tGrISjGlmJ6Me5fZ8WK
RHrNzxr9O3lbzEjFjU4oEkHNYofqtzVlhYJMvoVCM3dGcD1wuJCBfzvf5rgrgGvF
6UmU/Zi9KOqk9R1LeAlNw+wCIB4fHqYou1/8zRjyYd8a3rI6NEacTfTBAmaDNdWB
EySHYVnCWOx1kuPrAL8vtzCP8VFXDl914PB1qi8ULzUwZqshkby2KrlnQGvH9U0B
w9FrGJ13N8tQMKCdbDmLoQdlLX9cYN/rFd3adyiQFOZgDGf/Cgrh6Z7qNL5gu9tz
fTB8nSRvPqQOp2fd2JNMi56TOzj7cOYlpIvXFUL+D9rXqnY1DHDMDjWfHLvz5fbD
0pLqdrl40Olugf5lMCie+n9RwoIBeXVc20I7q05ndrmnF730o+CjvmZpO1+6OwyG
ElBmU9CoWjGK4FLZTit8hwr4YjfTEK84TCHlNcX2EjD0t8TvX7CddkU+GxckAKXG
UrAMiUOzXoGsclW7Wn1J6+f4cQI2kkmSyI6vkUJGdTrvBWmq+D5emEyEjVHVYmuw
z5s892Vvz17Kri5KEF7Lk4+Xiz3znTVOVYd/43SBv5YGK7z+sbthkhGEiXLjnaIK
eucQg4PzPIG50By4TgIRlTveU4j1P4HvxZvqL1SpfqXRQczH1G0JZ+DvcYyUdrhh
kDGHilovaRgjqzV/BDjA6T6SctF9xaGCNAt4y7sIyv83sJHAoTLdCjEUDrsQ32ha
8BLWkdZ5MlXXLdp5jklAR/6oDsKguqB1TXntXRd7sg8rP+fERzLcbZs8L+lEyrNx
YMQTrviSwVRlN1XZweKUKhDWmI1GQOfMEuoS0KX5Av1YgZGbJhs1wwYOWh451wHQ
qi05VSJHcQO2K00O3WEXBPeuiotEVhoiAZJGc8zn9xLuiWrN/HyD9Mss6u2D0k0u
+y+UdlnHs/s95KMQJgH4m2sMgGDSnaYLnhK1v2xnKl88kgBwjT8X3udDywM1Z95T
qVkBAbSooFrQKF4oKUCwVR3m/hAIW2VBz5wg2HjANG5vi4peHUghAMl8mVuS7Y44
ElhaV/xB9J+jUwe96TaoPxTqD6EHBPNgeNf1pRwA25OrevGwW9MPjRjy3MDiegYu
BfVUBkYKVN7HSwGBl9BNuFKpt4qh42aIAHWtTHziiJUJ0Qe3YOHqVdIVUJrfHO36
CXW+HOAhlR5GjJ6gcooW15y1H2ykWg769bxK44RchBfvJs5HiM2UqLN+nz0CCTcM
UdeLXNCrfVpNJ8d7yxZpV+x5qUsBIWzZpGHVBA3Tn+9RAk3wObfz/IGPfaDpYuXk
gWjQIxIGoWamK/a3MFDIsUN2cN7N+JuqxLBTffMhyGTarcx7j7RqFjlAT9xleJJU
QaBCVHCLmWmXcLb17ba2aiHdcpZziyTZcWatUiPBFh37rxQemF5nXbznNky12Pyq
MImSIXG/mLO7XheQSfSWg81A+0gDxALUOOItTFvMlo/zU7j6am1PXLzbZvz0vgY+
AqG+QKgnNXRjvLiPKKpb+25Pgi2ziyjQEjdVItq6BUFShm4B2L3ERNcwW94KMkjV
NfleXjnY1PfWtXjI8uwN57J6HyjsXxsTXx5TtSHB7deA0spOtNsSNze1BHgcdZQW
cl1iMrvABrd8OT+uNtaHx5ECgDuk7zuzkwnPLVWXkuLD5gEjg4G4nn9XxjOe8No7
GjrJ0B3DOsY1lrTEhS4VzyGZqbbyTeXW7BxM+9Liij+gYVxAkGwUJhl9ghUPt1hQ
F6PLtJTYB89gaL1o12rPdVGMMxWR158yoHbNpoaCOZeNWGY2FHwXGybhuQG3a7fF
hnu5YsJmH9GAM9oD77xgKYLam2WyDQkoBZqjSMIvMg0dj+O/D333kxZZdwk7RUIy
Xp6rpwdfcwzBddQucJHauU06SDZvS4eWaVfMbxS33RiKXOh6JiORCu/5nBkOqDGG
FTY6rKo/xwj5iXZjwD0UbdkkmIIsV322IaM7mI/76FYLIFQ3KzZ0XJpNm5rN069f
JybDGiZXgjnbYvCjHAkpO/lXpbCwqZDQJc4+/h/hf+x2rLlVkIYRTTOuc0J5p2kI
vIMm6cRS9aSQqaBv+UZY2EeVkNsW9SBqhFSLwAxuBWsIlRwp24b9fFwhTnIVYc8W
zaZqMis8sCJfqZ+Tga0St8bLf6vfeEIlSernNiz27Y9Q8F3Jjo3rTTkm343HclEj
fDDRJzzgFi8C4V3WKsEqprZI8yY1irDy1z4Ja+2gxddootvQ0XUQqRxkl0O5WpfX
XUlK5O9EvHFZgpd7tgSPoJfIp5I0gzJJ2Rd/qA0k9KAt3tOEY3ZT2uyx1xIZedZa
6SB+IrSZl8YavD6+IybvFi56I7CRrbHdqaqTy6c4aKiumb+1RpNoaV23XSs0bG/U
2bL2c/6jnNOrtT2ebSNdeZUVRKAqCiJc/D4dn6JpzEbInFzl9RVYxi0BI0tibUA2
yhFGABkskSOJ0FKtwPhBvnwwwGZNq2o4sKIgocrk/guQ11Vx0XKqRzvrB+pe0GPD
Dssz191UNoT92FUSSq27qbiB3HmaEJ/34ngYbwWgl/GACxMyE2kS/7Iotqo/niRh
9wmfi+YXyKUBuQFmQglw7jSZQYMKa+TgmBbqvKTW51W/FENR0USbA6IxpYbZNrn7
gxN9M4TpwezDcpC6Ix+bdbZM3W0B8RIAme/Qba7yKeoU1CbtOaP1Y+imxu3zMIwu
rp6F3BmwsInKOFNQ+MugRPJMP6O9yud9q5FjbFzo0gXJT+qfZdoDGN896I6CdvuH
MYVw5XES+0+5PYh4cKLq1OoP2kxxP7XESlBcDvsMFCG96cRZDaacQOqaybZRi/eB
hfdxc6fPScBTgwId01X87kc97n1Sho3X7GGPr/Qix25kjlU2nDJp/PxHq/Len0t+
G9Iq54tTG+CpgxL9C41+KH9WbaHVgnYH/No9+RNA4gB0zUrrlTTerpsX39UZQ52s
BnRuJ3BSSjnvYeHPy3LfgYWSEzofBd6+7EMPLIN+VJEo013uef82Vr5iPf3nIJvY
8WvA5ZxW2ZboDC0wl69KnLN6k8RlzR8ppOF4Ji2vGFvWkZnG/7aILVNYvN2KLD4p
I06P3eoRHq4iQnykM12zD8LQURSrKHVEiArrEfO8L2CmikXZlMmhWkl0qcYo9hKw
IdA5Euv5AWQpq1kmKpeS03KoysmyrBuuOYGo16cZJNO93wMBv5pNasUrcW58hH25
uyxCpoDABeTgHbnZDe+NhmnQQi5CregiMTPW2UF/5wwayzspX9+awrh2kSS5cVpt
CsmY1rAx7bi07yYjAESFgBzsbCFCmvOUacw82yJjEc7/ws3FKwW5YgzYknlwLmDn
oKJmxThOiujM8PmBbHvADANfmTzs9DopNRlVh8iU5/dwtFZWTav5XdsuOjHeNGx2
NHn/k9EDW94nE14XQgV1skgeekTGHs4fjcy5t9HxlCznbeSV5zJ9dWudg4QO0WAz
aG/dZ/E6H2tPL2/edivPseS0NY9X3joMQqUHb2WgUSv1Yu5YhU2aTuU5z50SwWH3
VQIjKErhtl9rO8DygffLDUUDutHTQZBW+FGyEPKDPai93Dm2m9lGJspRDuSsPZjt
cvEr1deJRV/J3qe7xO067zPGHpyGT4v3S6hwjAZBMoHjHC5NnlYeW1dIMV4q1vz6
aHhDPzvqTxNTAw3rBlJb2q5NQq+Fx6b9o2QH0Kj0YVNBxPKT5EPrq0PucTK3DwYL
8NOy4id/a1iTWN+vE5d7ce2KznXcb3gMP0Lw5nRGhhSR2GChKofoH11q9P2es4Wi
Bw/hQ4cqVbPkgcj2SC7c/tB26zbT2WjHqoH8sdQMJDsx0/MFqAhlSP/o27xhHY2b
wDi1GwnKWgJV/zAVGKwkpeJTKPmeLFJBefdLEnQF2YfToD+A7FEfEhXrnFYI2X4f
H78I4CrmNX9JWr8Vk1KOwQX9M77iP+5xh+usoFFTijEoL+CE6hccDl5FT56LLkPc
K+dcyuZV5Uw9/JNUtoWE5rHIJz0CEITDTwf+w26pKFL+zKwWU9wUqYAlJauKAPOL
x2rskMQ0LbnBoxxKibjRZRbXMQLm6wml6pUdUAAwgJaHi2t3BGu16TBH9Ygt67ml
i4P6tap/ss6/cXdPI/susZ5iBKonfptVHBiuBvsOY19NB+V2gmVcUo946Wz+eASU
CvIGixeW6QP/Gglch0/3PFpR7QSjKdPOhg8KTUYyiF3JUwKQ803VOxPl0pRjRjBw
c8EStvu+JrfEGFwwevC5Uo9ctc1bandYlMGGXoaGy0CzpbVo3XlH5QlTv3U1qz3V
vGfZEMlMVMQUHwtexUPOZfk3eHjdcMuNMtf3gz5xgyTzj0l5glQ4+2JRNrXf+GW8
LuTX+ty7tU/hgis7llFJFyvYIunYA85CvlOv85F8ifh0gUlNackr3BVFH0joFlBh
9oNKJzbCFMs4K1ZLYsrgkzmU1LvqdRCVTDF5tCaLKwPjzDFfD8+C1Ef4yz+ro1vm
PqWEIQoc40VNJX02EmywPABjoUgbbfrjQFvphUu7AxH94poOnSEq8x7I2eMkAN6f
t91oCTuDgd3oySK0DidMjK8idpdMzk1o8+uxI53g4u6SdeIWiQeJPtTtM7fJQqvI
AZzHrGfGSf4tjutUTzzuIHYdwJ+5rowNYf7A2rqCCohE8SquOrPVTJGWgN8j6a05
7kwenWrJ6+3llbpZU2b8HD5N34MQERnWFiy4s5AwUqMo7rL6qsu0cvr4h5zlyjmD
EVapx+midpeFOpCAQYPB+KVZOT6yR8ggsMjoAnvMlxFlj4TK+JVhPdGfyQ3Xs2kd
WfPlQF48b9r+Qkm6k48Tyr4TXd/6HH5TYukUN7hGVBx4ypOwLRVyTRGj2+o0/cnH
ULbTe/j74glIr0KC9JXVo36ZQY52UVhB/zZW9NhP69iwth9UmhDcsiPkvgKdWTe9
uuwv4PD75oVgBoE5OQGjAgD5ewEo9gr5ert+XDnS0FB+sc+FsN3QiwalXLtb7hGw
g1hOovZ0E9nVLc/5s3OkVPtxfOt9k3QsQmliHpT2Cin4AOFgMtTxyIuhrQxzDl2x
4j0Hs1JgaXsS74cgdWx+YNKUPQnNvjUCiI5dDR6sPyBLdsfsG6IevAqBMZIsC1aH
1fJX7LSrDtE/KtqsskN+91EVAczAExncpBs7qvH1eUJh+sSaiLGxlsfbngOyswRl
d9/bHKrU5gmf5SYbVdSygJhK5fktaBCwmiis4AnJ9B2H6LpyTwVIxjhEhNqJX0C8
7+SCkSFgOa3oggAXKL4nlGzNUa3hJrkQFJSonQt/mCE0f9tblA8Vh4Kbv9nzK+Ip
hDbxn2iRwWkk8U0Tkz/Fm7+AaEwhqccxoBYdoqSyuDgzC2o243zmu+07gKNjZnM6
kxIwbKNKGtBxE+NQWbNW6jJE3ms/DUKhmeXGIHODlfCpLFjQidOpvMNsFC3jG8O4
sfcPqMK1hLeEUD1fyqPEGmUZR6SdLv9Jh3PUqYdZXiYRC+VSW7hXCbHRSvZOL/VU
qVx8io4Ual36c51QeURjE4egX3AZ7q6rltJkZt8bC6XqyM2w1/9f8FEZTNvW1Zhf
zGfBSkFLP9XS1cuw5nCx4AwJgvE5+fThEgwzfJGrYQ3mTUMb491JWntiw9YO3Xtt
isXjYFhIVrtB5GRDb/P5sa9cYxizhvzgEo1BVOvHj+de0gMwKIKQxJupi9XEivNP
Zd8yLUAuqV20pAyV8GjeiMhp5zK0Mo82bh2mY3HadJeHDP+a28PeFDgBhlFnDXum
mjfnqrjUkmuK6ZYkAIv9cO21rXR0GJTjways28kvEmmCTOiP/DfqQnP3u3T2wsNp
lpOHxJ/kzQ/vQ13TOBbSgCnk7+hbASVUXExdg3e3jrIaViMBMdVLwYuFl1FmZEAH
BnW3Bw4mlqbwOFEkDVL1mMrfsfgyNZyg4jPdOonywRm97OT9s0b75v3NPSEd9UXN
cKY37A90yhgYdHCjDElzj/Zxae6icnjYbOmxhoES6UoKmN8441zG3x7OEm3sthDg
jkxKctSspr064D+W+Sc9MA6JttCNHlcHOJYwKfb1eZyofBGC+Z75EnV0vHOHFxa/
NPb5dhreeGqemNLpsJ2/ogiDZKw0lvklu6I3awoBGGsF/GKhM2SqKsBi0PiPEltZ
9jGZUOW9rBDn6koQmA9UHDVuYhaWmphR/x8OAQK3SpdoctvxsD5AbzuuomGHgP0B
WmZ1CgZUpOLB2nVS+Olo3HKHF2WBJqS+8LrvF4QVoDE6bYrEs1KaLMcAJ2ShR8n0
wHeFQKKv1pwphbTFKr/sazHODVYH2fQtCVuJW8voB2nstl95uWhfcUuFOVeXhP/b
P+IOQ/2E+US92zGGzbDY0x3uORYWY2GYC2Z/XlnLsMk9mAfZc9qWJwBV3c8/qW4G
0vYtnNTQ5sxZNSp3xMp1Yr9pyJ1LujjTuFcAEoK77FFi2IljYCaCWxr+f8NS5qnQ
+MJeye1nfqnGbOl899zDIlMDdKuBQ9CMU2PqKLrkrNzBBuQ0OUoiNc+C1RNSg3gD
ycLMY9L/osD6imOrsUfka/w1Qpwnt4N4I5KoKNx2gbpeWnwocfGWppnQlnJh8fqa
cR7EuqlPuiEqkMkhbm/bCPcU9Wvcph7mIqXSFdkpnu7HgXF6S3M4bwd8gJb1Xkk1
4N+oP7sMBzOU8ykYRUni6bDOo/jBPX4jo9IXBkmIHZzZQP6yyxyjMKO1OQQHyesO
acnQssA8lTSj8qjOIgLnCWhS/RTmypr196jEefM7QTCLpdz3wwtge/xxetzUVG8L
YYvnjzXmvhKs0b86hcO1rMXfvWWRpS0NaK+9bl15jqsb3cJhy4LyeMHwNLWZvurj
EbMkEDQ9g4qN/jlbguBkV9AQwaV5xRW50D5dfpOHcLSAq3y99nFb5THFF9MDVA9T
urXjJy3obrNUV0DY8li2HDkVvJfN8GVxRVSop3B3oi/JnYRHCzOIw4/+PA7wZWxQ
h8B5+MuUaQfA+L6lR3vHikP6qIMf5ZpoGs/7y+d8rjGWCS16Kq2w8r6GabanuDSs
ukis1lIjsJ/sUdvTN3/YkfxNRiUabaW7rj7UIOG52Vbm8srZ6isbQS51DWiruTb5
X2ZVDObFljPn/Ft7OMG3Hl1cTSYovApLUvx2CuGg4v0eHJBVtwjdfxyZAhlCijcB
gfT2o37JCmrhcm/XW1VOyqKDVwJWJKHX6ho2KTFyg2mqeX7YLmqreYe4/IfTIiqv
pegnMl3KILzal0/r1v4uuVl6+uXDvjsZZRaKjDeJmCvKJmqpLrjiXyiXukuR61OZ
Gz5kdjFzowfmhOOiSR5mXauWMVuqmDGTYmJCG3XkX1PfFYh1oOvrNeXS2jgs0gTd
hw7yKUj8+YN8iGyiwlEA1/Sif0LUwmr2tFYLjN48GY/jCDzDv0DkpK9Zt//KvMIo
oXdS7ULK2G5DYFvYJBMp3lq5EmiMjBSWVar7hBAVrjddQvpXQttPeE0wr6xzpLu2
O6aqTYxhBakANMyTL1vmIK5FDpImY9HbiCqJ6DQEVcmYqD4QSQCCknJzOP9Spcre
XhttxPfzf240Cgwu82z3cOo1lvRrxNJze4HCGAd5ovg6HsuWcul0Mhp6p/bbP7wh
P67ZpckTwofGoCLqA3wuAOmn9SZx7rp7w6bZLHFW8M988HpjusICnd4doOpXiN00
M9N8C0YzrZs4lojJGKy1V3noAXp4aFV4pQAMRr+MIwy6vsdg76OMXTNvI4CMknqC
+55gy/XeygraQ4eBVvcGbdeMUWBq/UwDFmAtwnFYGydOPOE6MoxI/jE7maIYk3i0
KotVeKEM2vJy8pg8yThu/p8YQaKu4Rtit8UZyxw3jHv08LsCRpOuixyFyzqDUwdK
cavRrhZkPpfJ2Ndhd4g3LYGz9dq48RJvOzYdR8682HJ6/qRAjKeJLf1YUrGTHfto
Ua1kgiUF9Xvm9UN8djW0+1EoPYTQPPNfGJnQuZi6FqOA1r/U1f7lZpljQKmP99dr
tOekUwY+N5VifX5IhKgA00zBQaaKlXsy8dSvUcNzm/lGmwRe+6w+i4os8EZ2fvHZ
ECd+NL16Yk4PgO7dpTXm7GfC9l+JrQCFgI4rxYKwJLtDgoM7NL4Yh9bqKFp/+sOd
Wd249b+jdmw77Xe9FyOC472PPXcrONW8ERPlSpKyu5oPoaqoQu7ywFzD02N+/E1N
WgvzdW7cXll3wN+54jDVJgd2oFjETCnp13uOc16b1uAPul7YKlNIgO1y95cZLK2k
ze1IEHvru2snvOw/eARCh5w7OPI9xcVU+0FS4TIdocbdzR/T9ex8+K3XiGNx/fD8
/SfcY07JI+vYTgsj4sx3ytj0+QUaAqjetHnDXQg0ef6gSzIWRz8TeBAdfNnvASRu
rpR69XFhw0unyOjPUg/iZNGSTNzgyTeDWPXxF9Eynbd/B1kmlcojzdkCoT4JTKql
DNYBTalgws9aGJefz3frcdbsCIM2sLGCguq1wKn7TgF/7M+vA89wYWi+JOaqTUh3
Oo+2zqgol3egUJZ6e3gmXE2XpKXw5SFeFWOFeJSAqngHGRef941Ubo8B1sSgWCHa
oe0JD2oYbt/EOsKSiIL188WpO7yx9rpO0jUQsdDTalQDlgaLORlWesgYx8T+hL3z
twDDv92l1urh+18pHJdJ5VFyc4pvEWsa8dp/UUJELGrDBT3f9C47zIy8V3aQcbJa
Dd4V0WSWy9rvQXv1J2vaHiO7MaBuUAiMUrZ2xajwnCK2zgsOCp6OjYLCX19B3Bey
QXnH5fs3K9xWFD45cVo5tvphfMzWAvl83HSQxhwyBDeI/ozbJo+8SgkDHPQJ0cXN
w+EIYoXmOj+pMXqJ8xhhm99CqH6A56IuWKjpXssK3IuxRFYCoUdqlf8/18bf56cQ
x8qy+r/Q0orY0fE6xVHzA8e0MXPVGYnyLZPhc005/YkgiWSIRZnPg1UpriD8Z5uJ
U614RLurFv0OsCYn1Fbj8xfO/KYCqTEzV+CGy47m+H056XuGr3dCfMvekMPNxc6G
kMDpOD24NJ6QsLfRYAiW2AcuwGyVDwMxxTY1f3VMwrjM/jWBrfShhin+mXj7qt2G
VNsrrnH+U5QY2puJG1+6cLV8QpSmxpzO7fQRde2AZ6qMdHGnWvEdfI+vATzgETe5
Tcaw+YQV3S+CcRsvnk5hYn1DK7uNICGxqmxnq+c583m8bMWfhzY9JK5MqKGIVFfU
e4LBBRVMPvrRf5vx1jeyZJflbdFi1KRUHXmn5hkpq+fcRUk91KzdPLaq9hqKZPSR
FSe04WjEt9Rzr07e4bTXIiJ3/oxngYk48OxmOXTsU56nYR312NqHN9DtIWQa6E1i
roJ85XQk/ZCp7E1M5m1vfQG5wdw994qHo1Rt1c5lxRyJpXbea5PyjY1v7wAQA8O+
Oj7+gwb3SMEvG3mByA3qduWKd/fhjtuMpJ6VOZGGX0TtE1cLZregJgBAE5U7Q1px
SXXmP+eJkFnfkSzdsqPocFjyOIEM4bG0kZ6MHUNlFN2ZUFOZnZwhwV6sxVwIUlPt
5Bfr88sMQPe8YXGyo30olBfNUKs2ss0VrdUB/Hz7LeB1UEwYKUhndrF6NlJTDWdJ
1eh0a+tMBdjX6S2Gvlr0IpuijH3JCcJoDju/z0kPIhZ3407wt9EnjTedjXxjZOkJ
P2bqHPHeQFOrnJD9bCRwUhiUTbMNZe4q1A8lfL/Qg8XwiNe6MbeEoTutCw7xIDt4
AKhtWs0EdWUqRbyrDF/b3gDTgzF14jQ06Gv9RBcjEJ7XHIRRA2y5kLQV7vpbtKf+
ltS7EdBGRxg4WyFJ9z9wvUBqRrWFfyX6YLhb7+0pUBQqPPAi/ewa7pY+RAHxaEf1
T9PUrT8k3UCZ5yRvBwDWfQiQC14bjOY91ko6zPQWiHJcgsz+41r2ATaLLHclWE5r
kMBI9hBuTa021dRGCvd9Avxa3L3mztDGj9SCIpQ8V5HntBDekkK97kXATyhwuEua
/8U+8c03NrZEPOsgmQMA4wpdTpDaBbP22Lk/LFD7DZMrIK6xTITB8JQM0ld0o9zS
tyPRlc1UdTOUA32IU75WSws3Dkn6ff+rkk6MhveixxXsp8pFEPOvdCWiNrwPv3pe
0ZFPl48fS58SRhp7pwEwZs0jRazKf44ryKVTzFHXbl7odh1vEkHuG0z9fB7JtyD1
b5V7cYEX5dDX0rh2wAg6npPKfb8BPcg64/naKhGqi2VeXbVbF7e2hbFNMN1+KA21
8W+ZRWDFkm8F+RCRsi9XZTG0mE48kpavsU710785GngiihJrHOXrh2/WXIYZbzb8
IFuTk+f+6ozV0UNIcHTebMgbk8jX2fv8m0CASmJ39VMtMv3Wg9jWGRtc3rAwVVIg
/6a1u/y+TDuuR2/kIl/41DV+mVdHTjU+o2oa26I3vqaBQ2wdkVrVwpFkvQDQ1DrA
aQLncVIdSpx7Vbl23hyvYcz6slSwLvk97hP383uQ4tCeC9cTxgs/LJ2G3yCqdffl
AeBwoM+CgpVBbex5+8XMF6JnN89O7r3iwwV3wSvFXvnTAbWaW5OZA4zAvNgHaixb
lyj5Y1rMMKomOcZKBNZ7KGsVd+vcPU8ALlmy0wMTL0cxHQAXjfgf3P/kx7iQyI7O
I3AhMxIcy2kbfGGygqfMjxHl+lVEm83a+PUFb+3ZOoYGkX8wtlsd79PUJZmdvfsy
Ga7M2Ixonz6S1igLeWntc/ZR5+JUMO+fo3XO35KIQt0HaajZwXRExx4VplCoLntm
yGLskWyUufM7YKCRsFPclafQUV0b1StL3Rsge43TZlrxJOOR1gzfy4IX58mm2lWN
f546g23bmBmlO/W+5k1dmiNDTozRa2c5f3f1Yeh6redNDvdLi7H6oG5Utd/ER6Iz
w8JM2qJu58yylQDXq2XDHQdTjfdusymoo0BhonfYIZ6D0GxTUDVMhLcgkDSEgvQd
M8V0oY9bggNFQK1vi3dvSZ2sk8gkNU8SqLG//J26ln2hYFo3yf9q82qEV/EUdJEY
1Ekpl55f8kRSo6IVKWzS+dsY2Rc7l6uENj4E9AEL2VWCO/4wEeRiGuFf+ZDJ1Fry
zxILk/6sAHhDpQA8OAR0OjiWnH59S7/UxktgK6bFGE8VKdEgkjjCVmNZL7BxjCKB
Hj3nFNiG2MqZxT4WcazT0OMSIbue5GD+aATC4GhSrqsytGOBmqefQuPEwbaLyzbj
MpKu6DRXiFBT20Gdv9S+mdXEfhQXkm9KhKbMl60LLQAxtjLWay2zV7GVasqBNYTC
JAJBxkr3dC9zbCB6CAXz/gyZuxK1rPwFkPcktNJZYRgjW30PeJ8+53q163aBV59J
30NxnJohp3JAaai5WBp0SYs+PZxfOafQcm/Ff9MI9uVU8doO/MExwq5hXyICJVWp
F4hY/JDxR8m6KmN+B3rTUpJaU2OaxJD+vq0qzmeS5N6wuxMikC7RlZCxY2D2NaXO
Y2blCBbQI6i/z9zUnzWfG7/zY//ZoC3c4eDkPTjJpYDVYF5IYM57wXcW6uYE595U
+TDwmPrqIT/1O9N9CKZR2XspSraI2/FZk9pr45BXUYtrgrv9xLgnFTSjaJrh2B5+
EImSaVnLUkjFIeDz0D9O+EGYXgeLqzarVIljP5JWhqJGYxp9muTg6N1QhUoDCDUO
QMTezn2WD1vt7I/3vMpwUp3nn4P2WICdKZK9FCzFYZL4j+0XqeSPSpf2YYp71j3w
Y5ogfsf+7sWfSWK2G18a8/e96y+rkJR8va4eVFxKwcXiBKT7okwfMfUNZL8DtcuA
C056xi0SZdHUePQAZQ0jAXcpb2TI3x2yGkLQX+VV1xelCv1OaM3rksb2ks/IOq09
9nUTm1WykocC/nikvEdcOO2VIjW3hORT88ZWS0VHunGMlsi/ZOoGEoc5WKT6iYh5
Tk8N8D6sUyaF1PkKkb+b0a9UUU0HRW1pPAb/9VNptpYC46sNR3WlkJ9TY0tuNP9N
gXj4FW+pxQK9FIboFZfkcHNHYXJ2KNX/Ar3vh20bcoPLvQ+Vg6/18hrU45Lbqk5D
93rDYEEKYFxI+Ju06T4DStHtL0j80lKZWR8zfAh8Wx86rA1+9IFUBGwdVlAR6vrC
XaHTHk3UumpJdZfOXrQglLvLOFKZgmbx/SH+8GOLHziw9PuS0rNQ7/kuwTsxEqvh
TDgexue1jjWw8CllA7+Bigk+EKx1ldbZ4XfBY/dqSESG4bV47GLH4SaJjaD+sFYx
gtChvUClRzaYAxPqO1/inWQJnbLPW+hN91ZSo8hRKKwx9pJ3GpuWDfJ70GjKZT+K
YxbRVgqnqg4v1bqmwWW2B9wbDNgBM+FnZXtkffH1BR4YRyJqi6nwRJURR38qpQ3T
APNoiSKsNvWtDM8gnOxCiBceNp/Eo7fwv68J/xhYoGtb/tVic6RzYBLCdt/Nn4EC
1+byaPrtlXNPIb0ygR6SFh06jVSlnwwzpSCOa5a7CMmZ0frwT0Kpf5L2WXcjtwcz
1QuCFIXwRiQ6oKFa4M6cNhae2ow4omHu9af7V3vbEwX7QEaEFXBr25YKiVQoWQr7
KVKb5wsuCvdkeSW3blGQpf9bw8Rv9XuZ65DPbK0wBrdQgRFll0uaIwmdpfyFVkcl
AjmUY/vHPXYoadhFoyrODPyteYCO+L7Y3AKcrPDFGtadG13lfaCoez7rjxjUToKZ
MGHAo6ltxeYe8XZ3gF0DCo1kTpaij/QXYZqUTClcOnj0c7eXMRcE55RqAWXuJ/sa
DEaeMI9VXLS6WVQATB15923dYPFQzsmw12DL0Mv57JPjgY8+KuHJzX7kBPcS0aWw
KnGz0ctGtnwFTnD/07O4Wr2eW+D8UtJ0Tj5AP7HJyy2aJqDpcU4cla9r/LuQNRst
I87ZfLUuzQi/KJoYk4VDJf4bS9espn6f0wN5ygfy2wwE7nptCDRyzl3jQOhUxwDO
HPQ+MR1X2x7A4pykT4Cy2p5XNPXUyHxLp0AaJgdbAClvZ+lkjcXloMFu/8IdjRNU
/CxmEFGiftPG2XH5seYyeCCIBcM2RT8/XimnyWLTFbmiiJr9EInVGlvakaUS+e58
ac5ckasOgBetpwzFrv1cHfwRW6qQP6hWrh3IEqV/Do1sgmEqSGr2i1IrNbjiXDwN
3jvI6jUXTR6PCWKClTse/JOerbVmIC0xdTWLVy5XuxjKg0ddRwyoxCbEBrK9CRtQ
3zpbMa13/cwt+0WeN7n6DD4N6M33vJKtxnWcpOzyjtS3GZ3xmSQZT8axdVTbL2sZ
42ByJsyppa7fbpnXMOd8PvNR6kYopY5d2WoV0dkCvUiPf/Tgk6VWCViSsIQMMMLR
coWmPSg2/qufD9kZpM98EP78Hr9uoN84ODltSpehKY1/H1yIrSpv5R3BD+1TFRVm
MXMrDubCD+u1Zy7aMgg1zALVrCinLGFQTdINaPbMbc2jNtoWba3OVv5QdO6OTIgB
o9/1mHcW1x/O89XXGms/BL2xgVvJ2D7KFcqks3NiWCZtrA5tgowG8VOqGuG/r1Jw
abWpUsdjktzVeLsO0dM32rRB8RnYYdu9U6bt0ZNh8CcnWLesDhrmtwhfyez1NH64
nwc/HRtsAyOZ5wqVTbz6AYKMiTqTtCFGV8Hzq8ZOilEFc6e1nh5PQ/Nj2GQLVRa2
mVKliO3+F9G4b3mjH8EW0vG3cDPNn4q7DvIaX//PrEinCxs772YfAiDIvoBhGVPO
sSowwgfx8qRb1yBfYF7WNW7FLsPN3W3ScOnhMF8B0ZK6dB4txy+nVJ1EOhvT4yJ4
25AW913rwOBlm/ajWmRpx1Bj4dvr/BB/KlLPbJYARlms7OtwqqG+j/xdV+EeH8Zt
MbsdPzLvsECgAVqwIikd9mMhIvVxvPrH7edYa76NjS0w9I8JoHTG+vSPS6xdmJol
ldfmZSvfE0vnV/6VszCiXYBu/JEUYYjy6313pzxTHsJdw/k26IjFJDkxMRid25yN
KY3XV96k0s52R1aIQF6iKPqw44WZc9WUEYGpBT/4GuHYvTnSlaspDfgrwybpElAQ
IOTrvFMHvett2v5qN6mBSKr3Wr4hOADb1ayP7QMW0NP19SGumCzhHgx9/f/vWcUs
KKUNuLu9LsG+OClGteLYOnepzJR5C6alQf8NZS/9tknzig/JrXAhRTWblPN0eEhw
1W6kdwV9XbgFVntnMWe97KUQdmk33hfjG2xVayaIxTbpo7ZmCw9KuvfY9Zf0ueeU
6KvwYzQxj9IJk3oJ95udfHlYmBmu+2a9nGaUCmxPAQNr/AhIuc5UM0mt/d9SNjYG
saR4lKhWpIEgXWt+mcr63i6n7c5ocEWnPFT0n+tN/oVrZMqoIUVk9b24tQVaIhXn
quPsgJkOb8ozJcCc463Q+33yw2C0P2l0LVnxkE1FPzYFBE80H8XXuKjVAg37WbMX
zwyoYd92pWXJkq2cKUZkviA/XrysYwh08g7jMLdTe54zuJTIeod3Y+BjqDz0ZkOp
e7XMw71YY+UaNgWIajlx0HQwbsDOFJylKn3jt7Lx5i8dqzwstANGLEVwuOprYIxe
mNldT8OfN/yYZk6FnmIuHAH348nNXkd7jNVTLl9M07vKxwDvEVWkmYRAQna5cz59
/8jP2dazeXoKSfCU//ZmRKYfaCjDZElyL8QrfagpfxQQyTRviHJKUbzfHu8GD1PP
NhHBIbK2wluBC57cbN0w7FOdYo0Hx6AxQcP72e96flCgsxldbI8/70YNjdVkWD4c
PYsm/rLxHOGoFWs/XNJXjYfJZj89T/q4k9jD3s9uA3AzOEmwe+89SXgy1oAgcgql
JINUaK4FIsAtA5unXsyGIeo9VIYNcn61FpeKycnCNJJoocgWmBeVvgl8CBLPQt+6
XXQxcxdU7deppl3BUzLwZUjUslKbU0e8WK5PdXmJLYmKX966lHnOAZ83oChKhiar
oGkS3X/69QvxCXYOxoTs6NcmnLHUTE13KJNCGSHGww8G1Sy7uQl9nJaicQJYhoRA
20mbkIHIIVPIJB4dH7H4VSDii1/nKsU0v0rFasplCFdAIHFVTd5Qu6j46tC/IJ8v
5s6SfPGoqV9EVUMsPjPRpa3or6PZEqclgD7pFf2GPAEHm56VZJ+TKn6AmsMGbRRR
GJ1EXpZcltn201O8gDq8s5kK0FfwsiAiKY817QN9Hhm0b1ZF6VeDaGdA3ZZOg2Sb
jCtly/kG7E72Xk/NUmnJ7MF25IZ9xDztugb+sw6Qs2f4RcqfmZ/pRhleHClQxRuS
oBPvQBgF1VPHtFmDsoqpztn9474eVPKLNqDqwozsE4ntgDW0SqKDHhe0/+dgpWt7
kZmC//4ngHVPItJwkTX5+CgrlA9s2Vqaq+ByoH1fvzPAIXPXFHqI5QVMMy7R2UjT
cRVy8wOioruIYfh7kbMbaLtTKrpvMoGdTHspGi9/QS7PQQ1iW9WhbO845ooCjqtN
mEvE8c6B83MPoNOu6DrwbmAVGbSMbCAaNrcJK+YUNZ1YnlzR1uJCHIyxQWR93Npf
6lThEiL94YJksoSuuZAVelKQrBlmw+11EAXY7N5V/CZGp//RgzTDlwOLbG3+lqae
Skuvey3rut3GWSBX7CX365UO7G2iBKGYrKGXdR4leYXS8CaPXYTy7BnDFyEUQ8o0
5+HHxNqp+W1G1GwpTbghRPuJLlc4K4TlQnXlZBh9od+3FosWq43IS4mg2kVkapkO
ALtrvhtBA81ilqiBaArBwHTRaE32Wkf2Kr7CMhuwnSCzdCCpRnYrh8YnnGD4WTSG
oWynD1l/fF+rtroIt8q14cF4CECNOHRL4ieWlaSM5JsiFNRcTqQH/3iuLZ2L6vTI
cEO8eXC7Q1HPHynxaNm+f1DPfQ9P3ha/8qn4FTIvBzFeyL6mx1kK8rk3RL14DLJI
uyZYO+y5OqrttgjSNnzCmbVot5RvhP0d/0tmhA0VYMHvnSrkelhMmhAD7umfhN7c
rw+jB1Mm8sMGs+1Wy+RGM9hW+NeYs1+rE5EOwCPqYh3Ffmv0PYt2l8iTWLR4MwQ1
rghEI9SLFKknG99vOqreuHgx1Qtcz6GyfT58f/GxHbmSCIGtv2rhqiH7MzGoAodC
5jVKYec/exWG5Zg5YdPy6fssvtX/rNZZZH0TpeROn4l9i2Hc/bQvKZMFKFVXIBs/
q+PTl06IO356Yhrtlv5UwRRAetCEsLU3RgUuHhPOd27/drGXUEVyTyQbvL9VjKdc
ecvrX+ZFQZz+/LjhdyKpJMlJ+3b/hDad7iCu/ZXHHwqJadTuawM3v/nvSf6BFB62
flnjo6RD60V55MAkMcrKGBwGphOnP1zmre6a00cmsOnWKSDTGiM4Z1GObaliulyZ
1B+/+pkupSk6OcgX2VRw98P7q2WtmAMDblh1eJqDqeU1gXriAFn5vCpTIpIGKyAH
n49XDBQWedxkh1p1tabQzFqNZYxBqLG5D7A8g5Pz5fHcX0phFcz/CxygxdwpEmgQ
m5K41abhq8ROb0wVWXmEmrMoel65CFP+UHIaZD2qevWj5szYwzWX9wi3KqOkm/FK
Unzzie495f7p4dgiXXBvom24iBn5HVY3mev3GY+mki61eaQfWq1KF4y7V30tBkte
3QEsf1dg4GzBVqZzZdbe5MJzI14lKqV8IMivzeYFPJNMACLc4koK15u/sllbl8dS
TKSoBGOxFgraNMfCT76Kz4qIDmyUMTmrQX3iuD/otFzdOaOKqDN7k5GPupXWoG1a
sHIp4qtRRzyUTNCJscFVMfNG2fc7NGf9iX5cNzsoCH1rZU02oqN9vmUFb5nxagOt
sLfjvrw9FmEV8h26ja1gy6DWRy3I3gtSul3fBjvr4S4ZZ4fM9A4A0JiRbttotyR0
DjRFNEgS6Dr4tbWMWzkQUnAGQBdZkYXs5arQ7VJaJQawRVAHxv9zA8ioKvit9toO
XjzQ0qXg3Mi/FrKp6D+OsLXJoS1bda0KdcuYhu6gq8Xn/T/6cdWkWZXPjeMrBJOe
B2vPwdxk/BJ1/byThigPP6icQL9UP+R9005pabJeQSdghB6IMbgkKrL9kV6mFlwL
Au7M0zRKuyd0XkERFN1eD0Y6DmVye2zekfl8tn+13yoh5/mpXIpGarkPloOq8Ic6
EZyHotcMut1rxrCMecQ0FeZ07NVgKY/TmM9htIUhrPDebc7YPKIdSrLpQVafsG7m
YO0rFdbYmBXZ1gG6zBZHoXyQzt2VRlD7B6wWjYdFpHnOQ8iI3FPn/Q4No4t05m7P
/73WSOA27zfMC0OsyRiTq/V4sYrYvEKpGmxdwT4XwSY/hVP2FNEP0uyCFFn5xxVd
CoR1HeR4bZJJxVpMF0W7WMVi1tuoQJwGYKHxt6PHijrJkJQDYxcKKYM/02zWKjkG
F7hmz8xWkbMYbMIpcow7dM85AwjKLB1D2ubNNCl9JfCg7DLF7xTS1HZPDm6uAmjl
petb7njBFJpRiJRjgkv1YiWKo6naMapgfBxEIrDQ9Y/cnljV3yvF0ezOCX+tZ7h9
kCApKKm17IT8212DjbdeIbmA0f7UEoQAW5P3O10zlywjTp4ltnLUBHC72c/hLWhR
WmC5ROcdaIqlObfU+5oO8w==
`protect end_protected