`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5408 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
XDmUU01KuyTGZ0KfD/yCUy0pnXIRTRHDFiiota/NTtlG4bzo6vmsilZXI0IM3j8P
oHkJALbaeJgKvCUn2NaeyJTz+v6xu1NJc6CloQQGWYFS/VQq2OPW+rC8vKCfySPI
bRJHUMYNdXaEWhdPC0M+yEefbiqjWhXrcQQDVDyRuayHD8aCqPWAmtS7YzIyLtXb
oGBqyCoVMJ43/cQr7azuCqHczLU84K/2rw2M3FjhJO0B9Xj32sj1KZYuEDf246Z7
9xqxb744JE0z2W1qO49j4QcuHjUyaqrtaVvyVmj2ZlU5MQHIxFFj+Zeo7XYQfTwP
z3hgMFEVXPUfxT5eJpwyKdQEq/D+o8oXF3H/s75wKKGF9w7V+RNmsFMSnXG1h5ft
pEppabEhB7Bh/3O36qzvFkj1bqJnios4zPF2R8AF64BmUQBhSw7iTGEs4r/HziLy
9nh3HguZLo6UsEjGe4qf7k0sf6O4QP08Gun2xR03tBXxnbdyZUqh7r+LWvRi3Pzm
AIXajbPoLrF58rE8O+0upOvjTrC/V+CVh7UBgezGxmfkmhw8c8pGb12kNuFyUS2f
ogXOl5EjGgMa6C4aYsM3ezlZIm8fCBKODWouEUYfBfOueT5uG7u70ImqQz+RsmY8
h4Yqit0k15aKnMrOUnGOzJV4kD7mQEqf2a8uEQbqg3TWds65uN6MCBxcnlpIy8aN
6WQf3fZBeuLL0EGA/7eeRQZkkvj85EQEoM/M38SvhKb54O2RXGVTYD1866oMI+kN
mCfzk5/drJ1NXoXqPhBUX4xPWqpA2UtfYt5qnaFy+hKsFqzi7lWlklxAqelDgBKw
F4wxaJnRpMUqP/OJ0S2N69eZxYieG2geTqZSG1gYao+x2HdUKwm47QWlinPkMotY
AhdUTD+ACR2ZlOeZwH3p3SJSCSnYG4HDgwr948fvp3PJZRWedySzDtBjgGxcsZI7
owxbW+pSzlf+gsqLpNrg/yWOhM/X/SKSj3NL5srietc44ToJTEsjcFNRHjznyOb+
Ut3dl60FUnb1Mo8W5ZIi1rX88aCflEWPpELZfZ2v8IP3P8LX/oZ/oWECTJGuy0uX
IE1LwTQb71wOj8CVx2MsF49PbJfXnSKwkbUofdZP+bDtIAkSW3qva9zvasmSWRN0
/7rMwLFFTp+MIfhpqVPGUKkA9WKRWSEHdFglS2+9BzQqHdh1LGDyHgFcwrKWvExP
+VJHCC9HQQkzyEzoPNePIr8XE3miXYjS9TDpxQQIN29KpYIjbEUwos2VPGVoRppd
A2BHLJ2hu/TfQ88IScgdNX6aAMBkmNYgNgqXKfjdKux0VBmC4Utm6qvS1bwJ9LuD
U35JhFR4Yop1PZ3OZNZglOM9UewhKb22I8dEp6M+JJ+T2TIej0z0u6NaxP4PsZsq
I1+kN03PUB3igQfbNdjarl18+agWAn9VoDdF/JsMSthKxtRVYkqhnyQLu2YFGmhm
2qtIKnuLC06OBgXE2qa65oQ6nSD+l3mBgyvVZGPNHcw9+nxtekGsuR7ax9gjjRf5
C3b6EJ/3BY/pO+rgNNY3na62KzwQTUL3ivPWfEnG5AMIbKsq9L1HcfKWeC0fgQvQ
KJlX3uyZ55QViPKZ/Yb6H9rO8Ez9wVKH7fT3okqynqbTmFXmwxKptBq5V9pqOuFu
wEDQxuuxX04Hmj57WmLnSJ3V3oMyK/c/o6CxDm/TwHs8vR8qeZNECNFUXoAz/Tvu
nW+THMViTp+b/MVKFwa0VSrt6LphsrZAbDS2fU5zBYQrz4tSHBLM5UYlhSDJNRcA
ZPKLqdgDTjfzIPQASGjVmYO9l6Qm1bt5YzwfHBnW1Q+bVl0H5NrG0/FxDoPbVQpT
o82CjvtUZZvptE89GWWyVP8PzwL0GxXy6UJ/o54pi596lX0ueDmzlSeXh3DelTaa
w3Yx4dQhhd4HQY+Zyoy2ua4ymkNtxsoopUT3DgB2jtUPXP4K/T/uMRzrH7NbV93p
JtY8fw21vQMXm1BYtwwFPKCKokjIqpVPNhaPLgR0tsDX5yiewliPd/J5FRq9u+cW
wGobrdGXlESzhXWn+XrxyC5F4gc0HOypo6ujTXcNsOqZSf+P72yAVASxOQgMuY3c
j9DS4/pg2hH1LSsvQY/mNJmrRmcr6OXY/ZI+BP1awqRvYAzYLIM8vet5IKjaigKk
WdtcNAigc16rAhzrHK5xv+f3lujOXZvKUNysy/Mo3pij+ijzOA9UuwIGySD2xwV0
PM1LLwBEbkmZ+B5Z+CWdWyBa2qvYR9at/e++4CeB9LiSHzUcv2/sAaP1ubFh4nAM
aQtTfk0iRbn1jImyBoJoNxIgtC8vTxlPFk9nMaEj+2c/Gb1t0m/EkuwVX1SQkdY0
FA7v+zMtB1Fzzmj2ffSBvJqMhsTIThoX2MpIhoByTHzED+V3vQIY8AMHi9gEDyua
/98S8aXalsIrpqs7dTC1iLpr5K5198e+97Ejw4R2quEj7hpiLT5I8WeQybiOjiKV
fI14D9TxhLmuU1D+iyUpUPYEJRMZIbu5mNDS6470Sjl6Unj1zkIAnNvXdLgKEYB7
oou8bzJkB30eMc7eT3a+aM/6vqobTyFaqWAuDk1OsJAw6AFQsUEKFVEOxUSJupJR
sWIoiEl7Hgsyz1Wp6Wlnj6q1ZTnw9dyvcKc79BdyCIqlZccBpMhQvJmtU1+WqS30
IwYvCv9/U+rFczudKmf2I5q19/2Q3szwT7ecW0EILcNlI5TB0BKOz4EB+6yZ9kFm
tm6SOwSweZtN8+bDjodYH5VV9buVMBn8W+Z9jWPP7RidTXMF7GZlRVZ113rgwsFo
P39Sn4nBFfcCV9o2Eo2Mn/P4RxRBkI18OAMWkQg7Nb+a0rcqlm4Hfuw/sP0tb0F6
2yGpK4dP29oWG2rV1L1KkeYxb7vGJdCD+C02TVDl6brNVgr4POp9EO4P7FRg/0W7
BvTjpdQ8qyHEzzGzICKVaIsd17b3vyzYNmYIhg5bIFpRTqycx2fip2UjhdNPI+4T
ggwAO3pCleKcTjiVnVz23hcb0LpLRw2SG0oYFGW64mtE8tqVsir17LIZ9iuA36qK
v38H/s+yXpdvPyXoEeGcaeP/miZNwK1UAh+MWuIEjV5ZB+IxtvbVQ7gN2fvA4V6l
VbqQvOAMQoLOl7WOk3fXmQ7oN89X9jlCSZlCcXql0ZP8Cm0l6UMTY5Wx7CSZcVn5
hhpEBqltvPv7fSw8iNwYiWO4DEj+js5BM/YSqKBQJN38eEyiJrSa8qIdu4Nerk3Z
ox59rqpuEGtEBhDJRKBJejo9DCpQrb7/P4A6kWJNoTOcCWSCq9yLIY01+8IaLWkk
Oo1ZVmFvKEPJJO3O9bquAhyMUOjHXsDV1JGBZCe0o58TlKAv03ZfDZbbm+A2Pe4Q
Zoje+92abzKgY83l0rpLdiP69QtU7C7OtolubtSAa0xiQ0xqb4ZdzMQYociRkJuS
+YfzcRsK68TcCUWKqf9icPbQ5czjVw/LVP6PL30xSOZSnUdCIG+W2ea52WejmBSa
vFmem3bTeZxka6BCkmps/8AyyYfbMdYJYVk8Ki2V3wRqzRn2561T+OntFa7HWN0t
2p/4L4ZmuP2/PeU0SWJuLswxZVyvUMZXjcWPnYSDSpD2JZDAW0wyY+Ms1glNtMHe
9+21/WmQEYHf5+DIRQnVtHK44KAqDapnhgGhinFKB5k8sGE44K1x1pizboAZlQRI
Mi2+pPcQxIo1maeVJIguPwr6+ZI0K9XXjiX1M5xBD2LHrQNafYgsZRxyBCj/oifO
ssp74p74+7Le7VcSUpmdrQ4dvxO9GzrsddNRJSCS7Qdzw0xOR+ABMCr61bZarqbL
ILWCD034VwUx+DwA+qx0Vop6AzCgiOX/L+vqtX1uPlJL3rrRcWMmRLCjQxiSK7+q
IfRgtiQ1Id1q+EHP3M9FKAJuVrcJh/+UUXbkvfjL9It2VxH8YgT91S24YsOOS+dJ
ai32+i17H1PWD2YrHiCYQK+qZ4OXJgJamBFz42DFVyHm3Qpv5cmZpx8KnvtUomqz
JyJf2Eb1bDVfNlIPopFPPUb95vX2/SQDQ2Q/i/vLjiwtLjHYPvy0OplrwUvXxNWb
CG1icoLU9Uy9nOP+cQMR/L8ExGrMDDzJdSz3xBQpPpTeqeySILq1YIktoZ1CoSIB
DPBV+srbR5rjfRZS16WqtTCG6cuxW5yqUani+lHnR609CFXroLgG2g8XInXLO4s5
vfo3B6Jx//1VmusZodoNvY9BeR131y3NtMRmARDblTHkX05qh5BX71n8UU0WSY9l
iDpbkdkMaVEBK67Dt7GSRH5eQN7w5YWWmBuXzvy4G/jXv6g4B6oF0cizWbg35Oer
VinK2Br8mgUSTmc1SIQjHTf32SStJFl3sDlZAprth+rshtMuWzEobsZzSIGmwbhF
wm4NyohQ1BnZTmczq/cjMIkWmE3Ngdx3dMshvbZzJxeBhBtYIiHbgYTXHZnSOyIF
5gqEl6gJ86wfyJpWPy0tx996J4Kjf+KmNPgq/+FCXJ1VuiJ8rmz8qDy0zwYYZ6tz
toIsUA/+bpO1qH+WbpNFmuZXna5lfR4sTmT+7w7T41sPNsSlBaNupP0bqEK8rHrd
oc6wvNB4aY8EEkq/RPMqrvxQ+VUsJjPfnNesJx3XKx8rf18DaFGetkQWgHAvF8+P
rFyf2yY6qsvvyCTAg72f2Zvn/4d9ka3fO473poW/WoOctM3NMG3Tnz/y3xA7a0hw
w84kakfbXSgq+nsG3xuZUVdHDnBkJKOPowc2zqmJ3hJEZ+YT8SYj6dCn0ozhXp4F
LyMu47hsLsglzxkrkMieFXsN03o2HQhzZN/V5szwUxLk8sKFIS4Fq9Rgdy3yeHYF
icLQs2BjLamH5TFIP7FpF+ZiCNAZuGm1Mo8l1/yaa9KZEmgvJLsX6+0ahYAStQnD
zqkopLNLgtnPVJ9w3P9w3B6YdNm28QA9CBwOjv+Moj5b/MHKz+YdcOtzE7mLeipv
1Ws4WvQg8UkUWcEA1uWttWvnTapTOTAKZADSuJSCEnZAWH0pjBtPdTcK497868km
gtb20mCKrKK8MtDLxGHiaHyaU3RsYZYmol2rscwqNXOUuPi8sbbZs2p63QsyOjgJ
l9CKb8CkgPwf0o9XJeNqvjmuCtRLXwWiJ86bV0TqJAv+/d69dwKdkDgi8wYk9ks4
PdDFi3OAyfBI52QSR7jKu4Z4E3rIg0VARRRX3yjBRa8uVX/yAgEfCz2+yFUtccUX
Ppb1adOhhLkFsQAd4+jn26iMMRGIUjiqUak7PsTSYt7XIPO0PojIAwX7spGAUA/2
ell2n4UVKyJUcUK9KLEreQjtHL85j+1jk2hQJSLwQNWlz/tUycnwRMnZN5d/ZqlZ
MSj/8tvfoobocchmDqVwabaPA5J8oWuwGgPgKU1elNHgPtSZBFNDJtfLcTnRWkEe
Y+RwA0WoRVIU+dyZC0LMOa2pMunopTnizNSiQzOpggR+p6u2i1TwxhhAOXtVPwA2
m3NQ1MWGNoiGG3ZNthVNr93LteRGMJDSv6mSIWVuHpZnxU8ga6qrJR6BuMnQfLwi
/H4BeUObWsfQ5R7oryjM4THWIJXUoQf+wCONBsk75cg3tjI0NpS0M/9YMcr+/IV4
8ujgi5oS1iKhSK0g+anc/q9mS4zxTNh5iWY/Gbvwk23FGfqpkMgtfmpt1LC+l7Ck
9u/9hA3XcMcYj6/M9JgLsW9y/UrfOWvxbVqKs6HI0aM9GZYYOKtW3HYBw29kwjDQ
/+3T0hI7UFBBnJAGCqeBEwv4ZMPr+rNRUdSyeC9tupa9pP6TJ/r49yPIxVV5k9mT
F6KXL1m9W51tWNuaRqKpikDqIsoQQO7cILdEVk9HlvSIU0J4+r+uq9ux6rTzJN08
fdl/Q6QRaZjQE5NXCFzGI0esnY76dM3a6vSd/xX2ldnaTz5CPA1Lg3jKtaSztIxt
Hye/lrC/1tBFYsgJAeSLT2RXMjqqKMcgapjQBuuB3pzjLB4xYzC0Xb5tcO9ZTkg2
jMjCj8nePpWJ7EweBvugbFhSqmHiUtPQoRcy8vFj8zb9wpXeNqIgpmKiveSSfNfA
XtKwDaAvlG/tow6t9ny2Y6gl6pt7z4WiQeRw+gUQLHt69m8yasS4ie2pcLKum/8s
j/1eBmvHaOwr7ayZyw+jSa5gMAqLquWP91A3wnbaOIdyJVFJYVVMZW0qGflrU/U4
bYzOL8/xtbBFeTzz9iGCD8cuR5J4FWco2AoFBmepSvMoU0BaE1LcQbpdGxzIUB3y
y8v5NsdQC80ED7S7R2sz7lbbEWs5hDeSmExtxLS6uWGne6r83q0nq7LjpoM2E24f
47N1kQK2Gh8TcfD3FtHCU6RQWChKy88+aVZt8cxhtTq+CAIwSPJdjB2geXMOv1x7
58wDdJy4AdcFvatdbrfRqdkM9hEV3rolS97A/+D7aud/vUNC/q3NPviPkhzcgIYy
7bidbj0SylgW5Y0RKBLt9zYvE0HIGeBkw+JEJE6VWq7BLSfqjOnL3Rftos10dFW7
HI2SlkHjRmY28hYJ7WfESUK3im23pAqDg33uFZehhVcF14JPZqqMVSv0JLNDbDzq
22iFkrveYifnRqcOXK1l04OM+BCoJSVCXhalzoptUWqi3PVTalKvpAqg02B8TIkG
Fxdpa6tasbvT95+Mzw6Iusm2CfWAxxUwl8I6WHDrEZ41RMoazUdXDFvrjvke2zKe
q8t7GI8O9RD55lXvdw1Vx4quno0z278aPKF5OD6rRLoVyJVZpIMSEDGWR5fzwA2H
YmBxtgiKCQzBYHOe0CNVqFBtTzKfVXlPioowIw5cWeGOARrzkOvTvcNM9+bqjyRj
duLouSLS4eRpMn5jdpX73bFBESoDIMHXTtJipHOlJwTKe3FFQbeFpBJqgqRe4YqG
BufOH6Ub6y2/MY6SJM1dmvqk8sWcqc0Oaxp9mNfO+oJJN/yFqMigVIhZyFVXAoKv
OnUIaNABQYNvh9NeicRNTU1KsMJMaB99dnSl1ZDEiduA9Jc+RrwW3d1Aipm4uZcD
oNvO86CtlLxhHssneZQb7FZ8HlSTKYLffIZU8kwNUSw=
`protect end_protected