`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 29664 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
/vEkqJfyK/81z5lf9X8oFQfajlHdKRylTyG5OjRjGcyOcNYr6aV7x1MeAUP8UOBz
5ZzjDHEuLjLU0yKFNz7jPhVjyJmTd3JfaJYHINqnqJvJGD2zDtrSyl86HQ6rRvAB
c3NH+unoYfu13+7tT9Ir1/rPhlW3PaB11qrb+ua5RhrZ58bzh+tj6Eni9ZhVVs+g
ibNIaHEX6KPKdKxkh0VxSBKVZbhpj2TIEzy7LcwUSCYWkQp3tlcdgjOvenM1p6Qv
zI3fD5TY78VfVnR1x9D039dtvspVK2O4fZeFO2I1hahOxHQCdjnoZYqgGIitYyXi
d8WbGgBt7pTNs01n+5ajk3g655T5yJuPYAwev/ULOuZ+wOfoc3o26NtwJsmX1T6R
0yt5oXMu6dw8gomPR11PnKkCL6cm0Vx5BQRxibY+lpkudIirZJ+fJVycr+6UiqbN
BJ9cObn6BrPkuQ/3ZuWMWoPbVSB/+5+MFEMGqLXIqeRjS4P5xk1Z7aIQ5CMQbPOb
WttiBCHVTJVB8SHbzmHREoRvY8auY8ebZg2IVoKu8bk7dhUpOPmPzdJlPqiNqDQ9
ATPyrfO7SKXPPoeWWpld3JclEw8+LbwVybcanVDiVS8wCU94IOqPDOdIdmd4Cqk3
+J77QueQxec59f8EGyUA655fYLRpdPxrqlh6SEYriXkup6VUXxYGAQ5eUTYaIoi7
f6bTO4D1prPqcZgNhcqc3MtIc4OddaZ91UQX6PA/b3q/HPTFbG9hxe2VhkVW2tw3
+dyCrN2/6VFdgfnYfiwQrD9j8YO8rhuSM+xDaz47o/OGTI8hd/S50SwoA9rjQL55
gJ2EYwXq+KaRhbG8oJDLQYyDhmKgFu5ekWtKyiC6oRAnUkwGsmtPGVu+72vkOW9C
jjqJyKbuTe5JOM4XzLkD//bvsGC1/C7SdZ8d8c0L9AC3vQ9pe6FO/V3CdBuExhy/
5VHGM8di6Hp5TQVnv0MpJZGQf7k/T0NSso7dz1gS4icBjQEN6EilWZ/7QGxi0ds1
ade+6Svp5WaRyeTwEeTU4xjh6eSePyU18ZhASrOlf/O+CAsirGlxrQLlBVRkHnjl
z89PpROIbaDqnZ5uW/5Pkg6N3/IyT6iebcBDdlV59tSftcspfaL6oLgX1jItC3Y1
LUKrbWRhijdEVKK0LaRBClZaK0/jzajhTZnsY4Zs2CivAtIzMN01AGJJ5EYl1w4U
ro/e3yPb1lFY+c94jeEIF7WQA75mKT4taNVzscejtPBbpJPt59N8ZjxUxZ7yOqOZ
k05LUYr/Txb7w9cbFVVuzU4aoc93jRznB+letk7SsztR6iekZKkCsxdBKsLi59EO
bMv2fxHzOj9wZuaOkzqgi6vt42thnbodG0hTn2o2ukkqGlDR0KTHwJdzHDN8FmKH
x4a8TncR3C2bgKVCVd7L09gFT8onPkwoyMGcIA3W5LXWMuf1ROROJeaf5jGwTwjl
iHRwvKslPgs56BXCODTkBnMBCp/QzT18xQsNJHTzhpkPFoI/S8NMxOSH5TOZVhXK
pS9Dcw0yWS3ZXRfwPeQiO+fkJb/UKeUx7anmwFLW225Ma1p4C3UbPCyM8J+BWuhH
xYAYqh4X2cZyr/+TdDAozcw0Cikmkx0pgRePKDY8DOIB0g42DbKLs/MjlRPhZaOw
8U5S7STa/7vZ5QjtSEO1itYFChAkkrtfq66okmF5j/Q487MaIYgF9LXa8CwC+AbB
oJVUCmWpr/8mSUGx4ViU7VZEF96f9IOlSMRPf+1uutghyUIllF18LaX4qdbFixry
ASoqN7sVa3LRh8l6EstLoDq1xQ+hIYIyTp1ydL+s3zcw4ERSnWC3pOtux+kE9fma
RdhucrTeKmLW5jXEGXdvQALRcVJ4GaNx2qvLHvXcpyItORpxDym3ZmciYfbSRpwj
SPZX5cxegRARDxrMpelE4nCJQUDfr1UV9oOkfQjHvIynGt62tilG8kfQ6oCRbm3Y
C+bjd4AUeAm9m5JbkqDE2RQ9N0sZNTtG0mbe6L673NhUx4Rsv/q1MBoEqZpK5Nds
2CqX7UDrekR2HdPiafiPMmXG69Q68vL9ENn6rnqEmWsawEc1SjFHe9BjjNpDGgc/
mWfBH1gTNXvqnPgpnAJMhGe+3OyQ1WHgU7lqsqQHpmT/dnMZUPgMAbZOdSG5AkP9
Jx/i9tf4NJjCWY1Nnu+/cYjtZ8QBNkYMsXq03aYKw1KY9cGAX34oMytfVAzrQELc
53qRvqKXQVJfSXct0YD1l9/UlbfgOcFgrYK6fB/qrVhbTWisNmRe1uKeGk6Y9LGg
YdYneYLiNOxkyLCgFo77EQQU5DHWtovdgUSGDkmdEbQCDq59PiYRNUOyCTqcymeC
pAQLM98ZHi63PKR9UIHEkzlKeEa6UWP984wcrsCCcx2/mL1maTjnCG89XeBFIhFf
4fkgtwj0WcSG7acbZA6KW8J4Pnk+U012qaP6flKla1oN3lMkmwrohg6q2IT0W3OP
lUDFJqxaFBlalnQIJAx4veCkiDs8nFB94Ifk0TkKLYNtxi1gx67cfDXkGejfSelR
z8M/Han35nCLxOpqYGu+TQ/GoiwOFa5JlS5c1pGpDLkLJvvZfomjVYJAx6YWm7QE
hliBLDWfJxQDLLvv0HOQf6LAlKhfz4koh3sVaYljf6InqcldwVraRxPVf+qKXTnG
98jYUe4CSuwi2YbrN2xqt+WsY9wUiPfw/4OXqZju0742f/CUCDgF43Q5BMy6KaO+
ODqg4MgplgZUHcHwg7UxyqImFeGR/mdHppYOMedCVc15hq55hZ+FrptDeGUEHJ4F
RwMYMaTkQgnFrK3LzlCq/28owSucFWHtua5QZcioSG9x7gXdi71vDPfIGsCLGqYV
dNnvVUF7RKP+UD59eTtF7IZtwXxjSX2P6tGSbnWu/wvuX5KmSMoFwSxoe6y0Hyos
24/rzN/7Tnt4YD+Ill0HZctQ+YFdGNeTWOu1B+2AhuF3NwoZRSw6T81eDoOklxw3
1TZsxkQfcFKSi9DJg11pTnVWyZ/F+CARIcsFREoq/G3jBRpYlNGeXIR1gnNM5H3p
p1fRtM0ckVM5QXOAnfQZ2bux7Qs63Ki6ecgE713BZXKGZwrAMc4eRVTd+CZ256zC
SrDeDC0iOEyTI2dhFbHFpg4SKUBJhuMKdYczZORo9PdVpvQiO70xEIhif6IzZs+F
iPPTZKTSWZjrNNjTAztB6cofnsESySs+Wew6trZLm0OK/T0vbIfuSSJCziGE5/dL
tKIKYgRbUj4kghRqxjErdef8oXSVHYWSZIPuGKLWKEalJWJvsToURrYP37s+G+wC
7vuzh7FsDHLapPGPMhAv6W29eJT6YgNZmUxgtN0sj/bHBnhOY7gba5CdS0w5mRjn
Y8DyljMmtE7qgvehQBD5e2zPfz2+kbccgop0DKn7YhC9dzHY/oMtQz8mfn7mfEy5
2D22NKJJjcF4B804x9MrHmvtNtdgxY9SsCrObGxl18cp/Bu8DzxhKi/wYGfemgMO
x2O/fE3RUBImeFPjeGpL/v4RpOsJigGx0uv/qyWdJPh08qYnrjO/rc0e7b3EMqm1
lstAnhtD3dJ+8HMkYHncriPN5vkyjissOnMFdtuWTzyU/LzX4zTq2cIYl6LORXRg
YKokhA5tHgBgq8LWAVToFOCQIKOAZt5Pnsha/qzgQzigfDINswsFxLBNZftbSGyv
EthFDfM6b9LWhTGUpvKpT+1vEKkR2VMVt+/LyByL2o8Ncxmm736JK3jlB9OhdLca
Rqz0lGafZpGAXR+Fozf8bR8QZolHGKCvA54O+2E0swLaL7Rc/q4G+KndnFIFO8XR
PqdXBt++sMcF4dRL+UpwuGRdQi2gAvRRBmYyod04DnoGS4vVVe5iCK5dgudxnF5z
hMxNnFlamOfwBPl9Yb0R/OtypLiWQlVpnDd86kY3LG2NJnrIxzsertIALHLSHpxN
X+ZCHsaZq4dX7R4R5yZZVPPD+szDwCtqoSlr4//S3Ljf6OzDt5le9+gytxhf2+7c
M9jxB84pnLmaXpktBw8a/d3j7dQxznIqsEjZGFdsY1CjMa9PFzYdC+I4VXHKTJoA
ECWCGZdGt2xuihxxtD33AemxsTr3cy4iFFVNpShNbbVAYAxYR0KrkwGVkhFkDTrs
oX8Gfd/YBtMf08zUQr2SSkDVLt3TesjuhZTMxEcpJyc69CTPEr2Kqf8+BE98oGBl
XZ6XclsnfRefgQq6B5KngAApNg8QQcgtSwav23DOWOpdnZ1bj0XeO6anSIjMoFLZ
x+umrvzDIsqyHnxnpDG7IbkS6Ota2HAPElYX3CEC9BWGDDVyChNXbw2eJTbA+5TT
eaVOtq504sLE9iImwQhX99WWwnOtLXu5pEOjG9Xvi7JPLoH5Xpiq81S8tUJOs6W+
itn58tA0I0mDRbema0ELncO29aMJTO8b3FjoBK427vr3WdPEMQUxIOMkCSU0GG8o
bJ1R2qyAX455cPniKnjpd+7+No5T+zdYCe/Ci16R57e/vfWyptzEZWCwuFKL8XDT
S9mTCox0KDrDFBMxmPiRP+sTU+9EDzw7oOkMhjTt7bdGTeBjDNTzWj3NzMKgLkTP
+NgPbD3SQtRgxlLaOCGTWPVS+UH4FiV2DZvjkItZf/4D0xoPmfd/OzHM4o4sIz6B
kv0PvIR517xnH+BUrcWpr0GAmjaBmpi5Npi4n0zlUVLyOjLiKQh5NivofOCtiVMK
xW8iJ2WqjkHQ4jlz94Ox8pesSXw48mjdXMJJAcGjWkE/L3B7nHBwir1e0EhS5lFQ
oZQLctHppiPCm5ZgaG9Pm7Ao3udxCVneCF9qiGESEgLt/y9ERE7n2wiZTir4bTPC
CDlTA4P59BxMHzynSCgLUOXk7dw+KUK2gP/M5sszzoc+gwNns7iouxtu/pUy/bqr
6HCAQmfTJbp4pXGjMSGezfSfSUO1KrzXbd7czUn8JoIV4ra0aqYYveAoQKYordnu
aduk9u95HDsO9SXR22DXUBzhD00GVnPdU4/DkVveHctHRQ5LYAFsUl0g1NapcQvs
lh0iMPk9a1WLU0WUHZ66ZHKx22DDhYTvPRO5kA37ZDpj+L1Fue3Y3V3VjlAzo1Is
ylV+5nGiEB54xGgPfwRrBun6ThH+uNO97Z9G/ilzf3++nLulTBb6+w1rS+KSKu5R
yLO9deLMjrQoGSBrmWy7ZPLNXZIwgyEH/4K/Bg8jwHLyMVIt10PCHXJJGFqQchal
2aTDTh+zwpCFvurNoTZ6vrtGuTfb+k5RPmX2258sLiBwlB26UENM9/uYrCJkEXbf
7jo20LYpgc7Ns3XwKrkgWvfL73Qdr7vJkW3FkoRfoEn1Z9VukE3Vf19wbwg9fcfX
+ifwGdPd1GHb6oD8feUG4TpnvQIerTq5ERwggABONBGdHP4PSo0bf2EJ5A04XXPc
2uMyOvXvoMS3PG8mAy4yQbgxS/Q7RuH2wh0fNykLN1hV40cmYOsMQzOc01vWUw0E
n6SFWxPeXj/IolhWebuZZ0wCfOE/YZNCIAjBPfMF/4mKHFIXqogjmIog+X/802Da
EI6ATQxKozsFdbxadaaG9w9371j5bv9fRxtuLK1OaAdhFMEGh2Oozs0Dw1HC5l2o
yEjXtuvK8qF6aJNWLCQCLxbORkVo1MLTbnqAELGsgSjyBNB+zrTNy3Yn2S4490gO
cTHJi/mT3g2wsSQZ+ue3rDV5Vu331zqpV5R38AXfEXFVkdUXeJRiglnLgNooZbKN
clL1ZxNtbW2E25WUnHipDFAalzapM1E02AFkL5DXzg1myLAw6u1iMseU+7PEtt00
jb2euIMczW9xOLSBnVI4LVYPCVrgkm4Hhtq8nfu3iJBZ7M04doDDvi398gaphg3e
1Lzg+XNHvSiHjKsBD+rlYAyIpLBRBENIOLyVR2vgE8k7qdeZIvLbnm61EZJfR4xS
liaJ/RM57M0jqMs8aOIBR9T9SBTO0F2yO+B5YSpp3omRpw01aO72fQHHxjHioV5r
pS0lrfdynWmIo+9essluDZSagsdC7ReyKdk6MaFlOLorzYBCJaOw1hB6/m0UEhfG
Q5msSM1TwfJoqLVluRJZboQUMD2Ttxd8FS3cAcRzx7ZGW9fcESQE1fLijDKnN/s5
FAEZua3E12bfZlym650FJzaw1N16cG92spYfJntZSfE6iB9gnNCw528BIDBcMTvo
hsx+n8QY6znFkrsCcOUmhMy95MZz4eqMFRLd4YNjIzDGAnoEgIsFKsnZ2bYeB2I0
8OuhJ9qO2FWTcbxNZchAfilXZWz5XPdlTBa4bAKDvlLr+JS9iml65KD0BCDNQRJx
GoLAP6XtWd9isdahIKVu9KL4c0YoZKGYcTMgee+1YpLQliT2kN1geB71CqTuz4Xl
mlWydhvB5dq10t7wFGmkO/C/0dQsZNBY/7HvgbAsF480UUfAC7HLP84Bp/gO0qHx
XZHzct4YSLhEj2NFRSRGx4C4hDmILRMgYiXEPmkYxcRQJGfr7huNNofDGXujUQlb
HUbjEzcNDnsRITYgWdCYCosKscKVx37qyF+IfHVU26C4mDUBeDcsdHBvyjDHOwR6
eGx4pBKf/vHCr81rHZz8l8Pz59Is83XxvBHk/JKYbrMSXaTWcClhS6rz/bJrFtP7
YfW3EfEctGir1FgIGSl6DKUeEBq0gcWoeyqihUqZmTgkTWZMl6mjDQaHJY2AFo8p
luHIx1pbq2/J5toJe7CXsGxuzJdAfh6jMi/SB96KJjlRKLIcjCPJmwZQmoTS1wpK
l7lc1RfnIO9EVmnP5UocEA4PX7TnoNTcUhfzLP40aCFcUpYYNQSn+FWEfQUrCFCY
rvgSVOjNSNp7vK5w/bMDXJyVyoe705GejHN9/cS/DoUymqxjvu3+T3leXHe5Z6EA
G3hF7LdkCFZEJk+m01M7gIJaH8b/4k+zVJXDDIXXoBrrkqVY5L/+HxvaUzyNdik0
wlVPkHD2WwSbvjKySOFTBOVzfU+aNPw/mm3g3Pcu03iE4foRUBUB4695bm8B6uai
f1z/NMiygP+2CYdYMemg/dMFO7qEovSAs2NXFe6S0MQD4SoSe6407hMmDnWQ6vUk
5MbRX2+qIewGydrgAGqR0t342JexAP94/88t6nHdwL9ENEiokz7alMlJTodaRb07
xK/oQxBoZtAqgjzTaCK/XBWxLEhoNUuhDfIJHbtLpSzPGxu7KU1MAnkfttrAuPS5
1I4rwYzCOQF5uI5juqXCmE3I/yWE3gSeqmzSoKewhnZU5nE4rmf15Y0cWJje2qP2
w2bua3vVvG+vKfm6TJ/pQ1FU2JKpGEQrDh5WFXUYkyhWNrJFQtXTQEmqUn8IrT3h
1hVX/E9SWb7kKT+KJAw1/LRKGRguRXtr0FP2wJtTJbZOA7wh8nrzwD5cdCtodKf/
45kepdyFSmDUei9cytKehcBevQJUnto+vzlILimkHHNvQhDJMPParlqMPfJGVxQO
Nd7t/US8bF45qf9ZRPIC3t9n9AdMvKbYnRxKLvdDaB4lyEWMXxWGGcObv/m/isi4
dJiKJL9bvG/5ClgVojWCBm3eJzR/SLk1i1wq/vHnpX6FWtOa0JA9yjfsHuQ5Xzi6
Rsie0z1XaLVcH78eNg1SEf6xt+2ye4PtonuHNJczNUJfS5reZAlqBpNGYP5a+P4b
LJg3SSqIKliQ4QDHbWC8P+dw0Sb+tzLcneVzt5l/DgDmfKFjmhXFxtRU2sSP80QV
LJXB6YqwlKqMusM2eG3P4d3oWW+LyZpg2U4oCc8qDSjgVjpld8vz/HRpPW9tdZOO
EAE51T1HHeiVtklc0pYFj5NbmPTOfz2fI8jDTTeqC6Wj/aPf67mRnGrNrDNwSrjA
yMFGbkiMom4Wd+NKcCuvgqm2XRSVaiwNkfJenJFv+FR0A3UVlcyx8JIt/xuB8gHj
kMd3i19Ft7Zse0Xcd4kO9kUl6KpyDMkbabUZLY8G031JzJzadnzu4ZQWlIPrxMwL
uqTix2bPOEqLRSr9PrRAiB4r3IiRd4G2H44fmVOZkYOf/5hWq/VhSOAuoxwu3pQE
gwFNvCVl5hJSz8au8FsEj+cYfxOpbfANpH8o+BS5YLHu2FLfAvvZcsFZvBdEJJE3
DBR3T14ZFBY6t5wt/lCSLFYIJDA9G/aU4SbToNA8orOAeOnqZl6u/vfVs5RXobPr
eDVO5jkDG+IThFnjEHE3+60/RRr8+iXRAxPEGhDF5RkHG5HtnhXiK4SUAr9Jt3OZ
nr4A4N37ZJRw0H/0K92Ag2N20X7vWCbwjeEEZZWuaCMiRNhZFgWilB1QF7T3yMST
7s80Wi0BvSwmheisB/CRg/OCwDePuOitEdW7xUSHyIcvRHElTM7Zbz/lYIsOed/B
nu7MtU6uNesLuZHKfrME6SW3HyThYcaVc5d9MOiA5WXzQ6TsvSueujIuR/G0bw8j
wzvmpEd/UvkHhwlKnnkaIXBeZIMVL/1DJR1QAejO9aYXFn9VHE3l4byQ9A41z1MJ
mNVVzLXE7brAwlcGr+Rwim1BaMUTDsdM+AHIcdxWK5oI6GAvG71tvbdCw86jtuIy
QnHIrRT9K5gZPhTtDZBTlzkK+3G7zVZHpuK6or54xYCJyWkzFdkiCWynhvR4DI3e
cviSO18F2RY2v31aUEieDAKahA4L4Fw4RfHqaCX6H5CvqhNINrcr6ncfdC9Klu71
g9eLiug4wXLGU/anWa18FqqJZqI1iNixeiw2kFBVEVy4f3CKEoc7xQ527ed9oLLT
E5Sl9zJsvPx1JEVNNKegdVcv/Jqu/8LDXNN//BpC814eqQc0zClWLomX87haLXqX
QJ8t9NzBPr9qOGUv+BTHxm1wuXniVzgjulGh7RnS23ZIL7GBgxBMxa7VDed7ek7y
nhQCDMHJCIe+LTQBLZIydFIe3xvh7GDTDe+Ug0PB6ApTd/0FxMGf9grMMil2He1i
xt6lPLEjZbrdyWtB5JsJk+99RGIdMzLOd/jDMk/KE8b9KhrWfGLUGHDNzui15gan
/4TUgrfrawZmZvSloLNA6mNXbnEZSJQ4oiSBE6NC9kSo50MRMADFzE5BV146OhVm
aXpryZ2mR+CHUc2dQvkHMTOk/0kaGEgNgeE5bqDF+zdqtltTFiDsC1Uu2wMivMjb
LP0E2zYtyX1hzhZi5RnVsE1nqSItX+rN89AtmgEpiCzquqM5ajErsd9taHIuDzf2
0ro0hSiCn/z/+2Ab/9rJdfwZbau/eVBSUsx2kPqzQvoPP+tdPCTitY2JzDUFJPql
pHMRb7IdYxiXiACB2OEaqZDhSSuAUm75mJf+sEv1aaE1vi54FT/QGKaLLk27eJLa
WlAps2VRPf8uFIpvEPayyxsOK2faxAakYhJDgLRUayoyqyxe4g9z9Po90rWFDYq0
tGDrRR3le78/h3gMHvJdVPiHsIT70GEsroU2Kb9EKbuB4dTgMG4sa9cifGDtrZGs
0QqsgGqtW4JNptjrGieMihjcMhWwf9euiOOYhC9Fl9GQFkRGgSd661yE3s8wUhwE
Fi7PnfKRhwGypMgavGU/j6SgLKpzuO6rIIIrbq7oqVW5VxRFnvpqjR1wfzBGH7Dj
5Nr1V0+3MbPDP6IZpLT0W68Y4fQd5rTXm+9eVrr1sh+hHHkf3mtgyLxJLc622kxy
72ZxWMmXeINfbvEiDohkHUAuTVjonch746pEx6lkfUzgx9KEWt7dOhvM8Tej1dVh
3ITBksNkibbwSMPh2XrmpEOJ/APnGSQMzx5ntUZc5HTmVdUoQ4TdzWxfzGylcWTb
4whkgu4hMNfw6enhcZjS+lc7GYhPnibj7wiHRev909nxWwcK0bD57J8pAf/gnwtZ
dqPgaF0TuD0IJkUgvDnAlvlw/bUf0IPVmgFY/fn0jUkS2dJhRV5CjByqKqwURdVT
cGSE3FS9jTQkjXLD9/KYZbfL8NSKkKDUMK12j0i0wgQGWB8K5DPHCULlSzecJHbZ
f3/PYKfH0J/gf7kcI63Lo2i+iNCKcxfs9n/pfdhfn9DGyNnf1TskTTN/LwMDT1ru
axxF2X12RO772Izo8oSxiKeEdtHyUOExJGuszm6Bx8qgCOQWBWnMX5oOjuuyLkV6
nf9njrW57vVaBBJ1wZFyeMP3r4yclnXH9LxC3lERd6WBexLwwqQXLbLY1tiA9UR9
dnxZ8gLjXut7GPIKifvGPA+D374WQeF/rP0vr1WmM1N4Z+sSERKPITDQrWGRwGok
iYNu4zcQLrfT9/rQ0fp2i4JJTkr5m77VB2vbMMkgJFz1pdN7QhOKsnj2QjyCu1vT
+nMchCyjBnvX4uXbhsnUxTGRKoWayCMbRsm8uY9yQZ5aTiffPxocTa7PuXQWGKk2
v2aflDteAz5TgIuF2Rhbd1T+PkL30zcKjLebcS+Vi7THtzVvVDCEM3B3s2Pi/gpu
Argtczy9f6WIOJQEOLEZ+8s1dgdhtu2aI+zXp84CfRhaeUfpCbcMrcMGqWJVkqCX
lShaAhDKBr+wZsivNRD4crSSAbjgQFz+C2aErL+qHzb/pgO86RVnBSJetP7ATPaq
OJUOoFUjb+JrsY1Jl3V5Nwd9KO9ZTVW88C2NyUH0THsmzLh6SJ0VMS32GBlSE1IN
Ij1czlRZ0ExlCY4um1Yc9AO1s45+RZO+oaSXmxKGyIRR0UpW61+pxgrGlBScWdb3
N/XA9oOrAILc0QcO4RO/Qy8ggS9xdssaXVpB/y5hV9iBwnOzmrtbhjCh2F+kLJOv
jRfx4BKTCvuh5QNEA/VUPQZ4lXzJX3QxSq0pXEYK/r7eBQYC5S/9dmDOkTcR++x3
26d3aV1BojhRmWXVV1N8gb+snqg6c3HaHNslKCd842oA/FBcTfnsl03HgnCFo7E2
0yPff/PNE4hp7Y+tgPmZfxlupFpeRb3ACRyUZynnl3eeJRO+jWhuM+EZ4vl+gssV
DgLTl0qq/BJxxI8ppPasrLsqVVpFC2lznAhA/sZPU+GDyE31tNUCB6t03Klx9DjK
zlWp/xcs5i1sr598rrvLKeLVztLtsAtxZG50W/eZ4ztE8iwVQtGE7d9bPl0kOVr+
pYvBQPVNbMySwmtPHoulFbuSEOPODLA+axFwDUcO5f3fN5WHYZCS5uKzCEjGm2c5
onRkspZg/ppBPoSoA3knCFGab5gjxuD+doVBeaeFUZDsiqcBjoQrgpt/rNX1vuQ3
0K/t8naFPKeuVnhJVTU8S10o1OgNlx+kSblLbwkrCpqwwc+qypxv5awWUDp+oIBd
pal3sivPf5zpIaCzZYNPuxb2e2dotS4pZy7ugwziMgLQ2KBM6CNHq0Eb4fSgCk1g
MpwP/s2uMbO2FlItChIVyuDN1ErdbeyLmG12r1GRlW6zMxEEBiSpbQ4URoW+Qke4
xE0UqdOOqyxu3RP1txf8VGnhCKPub/0hV+xxiMX1o5jY9eQ0WxtjUv/NqSt0JU8f
VW5dweVn5gFJGOJ8GCSTU74tD4U38vmR4OeYb9Mh04B4w6XEKQVJoriGtGhbH939
pbKWXVvJpTP9t6+skuAXeQUXe89BGCOIBXW5nY26mE+PCaHk6KVbpLADakTyrrJq
s2y4wupCZPO1V8ZRsOjESjqPOAEvdL9Geg9lO2ZIoXTNphXdgaQgz4wtvKwdHXMK
Uws+l6IZp6ZOciwiBxA4xdKFUtp18y8z8IVd8PPtosD7lQAVZjCQZ5JmW7/uYBhe
FUE5a7k5TNiO1C0i+xMlsNrOIbpGKNWlFfd2cbDrLFYJhqudkTjtJ8XT+De1/0pV
T/TStQa+pToI32sWHYlGzi09+Yrm/kU0+ixXhl5xaMVZRQBdkaEYOWaj8XeNyX5V
9Sx1B4z40hWE5dFxZJTjx9+sTqG9AHUbWfpLYEvn+LxskFt9amYWgwqRgVlt4tt4
6MkT7aVqbyVCZaSKOYY6AQ392U1a/nWldXF5ZFe88fm/f41d9EkSHBzg2aGFQ7qm
aGaKbubqrpBAqgIUcAS6XE9EdYcz1yfe2lq9Ni4km9LOSuFrIgQWfysLPJ6Cj9d4
EXI+4IsBN6rAL7Nss5IgK7zpujxoagwmQ9paT6SU0omokpuN3vFwxX98i9wtdOdp
T1Wc915rNW9mGghYpU/cSkBcuErdq6M9mmsSTYue1XePlqc1BoWni3vGJ1MZ8T4s
XFFbeguv9XakpJudMrslQqkaK9oOzoQiszJ9uGBU9ipzwvATkvFCR5GirWO4AAep
HfgdeWgdaL47G6vxda+FC+IPI3uPqW3vkJgmi6ecXTZ0beU2ZJTdr5ARdwGdIfHW
RtqW1z46R0fiDeitd0s0qmR+fu3/qwt1if4dA8h+E21NvmelsUIEloAYd4ViQtbH
yOqDpbsksStBVKztTicZmHy5rAV7twCGhiteGXyoOhIWAcgDW8+fnxJurU8snDb+
W0EMaxL/sXOIWS7de6IGtLKVOvu/x5IYAMmBzW/CxKdhlmV6iAl4jd9j6ZsYHpN6
gxuWDtQ+dVMKSdyTXUN9lPNoh1fmu1YyOHPrPvUpcVwHXSv1N1lZ6QQ/KJSoqQw+
XNL7Dz5UUSol7TeU1DTxdiW04Hj98vUzSfGuNEkSaQUkO08IUizkBDQ+ALkUpUAc
gwulaWMDFcZTYzY0DI4KxgiuIlIqE1nK3JzY6ErKWtXi/FaBQmYglv9fy6yKS71Z
yZfQnPU8lfZxEBE/37MTzAgCbUsrNlYluBUU8DnBINWiYEBK8ch0w120W88SHbbN
wk1D6+CgntDoJpdk0IxTeArZQ7yZeUFOaT49SehzF5bObtLaF10va1g1fy59ua2t
YxoLLskO+vB1Uk2Lpny6f1WzlSir0ZQI5Fx6x+ldfn0Z78VdcbQ/E7iwYht/RnKD
LHagDESO4HN5UZ6QFCNu0OtB6FITjQlv+fhftg48fBVVOz0WsZQirgED+dzSBPYD
JFmiEmW85I0ePpuYsnq/4IuVCuA2LXcmBGdNYrjXckCTJhL08WcfyxI1k17bxwJP
iwCYlLi4srUIwnjGQdsjfKuWOx1JriERkxkQth2+zJvBSVjT5eiOy7I24rMPX/tX
glBc9hpwc+H7MlgnAEEM3wwuxrF2GBqskIiEN2YhNN2Sp52PHnIlXXpOZuQ8IeL7
dUK2H+fgAZl+QXZ1Gdc1JdS4ver56klDNtmG7vf5xNcQImEWpHzGOwfxflr3UsqG
2A3yiqVZeu7Va6izQ0ZtAKhmKqQFjiFH1UMzr8uwL+eHgUeTwhTwk0pI4p3ZFHAi
JNeoDQXRVeD0TSQCkVfMBfT1qi7n5NUPUt5nA4ItZz+629K+14omn7J9YqfuEgHg
wyksA0QvMe+lsXOfe6Q+FL0eW3huC+Z7MZJy4sRbuXP6MBWUpbbfbgbDfW4Il0XH
5P+ruaGJZacOPwevovvVnGNTdSfKJ72B+sCX6CgoaFopI+FxtqyUw5j3XBNgFcdX
ux9A24U8gYPuLpNAOO/J9QzZzGrdooYd2gKQjdd9u5zk9FufFNLVnuumSkXrAemp
UFvh2aU1w+xPhabG1oTENKdAkDLFTk78GRBqPwnjPql9r/6EvEF4qIPxRjLpKptn
nE7IcvkB1v47ey96kHU5AAUQB0HUIJaTi/F8JV9Ss++K8vxf7KYJPtmvs2lebCXF
X8hXF9BDFUx8NXKjQZ1jFIZG17RP4aJjaZ7CqrOX0ZGgLKz45rYuz59oaga3td9l
aLa6YqMhmNaDt5ii6BaSLwwVZM1pqnZ+hspHC5o68bDJn5CrpvFcPhJayGEygcoI
U2cSa4PmElTG0o8Osmuf2Q8XC2q72DToRZuciYYvJuDpXUrPw8YNbgvvRvyk9DkM
+8jX5kJWbqNFhvVizpmgUG7IEtthReXWyBM+UW1ij/Lv+1YHOjQuyJ4Ct4MRzISW
n96fM4JNqz8OVxe/2g2+t9pPaRbzwVH7XqD4jPmMDFpeHiQJbvYLuWEuA3gGxPL7
9rYDAVlVdZgSoA1U/wWNMkzCTN/GSNoAgpaf/oBQUTF4CYYpMaWrdma6VQE4cqfv
xCGMFKCB4g5b+l0mV2e+XT75ENUKJMZRnbYlRChz16EAkm4UFBjc8qOp7DXHMxmv
aqpKrp+63BvpC/uTAInRTwESCunHFEggsE8oS9pl23nqCdJKJresgxIGsiKLrlkF
7MRfjP/DU1olnHkijEcx9NmlDN4DaO9+5iU8GpSFa0dEZHsQ2YBODuJLDjub9XGK
UkhXcMnylNdFgrO9O7ipcECMk8SdRbTRh6jYhYpXoLFgH5BEYngMtApqAnC4XsLN
kYyN/z9skOxqmep2T0pj6uCxDnO7Fj7dZ9NOYJQV3niBoVoyEGiiblDW0VWnZE6r
3HP22jF6KmlbL9oNBh9fXjSVfc5dLmW9kLE/vFCIuJwq6i2feVWGWegwSXOtOnIK
3dc9mNA2nc+DT8XdodY/4DgX7bNNQEge4qTwsLFaRr5ol9MQJhiJG+EMgeNZhZfL
jUSbynFYYsk7+CytQKRwUdfwFXuQufdDF3xvKpxRNcmjJ/lzAceiqCVZ+yeRJWrH
W82s/YFn0VrV7K/omka8BhCrE0EQdGBAIzk/2xa0Ao2iWWw2Noar2Hbg2qv2jO/0
B01L4uiuGgfp5Opv24VIFyXn64fYjJKmIoGV8w1S7Po7zSK0sjN+Wm7uPCgaa+x9
OCjtDFSjexREVcrAENIFcqLGs/FQVYsRsntVhvXgOTIB9RF8hu0+OtfdJMZ9KyhE
VWzwf2EWmrOB0GidA1vujEmHBSsShzb5NMTyFV6lGPATETizO2kwDsXuTqyhMWrd
x4l/ywmWe98NcBfR9i9PT3Ws82RMRzS17+lMJdjQGl6PdK7oonikdijdo78NWjZX
0fykAK+zgxvlIDhivaH+mZrqDt/Uhxv3IDmRjc05lP1WXxsRVhGxsFZADbbkIyTR
IhGedkHvWee64s9DqS3TTJknaeiboBtQF8dQZh/j/0TFtqETKqUb67118ovOw55c
Op2+vZvbKKaIdDgUlWof4j2ILyYhVsHYS0fcVd/5nGbaDvpXoUDmUdCmXChJ+vWQ
dzQSYXzIKJYPJdf2WI1UaEAtaV0zCWdeUMgFbpwt2nWZ5wBS4nmghGfUkgSHOSyn
WEjM5Rv5uLrZ8An4IGigSu2zTvbhpkQm2+Y8elwHV5XN/uNoxp51ZdJjp7eA4C9S
SIA1DmbfDt4DRiNTES4Rng1QallAf7xeGdnUxPNZ6eSF/O9AtZR+lFf2+Nc566Kx
IoJeoM86pHNXVcdchOcyQ607D8bIaVSP/DD07KileHZirVI3MnO3x49y/pvRX0Sf
+3PMvdEwu4FARCxTaHsVars37Lnzww7jEIKM51dZe2W+Tt0Rq5ZZANZDYYa64MUl
FxBpkbqz9aN9JdSbmjYVFUyva27H6RY08koMOoYkGbiYq8DZnDA1wXp9jODBGD12
i5xzwWR6HDRrBrQSJUw4OeM4hWqwycoN6o8/OE8Be5xeou0uhB0du8ew+0WlL+1F
8bcAxyL36dg6yrGM6cPNYLYSk6Kms0DcjF5qUgdAX3xCPFx+bjo4wsX/QWyqidgb
typJhDzLCe90j4iOi6xTJoWdbE3cAsFQklAeC+5AxcLTvbFHdC/EL1kfhgbvpE4n
iNfsdnZMKgNW/xPaNPKo0SOAp5kTiAlfdmMLCTfOROH3uLIRDA7FT3jL9CBWYogx
SJXno5YFmCGvj4MrKdn0NvSram8NQxEkQ/A5selWnPMdVqTB+6HrnjU+uVeoU35L
XZeHGixGRLB2diOVmuc+sXRfvNW0FyIr74xK6G8/oE1wSN31fHMXRzqbXGYsy+VY
uvQyydYnRYCeUP5K/3FHaEFWs4gU8kxP3I0sPgg4j0p7q4N804haIVV9mng2COCd
ONeGo0dGzfzyIr+fnQX+B263LWcRjuAB+OoyF6VMAu8uKPif9jz7ZxAe+7Oc90Fd
xKJ5u20CcibkD8Hw9XRBVTwr8Gexh4r24N7IV82cA/J/++ifw3NI6ydxXXN8zpgo
T5d4ncF3PcvgK/6nP1ygtEDH97ubsOxgOHjBQOPPDfuQo5go3yScfJO4nVBCm8gy
Hp/zYM2DisJgamPalVJF0s3WXbI+B6qoElm1m42oXrvhfzun8EIBIdgKSYCAt4EC
yfZ9V3mDYhDqu0pVszpzm4NHrNSbJaBlcTLRNK6aXHlsuzsjf7FBs59Y2RdIjgxb
nsq3bcKXhu+BMy7F6hqWHIk0+rS8a6x/cjCtrJyNZJeg++OXWD9p32lKVmo1+Agr
Sp3ykbYk3B/zoiWQsezd0H/0bTlMuoTLMlVFZDrsGmjspvLdW1BoNIfwkTZeiE7a
2DgV1t2jcv1qkO+v5yj6R59jpcBew0DMminorslFz8jVv/psxbG6a/Yf/BTrxB2j
rbcmr0zhNUuhb8zf6bBBRLygOWYUhs94TulyLfsVQB1B0/rLLqegjQQ4qN4BlkyT
S1/k3Xc4904prCh+XaeeRLU2zzohg7d6cELMQcX4/xWD7HqoQSuOYKCMAKdbOAcj
4rFbAKqx+h9dTazqbe0PU0CWM9sqAUCw7ihwZlZATK/Vw3OyXhxpv/Pcgy7Jb7/U
JZXwtj+KxNkS5Pr1lOPsOp595646tseKZuovNNK5fHbGq9JKW8ld04J6XGwnKpSH
Bq9GkfceTDX8xvj3hnQ67OZr54vdxVO6Q1pITsgTWLBD1oXJ9XEY/C1VeqjVRs0L
cKQU5bR/6bHxuCUWBsXUGW6YD+s3BfYZQEuMAOJ9CBd6sqPzrNErSSrUD+b+CX22
cCC160IjyevbRBvtsqkwWR4kHkBEUUyb/BlUf9o5q20Pw1+p+vkRv0A9YMb8eBEh
ISyd5xDSl/NVsvJ3o17jjTEyJHc1Y8VQGdD1oKBaMquivvtFmSbwqIC8bWMSVq9d
6fZmdItGyFU32w8Pda4g9uK+0INS33gwLsnm2pnzLxAv0Q3TBAFD+V2svQvc+wAx
Lc++hJ+NNspTJ1FZli5jK96nqcJ85pAm75mmc+9NX+kK86Lu9r9vtYUIah0yjlWP
jHO6EKhn3dHqDJ57dHQlXXJgLAa3Kef9NFHNmh7C8wW00uuL4ETUpoJKOuhhurbK
dOyqT1qL+j839X66XEEFTc+KurEbJq7qDTcFdQ6EIJNKEenyI9YxHfN2f2SmzHzT
Up3EI9LV5QboRTwD7V3WtQOPOh5HwA+1PtvE35Rm0whJqflsm2kg8h6RH878sOZ5
QCnDw9x+n2qAWD1HXHx8s+Zvs8BrCFC4mVj5cG5MIswdmoj/yPw2mzJchH2qP7hE
xuDMuaD21MshNo8My5wMLPNp6WTQRacpM9s4mQ2dy4eWQU9/RFSGnXHSQ+KIAZpG
yq/umJoQYMXvGOH31+gcmyk5LBeR6v55Tdh+p3vbHu4cuELUc0nIs7IJQpFOQgbN
nfl4TrPIG+C2zuItubb2mnuJdg89XJWxPIbCpWgyFphYj8ud3+vzJweYy/GxNLrx
QoYEtFJJeQIOw+rXWgTVPEA0kKuMPCp8+rFwy8ElnMRFJmsEBxSmEwWA2FX5L24+
8+SlnekgkAcI5m8E0HX+Alc8W1XaEo4e6wWOYfYpe/QSB1/3IXqsVBGKWJSYWwt8
0HrYiFugzB43cVk3WpMbHZUVmE3CIEFby7JKDff9q60Sr81DK0TYlreadgeBzVcn
LRKKM9DDdQmDDxPbA6zimXsScbTTKf1VKPtQxNqrBrl9kvItjwlVBaf0H468pEgI
N7b0gmegF+CA5QtakH/VaoYzoE5o4/09uz2AxFP+m6eAKO9UGMCbNrj/TtYSDFcB
/N7L2e2bKXHMbCDXiXglzfbTOZJOT7F2VVjl1/dfpfvjvqf20KTypI01dvoI3yqv
bkgZO68cj5euZ5XFIj9pjOjwK7s3wnpF4duojkMKuMZxH+ulmMWgHyagSXR/HZX3
BtX47re+enpWi5grpY9t5C78nxS5UnPI8GmIrZ8qBbS8Yw44nt7DjbGL+xIW2YFB
CcCzKc06vwNlYI7BNxigRsWCPlvDSZ9oeSDMkh/PjbaJ3XodA/rjpKw+ICJsjV1Y
Me2pEptNSVg2UNctPaC6Rrlx85QhdFEgF1iqCksoLdvyNe8vBJyz3yGIoI4crDOM
JCxtT3ww7nQFjC3YlwOiYyrtaDnit+TNkCSxm84ydfz/xrT9XsuQqM32kKVa2bLL
kw9DoNWXQDP2jV6WEUSrqLAZkhaIsfzjB/GrtMla7qguZz0mQT1qKvZ7g6r8yLJA
Stch4KVCGKuEwlWgJhPS+vjV6I62kvS6CGzWjuU03fhZcE77bZGDG+D7+NF0oyca
eMWstRvy4Wond5MOPJ1+sATHgD5LX1VcVw6Z76xocoHxa6iGWOiLGQdq4bOznv/g
B9Oen1U4RXae/v4SvWW50C2qCqJlNyE3t0rZ5eQdg/T5L53AH5o1VQb61LRv/86a
zkNCAhKAXhwd7M06izqU5RIJeeCYSElQ0ubSCnlFvctEy5hRf+tQORgKK4bzQqJ1
2hr4KzTSkOrRwbvVjUcPfUwpA6YOB9Tr+OV4K/nlKGHTwQjYz4aIMqJ54XiDqlZM
E99JrYYeWdeKB14S7cOxX9NwhiEfZDcXU8qlp/Ad4q+/gPL668DNQAuCQkUvnCe3
dRQc8QlWKajjeho7KKppef+sPjJGykEoIu/oe74R7LaMzHSxhgvuQl1MjowaAIct
oKuLTUG4C4LYZw1u7Y9crt+ZCg8sUID/CICVVliBkUxl/1ScJA2fyjjxZZN7PyVy
QF5sMIMRdOcsnIsRh6sJTa69Uz8V8z3drv4lCSORb/WE8Ll0sI+E3wMaomw9IPAi
f+hhn7EUC5m9Q8rz3s8EBTOQOxRMziqZPpWSvUwwXpJHuyariZ2qy+UzTWurgzyF
lv//BIOljrkISqf0GAzBp+3L1urQ/KRzXoIQ04S9QP2V61+S5hBZOIbXLBLjaUra
lm6o8YpOEVEfrTi6RlkemIOy3pyMWbsiPvB+wn9gpc+UivrdI9dcjnGluaxaYIsF
ndWHgaA7/WXqfDStjiOjUSGYo/mH0hgyPsqtERx7Oe4jUFyomLY7LidwPyfab0Ew
sIaNp5A64HsQUAWQCFf4pxzhxYx1kP8ieJ6YIbJm4NC8MCNk8BwpuZGAHjxWzX5J
8riKjdJvnN9XH7t4h//QCuP1WwDba4vHYQ3RowkI0Dqa1RSMHnlvDfly+z42deuk
NTvkVrRGxKpvnKo54BraLUQje7gpT+PpEKlOwekeKiFPaaG1lA+C0zpCBx4jwznP
rX/fe+HnjRqRSWTPOMUPSYn/zzlI9oX6ahc0BS5xTVYHh3WxEncHQGxMa7koPjXH
bTsFenRl3sJHWzMEa8y8kt33GlcoGq8llSKN1Ad008b0XmjPrIt4bzAymvVBHWMZ
qpDoz9LwCnB9gWCq0CbEI3N2jk4HukOwPG2qt79n6TJPjViqkeyvEWclLlodMMZt
O/5RYf0ZS9s5rhPZin6g4N4h6RukA3S6LpDj3ift12KEhfhEU0ItvR2VvnwIPAQO
dlQIq8veL+APiy16CYdiboVM9Xr9q0Gz/vJDFRjL6m/OcfzdDpQlOi1fkNcpKO8r
dtnET6TOhtgn3C4WJDTipKZky0u3JWuHbkCZebJXUp1DSc+mEnCGOgPh5APJqyaH
adR5yFJGq2EQME0HUaO/sB6twBQn64snX0VO6To54YUtcft05/RyEEhyCrOLZ/m1
N70PLAGdDR7+S0XhtVVsPr4Um4UkYlRtcTjFvPbesGWk/9+2pJYF5s1ELy3bH0yt
13axJbJZgPZuyzqCC4EDkENuw9f2vTWZmAuhHZNtBo67TvnW+lJyfwYiDO9d26CJ
ClbTb+rFFpCKSPhPbxg1wPyUUV5lQwUfZ8zAUUF8LsMWAX+AoZjXG9K+iz2pXLte
YveoY6OGh1ai1d0Z+Ws1DZXz5jkiO1T9lBpEjLHf7Htqwle3vujJP1InWqxTnFHS
AJHcXyBAcvriY59/fqf0mcPtIX7+WGtnImbGVokn0aH7EYQ/5m/mhiNrA4o8y1RG
PnHPAk1tHhH3wa/FmLfujT7nfxylcsLY2+QymKKg6Skd36NVEJtE+pRZnO0UxT3b
BpYzUXLNZjlhPT+H7SRYA0XHlA5KdgZMLXv/phLVAWFd+XaFI96D6ECt1bLZBzzU
YvYW2q/EATeDmwHvcIOY6mMjAKS/WsDvTxDAUdJYYvhXRnqsulUxiYri3adUctBQ
Z1mTAT6fjjV9Tr//HT4xEjG/CeYXknf+erD+61Rb0TY1rgrtzzjAsS9HzZqKphLP
9dYX5r9+hq0nhQqiKw/Cx1nokaDoozuc/VlcIkRysANQ4tSzS2iJecNLETTzGhmG
achrxv8JYBwix1mu+HJXraBVEipJ1PnBj7KN9fRlpU7VEpXMmTBdVX4d+YY+LOQV
xYgwHuevRj2i3/V783063ubnVwBW9G7eVsfjTjRIM+o/KAjHaK+D8WJVeGX+luc7
08wYA3HoAy1Bve3ShDLVBSMPbIvYaAVXxcvog9VXNVCzFV4ukFMHHTgagC0gSd0f
gHgTyTGhUtS3TP1BzUa/ddN1RjA+fzYhgxG2ijYh87ej+l960Z0/qvYcfiIkzdkg
IphuDWIP9Bu6fGbdYI9rwV2hAjN7WaTHv1vOb2lHBL1W/QHL9g/7+/DoLDMuwrHU
mFpggxBoXvWnDM7ObAD4OE2fBukLSDQe/xXKWk+G4XOhiC2qVNcai/o4A3SwNM9d
n6B0jQZ8fKd8XMnIJ9AvIy3QKIyyXiFX4V9boTxGFYDAaV0FGgVdZXZudcLrx2L3
SDtY448bRTiYqzoBlqz56rBC9DXDA6KbAj+bmrGkzuSp9bXD2zBMsUBB0+UTflJw
7iWxOwbGFAXonw4KLPXvFvF19zfmPeVr9e4nYpbXJSTPTg+uWUg+gFceKZyvRYoh
MJr6cFVdVj4EpynmPflekgjv1phKLAqaSVEoF/hpZZV33EO1/bnfdosRE19AI63f
WeC7yHRShzoXOAPAtv1rIiIEtQosUk+DlasgroKZrdVeKEQtjQsOl6EfKfDFZppb
JymBuGn5JlvEGZU9QipRf2LnZtRFYx+IaQeqhOYKW7K9AoYRBwgafYdSdagbELIe
0stPKUqV3409u+Rpo3nUNo1HW1mYt1HbildD4mKd7469UE8vTOKhlJD8bU/i6XWm
Ef+udSbkcSuwxW62rDBlUIQu3swMbT4Bcv5rLMkBBuEL30BS01EJ6JpBkYko/z3y
3kJafVrrzi27p5wryp4JgVGZdZtT+dsHbPHGyK3UuqYj78SWA2mnvPf1I1NQW0Fk
6qqwZLXoKZ0fNFitt5nFJ8GF44T20CNgrPvD4QAQ6pbo6Ok1vytCNKx1HkYqzS1v
Xzc0SE/p0/uwWFspY6YioeHGqWKU8pQcPwDgB5Y2AD9vKAcBvVw+hahd/B4GwW+X
GJEtCRhI2U0caC69EC7StTGcNye/KvnZmrk3I8+kod/hVGsWr0I/kptbC/qDzB66
SNYAVFCamjTPF5ypjtfwvbUDg356e4ljguPL0OUzD0KXFO+nELxbNqSuuI5SYSa+
7EeXVRfWp4JK3cKj33bQODhkSr5F9RRS0c+sfou2EsGhKweRTVFpeEV/UuhKAxKA
xWaU4z81ZK/gHawlwvW3dFDDVVB258osPiM3RNxHAOUQ+ykaGvuXFq9LniC1OfHV
p0K3Ck4wbBx/c4GVvlEDuFpcF4SDPIK6DLMBUIta1rTZuftM1y4vo8ofUnzZ1x/e
86ryVK9fTH43PSL5sWok5uHaBF3emoWGa2Iv5MKNc3OoQ6ZzvX+Wwr1fCVMtTt1e
LmfhS0V31inGFh6VUFB1CrtCHTgXOyJ7A/gNT5rNk9ofJvE2iYryH15x/BmIC8az
8kQQ/OGWRvue2CaKXSKScxwb7Ccl2xLlYQjV6AtF/iMDDaTfWQfNKWeiRSGacskc
Upn8uWgKw3VQYPMJz/Jiy/RY5pDfr5PdGzsUNbLgGWsfHc1rtqbLDKlSbsmEEyJp
qEwZf88zZmLONw1K9cV0G7KFCMfCCt3pkLfHN+8EM6uZ/yLhE80b1/FOsXugNjYX
4rDFJqMIi47HtzL4+Kv46INSvDSRc4qF+LvDLspbvkf8zL4l7DFjq0ZkGl7wqswX
69+JiID2W9Ie1fu+suygFF5tWm10UkXfXf9BAkWUckSvMYnSwgo8HWPYNlE8aM5J
oNhuGkRHq0TpXriD64sbptlVH5eJOZp8sdue9ZGHC0JWIqNCte4bKUUiY+BSMWJp
ZbQri5t3g4EI427Uu4dzaZjQe9SEqoMLpvw7hORr6kF5fj7CiwK58RiuvYh7ktT2
pQjLbKG/Vu21qKXj4rK2dM6x0Y9u0wzW3b2IrhKhEHc0Dh5LdKjfsSbIiz2deERe
ApXzFlAsZbnLH12oEruq45mRc4/whOyPayTreNksqL1hNqr6XdgxQGg9CKvL46qS
6Vk0iguT9O8zzgNO8VgxrvESi3f2osmWDlKu1+iXy2eKgjKtcrMc5QiiK0tXAMxE
MbXorRbMzmMYIX+vTilPQu+QME5qgluKdpF7heO+mqk8yEzQb0IXy1Vqemi6F3mS
qEJjLQYfikzn85copU9JqKTeijwB7wNVNEHwiVvt2bcSaDCNOjVhWK+Xm12Vrg8e
K06DfT2OI1Rgl1KfCgYjPNxb/x3zQEFe5BV873L7ZPjOUPhf8fo0stPeoeOQall5
OUADeKIEgYc1a5uOeXyWnYjFzeQNtJjIa61o6QbCCFIHtNGHrvK3qps7OgwrcwPS
oZvH6Ka9ijkCORQiDSHZqST31t2kb9lfwXUhUSJLT+lAOIai8GFzeifrM0GvYAZo
3kMvLdCsRWW3QB/TZB24jhmBjo9o+MLgkdXBJYY0HbSC+tEuN9prwCAVIIatk1ay
SkLNDBQQuaChPqKmsadXZeJCEpf9awXk4ireab5BpgHOZCXHfGfJWx6QcfZkQS0b
B0ai8RCQ5rbRB1vmyeuD2ENuUGzeN73VN9AGjtZSpf+JTX9JbVXAAo3s/LakZrV3
Cl5jsnueu6ErIKiIoQleR+QYBt865inTNeOZodxuZoIkBLKiz0SFjIv26NMG8xlJ
689/tvsyN4ntBvMbdXuIXgeIIByk0hwvW2WmXfH2luCRIDZ7D2yZGKlFwUSyWBxh
45I6QW2lFqd8JcFNvt5aF6EV+OthEPqOoSZ/iZHHKOXXvuHZiWtob/C7dy9YR2jd
2hvW7x++CiwT7eN1T6/CA15To5PnYPdfqP+4XwUfEcIFVO9CCLowI1lL7yxg3bGn
4UUPz1NRH3e+MKE0HQ5C1cizitp9E0eAecVWvql7myahocgXVY9SfAU6AdEQg2s9
/kLnQ3ArhcJK9Dgn6MSsQxzemKZNIbXLuW3QQjR59r/IUTPxKKVDi8E8KXlrvf7g
UwUGEq4vaCbZfsV/5cW6xWVaXVZFgLDbohKRxsZBsWWlaT5GouGrJCmngRN37DTN
CoV6p8UTXfrVbD05oV83nxM0LzisylnNhuLCCFbeggZRYzOZ2omICFci1dTcRs/z
7hKyo77XBo3WniLd60NtIu2cb6JfBzjDRtbpLdmJbvvsV/yRNZCgTTGbfd5SOTx5
tugMOn5AP0uKn7lD1czh1t5vOAflt5hTAddFFAdh68lB2K/xLmTeLkDZLWeFHGMt
2yHYlNrmrU+vCACDj9363qCD0u2ljUf3ZFkrQs5leL7dcdphHsp1VUwfvfpAFIbv
Yt/3ZGfnXaA2KDfB7FBehyczpiIr9tXKZB6nI9xRdd/v9X77v123hD3kaOnwQTXo
AeYYwy5Qn+PWNlQVovXLeix4X2+8KbV5JWxBWTNMnIzBWAUAX5CbITwIi41wNmf6
DhdqpI0aMef0EnH3ScFq02LWwF5lVEDcfHHSJY97f9t3ojeCdSfPHH906kguvpUu
2CoGb83LkI/dyUd/ytHmDKHpKUoXMKyvwx7Yq9SbALh0unjTuxr69+bmQp3Mxh99
OTT+FeWKN+jw+eeOaQi26stoGsDtEFnqKTZBNAKt58qgdGH8E0yoVzKGKH8c6BA3
1SUlzM1U1tWbESEaF16v4A4OygnGynv5SGd9zK1ffAl7F4QUInzON5iwd59eyDHF
sxAoWYWn5tGZdJW5C2QPqECcXxJ6y/ewYpEoEIW0BooQSExTzAYvASP34l6s09+4
yG5+n3Kd6sX8Co2V3g01P4CbgFkpNDyT/OnI1507KN7HoP9RNUK0jyAch2VSCJEQ
lXbf/6xpwqG4nfEmlZp4HQk/LGACnnc0AwrWaZ+Bq0rdZgDwdfvesiCj78Iil6Ti
QVf9ndSby/r7KIXXzkRF/Aft3xGloQXYVx7fSyxzqYMcvf75YWYCBBOZeBUBuzp5
BLveDAgawGDt2zpiWVPQQMtdYUM4sNOZgmhBX1hx9HSQbnaS+7pCl40xg/vph0zp
hmyBvlZ5OvJSpB2AUl3E07YiO2AlVPtOSNNEOqVyUcpSUykSHm2I83U9YWRlN8/6
7k/bejjTs5/tYrhd178AaWgYEYxnXPgjP3Dw60SxQUa0UwDA0WpcFeLdojLbWXez
QHXgKeD60hKwV8kqMjv0LbStEuDHl7w36uzgYOknPQLxS36Ul55kQ9w66vAmSrRW
wASMnWgIR4H/pFQRLjry4i+PonzJil+VjFbGHBFxB/MN8Gm00winrwzzzGL2VK8Y
A3XNbuZv0W4NA6fVxc0uzZ8K2M5bbzyZOqU/62wi4nUStP5xIQzllLVpJiVEnHWQ
+O2i1KOkgRbzy1G2rIwRJ4bA/g3hAZUzlv8zIw+B0CFq6I8X1Gzm8sO+T8c8uVAl
SfoavBKVteyaZp6JTREdtt+1gBC2xOUvmXSS/l0L1dbhviuW6LlR6jG6k7VHzZFj
z2wDEQoAplJa4l3j4EV4xCXq0Wea9jWZixsqx0Hb32l6atQSH7FXssZpjpnYjRIz
Nw2s87r4lDGwS/NcYytEzLlocWWpsGO9pV0iJlk+/r/LBrNGL9g+h89Zfeo5B740
wqgsSVsL/Swo+MUfOQOUDNPJJMzXz2Fz3YPzDr0g7M3yq/IKLGyG3VRlvutsq0Va
9XR3KEzPkxTX3YbAIr2IBNJih3GxGOukfbBBiEGiaIn6k/5+BYfBEDkL7goVnJMP
h5Muay0ZcopE/itRU596zvJmzF3tXDUbBysiI5mlLTbJ11KZndKTM3UQ/qV6ktKz
lgVxMpUZafS7H3YDk9tHst4oei8u6izM0fNvshBBPTPoJUeXVUokW94lFZkK47BN
mpKPJDCWyg0h/FHaopaH4YpeNMB4oZb0PtSHcD+63JnhJjSBIvcnyf3gUIvPcfcy
hL8BwwZxA90xpAmkRCY8wluQxnh0WTywfbSvsVgg01n9J4jadwkSkRrANUuvDa0a
cDNeerukYqyjRNCJI86JceBK6mno2SfLUvGZYydaTe6XeR+IaYnla955jtIoyJa/
sO/eKfYmr0Cy3D6j086JnRXMCIO9yVxZKqVcFkQOiDzBwb2rqdK5dNjUwHJPwoo5
BZQZ05o/dkcTAIu4ZnyvIEM+b6AtXnZT04dU7IdA9wyZvIqBQ1oTeNRKimbcM0+f
sLfxw9rZLQLfpAcC/AYMYiW/8Axfon3e/ju5kTxOKMlU5VKjrxyW8nBoB7B9hiF9
sxK6ZxcajH7OCuQXYPh49TcOPnhKxL7HOc4r3fPqEKWvwppAZJV6lMP2+RO3aLjC
n1i4mTfIYPIqHr0DsuKjptbiNMDmABjx2VYqd6CvU2h2iuDaNWdGRitUdFusVgtj
1zAqdxUIIb+ZhH1SzIE/XeHJ+ikaNf5wVG+dGdDb6ZQytU2tJlULv+Vp30dYRNVa
NE/W4YmQJ3C/aSCGhy3vSqVjoT+G/M+jJhMhk5Y8LvCW/BH3xVcKQ3/M7ivMphAN
mUueRYVM6jDHVcAQYU6+pS6Z5347I3yai/2b4cOQTuIToyAi7aQm6XNf2KX2l185
7yn4SN/Jtp15/Peg1anqwMTD9RxFlcG9JPjudaJNLkb7tZCFmmQMT0Dr0CWbtt48
a8KhlOkb32PLBh7pUuO695itVvJ7AKnp6ztHhIlE/Sw0vML7UEaORd4Qf8DRKj/U
X61tnygVO6q0U0erMkIAWqqiGBfA3YuyDN0cUACoRT6LujMbh3DcXdQ8Pkh7/P3h
VVyBznAuWxtBx3H2PtjJodwhqYRACCGGavE3GPBG1flGuQhRFKXXOfKbt+B2Ozm2
5X1xz3bsA0gWCORuSbpFPgbUomYVdJw8nCLddHV51EOUiuUoQxhn7Ji5TrM/ka+Q
4popYhpTZrO6dJLIVNqvximSrETDtOF5t27WidgxW7rrkbIXYhOpnmYh9V1p55n1
CI1sxBxpxTOZDuhXntrsOwTf/tjETezP64JmieG+FFvsApus1b2alrcY5rk7++p3
mK1df7GF0sIswWXTylgvixNycc6nkXgq2M0hxdx/I/ItOnZt9Gng/evEwluyeJdc
AMBajuHf3HBfKkfY4iwZ2272vqGZ3EMQZFPgGAjMPHdM0Kqvx4KetQhPiz2sJsWc
gZbnUAgYNiTcdWfedwggjl6RxGHW3sX9OxpoXYARXpeklYEF+F5KEBttM6n3WLBb
oIcMMsl2q76HgWT/0WHNbbmryiXb5BGFWyhJ0GINRl3Wcn1TSYbnE1gDZc00QQ6/
tBRxFPB6uCfnRATr+VjiZwPiQOOnIaI01/F+2vFexQ5TONRYbcEhLRwKRaGQP+I7
bz47yF/KsctXcWHrnoLRup9iuusiawpC4sc2CUjTXsHDUmmXaLlbepgZPh+RMnEO
HBPETmJIDcMnKsS37+naWzOeu7ddOkRNWF3TEaGQLqYivzzppWQ0s21kkBiKXz8B
m3eKf4E0xkJtk896pRKZ1fZVoZ/qoCrvOyNENwlAeDQuglhJXv2qflfgMx+vuZta
xgRE/3zM3QOPiIsUTlmZ4LY7lTte8/7ZlGUOTXFr+3sCCBf+3NDaZ4Zxy7oW/7Ba
WAOF4oIwEe1y4gXc3kB3TEY3a6bOoEIPVsEY7U1rcTHbh0S/h0XA/DXA9jcDPKov
4SU03k9Yhw6zi8QCVszh6ucC3o+z/Sp8vxir2EQ6cx86a4jlfG2EKod4u+PTXzCl
VsTDTbAdZpyD1KcGxLdcbOTY+JwpZFk4mTaJBhv8AVTcWlvWYEveZ2gmuTKYONmA
RjqEr1ZA1DZWL8AeKWXXDxBDym79ZII0fqNUZwvjyuZu0Kn/mA68QkLB6or+tZE5
rde65Bf1ZxK1fOGxZhriwWURex7XbkFp/49DxuRWf7cw3wh79F8ZgxrMROlk22E9
AddfZk2V2GhEkY3wvBU1siZYEKRF3sCow0mBklxZlG5kcvFTbvSq+Z2gIHrw4+iT
z4WhUwDq6rYMwZt3imxpIneGzPOdnTRGfd/5tEjATuHeQ2b2a7WNZ9i/wjmxG2rX
lqVqGn7tDZJiTHIPmaq8bG5FMNhK29ZIdt2gxnYLZMOyHK7g2uqK5ujoHG1PI3Sb
ThhSTl1xhKpdmXQjfUe4oEwKQ3WsYx7tIdByGUqLa3Vi8pEz/jFzq9TqiIQWv+b7
1h19LBsAYYN7FKf8QSd+CIW7eAujhCNWR2wz2OiCrDTiFapofKOX92R/6PqO0W9i
yd3ThHffIsFEiAPH+B8HeEXFmVHxATdp/IYIDABVVJSPjx10zig0GDK5vCLFBtkx
zG4rsffU6qbNWr/JegmCXi7PhSXahraQBFQRVoMwKDTmbC3XtnQJBqXeQkzlRdlw
vZ2xY624/DPyxPRrIJrV7ShY5cTTriYxCZVmJ21U0i8RdLwYnjPm7tXU+8G+C+lE
tm4Tt7L5h1CndKocG4GQiWv0fuGT3Q4kzsDpRVtpnS9924LaPdeZavaExJOcxi+t
zitYeN6wMkHvCuhsB4DWUUiTVbxY04Mxxrz+1ajvUpZLQrG0YuVV0jzgSzx2dbfa
iEpxzI/2oLk/k4uh1B3m4GqsO6AMb2XDn8fiRKwV+c8b97WNRLGb3BNF9/sRgUBo
lcAyigIWyQduJ9DOKQLntd2nZl35fwC/W4otuosYFIN4MDIH0XSzv5iJGFr2DfaF
t/U6Uu7W2S34EZVTrV91Qb5BMs3d1p8393VhMTzC8ISWI9pHLBLQ+1OJ8Id/FW4G
PuYn0tTs74EYv5MDNBSva9ZuidPT/cd790eJlWHpN/B7FPYPeHn5gWbU/O7ZiIXf
Liwa/sBsR041yHVrXEFWgedg9FXmSG1T6PhIJxfGEMdHVH/h4Fltj2SSOD+WQJ/5
P5wgjxW2D8bq+hpnbrPBdRBUOm2TFfZOV56r2T6C88TS5vRhzjHBpGcutJcOGcXz
GPMZ2TmYamHd46+pcF9reIDyHNrCjNCUgR8wRcdlmtMJUH1I1nfS//wNLsEeslYp
ajjV4iD+t7EoCFL7D1c3C5BT4caazkxt+meoqTYDuHREXPmYT8YwuCtWiA2qtyT8
VOWh7flFgVtNM1ikqjfpmEZ4eJC+lgZ2c3PZ2VmSaVaoDlfJ/5Bn2Vkmd2pc1XO7
XYeZy4/4BErsZ8eIyA/Ib4UapPuBEG6N5oZXH1K3CHX/qPSBiCueNxCLC6eFLVOW
pIPN1+Uxryc50jR2d0Nrb/t36LekSQMjcAaJzSoJmxSWaTxZ8eW6+BU1V9lnnBR1
ypiInxo1TkuabZb0xH74ctIA0t59e+oSx72DpKn5xbpwWxc0jws47dKLo1WbrmPJ
2kBctnI+K+9UkHAqgJEwNe8tpqAQ4Zs7gEWsbcTjoFzcmeVaWHppdCPkALYlwyJO
FdWSoZc8cgqCU3/shGgUDeJqXSZDh8Sjtn5EwxkazqDBRD6Nrex8fZzjPVHcRV+2
Mo1j5ykHIFyyT/I+QCVHdIT4njjYuBINndrFjeIH5QQySXb7Qht7ASPjTi1l/CFQ
HjqAMZr82yIl5WFMEP4vpSAtvYpKRF98kJRuVJfJITFNOszXR/9E7wgBxoOFFtWS
QmetW1vFuoXRq1Z8oeLNWhBVMbzH0hfXO+apoZLg2GkQ0oyZmUfuFNfwfSNUXcND
V5WlEKjpMgph451z52D7FPx1TUx1ig6kZPteyTIApTyo0C9QLYaLdJTNB3SeY1aR
S1GrCKivH1KNPAL8E94ealgHKgRbtMp3LseRM12ilftiwTM63c6sAhamltaopB7u
iLa7fAUFW0hjOi/vucgFaJjbVNOHy9KjV3dvANoh6G6u8G2Cq/GJ+LFFLGHFoXOS
LEO3Y38AXSe2iz/lyvql11y61WDyrZdPoWjTW4sqEtT6RUOxEVCyT/PaUmESxJ37
Ky/NYCVhFQ6rbyy3xgs9UwcBOSMuVcB8RQEQtPkn24VfsXjrrUmotn/5w1sG5EcU
o5vd1xBr+bvvwhXhlzQvahMjDLrGYXod8yUPUYbi3bQzfXipVS8JEL9/mtHWWMNN
JEZLwWM3waCJ5TMQCsgOC94e6mK9T/9yNKD5ejoAhJc2AgKCMVkWAokb9BU2PGZ7
T//+SqXJ9fprgucI7ePnWBR1ZiA6MnNW8Fid1mrfD4Q8v51YHOraYqjukXP4LUzM
i7LUpoVM5izmS/vwrNjlzeN6c3luroq1/mht2VOE3lCbHHlzS4/4n4Tz5C/02OZi
MfvyhT5mvcYVzc4+X/H6NUlnhNHPIsRNR6Y+lMPkmsR8D1mapAyT94WdyPPwCCX2
FsIjZ2Uy/cuhNMECUy3/uY9R1Fkr6Cl7IBGmzJLm0UZ/Oq8S0mlUStT6jkwbirjQ
CwFvEgqHK35ew80MiS7exGL0ax1XyYP5lX94oKib4P1bcmDlxpivburyhoZAqyqS
gR5hhspI6+F23r75qjuzq09wdTNy86UnUWdDijn5yOtV+VnkuQHe9pysbz3YQN+I
aamMDlOHZyzQrGqJ6L0uau+y4XT4B5KyO43J3KIwu00sEqvF8r0C6JhEMnTsBzp2
uVNdMh3NwQVCQ/a2xJbbZibbQNPZkoRZeRC4RGAJD/5Kz1EbtXL+5enPvjei+N5C
4s6coKl7k6tUp5UofdHTXJxU58Ek688Q1IyT7MYnOCMlmgiRxLREnfsU6VHifcwH
vThyY7Qq7og0yJ5Vub50/lgdg+VvNMIayRavspSIom76jdjQS/pLPazJc1iFBcdB
YzTV8cOrEjCs+BjynTwwik6o2ahSSNhd1KWLdtA1HR8ke1OjE7nvft/agO8MG+VG
bgKbppl3xQ7Xt6fTeE1HA9n6wsVI5x5uEAOmwGdWMNWruxjT9zdFA2/Un1zGGa0/
nZNqD2VROafSrNWsNy8HvJAR1Tc9uDNNxIvDDUix2r6f4nEylh/do10qEULRf8mV
i/J7+JPsZkm9065mZUzQzEIefMzdMzferrVx8uMlgkfBmlL6z7XKtG83QrUpcqLr
Uh7DfHDuCtJZppDRSF+d9zQC8JC/N7wosmu1y7b/Vj9mp18u/rPGrl6kkZszMt6U
lKqJk5UleRJLKwxhd2xFD31cNyHSktkYXCJb3NaiMzRu0NpT310Mx8Kq4iXMROKo
CXLSTFMASaimw6f8QDW3iax4GVH8qn/exDcntZESd6V4Q0+7CJDNh8vZjZaoQ1kL
Nvv498c2SAQB+jWlt624gkoIrNeMUkcfo9qFJhRm6I/IB6JUy0sZ3Z3eoimEt3iu
C4KASxDWTMNdKRgwaocc7ZJxv9q6+9Z6k4mBBLE6OSaDTRlPUYtstEkH747cArb8
LvVNDWaf8pk5lCURk2HzD0exuN6dRq28cewuJ3e9pRhnYUvTM6PYV1/0u6E9z9b1
LF2XN9yeSdB3MhGZ93YA/dt5Feat0OPMlXjZM4aCpV8l7dJQRbXV0TCJTKQhVRb9
1vbieHbDYaLrjACriC/bX+liO3RoFLy++QuODPPb5Qc97Wg0oRJo1NepYZXroI1Z
Wq9aoeEja6O44JgCsBiHdqpZoVClG9jPgGTjcTCM6LeyZomCuwJF3DFZBDCtMIKQ
VRA8QshAJu8xP8m4ZskDfU0S7+qu1nwQ4P8zySk0kodRVXqczC644Ux8UN1govZy
VYnA1mE704zZ6eD/Bq5Qc1ZaJjgKDiW1W+PaK35fdZSGYGs1OMHCbRmm/ocijrCH
9HGxB3VVL6Wz3XJpj5Z8OgxOwqqqgym5gXys2BatUq4H4WZl6meTooR5ujib5Ugj
iwKP3N6+nKg+P6kYh4HXvAX3j9BHt/XcVADwykrvG3PyZb52PYCO+sszYcpDvx3h
wiX4qK18Sf1lqRps0FHlB2JQd6llpNAfPGa9ZSrwL+0Vu4rU0JvKPQ0xLGXxxmDa
OLx+WBAjrbBoNihVzdyKKL58EF2hslbzjzvXM2AaXstuFgpfMVb7M4EFuMMSnXJL
KWS6j/BNqnLUGnnOqUfjDgO5rDL6CVijdCNaOAggY/VqUSXbpTiSPAlzNXovzVgB
L5PaBZA7ag7XhK97f0AFxzqxttqIGfH9GKnu35+8bScbKRiI27NFo2wpJdd0tIts
Kl8FcPTPyQHkwMgaDRAQApo7ia2Nd0890YMiPtoDVyWcKz5eDeMzO2iFw6AZT4y0
0dLichOYppNTiBYkbNiAZW4k7svwzCiWrbSIU754l+xM5Eps/ktlJB8BCEghVV3B
v+vOGxRbGZyLp4Neq+erpca4r614YW9sBH0W7xZo0052ui6B+Wsdp2KapnRuYOnY
YAtIUt/9NCkAvsTTFaaw30rjgI8gjTsdmfFQ6sUl7/ei3l7tZM7hoxqEl7/TVpew
KptK11Tooj2T388whk/m9yXK2yKEf3FMYVnDV7GvO7xDJUBLzP2BsM8mYqTaWHDL
W0Aod4mDJV/f1G7jjB4PgiNVllOveB3zG8UrO6KM+c7Uqlt9gPBEBSKrrMD6QCUx
Ekfk11/v5+NrI7o8PDRweGf7phlY1ae4yx9Dou92NZg1tHUe4h3UySSUkuzxPtUs
2a0xQiNCMjxwnLNEK/TpUkx/duAa3zq7QcvYiK0GRYFKuwEWmMHylxQvcO/RehKl
vcvcm5P/P2JROY/ddmGOUq8TjxKHhfD9ORKkT7KbkCrDsurFHsUANEVMlfGfMtFz
4kZfO+d9V6tvrbmq1eQ0yrKPmvm7YJxL/EQJ4lPWoIGZLU0F/1ymdg/psK6z35XZ
b959fjIJra0O5fc71iUEQfbXrSaKN8uuF0DYwsnkr0Youxlkf9+nruMk8zGP2bls
Kjqvgv9ZFvOoXGasNqHzm9EIxKcUFF3W6Ve6vuNNvRjl/4jC9LLKj14UxIyI9yAX
Zvl4nyoKkF3FfBzmyGiuNqO3JN+iVDVwiL2/A6NrG0xx/5V5u3UHs6EdpsNCAJWF
3C85CnYRp2Vq4+gY6XZNe0FJaSWtWiMNWUQYhlkOMCHC9MmQsPOrQ6mA7ZajXy5v
rPfqQthGAFyCq/BLUm11LZBoFCyMcNjb1BXzNv8hAtwf5HFjyi7BCpoqaikQcY80
4sLGGx9c9QoVlhbMdKkV4ws32GLJ87b6+K5cNYQ9FFjB7DxGqNjeQn0SibO81cyv
G6ApEc9GP3aHyu7eNe5DhLeO6DzClFLJVIDbuX5G4Vp/e4J2mTuPqfD4ZZyqp45D
iakkrwjo9zM8KR4+tEo5LVmT3h+94/TCfF2V2T+i7EelVj7oZgtzd7+/xHNafELg
GhSsT2ZVrfIHTcEozxCX2S2H6urw5cjGimAjj+I+XNspWKNJq0szmHOo6zKcUgJK
m5QVtBhjrCZdqFRX+TC7tvEia9+B5MdidsLk4AAiWdiA5NgkjBCrsXDFwRkgL2+1
kD9AipN6obvJ/2+27hYUx41V6ahL9eu8IepMg9I4xN4lJ+Zwq2/oPMsCp5D/XQER
alpvNBhDbzHrdzsddMUfzCOjsAstDZe4+rybgNqCDZrMEoL2Q8oaht2YgVV4sB0H
qB2A7jGTwexHkL6OX7r7s5bYJ9i/EPE1qsVtIYlkjKQ00Ya3iy485iNzimGo6ADC
WHx5Rfz2zX75CrsI001msQPATwPR+pxLWNjdSQXKt7hGUcEvt7amY+Hz1E/KaOL9
sxIUnLgXpsNoRYYwD8OasOPoKWabq5rhNommGQrqbOcIdThTiRanCb3i9F1ZPxal
9PEKpr+UjOL7gpVbbQn7MsVIwHlg3kldMftxDSAAo5MFW0sM+siKgHgX9lhr5m/y
vGxBZeDw+jUi+z3Eqb20HHLW0jNd8sowpzclLlFcYvyA2j1EKJYGllcOmP44/0G+
mCnx0bCSjaOjFbrmxYR2kmHy2k3bRKYH2IWQ724aCqQtTkHMnTAM4obWVwHzXKY2
U5FA/LE2TM7qu3EP7tlaJyLTyp66wOiygQTVtHd5OLAdT/d+fEsG7yCPt4PUow90
kVwNtIoOpXikqzVLxOwYj5jcjysqWA9H2boNPf6B1aBGasbl2Wp8WH1xW01NJb/m
kGcEdktEzKNmHP3zXvVK7KXSaUrfATlb4IR0hMEMkCcS1F6muUrimzmeUyaEG9S6
9bcRD8oJ+QMJ+j74XCA0utUcVMGXepZfWlpock2MsyRLe/7Gyt8D4a41n1O9Xq1a
xMn2+qTK1bMxhZ8+MAnuvzR1Nw/y6Crs9QMoXhpO1vcCfMvTHbtawKgwd5zfWxev
dJjE2aCIZcYuHS1pEPPIazT/8ysfpDt/pQHNuwuiXB/VY6jmMrCiU/66PiaQfuUh
SyFjoy1HxadB6vq0NLe3O/yBNs8OXWdx3vhVhLjSdF+j/wtdChbZ3NSUP8UK+Krk
1+GssNeaLGEtjGWyXpyxOXBITuYIi/OmIAm3HUJwo75PFrwScxoR/DRcIANUwCoI
fFZPdasFsGUVK4FjvAGtqXgU0k1kZ6p3DZ3VYoh4jC7HF0c5DNuQTYgZZrwizwm5
DeGzx7Cp8ur1nIYMM7Ca34V6Ye8AXhIJm655ddYsKt+rs4norew1zn23T555p8ZI
Th7xfrkBAtUyHNB97tnthAlTTH36o46IaPdVahVsUz61QM8mUfCnsP5ututiKWPv
2e/gYG5GbGiLoAMwCiGMBrMVk2vBKgH7nOJ5xcEro7eM+ky3I1AztEFM97+gLQtJ
9PIlngVo36KgR67IJT0nLnM9CvM5/uBxm355vWGlJk9fvqWjGOH1Uj4hHrquwR/h
3mhSF1jz/uzFIR1PsRK17/uR0LTe7Q1vRtf8XN10u1Vmdo9aahZl9Dik++T3/VmO
AuftuGIreFpYeiPwgwioJFlhodcTRbp8rwAz02bU9qlYlTrR3kM/yFk4boTrU59m
o45UldSi60emPabyd7UeSdLucVzISWijQXQeOv2ID3QjxPIpBU6/WyURDApFLRmM
xIHm//k5qIE0AbrXSvkzJt4mETAOc50dFcW/xQ3LW/0PgAUJeXsgRbMLi84mT2nT
IWdub2EUQeNcAn1ItMVc20yLVk+B1qqK5DRu05NVwnrC6bW3RPlUXZO99n6AL7d7
qeTv0HuS2oA0s3/7t5bhgA7LbHJIFA8uaPBcNsCp1JmulvrP/nTRW+mVWYrFyW+g
CXSM4o/PsqRy5v+vUViiZKejWy2/AYk8ZiSANbndJlbzvXNF9jaPPapPL9Vethb4
564I5jpy6yZcVIdhEJItogc8T7wcna55aiz51Hht52bUBpMFgnRjKo3k7lCMpLsZ
WCK0W3iEmT5JLwLkol9EMHvp3LbrQGg+qoDCgA8pIkOX3yB6mXXbi/dX/o6GSNNd
JnsyTKrkchXCSBSRclUeOgI6T60BRHGNsQVEfqUnVbaqZ4nar/KvwQPCnHfPdN4w
53LlvhEoB7aAxks90CzWkLy3Tj1w+qhFqf/qucPkkEf4nRQricd1MWTUMwmdUHj/
Nv0OvPoK9n8myUsAOuaj+npZXIlFEIMWqYg0iA+h4xtO+g5Tu1WyWKY1Zk55GZDl
BuLwI8QKdaUcAVNn/KqJlk3030B94ncHZevu31nQwEh6d3bkzwlCy9HZyCkb4mfb
kazLIZRsF7igvGwcuWZV+U9uG3d4cA45POrZw9ZbVf1VW4cujzeaJ9nk4sdXBE00
0ZbnQm4v076GGzGRxfzG6mcEQDBdaKz05mJ43ieKk1GWCtb7W5J6ndGcS4xJAj4P
csLfawmEzrLb1AREgycK24o9rq+NQ0r2gjmHnbpBTxZ67ogZxbwrWjRaegsW4eYu
HCASBbowbz2lYdMQPR2xM1GQfXiCSDnm6LepfvISRlaVaVhjiSsVsJaTTCcRTJw4
KVfuk9nSImhwZdOb4WIE8l7zYrdOoqlutNMLcpYfZ+PNdv/YsZncdesHXbD7TKRZ
llMfKpy+CvqxFm+SR38bn9CI/ji8mY+vl8YOE0l9eQhgj+n8CYIOjZda08981L4Q
VAkcqedzxaW0D+HAwlnu1vUcauBhEArFeiTG4gDqkrdWFs9KKIJvMcSLaf+DA1w6
X/6mwlFBMWMREEQIas9JNWmKhRr9SNt3uhSuaH46j9cbEHi7ecGhg3voCe8xUNCh
2bkidlK3+ilNeZMQbkWddXUPbNFYt5EDEehpKQ2RAiaES7MRNsGVHtxSm9OMybdB
yc6p6Vm6Gglqdvn6UM7Qc2IBd6nmZexUXT3GhoQCzQcaYdvRT6W4RlPdT5cn/uJM
CSWNELBUWEL767iNz/wKFlFD+yaWr5c7TkUN08ZLzzYvDFZmfwPzUkjbOeVXmqoj
DmYUhx5DHpMohTUDd8mEmtwCPznqkvGuUKb1VkA+fzsWtgVFc2jcxE2AIiIixMyO
zv7CzlHB6Eg5jnnawu3H5OBACm6CYnYGFLiiyureFxl0K65sGcjJtThipAtgQ0Y1
BbmfLkz2tRrMxMhgA6ICCXlmRVKKwn7aI/GhFIUCs3s+LYXTWEbfn9IPVGTm2z02
gF34mi13sJDei1itfJMGaW16aa658bAS+OhRtA9XQ4eKbXKdl0YblG41wDMdAcaX
kaUm4aj2gDAnF9WmiZ+UAoqJ1eUD5sY0UwT/jeP8RvSV86jcgJlhNJjJpfQbdMo/
0liKJXAHKEZ9i4H8DBD79WIJUmq7c8ah5nPvoVnGuMt63yMTG3tklg7BWysu0FOV
DtG058fjUSZ0wi/0Xd20+s4GFdiRs1Z3sYp6FMZV0C4IcVaSoL+zVFbtIoIT22MR
/xPavRGPRsjQHvu+d/KIKAy4XEPmQxXEZZt/gYzmQSo4CW1wvl/d5afICLgTOzra
cRIHO2p4Boha085/PJFANveazO7m1ldCD4L/jiN6oCaSLPpnvlLLLfY6JEJtQBsk
ps5QrHRPURPSV2DljdNpDe4lkBW+KKlHFjqrUlAqsYSQT8prOu2AB5ZaOFeyBVla
SGq8OJ0X2tH908iH5IkCWm/lcYWvAZYunY0onk8hQcDHpNiXboeGsyJbpnUyCfsR
Hs9yeX+P+37YveS5viIxF7ZfWKTj/ofIVtpDVl1+nOR20dn+3rw5EJXT4j6kj/h5
wYAsX4F05rU2HwuBXHf3+12jb8W7fc5DXhIYIw2lDzP8L5wo+Osy5TXBZ7HZVsYn
IfMGAeRR5InaiVa6rb9fhENKRV+56hNRvD69WcQgEahthM93AHSEfnRdGyLAb4py
mheePkBCn9BF/R4fSUcVJRZ/Ln9E1yZY5vMHj27fQkghbGHwckIJz5MFLPElush3
iU9m0eDRDeiBRigPG06Z0lUfgXw1czzZaJy7PZEp5BHmGrDsw1s4y1js+3ofnDot
nbF2vOZgMshDB8ddGOvZBVbAn4yKMOHqhBfFOorn3T47ywZoybiqygQDA2SSzntb
CGRQhdTNd82YXMR0NrNWA7XFdoE7UpuLnLguDOg66VW8oPSrVYt+jbfesLE5bHf5
Fg93LqOCjIhjY+8RXBqQIhzmWrThps2aStUgrGXWvfVYNAUyUpFC9tOSvSZyvc0T
/Kb8Cp3DvseptpN+1guLRi1RkDn7kCH7YnnigM3NF0bFLmMU5ufm4eYWuWpGd4RW
Tf97S6DJNAY1ymsO6oXn5I8eOToLu7m0StBVifH9snoN8WAr1WwXtjwJ/DquMjjT
9Z0FaezAgE3zlnG3AM48Bk+qdgxJpbpFswn89q3lw2k4j4I4c/YiU/9uPy3kCe/F
JxQfYOSYPFjiq1/i+U4iN2yoczd0K1emFWdd33YSTxOYfbueYqyPW5YbWl8BEK0f
j/hPpeLuqsyD+0T2ZgdkaQuCYsPR4tjLKUBdJsXrFLjA5jc/Ol4eKefASlacJYJN
mFSAOMKCyVc8s4TY8VXISvbt2qt5UR98Upv32EE8roeVvYzNVij/xbZirS2ST6BJ
lryijKpNIWLbkq2zOFhXJ35wgj0Lyp5esRpMuXrlgFXPsBcRXrkkGgGrPZxpaSxU
gpJwT/bc4/TTRRhz1XoZHdt3hKog+bsHRBEIoUkywmhw9hpxkKrziPTR0Rv4N3Ba
tNWqL7xN9KKqEvWrfqaFvGd6z0lnHJ953UKNNleOiR8oPt6lGWli2BbFd2UpOe0o
HbukXw3fSIUBVse9dEQt9nXkhm2F46684aOeOyfrmg1n9eiD7PZ6Am3ANH6wt3VI
9l01M8sDcF8Q9NDLct56iN4Ol0bxgoMrI6om08fk28aYxtETs1pPrhERep2Urjcg
Ym0/MqNbjxAjBtK9DzlKm2apHxMhRVBRckkP2oOTJtZ8mIHlZYcAToTDPaMaueQ4
iXw+sRZeXKzmxgRtpsU/NBuJ5UoHclAzH7Cfd2jun7sRBazpKKo2oKTMNsGWkNSc
OCgG30shpHhe3Lk7kmPn41A2T/57/hziS3M+DBPC+ZJdt13APg6mjH3vdwm7I1EE
QL6bT2Xz+xcmCpV/5XS/xBs/PJTkj8r0N8WL6jYu1jIlZgn+s98AyyB8/LeKFvd9
JxeQd2ghet5PxqpBYOt4EKCN9pB3G/UJcRTrJhPIuPlDi+9PE92uMdsHL7vnufEW
yhPyQKIU64nnkyeDlGPmnvSCM73SGADPJyUMaBzX076iCDvafCXFSJI3EhcfPkzW
tJsxEgM1gIK96n+yIemEEAVATHK0G6pwayNS1/+1Zkni/i4KkCKbgZ6DRsqFdrpN
YSn5xrsEqQzBIW0rId8YgkkHT0TSz2Ld8D+bbm0dyvPOLrrOjO1n7n5pANfnUf8K
WAZEsuwEZ6MKsxxGp95u0Ny7cIuxo01NI682UEpMyMUlFit0e/YcJ+A93ZVbYSld
41OINv2BcL5CU+p3Kt/kOpLuNzMEZlldKBEHEkwsiuThquLDpENDUL2NimEnDv+t
Bvnv/SViLm7XC8ZveG4eoJNDH9Mtr1lYPOnwGVYdlucBz/GqjEkNKXGicQw8J2n3
CFX7kBqmxxzi0N9jSzz72ezTe6ciek62By20vOcaq/UrNOc+Hem8LPcSF+1x9UIX
RRVOMlHLfSmJU7PRVpuJujMXaTPdgi2zel+5h0T4mMD/9OCmhsUNAe6Lx4IWHt1u
/qkM+xUslr5vjEtM70rRjj52f5LCd0/gf4V+5MNrC04F/PyhQYMQx/4g2qPri0ic
bLrZMp7DkQgYR/VbGunyKpUyzEuUvGf9ddgq190c1fRjdaSB3qhosr5bwOWID6Ub
ErpGzz4gZ+QapjnrDcIvrVEfi1C1QafdpHj85OCofPaHV6pLTeKRK8G+AAVsGp8E
5dhQFCkgC7iew4GYruPsMdnSFJQOJSLWbLaoR+fXlqJvVbsxssu5esiXyt6Hl7fg
d9TrCd/KubKH+V3rdoGBxWaAl663xm8vEe+6nNv2cm2ftL3K3/5zaCzp8RYoavUw
ayNFZmS5sPV8kF6ccekgwoNRpvDe3KXrn9WkVh/C6xcyYMp4GaUVrhbjFKXtiNvS
aK+i/sRTv+5qStNHpnun5vCuDAs+pbpvMwjuCofyyngZnQwkB/9Ya/8cgq3RS4tg
ALP/13K7zOf28qGfXb63Urpe+IJc0kF+DUnwTeNV0FSgxvJCBumJUzLZve9J/taO
6jY9W/IR+2jZcaKwSMa87I2hDB213mdQ5zaONbWAc1t90JZW9+Iwq0gLavCixg/D
aXfY8zUrhGdbcFp8e957+gXVW9OuSxq61oFZtx/ywd7LJ2wBP22uCh2E7ftqo/Wj
PMYNQtTUEpMDAD4KSA5syUrHGH/4Guk1WlF/XMPUtdvi0UQ26ldDdp6q0DpSNeda
LJ11TAHPX40IN/gd2s+6cibmwnMVLpWT9esPnI+9d6e4tuPcn/Qxwrxw1uzFLs9/
NQbVSkR28sdD9KVEaLvVShOa27AdusceghIkCt+HAJNVf5j4djqg4PcJViGgeoJe
jlS5YSjCQ1qlQTrRZfT7jTGXNKNZi6uCzOs9L9FNdJXFIVbAwZRuFb/ZZsLh8YLR
WXHKITyF/4yuM6rhRenQ3BNFmuyp9/xcwpWMdfZ6ug3yX0wqHtoJEsmPwQJclEPN
ICInQKupbeGDu5Wuuv3jfYg2t/nNf5M7hTBPX3HoZ0b5fzymDVNePZd28WrQz/sJ
`protect end_protected