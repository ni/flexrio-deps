`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4816 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhBNVMbsl6PTB5/ApNH6uD+DikcqmKlY6aIDJdxactegY
AxVO9v0riIv3Q5ik2YxLJOlL0IidSVjGCiQjzimpEG4jKXxzHibLTOKI+N8VHIjP
pTj8N+4qNvzj2hgWhi1h6yJ8Gtkwl2/jjWP1ZTjqutLaJlHJj+4gux7sVmIEqDOA
MhDx/utau0E/i7EHoBbXTvBU7saBdIUbrSe+206wSQCJ7ZCUmH2COtjSEmwIOtEI
wHO/LNSLvY4DlVGY8fmsjewwIGwuWVGHIHZ/eMxnNy1Dl0ttnbI4kGVM83h0XhtG
z3oMf86GyXPUSxe55O6BFPrTRWrmRMLG41JRwLkhhrxO21xgXUQ9FqotZnMmo+k0
ZEje9WKurIE9YqwWFeDpckKq0c9tbZXSxtgu1Jygme9V6oI/Cd2CVRVLhabsGszw
bKhz1kF+xgod8xIfw+vs3lSJbNG2bTw/p68FNcsNGqowDVqkXC0DmW/1jMqCI5qI
re9te2SedgbRVBBmW7oo0mGcxcqTiReSfdoUcqQN217HjSsmpvpyXAjT0CGK+OP5
ifXITMDBZsBuVFO0L1tHBTce6PR2bsGxUAxjKK4lsOmSnYtCU5eme1XfGed55gu1
iO02op5Y9Qg89G7+lhHDzqJPtD/rT3+dTFdBifEm+DqWj0x17smczdEUpXrtrw1D
D5cEy3ZOVhqezUU/qRA3CewTSEaGFXRyaVOXHb07tpBsCbcZmaVCddbUOUamEMF5
0Rzgqpydou7rpFu+k3vZlS4ss6bxcOT+w28unfM+qN8/plNhvUJH8N2JuTO3NiDr
bFntamMSvBTmGn7OkV0Gz7l8DGFO6u3py6vcl/8Y1oPhaf2ML41aJ9e73+KufHCq
SD7DMNfFq9cKoYGgGY1W9EHzBPUhd3SxtxhiKtu5Lt2d7efSY7NTzfXRswzE1h+M
YVMUkO7NeMul281af3kvdy+o7LSwBEm5kvWF6kj5dXr8Cn2gkiY8DyXZLt0wAzj6
uKNL79rUadvGnuZWzgWlwWEZqayZuWc9pxbecfW1AocCMzVBfZ7hFohQE2V04IMS
/2uilrMx1SRm+amQ3lwoXLR3uI5BO5oMEap9Aij/HEoFn59nC/1niRKmtRJH5dLa
f/V+hlgth4Ih27knVjStXMemPHSPhVXeD4ly8PpSeKdQxhW1/68s3FzI2v8gD+Hj
MGO+ZV3NMaEENtAoGwNyYlHSm8Gu2kA4TzaeHwsFhoT4ATysH4rTT6PMK1HfTSjj
B1yMCmDPBf81Xw1sRpj7A5Fh3iAe2YMXSHLh2UP4W2LzA/77VWZUQgBg83srWJep
ou6fhkzdziSI7Qm6gVuK10+Fjbw1EnvpUWLo5uEh7BFrP6bj9WnAMZT0bilCu/lp
n7JOcCfw2OMlJ2+nkjrlTujW+F4LInKJHvWI7iKZw089etx8Nk6qri8FFNZf3M5u
ZQ5HvIvjaHzEJ0gQ4QmO0aq+MIJebZOahY9TM5Yr73QIb/VGpXgYFEZozOtylhHS
x8IUg6H/UNQyxih/EZHOOajsoaSsdyJXR6dLgWC4XWoxokuEc1RTeDnRKuWBIvpy
cZUt3bzwik1ng/UAiuI6RBlIWUS7TC0Adm+OMFBAVi5m1D9NI8xwUSCSeQZn0LYV
lDcynPLLAxADdahihZQh68xg/jviZtUDpRwJAo58zWxWjvriHCxRZYaz1WLvrrIT
Jq7eFDmVN8qUizJRVOfh4BcVufQ26t4bEQpF0hABiyT8TRemZXSw0s+Fi8F7tyni
ezwIFFRTr7P/Xh/bOJ5n5WgegUMxrWGgAjsOLFYiRfFTdchtv57y1N6+doiJ04/L
pZE6+EQZo7RpOzVw7jxsOox9+OGoCdaUpOsg0a58LgWh7gne+nPGABvx5GsxXUoi
aNGfh/Z1DgH4MrRlsIWVVozc40Gxbl6kOk+1cCvQE0qIQhD6GXDNn1xeSQX+ixHh
WWCxveY8489aoyIfhskIDS7P6VgblcItdOS1Jt2FZvIVRmoc86Z62YqZ+/ENBihK
Dw9x1IPAOtUjEFGJySlV/RK/TuuiNfk/L2+e14mx+utBWVcWK96S78JXhCZlx9QS
rE84r/KaJ6hH6oIMV1GJ2GSk2+DD95ohvbZKpLHvnCct13zx+oskFYprEO4sB4f1
07o+d/hOkgtGEzrKaETZZbgK62jqp0ZEoEK89Wx2TuMXbdhTdyixQxo0kEi5k5Is
8S1vpP4gDHPO4VVEhHDQWa/UqWzc1+Bg2B3fJ9Xe1bv/OWgA5z9ZZNmsr0kmxN+X
N3DEsk6jEKi7Auyv9AZGOxWUO5GZrCajWZtGJy5eXgaeJhcCOytXq3MmH6oFxuOX
+yYsbtc9p0N91Qoq/Le5+fBp9LnKQMDIqsPxrySHf3NPuHDP4fQXF+4VzhLB5giT
JCryCdWmPlYIsVckdibahbqVbt3IIqMVsUVUihOwJogr02kU2HUBjG/RHoHbYJnw
BQdc6PZsVIYRcf7+tENQ9BtP9Nwt2Pg9csSdyXRmvEeu4pFsiLv1Xr9aMqWj7vY9
c+aNatjmY+IYMOgnf8UAlITWuyZWE9C6bOqiXCVEg7gPEx3O0wPXYo+PA8r5jvid
YgycwRluTzgCU+49dku47OmzwlITmghZ7zldjTGp18Ns91g7xw3naavzC9bb0Tev
3qrSk245zn5x9fPPKo7R2Oo5hl6ja2AYfkxhdHLJDmSQNw1RvXxC3p6pFctEcyzT
h3RpvL8BhOXfJxXHfWYD7O0vqE8VlT8jk3mSlk+HBe8ZIF1ZJf22AB96PvTDGmW+
U33zm95xKhCIoiEPR96WPaX//ed1oFgDpRkfvFGzwl+CKevkpG1aKRUKLXqr2W0l
Rsd1XxWuXF5rM4d9c3Nfy57xjhWP/za1z9qaYQzTgeptxvTdeA66rxbf69VVskue
v+K0JCy1icF/XdwZkmYgyQ3pw0/UqLz1PM61xBtoddVAXL4AcgLwWblZcJZ3ys6Y
vEChsM0Vl/IGprTekfhROFq91ssC5Pmyyx32xzKoy815TVqzX6wuxZKM9dA21DpN
s0u0bZWw7/QnxI8muLQXjn10brow5OoRyQoTnE0AsmcB+XDD9QGO03uLNW2z2O8P
Am8n2TXjFIKwBya8ZiOQTKBsIj0bk33eu7Em4huCK36NYgPiVu4ZGqNcOB0pNnOn
/mwnFUNNysrQvAg0QxLTc1O+TfjNwKWD8h3gvVBUOLc2Xe/EFSC7/0aUzGBk/wG0
HDPZg0ugcxIxv1YmXPFVJQYG69wBEaFjpTBTG9/VhLsxGU22iE9gA9e2rzjySes6
7zeU12vc7s6WDFRohZHT0AHVN3XhlsUi/WRoKa7JXp7c4TgBfxaXMt1g0mq//OqM
Ud4JYaiMHDzECu1bbSt82EN49Nxppwg5GEHnhK+GoyQfY9lQuxL7QINzRJdlKHHh
Ti+VN2Eh+ZN5UVixD/tYkUcBcPo9HKxj7vmk82+Ta4PXZPe5Cf6zlVv//4SIi8Pl
E0OaiLc4sxaESwPBtY3QJq0fpCXpsIxP0Tcrgrsy7h71TKITNVB0ODEFPJUUCHoT
CIfpK4GCGnNWzYHQT4/pSU7l1iyj/VuK9E7slyUlDyZH78HovCzGPkh2tV0WqVKO
HWSkHsxG2RY7rHf7KPZFZFx66vgb+whJgpANJ84DbjJYOHoOOl/RWoNFTVhiH5q0
7UeEVuOYcd9oNyRYAQnX9pUwzGZIAbijJnWGAJTlhro0y/DU3RHfaRNQxSey2Avu
ZThGcvj/UNVsEzj7BwJVPfgP/eS+AISc/b0e1NF1clG6xNBZkzZanFiKwOzDZYsT
zvLhLldUwZafmrDa9rMleYa6XYuxeJOByoiYA6RwU2lWc8hjQAslZTZYnFIYzqu7
aBNPQZT4JE6Ygbr+hnf3xn4crbIpm89xdOIA8S1lWxeGgFZEYh5poOfC5ObMC6ap
BlteXoAKOXrCvwki/JJeZLsMONw3u/7YO1Qs2o831wAC5wvxBqu492C4TWSCEzU+
Cr8rIY710D4RK3+WzYGqsYmZLv++CI9ZpwkRVGYwIRX9mcTZ1b97pIHXiUd6zFNl
oqrj2PxNHijZQqOvkVZFeJTUjWd3eiYTM+rvJ+JyDgRPHoxKmLr65fuXF/k/QHNa
PV/+Nv1vLoCIYzRRywbtBMJauXMgaVkTAgNI1QpEEHRLeFZ31M1CsF84kLMTHg3P
N7vRv2HA84iJ1LJzuibO08c36QTUi5v/Z+C7eRWSM50SPK+TohYRvrZfyOImYamx
s6SuasFhJdQCOqDZ7+ZPPuNns6Dsk+7By1ZPI5bC088n5+111Yn0L7so8UqnQYXj
8+ELzeZq5mdwcLk7hjIwdgfYAVCSQDIjebzuUpxLZzB25idPsQiw0wboziC8OcCW
DvdkQbJlNbqPS9qt+bLpRLXuHSRellVDDThsIGPBFQ/Su1nJRrYVddAa3O7wU+DJ
AkZPdx0LfWro9lxG9xxVmdAlZweIwocmSro19gLg8ff7l0YlgV2yhvDjwYPOm4Yz
lnGuHdBcGBnpvTaEozTXRQD3mBQSuwlp7ql4NUNJv6ITDpv+bI/WbcdnYddyzBcu
t7Qx8ej/fs5iYNfte8Q5JMKBZiyOIjBvwhvXsblw9uJKyc9VkHtzO28K+EocCQia
AxstXxI//JdiLP6RQNEF3qr1g7zUnHBNeMAYg2EIMAdVSvO6Ywlwv6wAMcLJ5Sb3
sL3isfPkXxaxsrsaO/M6jLT04rD4IlkfLtFadujLgtSBeQiU7enLHqbVxKwvmD7K
cztp9E+qqUbJsdDNYieJJGf44by5Qch6h8JDQ2ACUdf6rUEFRW0e+9ZEp9V0XqD/
C16b5/saclRwObpdywpxIAmMKY46DtBzaYKOPobr1LggT7ELIwogG9YnHhJv0wYi
wOoZiTy6rzigKmNT8pchGMT6k/lUisZ9YqUlK/abeqAg+5V4G6Dw8++g6M+QEMG+
6URGWlUbADFRUMBfyeBMknfJQTy/F5esUspyZtgrFTWxaTk9BIUQWERT7+nWWFav
0pRaW42GyTkD/yULVb+2P63c9/+Sk0rVwKaL6p6ebfoz/PIuT9LYn6bdUtehhi+/
D/RTLIlNECrMIJb19Td4t1X4UJGIfeSx+z+WLElgviTL9jfJJRgCkbiwrtABC3UC
+c/NLdS7mPvXIc2DUwzt/OFa1jLS2+Xc3qbTvUd86aiD357xbxe3pA/UH/mrmGWc
5jXwPyOgEahJ9tlXFa578SE2s3QAiHzTdulyKHsYC4qKR0IAU2p7IjjMHr2nvHWZ
gGbnWi/rarhuWSC2xm+lzxDPMYJkqMlaqN9qyAmtucHInO3PAMTBACTwklZRziX9
Rtln32ZOfR50x0iJ5WOWp3OoYSeiCQkCtgT6ZsRpksEiU21JDQ9YorMhWEbYXLEo
0BZtcl8+O3cNjeSXpE15HhfbEQwVEINKhO+NQPzBX9adjftZFgBIooCrDYHHYusU
U0Bqw6fPUiX21KMMRsTy8OcH0YjaJ5sBWzayN7Z+DC2dOlGslYOtW+8RXsbpehxL
Oc2yTYr2zQoTddN1670YmkmpiSpsfLw5Fzc8Oa4cm+zPOa/0VooLs7/VGtVeqk12
isvT93jS5kmsKCLuvGsLSrOmw+OtnH9lBwXd2mqYxiruoEvfNJFq/R1zWTXLyxwq
5HhYUsD99z0zvVn2bp5YfzZ6nNZu2MvfWs1PAAzYuB5SIohv99cVRUInqEUDCp8R
+ClGZVHS6N2n1b/X6byw5b4GTMpEoeRtSsq/PNnCUf226C8IGQmfRUt4Muzmc9LS
y2II412gf8jkXZ//PyY7Rp1p0cTgKzmEVU8CwePGeA/HUC1I5GJzw0ps9TEQ8z55
uaonP1zjvWktBPquwluaQM8mId/H6EIc7ShDP1Sg/18xv4jbVb30H3fD33Kd9FSu
xhD+l0xs7NnpZg+qlmqsCXoYbwEI5YgP4Wi8xQ30lFvtHnQ4TsXJcVHO/NxR+BvI
P1idoKuHMNK79cED+RG/SIvPy6h+R1LpPd6oQo8pMg0iAWRVz/1CQENNavwFzpvL
ABAlivdFmh6DTuwHczDdlLDhaYcfmJadB31siAWcr9GFfFPdVi1bHyWUCZ3OgWI6
EiV7uMHApoYxykqcw9Un1w2BlBBq9BClmZlhFg/fAyXv7j9HMO87jjtN9XunJIu0
/twj8DT3JWyPwOYqqroJ9f4XTwNP2DCJzObFKWT8d3TnBrKdDB8WDKWmi8ygMx08
q9YPX0JvhcJofIrHBT0NAw==
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4816 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/T97rZhQva68T7JOm4bkq25
b4BW57ADAHEm2yg/Vzsfl7TOuMe4xzV7rdHsSWg325uIR/ZdH9u5yMIWipIMzSW1
9S6ZrSagwJA3aw4LVbUV2EwlMscfwDRV+nfP6la4H4ufcZz6rGZA8SOP/DmnmO97
MtyATwuquaaXCQK8SaHCpg9HuY7nAUSon4JxEUn/T+z3gsg7huk6fh0XTG4G9emT
6/SpesXZ7r754MGWIIj2vtJsJ97roS43XpkZuTsIQdyst6u+EGqvHkjn1lFki0xl
yxLBN/vzLvHh7Mr9g4MXvuKHjnT05wd+X0J9dp/dn5Isecr5XkLVc4DdWqAi4XKS
xrp9QEbR6kh1GNv+/oVlQZbwUlaKpVVv64yf/6At5QX/cilDfNPHAp+/CDS5/nNf
VMWgET8rvVajafoUV5T7MuxWXaemhwgG65X8p8FftfsNXViVyrdA/kA3fzQAN8Q2
mEVhl8yyzk5ZJCEM+4HvCc02DK9+udZEyTuhVKCb6Y/6M2wR6W7cJkIwdkvmXnHE
oTIvE/AtqzfNyNn8PYX/8mBEuEl+P4suBSxa1nsyPiS6+YUFTgTQH9pBk8LdS84n
iaHw7teaVhApN0i8Sl7utbded86SlPpDjcPPN5CHbjjUxQgeAY67bCXW6JXQIOkE
sh7L9AgUNeyH9dpfkNqFDWezWb0CQj5Wqt6YuRWiaXh5n9gFvQz7HrzC0tdGj9pl
zbMhThTHdgeSxP4/whtyB+ye3nrPVQFtFmGChqMeXOWLeQJiJ1skAmlYNh3n+jPN
HPM8AOtv6dyil87g7AGpFSAevriJ8px6lZYaKT63plsElUjcSwWrla3tlSwuMaOp
f8oboO9yNMZ3/rrb158wex3LXM15tcPHNDY5+4Jvj8bR94rF97VCKtr+OhcbQdJW
xJN85exlfbIj5EKUosw0upiBG9luK1tT9JJ15oX/a6dGA/nx9PSJwOcG2WOXmxy+
9qLKV5yA4uUB2HfOrHfnOnxJVV+Gm/Tluep9bAQsFf2kG5Or3aBT1y1yFeFfDhJ4
VgeExWpn2z7gAAAEe+IYMnRpZZMhZH59iYxVBdawGn2dUfKdZqArrx3eLJhoDz6w
gnqUxuiGVYx1OnzdxBxf2gWnbsLOilUVZmwhqQosnPY1afjJMI95xUkfvtTTq2aA
rix5Nc7MW9IUNJ5bPRkXac3itnbPCmGxzjPZq3B+KnovrAKRrGfDe1tsUmvqYC3a
99oyBLTN/rgccCX59wibZ4/idDk/BK0sb6lG/kqntwvTPKPx0ha8D3Jxc5aVZTqU
epXkKrq4phgP0QEWZdSHiCgWKbrRRM+C0StkVbyLeI5moQVDQRtVv66wvTLKaO4d
HnuGbD1lkbYjA17QD8ezjVL5BRrDAS45yoOKBdKkG4m2IS9Y/Tu1FdS8lV7/eWXc
JOGsWUfMmfFd0i5QFfZxDGsTr0zWJG5EjrjF75nNTO6MsnMClGX1R6Q+xX+z3d8o
p6+hAJ7oX00DH3v+CgptIFJ5/o/Oyrkrhz1z3lMXOAC3xAE7FvBXRo52LZR8eBqO
CEckEulGdDZFGKETGHbD3X8El9GjgmIS13iIDgI+fMFZTkGnt521wakdhhwct/vm
tF4wH5G+Xt0FwcOfVSkar8YCB1/lAzjqwM6Rt22eiuooe7O9JfszHroFdrufd586
FmqR9UlYddbickYqJkBhj83/7EqGq+Ah8XkfFx5cfRGPYUNzNAzozS4pr9idVQmn
mWK3Az8EgsTbQOkspnKZeCANK1gNt220mYa1o6h+rn+cJOkDo8CrJ/CbAkkMX8g2
fdhNnyqxeMmXP186bcEndf1sb+XpvLXi9ReAmUypJSEEafAAuZf8B5iUnp+wxuix
uBtIjpQBJzPYbYNPlyQcJ4WuP6F/sEtlWnS/SnYAvE41rrlRDwnlNJNUh1ycqaSq
uJIWTapFuB8aQysg8plLawG+TAkvnlrLcvyVpRKpiSGVu9e3p7RlpdLdtGk20oPX
cLNO0IBKzzM8K/q7thDVcw1RO1mQqOvX2zgngwAJ2hVSMLb5wezblnA45tOHxvWb
O+kiAl5Oq/4s9drMEGlo/h+GJmg2Ld1hAM0nTaQ5b4b8zDnEGh51ZLjotyfdSj+/
gywC7RA9kftkQ3zA2UQJyzhJvi7AFVP4Q/lIe3COL/0i2VrsSfv0ftdYqFavwCRN
Mu1/af2wVE9cTM5sCU0F3BDcCOQ9It0jrsI3UTziShASyun55X34UMnhnu2yw/+v
RrPs4L2+KxuCaiZTezczhFGAT7sfWX/58WYqt9Tubva68YDXnTrhSOw8v4TR1tH8
YF/pB2zxWsmOE7so+rSrO6hLopPAT17aGx0YjzUID3nKGRccr2H/bblwkOYwhWGS
cFTV/g5OtBGpaeTiiTtgcU8Ok/x217q+rfCNIhhwEtYPVDf4djAS+7/kQTzAvZvN
O597wRbCcJYTNn90NYDEZta2MuxbheJMVI+k71KrAT2urSE7qqTxrC9bQvgi+veD
1pZXLyEdPdkKvXvYLrwyZvAMTMXlOubTIKVi0X2oRM21PIcNhbmddvwSstBZ6XZw
KoEn+EYxjZMUx0mcJ49eb5kugS/chGcKtWKrB9dDHusEAoZqyDchU1wDq5VnNivX
DdyOl3KGtEna8nKEvaS7xpOgXSGel5zpzRSFtkczPzvrNzUcQ/W6dv9dI3yng4sg
EwBKexew/am1P/wVMPzEhLsES02Ee/zW4Bz/mUhDiHgMSm6CG5qydLFs+ZiNYcg1
KERDzDKgOUw7o085Yb7y81DOZ2sOQf0EJRc5GlNXWcSOgDnW1tC+l7qdLnKlgQ7R
S2eYOvGHAyPC3iwcsOxKnyvUMmhtmLw7U2gQ/IrKqwD3AMawhOlNqm3pIxuy13wc
p0cgf90eRVcfc76RIIesx9374+m4d9FLyPFAk1WaYHtkPtktXdz0JOuPqOrv5PsY
lJSyecIMoPTTSrHlPvZwstrJMvBPqBUL85XEWL6Gt6bknYds/LuXL6Tv5S3SnbEZ
xg6XgHUHXUlmaf5pYVg6WlDXh843c+2n/WhIeKGAqBSEiPKMLAj2sq6qjOtsSgZY
e6g8rd+8S/MwiyV2rkciRP8kaT1/2qfU+bvpKJagvwJaKeqq86n01EuCOmJMWYoM
2JqCN0W07MOSCo78M0BuU9vlGiP1Ri/O2DhUGxfct5Hghx2/MIin1tM1Y925ZQiI
uaAR0LJpXbk1SewMbgrzmu6uikQKtGd+ASwGcfN5Ehc9ZvhEe/ffqRVWbZdZ2RBA
2SIwzKzwZb4rAcdTEK/IkhfzYZYlBtzO127bVnPbG8zqfJAWFnJTqT2nz+Sb9nfb
5ZQw9nnWuGiEdmiJNnbfy5F5HDR93OLqhLJTFfteZL8viYGTAGoM7IsQR2PX+D1q
G1YZCjNRVHpFJOArqx8UrdsSDpCMXczu9Uh+sqOkQ+s6D3dBrm140oqDaQRsVDwZ
UvcWlM/+6NJiATl7LYEbWX5S5/tgkz10ZJA3hPEPMzLynrWA2JEAlGG1EzsUQ5WM
8eKN/gNhEZQ3Ukz8WFeZQ6p2AbqDAic5AonfiwzKdyeEmhiYE7FbUFNYvf2wsezp
dAr4eoVi0bL1/uTDrS0xSGZSyE8EKBzyRqA8qAfECJRIKCafqDBHnZYYuZzDY8kH
qji6FiPnoGle2+Pcf0CuoaDiF1hnTNEwDeTnuatwW0rX2kYUBDCl+k2VpSk2Umt0
AtqKmsxSR1bccB3A40EpmEEIXCN+xOtePR+LqtkA39e3lm0b/i50/o0xKojSXMDG
giRLinTTmznGEueAPZFarQ4aMVwS89w5jRsJNVyipdkgZtkUDNqEdjG2dGsR9F1p
0jWsyZSIH5HjZIu5sHeTxW+5gXTJY4rZ0Iy46JUXCUjMqZbhH7zWyvlCafaZGPdr
dq7D3Rm3rMwvdBZzRijUtyQNjoywXA8nYYU13irx/4gHBY9HJu6V7V5E7YCQ/6fb
tjOP/wxz7p0kbaYynU60L4OZTRiXHjcNkfl25nflisQXNWeiTBq1yXYzg3Io6H4j
VTw4U++SkbTPZiYmzGqG/M44mTqqaXE3j1Y1cmpg2i2t5o+yLgb5UoMmFUWc7btr
D2PuuiSbaJ2yJfKe502S7sPe5f16zGxkagDV2Bkm2Mzj6JAd5N8jl7nQst+m7f/k
XZ4X1tri+V8p2InYMh2Aum392+uxGdDNLV+ZTwvg/pEhpVv/cLjAugTIO28DpYBx
GrYQiaAv6Ou87byQThXYHWneApl0dxHwDEcrwL6WwRtpjMq6Sbx6Dz1XSm9mBe4r
sQ7TtePSLT8rIfLInfEEIQ5BtuxZobOIdIyFvHsuwVtlHNIogyFY4qac459LkcaF
6x6WyN8TedsPF+BrEmDSxX894SNrbfDLqc3xS0QyHyasVv70OSA8LefyS9roisHE
XKkaFklUjNemFPXrt8ChbwZhUYUefuf9JDlzRUO8QkLFLTr18ax5y92PLzRa63AW
emupsaTHcwOmabjifRBhtia1e/1JFm1ytB6Thz/pBUwIC3xXxaEU09t2gVW11HEP
GFzKu78k+diY5ZmrV7GzIARI+NHshD2GHgr9atGaOhNrdTvjrrpZMBuM4vhqysVm
btlZg+rgNUUtrpZTZA0HR12K+OecakI8ClJcSACcAyIooCxIAKY2THKvnPG+XFJ8
WLpd9ok6AoSinT1XtHipdr4R4aC5Y8GDP6CHfXoOX5UE+6dgdEU8A1JYML3p9oJk
nKIpoww0HsDP1Zy0KjM0q7qeh2iifSi9rk9yBdf5P5qCqHNmEAahHuBsh/sNAxBi
XS+X0/riKOt11CSGnMYYt33FWf6zzN6OAwPgb8oTyJLOuEDfVnPkd4KvvgbCPHzK
7KApztPyDXyzWaCzBrnXbTK0TrqJvRnt+0IUMK/t1WXbhK7oX/bk8ZO6cZuEiLKR
WBm0ep9qH4KyfvxGMcVkgbklg8gg9ie1fm9zXbLl4X0mww48JocsBPMPEZ8TJpJY
srsmSIdRBcko9lcpFYTF40JiN8MKea+U4E+uWOFu4yAvqk/+UhFRagtqRo8WVF2O
4/KqHG8f8LdPUr0gk9OYA/Nh4fh6F1zRdgF/a6yaZYgonV93wvSrIcQP79Z16PHk
EuH5jmbV1HXfoZcGvziOEuEkuemHnuJAXnzsctu9+q4fgrQ8uGHOYhYggQ+BEmxb
D86bkj3lHWAOjdjaicO0TP/YM9kn2qGMIzADp0f7MLZZ5HtcONp6OH1uK9/q+D6D
pyvU86EugrJrfBz6QJu/xOzJ7poeT9TUprgV46uiiyaNvrQOardzfeBzJAFe0lk7
cEcO89mRUjKOlTHL1Zk0CbzZ5x9r9hag1Uz276pcc5qcRE29ckMXlSwBbiI8DKb6
sl/wC+zNX3qAD6hVeJne6ShaAheeWhMFvGGFPEEvhBV3QHubuJ+d+dqLFtx1BGRK
R4u6fOcJEEUTp0fJXJJzLoehGcmzdPX2rnwQbWEnkkmq9ZnK1mrm68geFKYys0nA
1Hi4+Jlhxy9vkiQTfOeZOHnaUIhouoMxE209DrNEH3ZkPklYHGCKTyz4qtxd7+ZY
wabibElUeE4NuFllwIqTiEE6Axw+DTGlp7yIOIFDFJW7LmsTnEfJW+NHJe/xJ3c1
xk225xCrhLPWCkqH8tpI1O9SjI/whBXz8880JxQGehQ5sMqj/Oj+WJ0dQUBX5w5T
x3VvufSbvtGJ/+i5h+J2jPPMim+1NvNV9StzHsoMnJX+9LtBpSl34eVEEapwjk0T
vy3dDp0cqze1PbvYWKPt7xJJX2sa2x6hIY09BMR2VLYckJCnsRnQa0B+ftYxMnvn
nqGVyy4eYJS0UgpMSP+r4rCILpWqDIjGrRau2whGFZfZcaYa11/Khx40sVWJ73T9
QbTvrwLZEKta66yhuE8YMyxrHn2GEHqeD7Rr+3bCoVB2OdCdIooUtydwxTbDyN3t
tr/V/Nvk9ywxwXi4qLocN39sWfKTURWVAf1FPVJ+o4L3Vkp9oDppWkqKcEG8Pizl
UMMdMT1VZSdgXXRfsqjuLnh4/RPZQ7zTlbKw2z+5TdB0KW8/ylz34t4oSVMUqUk2
HyaGTl0rllpXm2nSnkkWfmI8Fyw9htxdA9pTENXqieLlKdvFvJb8a9MbEbzKq9Zo
ydH8Gf1+ZJL8HnuLUPj0hQtd9UG38Iz/eYbMHuzpyYMDQpIhnV1QURySaSYZUSUX
auNyrwT7wXaZv7GIxAk/Gmrn7n+SjNGhIrcwFqyWKe6bCeGL2Ygnod9KFVjNzfsn
vNYXREKSe7nRib2/mUFEQA==
>>>>>>> main
`protect end_protected