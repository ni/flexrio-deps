`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2320 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
MZ/g83zWCQxCIBtfOHnYyf1Xbeq+ur8QQXlQmzDDF3H0wazoy9CSpgA/PphQrYtt
qsVTw62ilrjAEya2qrMYtQmOWHeNwcqmVFRj46mR84nbmzFcsb11Twq81vJNExdm
BljMLRZ++ewNImP61625/gHK1ZAkA4iYApG/MbW5T26SP56FlN277MA73FOk9JAr
5CjHGJ4O23a18xe7ZFTjrh6IF1KB0hxji9lfghJPph9zEZlCKG6OKSOfNtZAIA9B
QWm9247/0eZ0GbuRfIAzvfZ7piWo5NRLclO68mJJcSjAyX95WzXROEU70hympznF
n8Bc9b1geC6vKtu14G0EGuqp+5tJzt8f5qV4MCUaQrYpzofLnftr4u80mRKA2X+R
GcLCcmKNeEe6baAh0QxNhGGIokz6P8FZx+MvqqIIGZbz3Hj2gULi8HWshKzeJAoX
JPQkCWDZc5T+NBsZjd3fG9K4oZpRlrR00IdK1MdN+uSYwjbqHVGUFiJx4xwYjdyb
bzuwOXQyBQUyQ8/XJkBNlzwU4V+6h5PuCNx3m6Xb7hnX09+0+inEdgX7SGD+fKop
9wKuLskSUcW1WsYv6grj+8o1GJzVdcUC1yzCPWpkgRjrJuyPK5tUup7pnolaS//h
b5+6SwHrcNQInH9FOZdAVrd0Cj1MEtQ8hLhg5aJOg9CI4/ukflwu4KvcheCIO8xM
DY8Ma0uBYwIiN56urufxVb1Z96gC0UG/EdoBqQSRy+F7DzqnWu73XeQOYDORYQwq
hAgL+RRniqBf1+rlD0yYewvpHWZGquDKXv2QXKuUHcna62XCvCu+6MxkFBcJw1j3
1lHqUaC8qTxtcdYeHVBJJRiRwEXg0qAvRach344wCU/WUfhyf5yWV3SyARYHrJ0k
J4Dq9+myk5LywR+FmTcSUAeotFcVBYKoYehVVCp2qQOC/2h/BiGB1OGDLE+D0JGT
u2iiH+wZE6gjXT60wLTBdbWXKNP1Mbl/TzEsliocjIeC5p+phwbyGUg6DQRDO0jl
+lGR1qGzgHolyYzdOvaJRi/KxmlH0/grOLFsE4Alu6O4QXXje4+Xlg0mKrAXySJ9
qpsoyAZL+HAlGtQOoh1Egqikp8v4CR5CurbgAPRoZPmA9x7tDFiHm872bg3QO30e
G7ne8d0eDldDAHCCSLUrVzT2Xuld1gLsALGhpdbd3QSP7f5365piXXtm2Jo2e5yB
iz4UUIivnM9NowQQV63X0Wsu6i4jJayscJ7jf5cCVYEf+lMbJDdcgtay5nyuCFVv
+MZS3o1VoHhfUEBMqgrcuowuaN1tld7FXc7FjrE3x41Q5MlVEFllXmNDNKj2Yq6Y
wFi5h0oydBPyg5s4axSH9dW/cXH+ZxjCXnINLh8hNr/S2ubLSrJEuyHqEvUmY3MS
w3xyrLvcHxd1VTf1nUJORgeMZgEPJrVviJiunU/2tXspRm1jcQt5151j7ZAtxwo5
6eecAly8ExsK+5DB3QbcVrL0AXyZlg7b0ABMmvnRlcthewncFVB7ZA6Um81OhgmD
Ef+bl/3mnG/9DT3OXHi0sSIQw5RCSlCjiGoyCxxpfJ8cH6S+LKThnRKaSXlpTnCI
aDdJmH3v5+kLBXLlClU8JcAdyQF3dUC2EIQLDd0xz1JTqigp4VJ8PrwJ9SKjPyUn
pBetEX7HQvvHOa/TWrhiL3c8m1ieueXiElSvISb1k3CezRAEgoaX9ccmLjVW6Q+J
UrdLLQIE9PRKFTQgJjpoUhg2mw03QLLCDi2tA+ciOWJXO1qItfltiVnae/w41dSd
EGUfnEaChgn4MET3Vx/2suC2mzpnL1HdBrLjW3euEXHkd5TNyfEt50gbI1vXsXhF
9KW4xxO8AfQ6SQoMDinn79E3z6p9GbHO1ZU+ze91wKMtjQiiBYE8Z7IHgzqeHHEX
6X8MIimuP3SMCAot5SptG9++Zh2bwfSXeOUcqr+edEQwMowBP7yDPV/GnpfDB55i
O6HVRs4T8658T0wxPXkWkzWc4Mn6c+nv6OrdzHPXWP1Mn6kolfP+RQ1Nr56L2C9z
B70pLarTGtNTkM6h0BjmyDk8oub1sbXkoCHcunS5KOaICMbZJ6YzRXCzYRUMLfEG
c72OqNfk+XZMAHZiwtddt2h2XcduLQU5IirzQlq941Zwp+rPjmVb35a266vygg3h
Rh35ODon8AEeV5OkPKWKjK+tsWo7jDz2l2sLGloMpUnbwiaiQAAZvCm+HjAI2Thv
eoPGN2dhU9x8wcn6L2LOk3rPHFmw4w1bTBcuR528Bk4fWRf5EGpt0zs68mlc5B0M
o2Le17OP+zETIDz0ierQYPfC1oJyM2oY6hSeKfmveCK3goFuwhp1isTgcBg/a2ZL
RnfjTLDx+D8JZrXzahs61/ESDf9AKDBCNA/cBqhybJzyyn4vVhfllpA2A+cnBOak
g8JDBWl66etbOoNDEPZd8WeC3NMq2VvbFCvKnrASS1fZNViKr/cKqaDcoZlBQod4
l5eH7G6lmw+esGPT7FGBRzjZdIwsgdGNdF21oUMS+SWBdLb+umljfeyZupP/N75H
HDr0nbtz5tdXJOH9tBpwzp5tP17YD6CDCfUwaBfZdRbCs8AlsjhbCh7KNY9VGU5P
ZijTlzh8j4LuFyRSL/cq/asHKkEU+1mBaHBdn1jhWZWx9eno5+0GKa52EMWbGv7m
mmXA6MkgFNsC8NdBF4KdwnnOttjDqkB2MYTKHGnVryAbAW7ZHetJK8FmjWW/RZAY
uJ59aRkZcKgtLCQfQJ8TY6894Oc0K/AlfPyEQgNyYPCm+QFQpINEnG4CdliasP8B
5ATHH86AHyoZrxdsMfCFK1thZtmuYnavOiRl5hyejtmn4Bts6InyVS4dTW+jJeFm
5ZUzuk1SQwir65UbXSIBdnonAFmuX56Ibre4GBxRNU+prQ1zHQkdpYfcFYHuB4sE
8KRzXr3BxTGkcbTOpeTsPA==
`protect end_protected