`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 27696 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0gQgIG1mJzulW1XOK5NnZR8
C8XqDUtXW7uOWTnSVqbIbqEOpZKTOgVl77d5PaqMKeZBiczeCj+0qA9vPd6eII0o
DMQzg7XbKyHiDlO/gHStnRO68LnC6ywhPtJC/S9+EPHd5MbqCe5eeyBOVnCPo9R2
XZhRDrsGEMz83YyoHPFpSq10qDFcZWzuMjdLAunBl8NRWJZXF/P4WSaxOKBq841J
OOQe5jO+rnmMpOjeN3ws/tKeOLlSrlU2fMHNAOuQwwTCuggW8F6cDDhKkLJfvmgh
rqDu8nCbGInzQbk8DRPC+ZhRfyfzzUf6quu/KEQsiXSRGZsONlbeYpafDFoJyskm
a1jrS+4irDmwFSD7wCmBq1diQDGHlh9MI5TvtLvv7cfbZGdQgsV63v71FOcZoJp2
mEnHNIRjqmCwlM+pMSG93rT+Ot8I6V5bPO1AeuUMDc3vGZYNEw6Hhs1PLCm5vIL6
BkJHl/9DCyx6YLIrvIWNK9TF5W5TcogJjkuYVhcYydaMWzgzPnRFOuCps+EGwD4u
NfnfhFJECozHInttDlE6NgoLOGZQmiO9QNpwn9WNyvso+hYeD9kvBKIYq92DWhJZ
uZZS0IVu0kzXOTmlC9eLOkFihFUc4uSYgpP+pTxoTILlPqwvdRNGliBSOr8RLRfx
c6MOXL2Zw8/57vY71bZNCvxzf+E7FDo7kwsaebFKrTN1yScxvu9sbHnOU8bm6iHe
XWg90Pe8/Xz0NKAeWTnk/Bt92Morr8YzDdGmkwXZcRLtJJOhqO+ej6KBMAeCJi/W
x9IY/wR4GUiUkmJSPUqVVd7hIPCP/85grzBM8HPZ87l7joPCBgEcHMJo6Zqx7q2v
nBGoHOXYSIgL/6AVXwQJN5ePxE45MDcYKniyCNPRAlL7ei+0yxKcrzBtCZ+zAAld
llsxOOgWK2NNpotVmrb+tdJ3xHeUHlqNHlsB4py7vmCA/cVXL+862PI0uMIqwGbG
M/uJbnhw/hEzuv1/vNErQ0HC75EkPvVJa1RaBJJISylyxO0GEhYjfMyU1XygQFX3
xTHQ+QYhF3fNJtcwpL07MVnaaI5C/BjEsZvBRWJQIv4V19633cE62k5CPAT4i3nV
wsgfXgN7VMSrE+QvO929h7MD9gY3bAAu9RmwWyvXyB9fnzaZf3H5IVKqoL6kspNo
3fOfl0MRhstquoPS9EE0neqA+LFKmLyNfuKEuSWl1pszG9RaIiEqofTXLBAitsBb
2uIrW1wencSc3ZkHNhG/Ppf6wTl9ppKikXhL7/eTU9gt725ZzLhvq5cI4h3b+UzD
K2Hw7U/gqvVmVhWpHO7G3usLHdMLd71XWKP6zaz1BKCYle9kh1pTm8f5GkU8AKjz
l0bvzDik12TB9pPq58F8O0G9cQHWoFp78tiWEtEpZ8+MnwpZFReEfRqKcwQ/IIxS
mHU+oNM/w01uDLqfb9/tDlqbBNc694TvHiGA+rX+o6JYtidfFLepnwB+Bj2U2bWF
usnD+LEj2UAInh/+PUKbT2WTqzPLGyOfNJEJBnFl27PkjnBtCtctaH4sp5Gl8Tio
zHLgkTLY/bN6IRCJG+Ud/aPTyci+mIc8yO4Lprh/QErOJ58aOVJdZfFitJ7nqwhS
YVZLQm7xpLTuCbn3R/k0QIcXlLZPovVxX5Qh+okx3+mLBoQ5n2HirsCQi+kvAPdb
w+vh48Mx8sagwfoa+T3yXnU8PcOzLwPDu1bRw965dmzd8fqZ06lDCCBnME/AmAt0
SH9nRBMZuHboNulRJ1HDWJ7wuZ6MUeVBtNYc8+jjZL7tK7rzw9GLT4TPMIITZ/oO
MVT0sfu8BrcADYrIymgj6xgusVEyly0KEH4+0UbPYLrZBP4E/h/LuH3z12ihcvZb
CUdbP9ANkWorFV5u3sRQBlNWL3rzDLQlQcbFmtgRWwebRdk4PAVE+G7fEWe/FHZ3
GQsnmsZqmKiJsJwItUlpcuI2xIdSZqJvDVvrJEMi3662+g7mHpvxfTLonHTUsH9q
EGcn5xlbAL/RNxbuoRMR6oWDaLDcQykSyUZ5Z79Cp5cn+AcUW2ERZO80fekOnXPh
Ele/y/bKCTnWFIxx8Frrux+lSXqywf+Qlg7i98ypZPsldv6s9drQlmuyICy/Wput
Ut4BM3fFHyJCAdxpwWJdWUAtREZ72sT1H53e255219U+fEtO5aYkHZ0rBvfB9/MJ
sLCIwjAzMR9ABHkZpbBs0jBhY+KYBydkuj/uNsDq3R8yZrlR4c9TYxWr5dx96kEY
+hHqAxP4HUJ3TUu9iKEJwF/pH0gUoWv4IE4LaknSDSZ0bYprh2VoWReqf0m4T/Os
mad9VWJuVOezb0VEZVWS1tSgFV0E4Y2OKe4h/GrOnaaG/5aek3FKZHQT2TiWW0Wl
Ymw26S3znGRfXvDpM7KNO2HnYaq1NwbxZCo0vu1+MikHWBh/B79Uczx1jtDBneDp
PWFE7egic2PxoWzuZUZXBasoOA+1Ky9IMjV9N6tEvUJz1xRm+PbzfASokENuL2xK
rzOVs5rtjiZCM+c8pMp585lyIXn410k5Cl5CL5yTF/b4VySBjekwc21wJriE7hxT
UsqZKrD341/fWLkR4VhlBJNrAFyJurvcV1Z0S3LQlTqOfOYq3CPcvPqFQEBtA1Mq
fUWBVsBrs5hCagWMY014nQMp2H+wRT2j+CbEF7+/V61sVZxcZFidvPcohRcaRmZQ
emeT3muyoPCMNjh9MvDg2ZD0T2N4lp16rvBgzqc4A06UmQh3H5IJ5+Ovraqk1mTn
tBm5wmydGpqHd1OI7/CnxGvvnOC3sFW9+muUyYbU3sJhTpEkArrsT6fP4hI2dGIt
UbhNk08EdOGbMgcoHmf2XcMHJtMEmqCMpRoGSOjZD87hv+8ZIBpl3y3TumzXWbdF
YbsdkIuobv/lqhToH6Wp3Y89/Kke4EZvoeQ5kAglNckKGqh/N9cCjSqzd/ErsJGD
aB2W2vbqKCbd4v1pqTlGWQbmENya/XFzs7zmymbYIDSFiMphQWkRCXaHhRlvecbg
LUY0hwQrpysDxZ8lnDy+0iZb9ODZJG7NmOizhogGLoFy1UW+CjsEhBa9r1mnxX33
yl+fvqWWAPRunPdlMZvAtN5geAUvi5keL1+vI2XV8+OSonCCGAIHKs8BrDntW8zb
cqCHcScfUUZay8Sr4Xqygn8i5MnQa9dwRVRsOdnEusML3NdhmsvqVP7PLOnKwxXJ
vauNy9rxgpc4vqpiDO8S+Yf8fHzw9uIaqqz4VGNm6ymljdJpj626gqMBVS0phAP2
SnQDk2/ngaM/8WJUN3Lf9+KJBWk/Jd2qefdJ96z3jR0j4OgLZ4fojSpjSod1QUzE
o0E0prhpTtk0G75Pd/zX5FKHL92B55WNFcJNBTmqfYSPlOxg475F8lUAWffUfWzD
Ea5nDTjXMB2jK74TMFgA2IqqoyhLAjeUvSA9SfvK0XNo3PsT3ZOi78kl7nUsQ5Gn
Y3RQskGHlDnyYDP3/4zd+LJvNy420VIuy9PigEOP1fXIK4/QHKgoXUvVROYZs9BU
rdIRhbL9P+2AZY74nXm49YBeXlX0effWCreribok2t+VdU5fM/PDqYYEvXTqTrQC
gmt5t1Lu5d7eLwVrjPkmVPH+jqasf6ZU205UXnteDJtJxYnOJ6aZn1P3pOV1xR4A
5MEFShW7rwrE1DQHjsIiuarBkG35QAJYbZ6nnMbyHFDr+odwlGoDiNzhJfeDY8lK
H2oLtxsV7oKaNiAilhB68mvXQuYt79NG1MRJVvKAqVkJsbAZCZVVNQmUq9tY9bga
nRAs1zfFUAv0VA7e2QcbQOX0CoBTd4oz/Nw9LFp6zE8sKoYM0q+Qp6clTf5HcFgh
80ChkiE/OLxRFNm3kGAjy9UQ69v0JKGIGraMWVS80GKKqu9qos0CI8OHwpZ4vM/H
cFXS09E9Nd6/dkNTeOUrzwKu8+uWI7nJl/HTKxibHLsp00lgTkdTY4iBhnJG4eHI
aXyX0YFPJNp3Tv4hIhwRL7H/LP6VHYYaw0QdjxuU7OVHg5G6HTEEWZkFzMC3IxV0
mWQcu80HB9PQVK6n5zs9S9rKTY24ojV6YYbKQ0Gtq0hyGloJq4CUT42419Vthtey
ivzOah5JMiJdnC4akk/migvCNtLpJnTFtnJpc4CalRDSg8+ogk7/6Ii/kGgrAuaf
xzJ2QAwYIquhSyh4ahfLmx/0GNIkQnnCXGWrQHhLxm3L8KzvMu/CWMRp5+rKyu+W
4YNjzd5g4WWuy3i0jL7zIHe1nyMxq+pKJs/QqxArPKEuVfrUhHFTd3LFOa9GQ2Se
h9yg+Kkph56XOifE3gujZemxaEGPtpxAgzx0mgrs7y7nBs8gzz/Ke+waBSuIAqY9
Uz6l4BxaE1aIr2UUKVrrpLr+9VBRiohd6NMLJaIhXf22L2SHmVWLw66ZM8okxPlu
WGHnZo+ncVrUVvTCkB6sm8+t5f1Egb01a9ts7QADx/2tmLMRR/4womvAKpcubd78
H33OfYUXT+Zs4J3t7WxWBxvT+Jt5HwiWggT3imr45bRz5uB1UCyq+eo0nmDYcCk2
LgXvN6CwaVOyijZxVsPTLdOzX+6nfGZ3BBDuD6TluMwlKMXnIWyodhTLAAISjLyE
z55Js3OE48voAkg82P5Lxm0qj8ciO4NY/oSg9zr9d/C4pseTiUmeLUdInDvFbphG
lSqUCdEDVScD5oMh5DDNSk5PJn2BQbgfiq6rZuOJR6kg+fyVFnPX+BllT7gb2+bw
/esnsA7srn5MIzuix5Aqm0CS/JZvNQWxWw4Vm2DwPlC73J3kz+srAbBHgOQRyhTC
zi8L1apjVN/TV9j63RSii2ghJ2tfToTxGXdzIJbEdyOAjTr6WsXKGFidAyacwWPI
ozxlKMP7X/PViV64J5skm9ZMOX4hKa2bz26qP9OypQUuhEL1S/42Ve8IqDBeEk3q
FpGVpimb1o40ciIjXvhg6b80ptHBey8mmD0KW0sXm5q1pLNr/SGpQnHu2IVqN35T
WBE9ZZIqvYt+pBmzpkSONWwP6N7/yyPZhmAoR3J03ZFUOI5PMkJO3yFPC0Guzdrz
bWIcHJtowidFRXq0I9GLAVUeIpLJH4aa1aJlIynmD4pJz9uEFgBtXCZjKoFoN/V4
x7BqN/Z8ieCMQPS7uJEzB+7GYQR027JJSHGGJtcjzo7slhLgPJiiXn5KU92/riZ1
+UtrTi0NbV3TXusJavbrTvlHAINxW2a8UyBLfnkx5VqhcXXKMxv/0+JRAzXHiOCE
CDvvL5vbcKFTArR1VtYMv1m17mXaFLO6fu1YMLXNDFc+T1xU2FyMy5C7RTIoGXUX
mpHuAMvpp/TN/Gj2Enap/VSwKFzzCLN1JaiecZoPfSaeDUyXWmarn+z8hBWruP90
fVxg5pEaIwiHesjLuhFPDZgX+cP3d6aLcCSxVotJM6YquXFx+oIT+ARVBaFMch6e
9VdOQVQDqLcWUXmoMoV074iHiYGdLk9J4liqb+ULdOJtYip1AT1onl34UOCQuQRQ
D+3V+sV/ufAFux1L6vzTgc+hs1pphFncu5NEYcFhs1+fdKOKk2kxpiDeAk/iH+Iw
P97od2ecV4F2CSUjkQGC43zbFxHlqn0qkB0of0phoUtPTI0wFyZfcHUTESFHWUqD
2Y5CvscOj7bOEEMeqvwb9AgRvbv6i717x7+kikRwzmi4/610XzSFSEhcqFsmq6VJ
Ouiw+lkU7Du6zrQ7UboLge8NcKHppKj96BMiPDx4gH0t93oNEJaT7P+xhNywipPt
0LtdaGzl2HX2wSBTqygfFHZKVHUKSi+X9rn6ES4XJeBZvoT/r73UHT5ot107eujx
Ipu31tGv1eWTD9eRYqCqol3XAV2aA8Sa/Um4gX86iUTM/UVsTkCGX3N+5LmVQna4
3m5cRvwf5I5jntYfeowNZEewdRbK2d0bYD3ju8S464KYmiltkN7bMYrgtarUx7Q0
LlVycwLDJ2PhB0eNDFkrtRErIoAWDj6uu8pzWmYwIlFPQw1vAYMaDHjfIUlAzrWC
Sh30k53Qlg+Ngxt1wksisfhAjBlkqc52koVod7PQPsgc3av66EmtYkGQQsSnPtaJ
L8ddbGpB4wIE31pkN05iInHUFty40E9Zl349lS5XHdto7/00JaVnONFaPh0yC+AH
4j1tBWHQJGJ3SDU8+qOO+ZrIJHkbsCsHuoPD1h9o+HkItA+GObESNw/7fcJOZ0Yg
bqT6mtOIKmwRevk9IgITw/KkBwMQV3Av0S9XirWzDlHYVV8FxxjS8V05mlPsKOiO
LrFXfEwkDG16RPLQurZTqd8hMLuPRe6TkcvFmsFvoHozs13M9o4BxrXtF3HBHaGe
QhW83INQR8n0XvdJIQdVvDtQOrEfb7bL8iAqbj8cmcqHEa61T0in2nConVCLTyXd
Qi37619rAA9uY/u5RTMO6KgY8SiFaDcOKua457WMANE1aRPtgx0L2nCz4e6eSmLu
/AEfeIsHSqg4GFQ1A+ghN9eNcUY2NrOC8LwyDxDhhrh5a2U3CdyF2Byvi8efZDmq
dPx4/fgawoTjp1n/bnkTRbPd2fTgnCU+E0VmqAw+bAdx/UuFbkzsnwcMxQtwp7PB
gjYjKh4Jzul6/ZXCXdggOddIgwFlO9L8nwLdRs1ZLNsIKSYPH9qsIYw+EP1oU1cW
DFTCJ/B/kQWKsOqVUhojrTYlUUyEWVhhm8mpGKKj5lSOflys7duRoC3oZpHQwW5O
Z51OBYSGqyx5dHUcDa4e1NE21OTn6a+hcbAt6IPaki7wegOIq3P3gq8jDLGVsgcQ
XYAbipAs5mRzcu6VT53rlamZtq4goyDUmFhAOSwmwp5E5tqqCDtgckCGG/hxzUjD
tq9mQ02HZ/B1qxlQejQ+YwKK07P48gz4O4ENzt/3L+DL7Q+MMIUmKkt/qkE+q5rg
8OCZy99cpqwkao0lfKmZ8ibkYLY2oaC+lVSeP18kDAvBPhYHrDK0LskFE/K/NrZ2
PXYOlVVIs4fDgUxyd0QhLpYoFaoXrlh0dtq+GBvQpmfVbidzE79VdMHFdhpGebxO
fNdAL1N9wnmQ1I2O8D+bNk/SB6NzOkkr0jTIQ+/0SYVRhB5wDtry1vuvLTPfyDGI
Ws2p0iq2E+IcPGB+1d2T/5p29YnQn93O2z9Bm15wWp71C9GuSiQBgXkAFioGV2qL
qJNq2ye28I/bh1ssGPeNPSJChc3EimblD7XLLUqbA/yBA5TfJnZK4MYeqhK3AgJm
HczIxHWLpbg279n9PFftyzOpAX7EffLpZrT4RUa24kO9kBlLYXjJD+WSfeIjWNE2
6m7VwS1zuL27JrsrTmDASybmn2Xa7YYWJh/3wR3vJW3ixHLi2tB7OkD7L215JK3R
1xLp9WHLAup1V4ZuKxIWhWNci2gPBFcUtaPG7zRqcnfe93H9xjxvjp5CZBqlzV5i
GnrHmlANCk9UxsnWP0c1QsV2GeSDno4jy6Id2RO8mvbmg6mbKS36O62yk0tBJkqr
UkWvjka08i+PgjvrVND5wCKrvqx1A2WF6l/MzXfg2WlxavDewaljA4k0Uhk5ru51
jCPGRkt2OyiIhaOQ9Ii8dekwJECTxki4hUvM3MF0D2la0shqEs8vKY66/DT7eg6U
QwuLs5wrELZnpiEN3FVjrXPYTEKKH7BmzVWJ/3qxg3m19L30yvZJ60q0I0RBNfE6
UjYnEme7fvcyAYAJpLkRO0RwprsmyItKzgA6y0juCOXDRKzJpX62ASF3Uwza+Lol
Fwd0m/0CiSKGEYRg7UUqb1zKJsiw6RqxnEdR86RGyl2IVVOuv0w3nPiEvGl2Wa/t
5Exi7cMs/OSdsCpw5mkWtDDuu3waUjtU1xpAkwWm2eMBmEx4fEz2NijXVhakDTjS
z21lUgr48gZL/2A0kKy9tfgZLjAd3YFqhlHGH9N1m/6Dz3StNBCPkPyOt2evnt2a
WWjqyaNUMQndPV/iRro9oajmHCDOE8MzXZ29y/3YNPGx7A6k7GI7m24bkv6SxMxF
TXr/4zb1DkjcppoBTQwFqVjKUNhKKOyeDsMX1DgNQPNgTtrcS47JtPIG++O0Gk8P
enLmwiSV8CgX/pX5n1snT9vC75HLmL3EEE9rX7exFcvyszTzBqvBu8GlJ3ul3dAM
CESlkeTt6650AXfkgoH35e0Xq5csftf+yfna5aIc2WX2fvkhhJ2joMWTuYit1uQ9
vcGRGw0W5mQfQf0zMOFJrwZ+qgrHS1LqEYttvPCM1Ho34nESLCrfXpGwkQ7IlqZI
isHxKTdqfBWYaDG+g01LvtqBgSyAsGvYDqDJKz6s94PI8kRKKmi6FguiSNnTCxhz
q5BVEDnQiaXjYio5QYcEs9gFjjh/Qml+WAnIZ1Z3ev8qvrsmJxSGR3DzNd0bAHJw
kvW4Qsb9K+3p462zJOn0+VHHcZBc8m2Fjzu89W7+SqtF/1N37Oge3Pa1TWvLqgvL
OCchEg4CcC3s3Kt/AA3yB4bm2iyW+SZE/9NAhXF2E6U8CNCrjm5iqIirS2Sbf1TP
R4AOUye6DMKnx9Rop/HE+x5Sb9chocDp19rEdzRMYWgOjOhu7yLkNZ32CsQLQRQJ
DKFpUVMquvMCOmlEeiFn8pqwmceosJ+2VSqvOrGQymagIeVrE7c8PIMwKVm8tnY6
ySW4fr06wA6keZB4LjwyO/WHrH6UVBHitQATXN7VwAjE+fjKATsuIkAd0C4sQpHL
HW2UqAf4MhOFp44ESzbQ92qmcyRfrh8Hy6FBkEWipooSmI9MeF61ovZ3CEayT+SX
iLDtHjz2vjB4m1kID+csXvdKB1eDvC3x/c8wYjWkDggCEDZ7P6G9dnvWle2A3rOR
sPdzccLJXpkZfMbi9xAQrf6vEp00AkWp1yE8p1brR69iwYTcKR2/7JWblgOieRwS
eJLrEbkah97clXqlWKHfyyh4dKWM/5ODDIQ+gqpEAGYPHGvcqw/9HMZbObxSU1gj
6PsD1dsAJ/JlmoN9Wq3IBpZHxUzOaXhxSZdRxb2TOjkQ18SW0/U6Q2j/maRnEfev
s8XLMWec/NTN0Vtvjq0+uwn5FvdSxIOVEVVkGEtS2dyspe/M+IBaZwHQq1EtIir9
IFrovTpkHOT/bEdEcn9R5iTa0Freqh3RF4Dvf72+VX+gldYbx/KP0V4ayOjEnMhJ
9wnzZpsa0TuFoqCVJEOTYo35Eh7RgGii8W+Lf0Ppkk2y33dqP+SOkvd8AN8tggEj
c3p5EnXMx8Y84Y8adW88PF5unyVGMCvcZHQcdFEDXmSiM6crrWKkhCJNxyFv6T2R
YdndPIOCRKoq9B+REhRslamqDkbBKeHca3Nye7cVEtRtktwz1DQpHoFUEVjRvduJ
g9iBiSa5Fyu2YOZ6CXYclQeH0B4Rbj0SRHfFhDEP8Tsd4RFPLCPF7Fji+XVFiIY9
+X+YnMlBFWFpmIyj9P4LSEj5Rgs9Qpd/Lneyl/XovQQqqBq6hqJVC0O+FmuoNxZG
hhaJF/HM3cmjvzHlpthrZxOFg5PBEIByrHnN0BUprdyU47DIscqLU6DstC6wYzMh
L479g1Y+pyERbyb5gePHraL9xSWRO8JULnrZWto4ckuD8QjfNZpgHusc8Zkdr7O7
xBXZgrXELW4YqA0ECCKPTKc/gP14FZaFQER0rud2UhhFDGkP1oTp67dj8Ifz0eYa
7Olq253wgn7uvRklLJWnMlVNqgwU6JZv0jiVB2gmOX4UKCCfoOUbVybJYd3sz/9S
B0h8wcQkOybZ8GEeHDD35+W6cuZqzyiFxpeyzOGCrcxu0/xOJgW3cR3V4nW9xOjA
uZ3diaDlRYYt5wNZ0AK2ZdE30berK05j1kxUwiMg6GpO2S4Sx4R7w/QH0Y4il1HE
tzCOEtB/f39X9h2mZWXfBJh/qZgUQOLXOpFIz6GSvQ2KX1n/kwKSbUPQBR2QBHfx
8YCm8QpCh6dhAmR617B3tEFsfR06HqSdnkKV8VX3JhxU/8yUpt8WVnWDapvvIKaL
EckA4MjgFe9EUuOdoyd2AKL0FAL/4rAsFBq2oIcW6nkaWbmm/pBf7TnzSjQciwMp
oJK2hncbS17z10emaPFzvP/i1NM74nxsWAsVr0MSLgsetari/QV27Z7boLmyEdCm
jukcnfryyXxghJDAdN+UKFKw40dLNrzJsqsOV0ysocp4CcAL27BVjMUUIY1ojous
YexigR52eR8ol5lBlTB4DSMU8MgTRuM3sqG6aD9FbLpNrR89e/ltZvulvH0K1wgp
pXeuOfl++hJL4f5+nU0oniv6lOdL3U/q1JcEjKZAa2z3JoOsFhx/5fWud9Dy2UJb
UB83c7AiB8aov3SIVsa0bMRpAHhHrUnMkkyvARscFgYxOsvd5cRul9KMGQLSDERn
scBFgIPyu1JmFNOrciLzFbbF7wEZIEFPGQRtnGRqrBKL0EO9q8cl2IlDT0I3uT/P
vf0g6FAoj4YxJySK0vbyS0DtVWQHW504XFlhm/v45iMlh4QQB7fFe59EPYemUMPd
fHhCC+PVOwPc9U5egcc8PFbHvAeEQLPvIPlfDmvxVRopsfuGE8XUpM/WqWIUyLkq
T25q9mOnV6q677NgbWPZ8xanyWuXwyBA0hQh3YakalPHJ8huaLRBoD8eViFGHc1B
1wpccz5Ub2kuydEQd9k2FrA2WNbeDacrJjSu8Ue9Mcyl69LKGLOhD6Z3prH4G72B
AU11CnqFcn4L2WLTv5LjCqmPaB49azYWwa6qeDeO70ddN4wU/Xjr1YNsin1osmtG
TDlDFdDJvXiKkSG3kQFUFm6sdp6IDAhYpp41aooit0Igc7FcKHaAap+nWOReB3Cw
Dktb1XCaa+F/Vov3t4CPYzznSS0F70b+JgmWK64osqpERbrAzsZpXtK9ME4E5GQH
Ny47V3bPZGoxREmtyVBzjbGd3sMVzqeH3nUW5PkoyMd95dNp+O+vAm9JAnFlllqp
rQ8XAZeuyPBVlosoyz/a/y0lOUIdsbzrrEdTs7wSBdKr8/MdONvjPuecEmJB+Stq
na+S7qoGeB+YsM3qCqoE4DaO6kRw4KzBzW6ZHs+gKuISvQ8DgxtbsNq7KYjVDkoQ
tjiz8XtPMuiyHmjDgEJOfJ2RuJhud7JwnE6bWmhD2h2pAtxD61GqAXM1EZ8m5/zC
p7awd8oyu1HyYmxsEHqF7YP7kpjdWJImB5DdHcAFS2GpplZrBJI9fC6/Ah1t39Fn
3UdmmLHavawDEo5eK/uLENc9Ic185kt3mtPhmbUCB1ba5CFn15brSYpo2bNkjqIr
bTLGrVMtxR5YRCyzBgShSmbxYU1u0RQ6tkxHdMDIOEecQkP9POPZYG7J7IvbmHm9
BYvENlCGOfECtaw0KQ2kF3LRrxUNUWLoHayra0XbRyM8DfRyzYu4RqLLOcasip5d
VqinQVBRNq9Am7gAqlRLf6QIaVbqMEGAaCCYW/379kaizN6altEWVtRuhb2yyet0
H4ZTiF0N53aALSQ3FmomGZFQQ7HUgBJdoldIjxq6npne2FbYzknUJQsGcul3yY0K
4NWmEOSPJMHIl7UVSOAmAr27j58fPOXib9dJulBPBfa2n96fjgaVPvvv/h6TRLyN
cvptWVwzL3SstVL2/vyrEbvS11j7YOp3vHDDK4VzDnIbj3iVlepacv16CBPmzzlg
pyyHy4K9v+vEAVzkBWrRBWF5KoYNz68IXadjU3vq+sPZA3o6Q4asRSphTemr0x16
wuxKAYcPSyDXMq43Cj2xxOl4qazFBZxkYvoUrBel+PD7/Dshi6IizYCDkInEc4sV
yx0QsQSv2ubg9SfDPeereMuiPSxJZJAeBlSpLGrOa/RB0ZLfNml+qwuGemAKhP1n
JvVO94kWJpITivwps74ANtNkWSxL+Bltqe+20zUxyVeXFUNdxHEubYZSF4rscD5E
jDZA7Crcj7tjQCMUWsrUpF6YsQ32JKxiUl9UzB2VVwRsEGfDr6N0q/921UKWTnNA
w2V849+2gUbqBF2guK4DV2FFzs1tHrr2ksLq1g75msWpyCPbFv0gXDHq/PfG+Q31
O25rgSWq+XNGYAA6WEOuT3Pvs5vba6kqMOYKkVTXW68g9YxGATQMCMU6WYaGwkFo
rHFWbp40hvFhPXlwyzbhVZ11yzMeZjB60BYMLfl7gdZqJvYKsYab+y6d5te+db30
+Yt3rLSWOQVw0jvAhFl+ZRaQuPdZxk1Mo0/HiR+RKu2pEDzqu36ITIkzPFVnwYZW
N5Ehl8/ZMpJQ+HccY2hrt5FqZuvy7QfBKlBW8AN5J6aFLyS/uFGP/fNSiI7/HDTR
/VAJPPxPG2liFJ9Ny+sGsrXR+yisXjiscrbjywjiNvyy84yS6fNiB+bqjL/CeKDM
xqicbvNiqoh4u4ICNR8mc2YHABBJX0QWURy6IcKQBB1+KSmzYnVEOTekEFJHV0eB
x6a2K7yuXREqz6SJp/VetwT8a//XaONuoJkqPRniWhe9pKCQOXmtkcL1q1JkLLLA
YSDao/o5yQOT7J3fAyfro1x9081Z7S3N/QTSF311qcIqCBH5M3WTFg/ze/tEUKjQ
hCha1s/ZxOQNO21qBw2n+MhNzYUQ7rBH4lmLUBWmITuKnnxbRn7TXhMBN42QKGid
BJv/1sy11QYE6gHx+EFGEeS8YJx4tMTCf2oUZ3gM44Qz2sgxuu3NbrquFD++Ro5I
QTHTeHOcCBcVjA/aPRQZkNZaSSAxu6Q1UtATEL4ZhBLk+XAOoKj7lN+5tpOZ/WL1
EW79Cdtt6vBT66hDTokTU8Qoy48X0ykHu9I7OYSL6w754Ypwr92BT5j94UjL3xhv
sexY6lVDybnzEZOxpoH9JOUHJIHIdXl0hpTCk9jcjElhhCFgqG9tK+H1rlCU5uTz
fdgqSKKvjyWDcZM7n99jrjwG6rkhJKF/SKUXt0/PhjKVzdq4gcfIMbk8XoPHnrWK
FWBGK+KmEeOswMRlncvLpkQcmGBzWlglTQxt10g7efME71EIEj4kuMhLsdcdc2Qr
K0lkO8BjcXkRg1auWfjpqJQhFwxviztpx/QQcrE/ONHmz29UFtaiaehr98LzBino
HFn8Y927LguFB/UvDs7Wksh2jX27/cbgiMk60TRIkAgM1B0qVf97c9K2zr3dX6PA
ofad6MF3pUyiuB9PviNgmgPILDyC+kGuSFEanSiREKuBEylyitKbpOiIY5t9umyP
pFrbxr1534x5ZwjOmJwxeNgFIMJ8/Os7Tg6VAmKaNCTaBXnMUDaJW4b9qnCr0e5N
/hOafEuGdEODW8whyoewxuCznkHskqjR0CP4QQjOi/sap01hPh794q1YfGEL1/BR
I33GLhq19OS04geBBhuaygsNBh7reQB2D3Xrh6bFb7gJdroT8zt4+IN/c4ibBArU
tp69YkS9wqwucCxi3gVk+QeEJB9veynlnYQSxt5ezl1iOHLg6Ha3+yIF+XW//0G5
mbdABaqDfarmQ9diNzcUYlg0JOStFxGQxSqaEBuqAFJJuJ7v6RG0+eMVjyVoPAw/
xYKPNck+VBCMLEPM/NFHxn58gWPWbMcXxw3DhwlhZGcMGYVWDjgg4KdH7viXxy7Y
A7CS0n7eqn48DBT7kyjc/YHm8/nwR0dzcvS3/0AQ4yLWYrf9BV0ecDPzonTPGt3r
O6b1PsbC4lhAbf/HyRVOIA32pCOGEI44nHdk3gT+TYabiq/dhw9fNK0/NoZ3Nf8Z
gXikYw75iZdVUefRCfjyTpOdJ3sIBcZwmSXfZRDzQEjQgwdWK1+cEgZk38WYIuW4
NNi4iiMbcW/s+RBGf9IYcxK5DWeRqKW810ZX1tPgTIK5OtzASGYRKvlIaxo/cV3e
lHpMv8fEw/XnCvq7CPgzhkFKRtuWVNkL7ihGk1M9S/86l/hqv/T4JZYhG9FnkLIA
30cTQTsn0sVCoAvs3RiP1+bvyZXU+s21I2VAvo2w9ORuw+cbJ9UsAh+XrwJ5dQOS
er5SU7Cr6Rd/L7ZRZQVrI+g/PNVAFPJLKCVeTY0itMCkYwKThpVMC/DZvHw+xtrv
0AlfK41m+bwxvwPLevIetD+wEG7gtGmII9VeBeV0HV6mTSD25559FA5vsbDX8pYA
p1KDIR8dDMe17Apma67NUgUZzBOv4HmCgivbVImOm9DoNFxC/I01EVGeyacMXykW
Hv3Vva7AiBLg+cjezjvcf10+gf/pbWDJN/I375Mqy76IlSjmSf/liXvIyBTgtCQZ
3pH2MaLMrFgEaE5C7HedwFIAs9q+gItTx1R33hwz6bAjZZ+24a9GNAX2pnk4ektA
5WWgFY9VlCTUf3L8JffLXU4KlvJ8fTZnL+1qmLYdVOzwITdEaTbMEXlz6n6NX0EO
xT3b+/0ISW3f9QxYgHeiZo20Zy+svl7S9r9HQTPO2iuJQo+lyU/k4Njm1GOaPloE
ulPz6hUb+ECSD4Igt7UwrZW5hv218/mZC+wGlZEGpD8bSxMcWsDIkqwZftZulYG0
WsWYxeR7Vpw/qSo6cKLQJY1QToftxIbMMULW7Hsy4JLMNk8roWfzI0t+77UfKoUj
Ik76NSziuxqOXjRQDVRaPn6OSgd9jl1j+mmL3uIuY51PqGrkrHyDySqvHRK/9fQQ
csVIwXHr6qjEfBja69cHIfLUzrjyWwHxxsj+IGC+PUA2IT3leu/25gZPD7wj/ImJ
Hf3JQJ++xhW97pINBH/Ffm3whgS2nKFN6Ch+bHA2KsgtAXVaAOTnYYKBxeQlLydh
fxU5gBlrkh9yknenhanJ3JZgGQlApJbWKGcjyP3vR3FKkiXdjljliScnM/yvpW0s
TNzIpBoE2RkiK+wIOQlZhpy609GiiW1U1sWh9iiXRZpn5ZlO/joofcgy0tNly5Bp
haAhWdu40rJG2c9WvfcqLSNC8k0sG9CGw3/8Duq7rt0SdYEjcabsQwnLZSY1p1Ev
YgyThPTKO1/6cAiGv3j1agM8zoX7o8nyKrnaXfsn/iveJfbZ71jlm97ai/3qp0SB
X28XY5rt61YCVlAanJLjc4zWQWyUu/4ehwvTOAQ5YpvKH3l5LY4JxvO+UpoB4DmA
tTdecQwOnxyew4PSmR0LY+VtDBGib97/FI9QajpuDz0vEx/HRSs/bTxkfsXPOV2q
AJTanigEZiijsKT4I6cz7z+jj012jh5YhipUIea7WoXsQfdo4/OuDCWvg70liTkp
XrN8/2Zn7x6iMbwkQN2OCGFluAms6oKEVOKth5lNhhUbqAgEcPeMNNnXR8x8e6Ah
cYkhwOb4PWmO1rsT1ahPpAoPVzAgr2vgmRieSAV6nwx7qRauYJGVfrmyzau1Zxct
jDKNH6z1hUnHN5O+NeOHgeldFrJT3ExrNnqPSoE62iKYlxbylc4m5m0o7jhN0wDU
QDVFzQqB3GduH6l4cGDDRj36LVMqD9pnesRSZTUxyGbWiT+nHeX3zLVHerrn2/ZH
T69ndwRTrvLy+q9Aw92Wswdl1h6DjISflcB7UoxJdMs6wmVCifpQpBKruC10hE0a
Jd9larjbvUnvKQ3h7rrEBUDB88FzrEOJq+RXCvryoRJlwLE3g+I25btYnAMDq9s2
4YUHwoLSasfBcmiUsjYyHM3fq8wxi50bbo4S1uVVUuLikIQRFQPLeJ2Ug7aPZLKr
OrjOorA4RLzNUsLUMjnl4nz6VBcQjKJf4Q9KabC1us1TsbdcDTOWS3ralGLrf25K
0sxxJFDTdgBpRbdBCWJ5CKFfZHvxxbavmeOfrHrS5mB0UTKLLC+QG36z4smS4WKx
Ki6nqKjcGl9gsk/7sFbgQL+mVgZ9PWPu5oC7t3T7+paK6ZfTUiOTjaMMxhbqUY/h
xT3JzEswie2MAo6ixYFVBpVW5AqM7E/gdLa6lWLz71u3lPAr+Y5oTlTgqeC///S9
ulsh2ckj68bC3afw/k9Z9nNG7wWzV1lv18Lgo+LrglZNLgmjCtYqwWr7UIFvR5jp
gkG6eZLx0e6JC/ofPBlkoJFZFIOpP7lpaSlNSE85rHqxpgPdRlins5aRgkcjeTxz
qRnfQgUixooJZ/SOEXyhe46RW1SLNAIbjk2vFN1+POYeqcefU780XHvVF4NK7tfi
qW91ceoryBto0wILgLGSagWT8f3JWpdrVwZlgTCSKRTuHtNpotUhJ3AbfZfO/aYD
oDowouCFtbGV41Q1l7tPa3LLpoqc/zKlzfR8qG23JULif040MRWTmRibQVufpLGv
94YvwZ7qSq8nU+4X/roXa5h+oqAd036rCQ1kbTV4/M5tsBgGVNcs0AARvAc8gebp
ItLKvA66oRaVPDXsVzB3lCaQiltQYKD6F49eXnavmF7x8/ujapMvzl1jRffWqTzt
wee9NEA37abl5tXXFixikjJ9E2hltoX0WGV1WbqmFKkK6j+nYXvMQd1GuUI7j2o7
Gg6BLEmkb1LpIPq4mPFo73A8ALz2a6cKXM8wnNqT6eXdB5S6BCe9ayGir2juXpa3
r6I5vFaih2j+Ftad6wvcJNz+vofOTMOCgLiKxFTHNUN5YdSpuVG1vaioMDMXbQU8
jQIek7GIDtGDlm2ZhKXS+20d7Vm1HGElRMnN73P73ZFsCxaWchUkl2WYQO4UC+NA
au+ezVZGey3LPwW1FaUCWlzmT57ZWIiuOvkGBFjM91JaJVrzTEq5logzOPG8s13t
wlNdItHg/4rHWckWSHVkw2BoBCl/sP/2HfKBn8a17PPbAh+R1GObvzxv4rlilDDi
EyqIoN5Zg7Jj/bCIL3mTOLA8e0m2R0GjwZYj21q0Co/qcdmZ9h4wkN4++u/tqHHk
z8d17eUW9CkaNlZuenr6DsB6F0AOoFTEaQh8Bxe+ZtQqME2KAO+Fot5Bg5EAds8p
Tky/E21jFQO6txiXKFgx72MHFKCqfoEMJB2XKP256vj37I2e6WvtRAZ0iCPnXzkE
abW70i+ShLilQ3b6eOBsJfwQjZ0LwjB2V9WXxEIxaOvY5lkS0QY5CH0OztLctnbO
Lu0JKMJf2q/bYTGoxC+SXWL8A9rwSh4G35pIiCFWpplE2A/8/+f74kp1UsAh0Tqh
DDzYv4CssZ8gwUSj+7WkZbWH9Ot2gcxgNgf6hQ0WGQEgz0upDUhfifN2iKD5h+Aj
ec7hoOFUzs8J7ZafYnwQzGoZUGY54uPdY3i9IE/96NCbk4IJHODFAtjLKxzJFT3h
r9z88PIGh6cHXP5XE56XdGzEtzTSodorFkIboFB9GRXZWyqpCVjzGMvIGBsJQJFr
Tvnw/6/eBLXXByTCY/zHiVTgDMh4Xcrn+X41cvSAzmccmp20+J8IYNZZIkTzu97q
N2vsWYaDc+zRFQTdf1wsLwrfQJpbgQaFWIG5a7w5btV5IT3rjv+VzIkSvyVCARTa
nCMnJs607og2H+f69mOBlZ7ZhdTijShuWOkZ5YiaETyMduyEaKVdRqKYyCOoLcee
wdJjCHW3QIId8ZGZRGTadDbPBItMfXAYI+3vY603d5MNxbRNhrBH42eV/zkTnO1u
zpUBIFKstEbzSHrZ7KGcpJ4pqUsm/gaIBem8Ut19oM3IlOCKZ572B15jQfE7v6Y9
3tFqInxpI1ZKz6rURBq5r+xcHlr7gzv++zxmMLeXAQgoQul6UWgRbQkP31RulrBU
Wkqc2rW1oAQfyafcB6YyCIAh5MlKTpPhNe1ZEd2x2vORLuFscfF2Ac6qNzw87iWj
85iQpBz0yaVTRg5cCJDiCma9o8c7R9HuD6a8A5tPj0ugqgptMCCHpyJGnG/3RIB6
GdecS4+IXzzpCzG8KpE0EhT75TPlKmq2bR+mfUWJOpHSBeCCVcrXFUU91xAiIILd
YxxiApCXUHGrNDClBn8DYccyl6r5SCjMjrnA1FGs7VFOBS6oFAt9VXJZ18gWJbX6
7cREBEKZaJwhr82+FX7E/+5F4Qw67Kw02w2F/VAmgmPTHUyY9SIRmJnts7NtmiMS
G141Lk7POBu6hZxQAJukvpEGVyjP46dub3CJIjJ+3c6rzwJudGnSaxRyLVHd99Bd
m+m/QZw3QQW257pW3IA+C9W3cbrUFozqXKhW0bRA8wybzB0JrTfMfJbO/wyA+Mft
7GjwWPkC3LFwIg3e1BBMTep5U450iVNtNybQZhCOtCAjnoMDF1lWkMSmc3AKH/yH
7ahspkYVm82b0XQhz61xAQ0w99Cgfb1vxCTViLdc01krmQ4QrIZVrr0JDsXxUoKD
k/BrG9sf0bNyBgQnmUfgEjLD7JrDLWS4ev8L9RD0HPaqmsxcZK+0IuktPhjFfcmO
e177pxaJI29AtbnPknR0YlJ8+js5KSugJtQZZXP11yhZ9MljfhTudBVanCdaY5iu
VD0/ynv6Bh3+OpBlaf2xaTrzyDHdrhrqEaIcumH3Y1qnZDGzbgK/UMtbsSDxrRAu
FORk1Bkq0R/Nv6313JzTawN4H1EqbOSYL5ZEdJSk2W26mz2XQe575xmadSpvv83D
nmfV9vMxtJFGr826Ng6x/bh3yJ+eLou9qavgf/hZhQ1zg2qHpg87rqkQLf/rkhbU
DEuYlHmf++5JZwky2e0IxUSFyZSzO/7i9n1AegxS8tV2uEZGpKja8YAiq9gzxzG+
6jGIJvn7n+DMvsOkN8Qfy8C6chDG6EKy67vw53DSpAuoRzjlmISjk3b1Y5W6U9g9
DHY+xECz9IkqmVU70tTbsO+JcIv/+nPNytbUyKyFPhgq4c9uS8PunoSuyQ15eg/p
WVIsQYgV+xhafmgpNVmHdk81TnvYilmSJQS7kIqv2tJXP8yoNqjGxgN5DgsSUsXI
NFToAh0lqZ44cQHtKOeLGExPnR3Kq6hEngMPsp231I1mTYktfKuX9nKvn9JMrNDl
4ZhWTSTW0zoF9kPPSFzB4EeM+7RUOlzbJeOEbHeJpKe1THGRkYw9xCQ8SQjjdcoP
zFVCEszYNQTH6aMxBaHrDoRB7U1qvkDI8AGDKOPTAALgLUxyqkZBk5H+MFKpauc4
XzcSyUn8VPi5Ds285Rwqf30VTZKDCB/VzZDRtS34rITJ86rHV2y8Gp6DwLJGylE5
b1qhnJ2mf++ERX2bcAhsP4jPpn4GSt3B50xvyJzOrjyduPwcMv8Zg0JKK+MUB24F
PWIX4gNo4nWXV9TwtgkEJVvdgJfcIE6+pf/uXSqELmsBIJx/iZIPKSCkuFepl8Zw
+X6+piSfFRrsxvWAvsgFx9cPdHDfDxXkRp2oKrekAKvfUiArPMIFCXAzgw282MNw
yO3xAMagzXydbGC6cqEr/+qJMfFCYJ2/KBpvYf3dI0wUk0EzIUdRkeHn2PUHBdoB
krA1IGmMDSW88e7oWgQRSZjnw88p8R4xCSbb6WsiPUFyjqsF+6gKVewg0D5klvXE
g2/FTMejLv78/RfAAUgcAbRQ3rzku71M7PCGf0/wCc5tlVjbeTgrgql9EVwQZkv9
QX9k9CMLbuNf1GEr0xPk79GF1esZh3MqcRQbpu6AlDoXoMbiNxa90xGWCX886DWJ
03mk9ZZqFxrFqA4jpacghHISLGnkoEMDVB199KBv5N5LlHYht9VkfLQluUkP2uzc
IDrFlubzPZUCmkoy4jiCugg3D7ibVRUsNDtv1p5dof9AA7JUj9zD7VzNu1eGH+g2
8/gTx1okypGv72/ykXSm6lCqVmPn3VezS56/coP6Ku/D/fyDzhZwCbZ5whQBHItK
/oo4IbVXZWLdTOnXYu5trx3fEnaJ8VcheNTuK98GGVLq658eH1OzAh4MSPXqVUfc
+TqavzjHzfFiHbO8WCX5dsUAAbkA7S3uUPLrJTH9IJMEsS1bZUuIAHHZBHozE9kq
Sk5xL/F3xydTnWuaaKFpvijIUVS/8j1L5Ia3CC8Ma5z1BO94ha45AgzGA7rIskMA
AfrDGW1HuL1/kjWHz1XHPdVnOv8aRBb0jqrJeigPt/Zn27J2GBcXgGusU1ggAi6H
GpGDM2jIdHfCmL3ORq2nl5C2yHiyQPbWsFV2xPduQGbB38u1Q8j82E2VfXkop2rA
4e2Yyc4qTYKIetGwBbU37JTSggQ+4W1bVcHA9aI2Kvfs83MjGsoOZuGSGEM7fDxi
uxCn8H2vQXZlRQNc4Z/p9NnuA8Zv0ghP5JhCni0qYXe0mYfxTwnWAHyfZlKhuWqF
wR/9Dhk9eXDyYZKxrdJk4evXndv83a2f45KxcPWAIxcOsF9jhG/3mf3WUkdj0ugO
EYUNHIgoHRxD2WZ9NsFagrrMB0Yz4Ro6Iqn5+M78luqRILfAky8+FAksE296mNEh
MUMxh1rKaNEEUwk8g5+79qsJW8FaH4Qni2aJLxNGgJxQrmaoK+LiTDTSvdmFOU4W
1Shd2FHaoqMZJ1uqQn0nMpgGL8ydqWN6eqqPMWkOP+tMvCnkB//2KCtPa65NluKb
C/PtTzc9akQKdRXRk1ZA2HlzTO5mENHCZMcsPgGpT11eEV67Iu71TuXME//b9pGa
PCoo3ekVVIu5jxIONi9HG+RC+UzRXacKyCJ3dgRnFffP8v4M7gaVVFV8b7TETbOw
WL/w7jSI25zyxZjyO+y6ZXwRmbad4txWAHaUVSj+nTXm/CTeI8JOQXH9k4GaB/SF
mpkMsjz4zr/Bod8dfZkrw3ENOgRxwGgJ1Zddtfed6L8QL6IemrsWEvDjgZbi5IYS
7gHaDuwubx0rqmImpHJsAvnHK1HVQ2uRAjCxX0FVMa7CXPWBWBGQe01YEga2vhNu
Ya+XtjVZFWw+kMFmWhSYwUW5H6YaM6DyP9NX6hAwH+lCuNKXSPPLxTuU4rY5HMEu
tHZWMGtNaPN5bv5hFyt9YFtF5wBKApQoUGv+jmHYUXMwvNm3hQVQyK05GgQUe5n7
cvxuTfeZmyryCjvmCqgAzBqO5W2LD7mwlYf2TLCziBc6BFX/brR4zzA7f6+jiUyC
n9ly97kZefujjeoEmMB/qcFWBLXxdFudhv7gTSTjDoMcz/NyiR+IsVscEMIlJRMa
9kxdvleC6CnEv3EvnE8uZ3981rMmpLjDLrqzaNf3lP2nED9SfYfVy6lroQk5qV/G
x+rIH/NgIHpNuyLEZy01T388SDL5xr4q56eq7jAQSYMzzACwDzxP3YFPc8czKUyv
hMrVpaJcLIN+SBHBqziiti0EKJTTHWOpu1m4Y9QHei4P32/1RE/bGj0/+MzyASZJ
4WvzuOOlRD3s3iokY/eyrP9hXX63c2X4A1qr5skpSXYTJ1OsgnFTRb6oVHyVakEv
h/9MIpLe+YnqICCzCrge1bMvzVk4o/YB03Uap5JZfxYhQz03ieV52mFpR/aNBKjV
Ii7oGCrE5ZAIFrf+mgy1DJmvBqAIm54+Xho2HJTLBcHPAe3LY7ymayE4jO6GePb9
Udlok93fXDBfwvtH3vRH0V89LXZAFLAhbefSTpuSxYGOYO1Z+ejWA90auqNNzrf8
iWYIS29i4/iMuIiLU2pOJdjjpmoM65Y8YABJhs1b4CA6lSJ0ijjjV4uR6jbTO5f0
U/n8LSrx8JAgF7mgorHXOgNjbPOhoEhsl9tx5fJ0XF58uW7ImIuBB7DseWOKT2qk
oQDIZou5Wu2DCtgWTCFQ0H4mlqbdDIN+EIqTT39ldaZcLOU0/C/Fu/3Ws24g/rnt
CUEsDiViDKhiYdFZyaughK2iynh4/+SwD6RtAtu6LYwlpp7hUnSwUfhq6TU7iicU
kYO9rHng2iQVqpKfA6V/NOmhW+LNWeW4/+Qo3H0J00GHJ3iNaLFi0XIdML2EOAco
OTpeDf6PZoY8QP1silBcGLoJ2k37x9g+JdSlmvDRPGKdzZn+h04FApS7MPH1Ak5Z
5ibkRkuH7YJ3zVENX6xuw1Yd1Ervtz6HpNRdGkXFYn6CYU+8uT82iUl0UwkJ8k0z
x7VJxk1qyT7xIKr6Aqt1fW2NAfXAAR7CirRy7ERHlmJZgOQBzlmufnR8bL2LZprT
JiPSvScTopmfgANoW6n1oWFWGx7FDlEPaIhXzFj6Zkq47iqsa+DRBaWVGBidRmC9
4AgqmMCP5w+JS9nyEkwGVv+vtVuFzDFSuuNwHVxOAB+yEAnpsHZGiG58B1pvs8HD
NDkqczQad7WnvbrwyjdIWfjhF0ShklLYMCVBIp523MNPAWwCgV/l9JpzQrzFLTAp
EXWAZ01qYLwHfrWur4bOG05e+IxICoVHfnqXheN0OOWDwCqDKmrWsBFTOubWkXcU
rjTj4janWw4B06osTE4tJD2wsOvlxc0ywl77utOmSRzMd1PBql1rP8QUn8sN5Wam
EbKbJEHQxVs5VGZhAVN5glbP6z3vhfYte/5WwBMpeljpif1dRV2pqaKwWpeWpRnp
xbByVgZGfipA1BnRmY7iH+YYzZzGSh8xx/cp7SYkqzmgI4GB9oH1EgdB7kpHXyeh
Qq2dKeYQ7yzxnQj2QflP7H8UHpnHUfAmKdSRsSQRQ0q1v2ANzVsTp+M5yh2+J+Ee
8Aed63YQfl84daA4Pkh+LNaLvAafy+I2Rlw9I4+DVQW2bR4FyeZsliDkMsyCeCF9
CCBKw+dnKiajv2MgyuK85onjR/5kXqen15vBqQvk8oGo84no1/vMfXjVDvUmyYVl
a+lulSbPkm58UqYCe7PAI7UodoPISzzYglUi/U1NgEEw7R9O4aF4yTHLiKtrcXoQ
hEwVuLztF0rNDtkpaxmUxfIgGWK9bfGtchG/7n2xVy22st3hsYLd8pMfk88GP6XU
ayn9YERII7VMrpZGY+RbA0rro6erbMTOpa84yl4Q0U4FwaAZp+4cTHzaHvfFvbbf
ClqxOrYpVrOaNKXHUBAt9h/D8Tmi0qbWzkfTfWEclL3wI4qYhEWN0cxM4kZSZc+d
zFmg3OE+LfphQT6xBdOFgRQTh3v5GzT2GoMTnIvFR1vRB/IP/23LYar1DyqCO4M9
sjw3yUYhT4QMtbHJqVbdJ/4bjbY4lm7K5cD1eDoFl0OaONVJjdTNexaJT1Tlz5hu
qIQOmb3yDcyj1BtWLUJo3udwMk49AdsNBira7F9fQlC0J2RbniinOXvnDpFfVlh7
PFsyoPn1AFKcar2mU5M95/QEHfPV452sN0wUVLOmie/fgmtEroQ2P1blIVxkH6AP
ZvoM0cythu+l3lnDlwjLuV9P4tcBZCt8CmL2oqSMrc8XNFAEa3zjEGVMFqBPvqN7
e8BblAvgvZNQkDcFPUVGke0YB+JiHWwuMxSF5iv9cE9Tycbf3Ah/hIgdkCCQobq7
7A3PLtm3Z2FmqVQKWDSJ+WhZTNoyxIR9t4vkd2939oQiymR6fTdVHvYJLANOBBkS
I5fpT3iMZL+RNslHf4L6dRd5POoUvDTzmzgtwt70xS8LC50A8zQjTQtcTLjEjYNj
1KXE9ZBfTbcj/Lyc5xYlQZ+jwf6UK/VXBoKLN8nbnhXWFLuEnlwZw1+QRALe5dBP
nt8o9vyuBUmFfWNPjHNgtR5RLEE/Gp3i98S4Z5tIfTkKehdcaQxI6IFLEXCJbXuz
UCkPFR14491j5/w6Xqtc/UjoviOm1Rv1EZI1FTywwBqlD/lgas22LPWrIqiDXphn
JYcS8sq6E++Km2GLbgbVsgKJHLIr9OSrMiQgpIGrM/LKpuBDGR5o2x4QtqizudqG
mxE/S/yAUtkEKrkc4U8zAXDFy7AblgClYUdxQmyh6hemMxA+gxoe5uwMqEVgGH/K
IOmE75zPJ2k8HF2ILcP5SaPU2F0hV4KuQedZknN8LT64bGygOZQevUrf5GJfhp2k
RjFyFMaOh+ZOtGoaWqOBtI71rSZV1l4Cu1jDPyYU18wuxHVoeRxTAy0in5TqR8B6
ukG+SJIX5L3XEdVkTuKNXUEyyqBTI+SnA35cFlugoYeEnjdlXhkj0tw1klb3QhqU
mGyNVVWHFEJvVVcnqFIwC0/d6U+2mkpfNnwo9GJf3ORK7HuFnNz8gyPoK9ZIYdRA
HWmmJSUnjEZon996Tr2NvcWEzSQm1mqul00qPJ/MKHCHwKiq21qQrObRTRPNEjho
vzMszzfMX8dP9FqqytB+yAalBcDdKHKZ1Ry+nleZ+hzZNxybCPYb2oFjw+PCzD1W
TjRcFzk/DPv04nA/swfQNx5wIsLQZ+pd1Wg57ID4nHydrObT1d3h6D1tyYmCuQHF
D/SNFX16dxM9y47sTdkrMP1ksd5zl4g87d9eez3aortsrCe1vjaBJGrT+KKWbcFW
fIVV0ll7FwaBos5DK6IItPqL56n6ed9HqRq++ypWkCidJp7SJzEc7CTUabEgUT9v
2MZbpsh4yyUH1kc6jAIb60mWVi4cm3k1hcV6WloB8NroaIcAM1bi/Pwk/nIyrETN
dH6PF5O12vBhigys2SrG4lHTdk8uhbjl1yaLruUd+SuTHwU3Z/8lDSordyXdN8Jt
loXDDALIETexj8ALxje/t0ibef1rFPWwpztZt8lQ1OpkieRIGoTso4LJEK52F5a4
+WUjisw1EznAdIkJs6iQSyPILnAKl4v08SH6T+Ola/3YGbGdYXwPoPTfHVIIT58/
OWiaC5BMb3KAG9lhdLKkIhNAZ5/KS1gX8JsOpVa51QzXLMrlvMxpz3DXZE/sfmXG
aYGzcDQemrTztSsNIIu11/6GKNhW8yo6y3i5C6QnvY8Ud5BHrtHBybAZ004dMb36
wPXks1pWzbIj2rDQhM/aGZ+juvOJgqKaxvxF3VgpNT00Kpij/K5D2ppDC+RDHbxe
2wI7UxTJp/PoN3BXgnwboKw98VRHiryhq8mxGKs5GOevVi+NVR7z4C3dwZzYaxkK
kDMSlfmbpfqtSj8xFLuChuF0YvRWq5zOHtofolqRoK75DphY0LAai2jhTiE2gvVU
+sJlqPW5ua3nOe2b92UM6Hw4U1NXj2LD5lcdzmBgPHhHSC6P+S5qVt3N36OZDOzH
iXyda8h9L47ggStiquuTp/7eoa9nyUoQgvcbwLDb+5M9J8jjgE9kB8tgbS2juE/t
yVGcuKodPF9hqI5jxF9Yf0SaT86TZtbe0X1r9rCBtoMsFs9aULbEIaiCiieYBvP7
7vhSUdhKroL0ENhq+kpz4ji7MqK5XBZZJfy3C7jcme/hLF8x+TEkS2fmfL2a6owj
q5AoeL0U8zywYpHEDEv2ALBDJihsNCu+cy52ED1g8Ix3E90LYtik/yo5q0jU9vfi
uQIx1m1mdC4Nuv46ajn0xjYCeVfKK9LJjBQ/uEfVBQHN1YjC4eF1Xfkl1ZeH56rc
WIt82+/qHhmGCtW6MLa11uvqAqgQVEPCo+sAl+OeKJxD88pV0zg+RetT8z67xyEB
SeSWyc/RJHgeSQjhUtZX6EG2trcsB0S2/pKBECuUZ6sAscFPR2iPkGv1dP0iKsSK
ggqydKJrh1JELsDgFTgLXYwh1y6LXBoVKHSiALL+YHwsWtFFtWZ5l+hV3TG9nduC
KMz+YJC1OD5pK3SPZ78SR2kiEqEoCmzCjYAJu6eC6GQWwuYdNJAk2vHh1UB/Pdp/
qRI5rgzAdGFJHVLhW49pu2hQ8N6fbPRrtXSXzT1/rKVGCVwmb+34o8w90/KNVAc9
aiWaXkLocGS160dC4LmulhTNX6CroVVg2++fVvAwCXIOC+H+3E9VDlOS87bsd7xz
S2txC52GWVH0CXJcWlfHCMjHdmIODQ34bl31WhdUA313J9JkOOci0gfTW02Hfrj3
B56dYR6eZN/0XYKiUUm8GhDk3OQcHgnMDxcZZldxdzg9SCN69j6yVTAw4GgAl7/5
7TSS0Ye11cihUz9YnvVhCtp/ldtIv+XJKLQHtljycf12o4BBuuDJPu6gI0N4cPzd
fUftSFp00Cc5PRmJaRjTH+XHKmEIWPVcRWIvbm1yWK+yRCss0MDpKP54G505b8JS
LzzJ1ppMekxu28ugCxitf7Tu1Y28EACVttF7v8V4oG6FZKKAGfFAnSvnLXSUghWj
ZP2OaI4a51eDJGm4N/ClOLhdi2OEzgLqRLEi8jZRGGe0yRWXa6ZwGYsjfzwz8azs
c5DqGdC50HkkxtzRt8sWLFgmAXWcIxTUOyn4LLlhI1GGFrRyM9BbyIuXi5OfZsS1
Fn5wm5MXSaiB3UhtbYx5/HSIBqzTTuvwnLCY+1gJauVkz/ZyHOE/aGFuza2AkfOv
7OOAuq+CdCQfah75lrhMQJnunFCyqiM1V2rfSdViMDAbAQvH4Yc42Ch1Mu27M4GO
qu63VyKN7N0cwxRlkEDnvffame/iX41XzY42OjMA5NlJIUbe0Wq90QAU2n1e/u3/
fxrU8a1x5Xb7OvQ2k1fa68C3daaptEU7cW0YVDQJEgU3VLjUjj7y8DJTwusAZp8l
0zuY8vRhfUI32DFUYR2wj02VW4JBSjrbrjhP9jkiN5PXmD8xJCmOQsdsYKAkjxyy
F7OsbW070mMmbycUpu98r4Kr2YM3yuSaoNe//0Dcb3wH8fimWV8dhhT46CqMyI7c
f7txMSnKzJXtHOk0vweSAVr+mojIl6lsOK8TkOZjUIj27WhQS3Y9VgE6jlgPYzH+
QxYLwYH8LUd+O+gR4ah42wTsjOZgxOgFVLbF3T6trWXhxIkWGbNsvTOgDW1Poj9B
aUTSY1WENwD2HGI6mV60Q9AJkq2MqT5CBEs4dw5zLDmgMX4Jn5Det1Z0xUSHaeU5
8ao/5OyPhaWTN0xVYj0kbVI7S5sxeYVcVVe8NNYsXpaUr4jrSNJVz5Xhyw3dR8Pu
bp/Xp6ovA01aoptL0UF4wudzPvnArFSYlcEGxdN1Nj+O8VLCcMG6V+fMMiIwtSI+
MWrulopwD0nIQ9WuNpO0yOO6J31boWNXj2QBR68eqjhquGQtUczLdOdSX4e2wZU4
d3cj04ayBurO1Sfvtp9hvsso3f43X+smrOhT9GcNvLJ12rebAfYe8WBI+ifQKzNQ
2yh/i4iVAeLGE42dewQMsd6aqdc0LeB/fVjJijSoC3PdL7Xpy+hdVo++hxF1brqg
5Ytig34sFKIVQy+LcWlNIiY6EK0j9Zb4iZJenl+wsxXRjkFmw9OemS4zDP7qNt/d
ji/Zvsjw/PZhseqyMEKzJywm/ksjTJbQF+/jYGYZJkUBnsntM/MWzrHylxFN3sig
RafV241n4xYow9Qj1pJbSbMjxGIQNqbrw8R+gxLaljeeNgDXLcM5DtPzUmwLP+px
ExvXJfLsClXF2NFVXJY56VoftwIEB6bpPf3GA32qvguH8xmy35ND0xrrNwMePHXb
YTiozUJqaW7/213Vx60zvUnfR5AfYn75gsI+2CZ9IhNEJ1S2Vsger7o7JnfrYuAR
wpolg1Aka2s3J7TYfxt0p/gnqK4TmZ83SmIT10mJGgQmO95HeY5vqx9+yhikgLHs
fO+pA2F4Krbf2WnCdTzqawkKQ6NRgCIzBeED4Y/a5lrL0bKYvM/oZZkC3U+CtPVc
HwQlXeo+n+OWrLs10QjkS7u4XAWt/IoWtK4yerKnB94FPoJglEuyxL8YcOFH7xxo
2rqFGvgGnlZdvwJQiLZKsipdNVT2HMQec7HiZgsa693abOxlLVG982vkgJvlhjCR
2fCm+NYM2l8H2/gCoW+7Bk0gM2HitGS7VdSwqjwccg3WqcxKE6hrhLCg7q/DDh4T
L+SSHokpHo5fXuxGZ0iKH3swPlMf25mkM9QXAHgFCWmzZu4al9KocxTmyM6XGTfj
9dzE8Gn+GFcm8T3Ki4o7hErNfRdu7Iy8vro7+SLzD2ho72BqYAETc5h83Yp2kFYw
YV8aqeZCyK8SNM1uD+0EDRo8c/vXNywVNjcda3P4L92FnatWMp3Ptoiksn/l9a1+
dtemvIYcci8piKfxu8yqCww+zB3wzZuxOx4kcj6l1Bgx+xTOy/FJgGEcVGrRMnzC
TKlJZlRlYcQ7QTu3dbYz9uiNWwuSINK+rIKhe8n5dCKFYSm3xdit4b9LSgre5zgl
EmUpVDwSl/zK7VQzpNAaS9jh0EBLDWOI3r1Fn/cU0jTKA9Ma54q3jMnxU1OtK+WT
lLQtlEt3VquxgHLE9K8rbzZlDAiRoBDZHRIfG1iUFrLOjbHwVzmDtkaJt9fz4RyC
AqYRHcJkb5xhbrPXOl63u1wOTNs1etgFOyEuolemXxltvs14i8C5o3j0woWiZVGh
RmoRU2EjdtnM6gufhCazOPZshmo1Qt3IBuEsFv9EprywquJx20nb80HyOr4BmADI
pmO2BCBAkq9tLJKTuRCLSRYOI0q+XFRmI5c/iJjXb7D8EgP2fpXc5VHYzXaOWaww
kRGVzgmq/rkdIFdQ2MvFksBrbKxaN8nQS+mIomvnCLd8AFbzjGeq8kEBcwC/08B4
2KSPC5osJW6ClcNJajEq8JOr9ofIqt9KxG4AgkWMuAFniBC05gC7u3cE2/vdOBNY
bOz6A/hfFceLXNKXq8s6yLe1Xvv5d9pRVpcn78fdfZ81S0TX4+VTb1qUqc8j6W17
1jXcXs7ElorL7Ui9SUj+Lluw1yc2fA1C3SE2ZaypefW7zeV8Vx9Hw9IDKJoyHa1y
yXyzHv5wm3PJJ94rRShsh58WnCYId4c0/AqO77AtvqlqT2Jnk51/BT6cB0QCYKaj
Mjx5yL79ST0l9faRUYEuCKzGDsIHA73ZibpLqqhfoOy+y4nHUmhsTTXiIN29Etqx
96ONGWY2cI/6naN8Z0CYfnSOATlgYn/J/lzV7+cCR1p5W2wHXObrttX571Uup8pR
fv5aG2DOutClKmO6Ha3vuyzTxRunSoflxKxZAEYogXrX1VcJB8b/GUsE8/peqXop
zXBIOfnecrhSuUsHSeGPFFqNwHFKuEUIn2yTh4PapmpmUxLRPdZE2u5Z4eMIO3KJ
Re11d/LMDHtHoYc+KkjTvpjd6a4fWcKWQ+UXRjahNtperTu61zEIuPgBMEKkLfvr
0uhEsSYnw9Z0o5Ho3bamojWNjP3HoPkoluE9T/5zS7yusgUrG2a70Vun640zOslP
oIibAznnJX6a5B8D0SNm9TsRuQj/orF4UsJEuGjPHri/0MqgbP+Gyo6AZ9eo1QV+
qAIk5g+uX2zmMVZtyybD7hbXt3C2SZXogoBkMQq0MzVQ7v1bjElzWHQq+8wb+viK
1qLvKc4SwC3iTrMY+h5op/6iTREe1mDYHCpRU+FCr9mCQCB4vOeoWWZSLyzaIWe+
v/vh9yhYYUXm5dhwBbqdBrBFMiI1NKQKvvRBsawyIC2wdV8FbynZ0QO4An1x7s4X
/9bAe7IgCvPtqVYiBvw4LTf/1aEXXGRZDWCDMmC3uPKA6ikS1PPSI+WxG5w37/5K
nOQni+Mu6HFMkB41dO+FMYucqhwroJ3gIiWvdYfSrW7e1WOGDQkihURnFmH36Wdu
tRD/kCI+7snLl/6UgooeYhWt8Z/65ROsSyzi8a7opDN7ZyfA7b1OKdbnL8G2lEsU
O3IavN5mjt4ZPMMqxFW1dE0Dkb3NSV6u3+TE+nd4vzajvWN1G8hdssiEbnD9zrpB
t/+IuO64ndJ97LLmzzj6nEKaYPYhaggAa6MxhZ5ofNyKrnygqyxJjZV6y71nffN0
aEFy0GYYmxMmL8zwmI9NterRns8Vwhm2CwVm3VTstkHjJ38VJgG4ueEdu+TFzj4R
KJZZWyIDg/FebE6l88ffYbRnscxrEJzgb9k8HP5BOcjTzjEsjmhKg1ueVRRxJcWR
/8OaXbrZqhZiBxzGr6HVQsuvoav8mHrRdsknOZjstjJoiPDOqulezYKQnb+rKVpW
50Vk0VfT3qovSNByJdECWT/ZipXXycPGZWAbPnMj8WVkjrDFLO1ImyPvQdS01o4w
DKZlBmmXLWrV/THiN86dWCs6UqDYX7rFqe7ydQdJ64essgY5nLmNwQdmuTJ48KcF
Sdg5PmfUHWBBJO7ygMSlUqdG19lqZdXO5jd8hBiESxe08KKlXbonOvFfD2vKeKQW
nFZaVjRkWP4P6XdHLM4CLQoyPw1T0n3tD3HpPKtRS0zlBU2RJxEMVLH6/4Mrw47V
mI/pAv93CGmo23poUv+alstJlgO56/9ZPi3spL7PyFIPgsv7d33vKQDDHDMDSbiC
24m4QhxOzK3Uf8OSgpFukjpzo5uhKAVMh9XJeLA1Qy+ieMYUcaY4Sd/QvEdTl0OC
el0WDJ2iA0yNsWSjm4yNg19HYKGyVAPoMQprlvXzTW8vzulm/yOURUC7p/JtGEeR
6zIr8hLXBCaCSod82lAxn/Ci/d8AmJ4JGL2fyNnsiUur+fw7sUYuYZsnGv+CEZJx
qLRUQul8eZJzmVgzx0SqtzR7ERawr4guylCkf8UJv6aRCeJVFEvJ7LeMhosG1w24
aMs5qNqxXtUbQnIgV83rIMQ3VULBaWvXB6HZDPdlhbmW85cl1Afq9pc16rh4hv5s
TrmZtpju+Ez1iSXW6/5gK99tolamb8dieId6gEIkAP9M2dguQ74mx9K4hMVn9ieu
zJ75MgE1a2V/l3BrMiy9IS6ycc3dx1rrnusUQQJKvYZ6tYETi3CK94gi0KsDXAAA
t8iVFlwyBrqDvVVWZmnhqGxzAEpuL/jFtOOQSkesdxJQM5Dl571bv8149P7/wCHd
Bamzlpa8HU5YMtigSyBz2OKSIk1Do0ZO6SQXcq3dOi8EdcZveBC0FJBqCeV1FEWG
GVCI0QphQCeT7Ncgmf+nHDeOYZMD2DHKDs4eSi05UZ89+mWu3FOYEBkAFxxpAxbT
6UcGx5/AbJgnPLzCJvCBfS6hfZ31IcAIBAQYjD4oNfIhtfV9p+CtmOWsjp4J5Fbe
9oc5/bhKGrPDJSJzilAutX55sR8hoFBXLX9NSDwcvFBoJXGhlzX8wk+CpMAR5SjH
aDKbDh5aqhAX6+Fq6+e0FzbZVzgWpNuHgPZaGElHJMTpDYQ/wBcOM7c4NshRj/zQ
nfJ4zK6BCXTIaCqOVSeNMs5DGU5v7Ck2FhYknpROUsCyOWmR5ByZX0gdf2dZIPPf
bW+zz1M3GfDFt+JMpl0MZ+0BtaFB2ymiOO8Otlf0kyW9DrsNxQBU/4XOwQrVhIlV
kE3CAARqOKx4+mORPavts6ZksMXHdIUa6tRfoniZcMqf0XOFWcz+kbAnnrtCAMiJ
UqqAc+HDRYUcvGvyFuLnk63GzYSRR424H6LGRvwYygYkskUdDPAQ/OQMX/UZ89xQ
mbW3E9CRkOwgfZyM1lkbskhPjDekMXacs2JssXfalwU0bgCsbbzfa0NeF6rgkc5B
Wf+IobTD7FpFqpOvL62Cped0gdXSIuJmn/I87zSFf+/dB78xxW7w/9TwD+QKwute
05Ej+t0mAum+HNDq/+RMAlVTfHIrOXqLadls7y0C3nRHQNRG38zop0MuGBL61MRF
xt8b9XvhoMoSgFqF4LncBwMi6ezjh8CjAwJ0++fqR+1m/3Jva4+54AcqOhRUad+F
jXwi31qOFe7GyNQEyK5+Ijyu0iAzW0L7FiB8QLZrcjkOTyEbJTlUmIDUkIPa8kDN
84AgMXBrsUc3wJJIQ+Sy7l856O13AHK7Sc2n5pO6SxEeDTd/kkRXxyAM/qWlhULU
rDfsnHcLbcGO0ixMJ+A4WAnPbGQEOs2C4ucmXleMdcXhdsMr/6SNpXodjk9/W63t
Wyxoz+sH5ROrd7Fhc0nUi7ACkbHTE2n9XSS63PjhvI3LlH/i26RzU0lHtVQqEbDS
g+VCmlHRc1QthVlI+8QgicyROTWfQHKPaUSJcwH5zPSry1SYC3r7AKCY5cRO2I0L
Mm2ys25RA42lmRSjy9k3crOwa0wX9n3bk1rRdeZc8CjpzzE+hdZw/9m26NnyvxOy
Hprlf91xGywkAN/72wFXZq97SyNVdqyjRHZ/R8MZtsiPAyTgjAOzBkismozZzh36
/Q9P8Ax4sj8Ec4X16Ztzer+0NQpJw1biuSUYQkgMijCak1SZ/gKtFLdZMM67rkNP
OTlmWpDMc4cbOfM7tOTqEIcovvK11zUvZjImxi1ll4K9IIV6JterUVK1O9OSUN9a
r51oeSwc8nV6AwGaBmhnfvoW5GgomDPExOrgOdxKWcJlGwn/JlMJQb8IDeOaEnOm
DA/nqiwnrcDgk4mre3urvUlYaFhnE0+rp9zLEdbUPYLXAV6CF6KrLwQ6CjrtwpWE
C0hOGwIiygfzACGszThiz7ydxPgvANBWR6Ck1dBpyPCXAbJafWMdyn63wc9Td3uJ
myUSiqtSrsjom6JPkZu/PCxhk/rdYo5zQ8O0C8Vk/4V750RnnqRcK/PL054oIaG8
+YWr7CUd1jLf9cxKR1T5G+0gsH5qD9JV9c5rkj/MpiWfeTVCSBGH7+hQzGgaXNz7
4g8ldQcLTUBay6ZS1ORx49xrGo8by3I175NNa0GHNPqTpe38FmfU1O1Zd38tc7vj
Bo1Gy/PFhuqGowp6l0441oZAwFBgjVdrZgmcf2hymsmSr3anvvaZi1QxtokxWbSt
3UBSIqn+gu6wbRMBau0WuiSzZBeSZKvvdiDLGEf7AL1WuIwfxlcQjM5EMdS9/U94
myIIB8tRFhhgpAIDfqLWOT4F12wcLZVc612APssDHlwzwxjcapi7x/kx7rdDmObm
Y/wA5Wt3BahSzEJUIuK09lv2hhKsU0GzWUBjoJwG8w2NiMWbgGf403Ct5BxSDtwv
PQVhsY69huVcHsSPLRfpZjiPT0XF1e5fz3i9MK3cz0Cw32ODE74SVULSh8tNJ4qX
WRTqiMrwKlYgP9ne0ICK94Z6Wl1MgWwz2x89imlV95AWtbEjk9sVaeyvRTfxcazK
SibARuAk0O4cHmtb6XxzIQ7l2nE0XPMF/zmDWcLL5SUhrGLu5Sp3EoTneQCMOwhy
mHeU5NGJ5yn04ajV8Iu3hKUIEFeSZjDknQe1gvpGLCC8vpw0aDsuw2CqVHx8Rnga
oK+qH4SDoVrAFBrIH8YhmLFJHN+bUQGGMm0efrgJz05I9GM0t5E4Y/BGxnJ/pqu4
V68oavEf90r6lXo84KvADuh6nIEFmMrEhZTSWfD+kpcoyoUC4xzEpLJs0mx/PLy4
UvDq2hRnaVZ+YTjsp08+JJ17XW7/wEcz0EwKZhnjAnjz+VZf5OHM4f1Bl45FrChF
F+z+mMtgDHrdJS4iKlng+vZThmtq+rQCy6p2hpaMOfNQdHehPNx7fuum03IKDc8Y
Hk5LUO9rQMvHSy3kppIX6sr+8DqxuMcGlwwICTd/XN79ZVjQcWGXIdwMgp17Kmja
0RnfawM8ubxlAxobm60jARsg0hukvMRB+tUvaOqpJfIiJhU7MkfSZA5kgFg3nhOC
3aS0+jeQfrsB4573ORX+/JknDXqjzvLU4XSN9CWr2GlxgV3/lE1kTHzQovmLIJES
laVhepfIHz184zp6IbynaccTNYg4US+/O2+aAJxDPiAdvJbOA46hWMMzd910HrsY
RnU8sWTGVpBk5qNG+m82Yb6/vtu8r1q6OCTGj8oYwGG3jK2v/oAajX5tv9LhapDK
QCSBF+Hw+rjIdK/bR6pSPOxdQEcvPMyTihGdGewa/tSS380lbKK0B/jpFTYil6tg
RntLe3aXZg5cYDxDH12IDulE1kyxKzyB846wNMtaU5J154S+BT/f5S3lE1FBQs8z
KTsu6lv/8Z9c8QRYN8z4MB3l1VNYktoQUdiSQFqIGaZMtAwEK48itNT2tBf2rJgj
YeaAexh52UPLHCCnmRjYp98iU9agDq1X5etKy78QR1CI1YmiNvTpUf+mM+Qf9GMc
EkeArFfk95cNeQWU4UX5nYhhc4ndcov2AlplXW1JSgXolDuV8FZ4XWEnOIVInViE
mb2q1Fg2AwO1VreA+eWoEtpHscNbtqqLNLXLxTu0H0l2IOwDcMr9CnpSitT/5yUs
mTXAhhGv6gXwS1OnlxLtU9FNBfckqMAJEXe8g380o0MiGS9o0X7yx/VtiiMKPzGP
anPIH7QOB3EnphEy2vFHGfngBKDsY28ypfuPcft9KNvQVjcWx3ejadUBN5/xOGrY
xieTorkWawZS0PZOX18FVUjTDFpOXaKroO5bBcD0u9GHstHMpn/DnEBWxICZuY4g
ZaRDdtA4l/zY4lE6umQCw2hfbmDPzoHvZf2jpkdFQz3zuVF9nefYBJOI03QXKiTh
+epVjRxRDkYiJRmb3Wxgv21FmgaK5ovtIw2/pnC9EpBA09jTnCYqevsFWEaX2BEa
d0clppV9bqnbDw7e4hwbkFW9G6cAw3DetlzXhAHRvIv5khs+vwsRzPaQzIFGRY7N
v91lX9GyWi5B1Xj1JcbcrOyKkAb5gSnsHYEPD9RYNc1Qht4O1Y+FGtUOB4Qe2Gf3
qV75IFdgWRW3oxJ55dixfr9UWhK50PDFjkog0LJXLW4d9ZA5RnaoPRILnNTdU2d6
0Ey3i8a2srkTVxtwAbTKLbCjPZZr4gchhxAbRcPSVOP6HElPZq4Q93wO4jx98Ipp
tmaoDRYePEBQBlt9S2FnXhpQtP0Uo3BfisAHS3qdZD4ge93F3AwHXVNLjHijEo3F
VLnGkslVwxbLe5Guv6uyKKtW8R+aurlLuWMv+V/7sePZG1nYg2NynlsaEEStdYKe
FOphlGmxxtY7gziJmLV79EuG3v3HUh+cCOIPwedqo6/bxXyB1xqDFyLGxfSShYfz
An3Ktnuo48/ywBhRdtxbAcfJ95FbhOeX8qorGgE6jvWFNPsHaQjdEdA0Gkawh6pD
y4hKzoIf5zcdoUCZE0zdlwYuBMgVtc97JsIdTQZMSixJBJS7+nquwILE1teGOeR5
u3BD3+lOhRyrmhfOUdHNOLk5UfmwDb5dZrH1dz0Fz70ooODUzVmhhsOpemiAkmhc
1wrWd5sY+lPoX1M3w4meVc2D/kdIG7S+KpIqZiaZjhlZLqBNgpWL17MKxmd2/izi
3vHbGHln3wuTS+MpACZcbKHztiF1Ms03FesxwXiJ85k9nfP24Lv967fHjY2RHvOB
JyZhCMSwfeaQTQfbjB6461UEzEFFsxW/hLbuXS2+kWrvSzvXoiCQfspJc7mKva/v
MHSjV5NKV8C7EnAAOgMQHLzEP6RsAYeeReTDsxcaUNIBtNXiOuKrPP43PzUYyFjM
kcngGejfyv+cZuS1lkSO5B9PQg8g5vxOa14hFLtAdrnJQ2t5J9qKdtk+tRRenD8d
D1hfLzYCY35ykaNFDFTbAP7gVZQn+V4tXXaDii84aAHoEFMLnvoMZhLbw99PC1np
XyDyKCiCKEjAXR1aFlCS68NOWnXW08hWH6X+Msy7HKAVBRUZc+qgf0QEBBUPTqhx
jEG8Zk5Ky/faBJIt3xFi7BitYox96vR6uS3ysjhPwQd9dvPX3xOrnNXDsV+boNTL
eGeSUJ/fAND7JLoo2qpIokGNsE5G5bnF86atJJ7k6K5yi03EvHzr8tnHm+tbGfI8
d+pTdVbhOfBUIGj3glH7OKTTkJEHYg0sdPen3wi7CClVFls28fTvwdx0+4ak5P/D
wvE681HgrMrT0TupMIpIZmjC+Xy4zZz6gF9kVEAgmk0LWuWgWKCx4oCzEbM5kVbN
TeKPuuwr7P9LNf6ySvuYb/47P7gtuG2OzBVy1bvFOefE+BSNgvHBYh3uH1ZcbbWL
h7mn/NUJfdxfcrBf2Ddpgezw6chgS0ahvZ9WxcN0miPMJImpeqUs60LUhTXxXysC
uGctUw2vHsVSCFXvrF1KsAyjGBW1ZVlUK1fcdN9qo53m1hbthLOmHjdJnWCtiMJ1
A2NfCO2RzZNaR+GFCVSjWOOlfi+LtkpZMW75TYhCS7N/pPjudl04kRUG50rHtzrq
opdiQkfH5ah6tZneH0qFwdTlcjoy/0z6AS1lb5x9j8k4+P9EhpLqzFPwR3pgjb9q
9w1ACVRFSdnkHaLtZpiRbWX9Y85eqLhc6FQlMncZOejVxpLFHASA2cwcbil5Zlf9
lfCH2cbP1dRQ8ReGxPDjRK57GtMjcARfJVLUeiJEdMWMCHReyejOEmUfCaGwEbMl
4Sm7tgRsFJXQcylGROK69EJMlAEwh35o8cGe1rHrP+/3Q4K9Uprsz61aHCggw/OM
GFLLaf3aXT69jRiFnjXS7FAqeYNvjpVsTUisMl3HBbxt0hekvfXjE31kdR36HPku
8xZKGONWq+1MTyyeRpSsSrHIV1P843+/yKQI4sjOUuje5bnr4IUWxOS1bAOjalKa
U1eBRSPE5cbEvZ5W6ObZOb0NyxBv85HKLxddGULJjjgeGfPthaoRKK8bwGVxosme
giwdcFmjNfYuR7MhTsPdGTlF5ebn1ZVji26Kzc6Wb0VhEDQevHSlu0mnoSlYyxON
yHdosKOwXewm0zYuD6eRTxSh2kJ61hGd91PdZ2PrwHbO0iA6lirP3wZmnjUKlvyw
JwReP5/HirTLYrSgAlFOGrlkYhHYUa/6HeEz1k8DedrQ7YkoO9hbhVpCi8A2pcOq
Kpq8JmtL+DydiWaXQsbjgkS4sX+Awy4ocLmu2HjE0D/PNHGnbsdJ5mCow/48z9FF
jeh5RgS4MviqagmUPsMq2+1cPzKdQotTd6PCjQJ2yeHs20h/kEI8yPDVuz5xdfCt
TkIrOnmHfITHAR0oOSEFXw8iBYHdC2k2UOwGB26FfD3oNteqw6NtPKdXPZqi0wyL
wzJp3KIXTfULPAVLo0QJE/TqE3J//+WMN5t1Xqhdj+refPn+M8pINzy4DB1ySMTV
SpmsFu7CB8qM7IdZuP/bG9E9vLeqLm7HpVIbvyhKp+mwo6wKovD7xhyVe3Q8i7Mv
DtAw9VIDjDtn9lZwKfp1T1Q2AHzem9U+qlR5pfFHg2MU/XOevwMwz/mjLX+yB5BS
Vkcq2ABE1aDKwsF8u5v+XvWBr9vprEZxmdCU3z9gzab3DemA/JndaVL+exG2PWPa
x6KiLmzBRsq/N2XNTpZvzP0ptVjILYp5K0cFIyvrixbHDfkF/KhlqoV9wjuvMGf7
`protect end_protected