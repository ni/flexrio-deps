`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 57664 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
we8OvAuq+6JGAI1WqVfcIPa61hiAr2MPjoarw6Hja4LqVvkXUPHhneLWLC9ldEZH
94HwsrE7jOpkEjrbh4bLu3iQwbcrIBEUhyZqERiSC5oKymDINrA9kdklXYOfLIS9
rllggmm8e9BbRsthhNF20CeQ3z+G10TVgz5cmhXKny6YtLubdhhbsolvUdtPtcVE
yoviYVqle1R+LCrtj+Xecbs98EnrKYwIOTQ9YZIAnd9MJVireYCSlDMa0Ai2kxf5
hd1vDjhUPBTb/KBXRAVxejvysn+zu+PYiolN/rEg05zYTNzTm9P97yWRoZ2p6wMo
1uIxrW13GudZ9HlCJAo2EhpRacXNLZdSgRaJc6L0vHrSSTbzaHeah2H7zLnp3ZM3
cvoHyww4tQ9wLS6u3ZUABiujSM6PdW+Fk7nuuJNkNVimLUk/Oyl8Gqb75tB5lUxd
6ZAHLuHrc7ISo3FnDfM39kDRIPo/1qgdhrvxLvWUYszrDT+7LgnErRLXPeg5qbqP
UcUhGMvXcpSxiL+piQYOncA003/gCoSfLfKv09J5wrxGWSpXn4eWKzOznJV8mCi4
kyZpv8+2a0rkIQqFqK/NV/ONMegQY5etdQQb+zTZaI9Xw4ct5v85N/iXyxyLv+k3
YLr7Cl/sBXLd7Q9Nhvtz8twhtO7DuMIBc9Ly10O4QR+4sqC2nIqquEg4fSu5iLAf
jXVJCnZyiiPe2YRGubnpd03np304hgGOJ4sFgjGxoqDKHHs3VAzRghK+L2j5wXlY
BDtMAN97boufEDGB038hIo8PYYtj4jLBIoBjX9TaR6wuHkrXZ2mqsd7/Y3G9OuRV
j9NVrF7oBF+dc6u+VXP3RrFgvgePIulgtE+Amb79z1zkGb3r0MlafvhDZ12CfrQr
aT5LqcDH2GIkDHwVGyEm3fymj+1xl/7jajhd1KibgxY4f60A1wjQM7R0wCSnMeRT
PFwiWuNU1hSysRL4ntrZQDrcQ6icv7Qm0+IbvglzlRT4MZ862wyqDYqXVyWngSLF
XCSk6pXLOxCM/q1GZsoo6xfYcIKj9hTppSHERyc/h13SDD1y9uvJkKk/a+e5ATIw
wMV0DrKlDLSn98lO26CC3BpBvfL8lBuvKCpjEfut1/oov2erxEohqbSf2LmotUue
DH+SHiDyWfn3C+wSQFSgRJ2eiWMhiX3X61Dv/mA+nFDwUgQ5mRaJLE3pZB1WyJfD
CmAvl++W9IWL/jA+ruz5jG7SN4MC0BVfDVgKsyFSVssxGcYKK7UhC+Re3I/0n+iK
FVLpPXL236NHgxlhTsRRRcW8XFCRD90yjr1NFOw+wDqlzSbs4JyTnhoQPrsLP8Ax
e/1tju1uSnp0eIAdFiJwj5xHvQpBV0qFuYc3+q0UFq2l5yegvoY1wdx+nlc98ZR7
0wqP1IUzkQT6kBsWVpPgkd6sICQCQwrcnwU7Z5UxPWRd66hrniE3H23K6nvZFgPf
cAKW8d15HNMFuar0RzARFsB1jsh3m+43PZQxqpHIG8N5O1mOr+n4dQbP9LBQuSi4
GqOlv5RNstX88WeazRWbROOiyeMCi/IXLKZNyK4/iQaTrACkZUwpaWydkfGhpzdu
WdxvHBX1Jt/EfmFJaxfrveBddZiw2sf+hVz44mQBujVJWDiyK8bhoq2ZdtnRrJer
8As6lt3qLCGTIdgawFYmouj6K75mP1X1NUu8Gk7EVY/Xc/5ZgJdfuUGAQg89PyiJ
ZkOR79pbr8tW67h2KkRo7MeKYVPiVLyRWbRSJw+CTwJRKmp5b3t3c0nIXth9BCqb
LNPHDbmkHiEel47dvwBU7K6YTz0G4L3O0HOF+MQWm5XCu7IeErnettkwkI1I+lIe
S1TCQ66Dso1bDEQzCh7VCfl6QT383Vu4qTDGr8gEkSN+LLjCoZ7eW67q/jHO9S9g
ZsUyTObgqIFRHYrrTeE2IQ2s1ZiLstk9xHFbgoEu6dv/GKAreyom6itnDB2ttM9c
VZdKpF+RweoXC84LYpxebV2+aJIPhu9/WNYVp/0kxCu10zK7tSuDW1OlpYz3aE4k
a4CLzv5Nphap+vbyigwrJ6rO6faxobmF05EP5vE4BUCtiuqTL4YSCX+TdKhVXTFf
9hSHpTe+qSM2wKngEL56QQd5Gg9JbDa6jhxFfVf0CmUF98KbC8qKWE+/y7N9pYBr
M73c/NrEMZOiFHWpWbcVx5dn1qmdZaXZ6aDRMJBoHWmPDk1TX4zWYttMCDFfxMUj
HeYqV/lL3oVGMt2JowxEgu9L5QDB1LbwJRgkrAXynJR+bwomVXwR6Uz5w/ZneCPC
wHoIq5TRH7d9a5tP8GMoa5L7X64mM4ttxjermVXSmnm2wjJ3I+j9I06nc+r6em7C
grokbWkHjG7zm7Y5F6MY6nByhrUe5SxAVDE5L9OwB4hAhBMvOd7ntyPpGOs+/nUV
4hrvITtSHPrkuuPGkJZlonvKFi04VGTVjWBfn00eRcijzFnjM+LlHnGRIB8jhsSp
23jq7JTr17rTyIct/7cwSHa26DREwndyoengkdl9cTPjsYwUFWvYD98Zc9XdjnJb
6KDJoxCY1OiQrtzGK07laY8r3bmiEoeL1t0jrH6IoBjp5cJVMjOyTkfr2maoK72p
vgvb7kdKGrB4/v1cK9BQW0YwBZVNL5z0j3pJKShNkrc6PATwLWAs5swo6+zXZKqS
lXBOfWH/CvP4hUaJ/2GTdvEHGdEPjqgaSvXQMYxSL5Ay3t8cCiMW4iDTRWgPYAGW
ZJ7LDvGzoa9mSpdgLHNJt2/4NpU82hWre4ZSCf6fXB+AsyM4+EqlTpLPtcpJUOf8
RSZKkycuhUVO8qICr3EWmuuMw8XoyPiSJGYAkFw8MT4bHtWrlwkLXLFPTyU729ri
BQKB3zGG8Wgb0suM5dpYhMNzo3My1uvU5sbNfXPOXCmocSbwGHJ0FiSPiGTuDhDu
dvYCon5Y7ZnqwSWKnLXdNFz6/g0fuiScRpB5qSNvGY28EizpV0YmSZNdaDFu8PY5
F7YVHWlAYm7OaIk7TSK9zOAW+uGAX8uXRAJMkeIoilHGhtTV/HVYSeuGuw/N+zGi
J+WtSNXeoHOrZ2JrEzsaB8MjtHQrVSaTotTrS3HnHHV3Q6AmAtSEXz7Z/G1q8lmo
kCPPj6HViIyBIaisc+FBruWxJV0uLAXBtQUE/UolWsvVP1kPJLF0kD+ba7QhmhJR
H0qHVoK184gRlhLUr7DZ0K5ljtNDXfCDycC8ApTe7AcTvsy3vZJaopkwlyZcfw7I
BnLrWOeeaeF91jkVIoFc3wqgY+r/H6LrW1/vcaf3B72oFFpP5LUu5CGlw1bKbotP
IQxw95LGy9AlR6P/y2I04hagsZ4SyNCLGDPVn+rlIH+aq/QdJ6p5l5aKzLpBRFrM
qktD99eBkHSLnm4ETtPsDqJuSnqp7CC1qdXEMgoqOZciyQi5bBkGkEILU690I8XJ
MenpBdudDb6x/FPuoMCRXDmJki9+RJUeHCz9T+36QCbYmmjlLg58fE5MrOdDcm46
v3pjC+DpWsV7S3uNQ1eGSsgJYj+Yhv3ShfObi/Aaii6phcvcUESNG6Fg61p1G+yr
YsvpgexZS79Hcs2HkY3rUMA/G3DjgeEeRGPHOxvqXuXKtGtdw1pymSzZ7ivUoZcb
xGcMyE9ZUKeg+re8hUq5Sl/lykAVtUnZ7mzb8n+OFngu70O3/UL3sKSIAb27LTTT
z5aOvocrlcD1cZZzBScbQUYq5aRl2QzfAtv/CNoshXeOipZ4V+xWDuxOHYi6lPEc
jLazdVr3FdqBciCIELYXOtenkUp1vXWN/RIXfMXZLa4cZk8z2OHWbEvBRGbhhYgO
MsdlCvNGbpHPqxUQhIbuj836pIbHqUKYGJi9KTH3jfe5occdoWwhKJIs0ptqukaM
rWltxhuh3FNbWr2tizpJhjHq/msVOVMjzeiKI9zsDkKt5oLA9Hd10T6UrN2l70EY
ljN554Gt4Oy18XFQB9ZqklTic9jKCrAlYSaNj9M1WqioHrKbm4U8NFNjOHm5yAul
M0pR5rj3hc9UWX0U/wQQ5NYoV5oY+oc7YrZJfTKp/GMFcWq8DrV+iFqQnA+EDdiR
SXLr/tROmsU+KCyLbfWrJiA3wxJHQmsMF2Nux5+xN3OTv0cQhhG2pzAQfjU7af7a
hwMvKErD9a/6OoPl8WnMakgQW65eh8M+65esxsSc5W2awNF63EprR35POqInl2Vc
aEoe5AH4XR90U9T3VERfXbVw2Yv0UgumlxqwFuLTVw32wtE52Q8HnBh+Y/Wz/8qn
NoTDCeMZzgZoDowy70UuuhNtVp62vJH3JHXTMv5SBDMsGcLraksDofGQT4BnWaBd
zwVSE45f5Dt2jB/du2NdKFbc9/xdkFtfQGfHhR9J/PvMmWsqH/tbox1khFONs2c+
DkJ6WKfv75/T8WhmPFri5bzI2PdDsMQyQ/XhsVBKXpsJfrl3rXhMBhxE6/KxLtjF
BMRSmvpPwdKEmjAOuiyld1M5G/0jyxBumRB8jpKU0O6c/Ts05fax3P3G/RBTbk9N
eYBsFJUXaQc8psZWj+Txre1F+QYErrqdtJZdfRkLQsk1DaU28saKbOXwfy5wH5NB
lOaHvduXHUHMHE+JpbMMA3DBWCpsYCrwtd5zNwtCWJHE4TzEyOahdL979+6SdRmu
3BGc6tmm0V/KcIA2ui+MmO0ghf4Rx+uz+ewX/K3iigN7b1ojQ/Y+DEEwq+bCydFG
8fCPKsURf3cFaHHdtehHcVWGP5u88z5IZFhpydTSEERR1AlFMmYS5Kpn4JFTeyOi
sqffdItOx80UWttEhzVwNlTtEFN4ikt8AhgAsPlUfmwV+D2HPE3cDlfwD5skRABF
MFYjiZJ4nBNdk7tcezFG46uJvtGpVzEMlbAiOHOSnsOJPK/VlEhoE3MbNwdmgb+s
nDknqpHCGMIac+b58S+qejf4KlH5m2FlL0m/5zbu9cXJNdnt76cEEjzx62jGMt4k
0f7m9QUYig2r8s0cMNdQMNiogG4uUcvHau9MqCNYvbPuiJ/nhi6QJrpp6ZFSE0ne
H7WJIrNAhl+9/UMU3iPzlh7JhZ8HJvzmO3SlZIdwq0R0C08f6W9h3xHTEQwUCobp
D+TKKOCyWY04c1jZjQGtqBnolVaMw5dbaEofBDJ5VBXCjHF2Z6ho9EWkruv0LtKp
weqcFoP4lSbZSJbe1IiegGZHA2+Pf3rLb8raFPszIFBwAQ16imB/omBlhToYVTXR
iUSDlPtOuP4dVDVHoz8f5qBDiokuNuv8DXsFPRgyO1AW7M2ORlaYXn6RpsXJFTuL
rLQoLfFgIFaDFfbrLDJ4O6ThxPMAlzF0UudG12ycofjeoPjUmW1BAGHe1gtMnwLB
4VHFM1W38IfJjRUucY9zsAuMMLVc2gs8o82J8DzQ8WvCG1fCSZcH27naakreUGFO
BNaTy9cZni4JPdwgilz7FQ+E4fgnVukGb19gVxemg0a4xgg6uRWdXkXebIrWMnOK
DWezm41uuC5Mr/VoRUnNGqp/SXnnenyuCR50TXOFKlOjc0V7ZgTupUe8wJGhPSjL
jkosmiGlRFIOI7nsv0HTVNLdlRKCnjrPReLwJ+1IqT/0aXHrQTScGGJDCBpUrb17
CPqX3ZwY1S9Dunkm3zqpvRmmFT5PdUE95enW9RWZQRV3GKsMtMkzF+3wqoLL12NU
j77KJB80RUY9ARdnkbpxmqJ66k02UCcuHI3RKv2eNLKw644L7RNlUhuhzzqkRjq/
bXOlXBQN1TwVUER2p2mJj6iOWTEH707QJo1gNAgR92fZVkRTS4rP4p4tk8EIkebB
/kuxRZaLJ3lGMfU2sQPwqJOtB6JyojZAN5BVZltKBK/aHKr2U+ivopeX8jp4Ji6k
u5EhlpPkjRpBDRUX8dcdaRTucA2TuaZe4pO8fkAw6QYbGAo8PhSZBMjQFO6rPskX
cI1oX3R503rwC62OjdXI75seUDTebWKrTtPs9ce780whlAr3djgnIMpv20/Bovim
bQ32oPFpPxe+xTVOh11wnKPpvVQ/V2h5/e2b56rWnVG/nw/+sPeCNk0NkUZn5s3W
ZlNw38E/9yU96s7XpBd2ENkicWiSSXULOHnxbEeG4S0/x/O3VJ58aNfELvR3lvxL
xVB9ejyYFcbgqWyQLvfyRDr0x43i9mKOXg/3/M1pl86XrkUq3pqZ0qv0yr65kwGI
/wSLDhiaTqKppaiNhnMYECAOoQovsBicLnxYowRjKTOoDPGtf2og2cUGB5K0x9It
kRepwUB25wJ/JP8UJpaAtCYVFuIUq0T4CXJbs2Yxn1IybXOZJfKTxc7h8cEbWn+i
sCpyVwfHyeK37aEMBe4rZcze91yvU0W6ab8X9nVqnSyQoheRixLOM+YYk2nxv9GJ
6JE83Hf2uhoyI8zXjxQ+hE8a4O16hH0MOBb6Yty30xXaMHpPGcQAUVfFWZKoeyCM
7K5QuRxtBgCfpVxlckKu/fckoULIwahZE+iyt/vxLDCWeShAXExEa4fvxpC55Po1
hbohE7RE77usQcQe9XfSkFjW81EZkz+35BKwU/go6p6p3u6Xje4D9PXc+eQa7j+O
IbPh+e8JeStScnbyj0DEO5KBh3RSk749uLFE01IVl7TEX/5i96Sr7PV5FRklYchT
VUZzJGA/VPeRNcpnwpSMHtJTkGn9CzHM3vxZfwZha6b3QwSEJ8Ee9VKicKyBzSoJ
x0h1nr12acO2UQnpFZ2GFkONbfYhuY+474rladJiOOU5kFfGbi/MUIsvkfJc/G7a
waZ+l0kRJI1O8Ts8b8saJ24ukVwqHrzryjxrcRjWJv6Uu5q75vOVmDAqGUgW5n+y
mtRyEU/pAiY07T6RlZujOowfq4jREU1REa+h0hfRsG3USl9GCiPgCrfqDpXUVeB4
0UgzLDHfb1wNTcFFwHY0rlIbvl44SjPKUN8E0Hmsfkzxss2cvIZprzYnzbnpCfBo
7e1sqQf6iXzcgSi39KQ6HCapsatdX2CgQc9//l+B+6hop8aP9PHjhjH66WcrBRbp
IpL3S/RE2JURBwVI48snIa7rjSuBUkxYlcEcQNMb8AzQIPCd+btqSSenj9Ke5Caz
xCR5iBWs6XlGOT3QB7FzoCCiJ3e9pBrFKUrRP8Z4rwrvsFmUsMxV0uzdOR1qBPLV
B9SnOD4k8DQu9PunrBvwiBHLVRLUkwGrYoVXSv17rY2Z8lSgwr++c4MnqXuZguzE
UWvAGZztffrXRpy01hVaoOL1oFRKGEd8XzZ8iVn4a6tnMoX/tGv4CF/V+5kg8+aV
1stOyFMUM8lBN1rMfsdhaEDAtnhqPc0kd77XdBafwQgwCx4XhhHX3PX8qSfRzYNd
Mk0n4aVK+lm2M62UVvMakvPa4NP31DjKZqNGSeNnPGJ4mAYYsfoNIYObW6saMzyu
vIgLUAbUmTxvZklBiqiKfCATD1gcnrk+FDM3msR7omT5vQkrxB+oPY2jNlWcUMNI
Cs6LfPvxYL629Qil4WOB0Rg/q4lBvh7/s/a/f4nqjNxuODWJzQk1gUyp4XCUcsCX
RVcJymq0VocdHfJxLIBlvNmB0YAdou5fgeaHD0rKNJxJGvKDapZojG/L7M7bQ+Jo
hA6MrW35tqd6k+wyKRnDx1uOQEKxYXoca+DEPP78VjMbUsQRudxQ8cAxTzmPj/Aw
TVqgN7X+Tq02GRX1iSZNF9clH7q2Q9bCwHu1lYFaGsiE4QkYdjwdi1AIzR7kBArW
li5IZK78iUYNmiycNPlBfuSOc8lmIKTlHZwhL1rT96Xyozdce3ttOZ+l5BzO3FXK
LR0qe3VH2Gcv3Fy71r5bvSDYCsSCploXWdQofLAAAKiKfeFRfQcDZxDONFfOnXlc
wnC9+zjF+87c3hcsGSHcqZYWcFSUs3gizwUo19dp1rEm4Fid7uGoTQtTsAjdiclm
nxMq9jb1Pww5/jfL1iENDDg58t7xZnr3Sp8R4nAK5n7A80sNqEQTbSY8ew0jXURY
JaGZ7Xs/SixDMujWDg2p6Tm5v1E54Ip3ZCzL2bM2wz8y0JMJxDdoTxXQEuaIX66W
eZ+3hyUCO2pxj5h0NTwpelzwLXqX8amPSAVdbpzCYmCp7Aiu8r+Q6iooPYaL1MHH
y3nZ1j+23CLnc8/XYXYb/qsXaKx0hMmvSNooConUrFFTuV6EPSAjR23K+pZiV3ZX
OvKVqFE7CqbxEAGHDJRZpNmpqPytKNl0V5OB1TGk4mxFaIddQcGBVUxQVEDWQvPU
hvgWnre+gusH5F5GJedV3oll/DrHEciZtiFW3Tk2sO9/xkoWwhszRo/ZlDU3DfIX
lS/N5qjD1DwyLHE8fmk/jK97jURwI+s5syfpZrJZFE1SqAbbrVTJ8wRumgosTv09
KsphKj1oKkTUyXz50bS/mQDvKixaDZn3bSmnHrlRPHIV+ru3sWMdNaCQVqT0WFv9
bVOx17j5nR56jHRS/THos5mkAnuXLWY/g4y8piHP7x4jsBIsUEKaiaGgWXTEpgMC
o50xllYlN3b7TNqDou9lBuHXarA7ZalkSrkB1OFaF8RPx+kUrlHVCm6hhvfONcju
mE08UWSzmR8j1E20qEmSykuPc7Oayb3kf51hXJJzHC0UEAOvtBCdrtsPyCcOda/R
WgAiYyJLUBXtCW1xwbUq/g6XtGmw/pw6rrGxjd2mXu90qj8J+jYhl3gU5f5g5cuO
WpOWOBchXAR2MTCDKID8bQF1UJpjPWuEwz6knPVqqOl+OQPHXjM3XKGUvAxs0ma4
YWMtpOgclIigjFgF2wBl/G67yy9vFr4LRvS1lktdNl9R0OWLj3H40Uxt7mhXj5Lq
kMRhlEKuofsvS04JacKvsvHnyTVPpBHCr3BmNJkk20IvIaoxlli1ZZPItYCFkhYr
NB9x4iqFflKHKW6m10HhOVyYyCBNk+V+thnVwftHoJtsXusreBq1vAnAsygWQ17P
+SbR/ZUHLHyk2/dbW8RXf11WVixyJq/P8AzkbWmWjBTv11gUHo8jJuWbEhTlQRqO
cqnmeZriKLIyhU1cqgFkK5DlgkOHOAT+qiju/lTzwiqGbBSKOaVC14q5AB+8JpjC
mxjZRIT8nwTj/d9f5AoDgXuSLwEiIRxzAa6QxAwwY+J6s2PE5JJqtvcjELM+/FC/
cvFqR/ktxRYOO++Du5CR061y4KzpMLt6ZYSVCFbDS6eX1G9g62Y15EkevSS0p1Gs
JmtaJCPr49niez+k3OAA8iVwHv/1CeGlXsdqe6nDXpOaV/ZUmWiAV6u37EXHnxO7
kzDp3WdlqlaD5Am+miowWvDwKBR8O8B3Klk02FQyotN7pxL6Ad2dh7NIRQ7MQkWr
eVZZD2uA8VExvwcAbBr0QfzRNNHo83KZCINXUTfn5cqxzVZo2p0OpTyhiW1zicOJ
ir7euzWW45LUqDoczJokUaz+sg4eDUQ1BWgOUZgJ9P/CQI52aFHzRjaxROdezyTT
ToSKe5mJT2sWGrTMTguEHAo2w/bfRNcGBXqprL6TDE1JRrMtjRd4xbnDrb2tC3eJ
Vv1M7LnXih2+7LAx+t4xllJLsoi9vRQ1nIpHMlUPo89Z4EwRIwTh+w8drb/Ha6JT
suWZmpvF/cyw4puz6rBc+NFBuOxqHewHLUixlsXF+MDc7PdX+e0ej9x2PB106jYZ
mh5YMJyRhEzOLbWq/aVLymyGYwPDiaF0p0dwuR3fNGOY7vKvQlDgaTvDrdXXUwY0
5gE0S1LO1mO+pxiXOhWke/aqT8oLmf79tDHhvJaosdjNNqyWSWwv8ZhwZnoC/M1k
fZCNxVD+Ak3xNQXVCUGbXFe/96RpkP3uzBdQmM5++vccmoEVEMNjWjaLrIl41TdH
5l2UOSF3aIjWiF6vKqZj/zOpAhaXuZl7Cj8NGaf/6tNffJzksKQetTqnKvLQ9k8l
oP6aUKTnG00imN5dl4dEuapEVbUs/hdD5xPVELd8plqNY8CuKc7PPtEZ0SpGDEPn
xDdESxduaDJZM1ZHCQDFeD0pkqN87Q8E4W6A1Kzs67Fn9QZULhxA2pnjYNcEsp7Y
wFaaYusLv60gzrXUSiw/9sFMymLIZFrw0bEkEFl52crmA47L9hj+onTEKhdaPqCw
ZxP2uiT1Hhf0FEIYGMFGm2ajXAU7squqaFB/XECBCmZJr6sC6T6kciqed/JJbVvQ
KRLTrUOknpR6C7Cpead0y+x413YjE/Drl0EMEW8BU07+zQ9v8WgeMwni0A/559Ki
ZzTEOweQymc1EQ91Td4fZIuyOqXCyVfqxRnG1PBMKwmDe9+gL2x9KvgVg4btsMmu
5WlkciNjLyJpyu+GyHrut03ZnzbGC/X/Fc3c24NCYnQp3WfVeIGdlgBw4+gy9MZE
2ilB8pn1uQJ9vi4R66L1fur/S4krLI5BJ3yfG0n7VmocP2WyRZg6ZPNb2TnygIm0
MVlTxZyC+I08pnKQhmoxrWGF+q/kKVBunoXc5fTEm9VrycHoENCZmhoAu1GyyZDI
U4bQ2g+rAMLolGtiYGWwCIm/3qpHu148BTW3BxDSrdsiQF9Q/qZ7xBVl2XpZS95S
5/MnhTwdh994kvan2pkmxjAkNiqcLaQLwZKv5u31fSQTQxT9iS/oZU9lxPGJi8FT
QU0x3aS7lryCKgS0OkKp86Vt4A04HEznM6gEx56JPWUzw+FzTfNiWo3ZBCWd/OW4
0n1Dw37DhPhubn9BgfkisFb6uSWJ/k4LW9ARA21+IXse1l0ljB8lE4A2qRcb8x7P
b0hTNKRY0G6Vma1kL66rsRCqab5tobIsW7245xW6gM2G2mhSwfZ9xYuqPrGG6jJe
6w/Efin0L+InsC5CdNwbHuJtSvf1o3tM7vl2pkUcatutWbjlHhcUhnWSzgVhB0Lc
gVHAKOKBuTo8vMiCKlQKLB75mOFAjc2OG7lbsaod1TOQ20bJLhTUVe9gXV4Yj0mj
zkC9OnK18hb5Gg+RzVgraBkX/WwjZtj+sRoJHR13RZTaoeUOcTIRIYrDQHnmLzc8
EniYK/ZkSeD9d3I9aKNiFr94xenoyBQrdvhEBzbQcDqSRmv8NvlFzFu/XLqNFpCd
V6MCeuyhZpBfj4zkDWdwo6ym134Oc6v+QvQrvulTjgafiOjDduHZlMPjvFsYQGA0
7A/cadnxA+6pVvKsRC+EdgmU6JUy/ldDAVLKATGkdlj6WhYmtHVZTlSZ1Xq9wWx3
P/1wLnVZOVW5aWPw8OtbvR8TWzVlve/jzdLDQRivVMl3I0qZCPbJY3ZOwRahGt5j
BWEzPocP4M9+0ooxnhw0Iy/UtyxJZw6fpDGWIwgVyPHJLNhNSkue1B62LtDKJnLU
/tsnj05rtptkVtUd56jXYgM2CX3TE/zvbq8pRVhbo7hg21+tnPph5KaQcclqgFDY
w1WhVJQdr8AkzgT7A/d5kSGQ5SdxwB5VOc5xlEobCDysJjGgGkcJh24wNgioWTgY
q1wZDbhRUQvv8SiRejf+HgsBTXX3mUzDF65R0+/C3awX6W8HEQum6cvk4/WkCvpX
9mwfwp6s1zVql0OdmABzev0wQaOoloFoN1T1sP4VSZVpPP7g/JzKjkJw3FqKFq8w
OP3NUsfXvJW844wJFZhinm99qfoiNTpgwR6KOqz0rVWXa0kagWNF2G8aDUnZN1sw
vU7K0Zj1IIQ5NlUVG5Gee7Ha7z8fTGuchdf/e70c2jyjBJhI607bCzFZBq046+Y+
WXLDjKIdHHY1Cq4mcy4l9p16oHI+emeKbiyPzNODJLPU14MbKzTvgGZsH+5aXwB9
TfXkogUlFFtdzHAxKo4WzfQW7Y59yivk7Ko3P3z9bD5qG1GE8UDd/dxdWa/G/zIx
LYMIu8HLY3sffkcju8nB2T7eJlBkkAEd3EyW8fPFb1dCC3498ZvuIOzAoci+gFux
nW4iSm7VqdOyxNHANx2n7x+GZS5a/AXBO5+F4VjkLW+G/8BH4xyra0dIg/p9KigJ
c6wp0mf0eXEv/6sPCMtZNPMnNnHTVPzgffpyzb9/CtJ5QiO71fX0h1/5+a2ShUM6
utvC0CKjJuXrdh/j16/pbSLo7MMwkpb/M+SMa8xHeRcW8p4jcdle7gHwuB8iRuLJ
ExOlyOyNmmbEQLF6cqbHDwZXiUqBzVSTQrkpXsqQ6v7O7JMkRTQP6D+uukog5i8z
mYEhX9MnfmtKpoykrNKM78F/nnlMrrUi0CYh1WggI54xIKp8/aZm/s9SelSC3Z6+
pZOE1xE5G1MxC7dSuar6Y3IHfNND7HcI1FRT+2jFVGJ238Hne9w5oViZL3deWXaS
SWJLcU0lrDAxzuAtfSFf+F62iJr41v7o3FCyXiQEO78LIiTx7cbE+U3zNBa8HQh7
qmuyEAKhEOZyNz74GcThqJmpt8Tc5SnmiYNZwggTaniasPZin5EdVR8uRpqWeWH8
Jh/mVMBZ71L2zoT5qUENW4YXfz/W6i0sLLO2b6c8jac7OhLZOP1r+MZIR0UTTKf4
JdirzHetmkE+HIcGTnfxEmzJ4+UrPPqwb+ifi5c1k79UE9FKSsDqN5uRohmSlWqL
2x0sfFGi/b4BWSYT/kdDEqM9SzUjctQXbmcgWdHwuMs+SjJIx7mcrDfoscKY3aZ3
OOA1t0mJLbSZtrfHv5U8I5xidONLbFsOKGLcCvvf/C2kjkAbHSCdCYBe1VynNmk2
jpCeiYh/TVlaOwhVNSc+XE8NeYDA/BbowDwSNb9lnyBqNrc6ZYxFaEyQ3nk47B3U
HDr7oXJqXfNiTP+ac9+l8M5f1Y+47lQhE1vB3no5R/0re+wRKdXH5/xLZ0zcK0EU
A/XILrbjxq7rf7ow6tCiwK0e0+2lODsYo6t9LrkdHf+SpjaJQFst+G3L/Cuum4Tw
83YJ2H2UDZhmtfEH10aXMTrXJe5/ayEeuR/ajRFBpx8r9ouOCCb9RJapMcqcWLop
kqK2NDAj2U8O3Mg940GoTCBmTC/IT+xacZxKIaM34CfSmGdAMt33gOSFVJgWNwE+
+zhKs/OlMinS/FwF6etfsksomXf13j8AGi8ZLACeA80YU+Mr3NkbFMb+yRiA1LdP
TmItEjL+ANlf0ue6sH1lZx+IQNdfVuvNePsB14zltX8mZtDFuJPXchNCkNRheIvF
abnwhfiLOeckGVVmXctc4Qi5pqdWljVnGa+BP80fQ3QdGE1WwE6gB6HBTgEEp3Y/
OvGfaUXvkURt+eIBSn9+7NEISJLsonmeDC+QsIVnhJD2i5RpuRKTXmEqC+g72kb0
tPeRkm+v4EzyE0WX0BBvxejj/Mkk74XX1sNd7L5zP176ZORzIV9iC1F/0ofZtAIG
Y53/OehBKJU9TC7p62YYWpUKTw+MFADQMNRTDF2m4Z/yL7qwg6v8s375U0EuTfVg
iv4RGUA6Hy2DQEP8M3DKvJPUyjZZMDI27VB2EEJmVzlmb4boeRosGQR/yNmjqHHF
OAEgYZ2NqfnCIEDcK/RuqmkSGYDC9knL4nt0PlT4Byzg5WtZpFS4Fkws5uekRPnP
+Ijg8SFVbJj1Dhv0xNlQHhE5SjJUA11d2ae5jbSDJhAwdynMWoBpGtfss0RWrgNh
2i/j9FFEdJNNH+8dvbO+zC7o8jIyfMx92FKFyRjUV/gJFANYDUqfqQrcUh3Sj11W
uKUXA6M+f522noSu3IqNpuYvTOT/W4EOtEsqSC8e0oeAdDfzf/saTsfGusVn1WcF
Pq1BtFWwpE2hyUbBw3F3/4ybi1qUNjjUxFf9z6CYvJMKsYgJsflUfSMkdBbP9I1r
dDZzcfMlCPk5qOQCgbon+esuSUyfeVbm1Qca1BaZKU4l0809dHbvXIGfv69nVoyx
YAmzHLMOrqvouZ/09y9VQOVNRsjxda3xS/mUoqtL+5VZGoJRpSMuLJ6FtC5F+aho
74s/rvV0y6d4oT75s7HeCpMKlOBwmAb80cu68uLT0jseJCLth0WnGsV1HjAEOCJw
RCg03C7QBGdNJE802fh/forPRfYGz+YUiG78FmcZu9uYWF4eQoVPN9CmBJqjLXN1
lMNQOOUkdCv08ScYxANt1xjEQaisMer3Vbrs6Cu0f3/MA9xSVWszpFlOgU7SOaAu
/cq7S4QbSPWb3uXu5mNshuBuKa5jNqOS/2POBeDtjTP0W+rJF/Y+NaHcqeKz+lKj
9UUfYwxnJmmw2CQVLwUZklB8KJqb2BMgCOPPqH0XH65XOdS6BnRZCl6btc9+g5h2
PJiAGInCsxA5BgNxhnG7Wk4fXH4YK1XkEXQv5TZugES/vxVYjfemPd9aZaGbcO7W
iFzI2pVzdJBYXEsR8jGxbg0fzYyV4pHqE1znzjHnSBNKKI0QpzCS9pzVxCnlralj
lB2MlbP0GGHnNrEoExc594p6XlNJH2BF4B6+9l6QXBkzGx7YocWx1d5GqEpdC9l/
lkV0FNfjp6AhHZupUMPAmVLiOjoV4B3zHiKlkdEE9C3laJOXJi/hU4en9VVU8Ttd
tL2X4jj+Z90J8WE/BmyP1JvtmWrlRvLwTEj9bkSNQ74gRDD7FOWNe+ZS44ny3LTX
7QCC1VPBuzK/4NDH/QcwzxaRBloRk+lkBv4fzXKxi+F1Koehhs+oSVts1MMz2Ejr
pqKiilJxTbJJLf6/htJCsHwDmQ63I8nf7i74USbT5xbIBa/feLbRFVZ9hs/IGxPV
YH22BnSQNJWG/VJyN2AOQkoKFkeoP/GeBnxpA1cfZK5Pdu4FsC/qquMDgfioJET5
JqQ/GdNy0LAYqMwep+uHwR/l7NIYXRd7gyJfDo5OT+rttD3UaOx8dyh6e187NkhH
vgDeo0N+Pzv09cdhKQvbmawXTT+LUQXjoohbyIgPYNvrq8oG76qzX8OxoXlxP0wP
JPOcHcCcdgSrnrO40R3WAr4o2fmrOgqfKaFOfYckbm0zOUD3JkpsuVyElwmVzUd4
crwAq9bKJ8+G7LhvgoQpmMXLfD1f0EJjcMjgTArD1Rtz4G4GuH4w6KkTYLURdNlB
WijhA1vbpc8qajTMiv3GK3NYZCtoxT64aMtFeCglA5wnrcv/OEyCj6UDvajkoXuI
VLec1yGJ1fcEvJA7F3rJ3glfNOcpYqSXjrK77AEP8yFKw7+SAFEJZChsdWItpZ8G
+YH58zuY06Q9bxaMRfGx3P31Aol37SvMREprDFGqXGLSMGKQh+zbHas2/FVPNW1G
N5o6ZNz71hQ7soqiUvz4h6I3dcWfiQVL3+2+Ohc7VRLtUpNKu3B0BO5+oxmXWy64
wz+8ctj93rtdMyWuzUOjUnoOIcamgL3/XZ/7gWs7IuFiKaWlg+cXx6xwvSA3kkdb
rTTcfSPLsjFtz5QQHj21L8CyTW+RZFwB5KLCLCvAPS+B70zPO7DU+43Bdf2/XlXv
HGmy2/Z7YbIFswuvlTBYF6b5L4MU1w8StoVDiYPwMFn+r99Bacin64+TlwcEs7rG
cIR4aep9zhIZXk81nf3Ez/IY8GnzmhR9VkMMneV3IYwLVrBKePOjCSYJA5vKaGxi
frPspLV9uZjAiQAp/PF4lLiwXhDeqO1MTjE/g07J+c4B+HbGjUHBNDSWjxbDTAkw
Yk2qpab5KMKzG3fl/lzM0MB0wqcbaPP6iB3OdM0FI0rtcMaczfAv4kp3qf3nkFlj
pk1mHf2/5nMUfuAqa1qK1txq7sCXW4r+NF8YjjKXLjK7tKLpsnJN+r0CAXDRBl+0
Dh8GYjFrEJXkOex9OUYs+IhVaxGhlumLMon6SpnvQioT50iX1ccV+lsZR8bVc8eO
+oA0XFV2nwp7a8z9R15Oinif7OFcBGXLP3uy8qlWpa64ekRLR32VioB+yKWaMJ/g
z5a+L3Gf4p5oEqeQXfGmPMz6CYxAeBSLBt8hIlZfa5mjhbGMOGGXLII6XSWVQHXZ
po5uxEcy+hwB+IDVZntZK2qMgmEGxYXExoLq0hA9Kmp1qnu7ren01FzdxuaWcZgY
0mo6unmXTdeHXt3tSjmTNTeGJJrMQFrhxxfPo9H8tlaAaEwM7a8gGJtdJPm9jqr5
pYmCOZxxf2nMPAyZGMNZ1pCqmBEeCcGZwiiDRwAxmnDLk7KaRcDP3pTzv6WSUxVK
MoLqPU4m9YLorbxRG88oM4MYrHdkCAH8UWXhHxwOLAz4XoDmFApn/PrU0eDORmQz
vCZnqyI4DlJPtKazVJwoyl7vKcRtgXFpyuZ7rYneY7iPizFJ0PSCn0TB0Vm865YS
ZjUtZQTYTvsbZGruXtU+iJ0gS/NWTT5oEqHYBYW8C5mpR0p9+XwTB+Ke6gD6ue5g
hZskCuWgTCctCZnHDsG77wM+/2SjW+GQGDWoQ0xqMQBUumjS8bfRr77xRLXnr8xh
rHTeUBtLw2meBJSxpBPJ9o+AakKzuvE7GvNx7LdbysWcXj7fPeDh2/X+p6OdMLIG
3qKD3NmWfY3iMVqGtZFWVMKG6qao0v6ol+zDhCeYjEVfFEDWal9fUhV0koZgdrqw
Xaqm1QZpQe/XbuM4K9ZtKAV2pjgwcSiVhTfQJa0EZce2uKjf5yhrFuNyb11mh/fb
YmFPc8sk0oyWD0keDsM4/fxsWf2RmcTcwH2biruc/eIkUmbmAdstZs5qfRpTp/+k
GB3GNRNOOMf10Hd1j8XpdMojEQjhiVPwTV0ZKoCKXzWs2RgY0mogeJA27afzq4dC
oreumIoRt4wzR3H+s+a4063sNKpMbqhZZWNX+6YU4BZ1swSgZFNKdm0rrs0296Qr
Db43bcbtgYoWLfFRNMYc81/JHHgOcrbtAi2msSExYNhUVUclVN6q93qkl9WL2Jur
9NuZjQ9hBXmOnyutHSEdKBUmaQ1FUTmlG2CyIe6K/hKda3+1H5nWWxfQVfxqK6fY
T1oi7S80qbjfEjQ7Bt1e5X2TevVRwvAi+HHSyzvVwZysuUXOb8oBc7/YpB+uG3UX
r9e1hGZI92PY4K6Zc4zjg57vDDHv/EJinGuWf82toG12VMHp2mYEQuNd91BH8A6a
mn+qxQrQbMSUzXZpVltr48UNq8FG6VLbYsSVqk7dA4VO2Kl9SvsJDS7glQ/YSmi3
j0XWs7YOu6onOkexGW+UYxjPVzkRCS0nPSRKq6P8GtxFYdltzApZMt+VCZNieaPB
1zb82m1XQj7e0tUIV+f5P4ZMRLFOSDZMbxLgjoJ2TRIwuAQusznoDp+tPAg341Tb
NIJtG3CabU26JMRr4q5MZpV3Z5ZdyXQ/KopUpHIhSmAVIn0mel8xV0R1Gg+Xxbs0
K9Mxd2yIW5N9P55p07EcrlVqE6qPD7CNthzX6VXKZDlsqKVZD0kSvGrBYDvF/7hN
Ef6UmBTX+AR1jzUPhIojBZ2WkjiOUhj5ru01Hc4dB+S/HoH6mNzr/xSCof4tmSNg
84j3hxFDSXGqDEiV2NvVnhYg4QHtVoMrLJnYJZQTWefLg2oaa4lHMN8iqJFTomKZ
Pgrba4XxJ29NRg+AZultLTAmAsLRw518sdao6wuif5ee61t3Hhdlwqlxrn/uQvPQ
8HDpuuZuO18Y8K5Oc/8ovb7iUXaxiJ6BvD4p1qI3MEKuEBoFzlB4y7c1it4tOFK6
p6+43kI2LmMT2mD9EBrTO4m6f7hpbPN0Uws6k8rmkYF5fZP1kgKlZOAiAonpKAqP
IOZNRlw0vX/zCMInDDMMVJEnCsmeIjKeepZHTd+64p1nq5VcvqE0AZf8hzBzSFGz
oyp8QTfgqSIK+xh4XMlsEiah2IAcNgRDqLcMaGGjYG6aw0ffw0EzbrimjOrolG6s
Y5uaxouXwCl2zqhk41vbKdWkg1yfagQQKceCifM5QeZkldcogBZf9WKojJ1axAC+
IlXg8mgtaRG1U9guFxtulgpYK0wLDmla4AmZlQ8dCWe1qYDi/GogOkE2TbEY+WS6
VAgJl7NrLmd+Bf4zSRqW8wGAO1KqeiBQNg5Kv42cwadVL/w7D7pJLoQkfl6+0d1U
hV2LJ7/PZe7UaGhwu7OPzmrHif6PHe7hzae2OXWL/LW8a2gOQ7LFGv52+6AIXdUl
zPdCwMEkr3WoBCzEl1dIC6FDLbDM0HIy+oSfOkETXcIIYkFSW1BwDIlPbD//83VW
q42IQ82W4updAG1+PwoQC/+gje/6zHOWjl0joU1as+va9QzeROvvQod9AFx4KXhH
nhMrJF4rbxFGvpmiANxnrFFIgw2CHSp7dtYodqwDVpME+j88sBCpXuxtLkk4RVrO
UYzQkWjJf6xKNzvwrfUArgoZBwMD3+/sse16jgrCvni94lK6b6sn5NOm90lrgrN5
Tnb9KytnZIQqu5qf39gkwmV5R+T9283BI05gJMe8TEmMEEuWqWWrYjd2aGzADQh5
h3wzMBD5/ns/EQXHZsTbb/+cv+vWsrHVpXGl8oAI/8tepRpTm2kKhXQZrcFzdZFK
tlKIYx8lDiYNoejXyOvD8/VajvorSEh8yYWyYZ9AFVsnmPLjlfFEVanrIin8Zf/x
JIBuIrgN2VYe/gI6s0zRXCi25wgfyIIaRXKwI0WbwT3pQGl4+zWuv2HVSHSBf9KQ
8f3lFIGnCoszMFuGsX+cRbNpc4bSDjCW6KHo3J529tkdlcUbGnuwkyCXdcNYtR1K
K2Az3vRvCPGMHNkgOqzFeHk5OrShREnoEFS4wz3BEbfDlgV2y1luf6d5XUZ1KXwW
6dKXBo4A9LKHNa8WPBzjOkcvL9rkrEPwSCRo+E+zKV6Uj8Y2mTPDkR+WAvBlMQfS
RU4Cu5M6AwfpNgbYq9A+zR9ki3I5Ssv2ziwZSzZeYVhCon0qeeX/F+scAFBH9OKN
9DFTbGW609Wn070v9tAbJj0BY3XkHYv8d97SDPuIohFz5niM6shoFZvNIa7gb6Kn
05v6fTRcCC0PN4M24nm5joDonTDWqhjnVnVPBC7WKhuB2EuiWbjJrDGro20puzDz
PCMRthGQdECVk34gNXw0vgMX08QBVnL7YjC8a+36zdjABbcr4v/ih4P3CmMfmcL/
CRLkwr8fEU1ZUVPBV4VonbfzzkMe7Oa3tvqtl7+E7vnl/cKaX8seeuemKjW53WoO
07Uj/0GPU2iwuqGUVR441UgGZLUhiqEj3UYxkB1qyiaCyBYcrMfJxLZGLMXZ5mHO
Lo9n3UELRF9PlwrZRHt7zSlVfkei/Yf4lBOJKbnJsw7gqvDdn08RZKOewiYKc0PQ
tdV6CnKR7tShaS6H1YNvq65ordpxuUCeM+0l1aBhHRu6RUHfx5Ft79jWsNqs++A9
GCn0rp1ykz9eC4RUl5n4Tsgxtky9HGgudy37kvJKEqoGiMEDckRAGxM2qx2lvi5K
JmWeAlmGMt7V9hxF5evx2SFRPcL+wYq36cV6+RB1gTMKPa9wLZrwaNPTguMqepMS
GxV/K4U6DAE0e7bat9xH08Sae+1uNYxPDbiH3PRgVSbRij7tnm2IASP7QNrsFGKk
8OkP/0dVrnxxUoPhVxj1nw4/VnGp4lF2az+ryfqfGxzykZlmguAAlX3RUQVTySaT
TZGdwcbmPq7NBBSIkI0npX9n/CzqkrZ0TkDCJKJHroYsWjKvCaGXUBOs/Q0hrDYl
/UOSSL2ii64/HUpJQcglb0ro9a+USjEoWKFaobj4YKxV4o2XG/9tfAHuFBiBWEWf
tdxfsyvwXBK0Wk16qv7gNs6m5XJ1qzh7AmUN6jKnPUEJ1ufruk9P2d6cgZmnWZ57
2D4SM+ChdpVmgFU8GExEL2/uYB+Nvee6hPqre+w9K0TyHwl1+epa6wjIhN3+Vmi0
Zjm+JhQ4Y2bwRis9SNR3EU13cnc/4Jlmo+jBuNZMzbHsdzoPkT9uieHpseqCWHe1
ppWLCrXJzmDfA3H5xiFBF+ueSyv75jsOXuQSM7uYFTwdHqv4cRdusw8LLtkmYEKr
xUH7EbkTusfuCSrk3/CSHPzqQXvSRxVM3m0CFHAa4wztq9Sx9HT82DGWmz66gGTK
MlXACrDMTEACFx0zKYpMBMVb1Em4GFdxj9uF3plBQptJOuUxuRCon9RGPP2KwqZD
XMA0qZc9a9d5B2V/GfMpsXSkVfETjw0eAwOnj+UK02Q0SrUkS34zonlSb1xbTuCJ
7W5PcUiENG+kXrYInnKpnWLc31Ppv0rvrJw0hAhegCvLGOgLFkMVRIujR6U/vGRU
mbZZj5wFbnWga2AJZFFJaolqw9tSv8XwSJT7+BXJCMvfJHojL2VBxZPuA4fScFpU
z5TlXcARO1qdhmrv9RXtO/KJ76u/kfVGpytJuSy2Drjz5DFlNjE94YPdOX4Dt0Pc
hBuXxJUL9xEm/+z2Kv8UIBZaZvN2kKbXcZO++TyKPjpz4Gm2rjH5gx180AafS9Rr
abJvgvsfZKlB4k3G7M3xsdfMdKlhNGc+NTBYB6Z+r/txfj5XL7M31JfF10STcHq4
6xs8uP76UMZkj5+jLVo4XsN09YorppRCN7bUVpR9/M/ztoHYlM03WuWM1/sxf/rm
hvz7uztAwv8kAliwGs7JoMCATL38rTYSmCV7xetyCUxKt1+jC/kk1rm7FZ2VNeMV
8swkwiGKUo6V0WpNbTFyrFQ+Ea1i4SFxbla9Wtk2jlUr0mL4Wu48bQnNy5GeKyS/
7d45n33jgTz64TJvszzBm2ezB4Zo82LTMj3FrsnJy/hGllDPjn0SfkjqVS0HjJPv
hY08DIo1eTzx5J//V31mvcwRJEUiiCgxsFe/1lXSbaDTtDQr3Ht3mu6emzTiaDFH
+fENOxNMj3AdE5Lec1Tt5gXzJ+8FyErNWaIKg6Pd4p8O3vYbWMnXMoj2gO3iyAzc
4y5UPuPVOSI6D7JN9vkC6Reel4CQwp+BHjypYHwW6s7YfAY4cT+5oETkceXygrOT
aFUX819uvesZpo0niLBuAgXd3g+fplPgzeC+EuGWKYxP3G8ZxGF5Y/ZZXjm0NQRm
kCZSH3cEZiDRaYbj4t+C48ydwzhJ9qAiZ4XSNXjoRcHbGVpRUTyhI3vCtBXJHwKK
E9P2GPQpqgmzG0zJw1HcJ04BzWIY+cA1eqP4QuKpTaBUOP/5lAWy8wj50rep5LnL
xAjR/yzqCvDjEflNN4/Esl/pa3uhk4Uj8wOftA7m+bzWkY8NdSfLhw3BAr89oo+d
lbXHypexJnhm1/3imx0VlJUuk9bPDDI5ulgK+Iy94bhmt1fJfePhrZpiyUS22GHh
oSmdCtTF87Ooebv2twpmkCV9srl7k86oH0bPGNdtFTlWy18bNCG7XmTXJbwg+bCX
NC1xF8D+aaF6dreh2LgZxbxfvh24zR/pCLBMyVFsNLeJU4pOWzF40YEglgFKg5NN
viPOOx/rjhx2qdMMvUIc+gI0JZXBX4bKC9m4M/zTz+PWSpPeIdchTrNl+V3WlnDE
eD7PhCuXx/agsuFUTSzmsYOpqGIFFb0QoR+OG2X7rFTiyz0ALr5//2s0J56imApy
0QeQF9+sycVMkofOZEEpXDAl06dFbWOAldwN+ywSjwG4nLon0aLoPIsfAeNOuNqP
/GeZ9TD8F9uleYBC2VSnZtFk6yyXuEqp0aJ5cUiRfAgDOIu8Xbvi1rxho7tEhBHe
MZJxypg06bZ4g1R7s1csP6rZ30XoEKdNNss6jQfPI9ucHsQwF5J70yVduSa0zeUR
ws++864XK6DwhasfwVZVYQUOPHHrYEWX0xeFtGVxkglJrVsx9HfF1nBUFuOeE5PS
keATurbYP+KyRLe55BsYJF4SEVOajzBN7r5PxtNmMueXYUu1SQGkx0msS5bi7jpx
AbnZfgY87GdySDY0cW6WhybRugSeXHbxZHtlNVe6M7MKlSa4IEvIbv9Rh/sQtGUk
K0HSRAMWKab4ieL63TjuU9UMbHNfHl+iE/KHnhnNGOd22Pv9J9r5cvJrVHzsQySX
hIMPbwx3sw1znMcX2IQEThYITS8AyRwmi5C9kPcNkH2+Bb86U5KrQWM/EeUzCQV9
64ZsX3YH58YB3YUKmZcTFpYsg7bnpMgJtrnEP2MpsvoeVZROqPZCXYAv4OfBTgP8
MVzyedpFTXciz47iQJanTPRu0cNvKEKJf/7ppUSdlhb3o0/8s9zLNEeiKlIPnekK
sGcXj138FeRclVoOsdSMsQAb1FKgnxzFwNTasO2HEKYv+vwM2+oOdyXuiSsT59B4
63uGh26ySNGy30TukZnoejgFigaUB7GH9SFs+wmfC11hfiHuYmoj1Gq44OsnBEdp
UOtSJfgjORrvNyTIIPvaIUr7WCxUOIyukqKpLkW8FvY0XhbfC3AeWKnjCo1qn1j3
eCrBStwFXq3kLCnsZntDl0g5UCSRmCYqoFz/J4v4M1sUFnXQIgjI99i/lrPVg4/M
1kNfpvE9tL7uTBaf/DgupjIwFA/KqGJ8kD1y5mJgh6rHAVDKBKd93Fgo7x7WcXgL
pXX5lOynycnfVgAXgSs+Q1zgHEgZh6B7M4i36E9iJzvxXja+SjY3o6493ob+ID7a
5Ksir1AzVtF5jhFKa6S/UVdqlEA4oYhUnlQppFN/P6BXu0QELhRTTfEHaS3snSxA
uKF5bQNOdv/Cg4di8ZqbdGRqOxgpHGtSZgQ7zrxRl9sCEo3F8TiIhaAnMHHLOLH2
vVum4Sfj3AWTeS4DilgCBiU35DRDBq5F7Dsp6SfrferUgGQA+kbOaf8pQQmdpWC5
QNi1+OkAgiUqqnMs1lkIYYpmcU+sUe/Sszw6zJuEdxIgylYaRRh6MhMCmI8379ng
uEU3iOmlPy/dyiVh0rq6zC08jO1RU6ii3V5OZi8WEbxLir2XiPM5W3J7yBAZsMf1
I1XCEvNqGo65xqgFcE8o/bXn1QhmZlfZ9fNAPDaa3tEqAj1neS+HiMGVO34H0fXf
Va35lyH5fQHw/qx94KSvVRUGtNBhFDnPWQLdzoFHhGIMo1sR/fWEBjahHuQIIzlM
QVt6zfeOvyerwpSO4pWZDHjIKRpvekg2vzKKKeQngivL4iRjIM7ZHfHlxELWOVRG
fX72fwq0iKldoz2P10xADH8ycUaH/9i5ZCkH7guC1pgwGFgpqx1psg2oaJyu9CPJ
LxerB5Y9paLCxdoZrY2AWn4gaOZFwAOQw32AvOIMmLR9R1WCq62m4pPOKUendRSX
NPzyGsCK2L7uFSoF7+B/y63ug0P/m1/68tJwNE7lJ6JanwRkbhSsAULGnTznwlt4
y2uzdJx1zvChl/MmRcVzcSiwDFPx2sg+qYTfvXj3puMsiitlYPvb8dgqaRMdQKUk
KRaGfjj8TRiHfXAzSz+H2mv9l3tkVTHfNIK4AHSXlrOa4fBjA2hV4Q3DoNAeMPI9
ssrUjw1JwU0yZbncSryBc1K7NfZ7NDJWRwrl+T5yeKigsT9dr9YAhbKZ+Jz1lcT/
p2NVHLOSDfgPnWjASF3wjYc1BXxyW4b26Z9jlv5HhTdra4db5B5Exdc3IsHDEpny
2RXZeAS/Cx7vjspWhHYU0kuAjmlllMpKhogyN7QIUL49wVoEx4d5QCCI2Rf94dB/
arzzyghR7mLa6G2bWgd4rRGmauKIc3iRAtbBmmGwnsXZnYyOAX46V/v0OuEsHRWW
IkQFwbTSLavWukGJrtOgWW1A7Pg3V707DmjksqDpRoypvO9BNxWRBBx7pxTEyezk
v+eiJ0a2+XuLcB2h7BtyYQnwvDCecV0F3kqItcJLqFSvtS+Fs+lAmfmX0oRK06Zj
oMgxNLb3fk8bpPsAUG5e3kpqSHQZfYFn+0dZFdOIB+o/sBFiughbW1XT4VZM936d
3uiPkIuC5l4f/qeXB/1UhVthjusGpaDD1DCu7FZxbHZnhHLmL2chwinw0fy/AX36
ZAOU2NVgYsMLglRlXFULjsE1IMX4/ob6LiQj+lr6X6Gmo+99xLgfCEtl4OD9ec8V
uKXZqNY7+nyIjm7UUX9GLVTrIHxAGanJlmGP/7PLbyzIqXUTZxygoQiraMQAVd9A
VQX/3o7FWl5YHNKdWagcXuFOtStjKHht/umz5X5hXeuIjiCDJMmN7Ku4+cn8aSxQ
oEIDgemfNEVzhLpR634NKBKWJUZ5NDhyYSqgvuvbEp19X3HFpXcTISazDq7ghVFT
RaJK3E7TOp0lKmVxND+rMsFJtfxRyjSbeNtKOpSYWDBDOf/ufT7mzJSToTvfz7F2
ghdnO4DiaiydEthD28v0Mn/Vhit0BJHABr+M4es6S4PN2XowCRRJWQ394t7TJBGh
hMyB5BDXy/EooECm/w/DZhrFOIjxkHmRrMF5NKA8cbs7oiGNLLwgbuXZHuUUnrbG
EPQuZOe+JWBZcA3T/VKy++M4rU2XoYXICxGzgcva4y+hhBH7tI5Y9WYhWfsFku6b
EqtMpj1Gm8sk3NzhgDuZdNJITOJZhp8L5H9HKDWK+RMM7we1QdT1MKG7MAMzzx0g
AqGwgjZZ7s+2Uoz4Z/6ZJjYxeFV7HbZVURMazmqUN9K3vCtIRSg81iSDCxYchX+6
vi9MlnWelGKN8vTPmgn1FEwqHN9FBGVzvE9UMv3bCQdFTTd5WfDlrEVruOmG8p8P
lCJhrfoQ+PvNgRMHRtUTMMNShdMc9WPf3Eg+wgtv/Qg5FMeRK2VBdkcURW/SEHM1
F6VeMdDbVSi7zGvdrj8rXTD2wBtvp0jP84AzMTCJKCW1+b20LHjwVeN50vIjMFej
fIdYFCFq11c9p6ATTlZmNMW8hdQtq++Swx15Qvr4Rp8GiQyGOwS3lAbUgu1GX9cw
aZ7lwx8Gc24piTEoKfzhZeJ0ivoS86jFGhGH/4BBYUqPUbm5xiBiREIr/jdhaSpY
Do+ObvSHvMAyvionhOQAWLei8Gw/L6x8L62xDTovYciCH2VBdYs8eLBeGqDVlpwk
VUmDkMi7flX6rDD/2mIgGZPOg2s7Un7nCQuUYZm3AztpjO+Z62m9XX8hvEhMmnqM
s0QIbUUGUiHBqE/dbZSFYmJb8c3d3XicB2746vdea/qeYBWUf9Dr2h+18MQ610vH
1AsUzY3a0KmxsC3u81pehjaTKNQRYIecfeY+2jbaKQgqf8W5ZMCE3dg9Zy2QG4t1
fM3MVMsQ+FCmdCHjqrOiVfpFtYBPowKTi2LtLyWtu/0dMafXn4TGHx4Ag43HCDdq
faR1mMmWA+65N6zRFBDl80BNPZmajC+qA9ACpi2SR4eJDMdlh2sOJwtCQYbSsDwN
TZ4TTmzOEqLwSac0+waJW2Hmzli2kHH1CvYoOofCtN9CcYs56PRh3t36uplUPpbJ
XxoXjbTKDBMd8XcQ95rdZV6vZuSjkVt5TEUH4YIFCLIA55fVhSDaKX7McVs1n6tZ
IeD2i/H2tHyc8eO1p0A/Cq32mIEk8Mmz2W5Rh1seouip4VjXKZP1Vb3mUTHlYGeN
qpEcItjxcbHrmcKBUQYxAmk361luFGh1j9WTEZGFMp1Ao2GVmT5Xf4cSM1atie2K
wZuTqy+kTkyL+YKTechkm6vu4H7Nv+QHKO3x1dRVffi9keML5exETVMZu7xLDdhM
IWiSTj+8662allVErhShHeZTVRKgEG17acuS8WJJh3N3Xqhl58EunefaHD97pXc2
ymOvqAZ4dZY0Gm0KHuy+lcKbbHjPAEZF9otkL2nBjboTe4v/NW8eji5DApyVpFVt
rzHDQxSbAO3C3RFtwdV7Uq0nwQYKgogvRoWFADHjZvqkpXOeRgFCVIeytBPV8Gd0
zzHxp6kfCZpPrzwSBRAJ44Mzi0wF79OSAdwaKXQPiYkDhB/zS7qyOhPv1uA1iyQP
yXNgTO9/2HPA04moyDqQo11T9M73YxrXincMc+V+5tm5QVvlJ9W7PiBi49vW/ryX
ztnW5QCWJwB2k4m04cQph+Ow5SsKi0TIJgPm2WU3QBmm+gC7soyOClTWuA54Kgen
HMUJGj2odcnSAlp4aoGNTL4Pf1XJdCo/IrqoxaWGH98YNmW6pfPuLSVAa2CfxCZM
56Vx3n6nao3M9MeOm4JDpLV6cRNAcFRa7utR45uuXp9nw4MGmwi+Vig3bYB3FEQK
gk55+IKwYl7ICYZUBHBZTOIxAbcbR+bS+0RrrLVaMAKWoeCeFtEV5NAPP4/UfPhv
uAisMKCm58bDCRL3E5+wXWOXpJSfz5EbMHSlbeSw8XGdBNOQuT+mJ2uXM4UJg7DT
i34ndq9tYTDUB7zLc74hf42CPONCigG/OY8xufuBmu9YyouowFXzxfIyOxRZ71vr
a+8MxZlZqyJ5W4oXbq9YTF5cA7SG5wnHIsE6YoAebwdMoWaPq4uZ6pmlXZ3ZmA6S
bBNjrQz+V/Y1NUCO4R7BtlkFZih4lBCYYEyYPtqZeH8se7zcFkW5OG2r1wk2zBAr
A8IUkq/240w36hD9gXRyUo6N5XBdzxfNEpXvULnWUTGzjHGIC6ucBtQ93+X4QXLY
h3zyMwlIz1qJ8VhR0aejOhlbC5czU6UGfW2H/evg8wd8b6L4WqkQqhoZqX59t+Gq
gEPq41uv2oZxQ0zu77zxYsrnCcdrRHVdN+HbSNeh0ZwFBCq7oB9kxzzkGim1OcIA
H/VGtszlw/NFDYIZrFrZC4rvem4Jbqwr3glj/WaaJmvVA2qOxlKSBXVGmllICTZ9
1+F/tYW7KUA60mQnCsHsi1tHWq8/ep670Fv6p9e5fneCuBOrn0eb+1mIFULnELVT
bMSk1XxOoSXbE7hrAdlBp6cSW3/dj/y0Am/bMX0bSma4veisisnwx6oiDfa5EQ8t
nfMMvl8hW1hLBWSdu6Bc4USPsuwskkdHYT6cg2ndynAHuv5UViAczvge1MwjTYx6
wrX8GvqfWuJNXDthyY0dTXRp/3R8qQR7zLKb8qaoTw7UL34jO/9OqKDb0AYmIJj3
CMLNgAJAgpSGZUv46S2Frv3NQkRXeOltCIVMVNdPQrBcVTFiaoUvoyZj20Wi4bY6
Fc/bNVVyt29lvlBP4VG0C2Wo3p+xz76+5djCU5DoQNrhwKvTUjIrz4KRT6vfKAw4
qEgADten37qlXws13Y8L9K6jGDjSdbqM5EtCrq1ykgxnTe/HkMgHd6TeiWM3OLg5
AAykrKhwOctDH543+dIIhDG4hQoSED0MoYA9ofDOTjs3Z/7SJuuUKaR3m41/VGtM
TUfhWHA01rn7petiJMzSrW+dMiXtrMqo2z6hbsO/vMwhjuv+lu+hhKtDwhzUvWAl
wsE8/tWz8pe6Q3oeN78tXbJeFRAnXiyZKzQp9UDAasA7wVY+JjmLHJm2mbZlDA+r
z3zKImKw5ncwUAg/B3q3aD9T2b3GOMXpRzad9O5pkeH/nvwpAH2tV9lPNrAcALji
7uL/AvyvHeGW/Of86jJ7jey1+1RdJYuLztPGwxR7bbqh2kY72JHPlGoXduM6jNGz
Hr5SlJAi/4DRvDgXYj7xJQ2OfKxjhosI2fqfPBKu//sx9isauln3z/pJy7Quk7dn
UuVMRLXcTNc+o/0Jvb+zXFCvDbA6Np6pMgUwcrNR65qVuk5UDdmqQh0EvenQ6ZJL
4blpwFhjFNjZxhmahybjk/JQLJpfxb9aDiQ1NnOeFSl2EXDvRt896kwemfHdS5fd
X0eMyHugr/5mBJYVBqmPIrME3OOsoadUYDJfPx4sQNKEHxYyIX+ZUaiuQOpuM8YJ
oSQwqX1LUIXcESY02cxQbL4b4aOThbhnWv8odb+Tdo4z039cfF8HsV7e7UQLU4Ds
esbkRF+huO9yaDP4/C+Ufp+S9qp4dkdxs/cUVMvs8GfM/CwULQ+edF0tzmEXi2CC
AUdgP37ST9Xg1JihkHeIGRH9J3ivWBixPxjm0nRjQuSxYWhNZcmoUny06d/HSspY
3yGAUF5DhJgh3emW/iMh6h6wI5Fd2F88HN8ob1HU0T6yieewwFu/TVo+9dPJGP+W
mHOgjDX6zmEqbfFMCizKttQ8oKGSUY6x+35wmoFJU85B3jPa9A+VAvh/pORyitdz
Ti+WBnz3051zK4HyOrfaKxq7Noy7ttbl/VQK4nJGV9aeHWD6R8OloJsKI9WTGd7V
ES507X0WrUNVA77orpIle182NF8vAv8LxERmmG1A7+fCSI+cY9JTte3lYzVJ0+EE
NJnPuYz9f7+7kLOngqQ6PvQgybE6EtIaGP/xWWTT6PVMFGnSJ2mLTX8JsPEvxtlj
17zx68DjvBVzU2hJqkElG4CsgIJ+9W57e7kcGQ3bnm84ku23wPO4t9bsoIJAuEov
Pr25oVM4trBQme9Rawv1uCVfUvLtWKoLEqC/lhwSuL1FAo/HmSESFNd5o6twL+iF
TZnWjLzlnyWMuh/kcm8Ekw8YSwXEYalWtemBBCAAkh3mfqp4lp0oioIZbx1c4PQU
Xc9OVjOp6cSZ4T9psnHrRT8T7v6PxcDQfOMHivbUCNp34YLjLulf2a76Px0wxqWp
l2cobiwjXeRYyi1YSoqEnsMSYueB9C7zXY5UfaWU1ryUpLuxWm88FHPCTQOW6zGV
ekkoSWGcrWttH/4XdfNbzRz9/3/tylueFc473EuTg22juiMmLgdpg6zFAfJcFWxg
em/V1Lf+sp17DlYeI7vdiuXHhAWqNW3Wfh8SmQdVuQtP8f6HIY96qOhFx0upeQPn
Tvsz1scju70trXF+8T851ZMdbJ5r86RBQEv6aDb/DAsnefYFCpRklffJd6Qm+xeO
qkN+NyYrk4PgbOY4L/me5c0jQwIz6rLCrG9Wumo8d9f9yhdh6YONvHS/sEe85xsJ
fUyk+dJl3kYnqWvtluPI/5d77jp8pxJeSjaIRxYePdY+jhlMW9JZtEFYURWawsU9
ddejeSB0gL0twHwyiCFyi6zeGq7ri6BgBxC3YluYp0EZdnBrJRjOJWTgC+t0v+uK
KzwXxDMb5EG1AVUSBBbog2+up3nbmFtTWXmoWurlwEjyYXtCfzCBe1zvte/CzuiP
+sLcff9vh3ZTsCCKYGnCEfKe1TakThAixpGZPa0RhECwT86EWN2+Zdmvmdin13JB
z6+MTp+ue61z0M3xxO5J8+dM5C0pvCovtW1GiebKkCFobsFZ4xMj9SZN1bHEL/rj
v+SXGv/GjcoYcNCBRl88wDaLOeOZV4iRc9TJIbWfFZ/PwcCJhVA7feKjMsz2tih1
Kl8PRglcl/qAJzmWRsxCxiBZaXOQYx+B3915l0MUYsgFZ00HugwLvILg1P2Hqs1b
97ycMsvaTCn4Iv5+GmZXATPgUcOth8CIbj1zdot4EPiLs69sEV2Zy/QJjYxvR+s3
bpKRc7b86Rybc1H/JUxz3IAXX3gbLHRfx0HKFZOTc7RM9Vzwn42dNwvKxH+cOcc5
mvgZb4JAT3zEPgLHJYA5vefVKu9IWXtPgdT/oNAEJoqwWSQ+wl0gC2Zzan2KTl1G
wLSsoBdt/l1/uZBRAndiECbyR+XbnE9jRfFqPfSO4RWZriWYCibBsRN2MPj6QNIs
ZQ84AwoHX+Y5wAJp7x87G7Zo5QJdT/MbCjpfBKSx9by7K4Pw2lgZPlyj1mATQyDr
UuZS2I36S8KD7JPyF8yrPc/G8+Y3PcWii3BX9Ipd6Rq/WPTHM3wIRO3R0r8/4QHA
VXkiG0PcKj2FCqWTbpnHRM78pG+Gwo9wR+FJ6zfKWYu4/Mp0HNGlzD8SbQ6rWLub
+Y9DPDgPxSjiTUI/nzmX5pCWJDWYHVGcn9i5rmWnuEgRP59vxDPFqz7uz3rdIGEA
OtAcBs7pvYghAP+VAW4PWOW1fbUi2UedW5H/jENwzyVdlJ+VzLMfM1Qj8nR7RwIs
AdlVH9vhmlUPhoDjjBLVnWOjKG+tZqOMTZhRWIckNG4c9wC4+ISHfD/tGKzsGHqk
VfMen2sBzZfgKCsrBpeCVbHbnFqYgKGnUtyvRLJESq8nKZ6PeIAnkcax4Z/ZIA6S
GyT3sMBa2/ufw+On1scvsTq9G6ZJDviEKRi6wsmizCHpFXbd3BmahtGC8dGHNjQQ
QIVHyT/v36KSGb4+mx1txQhn+7C/jPbkGEQbfz+6UOIdPHaoqI+eWWZzfIH+33v8
0lzLNksbX/+X5yqtdemqU+67mw1Scdja4EzEjdOmn3ri6mp7FcQ++n9Y8hDITlj5
/uRNjA0qNNZULKO4iahAPLB1nZSq35GXoxXxJLPRa+Z5BZXVPRpHl5Nac+84vxZ6
jaexwhTXHQd2HSDssCNzbk8tGYx5EoctgE8aCDH6Cr33AWYwPNMMKsBRBgdUHMkW
qs5ZfDya9qZtGRuJ1vk6k4Q1E6qgZLN4hs/pzq4I7hTccG3E60x9MZvIKZqjoeVA
trSAERjvuWFcACoFUEQnkyqPUk7zxnHttakP2ri+P5cYebcwlr7BEthwhkVaqIrr
AccKhJtgvk9FdvZtlll0gABfC2bDktSnFCgG2DcFsuv5BeIDtvQ+qwJZztwmsHVi
JAOCx/Q6/3oELs4YZNDkwtvo9LrokFxcFg4wuMddAu0CGRpd1tedCLMLPH1fVhM8
6m2pHSjpS3j0b/F7ZOouUKd3Ek6WMGyrMsIfxecg8RPoHZXF3uLcA6QpvHQTuSGh
tcCEDxpOD0sn4UJzh99dDWoiqK4dnOAGCC6thHAEd+iQwIf0+3o2QiVGYrJngJZK
YjWIKScJLM3EiV/VFUUrmocZT5pUx/oSNC8/C9iGMNQl+hjXigKTVe5/olEeqyXS
BSrUJk82s+/ECUxesliUomb44N6r37ZCLb50GBKuSLEpYogHwpaDPRnsD4BYjRAT
nzPLsZbnuF5jZOG1hdsDOxMJg3LzjkR9Oalf/jnOGQu2IbY2X/grpLn2T/cE+9Q+
kNUh/CgQ8kAHJNvXmfiFF1aMom9bxWteqJxS0RoqM40JfqTt7H6gQIf1emK9hMdd
kEQeVmoEUcurozA0sGnmUygzRibWHbFBHnPhocv/sRHxXLvUd13BE75o8w0elbGS
ICIdtl7i9aOPSnnL2Ct1V1lmenr5KotY/i2lc34mpj3kxQtHfykyBBxold8BYE/0
o3MZ2XCLRRdPUhmHV9qZxMgqk2OlnsrGwzrGWItbS7fXN5or3dFNsY/zmePmT06j
jisJ6ipZ3XH+5J90skaVfPRsoPVHn5uCO3wmSoWbF5yqUxgyJpNtVrMNHJIqMXQt
QBCMc2Wz5l2BYBnslLZ7h70ZlDuSOxARC8u+aWUZ+c5TB6Kda9EpbOMuglOUXWpN
1PhwSJXOsccNH3bvHuLbl/BEjL94+rhH4U32qrtDPTpUDIDzHFYglXlFFQq3khHh
K7b20MW1eyogd/BC0oyxFfyV/PswfVJh8wHzl6BIXPthmtFMLmkbqSI35Qfx/Jf3
YTkm38ApLz6FqXJoegE8z8lG2VKLtFueAAQkJ2goBUEFbtTHnYFR6kw7INk7zhS1
kT2MR0FfgXG8Ks9/42ZNo43eHQDeAQGlw1At/DDm5GXPPfmWYQ22/lI3QUlXWm9a
ECq0dwXTUEOOUC+lIiOG4ByDdK099P6EhID6SQVHlReWAlrX0/GW58DEe1vefU6v
pFXY6WLGOW0owvP2X52dII6ecrTAZSewkpknQaFynFoKnY7XCYg296StVMrrmaFy
XI2KFWqYX/JLYwdIpmpcKpvvxbR3y+3sTjLexhw9nFxMefZ8hEZ8p2flhMmvJ4Pn
T50sG/DuOcX/IEDMCg0vygqvNgjkJmmUPZX3KYutLTRW5mxrpz1gtG+Ijr7GEfsb
8zrxW7EqFnS/AmIK+WSVWQok4R3nJNQZ6cTyAZmnaOlvKUAIfIkZYU4r6LbZzsSV
er9IHuNwKgfabKmpRc8bUGyshYhdJ9nV9qOPYDMwkq87wa8ckHRwa61Hj7YRiXAD
WMBMsGUzNSg8uHPprKOBidA1dUuM7qxG5614iBqATCLd+3mfIk7HEPPqfMWBr8qB
tCf4dQMrbZqlfxzhmzODV+AAql6bZS0QXmlOpBovT2BabmbHKV2JhmYrxDBa5GQH
JW1zQrVjRqgQQd8Ba0hfNsXyT6aHTj1kyo8ikLcZnF3m4PyaBHTSZkqglIGCD01d
uO94ejOezLbEIT0eWz8Miby46rfat1HNe5PL8eSGbR/Jn8rZm7HjUjnHhEQ9lJQ/
ed7dCAN6tITTbAO7p+9isrBxr8ti9jVYixhZAXIoygC72yTbFIKQtBKTvnPIspG+
Fda54vle/9Zizznk/P9jqFtQfEtf+gb8x1AWl0Vjeh9iOL0n9jl6qkDNBBf1YTTc
wAUkkj/j2CIkzVNveejQdGIs405NrV0yFGNi0RTcouJwhTFVeM2ek2LJcKxLPAwV
a/G5roYxmyiQLvmxbuQ4ar3niFI3rq3jtGKWSR3DHB4S3uLq+YqA3QR4zEQ+hJ4X
9p6WOmD0WU2JduwLa3qkg9Db+JqT1WiaRI/S5sK+kwodFmwXUxYAz51mAklm6y1z
8NPnd0+lH9XBgf1XRw40x5YapEhEOsMi8BEEUwsfZtklIO7P3tK+H0AEvfEN6dXE
3VJQSnYGhs8zdadq2JrcTKxUtzFqUWyp2F0cNACd8IcaGCY3IDXy0ViJHJJXs0Tx
FmVbpt8/YPfZWTpLRvDrfYD9Vugqam+ApaXvsbCEIibwDCuZWfxH4PPvOdgoNBXJ
6kEy6SGNB9KmDe4G7EixUVDZwB8BXFAdPfmuvLGQiVSXwtZhflj+hUYZeIZE4txl
XfvQPord/ug9zqgzDPHnoeGllIy5COe37+4NlhAzoXn5NsmbGV5qRKkS4Riq4Gy+
3zLcaFYDBwlVs5cBJk9JcyCTd7zcRkNq64ZoB83u0GEWcynfxqoQ4TbI3So8iqE+
iQjVkrvAnQqonYpRLNMnwCMzoL9Ze96r8v4qpceYiUw4gT1/zKFQ5dtak/zFwIcz
jGGtAvF4obhsQGVsdnTMtlw18Bw3RMJrs2zIHdW57NTFaWQnqOuxElx1fPQRfkm0
9I8NWeM6/DMk1uLrxSZ22F5xbhMc7zDuSQLMvwY6ZV6wSvxeiwWSEcX2P8Ki85F5
JY51K5NFRh0OcU2zGfUpuzeoAQhxdbEZy2pDNXk2R6YXvzg4ylJo62FGHqIwS3Ss
mfP359DSg3lQ2j4XBFuhP4T9GOwBgg2NWuuEvnEgALmXWRTk5228uF0i5L74DQyS
iB5wIFJXH6MyLEhqi08mSX2jsTGymCAAtS4Wr0V26SQyueHidSfATL4rtMqvOz/g
PnwJwE+Dy/T5GUbQ+BfX42UB8g3s8RytnQelpLaNVOdndJgC7OK35WcHmhzDpSPw
4JrxbbxuyqCYBUS0C/JdNMSmw3Aqlz1SehBIDAEEYURPujJz47QJhyCXdzno9maF
n7jDNeKEt06iwVvv1cbXki4UuQX2MUojOjCNzotS7w5uR5dkfC1KLZHmYbU3a/aA
SzY4XDAxDJF+0wW9faeYmKTCNeaSHs/YRHqHm5p7Lx6vIMxLoWQaxwpSChMVCCqW
/6XtNtyoKtFhqAdfpQ6XWuvzFpxmv2r/EEHElyI1mU8cg3FDA0z3PQMD7wZVd6OG
SLJodK/Cs1tRUmIzS+rM5P0W4O/kl/kc0gsTJrvpYaBnjoMf5MeRMYpmTJDn7ybq
8XXxdCEsDcLTn7vLVOSf+7w6Rfjn/Gssv3W+NUwoGJt/u92HQlCiPZkmECHpM6Y1
QgG4DfDBT6qLvIX96DcbDyTb4YTnPFe26l3JknB7IzJNM4obZxOaHOluPw5RR+KO
dmiZ7PT6fJRqVoz5qFcLCv0cbDrSwKTMLRCqp0NXm54g+/eCguKHo9+RVpdc66l+
D046I9tpeD2KhPssLipBWOFseUu5ssFBy8ZIrJ2wpoRnwOXglgFV8rCOx28SoogU
DJV/sAPfan8Cyy3+qifBV32VXGeO+Zo2885jtgmYnG2jOziDPISXaHyF++/5P5Jn
+UoCNkD41j7JErn4Ql6vf9ZKYWDHICgAVO4eIZbrueSkt6tV+Ze+h25LiO5mRqfR
dvVsIqpXkZUTjDOejNqC6KpkBKrJTZHMWB5VDSt5kypzOjbuS7y9ADyuDp/cPxnx
dnBZPFFVZLimQ4lkjNIzkcjgrs98puanO6RfaBtXgcC1MH7XjScdNXUdifIsjgxo
530DLhb6ZYIEH8RG/imQRbzdaixhvdmNkG3UdNyFAulFIbw18P6z6O1UnDyvy5ZV
RUUWoYdYqUZghmy6QrFzv+saBg1+Wb1OiHLZSeymJuKz7pIeCFHftvHG39r1hmCG
VmH5dlqmRRsAJFmPZn//TgNyuzsz4jfFALYLwyfzvukSoYrw7DmAts9vt1upXuJy
MoBD0IXW2MTvqaDyuVm1mlOaf+8uMs9g6N0mWNuTMGeraDUkWKKKLtlGHDFxf7wg
DJB4kFl9+ZJMohwKALtWSTbvzqlcumWpeD8xrgeVOpR5B8WWX7tT/uTo4hvLRwt9
LAALS7vIZymuTj2cdjvxQd3GBv4LZlJKVxybMLlaTDqJfvAVJUJGGGdDzAtqjMEq
xcquYL7jREExXPNEOXZuyNlKPxDF2SnemAll33Tjy2UVON/Gg9LHOT//zhAOfC+D
p3iyUSIYuRQqD6Tv7gVLGaQj9kox9IjtY+Z8Z8a/A03wJ8d9n74c6o9xXNpm13MM
I6TmvIzU0jVt+C9n4zazR8Z93gZzG3gwX1iFitAIGIHo7GVMufK7H0+yalVyYihy
T5Oyv3zQMdEX6gIJTXXkRrBhOv6gIPomHqpgXtbARblAB1WSGPhILS+pgLI7Uz4z
CvknjKLyN5fwiWCfX+gcm7WXRglydA2t1b9IrIxXWIPmymF8FwoXE+fTdR2cDX7Q
TYVLOWo98Sg73F1wKxZPiceE+R0jMj+OFTt4g3TAyh9YoQI75LKbX5BMKkx2fefs
JsPyoAcJUikT0x+DimAyw1578ry/gquxaQBTHkUygbFQLVpkerFK48GZ7PiJVcRT
mJ5rT0RNiMZGx+5jj3QRdYUYMgHChMj3Y8eFeCMVMOUHl8e/Gfufzotvj826QK/n
atoAEYm5YUmkOeVz+WUiqooLbNsHExgKBiXFILFGMSW78rdU2B7IDNp8L/MiALhl
nMBY6TFPK5ghYr24eY/wgOW8uBQUEC3g5Iw435z9FRAD84K/zxyMzi3+Ml3tcd11
gFLlr2scQlivtt/HQRofUkTeG45mBL4xQUN/GOg1JJdxli9/OsmqXaNy8rwsgFol
xCYGxezn4g7KTx18lKJSnMudg1+V2lGqAw5n5hEx9PoJNvq/xheAd2F0rmI3ZyD6
jRtjVFPUN06eo7scKJt6rYRVFVkFB1MakY82DBkaeXOZ0BF8CAgG0QXTMcfBu+dA
RYdCXyAURQx9IhWsxnokmmlPE2LAX8Gw4QC3uIGVOMjc1PbMuBR7c6ALxBjGt1W8
xCtjIwSVkHcnrg3j1RBOkq9ybBsgxuCt0g2hm3b56skgmjaOUzaH5+GvIKV9yUYm
pN4M7gr0sgcjCF6TA7LFoTVJCi2sYDPQ5JGBiroXI2Qwx2MFj07MvZigc3zV10Ue
ziNR/tkZ29HwtnBpHYLTxoeE7L5fwJ8xC/Fp6ljMdVrcPftNH6pt+liZmdR29/1C
spU0wMSaGuFkxiTp1NJ3xsVu1+pqq022I5tDUm44BnBX6VBB5xncRK8Dii4CBXpy
mVPocqdvRbvYQxeIG380OPTCbzGmW2w8E4C9ZUxkl8t2tQ1umvOSkMk+gZ/SjIQC
iOzIAS5/OwIaAS05DT1nToEGUj7WWbxuxx9qEng4yS+uVHPVZkqzYWcqiCXN+Zup
iHokGft0cSCYwlnar8qftlSPaWFNjxLsPw3UbYqmU9SWjVdqBbkVtgaCApNJLKKS
C7lZo3+mCgNFw+/EpHbCKFcl3fL/Sj3UQdWoaB10mZqm9rdGxaChPx9nUwRFDYKV
UOmcSYCFyzjMR51GEjQ9R4bZvZYes7GiyOm9ERSuBCVZgv74gUh+tGxWGAH2n48l
gdrBKV0I5hz+lsnj+HpJ/XqW5sqgaAzXtECz+9Z7gL+GVMCqFL1E6B+jQAQWiI4l
UHB1Q/49OdooAHX9Z13Xct4sDbhv3lcCWEePn/4juGFvuqWgnFDfoZOx/7ZJDjmH
exHhtsrNbb+R8AiG/iTQ5qrrqVcf3ELomXe+hJDPYuq+9LIuQOp5WIwZq0P/h/HI
GZCSQRGhhTqWIcbxiZ2c8rUfU+RFkYsGnr3I1THKrZxtaiYCbLO1jXBW/Meo7T13
9PZVjJ4gETJmD5jk++9DH7d6BIysYfQcVlQdmIvBgYXzU4aNKXs/+wwfLBTqUuAi
265POQH5XI6Xysse29HfIEQ6VRiCA8/gpGMR3a/S9o5MrlGn1mkYfUCgZFPc2DBl
rO8zDD3gNcSpYKeBkXZI3svgS07krMPpPx7YvFYl86Q5h3KppWH7MhwOQ7beEo6a
gXWxjnG1EfrtNnbq/VI1C5ZCCnrycW8Vnj+r/bn5Br1J/qXRNP4z5YnFbl3qx5L3
AZfkfVwOg3eZvEiVrZFmYxtArBqP0vejnRWrs0m1dgZ9xxASEFhVqZuY4+QRx+lX
Lk6aXz9JJXbZbK0+AG+R7h5j8sRNdswjG1UOCm+fZuFo2q34XoywUY1Taa9OrUf7
x772R3Vaipdh5LobS16aEF3woS+SPc3Hc9SCBBwtzGcXCfKNW3wl0x+1YTKxjo4f
ddCi5XTjOwJe3XTd2Ucw7wYRBRbAf5iVs8vW47tYhOXeh7iUowreAGm2ODq4xiQ1
S/Zqekt2Sj2rAtEPCKTkfyFWYhb2xw0YFgeWTKNEzQc59xHcJGIO4G2VY34yUeMi
+FO4H4Fa/RCWJTkPAlRp3DJ0UuuWugm59uFii3ay5OITvBtBzCv1FmWF7UVNEv9h
VjWGBvjAMEHuy473tvwGutU4cmUwWpfxPbWHp+PthLzFW3qvbWT454mGDkd4OfgQ
PLV9odVzLQA2nu41gkHDB+DAopeX7IVhQhunseUwfoYdIdMj820zSBcF6/G0dRtj
iDaMdE7ph94jrCYBBs3ijqgO0ezauuAc0+arezgjBErsicT27D3a/xmtZfWcS/1T
ktKWfRr1X1sQECMd++/iTXvuXqlhWx79QUcmhRbGD/480SEXTv95CszZyzl4sIx1
O9um58XgQd2/f3GchwT5YDzck0T053o5/oOc27tGVspnqvfdkFRMBlEg+nuOXUWB
jGF9DsGbrcv4IppxBEU8U+k/kJiupLFnR7BXi6Apy7+vBEtd1IVVQ6l31yHt6eTj
i7mSFqWZK7n9ayRNfj1WcTEOeQgZoMKIn1vbpAzgtt5P9wltaZcdN5D3Un2laDZ7
PC3a8G3TCKygUDbv2M+wgx/+dYyXQZzEYpLDugbbeSi45B/4cJQAjE3n4ao/vExE
b6WygfJFohCqf0fa8Lg8VMPveoYXgfMn5f0jCqw7gcUpqx3DVC9pZvYYta43btzQ
Qjs7HldanRTs6Kgr8Iy1ZXWy8aRUVSAxtblLHUc6YVX11rUUzWACetlKNkmzgeWx
FA0z649yKsulg+umbhZ7KilhGR3iXTuhYTjOMO4G+Lo6J9aGHOnfrO7OgZFnC/Q6
wJ89mbuWPVfk+OQmvETy2zzXIznhFuviIJpk4CWYZnr9Xj6wmzU1asZCOaA4VBs0
Sspam/AzCd8nMd48uccmPilt95oqJ5/zhqv7GFgU8RNLr8IKa7jTVzpMEcCibXbg
tfbMFKtg38VP2D3zO6LxrlSrDE6xq5n+O1w2R7BDUVCgsttTJjPDry3ETgRsLghN
jpLGhIvQsSc2QszfGD/s6/UOdGLlBLdTz2kmaJgGTfdU05jGl1FPQJiD8Ju3zPBT
T+i+D+61HWieugA+sf/TxsC0bKOTMMhCZjTjJPjInAVOLTM2p/Yh3xwobCHbpTbl
glU5IY9lYYSN3JNjZW2ReuqFPGHiU1f8vMWtCyXl8GKX8VLlAu0y+7FCO6dN4esI
JXJbJ0XGpA16C4k/q9H/1H2suhfHxdVNDM68dcJ02h1ysTueyelYiIfEe8F6iBMN
6kpWh8/3Pd1bqXbVaISYPGNvjw5r389jLecJr2v0/qj1IFCVP/PR6jtlx3exxsAJ
rJwGg66JB+IbwrV5tVf+1zi3kcTYYjN5k+4IykXGHzPnrQcf1yoNk7K9xeg9hOz0
btVVZGLzo48aG7vmOJcSvvprbwzwLmOUHkDrxASyvTpgl/E7CZERgNFvRcHUCFgd
6GeJKlkHYDyAUJN+vDjnWLHfnQNPxA0i5dUZBOCflEoiPVFd03ROMqVEDy2DxDGt
zaMaW9/aO5EZnmkC7ndRFEmgTZYV8rQ6wr2UMngjCYyuTszoeT0LJ8I7xQIpLq0m
UW3MxNhBE0rqG47R9WbISbKV87DPbb+AHe/oeZUOy204FLL8VjsGRq8ZxLWsY+Qm
uI/h6ReXOUwZhe4U86E+hVZWInHy06PCpuuRy08m4QiddPXEwj9N6sWlR4UgbP/4
2nujKDR840qn7GNe6ayuEtPF+Lyf9ctzLUQk27hGri+FM4S8VbUOgWeH9iqpPkmK
HjYXhi9+zMn1yUawqeFrp7j848GYewUmIqjvciz4yzl+cf9Awvm7tNVJhOwKSJ5h
RYQaCm5HKXdPSZoJ0PMQQFf51Th9t86c1DmOoknyBsZqEv1Rp6FXlSNf+mfmfrMI
0M/E3TAJtOiyEZmu2S+cetafjiBp8LOH/5l6QORJC8DuniiLgy413zeihlz2SFVd
ph+tkCsk4Ts2X1DO5ka73Phkmg5CQl4LqD4ak4hAxDRSobFyb5cX+vpUBOAKiof5
8ldR2mEhujxzKcIxteUT2xkO9KI2GvF4Fwt8eShreK5ezcZ+HlwHitXpBdajcDlD
R5IspXgDF7L32HjkNjjbpX/0Ek9DDSERC4uLbhbTIB7FwWNdg9TIYIqDQz9j23hn
0sMU/BpImPiV6U8UpbQYy1slgVbqyG678oqRPOjInwQ/C7UDOk6cM5XnjrADGWLA
m9MK5pPnvcPilSoJo4Cj3ze0fptdjQHZYyKiWCAzaH52BYC18ZLSRJfilqgYT/PN
DbcR2XmJaSAlKMHVYRHqzNE7eqd8INSN31ugYICN/lgUSe1MGaacErSshfbZJKt6
TomlJmxhDsyhsRSCetWD9I9iogLFRgZTdBd36P7oD6gSbYNNUEx8g3stNindsWkJ
98cH5B+W4XWpYlKozoTUZBN8RIduuOYQ5eTFWwPLiarbwAd3qIHJls2D/JgI/QAM
UPqydBr3Ruefc7NtCaUNOPc3F/yjM3Ga/NePTyisJ5DRPnlrwtSJpNVlIe30T4bB
Ekz8UyhDQr1QmOsqaBEPF0TuG16kr3Qy7mg4SL8Bu9QtMfBkjkPPhubhTE6Id7G0
8873vCNR+XCaXulNqLkOmmfStz/o7Pg1553gJ1vT9IRvPtpUQERFs3uJxipsH6O2
7ssRu71V+4euMQAxnTX18MQOEY+R4y503iYPuh4K4Watdtt6aXisBq2kVzWkqcZA
mV388U505/oHIuIUNoRHAzV+WeaZSlUBFU/Oq7TV73WCveOCMaMoEH120KVg+UMD
6l+WLsiZSE2FQZSJ1xnlPdRv4Nj1tFZZ3O1Fukhi/yyLt+meI74F+0qKIrhbr247
IOLEDUQifuVDfgsF9HJOPyvCiwMg+xwQshc/H7ojg+m7kZRmdfFTJJmz4E5/WjMn
p5ABjmI4v++aLhCd0eUHYccv4VBbO9Ogy+LfWSEXW2sOPYneiI3OxsW0RLohYk0S
IHeNk8wpdzufEjb/N/+s02SFMy5AYq+lVLD/EXvFu2uVGn3KMameZ/FoFy+2IYMn
UzajS/he68gSj2GI/5Dcia+eTalmobcRKZKvHNqDIiU+WrdSx+RkccIVUPI9oKu9
V9UcLv80TdBBOw3Gw4F7ZKAVO+uA8/fg/nM/GazkuuPzY6F8y9O0IVdPoHCgwdM1
kZffsVluByFLjHIMmqNg0mYM98k3bOAjwj3vDfY4qB+4K3OSzbtoKEZ5ygOMm3MI
/zQQSVqwZs3eKeVMAj6UFNM96KNPqQdgEV9x848+KH5haKumPQelaS1nfKA/+qtN
WNa4lPLpWjCIDmKOviIt6f1IN5EXjiw9TQPhpxIP5SKgzFyx+o+1jxdzjauZMUfk
vpwEe6FtSPVhGqWpCJD3Pvk/8JBxzjyLb5DrkdXBVoQzp6iaS3vlCTScOVwryShp
IwVgUZ9KjCJzAjjcaoRuD2O+vAPKfzpcfo12Qbn0QQicY7NFQcbLmPBirPUWedYY
UOd3qix8FC2vRYd4KWm6J6EZvcBkqGbCHZUYYjZdozEfKS/v3Te20v7adxeGR7CC
Y+z25SLim/UQia7wcGjs0svS9b5ua6wxm/qLvETEFrKImvcYSOfgKkeis35Jg6Zv
6m+uzTrljOWgvBI7X2jUBYOvIvU1tGNwqmm3O2H4iMWHOeLdh+bN8P52l1ug9Iep
w2xVkwHbR0x0GCBmSj057JUYvwKXifX6rQVsyhsycRddlsLYEb7scohiHshws8rX
qVR1zFLoyeYm5bPhrgIORjFSu99VErQJIylpjCTzL9jWSMWhD/79V4rNvy9VkB46
LQEsizLC+NzevUN6PpgxCINRHg4waivsKUGzzLAn5bJtm7AyeQeTGrD2/vnE1Cmz
gdzh4o6lCm7Ork1dfeKYDtfvaTCvWh1/cSZlBjXnpZyKXvfcs6V/g/EAAz0gu8Xs
2g6fiNLTAWzPTG9SrY9SPW8H39x2DIDjKd5j1UyugV+UugPlrLAzOr3vetFKSf/t
zhBZS2ebPWFGFMQNY5ljiQKkHMHboW0JHYytVmkjcpItCfS8qhUt37+j4acvL92h
byQycEEQ2cRpyOyjwnCz4FelGiAOQ+A0l5CHFtYCvHw5rKvs5k1t160oYpL3ZQ6d
K4l2rri744myRIduyuRLafOL96JbwHTf6VXlwvruGvQMTkP8x7FzDOU7xfGvbWzF
HgNdAEz/4SY2DZdJkvz3SQpFET4n9s/mKqHz1chjRtzyNWH+jy63JsOMNDnR30ta
v2lOMO0SPg+gc2bVhLTGu6ZJ26rTpMSPm5RLeIAFJ7nazMHd0TPQhNVf0/5LWrGw
4vDPwID8BEfQLKLCKRA6IHIGaa7ZnDluGZKT6RwIdux93Pq+Flw8eZj/s4Y2mBBx
S9dSsA8se3aKOTXWjQEVfF5AMhbnk9RR9xV01xzsghSn0Kx8fBEt6gz40SXGe4qi
mEayMg5kracOHeUxCZ+s1uA7DXtB+DpKjOlYUw24TiOgkGBx7soWQ2/07PvvpJf1
9YzMCL+FRlaaZTqW5UVKE/75odGJDTg+u3+Y8tVn2UAPpqxKRIkGMaMzdXx+Cdij
Dwrr2pZv9po7/b/CLc5MhsU+CHv8rNcLqdLypufVRXhz23cV8Mu3BYaK6NkLWMjC
tggz+LHGaUSxl55MTuky6MW18GIwqCFJl9xfbTeUU165n1b3Umr+/OExLdH9GVfp
sMh1VZnrPpIQbAZIN8oE1Ty6mRSsTQT25xKzozkViwf3jglxF5lls9NPjPq016+e
2lTfI+euTnvFAkEGI7yYiwpUOykeSktLJXib6MVH3+CDPT0BkqVOWIptkEi2mWOk
t6f6tB+6zi6vLKF1qAv3Sqj39gaE08MzUqI1VAOX/EpgQdEvzdNMuTjkBCS5gM0o
yWUfE9z5bf/8W5k+wpHchLEx91Ei6tFqLsTDD9xjMbmWjbGD636tL30IEVW9ZX3d
09uoB1s1tuhWG5b8nZFlFxYP8+ZbkoKLr8J7TkxkG/KAYxpujg9+jUcPdz1cVUtc
7Q0zikWPRLD1jGuVSoYu/nGEpzgI+3JJld+4c2IOjLKETgdmOuwT3EmI/o4RyqfU
bi5t3s4FjxDYeVz+CpE18Yt1aa2Jk0nH1affuZdxHm7Z09q+eEQhQAOlDiRDtpbL
eomDZapviOxxSkOTQwwASJZfRRE0StlOra+di0/+MgLu1YKjgLM1/leRUba8HyoO
cMxr+Cuy5hGHLTkZxw7thc062Eq+rI5VmE0t56KlYaN/4TWJ1CEsUnjwqh8YCMtm
82Ff6o4hM/L8gIKrrT9GUfhnG7GxIHOuyXHOW/KRn16zvGXnG7Z6VZi57n1y4O5z
b1u3Q96QillpH5zCdEQM8BIfl1Q+58IKdVlGvP0VMwvx/X858uOVZ20HiHMLsGmY
Ayf9lt3xF4/fqYXx3toglAVc56VJRyKjsexe/KRR8Ra3vAzTHz7EvkYHe8z/QhO+
NLeGOD3VGD2GRxBG4wqu6nz5u3cvc2+wuM+4FreddNfhxDGWYa4Heq+q4TVeygQ3
eKXX1+I2Hp55hgqVSA5VbyZPt87TgtUxyXiecWYjtTnT/Jo9nz/QJGU2s9CIlZ0l
JwphBsk3wXy2M1QC+5e2hy/EeXVYhrrfLJzPNNeeFi4R/LA/QmL1cHZx9Qc6lQSs
rQ/fWSPuglEWDDHVDlxKQq5Yur/Z8Wm6BgFmHm8M30HdmvujTdEaJw60lHd8fLsi
o1NngumFXWlW8CO28xwwIoP4fOSlGM8MCBSeuBJyBSn4pT/rrhwzCldc9y3R44g2
agAGMBNP3nr9IzB+UywTHRAzz3OFEziH+pTfVCbljkewBh37mgWqIz+2rypoJF6a
01ZQwL0i/6AuIPyKg0gvjZ31FImGVd2o2ALawhH6r4tkPangM+gJLXCNeduRZZ9l
OJrl/YY7LGW+RBuY7+ih9vuvoQVQs1gb0UNTti6/D1wBGDH0PuUXRnVvXBI987rT
qo9lxSBTKT40PQSV5/c5TY4DCyA6++h8lkGvls8NtvfEBa/YVG2XbF6pCb1a6Rh9
JzzabSdLnIkSixf9DdxxtqQaKEn1IxWYuGOr6bcAQrucmYWRQpXyCWKE02Ti6t8s
Dl9whZ+goB41Ah7Vm6iThuyR2uCqtS2PlyS0iZKBO4olCQ1baD+ndbkLEU7OBErX
ky0gWPZRvKd9YGlMCDgG7ihtCOgY6B3bFhb1Ea3ZLXeGFA5DVqke1bw+knhqtiBA
pNZNFExeA/e58MdH7gOH4A/8a6n/e5kg2VaNG3S80EgL4I3EKCC201IxybaA3HT3
IMTCcWu/JCtz0JLvNW/To7vtizPITU3ic79mg73OI8NzTHB85X5CkKDtD/bC2jTc
tDALfZVOApo5fp4JcNiA9L7lzTy1OGUaOJid0DmfLXHNgSlgcUActQWstc2NWhVV
FlUbl7Cz8rRGGqu/R4DdIDKV/c5rfe76UC2dtpXFLZOHeh/e96/VXRixsTAlBGhM
aUs4wmyXq/P+glIfgDbLEFAPcGr+uVb9ktBXz4KDEajPrwqmTKQTRM/JVo25qeIC
EmdJx34H34s3bAN9c1zZZIUpEAwa/cqR+DjTBjnHvcrDs5Thre4rDZL4xI9i1suP
X7EY1YyuT6drYj2OhOq2TyVKh/1ojG3k9j4et0xe8L90R3Pyvb81+nXr5z2kR3JH
wBqtillOxBj2QIRmq+IREdStvTn6iiwYpfdWpUPlvBUITW48FPePv5ip8e6GA9iu
Eo9FYXAUIPctOlOm5BIW1c0sa3zeqLXFrFoke7SNpbGfuT0w/jtxYLDR1T9JH57T
6L6KDH5GoOx51Ama3eXTnbqUJIQgQ/0+20WvIg9DFpj2uVijjCNaPJbgkJ7urMKF
WmT13IirkAwNeXf5a3aXas5lQfMh+252w9KyJo0PuagmXZg4ZtKJ4tbQh4o2HsZP
7Ci/JNGqFhOjRD8cHua0okiFdX0heyhWIuEmX0C2nnAX4yfAGkCzTuLiowyp78aZ
ZcdigJJeSGWmHyVbIA7g+9k2vIDGnAka9lR1OmYAFCbYVyVUkzP1arNSm5ZTaYyz
zkKIVmfdTF+pCth5vpXGxjgiND6uHL0WTnrBjWnk3mIWpr3c165K130Yv4WV8DJu
a+Ewds3VLqIhRMbpabzKTiYYGqfIP5hzDQFS/RtAZXgf8nmvU6y/Le7H5fK6uwxY
eKiF3+aTNdrEiP5BJxpQ8bWneaHAluozey/knV9hiB4Ejwzk0MjQe4gteB+9MdcC
wOVrxxStK875NbIkmMDA1hLJFfhXWIUAateOALDh5A1HHrNrQUYkxf3rGIXfmIi+
fQBW75p2cf5I+jwS3xDZgSxZDtG7WKuOjnSuA30e3D8iQyP7z4bYsNyjfshHei4J
jMiiwm7de4nkgGr2WhekMeDW3TG6r4atbw9ExmBstvsqBo/ct1KUptlMuzNkhUrW
f54S+xyQsYVLEXf/Z847bTSRQFaH402eO7L9pSt5kCfq2eHd4RxQANxNQfkxNDa1
RWFXKbXuiE0jknC1YWlKXIssC593yP4SLvROQmsIep75gQd/xqgh7G9NtbDr/raY
mfZNgsgnajU3JYgWb96PL8KXyhVtbpATUt5GI5SIRK2JSQ4eegOoDfRK5ZP8ox/t
oLs0STX7ideGJAsMCZArN4mZ31ikLZAdhfdgP3Oj5nBQDv5XQytab3YYI6RyOkif
1jiMR82X3ab4O+AVz8XVU6KAo/47R8SRL6lPfxOPUHW/WU9YZETTYA+4AVKnUeJH
A03OYzP9TCSZUmg0qRixRFHVMy3xM29OgIc9PPZr4ZS0N9mquH9N/7YCRSvKHise
M0dNDcVGEvnBQ1jNLFuKU7gpJ+uWHAtpexkRdreO+vgf9EWr8X+74Oo9tvJPTa9R
XKRK7VzWdQt0YX3HaAxe/CNiFMiUUc9u+IOzFbCtFjShNbBbx0luCIorztGOBxFW
UT9AfhdSVawBu+WEhyqL4ngVxDi9AsEiNLtwo01xI3lQVZl5skJhRtIDaKFVU/rk
Eu7/ODaOQvn0v6SSyR11XCrczQBq/TgIlCXUOCXH6dxrFwkiGKG/McufCV+u3ngY
f1uhXnOQ+5GxhA9bBhv/mleRV/XSEAu3tNCkIT1lMCz5nE7W8IHFKy3cjaKTdZOR
tb7HRGbrc41k/U+uCmKWCgckS5DZt88vvA7PFKwz1nxJ7RaiU28OVll+LPYp4qYi
rI8AmjTQi6oAyotL68oQrxhMM4jODu2Kd5fiH7OuhLJbtGueSQaxaaGT6vGAGvNT
Dc6KkCQHNBPGkzpOZRcfXSYNqPJxl0JdRbSCZbGgEUVyXJY2uAEsbhynxpg4cDv3
l9Iwop6UXeBV87wMb+AUohFRoUsiZVC4KsiC74jFCfpIfsYQSRqYswmv7xw47Vh/
3dMVdi8eox2vt34uVLYMH9ARMebT5qqqnJouFz+TtIUt67mHY+O+xfpn8F3bzt9b
OwuXoBmKft8/0MDz0kBboMZirGipcgTo9pAplDjLIlTxpc7Crw5sMmJUiuMNYnHA
qiw6tq8j4o1Vb8Gr4uCSgBpKVcCZTb0ZUHuvzB7ecdI+4P6+dRkDkDhEKmyeVKuT
SVdcqobgaKxHtpH890IyXtO1vEknN/RiWXKCuvx8xY4pkUBVNSLHYWaLhrUj13R5
GGTu7DXaie7/SgJ7LJwbdzGU85LOZvmJRqI/on2wNrOTeWBBlMzU6fp6SrWWDODL
U6wrxh+lbFcpfIJoh+ByEysxE2pWhA+o2HBvwME+SNIm608iTzox/qHmGKomtxIw
80RDXbHuJ2RnU4mYHj1wQnvSZfbTQm2OgMIv6uCFVpTGUFc/U4E5jsUADpzidIXV
vAXVJdTfyUiWDq/4cf8qlCAGRx9Po5cNn8GRoQAzdcLHxLfOWnDkmrC7oV0PAxe8
JcoSgiBcAV658gyWLyxZduwVopPWBQkFpvLfFBxGRxmA5vlgh2ktyG7oC8HseUjG
Qtym8HiLXCUOxu6R2IRtw/7Srr8VUpaLOsCuBqdvfOh7KNuamByShBCbSeBp5tRD
kt1EuoHol9pt/oeC7VMyqlCeJPD8asxQHkbiuuBoOXa2zitlvT+sZq30m1N8lROl
DnHhXmc130Dv+LhozKtnTaH1pZPTA3Fms5CqYxNH5gkWa4yGVsl3+gQf72a0f0se
+GBaRT0r2C1+VmU8KqCVxcQzSufnehe8I1CQRnmvbjqRluYnWxck+MNXZQhj4XaP
iQJ2AfdACT4uDJQrKLBLMy0J5XQvO4uLXyOIPuRleTE3HBwrQ9Kqn7FfIM2WNJBz
i41sWvNw453adfHaAHRkiQcPV1jPS3mbQoyCg1hr7229xq5OaRR34LDb9GDRHxIZ
AfAbbm2THSEI3OGLVriz9CRIaD8IjFGZA8gf2LWPNBiluLSjCUH+FuWSgjsjieat
TlZBKSKm+zTct/wq1Zjtli8M3IkuEzN/HJgGADhdAwjJZxjnPLVkulwGHG1hHHjS
C/03olpBpiCruL4erUIXmKoSiOhNwwNTG9/kPjhytjmMiPN0MWidwxoADkpzD1GB
mhck5KdhwtIsAv3JBDeE0JFP8SxX8W6m7R44PkLa+QrKYpMleRLNxUEZYaFERzUt
sjkqdkajLa9owLuJUahugDMFMZ0qtQj2LFz0OLsCPyYFEbpYiWdE0zXU6GeRW/1k
Lnu/YUTpyT4HBHM0cA3kLOGsHbnkq3EVenFWMRW8Oe0f0nFu4AHU/43MjAVETBya
ZjyRacDprm2e08pDC+Mi4JALeuGdsTRa2OKjL2SlU7jBc143gUC5WEdyqm075ALD
tD7uae6BcD5mURqitGNecRNSOX6xjnKBws+blVqptQMS2cRVr57XzN/Fyq6HycLi
OAyn9Y7GV4IMajlTHHQlyaD5SB//gahVlwP5PdOlZ4DZPdJSOmTrODC8GbtSJcAy
680v0iJIJWe7COQY4fbhRK3RLaErawBopiKPF6zq4PvXaQwW2/K5BUnup2IlE1eq
Lmsw2KeDRLSaYmJoOOE5cvI/9LLgPstlbvI2iTRi8174gDq7ZyNG+auRlFvZTU2r
txqS4jv80yL896NkVlZf2NI3fH9VToxzCHDQlOL5SU5qpnQ+0f1uuiMKYGOi5AoD
NMUx5oPb2kTDbaPU4/QdbjzwwmMW68qNuzjFusvp4NjnBgSUO2CiRnSWlo/FWl8D
i1HgZrKprWWddE+hM+U9/37Q/GNc/+/a+LqCoxhfMcQIZGk/90GSVKHTEYOsICsZ
xRLTDv2lcc8IvXIdkcx3KxRAphn06OusnlWtgQmWBX+K1g6u/tzCd59gLZFXaXWT
qjs+qQpEXM7yn8+uwUKv3ghORwDRrr+3yun54Q14BuQ+9DpK5xedXC1nHA6M1VHA
I7oyLCdRdC5JSYk0Y5I0WWEcg1pwMuifYZWJ7g8j2HPlcYcJ7xpF9+v6QcbHnZLm
oVPzAk1gfC+LNm7qxbt0jcARCMldjMsw+Bt2P5WEM7v410Ee+tfYsBGd7nTg3cN2
HkkC+LTwXmlmTyh7ZdI1uq4Q4NOXqPMIlUtpvZ6OoMy1HEExFS7ENcyUpXtelb92
BSOzCGOJ195BYH2XyphsncQNt8cfwyiRLPfeEhM1ODVvZDcDRd0eoUrimicsO1nj
e9M7jZ+FA0OL0PM+VoGhCGsQdLWZerh7C0g1KGiqVY+nnJ/ZSE3UY08LLKYOsKp+
7L7K86ElxCj+tD9pVntyzIB/5K21dS90/5HA0ZABOotT9/pAgglHy30Q905vPMzN
9Xh0XjIgHr4jnDbVfhmL9aUd7KPIqBfRT8DgRzMCqVPwD2wcaoEbLMlSAnRM6C/c
IiHXsmWJbqJ62BSlIMDiEXSkx9JijsEaYtW1WWUGG7bPG02UA4RKSJyCq/VnM4ml
cb8bX5hddF17+H0Y/aMsjYdYIlbcfGQY3M4cpuOMQ38FcbBk6aOxJnElMu+ZNCU8
giSrdIir2xEtAt/Ytrrvh8z3vFasvcYS7p1k+yic5nyyzQJ4Hb4CuhwzB5xMciTB
ziWWyyAD591o/YR30+n4z0ugpkt4Bx/K7Of79cNVpWI4e+WDsGwPApdjJ3j2xBHC
dxsaPf+XdQOf3FCBs72PRh/HlDVSKbqj9EMr12DzjvSwSD7zYwsI21Z8UcyAuZ+8
wC7k9kUKIfK59C8vrJGzyw+aUEpkabF9FKjlJORSAQUGXI7VUIr7wBBE2Obv1mOV
FzhfUcW6d7i7WeGjEC2fjtbHq3H88VacUjTLFZGY7F+bxKL3YLyuTw8Mso3ouJmx
vk/iD9eYfRDEJ00lGIV09StV0Kkb6oWSXGSCUSVpcBwNPdCrqObWxDFXzWU+2Oa7
UNpSrEDkx8I9jdyytTu3Gx4dhqMiUihfxlCdGaWGuhJNJbGnDqWMiwUUW4wYLPp2
0H0TGRBuzpRnQlTNYsymVHwGh27Dzcwuc4KKntGYFxXlguLzFm2j/zh71uAIrYNp
7+9e5egW62kuuPfcIvUDpjC4nbF1joHPq+6jEvifuLajpfsHJZyA40ULwLQC9Z4l
t6A3cIgk3ORG41ZI7VAFWlTa5yZSSA6vpimbvBmkdNyVzI5zXaJ9dPo+ZEPIePgq
SB+8o4exm8SWdsNRrZWhb8IZd539HeqyA+W9JcWktcBUGDxdglk2G4PU+zestgda
90cJ2Hz2hrfWJ/OT17nsE/zhv86S4oooKn6zKPh8wONyfX3toRGMQiSPEzukAua0
N4iX3ugPeWrV3TUYyIZnyVC7a4md65Cvwga4xokKAdhIYeA2zVy4ZxYrMcYylgql
GytTn/n470feFK7iCNFBhzZ6wG30dwxgXkLuB7zzAbODP5d21lFERm6oCDB3h07G
sIkHtziEODL+Ngu4gI+X32sNfz4Lp8GUvboVUzZqE2f6s+z7DfWINObcnlEd5zW4
DR86hs8Auy5VglpcMdUS8KZeY6jruPktCIzcbW4Fw12+BeASnxPbUwlX3W+IaY9L
rZSDW/eZjy6pdIZ8djBYLg99D0CaiuV3Np/J7NY8sgTwdEkPx7A5ugZyXieZxXF0
etAj3+QvCy9KPAzfIvGxlowAq3o2kren4ivCnhvysdc8gXaBJldGt88VdwkS3QLP
57msguTUgSYnaRpTcGYpJN9mzURWdgeiQf1YuIaxbcj6GRgxIxaoSBm09b9cBFzS
k5Om23k6Q0y8xMaYQZrHBed5LzBqzUGEAeuWT9mOiF4dUL0O10wmlp6A8pUZ860z
3ajvJgEmTsCkSZwHt627lGWBFmRtufiTgBD0PEaPWXXxyMMeGy5sjDtuU3NZsXBv
ndVjE4YM41rAQVbcI/yWtS7o23ZRzPF8RwTwSHlPpzQxPu7u2wqpCwsmCIeg+k/4
FJy1TBS5lRIota/ALQPrI1nR463TNEIXSe7n1IG4gjMxum5bPm3Mc+idKBGRIFHx
GUofzKCwMLm8+7Irfy0FGEO+WGaIb520Eqj2YBcdc+3622J/+Yx1lgVIwI9E5PN+
wQtu81jdisHe+falVhELNETzE2WNIk/3pHTKUsHm8QEJExx173hgCYxpc7mMqSwd
/wyYipNxlY9DEM/NcDzEuVb+ikX6Tu2FppLM1l208/h3M8WR0YbMPNl9FsvksJiP
841KZ9gVgxW7DaShdbGZwH07QARKkpXQUZkPvk0W3sSXi25k6Tj10OT0O1tegMHG
3m5OnDYQHu36ZtbfbTUnRYH0XivvTtQELJN2RfOqhC0ApRDEsPlO5xHoEdlD5IDU
KGyQXqrPe2Eu/uTs8yUxLsVyBB21OQbRvwZv8y4g36YN/2czkMExsmL5vesDL46H
pFs7DA0ecysVZLlRjZyBSLOWpxKUEM5NU+JxZOdE9vg5kmwio2zeV2tCeIKIt4Gw
f5xgjrl1Beo77DTvTTfZyp2HP0IndB8Z1rLgvKmugCgMdW9MVgpv/vU1XlMu6J6A
3Ll7mWA70ATUiBcTJfe9MIjHfwXURgjzxjAI0woxPOwCd0TQJHbJ8Yw2qHBz4UiA
ixZhiM7+pmfkSM2LSuqK9ip/ne7zGgpDN4KXv8SYLoZntO0E481dSjslS5rvEjed
Wp57JohcPdVhdK17OoLBG2awXeas9/EEQ205VIN0B7y8Da1JsdbjawT4GAVbcu6I
rHdaGe+0OcVSkBL3AWYfhtXy/1904+kG4H4IMBwmkTv3CghfcNicP/cvQ+dN1TF8
Omj6O5J0f1fYR2OfTtx+dx7RgDtQlUsTqdDf9UZY+2w8CSA0Xk329jVcNMtipOVM
/fgiMUUF5G1hHEs35x7LxYr+0BW+hqpppZIn1ZCOeB4Zn1Q4qOECcHo581Ksjs3v
xplXDtORyTKqyy/Qf0qCJlH6LKDUh6Qgk2jD/UALZBOtEHsaELkVD7WB06C2lBKt
snVlDFuAm5hmXd/9wt9wuh4OAKHR49iCJHSrAGzJfE1VYQHqdKYSx9NWxPie+e2S
+DvF17sRuiKyfxR4Ey3hd7gq8c7DTK7tC94v1l6Zy2zn/2HlBzy5peGI83XDBumz
koShe3zLV7UOjkZ3gJtWtXbRisDvoPM9uYyQyaKPmPr1QbgQ9tVicUwafGt9U8cw
WXHWY+i1KmjngiAMUUDhfIup6YvgGVhazhYjER5QuSWDH+z17nXT9G9X4YkOsMkA
ruxEAKRrHdvQBuZ1ffalBcZALfapHRNI5hd/qtSAPvDoSXhimGBe23kvBqyw8wcW
7kX/CDnVH1fPaaw2X4uvERymH0py1q2LD8XaybVBUKg9GvyJeQUWs44mMpzUGQAJ
95RUORzEpKYql0StGJQh5sBphsMJl3heaoKvGg+gvfcRXmC7Vr6FAqIjII9vnYdH
1B4E5W5nRMaogu+D+t62TiqkIAG/IkhRoTz0i5T4LpeQpLmUKTsjbRjbxlMcA6vP
qy3kPCqOrSvrsY+EeOBrrHLwOABl88k3UEDgPFxFmWfQHOVnJCRSFbTw+iSYew6P
K9Ek4PfLr5Jp3u8Kbh0KLBHLGt1HrMBqlOR5c5zrl2ZA32wOB0YbEhOGS7wGdYb5
RD4tJj4Uww5WeCpGB8Yitcm4ayqHvWhEowyKV4eLRk2QgC/JgLukAG/waC8lVbsc
B3jIMgGt0zwDAV8hNwIkqojP7ke56RHhLL2kqxZsaBUlZ2A90z3km0DzwFMp8xLr
kjpr8zL3/0YuTJEoXb0yj5RqaoveTdJD4SGQ24WTMnhZw4ad3JhFtBG1sdZkXCki
8eLKCHOHFBfb3lW87jvZaPvuBzolRZ+ie1T2vkfDkgNHLAkS3B+u9d4KMgMLDN8W
e6FYEPmBLGEQfsAdLzlc0vCHI9OsI5iJGx2V88NijF6aYt7QhyGyJvWtEtzHvz2H
j+vA4ez11x8r61tmNP10r0AB+7irMNjLUipUT6K7Q+P1J3OQtVRFFln6ECjj6Hyc
v/b+QsBhP8cFDQd2QjUJblO0TpxFLgZoiMQf3km7OOvkzMaJkxDJ/b1sTbG9JC9b
itdyvRPfR27FISRE7gajGQYt4MhGumNqeNdctCA0i3G8Z9BUp44eRutsaUAlf7SM
xNJ2ujRrWNLW5uO+WOCjL/aJ/4ttgIyfbvvJX/y/zvHUOCqp/iYHg9ENcjZibRs4
FZzsxLYyxdPIU+5FxtdORRdQQiZWer/lWYGIXnAefRmyVkJ0kqNotVGlOkUT4BOA
9ZXGPvT48i5F2l7Hqq0X7xtJRADyGBS+HchabpNbjrYZr+lADsZ4muvUJVrrAwzj
dJYr+vd/GTNZkH9hOeKtgxBGCHBrop228sMRhDrC7HcrhZui+wN/bvdBOnOXUyoV
UDF23jSe6FXoMDd9q3/N3U7+j9DJFi7hyVC5hnWYlHv20c/+IF9G4Q0/SkNjxrYU
JcpHUfp65V1yNK71E5Hc6acsk+wtuyY7bkTfoYf7VtB0+xE4MgBnCU6Tk6akXLAE
VytPFtQ6/qTFFUpP9gub9PNnB4NOyxghkbCVmuRQ0qgo+uuuhzGNqx75a3zJH2NP
7iNyx7ZFz2ZoVSokOGRG99123gRLDx7j2v7WzDwsdfER2zHz6AzpIAEEDXsYEUCW
x+ILUwWUBM2Ert1ivPvHYCOLVl/FdftgK6FZ8AaShWYmmkFR6AORYUQKRZ8btzqr
nzgS9ApvFSsRrlHXhfhWthUekmHNnqnmHC+aTv5RrOrSZ+wvNy+kKcafPIZxKYde
D573SC+c7PvFNW0YrSylVO4qwCNikxpCd5qO44opjMe4UajnOnlfUR+ph0YApZ0c
qER3Tq0rMyUFk5J8gn0wDQcjmxieV4lkR96QtbLibiqME2nF22sL7FIf3olInDuf
wA7D97cL/U5aZHedF4vzob7cFUJoEInF6zWUDUAdubYEy1zEJfKCsnhOu7frRaeb
qlXimmG0PpYLXKuXBGfg+ffbixgMZa5ZOLhwE1n19DuZXnPX35o/axwkHwxEsjtc
+hFoewn3Eb6MO8vXof/ost3hMzD0Ejz1+Ksz5PQ8109mnynluukATUTyhi43pQZo
5alSDTlGCdRur0JCDvl34SkLBCTzHAZGXI1h0yzFf5bimD6aFS1KgltwthScrn/K
a6/7Vdi4YvbYhT1OTg7fy+omasfDZwyMbAtHHaK4dOoVsciZgztQePZVDljuS9lA
uxAZmizSW3WSvqALG8qGJlkC/IuKjZ0jnNuljw3vPIw1bFpmEwtMOaAA/CqdEw58
i2JRF1p/xPkEX9kXM/HJcXHBniT5oHkVS5Hq4Mondpd2sQWHQ9NhtnVvW3Q5ewdf
inAX2kqLE8KBhdBhxKqghzOndk0dltswQv8dLGHUnXcvsBu3c3xBjW+L8hxDwbRS
SVijrJZLXF8qsM5Q++1j1mPuxhg6GSTas/XTicJVeoWWnzKUjT0Iqlnajpuj9Vz/
YgrvTTTMLRv+f9xgZhVApoPp4I8m8JoSqlqFriOGGl8Zdpmdvkxr45jb9wEOyv2p
t8UlfP0vy3WFXZN8SQRxKfvhzt5guG98JEhhQHtKP0s/yupuAE7E8oU+huUCYsq9
J4vqy8e6jhnHA0FjM9PWD5k3gpUSWAdR1H/UMwfYVZZcFQALl8JWgr9oi10orIoA
TvwO3dZKEQWXG/bTNyXygIfXwTHFdZ0L9gOQT40Ua5OiOzT1bQMsSxr2sR4Sdi3q
Fv80aWJjd2U5Kq88qVikWO+tMwth+EdOCAsgme0jF9frOerHVQ/bi7rYb/MTEcSg
EfldZPTBqzguBnw9Dznj8CDHh65/zRDIBbWWdojSaSBThuwL88fk9ZvHjfcQwHdK
jt4TUb7aYFDU7no/CpG1TnWC7Lt2XEVRO6QGIqykceWXk2nGTHbHNUA+9JBIKGGV
H5Pw8Wkdda4hDTTzetcuopbO43BXz4RnmAQpG/npA9Eam4iJepabk+MfqfR3R2PI
6/Jg+W0IZYkIVi1NXAIWibP0UG7Eq2v+kU16UzDO+/W+Sl9/tNlJH8XNfqBrgfqz
85pnLIyF426fF0hbTiv40zzG/KS4BlPZFkeHFv7n0YxllSgK8UncADQGY8cVGCpM
jqMnNasruidIjwXIVM85FvC1OiexPlvre6tVoaBTQ2AhP/DlIIht9JXq+NYAus7n
FwBzf+D29Cw2qAKjyPlWu0iiKopN49ZsccPL2AxNMb4A5Na0L74/AoCn7MwOibNS
lI7m63wOfYKhMcMKpjoMmnF2EDKlFXBgvQIyrwwUyGxIr4yWXP+ZbbusAir+HxfZ
NCZYbqBp2xM7c5AFFdkVMEvXhJ4XEE3pbyC4o1nGfe92MY8y4zipH8UMzC/s+vyh
umkhCgfnBD9MG4OJWr5XuDF4fVqqAe2UzOoKqiRbspOxfGk97rgugMxyHbGzvU3n
vipnqMmVUnsa1+9eqCpIxXR8qgZAtkwjLpI+KHYdHYPPPUA5Wl69v5NZdMTDjhrD
j4e7Ah0quMpfT3NbSkH0t7W5oQkw1ck6lgNyGYlje1y5XBDVCbqjYaMo/1qsV185
QzMfokRpgojdOBxvIsIqrO2A/bz/IGKAw6d9/N3UE+BevUDQFxe85i2cizAmNM7t
qC8uCMiFMYGGMhgu233UqLoVtH0xRgVCoMHQk4eCjKMmEtjlXqgRQyty6Y+kISdB
kFyyq6sSpXB5ODpEysw0NGviPIBLYQsYD+MDxVLA+P0XrynJP6uhIn9+hJKye2vu
uWnf6GW4zE1Y3hIhYI/kB1xsHEtqXDY6mbwqN8fSE2NJdwFoK3P8BrQiWfw3dQ9A
t9D6fJYwjHrxI6A3EYMnSBzLwmq88/yw2+JqaB5Z7it/WqlRKmnx+8JZ98ZfCRsc
sAC60phOjj7idmAmw8CXIVu4FQOYpucJn6fgJ1cM5wbNotQDIgHHPsR8z2FqFXeC
UYuoClSbhsG6U45CYGTW5fn6KT2oDs9hqacXF9ALPLI8g85U/pIGJRdmH5yWRhEs
Sx2HcsiDZhNdHxEJlTV8VhMtOTMF/X80dyKUnPiMemsEFlkfYbZAF1VyQKqkEf+T
7C3WHW//E4r5NYE/IDSxJ5NPf369TUnni+lNawwwkXJHztqA+do5hDWEJ+kAyk+3
5L5DyvZ6r9KH6mQ6ZMCbMWGB/z8PXqPdbrRMnaxFcHj6LsW+HF0zrc3MkDONiYTA
+fXeQpZoEihfDxZ6DaUzLUmc6aHvRVTzUq2pGLNdQ3ieum76P9uidGey9N8tdf/X
4v4nzID8a7wDRhhUgAJ+WirD+YjlqCSHNjdfO18t17CW3zAlW9d3RWTDRPPg6oLF
9CC5lXCHdQPafI4nwmXQb5WTAgZm0oBqNPEF2g+5azICFEgwhsnr2wVAqg89EexK
0IBqa/2xjl+AC3cyVOgAHbpZYirDpOXqGILDKR+Fqu/rybxfhSsTDkAha+oNQ0ij
Fj5PgTycuZ3i4teo8VrQKzBNGXoCgFPZBGl84alwM9e621tk8HMmdP/00Wbz376h
PD8t3LiLQawRQyPcMQccZjbAcLt8Cq2W5OiUYaxCRJsDqpYOXuoOiBTxrCho5rWu
f3ODLfo5C5DtLOV8A8cKuI3t3Axy81tJAi6uDMNSv8Mu0qiGcqugEAN5L7cL6hbn
LkwcqQ+QQNuB2RIo52WRlVnT7zc9IB8a2Az0YlFk/FIvzDd3HexIl4YK6XuYMNjC
LNnhT5hyJdGLMc/IkJQpBYfngcZgtb0g4H/8kZM+5uue1xLmK5retWH8ljQk0XwQ
XYimA85shXGE4ZATa3nVFwDvAmF510J1JkaQG7o/bbdYOmY+kPSdfeWgYKj2K9Ht
IVj0HnfX5MviSRUQqqZYIlqrYoJiY+mWJBnt3S7wugNZyu4dF1FzBFpaekmJhdfW
W7Vwzkyu1hg4aFiUqry5zY2UDT6ojZV/40NlrOALss+no+IENGN993sxc2N1EPq8
9fwrfVmjOwjRSPP4bRPg8OfihDeIV+mWgwyR+yhSKhlJoG7gJOz1gX3S7aDEgF2v
j5u2z7fKHRhMSDH40XLzHM5j8fD/k3Mpyu4+uwLuEjQmbNQ3iWEWlItG6ATjtfuB
lrcq+3s9gKaqiaux0SAUfRoAuhdZDUY0HfwCuBvwqZhG/b5QvI/vJkDPirS/ReO2
BNPFWAKd/3OMpBKbY32sIGaNuSbZWz7/1xqAi3oB0VrRwmOuxteD7dN5dsUyOoQZ
96yog8P75lKr/nSWGX+Nmt+C22nfszvFQ0lqdTchDII1+eYftnGKW8p7Of6mln2w
BnreIfvedB3+zLNWAajjF+565gk+o7oybTsG5nptvTzeU5DuldXmxWu2Qr3JZ+xp
5+UrHg6dH47Ojs38i6Ylht4FicVSM0rxhq+FPaZ28WLAuFR8FuFZnMNbxsaUxfpA
Iz7w59ZzRrBByLTw1jV4UiuXU/PFPga96Sw5VR/+FQMBc2InXx5I1M/+77DfN8xr
LIvpamNkmNmlxIwH1bcBTdhhR4idpP6PZCwjZInM6NYHezfAtuVF/6UdSmaaE9M0
qdWayPPmKoYbSZzCLWeAAby3u/GbYtfGVMl9F2SCZGPveywmGzPnfKz8hBSFWp4s
f7AqEUmyYmM0CLxwK3/ELN49WTUZ6NLVsgHnJVkIivn5wvcxBYkCHnupNTXpVvB4
ZHFP5OJxyk1HbhwOLN+K4xFEEKrzsBndoOYa07b0eCRS7YpFqCpOu8E2d/gKAUyg
IzOgroyDK/KB5zSeV6lnnWUq1DTRFDzdpV38mWoarjdfTuSJKYji/juPHypB4rqp
DAyJYqLxADDmhrAuCcGQbzumFspDAEn4qBS7KfJA0qmm/L7K/J/myoq9AWyv9OFw
CMZ/k2NQV/A01p/maI8vklvLV4ocNU8I2zbQq8XbDxUOPQr7m0d3aIH5U5UGW/Gt
DdEHQycTIowQFhbtJaxf6fIrx1O1BqX7Gtb4IXY6m9Fgnw5+2RVo7DWWMqDuzH3b
2WxWQqZifg3N76ZSKXVlowCZC24oXNBXm/Cl+mYKAzCOplPx/aapOWE4vXeo2z4H
+57FJSAXsHy2vZatazl6dL4J1+gWpMpZzlSlQKrDuiTKmJUig+OIFs1JhPgImXeM
4+U3rVps41/ttDdgTCcIdbfO/hKtSghW6HQlApx/tBc41SK5KC10q9uaOj+eu0O6
Eg8kvBUuqPzMd8SdNpSz0wUxPwa5KqvIZu7NXozBineklZBdjEdg5zlGuq4OEkUr
VzMSRF33cmKIudAen6qGo+GYGamPYaNze2xnF6T3Yc3BljPHhoxhd9Y3IrqgRsiL
C6Ff3D6bGMN5+wyv8hCqG0PM3kc9zKZuJMEuU5omg+IqLoTxAzgz/s4QxLIBFAKA
E8h6P7LaBSakVJEbPdLJhZlGoIJS98tY9v19kkxjsu6D8D/Om35cRrWwDIeRufmJ
j07RGYY8hJjLifoiNkWt1V8V23pQLljkVeQ7shX0xBzTj4m4F6gRoM+KAlyOqP8U
BH3TKyXnu5704gst2uyYlXIYW5xYomjroI2bXgxyce8magZQRvobFO2pasQBIB+6
RZJly/VoipbSHj2mDlLke/U0D14/BtPh5oopeLUUpJL//TI0uLCTVRavSyK0vVCs
Uy9IqwBcodVygEThea/rA6T5m825oFuC/htEhI86UbM4l0y7s3OydHKrTk+E407l
cxQF/OvaSuOLOWE0MOg2Uh43c0cdBHcOAP1oKutaaXJbSlUY0Ex7M+vuWArmyqg4
/WSxF8MXt7sF6QgfeBni4s7hrvIHvAEhvOEfZUQMmyZgkPgKkt+M14vU9LI/kUOz
Ov2KXlPZEiLTymI+Zf2HYeR+0wkUjxIgp7kY50SAwI9OQFnjXxCRChRbYMy/AwVZ
Yzx63tuSho3oQrIBwHzFRGLVmoc+7PEIivD1rA6LoMf8MQa67zHKM3C/LhCxzy3C
8UsIG3q0eQUZOXMfgkrtcQ3pw5e8kbOh8bRP3eKQ28mrTkS08A2bsoA+SRlvJHOc
pADUVO+ZVlsNuUs1g0JipuUZPZ43Lh1PwlrJR/fIh9XSW04pgV6tp/uTzG0vxH3w
cqIGlqLyeQ8KcuFrh2yT/8OvX8d08fyNdk2JAkb3zHzwkHETMsfCdkJC7p77pOfm
UT0ZwRlSkHXXtzaSVqJQRZjDeeREVvVRkdArnOYv+/3QRLrb1GdLTZVrhRlFilmD
pBuH4e78lryUo+opyG0H8NinIIVe16rnYsIoxUZ0rACmAuqqDjexn6yvXQ4JBbil
q4UmNh+62w1F86ZrwCGY/BCWEde+BcR9wh5F3uS0qLhsXqdVyU1jfZrbg/yOmL8R
ECQwdwvFgcl1tcWTgxo4p7iei0xI/MMojNaexHYgeGJ67qR1Ef7Y2A+nEm38yIeW
g818WK+WJ/C+n/QqKAil2ws/FeT90V2cu9QKCysZ5bdjxAoqNJJ9TADNRrgziozK
5y7uvF47gKZ+0vKfefuiTFD1jmhFHkC4i/PWFBl2eb+kJTb256AAH9BVeHfjrGpj
ODfi0lWEGWt42FDnw/HP6u8boHg839hWkg/57/1agwDj7yPHDCNwuYHi14EG4560
0PlCmktuj0KEBTOuVAFVykMODI3G3wJheTHlL8OrwJ4wtCrGB8QP/cnUkE25E01e
J/JuHsYPxmU9a/E4n7LPBZQljTxAK7hcgGkK8rUEfTGZL2T2wpfoJ3eIaqMC0RXD
biEu2wLJtcsl7GmODzxhWLuuVjD99mdrfQotRFVfM85HhdC9fk1hx4kmQMejj7ud
HGB0JhhE6DmphvaR7o5EEwC75TzFuGxPlHICUfUyJ8DrGLTXHPQ+H3ojcz+tJPOr
/NBJ37iCYXdG32+5nG1Zbxe7h3PnZ4ALRi+MmAYlg/JGxCdVOonK1uS6iXMAF/be
JRBdTihlaq/07hvV2+HRFDnJ1QmCdczTyrWQnRk3odGLDLwpm7vt+Qxgvh+nAuvW
Vzz7El1R409a18q6wYrQ26EfSYv2lck2KEg6ddOIYYAhR3G1aU1W5gbwA4GN0oFp
N9l5ppQruJE3kPpPpPam1eCsSIh0ac8VxeJ75zgJDd/BR7eojqewa/sbLz+UWw3D
ZAxjZZToel8Ma29UpAgCSTBVQPyNJ57mqaxpJGi0knT655xUoNimFfHnGCwpGX9c
c4WQBk2FQGtmOVk/UCzKnbduMcD0nNGw72V1pHViOU0g4kJpgi0/BCIRl2pEy19W
Gj9r9uvup6po7ncjwfV5S+oG+ARDiFqiYi/nxPAKF9RQppzt8TkgE+eZBLKCShLi
WITwWk4pQkPfj53M9Jgph4CD0DdwniVXLN7OSAx2Yy1q+VAnc//L/akohXVb10u+
eTDMapnbpCjlhNiMvaueNyfzLIHjtJSCnDR6lOqXBicrckSNu5pTafymzEMjvJZ+
vGjLJTTE1W3ZAgzdOYQX4WSqGpddvCPtXueGD7qoRUuzSy35llbrfSmoVyQ3X1uK
f0OAwtQ4P5UxIFcgAAhhmjvnlk7DNzl6v/rDdu5yMS/QLt0tYTmMw1RKUWU+v3KG
mINnAR1J2cF+42K9apebJgqOHgVXxvxRsweSdYhC3aR3qOOVcyY+3lAwSEWBH/wt
N7UmZWhrzqc4VHdCDGfLI7q7EuPYog3MuWn+WNnGhhp8tRRIP8AwfmiyYhzGnhEW
bcGVrIDsKKy3AJOiiIWZ/4qUYXc4t9p/2IO+Mon5vvDlHxnmTTKO5JRdHHzfiPxq
7oYjenkKPqNB1IMIAH6TQDdtmtFfXbqrv2cnqL6dBtlpv2e6eX7to6K06v8Ltp16
DxKb3Ucnd0o392C8WDXCCVuCH74gmifhNIY/lEJNcRMuBx+dfgkGCMxE6cxfSbWP
iiu6vaPbUJEWIsL5Yh6YyC//O5sM9Nc1xBs7NJ9bLSuOHhKMUFKdRcNlVi/CotaJ
vRUGNmM3Q6oaBoQKdMawItfQSecGAAWjYqQsl4y8Em4TC+iCFXdmCMGJFhyAwYef
z+3OV2Auh24xLOiYBUfUbZ1YVuObStTDrBZwNPGKJOtctUwiC2Xf2LP5SIQiYAyB
qUbHxH7DUuueiJ9fZDwyBjJ7TYuRLfVYRbi/JK5T6BrzLb2lkZboaQkBbxJnnlg9
oxVEFt+X/q/bNd8JM83Osw63iZqO5GsniEjRPArvMwwAv9cCxkggkPQ1oSqmhTn4
CGlo2Da8ve6cqnMKM6qAR+NoF6eKs32Ia6ieTu9z+cSoCpPnS4dgLdyTnrGQwgmK
fr9c2JZL01wByk9XLtb/hRiBRRVihhtNgammN+upUDUvZE7stlmbTvpRY5t/p3Gj
0GWIFnMFpZwMIf5TcFeUaXa1G+4C4ghTwl0xUJe+1NmPWdPu9nOHA592kTf2bU/k
5mcfVbJXUYJFpjz2PuQSPtNjJOS5r6sbg4YFRX6pZ6CcF1xUWnhMduTzr5DDWSAd
gya0lqd56ENojlUqSyIUJivemSVkqovzrpzZgu3s297D9B6iqVUR8kvPEPp8Mc/E
VNlwMDLQr/ij2zD0fJit05Rz7XdT7hZEgjMuhvmRBzetTj9N0KkZZKLLQKHX2Rdh
qrlEI8f1vBxLz8ylxJryonvBTlil9gvpYXNH8RLFGuwFcEtz+C4V71WxoQPpH14m
LlMV5RqLVsLcZPvscA62e5JmNcTGcqwEIrPrytJwLwz26edyC2V3HbKXahstQgcL
fTlHEoL71N1Zkdb6ztzjBmJAJh5/zP0if7cZ2GRjsLx1w9S1aQcemzdAPLuIJIsS
dUJzTG+PJKWBhf5h7+2ihrn6NRQXQtJyL6TlGsqZ/R+m4p7MUZ3vMb1Vbc+9XUJE
bccelhnXvCTJQF/8tdrQxi0DFwlceacLcuFDwb3reaSSMDtprzidgyZ9yB4mGP8i
CMgaR91eI6aRQjvf58B7E1rUCQEdt/M7QqzHjY51E9zOpSB4VRy72sUpM7qWfPAu
U0jzBMC+G86OaaZjEbnmc+JoC91ONuDZ3GccFQdE7Q/SIXrdBG7bNHIxRwFAGERR
jCkMvvhueYbUKrIaAzKmd3Fn1Uj2uXvhBGeYrc7HQvCspMWzRzBM73KkAqQ+72TI
9Ucd9loGj2sCLDSvbccGfn9S43M2chaw80aQfZc6tKmBBkGqae9tk4v7xo2MJW3h
rpuuleX7pP2IstWDopiwAZ17eOwiVpUu7d+FylEm3e9HXyojsT1eFht+VykSUIQC
TcOYLl/HGfz0GqUUlJVPTIG78hw5vM+dqUKWoT4VldGoeKKj4MCxZHjwppQjBxC5
JLbBEGAZNg0yIcVqIEEN281+q6xLVZ/PWPcLWTT7SWXp0E/snyW0IhMbhs0nXeMb
6x/LWf1I4UIunRVKunL98MvgB6yJJZZWSaeAn65u1/LbwunQen8M8newavNd3m23
1qF8e/m8PXkAhpKf5yqR8HVyFLfMhq+3iXuKwxKiJh42mVoCCxiir0ZBQBb3waQh
hToB4UHJUPqRXS6W+YQDjl8h2n6vAZ5VxAgofmsz6Ll1spEowpmU8ATzs91ywKal
S9fvoGCJLgiNciHNyDoMHd+e9ny5TLLXwfvqW62g8ThRoePkfiDLAQHcna6bgWOG
g2JlO92VxVtGYYQCmezx2EsJ1eeOpzca9kBZ4p2ier0hN5WUy3p3nxNW9TeL0Vbp
cggE7AoQwti3IoWkHJfoF4RKlS/YlinEfEkaXPO6IgpwAroVKLW+6vgvhGJXbm1H
EXZIzSM2RPESQMQBoulFPNOOOJysMHHO/E2vfD6U0ue0aIQXFKEfygjokOt8fhFt
16D1cwcdNomRoWLW7xCy0/SFIViXcFeH/UUl5zj4M8o+I0MDNGegPIsNSvH5lrub
QykkS8x9Mpq8qaANc4Mh0LDUKTByrUh4fTqSgDbbcxLBmMySkvQNuRY1sbLEZ/S4
3DSg8xdL4U/BhjdQw8J9Vlq7VV4sU29yYYYAhyDvMEnKBMiqzWfG+J+9cWVnrSBs
V5SmvoS+RlyePiHZ3FEsp3rqTRyL3XBWgKHwg/z4MyQqW2n5727KIo9Wd8UIl1Yg
jdEh6wcOrvAXRyrS5hCIObMqX1COvV7o+4ZcepKmV2dzXewGbsql8PyQBKJW3P0m
VRjTuQVnvnny43r1DJMEX66XXfxBnrPzDgizBWLCBJbvxaR5yY/W/cbQmd52AvMD
1quIroJxEr1TSMjW7yZoXjcTBdN+EQx+cQp84H9e1YfMJZ6X463LfABuL7jf4NTr
xNmgvvWSYv/qHyPbHz3vOENgyhS5IP8D4luAKsSBA78y9Sz9geDIpCNW+s42HuTu
sFSv9AUbw7BVob5AZDeFQMVAmDb/4YDW6lHX07nj8RBasm3JhKqIMZEKIE7Q1yrX
DewAUDjiVYYWeVqFEtBuG7K0L3YzpfSMZ1VyPvUco3Co/9SnsVn/Wht9Q2IZMD3O
hY0FKeE0LJs/Z8p8i5ksu5gDjiAwRVokiVwzXIthc9gjYjSYcOLPGcCIBlvkKh16
3bVI0111hxftv+ucIxydZYvLbLzWzmzZzcNK//9V+1nrNK8LUrQ+Ko7IHyjqVVKm
ULfpJIrHe0Q9tDlTu+ytnpsqkV9HtVM3KIR1T2zMPCj1xea2kp4/X1wNkEtShJXj
AnzVFmII3gCCrCz2zrcndqOxTUwzwo/iVsMlH0NykWCsh8OXZXfSf4DqGB40YkRc
SNLtHpC0fOjT4/45zQ/9lAYzzJjgddlOvmsoGJy/s9B/5j3E0MRORaTO8WjNZrTZ
ZfrT5sHW/EHJbwahm7HrKzlzNvdE6mByaGJRMjg7UqJvEl5YnC3w9da71G6s30IZ
gqqBlc6fUvbISdFWKLCPXYzpni6O4iUWXE9y1ZjaFpxrSr5U4ipsA5/CdpfhND1V
FL0lJ0N3vg9/yJu1xDgBQlrq1m08bz5Z2dgiB+NwaWq9UWTkOtF3ynGhUKd3nvD/
D14YDZw63aQ8cgN1Z9xTG4byPADd9ABgKJa0Gt13tMeUuqERYbDdL73n7pmZ8rAI
iO8uCFVqOrgdzUl0j26vwtWTM3BAbo6OO0wb6wRX/wJ2sB0gEJgipmiwCAS08Pg6
cLWauyd0VEZ/NhIDn9U34dKVUqNebUSFL1XNnT/fM7FMIBAuyXHtYq0KyMaMdaoy
D0RzzkafCAJlAYUxhfwIEWcFtHS/8RNwYNA9AhdlJLL9weACV7w0nyXDxgZW0LpP
ZOzveQrTTbu99YdBgChwUMjfIkAx03vITEcVzkALfS53sqr8fHBLWoSvuS/P/+7C
hRXuroZ89HhrDlHKR2hyw/XhaDVyYNLCy7QGRjos7Mec+U0/rmeTwomIXyo8SBrr
q3NVXt8o6eZ0x4Irea0kgov2KQHh9o38J8jJyUcB3ARkNkhGcvLPV3l825Ub1rsj
hCRFSovoedqnmxnDKQGn3JXIPJ9SAqgb3qSwNjf8rQVuGvN+G1Cwn6X7bj8Oakl5
E9Ro5p9HNYGqISUds9Vq8C04gYMefLLrDz6oYCDwJk7d1Ejfsda0LjPgZ7K0QxC5
i8rlS+xS/aE8nhWfMjQZji5WnHqbpvTfA0Y+xtHvyyjJHUj3YE6EqvxayF6PJOu8
7wtZjG9xU7re4ozDdhuSYvMj5nGcqQzeVjIXNbGSQ3u8CDdJbdFWDe1s0Jw2FPJ/
TEfM6eTA9a8M5iY8czdlNXmWIpbUVZ0H6eQ/3lv7y9W5a9Xyk71RnvTZiaPgNl84
azf+6X3tM1bwaHzKlCWOuaA8ux11AXQYpazi7YfWVck3zDZNVq0P4Mq9HulnGpVs
4YyvJjuUcAeSIL8ditqzcWEZ82zykUm6wtOJx48yXJduONpzoxQpGn/1ywN1XFAH
VIvcSkHdDJej5stt1UDdK86x5uzVAKfvUd2I1eWoKJNqgOZF3nHnaRAMZnamtbdb
u1iPGHiRz3qgeAc12WM344Hm3mxE0MM8fVEc7UqZfgnxjod3vsJ531OsjZM7W/ly
2oJ0uUBItE7KR8awNolPM+luARYoUR24cbnT4Gex5fkv7O6+RsnsHyFDrLZmiuFe
kY9tL+/MX96U7Juxkq0todgMo3gIHz5vWj7p3Maq3pW99pnnCZM65ZQ0vKKLZjjX
kq3fxRRECoKAr07e5A3q4+liCcHxVn4MX3Txh01fhtT6JxRX2mf8ImYb5Fi0Nv48
tIsJSrT6/jeajknVTiIYuEyKJu+SNjmzpyW2jbCULCKT6aDG+eGQcWKtDsoHseI3
KHmf+WcK7egjKTQrbfDoqsjVBhzKtCChMOPkU5HIKeTWjkTW2exNAExJNG1WhWY7
11JN/E7mImFM6fj29F3vl0nn7vtAnEgjk8fGrtJ3CEH5hKjo4Ih377qEmK85/zgQ
d4AjkODbX1JmPxajdnwqXE+ANrrpic/m/bnz0HdKB+DsSViSfkp6sHLHl76iSB1e
QOzz33KuOOLE4QbqOAfxe4pVg+dEiYSYCpLJB3HGjeVpcgDzDA//UzPQdmRp0lPR
jflBoHzGMk2R7fr+6jZAj5/j1fgCklO35wG7yHbyGzzNJhTu9yGKSP4AAsXQEgVn
3Vqg5gduoffZWVLKoRySqfhQcE4f3CpcbnkSDddebxJQrav1QFWzDBPGHG7an5CQ
9Ow9I3/FUeGG2UJT4yDtlsok0MMqXkMQteIrMtH24ereSgxhWx7xfmS++Wwn4cUo
/5lhC1Y8U2ZLWagT+pEDhGoVkjpPvjKA+z4geoEpZ6As45vZSVQnmfPyQTZ9FLWe
dlIt/BXCdVElEvKjos02VhkfnFUS4gShBD/8LYptT/AlpbCnzp/2xGS74U6HAUmP
8moVF9nlnTaEFRXq/cEriIxk/wx9p1clfm0bLJ42kO/qX/w+znwV4ksVotQSKzlf
DjYd9jzF7MjVOX8ZnrH/PXvDvp67KJ3dadRYnoui+gGkP9/MlHPRAJd/c88YU7CT
NHdnq6ZC45WPoBhubYFUW6bgcvYuemLA+SBu64r/SUCiQt+ictG5b3SytMQ7KG+R
QVPvzdEifg8qaOzgOibQ1i8YUS76YDXmLBafObzVXNRk0kOPflBSobfm/v89PLSo
CFIZvalK7qy9ryRfpVb50gt42f+zWtz1OG+dnvzsVb3Lbsfaxdw7bTdzRnBXXtxs
kDQ3ekuLewuv92VYYm595BVIZzgztSbVODuaNeCCmqO+vsq2ZlcdeQzW2uG5TrBI
OZRxaSSSsE1D522dS4ONCa+6K2qO5YzBTzcAgvj9Lv8+bKgm3Dh7KaKaITW/hQt/
JLkpIpw3jQJDEtMitlQIP1z+4GlI//93d5uwkdH+70CREYt2HZxSBOx0bXO4Xsgx
rTJNpDLB0d+VSvx/x71KhX26Fme52SLTt+8tZ5cnJJXKdwLAyPEhkN2SrBveQQUA
Fce7RaEbLou9GySXoOVfLOLuA9Uf2I8iVIWYz9zvhZ9RYufyLBwPWJVvWlNVcE5w
UB2YtpOgM44fi35dQslwHRUg2uorS/0yGH3TOBuImLmzrF8kbfC5QC5C7hOteOz8
3YgBOpSbxuxFkJ/bRk/Rl9P9V1C3dki1izT6UKIP0PWiwmQA7X6wSWnkUnry25KY
/o+pw8eP1IaELNJl9vlPQles/WKdK9CuqjDutNz+cTZ0ceTJeQSnHUEvUJsfIdgD
MvNwkELnFhhq2v7e55Dx27lpoBQ2ZJilxADBAS7c7skK9AXkuD3vsGbU5656S3gt
7+QhuggemhjeyKK0Vgumdllak34OycVEkvAyXH9ogsIXr7fwj1nSks6dS0R0viBj
47ThmsFYq57FKAM9flUFpOPHLTF7G0digyVaG6Dcb6YkU3rSOS/Rt4IqYEdZJ4ge
TTL6UxMji8BI7j7lGkuA+ZKvuoz3twnK4j5CgMazmPNnJc5eCGzaFwpSTudia0q+
vFQlzYom8xOtNDs3ygAttNKx1nccomaB/xaJXECQRCiEqsO0PyvI2A2Q3gWrNveY
focHOMWz1TU8LoqeijkWtd2WASR+lrTxRM6eke49hDFBOyGsWrvEXY+T43RFnqFQ
Xdzx82nzzNiCn4TkhUnd/VuSyDn6vm9bivJDrAKGrdgeshTeH3fQ9kFGFR8sodiD
Y7oFr4JH28NpgYNPlMGaK3spuUq/VO5wjafi1HoucyGJUpZnYHTzlWTf+2+5xFDt
OOvDQ4yxytvdtSo+RVtyAmgIadNy0T+mUJi43LELtvqudCZey+T1hwjpWrhOj8i9
DTBQ4u+OSejHnV7Tk8WnoO9mjnBtyzfxKFLsJ2eqMOOpzguyJrQWHZzLUsiw0Rit
P0tT/ofjct9jnFicSQCei9LlJnt67RKT9hvG+ctBqkzpvezpWV3r6cukjEu2Wxks
fzxndoKzvFD3eGBRXnXwXRuUj0/4V01R+d76Vxe0wI3RKpA9Ft1fR5KbRJkyMeMO
UVWAJriC5CQ2dXGiMdpSWzpFm/SdFgqIyIEdTHeTlnUbFbbxe681h6kMyeTClx1D
VmpaduXxei5N/tD7e3JKI4Mk9EqSDqqyYXpzELl14Q/aA8zM1dtCiBkloJgkrxKL
LSGBYjYib8Uk/XgAm/c1EoV7efdW9FkuhrqE1SzfB9AhYJqpXaKzO+9wh3VoDgV/
at/Cg2oE2rCzzuevPAiE4l2j8smnpJTbXUayehyWZ0r4zLNpBeDdB/B6iSe/EM+H
qKOcEgbhFqe+W4ZF0LAPRrKC8tg9B3fTY6teF/D8/tdENvXQBuGsFxKngzhkmsnH
ATPvY2YAetYcnzZbAJJ0Drmrmnr5y4b8Gc95UQKez9keV5XQ3z4sYOBlZZRKtHdk
LaXlLAghxFEsFBcgOc1du8slFEUURGERmraz5vponYCcjSsTGbHrtQ429tb93trd
4MUM1//v3V6yEY+r2Hd7kL7TUoRxHknJa0Z883rPlAPTvJfTJ/N1XFj9WHE9deUQ
c1bGzKWhY0hNwzD+VpGhryiI9beu51TBE2RsUFHC1us0W8wZEanNVamoU46TTuKw
dez1uPd71wECfy57XCtNcGIqckhdCmXl3TjegFFigecR+3T8K+net+Evz+roLGWN
T+aj1PjlXkg+5ap6fdzyUrdwuGVBHbJTDeEBvvugw+qnwVxjGkJ/mla2EqScDLn1
H19/NwWD624g8a+TYfIsoI4fwOPt1Gdba/tmBV+5ssBAMWnhEZQfLjQvlkeUdVhb
oUbj//wzQ8+5ElgaTE72Z62JxE9oXPOXEKS7O+Vz76YWfoetUBLm1cEGJjEbkCnI
TjMqnbSgRztVU1K45g/6StG2tWd1nfJ+E4aaQuP2zU1gBG1VxwU4jY4oYCeFfVHi
WG9evwECzzgS60GYG4ZJUmzih72isusH6bH3JBkJCvqEfT7UoMKv3hMvWl1NbYWZ
kA/HfVNd4DJFsDvkjaleO0SYVkuEIaDZ3D9FcLac6VT1vg+prktz0E/o9bYEJHfb
VMFS4Y10vicYmOSPzZFVIz71gorcfF9U9sf/gXaSpT7phcgJH9k4iK8iyO6EzZBv
m+dizrI4wj0BgfV37sG8GpXCQHZvDCKK5JtdmqwmnhWcXwcJLgsqWJHaADTn886B
vpqDjUbmdsl6eRS2sm8+OgWw7IdcMnJRIzDEdOvdiPcMnxyO8batdJ2j/8Otjur5
LeWEoBQiCXFX1Gi87ru+WgYhzYby2P4ojH3NOvrcw79lOY0yy9YRS3/QYmNpQOAg
Va6X2DrEm/zsTMNcp43nTPslhPNf2ZqZN3WEO6eRBuU/1d+ldn8L8JdKoxKhdmaa
89qF7HsSN70g8k5bcvGC9+P+FeZJ01yMLvSlvc38t4qexokc0aQDo5YR0RN3hvjZ
alSMzlC7ZacuwT10OFlmf1zDCbU+qgkNWQqSr9XPzWUZjj9SyTzBFityqldWbfSe
uUku24p8580rHOXy2cLquQ1F8wX8VhUJcas+YBk7GGadw5gj0jfLNHTbNIlTBLJo
dUBwXbjrXdPfd7X7B38F1wh8/Rt94SN6dj0lhjmoUFqChkuNI4ajb9n1LqvKsrRK
GJk8gEXdqrVyWpfYVHLaaGOyxb8guonMvK6iPKm/h35UGkc0MYl5ntwTuZHhS72M
aEEM5gT2iSArCHjf7g22yyZ06WRLdyq0ofOEcbyR7Y5eL8c3WAoTe6dHKyID7qU2
QZvo2HED3C3Cx23G6rUvDvHaES7pW9qfmYZ+tAXVC0HAXJhIo+gtNcej9sYU7bzY
3ZazvCHRIqfydzws4MPLJlB8gPJvz1e0rIgY7k0llRDE7/wqLmm1+E/6aLiENoG6
e+nxWaP2bdK5It+TGFEwejWYp6fRUPciTEZJKLoYcP+IzsyVl1o7RF/Kr+gCWHOe
LjgNzM3388CrgoQKqocaJQoR/qSls71SWFZZZJKK8iT+VjLcU12mpPBNBgzF+r0q
UNUQ1WCCirIJZNy/smC++wi6y1cAkjUiYI9NNyq9xNGeDsEa3p9r5btlMukaQoZp
JTnFfwopWErNTaPk4dIKntO79Q+b3z7pXOFnkMN17YjFK7+VGW/t5B3H3siNv58U
QAiQ0P8L0aTPKeSQjIb8/9Xs3N89eObloxEYFSdAIOzWE5g+ceYYW5WoesfHR6jd
FuJ/vT+i1eS3DgX1PZkJFcGj+YNYM3//BD0hawt7/G+j/ZkM1uR60PBw7IQ+nqGn
Ntxb3DoZ3BD9BH1kITDx3UmJz0AaL0i00LCg8ZkXq3CFifxHKDcqjU1KEc+PkKOW
iRC2+a1HHK+LgH40pXkwCEpayr8FzsOzgDK7pGApARwnqOlkiuMcUNZ/LOLc2kJH
di9/OA/2cm4p/2gQ+I+5pVGwgwkZ/LfSco/uZ/bUC5dytj3DnG3wIR08ykFh7ebV
hLxfpYGfpo487bvtzpZWgRFH3SrK0atckdzsOT+DTxBD+LHnPTFfR+Bx45aIA23o
fMN1xwu4N8pXvTNKKO/MiLvlaDbkqZR3m2ChWeFH720rfX9WEx/5uMS+kNg/ubdP
34osZWObSZNTwuSGaeq0Fk9bzMtL68vZXVdsL/uoWRcOsMO8PIQ1uguCD624qFoG
1aTKp+ttHOEQhIbdeXrITIKKQkuuGAi4dpohhEy/B28yDJswy+mN7/c4DGE+Mh65
oaV4SBL5rKg6Z5jPWkuvyCq2AKC3EjPHW7NcWh8H+3+fhZBY1iCuWbX0gEsbMtr4
5hZebzSuR+BnTIpp4jFn3LRJ4r5MMJteZ6A6KdnuDMklD4aE4oCVBB9DbUdDCUUa
vGE/o4WwltTOSLFzJ/7dPTCUU0JCymNUGdyiWzQRuz4X7+PvRfElwWMf3sOzOkrX
vm/MUG16pYT/a8EK03mPoIlGIdWLnwHZ/HFvkIK1r3fiHoy2INNIm/PnUyGWXRMa
Ns+4hN4m/A54VVENf+fM48kmSPkGI/t84ah8wHuOZSlSxx+r0fEjHswc7tyr3Swt
PehtkBa0HA8rC9WzAC3sC8fRHi9xL0LIENoxyPV8fIxpVaQ//KYU1OO50SxAoaRQ
I7takUETVU+T+zCyJro17V/DqGmk4V3oEaNnHHyby5oBKEDaJXcvVqbMD/Hz/52P
GQcxmLh5WnKTaCap+DBGtMmUoLobqdc2DU6HNJyNeZMCU2sDfiPDMwz9UU9mdHtJ
vm0Kdv/IVgijsp8vrhLQP+o34PNlDpf2NfSQdam3Eq+LEdS+aCgld2EBwGRvoCmF
W6voAMYYaznK/lp5A9fPPdBW98r7wlPsfA0Y40WLxq433kDdYVSFY3UR9EBB5vdW
LhPoQ1V6M+dfvk7LVNfsNr81dI0RXZPYuv5M/jOqakdrDDpL6v/A4jIc4sqPO51K
HegbCNe3JiD38XsRfnI9H6xUAvy1F3ncUqbkQtYC0nmDbdTSXjYW7rLB7j+ttxf3
2qYsmiS8cpz6ydvYfU9XkVl1IaWHP1eTyPBD4fCzoavDO0Tgex9iaapqxam+ybNz
aCi/cZsJS88jSOKOupJOxFgX7ELiBMljSdhyiqKhFWXupkq1VdkpKoQma27arlCi
/qfRHNnnzwxYQ6IqNQg4BkvFbzfccPo1CQe3044uo0pKqIsXBdqGXR17vQXp3Sps
Zj5HwLLVaZ9KghrZKh1oM5eJ0z9U12p40/lTbrqLWXIHGmvGwe7Yrk61ZDuBXaMR
Vz1eSX+kjYN66SI5zsp3evsHVS13BX/lWJc/JLa0etZMcO3f78ugEwZ9KfETkL3h
BFcbPczaL8YqDmAg7kFsAslLgr5UgqjPE8tSUBg8n00HDzZuG3aj7JYmkfIcjmRL
KQOrM7qm8mGnh5D9rLOs9vvr0jKbWF+Zn+EkOx8dWxDgfCdarx6pG0iuOj8LZM1r
MVcLHKPCMeMnKKC71sJ2qMtk5P5fKjkqbkgQP1ScBavBgw7Tsiy3zz6OBsvg7imO
WWwjGInKmXgE7Loif4IlHsq4EGj1Eve40GnG/oCBVGGnvUsAiDkgdzq8kE9rUDN/
VKb1Xs22MW+mNYyP8ksfeFIxw1oxgXhYpRV8YKJu++jEfm2LodyjnUPvUaWyjXT9
CagtGqJs6/i/uWDZGSC4+JQYidqbFYTQeNtU8WfhUzSlxhxmB5oo6+p19xcvu6cc
vB1nRHJq0xzkY60UC/QBZ3xRHC9FYkVSr0aIXuh9+Qv9dCkcl5E3+Vg++HaKRDnY
apbf6wwI8dZBE7VzD3cpaL/tUsMjdafwmgS2YqnrmrXiIjApLWkMhhuORXt0ypWY
u0ifAoP8m4eqlii5+QyrbLa4yF4jpwqyu8yeNRTBOPrOKQNuM2XnVlOpTZ2rID08
rtMDZDfXMqyMdWH1ZtSoTkyjwPvfDrjaze1gsYS/ETfquGa7Yti8H/X0RDNUBtor
Z3KFQ9LjJdlMCw7Yfa4sFFcCOy1iCwGrdXJ7kVoiwY5YieEgw7hxPu8CzJdvM7B7
RC5nPvDMHOv4Wyv070iYQOfFuBOKctn5gusOnhHHybaK98eezxCUvXUzgyE5Y/bG
Bjve1cJwgP672POUkv6tIvIdR5b4DA48LajGlyvzWLfEXTL6aQFQR36epdkNpB+H
7MRnwfSTMC8BppWVcOA0Hzljz5Vwm8SO8+OqfBfTWxulJgRl2u+EfhGq44zs/VcE
MiGeTehj8jndJMqSnscx58SusqDgHJ7XNurqygPfyHlue8wvKsbdt/2zvLNRm4r6
zSx3H8UEu9JbSr0jZMkINpKNzkUdp0dD/0HdX9cmtlMZkau4pyDljVmAGhCfqm8I
1N27QJDnf03ue11eV+4yqJHxzE3QPtlVrb/ek+y+XBpnU+FQc+iBtW8Um36fsD4A
MnG98ouO12TfqB+pYMrMDteXFpk3qyZlwNAjfAJpgG2nGeeowCLIU3qYHZdnvUhk
t6TUy19aDv0MszSr+eWOfTNDX9jCermOtfKssmgcwcsqvnqrF4S0M5p+aQezQ43i
a8OBD0zjLIdMPOKX8y6Lt64ynvPDYiFeMXd5ZODL6Bcj6eF0npbwKW0f07pGE0Ag
+UKHRVVVezK371lT3TBGGgkE3EfnqiI6KWmZkHYgDI+nndOQnmQXvaSsQWL7UsiO
Kmt/9maeQKAMvQQMHIWmdmLkYJiyCup8fYZYKGyw2CbusnQgvq5V4+bC6/FPVkYJ
el8tfhl+uGZQ5gM7EXNa58QUTBd+gWSswowiKILwmFxe0txU1W4HpgrTCHr9wqyf
zIxGe5J/p63amcf/PgU407HytB3CJqD2MnHnBkrOxffwM66ohSnyNFiRV81BE/Ci
r5ecvr/CRVYq8vghfk6vHefDFaC0P+moji6iCTKPQTfTkXNAswxbG8TcHgJoERNh
0Gr2vpst2tvpzMVy86LBAK2/czrPMevf+qabZ6jENR4eFp1mGq2swdtffV/rZBEP
s6o+6UALEtgBcIOcxE4S8aF/BlZugKzl1YBMgu2OUXsLTt7Kn0Uwgm4TIIvB7syz
XOMb/nOvUbhhLU+ezreX+uHKZR2UJl6bCE0P7iIR7ijmAfRd5MncEaz/f4A5zpeA
ZKbUc+lMRpg002BxXINSPd4VmmvvIh33D3FNvLW8mNaFVesCW6dcDPtP1jO3x+Ke
iSgxk+UaBNfg1GMcPKlKDImRr8AU/kOw0wiHK091g0QxhSDXVC5xd3rv4QSRP+4e
EqQl6kFeU3XyJfx8jwWPLh9WbcwlSQCWWsetwNhtMUruCkh0fGSS+ruFYan4aXYe
RJ6+8UEJi/HT/Sa3YJLXX35xoyexiOZx7WHhaw/dR4FLaiZ1W101AGgvQCNWCsMa
v4qCtmtqI1zo/qDYxECTV6cT6krbqASMA9b2agSeFD5LePVgziAnf3w4Jr8Ps0cq
zRv1leUnM2N5dalWEbCSYeLgM3uJmbEFi7HAvW8/VG0J0OzXbJ70sQAKNl4Uxt+K
C0WUeFGLA/R7je89lbxnkk7oFi3pqrU41nJT17UGndC82f/j7BNsRVxIs7wyP+MV
hzs4u2NX3yBdD0JJT9GA3N6m21KbSEsJdAU/ov4iW4NKwzyV7NOegedLsf4+t4H0
6eQoK52HX2+3vnL58p7i2nV7DaDmeSYZXKOq/g+M8ro1gDyqLZ7P65YxPeikuRKV
xCtHRAuuQf5LIC6b48LS6RzT2lf19CNltztUsisJIrgMY/nW+zPlhkgbTgsSksFD
X51ImcerKSrmg7fUrSaQ8PjkIERp5JphgtACVcsO7W664/Si3cg6Ak8UuRdbo1b1
DnVDA0u4tJqivN06iZ1XCdrkEkXEBkI35TkAA8lbhY9D6QygFZPxiVyabJEFhh26
vYQ2pf77bSJCJ+tZ8yX5GdivigyDma79xDATcbCbMT2gjFaxcGPosnVHxXrQmkp5
60Y+SjammR1DSqNtyBJeWVGBvRisy7TEWRKuNJ0Lv40bFDwQ40Yn59oIo+CkR7dv
an7iPbzJJSX/jNG+twEMHb6BJNImM3fJiug4eXg/sm+3RkIcisysKzr6K6yCQalH
KZF/boNW/HRVGMsKTa77HHKq9vwU9s8ylEC8+Ium/0mlc2J8sdwARTr2/b/rFAyd
itHoMgpEOYGhmuYctSHDfHWPdLzB6gQlmdwWzsHlLt82mSk96Nm/YOp3E/IDkXkn
pJGCDRBtivABN6ODjgv7q6G0kL4s1ro13QlkTk4ghxdM8oIjG+G4nEnP8uB9HuOE
6yo7K3LR+VjxI67hxb6RmkugNTZb411QJI8DQMH7ftPOLFqVQ6fIJhqoSL1bHhSg
LZPScVf2DPkZ4GLdXTbwwrTSRh1/M8G3RNl3Pc4jsksNaHig5T61HLml4A0yw/EP
m9S4aEIxESARwtBPhMZ1y4anW/chvlMqO3jjntlXXkLWlGG26jteffPnrnHiOle0
tJNUguDrk/zAXeL570typD+tquC6Y+WFkb/8crTG9aELl3xgQdpf5hv5CiXyMcLx
60Z2n+zucYOhXMVO7Z+r76TWwnGkpwMSQ11RpuJwQadzUAGbaNz9/ImkSfXPfdQQ
qQMcOHCTTL60+hqk1uw2zINx3RymTPUHya1ZGz1JIdP7GfuqJSShxYC9UtXYaj+k
+XXItKcb4yDBMVzsz9oX/z9qlZ1/Hc33IP21RaFAbAmWRrPK8DRhZ0J6aahKDYY3
umvyfQEPjFFdvfcR4Y5wZp9/6b47kxcVqO79HhKLy2PqJI1x/p1m/hz/uSTajMdO
l5fWfewiewGxYuaDvsc71Ypk4f60Vp0zvsRUOZH+xl5fwgqUBdmnAWuGKyHsN6mG
ypP8WgsjPdmMYC4kjzI4LlCoZDTCWm+IHcaLl2dmcX1aXnKCsePTICBmO2egBNj6
B8OdnhdTImlqk7g0lPL1CPJs0J4UucqoWexPHjibtN2ve2w36T7MyJ0N2D+sq3bE
2lqH2aCpoa2W56hK8XKRlCPNsh9i/SDTQ69GLf40HzV8TTjxtq7cA+aHQi6f7PfL
23Wto5sU3FdHHCzSwNS1gn3bSXmvng+bdBPyhDA10Wcf9dl99tV7amzZ0frk2oRi
jR2h6Wkj7zPnrCT1OyTGU4iBxj/i/w+iMEuKNqWS3a6LyYKQbEOSOOpX4fJjHj63
UTO5TkV2L3tBj2lNDrri+4r5jtqOTFJ9uUkwJuUBgPQJCHnwGJVuMOznJE8Y04rX
A9v7FFUM9z5i/2LlOkUQRyGRdeEYM4BhE5hSCpDOf5FS6XCoaK8kqbpS8mMIuQKR
Nf4bSGdiKW7yzEHq8tfrIMHNXuWD7v61t6Jko2iFEQpezBEkIhY/e/ckVfnUEI94
yogk3doHxEaixvAc3xVfK24ZsgxPVpndWbB0M1UBHLYnsAnoBLIQcJ54EZYCcuBb
jWddmP+CU3zaQ7JZGnvh2UM4hVL/Otypc0MUf7yr1lIlmyPloTNYsSTo4RGdkz+n
ACH6OP0uFEdptZrSTz1Q3SMzJpk/xwrD95vfA5Flo9HyWh0Kmrz7IPqhvjRWQTKl
TOxRUfywYXjK78TieEye0iIcfgZYOkYzOQHTiB6+gZJOC9TOUTXwJAiMqhkSzUh6
vjearTj/91Ot6D+EaASad6VDCP3BhQ2r0U0aRZ6q83b/2MeiJlS0panUZaVGRJPw
Mnc22GsnnzmiPzo+O/RZORAYzmsyXLDV8FYYvNJ0a0/cSpNsXUPuDZDG90VQJUro
aSGd8IqvfmxjoOdeulKJNul1hOwpBF7ibal/uUHpPnObPJSNCeQHZHNcUisfPSNl
WRweoKVO/p600eya9+KYOuFm/t3j/XrK4BdDxXZujWYBW3IUQc8eWoHUfuGRRSNA
z+29Z0x2oBxuBYy0wNEYifw0jHWlP0xHQEwdrkQxwidcEm6VgZ87E31+1Q9tkNRo
ZMEr1dtfg9nKZoeNp9vCF62H2c2jYZFDtRkau/obau0dlqzU9/pP4IELBlsNc5Fo
IkXfgjQDGppLg+tDn7fjLKTr2J6iPFPL29diw4ZSdG4WS9Z2DKweRawERr5qk8zx
LVTOCHpsRiVUNezdFyd4xKHY0FlBt8vijKjXvVtEm+gnP57HAZgvxr0r3n5KF8YM
F4Fhy4TBEfzAMw5l15EFEPI7Vhky0SX9MV94J5KihBVAYF9MYkWRe+/BAyxfaEwg
LBAPszcMNyqW8h0PyfGw5heS99aiNEsZLeB0X3IXV3Ki+arQcaYnPaznjVATNS36
BLXhSa4DbEcQqNKmwFmVAI+XZGlbIDxNPMGNhPa68JzoMHxCwENQRYsSkhSTEnz1
IDZXKUVYEUj3BxLXRhYSC0ZlH0az6Dr2jcbcRsfeWuY0xOG+B3rGyqdq8rRFdbwf
8eRsgGtU3FbVohISfbLW8Z97CR81738nixraJvkjtSW0BV+IstUlarwUz6/VAyiX
s+bbgIvy5UoqgFhpssJkgFRmP84cLvlK9W9uCuzTmV/uU/xBfn1w0zlIPI9T8ysw
qOo2u/qColsuYC5jQnULK161RiWcagmFh1ZcbM/pkcmlEQYUt4XW6Itm1EBe8u3L
3inb3TUE+HHXcTm5lSEE2KDcwFaA7gRP8DGbENvF6v1Pf7f0wjZc4mPutyg/vcto
XyrYZ9OW7lol9xBxrwSjo4I5QD/QFqaUqArrkxt6Shc5k14pxSwTWxydoCq66XW2
cR+x9f3DXRsoGYLOWQUKbBVDcQyxaq6YgLaZMwViE6J6tMN1mUrdEd7YzWOl3N/w
KlRuzXWj2eEjVIqW46fiAdr1Ofe97D73oJ2Ml2SNRlFskEehpX+ChBhq7RBTXLnA
qh9vge/lyGs+p7+9K+cYDwpRpYab6u+KrUWHErydEoIe+ODjsVTG7hzalOSUJJBj
vIjnkVtnYVUhlM2vQLPOl0yfsI/Z0O5aPBWlrIM+Ic4Xs7siFZVeZT93eqVIlLft
GW11T43+m8mCfMhXCgF2GKWOGe31ecIlOONScw4HvFyQsUFgQUBsBYFRV9HUuNfZ
hdj3YicnhwaUCAllwqhiXMqaCpCz/xdg6nA9/3h6leuQEf2qiAWCY71ecqyiuQUv
V28QbFXylAGrRJA+tqymPoGctb18fJXMBZG4NLikTy4b2rXwofKCeZ0MAi1UIx1+
Szq1H4bpdRFLFnB09plxMhYSHTE/ZUtuis/PZ4uJ/dhsaj02n7fHQRZVOQlNgyOK
SZ/h4F2uSntoh6jLJSawqpVWzxxZ0N4EP3V7ovl++ccLSSbpop2jvfNRttsDEmkY
d3NdPp4skx8KE6swzgxrDg1T6D0WscMRIFIcJg6mnDWkRcUmQHjbWDDcc7ANB6e6
a2XgyUEwWajgZAipQPnLubPlpRozpGZ4SZv/HNsUkiqI6Zeqx3MUHsfotQkmGeup
3UR39W3VT38ErAY2W71wdYV9hGnKpYl1E0K3+EeWsnfb3g2TJn2+yqId7GQ4+uee
LdN6EkcSCOg1iYQy748SgjGbqQWRB+29zmGCaSCk3D0OdvL/Zpl938f8KLkB5esV
6UqwUbO41amWHi3M3WJKQ7L2thHx/YpXEZV1g2PSqcL0xLVRrlmT38ezHJgg86tp
8EKelnqrpcKU65b6V2V2jUb9qZQzS9HZCbXBOs+rMW/no3ld5WBwvG1yrqBAsF2m
PoffbnEkSMBlIqUuns/KkNU90+eWX2Dz6Dlic2W7FNZOAcsO8kbqtP4oP8fNNi7M
B/+JSO/coqYAsOvToHky+pV+Wg9TnoEaXOXQj6NDxVdOeMQxSPs1o9R+HPbVduDb
K8eVb6Tq1F2zLpQo1oul2AzYcveI902PVjJ+8h6OvLnjiE2rs1VfT3tqSLbeDTmu
jAUOHsZon2xqpAO7TUrP4O0pF1+JVPl/HhMY0OaE93+5q7xhX7S7GNA849maALj5
uZetyikm8GbNA73b8HaPDk/WWiURpAKh6sxeS3mLmOn6DBvZNbNVqXK3obgaLrf5
SJ4Y0+46ZAgtLq3XqDqluny6/ugUAuoaHXLsTPNJFsYC0bPGqABK8C9twEtBILGK
qX0I6r04JuZNME6wBNCfv48hwx75OjvA8998W6vvSmjjQWhbjvcHc8TqmpXq4FSI
wKrnSrryqF1xBT2m69OexrB+i08YjTS4sqGCfKecttNfRF5uURApQCjzyQHcwguK
5+V4bB2BiuQBmePgWVMI19w26QC3R3dAGHjT5daabXkzYsibAAYbLRR6HzW4dX9o
ZhiB9jPxNjtIUy5l/tA53TBeLXag1WXOkkaC0VcYQJc5USd4I63L84T4a2jKURpe
gp+4UG1iRDofrvhA2d30N2Ecumi3RWgwWHcFEtOkdxgUFOy1V5oujRUwwuCLwk2k
H133Qak0ZjUkryt6jl2wDCICa+gAbzO8rrWnxYFINQXmMy97CA1XP3AEBaVVgi88
CDUN+daynKsSIWRjtJjAaCbRwhyHvcx8TkrSTFH19N9GGgPwZTW5QhRfsXyHf8hO
Hxl6PKQwa9fZm9vJEwOZogZmMr506vM0/C1MyG7RHjjt3CvNtR4cddUKOkytpAF7
Ba8yA2cGw2YPqiEZixHXTfQi6wocZddk5a9pB1a4yHvIAIAHe6HYU5aJ5spmnmky
Xn1ZM44NbiGxEKX9WMEvVODP9JPNkjT/5r5STjp7CYK4SgGnpd6hfxSOr3JLBr2b
L+nkqbs1zuhLZgO7W2fyw/LhJE6jW4XB3K/sN8PHt37CtqZSRyqJGOwHH+OQ+SRo
MpQ9WAs/Xty7wZG3fKfxyFhp5oJWB4do8M/T9JT90+t8TtPLQbaqEDYvBaNO6qXT
pamLBDJgtKd4C/BYY84whoa4oKXEizqcynBoWEMDdgZ6XhkZ8y/Qi2q7a2DJSSox
PuiDkFdNNVcfYA+qYH4uVA==
`protect end_protected