<<<<<<< HEAD:flexrio_deps/PkgFlexRioAxiStream.vhd
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4128 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
9dKN2lpiqz5lCmPQNhR1VpIaRZWE3AoMDCwbh18rWZdSQWq04pT9JDz+oHfriK+P
B5Jr8tiJUbTR7y5GLNIuETU5nrvXXt1EnEgNrwn3FZMpuIQABhL85XHQ5QgtJoOa
H68wqcpMHKbsGtk4rzpZZPqAJySGIx6hc8fclpDO5u9M00g1Hehv9oa4M41Jrj2a
bVmRPHs5jHd/uIGc65yz/CBFZlU8R54GW7BJ1w32JgGT5vN9T8JM36kIiYhOWRfE
jrp3G2G5Ilp65TuAr+KeVNVGETea3GgkniavlMjAE7e5/K45K5Q1oQ5wGhfAfZuT
YJfnr7owBrhlkZSeZlk78RRxZvGrtYIzumvdShMLxv2QUSH6uJsgEhsamn4TEjVj
jNiCcJOn5Br+Y9hbJk4JJlnBqgn05BM2twz+xqrlyrq+vlQkrvd7MWQJFnYnMNCQ
glkBnZ+B2ZM0dr2jl8fGo3sHcX21bW+QwJzuxBSWG821Wql8UDGdrC8yJv2voBTJ
DtZTPCoKRbrYji6PPqE2FgwryAb9U+vOGA6SESkd9vpHGDT3KHa1OmoFwQwgKPnZ
gN9W13BtqyxlBYDcFsBkBtrWwtSittoSUYphBCRmxVpvUtBgQXbEuI1JEGZWcDwO
z3FbwhccsS4SyXcFjCG9jFEyP+4c5eekKzZKCVz2nKXotvrHix7wfI+wYR2Z8rLW
AGr19VCnYX8y4kIJRaqoCbLyU9eo4pGG3X37N7A56ieyLtNNiwb/xceUXkxzhmqR
Apgu+hNHxHyVsV6+wfwnIC4zxo9/5FkBkpzDqtz7V4mlfljRM1zdf40mapU1Cod7
At8LouZW+oAX2zRVxJNAv7ShN46dw1F1SIlpuSH6p7XhlaYOcKnpuSvz3VD6CcH6
AXgAIhVS4RdX9An3VC76jB+Ig24ta6AMN6hyBj/NFcInhIp7JKde1QsEHMN1Sygm
lmfW/4zAlFouA0qKILzhbqq975RGV3P7M+yL0nGON8s/giDXbkctrWBsT0w3Q26e
rer1XOCj//6Fibc8vQvICT1Y6La7IY09NQSrgOjOE41DDKVUqNO547LVk66cMQRX
wtBb9+6sHhldoRMJWQDBq10oWSMQnl1gI2t0x/MRhGkkIlHHTskUNjaKdUvmoaYJ
AtaJLVN4gMcmnQ+q55DMJCJ687X+wipkZ2jMTdgjGzJRXXnkafM5TNTmZ3II5tpW
LsZn4wt7fRwG2WksQDZ8di7GD21vfsdsj7VUkaqoMK32G2M1IzYaltsA+LPk/ART
8GGpvgsTwRc4hOXliY5YMRs52t8Rd723lJ6BWAM5Vr5q/7xWO9ndseElkoomtyfQ
ExHTu6mjj3WJeDEbACrAfwsO91/ryJR5A5tMJo3tcRftyi7WCzHdEYJZ0etJ8fUm
BzQZ4HVKfJ4TnJn0DPI1y55ffUVoQZagzZ0+/e+RSDHv5omy64cnICozGjO/Wv+c
vp/z4WNRodLG/MAqjTlW3RRTMAgL94esuvNhYimDktRLr/nUE5LDsKPkdVxO9ySN
MkP4Csd24IS+45mUN4f1T8d7yWgJ219rZrQp04t8txbZb5RZs5xi952yGjSH5wt0
EUyyXPPEuy5TL8kBniBBWLZDHfXo7qF+P4bvndIAha88/c5UZOPCnupVTVNk8fyj
owhFPtfZcLodYdLnqA/gyIrzlNAXfymCVu30jRJHxu2FR1GMIlMlmyfw1MkorlT7
b2UzQTnmqtZHBnqHLRQ+Tud7/RTyBhQ9uVYFQOA1F1kIF+2huS6pi/PSda+24z8O
4amn+ov+iKmFKcBYA3T56FnlGTTuuupkv1JsSg74s/esf50lJ+AEpG7pV9/iNxBa
61YJ2yhfLYwU5xvDvDOgQTKmYQQy8cs1GnqWfoXLjnGbgTpd38KmdtcYgLHR6HyR
ZC3OzNqKuOXOVG8q93qmJGin/yWhuDqSg7G06E51zTwI5u2hI07CremezJ4oKDRO
lfHxftN1IWEM1UhByAj/eyW68eG4xAZXzfjKj945/Q+WGJ/MRskXSlQQNpIJD8o8
xHtdkDZn9n1lHQfmHR1L0vEwdPSiw3rrfWrV5fuB8ZpeN7YFlFawolDnz3bqfh4d
gfCS73/YPKXp7fE68LB+pEhp2ca6jkPHK8l9q9NcHwDvmkGNi0JuRvXLJz07OAXP
0yu+bxHt0iidWMMyzlg4ONOlSveSDO28zPM7DO7LbDasBGNsjHN/1sKxgBkoNKfO
aHfNbnvj2gQAvvxEE/VLj10IBe2tEKcvVPHat7rAEq8jwc3p9J0LIs77fPIiULnC
B9Aj7KOvHKwWHS3H+mJBu2LVJg91SyOMEXrkyXP9ejPj69CBz5d07kiMnlSDX6p+
J8YZG151nfi3U/+KD0/+B7JpbqJL6XSm10ene+TfNJSLcAj13xg9B+w0pg3GnrxO
iqOivgrG+T42je1UFO0SEEoD2Bm0WiSEKVtsStT/eoJ8hLaYy7Pp8FKWvZ/EODNH
uBgx7iS5QWIGY9i8Ff1BYBWRXWzwZF4FBkpjXFwb/geCJXYMjzfpR4AYzbZ4j/4u
36A1ufLuWGT6gez3RLBM2DXbOfo1knSjpM52d88ss+y0u27ddK5cIe3c2uuiufwo
j4Cg1w379kAuQlSluLm8Vkx5peY2Ee45+YGcscpnZQG45/ZFnBkSiaqMOe1KYs7J
qD7AkzqZDPkWYQiGNI/PY7F4k1Ij/Vg6IBWg1sZwifZqVAn3lyFivFgWtbDsdo3L
XSaqk4DOMxTfySmJH328FU1TY8N+y7YK5lXU/p6wTPTnttX/Fv96HOScYfsEV0pm
Tp4OoYOb0s6GseHC5XilWLOSJCiYkJ8BPDTQC0EZGuhIAgf1jyOnI19bbFbXjyP+
oN1e4pPpUtyL/HiWYkUfhrBNQZS+QdoHBN/PtBRoSAJDxxhxdcrerpF3klvhEfn+
rd3KA4cPpqNtguJ3+KbltJSvt7nmfdCCkcfSCd8CuxnT6mnU0bPstMDVXtVvUE2R
7Hg4iQo5Fy2nzjO7AA4Kvo1NhyOjCaASpBDGfMpe8sVHfFlm1v3lgQ98C4CvPjmi
pD1Od4vWHfh2ByGBh0q4DMUg/8AiLtcUN+YDW1NgbfvWkP2ofJwNdFtvgpm2aJLk
nQxNz92AwRIZPJpYYgLrXGoaLkImrS1rmoAo/f5H1hnG1llX5UtaBFC6Dzx/nqsa
QG7WuTJFqv9jXzoqpnlSj4GPNG/6JQRNQUadO1Tj2Rekdrs4cCO1/NCG0e35aq69
0+GJKLCbZhLN6I91EDCd05z+ETo5D6D8e2WOzqzA3c5WdyPR6JKVP063Wdd2GlFl
X1NNro8Z5J/DD9upHuSzZ6JX4kVVgC4jGDxZu5etl/ieNe/mo+6Zcd4OQ12Oer9l
KjgnidUacQK/gh6q6EvouCfMgWScGr1216FFfU/LS5BHHf4RjbuipMek80BJyuvV
lLxx4vy3SIJsqcPkLzihvN6ehpjuzVS5wqLo07UiDV2Bvl/uWMNRR95JiJKNV+fz
8tr0jEufcQy5Uk6RZ6enZQ/qQRse+S8lHwHWtLo0OUOFP4GwcACI2axc9Kc6avPx
d3ji7hVbyoL0c36jJuYAz+gmrekf9LixSrN7HhaEn/2QdXYxNzcoMN666cuMr4kg
+F56Kl8njKdHtBX3bHDJV34HtiIOA2IYSIN2SWgVfBI4it1Kn0IPIoeP6goRA8TK
Xuj+LPX90hzkSOq4RthbKatmiocEKsEOVCBY4YhcXDIlC2E5ou95K3kKW+q184cG
DGkpR8UoJ+nJWSsYIMs9zKNCh9EhZN3iiG7CGK+AO0Ah+wvmNUp99z4tlwF5Cmbp
3pwg7sRAPLTI579G/+7YJj6PRpq+J6VFRfsuLNVmIAQV/vc/iqA+5tLMv947CuTp
bSdqvxFbua0lhsM3fdFhG9Ks0S+dSDlZ8BmDJnstGKb/TPh/EBSG024KInvE23+x
Vs0poO9UnjGiuxyD8Ez/AhCh7x93E81QFCq4ZCNdP1pDlu2RCL5ARFXJGAPs1Jg+
br3Y7jYav5LlBzpT2fhXwkvw43gT92lrCb5w///hwUd+guDPaQhVGQMnAlcp/SkB
p6bbmmOwPb2j7exCP2SSVJdJPbFIXS+CH0iQd76dbVCvgtsBN4HbKp2p16/2TdUl
bQnZSnLKfa/Dh+bjg1GxndOocN5TdPfTSZ9+4mc1DR9p0E1cLV7BPli0/VfFizYO
E1kb9mxlP2rgKeI7nDMkKW0gcAjhjHtGUHDTQMwGwfsxPfrRwj4Cx/gJghbi/6si
3VyM3LYPDeKK/R7uyZIM96J2JWcRsPzmIqzm9EzZ7PYJFfmFcOKHiCNJL3xMUR06
yVO3zS07UP4o/1VLxoQxGLCt6VWFjsJ9LzLIPaKy6rEjmH6lQosCd186cQJaLcXC
NSzZRsVFTTihmTtYWUfj7kbW2bn6LSAxNBJTSyKLewEqZsfnmH93KBIRF2D5Gzru
DS6Ioqrs+L7i+h5O45nu9w4GY5RK0gOR82Opt3rlTYkAI5cY0qrSR5Ne4vB6eCyZ
jHimx7p+HkBDTENDPCnzqEdGmX5Isj3c3W04oRJsPj2zoBCQHfn8o2IAa2rUQFeg
NpWXJCgp7af/CkISHPD93GaF+nDdLxZlRRgbqiPydDj115JfeK6CYeg3QRQnVenO
9jjHIS9V8eoNwEHcdEl1Jrg0SEFV75zvUpBkD6tjEL3kzD92TFvgki0qkta1Uc4W
QRBbLozwoe1a2M5hL5aYYSwDYHG/tEBqaef5DKD959oH//LNdNeV0xhUecmj7kk2
VXNCFcPMrP3TISNY/MFQJaLVth5d6ZQUuCwl31yrQIO7ifO1oIez8nEJuH25T9gX
/Z2+eZwE+PBMMRW5mUoqqNsOyo/Fqpr44lnT1c+lImhpNoJTqtbxEEmfFuxJeN9y
EtOR5VO5T9yTRQH5x4vXAExpcMqc97vf2YIXIaZ1wDAnR6iBvKszUBnmy9gf3nhE
yjak3V3J8X/cxMcFVDFo3kPaRRj/Om+pYexaAidFpVjsFAtz8Mc12cpzM4YD4Tl1
sh7cBW326er1Eu61NY5Gk33uFfJGeWb1G5Tw8oe3BFdWUdxDwhOouAzbpdZ9WClU
GMIntlS9C4ik60ldK/Pup19L3kDGRvAK7ebg6oLhMNxXGVtfnuCa15m9cANBEgDk
5wowKlqSIfzmvMV2hbMnODDUg52mHBaWNPAM2iCOuCGTejBPqB6a8kehsZvtNeIk
i3QOgDnAUUFfBh8BIrRsy9RWJujbVPDZ6brXjo6+Nc7QrDDJLMq/axhlt3wLyKn6
L0DmUH1q26pLhgsRQDDngVTVw8HdKW7YmphcTJ6DB9X1Eji5NavPzvYGvEm6pUD5
=======
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4128 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
oRlhLo7s07tMU+91cKr0qCayMaM7WFQ3ALBbAhCuUrVTHBoAqmg0eRMCbFmMtD39
s0cpe8N3l3vjpobeODaYz/KVZFUYjkWbgiz3AO/ybZshNjUGXlio1/zpopUtxstJ
Pw6biEAvS09iDtUcRajXn4w/4S2AJwW11IlF1uqgpyaGaDdAOAQS1hbDLA51STjd
zOuYHcsxi6up2s6N0Qat/dUWIVJny47IqnnQErGgXs9MfBy01vgN2NatstIDcsYW
4Q8f3YJFRER3fQKnpGUP/ZcYqmZiP80U/u3orPmbB01urzuFSrNDDnFM+Em6Xt6M
rGvv3mXstBk8a9L4+5hO+XZEfxvwsokS65Xnv+XtCk94kgRCC0YnPTP9+B3HXVKs
giv57U3GExLQJTmgssR5jiBMudDh9PbYpQ9TsnLYUeFFUDG10LZQfXDTZ71Mpv3p
BkmpWwDyYUJZXxBEDEcNfs67zW7/AF+jegxDhxE6ZOkP65ktPTPRUOCw/dCxraUl
T4YfqaefLjKDqyM+ysMs0rIsBIFe+LpIz+rgEEV8Z+MpOertBV0nzfxHckH80MT4
JuSHbbUVbB7MAcJl2ffU8uLwTGW7Y5H92BZ9S+xrdJXDBtG9qhBNJUGawL+LdNRg
NP2dApfeDZ0xq4hqwuTOHfwpqsNptPJ+AardxT5et3qGbhHsZBWngMI/FOQVanAK
nM8jSkdem/3QWOaTJ6PSJaQhtC0CfOimvEfYrKEkAxk5vInq9/hgHJzQg+bAwbAf
GrzORiA+Difm7IsBbesTlFLMSM0HTrgqhGPWFjnNNK1DWWcLKBD0U/nGsDYG/ZGu
NW4jpufHSN9xIE82975ahOdTWyGpJdJ1UiWD+ru+PsCzHdmcaEOOa2ZEbvv40tyy
9vMRuJljfyh7sCQ/tVGoZGKYLhAwQpidcTKsayMwJJWh98JyqPb/RjZQRxBxrlMU
+DOlkO2QG8s38vJ0X+rbWyAEco7ko8Cq3fVXnqgSNezaBGysquFINJVM+BXHdHu8
eDL1lDgJaX8D6AQKed81X0IVxv8KIsj5PlDjqHVp1G6tmIXfxKXUayKl4hpNZufz
420Mnme+OB2cMtRbRv6SI6yaGMIOpjMxXuiUjDd2gA5JGFGW3k1OGhW7oPCYhB/V
s6/jOLkAwderz31jdMjBzpGDQ5v8WzPP9NNQqvya5JRr5qpEN/rTRnypNJlz276W
Anh5++t7TV8OEo/YVtgkG5ZBzZDWBzKZ2n9+UVnkc/v/f+kWWyiwe00ehAKuM0bL
h2nytsSzlBs0hmXfTSXS/1OVbcZX5ABFWZGreu11vtQuWB8zimrn1cVeXYmiXW1a
w4+/HI7Ihfa9uhBGtapbO+SwTFfbwkwTGp2PWVXnxeALJWfeYhwxX+NgpIhq745s
VlCCAxb7IATjBCEIfj4htDpw052PdPNoZIL1LiCiSSHDc6X7utAAXu6cJdcJh8IO
zpn0avUsWai6/6Ii60Mi+CFzqm2q3lzxdDeCFN0wYASR9oMsWQqbh4uDKtHemP8b
gPD2YphBSNuv4KpoqNCpGtF6wGvPW4W3vRDQBpmCQVz+Dz3CbufIO65u/t9/Jpqe
qiEiVGvsA89bvC/LVvU0P6lzoTEBzCZB+2gqjWktM0FHxvWdq+c+g0MChgmaLn1P
yCaCS1Iog89gdRNIQqzAF6+2jk1Nn4G+tvyBV01Dc6wNtsgCEAZ3FATRNj/ob2e2
kH/OJ1wPU+JSwocujlU6gTPyg2CYQAc2e75TdmKR8HbTzthkOARq73KETPAyjRT1
k9eCOa/c3VqQMxEXruWFwVEFj4Je/j8CTyiRv/j+FOTPvDJtA1mi7p7+UzwLM9W6
ofKtF09asF5zaaQ4Uzk+PAkKX8roW2SwE4YR0+cxRmQNYxxsGYDlZVDcD/PL+AkG
VOzGYezuWVVQZHoqlWmfx1YHspSvGe1KoCUBvzfD/KoCqVzv2N61kaM6TlfAZstf
SzSK4w2H0fh475HlZjrpS+X8kmdmKkKY0z6Dz8t/zH0jKDgCKDi9hJpTVsrI4Dh/
UxB0DU4WxURUXIhdqjukxkt6Xf2EJIZbdAMNfiMNScKGHnZuvkD818VO3rm/niaR
AHHWkG3ftYveFNoUmUBxT5JcUCmPnkKKzqAbd2giw0a0JO4MZUjUMIAS8SKTKCwG
E94qUXZCdYKP7jdTEjq+HDtzI5+IpGzAieYt248pK7/sAQfw0ebRXiDI1H+sTd5A
7oDpCKsvpaUyIg8ksCjWBYIEjh2Jow7H7TCdO3sCjl3no7YIlTWMKVvl2hLKhwY6
BJNF+Ld3475oVvtiFpV9NCPXtcKb7gGXMCYtqnVfdmAeIhSmrZ8OoEUBYwkx950Z
p5eZ4RWxpRfynguTG0yDqZ74MUGrpV4rirNOMSojtPfA1zjp5U2028h3rjiELk4v
dd8xA0kEOV7WCdFdbXXRIROS4Ww/tqyLbAvwRk6TXzV0JpBFAWvndS/GDlFDxEJ6
csZ1a9wiJOUIZc2XL1TmRses/M6thlfG7Yg72ZqNZjSFwVENq7qWSX7VV+X98pKR
tIvW0kyJTIG7LFyV8LRnhgMFOL3ewx4svBxC/PTTHkagS7FvFmKQJLLx8cbHgldm
KCM4dBiRHLpjH7DNun9ttRihA8/ZO8CKcdo1mOiwi/fjboTOEMC3SDlg1Ohyo3uQ
Q+X0a9LsmBcleitrRxEVmfOUoRWdwPoRo9Wckwp03oR1Af7XFtliiBLWL+rFS9Xt
UCT6K/X1af8f1lQ+rySt4mXHyJ+/rsLKMYVkVysgP42iPRXsfnKtnW33Xfju5RlV
M/gYM43GB3wyILlUUiW2mLaLHjA1aiU8nnAyw5eJ/f/Gnq8d0dTmSqjfGgkMN5KD
MhzSVYZyuZQ6ILYlXA4S2Q2VhehFylFwesDV5dAef1zLAAVBc5bgXsqGrPdRPeEP
rT9VCVz+zQPowrsY13vrVYES0XeBGNRkN2Mxt7TuHSzGlzvUfmj9pbfqI4YOJTsC
Mc4cH58E5kEvZganKOUbbRCu7IPTgYNvuKwFe7Co1L83nxOuHFC0Yfr2sukT8wTe
ANi9IVo4WIHtHdXjnEbgv7Mxj/VbbfWN3XTzcrVXkArK7UWDBnDtmGey66mRuKJC
RETQ4H+6Yfw2q5+Z6r7c6zA6cSVMcQ1ITFIyBzNAMTh9ci8YxaOC5wkoWKKW/LIo
pXpEuv1fadOxNt4K5zDvks2W89fOSbj32lFxwj4z57km7VWs6DmYQZz68LUVAPJM
zim7FJu9/ADBN5TgEETeFDuyQ1emeednYkifW1sVjFeG0FSLs7mzqSOqHE8Ih3JW
PX3Uow2tvTVzViaOoLKC6+353CXR5E5SzxokXZ0+CKT4jYlmrwKr8o+OrLqGb/UO
Ts2KN623gjBwd9dLy7aTsxQlYrJCOAjadQqNRGjq/tVQH1KQykPBzD41X26w/L4y
hqnljo0u12hjGMC/55NgeGU37VVyUzleK47HEidhqXD7jFKAdBaVpm8tQUDAB3h4
QSgQSkSAix0eLSzQxu1nOGQjtrFhhu0ZdckGKMzgzbCGyt0VPvlrK2/BT6vUna1j
5O8Pb8wm69oYi1Lb9ap9Yq2lB2WWe1lW/g8PsfRgNhggRFvY578acAgOsaO5RFAh
vkBIxS+Z5NG0U6PkSfaLQMfTySIAtBJQpB9GNEtbqmqtyUrxqKRMX1KUXWWjF8ve
hZAHNRGqB+f0+NIt7jcxmnuCEXzZcczYp8BPaSYsOZ3MwbztjeYmdguoze8oQMj5
LtkKSXFVl0qgdt0Bnl0y4wVANuO++rnktIdMa0dKOjtHKzaBkIosG3aJDQ3LQ+/b
LbsecqEqw/tBfdr53RqXIBh3qjyx/TatTkXmec0AA+OOAsjHV8ShZ8Cl/pO6lR3Y
medEUt7AtH8jggWYxrC7bD21ELbQ28dW0OoFSumubnTPgSnUlE31qQ3OgN6ChdNI
5Cn4V5A8zsMb1Sh9WD6oCaToaz2XsiyEE/VbpVjWq7CjAk8aHNbJE8Vu3gaZ5MrT
yafxQK8NBOEP4OQOyaCBJi23h6j1ZZ3RPxICco05e6msephePaotsV7YceWT45tH
stL05bJulerG9A+qGLclKDvWUCrtDJO4Yl+TgmwOdGosrXeaO0xbH+kEpONhQHDN
rmA1VEK8/qYLHjJKVWQva33ajNZblI76At+mSQs1mEXrqNFKRb4v5BRAwjeZjSVc
03paOTi411tJB2IfWWVZk6LCysAWisb+PMi6hGCg4n/2vZfiOLF/LcE71QDEH+a7
FdfCbQiQ53J4g3XAxDBFWVPTHjuGeZrFSpAmn5w6Cyr1bCizB0ME58xWEaxiEeIY
9zdUxe8EbNhtVT586nA3vy6Aa4Ic5GywpbeGymHr4bVm145vjyiNskbVNy0o4nMF
JPJ1mWkEZ3oiJ3jOEtPt1elIwcWWs9CO0nG7NEANObk5hvuSPWSKJdzMHaZorWZo
8qE2j0bU69Vm6dubBH9OKxvaQ/7zYJR4F/0J6Mom1eLaj9v4K5xTygTi0qHG2Qdk
qPunLbcSMWGYJndHLDKqFg7nMbXdY3Ow3wZmYoKdO68Htm6onbEFaZAcyIysLekv
IMPJxvjTH+fLnJO1qASZgjTx0OJLp8VQy7PyCa7CYB9VIRWl8xCIn0J1SKKgiwGg
bvoVjFoYPkycMehSzjNYG6M5I5G8VpTM0cBzwlwh59epqtCr+GRJjMuE+u8ZzTBw
Op8NJYWm+VIaHxC9WnKdN6sgG39unCqAS0I3+yR9KvrBF8Pm5jWRWNLHWc6Sh8PV
LTHwnnsbizNk8ZFYjcnDt5V+J9ftbCuwMO0aQZ4wbEUYvTNKdEHV01E+e8ErMQ6l
96eI+1UMjtuyEJqIzpN/Y1Egxb6O2Rczz6hI7AR7O69ZjvUPKxefxW0evpEtN+FW
RhWkM/cYW1un3NzyLzlBmr1iJH4a1q5FIrngiSCRd2vkZR4EmgJbUHzNTJRaq8LU
pknTNecbaG8dKWBlNCCMKJas1hnfsUv1YrMJEnnF8Xhav7LMqN0RL/qlhAXJ48sq
bXPlHSVaW46u/fC4SoAFU8ICMqE2F64YQ1E/oAzoP6YOjcsL7fvia4auNoUcEHu7
ZY9Aol0uYP1eiohQMerVLcEkbwoqXT/oqdNPxjRgRnjhm4wrB6FuwqCIe3FWJYsW
jCy4klzTBS75VOLU28IhH8ACbBKuITF4gPCXzdwc6p3NbrzwQtp5RaowSdPTObua
a/SIunX3aaT8tg3YguqkbjKbDSZz+0wPjHYtCPK8hsZW9/dzpTZINsntlkCWDCYk
d60eogeOzl0SNMPV8aSvICfL2+qwQeLr9ypOc38TyWQBdvH+IC5CgkLoRqgWVhBo
>>>>>>> 426889eb8ce467b9c9a9f74dd4af433c5046285c:deps/flexrio_deps/PkgFlexRioAxiStream.vhd
`protect end_protected