`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6848 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRu5USVS7579wHpheYeWNqWFqZEm15wTQ436jZJWl2c+D
Htzd7ds2HQDtAIClM39VrZ4FrJekT3UVRl1wR9wXDTuNY7HvRIxNUV7LFZb6IPTU
qrusQW87J+XWxIXEeznL1TvBruHfhdftqTcw5bZS9JYdb9GzoxwiAlZ5dsPi9bvq
mBsF0lEAQsX/OETRpgxCxJB+fiDHJjK31qVXauGqgJRAVBEUqkMD3V8m31T246S2
129P0qCSOj71mmiDkYyKlQGn+OLeFm260OLgee2+Fr7eISD+TiRktjYXIAThqi9j
wvWByxng1v5pJf6I6R+qbPrxaxuiBsyjgP5pbiRBG+XjFXiLlCBwbPG/WGupl8Jb
dGiL92gYaHtSdcSoZ4CYoa/kiirplcccttZ3/qtdcNTgmWBCd6iLq/zFyVYPR3m5
AN0eePlZ9/416zQTQf6l0l1jC3zHWNHVx+rF7zycE71lxouk8GCejiWhYet/dlTY
eVksCaMi0KuuvmNRvpJdc9hM06O7RfIXWMhE7l2HaT/t9KWgyyJ3mGZJdzWqasGC
YQC4y51AX6U+QySqTubGzkacLDyv9dR0kEeJXK6+XMWj7ZqVzx+46Nh48PyTNUvR
+gq0dK5Oe9KPJt8Qdyowj5REZkG3Gasmzq5NKrYkNpbYsvpLWXOFZN4Bk55B/YXV
V/7Tw/m0812x1EnqSoBtlfNE6gi4M03DxE5pz/ootRNf1UFDvI91pGIcdZ+oddQK
vud4GKePzVmz1MM9ph+6QK4STVsC4SqOd2zIt61AMVmSmDP8lhTAxF3/hlDV3GrK
rkwHdOO0s1TkY7jrfW7j6lbV6qJ6bfzOV1Cd1cJkwYeL/qvbEZg+5GXMzi4Y9miq
n2jgDG1kCI8OtZ9qPbgGDmaUK8LEYwhY3oskPjDbr2N1fX9IoGOKQIZaRxRkVEhh
2kDWpfmksGxno9aKBHHbov5iugrF5QRqLsUqyxBRIHVWDZExu7vYfy7Nnk0uS5aI
iWw8iQ2uww++y+ZgHsVCffyirDXdLJGlx/3yaa/P1Ku1/78b7xtAsYksiB468J87
/Mgkl0EymY/omjdZxCBq/H73ZhjoBxvOEIOClTIdLZRcUvOPguMwuO80rgxreEIg
fJZISGkJZQZTY29kTWHY1z2iPg7YdlZNq0UemvL2SEIZ/eIWJxfwS46DWTmwivtj
da3RCazxfQ54o1yZcF8JKoPjllOUMunBu2wl8hfSS8Kz0uNYq810Z1l8PDRnI1AK
4JWwl+5KKxeo6Ae6pj6ebIQKTfx/qgM7Z6qbdlaibKIuQFM2H/o9hHAqdgvhVBvP
cHQf5tujWYj8tBwkemaWxi+iV1S+3Bi1W2EniR7w0wmq1C0f+wi6BQFcT+bNt7gF
TnFy65o3MWnwSfkY5bLNzA/0Z9k5HM/T59Qu06eU1zeVeEef2F8wif7k9A8hsSeI
JTGthveoOG1+9+H8ZeQzEliH3etik5GxeKUifLJAggtJPN1dVX7e1pFOZAnNJztF
lrMA5bkyh5lTXOfJg8mDZize+hbVzdnBUQWCaTVT/DiBLm6mWKI9hI28X030h7Tz
jKhvYab++7idfg6bGV4nRC3PYlhdbxeJczkUOEu0vgqe4cfDhW/ugo29HF4U8tZU
x5i9km3vbIyOXEvuO9DhHFr+HMCKLcDXwEqMNzSk3xW93fezkZbPEIaS+Nt3qntz
gCg53asq+mWtn7149ZN3MOgIJD/NpA8vzubtOEbEmAGfc9IfcThI+DcoODhxI4hP
6surcsnrff761fSH6cy22jccMGwi7MKRC/Vy293afxdWk971cFUpyIRU+itnHKpr
cXWHzbO74n1ZEVBKzcnW041ZkqUJGK3kRPh3V4jkY8NX+s63oQMcyXAkyetjYfx0
Dpmt2gct4/i1bdQCwqESssKk4jbnrRq1ZQtPHLb1LpuV4fXkfHmNMHtihiR2mjdi
qh9om2sFQge00J50vbbOekqP/udRGZI8nNm49cY1S1AZbINOmDF35p14jJcWVp/k
bQezf0xtuwSUx7j+KoJMiWBA7EkSBJJypldHiJRkwgeO9pdZZGsKOg8G7fNVzgCS
xQQtx7pfFNC3tV1nAMtYakboNlbuGLlFTwNTrJSAlzi5OAnRr3K1/9/1NV6UmfU1
cchLy8VgSmDPiF7gkTfFx26H15RuBso0QNkkUGexc2hxg7eqTQ8W/20ywOPfGssV
iERB+x/fM6E367m5tdap+OTYcpJJiBzSLCUICAtcJMrj1Ra3+LV8Co68q858bCaL
kvSOk46iT2Bh5GyYGWIluAITlAgGGaKcPynal2L/kaelcDx7gvoJ+2D1C/q1tqAi
TZMreH/dNZXZlJfS5s9iz5VfA2zwMPRcLge3M/KLDv1y3KIev+igiuuqZTMH76zl
Bad2IyLzKeEuiJnK6QcaRdlRqEhyOyRhbxsTT9eo+vclMKvNOqBMD96A/weusmNa
venIs6hu/GJ3pzz/2xsTxRA8a5crc9n174ITFvHyFtqyxGv4o9GwIU77oWFtJzjt
LhJzgzUgH9pjLcY6ocOBsVzPlQSmfKQnRAxLNn50T8me/2DRNhE0wdGHkav5TKBH
sSd/Cj7ohIu9URJ1+WIk1rQXfL6wNZEB+uU7m1lrU2hi9e9yghi7cetxqqGfN9+d
RsHAJoKXZFLlBp/NBEJqKeUaC6jjhJI4ckWTskzfA/K14BhY2RINcUzEweus03mc
vZfYUkJXVDFpDCdT6WyDnCl0rNynZrc0jYMu0SkSGHPdYmVJXSwAqXRVP9IVdhbm
dsO/hVY2/wBzLalugU0hjwRUATkmNjD5mUqw65Lq/b4LBEswMrBK0wzAc9e9+xxg
iBgUvNkIXFfzAjUXH7HraIAo1Vhi+8K5qIs1Eysg495XGx9197Az1CQ2v9Y3L59/
eXlqF22cxmkd663CrL9l8q/vdfs/mKR2AEJoOg5+fo3PDmLRBD6AqUsTE4kqlvFM
xlgiFsdnJsQY80xtIW9jRBxz+oMvhS2jypRnxJkJo5OgjTC4LLsNuL4/Fpw3P8Oi
MP5p4eEsgpv1r4Ft38z0x0B/MMnNmZWUonwDIn/3A4D0LuG51Oqm3C9ZTh4H52y+
8XQbg34WateU8RP9sBVe7ZY9jaiEbaxROYk7BqoBpwWGc6icPv5oflq1k6KD5tPD
FQt0zToUCv76iHbKftVS2IOHuic/6b1BqypJLVVsxD2IbcbJ++iAgEmFgXe5u4EF
U3dz8WvC/99xjlVSVTXmkXHMuuPoZDwPh3ClFJKdchN23iKZ0y2HqYZDtTb2QID+
LD98bMnybCEaN/3D1o5Nb9TQSWwGpE6GLVMxYGx7wyQvoncMEchSm2xE7TSU8DpB
AlbfSGeabCOtw0Oq8rJdPFfizyMwI28IvDqjVW/SfwWU5PF6yN8jvTG8KMnXO1np
2REvGt/yg2CRNRzYLQP9W7xzBQSrg52Ca94KusqhsMB5nl7PIqNNNPlqAQj0GYU9
pp6W3VPTC33R+065/joke090psn/6ePiJoUzcHUlelKxdu2/1pnUGTysaHFKPfd7
LluInVahcLp8j6jhuBIbgogjO0RH5XcD7E/xYnzis1AzWnJtbuvKA2R0g1O/VHwE
4G79n/oLvug+zRykdprGD4r5yg9hpRQXY59gLNwd+07iQkoQ02aV/gz+IGZKSs1u
gNgOC9Yi/sCPeNwOqSUd2SyeVKE8k8ccT5jjfh8pmGXq8MUqe0mx5vfNoEoI325c
1pu6og1DRWps/rQ+nuKeNb0/2UxZA9WA43g1pqztS7Fak5BvUe5R/kVZkpS9wZ7C
Wy6Wh2ncxETX56JaXGUKPuObZNvjHBANJdo2TKO3m5G9Jnj8qwn9B3h83btat940
jiUjPv/nJf5WZ37EpFtpt5RJ/n0vKq0po7/M6jXXpnzShdsz6NkURA5446GGkPZE
FFAYIGgCbjZg+GkjzMLFQmcAjVED9fg/3tYxdX6eFrnyOvNbp0j4v5fpDNuvua9V
tm415wjb+ZLr0c8S3FEAA0taDIgFFrAEqhMtAkvPveqpRG47zxtZhug8rnG01xcm
WeTNTYOk/Jbc3gCmmgEnGYF6IGlfND6mEM/CMBxevZ+k+LSw1MCvCBYehM1GFEgF
7WRTRsXFa8Ti/B1JWRKwyvn3ku/iAf2jSiPv6Gulrq2RevNkggor0XCQmrpEs+Si
NbFn6/iYBlsMXQwyd34YcpSs4r3lDOkqOAm3DQRshRLArUkxCB6FV7BC4SNTop1n
0EZ7FmQWkVK12geBHajqBOX0+XEL8ovzbOXV7tVjR4T8n9Rw7WIvL+mUK8G3zz/K
Uzr4OfhDuzzk0VtOHAGIsAoO4LV7fM7B0ABO81uEwIpHvHo4nKJJqgA043OLyBXK
21a7BIEQ0yYGZF8gFJw0CdKz6fAJHN+A5cBDY+I/kxIgmCItW3rGBhyI4+U8qxX/
R9LiGSDFSRDWbMQg94Y8JNH58kFpRRu9jYYWCInFTacd0f5y0uQF4u+r7NTGh9oI
WhqODKD/gOH8kOL0pU6POeUL+j40BY04RuX3eK51oUJ3GWWNsRpTm0tprf9ujMfx
0HdSpcdSfQeHRvro9LQnQKo/bJ65tPb4C6702wsZYo0R+Qch+wCaC4f/j+lRlx3w
56d2ufWbuxrmIPNDjDC8gzZXZZD2Vla1aB2lUCCJJp/cpCwMTSWKHp/Oh6ZZ863e
U11U/Cb9Kh9MfFZ1T1CxhzXg6gj+nXhxeE2OvZhmoNDYISIcsHkpDLSBFcRDpMMh
3su6QAMpqYVamFtnoADS1KTV4yZZdZK6eoO8QBDLd9Q/q2Rh+q/w5I0lj3WjuRwc
5ZuSAgvfGJCkOEeca3gAJJD0BQpO9cZFLyJD5BMQsDTG9mIqCNZCEUPLoAjiE4jX
GB5ngjCNqWE+4Pu62ajYWUR5R9uxx3ZXW0otkVB8fnlsyQtgRfGcz9OYweTSAWUK
GCZaWMu6wcMXBVLKLcd3Fau7gi6oKvjrdK5IVIwcOa3iF/wIRdQf2dh/Zj2DjhrG
VGeXUknWrtTHCRgJTMKfqENWFuag1AqYZYYY4J5+aEy8yapF6/FM1a6Suth+IcaH
qK2/LJaaLRIyJot1mZLTnWH0rAaWYJ6UFhF+eg2pZNOfozmymAqgt8WkJUoX+L2N
e+kG4Tkxxz6ADhgJrBgKbbKUfltyd5W9UoTyTdsU/OaCWx3zz87iPrcEFPUFFj6r
jfsA/xjGcraO+maz0EnYUqs5RLkJakZXJxOIabj1Gl7y5/Mw/ZT2DBINoKFMvup/
m56rkHqPxOjO/kTUtxvP6khkB2qgiDLql3EJN2iBtxB8AvfXGJH4PQ6UWPOM7P+s
3bMG4oB/mqQu74VmaCGnM8lQwg5vbbXCjE1usEwo8Qqr1T3l+e6TOXUjY+F26Jup
UPGfQdSjd+uWYXH1XFXpGqaQXeUXgDeJREITz50b7s8s7xhuT23/mNHFzZqebnL6
lJlHdOjYCQFoeccRoC61YJgY1m6+OiATwL3ZIG3t/vkSrwnCg7xXEh4Obxx2vTVW
q5ph/J0Voz+4tDk1vm9j2fYGQdYAme0qBXXgfrxWXbbDrghlRvfabUwpiNNXHMT7
ZlUcR/VcC8172gFb8IOfm8HZR5ZfOsn+htKiG0eZR43cpL0Iv5kcD1d0lYfgdCL+
tfT2MMOvoZLrtWpZj9GFyYRJr49yqz5CaZ9atlqY9/RDhXdecIgM2PUN3OF5AsWi
ss95SPPQB5WsyvB3taxfU+Mlw5NPnF8LhF/dS/KttQ6bQ5kPhpRx3LjZVb8cUQG6
Z3NZXf809Jz9lHexaOLhfp65lGLV4JuWdWyeFwlWp/GmMuErG9XqK1HVsqK7CWll
aV/Lr8UadNliGGNRYQJe30havezHJ6lWA2RULOJMumGb3+QSM4vCScWkOsAtw2Sj
ZF7vZAE9BduLI1lpWREgKF2DfKTCn35woox6/Y98MCFiRuXq1O+zhbgahyVP45q6
4ssEk2UM8D/lXW2K95exyGmfLWojEAM/szvsoDNFVbQYxqFt2+vwg9NvN9ECushp
4uTYgcla2pJGzpWrB0wJ6bXrd6SY5JhsHFlY89G+B7cbqDHo09fStUTkCW65ox+D
NPX2yaeC6am7gPboq0KGQjDXY1hgW7zMVadA8WzCpLKy9Ph9uzKWCBQB3G97+ur6
jSsTNshmvCjjGa6NovyJWGDgaLt4dWs6kXSVG14WIURicYny5lYgEt1Cyc5X58DV
0GVWWNyq2UnFLBG5uKPaq44A0dk+fcoW5B8Z+b7yAEsf1HhhqNuYUrHLvk3i5Zvl
FcJAQix4muN/IPqvPACqg8xjEWQIjWJkCscx+aa5/xLaJABbdZ/hje7WkmLl0yPB
IiwpNI5uFV5/JHIpeJNqCUXnkMB0Vaw6ZTRAGLX8ry7pO0hGSszgW09KvOywGug4
0sgfSdbscz0znGi4FeGXvk5dlYQY7bTYfvrAwhvEbAadrl2i+mqvt3L9a4qEeRD8
ZM1g18McN6xDuOmnrb+t0co7RUMDs8ZavYynAJcYhrHG1ns7yiB6crGDX7YBBA9g
pzJ02pXVHCsAAnpbaDGb/aLJr+JSm2k+SnpskgVvuXChxPVSAuR7Y00+yDFPaAQP
wr73H3Q3AYsy8mZgGsUmZdpPMmkXLkRckleQu0IeK72gRqnBR5z1URTeg9AZiDUh
OTFRI5i7Ux/AUNTNnq95CvgsPigivpkfh1VlSbFBqh4L07FEytl1StuIjeiBfOhb
7omDQODaefSIKSTVj5CLlxHs6SlNESJGsq05brUMd+7Uvfq9jY3xcrgW92ca3QkU
rrZ3f6BFpOV7mqAxyZhvG3CglSp52XKLP0MsdVnJExy8/ubulzFWj0ktL2joSL6S
JBJOHbe50e/S6cec+HTbaoGNRL7isUusGBHZNzyAiaMiQaXQ7QXPYY0PgNkGu5K7
zU4yj9VfqBRMLL9rDIx8NoxCMqvW1ZvMOX2xxmhAV20tqrY9U462wuT+5C9TUD/J
k7cRQsjknzX9Ho996nbDUszlNYOlGVkDyqkdO5DzEntM7yPwqCdEjsCb99X7B+mx
3p3A5DeoR3AWFgHiVHoBeNDYzOaJbflzUa5VNpYkWo6tfmZzcNjWdTYMIouovHtz
EIH/untWxwJt+zCNq2zdR2fLHp0sAPsgSvxZ0QeMpzUMjGtab1zkJhCQRK8EPt8/
rWJNNGVXjEt4jaFULVUhoh8tL0zvaVTqdnQ1TKnNn+sg0/3Lhfoph0M0SF9nfxf3
osMIfUzmuq1NX0J8JPq0PauAXDmvrmpEmjzElxiBZDb2m3JUvToNq5srCSXZZIaA
LlPuaysLN9YFK91sEyCqIXcjQeIZpEQulfR9PALfNlJNSMvg3aKqKfikQtK8g6/L
WEuQVyF+HSNaPeEup/7C6cIWqHg9vbD9n4GCJRk34kyP2TbuoguSHGkuOv92MKbh
VmA7eLdgncS7mi6wdGcCREQC4uZznP1nolIE0TMMbqRc3KZq6kGzc3TyXZqUa+mJ
Au3zQ+0g3+E8wxWiIwW1H7U0Ivrr/2g0KilMWQg+U7eyDSXpWvBsrNvDSGyBLMHd
AWz54c8SrK+pmHYIZOSqyuGOp1b4uyzFcy5HQjD1fYsfjg9MBXF8X4jAOuWbpNv8
7eXbcK5aBZLqkFGArSBNHI3Nu9T0xv3FkR9zFbsJdRmUn+VYCM8szg5VeHYbo+Ax
eUXgpaZJ8zCpSDpCbdLjYjHjwdDthWqBuY6LSrYq0i+4PSdrK3j9aetWObYTA0Wd
p42OQ9+KI5RyC3VjudonBygpCyMs1VumAjGYx5E3U8djUWa2E5/BKaq5eXVPGrq/
EVLAkQ4juhY0lR+q2od3gaff+rfjcUJTeLB/NCuAvS/yFS2CBd+nFrIKdi/c8SsG
RBqiESutrEn1kJIpb55MZ5uzLbv4NP4y7VLO6XIPp00Ko1MJ5P9Hj7rw/1OWvIMZ
KzRYUo0b8ojWSkx9de4XNB4KIucXEg1r9ug/liWGLEKvcmF5CCmZ4KQ3S0g7fG+4
FO71AZlyj0lbwgU1fpG2T4czqqneffQrSQe9p7S5m5vUqX3TpWwrlYLrc68Mi5b6
SvL1pWUY+dmemwgT2RJi2OEjpBlVvKNTD9jqGyqN8kOqcJhn5ffsYF6uZGZf68UN
py41rM45w51DThjTRlqdr6m8GhVf4/wMmBDxYZFoZzh64NdDbsA57phtOmtRDsP6
owK2bmUHxM8tmAXsanIj99JY82b7gjjlNvJscmreXwdkgsTT0m7jnrfutNsN8lSy
WVvRxrr3NaFG6Loh6INhP0RISfwO/gDs6u7ydrBOnCLfQM9th+eDbkDa68hrpTqF
QEZYY4akOqqLy/rKUa+a2n52yw3EUCmgWqiQ/fHTneamNokEjtrleuCNFG1hDomX
siFbSdx/vCkAJ5oGlPsM9MbUA7jONGXSgWf7cOHg3LwK/98m9+NGhGfY8tLr5BKc
6Qbr9diI/M00CsWBqV359XLZEFJBxRUm4xQoKNRiwv/gB7NoKqufAt65skJLhj27
9pnQUcdHHLLreTSH+xwCWmcw8ox+5juKNt3kL2FyzIAeBZbqu2s1IU/xMI1yL7b8
BABumseJm/pcuu8OXYaGUq6ctjBlH3wB559xVDRI7HHJHDdJQHSwfBlqlCv573kF
+v2TOUJWYS2ebuIqdklEZ9gfudyMAMHgns6NPwTiSCZvDJw7fhpqk5BLh+tagyxE
3DNcmGIo8oESFhGqamC1uXMPZYu3nuSs9HtuHSxAFqAds3Ara5vj487oFT3ssf/x
93a+MmFI9yXw7BZtJM3w74xZGF2XNRQTgb3bc6qpqgWAr3h2Uuu1Vu6gb+Nwq7rH
PxgDX2MG7eijCoD3Xv37VkdRiZu/I3xCcHyST3RGlP5Dl1iAgZUnJToRqwFIZqJL
ZK9Y/UJmkH5eAPJztnlKN/D8kTLl1crvvK6OvW1HVfI=
`protect end_protected