`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 99312 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
UPwNTJpYF6a2TR8YjJWNOg7oIGQg7l+s2vQ0mzOxodwdVvmUaG+eQ4YWXHBM8HWH
xJKBE3HUJMMSexUSvM9CZ6msog1Ml+yn9Fh++TuBhNhjMq2GtQ4crGWI4sz79TNS
A8PQhhwdOE8yR4f7uqH8pI8+w8s3hEGjmrfTLhvCW7UPVKJfjbOTKGv3p3/FpKes
ZJ6inyumud7CxohysRSQuqsAKb+DduF8ZZw/zfaSJ09aTofmPfE1AuFVyUIbPqQS
Kke6epkJkCiI0IfajfupHwNkwhZRA8Df5nhxuti0lbxeYLcGBtp6tSbATzPpBk9M
yts/OPIYCPVxK5aXM/XkQVFi25lZLsok1YsfGAe5l2ll2fX4TSiW3GT0vqj37nB1
iOPnjgiHRSLQG1j4Gx8tmgfrgGgeOldxsUJrN+Pue7XpuIVA9QlGr7FiTDwAQZfz
pOkuA77vQRR6+C8JYpMQcb6GQkrdQKrJZj72Uv6/TesMq2tF2vFWAVa61A15i6d3
FDU51Q84vehqTgcP7LQGXUMq9HKAUeaYAUtip+HgD9YBDfSrJyWb/eYDTBEr9E6P
fhCDBxd48Vxcpeg7GfHEsL3/338lykWUz4YNLkKu84qYgMy9vcdJ2m1HqCpZzb+O
4tPyKZ4v+CgG/ZdZGw2S+p6DB5uNmhZIPaEzD6yT1r74z3Og0/Pux5o4+4CxymtK
fyrgIZXGyrk4Qq3r+GHDBdaJHHS+aLErffhmi5636qGOa2d2kNZStP32JtpFxRex
xCTZujnhqMjUxgYfna+nX7krknrF0kbC4Q3jy9qil252Kq+mnL2gXqhQ/HvGkLus
JLp7mIITyz//yJqr6qJZ7Vaq4QFuWoYZ6mZHfIPIV0ORxLPVN6PxleiJBp/2LXX2
lKFvbzr8oiWffufaLnnPrvUeVyb7AhKXYFhHCSDDLKdX9cRRktLdNMn+VSFHYpUD
n8iTfao8IJFz+pkGeia8ASGGNUjLo4OiEQMWJ9P0k1SSlzBDt2JtwSn24fandkm2
c+f8x9K4qdNBqKzj/EvMmZwe6TZbGhw92xtrqvzafyF1G63J72YECFxLv3zmQklV
S3j6jz6HOa0oYPdehJIqcKuyn3/6ChLsIKc43xzP1XSUY90TQWnnJVMClwR+GHss
TTxjE7Tr4Nr/NxfMaXiuTMYNpMJA/HQV8z6tyFx39y939Si/idsKBn8JdhNDC0Qu
cKPY/jonc5vVcT3tg/F+iLVHpdmumX06mhKyBEfYI54rMxBxo655OeD09BWsUHes
k/PgUOoY0CAOMcWsqYmLNx7qLsWgvfJ4lVM2EwBC5lYZfmsEGYw3+a0ppKnDi6Ge
JfrNWWwSfhdDX25KaxrKCnRzwEoqgr85eEG5Qn9Tte7NuVSoZn82IjeiWp6B6X4R
iLgmp9E0dyCbGIc1QsWq+dmz0ltzI+k8ggBhfrfQ6wyeKHGBFfpjYbdY+P8svDpA
ldSUUqiL2jLy/BRRqv8QRhFWCt3MMph0jK70yoJ7br0FTh0CLMhKuwW5JuDEgwSx
Z9/EyueTrgS9QYX9ST8UMmUKSlLn6xHu9j+nQXkZUJJ/kaHcS2tbvtwEdPLPto6f
VwF4j5hsl0CK2YC605PddLX5/FKzIxLX9qF8grYSMm2Vws1LOWxvvfZV/eFpY0cA
2JzgTwyJq/y5sxyFb7vKiSGKuWsCo7oXpin+DhfzssjUjfwWSsuW18j53UAXDWM2
jJi2N3LwWbr0xUvp46z639AyxItLtSfUqy5/4omGi54EJBHQSWkye5bh0ziwhpmG
cjvSnbuQBmhmZTPGBh6lP3QaSF6h2gJ8PZNaW6T1IG1GHZK4Mp5RikHnDc+v1XCJ
pc6ysFxXvoqPVKZkOcU86Om8lw2FaMvnYnl2rr7XkEMWvsSRRGgoZZ1KC++iKU9/
d9fRiEMkDT9Fat0OzdU1uHlxpF0fUUCYuJD8QsJ0r12RnJSoSJ7AnNA+R1dRpCc/
JV2b7sQMBz11T+QUhdVWimsCiHMLDdpmeRs3HIpF3Z3T/pusM+XX+sxmLep+PyYn
WTeTodrRzaQpwCtHAxWnSwNqurJKMCCXZXUawlSET9tkxs/ApKtQ3IeKhpvlMveu
WRo/PJbz37yscGBIt/M0MWGuLIF7F/2+4L+bA9aV39AZ6xZCmAy2mmxCTTvEx4kF
5Jvzm/QIu1ZNXa1IH3JLco2amE9GaEr6WnSFUo3eaC7XqOI/9eBkVV/YLgyCCF5j
VFJuuqEYt4yHPxuqPUDhPM9UPwuWiyPiRkXOalUz3pRJOCDo0bduLG8usmMmXb+e
5hATzHXwtfcZdalka/J7CVVFHKw+PUwtG6PVaeflgi72qHIKuXWRtxet4KSO6xz8
l2eLhPUQP/oXlLqHiDo92X0fBxTfEgpKT2ecPndaYWJQ7S88Z5mk9lWKoYqNrbTS
/owD5ialzaJD53QO9SKo8J3n6S7pYQ4BTJDwTannfV1u6jGZqVlLW08mheNneUWp
SjWrs8mfyd9GQj6w8MVe/jZVfRFOcl/RaoRK1P2zLO0Wu6RIjTN2+I2KbPufSyRN
LMO1RRiUDSmGeKEGgzrO+O2IpVIwz3UbgQl3VGkkEwOrRDv9osjUg7LmAk59KqkI
TaYnXVxobYXdTNFjQADJHj16zwwrZuPm/Lphr9z8C8WXT3Z1cbHQXEuYuSUo5FqQ
hOFdpqS4um5oW0GHG+0NEl3a0DUwBVYmR/hBvP7O6rEq178KtRQ1xGqz4RadPAdT
cy5d6TN5ElNFXDWvFxuzpkojePX97UlUzUx9Xmk6U6zjkgqmys30mtehRIjXuhqy
WfXipPWQSYaFY43nWpH3V3iiWusbXNbL6eYbQDpI6PqVxsykTTsoYmHpW3ooNrOc
gC13Uj9b1kyJb4NpV+0hLp0OZNeGZabduzHcaDqQQMpTooWMBzsRhff0cvEG/LMx
CXfZwRZ+t6u3P3glYmtNUInKngVb90OmhpA0EHvAy8DSPD4nGl/5mJDZKrGLOYoR
loy3CxphWrTUDl2HXabXeRgGu1Nh4u7wTu0Zmh2TVrd0Hbbrk/VLlNbtgXIcOSGL
wRJ3iKk8dBAcxia+7rSH1W91oTUtDGqv54gahuq92xuUwFUMJbyNqvKw9SG55oRr
ue6HSZzXtoZqJ29cfDfbOI5OlY3shFtG1RtCnYqLuc/Pp79OH21amNwdZx+AWjU/
/OpjmFQU1gPeo35cR42mGm/trpXWBrbe8c5YHrdHxg1fuyqah8n1dOsg9+GAo13I
DcdanQ+BqcgpZzBhZPKTjdn2lVKIn6uxz8q6oJHIQpsLShsoB4YxRPGX2UBEXAxP
3gkmVcpuaJAIpDHvPFyGsDLUd/vZJVEIrqxQyFV15QNF5pTm5ZUNItOg8J1CNvwN
v2gQ3SpWHJkdBJoZzd2EBASOwHGuZM7c45JKyLjlnrIqqP+OjISYIV2U5B5fRjpx
IgE772HqdiQRsOsfEpn7yURLg2mna3QCWDiwu+3JnLHQy7ISS+DpghLZ/7lb8AGj
hZCrwRZwESXWA+S+BVBzhxNR21EtaHklMym5MSGVk11lQmtT5HwlK/O2RJQ+k5T1
rRULunPfIPz4pIuiRSOwN33Mj6dbtO3Xpqmbz021MUgMX6PIRGVSE6Y7+Nd88a/2
bSxNG5wxhy6UbuT02E5DB/VSJ2oHaFOyaj0Ugnu/YAgR76rBxQRqOp3cPgM44f/y
tA5vQO3LMzamq20bwd+Yf/KugbcMrUwFXS2WC001ac+RtetEC3QHCz5TsZQEg3vp
fZjfaDCV2qYuqxvk09ttmVoqOaIB6UwKLwrMvU0ppmlK3pD5HzUUQ+IJ8R+V+4yp
iz0JqTsoQcrRkK4kZyM5mS4c0GiEQGt0FtrfHtqvslh47MmO+T8/0fYDrAP2ayb9
tC27U9vxhR8McPNNqQ91Fp8Zr+f7rZodQIvvINyvf7YpD5S/HKjWOVkCYaJhloOs
zZcOPWUhmnI4Z49bibdFgm9BxaJolFwqm7MsFAnOry/c0I0klfvX2SVI87xvMlGw
blBc90JUZEJPMmcmh0n09NFMZSUgY8yYf4+czFiepubR4NPcOJhd9CmgvZPUd+xi
nHlbVcwcsxB92z81DATqR/o7A3l5z1GcON3kQnYa4TcqPyAiw7HbsGDILo7GBHkr
VnpSy8BsrJQAePwr+Cqr1DovTuqqZVoeTJCPd0LWgqLfSMPLzT/7Xt7OVO+TUvhT
5SJ5e01c6zFIQvoRpKTQUZNptEVUlQjMG5OtLjbNfDET1hb87JrpFamNqUQUmwUH
xrroF1gu9x42eMZDDwsfzMipjQUqKmhVAoj2Mp3rMCPEd96bijCpfueq8cFYUKa1
VmAOVBNO4NXp6ShhI/CrIOKmlASMhIXqOKBTdML0b3HMFICGJ5bJk93FqYLiAKep
lnK9BLXm319bMCyvIZgUO9b+ZJRcra+eam3JzQgF37bTuKL7rkQ4JnqC2rOupQ8+
TYGLBAPigGlRxuGeTYM6e5RKEQzLT5htBs9qV1FumsIfTVt0EFPmXjxaNERGRwp+
Af832iTQWT30s8Pl0oHYN9V44aYmyE02yGVzeadAgmhDEyy5kxJPH2ukKzD7CaR8
fXsQ7pNpYmlSb6anfc3LpJwBAAifMUL6LGvGpftPxlj7UXAMqe9S1n28wC0C8uM2
wdPb5hqtr6AJzppWSfjJWAHitZwrTc2c0ck1rKaXTau2CmKVB+mjYWyFLLpB7Xqd
6FNMfmTybBJ4nl8rIBBiAwvmzK7zUtdM3saD6eoNxTNbUvwc/tb4UPJKwowPRooW
5zeOyZsGodCJwPr0do1gdfpCPIps2ud0y8XSCV5IMghQfyTA3wkSIRym/3lvCqE/
3XnWH7iukr3PN0uyqxGTYbSBfyBGk9/JXIpK8+fXoJZztplUugTrtsVXyT5jbuXK
3cH7wfJJCI+ki4Zxs++wxS1k8apJcyStOovGfem72YDi5+xd9y6p9Q8OEjs6LJ68
roFJyUaK76hvaI9nh2zI9HL/uoO0cuUFeflBJkFLEIyPe7B0yDy/0RBR/KK3Y8OM
6o2v/SZhJqfiBodtZ/rV0hO+gFGFVBBXix1+p9+gX9UoIRquVGDVbq+MBPVDI7Vi
TCqCVA/FAksxYOf5+9ofzZk0esQGhowb7FJyX6AcanaMlZNVTjWnBFK2GEfht6Tk
+AypyZEVU1krtyZRJJK/8ioRtuFel2Xta9Hb+OyRSO0F6EW7lzwZPlH/Hpjo1keI
32ddItLVIOqT9mz0/Rv3Ez2Wl+GntLkYW0uSOTKDB25ox/1msDgZfZFLqtEV9eDi
AuG5dZIGmRoCkXi3vw0zzdP6hZNpUJbXNJyS3ZdWF7gCHRofPPU0REI1VHjS11vi
rCJ/C69FtHf/MPB3dvSwggg0wyEYB8XW4dA9FrIWmJZU0F92odO8Nw+oyJv6r8dM
rEGCILHxhw+k82sWqo8LpWsRcPVHxcIJr1Hmf/irounYsT0tKBaO9l44GeKw2mml
DpIkfODvm+PaUHrhfbLLDEUMSU4wN6WQzq3k1EkbBHBN9KH8TIkY78HXeuaSLjIM
+Uye0ay7rsJIAYEdLTHnqql3vLCit/Zn4wKizTq5eXuPsshHmQZxLu0K9/OgC1Yd
bf52VXW7qTofmJWnu5uM6eveI+EdHwH5i7195Bojk/FzHzJSlwYGd6gPISXHJ2U0
1zJ5GMin8OMa44zyw2GK+L3QrEef4qSWWmURZG3ldt2iRfrDQs0oE/5hzS+d/WYo
sM0CaarvvS31s6ScLGW32L0plBLw3T/v7EGqtjcVru4cupY1KE38sRydLcxByFCo
cjQsoLh13y3KgyXjWHHG/1mLHY/psqmhq/HQW0NK6WIOWAbO28UD7GrkfaQpws0b
Gsyjbqcdyj2EYop6HdAe5zoVCYItdaxJGZZmvAo2uwFyo7JI17gAT/6BU7KDxqS/
f5O6kM7Wkn7HAH2sPL6pdTCCqoR1bTuL3SmPQqI51UvhUOjTK1rQ9JybhlJ4h2Iq
Yk2lDElEDBZm9ycQ1tkL0y2EwgzVpXsC+U0NLw60oIDh0GZRU0EJuTYbiRD9kpTH
w5mSGB4vHN269o2WJ3811U6aYS3mPXy7Robu/0mOUCYPzLXqRKjpsBEF2hBrb1Ki
xpGUP86KuKj8OGuM/feFoX98s8OLGojT+ObQPEPkvh6wfxtvf4BzuNnOcE8gY+km
7HrbSoZcfPmEhp7qIFKM7MJGCFnSZ7WJQpfxkQ3JHC4Mts0asOlX7e8n9pqhGmg/
hpO53NzeFdkwLuOTUs+tQQE4Qv+MK7+OX5zl3LeE2IEBD4Je5cqEQkyN3GLhToJj
3o/hBdjICQG+9X65YwMrFNrpxFXrOG2ZyCtWcJVcAwjgPyqBIziCiVe2cXXl7zEW
pNHGF4zDI9jlr6wlHxVSWd8wY4ym6bxjnr9+UMTSOg7ntcjDUuEvf1638LiidaT1
oNfUTcPV6+hdhZzArDqTAbQVzy0m5IP2TvAl6F8h9BJWqT0ZTQG9XkF6ZxHglQUx
dAhr4o7G76RR9TUsq23jQvIt0JQ3IAPhQWs6+wNTD2onjT0ooTcuVgMX+v0X7qhW
yWBIojT1suXpx1JV1IHEQiQxZHoHMBl10ZlbfoYBiA6XFbGCagCIXibDfpcSfvP1
WTwEvtgmHLFql18S+n4KXHBuWVAborisAF9P6R6tYJ7sRHufPYfW8/74LjUpJrwX
ye1mTzRrg82NALmVkb0jOii521BW8y5TsWQIg2I0umRnjgw06uH1+sMUDuNEirNE
2IMkyqP0bUj09EoX6mZa+qrN43ak9sXaKakNlgVZa6xIuAulScAXMXyxEPMAbLgv
jKPQFdGRQnCMfRbTwcq5Z0AIWMg6febNDRs5j0Oxl7hFDs6D7Q1Y2cRqwVLwZzV3
mlrpIFqB9AVTlw7BmH0llxyDE+bg/brusRKgCUgcBhLxiYe6M4d1WWhZkKZrvgeb
Yh1uA0i4vLgoKqRawgy5trcQ0t5SzO15x09z7V189uMZb2JcTIXL5yRJy7jdBbba
/9wCb4A0sOWhN09ebFv3nXv9AeW1L/qs1RN+iGhHAfj38elHAk5xjgA03QoNk8Au
8rMzp3deKBj24WmVUwDKuTqhSBqGNNMK04nryW56IOQ5NIMD/hDoG0iuT+YmRLjx
TMmUG9MxgSJWtmcLCWbPmYywEMbDAXR+N7EOWkGVDa1lqr0VB0V+Xz5e0IIn3Fsc
O7iUbrFJO861cW/4DGgluQ7fq00ooqC8DbJ/w/VFijER3Zq/x6UoL7z/rtLtXr8l
TqpljPtKLxcezHwgiPFeQFQO3Dyx4lOZnP3bgtQW2VaMsP5sP3YxbugY98BtJZoI
XGe8y3N3cvtgdkur0myhaOuUHcXGW89cNNahGF5GuAuQmaSdLoiEhg5a0BJuX4FL
lcsxCsHJElEMtTmh3VHPTjhslqim0UK9BVdPPdTdGhLiRPUM1ejxIEaem0bGf+6y
DmcGzRF6k4hckvD605eWF0HA3782b7zx97mtk4HeBAlGSE5hEB/gv2zkYyqD/G9K
XbTfWyQ/arvRtyHly8fisxDIDADTJyhRXvtdkxAwH/WXSc5wtiTJ7eS/BNykLsFj
o5O8KZCTh8cQcwlJDOpDzHzxIi7BZV2D8EM3Wkc2YTUDdttRWrXDqubW/KwxV2E5
/ILmLohXSlBFV9LVtEwA82WcT6n9WdLZrzmThIc0Od/SQold8kM7fzyyQ81ByGuW
9+JGPcv+NI1EzUP/T9cFnDrg4FOn8beDw0/CvwOw6ZCGjowMFgs2gE0yyD6hMvuS
XBIynHg9S0+jYhol+XgwoY0M8V/pHkXx8CKcwlFOm7HtKjVst2J1zCRnKV25WoRx
Bv92/jr/2j7bDD0N3M8KNGU1VM9A+QazPzaGWlrRcrbly529PF9SexY1FTSpz2kb
awMcQ7sBGzdhidJoiuWq/Md39eXeNCW1eG92wUPKsrkG3Jl9J2MxT4wt54d+boYv
W11bUAHV9j/QIHOEm1wHaRcriIcrKiOUpz0lteGnl1SKkvW2D3FG8l7r4UjTjV82
XuxrfQylrc4SADQzwMY3oC0Ee12D7M40hpWLZ1I9ZKNuVk0BossEeHEIGx4maeO8
vzTdMSXmHLKVfMjqFEl4jeUNOUiHS3R6TngRfKUk5UiVKayKVr1CJT2//KLzRGDr
riYoRktfeopjOq58HeMvGa0JpqMUb/+/JK8Jrx9qJD3z13LJuBWXWNAlvfhxwzwK
DsALsXE/8c4s1Ddk+tY9kIUn/dMP1lBOpXhABFctJBkLLnCqE9I66O+RXtiGXp5F
RMjkHX5sSMFloEnGhMhyAoOg9hwBpzzXHlUwg12czgvm+RVOxoj9xpnviUbzxZZ3
/wh2NUs6s0jIX6X2syPJVETJGQuZTXN/awCa6jDhq7a6y1NgN+KNq6EUvRNzLU8S
AWBw9T7Jg7SVE3K+IsTy2WD9o3Iss392hbS0fiWJK3adWIbBIAq64ovNImb/byj4
JaRa4ySnS5cV+bSr96nHPfiRqf5rpi9bKSU4WqsWSaOtE6ikWkM2ebr1Vs3COMv7
kxBNdjqVhECJMVL0KC1GMdB4YItWKYRpcLy3Q6KBElVGJg5tU7CBc3f1p5lbVFCo
+t909VHHRMueKJV9FkYdXHM7e5xQrbRzQ4AgMe1UkpmQVVOQS1nXSVVpYhE/BUJ2
JH2FlEbSQ99BEAWEEE+kQCKEKzy+/t8Zhhdx9KEyeBnIVlU3sNGGeJaX6+wOar9a
VidEb2v57orjrshrWMHaLgG+8LHU4gzAWcUUpaIEyc4gNad8Xjs8C/fmeKGIKhCv
n9MGPq8Vqij8zmvPlJ24LQvEQNoqEXnIi0c6mhPM8+LIUNWORtpnqluYcE+nWtJ6
jflAtGEjop/KLSW5aG0RcGSBDZEAy/gYYJSQE2AMNcNVlwsf+mLlLc/PJ3rwmzXd
19cYHfbMrYFh9tiEk2ChfXtrVM3iYwZl0UJASPNXyBEWb/0Lx9tMRGBqFe/lvoUR
ff+FtuR3oY4ALenUGAi4FgdQDMlA1mSTh0yMpigIFM/OIedboELjExJj6cchXK5d
xlrQ/4BlIINNjEMDBa4gdWjPXM9T6GCeT0U0upvwIihZ0tF4sZsR3fRXg2q07fLe
YHI9y4otJfTehxRG8T+oDViDuU0IYNCY1TkPkoj9CXnam7mq5q9xkRVDjz50g3Bs
LqXQ8mSFJQlnNRtyEZrTvMqFNbA0R5PbJNGAoybCBfLMbYRXeDznsHmMr5E5eVKA
INjcqNNvBJl2RdRCsR4hijBPwCLzKligAoD7Mzd4HotlsgWHSDXz//MkyQsvzzDf
OU1/LBeJtd7TKOs/w87NZV7Fv+D+DEgvJKYVekXst2Go/LPY4yR4AiudxWLs9nxo
r2oRXzuTzRqQFIGyDTtbOKJZ4AZsAZM4T44RLb5qoSnX3/YubgusN2tSSFobA7ZQ
9GK2EhRLcY72aOGpZ2oUKA6+V+09CNWFKzFwRgPQDgz4cv9Lj6JdqWNp3Ly00KfG
kUGOHMBchZJgNK7WFZTvNIS5Njr6pT5ZfOsgk6U9LmVOLEQmA0XNBXNK8wBJzOks
2qj3iIsmKd33ZJoRwtbc+xfblObWZdfbamk97KpM7Jl4SMhLFksan92LQ7PJUIuX
Str4hlfq9i0H26W2bLts7xT7n+jqIinHJDVeJRlNbgDQDIE70TNQgUgdFrLPsr3s
8jIIzEjap7VR3qBh2azGWfNh2c2UiLWGjQDBQuDUpMFbHSbEPNq6ACCaFvzVmV6Y
s688VnK+Y/ANeR3577k5GhbvefqorwRkwbpOCfPA6bMKidjGw+RqmjRt4r7jnpMy
fNXAFvkaLEWMIpJy6hLq3OgCjUjRNhq0HWmVM9pe64wm+s/XaGvFWs0Uc21TLgmG
34L0Oj13UeSWqiwl/sspkcXWEHw81ivoGW7gdIb3HJS9AvonaUn6eeS9C6WAhzFU
gAoHSy42FARlkd83HEjgDwk+tD38/4tdDOp1jMzgjAHDFo3/I/p2gAs5kZQFv/7K
R845sIW5TjIn/9anhgVpzioFzUmyb4c5PQJ8vmwsxYKWwrehISkyH5307JY2VPTp
hJv4uVieIA6qdTUerRoRkF5EcL+3pIqU7eGPpIGSUIfW3ooPZPJdojXQdTmntTQa
fZp9r4iGUvV8YW3gx31s8Oxk76g74+y+Sd3ilTljhriVekNR3efCASfTiFoUUuyw
NKtHRVk0eoNpsbC1RD/eOGOVCdl9QQWvxcl9+kzkDVnDq04Cy0gWie+4Gyy7z/gm
SsEnG7W1yG4UvaDuAZ9a8kgO9Tj5F1/dY1zU9imlGleWdhbboBhT5USEHLIemz8K
WrpI/Kzki6+dvLGqLyt5R9S9g9Jb3zUHWX4YLHciTgkYW8TUlPXbWCNFFPYRnipq
8wd//tGos66HNyfcGy0Tba1/YVoIRAbU6xPuMOsHG0WEnk7DrCS4eKqk9TFW26mZ
vKwQ7WaTM0wxuIN+4hjo9ZdxOeHe3pcBe/IF3LGd0f98isFHz3FTldx65KrPNSAt
jKle4NJw7h+pFORZQGeZ3Xj/T1qpd4B61o/nzfn3nFCiyAUcfGQRTxm6Qwi1HDtc
AJEI/UBH0037pZQgvE3xHAgmslM75jgq0wMpN5jdEIoll41ubonuMyTTTN6XRERQ
2pDYrkB0TJQi0ukuAX0UkaTeCvZYiEydwnG4OH82rUZQX7jDbonCyBNw0eNxb9L9
p6FybjrrNWd+mRZdIBqrb6nMNivYqPdxXCI1u3+6XMA4BiFP/gdOLOcvJQXeTLnL
k/BqnsiWy9zz8qppnbMmlyUP7CFNVxhnp9DLgyBfc1Lnc+TFCPVFd97lyPe+97xa
cW7ZIbBncD+jQmOWbaFetB3YRdD6HZtRnD45Il9WZ8V0G+k17N9PgfYm6+u85uV+
qFYwRd8FdvNipPeMTnzYZ1WV3JiUH1eZLR2NPNFGbUK/WWdraoiLPtElCcXBjJnu
umjvMHY3OsQVALzZJim5LEfUj9/iXm2frwJbKQv0wSE6N2J/NTbQSLjAJcoL2Q7P
r5P6PFQKgnREAy11PTbTRH/KLfw/nVl+itOMS5Du4TDz+N/hDoHuxuJmVwUf/q1K
MpURHDWoKO9xQsS75CBuDvM4RqEpdMFITrbX8qTG8sWyYjUgrWPpjBn7AIoQPuzJ
k9U5CuOuEvKeq7xEm5ohEjkp2Maa983ccIsKgtn1Qj2nqBlw7vGmx8Fy8kuJIOCH
pHTYvFn+VFuTY/zFQVe+bx4i56UmpTTF0dJUJ5D+/7bwRv+eBJcX6a7zC4PkYPau
5O1+piM1A8rc25eKAOsopNDqPJBVCy8Fq825UKgvgLGFOsMAx8YYCfwNf0oDomEH
YoAnt+b+xWZAFC5nx3xEf65QvziqjhyHmOIIqTXoeWY+yw4gp23kUqt2cP2d16zJ
nFxbEyd+cJf/JMi3XfSMmhb8CSf6tW/6uJ6XEfT2eBIy9T9nkBfNNzdwOjLbgtU1
JBHEWYnAhKrEviFKxuQmoWoFuV17/fBOGayUxR0/V8U+flLIZFjbHxvUSaVexBWZ
TGD0Db293G9PfAUDDA8be2NN+mMIwqAg/7EoSDSoaHKKfGR5kCa7m7SE+nsbrlYF
c9khvKJ2EJFbbwpFqstTbGJq1iDfqHpV/3lB+f0Ezxc8DhTgry2vlMLYaUyjKMqP
lXDgNKPl/5E38cI2/RdT/fk/gym3wpVe2HhJ23FoBeeeKzsAwowJEX6gm0duCPni
jT/UzXjS45CyLDRSaDo2gbRhyzRMWVEz8cnZyAvG3WuUuMvdGkWSwnfJ21g1qmUs
7kfSWK8NciA4yigioYLkW3Gx12oZRR8RmiHlm8JHASZ088iKCt6le+GmPDXZ2bM/
U0evxX5D7Cl+a463I0APC715Pb8pxEJXhwLWtq1Ie9cL3Fy0g4JWeZu0pFSoc8kR
AzecleMXhcvyHFPdOVrYNdufmwfSdp3xwBmYCcgQ/CaPCVX5/Y+mlTXQhWbxr2mj
DOeMXEAepD4F80nsyeEL6IW5xmG3Szbof/5vE4Zq9iTHM9tVOWU0yntDp2JTg0W8
K4ULkyWDeSmQ4gKiPJUQaP12R84F701BG1OhAmBaATNYcW+rsXdY7CmlAY/Xdz1B
9YQDiRpaUmog4UY1ywn6vePVX7ZhZhLOwlgcOCimDsPaYG4Lwv5e0CGDXyffDdVc
BfsvUSLyt5t/gDHxWS1R9Xmvt2D0rErGWyJla1SOqyCMXsf+uCFZ4JSRtPwbEG56
tfIMhrsyefZYw9doVn5mMWku9uDkpW377xL+MFwVuc3LjZS4PlFa/odgz3Hnl0ej
N1jcWq8Bw2W78ajXaLkh8oQPYoQW5cvlauKpopgzjjEPHvas04hRiO8fSpWnoLz7
zLVl2q5/VMVkvShmD0iDAsetnWLuYdAWzNrVvpVGCRyKSH1LPHhxzdA/+tKT31l6
RL8BKPQ+dGh30wG6w8xAo6IKg4W08xhhlaLm7lnU6imCSNMqUssqEPA5vFtFOx87
qs5Fly7y1piN1JeoS331hByHoBMmH8uNY56DDpIv6xFC36K4+05qGRPaF/zZAJfk
EhFEgvUiUQR8B5qDpwWvZC7Q+brls8VBsoQgPFWTTF7INHvck+S6UQTZYf4FhqUQ
0rmJiT8TB/qJl8FMZ8CzJQ2CFOu/0cSNDF6cEZ9s6dLjjSavrpHXyIelh6/C7Lmr
mwC6Tm53G+IWc4adeY5/mRQba5HuJ8yoD1Rf/xIhx3/OumcCBzynd0HO2xGHCbm+
KfBPDC/SoipMk/YEsps03Uv9NxERAMtelpPdKhotxXLX0McyGqlDv5on2QhCNryV
JFmm/aDbbd8oByFWmJ9VC7SRosm5XN1vCjCsAASX+6TY68VcHLSzLE91PFjlS1u8
5whMQEJ7Bx/I2w4mrWwl8Yf0Qn2yVWrhj+fBTDhNI+0rOF0lSJ0L9jkkJhc5JMer
00XuRXdaZm8DBVwH7nvvOOgo2Y6HPtDXxHRsI7cr05CUgVRbyMbWiXV69eu2vozd
UPfnyvGA2Ap/+PmidvFdu4TZCGNqkcwl/3a2RIDV4GAilBSjj1VbfhQwRZYqH0az
ZLBAQc0hJjyJazR8oHWKizQhb7GlKHRnk2mdJyAWUmV6jyF3VNV9bQsRiCItlmz8
rA6tR6q3pA54uGG/GgHGNhuIdFGPT8ppXuMXg8R6sBEXLXON52vPrmknXMMSU8pQ
9Ut3nZ+AwCpiMP4jXoj+5IzvzWjfh4C1XqcgdXyzGjtqm45psdALwXIYwhX9VubZ
9Aqk5ota8m4/HNkM1NrbbY+XR7W/3cunkIGv5J5UCquf30D3YET7pvuymJrl805Y
pYY8w3DkcFDKHoGY/cAGUOywiMlBgrLPLJ/km/iYkqZn3qC4Y+zb9OGWOd9rF1NM
9HXvvwU0ydlMitt6u175mlqekXi6pchXKl4V+4admA2xTHA2XKRSJy+9cFOcuIRX
1q8N5VJmPXU/7UhE5R+vZKetrCpU95PtMJLN7MK5d/N0aJ5UVMtpuT6WlXntvFis
0y5YrZ0r9o1c3JyLD74483Nj3L3C3ILtJ03XF6ZaSX2ABo1UiaAZ5QhBN/HEvdPa
1OI5+5hRTzB7LRZO0ga2nJVw35XOk5S1zDYyglwyyVXMQQ7CoIuGjRPby7n8KGOQ
FLilHN3FqI+EvcHFnoKYtHeWNuEaupoztRsASjgrObHPOIwD6/il5I8o/MH57poL
YrlaVmbeFVw4AdX4n2XZlwo96LPlS2ST9TZbyfnNLuteOlhqXEtuiXsUbnUFAf9R
QFTBLaXdbT77Ur8shgCFTEwJcSnZGkTLXUkHMO8PyXtPs7vTQ6AmEL361MTF8Mnk
2ZMXZwkBPdYNIMLIKEA+/Q6A0plmk2LFJps0mAIBd3NcSuGcXTLigHdxkf403G2b
GSr16ESAC0DkNMBffIefJKFvGXzfwNMJB8y0aiB4rs6F9meOkby+M37Pj4ZAS3Tq
tY+G1OvRDEJaT7zfwdlYyZ8cAXtazh0vNaFGHpxUoxCFuLXCz8pdSX6ENJAsuHTW
gKkfOC48HcGeee4fzg3g5bioo3UlC6YaysWxntfQ/sKkSMiUDacHarixGJaZCWDE
mSE2RwUmYbjjC2HBPORxd7zFar8VWlVs/2PoDZ4nmvGXICai8/Ig8jPZ1Uf6jNOl
lNdtifd/GlWBL8FnB6eccrrt8EEdWeTUEzAA/vgVhQ3NPcIauXsQctvJQc2jaQX1
BGANPtoxm8bH1EsPfeX+p7+EW4fNwc6J9LTBbWn/n0ABH4dRgMEiwo1tPgZRFTHs
BgbD3q1xhi+LTQmizpuPoUIG38LeX6mQYti+MQUkiNUkTi8D+BTpLSE91He/SIvC
EBi1V3ayZC+x/4ZHJ4PxeyAPw/8lwnOqtQJaG1kMDgO8KD0LJGtBYsM+TF/wNNDN
w/vebGzOE7OSTKAGyQc6njFJk/x5zWwgQVn3ZydwNW+eWGjKENDihLZirT3lVabw
yqSXmAaeUzAr0sTn363q+Cf5oSxG9TmoYoXwnXBtgJCQTfTF+XUq4z3Qo3E4LMce
UaMPGL4GourlX1pdwKg6xFg0734c9P5nqewUGD6CV8JNbjoJoGffLbmyPP8O3lXu
Lhk93x+DmCeDn54ChUIEwSW918WHnjlwOsIVHPDyOkWVi77en8+mfPxjgxoxMgBF
QvvQHIAm20g7Ux5WUyICR2Y5UBQGBod4lyYrUdZOL3QYMLr81bQ+0GQ3KbN7uARp
zj2oCpI8+0wOpPKj2LXDFi+Ji+8JAJmeuz83vXtHtSwLZeT7d5SMcMRZItOP0GJ+
ABZy0A6rREE7aWMPt5pu3wEsZzgWaINXDAOy12sunwtNUWEFLkpaZKDTg31FHRxq
B5XQrHqHFRrZpFiAccB0o7O8AknGfVWZNUwxa1J2xgRZpgUA7KP8w+hrYeItBO0O
WV7EKtGLJ1gOB3LkjjyKa12dadK5Jcln3ViyvwFAKEMMUSAw2C+N8VaMPGLFMNIY
cUizQFujfn+pSNVr3T+OCXdno2McmzHUNEYAezT0Gd81jPC1rXzdmR6QYn5Gjjk2
GDk172zpPSuMNF500SiQ89lKEnufYwUBGjHh4jCBLCE45Li5yHDRQAVKMUyjWOPT
n6kzgWP8DiIOBI4bHYhX/FKDKS2HPs23j9PZKdP+oX7LNc95/9uEchPFBSPZdoXz
jhMpwZd/iJggO0gRy/hF0Xba2G9QcW0sNBk5C4c0UoZ7EA8I3oSmpnKh+4kSgNNg
JNozNKuRhseQYboWiVsaJGFJrGwfjGP5NKENXccLFieyBtSoqpNrW3RUx76iaT5F
RTw4Fv1a3Lalyec40MINU8dDmqcJOCGsL2ntcR6DykB5YF7H4Cw+xHbSDJ+CxOW0
GQPtZwDP4/AsPnU0hjtVB0v+d48+ycC/GYBW62EBhgzcQADHrjpBcUuMnN84KNiZ
GS4k+LGPHVpZpCv0ptyhew0uG6IuRUlek1PjLX7HLVrQgNeuFLZxIvr6Irdpnmd3
OPCQ/eR0Gva1K53GFHnxPsU4qqwG8ojvh68tlMzRD7NePmIn16a6YJ9GVb5FIkrQ
q/d8+iBg4z5X1vNY7XcR9AHBvInMAplCzakqJUMWrLcjrJQve8h6DUldD2Nfj8OK
JnRDBHgK1n8PONqKGg4uPtAsy4xU8CT9aFmN1CnCCC1Ocf/JtYDsDr4NsfVm177i
bBMxKp4Bcxi3qNjAelYMOjf0rgvBKU0j0Pkf/iKY0UR5hypnAcYe0IXfqzNkE8GR
qfOq2KlyBCstop5MFaupUi3qQGYJRnNQjv2b4EUfl9N5IKAJvidSo0SWCTswOiXE
VZdxPQDQ2LcO+6+XxhCRnzUEtYSuqXwuyDk8c4E7poECHAh42/SKfpW1P5RDzMlC
syTvsVXalJJlRd2a99lNFu9/r+gDJFYHklJQMdYLAqsv4ekURGvgctH3oX/G0EHF
wdXpD7v1eyuaY3vzCKT531//ZRXKbt+hViUppNVJCrNbwB9QsST0YuY7bQ1a/iKg
ITywnWL+gS7uotL6QnSHR7IyuzwiHPTAegld4rpVtl6uee+/WFYbCPkEdHAQN6Fo
RSIh/Veu1Ee8zVLAWryWQR//2/D7hca9h34Aheg3a7GId6kujx13q6j25guiFsyY
5AwlnK9hG1R0xF7dSC4uWgDitECM6PDcrBccPtU59NJin8XFx/vLEoAia6Jx4U10
ItdbeP/CuEDhzKJfqJysh1lyGvBPKGiPPiLCy5BX5kPmLljUfiJEPAC7jQhfUeop
B4k/eUJ8jE0uB4wNi4oGARP6RDD6wPJEdsCGnB2pZoxrBPbc8oWEjnEadaOjFDoT
8M1c5jkX9xLF9CZ1OZ6d17iP7msPjPtbeHnIopJZC7bEm7NFC9l7V9SpdSoqOTCv
n7j4vZin/EnYCnRLF85pM73O/4n0ZWgCTMLBftMGruVyWpK9++S8PAcZi5R2JYG1
s1ZgSYDk1grTE0S1RlN7p4f6u2mldSH6KXOozp+jVxJBovzHQFDEnw2WcykE8KmA
teSm56ivfoBme/j8r8h+GCRurVVvyvsG2GdnGm/zwZ8N58P5MKb6X0IRSH2FCKeV
2E8prC8mtMsUkfkqCdXlBVLwCJabuxhkXbDRmd0aYeW5MfIYBeX+mpMyLM2isnSk
TL7yeIfMZfLCWqsgND+NZ2TQgShAA9edvET/PRwS86DZXmcMV/j7yHGbxrRwViwD
g+XElXJ/2symsZzpF36Jt91P0vVAZOwftU0kVsvkLgpBflTgUdcTg+4DjL9upoCj
nQdAB5rAQiVLK4vl7wSIj717RoOv1qhF6YzvcV6RpyYY/NEzF8w3ynXhreLemB2M
cQXK2tLUWTp/EjaIa0XPSrnofsJFA/1DXxNmXF7NwV7w/6uGuVZiIH/0V3Ayx7/j
PqX0XL+VrJaduubM4wH4k24Cpek8zONhbozCulRh0nsENqSdSAJe2N8xBh+61N49
GJ/jv9WFTbSvb5m9sdZ2bXA7wU8zbTjmtiRlmg8NG2wVoRrQ5xLKErCBxiHzmqxI
RYy7gidgxq9Olo1v9g6xz/oFK40m68X9ulhCAunQGJM8lwQ8f4w3B3HgzfFcsYjW
h/kSPUjkhmmtQZL0FTfNiMcRtHrZNrtAGLTcd5mEbaGw9rSCA1Clj3JGBT4xrAwY
dK0aCGLwtFc8fLE2/LEV2zN1i+Amf1Wii/dOanoocywy/D1VIZ30a9awkAWucXtp
JbDGwurFwD5GXlhF8uqnumvxuYRtLAoy7Xe2holH5L77RUML1c+ZQvDCLkTw3Iqn
hVSHuHsWalAj7KwQvqHT/Hse8tmnIERw0doXhFJznqjXF+gsO1BGw8D86dvQHyhQ
XfEyOTxrAYxEfc2vgP2RZzxQZMuEsoLs1Wowt2iUaYA4TpLNDrA4Ej2a1mQSk0cE
FNaF/AU+Oc/5ST8eAS0afaszo6l5lwGtc1kCHdKpt9o2btmwV0Dt5t/pmNsEIlMp
Lk4hhHk0jxT/zlg30/yXSoAAwZQNmzYFsqlQoiT4/2Jf+sfGw7KDHZHymHzKAdAS
6uo2XaMOtw2EQKSwCzXZwvOnNhxI1gA3eVrHzfRybinpPgbMCW+DJTGBVpfiA4ym
Ut8NRYNhcgWYNLiv/uwGoqB4pU4BoNTuK3upM1iScHhp7qjGTXEPIOX9DNS7uj53
TY7CNxnypjES+FIsiMcs7VauV2M6fVqBPRvDe5Frn5r1iCMk1XTldetOeXmANNTc
XolbtJlGRe31ZtPVumPbG3LS/G+OCyzBEJ2utfou152sNMivAH6ZvOfmLSXQi81O
KZ3NaX+10SvyqtLw0exOcR2HVUmNAgphYLMy13T+7InVNccQiIipvQlLKz55hXoh
6+hRIlbou4emihaxZV7NhmEbiY+FzLVD+jfsEK1tAek2sfZJwwuGucd9ttJ7qZlU
wFMfx7p/lcY3p6GzqZ6gv/U5me+wJOGOtw6HsSG2tHcWGy8TA48iDDZklSeoJQZi
+w0sXXLiiTTk7sqzVYkaAXHsMp0m/rD46qUBy0ABoyKFolSMm8hA834SuEV0AAHP
LUDs9nQvb8RDM7c3UZRr1oShREu1xPV+rzBorg1zEAzgNMsm3czkN+wW8k55WHo/
zw4dJ2va0Fmjk78BOoUEB5BZAKZ2guvSm2B62OwE2WNOFoiYDOV/ZVRfYz+j0a8F
x1JNYQ/iDvy14Vp/23KAEmKtNOqGlt1b5zWC9a1+3d7urcAHtIEvMzW/aQl+kGyT
JEHiArheH2hacGm9gKSZ68wl5J+iL9FzkTcRaZKzE+jf4DFWu34qsnQEflnclK8S
IXAHIdhkbK9drH9FaRQFz99jPdt08wE78g3bdNA0gwLIfMog7EtTwfGSDIQgWt01
YbKWPWG4JD7LJEyFXAZnKGZgXbmFWGg35Pz6JjRtwBn7QsZ0iOeFYngTcTyYpGAK
L+9hO5UmWELqAyTuUKdf2fTkxcPbCUFqC+bo1+SefC/1ZdNqARdCtcj8qIpPXuDT
tE4JrqrUT+2QaiW9DR3D5FHdEyb56BvAIxbQr1t+A5x9Nl/z29ZnMe1usMjE+Zi8
RVSpTCTOBMtRYY1lCd8pzkohnCO5UEPN4o8Mcrye6rSZ3nBAGiTHseroqMc8d3I+
vMd/uNqMeBsRbOf5MobDXN4bj5dUUaWhIrx2UdBCG8ONPhphEoh/FUOnuIutKYiG
AbrlVuGtUl0QHd1wXl6mjdK3v7ANCNFcwaPD1AkFdSODUuHOBMdUuYkv3fAmmqhr
lla4qYzhM0ia6ntHeeU7natWaatkFuw4Si2vEVdpA9E4iApqszqGoAfE+n40uvOg
4q4ETHHUuPX88CwOTXqL2sYCfzYbEJAA3Fq55Zpwu2FXH0mS/MQyVQWbAKqdIRdq
I8qF0L8J9M1SoN87Bgd0XxnWW8XQ8PpYRr0JaymtNNYxQjPS7q1myCp5JYfOERcd
FipdMno4yj+Sya055i8mTaPEjKZuVpYiZC/iLYzU0DFkyBlOed8T1LbnwAKqQgYA
LyeolU5L/+zZmK0pk+n8OTbyN4uKrq6pw+WdKnB4n1gXENLHWd9p+2IcReqFemdd
QTZ1Esw1qYvPRvNPx1Ex9YmF1Jes5oPaTjkL1lGNdXMygvTkSkAPALr2TwzUEgRm
0/h6LIHwlWQdDEeycbv04cmCpyCXweZACJFMWfy7a6OsTMaAJ10PABhJ6Lr1Wc18
DcmpezHkIkVglIzmnmwFybe7RK1alX9RuNmyFaIHi4lgqQXkcqT1Ema7r8w8cXGA
g2ltl5K6ey4cepOdpQqRD3f5VC5MoUcamOPBYiZTrwWNSClS37LWWdPhPn7g7BRG
o0AE0EpwfsLa2Mjt5D/h5Jbg9skak79l6Ia7iSMIrS/MXEwtoeH2amgItHSNDUWI
fsZH6wVPVJgBnI6amp1UP9+NAlfrpGIf8okgdKkVJUX2UYCsBChcOMSixgiBt/a1
+JHTZj4Lpgy9hWpr9VV6CoE4CpUW5/1yNtXIoR+rM2dW18/9MGtNCWBboThZAqsX
kyEZiaOYPG9aO2qr+Wvg3cdGLsoiXkLTDGw1vk4bzjaQRe9naB/jjDQmTpGfwTqa
1t/Q4LY5mCYHnkOoJqGTOsa4Gbm54Bd7rjZ8jkvZD1uBtEohOd8QP/Zd2l4YXRnu
PdIcvCJ+t0DM08ylYcaMIhuvZ1lZFJrQIKz3ovuPK466xzq/2fZEeM7dF9vkpkcX
pJRgW17uVrPKe2qZQmmJPtPmp21EyZfvq8OmjwF/NbDEuLCxSQ0CE6CqLICGeGyd
6QrBzNvjWwNSgzykhRMks/X8Ha18DJ7Z/1Mm2BN5m33fiadM8XYN30YqyDdEamSJ
LaFnXH4ofrSG3BULHm0VKYvMLj16thNp1HoY3c7NlbsiDnMi+U2g2n/UEMTbMlbA
kyiSkvnbHSLAjPVwdjwHRZz7K4VB5Ej3Y1i0oFgy1nVOGSSM5vl9YuHhxEO0yyJb
suSJ+j4j26iDIqElLU00D4wiiHS+FsE0cJ8IH9p8O3fiuQ5VuCpCXlz7yHeBBDNC
JZfkVR5Mx/HV0Lb7tdBQHa651cwu+I63XT8LmWtFaCoHURPFLFOR+S5ZpkFcUkIL
CxJab744cUIsIECzbLS6Vqd5Tp03i0fS0djHz2Izu7McfD3xJt+cs3iLWp9shP0g
SvP3R25fsCOdd8dj16C1nN6sVRaE+xTBJ1HChmOoAACs2BAbQw4McsoHDKnKxbwl
uASIAkr0U+YLkWNQN8fC88cL8lrtNy67l/4fT6IxKl7EdnFmu+xnvJ3Ph89skyE9
IsKkPi0dY0VuCamKO0UeOioHnj/BZOGj6Qz4IYjs9lF2Fp7+YzmwCsjUH8tyz0np
5MnqPZmGAT+r44mGegmj65ychapI70ubZ3vDLtmrXJpyC0+WDMPFGWTFwc+iRfpv
qXOhYXGaNZJqQBpGGnr2N6NVLLq1rcxLBoNIv8eNquyBzf0OxGYlgnuCwQTkw0PW
f1uok4SfAK4ZYAfgbmJQ+WIKx0xEpmOawNyZPX7Ptj2XeCinuqc/Kx41sUyX0MRl
mjtG90U27NMNXJYWDlmoYUYL5V4aD0is4Pm+E/AdnC+fLo7M3cDz1bYUE4aJQxNB
Qr10M0ldLvrbpKIt9SPDvRD7rDkeaAO6uF5JA+qDr1ogumdV5ILi1++X6AL/HXG7
0kKHXy0iZssuYNUGg+zI6GoHrvYgdORNKSfRnfSI6GZikzXvSlL9pF9HkFM0hQuP
INMiTMQc+rRUFPlAwhdYpJx7CZOP/2wsndxeTNliqIMc38mYAkLmwBO0GFCNB9g0
dBToLDeBT5OV6PN9WdlOptrVLQA4GDBTQ2kUxTGU/+JAWZJIlTW3o+RY3pp6lGSa
uOq83t///4415rn7FMw9rRP1O5SINU2hcd93gRZCvTBloEG2DbwtBl++KSCUiwXl
stOAdONes9cHeorpWoGk/ELdshmfLuzgb/vhszXL0hx5+jqS7U0GylzWUzNzus2W
7oYTIvNE44etXfSjNF5nUcAlXimYaf6XewJpSNfcQTDPgetL8E11HCtsDtbqG/uJ
ASa2E1jIeDgbDYW7pdKOkdsKI6wQf0hX6ueXLSCifiZMEHk3cf/FK/bcUFp5SIFu
kInJ+dg7CA3guR74BxJ1yCmittQEfN/rbtBtBlH+lc0hWn5exsxPfcCbFdVZpTfk
pj9Uyce3MDEMZNeyex5A+zeb4zDY0G7qMrO3Shi5lKxpJs/bguTffOp4romJ4iK5
TFr2c3nv2QEjsPpa3EQn4Zr82fF7D2SZ6bZeVJdYJDYBkSxihHkbHt5IiO373v4Z
MtjXT0g1Qg101mlX5K1Q9SUU7exsu8ecvVVhm11Ds84lOqmRldl6QJz3XCq5S7km
K731G1bmbTflORuR2XwT3My4SL0uAc+phxQIOkYrO/nw8HkrxRKbR8VThqnqT3z1
/8cJJk3pT/JDWKUkLnmLIFDcrThQ/+BzePLmO5ZCW2ei+kviLaPC/Na9wfz5XdDl
tlE0FBB+25geggVqGXQuFiZtClmLB2mgwXkcUi3yWpbReR0dsbggc3mX7LIjjXnW
n1x3tt2zSbJJbeO7fmz7yfE/vVN0uV1RHPpIwcUa3oSKP0NF4Wdaa7CUbYxUDXfJ
areDTyfovuRdahz3ksXPqKjKMjWV0UAbdxbj4Q49zyKb4RUyit4IxbHOcw0OgMF7
uNT2ljd/bzSAq7Ayo5XRhC8qw+StSP8yZxpoL3e+jWbquxOwpDbejHBw6IhdnAOb
m/62QVhHTdHM9QVDP+yYHYmlJsUCGhrHFh91BEgl+ywEv1KSfxmfWyY3Ls14mr4c
/IvqByl9AQqlw+Thu/utoj5KateItRU53qGrxWyEajq25HjxtPjMg6WuJElVdCJq
0dRmzwOZq1BtofFbeLI/qOdv9oZn/EdRt86K6p+fJKE3SByfO49252/3jIn7eDuL
TM3kaMXnBB8uwquUlemr9+QImOHHtfpLq7N+xPL3R2QMhlPOpuRVpJ6jwiZaIwqK
fdfLHoiUe0xuMRSdYO0zBo5f6L68KHP5nvCsskmbI6+jy+jjCrXpY1mMwV2b3lOl
s0Mufl6NbtrU10cUQcjeeaep9DBzbFhDJEFleALSiXhLyVSJbuTmHgzN0R5a1GLZ
LfHq7HQ08nJV2RfDI8AL7D/OGXxv29rEAP4eKt7yplPnUxasIi/ait6u1Nie1Od3
UjnaAAE1gmaqvzhzOxe+e8Lc7Nm82zw8Tfv/3WYInoJBEYokIJgS2NnNGuOD/j9U
YQx0d6aQodlWHmocdGxQJPPhBJr+IwDzEWX7b9ILXoYtPyEcJNmmho2Z7jRUm7TR
rSMVPy9Ufa0+t28k7HCvIr3ZWqSj05eeY85l9NnmAVrP701Ww/pgNkGPMeUEQMsv
FjzlVPfw7VWo5esFlJYJBvF7EdzfRaZvD42gmZAKmXxUHA2H0bWE6H0iYRaMNSS1
4ENBoQ84244rwP/bfMY0nN0+Ou4jhnvYKlogvS9avWYLVerVvkvkDFNJ6yKRIE8y
x5fjUIiuycXNZVG6jwdgM0P1gur09eItrX2SvIp7L/ESdkDP80JqoRRc8PGrgJO5
07R1kEuxAYJ78yiL/PkbGmiOnGw+ya33nlTzVKEmJZukoTl+kzW7c4fNz+qlqwLi
aI7TNN1wgNafqcXab0c4+6mZk5OGmdnravx9IBx4ML269GW38jE9Fbtsas19meAa
GWuVSc5xazwwba1rOtQN6maVlpnwIkTcp2gvg6haIbzhRMLJxH4qaZDhuIEZJVum
4MEa1ErTg4ORQ6cKi4cH6fkabbshM6QsF3pmIlqLfCKVMJuuAma7j/dJh1DvCYaW
Vjjxn8KsjPSJxuxiEYd24JN3oM4Z98RGIo4j71vBv2tzHaGJWT46O9cO1aB9AA2p
hSmpC3j997s9CatJ3wxmBr/Fd1jqSyjEhrtCI+MxDjPItVcujMDvIBS1Qrd9uoMR
BXMUNoVWXeh+EnTSxxzxGZrz+YRoGREDR5c4me0m7UK0CrRkbldpBaM0rtKql5Sm
BpTGtGX1PoS7rEZwcXg1WCBkPz6qdVka3Visq6Ym8zyFofEFtH/lUxwUyyGVbzUt
+kYvHL3z3WsGbwqbuhzcWXfPXn0WNdj8F363Hu5gBDJGhFFHENjEm/SGVJ1ssds0
SAVcO1nuKX4u1v5atCeq7D5PyEi8koTAAEHye8YVdKPliVag8iEXfsc9HZqjDu8Z
Js1uSmWRv6IN8utaGg3YM14y3ARAfH8DXpLA41K6W5S6cI8MzrMlJH0gtorMMspz
dBrcTcu7eP2/cVfnmF6tq1FJeRc9ivUFfd9ZM3LhPCIHOLkjy53aVta90XCUs7uX
uOJCu1bScCi2oo0Djg/TG6uGrChTD9nFC4ptNjvz4IGiaEY5SpQ84/1qCwtv4zNY
UcYvXckue4/IEAcY/EA79yBHqTRXgUJHPVdlpS6RfXziAOKIczuLlM/I7Cp+whfY
byt7yAfIQDwbZSrBkGmoIyq1Gz+telZe0J3QYBnMBXW3MGcHiNHhl7vtKx4EmgYq
rf+mP2idJNRuOdq4zpnjCDD/OccN8XLZLp7iPgtkCUH/pXIc/1EGykxua+B+rW5c
EY98NKcaAuipMukj4md4LrprtlaI/uV0jwUOsQNkWpIxnfYEhKPm76jRZ5F6YiH6
37hl175IpOO7Rq4wuXg3EL0pWGmE0DeR/ChKk2VyyWokmSYcgpjBPQVopSdEYDAR
igU0Tc5cAhwe3FcCtzvELVUwyh+3j6DWSfbXqT0lK6i23/VBwVqhHhwyFWLV++/D
1Jagx/ii93Jbbj/6HFGt4oF9tprPITxMsFl6160hztQm5VlWyiRi0tLdkAOeWMj3
zNy7cZidljqWykdkx5aNJB3Qc547brIE+FmYKYPUu6EU9NB5Fhqe+M1jJFb8F4qd
Oi/SO3OkZ5sjxuLQwKbUWVUkBDnhJP73D7W3o0p6IfPQwvP1FB/yloI9P++gU7EE
9kZvUG4BCwbW35oVkLhGlCX+15y30sOATlshW7rdqiGEvJybnqAj3bsMs3+IjjeL
nqkwCRmEsAgZrn3ubAGlzj8Rjwy6rjlxDE/swZwT8ensJx4RFDaSuLgCnoDpomiJ
1RGeHix3gNZfEonM9GBCi4zW1Il5IwdxK2cZL0MmFP7Yv8CQheyNyhzkz46ZnEN/
NQcWqjPJewyN/xjVFoVroDLFLM52EcQwh2JMmjB/V2v2EDmqxjhyr2kguWezhjh4
tHLm5eFwR6eZCwzkf1wViN7q2Spt1FbpS8K8itk8nmggY2AUHBUAPwg3NHI4KQAC
zOUU7Akbj+wYyYgq09dsQFDSDjB7j4p6q+rMUJ6BYmawD/QGjD8sUvEgG0vb5VDY
sWriiDnRmJj8BYLsa6NVMVYWtiIi1nlKxJ6VKyICNcxh6OGGZgBlcAUSZD7GQ8Qn
9r+9u6JZ3DmLIQ179FKo4lyiiv/0hKO6Cv0GagbW0JJxvCCTBRYj7tZUEPyPS4GJ
FXkcbk6UGMWaKDvdhyP2Y2fkwpaC9ed7ilOVntbcX8r00q63tJbqy92G5K8gliK/
boThcnCEmyBa1LU+RtTiIu+SVIB1+oKLZsPLzqCkFuNFJ34rFn72qiMqE8GvBN+e
F31KvEutbmvF9sjnZRATI+xNoHngvVnB1ZJJjMw3+nK7jkxb1JDb2JbrZwyRi5nC
WL5X3/kCOV5bO0C3VCF7flHJsHPL3vUcZryB27rqTsa5ZOCCHe4aFbb5+TFry+E2
l6FDczx2oXW27+7QoFaqw/p88Xat0+80AuUAKqPpibVaQ5MHh+iaoAoKRRQ0WRPB
MtlIxqYd6dpT80dcOGPKydrgu17EzMxou5pq1LjGWcxGiC1e+DQYL8ZD42zhuupi
ImOdago2PcpXib1t4PvibJWndY/OE52ng0/LQTA/cEU2MRY9b6sVfw8KSIDtVcX+
KxYixnE/q2VVaWOMkWNl1ZS1IVzy/kivu1ral4OQFY9UqPcxQRgw4Ilsv9fyGF7x
qposw5xx2lWh2B6x9St2PeDDUsVwymfKaevFESrSwVj+LcRjnj1JSZXzoLX6cSJ/
tFwryX+GAyAt3MKnq3VUudQdzfQAtYc+AhzYuNuHLbXnLYrIQ8zc2oVPViEpIZE0
ZFNjI+NkeKnj77BHNpScEAKnsU+Vf0/RrRHzKkMSHiGBufYwyNPDrQbDF3dC9Hts
7fXrM/MLceqRcLiuPflqLJQqrFXZdRWLLOsS/fKwTt4sveG3IM83+XuOVClkE1QY
iJsXCbpLL1kHh5p4LmbsBDOrSJVnh0h34Iv1zZa6/PENL7ZaSpBu8bp5kZAZacSg
QLsMtmT5GJyRGbdRh5yMUyFdohML58w+j1tksiKeJY+l/ZXkTuFxRaNtNRBsHoGr
HZ5JsDy/H3aqMafEyE9pv3FWcot4IAzS2nR2FXn2w/UrF0UDNs7bGgghkE2xSVJg
OJIFWauuqfF863uJyaRxHoOLrXiU2n1C1BUzZ6sssrBfBrSQF4vOdrSn45gMuUJY
DfCrv2cFXwfV4IhtBfv2PVUEUu9joaxYfRjqiBfgJEwUrVYMQvurbuXaf/fwpoOP
FLchDsbjm+TL9Olika5WoHFFdOYkGfBdby/q7D7vfV2PiCbs8MCabOE8gl3BPGZw
i051cKhy0JvBxAsGSJ8i6VVwAubbO6qIfzxCP1/9OtkxO0Lp05J4wp5gWt1gDGUO
knVUMrm/wwMqX0xL5xx2qcJdEIcT/u3oRb/Zhuba+t25Jbt1BCgj2lOEG3ZGtBOQ
nL9RTvZfXZ/lfUcAtaDrOgUV6bxjXsoo6xdoL7o9t8wWQkNxzpUTg/0haq33jaP2
3skcdXpFlNs+IWotylQ1lRPW78H2sDTHgL203iDoaVQ7XrfIH5pyZZ684lz/G2zR
dsH6XA1BSw4rg512xWRn/QVhFkxhN4TLRoZLIWL23RMTb3nGXzhHipZ6HvH4bzOK
l+UpbZmNlvjog80eV0nvSfA9fjihqcbjf3JhgwETIaQS7U3uy8nJ6FcNIFjkld5A
mQ0FA3iFLjPzXFQqvtIzYE1d6oxIunCQepNqRwnG6i1DfRAQNFOCXJmkO9GEV87Z
0twV9r8eTOd+XqtHesfgjCa5u6nr07FSAguI4Z2lLevVqS7+3I2/PEsRmfx4lj2F
b+R6bIyJVE7VcajPhM5cC84NI6N7EJe3YWeTxbqAGAijIxrWMSA/VPVWhrWeItfY
BWshHukLMMMJIS+P8XmFOflk5gAfm1ceS5fum/Sf0Dv0DaTjsZAdHehRchQMSLw0
I9iJewsVf8XnvErr9AgK1wdElD4TEZos+/jfJ/hGGK77/FZKaMhVPmw+rnkzV0PW
fZuKx9cXp+L0Wq6kedgTQep/WUNg4oEnFaCmU2pTnC7Gxh69O2kFgYR1xPx3vd2I
ifK8nQ4D4RKJTabQC0JU6s7/ofPDuPZPeqso5AcR88yp9pv1iH1sisZSVp9J08u6
2E59Sp1Y2/P4i/hljTskICIX1oMLQ9Mhb6nKTAYLcnC1N5xbDJ6ve2/A+e79r2Q7
ouDUw4AwAohOX9BZ3U/qzb/ScR+yKAhGUYk/hLXqM2ONiimAsjGO0KA7RpRg6eYI
LV8UbXY1VhQppOeKi5e3ziyEbFVKqSvEZTFBxGg17IVvuxfqfk63F6vQ92omtjhx
lp/MKHjkxHhjVaAZJnyw332jh0Fzy94GdZ1Kvg8QJyhSf1xc3LJEd9t8QFv2Y1dI
AhtPYfBPLFBkcV/wxAg+wyGP4155socfQss95aRgiGBcIqtVvd5JKO01++da3r2v
2DvFd79QB8fhYgn8GpaKx3bhrNL5mVLFSdtcRBdozELU2b7VUftab04nGjo5Kwqj
vg1eHA1oQJQxDPRRAjaZlPgVP6Qtw7NM/JbRboWpfNXqIc9rQUHHlWlB12zrfTos
/cv/ReCA1Eg7X8wir5vsK5yYQzWCS5m7lvWgVqumyHJ75e/UbG5ayCgoZ4jOQjuK
RCeCICwL5WYYmL1gK9O9Nw6oLiXdzJDa5AVWFOFb4IWpIIPFkr2vQk2pbgKg7lFS
66eRFQfxqTYD9RiwX/LDmSyGX86mUyLq2ecxikmNRvmztKXBjKuyfZY5h8+ie2Cj
zZrqe6QM3x7CIfYWAjPkGjtkzQhQ9/93LJuct4ykBEGh1/WBvaiB5nrA6DiuDTz0
U3/u7WxYEna4mlrv1cuP+6nsfxQCuF8jSgExQaRniMYvUmJwjWdNE3Tf6HEvqzic
sD7i5Rrb7vBHE6FOk4cBHwRiBapke/SI14iFc9VVe3YX7UuK3zT3QBNMPerh93hw
8JRug4bM3s3x34bM7S4YRxFbljko30mZL7qmSSjX6kMOQA9nd1m88e1230B12kgF
kCCpN2vKgctXCB//Y+Y/eka3QjNFVZu35cJnyvORXn5dioXVUcWgMxIx+sc26Dgq
rbCdLkY3au9dpRSay3YuA1QYibIlvaAPgWt5IQeYdbbhM9v13j4aJNMikQPoSXx4
oQsldW7/tA+g8HxhCGnRhzzHwPaER9ShG8dPPUH5uXhNq844lLJkYrgPurwSi62O
jueGEyNQ7pGXDcPeXSTCEDADNCRuyFmLzoMiFtn8GCfZyDjZk2uN7URlAo1Ly4Qu
HK3WjwUMSfLnuxlVyirqoPrM3k/E1iV1x1a0OC1ku3/kJJlBZo2Api6MjvdKDpXE
cSuEGshOwjVlkaD2xcG/d1VK4XF20lMe06m+G6cz4vA7f1WxB2/FomBzqk/AN2S2
V1Ur4pLbNdIbeFy0ghBTmN3zDp0XraNBWFhuRYuBJ/4uAfxUkBxkK6zdmWVZW3WW
y06fM4akCcWN27KF7df6xX0E5U8zvDxUKX7N5soe413DK9EvMYSWpSQDOHpovXrY
XpiZBEO4xclrHLE6TT3AaIIAwOpFWgyk8ou1CZikjLnISqC4wW1aIRQzoL7sZxt4
KNatnZCJmD5HysI9CPBulsM68g7d8AGCKqClQW5s52WGtZfgcf3PffKm0KUWFI/C
wdGt8PMIWk5ycT9frteLVYdph48XyQCf6ZnynBrckk16KtLHYtr0Tq1CE8HwwVIi
XBqmo3f5IrY+smm71vMz5beVPV9puBN06rJv9b6Pma5g2u87dvSTHktV1OL+Wbvz
o7kCAhWu9vH0UnWtRkuEsKt+4zPKXsuZAz0RUezYPQoGKHl033mVlWYqgYHrsE0i
pJI6Pvslr46yiQBkX4R+MJ0WpKPl8Ap/C0FAeoG+Ta4zLEsnQLVfRtjkbEKpe9K/
2tGbUBCoswzUt9RHh+719nL4JAeqzg5LPGZK5fYLeF1MEmzcvxW4QuyKEDPm0sjg
Fjk5QULF++ZKUg95LPTHITCCD7ftPQ40X7hBs980urJT38Bkn7r2muyCSkjJTQJX
2m8TJtYaGN/iRkfgLYdz+gLXDnJuEwSphBm57X10nvYi70NIotyx89V3gzHpfCln
Ps0oN8o/a+f3LTGGUawvvuuHMRjKaN7z5+u/n1HQNtv4b9SojRnx7A1rPtgEj1cv
BPVO8a8VhSu54inVqIH5TdCeFPdfafYnGkltLLbC4gHKjVaSLAw74gjFbDpWvK4+
kWFKQTgYqG8AAHiQiMnlIY14ZgOZ4L+sg1J/HXoV6EBtpeRqP9V8uYspLv9JR9fz
vkwDx7woqLgtBSTWBJi41TNZvSn/4mEONq65rAtL2ZC/eRO661n60445vF9pPWo8
LUB+MRoziXli7U1pEBVd3LTx6QvFG+ssH3wGWQ+SzkPewcanbtf7GkbxX37gy/sz
NfZtzErRNRtGqv1LGRvRgBRlqI81Q/08dZZ0YLVPccg0xOx4s3l+jcR4jM9Z7Weg
75bg3lOK7qqJ7F25UuNLds9FxBtSSNPCxMJgzM5JBg5ak1TjF5hvWZea9GdhfIGQ
40LyU8wpZOxK8wAU5UXTqC3DixczOvt6bEIWtQ+Krqpy7po25n4Vd70IlTIqm4qV
nGOH/0UmqzE/pu9v0WUEtrGTYaTGXdvx3FNWHgk7qwmYmh3vwLsq3Kmzh8MbBzke
h0FSE5rBpLYO/9owLEY0HQUmK9FawBDZwyNY4+MRIFbzu3qYAxBTrNrZxCpHXpVa
Ig1AubgY33osPTyzhrHSxA2PqU57Lt3FYG8gWrRn2jFczVr3ugJG5Jc7dxla3Hd6
OqN1mFk31m89aUmwnhpkz2+kfTsXbobDsqok+K6pCJXcPMLmBo0HAK94RyZJmr5C
ed/8dHXUyIHhmLjhMTmhf4cpdZ+l3pYy5fcPnpYY6yHrYwmHD0SbKbelU5SsSk75
45d3TMM5Wth8kGmjFW99TkSRX4i09C06I6sP3jOUS5+dkKOkr7RI0NNFgEIeFusG
0kxVkU5j1e28BNlUR/Lhk1JZ1Fs4hufrD8kzAb4wq1WZ2d0MY6tE/t5TwFuNa1y1
YTfi3hka1T3WHLNGn1dfq+OVuwT5NjJp50+Nxi2SfzUWDc6a8n4F8r3LKtzNwzk2
lAQkZexwDMC4/1OQnP2Pxgsvz/QSLI38rtticcrGdWll2C61BfgXnDZsMpfbdviZ
Sy8cplGCby5taeGd31hM6dB7WMI+4a6kZfXOL9DjBFU5lx31w11vECtwhq+zDWqo
uHYLR0l6JaMQkOXYGSh+nRILoG1prtNloxLbA8iRun+Y/axHskeiWZdBe/P0cpFP
GAVEdnX4FPOJZCqqUiuzhcuzw86jzXD2vYeH93HSV91dwjCILJfc2DxBhmv5tc/D
is9T4Cx1pmLZ/0EdNh6i1BDI2Td65ICvZmUWfkFNF4/OrGKfsp8U2wkaTsbtZqDO
TAMtaY75HhKuU3QSChWMi8atCj4xwn/qy/aNP7EmLoKPPp7kDc9gupzwB1Dus+Ux
tea0gr/ykdD9BSFB1y4pYIuyp9MBl3WxArXqlfGO85OSY188sRpAWOiDKU8h9uhy
F+afdzIznBXNLEzTp/HXh1/AzXaGQECLQhv6p/ZQCfEK0k3Ca8Sdo3YnYCONri5V
tpoCltB1kJKFPwCdt6gg9WW+VXUi4g4+ieRF1AdKy2paLah1hy5ODKCpQdVVjiOg
RnXZdIYTbp3Kap5FpinKqtDo0UQ+bcFMcAC818fT3MQri8snwwNUrOP+icOs+nZu
L+OzrTU24x4/oOqWkMh4re5qGPDq73R9m7dDNOxVQsMSxtpS4QrTqPRqmcceBN/q
0Rfbta4d2ax+YcC7KbesLkIXqcVM/Mna5Al9JN0dt8ifd5PVjbkZlY/wEKvy38n/
0vijLpzF4TC6wXFlPPUbgdOKXP+WotxB8hBaZSUlhQDh/QxjCrYJYqJzOi5efxYU
djVTIVRbAW696lLrEajwKsb9XgRMCTcJt7d9LIxmsPUZW2wIjDdUKLzz6fFB1oKo
sh3fdk4gbBz3KmDQxAl6RVuPomLXavc+EHR2o3Oi7w5vc7826D/Evjj7tGNlsn4t
WBV+TjNSNuS3iyYhnD8iBXO0KI/l1WwlkVfNqqlURXfkAUrF//BWc01RcOskD7by
xynMF3ERgkY6gTCGQV8S090q7/HnwkPQt9meZ8ea3MPoXT6CS/Wv/6PScmM4K65J
rcpRqNAJwCLBqC+jNBMCSn0WX4s0sKzYR38K2M9gPnS0IMba/gtqTw8rgMJYh8q+
WqVYy2TL6adxWvQ+RCT10fS4Gvzsub3sJjc+Md/PdrWiht0rVAl8tkqyKS1Zgbsx
gU63usEGUDFdlBSyAc6oWqNvd1hNVeYWOBh48nP5NA3j/1KolIoiju5tfQPPWC8Q
QxiJAXbhc+M9l0pEgiZs3s11D0xtAszEkuQBH3wtuOORirvPREYgRD9j/oUGCAjq
3Itl/4xyCRF6Ej9nmtd1Z4e5gt6s4U16ILH2528c97zxLU0BRpKn+yd1nm5jriEY
KqKV7mtkuLwQzaQD5YlQnmfqhmeJIL7L6lCH1LlqF6jaQYEVsHkeDwCwlXybkke8
TxYgIrx7YcFcy7L/EYt//MvllX4WbCLYNl9Nu42EYKnX9xHQBp19egF0zz4DwWBG
fnxXAJ4FvHP0l/xQkq1XWJdjimee2bUQiNnN/e0YF2iw+BaeRzMRehM2HuICaMzl
uG8T706QVkPCWf/Rq2OnUnwir+eKvU3g2kG3sgPq2+9v1OTWPSUoakm+w1Qg+gu4
f3FSca/c8NH78PHETWQ0/WUiSI/iRZ9ZCH0ucZtdWCmElT4zvqc7V8L4gKmq6DpY
Lv/4Rt9cOAE3xT1+f9xLKqLH+Is8IYNCee3eaFS742h6f4ZBSkkcxj/MyIfF+FW+
27mQlN9ESgrKvFrMffzctYw3jN0V1GsYO9aboDTRVV6PRs/5o8M48GgyBnmdoG7D
y1UXVBhflloyPPqcRFSuprhPdkoRVperJDPb24i4jPk/oAHsRbYnMQpIr4GTMO4i
GQ/orswQviGAp7QJuGY4/u4rPTMLvYTjtJ8cgBBYQqtUJVBeTtQLirWo0GBW/J8W
l2RMy5fLkdnGSdodZa4ypmKmOPDNb5x4xAVP+rd/DkM/WuI9bGRWilsmS40H+G+U
+HG1FRRjOBWVil+eSJJlWHKYYn1fDiT9gJvqkYMD0d6E0QV9+1dqXXLlJW7dQ4U1
Kcm6RhSO4+ALelOqNtWH9OarXWpDikrKDCR47ZMQ+se90Io0YGR3vVw4A7hbrLes
tkU1uAJ8Ibk0DjOCLxaka93cjsDhBLb7Ypm57euIcotKKYx2rKifkqyplVGAK53W
RljuQsX2GoZNpvBsh4H/PJxaRLFAKkDOx7aBm/Eq02KqOqp9WXCU0/R5bMupzMpC
ZiXYutRFNIwxOSeUASINyTl1/+Rv7rnDnPDeGimPWs2ZSmY6WqRYewUGiVe8RSrg
pwNNJ6U/zmULOvSrleAyLP1sW7/OAYrJ3FdM3TLfyPExJ/nb7MXKtmRHdnmaVH8O
BYA+9OfuXQKnUTtj3riKIzkryQJjfFBbkmwIMbReMGrdT6sO8JQ7rZ82WYz14yoQ
T3suaovysQN5sQZSbG15vBXY5VG7BGskPq5yWt+Vk12hEHttL4EgQYJsWLwKxCWv
ErvBaeix3Eq302uPfmStIz3CoWdyC+yNwr1lUU7rbzvDjp75L9ivqWLO8SPeLqmP
KFsOwxqXQC/oS5s1MEDgFgeMHwXo/cD3CEcr4s0CkUuU7sGHgvdP26DdYbt7zwNd
288Ii+mfR6msQnHgiiP5xjLthwthONFQaj6FSVUIhU1Td5aUpdQfMh5PfarXGYDe
zQnvQdr67jv2x23WaFs30/RJuZdkgqVkExwkBUpch5JlmDTSUQQSvjofJRwrEXcr
Ge2vRWLyEtNX6h66qaCrHucIjfV0WPJYwjy1ssA7Nq1/JnUqRRkq4BfvmBjg12ah
ZSG1hQ5qd0u0LxVQ2of4/Mh57FTYWWac+mNU8510rlZqtgfGr2WJAkKVDPMTLKVa
//i4HrZHxUHNubnD5L9K2PyU7Q2n69pOvjlevJjlTaTRJsaSuSZsxSdTCynYUC1p
wGI18l+4yzRoMJ1V4/FX30nJhd0PlWcTQ2Rj1Xq/5+pk1YZTFmy5CaC6Gp2gda9i
j8G88dW53ORT4ts6C5grYYHw814HHwOwP8+zbogdkfn19wzE2/1oExKxlOXt82Zp
+4oNEvLrHIMBBWRK2vmswETJIn4UQ34cjIn3htkwKGmyaQ8H+Ae6ytJisH77RRK6
GBV+OFgoef8BxSDWdgn6aEfmGRwh524KvqS+BGi7QzgG5meM6aiepVDC2O2eekC6
9xxg1T6RpwJ1waa98VOBIreMB1wGTjuua0UulPFiKmg1vTPXdg7J/SNRo/cKRQFR
4TNuho1hKdyOzAe8qVcHBz78f4mrYxUUFPWldZjJYWAGl2D5Ezg7rlIXmMh+d6Le
eMUVUeoqhWTyMWiw1HS0riyucPWAAb5vee9xvYIduF09DXE/p1jfyFKusCFgiPfZ
mu+QGd3T/K7PECU9rmzuvvq1Z1YqcFYQaFAA/9mjuy0fRcNaNtoRhbcO1aqpd9JG
kgGsi9jccARGiB5vqydYUDLQ+OOv51xl8iMUsj7pSo0hLfJFQgG5flKbAhb9owa5
TWnP69n3Dk7iDPklw6nUxGackV5UxE08LY6FV9mgmYwjcBSmi3wFOE3krGt1yFav
CvzMja1Zo7UghxQZzDrIqSmdPpH+sETVBqALLQ7EpFR174Yj2MKB8jU7Z7RJpm/m
oR5k07AUnZ0er2A0G5/rUjyR7hsB3QA3KJGGt7gubmAZULOc4N0NIf2c964i10mM
eQ5Cgn9ndRPj6lFeEEv267Kra3Dmx4neGrj3bC+4Nj8AXtouxJYIazHgIG40OmOk
4PmHm/QxQpMqHPqIs5tpEJOSNRwDV3k2JkQf8CSGQ4sI7ssCOgyg3AOZWYOKCNlR
/kknkQFWcK15H9OTxN1lwsgubg33yBBM7vyec8FDEX5iPpRCWrfWTo3h80wzw/8o
JPuxEwRDzKZQxEtSEVKBxegHY9PyEwbAm40Ylym4vfOFYV9nqu5m49mWYqUxBWjS
wJY9x0hVw7QFZOu3vAiFJIOKQL0/cpG2yR7ZgVQPt+Ai69fcwT0euI8SQO7oXoZN
PZrLcs/1PwLRweT6fN44+1Bgqg05HTgSnfbVLC/jrGX5Lq3icWnvFNZwTHPRbiRq
wDB7hILoVHQwE6kOr+n2IY6lTzPU0spMPZEGeYkxCbFjk8e4buEN/hLEeZkwyAGO
mS+5+H6d1X3QPKYWf1niYOPSl7AlP5EIGfETE3OTVcGkh8LpGS738V8hHMRI3guW
io89wOR6YKp/Iwl0hlG3Nw4BGo1KwJWFF5HweQoIZme9WULjGHPwi7qhyKHkSRK7
6ZPGGWxISmC2RT8Myufp5+K6jLB9GsO5L7XTMgfb3HN5PkLnSp0acgj/SQJ3oemj
knR2yak4BTljZBedOFP7z6n8i81r8Kgkth6qKiGbUbeZ7qcYI2pgHbuRWdg1NHPU
d8O8XdC8zARPV+Rkpoyc3Pg1YbLDjCZwx5L1X9sFxOHXIyT5/GHhsUy6TynYEUZC
1j6KH5dcpCJ+LaaNTiVnBiDiQB/BfYI87SlxVUYUZnJ3JlmW2xSX7pUS1rqLL6Md
v3uT+F7a+ZB9CKXOvRSv1oLPuJIlQD4i9WggVfxWBhzrdArzzPZ5qz23Pw25xtD9
qkpx9EwBEcYvgcsdvcEK/bPOj7ewEJKknw93fwbv2j3LhQvZS3W8Y5lQU2OkXqcG
uzf7btTIp0IAhZDB11oKhSVmvPJCvfQsN6MykDz8j+MLdoLBYh4Naa+Z/HZuLeGx
I8I4XSdpuXLOJrjReCvIqIfOZ2KS+tqvZtasgtr/qG3C4Gt8WVc0avPyYIwglozX
IT4y9UbwhPTOIwKYb1nsIRXFfh8SCxrgNCavSPUhbe1GJ4lYDXHBaA9xhBTYb0rE
n3qI8DhRtxuH1uSQnCBiJoYyJS5K9yOoRJWaHESHogWBEA/YIFnZRoW0rG+P0Xjb
5hGoxFWP6cCdP6e/l2zVqrfvuHoD/r9AFomfFHLCdNLpu1mWAYf7AdsTomzyEgUC
wgxOPmnIoFHZ1xV4QM4UlD9JhK2xfpcpFgn1q0YsAWvH/E4y01MSKuHZyKE1hF1k
RBHmtoic0e94w7kJ/j1SzSAoEuIGS11UqovF5n5pKei3qMSEO71hb/Q4ftO+kGcP
wHQdkoyA7+x6+IcRroOuO7gUdLgACFZmPnEKhMmza1DlTLZ7IUNb1wri+1fAYneL
gtno35w+P36JDJeIsf3L9TpsD/MOza+8OZwWBdwujA7WKKutKrYGQfwetFlA9PYN
agR92eEOQSDHcvGT5CB74+z2DpAF7ewROujVSRlB2swKvTv+V3F0cnh75OKCrqdZ
3tIPr8nSRYmsWtkXnDjeidL9pbaOnRZGy/YeuvyyGHEY2Laj0kQ0jtPxlur/lCjr
wRoD9pBdHTo9UZxvFzFkwyyTqMLrf5zZ41n/34uAitifZZwulCEYUNvZAYv70cDq
n1tPMtVw4zGAwOz+wg9M7DtL5uOQecX6D9fCqVfRHukFu3fvXtfAxbFR6tJGI4Ny
sWrzA8/UP4r3t1hcXb3TwpAV7b6xC/4jFTwcN0O9hNECqr01+XxSA9cGj3k73/C3
oiEq/28i4bF/iCcn+V87re7wfvTLxIti+eviMpn0WAUtehh/qCbpBlCvloYY78+K
T93qgCOKrUUHxXUSjuayI9RqSEtTkxowKFmH32ncz1IcOigAL8YSZV5ZVcdbbhrg
mo6uNEruZD+ZlM0Q4IfPGWUBLQYnyI0oHb7EBHmDRV2AXk/ToRxlVezwAgn+aet4
f/KHvQGkDNY5vYX8SxMB6RM739I6+o+v7jBp8ampfokOnyqNbspAYMmf/kwDdppD
a6NthkQlNrhSvJIu4G1vCevE0vYmP5Rvk1HOYBtjUYu9H7wdrjXFcGt7QvucjqUL
toN+PlweEmfvN9YSQAXsE+r0hDXRdPCCRpfiRZ+Y1Rk2p/0lQ5HueJDihUGp2EaV
IOmMbDGRP34ePQPZJS8PNJxWXYrOFGtezg+fZwA9TdJUwbM6MCyBt4WhKYIOhPqi
3K54rIC/9++dGaCyfSkbOsbHgXbSEtMjulqcZycouCshGdLL9ncjk1iX0L9VKwkA
hHGrgtsDhWzR8/GVJwsMBkhwiC5gryy0803ikj7U7rBoUQjhdGdJBANeW0Eeuqa0
tjP9Rx9Dhr3f9Al+ehYQo/CozNvWTo3QMhStCqZ25X41ciubMk2XCsMRCRoAjGVT
X+XPVDRSaqub1kGydJEUR5CxBVlIxK3E18SpdJ71un+HHHuL9dE3Q2+XIApNdtpp
bomnu6Iy2L+m272mW7V18Wiz890DllboZLLi6EQUUM4jeSYfKOfEFFCjMQ9nT9c7
Dft/2AgmrolJ8xHN7yb3XcqvAWLdscDC62qwzkBb9rj5rhoRq6DMuYcW4dOMMEq8
hTBgYB/QUFEGCgnsnBBWpjxpFX1+Ons21yybvym7WJNBh3CQDTV5+mUBRihqHtDm
ZrCcBI3DSM33WJIh7l/evNXZYq4AXmf4qyvSop5iZnIgFdEh/e2CQY9J+3gQ9kJ3
7L2Xta2zOg5X+WDyGJ20AWJO8dowReQK6FXAEQThPyMZf2GypUmT/sQHoX0ojz9g
DELFRfHEpWiYUmS3eAxXkgjJXw8IGmfZ8FJVwAzKvB3RFAbt0Q+LOkhcixV9/FzW
WgBf/Kj6SPu4+PibAAJDqQlLcsFpHyjv2oUtxL6qsP5N/IEofENMmsgrOBQXB/0i
4dpUYJGN4Ljw/sqpY8mDpqbn2n8qqon2vLYuYS/pBZKmSspXb+FLXx/8MckMYBEU
GKE2NcQm6THbmZd+l0K9ffEpe1UzBrVeAXIpNCVLERDp4zQO9jp3JhGiDmpiBlq9
dabciBCzwAQIulLar7Nen0j7OX8vSqEfzPmVX38ywhqDNouvbUo6dbIKBCe6cOYT
F5eCMVosA8qvlHe9c2FidY6n/yHE2EvvBSlHkMN6q9Z7V/esmZMACRGnlvPKeiF6
o51alMyfuAkgr9dFMRshCRBhNvS/su7MB5QDnL9eAcTE6riAQJE0VZ5xMtAbg+xh
AHeTq2s5f5iqJc84WtlF9gl0c2pID3JWPVDpIiQ42W1Qf9B2QJjZ1ycrG6oIG41H
tUlvtq+Ixv/Z+TNDvPK2o517k1c3LrDrSgL4B2YLBaWQoHh3tznfh1MvJWPlQbVg
xlbxSZWnBgb9lslvF0ocHSFrQOEVsxJchh9nsJ15GQ/yX2DzTxeUZ5DlycCedn0H
DmDZMhchslEc4MNEnX19nBu06m1Pr5hUtjP4Th/UstbOmKb9RQbEgwJEGyP2IgBr
PqmjJ9Qm9Fq5mU08ReQ1pNP4kNJlp5xdDti+llHqePzjss966rJpLfAvfrum7E5R
K+x5mPsiUNciBOwI7BH2sD9IspNNymd+R1NcS+PnKUkKPC5I5qYqVuxdPyU/hhfg
GNruG5hbJqXtR6B9V23dj//8uBvuFYi5ibvD+LJ5M7sIwakgr0ggH5Tc4PDhRaW7
84JVdM46B7Q2E5odVyi1bSEjFP+m6qPVc49EXwUzJOdJxzyHTkxjJdGxK6jXjhGL
XznFgYaBWT2ImiK+dMQJHs3AVbfD6DbDt7JnZuJUUGHfA0M1WometDeh7g+yAfK4
l3VoZ3qQ+nceQDFNjNmuLahZex3mo+WOZ1/rcM1JwvBbvwUj3OSWxO8RgypTnc4u
+uc0iWKsLeW0GQO1jHWT+elEIabA4YLEBTJAFJuMkf1tCcTRZedV3OQTdbkkSvhA
aoZykeghSoPIWGn1eW5UUg8uabRg9Q8JnVzEmDa6ktbvjL+LAuiqskF2EHIoayUt
wxU6J+mtZsWemmIy3W9eUHgdNo8Qfg3IXY80Ggk1A+/5LtWHLoxZ96Z/KQIGm0Tq
eoTvi+eJV1Kd5z59MPxseybsqDKzJ2sXIqgwKd1vmQSGN6N+s/uBg77nsOlkmNfp
Dh2efExkXmYV31oQr4x+fZ/Vwv1OPIevSGeZNu13E4OdpcYs8UR4GnnhPJT0le2s
sjVqBP3JNczxuH4iPRJOa++qz7QQ/fIOJAHdhI5EFcZJ0GAfd297rjNblK3ksOww
ZFWgmn20R6I5Wdz6hpSC2j7kvEgfrX/NzAl1GovwADYGPU3lqhzzqo7LRDMy4OdR
oWsoUc1/uVagbyr+mU47yu9E88w7+5JOfP5VK3ywqDvgGqr85j1ebVo9tcz56s8D
K8nD1DxWnH9Lfc+QTIZdcmxsNqfDtOmNga9BhZJSWRMQMcfcE8vSdcFzKDTBCxuY
+j9lBbAa32piOkG5n6Azv6S3/UQAngw0ty0Ibhd7a6KKKAAspjxw3ynTUD9nxZOy
NlxowzfAIyr650X8XPH83mL0p9X7DoBbRFSqHqPThex0eB3pFTYQJFE66po9TsSV
hQcYx2UWBSb4aObtazhQnXT7zmaSviPPl4ECH5lerDnyICATZpezTPl1PPK2XS68
32ZagpniXcrm7fwIKfPgY2GyDwu19Tp6aY5tzp8r9dKyC+36bu6mCH6Kp748A+dx
LmFllMW8HBagniQyNAjuc1/xycmD8IayyI2Mg+SEfgxYyO30LqjoW8F70TrdyI+u
M789F5r5SAET7v2swElh4yEuIQaXakRoOrQrZD6jXlmapc0JlwF5HeWkSw8eMPSO
j8zTV77833oHE+gKQeFwISI+s+BLQ3WgvV0499lW7s7gDWAUAf04c5vtiMV1eWC8
Ak+zV65TavQlVbc+/Gt0susmRcIItlSEakypRd6aKUCgEiwy39t1k+uSPxB/Ml/z
A3yI8fZQhu78OpEx/MLWVAzAbzgv3s/eqGzOiACikaLQL0BLqiOGVEaW6d1hxd/O
QLpPn6MyPSMOJftsJ1N36ImPxtq5x5D6q8Fa8CQY7t9qDWKKI6QpulI8NmMc0LyK
WxtnptmKwyZM3XXS/HoNm6nVkjiam0RI209VQmhUruacni2ba/GB48eRk9TV1VJE
KikpkLCoebjJwgCM9H9egCoTzFYynBNFQ+D6uvqQ6u5lYPwDvhoKu5yd4r6cho+3
flD8w7P1EZqcmkD4j5+M63Tf0xzwKHQ4fea1q4PLFJLe1MCfUrlnyexeq2Y6Av0q
UxuRI1TonkpPT1WdCzd3fGirub1Shoh2P6Xf9Mi40Zqa5uct95ms3ZAjTFwVPnU6
DXEMxkiZEztTcI86AVqK5ek56gY7k4tpgh5nw8NRGbvP0h33JYwjjBx0AILTUlKo
lgDfww9yr3GKUBkhAsf+p5kLYZh7WqeXzQCjuusUr/ht3idwJPDA4AT5KdzzxtIQ
KvQvCsUz7vVljita6OkGpbepMZdNXX/YPeiob/NxVhUVlVVsFF3yfgP+v5a/a5Df
eIyWMW6R0bf7mULBJwBCV1hDXWDOWwbuQrIgwaEMpew5gd7N5K/qMSUGxH/Hq/cj
vkvGvo2IQFWV4KSdEKcgq5ZC7gh0h18TGIaBLGD5c3hAONlWs1uV2Re7hEID1db9
qXTekElbj1xwXYSeCSjwuIKSOKZqbLVj+kxLIP1SxZHwCfGz3gu5VmJN/d/epCW+
xk6j4wEzvDmjNFWt4uA/T6mVtPirkmRB7GxBPBpV4c1Zb4GdBM14q79U7SBKBm9T
vy1rl7VDdFlj+/tVIZGTAvuSxp7MPD2dbIJjQbZt+oNj/W6Gf69nQa9YNUcrpRsP
jC6cZTw9tTojpDNOr/2KW2jvd+Kj7CGsj+/UJutREfY/MwR2Q4WAjzI/LRK2g02Y
nPpYJle1LaQmegWVPDusrx4HsJt3y9YLEHG7pRwh8FeoBFxfAjuasgQw6ytw2L1s
XoCReCk7CP0NKNb8iq+HoBc+ooLor5wZCglVckJuWCbnHZ/6HaTJkt12yCwAU3u3
+0bVnMdSGZzL7apLu66STu0TQnEzeiYwz6OjxJnj2+3uxrBzHcw3VTaIKzNEvMpZ
Iga91nlky8VjkPt8Gtox+5E8e90FjVYZ4Wux336bbII8hY4m0zp5cIvDpw5PiERs
Y0afCVRI30yAiiYA5YcdQqVicF7zQdok94i2l0SIE0l4ceVASu3IWkt/9RBDmxKN
Uf9Uas66y4VVpEhIX4o0oqNOS9AX+Gh4YmCjV20TdLUP5utgf3mzfabwCwnvPAf9
u42DQorkivDZBvq3a5mnA4bkWj7kNIgmYvXwv2kJXfFTNgZ/eB3zLasxjI62iVF1
0s5hvXf1N8wsCxWu9Zju0RfENchtRgeCS8nIbkn//vAiuMf4Ds/jcFUqkt0L7tJw
7PHAdZtKkzphg5wLSNBMtW0x/fQSwUA/1u4tvQhC+3AUegLbUg9Vk+qtjpAJ3fUx
IVaNy5sSKH/Aeg3lQ7l7C0GcsKqeoISI7+ClgIN9DbrJEmiNY8IEDMSTQT4Wh4lz
PLyhj/pPN1IHoKEHqfIGXjUdcIz5HwVnvQbQ4rNGYsv21qyVtbwwFH48ZqYf08wY
4txO2zWfhHnyNxB9NDOZ32obqGN/7m6LsbtJem8Y4niiKxalBkBZ6JcARgiBI3We
j2CVRv0FcnmabSIHjEIZ/ePNBAUZPVloQNXIcrc/3KYVP9lc8wZ+QeE6jWL6MZTe
x00QsDOSDqdxEmhTHo34EzBla1XmQOO549LHFs9PoLx6DtaPoQxfSIrTGB0VDe+1
Xs+X6QpC3AP7EY6J9WKg4jLu1g6aHhRJy03Wn2Ro7AcOFnBqxwkTCV0TQ9XH6Ju/
FDDTfHyzU915TYF7dl6J37/OmxSyeKVrlzpOrBa4mvji+PFrdSEXUycKOE0b77+T
X/9cNLq7vl1GUCKhDQUDJKD9o278nfDf+0LiWX678b4kjYM7D8Ap/KkU9A6YAR8H
aJV2EE1aYC+4ex3aQ9FNp7aXLwzR01l8OKp4IQ3zfDepLF+ZQwc99AcXrJem1f27
aAbuqW1xA3EoTyTk5p7i7CIxdozFrUjdvRae38lyTlce/rLwRaR8YuxK90/FsDPs
UO/tW8ihTXw8vNmzQzgAEMmntztc8vg9kjq+9NQkktKycfD7wU87anuinDqWRuJN
/cKaGIlCxe2aMTIcq9sgoY4IZVUqOLD7tUNcZGYGRJ0dLjZRaSDXdBgRXEaKp4wE
EINQhHuuZqtf0SA9Mgn99gdC7vY7egCVby4+fA2E2sUn3KRDvD0S5m4Df4+sHvxn
cTI8bUB7LwpIRigBSpVBbscZHrW5tSKuoWycvLwfiSyqDHsFgfS69f9Qu/fBAU/G
yzKLtrGHnBUQrFevdwiiz7mOxeRDHOoVPFhMwQZkpm1LJQXiJxyvobYX+b81/ZLO
cqXrwMO1qEqizvi3gh+1ncsreDpfI2IPfO1e6eK+HEUJZn8rs6Kes2imFndjA0oy
/8ppfjo4MaKyYe/it6cOadxLdpA36ro8Q9lynK/njWE5Akwv2Ye2yKeAYPDwz9cs
OFj+iaB9sdG45y6GaHyrAvtv7DBlD909B/VUuEB9btbV5Mifc6fy87FbhbM7zkDt
lEl7USx8QXhVTmbYNkYys3FjITuyVs+7xuNJAPbmgb6uN9iP9UqAYdqRW/JZYlUA
GFQ0Nb1NlOPO6l10cHSbrlgmxbOP9kczG0ACuM+8CxhuKeP8fbIFelZPYojM9bKH
wz2MngE6AUHN8sZq1SkhB6sl8n9xcUgZ93K3UFQKbz87WcTY8d59U1Exa248vJpG
Gge8QiuxwIEIZTFIxKt3RSwr3+7N33aYNReqc4B2LR2IIxmJT8ZF/6V44MPi9nxK
yI5f+hjSP+pXOLZIrSsfd94s0lqxKkGsIT9P3eQE8i/CotF2EC37M/XmFaJoNw2S
JiGk0pKYjsRr3eztYBNlYHrvw7GxzW2jk7zMN1oIlGFwZbstE6Sh0LmoPL8Au0T5
wM3KU3cGteYE2GiVIT8iWKq42z5Dsq3GPkDDNRJZYjbX1EUw92dyJI48JeWQ4bNh
xqfYoT0enLz7YMJ/MNQseCUJEHM+KEtppdCxvESlrLm9UuXFhTI15HysVJuCn9k9
nSDdfZfV0k0xucEEXuWpreq7KPQg6uFIz6IFS2uEY4pGwwjH8ZXqjhY7B0IyhacQ
ZPbBvLkcApFvEtBLTYhVKb9fqBKo+BA4EuQO8j7EjPWW/EgQp5j40bkyCvPAq9LB
r/+2hnfcfmHfDaFLlj4jdIp/kXmx/mCzTSisebdEdTcqt5s4NHKTk++izP1A10mb
2auyfozjIWUxZKLv1KFp7i2icQ3atVu3CIUsZr2HPw84VVvQX8UxXtjwPj4P52T6
M/wNcFmEU35Y9i42KKNE9gv8TiBW7Et49M0HrfAxDpnTWx9Fpv0lKpxHlrihBXhM
VqGOXS62hterBdvOaid0uJXYgDsHN0rMQ5iRWcs7frLCudIABklTOqiKS3T3RhP0
nSAMXT4o9mD8hSwgiaQMvFk58FTyIkHBEb8FFqnHLPsDat++8FHZEnXrWNrXp/Nn
sn+4ERGwXbmAHXjixFm6xDWdh1HsKbUb6imqwc/2AN3VxrMikYLozMtHhABDlSWz
YehXsfhfj6UuMNTiRfYVlg2zI/lDxIB3zxTj+VBFbTncFvg/uuS2N7pSlICrdC93
47s0AedIYAmX7Tm9W2KnnDyViR+wwIjGW73TgdBGkRTk0FxwHYoO1bZ5vmcGHxiG
59OO+y4gVIS//iZBU4jWqYLRP0/ZAuNC/0ndG6LF1SaJVNRaBrng12fWQP0EkDc3
1BmuwJgH77SNDbzu4VM6257DDNwBGnI2BDSlha9eMmKeDj0uXgi2TGXyjVP2JjFJ
gO3BSTSVYWOKvY16FlicEf5RNu/4I9f1bg45RbeyICj9fltzOBDavs3HEHBo3pv7
xa47OFiy+RsqBOKXdpyvkQDINw1DR2sHqTrK4m6pjOg0ch+NByVeqG6Kp+EQ1kmv
ikXv8AxzQ4TxQIG1kwS3cAz/zDfnDm5UUcvEuMchUa+kis2v7g94Unn0MPO8cyfv
uWgfsX3y4/8nMIH2PyduxPwzqCdB8ULqzOgwFqZStXoeeUZ+RyaMY/MhAwOout/V
mEvTIqENvWddg7/x1pkSkCBNHxH8XTXbKR0WavMtRr9X79GgMoPVGeNWJNmLgggE
W8b7/8JgcVL0f59k0QQDqkDbv8hT3Cxoy5JGTUhXnXNKFICRfv2fq4oTFCjXShU2
AzGqDk5kV0+R+hQs2v6519jlN/nWJlEy8YMzxOh5QrDuo0QVAqGcxNYsP2hq1jE+
3sYyEvNFXefefn+ETGkfz6cPaA4PwZMB1oUDOW+g8N444JQqCnztHLPakYsHwUtP
PTE7WIA032MCjjOANoFAydK8gLOuIt/Xtvjvp6MqBpwV/DEp4d9suLfk2WXUSA7h
zZ3FTm0ps+ido1O1ZpjZcBc/z4U3bpKBD+bWNnJ+cfeI9EAQE9WZh9cWEAiFL1L0
SVvHnx2rvSMZnjImn8osJA0fo4zxoDS8dBTxzK9J2sH+bCJnUmL6dBh0WpHKoi/D
QTMCsUoqv1QyQFSJA2fZBtd4hq464r/5UgLgpIgEFB5OEoVGiv/TIjHdJ8mdQjry
uO4kYIPMyADN36SZGOiy+JJCfB7iwUULsIFcUmMcnIxnqrLTRJ1m+1NIVmYs6Lap
Pv500wQfNBMT2oeZj+BrviylRpOBusUcQKUM9Fc8oh+sPebrM8E2EmUN1JhIRzsz
Zv4fJvFvwCpphWygCDg1p+fIhPuUYUQji4Y6XsENqE3Br1e7vk+n1d22jx37Qng0
d8ye/MQzFiacqjzCR0aEtei/e8u4LAsI/mYamwt1nLxMQQjQsqjryHl+8CzP4M0/
VZYUn/dX2Gl56LxGrGtCuUQusmTCxRisR+X8YiteAXFhfm7IqFDpAmUtlel5ahMT
mJtHMaZMjwZB8mcnLw8KDBuPOe9o7ogm10HIqAoow6K8dMMghfLFY9Gu9v93/8p5
8/9Vun1MIb3m730eFd15/0gp3lZhcTTU8gHjSy5+4mNnGoS+9domxHc8vZxJaS2A
I2kDD4VwLBxZM4QxR18iNWWXRkAVRWHMu6tXG5GiBfBeyTQ6Xlt8uUev09XZHzbc
VVwywt1cf/AtijNplmf1fikpT6WsOJqM/h8FLqJBdQsbY1pgN6prevEFUwfKAteo
qMCztHx3lw31ELwoCFnFluWJOGmBnFkh/T/bXnGnBFzrr1M8YJCTtKWxnrVrPVmh
ksLcO8I2rXPMnLI2ou8xIXxT21qq95DHMGdbWdf0g4InjLjcO9wVOelHv9Le+gJD
gfzUc66/w7/KMc97a4rKtxw81k0aIsBTOMOuCy1NeM/hkrkvGchT3iQ/QCHTq7+P
Qvfddoc2/hp1HIjUJr4tKj7NxOi+Ff8aAAJ6VZhQ68EJ/fM9+zXyUYSasYXTVpOM
rFM6793vEJ1wHVSzoIpQ8He4fDdtrgWJ0r1QGLZ9IC2Jtr8OdKhYlHioack+0X8W
t56Occmv5gUJGJQFNnj8tg7/NrJ2rHJULfCI7ndz4GZsxK5RQEW1wiIpztn9oPFu
JGwpHVs2fBIXl3BTSOLwArjDNf419lBt8FJLcJqWN78NqL5cVveIH/fPpNlx/Owe
BgR5F0AOcpF84O/VHh1/0NNcT6nyaOARTjXEM6WM7RA2RLzhDJzkd6DiKEbEDai8
XAItNnT/6Dt6j4lhlOWbWv1NFVePoHdmxUwouDJiE0cUJOXFweCTck0wRbxBfCsW
TXxAyyvno327HdUv8uXkuzYzJouYl3YkJDDRVdBZjSm/vGhmELLwkQupKiTKJgtF
Oprpv3poCQ3rKbf2Kkk+Kf7eGmmTRotVou0eIiSCgFLgxYEcSXmezmeskIu6lgm2
PelmeeisXTar1UlX4RtXuRKVvO/sMyzqFiDbY2Rp6YhtuH315eJMvdyHMglX9Kyi
V00ztgb14vRVHUjTOF26UoHzScsSUJdEriBiYbSSifsuelxVtk+jjK2vuow45RfO
3619CfR9j4ds4s6rgkw7ulz1pk+isvsQM0ZEL3yfs+FHZXQx0Rr8F5oiEFqNOtmd
VN9ipLc05C+i1CrZvVMPxI8ETEuQIrHVbqsjTY27+T7XR5xCqdXM1i4cIX9OP6Gg
2WaK9Cf0g4NzyB0xuHs5ru97JX+XnixDbL77IFl9ijTwOodl+OxmC1W//5ZyHZEO
lBDJ+pLD5X6dhWQx2zpv1doqsoB31mOYiBq0gKaHaujnRcKZS7VNCikbFnLrmhDH
LNziwJ6mbTPXaPX0sDkFp9nmKGbMsM7wxbTNuARBXV/ftJKdI3CoRqXI3NAHloYi
DczbDpcazc3VpoI8mSOEH6mRojGp9rX33BRT2TJxpzY3g3LdEXHRs429o2NTnwnd
uiyGPmeyJ+lYFy/dMZq6zEcbNlyd2QFLrEaRAP8j22Bk0iiA3eOIcmqqGhxZ+mSO
nOU5ratt/xD57wadpdW1MVi48tZpPnOlNW7mn6gFytQZaJq3p4HZGgYTRxjVXkRD
Fl00G+Y2oGk8KsP5/PIcq9wV6De5Az28KF/vutrNHundOC3rFVaozGJGLCNjT/RW
BUZoJcNH4ahH9KWZMNBTaU7MMLePIfP1Tk8OvM6ej257qmJbZl+aX1onBesxS2rB
9ypENEBVVbVvZQq5Z39ZwfjpnsHd4vOyKwLU2amcJkOCXapMdmMZPZNsPj8c8ueH
HnROa+qWv+5GZhgCCfu28vcsd4ix0T34nnOrzUUCHW1zvN/qIVHxrCGrG5KyhOlC
OoQ63/KdH3VgErOzQfPVUX2j0/j46ZgFNwiPO/sv3vceYI2o073qH1w8/5Bw0ewT
g3vpiDm/AORaP+HaASvPQzw42iZJPLJmKdLrE3MEu1LhxHovz+e0K06e/h1pcrMV
8qb68S7yxmOkanSWwTK/wJSPMjloZAq4JYHCL4g/EV7CGoG5uWrhAWWnXOCAulsY
NgCv5dp/wXEoP3wwM/vo0XUI640ruCwwsk5CW4qwb0nDBZiNRKH+moL/ngDA+u9v
9tFf2sn8teDoqZg1YwgDOIoi1+nLu0/EQvOFZ3zZXQc/y9Wj7ZmBDfvtKx8Y1Aj9
uPCLbI3SwbsATFn7npVR/Scs/1hu7woXEMyu/SzK5yJltom+TbPt8fjDxTT54RPr
9d+QcX2eSpIz4wV89p7CN3IiciYhMz9v+Jma308VmkmnIq0p+rxZrheUdibx9i5F
XUv0ZRlYf7ArdQgPVQuCxkIuiqPlh5j4eYhs9JjIS6nZle1Fn8c6QFwSL+L0ePVU
nzfola/TbGt8tOdwZWT8Cei2B5TsoxCeR7KMZid3aSQ8Ak1JxqBcz7GWTONuLxWx
xdWlucPszT98XDCB2ufocyYClt054CreM3kYlroF8yAYQOGzue7hveTO+73A0+By
qhhi3kEeuTdgCe9Ak/SMWxlRkb7Igs02KXTLWC/7UN1Z7564nImcEmXaa1pZjRwO
6QOBRjMpoLjB8wMYOqAHQnw9hbrK4iAA3D3e7UwouFYgDQPxyQQTxmskQ9WmUQPz
jyDCO4e0xwhSLJ4XH/Q7x/ZczbmSkzDCJ/5kd+me+OHof3qtJUXBH9tESONk3g5N
Tg9xgDyEqVfIOTv/g2c2kPgQYHjG2RhNSQP+enjYyVTEk7Us7rHOvpOzpOGzWB0Q
7gaUkYHprCoI34SXnNz/3ew5kCdKiMW10nV6/h5O4JoVf0fvoYubC4uYbljE0Fzc
7v45MmFL2anFlLqYRu/DNsgSjt6tjaxxKECpyRmRbUG3iAQ9kwY3zOSJmj4efmA8
o3+yItAyOXUVgkV2wkcQFsD57RJYZWmojamltgHptKQtetC8NRya0Si1MYcQHfr6
vK6Eob9QDZXaGgsJAO+InwTfFwsi5nrLzgcNImMnJTj3j9Ou66N/BLPxqw6ps3U3
FnZsXWaoehAd04yci2WQHArVkd1Pa5TqveUOhqMBLbFj0LkGRBsj0WZt3I5FHVY8
ME7PPbxi+hs8QrzFfCwOYPzz8WeTpOQZDRX+v2E971CqxD1dwrXvDtoQMrBFCh5g
c2EvsmC++hgQ1XvBzqTpbNR1uC11WtXfOz9v2EXi0ZqaVzByvA+og9/LHVvFGZ1y
2nUqrak5dAAJzWOKl9cnwopWH5LG3lExPPAFfDvbEuTk+06L6odbndxtZySwovQo
rMzB0ST43xbinv+d5hj9QT0YK/5MnYbQZchXKweyvAYLf6BOIPicCK4dVZn1aTTu
CWtSdBuTyJvrUIzcgqZNmUGCZi6pmSa8GE4L+u5OA4gTXp1XsW8SgPD/po0gy95E
j8tAS3PdGhqJZiM/OlDuXd9v1pnKmZ0OwH9ecDKmhLOB6+3itpPJFTXnxQiw1uGB
Q6URNyaswhwDzlg/YCMdhz+Yx2bC2cAmlqEKVBuHDzMQFnXMnyeRyrDlcV28Fjd8
H+Sw29Y/A9iBNxE/oE9kVNsvO/fO7iEWbVuVhAEeboJvgBZl36tFpr/085rYT5YX
1jrKo8b7oQq1DJyFlyiOdPUAt1O1i2UWlYnZfqX0gsrHqFuz4neLHjH1zBMQZpM4
8gerHIuxKykhCQa9rh/Sii69zQ0nrFWJOo1MUgxdv973ymZ9Qsd/+VKmE5uw//Q+
et/q9rN60dOfg4A+aRbarNeSVehr+YG0k7FWXkvjFEilj0oiGLPf8R2mF4fMJZVN
7vVuulIHEHyaPLoYxsqFeSNtRvf9CUTZhmiy1d1xMmxZNcOOc33fFY+s0BgtmXyP
LkpRFkmYUhTLnUklUSMbvrCZUljHat62ImFMjWXgQ2riUg1yCBtEBoqgXx7JJ4MU
+KuF8UPKzlQKv3shCN1+hKCQrmgGsmurlNOTXWjqQ8J91c04ca+k9bu2tNkyqwCX
ekn8Z3KrOvSsv6vLe3qpaNLATRqY8sNIGGv9IgaczaY4W2JEwI72twj8Vf+3cJcs
SmDMuFI2k05bq1CA+VZ0PsnKJRqO1OgguSKJza01kSBedP987WKiQdcgosyXXWC/
Q/QcjL6h6TNzjECLcRqZDyQmItNJjlAliapbUCzIoIGHitF7dGbtxbU/j238xvsI
X+u7qwiZlKZkx6K/iP/v1EqIzVSq0EhJLnH9mM4Q/cb41apyZDyf0r3siMp8V9Y+
cx35pjoKRut0VwBVhZ0xeplI+8ziaOZe6qFkE3Ggdh7fdd4snZcrtU4mPnbHwe5+
sgXBnGb09xg0shsQAuGrF+rTuRXjTacxggSJaWjoFDN+Qj9b9Ed+KVp1QPq9nmtN
k0mKOc2yj3AtYx6J+CZJ5KmOj5MZ8QhwynUoLpw3Q814qfmBE53ckSVYX/Bgx27t
tyKquaMStgpdzhHCgaK3GZo1rwR+PFWWG/9m8tVfw2J5YP0g/jx9uEEQMttaUt0K
ffed+EfQveugYUxcyTAgAdwHI2UkarIb4nCsqpa1CU7irJVV8H7F/23A9FXa8vp+
83de9aBzSrqeig1SLSsfedgkhvNOWcfI9M1bls8Bm/XtIROZJ4KTwTYDxgt6V97X
Ffo5aFW9Ocig2GRi5hqYQ1bEk15BWa3vFJVZLCUc6xEn+vLFBb7wcD+yOMeem67n
/fXDdWCoJgDDRsa0OzHI1rqIzJUfBH6t1rb2YoU27qQYv3bbEWnqo0jcBe+3sG4o
pBnYg4kOI2Qvr0Zdh4AVUrtECfpWjqDntO477SLNuPEqznCDLvvNegB62oDQsZ4i
7yfnJKQ4+Zs1YaAjP3zBJrnf+EG0/DPXTshqBP5gHCtMkGkdocoQs2WOS7Dnlr9P
6pC+vQvg4diBCQo5+CY6L/eQHgRL092bUjrmxKJwSElzTRuINTUv9iCjDZy03pMx
2vnrU0RqGGXv9stfI2E0g8o5feHN1Iwr7rX9N+1lWdZ2SgWmO2QnlWDCXI76UCc3
Pk/vK+yUvAfF8zcd8MdGDnoQQNLy4V5WcstF7etUcxxFNwwd6cet3yXKY7BBTGS8
qgy+/Fz3Jiwr2SBm8yJuPWhpL5dD/tUwwbbTx+LfSFwgZhIIp5WffO+nlWGvh8lY
ymu1tF3gSGgVkCXQ1TW1MEK+XaSzi3QBSlogTfKTLoVl/r3/lNzlrPkJ6MkakBbP
/1Xv7d/D+b5Z7LlN/gWpqBzeMt7oC9CDWrcfpPXZoLNWaQBnlTzIW26vS9MrKXZ9
6VRVkZoASINwIbsxXDqWfjgpT5hL44/VQt7ku4+IeMeOO5KwDkcH4/Igta/QGPNN
WUbUVGSqCZMs9PmBxApG2mW5Oa/bYm0rguFCfv9Y0YBfenySAZREP1oTn1auntwl
9IPLevwBgjPVu4qBz7ySOos6egCUqQzZ8TkOf5cMEzCKhZLCZTimJh9CHD1vL3KI
Oep3M6OI/fNBjCOh0gI0edhalGJUVXY4oc+35JTeChnmPj9tjPnhW/7NxnkvFVT2
eqkdxcsmnATWjKRkBKc6GAPv4ZhvLc+c9OSFYKzqyihYj+2kGwGlmZ54HGQOiWcK
vYDTTfya0ZHarXagnP0ytokWLo7fGZkuTsu3KfaOidYFwt7gkR3uR+qXGEh1JQq4
gRuFUmms8fDGwVTm0y67gbLPaaR1tfjFC5OI2HMNVrX8HTJ40ONNZ+VVp1Td+z+X
UGu/tOeqapEM7Rq3XV0HR4BbiL8H4JO/4Zouk65AwM758eiC0NMcAAIDNkJwwDly
kOsD+s3tRycOwIIAOBHdVHIUgmI4Y+DUDQjmAj/VVM3jVdcds+vfDjpavTs9RAQH
IcF7UA0u/r8sAWS62dqiNrcE+6eyYshGcHInK8fPGmfbQMN1YUD/B395a27gJhlg
7TaeP4GjqDQZX1ZCmcHuTXvrjoq6eM0jupwsNq1wBRw6xjCqaZRlu89oWmfe/+g0
qctk90QvpMiyKGReCIDPrjcBPe0h/XeliXneTBt1pXpBlof8O1xtq/oMFMlY/jtJ
1GnTJ1fjsoeM354b5hplOL48GhoszrulHtYynORJmZ3hfIaCFjRw63LDygT4TK8B
DfhsClJOXfpE7qCAsrQe9ZMhLeWNSWh8phvRdHXi49X3oP+Ja86Vl07p/8BNyVAp
nfZIGIRgl5+btdJKGVAjumWQdBM8qV+EqUex+/BME4cAQxbQt2VQKqVtYR39sv7R
11gt6KUKJLO7bawemgHu0+lP33z8OaLHJMYAb64t34CTKwjMieFzdcTk+AijmnPP
7bIBf4+lJq9xx0YWJgYeoa3BYAbpSf/wjskSeJpHSjKvSQyB5bruzm5qh6XVSYMi
kenaSfaHumdAIwMo0S2InOB4XBFCGUxZ0dwadP7CflEJOMTXD8slCL6U+D7QKseS
E8eBmNjbmRpQiDPuZ/OYA3HLFw8+zOO7lAgdgFq3MAGfom68M9h46RmSotRkf6EX
ygGC0IP1GtFafMWpE4eOMJNabmT4s+Rp4NC1FM6HgGA9LRpnzIow2m72Che2R5Nn
z71G3yjHpw9Zf/RnI9nK6KN++6hydZxYamvymf4nnrdb7bkbCwUEjruV8AN8nBiY
EMvHvATXfLFMf8oQ12GM+b/WV0ylbso06VLHPLWJ6Zu4fRIgP+k5zb6RVmk70VPA
ZGXhbnh2fiIoW7wrU3WYP/ONXM2ncUx0xDb1W7MWGb0mHCD2/5xYwzm48dW0MjW9
wkErOE0AYQrpP3tjpgz2kWOl24qyBxR9o44Oa/lmW4filLl3B2FA53Ooq7vJHlJX
sztn90+zTwGqIy4AV8SIhXEkjaDcApJ7ykiAIqfc6gmjsIuMYiyz0RMA68b8oIcC
PzYoUvoBCsTcutTfMjWuAqhQE7L+u5jwZ2W9yNprELDU7MRGRtECHrg0d5Yt/OXX
2V1GauhLSaM1NLvwl9S5RwVu+eGqm8zON69SSiJ5O8CuI3GhFkREvZbIrHgOZkXh
i/zD3tjPG2NMeyzT8xw4xzxjkLXNFLujihTZ7wleF6QPqxeRZaqbjzWhQMIbmvZ+
juio2H/Q1Vr2/vj5ptMhwoL76KjpW7Kv5HI31LkKTaw8W9NxobkgXh/m0gkoUPv/
dhmayLF1Xv2/qbse0aU3m6osWbhg7Brh65B4HGr9+WXWyzqg7Fz/GGFdrzsCIvJt
0cFEKSiYj4189LDE7QgDFZ8swE5DVLCEsVASgQT8gRSAgjxZdBjIhNv30zpma9Mm
SHtTobwBLy+PwN2fqo8KMeS63u4ZdssPqe0T7ZdGmFC2Hnu+JrH8M+/LtZ6695cm
EwkfLIALpzEG+TgLly6sZ8rzmxmLbpn6l9x5/v5LPc23tFge+VsTP2DyG8pApwcK
j9dsRFGydveO0vtRPFUhtneos7R6H6W5sMRu022IyDJ1RqtJmOoAzAS7G1LbRXTe
H1Prhw1L1EWEIPODoyieccbeshtQ91nFdO439eRNbPJZmbJviCI4EIj1vA7ncVe0
Ys3WahU89Ap8KKo6YGkxxwrc+/14dt7ZAgTFsOZ3cSilX8zLMsgFmV9euSDTSFMU
Cra0nzf3i7GaItqS1sZiQQ9Uq2ySfRBrBgkXaUMKDk1K3LBhddH/aJP1KksqhRBm
X9WFgESYhlOW0dJmjdSJi+bICnaUTKyW9mr+0RadlILxx8SWgbjuOqtZ1Yji7pxG
/hDz9hCxK0Cs2S0vEjlmpShcP2UsOUnDSrMA+I/89CGKjjl0IQkTpToO8Umoy4fN
XwrVsQurWrXSOibDS4rKwxenlC3/BOilurreR3trnmFAAuZZqS8iqVAxj+0WDuDp
7BDMHgwbVoC3T4VxiLRRLsb+ll1VSw3w+5YPLPe//hf3x6QEjlsDoMzCjz4+/C4J
gaGW57EVf2E29iAeZTggw2l6C2yyHFzLpzZk+MC9y+7A6vd1jbsjSlSHIOG49GSf
yiqlkA2Z0dATXNe126l/ijQfEKvvy6ImmGZhZ2RJYzKo4jr5mJ+XI97yt8H5h7zl
fuMpF6e8hGd1atXtWAfTvMTclRxu2GazYPP528FBUA0FS3eSmVkXmADTup38Dje3
m3NqDHb39Iq8u0HQL9laJ8RJAawFJ+0R0YtXxKa8tu5LAdnY6F9Rj0+rQPD63UHY
iQv9fhK6/kM+etr2N4ryBkObjxRKQ+oBEJuHQNdgZMMCQre7SnDgCIApJPviEF3Q
/+7YBZgv6BzG6iCZwWHIooqdWH+IsiksuvJfV/gNA2/lRhp+uzbkVMeR1oFX8sqf
N8oAdahtoDdm+L+GZ2oBDFILE1ltS7Ac8Lz2UYBUot0tE7vvmSIvktGYwxYUS4k9
SAr+wamYSpg6I4x0L0rmCwjUNbyNVPixxUioDg4vUo8RNq51WcpdwEYP0wK2nomb
iyxFaI+0k0K0dgy7gqMygGOBcUCdZ0JFk9I1TW56HH3bS4o+TsXlHVlKfavyM7GV
zBdRxJ5+FYd6+EFDOy9ZfWwhRKfj/vithdn4RJSEp9o1qVT9zyG3IHj44syxUVy9
2ZwIlFif15qxV9oNFDp0j4R9R4SsnY992RiEaL9L001mTE2WaMCrgXBrhP8I4MU0
oIL6P+p57eRYoaPC7k7Ru2a9uBCeeFteBpnLloxNeqjsdWzj+7mNwmI64+VAdIc8
YaUKaVWncjbKZA/R/M0ZHin9u1pV4GVIMb0T5EJlRSTDyfJAr233bESVPcNKBaCo
CxrfT23vnK1IaJGygdWOXKzS1EW0eS/LmgJwymWvXiyGzL9dgYooOErU4oXUny74
uw5BbMIInUZo/zZeRDkHTB3NifUkrsbN9gnRQ4d0xgqPgeT11Q4QZZgMteX7/4D0
s4zoDbnt+L50G6xCr8l2bz1ZESxJerq7cMUqI11jC84raChOhuTG/mVJBv9GTtX6
dDFQ8G9f6dAAl3ThwsD9nDenrcXYXWcYzD1wFw1bxw+GJVvRmVQee4MUmaJ5Lid+
tWhO8QmS+QMSDYrwrUeq2TcZEizvB0fGXxyYTLeOtMXjb22Eksa+y3nVDDSw39Eb
w302hr4z26qB5dTxYVznme0k5KYKbV6IZDyni7IKScTUe125Aatf9XsJQLssc6ZC
XXS7rh7C7Y4pxfh6TFCdDwSBLPo68oVgc5VqkvqgRORCiarZTbuep5ZsJ6hG3KN6
xEsyEdxxnXMXs1rU2obfTNUD0L/lAZzwWeZN2IxezbPD05eyDLb5SLQmMnCBZrpT
khHEy+D8sF46ECW9UFXBj/ECQ7uqqktPWtNaewT3Zi/BbjSqUgqnZhmC8Nd9Ic/N
zsR6dyCJpCFTX+WGj+d9OYz+H19XPM8kv5PiZiDNmDiQpDziGAMXOI4BqeGTYxQG
4fbKQ5cBA/dV5x0GZ1qxXRhrV8wFr4jPCBrUDWYfUhVjsT/AMmTyw31+58iSXyle
+MYOtK9+lS+1GqNGWe90tMwb0hIqEhroSFdvmg0VVuqqWb7Ub7fv3+DLpXTEWcWm
akTzpLRi4/5zBLhiH0Bms9fZrspEvS86HPlakb0m3U6MyfBe+v8FtvSvURZ11ZGP
IIcUeYPA9y3WCL0TcwM3NZQaamQNW0JPCnEvNTcR4rO26QyryQwOHDaB4tAILCJo
M8Xmh/qG6FhXymTUUPKA2Wi0sIf+9k+8Yicmbhg1mIcWTVMokd2WTu9w6Lyq8Nhn
Ey/pBlwuRJ/XfQpnfSVOENBI5LHCbQXf9Jj5Q8aGy6rBavMxpu3DfUEH3usv0Ety
ZpLkFH7464WK4yzTR7VmdpuOZvgYgTMcqAN4nCHbe2G35mWvW/DjwAeveX5REov4
pWU96NUqeMZy54FdKRo2fBCStVwWz/8PA8BOfsJkpNhKjrqGLGAHaq/ly8u4VxFo
TL/Fe6PuS2FCQExvEiramWbgwoYtetv2FK2uDWMMUNavHwynI21x+iG0mA16HHKV
hdXieI2JseJnFn0QMaPS6IFbO+lZqIV+gvHv7fe2FXcROU2pRiY8OWDLkvBeo0+u
bxTPFwatET5kKMgUOv0gYKmSnr+K8btSi3452abXQR2eHPg0LRyjLbhlGqc10YYH
uhZv2UTtJ0ivN/xKoBukcBfkLHiHfIjxUp65OUMBlTaBrVkDoAjhCbt6U7h3yTwo
3iTuEId8ySA9b7Z6dz+6Q9XshF3C23xf9XJL6zCi8eQZPEPmXJ+BiCo5gQdoOh7c
P0HGhlS/Kg4Dn6xyxUXQwsmsyWq7VhZD1MU58a0f19NKZQ2RyUYdFHMxk/A5qkz9
UXR1F+k66nPcbSM/LmzQ4LTOHw7A2qYCNm5P8I+PoH8L8zxhwA+8YC3Gu0RM9mDp
aaJ5D2/it6Yc+kacH5jt2aGKLVLyvWkuln6hTmQCbHaNQgWYPVjv5iIzoqXXINcB
XXN/J7VPElb4KMr7Zh4PoU7eXtbFIWUg3aqEHgsL6ThrxOGPnDPPRJEsLxSH5dId
Datai4yF8i8UK49hPhotKrRjFr0S5E4u7IkpBHGI3i2HNyRAmiOjaqwBD6tFFmML
j5ZRnypINdd8yOBd4rVFEuTWj5HqoGmE7HeF+keVe6F2IZTKcurIYrvPpuMlTQUg
Z+7y19wtko+0RjqnjeLo7inOPsFbaEBcGUEYuUsvD0O1ZRaB52hguMDIOQ3hhftD
GffcYtBfqzid1AVLvMEAjOuDGeWYL2GohjQwfb+HanrGSl6TZuJ8Fl/+XxBmPeGH
G1Rg80SM8M4jU0XbNYasGujfKBEOMsmDrBxz63jSPagSo33bs1pqYnQOpmqg3Isc
aDfaY16ux0KeHIsLTM+/BpSOEJYDTCuclBHVmSmp0GxMwQ0U78Hv9yAuF2ExTuVY
mO3btiBzagye3DqT2kxwbU4Plr9weDxneVgi0imlK/gAooPbnQaXW4OAB9vHiXEO
P6lG1hOQ2kGZ/b+K6f8Njn0dbQK/9JhMsAs1hMPF9CD6jahqqxlayWk6vZ6ZL4uc
tyDNMdOjH3HRu7vLAQyiRs/eTv/JTx6utbmXc3ryke8aqLit/xHIL2B6+6iHthR5
4r1z/1Rcu8Pm9vI877r9hl7FJ+Q9Aapn9T+Qakx0Kqo/kEKTM3tcEoHlTY5NfMvl
5eeKGjybkbIE7EIKtdME1++TVMYqJZnHF3M6DdyhtI9jaYneNgr2lgbOuCh1tzvI
korQJayvlWLAahuO0rouJySGMimFXO9Te2OqPphQPvi3ZYBwwL7uNnK6mIty2Hd+
QP73E9a1GqMF1miVhMDBRpnJX1jIrJZCwthKi5bUNs0SePw6281tvvWhLf30F03l
dCLoYsN15wXSL6KKEqd/WUEAijOmxFUanb8PV3Kc4sz067pYSZSZ/w2pRsUM9/Fn
Vet/usghgcR2S0kqAfmMQtQFZ27AI8gVeOFS1X+py/UNUBWAsqpo7cq1lyt5i2H2
6v92uhr/MkxqhTmy4aJuGT9RqEdda4bDQ2ux4DWT8haTKDcf2NoIrBJ/cbq7E6g3
obR5tXKsfdPSdoFoxc0uexfi4Hy4hVvsa/xpnNR9UVSqd2O7C3i6ptMvevImng1C
W9LQctQaZZvU/3v4NrLSCo5PQFFxc4NfYtA9dd8cPpifck2ikLamJSO+C8guucls
V/C4jTzUtD7gHp40C+c+cCIVRi3t6byGidKOBVQ9niHhO+UR0w28y6Cr6mBZtEho
VATifobaoXgmTE/Wkd/dyJM/4tpoc6AXY/XOATTYZvZRD5RP+V4CDT8QZcvTextq
cEHSJZJiLF1qCCow/Mq7h1YkCCJRrASRyhdn+GZZHlh9eQQSYpd5Lvgm+jw6MB2Y
qlwsLTkqxCCETtKn2zcp344040eXdXu4eKlg0z7jf/PCx0fQKUwRHkLEn9tN7/p7
OT2cEeBbEJxVMYrRmaULAnw81YN2j1qwsJke8KMOVf9G9uJwrZVFeY3fIrZcae3O
7R6Asq31ogKgC+DlkrjCXF1BzrOs6qwauaBOOqVOdRoaKz/lImxm22eqHxwQQBJ6
H00tdf9N4bvHpptBDNpTR3dKR6bdFtagLt7nrd/AKdVn5kbOOfx8J3tpCsF5OU2A
WSi3EWqxFCWStime3VzA4Eb+egKp8y++SCEP9JsAwPtFPm0xFRjXZrTw0GgLlgR6
hH3pjq9CtgGv1mQCeOlYp6nYsg+QYJn+lfG1gWWYTriOpI46eG6vWVHdiWdaanmS
+vLU2XcCOihaFLxQWK0NIoJvOP5soLHICsRnaTWkyH+v78qBK797tAXOBiTWUcHx
A4mMU0kGmzMNe9fh+RXR3PBKI+BU80WVlbLOwg5yDy1MLZVUjpM8gQm0CqjKfiQo
0lLufUwm8qfopo/tvv/ysaszwaevy3tE8oglBqz3wFSJglCGd+kzIzF8FKrGRVgy
C74YTqUTyGjrds5FVdDS5FoY21qa+BqhCcI6mWpGKooCeUsMbTWmJKNGL7JlUV9d
j3c7Oej4GeS9LzuYwacAW86xdr8q8/3qHCrVZoDhBKaV8ufG3g2SQjk+4WaMxenz
2ACQt+ZAI+YTcPX1OPgjkXIU95pwnu5sINmNU1IQRt2+TitlZhinJdroImvbXi5G
EP2gkc2V3NwioCNbKU2+cNtgvWEgZR4MGRfYmItln8+DE4XOX2w37ASevljtGC5b
xTezvXYtvciXQN92ILPKCcdqbkgHeE0hAPMSYHIKhkUMV8qNoEC0fhHUNibOC01T
b8Iear8xKViGYMGO1lD/holI/v4k84Qv/cDjuRp0egAfmCAQToWpVEwNs6yZ7Emt
Mp/PxJw/zJmJi8ffZos/VouGJSx3NnGvlD9ehIZC8S1LFmYI7IE+goY0duFdCWPH
csLm00b2epDebBKN7G4uIIjV7jcWI/VrzQKTkHXaLvqOWb40Xsje+vXCQTXReUi5
yDB/jM/C4yaqFNM6fKut2dJf9onzl28ShiwGdfTn0zjYyCkvfKkVViMeB5U7yF9r
MTNtx1n75rNjCXITJX//k3cTYm8Sbd8SWZUW0RmGu23DeBx0qHqcs4jmNzBb+PPF
Qh0BUOdk0SJN6bErxms2k+F1whxwuj/auQLnRP5YmRliGrQiyKfQm5XS/R0fH4mF
7+Lg+crrYLhNO05ucEYTs1HGagmIBC9aNlmWNsUWTslskRdBR0F9OATyHxqeb2Nb
mxBeUJEd8tBVpbHNUVvb+pm5VmG+ZGPvoyoE0R5wU1h0qnb/x6uOVHfqBdXjUozR
mkZYooYh7WIOEc/cAFj6QViTYjPGE214Vfgsh7HBsXbvt9fDOW25nbB6sDEzF2m0
06BvtIdkai0NImSsA09RiW1DSnAGkt2feIA+QeO29hajiNGf6MCxpVb/RoPptBRS
akULAYG89mJv0OzCYQsCoywcE5P9oG5BkY7U89UJsELOpyBXgnFnJLD9MyV0FgeU
QXgLS3jCbBb+tTv9/WBVkJP3lnBtF5f9o5yLkxJsuFIoWfAdmC2RA3gvTKKcX20o
WV7IYhL9Y042GYIFu0nbf9VbBdb6D+qe2Vjw8QT5k3MwLmqb/KrhPedGawtPI4iU
8Mw06akSu/DEeaoN08AM+XEc3es/08Ga5KubEel3HjDJuA7Ji9m1WJlRtOBnVwTg
YwPoG9sR9TR6mh6lrsX+nY5K422egqU7e64OlH7dIAmejF/PAmu06LwIDeV84D1R
8ATcS3ehNzOCAcsKksnwwe6ZTf0KU0I1gds9fY6LbUinvepGXcTf6BSwcYaW+gyP
GEb4B7MMEI20CQJQlLpekpPG2m3R5CVUhj9gbxJsAym3VQZ8HiJpH4URHwjSA3g5
9XzdwtSbk1g5U1TG99rf1oNwb9/Pe4sL6EIdryk63XvQbJLTsaubdO1kpyFrI7qx
JA0XqVpzdStbDTtLEpSRu3yZXcDDxr/j13MCvyYJlVZMrqXosoJUI7YpTEW06pSi
DZBKYNHJnrroB5ZIHiJkYFF7UK1AD1cZZB/iIKN1n/ZQkKKYHmP25O+4ig9NdjCQ
TNfvDVYtfHg2NNHGQtYktqHWHkxF7YqWMvgZNcZnwvfb5G88e1HWeNeQ640DpgRO
cLrBep94gCutNZxFukbs9SmwY96QhaZUP36Gdvb/5KB8OS5SFDGCwYSJ4oW2cJfX
Gie4S535kNH6hhhXHFLnW+yYDf1frCUzQJJW4za8RV6LbkRI8KDr5HeeNJgt15nk
Ppj1bcoDXyOO0XLZoeePobudn3sjTf4e+QV8CfCBFFCq8RJ3l1HO0Gup7+8vck+w
2diwM1XDQfuSlyL9uT9zZX5bK6EWSWfQ4UfmFIKdZGewsGEhaR3kMMksiNS9NW4i
R8BYbfTgbu7zSEKt8M9vHA0iGdvfWB1KGpUSaGH2upN+NNUHqaR/3NJpIZtTg9we
IriU3Gtv3BJcrhEvYZlOikw+GIu4kYF1raqgDItnJ17qQoNVAFS3+EooS8VDj+k6
GrcKiWPMTvH6/CvRZCy+DgNj1LeRwis6aycgONu0zrvPWGg/nKydAqXp2x2aJg0B
Z5qr4a7mxnBP/i4dU3LHyzvVu38LRBKxKIw7QwdeX7c+mkemARD0rVbE7D1dZJO4
HX0ejoktHGYA43qCoHaccFWxOpK9GB8pqb4J0j5g27Ofv1LLtjUip9ZjVSm33vL1
sq23V8qKQqVH/nJ4ISynXn6nxb+k0JfI6JDC+2fdOf8YmDIb6fEbDufSNYfhzUOw
tcnf7Ujdhee5OpNimTCDxBKDAcXY3OXmS95PTC6Xx3WfDc3ckJy6qNq+JZqKagd5
+Z/iznwhgV2NLg65sCcsSXSvj8Gl4bnPLLgixlMqu7i/xek3VzbMw649fMVcgPma
eLw0QyxHKUOrSlEAObAxwkv2/xHsCngmdozPOFKGCCzyJRrmjJGQUjQzyA5T6UFO
vytgcDOrvOIZQE+Mw51t6icSICVo6hAXpfzv71T32p9d6xftQ0LM3fd5LP85RRh6
8nyoIARSLwIaycTGilYPKcBvhtP098uOlocMVKOngeTXBxjEuRrsywvrcLjjBus0
E7WCdH8V6q4nivBRpVdcHW9ehM9J7iE18a+axqPZ68nj6fdL0Unk35QUDlxQTr4j
Zi6YY8vWOaTicvUUMQksorCsLvMXPeu9iMWozGKSH85XzZPIk8Yfx3hapw8E6FvZ
h0/yijKww5sqfVgksblSDnMdbrKTYqncb6B9UClgmxG3MyDNPCv7fZzGtbh855Ud
8SsQgAi688b/2xxKDELaB++RqceVVp7TX3JZl6px4X/0R+9XHL67oWXDMtKk7z32
tuPHoYh/Vs1NuzEMYfe+RmF/ex+kGIddoUzEvrv/x3IFYMQaf9t16iWp+SoUYsLL
7evnfDuQ0zAT4/OXKn4zZChLzZxX3+RevVsBt6D9ympmPo5GGrJS3kPycWyk838Q
iZYQMdQHvNr1bKurdHwDjt47nfSPvieSUnxXaz5NzI8cn/JKFHU/hPEo5LHna6ue
5zoJVopfF1CH/UT3+6d0z942e2ACwr5hJosXnBVw1wHCfjZ0qDnLD8tekVFNRH3d
Ry+UJKyEpTPP73G/yV6XQ0E7LwSMCXVrhLWFiStRxiKhYTzVJReGC4JNus3OVimH
Md0pNZdWf9CU6unJ7xCHXe7fotIKFm1u6GDWo+/qlonMph32I4UGZtbf6d7tLxFy
U0eV5TU7YQbYgDHXbXJ0ZFQ9OxvmktE8kurbadOgoi5hJEB6HUJuHwt/pb5ACmTt
OyIqpICdAak8AZGKLKJVXFG7CEXHp74dl5p+HsMdX5uV/zyya4hbpeCNQ7xcHcYj
Y1Mf/xOP5PLG6ZppAsNpGo7axZ3bKp0P+fEQMtFbXTKK8YsL/oQri9KBuI5nRJFR
Onf68VPXXw2CEesW7AvB8Nyyc39Vo70wzgD8UMBCP5IMbMuP3b74WxoV0r+eHBIt
2A75+f1EmMEZXg9zqKdobXGs0d/IqjWptAl5q81NPpGGyCk8J0cm/gjJMcjYfuzq
T70ZsLJXkicTorrTp4s4pu1Jnelc8xoq+VMu6+WxSNgb0188bqpyYMuhbpPVvI7j
FciYIMJoVOcnRVETbI4pSmJcfPaQXLv+o5FtBGR1CcrzWZCbV/AuG5X3cB3rwz9d
vItE+07/C0bXLSSMsQ05DA4mYgrIG8vjQcy6wgsh9PQTBAVpzCbXyH+daTbEYBMS
VkltygHg2p8YB4A6uPq9SHqgtemRx5UIVBGvEVNwUDE9BerQn049VREwwJWNFjv3
PIPbUqMSFjI1c+8DHfT+DaEwUMMzqi7nbs7IAC5BLsqyXvH2wV2WbDcXbMUYQshU
o2EvjqxjeYv6YIJqYkQUk9qq/quew8ByBjDl6ZrjLGJEUIXQKJIlIWKIFGfEJ8xP
WoN+vZVplxMGznSFSgwlJN3nd91RmKcwWjhCfCe8CIVwVMzeCvUkx5bN0y/ZfT5h
8ACLnkufe7GUJC2P+MVIhcPZWEN3LhNb0dfNh9uHAQPT4nwfz2ILk1HNmySpmgJs
Gt9Xs57IIhr1S0dULP8upz3KZ5mrppKXJuwynm0p7QEIcb9OrQM094d+K6KTwHjb
KgcZoFaQfzkApx+HyW+pPSj/EA9VGbvEi5c6c9w5w4IAtOS49huTPViOWykJijUX
fjVEgypCLnxUBoxVfpmT2A1/ciY54BayVe+XWylxG4rJDBFNnQqKV3n1dFr4IWI/
UKYDJoqGNzts5g1kRMRvCJUxKqy7s1SJEXzB3R4DlJ5rBVeFnMY3qyYkqC7+tPhe
0AXqMUvRGkHyIkPih0IBwmE5FvMRFz3yzGr11kbnnV5TIRo1C6U7Ke8EW1UNosrL
JMpMqyymmFFCrbsNUmt0vMKINwXMYqQ7aUvkQBCNv5LDfcplqVQqsgQzaY9uBnnI
9zQMvyCA2S754kzaCXdd11XxYZXlVfO/3uy6xHgfGKKXUhwhqBSWJ0LAmVksB0wW
RwH6C28F2JsU6F3FH35e8C36DgK5VqemoDPevkrL+pTbzBmT83ErMWcYea0QIEcM
tKL7bCAySjw17zhaoX7kxZVHu+VFgQ1nvWJg30d0I5YqdIMaXoDh61j8v41u5jY4
GTBzmhY2ARtPJ+9m8vpr2NASLTmFQYXfGt/p+LBXap85Hx6BrSpAl+RAqQeQQA3p
1p7RT37Np7zKEHqbG0P+ZOC6mqyZV677Oj95uc1EguNQMEKDqJ8Vlb7XSxE0LjPF
ZLN87pa1Hvelrn+EOYfUhlfMemvb5aAV0y4cB1aOJQWaBqqX1MgLOlKn/ajVKJjR
ntTydNen3PBoDnUCYRACgchzP85hZtWUx15WqBDVvEFhPzV5RxXymJIFWu4BlPkw
L8TWsxcp1sIV94JD0sn7SGCnDA0kKGMkdl+awzHukIe1BMtmPO9DHQGO2SJ+sXxm
3m2syhOV2N5yTYuvY20e6NA2IPDYIk4aw/EWmhJlnynwGiby/rOjdQI85v4Tfexj
gDda9vHM+qShiI26UHCEbR/N4rMeZiMsAW0DuRvS8dOKir9tV3ux3Vtx1Jban4K3
a6yshTygFQ1CCyhabFpMZvLSqiLA0EYM1GiwVZ6sdmyvV+6klQRR7rGl2Au2KKEi
wmLyDlrZ69WTquGMamN+wkGOMSeHTf8XY9yQqQfvF27LIVYLXJ/zx/dKjEEoMkFb
iM9FB6cxZVzWCQll36N1ILMUTLG1ux686pZRXGBFwxA8nbNnnGsS1y3HtEMUPkBM
ieNGU86jXpNPeAYyhjyVX6sI6CYT69M9AI28Jdzq4MHPZHCzRrh449qv2NJH48Y2
h248tUKHLLOb1GZsVz8rtLRqochjucvcgn8/osTfyxT1TPioav92Me8ki6akUxkR
HyW/zTr4YBBm/dqaKaIm2CmUO4h5j8f6BVxh1USXsgYHMjqxkQuPqUobocK0h/PJ
f//7Y7tDJDEX03Vz0DSFChhn78LCZ87d9YUMcqQ80hzXhxIhCDb+/Iw/A4JOyWuO
RBjIK/cHMr8EymWsYOFGe8PuhOaWYW7WIjUuNg+ZVVv8NTjdMfwlYOsAkiukktg1
EBen3LGnU7n/FA79a+dNWsSHyEmqXNwxERH7r4UJtW3gncrg3JWqaUff5ywDzBcX
kWOapK24jQVlZdcb0e5SQZ0u/+Zq2vJO296hI9r8e2hJNnNYq9daLTutpZi0tVL5
AKsBu4snfy/LUJoJIFRmoKQJjRZPJarH973ZF+H41dVulQhvVREK18E3adGb8I9y
dBa7oG0SolaorwV5sLHcmrFg+W8Zkzh3de2i7O+kyptahXdqCyg2GB4iz8iE2Rut
XP1KZcpjpTZDltarU+RZCMX2s0IVw9Rt30kJfiYZ+ZmVoYdvey/Fi3k6c9oTCBD4
pEuNrbmTDYCBeYAmFZb6hg85l8U4UaqOTsTKaj34sCRwZ5wcxCku1SPdh8pLH0Ir
xZdFWxa2LvlRN0fiYMtSO+J99tHtnz49QpvwaaTp9PZCTAkKH9VdxC6nPA86UQYB
UCz8XtMaBlUzIujbj+kdPqBIpB5NlEppQkXl7GsWYjQ+LOEWhEAy8IIb+uYspj0u
VWR8YHoO0+0VJbJdxyTuBL54TktRt3FDalKlLLT4DnzkCM5cGzaVBnB12FOf0Utx
dT8/HzNMZo/sYsOjk2CUnzM4PoC7kAZZqLeKkC5LvfDYPc6tBm7DX9ZohqZ2PZny
PA7Ff1ELABsdWUQOoSayoyqoMLyHU3HqpCc/9fdZgfVZiyOFjIl9dhSnYZ11gnaS
ylliK9pAjLjtqjluZuExl7jgz0E5gH1Z0ioLne3yvLfNXl4n55bdyVlvinTYKW6F
UTBNUVXwm9TQKXUDFESbkv0uZQlezGmL7PxkOiTjlFuwz6SRfoYq70TR7nA3mqQA
CvcWThMHbaRuVgahmorHfRffpNZcDDdyyoyGOrwOZdGwtxhoQ4i2G773QXnhJ6wC
BKhkEKpEdeCq98L+rVm56e+ve+AYyK2krFxr87PRUGjB1DzLQibbiYbP6hQBNZfz
L+UF+jA/4BVcICxjlbk+QhyS+q4cLhIRtl7VRkE02aXOZfKQFo3CQcZ8Jvuwurl9
tUNCWz94yQP5BUDsGrebV2xFYwAPI+Xm54j+e2xdtpThFw8zhnEV9n+4YJrviOXv
Ndf7HfgY2WbR1tYuLLWOvOe3Iq8wYtx85gXAlRa4oKaraStcQFTZfDywXhINrCfk
dM1aEdlh0ugmQqaCLc3M4htoe4V3TTFLutukd1795DYMODvQKtBG6kG8hMDQ+wA/
8i2+fx5zXOCwTE/JBXkISrKByJ4XCOYTbZbxzgdEn/r9ekQiRpKK1uiRBr0lnlE9
9EBc6Pe89qIi43PXcymmgWT7mD0ix7Fth4yoCFngbSB6BrSPRyqvSHgNtUl5dIZt
jCC0BjLfqUYJ3QbJBGjqLPVDfDsaDWLYJtuMyxK+Go/MOr1TtB1Eg9BKWzpvMU4X
+Db7re6fyYIrIALgmPbOFmYy+sOw9aa03xq/mSSzRoWDfKZH+G/pcTLu8W89U/St
Qvd3wfB+e23olC7gfu9pW5GXJxKcyww1Tc1KizAWgQH0UbOOupV6Q+DzP5p4H6hE
rpwhT/ahTjGRJkvpVNjvSEU+yw/VNxGCTnFDtoyVii0gIF62GR49XGtVVJ4hfbRF
/rgPNboVfDnpIIUYBaxAwRtA0jh9IDBhxXNwiSwHvotHnz5uffyQS4Jod7oqvMPM
LcWcOsMMz1jpr3rspDuLjX8WR1i8MHIah+iqX0hw14XT1eZeq6Y1sshDDNW1vxLW
Br0BkmqfDQbnk27Q54P//FmLUQZKJ50+mtnM78DfaqSrq5KRuHi3VNM5pFkyUhEj
8sAeUiietTmw6oCMjOwA5EwvTFS9J2TrjCGG7FzfiyTBWXw/qImd/Wh7vbX1Q0Zv
uNigIjChKyRC6ad/peGiYSGHU3bZTM0PYdlh7A6gd86j5MT1L+bJZ42pWaaAr//z
sb6NODREAWzJEVElGw4TdYL0NZjJJKgKGbn65KUvRcdt3UfwwlT8xUnDZDNFcpMA
NmctzQ2v72B6z/AdPPPY2p5Jag5a8+Vw7Q772BkXvjgyCU2svmdGKeJ7PI4xOrEG
CLdA4d1wwKmK2djnrtY8R3bDMRUWjn/NNKB/nLtyxR+KPOXVCz+tm9wupRdWM1qB
LYL9iSSlgHJLN5mT7L+jVn9UHJjhvBed3ObqX5VRBWqObm6VGqm1ErHYgOUSBsVP
WQr8kGh2iu1pyIzkS/dHV+l1GZL/rs7jtHb1rHaftAN32Mvur5pTLtjtcZ1aiIQc
fKbXy70uxzzEzL6M7bjtsr/KAUC5ikj5xkLyBklrLDn5gkRWpeijMXw0xam3a+Tu
IPnephiy7583GWIufgPMLn5TNUfA1ysk51/GSISi60v+g4pdBKrc3KjW+69JtByl
NDO+3gwXb5iThkH+ohHpWo2uaya+BwOpEAXactRoASQU4RszwLCeiGfP/NYequjQ
ioNYOs8cfRPScOfcr47mZaEjifasMKM2yH1hR9DOzo4maOjYX/kcLd8MXD+qLfeE
0/KOHdun82saViLJn4ZYFyznU+Z+j7KAS5InITGoE9VxWFNwLRL67J1eA2wBSbU6
VsHvdQ2fZ8a34E7kdjrnGdKWlEmfvHyUQa+FWihfxGwmYYLO/HtnyTBPvDpUfCop
27/cN7weq7Ps+oZ/RyRH/JlDKRLNnpHDsyT7J8iPvg9vqND8l3MEJR4B5zypAiej
fhFyTi+UW72o2DEjjvefr93017KUKwXGI6ug9NWuopBtLlxk1Qc27ElEbghi4Sc9
v9HNrJee1Gfr89lzpXjh7sU4fKLeqiiFaVy0ZhBqQZ6fAbvFcwNLZaFnmlNds2Pn
HwDjE+cNpw3Vg/iuq3FHpdpd6ZdfLaD2H3+MH+eeQ4ePbgTMXDtKBf/LadpeL286
d1kWYjt37C1hTETjkz9sqJyDfQMDnnKqhdfsGXtWC7lkEmGyqC2ueU8HkWPR5Dsl
GEjBcGKsIe0UokociI3b87woxXVTgT2XTbhYTGshjw0nBwxsF80nty4RJzRXU7PV
lRN4HAvIxYms79dtf0J/kUdK8/FOYx4u2f6pvCXb+Kbjl37sxHQXDQfttpKskPPD
wiZ1VouhYC2GZfiS3+hYP0ppfumVeYltQ33e+Lyn8e5NyKJsYTEAHQeB5fiNMNRe
k2vK+1EP4jUj3Qiv3CiTxi0u5dpn6nivQdqFMjDJRW70rMJLZ85kEmGEnCkV2SWV
iqlbjIjsjmImN/d0Y8akCANVhJ+rU40rUBnpFKrH9Sp0zbyrb9L8u/gdxiKm42gZ
G6PAeJmzEAzTswJH4EUp0gypMIXxPcO0kapBoDLD+Vs93r0Pe8pyUNVoN5BoWzi5
Mn5sy/SeyKfMkGGbzujj+E1FYwxBhhcQJRXNgnvqrGo6/WO/GMijJhJa0xFxIvZc
0ETZcilj83mzpSFz1Gbnb6fjuR7339+wLAkZqkk4lcZFbDl1aXvlarHb2NImWRzM
vxeVQNzX6PUdMgC0ZC5gjK8vMIomhfysgUEwJ7zJRfucVRlvH8DO++g4koFHdc2e
LjxB2Al6c4TG3P768LFnR2gNXfydLkgHfAAjXJg3/BzxOQqN/Uf72wbL58p6Ls+m
lpgfeGgwfZj0O9kJVqpkOxPY8FudyrjuW0VKaiAivWjjpg+1h4rn5oxQHMDaKBVq
sBhcHFlL/+GL7dweBsYL0PtO8DOvcE0GmUOSzTehWGjNoiX2zWUFMwuH24U6p99Z
iKinUlTA8PvrJj5/JEB3bK4og+k61YK9WNQ6Y0WPdbX9sUu/mWMN1yM5vHSH2rSj
NHeXdgA6ksRUSu26kcPWxT4ZDzCLzULEGvAHpUS86YHMXqVNJ+2eOGuj/FOhsjmV
PzSGSOriC4HIdB/YoPnbY4QMLQBC5zXnBolvcRVwntBJi/zOFKeU7gv9SWhS3U3G
u4IkQE/jJoz4odorcdWiMEbNUhUyaQQQc+VeAkEarGKxLoR5tE7Dky+WuML4PAMs
yrfLJZOHARnL7PasWlot2UbsH6fEM5Icnpo5/n19I4aEQ45rndztGFPDDRRbXyr6
kCyre+Xh8//H0GJM/Qho4YwB03zDjXp4lkT0nhu9RlOvF7v2o2IeOLG0lRNQZ5YH
HK0Qda1vvwteiAwmHZc8uo5QsWVqd834m605uFfDrqSRVAyfhfCGHJlkVcnODL2e
uhOCZyyXrQFuVT7T87NKUATD9836qYdnAPaEG7AFJZs6dXp7gQrTkUunMZT5wl9T
wPVvday+Wyl6VsrG96+NBSpJIWYJrwOmWJfpkKRMRHL0tPBeFYPu80/e/QHC9Rt7
bJ5sX1VPuC2Mvo3D3kEXZI0XKifhrf6iAvq4N+ITCkJkjyqbU27GpiDkGs0Q7p6W
oVDB/8JPaczyDw2AsSqxm03b0rbb31kzUX/T0VShRuQPagrUNft1aR+tIEC+S7AQ
qxjPh/lH6ik9iboO+Uk1yCNDF5Z3vtBSj0PH8O6iTFw/KoFMb+KwKH5so9mWd8W5
kOXUGxEh+k5Zr24fRFT3egXXUWrXD5oirToZkVPvULEiopwE7QyEnM4U2zI3BmGj
ykLeh0L9I61WBFau9veGnr3q7FFU9c+bvM5VulVhpZF3s/SUA/qCyRQqZD4Kr8IF
5BC5iFYE+gclnXh1p0WW7Yl1Sb1d+sNjyQQfSWDBZLy9dsCv/3TvJfwCYklJs3jk
3VrHrxXRT7qDHnJ2CcDpcxWpQYa+5OzxdJlDEG7HQdkW75h6NUJh2/F46RIeYlZN
f5ETX8zvqq+94XtWyUwlTMetH7LSFdTi3E4ucOTPhoIhMWqtH8btvnkGSplxHuPr
AOs48Wt2GqsMfnGXu887F+GkGfkl62Jlg7vw4yQacr9CagikUH2pXlifnJykFvc8
J1A4UYx5lPHGrVrf98f5HyGbXoHKmGpciAzAsKrqibhYkH6ogBXcx5sa3jKaNQBU
9pwH5wKL2a1ej0XpWZj+ZEeAHy/DbFsNKCVgOBJBZVccovuUrfWwqZ7qzIlkfCId
1V+tb50KhB60Py04ZeQ4yN84ZcLRcswHGv7q6ZITKHZ+6OZ/iKxvoV5bVaBzHfJj
XHFAX8Rj/5YIwoZQuLkCO/YLaDZ0OnY0PyQ0fb63iB1pv/oyHXilTRfUodrVTFwR
EBTNJcPHdUuaaISKgWpMsMutzH9ZL0evLV85pEYjC1JMQfMvc6fQ7yEauTI/aoZE
3Sz5e5+AO5+iqgEnkpq5f5oFpSYYF7+8HydzNd6LYy8V7ls+BtDqIbq9wZpwymdb
876hxmkKZ+2WRY4Kx5G7oYjRgo+KzYgQqZhVKx70Mtiu1A0A6EIPyVcBC5ZemYOZ
E2LHR4uy+OdfLwlbxv5XFon7IiJDbh5cFXW4wVFYDP1kbdT6FTkJe2rT3DbIgf6s
TZxJwIk9YzsLmAWfxmx2suV7uEVOyRvBcuxov7w1VgdzfwY1IUyILz2Hnk4X54Id
XVGhbEUVAvO3OR8ZR+UWSer0y6xXUPjYj+cIpB1NVaU9ll+ZWzJaAYtsukBvPbS5
HQD/PzWXHPeLFxg7cwA3wwp2r1W9i0RhV503YcYGT9miZ6jjR4SIOybEdMDZWCNv
qFb8Z13ccV3pVV6siB2tXx0OuXiDNdOwtgXoV9NYAJmOA6DA9n7R7D+opNukrAF1
Xl5KU1hxGi/MhMr3pcbvQOGRcoGPA3d7TfZe8B5dGkca/VkBy3IoLL3K9XHtdqJM
MizMb2Di1Yh+obzcRj9ZAYCEQXRabUVzHgXpC8zA7lAgxUeUUPx2UdkgInAG3s81
YZLI1sTnUnKAIPXsuY16avlw+dfna28Gy/zrma+GeHx1liaOKERfuvpp1C9xZC47
mWXuZDnh6radrQ+FtuZ4rgFO1wADKYUsfd9KWS6O6TJzP3g+bnXBYFN2rwE8zw1q
HBPmGzEayzAs3XRz9IGWdLAPzqiWGUEOVDZTkUfPL2TcFvbYrHy/fDTCDwn+4b6t
vvdLTzyDXbW3BxPwRU5VHJMvvLk7tzTmR13k/Z25HGDGDnRzZa8071CcW9HybCHX
CVL76aUmV28ovZnPb6GMTXHChd4pjPqtvC8JBCrMvzTv2m6TElvXXp0aqMAm9N4z
42NXOeQvDm0TKArEK0GWJS10oUe4ejWT+kqEgCen+f88mLzuvMdS9LJjXF2cVVbz
/ikWiozA8M5xZR0GTk2tYjbIQYgWL2LYOxZvHUqhHC87kfa4M+je+Wyvz5AIgMbb
VZOxClSKAINlrEF86ztxsYXu1jfpGkgs1F2OndxJx4GWeq1JcLz/X3ndyjHxYnmV
WQa+3ILZC+z15rBwcbFOcuSA2vV+eVBgWHpQrrqTSCdfwXvlxbmDY8Uj2HESKwzG
R8I7gzxsuyA1PnVeqqxGav+Dm0eVq9nSkRsC5aDBNtr2Rzc7osVd8QFwh7qizC/Y
PBWpUa2T/wCK4EMCo5l+f6+rnpg86+wfUcCM1SPPcQBYFcTmlezkYkjWALZWWYHU
X8EWGPSfiICZDppWovzf986lao7KCo43KVGkjLlCsY0I8dYj3VGED3E/E8mHj6pQ
ulDt1a+a8AGurT4NdRPglVMVcjHqHl5ixiigmAmXuQoxibzUP95jcsNy+LPqwjpg
DsMvj0rHE2PFT+joBAEqqgPWXyCmN/wRw/e7+C2XNszLB144eRth7JEhkkKqptTq
7Lo36oeZINHsiZPBamPd0k1YU7jNxvH4NxE+bEmWRL9cdce3XvT7YLEJE/adzYPu
GerNZNIQN5e0C0QRnRUCjb7QVHfbeba1G676RJ5F3FNqNJalgYKSTBo6mjL6v7jI
Rsm3izVEFudNiJBD8LdCrS9F+F7s/MlegQ3K2iPCAWHxi+3NaiGAAagZSY/c3yD/
2b6L3cDrtBy+OZseyhGNCIUXR+X3aCLbSbMnL773Ad+IIKac8sHgEidIrWNeBp/o
wd5SHkkt7pV55kpvfv5DaJmU0txSUcu1QT4O8ZyNP7Lx3jSC0UTBEtQnnsMh2TDs
l0SQzEOyg/6QguT4X2/WxgojYgj/wKmoCXjW78SJ62a6YpWixhb232P5Mk7F16cy
ZeU0draHgg/0nQtb9tWIp+nWGMkBP/LZwbWcEaYlYTp1uvdAtVAEy8iZJakAegwP
iWtexwkt6MFSsh2W2I31HthRY3SsFEq2KC4M+OOy3gaDuXOmBM/P0Id5IdD6bEbX
NqS1YZypUQ/k9SDBbmYpCKjtejjs4cy9CMsTCHDyk5A4LP8ugSuZKzoqIOcPySRz
HpUgoEe55Kp9YX3t9cB2eT1jaIA4sLE2H+KKlC5xOqAAS0tjyLPnklazZ1i3rZr4
kO4y4X0vD/O4wTmTgw8rpcTp2BgyO4BFsAiWOFwulYisJh4nJG4kXB1wbKm6pvYU
A7Z8/d7OzPx5HBHbW/mDJc48xWOQWH68bb63N1LOjWQHTEgJTWAyGkkugTIj1c5F
pFMpVuDdK3BM7/BUefE+oD6grf4Z8ZQZcTiZYs8H6hoj7tnplH9bSixfPiN2iqnm
H3VImrEZqaqedyAYH0yTs7a6ISbGMTqlQNLSBXslmKxxjQbPjM8NVWpCKREDlkoF
QeyyyB4pVX5j4fKul6FRWwYD+JwAoMsM7eD+yYXSwmXD8ruSa9O4O6zn8ep1tFRc
7CwRCq3b+YJuxgAIbGwxe8j4fQxC/ZS7HAqtKeQbiZQtL/+0m1LGiDtM9Bsc4HI2
iflEFDDTXW84+23XCj/p2ehDc+jzK+mBUVS1w6rFLKDMa5v5HlTYe/d23woQ1I+H
PGb4izB4YXSMmBc5366eDV7W3/XVgRiZ74flPnIbJB6cPKSDiT8W0d4TTpozwA/k
iNllPvyaud6j62JS2OlV4yj4e7qYPW+DeSkDTLL73dHi+6EYBGOFghYkElhB2ruv
7juulyXlxN2ouGOpNIpUtnaXGfeoEnyDDhtDrjRJmb1GetFxenujH+OPnY1LTJKH
cNjyn+vhiMs1Yt4x9XvsIaCkThF6q197iET6jZdtr73GdLD9F6xMQk1OgvkcwD6U
YU1CrgUB4sDFQPIbVyfWIh0ehVjbJzShfJoan6wBpwLSUWDF7lrfR7ejc22l09TF
w4j6+pEqGA6msAr40r7Mmq1ECNDmqQRAILvfXraUZQI3/2i3VtSKsDHjG2DOs5AL
HUX5uCu8v+V/onFTr7I/mK1+K9VMn2is60ToAeX/UxWsx5/UD+f/jixFgCOvyxd9
uXbZ957079z36ITBUTRZF9QFR1r7ZNKnIRsCq2JkMyIWyrMk3BhZdC5lhC09ESr/
8WLu0tXc5f1fjxw21OD4LNzeFZVu/iKtRalDYLfIW828oTCPeOtLy6MxaQfGiKTj
/BRmIp7bxAiIRGiPq07eP6FuJuTothFYT4CsU2KQODm3Do38+vHtbnP9J9aqUrgK
uKZD7W+GqrVTLSy1K3d9PiBax2FSxXgGYOxp9yFkfFLuFpdozCeVnEKEiu8MfoRl
RyRksTuL5tHG2mAzzoZRme13693c+HdoZGLRJP4xwSHIQWyEEoNpob9IJP3Po8gp
Ctm9QUlMBIc5Vy0MdreQmD4FPfo8Jq72Zt1f0b9ZVAl3S3CTX5eMIXb3UHqXoyh+
qMXQur5h4wvmY60Gsehz/jakdD8DcVCZODFhu1BIW0Bpr+s7Rc8/X+J7FqtHMKUa
YCdCdx5gK3qWe87K5YqZrnGMf9/z0CdPukFM5SJtcs3Eb/a52Yyr7kcenJOVfrJp
12Dush/rk3NXmcUvA0F7A/oOjpXRZuirRIugeurQbAvZdFs1nj/Px5AQw3zt+EuA
SeHY11Le9+m6BbtpzSSfd1yw/92ps32CDDgd544/OFGpyeXPspE2nDduMla8LOOG
rt4K5JQI5MNZPOSO828PeqGwgJRtaPz00RSGNUVLQIPF/MRl4XpL8cTmR7kUd789
w59rhswO+bsE9Nvl4E2vNMbiNeOIVrV5GJ+9tvU7PxUFj95/hHWWqpp21RbrY6/l
E3mWxwWl2kaDNez5DVhffP42sfU69L1lKDE75rhep+zd4XhgoxnXy7/R11itMKsM
vLSAUZkb/cPQKoiHalV3AcrVZ6Ajge7XSIxtkbJ2Ougyjf0omm/GXwH5nGA/wHfp
T9yAGjUQ00Ulfa60xlE2bLQCce8ecDCjqnvg6AaHQtFApNW1RllELGK81oJt1iI8
Ch/rk4ogeuTDXTmp5swhX1hpNy/QU4UoWQ7TmqgR8WVu+s4M3YuSs5Ww7UI0a34F
qvP9ibmWuWx4dMVBdtSBy0p3tavAkc5yy06BJCNKq6HZAxPQ5P9U8paNKnTM3ojG
nij8788+uUH0/C4Xcw7/Urq8XHcaskIIBz70wYy/tdH96v6QsPlFk5B+GC2lSJmn
8piQPbgOZEcQgYFBR+xIaHsyNasACJUCXT/xAvAoVZPI46+2ohN57ZUstgfAwpHf
o5a3pr7vObicikJ6kYwFVIaEL88IgL1ba/nRXs4zt4HpiQChlUiAtH39lmoCGnpA
+FxwoRMKuQjCjlvUGgLkSKre6nfn6dgLBTDJGr/n/J1/30pH9ZGwh20FHfd7Usbb
Fz3selFpdnUp7Q7GwPlmN1KgySVlThWyj/OzzFAJTbBippFRFK5pkUAW7G+w/Wvf
6KHL1XrFg4st52yWSG15trwj7knUGqcD8XVprdCStRFVi2yE0x93b0li3vO7vBQO
6P5Njncf7C/NgPkrBEqmRiZDEebZQWqEml1/83OvccgumbhJ7DKyL2bXgFXiwTXC
xRKYf/qwo8+mCgW332HnNXDuZsyrG62akZciW1stWdw/8VX+KETjbIPxFt1Mur7i
MTlIuXFgSEo2lkoJl0xt/p34XufWSYPl9XujIOaSBzFmJn1cKflair2uA56GECLk
h+GFVKjAjcrF9JHeEd4fwPZouRa2iacBWlTENp4rg/7gpcSODYDM3Vez7NOriUp3
9vmeqAOxDh3+q8P2+qdySiAvxVFvW1qwVp1Y5yzc1lt5psvEJiDOxxu1joawm3W9
86ugjG5kARkUUW/FPHnrRDJi8bAqBEBPKRmgZSIMvgaaMf0ie0ZWEuvoiMdfqfHV
C/byJ4JHyCORdJDctL86AQ/6IrO1L6bDiZhPjDKtqFZWjLB6gWC0ZyYRxMMSkSsp
7sqW5htX47FIIMXQOTcLuvbuALAzbpGGGpxQ04kb7hgAZQSiueI8tAEroziaOMw4
Rwakcumj/p9mzWFuV6RyCPqQVUnCit1dW2kczPwqMywjEsY0m27rfWnQcsmYNxCr
KcVD2ZMyW8wRUEr/zROjmFCG+R9tjedmdNE/I8uvk2f5tp84Rf2bRhPief/a06Gb
OwFC9gdd8jpdTnGiNi4QtCGb/JAK9/E2YGSc3jcF6llSUMkxYHLywOuPPI2keFGO
3OUP/Q5/lHEhUiYeGc9nRcmdYvfWU/vO3UnBOgDEuKd+arDOCKExCT1OihEPwh4w
K3dGkG3ZqMZd6YoIsjaKXCX4JHz6SXnsbcUmila5fiEwinTrgMcjyEFI2QtZeCi6
uhS61xXo/LB22CSnTptGgTbbEW4hOtRCKUkWFF96X/kCCcaq8Uq/lNwQFy37NcG4
vy9Ylhwz4yS9oYaAh8LYplAkm8WzDsh6BnBwjkCPAbSiQxKsS8AKtnj77gxIGMWJ
ZczDsfSBLVmoZdpSg+xrRry4U6r44cWhfQuabLErb4EjznMvcnqWNCn7CjnnDGMb
KrZivKsv3vJCsqtMvmvF0WStSr3hJ9T1SIjjTBr+CVo4CiwFeKNeuW07BdG+DtzS
9siQ6RgJ3PDsAFW/tZ8lyckY5cc3Up6G6v85Nb/F5wI7otIBQktskKwvNitpEdAj
kdNvy4Ww1zJd3MQM42Zz0LTlNQp8BbC1i0bikImEO8uakBxhDcY6YIHs3pogZABg
mKLga8YOksJEQKx5U+A4VSHqirXAHiDo3/uaoAaf2b3f3LRQ9WKb9uYOK00Oh8vh
jW0oegc/KP54pUgQz8W63lz7dM49QWGKCY4iHoZA+ntmA8ZBszB6Z/4mSpTtkB2R
rgLc3SFIWxuTYySX2cuMHkolRUMvCnK0leUZbiN5ogaCT2AK7wmFjJMlnDXNV5mZ
+RgeUr6YqtY8TkxJwCC8QaCUetlQFfPhhupWohyJO/V2fXOFgnKmeix6vNFuaQzd
UlHS635wOvD7bHWkIS5TjvMVMc++PDBvinTM3QlBnlOEJS/wPp6nui+oSZ+CdcLr
Ehs6n04t+QfQE1cA9URli0Js5CDStYPwQs59a9a0E+ABct4z5BQk+/UdLZpvM+BF
bUs61jFUU2OLzhAL0pg/aQyrdVYeJADWBIHzxg8Shh5R27bMVxbEM41jXnnBrYDM
b6RbWX6njI/WXbNYVQbLQOFOrJ+7Vvlf6mCxI3j6hnkJzXIx+XqTWHCsf+n88zHH
BIAmdLr3wk9PQcpOGyp/Uim8Zip4kmo68D5OBy+L9aLrQuWHZz0l0434Lh6irWsa
eYDt6F55iXPw7BU0Vg2oKMjvtcW3PD45W7qLs6DjjhIkedHDrS2j0G97/cJKjQjv
Q8YQAkSUA/KCVy45hZjIKwY2SE2kyknxTua4qXp96XxfIz5mqxfnnoBpqWwwy8Cv
fxcxixjnSLzVE5WiZxz4GYa50PMJX5W+TYwi6zZwrR9fHkYDMsdXwqQ7ahMAJPNu
2/3gKLXTYkPcGgg9wATaQN4V0lX1nN/Oetn6EpYcoS+9qVFrdqXSPwSvWhRjYy2Q
AteKogQWvNiDl0LhBc7OJqaAZCIHnVcH19rfmHZgByuA8q0z7NHBRQW8WrMuVvQt
IcFE7ipJtj1Ow9fVQ3D/juS5olBhJMWmRYVJZAQ0wpwhCBIFD5WQ+yPVmELZcrPH
uflTodjPHsb22tEDW7fEqP7fC3u2L1unq7P5NduhisnkFbQJAgvDXZ2kqCZq8Avr
2+bhuELyBWC//uuCj1i+n1NnLu6t+KrTosBlRcIUEiTM+q3z1at90Jvurx9EywtH
L9jL9SPxMmtVApvygzcKwYKGo89H8Df27fsLw3YHybd2BuCTravN3h3i6KzaTkWP
xLJ6TFZ7aVWdkYamUxeXxYkhxGof0um0V8Vp85g1EPq8k/U8rRNUC6xcG9Xmqzgc
uSgnnZVvV/OwezqlVqZMT/4QDQ5iC83B8pFhfrCZfGTDWCLcGjybCgDm8K0+S4hE
/G1O1DwfXG5Uw7Fw1kRD0dddIjNlcPBXuqEHCNMkBTruT5kbBqhRUz3ghh0ZoYx5
o+M/pLlghZanAM2hbAt9rgMuniCOlyL0GOwfRMWxVfD9ygMs8iGjf7dLl7ZQrCQN
eXcTF13gh3CV5rCNgHc/1mGTDxDVRObNVnireThu8fvLbD0CEJnhy07vdi68CpZ6
Y0EWVDqu1GYO4HpAtLuSfxelRNIh5+PVHLTp131x5E9rERXAqKSEm02PPzZ4CJSc
OgOfyyKmAnOUzhdehcPUaeaCO+cLLZ3BA4uC/PuRBGyRdR0X0+sgay2RnzoQHoq0
RGe47SQJR45bCocyD7CBGVNVUDZAb8tyPAE0a52EnaU8WX+9DDdvEThFOq14B5f3
gHN5esFM9PAp8/0+cllgGvM5IlORfX4zKT6Jz4IOzD81QauTdy0Zkz9mfSzJwmPn
fzFjPzqjmlPPahGlhXWqKAyWVmDCKU+p9PNyza9MyJzReRk0izyD12HEl/gQREw/
3MRRW0xbVeZuPTwNYXXJx82zecFiluSBY660JJDe0Q0QEIgbZk6q0UjWYRY/QCVN
vg32IY5R+0c5dO0f1MgTvg+UMpxM0ZJ+gWpc9lTZ+vEwK/Pr7Le+343XIjI/ai7X
GdOd/jFUevqGLBb1zt/aqfsydGKD0+Bsnpj/l8Z1BzAHVq8+YgKx7JiFbxpvDHkH
0cIU0WbfSH+dAMCPMOZDC+yGSW/PddPyNUPzOxE9cRdVpktVsr6yrknaR3gladzB
baM7kMAQgqgFzK8YmFXzhzvV6JEh0RK6g2ThMIDLEe0g/1RN8RIJgN/OlEl76N/D
1lez9Kzt+4NBPRJWmFGnLWlUCU4qzCSuSCoO10Tcii5SYM8iEOvKXNMJGyy9exSw
T7ytmRA7wHxB4DDXHPL56QcZrd8/wRpS1fecs0+EfVRMf6mqoQPan/0vhoQ9/Qmg
O568pBIrjUWckSST26FlXF1yPAqyRczeObCeJ+/cRPIMvOpd4MeGGf8PsZg3eXkh
lOA6uucYoo+FaSNYGxFoy1un6YSv7wzYLk6m8WGR7Ph1HEkHtfkdXZIGHIN/JUwb
1xuW8wxDQPVZEhsTeecrXkIjSMZ2Vbvfc7Q9v7yH3cZ2UrIRK0sB+1sBH0VctlAk
wtn+WnqQSqIHFTZOmNy57mdDSc+2jdCNFWlFkmPkCBMinuZ2eoi1bPqBFYBQsW5M
eEkQn+1E+WmESrUfmdE6GFSgZaGbZUTiaNMFmFrrtT5phH9s3vpioJVhiuWMgecd
Idb/FFuJRFy5OJQbO6nzHs0TpgSfmU8NymoJa4Bu/MmcCh3nEDaRpUpszDPLdX/+
22mbpGXE83gBKVqmZtbCA8Ew+MOAEcPyYApkJhWJtuZ5QFntOtrNE3/1fqgbDupF
vvBAu4YEJ46HEYvuoHjzTRKgsruTgJbQmxlNoBq4W60q06QdjmEjtwAGia+KFOLW
3NdIC7kUdkUA52BLNhQxwgLID73KIuKACe+CjKDNQzHmApk3VBceEvzwWIj/+uNZ
HwmSVF27bHh0cD2tx6PKHQQfs6Ka4dZ6ZoyVm3kQaOus7HPJjdYW6y/4I3hhWv6i
oQS37KCJSkvTXwfKgihLaOBj/KTkp262aJJRcRw9OebQwx8qqIw+gyPNWgCHiI5W
NdsvwT2QtSzgO0CmWHjzDaEuJJRERU+yJqe58OkYD+0Y/NAmjziW9DfRtkCUXMMy
1zNEKOvDWqkrzbmYvxfbQDC/luv4Uqun6UQMa+rinulyU51n7gTiTY3cUpGMGUwZ
WS+1nGGjYDfCSfQkQJRGJ7fJ4fC85+1G254iqAt0Z/oCdZHBsrHThPZwSdpJKikb
ocSaELLU2iXas3fIxN9MxuEjby9UhquA0peCpGZ4RWFe4w/YeU5761ub7Bvm2Ufk
VeF/dCIrbjvXS7miMLbi6m/ldCbb6QBPb3hic8Jyn7CzQENjI1EkGC6tDAfFZ1JP
S50eEXIjoJ6n2ucoBBQ8nmh93+CCzAtezDvp5ICdpDy1zIKgnro3brydpWvMXAcT
5ZXMOYSYbiCPZ+nPT2eE/u1DS7fU8gLzWtufWD7l7KQS319q06bd/i6h+Kcwu5rn
47w2xJW770FFl9GQWbAO1aDdDwt0AGRf5+savP82J0eZ6NLFwrCSx1zmlu4wGyGN
wOMeJcx3koWkM9meW76Jfx4PjrxNOBZ0+oP9jXJL8bsRgwocKkmExgLYSxPyAyfw
8d69zx3aPpKmqSFmsKJHnGrDG5O6Va5onIU9Tw/V7hHpzZipPdD9MYcfGxUBbxLF
figm/doYRVY90hjJyUmk9E1rS1jXvtqPGKVr2A/B6eHAzskQA2KYnXmEyL03hv3j
4T2YbdXLy4zkDUV0RgzKD8ON3tpGAGAAV7w+CB/Huz5Xn8LxRJNzsxISddTABi3A
C5YqOARvfjFUhFBF4ja4EVY++MBSgaL4ykNpf/5dLHPXKo1EuxX7EyfHYgN68pt/
y2yhxMqWQsbQ4wBk5EeUA3w8c7q6RFYL7Hp2aY8F8fVAG6EF8Fca9Ngb8k+QdVtd
gKwi3dbMwwMSijUA7VB6dsy+8m2sW4C5XbgLY4QBdtvUEdVgtFd7Ym0MdI9kqjgd
xHAFXIYCZvquzwaf6fUa4T8G9xmCWhAsEayn4CuM4Xm90WtUgBs1KvhW1un4K+gL
0dNrDjbK0VP2YmkBUQQDFPPM4/fDrFejLyBFcVBkRGXjbZnzH/56HmdBlqRVMhXh
YoFyjZVagrdzn9gkEvMql5TPk6OL7nQKK6RAK4e97iMU7DcP5foEYLy2bTWS9pw8
gF9QWNkCOIhF8QKSpOILjUrPFCM/MZobwTLxCtWMIQd/T6prb0aJhYltS39jgD1S
zh+Xe8pPzhrQvtjZ4MMO2kh/CUdRkfPvj9EtcMX6MQd30sadiYpBhJcDnCRJftcw
hgFJSdsf2gU/vuFCmj1hGaYXBvXeIh/fwZ5XEuL+qauSkAABKDZAcVc0A9cJxuw2
tiRfJ2tAmZL47CD31DUFDJ3dVJGNG08ez9+Ht5S32KeTMT+zCvWPk9uDw00kz2G6
JZuLQehx45mRHKUETdSmhrirDnj14gJaF6xhOFEMIfhYYoNd9Cb9kgYH0vlQ0h/k
+xtka3lj7K77ZC+vZL7VR1oTQ7bWZQIeRHY0lHNNDRxamM3+XY37VZHL0SYloc5V
pthYVMVvpMLUE3OIjR61sS77Rs4PE8xlDl7FAiOu+LSGqqf2L3b/+DHeYO6/jXCj
aTfS6wHY93K057J0/Wi5JxkZwrYgnKFMxgcX37Hg8wrbtGBvFm3fGo8IkdN8U985
JHctehInjXE2TkFJ16DN1vnyDLMmDthUPxSNCbHRAxLOgNKKdNnEMK3frR+AifaA
RTovlOQ/zllqxH3wMuUmXkRRtxo4gj1yIM7gLZJ1hMbI0UUyTU/F3e5Pqyfqal0C
V+uEEanDY/Hu0PkX+SICYZB2aQyXPPwG1HpBr2lGzYcnE50r9QGgm8VPz0i7eLGo
JdM7a8VVrKmS6YsIe+NvsDzywD1dBPikZZ7nvuu+VG9Rl2dc7GW75KGlfbohrKzr
VjayM5FxY3NUCw4LwnF8E2aDgkWYk6wLBCLSCz3r/xpeSKgh+bPo/dukt+ZipcsG
oRgNUdSwZCmg9cHNH/BgpwqC0wFcNX9I6bHb2D42JPc3hjI/E6t6MvhZvZQfYMKw
7lt7nYRESWtizf1AiHd86H3gEZejgYA94YmHwbc7VM91YFETIdmqPp5WV+LelXXz
0Q7qdjTmbyu+pDO/ZUVqUZfmG3Uaa48LCrhVnY0+NH3dXeYYnRDxUDl8KnAOfwBV
04ccki5FlmPUsosf/MsPNLKich9QXZsO/da/QC942FIrrK86DBoBjNSnUucQVGQE
aBwphBnf9OW7EF+qpPjsLctURzA5cqdZZ2O/Ihn/qOnWuq2Joj6XZIYfEdVsVRHU
GmWOGOi5Wl20R0mXIeL/8dNuG7ODlVRyzDMbLtjLdJITQA6sVDMlLd9WCyV1DjLe
mZsV3m1gfrmJyWFRO2TlOLsG2vOq45z/IcCtyocFhwNTZmi68glAoJV/vK4V3isG
WN8w2CcZSTAMhhwYAsQwsIJXDOs2OnoI7TTN6/hpjEf6BO2E65d45sQ0gV3jxyBQ
tDZjr4JF8YsuVhdx17AUUtK7mdrIBOF0AWyJgii3ZdIDCE9BiiYyIPDA1gC/TUpK
iZxgLcEkQqI3G6PQoiDGUGNF0aflz6De1loJhUlIEimo5Bb76gDDAErfPtHOVNPt
Bp9i72s7QuQMHGUoy7cQrhro7+W7vb5kIUhBFsdmL/2VkUMraGmd/qT91NfqAwZ2
u2Ll33rRTXzPYdKm3X/NcxmaAX3h1BdyJJujvIc4JThW95sWqyRXs6Nk/1sqlTCH
43KeDa+19IQuVtuh/7voBUvZPDV0G+J0teJKnqNiEPbWc6xuuIS9UId7f7rqvfxn
0oFLwXr197inKwZ7hdG8bcAVv0itaBKnR77qv1VOrfCM/3Iic/KUJprFAA92k8HN
ue5er2/fWeoPh9JvYbB/2ZHn637NvrrJx6dlXGSM0CDQ29UDkeDhLeRCytibIMSu
pB569jUHzXS+GhI0xG8O5I0dd8EXqjEzt2Lx/vZYOPjPZ7ycocRF0EV261J2MJZo
RdNriK4iH2zq2wGbDbH5MobBn9pi/cWvSQ2UTSgu6Z/RX+dOFl32phqIzM4J80fY
ZRuJkju2pD7CukXLluxhdzAuI7DU6c1gvb9WHThTo2EjtboY3e7uITYCEoDeQXvo
MwuQ7Pss168s4eKSARSJK5x1RXk/vqO/DAB+XPnFo6POqYOvSzpqvrB6bI18yAQp
77MbFMGaid6gPBMjtqlazRsmi7LZMe7MFAZR6qlPGbpYAEJcHvUuhwCXF4HmeqP7
M7/lenxgac95jJsg+SRTZIAZrlu2dxm+bkTv3Xo0B2NW8xKaBB6DgGhjYJsYFcii
pHQBua1gEAR/alttC3a0YMA27ugyfMwlHsodCQI5iXosnHS1mK1tu3FUmn4+r/qu
IGLTV0RUg4oLFX+EFFmI6zwT+wLmJV/0LH1fXILQwn2KjORmOOM/YCZ5UTZmYt9u
PevebYumXpr1Y6fUJb2O0X3RmDWbPUOHZ6HPD5MNEGVOQNncc1Xj730TKwlBgPnN
/i7swJqttTqfLw3zjfcJ2zjZeWgLnyj98jpXVGyPJRSwnhp571YH3882sjAJEqsP
Xa3vQ6vjfervS6+6mbdWd458rEQPriuwcWTB6J/0YXkF6rOPFwM0AopzkJfdNKJw
waAu4lqnPvF81HkVO6854sH9YBAhmFMe7g9k+emoW/0VvcUc54aGofbXgAY/D5/Y
6b5En25yHe4VHdE7i965Gi1DTkkllofyO6y2Uz6xPDcFM6UuKcv+DBjasn2UzLFR
/A8e/A1sxZNORpOpXUOPG+V2chRNh90Qt6PvT8GQ2mqrJdjUJA0+xhp8qseOHHWx
ujqE32JVrvZfi12h34sfKA2qiHBC9ighjBsA3eTa9Cs9GD23vrEfUFkAFODKngQP
VF7cSv3UPUkghreIflMIyvjVHxfxLLVvxx/oMunRtUoR8Bv8kwI+PgU7zT2oS/oU
MQHVoY77C+78qD+fGVoKPAcbVcCG/R1dNTwd91erEOJjZf7kJq7FHSFGwiakG+fh
aXnLGBHpfhGQNDAuKEhUe/5l/UOefMHF2bd5q+0oYFKU1eLth5WB9cDrYrMfj92m
TPzQSMI/mGchQwO/KKRa4PiNx7GGygFdic71yd/5jUeqFQdN244GWvQU4vka8Ape
HPlEGFL6XvKB5Ejm2SbwKJOAG/3vqoq7t3uhkykfVVU53+iN1rubMK6JpKVk+zNr
PiTNlXfh7h5NiM7QqPhn/ls8bbB7s3ZQKAR1cafP1fAe1vBOBLXY9POFgM9iVOZC
iyhOkKFefhVJiz1SA/CkfUxiy67pZ79h6N6aQ3ykzW5KuTgApM2dCmil7wBknJKC
z0PRJIPa7O3UCJjralkl8LCNYusUPLEWFEq3UgWNc5uZm4JZYHPWrpgmV85EJNEm
iCBGycUvDCBwNwS9kGZTgt76V3Th6Aw1LxU2fSKU8nA3dmUl0v1siyR6lgk6FYqe
FJkMwWdqAHhosGYLwZU+Yz6jt+RwTo17M/GFlY5t7H3cU/5/OH7FalNdF2NcBhXv
UgbJJta0vjFgxE21S0v6TpRx2uDLSu2c16BEQb642rKrxDI6weqFjQC6nK9PUpRQ
Gq0kT06DUjEuvr4ceFIPs2MJrS6nJrTfPkmV0qyfb+HlM8RzLqG2sDm9jzkJ3qBO
/zwHYD7wl6RMRfX9Do5ODrMd6wME+jc+ksj6SscWgd0cbEDQVqGkZueCSLkGgk1L
DSEUVqcR7GmUFP5mFqJRMsyCD3HnTyA2jLMsmdiHpGgTTmtxL1BmeAFxAZYEN80V
0hQ+6d8y4BGmRRlA/JLQGBypmSVYEBusbOQ4ILGabXo70qNKt92gmMQsxScGCFmF
Qj2YM+tLZCun2r2JZrJ52OxzZj69aUU7SFUVaRn0RLHPRwq8EIq6ZkohxdpYEIJD
W5PaUuSR5BJriMqfImn/OjLARzdm96IU2iB97PUqIb2BO0SSmsoEA7fQu/NrII9x
PKv2Aio2LRGWgaPehU2/AbUfpfcU7u+LgR1uO00ZD5+KNjftOLOtg8z5S0C+7rfd
UlaKcpHcRRcsUE2VlYjvwGm/jwvx90zIMjMmT8huCzuFt44tHTiK1a+XxGNRGTQh
jPLML45cZQd2pPK/KsJ6lJbwrPgVXIaQ2ebigLDhYdHAPGaHanv2h6LVR/3YnkCt
Y7yPpPJwCV9xiAHiBuLhLzzt9/oTmrpNSPLMp4n1g0unDzdMaNteYqPGqvzIvOeE
3IcNLyoCahYipb0xnTc6TkbGEZZ89qc4+4cUHbmFVuAHjMWppR5QqUVLAUK/VrTO
DS8tHkM+yaG5Do/un352P0wxQzy48Z24Nv3otLsRbzSSKsb7AMBz+LHlVDn+g0Wh
4p3kqO5MggtOv4/eQEfpeYmHCgMsyEjPWw7RVP4MtPJ36DWOrt3VqcvETjh0ISou
26lb7Wjyv7I2Rz1s9trSf7uslIPdHGX3CEww7cLGN62nNNva37/x1u1NAluIAmI3
ekwji2th7ANTP3EJvSe6RhtC2I+wSWf+4jXGE+GBAD4GCiMNRpoF9WrEU6n1ZvYr
2nfDuQA8/48utEWc/311fdc4XxEP6ZO/3sQJyHHaE8z8FnP73KXjN2CKmTxCtsb9
sJhQgyqbJq3bALX2JoVgdaXH1InyohnzDEVZ0wITCkfkasPXKU+tF6XpCW+bd8My
ZjL5MPG2LK2owoKvwP5XYN/yfrXI/+HY5h3NYniy6ItojurJa8gnHyyMTvGrtl+x
VjY8GBhSTCVnkIMcbKqTi+3w+1yahRs0F+8AmReNqKd29Q4Xom6wECPbSzXw3/1v
boh57xpD/BxfzXdwqDhGAYIGfv0URW4q8aLB9fisOUZc+Vbvw1B6eZxxmyBbt4Im
OmH3B42uKK0jBHhdsMUdAdB5j7i3dvWeYTJlXF5ZCNu7JHZj1Rt5velol1gpnOzE
fBd2MtTohdcarW4NXb9KDnIYSvYHwtm2JRQYBSrOYUXMqfJB5VJKYmn3NpGNDlgk
PMrieEmcmP+p4U1FkWVy/bnegHAuhIiLkO/mMftkInkBUHdrb20MJlKO6NDVsrWN
bwI/ey95Gc0sZVhlKT3VSo0WLkBXzAljlzIYG+5scGO4axDmKr6IkbEbhSKmBIut
zBEJivr3YEBjr70zuLsV1QPeQuDHM/K0YYYF7wAH/9IdJdEOiaeM7+8vmfaag9Md
7dGGMTc66JWsmVWzOA6yDzJuio76YUhuvpg4+mjjm3W1w0JVCmN1KDbfn1qbCXV/
r2+EuVJ2wW3DF5DdDBxsyw5y3jnW5PRQWu+3mcO6hYzCIxr43OAS/hs9MAo6Oa7y
7iirLHPfu57nQLoJF3Gdfh+Qs1Y2RqMlS3mBSGTVsudNm27b7WC2md9tXlzACxMi
WRjr4Door90gjTJLemgP6F7W7bRuxSSyrrCIeokJx5wNnjiTBGDmTIQO4WnUcqX8
tHG/vJB6WB9KKbL3Wf46FiDRTTnmgz5Y0WkaR9k33nZXqPw6ZuzfMPq1KaEbO068
jSR6ox4vUIg6DHwFils0rTWem+0DakzsrfgMegIyY/AC6sXdtCi0zU+HhpuUFA5K
l3DcJW5UY/wHHudrChT44oGMd49zOcw6WV/6fKwhuT92U31hVUwr+uZRWHVUqgSO
8Xivbafylbk/2PAmclu6v9OmHx9aIacm/BsJTlnaHMlBoGLQ9c7AM/HQxg8jiaq2
xQWt0tVl2SmnB488FpWOO45BH8dlnV0IgTqgeZQ4omTpaHfa0OT6tDVfFkzYMZ33
wzDrqOOFtc9JNE46Y/OEsRYJ4T4R/GJpnJt+flGFGxcaTAnwl7GOyad8FPXNdun5
vfxGCUu48EYEnceRuZIRTLHtW8XeYXeH8+V/MxbfHUUZFVah0NJaykNevYWfJzc1
hcq1Fms/U9LDCJQeO8Tvru5Rjb9ry1VWDjRy+y0IRRGa2iMFzdzGFbPSSiQzcoBi
KCdBDlwnrmD26UVvzetBDJzozVmDyALGEdI4GyFiML7Lo3/22yF6uEn3zKXPKABa
S1m+BcdqPLO/aQSM0p9PZE2Nir6wp0P3DfYsJXd7etkR3+imHtcZapVPzrZLKZqh
XGYi2vsJzhOgm27Hw3+6BlXhr1xHKwbFB6T4hclBWzTQgdrnanzBqxyFYieIqWYt
AhsuBWTYU8o9FGVc4s2DZsXf9XYXFIfIUsO85PSIdwNZzzRVNILl0kuwy4dMGk0y
F0ukG090ssqD4uqK499/AuOzKPy4wyxCBc3KATELLpuJgNYaCitWvhC147kIr8H2
K1/0pJBshrU6BWOxY44LytTu0FrKHknwNAfsJhIjaTXWHD/ikJFh4RJdA5H5XNWu
oCEZE5rg3bx2cY8Yic0/jPSw8yc5LpbO3le+nI0FzgFZJOEUawDuY75Noo+Zcy3Z
kOCtzW5Whe4z3IG5deFcFaAG83zFrQ56xFwkdnyaZzN6VxQr3ZwbdbMneizijhB3
qFu9hHY86TKM3e7DFqm9tKtvVeblC1MrzDEtuaQyynSijSjWihuaKOMO3/O0zfp6
6YpFHRM9qIqGxl0DoIEzLKrPTpjNpanpKsaO11AkayLbVYRCw2r3VlntdwlefP1X
Nl/+xYw/JmIAd8bUGLPs+vZGluRJyAyv7/MgPSfQ40LvTs7vZg9zb4qf8MulOOOV
ODhzoZQq3DUSo05v0qsgEts2cIVFAJ8GOLtO8gIv570+uMZmVTfLdWQDOB1rA9pY
6DMp/QUugDdtu8oXltGo1XsyBqlIHCdKoh9YGuSsY8cgrvrAR0rf7jLc9jARa1GI
6JD0r40IE8wPiCrHIZnX802nqco8bpMBTybYFRKYBPCM+OPCThDeGYckq6M0WL1l
jsd06YKaTM16DPHXuchQObJaiC5nT0GhyV9iVSIR8Fz1qnOZg8vlIDp7BhS9OI+F
URIJiDluzIxR0VNMRh3J8x3T0KAR5bUQEqbeL7zlA2D5k6x5iVUih9RDhcKk0h5i
c7ATjhsSlAfwAMmex/Ql0KfNZ+0XvqS0ciWIVWqWhb1OLSac+0ecPV3LsPNW8j/S
ZhCvJghaFBchgkehVoGaGslK+d8LkvV3tJ8uxguHslCTWsMuyAAAeMhlhPSGoyGr
4gHmhFNI3QeNNQHWHp003tIztmDh4No0csau3t8DTMy8+IXgNihwf6Nl8jj5RRdM
Dq5X7EJwwQOdNb8SuEU1gO1Ch5uocIZrW+ckKZqE2a3e7BlAO58AbeOqs0cAjzQ9
HDEiMjaA8rpbcsLPq3o/bC2BfJn9InZRijeuKIw8TSFMXbEh/H02Ji0ZFZk3higU
jlMvLiQUjy9EJC0XytdDoNzo2/AJdxY+AWaPrR5s8b0Z5WGMBZqCWTwaCkP3nsBW
wE5xUMwkDIWbrvjXrPEeGXH5Mh+fy6XZps+kiUGEaXZwW1arcG8JoE8shIvQjZgR
Xlsc2o3ZpYlWfpO/iShbo26HzycP83enoVnZNHeHnljdISPj+fsQVjs8o/93y8pW
/tL/X1dhDuhDAuPa504hnm7AojPQT9hkwRSBNQj2c/fTVygXR9779/Dj8L0V52JW
qxh3MhO30jVwBCUcEAav9SokH+xilU196C3tTWSgIYr2o/YBSWa3sFxiSA1kfpcH
EDV4udB9HPd1DuoTFI1DD3YzZvkC8MDU9pmRs8AqsPvn0NacdGacZKlXuMaIKBxx
AEnLB8LwMj/RbZYRKI8RruhMGjozZTiV0TXAHzwCA/itqQywl4NJ2ySbN3mC9+jh
hkWX9thrqpv7trsRF1ECRWrz82Y0HzxlkvDTE0Bl4tTuPtz9mbdkJiWce/oqstcl
WIw/ITlWL93tL38SspTwA/HDv7aNEgii3rLIGFhb2/k05TbjVb3C4NQ4x5/ebSyw
ss5ovGjTnkgW7YfAbGztPirnbLeVdyDYdhOOtvzWPktWg6wlrK+GtLnuSFabSiKY
UyYbMKTxpeyxs3KoVIJVl1qptP+amrrhekBde2CkWg1VqWutiilO3FixDjXsKT4s
o4RdX/4hwTy3BKLtC/E/8KmBa+DbgczDx0npBTBWUvpVvLBdNkbkrrM293sMR/Z2
5gj8uyIkYhbBIfTYENsqoxHGII4tu75+6jEJpH8CxXSTocuKs8mslGBk1rsD8qCz
KJfS1PqbtE7X+NNDbofHFivHHB3FuGdSLabWsh9RNpzyOOmiRD9jaxEEpR/cDGze
EOrXa0/2IzdCt/zMBh4NVoSHXxA7TB6JtbvyIYk1Gj3mifPIM+qeCvdlgYY5OOZz
YDxyFBIrPlWaC2QsT9c868l6jteL7P6hIlOpGdGsGkgT4j+yBTyvLC27++XnXh+u
uUMwZNqdE80DgoIMQdacOhXHdTQ3XIxMuhLpV4LPPVLHBaVK6oczValQm6Yg8663
mcjGswirvRplNqOuSsR5WzLFlTPPgopqEncNFG3JQbsyxQkCwhr6/VRkJYXoHZpI
90O310C6NtpXND5kbk1g1v23QfeMgOV/vnf4o8arMMO/Bw0xq8ufv6wAQPWnCtBq
R8TIzh4jGeW8w8ML7pzXlM1z6UAouz0NnoBifa2EdD4HwLJUO90LiaQSBlj/VHVV
ZNpWGjj7dU+L4/AGdNnwciOs2tMfK7yEC76JyfgexP9cLBOhiIo1IC6kTe3zZvZ/
Tl1QNNqobgUZ1B/EpilO7AlXUR1hZoR85/YS/sFYASEURLbVWAW+oWjvMTqal9Zp
dAJ+Z4e8RemDqG/dYrgWwyaKWSibs8Em553Mst5FS0YMEu6TGoiEYyZ4VBzGxeoP
f+jreZqfB/venKjjT2YyMpIk4b5nRMJA0BTwo9TFFqBeZc8beEj9pkHuOYRITOgh
2cPtAfKY1/Ia/Yc+wXG7GjHG43WVnP/NyYVdTgtzL9Mw+oSv69ddPoZeZHnlpeXl
MJ0we5Oi2d4jrte+LMl1KAxmLFPeeejg9Kb2FeLV9Ipx13ABAhsUwOT0pp+MPnsh
OItnqSkRv+YjWukv9NqXpcp+Scy7rtcnnB+kd/b/zlmg1mNIi7Io8b9FN6NtQiIz
EgIK6kHVr7Giju0GRQyR8cSsj5c06U3gPiHa132iy74ytIb6nzip0R3T5CZZf2MJ
/5PneoTamOe9GILDMCEcJN0yk0sh79xqaHAjvd6CPSrI68aUq690+BN1+E9xOicu
D6tx80puYfraOodQLI+GYBpPoZ1Y8mEk0vhNp8E8+SKqpa57TjR816Axfqgr+yFt
iDkI8I92dLb6k7EmHVr/zDJkktJihXl1JZD6BO4XGQCTfPOCrWfd7Ea8YxVepC9c
6iQRZvqCt7OlunZ6/szTMPdHyIQxI9T0b1vM0A5NfPR6fCqPz875M3pjdJWnN3H5
oDBQ1/7Oa3ne8NQff/9ZsVuJLIk/0F3YN6YoHI/Bj5ZvhXzNkLDUqkhyWzUQ5klw
WOpSk7mtmFfzgoJCfEyWOvZhRhlHv1pS7TfxdhLMTFj00CoYclHx5RAAJt3PLW3W
WxAnkP8SOmEbPFKh1ggWkyNowtHEObk/tqRd1PPA+akw3OnrdWiySEMRpEKSt0rl
sJR6Cl83OZ1TSvwXGdjeS+o0qyWlXoaRkoxtNsAhhE9BvmrB33YnN/8kJgkoE7c1
qQC6ATWtvKCKAvanyfMb0ViMR5lNBGogRc1luAr9X54t3+IdrfJ7E6zEczydqKV6
7/7Cv7uTqlNbph9xRTXHHdKSqxMQs7/LxwL33A4qGF5dA8c90pL5jNS6x7GbqWxW
p3qTh02PVxZES3pl63oV6YWSG2UmrsSwHOfECAmJYVD+dBKkBYREJiOPSeI3VqUZ
3fzU8+2ZuBND8//9tqt6Y+/RRSxXxMCRcUNko4FMZ8ukU7ZoJ3jz+qvXwryttzui
641AFSJSD8OgmLLti/06jDaK3JP3e6b2mFPgM3ED0Zvl5TuCk0XEguKVhRsFH1Kb
bgH+qpgnKqP5Ca+mPtp7inEgDZgMZORF0cG1SztDvZ80cC6gZbbjjLmVVYTLmG2c
wbgvY0/lDrNANOLyQXEb4J4D+Uq8UaC2hTR8K1x4neY8Kov7zueCJETMZdLuj8P1
3yCTdKor2uXFuagt+M4B0nARtfRJ/uA8WYcuTIVjIgGvlihzUcnuNXPDrGG3Pt4T
PGCWk1ZnuaigC6cm/P9UrwpQxI9lxwcv0iq38uzjVlheXJH+BX3fy20lvrwvGCXx
XzE3mvLM6GFH7x7eXTmEviv3WgT2js45NN+zdAvOAqa0kZnLhwmB4B2byma7WLAV
JcS4Aergc2I8CU0/3SAbb9Jell7ryoKHlttQ43Qx/iodWBOLZiVY6JnKdCo+/vwg
OyWSKxF7uj3yCAP6Wf2F/NXuQxdniJhKGvJ5OTQ0i8VTDGo3PzMQTryCmz+bF71G
LrdezVHGwCcOinnWAtzAVpgNYPuxcY5RI2tNKfSjYSWUZi0nU8/6KyJJPVVAn/8K
7Ez0/xWARxZ9kVyMRV5I1luK5rFp71rPeH2JWBKrRjIwUDV8xDEOSpeMOIdwP3CJ
SEwGZeqDbJV5QsrAJMCQC1dtz574bJKO15vMUsF7z4R3GNYuBACQO85f7XnJZz4e
VqSUbQYxd3qJE5q0YiWXS7n6A8AreBpx8hZ6BNUijY84s114ulLEBIFamS71mpPd
qpABKtLMxNjXxSewXJGKLa1O8Gt6880qVs/IIgXbUiZuJ+scf0eljSuEWG55qAb9
F54VpC8AlSgGJCc4KDzSPDPdDevKfy03AwQ50Pw0K5ZUlBjhS/ZAwE5peXKekxyC
1YU1KCZ+OisAfmd4vRhcwU6Dx1Fthiqil1pSRcgIcRrSL2R2fPi6Ue/riXP/Rn4P
upYM4v5QGM2dic401bpe8LbUz3yBm01Umuv0bViwCWt9w6nxqSLoytaxuYmcS7Hi
cX5raCStixNeTTMQ2I9g7iA2QBpCUrJL1ELP6DDG2zK78Bu7F8mSQqpIFIkDvoGD
0cBPvXEL22uaFheSgLGqabHwJugUxa1Xe0N6RVSeIR8XyZjEiorPFn8GPUD9IGl1
xf909pEbON9KdAi6SXjfoZguC+lge+vhOU81z412QOtuSXtCnBYYnnvZlVhqDzvo
/iSk8d0PmqPHJzuOVJPedXvhLjQVFclMUNr9USYdS9R7F6bGSSKMxoFUA/0exK39
f68H3MZMxRWqJ+sk58HvXbJ82ONEyX9JOXaknKbpsgwLWBMlZhuBg2btMosZKUK7
PlglHtFLWiVFl1/irBCU9EhGvp+cDYDo6MOjE1O4oqgJTCM89jllpkaF7Txl+Ivo
xCtV2iMo1l4NVtnuypknExqsEqtLYMffxTfJYrPSFEzebsOx+leS7Azh5G4TX67j
fSLglvhN6ZGIEeTdAtzo+GAGL2oZ0f3R+5rMAuFWAKcJDPP4AkK3xl9Ab9icVvCq
qpmRv7c6RpaygAkJragBM8Hmo4DnFSHzMDT7+feJTcriVqMnCIK65r3ke9I3XE0s
ZozybpCnXvHnfeqPgophp1rhXtmCivwk+UelwSc8Sm3W7hZjE6NPgYOQ7U+cqVJ4
mPcPQRuSwV99PUBsIvEcDeTmK7uCKnU7rVwRc9iG03HOVA7vJoMVYxjydxvmiX8s
J7Cy76IsJeHE142Obopo02RNr4S5hpua2+HDgATQWQ3YJ+QHROVLKjPRvRbLwIDG
8mfqK+LbFFHIqU83KA6aqMC1ZQdTsTjQMvc3k871v1dB/m8OxKNFxRv0uCh8lwzB
/953I9H27xyf4A6N27+860A2g45tqlr7jcFWTZNJRx1vnKPd2WHEDAYOEady+7iD
8l5ngUTndDRCgm2ZsueLqlmX3ubq4oT/yKa4s1kqolq916o0E3N/XGA73js/gIiR
md73berV0mkWRXIntHr24U6zDbaHsHRxaqpFSb/hxajkxxP7bjUgV3yDHZ3maq//
PpSSqkKDy5iGDVE7qrm1sXNQC5sYvEXjq1//aL9ZsKezBaG3En7qbhcsHbiDRMEo
hA7S2L1cRv08fyS4SQ0xk4dgzG2ynFuefwSYcocKwqXsoRJjVT80T57j5cR+UUUe
pbihJLoI+lb4sEvaaYjq5zqggZK5TKL7t+3B290m/0j/4Wmpe//p7HYrPryU+3Za
GjMq4cHaywfgVH4O3B8AtE70xzPVE/6BhFksQOrFKjKyrFvj+P+w+u60qCv4gAp+
PCFYKgUxTObZzmMuGT3taJjTFUbyEMyH1E62oCvNjYh9AKbbSPV5eFZguhW4/1gI
/NPz/1bIekAVZWK3U5KJc8NRLHDukJZ/ywVCFp+7313ucfyycM190/nKc8j0/2Bd
02vDM3mx7fXO73u7UN3Y85ylLZkV0Qr9cgwEocSXJZ1ouHUCITIcY69K2KBXSu0j
HWPNZDhcTcYy0M4Z+NpSMoWNuuZZzkN6CjjPYzyf13E9i9z8JvNIipq0mp9e050J
/DYkH8hmGYqHr3y3e7Ovf5s3gXtWI5YkAMmQ8NSinJyw4NR3wwr5I3rAKTV4X+Cy
oLFRc9bQzmfPz061a6/3Vi+HCbokh5K2n1Ve9YQ4KZaLWNWsJo5qDipsTOImZCgN
gL/z7xtt3WschTmvAaW1QSAEP7BTI3XQ175IXqgvqrG6AycsVMvjvOSBWLxouEHJ
uBt05QRfdJnOBjKzQV/6kgVxfZ0US6OmA9BGRGp6TWH357MUSnCTEtAPpbeNpJsP
KrG2MOD52jVrDt91csypm1Nd2X1tcvH4gz9UschEPfGARbGnTZfpKwZR5KzpGU18
tLSJOuTpJOZ10PaWQqzKL7jgQ76GyknSYsNSx+U4aomQ6zi8ms7LuxtvqC6+6LVf
fgF2Y32t4d2LBVHwEACpwNUrBS989LPn12mWinZg14zcIkoq//Qo0B/eZyIaLTFj
uXuqBpr4oCpBazXZ9+o3mtfkT6hNWjF1E5aOcrXBlxrozUC8YgZaww6I5orV4dwh
LOnt5k9+IPX/ilObiGKLFSMwV/3Sx08y6nxzaN4MqLZGvfP6z+NtZHwggS0ZbWGK
kki5Jae6KSIUIXDskF/sX7L6oyPPnF4+k1oxRMZMZIq+97dUqIWo2SqulCfSPP32
C0fSh2o8KINepKFoGqzKMdvD0GdN2siotFiGnQ9fpdkPvK5lvbvO6CVdS62PF233
jSpNokewnEDslepUqozBTBSZlrCdafNRkewT92y98fDmn4PNJHkiPUkyhGzpQjbg
4den3ZkvDRzzIRo7CBD4ySrzMT4d6jyfEzFrlhKMEc8oX//8r/8AZnc8kjXsHE/x
sFyJSvXN3EOyBthyvQGSUZ/GxVrWgXo3ORtf3UuGIRoS4l/H1Hy6Q3lz5huJuRHM
GaTSJYLGJs9mjxN9x7O8bpqxELHfibf0FKplkwrrQjsIADU423x/tLPezTWUtlkM
Xs9JuojwhkWaFtgLprDB9dfgArDkK92H9WyHy3hlyWOXBiU3b5bS/h0I7TY3lID9
AazNstH8e+cdTWLqWUoEePeOTC06EQReYuxJPTywLzD5ziiXKp4CL9fl6wRjSh3Z
mF1ZgI1TeRZFB++9hYAhfz6/a7tD5V8U7fDcw6SCkBNUfuB27hbQZ45LhipaE298
/hFAtNJtVxPM7PsBRkNHpbkPYyMm10FtCufAE0L+GKmnXFeE3pM5x55JxJKdf3ZZ
XsROk+tajJqtuXR2FIN/GpJ9eo40UZqUijANaF1y5992vcagvJBvMeGtZQZ+A1OZ
6QcpDEYg8oIMU5aEgxChqhhBvfTMHOcxa/sIkjkeFKgmw7bisMn9lbp84rfid9dA
3JDD0WBCc5k6OE0NGs/JftbmnoCWlVdL/CF9XCNhAm/f81Y9XRsivu3XA9kYFCUH
jbUXiW1T1Vt567E9M4lT3DaB2bvh90Xnu65iLsRELP07mUWJ7YKoEOLg8vJS2bVL
3e1g0ErPEODYrlnBON8OvKgFlLM+lhw+AKiGQtYPAD+HgYd7b3ydl/q5HvyZwdCh
SXT7yfzBJY3uqZsKbvGcoosOQqQ/ZHV2UHqhOH5vwXS+jMes3jEnn2oOm+cpjGrp
7CJlwA/0MmySiK+LTgf4AT7PPEsNjAYcjOkXdMvIMm+sj38QaeHBLPjQXoZPtyKH
gpFZogp6kg33pVNTieNcYV/y/nm18tVf8ckaWdzZmPhE0F6Hq3nQB34k511vB9mM
rA+A6+1cwXPfGXsAeWwRSrznULOfw2w0xXGEuv4IUgtYywCSV7z8hh/ekgGSB2hT
YNevx1my8dd+0d5MjzQY4qwZVfcZzzRPk9Kj6PYDyY1Ru8PKsQfTgmTllYS1Be9w
k4d2HNe242Dk7A4SRKayqK0W2TaEXUV0JzvuVXztzgnXPBQAgU41KvR97I37RMBj
/RBQPblFAyiuQWi9PgO0cu5R720EQrvPQ8+mJX4zbAcHcf8P7SWI5plCnAcr4hBn
x/qSq+m6lWJ1hUTIhxjmGciq3y/gWI1jCBrxqH4ttI0D1kbjgtrPmuPi4aa6Dn8U
nKWWlW982CSmoISlSyNcIlL8AH/muEP59/5uHej95tbZcImCZoH8zJxmCJJ0NSBn
5MVdO5LDcNQrEHH79tlj+EVu5jsQiIl2YAEk7F2VlM7f78XEQgLR36ERZMqKggAG
a3kXCBj0r6zwtO4tqM1W//N6FERbFvYQd+wsVFS0LIHLqCWj2NAQVpesH53w1koI
aVkf+v6aijB39H5pEWLnphwC/tM7wQAN+UE3U7Xpy+82RzIzwK7z8uGVoUVuv2Te
t5w3jUqL05jkiIN8N7gXLYsFQEOf9lAFU7AU90GPkK2LojII9D3ZwmIPFqgCwtp/
5TjuG+MrkXDIWou7bhpoLWPZ/5ijig6pz4cDkBm90ZoG0fR01IJEuz5gSijeRtof
ukdttBpPzwDXAXN/ULhT0Ji51/qaPq0mKc4Kc+ZuX8akFUCluXxCyogO6SNi9vRS
ng4yhj/fDIoY0FCf1glLU6yeazJIL69qTCZX6Uf43LsrJbMAwBuNB6AaCBdOcnbD
3+RnSdyMmHY5guW0JEjt2trf3t1FGOiIkn4Hvjdtgh5DIkP3yYDXK3hHBGWP1S7Y
EYc0XMpE5GJ1LUIojNv6MC/QCW6AssEpk/AlaTx7ZxzxkmNM8wIgggT2fH2ktSW4
m1kEYpa7YTguDXSeNDQM82U0OZ8a24JadYT+VUtFLts1iesZsRjQLV1CEvH+fI4k
eoHJBvIgXlgwRIZG8wUQKnXedzX9RdJgafnbXa+8cV4bta29nyooSnLtYQ9+5O+i
uZyJPt+5GYA5LtDvIoXA183G02VqBSoYChgL0m9XHehvgXNGkV8Onw6mOK7c3v4N
bFpC8aeKRnS0gK51luzXExOl1xFtI0oiKWAM4FNW5E3e1JAGaIq3uDCrxOQ7YLlQ
T8Mp025nno2lFf5iCdAm44/52jcl9ECEjGCDsFY8zrDTjzXJE0QBXANWp+e9d5Jv
2o2chKhfxcbJbjaNQ7g0FSzWHEfxeGq3XwfTvR4wCcEfKC7cn3rHoM9zJwnub6LO
XInJiwx1GOdyfVUZci9QC5kC9a1/F4VrXRGXoaUg6JN13nN4t3lcSY+FhzD9LhEK
ncbeCHSR2l783K3pUL+Mk3DtoKTlYC8/Ppusx0LyNx35PmA+/6CeVVZRzj/SDJfS
ihwoN0L+St90hvUSTrDk1EVuH4pf9bgNk1ek8a/mTI1BtmB4VKsN8gfMbxU41esK
tkfgrFZNAmhKs6qlmuB8793aOvNsiXO8DbnfVG4VNEnuVxNI8BmS9eJL7XhCmT2y
maipLaAQeZg8cEM3e/OLHf+U6VjNmHT0cZTXzHm1c/JPmilj27klAMCr1Gm6mk3I
XqyeCLjqTrjSh8hdT4zrPhoX1v2Wq5+QGhzi8+zEt0AZ6gAGiQtUxIs8f/vorBj5
jrAnlyHvS+Jay/DehUeBzOPG7UQ1zLJ4MtdujJO15+kerrawq05fN1JGmgDn+pY5
p/hJguwvfqXZQLFft6bHRTt5CakLwR4HgFC5bBuEFs1GUMkDr1rD0vil4l1SSNzZ
xmniUaKFpjsHBwAGHP8QGtuW6gohutNZ32SAns3A+enXRqyzdxtap9lK51WEuoNU
790zPVLE+oLctaXBTLyEYQ+dRPCr4WlMaglnVN4UXEoBPdG54yzxRV0oH0kjjCLF
ytJXtbrtulSUWsG2sM/AWYA86g6EA6XoacVzZPI8uSOQ4ielYaWvSnXecVU7f8Qs
K176VdmczyZcTvibf1ttTRXHzS/l3vqhLJ874+CqCoSrz5mswslndln8jlb6c54j
/kD/oM+oVwgpXK5eqwi+/DkLhc8y9VVd/64l7KIuAVSTjhzht+G/4UwGMvDZW1Vm
/enApiDwrEzCJi4guz43bt3nVgaAiCM1ASwWguOneUNA6UScKgRdB1iROyv3Rs58
Fjg8Bo6SJvzbcCJlxPWNITeLUhv3is6MXXcVdEqjgQRjkrLnAb3lK2egme/PkUZf
gIiRnbYINT4R7hvMYJRNDbTZ7N3POtKFZh2RE1iOos7e96kQrIMXGjAExk7rifl0
0sRRpSqElt73cEbW4mdo5JtsUeFrRvsfFB83sFQV/5mG3IcjHt15mPUk2sPJ/T52
V0QePHNBn/9SoJbM4x3wosw1hCrM7K410HFP0cXUaWQt71ROmta2b7DLQRS9iWTZ
45kEjzRUbCkweC322SxtBNvLndfGyQfiUytHx9fhadUe4v1SppLjWUUEjwCJdUO3
BuM9gXu+3JwF40WFC+6Iz8nEQi1lV3LrQl57WgrjkVHwzKSQ79TrCxrw2JGIekJs
tIEOXDdt/2W446v0xg53MRPnBNcly5gZDx5CK6JOY6/x77WBTU0k6p2Mw9sR9x3+
AmgS74i7n1drHmRgYjL5Lgsj0VWquZ1b/q6pzJdsIRdrkCLhHVpAxnjdTwSkqXPt
pb4WXofsDKd0zzY7SY31JnSFcXBgQpJjrZFdpDZilYBszbTRiSykV9lhcMkzLVpR
V8joUii0mPadHC9aK4VDHDdbYC69NYpIJaQYepovf/LZjwJf+RJ59rhvkGToaVIg
eBtoZIzeKwECZFHWmE4fqLzK2FSlDYnzTENH/tSAAnpETDr25ift72LTSDvManEM
+pzXZq3AsfG6mZz/yWEOAwFvOyoKF/8740Tjsq1oW3Oqrp0BhJMzwtSvrEHj+nUb
3YcPbuE/q+sXjfjZA8phOG9MI03L8BJ760LLLR/Qygz53N2cw9YoGlq0sDIvA1Bo
2QDlIxET9eSXgARA3iJIHS5ge6J0P0gmjVo+0YpYcv0hsnQ5rknHRpWU7MBgP/nj
sMOq0VrqbNZBFX6wVSPYz8HoINEjb9X/BIXqe0sauaNYMNC/M/0WclSMgGYC8+aT
V5VjJPRbG/LUBEtoV3h09UBaus3LawWjksRw2FyyB7xgG8ONmaMVC3yG41hmQg4n
XViW4f2vQ229y6+8itnNK+h5YwobYQkqgCee4Ps+Yoa5VP8XYEbpAiPx1yaIZ/Cu
xJ4axmEQb825frIgYhYzCl5YrdswZ1VbQ8EUvx0cbej93EjnkGokaKmCxniaZ2Cr
RM6UQjUMzU2TbXfJ2+e07nFMIIzzM/eZ/SNo7EVBfMxRO7m2je/ZCWzmR3MjFcCE
uvN1ISOgJDdeVrGcdmAAURAQgd2AIUNpDTUa/U9TdJUTu3RxNXJiXBNQPFiHDljO
t8OVZMcfFnYrh03OlP2EHLdSitNwHYUF0wrViChANVE/RnLLSMz4RPQZgsEEfcne
UkVIoDsTsW0/X9ZJ1iWyvrjmFT9QETD6rewl8wZ2HROur/okITNDNthYgncXMjO0
WPqdjVQjr6rG15x6uDh/li5jLAMIy7HnRwhH/BBNYr1DUuqONwwV07Xw08x7ogBw
OF2kYN1ZiSYC9oduhxITwnt2T7S++1UCI4f7Nb1mZr97ag+fAMZXLkTuIx3bO1KR
yBFhqCqzZAxE0kbEs/8DodYxlRx3VqL9YYTtW6v2HJAhsS9sBdse2Kckn7Ve8Wvn
FLNFQO0FQ7LjmK5eTnyzzv3pN6QMzjRbdy9Hg/VtZVuXEWPp4orE6UlIj74/njkh
Nm/P1UZQAe3CffYVHqnMN+p+2H4WO6BzcIt96o/0uXo+/2M7eneQTqOllQPHblew
ybMEXC0jeAMVNQwSzliQbowdHkYvxxuqa+stvmnOrtpdNbwWi2pBtZkMK1Cpw0Zj
bhuaDGmKLgO5PZ1jDpA9kEQtf6/HWE0mthu5/vYvCHk/UUrDmyV0FqtnypVVHoq7
e8nv5uBlkLBKbW6plrC9QmcRKHfyXu1QRekWYs1MMphmr22QKNCPhKta6REFgP/r
yB5QF4k9ffidaFkh2RooXCpBSCnX6ullwHjZcSyYS3GTI5w+Rs3X2ApNmKOnc4BT
3TM4V8F/cr2Y/Zm64KCYmi48IHeZAFT8gRvlgHGBQldkeJmjtQF9tuCv6US+0vrg
WlJaJwsoHTg5CfoQhLrvDEuJyJRnV14u9kOwanbK6VH01Mo5uYqyOXnIo6JVwBe9
HXLtFkerhO++Ewij9/GlA3UufhhIjiDc50lU2SM+whzbjFm7AnUTZURrEpw2vXHW
6I4aOivtWhGIA4tXXWmPCQqNTvOz3/Nlq18xfyM40Sl2K2B1bkbVKmq7H05n741e
aFgIzTpFRQ+Hr01ApyXc70j8edN705LH6eRGirPJMwi6EfhOf/vPn/T5gr2iUuFv
XQTO0yzTR7ux40Nlfzi5+givB0pMpcJVGXLkk+g7g1UsLm06tplfiuiA6YF19nPx
9scZK40dSd9DDbhrRSS/bfQnZRLRGvF01s4J2AeeQp2sMLPtnLt1wt2bKXeAovFl
UOxBHdfaFK1Ea6BWgB+Ol3NKuB8u7ZG7ycPAyWhPC0tkaYtRqR9grc9/dBc0gvVp
z6yBnM+pzNqqTqEZuW2asWU0AGAmZJVRj7sh4wFshHUo5s03LB+YtHk8kVngR5UF
ezRGsGBUg1fglRErhd6CNIte8mDloI93hmtGeEyfHHU1v34E2lZ+E5e68hmIZHrM
qzrhTnwbcUyMWkl1gXbwlaN8E7edHR9y2mbD6ygYyWuhkS++gNh2+wQSt6Cb37gT
e+rdvrpw+qgPwyLUkJka8NPqwpDPv4RSdYucP8fhFbktduVX9DXDsz4azqR+qSCZ
/AoXA37GdHpYcL/Wwe82jDlkpNLzy0ZNhtiJYet/W+oeyctvEl63a8dbxUQRSqO6
hsfUeiAA40S0PsHPk72GzM0YnUmt0kgUpPkFRbsVCMOYGtVg1Peb8IqAJaPZgjIi
2ZYrmYxorBbKjl/8lCVXKkB6CoNuMGYuNVIjIj5mDW85ev56Lfq9QGJ9r3YUHWwj
UdS/0cb5GlZZDQvXjYLPobXMuOc3OEJcVIX+wac+ic4JSgnPeqxYVQXnP0TKUivc
Bjscse1uT0xhNaKWusiaHf0rXvkAGocQuAvKJTj4hl/1h7rxv55j1PAv/083/TVC
B+/8ot8JhJ3ZKgVGMxI8/idXyEEe8CpHdBOTt4R3/fRavW+Ws0pUiCHJ9z7EmisZ
AJkuhZuReX470JpUz+0h5ZNmXJi2vFRvWqGBlJFkN4kVUVd4U8K/qVO1HT8F0z1D
ZL26Ny3nY1RP+IYRZ/x15i8kD9LCSOJSuyRs2VgUJfOUpsOSIgOGidpUX2HxH9Tl
eyBRCKTapjRTBtN90vyDzmKRmaV4AwtZ78zPATdd4Y5SI01iRe70zqjVcUf1YTAq
tqF0PBnRkvyjs5aWRY96cLvMQ+OsfL+qpi+MIOwYR3/0POm0CZwIH4vRw1g3b8+7
WOVbfx6+xJDryOQ0+tbmMNWmhQrMdmI6hdyZXqpYrJXc4v5PMVuIPl4A4d2k4GRf
hR/uE9v8BZnJr43/8KyR4HyD4foLciwALg+LDy5U65Y8XW0v8epvJFxGeUFuPC7w
eK/004rUU7PscxazLfEmUpD/ZnofElIgvrpwMqZRL8BL24ZFVSMkIq3sWFg9muTY
Jj4ILxSk6h/IPmoEnuI2IN2nK6mYxOG6iRHIj7dgbQusayFCNa05Ym3HOVyKiVkx
/8zWqxEhhjD6ERicUQclNKF7gu/tk3OtK/elovirIB4djaNAxM7hf2CiF3WMTPaS
UNa2XO+p/Ng5dD4MrcoQxoCfJe2DDA59CjvsVZ10GsUtuTs3Uh81GJnGb1PgdtS6
hvod2eeJFh8kOx8zfMjmpxEHzhm7MRRvsr2dCduhirHDa+Dcvc2lhO5D2/V9Mp3c
xBOhThuJOK09CxPB79wkUJ0kOlYxI6lj+8hYbZ8PS6yzlg43R4hcUfjiibCwx5RB
LelAToutfZdoxtTUJOyGnk6hd3DkyRcwcs+t8cKeXvEVo7BtQwGCl1p+62a9n0oO
VEU348U2rXMoxsA7jWsX2SGq3m32u3pi3KthaJhOkVL8MW5bi6JPcM9tksga5pQO
s3qzwknQ4wOapV7MpU7ZV5xXOsCGEKoifLuRFEvbL2gKpzOK2ZY5vMEe0a1kn832
VJG4XDBLyYef2xo2DUnO3td5gJbNVyfBc+qj+iPSwB4X4MN4VtyBlSGt9Rm4qEAF
vwR78iDtM0LpK3onA63J5Xgk5m+XAH97Uo/8XDDGc5KyU2ntcN+pPc7MAXa7DF6I
wONn3UZR2bSFBKO9n6maWmm+vSDoXQ7YWCzU8RGvT/xTiKFqzt2b6KJhwDhv0pRK
Es3WyYt69DT2yLzPcvw9qSyxp+5Vfa6CYyf7f4WD6xPigK6e0YK/U25c6q3EwVeJ
42TgMGwSoOaBrYFrf1t+guDOXRlvRFRRcqI2TAeKHB/ekzZ0o4rwOjrfmp0XfZso
oqOp67+zZE3/eN+bEY/UHToLsyctlyurwWzsRkwRM5yW/6Q67wnBe39eYUPKT5qM
tnovwerT/SO0aZffSVRTKj6B+e5z/n+FEQ4Jc4MnhAXxlU0dIJgEOUHQ4t4cTuiX
Q9P2ZacedzrspGpVyuc25KfnEkexIbiqnQsAuCBttxCyWMEXO4PaIAZ2rwBjGkKk
mwPtpMJmcLRzhl09ikLsuRxigEbHowAGwWyaMHqlE9KgSOtB1rdLGLUHxXwww7Pu
Nw/zK/lNYJ6OgSofDnqNyEYS/R6gpvP92kxjb4pDr9i62dtgRvueGX03Lf6fc2lm
WAJwMy8aIyjY8HDjsR5oxv/1m/hWdQNrwDIqpMBd5rOSeLdDllWxsHclD5ds50EC
JSiNTstTFG68y8m4qxk1H0LzQZ8dr19A4/FwCztwOVpzIR/7NjrNc0W/UQed9m3C
N9sHivhIBGnCFOQaqpRv02My4KtLoglMqTeshz40UzhcYFzcQ/iAApHU5b7GRTYi
t/Ly3D3iLlHWhb3asGUztCozm1TBMMF/dv2VUZzzEukYNOxNyK7ZbYrWhowLb+Ly
XxMwM/Jf3MgXnyxOUMo5UMnyHzbpzPDv3F7/lX2SMTGs4iiG2UiQPChPBame8O/z
mJljSpRx1gqFuNt2SI6u0vdQ8DMSGtbMct8LD1heBh0Lo5DAP8BVMPrau02d5ymc
njv6VDutXenpYinhb/6FU2zxcuu+wFd7WeNoCC/Ts/Fed74cCNAzZIn31y34j8Kl
bBqoaG1qAG7FGeNTp6mRp9HGG7haxy4y3/V8t46hOCvYu6wk6NNbMREh2yjbpTJu
RwEtqMTYxZaiEwFMr9tbJiffs585xg6s4p5LeWFIY8yPiCq1+AwhAdTP8jJZvW4g
5a61EX7DliB2ju2KyGAZgKAUJQb6F3z2kOJGRmWM84OiGSCdItAmAaL5MAqBYZAG
MvY3eY7Q3EVgZTDx+40WKPlTJbfrSGD/Hl0fT1QpIZ7hoqXO2bKz2PvFrm6JTOKW
2Fc8MpHmVRyMQgmdP7ROUWDL0vefAjzFKzQoabRaPa2KS0JQuhsaMrm6hs2foRQh
1uFIaJgTiX/5qwFLM5j0PERTe1KvlEolpv2F3my27fFR0UCs4bbkK8RA4PNDmGKT
hzp2/P4jMPG15nUPpuSHax7+eGKKQ/o5Ek1w36vxVSqiz8HZohFi3iXszOi7kmcY
E4uNUcn8UdYWpbwZUQ4/yjTC5/76hxLGhjmYmk9UV8n0cEJOJoYt6JifcxbiG/Nh
JmsmG89OyaZIDXLChamvDqmH70ELdPYoHToiPQ0ORoUcuPHxXxka6DpRb6Vu6CD8
6eqaNl9O3kN42EbBImys+PbPjYJauqVaNGa4D8vCMhMBBseVFKGZKq1I6vTP5fd/
WFzvR09AAkS3/cG54neJBZi3kIHM0ZT4qBEPjcdXWhddz1G6L7MYzg0RIlDv5ZLc
BhYdRBBXk2rGDXgxLIU7dMHlEp9NpkYHsrCeBJBS8p1GUXfs+BDPLb7OgL92QpM6
pFy6tAsAXUt48HIYu0VERZlzWHWgxseFLYQj8eiUBgYb2XCqjpxQxfs30E5KmTdv
dNLX+9QhEmKKuNTxQ630Qy1usasKZzLTM0de0VFEdM7hXSu2vtzQ0U9g2tzFRvuA
I0lwKMlefhVb+cwOGBxP791K1eD/EzZp5hK2L9xsIvw8LV/iIilcQo1xPJzlpqfQ
3VjWodv8vj5KutFS5tOaft2cBdbHVz3ua1txQtKHjsXQ7jh1U3fQVbkONMck1mVC
pwW8PSgA6zSeAwcV+sgCgJ6hXeZOfrntTeXeESSpYXsBJyo4jnn3R9mxsesT9ZJp
sLyMahV6HwZ5h3MTsPhquO7GzPaz/6Z3DAcCHYytqCdA+tNyKzX98/bQaJkIEYwZ
9oVQopRkVnVNT0jpAosePRMsalHI7x0X6jn0K8Dq5Bot2KwsDfLFUW2AVunvNXxy
ggmYQCQ4wVFG7rnAUV1p6bs1+YsaSnyQHjq+ZmNgXxYkcuHDlOm9PYGnrvAhy2X8
yruS0381h4qBvdLpPmwGbClUelhRabjw55H6ddh4YQyBTlEslRDGIwYs807xc5jI
8Ftk3xmd3/HJWh8QDXUftNV2i4L6F+L4cRwDbhZCLpemfUKixiKZRS869d3Au54z
HpTYp61K7MYlIMzaKY83imb/v6VPyBjsAas3zRqOH8T71W8nl9ZwjP+J4hI+XeLn
+cCnfngx3I0U8fk0FmcZP4RDzvuL6zlBIrA1NCFDZncYKcdhl7DxpUwx8vbSSjwo
KmXFGtV2lhLQDKoBLEVQnFXcQdd4scNNx25jxjCjsrLdLsyCyANS6Njwp78orMY+
o0mlX8rMJhGuEoCBN8dQ+epCi5eOWSDafUDa4otQl9RgYU9w9b3Dlh1duSInkmsL
T6/fNLcu+fLnOz3RWNQD37mqrOuhxzpBLC8WNp/HyLhr9EIdVxfxA+e8NgDm3Un4
9KHxMfhRClVl2mGrJJlx2tMdFOGCc2WYJ+KemJ7ishVscVxKBgjY1LbyO5exi5RH
2dYGLRzJnWcdwR6DFdXDhoK7wstn+nt9Yrb3NCYXngSJfac2HcoxLk2b+S08JBmh
VFyr2xzYqCeTyKjzQA7/stV2Ff78CoquRPHzVxWOcTqkONNrzHqtlfZthqBQe/rz
a49QHvsO2puzgZPamV+fH5GPcBrl9UCsu+Ma9y85znpGK2EpXycKDJZnvOOobGOA
orre0kAoNnqrIh68OY4apWX+betbZB+MWQwBBkf6fVxqTRlEtn0rwlN1upJs16qp
lgbdWSnQKqfbJfRi5R8PCWu2jmFvDTjyA+BXg7l+GnFzT29G+IW+m7SRthc3BEPP
6LPfHTKYsPz80M5P6IYSbugg3Qs5b/SOtFba/Eet16+kKth2RkNv4P64Es8+T1nl
iD83LWFWazmcLzIIy4SgTrXVloH+5ZevlNQgBoXyngBPMMLCdO4BGS31vxmCF13I
2zeO7DdKeydcxipoXHR3xsICDwReRfLtgHhe/uaaZtinKQMenk0u/CmRzMwMgS4w
vIkiU+H0hb4Z9f5uejDkotPgHI91THX5hJYnkxjRhTtg694WyqvpCeslbCtyssHE
1KrQOeEff+UECC6V3O7eXdVZMbY5Rz6Ufi9RcE6hIjyQ76oIda0x0FbXuFVfX2T1
57nps4NYblB1NKo60Ex4KN/yvE2Y1pFN8JwZPPrjDVBqvJrSdrNKvzoLjs7kPIc3
Lo1vfC34ZSozWCq+JBfC8j752LuKN7QUdyuUcU/YTCzq+aJOnkXm0+DtNhBEsflB
ey3H0LV4uG3zvpfO0fB03clPTv2E7I6smd1BqJZE2W9UzVsjww6dwqcrXUuefyyM
QJF79ea6roaTjqm2uxwvg65aOGKujF1ZvyHneB9LOlVWdHum8xrb0qSWcJ81sta5
r9WlyJeBibFgU3x/E6ATiHjsCxQHrsxcIj6c3wtBpu/LZmwIkoPSSVQYQDXEWzgl
jSK1AcsTNZfdrRaYov9ASodMsp4KapxoQgdNmeH1+8T6T9X/jV+0ApMDIsVnDXYf
Lamjar+sg9/8Wytvy7dGGDssGhCjutliZm9db8pMUjC1zv71cwuY8Uqul6dX484E
3O+gMNmlYSaxWgquEUc1HP44fmrcTbs1mz5WB6hbSF0FdAYfgsvvCTAKnFv1usqa
RzSFPC8QcXzLmtTPqzqF1Mn+eD0rqwLJ2ZULb1ZyL4hKTNdeXa8CpZ4JgDu4x3Q+
EsQj1ihwSgJerQM2cRRWUZk8R/ekBVTj53/o/8dtzNhuLj8xZKJ7a3JhJFQZqVWp
IhnApgeMTRbd65xeXAxcKGdslPyKEL5POLYXkH9kghmh34L3bZg2OYA42fTtnsih
cj0VkamctyLJPDnEGSEg+a2+aqm9Vx+jZ0rToKM7oGy8ZcXHJGXzcv1pGS/wKptl
7ctAbpBD4pPmnKjoqMtE7KW6rPbnD5NNJH/+wvitfp4nK4Kz6hxV/LQBqShH2EPs
NTlyRl0XOTecw3u/X9VffRZ5lFSXreMkabH1ifNlE9UoCwBqH/uCOL4Hw1nI+vk+
DAZM775RGmz9e7iJuTYqrM/EC2rxj+Qsvfw0GMRP7YqsQe8wL/OeIIh8Em2s9H2E
8idZIjBlhtEa3O5XV/ok7COX161U4RTW/94Hy7q6uYVG/DE0guf2/uEriifJ8dvt
x1owwXKgWnud2svcWNGzwIJWxXd4sKaK0Cn5nFs97eXyBvs/dhtcDOhVRjyd6tni
X980WvP1Dxo3ldf4YK65cc7YCMbmZEw2tC2wQPEvGOaFDcWeLSMR+2atmdKev7+z
Nk5LfWeXc9iK392SM+0oIurnKIQSBJRdLgXIIHJH8oY3b4VFVAe6B7hVQN0FtpRn
b03MlB7X58de8j5fbxjnpcfEamQaiCiNETtNXe/+1OR2DR4dpj72sS6mOagLj7tX
feYK0ZSAEKuNKWtYkmUaCJbfKO+DwGrxoBSXFessgZJFLkm/ffEC4DJ7d/D/aaEx
WnYoylSLlyvItRqkhRKdBvawTudHPX3pEThbX9lOeqwn4F07p1ZAL0TiGAR3tIfq
8osEMioY7dkyYd0QL1BVtNDPh2Ws1hD6FiptFS8iTTpjgF0WQcPuMCULMS/EhiKf
UYXyLaIDPeZYpsgamVMWCXY41rp5AtShevYyh4EDtMSAk9SUxes0F7EUkuyLPS10
f+WPWuoS3TIRs1W0UzCzfD+OHLIcbKlGbuXV2zyqDo1JXi/QI6p70Aq6uM983nSQ
hlQ7WyTnemJkdo5o9Zes63xgQjTDYhiUejx14bTxJeM+m52RH1uNPUowMVa7W1nJ
TCW50VvtAwFTQq2pM8oaFDUINKGeJ3cAR+a/gAOMfS4BZ2QjOIS2x1AxF2Kg9AF+
030E/dWHHupVedKqGuMts5nHDb6vC0rDFGzSo5A9P653HjeByuBa7BUfGg+p/btW
qb1r20hTfctLgHB8ZeLsT4e/MbZT+CxKxuXnbo4YNb6A7wtOGXU5TCY51UuMNVrg
+CBiIUK7LPKPaL0pg03AVb5CMbDS/hN35ZX83ueCzsfNQxu1mPELlkWFiaK4heHN
kRlONCQ4l2rgVNysW6wlvR/z9RhEPphOGbFVK9dL+6jCiHtiOIboXyIHUPY+LX9c
tW7jvo9286utfuQ38osK25mzi4XqMBbwlZmyqi2Tcl+K+NOGZ8JQpt6ekRX2wrAT
yUPvA/IUkT71Xig/TxW7HiksjghwPBAIfkEuoQVma92a3B+TYy9vp9j82YC+mMFW
fBqf+lRxQCLlHM0SHo82ory0IZ+anNTLy94zsQ+aftPzyc+33kE+QU0cwOb3OWZT
VGebsHCTO5XQycp6d9dzGueIu9UYEQz+1HSmULmH92bLAMI7vi+QB6Do0lMbEkP4
3N6K78qClsxNODiY3O0vSlGQQEBhFSmNtaCu9ziZnw8TBHQkEgAQ4uou/GaYUjwn
U9zWIpNKdbHdbwkLtizASWoIbT4F8bliL7IFYYSqTd3zxup6b0A2IW7G4q4QijG2
12qD4okFlmITDD88izgLsrfyiCE7w0Yg+SABP5gDeLSws/4LFlZ6lez+4Bh9qotL
790p4a8bU2CrnqlENO+oSu4u13nSQt1/TsyO0SE/3EoBleQfewuJ1XHdVFrfVqgj
035FyoOn4m4UDoWmASkvmoWF8sLKzQuTEZwMnlSPC5a7Dw6+0KZErdWisTYAHb2D
QuFQkuBhmjq9hHkGYUvy1Me4DFDPAvvpJPlNBIcGePDJEyMwMqAa4zNHbi/ykPTD
K7CqvjgMyBKw64WMiUZhTYzAx0TvTQhmfx37gnqu6/o4nRHacDWFV34osQd7Fg8y
o/VkH+ZwmPhcNFx8wvSIIT7gtPYxxOrzznhsKdEiL2oNKHEWRi4K7CUEK/GFPFKZ
Ak/vVkx2ODETViDpnJsHQhGJRU/3VMP7eR4KnnJCX5XoEUmjDEZMQQzB6V6EMbmf
BmsLXLNpGNJ7Uhbd2uOjSVyoqMnjc5bdsQGCiyruw+2MrDtk3aeTcpzgeiIduaMH
1bP+lHzgvfKTWrTVcCpxwCAiA0/0ZSMVemWk0Km4Ua+J5DvHQtQ1tlfgLJ6d3JAG
IpmT34kHIKaX4T5pLFPCcgCrtBDh3zeE3IysjahktkAlPV5DTRzlc2/IP3zIxrqL
qPMtBkuLByF1aZXc946mjZUyPaYgM9l83OUVe6NZHvUUIi59ACeG38s284+hzEeq
RtMmXBKPTMGDX5o8FyxWcmegSgzNZAkAcPClRPDydHtuaXqKHtcjlYbzps1a5JnB
foHjN9opseNLtK/+mkEPAGxY/bqvLg+FwG2ug/PXNxjhDLy+9XGNHcu7JUqPJHaF
nZk7U/bxfU8sNQw7ViA8GEgMwgbUAYOOy4uoRkKiVKzNjch6NmwojRhoYBJVMCZV
mx6F0zkKv0f6GhHt1fggxNBitvouMgoLLBcX/vfU5L+P3EG6ALKtgf+8skHmNUb4
GdogNubGDKvmENgNSuCJFFnEmk/q2V0dreDVrwtspPF3y6CYvvnehpPtjiGL0ROH
rNKEAXTkZ/w5A6Rp6CK0btp+zVZkqlvpzX1FkVeUv4PF1+W2Xz5JigmwKQunoYBJ
SRKgtGk5aejOAAxY9Cal5iQyIbTolY0kVN9U8VlzV7su/dUc4eHMouCQdcnxD60c
/kgqRAEVc3LJmGHpzPIf4vtZBUUQeqOHlLqJo8lEiQu1h1YGDCjK6rG4cP4erNKM
Kij6rnTjALbM8kpHPsMa6VBa93skk51kIgklxIe++3DODArClUimwcHjcCix/N5N
IsyXrGDbkBabmVgpefI2Nkf3VH5B5soLMw1n95qVJAioZuUr0tekDhRcM3hmtU2F
r5x6UUQZl8nAa0r0pYho1U0TTEqiyLyqeAJJS0eEIZZwi9gzadn0hKiRczx3gSHZ
isdrf5sTMnOBKIFS/ZYJhWdre+MHIZ0NRIuRxgvufHP9b6mRSE6ah2wojuw9sO5P
lm5lwKDWWaJPIaptPB65+2Gy16SZgCIVW2CtbjOiunSJ/j/FW6cIkV8WWZgcBLqE
WF1uWCODDs+2Kqf774dg9HG1nR6pE/fHoWjnqWmmEoysKEvsjul5m/jyAUehSTK1
u6GHcfzpu7gJ/caYZQbhv5svPZPUE6fHpE/jGGxHvaY0FWdYc7aOKibvVl5j2eJO
YRKJIFO1bl+lNXO6vx1WhgjIxVJYWv/QGcxlMQNH95rOY9HAzTrQisDjVnRY8sPg
BlDsj4LLQ9X8wUE6RkL1LFYrWKOj0H/fZnXcY0edkTMtVlM1tBjdYwhIEIvgY2iE
7k0g3b1DQvIbX2oteorSEmoNpaD/f3nqVtrrIJKgHhOVLNJAaPpYve1lIExftviw
z03eYL5HMFIbsDqpvpc6+xfdWpliI16UKN3jeel1Mtr3h29FH/lfW0gxcrKoCm3c
bIMwZl7FRJqoX1jo5NCvaG/d8S21yUMMA3uhZjS0u9bxPtGiRm0+Pv+dCuMSvY3I
2vGOvHGQNDXkoNphEphUqlHBywnQEgzD+Z/anRjO8qCvw9nSGmkGGt+fxWeL4fOj
lGnsxwFhzZ52y1Dleu2kaKMDffIztJh9jbHCMiolxlE9crcbbN/jigHeKrTAWIVo
YJ6ObT/Q8Sm9/ZjXNqV81F0rTNwOmSSDo8yRo93XQiVQZtMsF+Ml249piEL5BAMG
TS0scPuOU3eLm9K+q8GSEh/uKWEhbYjBZYH7TSPXp0sNjqZRRJGxuvghJ7aKxB+d
JjVBgGIoB/uPotUD/Ws9XdE+dlqzQPeQ925OgyuAibOfmxY6n7xzUSpKoVFa/zG6
pMNzkdYMqDih84yOo+7k2dce2v/nud+n6Y5xGoVR0MzfwvT1uSM/Nxm3qYvWDUcc
fHxvvTStJgEdI1pe0Vl0sEgeaUb4H2ZWwtFK9PNkT1JbaW6x5PxC/Jaywvyg68pP
YjnoCYnETFW/WolP8rvSOUiQTOkf08AcljN2+//wnPIaP5ryTpTeGSkV8w/ielVQ
9js9vt6f0EGZ2vFlbGNPqNivOgWFuuDXfZfHx9xSvKTwDFEGHsuuifLOLrGPzkK9
8jnA/KYqhxy/EfI/KMyWcf60rYGchgnICC/6mrOZaaDbyjPmX4kTS3TvGJeKQGpO
tzQpS3qKNJlO3unkAZnxUHVKdaqku/ZouhmSIsccIgOlrYfXRh4LGWHqfiefx9Eb
lJ+qcNaNhqiQqRKvnNkj2GLvCdiZBdcckhfKIYJAaEDUWTgUVEWaUfW+64YbxDyC
pi+7JP66tjUqEvwwJimJqlZSlPjvyADzAQ7QmFVCaPuqcBnXakk/9AqLcHXo4ZJb
IG2+tFWZ/YKco/iat1m+60XAYCmrKCm4byVh/k23w+yVI7T8S3iWHNQf1xu1FdF4
MUSh0dbVt8MN2kNVCCUQOnGnhcoRLCXVHFDUnOWWFLDlnPBLWrDFtp5FVFEYOawh
a8rW/3iWVAaglLExL73ZUQwJ8CHyeaPjA+OogfmWy1s14ixpn98b/u/4duj/lN9O
lD/EiN1yHFvzW4WEFNSEs6gfkmushSJFWkwoQYs855agZqNKV0oIaXfDeu2zqXUV
D23dG6crFkRZSc1uD3a1QbL4BaJQadYoaTbUzmNugxQRmWRMW2cLWWDkU6Ym/kYi
y1vRpy+2lnZBfxfVUpD7W1Sv5ga63e41Weu78dX4MgcsNczv2mCa43XG9EuudYr0
lwoUl8mbxLax3ZMusWEbiBiGnnt4hHQjLhl63Vo5lWqV+7SSDTqtu4nje+mnaXut
T+lEoeru5fb+Lwz7zj97f+Q47P/520FnrNUMcmTpyEJcFm4g5S5+kUQYOdG8Goq3
cG/eH0H2wFmVdh1Q+Ea9wcBuBTBZuh4Dq7jJiZV+TE6qsxXcBpt2uMeF7YVhbjwS
PbriCuiip+8jJmerRrtsJ5CC9eNmSxncW4dnoNRNdTYv7el886a0SrjWczowUsuz
ohqCRKL78XQ3TFIuAB1kk90HELPpi/2+Ad9W2ErHEMNeuX7fc8UU41no/Q/ILPNH
WvUyxAQNFW4uEJ9oAxpR2WULk8HFNESrd/qUAZGVcJvJP7TiBhintrEwgnhQ9fti
kqoaxo1vLOf4z3LfprXdkIQXH0Tn+lXySfU8PoHrPo3f5ebPxQGIXUQZLY6ptEN8
WpQbG49QP2klgPyTID39I21zgairFrdrJOi2KffRP31B/0GD5LTSkxSbtkaFu4+I
Lk2Z9WOrcePvJF6961Q/hUR6MVFWcc6rlC7jzQ44vAta7qwvxbzMJzL4cY5Ec9zp
7dc/bBCRjDi9IXj3WqHnGnzjN6BL80sPJ2sPFVy9Rrc1nd4Y+c22sQf5MZ5qPpsc
FYz61/rkYlh/lWFkpDZ5/jH3EoGhi4Om4BVcLo2YGAWgfYuzqeo+ZpR0I7A2Fik5
D2Q1ohkAbvzVGzI9nY2HFwn3MI+APUoFLhvjLCSkihfYQDT3v8k/egppeJoOlQIN
aDkpn6Zqi6T4TJCm4chQtbU66V6S//BMukqWfLpfIqot4ODWdw/67DmlWUnZ1ivE
7PEDKoN909gWgStjEWt+2ag6ORuMHi7k+AINgelGvCDhX1Rq1GJjaJPXjFVpNK9h
sG62SKgYmV9Kh9M7kP3U1n8mE9quM54+FQqmckgh5Hk34pMhnUkrNGJbqSi2QwOO
uYiOXFSY0JQmtVjQ67eDCQkXyKw/vcZLPQpogbgZU5ArJKW3g9xdhj8ww7OIjZiW
G4g7EByvQRWgERfc4tb7TwFfkbBqncyxABwT9hHYpdJnikoFKhJzJeR+TspMF5VN
pC518FG6xAH8nKleHLtzs4LZI4U9BSCjr0j2u3TouYnpXOXC722HCZf/X0H6REZh
N+/OV3/axb42TI/rsd5kKvenRxI0OxArcxSwK1sJUnPVRceHIwgUb1vTgweNXYR+
nh7sVZcgFA5FY0ZWMuBmx+eNrjPnkiJt4B8FfT+RWRqRcu7Jzw3PXR1EPFjBw6BR
//tyAIX/5+j0ChF3Ar1io//Wu5zo1hhtiO2MMwh7bLncoarxhgkkZ80MEw4VC0SJ
pzZ0mS8kZy/8PMFClIvsWIAq7EasD0G3+F2+r1rU4fjET+vVLZx6BcH0QerZxRIL
8dhp0ws+QAHgyWoUn1pb0gmMRycYOBngXJpdMTLhAWYKAGUNL5rySV/RWHaL+qzu
Bvf6YcDQOpVQYsA5HKgUz9lrPNn7kXwdHlKEEwEE6ZClpz91uKoU0leD/ObyDm8+
WK15U6WKVh0seHmD6fak+4nKOp3mrW189B71DrmeVAQ0uXTnFCZ0FztBb5miJ3Ot
meScN0u4qodf0bXsHngMOzsVP/AYf2FBEOWN+59fzYIoSD6rOcRbASOYlATxhT9m
f3GcAMOzn9bfuGHTxwRbYLWKqNWk32YxAdAXFtMPi7feU/IGKNq49z66jn7NGfsH
OCjnEMNDAXF3vFDmqyEvb3pbCTc4XoOUl2ybSa1F/9EV0FOx2AIi2inmxu63qoVK
3i/kgvMamXQ5CLpOkSMn0urebS73WXlKYUMZ195nMaRun95R3c/fM7quR0ME32vT
JAYQD3R0XYBf/jhxeoCXMARB4h/FpOWPFOeNysSV60g/mbojb6MOLeHhTO2Xsk8Y
N1XCw1e8rdqxm0lPLCybB4cIaJ9NPowTZmDn284BLxz/5z1RFzEQWhpk5c0GCFAu
B2hLSFssJoa2W4W8FXshVHnf6HRX9uMogYP+hvSsb8h80f3OP92hsdkauKZm6KYd
X/nHe6RTeu+4rlSM4b1XtSGCtqQeOV7dV5nVdrCBtVCIhC+4eOVjoi63HcP+FjvZ
vNkws8I1gYUsFPDB+/QnGhDSO+dOums//IJPpZmthUQvqV7ro4y/0vaAFxqSs9+S
hxFtYnyy6M4EgVUohCbIbCD9Uzw+QdpHdrnun2+xDD19BYIUKavy2+yZc8afZNad
FFWVl/kfeqoYSHTZkLMDtCUFmWiZQ4z9zfocbHXhPAMW7hMFelLJF+db3riPzDDg
mUBdTD8q8Bn+ZL9QofdTJscQl0b/Bxw758Xc24tGh366PT4TOSUUeeWZvD7hAXBw
P6fbvInT40tZo+k9lW8FZXIi7NCGsnZ49jUWFAKEwgMmAsjW/FffsM4tg+RnTKxR
rS4YpkZkL5BADXdJo35sWLPO3LGyltPF7m73OM8wZy36ZNmxj+di0o/+mfEgrfd8
oNSOrcdK0puTxPXR7BDHKJrAJZqckScLpSC1j1gJui/Cxo7hHHdC0HZN2Y9Cxyge
JoCdklgeH+/kHgsv87v2gippw3Vlc7vaUnGR4KF7KFdj6DOaF/R4vHtAgWtshWx+
k5yjgWv6zBQ2Qb1L5FLMmJmMGWzsAh9QaBnBjs29j5Jzb76pWMGom46R7lyAQXef
W+oFEyEtQZvAwRun+tiEn6b/1RS21J0DVAH95VvK+fP/Z6E3ujh6/0QkFEZ0mISJ
xzIGPq5Oy13gTYUI50TeK9ArQGn2YzIZp9j69T5AEyZabB7JTScv2vleV6aweKCp
I2GS/vvipWI12mbaOwyGfGXqplJbvo1A602ftDwkwStFNKBy7m8xunCv8HDbEOj5
cVbXNETv+4x64RhxDEuIy3PwtY5K50ZnywNUs2KxBIADTy5UuXn0/PjEvAJM7psF
FBZobpJiYg+hPLaNO/5DjSYcpaHuH+V2j8fVH/yU1eDU5v9BuH+EDeC/SzVTZ6mA
kJb4+6WrVGQwBethRqIC5xUaOUjJJvPRBXJozyz+YciTNcE2t6E8YZIjE0YylxN7
OUkYC+onXq9QSrIrbdJLf/tAgbOfbHL8ph7i/uTyjTkxLN0ls5CA7tLQulW4SjEg
BWBRSKguT/X9VY7dsZJlWQnyFft1IWj6Upddt4dOJTq8mpMzXhUL/Fy0B0TD/eP8
qBbm3Nh2XADwwY5J1jWDOUNwRjxxB5jaRre26zDS9g10QUNad/YnhojIiqdJRZT4
S+nXuBiavfjydcS8oL0GFte05TiBMO9QUsTOvE9awKFw3Rcz5sorYlMNO6aA5JNe
Dvsj1yUC4F2CWTfgntaYxbJ90FaAXqUNdykzFe3YP9/owfoT9wpgQtzcywU8+BJY
obqrOrrOAaOv3an1g6s+XsxEIvy9VQx2vjl2bESXicCfA93jZGCysw3S0UYnAfFJ
infXe/OTlUe76wRX0ceC6hLwMjmIOvf9wvI8b01wdsxjTXNwLOxcdfjqCXVqYuXt
nxxG6FWPHHPCn5KW3AodMdItT+102dvXWCHvIMHnHjEBqEsJSZFD8GBuyZh0cO7O
iGYWy64sQZFtkkCdECunQibWOk08vuDWNQhV3MUyXBWDagze8ZcgFaXI+GBmlygA
4ywlt6Pr+I+QWUNB32E7UFTk6IUy8RNCMzmyvUJzpjp03kfweePLCPD4rF1bwccQ
w/MNuxHgsWzY+CQg+G97CFbNKiPFJM5wfZHwyRZ9S6atjZvnMPne9o2TLKZKSdfa
zDrzDzk4gqJ4bvY9LB27XhvSdcc5K5YKKNiPRw24Vq96e01ClonDaEayoAG21X21
egGyrtjf4DArnRLfUb21NzdnWMEH6M4WFx4NxYaN51Q5fURmgmD0cakpEM2bjZNf
rt3eGpl+4UW2X66PqCxZaC9MnxyCsNTnNlpIC+Pc7h0q0WAxyWxPEYZh/Kq8FePX
7vsvqs0KXG0eQ8gBs+952Lu33zcqBPY6U9A8yakocS5m3aUde3ZS2x5ZaP2+Fps9
ndRtg3KUhkvUhBiwwgCa8pODU9kym0FqJT7Riru6IkTZspdkiefukqgBu2mi9Dde
3SEfJMFHspiEc/0gvseUugsQo4TqJTClzdBTGEpyGjGztj1IxBCcBndeIQh1mXb2
eXZb3z/lIp+LvIiWCn2RAoicHbrfkE+x+WLecRaDMg7XAQjq/Hy5v4RbggAMe9h4
SW1c8gn70CSmVkD7jjUxM54aIQY7AzmhVm5NPGr7+XIIu6b0DDSWkMgpPAsIgulO
k3O3DIQDN98/VPAdLPiJMIeISOkCIOhF1c1eIkTqQZuaW7Oc+PNLsRA0dX21989+
KvYz3ZkBChGVJ1KXpYvFfa9rVcSYa5ruC1yvDsuIYisu7LE06e+VPlCN8BXAE5vC
X7FmfyckezsCQY2jzTb3aySa+LpvHe5iqOaBHDTq/qc6B3QrjFmbZqKpLTNce8cx
UUGnxhjsXtmkd1Uo+jmRISzvqKsPSF1xT1ZCW1iBCCT3YQf9OAVlvbP+QdxwYldA
wAKtqBeL+xxOJ+9D/B23PMMZf4N8KdX+yIUJwFGtYuTA0l5dny9Ll189Oe4zMHQv
yj+t+23VFKtMO7c26mnqseEyPBARaQ5sM34AM1s8tpGLPoVQj9pC0BzAO1lsFk7a
UhGubcsLUPYgD0kxvdlKRqS+z/TBF/obhQ8dYCLqqsFOdN3SmvkLtufPDdizaUOH
6Qo6WwXDjqDfGHlIg0w9qrqEQTwDNshCLzEjKdLUfiJjIeCd6FIlhr5C/YZr6ej4
Y7Oo6DG6WQX1ldOG7VI29TW40KSYlvohlIv8Fyj5fLZk19eTYVZkXkAlD2g5iQ8U
mL2HiUDYaO4UkTfwXy1FlBZJ53FLRmKulBxk4lcCcv1R7Z8TJ3ukjrH+bzcT7/XT
1oik4xSXajFPNivfN0NONmmDPZ5kNDm4SjCPtdVoAftY+JnABwt2iVT3n8fV9FD9
VqZeut1kPiXAge7gxvcsW5qJp5FYrXvj62ITfHiPpmSf1U1vVuL7Q0+z9izir7Sf
pWwk4/3xwGQ54iYU7wDZABFWKUN777J+q1FUJonIxk+PC4dL71gdTG6AsHVZlfmP
Og1KfLAj7FogbTdiTKy0tYz2HwjUwJ6ZwO3U04KScFiqOkgbXfuItZEK8uDnkgw3
oBQsagjE47hOtHLvuuAJoYPenP5MErUSXkOMV1ZxRi3Tyh35ie5Vfmx6PVP5boJJ
6P1PWD7OYdkWSsXC98AGOIK4qITmT6iR4SBJ3G+aptA3rI4ytaB910WpRCT714FY
WN6SbUcpRUUJYRtdx2XH43Tq7SzveQT8DD2OdiH74jPWmJA5X+jJbsTA78QDJeOS
ZJQHSeTEC2A3A2io8Zm0Ga8QWwG1XC4hGETa78NIPMW+vdC2Bmms2SC0RbzEoliO
yt3zc8Jjg82nZtK8wXbNwAUwsnuXYJA4O1/pU4fI+jxXCERjBxa6EhGUuI2nHTPm
PvI1NyA2HvC7BDrm6I3Bin93VUEbcxyiSrI+UuX8YWDOloXA7twW774OB+Bj/yMa
huaZiPiyzFpOp62e5VCLXOvk0RdwWpp98ftwxny6nWGpsZ6GTwQUZtqQ5S2LN0tU
Qt8V9O+I2ku0N0umxqt9xWTtX/sVPiZSKYDiebD7dLEhSucBshj5nPCTG/PKDjYC
xlFvRUvsT0NSrYQ43Ntz/I0sAD8yBz0OiOkqHhuWXiBu1yHSnCewjPtq+ktCWhek
DeYxG7Yqd5jz1azf466CGtn1hewmvTVt8SsQT7d6T8LBaQs+3AdYFnyRP/hd9q0h
0kASdmb7n2c0pHkJExDUU9bulaprBc5CvCLs8TV85nACQvgzwyHnZiUG1cdYgmVO
4ge1Nuwc8hkgqXG/CSSRS1DzEN85uwmCG8LSh99816TFU7GRZ7xJUT5MgqgvS4Ap
tiDpQl5QBpvv4gjhTLlJzq8Y91Llf5Y/SKSWHRIWYr1tsCOAdDACYO+Yfj+e77ih
eb9Nm+tUSQSagSydvUJZpGCo9JSeH/Yk5qBU3P6IC1gXcw8ypAVs0IBsWkW0vydN
eiyoCJunFc02SPTL8GoNcK+VXIH49as872H7VLsRCg0TggTZFSgrwm/2cqs36IEt
8sfcLO47C0zFGhDRkm7L1T9CQi3j6WE3jHHazIE2Hw9/e/0gs8t5+HQUQbgVWn1v
lE2dJ+J2WvozKrwl4VYcNsLFnegtRuGkUrycUdXh88mng2yj8mHJHCghmg5S7RRX
i8cTrbeEwcP7Ppvs6SQuVMAy6g2E89QYwXDUzGmYLvz7dnN/8a5ZXdTDsb64Rohs
LtoKqrPbeE/EtejRo9bTHuCxWd/hR54DLuupr80XWqt5KKxzPMDHrERNgxvgq+3j
Szyv+qRNJ8KH7BwLPvkHjRENjdcZwLtuee9u/BBJm2BsMCiR8tlkfx0qlZ5YV1J7
0+PGrccntmHb5OPooYI3plO+y1WRsO9Ho5c38EwA9qWbV6SP340BngXc52RgKtAz
syQTIIIyu8o5gcOssnkaUEVMIelLW9bzNPfIe7x2nDngZKTv8zLaqkcyTGhEoGty
0F46u7mZ2ib0bRAGNn42S9K9rBUaYLpRxnIvHyQd0DRzICjKSN9tsaLW3CcI7fkY
wcilyZ1ejm1EfiYxd+rvsjpix7mfZhuH2/9pMHOIAx1RcGlrEWloQHt3aD7NqIAe
RiC2X1m+n8qitf7PZgrGJyKQbyOMGxjAWB0QStcqFe9AaBetmEEJxHSTgxWNKtJV
anlHGHE8uluvHRUfTvoSHVpkvHxo1wMZSSUZgcb4UQ9zLmpWAvHPrhFZIDLit2GN
TeBAWSe10JerSv0+63fE/5kThIrG4PsBx+KOSnA07IlMtOWXVJo+hy/jrgU8y7Ix
crhXOkiH22CXlJCOSkNyHzU49b8dANu1ryP9+fZ+EHg9hg8zfm7t0dObtB6GNI5s
qQe/4skxfGl69Qt7Szrbj5YFGs0U02F9VXEo+13WQND9BGxVW19kUBMu8m8RRwRF
9h+UC0rfpvrlKHiGRlL4Pob53sbV4RT4Bktb7q9piQzgS46lwz5Y8xlzygBkUSCe
/qiRVNqEB6sA/GTH+qO1LZdXgum1TY1tDUcbUSIeGTEeIwdIvTHFbAXPBpJPsdDv
W7Bv/H3brqXDiT/sLTDnwcNHW3FHY33PFpOgFUcdl6EyMPjAKNCtRbg9uSecrwKK
N6U4giTSPbx9jSd8I2d24Kf0FooIRh+WjNXcVAXecieA9PD5Cd3f4oVB2WO2/zkM
Z4rquUmzemCtMt/x9VvqEFH+zg5/5G/LiWwu/GEse67YLCDw5bbL7/N0mXHKTJGA
L/5WhzWa3Jtg6jDLPAJm5lHthvoUb4yW/bfh8p1smDnJHiQOOdzgkhV8xpvYyqBn
IJWjQVFf6kUad6FqjaUxgjgAb2JZxtZJ6GsRnb7ioQck+q0phKcjNM29IVR/McZ+
PcsAW1rufGD47smkeekzLFnTkn85309JFPiVXlY1aulhx+ldEikZ8HEGH11Is29z
DrbkpNQXWs6gwFdFy3cbGVxXYCe+AbqmxZX8MlcqSM2GyDDGiYdbkMstFqeAIeX3
GkSSio/beAimlnFcY2DIfOvMAtbue/aJppOMcbDd/6qpfG3sjxuHto45R2Bf25yx
v+F7LZPuaJznxXtKvmoX+tGfFZmidp10tRvh21m8MnEGGHkoEWhrTUcB5JmvwPa7
5S85VBwUCNjq27SNOemYef9RVNUfL5EF9KglDTqn6pmqDthXtjEXL+qRszZR6x93
IPzPtP3YX9p+002t4vW9mlBFy9lQcQW0HWp36zKOMZtXuRa+Xs/TOiLWuf9BzNm6
It5a7Qs31J6IHunW+dx8Vs1iAaKJOBSgcTXiPZ/bsWX+3O7MyJE7D+Rc4UpecmcR
HWIrIKuNEQ0GBHw7nzdC/ova7JEtZxF2OV4EwdD2drDEZVokNj5Eivb3EE8UhYBl
LcykBHVZPD6wcSUTWEMUgngQl+VvaF80xjRwaTPdT3GltwMcdKf+MCh382Kub9Hx
UzgvMdHDw/WNmJ/N6QhHa6PVVelkqVFBru5nf3uR5OVH9PeAGdYdTQlHql18UY8s
+LEgFMBe+vngvM4RQjUzl2cXMNuOxBUyKaUq/9O15EzoKNf+F7vRQ2wLY07XxIsU
HciatTJ80iw6rYOkbSE5D05VdP2eIt8J8Tg1QhpQmcuA6wUUe51CVd6jbFLJkpZD
dUHV/kuKoZxSHX+bY7t8zFe+nEmBgZ4/dFKto8cBv5ypzYrmJVAzaeUeZHlWT9jd
s0QFYnGMpQvd3hMPeRq1p+rEF4B5OGfB0aRpqkVu9wGhzVHBW4lksgysEZc8E0cS
psEquwZRgRLN119HpDWCk+PwTFFMFjGTgN6WqUe77wmlTW6M8WT/ud1x7u+D2X9S
VLQE+XD3SSYQOOP5ByACceuNvAVsf01E+66TqCrDRSjU/ebPXsluiw8KbrCAOrwq
ZVlYTYcQkWUHJ0LkrXlsFWxzf0KBZmU03fFI9uZJZfGvkC38N4+4+nrvAzlgIIbx
DuhQhuZrg7yCLG6Y2f1uaJQk97QW+2Eo0kjGV+oMSzM0P7jfF5xP5Vi2kBE8m062
uMORqvE+vvbifsa1yB6+gDYNuNKt+YV07RhvcSbqzVhCTU9D0TsG6O8S/oHbWZlN
THADS8K3Cyh64MlAZQNI2MZl+KEim+uibSNd5cuzJ0FZdiNvDM8Fr0j9XfeU6MWu
lzB8ho5tMNWEW3LE4TpsJLTjw77Qy2ojEZxdAgxvoquMNA1rZqI8PgmCRwMt+yEd
F6Rhoke/S+vZEI5jNVbSATrAa2MS0UCuevo5CtlFdXg9ASRzb8CUiKuXA6059rM+
Zb6shYcbQRvck5mihV51hRgXTKkA4V4fYYfCG9TaA0LcsJ3+n55G+wQCkWD/gj2o
AMPDQEgxXh5H7l27Xy2R8m257BcmIEp0eTjBCngfmXL7z3dVH9w7f5ZA67XeUYz8
c5T0VPd/qY2bOYXI8BwWlX2tTXy/+QYu1MV4apLLDhT+FVQKYZCdzwFt3aGC2koh
IzvWPgzRaw7lFxMqGk5rN8Az+/sokXiZJNwWMzHK/PtO4sBBxmbJdETL3mRroal2
j4JecbvCUwf7lsIaZpSMnWaZqdBO1i5Q3WCpkvlvGwMZMvzxDndICfkBhRPg2HcB
Xmvdml+FFOEed8UZKY1/KBmQhQp8SXkiRWGERvAChRYnlC69mmpGzlkcB9kY/KqZ
1ezUdylyyv77lnuULRD6JynuQSX8GMRjK/X9ND+IxCENV9W5rqrSFP0Y3pmq01YS
JfZ+IwCUdgdX1sI3uaRa2jmQ2Fmw4qMHrdE88O+JjAhzl/9YcaQ7qG0mxlbabfYn
GBCl0WwWkiiTn7+seEPDtrP8eenE17cfvOCECZwRYs6X23NcFHMdoJ3j3QBnl+WY
fPrF5HffIQkBI3y819h1yxI8MqueUlkMfuEXm8MkKIMGpRa4+dE7LjrKrrYoWped
8XpFVzODUL65YWia/Zsn7IIbjLVqzUN7EpqsEj6fd1z4+EXZ4SpH1k2I8UW7EoRV
NdsZoumT5tJOmyfVOwjpDBjz+1tYIUUZaYsFUV1aqbnphm3JvDEoi34ScA0o7J+Y
4S5zxYNv5ZacNE0JU2k3bnMWSMuRTm1kQ3WLmOeu0+2zceI7MU/l88cm5ptDbNCT
dhc++aZEpF/FCj3BOH8YdmxAepfTu8mrffbXglm7DIxmvehRZqpmhglZ4C+TxWZz
ubD/ITVrYx1dPh1OG138t/PNUyeC45unofCP4biDj+tWIBMWmqcfq7E1TIacZ3Ug
uqMM+fLXBIMXAapjnsz0XuPbWNI6ngAW12j6vV5wn7qDt0vNXf5/P/PzZKYkoUBq
lQSPak13k1+7WYoj+5r1ZnfstRB2j6kFMixa9b2o20czw/pZ0EbD6HPgSU2Lt/Lj
9yaKf3wIfTh9YpIw1UqbNgY1ucZHQPDTet+TbZDiXYsTCvOFMlHbD3Rw8iwo/oZb
7vJE3DGV2rBCyggM/+u532dZHju9WW5ZSZYJWm6cxNZE1asq+utFz19MT9kwVihe
hHuqcFlHKDuO3HHW5rdjzGK3Fzz78N/neaC6ABwxbh8MkeDOSv2VroS31qMcYc+h
aHzqi5o20fzkp3cxlcGgABFgB7dzpZKZZloYiOfoVSyoap3+ojGZeQ60uy19xrsh
Kg6TWcNt1k4COVqQiM55N51Y1ffnWh3bgE8nWDL++XQYHeI9p2OzPndhQaJSS9vJ
uv9prHCBFJcidFgLu4TVSQbCF3ErbmAMZ5REXCJIQsv/Tbj44v/Sf2bHOfSe7Xvq
rCBDUOq0V/3Jv7x9+aK5hCnANnpj9sb7j3EuP+EZm0hIvDk574Y7KQFfohrUWsaT
iGyxa1gK4EK4U3HHQk1l9B3uvkUgu+orQ3F9U3aconViNM+4KMoR1lAJwPqfUcXv
FZYawh4+hz9qskfmlhoiAwqGzsoZ2Y281qcGlydlxeizD8jmSUDeFXEW1nf8TNAQ
VC/Q//0xu2DjnoyIXR+5/s2oD2j538fZY+gShFDAU9Q/pP9ZlQ7wXKl3TqdiHizb
clrDhleeDv/jVMk0pkI9A6HHSG7zThNXqb0j2SGTw00yPMbGQczDC/ja4klnXDv1
z+9+YrKDGLpBbUKZr61fFZCl2dVZdm+hTToh1mrJlVeNuj3+Cq9/nK0fB8jcACIw
X1P3aVSGZFKu1pI9Gdkiq5iYPRtRsj6zyN2kVnxn6AxP98A0qTSPnxfP7hqPn2Iw
19vL+uOMU/y9FYvFeFhov11cnuW1XstY2Z1cKdRrDt5s+0eiwUM4heBeob9M7fKF
sFFl0Iifv4RMzuGChZFhB8G2bLEU8VDECmsuNp3lz3u5E/byT79kWMQ9rjyaY6rL
Gdfnws+4o3Ko+CuOg698ymTZbExu33wzrFPWIAvOAXdgXZumeZkk102Qqp5OkqBh
OdFTjcblcQjRFVtXvWNN7tZx95rHPyf8ESzebUFFG6Obhl+mV+0zxIZTcRUe9BUP
Kx5hvq2zhIycMUOEYGUEtXkmiaw+OvuFAlt+px/fhlh7UV6Kbsbwd+Cvrwlh2pKJ
+g+KXgB9LDlUn26Gy44DUmTlOXGN/ltYbHSX8OA7Wp9bCA+snj+ukWoXx+VGf8iE
yAsROCCXXYm+5rRVA9U0KdSX6jey8Rti56Xoht64cpazOOMrb5p8yh5jIb6dMh4m
xNISGm4WjeAeNh4QjyaFFhJrIiSw+qINQzwVhSTgjzRHdRsWpPdd3AcOzbrVm6iC
QOJQK+TnqC+XO4PXidOm7YZw9R7Z89uUZfKMNy79J0etTEHoZXMQWG2PirqzJA+P
1IMGki7obWKd1+NXMQ8aeGrECwykDh/e1OWkzt26sSHSv8AbYd1SxNG9qAaoa1o8
nhzE6sVBM+BT3I/Xhdw7SrI4YyHjQIlFd3m2rMiSyzjhEh8EKaCIOAnl8FffhWbo
yFTsgrqpUiQJhlLIC6Kychrw6kOBnpuCa+XDZxCxTR8hugUUTAMWb+V3PTMMrvdQ
WwcFasVKB/80/Gbtk95ljAaPeSQrqx/GNO9D2Z2LnMrLG4EW+AoJXGrhQFHcqgi+
uXg6nzk2MoV7+7hWyjLb6WV35gtO6jgjswNO8CBo8uk00AxNhCLM4F+TdhXOxjZ8
z01a0MBxDiuqYc7pRZ6GdfD7hguvCIfGcVSG8n6ujQ13FLCNBN5NPj1DqWPxI6Kk
7dHXmMSWEDNq4KNuc9bYL95t9OixgPZrOkIFPnstWsGAo/JcExS59VVYZfpz1P9z
CJ+QZLEy824LXSjgYD7qkZ1rxBWjcMxh76Azgb8mQJcp5SyWlEGfW6v5SR0IuGKr
Exyyqy+6Qgjnh5Iv4zhs66GY19yC/TC/rNzGL5UzuaCoYclRbyi5Rk8+q9cVNZJi
rpmHZTcmujgajN4UqQZ2mUAoxnZgElL/06gcyhkqc7X3TQVFo/D1YVr/9DVPBeUl
pNFY50CiUsB+pqCMnNur2uERGDP5CJz+a0m9YRWWu3q9FJpNI7Ojy0e2I/d00ZBH
sCvhUlVi07RE5DQVsy+Wg8IZqFDvSBOsTnVMlpAzKkCc2ix1MtXWyYDdpfX95rRm
nHaY77DRBnpUw98DPL2Ip0xJRToRTfA0SDhegXNJ00/KF1llZrv8O5XOxkD2TxTT
P2iPdH2r/MaCyN5XiA6Uuh/WRN1fippBijU3kKNrT47o9UXv2ONey5aNyQuCwFm8
Pf/QEXz2sFOxs6HG/6ehfthFgh1ZDWaMFmDfx2BUJz24vmCsVwztN64WvDQGNhit
o2iMA+xaFIIlZPzbJ+CZ/xN6H0cQTExymyuSF1E2+89lSkeoZ6tNPbKISKDU/f+M
KndleobJNqOv6owDYzaoQ34rmX317iuCtBJwF6vUpLF8zXR6IZQEE1AsXLFWTxsU
gCqEtP/gcdei14XFHB0CpNSsSatgoa0bVUluJw/UufHfJ4kgrXO8DmpVBx3SEcTC
Rn1ZL3V1pdWSm/cwYdBLhIQiFCa9nJPRyA5rURjcI8uFXUxpdOstuZDfdhn2n/O6
W4g4w1zVEKeo+aOVNNJo2pgcCLEluc6MU16KK4Uv9o18q0Ocr0X0Njv92rNw48Jf
tGTOidjdjU1tlvh3yjP7s9wjUOLXDBQV1E9MTGT54b0758wkUOvQR/62Ohb1uohf
75PIRvP7Ace37G9057rXllUYqpT6SqCkmcxREKLbb+cRZJ9fDWinZWg65Mn0W2d7
Ofm2MwTS59yq3q1Vk4TCPstKEZC/DBmRwPNtG9NR8NXanh7/w7qzV8nP0YuVRBs0
PuNU5d2IjTsAD6OZXviiOKSmedRE5N0AeGWLUISzJ5L9Zn4l7GYZCFqyBO/ii37t
JFLv6ZOi9HO1O2YBlsAd55GVXCKU32nRg5IWJ3qUm82TRI8TW+qRD6BCQ90xoD9k
cP+nhPtIkMZOvOOEegSWTNX/JytCg11zqf48cyqwZee4CLfdBwvk8wuGh9ZSf7kh
fihgQjlAZTBcXiCW7TkiNe9Sjt7MOmaxoXyAUaNDvvFwkfkHiwyb4jO4/FHM3xHN
Kiacp/8Gz4kqQxD9Nc5axNoz3Ki5wpbRcKFbrsPdlulpShlItDPjs8zzHcaE8AAs
oWKwU85PlSRcepDTmRnUvBQ2locNusl0Dwn758B2i83cbR9+cI7Kx7r7jjlLpCgx
y+HYJuFikBPjXHiirQoH+W5ByeZRvMFIuHbhl7sKXISUVQ9uSvLNpFpIAwicw5Et
ym1wOTol9y29wKkGZkMAGgEyWbIex5Uc/QeOpcULwXL6IuAvysv9zWVIMhKF4adh
BoQFY9+4pWm7c1QQL/nhp8/FfQpteQdJ5N6x/Ugwg2nEVogwBpzonIY+8IlFQtDA
fh0RjxTzNe+y//pukls7VwiwYrGwUH+xqdQUEy9/rmIkxWRU4nDWOWmNhgXEE7ad
n0C4/yrQlzenIUgAHztiU+wXw/RrduAg7NzqRRxAgE85/KQznVPG5A5T+m/lS62H
7qKb0qQ9CxpnM8X+ZtOqTFvgH5LHtmBd1+w4Z+Pn0pD7xOmTlO269fDHJE65nl+f
zz2vJ2W4cBPUMNwqCzjDTQeYQE2Fplsg9JNKfFIaPcsORKbAUeGZzpILQ1eRGm68
8th9MyFNDzF0OTb7In88gI5WEOCDaz7qCCNeLjMCDDfkpZc1xUmGpe7KcEXABzGx
5M2pIS+FSBwhSujQowZZsjY0h2oPTJiRGWeKQrOKviDrKIepQADtVrshq4/IJv2a
wKk7hYN+elyCB4x3x2FbVTHNJXz7YcIYVO+mSZFMQjZ8dOw/35iYhGOPvIUqVSdZ
bcWnEvRqDs59eVHJHoc2GZA9FUUAFPwKBCLIlEciSLrvlbPMjjAA3vuJ+1A0ILux
1eqdQEuLH5w7X6dj0WOc6DNRVPKj0c1lxhInVSd/CYY13c4yqFDApVCqkW5zomX4
GayNF2Kkxeig0tRqDlOUezow+aLNXsz82aJeYmgqDlhD6uFGMf4dHpO8I54VByw0
25Pjd9hJwf+hA9bc7boJI1tZ0HDRNiwye/ggXdiWw7nShCncrMLgJ44y5u0GNEfj
vJ5YOWUFYKeP7WmjQYjoiC9miKl+hTmLFgpS02IHK5HxQ83std3q3YPddVGTgteZ
Ynx53+7GqwxsxGtsu1bW3brSZoF7Lb0N7d74umwk4GhOwYnhjfKMO3OIt9pD6AOc
TeRxp5mRXZpB8zM+XCLNRzaXPpMlBTO6etK530TUst4knrvqsjTsKYfrS1B/Di/O
B7aOfYmIlzwn27IfL7c2IXSSoDr12KTLz/bDj60zA27E9fUfcwuExStsuMC4uTa2
YHPui1iG3NDLR3ontgkFPsoGES+CaMB+yrgdTkyytqjYEuRTXDGnm0Qyn/PHymIT
fXpb/eJUhREBF/OIltjYSJO+YfyQZKdX7vNspeXnwsMGpTob+h5zEpAKRRJRKJe6
wI7ue9Mj8ABn4XnrYFZRgXHVWHwnSTmkz4VMhhHKnn+8J1upXccJM/6qfjdgo3WK
swnd11Q1EsQnpk9HTsKT+fmJV3PUstpOg33GotO7hiBKSQHqHPZGZTuOuSod0jhp
319nqsi0kgLMP0L0RtXttBcU5uchlsaeV7A9Fel/jRufjH2CbHvY1CC4NGPm3Byn
4mnbLD06yxFTV5tURah6TFbvKHHbN6HX7NSkV/VJkWLnNQryMBmowp4d+NsLkQgN
WPWWlnmzYLYbEJR4YxoOuu4GP4Q24GzNNrxMiAz0GhNOASPD+KG1MLvk16cwoEbX
N9EvQc5/d1RUg0U7TdrlS3Ed0zl4YzUaWNn4sICa3H4EM1IZvm7RHx4tCn9C4ytd
XA29oMCTFXiZF5EgOPdU1bPH6optyWkxZrmgw1m44XNIZyM38wnLA+TLQtXWEMsB
xrHmx/q0U5zqH+iui8V2rntrmMlmtjI/fxfza9ghhT7BENXm1q7Or0V+ROTlTQFi
yOW0k71UZvPFRMW2pg6+K3dHe6x+2Ke0Kvn9IKZotxeiSQFzsedUUJpN8Z+VZCLW
GRMEFXDMy3z4JaVDzLCP4czXi4WlVBnv1blNystuj6QRtnt/leBvvJoM0QFN7+4w
924O48tFplH4V+JzL9IEcskUDfm7Qe6tmvIRHwtRGSQlUB5vk5YBeBNxh5Z2u/Kc
wH+/MtcAIfD3TmtF0Tj17mArmFpkNREuOazthNJstC4Y+vhCHP04lRkSZ2A1Baib
s9d6OHTKZhiqDBW/Mv9LD4Xy3MRKwa1DIO4md5U4+AE2FtKEy3Jl1+0OjRL6vWLX
DlHGrVl7DK8/B2frH/9g9uxUrUnBbvgAIhSXocIWsGW7+Cf/M5ekzkT8r0dyTkhD
ye3UdRY+HGsNqZSdLCyPxVRLcM2mi6ylWpYcYuq8y3lEYAaBIZVwo2I89Dney0Fe
b2n+rcUsz2XNt3L2sXe8dYCFqaHl2g6Rp2LYiU59bTV45Re2f7UnL3mOpoDiWDYD
ykeolztZ4NSOZS7wtJGK8NSPf/ohwU3W+zEeum5PClpjzejw92ovxpiKcwq5qNxk
Iaypm2Xa/qYRaCQlxC35JOdjmP7Th/z4SEA9KING+fG5ArpjZSkjNXfR/Y2/7Vxc
SM8YCKr46QGQNXRftj/hYM9Upqk3CsduncS+wCvwFr+v7bvJaNXLdp/JeoW4s2R5
5gGiE6JZQz9vcOmqYnJPo0JDBXuHrQVxN9p+BGcaSukwPYS7XAYsC8NtgD6Aat5z
VfoE1YN1Ch3EVkMRNSpdg8u2xkWRFqHgu5eO7C25vrw8HOfFBowHKWwZ3t7BMQKC
6XwhRp2N+/nHQ2jU36eKJGBgmZYkwQS0ttKS9J8PNEFA6ETT9iDBMEYqvwYwPzZ/
ZxywzYc0CqePE+EK07Q1HNcinSBjpvtu80WDiNZ4YSeGqQeztvjVdgrE++0O8l7a
lnmWgxFbhkczcJOCN5MUKVOEdvkLyYUZ7MFetQ8LiDMQnDxKUgiQYK3TyMk6xi2i
V2ZuNK/UGXAktln84D9fr4zuc85HHW7oWCx60mXMcT39DffCh5UTayn1WpgwmNu6
Rfb2nb2toZTNLYm0W7nM9iaiA+NvR9tAo9oLwp3pXU7W04a7eD63/lRsDj0Hf1a+
K80Azi+bNvFLM93GqBte14X4J9nE3ayUwewfqNpAV4lGcDbz6Hy18jNNCu+nKc1j
hhlKQUNsKDzLYbIwnF4V3dKJ+5G8rAEwl2Bs9fGJVzT9iov5V+OIhcfI+4c+rnnR
4aX0ktEiBDICxfIc5lD6vFkJ1Eu0y2Kb9Nbl+3BoVE9/DKPvj0kKPGb5GXEtksb0
wVh3tQGx2rPuo5pHZFNM5RoUUOkOPpDmPBAqDCyJ6nUbB5+ANJsdBjEG9zJ7N5j0
2QKhYOxbiFgZGV5Ta2VPBHpw3fiCmR0qmDfwfVe0DYDJXkw7WDVbe8R0lTMOgPtt
cjgjcw6TJK//PQIZA8awgzYLuvwPVivoP0L5gphVDHODi4Bc7fGuh/ueHdp8O0Yw
1JUIC7BELpsG20JNhS+/DgeAL8xHGBP0Jgwdn4sbNi/zLYW1Tfzf1+GBxvC1fqxZ
QidEcFmG8rz43HBu7WZy4gH7TWlG+EKSBy47fQMgCBSb+KlLBavRCxskLgNVZq5r
wBHMaZBQpDLyDz8cbL7/RDM3zVkCXCklmJeefDw6ueZwOcftGGQpnXZpEaHpfEjl
gZffWByxg1beG8hJ5eVsVY5frc2Eas7qMIN7lzf0dhMq5NqFh65zXQGFtpeMFi5z
NWJ0zAg6gjEeNJmGxbkzhI1C/bEhQVNMG8wRuFYVkpCZN7Wdw3vEXZlyu5IlMUja
xI1Vv6mYK/VhAVAJEiI4//dresfcVbrsCxAioeMmFTdwWlKwsboPa5g/ttKM1EMN
YARmOmHcL/fHuo3SSCWwQoEdzubxV7n5IZPvy2Pl4ZSCEn2uT0DWcZwZUGMNRUFb
ZY8QcgdtZUjJb0TYg4CATCa+GDm/Q5jJ+DTOBvjjAKCw+sm2hGOz5lHicq173dSV
13l0Q25GlLH8BijcEjSeVldP8MyqXnITwyi8wng2FeiaWwCARau30ddqRnGgHJcF
sZZkxN4nvLXt4MFbBWdDBIYwUsPIimmK8mQ+rD5foOgqUY2neAKkEictu4xUssbW
wzuO/W+ofDGBRWckgF+w1VfMpegsQvUTFvbuoXUqlhT+5o7B5Vgl+0hPXjQOeuWO
3i/8UPM/e1kDXxFrOWY5KJI0P0gOKcxlc/titWlodQP8I20C5yb8pz2ueKVEvACb
ZTzAZwDOGZgcLO+mgZdPxI4PwOpwOlYOKWqbVqs14Q3ZKplqyEknLebfXgU9VVSC
VQYuva0gZo2zqIV1dhFqvDkRfi0BCx212gE41XOw/o5QN7LDxUHZ7GNOF9fNqjcy
MYMrHEndKKQnBtst22jZ7B878YDt6q+NJ3QIYMU3I0Us6KWlttpihzeJL/x/PkGo
I8CiD8RJ75B2o++Az8Qbo8/s5WIjX/XYw8WFquU+apXxkAtZwhyha/QjrQFFnwKk
fzrpN29b3G30ZLNpUKpqzh6Fc+UKWjsv8JFaXYo3Sre/ONGjU7MR0RElATe30m0M
Kj++mfprsvydin6y7HMqaohGWK8wdr9ope+zVDCHiU7G3euXQf/a4Z5jaBdLJb0K
rzYLzXtoYEH4aBxwsmTnc1XDCFZhMdoBAYCENUbUVC513nPg5hC1coDI6wF/yHLE
il5D4jIXxxQvgDjCBIgkp78qwd8h923J28OuU0G+shSmaAhrva8LzukHE/06aILQ
TSCKpg5a7/Axjw/90dmMqZJQl9uNkAyJOWNY0uQYcLkF3ReEBB7R6t6cFDz4jPqB
8Pqdt5+qMIfwliLA4eg7CSHFkOZI6EKipmMjztL9v7kRtl9Es8ntzu2E3mhzQPio
8wRDqqzZw5EGB5u7U95j64A+y5z9l68wGVhkPuDVWpIofF8psJsk2QgLx9PHPANQ
2rot6F6GhP2GB2Vvma09+zfRQYvq0J/JrSoWSuAtnrJrJBVLwEtk3hWHjY8WNQHO
6n6GDGSFcw188e90Gd6UwCrWdbhAQ3UDsf/W6ctsyEAeSp/Q1Togvhdyz5PcZ+px
KGrTBSk6DtNbeK0Rd9hyFOz7Hm5uIY6TmJRxqa93KotGPLSDKN3xHekbLT+NjNLh
kWwVVsPT5hLykCWMIqAce+qzPXgt4RzCf9xHnQT4PyI5MFhnqlP0oh/1aheAGpoA
Gex3pg9OL+MDREIqOOZ5vssMdNRiON7OPLuaoFaE4ZQbqDW3/SLsBq2ZC53XbRnN
kAeZ8h3VZBAw0P/KCT6bBXItY0Qow2zP7m1qINodm9qnGnYYfXkKDkscU1nBBxmW
J+p0o+K22KrqAK1kEbSQ1NtL6A8dt82qA5XD+JRR+hGlb1pT85DPgYb2kBDVkgWG
VbMSCt6mtkVZRSkE/N6lHq0pva0DwQi/o498T7jimAuiocbEOEjfHifVxWBTdS+P
o5pzsWNZPhOKE3D6NEyzjUPcooNwIxJBCSwRVBkNz0oqWw8uXoJ14irapzl6tcOv
GdrV3N2Dy0E8ip3EymRJKK6ZMB3OrauTF2sJvu/wV1Ay1Wc7Zt9uJ+EtqhCNV4O2
JCOcN6pq9AkDW0QMoDvi8XNEAM49+zMRkubEGI0NFzGiskp7hwr9d3MAW4AnTurN
j8DaKj7+lzpzIqf5rdc65bhZXs2Jj7oli3l96qzLNorkWtE6O3VklcBfRouf73ds
zrNlAsox4lrdKR09DD+n7vmuk5WFMUZFHP7agJK6dJ+p9Ev3BMA/yMan3R4AiD9t
0N/BH5Barwoh/rGRaJTw8jQfWv7WCukCbcr6X71N6oAqQBRwWAsPsyQHpNkX8paE
uUXFTzHQc+5d8F3nYP/T5o5sThO0yt0e+LLLeM9Ami+NY8MRaN12J1kyLQDYxV20
Hts8MQN4wuMjWT2facYgqUCmLr7umxm3a1PQtOyNIqT7tOXqw1i1yWQ6TpNJEEU+
izb1xKU5aG4b8t+Jt9s6jlNqdZGBDTn2sMSvNNq9JBNygW6uii9AMGgvKfcv9XrP
a3/Oy4a3n8Vk1sTZVgagPqRifNVozeEAHwwrKOsMMYgRgvF/uWdpI+1Xo7hlBAkH
DH6+eOguEYT2CyKbaNQtzoj0bej0RlHxfjpPOO2SllqR9u2bHdjw5OkjXyhROCAc
B73lcsDZMuV01PACUpMDByksMH3ghIFWpbtesykDcjQL4D2ltzPvLJ8OwdbmbRZq
aZGPONuHtfr0Pn/UkktmC2cGF82hPQ0rsCiFI/tXyEMYwHiKA1uHWG9dpPezvc5T
hA5YM0sG9SQb8SC87LL9tTOHEDgFxvtb3/JTCPgJAc6Pzkfg7LJKmni3CZ0JCoCW
JPRLxzWj9V+Yb8sPQcpfw9lexv1wrPVss/za2K8a1c9FMw8RfTuAzuALMYbrUh0T
+TxX5xn9e1cQkq531vIOgqa2MmNPmynL6PEARtaaMFn8mWlnrlZk/dEd8aFSpFxS
jrnhie2SeJRPYxdudB6rxjSkrsDqmly0YpgsNhr7F5wdcsSHIbDelVRTqYwXShCm
ae1z1DPNrDkj+84eyH3fxELyFygdIZL2aKEiwJsmxC6vJj9ae7NPjUrVHYWMVINz
VUtToOkoI+NL38w5hkM1jJSM0I/UWSOX+K4bH2R+/VsOwIMBb09O1i41qeQLsQGl
Arbwg+p6WG6Ae5zlG5w0k0QesFsC97N4KkSdiH8iaqoEOVqJN5cyv5Z9dyN9uY8a
E7rq7jjF2EXhFJd1soEhUmAC2fqGXFaS/YDLHCm13jmVug38LVY1UbjkBhDh1tpB
dV5VHQPTHQKDQrRBEcEV/545n4P4WeQW74CLXj9ZOaXdFkbvr/o+Dk8TbWphJWDc
A6blsQrLB+3rExAzf2FhZGD970oIFekpNh9Qcdn+h+xiNJ8ODUedb7MVeV9LJWK6
/mNVeUx3KstMkRZuufQ8pDtnMnMuOotUxJ+q9r8C1gerJRs4pLHuFZLnegqRV+SH
LG9rffkRgerap5DvaEn47oi1vaAClm2bYVBY2Cm902YCl7jhbz3Ws80WgHNvt8Wo
ClCevcQMFw4d0l9QEjjAbW+8dilnd/pob5T4yHGQebhP0IImR2lKVEwAbuTTMc9j
zbsnz+wo1FLziq+Dq+VLFYh2bjkl8y74ytiS2XrmExpDA7daHLbtf6z/+BdkJ/6D
g9mQ92XXG1PbzUTMYrGQe/HEii6GRRRuhhXf74+fYoAit0zbviLjGHlkP+UWZDb+
YyhEcm+Cfz+YaLNR2vmadWrwdPUyn7oYVu+LwVxm7Tm3VujV+RIfwfk78bFzWgO0
P+uDbjBHvCXcEjUhErxz7qrwvrLHPm83F81iKlc8a0gh8W+MTp7tmgtmfPzDV7kC
uxQp4f/uwn4V1RFsjLowVSS77SxPD5fsJYUI1wSn13C3NhbBh7Fxy3GKMr2XpEuo
FdaE8L82ZQInq5udy4U3siOtSsWCX3WAPyUCyD4udmJWlsFiqVYX+5UZAR6wrqke
6ZISgC9acwOI/DJuKyydJXC4EzLu4FDNz6zfBNmctJMvhs7jzMlCAvEr8lFj50Hw
QTMsoTUNQYAPM1fULqE2hPQdtUf5OJoV3weyCUgBBx7GnCpHknivVAKQyiTGvTle
98pDGN2e4Ve+GeMBMfdvd2F1T6gbPHOqVUelAvOOSPhYewI4Cd+IKqgojFOF/v9I
xzSweJULSb+axPl9wSr0CWLnx6EsfiJcaxgmszSuZMAZt5Dvrqud1ZkFuPKCgDZ/
WVFB673PXhxQcwYnrL8FQZqHuk7NFjEbl1XOGBz7SqKNw/MflPyA7z+gdgqhrHSU
MLdvwa/K9G+FynipB+aPm9+sH3aCju31e/rT/WEuj37b6wuu9anCC1fMyoAgQDzB
6YNO/wRRl29aIN+1r5caOgaY5yWTuh319ujT/xA2kY04G3BnPhupTotyNwRUx9SJ
bv+3HABafl43cPNXoZrCu4iMHEIDaUUt3NNx4YcKQBkjHyFS1yjD6j8gp+U9a54I
iiRxyFPij0Zut8bKRr4Jik0CLbs7UXT14bOh6bVkUAmcYKKaihj/I5URgJAXDdiM
h8FsXgAsiaVF22mnmC3DMmUroTZr56gk41PN7LlNU39CVcIO1n72/YHXlKPaA61y
6hro4e/9i31sRCCcHt4TKCNtvPUo4oXA2OHIzkQ/vnF0ji+Ott8aB/AhCmse+LCn
H3GcmEo6Nk+2jiBnG8H4iL6PPZ1u+Af+Pca6QtMn6o00gkP4b04Wp5sQUdSulyS6
Osa1EmrEZ4vrjbepwOJL4UcLbyzzu7F8PDYigmwg3ukeKg1dm/8ASQM7eaKmQEgM
Stxgs+LGIcPCVEsjzvwllHaY4cW4WetR1oQjEBMOclpT1xuFMe6RYv8DL6wBReVG
Ae1r5yBH/Ze62ehBrn+OSlm2EkQ4mf5a1jppWFzks6nAFZhWJkdDrSUSTjtUU4mJ
CaprviFUv51tk7JbOt75+4esSnNCwJrEKlRpYsZ6rKev2gfbv7bNz/BOQOIZNRMk
1IgYEcNXAqWbRW/s5UUhq9ei5OwC4dQez+7LWFSkdnsZ/B0kMeWbQP0mfG6kxI1y
SEA42l9Y3T/8CmnIqvTWfKg+sVnvl1te34sarw+OJOJRWvkp0J+n/98cscZN9fn+
1jeNuTryHF4Lc3TXdv3ZLvBxvLLtQYLDAbqh/reyCoLvWnNEQXCmNCFnJatArgfI
HqbHwZNhdK24jKignbAAJsNNefzyx1b6m48tghnpZsjOdmMkZlOGZEJ7969dPc71
G8dizuNKe9dw/H98uBmzNw5mtMtlYkDLPFdP4r5Ot8eVo6KyLJV/pqVQuEyKLQn2
eJ/f6+ll1eA9QGTWmodOhDZNMDMOymofBEONqo6II9DpG2qn37ruRo40akQoiW01
BGTmBEMJrg8ZjqLUmwwITnOf/kd+UKGmu9HNeGchJJjBYaEM8Oljc+L0v2ctDAfZ
+K60oHCTK1HA6+GPKuhHaS8IHWU+OzsZGXec2fd8QQc2HkGtAnJn2bVc12TqYqOb
2g24IWBZRCEO6SbBay2JO9ynGdceUhc86Fv2FpeiOTW7ZvgowrxSMARJLe97aWL6
hFh/7Nl7u/D50y9s7pSygLXyXdNTQq6Z7UC+7V6obOFDAsEYZImTV7YyZWjUWTsN
fZelAp2Hj1msAhzXgVWqSXICBdDBBZqVaoUUwQbA7JwGaOUbrWw7UZilvKFfdyh5
ib1wEqcnqoSHmH8SwMrtHxnzsUOk7AJ7qfMVy65TcZHmvIrhhE/QWRNJwmKkoHUN
K7PO6i93iJYNkajguPNjioBt1KatzhujBNjTPEYzpTBi0UG3PM7XWRLZcWlWU0pb
j+L3sX93xbWntHxWhWWqxp4kEZAgxmyhG3Y9G4su5aht4bfJXWGpqgaQUR88SMwZ
m3DUguPT8UtjOrdJ6tMoYdP9Cmb6TQEH3Mr4X2vBAaPvBuOba42IKJvoV34tbADF
tsWbWgfUrIDjh+XbhFLzTWQVv7UCzBCvHGyOa+jpOZthciM9EuMqWAcVZZDvMOTb
oZQsiL1hivokCnilnjGoE59IuIWQRGBx3oTMJ48b5LRLsfdsj0PJJ1UTaNOBFkXA
uefJfgoTUc28HwNQ2l/JUaeHUTxMMCqmPI9IWKwKDu/Wgg4Qnk/Vbs8RUrvhcFHb
5+LKFdCIkY2NA0FhNC/OzTwzUuBD7P9Pk1dHU0N3MFXq/c394duryGI6kfQvAdLJ
xUxWpjgxkpCEAqDyEWGYFA4wENjE2f/5G/n9CZEdKY3yLxXdlZCYC1RunTcrFeg5
sMZSlNSZj0Swq5Zjv5DRuS0VvK7bF/8WxdoYlGm3Rcfg7wKE9BuwCG2bLxxw5WpQ
1wUNg/Xnz3h8lCFGwVpH5/Zf2eG4mk8KrA+joAqJmkkMTPyiIE4rZ2ndp7Zt8d0/
hiHwBml+5jDgHvngqhJO/TqIvwfl2za3W2N8SszK7W6SnbhKxs3ymq0DPdmyXPDZ
/KFZiEnB6gZUY0qrr3RPTHC8vv/PN+GT+5J7UsjdrNxkLD6mFqGNk7Jzh0JgNLeM
cSgKJbhz5gGJC+0UfeTl/6swrYhkF6++XQyj7+ZkSr58lfyFFHo83t1lmQhapUeY
WnY/MoDrXL12naSnwLJ6R4NleOwF9JLaP1AhGczJNsPzQlkFmWnzRnhqM8LYjA+v
rkuPHesPFrtVZagAIBDd/GzOviQKV7mJ76pc39+p/XPH2qX+XQifnW0yvEZcEYBR
IVAJqVofUx1d+8EW3dengHX8e/VNemRYEU2Ktbts1A3qx486CtPzMNWxX3Y/EVi/
6zpx+DKMsPad2L851RSBb5lsVMkREk/UnZkDc0+N9zUPK7X64E8SVviMi/IZ2r8F
e5+9KZAwXP45WbUg2IL+bUblPWYb7/R689ezUHTnFmx7CrfMW9YKlrxRhgpMUzea
VOpGWHWJ6Pia2wYl9F9MylsN6UL+LCRlTKTDrY9rhwYZJT7iUG3zbnUvIqszwEWI
7qUfN4eJdTQ+H7vKKk4VPUr/DVpn/1xlr8KuL1h7+gxJv5AAqQaZ+BQE9Ny53QmB
Da93LzOoO7PZILYjJuzZMHffwQE91Ydj2p4N6LujDennnDzyzW8cC3MCRwYkCehU
8HoMd9kUyA4IAAtVZ03Y6OkvHzdE432w06XIGWWnOM6prypvu9FfrinlniVVTgQR
zyVRHc6n3zuNC+1pAjeEwO7lAwGs1zb0fWGn/dRoslZjQCWNuZ0MKFRiTTggEAJR
6OuuZ/OMoaBLTPeWwIwQf1rID7qWF8HmUDmCPXafvsfshFUsNlS18+QX6eYBUSKY
5FQF28Xwz3DDkatJtTOkdR1qn3uMCjHnwWvpBdqsqlscIWCZm7a7vZ8eFqXZRtnz
Hum4GKTbCpQIRJNJlfWacqdFKMMQNm1+xuZBiePBT3/glIMsnBXGNBxhO/CuV1i8
mFEOuK5MWzbJLVivFJnT9EPLTUvkNV0IDIzyttsyXBGqzyQ4quJXCm/OTZJ0YPTD
YbHQ4L4NtpQy2yi+9S6ypKu40W6hbquEIrMLNKzz8in5ElqR9Ryi7xhXhlZSAL15
gXjfyDUBsEId7iV5DsAfPfqCCLSMTEzNhIUaIEib00zwIeAxfQ5X/U5j2UZLflwu
wbvWkn7zgyuMl4doqCmHyqYnlMYP8xA5j17eweI1ULM+3OT/Q57dez+jdtDhtYWs
TxJQSkeK42zmsdcf26NX/69U8JL6fPkmyChu7o0cJ7mO9S/XvmeDzLsJVM4vkceM
jr24Y+gJDsAinSiLDHo+7DN7GMwdqLisFgioA66TnhcXzeuC/UywwRfTVWPfcS4z
Z0ElHSvMdvPqXVCEiE4u01qND1UBHgU+TMlXUxu6IY1bnZZUYqU+8lpScEvk9rl9
yLPhI4NdXsmbtvVD3i9wgos8tMaR6bRW30r6mKIVoIMgz3Lyke+5ZI0GO7FVe2Ac
vevGnYvazMB06PPXmgM9zMrI4AfciQMO3Wg7N///4Y+y0zHGv0akgrTw3yaIC/+c
rDFz/liw7w6I5PtW8FnRaV/0lS7qmmApxts8foIEEeLGhTPEr2vZHiL0XYB4kaoh
Xr5gN2FBVusnXHvOE9k6yCL4TXJgQg0CGbZakQY65MNCpv3pbO1oHowQZu5nFpgX
S8HZMuqT8PRv0ZVarFzDOYr7Xd/IgRiizGvOKK5CL7PWGICEG3qQhgPxNG5KEZIh
l8FQXDiuYouX6a/eufrEtQzO1WPgoxTPbyndXk7Nrvy7fh8gRr3KnB9nDjkk+r6H
XmS1QSQiEUt57OKqsS3nGT6gn/PHE3/v6ZYEFUdGqNfaJJDKmHwZeIkmGvWXlO0N
Kl1deUq8SPuGZhr84cDEJI9Xs3h3bOYC1EMj95IlYHN3CDc4g9XU7EoXjtLBXFSI
1Evh6EItljNAnWF/JchbsvCHALzRsTWUt+pL1kgG58sNGEGukRY55J7hPFNUFv6k
+6JbEqK/ZflfiJqJiFmeuXEtQ1FDBMhqZu5Stp3gtMpXH8AUL1SNzYsCgjq2tVPK
DtVavz45CfQeDT+zh6kbF4e8U4IXv3hCW1tapSahiTY+wDidw1br+6/9V6CwXdr4
+Sra6+CzUDapfmx0Tbi+JVNViMo4rSKinReMok+zo1L9suPps53a6RtC7AheeF/7
Mkq2SfD3AtwK7+X+0X/8KvgSO+w+7FjWpdNcB0+qNeiuYwL8puek03Nm9NDK38VO
+xz0LC5mkAg3saFgFsyJgzuk1JfgO6Fr4ym2w/B1Z9hJexbKJ39IqWwXNLOW87IZ
3uuRDxPKDMksfqTDQyPx9eSjXj83osvlwfDvYHSCdxg23kJaciLmk4Lncvz3o9oh
2pO1weE0j4Fpsokv5YpLizMDXNUFsbs3vDoDhMoMpRcpQ/XIhCUhJtfpgrCVEayy
JvLYJROR7fwLDnC7T9+QIIdEio4rZrmcdSnyQ65zaoaQpK0wxL3SkAkmLyD53FPQ
HK3WlJIEX1n0k6BTsTO8Y8AZqBkWlJVTbPjOpvK8+2uHufJwDs7zbJZz7b46bXOo
wx8wcIPTClLvDGM0mNByt8ScAu3nRlHdxJsuz5jSEj7ffAa2jQYqtTZhCdEMlmxr
ZrZWt9kNNZhTUUqigBeVvs0G4bkSHMQn74Fd1wq9fJCRDZI4tOl5eJwlUTEzvKdc
7R2dHPce5k/VWdn1UHL9sC7CizXW/q5+RTQZ+dvl9Ns53RjenZL2u43LERavdi/X
pTV68cjmsfczz/oXy7EHIVjVZE7u4mArWl6bsiC8Hm0qVs6FRIKhuvvNDkd9OPCV
vDsb8BFLB3cx+JEA8Ubnma1DWvtT+k0y+leGWH0hCgEQofE6lxlRDx4v9FHLL+Ho
nwWOKPCQtsfPMtFKY57Df8sThbinvtktNQe452Gvds4/EZb5JS26w7CQ8VdiT0J3
uF5iy167GrKJNKG0eB+s/HfGXZrfAuyuFYf0sTS5ivI1JlP3Wz0/ch+6KZ1NcKOY
7DXh+Y/pL5R+DLkcgPnZFeuH39aCRIQRvvW3OiR1caAOWl6uYkI1scfJ7PbAqfET
KnvSg/2KE0Rq0LVv/Icv1haqPOxfo1xae93FsW+98YUecZj9gQpaWfyxgcVtbvns
zmawgNl5y2s5W17+lVWIKgFbljrrPVQHRSk9yqRx3xgdlkiEY/UgH+3GveQf5K/N
DHKygWZgTGkvRcmZB9pQ/VCHFLwI5Q+Otq77t2rio5rdDiJtfntutHUha8/cqObr
CXjb8BnPgD93W87UHUBsa3wcICgz1FNXfjQUYxVLzf649gel48z6kJotXwVeoqxV
`protect end_protected