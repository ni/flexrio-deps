`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 22016 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
hRRAlfE1xLfeNfywbrz10Jc2CogrsXRaYqxl8lra5/9ForcCYFcWwGHS1kFDKN+9
O+DlxN7KcTNU5QzZFZsUvoZOReXo7eadnymFf6dDO0HpcEIcaZ5csObs/Q4H3jdm
9bGvVLyO1hovIAtBJz5/+42tfGvfWApObp9CeJ/ZO4FLFQY5FikHdAXaYeaj5XBq
cfFjW2HnOTX0nSk3df8cbgnnDOaPOoqrGtFttx41Job1kpAXAaYWeZ4IkzlZ1uZd
Js4ys46qUBNpzxH3w29cPk2u/dfb5eSWP+J4N1ibfzM+hTVXoA9Jr1fV55ddWsSp
on4QSZ6wfuKyCoNi5UrIsnWphLVWH8kg93Kmn1u4KUYfnWVrYIxk+OQSeJL/3XGG
65NAXjytW/n4X7nlK74V6avONG9M95uUMTAZc02Bj0u/k3HBALY2Z8Pzg0ZbB7g+
BS77XByoc7c5qveYR4AcJvvjiP9bl+wjWOBtP2j7Kr2QQQA/ZOfwY1xFo83CWWX+
X+bRJnBBUoBTvoNzVpf20tiFve+bq1Jrj8ikd3FzB7qxeIiSGqu4LEnfuJ7yZamW
ggHoW6gYoa/lYXppf5r+Z6G5D/xKrCur/9TZaxHqHoeYT4gGnGDkMiD7yB0FiSyQ
Laic/zkgT2M+yvbBjboXFne3PZqFzFGM0ItxpMoVVZS+QqT2LXoUE5GdwZC7cuNS
+PPvBP35LRIq/UOqwV89S4nOBNc8YTBs7GDeJCg1A4Nw3XMav1kX5wHnVtSXp/Du
GcBuTbpiAbKO3b6EiSxh8wy6UEShw1ewb3YT3XxhqXRkamZ4pRC5HQV7Ml4ihOVh
Rf0T9mQ3txUXs0W5bPTAvX8wYtIIfau6AzsF1teRv+p5T7lSSLtAkIpqZE27adEK
nRNPxxYZZIackvUWnBZmAorJSIL0rtcdruhfhVWiPUwN2iCU54V86nj0tCYEWPy1
Id5OIZY1gEEz5hHEkHVJe+PbZ1rf6gdio8l6k3s1JogOPYtMLfbGyo9o3AUeNGIW
OSAvuvWXgUNaRtuG+/2HKAmDH+Q0Sc2g8nVPzydPpxPNg4RjCA8A+QoRVUFCcOqQ
i8wT4oVYNgCuw5fc0h4zDqaSK88DYcerAClmln0BGMLbP4SFfBo5qBnubLQkIQI5
HEHPFxcJ6Nqcj1noO0Z9Eprn/fScmA2mIvf2AibVlUcr7pNPtCVkvm1qfTIzfq7l
BM5uj40s2vBmdaUwgIDrzm+IB+OTrQE48uW8uRE/Jw3uX5sUwrf4/ACq5cEPMo0k
dJlQE39sTZuTEbc4fr/+TrDAZAxscdnTtRNVEibCDbqfZcP7642IGbEn+qRJGC1w
UOtkOEj9s3ya+wzGApKGZh2mT5TTl64IWzS1UnMAxINWWqcc3p949NY5Y9c2X25/
jvoyMQMn0HDL7Qer/tvoaRfrw0yxIAGlTWiKRZ65gwnWdpRBLoMcFH4TAThWInOU
3GQyvGzBpGVl6TyvC0HjZQkepRYl+UgZuvH/mYxccRMGJvVwCfqncWkdxYcSe94F
O835/FH13FIS432O5NWuqX7UyiI8iI5m2v2+SzwXq/qgUoK7URcEGEFHlZFxVQof
+kGZjIpZ/hLx9WZB2Xn4To8msB5IEIlKtrdxRXHr2sB2Bap+ns1haTTDE9q5Artm
12Y+msio1G3IEfkK0q7+4S/8PoOq/5ypcOkN6eQoOMJ0uGJ/MnFIzUUTKOiHIlQ/
oaaMBCrkY0hEv4DOIsqwaz+56XssngnU+bncB26j1/CV9e2JQ4yEDoMsWRXIQvKF
GSjtqz7Ut8UVDSBpnwDS9a+b0xhb5DvjwGGx04HRdzKAC6dMpEkE0Qh9MwVuhfb4
VkYAYcybRSEnkIzZJg8e38bt+1S5F+RugWfK/FnNTiHfQ2DKIAhcAqZafBw8MwbU
fCYBDwrOP5pS+XrCN4RucN4M63uH53LAKUG2iGne7aDYXx4iNMat0es/EWaOA6ld
uWdaoISMBNhkC+Iv96eq7TChzVmvEV1xAOKL88wg8cRYmelQRU+7tndxMvEnuZFL
ZOT5UG/DQmE6CbNQNAAzQPoQ2awxRLRXGBOZmXWfmsrf/g5HG3UchOzLVXenobGo
SawI7QXilWmhS0CThd8Nff7OEx3ETz8D7cj9Hdv+UuoSGE58mvQi1hDMQ6vMjulm
pRW5V6djRx4K4iD6yg9pxkUZCa52MY84eLOWOrofwnqZGwPTDS9kPCX5Cb+OPNwt
ZA7gctPoisLmVTZsJOula8lge81ARjxBUf9Ie97aNRy6tuqK7UeR0n0mdfz2q/9p
XqGfrn7b1R0JXDvM2M6JFkE7yzefTQSzZta0wgwik+YEbIGdrIt2yOPvluykJGCa
dyr7boM2K+uxqTbEfTvgsgz1llYNHoPISz3UGqpT55/QJSwx962RY6u+MfbT4iZM
Tu9pmYG8rQLtX4F82kgAwXTvzBEm/652uopOGlCGD+9Yg6ctfg/8MuxNTolEHvTS
qTYP4WRYiQAujcTmDkuI1AjHGAy8dIUl10SFLcsv3QP1BC7BQUtSd1+3oI4Aea0e
nfZjlDp9kNOfyZ6/hZrMApLe7DbX35roaM7nVIx2tKCKxG7ks64bYY8bpnPLAdhR
9ikF7huYIFstu5qwphMOHqkvkm0IfUW5Ixamplby1AlIyslQbaJqCr/frIj9ZJcn
EfMgwXghekBuups5+Reusc41yxVK4HAAhN8TACRVjChgnasr/f/9YHwNRegKROuA
WakQGrrWhwthVW+H7rqb4eaftjB2nklzy+4U25ssXcT3Ka0e4a77MPwycfzAsrY0
KVWBdhKyHeENEROFStcvqcxkWgC5zP924hARgfefym/mN1yTj7hARKXqoSdf88Tn
Ka4JLh+oHD8D+M9R4zLZW13znVcorZNMOwMrtiqWQ8HiQYnAe8O15v8hXlb3yPHX
iZrcjWIzAJL5jDxo+/9JlJ9Y1Hb2IlNKDo6YmB497d6+ZNHUajbteIgLg6UkFbw+
ap7NHyQHV023PaI5n0cprzM+ZTLXq+g2x76TvnsWHOlUxpl7qGeY4iYF4xUoKuJb
iTo6UzWPqJIwW6pnc/79INWZGNM15NYuk9fyfGDBMks8hJTJqqUbJlFoZdv96+1M
bCE2w4P+w5KiudTpEwEdyxXU7QZIgdrQZi42X/0ZvRjGn3vf2/PMKyNbLlk7dwdd
YNs0bE2Z+PZidJP15cZbWfhOOzxuVoC2mY0jOXpFvZW2vQLLq5m+pyh3dpRazfPn
krPa/r8eMXX06m3cyO6F37FEnmHHM/HvS7d3wGbAzCGWyY5hS8mxOdKZEbSpymK8
B1RBZt+99hcdZi6VSUEvXwplro8pwqHgPjzkkubeGqhatLqKUbpYk4zQsx32yFWE
J/yjLLmlaxw5pIAAorjtfA/VhOP+/s7VaPuL9Y10e+KJ2Inst02dsE+De1EQqGGT
puIzeyxCpyAh5ci6hJK/8Pcu8OKig/NEgV11Xmmvt+mHH65zSpCQC6ellCQOSDdp
wfINvO+ijBg89bYSDsW0U1KKnczoOzbm1I1lQsCXwRJp/HtDnIr2PtZjxYOK3zar
j9FM7IbIbUnt80fSKaLloB0oi+6fa8RfFsQpfPjRFTbmO8KdpJI4HhkTa1b1vtIm
32GdEyjljH4SFB/F2S02/HG5eXA0AYGp2JUchm6xrK/jrond29WBHfqA6n6+eQFM
/Lh+waebi+vTneuQRXLsgfdu2c0q1fAJVy3rYrATZP+8jmi6gFidg1T1cwJ/e4s/
1zkG1+YXxSe7nDojArfTCxRZWyFPU8hGFwnnWTjVZoq1WTByqqBL2KVV1Gzyt/Ia
o7V9RHaOLcg4YyZ41viR1iDsO59xng6Ukry52E2ZZQPBgsocuyryI2R0uD+G9RV6
in3+ygWrOi07thYfxXHxtLnhKe6MLWHsw86UhRvalNdNINgmKvq6FhsSdX17+uwm
6Mw4RD8GLoBZnASQ2vUmBbdBSHqun3SAHdHUdIlW2K1KNEGaDGTYr8ct2ilB2Ulr
npe4O9E8tQtFaRci+21Jv2FTLsmCI11V6qAXMkTbUdfRgW7W17AU9Si/bnpiMYrQ
8q7nJVY1amwtVZKL7cVfWfoV9Y7x2MyYQIdtNG6F4tRFodw6B3PGn2BFsLvo1MEf
u0APe+1Tyl7c4/qnujHdH/3+e1xUmRerh0J2W7ExbAz8e5NuAXu0bjLrYJGdxRg5
gz9bzUIw3FjuFIGIN1lVlJMGdKhhneFdnaK7HMlihSKN5Q1YJr9vSYsf7nP3T7Mu
u1gm/SuCGemtW+kwdeQFVimhRRLOHBrVrp9BOefrlJL9Cjk2B8RrAVf01H6Zpkjk
R72DPlKn69xwPtR1YtOsildNTl9qjgPkd4jy0qmSvTQd62komyhLIkXbcs4/Ru8m
/fvBqdc8jGG8GIoPaGvqBZ6AgPzaZvkxsI0ziMOrsbHsDCrhmoAerS4v8DT9NxqP
TCMk90+3OwBdch3e/cK/UZeMiSJqRj5Vi6DcEANjCiBU5scCPH0cpCw8xCukth/6
rKOjWS6dd7R57ciNhM2VMnc8jLoAXHfFtAXj5MvTh4G36Mo0bxLx+U1PiYlbZ8Kh
b4kg3VvwCI/wZLBAaKoRoZeQoPy7pBzXDz5VENSVLaQHc5GtwKMjv3o6B0V+yKBV
ZgYcnKO26C/XR7cD133zMufbeHH9xftUJ6edTZ90Mb3DUlA7zMbDIKTQNPs1NDig
zVxngMkMaSxLbrVUbOgpXjXMmYCmyiSDqMzCAl/dr5rRvjj0HRphpsCiNURa9Dhm
QYm6jI6Mot52gtAIzqn+pAaaAI5wlxoIabiwxrqvu+PiOfoXq/mfY152VuiCscUx
GXjLxlFfi33J6/R87B9xhuB4ZNITkjPy6AHcLHTSwXk2XJjlX5TQNb8mjInDF3Ze
AyFYGSbxJ5uRlR53e3peP+KPTOr92FQzQzymwGjuF+Z82AHvd7Lqldg1sCdgjjq5
9ajbXnnv+hvQRtOmju6wfHDnxq1sa3yU9EB1f3sLIUrzMPxLr0a6YQbVXGatHjXy
7UhoP0q878N8KH2nfQQGEElzaKVMoA6g0/TVtxKXSz911ozzYXs3snQQ2khW+JhD
xGaXLTvHTr56vYNymGF1sjuytMpdrV3J8PgVBUSRD/B1ffjYDdDLX3A8OZ93vTjJ
/rjmNEcWTaOlYbqUBvWiZ+MPP20zS7vshucqzMYqYA1MvYz+lBTvXt9fDOygR9OX
EG+x4bm1NvHkKf/lFd4LjSsAdUxYe5ZERmSoQZyD7ky4xmmnrMrgRZ5vxU3f5pJC
ZPkxwUY0c5kcQ4JrQ43kYXZD0hVHcIYp3bOyXA/eL5eD7+LiDFat019oYttxVwQD
zZUOjdFShNVwjKKRrF3lhJ2KSbYsGW44/kZMPqOrjMyU9oHowhHWDA5cfFUSURS5
4lOZwRPD+qJIIob2ykTdixsOL21H6OSG0pZPuYgT9hw4tRPB5CSDNIDSqNeDwb+T
VJRxeUw+ke/W+GGY9pXg09KjmjXKwMagLf5l6bTVHOanHxdtcRNhUAKmO9Y2BZk4
XpTtQXzSmA1iRoNeK7Mw5mohQLdHzWDmkaqeAotGua3X3a5bZu/jjEux8CbcujJ5
2CwZgxEPHJqIDkQGcpnZrlPU1mY6ehSkT16UBYtoYDXKSJUMquWUG/5f7C5ZwQg6
xTQJTqcLxoaWbht+KteIwE/Zx++2ktvZhRyYCGKQmeEsnZhE7WLK4KpjeQDGLhbV
ToTnoD20uUsosF3KPbGhNlI5Ik3aWXhMj1LtzsGi3pIcvZP4O751sm+u8Kkdbil0
0RdFE+HEB4nY+J3azurCQSATSGqNBeD2PXDxfIUagBayXBXrObxlIb1N7HD8qhsc
3IIv98fm2/KvwgDsp7/6FFNpLu2Y3XfCOEcVthY77hnbkCxe/GBM76UilKeJzZF1
roLKqfR8RXrUX/dnUxrD3j67QVsm9SVCSNlyc0R7eBbcs2+/rIvqDHXo5Cimnkhz
xTVaq7XMbdpq2kjYMq9FBFEscUuRiYiZZAXX4LtlcX+qvlZmuu5+DG8ZVRCFsktz
f0pacCHt0dTN4zUPD81cQgBjgk3k/iVV3Ch+5UJLoWPzoG7Cli5pXfzOoEsznH+D
6lqVkgyfDt1Y3c1AH18MDbF0O/85Jigniq2qXCu61pimMt+ONZOTW43+XOxVI5lU
bM4oibIXG6JoaILhoHlehBuG4p+era2wMl9snUM1BdFWVs92ATc0hyXvCo72XWtJ
X609yKl0FTBjSp7LTJz9JU/b7DfQcCd5JGSMC0NkasPwukzk/IxT/hDoUgSwQTWO
wr+ED4eby47eq9miI8AKTct03+xkNyUd3rvvMmIbcrY984TCySOXB+J6bKIkutv9
dAR/jUT1PhV3CT1JTrtbK9dBWgJa1ADTWiRzx941Xz7b9EUhLwcLiI5bSdo1sGD3
CYuDO89JLgoe79M7HhYoqSS+tTSFMC40JYqAY+iD+EYkXqkjhY11t5xkgdUE3hsw
7sEpoLINzkytR4s0UBf6RCn9RFvb1zfxdK9APjqeBj78Xf4IrwwFbaGXoHv4KdER
g4XggVlfulw9iuudOzyqLojJ6QAIiWcChHjP8WrMP7ie+0mtWmxl2ebHRbs3k57W
exRDuXimvASaQyVls0iTk41aKbPUVVliKNsdymYDAlB0TBi5BGK/XRU0g11JePfE
PXIwF5gF7+oD7YPLnvoCJjoooL3sYPNH9NZyYF8HvB/h6hFF/DNTBpCqNjNARrWR
rWMmRXEPYvj/hT66mRcflL3qKCp5GQtxxCux9WihFUqPYDWJjVyPmDhZ51De2v3C
1/Fze+6savr3KUuLWU/d+CDbXYSpxxlMUgZEHbIY5nQeEYV5XMbVj1Bcs4YVYy94
4BNK1H3fy6EqkW8CWE+e67+mIklh87J66g1bMENOp0fOm85nU42Uy7cHti1b4pi7
cciQTYRlGnsGX30L9dDspNdP5VR+RrUQgVfVUcBXbnExcahZpcm90tL6QkHRca0Y
+lNv4yGSjFHwWQ0sZAnxYTYlzEOBi2+5CV8iLDGki9/k+fqkkhIbk0TVxX3Nhkxm
xC0jC57HLiTLr63303b6KxfG3uAF9TzHHYyxgWTxieh1bquPDzWoUu9HqhnShmbC
Maj8f+cHQAJvkMsKRRAB+SpfvfoLy1j/PhU5CD8Q+zT2TVrzRSpjlKLLjK55h234
D6Od1fXpEIRMUJ58eAGwStjWOWLM3N9+tTGmUMfUzbcvAp5GJxfc2e0TmHecgoc9
fBCzi7VghPffqDGo5JkWvR29sWztRww7ZMEW7+9oH4rB48vmOo4ozXDY+705iWxg
KyypF4T3Fg1eyn74zup054e2SE3Bmm0Wx/XL7K2drzM5P8IM7cIF5G+p6BGVTdD6
nAN84ybSVnwbIrV9ZKs1MURn+BKOFC7ANg/12hmGqf33ZzYiCi2f/82amwbRYqnd
+v0m3xsxysnYBbdfDIjQRtNDNp4vKGVeqC93VulcXF42W5VV7xRwJhCt52aPnwPg
b8HbLhUv9gT8eJ2r2y4Pm5MKzadmNI3IOWPtnk3D55k/0+cJUZbmALLhL84NvMYX
UCQRzQPDJhafBBQMWSjzj6h4VUlRuPbiUkRpJpcnjNDjRkHiMErsnrMCdIcrubH7
xtuD6wCCoG2GjU3h991eodLEOohMlhGgJQz9Na936AHH81kT1kSF82ISRe0/XhZS
bGoZDsWzEe+M+mD0ntH2WY2IYJllUXHlmx3NxOnirOwikdrPcwvPZxbm9dhLeqiC
7LdwnoH1xIsoxxsbzNtb40CHTRcMVBzpZt0tY4m71PKu+m8x3ykSAG/Qfq9N9ACf
c9NLioHJ2wsQkTryH3bwbum/J/SuX5YBf7AZk93ndyOvS4TRpExMlW+RD2Ux03a6
hjaCnHCpKcqQXj/m0ju4QH6NYTdMqHLvrKJuyNUStgWIuCHElmJnj+zWc1Ht9bsg
L1crvdIl0WTGDnHkUUBw6tYiNc+4WEQTv1eyYvViTtkU6QiGIyqt8hivaYy8bmlp
stusFZc96LYcmf28Ndb+g4cvI/kj4C8qupTHmYFNOulxdkOVF4p1sKV/+ckLJeTO
knb+cgKk/l1+vOQ0htyKaLQgVsx+9GfmfBU2IrjkXDfKwd+T+X9ITiKnnOvxmyt4
AmtrTLL7GZ6rCN5sDcWq1AT0VW4yB5PYpQI2yab6ax5iQbIQQrVJOQMlx0KQ/n7k
X7S3pQXHMz2Yes33cN8H+07DRfD+ox6gYGWhuvTNs7nE5zP3oq8dQ6FP1DPu10KW
Ukl48B4PrltWFSS/7hXkNkHcfltgYMP/NQMCBOswMPQEGeOgJ4HkssH/PZIag1xA
WfVvF143b7KCEq8cjeyudGaZs8B1YVFKMEBG1CdwHB1cS/PrVaV5Jtcm8GoUMHxH
lrFG2RF9ikYMStbW8TTE6RoMpNY9Yre1FXCg8z0WUfZGdSHcSZz0THtISsP2KijU
smkqT46B8bBiV2btkuZgye6FrTA+s2simPNjBAGmFm26AFbzhicP7ylKy1+uxNcy
MVZtMfwYlMQfShtIk6sQZK0V0HYIxQYwi2KnbFCrW7no+u8qWWXnOYeAXtuSx2XV
hIHW5h6GXFBQtIe9yxRIj83Aq8eMXslQ3MY1t4hs+H/QksUI5LC9/8d9CtrKL0cc
fFz63FMJSmlA4v6RsMkbSnd5+Bm0M44OwkBtUv+HbSEU0XqJUOnlAKwqBmTmM0jY
GFSh7djXTkm938bFnPRj6JFjrP2II7sJ3L1umMlvQtcUADR09Xuo91NySKWJo2sL
cSeNdLoyDndGVP9zHUz4O0OmMyXKTn7n88/xLIqrqfQwzsWNjNIK4dU+DFZqcmZU
gHmGK1CmsFJx44x8MI+/KFFkgNAh60YoMx1RhVXLYqBwSWaLjUQMJ2RWnA0Xznmw
DnE0/9D82qxtJVyKpP1H3AupHHKYl6bXuG/uKhINCU8Bu5TaBNeTv/Vu2Wm/YPUB
jA+KQpB3AmclKAFZYuYQdXgbkTOirMbHllWQrbgtSwnczvfQa+DF+KjzfMHix736
wFHHSDoQAWyaqW54EDHmJvbQeF2rHT67F9TivaAaq7eFxCXIaqXkU1ex91jQZuMM
5EFw+4sN97qNSVx6fpaRD5zkccc04dCme2dIP3T2wLWIeulQ211rN4jMD9dfOxKD
rPKFwAERdHH5165xENDjZTK4pUjYjust/sP1pAynkQnqf5VdnL8zQk5zL00zIViD
Go+YDaRuBNXPY86vcwsWKZAHQNs8/GBbkW9ZeD8iMisubdm5LXF81ERUXvRh32Jd
QipeW8pWEMrXW8R6zntTh9cRwhXpaTlJJvSi1tclDCOlpmDJhhaqmYcoC9szRC7M
ZElGGBCKKuQHWJyM+BEYSvsR01RL1vvS0et6J5hvDDZK3Vsb0ARwdM+/Ag4Am8mx
CAFA+WHSeXEy3PfYOifwRGT0xgLImUlSE9KJA1XFkhOeFleuVu/ofTQ3yqW2p3ZE
vMLNygnTvlVcDESxn/BLxqgEUicU4WVQm/ZivOWw0Iqesma705IrsBj2j+395ZBa
21WvVrFhozx3lme3FXwnohKRyg+efSgqTZRJNawu2WrFOTQlSKNkr7uQ6sRDTQB1
KO0czdkbI6Nu23fHoYXSleFW3Ex4K13QNSJCIBLAB/yjYcc7y57S+Bw/nJbg1UAG
/XNBF9BicBjiZJ1n+H/t0VByS38hZ5jkCW7xKSBWaG6lZhEmca/GxFC44qtf+i9L
6OQO1PsApoZRWaGjTyCcm1m9/jszH+wtOpAvApGAMiQZrfRHV0KEUZTE//wt0Cbx
L8OsyGCC7iDT6E8ubh/xAXtCF2tLXYh5x1hyqt8aoPpeSa0ELrmb/02++LdQD8RD
ZiEBH6Hxa7lfQei1MXy5bA5xgwIeC0s3tpVznFy/Dp7KTpwolieLFW+GSs9b4++g
hv5QrJv20GtpPe38eSqJIr/5VskMauPp8eewl/+GdrjQqa1AmcuQlropq6XH//aQ
deoecJukfLKaIVyuyW45qc+OhhfYk956aWX7BjwwUhL3Fe0bt0HOZ9Vvn8NsRiFB
gR0vwAovrD3LrdSJnOExHdmLSBtM+zNDGtZAhah5IzLNwj4YBGZKIcNxbc8lN0nV
qep6naOWjsv5jOfiGUCvXk8mE9s4vM4567yjzKeQXw2NN1img7xcqmbT73r9mYqm
u+G/67zmGFOdVmjZdNxSBre1hDLe4RbFBpQVUA2lczEu0UOOdCSJ+LkIQwdS2Pk5
dlkSSEfVJr5/JtdQEat062+2yOboNeq3g+xt5CddAAq3h2hYJUnCrFpiDRXeAgHD
ouDWwqjuDpt//U5IOtBERuJbskN6HaykOWMmjx0l2Nt1qM08CVzei6VUSlJ+4pb2
1aWki4belBITXbvHLXEm2CYcgfags7N7OxZN9cTD8wbECWcqlQvQa1vyhDDLjDIn
qSjP3UFAHPXPtBrVU26oq7AZVJpr9vMaY6MpSWoLz/phbZCRi+aatjVWk8EV6wo6
I1qUmcILNTQ/lIa7YFBdirfw+9jpgMiSBHzQ2mq9Nh7ZPAxu9xUnpsO7ioUkKu1n
m2fG4lt49znhwV78rw42lu7ZKyttUQ8ldL8KIF1+ohQQrEEl+66UuqnnprHsJ2Kw
k9yaDWkiLC+Yn8DEGyfEKpdEfsPZBPhBnqrb2tT2/TmpeQZq/jEsg23PUsiVpogt
3bJ6tdAYGzS285HpM5qUi4n9dRTRy++fUgczAfWjCKGw4X5mZYrFsu0/H+sKTIhj
KbQ/3E8vHzt/FNYZxtmk9DJstPxidWH9dAX+p0Y1Cb07GHmT3f9IOLur/LAY/1f5
+fam+8vNz8CQnijY9G/a/4hylFs1PsPZF2q7QYw8VdsbrPN+NQYbXqMnUac31KNI
axSGkSyKf6Dl0zPk9VbGRyGxRvZ9Yp+BH22yQvxH8zXN25wqPPwEyJAXBwxLLEU5
DerT0/E4Zxs+VUqdWi00EU3Y4PspcxRVLJWqa+VwkuBaYSs9qsL4H7vJ5GK8adEz
a/o8hxvO7p7cPwZx6nBtncET93Kus765Xe9jHUS5AxWjaAxJ6YibsDB7/Uh0y0c3
xqyJtqLopz/X0HNjUCN3xTzbzgPu7ntH0fn3GYt84A6U1vgFV1kFk3nQO/9xEVsm
Il2dKZt1p9SZG/L0JHKDhnz+IAFSn6G78A8ca7TEXdNMbbZmsOiT9cd596Oahos6
j/mRtKzSnCKGnIphDRTV1MLMHQrgKB5XKxxqy6A9kTzwkHS7ezmumZvi5ddfxTo+
lhpHKxJaBj9QqirYqBlFmbOJ8hg3NHojpzw60H+hOv4jXhwa5xZbuEe6rupbRw9z
l1jTvXVfOhQ66tLBABu8thGSt1hvdAEl0l0EFi6/OZWe5LjIE0Wz10BYMEiqImar
aA3y4y3tsI69zAXAJvrmMtL+kY63TY91Th7bqphs/+LHFkKInRDv36RUqaVrqJTE
SnYGAjzckSqGx0F5pWa7mrPRaOBKQafH462UgCWFHg0Mkw6iW+ixnc4IYGRvFu6v
L0eLN6IBhdH2kXX8O3FOLwcasy/XE8wcZQ50hurt+MtVq6bgNzaIV5i0ppaAudh5
x1FQTRxJn6OcNacU+TUup8p3R7gh3kPeFG3oxvN84wV1IkxAhXOVp98ajaNgMyIG
JvZ44D0ArIoFRflrhA6hWWZyXXyUiq5MSAAaztga4aTc9Ps8vY2ypJrxLQYUJGtz
Q57AONEqJ7ITfwT7cH0l3tM1Bsl4Hk4qjfiTze3JhC3vUx+LVkjR564/Mi4lTJab
h9BxJXl9waWwKvzo9OQEsAbBtBZC7q2ybOhooGUM7dAyEpMax8qVrNTdZmMFMUwl
9clneNEu0HPotfZgkKe+EhhqioJG1cl/VQn8VIC9W49Zlb2IBzopMKPWHm7nP8vt
Lh4ygwMioZX6KJHNabhw8GtkGmG8wDPO0H+JsdyKNhRJmvj64gRT6RF8xPOo7edb
zlAj9qq6prBBnMINXYiabGKtAcHWrUSdf94oRz+SPSlpIVP2r6H0C717ZzsqViYo
bqqw8b9/+5CHe6AEbvbBSurOKzqo7ZQOFPGB1tKpP1beElHGN7P6GbrNgDn0nrdE
Ga7VbGMMVPO6XSWP+hf/j2JQFVLvwdMtsRuXVOA8l4w5S7Mo8e6GMg7Ukn8qTzAy
07QbRfOiLx2boPdw5X/lvQLRVJs+bV9PDjJKkFom7BU7XPPwC4SuMFExd5dNlDY2
FDpGQ6l0HmaVuD5tv99mCsjI3YjvIXRvnyBtSbJxZYeSj/FfVsvdM6+yDasfKVna
tvA22t4oYP0PnP7eNepmsWXhOp72IALxoZrsS5drKHgPW2ZRUrOG+O4z5vIn1xnD
ORSkNrjki3bgZOTDV1Yhz4odDEV1iRS7lvQwkw9pHq1OEVLW/2DrhqZiOymlIbm3
Ijl+AFv6cXU5MXuGwxUDBlVtLAvxXzF/D/No23ZfEvmfMxE7QNlFeCz5vhSGnnml
zEkanPVguTkqs2cW86WTTa1AthN/nUZJ7Cxxde8PdKBLTKPAPmOQKE0aTcoqj8xm
wabpW+Db3PUoqtgXVM6cre/F0D69D6Nhe0dsPwCQv0XraFC6QwbGocVQ+PjQJmge
xGa/Cgcwu5+QxITnrP//zWUXtApc293R97bfZUH0w0LpyQPHZGHgoXE9lPKoIBXg
rN+DLzVjoGSSWxPo1UainV9azOF8JQKjYsesEDJsY0X0BriRH47CaaPYRvfXJJYV
C7LjtmYMbXkmEidBUMpfA+kqwOCQ6TSblIUTl1MJH5pIBqhRlMPgbFBz8t4b1LL8
d0UHBJlsxfkO3GWdsqma5ujHXBV8kNXXeORlUuhEK4ex5R/+HiDhQAncsue9SzXT
mGwuda6rSDtN18c3x+iX/sfIfiAp+7/Os3/4lrOwuO5vyGC7liez8YNWgwmIBalM
WSPL6JCRcGOs75MNM1DzHu7ytfkiLtKXOm+1oDHBs0mes3ltzuS+NdXHafdaLmiX
uCMJ2J6xdxjYy+2Pyc4p0Bi/r85G4kh33qAy2JsLP3J6ro6PTg+d+baE6W/55Da9
WqFd1E5iwtf8wy6rigT+hmvIMB1wPgtXT/GEWFur45DxlnekkxkwQz58faFiq4CK
b/pv1l5GPEakJiox5v8HMrN+ivphzjgl/58TCSylROYEyxpGEGKJwPdPW/tG1hHv
HpveaWTa8hGw2qKN3FZPti0swj8ZkPPBNy9RC3JnLTcQZbtdeRbcc/WF8iPipwK2
M1MD8iKmwdeszPTHl+YMyL8DqoobYz443BZnTqIcoQhxbXWxlVtS6KISB8PN8hXo
O/cibTYKvBKvcmOyEtYFw0LUVIXoqgf9xiEjE/vxirtZwTRPfmdH0V8N4QiY1puj
ZhqRJLbKyHhHd6QB4DmDNoHGKy3/D7y1qTBMVJnmbKBXzFGwWt9Dez/bgjUhkksl
QOkwqyEZMJRHtdMecJwOuOJ8cjDeLA2Ito3OidoqexCQU5nMY8Jt47N6PH9ZNfWw
x3sa4awyLrCHste+OHbG7gr8cGPOij80x7bVKx1eIfNRglptmDQdqFzR8LAR2405
W0va+TfdFmg/a7GExJvWxysmpysj98q7+MwI6IG3DrKKlO9wYO7WQHrnfn6vUhAd
A9lZ+q6M03i0ESfVz6J/BTZvBeBCnM41DuHguoKCFhMAoRGTxsePNtgVoT6dVt/I
fyDuONSeHfXrUerORALh63aJIzHNxYxx/cxJomlFoOXUNI3XebNX1W/bLjUsNJ3f
sJz/YbM9pkwiZwlcyYfUC3Vcdu8dmWtARx98USmIGiPjxbXxZHOt22uWHQfMLR86
RdzcLAxn9QOOEh2nefs6DcZ9PG1cHQNRk3vEH20irb+OtSN0XKQwLVIKBydSDgxQ
qcD9adY8DFx7P+uHGPjo2lkb1OzIeYglbJmhmN6qrIqoazs+H7vcdV+IqQ01+JfI
2NWLOvxFPqVSAUnNr3mBmVipKrXXwfEqyEENiNJmFCbT6fLdU/wIXoaf5pukCz7K
TxcrD0Z6a2OhpHMANe66y6CCjaCcHZEZMXzQPXu933yllI9eYGxVNIVXpmK73Tr3
TSeNGOZwC+jB6+Go8pMPdQydicCOzTkb19rsZugTVQM/CQuQ5rCPsF7lZHJRzTb0
0HPBTIHmOWOXrH9Ra9Sz7FBjaekBzOQZOq7lKYXWLDP2OIgBzmlb1uXZMrxf1jxS
tcS4/gDf3v/cd3MaL2ths+/ewyQZI/KP6PYDZA+6m+UuWiLzu6taX0zSlASHUMpO
fNwuG9bX6tSyYe9ELYZZxt98QRNqUL5Yi9GX7GHrERzuN++d+mrTM54qI4QNrPk9
liX0Xub3UBNGbx9dEmiwqB695Dcrg3xr6z0W5w/E4lYVKiVkAFkFJTAw5/k4izIG
5b7hRCmX2pOg6ZF5qy+Y/T5C36fzvv3QKmdhimlTabocxDSVxWUgoDZwampEZq3C
XkLKmc36irXV4DW2hxs6LV72fgrQWixDfVH9JzzqG4eGeJKgPPH0rIlCRb4jRS93
khTh5tJ4DvZThXVAE4xv3pIJH/jPK3TF6wQp4WoY3N10S1LRloKoaiag/HVbSkU5
SN1ATKBMc2SRbD9KyfDKFjb5s4JroyZ+uJ6Lb3G+639ieCLkkM8hQVyBGx5zeNFj
o7OCTf8Mm82gtL8Blawd8LTGDoZ0A7oUQLFZIiTEU7PXWm+fmeAP/aTmSkOTtrwp
T5OPkommYVA91Xl6sq3JTTFkNqorHbDWGI0fOMGtqrzBVnjRZvFTVoL7Iq9IDJYz
VKUJZJHG08z4dE7CXLbnBTeeUGOL3iABF9cD+I7/vsMH51+DRv6ZtuYV10eBsVWB
7KSK/NFVNJlIwKT1dznYnom3WVPKtaBvDOUkLgmZ40VRw/S+5CuVXHgoA84MwhJP
7MU7Uqa0lIYPIvqTWfSLBFBoJlvrQyRz7oesl/7kMr9/IzmRMS5dYhliOqWk6Uhs
DOMbhajR3fLFAzcg7KujXxP+Lg4HSoAiJnCOSnSGnOG/g1UFsd1AtpK6/aHQTlSU
QhMKxI6aWSQ14IrTCDE0B2zn7wDq/p2FuvNemxBbK0F0hRsivi8iiG5syhe21H7P
r6prjw9BPzrS6IOphCxYFNP8sYq3g1rqApMIwpbl8OEyfhLnHymdWQiLdfwot310
o/DxZtnYndYhXEsCLK668jpb5w7xACqJ0tb4zAzQkxoyz5M5dFs7v5INYImnTB7Z
L7M5tTXhUNUwTNvNxJRKjYJRXI6GTlZ02yZuRP3vnfbRBsHJORwuJxfhTHqAzA75
QqHwc8rf5mr1sMCr19KaTaGLyCBtqg4s1T4ZyFEiWnDx3iS8RFcwZT/tV/dGyN96
UgnrKPE+bjUDdK3XE/FuflGji1W6FlNWYxQyG0zmJpK+LjlWhqZ+jH+376c5f9Ri
ptEAL9UaZ1hdkLKfIhVoLprDY+nMV3lKYlF1xVTbj6lyh1gsOOC87gz5D2anqRqT
Hqu18VvVUY1xKvczVvU3Q7y1aLG3C7wLW7oI4Meqlt34JHNKaketAVNg94iyOTjM
NVXqX20fdAIGh9N28G7Ow3DIMfC7mau8aA6HQLWK3W7n6lZVmqcImZSwyEjhxL/e
TBZn6EcMjYr6tBA4NAtwor3Fvm8H4xvCxzOKtyl/Y21wndayd4qHx2c8adlRzJ7u
QDuAx+UEmIZjM62Hv8wfKeIlel7LkBnniICFp9ARWtS0Rket2qjWwTtiFFgl2vL9
EhU5BVFFyjHbwb1N4wuPt+O0XYUMHA8kX4rQtPMUAuI1N/CvGNBLZrpvlNArxX22
RPG8j+KjJgOU4rj1gf5AZN1370+dvLkZdd++p4rYTvuwnieKl1U1mVQUUxnQ7Xf2
8czQeAl342oa9WNgoXhI109VOUv09gGQIdipGakMW45JE0TjOXOvWHeM0qJ5BuMB
VP5N16M6yw3IOSj8TshcDmClRiRo82q5+u4a19Gphe5/pKCHT9DpmNwDc9BB6Hc0
r5u4tMXjelHJcfTQEnhiODedpfYqvfrd4G7t72EQP74RANeoFPH/i/t/mnEXN9Dp
RM6ZmBV87V+wqRe1klCJgWtmXw3RLTaR/QL1a6R4uod/vXtowUHb9yuA+A7gKKLn
/K9JCcY1bEwJDmEKAH5nne384S0iOo8MXVyM96u1uhG3tE80NouJaOBOzdPiZs9U
Lvn5vEp0KvOzhGZDaPd8TqtPPEk4A/vrRB2C1N01+iMn8F3qiElh+Aq4/VT7F7MB
BHst39v27MF8a0QDJsNP0UnlZD2H40YhokJ6eQUidUdr8Njh9n/K28G027Nk05s2
6dL4xKhkbT4SOajIvkfZb0dd0a5dBV35tN5d+/nqHS650lDCWE2cIdpO0HAE+ffQ
zlH+5pnP4RQo6SK6fT3l7ua7zNXIo0i4EF3MUapkbMSQc1Q77IgzesOjbiif7Nyb
8eifE9khgrGGMjkbOW2JIm83mmTZ20jteqnS6JbO88gUgKERxyx6FCojqYCgDKMZ
itzXYKK860gItrdfipiEHc5EW39QD/wka/tx0ZC4PQHbS66SYb+4kFJNDePpnJLo
WSESiCpf+94Gq2BFLnenDvVsgYMMcYUBH10GE6dHsq50ZogZLxxSBJT3fkLmFaFw
ffcyIFdidnLmNuX6n95jbkSBKVAkoXgvlDbljU6gPHxCgYcCxzweGnbF62hAUBFF
rvTjmK8lx0cD8lYZL/DI4A3DHITVui2eRWo56hdmak8CBX4kilcI31jyY3Mz0JAP
Mh+F5bMKeI5RLhVj6LpmP/j97pR850nDlrJ6JVCK4fkOO1C5Z2znja1Qfzq86RIy
t63+O4y1Heyc+7lk5jfArKu/AOkQr1FTBlQr3L/MOXPaX6GbogOTSrNly6BTQyRw
i38FT9VE2f8jQR2mHwJbiTcvudWJva6ddWON5q8ZqICzPbWdYnyow9aGflsBGQVD
kMc7Qr3+ioLo37VXczkVLKe5Wy5iOigpILjX9d958lA+E9KhhnNTVWJo2mt4p2cs
7+vR4Wm89Jjj7d2ASdvoxzDntWVA5FlZVNLe4WfIdyuqggse7Q2LSXaRr1uSr3I/
0Jli473yG98mvXfbrL0qN5T+0nW4yYxjPkXeQF2fo1mJX+9xCcEWqaC0ZHjw13Km
O3FyYpMKtAQU7n6L56Pfs3tdRN6b7RDzmj+ihftXIRirawXjitQhk9YSEP6OYD4Y
wPmZtV7afY8cJqTCy3D1GQZ0TGw6HXP6QuUqjlSOOvA0V6m+a48edEYNnN3rsCjJ
+zhpNViVOqXHURQjZdzO+Jeod4OypIDH8GH8if14DDMC08PYFyrR4WGwiHXLBr0X
I1MGxft7fuLP8ymA7p2Or46UhZXtpQIlca0TCAW0dlCJGXYRsx/rI7fCA0FYfO/k
khLL7YbuWkYM4VrPHTl2v+emBkxNKSEswbwxeParI8v942+tWivql6DySRQ9eHca
zmxQLoKlviOlD6yMd3OzmgdNpKthM4Hks9UTUA78InIdL1LHQ3w03ZpNERQnYzP7
JFJn2PCRp4lhPfI9OfULIDrUVASj7vIbYJl3zse9sJSSfO5mFH6yi0On98H5NbfT
8b9YtfCdOfEircPAjmNl0Pt2xtZzSC3N76gS9sW/C2k4OzbuRnGej9Do76meh2V1
7uMbYkKSbGb1tFLdCy3309/Hkc+cP2znFSrIJ2qt3rJmgxoM3mr+EDv4t7R2FfDK
lT/wL+dxy8svj/jBeTey9ouAW9MPGUlv27xG3lswzVDX7KbmhYzIxrCFXLOliKSc
jr45UWOPqcjGcFUDpRfvDk2oWIEq051Mc2v3W7UO2ZZNoRofwjHLqjV/eDM4IVJD
k5UvLBbHwss0HJq498Hv8cNDOW5IVJIXJhu2dYSxQyBk2jtGnQffc9IiCvMieTTB
4thc+AbAp7Pycm/p20648A2EcJgZZuzLkaFBiJnF3Ogd48vlGCRRPXMarGNqcX7+
aePpbzkXyhA1JE8qJ+dTDTYHf8WCCroBKPgBKgBdV8R5KjJ8uOCOLYEl/fPOjCZq
ihtcGeYDuGTjb3nitLCfmpTdZFGrYES95InxogFvcFKuJOoIplEkMKC+E5L5KtQ0
x5vYSn6ByPsX0NkTRXzswkuNkGAXTEv18rb2Mr4iGoj8Tzm2UlJrSdqmnmDfTfsu
1xXgh6MVxI3z2M5V9vIrstoCbymFqIZkfDop3CC667zHxsQOnfCV8lvr8LU/3R6R
aMczoG7xFGXnRsiGizyy6CBXS1+9VaG4Gra4OH7PrdmaG2NKghnZpHtDvzsXFiXu
urlop3rmFISADGrv7k/seTWZ/8oehkZUp9L+SGlfTYE9bpTueWKte43UZCsGP9fV
b8znXNaVcmfpzbHyigpc375K3b8NzT0GDKZDGRe3kq2pEOw9lcYnskguMtZgAuvz
vkJpsckq9NCHLMlzWrbBQc94PoHpBCKzNI+V9xIB84QZw+auVoxQw047d4tUQ+02
eW6Tw89ZNC28nwYAKw225GumDLs2yxpa/XT6C+7BsFePXAjUyPJqbOGw6nCc7d2+
/17WBuK4sb4nFH3x9QHFEMVey3SZx//vvSSm1LOA+mfuJAhSaTxoteb2C0iI+gnQ
VEl3tGsttbLCOPsHoQSC8bJE6vf8cBDgseexyaBczr4eUNuTgMzP0Khs/k/NnCOC
YNHpk3TRfoHdMHPiD6CyOL2XCU+ZSkj72S0ARm+puML33o8mDOibwkmRD5CqfNLh
4m91LDkMmWGX8wHlp7LLfy/WTt+UIjoKvB2KbM/StcNK89ONRIinTQ9SNKEVJhxF
6uqPAIbC+bWp1A9q8uuhXYl7j0uuiEeM96qXtIqzY2TLRf3CbviX+HPgn61t5HLH
yfBhgLQ51hMyy+WEXJhuXom0o0AcpEDeAWy2M/D7Y0t092PeEgLEODmSBPUrJ1MG
hz/b56xnIEOf2bZDHPYDDAMbOQJXCKGIXe3DzK9k68QLgdatxE9LgN5UkgFwuP0F
G/hpGx6Zlv2fdtx6XqlCMvLN1GJNqXI/XnLkeyaOqdWMG6xKWJYBNV3dJVtkSrL7
9twi0Z2vVywyhfiyBA+zvlvF7jd88mLNchNsHNTsh/y7MfYhKxAu3QfxPmQAvrVP
LZdeYWZQ2Ua90D8Zoh1S3zw8FxHz9vrnNZCGV4focIsgD2uow7dkS3j/JSQwXQ/+
aMee9P28FUBQVCj1n3qiDsDGsNS5cecRE5LSCA4a4HHhBfvJXQuZgm3D81RBQHWs
QdaWvZ4IDlb/vLpQukb2F67wpLxGITSBjexf9cseCVsmAiuLBM5qmEeUSVpN6TXP
53zk7Py8rdg6nqf5uDnRgRSW0P3n5DxccU+wkn8N1tO9rPetQ1fN3cKyOGlUsV1V
fPuhOYE+XpxpirdTV6WVnrV2wult6x9d2gPOMGZTPYJnJuc2Rt4GjVW6ykarWEzn
4dpiTQ8tZlakhZgZx+n3fI9aFlOME/SBjqJHOrLlEygoSLcMWpfhOU7xi0MySDl2
oIOg9VLhvYi7IrHXxa/acfTUaAiW+cZKjAjpEETgv6kOaPPoQrBhUCYMYCG2eS+X
5RxoC4jDP0hN9GN37KkCwmMG8NUnys0ca6lrYyYP8LyWsdDvVOUrHdYUo3SaygGY
/pIV023iZd3Uzxw/zeqGSBicp+if39bkmoHx9eMo5hRB3JxRFXDlYpvdJPwk+UCj
b8ROs9W0CzAI+JinJKscvKxlVzFI7/rnRbVIIuzlK/nmxHjNnUrOEMwKwLvKF1gh
zkfpaWMp2eA2F/FNTsM3rWFxh6XN8OZ7KHeKtwU/41HJ3lmq0hvT0dxE/pWKLmix
30myqvUveownFzLe1HW1GJu4urHsZqFRe1LfcJolpRU/Az3cD5i+6MZ46J+AyPBf
IjSnwlEljbdkLJu4BewnUk0qdlgJYfrbsliLXPuOH6dPG+A9IlVkD0y2Rkzi5k0y
m6LTDEurrXhjxHoc9inAWW79MY9v18fOmkG7IpWwWbWGgLjWPLsP9Q0MNb4tDv8m
e93KYrkmYkpZVKxIbdxFbwWgWXhuwocIIv5kGEMVM7rzeYOEEebgah+SNi8FWxRJ
1d2jnuHq3hCn8TXX4/75BSwp+WFV2yYrz70W5Bc+vTerDmsBEa1kBKxygEdvvYFy
/YT6LzAHGd6sE0ItjrfPiN6Mwl8R6wybYubbPbgQIkSjDBbhBprH1N5hue6KqqjA
uU7DBjhiyvrHYT22TuYaycQSLC8ovGpWduu5n9gex6zv7NjeEV0+XsaNl895IpwH
MK4c5qFc1VvakO3qzUb/gFIwuGuauvz1TYEU2x1SFqmjHQ4LgelDRswdYeIfKKtO
fsl9fFhZC7HE/PRRgWCRFt8+s1Hn1Yb7UBi3MnPJ6IH21xsOOc/zXoZiqsMz7rT0
69HhH6omhHUiwIMkspThavAp3i7H7ZVkVXQae8wGFQLl1zi7uUAMoMkv3vY6YnaP
w3n+kMHu51zzwrQGxGLthAHooyqvc9Md8D97v6MzMG/SWzqRH04nlWyajQJtWMUB
aQlCzB09KvmcBZ1/+A2PeNtw8gU0y89mPG1m4BmifLcGD/1q697Rp1oxCrTy/zdE
SiEKMEEM3voaltnK51zHbDmGFEJa58MwqXhHGOqoVD6ZRy2eQnDec7RSeE4HWLb0
vKULPwdDO31MsU8e34l+/BoUzZTv7N1nim3ZIvEbLj5PhPAMkmliOgloUk79aR9Z
uZ3WCwSnl593j0pWj4/6PNg7j0h9RKYvBYm54NjZWb/eicNBHt7xdNcQ7Zg0RLts
6ByEH9jOk8oDyVRg6Vl3+F8AGeAjaQpEj2oxLydHtL3Zfxk5nmjKrsrbM8+qgyu3
TtpGDMJoUqzEeRBSILV1KxI/abvLAS07UJxZRHEQpq+EN4hp/P0/aTWojuLdcsb2
LarMy6tc0BXo8nqAE1xRzWlvZNHZdBBn02lKywnAwus50mK/XE8sXiBE79oyQLzx
cENDNeVsedSUwX+x/XgQjTd0rGqApIquISRDp42fTiHNISDp0HIac24DwHarWSPt
xbZqrbhh82yHHI6fbwNa4o6fyT7ZU/9NOqW/2fcNZ7JmyepGJfP+HbmyfNsey9Ji
vCIU9a6cgG5cMi3eeYIKYMJXpHRqM0gC3hkM6fAbO9iCyJuCOmY8uRcJNzUmvhx1
KlNa5Xr2f7M0XRfbF8oBOMrVGU9NztxGDYLmeNX2NA6OsYmJ+R1FJUW48r+u0Uyb
IwuTsbkW5CKFM1UNdKSOvKYrRT0jXCPkYTusnPZjxE3ogSse9YOiSawPyD016slP
nGjNABMaL6hSiBDOPk1wrg3Luco5VlgrOzhxfjMNPb9BeZUfdzxfV2h2mOF8biv+
Q+nl/ZywJk4pvjmBBwhVajLCPqV4ZT32SbeYGo4rYd8WNPqDdsMkGJrxOFWsZcjD
RJW5RZGVYPg3sVxabB+gUnsAimKa+3NjNWX9sfPkCNg82K913YSCmXU6szGFscbI
AmYjG2GblMgVoTtj+2ssX77LxB0jx6/JacamNFD3jt9PC3sbRXzD96E2djkuehtj
sFFdhrU/yEwBTLC27H2T1/hQ/HvafX2c2rpM2OhnjqYmaVMKOkA3D2/9g9ic4oHb
TVmNo3nCCzCtOqGUNqJCJaENOVO33NpX8YLj1IbUT2IQq13BO9BPzs3KgjDJc0B5
dKX9GEJxLHpY2KKhFOMZQCwm8YgtuB78UOd8tL2GhVR26JPbRKffLClK1KzYlhJG
x20FCzmLtw67LFbEfb1mVftTA0ht/BqKyrUVAJfOl5F2U4IeXGqGxzUCqMR6nO+F
iOXv71jh39Y1nafP2LajkPi88MJ7bPINx89klOtiD8cXUl68aBvJjOmqvDxIh1Zj
VkKfrOtw0FYSNUw4/JPltG1uvS99pa07rzyzU/DauHB/2E8hE2QaqKcfwb0jvafs
fmOV7it6D3op/KfgXmIeWdtmql2H7C39oNCTac57SXMoz2SwMXkk2zVbnfZtckIw
ZICfQvHuS8R9gk9L5jDTPBGrMbfpG1Bia8RH7CFqM19xyhzTx+Yg4d2JHNd0WTK1
iCCmkiMI+oN6yZYjcNHPKvGupzJPg5oYxlbEjwzrUVcW1tKMCS36s76ogAYjk7zR
JW2qdyWKE1TaOPSjJvQ986EJgHqBjvG4WH/TEITz6bKgmZGNNfOKsKNtT0u365wo
YdHoy4m0bHefvm+ydNv2EcbZ4AOYMISL4FMfLD1ikXJPW5p671h2abcuq8z9DaAr
QPTPo0NjxdQo1X/hTy42E6Q+aA28LW8phFNGp79F6aG4hhVRANJWslmkKSxRs/S7
uOve6sYW9lCVvNdUgN++iRsNXsHQyoWxW6hb5t7jV6en2VeZEF9kNx14Zj1NH9Ua
crTRvKkqVY/Dl2Tyq7547bb2DSHkEH4H+l/rimsZpVrlIAHxp9WctNlyiCj3Fx1e
wQNqEeACiaZV1jd3xsg0c3JM7VyJ5qWCpySSkm2QhlWbVDCIZJf1TkLkpPhM2i5u
7fFD+hNqCxNzWnXQg2zOhg92WcCmq/RWi3NlPXjFCn1rwM4EuRew16VoERN2J0rg
sPBqYk5kE4JNioLBwIwTaxeJG+gLOWnJ/lcK59xqXqdI0VvL+WeqV+oDTBcz1bnz
5WF+pHOtbLTyHVB2qzqG2HZ5Y8sbf00bnDvRA0XxsiX5YTFeKDmnr+MADhz8zwMb
MDWYMDafagM/GcXSKhCaAWWXNefj4ND7ktFTWZo/Ll+Bv9rtcoNCFiL+UEDZ/aHQ
LTEVV/QhPJqPvmewPj4RfyJW3qCo9oDHEaK0LJhqUruR4LpT5m0zRJ+1Im/gVQUM
o8qlesEsYOF4I4vkhPsI7kQi5LhNzdJOF17wzHtDwzkcbs57bGfufDgm1xrVDIy7
uFWNngrusPgK12kJyUNIdzQXnesBbzYLFHmbW3QeUAM2359NhLFcgRUT62ZaVwfj
C7ZpbdytgHh8CAEKbbUzDGTt6m2fUR7x5IgSXD8HHTQdUZ132hBYdB89qwEQSlk4
+F8xFgcyPytMfIynEvq29JJcBx95ORS6Eif8iLM9jIP7wLeJrsIRPlH82rOyjOd9
iz9c2yGWOY/eGmkvxIze0umh8id5KsZtHTLAMd67HG7H0pWWmYo1LVdpmVDyNoAk
QV386GRVPjW/rREHLsKo2WaWCAOvrQfA8tbRptODsGRhWESi8UmVPnSkMcSHcYtG
glSprggwptxi2NjemiTZm7+ko+o88ZhX0ZL0HP9o5OXxxgSVn3v7wv1rk5Giw0Tr
eAR580315O4AZqV9jBTaai4DJXXWfcxW4pC2SoBqOd1I7Bp0mG7YfKHG98YYrB2r
8wC7i7EfA5Pnb3eRrhmMThR0REdt0fcBBCCj0jBYwTNRBuPb4+4waUYQjl3od/Qe
V0z/RLsy+NEZCFugLZVnmTeuW7fm4BEWfIbcjOi/yMAHpn1mtwuiJL0J+8DEGnvb
FM+LUCt/vTfhng/8nJzv6Qr5MdVbQbKi70FWomxKiiGevajyT8EqEEGDbEptqwTf
Jx4fvuAJP082Kns4hsXCur/xq2u4UM+DqrCqn/wREglFwMUhYbFdMTJbScMA4CxH
e38gEV59K/K9dLG1eU7pQdaKZQYIDsbHlRupl8wd7v54jdCqCEhaQhSibDqyUGyh
S7Q4+Mx4xEm+xogIdDLoMUTPIBHeKd1NKN5ayWaw90hwYu3CwuoI0IbPvfHP2cg8
/aubTE6Qq4B7+oc36lWTxeFtYS4gW4H+c5DNG8d0u4PTFT9eS/UNp+nKA/V3u1un
hpI52tOhMrCvAEf4UIEsS5Qe6l28UWeM0XZ13JjKHWifWoQ0i8asIEzze7o3clsr
UL9A2JlcePRG6P7rloOlOlCEHmaRm36kOIcflHNdz4cM23r/ovFfTM01S783SVII
q5kHQdUsEG4YrYeWsIuNrUqDXAbg3t15mdT7uQB/pUqKrJryabgcvCrjztmXLrWD
QdliD2VQSk72A+AQ0642MHcpj+bP0Bj17f+r2CCiVeecwwUZsCIJFkh6i4GAupdb
tOZ5KdLgB6USkmVs4srWDDF4q98QTEMkbRXfAhF/BlnJyoFS0pr2smh6UgYUkRsF
Ajk2VXjkX0IPNiqCoehRq2BGTyxtpFL+XCUBHP2K0N4WiSme2eHEvm/FX9pg0CRk
m8TYsRD6bEU/+7M7HmI92dIMhnW9uw1BgBjaEZ7oGr94plK3ETHJ0QKrx8l1ztdJ
LHzFr2uEnuYF0cVh37ME1rkZEBrJSpmeo2oZDuzN/DHCWD6GzC2JrJFZaMubqP3M
tJGyAMhvgeZ1XyF/MV77isLqjCzPH3ufYD9NiV+TI5sfQBZRWT5ImMGUEQH8yrhd
vt71OQHlFNoTifNxFpON/DX3Iu1CxkqDJwAg0fOOke5lRo/5hNBs64NhpQs7/ZaS
E2l8SSOylqeP4AEOweoW59EY6qqCV0KfrPkBIin1tthzAd49yYIH54xWUpcCMn35
ZWxfQ8Zt58PLxlLRdQoAsIyaMH19manHgEoG0Sq7KsSEPn4xUa+LVjwszlLsL64J
XzSSi0bzJ15GcmZvvgNPt1td+7B6fxh5YZTH5ASp3+fGDp47pI4iG+S3nSErOder
9T3pXNRuxIsGYf1ry0j7ArUf7Wg1bdREtRWlD1nyElFvAW7IviZp4xZb/9iHcN3f
eT0HAkYIYxAcRdjccFt+Ok//iAh44nSoSzjzFTLfLRKgQzHtxS3ciMkxhzsDh76Y
CGmr6uP1XbXdOBEpfrV18lkC+aqYkO2Ez6AScckMVNoLOhcGlztDcGQvKBuej69M
NSqos69IXzxWqLkc6mrf4uZG/zqjgIeuddBR8X6ZEgWTj9Vcdm7BNwk3t6jKhc/3
LI075JX9SHl2ywCJh8agHZuQqwhtLvee9isG/02UX+hJzShBvIV1/TsdoqwdIpsU
CtHpRVj9IohKzEgNKP0jSb6ju4duZ+uGI541e42fuQaES1EZ8HUfYzo36ihbvWZ5
qpshY0O6fyqcvjZQL92RRCacXdsYdwewLV4Ns5KCmdVdM1b+1to9FsJHZbcdq2+2
3VQsvN7iOqX+E5aRbHhXbil0bPBPFY+/CtMt6T6Qpq1Jd7RrgwD3oU+TS27qXD49
kyg5Fj+p7bTt562S5KdhxMNFrWj0f1yumhaO7zgMYxlbmMdjx3OIyYafkmOmnp6S
D9/CA9o5jgVCJ0V78e2Eh8JF4oXsr0hoyfFKIcL8sxzjQ00/WeWb+FIzYXEWwcaN
OrtpBxhecSaYxuiHXHzUE4Jqf8iodqQ//ndVrFcEZCLXrow9uipI9djmQsODWMD4
Sq0lHy+oH1zaleTBYRbcb4lLw/qfNQXjBjYBZvYk74CDVWlvSbHELqPapbKONS2A
rJlAni2HgovugkIproeHsLd8RUudZtg9urVyrne+NSE0iKvCmY0tWGWx8yaVg2eU
YVIO1Wa6XAtcajWXsHpIhyCypl/7e18amLronsX4YavPQ6CNX1BgjPxwNsrQsEZp
ZibhQchoEJ6g2QcQLzzMbJ76bkWPxkJ7+f9ruwWSuDflPrKFyTfowEfTh1H+CBym
OFrlhJNJpQBS1RWKLwTsy+jjWduFTK2Q/kMxYnij3aoAMrwLXEPvW316WTcT9BpF
3VhoxfAAA6eMK2v3nnhPnTp47PbmTkqBn7A/8rljbjxG5pkZnNXsNKCsOfFFNcPq
UegV0YqjK9GjcxP9O/LJ2WIVrL9RVapez6xZl0WDjl+5jPsihHqp8kY973KRhhA6
W7XWeNdAzQvkSWLVVtKRPfJbqOxPMAtK/uyOVaUQrML4KwFGF11Ugdh3wNHSkSME
68XT3WU7CvC5lrcdOuXTEUqZzKLCTuY706tAF+k9ydSrnVKzQsHTChGF8Ig4cjqr
OfTnZFQTXYeKSR7tj3nj/IA4bMyqJzwonwbCiRki/gvPyKPsx5IDCSv765hXOU/u
Bf/XFRupgJe94+OJ/c6b/UbQfI30z77h+gM9/WguzjZb08ndoz9Ukd4rhgFxEefD
erL3hrOOF8QKkKchp1eHJsqq6kZi1RpZG4lqhV3lX5FrhJooXxv86wGN1VUP62Vn
HpRPbXRfIO69yrs/jfgsdWgTNyDgZeRYL0HN5rSFLR/8NFtJPhZChD3Vs0ttulhI
ABSdbHx/teeFrVg7WUpNOnXLPNrvcZ+HGwI0lPRa6QbZ0nRVcPG2KN3tZlk8wpdi
rc5jC/CYJi0shZUJXIpo6iKv8ymTeLVWNXETjF1WK3I6xbFUqbWp+vu/xKgyVp9O
6FlVYJOFKY/aiuRUnzBG6pPEYsY3XfZ5WItiNaUQXosPo+MTs3RdgtN8/1GNY+/F
btpv47Ba4MWGH71ZJZOWTbnOoMliVhmjukqDDjY2GTlIvoOhVjBNUsSMpdbbCjca
OaqRwRZ9hsSt317lwYRQxzJkf27b04EoHyfQNzCzCCBhFJHTij3doj2dPTFCJ0Jt
C4NYoD4hnpxk92v2fhAPoUMi07vEu7lb1aHF0xyn+dJXBz+bOU9DwnRfPWzD1zkx
JKNANLp246PmLQn5HbABgZcA/NhG+jnVpP9nxkC+CrqWg1uJ0P5L7eQ7m3TMfU2J
OeNb2DxfWDn2eUes3ITY2JwDMH8gJD6Qa2H1nc0a4WCOiu95ZJnC6ztrEQEsqwSo
36abdNZFZKs9XOZRbQ7eW3Y/q1Qxi1jokoWh4ZTtB8TH5b6uBfpDNyOZljNzXlAQ
iVJUD2Uy4uIwLWdex0CzfASpo39t1gf6muzRsoeOGzutMEWonZQAF64Mf9cjZX7g
gnGT1m/ZLUuVshc8680wqp0oi2oqmW0wAhi3E9fvN0eP4ZsUMDKXjHnPcWRx0Jq8
cFaI6PX1qwmdDSHjcDzg+IUpJUTAh0FfOO/ycv4D6mscQ7bJEJvxvNP6UzIIYjNk
jGYslRNKB+LlH8wJNCfArWGJDzoxmsLd4fMquQwXU20x73kCGrvtJlpwdBYfLsiT
oiAB4r5UA89fLsavUdDagugFtmqUf3y/InwUXzmwlM+gb5gTaWc2Lfj1d9n5Vtu/
n9lzYWq3aiby6sS/ibYnggZo5Mul0tzQiWamrGPR6ZISJtWhdn8fpThfq0goBE4y
q/J4EcUvqF8I0Qz4Jdq6VAFiUMFlQ8Ectia+RA/ObK5BqfJ0YxYZd8qZ7gwNeu4K
YYd/5lM1QJSFySa/LrcNybRZA5j7mqs7Rfh2kVOMuUfVQ4qk3gpUaC6Q3X/ddsKM
Ga2kqurqYWvrR13Sq04W/RTaSMS6muPR/p95vEHZfXZ9vU+nGn8VzffrNGq6Yhnp
pqwcVNL7YIEtt7z5XAUKZ9Z8JvWs3mtsJkv8bAizYGpglQOi1WWgH4x4C17Byykx
ZoXpZlhXYdy4mVylW8pleoIddwr4k28zvu49LY4Z/d/UTsKwpmE0AHd6nC3We+Py
pd32p8WIAIGqk34SQA5943LAJNUSahEwKx+54UMBkScd7fmiAI5iSyWJPSuN9Z/Z
I0YXGLwwuQXFPmLfjWCjkMdWSUI279AFi/GfQ5hZf0snMUYnrGYgRbAa0bimlWce
k4wu/hLLBAlYd3hLe8eicXnL1VjLschwi6O1dTRYl075RkoHyUSGCTMcL87ILmqN
vENHSF767M6ew+yULUOyMMF+60kZsOvPnlO1qhYuVQS9Udj3I+YLQKzolIhcTZ9Q
uPu8+YF4wmySI4OrIp1h+IlVv9geV6Jb3mrr4zNJOMwJBACBOP77oqOofCW0RagJ
DwosTMCLZhr/D4iLvbPfIHzWcn7FJLPHxf704natyjJzJNJPRjtINvp3EMbiyYPB
1DonqgYh9xcP+QKRTblBgbBx/IHxxT1htdh9e3feUB2x+AXgmSOIr6zXVsvMXpdh
uBpaAe+csl5MceEt5hqV6gF3noIKtyMJPwvTFWx0MyvLenvlH13/tKuQ9VWYVVuE
ryk5DDs29QlBCuvwNEnkHe/SILs8Ut0ch3W0DRD4aAshmb9R2OT4oNcoCgsSuNfR
0AwgCxTn7OkeFkc5jbXfjDpv4pr9KDYNN78/SNll1nyUADHBAipym0ldKWpDeqRQ
8ouQbuKf+mUrx3nzlmY6Glk8taNVYy3wesriMDzVUDOor2T7KpWas7L1s/meXzsX
IzoLIzYoRKTZjtfDO4bFGo8zs+YBOY7s6Nx3boYfuhcU7m7h2kxhHIRnSzl5FmJD
XcpwbO1KFrQM2nutN7fFRrW+ZDR7Qw57gPoNIqqV0byqlk/3VoIgY5yuaR7CYHcz
kwcM4Mztqh6sCaCb8TdTG2Tmiwf4Yo2wLGMp+eO6OfzZ8O07nopnk6wa9QUHgQWe
AmM3MohLrpsmsAPtAqb59UQQTB7xfJYLlzwAz5vwe24X1rtDnwID5rhd9U1kDi2t
6xn1B09ZDZMId+u+Y+xCAROcnkIhu4bRJPE1KHiOowRO2bD34tHok4ZNVtrHq2xj
F30REMcvriEvmBtaOC432t3li9qimull7sVWjoXNU0Iu79BnS80hoj5UNX+oIV86
MapqCI/GWLBbJc8EO8qnrP4bTcDNRQjcWaTzCbZYhxz2eIVjiB3c8iTDXGUkFI6S
oHHOhhoYTk56m4PNMBLBUC+grzoLflpXUwIOsB0DBrPhQQGi6r4wUOxTP/BPrEyy
+jERJXO+CXupqV5sdy1gcdPjT/R6fPVuaNCCL+pzRbZCZnmOmZkYzRMnchwpfWsN
JLtYCaa7tOSkvZNG4QJUnWBYTEV77oVjHsUabYiky3H8iLIBUiRYMjYEWnKkLkeN
vGlOw2xQovHuaAM2GCqyGVKaNZi2faGC5yW5QOg7H/OrDvYuji2fuQbnXIRF4A9S
53YS4bFX5QLRHZk7XS1OheH9QWqZs4PCDg+pCob2uVmMbNU2XqXayV0XvAn+IO0H
pCpd3D6RhklonR/O4l6E/euD1waUmnF2bFrTVb1FxzOPXetlaqjCnUu73bgQjRGw
tK9ra/kLtJvpcxkzcIKQ9hIBeXflH3iBbFScrtU1BVB7BuOdMVfxR+Phm9AajadM
3+cMkYbaZbimDLyEDdZWuLoRBo/SwaluSG+p6JnCtwBiTUXWfKbmZSrzkCwkeu4y
5w5dNZHAUFuCvK1NyRbbIRjjw5K76jz94mOCHOLgQCs=
`protect end_protected