-- 
-- This file was automatically processed for release on GitHub
-- All comments were removed and this header was added
-- 
-- 
-- (c) 2025 Copyright National Instruments Corporation
-- 
-- SPDX-License-Identifier: MIT
-- 
-- 

























package PkgBaRegPortConfig is

  
  
  

  
  
  constant kBaRegPortAddressWidthConfig : natural := 28;
  constant kBaRegPortDataWidthConfig    : natural := 64;

end PkgBaRegPortConfig;