`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2864 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMWORzZC7bo0toZS2Zods6Xs
yljw+BvqICQb54hGe2JGpN918fPsJVIveSUetI1VMplMqnd9E2G7yni8di45/T69
CM8lHvWZ8gPdCtD0w0v+QL8nPPDMpXyhEacd5mYV4oV0drRZK9/k7y01o9GiLnYg
oELXL0PrkXsVwLV5Dg2LBQj1idHhQM4o+6p6yYXFW6BcCtQj+iP9JFBbl71D9CFn
kZg7zcFd/9oNnGn31x8jOlzKrrW61FaYyey7Pbc+YTP4LAATJBUrIcqkEn9PaPTD
BOrOH3d9Yyq5lZ2SMjKK+W3KrAWi29qDgKjMa6m9lvv3dRyD51OQHlSe7EByY2sJ
oM2sndxD0mD5kGz8jUkQMsnqUboJ+0m0XmkIb1/St7DUKMDBDeUmaIx34PFUgidA
FmbJPZG/oJeLcaWOCvbskxQyatDxIbLIRQtk1/HPI7cvo7C/bPk+d4kVLwW65l14
1Lyvx65V+3YXwj6l7NGTSEoYil4h78+KebKRAEUG/nbf1FNZ20pvAQ5qkUytbqY3
qtA/p5ZZrhwvm2QWFpcrZQYqBeiIrQnpkYl10h5x+oVgFiHveSX3UEZdlDqiflgH
xBYbaZc48U6ENKI9SvuFXDY2q5nEIb+bJGBrQTwSCv0i+zGCrNQCgng+P3CfvKRO
pItB4vSUEsazJzeEtah/mhIrn/SMyw4XtUPCRPozKDC0h2n6rxlnahQKVL5TLjWd
9cW96jDd0b+XZWPiubhrAuLDMR04EKhziXQk5j3tyRUGS6wOgIVK01QfvbePmPrt
xFhOmIgw/+34wDPBi4kWtOnMlJaSN8l6gwvm2njsfZIOx+fqe0thQtBhb6vQtXyi
4acriEJFeYsEGYta7OZVuxu3fn8/3a6WAAWld5x91B9JToVnnDAyB1mqHWLi8rDW
78axARzgUHc3u9Fx1qDc+DiA38+K4+jNhKRENrUctbn5OAlDmS501M/t/7mP4XIc
Hg1NPDwEjU7AhOnhdw6wBz6Ptn74A/73fDtu1Xgu6dHmtnf3nbwPR8QzXozhUw0Y
Ue/Tz82bZ4hjUxCDmCjtIe64awgNIP8bomnAV9wTyYymFks+S7tKMe+vSek7MSBK
3mukJ3pwx4CS0hMSssFlPql2MLUTIl90/96lLoMo9c2yRddYTRqtfHSe2d4IGNqR
FIuODx3xfBkD8zUIk8BH1G8est9sRgljjdmIRaMUl8sUQVC6i3rVPvEDfbiHQ4aR
m/BIE0PzIHdVrt6fjfoxLBj4gvhqjie27YXfIuO0WR2FVlQDaIyYOJYC2u/wnke4
VDU6nPdQpQ8rLWQoq3n5g6qiNkUGqxDCsMRFJrg4wsN+gl46+oq9s+s1jKovPH2f
ublU++hhvX7ruAAD9C5yI1hqOM1liZVlIF9s1iDtVQ/AUP7WOTfdffScGTcC75OO
Md2nStsrAS7NKRcSnStRU3Fyt2TXocxn6sXQ3KYC6wlzj8RgWuZk8nu4E9eZT+x5
PtV5hWdRL1sxudyxvcL/usuzOnFirtRVqlmoz498EM596+I81twgm3GbujRzv1kz
HU8xPRwxt3N0D4+oeRr/l4AEmBS0ON6SR7Zz0+MHH9CyX1fBwR9w91vwusdl1746
Virt25l4ToO0FkLBW+zRXgDJi0pPHUOIToMgJZqNXI6ipUI7StR1Ls8BW9hJPnTU
6404no2YpmD/2Q993uWYoBnLCEkb/MQ+g1vmqR+QXUFUa06OQ3rr6QlHmbNUlIrk
PS/1lFYuwYRMt3AICYs8VIvFdI0oE8v4RkavfK9VhkRtFoW5p4FdN60iOfev0d8e
BXQVd3uxMv8nmXeEmqxUh4JjFA1REbezb9oOIfR5MZ1ao8qZt74F3SUIayvyXLrJ
GSA/7uX4SorNpYOIQyVC8ibjGg4mO7brRYqBevkK4bK8Z9wLwhfgMpY+rG/eczUE
n6bX9Tq9KEY0IFRMsjmR8XKtiSSsAXS6fLnD2DLftQw+BpBxomRcfgYDROIVXxoc
4VEPuban+elBV0UuwADFHqgKAqkdSvOC9fL2auBpIETChjFDGeVB9jQ1TCpN6jVl
LP7irT0YfL6ABdnXNIrIQNXwJ5nzSbc8cOf21eSNcdURornavDVnp4N7S8eoiwKz
3fWUoTevuznwBjB4GqjJKK9KYw1omrxU/B7T+ay7wwq5UA0AsB65zWLxUyjf5yQO
ahOuhs9Q9ZQikWutqZ8cB16DL1FJLg0hfw02kcTVgKE31laBOB1BaRk6oR1x2mzO
yWS+2ibeNByf75kcxBrgHQCxDViTjHRQvd3wnSQ7L+QZsm5XHpJ8m8NxoWGePOCy
TtZ/vuJ+pLw3Os4HHm6WFau3hf3bGHqL8bAN3T9lacJhGPOgQlyfE3zM+TAD1Hkk
0jdFCYn7/qyXcceXk3YczqOXgQYZRa9QJJYRpDS8kddHceqJPrgsIecUVSwI1U16
zWpXclh6Kyt5WM8WuCck+76RXMnMJS4RhSUp3fK/MKQzdcuQewyN1vA8suj25amA
OPaEE3wAiX5ymB5hacokiIuTqrST0muYAAqlLMOggfx11wLoFwkRu9orolfit0Jx
ZOXqmlQIa8dH5wzSLMro7NbP2nBun7cJOy1hkRyEHkzJJZqxtiyZGYWUyKcFZPt/
Rx8x7gkoOAmC+voYJ8HlANFJVcsf4rzfr/iUutyAeSBAKf64iEMMsWyuccFWFazt
+Rf/578ZCiVjdefPaue2l1lwRk4pRpt442V+BZbA1HQyp4u3vY1Pqxj5Xbe8cZRe
Y29S7lYhqJV3CXXc4gSNYv4EA25lr9o4wPePCxwuZRPXaAFqoq49H7pTBZWTEWRm
8vFJkTxJga6rLavz1rp59punFRpJOsA1Pv+kF3lssgqMnrkEq/yJIKz7ZXRpUGsO
FsokSDwMo7rFkisyx8QIcJq5lUE9y1nOyibHSHRphH+OgA+vI3SZdvWwglYQZZGG
yhihXrgSLXugbAZt9IwgU1DDwnwLvKd60k+2LzMS3XWifQ2IpzP8uZIdslXdU6Dm
2Yvg7dOSnL1XoH14qVWWN8onKI2qgRR85G3EYQvDejELs2OpLj7hG0+w+rOW4Km4
0aDQR/Jh8feQbqsViFmXpFO2Nfs3+hNgYg2lXnqugPya2hMCRg/F+DRCVqY1Pgf8
bmRpPUbOgstUGAaxrsk1INsWDmCsGvisJxx0jUYbqcLR/pdN4LqCS61871ziisJD
GgAZeFHpe35xRAhRrZvVb9R09fWE7IRJz90rnWgvE23lmskQ8EIA1O4/UkdYshrR
lv62DdWU77o51D49EnXOi6027mUe/l+gzx/ScYe1eMiRz7CwF64qYY2KkJCYSkOx
avGvI0bLHQULEche1YIzpL0opHqT5SIdAlR0b7wpvWcR4GzxrlgsNgLPj1zVcgV8
5QXCCswiZbfVLCjXJ49lokjy4flbK8bWmxc+lsGQPYawCRuFprOaLUvSg3BuAyw0
mTcKu0BXPrPWuyDGg/k44p3lsqkYc24GHuVsCQKluR8YjrGKUsjrb2Ab0O9szV6y
Vs31vJqILVh66fDucveeCVGjcDPRlNhhnA4sZZjYY/IwDHIpYva3sKPwSJ0yHADF
0/WblwIZMuYMi9k+SftUobJlEzv7ZJdBikSOO820DEhHk6ub3j1bUpndgo3XLfPw
w9VpaQn8LqmQ0E7SngyrFTusp9+vj4GJyRE/vRasWkI=
`protect end_protected