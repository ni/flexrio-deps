`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 37808 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
UPwNTJpYF6a2TR8YjJWNOmRRQyWejcS4dqBecDS2DcKRN54jub/HuNzQ8MJsKxVv
vnPd+BpLNRYAWwe2Q/L7obyN7yvLQSUtZDcX4eu5lIE+jmCGzoVeml4pitxphOVK
/iZnY/Eu0HKa1jNC09UKElAgzUqMkWJIYHQS0q5C5Yv6NPczooh60l0YGmnqwwJe
EJKlBl0lsTvtL8JJJM5MJzxVBYAoGyuuZRZNXGtB4fD5A9aGUBoe7+iXCevNHBLZ
8TFFzdUG11nyUZlzuG1l1nWxSYGx0GKoS8/Tac11tuBPRWFSxAc51eyPPvXdnaJb
O/a2SNdpTtapCp79kFh4ur+ffMO5q0NUneYRMIuwiVTDbuOZpCv75SZqxIqNWKUq
3BQBzoeS7AERLK7D/2X/VuVUNi8yjIXFGl4J11LYRkXvGYWyvugpACfchWr3dmrb
GjVwxbEc66rvC+627bh9PSFEpiPOOgAERnkIEEruztqLihichx0y4fz/dOyRGHpc
p3WJTsOIInCHW9hCg3Q2heT5xUquNIklrxN2Cjm+ITkngr8sR/kpkZi2num3sJa0
0VHNr4YoeorXmwuIwbqWlHbBPCdJ4ZPZf+wohujCXDLWk7M04+TXJlcMq6lwJzim
u7MX1tsmoh7ohgEYNZWcRJt+Sar1v95vW1S3L9DmylkGoqB2kMgtTwGADluz+EmZ
2ehD2Z0yGmzMYlsncTGBf9hC+iOUUerYgUNM8Bmd3xHL2IgD8gNIr5ZzouFuKXZr
+W3YIyfsGkSXTa+8zbSUXnpzKxhEi5O5LGWDYHjTaOpUlu71C3YLJQ4xOooRC/iw
f83hj2H0nY3HAs7wdi+OQZQ4X12hx1Au8fFVJHLr02mrnlE+fJ1yYWDvMVmtQpUm
kkNBgw/bW8xBWEHB7PZ/fAnVlGND+PgrGG0a0zuMyr5pvFOO9xu8SNPRaMrv0YBQ
CRACmLUjIljUhK/Gz85Jo0sTRHIw5dGov//HiwScDp3qTBHe5u1345d4vwdU6o2E
uPN0PLmJu11g0TQGuxYeRTE5d3f/8k48G8XTn3sRjZ/g9DYOq5Rvl+rwnOm1dPPZ
E34fbHESQlKTaZSBZkPJsLqSKQkKq/7E1So/BY/Xs9GtrAyl/89L6IrSxBQzFgZf
lcsIYYFtGEfbo0b4AdRTRgsLVbk0lcqYr8zVwfHvH6ZBp4P2u0uzLr9Pfj3nyeel
ApGlz0luZnqV1Xgs8ZzGVXXTUswXAGaT/zyYJBniPCJkIkaST+ESQ+Z8+zzAQytZ
hMxb8PhQR+Jfhuph/TMKS7V2NIVQI4oCkYfUGXetBCBLNdJHb/0ACA4j7cDrur4g
xaftWhMB5w3gt7AxepBcnyfCbKsajNEufvaXjt4TwKMNWfCrZOdhlCD33Q46U83A
QG/uBgWclS5ExHlKUxDVm5u697DyWOsbBmqJKI8d1dcK8cA2OqZp6n+kRweRNvE+
/xEXAb1a7eWrRCtxhB43uED0Jo4hl31VATux+lm3RuhyTJS4Kalli0QPE7kUMvF9
MfuUE/pnqQCQRCKv01DRdbNOXDgVoumYlnTBMedtQuHV6O8HlSxmlFo/7PvgxbAw
rDmqb5Xj0NGzmYTS8iRsE35Ejlp3kmEaV9HnAl/mun0bClAtG8wyjQx0CU8YZqkx
Jv+oaT0lBEYiS+3viENGaYXx/u4c23HsRT/DGdvM+iUKCM35Dc16HU/PIvGiFYPl
2mwkFhBPIlEkUn5FQmlj+bgYe7ID67coIUWCLjlxSy9iWtRAg7FHARehm3NBgV/k
zPzjVT48YEeyQt08U1pFUXDpDvsh00zbY8eAa/8UvlX2GMrkW7ff+QgK9wgArvDQ
550drEC9855sEbU2XKF21cU8RTNvTgN2UnJfsng2QrMyzS87QoaUiALSpJTpNwFF
uJ3X+E1mEZ+EbTmTtqnT0we4g9njHRHSZD9nRnEq//YEhtyS5Swh51DIJDMoCTXC
bVL5+LydvwI/1QHaIZ7FZDcpFahr3O0dnrhz61ky6SUweCCCKopCFKmMywaPtmD8
+jwH6XLVnel/ZiGj3GY9xvZ4mc+g8RYSVP2JcvSkqvHkyDgu5U9Hf7UAsNCepRtc
Qb4XHIsSfwTl1YZIXrm6EirrrpeYtonxu9qpEPBp+U+Si/kiJyDLNk3zQZK/GVgH
SNaquO4pS+KsHo7JXvAwta08mJI3KmbR9gY+4OMsax6DsdWlZSTUXX70rKlHtLwb
8wGGC771DBq5lMuHtuRaidIGE2T6PEXFONgtx5qAv/3UTs9jFBqh4fpt5iRpgGME
137DitMqkXm0LGK4X1EIZwixoIHlxqBzaCKWizz59M/KMBtyPrYyZnfiua1fEe9S
dxA7kVWauB9bKY3qpG5zZKb37Tb0Mw5XeTA1CKtz3rXGghr6zPDM2bfXHAiNBJTw
urcNT12o624ZNqpt5+lhp6QlniMx1+db17UASsxFgKV5wSOeMKrm0iZMuUDbAESd
pdKroaG3Vddx5HNKMO5Ff8lAPQkgCtOV0SsqzlUX1XP/wXKzueeKV23ks4kM30vq
SkQ5autIwTiZghqr3YXL1ajPbGmQ+RqknDtWixWvJAFalS/KkHR8aAU0kA5Gwi5o
TbRAkWXIue2guzLwZLGqFyKqLFq+Iptip00iYN5KkUN2VLz+pXlnNmO2nAafZQOo
xpFY8rewop4A5a5tjmKfLWbrhs/3ELnfslwvvhSlqjYr6N/CP7nrk7XDD6ya05rK
7k9IoYDhPZCTp65RxTQr8s1NGwhYBclq/Yqx/nI8/v86/zUofYBVFCse4uCTTOKf
wCkT1bmXMKLqy+RvqI9Yu2dM8lexpYgWNrViv9lYSyzyvl7DmgYttJ/tDvvf1J8W
kuQlE/k/jhf6fH14AUlDdoXZ+emfR6WA+s+b0R/lJl/Q7XSWO4tSvZ3Zy8ONjo37
hD+B0zIrxhgdoRfJWYikiK8oNTvMGxANzZigE3SINAo8CLySjYqW6CUtwssZUgxz
w+YiGUpFzrrji2MPFRckaeh7GaR0GWSraamGX7bAu/k3FhuvmSCyJ9tjoQtKQYpf
TXnQ/s9Xud7nCl5+KZwydxiqU5NbkAWnRB+cOR2NM8rPhBSj1t23z09yY3FK7tmh
9yz/9tFWSKFVDev+PkSoPWlVbByfrG793+kHC5I8tujWzMhkUQPkicLHij45SM8r
RpXZRJrY0FkZ642PaLq9DbyLQhShWCeBeXSctS57xIm0kd2Y8yaK1q397vewkvx/
Gr6+grHPtSeMtrDLh7DyOQkUvp09Z2ro2kCUvGsCCCioqjDgCOPxBg+v/bLIQhLH
itmNE1RxjgBpTpq5ZgdYdtgC+pJxKY+t/wD0Eo9kWkjyEE0lsqFexDFXPnbUuwlr
13BjdEqwW8Udw9gFT3B7IIhd9ha/hjmFj6R0YCEtv7EANhGPd8oUpiq6OaUbT5Mg
w5XNjklxiXwxr/+odmZrnyw0JLthcJChRMidLrIWPz5XfQNmujaE/Fk+B+a4Dv2T
ZMxuv11JB3FFu6lLBphW6yxBxNNa8RxHMvoHfHMPJvCnrEid1uyT3c3kT9Iu9c9o
pANBs5AQsuHAH2D5f7C+eDgy+nm3/gigSKLVgm56VGzIU3+JypHbFPBtBCAaBBK/
w78atkIBm/k/rCmWyUh4RXAYvpb7mJ+uB/aWOnOUpygOvIgIT7iQ1aBiLqjsGFa3
BicmHWXNlGyuA+Wfgm5meojY2GDdaIBiK4FnhvNsoVgxX0GmPhSdKGmXYPNCPb/M
mceXipez6VnpuTrn02KTPhPgKQwhVqoQ/QoS9JUF2+ACnI7nQr7Zozc8F4FAHdd4
WIAgm0LXT7q7a9zlKiJwnASFjPWmywJaOBx87U06vYhXQv9yP/4cDrRm7zO+saqZ
Y5d3dX8VPEqYqnTGtJ7BCJSMjs9aVgYwsE+9t/C8sF46RqAT75fgfkqd+zcFBMo7
Vy77cD5pV9K5brucHppBaK2MVy8uDUNcUI4kj+htpsJpC4ri6OkqpvmHo9DWEM1g
Mh89HzS2ZB9WzskceshQ5L5RMqrAxwzDS+T0MK6tCHVhsBKYt/IawWyOslnOS5HT
Xatpk10nZojaXtkTZ2gmzlP52MllKixS+SHaAI31IIPCLadkuBW+wR4vsEvdvg6g
3/aCu3YvTbyy0KOPxaupHE9pupnuUwqj92m2XQCx9xFqknjGo50/s1q2H0s2UbLa
gHKTVDKA+ciNWyis6Whz1JfIZkbGG7PYBBZLNPm29JLSn9ix6E26H3F1h6EG13SU
veh3K0UvBUuLlRaBg/VgXs9KYsLMW4JgTAzowOc4DEL5rKoGAj+Fp33BMpm3zO5t
iZf4SmYGBqxKAxsNyUUFFQ1QT+zAaId/1gHlAOnY9uPVgVGlw0p6sjGKASN7h1PZ
THR7Ffo3iLjTqUm9kBasTmiIn75CUkjCYafTTjEtcXDwJipGUcgpKo4Ttixoora2
124NyOru4IVQIawlKedRwdI+dWArBgK1jHf2/juqqw+yPmOpz21cw1URc9z4yhMf
WzOxcsEfcDSPXIroxpxKZbGkgP9Y/g/bOTL9Rc1cFGzfDFnUjEHHFQ8mC1AJaQIz
h3ov6wftKQrbOPiIQ/7o4oTawDJegSvuaizFqnJGtZrVgpbj3HwUHdwytGeSQgK+
EXr7mD8TKc1jviiiD05wZjL4Acr4CNFWfkLYHNaqfj5tmBf6C//NPI5jqtMiafQa
DD7o6xFaMnnLC3H9WwBtOy3ySZhyR7IMcFLnjHZ1t9dbplZpEs1xIUqejftHUE/+
kJngR8VsaLpnb0OuxzChxX9XnzpbwYFDs4efTkgMQ6SHHpah39Iu4GDlQR3sPvkG
4cDwgkhYx+B3XntrqLGrqZrv6uhl4rtrSQ3xPzkyZ5Ib2cxVXFm9Sf6bfe5hH3KT
mQeBJums6sOiIBTpC/uFSDjkhC6QwlL5g8nJWPRMt0gDyAvf92z2TYHRS7JCLSQq
lLXbRhr76poLe/a4FCrWQTE1MrXBCJJ0X2vkZuHNBDKR2V1qQOJ3Kih4rLd9SskU
cVI4aDO6xjiUHklomiJgCRDDaHtf4zmoTKO2qxQjRQtsj5539qC/u5OaRexr7YPg
+jmhOFuiiKVOmjBD4WKLVV30mZxUPTM5EjtiHg/8Hg3+5Yz7u3ojdCgt2sPwGEbf
JuLzn86zxEqHyhooC5e3pORa5eII4O5ZJJqcg2WD95AALV/XnkRjFkvwUM6UX/GV
WtWr7cNMg4yMWvivILpwspcQ31jtliQkJpQfSHMQIHbe4+EtonR75Nh4mwnNZFmB
roWC/NiAIyZB2QDKv8Zj1aLJMC+Pvdy2ptt34ibVD2smDismRJEGVcdjefxkLd2i
CuKJzef+ZBCh696suu2fA2Y7xXtuvny7CFkKUl6hNZwIblIj/6sUabLtDv2RXulu
k9rE091V35uoH5dDGkgaTq9fASyDEfkJC8vTBPkzg9TnYAYNMXZJHMY3JfNMX0GM
PU4TiZv+u1YcCd0+DPP10DNPYgudtxoXs4q3+4Afw++V0ovrGTejR/lkbmMoRbED
OIsETuCX5nwFekUUc29y2jt3Epwo98I+rxSoW+2cXFgDvG3/a7Pcb5oMuOKtg8ox
R6kPRuIUjgcQ7OuOm98mfudyXPG1Y82tAFTCx99XXFn+LOP360/dVSc7HsMy+r1C
6ObJJ/Skq6osPjzT/eOSxW5v7Lp6RDI9KxnNPAdSJcZsL4MCZQpqPkjh6wy7lFf3
YFP3z186+pTFtO7xZcxokvCXRkK03/sqZseVa8eciwz3aKmpdPSOu6npcbxVen41
Nzb55lAovQnMoo+P2sE13mXgLeOjUQBBsLLU5CQwpCa7GrYlbIHziQkwjdSN6yvR
+Uhfbnh0DeCQDzA1ansLbJqOeap6gpgpc1NKn7/xaN4MKxW+MXcqsoF4bxXCa6zH
GhyxTdWpgxiDCjw29TUvog94mkDW4YTXmP5mcm41LsizWvi5CFpEiGchkeI83GLC
wiBNYrPEvLLoWYq971/9NiZ0i4Rag3d5oon7pedNeR9NPLDd7kqlF8HNlctPCg3t
eqUpBYjJTnge4SIQaZrq5IaXhgeyPinpcYD73kx8DFvBvKW3FiSfmu7/9b79bK8o
3wU6BzDcHTF/HVeyFNfOaogszv8f/gMzYPMOiIpqUQrfbO+xOaprGX+VvsxlfGWb
/e0E9wRCfNI6x6I6STjfbfohFX4SW8ET/A051SN/4wE53OrNRIoYl+pVg3chTtxt
qjuCYefA0VRaKe3Ujg6NMnBdUUX4J4bj+P1iA+Ocgi6kBdR6J4UjdRH7kvq7MAPy
rw1UREqOObHyHXerefaxpNwrHD4nUCMZVvrHSVetVre70+NVwP8jZL6+okkRFQmr
vy+mXRUHbxFGHzVlo3K560A1QGbvzNzWzKKOYk7dcNoKe4Zms+UiX2rfNaXkgU5g
BzZykChKq9sbSz2rG5elji2Yf+q21U5+2uYkDreKu8Jf1NoAXLeJ/DXwdlhnojou
4Rvni84W6CjttsL3abxzn+wiSlG3uiiBkSpUtLthXWuQswHs+frXLKQhYqQp5IdT
Nt+TOWilNWw3Ep4ZjrCy5k84HL1gcZt3Jj8y8nTBKaF+l3k6TbZeEBid/qPToojL
LhnxcLEymucE+CB9COabAj5Ao+w0c6K8M2RJoKolP2OxFcKZWyDygFvrtX+KizS9
rSbtnI2BlQJSKFaB0rVdiWJiuAZ6Z2fn4MK6hNfqu3Jlek5r1zBl+s0sPv9AYFKO
ZTY7hc/RRWoOnhTxZRs7Ky0LZBhS6nDVGOrI5bE6SE4C1SzzPY3EnO5YhrJQ08QX
+DRaL/LnfDAyjo+q+EUBuHVa8glW1coFKdylFlSWVTiQOzwMCroRCJ1ymRZ9h7LN
ZUvBgeFvS27EAchMKDaQXvhbURJDwxfMddnNxHlM29YmXZLMpYkDIQhBo1ltCbLY
1qmQLGwIlGJAZ3j4hjKv5tnPdaVkdBeLIrQgUNTablLM4d2YPLHVZ1YUDGw3ADLH
QBuV9OSe+o04dsARhNmVV5UGe4WLFXVQtrmCtMweptlryTq1GamihePHCUd2rLGd
IWNldC753YPrEduu/qeqE5nfe2Kzq1yBa/cEgM3B4umcP8WaFEQaVyKRQ24ovl87
nkehxBQJ+UdA1G8OcnFrSzXqvqxC+3Tyf0UQhaNX0nbesun98bNm+vPyzVPG7Xub
DoolAEMHoYFmM6ODeEalIS/hB8TmPbUSSuVrj9G9CSPZU+O6LOWZ6iLnyKU706M7
Lk/1WNuaMJRCw6SWpqXW4WuZDjGOBNPClt7/XvRuvB3Xg+Vx8ApecpO4wb5zD8nE
5fLJp7oH8EIYHpxOF4TisxDiyoqndHi3i9EWKdc/0wYBlnmT9bmiedBdt7ps0ZvF
WztAwI8M3a+dxOjl9lLyrcdQD73XWIt3fXp/hDT4+zQqpVIkd0wF57794Ps9ar9Y
2iJpP3/kPTgz3KQFfZXWBBocpJbvdUmrgFnq50dTq6w3ha2oOlbCOINBIwDHZaqB
gahOMepA7qX9MVG74mf/yL8AmXeqKciDOVMtyoXLx3Qc/48orU0GnRn+NDVvfcib
0KG3asdu73SPTnepX+75euksw+pTr9PjoklTp+CjiOfQ99E3vqwkLvBtS4ORe1Wy
fcMOKu5+o/JRqBmqBNirMGhje3IyXRzRHkXbmTFXWqjcpL43uesQ4jySlXouZfWY
euGze3qVXy3Mazv9UIQ468RfH1uekCAMwebruRlBDR5LlDpRcGqhA0+ftESwWmWL
JdbDGlUDWC1JG8gi/IK/Z+icuedkdBJ4unNOPFTOUzJEl5ZB9iK0WRDQIstFJjum
THj6KnAbhnsM0vWx7k9OMaPaXSuFQ1/zxF5PaoylYsfYqLt+4O9AArv9pn2E5W1Z
3Df15ElVQNb6gxJCEn/domF997149c4DBhar5AQBIlSIEyz1uagSY3XxZsNICFv1
eegadsLaZ8illgNeY8L8no8n7k+TYdKbfPfgPMvHwmZo/iRoDZaAXCCrdPkNCudl
GsQptKllP5T3FNsKSkAyR2lEzjC+H6AKM6onxzkVXSzuZGq1imUkmwMebFEtaTWO
M47GCDpxKfVt+u6FpeWCchV9C0UXpODEEN4bG7zC9o8vbzH+vQ5MoLFtuC9zwquJ
XSdByu6dSTg7F3NwULCOSw1YCd82sMIv+1pv959dGT6xN+A2qIjuOdPjayh2CvLr
PpkOcHY5mKeMPZvzpru4px8GtRAC4H4xasJ95AI1w5VXjpnkk2evxBXQL59s9j42
o08Qfq/1DYPcG2UadOMa6iopyyG4eFSXxz9BqnhrNe4sntU+KJa7C9YniD0RIIBl
skhwVbC0+nlrFHihVFOjs94E8zuCae2DWoeKrH9T1guEQuyw1LWbPS6FhT+bPSDo
DkLWbrc/aNscdXC9FF07AnS1106q1cowBK0Np0V5pHlrn3yQnHHlb3Uv+eZJotzq
tOpDDmzKLZ+jYxRgQiCelYWGBlSBTYgWTFdP+UDD5ZUvnbTYtZakom3JrPfhdd/s
QJ8X5+TNUrmbA8vfkgpFP0mX52WrXJqo8+8anwD4eb0pFaGVHK/JWugftS27O4nx
a5sS87xSgTRXTEA+usEH03Hf35wRW5sDKHcRvpMRJNA5b8QXZBUHUsiBETkCY1gQ
Ili6VQouBUh/bCN6q0ZZIrzH2tJ9zjPiSgOduVJ023VA2sb5q9VpW/+hvYzhYaBC
lWNPk+v2otRBljhuiLefPIGC75GwQ1IxPRmw37fMpAV1kpiNKLpUC/+B5vksE3fm
GNXM2D8s/IJOOMXX5XDeXnM5Meccq01/1xJ2EWMTEzRJfNBlksaI9aU+Nc3Q4t7U
s6y69VvvLd27D8yxwN/SowHxUxg28EJiyvi1VAcamwCzjZcuMtQrdOGbG7UJucjo
h0aMRKjz5Gh8vOG9vOvoqEof7OImBG1p9dfmWujkXsXUrYNMhq41zcjoSvDrO99t
je6tv0VBgqRTMgskzH0TB48YdQcvJM7294SZunJJKCA1twJ1j7bkQ8K4Gx9/gEcI
Txn5uXQGCs7gmzZZXujLy6P9v1tbm4wOuSTb+3A2IuCX71L9U9NK6vCSaW5hUKRE
03wQB52x9ybgECcwtJNgsYvPbVgx2zvm3FSNcWYdUZVBk/V3fjkpKnAaF1Fnrjkj
ChRGKItTKuKol9eoC1AWepJLjKUQOhDS3jWtbOWkbjkJydkmnVhcVbLYEb+Fd9Bf
hjnHUsge+hFxxK27uYH3PmIY2ayoGKCiEkxGffWICvxlFgiat/ZAiVEt5l5VVKaU
J/rJSxbVOIDFwk5SdrnJqvliPyjB69qv6FxzIznGqkvuqCo4Ckm0nmOykW4Au6hf
8w67oZVyPXZSJLW0P9ct+aKa2pOknSUxZtoqWH10R6hBUMtYehdmKKe/4RUGfQBL
U9uuHuPSSwz3vMwCHwKbTYQ7eEWcy/GeTG12FxTgLyYzWnoQKLYDb+dfT3Y7b3K3
ZSAFKQ2s5HOcKcyUFmR03Xb3BF/Lb6hGptW2nT7xtQvBeewCiKGLnru3npbicaN+
HwM0FPePgKtIcD/CvQ69QeBs86X/2IGBn+RYvXUGAF2RM/MsSMiRrXV4ZQgNcIQl
WEnlMhWztzU27B2ICjvnzY/IKviaRyjwpUz9y4/bHqyCDiicQpGDy3gV+fN13mcK
jz12kBUR446Zo6jcsPlQFENc5b4g8bRvJ2jzwBExzKJKVyqFZ/vvwI6bif8p1Epo
dFlE1Xnnf3uH8EjVWcZFIfXkkoq+eSeXU4PrSuvhMBZVbgbg93GTu5vWpwGtuO92
iejHB3KJ2FvbiwPlEonaODsEAOEXt/5s+y+uWd53a51U74uaN+cRyf9195/JnWcR
4G7JUaC4AjwXj1apa3afMyYn1tlXFM6WioUxu0C8HnS+sz96ueIMNoOWg4uKW2WS
JiTRJ+P6HJllgK68W+40gUzUFNL+MOTQoO4uJI27hXfqE+A1L41yd6CVvIh6ZLD5
oRSgIFBrd9N80s9LGcjrZLrEOv3iu3iF92l9Aq8DYeY0wEZbdOUqlD6qjvOdr6yq
1Zy9sGrXLlNcv6AbonG9DMfpihYUBJ6LyFsEUrVN2793i94dF7iIOKx8NVbtCjFn
l3ynooQ/4nyra183QHf1E35DQ2rgyHDuVfjqoz6GErY0otz61nucl52AfVmxv00V
hUjWQk5h44e4VMPLselOU24zlHfJk1viZjbJrMBLM90vG1I3541Mm8Tf7dauWi/G
ZHpAJP8ZnkJe4PyHcFtOYAf/b50DTwn3HMG+HYAnFx/lX1WyzuN6IfyD05hb1B07
0Dbdps7HSUo1BxvGX10nSubqYNIBfp8aRpMBcaEgUFxacug+cEN3YR9hs7SOOR/+
xkDC865lpykkOEPlt3fAzaZfaIeqM5mDeA8B4PNV8r/xSmUFf122qSMJBa7Q+z+Y
b11LEfuDe2G4MCeVPunS4f9V4Nv5X/L98XYlaZO/mc6pPET5rp6Wyw/4+NPkBKel
/yNqnoP4wDDi3z7gONhojyao4e6kqFV6Sl/gqX/FcmaBmUuRD943AxWOFeFnW5rr
/E8JdbcRuuf00tQkG/5gbxgSkRuwiOCj/tShbAeuBtWKO8xGtMd1tHWSOeXJZ/jn
pCTg9gNFZwttDo36z3YH7DB464OLdrrvgiqu7LkqZjmeyxFg8Md8QkqzVj0RltcH
h2NtPzbg19wAmqVBJQz+za5SnAl4SFBEsBuPX/kjvZQdCXFsv0RWYboUfGmQqXma
lKe5543TzFB5V/j7Pny7IKGNE0l2ZehPtFT9lzkWzDqzOYsisS9XLoO7CCUUbEoZ
TZjcbuCrI2p+4ldbD+8Qxk2Ge7gkI7DG5ipdvKNpDxUo5fqLSPepdMS7YDRJxR9D
bdon+FwudbnrTCP8MQx5qdsiQFOYX2oL6ny8otsJCFO0GwDzsHhaGg68aYCd97RG
PM5zNipL4Ac2IJOvseYSWXZWWVkba213nbQTO7KC/Dov72ZbKPq4wbE2wSxVqlfG
ziH0u1n83Rd2LqJTIAldr5Qx3elFHdOQhI+tDgU1iaqFFibEyqJvIvOp4FlF4sMN
tdqBw2Ab3Jng7HEQAQiIrPCD7Hjat3Nl5iRlXPcNs5o/Ym7tovpF/w3uiWr34zrg
GrY/X+PCwIWL2/7bzgWLheYkJJ18mQK03BNutISG1xqDVcPLgCxY+3ZAo4VtUdRW
yr/9pRMb218t9Dp0gbjnkQg0jxwdipF2j54OdKVdlsRBzdocu6t40vviVM3mE+YA
GOAgRAGwmfwyX5L8LtOWZA/jbYDG18OyjkiLRFOuQlElmWLi6sYkXZorLczXJg00
c8O+45yuZTC9fk/PZDFPHwrB4xRx4wel2ZQqGP2Ua42IFcstntJGpcf5tLlbU5v2
lqlG83mlRkBJx5qe1JXEaqgM7QH6BJtaLeWAG2T6MyXKk1+OPbna7aKLLcmHIKzG
uuKlobUeGQLzcDfrVHx9NBr/QlnHLKNMTA/W7A9qIwKGRLLq6nR/wuOS+uPTMjGb
CS8BD73Y4aKTbUkOR8pdk8JX16VxPothr8dvUnlDCr+ic+/6EL+6jigwno0F1AC1
+66ZsPwjOJ1Q17ptS4Gs5bc3ePFaVhgoNfZoD6Q68JXzn79FOUvNfJCQgleqt7CO
jMoovaxGS/N9ozZBKVRYjqb9lrOLC0k0khwyCSZnzZqo9ll9STfkqg6vuITTLiGa
Y3RiPQwRINYpKJWpJ3v5KjJe0kYldr0HoYRnMBu4sTe3qW96vED43/4eBgHjlX2G
dqsyxK3C0e7xfhmJg5caD/gZHIAxauFyh5GXU2LnMlVo+GcyYKs5PTdGG0/15C7I
rrWTh64y4xAPXbTYYjGb/4hALfl0wHGemv3/Gj0mThGB3V7i7BOIVbWkjF2BFoY3
enPBM9EWgOUGqXJNbvoE1gAEy/kwAAoFFat8U8V67ExOLP5W5xdio3R50t3qA0+l
eq04o233/D8w5Qm1ISmDbkTpGdnGvdlTPVFcuamd9OYVqlmMSGsZIdLcZS1KWaUj
I3wBMZk4R5sBZjAvmLJk0xQcG3PcFM9qZp0MTsRSeSQxZBHz+/x1UFwTRyFQ6E8v
124QTTWtvBx0xT01VoT4xrldLeL1Fok40RC9Mjapf9fC6Nlp2R+WDr2UnVwrZrcM
Xpy7GZNzfYzmnj7Pv8LCB/i2rmvAYJL5ec2/uUP9jqq7+ylobkPh50U4SSZ42kvs
9E43ZjdhxRK1hUzcAnAAMj6DFv+b0OmypoK7nyO9BRXkekXqqsC0gOsjQX79/OU5
/AM3h4hHGtNbFBrYl2FarDikhPTX4qeKL6AAslSj3KtfN3j2hWT8mlPD3wZed14u
EwCYKsbrch+hLABjmHagsiCMYXPOpHu/msfcWVL0f6vYhm4EmsDccvjzhNdp7ls8
os2KeGqYBsGqFh5tGMHG9Wt60wG2tZw0akpBss2AbuA95uFZm1Vv9u0nqsJkqN8W
tZYqvVDlcTH3hjAFyxna/snI2GafH4ZX/DfaaMKbUOk/FKHKVtKCKzOiSS5TuegQ
7d2IGlXfVIqwCJ6UIG+2p68ozW01eoHEkWO+zSg8IKlEgdRitdgdehTcfGtYgEwT
M4QgIwFwDC5aBeI1HMsnNNqJuvTZCuICtvBcLi2nkfoNsagEQtssTuIZf9EtHfWo
9CxEDnT+LxM5gPUw0NNZYtp7dR1lfVxoUaDr+h80jE8Dq1dsaiuIuHBtgS+NwV1Q
TyFW3qsIOVwNXjjU86sZ2j0Ex7HlNm+hwSg8vKDOR27VYW7fGACjjIM6PZGszjPq
76/+ik4gTW/j4m1hQZapTyBuYOF0Jyo+hqTwUBmAlSTPFPUhJuI3Wfize60XuI8N
8kuQhQmCAXZuER0YO4ACWXp6xkxrnH4kTtAc8BsPE6ETFhVXVHAKDA6ApPV0MTUb
CVw0bj9zVPiL+AfutVT7f7jZKkCd51fkjIfZaPm2tKf7dUBDHUT27apepUeZFUCu
Z39o37IHatS2e7Kzf3UWkST/GYbExA+OV9H2Ny/mQKNfSi2pVzfAKfnwNAlxTK1+
6r1We4fhy1P4GtaYch1ajzjx0QKCKfYi8gA5ho9UXL6H2k74aToVIsEtGm0Bz1jB
vjlvcmljSYEvoRL+75m9LYaNxwX07iTzeIyqL75WJRwrhEP/aws4hKeAP9OHwkUP
plOlo94vg0VyFHMhfyzDzZojKJ8VNZr4jf0o7a5vX4Sn7yYStIXQ2WBxeOTk8/PN
QmXvVx6qL2t2uBxd40/vuffpX5r0c8j3W6bmymu7YUxeQGFW4NJgNv57s5cgjF8q
8gdkykbFTQwEXiix58wkDLgsEFv2jDjvata08sNwF13sCf7MQNTwasFYGLyV7XR2
3bVtPkx6gqmp2G9KBayFeWjMYQLd/6F7jz1oc4ZZAQGF6mYWvmk/+yRaCGhSFOW8
oOH1cUmFyu4QapqGexR1g8sPxo3jotfrKpv6vnZzxqilcRryox2+Hdir4wyWEjlm
My+jkgBf6VvPoDBp3eABqxyGRThq7Fv7Iyn4IvlMceaKNvzfn2y7aXjfzOMkGUix
XIG+0pUWnDOL1RnjRq+KQeBIFaGYrWzEbN8oFTaSRKrExbsQ8H71PBVD/IOkYEFp
6TOCQ4+74pbS97QUvqL2NSaFiCJbVAoAfP2mHyB8YLdaTvckOyUivmgNQiPTGs1Z
jnpeBvsA+noSPQFePXQ7hx6wSZtDvEXTX65PY3EZ+0gXiJ5z9uvoEfpo87mJSm3R
AjUwwPao/LngYE2LuA06/pYSwF24LsHO7NHGlJKhKzWdjzS4ez6kcpQ2rrk3YK7v
ipt7ZPKfVUaL7CwLf50PvR3Wma2yJkv27QyX/CoSJITma6TjEdUwgZTTk7+RCd1Q
v7Je1vO9wVYN6ndHkCzo4/vn5PVAj6DOrQqhN3rIs7iUHFjU4+TgN3EiHXKfsElA
A26q91iqKUZ1rNo/3TERwnk5btHPEzPT/ZohkOYsZovts31KtIECCl8BClJB3x1/
SDeDOebjJKkKjythz19QAMiVndbIzUdDr8N3r52E08B7N0ah8KHjBC7rnKCdxf28
QsD/ca9gHs3LOwNWVJxTLE/ZhvGFoYBgexr+1HvmSudH5QeIaVZbMBRCbZO3+cSk
eDCnxb3mkXJ7ZCSpLRW4wRXMhvOe+CLDrkSAmi0Zv2FZTbXVPpqCRhHQkN8YzlX7
c+hlDzVnkjpy4fdvwfkClOHmSVYGF20D7EqOeB32bSMk7uGLU7v26SsiyciZO7YA
SNl8pIF2dShZk4Ng3wy265HrTox8ZbSDygoQGGnHuDTiDEPJ9PcvKm8bMJtqnxop
dWG9D1MCeRxsfzxryUsR29qPbV9IqZw6BmoSj+BpNWreg/LPmYNmxA4rwaSpW/VO
AqasNxH1uOHC2PVIiyfkga9oe3y5s0/M1s+Fh91vZbi7nxprzcZKNE/YupTzQSuS
sA4VHcamkg+D1uA+YEPVHGuHz/d+vepW20949wHvnrCaqDi0Dcsxsfx5pD3UNFzn
RHuyLXLcmGWxqLQosQtJTC+55h7yrlso6+2wT85IfOmz+tSToN7dAg+gMDG6blCo
W4W9+HuB2R22onofesFchpAFP5BaydJKDFGLLX31gHkCjKaYRZhvAbDq02/J+E2h
btSHh1CyRnjPJzVDMbadqjHpGZJddUEn0lIO36FTzy42sAZ9BblIoXpFqJUk5LgO
z+sxYB4OkBg/qU/Pm6WvGuGKXY/I5RWM3ya5tGU1hIzQLWY+qRuYda+aD3wCerJS
rgbx+WkIuzH3dar2XqYX91kjL8t5wGBUyxeF5RRnqdocCKlCUXOWLFFdwf+zaqQW
cSK6LR7UF2wgzgfXUjTsBb19FsS9eqQIGNZcVX0r/LuzkiD9TQwP5zk4HuY6fRJR
k38YbJFcdQflDp+dfTn+FqwJ4RSfFa2W/8WuOErBfotmnEHvbT9CTepRLbbAU+Ea
ksD7vUa9SZXT4hJPtgbSddEbmKWcsu2duYJlvnwiQzyGVhjgFqV53SumJAODge/p
dI08O3/0NHw4Mbm6XBazeTbxeqzPsyF6UdKLPONy24e5gZg72/wtRV+es24JjzeW
K7xbHOjc83uHgcMHv3lz/p3yiaIK6o2O8NUnqjEiW+RFYLaJAha0+4RazwIbbHgY
A3oeW1ux+a64U8/mZfrwjmSyD1YCpV14Kw0ivMFyG5vv5iTsTQYt7mdmDUxhRFWO
S9E2XN6N4YM2QiUdMGTC/Iq9jvjyz4RDzgkAeJ+ar3eJoTwlCZuZW9NqB2dNhM7r
3TAF1Bk64WBQDyfXg9LjnopTPjpl29nuTWg+BuD71lRajtg5QT1isJfF0/NBWtOg
ZZ8+PY7x3eHyiC9uQeOc9NGgq4BOTAtiU9+ChL8tDgOnTSXH+6Ru3taZioVmahxz
BIwRuunZlAJeEar5vZ/ySlWs2p86x7zHtQaQT914MVnTooimjC/eh1KmJjIRWg7c
GjCmlosFTSRMPsZYmJltmY+5UU3INcrCpWC6pFU/LQ0qp2tYBJcYKJwtakydRqvx
3EyUFxSmSYfDZACYX2MlJAgpDWaWj+lWCLT83m8IWAFNAsuHjeZqHUSFWXuDm7It
lgslpjNlwMSnEw1/6IScZmGAtG1ebHCQixGo69CI6YEDw0TI2LxiBKc984bw4GmR
4Z6V55N+rhVNw7nHRjKVd4BqfYbclTOryHQpqVaF7ilKOMEJxY6snsY/Ip/lu2bG
Ey8IbmZIlxd92/mhcv8kpILVHa8Air5gp47rzv+1oeYMvVFIhMc3pXlhcgaQvN3x
ax+9cuZXEck8DtngEOelROr0heV/WzbV07zSlpvU9VU6F+Hr6tkloJFYSaNQ5KN+
8XklNc0SsdFxN1TnaFNnPS/qPZBkFgUhTieNZ9biO61sIKZ7M7VaxAxhp14CZ+gQ
z+D7z5zt5uGqe9WljeiGtKcZsDxWDjoV7QVI2pg7ssNWGlY+wvOkmtqz7dHPbGYv
pt6AeEerQrLXNLeIpjfzjo8Xyqhc4TbWKmD3bDqMLGE6OVfWmpGqVBbgONK+wcqv
QQGmIOpTSR030Jeb0YS5vkgLfij9Qo7zxrG9DikQvEeUuM1WUCMwMeJRm8ik5xeU
wesjJmOXaVG+7Ch1RwKLNO1nt4qFgQRZLGQghbBR8xRNu5UeZ1HqSLM8QHCBPT64
PFEbLPmY4ywQSKAu3QPusiplHrPdjT+JPQjB1YjH3id76SkApKTOYb/CA+j6t2qO
aEJ9SkCCHSTr9hSLWTJjB4Ft/Pn19CqSovNRHrMiONxofz7UvyAVJOS/S0UuMCP5
0auCFpfdHI/zaoxeEKybLlN6BvnS6onfFP7my9nZlKOMnIZwOQIWAAdWx+nsS+nu
RWKR1ohlFu9oDzzT0x39ZFJ596QkSD1OtKMeIg5AClHmuI9iUeRVY4sc3JRPSPm5
Zq6RIO950ORBgpvukg9b1xVVtVC5CmyL/DLJsVXLpnzw//5mWrt4YVzkbNuuDNlf
a2fy2jZmuWtRhBVKpqvzB3AB4OMkgJx46ZoWtJIjVX+85pplFhKZM0defWv5L5Ma
4FgZVO5HyfNPzO/AHNj9ChtL8VUvq7/tLg3beSmdUmhS4sV7m7i2sAMRUC6IIqbX
ww6zHXWOqKlp+arIaZTk2UpqHpKP4ruqC7Qgyw40TSeaTzKIDQry8fTtXsA9hZQ6
gqm6khZwAn2BJX4l2D18xPd514mKeMOc1KVofegXOrp5AciVztyRBzrZA+iMb666
e99fDXeQyJe5AqPFQ0T5ixjER4E7jqC6FnYAd65tPP5lLXHM/O300Jz/RAcMSiM2
2Lt4Mr7ibBg5VtuLKW9FPGzHBE8mpIKqdB+y1c0OOS0lOM3VGevOpZapa4QLbTgq
yFTZcHh7aeAiOIwqToQkn1lINX5AJ504f4rRtAxyrIbVPDNLA0Ccz/vdAJrz/KPl
VN/yxvOwzcFlUuL5FQRjscpTivBmeZDAo92UTpxa9Bbqrhnn8NsOtIOCbAXElG6f
h5csn3RFCDkyhYgjxJBzrEp7iUtVnpHDXGhhyXAxyCnfxnH1E2Z0zOJLSST1bKA/
h+lfQpidGNINCPg817K27JB6ue9ZnTZs0XW+CeWPondMc0579yTKxd36rONc+5gj
DAXb3DUTSwhL3+VgFAwYg98QfZDFc0KKZxyhl0AJm+LNhZI3HHMOH4RYINOcdNII
AewEAsZCqUQnCPWQ6u/TwhYKFUviUUK0CsA4T0KvpNXs2NxhHww/M5nV5h7zK20m
vraTh6cCRZ+l6YSdodxk5+B+n9rzztWw0YlHvQ2U+OHfnj8XZSH8+48cF4tHKhIy
7/0Wh3aHEF6niesandOYNnGX66yzPvqZUSs2weAHbMDF6Giqe+a6i4J+c/SGJsuR
BZ+twGUC1Ezch3dHwRr9pIvags6dVIvqQh6IroWz1v/JgqAy4gq1DRillR7yphdN
sOnA6oK8HMsYl3fN9Cqiyj08D3LJHCP5TqRKdQ+mqO/IJFc1VXkQQ4kcA83yEX0F
d0GtbQWmwgOoT6ZcjiOuPdpBVMb/q2MuebxStvgwuEyEYaISkViB/eNvR3cucMna
5Iq3ls4MN5sM4vHH83K+SCeLv85q5po60Yj6u78TUl7d/ZlTSwR7IcH2ItOoWELZ
zDOUvSOa0xlovSgjS+ZmaIrWGPaQs4PlgNGktOaneAAzK+uhiVp+XSQJeX7ElFWI
06yONOfia5eS8yKS5FYD/n3OmNhyiG+lE2FzZEOWdY+pRChph6adTCdlx/GJqkLC
2ynRYzOuLZZtp3TChCDqW45Idy/Gkn73WVUEC/75pLxMoDOgGTqxQwfuBkbP4WMh
aSJ1q/0oynv3b0qQDOCyBnmUb2xgnIqo63nb0LOIXoDgm08FshYUg8HGwAPh13Iu
VyGShsCGAz/EOSbxqVKWvxfylGIkPr2VVVLuwgTwaqN+Wranbqej42VgRdvCf8t/
9jjCPH1mg60IGBOFf13w2mC0vcEiOEZwPYRhBX72o9zE+LvtZPgUkUcPGRSoT816
jk75+/b32fwdDxDCev17aaoDHdxwugitBo0DqpVupX+DBpm42w8bhlQUXn8s4JID
Cl1K5YiksnGYp1MrOtwhRo3FJNFro6khXad+o8gfrkoPpZGpn1SrSq/w3sSTemne
rJkoI2LUsBnZof+BShcEM3978d/BKdvljm//GB8XvgWXPT5Yl3FIu6OlnD5E8B+T
yfQJNDhU/IsIZdp5iVo0+FsjSL8G6+JwHZ2mBsReJONFJEurpICey7eXwVjE035W
MVmSHAVLBQYMLgbym0aUlj1TJTGvOoV/veYSzofJ7pkainbmZP9pIlkCC/D482YH
UpvTErXIuMyr88iWuorri6CiMaO9d86LMy5M1gcEGrjWMagK6KvqeUEumKILKZmA
jvGG8zSQToigfpM6FwgPjIEy5DTb2ZcHUmFhSC6krrpnfGEWUCv5P0+YPa+j/Y9N
tLauf5qq00tXrveGb6uGq4Q7riJs1Qzo2nsezy4I1zmRovpNVCVPLNEfheo1COLf
b5ZdtPu4VVz1uN5HX6Cp0lTtoGi3sHMKUfUDwMH61LLX9b0LnsYSuOzStkDaBr5/
meiBMFLPv6GrZRewEFKHItKGc3DozIqa9atXtfVf8HyNQUipfUgCMLUucg6sHPdd
Aw64tla32PfuXEj4iiWkqaz5QiC6qgsAtHn+Jeayt9FzuK0V2V+Qkuy6jckwdGGg
ZTIUo7mkiMzPGCZLRtwA/4eVrbUDgEnFxIsFLjUhcFUqJgUaHNQMZZko7OPVxG42
tKENXPC+lr6GB/XL+KrS9Y559rBJaJiOPIgdtHU1dz9HHxqNP+lk6p0SR6DHG9Iw
ZEPOHuKdaXPWn3mZ1dh825rrTrGaEFA40MnPP7lgEpVafsTzWPOratBb8m/tliWl
AMmHoUZBPfPWxopz4rxyh3PXg8JJhN9I61z2gOMRA1RJqvSGq+TTWCTRjVumTAHc
Osgvi+1Dr182icm7z+Akr82KAQZXILE5KhuJ8hJElln51axyxa0KI+XLmFWKDmln
IoNPdPool/uNQzwZkLDqqoxZ+UfhL9L3r3Zd+RV1A1XEpKzXcLZi2VBNyK0IF09o
S4XJFoZ7pfI/oKgzyaqhckrTUYWgbl+z+o+J4JR0dAtzMrw2329HwCDYP5OHWr5O
VH4FwMy0eM6k/jR1NrBimoPODLBKpYPsrNUJBg6m9pv+iPCIYIYMyNeuav1HaGmu
5U4rAP0Nv19CJ+PWLai6Wam+M6bSt4QVfyd4EyVo8rqTy2yCdQW1tO07J32d5D70
Y7+eVsojT6XDPluflBXYPQ2RrrtscwQoEaQ2t0IBAcq9EtZ/zYnO87pHgnp4Jdhn
XF37Hf1pg4kbU1f4GZWivqLznw9aJ+DK9AIkJFMEDnSG3s25ksbn3/G3ggYwoF+X
rybAJovrySlzmI6OV8qJmuK0B8O1RxgzeUO+xuAQaxb96+Ot6xY8k/wdpy6la6Zk
MdyN0zFQh5O7hKp4fUxoWqMhV9Yh7+2qXXzOtOO+4okgMbDkCGDxPvdiVrmolfMV
NyqZJCzje9BnzcHpaePsYZnaiGh8e11+BL+Q6flZPWkZOTV7NHVQQ7+OGhn4B8+k
peLzeZ6likYKeH1oAGaWFkNt2M88nK37Ko3s5rcYACxj0WVgJSBz/lLjogZTiy2x
BwOw+qApeJhWLxn73W4tFLbj7V1vfEJYUybcsGg1/Ebpi8WBaxducCkiY2oemPN8
3p6UKG6JRthi0Efq79cZPK3cI0zKiP+40/PhMkGhl3kSQ8acBdkysBJks7v6U/+q
H1OXO1TmSGTmk7xMMcCa1t3F0oY9VCUecq7SHfe4vHY5Qa5XDmxTvhmPBWPiIxiJ
StoCSXU+leCfhxlIxVnEmqOncesRUmzRNS3GxHiDQVjqlWkipRbsGVBR0OlZGeOx
tgqBna2+S497Kq+/zpa8wBVMUiK7YLP0dAB6hP6RzVZ1nBfcG91z1ii9J2xDo9HI
ND6am2bzAcd5T6gRoqpsZpVT+E/7SBUOlIFKOPA3RLAABxIiCuk96xn4yctDkg9G
fjIat0/oTODNWgoHvZExHQ9MfHKpFnlTkw5/XqkPH4gPp0/+Z0kkGajgy1YvW8Pt
Dthei8LG7N+ErOo2CcyBjLxUT4MAuXfVG7gwOEcHMh5yYcIGTPmEEm0jmjyId0JA
+sbtK4kkzRTQheCnTyJRnfLmUt7mPSMg4X8FG5WF+dXw4afLuoauTAZ4WxDpXaja
Oi864Xa3UJlh1xP5wvwnj4YFYLM2h/DdC3UyWVnu9RueG8Bro+C+1F/SlVZ8Dled
tvVGbhy+4i/k95CNokhpcEcjdSk0mnY8t0pJmz+so8C+YRX0Xkb/xlk+qfRrJ23D
pfm6vReb+OxuSHcp8aX3xpR1vfDxOjQYO1Pd4L2M7VyOeac6I3NqcbCVWx2ceGPM
T0hTyTcPbOAJaOSSZ6tK3KCTgGUt+ybIcAmPgvayKO7wUVYNLQ34vnlxvn3T/Eh0
Dcr8ryT8o1hAjQxkdK3UAP6jUSNESFvWpiegjP7eS6xDll5j+i9rtSdCrWuEV9dq
mgO9pYHAO5GOQOyU4xBFEK99p+i42vYgzEscr8UcR2Z+zIzCDFrpRr35dpjt5BRo
st1SVW2VCyUJWUxLO37XLaDis9E1pVK5nKsrcP//Au7bA6yLhmW0E/q70GbF+Hob
eEx1doDFdLeNpmtapGlM8/L6dc6y6IijWqti0xzDzNVL9+1bMDtoaJ7xfWgRlrdH
BeNnHsqJi9fMu7VQRGNZEyxqgB8HITOWVQfuJlUpAdxeq5J+pbyFIf5fgHo3+Htb
a7CutNfLGGTp5Jhf2TgRQeZNT5iVzd3SH6vYEst8mLBfh8YXO4TjxT3PrrqgRzlG
AqbcphN3wtfXZvn8etxyExNMDrYMB/tVIfnVmJeo92JwHcw7bdMaTJIBz3g4zxaE
m5YMP775nNS2TA18lhP4jL3ZRSppZL7k2PKolLgQwzegW+a6vnSVKL4vmcYOSfY/
Wgpo6MeZMfiI8TfxFbc9L+lhLxdZyht2se8pSkrLE6ysg5ZnD8M5iqSHGdwW4yJ6
1mrxTJ/AOSsMWK8d4x1NSB0EYgGeLse5qCiJFITmJhanLEI1fXPKegd53G/mgEFD
qT96AWLEVl6zaC+7JahdO5qf5605j7GufFX5NciyR/gwScCmKj4wXYhoNBlReLIj
nKiNYPLYWbf9X9DlqKXSIAX/82fqSxolOT2HfDQBRHbshtys7mBJFuhlwvXPrbeq
CfAwW52bvy52O5+4LX691PVsx71Wk7pFLMLkt1AlaM6wMjHF3XCUYDrAzrQL6iDQ
yVWYY3AKRscMe68yhRt2WwtJy9vIcJ7pojIG3UQNm6kfXh7YAp2zExvcPvyRtHSO
BATpkISIXS1PlylzXCdB3tvlPzABHyTu2qW1NOaLbD1HP/OZMOcFXlYgsliw05+X
mUAZ9gOHp7muvOsS3jcUKnuoWloZp37UrG4YzGZ5IEte0at4XoCGJtOQobXEyUUy
vqABGI6GBoX7/0MbuewWZpOTu7+Zif4OzrhzfJUNPkcwsl2/iXpER2JvE/tRmHCX
w3tJ4obDLcbiGmmZB8e9bcRi2CDcb4+dwtrwD9hUbM7Z3vIoyYFio+s/JIC6faxx
iF4DyhylVUMBDqLW0ikf0wQGQ9k41/o6Nq0nmfv5Y5EXvZc37c6JOF/O20WXm06l
OKiQ8H3bfpQMApu4ujrbn7zEFED1fTjgp2olg3/kJDqEr3cHA9FyzLfJEwYHY6sS
2RuXeqvPwCUUjF4le4T3lgFoC2IEY+39SnZw3tZeTJDl3SUkMWl8LR7cw9wQpY6A
gKEYjHITIUgVkXAzafO6ACoQwhOidd/m34yiJ+1LaoMUa7m+vy6KkSlU3fV+9+zG
y+MsBh8G55BtDDDVHeuIGfajNWFSG5MAuRt4Vp+tsoM2se6rzdeMqyuNwfhYaFRa
ESwnl6qJATTQYzbfb4ZoKYDJyoWa5P0kUW7RsdegfojQG23vc1659nCLaIAGdSHt
zJgwkboJNRbaqhm7ob5mvew3iGGTLiEi/UGxaaqhgJ13PO/61zQCt4wnkHzfYX8n
2Uare5S41bEUlcMt0rern9XUiHCvNP4wiWEJ1p/AYCRhKAxcOMRWxZ74/+eru+iJ
iYZcA9B7ul93acC3u1umM/u36n1trbn5Faa3ENEYIk3WGoVCOuVQr7K+aLu9OPQo
AIz3+XSjjWoOa1UEpqizxBrY2KBF5vyAeq02SKOpomXVDNLcBJKkd938gMQ7I03n
fj7qzMkvaMfU7h+Dnl287WnCu7Z8h6c2fbjG2+Hm+YejQVIpkqX6Pep8fN8fV/9g
kqeRVDNQx8F/4X7srAVvpqzopsAi2+eyPSEbe69usFY6I/HwzkzaDHvMIf02KwB+
kbwCPyk8n5IBlFA1e64BERr5yWknUP2GYgqf8NaahRj5S8zIcV+SLfzlagn0j+DU
+H9Dan+xrdBnIxWFeb5PtDbHHItQDMrL/y7MTB3NQz3NP5uV5GBOcoTJ4GDA6bk+
VwpxfczDhzf+0haqTddCnivmSTxQu5LsXwhDRenHy+7Pa0k45RQnX9IRwcWM6jae
ZzGDks3BmkaekaXQTsOyLHiAqzkO2HbWlnf+CSXA7DvZj0mMmgG4uA3kZCZeqTDz
bT1ySfsVWdRv0K7CzjcI5i3uRBVCEb26GgkbAklK7W6DxCwRaeB6+Ec0dXOsx6d0
xfsnNbixPt0dFnnNJ3HtauJYjPP2q9TPPUw5O0fjEzacVjM23a7XL4brFK+TSpTP
u3V505KWloq5KeueYzu2EgFcopl4E9Z7sbK3RGUz/CmoO93B1r9QgTgXyCMR2jGU
p0U99eD1e8wQNQ8iZSAYPdyNENR3ZwRgJoNtRjuloKByRnvZv+NWhm4dozvxJcX6
9J0APFo7+YNnjMzjinL9zzCpqEyuPvhzbZL6kqOA7weKjAlDTZYBTYPLUweRe1Jm
1etZihihadFTC5K/Qxi91zOtac3gMC9W9+5OXpJ7eKRpi/9TArfaa53vKZTNGMtq
T3h+XoQffeyt6t5fss7UJvLrN3o/Z2ZEk0fq1DNRcnagH7XsGrlVgZo3pb59rTnU
pp3aMp6tA+XmoJ81N6fbsLKsF+OBIW+Dcnp0MsPOudUKdUwGk/jTcgVdex8pA2yl
VecAeRffPgVEJG/vCj6yTTab71QU9y/sLK98kV24da2nmICFQmEpsKnSoO5IwCLD
5IiG1BaZSVJoLhv1CHoaBuQUe8FV7WVblhpCXWJ1WhtxF/9gNi2ZFKPFeoqAKdj5
siE+cHU+4bk8vbHBgtEbU05kUra7Yz07Qh5YjNQHjx9KYAhK4eM7Swb0kHUBGinD
ee8lj/z/pTdLueWO1mR8Xt6+bj2O3rdke3iApolrbeMQsr2pGBb9Bnf0SPxPQYKM
KUtQT5Gsc1fDWteEsXeUK/7+Nyq7yPLDo+Yf4wKTta6vNpCLUD8vwwIH2E/k/USF
47F1yptB8N3Y2PSbXL6pO0k3iwX1Nn3oDl1k3vaBuYzSQ6bpkvFlkkCRCU/NjXDZ
uMsRAwUwjmm3OCLeP09TtO3h3vqBM66muPsPxrfHbt8+UUyt797vrkraGKuwT61X
TQzaatcLa/DhO748H6sc9Rx6bOVEsn+OWAWyIITB3rNnqqWSGmQAD3uyoYpLAW+M
PNbzR9q7/Nu08SaU7xQUVtNiPeO1wQIIAgkeMS9gno1pB/Q27LIXONdaO9LPYXou
36McpsRUAGhPcRRgi2dd84TXEtsixhT8ixPW9IzeeB4eBOD1WNDUcjuHeOK87Vfs
GZHtuWvwuFxAjmtV0TWxP1iId95Q5yaaWrNkXeRqkRgijWcLT9Fp7Y9V3ieGyC+7
qcW0ytRlphadbckQos3til6iyrEUxuQOJ+n/R1X42YO2UhWtu6N607KvCG1+65cy
3ID5qPES1NPxOyEfmVXjiaRrcFsPuRwlYJBmZm0hlcXVpUhtUcGfqXHgnk7cUGer
Z5rpajgw+s0sPSfAK4Ak8LBaEByL6vMB7ZLNmmJ1Br3ndKE41q0hp3ch27Uo4gbq
NMf0S1NZQJXKAUvQXCpylA/dlgeCCtzZL9sVio6rpgEZDkarZOQMvsXFSFknO6fP
CufSKoe6O1NVW87IryIV88JEhKE219HOCaH7/2a+uV8Qr8nbjpFZFU/B2wYLsenV
CdhDFAgjc2nu1ObsDacnpw/B7nXyhX7rb6H05qV4IWQOpRjIdx5Sq8XyQeFimgBS
HJBNgfDeHzMrRNytfM0CJM7QydoPXrgKUfJcAYi38XnjbKWEhObRP2tFWnhUIs2p
hHRj9zr+jzNynHdmpHwZuASPpKZ/36ormAUZrfWd8NwjOnv0mO0w+yjMwnQyIHBe
Ng3q/I8M4JOxgHBUxycEn8UJ2grSKwfPL4UbHzAxTqMauLoDHUTogjcx8oA9+UbC
ORby7LdviKcYpJcPFjGr4eYQfaNtq8Ll9eBmumIVy3DNI9zQEjZn6wsv/rM+JjL4
x6GBGH0+rSCeWQnBki8mYfQtc+Le88fHBdjXnwbdXuCULurxKIql17x2wFH24C4M
N9WAWt6OVLK+a/ubvYcDRkzwfhVugPqDKzYMX1h0hkTc0C5PG78zzdCz4O4S6cXj
k1dgnIV4cI2rKO1PScOkc5Hpy55MPVKXSiLx4Ufd2uvNvrBJOSp40Pm73rGCM++j
7szWwal0qkLNB4LlMKynQAbikGu6xpW4f69BuMkBtOOJqRffBHPg15w/+xhHIJ4d
S81mKhzCRUcHWxDWgrcTdPbgZBp4ym7w34z8qS45cztCEFV7ScrnOH/I4C8UkEct
9P2T7BzmJNFh3mJVOZSIF92kdmLvar80h0IWTUdPvSXj6btTf+jvAQvK1xMhJbgj
NRi9w2fPd9CJ3metJMJ6J0o41B7vQR+uvk2N6bJW3w+rA5m5hNe9dqTw3rWOyxnm
YyagDW3pRxzJa1tg7EYWwQtMzuVQkAN84KF4KnXVJDU51XXH2WLALlUoKhs8MGM5
8MtYqU2oiSt0If+/X1LTHmS3Y5p0odF394c4fuM1XdD8yMFd7n1PvdQ0+pabulLS
YwKu9R4aaxz5l9UpURuvulH1Cla/DpP1D0rnNley/eiUaev6CYNTKkmOOKO5xw1n
HsMf9Fkdn1BKdIJiRPtT7JdcrEAhu99CUS8JdaLZHN40XmDyMNo5SiYz1xHviN0D
ZQeP7qH4A1acPmtVAyMEPUMwJkdyStKdHLZlQ20xSfGW3WulSKAgmdYjSaBB9dcD
+S4tO1l0Id4NvmrUKBEQLLuXsuBN+LyjykDVIE6BeLO3RMkfqwpMTlBH9IP4pnd7
A/oFc1Bb2Fer45h8y/hPY+iYqHIc6sZFnxdqfiQtovUYiE9HonwAs+EwRj3NTbPD
XCUpF4hnNVG8iicmqn4YG+jvyAvzoSgpvpvzm8StGRqtLl1jsYU2lXRUhDFIk1/X
3aUUltsJWm4I/DHW6Ag5gSEhO67A6ZGBy5v5BqwzXlmxaZWOFtKmFoGwqJ5ISbu1
4p+GOMB/5wi7L/xsWQCryRfQyRhQ5iUhsA/Oz1LOrmTl+Z2dhuBVm+fz6r6vSXS4
tN2wbSVim8T5gIGKKOsV8Rzr9gO/D/hEEETq4NLWZxogva8ZWZXQZXFDbdlXc9Af
u6VMzVXcGvIjcuwxe06aU3eVuo5CSJLePm+SHue4eW+a4p6oIpqSJO3v4W+rUJwh
e2XY4dhBiI7FWpc8JfXkuFPqMEGMTFHwoNv+/O1Tq9HT80J8xZnvptKbztdmUOb5
fevIQXngHFrCsFOyFT9eUw/TbXxf65Km2QpJl45FlD0MwXZEf1UchefsbRNDrGhS
dEZ7dV/vHmOzpDjABLckXR12iUwFZ0HP9LpV5MgnhEFFhlvboaMPiW3gSqAKk2cd
jRDhBzYNWAJb11neITC5ohpVmrZLQvg3hrjximDELkxvnTMZw6dS/KRLfy2X094z
LJxRbJJkJy0FcuHp89tvjv/RIs/a8lg9PoUVsHq/zpb1bLzvdjZrGtFZZb/+n5FK
iIE/kObeEtMjO3mMbSsSDbw3MJHO48iClzZW6egzC53LyzAmIOdl6vDk5pQ3aqoL
anc4lDVl7nUoLlbw0SclXKCEJo996pENm9kbg64VXUjXI3q3JwqAK2Q4MCr69x4V
7YpvWFe4Hj9XsBKHP0+gN+eg13B9/oJg1WnbJtuCsEkxJ9trYqtbK8+b5xXchXBP
kwmEQGQkjw2pttjvaVEsKxDKjfhDCZ+oD7ZZKGVKAfdNQNTelvEnVo1F802xrJJB
YGX/hKIlOiVJkfVnFInY7AKiDQ75yq9kb5pgRYHqFfUZsSZ6tXj60beFHT4VEu1e
qRLEJFR/YcocNfgDNax0SMnvFTJDCk5J8BUqzmaoBFg0kzy7Rb8s5Y3ahidB7kAl
7gWBhzrvdsc5NeeiyHEEJpGVJfzHM2fnzm5o7htd7VtUt8q35Cg8TZkrjtyzh5DD
iW04FGSKbWqw3wVcGTAaJ4AS9krWfAE69/ts81SAT6pJdFD/wn+Q75WUtDAgsD0X
Bx9Z3CEgdJMy4mVZLyPV5bbHgXJP81IMM0a/dl08nzK8+ixfhHaSQCbqxarTRbT8
D6Rnf/zcFfLlOvi9nSmsFT2WfsJNi80M80BD30KK2IBsGQjb2XohOKP10Qm67l6r
D3lVK8mE6cqRquRPp+xozK/r97Y5zNpq0lVYANGWisq1GQxMcRzabZKfGtvCJ3u8
404rz328SoE3K4EvND+dmrX7FwfhSo7vM3ZCEaEfwyNzM5ocUkgwQMCsLbLlxbLm
6pI1skS0kINlBjpkt5ocEZGi09AxZ8k2jt4k2bp1aUD8rpYrp+KJ2k8xyNbKLUGc
L0q0jRyi83k/bpxKWTT1h0RDlEXK6fmTvrGDfiZ14nSrkQpxc16ssC0nILipauFO
K+81gBm3XprCdJ2nhVbQHmBUFa6Md/usRosVBufYqDHe5HZP9e2KUmC0pncoOntX
ZjABi8PM902xBqlAprvOdKwqsXnpn0xHHzMfZhPP0DahtrEDPrbqda+Fz+O5IeSK
xvdO0fC56rN7ic3RJyANQ2mEtaxMgLjmfNleY0yWApPGNDYzvP/wzfXjsXRbDeyh
Maxp022DJw8qwHne+fzhriV7YGFRayuuW0f3HTlLHbW/gfsIoYJ3sImHX2kwpJJb
IangX12S9EasgfkZuCTxosDlPUAgKzKiclwRwEjWXhlGUyEitYIfGUTD4FXbTa4o
Chj8OX50JIBzNBDKz8TJ7VZF+/AZfyy74uS1r1Xqtja/5ecRDlCC/cBnXNhZXirD
kJ4n7le5lNakNf0nUqf5jbBgAHE0CblcEopCU1AThhut8i5m8FrCxlpuO8UCeGYM
xHgIeGEIUfr3cruG/mOvx29aiDsuwo1qQwHf5156MFX+ZzO0C3JDtKflr+nudbNw
BW3aWv1aMptYe63DR0KWxDBVlmFSm+iz1CKoMpkbC1Hljbfm8Pj0fLTgZROm9r2u
pCHnmKOZ4RI0deFOu04PngggRQ536w9eZiDXHngDCZtNqz7/4wNQvKXn7yBWgD4a
w2aZC1wEooh+LpXLaeqmu0WFpVY3T61J2d5xJ3opeiNItvzzvaoW9YGFw/gQNB1N
8xCinHAD5dJSYbuBtrribs0+uUUFsCQJpZuJ3ZYFs0JHqI5EKY1ralEpjTe8toQX
anAagy7dmUNhFlTtMAJagaEoc/GLtF18G3k8UWoYK8RjAWvDqtXGdu84XRv1175y
5xJ5C+vFz2zYg9qj+lZ7Q8KwiiegwkC0iS+E12DsjP9S/b7iGIEpPaVZV0wvjhsG
+iLT6B5VMs9oV7kFYSCZW3oCHT3wIYmoVvZwhc14AklKr7RBeWVZiQrDy1G4nNJf
QUelnNOrjI2Tvb2PNv1MICUqI4HbsRta9CSifRnZ+zWyOyk59IgM2QUI17ILzUh7
PhQ/VA/sd9iY0cd72iQaKjymiaf2JXwfoHQJTlTjAsJlOcolPfYL5RyO2Jz36sA8
RRfv+WrMGSrx1jmdb4dMEtVRGWHZX2UXoCXJ+eGSNOYNkhiliyww5mFlicgGQGqS
M5mvCRggGYdzMhLRj1JrG91zRwPdttinPUA0PsDelIrlBm7j7vNbMMVnHxyUBu56
JDASQrrVs09PiK/H3uXQ4ZLq3KNWs+iq0BYr5+Ug7OVzbPGJuyjBZZJXpWtoqZuY
XW0aKS6Lff4EYV0niUuZOmc2wASfNP7r0tXkdCqWb7n13FfYScNyRBUC3WDOVogc
G26F1HD7t3TtK7UnTEKUO55M1o8FGKuiJidfwKtUMmvroswe9spZc500o42E2dr6
uddVYyRdg+zYQzJIcbwKWWx1E0jQHgOIuCpow0w7qdCyAxlJuTBhuKZotDKkxVsv
D2VyGA2JLrrOCUDEjLCYMvPKDNMud+MS26hOwPfCR2+ObMYmKr1Aek6eGpCMJznY
fyz5SRR/YDFIYnY+OSt3u2nyUQJJ+vA/hpzSJDoHvToR6H2PzRROzEDZ0tC6RbDv
OSwoX4agJ34nIeTPBLkzzF+SGCq9WC/xPDyw5043rI1pFUJqkl/NQQ5Ur2kMD0yg
5bxno5IDzQgsAmblSeJpIIycTY8qMZ6XMeU21/hZxy+heTgB0lm70rA7FBV1xN0+
PxX5pYqN+hizsUcF24u6bIMsRfipt2iGIiEMmupLcujcCwsalUkIbqgn7NJeJGdg
804ZzEOemV4iYp1bv/axx7akzMLzMTL0umKF01ZouUU53UEFFeYOU/3XwWitV+wv
hwKAmUUNFfY1mOaumeBdeHpY7El4oEFxZWFGcy9xvDpBXUnSalBOX+ZMIuLVPnfy
eR73CrNVyhhLFvnem+I81m9xa7EsC6m8V5Mc4ylfLhQgstBxx9iFvO9gz3TpEs/k
/pcywF/bBkaejGBhu4yAkzG1WOkPNB1ueEY6LVLSS9hW8Bw6FtmHp2cy0eQqt7sf
E+Bap/IVXdDbj+B5iAkU5+QkeYNmINhVo3GYeLLh9xbZioqUeYYwZt+T0nys3eXW
VjrBd7S//OYukYoCvQvT7OQTZB1U/lDKeLOi/QogOeqRME1mPKoNq/WUlsT6g1NF
QG+0VGuzsHNVMWB52r0GyPjdPW6JkiVc/yFG/FzWNVGii0IuT/fBaSrlp0VKsJgY
LFRqRxxrMDrHYGfwTxImoZqkorcIyEYrMD8E5DC39obEwkt/EU3E1RFY9rtXjPn3
pB5HgVueP1AjQey+OtgoBpgG4tImVl3yGtWzyDzpCnKN3dQHr+eChqMUBYrhaVCS
YFPtMKKIbwD4bkFd86BIexxYlWYCbEDipF26F9qI4Yg9O2LF+bOp0frWfEQ3VTgA
y8u4hlC01ZwGfN+0X11w35bDgrrBcrLKo4kd54yZ4g8ycuK4tQ12aMn7M5DD0cIq
VcoCfA2V5o/fi1tBKexa2X+zNJQtBG5eo6mWck+j2gD2Np43q3p53JkNqdwz0XqM
a7kMJKh8X4rP68mLSgOhPr5sNHMdfHR82cKFunkRhiTwYI44LL6GILr90x/Gjgxl
nNHlOhfuKY3C/YJyOof3TLZV6PtIeR2OY41J+7SUUr1SuMMxa6lalKTRnO8kEFX1
vt2uU0fnfNTDUjmesF5Fmes2JO3ro33BPJcfm5FlLYDYAm0XWblafwFBXJx42tTZ
RTI4YCLM75U1vv7fyaA8C6xeq50JsKJEnBT9lnDQCpvJMtDlHp3rlDEu813RwLk8
08Lfm3h0VLZ/ea5NAqFKslMI7/nw2GWYgZ285YKt8qPlmOJS+xa3ErE44AnwSvzC
kSSByiD2YObFUYxZGvPJKfT/pXlHdGxy1L/8Y8byqEsvxlXRzFB2kLlNmwx51J0k
yMyFHV0x1w2Asw18K5JlOTQW5vTx3H0pv8u/QizvyY5MmEwAk4hspdIEuc613rle
cBDqbUSyvA8Ue8FEdA3h4awosDwSLFeiEaDuSw2H6t81vYWyjilwi+ZMJ3gNW9a1
Xf2GZK/5Ys8COlUwi9CNRnUuFQrOZe1MhDwJnohUL8XLSyFYoBsbeeMK+xFUhb2N
pxNuQ3IN4AhDWp8jj3S2M9/HcawSc8bfL+5CMcB7rdZnVMw03wj1y7f5LsuXq4v7
whVwN2BTUZjc1uQw9TgqiOU3TxNQnncUp1DDoHd3PEi0zOXUDG4wnjClUhcU3Tbp
RfgBJzE0FSs2VF/J7LavJryfWgOzyaZgMAvRsxuEgYTZBR2VNYqgvqqEcn6jLoK8
pvLxY32CrxlXmYy80zdrJci/1CIEOTVPSOQ0QWd3Rg9Q5ugaZyqh0FYUbOLsEVHE
eH/WTfaP5C+zS1vWB/eDDIv8Fis0e19BhYK2CTPRHAhSxopxb5F9PY3rc3h6Vpcw
NBHYoZaxwXZURgqVYKXE/TjH1HEyDabMS3lmyo4g17WaVuVycQxLbERJdEx9OUKi
kEk0O7Ei2AXgU7EWmcelK8YFUBs02WarN8Dp2FsTp4fNKxsjgaChVeStfzDv8hsu
cx77e/dmLLEygrB4x4p7LeJnPlQgoHgbtCdBewVP14gnr4+mIiuk1Y5ezXwbzxgS
ZLpsZdjeqoRP0QYG6T7P67S/s4v40hk9l5MKY5PPCU23xSbXLsQZCIXSM/IZLCgK
o9naZnmYtsJ+IYGq04ZrG+jO2Vtiks6eQ59zLmXz9IZzivk395hXkUlFteIVz0KY
Rdmq6V7OLdvZr+5+NFENVDp3mJjZQHkXJqGP8G/f04c76dZNtf74rOhKQZRgFqRR
1oDpfmNxtkyjaXFCRuN6P+X7Ba+vm18oQKJj78G2zdnpskPfDYZmT52lu9/lew0R
vUAVWlA0AhNKF6Mw2C5dsPC1nhP8oaAIR3knEELHdaR77R8WCLEzu7LV94uyQWEh
oOHlOVrC+71RSOdhuim5aRwpbV5SQ45LbDkYUZLoT/+AqZuKiIy3RGNkdTYUtoYM
V+qskqEsqnQCIIeubuFn3O19arexVrOKMLy6NowHNJyi3gllEuhy+Dz5/CsBIIRZ
YplYXz+S3e19i5PhCH+liy94Mr0uq62rnbj+2eToWe1F46VjqY2apVvAiGj0usKt
+O/CIRm2TXw4SjInCuk12jc0zZhVEEbgK+0lBRVMgeh77x7oxaky9UQwDYxG/oz5
prX+FzEI0yHA3mvu6tAMCRuw3G6CjVwBTP99P+No4aAiJ/2eMvtBwsNyZAdswxqq
xvN5YnbctKeR/drqWgAvi3DRBFvHhez5ajcG6dezb8r2H1QMIRpqhCl8Uf3iJbXk
kOjA9izp+Jjn9vh9dvY0zdI9cayMfuTkJvBa2MAoVWIDkcoUO1A3kCCMQ0QX5hTC
IiQIEsmxi7WDUWRLWbLwfGigt8WzLDOEexDJ8/LdHCn4FupCe9irs7K3QMA206ww
m8aR0RbWmgK/C0CwnnH8dxFxbEBET9x3/RGTg7rChNQzJMXaOrQd0r2zDld2C7tK
cWYnOgpSivOF57kDh3VzR+HkSAt9wHrWEojYAl697E0Sr6MJsqGyYyCV4FoVH/sB
3/hM0LZSNi/x+EVEeE4/rKuOtdHSpw/WfJjfZcNl+m/ZsARs4oPAs2OE1kwRCYcz
DQOfji6fPDZF4Fu6HgBKU8EVcqQidUSAqeyqY9LMLbH9mO2d1Hfo6RpEapaPKo3n
ESZoXwZ0F1mY9mLV54siFUCqRmMWJ1JMvRTPPQPbTzn4W3V/09SAzaG6FbF+vOTc
Z7aU3Iw/7OHD7zXZ245lI4AZa3Qsx84lm9cvrRDGfYdnbXyfsTt8IlegWGcfLOiL
OmGQORvCtIuKIJDFN9ILJAnc7yA4y+TGssgV6dsYR5gMUhpbSTCjGITbHfOn55iG
QB8gwyZ5vYixTehEXbMPWBe+cz4IrP/ASnVgWHE1yHzth/U+OZ2JMMRgV5Ifz2X2
NJWtSWcm8GjKlQ12sEWOfZdLLpzPr7Q2r3XQ7trtB2+d/hbedByu0DtWTl9KGm2X
Qy1W9QTc8c+l143BuerxP3m0d8UACB/ltGstb0tjSAdETv+54wrM7yeTDGf9FLyo
bOisugu2NvIDaS4v1vpKVQrh70pKXGWJ+0AQtBsaEkHwSUKC+pKhdyE2pc3vEIxq
C/iVafcKt7atOUy8823PWatKHOqNJ0aoq/TRP9DXpLRfLSt3KFTjeDqt5+7OEVsH
eD2n0IUSoUm0CEARrU4T5de2hP7BzaaoDzxnZCfygayG5oKdrQFCAMBdmu+dCGk4
qpiEb5jLfmpAcZ4uZJCeEp1kiak1kQ4Qg0b3jSVoRnd+RX5S210Ob46O0Fu1KcdB
7uU/YkxsxY6DUjcYpmyVVHYoS4Rms8h5Jklm9I+AoD5DXU6nse93xBdmQ0+wMdb5
6igqRREj7E5f0Qw3lk0FnGd8+XisdiFZ+EiBGZc9aqYRGZLLCRA/NAJfC9+PA0ij
/Qf3pAM3viXW6rbu1dDiJij+Hc+9HfPz3ytd8att4qmmwGPlloEbSV4JxKMCjd1o
6+t7b7vXoybZuLEAmHhGGLqbDIDbuDTRxSZLdc0Kn4Xqj/ExcXJHOB/M/8CmOdBx
jImkoGWw5T3TywFKF8MWAh/rxcxS2hlpfyxWGEW81WrrcpiwHpGZfQIW515mbwmW
OyzdTAIXNAKicFfmiPlHZfsoRcmPLmXDdRSUtXDhrOjlvJLOPMgh9mEmIYFpYhol
mxa0XUe3f/cwtLqID4y76DWXN/uVkEAp45XHzeKyCVo25kNE6P5SByiy806d2xoa
RZS+BnqRM55hLEsICTa1IkbIP5IuPT+A8myT/1V484TDoCrmMnRhBIp3g/g+jvLI
fvtWHgiS4As824UP5flr3xTStv0pyOFjB9cOlmKVSC8Ku9/PJTk2jvXVbEdjNG68
o2rwVMo5o+FCDvLOWcZr/gAbG7uiG3m6PCfWS1p1Nqj62IIRpapWjlK0CC/Vawlm
p3zREW9X12YlBIV+fTsQQEggU7BWUCZA7C9vYZOK+2Ij09UB1YpP3zLTaWKl5dT/
3ASmm9caCQ6KLfGINwzalz1WFCmJxm4i10Izc4V2cH+pekg97yYKbWEJdRwQ6UQ3
h8mmdyT1Onq0jMoSOj2hSUxfKz4S59UiJflClDSPwHGQRkcQdGf14AacMKZ0Fs4K
kRpe1+t8PGmY5C6COXv+ySagzlpNV9jJRanKFyhypPMBr3N/RrciK4juFsMYQ/HM
Z+BAEWJq55oeX2cj30rqBoJlYmXu5ygH+xqVNsMb0QtJrn/CsZWEyrJPxIlWp8x9
lrN+rZS6n+1Ue4/Yf85ZPoGGy04Bw3TUgevEEFEbUrKrhIlg6DU32Iu+V6uNqTKN
OhxjOmBw5WS/RX9s6NxxIkIq4qR9GG0ENEk/oiPtx99pjs04XDqcG5VTPPBVrquq
dr7NUzlXFPjBbHLteen2KK1Z/wdnXQI+N+b3pKEJLHZ9o0My25vcKqf4l78+Jv9A
gETfgOFuy/mPNnqox8+DsiYpi/Zkc780wbMKaSZ5QHnJ5tWScQLkRHCGPnAty+6t
hYTUjs9g94nXJR/Z3QO0CBjmn9+n2i0TfSfv/0YcgD/OmMZSM1n0zfj7mROzfqFh
tWkSt9DTGz7eHPuxH6voGW8DFxMHrDdMmfOsvBf2lxmxUwSwSvPNS1VPBnPs7vJf
mzy96IMyApWiJMw0Fy3p+EpGMhI3ogW6cpuDRjqtrb3iuclYtweGROrBP6rnWZKu
2sNgyd3VxLEYuGwQBbFSCXA0O1xMllY26U0fpoM2pXiHF16StmYRIh69xLjJZqAy
0xMbic/dk0kL8metR8OIWUzMyr5afTYx3csaBPDQ/hneTrfzNhCzVZ/Q+YTPPxgi
JMWmvBqCy6Tscvv0mlTh4Liv0EHuTov5A48MG0Y97GufYleHKRbaLw+va/M6xTx2
AlY8/o/U79dDObogkQ1nV0vOKusSRCu7pdoMACXLBhRVp5t6Z5M/CNmo7ItvdFUh
Is51s12lepTdUZZmOXP0qVxG9X39eg0cRuYTmxMSN5kd7G8lVas3eZeI+uIDKzWj
N4AoN/IF1Ns5wzLKjeSDZEUL9EUsypeAD0UsIx3mnYoOHvF2VqAOpAJc3Jz7/Wo2
PUk9fXXkVyByLW1DIxTPeEcgF80GAoYDo1fHRA0CercBLE3qrCti6uB1qf0A4/n2
XzJJi6egj2z+f4Ut7zZmYVpmBz+ti3eTqAWjvVJgV+QBnP4GFun6iRdeHfq3lT+P
23Vsu33whYuRo3FXlUAMvpYHbEG3mhQ4E7k1cbteBeSLFVAkNiLFOauv6bHHpMdh
LzeLpAoncP8ChmBnkk9AuwvvNuUJDI9Ho9PuF82+ByIJ8KpUyjXFpy2TNv/Lybu/
9SOTLYMEh63T+BBUTl6YFWkUaDGZ4kevsdi6hUU7gL4Ab895wsekwioQL/FT0IEI
e711WmUD3ZwyDnZvgRiqviBBasIUUKVKtjYm5DT4zD1zDBkKu0qdUfJohSBDIVVd
uGmWDKPepGXHkQNlmedhvG0HJR9yxC3L5tHuQ9pJpnbo8xelOgHSMtaqjsbgHiUP
oU+Oq2IR29zUhsxjc7fhuhbAlgP8y3y9qv2GcxvEV4xLFyj9yl+ZoXaX4cdAy9SK
otgoj0JJeF7+fAh912PmMOBw//0aSAstSagmCYYaD7Jo6IEaSXneWPqPbXnjGFgw
3m/D+ZGI3iBidFQdXHYJEdbnXySqsozWOKRaFkllzaq+ADbhFoQBhVVl0ZlaABa8
ozeLXNA4M8V//G9q0nzA2VQVC1qtrdzyNzrYq+HJsrThh5zV0HfHhi988Uz6LZ2B
jEqtbgJT9JiJQ3bqC3Hm6P+PKl2sbRuFqgvY1I394AQvDJce0gMUC8TLu1dx/fAx
hqDSMO+uFqD6X21X8jl8CNkET/gNcoRGiWcABfeWQQokKpwgEbLVUow7JuX0+ESO
stLn5QHWBC+rsdgmJusCi0o+fVkJFw2h+kL6ZkF1rYOBB5lRTsJeVmKdF3AqV00Y
5+ZMLzvG/TyOyMZw88EtkD6kCWPCj5GxEx5Q0eOlu0Q4OZ5N5KdSqPKnUG3X6viW
jBkRJuGHmCjkofKQ2xyUdZX6dgo4QhjaT1py75vA+DZc6kBxh3Cbej+PF0xO5uJH
iCN3XtAOwM8T3fhnTe6S8NiR22unrazRtmZJogNMk4wLn9E1ji0ryAeZZ72+n9Mi
sVNwBFrGoRMF5+QQ94QzzSqC5o/KImEVQMtpd6ZcszxH80Zmo6VUxgA44gF+6+zA
VkIjdi4PvBbW0YxyaYWzGj0rn6WJlQDRovL6JFH/Q9SDQgJX63JKRXJ480tUlfVp
LHAG2006bRpkfZzJJfPWZPuuDCCqsLTiNn4lqvOpd58Q37Se5J1rPH80DkQmZoX/
eWz+cGlqRMrjxZ+gEYfeA0KjDk0H/WW0yBPZS0MtzKOtZD5zNQwHoeEsP2qUR5W8
JUD8tLAaGWr3bX2L5/eMcpaAkuj45gD4y9c+tnNIyQjH/RyqdjT2Nb/9bdAl1jfi
vWSbO7Zxqq7XxAKPVIFV9xRyG08la+vFNznuEQtq3AyD19FR9Tc71wkYAsqYK2Uc
h+hnsodO0rq4pvWJU90qrAafdPq3FqfMzP5nCJc8+LjQ15mXXw2lt36no4KY/55i
FfQI69LWipoRWniUq3JYlyKDUcwBujp0JUaC13l5vrzCyBILYs81q8goHgxVnlGG
II4jXQLyFEzZY/I4BGG7risf19JsA2i+LKlp+5J7BbwAe5ec06nAIaLz/F+PH5uL
haHerOUh7dejukgQ504rUF1rekkG0UlZaXrpm6te7eEgcABUElPb7c9lR2IYMkO+
1Lf8S9uhDKrRa/K78uVbT//7+BErxtuKvkK9H1DnKSJIO/LTLUhYdiAPM1IfYj4v
Gddhob2hm3pmQGIwlNut5GYilCvJkshALcNB85cn7p56bytB9Ojz/XGD0PCFloVR
kZR2LMwhujPNvqBaPsDxxX0O4JenHgHYn6egj1HZJbYv/RGJmlv2dOXuSTd/IIUh
0qbj66n8wHsnM04DzgqNxFA1QsS8R/+8Ct8qKZF1TH/G8k9NCFH54U9QISLOazRv
r6wpkN5XZKRCg7ZNtTIr1CCqoPsdLLKjf2Kj0N2m8LbmyUnq84dIMHDWzEySOKDY
txtb036XLBjVjs7S/ntUUeAlwbCXqSBHG3YCNfoqcA7JF2MeJwj91B1UsantKTR+
PGbb5RrO5OwZRoE4kJZq+/yxAybkH/z66el+ZoNSFNnPUvZm4AZKee1Jvk/6QU5Q
UQ8x4x0rHtsKK1o9Rn4H4kb6nm80K5qrI3MwZlQ4isFE9JJk+mQXsrKMNgqndCis
0mRLP5kaE9l1tFZ/jwxOlPB7ctMpmEHw0mHMQn5UdZF0DVTT5mg0A7lxPYX1lJxA
ilYGKhLxDU+xxcleeuLEwCttFO+Va9jrGw2RTF4Bs4pP5upUJKY+w1monuFbt+L9
qqUJeSfR0hdprIOQ1N+PqKJ+Uktwq3JYx93yPnsq84y5qkcSgo7jP/ecMgxP+exa
5BRFSRqP8y/GGB2ptOa0IrUeFmvYoz9Jz5fqBGnk4/YgHg8d/egv2UxddUocZoih
ovubQkKNqwuyOat973cyLzBPO8Nf7kHOZsShh3/gpqoHzheiCKBR3Ke0PxUMx5py
5zYyHNvdW2DUidvQTm0QTofMcp4Ko2Yzzl3ufsBwNEn7qz3qTlbIiVkEJQ9nTSV6
y3arTjRRtnuV9wbC0Gn1k4OT3bJ0RFAwIHDZCox6EBKzVVUB4nuwo4iqV0tryiVQ
J45EwEi/5NuVl4YfQvvK9e23lyCmQWUCC6dFqO/cF4SLpbxaHCTpW7dvPLpyLGcg
utPYenP6i/cBBE0WPG1b4A48Qu57S8Czu05A88N9JqA8t45VQA4c4offUqrs1hFR
TYrungDduq4G+mTDSJ1Tt1ZYmDg7KP5MByFINL/x4NQRc0v+CoVIf+D3YQlewxKJ
MpU6q6EYAD40m6KDqshGZQTG/I7T4oR4Jn/oh4LoUu2rRKjh09eRBMSkg6KsGznO
JMvTN3v3puzWNPb2U8wBfl85ItxEMlBa9G7QCfo+yZD9YI30AUgJCUR3bV6Anxm5
BBUdHiWS10cBCD50R5eq6G7ry/oBxDF3RD5J2ivezF/w8VZ/gQCBAXzQb4kXWTVw
1uk0p2KUaGLfehzL6yAYNrJftXC/UTY/Z29h/82Pqaybf2Tk63C/81DTyQVGJxCL
5v7p0hP6qSfqjSgDrIJRIY1221DxB4UBr182evApBvnhxjVPsL1qId/ig1UDGz1L
dMOlXvwFUYHaYJ1N367GuVkeyJrCNsCI2ZL1P2ZtryFqcORuaiFK2IOgZ9hEZbC4
6z7UbWw/9ZLOdtT8ZPKVCMsTd8nTSteGMBvTO/llhR9R6RL+NmryHcfFT2ihzX0c
WgTZ1CEAqA3wOWmPxecQCpaesMzutdutO4Vq0SpSQzaSjbN4611kHUdX+Kf1LfJU
WoI7h0pNgjE1r7Gaj4XSpTxbhNmFDdustlWg12PtCUYC36xlzlXeDQDkoFc+WP63
3p1qnjxfTrSJ5+RpOE8EZL7GZMTenYg5R6aonylUndLwJEPsRZBXgZUvzyaTNeD9
o5wMrDPGRf+D7mpXdjwj3muT0sqE0vwD/p2pILQrGt7Mp2zuQkYY+AZv3av1ItQg
tDvLGX7upZroOOUw2w6hNRVYusTKOKFn77dM2Xek/VmeewDFbLOemx4XJPRqBPi9
E784zH93YUU6JpwWHeSmOk8bW/Fs9z4ZmFD9zOM1chEIL9Qohys0EPjrQT291KC3
63hnI/EmfOmuR8UKcxR7ZG6lych0A58f/37au4/PzWTBoXFezbLdHRaMIsbwnAM9
83vfkEx7ZIIZwFGxKYc8dDjU+s1h+IKPzgj/iKd9c+GZhQJWoSn0d7NF2+CvBpFM
2S3yU2oSAA47JWMEXbufNbxsqvtRnmn/5aZEsVTQ8oY1S1htBLZxDwILtqQsFe7h
mfUHGkCl4HgEDqLfnmz+q30+e8VPa3+kurazZSb9PU2YZ9ht6yUlbJp4t9mQZ0Of
bEcAl+yAO4endI1H+ACucf+F5Lpy+Ix9RTxwXnXDkCExlAVLNuI/GKZkqtNTvnri
LNMKOfKopMpZgZz0oqzJOSFkenKLUbTMi7hsBy8UvgWeBFrGmoaqkwFT0gT+tBzB
nw4QN0F7x7oNHn2arhZcBQe98KJamUZpUVHIrRQFKfATAGweQfuFDWhyZwcBo71n
7+SNLNJZZeLoUwQ/qim0d39VmB0ombRylr1hsH5DHdOrbDzrZSF8MTXv2EKSv5ik
BmtdHJVxhw2za6mt3yeZbVkGgp25PYM2zimNJ5w1xsXQMiyKzq+rp3kHSaOeKNwe
0oMBBURmAWN9kmpVl+EPnlm0udbZm6jDtMXKrSM3gdr6h+R0hLJKwbQF9tQAehcX
DXg9wB6YzEF3mfXzig8njS0v0/D2I/hQx1Rx/ZvjUxpAj4RPFyzievhKe3HCAfaS
8urUYo2KEWQjJYOue/r9x+IBtXJcSOndrleL22sZFyZBl/fZ/hwUXc2HZvUoHFMQ
bptbiYbkearvlQPLg7RWus1LMhmOv7YgoiHr2pKtWr1g4Gw4MJXW42JaQHq8MaaB
0Vi1jXmhIHY2vcakA4kHF35lbkUl1NgV+wesZaq0RSFQcJW2eHuonMZfEEzz1ECg
rT4Fo2L3cJIULc29MUgP7wRN4uLHl/pxe9mzrRJ5XVL3o45Zt9wolIjhs7yd3iKG
dAU1srj5bAWKhOoprsNqPmrjk0BXoPTwzPHlJ6M351aqTFQix3B3vNnqb23kS0sC
gGG4GKd8hmuHP9wV1QjgYDJpzaCNeWJfaItlCa0KIuqkLR2xbgLJys8mfkqaE+TL
zC/w33hTN1jP2lnaREeSFnSJwclls675kT7foINLqoInSKoKvd5GWGlT3W6e+g7e
RUs26jl0uzgDUUDcwdtdwZ+3L4TJyId/8/i/AubYf04tHckmhseDbr03BVwbB/kY
u6V0cTTTIeT0ws1UfgTV23lHusnUmXS1c09mtze/+TK2pIiffTIIMv8Q2gh0c28K
PSdpnFeYB2bhsAV+piWyihWxVtwo86X5p1AGFqOlhAHckU7NuBdI6vPIpR7s6+eZ
TezocVb9HVxpEeImtvIBsRt4oHpxzXX/RtZrm9CKJHh2WxCti9W9cEetdMabiuiw
5md3So07aLP+0IeBkNDa0hGj5wz0BS1VZF1aqRPSwBoTYR7q9qQPomVgQNnII6Nw
+r9vjwDXesR1hxvaEPbLazN5ZGoiD/9QTztxtzX119gxuQEHSIEGtQZyT5RVIYx3
qSW3KEOBK0+VZ5jUVP/YfCHJZgtIV/cPEgtQRxz+YIA1tFtWjGcPr6wc1lL5SrqF
XJtUeHWnKGsmxQhSHx6RMQoGzzrHLCrDAvqcJMKM1mUllO2BdOdPCLSld9s1z7jB
Gd7LBmq3fSlmBCPP502iBbFLzYL2sZm9FBOai6tSjinp5OoULQJZTfwLcepxL1Ae
BP6dC51Ldz5S/BM1t1Cy8F7yxTjJu7kYl/2zI5UyfaU1ndl2MJi5Hy2hY8tEywPs
qKPrdm5qDcOvaow5N3UTkkVowFWjZv8snG22wPDbYE32n0+Vp1u+Ic+IezFyE9dA
og+av6BuLZoCtla3heki5ykXMY+LddhRirULenZ2EJVPfZ69DYvCwl28sOrMKaqB
2CD4Mnhs3qitI1T13u/Jdu6uY3h8WfAxmJGAc7CxAV9Hlw3Sw/73hboq2iCixrnW
22BbNoNY5GwgInEL50Kxhnad/5CY6jQOJVZyhZbPT/K8lezeLOrK63sAUt/DSOS6
E9iyxVIJ/66dXAWZ632WCK1uM0g/ugOY59UdSzrVYov9ZXhDIWEBPqsuyUxmqhPa
ac+FPjdRLMHms011Q9OfXFl3mCJG17mTOYPL7cABBEXojTjxZDktr6tTwA1hsn6l
JVE+U2x4UXj6I5I+Usqe7j6UQGke1CQEhls+n4pPeBHu7TmB0Sp594IPoDfqFT3E
kzlf8l0sLrwgzeNymBL0PZdW6UzWZVQsKT6tv6pSJ01nBOj5g2hrNvHVyvK21CPF
6ZzJhhfWKLekXfyAgAoG6RrCgAQ81M0nHkCzhEUm9cqwVAwiNVvMf1LZHANHD1Gn
If9xUccWR+uyFIONn1p9Slx1cWvYMFifmm9TlfrMtPJ/8Ve0tYuGdMLXZh1JaTq0
Xh0k/xim+8i2XrljZhvMffKPO5UYWjZfeLeGHTVYWVoLF+QWp/MA36WRj+7mq8Gi
XdRyB0cNE5GSXMDCGS3MdqPXuojNlZptdpMdWbkdUpoi5Gc9D8tKOhB+pPmmt9vK
l+yD565K816bHJiHETSWjrCoeqMTjfydxZfJa2Yxq4957W0cME0Sgu2EzeUm575+
rzf1jhuzzl/WaZXJpu6VBsggiIoojXoGMwNZSBnnqFHqvON42NApD3pn2c8eUjYg
IhQ8OLszgz9m3dxprP7+vtu0FHYliuNIx96OHCbgAvlP+LMWYGpCbbWUm2iw4KdL
AEkd5KNj+Gc6pZIWGGqNhSFarh50FIWNm8PQfUF7sRlOApFpLugBguRs+obwSGju
2ipIS13X99CQOjWdNLeYqZZGOES0HUW8Op+gxyTfC0BCfeBRLSo3pOXnFonzigr0
eLCCLGNVQpnDQNeMTr/eQUdiYAhFBWZEs/3OiJZl1I+NnVjhm8SqX/Tp/+eqeCmq
hZoK28u+Lp36B0BTZx/sFss6sdS+MO2bQTJgt7hCD72R3CPmuwAIdRXYlTjY5m02
ii/VQlHTv9jk//AeBZAildjVBJ4ihvxBArfDjIRIsgiCgIogXpWjFA6luODAu4ss
3aq+SaK2fqd0OJ+IBSWk70rjQPOJIFF/0UNPLp6OX8TIB2cnLFb/mN6TEj8chMTT
g8iTRHUle+Ue42mVVeMuWRP4L8n3+6Sn6iAahebuU5UL1tVKNY+dNPP1nZm9ZkDd
2OW+i+BKksIdWyQP9Sk6lEzaBkEn1ivJnJnb6O3g662U0cAdbhUh02v1GmTK0lLC
TCxMHjU7Aqcn7xgUqptDiWrW1aggUAVc3jgQbP20vfsjq7HyrhkwnVq5l6Dk9ax9
BGDwq1G8GRHw1wjuKHoiWW27n4ekAjGBWDmCSP2hRYOLgK/L/7IRsQTlIBUYGRH1
t/2hHhWO6zd+YCrpZlnfxYuRXnCCck8CdHiCdgIMWPft7yecRzThRz+uaEEcC2Qk
U4Qt0xpJ4I/Du9XX+e3lIkGZ2Uulb+f+M70XxoQ/DyEqfFXxuCukCN4+9elCCqnN
pANLtvlC9sW3KekYXrWzVx4dNnGcEaFYZKmDRcwWOl89QuJhlFcfnbOj3loXTuHl
QBlDIjpV8N1kNR4dxY9aDFHgZ/8z+UScNvx5J8GdwgIhym9iMiO/N3CFXYMBV95U
hvkb6vw1w+YU5VUKEcj2feXdxo9pBwCuVaNGYAJHpUe9+AgvxwZ+PVYA9dCPzMAT
JRKKu+2GsHdh8nBJhQ1zs0m6ddQy/AEFDHkObrhOIkayQdECWduEY+gLYttPwbxc
ExTs9u4ACil5+JzWuFnyyjtnampxJH94i32ql/w67m0GSQ6IkBPNZ5I6yqrIX1Bm
HJ7ewxaZQ5nAXqbuhYy+tjMzjij6eZ6/o5EFPlJgTdzM5GuryYnCC7zyYuR3HjE6
+AON17xl5QAL0pJygqpfqessuA1574MoXKtPmgx1vOnTXIQhADj8v7OMW1Tt9ipl
zBWF7cFwUVV7dsbgj34S7ucf30XrKpuxzl9yh6IfYA2iWnGtRFF2o4rE/3zSjcqd
J8x0ylih30H0+cwg67VSxQEAdbqSgiMpDtKdzUWyZ/Nb9TXvHp+DTh4Y/Hhvh98E
kBhUusPc6AA3N2kS9oFOObJTEZw4YQMBeq2btO5Bfre0LXDkaY4Fws8k3jq+AP7K
spxGS4J2MlOZPZdfYwoWXoNLswRovqIsAKHmFpq5WvpUHw2Jj3zAc0z7UOOs6KBl
qSpqOPC3Sn0reiHBJ6s6Z7dFYho2KdmubwCpcSH9UzkUmEaTbUcWZ2Xxq2+tSqe/
8x3cgTPxTy7clir4U8WA6HBrGEQlUhHZ1ebP/X6NIzLr/CesRCP7RZW7e2ud6SBt
xlQ3aMX7mzK45u4vjhRTYzos+FgRbDJSm1d6rOp28S9Ge24b0PhxpHtAoWWw87Eo
16MNFOqmUWPOGK29cGqjp8wiexZtlqPAGICg+4hYI1vlA2eea8OLmIHG2dfsYGzV
iKRgICIV1CVpNDu4901iH0tSuMJyAQ0qMy+SnYY//Xbj3BUnExb1UM3oefLV8S9V
EifGUJ/gCHMxr44x2HhCzqYv+S+IbOVqaonKejQA3TXxFgwm6WO43+o8YXjSGppu
KXFFNRUVcUKrGf3eJKp94+h76NVy6NJfz4v41beLSzZ9dxOMRwCq/ZNgdAiDlSRF
Va1SaHUXE+iWFtFCvY3njtg4WISSFUytMv6aRhtJHTX3xoGikyvV2PqN5nz459N4
EA8bdsojXGF1uvY+1RDxoWE08rf4SsV0GQnzNxoluqu4k5myiZhxo9e7NiF4n9wy
FE9/ylk6dvtP0WkDjH2N2xA36IJcq8gbBX8bQlHlufT1uL6UEUU3TAcf8/xmdSjj
mEELOAMpheQIIEpjeHJ0ssqlDPsxIK4IKakKQFlSQU52LkCru2hD8oWN5YQvxcQd
RFfXxkpW56nXLbBISXX2mMdEPoTYa+vdhzD36Q+T/YK+3En0FB1y3DJs3IacNa2i
aXaxex1yMxrBPfD6Zt9PWk8DF+dhd7WbeUHVqBf+QcWpppfWx3Qr4hd/UQNjqHqv
6NhBkVq7pY5XpfUz2vM2s7cfx1ZIxyMnYqg5QFNj0D1rBFRtoNkA3FGZ3nu1mach
Yn6u2wtZ4C6m2jMsXY0uLH7jcX2ezlawkPOKh5yWDc4VWKy7cYwxYWWMxXn4y9kp
JJxI4VepLVHV3gVdo3WcIFTC4FiaLWSRKO9WosL2I15bvMVohVEJ+jFrkbuUMoNl
+is83eNyL9pheU8a4voBPsvzdoK9KLGwVk//dwgZmLi1g961IVndbnxQkE/9pm4M
Kh2rkCMuky3BwPufIoVQSolqaI3busN+DYPwfB2ooP5RCOFOctoMHvuk6FpR56LH
A2oXUIvbyb+gSkV/dEgElQ5gJBABFW/hqom2YJgIrwGayAkmi8NzOf9/Gmum9rq1
wmgT3fxUxTNu9CWjw2DnR89lU9doS/jcdvRXZcB9WLH/srOIw9B7dpoAC3k89h7v
QXrbRfQ8HZ/pWZRn5/YFxvkkxh2qxprUrjr9FdBdCoKoYf67gWmN9UrSbOxyFWqC
yX7cWpvoaDmSpM+H5uaLQYo+nDhJe8lVjD1FMds9oGyNz1JB2deTm/q3ltBJBXSL
EGYCpKLxyKa88kOONbuCWrrssUkl1bm3cz6ab9t9af+bxprGpWiUQezpnZ7Ss+n/
ZYxxti3OA3u4ipjs+t6YcdpfISDTWeqXh/qZq36b68p7QVbNXy7pcnaLGtOfRX8D
QJjzWA1a93fPJLOhUrXpzcuhm/2cK5l2sG3S4T33w4vqhGmkLxYIZEY6+7q2MvSg
nm+PPSu7pzaUAK4n9M3m8LYOJkEveyvGN56IT+SGxdXkbkbHwcW70eKQZvAVBVeX
edkyk4J/lS29VRq467/OSnxCp2qjdm8Pv3w3FvYBfoO+H6MN+KjOhFxGUoQHBDht
KqObFnl4XyxWwo32mpiaIeLAmXzHc4yBPr6RHa1S9bVIDdCDcqVzDmOeFJd8MYrd
n+0wpf0KXNbcpnpdaQg5MF0XkTlWsrdCcq+h93PeaZhZBplFJ50u7ixcPbGqJXWk
KIxmAEMzRzCbin65p58BiOJtmlreoeixiZk+CwQiueW8H4AXFgJGQEc9Z6xWe5MM
WyfTkLbNKjH2HpaexCUWyP/HkV4bkh6eHOd+gSnCU5LEfXT4kG2VcaR3oJDJCOYa
1W0aNwzTPJSALIDlDToxc6U0bjY8O2GQfceAEpW5TpEOjjE/ujzwYBJdbWR7B7QK
ldR6TJsCRcHHCRThCeEgjQUYVAT0NVsa/Otn3DUH9N2Tk3kz6mhWBbgk4AlZBXko
/qeafpOE/QnjOInJ0i9RcF9ZTJBjGLyzBfWPPVzQYwEt5FHuAZBXJKob5oMPJ9/w
RHEOQr+lZ6mbdLjWzeAgV8r/cNlDDIJCt6prVj5I/19ZUOJ4sDDiJSw5X4B4eq7k
VORNthORhdrp8byxGDJ6tktI/4/gqYWCfff592L1FGBQhawjmnjjr0IR8XyBDPff
1rPuvanGf+6Zly4Jf0BfgvINwg6fNLWte5h0l1f0c6OOdx5faoqFbXOrTua1PPDY
YOsoB2xImvzVAj2ni7zUu4tzkGwlU0XIADCQzrQDAUiIljELrKQWtEtC6BJUERzT
JtPyNAzn0ZZx6oPzDcLN4CPfeEC4Tf8QAZmQuQHmpXRQJ0oH4o3JlmWDIgUngIg8
HxGN40KqTpdqvk1nJHisxEb9c/fKAVVmNcAmulbRcjqxx6LZAErAdyGWU4Fe5dya
i7GxTD6EuG5++Z4/4GO0P358fTBlcJIH4Mxqd1rPQ1nEX+SVXWOnd/2yS9HTs2HG
q65HTgcdL1c9BjTDVyF3QlHzzAmx8D6W8rVfFlV48et5VQTkYno/G05rB0sWrCpm
D2g0o9arns2r/vG+1w1Gp68cb3FCGtyMkMajfmcgbSu4YVLeHW+qtIDgQ4vgFJQ3
8RrpKmFbHwGJ86MVxURX1CDSv0NXiGYdZTPrcusDxLu9AaUePyNWSoiCF8nEySjs
JUA0zq1Md6ZTJFsf67OMbzVoo3Kpfr3JvuXea1mEg113XueG9SjzDJRwHKKYcxUa
CpTpGobp6hNvs7ptOttr38IPie80+JMi4EmsPK/1StiYaM9OwDmsc0YJvmS6eVf0
OzMiXuRoa8ZXZcDtE81m0mNN8vEj15bwZHIPPWoYMl9DhAmt4dSDUZObHEv2Dg9c
JIAnYwoEBguNT5F90jGp6XnJSOvy1gwqxGDXeShFJTgIcSSWZBij6PJ4RbLzOP/e
Fxz9Al1ajZGr+FbuBiTkUhNA1fb9pRx+UEDJZTLf01O+xKKoacGUDa0Wg419iAu7
4WfZKiBqkNRU/plG7SYquBl61gZWyFDm9EjTGv52+16GbFMB6mB9xwofcT3YEpsR
uKF5g7B+FCFYUyEt2zUCXZHAH/hpjxv3Rs/cGHpegLouZHQoCETFYIVpZt4jJ64W
Uz0c0y+UM6SiL4UrC4cWEg8qxfHnSbeymHhVekq74Kv74KKYQb6uoXn7juMqerD9
jsd5+wKh46B1728juApqwnvtb1EIU5ngqTiIIZcEFuZ5eSo34sliOIeyoQDxWAw+
/DKrb2cZExwSArfAITpXRn4jCUUgCGOm1h32nGXiES/jW5XZcfWvJYmyJZbD5Uw+
WyFmOv47QkNTEUyl3/p9YyesEsK+2NMRRsRfZu+GCjgLTkjEDNXFO0ngDTHg0niu
QRN3Twt247Mpjf6/HIrbdGoU+/cK227qafBgJzphasfKpKXWXfH/Qjxj1Lu2pkzK
6XvsQEU9NIHSsgkP9lfYC4xV2Tf5QeW0m+bl+2y/QIf6Vb1OI4TTHJiq+v0iyEM6
LjL61hiIGhFsBHNVuwitI4OaVxNTfti9i4RHzyhDcU7u1a7e4R+2F0x6/2Lj5bGx
PaB5Lokbnck7iRPaTMCbeIUVfG8SQcAFZT5O6hCBUS/NFT6ESok5MYvVIoqf2WYF
23ATWTlpWLNq87SWGG8r6yDpwBq+c7SpMYDDzcFozN/JVuj60bW/JhpihZC7SjFY
2yHXAKc+LVg3rL61vimaH/QWTFYUDAIvtV2uCs/UF92/HwuGPoJapOP+WuBuf0BJ
dQdC8yTbNjb7RVrnrp5jXj8pMT5G2sq7Ja/TbHkemEBgeTx2t3nINyklCCClRk1q
5Dbrm67f2J8rwZQmbdNORfVjRLGf4NlCfpWDmq0sBTkJN3gUt+58ZRZ5IBTXDLeO
0hQnYwSeUy/PCO02YOpqKccbp+IjEvRdCuWy3WaVyUqG/p3gRAnynsSqXGa+bxl3
F+aq6MzGqTziKiHkmy/ToCjw5/35lr3AmmrUEWNKFhkWNSsmQvmB5Jo8VpHM/Gz1
xAH6uSmnEMHZTUuNNw001G9DHolkUWCaTaPl0MZArfebBPF7U1xDilWyh/ZOhWBb
wEq/+W+ix6zyeO4JgGIMNZTUrj+efmRi1UKxs9C8ZMI5uRmmr+kMeuJD7U+N/aHr
XHGRYc/7+nJOd9VinNkNImoHNkKVaAkSSy3rqdcTNQZZTM2dkZOyH98UATBSn9dj
pqn0d2GuEr8yKjGPDGcYIKc0g4WeVLh0McQKYHDxQcvB4xTSzUhuSooEVX9argbP
GM9HV7BXQ2sWtLGwtvZcSq3tTjLRdn1Lf2ID6G5K9wRyf72w13y45VQ0U0Qnb0IN
MNVFb7VCk7Z89Ai5nNEtj/G1xZJxQ5REZXDuB4bWvLSiPDKpf5t9McnNGrH+Odp2
Rlil3jL7PJxDDpgde7QmkjcPJTC9mjRiCs5EpZgCAnFhtiL/+LsNhIsTeS49vzmL
nLw1M8pz/hseOQhM0QoCYkgF1AhyQqH4QeYe9f7YkmBf6+qY0XBkWU9tUTgWlCaG
j0HTGWcweOVzZK5q/j1BXsS3sudDTfFU/AB/oSQIiAVSGyw9J7ip6zOQ9XTgzqxB
WMIyldEdg7x7s24s150MM/V2y5coAKtBdxG0D2wxVWpmA30noJ8XdpvJSnrpRcZK
Cxj3vUZ1wzUTzGUMAV9NlI0IRiOaH7Q/JjR9Ed5POR6NcD+AywymrYhXXyKHw+72
rpiTMS8ZBgFEKqWfnBXPtye5FnZ0eTjGh94biCPKbC8t/xpFe9GqwaF0abdjED3O
3oAVIJWriDhRxRVLvirdRv0WXLGKhGnvt7oPMYhMZaQx8+DPpwedp1c2vqRRtQxU
BbskRKJ0qKQ2cq3vkmi3gW4GFGPiAVUaYtSjc0CrvSQbWa8UmWEf3kWH610UBoz5
FbTtfaVQzRPXSE4uMUsCg8iywH6ZhqgDSOTTD4DDZo15/NW0oo7Op6RLeAtnokUa
7R59A8GIIdydvDwllzixcq+JaGSEePMEJLKxgoL7DoVG/0NfeEWZ/gLSMW0Za+HR
wxV/okEOb7XV2Wu05L6H8XFnEeN4VeSOqF7KMD7m+a8KF6QD6ZIPG2OvWJ3WXzUM
frmisSxGavqVZ8TvKIs96nRvKO9scm3BGVAStbg1qtmBrdzZlIMSGCC4xgYkNdpL
SbTzNTHBtIViUFgya8ZU23hco0WLttcMrFOJ9l06g3ea0c9m2uobcr4nowixK8dh
CDZYdRayYwp/aPW3DiBC0QThwmXFZke/njuY7gS5Acj6n5EHDXU6K2xRP6fV7Zgt
sMmGKC5IQKE0qTf8nYiYydR7zNf/rQFJq98lmWeGzKd5bSCOhbjZuEKDZReJRdy/
rZCZtr0zNUVKzP5xmob+V2FlfjHBwAYp9SDi5gXehnhN0urXalqBBBb/a8tO1wB5
c0JUdE9IJsJFJFmjl+mS0jtwzekTquMEdcGfj34mSJTsd0T7vArdRQjrOGOYeIxe
drgQ2MpYO5Q8ow7nqQ6BTU/TDg4aQtPpQ89WFLR6wiZujJ+1HwQz2vRPt4m88AmG
0X8h/+QG2DrQegl4pWKS22q5Z89r96BRP9zouw8HPgUWlvp8ARvUvkZlyiSKaPWV
hgBTPj99v0N46kd4QfMDLQNPBpgbekdQDbxrzMf8tO+3/8zWfUZoz4+uqJ8ENVgx
MMozncUGWgyKMstUaLQ3YHoI7fIfMJTdT1Z4kpb92otFhrEPMxS4FRD6Dcr+Dcro
GIO/TXEjH+tw0quv6J6wzVhngPS/EWGR7g56JE0gQFQDpJ3U/RWlTIIMmhwhPOEE
BBk02uerirN3kfeFXqFx4rwW00hyDgcrf2FoNgngH7NvoPAhf7sL7pNp8YE3g88G
iujSlrPN2UqunIB/XMv4W6QwldfkXnfXqFNWJfvfgU1oSb2lz5o3JrWAAuBOEShG
yJwveEWRLZRE0ZIkmZfCCODaUGyebPKEInX4iG2+DqMVs8eXRSSPo7YYucAqU1En
gjwcHZPrj/4vkC8YpbBLu/7vx2zXfGVgxVUjdjwrrrIGgMEM4MEFhbr5RPHKNOFG
CpWnk3oZFsU2xkKfpr5husBR7XeNN8WFhb1b95g6zCw0N2Gqci13aK0JsPMKmKXm
w6qS04KDWNFvBZBZxneBpW15RHXi58HTSvKrpQ3w0gudD3Mf3yUYzOGGrtU3FC2g
TKslQ8KboN+FmVmPU8iLpa87Wh6KjW8gdnC152svTighi4ma0ay9NxcqtykHdWlC
nq6uOZc3fQ0iv6eV3bnhr/I5+x5ys3cYGOFtGgTyBIOMSR9ek7XaeuZTLtEu1ALd
LkK1nt4LPqNFA1t8wO7gI0WgO/cYKvUdrJrQZimk9H304LkNhsodhETW9UJepxZB
NqgT9Z2OANh4FPfnhCjUSv/LG+WR3HR35OIyE+7c/EZ4cFjb+BRTNWJEZVb+5U/N
n2017QdaYwUOQXIkARCz1mzOEhuoa4AyTqtdOzNMR6u1CKBZWX3VQt0VDR02x92K
N5e/G6NyWiZ1MyBsNZiPDOpb1FaOcqDhAMRUjuKATKEa8N/wguKNdfVPrTse+Aen
nXkgFp6sMlj2orr17JDMJ2vuaMRrYXAzCNMGI7MIa54u2rBzUL9Tvvkk1X9VSZ6q
jjwDVwZssmD0TGo/68g8lgoxQiyW/LOk9+GKsszhd+fi12i+A6UxqpiKnAQGzwpQ
3VdPiTAVpOvltSFQKd88Fu81gBFABrcPnIwc/bA6Q9430Uadl/EuenYbFAYlqf0Z
7Y7NGFZDvGkh8TXfCh1126nhflILXpxJ+V2ybyOlTQEMwWWURPnaGrTqkrxT8Awq
mA184jfPm1MvQdybsro9319rIt8jE2Fyp/9SrN+n5Nkpy9eJUEbwtwp7c4cYY+9g
u1j/fO/ZeKnoHPLq9QgUsXS/Mecab3TwUH/nsetEVjPj3bLbZUMR85rUFHJIbKij
aCLlRtyPv6jE6Ob3KPNyhQ0YVIOxOv4fpCF4zntYQQFI9hCLEDYQ7+8bYz26nfpI
IDgf4w64JhE2xm3oSV0c7NFCWUQHF4K5KA/osjgs5ccTrfEuOLjSv3FZZjDxOqXn
KShClrhetZqLssGANpqbEt0+kK0keEwS5UAcZn1sQHrWizw8scvBXNZuHp2axHh8
bvqSUGwJKrw9dQIC5Y8HBKPWrAKsphwDPNXLhqLQoBI314yQFc8I8JeaolKf0u7O
6p27+XYZ4GgN6KWFbYTr6N0fo6XMaS/+R+5rjLjYpjSCeHAQLUXeIsPeDS3lVYcB
qsvVr4OXTkmCAm42nv0r7lCeEzfDIC5Lp/r8TpmOPGn+5ilZykiJCDNNmiVOsnb/
vUcGdtIqXzdwcSxXUCxTspJ9Glw+DhUuGym1JZSNpANLL70nDR6wrTV4EeSGICU1
UTnplXu62Yx9sXGMLsyKOqycOmYpb8fUvk3UkS0va1b7VeLdw2WhTq3/sSNF8TQv
v/oFMIWZOWs2hk5nMYGWqyDM8E29xwee8FNuv6qyrWxbWAZkIBkuraiNne35aCBr
HCorZx7v7FvKflRuMswl1X8Pd+4NKyzPEoXyZotaxqG/RqKe0evtv789TOR9+yt5
sZ5v/upFM6dl7yhprW+gQvAys0Jtr/v7FM1DFK72U6bQLpiyOLQgnRNoF14cg7ac
LgJdd4mQ/kp6J+7kaZ/Cj1Rj7U7DAuzXqb9qVMmsgXOpjXa0eohD0OTzM5067VU+
tAp0yhSUWdGoLEpHZExRqaNBxNZ7pBhwlLckY2uu0bXvo1GnoCbMU6/DvZ8qnVsw
1LXhHVBzOly9MwslaDzY/SNS7v6Dmvx6wj/WhS0pOKy/4RLlXe4El6b//k9T+RkK
b/4fIKOm4Xq28SCyA9XI42P/8aZm+xmLTtb0XX2WJkezWbL33PMCyYJt1PeRJ/I7
pTXUPWX349TnskU6zsUlt3/BPF83mxv7gD5GL8zjNSc=
`protect end_protected