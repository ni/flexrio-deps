`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 35344 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
lmOQgIOM5jiJrGbWpsW/8q8PDtkiOLeqWQzJK/pqHcbSP2osfR2PMFctf7JM+Qog
weJLSdcKVQgGHIC2x8Fphk84zitG/9+PMPa5XQMOnEtSYfsVLrM3sBtMnZNMkCFz
bn973PUNc1LoacGk6brQGRqQFDg+lDaqHDknLGWnJ0kahvoRuPmqkQncF4aoQW8Q
YjVQTw/J1pOVMEKJRe4NO+45pCgk8p9chmUKCZZYNKtLescmy9ggkruXXPr4ZdZ3
zA0H59HV7ae1Uosb4HzuLZvH82FPWajnqD5xMI2NX6gtSJHzSj0Pu63PkOQlAogD
+ml/s1Z2BIPiSq/EcxxQx9NqA2I6rVa/0eSrQU1VdkEtyaj2OkuBztQNydBuOXhb
YPvonazyeGtPygVtXYGaxDr3PvewXeUWa/+khayqz/vyuZ6FZy+DYp2tRsfVk8n7
jevYU7bC3a+A/Us0/Nx2C9b5K9xDd20RK4l/TXA2Cs5TXidY9g2vZPq9nRJHbBIy
V2OkKhDtIjpwxxlXFgdrTY/aGXJhJwsOQ0PODdj+2sb4RlCVuG2hhww1Vl0e0MhA
HjEs78BxbYe1EUK7b4yEBveT6D2XVfk7ji6wtGolRwvk5eGSFbwPDO49lzDUMwUR
X6KlPmSGaLy5qeOBdqFKG8wrewA/a2N5bkI2cWSTDlEv1n4DGdjKLwSobfoMN6x/
/2aLMyMmkwoXxmfZIS5R55f58NUo+ph+mMX6DlczOuz4hKi4LclmkJILHFxQrVIU
T2l7wLMoTjROq/MMiDWnG+aDK60trtbfuWRcRWsVWEp6VrtQSOyQo071AwJaeRJL
BU+J7Uym9Q2y6ciCm0ucaq0o7LwhsIUqGavSO7fs1gVUV473/wyj8B2LRc3gP//4
zk9DaR35UV9qoKyuZ9wBYy9rVXY0yZ3kZMafs3dD2gPUf5zlTFPok98f0zJ3jJts
OOq+L1pmQnMAeqX2qwOQ6343kWBYnE8Fhzij0nzaaOPf2Cv7xPzrIrQikJITsSXt
tF9c6V00ucEwaIZy+6lbkyd+yeyyCu6ZvGZ7eYxPq3hT0ANVnxBBKZl0RGUlabBr
vPT35LREwYyn6WDYvENyPf8d/SkEoOuidG+ZF9CrCt1FOUt4bFPhYjLyS/Tk4vqB
n+9MsjQnmvTggI4UlDiq9TVxFfCLnTY0KbyZUFRIogC4Dh2Hu3JtX3drVtYb04y5
hvVzjpmt2o9l/o0WbbuAQ0ZwQ/vH7AdNlTMKU30+C/TyLUte6fXgGjhL2d3pFHTf
hJ2p1SQCFR152Jn1tzDdRL86caT+omzvf6p5etn5wyGFwRqhb86yE2XhKNFi6q7a
FLLA/guAohvoSpaW1xZfZb9SI2GHyQTlcjyHt8vOeUxxRQqnZ8QL3YckMahtBa5e
qqHJ6/oVvF0iS5fCTH5NZBC5u+C+RCA63/klwMxZ7B+xOW303XcDv0f0aN0D06DU
XzhVgIG7+30oNQpfPWIDlkLbPNPcqKoLz/RRAaGNybOawzjY7NYVWAjZMvbxRDHl
PD2rVSUEDSXO2XlRGAdJdxyvg8y9KKz2LFPvpjpkrMA7XcvyUsZXzpl9OZXTTjj0
DJq0mnSkWxnwwsB4sUdtxL0/PiZsAm9zroCvJd4UumgztBp5xq5sEG9x8rLS7R9S
D9O8b/+NpSi8Bhb0jAjZ9saGrx8b5scB+XN9Wmack11hTcJFfSjwxqcVtzxTHrq6
Af7khLdu5q0FfWz9yfo4aUxZhJqLZEqadq7vU+OWmyg/v0jS3tt1DK4yO/pmYQyb
+id5l7CeoMIQDvXfrvYCqCcGAhSB+Zhl46VH0csEle8C+9Q4CYpQDlk7nWFmJ7zM
CLHR9knu/g5DtoqSRw/ucZTZ6hxvvw+LAhKYvkuARPEfFqFhb+KfR7q8Ffa3Muqa
EgQplZfG1OMMWdTLagdhFJH01C2ccUVQuNI025opAVuoV8FEZHOCARNyAmJ2KEgH
LCYn3BdGeaaLd4PyvlDzYvFd2T1SQq41SXaDNy03vYMjR2XCDpqPl6gs5R+ojttX
ebw1D+lVK8/7Qp6evYWXqzodkGkLvHYpCTh7Mjzz9qoGwQzMFJ7R/UQJCUNC5Al+
jckZNCz24rjwwyO3wwoLq91UhMXC/w+oXzGymTWk0dd5LcnCdt+v1YXroagat2LI
XdevDNl6cOx4So/Fx0uZ7Erb+4axcTygEaq4txyp/dniXZFR1ti7N32j7F7QTKxz
kNYDbyT9Iqvtm8E02BOQRCbA6ajhOlbE+1n4xUDq28o2t9M5SpDK5satGGRiSZRf
BBdiSp8TItH1rtZWt2v+8eKyp/qBaabwhIgiu7uvPhaZAIBOp9P1Rx7Y9EPEAqZP
6gi2JnDx08OGcm/XFsA8fDueDI2adPW9Q9d4pfVtQ7VQUhqjnXb7MlMkZRrpJ4Pt
kRyicRfvCiZu7+ze+JCypqihWgkr4+qPCAsxalHltIXSj/vIPV6gYfH3MRsHVyF6
4sPYILmszjfmMrdkj4vh744kYQidXGRKetdR0ju7VmrwQqORs6l7JQ+BbWMJFfzp
h+hotREASr9CqYqFwJSuEveBmlyeIW0ckMRYIWKOUxzbWVVQEKn0/a0FRDYCauvV
ogBLN30WXS2CtKWTbVaNkFI2y3Ba1rmMJB96gTT3eZmSOCgMm3dWOfb1jB1o5bWU
c/jhOyqCYDJunECgKfR7qWS0sSkfjiefM3YhoSIYeoFaDoNMQu//bhdB5NPsxpXa
BlrHUHfZlJnRV2Z+y0UkMl502z7wHq6qpT3rWZAIEnOR+Xn395VDcGkMm6cTa397
9bT+XlrXBGucN7gGRbdOJMsrTNlA9Q+3rVG3n6u3oxCx27czvmb3noq1nFFypb6J
MfBsUgGsI8ZtYxUFylyrBhgL4y1kmAFjowip3RuoKJRkVJUlbLnsq+Ai4EXdmqAS
btiKhCLEv73KwcMKWE9fI7DXhIJWnnxFawNtK03M74oW8LIwuA1tjFe6+08aRIuS
/1fQfVCwoRHDOL/mLEtCTjkiUyrF96yIfBiV71MDga8BRj6n+AUczN29PJthstyJ
zzHM4L53u6uv6OMFzXy7eI5mDv59eR6OZJatrP8xGSqAzELfUu2ztQ3xI8/2xGKP
jq1x0a5wUdCISFKOa4xkHuNChQHIwMUbUBzphas9LK3zqdzlN9JMVVWuCbLOkY3J
Q4S+JhWm5Pn2CrG14a+TYtD/KpkwwtS3GV+hWQ4apKdQEeja+ivFqqTkQ5n5yU2D
Xl94HwVV27NQJoPoBHXSnBrP+6JtjFMttydIym7W3UGINKk/IVM6jRWdyNDnsZHl
TlGtzd9Uu9/ZWeDFBb4S9vd6V9X68lfRHnnNXMBoN64qTaW4jbK0bPIDjTrUv/Dy
lUaURJkpDhA09ccJHGf76yQZzE7X8eV9MvZdn+2K4jgUyZ9L6UlD3pjVZufp0WXR
XcFLUPLpMuaGxBTqb9u/yl7Yt+leyjG3nzztK8qDFvteNfJahs2kHtP//RQeCqLE
o6IRdBED5zJ75qZQeXgc+2zr87HK/jgjIVi/Ex2C0x+USuoXjoCeZfKr+grlyIWi
OOYo/uSMsI0pSDXBw1P3zcoL0h/hbzIsf0OvLczUpsTJs+nnpu7G56wK8DZQmf39
bTOIjT0a8tAKz7OHq9v18nJ46WF6pCl3OKbqK3gR2/+WnBFZerTfvV1MRs0EgiZx
5xu9Qhp6RcP9yR3JQf0AUYYviMNNdHprDIYWd69PoDbY9EBYfm7nptR1SQxLEesG
Tdg2TWbDflIyjqH2mX64GzoZJABkKqAoJPjIy5CqHTRJTcAcRCTfr8zcbqNGjR3o
trrz45z2e/I2+Ylu28makLvccmdeOEvSD0CznN3cslR48Zf40JcFtVCFF9Qdjbzh
JjP7WP23NSH+R7rYP1cwkTAC0rL4wBbsYf/9kKlB4egh8FEVIe+oPw7AcSuZaIHD
FzMsIIG88L/AbsdSXmfzfLhjKEC0ZeKOcCx97e1wzdIDpHT9ouY+Iq6mKGfir7a9
jMD9qzkQyDfpQZ6NWn6rhxoiJJk/M0m7jYFTBfjpODn43v5YCKngEi1UIJ1vK/qQ
nkYVSlF3Z/E6iMC3NTwTpD9fNAlbJSml4WSjHQCPBm8OfOPs0Zya4CZNRt9aZ1mT
0WlxzgujEOy93wNYKCN0eWb5X2NydSaPxDe9UTrUoGCywPSmsR1pwcwz5cMjmJyU
Klhywd1mPMyoDEz2bMxYBlYWipxcmOtl4JspYjGLE7nGX746P1vX97Zy2/kt8B7T
vonaRg9PWMSKm+eELKnGFSRbiVpFW/Gw7ET58nRQmmAr1SslVPhMq/cB0EbaFYPD
WVa9MDDK5p2IqxTCN86C///mk4rCiVSA2oI6pprtEBmky4ySV5s32D/+QUkTwQE1
Vjv/PZX61vB1+WYh815bPECgXczf91FKJbCalkX6ZaKlKc3vDgSNPBKN67jFYOff
zpltuw2KKhuY8fE/vOlOr4nsDq22bKeBz2K/uWa9a2SpPUofQ511Wsi4DZLhat+0
UpTTzd9X2WGEIWR12a4sFRNygsy9oUDebT0GAkKn263+FXfY5r8Od7iMDCKZx3dZ
9dXOxVa3lDeM/RBl1xn6Hj4knGIyS34Iq0iU+4owBX3syzpgBGbGiQn9TcjC3QB6
51Fdj4hWo2VL5k4JpDag3i9KyGB00F9jIIx0DDfjA3ekVp1HZx4B9zcEhGxYw52t
qfGtiGpvH3PtB7pBm0SjJDRsCkOWdXrcEEjDHnVm48BgaY27XrIbLJDBRcqMQWXm
ZHlqc7gcO/pz4N0nfMGe/0pDN0G+X/eAMH19RRyHg9mpC3RW+O5/BrIb/pHjxqGC
vIrpyg+ctK314m+oUSgJV7TpJC4a+O3OCiDjthkp54Vy2jS5SpuwEEvOBBVg1J/Z
CtBDmbQQPE1IUcMjd3/f+Q1nf6ElVfRryWNqik0pmcGRJc9n8Si6onzE3hH3bFlU
ioy7nzP+LdiT7xaX0bk9YzVOOj3uhL4g4GYZOBthtTD38XBgx21YpJvAre1WyNDY
y+CbFjoedizgmiVeN5/mq7YiCQXXqk0xX2xd1qEw6SCn0cznvDm1I68tXWAupn5t
WDeUZT9M/cSDAtJ6+jA9MWWinlkyb0YCY3bmcQXJRBsFDuZBQrlRjCaphja4Hfjo
wUwjuCM5vC87YISV3jH/Zxbon6fLpIlMZsiOv5cR8F7GwqYNGl9kN2GHrK2K/hMS
j9MQ+H7m+m95uf7RHT9WQTXULv530BQDylr8deXU2HPzqiYosKRd7Ycv6PhLmfXp
dK1ujUBVgHQ386XMGr5fN5dQnLlKl4++VURpRca0r4QTq3DMMRKAnQsJnBL9OUVL
+s64rgeXVtcAOVGlK3Ss+eaKDt1HAktCtBVe8KSK8YxddRMkEWm+7zeXsmvTnGr2
XkruOuhUsHwU4ds0NqqTQDPGFTfO5MuGUMbSfwbdrGM9/6LPzsUfpZhpTEyfU2GT
ba415IwQR8HBe5W86aCA2kLclkhrMUZDlKoRh+b1VbWxkuIdsz2BgJgtfom84kTU
13O++3nl83VK6z7GZ+fgShiuBbyc2A2FimxwxrHpYDwHQYDbkL0Ykap1LF/8YmhU
Ojn49TAO5zbs3kgRaWYiXOA9nsNaUXCOOXaP4MKa2G4po68MeAfHPC3yZPmDjUbu
zXVmWsKTWHAoQ9cqzXN29zZNb2sQQhKAvr/VgD/am/Mjz3olCVzQh2zzKQe1Aj78
w0YEtSS5wpnXCnyWDQteGjLvZemrPfDArv1ZioH2XxEAPzPeR35K/zF6Mhvb1mnc
iGjIu3GPxBLju2thzYyNy9mbWpF6/AJRcqdb0lL3QzOsGM4CiZalz7hhkxjTWcYs
mU5yIjXIoYvkwFHIloTfv2g9FyEn76rR6/MoJvY4FvoWh1xTtLlh/wfr4z8mxF2b
aS+BcvEiTPUYQwYZbQe/BiLC3dyv8i8lkaVmpGwrwStiE+Th7tQcXOhNAunESc2A
7jzoQ+TDFOX6b4Bk03CE6Q/vY182BK/qj+03JO1+8jaZY8C68CkCSJCtt1iiz6n9
NhPG8xVdYnrzCS8x0+wTXFPswsbfp4Ee4AD1Z/93aCLiqH7m5pXf0I598ROSYzZT
SN+KT363keKoDhmjXSt7CEHqdBWID/K5l9VPWe0uYCGHYLAgVhPTvh0aTs0O4jHQ
OIWf/aSR/LmRcg74MM61eV2uT9dWmN1OQNGQD3yzn8xeZRTetF8UQOWo/nm4UT85
fiYNlFScVn23++W8TZbjdEdKj0wbwyqfrQC+1wjTU4DKGwnOEfG51G4HQLh80S5X
7xKUbHy1SEh7D/aiOybuTtaG4YFRQ5hbfLwsLp8vsmpWdNmShHHwmanuXEBuXles
t4eKl0mEfp+cH+Dmpv5Qya37r1JM3FwIOCtPovjj5RwKID5c2PJlHN+Y43FUgTwP
S8T/SWk2t7BmUvKzurx8YHrvhplzk+7QLvMTfpHsVx0FWejLREX+5qdnWWCiRWB0
zjtzMJnS7ToE8T/PP0NP+Xy3ZTfRg5EydBh0vgxvwpvHXpRfbwcaH19UODMHxFY8
3VAi1DG/AikTFrv2y9iJxlSFfh78AC+W0DlGSpogZLNjR6FpZSCOYFR4toUEKYvK
Xy9EQaWdkZfzqxoo+6HBg+reHpNVlRyDoa8bqRlB/mXYj9Sc6x2u6t3wFX1XF9Vh
F/nJT3BekRQzH23NKlFRyxcBMJgr+Mmmnl/twqPcujXxV99Oxl5MKJwLG0AXWLhl
oyGNlLra/lgXE5UyERcHZrnTHM30ql2kzMG3ceiYDq8l9ubFzxVQ0jCqsHtlzxER
2l41Zjm1ScBjIfCvv9sFQVBDw0ZQ3cgjNgU2lPkALrZkkgQE2H8nuPEDVXqdxCGK
bMqGjFMas7Q6MJhCAPlcOX4Ml8KTgQiJFE+gPzhlKmOpdg/NbEuBEwFcItFT22vo
r5ithI5vsybsZYfI56S3K7EaPfOvpdL6Iqt9OE6HDF4EKVSRljS5iGr9iLMXMIMy
tYhQef15IvsubJ6bOjqhfuGdJ8/aZ6GQ9SawEmDBvlUjsjVCtI/1h6t1KBib9d49
TAsWY38eFIJQ7p+zlJuHTLluJUoKidkQ6YAEhGDnYwdm/mqJgOACQrnzjhTzjhDs
BV+PALMcOFCMZRyFjaFNPUJu3jCOA4pepFMu/4ONpMLX24O2crfejCNbvx6hWYAy
Ixma1arxzkTFibu3OAskR7h5M2W2XgmRoa1Q2Ie90xVqo/3LHmOKQXOE31eZ/Bti
cXqguRY8GPj/aEdSe+eFJRrwA4+r9xdlHIHoXHfGjOCDzG+VN8pIgOcVrKvEZ5L/
TkxasXiAQIPj2wWgtqURNvnF+fDQ9hy7oZ1YkXBuB4Kk+RpFWZzt1pb04oXyIJFB
QmA1IK7HrasJtxecgw1LUd0w7maNeUGVG6eaNZ3EKRnIp6HmURs89rctG3udFTHw
zBeqDFb3Tj6IpH88B73GvNorkF2PRwi2bhQRZVLQu8dfAg6x/KktJXqS8+Kt7oIB
eJlMz4YFzoxYr902OxJ+IE/3BfR9Cj7FE/6hv0UFrtUIdDedyFFF85pqINXBsT7B
0cqY3TOEIi6FYPdbDm9jzh9qNVhxNMkESQ0l2clpy5b/qwigRtAbqwpJdb6As7bZ
cXiw61jQRtqxQF6KNkWqgtf8qLB1zbXjV8gMQMQSu+EDo/sHABFx22In/R/uVpdl
0D0boJ+kZS/mUlrBgBdrV99egUy81gDasr0e2gtdlXn41z9/NxEYHxm4zA3NR30m
aePuxFtQCe/7J5GncXE253YzQxQxhD3SYpq/xI9UB5JSG6cs0/RCcLqPzSZtC4Qy
bEqvS0VPIiCjg136KJ/Ai5jE0OcocoXg0e8EbJPSYObKps2NIJt93W8ZsEektXJE
2QxswuPTBOjkA0fqadDKmS9MytU5Syc0cBg03pB5cMscxlvviv7H8SKFJMzcmV91
ZJSmbxBKsljYvfLOmYnMeZMURTPSZjbh6UjMxj9Oag5xX1lLN9i9NGJ6M8dy6v3l
DcjWQtR6H+YIlzSkZEHUwwdAazJkb7kw5oSCCX1V542SrnkQAeu/o0AMLlA741HR
LiyNCQCAeeLXAbCN++Ovom4SyAa5OAS5ZRJkUAa9+rxowOhKRji7uhgUS8d5ZBmG
0z4q+xkiEvHB5NkYSxMcKznHtVWFNsim2u15AssJuGdPCSHBcaofrU2F1rVBQmkf
JETVfY8FnDsQmxVR4oQJpmN85QKJWETSR9F9wu/+nfjBnIFcR6lxIpB2/6R9L6m8
AzQS7V/irX7NB5Yb9dHQFhU2bke0dtE19k+vOodL534GFkWAVsxDBCXuRvNQm9AU
m5rpMeoLJTGFrtf+vLjFqBPQ5jsjz+0EXpfxTkOQaylzSQ18Ey0fmM4RBden2jzL
pMivGPJUxuJ9Ix+lM5cpDxMV7ueweX5CjlF/aVGVucuuU03KQd18wxZAKRh1FxW+
M5o5jkMWzJSLsIRoms2QKWGAe9Aa/nqxNL5MJGHm3OuECfPqwvCgICMUdTk1X+W7
WcPSHzOHjupjVrpMeES1z15cNG9CFs+00Kcl5LcBXx9J/5e1ksL7+l8PV1D7JprI
668vzL2UgwTTHTOJrQSNuBINIk/HFA6CJED65thXoMHoWjb54zu3dEDlBowSv0uo
F6XVHjeXsdGNIyu8ioAIlA3QOMa2KnTTLUQsN3leTLSzcuWl9SwOVC9ouby+4ad5
N/nXtpcQohv6gt473+kAENzvRPG/cAA/dTst1u/+7q2oxAIFNrkxTUU/V0eGzJ+5
HbiPqt/HmXg5Cn24etaiEc8QbfpG2Z4coGtaNB63a6lnDSSG19nlv3CuOK9rah7s
sMDT6CLl5iQuaXumWKq4S55imE/Q6azaycc8RMkLGzhgxokOJ1HLLU8OUEGFWpXT
Fa63djYgb3kr3RnELC21ACT/e4xnxcs8fCoR7nBClRcFfAY6JLcszRPEkqLVY4h4
0CNlSBANP4Bae3hPXgDNxSF48nu7/U+r484PEKiYc5Zt4w79OvKJWuMoIaol9vz7
GzWpFjuUM1yCPfEYDXDV4rpsfBjDS9fidIdcwSAgzCFQVrEWCUUzGPgprKst7h1G
der2ZtdXklGRMRTDFKtQdNnzefYL2X+kiE/RXLIHaCAa1Uw3tUQjpFr9a/zR/5/o
27KRJ2UKKE79RA0KeyrNQVGw7SKyziH7LDWijSkk3aJffLSjJR7cY8CGrx4RCRqa
YpklsEnOwOf03dIIFavNIpbvEUJQoiOc+VWzGGfGBK6HNT6d7IEs3VRY2LHtwst8
TtdnLppZmMJq0O75Wy/pjTKptFMnUL0PWTmS8QbOG6PbbfSp6DpfX3M1pZ+A+VxK
IY9MVr7rKw24BJE60WHciPBqnc+x6cM6oNqhHtfId6/5NCifJFIYtBVcHrY7hqiw
htUNYgZUiwYaDxL48GoHY48G76vi2Xhn5q4lArhDvlRKByxd9ZsAOLSrFRTnni6H
WotHS7PZX4w+4hRX9uVEu4mw5Kb0DUR7tT4NTOldZVdy8Pf8UxHmqKbg/SQGEBfo
ataVyNP9365PLSrWO0aKu71OBtB/G43C7KCAHcLOfqQPQ5iAifIH53fwmMG0oU5i
MzpjExhyCNUMOl5Z5ATKweKtAAM2u51rAtsGlKS7UyWSPjyzydlotZTCNHHb3GT1
mQl6hZLFm9VISU/yftKQvbWzwPUvGAn45Zjlac3/mNWCnRfJBnWNtmKUdCuUSCEm
Inx3n4cIeQ4WUbjqpWZqdLuMJlBiSJ+GfxRhKH6moCsCCqeg1OlOeGzJbU1DY9KO
x0hrzVxftZAJN/6XcMFMjAmy9VHdxcd9T522zgaDQsyx6ssExd/N2EK7T63rOkrT
KltogfVpbOPR7CjCcuqDy89MgbtdnO2Ac86kZGAfLTZWDYYdvfT6LkhomUgO4RVX
9DfUFJV0ck6ls/lGhHoHEEGT0SGGBah0OkNWdmLVHcNn+87qCjO+JF8bL0e166cT
rIoCV9AwlLaRygzFptV3/L6hB6Q8MfMxIuH6JiiOAu6Ua7mizA/pkZLfM2dAxHzc
9fEepEmEXuuiKsSWsJQxjWK8EUfHD8e3WZbxcmX6JJWTRMRzh6B+UwGUt/Jkr8jR
POyCC4j5/1WGF7rqyal7lOyk5ahOEoyFW9M27d+vNAqH2lhx/7JyMIT+qQs9iz8S
1xbXFKxaxtEYsWc78rUq0B/BI4nJYns3+VS/LzEQDM3kivInLQS+Bo9D+j7mWCii
pYnxrSMF3l4TQ4qDkwOvlxSMYY9N8mr0KYuniDTRk7+lPIuxP2jwkCKHoShUe0nr
IJmIrfOK+uj6Z/etqKzeYOkR4m0YtXgX0QTQHVfqKSEz/FyjFkF1L180q9uZ0P5j
rjmLkxM4a3/qR/RXGg/cq6NTzvSh1gY6KLKlzlQUujDG1HScOPM1Xxwb6VXaGWbg
zjaOJDAjZVC/rkABK62PYoKL8b64AZQorWJJKpBF162PfGiDIFoomSZ1bZbVU5rF
sQPivov4bPTHO9Tk5wAqq8EeNVom+11YQqoVABxGWv6jLzoFnA22D4jjGyNzMg+t
xzV7t0OO7cHhhIFmdf2Gm1fQpPy9UCccQNmZ08K/qxmXEUIJNiS0VXrMQrSIi3hV
Q0os9at+Pvp0nNh8CLwIiHCcpC4sOz4kP6VlE/A0/+49Df3IXh0fwYBpnD3ZK1lF
jqFs/l8sjjC335cWHdWMpPQIoocRPFwo3xL6n/aQadavjtsF5TKOFTLnMgc+hAwi
JRWIf5pqxkOUZRm7saHx+V+TPJXVH43SGUXrom8KcucFuAaYLyT0qbfWYwEaYtqn
gFrsJY2xmdoAvmR8osoJBX7UM+phvEbug6jQo8CtWSjIuUrhSVqa5A3NUdadL3tU
JcUh8NJ1M/gIWhtIpysHa6wNsLTUrzqY0q8UxVDf6k1br1amMHqlbMhzuXryxaui
qYWHJmEbIupPtFQBoy7GPrlTlDtKhCz8PlicoMptjErkce+EYobx+XavcBcamhkg
iGpQQR8KnMZ3HT0cfxYAJtFcXWRGa+cNUsJpiXH9tnuQ5EoNzyWf+Nxl8fZus5iB
a44GxMgn2bMLs2vGBiNCvEpALvtc/IvNp1yLAPaszm+eHbfnnqNQA7OpAvPsvggN
t/n84U8BcHDFt84dimwdE1BsBZaeOnNlPX82qcV8V04glog+EQvZx20jr+z2amSL
4I5fEJkGSjolTJW80Mryx/dMvjzENp2EnqkvNb4g54kDJiO4vMNe154T5FKgwOv7
Q2yf7gsZRVZP3knFa0Btmu2S6cG+bjZbpOrLJbSk8Y2Pl1QnE6qtu8ThQ02QFexc
4JBSgtikLfgRjABkNZJE1ug1qgfvLTaEUD1tElPDHQ7X9vJkddKyBXjcoQq2cElT
feQJ7LT9cRchjyJUj3N2visiKfkOclfRm42O4vuKgBoEIR679toY1zDSTUjjyjsr
MVYad0+mfXK7CKvIcboC6sNfFTNSHvaNS6sQH2DVnlnXieMvy+xpMv0bSGYDK/mB
9icKfmQ0aWkp1m721wxYXXnRzdh/311eFsD7VEa2sIIK2q1oeUn2n14JKPlZp/gM
25f3UKCK7eox8oiPskMSNNsVGFiEJWZpkWgQ+c3u/68IwVqTVu2Vh9DKlbviGMOY
CJqQc7aw6jDaAVObpCVX/mNOFacpWsWRRQy2MGr/bP2NRbJEPMXGueg4qJWVCDd6
AJoOMZ5Db4nrKErkOWwv/u56Wa6bWcEx7HwNcaqbS8rcI+TgP/JoSpjnwWP4/jDO
GsYVQf8Y/ocdiq46eghLi+pAP+nBp23cXTW8C1v2nlRGzKMGuGQZ8eO8mgKyAiy6
rr2WLivYq8u2+vAZQPUe47cqE3qD+UD4pVH60sJUP1ZJGv8vOGh1STgFmm3o/U3A
BTYktTkp3lshG0B8k+/2yz3TnldAqWsWMfAay8ijsprIlx6QaBsj6fgz5gKzmuDV
q3FNY7904VK0/bhYDLd9vsJmim42ai68dskCIbADbdvTI7CATp0JnU57sGVBjNC4
suL4qGP2omVEIU97VrubkPim8sHam0l+8McgVE2jeG8b9QgDu17nbwRlRmMcbmMj
nzQeG3o9m3K44pAaODzpPhkwKHpVVV8cKkWvipT3qJhNOhYmx5W/2RhV5+EWoxP0
o8Cr4J3Eb7uaeX5VQgc+sMmdD9KWK0lDgDmw2zGl0lIzsk6sKF7xPKax8cn7yyOO
h7R1SegPdF0p/iIs4bTVQvKHMbDkgjbOo71bTz/67fCGetOuF6xSOGjkNDaVkpV4
yNV4JMCaBfJeGGOtz+ezntB5HdYb5autiNslf2STIfLKaOq6fJGhjBGyd5yv88WI
tuNIkkVVuhIEIlHPG1xHDbLoLctCzCH4behi+EGhqF0k90EV8E2uMhMZ7Qi2WBAr
PaEoXuIbO2mg40Gf1qLisxl1Lb+5Ip6py8KAJgj9PMHvP+ThrFivElFp8NUfHawy
Ii6qVRKlDAXmoKjFfE+63zfNuyspwt3bVEtjgGNlChOyQcG9YvSp+bR98IJ1Te+V
GmTi1ToO31QeS1c1/o6FF4iDrkrj6iwpqKhw+c/5XmkqxI5wloGh+xcJWrIZ8F9f
TA0B/keqMVlcsxG5yVKGdIWY94J2o8+GHbZ6EqyIt+FMMM7fMEH4tNe+QBm4Ol2H
QqKbU3nfoZmxj+ReqmFjVpEmSxFaKtnWe9F4SC7MaR2G0Tz2WCF+ilM98wONQ/TE
JimuUSPDle3MUqL96AuUv97D6Cdwwv3rD5NSHI9iRVB5StvAc0N+D2blD+phkMDg
7kgLFVoLCUxjk3tmII36E/1TEh6ygrYmJdMQbIaaY5UMnxCnF6hWwujMovFT2FM3
2lJRHsvm8I0/e+Rsi20T8Z3oKOpb0ziMjPJeww2ASVgPkZqLmQIwUp9g0D/FMLWJ
fuFbWVdcC4e2VeQxArrYXl/RmX9lEirnr+KdU+QC63nEWT/D5ld9LnrH5XA3j+p+
IA5Uo4EklxSi0Zmyc9xVEg2o2BSFk+1RcDpTfMfwSq162XOXSFc96zUbgAD1B7IC
pjBS1g2rNkVzHB5TLpTWa+71AyHnPV/onCHGkowJPpA4sBucUhpRQi1R29UzsJyS
RMYCH/tQwE2ZOxNqoTG2gGLn86A0GxP3JbzTbt9VUHuMVR52azwJlTAPtu8RcPlA
E+SwEvzMHmhZ2LSLdX9GVN9Xo/HS2iOGMFHnviKf3JvsJJc2qMUqKo50Gix4Psz9
WjRAA1Jr97yR68JPYehD0gdAc16MZK+2P5wXdQ65NDFX9ZJBoOY9KDMg6ecCQjRV
QzsCrF7UphHmqwlp+Ja7Nss0bb3cD+xt0gR0enEHSnvEw/EeL4K8gXGjHE50prrl
f65QmyAsSTvzV2qIiwyHSHpttRE9Xw3hgSUir30cxrTk53M4FonMCaGeUq60JSfL
surUpT50ehJ/yyEq9AumcwiOBtXEnJ0fZ0Z7TX6Q8EfU9Vr/Ztfm0NdC8WFNNWpd
S9UQTrUYlyRnQ+B/0p/TsGED4YAUcq3D2VAh1ZD7kdVpeimmjOXkk38/v5OXqRir
GqdVTYangTxkIoPVLTpNrIvjK3tSVpS/EE3DEug1uBWVn4umNFZhbOl4KWz4gyWt
g4X/CT/VMH2ngxab1oIstoI66dO9R7PSgQvLSAEZT9sIfQaTXRsdLuc3C9ar5NHx
cfEP8ma6EOvGyYYq1gmNkm5V02kQgr6VNLqXFsf2GxDWSesli8BC/SjbOMgQKeKJ
0NzaPEFZKBBsKCPqDENMoBcaPHpFqU6BNAlrAGoIPnuZSuE0ijNomWN84qffvDnX
60iN6sxb7JpmeUV4FmzbqBfz/W0pkXYMpBTubOPSisj0gT/mNqW0Na7bJW4VHweG
8iNAF7IX2eo0DAjfUAA9jjxzgmW7E37U4PHcoMyIZQy1RxXx31I+aM1+NoiSTxrD
Fc2GOsEBA+J0Nk/uMlHvNlpBXBdA+IAGkI2xPaYg1QNRfbsMPgAg8xLTZiZqfUSZ
soc6jax9s90FnBERrYp7cb+EXEyiX1CalXAUMz8WUkn9tkNSSSYbmqFBwLIxgiz6
BZkyKSzLdUDv50xDgRlI7mjm3WfZiJnXSQrdzVweBNd/0A8A+ZG8iLxj9qOs7WLu
yN4qoPmkbAkuK3VtkLfAuYCxHq0TKmamCxp+A9kedpaQ0IMCdyBDJ5PTbnWxMpTz
8kz8C96cGH3nDUd2Lk172ABfmWUxFqqLL+zNQzr5jan9gAwiWijfiTDVSc82yvL3
s9ePSFSrxQVftKxiGnf5z3JXF7S3UOnkUZgDz75FEZuKg3FQg5Lhf4MYRMx5rm+z
e58bKMCfxaCAi/T7ryahyZGhOe2gGi2fr/UCG37xJeSo3bEGSlKgY1Vs95ddv3QK
1Zqod37Bqq0398YnoS+hOF1P3nC5vvMdEXHK/3vZc4InZBguoYJm/IZEVcVljEOD
xw3MYhfN3zNyjD4x8UZaOWmjYhOQ83lUgzvD2aysD6q3hxgSk0LbSCjc4L3xKnpW
R4opkkDHNbsmWLubp2G612sNWo5jKiTZn0vzIsA7PbGg4TCBT6Eph8QObmTPpRRS
fKlKTRTVly0ikX3/u/waPPzVpEMZVRt7LYDtB5KOhpbxBKFKA9KlstRYt2Kj5XvV
pdnwUT3OiS3r7m9cM+H4CeVYvQ58ogqDXxFTV1YLjqJTZ4hSHEnxSfspKUqWxeUf
1kG8IerU8HO1DLunz4bHYmyshbXJ21pBKL3mUEls1N0wPeMor0fo3LZQlj+FrWad
/bWaeB5XFGZuZP04l44puznXduPtsiVTWjiG2T5ARKT4DUys6B1yK2Qj0l4/e9SP
8Gn5D21CO/2QL9rM7j+BjRjmP6VzI1u0CTXlNERK7hD34FGF8u31Wp9/pfn1N4mp
GkKFQat9CxmWSkOkeXcD61kzB93euBVRAQvoQ31+rTemTj3zyr8Zmx3ZlhxL5YVz
x8BjsXHP8BlJ2N+QclnWWNWDPEd2gCKZUm7ktVBOe+JehO7KfFbfmedNJzC2XdTE
NJ8OR90torxP3A6lnGzvbszYZ49bFxTopBSWjFWuAsnpDWR/pbpsZG9z6BExtW0/
BYUh71IEFKtUadZkK1N7sDz6n89sgqt6eSs2O7bbbnbEXEt5JkASm/dS/mfAGgu8
0WcDZ7EVEjjOozN0ZIi/HgfXngY5dsDruShRc1Z1pBD7A2op4CHMCVCKD9sufCF+
gA7NZgfzgCga71ZszYJcxRXI5C9npwpOTzS5Xwv7GZGptp5rNpJVnRuCZlw0scdE
jvt2gsspeMWln4ymjy7eifbUrPs8h+lxkN8F5sjYqB6RyDWOGz61iZRVwkuvuIm5
mkI5++2+MLCu5X2oNCURcXF6rYiaq6Fgh1QQgAD8m4Ie54mrjYadTlRpSSCd2v2a
7BRQkQalApUuBuhVMbFZUoU4fp7J9cFKVRRFuTK5C8CngxJ9oDLiZG5LkrgAt2mh
T7X7gOaNIKMf0dyxEoX5I8JdSJ+EcqrCHTP93YGBrBo7rzm0ce9QSKzzhQ3vGDpB
pzWHh2xbWuYQJM7EP2IbEszX31oBj+K2g016UP2s4h2LyJmABKJl9n8gNbCC/cyg
mC5UOu8xu6hGaivuPvYTiSCmr/Pi4TfyT5TznscVyklsZXT8KHoa+hzu29syOiNL
a7+YdsHvwnrAfo4DS9avkOtoyI+dHs0iIfgkNUj97iJ8IqfxdMHEKJcJ2pRzrd6K
pZtwk6ub0ApGlt2Gq5+06wvQrEAYUatnDfDQqfEF/KaKyM0NCvHeO3E4o0gdgQ6M
8364JSHCxIEY2MBxcR1YqiqPGVEo5fNA7Q63bUDd5UhVP5G42eivdGT8eRhf8iRs
tXjbTo7dOfIh/1fkdIXHniWCAFxF/t/tuVSIVs2/hQwJ1/QQk+v03sMRp71dj8wL
Slgku11bjOn6gHsbbaF69QUxwnOjbd/zw+TDeMdwafIy+4hLaIVs1WECJTb8Xhgd
EsFs8IoJagCX+XZoKO8MZ1/Xln4KZ7qNiyjUjfI2/UTca0wcx9w1FGPZvDtLo2av
yAlG3ICs4tgpwxtDqcRGDHn6oiVZjnxnFDre9AxBClELmNvUnM7jFGhMn4oRbgod
yMr8k8/LO62ZXFea0J3Il/+r36m6XEg68PFtiCFdDS6VCs0SyIQhXap0juxNlj0h
PDeI8RBwSApG0wK/ExlWALUAGs53ndam5Cx17npNWsAGxiMrK05fXtW3JfrIZSYn
BsTWXl5gFUngjxgynOnuYOcZn2h5ST7AeBmpS5J2g5Nagrtnnn8WXtFKNRM/SJWK
pO4VrnRX3W6z3qnuh+61/a25p3jlzjd7uVCTRJ+JNJrg9X4+nTAve5R3Mg6ciI6i
UG5YVuvMDyN8qc0100fTSjykQ4cFsjIQcSY2UYUPg4aFf6SCSaQ+sVXf4FSLpY+N
VFaNxajNrjN6RQRB2x4dlxXu8mh6ctudgE7hCQFcuqn6n9ziQP/biCeX0JpLvfOb
wil3uL9pbkpVdUkulFkpDhqiBuenNlowCLJGMc9o9epkYjR105esfqxW0ZZL+8Fp
8z0atHF17MzzAl/zR2vWIGnudVZZOqatx0hYCFH/nipl/GLAgfnQYOe3EMsV+Vy0
hds6xG132tUd5vHal5sNjckAgvXJe5Wh5s5a5Crg5IaIF84GeoRIhmt76m09KYDp
dgc32P391txCS3R+/w4+usYiVDP3L7HtCIdBjndEsDsgOMPhgwH5uye7agrYJfiJ
s5KAUR6Z7/dHed2f8LwlN9BCWw6+I8BzSnmnenLD1SAPDuIJKgxBoUu3BbIqqzfO
Wy2rC0thRM5fUyD4MMmFwZTXBelBHVeSKaXyCWsf/aS6POGu1rb0iqQrax2v9rET
nLAr0DVw49V4WQ8E6D4wuDkxwJBZoUp+ML2DICUMWToiII8SY5ML141OoyJY/gxi
yveU4SOQkQqN+K+tNRLLsyzmkrpILFOZPNfVKz9xI37cqeE50woUabCR906GA1PJ
iXkhK8y2qKHkcVSmAs06ug63vOTBnWOSZKj+QVvQCQPLgNHK5xBEBj+/SiqP4AzE
xFK2nnC2EhBV7NKKCqsJwLVYP3C0DEIP9zXCg9DxoTICSpLw0ujPDd6KuELPQUPP
U/wBElqt8PImuHhmE5OR5S2Zu5d4rzcBDqXbJS+l69Gu4LmObGlMNnY3o+CDcSvf
kc6l5IU9J28q8UgwnVWhEM9KyF4idhCrNwXyeXI5kQcBWNmesEeAhkqrZaz9NanV
Vrth+sOqrwMEtjkZmM06oVywzPLs0q+90Y2kZlpDcPvD+DfIBecfCrW194s1gTrJ
zj5ARxOaUPO9sbzPLBaAcyoX7KZ9O4LbCgSWaUrsRcSNTFc6Ubj2czrsp+1MCdGj
B0KmUWE3LiuTQhWocApAAe0VnesWqCoVO6i22Snogf0Qjao63AFrQ/EC059lp9w2
Qbp5NNyQLwl6SveRZjALTcyFi3sv4jpZRGYuw4Yp+/ju6zxXILUbbZ+4vMHVzpTm
H8uKViJfX36l/guLiBAa0yVUCw/6hsFMep7FFxVYsIoppIXR+PCqdrTbxhgatWZ+
SCw4BOWyJOxQcVnoiGaw0AfrlBn7z2PgqW64u8qQPznPowFdqXdcatLssfjIOrb/
XnNvPItLKVfWgdGZXSD/KahWCqvvHEt7R85lIYT3PYI/p82gTV9N7o6J2NzjSOgJ
Uo+Y8mIUvXD6ZCWmHTJglnVzXMcRl6yOwX0QpGICuv+Y/D2/q4kXns9KuBlNogbd
kq7hIAwlTnOngbZFDlKIAFhAuUWd58Kq7eWob7KhdmW85GNVpgwMSR4ik+A6mXBu
IWO/+64h/iQvw+Y1k479hE03MNXFKYd/9I8n6Oao0WLWv2h/NPWPPnW1AVZzMIPu
GMMSlfDdsl/kZuTqCO31WWTUV6ycBaDs4JxO9xVHzhwRJv4wy2MX0q1SaF1MZoA/
lcm9bxa4IPImBi2y85LVX8bxj31Z74Es2MFRwIoxNY+XMQ/du+yPbESKbFTm4dsX
DbdyxtiNsQLqGjVt5NWthf2rU2FtaOo/o9PjyuXHKJ6JbmEKLWK9nGPrWJOiFC0i
JaQAXAWSOhrjeURLptGma/c2avoKMszNe3Ent7tpbzz4y6G8o79J5nfJ6o0JFUoS
m4QHN4fx9+IDeWHOe0FhgEUhs9QXSRRqmD8cn38RbJboVG3oHomhxW8grPKeYVoG
Usqsr3KrVFdhqLyrr63SERmRnEysWjs3u5AE64ofNYNL2k94dVykYkaAGcJdN8Ld
fdvC8HGy7hTzVu0mckAdVZ2fjrfQUYCAJ8iS6ddDLXHyWSqex0VR+CdKXvRkxLeE
JVxnCnpl4/IXRCK+g8Jx2oSbTfdlWAvuBkFzpyZzrRyzbol0m3kEYYxu6wDtQFi4
FdLgMVQ0rpF6giBukbTU8X7O3REzjGTE/C8kM2WrY2H8QLEqLmcu0e4Jj9FUnTUd
8Yz4iwagMX0sn5D049Kk8N82m9wt4ZO3z926FCUpaJYqgZIeMk0t+YJM/CvcyPy8
kx7vvgytMSH4uujUpYJKcIqaybYW4gGd0lcNSpx1tHc48yVz2uwkyd1uuIduNHQa
Ut+o0/Ol2BVoR+6gMBjKvD6HV2RzBXAwyyEaKuh43HcV7/LMtiiO8BTK1pjaJloF
PRQAm1S5UjkWvMGSD0s6mNr3mol5UNcuOAs8cynwhLjlzlf6f778s3Nn2hOtuZqG
TH1lv9Dy2RgC1IpMW00PXVTriQJ4g7dta61RKdxhlcY/IWIFo93CeW+QTXcvM3SM
AU0MMOwfGFRY6K2POQUC765Hq0RvZ8rz0vUZQ8lKB0qrFcUm9B5GBtTdYFUR+V+A
KsLQHBVG+VwXCjCpBGGndDgBKkY9SMtYl6iathyrgPh+eSNwjvRtQjsrsGaJ9p1p
kawQ9FyZmzeCyRl9Cl1934IuXtZJWUBqp7Lrl+y+XDGBFitnEGJyHw5MFPC8bV/i
ycKgzwsAMhuyBeUvBise+yaAFPiMqtiIoSIzDakTHBpDfInce+lAMQ0p/7C1Gxyj
fQ6RiKynAcj88yGfSVXZ0a8v97QWngxwqR2ThfdpUKML3oJ5AvOZhj1oatHu83/C
Jeme15d31uklKMdS7/w1AJzmqxL8OsgcYs/PViJqZePydL03j2typwS/0hA3X4Jf
Tx/rcm2RtGDzpeQlleikpH0I+SlX5UucuFIP9zOQEE1LC1JWOnpXFzfTpXIJgJPB
yBXaU/mx3I6oxS5H1LkLFcIRFANj5xunKNaXK/fBuRHayMTG0EHKYWZJYaONjbY3
kVPFPi6RSZYjW4Q7BW6c3RJvJAKhItt8wE1W+R8FDTW2Ll/5HBM3x4c9nGWjPx9F
wLr7Skl4J653/vX5oT+5s6JoCpf+rkpeUsBJmARQCKi1LH8DIYTOmru9vd54c1o9
trpSSoWwZdAu6t2rtsKwY5XJMLDKS+VawGdzVbkOvE1o16VgkDWR38Gw2afROfVe
oucWPkZWTB7eHLDTUXcC8tWTqWEpzXMEiIRHnexrBTCaMGKDdtWWYMWLPVjskL+1
otuXDQLPyaFJwJ8fVDc8piCbsmCVEbr2RCGJ2burZVZPSmmvA+mf1T4Srdyu5RJW
7ZjJq0Ha5yh648hOjt1s+lOLdjljv6abLuU6ooKN65bJLGrXSWLu4BhZgnouDrfh
xHJz1q7kWn56xetqI4Ogaj1PGNue1SlCgEgQ1bWI7b3kLpn7RsspvN+uI+FxolSb
CfbTcDvQLebJPaeeXQrwLxh56bGRywk/2fG9APBv/i1twXY3xWYYFd5UnkPMhHyy
RX/uHHMe9t4ZYYiQf6u9wKVDLQ5tcGjfUO7ZRhg8TWglzmzST/wZ7W3oHUrwC/dX
DNjBXW2Y01lu2dBSwZLTWMgok6ERoZyosZ6l+0aAh15VwsrW1AiDfW4OBQhza+60
jNsJQOm+5moRxAEPHt82jYVgSOhgtaexu5O8gwZ0CC+OB5K8vVNZfzzBcF1wvfAR
Tf3l4KzbGmoOtI63B6VDjaLuCeTihJnNpeRzoaYy5D4opw1XuIqhKuJW/Ilc9jac
jx05DP+MKRStDNEnMT1+6CjbsQu5KLbaiyg92JN8CSfAHW05kXT4eKqz9wOaRUya
orQLUQ/bkucRQ6Al/U4rlfYCQ3M1UlF/z03x42VgZ+RvMmXYw+y17HKV78FY8u3y
DnYTKvMu4nuHBR5EL3o+/krUNnUFRdewtenW+C229zukxwtZjO1XWiXSE1/9Np/n
0AFNp1wIROemWVbs3qPreTr/HgKZbetjhlXn847K4yAezeDlt5kA6KV8DbNNlHlC
2NNnc4F06Yjk6uV4Wuqs55+PA41tT8SryFy1B5a+VC48vDh9TDxmvelv+u16VWPU
TPdC0eoKmR6roKF4LV5eDjvaDAXAn9bSdrTklGfRI9z15Brpq+8KVYjd/HmhYbx4
eIL/dgVwF4Fr0ABw7B8eIsmztP2W3kvs4IaBa04qYHtkpG0Md4MkJKGsgMnXs6qI
p+Z6j4H47HSEhwKi9W2M9T/700x+k+8YWq3jhfVlgJiltyHNW/cGZeOtKgaHba+q
bnMmVQRS/vtldrasvpUsNnLOrvZHl9oPvRE0lSfo1Pvj7JisuIYIZ/AkuyO9U5LT
jDMMf+RH4ikxt82dPs03uOFc3NKp4RzH8G1jOb+l6JYz2Zu1P2Ee4o8E7scqUtOD
AMZxo68YKHTyyiba1e4mGdqIk6d0QCu7K1NsHLQ4oNmoYFsLqSIc5YfR0SzCv7Na
x/OAyTc8ny+/2P61/1PHndzKgdTdOu9dFQTwjs/B6pU2sor+rz/5K8Y0FbiFh8J/
HmTNIIjI8SkGdHbAGfdzqRhARKzsaeahiBBsdPBbnWc26qqf2T9YlhVZc1WIbw9j
wRRLBouHxIFV2selCRM62Arc1BLNMC7aUTAkS/iOazMAKCU5xVAvNcHjo2OGmVPS
whHLF1mYqkvJ/qFARq0pXQRxQA746XHWVh1KmLGd3kz/GfCxBtAI7vgZJ8Nq3UiC
6VEuD1ueadrFIKnybof5Mj14NMGWOztXl32H+zQJf5/uhNSdqlDCyiTxwkgA+qBs
uf9MFbDdKnN+DXg34PF+7G+CDGsyRq/4mx3S2shxjsiO3tm2vkB0q9k9Nc20TJuj
muvcN/wx8Mx4z7hem/guTCH+PFRNVAf+kOUPFUNkmBt3sTEn+Gec38t7OQdmv3Z+
BKzbR+G7SNb/q0Q3e0OmIFr2aBJ+XKnFTUdKUXvoETghQMdzoxHuTvgcG3qSn0h0
BI7EdQpZTPDIb+vED+vKEsblVrEbZ+Ng1ai3YV9vE8GrEbRZ4ZANR/mSLbzjqtui
AEDAW0OVnkBP/6VVfcRzqmGH0VDb2+100r4KeINkrphpt0dbtaL5LGktAKJBr18i
Fs0x79G5Mq48Dm0sTTa7fXJZgnN/Ua0QBaFDht5XX4/gGJWLNaSFxC82dO2dGeNX
rtSMHPmNMAG4palPh9p7Zy32DL7Dxxv0CJzmfBsZ58DZKJPunPb5uMdsK8dh3Ro5
kqjcDZTxDpRXGa5j6S8y2hJS1KZmc4ptfh5jn7Kh+40NAsXayj2xv55A48mDtAKY
SE0hGUSUU7PbkSzF7WcueoUNz9/nN3cwwFTniZll2dqvXdw2iRkkr+GjzDTttdso
KfCILLrrzBgE9eXEqaCRirouSGrvm4cgI/dfAvEFq8eiwn5s0y39ddkx6Rp2nBDo
Pd2FbFdpFvhX5Fu8TQPD2uR/uat6zqRWfnergRDWBkXvVZxzfJZsgXWQcJgFo51p
JotvjVKtYM84ZmQ5Wtn2WcnnE+SptlIyOybY2Ujf0Eqkoj8Z4z5U6MmS6bYJLCAC
JUKGtJsv32IcBCVna93tHmBtTJ03jAjfea02jhndoSqXcnBdKvGL8A6VfyWK99DE
F4bwq3s+vYtMlfAz155h7P/Wdey27D94KVRklH8Td0odVmDjtAohGiy6Io7jnGj3
+p4+cVkh3RhD8c46FWZwraZTuz5hB+PHvydKpwGyaYbsFFxJ/bJsoyGBzpN6RA50
Q+OXc09mkV8oIJiCH4yrtJv4iWHu2s/qE5nQaqfA9gujVVsZEyTlUAHVxccwEuJa
6IDrZ3R4/F5eIG+cJDPnkhroA/Lu3vhfNuIrhxH3iQ5c/vTWY5bLt2Nq2caaE4uV
f23lRUIVOJmk+M/Ls5FIE78OUgniuQrhN4A6uPW006ZQ4EVpyLmpyYuJwG/3fCqU
BRp/+/askqV2PUTofIXRT/C+u/T6GhHjlzOmh31XFFW/QnqgfwcwsacVE6n6+7nc
fbHfZcy6R204nlvwb73+DEthikecuRz8FzTannGaKagdugjIWLCtXeovYdb/xh5R
yrmrPCQVMUWL6Yn+CbQLmABDO65QhNgwpeM6paPVzsHqvoyHcj6cjn6nF8Zp2zq6
xLpMimtEaGJ9IsaevegwN5OyLg+bCC6nLT9FBQMQBowxAqg7F1V8kAV5o6gZsZa5
8v7eNWpmeh2+XnXUThWwtK4xUA8t9K5HEG9r4EPX0Nenck8znGA6CuWkttqJzHia
qjnu6uqHqs9NE+eIPjm8aAKfzkAlAbBpv2SWe/doeyJMzfn4vDJ0NjTSiNZ+BbT0
m+BpDg2IkXHH8I7slJ+2E2pgKLrQbwDXwD2znPUDBC6UXncrA4UJSfK0iJorpoKA
PTP6qBt3NIKxDpVecGfNoBaN3CkpNr0m/tSUgkPYPmfY3aAEok6aoJ5O9Y38NOhl
MuSVPiMZxz72iWA8B2NwL1g43/595r2NZeHOTk52eLdqZfMNujP802TTH/Rcsd56
M+b24vwV5J6+npXxOlZNXkw2N+0l3aUbU8uYHglxlhfTgM17qSWX68N5DfNxGp27
chtEeO6uroIwXQSAZkPnAZ1Rm5mAuU59SSor0+pDi73au8OnWibEH/SebGIEePC9
/SxEIEgGdxExUnL/gSOY+6DrZi+Hk6ADM7QdCfe+Wd79YrYfwHFx/BxaaoFLsbIt
c1LMfIcmJR0m0C3YLe1T4fs0QoccY0oJ8IYC56oI6vQOEBHcIfjLCBfVN49rPKBK
Zf6oUutwk5rkZhp/ni9FrrivArlK6BfLFObWETiLa+Rf8bvqPBYFeTCQy6Kcslqd
StiEqaVb53xj1r8tq8OJJwKNQfMLBlYew+SL+LvfXqtxn81R0BZ/aqww1UTwJZ2t
bUj1rUfVvI/6ynTob6F2IOEqg7J6FGisvHDn0sIPBO9x6rmRE4a57zpHur4Tt0Kq
UDoUTMKv7AY5eIOXDm5AbF5AJHqxfV9U0LFdDarzZBMX0Y+q3H4ZpsZKENFH9igW
BZEy83ZFkL4wKqDaklob3dMMZ5eE7ytFk8I1DwYalrSIhscWFpHmV7dJa7x8rpgY
oz/q8z/afhauwyBcGDYnVaa51PHMu3DI1LgsQI+fqL18OmxKAYT5eFVRKa64vGsT
0A5ZI/YqKUSPB2KEyYZibCqHtG7qRvyBtTC2Ly8dEhSOhoxL8pv8qp3vJlkhiqj2
i+yJ8h5yIj9WvRAAu+abtyVSmFiqUzejV1mKnyKXBZO+Ne99q5+EcPBwBpZbAlIo
Ud9VF0xTTCid1qIOZKyETdE727MX8eWuO08lqnhlJvfOLiv9sPf3c2PmdkyHhqQX
U964JGeZKr6bepobNjXkNoSuEg8uMRG8jRIlFkfbOJB6UK7SoVhv4gYBMgklnCvN
bYT1Taqpr+m4LWHqzyyUIpyZvkORXcgXKiCxlDCupLbGmAgXq0dRw85YPjul1sEG
klTxjFBTPOapp2QxgGIuIC3WhQB0RN5mFnIXzp8myFu7MmJ17uI01Rm2nJwaR2AG
nTgIus04mnzSEuKR3oc3LWC18RMQ9DY0qVmXYjM1ift/HoeJXAEIHfWJus+bwoFv
hu0ef+x5JHnk6tq1KZy9lV1bTZywSKeO1k6yOQix7Yul8E6I0v87PjJye/6c5MCs
O+ohAGNs5YvkNX5xjTOvPwN0P83rYLktjmD0ZQKNWywuSHvYLmgc/TEqchh4BmLP
V68EwJwvsN/RShxS5cLGSLLttcfE70mV7DPPgCf1R5ILkT1braxVrA/SP5CoY+8x
nUL0kRI76X0Oc8afTGvWG2SVqNSiPkpZD7NSPL2mqBEFbxejnlrkiPLmsaivAISh
G72ImHJ/zR1TiMMiM1E0oa3siZMXmD7UEyNgUJ3AhN7SVE6919+h/ZTYNHur/iyh
0+MlFXBMZdk1HwUYwuKXI5tsMTA7dJpbgFC+tkvbDj5Z+P+5+0bbjzkzweJjt4Vz
BSei0wg1t6j30vNlrtiyNdrmDQAgRJGaHkLmLO2JJH9AjhhZBW5LjpDpwcfp94Eu
P59m15vHN1TRGr9uRSPY5wn+TQRcA3oSp+zQUZeF2io64xs4IItOywWrfwqcDZGB
nIpb7HFzim0ezmOTyRqQEAcFkSVn3kw0NSIzEdLbwYVi0gVnet9lPwleEDJXGBHq
amU5eLsWNpawJVE5CZGurJd2bZkLSvFoaw7+FF368pqvdRpt8qoAIGmeLeXhKrtf
lXWw9HlHuXSmGz79m7mRIDfHAozB8xFUe32L2GAtLIpK4BhHCS1zmmFxQvBp5mbv
gvrn2jKDBhwSWD1VHOrHZDe6yIiuw8VKTlvPebTT7QgYo0dMZSSeeMcvcPT7HBfs
2rpBK8WGOq1fmqVIlwNw+xRyECLRQRfqOkeFeUPpge7ZXtiGomxkk9ursSChYdbi
9VXDc7JZ99pomPW5LZO3HMVtXzkzoASYtKtdbn865MNNeAzvJzi3jNBZxZWL8vhA
HqWUa+J5TYqWqdo7mRDpNnT3KaxeNcYo9KSWmj+5OEJFMfJEd1k2caoXabXj1XDl
tnSJeLRkGRkp/v0aKzL4NHJb1Le1wRFfY/tpvBd3HxmyqKetQ0AMmIHCHtsD7HFg
tFYc0nqG30kVG9pAZEAGgj7/z0aAi433zKhlza+SKBq3O3i135PqJEC0D04ax7wC
RQLhc8JnFf8MVwY2x5Uc7DJz0OV5bfWehkF3J7y/svuSDOq10/FMFtRnLZqAUWFe
Wu5ZYj4Ha4J37OOcNCrzqr+D+9nW3fbz1/CDMvqRGMYU+/4gv40Y6hBRUp8uxtvc
GqUG58okgrgEfp9Vl9PoFQjR/BhIM/LwVpxWZBSSkTpU4MT3TVIdd3cX27F0cvHd
jmZBJqTkm+97bifO27QFNmeVo/mDK5ml8DlSmc/16/6P6FOKXjOotWNIQXqlJbR8
YLhdSxTxxloURKIjDXteCMa9+pXYAfOCqvq3eaEq9vZvhJ3+coO7+t/hOZHghQ5T
rX2fymrXKU8wl7WuudhmU5XJGveMHxxbNFpG2Z9P+6t9N04Ytc7qOMlim62SXb3P
4xaGBtzg2za8N3firP3QpzRz2Ng1bDj7JLxPGvfdS44Bp2WtppVzsjZm+yugm/mw
ZP1rN2AKLQTaRs9oV57x3MRh7RkY/1H+f1zkkWgpwsW5VmfeY/Bz0bU/ncaweNBK
o+kmCGPmGHlEjrvewDRHt59nQnSThANtaORiSz1ykKCedS0Rf6s+8sVF2bajpNvs
LABoxPhzXlJuS5OOnnjai/Vyo+PXtGUqELb3DIUqQJdgnPd44RqjgGDwggCMpWQa
GcZUKIjRuH+pAaiUEPfTh13zpJ2kYFWUAQ1lGah7wqsAT8nZv3VyZwhUea8cAjs4
5t0sVbl78JSId+F+YtW35NXfIB9oqBxZBj0m1H9bFDt/3xU6P2bgKkGhKAxqMtI8
by22VjtW9dZTMMUSnbzPHN94xeisxZG+C2Hvj7TeMja3B52jjyc+ivL7l5zCdm8g
Ia+84FdvyxFpqShn/NpIash1sSBQXevRUX7Ks1dPeO/vCzMJYD/pUSVn7nlC+QPd
J/BSXxXazbMw0qCl0ydyW1WtNYK9H9HeLgQgUdyw/Z/aOhoxc9DozZ65VMSnhS5D
E0XK3dvjDaMhGBzTJsFxPIrOBfugdd7whNzOY33w47sRkUVQDCUTWSu7FKRMlafj
eOYV9QRN2aTbzvGf/s+GO+RuRYLXl93ZF1k66d9kOdkRLIp4BbcQ9bVS8R126UTX
GWSDA7MbHRJRGW3yXaohQeOBCCG3RUc2gwloSUC6ikjht4WtaCKPJ9zhqKiGkcnI
mu4aVeM/kVZ8ol5Sw5OUkt3PFvd2Df6z62DFs5Bcmdzp62bgy0Juio7e038mbE2t
hdOBZAUGK9eN9XoOMh/C5cT1hM6Qgt1EdAF86hy5BTNCcx+uO7Vy6JypMu/3mc5L
twVX27gKk1D+Pkaio3ZFlyMzDfWiwP92WTedNT4Ubg5jfo84pt0FiM271gmnSmHX
eDO1jp6DbRngsB0ZcuoBJFO+HCQqf23//PBtVfJAZC3e7k3gV0mpkZOzga8M+A6i
KSV3T5QMpWRXPaVVn/adEk8UF/yqy0Ibp4jVaWhgNuaLJ0FvjDjbjebATYJ0vkxy
4va/RSYFfQzfJ+QhhVjJ4Y9Rgm2gYUlza+UdIbLWxBqHZBU1qQhaQM3KLG0G17ee
XCjoOAb/l+z+dNMj7iwAkLs1U/I5BXX+zCiTrRmwYhcZBtnab0G1rhVTfAvR6uVK
DzZv/X47jVdJqrCucw4HgcllnlFpWPR6EWB0u7DmhGFgDWvYaZUG8w3jht+0mC+l
+QaPzg3hCFZCQLfaa/QTXdi5g9aMZ1HB2FHPQl5docpLqTndHivqUatY3K11MPRm
OG9wJR4eQl7DuSE8wBAIuQkXvqh6ZFX9GIKKAtKINiPdbF071961TxSUYGM/Xwro
z49fI0UZQPMjcg0tVFiJV2eaLZH5naadrA8E2cXbmwFZLbppyJtdR9u2tdAUu56m
0BMN0sLLLq3y4j5bAhb3Pko8087pQY/yeoyzYGcHH6VJW71XKqUfepj94Dn3VkQt
qGRNLNjV9nXtTJlUBnxSTFKET6QOhtyeNbf5Kym625LbQwZwGnWfnFSV8DYGSs5O
g3ka5+NR1Bc4JUiV8qKzcHSEqdj3RsvoqykFFPpOcNXXNTIF1Td2Dd4Pd7knrS1x
zCi2E/iSi6DyANY7obbtpkQ42hb4UjjR9Fgthktli8G6cydLYExZ5TW1CqJf1W5T
WZ76xzm6ePLeV3qUdmUHLe7XiLh21IadkzeDSAuajZhlpyM4NvBJ0EFDK0ADdHbS
qwYfH+4QqrR17kp6JJADWOq2J8fGT+07YkP8ClcJ0/eRPBsYkl2jSD2QKh83Y10V
BZl66Y3CSRmtECL0np3/VI2tQCmEuTiKjRTf5/wYsHyNNKXBIIHrhUEGF1ZyG5VV
LEFR+6OWCz9dszMUqC4C0adfsTC61lmA85RTZ2g2T6RaLrlaH1037i9jTp47djOG
cuuRETdIxW91dh05nkwim5oT6gE+8TNHT4ebQjGqz+9EgWLBtrongMEX/qBbjer0
D5x6qKBWHE0nJo2PZVsXb8tXmU6cxE7NYwkVjFUCdvxjiFayu/KECnxMow7yMr7i
ermHlytldmmO/utkkhUh5gOvEt5GdPbfGYeBvXlA8nRA/sKx3zHeb1b09MnCHgAQ
+cP8G0kVFC5KbrtQB7X4V1uRvSUfQaf2DfHDIOTkE+w8BhQqgwexfSuMhLJT0kh/
r2/m5l7hjR6SEUAu8Po0oKtIybYQSVKwUlpjy2I0H+ypNoxKeAWa5bPs6nLBALE0
3g8s3yd6DDydspaKrRBzy+ouICixouq2ouxyYuQJG8ENRhdMygKDlyAVBtKIW89Y
0SOMqr2IJLieOa5+HvhKZvVd+9oYHHEJQZ/519Uczhu1sKT6MXDs7duUPnNZzPXc
IAs+Ix/3k9/A8CBufRVvHMPfK3TS1uuvM9Q0M87ZMl+SKnxsnxmoCma+7YHlclws
0jzGwFKTXRGDKAlk/BzRq0TOa2y5COdABsTnvDHFwizJ8qPOam/RU9dLeSmMAi78
AnOXbCgacuDN/Erdc926YHPpas+V82Hi7d5bDkr+qW9GRP+qQLFnGzistGmZZeLZ
KS9BFNhwj9KkC0kQSIkKhXlJzqC2KNVMtYfq+if4X/5rKxqMNqZDwQ5eJLIAeeRU
FwTsRpdLIe5o6UdBBHwHFtzEdmMXWEYSl107NifJC9KrvD0XU6kBdeI/SR6MDBjk
nAYjRqM1Q/rIZjMuqOWafBve3JslVuXFIXr47conh4eoiA5PCMaIl76nzLUKGznN
MXkca2fB3nM44DF3pGsr5mtedcdINheeEkLHIiei5b+2zAvjUUVHdeFveTFaiIph
1v8b5Uq9MmwVB4K7cpXwhxKZROc0P9GjwCeUVHKpyq74oqbNuTA2cRNAsBhMfNJj
oiquhYPOinrnTuP7QCS0vRRpNsOSbrWKT4C1Mqit1gAyynaLjCi62hhYZZxt14zE
oEkqgT43pSgXl7eABaYVvz8MsX04CfzNONIa0RmgokW2IsLYW/Av6Ht3ydpHoYdh
/f/wSdhyyb42ZmkId6Dv+wJr5hnnj9NXB0/bIQrmVSUI49JgJ8keJ1pZKfSnfI3C
r/nS/w/GpOEa8xDnW6Lo+uWhQ9zKqrs3s9cGSO4eDil7GQCAKHoJcBHF7lJnWUhB
e26SoFnXGp60Rd9tZFB6vEps5haZRwoXUoq2p97G5gNr79oQmrl/Woze3iKSpmAB
cOTNztZUWAWNkfJLb/76cyJtBjumTLk6l8hgc4/pHd6rneC1QPSz5wulS5HYKfhC
Zxt8N00tizBuG9kpbLoLZfraMFpXIgNdJoXLwg4+MX6Mu1yWTYKu06yA+edWewcj
8MBJWsx0hm+C+7WG7xK6AsYCFNp6qJiKYFCjc58/Z+68/7U0lO+Bsboqd22nmz+1
Jwmx6BL4Bc8H0J38144sFwpNnMi50fYnaJdclVYy5IWlMcJx/Jmsuwftua3UlmSK
m7iJILSgvSMPU6oq+OmykbCW/LPGLMYCmE8PKiw2bZzncbr1qfg7SZVZCAdYVzLT
0Yk7n6+3VJvg23QN6CXeMTQlpUn7XjI40nuT+RSlwiPpuSxHXYYxEkkXbyOLuxp4
v34nioDn5WacO9f9iT7b9JDrLovKOaPD/LMKi45yqktnhUejGZNVOCf/4/WQ51pi
a1Vo2kPOlA9/00Xitb4jgQODhcA1AtI3dTBXSx5RomMwluAQtAh/4l9rHiwrOrJN
AkEjREd3xPiWeqazLQKuhb8jFpoJBylAPFD1c51HI3s8oHPPlwgOuDE8VgpUbY6f
+Eo9wijsRlq+jBKgjfKaWYVhiY6KhK+E5IDnhN/TzrFODwmXb7Kv3rBQVghbZJtB
JOPYkuCZ12e5c+w+8jkZK1eQejy8Dsqdtg9IaJ/JWEOlEHeRwW88NFATbjfglAAO
bXDeEO65qKdqSDwQv5NMhOs8S7IxT/IxCAXFEEc7sRlonCQTlAOv4z+5KBVK96o8
pT/Bp7TUX604GZmy01E5Buzm6+EfkLA5ixQmv0h4KsL93Ghu4MzVs8cBnuepTJYl
zqqIPWY6Nb3YdRk1eNY97AMt9n6Tm3BEFBGRmCOm/jjSPorMEvS3Y188tdpLKRwT
AfuU37seYKHhE58ilRweZdQzF59LL5/Bz+biQ7WHW2wCFsIKlnIjnkHs4+5v0MXd
SeA3CNGlUvgOIr7uA+/NKBO98RtbJnDF4DTBMcDHPv2QzUCQ4EpW3yfGRngUGODt
PijM9FPjfR6WNxu0nl/pIcU6PA8jb9Do/PMrQjJVF/vw8WJa1tmm78XJYeitWx7W
vBJR6f5U9zwAzx2/jj/1DTzjolLqpEC5i9PhbtbXknWJpJqzyr4o9/2Dxvmg9dAx
wWmhz5sK+LFVEmdXrxqnYrAlcTEsjiZ6HgBs8lsjRSs9UJojSQp3I0XY2YgK4jW8
4TLlyIJr/ElZE7+wgcsO1SEbNwCU8kb1Flmn0KKeZ/qkWGGi6wcMeOJB+dtGh8iV
435wo55l6OgXI/AXZYY/e6KKedmYzB5LZsPxPb3aTAZrtYj8EIl+BQkpBlX2Q8FU
sNNmg4vsqAsmSz3fTlN5/HauO8mNECPWkRpyqJ2DLvBb6LrIJYaYy/7cd+AIhnmE
k0Lr2rja3J/r1WzMPWgmgKQeEUvvl5XAAypY1DpnrrZAVI8or2/kDNqe0Hbg4649
I1WoW0buK17BBYMPsO+qNJ4tpTeMpAZCnN7WaSc+xvDW0KcOnHM4yNSsuf6L+a6V
nkkCrO2opzmH2n1q4k+4KYvATezpfWY/DgXDmb/CSYY1Sk7lZiNxPo/KDrvu88ga
oiA3H0YirAIlKmNrORLAiUCwdFHklGnw837JQ/TzE97KfraF2uV6Snj4FLBzr9cZ
bPDo1CED8B2q1+1TiKcuHGcW3FmJerDFh7dLLkEbnX2mqjcQ6MWJmYDlkhWmSeQh
+TY+Ah3TCzpl+U+fC9vMefDqxDYJ5GI/cKrVF/y8vG2nEs36kLRQyxkxTDMvXqYc
aPhW0+qL7oSMRDT1Nre+PkBhEKdO+VsYJYeFBPur0sif/NmLnebfp/6FiEsv6Fsa
z87zZU7v16VOXg+gVA3Kk/LKYjLS+52TzG6dePW2j6hrUpVG3MCsjabT9eSLeBYG
U9hQ2iuW+/qBlRut71zeYKyrt1m3ioPFxVopXOOmSV0RZXkXVoOkJ8VISBPSQvRY
S0mQXU6RolMbp0elegMG2D1wE9yJYkKrjdgcb1ks0QRV217nWwSqDy7kN9hkD0A4
MvSyow4dsGdKH352ap4dpxKrijV7EzqOmY6cNOYf5/14+dkDFhFERvXGeS2ae398
zhxwgum/wNxpaxr43hU1OPV6xV1+Szmy+GUIXpkB7IymKZsVwdQvAQNcJdlrUp0X
n+N6GsIimmGm4hE1gZrh7InAF+2SaVwl/Dv2oBROkdhtKi4DOeLEbXyiLWvdkqrK
IZTcOpe4Q3sNzwrCuMzHocJjaEXmqv1LIIO5lc6lft8gyS9WVGBU8cuw7BsL/LnX
u4OPr1o9g6chk3MNgeDhWO0wJBMHmTnN/AJz8Cp9n6k7YJExI/I1cMa8gzCSjNS4
cxGFwdf1gbSoNllZHyBNKPVVnlsAq8iyhVp7xY1NTgdmk9JXeydTGPZMtzAEOGBm
HJy5bn95e9+woiIki5htd1P5C4512Wib41bnprksCLpKpwiQSoykF23q2E5BRg0Y
5q+Lh41JT87X+NEip4sEgzquooLRNJ7jRyKsG9zFQcz7RhlqlFUOM/UDKLmbdXX7
PNrKIK3SwBfLOCoRxwTZWqYCkXCxpnpZROGZRQu9VcnNO+SDn/Bb2pXfMG+Ek+O8
M39MHhyuUX3I4apjwilNU8nCNMsT77gOao6af7ofdpIgnhGydRND9K0ZIDNA3bhQ
nPk5HdYU4nF0/VN44tTmM/NpPJAXv7meLsWtzpdvlVaysC3twc4Dl6Dt5hHn1ny9
0w7qleGn3Wd45q3mL44gN8srdhtUUv3uopuw/QQEmXst8pXjUcZIl92V822iYnA/
M7J3saPJl03iTgkG4S/wMAwpOSmrgTEs2VsHAs3WgFlnKMsx8lAnmAlPMnkrzKvD
p/KLHrJPMc4ge6y+WrWxzYixetP2QWyAyQ4SElRFAAGAP8pdmQjpm62Kn7xHz5WX
F7UfIvUcxrLk4mna33nf+JDHrf9LXFsm2RfgmVA3C0LCUXCco0wLKgkegdFS1dcw
cjrtOlNQbPmaLIwGd/Vw5WBqipwQ4+VHekUzsZolXgwTG/2EXxzNScPmjtAGTq7m
Dc7tL77snNQsAnMLwN0ku9z00/17eMEH7BwA/ekLX2yflDderoYRgZQSY6e7iWri
G4tyVCNt1pKdUK6LGGIQ0DsisqT7FmCY/JQ3c17iu9ydaOmjqAzENBPSLV8qOfJS
FWe6sR1Gefqnhi5czhFioKGQVwhaarIIEjn0MwXJ9xUkYHKVvTYesXP7FqNJItuo
sKt5h4iraN1vS5u5DdS53JTu5L5aoSFZoJ81zE1qvZk4Y1xIB07JxOVp8mAskBok
2PJvk7awH+UwjVbqykjIKolN+MifqX6IejRnnYeVbqcLbmCylw5Gcl4gUMhFJ7yM
0ZCGF1v+8XYcVO9soafrSPtdj7f7xSXFpAHLAABkCycs4dvfbykbatdU9BxKADW8
13bbFRgtu3JGgHKwVfqALo10TVLILMhQQ7oNIiau0IeCBKzcEpAB3Pq8ymajt3u3
WoNyvyRrauvrZWcd+x4dEr3Vz2nb5ZHJ7rWLgKqzSlvKzOgQhsOJVuLr2TCQ49N7
dgZ45N+fCyRt+YZycA5c0kaWjIg4fr8hYcNqCIY/MZYOeRAkfEyvJIYLzUlL+oxy
jjxmZOqCD2kTSZpwuaebWEHDBmsbYskia4wR39TcDf+huq7jsdh4KNr9LMTmJaw5
aO9sZ/cSn7gTSqgJEp8VXY9KBR+EnpjXfgvX3Mde8zaLn4A4wD2c8AGD52K6GHnb
ZOqdYKt8ses1MCXmBzxviJZEvD4IQttwALmj1vToiVRPVfSJ5HA/ilhihLB+MD5e
+/dJz74g95jJkFID7iADGFCifJPEYnWCB9vLmuU1LP9lrbRRlaH7l+Cb4v7QwxEv
mX2XC/Aiv3vlXKxHDpAPIoPxE/r/lfVfNNldqfswtSPFyrUZFNGDdI1u8751jBbg
vVxh2qd+UJwk0A5bsYKAPy2new/r/un76jEB0rmnTzy0RgOdnkvBggNIZUba5c2M
TqsjiwYpzmo3wF2dA7iuz1HgQEZGPFxCLqdj+hAtOli17X6R62QsQevytoz171xS
DndCGCJdd1/ygoHeXgw33n3X6ZyZCJB8fSadyWbKb4+xfnoBkEtdo40NVLs7bBKO
RwuArpS9Ten9BPgCNVv0wyyMGvv6lKp5qEfGK2TQigPZX9qbzzEJR2R0CsKeoNuh
RYoFx4hXdKYx/jV/8467eeyxMrzGcBOARZP7Qj4GebYb9MtGi/cBl8SHcihKMJCo
+XwblzpNpikRrGwcoqAs+iCdseWwfqnO8Vi2ZSKRA8up4pna8aYEw+Q9WeLs69gV
eEb0LdaIzdBGzCif5z5eGAaspoYCv2BNV08pnmM7A7KL/gCQZdHAr2cgEqLzm8a8
J3eN19EsOdXXsL84a+boAJN3vqM7m3srmWU88htH3U9swGDd61DTMgS3l1yBqPDA
3v/J/fjM3hLzwBl0RaObAIOP7PtaiWHDEhk6w/J5JQG6e0yl7rJ8HndVG09GZJ5K
jjAY6Ib5VCWsDGpatzbMsevyOip71sgKJGYwFRjZTjGVtlNyPIhRv+UZBMHyVcaR
As8wSXQvOkHSV43xB3cbRW+AxSwVuCa332s5OlRQ4WJocUjvkSqiQ5UayNBrscw/
tDRiCGLUUk2J4iQm5IanT0YRKj5NLyG8dJG/43EDrmKAaOeNhsqRAIM9EdljdgXN
HqrdyJUCKOzVRXdqlWoIZ1gJhLMarYq1pyBWfcwqo+FshN9dQ+xE+bkn2kcBFsMV
ou6do4yMY3LXebVrRpbwCP14WL34MF1pygtrD2sQLvY8Xc/6r20x79nlv6qgn4P/
bhtHIeedyUlthAmHOXUUwnivwPAttydgGEUD1e7bzRQuLqL3Fmaj3PDOoxFBDvjT
dPE99cot2sIYQ6MHRIEZH4A1AbotD2uOQESGsrr53k1T4RkpETY86W0LUk/Cpy5l
FybxLDTvlDqTCHYmLIRyuTl5sVvAUammsOj8p8pF/TPJhNZDPFpVXZLecgmkY7Ri
AFx06gXZpfqtGtJvQbxyeeaPyWIQcoxmuFQ+wQr1zXIaQD7OmcTpdjq1EKdsOs42
eyietEqFRD/7dTLmvtr3yGo71j8bsnLcByFLxnJWKCqNsReLWvK6GgLIzHwL86m2
zXB/HPC/KxEoh248OU4N0Xelr906GIhjifiaDgn2FClbbdBwJFxekdYtesSCDtlt
30YKywxa/z7Gtj1KIHdsO+M1QF+XYNL4wxBmyW8y0DY1+uAuZE/rZavWnpGD+Pdl
AAN3IgIykT5ZKqs2gqjU+K8SpM6a/l1dPUiT75UnqpdtwEUKyloHlRBMt5nkcpwz
AHPu5WoXByPo1gflzJdmvdC6k9XIqUJyZxfYjAr9ec3U0HCWVALHZYejbWEsxoeX
ufHUMN7w9ZAXK32NNEwkj28dPA8IRPm/LWOh9jhL4lvgSQ9INhjc9nR8jz1DtBnT
h8rVZ4wBDkIMbezxg3JyKw0zsC/a/QBJSC99ta/duq/N+NDrwGQqMEH6Mrv955Cw
fY5LbbG9PjauIA4XEssFUop5kudZVztoJfjlacoYyT3bsLkP66xYFxAzPPlrisR9
GGEzIWZx7AQYF6bQeF9GV3i6DeW4aIVUcKPLqhNVoMDfcF2xeSnbV1kkLpYeUnyU
lHhK7jekmFXRDbBe12l+6tW0ZbClfZd2kRWebb7B8BtD0LtXFiHFKt3dC/xif4BV
iZCiT3uqZfEL/JHu/UV2ga2Tw/9OGKxCjS+a26mQQnacJI6CPjCIAzQnlHvU2xcG
4pyKGPdeyB1fHJEDBvD3OkJdE2BeCItdde/QbtbjbrrR8QoTgeUsn4NmlVSRPspT
o2bXVekrmjTwV3THSdkbJbiGzeotEkE2XatmBLd8rBj4jh1rs/hmSqoF8di64UCP
paVOrONtm7B9xyndyXE3q+RO+QLKfrqX00rMAoQm+ra5sd+enkthUdQoPom1WMhe
Sz5VkgM8FWcwrMLr0taOQC0xtIgfMufXzRMORqXaf2l52E43OzZLnEIL7K3HHpbh
j7VaJrKvMnVjEN2R8o/c8HSmmXog52ZtOfzljkTtvKye4wy19cFa/XrmkOKKH8Eo
oKUE7YsvneWDuTVzz8VI3Pjc7FiZ7fO3KiCERf7qwBPecIdHB5y7+ctgZ0AcQr0B
VvZOs2Gp4Q81ZOI48rdx6ZnVQ+/9zLG5pt0GL5G0ACgqHBTJ6Tfl1OvC5cp4NtC7
Q/1MfqQ5Ow/o6Z1MqTs3zQL3QbFwwGEkF/r/u0//hw0Tm4D9IJRsGvxdY42Y2GX3
booal5uKu46scb1y4OvX2d7f818DvAgI2EohraoK9ohgnVIYdot3ivT2mDw0Izxu
dlZLwMCJ0CPIfz5/Jcdd7lfuHAmDVMkPGNYOW8zlFkZkn6FLYN9LMA9LQt+lXSJz
fFuBcgg6tT2SvNERNiHWOB5Zp/rHrCAITpngivRoS8fKd2pazkOfk3idN0HOKiY/
j2XXY2xd0xaaLP2zjCNrmReM4m5ww2jiuppsrRgVlV7mQS5hYH+FRB6c+uHAh7cl
B6767wzuPmrQwz7yF2FyFFKIzc2twNjnsdlazpWvD5SHrws5tHDH0SApWh247Wk8
Ow5MwanhHMkWamMzyh6qJk+CBv9QfYeC7wGplgkHddRneUJL0uk5Z3hzn6trcvJp
jZqTx3PVzDyRGvmqFWdeAox7u8w8fqpKG5QNhP0uCpooH+IokPxtz+U1JwuEy5ok
ulWIRitofH8OzpdpWirTPSvoV0622D3C0sGfLZ6cOsiD+L/D1lBGBaBvTXkQ2MGu
OR38v28NSU5UNvxeGcOpgbSKAHBIQyX6mC3C4VxgtNAyzzQbH1SEJW+MoojIqwKz
lJkgDTYsfomC4zKdWxKu3uSvhr3CsxWvnXsNwPOKl0A0k11mUovdWl9LT+ts2qRJ
j6JUjBGbtpw4agtbsRfJvudPWbrwIYXnJ4q/gqB4Ct9hqz9hNX32hwjOPBcsW2va
5/lhRFH1W9rNF6ZRM8a8fw8bQOSYx1NCXrHqPd/70lCyGhKc0B3mDXYYi48V9AXG
PxIZa0s+NzQJnFOwyTxVWpjJukRfSPgbBkZ2oCB2vfhzqvn4hZxdjVCkQDsF8cNZ
cqSxv+z/Xv6KO8he2+AmBxWfHqsuvHm7T/BIrlAlHTpEV0a8sgqdDREUJZRT6tIY
tT9Xu7+cdx3/4z2lZ7qa0GMUGmQFAP3BppMgLRhi05kCvg6XCRIIQPAa4iA0Fs/c
jorC04nhpr4/t/qy94MntObIBHSrdqo7MSqX9AQXGV6CP81RWKryMU81OsRhcRHv
AeZ+Me56l5gqlhL0gBFf/5dC6p82GAq9uldVk7rlSLna/YQeNJF1nKT/LWf8JLL/
ILKUMWOiQ1vreKmVLeG+3/7sTkIRtZC72OX3uV1+l330k5VsgOHeyjo5AKB77PgQ
VjQH7q6/gQ0b9VpcNOrCz9GSe7yeQWAaRHUIrFVEFPeNDOTO/qX08YlyjULk08p4
NMQg76m47Ap7RJfXhdk9LCo88XTdHH0O9W1kMpl65Pycs6sJCE6Jlmj88K0RbPx9
hwiS7DlPVJFHQKcjhb3Vx3y40QcZ/xDjv1lth9fcejyahdNDrnQnQ/NbJCU/BpWf
WB60hOxA4afJgEb8OYnpft/6KjXGWWTWdRxd3y2QDQSVBqr3rwwhloQL98pXJZAs
kAOdsPJYx/6YwAnT86IQGsr/alVJxbLaV7oct+nsnRj/zJD7pDBN4C5BJUVWhdld
7r7vghutNP8wNQ5hVGtcYgfjmIm9WmfTYWOIMA3gXW+fuwJ8+jKViOjtR37BZuMM
/CbewfXoXisVmOoH+PvdvnX+OVI07ukuUhLHLEcAAfZZRVAw5/qd70+h1A7Ezy7j
56Q5206S3kJDanUvgWARttYuXLwNZiX2tax4wUwEaPb1Izqlary5lW3+QCX3CsFZ
u/Uls8fFhjo9BmFN0sAgkE0lghSfOwhIvThGBWkaF1l0iu8KQBxNvMyQ2p3cxF78
1OfS8zPZVVzw/X7gchonQR6GKON3NhdHV2rrA7nDo8euQogdaNAMgscciTvjC+20
+9KPzPg6u7YjHS/QYfGR37XsSrGlzUDINkzFnYydvZi2uxVX1Fg1cIe4QofNfdUc
dAMnuS45YQ2jG93oig0fzHP6Xp2j+hrMDZrmw3oVSepOk4pO7jms5aWKmR50vqqV
CRogbnsxMbAMJ5aD0VSD90mTlGXDA3rnT+upAK9WvFNstpUlXGDHyCKdrJc0Wu6v
y6/UGvlXjTB3e9xtHKga8G0KydYIXRC4WZvhRGh0TBIFXS0l894oifZD7OcoTRi8
dPQzuuyiwT1fSDe3cTs5Od7aqzh3EW4lDE5NqjwhuRi1o2sQznKVVpkZ6bMJc7a6
+oh/tdVhuUOdfFMTnGzcdJN5ZGsmOGSo9kA/jb7hxAjFuZ1utqc8FAWPCmOnU+bi
OzOSMDP1Fdzb56bQfCAh3etQjwm4z18m0rD2gfIUgMpGXbJAHOjIm45SXNWjEo5D
LkmfBvzCWlbX28WsKPqVNKzx4vIcQPOdljMi9ypC2UG15hjRIBeJsgfw6VN0x3sl
l/rIpY/m68S7aceLxYqqD5Ia2tPtJkeP1FnMc9968miwxDrxhNrtc2DMFfjEV5/2
RlAG/0nhG16QLZFtfRmswjFh0J9HXlXgMeNVHZAu5qtuUmcWYNz/w7ow6Qd4r2X3
6x47GfRmKfIv8HBTifKyZVC8NA11CtJLrJaJHaS62sIvKt94AtYnEp2UECC3uhXs
dbqCkgJ6O8ukZLIF76+2ozhxhk0DLDjH3nbB+TmwYk1/tI/9BCKj2Jyp4QeXHYSb
FU+NhvHtp61W7/R2zX8z28hrjDrYrYWBDtCEAwXOmsFllbje1BEmFKaw1XMlO0g+
KLP50nKVEPJC7w8iQEHlCFb5xI9YSMDf6Yv6O5IVxCmZTZtNqKK4BF5ErS9HlpM0
lv+iTemi6OEPOAobCg7QkHUEQgZzczhTlM4tfHmGQxwdzP6CRIKmTYSn5TMpUkVr
VhETdR8WqeDQIRFnPb8ulsJJr3aFbcec/8LjJCjZ0VPiV9WN/NFBrte+IJzyA4oY
A4b7bLauorasupmHml0t1t2VBTSb0NhEvwazQrfPAMPjROPwliOV8yaDcMpmOv4L
Tqajcr5uCTKrzUmO7R7y9l2YJIeunmJTfSmS07KdnJzXAUbJs/zbXniJeCmLizMv
O/ydegXijLwzlTsRrv08lrYqv5Ze75ymEENi78jPS+dV29uL+3x9UIc0svdb1Qco
3Oi/vE2uZmC/zbgcwNTXNcH/mbG1oCMtTd9BlSuqdnLYTvFwBAJRadLyFjktiWBn
P/UxRfl/PRp0xpcCoQF+XEczCp9ySSMcWrqqsRwtetHyBs8rTUXs7C3nu+EGs8qy
niw5jQJYDC2HfRJsu9rfPb/5vf+jFxeJ+KddgBe3VJN6pO5m5wthvKXihbwM2z6h
XSznZLO09NnnxRusdi24AeWYwk/BE5eW3F1iqmFS/T/53asMGwgk9/ajCbjmDYnt
MpoQY/TCOWYnclatpXdO/BfRbnxQpgIUq3dgqPGjYJrYxlEjMvpy4eFZHJvF8SpN
EAHSz02RxllE560Wdn/bTz2Kef3PeYxLjx1spKR8Z3QMDy5IY8qiYJJAyyXQ9WDV
B6zeCFaC+92TkHj0YimFJyu16Erz/TYlN2CHH2oIGIgey0KTf7z3M6A9hgM3r1ao
GqoZolrIkRFggj1J2dx62gn3QoNAk+CEL1752jEx0Ra6yqxr330BQiq+T5sHUFLf
O4wJNZOZxtHG1xIZw04KS+tW1oU1SYZ9OsVCVIiXkZK171+Unc3ENM3EmuXWDtNU
bDRctR9J02DhJNZ553HummypdSTgSB2W97UXSVw4RDXlYJ7Q6W+AEmdnYhqoowbP
pKxbqZGXbx7nUAjhElDe4LYdaUxUXagm+llnPmwzAZxzn3YMoOXqtxwCrBtl+z13
BbU2MD0L018Ze+P0lbTymyi1u8bTqhj8XxQ3czfdDN2QDDZ+0DLYx6aKa+ZqW/Rp
pbo9a+pMxYfgRJR8ChqxIsm1ibd6m05jHg0g24HyKjgh4Y+UP8sod7bSI8bArgx+
Aje6abvksC5noo3eJvnRB2bNr0vfwF5/lOWd3AHt3nGAVgbtpmE11c/HKou4wif3
zBn4U+jKYnW7dBwpJhoTJMaVWPtHSllqsZFLgCj5m0kN4ZQ4h9/iTeA7KxmQBi+h
C81Dlxr449esu8qkeaOn5+eMDQvOKg2cHCQGrEhFYYkDDAEql6ry1fhFyM/Zj/S2
pj55Ur99oEuO+DHOEmShx9977MItw3Q2Ao2c+t+3k6PHhoLL7qOgg1G6almlzdJY
KjKO7g14MBuh6GjeyZu2wBqvH/zyIkAIImFX3RJudwkrFMCjKbTguE8kQ2jli2BA
7iNR82Ea8K9AAJ/dcL/9F0OQqDMaXnhOqesB2HhzSW1Ud8nJzcIljsE9ZHz1xqAR
4Zi53PfV4j8tKeZjBbP+jc4HuGgwQRIK4jqdl3XutNF9Hyx7df4v7z/aXSiRRs10
7D9x1mmF3cuKOwAxq84OSoUaF/TC5HpkBcVB9u6AkUjDXCSPW3rJYOzA3C2Xvi6D
2Iu6AtCIKKerqHG7mfUkas5OLxxYp9pZhy3JZCIlrAe/JtjzNPw8TRSrYfAHb7XR
0N7eXh3+EmInJc8CAzX4zsWfmBQReFx6gxCgh17teL/JbU/NCD/Bw2gCvddkdkaW
YBZV3l5gKiCxRw1g1l/RfZ4TMdJVv1ykCgOocF3Hn/PIfeYNJzKZbPtSYkvkN7jL
e/U/M2MotncUysXG/kYpB1ZDrjXQjhXJ0gJRpJZP45ElLqBe5pExcbGRH91Z5u8a
zHzSaSQ4Dftmx66c3TBaKEInSjH9HZRx2MOWLYT4AQ9tpZuKUr7IvLJjsCEgwS8g
oVMg9vhwaNZfTxjL1xeF0X1DWGQZS9RdRucoKmmcAwdHUVlBkZO8/O07KSMO0MgJ
WL1F0D44agS0C9imfsVEd17i+cX4r/WnSqMzqhHiZHBiUC3G8CTeBG0vb1nLbeAQ
A0p7QknBJ07GsOwP57++xuDhuCZBy6iYDORJfg/jJ1rMAayAKWXj0RZNpge66LbM
swUTvVPo5fFx4uCRpA5hAGKpSGKWxQ4k3pMvbJ7k+Vp0mYvA8eEwVEMGOxHE8gaX
CQc/GSw8JY53Yq/bhGJPDrsTc/DlxO6Raj/E3bk0l5n03kglZHvXongo0fRCwrPB
UjIAEfaaI7qvhgJx1b3RuAJsF8lPys5/R3QDZ8un/L4DTQstPqYzgSiw3WjTj6xj
rhmuK6cEGFbBNacclQFD9KPfA4WY8u5pta8mLdiDjOAWXeXjB0XrlCX0A9IkZwMd
Lw/SE3xfwRBGpsi7U68Rf996uXUWaDdLt+x44TJD7lV3Fj8Uuq6h6vEnEvPcD6Bd
ymyAkunH/00W1pHafCMFZP2UISWFFMWB8v5EkzXQPeVWtUm6Va3i0h5IjvqcZzff
T5ZUKZLuYsfm5N09pLC3h/GAoIlYecK+DafUEMPgN9QIUipTFixPh8rP3gihQKVQ
WqETYE71usLVcrnjR/IrhLwdqGTbHVnUmQg037H8tz55LrHDl05YTtaxDR2ww1D/
RtrGA3zY/VX9AE/5iZZijNBCs+R97lp7aqHAveavQtF2Y1Ax+C1nCqmIrSrWBwex
63/8iVoCl7+YH09kZ8H9EgM2kUfN/JUNLkkYr9smYDP0/BpbKJKCNzm/Onu+D08l
RFIMRXj3807ymsbUz8S0fkdeD0zEcDQvVNAsiYsaKGzQy55Eeoqzq/GGzGTXSoHH
k9NlIPz+297RsxAt8L2de0oKl4kuhud8RRE4fsSe99dzV1gEPI7AFG2/c+t/b728
anyHp25j+r9NO8rda9uhRgIagESPPXvrZ1gS76YqY+JmGN7SDEpF+CSnLswLt7v+
M4yxHc3VpDLQ7xNhFS0ZO0os4xkbiiBmL4zJfC8trpeqrpzrLqzoYIHJzlweMJzV
Cvn3m/ONjaljDb5pZrwzzUdAVeXQysBzzHTyBEXeE4DRttHs1z9eqHK3gVBgddss
qhvaJRtiF+lW1Ra6DtQSCXC4KePXkCQ9BvjpWnVr/E9WJu0dMT5CRZGn+YPmnpDn
qHH8ARXf3p3fwHuyUcb8ejyS2hTVzv5eHfIGrxdFiHzuy7JiTNC8e2PbZdA8z/S9
1P9wQWQp8hy0B5zSMGaYtd4eQPTPmeDNuRV2o4UNlWMU2D9MWSRzeuih0InhqDTV
O0KCcncnN0XlsEq17NwtQ8r4K/WpINaRdCcJIYJhFEkmi9zo7wy818rQ5J41YEj8
VbabFYY2Alw2ZY+bqFpXM+ZiyPj4hiwZxP01Y5pXgrGDQkjPcnlioCTSmdQI5NFz
AKneBny/bQTUdfgZKuQfVjm7Hbq5DgYganqqNshyF9q3S+jFtWe1hCG2k7f11LBN
e/A+cRC6SIwxx74v66Y0cZeMWfksS9s7R56fjHrlb/aGu6UX9H3hqwJlJBmIRhv4
IunO55P2OcAXt+R/FR6gNEQ5j3V/DQy6qEdQKWnIjGko3kIsQt9jgh45Pd+1Varx
KV96PjbhgkRC9WdBDssH9iVyo4c3vd6EPx0Su48c3b5i+dwUGkzJT6SLmiafPX/m
47riJc534kftNu9VhbeG45xMxYSK4Eirxe6b7RQrVk6rGTzL16LfdA2qGAGJbdvm
ok7937aOBEZpKm6hIIxKhUVIkiyiWAJ93J0FOBdwJtI8Kv+gldKf5fjG6XZei00E
KAIyrMpIZhvv+Ib5Xp9FlKsIgQp+U2YuOYlsAROREShsvrzl2o1bCuxewdUhVxWz
TL2BvS4buTL6T6Q7Q7Lsa3itr4rxFMGqG6TtNIUp+2m8tcIQ7hTzgxNhmx5O+ghj
7bn1OgWbHg7BW/gm4YG39Z55yypCin2TPGW+jPcBH/Lm+dsCt3bGS0/7G7PxlcML
Sjfe4HBaJ+YoxJQL39o0X9gl5de+lMkPHfOu6wosEO/Tcbpa1fm8nVnhFRnA2qUP
s+ql4ueQG0ZR58WbpLbpd3QxTSNSw4A3bha8w3URIjMECTxwP3M/h5FppYDggdUc
6cb5GaMCW9Dm6aI/3s2zLC3TSSkgtwldqDOJXrVOHxpl7i/cn9aSPRxttJBsBmny
oIIpgCUnMb+THlFmNOywtzJ6ia6ZWu1/jQAmnBTgeAAw1Vzl7cy9pnqZWBsNgT79
4Lj6ivlJk8cJHA+/2q94hteve+Dp2OsGRc/l95ny0bOf+cZ+WjJnRgcKZddE00D/
AKPSW+09IkDzQ7WsXNfBkkN0D1QOJdJ2qnXhXfKo6HBTGSYUZhSS7MsyMjehJ4Lg
wZY1HHP0Q3HZBjowLRJQ30wGys4H8atK760lRDIyxO35sJzcIjR5FxfFbYbtQOya
jOzl0Ynh0Z396BWtUXZdyECV+rV+K80nUrA3Q9BgS3pb0vLSSb5HEEp/wmMnWqv3
9/GHBkSMLcmPjMGdrVAsl0OljfW7O7Uv/sYl6qlZYwO4RVvXEHJZXE4xh2j+vzGq
+DcV3UuSh9u7gfWfZ/DYQRErOxPWROLTT8hF9TBjOD5CdrgMlc/BLgbMP/YTlpAz
qH075X1MgdHfAFtSqQbitT11EfCbcAMGWbZgNbtvtc7XnFt7wwdbwhT/BW+Fv2gO
I1yC7/D2cyTqP872IQwyucdQ85VjysraY+Nu9zquUge/4+Lt8rAB6wjvVh9gO1X8
SrzRQZmZlTLHHPgSy3p00nGussqtfrp05yB/M6LjIDeXOedUl0FOCjhZKrIjjoCT
uRCcZvVBezPspZVGpbUkyx9XOSDnFqTv5mXIMNzqwtryS6SnWAMKctXcoIPps+MQ
ZwCqIg/W8A+RCh1zJQ0G9OK7YIDxbrDP8w+IZ2/WW1A5x2dPSSLn2pTcIlXT56hL
fPPaPGmaGGgr57QZy8r+S4cUxUtvYtUpFkOajnu4abaoom9wLq+CHZ9zM+Jbd3OK
AO47ifoHRHiUBsSe/zfltH431R2PVpnTVIDFElh+NNupmjqG5yMwNpslYMKLXSDR
T9iA6Fpx9dKfEctKsIVN4BlYVgitsrJyMBZJFLU+xkB014eZUaR+k9J776cJEGq9
5MYthgZhsr/QO0iQBv2PAL1YXN1Xf5q7vtGEQSNcraQtlKaJPYLNCQK/iLxKyOEa
RFZPt28TlbrypflQoR/fk+q/34BpZkHkzVeywN9njxGB2MutJsqvpfHs0gyd0BIV
q5GO87pDKMuETa18iQ0onOuSmkzPbgliTB0CQaztI+E9cqdTX5iar9ls625E97UR
CIAPFlgFvnLsqss5gD8MSgF+bSkaPNdRmd9uqvwCzVd5XLcNGSt/9qXValtV4xi4
o2GVQjPZROd7wEfzgm2snovOgW8XbUJHEuOoq+ZoSxramlPER5GEYFfnAvXtW9ec
2mAJmudBdGxPYbm9EE2iTmcvTcouNf7vLRenoD3fKFjKM1uBXGmA2D4d1tpfqTtK
M6PMXd0Npn1JckYJDsawglO5SZXKR83MWWEfFMBY7ePaa0MBPIA4JFiHcFMmfegR
odsGrp1Ab523YNP2/lFZkQysNvQQSR3Q/zUj/OTAhUdIMj37oO0OpKIe/7IFYcyC
/Gvi8P1khY4Vz4kNDA75AYehHmTsn7FTNtK1i6Ps5s53mJMcyXXyGHWpmhLw0r+f
SH1OFMRk7FfJ6HG/Wpyh9fne9qzW7HUrvacMrU18WlcMIBUuwQdXXuTMpQKOSfvN
WetU6lG/dV9+UnK1YN6bGsqqTjxNx+bG/oy0lGjPzmJdYsTbC1uCIcO/JOqScehG
u4PTw3t4rO5rfTA+GMGiPpHyKZoT51rdB73KaKYTf4zpxmRatU7WGRzzy5uxtOJ+
CBDlONUC8sS++HobNY81T84MXirVXzqADdAKl/pOAZRaeNAw/eECvAqwznBysFLc
bft6obqPxM785k4KL1rXdRcBRsMB/efP0AFoRbuLb0I37XYgeKQ/LnHQB/JJwOne
Ef0lq8ciYuvwQt2xocYkP+tLuEYIqxDqiNZip9NyBJl43G0Y3R/80JUh93U/J40M
85R6vukIcqdNw10WGqfM09O43cuH3oxal4uImlPMnAZdRp3BmSW0y3r8parqFVRg
XVAramFVhBGUC1etLotAXucnwrFUV0m+MJ9gXcasLJezjPYWBKkcAnHuXBmfq3T7
oEekvee/lxiCikp399JbqJqsNnjdrlHxuDaWkZfSLHksomgaatO0f9t7OPKhdIOP
nTeWCQ3mKq7tYMROcgsJciNuJjFvrZS2rNjVvqDtef6Yz3MF1l9BQ/iN+ZjABelP
3GIZb7h6axDJiLNeuZ9U91XEWxo6jma3AeHi24rsMzfxRueQdfaMM3jk5FUdga6u
v1HBNpOCOI4b85+MLpwanhl1V+/yEqMOqVf3z1AA6VpSTIdvjfTCCHfk599pvgfY
13yfy69Jb7nnziueh8D0AnUfsS7aYHalz2ypzKw75Z9SGQwImxhZoIbzXLEyGDRK
Kqnk9CxoN1qFETkcV5q32UaIl++swhSYempNwJvZYazTJ7z+xKmw/Vb39gzTWbvk
sii5q91k+KXsZ0L5MmHNQio77e6i0ZMMFnMYvMxbz+f8O0qJuhXbITkMQn8Cl/41
cC7n86M6ex8/8fo5ecGUJyd0HAATNbnH3vgg8PUriWceKnH6CQEuTwsHYN+Mscm3
HLdXUOOVN/UlirPYpQl+AtyUTX24yQcP5s+rGa+FrTboYeUNkLtE2J0k6JpLWWe7
IlubBITeM8YwmtDihyTek/Q8kBi2l0PB7txYeueSesr+D/cAV5YgQJX3J09j43a8
lDVwdNeP4Wz/YkqaibtPx+weK3d8r7NF+kqlC637uR13E30GCmJB5uxK5Pn5qX/T
dA1ZSPoFJ5+q7QvszrdD95EZKiCGCzcxkFe0DpFS0KkVZcroOXRM4m6Z5d4cdQe+
oJU9Z031jwjTjdBI1rPStidB/ahK0fFTpovDydFCz5Ungprm+wkOQSDYRrQ6YY7X
P8EX111mU10urGFjdEs8LV9ydhf69P4NKw/x4dkbx9XvtSSuN04R9TPNXTFpSeDV
rLNyugZ+d60adf7F7Qm0eBAq468xoBJgLRmPUzixHsVTasrllbingwedh7+oTLV4
lyENXSHK0kWi6jjO7dRqe+qY3AwRBSWD5Nh5womeT3gWCfsGar7e8HS0BS+1nc4T
BPLT2d2QUtU1OhK/WxpvmlY4s7pcpXV+CMeBRNyccJ7MVD8rusJwbTVbrUGn26c2
ADjKjWGajlJYYyuTF8uksYlfafOFjNla6Qq/KYB61B9WKTLqoi4s7EDCxZv2MEiQ
DtvO81mIxJD0vPTv9L0yyA5kvwdzxHoM0uV6xUP7X7FMaavwonZj8ewr7/vK5l6g
HzpGo+cPSpHx5jx9k1NPFdUnk9s8kfclJXHwOgtw/vJxzPtbjrDX/PpvzhHie392
8bRKUBd5++ghbYYmvA0IcI3DjY8jDBe6Sx+it6YpF4E9P2uyvkChWYiQtHnUXhYs
aNwyW2Ms2wlnFCsAUa2T4mOCxVb4nC6XVA8ADSl6aLVRJ4IGMLdd9HyIGcgyot/c
TDlG2whjEn7kctVqHghDMuGHm6FomHr5moQIkmHgQwAc5ARcWDyp8jgoDLxjvHd4
1eGr6TdWsVjIx/EO7G6ZrL47Ln11qwBhBgdBdIntl248oHN3OSMYzHCmMUWTSaYW
2zW5+R63oO/FWnEZATpWNqmpLVVvpbEyymgEdJ+QseHJ6alyNGRZvvaJ1n/pQRlP
8LRR1uLcrkx8B4Y44V4n3txvTxfS1DFLDYLIW3JyYeFIbwbHz0MiGRnmLOFCxqv6
b3fEVjfVnV71KQuTMDqjBUII4obh008l3M9y4cRFa6uy2sNBW6er94H2znceO+6b
sbhK44YT1DkXql/rFBJtSdt+MTIpeyk5SXtPJNbFmQ/bcvSJbOYJW70mOkauiiwa
FJWXgC54E3JzImw1n/E2dCdGOdjkDAbXWflkRTBtRJ/zBLtzhSYsJvkdWj+OjcQ0
NQljOEkD02seAJPedFnxd2ai9YVxR2qktdTP1uyX85O0bh9BfuPZ8mdkWLQUoELr
+2bWt/EJYbHaYquOpu4+rVr2HAr3bGLh5jpSmD1YX3ZiGYNsWhnSEA9qUjEOpR/S
telBgNS7zc6iOCdfej6chYLub1rSdO9hkWCU8RRkjFcE8xtMAPmwS+DKAXaVxBpX
eOudr9ZrGKDu58uBXX+qfRM7Jq/szyw9u+RbIm1IwqY4IxyV6xUGFacIsrmL/a1K
yleA6qgMrvq9NUDaIarFy+Q179/k3JJE9s50f7GgzfEJqBZg0LZ1XDAjbUD+ufqU
szHP0NFntqYVbaUVppvI51qXRqMEOeDn8WTQ4KzKaHGIMgp14sE9SBULaK0WLjFH
e1Ai+aqymD5OgDZJDCpt9oNuVCTxKpCZYLVwmbHe3MoRL5h5/VDPtzIwAI8WZKuN
3bhCxGX5V/LtRESSC1IdDWw/r9mxZym3GGUP/djt2W6bnhvfdJq1sc1jAcbH3bBk
9QCaWDcwUE8H5CweCwJbRNWT8l35sWrmRZaxlpIZQFggdKVS3cVpx6JnmGFfaOCO
1vwjC1rtH2kttdXVLc7iJSmRNz3tclKfk+vlk7wEhw0lkHnQduZXzNSmeIJGQNRI
ocKyiKSRv6KLSV3Fr4T5qRRnwT5yxsmjLkDDsl5SdHD98rsu2WXnetIUMu+SJvR6
xq/f/pKWTG+UfLyBKtFre/ED0HfO5c9smWo2wzsQHmg+NwORWqeIv0uYUd9BhvTS
u7F5cBB/MGmV5Skkmjb/tyRaZA4JlyF79an+Kw5A7lN/6Y2rr/Fhs+eOynafX86x
8PuXZK+0VECI8Q9d/7TvMOr1YqJjL8MfNqwsVduRnaNNYMKgUTtuQJGKjmvTWQXy
uBJDN+neWDHgQ4fumQ4Xv9CGn3TUsfTV3sjj2C28jc05XUKb9PS8om7COaWQ7HNT
mwD/mKObdnI2zWdYc84NaNOD8WGKQlfe4Z0uK2tzRNQ8r5fi5pin5CoIoK/rbqeE
7KJGwsC421E361T+ag+OaJvCCoImz5eQrFvPNZqCgF6B7+aIQgxkaCw38aBPh76a
A3/ZLixn0waNAE7XAMN56w==
`protect end_protected