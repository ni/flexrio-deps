`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aMReDmrPskJscpWYThVKVItA5gecPPZO1R595p0GoIq1TSTG+UxXhmmUXc+VYHJ3
u/C3EW5qePLufxmXxmhmDnr9U8/cYC1zLfk44v/2OPb1TBrTsludEDQZdGNWeV9l
cPUMSIfZ0dHXN7L1M1E2XtgoTWQxf3VDHs7B7lU2y9Rdm/ibz0fWMow7op2nWdD8
gJ4QlNl3f9Oiotp1p8vz9RFzzZOF5gBBslZxcTF5+z4qO2W7+xLByngthWm+exIr
3Pzy8qyUo/m2DDwOz3VJSvSNm7RUq+0/yJNOOz3jr3j7ZyCj5OqT/jDAWjJSMH+i
2402Un+wDMOQxi21JLo3cA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="5R6K2aWI3OdbT2A+sz4o9+2XAInTqB1/cSw5W16RnA4="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
Gm/2BIZF5/H5qen8uQizPH9RftTuEE9mgEOF0SqeOKegtP64CfvEUnIxj/ahmIpA
6xUR2v2l7E5duaLZh39Mc1GYsfqE91NCPU5whLaBPg0UuX4cgTkO4cYbW/7yvcrd
4wavUfwXEp2VSiN7EVxL8RcZTSMSI0Jr/aojiilFqVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="TEmQtJ1Dsm7TOzpJk/CeTSSFx/zKExk04H6I8sT4Meg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 34752 )
`protect data_block
nvPqn26PC4XWLLQG0Fq8XsMTlhB4evbpiwGjZroFFLgtNlE6bBjdtwWsB89WW4j7
jNfYbKN4sBv0hDeMH0AAR+8g+TCqoX7yLdIUd7aGwBUZJr6FdDs2wTUxRkXFYNTL
eFlqjN2vMAZ04vmMXbY54ZiW4VYgLZVE4lFE9wKUDyjiAbcl9MDVNlS156vACxnC
jpwtuBSn9E0ZRncGt5AVBC7FN3rfyo+P27m6HgkAm4Lm/Rv+/y7lmNjeA4rNrouu
Cp/oynIixwcPUoGrcEx3VkRFz3zU+6ijeGPhsEpXQLcuholeQw5sPA9qHzw7VkId
0FZpM5xXnJ4zOalhfh1w0TjsSKL+T9lHPrl2jOm6xRVH3LpUhUqRaXfnv099YCNH
o7GwN29/9Yx/+ajcykNt/xbNkOWoO99bbbBWGb29yOrKqE4oJcCf+Kv9rqDz+Cjk
aS0iFc2VXfDoXpKcFZ1AGolI4Q9hQIo/ZSC9B+oPUpRHzw7Uzrd80LBntO1/F6LU
XJHVfdFNWNDi1ZFijy9uKjZIgwLBOHSsMFoBOPZesMpXNlsDI0Kru2NLQOQ51wQm
I1EKftYQueUVan/Y+7sMwtxvd1q1m98Jua3gWPd5TaQ9Oov2vyP5t3cQT6x7z8E3
bZNRv1b5McTbXDrV+agd4/0KtmTjoEM32K21AzgtVbbZC3zy9FjA6i7gaqFANKpR
+tQ19uEZGc2xZFceeIV+8PTqqUN9FSHTgeeDa00XBhlUjsS0Bq5ClcDOZxGw58YC
KmdwqhAib31r1jLTEEYunM9g3Ld5KyOfUJP9YmbCDcG3NKfsp8aR11h+aoFtEomT
0gGqqenRo10Qyiulr5J3QcYO7Jcj6draXE2vtiKnDiTnn/DaxpsrT2XHtcjNmDNr
NoHxdE1G/DC7UdxMlo/un+inNxVgIdfqcoREtxGm9W0Oj76SjwEANfJgciOJjt9G
Dkhm9Q+4N0ZiXiEyQWPCiIW/sXJkVUt50wmFjIl95911Jv5BeRHq3iQ7+GMEIsRh
VGC6IJWg/Az3nGh3YmeDW69EFf/VOiRpj0Gw+ENHOI1mswd2fNjeGHtDV3OFM8nl
/RWdKcyxOHn1ioExOndA8QzIhNcy/xXBRZq8c1Sq3bgetKoJiAvJG/RiTchkH1RO
VBmNeOY42scaKMolkYdZ0YpTXx1mBXF3GTHOOpasIsJPyKBrZSdRXtVsLxzXn4hw
XbS/H2IdD48KTY6lnpJKdMi95AXOzD7q2SHvbttISYrBEklUVSJ608ei6fz4OEg6
xpO7re09yhxCFrTPGjb/tX6AMAvHlFGBdjZsP4PRzpR5R4TKZKYIl7jSVKpsQ565
iHDZq4jvWox7+UEhdUtY6KupyAFEI05xwRzIvN7oQg+R9tpnCo3lElEECgiYxirw
zG3p8BrDVW1JiP+fZeRylDvsoKdExMNkWCt9+mboY+4X1y9ySjWakswMKvH28wLu
DI3OnH2MBosEQMdZW790SDWZGu1Dxn2zrTYUSPEtrji7bAz7Z+iL0LPjvf+MfgVO
IINl2GMx2BY6x4uEv5ckphRtgBpDlJPVXW9qr1e9Fv3BzunX56ldd0xRFVIxAf2K
kHIXerrGwCqXEshMrDRI49vg/D+kAe0uvsMlzd1hPUwKIPKvmd/X25gNKe2qfQJx
jDRzk7wLP/k0/frpu+jzaU70KjXrpO+nwdwkJ4iyVMsj7ii6w/W/56MQW1pFAGl0
JX42j52ME8HOgD5zZ9gSGt8axotfm0IBX2hRmjSKz6TOekmI1RY4Bre1Mqkj7tea
ghVIArW/o400o3mt16l9BctZNxC+m3Vsu6PlB+TL0R+UeTy6WUZvUs/DvjsnS3Hm
8uK1qVMOG0Uht4oAVzUwYf4HHceP/VK4PrrxZHMhWjOacNbisuz0fWslslTC3hDH
wAXErY1eosjLnfvldMMrG4K7AyVK7xdwY3yxDs0pWHHOyIFjjGZQaJA63W6DcIu6
jcFTQ5Oi1I2YwBOdHoPx334JoIBaeNbkEwUvRLosRwyWuywuy7bwL4YdFm9+lSp3
2/YilJya5Ye0sLiU6N14SVlwY7Bxi9BN8oTSwsQ6Ha14320NIOUrxL2Imkf2qjsh
YiRLwHwTBs2Y3tN0EPkbOFtVy2+PNCP7XPnde2UnbR2XQ5kKTo9ATBdZmHVrFcVv
eeh3h0DvZ7mYPinq2+fVDJU5YWlD24pr23LuYOyL+Ml+zpPLiKvcE/qmBxF7JNg6
6+hLmPNf4763mE41wCPbGvXpKAS6+IPwrphTx1nFYSkmaALNBMSZf1LVV5h3RKhQ
efjPnTYXHPUluWgYqcSTRIZxRYq9agN3puge6Vpl9lQm8Zsr9SIpg+MaGlTjQW4z
uKfACSSeeCoijISx+BS1UPhG7hUuho53OX4FRGtSP4SfSevO3A2UYKMF20AQ0qSS
YoF+ECYNX438bM72+9SXtv5wi+j9g7Ii8o6LO9d7r4HeLgPXu1Ke0YN3WCaWYhq7
89Ug94/ZWJObYq4Gpfhuui0gWtyWs72DkU+SJ9BRu0Tsrq8MF4R0gDWRuZw4wzsh
05hFDuCaUy91XnyqHe+5E6WiFCI84zAOvEe1U+UxSOGNfxNjMjixjDtLib+MCF2G
zGfVN/9T4b06/H0xMSRGGNKsetPOYEW481bFGBHhhxfRGncYIFQjU9dYO3wenoZ5
e1qWVqBZoRLqYCGDiq5nriRGtTkuZJ8sBf5vlef0o3s2Ah1273LR/+XI2y+cfr8K
swKEzb4L0gJR3X9kblecRnJiB8sR3NWQ/3tXM/kTC+HhXi3Oup0bkBP7qPaSh5HW
Gfu1mPObqcH6nsXbR5XutMA930Hr25PF3rukg2jZTYdsLPerqR1pLMyaj2aG6RF9
b7Dc6XRgm35FAM9W2GxD081fv/idQjBvHj7IEuZAcmPbp0vlSPj2vsuhGg0bpOrW
7eOozmArzlWFhsEqHj1oL+6YuaKrTgngAcAGws4dBT4hMcRzMn2b4pTPXsohAxVa
F4h8JaaKFy3U3/RvHaL9g6set9/UKsLTfIc5IWtRNWRpe+fCyuNbxM+gIyaPk7KV
Y4ZuiUENY4aHPyt4Cb/meapDnSw7mWOTgmQfDpu7qHgW0KJAqbMwPKninDgadPE1
evHUhQpl5If2G0Fo4g2FqoMnzxxUa0NF45CQiCKYXnZUDZAQv0faJ7o0C02C0RaL
Cylkv3C2CTu2bIZ9nGP50ji3+Ytfsfnv4ep+gTvlmeRnbrxmoWVsaFEETCP048SC
/II5A8njEDZ40HKRKPqo/jOOaSrqoxUotqMgX6jphKvL1Jipd1tskjDye5435A6e
JA+VFwlnawWKLART8wZ05WyXfJlZuAynNoDUORHvuxDJBPjfsp2hV3JExKl1vCrT
E64l72QbT5tIGrNdyh2KmECun+6ldvRMIK8WSV7wzu2mI3sRwv4BEQQihL/BIxsL
7NY1B4HkIZ9ylzXYMiwgDcJEB81pfmE1A7zmV7HU9seRFDh9Nkj0gwYfBafnvmR0
xkNvHO0gjJ4H1mR3cwzObSZHQCk6QRpdMuvsdg8nhUNv3xTHgd6Yka5knvKfNSsC
chV9fuAjgBlhEn3DPTCwAsWuD1ZgC7QlLmW4b/8WcJhFwMVEyxBNdkShAV6ogv6r
kSs5UCVahhOlNMD7S2PqIPSrm1gZCS1C4k+U4FzlX6QPYkhbZA7gamAUqjZvCrvb
Vq3O/FTLgXiUL8oYxfeLA+wEUnGPYMaVkR7Eh/CU9x3LeS4+nVsIL1f3FcD18Cw9
o4Vp8wvOG79/TC73X18/jPm8FWMJ8ZVtDxX8V1WG7X7biiduDa6YOeSwIY3SxyEx
1NC72F3Yo7U9aISq4iLEgpJcfJu9bi9YoQgLNF56HMTNSfy46rAHdbiANULghxMo
Mn/DcZTJKJh8Lt0Z6Mvw+JnYeHD89rAvIXHCMzxuhJ/E4CslMeaVCBoPuPggMr1x
fPUwoFLlsThQVxg+paZ65vFzhdh+tGJ7ExbCU5D1RCJM+bCMWaP/6UMBGf0/xeq9
YFqcKBHtzo6aJ26I3wuAPweBYnONMJFPFkbqg2aDrSrxZM2rzNdAatBPF8yxrB+j
QWuYYj+HmdcoHGjSzgBNpnEtR75jhALRXty2G2/2d7hNOR2+foosCRCbKZYIFgib
yPz0KcGzWerjrCyNhsOlz3NLoFYt0b1mrVhW2POI2FHrM359bcgNJWeQLTihAemt
YP3bjbcNY2KteSrHmCFQszhrb+i5nDrr6/NcKA8HKsQ22Ktfz/F2YRSwbysc1KjD
Y81+p4Fv616/DGr8Z3k+1+rmcajS25el/59Zu6iKjxomPB3qxJEV8aqFl6/QIvWM
TrFjJSO6bCXYbEpU4dXtbvJpNSQkUjW6gQ6FYLe4ayu7zTIyrJwO4b7vN/KWv5k4
KKHSNAG9C4iGh1mMwoQkZSwCpwnmM0hufSchZ/9roiNUPa8Fm1PyAhQ2+KNn/HdJ
KKyN1v6Fac6fkAcWQRIAd+aBd+067tiDZcTS93ZkGBoJbl3AkkCgOYD3H31IGtac
Xdt7or96mpa7WkB/3Z504l/skJGhDIHPAo+zaxnMeG2e8+BM74K8Mc+yoZjFKW76
yqfIW0U0zzgBJDu6V2wCO7X2oDKDfHxC0+ZJQpSiCDUeh+y6hNyFK0y8HICRHn3B
wmU9fSHOl6+UlU+m9XHsZv13obwrnRNbv7K3Qu6D+scqjVpTGVCMrhnVZCADjUNV
boBxlqh6zrM1geVN5oS6DLgl6NNwK752uRHgmiscCCogZaL7LRzzKcHQ3GKHBTmN
ZwCBcHxYIQbJvNHy5LIbAWuiu7YEd5fjE/HUcZrmqQphZ079nz1Zv3QPZs60wR+u
Va6ukIxSNtpN8VAxuHT011ptNiuihl5hvlsz8JXGLWp2dlu4AEj/t7JGF2EQHwcA
X+O/g64oZf3vITt+ilsQ1hYlgOuIzMo7VimyN2948fWthhohld8dmw8SBh38YROv
l7OFU1h6kBom0Aek1J3idYFQkzzZv8kCs8JpsJnh66JjTIJT4BSNtsRHOeBt6/Ta
XXzjp9RiFkjbZCWGtt7kZg992kUIw3XWBxWFs9Bujaj53xHWLOjvuBfceLAFCcbH
6jqpXC+deGmbvpigpFv17JFXZe7X3yBKGzHss/jcVNsHuphMh+hdElPaOXPx8BfJ
nUFNac/ddd4CemYLfFiiYAJHP8ticORcY4v6bJ38UH3vTXFWSFcqUxLlWxOpkXf5
IBb5dPlgeu9rCFBBL9CAQIMIO9AbGdgQqMyw5YZP6ZWMdJFJuUchcfbufxRT/QyW
vHPke3gBNI29xfa+m6Ifhz2UTFiVBaMDq/5bpIByca+k11DVWWCIHkOl78iIGDEa
goia6wxUSqgmYDZoJfDET5U2xu70y1GUPA1R9Lf+Se8nQ02QASpmHJNMHpJk/hFW
B3z7Fav7m1Xl8e3vdFCtIHKzivgtDfU8Y60RkarvtnRi2J9LC2E+uh5fJEse3X7p
oE7eIukpo91Gho44XpU/1WtPoGDipjPwdjJDZt9IoH9FXTqZmyVGWmyOvUtd9LqA
Y8oe86NO1qK7EN/Gi4yXmi1bxbFH+e5Bhs/NmcNoXkN/6phA1v6jns1JPLevYO4B
AXaWvbY7u/5iDs7/ht9C2vM9ERSfLDTGtZLzabnOmIel8SAkiZNiVFyAXi5BUDTY
S+ZG+/OSXwu0v4SsrPH1M442C2a3GQbVvTka+nLMG4V0/SjlUTC3rQPgLlJw1PED
3zxlIPun72a35aWNsOHByH0xcbLoECughUGBjOmtVeMh71xySCn+4qhTqB7rj4Cb
RsCeQP7j/9vxXmfBcgfBrTE3jAd+RCvShh1rx+SfyT59EX2sGxgiKwTGXi2lHRxV
WzrKGajnobXCAudxDGUReonhoXheR23zi7ITqk7xgw/5catHtl3XGwMIkVijPzGF
fFikCFYl/jVGQFZps+7Uj07adBK1bp3PRQv59WDNL4mlr8rMt4AH5RkRPy0zCUtA
u7wS33NrMRBomMFEIl4QKdeGwMgI2xCe/eAPbwyR+uuWvBd9qYiiBAX189AmiGm3
TC3rLsdPZ292FjwnO7aI4Qi7/Fl0br0MPMncTLZZxFwUKkSj0HsxUEcGwosf4nb5
OmXudw9i8OJ8u5mL2FkSQWcyf90SSpB7bxYcej45Nb1VOXN3JGRUwMbHPiHgMVjk
wM5o7BDRuEPJJ7pI3YNdTVc12j8KI5gl2mlI/TtuDu65IMJrbsN2YvKWnxbvEkJW
gecy1CKpkbvKdDPlRVeoItVLtG8E941o5EydS/HfJTw5Mqiq6H0JGFC5crABYiYB
V933nuE59Gv4PutwAe02z+EgbQwvB8aoplBSkvETRklouzcjCGF7Eo9NJlWrEZUe
LCapzWOC6AhcCcZXt43LG0LB+r3ueznhYGKTCI9O4lMsvZ0tMHUuYO9xil9Kr/rF
0yNw1Dhubg+Uzft4qMHMS+UKkgJaItQ9JnTS3AnqpwA5IazMWONg+uyi8Fvp4o4W
hkEy6FDb1vAb+1XorUt8Dom4MkezNnpMbila9ZNd9o0oPvCiHYwZJ2XfYkKjYNxz
zYyPErqIzT7D0cD2hmYjqoa7rfZvzL27lKvVPZM00B/WFfRTOZ4udKpReJWYoVbH
vBaoWJBBw0h3TufL6aYKJKaCJfzx4wka8S9jdDSPPNFfN1DYA0hEqfyJ8hcM2xp1
pk9+UhYdjj/r7kdmiX861vWPs62h7mM30oVNpOipITxLZX6IVoRne3LBxSsT3dkV
yy07nzo9itV88SnHCUeEWtwJvd0WBzwMLDZpgVN50of554sVlRvD4RN3tjxfogiE
vM357gVYaTyhFZq5uoIfl0U85WSk1Au6k4w4R99gqWiFS5v3NB8qmVctRW43QDUa
ciGpXgDmAy//XSWEg05l9wrmBcHrmAS+U30s0Dv8wuEmL2a305fKa0w/CQHl3mzz
eMJ7z+zxppbBTZONADSy+fG+tgOE2jpAAneJrlEopoC0pcGvJk5CLf5d+9iaZTdF
72tBmkBDgFEGNWl4fX+a+QyvM9A7chiHeOgotMp0H6HbJtgz38TdN7yyeok5SZHi
xYGNjYDVFYmVAKumy7xLKJDZ77/qFIT8oDQAJ5UXmtBnrmneA+XUSzQWUVMrqZdM
aAmya6jpgy4I3T/qC8irkhQBHk6EN9hZSqlMdYWremVyjonPcIbwc6lCZT35GteO
udJ//8XG2JTddYKU++l6AHmoNamj/QVRs5dHjfrQ2qij1vSFqDRASF+yQq7fFix1
usNXStd3h2XDCLJEaOYWNGn1Ay4Yd8Jlt7/16/ENodErHgwC3APX33wAxdYrgO9/
2Et5I1eym8lziaK/FZsWXnKc2mW+Zk3JDyjtP8tMGurNxcgdakpMRGbUEpM/E2wF
deWUDv9+LJYUf1lFufw4dqiIK1uR2CGaddCVBxAOB9VTjf9oCNqbO+xu6ovoWtzb
V2UpMX918EaHGmqDJcyqQRhRI4FG/EBxNxHxRZ/0ogGnDhyIJZXqHqBFl1yNQKSU
qpjEqZrfyTJ6LPDISRQcYAiDEEFu5fKLhK8dXDsn8Mmj7bW5BWm8wZqaBdaFILbV
T/lxOQWdqLNAH1Xz6kz4p3mROVPvG+/CACAqFQRn5VB4lzSPJdpEzUFGArrJ20Aq
W/0W539IKdjGgskuqqzK2g3QcLdHS/8VT6c6oLXX0syaWwEipZzUgS7iI/hBO/WK
EgMLagGDry766x+pvwaNzptzPs79/Om2uo9Oji1+nj+jWwr1Y2xnoyR9wXtBlyYG
wg2kojg9dsn7QrZvRnDbp/cPzT238WcRPaR5pbkKBdy7YkqJZ4OIiAhD+XvrTcMq
FTUkjnCRnWkgu4aJD4/c22daARz5zXD2WOgq4TjvL0PC08n//OOXvNONxRN+2N62
2BDOYVGReiwnb0fTbNr8axTIkD7Ff6/PYDB/sko+qBFdqg2LEHdlKy5Zup0tfvEs
tWZl88tu13vLikYKOpsyGB4+6yEV7dn+qJMMJTxIs2h4I16kSx6cAmqYTNDtVNzL
mYKB9RsgdJkY0AohIYigQSq6Z65IvsV+6HsEfzA4VXIk29u7cZnbcBNnnQRcGTOT
2hl83Rt0Vo8Nir046J928UtKRBizCr7LHN1cJ/YFDkrdhytTXJmLNv3SaUHdcPGC
CMImQQtUoVqPiERFAm4j72Jy6Sj7S9oIUeaEVomGD9xcZ/FRXHDojV5da6Jqo0xm
RWOFBB/aFG1lAyhg49MIsk6AJGHYYVdHaJ/SxBNdT7bAQ0OvwhnXFrWx7Q9W1UzH
WW8Ppo1UyfSvsBoPPG+BPCwaku3RsPw2ZC0Jq3+4GiIJHrKfnXEg7Dv5I4IAjuKU
bIXviDJZbAJKojgvWQB88imhfDiJKh3k7hja9GYvvcRYZI0nv3pQDSG/uXLKs8n3
NxpuAyS5p1cVLLkdb4QoHHZfbgnHwQOq7E5UAUhOKnUpc4mL8lPZvPnlAhDz34GD
T4BxEpZiTrJi4Kt+qltoU9Ots3QKPI9HZgFeUxXJwFFgOOKNmHryx3qzl7iS5aB4
ayyzRJWsqRgcEY5fBTKQvew78Qf1f70KHm+qZsLuQQndYYiyN0ATikExWcV93pjx
8IgndY42iLDkhhvTL9wk4r+/OokCUU0xuLCHMKDVUlGJRc6xuu1nyISKPp3V59ej
iyNScH8YwdxHchCOgqLDWNXYjkKENR/4D63EDuyL9KwgoOkDZY3j0HAuSxoYuXqY
zjW6hq3yKD39l4m8L4L6AFZG8JLn1R0Cj1McmBE4bAS6mzsKngKmUyM9/SRyqD6y
JCYvHe52PuU5pm30Y2BHXVcc5Ay/OB5y7xe+iEBO+n8q5eLZ2mUXe7JyoUEl1lwn
P6qc0t43ZCCfv/AQ+KtkjCUBQmneIVbO+Q0jyBW5DXeSxMF78eNabSPXfPuBX+r4
+8bI00/mEKZlGGTxVVgd4B7gTXNv7F2jWSA4+kFqmFv9c3GfOLxxgUgKUS+ZCj5h
VTpoCUq4iHpnioRYOqCVyeEhUaN+JGUpTtZOm1nSIzGSKwMD6xCU+OurK8se4TeP
D4Qf3vBxgPDOq/KT4lh1XdiggsRmGudVHeRLF8D7zlyEbI3ayfCVU/EL6FTPIF2+
PJXw95JafzScyJ1Tpi4c6cO8WnvTefH7HLADsLkxsS5/kIyLXQPT6oGkSP4wpyWu
84dUPS8mFn9lQA28/DTenNRZeed3+5ul1guwT+sKpITr99LRfXf/dPGpiMMt53ew
hjDPzYNbGhCmHbAKavtxZa/ZJMqMf8Qmmv8C5KemiNRx6zLMxJlrs6RXOHiphTwH
InehtG4+0atu8cL/K0HS7jDrvSWVCxqNyGxMT4hwpap/+61VRX+DEoWNERfIuooi
JqeGYURBL0Uwkg0Wons/Y3vEGgqAJ4RsVL0Ko971652rZ/yK8Y/elChE9VydbfOt
2SPqS/ZI6Vds/n8bTXqCq+hLvH3r2i6ZYHSZN59rAF+ioIWHVsNaWrR+EyTWXAck
7lCtIiziHcMd2JcUU7eFhb3oHxksD7eEpDRlEyZyZTc3dTiMP/NL35XV9Qprgfv/
So45ImUZAqQ2j3duj4shNoQrn/cWHrQzdEHygIL9AXt9OC0mQCIiy68kuHld78PW
wadzPDeNvVcDo6XuAR47dSqPQ5Tdsm45gtxzCzb2zjxag0qJSHR/GhdeJiT42Skg
sds8jFkb9lAI/lhzrIbI68B4OIeYK8N1LMELkCq0Ds7H+suVkFlIBWRQrTjxf44X
R5sCJVNQipMcS80Mcgm/tavo13wwnblpWfRYkUGUn0xg034+a3i+YIfx1lpmgjC8
cXXHUNLJg+f/qFhnIc9hzp5QyYweAHCATrDnfb1ka88TCzhTnOz9I5InY997JVYO
3E7axLquhySJqYfUQKPZK1+Ur8hNfKH/QuJhOWUO+GWSdQG1U9wpYtkionIKJTHV
dcWPBBJnwrbabJbL04YTqWM6AI9YCrWXcri0s/4HzPHiDQs8rfBVNAFibCOG92xB
fIazsvtUBYoWp73j42vg5VZM3g5bI/QU0UKaBzf+QEchtTGshsnMjhp03JHVoNKD
nqjzMB2i8LF4Vqy9FhS8mHqNSP4Ktgwsin9MkvGTZbAB8pnub7CHO2Z2aZrCjJjP
/kI13j+D2FAvuL/0OpB+AftsTKqSmSDnRWZAJZfjrJF4fD+KeeON8YYe1GamjtoA
6FErXsOPRqN/N5n0VWOhphJLrTmHvYKu1zZ++3uyns06JcjqvWAhhPsSHfNYbRao
NqYq0i2ZXvoYXNpe006GDb7/1ousreRPQqol0M3hMZtTdUOxuJfZADYXSCIlBaBN
PBIMMtQ6gGeVQufIyUU0TPugohkrQPbdakErgbwqGwr4lw7l55qa8xAZSYSrKV+Q
aPOVmLZabQUXwyrxKluvFYw7O0SqKOzVdLHfBabqN0HKxkRVahb5qp6fm5wlkaCC
MigeKtRWT8EgoKITTq10QFuDYRxqgUt4xhFliy1gBaWm+LIecYoCS4QAvhl/WOKn
Em88Ofn2buSyM/WFpYIrEnvAPpJPC0Im0y5QHmiOqhoeTjllzmaT/T5Q0wIVuf9V
OElzHjWjJ1YwrIq7CCa67AdqIQZnPjU0jlrKFq3LLLgJVVb/9pNuhxc/bAvaU2j4
1duMfIDXv9INDx25Q3KIDonpwwKbGOJOkYC7fsvRGgYJ0Wo5mSwcHDCrch9LgnyI
9vo2T9XTpylKlZHhJxFcUaK2TpJKE74+MWdSzF18eLBjtpmGtkuNM9tdC03n7DES
q8yN9B1PzglzeZCsiDz5I30Xe+PXyeM9X3XVIX38FwiX/ghkjXgfVgMLrWsArlPP
3+5VJSxcNy7NFz9ZUYLFPrU6pzdLdmJU4okaJqMjvwxZQHgEp7hv/9RekQR+6380
Qr5djKyMG/dPZpfELTvLzzNBf2CtGDQX6wrZuxqS4HFv7LKuVGxvIQr/yUeycCbt
l+CoUFdCB8LCD18abViEVsdCAc2XGO7/USraXYEpCwJZs5KXZmp73DI61lbIr9Xd
1RbLCzBCFJMNBvRWbjnhXSTT/vDC2SVSvmIbUb1dM56udL+vC5JjJt/zVH//+6z6
91qAj/ONfLGT8W+0kore6d9SxDnkZcIiCYLlODXpMjsPS5tCafkgDEWXh8wU/5jH
kseUQZ6B/FeGp4AGBVHgxkxDHYO2jLgC+yBPILn2JJOHjU5hBh7nvN2eRlVbmACp
AVfot8+SAZx4jjieGHqwD3uZvP/5DN26gidFl9hNdfMOJ+xaqWEfcoCTvGu6oJ3S
LL/KJJ7jMVLfehUwEi2PzJNaG/JCajaCwdTZ8TZHpBzC3SzLpctHPlRPuc3j+fHU
Wse7u1Sgp/6Y58sadFpJZ0r7xDWPlSpGgQm3fap9lI657RDYQQkvvkXH+B+T668e
Unp9xLqy5bY5j5aNAhuQR5HHTXM/fOHz5hMYAX/xs0kVU4Xb+eRnoBOelCthAG6L
0wXsQJh6vf20eemwtiQerDhZou7Yt3CwjVbnBNn5NhrVi/OezIvSShceuiL3lBvB
D3AlyNIX+iauOPYy/lhRpXE4FWdkn8JoqTt1GGlPfLnwosW9naTd0xaFG0ZCZuzZ
akb59xXpoeIKniDD1XypxegQ95ElFgiu1Ethsruh9yVgxiTotxoLihDUpYcnNUA3
uiKOih1Am62I5WCs401TP4KNIer6Vcm8Q061Bpu4h/HBZw6iXRsaRHApMwBBrHJ4
0up6Sve1bugztRaMQmrI5vv0Q85R+DkUxZcLrQkOL08OmIZjBnRlROwWZW6wOWjm
61WFcZlLQF2hKI4wQYxKhSA4rBGmSyBaayJhUZx60BvbtN4uZeq0hQOaKuCDNfVa
vMDPEXVXhircaLOto7U9io96eLbbjlmq9zsLpsO+IAQ0nYBiPqj1gPpGhKonSA4h
FhytoRsymkIkWxAv0IPZQMu/2FvLVcKUhBgFgRwMcFv59tvS42TU5Z7UVW1+TB2K
HPNMe3IotJl8s/5o/2S+TyJ4lYVXMgOcRLq/EK1o7iAcwhyO0AFOyBVil50W/WzE
t4InWnlGaE7mPYzBNSF+hHFtCwr8rlfpUwIGrfastOg/WMiK89arJTrTaCoh/38r
WSktplae2D6OR6ZLz+oB9XJ37bT3/U06FvANRz/ic/m2tFumpwzxp0QWeOTQeT+o
w7dxYJWBcpN7LXJdeP+x7cIIdTr8+c+0cXYn4hDxmm+MYqHgEtAM+4685W/lEtgs
pnVC3qmeq6iRLRNGZ0BRCuML39inpazhG3bBIxA7UOeEv7Celq2z0o1bfSVjGlVu
KCrSled0u0fhMO/3xGYLctPlOsDH2957Xb4bTITffcnBTGNV88FOJpUbrNBjs1b6
Qt0SyNo2+YKS0q3B/qbY4XDvqZUnwlXctkf4t6/rgz1N793AIqR4v3QgeMMLL62t
KNpFhoRoZZVqCDozl1ULlfCW6vFGiJpOzGcP/irh7zjjUf/qUT+OubWA9oCTdiHW
TAlPxhd4Xi31Ispb0gfCXIqlCJwcv+hf9Ez6PK5Wlto5I8JjDnlu+l8nyXTIapnl
p35JTbfJxbTumkYbsVpLMwT9GPD/sepb28YhmlvcJMzS/zLsOth1RiYfvX3Rh4tk
eFy7Yg0UtnuA5bbYNj2hYsl3tKQjyqf8qBrTZrXlo/UdtU4/ab885MgyDDSXX9Mn
NleJc3UyFXbQPkU7hpz1pa4eAH5maAHYDGfV/+PiTPWdwm7hnIWzxst+iQzC3aO5
OtWGsLwi4tC+qAuxRjzsuATGw5LFcp+NHLPvCdiVSNjHBJn0QJ19DgdjfUATPEW3
DyUsiEFQXJRG/nqXtFXlKZoeerdUYSbKIUYO8E6WIYgIvZtvSuAIawwaExp/4l5Y
2+a8nGUB6GOTvuZUgD8NDXnMmndx/+BJlg97s6IlDzwV32jstcvSI2WUEwJdAybY
6qbWmkncBlBKO1DY0k8LEuzIq7DZcVPoOyWfRNTXIwHCm6aL+Qvo8VqT2mwmSIWK
ygK/jf2wc0AnL46Qnjfm+bBf0JWO0/dspG5mtmT8sZmQCT6OfeckpHXaoNujrc/M
Cw7wmFzUHpGEw2JpsooKwhRYafpXTWsJKvyHNcXCH49lVyd07G7eGOsFIsWeXBcd
U6fkvCVU+3Hv5M9/ShjsOdbEJxn6rMW5CglbiG42Ukgds4bnLItOjY7BgpPklgyj
hcp+PO/zzvxiGPAkDtWUt+muZKxdK2PrLysbPYzSYMbjG80heIZ3qHZewVi6TAQo
fxnPJyIx//F3xTOpF5CktU788cQXw97AgESmLIsvJANRpaYFSfYStMZtK3tNvdQc
N4AxZyCZKYbocwkC/I862s++1vpEIgtVljZ5w2dKR14BtjZQqsS4q9eT9Wt+FvCW
u/gkGQ4VcZmtJgNvOHITvsqBL9BXhC92EDeXXUswl983NuiKgDLPsCF6DHNObCeJ
x+q4D9FZQl+d4nnGuoDEmZBj/eZztCopGfwrWkxPd7vBwDUi+9K9H9KKHgBS+xDf
SSxxQVReZOTILJ4WGU8TNQYuVDb2lVk872mMcTpo6i4crTfioEShNSfUDCyBPDe1
GcDmS4rGd0Kzb9Q7U9HghpWke9ACDx6u5SJvxWxgGwZ3MdUncu2zHKeHtHAGDkns
J+HxbyNmviPl+627vb2rinB9WPAAuUQRNjH+VqB2P8QjZzsvZEwZvBIbqw91pqoA
FNwSUzpb7garuYt6E8t9NfuQw17VlK88ciDoNBW1qfRk+ZeRJrYjMpvuTwi55Ojw
NsLRamkcVVnuXtA3TvqMihkdmRmUZEV71lXjeYkm//ouZf+DE7bUo+b6grIW0xrA
mEn3KGIwDiljpcsvgxcf5lCwp0bDDpZxEBLgWJPmlqcgON0dt33yNSpu7lmupmv+
puoUyXmptU3y4hFFEuc5K3AyiQlQAa+mRRVMm9MH+3bXdVH9LI0x2mfmMov9dHhP
MLY2hxNjLQ4yHZk3OSFhm6UlzwWzwEkhp6OqLkNwXHd8IzhRjTHbjRxxXZi891tr
0ILI2TWO7347xkbb6NeCmEho3vZwE6IURX9/NIn5f7QpwRGxWZpC1WytGRKoh2Ip
oOoEPBs5CtZ/GG0UhwTfI78n5u3ba/fBRZALe8Tk+33tW4EIlQrMgOftXXnYHPPk
RVb+sKP6TrjM1NNJUYNlBfQr71TAnJjukI+qYRaoSJNrVcjhCroBO+IGtWN0/+18
4ToQOs/owVvqfIF/Zk2JZb8WeIQElbcoJcGeqZx/Xwo9yKLwV3EFnbBEHHBtr3Pp
8y9vztsWJ2OLK0gbhKa6pScL2q8gaG4hygHH1VXklFhIwuMpSKKzH1WqB/vA3Ql8
cBZmJERaoTKkmxGrek/OXuX0ez+RCWZVDWAoiWRMpMF64iJlx0kfLf4MA5AH7z0R
MXTr8CqtvXdRR9s0ySNynSrksbplqqv5CpP1r6nH7/V1obfWnrXNhqg9Wm08VzzF
yiFgLbixD+Bjl6Y+xwBTi6VhyK3bOM/2GQ9VUaBnir1OvydnjL/GKpi6iMDQqVuF
Nlj3pZz+PyBGCIS9B9phSPOlaQnYUUEklklTCKD2tCPwWr8uKcv86svX1a+4d7Kd
LWBxf+12xXPVaFrJpb7iUi3muUbRU6GhD/rt1/RVmo/IBowRqgsh/7dsFOdAT9Tc
CGeF1ydp+sBHLbQHbV4QAnEeAilZcU9hmfcOBQNd8M13qOcxwedyQSsOECfMLHrk
race1SF8Z0J8UpZhQInQt7z5rojGM5QLmKKONyfzX/+7Wq9Px70x2ytNrWBgW/ZD
LWSFE7/HlVMYrBMUiUdtqhRYNW25hPf2SA2Oteq43ZkemnDgR/x/7blG4EG882gI
zb62KiysKT/8xbI1pP83g/b0WTRT49RZYuC2BgasBwzjDTAVFwiaAUMclVK64Es0
nqb/bcUu/euEKVwp2YlMkwhSF/oFcb7tcNevi181/LA7NhaQNSLFPzUIPHb7TTpv
zepKQzoruO5MlGwPIDDo4PUsGwM9pCOuZijWtR5BFsb5l9T8yU1kkVVNI2tbdM0U
/DnfPBTmqJfXh5dCTRA9iw8SPMT0xY6Fe+mzEm9ikv3GtdYR9dBuAIfDAKl8AlqX
BRhVYVSDY9R51dGzDcy9WbkNlBEzZFzNqX2n1LI/jREoG5YKBgW/aTYucackZtnV
gHPkm2CNzmpvcghS8SR7P20lZPYJRMfjjT7V8TILDt3uiehWoVu9NyErecKyM7u0
w8CHrLpqNybr09srOZcoM/8jah2md5V38W1OnPcPbQd6atS2N5y5B6wC1A5/kMsL
uHjWLg3Czr10jYqIZDIK43YVB4jnLdc3xV98DiwOx1A1w37Ubm9dHcLeBCeeI3Ym
N/colZKhoU3YjIh7zakU1xGe/dyulM0YUwYQFTzLhTDOwKclzybnMX+wYJFw5JX8
TSLejbztnatNgRCWGv/IVfjzWIynHWDfU1k5T+dGcodvT516nugq77Bx/gmM4ZTW
ES5DnkAcPGqojPjvvkjDAh2UlUNE+MwtosQgXhF0+gglCqiLu9XCPa1V6lbpQ/zR
OkH8IHhCO5VvwYxXfj4gMAWEe+F3ymx7B7cJW6xaRkLStLREbI7HdJkzQ4mLgyzq
AOB0Cs0mjuQTwVG+BO+PxvmL0PvqfM94X085nkIPzTKblKWLideZSdf7E+UsfeFE
llbaJ9KmKJMtjVVncxmCmvORu0cjb1dOZaY3cC8xYIMfpedJ/FptFHQwM1Y4DJD1
lEVjZEQM++m+wUHIve+qJ7K0ERzBwUV6KQzfsLbadPYMBQe/MSki/tmJ8Ynvvi/W
hV+3/bRwKG5znqr8kiA52DrF4+FdLgf+7lxbl1vSiGIKeN+vUnqPDPaxYa0dfXt0
ICiSCIZyEgQAmoXH71MH+m2C/zAEz/5uZl9QERDuIdWpJIMWnoZOvZS9xjLP/tXd
JWNXIG0sYEH/vMhj4SB5zaX/rf4pHAFZyZqV56BpAicTwDLYKMq9XcrxGpYdI2wN
o1lNG2dXfPF9414duFw4yiqjMEaTWUuACjwvlUdF6G4AELIbIgmXWcsJlUANylV2
RQFiM/VXUgbdVs6av0Ma7jHeZShNoLSw+xGUC7ZffmPjKwbjkm3yKMLfXk2Ypb3Y
N07yl0iqW3yQJiUQRtQn2UetCdYRAm1c1jv7YMNjYckV37aOwp/P5CNI1LSpA/vz
i4tR0FXAPdJKHG8JTHPQ09Mzb4EoU3kCs2A14zY5zwElthi1NUEl7eMDwImUGDFj
4XZ2aZFSNmAkHd1o3e4ieJAjlKlLg7mcUfm5+OT1BovpViji75tOgzmg5qBpVjE2
aYCzzYLXnBqMzTtvTw/eUzpuZ6SQWgSDUgHJLLQLVSrb9UZaxlMfxdqoU6UXChOC
clG2BVT4OyCN9pWjVk/hNwiOsL2PxKbQ6LKqSr0UwwLBEWJTLTu32VIsSfITYaik
RZtkFkZZ64+w1NXcxf+/pfrwECzrvdegtf5yiZgzAJyBbBEuWmZ50IJCFohUvIOT
OGVW2pXwzOcY7Nv7wgbBAETKIcYWqwLl+l2HK6v3hbz+LheuNht3oByUH4+2qawn
8ukBG1ntEmquCVzHk0tH+41Lug6GcSCPQEwa8M4Ou1rlpAzX3X0AFMZ4Tlork4D2
ke2iFPxdijJ8NaIqz8icj3JHeE9iOJYpEb7JCJovbu4NsZIOGdseRmF6qExztS6O
OE0O2k3zI8QfX5XVtTs0d1kA06b92grt8CAvDKYNG6dr9XxNbUjJBf3UhWdhvwlT
43S44T1q9TKpqFJkCUfvVH9Wv0Ak4dXiB2hPQwWY94guSivgloXJ1eL91aM8OcK8
QwzZ672RNvSQh6p+sYFXvyvWNnTBPK/C1vgurxj3Bsx70qaXPD5Q23Rb/HYps21C
m/LeAOP1OQFg2S1scBcQ749ZK4YLrQqPFPM/wTFTTGUJa/jIpIIQbxlECZk4CB/D
TFGRT7VfX4meZ3YV4qSW/T/4bMoKnVM66oh9IwCNvfJ9knFCiga17+5/AlOCTWUm
ItDEHRx9htE5mcryIJ4dmK1SX33EDdJ3Br7Ss5ZBiyqxh0gI31B7TcB4gy1SJbYS
aGgL4IqXe5Yie9219yX4QHchtSx9gv6zU+zXdOgWR/kyFuJ1jD/GN1aFCrqDzb3C
Cjw9esXN25SBDH7kYArd0hUk8Ga2a7Xo1UTZa/gwqPtIGhodJZjY3l03ueclm6+i
pCRfaC1awFYwOCjtGuoYyH0Wix5if/eRZPWMBzXze6TjpiH+EvYFJDYcPR43o73C
AsxdmaiHWKjHDDjZhrBhn5KIfkxppx8BIp+9TIMBclH6NvDxYUh/jFOnm+/kK4xi
hs7qGVClgElPdl2XHWZw/ZLxCTy9v+XkFr2OS8Mh9DM7BHAzYVJjjUpvAoLfjiL9
SCcFuNqQVfk/L9HazIxv/TjSHNoyJO2blIyMKO0BvHJfqFpiJ7gCGssSqIQlFJmd
CSWrBAp/sRtz/rWBgB9IMFsi0aLuD70AJFC4nxfPL9QidTpk/Xu9zN1tJMPHrw8i
gpyxt8VdqODDNg6nUepKANhnjm3wO33De4yx04JCoX0jSvyLxXOBFARfUx6IiWyl
XOUkVAWjJz1uZy3S9Wg4/GPx/7K+SBVufpCpilW3QlZmM4TwD9+PZEOJztXa1rOY
yHVzz/tv8RvoCwNIB3t9vFIJcBga4a2ONq0ak3VvEozoouF2f5FFNl8ptWveN9/R
B93L/95xALqDNVjlJcTVqW5MEteVwhya9IqLVYGoefRaZSGhx5QyrdOn2lkbhqEG
sSJrve7Va9TyV35T0R/a+UFbBGzFxpXV9vVS4lOKuHi3/FhtmB70dxI1FjdjJpFT
Q2TySII7Zi+mCicrAMimFoU8ziMP682mPYCWCUesVEFaJFbwA9bDMgbdZc28Z4O+
OJJgaxcOjiGtSXXBxp4ejnx8BCULJlnS8poPExeUfiBtg+mfeYPamXtH4nVelolT
MyNDlJS9Eq2/+OAYsSm0NzxIqgtGk9PXKo43Yeh+D6LeaNPTd7b5sCuh6gTRsSwJ
Rgq1Ytu5AFSeqoRkTkWAZJWVBYLihWuE7uGZ7XWFwiQo17aIR4mC65/IX+EaFlq2
m45NCdgedqKdq2GSIzY0tFOA2Cj5a3u2SL1eJS/lowSv4dZou5pQLjmXW+At1VHK
2RaWpUXEcTvloC3Ls5dVFQo3BPyh0YGSEAdBk9wr9+M6Kg6ZpSRWX91Msr6MoWh8
fALVviwpBPADLzjOWPP4MPDDYizP0ED9MXPpIIU6K5G4qNjvboCjZ38DUsRLdgcd
l1bPhfLrTzyEd6/nNALypScVkMeCtePnIb90PptrBVd/mmYVsGwAoFeXcE3OVgiz
OYQv2FKbmncSc0WPcbOvAVfI9UBGIG6xXDWR66d2mDlHREqqLVsVkp5Vqz0i54wn
DCG+gjPrtNmaiQmToxs8ovL2XPLSm8QcB31UT2n27EPUWUP0+Mb6nwSKSgSHfV7f
gC0xdi2KiG7abi20uCBS5YyxkKCShj7Sa94rjNQHU7GdZbl4Pk/HZ0wSvjb6CsOk
G52x4PhjgJKM5zSEhqej8CdOnd/NErmWjWurLV0/Gh4qE4iCos12oJ9rDTRtkLNO
9TiYecKFFji8tdmtdIvE2cBY+qW1lUISSnTQ6qzi6kczt3wRAj5Sty4/mHTvGtWM
zR14o54ptqsSJtOA5MppQ6AmtDcg+YwY0hSoGObkKFpkl1tcV1TrDd7cBsSY2Sgt
zsbWb1S0Stx2ox64rtNL5CGqHrX6VJO3CTwL9lH0CmXPX1htVqpHFSdnpMp02GqP
h78uax1oW9lagQgY4LdbZFVtAs3MsHMaQ5saug1kcY578IIkCV1kkBp4qAK79JII
xDqYECk/+YpVswfT9SEW4L2/mVWxaBOxN+6y5Mzs4zqDXjavvITAlFAT+XY4x+zW
a0uWVq9IhzAF5qGnNDgLTiQEfX97Kr5rOuXL9QuOm2lMwRBiZdX5A9agDNAADstV
wR6fuqWEPo43MviPOLjj7MKGsVdxCzgh1xTzn2eBVdL8/h1aN93WdnT8x4N4wO5Y
q+0BU/u5K53o3GmUqAkoAprRFXf+lommIKWEyUgxYPVep1+OxdhjMomR4UhNx/Na
Xej6XOzcGknBkjJqHzXlH6AZruaS0XGhRFv5MjIKKkElkq2J0uFt2sKlNjBKqBcj
+m6MOIF2EIFQAw6iYt0G+UIP19HjwPtIi8fANDz5F4KChyu0qAIbz2hl+vdJwFEB
T3LTQxKJ7KEe8+B6LGuK9jMj3aO750rWuDsR6H+l5hsF4EdRkeX4aKVxU9a66+Iu
9zw8oZxvmMMPo8rxo7THK0fTgo73BGbDA3iMbEPu0VLVaVsDgx6mCZwxDHmaO5/c
tFaQt1uCA3oiIyxkhgY8FjrkMPDQoJY+3ETIt48IT+AKhJVDSJIxE3Nwuk5wkDGi
70a4i9lntLwKTbXcZzJCcDmpeNG9ja38zXdw+JG0+B+0+4SmuynPQlBtLEFDLXBo
RcRuJgbsFank59ShG8LMsfTLhqs1e7J7nXq8QrrfDrf8NTbWrc8PjLYXHU9IvOuw
99WbtQKBP6JUjW/y1INe2DyZIPV0sn6gueH0D7VIicZtqazHJ+Z9l8iSINrIBMGy
8Z/tWiTMhKVkGhqVW7D7W63r3jzBHuFivxyoTWPt7dce9SFoqtZYQpo41DnzXvM4
gaaHtTIvpfrEpfkdUEcUtNJvcLMrXj/ajIjToS8POl2aTsAq2B1vI+nM8dbbfhz1
KlKsl1jkpXGDZ4UyNUqY/NAIxcMlxg94xjQcPRbjuydePrQgmA67WfSY1PL85trP
Et+NBgvJjerWgzvIjaacRBlYoIGmCV8osl7peeopryL8RecDVvkzdR7rnPMdkhEl
Tb6RDoWDJJlI12gR8lcfmHE/sULZ+r5kg7vvqgpnlpiBpnyjyyZ76VjvIQXqm5PH
6NKCRq1FztI9miutIkcPVU9XUyPpDvs0KdW/w/FKeuDW8xypeomTpefDhfa6l1cQ
54mgSviVu1N+zTJVKQJfoPs+O0raHdZKkVWaXhq55l/TRN/lIFQTWPeYIdOQg5I7
tDXzT7sSxRTMymNs9vkvAAzqg6bqUDk5ad1PH+2T6h0PdNg/me7Fc8OORW1kWlqJ
ezm163afHD5r1mBT6PkOV9mwP7JRaOFHpHhKRpLLJAMuLOv1g+NWfhsoQPUBOSN0
JWSxbR+ZXS5zn7RGAhaCb+0cDVK5B6iRlv6P9LpK/eVu+R0/NAd3eujxE7ZxhF4B
MrWV4sWrOR/a4+elk7ZI9Cx2PWLT4ONVXZdTSl77rIopnPTYup36K0M1ZO0Tyzev
jpBnGy0DTRHNkr5OF0eRksvvg1w9+cV5Pa/EJemaHuYJ/bakAv+SqicpW5nVk9Vk
mbfJW/zmC5RYPYhKZUdwrMHz9wVZq2Sy0ffmnk6JgqKi6OHdnxNazNAmaDv8eWgT
T6IkvqLzukiEfUPQSweVSdQOjc8vNRVpC5hHofo/vVEs8/giQDJqlW8yWRvTl9o3
DbRnCFEB4IFaarjXA8+Q/A+gJfEA96/so+4R4uuEbsszaCq4vTyZTZtjzT9Jqvfk
CIjrVs7mpxJBDe/1DmHDH3S1zo+Xz160msA5pNtRqKYE6hEe7cMVbnDr8aS6nX4p
xKqRCBNM3zh4fpxATEDjTlx2DYlgRwZcehHxIyKDcX993+C2HBWui0iV/esrQTOU
QDUn684W0JYXf+O7qynCkM1yPSBCa/mqYTahm1xkP+lVSWczgsUJvIpczlwzKei4
1UrVG2QEm7RfxghXaaki/PiUz456QVuoJoETMYtIsjF5oyr3DUimshgsQcOS+cc0
VA4UeMgt+AZcV/yJiXjbqfSEmQsqoJBJ8G3W0MbDpDIGt1vdb482VOrWfd7SUBHm
F6GI+xJwCawnGoIicU9lp9IZiam3K48uSDpRSskExlN4M5CHW3crARzRuZcDeLo2
wxviOBdT9Et+NZob4b/fD4EdfKfSrvgpEAJtF1TsYVpLW5XSG9bnO94o3m8QV6x9
bn6kaWAjzAQZMz2W5+MLk2ChUhcb80CYc/GwhYfNwmiLaeNcEmsHG1NvmcINOBXx
VtLvYjCP7mIBrocLoDv+JUzWLojgTMyHWwFzDw8wHoKxaKt6sX/qo3pi999QBOo7
cCUlILv3LAah70FXPGM29vVFBB4zqU41ZuziITOTzjO80kx63FmninqrAV/PA12l
8JA9l4abk/4VuQROzuvoEvU2SumfGrk0JWPEVGIay8w9wHWq3LuAlvIy4Wl4dT8y
fF7GjNtz7ssHdrV1FG8Ihc4TUSbyNSmaODLoRkThfnpYPg5BHHxE3CcB4lx0GDR9
M+4DBUf8G/AQEYzU5InGpviFnb0sasBHJebdjZHJliaUfYphBTeTdynD8HuZuzN5
nitFPHMh8i33fJCNBlpPTD/RjZ+lVZiq1AkNjqsRl4vww7DOmMKNJz1wEY20kncw
tEUUzs/67nzquUYSuVekoM7WJB4C8QKfHY1lqfaRvs8zHGFh7b6vytW7aC4/SRwp
oSEice94lpIvdL4JhivwraucwmDCF22SDoAhGi96Eq5mJodQ/iCnUVnwtuApf6BC
kh4LJg35ZzqhcJm7CdFKbr97ZWW0YmmdqC3w+4HOCxrdbtGDlKEijbjxlaoRH6IZ
je87meliPLCuQbAqyZClk5u+OYuhHXfWeqdBdZpzwbd+6UVMjNXFJbW1hd8WgfxI
ZZv9PyK10v2I4plG45dYrf/mUdl/yifuvk1Azn8jxltman0dIsAWw9Bh3oIuZfeC
8BV2lqEvtw48v+xF6/2320gnuGHN1EByJJk5k8Jw2iB8laQ8TQ8qdOhSFRhC7YOB
m+iV2Z+cFbLGCB+8LRfTnzKAsrGhfAjbsti1/eLDBXMNNFzPByhppjmyVxzH/RVb
ORqSxwzoy1rP2jvAVzPPAi3BPs3e0+ykBgWyAjfcWkI+aUbZb3f8bmtjO1n9eCky
UIQiKkVCWsU/mJP/VwhQwg0pgNyUKHjA/XL+buhb/eoI5RVMyM3npgpmIB0FM7uA
hA34h7j0lzDYC3Dn4u22ELiOoAIoBCz56otJYYeAK5MWM2C5BruMrM3YXvEwpFLk
wLX7HO3m7TDR1fyOr8t7SCjHKAm6sDgOLEfFxbQp+UygorUtz0cLdcZIxStUy3CC
AigFl0A/cfMZOOd/W8mFUXi3vhiTRgPAaGT1fLoeiiVkhyjV2EY6m9XT2Cw8EhNk
OT8aEq17b/QrjiwrIeUJQurI271hKEO2Y9Y8I2Q6YzIJWovpEiGWXbsNk/cGDMIx
e5J6zi4gGRITimy1E0Xr5uraO3UY24nmQzEbf5+5puEyjr3OyUrjDI+Bra2iUdRp
56Vu7U4tapoSadOyZ3NnQwm6Fm78mE6hrD3KPw+OsV7Z74a6dDn5FUWN+DUV34L7
MbtcQ5FGUoWxXx/2y0Z7wMC4X3sZgVd4zF7QZtuA5jlo8Pcpgq90egGQmRjr4wfa
GTeXr3rY3XjpK0z4J0tx95ujwIxv2RASl9EAichK9QoQc7jZ9vlGPWxLgfjnRTx2
1hPedR9NEdvUozniKRNayfADWnuKelk27Q86tpgv/kv73k6r33286pi+9bqt/vi4
tDQSxRsH17BkbrIdRV6cTj1b0JpSV6b3wQzbuqvVQOU/laJks7XRDow+1QWPrlH6
KWgl0CBIBxjfpRejq1XvRFj9ldEUZVDrD8zg99jFQXVwMflJ7t3ZsGTqklqYjYz4
OAoeV+IDmi0hRH4OsdfYmr+itiyfJoz7DB7+4R+Q8DkP58zD+psQsYFqoZpQSStQ
sk6zoNjFSFr4gvgtf1OmUZTMROYaI9yv5MxLYqRhOxN5t5VoratjoYKiaTqKWMiA
vMQ94XmwANqFzJ3jyKqGNlBzqaQQbPGYyGpCHSnNS4o37fhpDQW+AQCcjITlPhlx
fu9BROixxf8pf7ymdTqQg6dPC+NsY2NIegVkYi1hadVc0OEMg4PyuKtl/Nb+MJcL
gCwnN+8dsOh4LP70a3+/7HhZ9W8rxtBVA/lR4qA7gbuuzTNEaODY5UY356AaBwcf
Cuk0CLJXt/GJuDwgj67jV2d2LTwKQlG4symjfI8LcbkKYhB+JZWqyO0IFaF4l+h6
eoHHLojL/soZxMcOBzOG719l8VF7d7JBVQiy00uNJz5t9WR49L1RMfW1LQe48Ai+
R5WGCUO55lJ3M7OLBOazyYpRINuRSixTQxn6X2QbJ7IbJCDy3CpjgXh7iGY8pFze
xgxB+Knpyyh8CnuS3aIMHF+gVfZcaP6AklaMiEWK4D/felArTMBHjq1Hy0WQ4idB
IVm2m5QhfDTqlQ3zXe2wSsVefRqkC6TKx+2Tv2yzHXIAS5T51Wa41mbM5RJfrU9U
ZVOy9YTv/SOQoLbIJWreVbTXmAGn7XdYJ9MNq9FQiz9glRJnekr0ZzcfiQeqR74I
y6jNRMwGHGAmysiNyrwLqteLc2TQhMmKF9uS2MZbzQyjZ8xphv9slXtAFOCBTrnd
f2qL2sH3e/R4WTEfqTMeeEEiKw1jlOdSsK/qUlIikbWBSzc0ffbDtQ1SVchVWFVm
CUsgqi8x0rnELNtLK+fQl+gXjHXteeAzLVNoiYtrT37TgUE+aska7pe68SmQvAmD
6VLnWod3UrMb/25dvFHlj4OGcI0nd4GERdvTToJCRP6/8ciEb0HXx8wlc0TMu449
wWgL0UQBMMsj9XVUxIGNhQY77GiXpRladiW0rLqs0nM2UBFhZmcR/BZV+VDpDnYT
zgmn6vUR1HBVx6o+Rx5L0Q0NhsCej2L1uDfVqf+DmQJkTf9SwGU2YuvqK133C+2P
L12b8jSMKvjaiowXAP1cAe8G2KJYD2NAVkIG4SccmtddizGon75Em/Fo0qvPJltO
7X/Wnsecy36tsk48QKEYfLN5cHMYTHpu+IGQLTqYKSvhO2OQ/XSIYcwCshc1fitw
71qS+yBFwz0KfjFsfGeEbl6BLsuG1lQIWcejpGIxYqALOOEcLtNSs8xjYhfZ+eAL
9JX58IvVbk4b2sxnElukUyHM8nxh+cL0oPbjeNZSo18YBo8izStYfi3EZgYvfwjK
/3NtcF4i8VePRi4qHmrazLcAcN9aAN/iPXkMYKLl3HfhqUzo5O9liZxAfb8HQ+bv
gO6y6BLEDwU+M0qYl67QDUsTY4nDEuDYuVO20aGndCCIGK9uL0WgZNAqRIBFN8jT
+8nMtXJEerxcvRi1tiSlvem/VSFnxpEGzdQkI22tN5jXohIsMeWUILEgbT2CThzv
5phtbONtFmMGiRx/9R59UhWXI9g3J7Xt4eFix3xxSlDeaMnHZAJmLc3EI922o9iP
4zRNt0UkUoj4K0alJbAoJsa155EJwLwqHRsAgtYnYXRs7BfW4UkDkQ0LU+KKkLNC
rzooIofCiyprYxewML2WzGkQXz/J9tbbMVeWBECuBXMHAEjN08y4UhhBmhBM8mdf
YrzV451ymGXMMU3o6hlKTGmMvdHH95/+3mzn22SdeqxohzUotuE2W/v7u6Ogz2jo
Mm0ezcvvKaLNPPEE/hvYO5uh9WPyR764AGEKhPXWcjMBP3lsxaJ96adPAob+Ik/g
L2phd6JG1fhZ7zFyEkcszAY56QD1Mz6OvEbEjmfqViWo8unUpiBK5G7QNOt8XeK0
mgp69lLBgSghAGLFZY6pmsnH/LdT6MPhcjkR4RV7VtuFGpBZFlnc96yi4PpT/0w1
gqYiVv9s2hxkDlUQz468C/fyhDqMfH0REvdx2BJROXw8Nk38qi7dFAAzAys4KkUI
xWWV/VKRzi6tqlWP44ML0/7HLx5sl+gKAC+LCzgX4Nd9fXmca8FBgLkqIRF/3G+r
srSvaUEtV16XI6lH3RxpoPV39jCBbyIMqJnSTKtnZCl7QLLktE9hLBEmUU+bJhEU
y7fEKpqsdUZbQOHM4xLOuQMGe5d+xKmYVRoo+APgljXAeY590YuCZXmT86KiJWpd
KB4R1tyXSd8YdvQPJZAaeqJVAE2gGtRyQwa4d9NFnc/AdrrmAAmx2y8G/lCTf7K0
6BS2ZP3NGcCrQjhSo9C/cy6eIy5JAvpmSPud2pho2sLas4ezPKMYzS7OJHG1VOlp
aI8gnYTNp/YyKvPVP/TjRL/ZfwhdQNOaZKXKI7VcMlkvwPPUkzNF+Ku6TOtNtEf/
DgQRTJQ8jftt/5R8e7EjwvlQdFZ4Oi4u656dlyiUFEVCqC5OcZ4cWmag5lZaIDHf
d9xR97Vq1NPCT9uoBykqyuAiJsUe3ANVXw1IOystvrCe1T0A4rv0j7BPNlpWWADz
rLpSlIiJfx0HMPH6oZPr0JcHuhD86gkz4XKUg3d/oz5G02TT8hz+Sk3EGrKdAzJz
MfAfbUYrWmB+esWNMR6A6H+VIpEXk97wiNnS5bOJY7xmRIa7ayV+VmbeZbaGcvlw
1dOSXRR8QTX30OArHHas3hqq0IVkFoPDODnluc14sQtBqEzQiNJi1FXaJ/C8BSRg
lTZTQqryqE5tEUjAxnyHAcpW3ff7SapvsmTHEFnRzY1+h8Ai5hjUTajAh74NxA3S
inEEniM9aEIsFCJiEJfa0NC/lVkKeQxAXqC2yxPNUaFj+d73niqEGnSN8Pp/DMPH
Vd9GxSU1GMfWZbjnDxR9Kibeevo0k8ita5y6sauOqFbMZvYE2tEzgwEvnf2vB8le
/gw+DDti8EFsvZNCpROCjbWHlsk+1GvQXCwcfSum8LUzOvdbpHoVBAbFT1RiQGuG
k1RKOeR1KBXXkfv8Sb/QOA6xsMWxpI9RVOT1nAm1twwT2d401vF+LNIYN7xNer73
ZYNrkCVKkwcGA0BFj2eLrkPhJcDaxHYong5AtcXXcrlVFyz05NeJNjP/mlz9JISg
XubLKLkwl7PhE/D3FVMO8PEyQfSHsczECw94UCV489TZI8gBzCJs4Fx8hgII3dRK
fpES7VNUy4c0/zOzOuPSmMrgOgxJSC2HnII106TnbIqHm7x4u0e0GwtY49xjgAPI
bDeO99a1qwgEVcl6VOdpgIvTWJRG0qWhdMJnFPTJnAQbaTpsOVV4FLphRVkQvRuw
WlURnFdQtYbGU7eLxUPuoUvj6RdRg9VVTHgG65z0TXxgS6CD09dLvEUfPjVEXfhi
7kDIojamZeTIgUZ9dwxAhULKBcF3pd6Y1d3hzxvL1sG/XmEX+eukO1kFm80wjWuu
TQ0d+xR4na9u61WiZDR8v1Ecm8xwMUx+9aSfaOlil6y2WGmKyVIJW/ObFTKMLvJT
llUARoYB3B2ILounjLjchOOsYM4FsGBu3uFq5oy/bvZT4RD+MFy0j6hyeBa7KuyG
W+CAmGDomTy+oaVmc8aiHR9tSnDqn9ffWNxLqy2EYnDfoGUS9Us+HHVaKoMXJvMf
Eq6uT4Q2n+NkukOs4vfisY5wmsm2tUTF3fetYOcQhbfBGxG/4GpmHCdBYZPIZdNY
ngJje+wRyMpqe7ewpTmSNB5K9/ZqJs8mLLiSOqS2fImLvtjKgtFxheaSeqaGN7MI
mhT+mkwN6tyolUqFo17It3O/KhCje4EExFoGEBJ/5FifHpuKyZWDWjlIOy2mozwO
ZT6AUkrQqN+81YcClLgptB85v3cJMjf2M5fFfVIzsArZQMoU2grxbpWF+d34kGRI
M9+/3QIAC0iG3Axby3RJOOjjIpPMp5SvxMZ2HjpH1i1Kvlu97zim46g/4VTxF2G+
C818r3vlDusZd9uR7SShbit7Agiy54k2d33eQYcqJ5fsiYvynLEq4l5Mq6SAP3Cn
GO/+5Rau4/YchSyp+ILX2t1dYi7k4Jd9jWPpKRD/fCjunrqPR/Nrf+Zj1+Zp6MBw
9Bxe6F8/pXFd1zITPY3SrVx2Z/9XIUoSU3t9YncdDWn4wpHE41TEywdCu1onY6bW
N0x0soDTl4pl+9yEpMrWet7rzSOadki5gULlcu7z2eea2KoXF2hRcnos+EgzkXoM
8LxEbhK1UTWbmlQEMoG0D5V1kLfomni5nb82elDavETkb2flXmh6aZRcpjBLfRza
xOQtzUyT2bDxWcvNQQCKaTe4Viddvz/sv/HLoX8On1Gn3SStB8hrs/b9bsG6cq+P
QJU641d/4KGh2ECKXJb9+lT2U5FbZFwQoDzUV4P9PmnFZ/rEOrCI+j93y2EBCWBI
BRKz3LBI/jDuWnfHREqcvxFJBh5nZZC4SSGiOhYtgOe22t0Af41lomrawnyphOIh
YhdE2syGl2+Y73qGFqRoN+P2ffWpIsv9pfIccurSXSBA55NkaLROW5hqdqMaHp7/
IraamOaKHNzps7he2SDdwYY/PRKpQYCHEWEVfir5ANjUUxebnUykV+zloPtkbBBj
QuKmN1bSRX+fC0F55R6beU5AIASRC9JJUcTpPpGM/PWquqTX1EHtThwlFl1IYwTs
VIpsxGw9YoPFCrETa+ccQ5fVA7qfb2ehyzEXYR1d25YsumQ4lHC+VoYliHVZNqU9
0mevnBdFBJkc1aj3FNgVm9FZxw/Xg0NNRgNU8rMoL7ms6TyeRcjIdWiT+XIWEStx
B+3GHbaj4ryECIsuirYGY4+mwXUv+0rid1vSFR6UYTYpLlQf9MBK8IXrCII77K62
sBfTIdQtEy66iGqHXzu5/9+FTc6ZRDPUmCBgbe3o0XRT11RgMxaU+Fr6oMIr89oS
hkRWMQ56Wfgk5/V2isRzEvS0o9KUSQLMc79U8iTmScztI4TYvqTnKdEl2W9mROM1
BfpzJdXP8ZJs0mQWVdyhvyybJZ6MgJu8JbGs19GXH9E6GSvJPk3g/IGkXMNTfnU5
iNhCjKlCGN17h0YUXr4Y1Knaw8Yav0djgLFI/L4mk+fQty6VvC626LgRNypKd2zx
OHznoHjVYgn28kyP2Mlj3XJEKjf99pd8NkvUEvddpQh1tRJGqqemLLMPBSJzzBl6
StZwYHBbJtC1UawDu9BnCBUitKol58LUCarB3oiDRThhKR/aCD3EedLehcRdjrol
GVRRcP/FKcKLBJ+qu/KFFbnn9Y3C0SwXBStIqWJpf9Wp1nrcr6pvMMZm/AhVTgoq
H4fna/D0+u+EMIEOxn5lV1kONKy3Mwr9qa+/Dw9r6F99n3pTvUpcx7p+LhVaWC2V
/xIPoB6NfGLQrc8lPXxDj5YhAsAHtVHChjJraTqhxUbCOiWuk4nzS2pqeTgOLMIc
1eKGrsc8/3z16tNlVXbhEgYM1P3rd5pzN6gNj8EE1L3MgGjSdd1KztuPoIm01GCi
9usoCW/pII0p9wGJaU2wmhPhWNMlcyTKCbvGl0qP/Q6oy7Gx5GF8653j4GROzePk
+627NJ2cznx77H7R3AWQwFeScgbe+6TECVkr9KiHvoTn2LoqG1bznkb3rkyNA2Dv
/URlYJmKnXUqJXjR7vtgDlX5mtOU4sv72Pep26pw2WNCpkZFFY+617tLmEZjnLmg
RJrZIYhkFR/rQ6D0e+Wh1y+YgRxvLyf3dcwnvSgytdrgz2fjQGZDDKyy4xSxU7CB
iJy/SXTZZPaPgJrhuEPFfZp+cqxHIaoH9itwPrmhr7kdht7I92qNEYfg3G4TsziY
jrUhBu4lNaXVO4JV86iW2cHGklL//1XGX+eT6warUMoEHmTHT0rteOGCgUanGB0Y
OYjJUkssiXvUgdAl5NSJvV1d5F0I7UVnNs+VUWL/w+fylaykQKjd8veA25a+FZ3U
libYQxGdd1YxdkDN9B/FfrIDW6V1wz92bpVOG6yefTglFNMbW179raKHc8T4HbA3
2FuqEzeXeRmFhp1T1QlK6TCZOs7wVEQoeOy392Z7HlyElRJi6ozAgtr8gtSuW17F
UGB3iRZuOSZWFKoH+tL7aXmVMnlt9U8g9J+LRljZ9y+xmZqupBkmr4Zjw4/cd3ZH
ngZPV/RVnSEzMwls6D7w7lW9/WPSG7FmvGFmVPktSGBdIoHkdbiUXYD7ytfnjbfA
zMqznXmIYEUfpYZotNnZicYqYqdl3/IIpBVB6+RRm4aRG3USYblQRzHJFoBpzOcA
P1ivu3IKYPscSd+TDeiszY9SSgozEOKMT1OVvsYkOI9G04VG/nH0W0wnJV24iBa3
6F4KxgbeGWmRWxPFjQKP7VWYxlN7sZ87NF5/ZCxhZX6p/cKmRR8V1/G6sqYCy7RC
fTKgk2MBn5LyndpNdg2f1RDoqwYiFZiod5v5x0v0DDwMbwwO2bLmKl01sUo55hYa
Dz7x0JbOMssrf9SRiO72a3E2CukMAcNKhXfEwLUHwkCe/51nSpEkkd1WaeJx9axY
HpZZva81giUPhnl/Hi0orCZD+qco+L5G4lQ4TLqOUr7DM+ZWXpTb9VNdqZzq6DU5
HywXU8t2Dhx2uSD8Po/7u4wKceC5dK/mekACsfs2y3A3KlZcU9xmXvZWg5x2lEqD
8hDcJw0Tnm7ztmGVB0objwoXRmNPrb7hJyg0hvF66Xd8gKKj7JX1CzlNmUe8vK5l
UBKcGIsKHVCt87xbeYvHlTptG0nO+IGHTlB7AfsxG47JEJUDRnsdEaQ4DzF0Zh5j
su29IEiKpvr7fKIerPg5OKI/GQsgI1VFwaS++MDteYCvvVaC9fQARKoKuWza9iVZ
6c2cO5hmkC7uSSkEwE9Ia7Fas3XvLMzr46r0Feuc29KIPxQHzx5qa8/O9M69PaoI
dD9LhrRdyGRHEimlYfOZriK2VhGKnCu/uET3GNGAcl97JFFMh7sPHJwd/BpjZ+PT
boOzOwhyLcxmJQcs91dLp5CPTjkIsvF6NA96vjEWlKW5wlaY90qaeiTRKbSefBt+
EuBe+t3ooKaeGWgnx1Yj9CCgVctGwNaMjL9taxs/Fl7nAHuYONHC1y59M7It0Mey
xmXkicVwkUO9y0oS2z5hahu0P6MsLhFyXONu6DLc+ozOHeodfMjMbHfN1uIUQxdk
XysGUzwSFicQTDo3wxHSlz+idwJ+DM/pP/fyC8zVAHDYEwAZv24EnnaPu8n7GPCV
KCZSPG1mUs2u21Ej1m9D9a7VUNPHfFveeSOR/d+UPTyk7pUHjyTige1b3pH9bLbR
79SAZ4bDhnHr+yGrpLSq1hkr/jPpszQJp162xqiyVzeRSA3eiYRROr7qpu4ypPWK
pQTUOKP+7j23D3iRSH0QNiFEl1EsKBFUU8SQEy1w6mLy3FD5BNB/zRvgDCbbV8xQ
ZqV298/dNlCt5cvUBDX1ATqXvQntLLJCwZe2273gxQ0ADeowqezZrz6ZZataiakY
BxpgP1UcAETbJhFAP0SVNhtxBgn88eSL3gfBSP96P+x8dch7bfcabgm1j5gIM7dx
fn7AXp3xMBOesjUVwH0tAzZHbpzOYCmvkfbZ0Ro58nXEv5qald+tr+3QP+JwsdH7
kFFxI0blejqp7XLOg5PCTwV1iTEs93QU+UYVy7+3ACW78Ro7ZPc2jN3j4T5Fjbb3
eH1GUq0bxBc4Lxt+5VQA6y8nZDnYo4KSIQAJb9Qu5Ztba2jIoxnmG0sDJjT957lp
Wemnes9ldSRFvSwheXN1ip1b1CRrSyjljTKaD+tKJ0wUg1aCxiMMa0E0yybxQ/zn
of6zyPYYs5mIYeXaCxgtGJ+vXkASU4kq6k5EGSY7U6bccIvIJHZJwJwowTZ80QpM
8zYYZ94W12Iv1Ls/AqxE01Nh8/v6ONFyFEsUvP69NdapYS1OuvwXFUpWmEtwIQvE
IF3p9vxRYGKMHWvkNPiUejuFEA27xipdqKxtBmYtgH4qr/sphGtY5vH9Znv5hTw/
wTgIblDUTzkqmv98IcvNf0Zwd71848ByXjJ5JggvNVnsamboymTzqxdHgmlKOsiZ
thlYtxngzgTGj4fg8PwSiHN4tUZF8a6NeKinCY1aUJ5PbTTiotJvzhbZ8Ah1fVuC
FjgeyfWuM+0POupDTRst2KJ3EDW6pMY6mnCJQixCLBt+ekFDRzAkYVmgMIpwSujJ
4yo49rlxZLtLGQ6rmYSDbHF/QviWP6WJkUooPIFI2Sj4p709b/EdXrLPyWL02d2T
RsVRaqdpSXEIsYpJWur8MsEpf+uxylZV1jLPGnIuQY1WiaFVpmPiATZjp5D9G/6F
Dk9EyVamMsnGOBBxbRZ139GJD7Zao7EyfDvlcJJ79Meej3x/5AjP4KZ0v3pTKmzD
1baZGilNtN+VMGucEC/f3E1xIfaWJ/rcd2d/TWDDiFZcuXg3xflo/6WYsmAvPXsY
moI7mY2FSgQnAM5oiQjE6rUO+crR0INGWXgichJXCb4cpqV01a5qX+09oZwvJAWl
auOSMPDFI2u3eXk9Kigj6HSPKVSb+bpC1HeN7gONkXjfNeY+CgWD4IxXlqY2Y4E5
IvsfbTCCUlqncXB7l7SC6Rv9ZX4VVbsxc7uj1NrbflhC9o03Hmol3f1BPS3GSbSF
a+db04CHl5l7Vc9vwrIbesgw3JSvIUVR66xxdjds6c0Rbjy3OvcieogaskKXqKj7
5n9aVULKC+pBt6/+sgeQcrq+FGoeNZaprTm20bkYnUEy4Undwe3qpB8aKjYH0IuZ
xwmrcHPMEckZlfl/yFpSMEsAWqFFORRx9uVJgH9R+Q5H//S0BqGzqAI/GCdKuk7F
LOOUA+YP/RJB6WciK9a6s9rTBmaTn7EbvitwcF2/ZhMn0+66+hrX3qMHzfucY/Nw
mAgZOn6DViMnAWSR61GjZwsllAVLyeXqwqdWkbddtOnBQ21xRtIkcDubRKGVZZS4
fvSn+c30rxlRF0ogQIvgptPBirA7hcU717NJrpiTdGqIX8wjoHBj5yX2OvtrQcjQ
Q8iSE1+tHZYJVRn9dF63gLXPfpY1kyjOI4Bi2fgKpV02G0+TpG87mOShdN1CHvuJ
dZsRmWJ+5P+zrs14MbSUT6KjMsxwajut67+V+8LISc6UW6dRx3Em8kciXQxcBJ/Q
Ra1zkG7q7VaP1WgRN93yPXu6hvGVnVaWUs3zTXGAD+dP+1fMfwLA604rUPW9QiCD
ztJErBDcfzbAHN5mhE5urF3pCl3RBGZFpWQ/GDiE3YZ6w1ycQQ9YsNyHfL2ysABK
/WiQqjK4ep63Tr5EL2+t81bnFC6PXp6y+pTK/2chtqBwrlpxq6SGqWl79XAiJDHr
3wwpnZfSY87DpQQull5wleYlRtnY4O+HkBCTAa292VGs1BqB3ORNqdJU9ohsdq5O
rp6i+1actKxIDOfmfgKQAM09yzjNO31DTNZeJNBcXaZDazSFqgBuoYcWCBVD/+2e
wN9js42ul0wH8/xcaC8XXN1Jcgym++VLKi+H69sKxsdoMRJNOJCSo1xRPq4xsLEG
/ERrNity0uYTb5bObxG8WUyx9/wifCOQAOUX3T6Z/9lnYonSKHchNzirGu60lNba
dSyWTKjK86NF8QW39qo9yXKloM3gtbmerNnzbDMR0SsJYRdRs1lOhcU2jp0h7d84
v/oQNDyvQsUommftVSvo8tYcc+Xv3wVL3H2Pymd1GCMJ8nZAM8A07GgpgYqAibDn
givLkB9Icb6IGnUZ7ToP1YPa8ezibELQMz0UbtMZgylgT3PmYq5RQZz0wWBvdobd
y7y0SeXEL2peJ7yuha+1NWEyL9Yv9KpsKqrAzI5G6rwt7Zsd7/qrhhmlC5sRWQaF
I5iDoYQP6BqwJTQnc3Ypl5VQNIUGDMHYTPsJtfqsBt1C2txtybAUAtQEL+hJW9V1
zZJ3I1H2nQ/B+zmFR45vuhRW/sm1oQcMIjYpC+MMcMBhgyn695G+aDIhBnRkheU0
ViOYd/yvAYqQbE162GuH7xRxHma1Az5DGiqVzpGhB4wxCj4rHVeVA9GrFsckQn2m
jyPvL72dJrEjY7LsW5UX+k6Lqgq8lY4783UGTIoEj2Op3eanVutQ9ROfWSYoU/Ju
1wQ/fQcnNNn4i7ddcOepSR2RlG5AT86aosbklgxI4Qv4ymCUYSYXhXescWCLYNTu
TcqdZZEcU5EJac7wg+yACocqQ2R4GenyUDI3DFBqeBEbEn3HM0UxmR9NE540FWwB
wi+fU2SNlGUzTdPJtdeUrn2y8yXgQUnJivPdkToqYudqYCpgsvSM67qFh1oDzEkS
kiXlFSzSpIG3C2br6WBlxUXCtQFNJgOv36U3ktsCwje3KDDt7Z2uAIFQQmF+o2rr
QMZHcqwnJshoLlo/zR5j/bzlG3AvJQfnte2l9JhrE69xe/KebV/foIIUj/tklRJw
iahhqH1QoBVVfs/AWyi9ObxHO3thieF8jrkJ/SnGf1em4cm808DNFcDJTDVtEJN4
H0HyMK0YAUvGPAHf4WHnay9FaKkACRSHnE2rqJB2/JUOiGLN8hXkBcEcx1jJJbby
ECNZWjU0kX6cUkne9yvgFpwJeHxQdl/EIXPZbPMKEC7Rc3FWG7JvPee54yhjkAG2
lMd2XFbyFA8y8z4u0PltHDkBvmqRDyD2itEzSbwB6mHlApg8v+fGkYyZ562Q/eie
cuOuwwwaGYIwS+j7zjopey9yeTWPOgUxmWcZgwOyWHrQwK0Vwpo6IfZhtHw3Bmne
fl2adRZQnYduBCIHxs0hh4TSyqoIwuLtzxeNyuyB//7scKSD59bFpw1o5ehDKSch
iYCXpx5jbcHqimf63RPva5nuKLqJmbbVbcxT9PvUXAwxoPobW/NCuchqNvkLOC6g
9t2/+mUzkexPiF5jPwanV9StFWE53WAOjUy2Kra/ZNEgjdMtPloW0ShCOL54gkg2
PIqj2sZ/QBlipCQ1LNMIXwJh61fy7heo9KewKYetgAGSfr18q+elcSOECa195VMD
G2549PxGvKuPH/VwKOfdZzEcldbd+ZHk3RqQf7gfsz9MM/sJSzfgRjT7kdjanSzm
JkNS8O0fsHlKWPtRxGebfJtY8aP4TwPduXQXf7vElEu6ALlyu5Bec20CbtGkrSRI
NxbE5J6f0BuVCiJnP7q638+M3Rq5po763GIW7E4+XnykRDyRwFDtjUYGy0dXwrRZ
PGE+4g4+9gisjUPgo+iv8preIEwLefM8hAhB5w7XbXu65hJbKZbsMRmnwxYzT97c
xww6YqGuKpClepjIaB1yFlHger5FCohQGsmmPL9PT84OOFKMPbjP8SCXGKVwicz5
2SA3E3U+mV8WmeT/pYRy6OBVWf0hONAxmBq9FQN+JJKYayO+IF+SDMVzl4aF14oM
bWaFIeY7SfvwP3RuB4X3bWSk2fHvpBx91jMlcmqqOBolC7RNpNBI2WJS24pjQml7
GRaKt4tOgBfD7ja8qpWKm2M6JdnaVWusDZgvPP3Z4mYJGM3JQWIPy0U+yJOMO/UX
uGdbdI3vfol18cmwkLFqDIqpc7EhrdQX7kb9JBpVIZcB5YIfko9muVjTh0UAcg1k
s3SrcE3ioaUzLCqOVnkzHli6Vzv4SEt9u0pqjh3aHppVBOy/NIoTUV+Hq5P+QrTE
0O2U4yuiJSF4zjal6I3xbsdcBto6B3fnBP5MSCLKhTcjwPS2koJ9IvF8jd7x71Pc
Zu8CMKhM8jXxHBe8cmeK5APl2UHXvAvMxW1y/fnXME3l9Y5KzXUMmYFR94ovoGzR
K/g2BVe572VFVGr9cHGlU1ISTfIdTs9cdDNbcOPhDwejk8pllOOpIzP43kWAbf8E
TcYgSRrjy58CMkEeCCegNqNvH0IlFJD6ErTf0RcWkLq0Q/mb/CjrwvZ8mydm8n4R
7f8PmwcMTOqRJ4joOfdDgk7qN07pMctcl9UNbqFCcevHmilV42yn/IzO/2NntRkb
PiUgMoOyl7vV07llOXH2KzLu2Z7hUT7ZfzzZvhdL+n90HSPiwjzSEwNHizNVZd7i
Mp0fd2F+5E+0XjsVKwFW+7Mdi0yOypTftJ1RUlfTVGfXahuSIFtklSum7C/KwWj4
/mJu23Vrm8/WLNtpRyZFkdDz5ZMGdlQ15I5w6fPvN3CBI0HTdqGnb4P/bCdM+oeF
9AicZXbVa3MdAr9c6SvLvgAh77jX5jY0tf4kgy/uuPi6IKxiPfAZ0UOq+EBd4W0d
ZNSu23jlTGJ9hvPJ1kAqd+WaYVR9x9Dc2wEVAb70s/w3Eqw4MjQdR+duIM29zxsN
geXn/xtKGCYtr8xcQgsSFQb/hoWhzR1KFjxel4RSVA0OZ/fXEMyCoDQsBL9hE9Xd
VC5L0A56eh5zs6apT2f5v5bzpWyJN8/b98ZnbCbpd3ZZjmlZqf6riv/qrGebewGR
V2FR96QPXTMEhmaT9kKRqBV7d/DPGS5FDR1t50fm6bkUPFLfJfWK9vG9rfvu3FYn
cv698C4Y1bTVBJBeYb2dbiKztBy1F8iXEDgobHrg23SE2YYsMYWPf1dS64t68bkO
WPS4snDTcyo826CKGJE5MfnfL3ah6Rt48YyDCC+5S2c2Vg/ctfC9ER3E6eHiARON
PCNnZqIEDuaxJNj3ewnose8P4BCAzVWo5jY8i9QOyArqHyM8sohFzIVOtmqCtRFu
geAQitIr/tXcDXwsUDG3mtID0L1AOrxXCDXgvjcSt73ORmoWqZfQmmlnd3e9v6fM
GJgZSzdinbh08cGBLidG76r+HFo+cTEriQKsmro/VwllJtRZhFPAZ9z9uUdM7nig
G0/yjQniCwelgrJ2k9YelVLIK/Q8ROKyfc435rBdH3J49mecZOkYroLjE9Zw8XFt
uGhoikOFeHKtf7GcUfu5WvJ5bJhjB695ajmd1kpQm4QpDjl2eP+1olpNDNQdNa2W
OAv0sKyXheHGJGOtP8IX0e668w4ldCAN1bF3q/1AgZiTJwCkyZiqxahSMzp7L87L
xdCUzpNexozB4ZajnplyuqzdF3kXYPKY99/8IeFdaM224UZ+eZ9llV9ZYn4H9DRH
Li/JJVOe4Ma7fjrqf+/OIaZWYv9svUPSFzNJfZ+6T6cqq2UYwh7V7ooIyMVW2CRA
3G9eIHqBMUa12FEJfcNwdoaz164/MDVPYOUH3DCsjUdF5vMuliVDkHWkHtB9+Vuo
18tFWWcibPMvHWVNxDJCEEo8k10tkDj2RdV+l6M/DBGrf1D9YZoT4ktSBCw6iwo1
wLU9N+dcL/zaBFFfBpzyr7W9S9jLBeJpghfN61YAJceonf6proYrQOagpRGk3hKS
dL3ftl41NCBEAoYWAmJRzIyNGozj4EsxveXOV6LhVH2OzhuT5BX3R6Wxktlh8wP2
OmMjSgmb4CvlvuZfzp2wUwi8InxDWt3UHVSuaTKwFrUhsIG1g+4arWFhVEJ9S2tJ
SyMCCrF876CtaklKRpXCpQt/t1qiClb+Tl3aDa+eJE4UU59Mk5beBqryhAQEEpLM
+OB6FSFyMIgo2X19nkcEh1mL6KD/3GG+fVigqPOgrF9PhKxr+0oQNaxtWy27BUbh
F3C1qbp+WVwYmI1V65Hn8Y/IIu8aJ8IUmRcTDBjiC4PxMtUkFtmlSP6lWa7bPN15
dQQ+/5xZzzKZ1ksw1+Tbop/FpLM2HIrYDXHJMH/NmXA7FKYSOYG62/72RqnOtNf2
oWCT0DWAUMaE3X7RX8N5LqKjlXoU3TWKIJPUEbiZk/wGpRJOunnXCf5bM0d8y0HZ
zTRt9VE34CdSnaHU0dbSIXmQ4N3ZSlnUBPnvOPRY21AuhOTWZi+N2cUSizvE576Q
hOaEKXm2Y3SCP6J9HU7nJXzfIwAspYlk/xbfbvcdgrmRA9C8sYJRV8WYT0mIvIGQ
3trE99Fg15m7k957eMI66/pcSpKS7zxi64ZvVabR4hLFxb6mTJIsh4wPGBYlLWHL
4ValFbct08/bDEio6F+7QmXvJ1d7iavc3RMd5T4BiK3kxVe+mUZOC77s6hy4IWkw
hHzKYyfYSuEsSgQhuHa4LwrBQk1AW//xaeolP/QW+z+skhaKI1jhI9OxNW/ZD7ZJ
nETET6UMmoJ4Tyri3RhBHXvTss22l7KbBwjEF7pICeg7T0GQ/U3tMfDEGWpfKb6u
fP0MzZbj3h7vqbdujhlcYZM02m8Ib+gGdjtg69yXA93Vklfc+C9Oje9IdsuPgN+7
hepFLTdInclylbxbcSweCYcuXsP/vCN5txu8iNm7zhWCTXUOT2ojKk+AYttC5+kL
Wc+3u03LEYxeSXYArHGyi9GOtzihvNgmuS+ZtcQ2d7E56lLeint+8XTonNCx1uBa
Enr0FL0y4ovLmeTq5IApnE+FHsMdqkaGV9JQH0vvOFz0XwIl4yLSX9fmaEcwLIhR
JsVBw6eXEKbue12i/F4OE6LB3CqXQQLsxyR9jIi9h1ZG9n83FNSaCNgtkUvNSTNy
om1+Taw+wu+fQ09aJp/qFaETEKwVLcQsgXrFPahMz1OV1RI51z0byPlFoFhmp7ey
ENawrJkUCHXdVDw9SwaOH8TP5bREvsgaMIzdhtnQy6hsn3HdpFh2B7x1bIFJ/qKK
x4ebpZwcl81macnTICF/5uWd87OZIBrZ/QyImGRsHq2I5f0WhM9tzG3k4PTAbrmu
SxjPNSzH/3CNZNXxqDqdd1bwy86tRsfzG0b3qHsp4X7CfYsmikcsxS2TXd4k15t9
TSE7EBmxCTNJOa9xDw7xC8twMuzZqPuSasEjExOw5f2Bm8kkLh4wr3MUUvxC+GBf
YNAuO6TanHVU2aBafuz4io2rOX1efzdxux/34RKU5vdH63BrofrXIQ+vhDiafCb1
ILZ7ROtyvH4VXeMAMsLhwxBb+zQQP1aQHlhMOt/Dmgk5y+gmmdskuQ26FeSiSi7h
0MwBQ0yvkCjaRYzNSXVFgSvCCg9dqcBSaMHszyr7UvdbAkJjXanUDXv0QnyjimRJ
MMwi0TfSBcuAcy4t3Tcy/uW22S7+WshLAL+jY3R2CIsHP/Oqu/xiSR/i7hRvHhzP
viv1HDzAXl3PVnUtovjyMfsx2+U17UszLVdhuJt33s83o8vUhbZWTa1uqk8IdIxZ
95hh/g/ZnS5xvK3feKmEd/O97ZlxGTAP3xyJiReLN5AbqTusAY+5Mo5UceCOzMHg
usYWLhVbABJcErqVuFglXlXYQscrqqK8wUhUYjsr/ASD1xxq80Ue+E0LOIgT+8JQ
y3fPe5DqkcKA95sVEEeq5W8rUtm4uf8dj2/gqMx2CS8794Q9hooP2y8N2tFcyeYN
/uCJQjl8Vhp45mZDxG9zXNmyWOlGliyr9cKRh4QmPWZ6b+FyN1fs6++NBoo6vzEJ
SN5ctoAmJnNAg0UjCwHD3Eyz2ZI/njlm3+cyAM4rFY0/Pemmm7t3aW4znkCccdIj
lMS5e84J+N1/gja43Kl0g0M6ff9hpDy46gYPkId8Si7lbHxdIRIXJwstIZVyilqx
2AzON1eVHNGtPom6pH54mnyI17O2uS6vct+/kkJVxVqfkW+NNz8YilTytYbv0l75
ZUDr0dER/424Dh7U70zF/0KZJ1Y0E6VaqoJqbUHBYHtWoEgtbpU5P11VN+RPSvzF
LnUz9pPgEV6UBNg+fRBdvoPqaDn3/iNsNALphNzfuHQsOzZ+wqmGj2kpAoXoAhZz
yvXvSwJ6nvdVdGdzD3O3i5IwU+aEIl5P3Mf6YqBTCkJPwHOlIUol5zS5YwhxZJux
HrzutZ3l4vuzyByQ6gIjMKDW/FZOj+l3eGCfQe5c73bLXo3TYb0qVIDRH+jqCjhc
zZ0G/y0IbFB4Qy3rbqP0EeCTCsldwhYU9UpLDvRNQPBoX6/zL4U0gb7orDLmQPuS
DDZP6dgidIMPrAhl3gCSb63HlEKYbSTekvBqI0rSEsXESO9JC5Rz6gbvdWu6Qi6g
cOvJHuRx5zlRb+mB4FK2Y4S7oVAXjWJP0HAE0/bjKjbp2a1xG8D12fkkw0K0AoBk
g+/1Ya/WYAOXV2dArfo4AU3EDrAyifKqTHeu2apWPcLAiWIkKTWaEk2bWo+D2GS1
arOIn2Q265sF/57oJiBAid9nF4MlenrnbYSYk2kzJpXDO7c0QPWTXQQojtfoUkvz
TDDeJ0eUaegxjyWHzVhXY7Fc/ocwFHTsLz7yaAN0cTrRrk9zks34jmJTCg4NWbBB
RZf9Ak4+EoKBqPM6MRqWOmZvONGxFQ4af9EI/0B56ZRoa240mIg6xsWn9oqFuOjy
BIiHnTwGq0fzNP8C2/H/PzjMJISi/KaS5AIit04XLUEylsJpzw5jhQ9otqpLd5Wo
pJFnqwQ6u5vnm/Q6BPvqJ0A6A4W+89+e9p9LltkIEBGDAA23pmF6ptENv/gCK3IT
Uw8ltdNc0W5uPeqVu48Uyzey5/OCwpak5OBbIVRMeyTxNEyS3nnlrwsA0/XQhyeL
UbCiLmh0fL36Almdflu67Rrg/uClvMvve7I97zUZNp/TtO9tEwquIujhAXZDj3YK
UnSsuiyNaYfOU1LV3CLRtM/21/46sxMeBP/+/pkiU0f8/EmwtWYd2EviGkouRz4Z
4vo+5jdzY/EIp4e2SguNKPap2kaOlUbNvNXOaAWXBYCJeKx4RFW5HZAXg3BltZBV
9sBWDKOY/uyRsdirx6Jr6X3i80TlvwRiiZZ8Wxw9JCn7I/h9dMhHDdeRuXaAJO5N
qDs/wRYA8YkNFq+6S9R3jOuumSpoqWv68yn/zm1caq3/+pCi1feV1Bm/HYTrm1zg
73cf7VPNb89p1yMsrNSGXU6hQqAl+oS7BdsS1AybUFYIi2044sdL/13fOsMlWz1n
mKD7XPKfaq2ZBVZXHZW8ci+d37HrZesa/feCXNSGolv6QUa9mv8xZwtn0A33PnLD
6wOJ9IgKp643KJVVnAvbARr0X61KgUKCSk9F7KwxyJx5v/p8M3kbjNONNmwBshtq
Xp8J9pu3/rFzq+hf7yvjg/3BEtlzK0djyErR3Cc4cqKWaexIYwxHFSsMllakEGOl
XQShfcRPFGBSXz8r5XXZpwoD1QTMsXSsnlhL0TiLuiUKCeFls2TrKpDWmCKxFPXC
q7ZHcsJyPvBQDy9lS4/QHpRJHwDkKtxarmiNGm7Q0RDvMvY+i+z+TJ4SUKuhQdSs
zUDDHSTtlKfXST+XRykJY/7Cm7+vIrRA3LfdcWwPmOZCXhLDvSpEpnpWb4pZDvnN
OKqCRoCpkbOfaH53npyMGxbtkkHqXXYR/2pdCwYXkDzM9BbvpB8lEW+kDx7vvLG/
qwdYRFnk6EZoxZ6Z0AzTnS4pna4T7EO4xpe6Z6UTzdpJCkflmTQsgjXSjYsmqfqE
61PsF8dWYdSOZeKv6mjxE2C6nzQnvXQVa5SsdfvnnbBKBb/ZpabNrL0eIYF9giAK
Wq4/dHkiHBmUHYYDdPkRmbYDS9lYKopQWFSnuciqKo5l0l+kqeWW3MmYgeMDvs9Z
1MjjuFaSqiOXgVDUH93JFWaxq4kfywO5z5UlbsoobShtR+tfIbYjJnCH9cCE2z/H
I3TOmzS7wbp0/r4zdW2Huv4kBJo5glWtryzksOxq8iSswpGEosCZ7D/+4+lJx+ya
KrhkN8/ADiGPWTbk0SnjhojERCVw6h79p14CWKK3DuXhP0zKAXBuaHI4OGaMz10H
LS32BYuaAvw1dOc1aRImH084+IoAEmvHJwNc3OeH205onnzr+brKs1YrZ6MRQKaT
mkGimZY1WgI7k8oWHgly99eVXg0bxs58OO+9vwVHii+CxPoS1x2MKu41OAZafaQU
PSAQNBg+InhCnnWTRJPTTnZ5XbCLN2Z6A++ynvDmBNZTLJSIkHSa6/7NBG9y2bL5
yRJmsl4+V2a7ebfGvQ/UWDWU0KNp+0qcDf0Q6CzGmIG02ttKGtpGEcUi1gFO5kWC
jYc5qSuo1hlwZL8Eg+n1qIvZnjpNBWfB89nyK99ffiao4yTC2A9ynQ3cYT+MIIjj
/ntK/ChGmaB5OV6FymGWxa6ddQCYqRvXG4Q7Y4FRErdpV7lIza3+vplUg3AuGMvH
0lBxu9DNVbdfJaTDH6DROhspLQMw8Yt3Jy1iHlFrWGi0AXTApQIfWIudtXXz4EVM
Hu7p9DDfl+fMG2ozg+1aa1bXmCP/xkSQ2LLdkl60OU+QphG4sT71brjwOlXHWHNh
CdGoAyVN2wMk+0ZO7zNjxqOHRdabr94fYg9NMpKnyZxOCXuA0oaki/PJJoXCuFe6
9ZKW/eCvLsn6rQs6NbT5Brl+j+q38WiPZkDoi25j1FqHjb56odt59inCHRLymlJ0
s5+YqF26kAWAzEtQt0TeT5ScJ1V6mmHHOTFXKcBooV6z6//2t/iBj3kpnkAY8+2X
3PKycpTQwp6n9m7aJn7J4PknklEizOSankWuswOJOCCBfuxgqG8tyqGa0KNjnmNp
3jmQYE9/l5bYVyBe8x7Hhsnen/aJldSogl2zHMmkKw0nf+77tCiHIFQo2CUDdQbW
gdoMSrOCM7WAe+wIoYRvK5ix2MsOtW12o5bgmLz6h8j8nBjeOosETvzjl07w/OwF
028OvX0xxBxWjWOIhnZqU8khCUjIgDjN4jc5Yn61T6M4WQDyBJrLgVD32ULhFwuO
0eI0FhzcrVWfqmYcgKVYGVUrLcz4dzVHA7H+L1ADxt9pQV/N6NUpGVUN0PSyNem3
ty6QC2HtlhWXeRxC8V2Ls46sq7//4U/YJoFhD6YNunL0DVRkZH6hbhOzL9rkx/eb
/Bqp7Qy8TQiy4fciwCBTM53WhLrWPO4etv3RMCr4nIOtjvNkt/4P00Oip05pcDp3
ZRUGEr6dCjhi1LOvxkWfQ/nKinvrk3h6UkrexnJkQzX1aqeJjA8XJOTZ4YrWeqVV
8ZjP3dvWv2S8hqewOKOqFUyYV67a3MW7dgrxVl9AB4oNtbbYBg0/r6CMn/4ivA0D
cdWIjIABxfHY7QDsbErxc6cbWoatR0lb/W4AyTQ9FL4QSuoDjf8A1xBTD5wjIvR6
iCTaJcblNYFomuIkY2F3z9qwee8rYZSsqgpttKlMQloDuLHRd7I7WXIyWWzuQVq/
O3ILYe/ZnUxvuW+YP9VQB5gTkPtuZa+I1jT+PyC5GAfw53PVgGUVL0MlQtVN+XSf
KtgntAVyTMqmXg04C5hkbkIfX2jObm9EYv7wgkk5ffVREL9mp/HnQsEtRpIGqdxv
4t0bZeWKj2bVwxqdP84YZmEDSLf/BPfw/dRKMegAimbjEgrT3JW+k19t3uT30Ui3
at/87W7aBFR0hQ51B8+qqF7ApQsUuq6BYdBHKY+T7FEzDDLNIyusmJgVEyRVnhQU
Y+MH8B+rQakAd0XOX3yevJ69rmHjPa4hbtRXvTaY5x4iopE+NvTA2JHgnLLA3ehc
qP/eMTTUhc9rntlZ6emdInI+f6ae6mWaG3FEIWAoId8DosdGl1BccGmykFF6FQ2/
7rJzyzXKMbvwlnjBLx/plSa/yUOra46hAaekHo2V/2+GedIFtlfxqJv/vAyKm3wR
WG7Vm0IsWf6w+Ew5XpShijM4P6WjeAT5+/0UWBZ3ePaWgvrY0UIPe1Cpu2pVMmVw
fCX5As6TZKJwv2wtqEvU4/MGIB4JXG2PCafgQ1blsBVWCACmEjwB2ABPpHkkIny0
eFMPmXxgMNnm/Lc4cWmupesPPtF/DFFexf24omXzyMoCYJLkaPLITEkG02CTLY9J
V8aABot44CsjRtdV/cC5d99P6w/ykaMTMcZRgzl9Ro+j+0A3QVe/Me4Do+Q6L9l+
T94OeJaPcT48RYiCgx03K0bn1drFVo+1lr6kViIExsckZ7Ih5sFVaXCQRa27ABz8
jbU1XYjvKswsYytan2h/yov5/HCZRxC4HrLEM3xJAZdl8hwzq2N18yevkfkK5OKu
ZpczVABc+HngkwJV6KiZchKhtpMaJ38fcpGLYDG/TX3ttK0tJyQA1GC9bdhs6Jwp
zwEOV7D+5Hkuq9azCCTswm6E1LuZltKTLwlx/DpB/RzyHbatLjyFw9zWn+ryEVHO
Al5g4pVTg2OjwIHG5QdbLFNQQcqAkjJ40cEDSmtBktP38PL/08kwLvPNRHZ5NjIA
PnJ8rIL+3s+RY5C2d1lvMv5v1VT+m4UXnBguu/Up2JJmxSPTUPn1vekHjcgovUrs
s7EURIciJQtz/SZ1oB1avTJxqvzyoP+Y24CXosX6lB+tRenX42UXYnjtLog6DUcO
kmzdZud/YAH4K0fg8jbomtcXySrS7F8wsQGqTtpTykz2yvOzdgSkAV1EPlbQVU7t
OOzu5nMeZfZM2Eik23PpNN0qArHIL9n8uGNSLFychCQsRUBcY8tKvKqLm643R+Ft
mx23tL8gQ9LkHHsql8rebVQw/94cOgjgpb+GvSAGPQ4j76zMSq+MuWG09JiVTmDR
EQC6rU9K1M++ywahAbq4lYHJWWSZnYKE8OLX59XsGpm54J12HP8GpR48ceyBVnL2
EFZm1vxu/NUQ+eG7F8/4LQTJEAUHE4VtXKkLUN77XVBpA7ZkWq/BgibUNI1lEP8n
RoNkcS1RUiDYiFQSr8CtT+LSpvTocFYbXH2Kg/5nl76EO/SsTFHsogMfYUljk7UQ
lw6JwSHFffx8W3qDD0jp2gq/LNNRxZCtE8dJDrIbWnHhZITszQHXR2n+Iq/Dygqx
jWpZ7CCYE5ejFzrT1D8K/hkTJamPBw9wUgueONNxT/FxIKi/hCBisxuy+aCFh3mh
62ipdZ94rmX+Q3pCPq39s50mBp6mUL+ZF5h+IIfADpfUTAYakXVzIY0cj+4Q8f+v
rgX1XkHoCnsryLJbc3qdp3p908ZsZ+OzvqpmQ74ZyolScGvyo1GFfvuLXCt49ETF
DnCojRemEeAtwZc0sKIeEjRRJs2FlhCXgHZwKPIqT5H2glqa8ccule2MNMpPwszn
zAs5l5jGtShvQX3E3ZQB7u5pQRu4hBwST1vagdP27Eo0toaK+kgpi1U6wJWaULAT
tBFwTQi1DAodLb+1hyNSiCEfvGdCHuAD/BwvMOKqLofpMhgHSO2QHuC4IMEVLmgy
u3iWmz8j+NHZiaPEjJo+hSLk5Qy5DGm1RlL8yvhvAEeWyvRGUf0KJJ2vnLrC6/oI
WZyzGklLW5KNpwJA+E7BJQPjEHwaeFl3bRLFp3Ixm4NRViOrAi0aVEsxhD4/+7GW
LHbOF/0ogGMxcoeBK0XjvXaaRm7gj/BNNOT4XdsXzjHDBPnvPaYe0QzuXNzLdsxL
MH5pRMgC6/Pn8gcKQag/tioLu/bIaq4nwF3ZXRmw7YImTi6GaEbTeYwXDheobxeZ
lbLsysFUW1LttuDS1dKuWyMojgw9gpVP0+kLRZya8R4h0zLmqFT3DMC4RA6ZrnUc
box05Ztt60jH9jIxezu8Gw8lRtM+42bHr/xC0WMqkVuH+gqS1l6i/1ShXE3zHBVE
X0+bLc/Cg4fj6OYkuR16LKjCcL6UWfQdfTui6MCROfYamiuWwr7vgyuFAmnMgNUW
RX78CKZhcYTyd0nDOnIjD/VDXI/nsO5DvZbAuBJQZRDMv2IofzvXqYLU18gRiFKd
3cQddO0EYNK2YxN4x5BpurEyP8IIgLPzv5SwmabRWtHFuIBRRe7o8Q7VgALJ/D7L
KOzsEBJWVfm+sTxxDp7DfICSlsDGahVT8ZH7TnjeP5V6cZrXNTv5ghQMeMx3mhNn
VLT3Ty3589NmXxVxDV9r6RDyoYVI2SnyvpdG1YKYW3v+FGhPDYXU5ttlqgN7ocnr
Jw40C3esG2UqpyFAZ4yEmmeehNhJQ33UhmApR6CLrkKADJYwenEgaVrpnauduqb2
BL7P41bbvtFqgIXbHjjNvRqSDXoIP2iejTxvgpXnpGUG/npD9OfGV1XWlT5lFsWX
19I8u8qW/KpJ0ZtTWG0J2k7kjBIALuX1uVFpjPwQC5yW418Mn3zdwpUq7niLZVkR
oIIVUapoLF/uc8Z2c5pNPNbpivPkINKGy+l/Xr9Hq9Mr8TyJBk3OPFwmzN8gKE02
tzndQsYMQ7pR/5DQ1n03STe6cm/QQzyp6wAQe0M2qdR0r8cNh/8tG+j/MdWR750Z
zS6yM8lTDhdx5tWcEhxJ7B1+ZaJQEMOvjyi6CQ/xf+VuEN1hbPPzgDYyRjtEP+eQ
hPVRBA1QbXgNZGQZyw2fyXwZRnvP/zQoyfIvCLIl2uq3nVLZ5NPaYWdqw1OQua5d
NUGapHrN0mooEzFvK4n6RUTrZRmLtHrq1+zYJ77q1D+aZ6fgE88qoU0FlGQNwxCW
M5lwdOQATMKYqiSR9vGW3I9XId3N9mN6BtGOdAjR+QPH8xb96+6M2oZzM7ZoH9uU
pFOdx8XZ6rJwMvrXgLcyC7T1oMGoWW09p47jQ/ydsXHcYfblIWEN+ZrGzoQKZ21L
ORyaxDAXeO3V04KQHv9c4QC8/dDaGFxzPbtZoUkh/apdvYEaFaI8YaiPavuooc4h
ZXQ7rRzT7T9VhQxd/Xgh03bpt0nGYxZamJS0c5HulDHrr2FJYlNlPTTrSumWIhjF
hX9HqGZ1ijwkVhx3dJpCP/lsOgTihnjWDK4h0elG8MYQrM7Q3M8NSDh2+KC5R3eH
2T5JCGnblWrnJjWGOw8HEmazhEg533rZURyuuBqnMbt4OVuzHaJEPi0FcurKL3fG
S2FUa2VObF59L9/5C79SLR7eZrg3lwgFG+d+/vmsYhh+Nch0EQ4i/+6odGOsCSML
anNEOPFX8D1ElxbVUqmtpvhdDKdsO8d1HG5gEuHMXhy28AwwzyDRzekMkgnwn7nn
+PIhizRPAcYql5q31ODJH6OgQo+i+810M1KzXGjR1VP1EfrGPtxD00ZjXx7pSJlq
tSSwq57uasroaP11oUPiEoL2bgwGyhTQGViQGfK+eUyxOwL1fCju6kBl4EwWw1vf
i959f3WyzFTAJ4r3p6ibtnqIvMQGlpAuSK44iICgWPRAiy22Xi3S6AJ6HJX1DzIp
jqpp5K1aKXywP2jTWe1hvBpF/m4zGC71op5/KQRI1++m0SwJ4RyEdGdDQaQUwU00
LyglBrkiNx4Rnqknf/g/k1rgkX/WJWX0nlHTHcMsTQHOloV5qpJRuZVykCQeww3t
pAZhB4TYJCvZcDATHY+eURRZYrBkSCK/F+CQnYKPHU/o1/0FTaKmhdYKNFSPHAmf
L1cwiBTSCJtg+nIqP3xImjAIt/Z1ZYwhRCDssHhKmyK5VYTZpEm3X5KBS7JWe/Jz
kg9dhAMDsGk1L7cp6pgTYti3sWlNb9VZF9fS4ZUfC2GS80X6lzjWxpJRP+B6aN2D
FpIp3mpBg++g3eiQ9wSvfzKVfJscd62ly+nRKw2Pn107NfNRucT2do5L1DVY+2/D
C+xDjcDoc0BqRwiBn0YHqoOBePF7w7r1Fs5QuIRIc1woBOPXwRaMJu+ftY8G3lrC
sA95eE/pNilryU1SNrkeHKyORzGKvbeR8ZBAPi69VAPrLYj5fI/dUJZ6b2IkTLlH
`protect end_protected