`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24224 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
/vEkqJfyK/81z5lf9X8oFatn1sSwjEoDyA2afh56iCg6oIqBNYp0nC/oKYW6Ng1f
OjJDpRvYX7C6sjbteicMpLnn9kxC/C2PPY5MTVKXUcgku5PZye/QvIknzvRsGvBu
IIhrfEPusC5jOaFM1C1K02LBF2joaeFrxWJo53CJnCjXq7RC1yfUKBKXnU4L6kVh
NoHNXQvOn3OqffKg28W5mrXUzU/NvEAJRfqOn8rNl6D+nTPzEUpeuzZGwSFHf+xi
7kr7+b5SALjakO4Cafk0b+M9EGrszxjKfq17qscx2mBf6Uwr5yOOgQDsr7nQGVbB
rDDD+XDpm6oPQgw1LCG3dtebp5WJZWOAS8O3PmGFkGWqrWkgBDzVUZ8ZcJRCw3FA
jy+vxN+TEV5O9Tz340p0EIAH3aOwUcX+M/C/CyfcDQ3hqbBhZegbjZAHGEFX+U5w
wIQ+LepEyYpkgSZpipKX99/feMyj03rvDIgjLFj5hgBktE9Xzw2g5EZLTwtQRg8U
8YmPikCESzc8p6op7sQq0N2Ir24USquzIyO87q7SFcXwJdlGI7oJEhBX2Rr3VTsh
iH5Qiw13WDURVoFa9MBe92xGTnm/HSprLPJZnVqMD0xp2/VPS1PBe8xORhaVNafN
MG0eVIG6bUaEXuCQx9+V+ryKb+WR/3D2/h4LNwVCy/ddF5n7MSOjm8q/Xu4bRQ3j
8tdd8N7dOCfZyI/UfDjxttWV64F7fe9hTi16XXuokRqaWfHaoldN/M96dQ6MFMC/
qEMLVViEmHE5WE0YCzZ0KibSIJ1L7I3wWdpvMTnhbDJn2JhH+GStbAw5YoiLvQlY
jpEJBLt2/tz5Ce6qCo4WLPMywgFC6JSRaXSxENckEkFWXpWushAh6HR41y9CWbUU
TwXRR315+eSRcIxEuOKnM6jQtf6O3jZKUgRXW5qxj8Ayxu3L1TK2qdf+TX7ioOyI
DItpEoGDwzqI2i0mSjLiabyh9SdpAk8Qa1jAjmkYpNWGwT9b9X1X2zfkt+7nXYG0
72/VwPvxYTqB31lFWTzdTyTb6nf/etubk73QQt3HYSo/g2/PCJ+u4kr1bPluw/HH
3YErEF9+f7LbLLp2Xkw2FN/T19/KOAedqNIWcRdxa3DIBVMCoug5OuvAmLAlVaYU
RWvUesSaOVxrAMenVKF35XrBQ4EUj3lgt24UhFOxSP8CzafkodtEcmUA02Z7V+SU
YjwJWiEF+ewAL4O0r/C35QttIszGVYAsoZDZ+LTuD1VR+BNPsRrQsp3mJj1Pj2+W
4Snz1KOc4bae9eorVxnAVgPWEf9f96PJ4j3rWaYVW3tJ/tuGETSvRQKtSVdoE/YG
fmDAYTnojy7gYjNP8+qRfrIu6midTN7vDuEZCMOJWIqRaUVn3b8BiulqcEEo6WT3
+127APCnz1AIWCE/OfObA3JeD2vraBEkPV2dsXchLATv5DE9eS0wi9LUVEpCEjlT
/Rl+Uxp7Cb1dsdqCmzjVCsDps9tafbD8b6gS4Zk05RTnMlj3L1STyYcGO9njScBn
X9lNVi5uEIIKt+xnAJl7sW+ntyS3Uyc0bNuscbVD6KbdmzImR7ULQoK9NBtfJAmR
w+p233gEczTlFLJYJ6oo+FG9S2YcY2QOR03GZmNGoRTGmWu71fRP85tgNSNHS8BW
zcUCMgh64DQHQAE7SKT8PfcIniIxvEvBZWgBN1fvnSRSf0kjbx0vIvVTdQDFAwSV
KQv42RjbuhQ+NN6LH0FpLfnI+HCz7zAq8Uul6An1ecUY+OezbJv0/n1mWKJiu+qk
BdG0B+MUfJY4a+BgFjgB4xAfu9N+2meEdrB7qIKG/TpOgUVEZbQ/g10gWOUqGiOA
CEnKRkYqLr35dmXb9VNgM+0gQud/Hk4P+cXrDnwl69e2I3qyyqcoBLj50zzhSX2M
5IPoPmOVeV3bimtWuPRsjYk8vDPE1bgXSfeLmkyk92BcIUTulclMofqBceY8+PAj
3t9o5JB4Y9f/+dpTf3wQqUH9t1C5wHIm5sWE82hS0HStP12Wfa2SEqTevu5rbpvl
ytPEOKI9ggFNRBVbgZtGAtu/tGtdnI3jUWxmstNBt9sPn+R0Ej0QTclu5FnFXyHJ
X7pCvpK/n6NH0WgF04/N4Lh1CIgJ18UeRLKQL7ZGnJmnM7zyglpgdAy4Lmry4bqi
N1QHZDjH3gZrTKp+X+jCP8Qt6fQ2I9T4IYjJImr9AEiIBFn/a/xDe4WM6IO1N64e
Wj2FKf6jSs/4yWxbOHKi2a9MmF70m6aPK1Ky+kKqwJafx4ZbxJ/YYUB45afduZcz
K3asmQ0bwPcBX/AeEMb08SYg47y3zL3qzd4IID6IhKm+I6cg9gigP3GZ2vYENzMy
2XJRPe7LTTZvkA8BnEV9C9Kd9v79ssUCuTiyxFZvyp9A6MRXcy9WckHYU4txlW5N
JuR3DIkO9XG8NTno6fwo4QWMRgtor2WYHxFlIh8HfGXoyMWkiOfEl/DjomZXps+O
YWRFTfyAYXqXRwjugOmgl6eoJ8F+mThVazDiq7NSguHon0vUYHoT+QOPZjpdx3nV
pGz0JJqIZ95F3gFLeFmrBZir2wQMPgVF0BV1aZEHdpSiR62754W0tt2SlJe461vF
kUOZuRkHqdR9MJWP09XykE1XWWn7xUQm6mXqoJtEoH9fLhxVyFd72jnSwx5evj0i
w7vLNZbIj2OmXtBegP6ZIXPnxhDS1svvU6iN13al7Scb0rEN3RAjTU3OVy3Z07eV
+A8jVtBqw1yNNhWkAbHYGu9VFFq0i4OkKh5uVHtJ2XoBSngYTBHGoCnLF6/10KaD
I9EiMQsv8ZeaykLSWkFX+EOAL85iOch4waRUzt+ze/UWwg/HKqtf8Oe9wEpn0tnq
0i7v0tKq+mSl4RQYDRbcGrC/b3xIp+A3b6iULngO+v5+2rglKFtfx6Gov6XRZzR4
5rXBuGd4vsKxvS0W8jdNPhihO/Ql0DNzcqGbBrUZZ1EgNt502Gt6d3wAfjM7z7Sp
jsqv1wL7BEPOTMuHtKCJYj5hZa9qIoQifMCmZIkq1H/CqHG+f/sQn28ATk1oNxps
Ewn8uNkd6IHBg9cx03Rm7rkYvY9rhVYsKs0aUkKyvpEVQ4uaH1/4pgNXx7OyNxbu
LBFh+SZuDAj4q8Wz4zT1UKE3cTNnHBWQ1QvVDg4/H/Q7t7PK/3VV4/QFsZ2Q5Ono
BDpDNYOQD/0HoU3e9fMGzcSto8t7QaZwoIgYfcwcnH1u6t46UeNUXVvB/1JZlGQK
cGFC9YsBFz+eA6aUTK0C2Af9AzoyiFgY9Yho9y5Dr0yK9QRztAQ5hRbnOE47AVP4
S2WAsR7Yoa+MAahVgzHPP7H2p1s82xxz/YWx9aJmXxqG9OQVzNJWlJUbkbatLekB
ycjso3ZSUHWSxt1IBj7b8GlvO0ofhc/hnkMBw5ZUghLzy9rp264swgfVzabhAl9U
IG9bgY1Pvp+mpH5qbEWW+nXw3w7LxdYS+chiMvNxghh+vgygkbpRpN9RqLddG+pN
U6stRMxqN/7oIDXa3AXXg+ZyQq/pN8j70JtQbjTHgSoEuIGV2Ul1Lh9MB1t/asOs
DTZL3FZgXmw/a+0DZSeqqI3zcfVzh1HzdUfBWRhHZK3DSHKd7PF+JDu0bs7Akm/D
nATSrsvtsTs2xZoPYqaSAoGOQ5RnJvnp+QZ3eHGhEs9M4RlRdticRv/rlOWehrwT
zevmuhfB/AtCC1dEeFFiWIrgDBIs1WxmPK8IZb7G0olXEWW0Y87RtD2RPCHQhGU2
1KFNtoxTJyVg1wzoXQp6BsH9Sba3ATzpeqm7N0E94v+9TtClj52evfxgbCwVyUqC
bVSion6O99WHJDAM43QAb662NIQyVpGl0AKO/OyfjIyTVUGbTKziP2ivmdIITbKx
KphipcG+Hzjr+IfBzn/K6o2vLXq6GKKLoI+FaOWQLDwCC8r7pBT3/m1i+xu7GU8a
/Oq+niiGxVeyu6gC1Pv49cWU0/9k9VU6omnLGdIWArewVzKTsbjPm6rQO+6lrBsj
btlvR4Hg1sv3PGzka4sI/xLJYCZWat0vlYrQ9u+EoTI1hbstx0COSZCxFUiSshKz
bSOI8PL+1VBvsfdHwBh9w5P4UBuzRGjy3szJtsgksVhF9MWsZu4BtzfOP8r2T5Z/
bEs4bejp//Kz/N32k2qO+OmZ2YPkIUwwqWswG6JCbM87/udz1gxtBBFRMubASf94
Bz7CXFUob7H92geCKacdpAhfZh+BGwR/TckmINr9VOO3Cs12vq5/S6PXnwc76UqM
2H3H5GOGh9i6bG9I4iRsZ74R2jttNbOYOLfku/TsisMNWpiEdWdrmclesN1WlarJ
OhAccr5PSebRnr/qtG+RzmKMSYnwkzBcX9Tfc1cfDCuYzs55HZAlk6OU+MtO4ePD
FMt/0r4GIfOi9Q6POHRfU53Urx0hQjJDZ6iTtmvT71Ou9KdPfwhketLsaE6HciQ9
1r9Mit7Kps0hwLJdLbgk6C3yMuNkI5ROp888AhnEn6USr2yO/PPR+m70OYu+MA/B
dHCKbBEO6neTQ+G9M3qkjHT0iQphxIXro4Gq0aKhnBNmGa3sm0zOXUemDm2gDnV1
L2C7v+TFwZ2LqyrKsjn/pW6Gx68lhUqZYgTKrrR5VuQoQQ4xfB6/3tTaFgdtZsK5
ziNTVPUW6zE+LngJX+0ek0zBiKbR1ylRJn0uJMoKxZ1gwlZb32Ypsdu843qowdxa
X9Nia+XeSPju/VpYHUAeNf52Fv7sZpfe//bQwL3deLi4iv0MrMLEGjJlBlxTE4mD
TCUry3ScWaiPKGq1uSILgOdgxvl5hS2AKGmeoit+M0+RT2su7Sq1GOy4wCVR48kx
4BcNP2RcKHk8CsCSsVkK11411eJ51JCeAVV1anFA5KasQLdFkuq+MKiMRoy1HAPk
bwIoDOfehiTQcijqIFcYSqVq507+ASTk0333yK1sLc5pYvaecuvv55oTQ5ff7Xdc
TqV/raC3ODgV/cftLqD0W7juNpGwNI24ZClQjstZ13n/tBnLPXVJz4zScFQSoYH5
H0NO/DNroKR3q9IwMTRXv8rIJuHY5UtzP8gPVP/+3hgE2aj1dqlhK/cQBIf/60zI
9LzYLAwVR0P7RZEsapNE9sH1PFHwa7EEJX+yha+RZCT9QoKAR/rXoqI/I1ncL9LV
Xxsj+XxC0sEcfJOXVRLNcQXxbrj/ofqTYZdnu0HkWuKo6bFieb82ly0MsTjVxAdX
b6JMeOXlqzET3kgtWf7yuDUe00gjgmQtXMG+SmRTMtYQlXaCH1EKtOmb12S+gRr1
kcs9Rh4T5RpjuWBdAAHlycgp13aGTMou0oAAfL/hws0TpsKg2sxc5MCDk4SP1cYS
EhyVlCwfdIFsK9ST1Mpn8brE+j9HgnJFEuHKUnBDe4UXbwRQg1OIZgybGygX0X3Y
gM1B/1MW2Pe9pOKANH4dtLv2G6g4PZm4BTGNhx0Igack+nh4kzb1KvVpYdonh72d
aN0rQ9AlwUwhGyFHt36tjZPUqKwLhIyYNBBTPspFjsGEBPpGdgYKZ/Pcv3sbephp
0hbNe8iRoior7OgGWaX0xtyt41Q18h9dqlGv7cJCxm5ARxjLLGnU2OCdGezgZvKU
o/kaPN7J7ZAfsFEHAgMiZAl5QDYM2oFg9qeD22OimHHk2s6GidnrKZsYrjvQV79b
+VoN9JrM3ZXjXpBwtKutlwnC6lICKFNcGth+6fuptwFWFHe8+iedWDSSb/QlBMXw
3TcY+A61wrTaDIurV+LaI9Kq0JV3YiZNCUjuG4k4Qu97a72t9MHaYPLu6DPrQJ+1
U+GInu+byy0MZsHkDJjOBVwMK9dqNly/CZKJQufKHY60tek2Zr/DkjX3m6cM2I6l
VXBJbMKvSYdO1mKtd1tP5ds2KTldhv5G0JTydh/eYY1rjf38bvwvI1/ZL204wYr/
ygh2+xwpcxICc4fkLAKdCEAswVpxxTxmC+UWOOBbG1+mI1XzDYXGTk5tkNrNX21I
o0bcoE0gflt25OD4PDyUTsBC6PlKCqERwiQbALMWXvJadlBtXNoRwIHKrJ2/Y2B6
3FD46N99cEzTcycsTCYqPDTHuMJ6bOjAEgMly5KAW6sUyCryX5HzijNgJ62N8Zl6
tDcD0EWyUSdlCQ5AndWozyRzsGKu9984x1rflODGUONEAAKK4RhBqK5M0zHvPPFy
ngMNkz1Nb1oZSn855uej4wLrYx0NuL/BPX49C+qXT+3/Dkl5kIR267jA5k/VCXBA
fNqrzDizmb4CQ7IVnKMo1j/xKh3VC4U8A1SIb/CV4gmZ5UsCCSek0++hvaCypH5I
51MB4thN+d44fpWBhqFphNxO7ROT8vb5q7x8HwPd8pQyS+rMaX6HQ95kEVrG/7jn
uiLZt9r7O/O88Jz+Swh0E7aCMh9d4IcaYkC+xO2pn32MUNCS7gn4/6eMZaZCMijy
JzTPFyON5Aj9I+lwOpSNJHesTpljbTOP191LO3JM6bgkIdZQ5/k21NV156huUW7d
ATEDXmLFno9kk6AwUaWu9sR92ClGsmoOttNa0HVSGRDxowbJ3M5aG4cuQxCgZ61M
ZuwVJSz8IdUJZCEc7pNTbEKEEQa7HswyrIYybPAasXRk24oqlFBZ0nuwiKGns8Z0
lV/ZIxbtA92PtGtrk2dEGmxrKCDDvVrWUIEk9BAGGO3UOrFCDG6FFsn1H2zf4AwZ
wAQgMX6fn2aL9kEzboUQrjQ23bXgz8fe90qJ+fiMpNAAvczxHtCRmhM5InMKNAFd
NLtxvi4GDx54XUXBbXlGN6EiMqnQWmptH4EGIsMgkCY9MIGEus5rKXezqN+rEEHy
gbxy6zPHIayFexHjbmTiHP1jnO+UnyFqPw5bYpvo3aVuhoIrjBb/RXGQlQkI0/xK
3Z3EAGfNvuCSd85pUmqZXg173CCg5PpsgM5iSkMDt5twIc1dnDnSyzl2cr7OEt5N
ObxLB3B371gVbHToWV3rcFJY1GNCRDITkAkTYNz5i4WEcdarUhFf/4ekRLPOuwm3
ffmMX/kG4vbn6/tBdAgTQuzALqrS4+kPxlN0FUxmNf/nlFE/hlhzxM1Txhcz640S
gUL54WsIQ373BbdTZqQ9RgcwgKL0yfHa2jstp2eUNsM+zfm3HebboeaSzXlnKaJG
cKvDvxM55v/1F2yG5LR0qwOlYAEI787ovxWMi+td8HOKyeMKktY7go3z22ViFGh0
MjtqkIAi2jVBdTC3FBZJKTHdtIF2hPHV1LLvJgoCfBr7d9HsTOX9M2KHxukBHAHH
CGGP7iKwzddQVNME45Y593wJIRpwnjCEhgb4ZwFQ91zKxlHRJqP45/aQ1sBB83TU
6a+hWDOTw+Sv+voG9I1VnppTmebJpBINXtN4xxVt4DPBPXdC1Oh98JLFro5FXp6n
RFoYUQ8EN+Fs+Tx/pxJGeWenCij/KBzg7lWFhWhse8+c/oRey2M0WkwmULH6xPSx
LKwC9wnxl8WZupi5WP561GKoey6drePbBiGY6LA63AITL4tbK24S+XH8h9VOAkjs
y1UF9MEhk1mmmFK5UkLWa/xXv/rJEYKx1VCxe7OzcjKT7wHapNOcQtIUMa/3xPul
WM3gS3sjfDvEP05kwf2N0nN2KZYsUR3/I/CypJTX1yDGvWFd/9fQ9pXgG0O0lqhW
mvb9JTAc/vGO5bpTYLDfqZCUPcv6imJAby0Fe7X6x9rEWlJNfQtI9z/xh9V1nw37
6VJjnApzk0DeyZ6eQt/QQyi0MEOJovPWQxfp8XmpLB8ifNFyU3Mtv6Gu7/a8Urx7
N5JY9IPnX2SmjzB3mhoQg1aGf7+LYaxviTAR99CXT9ctj84/HC10Jx2hsqvRa6Y7
DemLhs+8KECh1G3WeDphLykz5S4EpQADZpTRf5xDm/DRRCuyK8w8ItVew7CRQFfX
153ZWNM2jC7IaLL2Yb01xpNtkNeqnnV+ikfcLRPa6jMb4elvie6O+Zk9/VtAb9zO
/7coDGFLp6vCS89y5aoUbWxrvf1anTxEIIjwGUamBySZ8vgDoRmBymllokhgIgeu
exVe4+sIAIUiDeua+WdjM9vgDnqCdmTkc+6l3WWPO3dGOoZrDQjltQLnH7IAT/JW
vwWVL+iT/sg0tkwE7Y5NfC9CSjNkZOvg2Zy00W3yZbazEvrrSAPeiSe8aSODZVAw
7h8oVakx2xYIS9U129wTo+QijO+6f2uBQ91SiiipzFaAtZ6fQIw3Xa6XWph0zs/l
v3TBQp4u5rn8IQ1kftskdnVVP3rk1bkblkE+vXXWf7mGOz1brkH8VmzlJIeVyhRv
thOLB+41zOndsdxcbkhXN4Qfpo6Tug9B7VEcF/ua5Zqs7Zov12YuhSjnPKF4Agu8
3zuYF9U39ojSq/0WHxZf6AROrY89nd2xli1H3aaIcCpWA7ptFFi/ZGe/+dyQcNIh
CwvMvhkNgSpV02ZCNvxbmdJaN+/1brRlOEurvC4HnMyFf8MZ/NEAJExhYTv9Oa7C
3T3fsV0p5wy5WpO8b8pdg3rkLVsscbV4Ahmtc/baWnV6IFUEQg8ubtRz6VnYQ7n1
dEkosrxvs4U18Xm2xtXWRU2YsjUigBKidXJqCku69yzN9/TZJwiYf2HMAc8FTBOe
oZOv4wDvYxLibV09ewChAR4hRUw64B7Z/hnjiRP1iNVVODJZj8g1aqruzvSi+Jbn
5k3A7CNxGHVduug7gKm5aeRcsk+bavuc4IMAV2GiJtyFS3oN3mJFysyr25n284Ut
p7b70ryFRx1FeFUJWxZBARPLcFPULTnxasHmQpd6SnfW6FZTXWmMMy/n1Cw15b4g
zJT2FxvU2MTtsBFB4vyD/WSSwm5K2pfBjpjt25F9qek2FOGIJjD/BEjIdi1G44tY
VKJOikpOJ4xykLhULBoA6c0M8XHyvqYdmEvDRWi+Q5kJ/kkk+KlDG4GFebGaae67
pS5lWY+OfhzhMnpsupiE8Jtqsn1vQReV377DOWBpFEXXdVP+VhZpIiYfVVFVwTE1
yhIKX+V3yYhNeTPQ7mm9oJ13TcQrXITpJ+glUqCv0R8jYqXFq5mh3fixvd30r8N/
cmovsCCtR/83GkCX+PvIQh52LUKPjJUzgIfSZgSBHOsWmCf103306TPcC4BbPIaa
TykFTig5Yg1cppMq9dma93L9KekMR0zuCCoU9IubMWVc+FO+dHaP14KXvsVkqNQS
YVp5yrU8K5HAHhW855Gv6PyCgaifuf9o0t3h4VnzPloBWuMNy58ahEt5Piv9Olw9
iaEYucAPw1hvhtODPbLeLrLBRfz6bKUEwRVwDMmH8zFoKPhDMbTy1B+iDf49y6lL
HuzfOs+voPnPYsGz6rmcGDSjMmUkI7QabOIcHRPmXOE6oE5AiPdLpiWMjAmEMZ5u
hmbBkMCjlj2R16efYFsF6QL5M+nepxFBnRdO6xUX2xXLraSktJgqtwVr9KfqJv++
tLahj8M7Lalj9S+OpnskSW/7bKG7qr7O5ticXTh6hL9Atj09q6GlVNIB6/bQA4wj
OE4ASGyCF+4VFHxUn2Kfmrbov615h9vuXcmNZGhE6YZ4z7qc3oLkGHcvmO/FaabW
aC418ucm14er+jBhFvmzievx2CKE8EgmFXCy9zZvv5hj76PDgZIpHawG6tZZnvSJ
5oNPGfru6t7fHowwoi9bkydDdHp3NngebdqO2N7+1DmF+nTOlWrdx7CoI6ATuY8R
Am/nIMevfPAtXwHrOSp5djQz8WYeRlAvuu7oeewHKPKlQc4mQsDc83pl1ppYyv5M
xESeh1mMRgMWSS/5I12+KfdwusOKrwjA1W5i5+LiQZfFKeGqY2ESHLFqqTZf7XfP
7SBOuv/wl+o+/wqvkJ/k83kM15x8Ha/KOu4AH9CIRI1u1cWOQXODnknede7WoWCd
BSs3iZQb5lOo8niDIn/ABjRCQ+0A15fG84hgF6ohnqKCFrOVhJIMICAxOsGCVhiv
2amy6jctmPG1iebKHJ4agLTqj7TtShp49a6w2Mwy6vjKFj4RRTARkj4ycyDSzUDn
mgiwsiAS3ex1E/ABA0SY95p+NHpSAg5lfMTC2+6TddOW1S+K2/6hBArky+aemRqU
vyLqNpcnzPnr07S7GnA3CxBJvp9UN6sl0ludi0GLTE8P+d+BzMp3X+vOFX+cREqm
JX8P0ZfOqzLAQT0v05Wpx1AIIJZW/L+nlw54UcXEblBmkaEai14t2KOE76lm7Lx3
hluZd+82nLIYZjYnSlD7IDTsfanl8BlS2We18TjaWV210Ob3g/yf0mbd299fPKxK
f+23y8eWRfCc4OdSFcrqMy7ZaWkWPHKycnhaHCSEOkO7ksc/UmMGjTvfKV1fP/ZB
1xjmGITyVkRh0/w2ut1Q3kcWpOBPo4LXejzWJXAfrPT56VfgHKqYH/6dEizY3KjT
rq0rCYyJvr+Ae83geTvrG48eZuwD/DF1m5KM4aaToGt24gppoSIHpUKmCE8Xedt+
h3TG3PpCjisNgn0i75NcczYX+nWvdNTe37Glop4cOJaq2wOwthMol4UDPHBsWAGf
pBugPid+9vyfLzpGaXeKl95D4fDu/vwbzChOgc6sJxRLDCV6Ezwev+kge7IIH98m
Zy7qQx/5gNLrpfEmRKTTBRLnuSNyjIHyAASIN6bZM8f6vrOTtzPSQq4v24oC490Y
CwohgUn1+EehUJDs7oMrXwhaRc04JeigA4snj7h2FcqCSVMcX1XNaR7KRtfPNh2A
seZd7kB98iLU/qbGPZ58z2nm4TDs4BcFTLZb3Vp+OrKmTO6rQDKRieJChMlddAym
X8n4FAENZXkuGthK16TvNFPOHQ1w7teK+sbuZPoscaDEdoRjh+WVGhvu5PiiR++j
LmXNLXE+HuwdaO6knLJeUD6l0s1eyoAaE2CcDCLKhyeQ71hxcXkpPtoc3oC5DwWn
SOfdi3kmah50DIMN+8ahuh9rA8R0SOmGlPEvBJ5T1CsTkgOBl/dNgZuuboQ2Yiio
rx9kBAeQhTKePjx7JQCS19FMiMYa5VtVktF1uuel6sJ63e7ABAYQU5q81A1RSGET
ovJsEtXr+TX3UyPOPM7x49SBtxP3DhXH2Db0UjFbkg2VAdk3nrF3027466MNfgCc
98lHCbU3JLKeexcPWRuVZBfeSmLz3yLcY11Otmimds5P4M+ILIIJNOoZxjI2f31X
eB2Bgcw8EgKm/DKNIE5czbq5y5M2cOYHgblxo6npCZNEpNIAmkiTE3xBUnYAP829
ZDbGafuexDf4M1R+3KykNUz3BnC/Cs132DbN/nPCjC2Bn+IszQEDQoswVYtKwfaX
ZVNgHz3oOLabl9BkarEDBFdHNWGu+ECmVi+Z1urivTr4itjvcGBhLIZOsrcF2GLI
oMZPa5IIisy3VRocqJEj3YIovVtTihCyw0sQGv/2dHyYcwS6feuK+jWhInwaAP85
ICufIeOH5kIZV6I4HsZFJ7JdxH+IJO2o14mPcbLIEEqy3fj9C8wCegZOYOJm7Ouw
910YuY6rDwIr0V1AnFn7clP2k//7iDx+7zeWyaf+kHY2NYH1O2LVzHv55m+p2rO8
k5XiBMibEYHwAfCDLZk9S9AQFVzYkWZKLNZG4UWLEo9uzROXqYuUyhXQbmOUFPOs
E0DS+2182VO9vbNEfwR2+48Zu++XqNfcc9otvehXOmMbKHyuHRfKIIBAad6gBjp0
k31fbOy1wNhUUZxKzOOGX/mfULYwO1KrMZ/w3tzm35yWV0wyBCCIbdvGp8wwYnM2
W2ki7uIzSn+lJQoslrJHahxElvBBgDUUF8hr4vzFUhNq2GQIDDYWd0HIDaTjbMba
uoGVL0Z+n+bWQQQsAQik3NNdfXABETGbcNUBfg1gNw0dkdmoK9Qzn6gza4k3ylXO
6x/F8PXggbuipmG4t0X7CKD1nscr60z+rh4ivMyxpbXuYyyJzYlHIjelk5NobMrC
8KQaiaBCAc5M/Ey3cvtaLBpMOL7A4hMgN1Rh45UL4cvKyDtBNjRZsp+ARgmaDKjd
JMsEDO4+2xh1Boxtw4bYoZmo9cJDm+LTQxOLUeSmfbA8sloH5jBQYROLfmz2PIXb
S06vRtvWvYaJyCRtSwsIYpkxORAjgB6cBlUHLGVIp04e30TWyx96Pg9vvWqFcD86
j7pCSB76Yx4cEa7fNjF/zM6jsZlcxihBIT6szy14f9XFdm1Mj6W/XueQJGgYhxMM
PS9nFoWCsP1wPaPUAxBjps18fXccQEmODDZVJ707AgPw7RU47RkrSfRmJyR5tWLV
ix+X4DQRaj7p+cqVLptENttAUywDnTmM4kQQhaAPitZPIChTttKC4wRagAgWeMs3
fr3twJ8oWOK54Bwe1Ho532lkT0oZxyomctMeunfuSSmZ2FhZJpu4bD2GdytFq3PG
0m+dQxktfHXfz4eDJzRrhEKtQXPylfp3V8ShbqlSWs0CuPjY4tG8dByDuNO1BxNO
MXi8205/FGVoM8Xj79CgCUq64sicGDFlt17rZzbE63FFvJloYrhaKM/wTdEZ+w/C
4BVhqZVuVJHW/2pK7N+atlMs4gNknr5OQbB0qvg2GS2bdxzj/VfBIUOio4pF/tAH
36qnf4Xf17sOBWQ54JGEiaPoWf6dC2I6x1OO6szB8h3uT+WfABRzvev2Wj4KuwqK
/uzw8ubE1aXdtmSUlsm+UjefCsrC30Y1C5dVWH+I1u15xTxBRDaDLa/hyi8pw3gF
LdwRLeJEeKRBgh9SKY6Rjp9zmwn2dWDCL5XiBJhOKO41pUHmJQv3CKDU6m90lx7q
MwRjmUPsBe8M+Oxq5SEotBAElw0UFdLDlxawxRiEyCXciZqG+maE8Oym0OwHul9C
R/G3HiBfentdcwfESMvWjPuyvPD++XF/szwJPULtm+Y9KpCd1Vi9Spukth5QbM97
NiJ1VFdITNMu23yRTp4t4Qj5ADLNDFkqs+ZUEWisfOwHEMOdxGNm3kK0sxp2TMyV
k5WmJhBOz8jya0VNFzGZCAu5dgpXmHl+SwN20xkUED/ashGA+9IMuI5RH9xhNmja
tHUER/tgJ6lkn1hQ5QuMvg+vSapQNY1K4Oh+VZl9qATCjBARZzF48GcLKbGQvykR
vBQQW6pXjxnwPG4/uk0Ebs4mwoVk6IMySEcyIegKA6KV4uZqozcHDcMdxqeJ3EEe
eLfyWOtXVQSaJ6v+vfCCxuF+pxN7/4eY/6Yk0hWQVscvEvOyXOIfd8k4jnYskepT
Z8vFW14IXwDXENwAWfPUM4B4nar84UFfcackpi7SVpI7johMx39Ojug/9J7AUJKB
hvy4IorDk/xEqCvIzQvNFzpWl8B0I7bLfrYstsCSBhBAHAC7gFe4QOwPHPK8yaj1
lTN650p6o3Sq3i0VdNgEnCYuEZ+8G5r2VYCslp2I3ZVnkmd6p2fJzO425cUZQDYo
3pK54qiqTg83BI/MuOIJCXHr9yj+BCu8SaGhD0pzZkmP8SdE7zLoWfYkdfRPMP4g
LXQP8Ku9Xt0u215V4BFa/3mNQMZCYk2xEl3vrxooYg/EniXPFKWcAPOAJeXyEaBB
1dxf0+4SOmaz+gzeAkkSlbDrsATSXSwIt9vFI78ZeutwDzkPLKtXkXmMwPtluV5H
gU2Yt9gbyC0kvU+QOrSKXApXcxvVz+A4pCmvWRlvaXQ+HOGl2ruNRT3HPaUVGNmx
+FEoVI5jFluVPMVUdp605T09tvp8KK2qpHzefcuT/6jm3PKldd7DbCecCDvdEYyN
BiUwv8+5RDeuz7tKxJdaQW+gpJKEK15vCmYAO0re1ZOZVYO/fGr9en91ksMisA3w
rrfqIudBXMszu3YFGeEhMI5JC15EW3bI2QT9wvAv/1Boju9CNryXpbTPPKvTPxRn
zU4B4FA2nRZ8Kip7UXbLUwIoIln+pcYkQonpRy6dKLyfLKzoKXZiNZEv/78JLfVL
GMsj1uMoEecwAvIQGxy25b/0AAj7MX2gV+dvQ7TrdBFnD0KCoUYy8DXnvHkFdQC7
o2O5o1WukEhssN0HNTGoTM/AB+zwt2Q6qRkipCxJjOLPVzerhCAjj1XMtUlPdefx
iUnLrtS5979/RT6keFus6vmRvj/tq9X1HeEZLJmHuGm1xWtaNK1ha/ZxZqUUG8aZ
yygQCYdCVyIOKERrPJ44rO3pKvzPWUW62SyvSyCsPorriG5yQk3DvVPC9LmkHrMR
/XswwU2/JJ0oN/+uAVwma/GXvNyXiXaKvxqn/WzpijHAfdnA+FvL4CAENp8h6Iie
IijQLHHq1i+ClVcEY+Yj5/2OhORIeNBpEEul05c7L1BP6+KXPHfHr4KFrGNcSEYd
qcROGOxjiJdW+YRSFgjTponlkRGO+GtRh/1ycjGccB9XnwJ/mbMu8ZPIo5LATr9k
bSi3VXCK7TwvYNyaGO73NjX9oSyuX/xmJWYuxE4X+KrpQuYf5LKsXzqjiQH8212d
bFtqrU+YEHt1ssydba0UwyykqHYD6WPKd55WluAi61Blh5DjnMLX3YyFo0XynlSn
2hmG2JK9s+4ZDtFjyi+cGtEIZ5DYsguncpf/hHAh953ivk2dZn+Y6PTkznO1/bdW
SvZbvSfvWKTe3gRlp/qYO0qIqojRj/6LISpmanEQv4xYevmTkrxTv0o+XoEjkfb7
X7Lt/scqtq4EHcOSet+0rSG2ZYP3AysGW2MGzd2rGHY0K5gAtiNF1Jk3slt257z1
lnOjyGlDJa5EDvJZuw8P5vMxaDwWf+ASlA0AAzSoNSxkGkdznqCzdPXsUf2XFGbc
BfEcLyjAWOvuJJKID7bUNOZsOR8LedOSjuXV1l8qnGYK9DiknqVQ4MLEY/+raJIu
TGaDul+X0xm3HDxRwV8xSws8VLEm/I5WFOCYe1LezZviI4wB3fONbB6KPe0bGDvb
PudUAWhJ4GfeYm9GArfbysEhzSpopdFneiCl33kD7gneYWpYBIMwNQzSwrea7djB
BA0OYBX5zORH0k6mVhMtEpNzx9N6bN9re6C+UTpgkz5ScRz2Vwj0SqFj3wWPl/Go
fBZc4jIHXRImnTSA4WWh8+Hly0CNxQNTumugBpx47WIGT923UurbmbevI9Q6xXBB
YmDt3jDK2HA/T5PFsU39IPOBDrEd4VGNF3glfAwh7hs518DvYPtwaQIPfeQIgla1
GHrgEtcOVuAI2/cR/meriaGB+Cxujj8cc02/XPaJNcdZTD+zVsv6vIwuTrJUmxVi
pVmX3FCiXjDN9WjnC/MxApbuA9YlIn775F+w8t5GGtNYCcq2RHpqODmqM81TsACm
o7NBmOT7pp2UVJyV0huRPbGFxhWHqqAH0L7lM20dZv07BhMSUFnn0wmsedGYw5hC
ruUVvOLB0J4Xz1zcCA4/vzbmAmIoo/QYctEmJLqLbwud0DuiIhtxuT9nBgsAXdon
ZSt+tna3wleb4SjIwJFMUjRVIW7aYo/9iqTXzJ8b2329a/Do0eyTguIk6TMoLUvM
gyx7RXcjaPngDqZmzII3CQ4I+j4nQSbjcZMnLynpUd61etQ3vuSoXD/Gr1FlCYtI
fCuphKeJvDchFTbFL33QdY4XUssb8ipO3dQOTOWA8ypuNix5gUW0CXxjmSEaTxid
D6kyysY+vzO9ok+156O+/eWfe7y/D6CT6beC9e0lViPNsMsBTnDjWgNqKQ1LaDxx
n1BdmIkqlhF6zAcgAhIKvbHL2wHtrkhUZD/z1ZgIPs8aWsfVtDbgBkDBdMeFM74V
dBM3SuhQmKarVZNXr9XJ6iFEXDBH5Ts6FICeUwO3NNhrL9s3YjLg9+syGZog3cNR
oU1ZsbF5jYJ1eS95FjBccJ6BuAULjqvXXVxBTg7Q5e23vZ1Mgo/B5ZkbKbKMDS5v
/QqMn82XOf+vYpo3NHaRb3y6kP082mxeosnMCOCIH33iU7QtMg2NjAE+oshjyBmA
2I86CCQFQjKR+3/mo+w1inI4Xe7AhQFTolSPidti7lztzel9cnJi6UKhH5i7qPu0
BwIHgTJ78O3JTFXZIHkH/RTLglFhR6oh7eYY+XgsQqxPO2R6icRG4HBQB6KVynam
u6qoV24yWXf0sP4ZujZKeZ1iAyWknHBh5SlaOc5hmtBQg+cbVYPc1tDL4LA5WOdw
9WmE+K6Ydgy+KNqFITtl8HskHx8SOu53SiBGXcDNCvJBgjPmdi3CAs0zyIf/ApVd
PvcQrfhQPfaGLZXH8YHE6QbJz+M9xamXJCxW4RgNNtVQWE8uVF6qbbvzj65isKqZ
ys3jk+8qbOd0ova4CCOucBE1S0Cx+VTOR2KP3SP4MGuQoCtgYy9BBPK3bZHkDdp+
KbsJap9o9eJaOuQG669IaEtS0kTFKJXNX+CUH//BteGxRaoRB+KzsbQZskVj2OqZ
sPL5CRCG6C002idaTI65IRYtkSUuWsFkDULcdiTgB2eOWq0tP0Uq7dvLI8DOp8D9
tJ1uRc/b8eoJyrNKDpAyYe4ZdjEyf+Q8CUZMo18+pW6x0jTeOcFS7Kp+mOTzLzkt
XZ32t7utdFCI8hW6CHes+gLT87hAUaaBagebfY8BWoHizurNWhNeVz5mlgGdv6NM
dWFxa1oxnG3SfAgFCC64zlUAU9fjs53Y3ME2qFM6mpfrBdhQjpWijnQizHwrgQVO
/X16UM/90ee96rM5ZfLIbRT0liGPcwZ5F5HxUffvv9em0lb5hJf0qoMYpwm/x2kJ
dK5P8wiLIC5Pjr06H0ftH4GjM9Cmv9+aLsE5CM4TWIIIb0SOfc5lNUbPGGqX8ODs
InM1n3Q5q9zviTdEXFQPUROinHKmsk5j6um1Rr1r8C3QSHxRcc9vqRBbGjwtPVNU
hxchP4nxNLQxi1aw/ldtLgfB4ytIG0zMA+qx0cwtdYQB5G0zh55cHRKNJlRkGvel
oFpiTCDVmUFWSCTIQ3B/TsycPUpCt2Fylk/wD1EGw/ReH6lxDy/cGms0mHDTyTTF
2uLqE+aBWru09MK8hIM3uXzJ2RXTgJ2b9UDqf/mLpqRuP1kRtgfMaWyCTgj9EuCs
35F2HN1axcO1KVNxhBMMLDvbydB1MK7DypAy83CxGlm3qvqe5n0UBXJU/ahkNm/e
k34T+kpMhySjUrtYQHRTwLTc0Z9/rDYd+EGVI5rX+d9yReNozFbbGxX5ScqYg/4C
+X2dRweuRLHSukinpWj/a65hD7VKTQAW25Cn0c20yKaft50jHXTwmRfNL9JsblQm
K/QaS1Kob8NuJ+9kagNQDm5hTMyqFEH/Ypb9uODzKFlEtcMrG0269xth2m3UE1VS
/7J2zN+7IxfQ59/8HLFfZZQ2DE1UfBQ1n70v0z9JjfhjPSIphvEJCcTfb9RV03h0
JBLw8sCTbmZCFSSo1DR+b+nEZgFxg/OxuT2GbTekqDEXTqeWIoUmq3PowQlg/o0q
oEeZCdlLfHSJT61hLrOpQtDqyBtag5toOqujG38n331WMaR7Z7kQJqyY4Oug+ITK
dxECWP04oFL42GqpREDUDjOImifWooQT8z+VeOOcMF1Wk26O4fPWPdnykiWOLcWV
vI3P8o72eGudZMgpd9QJJRIDtCWXP0hf8LoyzAagdPBQHyeLMUVQjjI/kIVpvMoy
D5+blyT8l617SWLuQP4jh5UEEV1o64rHZUtIdOKqtoNI325NgAK1p8Zg6sglgHFS
aF8d8nWpK+WdTmfajUPJTOwr11lJY4IS9SZ6/Cgzbdi09Q8Pp0tkc5T9CmRXZNiz
GV3clhudAmfJGxYxExPxMLvUMaEzFf4DqEm5xidMtj9pw831RpzjHc3JgyqFglzB
/Fv0aAgolXcjc1n6huQP6anJz0fjDXmkFNdH6tbgxiFnSbR5/WZaIeSe4J/pDBFi
Bkn3GyFmUIaWaOAJBKytLmLt+xIHqMte2jRAUPkqOB0aeiAfEv4gvRhQPY7OtI4n
H26jZHVXfPvNvaMg8eFCbEnhnE04OiwwFknXshwppkseBIIsw59rxXxAlFHgNLwu
UzHr/jQ1+r7E2v70r71ARiDueY73AsIrZP9hkhV2PHlUzXXVr86sLmKFVT5dvQps
hpGWoF2bquhpS4W2IeIiGo7i0KiYssWK2u3Yzvnlaw7Dz1FiiqAwh0ys/QvZkvKW
b7BnBweFnLshvv5nBGqp2ri3oMFZxoGNcyFtqss/U/MuJff/sFpvPJweyrw7sdBu
8gAAsNrV8osB9yX2tTefzCCeJ7YXj9Hh0c1x3q1vM7ykVmn7SZcRP4OmCclojGzC
PYd8qFX/t0LlUdnCFBQg/CPklJfq3BJH/p/BbAzpodpN2vN9kkj9o83PAXf1Fouk
Xe6SFo3q0mvyg3VrzHp/n90YUGX/gz97d/IfBUl8u4Tkn3anvtYY8F5xlDiBmY/F
q1cgSyFpkbMY6AuOjRxpsQZotogmI5lqupUscgXqN/6kj2wdwms86wbnI7QXhazJ
OCf2Eqy5WoFD1ed3ZGLTQ9DYiS926dflt1p2Yj9hITIjLiVvKube/wpne8tmFGTq
fazXLftkgxrsaPAAc0/pSYhvobP82/RPV1E7LPnE92RgoZAfwyhFeMrhxB3HqDhM
DOpxpKrdUJJdlG1RZQgI/6b2Bb6ie8ORxYOdjzKclQQ/r3B6JK8G7OkocM6XXuac
87ApXax98YsrxS6FQ+uZOySd/P1zfCCJ7GQk+S7i5Vd3/V4XmkGHLiT2vuKk24eN
t7yo+jfqgaHP50LcW62gZcRQSOLRh2hWqnO3ezaqmOMguk7FecK+UfZ2F/gyp4FU
lH1ddl3pnNwigfLaOTUAJozSnocSCzoIzc4ych1p7OdgWW7fbu/Sl62VsOSxPi5B
BVTO2KOPbJXkMfv3GnIZGWF/Fp+P4ysR+aedp50Y7hD1TnZU8hEqmV6PIxUmjJTd
4NBL6M70Ya8JipNJ3ugfhy+/UvAq4vtHMRuyNtj54X3Uz1wUC2KwrIszSRc07ne6
Fh/pe4apF7LGsDPvFiEl/2DVtBXIF7XI1OGErez5qOjW08XyRbxZjT8SIO8x6AML
5lmqBm5kKLE6Ppieni42WiDAinslhkEuhmuol8IcuiMuhxFFrE/oTMsMkTRKIKBt
8pWXMJK3DerpHJoMdzizOiE7Q0C4gLyT4q3EivM4scO4pHtSSNdMZUOQn4q8LpII
v7NlQN2Gi+zT+t8GHM+ppA+WRfwCQyXWpVs1zb8DzTVLNEaNw9p6886raF7vuUXg
KAFCRHgrxrVBWqSznh12bmGFoeRygudNz0Y95/t2j3l8QF8/Ee8GrnpWQViy3En+
x6iDHvuhQBuHjo+tzoyTNvB809DU4gF30gXzyOzvRetn2K2ePKl+pUmKCN0lvke1
EEvfvbwh349oT1jOOomttu2MVeJ75PfUcibfXkIUq3KWn+30XD/FCl+ScVrk/1yG
tVTXRYDOlLj7k5fhMJzPWKD0xAc6CyZkWLBY001W+UQd2MPzSMKMk/CEZbdDtuM9
ZDvDawfr5fQM/PzgjwuonJ1moyBLbN0DB5iNA3ZKIjl7QFf4o8DRMKjslatv4Hjz
4ExlXLTMIob446yaQFY/H8rTprjMoxJCktXJI4PUN/aaUHUrEGR5wLnKlcYtv5tt
mAjCaJPnHrVwMY2Ywulm0d/1MeL/PJBMvPIV3ebZtMRZIbGv6oXq1wCsNTvwitG9
acGwP2Rca8Qxxe0sKTJ0APsLQqjzAOiX4D6CYBTEaFveesiHEAM7SKFC6XJRWgkN
ruKVEcgt93C4xHDlA37PKvpsliNPYic5cbU4IBAW95oFzFcrzrSQVcgruLMHxnO1
MNk9Bq55f2lFffzJ2wd6/nqnxDLplXPQR/MUHv0nlnTypqsIpCFHt4kI1Y6W7+xa
yk8WEjwEXbs/AaVykIIDQ4RYCJa5CPdT+06sPY+RSd0yuKDm4aBgyBjCY3kw6g/f
UZTQmfHLX0bORlBUdt1ZVCJVaO4KEJh/WWB3y/UrRq0Hky5bGDvAY5EtwXxNN1OF
xoqnH9e7af64Wj2VmyOdPQLPlhZn6gesDaoiY9d9EZbeqotWIQjI07xNM2oj1LKu
zX6Jq0SdMM7EuJ9hMWNDyIj2TxcBprYcOoS6P8dR5OSWuBjBGS0OUL0K2I8Qbq1Q
+2ZS0+Dkd4iZ7Ypk59mqDSDntQJOLwB6vUglNC1rcy5FaM4waK49yWZxB+P8V2Tc
WIuzTNvAKVqpuFn4KQIh/JUczmMWxgTxDO/X5NX8sfQj5j/16pkuE3v9NnPvqpCJ
T2m2U00Mypf7HxOdPK4676XLnJmdZHzfvEYATEamvhpoeNUyVOW9iF/HwjVyd56G
TNKN3iFLcjkfv7ABwyc7bnGn4bqLksWxBXyFP/uNF974ptSFfHhNDwmNf4wtbLsp
7Bc9ZQqZ9jXpCoXA209EhCctQfpQrBjh1qa0lRO6sSklaDoRTfDQSW3Gijk0gosZ
RLLofh/TxYe2u5jP63GnPFb9y2ylJiuVYICKx4yR9aJgXILKIZ8lou/Pg+qpuB1a
z6OlxFpYMJUqKYl+XADl7Hytme6ELXK0jD+zsJlBgqMmPr4WvXn5+8bpMH6tN9CT
bGlwqV3cerk44yc5GlYUhpfVutgBFdRqZPxN7R5EEDs9XWCCk+VH+GLhjk5ABRso
LHqNMmEjqmVztKB5HBPkv+lATiP6MN03uHy4FxmloWSUu5LRtZ5mzX1C6+OtG7rM
17vWS2ztCoKnBNHyAkC/0XIaj9AXZM61BhnD6rUJmcEHbzq2NbKHpmWDrwf3u2j4
VQqtjP43R47uO8pLosNE4uPUTdtjWl8R05bqlMHKCK1MC7q7RbE3Sby/BYmvODf/
KoaUqkx8h/JT2Im77NqRZRf3gqPkJg4B5xwukvjCIiA8bxzmHliLixFZrFA0kcT8
oubGBKLWWhpFykQPNuhUO5NXBkDYxjfoCddl+32x+AT0yCGkGXXkUjH/qGAVRwYm
zRuh3mjo3VnI7KnreYaw2D7yldVemOvabqvtYly74NJYtEtm45bX9djXj9HrqkGC
lCyLR9vEDC9sXtXZbY9C+eigUGfjfLiysUAOOp/Fkuj0+pfZjVjfZsoDnrrV1CtQ
jJdcZwb1UuDtcIygIag8Ru4+IYtWSe/eOLM0wyU2Wp8G+/9QibytxrKEAgah1xnd
PZkeLk3sTdstzn/ChVDtTWod3y8j7IXqukXgucZWNZ4Tcu3V/jy0qmI0MMtQ4/0j
RCz0lybJ46YBp9DthsswPJSm1jIAGN5rsNfxnoWc3zPWIjn2ODd0NLUcOVSW4Nj5
jnXta5CalulL6pNPMZa6doeY4Ug/1aHeN5sI4fTyly1BjEHq3bkpYZALUbLwIWwI
hX7VBL7px0CIhB4zxGbyZiIobkSgvHJAIrHa5Fn0tEpNgSitjg6BoSmGp+fKIKpV
cWWt4IP27mC+51GE0Ll5IZoHBtTAZ6lmeGZi9qwp8n1b7bL7KWdcPjb82tu/mM0U
TeaMWAogw2+tYgUMokfs+gAxoUnqHKcosIVl/8ztb+Wzv9J2DwYsSkwU8kyFNF7Q
Qy6WEXA3QOj4d23Jb9e7qhvCnMmpW5MoU3h2on5NiDAL1HkWJn3wEws4mq1VxvF1
NEUxQPQLbJi83gf6gsJKXJbbHHK4BoLnBn6G61/4USRUokmz88RzbOsqp67ZZVzk
65btVSxgPr2cuOxs2MK1A+9STr6zxBfnM3dNHhlbQm/cU922Bqr4BxaEKkspoowH
uCDnc5iMHXeb7gQhtIaMjjz8nvjuEOfoHuon+VsTRHgGdAFLRw4ztI5UroSfPlNB
sjqlyEJ+po+ubrd1li8I+oXKymgGm6LdaKFvM34lKZ620PKBPEtxocr38BAdoejT
hvodaPjmt597cgTWCKvD5lpQLZR7ekYfAJ+KVX1yo9cBLa7iisaB+Mbigp+z2oSV
/Z9cAJvIdA2Glwa50oIBubCCTRz8RFvI4kzs36ZNkijLIwKuwdFDASmEh3XwJwTD
HwowlC88ITz91C2WwQavDkSdCbLyX0xBo70vrH9DHaawo+F5Inn7teWtGUooK4A/
aqVdVt/MTivl2m8a3waSDIvrpu1/Fdf4DzatxwcizBt2MF9vniFJrpyUhQLEPG2y
ZHWFV+0x708YBlGD+6OYV8GKZp5QSXqC1YeIqfwGQ1Fvq9kQM8LiEIkTgst2fAh9
N0WBrHauHt7hqPhdmRU0r9YXC54MOGYoNDA6x2a31R2uumer/Cvv4XlDNqD8+wOy
aF5LoNcrPnZlrL6WKQbp8BiUwzF7ey8pvPGe9Vf5Sx+f0ez8Q3FFCvqJrj6tOJ29
f2ZxHtGy08/B6zvpaw1sanpr9moWBjV/VQ/lN7swR9cn9VJMChkqaaZD9aWstFHc
hXMDsHIrASDKXQHqa5WzA406rB8TLFOeht3hwO4WSENgcUJzCMFZvQi86bK3RHIy
45yzbcsu1jVXGxFKjiASZ3Ounl+spzlsi5S08lWx7te0VS/Fm1ut2IGdjNDmXmgx
lom+kjJtjj3GPlSqu0ZILfnlPtXqfDDufP2aJZS4PMKPjv/21AT9gi7RU3+Xlbbm
2Mf9DU7C1NdkOORl06n1JafktuVvSFHV21IIyjLVMYC9JisNevdT3n76kwNcy+8n
MwaqClO81OmU7u3hkYb1fDIANB1AIiaoSPQQzoY/m2j3omCeXkksnIhlZtbjBQsI
A8LW8ntWAzE7O96TLAkXiuUonjfj99jSLYs/gozwVHjkEh6k+kDPA4Z2+L18sYuA
bnSn+ykf3n5j2Z02tRUrVqThGphQltKRRwO36rxbp3KFDs44xPzKdACfZFicaAs+
o1zKTF5INscI0H91wbTMOWNEL35a6d6ZrhLQcAawj/rTkBkbiWyLwVBRGmGPv/hG
0FkY3SQzFLgzB/XtDCvfEhx9aQl5QkGS3kUgXVgjZ15jMmVeLGKQU+Es/jN+TeLX
u4TEP3NxgUdJLPiSYmEN58jDgZkWPOkvC7qkAMBhuSheZn5D3ogC2dlcpOi7tp0+
qmWJrxLbpMh85MowtR7yEo/Z2+1wy5nfS1hm6wvGbgBwW2R6w1gN0wz2bDdAa9mH
MCOsouNwSsfOEXowJpg1B7uqlJDOwUvizGhQqeAwvHcB5XAkSrsGHfbTaOe4SyFz
buSCo6m4aM2NEHzenZa7XAZoDX3AzUg7gsS381CiuwS7p+LOXeLnRNnOxFvwAESt
2s7uJKcnlQ7VDjjg6h+4oNeceJAIyYJmmAR2JJ3q+BzEG5VBAbFoDf5ronTkLtDP
Yu4z1P/nIlrqmmhJNY1XEcdPxzisi+E0T9EuskwPvu2h3I/kPLDBStq/LDfQfBOX
bQfhRt1QV4sBCBSJUm++iVmeeFPQ5oX6xTa8ILmcBFJkdZl9ZSN+svN4onY+zdHH
Xu+Vrs475kTR0Oe0aBuq9lVaXn5Vv6Dbw8Uj+oE/1dxpFdFrdXKTetlo9Thnpj7C
chXtrLKD3NqCKWIZBCg6e6ir8CuvWqSVeESoyYhIXEzY0LSAx5ZA81xjSH1b5e0n
726SjDMqT1AhOF1nec5WolvJ3wVw4zYLOOa3PJmcw2gQBcfmtSgsRBtyoFxEoVmT
neqoMHcQE9ZTipAa3mAEcpbp5PcPCPIXKtfzKdeg7qXUMxrk8O6SLdadTW4xPH3Y
atVittNvzAhQ2hHmSnUzGuYcvdPDxjXGYdCgj2QXODnTXUmTeMcQmGc5gUHCQ20Z
PfhscFYuVZG65fcPztYwW6GbVztFuEsaFJuyfVejfVmQQADKjogfVfEGkx0uazt7
p/8LQ1Uw9idxEAPJCo0C24NAF2rzCxIxSyZaIzmuQ1cp55ptNGDdUL5FIoK6NeNN
aVlknca6pCK5rY32kbAWISw44Ygc4GQWccLq+fXXDK9WRMtcxSiIHxuVhulNWZy2
AyQNrVoO2w+OF18VCSqp/d4Dt+dUFC/ivHZ751w3VS2KcHEkLSYNXwvdh8lfXJji
vgFbZJj4RW1j+x+pZMt2TmJdS83n+kLe2LCKoleev9mZlApi9ktP6HlCLZ6mK5AS
lxJQrXPhJCRNfKE2TpjI/iSn9ziVD2KtToBvToUFE52lXVTInmjYI2glBxrETqkU
owBkqsnnnvMnrIFKLBZ88Y4T4+SSJT+o5xnPKr7fDmRrHnkn/WpTFS6DPVgcWfaU
J4KsmkyKWWIzk/cy+3hUcKsUq5uXl68Qn4SVgtNKMMTgKKooZ0BPh0zpx5e53uAZ
uvFy/SmkagGCZDu3DeMK/UitRJfw8A/j+TxeRpkcp7a/FafhzbhODTVe8+3LS2bb
ZcLMcIRzPLJdxSNFxB/qiU1Wed+MqsjBNoO80kBAJf+W64lhXhZI62/rIpnDfSG8
XXh1qezRlhZh5AgI5n9D66vTRevA8LZFFGmKn0auObZNBkAv0LzCfmCBhhaH5sVJ
CL4r0xeg+Zp6eQQWx8WntvsfbAVQDH9oTXCD7brO5DlSnExsQyQRPE6w4UOfvXM0
lQ23LGoaGWIS+pX87HLrkUacFl8ujMk/jTGCMD4kof9+4jQb7UKcnoayYzutGvuL
RuL6K+M3a1KcZGqYX/+Dyyn1UMGpFY5TVnv181euxv2y8pgVZo5hfiefVnqIXWPD
mFtWKpWHGk0gKKO4Emg96DN4vBzOAXOJWUdvzgK8aU64PhcB0353NsEWWbmYyB86
j3JFBeWxD+D96ZD7csBuQp9Tc0HchzxTvhiuoJK9rLdDg11rIGGLmbXmgOwJkCQN
uIuip6oOt9Vn7I0NO9vMz51nb424PPYjed+4gbEeHkefTIik8RCOHM6bz/dlonEe
ERpg3MqcLgv6twqKU9nGVAPmVjJlC9rP1lMLjj6yAFFbBEaNeLTdaPBlR9DC7Nj7
8d1Rwxu2Q8v9wQ10SOWSPEkrVHpEtt9Dnw3T0HUA26NbkfiViiIihxUu7/qYtXSd
zDXpwiWXkUbsaYbDitqNq+/sHDbx1H4fUvzgxjX8XbK+/eRzBclhd/c3DOzalu+Z
YUbPOrzCDR/HALe4TxrhSWo+ugPR03Z3pgN1BYLD9spQZ23/UlMrDnvZiBEQM7r1
0ge0n1lPWyq3G1+AAwCRKeFJMwGvS3AwsfH2PUlAYr8acJWMnLxHtIlnJZ9gVETV
eDA8A0n0mXKmTt2kmdvHEzROl2xOi2wrOW9WdNy5t3eZrHLUK0sJJE5j9JlG3OGE
w7kUj1puKNvopyzoTtgW/njEGO9kCyerGRC0tyi6qc7Vz4cvXy7JMJD9Ah4uS5r1
+oQ32bOdsEo8dhaXPlNKL7EU06Wn21GqvuXxopr/hqYTv91aCGw29BgFEB36xSew
BsU211DedcbL4QRzmuAidP/TC0i2dXTjGmzX81a0NdTuvQgk3+fzQRnvyKjnbyYH
Wdh5FJXzAAMhzP+7l5JNz9cWyCcida6UXBbwc++ZW2pf9Npr2pIYsD2DvSxTJsoG
FbX+ze017XlpkY+/PufT+jQxsSgJZXG87ljUTOcP1utbQ2oQ1beTHYRZwgCfl2eI
tYJYid4OvzntwO7XsJddi1wmsa27m67RflSJc9udRZrsK+l71JhMgCXor7e16EQG
8oxwqQMVv7j22HEA02WinoQsEY7pVrTcM0EjttfKrkhUaQlN2NLpyfKhEadtkXGy
CDL6ZK3jpGnEF0QwvGUBtC06Ci8YAjIKhn2ubGx6xOdmtCRspTlfPrYEpgbR/Hwq
Maru7geJYGiBDSszfZQO8motTAbJauURD95L2WiVJ7aGigXyLSHIcZGZfFQ6109f
sTUQHwTWUVhYT8u1XMcjvLBM5TXrmuE9kqYS3GoWYBh8EHzv8Ka143ZvCJpUNKfj
cqMMyC+rtAw0Ir4zBPF/9xw2Oc/CVuFaABpV7SzuuR+XBoO3RB8iXELP4neNQ7lM
d8gwGFIeQn4y+bJMjYA7lYiPhv6UJYKWQ3L2ccVEfNPKGxlhpSLV1p2Uct8EU5DZ
U1XpCsrKJMZ2BY6p4L5qnOJNgS1oAgccieh4biol0HLmXL+NMUikaaQYYopLwRIf
/9Hxa6P6W9RRrP5kRzWuSYdaMXXE5O/xYebsqNcKuWCcSllIZYVU9JVv20vCgnuV
1H9xsKPBrx69g5qUa01mZVx7HSak1SNv+05CSEfOa7fDNCstt68mQHH2xsGo4/y6
2mn1xGHh1y4ErHqk1WNd/Jhu7tE/mekQDuSt0twsxptcpt+vybdsb1kfa5z8s1zX
Ww8cy5R/HmzAGc5VU3bYoVO1nnDpHTLtsXUGp7XDkASc1QamWS3KuGtkvfLuB74K
fISyAsUZSTKfuwXZvLExyhbiG7OxHSU5Un7Eg1TswDq4JPOUkamXt65ezIsI0eyJ
kC1Ef07YRqvAVwRoTfy17jFcItoFpYifdRbgIcHVoI1qUpzq1TkzfE5MFcqjSdCR
dvq8j0pX5yGlRJnfzyaw6M0O4bUBQdKiSR1MOQmtl0uerAkatckgnfy5E+F1kUjI
/8EVHFg5gTCNLazhS7UGord0rhJX8nTQuhQ5+X8m2uv6MqrvNk4b+FLM9EgHnn2t
2BfUyvGwGEYOneLHXyAKL+mwAn+6jVZFlihhou5eUYAImwGrsn7Q2u3FTuk8XnIw
5VTnheLT5Rb6mA5lgr0doOC1kQkusLlk0KPiJDkU120yLkptrKYnwi3pbAj0qt6B
OT0ZPFmvOP40y+wBbnGlTtVx9o7nrXYlih7ZMkVZYkI382b98CGnT1CFB6AHTXgy
D48xAtcgOqJ+HcKpLMCFSBjEQHtSlJFa83vzDTVJ23DX2uKbIUdCTFPvO3Ol3E4n
9ivUc6cCRFpXi1o01XoF40ZtZd8RrT/u8rqKUKFr8Iavb+CM8bxikNHjMWcZyJSC
R+zVMdSY2wOCF7sFpcHKhiLJ8tfvXGs7LW6+9val8CQib58O9YKe6McfJ0FEqi/u
4nWsh++GBTzM+Pe9Tb+aB8bJbvOvl+gWSiv/+gnqBy3beE0A+ArRcgPzcWBH+ofh
9C+L+NKRDQX7IBHOUxp+p9cwvrwX0fMFYWC8HHuGEJzc6NpZp8yvg6JW7WTkgOGE
nTU5dIprFF6pMw3pm6dkClBiLBmWmaulkXnvAFVvjBbGciNLPskgN3IEriiCQWq1
8q954PDAv2cFZCs52b2npoxG9XE7VJ4djOn9mvK5Io21qpFH9clIpEYEhaZTP9XX
YMFnYW2NjmqOtzDHiUqcqisecFXY98qyN8ihgSx577HOaP6CX6wKCZ13UhRfiy58
2aTMhI2FKQvZlYgXt18+krwAQPlo8k44j8V/Tu64heyV4w+XeNNPqSmxTI1OcoOX
MkwzBjY7oaa94Um842COWWU7KjkBy8tBh39zOlhgjRPv3J3qTnkMUkqam3NS35U4
AUvRQFPc3iEMZfUmXTSGuYjb0eoFoDzxVg6dFO+VwsEJqB7semLxqSnxbXg4j0Zc
hH6D9QiGkUUQojHHhX9VAFCN6DN3xA2rEz4u0SQkbEst52yctGeX0nHadmcXJG8S
6tCjDNJEHMKZJNb/YcmEL/7ZrOg3FnoRrUlcfM/0vaMEJWHCA/EoZdhNH9V65eqC
uv5sXx5hpS+lFUa4C5mA4OPKpceFFgj2kT1bFrI95tgF17uyOcB9dAF3B6bRUtia
0+WxDDc1VMxKlgTxfwydNGN+aLXY0b5UOtICv4Txvy8F3Um/OaVsjCn4O0r7Dc0O
8VQ8GhqgB+XcRKiaMjoZ2MpCqOkPSks9Fu0qNTm6KqB4FZ4on3Bj8koTahaJpIpV
urC8bTakQCVCe0UxcUwiizXsOCDPqPEx7qGtkzvtb+0P+LK7GLMTyuy0nIBoNna5
WFkJTiSExWD/Oi83Q+cpwrHMOovpSuaJtXav8pvMiRG3gftIqbw1+0IYKH6tzMS2
DncO9cMev37g5z5ocVm6euhIiE/qsO07eIiX35lnsLOSNomE4laigtDbcJ5VFErV
mxdg3eCdlqvWQAuPkMl21byGhzACfqtzPSEI/dtMRSB78vS5oN3G3l/z/fS8v6xz
aOtd7q0UfcBX6z+v79kGdu1DuRgjIzrrcgWuuOvf/s8LvCTKWVyNN+mBC0it9vaT
vWB9lnNiy7aH3EevTS1Hj1pdNstzglLhHAiAW/Ma9niM9LO0gCUj25uK3sp3mWqQ
tAsn3uNdgCATb41F9IjBGre3afEyfro/0uCje/Q7BN7b2dS2qk44sDJvAlUTPaRp
hufetiqICs8RaGIIp1bfjyQsiLEn7D7P7wKQJkdYRMUbyOIwlXW/HN9lltuOK3Js
qO/Pw8cXFoKpK92gktDLZX2cb22vEZLKyHvIwAW67SIZEhg9h59xrdo4t1PHQRwc
864JkXvPwhxF65A0OQyqNgr2JiQSvXPc6eoyWCCUhzT0BNjaHpxjTeYrkGzEg4BJ
7njiGNuh7s+mOfZHcJbjiGb94HjUHZs3bnebDt8wKBvxlA+7rLeEbQN8c/nzSOMU
Jcr4tHznGzfXGkHHyr2D8qS6LkYsdfT9iler8V1NezGc4GXuW9Jitzo3wikD35vd
B9G8z9M4AdQnfx7pS7O/ynyopO4m+DDr7QTSqJ0yVaZI+0qVMj9hswb0TY4wq4d/
KX/RtcF2djyiR077KcyvZNFxRQTsJKdzHpxIdyPawtUMmfMVaKEJOaKnYyV1oe7b
5n7GYQ7R9FJQnqyKgd+c7z9uP5Cg/O7hXNPvTmh4ICj/HVlkq7UBV9MZjIu7dJ2M
33L8aBWAL8kIToYGq0/z80l3dzr1LY/puvxin0LG+3coXJi5nG45TkeUplCzVs0m
JrJDKCx773joZ00npj7Nq0a6/1DQk7+XTtWswOceT7dmObiUCXWWzKR+h3wIG34u
qtyka/1Q0l/8DmHXdNo/6ABTH0qSG28GBmAijWLUOErnRrEUwOGiuScc8jirgkWn
8NW6ijeBIsdZqXmHeaohHzVSPSLNipzQwPIoLh4yI85uT6GZ+xDYNX2m+USVeSF+
mdD+43Yx/8EGor58Dna3yvrxecEujQRebu1e/r/p9BqRoPNRytVCuprvDdpoS4c7
TVyX9CqVeoxkiKD76VyVghvoQawvjyplabCJ3kRnLzHMVCPTuKeBUlcKdu3IUjpc
3yvCpXKR2kPPptuA8LVG62l1pRMGO+z+7m2y/szveYkcb9wn43GSdZlNrXX/YZkX
q8QYhxBeV1gMykEjPpwkc4ruX38XzYlJr/zjyxVA3ZaRZ3+MWhMVTc3rWS19KiNK
qdF4j66+Pluzhr4r7lsU8E2juqQ42Ze8wczhipi+wY42maP49bA0GtpwGzz8Z6F2
D721gxFQHaBDOf5j3erwLOJW4Nn6wjGS8AOYU3sJu5Kyb+gF1SNXCYXYuHBSI8Li
PpJb7++61oP55T31QqavMAKwm0sTwg0rKCKV6yHSRzAVqj+EoShXu8m8vlfKU57+
RrVJgUkHQC3s0tBdbHJRTLJDZ83ARJ95llguZcUs+Wvpu0Ng3Fxdi/yggAan8dGI
RPAXmUhKnbbHuzZpFyLKpas+MPifAHwFVDJZXWxmn4ElWpPL0lwaIDMe6SXAoPC5
IG26XVrKl3jkbDzVMreN9z1zQKrFqKzmyVUR/IK1PwHKALuiWwmwBXCaprE+IhCm
ZfIVIvvwftNfXKLE+MkOb4W3DW2O/ActYnF/+XqVbXdeYXkUepk0qAATlqM+zYyY
8jBlOQ7SQlZ4j5NXw1wvFbq9B3ESkvFWlDgqDCb3TDNLxAVLgfZrPo+43kyc3BIX
IhpkZow752FpJn0FdsuDvOLK+bg5ize69YRYsp701Drk+dOlt+8h5ze1wgIgXjmI
BW//H2UnQQOBSUJ2CDrHX0xopslp7ZIfY9tuKd2bmgDZZldfOpsVasmo2Lx31AZW
2aAAdM5+YLZwLp2yEn3GWs4fePqJ4pDfXK6PbBqqqF25rjmoZeeuYI/sj8/Kp6jK
eMSZ8+v5tJW3iPcSc0ZdrPq5BmG8Odac06TqskmowhX6vAC5p91UOBeZt8rpI541
ETBgLO4VraLUA6amwOT0Yd8db0DTB3B9ZppIDQAqpf9+hl7VXiQTcAcYstLI65/E
iYbsxwCMwPYolM+Wyf7/z4EVdqwU0OSu6mQZD55NOWg/PGN3gkMQyxgAbPyIDs5q
mDoXlPTFlIBrWo0GnGjxQB4510AkgPRcQ65ULcN78nMJwe5PrW3NGq7SxTKwUs8I
Cgu9+UC71W1kPqQDy4nxjP0JNcLGZdInh5Kwx2iN/WQGjAO9O7uVycVjG1AK4GL2
L5f39b8niGgXadZeH5Tm9NHn+UoWEzWj0cyEUPJu4MJendpbkhDdapJf+vWU7I5S
oGDUPzURO66icJKrIO4ADS298avWgDQ5Bs/tlF2dCgBS4zdbPtc0dV7RYzpfxubt
jLyvoZa5+m3ZT1exAKwbIDytYF0GKmzkzzX0RHr8lViHIxvPu8+VferGB8uOX+Sx
frj+nDr5O7f79vwqg5CSyPY72D94coqUCZHDMDx21QKe4mmDi1ibPMnkmz51pK63
HCgXcam5cHFQZ7ISk3G1MH2DGZntmUqLEbe4BDk11pgteBnGNLG4n24W7N+n9/Od
2Td+VyxibgmgPYESBldgP7a4xN7pkV6n++IbCCWzxBktSXgozcJAjweHMRFCZfZe
gYqq+j+O4JuWS2hlGWtMVFseZp7USqGOceEX+QsAq/8fliIzoHqrhXLK9oh6pfcu
7y1RCsyAtzQUZ3JJZ92MLKoC5ytrbxPYbJ7MQQLpOovP5vCFPhER0FTjZZFH9Iww
KoMnEdcl5tmxlua2+LwuYNvOlGqJ8QfGPf1f8CYsqALnDxQh3DS5NWWrwb/0pQ2+
vwd/5fhVPStgGBKyuikzBVZHk7U0Ec3zQKPh2Y3VlPFA4gW9kZxYZEA/UxM3P4eb
Y+9/bBK3R3tcaOpgR8iqBHxRE9ut1OPUVvYr1bbNU9gBCrvGkcDYDCQFp0zlhno5
OXNd2KD4MXKNYVI7ELe6dvvyTGhdZ/Z1STGihg0tFJzT/BP3ZNVkiG1ecwzA1DTW
U8Net+3G76GUb6zVzbh7KYBupt/nWf/ztELG3O0Urb8NIOHy2O/Sw/ipxMZeUzUW
r+Pom2s2dgKc0emY1pIbGAVIajuEcowi5A6mRLi5d+3+rgH65beK/LRyk+g1QtEk
NvAPFblWpLJTRtybZCyWg0PpmOQdRCVXOMuj2wv10NyvYO3Eb77Bmf0iNOxBWQlL
wn24DctYdROnPQIrSKYx1fG/hTcK+ISc3BUyCRRR2YDfdx1307BpeKhujKEqxsJe
YiRO58EwXAGdjNZfNozK7Z/zTvtbRPb8y+RClqEG8eCj3KKIGKMSEBwgpruxjqs4
T0cye/ZEcl75ao8vnnqHODVUAb4b5/XZvLUQHe/GiOW7QygCI/TlbZmNzblp8TQB
+PrJfiVr4ZwRs/sRJzgm9pWkXcwm65rr2lgGiZG2Y3IeeE52Xk6s7tMrMRB8L1P9
ggSO8NhxhIofwsJdAQrAV+h7KUMcB0sEl5QOKvvCCxvIBtF3LjkzEU+CKDfmnxac
k8Dm5egRwMEYEJ10Hz3PrlZ5m+4i7t6719p8Dk20X38kSI8gDUlf/a8DY+Bwegwr
J5SA/qJEwsYmivrO/sjxMLxY2bUZ+p0pQlG4CpHLLMtNvL+05oOkoWoi1JdimmFG
izOFuI6DkFJewHMcx+CL6DplfG2DJDsYIrZ39SiNosMxOFvmSHLfOv+Gc7fjqxry
bcRTMjdkOQ+uICPlKooLxrqG2qxFC88r0ck8wBDGf3f29syD5y42bmplqasBsl2M
kYBzmEdo84nnr/4FlBQ/7w3G01btCbIz8+2ps1440jFxxU8CAw6lRGJNcEzRSXU7
CTmBoh/po1GsfQrfoS3pnu99+0CLDF12ebXRBMnNRR98SPGGilgh80GYM6rk6oBH
YWMZA7omw8eJhQv/xWV3WdUA4m/+AKIJxKWHL0VA1J3dfn4L6GSWBsI8Ol7cM8FE
4DC0RVNRL4y1CtQEzB3ZdElnSa72I0ilOnZIKqVLwhhxDtxEJTR3ygNeh1aN6RaD
P8mm5TojaNsiqY687EyUzwye3crJTvJoI32WLBaWnUcIZuFn8d4wby3Qp3/sLs56
++46XbSadKdpvrTjZ1OnFrNbEERgrUSGx2t2kzWcDOxIzsvPi/Eo1SwrgJiLK//o
9aV021Dxw/p7Ps5kst/sJIkAIsE5kk0Be+stuh2FlLA=
`protect end_protected