`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 19632 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
ZIICkMu+S2rq/yOQyqhpulo5ukDc/tRQVITd5MlhjyLpNK1qGEeSsK9RvWF2qigZ
0eYvg3oBMOm2UftfjO78516QH7AgwtzwdFecUup9uvJN4G0cjfw02tihQdN7PQP6
6ICtG+5RshvY5OSCbWpv6UKp4sWwa9L1kBpi8OKxtdBKpbAV67khtwdPvlt/2CP5
PmBYfaOb+6Br61Mc7KFAcbrb8LYf2UhISJc6Ew8FwumbJ8qr6kZs84nrfeG1c+V5
7eOKPyKI7KpraqO0svibWhDxVAM8dMOtFFx8cyWcCdOrV8nuIOFfziWRV2A8Vjl7
yo+lDyuaBgNUVhn2m+m09sk9KeJxCioozo15PUIkz3QY2+NJbi0dMy6NZp2xnEcB
vmlMcpXzkw0PTSGUZqf/DXrHMbbItJQF/OmUlQewWpdAelb9VH1/kGF3k/57BnzM
GgUy1ki3n7aE74XvHnHvCH4uqluHBb3z2GQn90II1V8tjLxUvjHPGs4/i5tb7X+C
hJqkp1ho0DZzOUBDX65mVZsjQCxYVhHsMaJBYQezwd0J9OoG6lavzAaIJ4ptrq3Q
EURty/1bKs0hVgv80HL8Hn9lmzce3Nbz+VlTPGxtlE+qgeG7pXaYq/4+R3Qd79h4
BwHDqoQsSt9bdgb+F3g1By1VkmzJ41kQ5kqlneaih7aPvaBM8mt/fuIgMnlGAlAk
qDDzy0O6psZy3dklHnUI2KKsglrAr/YK4a3IFF9HKTPqQJrBre+VD9pECxUkFxBR
xzcLe5cBjEHlCoSMnqmuvraBQf9Fl6Apj+Xgb70ddx1t5CmsZA4HIRBdqnkU5VEX
BRc4NrGV5gNN+70ZHc0GzAg8iiTBa32L3UCoW9tE0I5ldIfd7SKomFcsKy+50uf/
PryK2vcUvKodnSKLUAmnU4a/P3hO8/aBbsjAZ8Ma+xeXXRwM5Kkl96oxWIUwf8Ii
mkTRRd8DCppEmI0OHXrbx5GSNn1ApvvT3fl/ksfTiJHtp5Bc7K4+5CXTtpC5kOqh
R/H88JeezmHRoKcPElaNmtKNVf0yI8uPIQ5zQWk3+4NY4dtwbx/fSl8BLH0ATDE6
fEIFV77JKrqk7t3cdGcbXv8TRQZA3nDP79rQ0uG9Hmj7SqF/8eof5p6zRUlyKpiM
Qbmq+2Oiy7nf0m6IKoGk6JtymPUuUo4f6wwHne02Q2RAz/B+IHh6G4mPIOIVhXpi
n46ALBZXs3dRfdo9Ep5To2rzNHaML1kOJA9FQ6pCobDMdHbApNeWV4KieqrcGqNS
g6PAgfS7YFlNLmstg4MIwxwJm0kyEvKL+HD7/2LTJk+xjBrGJmEfqct9QkJUrkU8
RleoPC7Gz3OyrGmud4RRJcF/+PDMuIRMZzcjIKdROTHST75i/ROYnyzJ+p0pduYX
L/m9QVtUsQf+ii3fPP3lE6XrM4fGYlkoZEF5yWTXcRQ/fy9PfbsVsOvh/BKZWOJy
7p38O7KDpIakLHGm5MSRn0aKTzBiV8ayTkCgnCkPLBskDuL9xxSJJibNnWBfOoaG
BuLwLP2bZ+VgIrUbYIWOUCHh/iooLEYGcRbXXyw7kM4+dGViKnJ8MdpZUTmBmO9q
k3x+ZEsiAu6IHoaqFLbv7sB0uSkKiGVdhScpDikEyAEAvmX5qPFsZRXpUJmcnI4+
wI1HS4yxHk+Bk6AJIhXw0KWjpkx434UBxgJKNTaHKYDMHl6squJpeGoMPYHWaQzV
e6K9+6EioPDEJTKf4XtEGH/aHl4fs0BV/yjD3RfbtoCFiQiI+tV2BNyb19r2JFBL
c410d+ch+aTLIzbWeZ8ectv/39Zodgs5gokqh0fHZOtk1aomehCHp/qtldSX9BWK
4BkvhuPg42nubOpjibsiZz7ltmBEzC7WCZ1dZ1A3GpD9pcplUg4rBqpjyinvf6hv
1qwnNgsR/G0Xk6hpVKXj9+ciQei2V64AWZElb8n/6deznaBqBKqgY+TDefeeJWdJ
R79sVKlvO65vy97naUYCtofKr9Ndt5q+X0xZF+zeqhn71u4nXwtj8TXDnjAr2NMG
Cdg3NMOJZARPUJ7NxRs9KPGno1Pqdz0vjUeI9S0bV/LAZEV4zK8sYGZ18vSObtd3
dQ6vCpEOQ1NBG/pWLub9UC/sL8LcfV+pFAwR3hOlw+jSduQPOesd9jpNxAee3pTa
+fvmmTxSIOAYD6LhwRKR/BABjR++yBNZfp75Ioo0tJ4fAJdTQCvliR9yovbq//lX
VzMRt+s++1vvV+M2orxeWd/9yIChHzmw0ug1GUPVbcKZew6WsEDjVaaMEZd1q7Nt
X90Pg0yWXyJJL2GaE75p9JaZXqgrSfTA48dhbpRdbzsBvQAVMoVk/vEhbgzuL5+2
KWWlVQVw9kP4d1krdq4AeYQsXKhmTk5+upQJ/6hwiqGISFG0BQ4vMy9/3hFKsO/L
320uIR8I8GYqCxouLsGn6m/j212VcHU0IYf43B9lyE04aClQg0TZsAzuHZLqzxcS
kdT6Aeky1nqlkS2SsfYDVxFmQDgCF5Rq0ROg4/fuOapt+KhYoqzTkmkIP2TQ24dR
cykyradfD5ck2Od4zj6enWw2LjxEu+e7qDzQS5PCxSnuFLxPNdeJj1Y0E9Wko4uk
W/YOCVj8CeTkhMfHeaBHzK/GpVmqMGr7MAEb8KvAHRlh5kA2Vrx7WzHAfArd5+Kx
hgWG5tmWeHDRZHjlVgu+lI0a8aMi0BJSMZ83xs5ofgXThP/dUn/+6t/mI6H36rqk
nQDU2qlno8KrUpTyPzwpEnwUQOD40NLrtZ6PK6wHTmKuM2D5Id+C8bo6QWYd68Ix
H0TpM8FBE0ROERaej4iJUSoLDiy6NoCKolvQjd5XbnSAO8uudE6hEgZJ5odsOTV9
MLL1WxDHbe9tLlGpln7jhrvinH1J+nIeEVG3V5Pqb4D2M0/Pm0l7YONvMKT6kyKh
QVzvtMrHba/mskyVE6xOcOWUAsWC0QA/FRpDh5reN2sOR47F/O96dttRajjQgDis
PzUcp6sdWVUX63KrGI8PCq0LaP2MIPbMr3MFUVTcdAHvvOWdA6DBHc8FKPjGmd3c
6ak5nbfHBfK5UYamOIF2H2sVcn8YxD/aVARcJHaXoHo/Pb5VHgznrzNVlkWelUS5
ZicFIKUoOllBowj4Ktc4/wNPr9aCaw1g/6pL+vE2Y7iXClp47/WC8EbKoesVu7MR
jGg5vI3djJNayQY6ztzDqnPhDVqFwDWs8X3dboe27+EB5IWNHZjIVJXTNrU9UYp6
eWqre8BLIohYy7wnm9vZeKWzV8d/d6aSnvLEPn1/JJ3o48zlllTMpCzIPcbtBMmn
sQFs9vbR47D6eOOGRHvv4DEFMNlHdJDYYedrHf3Ujz4yvSB+nPET74lPc+wfghZl
Rd6rIyZQriPmX7KjIc042gB4DcfZHY6Lq9644lexAI2u/M1yws26F2wYOF8D8GbD
GiaPEtZKvkvj4/0d+nSwcONp9OhWCm8CtTBKtH4ahZJVhlmJOWSJGiPN3QsVYRUf
511/Aku40/1Msoa6G7Z+zi2YGINj3xt33WLq2pxrzGPgVfM2pBIhsmxAH+yy/LtT
4qGwFa0VShWh1YGaGY7je3kcWckDZuwCxSMFAFugiiUacVOvgOnIqTYxFint2bYm
IdWUYT6hYdeC7Av6szKVzJ9ZeU3B/WmjroTaBOhGDozT1Nh4B06IHDNzrYYInXK6
jX7zp/buiYz7+OyeDl/+g6NSHlDLQrRu1ROzvfL7x6DbMU1F3mc4zIB+uy4wmY+c
8cM5m6lZXj8kmmujijyMo6JVpdWZIA6S4hSnex5YWNUEZLR+f2t3537l7dkIQyyQ
9YRTi+74khx0A/q05fV1Hq/lq6rkVJmLybZEebVkkhXOxa3zU2ljdjV3WejWw4lO
aYt5R86VApDX/UnZnJs+39wYaKnMKBkEeoLxRrbfv+BRaupxlZ1ValOP78CnFWRJ
kZRPxnUbL6EnGRGjGlMdV0qtZ+3k9gwlimC3cb20sBcL/twJ10130JMYNOmXwRHV
Ah9bovph9x6N+b7xfzIjiYtDclmEMFipKxXKx7cYm2maxiEvbEOIjVhYcg3hs/cP
Ral4TuQxs6cjl+loAUPMl/Oeg76OKyjvD5kXOBRqzC5ZgnBB2fBTw3YSMuxXfaxj
0UznLHH8pYmVaOKZY342Vu8ehEGspCvTJH6GSsIcMa4w8iziK9oQMBuoSMenzarO
yfB8BjFspWZzR7/tJyD2nnN2U/NJ/KhlAc5kj5Z4qfvPHArDzTAUIJUtxVXRPVHY
supzB5FSxUhxqwiXoxonuXtO+AZq+rTtD/fY+yOV/W5a4THMEGMUti5GGf4rcf6Z
JSZyUFhJ+HY1rUNYbGQwedYNaxVW7MnGHgK4goU3J8JgU36lSKiv4uSYsbZxc9Sd
FF3G1mKFie8dBA27UhlZfuI7UwQHoy1Y4pG6g6+hWu4GXYOEkbemFOdfIgU8rl6S
TUez7hxGpU8+JiL2BGoeEs33zoxV758+F1ArsZZTgCY2aX3cSSG8uUVbIYiQjCOp
3y8bv6ZBFoezLiJXZFkuhZToXq7GrRXMDbwtmSmCZEeDvGAS/9ANUijOmnhX1iZY
xg4uzdgAzH21nTBsNGAnC4DeKtgtQnCI2m8NRAdfuonBtVYSorT5poD3nMk2rKpC
KZLhguWodpyRY48n4WrCEQzbRKwbRcOYcckQTFy8egq4d9rs2RAWrZRbBogQaGHS
VXiAty8rFJGbJGuPCPkWAlLJoXZrBe0CNuLgfSSmBEbVCGTuUUqWeik5ys4Y1i14
pRFfX1QqrPlM5xa3GaqkH91rhzzlpP5sHbpfJMcRmWM7oRBpEGZzx+HpYTFcCaB/
fjaXy5KQ1X3cGWzWr9BZaSOlgZDcaEg1wFA09y4NNI0E6l8BQ/HyxsMdG0o9Wyuq
KPqlzeqVVH3UDan/Og9xsjS4odOLW4p1+XhwTDEKh3+TP7GjaiuOzWt0QDxF2tZq
/o4vagJs7hwmvzbTqOQkjpmxqqZlJyiY1dLOqJ6ksG7oqBPZ4rkIeRAyauwonVVv
aHApJPcK7mEolUH74u2m2zzQjyWp4tWKFcR7pyn4EmMATVsptwU6FdVel8dOXSJ+
usF+7NMOhq3+ZCiabttnACbdQ5VdZVy598H22yFDsrrrhUm1KOG1XXaz/gYPBuT7
XTVxuLOQ5S2v6+ryG4M2Lh5icZuKDgfJ9agg8ZmQBuLiH8QW0TXKNz1wEdX0q+Aj
PbxP+nTR2H89ZXoVNVqmouDGPO6RWTE/N3ha7hTRjVPXtNSGhKQqfnEBd+ZM1uwL
IcD9QIbfITOL349F6dDycKG6xiiu8gPEGcSsVo0G7AKoM2Ux2YVmpPGRNnMkyrKf
nqAgj1RKLHhxHjE3pguCSdtkarqKHdvMRIsHzp+JR4uD2+Wyec0k4hYVG4jIkP0F
S/UvestprViC2UFMMDzv2RirDgUEfrhRFR+/iH2J3ojfbdv1G+AGqOvi88D7eTwc
Fj3CsuOkbBzwGwzyFCBkEZpzJEKiZu3AppG7U35HPOtl8D7OVa8Pcl/73GVxYqYK
ulYm85nHfmXo5K80GzBIcZJX3CinDE5fuosOXTSj50tzBTBnhyAvpxbJ2ITcM6IQ
FB21p/Qm1LRJGGfNmittVDMjwuwXbDxfMg5On6xyO36Q47fNMhgGCwUNSUZPodSh
cfwXq0sMn3e2PJxexjHcXX/2oZ9x9h9H/nySlb+MBfjMlBGvHQLE6oLvvulsOKCK
MtOnxMqW6aHtKlhS2LpIz+tG3X/CQxH8971oLmSiBohgFhUTiLlgzOu7tT5bq9Sf
OBeoRITVspltFQ2Xm0z+o0dtdbQiOE3Qk6+IvWoxsR49CDrRxRS/PcgVLhEwQIC4
ot9ONUnjdZin+dPZ0nV7SWRvvcVJYYPoMPeXoY7Bq2PLM5mEA3U1VzAQ9X0kixmi
Vh5zgc2UA0tgldfeaBZv2xC9OoSGz1Hw1Uu1Wn2P9cwdQ4roEWL4+Qw75Qn8dj8H
ZLIa08ogh0W5XzsrvInvncskdBHUYC5zKSBbl9IIWNrPo0EgUnOt31t8kMq1H9e5
HVes7ofFKmZpSssQStEtLxOjkfcriXjLOQw1vK1EeSj00iGFRFhq+/wcZohKA2eC
C014EtSO2YlyaDFbwPzxuT1v4PwBG1Om8FVgvl4i9F8bQfRliSF9KmTlVgDjfPOm
TIXjUUb/cB11n01AN90QCPltk56Rka5AwaOAT8UKvwsg7CIxZQTk1jL+drwbHW0u
PyX9Lq7AiixTXDrV+pzO1/qPouDZSq/RFXaJ62eh54E9wGNPovkZwgD/CIUWtj7d
Z1XuJnuxNBMjAcSQO8UaMO9XLlv+drF46rA6CCSdOSzbfInSa+5IwCkrByfCWnx+
porxbs4FlCjMSTm7Ja1VWPufY6MdoDaKOPDw8jIyE1XFFQ+zqhpm7g26X2qVH3La
CRtIhh82439wIhucwIQharNpDlMOYQBZFxVSVOCvWdTbY/ZLiGJF3BZVJ4kQ7r00
8gPH2nBAftx5OqAO3wi5qJpURqbnAIeI/9ZUGEjNVzZU7xrqRLFng4sxawIQH4A0
ClMzrCRN3br5svhroqPclxWJQMlAS0mduwOr9IWK8tiNsSVULta/s3mjbTIvY0cc
EWD92dL/nPSROR5wKlYBXyzTz5f8q6c5qa06Ua6x4XUvOD6MI43L74z5uO5gA3X0
Uto5DARDi3aNhhdBYJ5lqNpQFdGFxJsqt4io4fTQQr9lZopJTTKPliNFAuDPWNtZ
VzK/1dKKQsPSnJd2M+A4n/vCmTcdh157ommMLyr5fCbHUuuqXv/jdpApJudbsrpv
g3Ysh3nD+ktsmHQZwPpv1w5NJoU2GRks9G88Qxe7Zw7hiHxm9FBOgz+i/t0ffXzU
lut3vDmJrCuYZ4KRxHjPguM88wRvHe4p4N9EiBB4wFmyhMrnD+vx3B7zqo48OVxZ
xoSx1woM2AEzznLfGmWkwiiKwh17Sec+tVRdiG+CdT36EgYluOtO6lh2xsRffRkx
fqpEMoL8siiT/FVmScoLkD9aZGM22lsF2hcQg4TD9Fuqgz2w9UC74qlCjCgAlgte
vGo4L7a828aJO8BLEwR4h0rj4jnzVlFqpwVOPO5KjKeEfSnp/azrOus4NmMNH1o3
CmTvb82fOCl0eKEVfuQqv0SIw7fM1py2cluwKyShHiPnLq1aeM/5iAK4K+4hmSJG
KAf+vbT4J441jgkM9qE2LpBJEwTwVBefdY0P0FQgdILRV2Efl9IpMPHGdJx4p8id
BhONacUHF1i224MjvriJmF3SqaqBA7u+putVnPrc8Pq1ESNCXcHy2I8NhWhrCY+Z
t7qaZ4UjQhANLsnHNSZcvNiRmNGhGDUoRa8yoQkFr6oEFWPTkiDgSWUy69AYqDDr
f3GWoQPxtyE5ZSeA1ms/StcQgIupJlzXEW2B6wbp6P5b9ey11I6Wijue2N5jFxzA
W4/gWRxW9d34kj+6Bt6g5/b8V/c6QWBs7Q7y8DbbvqajN3QfB83bG5YT/kzCx68U
1hdHMYVsVS7Omv08MpOGKWUirBmSMHgzRdEiBcZfLMK0MV4N3Pd/1SAYvsiMFchF
A5T7E9typ0Z4BnrstagBTe/l/D0JnZ8qFjnuKqYzNSZsrF66iMQIJkYWt8Cm+Y/Q
BNvH17U/LxyhRO+Gj0WWblzvPejNXj4yVfrRMtnVNddpCgljjmRv8snG5LPKTkKc
5wP6UyhdDpgURazB3207/e7gZi4aw7A8DqB8M5WHpEsNauo/8kAkVj4A3lXBotKP
6MaJoLf/TT5srKIQBqRdc/ZBVYrkoyvA9F0TiQ3b5VMYdn0lb2XDdr8LtbvQ8ecU
bxn6J+myhuNzGcCUjhICrKjv98WeM1fBUn5BmHQsCxAkilfghdLXPTimDRNnVPP0
81U5CUxP5esyBET7dwIqvhd4/BBAXkO9dXTPECjabFqjBVBpAKkFEMox+iHnMXvj
G1AOT3dvXh/acv613mlKl63R556bKZejJ8ND6XFW2Q/f5SdqEqpijwHqU/Y3kfT4
DRahM47NGiS9vasVxgNEW5eZJ4AL29OCW2u+HA5qHYS6acCQo/0zswByZQIkbMUz
GDgoDOMFyzVifIUtPzvGBvP5B9Eyi63H0t6OQyroMSlLQhFzYpjcCvDLwaeh97fN
kvs+OkX/z5AGejsiTvEILlHKp6KFcWehmTK8Bq5dJiP43MKWF4fmAqGlsX/q/mZs
xOY8qAD4PTluTaO3RRok8NxqRlevm/cvMeAEPS3ah4zXtfL733FehlA4sQkqULRA
cleo9zaW01a9LLoM/FV0SKP2/Ev3rBpAqCGouzPHw7fDOGqux945dL7oQvAGEobR
3KGfnVIYKde1xPZ3A14AkkOIZHvHacZ8ewpHqh71zWR8Y8K3+xMwAMBgX7S5ua+k
wI5c6JopwSsuIo+WFPTpZZky1F25IWnutMc4qb1+3ZPWjp7J3eghQ7I7PNgeutRI
Sz5QAFBlQf6wMZqjvXBcTte9dePys02lZoG1K1v4OnmG1Upc2xMfV/VnMHU3uLi/
2WcmQufrHmkcVrWHIuSgXdg9zYNCDnwuRtmiBz99QtcQalqPwp1N2rConAM3tH4M
vg5qoty5Nw/sPDNrXgEkOWO+inxlINlkAr9gEp6rHuaNVjw72u0paW7TDMypGVPk
4l0btyCGrReuI1cEkCYxhwJW8rD0WWrPbQtMMV58k38uynNly9n/FamS5F1MervI
fFTt2wTncgk1G/FqJGs/IPRiVBmGTWESQHszS9j3L366EFzaW6s8ijsMhq7np22g
MbJy1NIDLGXHoAaWm27lneQLJGn4w66uhnoWO2QgqFIBHq53MprVOIZex0FSJSs8
BWcfRd7I72c4LYNsX92PLhiHeKZnx81JojFvj6+CgLhR86fdRu+gwTv4qZNFzssm
5/DmFKcalbdSSOemorzo6r+3tPs6RAQbZ0HLcdA/mOxrbggd3abArQ6bUOMFAbrF
64y02fWzxt2h8H79WVMt/tEo1q5voIUED4X76yUYpA1OuR3sgtaW3y5DCCaofJRO
5r+KzM3Bd3D9UhfjBiY4FB2WdrMC2CyNKzca+DurNAItcFRWsBMYN9s9W/5h//GC
bAgaqUVeuc40kiFW1MI1ZgyZ0fqNWt5sfn8Y2peJqAsmdSi1MvlxhghhNM/egS6K
7vHl9JQK2SshH2xkVdFCVqlS7B8lH6ax//uIyM8pwrczAL6f/ZowF9VroOyuzkDX
fUyC2SbPXQH2gFuuDrhblo74xWN4sERveKPRj6pavkXNwFIZWDRczFX2U0tqs08w
2OHfxOHUxav8z/hbmB8Se2akDRoxC5cihBymLLxiU57t3GFTPUD7oNdIrlv9jbmc
L80pyeXzNBa/w77Xx8xbCTSD14YnY8YdPYg2TYtYXe9DC0UuD8YXIqtR9BMkGdgV
VgQVFbqwW2OjOeLkgnVjQYkAD3v82rTwyyg0lIu0tLpTO8K8EzDC23W46YkfGYSG
G0RnVIhlshgvDLJ7js1Twhllwv843oPXyqBGibVljXM5CYCABLSNs6sHL+szjsjR
qV24BlOv/cJ2hyNPJLrmjg9RS0/fxH149Tj4+vMsZv7spQnWWFYR3/WPuyKDhhc0
6FA1BoEf23r+A5Nwh2t34hzfHbJvSTunZ80zZhbcUpU6IoykKWIT8hJ+/w9CjBGZ
u4PTjEb+2mc2iM6REPNh8EYplaUyQj5SEOdync7HBCuyoL1tdPQsafd7PIAOBSLM
myb1R42Vdi0+eV+nS7PzXqkQE1rxr8XYKY57LuxS+TxeZZnnp9GTSVesQCmsOKac
K2PXWKNh/nCYgRJO82C0HXq/py04Df6kL2DQkPDNasjJp69lQ8AsH1XhdDRNJY9I
iERnhPJwtnGzdO+WOEnlViEC/DNxm8F0eC6eXAl9kCjwbSkHS+oMvYnqZSRLyB2f
EeNoDenV6jXA7i3M5Kv/RyV7ZdpnzrXelWTWF+ClO+12F9h7fikNAsO+67z2aLSi
Vz78xXXZF8BiR9/5Z1UQdspqRji8FEU46NcwtN5XRvqMz2f8Pk7Y3icPUfJjHOTw
/RUTHt5oceDaCAbD6XLOB/vOpGNQm+Un+S4F2tkSNuHI2dcyEW7lHreGhEiIKtsQ
wWMneX3tqS5U3kwPQjyB2zpAnvC09kjN0jIO2HPN4fnIEYwyShO+kiiiv5wkO8Pv
927oMj2wAOHgpuhaOxJp0xcVwFfVQt2VbLobuG+8SSr/0tiAXOkdF4ZL2Hz8NltY
OL4gjyIeOvQ1pikE4FiPTIRnwt5OYmeip6SvKLzlX9aAf0dK1QbVHuul47s9TBgt
WzykbjchJwmUXVvD8xLqg2gb81IP8CG3JoP6JP5n7QLisKMo+b7MqT8nT4xc8alm
KX1+bogc2fiPRkMmiVBGdOi7oThklp+/aSPjFmzHGiYrKoKY8LoehKQBpqWSO0Rg
9eBIgm3lTQGYeanHZZgMBw5fKGVOPcMzcv/PCeFn3oBJMwxL/G8PAf9DyPObKR3A
JBZEx2qW+l5YPmDirr9zJc9mVWlrltmgS/roQfC+546cvoqCi6TouHv7AnfOAEzP
oahVW4XWOZwl/qD1NFKyOfSUh2T+eGCL8ijNU2wF5LZPV0wveIQvUNyIgTQiRvf1
ur6gfRG0Ko0QRdrlkZoWONT0SnIbMSOIXvxuEPgaOHf3zb4Yqc6o6z0XBgpZJ1EO
hp+4S2DcfnL167XB+CCcnF3Qc309KW8ZBb5bqeYodp0Z5PoX0P3EOg67zSTBPNNa
2q6X3AmfjvBAvTuk9qYxKiwFH6Se7skxNUE5RvPDPszISE74cL2HGxf1XF2Y7gOM
gSYQHxUFQu4xRYCb19+UtGPBbAJhjPEbIK/cQJA7m7YVjdsTMKZZHUzjnXVnAOdM
zZr1LyIZbxNc41rrwgyYSiCssuBZGU9xStkvDR94ngQyzGDW4sxwgVO0Ha9BY6Ox
R9NrzDXSgjUQdspnw9vPOwecRaFZGEaDYtdeSVQ1uMORJNbMaxIZss6I4IAYOUSA
Zl4Fu2PbSmQhMvicrtyuWicMVImwm6Ke8UGHp4p2iy86RU0u1JG0/HnBlFog7Kwc
EdmI3v9SBY5OhVnNsT3S4daLPqYT8RamwyI0J3HugMUCyH57QtRyOYFcJ1ieoIer
8aANXUihwM7A6vd186ofpY3kya/yjRxFdRG3qYkEiJGmigCYCg2OjO4rYdJSMTkr
bpLeybcWKlZrdsUwF1aucJdGzZBqbcKbuVsCtgd160hXDMAGdrKZL73a+ymmALjl
pBXr873unV4JI4fX4e+biC50MRWhEgaa+mhKALf4ho6ANMaCx7+SERao/tt0ScOz
yqFo7aA1oMvv7zgoyx0FbTT+xNUaRHItw4oCBOXf5DGSiGqgm4SxNlXBcU/NNozB
/V5Al/Eq0BxLM/mszU2HMN7UxgtV3tMShKmZ18fvLdUnxVCi1i+vsciwSW7R7Mye
0CfqyM5IZOUI9SAWhvWmecgrwJ/zG2zPBrf2kRhCz3+oXz/Ln3a6ZA0hUx2YkBRy
Tjq+Mm3q4BtGBKLtnUdRNL5znq9yoCCnJRUScmIzdRA1QL1vKpWsNyaf1zucnMPo
P6+c2DSK2p95JuQSg6y44a2okjAzSExVl8+qF5VupL2+DnLg1z2PrF2p5HOzd9Wt
z85SEOW6JuSQtDN1cFv15Sbrtwr5sK9qpa+4w2W+Z1TG+RyManQQJFbuzfk72vX6
3s5niNYmabWYCNKGjIm3DGEuWqOwgoIQkzGKt5G0/PeB3urbjErkTpwkSz1KmvSH
O7GPnB8wD3zbkvUwY1Z1lSnjJLC1FyPGTbMzq4EBoUT1X0wdlKm+HSFKcT2holQb
+GcPhkJ2sP5Kg2HElxvwN4MPhb/4e5iRqmI9XOqCNPYRCG6aRO3dVbZor6m+MzNb
+LUmoEFgjMwEjtzHcjo4s9lkvVBd6sVuD8cY3EzzEXE0RO8LX0SfyV/GQO2AGDJX
z7JeHvYlzV/VbCyEUQsyETN+znbszgYJyOQV7Qie6mOjQnPEfPpCe1GDaNLBV5V0
MWfuDEJRZuHeiSAwQY+qqus/Ps2nYneTdU79qHrec373F8cUFccguoK1Gl1FMyJj
/vUhLFZ6FtMkBXSC98WjyuLIAFCpQ9cb5ABr1CiN9cs0eEMd6T5836uB3JiTypxY
mer+WGmAx67S5Pfw0NP5ewwF3TXTFNA1pw6sL6m6fxPjTv16GXJ5Khqjdg+C6rkn
TnQlPoOhZMPRE+Fdhh7WdyRVr73RVyBz3XAljv4GLitFaUuvE6jDnvaQJImjgFmJ
/hP23Z+ZDjfcCZCF483QvGb8d3pOEy/wKfKG2837hcYCFdCX3wyxyxlaO6xE1f3F
wu5dyuLBw3UqbbuDpCYioKjx+NYqsFD2Dt/ZGcdPnPmqg49df4qOEWghUHPYJfqT
CC2XCFwHhNtVAjtBMzknzH3zUnzEHX2YoPi5P8qgBLEXXbTq+BYrfLCfuXGYlchZ
8yLlrLHlCtZP9CdcU525ReGp7cucRif0j+q4VdjEjgznm8yHMGFz/8BvpDslBFRm
88oiEP/zyyVbZyDjai9+me2FC0qtBGGye8Ob5EuAX1eXIsJPzAGBI0RKwieOwY8X
WpO5O+lJ2vieJFS1ndfWXs+H80iYxBt6HYGeVIPrWmKuS+z3+iIjFfXn8z2goMIC
jN7LND0d3sfcNScsI3px9JsU0bSbIXhmIX96cD8BeMw9ecpitckmohKgAt9EeC2S
InOtZbJQm3lVewjiH46gM1MJARrNgnll9SeHSTk+g4+wQxp6a4X1h8Btusx2Etw1
pBCjU5T4zLxTmUnaZ+/2fSHaOrvBWMmJ/kRN4j75VZ/Gb8RONiLOSMZ2QK+7z/nS
TO22k2bO/Lq04vIJphLv05qbQojHAZFytwwjiHM+kpZnV+5hua467ICiiFtPaVGL
cLhKFMknskWgcjqmnoucR9+LPSITFbAki3/zMzGZuBuzSVvjuNy5N7wOVwOvZM40
rAcBas1JA+c32fCfHaH7kL5UouK+SioqXbfznk9f0yyASJHOw18M3V/Xj0SexmCm
aCL03ZS3XF6BGNzvwPVemphGRvUkUoY55fvhmxVjsCaINZXg+6Ctl4TqeVzIdzXH
mcwrxwX19N0HLEHMVh5PJebenRRHHvNLWhIh50Fag0ilyoW3LQpSkrjqVjR1fQtv
XTgIGZM4qDjvSi4MdgMEsWP5h/Xq2RKD8EKwNBVCATJP5/8vemiRksdSNeMa0TqM
60DIKRVh2JSXKyBMQjTXmcZJHQAm1vYvhxAwE9eh4aSRZ4HunjKXO6l0AbfVySg3
He6YJ2H942QiosYx2zaM+3kZwy581Uoydvz1OPf0+PPATRzLuigrvFCKjzWZK3J4
sIFogBpoDTqwhID3KZT/MkirIYWxvJX/nchPphc4OYCSu0VXDqI7A7OqWWND+q2e
fhO6GBpEXOXlHYkD8ROxJeJH0Vb54VE8xk2hMzkym0ZuJ3Isyx7PV67jJSad4WrJ
gBERptMF2Ui5hHGIQ3Y3ufJv2wzPT1IboeQOSJyv4POyPSxkAbjOgl/+iJNw4Ig2
COtmTyk8KWew1/QaIifpeOnwI2rvwwXtmFZk/I9MCWs5zgGUWRok+M0xUupbX1Q9
KzGP7kS+3evLmmtjX4LATczvK0didV1EyqjdEZB1uZKl5PbMZPJIMK5NnCe3dyse
cLDROH+D2gWQqIsP8ukWH+dJK+i4OiYAZklXlypbmHfDJixS2VAu6eAL24UWS17l
J6bDWfsjMBSW6JCN68XLr5OUWfDBR+8bhHAMHosY96wbAPHl34n/sQnaKl9+zoke
pA/hBdlgqVeHexMjaD0QMosU9b6MqqdzC84P/j/F5TWEZKdRlBy9xSnS216+igtQ
sqK5C/qjjXIvGAps8v4U3F1m/S5L/TxSweTYZlH8ySaIlRUNYEso/pHtCBHkGq30
zkg2BJRi7V2LbeAGmH2PfGzkCeaQYNcae8hJ/jiL3btsZZWofDoHr5V3/8SyzRMI
zHhoSP8QpMPYcO+5C/vY02p3iA+fwRSHKcDeTLvO29gn6Jfrnq+knAY+GQNTlbtU
XZ77wsDJ//hKdtHO2f99kuMhKH2+FabLnP2JtooI5OVuW7NBUAZKHwSc/Jjs/7UB
x0g9OWlzmfp6SnfBoxeLFpb1QPrvDu1mUxcNCRBeqZICdePOWKkhmZkgwMNq0HAE
+DPzs3oMEvg9bdAIxnBNtwFk/wScSLWUkLV8f0mkVz7ILN+3pk0BSUqojIwJ4PwF
XSudwlTYhEWWDOLbDtXQD9s83OP8Md9RSVpt2tq/E/Wt16qZW8V9R/jA2x9hr00p
wRyAig6xvHU1i5IQQU2ng5bI3MRhzv5NWObJ1BMbgPnGrXdOa7x7aIEJGb7QHGkm
pgwsV6EVXnvzUBAxOOoY5+KlyapAMfGtgOC3xG9opa4tHZNQTIXAMPLwSUvyb3MF
oJPS1yuR18c2WxW1sQVrPplAmGWf2Qf4dRzI+Ig+k8I0qdJA75ylmym1HIuMW8j8
9NLxy6FFZvqLe1I2pR5CGOm+UzVQb3V5VW0EXF5d9bJHktvfBEShnfMU/vA8Rpdq
S7NEUewQtI0HiiN0Iim+hw0Z2WmyJKDFaiZ3c1fL1Vshrw2wNEDfIVU7wAN2k0ts
PNfJ/HVbUZuHT6qc027DIBiH95J8wvgZS4LE8idCE4J+GABlnEHecoaVxbcsUCmr
nCcgN4YpbXKiPFt2W3q7QaakNhUfdeFcL7I7DlegkbpVpkOkiEFRXAXWninulxme
i7fYEwJ6gSiKXBTgPkrAh0/+3Ftch5IiKOEPhMVbgaM1jrZPJTNUxplZQSmRxw2S
y//zKdO0gjSf8slY393E05h8+Ow6h7a81YCxVD/RDTOh5OGZpm0+FZvn0peGGZ9G
UyruElyjLLkygOaCYkWvHgEHBoLhFDMzepGjKxhwX40bk3r3PeLlpuMm9HxlP3Uv
IkYmI1MTII9NDreEGDP9P2NHbbvMhIGE7IB3DzuiXTmheyyrjBF7xiZU0VFRDfvX
pqO1qIxBL8+EjNNhcK6+1ivHxVTzbxEEwquUbCsslhg6Xak+sR7S4Sgrduo68vTe
zSCliO/VqL9t9cm/0tUtUgCgpQwdN5e2h0nxzDhHg3nX5MfRqwZQQhvklr7pEBHM
6WxbYhrR1GUbhWM3EhASwKpHM6ZMICLkAs2VxW3gq9x1a5eN0y3pqkkwOqpYnmU5
7I0xyi7mxCUfI8OA4T5OrD+f56KKFH4mwCFUvHEgChWXFV5RwOL8eGDXJ3GdYSIs
Hzcjoil+Zeo6VXasEoYDvbhCpxvOMmIWt14LyObEX1BFQWIjROKcmU6IWFEQ6Jar
0BAfG4j4DyvTG072NbPK7I40H5O3fVIKY1GrbDZ8vP5V74B7qxnm2tqH07EDP3NS
XkI+wS+g0YGWYWVcV64u1C9jnKB8UGzKE6w8zOFFddCxU57CxuOLHdVS8im3+LQd
OrlBmCOmWDUCOZTPGz1yP8cF7x9yMTjCc0f5fLcrK8Xf2JUijWG9BBgKvKso06wz
tff3ZSzQMFHaIsraONQYXt8QNa/pIR38nQEjEm801QzeC3LY/iz2kV4qsdDSwGM/
fd+4KIVkxgokQUVsbSsABR0HwQvbG6K6aJbY47crjCHPlI6ipYud5akrjrd5pVqf
+yoz0UOMbTKnjA+kPpTVPZeKf+Wq08xGWBu+HyWCqxSJ6u8kZaI/6tiizOw2pKqO
XgbKh/jhcrL6r3vkg53vlcASdeXXhimR5gq6hzjibhONDwbbw5t8EQn7td68goP0
8p9rtXlNovjQVttHVh2PLjIuylqktvUe0HxT6Hs1dP/Qcg49VCYJpH+twqZJ9d4V
97PWSAxrB4nDoLlb65gMJ97hpvbXJLNDS7x49ZAlCBe5KYbo8Gl491aJplCyvnYW
EzdY4VbRbh4jKGbGrCqmCPQxWtkZ8gf62i3DllaopxZtwvdrpsuz5dybReHMNHPc
F53fgcnpa0nLyO2BX+eoHMzWRpTOz41Sxvxr49ZoQkjhfvlfyVKbuOCSKBblD/Pk
TjwTdsVlzoW47CpxD3qcklq4og61oyjZPZTxq31d9WTpJjL0fi3Yl6ZGSwZtwX06
PAqc+HmS52dTA2FpJxamAq7NHoCTamez68YwskW57jQmzqPLVCfQ+N1ur3ow6IP5
eBWHj6x+fy7TWM+kv5vslu2pHEuXDcSXa+ZPmHa6V97vh33+nIm5Zk7oWmqo9dD8
to5F6f+Rsu4SCqjfzzrGoC81RpU/JdDtQVmJhjEsNHYOVRP6xvzJmUTlx0t3QHjt
f04IXVwFuNd1DU6mXkzM5wNGg50XGkN15CKRhb4uhqaWB+zvYR8cm0zR0Sotdvvm
IviAOylL8FToQ3HX390pFLYhgSBfroENTU8/HvFWCHBEvRd9A/m3KmkLWjHqTmAL
7uJtgXnx0FnwUBdcx1j6sWBOd6Z7LOYcg1hVfTwD3HPu+xo5WOaZihCr9A7cxIy9
fPonAuvQFBhi0vDBwvIZNSlTGWyGyl4xfrpO9lEBOeWBtrITCyFE5pZgAgtN8XJt
Ilc970rgNH4kgd54gMB8kyDytJFZTcMsfeGbjlycc3aTjGJWFl3L0yHw1fpjKLKD
jkE5iaOdKldZhq9+4VfzN7ZAKrN9wBViETCA2jtIvs6ix5Oy6y+ZAnPzWwSqYkz/
TlIQ4ZpUfq7CNCrJ7eBZ+Qb6YWUGXqV614i3sn8rDnamzrPSCR3AMS+n5s9LHr42
kWInyTAdo3HAxHSfinppLJJ1gfllcZviniBb9jRAxaWsNdpa2ZkPyFfMOc+mLTbd
04Tkiekkuwc1+EpIVVWaYtkyepZVpKYT7o/NtEZJRyY3paMV49XSBHNhwTETQm2z
FQAGzUuWR+dmXZ4+OqlZUWcqH9bOsW7NmLZnJEQ1+1xaGqib9GKfqn939m5HZEwI
sy+KRedCjAeMESKy76ZvW8egung7+JV3PCq7q/HGVO3o3zJypg66L8yTYHw7DneC
1ov9CkSimxvBB0/bH3tRf05iwBOmZtIJcYipLzg2dqBgN80EJR9/E07rnnf2Gqi4
Jd7ol60IEJroiAXhqXGd1XeU+4ypv/BNJFMvn1PcS7XTmD7qIptpyj0wqNnAJx/Z
q9QIcW1yzki7UfolnKmB2fdz5ELIonQyVnba2MQfg9U0HBmH8Be/3dsK4avYr0zT
/dwMK+ELV2+mP8Rxa0+J4oJ0WbZuHK+fwtPWlrbOGKE2W1jxyG0mQTy8kjOVKmio
pkUXrr5ZBrIwzTa79/w7vHXodLZtXyRWJig/W4sdjwb6JcxzyCC1k21bEUWWwOn0
U7+2UWdoRWP6bsjUEcqFMHJbRhMdOnOb5WnG+/NMlpmmIENorZ78yOLDuxR53UkT
7j64OMk1Y2o45r1JPp2Y2D9obAZve3zNFAx3wvUuBrZPFydcLxZ7/duSMHU1B0bb
z8MgWCcULMjnRdVIQZmLqtKqH54Wmyk+Ym1NiVvNCCkf5m8hLR3iCxdC+zb5n+2V
xtCJMEoNAtMHvSWi+w+a/RsZFm4txKFdutdef4D7xyyi31FQpGPs7fFvPNsyLktJ
Ii9qk3L1WkojC3DKBtvovwlfo4hyfj/sG4wFFWetHb3f4WnlRfMsWQq5c3vOLmHt
pg5mm8Ud3H2jnx1ePGjMt8hwGvGmofvj2ivwRikg6lJAdB4qvxkQsHIMHGCuHy7F
ZU8mtpWQ/E4BvQo8YsahA9Va6WPwXFuaaGeMI8uIgJUBCfQJQ58hxBGMhka3QXeA
9jNxsPMZvm8D9srmtxC4xnIyrzyzOQbZaNQWjUyRZqSDeU9ig0vaTuHBicjnhA7T
aJ0jjzd3h2ks0SwTkXgPPgvkGD7J3/UkLby7z+6x22L9C97Gbvt9OPRB2p5oMWru
OCZKGPpMv2F7Arwf0RJVFmW8JBoMMZE+3xC9LOlvHJ1BItS0f6j3PyDeIHdsLJtT
TI2qbpN2CFF0x3gzv8PTUB/NjvgyCeHl3YFoVpGEUIaO78n/jwNYmdI19pxyjMnb
I2uTwFYHCYFSge07ZySDS50MjJ/Y7h5wa5YEXNcVvPjtNj3LraaJz8VSI7OvJyVi
eLEpS2mVDluo1emIWQG91qL0SBCEYJt3UUVG1uk8bZ2D4i98jaLBSqqPQYhDBWyW
bLMdrR5DYJX/doaJt6CNHELgDMQ5t21vhcEH8XVAgeLjiFrZ46SLN5aESTeN7Fu5
rRho0Cb9A+YMvNIdskD1ofILqVrfLLyDV1i8TPXSH6y0bJ/KFHOS14VbEuhS8pYh
OlmKBg2Ec1eLbVUwJxxj3IslUEGbFKNYM9nZGnaTc3p9Tcdz7qTrNnFQYvPFLqb0
Z41Mzeq06iz4BN35DjQJgYYjngHz0EpTZ8oMfGtXlQNLKuxzPeKYEvNdyspTa+2N
V1I09oiZe3LY4IUieb8z62TZSLmxZosnrtX2wqT7YEMHgN0DB3lE1pYI9mWIni/v
KWDOcKj2TIaW1zXke6wTrJUJnsgoxCeGH314djTtKwxb+QKtaSZs2YnGWqMyKK1b
gUb0Z15cil3+ieVfAAPrhATI1BRG0mX0jzWqz6ISZh9ejH9jVWgjU7wDjcb/hz3z
LoKPccADD6+FyquYuEw7qa4ph5GXG2JhvIM96Ci9fZoZnA6A97MN3eJ4uGB1yKMu
LdNDTUqJhzvOehDgnC2erWagxSAlDoSDS9QmePKWB4o9Qspg3ipUUJBblXMgR2nd
p2qSXQYELUUrYQoFtoJ4bEjbF32kGTxhhOSZHhNFi9dkQ7hNqUZ8gOrJMu+mVPHb
zo1DbrLccv3ZoCmrwY0y7hszU8PLLo7LDFj6QfdSxSxy/9MoPKpBnZx3hKfDjGwF
5egRQakXoZbiByti7GCNmojXouobojWmYPPzdivlGTBlPasbThNhQoaNgPGSyTCV
UXiixot5s+Gus+23GQe+73D8HKm2BACgAi5IvnwpKBqvhV5fdopeHQvUkMg+jO3B
OChxg0E8Jmv90rpkfXOD3OulXgBmJxLDOwpd9bFnA7/w1A40+M9K7JVRmRk86ZDE
4mTUaZlHPJozGyNcDIqGRipq3M6+qQ3vnrPPmkvPAxhehT3RQ/BQhknvpCGMyp6R
RZqPkDPlRwI36g3s0ixEr7YerMYk1HnoOXiIVbkf3Ipo448/8kCNEcYB3k9Q3QJC
lkMR8R1UJ7iXXj884bgt5ZCNie/Mv9AFQLa3b9nZ3FoYiSR0Xa8ED1amrT/cfhil
GeRw/6QOpbCr/GtdkTXDDr7ee1IDe0hqXpwLXGRhZP/NABdX353xJ9OiARe80SO+
DPanqGz77gYa90f2N2hq4KScUifB2VGub7Ct1dzrrWMiwfz0f0i71G+WD/5NH18n
2iuxUzFSxkub6nCrmDBoWNafTEhabjt89ysIRZRMLl0KYt8WPWPv9F0kSQ9sm4Lz
dxJ/IRnnd+XoX+OCYU1szNEOuIEHiqmfP35KEe3aBUJNp9AHVhdxZ0FduWrOqoSE
czAG7O470tdvnYGfo51S3gnQU6mLKi2AG7pyFvH3s/pyqaTrRMrg370lG4mDQ44A
A62VzZ/DDfiHVPNixY/T4ggmRcwufotIpS4a1TH7DeqZfN8R7Tblfc71pGVsZP1K
DfOWRW0DNUQIx4hF1Hif0KT5i2K+7zl2uEMqiw3Q4VRwCqQhPd1G7dM+InWyW0b7
2HBq2Cgf0NGconSJT5z0Q8dNvifbsMt/KDrH3nfnz+Q+8oxAdRCbp2BQHhsBIXqp
dg2wrRQ5NLP2vDXYttXIMJeuy+GMVrlg2ZE+cWMHU1b02LTr1JI0108XD/wNbJaU
dNWAkeyCl4w0F5Yohk7YpNqRzCRnwgpKO/EKIOYuicUuWl1VFet2tYpZfYjkQPNO
jwbkI1NQXO+07hLwRZhccqNf3jkT7B+2wEsEemV30fEk1CIYgJ0ey1h97GqYzoSn
If+If9MLa2s7T8m/aeVNSEwQR7kvo7Ct2NsNkaFxshpOgMA1HDAvgq6P1DrSm9YV
XH+xUh1nz0YgxU11YwY6dw36yeDXDJlXs8oo5lhCu1zWTGKidRegBsYEHnA5fhI3
x2pTwwYme+l9p0R6klZY7bqqmntkKLbspsrRnh4e5NMBLYY4r38LXWzKxwlxLxct
usbPGFbt5U3xJ54PCB0ytPtlXn/JDMrY/4XBA7B5KxptEwEd1jGGayBLaCsr0nvp
Sw0fHEBNPNIoxjPRfXIcNDaFjigCs9JlCAUdDRjJk5TT12wj9Ynzh7xHsyb7RXQP
70IUjkjmc4p1eQUYnU8ds2qG1GrjYfeFGejwaHeAtyQvO2QwQdX3JUmlirODd1hT
ISSoJJ0AANQbzNFLyL+AkS/D0gMlrSts4aHre2HIAQhpfdJ4oE6rcvHTEv4nNePD
C9jkN808WlWoWMIvq+Dxfumun3POlUUSWytyVaccaW2ntnAo+KgmDaeWNBcU5yP6
BArDH9JhxwdzPpmtN7NsjHcLQVyxXkzqoV1eTwHJJKCXBJN2KzgzwhXj3HcUXYqt
Gvyrsq1RDygaF3ap8Ybbp9Ko8F9Q2UVf9rQvsbI3N8Rq/Y0Tz6rU3daD1ZeNP5FF
biOdQacNljPEMt/vh1/24/h+qB4Il02ASvf1QytsTBrIElbyg+KftxZrgdN1OhNw
GfkLjp/8uCbCBFyOdpbgjc37Lyinod2xhP+BQscrcyn8i52EKcehZ3f0UwsDo4yL
YtC/RKhMk/CmXbEqpKcy49m+GYqvioL6YOpYw5tfakM7Ooa6UfORuAci7M4f3yBX
/5kyXEp87hSmj/+W9BmgOIEQ6n979cMEyAH/eypstW5yked7ann2FbPN1x6KtqxQ
W1FeJbk6UaPgEoyORuzezD0XlQ0HFudAGVn66tktxVN4L/H4xi4SPiy25vC26TCK
hQgBsaxJzetdCMvSA0V6dT1nz7ojUmRD+9E1mIAJLcy3X/xaI1N8QTrpgWqfsx7k
EKZH9GuNMUd02zAlYYFY6MRq+js8x05K9lrc/bQezkhnj8YwNca5C4Wv0vQUnSAH
FIorbJ2e8xMk2OegECb1E+LXeqLXpMQLhUBi+wpQnbwoJShhESgXJe7S5u7r7LkQ
s8OIb5cFbB5gKArRoYh+vPXFjyWeWOduhxjZyfVnO7Uxsa8tfrV1aavYkrkTls8x
741/VTZteDJpiKi+tBGxGCCWqeZqn+pLLVNC2BlX3Xhg1MHCWuRqKXJwZ4NtlrCC
xje/V88KDQW3C094UAYoRPWZQjOpdKFI7BjMbMuJezfh77j0cdPhzyzpIgpJeOc7
PjWU+9CSJU4d+iLWtbxOZAEX3Q9uVjUAqKi93WNs0o7ur7mN453w45mjeGU0jqKV
cWNIEOMrfS4BQP0Qtx1EeQp88nGM4tGBrT84nTF/de7deirivmf0YPw+yWYYLMXM
vwlbejsTvH9CjWluO+NLhYdP3wdXtCiFgHVLAfjtbsV4omcjGaZd6NJeMkhzpyBF
NDx69zS6C0Fx7aUnR8rkkCDdygTJjf41odpv3M0RWGIL9Bb026Sh6gVcl2dJvaUg
Njm1FWtKQbsmJuiGJjawuzfEhppprB9thaiJAmy/fy4+/eKjeL4D9XCOwXSPN7Y+
SC9H/VnetzWBAplx/WKNgB+6UV+a8q9oSV0naH23teThHESZSKaIfzL9OjT9G4dA
rxlI3ZroaYemjEiLeW0JtYv5n5vZ/6vsnfTx7Ky1zSjSkot6SwDAqGVPMxnzzrkZ
vWxfFj5MfU6bFp9SnPpXm8mT2OVod3dmS6FY43cQIwcbmyG8j1t9WZ7N4bGLrICa
fjpaoE1mtchlYCvpzwzZwsuhK+7z+N6lVuGrHL0RjiVSRfO60XUDEiQIr1oNKD50
zMqwxQksnNcJkoPTEqreHBLay8UAa+2qzuvFEtKu2OAVp2s1SyJuMNjc91DHW3XA
HSjUtUc2nQVYf1Uod0srEw64Z0YCbkgnm7+i2Zv95nNle0TEfqb/jUQNgElhklS/
NSj4xEiZi0MdxhZ02aZq8UF2OH5+BSfDS/JbfaXaRwSVvsQ8myeTClW+VIo0iRaL
ElGeJaF5t1jXEzt62YV9FDqFKRWgn5A8Q7TtL9Fz/h5w66zvpMBGhmuYf4fpWIBJ
Taf0GMUaPpDCC5BxKijRZlilgbhcyFId5IToqeSAInf3RETGT33AdYzg51IjiKG/
ZD6+pTwU+5cK5+m+IB/5sRTCK6kVqAtUNcw4eaDhMuGrNfcegpSRo9wtsqFcVYlV
gpt1YJpji9PTcbyNEKkYAkk0Acn/UpR5E9ycqgPQoWsdZIrzGMgFZD2Mspj2Bs8N
vOVa+XnneRPWOtBMacyekGNlP2HlVgs7DVIPgNWx7w7okH9OjQkf66p5eFoZ0jd5
8yUiVZfwPjbXSqy6B3wOMpQalNx+SoupKVbsDS8b4pK+eLIOQkIfJNS9Ctn+oPbk
8eVOet1Li4GT0sLTlbxuE7CZaf2RSxlAt0H+nnj4/+RrCy5j61tUBLMGWghCc6NZ
oFHAbYC3UTEH6NjdGkPi9bdga8bvM2XCq/HZ+f+UVgTIQK+giusbashMg43hYOvz
J4jb/r6omKeMysyh7/OiHAtUOdtCOTROChfmzXm6LOZ581pP64/IFzfUy3MRynzG
29NfE9kLpWKkTWpwmTHOWL89PPCe57SEIeXObYC740sOhOq5h9owZzHsX9JQwGkb
JV4hBOQcihLwub9xqxaeOSviK9n9zGm30W5LKBDCe7FirQ0xS9rghA9SJ9p62/vX
mfjSxJfO8DHYPbd2dD1VRe1HOXU3dGwZe+sg5T5c+XsPAGaiKIFkreUwUs2EKLeo
/G1gcRTIkBwGV++RZSHBdQHr4OLfbOWx6P4xzEWMePSt+rR5kuFUYQQnVoYZfK/X
QxNxPJx5li2iMs44seABSPiaYatKE8w0YnksufV2KlSr8QLK7OeuQ/+5EThh6JEp
GtdX92j7tD1JhoFVttQ1Fdi8DZNZX4fa4J43+P4JkLJ3Z4MHq/le3M6wyXiVvmhC
aoMJkAP+N7weKjTrXUSkSjgN1gs0Tb8n1XooO4kmy+O23nytzKUNP53rKwrFLiyE
bOTR/YBfsPj8JRCkSeijhf4ViXLIrwkl41knvSY/AmXixdMHdojPPGvPQwZYW502
BTyK5MvLKmzKbSEgEEPQQ55eEq8ss9e0bUD02h9BMQbXFcypc+uQeB2JZCWJmlnm
uIz38zXjq9Pt/3SYeAGeWduYTtp/gJt3+FRDjpfp1rVVklNPumNY5U/zVcLQ9fWB
2uG3r0RQ5YIclQYSrQsCXBKYZj+JqyODA4bW2+vlqpXKD0hnL0WJu9RLn8kOdFxY
oPRirq5yaPWac94zVVOcmcIB3OHruV/4NMjot1wtuIjImGw4N0CyFdVnR/TVRPKH
EVH6noPAOZqF1fuTfIYvaKX7wGxKiK2+b7Ud4paK89L3qvr6Cal+0uxp6GcWkI2B
Jub7OeSnUdpfaq0XBcPpe682djSaOPBHSn5NfBqP6NoYIjl0fYIRY7e0rvkvncfJ
r1vTYWgqgESk/bLUL7JuCwUu1PnONHalUVUXLy0L5XmJiZwFIQe8IJRLMt3Z8AaD
/NzVX7WPL8wlFAokFmWShQWub2yl4vkirwkVc+pu+NKi0ZSmfIhOI7rrAyoOipS4
bExifvq6XgqbhmaL0voLUIqrrxaYLdOs0HOEadaRiDp6QZVdfX8F1lxU/arz4cqj
o6Cw6WAN2aV4FWKwK6qA9rN0Cev1KrXSsU47IG2VioVdksjfAK4I/Z6eiGFg0dxm
gULFjvjcGtHuN2OzpO00I8XbdgwdW2JjiZk4QrWD5X1Gyo1M3cRsgxZW1BZUbIP4
izilxjgblgnBuHWr6U698BzzmLLIjcXUzmkSZmryPkMvRIlpXW1rdOX+gaYUQEDt
tl5Q+M9CFuw0H1iqUtL4M3naKknAal/7iDkTAKXbYEd9R5yQkqiLGt3Pd9AJ0wzb
HOUJxUXhY4+OCuxAp9bGQ+r4qM/uCHivPK8onUsTx9QO0WxNmTnUxZdRO+qsh/Cg
88z8YI9cJibrFJJnlt/7ZB/5cEvaYr/4YzWqKQLjvh6J8TjXns4w9CElA8cUMRod
rxewP4OW2nysIvCDeHW1VzaC3p95OKx4j97WZ4LhYMajXvArmDC+skevjrJ+Xdyk
vy7u8eDrQTuozOCud9BsUd5C+UakFI5lEtZOVWkojM5y40wRc1CUmNobbfrhvW5w
McQCEmMNd4BfkkboNyWQpZ20RTJS86aGvNPwEtU9HgaRg1ifg20Pn0TSMg4t0EGW
auFjuqdgI+/LWDFOUesKVhhmloLj5Lgdlcqca7uOziqdebDErjZGYjoQarrCRBYA
al2onSEqBmxuI7qWwWvU/n9fG6mWRPnOwZO41+6aJilV5/aMpr0O5rza1eLiV1p0
OAuEOPynca4NpIcoy8hdWcpBnpZRBiFe0Fohh0HztVnNlz3SuES7A4w/865tq7kZ
0ZLiio9BRz42Xt2gU+rSJlwbGdtOtQPEjcNV9Gy7EdC2GSccLywU1V6bZ/+9hRci
N5EZUW3fB7Gb0MuW7AVCAfZwIJhpOT4S00dZsW5Rip74btn/o6jEWqAhcwC+kz5+
KNcX7F+wwBFiu81bmimPEaCwU/vl0uY8TM59JjCz/Lqc4Nl1O78DZ5zu2BDDasKf
cLXbfBbTeEeJ6v81z23Gi5ZXmRtBJ3Jl5PPR+7M7Ag7LZF2XPqGbrlruKuj7wBI8
/ZvqnUBy5hzskZpJhxfpHk0UNkExFZyuKBFSWgBWi5bq4YIY4mQiZ/ZoNFIMQxbs
S+GJhhf2yzfIRqYyUVJBPoxBmJlZJGLd1c41+woFIzKws1a03lhDwJHBwAnmtqoA
8D1/Slu8U1QZTyGke1ozayBkgqlp/rvrJUWli/x++DF9ezxVJ7/Rvqbj5hC81f4h
xetX7PKLpgGS/J2PSwVt+vzwytkUcZX99V/SBxgIoH2OgaLYgj3unzpbAdE2OpqQ
wp9PuFSPnx3nNilNKxzIZm6NZmpgBBH+2uN0MzQgXkO9Wb08qvxSGGvqcem8cNPa
+Cz5c5WpHYSASEnhgswBwGXo6OMeF1I4d+VJTnWfePRgx4bTCYymzxcEcrenKSVk
vmI7FTlnSYJNl3if6zF/xhQTx8D3bc/T0cl6BRsA0ckNc72FEeK2HWj34kiw3+Hq
7Lzp6GBF4OfAuI3dXLa6S84iMGN4qKhSDQqBQJK6rOKxutV7Flb93ROFPgk/KfsQ
Qqn7UCGKQbG6izKFdeRQ89VrwMRkTvlyQ/qcpnaUhRuVlYcPcVEiRjWkpgcrreNN
N3ThYjU11tnEAEEGk0s3rChh5DUgjM9mHP2JvIewpxN64Me/DXQ39DzCCX4YcYKJ
1jJCoASHn07aiNCKebmuGPu/lEsZ9Bv3tCYbeb6Sb1htSCETn4lllk6YmqN0aSPb
X3w/nhVriJ3HFCpo5vTEKda/CXT2WYRxKi6NAb8tAnZx2kbQPAPA1j31qiAShSVX
gkiPd/JJhYvcmKczaSQ1lkwtDKhwUGPdifovTYxbOqSUptvfsAUe/YY/BgN0hjts
LTZqPN+ndILeIufEIh2bGJJ8ul62XeCpf12yz7cxRpBy7hx6xdaSD0V3UzDK1gdW
PDVkSJ8XY6bYuzCXzhWCLa1LxtDcSDI2CDs/8be24sikTObnpDXnVr9rTrthaTJT
Zhk81T3cB7aaTGVH2LnywV1s4I/06TM4EMImCJR27Z3Y+bzIa5LTesZNwZaJ5sV9
Ujq3ECrw/4bCXMQTQoVT21qPXvTS2fucfvqLjTeIaK13L/qXvksPZplEojGVvnJh
/0ajDMZbInfMt4UiJ7lICUYmRHIqaCQ+fiJRXOwPH0tmfGIMZIHozJsVQIjUkFtp
7LE8/JIn/NRPWkTazT3as5tQz/w1eciYfHozur4dFB0VLgM/o40gUyBjSsvxz8mY
`protect end_protected