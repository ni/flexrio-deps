`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3328 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
ZIICkMu+S2rq/yOQyqhpujIRIfAH4yskBOkn5X0mi+tUc+IHM8Rt9JWDm+i/6XIM
w3LnnXXtL5vOS/DxcSGP1RA7CUJlBSsRyG7Yf/EUWV5Xr4ooRksRDErSQDhPuV0L
CDFrokP6QdE4vPqCMzxF8TojGzHLWzIl2W1i6rROt4mZ7YyY2WK0gE/pLyGmCJz8
RC6TnS1ISKMw6d3yvomo3ngw/JXloWZctqlIHcLu9R9ils0knKe5ITjRVqgQfyKU
bgn7tVw1CFGUuqRFoeBrlKkwpEX2u3HZgWNRXcfxAbCeJQQK7tZ8oFOWLkt0Qlmi
RkWb79uWiqQ51GZzzZrk6kT7NvHl2Pu9rElf/I9atFaGbXWugQpoF4gJnoNw0PrV
z8lQYBbwL+cePHzvFauzgneBS11P+AU7hwwlMloYgx6ZLGf6XAnfA86zC/5iDlkE
RuVAcehKX9evRSIOicUwYGeRfS3/MMFQjs5xH/M+5h08BQ2DWH1xHMaFdBPrLuSZ
kVdxB2CQGtvJ4gGaYdjZutfENcj9C1L92AoT7SfndAFTDfAEPBTlOLP833zWXccP
EmIOh7w15B7SrALrToVndbjN6mAzYdK2bdkKN6z5LZUJPZkczhl7RIQIYw8/nSlp
xmFhic82b2OJCs6tWY1quo1OPjBXKlIqunXKfOOsFbrg4KApXS6dC9cGi3iyoxSS
gRo++ayG3HrZnr5bhS0dFYB4u4h1P3WjpL+WauUgWSuOoarhSg12UXRkbmI2d4Cw
F/Gp8H7cForGqelvgLHYVpLIiwL0B123uPnXtakfhqoHSt0Amu6sVEqIXGBRwsmG
Ihx8JIxbHv/hoVLUBUZIfZ6qTOyTxtnLm838FnouxjCtJZ3UGF39sl9696+D1Fa/
GMemsiAMPeLHS8erANycsd+JrpwqEcrRz2xUNxqWtX9AvCD5ZV6427C13EjKnDdX
NL/4pW0z60VoImK1HeqG0Dg7CNzRN//+VUFXEwabsY0ZlxySV5IL1SJtfuEj/Jqa
SmmSqahs/7klsnFg/a0NPPhX6HOEaE1Y/PQG9fRXUfH0KVBKbc+fxo+4XHyHpqtI
qxc3+TZpT1OBeFaw1GMUwsLC3jkjbk59GLEvdtr13xAeS3R5zFTgYzXdXD1njeAT
FmLb+ktKjz4MqKEkgV1GDHYpVH59BhnPIRdve2XDW4hvP0SVM9bMULG6CxkjiwTC
tVxvQWnTk/jNajbzro+/3Mz2AGn5Epp0b8VxOTq7fHmT5MSTxNiVgKkF89LljQ1A
karkzp9Y/IumaPnPhwcwEqivGdGgbLHNh/c/nypjMGEfti2/1V1z2av6lA6Ub1kF
ODPFl5Am/N7Gz8g01cLGK2DCLrN6WBqL7PbAmgPxNslkRpc5Y6OJ2PEsamrcDR3/
ddHrxliw/HwYh0sCZqs0Ef4ZE2n+dOYdHjnsgsYbCko329TaA62at2KUbQEF0IWn
ieIPAfaf6Vr7uZfTilZ37UqFE9qMVyrAzrFLDHJ/TKYfu+MEPlEoutKkSm1cNJ2f
Xtxjkkl8mGV36/VkQOkKgFggjdiu49A1HTje5ASPdSCKCI2ShCo0/TisjWDqVyoS
5e0qczBZ5kUruttKdHj+ARWiF7HiHaKYFbPvvSVJRLzkfQ5VpaqoA3RxeH0g/csj
SFccr+n/n8CAhsLvucju4HdBG5z6Jl9kkF3E1fdgtDUMCP1i7UIgNlxGzrwyJVth
wNc8hbonEXbAAaoURB06jI6NLarx6fjgYDCY2fjYrEKDfTwmsRjl/Hy5DHFOtdlk
Zjn70PN0lhGc8cAFNEb8nB9bMDJTwnK8IXSwrEaQIs4W9c/9R4bzERKsDc7+iPNC
TjiE5BEqquIE0nWVI8NR9S3PooYCk7CUJFpMXt5mv64oM4a6nLd3U+jsUF4XL3Em
xG/coSqnvEganTUDBOXtK66NcgzVOg2LpDKRwprUJumOrcsc7sq0IcPjQN2f9vWz
+Rq60VMAyqDaxfZWXVDeMdaQOdI4sjOAi3xq6b3PsIBi39yXTDFIyMYPIF0006nR
JrcHLhMpy/ZI8RQccWSVzZZJtCnoSACYC1+rsrveSx3ERJDQt2VFYkm0uEMjV8vi
R1MZzxzoPXYCyW66KmE/HjSDL44LhzVRo7uT7w9OgrFaJCQT/5gBsdxkCc4rVCjU
3fq3qJdisDS62Va6c2FaA0uh2L0oNi1EpMzR19tkadbHZsWTdMLNojrkFIxwbdV9
D2qNGytp7vXdqdjJK86D8t4FHIZ4HrQHEi3ZAp6YRXSod6A1Jbyl4Yiefrdiiljq
ssTsJMcVfijHdqXCTxoeNr7ClB/nWJ3HBlZlHn2EYul9WctjJGxC+6QHzOxFBx1S
cdF8VOesbCpKfFDD2ux/cAUPNt4oDIFQxAs+4T62bPUq/mC2aX6Wy1GCf6v8ZfoC
sgm61i9BvVudtppvj/jt4iezM0Bo3nXHwFo6UHmqvL1ktCOL+79WgPLX7NOxYokY
VPFB/jIgTGXvmzYYp8K0Zvj1bZVcSS1YaQoN34MvgiySOO85B3f+vPTLpHs8heAI
7SHe443JVsb4C65v+/0mmnAxbAmzNUD8c3W6ad7iqzNE9i2upwRsMAp2hTUvKzft
AXMi5ZvxtY2d0IdqvX9VU2fk/wA00VzAMLnmy75aG6NR+W53uNPZgwHtmORWD66z
LrnCB0/YKgcKmme3cKC90bf/KFs3ANddIK1r6Qpiy6BbmmpM/JRoNDCWZkDCnxZ1
rpTClJPzkPrTsotZQC/4y72F3g2P035KLJMAeUlJtANzdxkEhocd+8vIwxYJazLY
sYC0dkyN2FG+Ew2QR4sglSdkdibdV6T8rXAFmUE8X9FH0BUF6xn0HN0450m5GyFQ
tQAf+yn03c3uiGDMOd/1d3XCWwcX6pOC//gbXryMJYMFEuFkxV/2jDh/zKHKJLfh
rU1bRx2RI0jJton7jUM58It0OPhHo510Zj5+227SuO8WtN0twd6HwDWvqIRzK1+N
TJoX8jbwgcLFW8lFkwlBjsfyN0oteM0cDLarcNGFT54boNyJ5vUEhXdiYUs3uDGc
t6W0QC6qbGmzs8GpgNiKFmeMGS8iL8D5yXBtZvi1xIC6BRNlMYq8NI2xky51eaUg
Es4bkxDp1Z+UlQOSRwJCflsDbYoUzzYy1LycDMEuri0NAcd1Q3EhflzzHlHfKMP4
wRoKwzbvxbeYapDyav4Jlf/Vv8hTVp1ECJjvNx7/3SWXck28yRQWDdHtbkd5K/59
TPskzISadk+28sBbDGDz4IgD3U7bj/5r5S298/g9+BmOGpEf20ddVoN+7VxPL3JZ
+8WqPbLxcRFab1eK92tcMDRUdykd9+XgEY/WOluNHurt09ziEACNYjXejyIFrKfw
MYiDDfjKnziWLPeV0TfxB9/NLK9ftUcS1SR0UG6WcRJTUGTOzvTpmr+m/oRP1VuU
wYJnevyEDGQ465SsZtQ25bYf/qTZP6rRCmbyzb9obawCER0KFO9jUpvnoDvhdsNG
e3713IFkoZgeb5owRbC6ZT9n7f/nb7fCiYhvvftrylLwAadHt6nu+imUYJi2FAG4
GIDAbbDqGViMp8QzTnhT49bc/j405H7md2WkdwxRYvggG/WBmD+HKjPKpIm6OCav
A3nSMlwNyqffOmZ4v5GNJdTEUEY//Zkug9vsWBzvlEoSkxFMapTalllFhT6+4ik1
rKUQbLg+iHUbYI7SEHCv2z2VAaqFnEtri2RbG+BVNGCHNmtpigoM2wIcI9mB1ipJ
Ui9CUvnPqbaMuKc6SP5ARlwQOtejQYmtNmJeVyb4Dz2uIeXWuvXifaSAk6/ILabB
ytCdAQqpVlS/ibAe/9r1sd2zlyZ/M6a2+m6Cwo26wxEkPo1wjXRKuFkcUfCTceSb
EKjVf2WsLF/+C0qNdy2bLr8vW7e9kepA6ajCmwIBoHBbNbcnNBHdJEj4POlkv46W
+zSkABDqQ/GzNOmuFZW9tig8uXlBKSOAQtBO7FAKJl2LMOboR3BrMjTJBdEiFHKY
dIo7cFRGrYTr4KKAax/Rnq1bT50cdN7oyO62UnBN5tTcIDQ6LcokkAv+Y6uiEND/
wiWPqJIs5AawlvKheRdhuB9M+ENfMDO7Gwp/Q0e5CEHEeL6vnV4wyEoNSrmcqqXq
xAkTLwSYL99QHLdtC1awl4YHm/+7/ecqV/xkgehNGEmEVXO8WmpbAEOPprANNdcm
TUV4PqkpjjhtxCtCye726wvAdVuSNQu4aGOnjS3VCF9tORKMafLMDAMTWLlsvZ1C
M1D4Y1QReQ2rnY0XHkIPRw==
`protect end_protected