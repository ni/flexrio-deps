`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 45040 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
gjQxfoUVC1+c91Q8h6upBg0vq44cZWSKgf1SozrjjBF04+DXjV7bb7E0mk5FBAOd
7gJGq0rVj1aW28oQNAKD4iHs/7Q+ZEzw+Z5r3TbhE8Mo5Ueg4AsDMjjXCcHKePK/
fasHhlaA2f5Y7jwffmSr3Ns4SrwMla1F+4M5JXYIOg1lvtiQHP0ypySKoPyMZgHx
tO3rmNwcc5ZEF9fL+4uI5EtII8f+miLkLhkb2eZ/e2fiMil8vRwjPejgyVytfXv/
JBx7F11ee6R//HcyNyD5Qd98kuorDB28B/ptEtU4hfQVhKujAGdGlldCby1TBYuL
xMsAUqswFkmddDhkhHZwAItJPeZ0XTocluFxUcuehanp7UmuA3LxTXidRxUyoH7R
6QpSw8x4lDw2eg1mqs/PHmTPNq6wAlQdjalO8FVg7IPdAqsfntoeOtlLFXxBZQtm
OP3qN46TO6A4wfHoAj7CtaEL0UahZSu++HXICgDLACTg43CeHghZwqbCWgzbKr3h
0AAjFaoA9ZThObnSDZA3EM0acDqxNs6JbImBe2QbMjRLPG3fUwDCcCnMCH89/tsJ
yKsVTERdRlLdX+jSclLLRzdrofgnT/ljbFPogP7nMJjxEW9WH6qpj58HsJ7hIo/3
YBA7IWbFT6QaRAd/wAM5H+6OwRxc1c2qdSaValQOUzeVXtVfbFa406tnvJAvK7pv
lOLRQvG/wtgF8SNYHEbJ0kL2xALxUEnUmCtR9mF9606/NZAiHxfS6aPBBnOntzjy
oFZokClAO9jC/ZcD5UmmLMqqKZx7ZbEyi9HpG1bkokD12kaeVFT1pB9E7W4aMdNY
WnH1pRSN8xHhnN4ZnclpoIJgAYZlVF/SP1VLLi8Mfs/gXtoCIx3AbW87Bt3NtRhe
R9Aiual1vB9gcMY3Ea6QKXjVSg7QFibxvXRa5P0x8PM0FoIwl3TWdjtbKvKlcNn/
80tGYtwiv+aA0qf0fL+tRMcTu60P0Ea+6N7UTFSeuJ6DqpLhKk29S/XLPz9Mi3oW
eG4uC8CrlZHRhS3LU+vTjrzGwk60gsZzkTY2jaCso5ea+9qxW+C1acXDjVNOYH4Z
+aI0PeNbmLIuQzlESlwPgqbTl8eL7YK7nICYumddCew5dCp/4vTT+J8Sr5W/pYHp
zHN14eWmLmQV9MarvfF8ln8e9vDAkHy5lZ3RL1A9rSoH0PqQ7WjJO7w8/PnwytuQ
pERbnIAQhf474CNfX0BZ9PT87UYkdeB8+ol/SKkplki7pGohMeI0bqH8bIpIKL+6
uSd76I3CGUeW3+R8VwlcInxOhpJ6Q8huCC1sqP+hGQkCHfnS5CzZD6tGnxoBFcZr
boL8EKcocVzmLYUcBavvbrZWruq9WPOK6aCLsnXLSmgZcSL8Y7RnkCjHkrGrWVxo
MapMgt0icTw6uFvBMgfeL2FIO73spNRgy9NkSdYn8MS8heizvOYunZ1qaA45d/Yi
u34oAkeYzNj5l2+SUyHW9PlLVmXNTRCoE9Z6cQWsIJp8os2YYXr+cFvTRjheIeCR
xUTgjpePfBKshbDYwwiJEMM5JoTp4j3aEVL+qT2/sZjeBl03jSB3wZs5IEh5GVMx
FrzZw8GRFb62z13kBbyEVbg2M4n/vG5EVKjZsYSaxoG4JrqWZ/M9HTrLt9mQsiyp
hrC8exFQmpxHvSwPxlUbTEkxhuodozznlhW8MvmzYXp8N+6PeMkSOWoafxpGzlUi
iNzReZWwK1iv3yfTnfvyXX7FPOHhLuU7eTAEU1RJGGDt1OEo5A9kDs4EubtTr/4I
Re0GmCs1m8OinLFIJ3uWTdL/795QZGY1nwj3m3dRtzrCT0v5h77KkJPqfqS4N/6p
TgogjCXts/MusjPTf4gXMeB5x8O73Eaw7iJOjaAc0zowcqD5Pmtih5/DLgXFNF5f
+UBRuit3R1+j4Io+KyT8WCN3IAsIjNToLfJ8ZzIFpQpTcD6FQaQ8i7Vc6q8ePxyg
JzGdiyFiTYlPam+/gAwR81NoP7CdP3VQenDiEV4B65x7UsvMxnweBIRI1CvIFdx5
QtWB6lngT6XmF7AJraY07Jt+u0laxTibVyji0c7JCDi2CeejVOdifTiciH6RS81T
SNqz9Pf/FaH4iMH9iMvNc2fuXjgONk8z3sfeEHa+M5aJB5hcgcoa9STpVU0ggwrU
63oICllQSXAcwMo3pbqyAwZ9HtMOyC51Ts9PKmQ4oSTkTsWQn4bfi34zMz1bQEED
MrxVNPOididmAZiD1oPnKZ3ADXcJvow//1Vo1x/yWyEv4zrKrguISHtecSjvDpKu
YwfUz9E4slj7F14A5UWNqF28C+U20pScaLG5QpaJ5EkjWxTCzD9yEXTp6/zamstn
Zzo09MOGbM5Ce7AaAfZpvficgynGBP4jq177iT06uIzP8zMJKplFnhSR8xjO+oXO
2XBIsz6X7UaMLoXyF5WpqyLm9Qu47OqpTTkxNNlqIpxxfigFhQg+SW6mYnX1snKl
3ImI4UxZttK7K9Lh2o5rfcpQKY43lyVc6qbr20IqOSuei271L2UiHEFDpY69SvYV
oibaPN4Mq2DqS8Ffu0fRN8M5zeoi9hT/8Hmua0BH1oh9ujLZoaoasX/CwleQakri
h4Z6+C9S/mGyRkJoMA54qhW3CSbtdYM39icKsAneYPLJk//wabxighNmLRgOru/z
jQeDXkpkzjhAW17ONrPoBaa1dsfETAXec93fshSDL+vQxlKYY0a8taTuuEwS9l0x
0mZHOs5IDU6RVLU4sDU7fUsKSghCfLfd7XA6APl7kQMMlg0z1THJHztA+764Lw3p
+7THn2zRHF4awR77N53U47c3uVhciqq7AzvuCWOetyyZKuoQMTRaJN1MXUHwwGjl
GaukQZDuQhZ0kK9xG7zufEwHGK1fps6m3e2Sn0dKwT9PjVOtO5BXy0gg5AvC+Yfc
8JiD3eGNkyeNK7V9vHCX77mfsh0hi1PW1PTCS6p/DMxn3+b9UuvhG50xzdWOJd3g
qqRtj19x0v19PHszlyPOnWPuqAGA2FkB+OwTeUSFAu8ftMeA3g3iN+QEFqGHxtGG
angviF027rLPBp6jP0PgI8WRDEt+7+hQGJ1Vd5iT5IsFvqHVpJT3CuGdsNBM9ekb
1c/GL7P5xucRtwr0mRIF7yBIJ6P2r8Y5kfR+ix9phbMt83C2L4S/uaE4xclzfu4K
W4ZX8Tc5Ab56MIHGBmVIS9qv+zYBOr7K0gVASOkv3oRB6tjIhcPldOX2HUmUnQIB
kn4ihBaAUjXFgw4hiB8UuKnugADyR48OSYlj5c/Tn/N1iOW8/onITnnOXhMh2WKF
9pB+Xd4jHp4r1roaaPoTumR5XdXbdMJrTTwXUGxU0UKSoCNMWwkKj6ituAQD7iFU
hMBzAaTEVSVXpeHL/MTO3vQi7pQqIkRmtHbQSU1dDltp1f8Cqx7QkGrBukZThIQ+
shkvTbWPfUhH9to6PPm4IXq1w6ElkholSeVJwKBY3f0g0JVl4EewAHQe96EYWRnJ
HAR+SECh9HZQQaKJ52x9XdbM/Kyw1IpknthC7yoIAPIySgZrAQ3V4NGAHMmNeOBh
6hYVgaf2kUShR3RKG0cSDPyJACymmoUW+z2XMywIwsO2/TnS6kWu3sD0Bs89AaTQ
ueYdi0hkXTWbtNCmGL/HB2pMEn5BctWjTp+/0OJewbMtJrgAFczbe56sZZu2yuZb
QtV10DP7JfjODVYvxm5fMStrYbrcFsFayCmLjcZ3+h+8TWLFHi8loAw4ulzeUjmO
eTr52g5K2DJXlrZLv9hBETqtVqszUdsRrrOIQt4BRoJf5XcenI/lOJMwDev3uqtB
FVhaXL2EscS1iTrwHYeAgKEJLUBDeHNhyKS8VDJDj0qBQg022Clj+xACZIgE73Vx
69tH1nK1iCt25NXFWGyMif/GavxuB3ddDaTZ+DqtjZCacNin3FvoOoUSE+yGrKXS
qNTUQfemYmsNqv9q/1/tfuPhmsJZsPcTb1+pL/j0kHNrPaxWRZ4S1O/xLMt/kgCo
qUYeNsX+BHBIQYPjW9wFUDkrF58s3k5X+IjX51JgN7AELrSRpCvs4b6YKI4ZEXPj
YIvKlTneap6r9C0AHk/m7zdP217F/23bYvOA9qEsG8830figXU2VVjq602ezfMH2
gy1YNgMw2eDGCDHGL8h5jzF7+S9dCdgv6MkqcibRW4eY6TD8XmYpyZyyCPTbBkpg
o7oG0DSvNVUzQaMn+6FQWC8GJaNyG9f+USUflYFLHsjVvwm3woWlkrXebQr72nb/
vEtxBss1qtttPZGxT5slJVy8ctRn0warrk3O29sWUKKi9EDxMtRCBTL14FngAYxu
CdpWHXPwdTCY2f0EBX2hDo3U87faIOgV7aN83rNqMcgMzOMSd1sayLn9clpb6Jb8
HMobO3HD8Z0VGD5xl83uC9vDkIPcX5oapAEPnvc+2wAQmhs4RsHWMfj3PqOD8aL6
vim4AODh2Fye3pd53V+zGiRUiAMjJBc6BUEIRIiESUwWiS8g4v1ypn+94ODuXrGw
mYRqvFwNX5qvBHmKGC6N+1YQxs0Yd4UpxzyYVvljtaN/S3L9rOOhl2Xs8eXzxFO9
pq5jnfFRgodNUuDptqqZjaJcvZhWvzT9Bvvv6pRoFi2BLwm5VVeMtRgeR/0kBQq6
VBpdUzwVAU+taXO+Q5SGIwDL//Nw+uWiLRDtBp8R9422mcLSY+xHEbnLnuPqlGIJ
K0jo9r9BdmYzQqq16BqzDwxWWRvbc2r3Wln7wZi1Zh0wUgq49tiuA8vIKpC+TZRh
Y8IGWfsLDLr31swdAcK/MjD0Z/q3DQ9kQeAXYawJJ9WRnsSo6dMbINR3OozgCbNm
w8/aJ+HzvlliCh5/g0i4CRQshd9Jr/k3qFYRGUjHaQNFoFSTlcw7URxZrLqTjNqV
3feNLG4j7HW0OQCH6qH3CASyzCUUjXcn2+06M5EqMTjbi3aLI5kQ3BPR6OaqKdRZ
KcQp2AG5WU6yhaYpLh30/zwhW+GogBjT/x21hefGwoKq9llC8kLLfK/RokB2eFiV
AKLy9bZ/id5ZAP8LTJpdlfz9s7JxkdkD0pNiJOCb1FmH2IBpC+xBm4M5gHK5SD4L
hrOD0kMdqKT/enNn9qhyEG1S//bVhaPyGGHVg7qOjo2YlPphnpGDaLwDNyrW4lhj
7kZEAlIDVGCWafv2t4J8xm3ROj/CLvuHkkql+awkWyjzYeaUDAXU8jUhOo/5yUqA
cuWEq7aw0APm0nJPPw0moff3+++hDg2lO0DLmC0FTj6pE3BjtIVLRdNX6g9El1C5
em2MYq+3+Df24hWumlZ0tqW5Xy0O28t375+a6jY5Ljr321VLRFaU0igSDQrqQ6Sd
cIyMNXZkES1DqzY17Ul9Zmx5uhD8tdoM3OmSt0lvfC2ytLyoOOf3akUGSbbQWrgE
IqSYMotMP6robHPuGzxoG4V4tAd/+FvOxz2HGk8AtEKl65LaF0zXQw0DIEGgP/l/
R0UFzRZP+zCksY9y7kkJ/fl1q3Dqnsc4uXdC8WWHfZcuNOAFRyVbCenoMMHEl/3q
+/TbbyY6vce5CBd//XoRcXRxEPE6MgL0981cDlcabrM0v+0aRNsd9GfsXUscwXgS
2Qx7xUCzSK/CLRDmbtXbRM/OYT+/HMz9umgTsae+UBbIkZcKizZE/ge53hW6UsVF
uTKBP51zJZIUJf58CMOo+hFjpM5ZKsEm9pVi5aYFCUNy2vVQjjnfVq1ikKdC3zvB
VEVZqCYOdDf6xz6DaMnJW+c/G5N0x3TFIp5RifnCzj6JFsdRMjO131S/6aOg6wFQ
HuY5yP8NFXu8rA2nTUTjDmRTpujkHnJrluzQ62t7AFulfEZiwaVu5gbG6YhhIZLj
mvNP6f/CZy2QQglmMlQoG74CGGY1H8Pjg0h9OnRSBA8yOkBcbWTMBvrXuWop3ktn
3YAOH2dNzSYhbuHT11/dzWzJIEri1X13OVkMc/IkalbYqmIaU8MYkTwutBAgM7Ci
6ZaVdj4C50fRBw0ZnB2kBfew2U2P8cdPLEGgEm43ZG0mYewAzn3PB5lLmCgCV3SA
bOrfmLjop62AkR+m8v2w4M6wUVtn6Xopg083R3L7ONou8i1to3iy5kOTosztaTgq
NPlE7o+KAYYwDossw3Uor3FdPqQEld63KS5KoX1wwvwYtwPmFSXx65CmFbXK/XYg
6w/kE+vZyU5sy5FiLHKB5SHDPOy2DVBGv5Dq2jA5rnL/FnXu9qzbD8A7qiOcMQtK
G6xYAFv4GfYaFSKp6TOTFLtYI7vZFhuUj1D7fo0MA59g1q/6Bja2dEgYJr6VHJug
brtzuJgWCnG3tZAoVrtwlu0KzMYO3Askdfgy4h2+V3XHWehmJ01x+Gj4X8LDVu9r
7b9OsJO4zGCjfepMzqLWLSalLo9XfpUdln19gJXbbeRQD7GsBOmhq9IckL9e6hLB
+FPd56dQvuYhuwkwGmJO4RvrXCJLcmfdrWwuyHZ8uqOmtiG3jzDuSChThxH/k28Q
Tk+Sl45o5/hMGyBQFwwH6w1H2xiDu+HleGM0sIQuskS7hHwBaKjw6dE4pv3TDTgr
MASvF/Vmb+35UTCD91bDgKYWgHv1SIkT2CU4MGCW/XWgECtGMmo+Z2IlZXjbammv
BMv41bqFTAZ5sMKzNLbqcUTB23FMFUkOJ0Fh3IA2+UfZEmIoG9giGH3iHBP6odHr
AAie09jomfsr2jn+hav6ar4P4nvdkY4HC9naBwcAwZZPmqqn4lxD3zG2A0mVBsTy
NSaxYmVWhlpRVqZwmFWFeNSgURKXFgXpqmwR/0n5F/vx1R39zDSN0OpLMPfeDB87
iwQrtzKFvBwk+PS3SXoCrlbpMSNhZ1Dwcwu0ZkYfFDUUjXoBY0fCRsPNbdzlXaWq
QwEh5CY+S7GpDQjrMtk0z1cgxOKx9R829W20huTXP+/FpbttQQ/HT4hnofPMJPwc
KkP0VRIdNFQ9N/0XRWD6Sbxm555KsQ169j8hsDwpMC834g3UBSQ/YWOCVNHC2AuS
IMKc6NP2cDM0IZYuo6tHiVnDQfE6UMWb6m9I+tTqaJarXrztgdR5v0t6ZQoeZYo8
Jr40k+v/ubcfqGIFib7eqfGxojMYm4lsCESdWKwSwfk8u6Y64TGjLRGCTBNTKQum
XelcH2ilDFdE6NMnSv5wGvYgsRMrNRVxPjqIokS/Yyxf9xZ+dCd6rWlPl0YPJwy3
BhpkU7Er3Wb2a2Ab8D+tDnQiT+jp3QRc1vSAsHvJE7uzBAwC12Kuuc/F8lkptUFf
Q8bmJ4Xo4Xa4i5M0iCVGtY6fSGuJzumpu31RKcKXNMV5Lx7K6Y6ngZgWahQwLeQR
zhK0rk15qS4knxVA+728jfwDXDLOhCzG/QgwuePGi6VPzfJn8bn2UdnZPvPy4p4X
eWftY5U9eVqaeBEPKTVI7McYufNUGuq7VIfZ473z2JkKU9ROBLt4FjWjSVcf8OVL
g2Ncwudcxvc1E9nMM0HhsWwAz4vyke0IiD1YlAguiboH1YTi94Ppq0bwea7rsoau
6ZDSr2LP005bBKQWmbs4ax6TIAkCyNY//NelCq/3yxPRa+q1je1oH+S++tbNFhCD
0FLP6rQOmTBvDMUm4tLM793bqdCHhrFAZvATDtMZa1zf8w6Ptncvx1Fq8EBSrjn4
gyxSaZfGeDbNcU3N3El5aEh3CCPz5BTvAOV0n8F5/5ycH+0DUY+lN2EiY53d66uw
0DGPNmwuWQFMtb0iWikN1BSlvhpwAzwGNM1mmFH7DTaexeogASQX1JYnKyMsgeqo
PomI7djvIuMkDlVO8+zDM9hjyQm0u8aCo9QMS8C+l7VgVcwZe+2rpSNU6BnoglDa
W/Kd6FIryvMuUA1giYq8+NCGTUwr6BK+IIb5n29vHoqcVLLoEqd1oSqWJYnwu/N8
afdcaKKtHLUB979mbSKlLA+aamLjCJkFf5RJa7gIem2fL1H9UnYRQC9q49SGYaKu
YzviQuEAM7HtMbcYWKzkrHE3mqBR7lyoCVv87npuX7gmOr72AZd5mTpKsXsGk/NL
hpmB4WsvVAeTUVkaUCU6P8eYxnR18WawXnXQaod86uEMcE3AWS6vts1NQE7cx0c4
hem9Ec8jSk/izSDlY+juhb4Et7oOh77Pgq1UnfOaGDANwNEi1QJ8R2pdGOyN2Nhu
5ZCHqceBU164qHWB00pOsGDzHuC2Mu1eWTk1H/BVSj+0F09eVFfMMASnBTefO+Cm
x2q6GOOp/KaVO6N9LXj9DGU8S/e4bkU7l7fFhpLZFYVv3P4sCIKFGKHgR4HrlFAF
0ZVfHH566MQuICLcYZj6+RS+ZTKQCkdwW3bCBDDVQ6A9i18E3dK3usZ3fk/3mz0L
1T40LsKxo/k+7+mhG6QWSh6P1rVtEt5Fk3GV3CfttIs3InrDaF1JEvFMlulaoLHF
5D5M5O3RDZqoxDrKKX8QVbTXqaN7ZXMQxTr+qDCuzOKY8nfXmis8PNEhqkP6WPGC
OBqgS6R6TL98szN+wrNU9x3WKfd5dbYcwkEiQddTvrlL3kMssFrQGMRxsNhuAww/
ADGy63USXnNGMRI/uDHAoWzivcMv0bnbe3Mf0a9APH9B7HC2vO2S3hDz0mhYaXI2
4HJfkQwB+/UPu0MfpjtUbvlW9zrkLPV//PgeFujGABI8FqpkJQjkYGyUOTp4DiAv
Hb3XFpwMjVyRZhM4+DuJGQKuCyKx4ngkevLmbEK09X9TW1ji1TQe76I9F+JUuoQ/
NZKuT82dZPn+9Xm7hHdpsPAocBm1nnSeSA6VhO7GtH4qBtCxqHoh84Xoh67o/c1q
jDZG3ptLTR74lyurQzYz5G0Ah3tQe2AuppN3e8N8qBUtR02A8O93vQQUmdzhpk6t
crQHmTSKAYvmPHyOSmncGUns9r9fEH8XEH1mPcPHdOr/wW+1bYHHpG0V3R4TAn+E
Fuf8q0ZbjQIFmoZxR+4AgcS68wJJVoPGpNiPRcpRiE8covnOjfC7UBoWPC84ZRjE
VWv9XSzepEUCd3w3Mr575JagA7bQ/qCcNwQjQqRS7uRZ+tvESmKemaVWvJz7pkxT
EotYgvODnRmpia8UhZNmsMDiiUwkEccqq7n3AvSn++ujqR4ys+AxHq7/L4G8XYye
jDIq0QA6LvPEz/+z+p6oqXFqausvZ1FUKJMptlg5/QsiheghttneehJRr/JCOL3k
lJtZfOmpZY60w/HEl2eGzHkwgPqWgb47w5k7tGBxGUAbPbiuEjU/ucf2Z6TIVniC
1OouUP6DehXjy+nApV/IVfPD9QnTySwy+QNf5JfL8yRY1gQ03nR7lyj2qeOEZZN8
TMC0Ox7HqL5IJgRt52j+DkLyTLwF5BwpyzFNmv5wEwsJ2FOcif5XZF0qjhR8zLQh
NFHGSl5XY9s25dUAdZzceE+H6PtXA+DCEnk/rSPL053Mz3+QxOIvfbdO9731L6oG
UGpwDYCIOW7f1MhvJcSaMh4mYp6pwL95T3sstfnEvH0Vi4u2yxLc9+9ahGP1//4o
Uj0DzEQPHxQBTcTuX5qxygcuzoWqZWfCgxXn6I5poeoicBFsKgybYiH31w3bN8Df
GiHzLFHdpTPOfgF2MqWSBOZoO7sSPYXp6LqJsiA/H4VXTKoUrLSFGpeJ+C+n9vOg
ccx1rud9Q18Wct58oFr6zLkWrDU1FCFxfVRqMGGPXIUSCc2eBp0eGDvTsqRBK3N2
06I4dfu9r39wPRk3ghZfUTyiWkUg9Hiso7baj+SutCdbv/hqL2VYO8t1349XsPA3
NPgGOPIjAO+pYGzM9cUalWB8JEGmoPhFb9koHWli+ZBiCqokQ8hiqGjDB+RQ9VuT
BmRcU5tuzSDaZ04L2qJgCfBMeWako8sMy2On+r0HpPJU0oH6nJclUyU2BFigBo1x
4C0ceMoFj+V7G0KMemySSnFQldngd1ND7y5gDBTAFgRN7B9hUHspWN0O0HHXTNJo
GW4JICB7kviA9f/fYfTZjegcc88tblEVvEs5DvhscxiQs7+x8z4CIwKOQoMZE172
MikQfYx+GHYTNjoRAFeYbjrhhEhdkKOj0L+YyNtZfauhEt51kfOmbX0OP55AGckw
Y+aBx68ka/B/77Kj3OhzQeq5J/FcDl+RMg3NJ0Cc8zCoqsJbyS092vPkRKEDCUxv
jsL3E+EvU9mu03NGUeANXalS3Kuc9ASBKNHREwSJA7IARicC+zTQuCEmD5RFxQ4C
gC2AGeZczp0TD6LvgN/ydKym1iqT6twDn8LWhLxxoVnTY0SQccbvf0RvbesqIrsO
XecDaZMFRO6Tx2o+dtGFUF1Q6HjuX4BdEJi6ussKPIeHNpQpNTwfn0BoAG3wK+l3
Vw2EfvRrOsGLzLHhN8kPKjIcyQ78cVmIwklLYVH1+a2HJu/9PELq5G8/My0bVsyS
xSdfkIozCmnURytjtB0515BRN4B7fO1KRSc9O6/rj5ebmI5gKd9wyeHdvMfnG04w
+DlOowVFllPGHmXtBaH7Il+/VOv4yM5ExbVBJZTbwEsXzYczwBN7m7gtsSAZcg+e
uRxiUUOIdw3DFRNbdoGjZfPsv3+hZ+Oef7hvD4nyTgW0m9SRto9vg5ZIrE8rJ8DB
wmC0HbmbZo2fjaIEwPZ8iD0JTFyr6xUT12SdZfvlodNr4nsZV6Ue8mWSgObNIa2z
VvGTw1Ln01mNE53gZLa3GbhnfaLgr+d0rOS6QimnfWobmejysxE1tIzbOMtPTU4n
W2u78hEec5zx8Mp35oIR65vGqUDEBpD9VUb8IaT/KDzXlSMCk+JCMgQyNS96riTZ
oAE35108+mE9S8ruDtiPmF25h0DjRSKLa/bqyImh4dkxiKB+3Sl7/8T2956EIgeK
uMi/EBvWmk8NO1CzYZkoRlePO7xNCMSNGtlHKlb/yqCbTJAe04gN5858H95H2Dt4
5v0XXU89S7ZfasRlANkd7Kve9UUbLdH/+Sff1XL3XK21TIZ1LDKfBKlpuF6qzlUC
3Vjovi/lXWGwwtJwUy1i5mxi8v40+I1nvv3YMTMWd4Rb0GbiYiCr2qKAV7DPutG8
2QNPZWoAfwj9eYfPyNQ8ezno/wi3zG34FAUa9VXJfn83Cd0tvsXESyCcsZKO3Ex5
Tu5LGtlzalzlvHz4XYDbtQffBCyuszteBIK7cn8SQF4rZhKXfgKuqOCXC/VzMk8o
XcMWWPsXX8kH2Vtq2Amu8ZAp2mcplRcY/Mt2G8MM9VWFsbEXoWsPaer5FfUdLO5A
zoRDBh5IztnRjNwK7tDAuVW4MFI1z6hXEULySR9o1ga68ncfozEZWHR6EpREFzag
uOmGLcv31nSVMMj4hhntRx9eLO84Ev3h/3EwXJh5SsR+qPp2z5w8UAL01Bq1mrEs
TrPFRCIeKzxCnkqNt85r3NdA8XxfbfhXvvMVu5z1SSO9Y+zWazwB/8yCn9bq5LGT
+PLmqC1IQomgo81A5S45DQZX2C4zoe63w/grzIXMUENLvJ2Pnuje/md7DmagY32E
YJe7ROW2iNKM2ZYzPk/ySYO+jkiZUfu0GuPpXcuA1nnQ6qgnMWWfr8TYu2tfk9TE
rj+Yeph4G6o022Dwzn+0NhStPcUcHPGD21u+wKg295McSZk5EZlJxnDlEB6r1zjA
KlJ2XeZCb+sWRZ50NJakA44u+BwyuhNd8xkN3s4pD09aFKJunPYXGK2SS9w+3GJB
VyBdp6D0Ja3br/etssibxEF4hEMFTzFV/yuf9MZAvHzPvj+lg0z4/1duO3HRXRFl
FRwW3izR3gMs2SFKy1LkhqnuHvnXE8I+WOKwSVUjqTnIaUAlc8TXpMx3Y29WNar1
c8LL6tqEwHoOHF7CIYLE3StqpEpKGlVLEEZm5jZu2rRASapyMuB3oFWAhPHbSniO
cCU/ZUYUleHSzzqctz76X6AGWLTPP+nvOCIkBjl7XxFhKNxdc1e8nW3MuGBlMhD5
vr+tPRNvhoaNl/ZAPKGUS5hlZtDW4OYpY1WWgpq2jgwe+si/bnd53KoQBJ6758l3
ZW6f31dHbHPCOL/oZUB7I0q6SADvcXorGC97F9WSkFmzo5AssXCTHnx8VTI855qY
1K/3Nger+e/IajygoRyGGTPdbWzY338dICOqyj7oJgVD/fM7+6xZoqaiANJsgzhA
hgSKg3hoDkuShY9ULdNvTdlkm2Uu/QvN/e6h7iwDojbZHLA9deHh1aCf+eJsV4mA
B6hzEekwoHWuYB4k2MLEnLAHTHZjvRC2d1/vt6WYJwaazB8R8RgyE6yJLSJcGhwu
sMAODc+fma502/DaMXX58zFlwlNQUmvhaSRVC1vwmwjuJ37kuymLdAHnU0uFOXJN
VkxmiAEmQbpMJSKNRTEhAAyLXSTZ8xJ5Rgsxprng1SvzMtYQ+uvAy3zhm5WRCR/a
A42gEcFK9+2fcdvuH8tahd71nukdZgtstdkNC9RFlfK2HNF4HptpSawwGSvOZlc/
f1z/mBS3hUDF2KFy9kdDGD/wKv4ZQpDkIFfm1q3rDmLWOZjtnhDigpiSNtxI+mNj
j8dIYpeHkah0RqRNEU/0ugBp6Cz7e7jdYD9govshxcc0JLDSFmas4/xOUZ6tzkSJ
4PX7OTo1UYHEveA4oeFOsQO7tXnmz3nxBiQwZditmulLIjhul/09LuAiFXe9hlkj
EE8zahYlzcZ8cPXoLtLsIuBbLdGUdpXnQFb1Gh5Ym+xpOHGYHzGGLmtKJuCX+6b5
dG46Fqe8B1RXu2wRhrWRNDxoCRraSpEFfSObx6Tzwaggp/AsJwu2NkUp9RBjzeqv
VEYz2eXL11ZwEZwA+ExktY21MQP7AgiW3pdMbwcONWRqDZcC8Y9R7bkUnwf1jGoN
IKKLZT83PkHqkQYgUtW+ozmY4iCtDOUgXkHnvLAOqDQ+tVFxqX3lJl3dkMSfRfKb
f/yNjJObKIoIQZcknb8uojm9PQzzLSdIwmDJn6VSjMrw4dUgoDvPHlnOZL9OIiJf
ujSFfnKgs9wpDvdmTU50X9Dgp6RcE86YjlFv3ChWCyNvGGlnJ8jL94zgUA9uhqTQ
RsQz938e+Gt5FqIJWg77PJBZNW+RxDzsIaRJDFPB8BwUeSNTCeLXJotd9ZzVIj9c
5+DHPEL0lfiE/Pmasq30Cv7vBYqIl122B57va0RxF0LvQbSjJWEHFnvPWIfEMj9i
v5tAruQVwF/xmhxBRs0wSd07lOUTXzxJjWreAzGYB//8VHf/9cDQkdl7m69xDwGR
pOPQyOhr/ypLUSzeNcMravic2d25XCVi+ZKbtUVh+vH/WRMdeLfR2hKAKYT3F0f0
/O5bc390JB++4ptYzZSXZYEF/qaPqOL8i1JAgnmfC5hvJ90U32Y+61Rl7ivOA5FT
zs8ipkqs01ZvX5LHfFGr0CfH7BUN1Z9W7RYhwJlBDWPSuTWRnpCX3B8GEk3G3AqI
jbhIbfOGE53nAt/B/x9F8pUsu8j0cMoksjll/04fiM235lSdHF/3k3HxZ9W5MWW3
4AR+FukBfUb0Yj4e3f/gpuel+tIA3yA3ERKvQwfCzSF5XGmRxY/SW6Dm4HNXscEE
xfwN2ULN2/a+EB1HsYztbGI9o4pMUywnMKI62T8hpxltMxHMQmy7WG/knsX0Q5Q/
CTxKgWke/tG/ZGBsJUY6xwjNpGxvDXIxYMVHcqOXsq4spIs7oyBVDjr81ubNElP7
9a2PJIwb8nEN/ZnGVUgQjv2VFxrYGoE3anBrXUBpQdUFE0OAKoQhi56n9pHsutIR
FsTSv7vdPBWcGCAfCz5/1cfgAgCsqnoGsslObED69Y7cncjazg0TIRRsy9nOcOsu
NGG8aJSK/zZypWf3cE1F2k1fEQtWovpTDdlMzkdvuM1D5JCAYZgJF26jy/F9zodd
OQkdR9Er1Ublid9BucARbeMQhNHpzXhoNweDPbGNfGIcbqW98NiZYlh1CHCxh8/U
NvHnP7o7Td/vq8g26WisEdr7//icrY4CzZZnGRfLqW+XuYNHFAxmorBUCo3eVk9G
XDTHpuYjlY5x2ltoppjzt6z8+XpswDEGw7yqV/RXgRV30pI6ua4cTPxBT7xov0Id
6fhxzVzys3bj59IJHvvTxSx5EG1kpZFA6h2t28krgds0D3jl6atrh+YiU4zk9DvH
l471TH5uw2CU2O4b4Vlm7QGje0WsIhEZ7iL+UFoGiByiULC9Tb0FU594QicWNr5r
ew/C73fZLDimpkenghdEUu2b4zeWf3I9KQR7DoIWa+ibG/xir9xdhsU9eNKMh8KZ
aAV8ZyI9GJzP788A2g8kX/IX+digKvADus9hInmoB6cUtyll4QopSvA1NVtMl2/y
6ILYDzPUhwvN321k1Ukc2jLBEct1IlJVPwPTZewJOt6+yCiuAlMp9CQIzOECXTPP
+r2vs1RdBau4Wg6n99aQetwrogmZL4tsueWYqwS3moZjcv7JaqkyfJ83GGe0cS/V
Vzf31WPXup9ZHxX3S3GAluntZbbSd/uvNIFABKesWINcdabfK+ntwN66/oXJP1Bz
b2gl8es3WN42Psn6cLhgaxe8PA+8xHWVYVVOivSiYVDWp5cRkQofkX6IpL2sm22U
jOQMzdsyk2VE46as4r+NDrrjUBd5JTWsOXeLtriNfIYIE+6XzMSYu6NRCwQ0J2tb
ZgG72SuxFUNso3vMGUDj30+zvhio35VPTZNQ/LgBfhgfN7609Hwgf/RDfE+FH57u
XroG/csg3ozcAjhhncWckvdff9hR9iVF0iSxrmzp14GQ6YQRs8PjWYhawpyz7ecC
rls9iWpH612S7TSGmWXdgkwRBfKoxJrXWiFCetL3kxSofLzbUHx0HsvT0SHCxO8L
xh82i9P7I7Enr22XUunnu3qtmc01W4V9XV3TtF0OG2srN9T9TA1TdkAEJSI2s/GA
eSoBK+WKmZTA6J0lg6TvrmbrCpaIpz671XJIwBqDJ+RjJjhJZL3A1V6eWjCggp0L
xwA9p9eCA2qk/18QzccWXaesiFvsJwmO7NKDi9NytLPeofCycq89nuB/yMaSSVKN
1uJF+3xnNvzbFMk+wBg06/Q1skt6IqZd6Dzk22LzJzbp1ss+e2al9ea7/ZfECqyJ
9kZY1w9HKk55vjWmbGQ45LnC+usj53GJQiDuGTaihw6asc4hnCWJdXarMN9cMaYa
wkthfj0al88Y43z2KN1PEc3XwVrBBUXVEwgenag/86Pzv/fvNnEMw52rOQ/Twk9t
v9dpk4bnIm7m8q7Zyp5B6b2mfPr7NeZQ1NDNldbl/b8Av6ErAmHw4t51Gq3eeZm5
EcFmLNlRSA4ZSxBx29riFbhKGJiDSKr4mgYkUdOIT6mZg/p8eHvBH1YjDCEDXu20
9i8xpHj6HJ4xA7Lu6T32+8YuEKto5nvkkz6MbxJW76YtAza8H0dcqZ07c9Eg9OPO
SQuvfxLBWasRmnMomS3FCanyj1za6E5vHLxQSNm8meDmWAT/C9n48GEMyL/a3L0l
wBc4rIwTZ1KNHFtHSFppdJoXzctpJPZeJhdB1Yo7RwBWV1dnk3ZZhaQaOO+TvL/7
hk/3utMWsXJ/FX6uaBBGH67u/EY82k86Xwl4dJybq7xIfzfDrmrDN0RyRyYI9/+T
u8l0idsLh++1st6yw0DWQsfbjY6xULqS5VA7LHW1in/s4GzPZz4jTvDOdYtU6B0Z
3UjO7qmoNvI887k0hO8rh5F2zUKjByg05FdrOMynBsBQWMjVG/I8g83VRazJAb0T
UWFee4Dalk6M994PJXN0+0m6R1KzZv1xA6/jVDuToVyj6UEyXky+7O/7jORWOgPV
fY4YVdaVVnQneyTX3zoZkdDx9M7WLF2DufxNYjMVY+nQqvI9XM7TWget55A7ND51
gbwKgYK/nrOi4S8bGS8RLcyvdh9e5Za1QRZ1MjWAHTyruC1Vby+XviINTUDD6bWS
5ipqYwePantEVXQ2QiqSKkug3PWEB4Y/8XlvJbESoR+NG+UveDYYm/AAWUYdhfyS
LKiQhTEzTeRsKCYXcxY0ET9U8xR6yUFggisNFzlRqDdGhATYxTNjrzoi7qZP7u2m
TSXMrJir2u23HYo5k9nT4SY/gs8ldBrtMKam95Ytyt6S6lJaOr+oYgQpICOB/BoI
htKMixni6MT9JreIC8t69wsN83oYx/NUxnbtT//+Y2HeNPZYp/TGO58Q6TbZI9Na
GkGIlC3VM2Bu8AdjvAjBKQ8JMXCIgDGO4jcFVSCqv+GeGh4GGVELzpGuG4Yp2QIv
BYJLEd8Jy6j8ZNl8JlXJR3Lcjp5ZdCuX816tJGASQBh8YUQqWITEuey80tTw4oIw
tvzY8x4eSyR20887MXA3USn+NxFrZxptqEBVYvRaFXC1Swm/jjfWVym1tGLgrisP
JvZcuiD1i6hC6Sjb5nBQOR3DXyDudIJFZBSC+/TC6cjM/MkaeWxdrDICxKZyNFrg
xr1QfPIwv+gOl+H+7C5qlaavC0bFFe3PcgJnqe5DGwLAA1nWJ1InrnseoX1RKIE6
K5284KiEOFSuGXHcjku2bH+wArdbTfHnQ4GzheThSmLAA3fS6WR6Xw6iAv+XTXXQ
tt2MwavDlVOOiDmpY/tp1QQbSIp6QpQl6rYqQfK2H0en+HyTDdXHTjH7G8FfKYUr
JZBKPcB+uMXsVYnSIHPNhRNapwizvOqm/riLwNXU/VjtHJF+bAdjPyWRzh1g+H6o
lzkocfzsw1aKioJFHdI3/9nEaW20FY6fVxBvBC0ffH6dea4YJ5xkfjo+rvYrLiLy
UwHqlte5j666Vkx2SmCMBdT7PXPoTe/MTs/0El0slXwSDIx/7/1PtcJpopEPm6D6
sUKy+UU6bwakQRkAoGV4Htvt01/0ss//0JlhUqm0CAjpL+Bk+WhWHkBM32FZDChg
jrfZdNOcTHHBktFXFPggZ3aXX+J46qqPgBa9CKfizt4LMCvUeRRaV3ojlOYdwyrA
+7oCEw6bHUGXsPwPCXhPf6T+SCrU5BE6rAHnNI04a6VLQ/XjBO1z9rDZXmZDa3K8
xlr5MszoQMSk71W/IVTi6+6HWF7w5VP+8L/nIUHh4z1pCRm1LX0tljV5e3QarFzF
lEI0yuD0NsfS3n4BPXe3hO4LG9HyM6v6Ds3U5xQCHZvT30h7Zb/dyw91TtbHr+o1
g+qioMkulfzyJR1hqnt/AcBSw9F0xDCRTojK2Cw9bDPBWBx/7+2JPTpWk3fx9FRw
6h02dVBa/mhwtcE46jIzet9g+8fKES60dR/WbzCA/W5l1PSShj+CnAiT0sA4Gb5T
OrCVvbyWSZZCXboL/Rdsy2jvqIaXDqlq4kbjV7xoqJAfmXDjdW6rRre1Z3zRmVfe
WbetH0HWnV4o5v5W+rUWUgeKMDfEMM0o0DmV6S/f4anhu6w7XsaS1ZXnboZ1uq4Q
q0xDKVLz8d052dh+51K2Zf/MI3tUCvUy8r9rKB+9Eoljr58QiEUJfoqR3faonhXw
63Ip+OQs+IVx4wCH4W+TaB9hkx9fP5YHIcd/MWGqqLRx7GBaj5muTcf4D7lCgTjK
Ipj8grosCQH6ITbvfMfURSqTDvGNcj39FUy5jb7i1FqIKVXZv1NyescJYhIuvuH4
AZi8gw4HslcF1gSSwzVy2GkfUj1WetdaTgDIh+x1ABvGy0NT/ctHEzf/IPg6u7kB
u69+2P10DVQO65TtGs96Wbh3fsIf9sufDuVHBmegUUZn0LZd5bvex3pga+WkikyL
jnfqOhCyb8uAwyBp2aSsUo/9BQunPKDH/WxD4VPsXDKYXMeWJPD9nO1v4l3rr2cK
GuPcR793WNxXwfbhpmRKPxJqyi9r+8zjjsJgdkKVzelc9jvZc64gm2lB8La17CBz
BKjUflcWGG74zHdIR0CtBc7IvVmJv/YXTdbKOzyX2R1FhmVdp4Ib6uxSNcVoj32B
O3FMIPk4kwa2JOJ8Jid7kkjTkwZKei+d1V7utn7vCKAJTpjdN9nm5D5wKrr/8lwn
7emz1+KtjFl+wjv7lvd3PxocwlHzm3LDm30q/TaOr1owAxPy3ByuopWprzS49MxT
Tex36FIKMV9mNweqM/KPYxcOUe3fLSv/8/9E+Uuu6KbRFMVH2mYNQg283RYU9VO/
t5BEmzTul1t026VS4483QmKNAiIZ7CWpLg4pprxQvPeYb7NGXJJqhqAQ9WJ6aRs5
mYMYz2FzKkvZLBRn5w77qyFC7iT0MCVZmxxO3s3Oxr6PggvRjQRzxadgHTV/4S+V
ozHp0PRhSBPhgSJijgVYMHQTODsZj46m3oeNy5ocmFXLrhFM/MlVoDx6ECdPZVq0
n67GtKqO/6mNtYp3D96v9y6rRNoqyhXUF2CucFIU/ESiYeE9fhsamTDYd81OhhAL
CERzAd6H/509L5UjHUl1eAQ0FHOPFEEEp9qvfz991egRGmuQ/SLhkL/Nb2PsejA9
m4vsUD+nOaPcDb3+2cJAwfCPnvD/HK7Sg6A3d35NHeRyjYZ0ML3dEmdyyboFmzrc
rdTCX7SXNcvUOwgFI4FbAAdhei1Ze5okTVgssoMgfFp0khJXS+eIU/sQMcvyne9z
36a5wd/raRoCx0VG6wLHM5Cmxo81KbQtPFfKVX5+e9DMNxXTsu+Jg8QqylRs7HpQ
cmNvQgnUDzk0iAfmbrmUkgmERZze4JIFs/PoAsJaCxbgfdp9M7j6cPaj+3CYKPuB
zrZ/lQ3BerEaZ24M8quNqZD4O0bM0iNyQKGs+Nrza1aJivzTvDQGsHYqygzzCUzI
a6koGomlMDnjZen2EJLdDjlRTzC5lX0sk1T3H42MVmHw5ZuOUAOuqutftT/2jvJ7
xrmr7DVA0sPAp/hYiTyJlJBK2uh06r6V/dyXnn4M2PseHXTZbfCyMRGs2sqLhA8a
F5Eb80Is3n2xpk1ETTZSfrnpaR8UmXJngTpwign1+wll70RTChyi6qSTTExZCqxN
31fIO2Ijbs526Vp7eET/cIej+zikwJWyw1oX1PFzaJdVyucOOtwRj0/58wVcaG9I
kvu5wpoIXFv3xL5/mNekOVhm5NpFM3A/F7JWjRKRvq0yUe17h19LnX5AN+zVCMk8
4hVAx+kqHaUNhLMSs4+foZceIGcFCAJheLdlt6LSxXtwBJ/1nwpnD0+K3ZPYdOJ+
wBwfEFFu2J8HYona8xxIqzhASiYtyOdvQ0QRfgeZg8i2nNJ28gU/C6yzJNEltFKI
giHK1OTHfJJkr0M1rFcMWxu3FI1B3BcQnR4KTvSE8nX0Drs4fzUgGcY0DkihbHEn
g2meXYAtOzYtjxx5r8e3iRBq5NFc4mbDOw+kpnOFLWMVWMdVTLaoMWrcU/c8wO1w
dSmKS54T0Z94MQ6Myw8FW9T6Yp37KhumdXgho/IzW0HWAWFJc2amc+ygm9mdxM2B
svPO3eajxHhN6odouLOIs/e04etiB13A5h3MFG0tIVu8Fs6lhmYJzFjyeXqkq53+
XxRaS9Bd8jINlcevZK9VogCKesJYkmQFd8GxLOjD27U/LYXVyNgXG8Wn4oJ/pwjL
RDEjiytp3qeJ77hTMzb823MOlmqXdsBx6r0vdZEyWldcM0AG/ou2VAgZAxY0/vR8
gPIap3cb9naRWSa1Ez250mGgUoep93ygYnRz4bujjxHAZYJNLNphtuT4sW/DVs3m
fukmA3AHvTczSoW092bC/npn7MuoYFReunc0/YlC7XZ1+XvgpU2cANGu/cQOdGxX
s8RVOpRxVvRfXJIJrMvhDVg3NUfi+BmVxPJ+q7+cjVI2IrUs0oTdcS9lEIMptJMb
B3H+F0VXwX2Bnodb9BkmKVHqYDbGJuJnoyUgIzrm4KK3tfe94QdI1fAAKhMrCeHN
KFwVaW8dQIVC/P4ump3qxYNLNHvCnjNKiyZ7LaoerAEVQxa//D2VK+KBe2vR7g9u
ZQINSvKAEiI4mB4qtJ4K3Qp0ogcfBpZZ8b4CSwv7/XnCkYKi0pOXN8+6aJk+y5aS
6HHXiVMc2gSot4+SZHiKrYuPLYPlz60MkdjePiVYT/rHc9QCRSv4uVbu3ZTuzrz9
mzwcGxFYA1cKiNyCucYT1Tgh3NW75D/KSa7aZbZtpg+gEZNXSuzAtbd+/AZBUw1v
wLMyVfUFpCgw+RoY2kVxShA13ECTfHMgJhzhSRndxZNWGia8ShQy/MYljDpr4LcN
N7oY7KHVzv/OUU3cXVQdr2P8FzJEXrP88gl+bxslxuMG2Vq/dznS5f70GuHQf5jb
wXkAR6g9S71MheUdWGr6KbmDvcLd6ljamXecTP2f5Q75+g8Xj5wKATjr1l4UCmM7
9v1xBtlmVj4BW3jvQdF0HekUntoFFryf2z/tnAtYN5y6+KLr8ksVxPk2aiV6rNuK
2wqAHaN7hXUGnI3sTaiSdzYFitWDzqOQBFsGM5aX3RefdrFWsNEdweElT/R7i1iQ
yGcxUYNauBghBBwo2qlTn0kn0gPvCZFHgws+P4hWih45Kf5hyJTH4FyiazMKxSeT
8V6E86kqyoCDUvcYDRSzQ6IGJpO52Syah1b8fIDQG393XyflgrTOmHEV/TybAvGD
5G05Sa3bFfj7ApJJF/DFp2G/f3f0OKUvoEoV3HJcYbmUIMb/8cB9clZTaV40JzRv
g2WBsFnQLHyXME749wSy0UN0+NbTZ7vwvLqY7+7KhOa234nFlJTelZNa1PX0m9PH
TM/1/djpCQMT3VkM5lVkbOQC5/3UGq1F7LM5XJCcBm36/WC1re65vn+i1G+65dCk
KyArH1R1EiBJhNLPML8Gwa3vu1V+F0rfLrAxR3+3LGR8MtI0UFmGBsvCtwlcqpVW
OnfoUUH7BOWFSUNobNdmygZn71xKQXXpC/z0+FswXphLFEvyM8OkPoLAPHABXVHa
S+wc55EOA4NBb4ma62mRRdhZkXabBlhdHpDHV62S7hbTth6x2jkD/uZ/iTt2O31t
M/ylTRetJnmEB+NhjEc9a6Nsb2rJSmDQ7EFdK6WoUaKMRSvpKGGu/82jrRox/nGr
3p9u2/md7muAbmw1htDHF+YtbSC060dCCa9rgWQ7aw2wQFN7Gy/03VT65TzSqEDB
mI2tW/JKZWq6OKt3HerXXCkf1LBHfA5GZBdd618zpkqsXwAfynZlrFNzJCtw7aQw
WUPysKk021jZHBXJDW0AMMMjpnFjeUyPSX5x8yg8MoCCg2GrhZpMCl8DfvJl9NCz
tXV8mkDywKnmeYegGUquNDO7og4W6jwh++55h7s4+W39aprFL3vSIhcZOanKIaYL
eDlcPUXwlZQOI7p7HCyv6yQ6XzlidZdbAcTFpyHWQ9F2eCfXdR0zoE4WnSLszxsf
4uFAugnE9KPaFyHvBcVyYdFtl0TFsAS5iDrkYek03ZlQmNjp7guw0l0+1SCTe3i0
Oxmwy3AKAGwPlwofKihcOyNZnvGo66Hct9MAw9Q/DDaoZ9wP2tqQYmzG0lZwz7nr
cYJr+eWvdIvDm3LMTgwsLp929zs2q8cd1vOe3T05VSIjU8J8x/IQmo/Za8AzQedK
OJG8cbU+NzhPDkFcxEzUPc6dzXB3H9Wda5MIzxSm0NyXEwr+iegtMhC+nxIbgGS2
B2hoFU6XjDh0YARgc5Palnx8MMYrJsbXGD400dnVeoX3mgViEhzKQsf/Yq4+fyob
0ZAHig8nzMIvNYvqdlf026gxUTtIM0X3z7Ck879LK0c1mRGD/8qOx/8pQ7Gwjep5
LW54hDctsUWfscX9ZpFMegKQJp1sswc5mC2m48/pI6AUoFSGbYU7xpXMolNyFV3H
60zu2T1IZGAVM7OVNVhXFzxdDCrETcIfVWmcV/OjTo1j7+URbrgY74RfAW4uBEL3
wlXslrKAF66UYjVaUj1gh2QMLNKh0ujshvPEowMGJqrqXdki4Kspr3falyi3bFys
HjpW9v9xklZ8MhczY/bZZ/MIVrmsoeJAL70pLnl3eg+DfLefjzZzGq5X3Z2OSTZL
4Jj9DFOnRm53PxRduHs95kwe5b/gnwTwDM8z8Qf3+RcsiHqL4aALeRO2OtyMl+/n
a92omyD/hQFBzBMFROc4ksS7VjqcdYP94ADQN5MyZkybQTCNm3+eYuEBm+V609Us
2K9mxYcGfsCI3iiS0R1rivJz2V2jKSFKFHh0ZwVxx/OO2G4RMduwMwP6Lnnysdoo
JBbj7UNR8N98EAWvCTJi4TGvKvAs6aeWpwXHrQG35bGRIMa7iCyTGM392LTOagVt
YC+MwYcyuvQUmBN85CnKJRqTWsEe2613YBt4XqmVDAbN9wYeRo5F3GxEMfM4+6gQ
ZQC/i1U7vp4ZBDJYym+3Y+8aYMQKglHXoKwZazONCNJeJtzGrYyEcR2btRR4Suo7
1FTjD02RKi70yuWPdVWWLQ/b0Ec3AviExiR6HaV/nPpYFLiRjXJTZxrKg231MUrB
FdP1tWD3Nx9olG5Sz19A3v03oRxLFbYAxkq9R6H5FJng+/WYuC3IYA9PMhXCXc42
JibZ6SWIHfeFhow94jGX+yymE7YK478ylrDuF5EWFgPxVz2lf3KtDDskwkulDWZW
bWHHrJIPegQCVkBm6qcYcRLEYJf39Yf9VieiOG/TsdydEqrN3Xbna4wJcaUjjptJ
FqRjjicvUj1HJaIGfGPTT3NE4N2AE6UMHpWhO71WzCSFQ3Ql0jFOfkxCQnD/8lRe
2X2kUYjsYUG3kQiy0cP3fSf0BGKwlPiSvViu6jY8c3FQfVlwJ4vYBHDYrHwxNE9O
WhiGUQPMX3DxuQukgP6PHek0ZENOlHCHx7yHjBfiuh1sA7gUvWJp4Qn2Iga4xb7a
EZH8jDQIyjhGw3o98zbHaMWcBLSNnKXdsvpmFzOM0NunYO/6delLCW0fZs67dQ0p
f9Ix5ZyTq+N5spQyhaZEko8VqDCrJll9AFzDuncoXiRew9eGqGCcVHVKZw9kA/2+
LOcTZJdCJjCUAru6N/k8UAy2WcWJvB7lKSY+6klLxfcZmKb/5lFWl3AnkFlveLVN
RXWcMD+kAtd3onDQOeoZ0d1OXt9EddRQVh+obzXcOOqTqfNiLxBEqx46QnYfK6EW
CYHjz+nEe+HnE/P59tnOQKmhYcHmgOYRErqxg5ff+g8VcAc9cy2canpX16OvQ+TV
Lf1MBcCi8a3yV2KzQZYX+r5f8whCqrLt2/cb12apA97F+HkjxBhnzPHcyBjpIUgu
oGdLEi6BMKx//UGUIyWal4l65QrlWoQtojhk6nZ0k7y5tDCq+jevPXJvCbpsMENR
sQQ26B/gqOwqY26ik/hha97O8kM/SrjzkI6ZJfR5ZGAKgjYQLpDAHkPpDwQFYM4a
csk44oL5uxIIAJ5+5TsXRVxzhgIe8eyqw9vs3L/27bEz4aYdBRuX3NyNGaHCv+w/
zyGwIhu+T+KYj2D6FXcOxpDV7q5uI90YuoFw3Xb1cm/rmlHxuS1Er8zOu1TsM2BM
z/l50qc4HBLqdWSIFKtH9qwXVbp3hRvalAQvqqlhpt9Gih+d2LO3JFnWMXrRUVSB
hp0XPKPDukLHDWicjOPAyQl0Ut+Bx8UFsIn3McuF/NFfuRE1OxpcD6WDzi70bkXY
XDvAVwTEN6CCs2RU1L69IY3xmnaq26+lkNtx/bf5yegfrQGl1IZYNwJkcQ1/fi/O
QWUZxCwDaZK2eiQkMMMWEn24P/okwD5LmDvOkkHQClEAidHbE5qDUb0qb2XIfUwI
UXUytzSoXgckro/NN3Qc5qryMJVAn8rN/xEm3gPwEH9pAEYu+q4QRfF1zRzzwKDl
cqksovozHlgyqS4ElNhEnBqYgMvglu3a3bZEfMvJNBZ1+jWJuMJxnmaeiMMCniKZ
c43uIITyrLzFSztjsFyzmtYnhytCBQvxEniF97vZAynZglJY1AJMKVw1z8rOBtv5
oP+4PfBquehnPe6Zw+wLoIvAqjZDeyo3D1Y7uKWJVqPEXz5bx1HLlIROEfUhjeCy
6do9ZHhDZmqShFpZ59PjMr7QIOEGKwoOS6M7qVKfcX565oyCXjk5I83wcwjx5MlS
t1hpzVpSH5hsfNjw2/jA9VZyg+8tmfIjYO7hf3JWl5niwxq8dD9ErAN/v2eScCCa
VNUrjsCUE4wmj/9QAI975EXj3BqkusHWdMOmFAFiOox+3lihSCBOaMSAz31kBbMo
4Z31g21iOlSEdXdyPSxRUStOqd+fru0QCwANsxMmwmdnRZPdgM0ObTTnLauOpJXb
GmlR9L2YEfFlLiKro353rJHNV4EbGN7HdbkTbOyS7/wxWxvZPIeXnMX28xXc2WMN
ag92AUfb2BmdDUq3SZrVNZDKdqtUChF/Hw5a7xjXo0tuwFVu8zLYECm44nJdw0EC
ZFhwQneOCDomHtlr7d8c6n5DyLcGEh6z7d5Wc9R2bbexT3W1l3il4a6t1aAp4V3Y
86K7b44NDqydHTSAL3C0xjDMxlX4aebv+2g7Q7KPD0mhx6+cBQsQevgpiTJAECo1
6/bsVVgy/4zAZlGldLvs11FB0c9CimLa3ypfCzOSo64I1CW2AEfOyegBMsomyKKo
L8zbjubwk9YthY0q8Scihd212meLXkz5DOEDc9P5msn370DeTkIvEgaQ3o179Fkq
CwEMs5WmGsrW8PZCsNKVE/Y4zau4hGbi+uoKNiWWKSlmH8p2aKGnjNN3DA4+LrBM
8EEWFfhtd+3bOsNaVFZzlVCngwd0jKwid3AukWZkVZLbemfS6P1dByHyHWQ42Rz5
mPiZmgIfRvixJXS6xffHcFG8edMbAVHPJ8ByL07YCe8tbmAg3ASgAZc3H/4lRnLc
IWQJb3GawKP0uxCHz5o1Itzz1Iy6VdPb2ryAzZcoeool0SuX5I+HcrVsmcgM4K0W
gRaobfr7vZF4RHbyCZPEdvn5dd+Y28vw8HRJgAZzrz56Q6CpZMvp64rRBWtOS1Qv
ZIu9T+Uo5VdIW0T+jK1IcqU7bARpi5tAoODNJ0Z3h51BmaC8l2cOMAliK/aVa6qr
4WUp4zbFPVbyX1qWFIMPmyLjq/p4bUOuv9lkgGqP5WkRpfv2EkpXsSRArI9YhjuA
Tg+5L20UaS2Sed+2BMSSJvjEPs9HuD+khdQflx+oW2fhBYmohSBoQ+kUvJquplLD
4P2Cmoa1rq5rgIWoObVvbu7J16LgrCXmnzrzacGXehM3C6wkX2rrqjsZT5o5Msc4
/abWU0j7Pi2ps/S3cIsZwf340pcS0gYw/qzfu5d4VAQSGzkXwVawBMc8FAYzJoQH
XRTPkXP7Jt1k/Q3Bcaoa/yFQRcdZGrCV81/QA4lhZXyACJJItqnoL+y8Jop6dtGw
lUkt7/Y1yaUQcY1K09Y2YxxDFmjAoMGu5pKdQxdBcLfN35DKhWfyB8QU9D2uyaaf
qrpAj3CSBt0ObtV7peIQRxRrdxyxvWTM7VJitcJzNzDGHeDm8xgHfBLdLBSmv/34
Pk5ZJ3vRJNLljyOyJJb4OWpSQYEqDSVp2n0yR2cZ42Yxx4p2GWMLJTuM3s6RYxfs
1DT/jgcyu+OFWn/5TIXurUOZus2ai2eOrhfSZoPzA0lJkkajOqlmiU/z+EanOe7h
fuoDAEUcM+Gh4WyBc55bx3iAN2CVDMzYnwM+VB4YvlpOOfBmYp2tp6Fr5k+b981X
Y2JRN2TXhA+HW49hZJAATQ8gcWCbznGgthsiYN3r+ICl2Sz0vEkYkcpiPyqAI7Dt
aHiJr2L6vwVSpgyFBj+gi8vOXHx6hY9mExq4I9oFydrPvZSWxFGuwJ6/Eye2JFVT
Qh3ZYIV9SZXCwfvAGhLdoUXI4u8zoJERM1bnBUVbPEN2nE8JM/6Y65O/2knIXJj8
6mDaTyJuDyAN9dLrxe+dlVFNB66cKwnYh9NtFPxOjlXpOGFkpHVghi/GGDDg9rGT
wxOpElTqMcW0YugO4BichyvRxQ2eTQZWCh7xD68fPtlNL80840AY3ush5GJlD5nz
Zoi4XW9dDTNfsQfsZ/2IS7bWbwI+fwgviWqpA9d+zn+wZfdhlo7ZHwGlvdDh6Wa7
s5goSDpzVhJrBIGr3CYTuOTCs0na6mCw5YGOdxNC4d7NeJ0CwYkbgf4WxQg40+kM
ke9OSXi96uz5ISpUEC4taxfskY9mrC9EcD6+eHldzJQBP7z47r4pyYC5cvjKclCF
YkGOTaWPKGYCl59n3BeIF0+ae4ZrZr4bI7IspaxCJI7PilA0f2DUpj6NFNLZiFpi
r4znpnJmCSM3RQI8E1rzzjYAOrvNy/QeMGnvPkn2e2FQM9OzSawwUAyJnJWhupLy
anu5kRgd66uTOPDojGy5fSXMfzrNqM8uqZJEAPDZwcBAEAPIZK+Vy2ZtzZomPILn
zZ6jMvLb+4bLiwZJFGdUq1UzsL1BrVVsohIsbGh8GLwytHZwcgfrSHcytLm3Xptd
obfPaTIR/mI2YXOaG8oZ3TzYH9UPQSbfGIfytlwooyU3VTS51CO765uxNlSPKFzC
/AGazjPThcJMGPyfMTQDjRTXumYKndaSFkiHN3N6Ke0RrAyNDUHFyXGYqgdwn+JS
34wJr/np3q0o3rGFKSR3xsKkQhNEI1O+momKkg8WiYqsT1jubovq9SCETzBSn62J
3oY5LvaMfkQ3PwT4LGSvR5B5XY4UqescQPohAoP9eQuISi0epHk/VwFIR4ynZAlh
Cwo7yCq5IiHCLxMkjro1PKKDk4+Yx0pqcEFT8WW5EI1vFNYi5CalEU8k1IHvxD40
9joYjQ3tv5+t5LDoxS6VvSeSkDsEJlsdqOkx90Z1ceQ0GnENh8mhAIegamEyHhm5
qmcKrwoD6KT9YTarCM/TfmrGQJN9mbyDs8rpanv488+ebbfsw3KXFpqfv3/WukRG
jNBdejYf7PR/jDLuqOPxMTtN0EpQ+lmMxT7qfM1c7wObGQvhVwLS/F+8944yddXd
31GFRtDMJ9sbHOV7s1fpj/lug8ZHvINitFnBTKwqpnhXNqFZcfVufge+KO3OjNed
6/4ZguRNDwRnhhSXx6wUdTGT5kQ6Gp1a8XFfz6Du7Na7RrLkdeOslSu8YFt+KK62
0duaJFseqsu1fepCviJVue7TTgUcH/6wL18YBdJ3CLgavRdk5HjlSTSlPljSaUo6
vY+Qd7uYalC37HCY5wYW9UpruW2Fvy6AaUS2c6GKs7hZWAt5mXUMHxGxE48AiyZu
9UGD38yFJ89/q8TP+QLq5h1zzv9Dw6IE2bMOIXCleGwoKE4iBCmblqqR7WKFTr85
kJ7OJEkKgb4hcBSQECM35t40kZ9ta69hkpCiiMarSQsBUxg6K8cnyCZFRntvKhwB
m3/f4CHcPb7g0w2O1w7UCU8oeMnX7nIy3MoKAjH6z/i+coEvTotCPHj5+eSIuG0g
08mSTXiSSDICQ7tZNngotjSVk+2Etydyi9P3p8E/e8IsRMN23I7B+gU2ljG7G9iq
6RuNR7DXWLRVKzNzuBkMcSLManWO8gz34SOb96X6D9QJgkq5MEdvMXndl7hdHXtE
pqjEhrGgO2w5cxAYIOFvEioXhSMkyoOHuS8BHDBiYA50NVtCO+wWEOwqGM9ofU/i
AK7nak4X8ksiKQzn0g/3RBkhgEg2jBJORh+kAT4ayu7L9/2NZ71PRhBN7u2URoJD
M7LWMe8+iBMX8KRE+E0ikJcR5kvgpt8bhRaPcoGcWrRzRrwoFv0SsR51NeXb7Aq1
QgfmJukhrfT195Xennp/n627AvPicBwuuvx/a/AFwZhkpJNpb/QVeciUtniITVe9
H3GhX/lXHqDswrmgM7hG8rouAUB7sk/5usNUMcarWj0aZDh74oKvnqo00Z2zHvJz
S4fyiAETHf3AdtHU11O1bBfH2Qbivbj+rmtJL1Iij5eQTGuR0A+raJ44IiMudXwl
MbfvNHfXLxuMo/O15C/YuDgjsi+NzHseoU/MlmQ1aM0apid+PxgSmCuLeFUmIVoX
LsDK5Jd+DfP4kPujSO9M3+86Crr4iv2XsIGUIJYPCaecLkY9wCNqsajWbjkMxrIk
p7psDrIFZZHturUG0ja38fW6Ko+wZhkjDBjziy8hrfzJK+ZixBVqFsYUf67YajvP
HZEF/vWAocP1OdqK/21kM2oGbe+0egkZRf11HGMS19/acIxO+LHaUnuD+KYzCUqM
4C/B4+kDNaa8/5g2k15cpgdZ/TIm7te0blGd5Vcgt8r91qOdjXtob4xrVGc40PMD
4d+Dtz9Cl8Ga2RB+YM8v4eH8Fi3DoGbBoDmMJ5SE9PptC5EREeaXukm6oKVubWYS
PPwfBQ3+6ysKUHGic8H5jZW1ZhHNR+fAZrZFsSnVeTVawADPldxpXAvX/wJvIdi7
KHJifn9R88MmdjryiJ0pC+LTfEWlP/JHfmzX7q4kBj2qj5kBmvqf9Ddpnl1AKeRO
HeMrRPJ62luNufYK5GyPRP8NsCvJ43IG36d6wTXyRm8n4vYNlraIc2sKy3OsHd0f
FVnTluaPp/ie4MVoOIHUEmaJLkTl1q+uFGPnn/79QxD09B3HnsGmppJ3YOBw6uCz
5epHHj9QyFWxAXQlfRxbJjpP77G13GCsVJK/YMfY55X3Y70D9lzTgwS+gr2MAMwS
WZ4X6IKRLMdpLlUy0spqZBNNmFBqXGo2+RY4zlQNATQYoGuP9D8Fv0x8wvYQJ9dB
9RPu9NxfOuSe2sXSfi/rH//Z96ZNEafPrzOgaYR4f5q7sXPDt1vOl9NM9BYJghjE
ZbaDvl8DhOoY8hi61PcU2hn4la4hgxICjvFj7BNqkQ/m7859Asu2LzVLt58YCJyx
utR7JiUvVHdbqXy2XrZ8yYoQOx3bMw2/7nk2jCmaujlHESxDtHBzFOYR6hQbvEJ/
PiLMzAkC3dfnYMuBvxI8GL+fhfSC9FKFNtAUPUImrye27xOKcLqdyYlOMUTD440L
6e0XIF/l0iM2goXLp/B/rO1M/lb7YO/oWUOt7BJHkDm6UBi96CjCK95AT4l4Jt50
TiMxxKyAy8YCwbgfEFXJ4R3+43zhH1/sRoy5L+arx2wivWs/VMkgCfQ/IYImhbdB
8SBlvsI2hpbInguni3zwb4MOyf3VWmWMqQ1Httx9VjGn4A5T8uaZoMGmKtjiC832
ElUnegn3dTUu3bftx4R6k2SDYX/Do0fUygAQyZOlLQ3NrmOZaEWZVU9vDFwIcDIw
NeNaLV2zYkfbjkDO79UoYpzHWEgfmUVl7Vw3GbsazMEU3wgAX5kKFJwiOAfV+tt/
NTfOmbFg3glGYLBiXSmwuemUotp6BZdmjgiQE+SwLxNxee0+p3s8rrYdSLbFI/2H
2JB7LDyQcJKx/LHOn4dWYt0YIkhZfD5jvvZofm1+Na/XjZBs/H2hBz9MzJrg5vHN
VfP7glA3OxMeJRwQKlFqGHRednRMM0wngD+GcsESiFo80zKMY0rb5zOR5C0G4aC4
b8FMlTiOT37fsVRx4Z6ikz3sxmQxkGXOYbPTOvtQNtGzSTI8mBbAk34u/4ZoPVBl
GgEr9NlD/imy3MufdWgY/bhya40y7OlfGfTGISk7an0mDK3k5vJ1YMLocMrjxJlC
jiBdZwhBZnTpxtJSbqQ3t7hw/uPMyuSVuG+iWlxxREw2nS2hfiJoigqD3nb0hmlE
rzjSUWPqgrTq4ZbRPDYtfJGd4DmlWPte0Io2PuUwXvUYEPYXEBWWzwhE5JRK6FDG
HLxO9rrAzJcSiW/bUnpBNu97nSUons4fAFHvdQJfwJIcPd0KuRGKf8BpTqPgDz1g
F8N6px71Szg0d/2O18PwUDR2pwUk8yfZRwphOkOH+7EmvJIogp7+O7AVLV4UeErX
In4gf4Nk8cfxY0dK7Qw+Twvot7mXVFMwP41qf9GroFCLTg7xdZ0w7ky1OfyZwINU
nt/mULzFKiJs95S/bWB6PkujD14UxxAY2LJtP/gB83tLe6+UpmsJFGUnSsn/Zhot
N+OlbDp5+66iS8yOqibtkVTcX5C7/msxltrcwJ1DopzCGuToOd1PnkPXc3AuHzDJ
mqQyYGs4KcN45/Cw4tjZTJjKw9vcE7Lqz2RngTukmpoEZvDRpPcaDf59ovNKK9qq
X6vXNxQGGTNyodTB+L4RmUIB3W9vUGBwpM5fOh+YiO3BYKNjA3O3wj0dzp1LMkO3
Hqa8bNng/iN3curzeeYa+u1YXYs841z5AnAUvv1aRLMM6tEWUlKc98XiTApjRYNa
CyAkzvHgx6fvgAAbTrgkc1EoBr72ApJstJTvnln1TybOSyaL+vLx/Gl+3iSblTmv
Ty+Bnm0eDGcEVAY3uwFbIjLsFar/fs67iEXhV9Tv3QoYtsLJmAS+HfFnB3V9CC7v
i0dQdikSEjyd/V35Hi9VWz/AHt55d2bhOOvOLflcbju8dDDDbCSaocX8wkZfiSqo
mqJZnkBMA61GONlaURsgqOEMnlmV3zLzGrJ3mrT9eR9piyJw6MiFw9gR3IVCZaY7
rNA+1p0GVsaiU9VTvgkGp3/5Vj/Vfuc277UzoUwLLjWJ/IY0fD27PEfvM6HAgfhW
rKfOwp7ei4KErp5JGXuTIvMinvCpnTp+W9I7PcFiel0hJyrs/dp7DMwcFazJTy0l
HtFVPeKFfAA8tmK1/RqvedNtMHSGFlMg3WVD1XYYsK/Zs/0OhX2wziICBCQoScdA
uxwq8e4ZjOxVo44WwTD0Nk42877Kxt2URebf6NwWj0f4p1BQSGOzSeLhkGinFR9r
z5BcMD6DcQd3BzEVQgw2dhWKxsI7VRm6wYIqJH3L30hFtcyyZCMSrNXOU6wdJIO0
I5oXx1UB769UKvNe09iFQ7+rIcLNWXiI3u8Aick+zQ60A+DAe8UZUA7pc1De1S6t
f+Z/IQNii68N7Oxi+R48s0wq27ARvY4x7sHdxgEAt07oyVqO4sQk1TjLJj8UyLED
vweyrhfKcZBeZoYuC1tVNJgIHehdDIso0Z0iPrFPRmc/Ksq/DYrsTI4mChBBf0+U
0QjUn6iaWYRr7ScsW99291Tna7cNkIl1Z37oayLBedX54KuGRE950yhRNailA6kx
ya8G0gzmb+SzBUJtPaH0pXE8ilExiHbavNoOAP3Vppt8gA/fli17gYgg87lpg07R
onR5kDQRFsfndsnNlLNc42bIzRZks+T5zI23wpd74LBfrdJdq40vD8/UJJI8/JU3
Q+HhUd5/C0w9jiWa+Dpy8/YDXAfe33z98wR+J31VUvJbcio+xrnwV/HbkgMAoFqN
Dq3L1MgGi6JoPqShSxFpPmFWanJgoVGVCcc7n9IowVVmD3Bebo/tldLyPejZ4mDZ
jA5pt+TluSFoaNyHexs7O76M4A5AaVf8dkM/1M4Ta5kwyoZSJ6vZ3JWF9Dr2uvcU
pPFyExZfnbAjGrkzS/sLXAgboZjB9E9YX/gNQwH8mZUfTbrcoCsWv5aTadLsVicX
82rufzhlfcHOoRMg1qITzkevMtZSyVfscMI3w2U7GpFKImiYzSfs1vulq3l+8iro
XefIpPWjG15zcD1c9P+kbZLta8iZXypODbrgTQMFIEHpyWZZcND4L7Zx5ZvDL/IO
+brr4BIN/YoI7XAIvnMilIzDbVP6RFJNtRjg+azjhMD1xfR1JCf41UNuRjVxrdRe
C+RxQenx20WTTw90nDnJqj+8NUEeOg3tFcpfRL02EnvvrwcmMzsx0IYEG6WjQQQ+
R6MWA2JRf36uAcXnmPnpROTOG/stxxiH0AXWYReb0L7qE2pb0PKI+BuRKAIUZQFB
E9IvTLC4sNn9DtszMq38U99rBG0TYYvGs95hJYJxHeSxENeo1SQ4b6VbWs1rDPTz
psEKhxnfOIKYOtlJhKmvFFUXavZVHRsuVPog2n6Ilep+EBw5i3cPr/OYwtNuCyzK
f2mUpgwEpEca5kc8ggO0d94id7AKVotfzZukHmb1O0Cmj9ivzVROEtPYiwzMs5bc
sJuCLvRBiwP2WSa6Dz/XnpfBjCusNYUErjsP8k1ABKRG0wWle3V1JqwxEcY7U+n1
RzNwqvfORG2dym/UmhtU3TV2dwzszQZAj+GQKGmxE0mq4CQECP5PX6MFQZOc2ewy
se+c8egV8lxzb7oZr9/xHHbd/mAzuGkWARWd7bAZa/aCGzjzlFd5Zztf9KkXcaq7
eI2M/6PE/F/e2hUg/Qwhwuu+RnSG38stAUSY/JF51VS0NqPufyhoBveLJ4CtZ4Hl
u1X529k2yVGFtn3x5oYpSCUSs04/RGoCBRtX/HwrepO7m23WOr5j15IHV1Otndls
JtqcGPg7i44d2LnG7V/I88zXG0lLCGmyZf4Gbf4ejKQXm+HR5ny22+F8QXiZjBJE
ToEdpMrKJcVOs0l/QYUvVM2ISvIIH8n8HI9Az/pjk08QU8BXp+GxB3VeZTfZvdPp
wFkLuEm/GxAwS0vCEmSXUXCSchoW/ziG1tapV3i/sPaT1Na1E01rNsCNguh8wx6H
+tNkzcJ0vOBdBmi1ACPv7GbUC+stVMR3yYyaEtLihg4v/Ovu3Lh4J8vYpzMixUv/
lacpdjrZqj02kSNnKAdbzwltcebVVw/yGCicb5wQuElX0AfS0zKTO5RFlgIUeMfH
/RAdpX+CSBj8maorUw9ugQFQDFV3YeihG9ez+RcNzt0xGCT43mRLK0c3PHBHY+nY
CM4BXwl+hyFYQ9JCdo+br4mnFtnT5f3HUGUOZh4Dz38s0uVbFGnmF/wNQogyArnQ
M+k1tu0Wegny6ACXAcW/y5SkPM5A56UcUtFppAaVWTtb2q5ffNAvlAH/mB4l4mlu
ClTiNZNLqO1JuXLguY1tEY27ypvQ9JnhNlj/8YCFeSsBJpvtNFddBJxIy4KeY5Yp
QXN4xkwnjnakjAaApTm6P52xGqnGtrJVkn2EQGHvHeNQTrWnaKsyrvKH0ZcAGTH8
rLAs80QHwCqmC7Dij1UhP+Ib6G74xHnbpFkzD2ulzQNcHTmjnMYFdz5jvb17Fp4W
mGy8QAennvG5linB+KlNt2A8+IpVTOdxU1D8+E92G0bygheSb5NFpSY1n/LUv+WX
vehXkGdbnRz1wqagZc7BlxYpQMFvOplOQP2Izl90DNfCxk4FTnvz4K5yO4gyUpSa
08M8V/iLdiqrBtZy50ZEAGtJWJJ4jHBr51gs5SAibd5EIDAq2MAMZxR3nTrCMo8q
RP2SOAjsJqiI1kTRlIRUzQGD9DSOZ+AOysDs6Pw1TSy4c8PpvHtiVu5CjU/gw0K5
T6GMU4kq0wQ6Ey4j+CWu1jkLfMis2h6zex/wr1oSOz+XtgglBzN2Zd6m8h1Rqoz3
7HWGXKKdD7pEBiaAkeKBKGds/swtZMu+RJjjM9EZnkZ6aHMEFRHe7V749PY3Uj1D
dGq2nx1EIQHc8F4v2USnFc0RC1XUKYbptgev1eywEqKz4ULw+/baZ9ekNcQ6KLoa
2kz7B64h27Xj5SOoOok+hMuosGgCALHXEugGRr8/zkCcHsMXUNTXHH3ZGj9aXtzT
3BKqca7oJMZKzrPI9DLd7Hx6NHBPosYL5gciAgbR718PjtlkcHBNx6CIkVQa1HvZ
METfKeZRhLk14TZLUbGAYHiy1Xdh1IbQsVM5QBumS/ELgu1tyztSbSLV9aKQrhcp
igZsvFCAI63uZbFqKiFkmhcdWLg2MVQB18d6VMNvAwQJGr8fHXviPWpq/W2VWJBd
x1/9itS5x0AKD6wOgbFrywzHZo+PzDw0n3m1NcSZGm+GLkeES8CmWet+FrTs9KBt
URc85Ox6N1g6WgM6vLRlsOJy5+tU2jnSHNpz6opGwRg7InZS1pJrrSirTlFp4DIB
zZr75CCEvJrOMfmzcb7hZsmctBwWr/RmM6M8dQ9g3RH3fAM44te8HqemRAHDPo+d
RvOHlHMXnstSzpOCppHuufiovv9liGp6KTuRztHCMal5LvFn0neGM7xRct/VuO48
ytZgkWCFRmgFq633uRb+RPnMZB5VXmnpyMTCOy5jVVz3aFVI+i17IZpC132orI76
6VjWT7jrqSV2dtlvs+kylaSeX9DvqoCF82tqbNya3H2w59Orm38+0FqKemWQxiNp
pfdkJscl49en8Asju1B0aj/0H9YetwuQbXSnFCpOoYMMJXF8K3QVzs4HHuLGygCW
aOlgcjEF3G1D5CYrj5CT658a8IXBYUxA8Cuqod/tF8KCYHO6FssKDndH+JTETdoc
VDQX9uXx4aivFW1vY20it06ZdYxlGiABtPfjckv4pZyeZA8YWoahRdDa25/GiB7l
tjkmSQu1BD1/YRYJjZdbyWNtDx9oWoGREH4uO0bgP/mvR1I8R3AtCCQ49Nm1+eSk
LhBJrQoJXigZWPGnhZ9Pz7kk2VTGVyUzJjUTBSAUwoWNUIhOUEONhGjIVVt1jJ/F
XFRuHvjCBtgMER4H4MqkyOA1BK3AoSr/liluK3qoaajRyy8J3IMfk/hsb4eO/Nr6
T4dfcvOQcWcHVYMWoj6lTcT6+5KQ0ugMnpjIKKSdQ9OZTa7LeOazThuhVUqUqPR3
LUNpuoZTycnT0X8FVUugRepN8D7PU0mE9N1PYOUVcX5hOv5fRU0+e/wvJ7b0wg6V
Brjpe+cjlkGuoIKNxg4+T/H/V1/1x6QmBSjQOpYSNfxAvyVh2lCnvqtMDwWcYiMB
BbfDCbRm6lUW6jQaf9zkFP6L/zABoBJo3a5Ds3YLUQi3vCCetgSUjn9P1UbIuJtH
eC/oiZQLiaVOWIB9WFcB64ds6uBYlxZHUhzXKCWDce26DezGTb3LexdoCSifo6b1
Jdq1CXxWp9POxP82Y20ESLY/qeIMUIOuO1IYioCGcP0PjEwauE1Ki+wqolYJE04g
VuqaI3lM0KV0cM7ZtsUU8zOGYRv663/djSsHb1/u9hJsJOicLKCL9qBqeC3htZLo
2CWzoyyqtOS9nyKHWEFycb6ZRYFMb5Hh6qHifsbzinm+1jofcj8UyolLTGarisGO
mwKBCyXHJIFLbCgebYvUWPUXA1F4EI/TT0wE2tJtmu6SRpl/OWMBcrFfar9PtI8G
cIWHVoLtu3cy2w8JnvFWOqOzckVZaJ+5HEA8ohhbaCC5e1fCpaaHCR2uYPRGV+s7
bpGg/0ujUZ+wzssYAGNNtZoAx+XUfAe96DDGZY6QE2bUIL2xSV2+lYb8Aez8OTjI
6gmboOBWBVxfoMI7g57fh/U8HuGSMeyvOqaN0EqGAu+01oqHkcKJ2zTCkIpumxfL
9bfKPfZXhJAKEd5weVk400hnb9gqyvYzfB0bIjIu+8TmhDv9nUFi66ehc5IPChWJ
8tltXpVEYxBiqroBfD9TsfSPoRXxMGi89ya6cxksAS/Dg2p5Ut5wxLnoIy0jJ1ti
mXyUZ5f+x5AioFxwkNrpdGrTN8eNUSTkFreGKmrmghUt9wgLW3czVt6y/y7mPVjH
GEYZ4BzdD3eoJQRFnI+cZ8RrWGdl6U7OxTZf6X0x1EkOKLLzFcnIKp/hQ2aPjgk3
wG2BZnu4rKVKUJRuVvxUvQ3A68p+YIvHTpPRPNG0kPmwP0TQdpIAEFF4bIoKRmDT
WEqNbHEYT1dmTwOf+oUvLJPUkzCMobQYGAYh59oGOWSrntAk/uBCicBXFwcb7rBX
eFC0/zhkBeB8I4Hnc5ZbMKtDnIzMB5rHuSFXEr9XYcyNZarnCMjhxbruWg9HFlxB
hycBp2ma/l8Zad9JD2ks/5bx10Riz/pCuBZ49l01G5OnwrlmxCEUklx4pF5+xAAn
vqsoAnUopUG17A59GEYfVTkeOXHfTFEbt/863BJdT61B0S0rfHuxJ2wWT5U4i8gV
e3ZGFnKVyKZ4Aybjd6BtT8CjO22haQw+lV4Zw/Med4RnJSaEA1/8MoP1yNifBLQF
Gbk3aEn3Irl3OHXNRHpIR1zfABnhY7M+LJIuMhxqmtAFafmvWr1X79CjHKKykrUg
+hB1ooTKazs9KkvbcS2t/0+smMehW6C8Lx7OGaq+SaGNbhglrbsM+4w0lkstr+6f
usigtS8hrHaertlocF6+Rw5vI2KT8FFhEKlMqpky9d8HikxYexD/XieVKGNlTTEM
VaHYToRt9RePpUB7ShOWmIEIbBfs9W1dgk17qnvsJ+CSIc5tvK0VXJY4WeasZRMA
2DOtuOD9w+Cwryeg7ad9thdwJGX//I0cY9iEoWoUkvyHQ4alzYE1VfTySxolHHUC
moO0kYT0jM6EbzgSPDZLA94/6NGv+gYE5KbDz0ucbs0jyfDTfHr7FcEsn/Sv+oZA
c1BqzrAVAjf9JCRx72Gg4VQUKYrMBWIuiEP9yzQya7kK23FBRN3O3BpTUKG8r0ty
rnNuX57cQTTWmfV2B8kGIcVAqWeukjxLoclDNfROzuo8gaWL+ddnYF7w5rrbW1iL
pM/eYb4me3ZerpTilccU0UJwGQXRlX2UQrftyQmSgOu2nUVoORL2tTcwf8NwG3iK
zGISWNWjEfauBViLj8rqm/900W9vVahosvEjrvNH5Das1upoT/U0/p2FgFBLbW2H
sODIAN/CzYkIFqm+268sYsVkCTCpCQ4wl5wTS2t+dT/dpxIYk3/bwLpTLGN7doP/
SyuTc+C3gkv/mK49aDTbjdlkpp9cO9qgU1DAnDf+jjJfCBnjYSoK9G/nSqlkLbe0
Zcl7E87mILA25WMDQZGvAyCInzkChxKOSseovk5js60M22pWyd0z36zoqfF0KEut
CQJ6YFwc4DXfci1UGaonW0Mt/L7FfsAqHoM+fWn39ctS1+74gsDkPezw+jp9NxZx
NTWTh6VmQP5cV8Ef08Sjjbu+Z9M/P/VxyDXAgJfpDVkfPW6YinhTcQxhutMxOFkn
0Pw075OX5GPqXTpoKua4o0YLf4CjSwxemmwUGwB4l3JWGSjwoLgWEj2RLMepnSjw
o6SV0c3HY+Dd98e1iUzDYZHhqPrA0rM77SsE2usHuI5xMBI07JSTYScQakPy8dJX
+8nN9Opdl6op+Ts/zlsKjtGGwBTdnPTJaxl6hM8VTbsJ7MSbk6igPJZMUerEvPzn
x30MWCl9GiONnSktL5nbQZLGOFFgoBOwh2TOH16TTn6cqjsLTMS3QDk4wZldfRYm
/rPM9aRRBqM8hYv3PsrKyLV74diBjGDfjOInHDG8gGgWKyM1s7NknixgeaTBVvTD
qORgXgY6N4fauGx6X3d3XzVEK0e/soZG/m0aP0XkvAaBOzflB0BxBNA58W1w03zj
SvUQI2wWGHNEnJFPoM/o8BcUdzo5suOcJcyDfLiE5D4yUncCCEu6nzvmhPClqQ5m
+SQ7ajLYybAqQ8lVJHCQrMmwi8UQ6Qjd9qtU7JjsCUptoQ6/cxrfUFbKlxlI6fz4
HMpIv6FXzL6M4piy43yhUbmpwzDzuC+57pSlfO+bB7h+kvEe1TXOYw+53Y+9yQYK
lAl4N99bV8D0Q2/oomBMCK+hH9NhEP7sTcH45vCsPEB3MhCi95qAy4CeaF3qunc1
wQNIjKb1+y+wMDVPij+Q59BmIAbZKRfIoJdDQ4r1HiwyFb/eZPyJE3c2TjsjpcDh
oS1qUFRYBn+PJb8XzmevbnKT3idV3gq5d4Ata+qF2qtmaf/XBbK/ZnRjf3oGwaNI
EBfQP4GlwB/EvD+xR2vf7SaAG1N78332cm+xAZVNVZnqb24kACVlIWZcJjD+JHeG
0n2lYx41EG2knreLZ909jtoOfFEcqmJUI/C9iUrGUY8dpMkm3PjgJI8pCywv3xXO
Zf+gkJGr/OaidlHizVOPRsRzXTAsNjMu87Vdo1pcKq/2dEKYCAkleYps5xifxiXw
Y69vVTx5QTyTAv9MlrGUxMhvi01Yk4dmvUvCs8huVh9f8EIsGZfbglLx1VoJRtMr
DmoLNPKpt+0LttOuKcRp/NABurJhg03ABMvi2Pxa4F0Fp4qzGdVuTlKjYEBHLyJb
DYqRis1bKySi+fG5OpgqCut5B+BT74C21nce8xUFVLvDLcdw9ANlUpsyPoSH6iPj
vsrhMeXkrvhFc/fiORkQL5XVPYgRE2Vjk80/TUudpeRqlzravUrn4NDD52BqpKFA
VT39hPOH42AISVK04TVxM1GHBfd6G2WXqdKNq80mYGoOLPl0zd7iOu7zA4mSd3W/
/203obFt5Vvoyqq8lrSS+rIk6iw8ZC+ZrQsQt8xWWUimX1EvfUnEHyZQMOMwz1Aa
hDTr4KAkCIH0lkR7DyY/1xIbvexIvj1UcE6ERV+UHPHJNeKCIJxBLnf5tVZ5QTLs
4OCvDkYFXGPtuQkQ2kjoi4NyklCKL661XeLn971EWpCkPPcE2NUSovK7vXR/UhrH
IDvNT9SI3vHz8omDumrQPLiBKXAqug8+2KovHZuaad5Y7OqGGgr2bqo7VpWD50U6
Mrxw3tSYeaB2JJjEHQVyC039q6tJ+TSe/uI1UzSCT5kk9gsWBKnggEuPOcWdOTSe
VQ0LtQ//YBKWVXCnuxXArCrGgcSF/Zq2d/qFSHndfioUTUzg9jfJPrMLDr4JuIm8
EuJXJRynct7T9ID8LMmtfWPbWZFODnMUNuom2TdUR9m944ghuli1gPBVCgPHga1z
+u8fpLEz50QSsg7dQLhI2O+q+dwycnOAJ7GfGq5cb8MbYRt9QRkeG5+duwbiLW93
OIIaL0zFigwP/N9vK7ksc2p4NBpfuYc/OAploTdr8vLHLkxYr28s54NSQz2RQxIu
ZUSHWHx4MsSjbCpa0vybCB7pXOWwPSYM7qb64PyTgvUbY55hkZrmssC6wQZ4G+Jy
qT5RML/emEsN7v/mw2lLG1jsmliaZwEi78huZ+MfQOL7wWVrdTL8l1/8WdmuCOmQ
bRKnNByZ7js32jwd6oDa6B03MjSioyofuSvRYHoNy3XypCTQCZjseisQsT7h1973
bMVbQisHG3VqvBmU+RlMJzDaQlrouO/GphrdJZBwpspdLFJrsxqNaPvcqdqHGSv2
9BgrTVkTiHCV69Rl0CZ35uW5Xvi7Um+H1TkvoGeLL/E2HZMEo0J87xz0Jpva5fpk
+urHO9R/XlMIDQsjQGuLx1uM/hxFen/Nhf7PKP9LQOKJ+Vjgfh1SBmsuNaUfz6CL
49Qs5oagvKbYQtvMfSH6TK6mgRFREC+OZYWtevE3aTGUtA3HYh72KV+nzhwX1BmZ
8o4eXOUrPbYJe+twNHar7B212Z+uKSBQhPqtHSTLfsnEkvTpf+UCeiE64tqlttS3
JC3enxZ9BRF4wsGiTrLsA5o1K+b+JfODTORxWkA2XtUX18r9wlBJrpvnfhdBIwQG
FmThmxvVK3MOLlW4uJ4kzCL/w3gd2+NMPpkh9Yga/bvZzSbm24NGNzUfyonFFsi1
actlqPc+z77Co732h5zwYERdVnnNEYOAsXmkjdxQ6hg1xmPCdFeYLAIqPhCfRjCF
X/fcqxwP0QzyWMRWzYR4IWYCi21ILmbkXBZ1z3wsGIdfd577tofHvSUQDob468fz
YD7vvr1yoPKDcmuiYPLDnH/r1WxCwYbImVCbXnV504DQo06RQmITqGDYNvm1C54+
zbwX0sxrxmRuP838vhCjs/gDP/Y0PfbfMd4Uynb39nyJZm3/uc+nxgGQqRDOJWEe
8+YwHoMrC/3z+LX35V0k76YSodLFH26RqD4ZpycMK2VXauEOAUK7l8S743sQx018
JxW1EL422ga1Az0fb7OYyJX6yPwVm+HeyQhTlxkGXg0mYFYvGpENc99nVqkgiFm5
F6O54Da6k6EvLlSeI153fO/4c/8th6h/QAczlMiqwGTwfERyU+3OKjZBWExELSF2
zEtL5kWr9riaiwOH+DCSmS9jOXbCUUejPeqe+DGBvEnjhORhLncGanmhcT6kZhvS
l2SkfAi+gNyPZd9b+Qc6De1cPsmriJbxekvDIYD7ngXrMLyFHB/1/rzDFO43jLiX
UwlfzQxVKQFeis1jlfyoSGn3oOZJT7YP8+WuNCpc0Tedi2BiC1b7xKshqMYD9Rg6
7PfLRVbfOQN5bGXW2msjYysEVvqkTF4T6dJuOhMvzq6ziD4K/WfZn3dL141g/1EX
rRKsAHCRI4hVmcxiYedIGR2xpq0nx6j0Qd29gQN6XLvXIuqjgUCAKJia+WsFHAwb
TXqFPBYT45CxdKOg5tkVWEoUc/ub+sWxRTokxQa3dhzrp2T1P0RiqJqAARjMlnxF
Z4NlmZMcLJbotfJudbYDFIxJXpnIaWfyA9kLeHKGr7zxgSdRfO91cPcQLiwNPf9B
yPD90v3m5cnDMb5Q9e0/Z5j/iBxX17Zmozina0WDdcv4pWyffpxxjh0iTlRVvK67
nDFYbSn4hkFYrPzZrkANcuDtdClU/xV/ijuhA3jFUNIzbg4mGf01bED6ezSAw67Y
2KbDMTTu1bAD2cU+tp6FGLAa99Dy5oXIN8IpOa2yA6njcuUxGxAyUaCep9Yof0Ph
9OEpvZ32Zi8niyVLwa50xQTpzfNmTVFz3BYyqjWzygVp5fATbEjR9powJOZ0AIqE
Ieu3nlwdp+IRuEemFD2I09f1zNfkCr/8z/zMwrHe2Vt4zehH4vwf3GhKgaER30mw
j2Pz28TFcuaL0sLueSffR9NnDjrqFSh2fmobUP0GodLIsxeJq1yDUduCJ0bCGWbP
1zmVzmRaujzyHbfYeXj7ed/skU0JrBmBZgguWLZXqSH5T3JNp5KvnLJmjdcHan21
is3jB9AkhHsarhZwjyOe+4i42wAqHyD+OeAggMjBfYn6/krmnlpXcEBsRqtoBX9E
Cu+1nuMDNfoMW4OAINo/WB1Ou5EN54gBB2Wu6y61+GTShdGLayabiEvCGipg4ge2
ojJCGp0auJ3N0dWFfsdUKQZvT4QPLbZpcfRaQycWi6i8UF2UitEdOE3+tr2Pt9I0
xKyK2O3Ix19JQMeTWFbG1FS0Qwmm+7erREedFQ3td0UYkDhGghN2o0KYg5t4d0cC
daJANwt/8Bw1hX+UD7LITftRP09F1iS+1Fe9VAcbY7RxLcGp2/vlmRZXauf3CZpI
1thTXHEyCcHTrp/2Qgo+hul8DpxPTqA05z6hEWhqdEJQC0kzNDUAoCECUsSl1f3x
2WEYZQWZNo4OFhY+dtUFW+ijwnnAwy9hsPqf0NgLV7dSS9B/66A97Q1sKZePndQM
F0OH0gPUbkFZ+/nfxGpM1NMf4JYgPu2TTdN1u/QusmdaxtJ8krIjlhnrD6ATNuWc
RzfFjLrtfOPHpxe6MpYVIrJKlLeyA89hTdAuLeIfQstQUDVJbLDTElvUy9zFMIva
j9b5SljVP8XvqGJvnLj/gi+arRVq/MxK/rLeV+Vz7WRnpomWtSBUohrD3pf5U2+h
jg/AHIJ50zO/G/F5oKE/SKpgdmtyZDs8eCKgulbSgUAJU/VhRvNjaaOiwRl6emBY
fmjodVs7iMcg0Z8whTes1eDHY3e8BjH5GFz6uSUV7fHGsuAHpCSvUREiJKKTbxRb
YAJW8x4e147bHWsx9ZaiZK75CV2JoVCJfmQdX8/AE5PVZxhD18Sm4jl5Gcw/ITvL
Tle4+GxGi/d4p8SR2MPhxqwPI6VGPAE0GbAipiGL8v2MFlgHUFh3xnmynuKNBlJQ
O31Cr6EoPhJqJTTUS1B7kniZoivOmzlcWEtaxrMHJxSFLJahy8VPVzO5G+x2qKB/
Q09UKc/L5sHXVQ/lzl1PqTIhsBlsxYKgSUW09jdIpGU9yASj7hTYAuoLMdRBwgRm
XqzdJnYsS5/WTdVy/torWCtaL2wQ95aTXhEjJ4af+/y/h3c+CYddJiJ9BjhE71HR
X4WGLdx6U37hK8MtAu4lfKf23cjRsyqfohPl7t+5GU8pRaQXR7Upj2syUK9btR80
4dicZSB1VNYUsH6nl5Q4L8icgat7OA4EVB58AMjzS+1tWi44p0YbVslNlZJwyxQ8
qiJCtwiBS2K5IqOLdXK77fHH9uVVZPmPffRVHldNrifqCkbKKdWkYUhRbnvT3UkU
HznxnmMaFcxRSdzDB1h/dn7HHEeXLxiaIQGi6fsO+0XBoBMCzSsYHKW/1PqnRAp9
YYn3/w58UP4Sb/GW2zxvcLtKygmTyuoJH0lD16CcU4w0aHzfzl/evJXxrOHnF5Le
veD++8ph4u3K/37coLHla3JNFE4Rvu3LNMiGFuvp9+U+oLwRWI6YIs6o3VJ6+iHS
zwvGdHvmBz8LvAl1b3ae+seG+sbGmkrGUlhr6QEE8EiEkKXQnWFCi9/SqojjkxPH
bxA1L9SZYV3vyDkOj+AJhn2oVzLuk71olMBhKB/akAqNxUF3Tsln7cvZXDpuyw6m
HevBKeqXMvfcHGHnanP1ioTHOE7a2do2jR7pIEeZj0nU/dVVP1t+dX6NGH6urq2s
lLhlDTFfqBYCnKs12CS8Ruz2xIssxy2UWT2Zm5v2SjQTgdej3X7e4FUuG48i7Yof
5Xru72DK1gKGs8z7lGPtNw9u1aXbxtZ5BCi89kNesIbEFlJ/jQociAxIUsIloR+6
SubLgcHx5DtkF9HJdmr5IDH9R1ybH+10frD4AQ0CxL69cjLIgxmPvIfZyB2xiqDZ
YBu6mmJj3MtjnxlBGBoQ+o1H/0yfUCPvb7leLdAZbpClwYrkBRji6ZrtjU7jY+/Z
z9H73WSPRs8MFahU579TwuWgteIowcEYqZkDdlFkPD/QYtC30K8JRdpFsXcB3QOD
ATqQ49u0TFhXGrAovf81psjginSAzHXRtPODtZrQkeDpKztW4awUl7M0Kst7mZTS
5xUtTjpKI0LwKyOyITiOx0nNgeDpMj1/OuK1maM6H9qj0GCFGlt0BNGWJO35mEcd
GpkJASmYTWKDz0g0Y/pl286R7FtSnn8/c46h+6xFKcRRG5HnkHaerTkU3khxv55I
hr+BY2I6iP6oXsY4VDvnSGFeUyY5v4TnMzI2Ojj7Y89NHVnmMVqdkUgUQewDcT+6
lgSrOYqCmIorrMTLLnUEUwCQtpD5aL9inFpo27duOS0bLZHaWy+mR91VqCc/AWeC
x4DuO46XIJN+3zAiu1U9uGipezdPxFlN62PsfGx86kAk+uYo7ptWjk8eTJrlwD1n
OUeSq0Z7A0PBS9ZoGwv7yObVHQdJ0RswC9EUli04Qytd1QUWlIEwS1vOnVk0rxnt
m6ESUunegRjpjzCG7fxgFG/9aR0y2riKSGQKRKy9UIDfcsWApIxYaqPpoCmwDWKa
gEpLhKTsiLaYVZdMzm5WUlAGCfO35IB5bVP6vL4dB88YenJNfDl0NLVs9hxSRs4o
q7vc8D2EXTCjNaY3+ixsXKJLdUFFe1dq62YveqN9olE6vtig1TPgmvnQxAgAc5tZ
JL4zcFjNb0G3V6owDSKtcuQgm1rLJmRwUFsF0p02XM9zghkL/ZzHmkbTpq5PSJlG
Sizq0O6MgGEXyTvhplVvRnOHTsY2sU2k3Ri2NJ2ulBDhiIda1UUTy65D+IJ2O2q4
zqKOAjnYQhcO19o4G19QnFcsZ7Cql5JMHKzzBIfWpeetQOgO3513/jmoFZEytFpe
fEBCQ8P3J5+wa02pUVAYjdgXiIxVf1mTw0kgD2lrty+8I1n6iT1FrJ25a2QYbHJe
wmdxaIwBxm9d1EazqAsvcP5Y9lx9kdROsj8QSsTxNwqcQ/dYIGSN9lPLDeSEAT42
PHneQCnNswH8Xyu5EJikX7jXvKlP7hngLhjawNI+gPQLUTfal2m7kwsRBMMRVNH0
CCaYuQ4RuJ9K6/bC+MJh4NiDahNdDS0ANei3s+6vvSgMcU2x+zzmeFo6xA5f16C2
2MeNIGNJ38BgmsHHcuxprrN6eOIxibq8krARiVUyiEcd35Tv+NEJZnszwGv9U63B
BtT+hjh6VQDmH8m/vtS2rhnGvK3omQQopmcvOehb27CLdNK+jTEhQM6Rby/POx7R
10q8egDZgrumcL2eH2j4ViaGb9o7uDN96RPrwJqAaI8Z7x9+Fdomt8S2rYVfs/qZ
KcCsuvRFWz+y5cYCM0L324vlifbw2bDkU51wqxPPXhdxmHXknuDvrivFBV2w5svq
6rJrEB4+wjM6QB0x8hNB5bO3FZtZGZ+nx8VGicov7iXf8sJy0Qj9sMAyZMRed98M
SgOspV19MflN2BqXFafuSQmJ8a8O6zR3XgodazcxCRpTlX8qk3MgOoiHcFwaQYXL
qiXfphxAibOBDpla/Wy1+uX39efggtB/KYMkLGyFH/L6khYxl1tRHSLcxTSe0K0w
z2aYR0pjJSe0QZTuEt/zK52L1wUgUZNqGddokuCAonFvDqgxgz7VaPf7rZX6mhs+
sRtS/9vTbz1MpSxMkVlDL1oXhcR5fVNU2yQNwk/JsZKr+wzb+Ik4V/YDrDMpC94o
U6hv7R5BRpTChPWZjknY7JU32kWd4xj6T9mlDujriUMzUsdRrD4RI/IxwzSSPFge
85WCBjrLI78Y48lW0vIgmcl2JeKiiMZ6kGg6ZOqKQ0DypjOyXZRXgFq8xRfKQQFE
DiTTwD32KCYwC4kzREAGYo4RlZ4CmHqi8hql27QDL5trtSILGPddfWRzrmujo+3S
8i2TK35GRxkYGoFnU7Xj8WBdIgx4/zAdikx37RFsxLobgUbF5L7oFXIYX9oHG7zK
4sK2SQEs+kUncUopippBuMmkm0+DoZGXcwVlQJkv6T4or4aE877kZFH4+DE4po7N
xSEybKw9UXmjn4PlRth/fbpHbRB7CxAf3dwRUm0JkDk9/Y6bU9VkkPUzH5+6ocp/
UzTgKIt6/DENZmjTJVXH7qz7vXwmNxx6592DgmWogfTtM+eEuGOANogPHfs90YP1
5uM1+8Fp5egEZaRQV2mam1Ud1MJE2XZcHhFQY9/EhYqQHCBnXNPx1gWHSxE5IJV8
eFHjqAu/8421zMktDWBGKL1PPL8I3G8+rTk5gIJJIJy+9MG0DvoSRlCcZg+RD5EN
F88YljROHm1prAqTdx6T7vqm+IeeUFZ7JAfws78nWb0+1O+LSH1dyXFJ1QUpaxAf
1Sa/tBOhgrQSfMkQTZEekFsApG51UPgE0B22Rhjt0Nygkpl2Vt5/ZHW6CLVbNiRw
5T6OLTdFiTdgq4SXgT92TTIFWx/xqCWYpALZgDrO71fMkgJ+A2TObnIj8NjREn0/
k7hfdEESMD4xAwAUXn+AMCpUEQw1coX96Pxmpn0XXqAy+SXLdKYND9DKy/As3GCh
9/mMXjAzMOZhzQZso1a44xUKWhkcESeNsacfxQ3nxr2GNKQy3tQ/6Zbq9qnjUpkB
ZbBx9Cm4H1ztDwH2BSlCQAjme0idNUa7+4GOJsM8PzPQrvQBJwRpoA7ig8cAO7GE
WrMoI3BHee5LrEI/IGRMAoivLqD8C/qnu+H5TBBI17c7vKU2UsewGn+1Zk3vTz4u
Z6W4iVcr3moT4JsgTKRjTgAloyqfpkZoR/HDWmjWWHe9PoIJQ3Nzh+SoAUk4/BXF
5ImlY9teRf+mvU/+aJPrwHJmOmMCrbRWVewmtqU9TZvYPy5YlZhGIZSqKS5wOAV8
8HgHkkCF+hESzTRGQ5oMlGwiwp9rRqNzKyjZwBte4/L87K/Z3CoPHBt8TFrfoqtG
puGWeCohEDxRzm0Caxgd85OHLZFKPL65mhRKg+0VKKR2OjmTkmMcekcg/BFIBRMe
Wz3pkfPA4ClFUizQzp4+TzsfMNECw/ysjHdD8HTcYgZcXXhIr+xxpweLZMntUVX5
/+7P/qio0DM/YR5d8k5ISS1k81z4MkAqieorqjYZSz1RPMysyKeUUlEfvcfaUMQu
PMHC/Ejd4xgpTq/izjGYgv6BQBpwpOFrcA0F2NsamvrGz4vNtes7fUWJee4M4+9f
1/T04VYCA5kkN3rFLTMjvYtmPVUcOc2HAZ55r1LAt2VlCzhciMhiwLHjYBXkmUAn
j/U8NELBT83wkK8jJfZeJj2BMA+xK135Sr6+hv/SgwLdGL7G8tI3B4nX6zgjG94H
NNoiLJqmfOnAHDaXFZrGPdBQeuvvlRwm4ISteSf+jsvET+OrVdzqyv/ZdDbM8Exn
Kg1KxgH+e+RztSAtyq82OOoIll1Ln0LSclfG5w2V2Y3X8FQJat8cghN3R/1j530X
cf07R3Nt/LQ72OE1j9wVT9kfXvGrI5qjgXHD56YBXzLkKoqrlYkiaVOtlf4Zsimi
d629JNBu59bASn6PYYx3NSa7zLJt6TSR+zGKE/0I216jdiRWndDJDEvxZMwcx0o7
lTodt/rV2xAtxfpngALgGeeua9saFtHrip0gJC/UbDMrerXpRMw0kZBmrH2KUEmS
cf7I9RKV6W74SMcsOP3lgc9qY00Xnom6cZ/USky5XXK6dnodAJET6bDRvuCv0wFf
l3MI4lSqBT8lcChmL/LpE/0XedWpq2zDUfVu/gz2cKr+igAQ/xLy+PPGqQ8rkc2a
qPolrnEntD7nxU1t5OcnVVbKY7QYnrIVyAa14O9e9NT2PpQd9pIVociFGrHaG5X1
rFyPXGaycK//zmK5DmisCcHYB1tn0wpnvK8YAf1eOO/NrI5gmpGnomLmQ7bnty85
t2mkgKFI+GH5O7bkEhtWQ1HqYNQ7CqZLkK3jZXZI/L+2FYtOpc6/eUdW6aO0YT9R
TsQbSsaLlxWgD+4UD5NFPSOm3FtmqmraHuL/qb453evUwIl6uF38wtjaslCyrxSX
wqnoCmA327psdYBjGJDc5hGFJBvuGOQlAR0Ha7jExOqddffHnjsagL95yYBorUJR
iGBOm//3fd8uUIp4iCg8hh+jirHLNqECuFlTe2vPADW9iOBPqeNzbGX34LVf80Mm
v6drJgWHKJBL00gWso7RM5QW7uqnT7vHRuB2ZTufkcjRA6naou2FiqRiVYpvo8xg
DhUMeFtYtCSLqRd4shp/7LkqAZzlDQjIdhfSDwgUOKg9drom9FciyORtydl54PeF
DgwQmv7ALB4/Kvmc627NkndNzp8qADBcfld/E/lLnwwFFW38EHktzrpiFQmAc3PG
cb+qvl5LC4OvqRdHUHbpQcqZv6w2Vcn2jntq5zYBDFlAHCZ936KycaMVYTSGKNnY
PpwtwJgZSBgmPLv8Rh5PVmxFNl+CMkAzs+lZQ+4hpIq7cqaGro+PCGv89LPRclpr
wS6op63eW3+pLv1pu3kfqn+9pM2Vcqg0nCKNem3DSHc73Axuiqk0cxCoy/bJ6XsZ
J62nnwAPRtdUsQxaWv8h62Hi2Im0y6ClKYm4SeiB78BC2i3agzWln8x9+QELTKGW
auKFeuLH62TPEjyklwFVkdwZTWUIrEdLCFF8oVUM3SybykkMJIB+868TbLmF0Fe8
7qBvMAZkEQC3FzP2+2NBN4Rc2R7EonjisRxjfjDtlexFP4ZGqhXBwjOdFMOU1xU5
49WNozVk06rUO4sHyFaXaylO/lLSb+wfmX1lXTh4o/OUW5PUWq8hKOHIKFnxDm3P
xds39pBsYCatSMy6Qu4NfeXU0/gT5KYa0niRhC81Eud7mtCqKV2fhbqGtH5MSicH
t6vdNSX9+VZn65jtC2G70O0jVOvUaIhH7ZWZQMzq+GewOt3MTizXO7lhWV2eFAw2
ErMieWFSwg9MLKz7Fd2AK3XJo0xZVbJNYDZQEPEN53WGOCtKSeyLf2LUrsDqs9fj
lgxF5j9awPaKr6caSJCECd90D9ZgipJvBT7NEnMIpwJIdqYWr/BzMMb5ey1nmsR2
XAmzRchOnt7sg/iAohrA4q/V8dQwXPvTA/Po3tNYPsmXwpJpCvKCVJdYVLxFGx9+
OgnVEvxcs/LyRPIbFnKqohYoYKaAm+40YZQyFJv5QANF0815BErke+je8fqPyub8
5FHnL5BFIy0xQ8jIFLC5fx96bjC3V39FUWlCRc7+nM6llxUCNTUuvt6RS+GD9Buk
qTQUv63W5CYrZDoQnC5Ax3a4tPKqR6l9Ttm2zdee81BWzQMSAM4VIljGK6kCsvh1
X44o6EXivfwbzareyVhK4HCw1KpYjMyxshB/GVViKtyifRl/brxtnZco+tI2y9Oz
N/aQc2MF542qtuvMtZe5bt9GxTUErCsyLXmUeJIFNrfRnWHFBufA2olDjUDp4eX1
LuudGqZbepdGpomn2agc4NY4Rmd9z1I8YttSesyESJl6nWTOgFp75Kb5QDjXvnSI
csERZNqPEeAIIIjX+xEmdWn9RaZzSgao+tv7hg80TGTR9WSkpfG5fCLnkzhUlp2p
9XsepE3cES9Cobck+FbKJkq6wF6WKAfeslRVM4ao1VawWRJFNmyEuh6nDNDrJPD1
AA81sWrmSOL0pFFHdWPTmdUlHFxrBnUrhZQStNKPsu+ROW7OMQPXg5fuLoAmLPiE
15DRmpu6i3Dd/bHNzLUmOu11VyzvgDr5TcxV5BGEav4gwS1mZDPSpYHoal2PLJkT
SDzPPumgTWp7yWzSZZsMvqDYmKywGB7NvWe+S2rOSNIZl/FGnFVIZr4FrT02Z3KI
fEtifuzT0AZP+0ZgCyk7nqyQQuSOoGnAwTYaGEh7Wdg0V6hpXJ4hDQZoFyzKrQu9
pWEOE2Kg1ildyQdbs0pg1qmgqBuIMq74T7QiRaKRAk0HDfJbRHzDtFGV93W0SX+u
CJQGKlxdyEnVoydT3lV2J1YVE+h3X8en9GO+8yEIxIp+n3osYDD+tRbsm4RBA80/
vmHvQPA8WoZy2aUR+KXJ1fp0oc1jHsHlS5vomdrSF0Km+6zGkVu1eJDiZUV/Ozss
X0/gXUqxelPMVmh4LgyOSzonnjZNuvL0ZGO7ecyj/afNVjH1QF9NWjrTBYvz2n0r
1ZPliF2NUyyfNlixzIcSr9Aq/YcEHFY3qVTnnu6wfak7FiMj3LBgu5KbCH6qPYCd
U42FwjbDjRW49rx3JNj5c+sCRPE5Yy65ikcdlhh9bwjgZkVpXfKnZKEDswXcCs/E
aFjNumjdSuf9yClun1WB7hQleGH5ffwLYhoJnnYHfyp6ELw2oEey9dTO7qTKe+jC
e5S28+J+kPOVaN1hloRODn+Fz9dJKGakmBtahXGGvOmDcCzdhOv7NUnnqB9U6Sw/
Z4k0DBNNO3nJbt4T/ER3osCI1gO18ojG977GShPU+jCV0IZ0/AM7fKvogOcyx6lz
wbs2XqVi11ImGHSLQy/8ZSzy9094hDsrGmmEQYepb83BT1UokGAS184r8HiP78TZ
UVW3tyk6ufUQ07sQve7VE5h3UK5D/mAfHaA7a4DeuQYTRpAo3rNP+AcgXodU7jZO
KXJ9AgieMl9UNtWg3PDK5sOyRvqHEGp2awgZtEBMsl8P54mE4YNQDVXmdD8PjWrW
VtmZDco9ng5b437ORb7RnaOl+eAYPvA/DHY5Cw21C9GQ9Q3Hlgwl0XTsiw+7E8Zl
STrgB85FRAoMtW4Fdr9H7r7bVJjaeAlZiJFCMJDHW1ikmnHFMEvr+b1wwDGfVYU1
34JHrWDqiBmaaLndWiPsUkmFGouAyfZEH5X8bygdTb3iKGMIdUkRZmUhRGyTRYNC
sBtIHdH7xNgfEfFHYH+h/UmH1u61fTldH6WRWio7OhkGnxmYcVO0MKsl8iCw8pIR
luhGewAGU1NbNlWC5edR1y2FR5chse/82XdxdI/gdy9S5mBrnNIaYpHQiJOLV4Nq
8HoH5eOhKK0B7QoLKo9NiUB4HQhW0PQSbvBExrv0iF8fnXMl+bCxSO7D9ugNkMhD
EEIA7rPCUtX3McVUmc7GUxXJ4DK/heiLS3D8NsUW4L+LeOomXvJGOeNqHF8WkpP8
kuPIlOyBcAO6AEF4WbmOgCTKFfABsqdc5b+A/gfbdInlo0SGqLmkSReSOQmOfYfo
/WZbfFMExfmENiFN9sv22DD5gvHHx4NsCWwL5Cn4xyxb27/VOZZBSTIu7FTb86Q3
yr6TaFPWU4YEp9Uhf3U04irv+TzUBB+ajgVqL+4KNll5Ip47+7HC1wjxgw2KmYay
BCIdmMBae2fKywLJsjXTIteq30B6GbG9Lgi+M756N1w5k+PYgQtUUbptekk8LuSl
6Fbf1plddXm183+/kRoBlanGPfIpcUMqW6oce03zGh/ybsIHQzlrmgKB9YbMWBTQ
4RCs2mGlCyMWXA0x5e7byVnRGJUTX+QWx+yU2iCQTNkctW0DdLUuY26FHP5BNUDQ
3yc6JyL3CzqOt/eD8FPv/wy2bF1wzgQ9e55HfI9r1W2KSL67Jwax+UT0gXuIFQ/o
EejGqnU/DSsK2NV1Ob0MU4+hgIIEeATWIUoE3JsqQRjMAWxyjI9/VO7KNzLdtJQO
ik1M77JmBqXJRQXvB6kD52gRV/TdsEb/K84ROaHofwezcaJbSnlKHVmyAs6tpByL
ZT0+VDHdpaVGzX5Aj5zA1U94ghuRsHkICvXDxtZ8mQUciPqRi+d6uAguekvr2T3n
zOlTN7FZbVr605EAtNUJ5KqqNc58DVY3QCnPxb2uV1iJ4DSU40VIWt4IHE+sftxY
a6dMnGg+FhRu+99/yi+9Z7e5b27vVLwUEzS7/GvdbtY1v0rS9rYwnRipu2vU1R3y
+rCw2Rg1p8BIxrRxvRo+AGfpciWcv8HcYoLt3EY+JDfU0UaIYidTT7M/QU6EqaWU
BqxSdq1N7Ix/mIO4a+Oqj4uvbqqkElVQ6xoIkII7Udrzeq0dWwaWCtQD6crQdo3J
lXQKfjd+TSJ95G1gZmbKxeGgVo6HNRODjwhjsBa1mgCncrjSNTRMtdJikCGNPmON
HQdDMElhxagJkVqG0NxVuSq0jYzU4sTyZbM0RrJX1+VQdk68TlmYPtHIcACR97MT
rAzccpJziAc2pUWdqV01rOiyfx1e6+ZF5700UxDdg8fjkr6dKO/Z3kPEXRPV118b
VzavlTtWL5MiJvko3h4+pdcGO3h226rsHHGNIS/rnn+xTTIWiEgU+EFGpy8rrk23
a3KTwfkOLo/Afv3FtkxiN9azSE9TS5BAxVd/brcNdMBt4VxnOH2xagBnpSuTIvAc
aHX45NZ6CsUJuY74pGjlwR7XcOiqdZLhTNUJJNR7G/+yxVCi1ph6/zur+8TLQEsm
Y9niKxD6/a3W45nUmMCcGqbW0yOSUA84cadwFxoCOrq10661V/LfrVo1V7ov1Nrl
BuuFG2am9fQQntznjmyAXg91XPiLqKLY5p652utuxbgOSRHv+bgAo4BnxvthWhgh
ilSn+/vy8ljX2JOSocgd6X4RaiQ+OxMPylNW2lS8w1tbEFXodFcplDHFkhe6zahZ
XhlXbrErOtR+PjVw9mQZMFMFka+QlA8aZWxNJTVnN5b3Ua6MxZn8E6IhpX3FXcOD
B+Nvt2BsWJkYqFwZjuvgNfbvsxkhuCfdk/XLBFjP4lFny1GyKZSPLEXbKC1QI9DL
2ZKMQgQ1PJRHEpws5sZ2hIooK4zlZlMZ6v7ylJKuR3UGQ4GhQjT1UBwTv4SMT5EL
fk2hFqeqjFmrdkXJ2dIPabWe0TpIbSIfA6Yr5zGGsb1oJJQ96BuOomASB/MBo9nq
3YPYwl/CM7E6c9Ej6YuYgZMk8fI+LQ5d+vQ8ymhaufSXsQxwdOO4/sLyYWVKXGNo
zORpQHRjzarA2vX35iV8eAfgY52uxSHRtUFInEvolZwyT6V7wSaSaaQUs5ARMWLW
J4Gz2E3sV2Axi8xpGDZkprVZAaX9O8o96xeq+NEEiwuI0aLA3vqieceZTM0vRmuK
NRWiJC4wQ55yu3Uu+qwWQiEJSpjCeoAhKqyCAO0f8dBEOWH1Nvysa8ISxGTSQV50
bvv35bUrGCC590oyIDivCibSMD3E5xn1dkvxaBv3enDUBtMoZbhbuv9GQn1UfzGV
uGmVuuPoAZ0dSSHrW1azp/kcQ45v0f7GKnRpTgG9htXG4Xvf8LWJAsWiQPd5rQwr
BfLIkJTJweemQwVowp6nsxdKKeFFwhA75HS48N7J18KbbGHYugkA1LnbxQtZxfVU
gJhLAygpczuAHv4OJXDUYHh4lRnekTEc+Cs8Gg4KQSjo2PY6j9jAZFkYhTcd201w
RyDfVOsiZGIWJkMOeeOJQ32LWFH7IP96eZPqEwWEUHxx/mt5E4/MsqERRQ8YgIt7
P8c02jUwjoHvk7I/Wr8Zbpd3rP67hMbqVUyVQYC6MYAtdp/SYocOiyWh4Tes7PDk
d5DNqdeIxUfP6BZScDwn55GRRBcKqyvBGFxI6WA9f6InWIx2nUVPKuivz8uH2sNr
dljyVuk4YJdry8WZ5vO8ZmpIkbaVX2Tpfq9jqHaWb6jnNutmuRDj1GoUWjO7H7NI
B9hiAfWyJsT08Snx80q96z94tQbaZgwJ8jeIdC21rOAr+L2d267ObC4KgLF5yUsi
R1mobojMYH7ANh5m9ca6FSWQaq6B4J5wfX0C3xDiipAgtcAYtIRU/9axUdCJY0l9
jRF7EaXB2vMa8t5nUqG4NdnKWTYUXtkw9g1SMZr68w7c/sEX6ifV6VV8haESc6KT
PeIvr3y1rmk6yNpl1JO1RV+63Q0Y1vrP/irqYyAqvYNXqcO5a7PRn2EsiixjaCyl
PVANQqsBZHWyDPa/OicAuRnExBYhLDCL/kOMopjMoT4L5qa34bpPLxlWXF27KDsy
+qp1I8/vjrf9FwICrLK7SY0B8MK/dOjum7+Q6Qe+3Dfk8Fp/0MVSy7oAHIGcfooq
WcRDDMQvW6OTUjOq3f7KCkB6FXHzP2WBDNr78lTQwAG4Wd878GF1FPNs5F1/yj4x
rOcBVuIFkvpLZwYTMVohdl+WdmH+uACFuh5TPjFPuru68Kwpe7jxiJdiERGFa9/s
fllkBpjGMxtYsKZJfAqfv4s93QSI9gtDJyLHq8qW/sA+gEP7GjfTNXw8IPfxNv9L
S2QEaPd47S8ZLm39SnK+Aqo/Ai3L8iv9cR24Rcuwi/UwyAPeumK4NMIJleYhD+Tr
WlqpL2bMkoJED9rkc0rBbG3IAx/ZVNOJWI4c4C8zaIxui+1O4ZvHkAstJ/RtuhLC
vWMhX0fmWXoGJnEQ3A8+G11azbqXnsuCbyhlN0fBOt71nZSMjmXfbzj6ZXS2MqS6
XwotEUcKwhArzpoG0c8+IYneuN3ciE/BwWLPVNqcnTHUPM0MkVQuzm9OA06SZK2t
bxJOlLaIdDnmZYs73mcyZVpigwGFaFugm+plcP4iTlehM5C2TUYTtukD/sZzLvPB
g7SQ9VPuJsxxF6JyxmKk6AcV56OIo+FOxEIrCpeMk81szZu+A9+a2AO+S8pqER1I
eO/dAobstXvJNF90NiPLBDLIkvt1COhEVaF9FSdZEkcQm9xwnWt9HQ1w/OByrx0z
hU4Eil/qTOwU9s1jtHIcC28QjTUVpr5Ahk4v9tXZAXjD9azB9woO4VkuM+9434i6
ZarNs+NDHv1aPc/SX3JSDe38T3SzMwzjEDZGq3C3cYZx9OQUGnDDSbBRt1G8RrrS
ILegKmbFBZ7cSxxR5lKpHuYd/cJhzvxUarmLBFoWHUdLbajDRXdi3MyuSzDULlgJ
EWe2ruJ5DRWsWbh7e540iiA7UEjyjPnPTMSSU4ck3aTZJHJu1U8VM3HLMv3tGieM
ZJx0pXZKqdc4AvRxC/tfUVpNxVNoJDigLU5VthZKqWgCN1KYXXcGFxLBDS/PMb1U
QKQU/fVLavmXF9cuTXEYaEzLZfruR+LzRf9BfTstT4syC7kaauioAtgwkHNyfzOR
NIn+sgc3F02r7ndJiZ0Ztecddt0Zzv9poueK8z1jRruTlzEtSpkLV3C8Bkh62u/k
JCpJWCAwpmiijON681sJLdoYZEl7NWRfy6TFYXNpo9WxYAyA8scOboie1E5Midk6
HaqS3Im0g6SNGj6MePZR57kfXzWTAIwhpIoIcfs2StQFHqqJjbuqPtAJKNJ0w8h8
xo6TuHZIeTI9qwv3O0nmnSPkj0kgVWw8hRL1AlzEYJ3LLDb1nQLt5z4HU92gOU2c
LbfzEjsWq7Tr1WJU41+ZegaDV8DU5THStjL6iufKJj4lvvXNZt4kZjo7ORvhslFv
U4CNu4j5wOR/mXempiL5soiU+vs0T1quJyLEWGoOZO6uPrAu7zFsFwJg8KeMiC20
sQV+Vmi1HHtrWAMlPEk0GVBbDPUWDDboWEOh2Ni/b4M24rBtG/kGtA1fW7hpwGyR
UXfdhTEuoJbN289ULxcBiJxNL6M/zrVbVMhbO/OU8fd9l/O2M+ORuUa7rlMOKvoy
xB73U8s1HXAHdRnDKDqy0VGTuWJ46onG7N9Rui3L0zvhNg22OVdwh+AK1zaHMrDM
3unRl7VF3R7yiD2w2E8aUxqi9KBRYWKloFEi3+1wdxS6pkZSAz8Qe4jrwkymnks7
By0q4jUUq5sXovQzMXKljtqY+xy/zsDa70HZa/PQURED3124t5oQ7Oga7/YkYmQg
/7jSF98cp33OB/7zf75CoPfVNDEfZS17U3o1T15mj7jJ0tUlKw7tSvsAPBAS9KjP
PHpe1atBe7fI0NdJ5NcLxiqvWA4E1hsNtXiuoqx0Y0xkM63WZH5P8qPvCahchfx8
OFE2QBycR6MazDTRIrWcRSIDIOS9fUSOd1BqgnuWaYkl0FUO+ECeyd+gr6f39RQ7
bAjzDpPkUrMuXL7CiKbfI0wlhfsy3yS0yM+VBRXudsokvChXMZVk0PyGI42CjmNa
KfFVqz9M60mNRLm3NoBh6NCnhgrvUvRLjL6dJMFz/TIL72DNM2mux8NtadZejgXG
ywxSouOLBFWsxR7YHve+CkvCP3exhYZSoaeiZtCy74+CSnFjPrryju78Toe9ZBiH
o6+A3Qh3cYHwd6wyVTPd2Shdpb/LD4EVjGC0SKh3877hCCMZ3q7DDuciLPJPdfdb
SemTMtiGVBImOydEi6LQmx5M7SzeX1ZL6yhvV8LN7g0mcL6AjrzOmWH8PxdAUXYD
rMHk+otB3lz55BujsPGqsshxcwjZ31igLgYF/qoXCgpPjNpdYAZ313g+tmvT90nD
cMHbR1bWo0htQgbjnMcgiaB6hbqGshDS2BRhZVEOKVokOoGK2gm1bShgPshvoxPR
ryjV7q5vk/qOlOOxphDGRlEXabxvBQuNAgbv5NBdSclU0SX/gZS8x6EFYs9urG+h
IvqLR6Iy+/FzMMEJn3pjQLDjaMhwIlnrP20CZj9zdbgocKsULYbOYpqLbcsiphG2
7R3Yk4dX7CnENjpTcx/+Gov0LceW8ze6SmiMwI7OrveG7dWK3VGREHoYXWtxWNMI
c1j1JEKCeZIpU6iggjn0+nkmPRlG+3AQ+XDwLw35KgsbJ5e0dfVGg4q76gfcyy7o
mb0bBzySjk7QmAa4L23PI3JcGnk1d3THFiPa0A4rk6dvgIaqSLiZAK3uTSWYDAK+
ziGGO21y+Aqu+QRZHw6nBXqAok6YrBe5CVJaw24r2752GYsyc7WQzd1lLcjCnM57
rQFONyo5MmjMyHgKTfDd9b5KRNk8bDvKgnqeDNkI+zpJd4MXDE90x5A65R1E5BGO
Gr1VL5LpyjXjpPhhcxUB8Fp7/WFzLcdFJlWiUq9U6vKxqVumNZJnffgrEL5I5s5d
p+cHQKB00KkuBUj7iWVSRV5/feiDiYuf1gJPV9EzbFDiuT32fbESEe/LCee2w40p
sLp4ZvWYfCwPkNJTU4N5CwMcLLmkVLFznXFAb4ZYuINgyspn93qwkXg6Ot7szjVL
fRUU/L/22jThTqHyUa96rBtIg0k6hXEyK3yD1rlfiFYRrpZsgYqZRrx7C65EQKhT
ZX2f8faEvsle9OJXUyoiiTwCPg04VifaCyX0bQuT3zkc4pJBSiSEdKsrnl73w1Ay
gl+rK4O4kMlooLqoPeIbeDs4bBLjfrn2+d7DIxYotHuNWwIGgcaRlqpeXxYRewCY
6xxyGCVRrly3/rQadL1ko9BO0sn3NPkT7AwjRDp48K9SqmVYc3Wsb3Pvl8wRCHkk
PUytYbOVnBwQfuA64y2yLhTF0zxHR0NDrFegVIPXGit+3ZUmfT3Cgt39bk5mBIs0
vUqY9UY407axjAfJCAyqljEqqhg5cBFO1L5kYhWpOtmhkErXGRy4jTSyQe+aqsTC
P/6sQMz/6gHO1zTL/rQxP9rRr2fQP81xZWfCqTQf25tvx+BNKYVQugTK5CA3cD1i
EJcXQlj5+r5QlghKYQzFA8Sn/H4Dp+vcOE68cj4JOHKlwArgQ9rdkBr/njfV+Zfz
ZmJDjJpepOHjwwt59M/8C0qrBC+GG8hjWgePaCcmZKPcrhuGE9gIUVqmcQr3BVWP
GQjLXqaWL/vYAMVMOv+YI+GtKh2QqKuoeCuVOEpm0BNJ0l8qmZBpr9oVAlHKKhrf
NKfocy1KQXjK1Fx+7phLjmawDwR7qti4pyLnIEQP2QsXUc5L/zkiyi4BIXeETCNq
hJ3+aaKYSoRbu5I8LR+GYS6E5FtiQ5Vmlh/s4yAIJ+PEwUFWnGhwEvRp4R6vEFgx
dRuoaKHfblPquPSqv+74J12gGtJ0g0QjnZQmNCKX3mgTqwuDvSC3GmIEyratd+21
RcMTzrLxbTvnI72kAG44+0GsQmlIRzKfu/3aOqFEr5XctBQJ14RTDnGOB45xeR3x
kXCIEkChUlqYOjgm4g9BjT6qTzRsfCP7hfo6q+qnDUU8ZYFfFMojPNDlioU7/m89
fP1IECj4YYWNU5Ns9RHDMiaDu+e5KopmaCnpxepvdSHSam6NyHWwsHRSsOS2o8ez
4JTGvko1NMiH3OHY2yZEFYbq5f0zc86QA0PJ+CZfxlpHOs17AbazTiho3LoEkV8D
cSA75cMVfJHyaGow/5dEnm37PQsjQX7EK9nWZMraF+vUL8c3uGqHJKmF47E4GkSo
NSnUe6YMeZ0pE5k2LrKKtFJ6dLj0sFflMBKrZzogqtbsy47yB360gf0p0g+KybcW
cjmSxjLKi62jvf5kcZv/KfWct3Bj2e8xa3jEzlAvIbG25RAh8Z3npTeyzkrOARMV
hf7vsaRDJrCts+DXHL2qOAEs7gGB7vNobJ2qC3ADnCyzevenId8dxq8pDIHoJIvv
TAm99HeCjatLYMvyK2X2dB60deto4ZCEQMtaLJMzVyLQ7an2SzN5U+KJ6LCnyEug
z6at9LyELtfgLL7wFHH4klKJ3sY8rNqmkq+YROhCnHIhUiRL5u/JAlWWkSx0Kvat
7/3MwD0CzCmx2alR0ZJp6MOeX25EhWBmngYSFauuuK/VJ/sa8R2SKflLaCJi7i1S
8zPLrgXG1iOWdh9xvXu2RElQYHBKY4NVEZ5FQ6j7IpOxhxSvd/iGuIyB+mXcd14B
hro6xEtZvcT7Y6wxVlm8AiZqlHzgPu0ppTrAule1f+SRqFjIl8ovqMt/zx6aRb3r
ayt5/h+Ecu893LCc6qzarPfFuUlgA8BejkuPcXCvN8Pfm9n2kG9C8JM0CIIbdLBq
sel/NzB9KGtsGzpoipyw8EtL7DcbOGQbmWF8SdDEZTlPczrAqJ0227eoBMspX0le
HNR+i/jlncBGAusE7RgwR8+yzdko6PZ+aTakooRRBAVD4uCWrss2H0Ncl8TPxxrK
ZncId5h6k06bcQBl3xNqjNwlJKvY7YH3pBeusE6UyNburxWzdtP+OjDT5XfOfx/e
rmoqezvold8wX7FgDmaD5BHXAD6X0/G83ACHcbDU01Qtg9i6pb3I5j0MKhsT9t4v
ae3P7TlecyPaiGQ3CESfOjCqQtxbXbpGv0j8BwS7MTwpDjWtJbDyE2vbbPRG0QAU
ZBcqtRvIVgwuWxmQgumCmuxFs4MnSc5XiCYYhtEgKVGT4NgmXLf/eKnhlC6NOI0F
PN/ze1U1yaNO+s68Gw0vU+GTLNCptLlDg6nfTa6UhEIXzXGoM3zc9WoQEQzxJ/Dc
xuOQlhGELHfP6rlYd2iq21qyiF4djHCDyLeHbQo6nCqZACQuYu+bO3CRjb/zm3ou
6ixkePi9PqW8O3MtMXja/LYI9WU7JnGXHK8jv0nvIRttOCiZoNvrEbSKGf96u3gT
DeC74vtNHN/ytTKh1LuXuzOTFLShqQ5djfl6P+qwoRIWSjmdSJmpwcKvm+pV1EqQ
P9QR9yFSEsZOEtL3Mpa6IMRch8oBMmHzLpjk/8x0Bonz8j75sAAZqmf+gqHAZX/J
7FJjbusHMqq6S2tJW98Dtx+yNcY/H7rA/poNQ7GTiMBXnmj2tg+WcfdPlnypru05
Uj6YSaGdj/MIhCLsxgNVx6X6X8dE9KWOZqUYDFc4MB2549uzYnxLNG/BMGDTX2v7
qmFjPAcDzUIuStz3WKPxw/ByvIG02Inkq6w5gShKVA6M7tswpYOfQkJ3cFe7jqzp
gYntFbhmS5Hl9eK8CIwgbKi1nS4WjNFHAK25k9BTUvKiVeZla9Yf8/VjPg8uZoya
uqocQTOUv6HC6V8d+dCmezAXOQYFhvdFVUP/CPcwn1htvjtNkdJ2ARWosCxy5jW+
DBdA3X4IkNWADVSUpb4LavSENvPCyuaW0ji01evi0viGkw4vfqaUu18xaOslbW77
4J4AhpkjcOTV/xPvJMY7kcP9QmnM3pWreHWAGNUakya9yu87aYfzgJ0GB9ZcKbQN
SEdPQqWjCh5kHWBQRQE5fGfjypI66lZlPalrz8wjeK2uhVocwX/sQNMvdUp8cw0p
ti5QwNYhQ4BYKa+zNraDI1CXsnDGPimLNSt9R+G1U4MGhHNAQ5WP9i0z4UAHjc8R
KM8oFJSYR+1eHfrefu3bvUjc0Nn6KPnHfOIk45gSIKN2fvEnjQlzlGBD8wG/Fgcw
m+RQizS2o74wH/H8oSnG4uk4voOrXuzajcvmQl62o+6/o3A7AHSCdL4vlVKmDvrh
486cpyJDrJriFR2Fix1VKJYIxy+6K5K+dpmUn+03Pr23ORZi1KCYDoXQcY1uLuIz
F2LM80eS5uyvYABR/ehe/iTZTncj0vvTzIwag+iZnWhiKbcWTkKn1ta7IF3noPhT
D+rITKFRkIOKgf90N/5RzmdEHlIBozEPNMoEzQlqjAiQazKwGAeffsH4GZro2Iuc
s0+raK5WNE8Ba9ynf5dtZFO623AHXx6exxkFUuFLPudgMuFFfsmV6KpT7Zw9I3HW
JmNHNq9oduztS99KQiTZdIxdfPmKliIULHntMPTtagLqcvbjboel6SM418JtWwaz
UJq9m4iHxXOW/xhjDj+ucFxdg7zVznvQasYeDaLIBSD3V2MbLnRFCCN1gn0BTvwf
IBdX6x57KQhP/7jlxbA0AuVqVayygDJckvF4EVtss4eee6+uDKc6aPA2hLx3XWwK
C8cI4C53t529wXFarWSu9JBRz+BhDy8OVKmmRwYxccGAxRQ5OB4/iMFcDb3NhCZG
/hgwLvtaJN6fmnRGJ+zanMc0d1w6x+wgDZ7l95HGC4OzyiCx2rlT7w3pc41QLVtZ
uRs/N+Z02ybFZaRyPm/fzaMeS1EmPqpHxB78CWWCfg909UaEbmJ1iBZvzDrr1eSK
msClHkZpOAf5Kridj82apOlUqelE8UFnfDY4cjfyvzOgYXF80JDWEEOvDNBO3IV/
1m3LOUnl73jZ3Ly2vS+esKTqiiRr6XXLQhmXOT2zrBzKAXmLNiEUlJUJh1E/3IBD
o77fZBUswKwqBxAooybVGV9GvuK6pPPDASAfSpip/22ab8mDWySPJ2iMPCeWwLhI
Wia7ZRlIF1ZP4Uz4T9Ug0k6oi3o5AHzWhjfhytmPS+M4m0ghMR8w3UP28au/yZVy
8+PrnaD0PtHh6aCRZCTIkLK5MjoT2uxGjgkoVVhu0/IFx3y2n2CU0Uvlk1h8MRMh
Z2QqW2zEBHSP0qK5q9x6z4EFy3BgeuMOuVLA6leihrUwIrj10ZotjtO2GJXdhJZ2
r5SAN5VmVQ6csUrGEfTN0+cQQKzxgMIWrc4ELT5hzptpZRDjqZlM38WCkdpajBBX
oGHR0qTS1IMVVbu8MiyUxGffJ+ziOsegVas3mDkK+J4EiioryLc9D+jhTnW9Mi+Y
eg9Z2Wy9c13sRIJEuRD3Tjeyyxh9uq3VN36BJwIP3+TGneX/kjQFl4qggQyV57e5
bLq5W0SgPCoWKwtUKCINQjIIf5BpXW94W/j3A48nTSF29Yk247aiUqQs9iUWPb5X
36pa49n7nMaroXlEIXztqw==
`protect end_protected