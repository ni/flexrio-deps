`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24384 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
ZIICkMu+S2rq/yOQyqhpuo/nFJzU+b1/WrbWSICZDy1joMPz8FfGg/Dr1egZFUet
GzeHeYrhjuRuUniQLVwQg585mOjQaw1qOkAprczckxLROwDSRjAva2+i7JnHaDe9
d+U7NHUB7NQqi2Jk9adAEpGC4IMN98W3+z2+biprPhKjVeCSSV1dmJykYE+6tEMR
BOuw66o6xT4iWGpufKmmDdKP8v6Te+k63tEjNeFUkde7HDIFLHJIoLavxoiFJATY
NUre7nuWhPGcJy9vEpT58SGQFebutdK8r02/EW28mw/ITBeK9KudRSHZgb1YemYo
j56kSbFVDo/wKzphr1elqb1tYSwrcvcBdG3ayzm1kRAieY3PEnU1zx1pq3GDxnPd
0h45UQZvO1HZcRSVYPAfCdCdblxpGzS4wo+5X11YiWkJuPQQuBOC+n7J7j1NzmGh
Eox4c7KW8HngUYFXZuyNxLfeJ34RIpsnFAhCfN+StcmClaLTQ5Q/bJ3ZPG0LNSU/
wOZk5qI16S0auZ5pwZCvgXV4sAig7yxIdGCjdAiPH+QREr9bVKQJpi0H07e9EucP
fcXYeKqW02aC5YF7x56Eubuf8pz8o3/58U6XT2oxynjAOWuI+O1xxiqsC43YpTAN
RvovGJtXebP4Q7/wbASl3V/Npo0jzGzOxldQ8hGUh2Mp5HWvGc36LBxMcQs999Uv
L4f99cqYzDSzVr4QL8zcMzWDF6rHq/d1iiCpm+63OwXtr4MmJcWBNjo5wuAO4aWF
HozUyLta0fL8q13dHMnq/wq0+BKwuACklrGp0iM6MeZcKyBHfPRKnOTx5nIMgOls
vYwBA+vE+2+gr0Hrt9ArVF3bcGPqekosQsep5Ha8XtBA4mh0+KPtTLQbMYIdAefG
e7YcHdxeZ9CpzX/+KUvvo0rhZVTzzql6lw9yr7zTS+2/1aYYSozUNuE9eGmyqy2Z
RpWZBc+lbbQUTy83PjUeQbQciQc+nsyi4x4SbiWd3Zt07uB8F6fJllhRgKsI510q
qCbJo5yZ5y/CF6YPKp7H2ZdNrX7+U0Ih1BVC05plphw/JghKxD6kwE9sJZkeO/Vf
xGs6otUCYG++LfSspaluWHWFXnRqb8ydSo/qmhQ+H5mj9XWKHRZY6jNkFl7FJayQ
cwYMIDQLpmTHpQ1zQEeu4gOJs/CCUK75ss+k/J3dTogIe0R/F96nYXq9DNu2DVIx
CEDVi8rj6mNaF0v+fH2ls6hFCTUMfLSXrS0ers5yTXArGPEkohKKJvUgg25Bhz9/
QCW+w9IWNRrZ1f1/1v7XwB0DWKDlQu4kJ8cknfeiu9N5aA8dilIF3YQnUFXZHByS
hcU5mEmcDT/OyPIh7HjnwalZOEjcZSpri3x87G1UHUAytwuQJTeGKySr3sFb5NLt
0x999BBZ7MOKdppOrsTvunTg/lk3NgzBhsjbF9QXK+lzV4wyRN9SjQMOYNEc+IKg
Jlpvl386+igQIqTvFKtmafaRduNzf/z/GjYOcIDhFFMwDqDDV0t8OC0YTHT+qU/G
t7rLcfCjjkm7Eva5Qh5ltkQWxHvoV6+3uPDnmLT8eSbLpQ9E8aN2Chc8PwVMKI0O
2kIRqtPc2cBTEBstYyrQTo9/8tnmfC994Jt4dcoYpRZ9E2pxnFBO8EqSLI85XP5O
RhFEfx9pS1hOwaHMoj4CDLPbIFSSKhO8dNVDSd6irvXOnC+8uNkyv9w4VDA5c56a
jlXUciI+a0kGd5frVcxiu/GKpmP592z/DG/UYYu8dCmVg3WmrXAfgum8CERQo5Td
Wvz4tD7KM9C70YXU3mQI5JT1a0uehom5r0ARh96s9862ABuLW4YSsGGnISiltrDx
GHzw84vC0sqvUN2nCs2MLTqviKLcVsarAUbg4IbS8pyfRnX+BuduTBNZ1vBX5x4a
EMPOiEzjKXux88k7rql9CdzhkP51/z7Rbu7juV+25Ay8LOLkqbB/r1lz+EtnEi2J
F/m+B/cR0dnuLSFaV8lLyxDGRbiC5zfnu7kaJmfzb1JD0rXjb3Bdprf2KxzW/Gkd
3Mbslx/JamPUXrur6JlADyotQzAyXr9oQf8haOqwidPfkqBgqq2WvW5qvaj3W8tQ
atFuF+QjthWSsamzY/RzlbA6PDIG0G1VPGVCcAF7dpkYs0Bapy2dQqQSiImlzgyS
zHjft0fVhSsTvOqz7UzofAcKUmIK5qyAhRK/fWLLAaxIdJdtwiFq4iHTl6o9f0r3
3YbTUerJc9hsywZ7ej8jp9sKtOt+jn/mnY0pqwXgeqffpnOkFvyRwqIrdvJ3GMGc
/QlBAMsPMmOadQaI5snLFfdzjaxsmoyMk2p8IUAQNm4Vk4k53HQprA+JGY2ILHhJ
wWsLnrMplMebA1EGOkR7m4FQjmCFk53ZNZxkvTtBXW41AC4tYjcIXukJ9fOmBfXo
Sm7sMM5tEJLml4woWGIj5ofX6t7maXCifDSMtepKdEcmkgv+jay5pfwf5447VZOM
hFn/St2YAlWukla9AFQ6JE6ZvCsIJoPmIGKeVbuDUbK138SSSVH+XEObHyA1nVFw
ab0JDroA1UVb2yRHylTecc7NiSg2D6ip6wGlbDOkLhvV0JDrPX2eHIWIfTJLLemg
zcGFIyMqvdcD8mlMGt3bkj+ghz7HcSyh4t+V+ljeEixuXjderhV5Tzni1NzmLaId
6mVgdKoq2wxqeJv81o31HMi2CQX+afG9xMZmPFDA6uFPTvtj4QX9HRjMMnJO1pM1
yf6xRLRu3pHcihJIRMs2rXnh2/UaUzdifYH9gVs775UJWwKcLZtZTLPbYQIbnv9A
nJFuk5DIH9YescYHIRlGyylcfdtONkdKbJ4FSeJzh/XPJ9bODPcjPl7L3MwOKv95
1wx1Q+uP1PA37p0lnFcxSCWiLkWz7+49S38s9XUqOiOYvLuPx6pf0kgnJL6f3QMP
EzbNVdAHVOA2dnsLa+aH6COLXdCsOLmIsPrS9rrt7BST1YRAP6X8EdUidujk1Z3s
fIbrju5mzBVckrfFvpgQ+Wdfe5LjVrABiX6JqEhSdPbgcdKRQmt9sxkpEnsrOntG
nO2Ar3eWNiPQVyO9RibEfRti6/aEtyXaHmgzrlnVnuT2nKo7NRUq2m50Qbsp4RoU
JUNJY/qGmYKg2cIND3GiZHVBk2rny8yG45LONQPq7Rgz6ike/EWhuTLWlAJ/9vnr
5+9f30D10Bhz8ny3CPdDCp7fDZWdERueVGTi2MCOTZ1BQiwgFbpOFgjuupxEuAgT
sons3dOjJ1a6bYkM8QooNTRGxxE88pbE8k0EgietorBGSqX5b4Sai+GXxgtsdBzf
Vofzr2UDQdkPS26uBPMDh9h6k7zTaLFcXPSeCYAKkxLhlvDpJ5Z47EkFKdTuw0g+
q9KFb6EX1d/sKF9XBdzkT4ALBO6RY5HZrtbgRnq4wP46ceoH5Ep8SgMYhTo/5eOh
tGI5msE138xmGxDFfMvy8KE8wQ0Q77TA46b+hcBKI7i/E1x+stJl5iablIJqKhS4
7M5h7BmkQs4lE6j0YexWwWS6Bk136sIe+fZ1IJAqcbXBDQvVx++iP6FguM0qELsk
k97cUEXtqmeNNN8BtIzjaq1wlECbVSRJnXZP+a38ofkh3zQGSHehGdNZkDYk1h7o
oT1k0uL2euC8rKm8UjpVBUg3btlpqDw9Cc3IeEwzsChqulKmtdH1JTYZYMwODMKW
vYCP06ldL+Zasc06JNa6f9vAvhGMqA8raBDG67XAh4NXYLBKe2vlM/yG2LOCSk7x
Q73PVakD0DlEB5ElE2pnNUwu3P5SQur9LS7kQxaqHTqyFgE2tlXe5AEzYhgMX/rB
NaHR6BqziO58tk8pctQ59DWvyaQltPfqKIG2fkAsK2KN90mmjJfhYymSB2qLihJG
84ETDh5I5dnWiIfhOD1VnsZl8+mldvZPteGCb6vUIScmJuq5J8BeiXn6hANFOVGn
P5h4qEzYhqF7RWHSLPQoQ2idO5ITC7yDGwxoA+vshWYPszK8ZRxq1A3uyocRHwrK
TTlk+HuawbCdUPFOfxXBnbY6PJRCOa8lYC7wxBsDdQrDpEw8V1KpUOoc7q8IKJIL
9LaflmINaub/JKB9DwGKaX+gg641XKpgPSuU6kJ1OMuEQveyDczkgujJ56hR5+YP
3z6b5z7srSJnPGTfDoZXgMGnWfsACpCEi5rLHkt2wkE0KtjhJo8kYRBPf8G49YQe
cnUmIFsBFavbtB1KPkU578ZpEke71DWZrFB0Ms1c6v70PW5XnijNCVtdpU1G8vb1
SzvZi/yL4p0NZaORTSDKyHhWgKpeQxhPq8D8PRsDBmrOVM8bozk6DUKeu2eMo4Fq
OOhVCMUpdl+imrlq0Vz5eKUEBtr6JzcqSrj6qQ2nyEZxFCPpi9nP8uG/HnzWJIS/
dp7DGkeMnxwQER8q97F7wPPs5n6CW06xJciG1oVxgWNM2wNTxOss7111oxcIDAIE
61sDt1UOMYpVmBx57CJFHa2rDTph81gdIKObYO/9Un2ciReS6F99prZ6iJoqVllQ
bnAoQOoasvcsBcfPJT1VECk0elz6p+42mRWanD9lt7i88wy0vawSrweNu6ofr0q6
Hlx50Oc5iJimVmCiepWoLS3W89IjsGGur/5iFlEu3GRM567P/TB9TscA+NDe1Kbb
Z9TZqchEesXo6UIgSir0XlI4OAmXzS2oivrBvIs14VfMom6keFV9xDtkdcN8PxPe
FQozNfxUFhG8aCbj+BT0hEyT/S0bCkdo/DQEHwoFUjxQbH5AyBEv4XpeUHEePb5t
Tk6Pdrr3FvY4Uth2MDfGu0oVT6y53u7XpgYjvZyGQOQcOrOtA45WW9qPZGNmtKJm
G61iwBD2Et+AIiQl96xKrHL1IFH9hLaFpHsuZWCXQEtsjMM4CP5aqa58yRAcek0k
iHzidqQE7wRRzjIgl+sv/8qi7ajLvBhfSx4hdkRTGaUe4tkx56rdIXMNEtt0Rd9U
ixui7P+CgRIgieMirUIawKVBtFcOTsKir3sHTdr8LOK3w2BJU0xEKo8OIDYPolNk
w4C/b5A6FygFskzlohzlLboOMgwbllhI6QQumdffQVj7yw805OG6UxQC19hfzQrq
LMbkrNUL8Igc8Hx2UH9ftTCbeQSJXHQJCfoah92ZJCfnB6/vLIDpIhrjnDdRHQdw
fyjNAmrsxY9MQdZwMGGzzfVO6f4JG1JT8HiHnF5oTr4TpnK818VcJnJym9R2IP54
2tHTWtwgcwBkbo67MfcZi2HwRmUWJaN3eF0hDSdOq/doNbJats0WVbz6gn7M2m1G
QBt3XqX9i++iVncPstQ7u+Rw2Hoij96uZ60wr6K4SX2xn71SIkJx5DAMAYVhEpQj
+KKvBaH5k6K14MK9M/UQh8uDs8WtdG5SyIm0JGO5yOkPKEOsSW7exoLJqzwfWLUT
6GXLaqhIkN67d3JDefwX4nsroTO4/+edi5gzNMq446Fa4ydXnmBMj9fHensEXcHL
7hcZ4Juh/bOJt2DMfpWbt26QfFYrILcJpoMpFF0rSSLAhEDWSoJ+zO2XpTIitjuA
usx88zlz+Fep37cVTrymPcdoSFnGgKgw7mStVXhuKqVpYqedPcTUVyMNzVxgWZ7K
J6zvNQ1cMt8tA78SUpuvZ3f4RjBQt1fR6iYvtI6yV7UcqYvFloAxmmARSBd0PWW5
OmNxTO+Ur7iLmBkDkbEICQ2Shjag/sNAwv3zbjklXlnwwSNuJPDWHhZEgjDEnrzf
EhTkwyPEQkyvjQc4CZuDTHZslBpEB1DAetg4u1Y4oRjTFp9T9z0ZsqonVpML5a1a
0X+hOyXgUMjvreE5o6LP2okwsRzdbRhfNG87lFCNlR3XqEQ88fbY4n13vX/r1n0b
+/FvtJgA15SalCqNgnbjadhWyFgAiSwuhx6wAHvbtu93Msjs1DcOcZP9A6AiSPk1
FLZrhyqC/CUg+1gDXGoFpltVl+DAS7qk+qfBqNK8P7eNJOhFG5fasJXsDADsMm9R
WPsb4FkCaca1DAOTS7avtnzfH36WZIiLD0fs6XxizNARgLASw1uAqLKHgYCdWYwg
W7WaWCPg0yTw+P4G5yG1M0xS/u7W7o2/p2BTy2USvAAif9dFPG8NPqBSOiI9/9me
qHH4+BsABZNPzKcQycNMWQ6JAiX0XghbCjyRDNqBT8gh3BBuCUoeFcVBAr6w60bB
kfbBTvOIwZ4duHAn+U/KplchJ3d1hyeupsxE04ABq9FQP82fCAPHZMb90l9dp2DT
Us8tW3XYeedtBtxXbhMBUf3kXxaj39zmn/FSTnjjYGORfVSoBODWDdtFLO6O79s+
hJdfYuQ7P9GU5gokWpyk/7NL684vNmk7vPKswG8zfndBlwql6Facr4HGGOaDD3Q7
SA0+cJZ1+M0+8cSXUASmkbpzOd3favtnK9k/N38JvuyzTZ5Gc7SWm1EqFSNgS2u9
gcaPEet9q0WcmbrQQkO8SAMlA4kLtjbh6OEZfNrVjTcUQhRjJSdujoAepb3koVtF
HnPwb2dz7x/8YshMgXoy/DgpMFNVx6+jhF0khSPSN3Dm3OVJ/QxeV2TxDwyvVakE
QjzmyV3KcUf6JC6Ad5b++9HRGQFeKJmLSDFimaP9wEhogesYDaSmvTn/Toxi5cXL
Hur+fcled+Mh6BeUi24qLWd26ko/NwEhfQSqArIoZQgaKp1RG9rNqkWZPgt0/Yxy
mU3sxasKCSjtgMpUS2Dbxo1nvK25NXUr4u0fmRxmnFRqaZY9iLRPPrplM0DVhXk/
59AsvrSxKfhgdqmGpfWM4i1YwXpI7RpDOaxz1shSQLsdHdFMdXQCrGe+rmsQa4A5
PUF4I8yr+E0b+Jscu1meHM//wWTrWsI/0sZpmJhhZNlbF5Z3tzB+fwCWk+TgSqVf
oHdjIfHfadZ1tlOWb3XmHwb5oKlHH5lwIt18gdmbrFdwhJRPJcyEky9XAAUhEDrq
hMwm9BKawaj3KXY00qyLSj0GcfoBYHEDd1o9Eiy8ioO3lJ3/Te2OJfVeUNnO0WXN
lO/F/b+iY31McRVCl0FFykUIjry+iKez2gPmWF636ORMSA4zPX5xZiRjUGriZAVU
kxXY7PUDUBxLdsPIQYNcwocnKhw8WLSvKT4H5oXjBymzw5/5YzXL1ATRYj1qQj8d
gSDwGAHloJNLX0i4W+zKd5ngfPyY7+YH03PmLN0Yp9hhPkxu4XFbmU+B6mEg1TXh
s7GWruT0swWJOa4yuK6bcqqI8clHBandhOnWSyASC5WZx4xNN7L7qjPxhrj4eewR
Fu8jCiTM2LpMlte5J0oe2CFZQTr0XQe+TbJO2H1ZIQRfDERL6r5/jnjGdUf5XfsU
/2F3QhbN2aaz7c1ctuuJ17HzKtqF0PoEhhynLPmq6UprFVUsht7tqPJ7B4wz2+by
BZzmpyeZ16GA8tlP7b2EFQfKq+DP4wmyG91x5LNGxERFqON37v3NIQJCdY8Njx8w
jDhtx+8YVpFqdUkNpjUjP+nTuZ9Ffnr1Hg+fXhyY1dxKhUZ4CDZJD9LRpVv1a/HY
HpBwp3Tkw42QmlsAT3ryvOBAUxlGhnYvwLyw8SbrdyUCAl1+Oo38pLLMJIvAxO8O
UHK23uyMtc/NIU+yHqobtYDHg6L0oqFt4BFldiCQBNkhLifwNeIE8ifySQzZB8cX
2fQCfrzcOE5v+1TZTGHVxUofIq4de+Uzw48JO9dx5lfQYRFoOWjE723wHv3k9I4s
n4lrvwP/QNrTNzwyAyQUl3WEkxDrHKMT5ySSXvVtw2V8YkgSaNGvQa4iS1ZQvIiq
0p+oMDxKzgxsdKH7e/EYhJzFQABvwUdprSwsvKHux5bNyMwFFAfcgtD4XpkgW/DV
ufno7f13KU9BMqgnpfHUs3PhYmmcap1f2K452AyFLh3UtM3scSUj3TReo87H9R+y
jGyeFm0KfXdD+El4civ9VuxedwSevggL4xcSI6Q8Ajp28ZKPVo5VY0+FrF3uPQHW
CibKp8dPS6Fljz0h/CtDOiJmRg32rdV+PdBDk/twd1Kxs99edjbS0rFHX7wFVekW
j9J4dDXkEr2c8UnBnbSnwk4tgalczae9J7GT6HPC87L+F2O6NiXqHmRgSY2Yhk5U
X4fnscV9j9CSmYnKhJrEkAUYzu8d58P/CQYjc1OC6pimSxs/MB5AuoGLOZCWt2VS
8Z/x+7kvffEjah9MIX/x6kKBi+06v/IPULCiQ5vzs3prq77fX3f+UEvuYGV5TxhP
rxaPwATx+IiFtiETeUamwb6uwtanG4OKkhTL3aKapsH8ljX5YdICeL6K2cJtDoLZ
iidDuNYwrp1CGLNKVzknrKmGg74pqJfRSDYfZptk/uwP4VYA6o5u7UF355gJz1dw
iS7irBPKaRt/PcUyD2YvaMYFJqKBdNAD4hcniGfZwKqGQaKA5b+n816nr9ElQhPX
rAB6/cekjkA0gO6m71v54rqyUdZ7hwSFepR2fBI415qPJSw7BWz4KWQrFSTOvvkY
/sdQhQ2MMcqxvCBnW+uGIcyLLVeuMMNSnifbSJgjb0953GeR4DmPT9sIN55HLR2r
58vv7TWhLhAl1Ba+66ADQRrUza4rHUx49W2YVb+dQhutm8gkbTn5xwr7FsIyja6f
NB/haPLaODqtzo4BpzE00sZf7vXRXiZOziKEMKEPBCe/mzeGvxrmS69gHjJCcsrx
BKhhqp0PbgEkcbFSFrCM8/7Jz18jZOEnPeWnyqTQwV3izoyD1+rdjmPKJZ5JZs3l
ztee//e+IphsATVmvKH6FkzjOWjpUQw6dnRJhE/fbtbTWLfjiBq1EtY2HUwIFOWs
DIzvJjsLRbiZbaVUYEoU0fnSFkBuGWwzvvP2d0lkzTBJlWshNOrNFKuQA63PvfnN
CywCyYzGdCcsryZ5C8IGic7HkJ+QGLTZ8Pv+znWSnRXACCg/4svOb6Pr2gfkQ/To
wtTAoS1Kd+eYdFUyd+VPU7z6/ifmmZcWHQ32UbR39haBrfD6F+GP5ge7q3MGaz6q
03DHuNFIwLVfgTQ8U8IZSDh6oCTD8dFKPusLYjLXmOR8N4hm6conZ/kCCfpzPfP6
qbH9xo77lGPJ/7E/6g4ZfgzrUQiV7Vlsm5/cmsU7NUrWfRwSRMJ97aikU5ZJEQzK
Sl8w1MFH7z8dWYDxmF7HoioHZh1Q8BHO1MditQqS28LarEh65C5rENQ00OuQX4eH
VW8Qq1ms/8mPCt7Cb8GeK/QFL/bfFc7n2WKCbsFXvWwmrNZx9BY6KP7BqsJYKNqY
19ClMFI5XvA77f5TC1rwd5Pk4jTPe3Ej3vYea7Id/Z0Jrf6kByzztw3YQ+rHcBXp
SqVS+6nRgwHkupeI37W/Ecsdo2H0POYT5jAJpk/ubcVnI0ISfc7AcmS68aRHWqG7
Waz/gZc90nBYel8EOzCxAKoCd01fPIl04ceBAoKCnwRVKZdtx4auXoH3LDu0ciDV
X08YCCQMzGG1NJt51dYSaOKpCLywBeAK9ZwMPPXinIKR8ckYdBMnJksoLXKgY1RU
0GLMqj6LknfOjd5i7pUca4M09ZCWO0qioOLDyEJtiIbsgRjOq58+i1mjB5UyEWfH
Y7nkfiFCQs4j2xwdmiyAi7Dx2Pqyg8Hw2Zv6dTbmQh39op3ErjJM0WVMQTyzBaKW
+yxD3PyNVXDYz1x1I3bsKZGRsQSIMWjg3hSArB82H8lvR3i1to38W5Yv87Qj3ty4
weQ5B2/tSKvZi35yPBOjiJ/HZ5QWD02YtnMN9Y0/A3LhJ8SvegMzzcztLOH8O0Fq
kjV/GavjJEgW4DQbC2mvrKwQb0XJ7VbS1Uiim3KwoKpSHymuBckpd7XPtFKOun31
gqHXWGMPqfWfgrUK4jvl5DPKNOGeNro6JublWHOtlRzLz7Ym98MQTm2ONnoZIv/J
MhVucco7hZrMjQ1wwr/BcLad/VHh3T77ykxLQclJUk3JTvIX/dChuWaDhtMNxjDv
AXuQGhwquhz1BL1xs2AyUCLBqZv+dRsnOe+JxPMpwmbOHrivTD87NLbW8J1Oc4DA
7oVAZOqlM++yLrObOp/ErrBc18HaWFB1vZitMnw0tB2CHgWBvxiUvk6KM8XRkx3K
qLnjD2CvOS+ddpAxcTMAFdh+Pz40Jvfqddy1zMGmikg41C3XxJlMJ3zcTkfAZgv6
vkLTeTf9REoRgdIvG3vx4Vu0ydTYx2ss/ko/88HjEmlNp1bKFt2jbnR2JdByOrdX
6iA0Ezn9kOOT7L4gd8OENq5wkmS1++d8MQdOpXhDuDd2MtPItqeUKxcD5zwmnQpF
vXT2hqsg8PmWiHqfCTw/ByWyqwe+MsZ2cGGEocHzpk7/Ly/mS/7v08iI24qIdS/c
r9rPywWJ7KDZNHB11aSJ/TCEyn3bkptafUpTnbkCDTgHEvcBkX0T9ub79qW/1dte
gDHWEmZ9hrDD9I7e5Avyn5rbbRVFogJy9JPVMEm3TvEnUBU1/Wg+lrN8vHgl+m9X
d6xEPmBTI7BjozGrd27sPBcBs+cOEM/HjSH8Q21MGuq2ihCawBCNUPeu7ldXLruB
tyI9s1iSLQjTqMFKOfqVmwdDaIVgG3mcZQpIP9ZQaN4ktaAASu8DaIiPpZ2rwD1r
yrXcFzLFS0tY0k/GAaXCjGBr457zSi5B8gPWIYT+/NZgAwKqWghWqGkIYcKbFiHI
dIVyXzxrvs/6PC5OIn3F2EDz06Vgew36vWsUG8D7VJ6uGrREB0lCeyntoDKuf3XH
DFO/sU3yO3kgyUgEe/7gxf6p4/GyNXQltmlUHHNAyWsf5nu94+hJ99o/XObk2iF6
1aBrJPWZQtqMMxSzkKoAqbpWVfO0Eod+xIpgpVKVJAXJPhRILGW5Fy6BkELEkvjx
9++v6StUUbpAsHEUa3pL9PrGvLBCBxGv8fYkFp5DOiGNmxm8ZYiUlfpwZEVxEjo5
e5hna5FRBCtMtEui+4gLjA3Ed2/LgYSqmxu6MGqfYj62lxbLnzqpivNuFqtnQRx3
pinap/lHYBIooK021t6cDf+dmuz3e1L3uZSEopPJouEd0mhzzYCXsws29YXAQYzj
iyUs5ca525xf//L8qZ2F1tONpBjamgCvk1hz5oiw9kosJPsB49xbrcoXudknymaA
pZ7TPwoKd2MYdt5/xNHvoJj87MyU9L4SUny0cyHluP6ik3wO9om25uLE1wQcTm+a
T6RFV42EcWNE/ApFgL7B04wIKnqJkyF1hKuWYqQmzxPzicTJ9RRcIXoytN93+z7c
mNCd2rcpsGV0Mkrdv2Rbpf+gpukU3ymhZ6tDGCiLYyaiRGvwmR7HpHujajwsUjAc
AupwsQwKye3AnRui6b9SgXKhVxlJICTMmRh2zaaGJV0OjgI4wrV4tdOZbGR04Nj3
P+2g8i4yBMnSgI6UcEt2waRve14gxXTTm+1R4we/X+UfyfC1lZ3ykFgY0cBgVupv
0mLzxwjlOcKlThX1d8qjv7FvqFhbWvvg3HmRhp7g0ORHNipubTqV2/V/gQRKRML+
vdLj0xFAdgb933BUOfSQPNqQFFXxLtC8U1qrRwxhlFo4ZJpXViSaOPt02jjD5HhL
kAGCpX0dvJGwz9KbAaVZYG3XAqF5fG8GpsWa88+e4izJvG/SWUSghY6oQuFx6743
A17KchziCuwiobBzc3vIQCbWLzGCYIjixThg9cCtqE167CesC4S336Vk6y4gsV8m
5835PimSHdDNgtOF3KmluEXjaJ1mTIYYb146baInpECvp6XJlFnbvAKw3tRgHtsa
U2g2SLW+xHOLWcP0zw7OFdjiI+yY7A4O/9Ux5uL+fe9dfmyF82rUZplG4Z/t8a0T
YKTSzIk1l5TL8UNk0acArRaKmP448/vZ36S3ooImt+3PDHlliwCfDCqfot+dMzVK
Lf5/OKie8PKzffattblTsV3SSTY/dE6np1bEDLJ3l5Qdp6E6LQAAMXpoHl/wlPw7
pLQQUa3BbpbjJciAK9ah38GDwTZy+OqF1lKUZcTAWJI5UT1U0RU1G2HWa0fyk4Gi
FgHi9eFcRtF7WblASKS1y6q+L04oUcgt8q0Q/Kf21PQIaeIu23K4QEdC5FrYH2lj
zQ1HAN99JqSgXCGPzO0dB9rUzClsalkafyq0GRPBxcyCoz8qFeHmCu7ENs6uObdC
YNAnFPGGCT4T9iP0V6vUewnjgFe5QprFqOq4kLRkouF3vtYcphu7GpCBEf/7FwNm
nvKt+yeQ18XF5KICyhI3TnOVk3iXFYLFp+dsmiBHh4dehp87VoAAn2d4SXq1c8Ao
r9673jEUZhn8RBd0rihK2zQC7SQqe3iU7+SnIukx6c+L8uEthuLQqqhlqwXQ1KDk
zdHT98dPjZ+dsZVsDpXQimKMyVksviJM/EEhFsxGo4Hm9QOLRSEUo8B466d7TYyu
vlE1LEWnGwOYkDuaD8OQHgcAsw/TVDWNd7nz8qol57DYTPQFnS7D9YBrwKKj7lPl
FN3dQCaIWt5WUnl7snPVno6ExKC/cbSRPWz5kYdNjxB5Kxo43r/Gm7QlpxJQO5bk
AJpFL3XXi/ZD35RYE/KWTlP8vX8WFR+lsqiQBQyLHA0I7T9Qyefy63ijV8ioPKUj
F0Lzm8/In6ob9LTeYLhsudkqwzj3EivKpNGOH8BuE+epAYIZ7wq6yFQm0kfDjsLy
VSrnihY6tZC/+covYrQbxdYpZoBSlqDVfUSqhQn+woWnmCL7V8hqvdNDsQDQiaDQ
MN9V+kmsiBg7mEcMRhZ8jYnGE0JEPM/dAR+G0s3bGS0hJDtfxRxJrmet+M/7/VBA
qeOXplLLv9gqoyzQAuo4Bz+axiZQpkpLhP99gqeZG/d3/nlTHrab+t1m94HZWnkM
YIKjy82J2tes1xhH9+f7brZKB4DQDT1l/2zXGkDoIhwnfv4etVIo7UfksiRXJbpW
TPl71zIMf/wJHyoN2PFm5ALqW9VXMiXCGlW5w5x+dCJVPogXVc2sDsozgG1Li3S9
mkelV9EIVw73uZ8vDwEWScLbFcGux/NRQ7Q/vNp2MujYiHlYo6kLCHcBIKH0sNcd
C1Xnl0sFPNdlas35yY38V9zj5IKKfKl7zXb5kdonrqzDgG8Mbt99lGJCspaKrKdm
FqYITTpPKp1v1v9HDnadXbhCowntXvG4waoUfJg4H6pTmXhlEVp4Cgqx9QubgwYe
DJywTssr3n+DYx4fFJBGEqIwLEFJOzMEeewZDO7AVUaHmZMXn4mCmBGWXgQe8sOr
JCIsDOKSchOZ3r4v0IoMnc9TMKtMNm8Y+be/XI44LDGLzQ2IZfsETtcDtIssU35z
UMcFyjI/FcAXH/O9uTRTxtNJCSDO5hes2Q2NgWYfoIqPDezl6GI89XIyCyoddCTv
qPX7OqBGgedrztSR6oefPeNZR9ZrJC5Vciaq988Ffemj5xuGo/09OZkFeg8/eqWV
J1aoGgTj6MzVPuqQjKYMdxnNiEBBCqzQ2+ZTIkqgE8P2chQiITvNM4H+oOk6vUGv
1tgWa9GxJtVWOtuc3GgYYrXFHx8C2fmRTqf19KXKtxgbybQTd9AjthDGHPTR7rdz
kg7uJHQJfwkFVipOiX/UazhlY/2KJdrmFxyy54UL+WxQiO6hoqtkhDAj+JIxz27Q
7ZakgHr8UlKEAneQQtMu4aTUvSOfO48fJZeLNUrkR451ULLZX9AjmLT0mmEq5D5u
/bc4x2C2xsnP+7voZkR7MPq2z0bQQm+9Sx5PUb+f9y8kX8a/f1SrHqe0/cPIaalV
Oyua3cFHvwtkw6f+tjWoVvRH74o6qr19GklXCZpx4S3kMHhBfAJuDtB39tF4ItZJ
gBOfShMCPZiM9DSbozVGBeDxiM/q0QqCWibSjJVWdXa/4cJCthtSOVTdNgqa6e/0
BQw+wJkItnq9dPlF1l7CKpxO8FYh0QHW1pLLtqaUhZmzS3rKeMwXK11ZB/FQ7q7A
tmc9HD9bB/6eqwZcr10j5SwK6aGU5Qritw4wOuyXPplv3Gvz09kqLgiNr47bvpKG
LcRKLYFxPJaCqs4m+xAdCyE35PiCHvN2NWYRTQC+kJXVYdSXpxK26Uu8LakkxdcS
oUm2N8+rk5D5IhMNQiRbns9RKFGSbrBPJzeEVzdyo7Z7YZvnlIulGsJAECAE/DV6
tCYsklkhRYbhZaZneqbiIgMybY3ky8qElpmN7/2Uyz48uwFfImuPx6EAt/Xcz/j1
bQNWqL1fIY87Li9XLwHi8QT6lTnu+1LQVgygIq59L+fLMtASfznak1btn2/DOi2B
dXuU78rjo7P5BmgtMlSlL0wihlHDOOJS0au+Yg9LcpgN5WXYFV8j5miY4ou9qfOu
F3BWhTceB2JSCvtYsG//tb6segRINj3Vmy9vHapxEsb08kk+/28gp/oJAYQRn31A
0NxyWxNCAym7iCfec6dl6ltDFImx7UkYPzXF2IH/R2m0G7mChA7ZuP7cyDMa0i6v
SUbpqGpTfVHRV8kL+9w/akFy5YsL7w4XTSfJSo+gzkfnNClHeYjcrMDGn6Nvb7BN
/WYYFSZI60Ue+utPtmECtZd2WeL2FfvlWf16wRRkZrjwho/8COTiVjVhbTA1edjT
vdHtwYUP6xvLcMp1I59+GtBdAFvYJ7aRxoROOcuWuvRpFBh9QvIE/taN40erADYc
/DBdefkleYFV+lCQmRca/pWQjTYsYY0iejBV1lP845Pba4mTYvNZkMgx9WKH+hcQ
Wqw4njF3xlbpwfqGeR2y9cfdpijQQgmP0HQYfstmizz7IWBRNy0RFIScrnZuttq8
uHPJLRsDnR4FeJHc/BkH/1L9ayW6vmeY9u2SVP4HeP4wRaZkZwWWlTlNdRz+F216
AR80x96iuAz5Mcyj45+cqWMcBpby3ZSxym6pQ5//a/hixLdH0UsTBrGQWa+Ya+6Q
oB10bVkr/EuW3EPPFNBwwpmTZRLWg/vM1D2wcM3AvFXyjiMy7Gfa6yTMyZ3f4t83
Mlzw5bL458W7EG+1WTuomXu46/LrYW04e8dHu5dY75Q9IoqknabyH33VZMzwqYAL
8mVvWoSfzbtLNAmFL4iPFcurxBZHaW+ZgIjQsaSnGURA54eZAVUh0E2vAYod63ng
NbQVd2klqF8jlkVn3G4bM8gLQmgOBeF5tdxonudxnWTWINM79S1lLDr2Ru7J1pRz
8NGJCL22TfqPB8M25ODLHD2juSiiUhAvi2P0AxFg1WMzh09rsiMgyHLaZQzJEinB
EpYulyquuu6Yv5wNOhQluOB2027Z17nJx4yP36RK72vxqxiLPRQoQ5IF6OFiJSm1
rAkOZPqierWTdM8xZuCclV/kOAB+AY6VwhJcbcQMPKFUK1Ljm4NDs7OaSSY/Ntp7
g4SQclEVLxSJnOnDiKQH88rQDQT0MX6KR7He/beL6/FiQBEmaTmUnzE3cnmQCEUd
YEWzZbQeA9JW1QtDZ5JUtsdiXwBx6OdYxqJu67zFl1LSDSBHGDft+fq2eurg6j0r
8kjgjE4p2TTweCVs2qSy91njUZ/WlYECOcIvIeYfLSS2Ntfd3IiJtKuzDuF+BOdK
4c5HJ1skgI4fGDyBOWLKSU7FDCP7nyg0Sr3zk7mVcHRb394W5omr4a3ZHjmZmxmP
QyVdzaJ55gGdFuRmROK4g82OLIOzckphmWCVy9Woe14bZGOnuK/NdyMbgTGgZM5O
WxWYaZXCmuELJY5+uNnAVfN9P//fW1GiAp4llOoLmoBYP0fqmfcfoMOok53/mCi5
rtkwH3af0N0kKFnAAOtf8En/V2PZ8J9mmFIFugug8Hqb9K1JGTQPMafZ7z8rM7hq
3wYR/MG6A7Xqkcu0awVisqtfRBXrd97VqpQlKQ3fwhphtp+8JbUe2zIEY859X6jL
pDsrw29AR/PG8zJFZhks9v2oEHfUYFsvesaP/c9Bt0T3nSxf4oqY2s6iAMbXWsI6
W5JUi4A1HH0xbWvnY1xi94vJsjvcqP/RMHSegu45Mu+6EqKlpQ7icQ7iGima9PYm
z+p9WHrfXhQYQF8Jt/GzUICNdnIJivNmRTh5e94I3kEe7jIHlq0bD31T4cyGizPA
mN3fjP1frDVL0b8Bomzv6RwZ2eqzzIGlnVwZukxPOUpLI3CgebtFF0FxQMbxSlyb
w+qDB+4eI9V62zZ+CwWTyNSd8bKE1+q8jK+M6DGapAYOOUN5a/wAH8csdeHS8hkc
0ufEJkI5Y3kFVXf6x2xA+ZMcciNvj1fmBunL+pp8ALZybuRckynJk53Cobg0oeV9
OLFa/kXJ0WiPsEVEWdOLXDvpz9B8cWHoBrQ0xZiSbSME7UxjRAmz6d6TwUCGfWNi
7qd7tSJOQO9ckgqdv2zDQ0hueN2guSBGI/H2sOcMVYjfMQFqV8Y7qwDGsk0Qckzp
JCNs9K1fgqEY9ftmc2+MKo5ZCVzOu+mfnrBcvVU0drxExhKvQ4KPrOExShh+YLeF
I9Yyq7iJaYhoQ8kvpJXdFehzMA0mifcDX0VnwMFS1yUaXKuwhoQhzq1xKQGHC10H
4pySx3jdpYxt3lJp/usF4ZEpSmlwUkYzSYZbRGpzpKsuLXJqBk0mOUtmpv8Q1aDe
0/LG3TK/oB1QuAI9bOJfJOOtZQ0+MRQVgh2bgYxfTxQpJbssYkVG8cAqZXP1o5WJ
Bs7YE1gv4cqPMZ/GN+NTetaFacQayyZVEQaFoutQ4SjznpiNLGCbM3QGfzieaj7a
QDMJ6s3U3OJGyu75gLs96mJdrc9ZPxixdjexYX7MEixmxsEyuSuKimz/+/i+Exoc
BpL9WPK9CCR7UfIth4zzx2isbMOvu3N6kEntZpJnRHvFJsb8apPT0m+Flcwxdc1b
ro9nTUE/i+r7qh/LeVm7OQygeaQuzXY40vmrvWVAzh5Nu9W5MaAmTX4Ckpmx4H0k
DKvfhVY3O3CJ2812aI64jC8oXR74OsAvBOSh3Sl+t0ch8uII/r1nuLrqOq+jHN6D
kvlJS1UcwnxarS2GP+Lcdd862KoWn0JVE86hzzs3Whn0oOtm3uzNpJNv0s9DLb4V
XG40Ufqo7DpSrwzK2t7/K+SJjrh8c6Aop6BmEisMqUhWESxG2nbnEOA8X+kv68L8
Q9h8zZhk9SNTTqtEP1eL96tBy1JRUDkzRyh1Lj4s2breeaQP5s/GoWsTxCmagGDJ
v8eJvLveYAxXKspM8GXJOP+3u01FQl3nI+f8bgZuMann33bQeJevr81S5hTa45Rt
ohzkx8Yw7dJ6r/fr5xpSvGwNaKb1Zh34XsZ2sRtXCLQIvONBjth7Qu98KMjFSbsd
WF5lXRBpQNxPajcA/BzAN+C3IOD1xMEsqYgqFZhkL1QszhpmvGCJSlAOAy9hIV1t
7bsQqjQ0utaGYwAHl/6Pj1G52WM5Gf1cleqSTqnwaTe9Rk7380W8qUw4v7ngnO8g
Gpt6E0A/PrBMo+YEY/4D3A+RNQqw3kL9pLq1AYCuD5gpR6vms5FzabYEV+0nZ9r1
fvgPYxcgnEEVwJ6jspotDo2e6/4kcuvz9BmlWtg3j/MZILwT6DblXyF9zZ4vy2C1
1x7unECz1XDdhdknZTHfbyrs4rx38k+LIJfwpIj/mU+zaTqJUDSEJtTBRsM5YXB0
88Xo2drcTPCbMDTvD2DRMwJN8fXlv10AgDHWF5kw9AqFYCwZlV01yiDR+k8fj6b4
BF8K+Scmuj2j1VazXLxf1Z5oe/xYNb4xmkHs67iknwPXtqPKPjInPGsIAxMh+H83
TR2lOpiB6tpR5ej4C11XphJG4U0bxPfxd8/rQiMdFjoFbWfMW+AyBF7MJjk+i6ZL
SHwtrirgXPDGtN7G9ST4GLZuynqPPR8qd5sWAeHS2ALUSc6N6THMJQw6RdTSrFbh
pm/yzzKMvMq8Kk4IZ3nON2KVsESJDAkcZnHn4fZ7B+cwqVrA/eZIDbFlIKYBjgqB
ru07px7Vq6qwgzqCcQYPGFVMpqg92m3LT2GjefdrEntQ01MgG4Y2Js86VCx4r6fB
l1FggQSxgTT4sK/fhthSX+ug61W/dus/8s142s3yLR/S7FSKlSExmHiV3TeN7Zri
pjCW1JyYIAZSuH+WDLLESVgIZxq8qU9qfwZmNt/DQc5ej879XWw6zdNWH3bvQqUo
T/56jkUxM9DbpfmArUFzv1Qm4KTrwJKFhqSC35F2gEYV5d5YVlfS8uB105jpp/oq
0gUR0pOIwCpPC4zoQWggmpzRYOtnmL6RBvDCq0mv6cUMBhoLQxmUqdpyvL2G+gry
XG0hM3uFPI6h3VUptdWy+W7iqpJVwlXKdcf5iZaJZ4gE7dXADPlUtGdrvAMuduQV
461LWsJluNoKQHYybalV5TsiynND2qUgkM5lK7oZIpewAhcTDrllxv/Nk8nvxEuD
Erd+1nxW+kDJJ9MlpnDeMjGSxxpQyKT5UMjaNPczo/WIAxA6sBkkawlo1hxiNowm
btjDIYBSgpgQMt/2Wfa3B0khfb/t4PdgcMqh7MdznKtA4gAdEMCIBWFApAEKygd8
ei2YKzyyvL3g2dVptZJc8poAU5tjz8ItB0BR/XXV20JIAO5wbg9Rz0lcLAqcmb7q
PznFno3piIUHE6OvMGfrqSytKTG7C9iwPZs0ErLVY1axrrwKR4ue8J+45akJR+5z
6/nh0coxO8FQFlZYrOYAvmjUDTP37LU9CMCaia3Y2gnmOMUwipJZs963O++DOiLK
+DBheLZk9xqjYYXmENW0ficlHtDhNlvGyaBhXpJYFpwyvgj3tyhTD1EI41g+8IOA
reG38+Lnfr1q1l1JjXgdcOPaXKXCs8Yi2KJd75VhCa/yCZ16hYtJjsdrmlx00xOF
RcyRgHxQmtel8fQn9cDopexs6w/7Kwo0A0rHDlrjZY6Icob3fhJtZvkOosRJgpNz
9RUyUN7H3bKFluFRp/uopUd0EWcfKNA0EOZ2GRiVBiWqRl5KdeYZUFQFGRUJEGMQ
tQxK2qwK9F4OHR+bsUB0iiqXfxYwq08gwLur/KSDheNy4tSixAPv5J0ayfrr7Zcp
amJELDI4EJj+Rbyj5I1Ov7tvCeVel3KsJZtXpELQtkdgpic7148LIeXhGCkDfTVJ
VwTNo0uk7yiqh897DpXMGmal0YZI4ScAL50aQCo9I0UfwXUQBu8DfWgk4E71o0Uj
sIr7OcDmD+k+78ng2p+BeSSZetaMONT3W++BrV+YJxq9i6xaD6wwRxKkfsc7g0Qg
RGVAjs/bYqyguvOfJdB/Vcvj42p9ycBhYg2/Emppbwx5pn589fua9wnBFexFe1pA
hag3toydVLeWICecCBFwhvJ5vUdCv7awiAMx2UqyoULkx++/aIwqdS5Gvk9b8zpb
NtokwiUGpJqruHg2i5aFMGMnGx1oCLNDI3Svq7kqr+45PtxvWx5ybwN2hLq9+rxt
uqENZMrWkQuONeq7OrNFvwq7Qz8rzaMApMw1vbBFszT/xY9LYS3s09FWHfp0w2aA
l3Qh3Xica3dX+7HB+TH5/aVwinfAOhO496vQpdH/s9NuVr167yt2X2wth68Jm1sS
Q1EDhQ3e53bZRjkIVvCdlECg741U49WfauXSO9+hbhCK1f21ZXjbDHvPPcvIw/1M
1Fl92nzHEpRInpXXb5ivdonnidXT3Rlbt2yvR4/HTFfqraT/2tmRS/LrpBsCQGoP
EjrsNGeyeiNlgjNzvTs+iPLd5rZDaMP9yjCJUtGTVLCOjGtJe5/NRjTKaSZ2Iswp
oVjXVj+VUBrzAzmxlMOyk1jJDY/iy7n3ANGV6ob3OQI8Q6/NoaQ5XuggCvm2f99s
i2A/TEgzseUHrgcUfedYJxEquG2KOK1BTxxgPhZRgxoLndadZuJ5W8s7Puq4PHXo
mBoo+fteiwx6WnEDPKsLrnRQw4qBSaRILRyqKVYfKh3FoVx6USlnSezJZFtkQL3j
kWLnGICD7GYlBVfQRthVtr5hIxRvIkjafSkgOU0lejgCek3w0MpNJk3innJNc2CS
PlNY6ThQ+cJSKsBZg2eVh6hQhOlOzPxRELJaUw4SBa9fL6eEo48j5T8L8upS/APs
2rqygpVd6VRI/a/tEc9VDin9YSoznnxiGx2L6z72NdMlOoEe+UyFwaVsL1HzWMxG
8+ClMFg70DaSCuUTUk4BBcUbVM6wg9WtoTeN9RAxVGsVLWDoSBKH/UmJQweHdU1x
TtzVAuT5JS4yJs1L17GF3k5whTrkD76hbk8XP7xzR41h7b0VVpYOWWMRu5s9tZkn
dv4GjTB0fDtORofy5Rw5FtKxwisbbN6tSWWBCIuh0Aab7J0xz8EtYiQQ0MLwLwn1
GHvZl9GZEt466VtU9yYK05ZpjtzUkmddekVOjDNIk/ZKTBgg05eBGY4dHdrMzFJ6
RiaVY4aBkEuj0q8gaIK8/QNXvWKF3KRe8qfXJgR1IPGolr/EKOuD+FMxjCMTxJ32
XfUtjuvCO81tcQcblOWdHMt0FRJesJO6MJzanJVWaXl3P0Jh0vTyM5AJSBrOhKFj
OdPMKpFYdyiBK6mZwZur0C1DpeNM+dZfOJQOFNeOhKqLGgsgBdG1NTzb5si82nK8
4twcQx/mXjrOEPGGuauuCLFPTsF3FPfJeBP9CJ9bdG4e+ZHvfPtlyTJfjft99f3m
jQir+M1zq37ek8K7LQu/9BUVaLA2nojvzh5KmYqjcmW7Ttv8ZEGKejTSEiqpXbAj
22WviCQx7RphodNq6JWGja3Q/YQM335qnbI7kWm9Zs063nh6KIWQ/y2daDtqbrwl
znYgh3rlC65yJhrZnfV3ipNaqzlo6XaE5cavVMIvYj9Nt98KEaqV53LPSYitH8bB
ApsyfLgT+cKOeo1XXVln85wloxolfgnQKZaF9PdZTtxZjMY3lvl4Xl4hH6x8vRTC
ILXuTouUzjEzqhO9whtkjtDn7mZMKCDB/R1ppMmrrbl+irhpDi6vxJ7ATPQ4BqmX
YNFGjXNNrljRfWciM8QySD8tQ6q4DaIDgqnxqiXyrpckJ96J67SHvnrfew/1JfAa
/XWY5zlQ30GwwBwR01gDWwhVyy1CMYy5BwSfNzb/PDnEoQxsmsM+1AajqPSFmQul
75otF4Merb5U/1mqACfA9NiXfgfXXu0HcXdnizhcrj6NbWvumPXNGiZdav9rCauY
ly8/VV4P6W2ZmezzMMGEq2oljVST9JcFRvhDCW456clYeDv0OojxmjoY5ybOlu6D
/9rgaOA0kn+8KLrboNVJcsCIxV1oOXqdALpvExHWTMqdoxeeXqXr2QStTby1zo9A
rSXfEB7jli0mfriN4s1teurvA6dHm7rEm6D+Fd+K9oDWjvyMk+jGgPogerHi1ony
kMtFkod7j5MvTBcZx37uBxObjev2g4e06R7ftHBJJVKOTiTT1DWcVOyezE9Uf7Kr
AR6FLFePjkczLDse0HrHF+upeO392O8WqYv8mv2sTjz4MfaP/RCldnQZXEmgcr+K
ynmvd5lEQysgWeB1Y/L04QQOAi9MfLdiU86G4040AsDhwoAO3BugO317Jx/Wdpls
ytoWodiIjs1cgvwB2boII5mFVH8VthRfpZCMaYkEbJaEHDIwFZ9BWS0AWTn1Uhwt
wLsTrPrb31CEI+XGyNcDipdIXf9uW6Uzcxty6rpMh04WPMuQSZlBy8gG0LK/O5Fn
hdCToZmW6yA1kK/ZmzwKLl+RqrFvn45wcuQceN+ZLxbex85RI8gR9N9YCsum6V4K
B95UHL4gbQWgAEhUivYZ1evK1gLP7KJweA2hu48v8ffsCGefBIKHYTfHWk5g+pV6
MZ80qIgZR/YvadiHqCZvR6K1eA7IW5FOsHSpJpL6bdmptKD1R2UeoJn8smUOXLlA
eXj4eSdIe0XhEuEfx9EViuNXRh/KqdzyVoRBAztgxvRFWH36auZcK0KWn2HRfBv9
2XrxYCUWJttECRtpv2GdI/aX/F7L1ydbcB4rE9D4tiY9vGV6hi5hbN/XaOray+2B
ckQbv61S0sk6eArlRWJSbsj5KaCheRpWwltHy53RMhMio6PcXeqqeddSEqe8qQzk
PNIJajEySuX4pbYx9l06NmqufZH249vrfpdPXZ+z/cctLuUQmG4aOTkgeNgZXusr
6r16WZdIMLv9NSq//o2XYL0wobbWXKfDcFQU7DI30SFDG/wurwaJT6BZn0nldQP4
u36Knr+VCYt3L3nAnXbU7Mh5YXIHOlRP4qKjdejniKe6ffC+wTntd+H0IHK0yHTj
2PJB5ft7Vq44l7s9bcrlRmBze+S1HnJAWriseuHHUl0oWZD6oqs/Rapddjkogcul
G26x8WZGZavHHiQGxaaelKlC+20F4XKGoWm7b5y6vB2tT7EOi5x+mqtkE7lA98wB
zVxL32lVZMZNyGYP+RiokNDRKO6f9wyD/cnbtYt22eVU0xTKlqcdByV9VTv5VmWF
9G6QsmgrbxRZduEkvEyHcb4ZN/jG8qqjTbX8d5HKbd4QHr49j/RtNg6Zq9w8RoNN
PTqpK+c1o11h2IV7ZdTtqudBbPhshpNNxldNFfz4lSj3e3/7btPVIyrroeyPY47G
DhxPqm/lpKfQiCt4jJUx7eo2yZ3a+nwKf2/isrTLIxInEsvryaUyb0RXOUWshWbH
ORywjiWAKC9HjugFYGkbWeE6iZaPftFPmkZPAXfr+1IRLz87kHknh40mSHFKaWiZ
1Mfy3nY7SK21FxVWxP3Bhft5Aq5uwIdEhk/9xmrIFVN1y+mc6D7kVTmdIovUdOo8
vL0Wsa0mdT+KF0v7onZxNhc4UOjwsrPR/GFTJRvx/7HfinvhK/IloRphXYmn4g+6
Le0+WuZIZjjwIB2RsySAsT99JdheUmUKX3fgVXJNub7UMKWZeUzVFW0qNfrUTV5U
VipQcjoLaldHUOm3ygeobS+GWGZzZSUyeAxUAyh/Z0I34eZ7wzELOPki3PtcNEAg
8NMbkSB7xjP1Q7XGMeZjbuOO8tRRkOUrWoQ1hBrLjns9jfWM6PWcbvT3hbNkvnw6
ceI6PosbHLB3K/U90ipnJEir4vnWrJA2zGvMupvw5xDT549dEqG7dJqXSXzQ8YWQ
S9HdMdRy4QIVqIhknz4zMRb21SvQkcWKGt0fSTI6lsevzIUDkibJied9C0sdhXaX
De0kB0Qry/gPI5FFl97OlV5S7Q9hA05Z+FCuJYSyye4nxF4Yu/dY2BdLvwaGF2+Y
pGdb/5ssdWDX5u8OwPPf+tSKwEcXgteN5EcGfWLr/fBoZEo76qfLhOR9UQimwCCf
Ys6JK2rBAhWTLFe5eBAe0Q2eOKIksX/07zb1HoIR2fV4bz+jjGaL/DKuroZI0YaI
utz31APqBdEVDAR4e9uXvdo5DDbkBmy5dFrtWqnF70gLzPtBCmAVzzZzv3xu2F/b
BbRrtoypC39BZTBueuRTghGKKLmHmrcRl8RDLpM5e617SV5zXTeouD57AAIrAxjy
Z86rtZ8DMwBGAnkPxe45Sr5J8kVu3ygHETgID1xx9K+mQTQelSr69S2at2XHWBXn
dALA6XelxN1QV/kVR13G8A5YSlGF1GTTswKf71qKgd/6DlrI3vBOTRrnxAqcoye8
F0RrNq0kwAPej8g88+fri25BQ3ab5nNbbaBK6trlw6dEvx/vWxDfEyowJtFv3XWf
gO5UXqYxaPdZERic4crgisWejNpyv6bIuy+wh+Q/MCGnk9+J/DjnNw/4AumtLYLl
+9iem0poScmLBMq7te1GU59x7InCuWCyKiqrCtKWXXe7wSgli0G31ouTaQxtgT6E
X7rAOp6d+SFnZqoA15o/xt+i5KIrLSya7atp7vxC5URWxOMcCTSRk097bRf1sB5g
iMwQLLo77xoX1EJq/E7RdLLLwQuFq6sUNhReJB2t30x/KViGo8EdAlAhRJWWmdLE
6DDrUoElRNgM+PUIjKtstUag3zHUkb/oZW2Z/olmR7BZM5TDAGPWdWgXQ37ySXbZ
HELFsueZQQ4yWCTFVtikyGVwgJPjkpKRqtgmgY/4njFUWSR9adN+DJXCVExklvAR
cbu1gmZzchXVYUD4NSfnErNL+LutEU9TlmWVHv1iggU4N7s2YBDywL1CUuOihWYz
emgxKpv5A8OO5matk+YdtUmoQvFlwuxyV+JclLuv4rXlPvon8CqpHnPSH2nlwi6e
AbCMZ4THXU+MShbZNfp1ZvVP7A1J63XyGs4fSNUs68m93HidKttOrvZRGyjY/bUU
xy7WyZLKugNPO+dQO3kfu1rTZiTVwb3s74CZHkt4/X4hv4SYZhF4rDWlv5582wuM
7oVq76gBHICBJ+dv3DsWrvhI8Ze7o8a12/Bu3XwVW01yGcCXcOY4qvYzSPBGGKmS
OMLgx3fukazYN32pQ2dHAFmI8LtANoKen7z0Oel/ms7Hw8fFO5XLrC7JGWOYR7lH
U6UnjQofGJhz0S5vzrpBZPBtBuCuik+9cR379dl6vDqSWm5lpE2kvChPhoTss/Ro
nMq3Cl9bn7bBnNvrBOObRCl+hIlZJ9duawfyE4BiOQfd0Xsm5AM4AMl5l0XfNNm9
hXpDqt1uVQqx199FMIaG4qn9siuM1uMlt1SwD2i+GhZ3EGsAPIXdrg2SHKkVvI/j
Cxw8MnG1S8W4+mZ0GE1IH9npfbvFzPBC+xj/h4Rl+OccjeQKctvj7BRiWcKoz5UD
2FTLwOvY9OJc+Yi2+rxIORbAliOeD2kEHGQfezdGcVRW/JAQ+zi/4Aeh5FSCNE6g
U/0VO2ZsrFncdUm5YhTeIBvepOJ5M17rktuRMld35eebEGty6AjrxlES3BT9adWM
J9DuoZ2wcGWhs8THBIys+q2xLDIbLgEmy5dvO/FJx8lyLv0e5NbhA5ie9jLnJpmb
8V6CPDUucK7rZoPFp38QPtBhvLvLLSd4MJdPWJ0DcSVZh32DFO+U/uYz9Oj/jIaJ
CibCXHMv1UQzsSSEilY874rdOIExn+s8kK1TQ1tmiIMot1ZsJZBwCnI1MMTqyoAJ
AhGTKZUJ9Aiay4qnGj20W8jkXlG6Q7Tvp8XvS7GFPA3VYCuMXDPPrz0j6A4io15p
2bgv1Esg3Catpl2eUTzOBuje9v8RaYAGKVkofsZsjoVw/VukiiSSHUorcyiwrvYe
cNdLtK5shGdqt7qwK3Xo7DS7++vn6nxmHQyqvD6YQPY0RzrEneIYtJf/s75k+6Mm
u/z0dtMAANRgO7wpDMzQ3yXx0myURa2cdUY7JWxLbsNx/5wFJuEeAgIkuL/zKHPW
wi55d9/2T7/NlkAxQfuJMvnzflY/va19sIGjWCsMwGrLUaHkMp06GtXztX+3DBxf
2S3ttlKJP/Zxi5Me+PsSMtYJTEr15zKfbkr0U4KZx3qydgTWVGnkgUkblc7UPcEC
KsF7Nb+FxWKhEkDySrJj1QWrxfKwfqrzWL/nNS0fF+e72OXfEhFj7kH9Uc25Rror
mIlSANYVjJ6J/JAFT9OVEI8OgzGe1u7u57A8eenYrW35vgQptDmp3gRp9pSSFDgR
eWzf2ioFaEN9YZQ3qrQGpYk+m6CSdqPde8sBoDwePaWLgB2PBUjpkk6rhA/7Nd2n
9RyXimpeFZxqF3CCSw0Io+XVJdeNoDX175TnPASBaxpgrBKmDo7/ERB2dZyRg0ls
knNVcIyDuYY44GOkHgHR3WZvIiX2xs5mEsrsYfzc3rAeMk23L0DWfhncs6GS0cCh
Mos071gWcGjy3xwbCLx/79zstRSyPCon20bWU0+fPqqMoGi3XpHqzNXja0wEztoM
tKJEQ/3s7oE8ZYPvCC70wtOJTi1CzgJ+khGSdzXN9l9/6nUmHsazyoQcqqGA5pso
ZuwNQuqw4jrw4+Tqa4UHVa28L80OuCSU+T1o78RvuML9U5VLP7PvSqHxPImVI0lK
sGfVOTyBdcKsOtcPi7LqT0w7iGR7IQsC16T38NNQZ+cLanp7GtFfsT7HzaWTEl49
y0tLKh4n8fIwSMK2slrZ5k+DqoAr5Uy6Ck0efmiTCo0lHxR8ZXlSdEo+EASHVhqZ
9kcaqzzmNiLTB3D/05ZcLVeRjmrrXAveimNr7CQqe5Xqahfi7h7lShUdReVE3eY2
MmQAdsTrmBtH+PyEZGG5xJrHpTp3ZuVQVDQF5CRptsHNKr+77EOduMBzYVLI6L0s
3Ji7yzOHyaC4K8yFz8iXcZWyjFieaGIHbIixTFJqf7BUpGTWwJ4r7yFBCzGKwf4E
p8sLHLPklf1FA0+bZJw/yyuC7L2ouZOsRa4bOJYwFLP146rRSE+UI9GfR01nqESw
CyR8r+Io10vRNHPqBhXxQF5W6jLYrtwrEsiryEu0ipqbRj0KDKHwMFOFgXNaGwSE
5ZCquF76QDwZCFuECJAmgYay2DOKhp/lNSZPM33CJahbZjUV/KSf4+FvomO7DZfs
0hcpMHsq6HyD0/ot9zmvkP/1cvIqik7+ygBbgPP+5qTIUzeY6JOc9ERhCXQJxRs9
EQX1idvH2/kLnEp6/3NqXkb20MIAPT8QXlqa3R3EVi1gjf+StNuaRjxWukgreUYK
mIBHBji3ntHYRcoxZSK9IYnfWNtybU4tH9t7jGodpHiMjJDhB01Q/qdrBgG2ESGX
8ss10fITpw79y//yrWwIr58HagtIG6FcsiYtm4C83V9u0oDbK3AGKU08JkHVDXt0
HD9hFNL1GHQtLK8Vn6ffW7EIRKtmwC207gdGYJadoQvMEvZYg0nlZBIDo+dRc/3+
7qZukAPJYUzDZnF6V2WT/VMtCcHNaia1w/33m/pRKl6NHlZ486FqJWSa6Yk55MEf
plJz7f4I63iJcTgnOaiCwiafTvCAbxh1nmcNbSAMpRx3VpaZmI68yaOGY6ehc+XF
7J02u1FMz7oOcZD0poiiFjZuwF+q9supfxxi3tctMc8YXX7sCxqLXS31hKcx+yd5
OnoEt3ROcDSV7sibLKkxLwZ7Wv9B2xBMqGqlQ4cH8X0AP2rzJWFgi1gWs2vrFpYC
oL2cbFzmmJgkwR6Lz1Hjp/IY+dxKR8SeiDV94AByM4GtBnyuP/OoFGz4T7HwI0uy
nC5BWeOW0cr83Y1GTgQLY1A0JgX/7BvYu+cACy90nh8rA+SJ2pHQdB9kLs1bib9e
2HGWnHXl95C8Ml/bn31wjbwhkz5nr/x9dIA8kouM5nzn7y7EhSBz6V+smJqKa3hy
AwyZvfJxQ3YQN6PJprO+U7gPNbWFukUKpqf/qDuS2IU7VlVlk/mL/r2HmbzXRwRt
slPsmevuz5un8a3XIpA9x6TMIrbuOerYwjbbukxfQpv9Lm6A662wZbSx5TYU2owx
XPp0d5KsUYqE7RFqlBpFQlKkCs8t3uFyRxBRc6s3eVx2T5Qw3eA0XmGFYKyINAsb
tXKpzVzDQYBeWVwX13a7bbHC2Dn7aP9bWcwnIfKzxouy76AHNG13JjVdL8EEu3IJ
ORShDB1GTzsaUFwXdBL0NPMR+ll1QFVtGszcJnE5zC++Jf2NA8Ym1fjpJIVHlZLk
rOJyXwb3mDGR+dhIPk2ZdC1YUDxdzA3Qqey058q5sJT9lk7S/dZNFUcAZ95T4ENI
1z1yJXTawAhUyq5n1NsnQRWZBrl8gKJYDInMKeovl+iAK/HFi6evmM39lynPkAOM
yRHaX0OJY5Kh2suOVt1EcFVCdDdyYnbOrWhI6Mo8a2aPda+m/7qiHplkaDNjP7HF
NljrnyHGOv9mqkju1W4s6ZdX981IyTj1l54ofcNCK/jAppOMxeZDPNe/HV2UxH6y
NIMKQtHB1w5RqIgyy8NMkdf2NX0qGnhdT9rC2oCyF3wBqsRNGCPrUeDTTxrO8lLU
mPPp5MvxyTqErsFdPrxJ1LMajR0yEYbYx51c2UOEa38b/a0kVR/CTLoAwupeL9zF
Z/Vo+bLJlXSjBjveD8B4oXRX8bHTCOXhIEYIHIcRpPFbrzgDKWq2/2On7K9Yu9Db
APkMQHpcQfC5X8syB2Jm8FY6ISnJe/h6UQqM06LJSTQE1ARK0JMvtcyrwqMBgP/1
0bEZ8BWnoqXhV+j/m9aZBorkife3XSBLSMF4dpShWqFOFSdiN3kzpCOZ9651yCKo
zOtV1FvEDQWsxCGa0j95XdfCipjD1qvHpK/XbM1ST2wSXhXS5YtIom7n21XxKmD3
+6+e5nBgE2L8Gr5zPJt0t1HPZ2JvglCOh7iDOTM8NYRSCIs6mLz/Qy0JOxxrwz3H
YCo9Knd9CUW+C6FP8dgPqrYBqaCnk77swZbubSJUuZQFLVTQwbvYxEYBxHYADj0R
Y8s86vV3PiAZaGzvLQcchEksf3DBVnTfiSPA5UQQnkf8YumDPANUjVZHnz9U0CrV
fqk8TZvTC0TuNY/lhNBnNznfUW+EV2Eq4BjDPbyVnTXMHP/3CQrRpuwyWnrDTW9R
BCWBFXhtCowKSlz3UA/0QaI+RIpA4Dr/rmGnHHSfRz97pMhHCLg+6vWMRT8XgUtd
ykGAa50KOJ5mY2MryydvQSb7pjszklc2a45wX7FlvibINFRELsHsTp6CFcp1/xNQ
uk1urDKE29iN3rnDLF3nVhpRZtWdByMZphbNRaMgXAox2AUUA0BTFI/hxXV/5cm4
kbjfojRhJTpNHWGLHpLeqjnzBNL8MVI3Iv/JJgkwQYWI1Zmzg6vQYXLDoyEIPRH1
pvhm+SVhjvj7dJ6OfVtiNVfMTRPl5npsNHQ+TqW+NVVIXBSgbm3U20Gwr34NSG4f
5M2ZgaJMpKjaCELve47hbzKYHEvS0Ve5L8HNZnxqPXvDGsm8B4CTNLDSMX1YFVNI
Au5gRX2ozGtSRrd9MiGLIHOeRuSJaTeVgVlhCzZruMVAHN+Kr1QFcZSr/cp/t4qH
PZUACAJYeHsWkg7bel3JfPpO1t+xpX59MoY570/Fdob46a8Ts7a57oMw+ANPN4xu
oKW5ciCIPs9DpEkNbeZXQuJs/AvFA7AkEbQfCXABwD0LWtCbUSASfyeFUi+NbxTN
YXHWavWLtneIbtlCBBEIO926tMbSC+muc2viv1nQsVIdSHHPHn+FFvLjQNbDpsDn
jkU7UR4lv8TUvw6Ek9J3bA6HviV2nZ8vzlRp0pd70/4Ag3TuoyAEL2Sj7li34xzZ
V1IdXiWDvjxh/q+iIp3rGd2J0XZ480KfXsihpRpFRRxBPIZG3hwQoCDBzMvm6m4X
s0G249ftzL6yGLzYCBniUeIhdhX3Tqos1TvadD2d6z3/YleEFy7ov1qfq1f+4M9U
jrM0ZbOnyZqlkpz4egRl5BHko5Z3go4+rq35I2eBZ2+eSFLWvTisVDvZuyIqMyqh
4hlYxujkH388jJguUL7T3AN5wzGiuv7I15tZDzEE4U9Ke/8HYEdC3cWJWJCbxLe2
OhRKkOxK/QK6P58pQuLyzCygG4Nu6vWlxZhxoBFlys+1/xmLFpdcxbtyJDOzHwCH
CBb1us8ipWlOu32Is+K0PlaGyxHBo5bbq87OV3iosz8TBlTlkHkHgnArlpn5Y0ib
ebqnULYlDqst+L86ja9Nwqn5YovRRqxxOgXzhggqTG7Cm7R3N6AwD3Nwiw9wDTO9
b8XASAwEvn5M/BAZ6Sp8gBD0PdJ1b2dw3JDQNCgsv08aTekvUlPhCN0KxVaQ3tqK
ackh+xzq/CvU3reKzi3Onpi9JioiYdbZrJMqOrAdRqFcIgUzrnfyFJAf1yGzJju9
m2YeB5wWToZoyN7WjRehbwkh5CbeT9/A4GkUDB1pgGWbjKrGSoo+u8sT6Kd9+rOh
Ruy5qvYTVUth2nDZP7At2VVx5GTME1fl7WHcJPz4naq2QLJmxrkRFHS5nE5pFVax
2Rtthj93SE2uEyaqsWwhXeeGNG4t0lTkSGXdndLgC3mtduxaEZEiNmTyUnkWO4RU
P6PHeZcUHmf0vHyHvrlr5mRYGJR2yeOZvgoITdQNUSoZ3vExctDt+n0HvUAyMWlD
MIhT4bRc23N1x8dKQIkqXECBpCT8d5oEwjf3Z5k+NHKqHMdorJaU/qf80LpW51I3
Sl6WsD5rdKEDGU2TqvOsFlmzAm8rJ8c7F4Dxd7XqwB1QzcMom5P0ZPGD61NX5Qrf
pJJrl4nL/VsdIEI3ysVhEl4TGXbkNZEyUAUXI2qxHSJHBTUbixYHNSmG1SbxLMe6
Os1JaUJnnGII653rqKmGpFrSXeRAvt+DkOH8B1u8YlCjMcEO/VJy8iA3+yLkqax+
Uj51wBDXQh76j/eR311HZLldFM8VpL43/Ux0ZF6xsPZ9p/2vlC3bDfNcrf6ChOXe
dC7MIIm3H50NKKZqGpZ6Rt2Eoxq1mwDhonjymOU5JiOGj2Jz5zqiNt2ZvYNHwXoB
OJmcpf9OHaXRlyVtIpLN4CFeIAokes6tEaYPv9/uUQILl72kP5C0JFMWauJ7Ja98
GziVoBvzZDO0lXxcP1U5pryGrMfsWQtYFOV5aJLY8lknJ+Kp6kHW96up0nejo7uF
laMdkd8zgEBCvnmyP5elro1FRrjog8ftuSGxskyoSUKd7R71USiPcWPcZbvPgs3m
Ubx3Nhf1fVMpquErVXIEDF9GITzZ8usyvGKUQVU2/8uXK/EfhdOfzGM23zNWTl+t
Q9lRK0JQgfsdknBTV5RWsLga/WX4SMmNZhN00SwbykQRQwZ/equ35WSxOX7JYsfj
l/stGPW1/69GN3NiKGMa9gX0c/Tdc48MuJZ+UlumA924TtfExIUICIYHX+tC/8Fv
uMyc8nlICOzL/11/7AyLfQynNmZ0hrhXXshFRMp9JyW5sz23jfFUM6w/I1+XLYIy
nF58IyUiOedFDF3qfr9wSTqZKIlBpidSzIIMtfmUZwEvgMiTUF/L01WeuUVXkw+v
9j+ybbpw5G/K7savBMYHw39OhXeLKpOPJ5WU6O4JefbeZZNFCWYmfo+mZuFSP27M
4haMwtFFUllrjCXyxcF8HyLjeVsvTYm+N4znhqe8O7C2MQFswcNIdd1lq9XAOqS1
IIRZ3S3alJ+endIxKrJCWHwUDmUQbGqQJC45le3YyKBotq9akQVHcbkxiinmHw0A
EaISfURQP3CPq5SSL2/j1XJXjGUvC2TysgrZmgTw6gRcl766tKG5mQgBfI9SfoiS
XZiJhOXEynpTgcL/aIyQagOaxBjSkYSaUbB1DnOou9yLuX2KHRra4q1kAqmcewZJ
5san+zO85usTTlyGJgsyNqlzmUHbErD1IxyM7xED8Tg6FaIH/3aXYc9wTHgvY8ZV
y40FEvA7ZML3+i4U9l06yAh/fFmOSSH56QXmw1mLKSwAM03fFDZHeaNxb7Wd+U4Y
9u+/EjJEpjZAuFBpgm/YKEt849fnXEwFHlHFP/Wkl5gWkWOexRbD43dbeClMGzVn
eAKbwr0Vt7UjZw8IbMbIgO2sUSjwXcdSMYAKqibpb27VfgJD9sSKWnJ7b/RTfuGP
toIiA7oeEytP7qZW4Qmhs+Lhl+e/AelUlZhVW76/U9po+m+ckaA5Xgi7GXFmJfnz
y4f8gOE3aiEiJDFehwFMxpSl09pQA57tgbFSoS2KBv7dgXMTJ5DGRSaFT5UXX95r
lSZgQsA5g0D6t0Kfc8s9xH3CWmWXUahI5g3pLwMiUlZCtloYJW0nSxmgShZGy+AC
KhlPkKi0M1AtfNEh8/nH02HiZ/+rjaY1YmeTPoYcnnRDzhqIKT0Z7GD4xTDUKKOm
GqlLF1Q9qnQKbooOvRworfH9RDyq786sP5JeRftvJKIoqsiNlJDYZsdtihGIgzi/
ri09TvVDbsoS+bzWa7Do/0ujeh0SyP/nd5t/EET2TkcsP5R3TL5o1oz+xiYyFikJ
KLhdJ9ygk2CsXqw5X5AKMt+9ZsdnHzt/qWDBuqIg2OWlRcbZYb3Vz6hJDYljBF/F
hMR/UI9+GRkHiDsg5M3HQa2zr2gWFRH7jE/TIvYaizahGWogobEdyRIKIKWB+Zg/
CFcu8SgmPCqXVZYDWz7ETuYl3qHvLhlsti84BAiJ26GqdZqxdmcCQqB+sLvHxHFB
L3V7KsvXVnK3ZTEio1l4epdCborCXDFah+P9bTvr3ve9zLan6OXuNZXXy2QxALbl
f9zPl+5lfG8rxq3rOiVurgcG/q1+UlcMbB4d3L441YkbVN76kvdefvKAFUTHswk1
LUzd9QqgSJ0SK7Z5lMhCXDQlyM0f8UhMiN3zqLjUlPwUUqBKsv7OzIaoAj8o9fDR
8b/6K3qSNacmKDRI6oVrT05WG7laZgsVOL9NJLGUdSVFzNzhdNAyfoGCUiHLfxHo
0HnbOUK9OrRHyr1angXtRxv35wgSnRHBiBBuvunc7E3tGXb6E5vPCMg8sj9ZfW0K
LAI8J9ldpDsmRCmutCFsdsA7+5JlkSQ1hRCeyMFdDVm5wkX0/1Jcxfr5M4Uc8QKd
0xKjh2fZXWQg+M6uBDZ7O/7r2jlh6iMgAK9GKsfSF87CKCk5UO2e2p0OjB2hQc3p
`protect end_protected