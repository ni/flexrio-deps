`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11328 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhNy6VWIb/c231w6GZGaUgwhUZXi7j8zUEO1Z7E9J3zs+
n5pb+7+qRdKaLN9hjD4guFRFg+no5bkBYlHATkQA/fp24EelXluh8psnF6ekBxtx
Ek0yCIlq1rzLmlDK7vfgVl1YeExulRE5vh+T+KJ3vBHFx6XtfnsMGOVXokqffOKC
SHwkUSqitTjoV0x76ZsTau5yepw0CHH+MZZwSk+uYNcUhrbzK9S2k3Ju3m8NERRr
uFC2Qz8V3c0y2PaqkrNA+QU1qO6hhX/B4x7J+aBsZXG4avJVTG6fFx1Dx20MW85q
Wj6rUTUZvVzcS/ZfvPMnjjeBdnqRos6MuYIx4v4NrY/Lt73xqUIWXfElBfL18aa6
KdImwWv3wHiaU47/1tsM+/CZbu54iTuU2fZLqQVGdYWryHssDAz3U5RJwe6+NBew
SQiSrR7URD2hdmDTeWo8kGGYe7vtbg1eJCbX7+Muyjf2v2G01BKpp8Uzn+xsosvs
KgqSzm02ZOOQ2C6AgaiDt+4EeZY7JrJWrVjJN2kBplZJV+wv+eEJV5Eb6LEmXsMw
IwL1+IUB+I4+9+zHqMAzCnHReHV6uYUNlQX5FMjPxQm2QBmSCgmLdt9ay6CdlUj5
2a5rP/Rzy6BQsfpRgPwU27lFOMgwjGkebUkOZOuIAeAJtYtQDZEv2lGBPhBBowL9
kYQw1VvVrk+MKhOKsYz+QZLG8ik3gebxHgwk5e9PWBPTlT4Dw6hryvhoNde+iBlo
Y53KdRwtlZnQr+imwm4bwx1LST5CK2qejOzh/x98xNEgF7+ddGfbaZ0YbKro1SMA
3EMGKUruWsskYMMr6c2ZZjv+IH9OSe2fPVdPYfHm1yeX2hN4qn6DfJbHAXB7TDa7
/LQ2oEIk2ezfkoj2aHBJRme77UfMgnoRhSb+sCvh/1q6oucaO47H2BAbVHbzPOyI
egucxNsdxgSDSusEj+dVOmux1bhBKjrqZU0fs+lMavo2u0VHvj7yCeMu9VEdCVNG
gAlIICBRO8XsOmpR32S52+IOZMvnbkI3DX6yC+KgpL18byUz7SfzL8bD6d3TtiQh
4yK3P34PHDHxweY2cljnmGZFNUOcqQitcks744CjX+L6tr0yiDjU+RI+xLk5t7mW
gY93Tn8userPhztXlOPY/gzqXy/XkFEYbrSW7XAfigvHL3wgAIdcCXDTJ2cfyPgl
km9NNwxxtOwjSwyV4raM6ABce4eh5YTa9qHc4khnGMESKP9HujRDlztZLc3mR2kj
oiH/aAYhCWxxEmAPH7IO4/TuKDcFow9nqxLLvcPKsZ+WK+f2OXhesSyaq9ifenPl
+BU74AQh1JQMXYKDGvocdk2Lw/9BNsnlfwNO19qL6PP4kqn1SIaskTH3ht87qvGh
5GCM3EVfjhGl5xOxtSUcaOZPQe+kcO9m7QJpiwPoSp5NiGhCaFL8aq0P23DU12j/
A/EjA1JYvkSUWGN2rGf8Tdf304eTNIpX9dF78ANnOLgD3kOLEsHqquDT8/fOoXo0
Wd9rxHpD0D2qupURod21SzlRswgfNJBFbnj+nWIIvNt/ErMeELIcQNT3JExh1L3z
PmMtRwYXVAbJK23gTUaCqdPcEmzsxiOGwYE+MUa/pLUdU2QiTOc8AYSnApAhvWgY
lSiHS6sJflBdJdDgL6C8zru7QTbcHdRX7ofTtLx+GrZJ/9QvvnfgKraY0k+IRnLM
6WOwT4ioMx9nN8fEvBmqwuO1TlKy6jmicqEWZ1q7RcW8i4xlOBBQRbZcOSUQ2m6c
T0HQL77/f8duAaHOkdCrhago4/0RXEn22F146Z67XwdF2WuFUgOh7NRMm5fvyXdX
N/RwBL3Qlo/3hxdjgOoQh3UozXPyL1GwTQdytbTbwt6TkIt1IocuznFIYa174aoq
llapI/dJ2hfn1RaOq2qfrsc/Vpu+4P20HXgttFJg0wDicwnxlhKw1fedWYWAdR67
0OIFQ99U1UQnJTU36xkIYHdVivZv9DHz32ML72M7vp7mTLbTmnwI6bN7kWGalt8/
rTYafTIZBhPj1NOrwyAONjeBds3fqsPz4ynDa30sYSOoipga6CCR9zCCUgkczh1a
WKZfKHfnNlJmzPELXpycvObOh0B8FJE9U3/xF8meP1sgiM2rw20veOR+8vRv0IxC
0XT23N4r3QOhUPS8WYwreJAZnhR4OyXVnhzC75UZ/y5EQKAQXk+qfV6usNvTFQRP
2ANzHcKWjmMUITeYIOK5toekVxPUFuT/+KHGmszvVUigwS92tvNZlcTXNfxGVDH/
NjLYvcb//Q/0FpUiMxeAxqf3fJiRDitU7upJsyHWqjSCFLT9hOoc8q4xk9f2AeVr
rJEgA/xApylwZJLX783DuhRtMdbzhe3a11Zfi17QJu0dbYGyYsTx+2GwBoMl6sph
TxMagB+oWQCoOFqTqQIn/1aoWCPlnhwBmxXPKz3QdoDHiHlbIIXSYZCNsm4DjL/6
Xees/ToYVZ1JsvmVVR2yt9utS4rJFXoDjVhK3IRWpFJWiOagAIVLXjYWPfAwb/Ge
LGuSHBt5UzHane+WTCcKCl5KReitYwdCc+1VqUzPdTcjD2cBLJW4sGQLKSPGL4+6
Aphf+q4xWeqp7V2ZACDxEIeYgWqUWQTOxNrw11p5oVops0rsK/6xwRbeYRVoXu7H
wc3XA4kHHM7JwVqLdVf7/iZFKTQx02GGYwUWKHn9ibw9f3wJdzPqyPQdUBjvCJLD
QDXOe4r1nMuL6nmTAZ3oIJI+rU4/StboahD9H0YB5iqjqBu8PJPl+NZHCSMJmiHL
dnrQB5mXnOPCGOI0CGWpLJXJChzpOKHJT/tus0z9oVUvuWf1UcEhaLzXDmSlPq1z
bTul0Ju73Fizvk69ZqkK+R0D1QWa8GYo7KstlCo25yTZd17yliXu/ih0Lk6E2rJS
VXgl0nKE7IqU6Lx+G7PveAgeA5xtFRfCOBPnBFUkM5wLrSw6PP1kVuP1fNMc3pEt
iwU+YUWmlgA1QsZ8v0us2HHbmjGmGhIcuo8qndn+aI7Zpf9F5GnwRc7cZQ8hmd1J
aRlFES9jdrkGwZrzduVm+gGo8h1ICOg3vhn48UAk0Kv/n1Ts202badCjI0WAs1M5
6OEVcx1UWY2/5DJecpWEiWt81Z7T2A3wZPSdxnkXRs24uv7tNMTQikwNSu2ioj7o
uTmRoAtP3USRqsNbUKdbMVZJImU3LNMZ0qR/8pinuqUTPZGLJAh221sUizDnCPQl
pL80eBQcKrcU/by2DobmKmMwT46P9zEQMNKRRKxp6skm8c9CbVobDooQQr2K3uMu
JRDIdaubZXdjMzsVYUhxjg0GgHddH4IqJ/A6o9GJteVqUkYBOxjXNeP3+5DEpT8s
ZUBmVU3isoQPDS467xMl+bCbdW9U/FgMMWMmSU73ue8YqXmDT/OEk9yj891mrLTB
PcENmHNSFTU8pt/PRa8AeU4wpLNuiE9jFIA4m6l1fBx0S/r9mTm0tIyV75fbYJVv
F3mCcXpguuuhUjO5JMmr8NzhlShZdg1FnmvCiRRNnQo/CvfjpIuuUtADdZZB2xET
y1PTkih2ZW57ngbboPCmtxYsjhxMD0nbojAL39MUzY9h3gJgeS/f7z7tVx6mg4sh
ghowz2Y0qLHswARttblUbiGQz3Row95zu47mBYuufV8Q14qa1lOolLxiQlOEcP9G
/1LpCDv1oUGASy9yJaLt88Cvwn6gX5tWaStEvPbsBqQPONXeAP1vyOxPdkbuImKF
w08x9u1vaJSF/zbIlfSijyQty5SaIf3v1hr2c8C7hRwKqVmTHu0bfxoGPdVGfGG/
pnZHKvCh0geOuCfQrBA5AvTN16f6xm1ciRvAzbxnUjZuTWqD/AjvJhvK5wSKV3EU
x/TsYyiMMkMLpS7VTQeEo54oTuOCJS2cBVdfplNIQ3r2blQ07DuMkhgHb8QTlu/O
Hcef02mWGpLAdgkyGPzRty3a8D5GOYqO7+VcnKQwNkxWNEuhm0ba6vDhsSAlJYKX
qg3Z1FT1Ff+RNjXXc1WdpAifWPV/8fblnm1iE6ESBLBZKo1Q/OmAU7tYRaytUAns
eY9ottDXY+yspyJ89VPf0KvWpFVf1ffsZ2Cw8MPAYyXDWnGA58kQ5vM8M9jppL0X
vr1elfR3PmLb2O+nAu9qrjLu7dshFN9OeBkh4NJzX2+v2eTa/G1x4RPHVuB3pflk
mJH2CXe9ZJl2cdoLsrMvYg+c0nZ/uvZBi90Mz0aXP0p7hb80QiXCx3eKrAlmFhLi
IF5YI8oo7R+3t0cilm98+fCClm5Eyi10xlmh3pjl6Do4n2r6cVAHfEE4KiJeguX1
DSWUcwSSG1cxp4tIQ6C2ELn0YOawY3vlnV22h0mlTD4lFnuT7iZPWUn1v9qiwwcP
OJfI7j17gznH+1znMEs7NQRifIsrgFfypaqeZkgWR02WLsNrbbpcJOANoVihoJ80
NxN0ZXPKgflgHnnb6Jik1ALlt5en71Dw62qwgA4G5aC/EqvbSl3gKAAaSnCjwLg/
+4D0Yhb9ROOH8ujNo6ncTEyjDSWmn7gNSP8aa7gpzoxg87nXsImX8MgBZxWh+NF9
xN2BXYZTOoX4cBvuGiZinrNnOrXOpv+RkxqFV6vi7iu/qR5itAHArFhF+bQxydTJ
sedabSbLwbwho+Q3d7dWiUqknRJ3lZbgM78aHzwIUzOUPoarL8SoWldwbfWPaM/L
PDgTU3TFel9rfpA6iiqZhpzeDq/dDyyFKIiEtA7NYUsGwQhta8i7yyFzOpmSUDTR
IjiGvxakUlK9k23PMywR+eAUdVRdpR49wNL0WBs6K9GDmAdTIgrp81OpHKWxfNg+
9EIaflQRzYeYxHzeaWI7guW49T2CqBlsDImFM2XquXNBO7DrUzgi32uVvnPcrtUK
7nVCfsju60ELpJZoPkWQX6WkY1DaA18BWI4GL02z3Gyn18KrhDy7NSKRYajKtt8u
hdXMK41auzjdScRyKzvtwU7B5MDOwV0IXpWKBytIcYfnpS8WXetRPrhtxSZaC6ll
WWMrUaRUxwCNDNrmiG2dS30bxd3Si2LxEjfLGw3k3BcPxsJxC3AFWYeWyfdNLrvd
M30psiiOSaTPkPjH0GYvUHaUJp4r8mYGHDO2P8ibU3DVn1gHsauB023igtI+vFtY
6u6w5m8d/hlOyop5HqTRAeXg/xOJZlbS5jFIDuPkw1EJmKqbMlnZHONVMqi/8wib
NPCCIIIf+G6JdH/UfGm7QU4u/5rg/bTb/q9OeKzhFY6UoSwA2rHXgpie7W9x5a1y
kFYTXvYCCFC3ItyrUE0Kwnlz9/nKn9ogxDKhcsnK3Ci5KJ56u807OdrJao0xCCHy
ooGjNRkSIMK0wlAyW9zEDtYDpyiccoTPdLwwSgCPvmC6Ypf7HbwqcjXAzw9k1Nvd
vC2JUr+Un93sIY7ekTAjKFbW6mVAZj7gh7zAAnDQxgMQrlgJE6cd1YKgXwDysX+J
BDe1n/Gap7PJaYM95T6nx/AjiLOMlK6XyhNbBvI0/td4kMXhrr8Y95cCQVJuZhsP
bXGVnXypdgan3M0dlh2XIDtk+bfVPzW7c8G3uFM5+6YWmT3PkxQaBWd7SxQKJWwQ
RGW5yF6JjJAy+9n2KqgiutwFZDT+C4i/nbPI4JOkBElA/A2y+rE1M/cyw6/CnyEK
BSEVI0mBzJefDixQ5zNZRAAPLN01aBTEq+t7G5y2HtU364l6Pkp8Y0Daf93Y0Z3m
wWZnpJA6XpNN1AMUc8Oqh73368RUASl8IiBbUdJe48NSFp+GIz25wk+zjobv9k7a
Zfax129Whb8mh2yk/pgNbcPgoZofyALJaapvr16ClJH/tAjD4sL++T9MxJUo6amZ
QhFQD3nWL9/dfBeN2VFtfOb+V8iQtGfZgUDnGFjm1r0TQ5aJC2vFinfqTaf52sbr
ueN8skBCvPfEvgMy+SYoeqS765XH4GVwphbsxz1cWyX/ebniVqNJ2AqtLV05ocs5
X20hEixu/IpGGUShZUrUKPDvbc/xwxa7cMN67Y9wTdgeLzzxgmOnhHkJv2Lgyvp5
FoJZLlcuV77YVLqHzlzQjJMVuOYTJSYnxjwNaxxNrNxOAysFNIiVC7eH6mdVUttc
6t1qKJPoYE6CR6B9rm3ZucdlYRyGfwv/OEGzZQxr1TNOu070k9Dmmb82aqSwOWm0
A3cNREV7CqAZ5dCd3+JLrPmrpxMGnUv+qyo1K/S24UiVdj4dXYai6oejwevpqiL4
sKaDqHveUJ9TnGswTStKerliiH3l/OEgEddjfetKbpUqdcsAl/KnsFXR+Cggomaz
KDBnwS4Jbemd9+WEuapBA3Koy2LrFKQAO+oOpk1uwRzXlF63IwxpPmPcPukY/d98
0htGKhbAZmtwo9ezZ3+3CVKT3fSbzDo3XeTGChQqhBFfr2I7N8GYf0Fxflte8M9w
ihEB3348zPLMYh/WPoALkeL7DyQFgfDPH4/wru8jElFtXOIIYvGRQoEHIOVKD9Lm
dPRQxcQ0EXN8+hsNozlgTQBoJHt+2G1xk9mFeDXe8Op7GwMmpUCuqGJ7U+DHAFw4
d9bF2dZQ7+Eu+XfECZ7CSxORpqO7WxxFGIcs9K4FIS/EUBQqe7BidWPsaSZZLVC2
G+QtN4p/7fjz++mWO3HK7uKQzhNaa1vM50MO7PBRKv7CaY20DAr+utCdZ7one4I/
VkaeFOMnzcV22IO3VY77ICgUDtYHxKZL241vTobpaNsZJwaJwrW0NTT76XtuBQS0
guhU5dRie7VxzJxo6Vx5vpk8KbzKPF4CEUOFCCpIkhwcGJMJX0FCEOm40WYa+IhG
zkuNQ7+LLHz2qWzcFrhdj0WXVsU2ToFmdPI3i3I6y83Z24S/DjRd9UMuwMUTVjF3
Z6NcbGfJdZhe/T6P1yDqJPAzYpIKztfPamtzWFH64N8DuU2CCpvVgYuGMjBS9GSq
0IlD5KW8BVxXqfycyX0YdMZ0lEaEOsZKxfDPAXuPAW30RWzIFR7gyQmGVzE7UMOP
eF1wM+zydF5o7zllbeXVil28cI04HighmLBBvV8q/tgwPi+ncvbOpeK0ttNsNyTX
GaZEu1rlUzHpnRkA1CwB8t2GR65rIIMzcYhn3I3XTPC3+Z24yGufP2i4GAS9Tceg
mYkviTv2AFRESp+1pdijudKnCsZKyPDj1I3Tnfu2gHXwJb7jI8qWhYSohNRZfS/G
JujYQg8cmjTboSQD5xeeuoBrXaqENVqiA13sjTIsUuQV2/6SfcXsfvLE4taVhY+j
7Ng2xaaIIIoT9PCA7YEoY9tac+jJ0n85b8yC6A/+3Lo35JNJXajF83E2K4XcTrzl
C5nlaiLoiYX4XkaTnwIPpUpUt4zV6HJSY0n13HcF3BLN9YSunzFayUVjve7dK5eD
z43kdhQx0G6wygwaH5VGAxNb7L23nmV08FMdizX7W4F9ncKYEln+5eYxMF3MZjwe
2HYbimVd5l/d57wukcBzFmlCztx+WLbMAv1zjBGSf9j+fIGy77WfOiTqjITczTh6
LmCzkVWvf7dIa8Gk+q5Y/fnuKAUWCiAkAHc8oV73sNCYxDCT3C8pIL2k/nX8o8mV
+bhZeQTeDljF1HKc6TgqnFEk38cToelNBBlywCGMeO/kxH8Oios8M/ieqtl0tGYY
mrY9lu+wkDGCJisHP+QaDhTKZX6PeuIaOL0lfuoDcjhcVAjUwQnVCbkdxodQyDHF
V7M+mNyXInJ5xmNSInq7dQS8PU9BGjA5N8oltyWbJrjCVzJrf8iYSh938dDLb4uX
i/XBk3RlBWOfXS2yd/lSgmzY8dM0tthupSoyt9Xf/1f/RxHv4cLeOvLLUCTJcWcA
o7KqQUZPWF42vEB6pAGGzQYEJQ/Bk/o11uKGFSICfxszsny0epKRo3SrL8c3u4mU
Kdd9GERdb8rV1sOLXPv4ZbTJMUHnRK7WpQSzC05ysMHgLhmkDdKEjW3s64Enmrqg
MOXhqRyLNIMOjJx1nuAomCkKtKWVsBa55JLnxOsDcC/XTlQP63Wm7/fwpuWHxtvq
2OX8gRF2vn0pJPYZWGPfCfdT8LAvKNeWMBUVeo0nG9d0FRqek/08dcB6zrLMgAht
0QpmfMImZ/cAvfUNAHndy/nmRzIEC+yjA7DRCJjTh3Ri60hOJ1puxZ2uC4ENa9CQ
0RiFLPUvlH2G1cLkA+NwbTDU27uwUvCH/BoND9SwQIO/SUbkEn9PZQgZVkHvbt+b
FnF8lHZWuX/u2w20CmX2lbmm+N8liQkSvhPIhAbOxzZpGXXZKHWVLk18yOhLaB9M
vNXMs9tT/qLcLGXjOB2c8crCCRbAr8vidF0Pwo8KSXD+vnTFKDlNP2VpuRc8TY4Q
imdnVONNfAcIGxtmiu2esj9bW6mzN/oiuIrzHh0uK7NFdAixNKAuaA75VvbjdSAB
H1BoUkPKU28NXtMxFijN3U72+P95EKT/8GoKn0sZy9/6XVxf0losnGCmDmCr/4v0
GD0avSrHyjIl72WxdWbsL9x9lwsPDaMw5zaN2HhHknuIQt/GjoGD5+tlHUcO8vjy
tT3KmSWtK7UPlQKEIR1Y+dsW+bs+t8ZQi22l5lVlxyDmqAZMVu1ZK7z+nxAfnOZO
Xpo/M/4+WqTUHB9fIfRqErIjCJQ8u4boygRyg+4PGs22YMhGBsfUqZcx/dc6MVCP
v7m3dJ9noPjCFxZ7lqdCTSTrL01D1igsWBimYa/2xyo3xxDTLxHAKYuZPvYmtyDG
vIUDte25ZpzFgiotxHPJIdJgYI0bwE+VCiz2nVE1Ttn2Y+q+327jbXUomoekB3uI
GUTWIV/xmyS+M1lyj7pjw4jsmYWX/rQpp+8yILICFgCGdX+C23uCtZQv4DTxe1IG
LWOqa5Y8HXciufHO9Mt4ufzcS3N7iYZar9lbT6RD/ook8zvhU0shnrgOpu8wBsAR
P19pkqRuorfWvwgf+E/OUD4xDGyNOhnMjs0qbF/yOXEM9HROtMLy8/wuy40/ae83
S7CEk25i1KC9Rp9yDv0iS2wr/jr7fE9o7+AAnIJ3Xxh9T93gr36vMEVg/ahw35xi
ZVnVCcRpcOdDyu/T68X9eaKJUAoH3DeZ19kSIJDCVYRpauR9OmTj2+LZxXpZJHnL
XAvo23ehF/NiEAVUmpS9+x8TGpZM9CtKRnyvxGpalrtFhHs1gysZpkZNlF4Z0SJR
UoqAkjeDOy+o1JLhiiRBZ/P58cOl1Bkl0fcWyxa0S8jMPzl4KJZ9PysagrzSjfkG
caGwwH7tDrg2s9LB/FZhkuSPEcalWkWzfpmr97kC3Z1a3TP6Y3AOOolQrI/HXg7s
iFTWOEFGtPJsJZxzBY3aFabtw5y7kWjeWo6he7RJyYdW+ax7LU/b6X87xxE33FnV
/8TDozz3DnsdM4jhQlTf1WOA3Be7XQcdzHwZy+KgQ9ZQH5zlsm2hOtIdok9A9RTH
9y6LlvhP6e/f5pBpZaKahKoyzr/OuMVTMRYLKQG18KQx4PkLanl3TqeRWmj7Turw
Y8DvKzNKEzxknHNyAcpv+SoFFchhVoJMTNQb8rpdw7AuzNE26VXql1wq/Vj7bJhr
mr9PQ1RVnbpXy7/698lTSB18E2danFPiFs7RBGSfURn5EVplfTU9zvxIHaehVcRm
/k9ZQdLXw9E07pa+Y7DpvLh17FCYjkO4ydTcjZW6W96zU5pu2ZRmIUdI1KrqY92M
px2NG1/xFMSAguZG8RjfAXti5uB+u1bsy+gLF5XC5sxCaralEnUAL73X9iQtvk0r
gW4MWoia6BFImqVnahuRMoFiMw8EYmoyjPbsVeG6pq5V6Dab/O8UqjxbP41Wcmjj
f02UUHPkQCA/zaigS0F6Y6AKcEbUES3NBO6j33/N8nFnxFlAC+m9Iy3sUD/kwvGf
VQXv1GNwjUUJqKWdss1Pbhgg8nIPqQWtL7G7SaRn6iUJiZbrasVifJeDGw+l2hmQ
Dg7K7Rp8KW1K0kKjXVOU0F1vREIBk4lWiwPTZFs0qVjU2HdKAsYMPoRikVq13t8j
S8mEg4kUrOX3vXwnE9ZnS/RtTXLcvykgbUSorM05QU/BDrMKLjANogYb5aFZ6gsZ
4OmxGUPCVhnVXTOiz+cG0rPWWKUvMCqO6fqf3yMGQX0qys8vvoK4+YI6FGPQBhNT
+WGlmQyEt69+eAoReZASVYxLoENumpbrHzAZGmVXDTpAjJvQxOyGIWgeaIhebWJz
lnVzRzWNgUBYKEHDdSmz2YgPG2J8XrcGF+OAnuUxNhgwMmGW5jcuhXac7Po/SGf9
RqccK6h1TYETN9yihPGKSboEvGNPfhWvQ8GimLLJ/qn0Mpr/QUdezJZKafCJAUBE
xqKSIvWbQ5478jpc88YwE0F+gUCONecndxUkEryz7qtIIKdyodpy6qW6m4tfuCou
ePlbPVOj3cB9jlkO/LHxPuxRvgyW6FTD3wXRzmd9NtyiYk7fwvlYiV63F1MuOfR/
u9qFnTSgZkaI1UYuMGW14m8tJgweh6zW6Xn7MQ82ljmTQ9tfey6AzZ47FpPlsJ0L
mqvbfJr/tFe7NmbzSc94CMjicIPFbo7VSKwn4rOOCVmxncs9RxfNYEUdDw3L3O+c
wGZYrQgzBsEwt03uRSKm7oj4f9povLyEgOgBgX/NzXhER4ATLn2Zexid3CVF3W5g
407KIqhNAAZ7wfKDWlcQfhI58OpzZRf/3KRNrkUOqfGPT4Nad3qG8/KxWrliH1am
Vwk5tu3q61UT7aVJNH0GYfZWguXjbA5W35ISn0Ilk8PbDe5Bi9+XZkVII/pQOFrP
F0Lg+KdQwL5nGbLr4N6ZuoIbm6pce20qsrCzJhlaotgX7iLXaqZSVqzrOzWWa3cc
2YTMxRuxSYjYnTXpeXc5vff7kl2bCpf64O6LJJc346U0wyah0g4QDv8ZoOLX2sFF
26Oh+LDCGnfDRWU12fWRph90HvGtcwkm09K6BiMy19XWcu5XSF7ZyLP/JvBhHtfB
Jvo6FNXnGgzKJ+YZXRBiXVGsqnbGEn2Zw/Cv/j3UWLL4tp4IDnZIqTlDByM6LNEW
sMjATCpKwxyhAGjHU42Ub1+Dk0KlEVlY23u6qUtUCb+zWnNCWH4cZtaK1BT3cLXD
Zn8Vvg76vRixACP4XXsOnoMIcOzW6Ye0FH3wn59yJEQv24BFtKFZ2NY9rpbsseAc
K5+leyozSTNVwqmnXfHbxaK/8o5Ut+d2M6kHw/XTem9z5s7/1vj/2Dg5JOyvS5Dd
VgT1VjcQyg+YcObRKGlfhMTxXoInm63duukZvVNuTzDdesTOz2csJaH9Xp3IUUb8
fhjziqorPwi3NbDL2X2H3qIDbzEuKgc5wUyBcsPOp43tHFyJOwvP29g0lGbHIe+m
Hs6crGoIuUTEsj2el2XvPmKBHN5bXH8V1tnoJbtDG98aj1K1tYkaBmi7qTRtLx1I
9WBLKiQgzirwGMcDfvuf+itA/EKpRfHe23W5qa0fTeVqDAc/As+Fh+B1ZV9A4+Wj
TPC40zE4f8jKRzNBfLzxcAjRbufgpyUEUDmJUe83lTW/0MzE9jgfBmZlzx0fgQJi
1BACGnul/xjwvI7sXoGK0odsaAuwG8Oc+NIuljJr3BpSLtRHR/fo+SxUqXwfdF2U
UX/OMvm5We/+p6BxLgZ181AeoUTdrKIj+RfRItkzaFvGOwKMtmS2rfv4vUrKlXUy
W7TtHw68t1PyfYeHMBL+tH6qfqiRKO8IW1UPyLs6PvJOuS4BuaPpJ+mFjWG8uKgZ
z4I0mUwbE5tsCs6qbbj4D0n0DP+lxZ+fE8U7ekITohuoPvKvygk9iMFseyXYPSSd
CtImZFcDKVIWuIBPq7ed9IHmJ4hMbUCDp3RIhzMMD/pUCSw3lh9Ikji4lZFj7df1
kKKVUvM2N4pcg1RiNHwlKgurefHzFwytz5uQJZ/qfN3QvLWAG3H0SiMOHfamOEJ0
Ns+vDBkR+hpfkyaGuBDYKbP8adjTxYpvDsFV1nbnK8wmLdWrrmMeeQGRuWrAZKvp
QkqoVLOgnq/Mg0nhJT4mE3k89bkUyQUtzb7t/IJKwI+bfrvqxY4TVV3KuYnOOM0Z
ecle7jPx8oWXD1r7g1sWlf6++gVq2XJdcUvf1IBNVOc8K/kbLP96L4kd6qpqbxax
wPpjr29wyJEdNSyIZkFmefIhb2scxHsq10I09QN6PFs3VVmIVC1DH86RXWsv8fs5
TaX+nOvVse/MILxWX2cKNHXFG6x8Xq92ZtCdG2pklm46iqHSnL9truYt6uf2lMM0
4Kuaw3EYK5NKVZCsiMIU9XCzWVpO9Rq/d3lkanIY6ECBRVxg//q2VomXPNN+/5qD
w+iGho4RV7faZKmodAeOO+T/P61efQotk7rQdTMtU2ePG5LN5qaldZYG/x7kN9jH
oZa/H0/TVZkDD8pc7c5XOgOtSt9kGkDMrZzOh2Wqn1xWZNKA0kWPRhtca3L1jdjm
heTyqspFHqV1+gOE62rbgle+VGyx6kdCk3GaTl0/iUmEVCZR87fovpkyJL5PC1XC
Y22PTp68HPYta4ZhrPJKgO5wPKtX+ROoG60iG6OL5GAHiL3F+QHuw2mEql+biRR4
nP32VE9dwmI8VV5yGkxVU+c1frIDcQXfaesaaHLfsAoQxF4wKEdcoXS3pI2BMcQL
JRn6SwWovBXN4ZIGiwM7MoGy6xsVv8dEKwp4SzLNQMw4Uk1KQ6WG616DTz+GqVSX
QZj5QSaiBfLnAlx8KmudDNCRSvuOrZbmFNDLvLspXwkqtF57dNJ5mmtTjUKuCQl/
NkUCKtPGBNZLD+QKdm3OcOgH/iRMn4piab8FAIBqw3uNgxgVlln6mn1FOSdKTAm6
2NFEZSjAIQfPbP/qeJa/2aArf0K9dne/Gae2rfiubkc9VQ94LwwsyOKQh6EE9JZ6
90AoYg8pDKSAYH+2vmfdW26si99iqHOHEdOuwmCgo6C1hgkdCXod7X2jpcu5UV9G
uE2CU359445CM0mzZl/oMaVXi8KgZg7xxRhX5hOq6g2zbLSXr97W3qkJNN6bbuh7
4aRPcZAq4KeCAZ7Zsr1HDAC1sC9WrzeugZ1tUADF9hFKiV6S3hcIQFEJxV8epY7n
4xRKZBUZu30Mzn6fsgyT7EPmu2b43D4BS04LeJM4PLfNWA1lLyNLRNI1OUc61Xdz
M3kdjfumZ2a5TAT4PaEMxNKtsNevBvDel03fmRVQ6VAF0UR4ELczt9JghzIgphPL
AjZS6LNGMc6Ki5M07NbNJnnx5UJGnkIAT2K9txvFF4MmtJuIklgpXGDhTMNowp6V
5GYhhy3epgzqcBSMux1hq8riYJL+x8zbQkLWAbeKGiUWSidNSQWEdLXujJoWqV7m
A0vE9u6HuLaXIC9qEayPKF3jlXH7Zqti8Jiz6cwF/iekyipf7Jmk1v1SQ+W4hmV9
JMDZQnAFL2H7bk1fpUwMztDD4Gs7loQm33LH2X2qtQMbMkEjNJGCDwhmVi/An6cN
c6epFIqy7D6bmssMIAh+ALVbcjkQ/ssPEaLGzsVgvk337cABpdAyImkeQt/9tbct
WTk5iP6D3r7cNwSGAyYm6g1XIoANIDfetyYxi+5EOJ55WyCq/70V8ItGQRYWR8a7
Ozc0hWuuDv/hOfQawdsPLxlPnjp+3HecCWO9KuDKOSDPoWWD4Y1m0B61Ncc8zYBy
6lrZ+K3pa9rGOOleq26Ayp6wGtZVYH3E4+4UYM+s1fssdoCV9XUHvC88ctIjI8IT
SoUuDHmR7Skhds6ma2VBxGjIN91K2r8i42XZV6dew7d5sJoZErYvGfHWcsTAyhIa
jFJ7yuG04pN1eKmkMeHg7L4F2q7VNWEGI2am0gHNdTuYYZSRYxeGsVIbSTinS+5t
9nuxpuMt9hlx1GGf0iBft00KU55OxVVa/RIrzLPQaMFW3+ws2w5HhbsKChwqxu+m
dVWa1DePZx3aLMsFF2rKl6HVNvQ+5dYu/HFkRES4zo7XtwMx2tDK00s48pLcPfQk
42ZmF+rtiRynKwlJURGBBz2cH/I9F7/fXh1ZOy2u+rU7ZVvsanowE0TUK0e2EjYL
YPrdKO+J7Qdl3M6gWW6aIbJyEJjABj9Kimi82i1g5dDXddXnvUGS6pwFAWruz9Z+
tMVegNJ8yZq+ECux7FMciGH1AYB/XO+oH13Kp29usTnUpfG24mMg7LlNmgSC/oXZ
oHBItp7h9pz6PaG9WbYMjeM1FSDecdlgyva60iMoNwNcj12H94ZBd5z609csblWf
Zf1mz2kr7OW0ZAucEeVBIMjTqAT1QcmgQOE7MA6LZqjfOPbFcpdD1I2J4OpQ2DRn
gUjSpat21kXhIZfS8B8yer7gaboB/nIvmjGpIsI9EYI9pkNL1ZLXhMGF1LlHtZY6
lUCgMOKm6mxutr/InKIG/hHBC3gDP7BWnHLMoOZo2bcjRX/LaPLX2B4mUtULQz+l
9nBjim8ROlnoHfdMGDZXOUpwSUBQhlACh+T9JLqhjp4EwC4r5nT7Wxws5ttjdpix
Uka/vm9q4pRW5TfIRcKQJdncSrS72ofZ1ZMWRwZZ/UoNrrt7Nb0U8M0222Nt0QjQ
924VXFV5by0P0a56t4KrPsZD3iMnmMD+AJ1Mg0EjeQIFuIMLWE+DOk1nkggJNO0J
N+qsJoKmXQInmgXqAuH/lD5RoZGk+Fr8l0kKSoKjMF9D3U9cN5nUUcGFo00bPsub
Yrr8UBs9zfJqGXHTtIQ1un6tU2CElMU4X43Y79fQfCt2MHCB6jT+4ih2N3yeHuBW
2aOzDpJDsQp+emEaUCZ2A3R6GN3ePMTffI3CMKsbgBrrGoSwBzz9lIU+U0LYw4J6
BXqeXzIMX2N/njW0VLngOAVyI9c/tsXmIRD/fBLF8/x5KYjwSvzU/17LKT6dY2ZL
c3nJThhCAcJ4DdYtfTiheP6uJll6fhauQCBI8A17N3ic9a2KfXSZkJZekYCP4gGi
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11328 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/T97rZhQva68T7JOm4bkq25
b4BW57ADAHEm2yg/Vzsfl/h2m1mlcHDJHfb+2YBIsHqL4fJ+b75Z/6eZddD7E7O/
JDeGKAGcCTmr1jOyIW+gkcG4rcbl4HmcM+9b/J5VrqBjDotf+3WU+0CJ5oAC17j4
rzaGBcGGnopBMxgpkgsz1VZCnnnCaY2mxJwDAcKabjQEloECe4I+Cd0ej5ZUbl7R
udzL9z8GXPQxFtQXf/TecyldRUMHTu/dQy8qa4nCj3FqQFRQWUPTh0n9CoR1fVEO
GGyBcRLgstfZ99OXlT6QOJI7Pc65RtnbiNxl6dWRiy/X7Dm8Fe/1xFI5JzYB3XfJ
hw3wC1+dNNAoanxOHB/dUXmyjfq4zIysNVkVdAIZN1Vaj2IvGkPh5KVMHBHejzGf
xqlSSy2wV5QJqDz1eM35D4zf2q8qeuO6F0qnuFaI6zLRt+fkYqAfw4NaskN3jyju
2hOHsAiMgEQuJgcq+oezBsulaahDS5bhFU6c0a2VxhRiPKmSbPfnQ+AGJHDW8Zvi
mIXoT4ovb5u0RMruvJ9++InnhQbS/s8CS4/X/hsvizsOoI8cnI9uNormK9lQwEo3
8khPoRdelZ3u4Dpnl1bdl03WDa51WXOQXH2dkcuHzwxrIyBvaPH2dmg2j+wO1YsL
T0B5TzsAKf72ozxqEI6Z/l5vTD+vzBroNJtPPrw28HUDRRnOItnZuhFGf8FYvWLE
nMbXAGqUriqxFnCAvlLjG4euGKHpD0Jz/IudB6cRAHHlDetmaZ+Ox5ajXBXVaeVT
oo6c6E/HhW10/NXR7eylp+tSRn7sxObO7A0S+ZLm6ThbcLZd//9NfJPQ59LDzYk9
KMIHNvak9t6Jw+HMAJRzHqcNosaizaKz8oSyT8EUk53uBSDYF+TbfMHezbgJNwIN
nfRyIGbpLUqFHGY5wfYZQn8C6yBdoKOm5nKmtKWc6KbHkG8p0bHQeYgQo4aTYKvN
dTOMXGB/SIvORSJfsGZJJ4n/+pmcq1wJrsUNQ81lWbPRBIePdpga11dHNu5ZFQjJ
PMkWpqaXZ/13lURbmMshzTQjOkLjZpnEeV7MlmJpe6IJ8/qa5dThhSmA8JxRhWCt
LSoTB5yNh+rmwwy6VZ65i/1UXqyg9MtKxmilC6T6wX1mbX1KQfzxsbbn0MCUvd/F
vwvvpGvjq2zoZ4W7+WvWRU9AFzjHpkwk5vQwsxmwYdkfRD5/jPrrlPgVxGvsG0sO
Ye1Axd8KbMa/AglkywwBuwEc0aMY5IupnqjSq4JeRcYuFSLoOLZniKVx/fuwNOTk
ehG6KilcbU3asnxVPsUjBT6PcpUAY+spbQ30nFJuVGXG7RkA8qswNjYoJDJwMvLq
4NT/eyQbyf8bP4q8xmioOJ/gxmvBSMX0uf3pUM1nvZoH23mLWkKgtrEYMc7e2F/x
rrOOwaWvkFZHWfM8LVJOfAZHWQd9pjakMCOnRgKPY1688qwUb+IicRwc3ptW/inc
XR9IC8cr3tw/2L7fwQnZCNVAyND2Iyh4yUFsBfDLpxQD0cICh9yZJxtRUSZzuy7C
iK26xujn0qh2MpeBbIJYBbdZtEIXXcZ0lVg6drgt4lRugUrgBKoJ/+ZOe/nOtGP8
VS509p2KZCOoCzchJhwiewPXTyhMFJZyD8psBJZZ7bcPaZkDqlqkPBIFSKUy5fwU
4QkLKqbbq4ftWnW8wCmU2JlfzB1XwGsMzKbaax8NBbzRWJqGX78uajrezUl9yK9N
RpuCxNRygipsKjXbEOD08rUaEfJxMdLVkR5Mbs7sEpW7yxn5tGiyxKqMcOz0gGLn
2/7vC15IpHorJNjzYF5dPqnyb5N64dWMwNmsXXFcZDYCWdx6vEVa9gYgkC65VvTb
LmMipOMD3uRs6I25TCTYT0KBMe9EmhoWWuez/zZaNnczd5kWP0df48oEUewoYEh2
ZgQxJAH1C9pMq9ArGM3hBjTOtUC1PotaIWcBJLI1XTgBYIJlE0hz2OvIlnwc7CXq
bHw6QV/uJkUNakwPt3RBUlxVxc2dbBJNABzgvpClytMGM//STt8FQP/utjQJWyDb
JxoC9cNQbWE6PhZsr1xIpruCjA3XOvzrr+quskb+oeZPNF55nw+q9D6X3zJ5d/hB
qsmpSZGSD/A6lPO++C8GZImqDF8JwL8k6qvIMx2umDKaHO7HafzQ03f7DVjK4OwG
zRq3pF1F7fOUL0zmEknD/ANa0ncqWcmeNj22XJZWi0OgL8MLkuHKoT5VltM22ljm
urqnJsCKY8NJ2EdVf64W5oJvqE6BRjN7fTY5N2ZxJlWnjar4EINQoVmVKHYZ55YN
IdiCS9jyfum6pMqjWP5DFS9njINtqeVOHjJGapxoKNZ4Mte6iJwend+hske2wNQt
aPgOIbxY2cU8DsxRh6IlTvCf4JXV+nTPLOZAaw7eAtst3Bpduv3EOQEIUbwKAfOd
U6eSYeKRK+hs9z2ido5pCIlzbnM13roW3AV4GoQ+FJ5l3FcLEwcZLSIgvf+lobDn
eCLhvOrpE+kigHhTscQDny01C1WA8ba8Xf6bCq0X5FJK57PDz+y07G7GPXgLDNg6
+UNvHfDwDZfD1NHezIKu+mxEmtg4e1lcSrmXTHny/jSSYK2MfTthuFV5QB3PcDKH
1zvnO4SJIaLvuq1gHs6Jyrd3tuToF93mj8pSZBHlr6EaSscxRFtiNngdENh8sYPv
9SOmJvLCq6xyQbe2Zw0TxkV5GZM5HT3qqa3y2XdGWeMO7WpK04D5Moy4qCs8a7hI
GQGVViasmr+DcXvMoBrrLQih9uGlaq1ili22zFnduFj9m0lNiaQG0bFjg4WfP9Sf
Pt8L5qQbAz+in26T+TgkYwdh7Vv7zm1kqzWSfo8aQq112VJMEW7MZFYDS0Q5ldGT
g4CnWNFoiy72HIjLLuwnY1f+AVfm+jjpl4rlxWuPgCUOXpmnL5ZM4dioS5S0aoyC
AXRaP5DoUaK6GV4fCjBuCbdbGY/dCJhADCKPIZ4582+/XQfpvO5/ktPWoxEtPl9o
9EBIJ/KQl/8nd3ITiZ2qpWa0QdMIbt3baZchZteZywde0Gf/DPKBA3VD/yrpCEDj
4zjuziGr19zGFJq4z5UODb1JDeTnEqt+54+GAPKn5u2ANi5tSyyYk8OQCaH39Yo3
KJiMhxNz2ga6edOnrcBEbtT0g8YlI4IM3xj4Ht9Xhl1l/pAIi0kVOq07qZCZ7iAR
yXoqQ79KTyDJVS2mTKoZ0sGpQ4R/QyWFtZs69PiV4A6OoK8WictGYytIHuy6FFdV
5asokUzr9YJMlph6Fn9SxPyaqKCkIVwCAxZIkNoMp/hI8ax7sPCabWOY7YRAj2BD
LBTUr7HDAOHzIaO828Odfu+gQwBVYe4SeQlII/OI/cI8wwCHFPGnS+W2cUfW/0Bt
bMgyCKTftAzBAnttiihaOhKdIvJzHO027t5G8oTckZ+dxPpt/5Rr9OdOfUiG/V/p
tVQzpHSHoJQirFyNUzSobk8SW8TUzFWdDCs39LgnXVITBcVocffSme4SMaseXb/2
hwFMcE4vBQN0lOB5WG67EPl910KW9w2D9EGWqGs/DTSHQhEHz6mDUQHEsg39kjgk
lzy8BTi6RFdv/IPmg47qqAUcd67KebWpK7rjRuw/vVbVX2bSajR8qaV9lpHsn09V
z7VgJtlsXkfZam7YQUTdpMs/uFI2k0YbEnL/S/Lm9y0KcXU27YSeE3kN1nvUu5DV
pXbxVotyDSf6lg1KUKWvRUCw4A7ZZacyUHo11Z0Gp3oyy9UoLqSuSL1or5LBlzqe
deE+fE/nTXczjbyJ1YcZpIkyostZvlhMRggtDUWxaphrshOeN5KNVhZsm+FuU+Q7
uDfELvkJDzYpcl+buKs3yqKA1EZ7jYx2yEh55lIHQqYBVCXj2Kb8NA6jkhZsCcSg
bFt4/JKVrygpvdq4em3qogJ7iAu6Gp+ttiX0aSm8+gzMvrscVh8IfPamu+eIIrwi
IWExqSeccnAmvxogbpLdaYpnfZ7LMuNk2Bi6w5eBjFfySvl0q9gz7M7WMIVzxGBt
NHT/iAmDrmhR2uwr3dfMDC2aMHhx3t94yW3IIxoJWbTQCS8q20KKrUSKSpNhPD4Y
bhwqWttNwjDWhZszWFi7z0rUlWN7kup9oFcK+lkIAl0u8W7M8XXbRBatwkm40bzo
l92EnsLOhmkCk9mgzzspNQ3iUHgVHy1GlKYEblC//Xx93/SJSk40tjqkPjoHqO86
eVP5usF/HId+J97GsiaRIMd6yfEL8TqQ2RlYzYRTyMyyRrHS7913pgrYPKBe4um3
I4banXIGfecpZsJ3hH/Zon4OOL5wgsSPg5+Q1SzmFH/653TwhvXxGju55Yfz7T88
TApHqMdGlgKO9o56SuEbdsC9kY++zSWZWP4DH12mnBTPTBWeDaXfDmRiXFiIZRV2
X8PEP4bB2J2UbzpRlifh0tP/oZCovo5FpKDXYjGrqkndBVNr4fjgNAo3mJHCOFYl
svuXVtFEboLAEDcxGOw2xUWi2GCyZj5dLJhkdRa89vJJuPVsUDFgq0q5BpFJy1Jn
XQL88pPX5shHf0bIsULnMr0NW8h9i85bEYCgxOnimp2V1SjXLtLZPs3165DXZt7A
O9A5tfcqOTUP7lBdht+D4S1kB2sKqhNsXWV/0AGWYNT0kZTqUtioi1sz6VWD9Wt1
kuoc7jU8LZuijnHAf1kch8Z7KDOhPuOhNADbyPECeN23g78hqaZQUu/WIieEUcQF
+y9UNHUR7GL1bXX3SgfEbCotJReBUTHAWlJsScLgRyg0NrQbG5CRtlivrIKvyS36
gcUe9PNlSvMvIhuc7K96nlpz2f7hv8eSAMZGru+NBIz9wsWxTZApg4qyernP73yG
ZXIs3tZO4H2ov8oJlqbNKpQ0UdMtWHeNS0iNVz24wCqNlBNp1UP+4qqgeOa9ccbV
ltLLEQQBn2RUeTf9e1JDegAo7BXWo99SowEM5sRmf57CJSaqyaF59cTJNNnZsSPN
XS0Q+u2ZIc9l3rA47isK9KqVsOvVTZ4Hoxa6cDpn+63u+ESIb8pw1oDzJW+p7MKW
zsqxTesYdb8sLEmb1F81LyCJCobnqidJc8LO4xQzq5OfsSHCrcRmpcB2CEB64wkc
e/VEgYzomoYBAkwqmbYqjbN5UNOMwlRLc2ZOlglv04oIDqrlbe12kkDZsxK47v1d
rxCxkhPWtEbwOE8OvJ4W0FtpYOJ/Of2NuYMuIk9+YdAaPS3Dujq7WKFL3tDhgmNI
bXTpr5n9zebbPkOyXDnmN84KlQOL9TIvKFBoHSnWmLCSQcPwCVmst8LHHmZ6IIQ+
EDumhkrgquP+uVem1ffKBBkot/rGoVe/qd4yryRF3n7SLfSyP+CzuxWXrgY45N0i
UsTdHnmBXNJcqFJP6T6Rf6HzMyiNBCHDSuIr2Q1GgsslPtdtAqn0GcYEmlrtjx6V
YHLuaYTNThcl18L5cEzysgHJnqcpuNl9AwRfh+Eaa+31456JYb5j6wUQ+KDLlbgv
HqAqV9yezpQYF/HHcZeVOQafmtC9Zw8cYMn6Z47QGitV0JT2aQ2M6c2Ke+njDaNN
6obkqXrJPVAQ1AieTU65ecYuMvvYrKv2CZ+W1IYOyyZzYY9xxRn9pITxyjDAuq2F
kTvooQJBrzWQfv70YIgjz1Vyt09Hmg0EBq2zccmUHu8nSFryVM0ZDJsDpk92Dwsq
UTZ8Swq5hXaT1kBhfx5ihysDQ6YJ/4myO+h7wH9n93f+PjMVclnvr/XKv0pV/Vwi
8XcAEc+emRmtDNzqOrDnVjlQFmjLi1BxwYQ3n4ufMWqBUqKx9aYbL/rFtV/nBJyq
UTEWnrS9EyR6yX1uYOQrkIEU6Nc7oXRWQEa1oce7UvNbcSfK15wzSEk7ETgKtaKo
zzRDNyhRpHOQoeFieFgyPJTfXQggc1GXgel+ZRAcKXCuyNDzdh4XDfUphXAkf0YY
ddoMmJ4B0zewp00xtMnd4rmmEzo3Z8/L+GenLAklpcBwmB4T0ZNrdQmseChIuhXb
qAyRTCr0XIEm9+7QDqAcLokU9q9w82OHpcJX5FLPFbmE1jVf2sG9gs74Z/riGZ7Q
+m6CG1UvNeUhom61OmDFYcmoVnZnNlytPzSRH6XNUa1R8fLUo07476iBD1WFKxAP
1dzQVRV2ufT9Y3aOIeeuNuWsFhconT0cG3MtmDT3JkbWeu4WVx+HQxIV6xqdR57o
OWfq7Au17LnFTgL62wOUq03QIWuu9eCF2H8OWd3ZkLtDKPsTzEzXjDb8MRJAh9Xe
tsX3LLp/uv4HiYEyBRq7mYlmV0DaBo7gJ5gbVhGD+LUL8RGSjIaCYczEJrUNt4z1
Gm7H7EjMPG98pYSvyhP1ojG21xtm62H8GzSC3fKdIUR9bsNkCP61DLymc1RYF56p
sfmkjDkESofZ8wkKTF2irZgEV+k6+6RqD44AnMT92dS+V1+yYlsjMxrTHVvMLtPF
gL5pwreoQ5Y0K1fvYSSR2jsmtTkwQONIpIZoCvKdz341Yl38sHsiQTXprwY7s2h/
GK0MiLdhY2UBLHOrTFvvmZNb4lXEzSqC9soxqchFaNG0xnHBFR9q4oZMInSuL5AD
7T2TDzKM6N7is/cIYPa1CZAydVuGR3OEo18PE81aUBxk33igGwUZd/Icas0qvouf
0XIufqnFZ0bWgZWJ/jQZewVxnQyEBI/pWuRI++1t80MWXRE0bKCPPsLXqTzTRqbA
CLGetKroFIp1qCAysslP3ruG0evrilhWrVxFA4orlNIVBb0wvLV5/iV4BS4Sz4+l
sLgfj4Y7qpbdmRpbFabSBjvqR5zbEuqgihT9k11sqkSZBg2uxXg1oTzmorkuDzD0
DPJniIgptcCFZRquh85mBe8X/+Pfmhh4Gk1TPk1c1o8QrgAestQfE8BnsvI4IqMF
moB28S3MFUUc2TFMsZkAs+QJoaPid6OJVfgAhyCoY8Kp7a8Cds0YwfLaJZxSHRt7
Bq/gYVxqERT5Jn2lHs6PrJts0i11yNT5pcv6Hd+GdRxOkdSqStTnGou24TvYKLEx
aQgzB/5iPsCE00hv54gksVF5/74vbCleV4H09Ml7uOCH+hcmJ8a7wAWtDD8Ql3IZ
NIcFvWfti1rHtgwzO33b/EJl53hRwZ/1bEDWz9wljfWtAu1QI19PWx+ZyXV3laPL
bdqJ8iIBKkdQxS2lQsYnV05x8g3JZeeVUnOoiWSr/xFBAWpuqDIwaSmJUN7hTMQY
bggTv9UW2DsVGwi/Ay7ds/oax2lDqbOm4nUUrImAFrA2C12q5UVok/5FDKMW9/yH
e56+9KG+jwVs71MFOpihkWpJGFtYNao9AhZbrWDFs+DelIjHvQvAdEOkmPJ5cxbh
pIH/GEPfTw3ogDjhcKjp1ytQ9acecUCqvdNKBa/yE+5TlFbacKb/1K+Eb4/pyvzS
JqQFhC+P/mnx7RadQFyco1JqJxugZLFridPWl0OSM7miHL236CiaJKdAztmYaWlA
wt0/Wk4W8zfBwQqWQQFBe7v2o3dhmXkhaUxHpL6gAntjBOiFDEHXmuvVrPRGXH0z
4ua37zeCGY2cbEBAXeyVmIvtptl2+GNo4oSV9JS/Sl+D0ARjh20OkPCDwXJcfI02
pYRCKoDtqxmRg9/T2LKnM4fG2cR5GpMtOEmhVeQ7DmNa43Xb6prDgZJMzqFsHDmz
yKT+/Sqjlo+Ub4AngNrv/K8dM2aPDtmBp8KO09ErjJGY3D3WLDFf1dxMjAD6LJGU
4hsEgIkQI8lAJt9d6Jd/AoIOfJq4wpY7ar/d+B5ij0ePpKWrPA7xRjoQrgcbilaX
ESDM3ANifLzSusgJVxQPj69JEjfQzMKYU9UKfan5ktz7OoQQQTroNVdYTXUh7ov1
D/+MHsJmo9yxOjGGADqC4vPonRwfzfY0BxJxuda5aNtwY142O2AlX56MRkF0u6VE
DA7OMozv5xqRd0FyVgX11CtC4c3F2qWJPmJW83nvBy/nOYtl/Zh+KV/GNpP5Zwfa
+kh9RRcSQ28y/CzuaiXjY2FCzn6qykXxkUWR1ykVha1ka1Nh9T2QiDTggxwaXKRe
M13tXG5GQA/pOnQCDkizNhWxAZMMTKK2BIBsFeR/MXgfagm62U1g+2ZP88jRLLim
CK5oCqxrX2395Xh+5mVoX1X7NGwpFZRntDO6Zv6KeF+Jf9dS9ANkDgC5zLzvbpe9
YuDelPTpXp62mAJ55Z3IIOD3GcK/KIeL39PKOo1fcgoa39tfqz4yLO/f8CewBzP1
Y0wg/swv7wB5SBrJZegXrXcP0Mn+K+92T1lNK/ksphiocye5SNdxmCnWm5PRFh7a
zuNnL5XaUFXBHqRPQ7V9YiQjGBUrqqBi17DacShj1vXGQeLFKosXS6BqCV+G45Hp
Mfn6YoXzzsU27SfCG1ueB9Z/LFSA13IA+PGIKUNTz5A0r7QF2drWjvwogvVe0ADB
nAyWKWYe2lNn3fsasNQmSt2Agk7SrCcOhC40xriWbtbqiiUVPgIFPTA8qYfqZry+
AGzJVC7zJZHGvWcfBueR/bgUSOMmGVqzMTUkJMtNbieIV2yC8yjYsDPQnJatIye4
OH1lmVob1zJFOeW4vKr2ABOXP1+YW7toxlWO9ZeDadQVUFUJjivgP1fmD0Q5YOXQ
xZoHImyNlJaH1Qa5J1fQ5Ib2FelstMnx4y0KcDGnxoVuDCCwZ85rmNoNF2uVNjJf
CIWRugjE4f0AymW3yzf4D6Xq0NQgLbRGfDs0+8P7nqW5St7AKzqQQ20LdHM4XmNG
MVqFXuPLTR6lirP6SNOdR1H/2ZbDnjvEu3mNEi7Lg7Crg3pZMVa8Z8yxzVw0h9QO
3pgnn9wMNDIigDBubnh2Gs5ZajSxb233oVYbUVPyfqVq4x6C1wyWjrBfRbIRiH+J
vflYse0754o5xt3gq/Xx4kyxBkDyz9P3IfjNfaX4zM+RDslzT0F5QrmrHrzLyDdd
bQa02NActaEatjSfH74N59Gw9gHkX9I8VpxEZGH6gPdd6AdiarzBX4dqCh8fO0Bk
yW7m6jbTsyrfzFQll/zlMrjZkks4MnDZnlmYvb/kgbbUr+2icU2dbkNi7Wu+UL7k
PtcDxvp3SGQbUOZPiu0//reo+fc9azHhKT8WvpiATFTJU7VNm/ot9yhjd1tin+DE
43u7eUOJqYAQYFzKXbRbtchrfPAo1sT6uh8sLfS/QFWDdAqGThYKydiAgN5nGdpc
JXPDRMSTkCR3oXkq0E4gp1DNG8AD7CuHVn6fnw4B1brpUbqe3G6S6J2qhFvHlDpV
5LiAI7i5D6zRHljwKrObf+fkzdVH7P8nC7DTsv+Ie5xdUaQayCTlFenWSkZnm6mE
gm8zBcoIGhd5amCQbFjBHpUwgRprlc3i9X3qIu6TLVCAEqfna6B6HO32R5ecFAwD
xkw2b7qevNTZ7j0jDuJVdTp4n9AcjFF/f04qIWvKk6JOdlifLzEQtcN70h4aW1kn
qN1GdILACO8PCiwEx4vbGeF+RSZ/jc2IvJpQuF15r9sK1QW/WSIrrcL/RYmHYJt8
nvu/OZfb4wC1SVP2kPJ8wFcRU5Ekc5y8efhmRRUwCOj1lmKeuZCHbA1qECblrkZZ
5lhL8QjyuLVGuv59L2WVC/IEpqgtvEPruky5H97XAhzI/RA2juhC/zQwndmfHgMC
Z5NtA4EoYExub9SREtZj3SHGj3ncisRqjCNhxFvDHiDMnlMkm/K8LMGYXSVaA6cm
Mc4J/BtUNJ/496SyhMboryCE0N7J+hX1H0+Koi8KUZZRtI/X8X+vD0wMLfrzGRNi
zfr6bYlcNnoFvCwy58IPPXwzrAaXgGEaQbRBWHJTWGeVHbSVGgR3TbG+CCdhw8DC
ylzUQCPmz72S+ci4JzEFaj6HR49F/1cs2b5dhq116njoWXXzqIaMVRGH4jbSZZ4x
mVHXajl/k+hNppc7ah2ER6LBQOT1YrM50RTwOdMzyiyL4kjOmzsMmt1dYeuzspXk
bpOGoJ2Bd3Yp7VCS/Dl/L/ubzrUcTtIN1YGL+ta6H3l307yK0zPNMxnUU4IApQk0
BkdB/xE3IxoTa92PGC4WhbbH2ZBm77O76CybJ+3ohqtzsBSpkCm2rvwalzHJ4gxL
TgH1urOpE8R349ABt/WmWfxw+u4DEesLeXVOMO27S8xskBm6B5SZtfD/UDOfx3mK
zNeOWKgEL780ANjFXBWmb20jYOBHqW7Bq/5TAMgBfowrRoyNTafYKFzBzS8lC6tb
MMZ8G1wnire/ApiGr1R1/puqbu1RRrh0G85WO16xYAKkP/EzSQfuBxXjvPoeZKGb
zZjPCgsPSSzQHYakJaFftGcZaATdrlNKIojWagX5Bud+di7VFuUGrZgn8RnfDCMa
XP0Jf8EkGL1eAVuZBfuGwvt7YGyxNyr/ZBLLPIPXhPwGK2eWgUsXw0SMuPgmbt+X
MWoTi7w2wNgz8GbaIPXRK8V7A+yKOvyAZyXjyp8BmzsopstFhmDEKZ3he1XMV9s3
4F4i7PzC4FxDlJYUzmIpb+EJ+rFRVmRr0puq+QbmFxJjaZ7Xw0HdrcuS8KekaC6Q
VbHS/O12brc5YRU9LpuYx+0drA8RpjbU9m3nsx7dxTBUbI65rUfIRdju0fToWflL
tv1C12iTSb70CueECW3kHy92alth0tSGauABwvcuaHkRPo5PWgvsVqmJxP2YBtI3
MYHPlfmMINdwxQmQbQJ7BNHgFe7ic6FGAWY1IlILSlf7uERTdL1h33Z6dGk1ZfJh
3is6b6Lu/a3YH68oBDWFauauo2du2VuguyCRNTBnTZ0hpl9J3RX4vD04YN5YS7Gb
AZ5F0aa1mI7jc4IxLNBSK2IV3JJ1PuwMOKv5Nv0w69ICp63/GILmRQghLVHLop74
ZotnkFJqmEL4VBbtiNKDSCbt4vgUHcBa4bJ2M9piZpKJhq/5zT88LRTEMn02IES4
CqeeudKC0uYAy20QYsch575Rk2ratBNrxNyuDIf+pUQzat3JrM5AS8IYYaVrwjMu
DyJUZuPHC/CFTYrJyBd1uvMyTTF7JcNscsTNgq4UeMokt/u6lV0Q7ek8FA9iaYvT
pfyBrjInxbyTZkOG3uWSziunU5fcojSfNPChbe+rN75GxtZBJ4RotQV4vCzBI16a
6v5RLpdbCHqnZv7rj2i7UddaZn+Evvx9Bp+Fssu7ijGEsEMw0tRF7GmACVXp0dOf
4nxOnvchyc5XS7la2sPxDO/B3jAtYt3f6mc09U84Rbtj3z9cOq4RYuFXN7K5pkr+
+hL4iUdt/77EzfR8/stXYU8R27j2/z4hqt9kYkyv3myBN/kAsJ/C0HpBd/08CQfv
/1Wa6j0X2mhKIACfQA/NuatR1AlMau+tMe5hOo9gL23BonES/WENHoFblwozJNwv
PtAwPiV/nhQHSoLYd5dG9ssvWwbUa3Bh+wbQNpyY0AXqZt4lyOjELSQEqdKA9+ha
NO/m5I1ql+mS7iFbhUMTOz1+xxyOunh2EQrvaSzyfJun18VByMKA9TR/bOenCplb
6Sc6jBOmZl3efcSMOvACfnt7rP6/m7rfwtzky7czbc/FCwZHZY7APTyQ9F7ZbCGP
TFGNBz+loBZ0lptR4r1SzQuKZB3Sq7hXl+yosyU+jUoXFF2DHySkurY6vOwaOjI2
qHRktuRXwf0Nfqu7S3s6iPSsW/Tm4MerCBdvDx4aQ1XG/wPaYGSeYXuSzuMWe7IL
7hufs2i0yv49KQsQTtxPxT/4DOUpmJp1uIMy0HicCUfHvmvDlLHs0vw0dJreyxfr
0xnYdmRJaVbzTyKziKt63JI8HziWPgRsqYUa1fZBpVoa6HICB+8PGZrQpr9inajX
xI1+/dK5JlMFG4m1x+CS4uAfFfR6I3YIMLishPpGi48lUDKDvexKde7nQVR2Mgs5
7uV//RSOL8CxQw1pDhB8x+/fQBwXwkiKQFJ7t6rStBCAlu0kaj0Wjkv8n0kmnBBF
vJESb49pu93w0SuLubqsJDyKcKe3vq+t/hHzhSeMX6rLvSKTtNCKRmM30LBt1iG9
J01kzrMNZupAajQ6Q+nIDtIvIE8t0fc14KStOz+CVu2B42n5mFjU6L/y1D4sdUMZ
yUlc0Z+o1YsT6N536MLhcpYLmRJICq6gDG0DmFQeXL/UtyHxd32jNuRBZmLjuGD+
00I2ynbVo3YAriB3CHnz9CFkHOKgJCHy7C3N7Dn8esFKN5TYfTTyciM7C1o3RDli
i/tngR3t0Gw/u+ke0Zz6+AQl5A2wiYlYRgv8nPV5r9IrCgEHSqlxgdJmepQXaq5Z
gwdwzwMkQPL7gm5/J1cuyK9PGSxyvgIVowkXSvCHdD2fM/6xw4YTIGdcCsLf/NJz
T6UqvtYmp6EM1fdqknGFsiVq9qc654Redf/15wUovXzKUdDOsnsMWNzM1KiExXHL
7WG6GjNh8ofpvK1nPzlNwQF8ue0ZdrYzOp/QMCOHaBupBWWYOqw9A86JghIOPoGQ
mu1gstv09ac9AEUyclAQLGJCdzEDyzrBKPxM1TVCqLp+zPQiLqjUpn1G1NqoZUlO
8hdg8GFIn6TEQDWD9pMUclRKHhfe9Gtn7vzlU3frl1wAWWZj0eew88aIhTxOkwg1
fE7K1VnDUUzB+QG3/+c/ViRWoyjPSFzX7cuuRiHxkeGqxYiPbTqw+Yk9pkRjlz6H
L04n/StgMvLJreaW5mraM9kABhu7aShNlDl0QnaFQXbq2EGulTB+MR7COwwrUZhl
+CciH0pJb9UyoPk++Q9b0nYHLPY+zffi+WZRTye3XW9xrHjWyHKYkmIu8qLwXI9x
192cCMD8Z2sA5INidsK9WF6JGXtXhEujucYkrizGAaLeq/dsvBLPPG//ejhozb8z
c8sn4o5vXnXHwf0ko2KgtyocW7KJoptH2gSuvv9IlAEmLHFSTIGY8oe44PJdq9z/
mnrlem3Pcg8LwDOeV1mJ1yJppChrL3D3U+LOUXpCTDfUpHZjnbpO1NjSEhKyup23
l2NnO86d0khxD8/xhCZyxR8U96UMFBorqM4jHSX42gWFXmDAbnQ01XkCg/m5p/jg
M2udLs7Zdec2nqpOgE2iQIlzlrke3enDpq1+W+bjx19M0lQUqmzHwOFljpH9V6SZ
vrFB89tY2ChUhJiGPcoFECQhQYVt3jy1quAMTTyPA4kNYl3Uh5TNrzyUu25ql+hI
1pXAi1sfBBK2qFFB2sh/OpiVLEoGKHKYDCdNxb2mc9wKLtTJyarCMLhzl6P5V1fd
n+A6y6HqzAQ7wFZQwq/BkgJwzPFPFb5ohswdL5EnPgtfWACv7T7b2m/v2/lzw+Ny
L85eJS8+MdMkjKzXBnwt77YWPVthXq1SBq37z9cixzc2iKa2duA47MddCb8HF/WE
5kx4tQLSxzYtAn9kHYEupE5XajpU3fxWcVVCj3lIQEmrSMRnc7sKD0hNQfWOrmy5
ulmRePZmyFbaCD6VuwqgqLv/4N3vFC2YaBrCjZAr8ClrqyT3gHg0iDJjTuwilf3s
4wflRYar/KRL6sK3ZukbmiQH09KxGxA3917PbX1xv3MwsS24nSzj4Rc3m4q19wro
+zMRBWuAq8y8uCLJ7bM/xGESd0ti3jj2srW+3uqNais4Ium/8ufVwoHJnVRhJbnN
wbKVbza0w9RIZe7PUyDTPdt7XHJigZhL27R+rUn3NMnIjRasckf3in/smI9X4pHk
Hdp/Rk9feaXFCAYsKI+w+IXC8NYWzjBYxHr2RSgwqWOJZRVt5xXih1D2nqd3sGZx
/Czte6sEkvNJ/hHa037ooAyLyrvLnxIElQ0RKgk1rk1XJk25BtB9GBVwu3i6Q5/y
3yimcui4kUwZm9Pl4Mas8XFR95Nn1KE1dcm+bYwOFx6UqMF8OrtJH/SyA3vvDyKI
1anDL77lMc+ng5MCa0rR+IBcSfkil4jJ06s5xIAGcc9hMNTiYHg8g5UoAPhvTBRI
7zqseBpCbSfkHrkjIsJjQMrW+Y7RtoSr87LVBnKhDsyRzKBy+cUDNMbddkyvw6dj
FCG8RToLc6fWGhwMylDWlviWs1c4jHKFfgkg3coceOXhL97sPSsEtJSbOY0khC95
qr7zhu4ac1ircI7I5DKzUbhsYooWKSXEaTJghtTsWJWdRYKuzwVVsxnfB/SJNgOC
Xc93l+MIt55Gd7NzYFjejNUKknaMWoQuO6vwILKQEJfZSaLluYR6C8LR+yfZlbFo
SW7PUgax4LaLWRdyzkB0AqJWIKeTknNTPhLA+k4tTjLqJoPhfqHo1+fyNyijl0hg
udI+IkX+sMWsteIWZwzO7SoJYoWOTh0BbhCiwfXrVzOIP0iKsTs4W62R6jg33BJ2
8b1PxbViwv+dJEugpMsnu3l7lwgr/alXInIJ58kEhVwdhgFzj+aNTXpYWL3x3Z10
JWS9U9Gad5H64/Rszwh/Y5Y7WocV5j33sOzOe7Vv16pwQWFhGBb7385Ee4OgKXJH
Y1ECtdyfihSG3rGutL+bsKc18kln2xOpB8uwQg4882q2gmiTJKTLqrSb5078LaOf
NRApvIGHFyhSkX9s5EavXgzFdpPBbwT4N1p/5feEaOPVmV6hqSGUioplwWRDEMe1
bS87RUt198VUTIvyCo8PZ5vQ4abG18U9fwANT/Wnuh4jnH9z4wddcPe0aHn0hC1w
yIv04cnd4+9oamcWIdDAjlwA8kaZbtU2wXCGsSOC5l1//2LhzhSoXu0NyiNOGm2T
CtwaUoXhNBM1jyo8e1SUguHjYEcsgROJWIWfPc1TasH3nl+D/V2A6DqiGzzznd/y
aYM8iQBG7wVw7LS5K1/b1sgrqJc7Hu3TK4Ahsroxusm4PV0X1knQ3SFk9Ljquv8G
9c/TkbAEulPZqWnet8l46UbjlYr+gj3q5oDy/sDr9kcl+flB21SZev9USVFiJ9V+
mxfklkqV6vQsYeDkXTFKiudd7GusgEtfglZ1UfxkphsqDuklPd7UIS0vu5cKUSME
>>>>>>> main
`protect end_protected