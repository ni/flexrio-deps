`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 13312 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
DmI0zUXpjr6rtg9EJrlnT9Vaz5p6WaYjikiX0c6CgV69BdZOibD5YTpLplVos40d
QCo6yY0mm8Pc2veKf355QpYktIlDiPtOvKKER5i8XxQNephGKDeSrZORmvI2CUBu
M2hbK0naC8blnkGAOTc1A6VHQL3tAH6/7Non23mG7xBblx3Bm8IXTtUCNO7qq3pL
MMbyu+fLdi+NjqrHLSgU+pui9c0sSzFcB2xQABCKFty0e2EQDobK0TghP1m8Vo9Q
0AYHUsqZ4EzdBy6RwL1P2qZImpW0f2eHgjk6RE6V96/PZWPOZlg0vpb/mS+jKva8
KotU4tXCa1jxOrmPsIu8vR4rg5+/VfZBJ9BZyDljIgeVzChDAxzc5u/kbPjRCQ74
gMynDcBC66ZBev0w10tXVu72kLylxFHu6PivxfS2LPHDSpe2+9I/jacwt7cMewg8
OthqklxuckawbylXkGrQOeAhRv+iOmR+9ILT4mIVD5Y2HM94MddsiYYlbuI265Ze
tpoUWZbtkMtpRz45t0zkN7xbkid1ZR8hDWYg6ZLhODbqKHVELsptgFWo+oMhbKgn
CtVIYNLdDFRFns1YBPpvGLuGgB7CLb9+S0gySHn81dUM1p8SLh0jPjkvK2VEbJXR
iIwn3pAfjEiqwefmwXhF/t1YUWtnkddZE+8OST4jh5hE9utdAx/xpUbC3CSrl5cR
MR5Bo2/JZ7bEusdF8aO+BBL44L4iVimqW06Sl3Gy+NVAU8gVELP4EkUktryz0Tuk
FTE2D833k9v3qHvldbK3Qnz1FOojYOy5JGWivdvc7wsFg3OrjhOgOzwLj5fQykU4
UkMlF5St7BoCe7luHXtPD8dtOR5H/XOfe/GkU4ibf8J/2dejhtMMOYPb+9BPIyvn
JF6Yijtfv7gLgt8aHbb+whEIebh080SK4sgplX1pLVhc/iNSH6xkfFRRRdcpSIZV
Th64LkDYVScjD7TNpfmL+XPImD4LtqCTnFx55Y/P9T9FM+hac3hcNTWfiAXTJl4U
ndpSDzxUMJh4IIwmjzbW79kP3G1LjtGs0E8BsnNEzjqihxIYOnJ4nB08SvcoeOga
0+n5IAZtICqIBPDOSUd8Y5W9FMwyvNH5SiNcOWKQ4ilPXrwK1n1E/2JJ28dKQDD7
Kf6nfTcOhjI+ZAs6cocgtLets6AstaM5ytMQ7ZrealfahqBm4LdYggZjPQqykjH5
SfXYiYv8DiumQxlTnhdfK4wUi16SN2EBF0DzcF+nMnVCXx9i7J3p/EHyPoBWi3xk
Lq3o0F18LX7xZlKMMMkQXeApKbIDq+2QJC407g9bEzaQ5xjaWBm/qEXSca75OCpD
OsiBIpHPAla3veunZJrBF5kM9WGpOnFfnAQWB594FLjZ/yLkXB/+Vg1pZOsnkGLq
mNNd7ejjzTdn2B84OQgGOIfXEHM5jYQUkuc9IvWkjcH/gVza9cCkd9PVZwrsYhXO
sfWs6l/z9xNsosfjbD3zcLbbiNx5cWpaoXMWQKM6CIGt+/eY0c9VE3lCUVVfJTz4
kdBOOdoV8AGFhAXcIbmdj1ma6Y/+C6QQGfZspgJiUeQ6+Z0p6REeHL/sLcuYXT+0
uldT5j6Lu3o3tcx6eXpfbk2kKxCuYmn8w1+961n4gRvnwVY4Zk/JiheO4HJaY25S
9Dn850Rw4wmvkkW0+N7Yh9Nah3kTP/rkjENkDGP+I/QCOG05hQyHPa/OqAxG8wxY
JpHnUETfPWrIU6tC8WzmUdSGgBNTNrPyY55qfvWgg/AwSv3DatGI0fDuJCMLoah6
T1EhUXgPRE9S81Bp/7OMhpQ36hnHD+L7LvUs2eB/eYrm9nNc1o+PZnRs6lFeQD6L
kEZHJtwQyDWdiIMN15ziJgw8jDv11XCAXvgDzOg7OPs1lcHiowSxYqaEr0VuyiXa
pxkGLVkVyupTeQbt7dkzqJ16V1hAU0pwrD67LwXiqVQcwPke1SyDmwqCFkYVzOKQ
PxECqEM0VdvpCk+l/2yUCXMjgRRYTbkakd/7c9AdhLHkkDApp81IDyiwPXdi8zeL
AQmTdJZtY+50QESe5+AAqVHFkddvAVDLfRerg+asZOlWyBv+DiFfZs7YkhnowmuI
aoRWt88z5BHWnHnOAlhydRmvI3MKTcCtAUQhszJoj9ufCoohb5qSZm1r1iZzqnXZ
K1NRpO70Dx3WsvOK9Ipw3ohsLoE1YV9fZWF5TXlorm8u1nyHrHtt2sJawYaZYtyZ
RJ5nhSRyR2pafI3szq6sTQHz3KX+e90uaYrRJrcVxyNDsx3nP4XbhDYAGvrnUWFR
1grcJSe5ND4ILQq5GGyRK10iQY1XAY+lfcAlCa64pDvo3kQyhigBGbCwRgOCslGs
lXov/3zFNevWsDm9i/7VDEgoY+iRlG4hMFxCdAuRYV4AxuuZiRx6eU9TMkFf9tss
aepplzWEEqrvW8mSXVgEB/sdgwHqEQLxNbk8TdHkJ//QT49PxOuw4ZrcIuWGAUWG
uMXL9Fy8OhDgC/MAPz1+ozAoIiU4LBRuDMACdYEsMMiYKJtsq4y8ganCwlyD/oNi
iHgKd+njtErsF2fj3sOJ3PzBc9/2gqOqHvY5hJc7/dpf/KoMbXZkFV0SLcYpWyU1
r5/MU8/njpyNEpcGcbahJLIbOputoaRCtI5GuPpX3+msd6TNCYLC+mSQoyg4etmL
bJbOLGjrVYLR8ycomV2LS+zsUmcYa62cr7Rvd8FJzDADhZB2X5dR/FbvbVBNkQPy
cA4fF28pU/dW2KmzFuomZpeBbAovSA9irqXA1NnmxvAeWDzHk7lCPvqjgELJHNIb
RetM2q4cpx9+syGo+JmalWZNDM8QzWrfxi9GsXJ8okpTN5VTesQILGPq7Lg+IMJi
O6YBd4qi6OlP22CACcIoQNGEseqguBrt5xGr9oddG+eYYAKe4bvFH/PJRaQNuAsy
X4Vee4F4LTgnxukeCoFD48CWAHscQ+6Pm5UkWgntNNu5Ne6b59/JLyh6kn/tmSse
C999CYh6ndyfFFMSMPkyRVS4loW7JzOIr2AOKbkx/KQqOA9e9yYTYaIlyZmqwMVV
3v+cPL4aV3bBToAyGD7WeltBYTybxvzxtPOqh0602Veqxu3Kcr6v4ORBhFFWAXhl
pGv2C2TFItiCCRpYVUTEFY7wlXdvakb2erFnjNviBlBiubSQHDXNCOXYr43CJvu7
DzaghkFpciQvIcUjV+btJsnNlsBXskHDmFjVdE3Us13/bNuOYEj/K2dOgzq23zuy
rTQUiMqE7KjFsQHCZOK2O3N8f49v4K/gZidSAj5ZDXRPRxlNTNxo+AVhxcXjzT1Z
dCbzfV6KTmZYMeocmuD1SEBsu/Dt25vas1DDyToi51AVMIPVuquDC7GC6Zhob72f
ickCzjmGnAWjgMgxxdIW3qmbvWi+ATnCa6yRhYHKtkAkC39sydVmaNI0G/VwbzSZ
Y9G3CJhgZHkrXCe5zsogYy+J/4Wppw+zNG0ctE+GV7o8yc+rzS1TUC2RdUl348Jz
ga2QLo1CSQIgFSnKvnB7FX75WE+Po74ddNIAfv9stdP+H5P8emyVCR0UU87rbnuX
FinSBb0QEK2gp9HMUn8Cz1kf++FImtqSlkoKNcPTQblJSd2d+nYTk0EY1xN5y9ee
vvxN0dsDhrMHJrfaT1Q8xFRnel64j7z0SXAdYr8SrSeOC203EAU3LDU0iCxwIg3Q
q8jJI0H2oa5xLN0G+EdhmthX4D7X/bQf1bfgvLrHkkUNmbEEo/jyTCgGj2aePNBc
ZdjktvNrqe/LRQITs/b2bdAIi9o15BRXdzER2+NnsA6pg5ZHH9Itsc3u1GlJlpSE
6BaC4FOHSwhHxJrptt9N3gOtL4pK1hoLeU97+/fOuR3N1OvkJdmWfKwtAnq+FD4G
i5m2pu5Vc3YxAlk68Oew/pr+dV3ZKHTIiw8YYLoeFVS0nrYARxUNgNZzGoQMht4r
JNXbP0zb6t4T5VPQhSQeubTC/tcCzpU1CnhYBKkseDup4vjIgXsbfJ4yt8zWdLJh
IxVdEpgupfDp3H+puM+8CsXLClMSx4cv5ty3dnk0+IS/q/2dYyvPxiOCNDZW6KvM
UbyVWqiq/vwhqA+6wi3hFjfy3ElVf5AoTDf1N7/TNb75eX5maDiPspKkvIzdRjoh
6CMzHXfO44L+LdRTR8vB9u8JuRX6e3Hb0MtJhpvF/wjR2QjIZCXquCfGyJ/fcOyg
d3Ulb1zLSx6ESNYGbQ7XuFNH9hiuqi7SDRIA9cgvHwYS6uT9RfC8D383C8/SuCSz
kdQNk2rjHUmRMgSL+i0P65XqdnAeVHpvZXXCCMIGw7Jl3wW0Un1PgXYbSXz7xLpd
fBDIgPBxw6y6OgGuNBWY2V+ECB0/K7tYOINc4l5Cnl0u360ZIYBtZJ25dgg+uZUs
JF1qy5wmwUGbHIPTsNYn9xbv0/sBzwuzlhs9obobxFB19nU4BWE1SA53Trnd4NLX
4+SMo/1/UYBsWC8dPI67ObYrQR9kYnsKlJ40r1HCrYNzkPiS3o8o/xp5P9gyfkF5
8COIMFJXv0qzUvrBGl/Ik6WO+4KP4GpPN4PkDi+gtnla8L32DhvNtdFNmLPWpYmU
Lf0BnDU+GG+qAWOP1WdK1YQlZVWcLfftzm109Mw7Ca+M5i2/M06V+sWwFl790XFM
ABJxIR+Xc6w1XOon0aNc6qlTqDAyqPk4LWB0t6897psJ7PxGIJhEC5ddNC3XmVbJ
tcVNDgmVqb+0Z5DTBM654jYhVIU7/TCxmk3Dlz1bpyK44ChYC6jvVTWJVxME7daN
HUu4xN3wRjgx46jjrqN+SUVT8LNhl4sZWC9+iWAEw1fgCfsusRtqvlHLw9/n7J2V
COAXZ2LFn1WMBK6KZl+7BKWCEMDMVmmcQNTdv2AZ4XG8N0dCoJYyItxu/zoqCmeb
HY/n0fwAAMIjaPnmTZ3j8mv6k76G0lBNpP62u9qUuLW6TlJrZ3VIG8q9uxjMMUyZ
9q1MXB0/qyWIgjAs8QcMFFTIzUeBbE+TfTOKxovU3erfqfrk6WR/SS2ols5uenM8
v1ALh4NYiUxrJlWupN9ZpPKQMuEIGQGLRRQeDReKqP5NE59XCqAmb+9IcPtPcLRX
xXwsimWFX95L+qSSTSsc+6qWfXz0atIXgRwwir7lcV4WJtbDVNJLqVamqjG3/X7I
UA/TPetHZWuhGyA1+i9VR9+ZFAoXDs9nXEvlJGZzCo1ct/5kLzwCPhZFW85EmsIe
yVb3W+iyyPuoeK3BJRXFJpoENUh9rDW0Gp7bxln39e8n9y+p7vb4GgR4YAn0Eq/N
sRCXMu29nqi4hoC7IbdmljcJ2XwwGx+Pm28J51IjreKVq5HSlgrEuAmhX/kFuI0W
w0JwZMM/VNkBfAQU0c0NCt9PdHj+Y7mmsxDVmBb3qrDSP1U6q7Jtw9AM+rzwRVOz
xATdyd89H9ZriepZ8SbF7Lno1ngPQYQsy2OdWaDICuX/Wuns4I/uD863snvrkNPA
PJKC4TPwgkp8Y9Q9ky1mI26NdGvgS0D1bmBJsQWzxmVclx9MHf6Iai4RDe5RtjwE
xHxPrMc3E7HQkaQ9QYvhPECoxrBDseaf4PLvEC9LmMXliG04p3qwrAGpjSm5TN4P
gZNqYV+ypLxVwL2wuxQ1vFGMrZVPnLLvFhATFIRvg4mXz5iLPCWQrFbjGaSVrtKb
GyPcSUpLB1RBXnlAoa+AW5TGlix6IC95GAVNwIu2mpOrcqxhzhnZYmV4AftqdbOM
E2JaOkIB1zTKeSAs8ha2V3HMWL4K4SinbBsqRJgKRDl1Nz1nnD98VRNq93EyBM4b
IDEFjlTpzXxlExu1n+VEMX/cBaa6/VfLULS2kg1PvXkdfVZRGClfQIlfAyYOMFQ9
H6sBEi4E75pXDn6NQGSA3PzSfilsQ0UhBJYpQzJpuqtCHefg88OcWxtgLBIGf2B8
PN/A6iXp24/S10CJ2k1dps1itsF4EJgVsuS9GU56dohWy157P9NIyfuZEkCtwJVe
KGKIku3u8hBCC2tbqyxaNlUjhpWzf9ODHpKlPa3pooQwNgA9y8zSSZYswhCgab2T
4HTUdz8yQHe6FgC2WyvM47BqKl56FE+Abmozhqs/2N/bMMHYF0cWonFDwYPTz2tH
PZuyZtNPr6S1aertGsY98g3sVneu4xzgS8HBiKf1DgYzI58xJcQS1sn26fID3FUK
/KDF1oTv4H12VLuxU7BCS1Y4liqoGW++W6u6AVrg3DtgBhCwhtNQR88IsOp86iQs
qWizENasoHjfw6//yod8nyk/y8/FvGMrAVhrloB5PZqXjajpoZHGTkxv3crAw/yr
eBw85voXtLHw8/ajex/VlOlaWxDhAb0OZXlIevbEfVSe2/RI66OrcufYOqBQEpQA
wlaI0jwCYB5YGM9xyT+DSJ/xYd5glVin7vfrhhR9LG70ONjwzu2ls+D4tbgh98+S
EaPEYyBIZRy7gVWeq3hLje3IFDbmmhJDa1+MEfvzdocRXSCMBOwCohUJ5jy1QCFk
OMgf+zwoVDAGQmLnXRCDW37S4mTuCox36THsdnaYmYx0UCcSCI8dh4i+zvupi/cs
xYdNv7JyebfjpNw61SWxYhu1kHTGx4qPvt0X4iglSrcr15cZejbXZPyIxPl3P3DY
lICvVCuBaLfZDN5uEkBTIqRjYk6LBBWz0yn7Mt46TRWU0SEYUCJzm1iJjXbRHuRQ
X2ZQrIRlMAItLcXNgDVvw/ZnkL129ka4FPTHi67bupYn8y5Ck7wthd1UhmzVN7Vi
3fBtRA03bQVoOEqdoRKfql9b+qoI98Grt8qyB6CfFum9IHZLjpIJBbd12Yvu2JWx
TLRCtU7PHVFpaR/CGDm105v8fsjA82qTZ0dj/rCBv6OAMLtcx8heE4K4X6U0SKLw
/jc86VIheJCKNFy3wJGD5X0C4z7a4zaUPr7ZfLKeE2GVvXy+0K9uqb/ZeSGZJ12x
W1QHp5SfaJ468oG1/Ih8BLg26c/u2O5NsfYKTXCTwh/lYFxPhhean35Cxh5uDj8n
1HJrvOmMhlaZaFt4VnKH1XDdoOKxgA2k5BfB4pKazNMaaY5rVLBPpAv4ek1PFNLh
MKEq1sv5sF7MavOpfvomvQim5hKEg3SuDNfldrPKxROFFeDf0epDqAHi3MpIdKXi
RtcnaoFQUlCWmnRndrKYg/FLtXmpEwuRi4mayTNEd37IvtprNiGNGbdI6NY+xCd4
w+zEtSyuV/1yZT0QIlUJ8BEQzWpF+YZwmqtzDCfz1IYFS4SthjX3tAi9xpCNlGfI
Ogm22Rjm6hXQOB8y5cPkMNwj6AYlw7lMB0gyY16z0KQQTN2dEQB+DCZi9w7GJ+cF
ncTwcyQB2s3nzq0ZJ2mkyAu6XQ7mJX+8ImO1bffZn+nUx/76xzFB2vEX5p245TFx
arTIfkM2nKUKZzT59nYLpSwIJki7+tzCMilw/SDcLqexxta4shSnNbpZ2bZXhGoa
3X4ufOzUYc4X/GIbHoqYoDf+4TtRWln3+B/6ZWaII7+GD0mmF0y9po849Ku6XpVG
4NNvpnABhjEfWX1sZbEz7MLN2jKiF4SA9NGb0ZGZS9N54+RjywaktNjf4+0pglPd
fmjYpZ+hPqdkali4I8D+SqNx9I6WLl3JQTT+MerdH1YezP+QdyIchqcYImYNKDhd
d7hRg+PZJRKRUzSn0GO1tNwanurq+exaU57SSH+DShvy+x/a9ZALAYHv68gGhql3
QsxrOrARj3n2TsOUPenNBPNqFc5KQ+KqTbYwhxychhY0lHQ5IQ+vKFeYGE7d0ZkM
Vt+odMCGneXIYHo9FHn4dr4WZ97rsFsxl2nAQ+d2uSbPlv1J02rhI9UP5o7CNLCr
E7wDygt8/wqnpUWO+mudMTk9Q3xuIMr5mf2jS0uPLjeFuhisasWcI/vwdXLOFNvf
6Ekgn7tKc5mlKWn7ySS8HV7ncvvnP6U77VKdfUo5B9KGqxbmIYn5D5fWoeZcj0Y0
N3YTnqwy8yQvsb1vSkJpcvTWwDqpp05lnojSurG1LaIk73tlCXMrNzqkmgp9hrlR
AxJVLCORQlxGMoalazxVVutvj7+57tNx9texEInjUHcZPPpoM3HSB42cIc3sAW3F
iz0Mjm7aVTkyDtBD72CfFZwYhbpCRCpGFS1o2eqP9XxzYOSaEwYRJ5X3Z7Z4q+Tj
22f56J6yk0TabsVFEli8oa6s40mVJtK2u49ALHmjXr9NfejtMG5f3NNrstydG6h9
BTnlQWRK7FPGnLhRqN0JP/MG1oTYF/drx/Z2XyKVx2HBFm1lK6Cg2Bfrox3Sqcfd
cfnHxI/CnzbN0Np9qGMUIC7MAvUOUmIMT1j6D97q8MPwNxJlXojRZ1bJfjyJ+Hl9
oaTgCM35tB9zEPQKogi1PlmH38ivXhK1wagCGMDn6zvkgJxcmmvCNgfIZpqu8YBX
Ysv6ENCObMy1IiDbGPJYq0r4ugm9vnerS1JyC8dUVNUX14Td3LDyg7eYYGFzF6Ga
6ORP7CbH5WgQjx+nvF2qurWSYrK1RSnXQL/Fcujz2SyrwF8VX38aLqZwn9FyHvzy
afOxtgs41lS+6OtIe9RENPssCs3SB0LBCwlhlqmaBpzFXnkgRezhT/jWM0hsnj+9
G2VbS+Tzj7Ab0oxLIlMcIx/YkxeX8jALYPpEyXRF9itErohltAGopv7c88P3Ve2Q
FvO3OBdVPcCKB4w6rDG23nQlobwNXNS4cptH8juT8dyKHrbqtGQN0musES6kLzHa
lv4dgD4HZRYJfUAqjwkSRjyKhbmbpEPKy7FRPVT2qXjbVqT/RbumGfY+IAawIT0u
j+s+UxuwUeSNEoaEpo8K0D1cHhY2gEo9FEY3n6Gu9l8Xx49n2T//6Wf6UHUIUxat
8DsXOL1ZYPzzGd3PNy1lnvHoViU7LstAr8m3V8DkBZHXPOe5R9wKVNE8mW0kAcio
45p+vpQbaSD8dp9BBx4LFUsH2cBlv7PyNxbMcBYNLVM5319IpyD/psCv0jKSk1ap
83DuHWi2FdzlU40/ce3sX6kfih2b1fWBtmta9S2vMIVGWfPIZ9Bvs7k6jbg+k9rO
KLsDr3Og7PHucUyLMA6GAJtZPzVN0cnPtugDSQO7NQeOIh7CH/CHbaq/YXMrCNYy
hLkegp2OVGvND6aBN+D9ZS6L4lNtHvUnK902oNHlW1TuYc7zSm+FncllrvMSJWOk
NaNTMCcM0wSPB2iU+rjnsKtW+VJwO8VaEl0Nny+OudluYaXGZ9tD5Y5NGSe7ETMc
3fP7NOFlOJ+txNJtj2C3LcdMkY5uO/1RDxPH1dIvqBqBH6HmXAexd7GShVyOr7lO
wXXeLe9jAeH269b3qyCcwpMhDTEa2mD1LmHhjFZUrz6Sq5rT7QueZckwlW2HGHDT
QqMjilHHaNMsB1v/eMpAuGEuIg6hzJFhNveJclCL7wHRpZ6erAxXvCY9PKTz8tLd
5T7/IUILVeTG++ysXDclvCH9/6uteDEfqxStD8Y7byqgV7mRYMwjvY4JCXt4U8+2
2HTKOaAMv3yCZKGXcE+sFqZmG4ocvW2ZHHf/z3MFVbClfW8O1QJir5wn8m4XPrp7
Hs5PLf5fQt4UVTbaPr66lqADWZa18k3pF2TPMKdLJpbfgnayzrWnr9BMtWg0yNLo
Cn0e99ZhOq2GP8h5JJfnp/0XbNyJg3/Ak2v4jVyxwwfE1lbuUveVgsIxvbQ/gYzE
jgtqv3mY4JKJvhdsL6q2IW0f64KJUmfdblCvEMbfvCZ5jwM374e/9W+jwQORTuYm
OnTIfKYtDqijOnoPEy/qdi4EqjXF/binDOuRdYvCkFPTUxCF/00H6C0VxcbR8ELV
WJvFbvDRT6ARZJaGJDrEbjuetB92fithy3O+MkD+2LbFtOSZz3JIR9zCTcxK7oZe
LwIJztIVj4RRoexS3icL8MqSSb8CAmRAmQv46lfWL7G0DV87u60GXnJ9diaugzQ1
iifPFXgZqzGd5t0Gx/MPvvFGZx7v7P6TEFZEtRaYPReqwhorPkb/v4GySHJXk5uQ
/sOm7IwVXfuzfPu7wHEbJ4ymwtUgOHyws0ii/uZgTynH6/N4yay99++vvialEE+Y
h2VSK8x2rLPVghUKClCNnlAFrSSw01MzRvKQ2SIoUp4QwgAoKbXPy2r1lJyYqfQa
+QK0IJE13nP/KLV1Wb/voywYIC8hInL0tsaMUob3GQVnqHng+vWTUj3dIwA66iFF
+8g+yQi7wIih0ZO2jZ9HBRRyEjnuTien92jcKw5VmEKY/zVLMmmUF3fWWTRVpD/2
gaeMVvBcq+vXhgf3BUVFP+ygsiPvCdcw62I5uWVq4G+wwB72cXMky5Z08Qsc1dNj
616SM83mkYBOnOdmydYIOgT99Au8QVDV33WtTK7WXvyHNC3ZndgecG728ctjBRs7
JR0LZkhgV/1KadccOwUkg5xv03EJ/fTvfvGqSiACl39frcgWwnxq6Ek9IDjPUTDt
se+Xetc52GlGHJV4LdiMO57B5PZ2fvA2OY3SeUZUJ6FS9jh1XJZ5fkJoMzDDDMNx
TN4VzaId1AbTSpQOjMEFoB6Ot1Cfo7P9IqLJHqVL6pkhx79pHacwDkhW8X77sCA0
Hg3VhiesSi/m5NyntwlOifVU8AZPj2t5RNCoI5BFSS0GpL5CJ79VtwKdXPCxBT+S
HygWIg32X8ZLQ4LygCoaMRLrN/pElB1k5bo0SffKFwq3r4ZmE2yMNcD4fOJ3hmoI
RVS9IOMAWawHPwahvhxsBoVtWnN2u5VLqiXZbXBKsaXBv+XkNXnvMq55dUkYhVUc
LZiiS8jw8OS3M+cDxqTdaopOC4w2Drh2vevnF6SNQY25fHFaoGcmGJRyt8vtflKS
nxJLwKL+vNBTBLc5iIzmv+bVILGGHcpMJmnxFWp9SvSjx8IEDOaG0Xe9tGrEmGxw
SYV04C1PasQa9VuUuF0iF/aIpRq5P2cRz+kpmt3ppOLMfTnv780+QG3bLrcsipxA
M88uhgd448Mv8Cilg5GuODX+byoJJH1zPcssXwXCrHOuBd9pSskNtuEt3wEUKOKa
bkf0zjoYLPcctzmO1G8iS48qMXThyKWnmip8KAiK5oJdsP6fNnoz4ds2LEqk+jSF
kyf4iJCF7w/wyP0ByuDoUrmCMT3us6nTpiUMfTNB5yIJcCPO2X9hhPq/i/REYAHq
Z5ki4iS3+zfC0vk5k9mImymlOmwtuZINBOnPboin8AApDodo2Etxli3EWFo6onDD
aSpAErA1PkW7wwf/fP66nKcc6qS/wphN5u4FKX1qrd4iTa1WUcew7BCq0ZnkQgSC
KPeqxUUWHqZQGdHzDYG+YANl+HRjZrB4JNJcPzYVvpzdykfRPdYLLEB598QYt2X6
i6rMie0q5O8WxJzw5P/B0OF2Zkh1TvZobMxVFD8lPIUDl+C84vquOVzKDUNLx8n8
STaqlNQJwdd51WOCnTDi2VS7dOrCGaNO0VQ3DZYyKHi4Yu40yvJxpOaJQiuBRyTG
crwLFM46T0V5VAmyJ3en+m8u2kgWKHbgzRzSUTZrcVvuSVMAxh4w1e3Yi8gl+7BM
Uxgg2fBnNK5DymAlQ/qErg53yTrQun4ckOJemLF/6xQ+r2wMU9L65vhLqSzzUFiC
ND28Sw04fdEk/+1XVlqYfPiacKveA/GdAOY58GTOCg4kBntVTWXySNLRYg7ezYkQ
zpGmhK4RabNG5DGhUFqLT0ZnSe8f7gf1ziylp3bvCmYKe9P3CyG9XIEHOVtEs94t
RqrQQzDBcDuG157/Aib0KCsYr9gy+02fLwCLOuMz0Uth/Xd0C/cOVWF4zdMhthXN
T3OoPlshNWcmRYpZBMCWf7nVGfbAcJlw5GZznY/w/OQNFkiWLlyd9hE1f2lpeYM2
WIYqfgyXTrR7fj/qRPNJsQcxb60Ma3983IpS7IxSq/eTYsTxaQy4v9dv8Tjnbkym
M6E+A1BlSjQsBFSHgQ0T9iaXyRtfwW0SsNm7CTEbbvjD60SYnGNwgJazq/UfSwph
U1Y78+7704GHU4dO/uk8nfdQR/GDW7G70WZ5wbQFWE9IMMbbb6zWYnc/wfffGW7c
UXxSM5+1Ha+n+foopp5JcyCOttc9VPJjOygDjc3IgCtU1+PBQ0qPaLl9jp2dRl8x
3PGGqoKlmtgh1tH3BpcrHDzhplfXNJCpBf02Mo9mqxuu52wl1D2QRuGgxT26IgCe
wZpXzM6QWw30ScrD30uJ4k/jWMTYA+sXgliL0jESNkfHIE/Ml4XOWAcMQHNZSRGa
LlMdo9AO5/U0Qecwy3m7l7KyKISoqQWy2+GFxkRk7JJysD3L4ykcviEv6pnRGD9U
fonMlMrqsyibeLZeZMRVIiRwsjXJC1/ujCMD6M9dXdBjg9gQr/WM8om9RFkiiu1f
IPe8macHgZ/7rdpiYfsgIfH6MbpCwiyc6SKC3xzNUv7J+jKVWgILybvQQ6BIIsQG
/sEFRgRSo+dzGX4Vt5yPpIu++GnvJ2I2EF/uWEb2Z4Z2UHKUH0tV6IMK8kktvDxD
mywM1SSCSrJD7eNIKVYjisladSXNk2djCJTVqn2bZjgvlufNeLnpnqR6VI+UmkUq
bPsR+DBJdLi7+7yFYXCln8bU/+CZBoAQoJGnNOFFw0tZwdAof+/WODZ076fX1NtY
OpIfy8e35PlXVGOfhHhRHjDDYiMg7WZdcfbeiRHSQ0SrKME710lbtohNygWo567u
cjdHF7zdS/ClZQJoYDopUQ7vSNQvUUJbx5iMEQ4K6iiF5R1t2SC+YxdIcydAEbEQ
rquBAHaTDpLPdsH1wUWySY4tTzvkTZMVXlqGNzPqYFYmG/lyTa5anQvhd+nPg0o+
D1JbQLWQJ5OzYzuO/duhMyEbarFggPUBgN7h+KEwm0e1hCjio1xrtrT86lKe0kH8
FXnzgolGun/hrjQzOcUaU87b5sqJaGgNct97a8vewhEKSsRSBVXEcfsoh61k5sKw
hd1HiGXEpT8NP8ITKhyxEbc3j2jTJItLTL8BYQ2F5UrPutsw+/3HIdeSM0WCmuGz
qzOd1Zw6JMXw3CuDOkk5C9+EC7p+toAPxwRCPymr558q1wyk98MT2ErJsggLeNDU
ji2zUaE4N5CCD7Pon44Z+ULqgWR2HxGlCkAZZkW86rkdkRY4d3HH+Wru1z+Bb4db
LmIpNbuxlbx0wzaNsW2UlLz+REe1J+l+CbH2kMoNpyrifGhKrsc5P831vG71Avff
9pnKE4jde+xnDEG/ObewRYN0V9oCOYO+DKCa1ZSSb1CcDgtyaH6gAg6GN/dsGXs1
auj3aJfIP1+cmIOaA6yfTVccV9jIdu0HX5C3/cKv6Q/HER5ad78KvO+rFjuv08K5
XcF+VvxpFZD/HfH5tGNxZHCfI5dJ3FVy1hqlzD7rQzQrFcF5y24ZHkUv3hkq/BGV
s1m1W7TpYAXGjuPd6QaT2HkTJnl8hHwcj5V8kzGxDWGinR6I+H80PAId3UcVjBNk
tXfyeYaFvYORo7axuD+atGDZRoM4KBeOWZM8TQ86lEMIMr4ki1eicOQa3W7PuDAL
AtjqyOxT0QZCG48Fq2KujwWsctpVYJCBJXj31AbZw/n/osJJcihpSGIa2HwTiTpx
UVe193iZ4u0IiYPuT1flDE5ybRL+2133fUCGn7tEeLRi9xkK5CVyrjZlel60X8RB
J1ZF8V4Mn1hdl+N0rmWhSqqdOKM7Trilb7qUtvPgDHLuVV0UOBSn4TrRe0KzuCqe
ZrZWLNWj/qOig6YAcDhzPFyhOOcHGvc689VBqGnwoegFFVnmvCAEiblEwojXrw2Y
WOTbeHwolXBDtyBNrgSbcTCEmVbh1dji7o2i/swLkZe7gy+FyEBn8TSvyyNoxRKa
isDxYMDXaxp3+9tgAFKidfZYUtGk7npEXpTZoRjc0EYekeAOJTeQOFaX57LsIMeH
RmPQAxWGqCW+vCF5nKX+gI6MJp9oGcVZbfj2ju0RETd4Jql1/tXESvCPwrNMgti7
RMjj4MGaHnWyW92x/Bw0cnVXUF/W4EnPdQkE+YtlW8n1vw6RWdYWKctGWh0bZP1D
2vNCph15/WXLTtmmsqeuprdJeeQ9MF/UT1Kr2+Yaqzy1jvoBdFs5xLzpOx9MyGPl
IoAqjJzsnMM705YITX1ENtSF0mLY8NnYTJmAq1186n8Xo/4PRF8N1bwi7b8UkW7w
qSk4ai4yp/82lrdZ86tDlt65q+N72Uzpw9o6Fw4bHy4aH5YMUe+IKg3P2kwIH2z2
EPvrotrCeu2ER2ZsAxbvGG4TyjutxGi1CD5M7SIA7NJBdXWXWRacLdPmqghRvGH4
IHjzTNJ1sVq2e69WOe3fb8yaJbtDVtHUQL/ayrVHy0TmmZCPSeCQO+LITzxgA9Sz
elNxfs5hMe4UBl7/BvkuiHAp7fa7OeahUflImLpyStWWfNG74bCwE6ehWdqgX2dN
PgiKKYRjKZ7WvFOKDaNkiRcNfd7/Cz91wTgQhx7A3gfA46zUwRbg5Qq/wtgHR/5l
fy/J+yaia3ZFONGiPPaGywpnhqCBX8O3JAVhlpMVJbvFaj7O3eDYDrKJiqv1InwC
KZdh6JN07faI+pNUemBc46P1PlJ3H8ymBu4uuuzzthaLPhzyHWvNj/mcP98KXy9U
cQXU9nLdSwYG/no5MMKU8pSvPQm+Zen7HGMKk0/eWlJOwbmh8I076FYFTvGH/wlw
RbeHagVGGfIc5QOCXWsqDKOHJpY9gdYYmQ9FLaiWVZ55wRX6xZMBjWeWibBZQCDM
JG4BD6ZzI/oa1Di7O0omCCjd/1Qa7G9l8jj1vroxnJaaibucS1BOToB/wfdMGDUx
KT3G7YBiC3P4aRXxMhbaWzX9kadlR7bhw6htYInIKbJT8PPBehpaJJaA7SF8urZQ
B5MYjgji3jdwYsKMNOaNGvTVX8Xo6DdH+6ubaXzIL6/SkoqnIdFjyF0JIzvKYsTa
z36wBerO5hvD0eTOXJkL/yS5fIIhwrK3Tj8uURUr8UcEAnil9a9tMghXK9qx29aS
l+UujuOLmNWKo61nixJqbTKcxvr4kZTbTusRvx7k1d1euRzB2SDRP/eHhOSyQpDA
3Bzu4+dof38acSw2GwqD+reblo0YwMO4QXiMdi3XQuubiNvohj7eNZ5xIMXcFqRs
08ljWH7blBjYMBopLiImBPGDXGWiIKjf4K9ganuBtAErFXPqdL5he1NiqczneBav
Yl8TwTRfAKQJBZcWEd1hvTwhOUrydMg8p0HzHj+SreF6aHVXOHX+542MSAibtLfn
RgTXNbkYH16jpnxe7koeC04A2g8NMLlurW70fDMDC4NjqZY8M9FcjzIrrRL3s0Cm
0nmbsNZY97H/HAUeHB48pRVHB71CjIQUXnZJVJWfV319zCoiX+6driIeWxEGMNK2
KgIW1jHWrUjg24ahIFW3XanDDHblNwNXXwiqqFFpb/WKrVoOKFRpIV6X/MxOKYVQ
xfb9oxNictNvcoeeiGrHNrrsDzytVZFPTlFQLOV0CgJyPl0WbHS7iiuMrYRL0grl
RLMM+t9pHr5C/QnzKsTugphkFeZkR/7JAMB4r05nNCFoln9ckMXnSTOjnmpTqpEc
kIVBT0kmENiOep6XplI/b3eeFqF136KVFYMPJLqPIF5fhl2VxPaFwMBsJUtzojqN
vW3yUFUtEbjSo3Lz5jzfvEQyJi1i6dN+IvFQKcgEMlAjK8OD8cNV8tHZOP0uDrWg
YDlnAQE4R37N3rjNZoB1y+0yLTZ1kjbjWtAyg3q3OQPl5dAAOXdSsL+u9gaNItcl
Q8vGi288399xwZzmu26H+Izj9oImDtPNlHBedacQRhIbmObVAdKu2IqTo3CxHvIZ
2ZGrYL40wyBPrXzx3jOuOr90DvldB+quQqAFr9kuemIp9RSABk8TTEktmHwNyaC4
TtW5G08sNiOKUfmCysWjXlb0axOR/5OZQpY5XXALwejTGEC4FA+Iapsq7fU3nHfW
veCcr4QvnySrha/vF53LnQYkCtLjhX6X9lRX0jh5tepz7xg9JoPqQIkjE45kENXK
+2oY2wWPLlgNU5MPYVBQVstORTm2zC4dCYSMIPQ2utzPaq2PilyAKDR44TbtP75a
X/CNLoF59OBlNVa8v6NZrGQhjNb4WxF7EEsUvP4VG0nuzpgP0+mdcZSWQ4mkdK3W
FSuowA+y2W0DVut3LLPlawEUcl7+pY0ersWIuDsp2Q3wm44QDNzShnq5XL+RkWYU
zjKxezhWWUPaf/RIy7pnIwiDvIq0ClV80IHc6EOpXYDlN+oqTuPiGkGaQX2pB257
Yg1jK7zUYWtr0SNgZjRD9YF7ypW7slJc7qWkDxMUGPcGb9ChCKedykM4gT/WbXUH
G6UwTRG939cWTuk3IXWFYk4yrLLMAKxJl9QsIKNJPCKDiVgjTxw9sQ+nf3VkbRAZ
ZMoFiUb//32X3QU4Oyuf9ldKXgocP4oIo7kM6W5AtGEhtmkVLufjkbaBd6Y7xzaK
R5mD7Vb1UcmUtXbKriq0YvvWBZ0LIvetWtbtY56dytSYuCTCM47eiPh8qQClfaqs
bEk6g7JcHhHrrmEI+NH9K1OHYI6g0zsMYlcvYEBamN7dHyVcCNpNBE77/iC+8LP3
zDvtKkq0q7goWhocCYGVPTh0xOcc88iEslJTAPCoN90MydyWQ3oOgQp/HDgiUfc1
WFqq2ZajnvQMDEJs9DIKu7kayAB5CQ9N6C/o+OVWRiYjehCjAAHlKFSGJ3J4pcMV
rWYPHp43bCWUBuEcZDFQ6GWpB2jNr9YqTkrK4zSLHlEeo/uOyzMEMl8O0EdE+5mX
K3R+J+QE28TEtjLGtRWKUsHfcZ9JPbeLIN2JGOus9xgqna77ZVDQxtBuPNEJ6TXL
MlrrSvMKUiI+64wfRfUHbaZ0nhCF0MAL8iROJSHGgAHJiOfSceBjDWyBkN9iUhJG
oDibhfSutAEN4HBfBnQJqOBczwTZvDRyLY5hcSiO/F1sS++GmFqDQR4lTgPmiAuE
doP/38tN7pxSJh0fR/Ks3ECSos78YNhkcyQ53VJmxAGBoIxJgo9Ff+qntT534l95
WinGYMg+8VE4MxxKLuxp4hxq0zwAQEt5YkrWl1Had6NX03tm1RGN6a2VALUxsqah
1q8XUeojOBMKRF44S1ZQv92Ajc6x2ziwCNQ0V0ZASBhytizHZk03DLkUaQHb39C+
EWxZgXJl8SiYxDNuuoRpClv9xD5fXSipriuw+VT9+JyxptKIpG5fsj6WLPchC+K0
Co18MLluNOO+NVbInO5n09S9kuX6omVEuqts+u04nPoBjfHmBiyzPSOEtHZe2Pnd
kAx20CTnAV2F25pP52+AoLozmE2il1eGLSISMbDSPh1EM71y7/k6QIxTkyCL1bnK
0harhk2DyebakHNY8WBKWzMxVNrbdKmB706tVa54231vu8TqsK/PTNjYdzJyn4vW
ecwRRo7jRz4KoA2GlwyvgB378TBAGrsszRAcHNY1M/YNr566WpZZchmgmyWNni9I
tiz7Myu32ix7FqlHCNY/Y2Cai2FePZDTzPUr76Ai60OdH2E+egoubIwQTAwl4JOG
Q84ce7/qftqQZ+jvLxfvoQ==
`protect end_protected