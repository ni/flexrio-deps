`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Jm2uGAVYfY7w9Y5qKstopObZuZAEY3b/Io3MSEcWLhjjnKulVhCBBYAEQrAzzGsT
vMbffkdZgjdXQUg8jOLJXSHZ0Dgbnob2vlppjZs3bgyHCF7MoJ35E+LOsaLimUA7
hlqStcK49hR1hdeBPr/OwfT3UeVrRtQyq0eJXQ1UksinX1G9Pz3/CmcGfTZ/C72x
p9icpt0bkY4/1I4GBvNCsA6FFKH947JqH27OPACiQQRW/K7JToQn+1uhWr3LA1od
lbVrWu8PdZi7zW9gK3jiW5GaPjwbYQGqeGFs3bTKBILjb7sYHxfxw7eDLVMAIu5D
W+OTIN4JiHiE1gCnNEvkSQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="pm+c2fYA/4JT1uhlJGVUubML8hZi8lME4xPobg/m8uM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
nBaXksR//iZ9fraC7WMJWWSrjqRXHxmM1Y0+KKN3b10NElDzVNMlR76DLrcnamFd
2n7uzsxWqhhJR5LBl98SXO3Y90J6BMbw+OBG/MFM/zUulxh2Si5YK5G9GCrG9gvZ
5JomxuZFDu9CzlWGTuRUt6FsE4Lr6sOL1P+hraQDpMk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="M8TXDiNa0BVMX1P60yIvW2WA9jKGGy8GtbuPknDnC9I="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 50560 )
`protect data_block
/5TNZvs8Nu0G+mfp7M8H+iVAGG3Mh5DYZ0Gn3rRNhV8b5CcJKgjQajrRoGl/gSxp
rBAhtT8Vd5eelHgtvBjpvFBA/EBUrRH6CG6pqRt9r2qUDt4UernbZbxC3BC14KYF
gLiaAkKLdB6NWFZG4rx6ag96XC/hAJnVVdmIEEnyW16bX3DCU08sNySu0qtMffQS
yPlI2cGLyGuQw4rTxOhHDDWMKN/IZxVWwSwyDSMa0W3/BZtNhzzSdwQAKK99Qb37
cilFgINo4L3S+bssU2PEGOZCKVszuEI8KdwMBDdD2k3y/8eSobKQlZGrgKeQq9/3
YEm8ULFDg/nqHGNjOacmEsMco6SylaW7zcj9w5ljJS9796SdRvCd/MstwaF8B0Ii
5hlusOW5G1NNhRLguv0gWhB15ckQH8BKApCYt+hhGEdbYaYyuiBVur62/+pDaeUo
UX1wS4e5DlHTdFCzKBsxYVa/dZh3IkNjQfxsJCm6xUA90RdueifL+hEhF43UVFXO
5fMc8bvNyrwnnZsWWAHOsgV0RsnPLacBhMNb1YOZv6x2GNntiUrxkhbD/yPRiQLg
j0YeLQ0nyzmaQXkV7/wmwXXbbWgpylt444hKiQuyk9hhU0N9AZOqv7tpt9gDExjI
VZ/3gQPF0RnMR5QCoUHqtT85CP0HBnQylE+ti2g/x25osqIdnY2jF0l5IhESYzFm
e9fzpTbqJUsiNWXHKiJza+i0eAcJLNoc0xfLPvIZk4Vn37CxkeqYV8Ft6Mor/2Iq
ICuNKEMMnL3i8cLiLzkfCtuh0ecmJjBxsdegJRlbbkW/HuoYir6I9W0k4Rjrx65w
hKRl7RmVBy8hZSgluvY2lq2NmeL71rQTWlD8JHhwHrpYiP413G2ZzVMPfBs1YAhx
fdLAeLyXNN3M+LKSWaGrU9yYJNPe3iYARBgIjBcNZisvjYfs6dzXJ4np57Ul2ros
4/THIh7vOhmvg5Vs2lPnDwQmkhp6xjqcC7jy+3e0OFXX69NziXabaPik5/nJWilu
hp9PpOQZL2JSoK/Wj4veqajD7kzgQzMTOBlkZbsL5LVj+Kgo4ezN3i2WUVc8zF+8
bj0bbCBx1+/j0MiL7l69BgKJ4CWkxZsHerfcEStta5h6lwq21D7SLjJRuiNSFMNq
2Gl1avWohXq2IPdmi3lUgVy366ffSYjTYbSpxwXF69TmpQFHpGMxlzu7t08hOWW4
4MguZ9TdwXC0x7PYS/Rn6CKOqjf5K1/1IMS58tJ69YkKnWQBLyai0WNDcndOCNYm
EtJVqCJ+1iDNz5QMpCv6k5Ke8Luf9f1GhWvdAGgVgg0MsJKWlHjJyuL73kPT2Fjd
S++9jZ4etZ0zSW/GF08Vu77DbfozjexjgIKdt7Fz50ahvYEOCWQr/zxsrQTCR0Av
OtzvOa/jSlctIe23nWm8M4BKrTBYysq2/gJb6zjE29PqaHCOJLkaFdDfIN6h3IF6
28bg4KHUfoBor5XxQ99kkZGtes/pMxrFKWyqzwEK7axv8OXT/hZ3okd2JAv2jRGl
WfM8M15Vm6FTRdAp1IG1dMovcuL3c1V7td2Ec/nMRj1xgpK2kxHuZfwAVAzPRM3j
ekXGLUxZmKqhN3oBGhm20cN10bb4DtyNAkYDfKqjMCh0SlWvo9cl2vR0tVJOe4kB
PaSrQICbpCihexZ1uroq0VsgMJNjngs+ODrDQGVTisL91fq1HIU42ZtINRyX3E+l
CT18p372N2XjmSKMlBO/igu8I4ypIJIBicqA6jJ6Qtyu6eMHaCHGXOm/jxRiIKco
o5cgy+cCOBRxCshw7bAfOB8wErZyjPQIMRoou6Z9EGygTfLW5ngHRTWVafvFiX+q
d/avy4hId4B2BDF4V2HQlLLyEk8a81gEgXpCG+VQTqsbjNdbrcRojte8VDHAFMsu
uvg8cXVhZo4jpV17vjbNNybmzpW8tvWb7Ar5jjCsZ8qPgdKwJh5xqC2dCTHPRi1r
19ncRaO5LodLWwhkMtUlt7lxzTDPKkqaDaU/utVnxXi8R4udeKr1C+TGbdKj0ZHB
znxeZdcRMlR9/z7PZSBjhrLRsa+/CpoqOaIcKIH9dERkpNc/YtXzJy6LSKh6jBn3
xAozMdOhkC+yccwKpfwIlASNVuI40wG2WrpEGWCEwhiuOneQIBXlA/l5fHk85mM4
Eo55ab0tgregCj5wd4+OsOE+4W+WtjP8dyiQSoyFhBsCOVDuuTRao4xo7mNqt0CX
14c+CHtN8CSgHKFT5tELpnQRGJpB6S1BRjF/jjyAqaUsKjWa0liFixTUV0R+jmqF
jndpn3GR8oAE3Fr8FdovrWunw1GbV5YLCbcyIIr4E1BbvvKRhdR18N3csQAP3Pjm
XuCh4moCg/9ikRcWPcAUIoTTv7QMYlgRzqRmJm5O9mHsnc66/sBlGKOFOspW9vg3
1ICjAqKI2bNcYaeF/I24eCh6cA9M0/Bf94v4YBRQbi6tQavq9G2PuLC/zrYaMrMQ
3NCZ/Nezkq3yboPKBvDRrHQCyWWvEv3tsVN1PlJ1eWtKt22k7/2jUbRr5iPwldd8
menWKwgE7iCTaoWbiutDmXv9Sj/yjRcw7CtpP5XDeTPBE7GCjLi3M/JQtv4L7l7I
bxixrxW4qDNm6TbOC5jL6ZHcAXTPJZnA/7VK5NeSMOCcNz0m6xj0sGLbM6Z2wvDh
3VFzSKkUIdWiDkjZOq05hMtmmc4HfIEB3rd/jXmbZMXO0jaOBZ0uhflIjB/HhIVh
tkX1ECnJmZN9MSSAOOojHg+nK7efiUspOpvWIVlcFTZPM9UIJl8sIRdDjG/lgrD8
JGTjhv4Jl3+VYligXAX5gkHR+wqYAtb5qbxPzwoHH5HfOAKooHQgaym3LdyIXFaZ
UEQd+11x0xspUJMB88btlP0DCJG7YZuGTkLKc2wgqglIfOYNVUyckSsi6s6K4fi1
Fh0RVFRB8T0ByT3Dz+Hw8BWkGgq9stYAkA9u6v+UffcHluPkUzpJQSYkxRrU4VCh
ffYphv00M9Qsz6uqLA+oOpp14qvxBbbu4g8h0+PSNAfKBxH3rWntSnoJQDvxSoV4
aoFApt3CkYXx/VeYdcNyT+R6sv+KNpVjXYT5jQs5MMIK6o3e5tTnVfTJMJG4JWVo
djOVevc8Tk4jKOpW1d3GGUryFrv9i9JfJoR7X8QrVAv9y0sO6YS7wV9NbbOgAEV8
K3qIrM+vSGjY/3U4qlNG0M9phxcvqCm6pbwSCIOUgGbVVwJQ9uLWfBCiGHLphjQe
OhTvOVFNJOWsSp8rqlKMTjl0WaV6zCvLNNADk54W6i+Eyw2GJK7RuA++mPnlqllE
4DePnRlUkFpISF5/57kK7OQjBQh4OhLNQBs/2BGi8QkYMYPIF9cEefJN8GfqjARG
ejpavmUDhnQcnidkKGh7XU98p44KPvrAImWetLTjJmVtIyhYa79zUBsKoi0Cl7UK
UFZh6Vu2S1r+yYTNOPhBASTbU96nDQtE2mOwoy8TyLDd7qceXf4lTHDnkkRzX3KS
HVHdfD9Kni63sm8n2Iyx2e96+OmUtoxNgWvD7X9Pd1bqB4LKmf6IQOum+xeE/zqk
vqo1ekdhjb4dKBBVgqdlSxJeInkbMqYer9Ii/y3NyrVtCWAjeRvhJ9GJih1TMRuf
JdSIqmv6akEb604O6nvzqivsnjbeFrtJhgT1BGNy4EjUlDami+hSgNIkpc1g6SdI
/y7+dB5hGyIjR6QNB66pnrugIeAlHmxUdnr5zcsdOYHBUHe+OmrNXXzdhBjlDnCf
Mo2EFHrvwFKSFt/CtMzbn9prbJe/E6+LP6DR4TIsqrxuRA+vQ3Z09Ck9euNfy5aC
KQmdiquXPbwc3t2SdVUaady0udXeqcCMk05II9tklRgFlhZl2JkzalnWhaLBbo9R
j37MjSC+TQfjnfuONeWulTyBGZX+K91QJHYZuA6aSOy8SL3ELqg5wqHh8QoFeH7Z
wIneVthbPdb5okPz6jo7bZvmz/Sr25ORdNuIq4G+OmPMdQDkrbKzmva8snIccaD9
A0rGMo+9uFTyDTb8aTVCXJmdqsbmLHvZMhoHmz1F9SV5CW0u/gPCYgAYLrvLq0zz
UBZPRzMXiE0ozNV2TP8JcKhynJmm2/V/G9NQl3iA0cU8CBIuQKJdzCkInOVHg061
JEw5/1+A+GUhKp0DhZgF4pC4UQDvB3DVuqptwp2LhcQPkvLVJwGYj1MJB/vsBR+n
JrJNZZApT/iysRwSIO7kKdIeZmdrE6wBn6TVrx1c2s2rpc0wZ+kKVr/A3+2ZyTwY
6aN03reQQ3B7mdPLrzWSO03JRjLZnswvSi8FT3Ch3FKtbNdasKvvBR346FMlRLMK
F+Ocy4Hr7YUi3/WhIRY+yckLrBy5QVCaGHm3cE5TnJBdnC3p4bsoLsIggsuB+PrH
mtMwN72J/erJbHihajpKYeVNdhj1SHqmEFwxgbJ72436qMAXz9xqaYMcOCMIQhza
sacMo9kOaaqvv7/eMX3lFJ7d/R1Wbsg+PtfAkOBetPdB2gx44QR1gOx5w7I7frQa
SPz5TNxD2V6uP3/X+kHWsZvdubqcMOpoLQzuUk+n5mmjzjWCaSGbK1Yh5sDW2LC1
vde+H8BqgWMMbi7i52F2jO9WUJpWXwdziqNec/Z8FeB3Gu4T5XnuHo66/8/+LAEq
5qz/6XVsXMhBVnjGOXcnEt+F5/q2eYmg06TAISTKTRK5mdsddDjWwpv7O/eBogzT
XsOATpnLSCZWiQ1iWDIQWeEIln68cTyZYx8eRyydg/OicdtsOEu6UFZJMERqHSiF
GmN8v014rpTu7mztNppS2BeBzfQHdL2azWhw/5NTaIi6oiuyzoZg4ZJp7B6xYDcw
Sub3bqY9E/I2i0/Tvw2DqxDs25WYhqfut6t9GcrmwSPbWtVFudjmwbVH1FITmHl6
bPitp1F7bTgc0FNLVKO8nC71rUqPKWtmzNg2bP2o6cTuqCbyuteE1xhQgeQteyvN
tYWrdb6WWvz1YJm4vz6l9k5xQQTUTD6mdxmaYwCCdMLMnYqYL9EMXU2btTa5yjbZ
OAvAZHYoSBNWZdwv2SIAx82oCI+2ccCKE2hLDXIIEH6+AqxKygBxlNy32lrDFKF4
UTeBse6MZp8iUXyaF8UGbPMaAD8FiwKWUTkTCWWh3Pg0ehnXXb/fwLNqmOggkkrt
hb6rP5M+cIN970JqKG16xJ9R9iReqAtrKU11EAQZxay8dPIGMNCpKVgo17qhM2gr
f8KYi88JcXhGfsQyRRek+xmtg8x+OHQrWzg2JEmsU7PjYd7i6akD5sDUX7lADF0V
PXADNMZFzHu3qYApM0Sip0VTxDCLoU8S5oKNBd5+LhTV12BmrbBlqSwgBQHujD6D
pSPAS18JiRHDkFzpJkowsyRFIvm2Fnc/x79NJaU2YrbwQxX/6uZwgTwYZsk3r9ml
d74sbjYXL8NrJcVeROleg6NEbO1U0aKevmXVy99tat/H8PmTR8c5zapbE4YachGz
9HtZkwxvQa3ZauFcOGhvA0Sm9Q0HPXAOKTnyo/+mWL1gT1aQ3P0oUnrBnCspWCW2
DrCBCKTm5Y21I+cXMGGAQmb9Gcu/J4gWhqhc7W7f6at+GcHeuv1gA2fEGdTAwa8J
cY3grPvw7PYSErPaF5QSuqrIrsN5qp+9lL92Ej0BamXtNrAVjW/Z5tct1QPFtQeC
jZHJIwbs+S7lMf7KTzpcv1Pt37hZH4FDCo5ShVA3eI0MKWcRyNWfGM3gCJmpmx2O
t/4zRyObEPB2/yKXgEZm2wWFaN3sUPYyHUKXhI/JGwI5Mn+DiUMJYZDPO8UPtz4N
dxaGA3akMHFmNSk3lH/yozZzWen1NF60gFNGSj7VJdir+CJGt58ccID8u0pibVL3
A2o/ps8XskxXSlI5NOjVr6sb8XQy4IFVVSHhBPhs3WZlQUpD5gOnDlPKXlhX5fRf
Rw4EfNK1I4KSTmq/8caWIjhnzMvXNhjWeQ926nN+83lrDwDQ2wN2AJqEeOWfTIfm
5cZASuy40is3AVov4fJMD1jfzftCPdfNGmgGesykbYLmsTAuIZ3kgWp9Jvsr/60n
ckuROdSGtDnTJtQS0XaDwi2PpRd/K9F4Oq2L5Cd/MAffEoH+ovbi7JlkERwPq6z9
8igq0TLnS1pPO2rXe4Z+d49fR3vZ3kiHhYpFfwLrct54fIsXSrJCr+MzAJQXQz8j
66/INFaCCOLZrNw//zn2wSyfLdaP9gPiHnHNlWeaXoqlz45VzK9xZrQtOyA9axpo
9BwWvIIxfB7VFlifDbws/1RCp0Hk5sBX0A5pkUzZVevRtCEUjLi5CKO7sQoutqZR
6hHcgdsIXhpqlHiQtIAAcdxNuMbYPBLS+DKl9/gBRTCfBqX/h0DZ6phowe8AlZR4
LcCUlf9eLiKZyEmNj8pdhdiTUe7HWJRT5fIAvRZRwfIGCV4GIKK8HqIlKGE92tcA
bszoN+2Zd/Qcz1STqQLVoXIQKjw43LHsmF/y8zWxgzEKsFZB4VBUYGF4x/jrerR8
lUDVyKmAfke8xWf2GDT1raJI9arSAX0i5zmL6qLNbimaC84NA9lv1wLyCdCB/RyC
wes+4DHjls8KCdgaPyyZhEyEMMs3VcVkIDfRhRzSeSAZYX2sxSXKutEhaqYMUnlx
NvlYvDle4JHG0yrj2bYu6CQgFn1N5Xn6fH4vD24PIZedp/PXFPsx0QTuziz/S+O+
llsl18zqPgtXuFkhcRnLPSaZ6ICmuY587HaXV/7v+2UWm2zThsUxTo7UeeysszIB
To2NS+n0PbyuRqkZjF3PY8YKC4mE5XSZZrmcJOwWIiJfBGwcmQmJ4VKuWqKFao0Z
EOknDQJ7UwwWSlbDzievvoQ50hnSTr3xk+dO0iy4xzL2qnCEDci6KTppoEUtOayY
9Dl5WUFxypP5XMtC8pabQGWPKg3VZEk68OZ3a/Mh6vTImB97vP8q0xvTENjxngs0
nHFzp/QlxvQ5m6ACwqWZtTO762PfqI6MecBF+ejioBE9lpBIEmk3RrENJsBmo3jN
1qe4ZdTXdDU2nWIqaBE0fuZ5LEBqxOguyI9aZ6Z7+LjD0F4MKX/9vXHDlxzWDfsM
8gUGH3F0pV955//Kn79Wz11jSd95SdHweVqeA+vRQdPtFRi0WE+uSP+n+YcvxYLp
gzkqUU4wCG6uL7fGTko+fRd5QhYzk3bU9AAafmkfsBnCDb5dfTDjVKHFczM3ODnm
X9TU0G131n5w8xEvvmvp9nAZRBRN0xssk8bEB68i4DFhQtTlMiEHKOtAzaU+fowJ
uv3MBwlbKNY7Om2LqYjR9cpz7pJRJbGtRYQ2feRCOiL9EknXevFmSLTtP/z1nhh8
nLFrEM3EH9yipj9P9zpBrB9LPAK9nHdNvf/nFg3sBkQ57JSyR7Lm0uFtRzr5A01h
H10J6N/c6sGaVv7MRfxSTAVCc/FO57m1MSohTWrMPRO+ut0MjUTuh+VimpvPiQHh
jk2gIUvW8WxkyDet3oL8nzaFACNyc8Qo2+EIL2Le2hC+9s5NT/lmAcFPfau4SMRF
7j1obyrEClyGxlay7J5unCLlIbvTsEIi6wcautmz5KBRxQ9zqavVGv31dnQep8V+
G3twKlBBCYccSsnM/eMzFBThRQ6uLdfYUqStzMWiqS2bCirRrI00bfWdHe0fUaDM
LqJAj9pOwSpq9lHd6DG2qhx/PZPnYgg5HgeZOESH8muTcxqUocTsjMw6q/zwnvXY
IIepLt04cx4SQ2Jex3GCoBog6Vm+lMoUmhAhhbq3mLPSOOkE8rB7CAVgh1To3Isg
SsXoB+OIaI2SpQ4X4aYa+D3TyuprECKhX6ZQ/cmb5hMjePP1LXbFTi9+MIO7ucUr
S7QcghupDQ9EJE9sAfnt9SqNMr9f+PzQRYQMCnTo4rlPD7Pe840vNkc2AjV6C6Ug
4LXqvU16H8LAF4nPzD7R1lQ9YitjdO7Uxznu0MnWp8DXLYL/HuX1elSXm56xzUWh
FIt+U8dBjhtjKjl1A9Q6OLTTOEdtbu++g42FC0/jKYiERkf2fsViwNjxgrTXW8c7
J4oO0llLQtj8A3DmC2moo/3LAZq38fQbVAMy2p1MRD8YdST6ARn/tT8T9fsGtqnf
WLRjdDd+g0jSi7sxDUt9N48YBuaWewK1oWgpaL7bVfvqGbI4iTv4aN28s5MjRupo
jnS32GYJS+VyfPFUEJrfLQIsT0EOiualOgQEIqX+11nnnlACoXrMibYvOM8AqCjj
5Nwf83BHPzvpJaAS5CleurDAGMQyCFG4d0sXBPcc8J91AiGNE0Dk8Mm6gSsvV5wk
kto9/zu+mdKR8mrPyyMW+yHQP803J8FvrJHdDkd1VVsn/v8nVAlCmgYWKvu1yoWh
VdXq68VdEIqVDNeV3J9iQ/KCrRjqjE3Voq6Eu2oenyW5RLnK4TIbkiZWuE6HmMy+
MAiHieozZhYa/ej3sfLBQjObe/di+y1ZdrIrtLWzdKyAUeQHZXt3Am4xR1rkwk+r
WR8+SMbWMP4YdUN8u/71JujCz2d+Lpr5f7lcShUxNnnGoxRZxh86WHWrY8NUB3yb
RY5lTkitNT+q756fpcPssBBv0UCkSs6ZwGaQ9MR1bm905oBucvGY0bi2OoDlb6Vi
5frD4/MKm/sVdQu9epMZrb/gUb9FXZyj1bnOYm9i4m9ocV/2RKpCOhGEt4ibzdO+
mZkHbZ9mBaEfXWpzPma23Ohv9wZHYpKikqnAnwxxm2TRYAvCmI22aThxt864rAwD
oro0aS/W11cPybsrLxN6sk0jN9cRZEiQ6RAdYb143PIRAnKB0lwMy+0nOUOp0MKD
op4iIUTARfaSCPIDe8bJWahfq6sVdPInzenywL/Wp2Ka1VhzXGcTPHyNVbPO6fS0
rD6jde1aVTd0S68/afBn/LaFZnYvp9YTs9GG77TjrdfjDNvJlLqbDMAIi2OXR03r
IDcgSZ88e4EYxuHRCNg4fkmcPuwGph2ZixEvLf5m1H8gtIegZRNotnO3DikCgz0n
qFoQTkO8mjf3VNSOoUT+XKcIa40vPaNvBIWYcFjw3uhw59gl1079tBjwKclQ1pYl
ggJlfaP1uLcdjpGkDWwdMuCkf1VOfEiUjIIf10EVkjtCCpb9+Ir7+iHAoNubCx9p
8s4b06ZRlPZl7bw3vwZIPAkUUHFBL30dv+5e2wEVh/kiY/KseiznbU2sDvo2ayY1
uM1rn92dpbIl0JSiyQFjc5w6R3P8R+6JHbqO2D/eT4ZXzvHnvEKTxY/uMGu/LGvD
0DNSLI7qSfwUpGYMQ0J5Af0zb4M8feQ8yNLZ35jtQOYfKRT/IYI9dVcH9l+H+YyB
aOSy1S64IdYsnSwIQvWc+k3qM/D+G08l0aXih95/m+PP05uPlHelXfbyLQWVpT6Z
+C7g1jVfCHJq+i6SdhYEY4Jxsmh32n0LOfLLfqw9hiSOY+sneSX+UEmW+k0KEVH8
LrXDPjmSWATuIedZzOqAnLtqMFs2RPJQLn1jKcxoWRK04m7THYE3XPh6R+nDCw6R
GeGkVJPzZl/p3/K+8UrTnF56KGOtY98yBCz/nit8l3twc4GS4iye222XGlbUGEo9
8JedMgQ4DeeAv2ZVtnt0NhW2Yh8d+tghkoRHBX4hRkfCs0Zae/dcChgW9GBnqGCE
k1E88KALlP9fWH13v/wWV+kRM5lxqLFbyOqqmXzr3yAssEjORt97bUHZfF4LTZPg
w9WZYvGC11vXDM/cmgu8Hi/TwSe8DtIib8nt1qon/uWzAxLfKHf20S/q84dKnY5j
xPi+70zUcUiqdL6qFxbuxH7CszboN3aOqPxnCT+N0TSHD/1HZB8vKKDpKofmnjxF
CwiROTEl8xVJFx3D6YD9pDmqxZqwN+kAvVBs/MEjVLvLPir+fv2H8UCnsAU+W4N0
DGC019GurTewOTKSbTUYd03uJ0lfg4utv30sZ8LjLnyPFjdQWXynqu8DzxjPF4Gn
GVw/BHWYtua0A2aAXaP1iRFO2LjwmcYcSs8FeUgEKwm5e0Glo/35EzyTbKMeJ2bR
nL/R3nNwG0wAeIVZhjex3fgybAakxbu/k/jfNHoQwUyp97YQNcyMkaO2nnXd9wKQ
glpAtfit78qhe/WeH6g6refOg7E59QjdJ6/ixolt/K5gQAgywPQiHQipn2qUeIU5
Hy2hid362ycHBylWGu57IJZGzQvwKOSx8MYOOqjf3J8ZTYFl55aACH89INw7V3A4
557TkxT2lTwXmdllfhyq8sPSazixnL1Zv7Escp7k4v/wwpQUuU9H3gVG7bBTaaYg
hjr1cCeUdWrTTil46n84snrZeSag/WhXomXR+hYsLz50F0TB9Tcg/YfF/6mh5292
sIK0tAh0hgdoKKryIzwfx6DllSUJBHb1eMGmWL0cP9ES3A3yjKcKFT83VOj0m6CX
+YlK7tzahR4OwEAEWq24yTyC2/T3fCJrolUCOZmf3McSoajdyhmVjgWpWmOHI8Rk
XDc88Wd9NGVQR73EBV8txP0goCmY9T7x0rjTZze7niTO+Gz1oDY4dDEOI4UG+cMH
+IaYENeu9JmsSJcjp0Tw/zn5zIyB0MpUKgX1MgZcZLHo1HFdOqr2a8jkOqyw79OB
gq1bk+warLOWyzaWhuywbRQNzeHBWi32EibxuxHHolvefJC5Epa4yJQyn9H/hHPT
p3YnS3QFZk8yg0DxaUYXxMzKN3bYhVmxrKgy86+tWEyYJVlcAolRiiepDuiiMSM5
n+2IhbB+8O57PWUunC3shWP3j4wKmUi8OuEzdZDAo5bsVmlEjffLvT9kh+30uOm1
FBwFPZnLl/DTKno7ZW6qWmjKSDT4HH3rvxsTIFwRaAazjJqlVQIk7gMf409lPcxV
T8sm26rOTPQxmQGVpnXZEzIc3mH1JZ16HexKFll+5P1v3dZOuUQzC8i8idZE6lAr
92rMF7OUfJGdx5OKWi8MpJaAjcz6IElAX/9DEiFZrevEkw9TIDpAQQigZz1ajm2L
CvxcEjMVdFIq39tu9EGRyzifuge6g+pPOAlF6K7LC57ZLBRGoFK9BeoxA4gMDeT9
0BlzlV8CMxWCwLLkEHln8gaeEKe588PckT9DDXERzShHXqgY3jPMq2vC57iZWbLN
2Fbj4IId0BAYBHh/pq6zg/+JKPdezSVWvKi7ybzeGk/qybDbT3lBnBWjpNaNl7QN
FxgAJmO8N2Us38+rVQ6kBOZJST2dRCRCQzEDyJvnY/DOEEflxAcllRD0ErJgzp2N
bdxaTlnYeQwS/T41aqlywD9SZ+RFIn8cI6hpy+49oUFGcj79ajBfgCiCOUx47siw
hRbFy530Nx1jLvqWdHIKAZiCkNjC724JDgI1oqqW6EQldA/qXTDMgGDZz2XoAYsq
2e4y7Nt9K4KbVaGQD7BIyICmRqQ0aR1HQJxEylQqkvnKynr8w7Z4NNkjVT9XsMK0
fj0Tlfeyj3Q4e13Ck1z5R0qGFQNSJJko+OqrCyWiudp3yNghZd/FNbe+ckpD7CJQ
BS/hxjqtal+DbRohwuyB9kKraZZjtTl0PUDumaVuZJDATKp3mLRYT/nneXPzlypK
ZXWztW4H+lmcy/abTakTfswQjEhWHy9agdxSls/OwB9rGoLWWgxJF/GHVwbdbM52
kvaupwJ1ZHRDDdKNhoHN1jsX2as++M84+730Qr/iba4AMYgxuPsPXzrgg85kiH/z
mPAIbZmvowPbd2hz5AbJbtBsZ6m5Zlr2Iy1N4Sf0lsqJnTKTnmITnkvYf3D7bHBD
iJRurKX0E5lo/oMXhGYCSyRyhj3iAkdQM4AGzySwby15uNSfI+hdmN8ee4KfAzbK
gC99u9OurgPASTBYp75EZi+NeGFhhxOwg3eO8iUZBIQYG7tx5DGKGC3oAdZeHlFT
uxDlmOCqjqbYNavuxDHX5NZcc+sRdEFbHVKwsMwV0qRPVwiH1uJW5zuvmHeXG2gJ
Xe0//rOGq8scZovqFHDxKSo0yKFaMH8jvhclpMJIYwZqHx7d4dRBE+9YGWqGlTil
fiGAlICUoA2d413QgpsG551/Xo5qGKhJMtVG3lttjabNDvVOoBYb4tIAOb+FlfFp
wlbvsxfuVbvCtI8+wyMDMi/1ezxNNt9BqYczXjj0rGKCMSoy3FRuGY5uJDvuftGH
+J/+PwjRDZ78zrnZtMQIPN8riQmWAZPzDMfKdRxoWLdZny++tmUILfEqqalR+RXY
0IvL143x88YBNI4Q9GzzjQmst5v2vw/3MLDvRqtGIlqANb+tPDUe8Yg8Ev6PLWr6
h+WaZdG7QhhFMZLKPfZyvTMk4lBO37NzeOMgYM6MgDrx/8v6U17TUL/Sh9hwjAzX
QLGuqR+TIAzePcl9cW0LESylDcetfqLCiAtCmTdKhaGKLmy0mMiXn8QITft0U1bO
BROQ+wxvoggsN+Nxto4bmzYxj34AsAStc/SxizTP0BOfJJtZoWMVZjqLozzm0iut
kFbrdahX85XguozpMdedM0uBMLxcy5UsqbYQyY87SHnlbPr5Y5zgMrw4tgZPYxDh
oGeGz/orbWUUWtQiPFqzGD5iEpCGvs+dZMOk2d7enKeXmNLj2bb3c623wZKIZQbu
CwW7e6H6fsHcn8bd6zdTEOIEnhVjLTcLZox1EeCYQRsPhTVyUmO/ICwVfvU+0Per
FEYcCXnf0kG37J7Hl5eoS/C1AHmSRyiF3QFHEwkAUle0HRURJY1ha6/5185mPiX6
3mOfSNNm3rSFe02povdgieNRqcX7fkotHCXRPuf8db2esq2ESTd55IxEWxd0zXIt
c2K4abKoitwubxdh/hWO2s5UK6/w+rcHowetrBEyopEBnt9Q1F7ijTmWbSEtvRAT
7J5yxkt9FZiu+e2rkIftBsssQ30iBcm3Wgo507OPWrXjQ+grH9N/UUxK4eLXUbF8
S1WRovZkix9UUoDBafQV6A4MdZfaAG4ry5g/2ICq/q5+HpHEEJ1Tbgr8nRhvZhdb
9Uyh98kFCe3L72hmdmfKPdqHv7/4KojhGxc/uQjf3RksDk11DLAmuZoLSF+KNjah
TYAP6PWoAu2at2i2/0+TVl0gjfWuJcQs2KhHKs9Pq/45lBunQKBe+D1hSczP0r8Y
M1gquSE6PWWCZD8+PdNIkWmKngBidu6y+PqriXYqDlhpuR4X2dp8xFWMVp+l6+5U
KAQxdHr1HD8GzVHHqcnfz5zvPAeMznWh90aloSDeAe5Qa3h5HZoBKKrwQYOEahDH
NApV3qZqshcDC+L4c7cnokLbTllSxxOYXSzwQx4p4nk0WaGUdqU+VEFH3M0v9hb0
lxDvpUUar5RG5v126wklu8GWzz2/AaWnnYEaTZTedxm8AYZ1zJasLz0pyjemMMdw
WntYGcK30Bxnku1v+4qxoqwPcbD3RWehHbISyG53ESH7xEQjFXY0Wg6sZsN1ibot
mu6oT4fN3Wb+KACC/Q87YFOzOGEHEYH/5QAUKRoNlVnwaZnu81cbFTm2xWs5HI5N
t8B69D8HBxLcAUawnhg4+HUDL1l7C2k5EIu4ida0Wvt3rqiyM6AgvdH11eV16ZOd
C0ez0pgb3gy8ZMocGrgjO3z8kYjuHWSb73Fj4AR80bQhj68Mh29g0FCb4McFcM7/
Jd/HOwG8370yMsGWPTznmNQojI6iTayIEsijPGdlKy4jBoWdqcfSxEA5oDZWxxH1
RzNdHuLbYMJWJUBkW5JTA1WRjE3A1Mc2G5jVWKRlUETozln2UqA9aJyK4f3WxcHg
1CZzxkbQzwS/J+Y8A0lR6jL7SN3IcBAbGKcTEq5PQEv3LUgwYq4YyE74K+o+GhtP
3dwqCkdvyYQTLsvI5TZ5KsLYnhNGRyGFla2cb5qY7ehFROHVy7d0FKM4Lfw/vt8a
DNt6ll6krYYpitw4P+31nDV6nH//O66Il9I7wWMSWhznPfH/YFh0nmbsm+OE9dHY
E+UwtGgpXE2wLswhYUNyc4znT2pPP0SWMTZeLczd81c3q3jg6YokvVrtQi+gUJ/3
9fFRYn7AeJCCs6WokjIq6HyIX+7mK1q20A7iGFtJtHIgPQmeRwt5CbpigbuSyDGv
VVRqyi8xHoNCBD9hZjNq1WUkngrn42RID6uNW82dNrejAfxNPAtWk/UN1qTasYh0
gqIX7+6xJegEUgNPfp6+AOBetoF91DqlOFAGVpg1mqavTASOR823yMtEqsOplTBt
ap3OcSAeiVkqwASHCrtw8OGsqX3wpOLLnplZAAX5LTR7c9QTNrq0hikzGmDNNB5D
J2PdY11+0lktgfFbIf/q9YWzMr6GkT/6raKU+J+PzNb3FQvUjEK2Ls1B/asZQTWU
8UOGv4pihIa1Vcea742ZC8RcmTQpwerl2WPv+JBF196A7ifJqVGZiIIEvCKHIVv6
u5RKJ4DCHJZW5SGDk99r5TOUBkKqtilNjoQa2r0FCDbnZ0XwrMq5f+4+fAyki6B2
OBAqgidDiCk/VWEw9MJJc3BKlt9/XMBP0dTnMPyT/6q8bN6QvhXuKsC2eu5Keafn
PLeqlXoLwuIKfbLDmiN2Zm8JfqOElvcB5+T6W9B7aZrH6XU9hbJT0KXkQD7zG/cQ
C8etR6GeDlxAo5uXpqfy5uuD2hoq8Ja4IT+DNEMBy24PhUOHF1RTDy1MaiK/FgyL
9OhcUMUt4i1oyZUQ+czRKY+VX62xB9nGHnGGEUUmyVyJTQVbxroKZnDixKdAdrHW
rP1RTOed4LeQP8R9V4/to/MJIFl/Xd3YF/ZGkABcta+X8ogEpB/QsiSTTDkAhOP9
uB/C/qZrGud9bQxA004kUur77vAXSKQb2eES3ijYFpUa2IejrVwKE6mVaTjCLng0
OuGrMqoDQ00sR+NLh4Z6TXiQntC6FRRESlsASW7dvEmawkTPsHNLRugV9SlXx90z
BpUsL8d15LJ3iP7THofQCYZ1anRl9yFyLvyDnIGvz/43cuDRujl1l/fszfEZAXZc
U0Gp5RNpM+w1WRcTJ8QtTpfcHxPCjexayOUbf8Q5IhQrH9fOsdyIz4fbk+5K2Xo7
TyuHxvOlwxahx7EwbaezfXsmZb11tmpiYlT+ptO1Iq5orlCJvhouItkNCrr/S6yx
gZq3N6wAZlQI+SNfB4WbXH0HKC/1okVUTKnLWhDgenMRf/vutZGreiq3j+r5uclE
NHn4/qYAhhS1Dt2NEs2SLPjXjGZXhtNXE1eRAfpLY+h4+GQ/fSU5eIYIWU83C3rP
9bjA6gKC8aHBJ/427laGJUFUj+URgrWWpmf2Rds83KxUUOr3+fsXA00ac3AFOSYw
59uxfqH4MOLCUYXk3DxKLTAWKe/XyGVSDmw+rH8CvbOba5Hw2gvQjNHgttGwC6FD
Ti18akxnzQAURFUqZcQTzLArFSB5tq/GHke6xKc2SQWGF66LDinywwNW+QrwmS94
aGnh5rGbxWAcJMYQ2Irm79cUxMPMZ/9a0+YBc97Yxn8YZHJeQrKCEHw3MmnzHBA6
yYXlDG4+iPDQlincAR8/ZvsJRym/xrB7VcHQNiPh3yNKFfWNENp6rw60BfG8AqjN
53AjyfCUGcl5b2qkhczYoKOYmb+Dj++wlUSyAM74eFAr+mZSzr4PMMFpk/+7BsrK
3geP3kZls8IDUy4FbQQQAF4P6Pe+ELVpHkGPhVDhitX4t93bAhxKmHC39y7czk//
LQfTBHqQIvka4IAUP5s6I+6tH7uFNqN8yZ4gw3P4SCmltSK3DJzqD8/xnNR3NVN/
Ayx4mlfreTDknZuuCQFw88p6A6IR6hdsRYdmXCpR1FUmUizyCF0dORD1qrLX8jPQ
ytZBIrfjE3aed7qgfCMaoZEyJl8aOkJ85tS+faqNC0YhMbhKqtKi1sF52Pe54wa6
rach2t6bOmo2NHAvxQ4II8AN2eAnV+Pmgl51gmToa80gM78UO94AoLhutjpFpUh8
3TctIGiPEzDQhrrqxBD9iyFqANkpiSUQ2I0CvwRDZJ+KLgRhYFIwBh/Do2sl4vI+
6ycP4ULS/koB6XZkQ3pd+yPmc3Gj1dFJGqpKrNRgdke6+C2FJXY+KUIaMEEJZCUp
CIwrgROnCsHJfoA+UU7+U8LKiRitdop7V/ZMorNHIOGLLU0G4GiIQCLIy9V9+LUQ
06lRsFmPdHgWwITULvP31Wr8/bU+5GetWIY4ZLBgpNcbSyhWuKm9xaWr9PUEvGUw
GmE+9FKJ3XIOVZ0IDuzIy6zXH4UI4bvJ1ZinD+oq0UCbnnxvcMfl/XxyZLIduet5
hFOemQS7/1U4Cwda6SbTVJzVjDlsnVziH6bzre8CcEXL6lefDHwpajzr/cPqFadH
yuHV+EYTHcyzSTevIlaALT7AxRAjBOBsmlWleNUoZwKpdJOd0jveZsr6L6Y9KTJg
3OsUgLectNFn7RKAvju/B+hsGRQoW5hpv7oAN7fZ8ZqdP3/d4RMQI2Yd2ocela/s
FpT0T/l4TnYGm+/KT9Na+BpEqmDfWj600Hligo4K1HpuZPj4qr+ClQWdMglLj5aS
hCJ4DwjvhFPtRdDv1v3XZdCT9fGdgkcZ1+Ms3F8MQ/2KKzf8+z7TrhUWJxizrhuB
GDgrbOBxpHrl5I1szP465D8OCu5Rl8fCi2+GerqSgkX1UWtYF3O+z7loOCrmipbk
zsySXgyW6/U49+3Rdzyl5fyK1wfy4ysLJAb1FMWWVoVckNgnvxHwjxJJsI0qLZL9
v5hY8GDznGx6apMJm5WkVvweRJDyl3VWoc1R+t8RgPNLGJUS8vQOBUa8FSbkTdrn
Tyv5fOxkClppNJSQoPZpRTMNxZ5odtVQRLGJtKfabVkRNzKo7qvfI7fFoEg6RomX
deGZgiaWr9MXyXb8dkmZlMZcdm2O92YAiMOHVAG5j8X/OE3F8ONZwmqMrTkIWCvM
TP5E0B8d7yeKRd8rzp9P6w41cuKIUJiC0v9beZ3nvkdjlidXDjzfktCNf+aPONgD
SAacIWU0GCYgNxEXGIOimyMi6wpjfg5UbyDBhT94DseTE7XZeQWbJWGO1iFXBK8V
WFMWLQQglf7OXGSkKVxDY4PpBb/5lk682YN1eLOagOb8agr5eS1+iuvYt1DKleQa
K09wL0tmC2HjxU081Ohsw5sRTjaEc+yVY3PKefZ1pDAX+OraMSeTh6OBTVomRWav
WgODhrWSUtx5Uf1Rx+6fy50LlSDRXujpqJxNhi1UGWx451kAfLok+FveLyPPHi0D
T7Ba/XaCs0BWIU46D33hoTOlHu0JCal+pwxeUkOYZjyNOQnhTuks+gpTiW4eTdgU
GlmUwM2DUBMvlXVw4arO1W/1uOG8gyUfG+eMsMB0V6zzwBt7rJfE30llnXCjOIDR
5a+oc8d3ATna+25Zu7zP5x4fcjWNKl1jAKHwsUFBxm1z05IydPv8ri9FsI/9F8+o
h9nDHL1zvwQaEUU3WmHZp4dCPaOY93b35AAN+dV9Pa0HWkVrxeAWPmtK55mBBwRJ
5oCX1+Xgcy/wXCXA3f5eDGLEyFB8Drh1inHlmWSUMNz08DaZigPWG/Woddjbo5Td
aA9KG5N+CI7x4zcCDL7Cs0Rygr14UuyYM76b/D8FCNCGc3RIwPt61Jz/52K+Z/Tz
P/+hHFOaxGy6D1pC7vd4WfXxBGswG1s6UEqjndShq0SyVn+ujm/Lk/e8eMeNxYvG
D0d4QgpfUTmsxai+RWAktl9upG63wI+IhT3WKWiLBQva94NWqzniInIjlOPbswPW
rKEt0ZupcRlrsbdr3LR+FinWWWjfYNAEHbvTDUCBytSX/yys3w20kde+feu/8aSh
ITtt0e8YvNRv34NSZaHe4XG2A8APXjwAATWFt7CjAxh4wl0P2mdkgrgb0W7AlA94
TQbsiJQ9RT7wGUQkARH0HzEtxCtzgztfaV5gFO53Xje719Pjkzy4HkSdz24Mb92a
RRGV7fgmgXCURWQ3/KfRsIrQU5eRKAMMEzugrtM1rgx/5oSlKyA3Hte+91PCcrDW
kXrQsYVtvgsW1ZruGeqmRLZA7wWapMX4vQg/bTVptVWDP0/nTDYoh217CHrhWJvS
SLX9+fM/m9Ns0I2MkZbieMxVgwXtmqYd5H3ilnBos5uvoPVM0ZeOs6/PNhd9PLyd
p/ODkOq2tobA86VLODPzuwKg1JnLm6/o2YY/xk63DrVv6z7LcPxNFcC2iv2ovPUN
/ZfuHcF6+FvGjObSNxdOhR7qxFaIDu/dAzSmQOj8WbH51KxfntEKB/J2stkYnqXl
9VwohJ0dAEYXjVv1/8+tCQ+9jnhZQUyg/2POLaKN6jdIgTvZVUEmfqqtJWbvvHTn
mPz5yi5zx/nMAR4KY5ZvWya8KM53edVvozfeLVj6S/wdLhnIecyRe5yhMX3rYgLG
RJUUztGrCmGxwwEEbiclKsNQ/Wq5tHLRwvbYqYYVTxwCJEgG1HCvZdXwMs1cafRH
wl+N4R9xio1KBoP1ktc/WXB+JibSCFGFNQSkoo/ZjkDP5fnz1GWSP5EeOjO6tEJz
g1qLe0ofkJdPqQHhIQwvtrEuhR5FMktZ9IrPNdmatfrUKSo9kcpyZBAnt82GVQKF
vSDs8bzlWAkWtnnYyc9i5F251UDt7W6Bx6Inp8UbgYnXWsaQIi9KOQj7zuAM+4Wo
CLY93MYGYdHnyH+diNyODon7uUUEbzdnvCuN3doOahwUP92YosDiWqCehMUnUkp1
dlzRgzYHSab+79UHQf8HA/GIXiAdwHgplF5Kv5Qo49/0cx4+DMSPRoPjxRaQtQft
VrBOPjqxJ2CkNke7zVr5QyNfRehoPjE2Ey+jSzFqIJWNLViVdQR5WTzBgw67+lcC
8lfR/p0wS9ypbBtOkB5OO1UXzB6iTllHzpAtbHuRD1Uzbbx8nOYUBHH9jkbsImp+
6qS/TX8PMg6r68Wl1zJ36RSA8PgKEcV78mTOrqfUJ6mXp4fS3ED/lXqV0/xIcEvD
D7/ofQB2LbGEZ0oGE2/p2mmzMas6IMMPGxX3ohp58Wf/ltf0n3MhFO+/A3m8RmC3
CkgaNocql4U9XDeFxXBc+e2QA0IgO6L+wtlU0qw5SHRbkw0E+AMvnffWHaMndlmv
PFtzfEInAIOFXOuHfX7jBLuRyp+Icnbyh70YltZyuKaxTtmRX8NvO7T/Jwre3vBx
m83gi2lp9bLQGSjDXb+txYg6BXEsxYsVwE1soC4llt5MCygMX2qWsLX7Ny8GM+8p
MaOHeL66YY9hv1X/GFMph24EfWOMDZLFo19dMgrx12NjnFzHar5E6q3R/r1FGKEg
t8tiOBSu13U8Ff8cpF0SQgw5zBaC9lpO01SO2ptgfQJAlWWrwkNgwXnGwQPIA9L2
5VJHuekPG8mPv/ZP6ltW9pA93KT6UzEPe9YJa1qtEr5+wzXAXnmYfn2iDCr5Kw1C
rxzmvxGy2JlucFoFXC293x//OTfXOp7h2xbdWouDc42zCoCySVyDZovSxj5l+7Q+
n6h7+OdhzY1zGICmJcTWkDOJlRS0MO+ongLOqE3xwCakdoEBG9tZI7IdZ+9xjwg8
QIeEyydmhnB1Pmmd6nuZFuAJxBLJCdg4ildiCXASf5iljH2wIu9/v7QTOV6j7gku
vhBvSlfnIwNYVSCO2TM6EhTs01130g+UeNNwtUiNEk+UwIMXmAiUXq45EXHHw5oE
IkDJO3QSEVvwfG+lqC4xoDADVBGwfHwm+fNoqU2WaIcfMD4NJ/9mKipaErJEkiw7
frdHopN/2n5cYABoPZ7PtFGVM7q9rJB59qwopGB/zywu71U/KfN5JK9nnLI4DgIk
kN3Vs7vRLjmAwRXPQUguAPJESUfzyLjwh6PgFuXZuEwwKjSJuurPs68+GtPlUi8Z
0+sCrCNH9S7z4Pnmj4t0hAm3HLvcqh5xsrVMVfxtP+nlKJqZUWyuMWEWo4jgRNZz
GdPWaMW7s0NKPgugNHHvqlkBdbpVhmOhsZw6pnk3A64UhxpFM9AUxUvq0tnHyxam
TZcA4VDd0MJfnnKBApTjl3b0q7l0DzL9Ev+q44Ip3cx1M1MpGEXkWZqVVpkrDKbv
3Q/fxPLQ1zlrdQfnI1FD+EYJg7bCD3TBFDvtjVu3gvArMj946vbuKo0u0gt3w3z4
xcRUyS1Qnfw0qHcMwRoGM7I8FW3EYiZiRPqgTpRIwUkN2FC5BjWS4gLL3sZCWuUM
FjzIAWBI3oyqxZI04AnAnMxNn6FANyG+iOqUpvyqjGuYoN/w3kDxL8JxWT7uwb8W
PNAf9Ab3Q9hESQyQOd2ppTlsKLdfYnlWokJDPT8UhpLvk9IKLoI3dKezjmNbuDVh
VPgYPcp23RA2RRB2fmLKt5luYDrwRsNiAm48jWlTRruWl4X1HgIuIDsDMBVT1Q9W
j1Ds13Npnl/NaZ9aU1yQgSLb0UC3IDuPOi2EV8iNLo5XSKTccsU1dlo8/VU7TjO/
zUbhCu8de0hAoT96qs+62tNBaqaAubtRiRpX0BTsU4n4ID03k8ZuYwdIFmBbN2p3
MxBSOwGCOU5Tm0ZWHgd2akscrdn4qpKJozDhcijBa1LJIIr+Q4OaqtX9EKlAhxqa
y6cszV5FbHZM0IAG33Un7r2g0Vz4VrnStvwltqgaypvoVjvBSc9VA7l3ytBwJpHB
sKI3dtikAEX/1WU8xfwinWlzfre3fl3oYzqAGXEATTJUM+vGuKPyEtWjhoNqACQL
wWuuHlWgs3mZHTMW35jVV8eDsi57YERd0DXgeiGkUvercovJ5qjmEa76bORqHnfG
Yma+XCFMRV2yV8o/JhQrz2l9npMpLnZb6vhbTaTtNJWLkOFelkmffVCrjcelBF/U
lwTNhwOnfd2Twfpnnz1xT8VO/FXKA0waFxXiF2FWeSk882fKHkVPqlE3Dax/anxD
ZvwMssC0W56ensTOXaAoXQUrEsml2oksK3jrdEJSskRjnoAn4X97s9myG/t8UXPa
9Aa6vY+YKReFSjptnxDDCRaO8IClH2ChCHlUJpm+9CTRXixgue+tpMZ/G97hWEdW
yGM6+i9EN/UeHlTJHt4OyORr80iISp0bhllJWgm9ASKQXBxaCzWxavixO6a0Qm9b
ebcfar/87hpfWUCds3mxV+Vakm8ZYqgSZA9E7SSIWre0+RDEIzNCICmH8h4jPclt
v8UXz08+x6HYmUk8H76QX/XPLjCm8Rw5Nwjzn+yCdRxe5teDUKHcJFcKpE5EK8Cs
gUMeJlbA1AYM8mPbkDbWPxAvpJDB+dX5pHHub9F9ns0BjJJFXbhlqmflLqwk6Zek
QZlSYJ2P1qH2twQSI4QuYzOSBcikPLKXTzO4QF1CHuJvHJ1cuMAlnL1CNt5NJzzP
7nRqXywgzVFaD04dOhCfUQIXDJlwY2CL7as3FrdSwM5zeL7Z3mz8sbsgQIPCXug3
exdXnIlJIvvmbgQUZPxznLPDGqmm38YQ+5SdSclXWUBzCNMFsW0L43k4LjN6AXdn
e8IwTW6bOJhIb1gp8OhwR3Wl8AtNLWQM05p78Zn1YEIXe6Z0n3r2vG46HLjI4om+
cKFA4MT43t3WaxotpHPPDb3ct80rPbgvn5UahZDf9YxUiRxUefaHY6A8zn39j/ed
3ShHWGIWi4zx/3x7jYJUnw7uzp2wDJLeuUrN+QsWm2D89dB//gm0lGNGXv5Fsurf
y74yRtyX8ZCYGitDlB4GB7C2RPbUtrCa9CqzjmgqBuZxhLyxR3XNYZ3hjsv9QOad
V+akWbweNXdzLLdxcdpLNH8NiBeBx5nQosZVvEzBXCISSt4fOkAibnimdcXfvOOT
XbTcrQJ3fFpvFgwKqLoXKRIn+IzM7UE1tbRV++zs6P+rhL+6NFrwFQ/bL/iQ/riM
FQpWSlHBHG4JFyIIE++DdY26QHLU/U7WUd4Ts5fzp8Rqntig97zL25egXDstNA09
sbtfdAQdbp48KTmI5+AxEKuUvMwP8jgl8ZLtWAAwNXkWyFQD4U+V+a1JG5nBss0o
m+kd5ufq1A3hx/1Rt7Uoj/2KkAQ2RlZIuTWUF5sC2xPPFYAdGaXVUgB7A0ukj4gJ
dZLhKqp78TaCBCb198W37OSEWZL8Cf4zzLqXdv9f11AUlSdhnXe8Bcuo4NQwRc8L
fGB5tYFStFUEPIOeJyVxEV5PpIFaf+yptpd/9EonB8MMejOnw27+/nJtfMU7WK+N
9wgGCfDySWLK0NeegjUwIwb6q8FcQSqBpxXBJ0qZFLZbYvyT+OpQtzYGejilg9DL
i674qfAfGIRpygjss+gRswXONSkwlm5bAJ07m/edTwN9ozi1nxC0Wc7ubWtcko6A
2RpTjGUnd+DWl98um7WskSH195oZ45gaxX6Q9YN8JH4xl0FpTwAuFTH6k+rteU3V
eUwtUhFRoCKNZ3qCqoIEEGCya7/3jdeThSktt6ows82BA8uSod99IXSx9iqJGaig
LlBfAYr65esnZCy7tc/zwqZg68M1HICcCHUrRD4BGDkyNYibuDvFeA5q7QvRFDOJ
M/FdpUmunva/0hqPk1wbmpxDgyp+r9NDLPbpxt/0a8vaxiS9iRwXcyswUf9CSsa0
hhZlHpMeO6vKi8p8wPgLrapg9qj2WQ3rxr4orb7Hog46W9sOVyuME6VgQhBtaeaH
qVn20oWXJ2lSSZ8OelmxvVQzkrwr3hCZAWHGTSX5LZEBUmRNIhIQYuTsHUvf68Zi
AFR+MoOtEzcivKSoWc2UGCApHGJrub/OV5PDt9g9mkZCBEmyigSdXkLtvVjhjLWd
KmX9G3jOHEwAC0aDNY4M+LYb/uJN4sXxsKbeuHGXOfz915nWworT6B4/dBIxY4Vs
pYnz3kekh/roX57DnqieetxDnkWjyneNH27zdq7419w6udrdYc8TeuoDE4+GNmP9
vUwTUqz249s/e5+eTUDQzpjS/dMFzCse5gHGIE06AWlRvT7grVqwBMyyVx3yNkqN
R0bhWqXS8cku02ORVn1JK6aOqJ/hXFtejZwXXyv9hwpBJjWw35EjWfW40FkxXCfe
TB7ckQuUlNEEJayXwq2tZ1ntEYA2FWpgTwakqKag2j2R6k/ifD6MfuA6XFDN7Zes
q9V1J+TISnoSFWanQbdbaFf1jvBq65N83QLD9ld61rAlEkdcjcKGNm7TeCXpd10v
emVr5/kf4rnGPqePmBckal+IhbFpe7zqdMJXX/GXkj5EPTivGfW5AyMPxKbbnb4y
w5mKYzwCRt+FzDS3x560QZO1JenboVqqySGMZEntQdFtuzDUdMwhUB6CdFCCCAaE
T/rk1ec8HgJkOr8DkmrzDYIw18On3ANebzwhZP8QSTtiGHkDEwZMRtMM96PydYNR
QqKncwdjpvj/3vK7nbf+4UqKR9KKru7Y+A6T9Phw11PdRfOwR871OMbtssZiU93y
3cGeJ8rP48/ZCabiCd54eAGqxl+E2rOMCdzEFm5jLmhjWK0fgIWVjXntOanH58hr
d7zRN1CRA5zlXeFM51LLLcs03yno5lNe3L7D3owzthUmpXUA33dUrbY8ezGMzQVH
7VQ8zAFcTopHtePAmDEi1Ho2MVwKHtni+jVle1z98m38C0pwPu7XIXg1NtfYSbe/
Eg3BKzJi7xRJ29R6lqP2e3QnqyvRaXpSoXGUCU5T4l3BRKLPg2Sfm5QkYj0Ol0bO
0+tOb5/DIBFnYoeDYK+IGJnOz5P1pOCGM4F+p1TS6dPZIuSpzB6H2NG7GlLAIs9V
3L1B0H7edLmQTSkvKC0ebD7w+k+ECYL2wZG18y8Ohy6D7TxMhuZUq0hAEf46lPOD
y4rHFe9WVizhPDvbPzs5RAXzR3zYPJGyLZiAwie+9XbkF/zHfyzTB83MRj8S9CFq
HAWK3kMnlJxyEfwINXSMMooQd9/M7J7MfVQW0oI49z09LlfjT9OBfpyOhaDXjTtf
xOyLpCwDbt0FJpb2stZcs/t8SOLIHaW37QdsBtmOtjl00WG9r0GRzqhKEPKjKUsg
jq88xPJcq9bI0qtOqOOSugPFbYQOHjdBPV036vYOXg9Ln3gys8jS45o6hAi5qZQx
GkYMeBbX4Ko6uP0oiTfC/t/l5qvta4l02vESkUMi/7j6CSDEf8zBlzhZETVD/5T7
Q+PprsalzaYReJ2u8qZKFi4G+M2NoFhvMK3c8QvmcZzbU9nKciDTGed3hkDHG76v
qE76huMZuDrOUVmRy64kVzN77pdrCf9tfGqo2G2YMPP36l17RN2uPSC5CQymi6EW
hBDKkBIGOl+cGa4IH6okfg3fWinDmLPGBippanlr4NL592EFt1cvIjTUv95EjluV
5YjzU2lmLAvZNhfNQsaDYzpYcy9eAWLDqkR7kywh07JSBI4/N3cwIizYuUVdcPqy
V8Agocpm4wdpEnuftXlbIvHQv343anWaZHN/Kub5fix2YYDg1KlHHkqkFg/QJEXv
OOM8sMR8cV6VnBRNEYhXKCWkOTRzODCBNueJRm8f/MY32K/RxvHKD5LWimGkbYhp
bbjPxXJ0JZuilzC+FBn9JrAZnfhTM+pmuWxhsWIwxJ9Eba0a42bbA4ex+hVo0PSF
OwwPGTLNalbcDLGX823sz3KMUWL/uMVvhmZztMTa+YHW0xqpPuMkiaLv4Yi4N1v0
c/i/F7mq1XdRxV4ngc9QG2nP4uG1S6CN1pgFJBtuXNFKDyGIuDJq3pd2MKaCMwkm
2zUaQQqA3cnJ2YpF2OEmxVszPIeRK+xfwNZ2Mf8AA+JoiQI1LejMyYgzWPaYvXkP
nLTDoWzA7aCtPvWeTj68WLidPePfvqjr7scRvViDJ3wHT1fv/LtHJD4Ot2oqPkav
wRftgQeGr33Zgex9kcQ8L0+/OzmTSLk7C0L11V6fEwWtiR6ZHedxwhjJhZQuz0/7
FGFk/n/ZtP81Fu/GQ7PxWY/N7/WeLWWANtm7Maorow2gIYhH6BYSz2PSinSpWExQ
C1+CWmTLQOtgyK3zybtvY3JhkYQ8givLeo0pmB7B539u/0C84ANPmfhKwwC7Jmwo
qdfrumbnIP61TL29rzG5URMlg9hn84Dc6bal5GNV9PL3W9+FNOysEK4q8ObrmQl5
9F+B2ldp4nifA5QWpZwQQFWNgkEsq6Bc38Xfa7qS1IJ6DfBkTyif+cV6+39imjgW
O11FilB79gYDsW21nzgGLJ5aZeIIVA+baryKTeEds+7E9Ny+74CEeF4/MH5NHUof
cxsINDvrKTAy/VFPfa0VRkZvqhQW9GnDmeIyhaD98qzv8hL3erqc8F3HgTxe/l91
8+V635IWhNcluifC3XkfqkkwPIiOCyKrWuLGRP7AWhMRvk4IlGba7IvPS7OcI1++
7qclzvtGm2qfV7yoNJWdSMTBiDi5JouDwgZvM4hBrg0zC72AgQ4zA9cOrxxgaHkG
JZchpooVEVg2ElQBLz9y3N3IPmmkGEdLflwNKOXbf0eZlzfviQd4FAFxrmIjd9Zv
RZ5SV37xVeAUfarw00t411eiymVSP1tb0nGz4BvG8QGrOsDFz8FXYw3LdOfwjveW
1/+UEkUFUnVzuFjDr93iWr7ECIEhy+CjDARdaiA4lg5NtPo7KYsAuNWSQ41KOnGQ
KHphx5zkSqkQn9OtuJgQGc6fXnfye+U3/Iurdd2HdBA17svmrzmI2iGFZjRL3q1Z
5vBd5gLUaiM2z/eA+2nUbYtx9zHT2hx8Yer0tKLoRTuabWyecD3mAJ69sYFrAHy/
NNpgd0vlIo6MGXnbD32pAzm0zp7HR6uOAVE94YcRbxVlkXBmS9D0JkgfA8dsa0+e
7TmCTnkaC2M6zv8RN9EKl3VJaobDUj0d+UNgLnMIgUNtOrJezO3LmKydgG2W0PHL
4Xx8MfyzNsnO/JmOiGL2hWJxw3qNnkeq/z0ASMeyriP2PaRJn6x/7HDi4uyFsaZe
1kbrpJ/T7AeBZB5PkGhyalaIN9q/MHFV1xzatkoWaz/F1LvVdOMv7EtJb/0yuNXX
d9XFYjboYLytxCpwxrVfCQSwr3aXSIG7UkbZPdvqk26yWRxYTwxnAGq8muEgRt/k
Q5gBu+H8fiAsQ9bD3Viu6FVwzaSqJrvJ9WYZcotkRjPv4pVyase3D1JGUfUe1kq/
0Za7HxIi8UNxqusbnlzzUPV8uaDyvlHJaQa12IOsKxgBg7o9MfBHAUCA+ZWM0z6C
G1kngz+xPGMoz4Bg66bopTJsISpfYh6+ysmFJ3+md1IYLsuDiraRl5nI2QIr29nt
aeG0FaHt87qdXiEcoY+XKVVmcXNkBhUezXhpsKtm5fgBKBwRy2US7xvl82vCOZ38
rLi2Cxh7wX1bQMxZh5oSh4OLOmb267DZtFGrB4UnPxpWvX0rs74AREenv2BOXfWO
4yRPcAHN1gEX16FpMTzZQbq6iZ0kM0WxfYtm5hEGpavi/93PwFIowdoSBvVDWjGp
9IROhkuEfAKVBJR5f5pWO46WdczwoqGly4IqEDXK5oHbwa79v5ocVAGu/OugBlKZ
0B2AunslemMv/SoP2QJRItdoY7YGO9YGiqubS8iOJOtXjFm7egGilU0GeyaMQHNQ
uyuq5q4zBLUTmhoc16a3WtYqEFp8DXZSgFI7qLURkvIU5MwTn4WK/bjZgvMPSVdL
inG0MzX/unFldweTnn0u1rNEq334fquwOjNkzR8XtC9rnrH9Hu0iVYdCFjS4Umvu
3QaoohEJF4Yjal8LH/BGh63Rq8slrjo0AWMzkR8u0PQahLG8c6gwksq/D5SwNlZq
j6Fn/RoPse3zPIokX55RdhRUYnVQisDvZuyQ/MoSL9J6vHCaiNi768l6t9qtJkqS
fKxXRZk1+xJEj88FI8Rye6t4xQ1UQNnkBc13phXYSCtpTn4T+VlRpRk3D/EAJUHP
cbE5kwQr2qKwTcuL8Y4ZT+o3KsqXuGcp8K4/ogyG+HfBC4c8CQNdsTbPr528lGSW
UnArVWD93umnau8NbzzvDv9gkDxcwQIj5XWJXsZ2NuEOc+Mf56EmnkbCycFrmHfU
kRhkhlzxojiNpNbghjSBGlCnUdBxdE335DIbnx6U0kpST/e0DOT/VAkFIHVpMOO4
S4p1BbXtyX1Y8Ktl0YiP2BWVfQrifGdMWw4lh0iVZ3IE5gU48qOIE1dTBpDWBBiE
lm6riyAf+N8tx3UkaIYgBHyNHa98QRLI506MjFwfnG/pU004L1/ODio2TY7tVbqE
Siev0vDisfPIRGgMF+AAAELU6xwqKGCevUDFJSQpVgXykwxWMuTgWttP9KoEJXZQ
cHCrytsLypLZP2kipQXBcOccN8K4xvaIwH3iG8hWkkQruODtWyqT4X/1BL7vtmSS
Q5EezOW9oSa9qoLrwpnPrk1BNyxgocS2C4iFhfKQg6ZdEBADM+zkgp74M2nkhpf2
ddMHuOUJp6xudHWkepcqV3NTRDSNzseGy6/84uVd8PR1obPF6mZuQ/XYP+mRWYK7
fSr6uhw2XrfmG9CdruiBK0SgsGpJbb9PcCHm/QEshJlKbDAquB+KDSM2Iu6lEghR
bUN9MxfQpBEfRhatJ2r7SDkzI4vVMSWt9Vt0SRPNzrcK53kkM2A+czv8x2+Rf3aq
xJPdEKmVyHHXoOqrNnxULs8kHoYoI9pbnWP//49XP9lH/3Vig/kzVHCSkfkzi1yY
/FCvR5txYaBEc7+D0v8BWmQMPHLIAy/9+s/8nQTlw2MNAxvefOpbLTzTy/SS8AOx
PiC5cUcvt5+P1Z77rDpsN3JbbFLpa/YVJ3orIzZNOgT/+2mOYmCNInfz+q7UkdZK
Es0hH8+ssMT5doDEZXjRggnvy0MG4LHF+FaWJWxl3/ZuANm/D155kAxxsmSevbhC
BtHq0cyrJnkaeliQtXsu/vLKTkWq4gW++5Lj2EUEgEoInJPRopgOKYe3pe+ZRItv
Jeuzbn5Lt+tKDnEmrTQkmzbgBxfBsMG0XvsW5eVkJlq8XiI3WU07vqfv8XoR7/jG
Yi2donsNxMBB1XTqOxKH0Bqad3aaoQW2sidwuXWMLi4fUeXVlvXaBqOuwxkT66Qq
4l69D2nnIhYCne8oOvOCAgXN/fWoxpjSnCnvi1nb+w4n/3In6sKE9G+myNown+mW
rAFK8lxvYDdKpcYWS1vojMqVsir/HsboFpguK+aCP/pTukrHNEnAvd+7WR/VJ5TR
4U+y7qhfsi/LVYDN0MlVnNA/PQgZHjokzjNPkpitExOrxf7yex4L0clMXJ61QvzC
/m9stELUvFLrTbXhuU2RAzes1Nq2tTdJxPaSixBCrWQ1oYFzyhZjJb1E6/cpAFgI
47W8Wax2PGiSZSBRU3noISckmNHJTrVgrniYj6rNea6CBW+DYCbSHggXWfwR9BQN
Nr/3VeY7dSJYkBF2xpbXEuYpHmkHA0BI/LkpMsMDDq2f9IRpxc4PB3p5eXcw2Q3R
3UGujitPe71J906Qi9I68NaEZ+8INCmWGE2GIyf68zS5btkxBJ37SJSr/QsQpB1U
2H6AwCVkO8tb4NfSFpMbHSg2HMNHxnZku5Rk1ff9Ynb1J3AyCNYCxgWsFlqvGcn/
iW/bEd8r0quA8PvOeE70es6KgN7gvx94FoezhLf153SWa+mNqJsv/IWPHH6akpdT
6by/ilZZ4PZ1QHAOzetV6JxR+0+STgI/NMCO7hgIyPMwMisWCw5K/33tNn4nJWwT
WFpGl5b3wAZxGBrZut7RbW/0k22roPz5DwQHZ7qB3x6lAg5d7KO/yG+tfKcC5cmF
xW8oq68SGmcvb28KtN72o6YH1iYaKEUR5qWpr6BCIBgVxQWATKyYOeKupvXweB/+
Ck5TfeFCW2dyw4nzcSrUyuq6xG6njXKznCWIyNsq4Rt6cuzpoAms1IsTqKMob61w
bbwEsEElQKDnNSDPAwtIKrBRvgfKaabDulZmahBYlywYh5+S6vOWXTAeAFWrl7lF
QrCXLiaYBU7c6HglF32OFKtuyUf8LeORVXZhKHkVKDA31+hAZwZREn72qazOHWfK
zwDwT9fCGrVNKHmdSvCDCG2rf3Bq9uOhhJW4YPKPcWoYIazPsJdpxV9UfI/P4lHM
lfTLmuPL2h8XvRKXUZFQShWFGkwSQyANEd+BXMDa2ker4JBiKWtMkgydm9TG0Mgy
UIDSVDGh9K0NtXfoo3/uZk+5mi+4xfpHmqlnp6fnFilR5PjWRnOWIl0uUVl/JVrg
eby+e31+u+TrJxbPNBtuFyXYsxuQADMzuD2xDnR2PE0ENZuDpV/1MpjxjMc+Ds3J
8oAymwNy4sqJBllyANY5J1Ia9nHNR/WodLmv2ZDFI2scP1iPJa3gH+jp3gPL4ZQx
f3Rri3PH4EYI2xKEloINwdVkK7AFUoTEx1TvAccVCRxH3vhBtnw2+Mx0oICzXIYQ
qIG9ytWSt4g5N5WfMbLXn3/CuF4oDe99d80qaL6noB0sSx+U1yNaUC9RANYtuVS5
JkEk9TdKtYo1urGY9s34mTUtfxE948MuIZ1rK6HHdBM+NOD0bGu2QcLZOdfA2l2m
J7ADDcsNwG9DS+PTlsW0xx12LTzg5kOwCVJZRdzwYYfRZr6nhSaB3E11Fy+jUBh9
PH4SG3ibN33XgoBjZeLqthc82jvZZ1G3HarzHF2hfC6i5tC5hMNkpeSouQOADxbS
I/5nNkJg3qiNLWeEHE72Ith/9YhyzxDw3W48NWEIP61dVkj6KHhjcQqNSvjt5Vwj
SSEh1jLyaiZl5kVc6aVJTL8zkHpCxfvd1J5kYzAgwC80m0RQMuKFW6cZZWPrzeWB
ZKVTVQMGDacqgoRVc//RsH7JeeMDiY4auQnaLcdroXjSz8XcL/AY2s5zd++3GkkT
6HE6/V+GIWUg5K5ujd8NHAaCqWzQKPp+jWMV3ZVAkkScIA6Cf+JABpi5M8FYoHeF
OPWPPP7Iha0UL5ZzJ/zSy8Ua8aHSYF/INiD2rYerqDOjVrLbDHobsuet+l733eZn
LahRyF9Av0mwkczgWH0a6OuM+uDCaQb00BZXTRNVC2F20Gzx3SkAmqPtnuH6ccUA
njRDNYy5M2vmo5DfMh5CDG/8KC/n6jpv3U0CRB4qCyzZAU29QhwLisWAQP1fDSr5
XM61JYVOY2C+Yfpj8PzNNyfocXGPx3oYW0UNzGY5hI747olikddoM0I1UkUwfsQ0
WOlTMucHRPb89vGWjoGtA6RELtHUArxkZzTnqwGH87Ki8ufOR/K5+/VD9PqDHeIr
jwDNWn2/Ep1qCgXdem2mOQeIAT0WiEvMqGVoGiB79c/qr80/hVT8V2JbRHJTi8fn
K4mRXPOO1Sp4YDsvP+ofoYkbSzJhJgdMuKUXhD1BYZI5J9WySRDj5W/033lOAsOG
x3vJfw2aVjh0pSbWtk7q3RkxdAd6NKb/+gkckl4IPdpzavCkqjOBZZiLXVMBmh4j
cO/i0vt1BXQIGF3ajW57o9+8TZh1mBDaoea1N8MvKcYC1vPf7Y0GWgRw3aJBdSn0
OOkI5wyC0QmkZ4PgzYZ5X/WBkvt+tAWHjfCHIqlv/WQutMVkGiZzKmVVPPzYcO42
lCjXl3d4k1/ZAIfrg/pKOs7kIxcSmrwCthCj+RHlPMzu3FXLPiV/WDyg6HV4liN7
l2lmTb3tZMvm/1yyNoW/iNPOoSD7h/xo/+8AiwXZviXJ5ahK37XUKshNW1MENPTv
36LQgtmi13Fvc9pMRwA3gYm9mcdsv6RuA/XVDMZFarX5cECUEEd8/BDY6OqrkOUx
4yUAoYK7j3jlQKLeilRYsfetClnTiqZ+vN8N2BQ6qeakE41JStcrAr8fRMcu4Cco
bvX/AxR1pKAvmQGNUHCFEi74d2fIfEjzSC3+Mcs22aIavq9l+5BNbptR//Nknyx4
uiB/pBYcgGsusORrDfs4gvyJA5V6CiLRetU+4azui0PF2fx9rquwFMEgfcS/5pPL
LliLLnOlFEsVnNfpJih4AtehfgLKP0Wd9mafQBQQyeHcqayESalufn3fjl/CwAWx
yecguafCefoKOr4AFhwa54kDSh4PQ/oWMryeoZhcmYyVhe2mbyIzba9tzzyMpZIP
7+JHHKj/kWeJkQptKC3JDJ3eB8qN1lr3AFWAYqhq9wpzQQeUVcfaKyRmTb6QdMBM
6T7rvRM3MPaExXFiXVtxhdXsXshW/hDpMuQ/o+XZgTQxQRfYpPKm6HPfhgACIXky
wf+/fV91toLAPd7jcbQV4TAUjMR3GWxbh+lE9ffv7R7lyZFOtxVFtg29QpUea+U2
y75n3q3PetVDrXUOUbc5OzqoyHj8HfxV0iXW6DnFvYlRZBEwouuDk0exXmIHsBZt
j0785hl5ic9gx+yyhLo7oN2iVwLWfKJUV4zetKLkG9+2RoCY4uzczd6NFUwB31/t
suChuGnWarZAvT5nLWvnr3us4slYx3B13wOA2A1GiGsIuyIEWlKcNkACEVv+DUnd
BSXGduLCQfR7SuKevpnZeHLROORvQPqyZs/UJtoV7p4LbsOZnnAMgpwFJWg4ZI5I
SO6vti90+SbaYUDgbeWffVDp1hthunT73oYmcC2WU8aNKprwTDVu8D9xPyYPO8fh
ONxdL/Qlfs5kZMYd1XT7bMxx8s+0DervIUHl4U3Lm+hPNBXKBgJJMmw3uuI07Me5
XUzHPomsmTDoKAVjxyD7uJZuyEefL5bnrGGxCnAAlq81X8CJ7xBsKH2vm1S9Dloj
9QTdzFiuP6SOPDKPjZp+RlgEbpzptPcOqIyHsYOQ2hqj/KM1Y8NU68cVprJ2NhOC
h0wfY4qZmkVGsSKANoWd8BkW3OlzkAwy/RwpgUuKWV+uxsH80N5J9ehrqtXI9Xf7
1OW6VDaUI4r404jZwRBoalp2BpnSbkXWV7aveFsIZntFDnOADXmCt9t0E7ouujDY
PRA/TqVo8ZSEA6IVqMIRIoW8tho68San4wnDurgQGxLdDGwwO/BmWFK+1UMP4Oc3
fTfAH6FypAQnRBGXMK/GGKmDpY55HTMPA6GQvb63fx8BIcV/Rffa7rcjVlA48TKf
hAWSss4BmTCzaVxeJUzh8veSZI0KS1/NkijVjw5SVJ1NTq8dXypfp//GNCCO1Sc4
1FIoeUa3CdieAknQzBzFXIYvxgg/zCCeFPjUf1oibSP/FC7Hj5AGehlih/twSRVd
13cSLS9mfgeeRHoSuPGQjocE0EskvtuijmmBMruj07wgPz4e1x4ee5RJai03lzQJ
RaB8cFsrAlIloN3yw/cxrIrtLUSwpZiDlqEEFhQM4OXg9hXEndP0tuN6eXniSC8k
hgLMR2pWXmVrSTPHB5Isd4cicNiz20y6kx8A1JCjA9RnybrQ/nbGe3l7Dx8Cq4lQ
YgdxatoawRkTbOW/uw6iDpKSwV8t1izD5DRGLRG2+6zVDLcqoQ+dVF3dU0bHQhLZ
Cs8ALTJ7aDxjvB4dTRYV3D6mMjRllD4VlZfKiBqBZTVAky2Rcd8H0yoDe5J+3LCy
DAxoFRoh9wWzw+jZwLE4LfBGhrl01+jipd7adrC00PRhHXI7FmfRmaLDT4PTCSpU
5qnC+U4poXXaeoZjNEorz9IsNyiIhtLCQMbAp+wdxmERlJX+UdrupO9wxATFASW4
mYTfZpwCzkzoCp0aoNQBME0DReydYiA0/FJ6JzAuikjL2PlPpcP2vdvmBOwrA7+t
s0G3iWRP5n9zlb8LMfGuIrqDJIsE88/8nB/xob+h5WIP2ALgmRVvG2UXAU7MXIJ2
6FUc1yCTBgI+yBdfKZY5BO2ASFhI9ZSBsPzKehZE9izMTsoW41VB5oz1T7b62c5m
hNp5/dvvH38ePhMuuIPaw2sbJDKBTPkJNbD2dozDABKEFqJPd/eUFxAz5l3XOy3v
vzCqdVM8hwa6QCMe3FTq0cntcZqWIVAryZUEPCCVjyGQhMxPEdkKEgfk6OSwfEdf
BwuTm+RcVmn/J3paySa5lf9bQsYc+mZCKdvvpW5LaCNA4ySf0czkBJfcFurdTF24
Y3GFQtuUBNzghjxkPFZwGwYvd75voiC/8r4IAxEVzEJLdbyQaz3cOYReEakNLlqW
VaiaXdwb2Bb5tch30ZNUT/ZkavI75BxZNTxtnqpX1FV+HqaLEeWQQBczY5PlVdno
xvPXbZaiV01tyEw46/EayrQSPWvX4fmdEiyRfVW6HcZH9qiqHCnQEAmlCpbpaxbN
j62lVPX7TDKp4/wsl4KuAs5mE7YYYeNIQ76Xp1fCqCBidBBcZZCmwNyNmFN+hEtO
/Qo+DMiJDsTXDyZjzs68S3THGvjGw84GSCIj/lRU9xmGqw40s322Cs/KGXxHpedf
1MaAxS6JIhbfwdAuqtFsNnhccvR0hQ5XwZNsIaIq2RM8pn9rvGkx88Bo7ukt3dDQ
660bxFYzG9qMfu4d1AnSFvcXK0UJWsBW+NTGl49Dt3IkEbRlNbxofOsPOmFHHqQv
W/rlu+bVpPEtyQrKfbokEZm2siGG5BHYGLpcLI0d9fOytREkyTn8o0HTij269+vY
MFje4KQ5+W86SuE4neT7cCp00FSgEZRq2NQlcgDCns9+wA6ApU9G/pf5Gzh/rLwL
nSdlk8f7cCGTvrPB5SpnLHKkyXFO9h7b+bbIUdAFNLtVP6J9hb7LtdQ+7AxTBBqd
6RTKKUzFBpVCUVab6VbxQJPnkHPc4j+jFAaDp2pBXSrkh2ChdpJzKsJwVnRductL
1knMNQ4ucThegyxztpL2SeFoXxiHNf8ZMKRD0L4k5qy24tNI0JQQW+CF6UyzqDzn
2thpS4Hul65fk7kXP4qHOqGXPWSWstHymXNLhbDCrvF2yYfzy3RZUm3dvvoFE/9y
RgoAG7uMwCtf2UoO9BeWIIrvjVOrpPqVuHfUpyyWAVqdpbTJ56XSqxyHSNjlVK2q
2x9xKAs5Qy9SFkYSQTgO1DRouQn2gA27wDwcs5wMx59D1OVTGs0OFqjpd8LZEbxw
oA/yRs0l7yuwMOVt+JCBEFUm1699BLahpCfhgmEdkdOyAPMdY6bFfiFJjk4AVZV3
nKLyfrxCxiIo3nO6rVI9S+jXk07A4m+S4znB9MfAoxbfwJnOjpGU34r8kYoXkImH
2zjzDQ68tlZzHHOeq/CP2vJeQyW6DMIwqRScHe1GvkAMtydqcYhAivFaL4ytCuTt
uOdt+qdV4M+8UKrwO64y1WllQMvUuzuBUONSaxebVNwM9F07SuWpQQXo631Cpq/K
sO3gp9yUcHW4AYJBEhv0Hnxf4zeVSg3QFeLGqP65KI12U7+0ir7DCfZnGm/sjdUj
+qeMwwIdp20qkteTAG33R5tUqahL1pnDwy7QrXVNOyPPxbjht6QNwu7d9yS2zPNa
xquh2qFadlXS9Yv6kWINXFBsRI48R3zvkeBc0uSgLtE3qpPrqAnrGNw7+zQFrGBn
2Q1ZZfqvtegcYzFFGOXYzXPIDtsWRmRtfPU3/gXwUrebc6P7+vDYt1ubZbqcsgS/
ksyHweHC2pVjd0ben9Qfg7SQ2ffwgAQt8iYOgAKeafm/hGhSLkaMEqp/LCGxNDan
39mZ6b3ZC9xPrsLZOdmOPMSwcslzBbBdOZVwtzHFlt2U5AS0BlNFETIs82LNpdfJ
Cife0N79EALhxtMzB80DBIDtIxe74BTpChplmFmbDprQUdexBQrw34I7Kj3St+Lq
T38s0Wr5bxpl1WsrxQgXpUmGlYGYHoWDlTUdyJU4sds0rxEhBtElIkrYohnXm1rH
eUGdnr7KEkafkAkL4z2arO90MhUek75qwwJwQXNnIvPSFnHpEidOdcQZvKqbm3TZ
dNJgRQY1FDBLXrnPc+aD0rxk+3kL6CSQMWDaVMrlP5BTb82wSk+LHLEnT+XqAqTS
qnJ7E/BcTMvcVYpbtW2lNlra93djyPf1KXHuDCQZVaCyBT8wNPqX+CziEEEXQHD5
24JAFV0CjDz/sXoiYvPUpoOuFdnP3LIcD9w3RRruUvfkQ4+aWRvIkF5UOyRAA8eU
Bf+hmNMcbPGSmOId9Ykz+Qqff2bhHLu/dEkBhO2jCZzwqzvnfwGSsKkGXck2iaAw
Mm1fMzW160QJrziKEianDTw1wi/x9OYrb5AnbO/NiGrvlfY7K/w26rHyrrJ7h/6p
SKwe2qwdcgTR9kt8PcpJ4zD4KZHn7O1TchwWRzRCatIF8jOCQ106InU29AvilUhi
1EqO6sHwAxraBGyRuBrbACdA8GKoHAgLl/aIeEGFhYNxhopuOQ4jWb6HH63/y+T8
xCQLfKCRMIivC2gJRmDYKqrkAe2yBKyBxiOpvBeQcrGHGEuIWEwSrgWYxlN1eyf5
aOtP5xQ+ClM4FBsmZVLGo2HVaCmx+TF+Jjp+R0wxY3XONBZHVP/zFFI75yV5YhFJ
8QOdA/v1T7n/01ajswntNuK9+GFc70Qx6p8PGvN1ZpSps8VOxzQMELz6Rt2QM7PB
Y7Xd38bWHl+xddsyAAIl1kRMdVkUp4lmr2teq9QlEgrNWab0mSK+hfS8d9CIJNsZ
4HO/7arQPsMFMOggmonhEC7kt+dnAWwEifgSyPS9NxPRhpTzHr1KzrC0WF0OtSCk
Z0tLR8m5Mlr0f4xx5VOc5nENa7eXvuQ2k1kPIFxwtvtLxOqu7djutDGtrBS8LdNl
H9OqWIg1mhHj5W1Axjg/VlvPlBwdiRExVJzwEEnUvhSGmYhy+LlgTY68GNX9urnZ
NgoGBy5FbHTF7ddm9UqeBOhtfK8XBv88YBn6FOyLrcwcplb4/Es3cgxqNBk1AUrr
s4Ut/9ar5fH7CNGAunDFV7D56077GxEavPw7ybmTpAuR6ilcymQeMKSDP+mxhuFy
WXTlBYtZ1X5kjH+IEW7fIQ+/qpfqJtWBDIXD8M9CdkDNDX4w7MdEcSWtyXJSsA1z
CnUeNO59xf0pyGXG/E0LJHn1yF+K0z9hyqFfgzmST+m1hPZH1IvYoPyrtIubfxQ1
3Wa0EhDh/vaYlD8umbBtB4Lt8NDkvdjCPEWgxk3wcbcJYDTl2UFcoz3abXsAkry8
JrwZhbJs/uqaa0s1OaYu4yXrUmK/ggFW+Ipg1vTISsxW8T2zQOeS+YnK6d96JQuO
tyU0d8hl9mAFDcMEJC8apZkMKeFXjl513K7ij1EJzyHOz/I04Zh/174QgkRwlzcC
mBlbaCcmviSKfWGyDYuri1fsLQYvhtCMWyGvd+8F0X45Fw5oz9UlPkd9WcQHgGcX
7UXCDRuaDO2mZNN5BQA9KK25B2jVleUKxFmCmEtf+Hxy+Dd5ID+B0wQobS5Jjnpt
qdM+mwFtKByAFso1uP7lrlSQj6PtZlSMdjMOajt0drgLyHIGgVowUyVMrD8w6FAs
zf5yQC06vOGMiAM6PWf31joeuKeydGL1eH4ZgS4n4erFq/5bKLXKIfTo8vYhmgXl
9tKie/PkCktFiglA81lUXUxswQISv4CDx0SqMyU6qOo42NPfO0PQS+ge+VNuM0Lx
+UVne/e73Z7OepaRALce9XwHYy1WOL8E+Nb6SAF3vfZka7hMj3gfXQDKCEZiBWea
dtPmJVlMCs+lXYdGiWNKPyTmp5uVylMYAajCdeVpWCEbkcIsHaZPJQMZX/mkrdVm
NemH62gox2M/RKCnzYGAHk48FI1CA15r2pfL7TJottCF318ozI9mi+ILWSm6jfUD
uTvPMjtu2tXSaxP7A9SpXlQGaXFQmvX4BkY1eDzRTbQXeVlp1TXtDryZbuzy1LpH
CpIifAzsTF4mdldQh8UeMfKMiRRCSU4m2bXpLnufuA+BbfxPkkndfdhdjuIKVTOc
AOHCAFn2TPvvei6G6uWyitp/0NOG7OuvFVOO9rKSWD79NlZtszp5yVf1DpOJS4tv
qESKuWdC3reE2mjLghLngFXa3una+cJD1fFgzgKeONc0yXWrEhCrgj3GBJTcwJ7Z
ygCibO1jzAWm6YkbNwApL7x8zELGz2mspgjabMrxGvfAcgOZfCYYSFAInN6Tb+IL
3u5qdfF/KOvGH8yAdCH4DJdLKorc/Ah/pxNcHzmRHm98PcnqADC2n62ND7HFnLwu
5MxO3TWlIrgzfy0UDEVepMusojqQD+J4s095Vecpq+C5r1GLN/aj/9I9RvQgUdfM
IHVckNTToMIMOxNPPTRsB944xpwYoJEe9wCaBY1meDFkeCGiaPmsR3LDxbLMvkc9
FnoUOYZOHUigFXsZ18MoYsx9eJltMCwW/aELjQPGFGvooIG5iGOPEhq001LTtKow
vKtRT1BjfdHrB1ou/6YwtniH/yhSaV3i5cD9SbiXqPQwgyBM33kr/Hc75U2Ttvp7
re/bhqU17iR+IO036ZLjSmqzWeenzP+R4WIKoRhR2R0Safjt6tenKMHJjcjPzPOn
rlkXR7/dAdHt70rZQJUFXwdTm/cq8hu8V53oB5RI4be1OtYQ+kiZhy3T58c6tlZi
EAnl5jSpr6wrc1E3IDhC5lEpJME+/Op7HBHX6go+TxBPbb+Jbm0Q+xNk++QF5R1U
MY68pG2NrFKIlbTx0pSwi5ZMGpKbto4rCRPSczq7beL1IGfNqwe43IyQgovbMJiJ
m8NdcXItqTSWFHQvfyJR3a0FGvi14xZsVImxVvkOdMECfzY66n8mPW+cwRV2wEEM
vaae5ZGOt8ANYF+Uw1oYRutXX7lDVZ5rJAG1lPorV+6a32cXaflm0tkQpnwe7mWS
tMlNDBEVUPi48xzvqnPN+KK9Xdgd7Qw6wGOOUYzmvtFXri3TNdUOeewV2U4r3bJZ
dqGDUSyHGO975VhYRZ4ykmfUMDwm2BWqCm6osru6nxGJ8GpsOWgnp0CXwAi/Jb+v
9p1cqNKfTUeDhH48NcJ4zbJn3RcKTmg1lchRY5i1wIZ8M7C5LXwTQlIr7eWIe6mN
wNNwVfNp3Cizm+y+pPVWGyBcSGOkIJ+4AGK0xE7jDMjDbaTyrju87uig5oCnPzAg
gsUt8YSKaYb1e1EA7tPSRUBBejxxzDW4k1/vX+9RYsKgHdyIyQqmAgul7A8tg6xn
cP3Ftd+mt2zkAjHTwliehcMOK8w6/tkdRAmGrjI2MU3PLfGCtxT7Ix5BUF5V/epo
euqU4OAbra2/toadSItH8nhmTIBxP0J40PuUH0AAkWf3zqseHdbeOzAf+WMtEehy
vNGZjnLRhBS+wMv9YIoNDnxiUKDBqFP9Hh22TGOtU1mkSgzYm29lgRgFFZynUsJf
gzb7BfS4FZrNJEjS3UL3XfYL0W+czfEhL8e6zdo3R1wLq8YBx1CAOcWuoeEadSKG
YoyABaPL4Q23jU6LK/vRqkiP/XYuTSw+SifXC9Wp98/umghPD9GP/urDAlFjbwQp
u5GKzlauGLjwZQst/kw0N4kHUoI8TPIVk7/YH+w3TchiVTFDyNQTexw9vR+kaAvl
BhW2idGphz4o008qPrR90FDNiRMy96xXtCBD2paO7PBlScMYjhGsGofQwQ9Ukmlv
wFY+EbD79Dqa5SuPUa43aUQfUuHowReB58YCG9EKcYMXH/fMsrSDmIl6qCWQZa62
G769FfMzEe7azcCDUGFpsqK3/nFNrhO42GLUuFubomrDg9a7JoEmQyizfv/CaNtn
tUCEUfADrd5ien79KngekK3zYPdHRGFbMxqamgjve+w/utis0PGeGaB0qrzSxr/g
l/kTD+wx4GHEbiYAf5lDYC/dFTYSNbzgR03umymXKQ5DIxbTYbmw7jwZOutieLUh
bEBcfNTFZDnY2tEK2QfgMNyz4fFT484x31ZjE+0x2froDRjOBq7ma50RSN8yGzmI
/dAPEpW7pUaO5VGHMmjLVmWZSADL3DFB5+umX6FsFsSZ+8vmyPoOb4GyMk7f4cy5
ChEVzXPlSBETbo9BEoWvtn7qMzeoz/3kwbIN/XsNMu8lJAvpp7SDIjkEh/W3ADCj
BEMezcFpn9Rh0zVjlBXpplwjQwzteOl9/CG5nuQop0sefvy8YOhghf62iNCAGL4R
91uT2zw+xOLVZEQrIhKsg5Fx9EkavAWBm7WTOdptOfx6WKsTtk4Wn9CdZCfy7hQY
b5Vvy7JNowDd3NdWxX/8k7xq9kIw7F0/d8ecSdzGP1kYYhWBCbGP1Lx5SIfuxBUi
72io6LixIfJYlBCgOfBrNRHP3COJ1+HUXckpPPRFhRaJjSiX2bDr7sd2bnwyd6B7
HN9yRm0E7Ayag8sDtZzfyhL85Oap0XVJeots5sks/JZQ6ky7jZ106+mgPJoLPQ17
leolglfqGUcu8jHgigl/xrtVrWYwrzD33IgMuiLHc3E2rLU9Cvl43o8MgUbrjvYl
PVE5BEP3bAtlbrp2NIiaOLWiaS2oWAdnN9xt6lTjVqCI8oTBZyWKASDm7H4Ps9xp
Eas/DOMU1CExXaXjPp9x4SdkYxuH/e73dQ8sbC2L1vqyynwwrfx1n72f2VpVsY+L
Kf23YlHauyrgVeEwNH9YGx/uBcAYpA1wEwsfCf0KMue7AY0A/40Nwru9jeOCtp10
ylTDGTN61RMM4/SCye8O0yWurXovPT+JVFhhLF+24p0zwjqQ632IP9qmfoW27d6a
4/Icel9gPjVjSm5HiPuBOiptYYkgcvfNOGYQtou/casgcFYpNSHPyhTXueoW1A3z
bScoUDWU25AVm184ZsbuboBdyYNhNi2A/m3rGS9cjOrcDay1Bpiffx4xkrN6v66F
YZB7o71NkdHQm8sXtl11xfbB8p6U+xSgrMF53PBW3pk/VNbtj1QyqP4GoRKViBDd
sBsAF0vkSAzVMNNIz1dGx32H7LBjwf7ryzfoszAtqfrBkUc8LbOZGqDVfZN9jsSJ
rVsmGRPBp1JUso5uK5tXSQDroki0wF7OPH3x7M78sL5o4RcgPnjBj2UMjJFn5WA/
Tz2WSeD5jYlafGkQDHTaUUJNQOaVbbYLueOs/ONCslNDPKQ8z1ZNoF3iy4O/5zPe
v+lSjV/93V1f9nijdVGJZHKFlikB7va+6vU5rYxILKEJ0HCF1lizLiUyRKWeCQ1z
kgovYGIANwibygZLQCsEWKZSKCD8CEF9eE3l1xBW1WlQQO/AfO55nNtPBsVzoJ8Z
u0YMtGDvNaNLeoWB1IrhRMCf7cg4mthNt5hvLZ56izmFBC4G0uNLiFi2qVLPHw1O
9M2vJbW830tgsanfk0UJMYIfn+/4WDQXBNC6ML6IoVbwTION7WNpkefg89YfsBvI
k51xIuVrTfWTfYG0ONFqgXzeYcUdbHgHVoqMnW4etaq0grflDBvREvBwMLrd65EY
br61PaUGM1oCr4v9xom2JFDVXA+9nWLOWfNSjkSPrJGCK9s1wzbnv3JDdfJzlLDh
2PZ4tee8fvDUxybJhCiXSHqnxcknR/ye0QjRLkDGo0Goo1Bzzt+q+Nc8HDvj5T2U
1fnHoHifNxP60zFM06g8BV5SGCQHKpJuD0phnRq2CbHW2J4lJFjCktGdlDx5MJuF
nr0RT1A8X2Z00eZTMQOWHe74RnZtJ3j193xHsUguc12vPrl0js8LSAp1mjxjU6N1
XV5finKyYdbdiAHFwGe86EBoziXImLaUeACzXrYzqFfuT7GuZseiFGFhKTW459u9
zdynKYS8hxt/ZiOSTMbyNHxt1mlVq389FPkYOXLzOjxUtwYw8d6JZSHpiqPy82hQ
WkGZxon/Hqb8UPR4l1OVynG5cubFXOU3WZIowkC/BWQ43LV2/dbKq+1Zmeemvfo8
HiGUYYpvTwoLCUrkeaNgTcoUATPgkNrhStPaJ2OLeT6lfTajoPkzsVf3rqW+C3N9
U0NF5Tl1drAPuzbxMPfEeZOsBWx4V+oePHRawWhB13r8n6WE7F//VD6q9ndK8oJi
N5uuK+K6EhnZr5vuspx9ZlNvB25DA8SI+b4AXajcydfmRy1dmxMfH1AHZsaJFxVS
jSYUOdNDXqlUPQQ0NZBWFnkt+e9x1it98V2sarHjvSVQfSYJ7Phtm6zDJo26YZLt
9QKeXWXeXnPu2fl9BqbEXgewhsFqm+cX2z8O1PYuiLKpEsyvq/Rcn2yWYs0bt6pZ
jGVlsFlUPtjPnfb++TrDED4kJpeb8q4hYGsJyu1SpJcl4l+B0ZBEcoS6ThuZ3NvG
N4PDLPLbEU4L5DkHzXkHPzp/cJTwdO28FqyoeCoUZBwRiX3rQk2XWXn/oUZtPz9T
FcIA2IE1fnq7aktrIFJTa9lnvCxsV7/2zsNBgmqSahKpSIcwEBR9t3hBxfqtIxFJ
axBmUEIH3OM1OG2hAFj96gv5zrERTm1K7ujnjBsULu7eBHlht9sSHUvSIASQDShW
YIm1fCCpmRNZbiRCTYVtLxoYzESWpTjE3Hmw3S4PaVNOhuK4d5ut5tsgfu1oP6zR
GGjQyB7HSPAPmXIXa+U3dqagonan3QRVkTMNCaQr6yoEPyCwPyIk5j8gR1xlfhaW
raPU670G02U6Rqkm8QIKyF426oDUVatu5Gr4vuYAN3ITMEfplFEFBvER+ZGtgyZf
uyp96lWyDU4tYrXMd5eCMV/rjE+u2MBqLKTgh/zaE5irMClx05mJwEObfA9Ix9GG
5FamsTkspG76DgQce0ZM4hqfFNAUU27wfa9DtlAC9l16c1+rXOnD/YtDQLVmg1MG
t34Z6AVbUAET1hOjRy/uEw8x22Itei686+5Rr+PsCrBXU9PoBFGQkW77T7NOfGKN
GdaXSnpqv+Sba0xsbaGbMoOoI+PjHH5gfXlDljdoZ9YFAiqmPsztJ0fzlz7YUcYO
3NKfy+2Bz7ASGAT+ri1DTDBNEG3FlepeFBsIDQYkuoyQdv7+r+23wFrTaabmtmDS
xh/CjogiNBwdW3Km6bob00luVAfuoBj1NR1TPMeHTPbdPVzVddnCnwUpMfQFPtQF
1qWMEvGoMp4891P5oU30ZAzuXH2JGMrOnFcGcnex+gjzBVQN3GE+IlCZL02U/UTj
slCLcC3BH4x6kJ4QItI5KFqr9Bl5L7HwXN1yYBiCuk14d2+KrrN5Uj6YEfdJgiJM
YMJyo9s+6vgJHhxTALfy1pqZtxPPHvB72t4yXbf8eqCnEKKW+6gLd9/43Yo04fyU
kJz/Qlnf1Apu/DsoS7A7BF8mDV4CUvBe7jDtwup+oYT1N5qACs1pPmygD5iG0Mni
FSC+a5sOp93gAnmb2RNGuNGhtjbrKW1eBnmJSCt5ApN4kmDLevgdvSlNW5DoFSd4
0n5ncP71/QNgdcBNepKuRdMvU2FizyBjmuP0PbZrsHZiW0jxeG4y5xiHMNCZypNx
p4mUVhAc1ImOc9ZYGn+HRZl28VNO/uhLgNBIWcWeMXYU1r2nna4DIAmdr53xLQv1
5KHMMdLTQEabi5wXAcTUZiA+FNLQ3b1E1Dst93PJ3k+hwwkVkSQMK8M5WklJVzRZ
Ds7HebAAysM+kZ7e7+zueurpHA0VXq6UgymD4BJn1UVHLmwmdtOQkS23cJyQVoMm
xLp2APzV8SwoEqKGnsn+cWsziruemyio60viYeWIQk3Z7BGSTjjMRrdXzyycHOAm
qdU0g72OYzI2vDs262TsfWpGc1pwGMxHpiW8KduOB3XBlBvMH9UclnUHCC66PKXg
62ll38mZGsB+5ZXUrb0K5nLPbcoQlR4REomFBEzcTMwTrLB291c8M+Sf/z/KIILO
q3O18WrWv9GzJyZqpopvrTQjbI6m4vr8fWcf2nFvkk4ZN879nyX5GtIJkcob9ZSc
FtHRkGez4F4nplV/6S/JWQv1hfmBjunEFOsLFv18+qPpElu/hdGuVuwd7IEEi8aI
CjYJO4J8B2+MJs1PKyyvDWgZb69h+ndXf0AsBWsOCPzDzOndDsmA7abANGHP8+eW
KHhHCVTS5ab2WRJPgVf4S/sP7MsJwDeE5CY6p347EZBddxiKbP3/2RLYHBvxhQr9
DAHW1INM/BPi84qnmqy34CV0i6yLqH1qErDNCdBvwluVzf/AxkJ8IGjwmLkqO5xH
OPmgo61eFQmGV0+1Koe/+jZ7U2Jnm6l6arsbQGellArTeVx6u9txbD/xxw/e0hw2
WnEpt+iB+l261ZsodSITeVgHsjWLplnwTPKzXHy/R5l1Rc/uJk9cDV5Ck8ebFsYs
yf0C9xtQFbNR4lTfWFxY5yukyTnba5A3/EUdBmwUoZyco4krw295u8jiBVKewqqD
4GxdqoegNhzuCQ/fqd9Ilht8M4ve94Q6750XLEr/qZlgq93mNlv4HVAjOpD1jdTR
e6KYV6nNzExgXncIhHfASCUL2RwvsY2u8ivJJK0W7/4+/Ex5MBuWRzyGQ9MM9iAN
q1ckUT8Fi1B6OriFsKTPufiPyH7TDJp7VNmIzBU6qm8L6Ql0Ev1zmCL3Jzr+9c0c
x5eHlqCg4KyGc8QHqSvxQq2xXzf6rZC7A2Le5vmCrtlcE3w3cqxibhslsW69doMa
Xv+fNTCz6D+IfLkXv0Sm1kfkZ+BYlSIIItHJy1yuh0p6/DSOMBojVMFwGTCoo67f
I5zQQmu9MnAoTY8acabk649Q0GONwlo8KxpMsAPJGnQKhS9X0+Yf3zrGQa+EhPMX
RxtzEEQzkn1ekozOyW35JvDFC8fwpLu7QMHgaaRsWHmL1UrB4JIWg4/5QyEfzbvy
VusyI/ICFnKDdu7RiaZDsCrK1M3Aezv2MwI8W02x/NeFRxN3RPMRHtbCNYOwDsQb
Dn7qN4ZhoSzasnBJRTQJ0e3uwIVBZmCcrgDdIJdfxRVme/DOlvU585jqzicnli3x
tUKlnjFYpgB2cv9vGeX3wioqK05yWpB2JjMrj5icZhiE19WNGfPLuLsCbQ7DwLSu
/ShgTkTB1WUBBzWAntNuen4tXeIsJ+b57JYdN6EtHx5Y0bSmQFW40C2tz/G1uUig
KY63whY/DOEW8svUpC6cbs3d0Ca6is3MARDpYa8e0mul2KPcR/FpJtVBmUUwIrEq
CPXDsetsIUNDzG0CO6uOonaFAr73Ax99lZGcgpzlTnfoXhR6rUlWZIOx39WvyT+t
f3ag6pTLeft37ioCHRGHYME1hETRuq+abgCcQYX7PElg66Wwr8ZKYY3yb1Q7mF/E
QuS4dmc3qw1XGpIO/6H8dnPMToyRyxV+mecbc4+Yy7YKtjyITzyHY+Y2lQC52CSq
GY0NMyjfPmG457tblSXhFUU2XF9b0jUN4h3L66T65SGl7Db6OEjYUnza25630A/U
o9hJs02VVnVwQSiEv3ZSEGMoCutyTq74Jfh5GnfWSVTKY5ZRoOvLbWwfcBaD+s23
YIqu95RuwIG2YRkDEk481KYuQvLxzMTrPiOtsFdz+5uuPAAdl3aWNfaS3PXVTskF
jqTHvs9KoSf9cfqwEXjRkACPaq1O6BEjOMMNMzXqMqMDxK4I5HVuXob8NRmtVz/O
WtsfJj9O1l36ak0NaSR/TwVnckZvrW/ySXwkYnpEOK6sQDa/uIBlKSJtGxhj697c
zoPlnKVROF8Jwa2Vo8HFy1ZPqmYLgQwYI5TKHxgjoOvpfFt5vLXRSfsowa9NAH1P
8zUR3ku4PZ//NJacDTcidK1220felhH9+Yy7MeEzgwzBZR5zTHtZDuH8Q7qYnqfh
gserJpQzn04HKGDiSvIqfqfsoRldXNSVw3ryAFLXN3AsKP2bZqaHFPeHZ86lBzFG
+3/dawJITCTxVhSLwZjKYXGeL4BBfcdmc92Dg+E8kxWTYDTpPJ/rwkR5c3beQH0o
P09p9bwoo73nxizrU2J8zThlWq394H0d32IQ8F4opRpt9jphRwog0hPJ1nOX9ksy
y5wbF6xpJ4GLWqXm6+oi2D+wsHSSxIrR+wS9R6TgcGAe/C1CZeOKczZmaJFhTPoY
FajCPln5wzPtNOOj0udDRoA36IiFEhEK9lXqA9BtEOo+aXxHVM/flRYsHZrC4ORQ
yt8+d9ZMoLvQD+CV8VKWWMjGir6VuVJlPY/SUNAbbY6u9AIGV9guUJ8doRkCU8b6
PrFfmS/KKfWqXhpJPKH5NFahZRPSTzSYzJ31yUm1zYqVeBRCVI2aCAkDAsuNz2G0
+yEFpeaLIKQXVAlGOdL2Kp26IRwNxVnTi00gT+SCyPmfvaceHIbuOlo0TY11Z9aH
fOr9m3yqf7Q/bciDftDFhLvTtbNkYeFdIz9d59aMeWYFAoUCP+/hpYocIicDhPBu
qza6o4HOgon/HV3pKn6XBJTZTgs+8gPYSzkEErnEQVVj+NKIXTNBvii9q+ce/iyD
z6qpvc+Hep34/q/3xTDZH46mYgVWvUp5TuoELmItD48OD1CRMXJES2ZPnVqfuzes
dX79EPx6pWJv4YqktPSz4BbeMiBPLBotOhdXiILDmjfVZ45WbMDUkdS5fQrw5YP/
K0L5/IePgIdWDr7Cwq4HG7ZTPNk2snB8PZC0yjjv/tK2QyO5/1XzmwL5KNigW0fu
PxCm0QaxDRB0akFjAY0k6oTdUGOLknEyxOjSUhL8v2+dUJbhkxiYXFPRTg3mVUTu
wa6pSVz2istRbhUkV/PuqgmXDzzmb7dRiNTOnaSF+UuOYbIgSpiZT4Pt5Ud29SsD
d5j1W/edS+cNVkVI8n1oybA0ZHSqGmsjm/VnASeF8aK5CwPC1IyNJ4Q8A+istk63
34YHXNoqoLR4g8efGVo7AO8bt+DHqLBHPdeGQlvPG02fyELX8i0PILDjF2qUp1b9
5Jd6cUr1TG06yz1C7iCJQAdQT7lbdROiw19bAe8elXRaci9wCrZ82uIMRV/u+lNn
PdG0tIq87wwIg+WSnTtIY61Muzu1h0ibfm0xufshyZYctA/lGJVAawV9sxCggCQq
1YcHYHS0bgPhJOIjYqEz45wRgptC7JnaDz0z9vrS8agYgzEsfOYML/LW5JuDMuz3
cDAS7SSneNqeQMjniqC6jY5W1xg+kDh7161I1yZXyGUbzk+9e/2JxeZ56gUCPp6J
XmaH9fAoprVJCjFn2+W08h2yLApUF8J79aQHLnlJaq/9K/pSbu9Lfw0obCAopPij
YCT/p/0ByL8JVPpaZcWUapxUL3F0SK2US2sMs6fsbF+Nz5728EBRNCZUOY5fIbWV
paRvTODfXlN3TAsqN6s6EbT+hSioq4CmQdJqZO7YdYOIJbll1DSqnYxfy+G0YcYA
DcU/AV2v4U1u+EIaZkQ60INgEzJJ9xZbTooWFHzb8AXE5Pa+wptRL/tUpnt1qQNi
sW54hxmzW5vfsQ4fn6LDtfpvlTIF/Zccx1bArwsSkpUKV+Io9Yyq24IgX6dTlq7K
juQiuPHvg/QuMtpnHZsyi9VsDgFnByU/07Ipe0Zwp9BAO5FPwbyttKrXF4kGOTcC
AkSTEate6yqv4ShYtQFCXvXVCNS1BUPjldL3yrM/CMZwyX1zcCZYnLORh3rpgsqm
19SSL32HPXzLtI6MrdkB7TFUQA1NeI5z0gLy9uVaFCb7pA9dQQW1/QbpJGcdPriF
pmHeDvgm32VhelbVsC3zu/E0VZJg+5qgbvzjoYKySMc1FZAgYht7EDyv+Z/78AdT
2lruFOujoPBMED6aVX3l5bQC/QkG8Go0bYufCVyu+1ICdL3O82fVahG0QKez2CHe
nTlemfrm6x3M81KJSKyS6dgVdio8i7VAfkHMutza6EqBRXqNVNUQzviB9qyfDo0v
ARtwinxlXZKUEumzC03tqSdMRnAEup1Pckn0MMDHOsI6Gi6ZRTmWtaaqhNH7k03n
S8rqzPwBdLYn5XbAlI0y4b7sRM5nZIMQxbEqhrD0uY9VMNPn4T8bG9LXgZoIZFms
U6W3iurxVnH5fY9/VY9/phGHYWSTOgV5m6uaElKFr667K9UNzQ0RFwInWkkkTz54
kR8UgpHLzFf/HB+lpq77nBNKTuIeqbeLstrmTjwPOHrF7eJOehIUJgzVQEYU2pgy
e9sy7RAugYhludrU8Mn5c3X9aQ4mBN/DWR2VWXsast2AA02hel6XySvCrVlVEnMb
vhca/ay24/zpX2Pjllanz2D9xqH11KQvreQNK64iJe/2AjG6+UiWy5SwboZycXkz
Q8F6V963bHegx3W2j8UvjNmy4+9s5IIU+xMcc/mhGNCnmZ+NFEpMWbMqs2WAEdHS
2ZWAIGrdeWBwAAta7DMTjWIQfXYxrPIK9YeStU60QNXlwTz1UAKsWlkvY3VHlS1j
1IoGYGJf6nJTcM4d1okBalZZilGkHw18JFxiUIqSYHgOktT2STdutBWcFaee7Kkl
H74jyPDsGLPRkPJ9+nnLAVSdDs30t2yDKS/waTfiS2CQPQGpRRen+p+UM2dSgVK3
G6asTRm55fN4yF/eVNcI2pNyBHXDSFq99sokduxHEQ9kfayv2kH1TGn+rg1DrxZ8
GJxvhirPidPz7dXq1/2gZ41Hh07ZJjgIV6xDPfyNMj7RtTqJG39AZfJ0ufErhM8u
6kweOC9Aa4wrA6BsaPMJO3/7xnTODC37Qkwnqd5oFDaqaeHIuPfPNhWrhNyBX4WU
jPQuEbCO5WnvhRxFZVSzxpBsqn6zkBHkwwWwl54ktxW5OpHPwBTT5V9nyuTSlxfS
AzbxLXju10IIzKww+n84MJbLZ6vbD9rBxos8vv7ktrLzHa+pizn+2tGwHQDjMBsi
j6jG1PSOZOjPrfP1I0egfDoi7Eam19cG8TZsl01IUNeHexX9ldl9eVgnqiChYSOP
p2zMtVb8icpQGBuy1U6Vn5RKujdh9d5GxTUJuvjO+AKnZ8MVgAmNZWPgbteQgTJH
nBdsyC8QojrAuD3MjiC5T6Rg46NvVLX/9MNxTa02sFdnLzSoJZSp+8IwaIJmyPAe
++cZzK4IZXd0y9sICA3RH5q6MFQMs/BJ9GZh3EHm3TZ54qJp2Vw55Me5JTHvJXe1
PcrpJuy1JZ/5nSOZyseEjeAp4J2pVurJYzaPQq29OBmGXu99CLk74BWFVAT5JExB
D/Ufm2hmk+59rIqbetHz6jjkTDBq7I7ZHhx1Stn9ts80d7MfFFRDemfIJ7uWc5pV
pqyAb7CKXFv5iXDlrAHdRq5aNWTVul3FpLIXwvz5V3QA+KaMk3B0T9uiKeITYvrn
gooGZ/2umRvTXMLLpgfsBJqqJpXSWlAOxneKYzzoSzKaOkm0eHqf413VCK3fCiXY
kzkJiTPXhG0OVyE7MEJ/535K/N6L8UHWEvYw22/CqgrqUlebtgNmlD5ok0mHMiqU
ylFWBIEYPYVOaV5ZgVl7Bt2sWY87pOQpKhUjNUev07F7HWKOJL+MoLVxmhlHi28O
DxIovrJTrDefSuT594958cr7862cq010NlUk6sw4v773tJGf5RgcOLQkqGe9jBDP
0FszLKu3tROiqs5jNiuWdgIO/o68J8d2ZxuZYz4aBg8vq0rZSkKm/56WIHYH3tfQ
o36c1Jyo9sr+P1eMiEgc3HqLYoLvh3VE/uDq80tD+m6pU/Vlk95ox7hinBfiS9wB
osY/sOjY/l8griQ48vYEKu07RcsVTfGa9LhRsINeiP6YpT4TJxSRxG8I/njfRMvD
m/ICE7ROloORSfSe4G2LAXbjUIYD8kECHfYGbBwdoql+dkfK+P3HhGvMoLt46cnq
V0XHDBmNVZKQCVM+o1HN1alnzfahEAdibHXXJTQUDXS8Eev6jj3VppTtxQy/nTEq
9+tvLUP4Odm8tRWwayWcX+jZuuQsiu4DVtyBKqmwsFGPL8SZfC6SRifaRgmVLoN6
EfhZT6yy30cqWRLPB98CHlANK8NCS7m41xb4trz/Eu908uiykaUxh3TC16To4p6i
gBaeou3LqznFx5UdvEJLmikgOIGxzjrn95C8POT/eZBqoe9ObH+AfBQ8pXLMbRKc
CptivHGpmrEpLM6kMBUTdQIZWUwTtDb3nrebeuTj8oFUEsVuFiy5QCTaxg43wzxk
FLlTLnTbsdc8RCJtbR4qCRylzRUXp1cHHc9V/EhGeib0IsaAhnU5FHrdTu6/1sEN
tfsvkNAh5vx9dVDENxIe5ulenkLpdSbrIcHUMC1aQIF6WpWah+cTSKpDpznm4X9U
95a1Ar7ypyL4iWlpFq5hEUJXR1ieyNQ+QAsmiZbHB2cAs0AnSG0orRBNoL1lg1O+
YQcVKFvnpH788MhbgLlm6T6yuSY8FxEyCVWwdOcy7BVoZ9N3jNPtv4611davcozK
aTdtiqT1jEcMm/a0Gl9UUSi3w3v5uKNAfSOrCRd43z2PcD8gPIKusNtS2I0oLduU
IG+Tx8NTIgx8AhUzn3RrKyuNK02JaRAWu4Hb7FsaoQGTxQd1RuxOTwwbvb947zAE
N1bWr4PWuux3RqHMQhL5rwn78S7eZwNMjM3KaKsOwgpD1bpUzIkLTqDvGfD1RCFw
CBCUVaU/rFs3XnBAvCCZ6FJVbq2KIQK0qaj68VGSb3A/kx/hMTXcmSqw7OnvaZa8
ZuLck+2Lfe04eGQlCZI4mTLnUykcjgBnX2Rx8IfHS6EJI8vwH5rnPD+WYRw8MYuV
RymsZvBOyGuvAZpDSjq6uByuD38VQr5f5WlVKwa0BoNR/RAh/U/VnocCohLAb9Nt
8kys8oFffgwZObm+miZyx2TknWSVS80Qw5oGKDgZVLE0+LqH8AJQVoKIP/Yj3nk4
j9MFWpLfFOoD0quF5yetGzrdOABsVCbl+igNMysN3lEiSHCaIk3J+CIxAg5OWcD4
Nbcck4uvrlUMyctaBRNE0HOOBOAHo/2Ykcx4jhyVU8r3MSJoDJ752HfEBMW88jt7
Ww/C798LrZay8DyAObo6QqwhzGtzLp1u39MUUHthsrF/G48EC08ItkH8vMpXgzK1
sc3zTZUzrtSDSUPwzNtdCbBWWCJnctkBAmnXeLpf3zMZMHgnHB72Rcq+VMeaaJB6
L5phGfAIB/nJGBSVgopXMVuqkdfcj3EBzTN144h5lI7SWG3mqDf3E4/zS2Qgy8F9
6fidMwS3zFAMfh/d7eHAEZdRkbnZsq1pzModA1F7DD2q77vG0o+831ZuGGp1Pknv
fCEXjJ5REaLceXhOGESpxkZBBHFIVmjSqVMpI/fXVg5xJMdZ2es+cHAMlHQUIiZf
THCchzmAZeFWGZIylvYv+gEfq9/To8DELGPQHdDqmllD0eIa9XeGgCD4tBf2kjoZ
0bSVVUrVDumQRTHapW1cKTO4QOjORWB3qd6/c9oeTiF1rDa5R8uzLi+73FPQX2yA
R2BQTPn8Md3zdGbtH1TZbiNmtTiPrjZCF4rN8CwIpUY6LBywOLiiCKpJOKF3OWTk
d85TpbtCe8XstBezEW1acNRUDIycfUBfr9WUldZHmRPvL868STHrlu0wRlWcSePg
tmHVZowauoxEOG/0OVDktVKzGsJPo6ITWLZlU3UM9BY05xDA9HV91DAnHv6EpbZ7
tP244+4AoB9GWlpTllMwKAZ7Cp+WMvqV+SttQYzdlzw7dqUeA9nF+1x9PwUG/5O9
STAPJstAepSGDzFLrvw6FOzhHNiEXrwVrMuBbh+gWLJ3k+K4VzEY5eRG1Lcy/bsD
mpjyHNdh7ptzrVzbuBncHBZNdlBLPAIYklgh4ptzoa0I23dBMzWyVMExpvZOgny5
EvSDvWJK06C940WxUg3M7S/RpY83L5ymgFc5Pk+xhBe2GD+pwrGNsMsi6EIiWd5t
5P7ktTBVSASpjaK0c/DxNlrAN948fGX1HNxC9ixKOD8XXj6ZZ8CPjRqtjzg4m9GT
H3WFcGp1SxS+bd91s8ysN8X1z+PlStJVFu3rkME9I3BcSJIZtCMeKrZs03JMG4VY
r76woVaVPjNIDrBjmzp0DArpkbxsK4GQvioe6eU0CAQIctskdNE4JhN6KH8exEwQ
VR8Vm39m5utEo9jN2wMgfyxkhN0oBSWy4TZ40TfQ53cXM06D6r627uQVkO5EGokn
zr1enaHC47fDoni1MDN/l6FMCxQXq2TBWosOfNwX2BYNuVh5IKmdpqbK/pocdO0L
WrxHi0pjzhqMvCHDQDBtmGxavMFqrQ4zBsWp1ZdkJE+NjQq623VvMjs6AsGnfURS
TX7QM8Yu1HFMsTzyc5uEThdpW5bj2ioLWvpCZSm4UVsVyU22OjHBmg3adGQNrLhL
OxZch4CKY7dq+heqSVVnRdNg+gbk0PFEQ4cviHrBEUFFLOoxdrHsAgX27UrVno4G
duXcawqT+eZOqXtdxqBZqT66U3bAr0uG7exOyOebnrlDv0JX+RSb0I9TQejtzEUc
9/GstkPrdJ0wJUkXEg7BkD9BX4hiIIUfHIT8IONaFezxeGUsOT1i38XifwB1J/0R
slhP0Wq/LS1S9WlRgYK78+EJCax4yZ/D3PlC8LxVPcXO5BV6NV4qGlj2tsRGSCsK
znOSiNH0C/Z51kazStSLXnwN9yUYsg24OHqjRCduQcTfHE+h+/a2E1sUmV9kcKng
2TxEqjGsipb4nMm1g7HzpzhVVDf+NivipMB3azFYwFJl/DrV18sQkLTaqm83SvQN
IiXm7im+S1t0khE46KyHWUR/Wt1BwNnp5BDEtNEbvi8LYyI//QqSUBkldymjRk0x
0E1u/ovbuxawoIK1Ty/ADkTj9reUqX72AntMBlWkbttjN2E1X75gWDgoY4TMNQ96
3ngF40K5r+PjfJCsaSXFCahYjlHl39VMjoPvFHXbRpIuzB2/Xac/K1wCnCgrhRLC
Z6FZ06TYSlNyy5JzsIEsHX/6PF7sIGNFRVQUodRaAsALeGciIOaVQ+A2ov8R5a9Z
/1dSoC7n66lnjL8FhcT1fP0nSmy40iGzqqmt0/4lKlX4x3ivsCP4dsi3zaLmBKk5
kRfx5c4uC/wyy8Eg5bU+mQR4/LSmbntSt3gIrNkGYMNKx2etMTgcVRbx3omLosNj
wG6aebZjyZdga1CuKHTx7bAVES2FQw8gPaRPUrxpfILXfcfluX5OHilZx3CQGEnF
v1xvRSh/walur8Ik2n7XIZ87i0BI+bjcLFzPnRZRMCbstSpkUQCz9oj5gSQdsiWL
JeoDsvgZX/7rukP5Z+BdcMkxjqB9EXw64LkVwpz5Y0cIqAHEBnKmPrzdO+A1pE2l
wKBIwEQ6vWjh+sxWh8fZSRTsSJAELWbyH9Z0aRcP7m/Fz5Z1UNLrkRQ0bXnOP7US
oLO3jSiw/Hr7SMb3OhPNljsFDO+PvOEuWMJljOIyonBRES1G8GyOy8hyQUTg5FXD
JhJKuMplRYuib64tYLJFsKcw4mLb8EXFb/gG4UigB0Edpgac77hRntSsLAbZZLcC
1VkfRCcUbIDcrYg+LpHrgIkgQhFRrVpfGhIJz0xLMG5/eTXzfz+QAmSLH7shK+iR
POExl2ns4Oi54EptSFe8AqEDnBZL9cFyXj26BVJx2ep3+19N4ONfdJWkRYUv0xKm
5KhAtAfo0ySsT7+2sJFTbhYxUGP3pGuAdqhbfh8KgLDN1MAdSfPhz3SLBhzk1CIy
hLJaGfHkhYzct3ERfAWPUxQKljfK8tPuyfw6pk9ZQoDYsOzrXDGH9IYXpJTQfF4M
guuHYV3o9HOHPNMx0Qa5bVFzjY1SxPag+z6LuGupabBa9ZdwMz5s+GDiZZG5LsYn
ZOoRXr/5dM9i8G5fHioJBlTDAs1ANDKFIKMBmlL0X7v0pDLNh74WboraVRU/JkpS
X1+qHZ12dEQtRJp+y5luKUEy7nd5wvxjhmGrZFxooE6HjrTE/wpu/a06nHZRfFrM
XuHGZhT1wEb4OMT/V+OrX25d5kAZyxfvPF7Vm5EwTax7Ng7TUODRq7vFqinQ1H6K
BJXrhR4v0ZZEEngsPVc0j76GXr7sNgvztEPRdQCxHRrkF/My8Y+eOGfB7UFvB11z
i4ucbqQwyXn+15aplwb4Pzb038s3LFG9r2+/AmPQuwl4Yowr7xcU0bY/ZVzOU0V9
IGZyOWIbAvWHA2fmMx57P5wt7tCj6UhftksC4e1a5j/RtMgaeS9sbanwNWrnK5Qx
sbg2pIJYOosJuMIuCA1FvDSkP8xHQyAPFHwqbzjn+TpVustHbUKDMsimmq9qcfDd
SyeweQAdSaNA48Uur8FikRNm3K8r5+RjKw1k4V1wQerjgIHMPhZJv8DjFfjJhrgO
ry2Vhyb5j8CpZoBtLo6v4tGm4Eqy5fPM37M79ScUrPPthAAX2LIG00CfkhgOUFAk
Suhe3tQ4LKP2hRx1lRulL5jzz47ABphbIjS5cYzmpyUXGs+/3Hk3Pi+BNdxk8L1b
k0vle8rSZAl7sO+qWtJZ/vGPuTlyVrbBLN+IpN2Rr2dg0ClM6JRd3nWS6Hot0t94
mjYSgQ6M7DZ1I2xpXuiV0G0/yvVInzq4BrzveSg5MBbHlSxiuORx2pOKmI6bVHe/
irwqD59XUFT5KJD3pOHg23s0A1FpwsNEo5Xd2r/vBkCgPu/DGzwE1XJWI3zbUVfb
6FAlMOacdd0EjDk7VYe7Sp60G1HxZAHSCI7Qbmgk5s/h9aMA2uANyLB2C32SFllj
G1hz6l0WwYRhxuTOjAx3vtetwzRuKelM23PHRzA64si/LB56xU73R6QGktVBWVTn
UAcxBrIId6m/2xbMBe3zcg3j9kgtL3gjdySiVnD8UFB17oHXw9m02hZ6kLRlJnIO
tbx0I8DNTpfdD2PooDyk3NmautPlIAD3xtyL10BS5FA8dErHfbehJV8pbsKsJjiQ
dcJXBjc77TbUN2AWzx1seXtXv1VAjebNh+1ImubiBfp/gzz6GraU+ZcLMgvjKNFr
Mqhpx27Rk5V/jRPFZV/jgziGWk6YRGWqe+AAEgYj/sRFq5dT9Erw+7VnIj4Bea2/
LxsoI/A4eF+62a8P73yJwgrByg8Q92Hgr21zk6QCbiXpYu6k2SKNBdzbYPgnzpPr
ZFpf+QFbmhnfdtMhDESZTxcL0IZB0Vv2D+oyRj9CVNveeXK1o2wp8mlGPr6OcQSN
KAgy2vPZOlAA2dS4FuwZc67GOr1SxkCYoZXG2TEeDY8ba1gvMOIuG1/v7lOYdM7s
F0BnD4ENwqZ6WeYG6uUNzR8fvkDRQqwCYKJ9EwNyRODDp/LSYYxgdw8VvBoFdbeT
dd1o/tgCFGBcDJJTvjRKd2LdHgXSPdPlSZqT7TOS1WObRDcFcb//Ikl90lTxAy9z
AcZHA8uf8suXu8x5E6qJxPUh7EK/nD/LDlCpFw2jKSv0OjmNLN7EAs3x5oZil5Qe
RFd/cFt1ppiRE9mECs7gBwZijcAsQWlipN838+W6SsWN5PLwESZExMWXYgw8C4MW
YRzsbD9q53V897yK+5jVfvvlPfEreGa1NaCUG4nxAAGdUq7EuirVHefoSyStLuIp
cyTR2IoJF4Z3W18Q2O/ofWQrlfl1fIKHj8ze5OeJ3QnSRxSZl++OQLicTAJsA6it
a5UjtMKbQBtpZMec1BethCtJ2a1NxFR+UPTQSYZOv3AKnj1ZOcTI7aS0j/PM7K0z
YT3fqLIop3prYuuS4hOOuBOsdTQY5K88QqFWD5x75somwXypIEJpNZqSaSouEdP8
ucOubO2BvqB97RpUOOTcX8l5A36oo7FFIgvqtSqZfhgUgH2vjixPPN/o/o111fYn
azTlClKrVOHLbdtaNgathXc1qTq82Zf1/9wYBjJR76+jqfjZk0G62zdTHK3inkwj
PmDU5lUHle5UKfmcsndEFZv0BSUBZJvbVRdnirHrTY40EzQo1+JgLFXIXeiUq7S+
wPkjuM83H8Hz+oC7EkBEyhCTGibDAroP8mKQVlT0V9OGrLV3JnGFiPKGSC9LEoHy
WXpir8HGG1VVxfGCK4juHByIabmBbihyEH8C7eunCITX64tVMpt+DuqJ9m42wRU9
qAJirAp7DLbpZatn7FwXXkm30cvkKmnH8/z2eRrwkjPCQqS0Is5Yet61ei+UE7rg
2f05fChMYntg5XZOi5WuexMGFYPTxIEeGtVADQ+EIRKPwedfghOgpj8mxXvHqBxe
ivyQDzrDq59ujTp66HeiE06mD8xmgjBmXUPC2UIv+WRvmqjjhCmularAdYGjsQHN
nO9XAO0icgl4xFswlu1uMcVVthGomP2fBFnmHySBXCo+ixVHYOLx+rUvM/GMpqdi
8XLNLp8zBt6jCEqIPN8+VQZImnuPWOiL3/t8pVpji7/UscfKEXWSECeU7CjjjIG5
EsLKU3Fuq8W6+f1ppTzj1nkvKacC6Ap/Be7fAeohaq13tcAYz/UtGwMMAs/wJfn/
3Z/Li5pdAjmwrb7OvT7Ag8OLs9ekxkgstzv75PLbpNB2A95jJvT/qtXRLcj7Yomu
9nvf9oouFYd4GlYERdfWKy0W6YarT+1Z6iD4lH2F0qIfwgJVMkyBErTcUL8HNI/J
MoVSItAn4Qv7KKuM1vecLp+S+clFT9Syt2HU9TVL+3hR7kX49GYrsC2GtJ/CqgOn
sta80qUhwqdMiT25gtWyjZ6qu7wXk1f3jcFFgxfjsD2F9l0XGO58K18sc0cx3HLo
b6NY1QSsNqemUT9y0hLUD6QBa6koYdZxP3sdkQLulYL20os+6cx8ortRIXgFBe6A
qi5FY3PmVccncZdi7uuex0r+IOCLOSKFA+keNurM9xrqJSF5l9BGmZ7L9/SKt52x
eNaFexg45HOJZlemIlXt9qRxYgnttgquv8NXnPeeAUwOi1v1E/JeaSs/3iJdIy21
rsERx+x4EuQaT9nYawCjz5H2bA/xbbPzp5rit2s0zNp08JmNnD9qpbTPXSqHKE65
R6NlwhiSVyrzjPQzWX1Nn4sbX7wSI5+0qDllIuuJ+r8Kyd/4gPJN8sgrnZXwpPSP
nBuPSKvLHLPVvTuyulS0OZKlf7MvNxN/6MMVZ4NuDI9dEaFuXVLDUFruvCiQd8kY
maQtbi/zK4ZpWUOLio5cegctE+cOaKEI/FMPpSpEKfUXBVJYifF/Q40T0U1NGPXS
ouDvXwOdwQSmlkW2Q923un6u6F8BEfMZGOo+f26iC7nl701QOCElBRssijdofEDQ
PNHbx3zb3sGPBv71u1kFXUSiZ80XpS1DPWWLSPeUv9V32A6RJwmWXEN9Gk+I5wdq
PJP0cGJE3V5HXhyvbXaERJ89BGo/xYddoKETzYrIOFOgaCVnhhjzaHmmgJ6JqJm2
Q8REID7GwO53S+lFFu931kG0GrU9fvZnRWd2B7MkTGlyCbQlm3JrW/jQtd4qipj6
oz1TNLoK69l2frBne2zo2eWCs21QzgMWvg2Lqx5pQo4OCGEr6KvMpXI0Bo6iqByN
YybOhXjOZAWfuHqO4cctu9UTsxxqQPV84xbNlvHx9TFiuJOcK/OXbtctq1MR4svZ
eQEqMLUgcgPoVQdqAngEuKZ/sA1X5eWmbIfnEIBIP2TZODiupfgpJnY3QrWlIGbB
UUC1iGDwAIzA6ug3hm7UpKmhaMR80p35AZPQCG/zA8Xt7OPHGyYcd00NkIW7XA7y
+Vm+gu3Qd6FAlQ+DZxu676oFgjaq4iJTu52lrN8SfuSGKU3ada1eVuyGH+a9n2pu
KiUnVDro/4zBUTxrbPJs3RoViwS+Hq790ZwgxJ09AmjW9xvvYx5QI3MxU8xyLJ55
TfA0JPLyxysSHEbPFqPo35MdkJDg2KNqUIsWp/xJg/7f6Y/ts67I5390Jg2zk5ea
7cB+3q8APqtIg6Z3mNhg1XyzfSQdsmyg/FkUDMq9I/PDSZdooTOhxqraOGMuS+sO
qKhKKTVO85+pNDBVExRjjOmMYng65UyMKfJe+8Dl03A/uVZ1gEcKuE9B08FOZ+rB
zFPuogAn+DLpoWdn5CcpiI9m6im0J+UKYWT13otjPwwnS3aDDtucss5PmH8L62Os
to6voUncU3GzseRaaQ2TqNtUPZo4TqWQosOqBwbxyeToA7wJTWn4/G5TWMrhpWud
nlNGFB2WBdHYPsDkx3dlfCXXbKeF5IfoqY+qEedvuGtplpylXKrINIG1rXTZazGc
zSdt+jsNuABNOxYmFbSYwQ9MdVZTfVJM9FNKk1cA7qrbpNv9Xisg3ka/gk+wl6Ah
QTKbgNK8JXvapAUEaLgJ2fdLSR7j3+WSG3+CbOphxrkHidNGFrSqRXJIWTmGxWPr
03JPRscKfsPQ8ArYxqO+Ma6dPmP8XlBJl1RW8HpxVjMzxkS5f+/8LoxcMGOOlsL8
3PVqIUMhx38F5yZqrUrn5YVcTtSsc9WYbHykcY3FgKl8wAAUKPe7LlskJAQoTMST
LQQd4eYbnf0etCWNKRAdtFixzK8AZ3i4vK1oJF2WF9FagavqJFabIZjdpR39AcUi
bpqA60vDrm7k24AOsreK4bvQs0zMvLhrMqbnTg24lOofdJDoLEdh3vouriM0Kauv
jhVXDkWzQiAYhJCj97DBckNGNd0/oowcUCIV95eEyXY5JqhLF7+52fvQXEtxc7hr
LBNFEfkyo/EIn3JYpQl5S73TlGt55OjAtF/sN0fy4kkWSkjWoQL0wWA/I/7Px6C1
JNKHOUWpJ4/65YtdklbXrGf78mYocHG3rmUOcbyDUW9rbFou1YmBeJBD0qOruX4q
zZKrfqAxh0tjspB9XkwTiclH8M128w80Myq79ThYOXv+hXzpZkzFLmv4UNoY5rbw
OZgW/MPcEAcQg4eIQAtL3A9LMlR36/QbV0zm37wf34mU28ejFXKyByWWqKuxuPz5
3gt6C3CWRtoGrX5PkEdLfdlb/zI0bMS/qulCMOwfHBVQYTq3vF2pcj5NDZn2O2vy
zPK0VLN4nJP7RnNuKpU6AyQ3v45IVSjE8yavf+VMaptXc2Qx+oXX3ejNmzOWvVaB
p4wIjYxebfu2O+c6Sl2cEgIDZicWPY0SadgxY+E3b/3/Rf1SBOvu1Q1cbXAWolLS
jIPYravbPQUvo5Y5zdiSExWBxhbKUD+ZFEWiely2pO/wGmOe/XnDrizlr9/85cSr
OMIIMt8NvuaxhZ+OoRP+UuW7tEj1oN3oROi3y1Uw3kMqxcYFbcaO0NISQMvedxeM
4oPS03yPWsW2v6a1fzAzfpmlZnC8vawO3smjFOGVNaO2R+LVcHyBZXuzjl1FDJHd
eyAzrsPEmiGMkxZCfSVHbYbyVUYZwpAyt8jMzidSDCQrDHvEKArexjRESGxw9qdS
pT7WFZZsL5TsK7w6m+3RCW0N/90nIAGW6+HSBPyjLiafA+f3GZarGjYgErUbh2d/
P5sdGCPzBRByUodIdmN6HavdwRWppchWXuVjYhQsDJNh2VQbwxGEoLMHDpDyVmje
KoBOB0dvZAXny2pnAECYcgOIElhNSdP3ZgvcCh9t2a1iEzgJIr9U2zQi8x4Av+/W
L5VITr65tV+MtiJfyWvBXoP0A7+hgHihr6w0ppMviPHshG88N80hwInvIioFOVpk
0J3o/5XNQppDJNGorFjzTaTulnZijn3xSwzprcEp3AVGIKjiQLsNWc1FYqzCx6k3
q2wdI+JVViwzx4+n3CuSkuStQLKaufc/QGZD7kO3g/HrN8Kj1gvjuZxbn/expbdg
nQN1SdnAKNC2OzHQeYtkwotZOoz2iODtw40Em+f3YrMUgD2aWnEMJCIL1HhUlW8J
+joKqs6x972xpdlDcCVaumaTqQtNe3sJ1MbEOKW81gtnANepw8cSTAXDSxeI5+Sd
vjDqM1wKrEoRyyyJgT6y7fRjR87ZV14EFHeIFN/chVyL5akPNBwQsY1LiHCx3YCo
XjPqSZRoj09xIIzzOrhBYTY1pp3DoEwLaQyAd2lsq5DdG/JPBrUqGq5Ggy1x9qrO
LubnOVXfgoqv4Be18XMxzJuaFBCivGx5eUAJMHL9sb/tIHPDYGFQ9jwaW4O8giX2
nV8vaXdQDA7prfyc1idHTPnfDK/qnPDjT+81lrgTcLAEOSKYHW6ufSI/6Z1Ch01U
7ldGm3lWH7mBAbfrl+Pe291BPrTCvNpfrSwwaVkTeArhscH7ROwdslrMMdr5x8nc
pUzMTvL7p43SJ8FdD/tWPKShSL/v3wzn/twiCc1Yzkb27DW2jSIsenbdny1GSpGX
Jq2MSE1cL6xm3e9X/sjiLygw3e44QMJNnz+Suv8VlHDEn1kS2qxfuEFcuyDbddzz
vYcFxIk4U6Cx5oQ0E0fYkCGB4AZbyUVYheZXycy6O+ycK8HyvdPN4pcOwNQwVMw8
N0uAF2c3hNGc2Gq8SQGlHWG5dkZslK1xUPxEy9BXEP8nThoPD4cbxdr0L/AGlI+U
eAiVmHlumJWJ41qsn/KOH6M3d4QU+ktphrwRYQyGYYXAgQ05qmLWxblQeq5VJhPl
3z4EQLG2zfajn8LfmGDRSzou/i0Xmsu7FDQiruBB9p5eH0UL/Byd3BYJxDOXEFji
Sy9djKF3m1RKujtg9a3O/0WO/z4cbVaMamU+auXhZjESQlsTmSpx2TaoiJ4Y3tVc
kCt+Diajcky4UTc+mzIpyrcru9wwn+y76zO/v/MeFReWicFXlzaMOkth43R6A5TK
Ci02EuT/JRAJQbTFLTpbtnCrqH7ZxQk9En18PhQTU0cpOhuQExrFG53RHpkuGjmy
e/+/ft5ifCxHXwUpZsmDXCLvzI5FU9JqAtFIsdJgr9ph3IGAu58mqPe0iPby454o
AXN5NSU5Xl4xu/rjhodmGeb5QBZixD4TaWEYFPFZkSRMnwE5f8HHPWX+AaA2ZWVw
2HtP/mHKyIOBfepzMrvINJlxCGVw1KkxDoHI9lU+5tIe/S6yyfGT4UsqUr4353SE
lWOMR73T9xm2G52EVwHvpjE1BBd3K/fpiy0S+uwzVhZHvLHGtdDyiGj6xmwMPzLe
ZCEFQlMY+sUNYdeHNCNeO7gq0HZ4tyZP/B8WE2cyiVQ0CXzXEqgDb4tmWCj71CKQ
JrHh9SBWoXGiicpwIDkPRWtYURTJlZaF5cDI1pBSs8h6d3E9L198+nxqEWAgEYS3
62h+xdrB3M+6c4YVwklF5dvpwWdoWqHLi0RA/wv30veQmuRlhesTEA2Xsr8N0/rY
AXU1ocVtjFaxMGpIB0C25dC3VqYsry/LGKvLBjDlOaOktN+46JjAVgIpbz/syMfQ
jnCVeILa7+y4X8lj35t628a3ANzAhmCICay281LNQUus5n20kVVLP3M+L6bJP3X1
ee8p7y4BqeuVx9TZgS8YkyYxmIOQMe6mCtCCioEgYkvK8eA3koyukRzhK3flRQqi
ITdWpkzZrSuArL0rg6YMRoFj+gqVPwiquJY1EYHkgTjn8WmI1A3q+5pRT9U3jF1K
AnixweuXMAOlXyrKooNmz9xungInHT0d6HIFyWsiziqrBPD08gdaw71OLlWeiYju
ASLiy12nuPcq3wzW93iJTuvfSgH9AKMpepjgd2DMQg11lOwMDnScMwU5K67i9tip
3C6tVNyu5pCDU2w7o5v2X3w0bcJ9HIuI0+A3+YMAZ4UJaDPLFdil6x7uCV1/rVKp
hPgxtaU/BLe0bEsRUCR0EkwlSzdz80Xu71opmrViSsklTn6mZz/NRRxT2AXiECqg
45eqO5StQge3ho2NbuNgXegmM5Lc/az7jczutcIlCIK98m1+/csdJRIf2AfAp+dL
ytl/LVXBdCV8ATjGXAWBDe0F1JF28bCpWYbdBxmOAqHBiKx+/s2XZqM+2uqA6eGV
NQ9EPrO/giE+66JMUeOCpVCsBMteTpB4HjihDICDsWLK2nFuD2Qb9AHdN4S5FgZQ
wBn6QVA8PbXo3CYCIK80A1cg+eMATYrIdqQs+MC/NS0pehtJySm2x7LG/AhlFAIq
NqpsS4f0vtTWHLHIL9IEbBBKg+KjnKK6ZJ/ca3rfHh66pdco6J4nJ3lbJ9CjlXP8
rpyJWgCXsp8u+dCg14xsqloy7lizkueNyksCIaRfFoLQYdp5Atg8hL4v7k2JjqfN
xypUKGy9YAW/soTkzhjLWFHh9rfoYHqIziMvTp4tPsK9A8BgS561ZIY8Wrnmg/DY
diP0CYzQR3zt+464kdRg+h0hANpIpmEl/mSs84njFIzANMpshV3KirCHk1ZkCCyX
Fi/6bjI293dHfG+/apwEPe4CWRcdOZOstDEmq3jRlPaAugmaooBddQSPKhnTAGxD
ym1r8E1e1drkus+lsheVOxF/UblRCSD2L8dr6aQ8YD3M+YLuU4T1S9Gd2edEvCNr
mDPfBSICn3k/OP376vN+XuhUt4uD0xKb/fyZ0CnfmA7mjrUgZfdEThxPwrd3MqGI
TCP3pXeWfACUJ1YshMP8GjBrNesgwOOYtEhCTEky9AcWw3q/q6licvUFYxNeAf0b
5sk20HhRWkUJ5GQs7Ilvua/KJBunTYiGzeLMmP+ESZsxst8FvO1PghISeb/xgDSC
JR8X30ZCON6M+NnL4ZHXkyz+H+EUIsY9fXEBvh2FZ8Oeoq4s6rTzRwdA0IKCJoav
zuokNC4Ioz/s76zZEGWV6v0U3OL4Gz9yjYL7gtP7gpnP0smpLzyOMWL46QPAfkto
TnmTA3+8INhJlkkZFQ1Pfs+Qu/+PlieR4qNz1SNw2bDeRYXtaIu8ILyUQytBGPMZ
AfZKe7AFRZzhwJu32fBblEy0uxs+CKvIcTAMLCPXsIKOuYdVrG+99Epi2UhBJyhx
64k2UmfCNKjyiHC9DpHa7hlUUhaGLqkHyHZOKxW8Xc3S14QFRfqz0tdpCqnfM8q/
SIsTZzgqkZDdVm9PGYxYTBl8YAmFUyxpW03wlsoYKX1IPVyDnzbaBMo52y9GYhkU
Us4uL196ASWVBPr+QYrcOZgRJ0CVRIO34kfYo22dPFXmmWj6jXQ3y59WwaG5/+7v
Tg3qUh/9PiV7oMlKLzqfz0+9+cEifIssj4+p0l485m1D6NSUHKiZbfGZ4NbXRNha
Y7eVEwU+nAjWZU2PrUlEntMvpW6r2x0IHFF5bGFk9lh33XHhL3nynALBGlLAuX2X
MGjz2Y3GiVfHJg+4j/cHnAUKujmXp0T16nHVOpqOo8DtPYeN4bC5R74Bu9aC1TDC
yYi7Cm0Vz29ARUCy740jogkSyNpfZ1P4HQ3yF7APY7/+PoTzzkMZAcSBAAdnAoPe
Gc8Z1tYX1cq4795nCbUCjRyVGzyvb1aqz+xxR4y6HiyJO6zmFrE5VOPHymk/5j29
Okz0fsIolKhD1/7u6V/MsrD1L1Oi3cBsiTEKcp1OZzDQjG/EMk2j8sC+N5K7FbPP
wLbmSkeCllkA9EI58p2Zn15N6WKPWVbwGEevGWqkqLzUYrkbYpSb7gaiGeo64Szx
Pgy+B6oIdhAaljursS7Cfn0QV1zh8QWsBB8xz3oibocmMi9EG2NQPNsqxSJbmrjL
plY381oQnOrrw3rklPu2XJeyIy18NAzH/U0gw4FL5fS43+2DA08wYWKYeESWoOGO
QzLs8KTfmwZtT/NeDHWvE3AgVRX8i2h5iPhc/YhcgFa4D/gZp3J2yGtdyQXBTfXL
8LfpPKiZB6Dayk8Sk89nA6hdn2f0uibl3Lgu93A5H/mA6O5D6Nh+AZn+S7C753ZA
RuVWY5W0S7EqQmgpe7dlTx1vtpJ/toF6fM+B7Dr7nDfdreXiJMUans1Yxq7Ixzgd
I3PR8Cf3lS3ImiARIT3pUWWMjfYA68kam+3YjEJb34e9zMbpqrXMOSRU9EqzEN/6
AGticBr91gzb0/6fjVAW8ZvlkzAKNyoRoV2OGceLdWEaYNef8I0T9vx4/nUjQmcC
Pwk2FRtGz/SYHt6nm3Eyd1LVyF/sp4xo2So6Hksg3iV104f0fS4ZVIzbsTdYFyZw
8cU7dy2tC75wkZQVxQRruM/8jP3sjM1YhqOCg5G5l6tFfZVgITki8eWCrtxyJn+R
UQfvg+hTe5BgMsowW4upxYfkCV9rvFWQ2941S8mw3FGZzdUIu73hJ+HpSeIxnH81
VUztpZ6xIrew7gu2IQ88TrgKQ1WwFRtQ4uqGse2QUh5CIZB614gwStGpE1XIivvO
FHG2xJ5WbI9oYnSgoZohT6fSoLrAsIET5vFIHeYfiuoWLQuXEuajMbVA/roEZAIh
EAAklMcq+OovNILYcVnovgFUUFqKlIokZ5MfL+fkUK/UlRV8l/BaxUfbvA6zvn6x
mI90c2CjoB7kGMw31+HqxthRSYI+xcGaR8fFJCPT9TpZFAN56zszymibvIJgzJDM
+vDOHaVLkPR67WHWH6ekI21t6EU6wNTYgOwjdgP8kV5UVj0LSjpC/LyzwW/FebFk
EIyn7SQQqicql3lDkjI1Ujd6nTUu4geDiWFR5wK2Dbk9YWtd0Q0UNZxBie9dnsbV
mPkpBAAC35r9k2hSoPkj3DnI6qUAul9a+QPyOUk2UKwhfp+iz9cikF933XqWq1aW
IW7LPaoBaVWxRq/Jhhnu9A60NYFOykdYLZKn5lICCtYNxbq3QZ1kz251UDZyQy2m
A1xf2L/Ze9C+zZ+MeuV8E86rmUjs2EELzgIsu3PVeruG1QepzwCdDwMR6bkx3d/C
QYOFbRRLaoh1ICFeDV3wvLSDTI45A9HdLpkDq3VEErSDKBa5ttevmcsnMxHA9dQT
oXOCdaHZaF8QQimX5vEBn5eYJfnp8Vg4Sl4qvDRBORK82vV02zxD0TLTNpjh3sx5
N3XXBWXK6Gzq1Ko7uTnWzFpXiUvGAfadLSXvzcmzF//RV4Yb+Gdg7xOYYHxmjg6l
quw5kVf6EW5ezqXFoV28F6VcGOfc1X7on0Cq7ZWWQFOSYuv7rg0N9O63dFAh/tMs
7NCd4YcqOIDtP/hR5M+HKdSq319/76kNXOGdaLslf6TmZARH3O+xnJ5YloAtXiaL
ygC1H0bFcu1pJwTGCCJ5rs2Fr6VWgeUY5qG2GPYJm7d16cDLRtH+0GfBY6UJLz5G
ryp6GAS/QSM2q3GMZsLT+VsVebUtEAomFzqpP1w/3uJDbkPeWHiz6BqYRPmanxUo
3Fq6UgRpoz6++Ny4oF6BharotIST6oFIUXODe49k+NN79kuIJvxYTO3km81+Ox7R
GH7zOmP1sMxWTrmO3sOymKlT6/ZdJxpKHvKl12r63fbWO2XcLkNmDQXA7ajb5zNM
FBmxyiG4Ve7vER6dGUX24+Z7RF5+aItDlNDc1nuot8ZnTEJK61wFCYHRmkTwoU3l
NKsROw8eGBretbe24SmrpC9YluwnGgiNM3J0qQdMZXmVMFk4NIcFTcvZorpntum0
43YqjdB/kPI9smNks8xPmAtTChKEbDIMZ0FVdqz7XwhIZ+67zbVI6afgrKPmjHeF
ZOwX2QpzcpATz6aRCTIcCe7/dMB5SSR6UpWyQ52VbRL7zk0F3rURky6Td1c92DQ7
rY7C+pe7hSuX9BU9P40OI0Tucd9QB0SGdLPy6/XHC+toktF4mkADDS4uXk9aWTcq
aFzMFdz4uVjiLvwEoxfv2EU4Zvs+pZGlFot3w979edH+Peuo73T26yj+Xh/cIzeg
/WheKr72DD6pw/4zMVAvMNmng/myuRlHF/nJKDeOlvAZcdLsX/fmPWWU+i2r1dJk
MjRdX7fgORhLdAEC9K3d37vdyEobTS0ovQWq5QvWIzIVYb0JvKaQeg4awjvHu8xw
mQ3fJsCzzHLgA1KgyebnC0VYfgc58syPGrVt1rBw85KSA9bzF2AXlTDMLfcq+bCa
f1T6p2eT7CqV+/Mij7kjJWD7ao7ImkFi1Rz3ZjtKFrNcl6ndFEvLNNIuu7N33VZX
+BSEMISLNUC8zlViQ6cXqI8VDTWcJzxzobGMW79wcqJ1CnIf0uPM9jrGeq78NPVt
Cl/uEtr4MksGGyloift4PtjEMu3lBuF76n8yO6tyWeyer0p/WsZEG3yy4Y5DDDGC
6HyxVuFcPAYvL+ycHmzF3mKaCH2TlK55wo4iQWvo1dyUd94mQAkBndqxdJdkjKyY
QvT9RgLwY2HviGpJxcv8tTipAgs0RdejIuz2jgSpnEYULyT5M+10W4k2ZU/7+RdU
/fY87dFeO4E+EaZhFZNZABJ2l/CJYND2BgMUOD29eXj5KGG385ekj0oo42ClE0CX
zZ53cACQYQF5++6OpduInLMf9OsxGEOrL5JBcYmHyI2Gncam3KDGnP2jcJgE0gTC
cXmIS2QfWfkW1LbG1zL2e5uuvmAHrefx/7QZhizfFu1Ir/ZIglMwvbkTroTaDhYm
LATt2VXmqL0FEB8ii2iLTmFlK86ZBi8sQTlzO9niKZY0k3Gj1babA8mWcRqPwij1
TxZmcOu3/vVFU3PfxTTw28BQbf3Ber5uuvZhFmBRBju2sUPBMjPnWUVbyM82FSA5
vIeXkRO2CABh3rPnD1bw1fNW097H7fpTS7O/xEqwXIf1BDBI3/lyFvE8UxJkg1qV
/rP21taab+JRHimF+UlgBomPbWV2TVOH+3evcqY2YifsDW1oIovXOQ/JM0KGCxsa
dAKgSa72orpoFr4jjH2Aikh4DC03Z8Nzm/zr/vMBRnnQUmRFVedw+uqqNCpGeP6Z
pxL9bemzwQA3Yd4iqYVgJpWtDSk/R/R9wTPD/2T1iEb4WYFavEU2T2rMBtjNb6xp
NYUOELr+rfSQkyDcfnPUwqXHzUpTfTCj7ECEwVo3HbsyVH+Gv04A19eygPu9CVH7
0v3DKdSwIg/YKeVDVew7AA0xfQcuGXzH7hYrBl9ExPSDtvc341VRqxaEZeZXqL/R
SXCBgDZSS34YDEebORB/eYOz656oMe2zlzLpnFQVny1eTtFzGlkX7YLnrK1hPOBU
mIVR/snUNJILxDDuqWSdVW0SKHIF0AfBH/YHFLmrXj/HkVDiH36hRpqLpAG0oYGf
jkrfQLHthTyXpNgRinVaRJs3BMUAlEBI+9NXVb1NXAq45h0jpascRZ4MMHJxATkF
cLCGDShFhZqt9Ge1HRneZlxGOqM975+/BF2NkupA7HJKP3mmeBQcAETo4I/jsuQD
NGTls+9V+sRGjcKj/r1zYBSubOY2wBZW6PLJM1CDpyVGu0azg8WyAVA7FA/fJfcH
xO1GeTjuynhADhRQscMOuwLFwOTYzZbYBnYRY8jUZcZsxEaaUF6HEv9dayjHUE0i
QN1HX00c3oAnJOsuSC7romB+sSsy60Ya5pbecVP76996fHgtXQ5+m5bclu4ySapq
CxxIJmMzbjm/ZDZKqG+hiBlMbR9iD5NJfsHdzDj/AiK0jlyD3+zMTkLBeZsWREaY
pTpRXG2UQbFJlrW3r/31KH5fkFeuWA9zx5B6UE4gBqavSML3rb3UBW7QUEz5q6kY
ogOna4zdHZJUxxjTcfXTU9QqDa2R7JtjZqT5n3EKonTRWGDYXI2n9MsCDiRDnSLE
Trrs0DWaKAQblAGjLuIsE/iluMBarobIksUVy1CVTKHqBkQBRJbdIBJlmscbmud6
aLGK7erD0iY77ZEXL1FqZCi+6gy7WuDq3SjjqGLuGsofPF3RAar17/ci9D4Mn6yQ
RGeR3X0Hzj308BtfPPCvNMzoAkpk5dTh5U4x0wBJPy2DYgB3Xzplf3G+gqxkh+sO
JxnL4vqw89sDp+PbXPKzpxC0Tp4EenSx5E9CKMBXUMkc+4iVPFnF42AYG/m2JTJG
/JppgLJv8zXXqFtceiGhgJNu6JJucM5z/sfWWKoebMDgbkz9inJZOOolLG709ICh
YYU45sT/08b4BJPj0D9IdJY64QJRhZu1PLdRXwPNekeib4xxEXArXEdcK1HCzvaA
U8x6Zik0NhXLDfT5SJ8OzdXsYgEKFKY0ROZo1UT+oGVmhO2PkICoFwzGRfSwQhVO
wzaJfCyD4WdY/bNUTp4xaKWAjrINkUDHOX6QNSj+X18J7NnOjV0wNExrACerdl6P
6NJsO89c54KgkDSNno6a+Iit/0rqJKCOpzi2gduUdOgxgNltCBAwQz/w0zSeHwR7
gZoLP7gxGjg4QCdf5CdMlbRekUxKUTa5epcdrYsQtG7Gs7v0I43rjEOeCz6kOaSq
prjBxIfaAT589IjE3A+FJNmsZmry4dKbkla+DG5uJVKMlScSbRFvrXkeukdLKR1F
yv+dROU6a2+TAjO0uqmesIHj8k08B7EsV5BsVzhwbxEJkhz69P8Z29By+Y9EFvsO
bgDu6JuzsZ9oArqqoP7w6B2/jonMFkBcqppZ1KV46dkrHbK2O9ipyC7QoVI6ua/P
B/zr4NJFn9uLWkQMmcmV104x0gXmuZsQmTgVvfnfLOJ62Z5GNZY9OQZHimZpl6eb
36aRf5UOXjd5Wqy8gY6TwwCBHpCCW+kYsQRwAOGvyXcNj/Ep/SUDXtxvIlHJyYZo
Df2Glmi/f/EtLVkeGkuTknCuqriezEhLyUgvTqJvIzBM3/G/YK1IPJMVKGn23IXa
9HymH/ZNonsEow13tBhktzv1cwFsgerxcs5ZBbALLAnr1QFieiChRUsQT9A2aP9J
EQiYoDLy1cMCX/kiskpmqHm0Ny3Fr76t4wMp8/rd22NN3XV2AwcAAOVu4LcsjkWf
B+qqGExZI9bndyYgjXxN5z2l3Q6M34qjpNMRGR+AmggK4ivVudHMYwy34RZSIKhg
zK2U8N2JnbpyQjjU8/e8hj6itf1V6nqXOwb77pvLS3I6m7cwlTu6diQV8ClccBbI
rylsFm1gdcLHiadkRZlb4AqC0IkEpsPukHS77vAwHKAUaomc8nEQUk5Hgx/8ic1M
JjuLyek8wYSx4D5GjbyfQ9QSaDVLxP3w8gpSr5dpy5bU7fLO0tk4L+jtYRmRycW9
tdslDIwO7lUascARm6Uagg==
`protect end_protected