`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
YATj3kULTF7Ty4ORuRfFpnT6YIk4rUPRrM74bVTnc4GjdV8oSnW5PtQkMCLOi558
1V+/wvDfc3y0Z8//ksX8sZm3JZWtrxUppw8c14g9Y7owiwp+JumRtO1zuk5xFbe3
0MMnIxxoTKLhyRJtAxElG8sbx8N21OWDGiOk0Xyd5CqAmk9dcOIbxzMjW/wndBXi
maijUdqS+5KiRCM9+Gsp6k/iEAa2LnYTt4WtjkmDD1P5jZKsiMgFck8WOqLymplZ
ml3TTfn1UlLNm/+zD3SFGP0kABAiUT8NK2xBPQ5UzQ6sMFPd/np8iUZ5u4QLTWOZ
hTrU9OSX7lOvRUo8pJ9vPg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="BzW6NOo8eyBw+CxsNNo4wIDxODIsVe0ft0K5tGuSUZw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
DhjJh9S2BY18dG77XPz3hsiSQ73+w0XqfJhD+f+lIDHHVjOB7CfC8ieNRTexgzn1
5W+qoqOEwenoVQtit9u3XViXJSRJ0wfUC5a9axblRNyD2mUbyfH9+f59nWqGkVOh
ieHxkA/DPprM70F3APxk51m7/gNSLICSvbONgLGndWc=
`protect rights_digest_method = "sha256"
`protect end_toolblock="L7NTNW/5Dqy+2kJZXKczEa3js87UJ8H00YWI+92sDHA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 50560 )
`protect data_block
6eHODtGLmq6ccbB074dgNWpdzW45i5jL0Nzx5wwM+RA0eeOHXxEV143NNyQGmZjT
bzHAi/6AyRCB4X9z0c4MjyrZE8GF4crbMH4T59xFHqVrQ4zXCea5w0kG5yvHgpKo
qe8DCPhYAB9sqzbPdPbHVlBUQa7ieAM2NCJqVHFP6IMMqfdVejrwYz5Bx+C72YkO
jz6KrkyV1w3soWk0L7aPWjoKpBHDaEPB7jD2MMexYYm1O8K6rFsdEfRBFZvfQW+s
NsCSRbmyPSY31Qw5kArajm4B4ZYkvKoQbi1AdAwMN8UgZeBUHpB8ApazPN6cdpbr
t/pXqUIuM7BRPZl0RlZUmm5lFUYZi/iOjF8S0mUJ2rhKJdAkSdp11PGs9FrqLpq5
dyBgbqY9sSwkPNhRFPqQisI0mmwEDA5fFNZAD5sXasyhxYg2Cw4Ab5W94k2rF3hM
YHgkmH3asdmx95u1Npye4csuRb7ulu0AmQLY3Qp2w1g2JQF8gTNhTZGcjrwfSnR/
Reh2DW9DVku8m/JSLjkhP383HW8qMKctHkW+klMfP20kVw4t28+MZYZXYBaAR0Y3
agZc8Ej4kQU51jOa9Xqd7Uo5Z9LGuaSxDdAyTu+aN3tcwRLaCxZLTJKn4x9Ap7td
pUoqcf/ec19wfg1iEiUaRPd6QBOZZxloMXqX06gv0HL8tDytSKbUxQtnWM8PhYFA
RjFC96B6Ol/uJMDEmnRvV99GspVHYRwT4pgYFlBY9Q/VOJq0XVjbNtH0tMN/9dMO
LFAxDDqawRIMJlQHP+ey8CksO4tKvJ4/I+HNtRbk9yINOKHBCh95kbKkN5oaBYzj
5T/xB3ulqRaCLhJXkU7Lt+Y6WaXsdBPIdhDDz+/7efsC84jb4qSoHU/nEnVJlCsn
FXylLIfKbXj+AnDVvxpu89AC/CXmPlfKVIW9zMK9arkMQVytH4jVPT6DgQo778AI
Wv2aJuZ/ugBeonB0vOKOcS5lwzypGV1j6dPk1koXgCboHqawRztzxv8ubrE3rKPW
2s5SumqU+2lzr7KqzDzHJ0lyhXu/NwR7nQxAI8LvPeGOcEnqrx8G2etQv+LvGQyF
bRFwbMLTgRfXqdy7N1j7h9tNgPXSfwkdU4J3msgAE42bpMLtN3VGZ0f/a9X/quvj
AhXmADDJ696WPvnohZDdWGuRPzqx/iv9fCk2J7bDJyZAqqjaQrCr7q7fvMizCi9a
6X2htna4rxKcRt5C5wxfTtwXWBnnrCv35BvdfyW4KFLqxHkOh05k0WM7FtbCmUmR
IOJOJR9UkCB98E0+7ZMhB+XgbWYP013j7iSCEMarRJt2S1zntRc53uwUoN/8bSyh
UinjGI3iN/q32KtvVk/UklWXhimYGrXO8mHAvmzg2c7RsqS0sj6KcO4X0Bgc/i9B
QySR1Fb6FETTkLOjOHfc02TVvq+JlySwov+LWZazsPph1Oh9peI0MoBuwaU6YD2J
IFXqhmd8Ba6LrvpYWJOtOL/kscmo07vAKX8iYeVNs/03Y2UW0FtVr5M3kp1dj5K2
I/J/rPGh9oHQ1G+WdPRJ7hMIqbZ5e1j5CSdiPgyAQ0EsT/nOm98BrQy7fGy771aa
IbYMmin0abBYxOezPmUgqJGR6eUyDocmirFnoHn5hUV1jteJzi4TS5xJwJCbpk7b
YWZEyU43g6SbPS2Q06mYrwhdPnjjMxFXH3iuGpAJsL9Ub9zqSurGd4d0EPzmcvsf
iiR3OvTKhfmjekpf6GZQiCosduBgKZ9yxcDd66QY88EkdktNwOTAYwtv411UYEej
cXJ5XgCStjGxfGefvjYED8nz/edC1i0v0L0r8TcN0Y2Xl5+nmWnwUT5fO/N6laPR
6lmRVf4udW30Sl7QN7ZiCdrNDOLKr/dzuyjG07g+khwtmzKMW3WxKaxNqzKEfXVU
KjZtL8iG12DV7On1IgcEp8eKTADMc9TdltdfSlpn6hk5JKUfy+T96xyhBx7Ut7S1
jO0Ge2uDd6d07oMW+7YZKdLaBwFrIjcEa/yCiL50N78dlT7o1kX9/hdlsf96do/2
BTOlJJ4czsV5eXQir2uJUQS8FtpwruSsJOsNic4dn5EnvBcdXVomfZbTIx0qddrM
ceNv0XfikrPZ801qFOdXF/FwunPHxaiRQThtCEvscG4+u1YKXHQqbGuy68u89UMF
DxiZZW8nXWJwv6zcEtvl6tNK7MKksI85RUfVw5VwKrHi5k88NSNB/dGXr9axf52y
k9+XzKM1P/308cAYI7fBQHq5m2G4LYoXmAV/B+UJhZXHVgODKpnrK8LBhd6Jya9E
7lsn5Y/9SVeg/TiQ1GiQZWsE2Sl2iLtcgc/FtEy8l1TVpDQngQi3csLBlp166/FN
hD9ThCGVnPEHHJE6EpGQ55kwuYEasO0o7qKTsgP73iQdhCKaaJntyKgw1wDJqyKV
iWU4n3LClJ6EnyYfUDwKUOGHGlTTcp/b2QLHqXhCXl5lbVUdcO9n/m7J5pKoSHZp
W4dnJnmH0wPJqDfgVLq1Ik16iH+8mYK1qQwX9tZv+9y4CCpDbALnVdDCgbzQ1x1s
YgP8Y8Xu3EkxuK5O/0iZHDNQT2Exc9w4J8kizHwoTtOE4Dkia1701aFFKEdKrcRU
z51Qvi2GMDyXzY47EhgrKI0HtxYyhSWW7Y5nGZretk6jsdcce6HHRtnmtPCN9PxK
V/GIIu34pKAIMPiDpluogeEIze9w1Yu5pDGFHBaOBEbEykN/bd+qLZEwNO/cFcXR
gQsrryo1KIJelF0wGiIyLjYDt2bhcOnIlCIqJ/HyhT9TwCfM5eS3pU/l3R3c+3Nn
bHAGxHLvBwcE2VvgpdVp7kOGMbS/coH1u+f5u3OFp//pLoAJ8NRo3eaHPa0KWJJV
sWYVcKw+uRlvu8+xYpDXrjwxX8MDauM8llynTUCDvdJd/09tL3zs+W/tEMqeYVbX
sIwuSy/BkdtXbSNX00gFq7cGoSn31/aEeltdOcPQS/w8csBG+9C6ODqH/nE6e0qR
dx3fzSup9KHQP8WufgfRX9XA2AJGKW18CEwZRrI63nTc+eErw993UBwWaNgtnoLw
e+RNBCkt2EIuovguMxPTFe5kq2jw7yJ99FUbn9J4veJCgySJYcOMP7lqHnH4mzFE
A0KWOL4U8emh4flbNiNYto0XBzPolbQ1H7KKJmA7RhHeDRr8scKhfvAnnScVW8I8
XE9lTtBDVFhHXpaTMSGjQfY6eSBWngRMU223uXxKG61gUgxfokiCAzG6cD6YNxLI
Qiw4udvhiGtbXdV+74oMy86mF666+g6ueyl/mDx6hr9e0pULpSJkFgycJhuEWXet
SbIaYrDqJcuEnmyR/XmqgfzR7XimMORjYOeRuknP8KQssXBSYtTg5CO6c2Z1ZWTv
i/bCmZZ92w9+LpGMcr3SDiPKTNfsagL8AdbiWM0KuWBOGLe1KMbYty4qu9lurUd6
HWZnWQaBIFznSXjEYzIfgedFL6F1BootUFrsvMs4WfTeYZyCClf0mE5jzOe6NV1e
JPLvy/zdLdrLQEYZoZvInO4s0mPsNd3WY+o4Fj8oV/fxChWKpOBCq7/wBrwGgUYY
G3eKVWeJaDjpor0uS4M5QDYFc6gdUHTHFWQDjDU+23xCfR6GnPxQykFCmjI8JGC6
vbDPWu8aBLKPUju5frkewueQXiXGBIHPT69Q1Dy6EC/TNJmr+Hsoc2jE9J8x60Ax
UIZ9RQQd70TkZeqgkot7dX+C4KpCO9J4tbvoj42mmjKSj/Ew9FSPQHixYltMS6Eq
o3wYfXDp4maAEZpgbzWw0KR186on3xsOrRR49Y6YnfxEETk/sUMP90DnzD2j+nnE
F1YXMmb2telB7M4jU9FrLId8H5FfMbRp9QAXoyhLQaJhuCxZWubrIwADnnan3uAH
azB1sv/68JNnVgaRo0Ef5AV81O3VnqhgPSe12V26TB3FGjjPe5ft++9WLxwV44PP
hVuIQjlxQ4FyrVi6Iwrhgibqk8Krp61ib+T3BlgOKPpvcGGO6/1ASjgXgPez4RCK
m+bcVmlWXc3VJ7LkrqvxbDg+/RQFDDiuPFfARW+Qt2C9Zhs3nnqhWvIZm+eg8UX2
GT8rj0sK03DAmRYEMqXDS5Scro7JDf73MFnEJ2LViSBfch3LAnKB9kFVBU0lJHPR
GxSAaISwplgx3L7ebgnKMJQEYQ/whu+2AD64u0vHs1MyuLlPgXbYnUTkmRagJT5E
OB4ReBq7G8zV3Ro36z0YSfqeIDxCBp/1M/+y2GfgBKbeY+QUNBFZm17i/cYCYZnd
JAZqhE+Fz+jTYepGOM1/LIo3+hUDcggFoX7rI6Qc71K5rG6Dj3FO9pK48OZ8uA7I
5cCyzcTSLdEJhhIEm2WuIElr5gtpUF0FWRQiCRsIJLDEuzCcMzD+AbOvCsXnWXVg
IdBQ21fKXfjuiznNI4EfGCA6LqmsuenMvEKmt5gbHoIbgAiFjv5n/+x8TauCL3ME
XzNHn0nQtwbvY9VXPadpO7/Z89miLHrpLvZieglQjxsUREpnWDRfxk/yqoKQyvao
jGh7B7N40tjw1kWXnEqP61hx9MX50NAQ5pP+gIu4mv5aC/VeVjfR4H38jgsaJbi8
A9hMXBhg4MeugP01LVVe4chR3nuS3x/7CFoHesIwklZR4PbS5ceAsc9OMfFVV2HV
FAOP6vvtCzN93TeRrIAB6zixcCBlvv5kOyVAW7w+jJ9816Do+8iyjyGyg1Nsn7vc
lsB0+bYk4VhebLYvsfe3d55zEepfqaGoGPlBTxFQbXj8XAvXo3h0KU0CaIzPQ3Gp
LkiSVyAQrHt/DSmFLLIF3Cz/5z/lCwR6ui7a6kOunim0KECyQBbJHzUHF2wHok93
YUr8mgIxyg5QSitVhqq9x/wGorOK8gYLxMZqwJcIlbN0lXWJwMzXpWk2CN8LIDFE
MZTds9w3RoUnM+uvVs4/8b4ENQNlI9zSKMMjw9+a9tQTLCK3h9ToSYL7juD+i8jH
VxnXRKfxpO18suBG6wnSNpYj9suYoI11zRYjfRMLtdhc3N7qbkIDxHA52SdKHjaT
5rjTq4VcN2dEjeypdbxB2/gVv24LapYrwFPZfbAiyr7G6rIGKCIW9N5CRgQ0eslZ
tompS//xsFEvDb6KlJc6Dy3hvYvoUzsZuJDbqRtzMLTbEvzYbDsb0xYiNWYo2Npe
I5IK0hFpF6RpJ+k2//Por4UPyMyZsKBcYrSh3U5xOj1f/y7eGXgE8+SOwz7a0MUI
AnjSGksjGLf1DhqDcl+cTgme1WXFKrdzyjnRp6bVbDHn47DNJRCdHxETWYEoI1vH
qNnwOxU1qrkPeNPSfVsvNs9YKnN1QIZ4rDFsFWlr6WyqhFpvFJbk480eq74bKk1G
vJVW63qlU6aD2aCCE2jz4purs/Va2+35SjHRTpb+xurql4SxGboluman1ublKAYl
Iw08F98SK9qGHgXs3h7Y4E3Ze+uGuSRNY+hIl1sbVnjnqozYMTvXFODz9JxASyWi
5lmcfFQijRaUtUUm3+2ChcDS7q6DIyzsfbviYvZLg8hZyaO0KgRpirrZ07cpW/K/
+7wzRTfTPLBeKZzXb3fPJYsH2dQ8fOwgM3MO2GrkclXPsNIjxq0GbYcjz3UIOQmj
Z6QmR4R6gU+TYt/8oBSc7HfALs9J0chR4iD6CFB52OPstdqAV7LiXNR4OoTP/qRR
O95EB6u9SXZvoOuiajCIic/CZBPY5f/X/AZQIdb3JypP+Ru84GJYW7ARh/xktaBm
Z5knNHM8RZGkvyy/BO8uuTP5dIaFiYsmtIdz6gewvADkNpRTK+7mWXqjSHy0+WpQ
s5utlAv012mmwy3NZHp4xccQ0dvguldFe57u+xeKxVMoQXmOzTnJaYrIaC6EN+3p
QX9+zwbgbzoQear66yop79oP3dBbIL0soa0ho7WohFdsyUNSuPdHUo5J0Mu4ovzI
1F9JgWGR6nPaZJMxfu1b1hVp0+Y2WS7mhk6s/g28stuHJ55B83WRfuPhaxJyUCE+
8RAAd9fBigdYV+i3T3xFQ2TjrD12tSwu3UaHoj3iIRJsDCk3HdwH41toXibPWb1+
cOadAZ6U2ovLZzxQergO81FDbLBsKrAQ0YUhujYI3wmM0gm/uLUO84aY8zjuIx6f
/JAw2McPtrAtrMXXNBsMUo27Kb9CWB9cB5pSzgJGL1mrUbdSl9coC5BpvtUzwxud
GqWo7hu27/UV6BMWb+8eI5WQ8Yj4rFkfeesyRDYDT566rI/0I5fLVWQp+meX+43r
Cev3fXV1NxZuod7X7JoRu4G/pq8IisOINt1YZCJo55mNAdp/wmi2WwgJBIXfhPx6
I5F2tfdCxfwPpk+NbV3L/7AwOdP24Uzkiq0SspuwgWIOx6X1MODB576A2toAJ/xm
+IAKps8GIfGG8IXeEzYT0Kg48f3AEyiIbHn7BplU+R6NkEKKx+Pw2Hi4vjHiaCW6
Nsp6/tpwS0raMaEZ0ZIzuDcO1NGZRmGe8wdPcOywqeUGSC8tUxYCBll7bmexwOKi
ekdZodoqSWOJCP5zqIrEgTVSWHgyFNxvERXI4R+kSZRCPk5KIEyM49gB4niei4HP
qk7Vvsd16ZLp41qbfC0TEvOZ0MFLvASiyp5c6LuTM/WH98j9e3EN3aqk+PDl+gDH
eQ0Y39tPq0fZvQMI10eohFuPoTtB8l03/0J22Jwj3SPTwdAQUEn8SqlZnbKd56fS
dQgsgXHQdzMSyO+dV57L8G1GTnevwx388Nnvw8t4pSXt2NQEXO2COD2awjebmHuD
Re3IdECT+qDclgooZ4JO+v56bcgq7r7HRdnT9+Q7V6y4DuFa8lmySfcVRMQVujQO
Z5wJtxk+zMxg7zdAh7pF9JImezawUSK+Rcabh/oQiV/o4mBXKWUzxMfldN1LuSlD
4DAKnKl6dWWhat0/bIi23ZlE+C8EtzyL4eFffmYykC8vE4gvXHZ1rRCTnpEGBhgR
f7bKUIRRmO9QZAJ/tHF4KA8i84CGdkbG/lsggMcOQPrMETY7EihPEik1PHA1YDnC
KTHIG6ldiTbF3rns8/vixhMGfjwmemfKjtPzN9eMKJstCvpE423jni8p+TBYzT4s
k7LecahDQizuWdtmoXncpsN0IQYAKGLB6dHskOSi35LHn4qq7zVpppNRSyTYmYOJ
EXXAwATO5FgQ2NeaIw2qPJz19QmS3Hn1dfKEXACBYsiUMZ1M4tbxgcMAHmOx12VE
Ft9ly7ii+aJJk5G6q8IqS5+918aXg9oeREXh+UODZabK5NlgOs0UbXmF5+yQkn0O
UB7X6xYCeexhndCd1Pe2SAayV2cpeRhT9nl5zw6Q8QboiMPovT1teF8lR/8QDUZd
Mge3rPKpywmRPePS5EdM+OdS2MxbchfZEMvtLqhnT09MWg9HuCelzl6lN31Rc1F0
5SPrJJZp8aF8WOnwekVBPtGtzrTFhCYBO3fpcLVnklEYlpxja5tkAankufCkCvNr
tg1zyJOpmXb7WUMN9EHs0Gqss48vEkx4Zyl4qLOt6OeKnR1yV9HMFTewaNHEJPj8
8jtr8yQrqA3VLIBIGQNPBJDP+5d5QN2vealklh8jCC1c1LfNdUitATsv5eKMh9e7
77eer7bRPyjxz20j5k/esC9Ss/4ZuHmW0hOVwYHRtE/BHPH4mUyAeQIOqyJzIC97
M//4FN6C5TcviMO5x/1cyFw5ty8b81IfHsnwlVAacJ/RVntfp0xnEx52MNrIGLlp
B/ZG+nAdJamU17zh40gc5/1qbGLscY5o4mDPk/H6/mmJKfmC+0nY53123OIt+2rF
I5FE5PwzDaMSYgLzMmvXGLu35w5AS3kkfmW81J347/qEJ2pbaBvuC+JNhsEfQKPB
8Gj4W2CCJCXFoldfKcx/ITK9jv0wJ/fQa/ofaL+kMC+QZnM9Qqo7KBQAA7tIfsR0
i/TiR7+YK6M+77bzG/MwH9jbVgsryARftAOUIRoX6Zwt4trrxYlfcsSmJaDZ0wsw
dkTEg3fyYkA0rrP/PNYWYu6nNOKKJur+QU7r/JkgQf9lHdx/FGLfwlnmOghtWUEz
+i4dPGLCvEypiNfQXj7nezE5Xx3YJCyaUyoJduLz4CszBZmsMYybJflylYXXDf9P
Z+1odvAI22YdwhpevveocSJa5C0bYk3CfITNoSQEi1if/tRbqQpMVzec5tCuuk8P
/bqghl3CIhVY1cm64wALBxCf2tJo0IWhckckJlSMfLUUh6EqcS9fxmmZcZ2t5jp3
jyWXGpgpxi3aQkM8+MCeJvGA8VVOZUdYBtFhphBhhrh7S1ABvOQoXi0P39Z3J2Og
TgjPGs5iM2zk6N1j0W1/W31s1tX/4d/jfWD9QxMztyU8sF0PwaDSQ28kFy+VKIYh
4zlXd/1U2N/IL6l7H6x2MyvZknw9KtKVwLbQqxslbkeRAYWAArrWvqPLgnAUNI1L
Nhy/LkVR+ARsFxoI68/BfS7a/fXrSZs4WSTpZuodDD3uhl7EEXHd9wcVJX9Z3Xsh
EQIPhK07TeKCGS4tfYJCu29IKhs4YF9q4o9FRBmz06LK4UCSTobGN6g6dMuty8OE
yA8S3lnWPHH4TtiWQu7L9Gg2uplgQUBoX0ghp+f0hU5bzUDs00m00M+/Pz05+dw1
nSyaLfnTA9CPMAM9TDbQ2LtSQQ2E6i+Cqb+dLW2Oibfxf+LPVohfcwBDRYPJhS/L
esiidlwvPOJyqXsRalnmpzZXOuM23O5TnGgZNBVpWOyaurk1vxkSrfdVlj7X1y2T
FweAf0lDY4IElzTEKmXNlFXPoWbT+XGXGqfKM2bXMWb3PuSkBL9NcXvw11ctOycL
4FYOHOEOR8qE5s1dvLvT5k2wDtdZbgt8DaUrRTB93hB/rhU+IWI7K3Mpab0oGvvH
pdbmEwmTA/0+4vIx6rGxjjVnh+Znm83Luq0PMZ3OtIgxe31J8kUJFI7F0Omel+li
mJAYQQavADXcFgydPA/G1MmGjNSDtaiiPa6rq3K1WAgQ04jJPaZYGMUXKxoTo1JH
R6Povb/P2EQINr968E9jutvztUbYYjsG657w911B96x6N1r841l2lxBsuUvyYWyS
myNE/zoofgHLjXnbJUzMzC9MeL0+tmT+URl1BbHexCD9AzPqWmRbn9ol8wgXlmX3
BoydZGa4hKYI0AEpW32vMkv6jqFqutSFPbPd6+pPXbSnMcOukdDp6W+khnJEiXEL
9V9T/HkF6sTeYrfJN+ktFDGUtPA6R3CyyHF5BSyrt7d2KZonYGPCgf2343hD1JLv
+KFPpgi2oPUDM6l5sYoZc66yFHlMsbeTvYVPxrS4i2gH0Rv/jsCK4fGLQPYjXMja
pCO/KZIgc29jlN7oH3w1otOh3fQkc2UkfpUnLW5Nbie6yUeuBy53u0bd4plUuRmj
52lOdh4znoGOj+QWYrxRJvaMHbPSmBiL3ItHKc+L5cQ6yxTuMgQIg1QgdLBWrAEQ
iQPGtPyZTfjddBRC0wSDctFs0Kuv0dKdOLyJt0leKWaET0O+gGnyZis+VXRuDYFy
vbcW6lfzZT6cBA8q9qHOfaPP3H1UPAoPYLBLLVaJqRx12Db2WRBnMd8zFCdyX1VW
HnMg51WeTOa7+4bJSh8SXlRm81nKhHcrf46kY1e2sfoIfFDWmFRi6ySk4yS1+p99
cjQjrVPx7gC6huYA2kWzArWdV7AzCN/+nk2fN+G9HeRDq55ZcMkIfVtlKsGGKXAb
CEltuz2tuxECGwrS55w/+XDFGvhxRG50bxKhjVrT+1SvOG7vRsF28hmFZnxEFzMU
3xHrX4HqW3yKFg8deQtNcPwfkibShH/UB5B3YNrCdZcErUt7Tc1sq9bsIaUL4tNl
+GU05x0ucF1jiCSCgW1SJhsNwcBxFIdFPSoRM6Ojjkf38QrDsELkRsahr0KsqQ3J
HDfv2ByTpxlucvtsdrWWtt+vq4WGXn2IeDlJq8KnOApB0M/PnyeVruV72XFnCdO4
ROsDscvkygN7QSI4I0djjhOqPHfrvR+irjwzznAamb2UGnzD3EolVVbzX7WRHnsc
OOOThykTKNDYfsJsl/JMvy6FNhTOze1UYHNs9N13R6M9Oy5f+91fRaXHExZdLOPz
Jifdk1bPi7S45PA6q+nlNAG279NHWIIEA4zZVyVlxnd+0BixnBlbarmGL31T0tIT
OjL9G+pV8MtwoV/bWpouW8cpvxPvj1VwKU8opzb6B46TYFOCtk12tSZnR/jShUSx
/frg+rnCBY+697F/aJYaSK5MOEWGikVnTMSm1/HZBt4TLOsVpoAFROG0VEi0q/sJ
xhA7S/cPsjC00gG+uzmzVMCLecGuj+rzKSUbhBFgrM64HDoR816svRbe7R+elI17
Nju/mZhqvsr/ccY4jJEhdhdN084DSWzATcu7R8N2lHawwopYyzwVg9l+hf9Hxj/n
8hbOHof1UJ3Zg2a1eQjFLx3ObdMp8PN8Fn2mez2d7dyfrXNuX4NXEMY3RgN1/WCS
NNYA/fetM5Ji9D1JdjHJIzWGP7qM+fDAUNJU4f5UEwSKMoiOgE+ewKoxxW/SFF50
lKMNqByWf0a7Io4oSsXwxgg+I3TjSeIN/ikkUmf/j63kma2jUcfazHcIPSN9iLKQ
0fpNLlkoNWB3RihIHh8Rdtz+hthO8+K8O5QlSD15ZLOtqthu5rixsXYBVNZuN8Q0
lzkEp+QXqG4eF3Q6AErmMAbx3kydoapS8s6sv6EC5zxDA7Z25cIYtsAbD0kEDgvO
pNetXYSyFbnBsBcr8eOMdJyeSWRW8tgaD4Hwb33lGCd//Ps+m1jCZAIjmEC4IrGW
lKeXlo9/t70yp/OgjPZ2QGEH+lH8W0EES2CRxsl9FNJFle6wM6XoM5uNxbP078Ee
tbYXvzV4nFr9QLNlEFQWvgFJ+gkVjwqQ726gIMWvXUusGXmNOVWvscDe1H2ATMmI
83cT52r+3sonxjImPk5QKWAOmNc7do2k9gri6Wn4f4RSfyusbSc3enjgcf8ES6T1
whbHJhjpvGKqkrFv2+s9gTuyF5BBWJKzqZQTH0RfF7/1u6FfM0M8db1M/Y5/vySl
asP+E5foh3ZOQ4Y4tDGwClx3iPc+u7JLvWaGGvEkcdLPW22PnxZQmETFrFF0/RqJ
3gX33lOtK1BsC6Jb2TyXZVRbNyZHsUATOzi6PvRk/8v6hCG0nheJaMqMQq2gsuCK
+cxXc/4HIBkS7ATJCh0tKp2Sy3++eIjkUCdOFdh8+UoKHgufy3KDfO8fLbHpP7jK
L2RC8cFOfpx9CuMyOkw8GH7tDsyEwyRKKVu/Siw/60PmJrY/dxkcke9zm2SFqmgV
MYPLRGv1y1vYRdXSzFMTNEMADrrDUMMlydNjF8D3GPvtht+iuBS/5Fe4dkZQzcq0
LG0/+ylbHWGGw8q7qcRUNgCKHYZ/Y6MRKGHSwaObIJ2YUtQdWYRZvwJiQblAJvzC
RUV9K0u6RN2ZYvt8dW+s2G1nedOLigFM2N3koXzXixRSqquF133c8AGQ7fMLuhoF
VZXHBdHFNihCsRfx2HFTLHdZKXkf4sWCIuDKclARN3qpokrIwPzZx4NVvNSaYgAE
g8NHY5PHBz5YBtTEZcJQWDhXYZvWDxbtzESnmQHF3c4wVi4sJqqL/tVyGpxt+igZ
FS9dWx54Bta+h6dpQISKIf7jg8mH/VpmDIU6RJM13YcLrmw0786ipEQR44kfK4Gz
JzkwDdfpRzlp7HDc+KVcbX+dpsI26GpLTXdVc8a/njGpi8uc78NxHQUbb7U/Y2ez
SCUARqeqvzvKK0BOhQLfsP3QN2mh1/V3U3YK+5L1kNlRVjxsGJUd0EB7swvFNtBv
MDVwpJSZpsGYi4OLuUwfCpDATaAifjpniWUAvZQoPC98GNdwUgeWgINtk1R0UboZ
HS4PU1q0OIVb+bDDcA8K/kEqVrnG/c3mexuORpQP+TjWMv9ww2aFg/rHc/0cRXuO
9BmywoV0GqS8wdwTCMxE5yWEiXa3mLIDT9OCs+DgsCDnyylwt9vybIuYV8K9hnhd
gsVB+WzqC3GN1ZF+ZzYy17ccBfG6+2mAYR8ttLTkTmzu/HzynNpoh9vtN7d0hfTa
zOCqGoHUI5YDvdHQwWHEHTSoo3VnJIITUlscEYCJiPg12j2G67Lf/5NHpXGalSFK
W8jrrdfllJCz3r3HQcNHQ2Mk8sxcU8HKfLNSSPrGpM3aY9ztoukSb0HXYKXn45AU
DMalwaqHlUuQca8Z9ccrEd+I11SOvynaOQATYWdHSsUV4IGUfIe2/QoJPz4BvqwT
Ng4y4F8cutURPnO0NAXZotMTcm1nncgDHFciGKOISzNdw5A/TVDgMvbXTczJ0m4q
aDsP2u5Zu6seyI9E43jNwme44PQUG23oAnYs9Kq5ai/xCe0elw5E3wEYzx3Iw1fx
Cw9cxOjWLpDJ/QV+CoTuM4T2U8rnu4Fd5D2MeQFV1rWBBa1J4wUJkpt1Nf3BG822
doahm44+x2BWd6r0pj0E5Y6wJaDU9LhSGg9NnWuAWT8J8BJrdIDlsBsQFzFlxfPy
+62MJHcMGOXjC3kkIgc+9hA5m9xzM4vVx+T/GZpCh8a+5P+KYEO3fpJASeZhLmoj
HbpuJn27mC3Ifr5+NtRqOFfZ1WY2wOjYufTjPyQ24/CGxtXcJOSSU9sHVbFUYmbC
oElMjRO/G1LlSXKTCovt+ZCrl1mYoue52qpgXwDXln0kRW7C9EBB01RTYQ25ARG7
dnulpCQ19FOIAc8Yq6hRr9K/Of8RrXIWCZ/duN9EiImCe4J09F56Vlsl+v8MN/G6
P0BJreAJcmY97SHuGiXhAUq3eQSxbC7yMAxCbJo+NNh0Xx7ruGzxCBhKIKDfJKYm
Kj1yM/Wn+RCSVz1nyjEcNx43HHiKia2CsEwZrnTFHBkAc8/YXPC+eSQRTYT/OQW2
azIyXvx8RV68aaTRIs0/PR0aoAYs+mNFUDpVf616lBWTETwrrHx/sWXAuoaPEOv7
2aAV56J9q5awbXEAgAS8UQyMM2T+sumoE9ItRryeEFOmAat0+f2NIsy16nqjm4lM
YnG3VyY8yqLZ1V+ikO+2HjhHJA4xHHZzumxT36whdYsSdjOX2BH2rzRRSKypOIch
Ugb9YBRsRt49Y690z4q0BlYri17JqHKnGqA/SzD7J0NtR/7HK+FGLafwBPpFrUkh
+oMvajpWfYVyYxzD0M8vlDhes0uBmgJ3EmpAgr/BGszGvfmsKXno2uP/2G0aeKA8
rbgo6zGEl/PJRPyORjNkBv3s5NWo61bjzPIaBYY6+9oFyvA41p3GOWKumIr7eq/t
KQFln2BibQRhOALQr9JAxb7ahWFbCnGIckAcRZoqkyge0lwM6WBEtiBBCXDg2oHR
UQjVZBmuOdXFbnsjp06B3iV/r2aDFKYSQUH2RO+PSRtNBc+ZmXF47f5s1WNREOLJ
kJzVQW1K78NpHk6oaR/+XyPYDQGmzKSCHLX0RFd9pQOKRmhP1zUksBUlil1/KjKe
LEw7uvhWcSZ+2G7sdd1e3UfwBB9rGC/iyIpMuSDgOY/S9WDBjQqj8tXF00wGMZal
eJjIX9AY56ufe0T34sEtmtQjpaWilZ1ZS+RsDkbCmZrznu4PawQa+pbsRkuCA/9M
Jdfs1jGf0AKS9+3r0DRR/Xc7jVZi17IdSFAqQHUbahwETZXsK/8vZGHt4X7xY1Pd
i5MLXMfHuWvTd9mJw7N4fH3YdehN+or8pSoMLmlV0jPin3pfnharojlnCEtFqmb+
8VO1Auuycqra9GeSBjtfh+s/mgIJBsSkWZC1VJ2JUvfZIk2TAX4BbzrRMggj7mNZ
337xY+MNcisV4qRfpCuDTPStJmkk5Qn6qFw6TM9jcYjNY/mhixnUzjLQ8bNaCbNi
wp77Szrs30y+nuBN4tfjHuuu1iX3bMYQE9b4Wy1Wh4L/KTutZ2q9UvieobT2F4XM
VL+V1QSDu7K8EnFZAU3R/+ee+KSPQI5YJgNqpE6SJs9BOqz2uzLx7w+nrae6tWD+
4zoyzHnkghnW7NvSGMMgDZGYdgq/YI5nbgVaW33Vpwlse516DaZ1FCrW/5WcrfIR
/Br2jIbaE6hc6Nd5uRBjewVLDNsGOjF/VG1cO3yioLUzhluWiB5vNWo7DcKwUkBX
RP8NsOhT+C2IGp61FVlpGownzYgckMqFhbEE3iaeXBVPfY3PLKIxyeHnNmoOuh8Y
UuH30DAKUXhhxn6fuXI4vuF4t+HiGQaQ1LWnveSqrYwtdTlcy8JQotoyxXahsTpS
gFM3aR8KUudyDtLzt2V4D2hblAPkFdeUQS7vKXMlri8HcHJiUClVGli6Wnffm1/1
I9l0jbgecDbp0A7NHFJ+QcE2HvPGkPMXhrUby0pK/vfRJ9PZx04fXF6xc0wnX9bo
sR7OHrqsvyGD888L/Dd0fKuTPBz937fVpROwxRHeY9sRHP3tUNruH3VxbGVDfa4w
sANBgAq0cXtalJ2apagNryV4YPqPST05we0kPdjI719qy5HqkuKw2v0oBryyRwYA
s8vdKUNlul0ARJEZIjDzdPBC+NXWJQtxk/bOeGfqIPRKmcNetmK2yv/RLxJAEALh
DxtRBaOh3C3IXqYEyFCWcCGoCV9YlCMKzLiOAuaz+yC8a5ZdZtsRlfsbbeFr5nl+
2h3Ou+LC/+VoeP6e/nZMCI5Wv7qCj+lCmDLx4sxZwKHN4u+1VLGrlNuQEspXKpJ1
7dhh9uIb8pDB0cg7BGIDduevkL/mmW7BIC1yx6vStTInBOdGYOI02VAFDblLRGFY
1/fvxD0d7nYPjSbatI8PJm9YGnisKFLQ0KW0Rdl1MtnuHaPLH7wRHMkltRGKYGNC
iHwMuuHyvCErqhyZF0HP8La16BSdciiAOo83t1Lr/hXoi+3UwL+qDqK2+hMPAK1r
IGBMThdGlPKRZPZJj3QNYAbCLc1dWQ5TavjAUjGor32bfWRDo0Gx+TzBlun84wrJ
kadVs8nhjlAnN01g2VYPkrbcFsFAwjtT4U4G2KGZNsA9C2wjuv3xNApXF8iyzU61
6VaoZSmQv2ZP5eXiEg0KDebo2OS6mTYsJxjLZ9IhPvpCMUUbmIqlq1oBzDn8pwti
xKO6GrNVd7cqZILZBFk+f2QhOXQwPRuxnCs0AI9iyCh7m4615pH3NbKvUVfvXEif
QKukS1ELfC5YCyjpcOwUFwgfySsaV77uCNitUJ3ShbUH59ok6esEoVi+8pWxVkNS
oZlT2EnGIsXViG87edgKhbLT8keztA6mP0ZYAAFBSeduLqtAnUaVknHpABRyp87d
rSmL6qB8h2vvSMVn1jCkaaKg5LGuxEH/pS24tL3CbMgQu/cGRBf+AKA8CRgnn0Je
l5jV7vGLNL3JCbKLtp8kZvy9to7gawNpn3CLPQ+3S11Gab1fX44Psqi6tGWKZ+UD
+jCyg+EmaFUB7iJY4+nNDdsGOZv6WzcrVoVhpUtC0pI8Qa4swTP0uYtC34scYDOi
MC8TilrOnni9MXid5Nvo3ylTgkU+hIWA8VDxFgpx8rcr+GYfVbSRrG72uvVyjb/q
LuoVjRnA9HnyfGvufWeRkpARXq4F2BkfPEWzNGWA5n4beYtGw5B78VaS/jcTULoM
IPAiXrN1ZhB/cXi1yZAhF3/PD8F8c+Lca9AKMWpN0jIRsX5kgdYZeKH0VNwjvYMB
dfBEmQJ2zbCwrlXR9P1cT+iJHYHIMB+gGia1w/Onq01aL4B0jpVdQqJxXT/4FwR4
NWM/zX3vXEpC9aerAHpgSj1r+hyhPodmWWyycvr1RiJ54MnJUxzB3gcXC4ApnPQx
jrDm03ZwR2hmBhPtDm5OXp1WBzv3/zHcSlAcfe2cv6NfLmGj4YJ6phFW0/av1LqS
Cbe4Bu9SB8mBMYEg+betuENfX3sUhaoD7LgNRPHhJ9ZdOHU85NLMU6SYwKVMlDkX
QmnujrtJvl2PGv7rtXhvqr2dI0GlVPwoWhTDxXySMGowHOEJ7fKnnvlvYFTJZdQz
l+vJELfWHHL4sMUm77uJ9RbZ4YSMzm8mA4CY5hsLO/VdngIaw0FHnr6efK8wB+Zs
ghdkVS+w0WklCjFlDCrtvu38DZSZOrcujws/ENS5XQLr55hRALFy1EIBCMaLCklp
gJR3HhH+iR8Msk8dzF3QXXYtH3uIwLclTRLyipygg85mbqDEKsmBk6VnWeKlBPxR
xLD2PCncdAMEGttREJZhINjlW03GbRg+Ds2Kf4x85T9Y4ppg4SrPUDglG0anlPM/
pEgNakVXSzX2jd20JFHChIEie2RY/9h2iKCtN7pjWScPRvSf5F6OksP8AswPbGek
x2u0mP4qTTf7TGlew2LjD603e8mF0jy7UV8R87B9Oz2U2S7HPHrMwAOF9gGoJ5np
7D4QKlhP3j05VHYwG1ieIxLJnmQ4sHJfnnVvyLkle9s+Mu7Wa9XvdxKh8ZDgd3/r
d0eVokVMkdPa8McsNNhJ54mpZk5zH0C0Lv8mFfZmDDvkjvWM3d1cKskh9oT5JRhW
Ro14nEksWWpeGlAXG5NDhngYKNnC5kAjUTSHOABGMJawMAEFCfC/sSdWDgPT0a9b
uIcglGfNjy1Csoaun5dj/PiC0z+K9WpIM+zjUDd3gyTreGaMZfnu/f/tB4MB/2Oy
Ch0eJuA6SfYzJyN3Qg4p6/n7dWqOUxybrZMDomdecsPY0DfFDjmwxaMwwg2H56W4
HY6DWl08eJdpz1vzMO+hwKQd5WomUKCWCSaaZXtKZQNW5OCRpx+CbYVVZbY5JFEc
Rl5g+P0i75SFuQDq7C/HBIsk3FyErqGTEu1Gx4x/DP2CcZ5qdVZkhCWSbafSb2IX
GbKxX2GvXy1zUrpw+U9byOY/MygBBQvU3gHWxA0SW1l2LJdbY8l1B3LxToDh3rgS
D+Q/k0maYNJvnEpxEC8Df0qOgovnaKxXgXi79Wkgmz3iJ9AnH6lE2zqtEMpmF+x+
JsBnBtM5OP8HlVP16GwGvjAUrwNO3uWoe6iwoV3dewZbnVmjMeFgExPP2rrmzmMO
aIzay+JLfgeyvznT0l/BWhwXQy7xEQp7dvOEVc+2d8By0eI3mUy9z/vIEPp9bpDN
wSs/8o5IbnINl7Dui43ZAteqMFljGosJVXfil5CL3P9yQ1mRyv7Mj1cs1tpjAWtX
XGfHLDZnBAP83iNsCXJ1BRPpeg8uqUkRjW0hT96J+s2X30npC3yRULIYiNXvFZ2F
myCg8Z4ON3KLHAJXzE3zOFSUzGlVS+tIPZhHjZaWNGygHaSKa8AlvmL2bb5NIK7H
jBLZKlQtLH6y3uDT55rPhCV3cBM8YL/GGUgk/JNFnLhmrXw5Xspjad7jSuF9xjbo
Pd0ce48VyBw0vyW+cmBWWVYFe5aRHuUNfQH5duERQ/pCZ52GHn06C0EL1DqrrdWY
SILi4kfTMLQGkie1Ow6Mdn4RyRzsjPcY8aK0X6FXBBxYVps+KF8DsYvbnK6Ip6MF
eyer7U/dqdWLuixyE18R2K9Am9I7UDpGD/fLtEIfvM326lP4aYUjsaS3KdA3K8wz
83KJYffMtBD0n4DXKaJOg64fRGiqwaknrt4vWm8AdnebpaE8uRfXeyLCkdqrl18n
zbAAsKAJe6vwNVqRxC0o1YS4xajz1/yaz7uU1BHCPsh41XB4p2JAqBgyKJMZFIjL
BsOntnegQ88U9F2haMGVMQB42XHajQpmD72/XperVgldoqvNNzlECkf2jTT9EBH4
lpt8uQA0g+mZ2ThdMJTQi8JXWEJKp+qNiT0eLwVO5xvgoRrFHn1YBpwW6IoQeuiV
3evWWf08tcY/ufjqUNwONK9qZ7QGv6Rmijij7JZUzhuUVTd/sjo50yoZE73p61R3
P2zWeXy2z3g49Wsf7JExJg+lBkPbkJnclEA4hS0jPQKjFzr1cK5m3LcYy3Hb7EPC
UkN7MJANfVStOztqwpGW9nAYQ9PNNjXaPgpP6rz8s31acWGG7rXaC0xn9NWJIpli
mUfQcgCz67UOvV4uU0IrZGepiK8cmP1uetL1ROQA+ZNswyId1SQZPBP1GYPiLpDY
ZnvyCCHzfSkWH4xWVEfERpEcTRHK49c98O2fVDg/RURwQ1oNMAfSe3fNwHGgLg4e
SdWKFOQHTcQHp9nRljJeAMvMcep9XrzqvUzx//tjdaAyxl6SX/Fo3UD5kMJtfvO/
uSDWutes5f2srdefA3hUM7wEfkW21yIqDjPG/U9q5XPxaP68TczBIviMBrDH8aZS
fhXl3ljBXkybZwQtgXZUTO5LcbF22WGFVazwwdAvdbFDXPLUGXZRg3UKquLxb96W
RwV3zx24Tla4f6IMQSr5UK4rq/b1hDmVMfqRsshwzXHR1XC1Vv3EG/ZeMeX4fBvK
KFlGaz1tdM2kEiEa/6wvQbQwkGfziq/8GXy6iwkgNSJV4M8N/T6OplArVnMZGlds
O9wfqKLYevAg+j688F8qA9s25wigScBuWXWt6j0tYGPW9WDAkBxDl8evu42FeXU5
mB3CTwttKkWnzTdrYR38q6/bTRWKK/PqGpmRRPmR0fhwIQpZ6qN1PCi8EZeAjO17
YyMeOZcwjNnqbQa22FCVM7p+2IVKfBUv9aGLkZxxa++riqi8Hvsp92xLvFQPe18C
//yB2+ldZOJtT7JWjIViDb9EUMn/o9YOE31pdg3c7zQzq79+zfxyo6ll7w4D/j5v
OhxMa823k641aJtnqWJbDZPU66dCEJ2pIwnjk68+4yiwO1cYVoSXuhRBKIkjhxDN
rotZH05k3o0NcbxP2HBc3TZRbxsGsU++mnQ8cfoTs5G5gDVpkwm7/o2Ebr5+QYzS
UpW/4aQDwgBe/enSliutA8XCDY/dO/oOWs5UDSvdcNqtIbE6JzKiJmvzCZraGjtj
YsvCueElarBE8LpN99Nq+GnglCTl8wEFNRta0H0hLHMIgvk0LIn8MamRjWiwB79m
XKjeTqU5Kydo4FMFFg4OoubFpGWPi3xehkQPbzkbzVaBIAuHDpXZoZUv4HGBnksE
g44wtu7nj+LBbtTlkpvk43+3tDlVlIQv6LctFCVban6sgfxnRmHS51UwKBUvgrW3
ZdDwNaeAYMqrWRzD/VLv16ohKKRDJ4SRM9bAvWc6TQ8tBfgXKCOHOBSuVOwMZrTc
fwtZLl5nc+hiFtvpb/9CN1OTR7uncCWWt5YeI4KwyKYM5Y0aa094FFNcwVCviuEK
Zb5S3w8L4kQuaJMxSVsd+Wgyut0I8h8rSgOOmnug+xFS4sPcWevVDHWbe1PKbB0u
/CBZ5DG1I0BaMMMRHx6sKXoXiAHrpqZeP4iCGs9TZDAThYVub6XSyOaiHWeDPHtU
KcEkr/PL3FR9mxsfxKlpUdknJ48CD7tHRDdlLDwccwPB70WhD1Ti3rXxYvQQSHWT
7E+JRFttLLCtgWiTAgDVRPEUgLBvwbFV3BoYcsGUbEtwoncN8ANYfTsgDW06CdFh
VXwN65wiTJqm4e5FbXoixr75kHNpWZx5+dJrpLaCqnUB0ZxqzcQ+c/qA0DcmmkLO
B0Rfwx82uKl5S8iG7pAkCXGV9t6QkEMxRsVyg4N8ZGwN7SDsIwCm9KTASDJKWrsG
8JFCa0BHgCSd+kYzki6akYzVbDHg89MyJ4gk8xgUNbVv4D13iTgIwepTUipCkE07
IticJ3C+O//V0ug2fhG5dBo3XhqBjvcYISovebkzjYOBhT81VVewgmJ4S0rnEbbi
oi4ZOxQ3ggGwQxcv2kyhN2IbiSmPZJWUm+s0GB5N0E8oEeZf5l3gGkQNJaqh5Evh
DjfHbea4gnBjf3TLXkFs/+KndSr4Dtd0QxREkHWGWgvSzv9XCfC65fiM7qP9Smm2
UvXKVj/c5/xIL6DX3MgUSi5tWb7LmkQo2ykb8TRxIKurC2US2dY1owgO/7TNr9IK
L9OnFI5Aliul9fmiV3rt3VTXjJCU1G/50FrIs3ihzRePXk09NcDiUBa6lQH30hZc
hu5RzEi+lFDiKkMvBVhEgi1hurpud5NLrRZe1Sk9YLuYho9GphNoMH3JR8aEWflq
nyHN0Apm2rwqzZsDuQvrye3NQ1ai4P2Amu65BKtTs017ZRE4Uzs1Fcm9HYplpYjd
M2IbCghJGusfTdiJ5O9asRKTDD9Y1OkADfjCrRno/6SH2q6Uv0lzJ9s2FbCcYKyg
ApCs97yGxjhRnTmQYxz8am+hRO9MO4aI/Jayp1YVKjKMPim4VC0rMY6cD9EzE/VI
5TtonIrxOU/1Miw6gzul92S6npjoV44LVeY4W1l17SaOSZMPjjfMCsZcvYo8bT9+
C5dsvL5uBHypS2iqe6BW0XWNx5zLvr3+KcDMWlM7eBPVjhPqcqwf+OhVR60HCebw
7I+xPIlus384lRD8V0wfOdiXqTQX6+XtpOSqwxhQGe2LabR9uvbc/WnfZ3Gcf+Df
tQyPrdLdNXhfvqsJxftJwDZ9HPXqWyaz1bvCJg8tU/xpwd1s5C5YgCe9InObgBVo
GP8H/+Qv08O6Jz+ExyPKN8oBnpdvZP0kwoKf92VRxOlB5pE5xF21G6jkZOdGZZKZ
NuKKZXKXfFxc671Z/R1A2S/GHqEzcZuPICgWMoGlyToWm07qnfsgiOPyhNUaGBBi
4lrbQvvqr6kieklwkO2SMK54PC8J7QsDhq6OxfokACEe0C9dArPooajUCOn1xNq6
vv1F0LiiHBHhE/Q9+mENY1aZmGkL/t6VlQCIsRmebJWCddQif6j3He2jJb3pzGB1
vhCSKhIqtpelnK7X3TB3RzCmcg8zoZNiDtzbz+DvuQcbQDd6KB4jhRtRsQxpAgQ/
LRbRI5dTJ0vkpHX78EKJBbb360UFzkDXmZoLB9GmqbWSB4MJESdp4CgBAabL/u+a
W0LLAQ6/EtpMpYnJjZ9hklFS59LoxT7Qa1OfMa/xQw3HjnqnuPKoR6nu6idb6LtK
z5kUlK2o2GIm7XKquqBQZEoxaWFH7v6ul7sj67XN8DMtFblh6wvC32OtUR5eFGe7
utSQCN7wrkqgDq0LOGbEyoY/9l41TP25RdeaUauY3p+Madu9vZ8azA3sig3eXUYI
N74gPdYD60aj+ptU2vnaICvbqqUz35cmQWJ/gDh3Pc+yINCbJNwAvZ7EAGyBdUjB
WYtDZhN33gBJ4u2UQQc5IOsdKf1GGccMgYLKvHbcMn9f5SvDrWTfMIImhcBwZlxb
dgqIYAtyNkQA5eRKVXMTQvF+Aa/M7FoFh0lXjx3ib6ynLypE8v8cCWhA8/m9c58i
lGjlzN+I7FDY+3EGOpp5J9vz1+BTqJBegpCvEa7i+TuokUbGcaHi34p5Limu/lOg
1/diVfr9VONouM9kGtbNS70Z/7DL2GQ0dvMPdpGKR/Ybo8nllyq12nK0qruqOHGQ
FGCNF47lCltpMQbzb2D7IGP0OHfeIuEwbVd7R43vTHo/RlCoetAgscQsMVzKdkvX
fSfwrqphWwwHNSRLvIRo8bSgEyHab8imzf32yKkXHn8fIfVOPCtBkln7tg+qQ3Tu
rZ00sU7dm7uH9ybQfubMSv1tvCJmMO0m9cTzTu/JiTCAeZKvzikcJ0/4sRKu3PE4
jIIDlhDS+mu3BKCPXT/TJmwKd3DhodfYy94JqlOBSwrV++EIVzq2Z3IXIQicoqdG
zKKC+U9Ksrhv7AQmYWLW/EYmwTH7l5Iu32HYK8d5TSL7pgEfx4vZlaw5fTqJvNQS
Tt+f9CDJ7G/DepTVffr9POiyE4zEBzGVv7VcaOwO9EaITVmRd4hXGWUrTpN8eXGd
Gykpxq20zP2AxFdfIhyZWHhI5/62tUhk1KVm40ymvrafCjnuvO7+AgfhXmDpU5gX
1EwiTYbsaxq1MTdFh+tIFz4TB9K/xYBsbYY/GjZhH81BQEau04nijiHOOAno39+v
7h0pd82R8r9q/kNjgoDu4KwFgNocrPUpUnZTA6hejuy589iZ8CEo8TKhRTk+n2WV
S1jgMkDJf6UXBUIh0mdOj/BKj4Kp71kygZtTmET+Xx0EYl576ZYPTipSZtoUUMsi
BUffS538wsgbqiVO6lQXfKRZoOi2oHh25T0mBKlvHJ+y6n0RZ0NntmOLZygXpoTF
8r+W/pDl0waYMrPVA9niUNogq2XonC1GsLbUFzUF80s7PrRP6cfVN/kP53iO4Lu6
HKP4/y/5p6dOGGh+Pn8cpzjds2QL6lkyh8h98QG5o0LyW4baJs7l0JxDWvwRF8Kp
wuw7cUXbckciF+GSCZJ3MRCYISKTLSq7JP7pTtzb0ASsehnxZtP3+uTzjLnpdAom
Lr90Ht4o7HUAgpf2SXHNytM1lpj/0pGsX60Rrnwya5YWbBtu+chcH/YuEOH6cJXU
onrGQfcSRMXoHHC9KJN+z9Vqu196XQRbK2VAKr8X1My4pLRDeL2ybvGpXUNz1c67
rl1AIt7evx9I6KgsXRYmVEYnnGiAEChJR5kYR/NCSDFp+FfLx1oHuYWixX+rRPN3
fZqmyUpck/ZF5HT5rBDnTewf0XIYQ+mt239yHq9hflhoRSIG2lwOj9SrTiUcNZNY
Tlh4mCCElaGpeHRBwOh3pp/OxyTAM65TiAYKSz4RgyWs4hbs70+aEG1MvM84HQae
oOQ9SoI0LOQRhjgBVFtjE2LWZd0UVXMbCwpoF14aRWsZA1MKGLzDftNC0dfkGBXu
eueRU+tchHxR1ckXKZZg+kXQgQR/8q08WiMQd1sqFHdiZsk0Z+2+r14FqN9HNVDC
Txowf7UxkLzOPJfZ1dLhTCA2Q15H62F75od7Wae98fD0N14UDqrMHmAYecT3kkbH
Has8H5qjAeUAMGgfWsERcNMzUg5F1W3AXGgutfTWFW7SpqG78F8AEdG8cruF8UUv
db9M7IQZCy0kqqIQ6tiWWpI7tLniwO/VFQxD0PRoAhfpwVHX/6Yrb4qzxjYmaw+Z
s2rFy4qN6XRRmcM09lERBHlj4tmxCa79gxdRCvbq0V3d0B9kJAk/sD+oq5/YO4lW
llOIwQODu9VMDtOkXD1cobmlnuBmLLio3GdBslET6fVicIy3KSaefkq546GR9Ceh
8j5xsSMNhs6sR5hF1Ah+OB4ThP1O/sLkbXHYwL9K9HFD6qeIhxRKCbud63TMOL3r
nV/fWFWDRVdL3rkCs8AEAMywAcx2P2MbIiFa8xKDsTUM/jAL4obKnDxk253JMJsu
fQi3PorXem0m+p4kCoEq2hF9j4ORZXFxLs1qU1HNbgu/xGhrNRhEUnjIoE/FCV05
isgSZZWyuFherC75krxj1uVyGoW3d8xlSAbN+B4pdGh2TX0oud5Y9tJcxW6fihZK
BL4279SMgKnvYziWA0oTMpdlYTJK1WYl6YZFbd+kuhJTcyvyhs2Qpe+uHtSLwjyz
jJTDkjtzY5gO54mdTHSKe9buuZzA1h7IezQI5yp2t9J9kkAgh2OPT0sDPg/kRnB6
VhvqSqT4MdPUblsFsKm/AvKjm00bcH/Ib9glSWcWh+bZal0nXaA6LJCQxp0rx16A
FJ/XEAWoUczYgtwRQEhddVv1jpLZHZ+Vk8WbXnTkVV2kvrPmPWeb2uP7mdUHMaA9
/DPhB0GoQlCJNn4KhNpVh7JvTjaAlXGGx5wJhgS4+Zku3Tv/CaJ2NkoTzL48V8rd
FWeM4MQhkoyBuZNitBVrRitPDQtXc794X4ojmUo1k7EjFoziSy0Y80pFVRkNrO/w
yCJDPW/RTADBUOo/Pgc/o6lk57qiUSOI08JwXSAXe724EXJ3qEZ2vvQTxpeHL5gc
hSgYNVk1/m94pDWl+ME4cf/UxMaK0mxB+rWJytVe9/G605edqIyC0I2jPCdIJxI0
4BwD66477M9mNgnv5aKFqGlmpaLkCvxHcDAYMeBt9Jk8SZ9hJtTjDMb4oZcdW3R5
o3VyFfLnF/5pmW80SiZNhDJjsOEI6jdggsi8Cv0L4cADV8lSpdKIViB0MbhD6kP5
wx9T57N5mQ+MGNgL0RtJIUOL0VpjIIjSIrM8oXP/fbZaSJ4KW7rMqPE/r3sbyQ02
HYaenIzciuPQB4gLhoNW9IJaGwCIzxNzcl8pP/lDWrbW5Qdt2jfnbQRwxeI0PEJf
LCvT2MwbZgtZhxr9G9+OSqYNFUvDSHUsKfmKpUmh8mOzf47CRxEMnr76TIsv1iv9
tlrgLh6vzJsP17Iq2ETRwQB/qKz+tRHv9ULAOxRagnQuPcnrDVMKJzYZhun/ea/8
1f4MoSnBd8Zjq3qy38xTXP5iQqa3405zG3c6vLH7s4zU6eqtSO+1hQlUVG4YuScK
zJxYsFxiRUcWg3Tks1TOXG4Yvz0mdgVP+QA3IhUceibW1PSiRe75KcRqpjKSttEN
wLoudHKCMJlfSb+PlnTn3Rpkxi1uDp9saqtsSAstASpLXqpAkENetCcbx5XCbNJN
4mFQVkca0gO7+0eJzeL37831pQkFsSeqCbqG7VLf2CFNE64TjQRW95Ihqxo8Cgge
kvaUEcN3/ghrb/LZD5eboQbiXJh4pZRa+ijqj56k8yRfDHDv3zAlFVY1QvgKcgar
RhOWKzRmMDcXM5qaYpYSwBclTe8W0z2+M9sy+iq9j4THhoDC7FRT6w7Xwuij4S6u
1n94mYxWRs1RK0XrPpgU3isR0Ljj6VHOfaTgp4it4BMpp6NSDlF9snUo6OjA2F3i
aJCkuiMYxbkqxCDH77bu+ukFJcizKqxJ0ddnI2wLBVsLt3YdU7Dcb45j5Hl9qylF
ENYvvZZYmutijMh7sirzJ3A78F+bfdY9TIulr/ob1okpcXhCMBbdhx7eio0W5KAW
McZnNJOSfM2ORVCgR5X+79iJZmKxhmfIwRmo29MuYUPuicL4iLG0VgXX9vNB4tW3
hoLUCuqD4ej3koDymVVdcA/LWs2NyugcHGU6HjQlkmzQ2x775eB9R5YJkEi/qZpU
TyHUgJ58iab9CahdtMqJTL94kG2Poudeejw9SRbzfb2ARk6OWSCXn4t8EEh/zxjD
A6mGm15uNXwWSojWzTSrXimV7yQHLRIbVXwXPLwGyf2TGL/tl43IBUxYE7mXZrAc
te3RmvtKgmpaMi/Lk+4nVK5mQ1/ik323HVWcMzlPU2/vD3sHhgBuCuxKlQft/can
KyH4MwvskNilH+XLelN/C3ee/PXx4AWSiP9dGRBOxpltABY8r1sQAF3tvo3Yellt
qegvEBpy7cGwd/BNTJtmib/2cfkk1UCqo/FNHyc7yhKw3BfDsYTJ5WMxHgQEzAh0
X9NyHKdgptyFMwfKKgaThPm4olzOpdFsrOs41GOxRR8uQeesUOfOPZbdqz7ZoM/5
5XD/hXbPNHnWTIbbSjhGBI8O+Kz1SXhRrZHNOcaxhN/Hlt/wwED85nNFLm/b3Ej8
NiST4Y2fDJL0R6ymcdu+MbORaxtP5PZhoV4lColTnRy7GEwwPVyM6D/c1/7pav5+
UdH9s3nIdcrChDGBTSddGkyF5/pj2zZzzA/FZDgI0ulVxMM/WBsImP02XlEjg2d3
GwaLchGg/4Z6HtYbjwVPGYMVly82kugaVnQk+U7jHk6zJ36qAwxTOdoq4wIZPS4n
xa2/wISY3XFr3nz2VLcVbZmeQJsgth5DS1uVx6S9HNLMbevEXWx41W286AWNIsm9
b2pQm2GxSWEpQ/oKpIxbSzjepH7ZFbLorbf/qYDS8wOVjr90LfrjVOJujLEAHq4g
6z+jRa6jM0DJi+cum1BZX5TqaHncHrfb6LaKIcajSfOeXUg3sCAWoykOCFHjOb9N
XYsvZPB09uDs0sq06kxR17F/9o4YvtV+KeFR7wj+eFXRtuzpWNbKhXoSOMXgH7sr
Gazsxq54+0y/3W4dh3U8R6gqOfR9hLJXMu+PrkZ7GbTTSeWM/t9lhiIDSDTTDRUD
l9Ytb025X9IR9zFDYOgjV2+kaw5C4gJ8u1fQ7kHLVVJ150LDblCvKoCAesPZoVlU
t662PbbfFbqe7ZIIyVGa+gI/Zun1gsEABh8/3Cl4PgvGMYokBYQdKEfbu5aCBC1k
vJtLlEqZJfyxb79ZQaojkN1+5qW+svGPRO5kboAqxG2g20kI/6y7BZqr2Mm33h5X
+8fJRtLcFuoitN3ML72xdiVULvQeg2XeffDNaFOjLFe34c0ploWr9e4MizqpXBJB
EPkhHf1apK07szz3IMI9OC/PWcI36wFj7XnAnx4Kr65seo4dJ073aMnByH/Khdhj
EdNPiOG/sRq3nJNHl1+fkPdS0ee10TsQKl+rQ8a+EH/naY0C+cGJNM0ipZst5rzm
vwh0mzmvh+yDeAjXmaLF3rmwOesA3TLcaY6q0o9cTJspAK13JvOatBOwUfgPSurB
EJ1/U2Hzr6q7E0q5OENWgSlqa9FYOonE2mljY2A/61mqNWncCBooWD+kCbx9jhzj
PIVtdgxPaIRNn4MMH0Jf7KlssPIeyK3Q7n8UXdtRibVUwtfg8229dxWk/E+kKNtQ
bBfbn9DEZy6xB2fjVirHRi9ig9+jIuT1+CxPKt8BWYvBp2SwOnMA/Fhj4rlIIS8J
V8b7ui9+xAxLT5PMykRNgU+QRGkrbzbxgYXEWEXq45f1TrJZX71JI7DR6Wt30WO5
ihQ/1pvep7bwCkS6G6AydXIgjvCWKUS8GdQP4FDXRR43624W+B0U46s1bfxJL+1C
WG2OBWuOs91pGjqFTgAY+6IUURm6lfI4KDK3dFNxR2QzHh8aK/KwlHz1TqfXJGji
xWceg4N7omAClzEx/Xl8s+Ai0sXSDK4sisvGCP3U1sDsM9ZG/GCviP0OZX6XcdeK
jlsk+F1L0yRxCk7qJHt0HeCaYkKFBe/7U+D+fug9k1lhNGyZ9oy5Axw1IyPI4jQK
LcPljFmUnLT9MflzGQo98vPSib+8aGpcuzpjHaiYBokMWVvdFX4ktgtp9Wxl706l
l0AgEVtF76sILHh0J04CX69VgGv41jYFvqDfiwpuYGm8Bp6M4NmEFOna74MD9oSL
3ZBm0+IVPP55rcKqRvwM3Mdaw3OP3R03YW3HnqC5wusMqMvkhqahhw/RQRAya81J
S3FB963VZVpPWA8bqRkMihTuJ0/C1jzhuVFiYDQjtbEaeRV9gvZ2M7ClkC5FOO7h
D2n0eNxhHLFRRVTaTl/gsuxbEaVS/cbq9X9rNYXJ52bwR6RIvXMiHw/MlsPAv30J
NU1SJRrJgAzzcy5dUIsbiDcxuLRbYB32HlHS4cvPphhs3qwwYFVuYNJT2TmwKgXL
rZEuFKTLqt34eAm+k3MDmD6HnQNlGb20sMNogT0N850tpJnmkpH5WIOmnahfA0vj
NqG8V7rO6anzgaoyg/rOY90vKLue37S5ccmGw/po1KOOMNvhb23uiZpNuWct+bH/
+EOqqA5UNOffuzWXk2/MOYBgsrckFhjrxgrhMrgR62QSW38rEOcx9fmJcrquv9Vw
ab3oTv+ikubI8q/MnYebPSgCz+zJnkT51IQpiGzD7AoEFUpwSSXojfKg5AzA4r+W
+HhuZoXCxng1JPhHlZaR5BEFswOglV61XOJNErJRVfQZDCYwK2G0DeWAtevCTUp/
9c7J37YxWWa492DRgaPuaXdI6KGR/MM4NzpkOxi9P6z3YclT+vL6PVmjzAYD/lTp
dfGpQgukaR400yECh7IEpiYeCQwDSL5bL1uaa0qPlt+dInhpQV/dy22mRnar25Rw
sqTFU5d1UhRKKSRm16xcbfB2CCfo62/pWOzAMWUwB/ab7Kju8lDjGtGhuPzQOhCf
osKSmrVu3GEiokKxMlOzofcXUgsPZuIXPq2s3zsUwcQEP/elLQ1F0KCTBxEI3B3b
SMpl/6bJtwnS/UynAkPr/NFDD3xKY64GeqIaS3ASZAM/aW6k1diI5ra2PwIlXMt5
DVhQ//y26zs3LzrY4u6+t1U4QD1kN027LpVkQg71fLgU3wPqMaD1OyqRdaz0i2UP
HIg61pt7CwtdkoFp72DYOp8iuDUUnqLPFflXm7MPLg0a+BzHQfyHIqDLPYhCll3R
EBTmZ6w+KMwYjuphpa9ggZTKv5XIr2BeSx2W7EusZa5bgB+MBii/BF8/T+dyBx7U
5JcfpsCMG8bQJeksWzqiXkrrJBFBdq1+baMsq5u6o0KFOWJ/V1fQpwK4/8pZfOwp
rqGJIzh02ok8PZN/SMHySd55j8tIBAxtPnU8770984K/4Iob6fYGXlA+WJSGXrqk
Y+DQ+WNsOLye+FdkJSocvtnqParsIB+pBSS7vvheFvyFaAh2/Uh9ocdzOGevUsgk
MxP2rqXYc5v+UTlr3CL8Wfsj8GSWMLnogmvzVVCbfkyQtuV2+d9FbrdodikhIYzU
N5vWUu3Vd/N8buQkije2+NIUg8hhQq819eMI/usN3G862aynJp6A2IT73rpS5zj5
IlOvOsvS3+WV5JnNHLLiS+K962hb1rdV8LRAwkRJ+Pr9s7JHI1kLH24YcJ1LWUzv
97gpZgQ9NxQNx62RO1g5X4y2ZHzH3jUGmWch3gUTUG+gma9EH1ZNdi+G7xfQySae
LjaqNDGdtMlJAm/2Qt/EriZVllwwB7+PodtqTgYLtGJNtt3Hsx0bnzuhrZNLKRL2
pFuPbXvxSLqvaCnYCeFheBoJQ5kPRhY3ukKpQR+3/ygqQz2KhQ8w0WiUNOIIVidS
oClKU23iu8IO35hjLupwDg+GpiBP9oOg7WWdtCvdSU1UtHBlygMR3iLen/3DETY0
MBGtQqDNMdXR6q3p5YnjJ6lXTrRQzXl7fOMpAyR7qzn9X3AWqERMOuNC/1p5Rvcn
jdG8oVlOwv2o3TaaCvKLuqMHW4txUcY/iYkLTRUCYSTbGWV5knU1lZkEYCKubLoQ
44O7uxJtHwofSmXDCHx9kVt544P5AEJlAc9c/AwtfsRCiwV77SLoFltDGb7WnxPu
tFz3YDR586+g4Ncd2irZw6QZHvuZoM7Bxck+kKq7znza7W6MnTN09YnbiZgI7Azk
1af4hMuk9zrLawIVkqZJ6Y5glySeCAW2/3wLfHhQIuuDqcmK6F6lKIva0W4BOyJx
DICXxU5wwm4SW1UidfdbUsGi31hklvw6EN3NotdiOSRLlJ8p/G2IeZm0tsoGO6ro
uAHQL4fI4ybNgsC6SZSnvUysH1LQrI7JD6gY8oiGdfenbummecpMEQen90yiJcpZ
t7Zut7pLUqiIANDbJ2VBCMoZ4KiLwTAVto8m85YKv+HPZO2ZfIuTA2+3pNyQZew7
0mjKd4ATVc76l4h8oZpvPMa3xQwv7LPQe8zuAAjeqhhzXo0ND2h+9gaZc+VGMN9r
UEGj4Z1abas2ZQSEnJKwiiFoAaGsFpVDp/XGwmWgfGEd8FIv3XlbCvVvPZq2Ot4/
M8+aVbhp2qTv6BT8IJ4Z/uXjtaNICT4KLfg7p0gVG0HPuJG0H+TacLzEzAMM7w/b
XjL4VHPrTJ2fU+lSPAb41TebDURW5Y2V13XdUlCiVdpuONlpuxaSz6Vr9gGpHhAf
eRRica497HXlTLuyB/x1U53LY7v65JYfWCq7murKjVKrpU61wfFQIWbAdxZ4B/o9
maiZIVYSA7dqkTHpmOFqPDTtJZ/xApYFiIlme6s3NZsYLx8v0c/Gg3eKS8Eq5G2s
unHgVlbK8K1eUuf4Xt00awU5fMKXzMhwtv00nQ5JTSPiJ/j6EnAwh+29c+zJt294
bgJZZnoAEwB3zTaEne4ghgPrj4u7eh6MIJFY4gNPq7qcT+T1gzJ3wehwjjr9rLBg
hcvg8EgEb+oTlEL498vSfTiBsZpcQ+H9bKkT3vqG66H5sRt8sKeStMdYXeXJ+m+a
kSzx8o5TB05Yf3X9OyiraxXg7VKwOHpG5rGilfhWooMTU83jyDdxx4sYTQAcMmA9
KPGr4MlPrvPtkJOQqz3Eu08kD3rcB3DuyZnRSKRcstlOKetXYTkphXCtgMi/Zv/B
OvAH/CiBIo2AV+jsQ/dhwzhq4NcrpU67egJ8BuWIBEBl07FMLGClugrlEE66pNXk
60aGOjdGKZUo8ckDUBg05OOHXbX8tAgFe53rVaBQWNs0egl1+VljvqTEAWgxQ5FL
/q/5ctAwcPTAidKxChDit3JKbtH6S7HGiQPNfImVtWXh8zgrElKQEtbGnlubpqI8
iAF0D+Kh/rf0J2j3lZQKrBOD1ZhZnIHsBag2G/nuIK9NzA4cOrFthXry1oObLIEz
w6w4LmhyKILU4WvIiNuRAZ8Nj02EEc5z7gXhrwPD6aVLYgjxdOy3dg8mfSfcSrfP
1k3KTcNxJA/APvKYEW86y6V67UEQHZrTmg527NefMY4X4uQ4PTWYdOnDE0SwYBdy
nbo6Bg/dmSBbP/Idm744GYk9h1kmtjC+8+aRmcAHVlAablQq7T2zqwogppJoyr3+
F2M0XHejVmDIdZHROcboP202Y2omU8mBnFvpsl9NrofbMfbhVM7R3D0TeCBiDzT7
Rag/IdOCurtd+KDmWS1TQ6T+6tVUqLB93Ut/g2GbHli1CjwOcD1R93OC1gzFbaZN
CEOI83AscEi2qojDxZYoKMc7vP8rL9+bVfrdZYBRgGlepPZVBbnFHEbzW5TYxXEx
zJWNzKsQ0o38s0iUX6JPAga62icMwWE0jb6xPRinh753XztODUyYY8O+31exu1fp
HGB5gt4pzF4GH4fiTPNkHlhpyO4ShwwE8zAm4eh6/OGhtCrjJsKjB3MvKIR5kMI7
lNJbdY6LmpLXWxDeXxVoJUXmd4JEE5lqo2EMn9a2t/o6dL7pnml0OTt3yMX50QkJ
qGVLiznSJ+rvGLDb5YkPSwg5ppLg0M6fhaTVP8eYcytLTOWTeErO4Hf5ulc2CCM9
Zzjc61YxkfziVNAMS8xprgXpqMpHtBBXY6w9UlHq/z5HuqbdwrLc9YSXx/w+SrZ9
qZLj5yR2edxOANt6FwowX0HNSezoxIb11g8h69qnS4h7eLQdzx+BKkUmLhRnehU2
ce462kEXGjB1FCMJXLlGv+a385x88XcPDnjKEDBu+mnJ/cvHL1IYxoJHTHvpvAIb
0dAYTGiZGSP6CC1AJwW9efCDeOjPL7WrOd4XIQcSlPfs9eph1BuydR6TaKan3zwD
6gjja3MyhJnjnFhJ9StTqlN0qcQftN3rxIu58DdzAlJFgXO430osbFetJL46qXh1
Kjs5rpv1EJI8Kd5njxXzTkH/pQ8NmnTZzu9Tjj8syOB2O3wI49OX6dOA6K4+TCs7
06kRuUbRQWrFzN2QzXnMfPer1BNyet3/fYINZvxNSqVSQmG9TlJ2QenT2IwKobLX
ZdcgaJWBLLB4TgbJndt0XY/Pvaw7kLYVT2/6RXLbbdf2uHRRWd3+1dj+WiqGFyOd
QK7lp9IqK095QVBFom2TCnP8A7/aXYp3gNVvnbFfJaC0/pofiYCIgy0TNqKlrYIi
+7b1AsXX3WaoRGycmLShzrmy7dhfSMSAwma6sXepriGV+k3hBCiV5P9WYB7l7hT3
9zP/6NO/Pxl516EXvW4D/kcEV4dqoRCDaTGYn7/sxGkZ+o6VFgN6n8UMLh1xQa5K
+6tMf54Ei1ByvpsxqAwiLeisQZzS0By+g45WJ5cTXgmIcAanAW7Zo2L/4BEMejVw
htClESh5VzklJ2MtkJbWxHnGt6jHX4YLaikWBg1JCTvj6Cr83B+bwDIJ1n2YYl7J
CCl649beMcsG3uq5OzgV77U+1HSwisUHYN/7pzLdFTJYYJ+E19Jyn4gUbbsc/+DY
hoJju5TmSXe6XGpCJNNE0a/g4IYrMTtn5LBB3dAZSam0XwPq91rb7tLANnvEllyz
KJuszThzwXXMWb2pasEQBdxs6Yfq5/SW4FvzrBmmBv9ETiWu999jlEARQ8sIhiIG
jnr1BqE2XPUMNVDID9R519LRWQ9OovUjeNob519eKyI7bXnznTstX7MNRhQflyeg
Yz5w+q8MAW5ewgCFldyeWsuPF8ri4yGeGJ6AELlHjc3X2QI7SvCUkXNiMlK5xlJj
yvbu1FRybom29p9c3DcqSMvXA0Iry7a4CW+aS5Bl5c2AXR0R6Wo7fMf9gMbekUaX
P5x46hi9JHMiquRow1ZPBMow8swDAXGmEgXJDRrVJD4/j5ahQcaGlKhPr3OYeB5L
DQ1yLLQPdOgvy1Pbm1PYScB1K9J0UhBCMCHddX7vUnt7osIZy8ulQbxQbV7/iPYz
YkJG45tvncUqye8ZIEHjAb+RSmrYy6U+XyeKMqEKCe5tR3k+tv+YOjXSSJ5CbXJd
RcYUsrH0cmWk76+dxs5XCMb9HP7QTKAqZ+SD6nyms31XEPPUooT6SCFJooiIV0bi
uDRmRQCdSTBWI6K/KP5jywdH0KZ8KJD6MFXSVGQ2EXCnSKWX0XJ+YAcEMsOv37Cv
TgLZBPEaWtZKVfA7k8Q21XVtrBsgOC6LnsI/DJTcPpEoOUa2Kd/WQjC5r6Xj1XdM
rqrp+LbimeKnE86ug8vg9T1IT6iIAuW8SyGGlwTbNfG1cFGgQl3G3DSzEDPHZT3H
3PH+UojUR+r4nhtAvegAePKDmOpBufgPlcpZOc5Jh3nCLq9Xfg5tCvaN4tXKfECr
2PPCaz560FBzsK6JSLB1nlc3u4MGaTvnTezb42yw2RQ7b8RZhalNw/b7i2fkTEMn
N3VCLgOPd6oDILY7Q8myx7VtLqgzTRDUN3/mv3G8p5sCQx12430v5WXtHdzdOWUl
38LW2U7anxF3vcGioqF30RPKRFD+KAGIvmr70K7XCVkrtFY32xWRWBGShhKXp/Xy
ChfUvL5DBrahndeukqx/BKQf5Z3ogzhnqM3Fh1kG0OvslGlLUrEsRWPogSYj2FbU
7FJDxRkrD0kTx/IBj7LFe/D4RhnjBbmpsVnWltkdRheypsg6WlyJsdAnw6mHn3ET
RBjb+S0RjB3DgG2V5ofBolv2Tcdk3dj7S9ZHG0a2CX+KlhWVfAeQF+3SJW3cKoaj
Jd1jseTF5N51hzOS001a2mD2XToWKWb0ejvaTLhzaAf74dVLorzVqA+srI4Dhfyq
Uqy+4sNLXl+4ATMXQham1MllTy3cRvWLN25XNbbPvAoF/r0bgvbAPJbkBBycO2p9
59ImeS0MRGa2ldKF41Hj0eVLwDtg7wyBxanDtV1uvT1O2JR14NPwzYqwAH3tGleR
ZBGHGYchTWI4xLRZo+RUoeJRYO8wMB+EQMt5rEDv3BhnMqsiSlfCFRIvTUAFNFZE
g3pxMhJkGnitt10QSA+85uyvcKi4YA87GODH/xVOKNUhIoS7pfDmVRAkiz3o02vw
rnDkPuVplLet/i70wF7hKtgTLxQ9nWh+mNfqjZlqAr6oTY4sdS0F8x+6rF/NKTi4
6K5sKFTJTGxzThNmRyBaOH6FSFXMCBlllYr5BeOMPfz1OSZGFyhHTWVcKATg2Y1E
B41hYTIbqQmUlCtPxHUkiHoRGn1SdMJLsLlI9lJVuUKiplIvHzLN6YXUjSmhdAZY
Mh+hOBYUEX7oQ+34apele3J/bYjt2osblY0R5PxhIiFfQkvCANRg5axHCSO4pUkD
UYrjirCEXOdzZJ2dKWhIhwVBCepfuQVio+sFgHEVm4apWMzcllbJNDrRyo84Mfz0
iBmvhPfa1JP0+xTDO16F0MA1B3iinzqK44EQhhtWt9XE7WUEJ4nq2HMPoyUiTEXW
xM7qlTbQaxjKr1G9VOZRhG7DMIP6fBidnfROp93YKmDFUisCi+d0NWjhJH7sDceT
j/2bJ5zmlCtyVdOwf+rNrWTCGW5baiFv13UOVSHRoCXhEvcDCuXULvG71BFEjyKC
4/lw2EL/NS1dD/OUGOkrINTOCUcN4ktPlH4o930ePKoon88RL4zkWIKx9gLlYPfP
rX88FYYuO9OY74D1+5IfeXr/Q5r14nLrJUzpb3ZSkP2NU0YsCgNzkU4X1ssYCEYS
ZW+flmJDdiNcggwPaDrwIakltqH4s0OuDx7f7d6EJdgurGLcSzV7GSSFsxQS+clC
AEPPNw/v5H7e/WaJxiQuvfA+IK7e6ljMdMzI/tBi/ZD91QJ6f5JjKxC9835zmgAy
vATImcrpaAOXVA+yjLsQtvs0w74cmEqeHkIM4kUT3L0iC/3nOgdiOFNc+S7tQUAo
T6k2dl0JlpvoTfyp9e0vAP+2hf32bAS9W0ItMD4ijS4fo30CliAGiF+2thjIsJG6
4di9Vp9kFdTZWfbPc419bKp/y50EydP5XrSUJpU04swECwe5K5F/bC4bBdX5MjDw
hUWLS+Eib8vCSpm+qtivqqVMrJtipXBvM+UTlIQr3vX2ueXy9WbYmk7qwFDjFDK5
1ZXIjTbWuQ/JvSLczIs7dSjGOiSmhnZAFXlIJf1eze8guIh+s5PCA5PyVI/+O1UG
Ut5XLuZe5ea9ExWZOU7jKCYy1FKKjoXE2PHWeppoSyEF5XBKlDeyZYSKLFLsKdbF
1+mFN613UeRjKiQhh7ByqU4RhjSQkz5F/G5Q1fahsBEvJ4T3ODx2TSlx9Z6ylRkA
R5wu2CmKdWJlxIb+KbyzJKQi3QGXpNlrwru3dCPUu3UCaItT+EJ5E6JNgzukm8Sl
pM+I7eMXjg+txnoxzr5ZX02pxYwQga+Ud6pzQ6pm8kFs4x9/niMK66DaDKyOrbmN
OzIhTy/IKrGdGtpj4t5lJT9H532TQTeU9IvuIqf7GfLoWSWT5RTt8oNEryzY8vGE
cujS7cgv4rpKjEVRWN11YQ5lNS8pvMI1qTyhXhTBfXezSnlsi6WtuUY9E8ZGMafL
kOCvmV5Se3X/ZQzqbu1N2b3EpO7m9N39SC9QtgMicuX5cMUtgJApQFLRb4SzmfgJ
NRlFoEkZ/oqI8bDFmmkBzVJ8mfqTDBrk81tKEfsRvZ2kJWv3Mazv0eoJOWS5e6ix
SpBRmm8VLMwCeZ1dnEjoH+CFByccGjvxRqbLXtGim8jpL5oYaFCaLkthSbNL69vV
duhSW+8uDfu2300+C6nZ2ECkAg7DkfNMU7WBnKejIBv+gFsIVFCd4ZpDLj7gz1Md
8PTFmnPeCZiu4xmPnOQe8TV82/DoVhuQFM7Tzsnvo4n9IJOmVu6Ezg4ePR3boy+b
iD+F7xtzSnWImT1GRhjy8nokQkUcDNF/ZQ2Zy/nyJcYM+7oFZhZgPTmNf8ZVW9B1
DaCBMSF3UC80Ws3HToCovCmd7ddHb0Vzdkb9ebdqnvNB/qA1Hbv7bm9bjw2JaA/S
xcXkkvg06gEPB1FxT2bggm9h6EooCszITTWBdSMA+ZXzgubl82fmKx49dmu2wSUF
JeTUKebL8N172ntn4NiRfNb+43RU7wXAKsJwL9qhMrCrajFSt3HVPvI6HPJd0SF1
c3xlW8jkSxj2TFhLpXips/XL0ijtawIoThdFGCY60s3rtCz1qX56ZwmOSNIc/B0A
HKUSdnMLpqKo4YoKCuG/hRwF7IJpb98uFlANmlf/qUPkJlrL5A/ngMh7U8i0tKrg
gxkBLn3tPMl3R8zTRop0VMOZXDmcG2PtNcI/rK4XI5SwgtjJYA6K2pMOqeOxaIcx
rSb5hGTVM05Cz/1+0O6bjhcgIFeZhHJ1OTjeBq08a2ktZszj2f1GBqVRN2NDCB36
0wAT5Dct/D01uLL6YU9w0yAAmOyJtlv9V9N+3mZtdCXFObp891nfzRkVvgR6OZAM
M/BRg+xHaOBk9OF64jqA6gdXhLuauOpDYIO1ATMPQRLCUx4ir8pwCcfU8qDnftFg
MJxt74nLX0z1HXvQ6/sejCZ3TKptdwmAX5ge3R8QdQ24MNHvnCIiZhvo+KhX37/c
2sNh5tm7x/8eax7i+o2UqgVau7wm+ad1vBkrkA/IdGHYJYfE7RraFPfx+eTEaS47
8dLxZrqDIEiy5jNSOM+zmxyFGAb1NRjqVm7SlTqQRiu3ElXYpv4YM/r47y+QG034
lRi18inQEI1mBeEFdO805BkQZCf09Vk9mihpCCyuAWjkv1bzeJLPiBwbqb2ELKfb
cgxzpqvO1q2zbbN2bfm86xhE2CHaeEtmvjvIFfD42IwXeyT9i8sLP++6Y8nMBdfI
ghHn09fMU13rlXLwl+CL4SLPss31Yt6KSE4/Rch/XdEm9yAxsIB1WkgiTJoaHA8l
Y94DUgzlZc0kxNA7YiE9tcLdj13fvr/YteGmK1pFQp9Rj7yWd9exKC5D3EWCY15z
m2bKUMIMGUVvFxsvlqEHMGZKbSEOuVzUDMqRwcoYZXHO1bv/OgJmXKgLmD0jFhZU
LD3vBla8CB6aLomenHGdv8/UBpCEsFnMj2GGnk114uP+SUZ8Rbu8tbxGD4dTXAqm
QBeAjGqon5VzMjo/nk3ceOvyaTrmFuSuk7tLOS3SSW5bgMas5n7a+j0EPw1Y0FOM
jMh1eiqwIhq3NfZbwtygJF0Z2MS0+g9fVvI+ADQcf94jME3T/BsiES8b+Au9jwmr
kF0WRG9Oy6yIxOIvJaIhED2MXEb9+TLyHb1Ie7oPqdDfctdw3mx2m38zG+RN6n2r
pjY9NKZOOjJeWo0umHoBT9WAnY/cmS8oP1j3f3tqvhLDV61Jl1C3Y0fxixftF8Fw
zeaHARYIEqc/LCB8MSDo9WgHoTS4ehGFIAm7xiUX6iZ6YYv0R10w9/n5IDg7evqR
/NqjP0JFESouWDQKWu0Rh/Yb8bF3I07RUNJNO3G+nYY9RG7NrG03pEIIGs6FqAq9
OWaEg/tivJIHPanhJgueCPOksWJzeyKbBlYLmSIEwxFgL/eVlIZNek2QXYYEqxVC
lsbFIyS7oUNRoC4SBsAKKIGN1CBylu9iXZd/wPNnkjx3XugDNyRNZI623J+gcU3i
htAJaBIAxkFmp6jfxg4atGionLB+DWpoemQ+bx0kiNxvewYft9Bhsv/pnnBkkLxf
865P1tf2Bi4OWX7k4dBzAEQL3nKb6DT6liuWQONkMLkoGCQjNWEtaHelYpwc3JiE
LkiEpYMUJZkbBRlyOTZ+a9kzCYgJ1jFzSsx4nXFspEfRTnOOQgvtk9qGIf86dVbX
YbM83/kIMZEU2e1ScR0TD1PjRXxeVru9eipb0htl/fnkYHROQtXLJcuSAUzuEu9V
Vy65z/odSWezl+/ISho9f4uDdzz/swRxOmfdx4Lnu3RzZfmuAE9yClyffD6fluq8
9GjZ+Y98MG4/HBAlEMSASPCczqXNtw/xUWbzZ/Tsd03lPTX/kLewATn/bf1JXTrJ
CDtPpV1aPxkfbliVteO/AK55MfJ9680v8p5t64aVTGACXL9ma2LTKdowZuNFLZ2Y
1APBJ22nVv7zOpXkZQ729BXXub1d4gp0+Fl/te2+4P/6/hU7iWaeovjDj3dF+wYy
TmBQCo7sq3v+haqclYHLH+Kk9uGYyiYC85fIPdxTFD5NC3AxMDs3cKZx8onpRotg
+zoK1KSO+KH0B6RXsV63aK+rwlNA7YSkJRach2vhSRQI9CphJ18o2RP99Nlgm9qW
ckM7DX2BObQWTEPuC9M6MkNBsYawTe7FV97KETY9NJnh6G+GuW9L0MI3OMg6aswI
H9ga2S4h8d3bXxwA1bhnnjlgTscc4pypZ4I5rvud+Ys1noPOPvAt0GCXu1PgIil3
yRvh3MpGvb8SYGlKWog+2byhgixImLGrf92JBFuwOyVSP8sJY7YfORfw1OHSjwor
/d39IoAckAbB7wFdnTxur+4IUT8ZU0D9OzM6lNtSKQnu1PhindmbvBAcXGjhcKUV
5n4d1AM5LQLKtAQGHe9Gx+D2yRTnYmqTq5W28k1fcw2UqG/Iq1sndqCoa0bzq0jw
8OaEgysygBo6vavHRrdq4apE6v9ld0K6RMfwGIdMbDUNzhcNrNJjAWwM/0b6WtK1
suvxuI3f/YUwyetenEIrtdYFtfo8qfp0cpFfWi8S0DrLssjZ1eKsvbrEM8IYOmP2
RzQ7AZhFikdrZ8/gmwa0vz+MyCsUo+6i2HnkWgaTj/5oq63cp97DMiuYcIJgYJ7b
9rxC522ypCZ/OUX+ZiSDj0j9a9PjyGYRIIge2mo4zy+WgiV4YvnxRP7GqMgbIcfR
LGgOHV1egkJryMtxYGkE9p3wS9DNv2q9q+wCL+/J8+sxiCmY8QCFSIs5d1mDI0EL
HCdYm97Y/ams3XyiFcLCTTrzULd+sjNvPs985upOM10XYSJtJhKOzSpaLHGeMxKR
85SZeCumjdAvDE6bEm8hFZpzbMyDQCeih1G80JXdWzw6lRPvOhAspxiZmDFF7nKB
YLc0rUAXGp4wkF3/zyFacSZ3BfucwWez7agU1zPxDVesP5wXzmQWuegG8AVuoWKn
Mw+oLE3F32njuhqKAZ8dhDN+wN3FXmxQAdOe9WcrAv4P2VN1J48kifAnYruh8lSG
PYgW7rP1G5wH1QJxaYD0WZoQ9EOq5GDeLEpq9oKiLw16JVqrxBeSGbEYqr5rhiIZ
oWlIexuS9nnuIi7ElFeC0cqAz2gf13yQJCFXk4/18hxTIWEhZnvSao6sc9gaAJPK
PpWOnbG7BufP3Em/lEG6Tx+ewk3b6xUOY0XcLliwawzPCaQa4e/DARct8oCO+ucC
EfibijUkXTVrtII3YpYYZbU9YPtqn+qb51eIhxnvuQaftJZ9EkeYVAMnLhhUh2kR
vPPrSusGwlFxlqYP+xE8J4BRoLSxCTet6QLjtK73fq7tP+FSWpZS7AmRfSVROfsI
e/enmjEbGUUHe3RWB/KXUHfRXfWN/me743NFzWArScdqgcjM5zQ3fzIfDGyFxwMD
X33RKt5gfpqJAN7MXvCudi24cBwjkwl5CxDAICFkVAjEXZDtnrBSXOR1OW3MutO+
pF1/4Yjv0jYPcZtm5/BKyUlP3qLMxZwU4Nomw6KX+14XbmUQpsmg4RGC3tZCvaR9
GCAWC4JtRYGJsloFnUnpoQ+AEeP+W7hqWiUrtn1rXxJKhEd8CWsnm0RZrHT7U4Zk
fLyJHttxA+O9ZPEVAbrFOKxjxVECCcUKNOHDII4Ho5LcT/RXiZUJzBKw9RWe0MLd
4s29g2jc/EpTKDUCgJIngS6+sHn6OVNs8u7TtTSEcbYwCNRvQHOAeuIoiQUb4jqw
sxIKt4ajV+YBA81fyDwGQ4Uv/ppIBYGVl4ty+BtVoca2QJ5Io0y1YH5oAILpW6+W
ZqX9i0sh0EbCgwn+N9QooXeF418FZVkL4F29IAYQdIeLymPcABHfkEVYtG0Vy65y
2WfkE1bZscdvWkHWfboCg7ouw2YXnC09uhpZBcradmX+Ho9+J4PGFiJV09WsGz4J
gKkb0CNg4v10BrQDlInpaF8//9j1GwhwKlmK55EfOERF4vtJrJygy9cKtQOQp2SL
KZpkBbFouVOuxjL7y0wudWDWEC1sJGOFf9i5mclr2INnS4tLoj9hp+vGjAE0YFq2
Qki+KVyDcE0BKwMUGTh/mj0gHrmPRz6f39+FAjst+IQqobuo7lCe8wK/QcO06QBC
FwYUdCdZTG4L5L5Kt35NAbQ9E55GO1/yQuPVnncONfPRisvTSiJpiNEm3263Shq7
0V109VoHYhx45zSdlPO+236o5070ZVArt0TU2mhH3z8oB7SuTLoqY806HbEi7hRv
PVxU4709WpGuZQ98b8FXQI7Ds6/ZIcNbbMxxwhTvrkvJEl9gili3UnlMAJDrJ5bm
N7YJRyihWS50FDkR+Hpzg765akbtMhFK4LHyApKLE3sA9N9EVxFbxiVQNRztHs7K
eZBSN8ovETX0ZLSJ/5oiRueprVnnydxkvzQ9a+NasDwFZYfcKtI/izPUzxKxDrIp
k83NV7o60JwqG2YKhXs+G7c7ckvby/tWllGrMsVbQKxclNVKMzI3113ZCyHdDN//
NCDXc85RyMnZh5hC6q5IhqqVeUj9yfvIsJOZ7IOCZwGxcnniHs5NPEuXlCDOANDd
34kN0NbvLbboYNK/cH64ap/FACml0bpkA++ONJqU/1dJpHGmCEQSN7rlvCO190cv
UyivjScSSrASDOlW0bzeJnDA3RLD6oZAOfyQ0yaSjz1W1XMr0g7+pbIpzF+X3XL0
woyM/7Baxm3u/M6GZrQIn/xyvIljLvLwvr9xLo87xhttuWsysrQZsoP0ykdce41K
htv1NUJ6oV1oqh19nG/b4i8g/CZUT98JaNwVkjmSsL97h4fVwtS93UHNrJV1y0qq
5l8RN5rYgb/S5Mbw260BQU9lpf89S6DO46Lak9rO0lMXlkvgjWTkpvrVaxOxX8Ro
4obi5Ay49OBu+up0m0wMlHf+WoTcugbNWT4mlR+Wb3CW83ZbXjIOkspFD5LKvcXd
MSqi59mfUnMDM6gvItef7+oHlXEd3iNTtSOhQBcXHP1lF2TNaLVbrtiSP7KOOKRy
VzKC4C0ZpOKpWqid03+JlVoZiDna4cpF0Z/VxXq5JjMeJ2eeEp56kDABwadJqV8O
h8AWFRSzmH5eeIhxKY6aGtRrmz+ASdNLQ+PSaHr9/KXdMwcXzDkxCm4DKL5eOtN4
Nt8UjMSsc8qOB2zTQ0kvsGovpFpHDtc4wWefqrulBQzjAi0lD1ccW/XUDZ4lQX0s
y+mvjm7BMXBuivMXbnjz4j4nklyMjXJ/eCBXkYo/SnCFLpRT395cG9pA0xW8wd8O
hV53dHNV7yHf6M2ugv2znNHzjEYtbJHezPj9H36G/06BOmEhq4xqnf9V7QOPtV/n
FgXKg+/QYcZ+9c4gpsFWI5b7ZnxsYOFSALqooNCpvPDduF9keFeaXNngsBNMgUl9
Z7lpi7DLRcQrHsxYYEScevu4UTi111zz+OH+VMlREJOCOXA7UMKBg7gYVHVGcbeK
bcqqfoiyZAqxNl5q2wodzdbTp6yLa9958ybjzz9mhV5vaqbmwM8T5W7+UigJvJDV
+KJPbzFWBSIYmGyIyDV0GraWOm6BTOOjQ7vMfoXQqU/nLX1yGntxYkPXaaQXWA4w
4D36LsrJYXFm6ITnj/R5i/IeBCpcChjUlvao8QPQgO+kx/Xqe1h4jPokp8BninG+
SZ8+xLKFZaM4NT1qZqYjVoJGhEJGzYaJffMFqN4CiNL9l/UfCIXG6PQxP/fT62NR
WHpEuYG2kWykW05d+ZkgLI4hkNZHkk4CizAtpp0fVXxt3H/NxJ9tZ55QW89m8G+1
fJloodLbjgpqyS6lDL/ruZwXbc6A9eW/0siRA3qd+0piNFalXcWTBDQM5m/3qnpn
FTpoFtCU12+mqzTdKcUGial/F/iFJwf//nim1l0SAnaO24VkQ8r8d9VYus4McKL3
ndK29jQItEXMGRvqbcO2VXs2Yk66qERD8+gzFMnBcg6flqa/RTc45rjQXwxq162Z
n3t6p87tTCqocg+N3W590e6FugVD/pMtMR85Y2T4RYJROWy816wtsznijnQIIq1b
92ZUjE9Lf2Hf2coHybjRVCUS4+h4Xv5e06nzf1pS14WbzW9ju4Oh+FyTJ1+nfGAA
9ucrnxQtoblOFtp2p2zVFH01KtTx8k7zc/QFPUe8x17Oo4hrCa7tGwAw+tixQHLn
qsdXhPp68dxiA9na4LBkGF++7F7pK6NUXhrQitpy8mpq1B5pjTuwlTz+uLAD+/ms
+oz2smfEdLbZVGwyIXUWmmt073/hMqy9SXTv+or8hWVbVcW6HbSW7Sgbpi+jcVtm
7G/kG9Fe1ozmL4OIV0kAUAZg5Qn/bUNskjiWW/0j8xSABBdsIY7i31ReblxieNFd
+Rc3O+6ZWOKyOQYSokhfzKbJlZa06tPS44Yp96JbodmoD1TGLFjJ0dO8/61HmVWz
GsNpX3Xzb/MS0A51UvJLoyT41C8Ejrhi6vIBQ/8O/yB+JVEPpJC1cdfgUjg/5acA
StTFAVtv43kgdGB2HynDeR46hjebRzjvYjC2Lmb05Zqiqt99d45yN+BdiMCwShat
RioGMACSLXOeYE4YX5jW/FRhdY0CZeE3sbTC6vXf67akUlIPKmz8hLb9RT+AGpGG
hQlnXU3wE0aiAR68Q8NQXTalqKBPnGDRvN+NN2vTotnt5SYhmJP0XSJu5T8IyU6a
s0cS9Jq/sohdkUCylzfSZeG2yPjZMtcpWztbLkMWHQJ86b9XdydNtVYEXEb7iEZ5
No6hBRHrno7ehGiBMxlcgQZmM1o7QXekXnfpgAI8Ajzmc4PkqgPpxfz3/FcxitaV
qRMJszDYKgxnssna6wNwhASDdSqfBM0L0ALNcRZ0OVnGQfxh9002GNAm1nZT41RS
epKm9gl4rVdLvMK9qfoap769MCDw1eIHZx+dOJ4ayJPMTeex81eBwx7HnZd60Jz2
nY+KxY45XdDEWKo/XPYuTpoL/KGgN1uMPatlmX9UJHEq1ELKrmzBi2rs0rNaqhvR
lyedrYRif7ZiN0JBAGyoGtx8iYTzY/X8w2fAnIeGy0VQmRael8jAUeiR3vAEkyTA
OSMjaHK9I4r3qpMWWce3qf/G1529DXaDhpGj56QPeW6WBP6Cl/03RDYExojF7SEo
K5N5T+pBMmi/8/t2kLneAtyf699qjABNGRhNfjxwRqBf5PVYRyyPogZIoxaqsbcN
01/5uvOPlrnqOe5CvNyJuOXaiHhV6WPvKpZMMwdvUhku8Vuz0/vQDgUb+D45D8gs
E3JYN1fhstxFpxsHRG9nfbdygrQbnrMufd6OHV0VEZOM05xxqYIxAjqup1lRUPmg
sErqRhO2wFIaufTjRAmZ9fbJRHnM0mJ9FxnF+oqCQjp7LAlpT038J7C18Wv98Q+z
LcduAONkHqRoEc8AuYpgxuBS0onnS5MbW+X7YkyMMlWpMEMuEcCRF24Z9DT0ZEnh
cOHTeCUIZNSIPQ9tjhOTkosQBChbaHYQHiul7ZqLzlnNYiPxa7lMXg9/mTRhi49O
GgrKVVHHQIrX3G29RCF2OsgnIJEvgqTa6ZS7hfgtJnbNg/6zUgum0wugFmOxjxgk
Pl9d4x61MhTRG3bclxylTYZ10lF18fCY7D/VeO741ywvt3za9av5bc+XsLl8BOci
En9mmmrD29NIZ0/DdAXrwE3wfWLdjQM20v6jRcMPlS3r6rlEdDpQJD+g/ZzVnmaO
X+iLkPYjfxUP0YbDzeRSiG3ClvCR+4ebdCf4kPiO2jIK4+0Y7ZC4XmSU6BE/p/3d
qeZxm2Ko7ecrRmPIkacfMFR4A/h1A59Xi84uvjPjRKp+rWhrCbhPhRUyVmv+Xmji
82GDsz073rzByzuf74nh+4HFNskpuumdrx+tY4SpMeC0UPGNhxfXh5768O+bWK2e
z2Ubls1a8H7PtDCOMwSEdnUwb6AzM0+dmAW1k5rqWLtKihxavuDnX+NNLqVI94gh
XgBP0vonWTtt8Tcpf7jte1oGTRbbBoLF+Wm2VhYrCHCax9HBuFRCFDwopa0u1rvz
i0tw0opnmyrnjME/uwYVJ4ZQyEH9eL7WaoXOvTiuv0aeo5fGVUk0pszZKIr+5VTq
7Ht16dJJICvkgKS6q4LeLi9UMvRu+iYvin8XFF5FKr2g/5Jf5iphgzqr310UF5Ti
41YdQOt4ZYR6zNQWZTXEGYULbHX0cCVkKhAP4nfDZlRbGMR0nYyZgcuWkNJ71c5/
mp2t6ILoYjQw7CEZgx3mhibNc5GANRXkdKoxieXyyx6xm423Kj41FWyUnBvHttSg
kqVc5F8UB/J87CdII1nskR+AZQnBQSxvXYVsalpT1xo4Znrv9e57vlTP/wg20fgG
GslWgWO7s0DUYZILYHJamge/s4tcTQtuB1gGdiSUL4zw3eYYoIu2p4db+TCKy9E4
OiHcSGOg8aiHs9gNfYlJ7omHO8p3nE9YI5xM2Vyl4DaR3zeYRDFckkAYHNRf2Er1
G2txb+/NjDgper8F8nZxU7M2qsurtd2J9aqe8devQAmIPOKIe9IutD0IekXmSpFB
5UCac9w4zbDxlm6yzUNC9eA8Dr3MeioyQeT0Nkt2kMTklrCw6X6feqk1ZyXI2Xio
nIbUn5HTQ2goZknSLP0V3/AAefgANg2Nzt+v6jLoxPreJMG2gvoyXm1nPc9BRZyV
iHG1JQvVn+vtZ+Z1MBe4pclFvtNhkZzdLaSHvoozFFyBb9djKE5/U8AG7pdwxGwN
PJiS1gOdOEUzoHOzznV90+YFKWhOepMLJ+tFD4mAEDd0v8rMjVtFapa5x5Sig2ak
VxaNVsVFKTDC5lwAB/AKpQOu8BhQaLgn5dsxTvQs5VQmT9unZApwTixbr/Tx03hM
ActDvZB1RjuqSeoHXGOLq/qhpSVgc/tIemO0eLLZkvGOStWDbCyQJ6QOrW5bCCs0
VT2d2tfYjQp74Rr7Q+Zlh5afU8jbpRQCTJmJ9FFzYf5rjmOiqIX6vi6jZMFZRGnn
KApReHOmp9peIFDJ1umg4csLOk3kvWUJdI+/J53GSb4XOZlI2sZOjUvZqGOhoav0
byvLMU2tc/8uKknS7azQfYtvjWJAkbMiyHHlpUltYRgqOlWEEloFThp5hbsZaN5Z
2tp8QfGkL0CciKis7QpZmHqhWuCmEtdLLXl6lSZWSjiKw5zRd2wAaNKb0tF/0hyE
KEQ6Kt94+qf1/wdgLl5M9h5btRPjz+fW4IQi8VoU1RlB+RgcOsYByLRpGIJzUElB
Ceu5W9QPy/OU7qXduAGgKILVuJLkiUF8uW4XiE89BZwB5dYDUCOSGmVCZggxWrn3
zBUKYtcr5tdKfDJIvGOY/AHj8qApgw5THEkAdTvKydfxUXLeiL8Co4OSMxeFJUiG
ypv81ulc6tyntKEQVJsguqziOeuZPmVwT1qUcCVw2f6MnRxGic1hDdKE19AGrGss
w22Vr/4XpZVWyx0/JGlkPpkg9GfL6EltlZ12LGSdrRC+yz5dPknR1Zmq9lMVcQvC
IeetiXx1Z2LPf6/EqO/w8GyEqaiaw76MTZXvhoBUobUA/xKJxbNwplSZsQ/vKhiS
wYmhV5xlSu4XJ1mdYHjtnqRqWzZN3VtLK4+2YiJCb7JOO7P3q1LfNN1xy2eq9y2H
uxXdSAefnBVDNiApfMmsc//nhKD17/w/zMbRq5Nws5bv6Yc9RIAsn6ACDDPVzZU8
Lx9oudgcgFj8e3TqGKbebGyO5BwXqL29KewnXTH+kh1rLoWGJVLHGqBeKZtvcDKR
RkYKbMeckwlVoUOD+MTimod2C53b3uxYzf9h4HoG6/pdVNJhsS3EDC7lRUeXVYtg
hUfoB0ZW/0cPhafoRz0Ftjx7dytxAtMgIb8wi9uNBxLHvQNplvz0AckLnx+nU01/
EdBIkeXCXYakqVNn78A9JKcYFXVbOwjHV/MVjcrrGgFMgtCQzEdkvqKNbIe0bL/J
4THhn7e0n6F56FSRMFKzDRPshHdKdBkRqiD/3oHQLviXI0V3z8DsaYiHJbZouCJo
8D8JTTpfx+qmBENkDEH3Z/ODm3STlStFKNvNzQvFMWOEc/DCQ/MZ3fMsA9S4vqmb
2RsLVRwIAkOClg3mXPux9awJQstxWLDq7YCL7sFO7BqbFppkZkGjlA/nTdm28bjz
9RTMUvhTCk2wTGuH7FaSUGD287EPibMSRL6vDG7NRpCPFLr7WL2lbE9hHqNfiP4V
DKsbKYHLHtGwoCD1AOIMv7L7+u95lf1dqTKI8VrJTHjYwPOi8p5wEkjr6/4/AoFP
vNmoyRpnHSf/ZMra7z/0Ad0kQ/R1Z37m29xw0gz10wCXHXloTp1ydYrivAHAj7Ry
dTdQpZ8/yZOnWbzmJkU7+LnWlDS1L3aT+VYqKryhLlyFLd13m++Oxd3e6EDE+WQT
460cfWd99Aix8lWGXrI47b4L8ahWs/icJOMqZNFV1vZ81v5ZJChnuxQIzcQWnZUh
RRTPBnIizxaq7BuPeGiJcqDvCb8X3CoPaO9QBly2t4JXdgf7H/p2ybzmDfB4Li5r
QTayYOsLaq4ktGjy2baNfEvBR9wozgHSvxJrXLJdzDnHAQ2Fel9T+tn+0RVlJVK2
uJzMvqX/d9d1VYETrOx04QiVPrSpZ8EFY1Vm0uK96gK91DPC7FdvXGrGrUMsiCpi
efXc4gLVxdt9OUmf2rp4VVF/wamHf3jDTcVW57Wq7Geyl8ucJcOpx76mEkPUqWGl
ypnhlp3dRG6fHiExP6Yu7nrwi4LwJj3iBCViEz7BynXc0ZQWxTmuArNH8EHSUi2a
EFre6CmIjYfDyYqWp2PvigqkltDwisBY0R0g2C28OrTOGo86H9AlUOc4QTSvZof6
927Olp3298LJQrRFfyNssFxd3mRml6T3febxyObgNKzkM94tc5MRHwX+9iLllZAI
uUu/NVjsZrhjYngzKHB0wGRRsgXPMaXdillCS807hCn0gqnWpOD4TbB+/PrOWrNw
1PWcXpaU1xH4822ezC42kAHkC1GY7nlzRwT/zvpcbMcS/rKlzecqiu5V1ltxV3wz
uaY87x8iSw/dwfT2tye5J7/MpfLntG9IzlUGzNdBpCNVTyOGr0VWyxS6CbHdVWW0
bqHnIZYI/U1E19grMwgQdn4q9v7U2bYvon0NbHPdBAmb8FQpBvyoAnCY1ZI2NCAw
5qOZyoacSOMea1NPaYnYmrZCC8ZuIO9S79XgJTEZgNzFKbUEsYFGB2EtXbQyPD4Y
Qww+S86BeJcSqZnsImqBcPy0tQRUtDIlOjb/eLi6//L3oFvYCv9jlNkwgQRSeMPK
5Cu/tXyKhbXBifp2izVnXzgoAlChEI+nso1BtsWft+BIeYY3zxAxWTaIJPhQ9SWt
ovw7ISYVemU/UvhwrYB2UB0Zf3NkkiBvNgh+p7qiGQoGOOQ9YnXqceW6I9VcbAZ5
znLOIfjnQX1mqpQAacFtasc8+4cn9rqP2I3K95Dl3BiOZrMmKmrHZbdXWQq7bwa+
dDQyek6IS912GMjHGuL4fnLcaa0ycHO198/uMXb5wYCIfBMG0ystxLHr436cFZv8
Sdf9nQ+FsX6sEiBqW4qambT0znIa1ZFAiyGu+pCXXYmjYuG3tRMNe2d7fguVfCLb
HNP/kHi6zEnfGPkmsWo3Tzk1h80wGjk0FXnv9XNoX9WSZf4d6CCZJ6UUACWhtQQA
BIYCe+4MjV4uKDKqXMFTq708eQg7UlH099AXsGBw+NeQ40Dcu+hdlFQDQf8LrKDQ
7fV/0ybc38tqZYbrzKwDQhVT/jbNKhct6phfrEFIId7fAxrH5LX+iwgkowDA/1cZ
nO8nb2GMI/Lxy0M8pQDGfItWTYhS1x3Zj18RIVm0U3cJZkftNcXdh65d4POyPipW
ovOsymGY55ejP0CJVO9ji5TGN3RivtbV7Ajaq65h3u/Fb+2iRE2YoSuPZkKqOtet
TFe2Z8e3K1Z/KOU/ClqEJXZ1qxDs6Kln/9EaA6BGJ2nbmSMj2RdOf7W11hluZ+k1
H2gVECpcyOgpu/yrMlRHvzUjX4j+PV617Z7e1Ol3uau/9G/Iz/t/MRnyFtAVFzKG
wr4uFu06IPOAnpfsFPr4aavr7yMPByoIE+SCHrngPioLR3w2y8kNYMByD3XdrKm9
8R/bsgX+5bLDcnp9DkEtnCAQZGM9QKza6mRalI8mYOkLFmlZ6c3sdXDDHs8eg9iN
7YHTdQ7tJwev3tbFnx4asDK375/PsNvY0/8BfIL+2WcPx2NTQUEeGH0eMqWe3poP
VnSlDPBWBWrvdzhx6S2XTSpdzWWAx4JRNLoZsYTyQ3RZW+SVWqzRvUk8y0xJpiF3
/p7S3agyPfPpJeVZQh8zUcq50BifImxNqV3tOcRDSG9iQl//RvsDa/wFB29PU/I0
n0aJ8HZiSoYfpic6nMV4id7byA8G/Q00tFrDqaircU3j0M0Dz+INTUDiI5CoB55G
Z4JhjEVhfDB9cYCv1x0jEpJMOlFYMKfWwsPTRdwhjTDdr3NhrNXti3q33Ey3DdFc
IyJZ7vtf6O6ydCuUpaE4ghkNscBID+MvbIzcBIbIOGyNKpUIdEweVgAQguMwJUsz
Qxev73ZKQ81fOPW0ivMm9b36K7Szn1Q64k1PN9U3wmUi37+Yu1ovkt2gq8PXwog0
Jrd5JwT7VyCNleXBokS/+UmxW5V9tcIH4ASha8ftzF/xJzCgTzYmgoeKXbIbqCd/
ZZWmthpPcJ0E6u25Prut/s9ZNXaJNWPF0BM0gicp+s9kfL2T3iDCxbX0Fk5+5OeG
W9YEp/cWxuKbjhM5kIZ3hKWd6pPt6m7CwISdFNi7XSgSgbFhxUIMSKee68vZTDW3
fIW8JL5AAcwK1y1OuRnPNhgKiOs5koN+/85NkXb/n2AuhzH6ucioM/OqG3pxqYHo
vemBYgAoojR89ltHEMCRAn47xY6AoDenz9HlmQ90B4/6cbZlXXVI23RtsPnr+INr
weOQRKQWp1onE8wBJLArwy4CGTWtAhozVK4TiIvzdDT/sszY/HYjypaM39lWONcM
cRg/fg1waiyW1ynkTEryJFU9gPfUWlL+XG9SWvSDui3kUCeMjxBNSI/n80zNp1QC
pe1qExZ0C3rfronql0UcrcobPhQM1X1ODHtpO0CnYX8rcvXapVNNYN0UNChAin69
RPGuBn0HVUfsBmgWDsGaBX9sOVyHCtCEA9FlbhD67n+JPp7AMibI2/MPpH2ikKXs
+3oJdUXd7+JhlPqThsJ+bGIuuRKmCFyUGcvxzZ6x6bQrlg163s4znGlBagiZiw6g
7Zc6UBFhOmIhp5HsvmC6zNeShMthOpv9KsmxbC5C+UKeMGC0D2ZCeGpHg+5Mw0ML
qBIIgQAfKE/0RNYOhohrGd3QJ8grRhcj028Pi9UoLgvqBkwUp7s0czlC6jZMd5DL
SPQ56lQTJRpbIpnLr/0XAnBwR7GHKXjWglywOyF2mnr2n9C3WlueNlql55c19/HX
TEkSOMT2dxv9efaqGNA5rTfdBsEA3zEiZ8j8F42ZZgddCgTbIxuGU/+WdJJ2lxeV
PSvWHcSGZ2nAJktH8dV8QrMRzcRAr2tI1Qp5EbU+duLGhSbjWUWckerdubh+6yLz
089yFJk+9dW2pwWJS1H4b/rJ0Idhz55Zaq3onjNfi8Z+tWXu5FAWddb1i3fPRH7N
c5FVHh+/zoH1uGc76vzYX3fcU8m95GN8XW41ty9rA95TDWztORNIVCRCbdkYzGiM
2rK15DPxgYwgDGQpNYdWZriVE8A8uZId+yKNl5I86xKFQ/nRuj0kIms0Spm1vf9l
eReFijIQ+3jRuG17rtVMrnScN23xCM7Adzojdn1PPguJdSiBpU15JlK9RId/hynI
1q4SCh5yE4g0uEZLiSstpMsqGIefEvTjr51uzW5U+V5B4wBEpqO2lGg5CqSXRxVt
9wCH5+qYUPL56UFQ8SYKLuNzSjvdTnf7NkwPvDVJQlFigFGH7P8jlgJBJ+PNSD0T
pDU90tSg88UZfvSEBcqq+0QtcMKhnrGnQ9TMFHxYh1sXL0HGz4qTfaPnz6/kGAat
zCqTSTGXLL2hez1SuXTQbLVh15BG43Qz/Cs9oV8HmTEQ+WOf9XxRjJGat8TtM8CF
zGgzVH/tR0MBzXYA0Vvf0aLzN4K0+BGEBrccWG9G9QwgsNADOCb1dxNcz5ZgXZrR
dcNL6ieXhk/i48ttAUqAtd8vhMshfUt7QJowH6pXLF9utEFCaTe7ymLrholni6Jr
FU8s4teOdwrM1HBJ//fVyZBoHks+3mB+O6Yex+P5PXo2YjmknJxYBvzmIgVg9iu3
VYxbigO7z2kKDa1Qyj2a2LMXoae7ANaifcPoDhyJnzlBzWh2zlj2uAW8CjUs/XTE
EGXPqNLVjjzeIWmOeYblxNKyJLyI/9ahDLDb2qHkZBWJEfutTFgMmhCN4QkYZaB8
5BBYRigPwpfpgw4rZdp6UyqdOywBlH03j4vORBKM46NG+xBcDbbt4ka9lPiilpYE
89NgFKMYbsW5DyPo/cS1IW836x0yXXcnyQesLAiwuGrEpAbLJmNKvYdFtwphq31c
yuv+WfDmHS4uKoEnN5yP3bz36E3x9NKs6Dm4f3xlvbQKMr1GA87ta0+r5b4mWfMg
26/eA0ytUglSlTsuTkg9ZNxosuPHYPXzTMrgZP8nxEIszh28nzPKhnsCTHsrGd/K
U3U8Cb9Q+/mvdaD40GA1AGbPxN6bMfSODGo0WJPbx4FOXB0fKVGljccLwJFYogLG
SrXQRtRRq1++9NHuhyx5Q5+MGrUP1IJx0294kTzWB4nwKI0bkw0JhqMtiFm2x2jA
oNVhT09MUyKkkxh7duJVz3ID6OO2SC7KpBuVcpJHHiwGxlNtkkRAIoIBcFiNB3/R
+M51u3Fjh6FmOfPNPinW/DqDikE3UXjyH0H0I88HDSI8gE3p8KjHs7Mi+kNxQgTI
DX4ZG53zTStWtsG0roXoeclOL6cKvxymeZS+f0H86FuMCYH8aU+zK7EeNPehu7UO
Ve1Lw8jjApUZZsSakxTI3bYf9C5ro/oQiw43b7ip4lOGtj02dtyF+WvQUe4Oxh9D
mDmmB/3+95Rl69DmsO60f1Y84G+S4F5gUMXe06JmBb9jT1TWNImR+rHN4nXjh0lG
szeSW/WKYdkh1FShVqjcAObw7dPzCdjKEN5pvzCSYoyUajI7OCxhwA+Hegrow9o7
arXCN57Z9CBZt/qJqhrDUH0dRwppgPvMdA7ThRImOH1hC9VWkkp2mN6BOOfHA0i2
JTofUIXgCSAZ6rqmdkC2Rkj7DPz2O8KPJsvCkabWugz87xwi8mQjaquqEwJgIn/h
dX4H8Y//fAcJme1EUCRmpiX2TkejSbLwKGyjdf7Iu90oUgE4CsZXuZAn3sxT63h+
tBjmWLyAiwwvC2GDt87tXd+261Vh9U4l4PaBcVe2xyQWcmCH4sCQ9immn+Zxc3cO
eXPJ6GsZzQNfAJCpYs3Is7lV7ljv057vlXWMmlkul9SECTdKe8byGpXpwBb6ESB4
XMF6O0QiG53yqkNz+AWatBU7sbE6YvjigtcJcxmmhyODWatzfDLO5B7XzeC+rBRl
/b9d5gTMRAkVWouv/C0Sm4nkC+ndHldBVRpBxAc5YZ9B8Sqe9i2zwI1njem5ftjC
y3AlWKLdXBesKb1ZSKfEGc5XyjmG2n7G8Cu568uANX1PjdUvtwgpxxUqsa/Qaj0x
Hs8q1W3i0h87DPWwErvbfXvz73dY72kmU9e7KZRstRPdohLvoBEBOUkIg+R344er
xJdrQbu1NsXVTiXc9+XnsdiiafLmWlS5ALdJ5lUz8Bajd25hQVQRwjre8RjPdBiX
W8aPD6yvLgaT2CAEy0GR5VCJfwmPwQPAp4MUUJsaSd80dOhkc/95/SPAJeSJ0Jv+
5bbLRRpfViXQ/30SFQM67TpGcMykICkKXIje545gJaJ+ZZB9WFZduJI4+4WpC/rv
b5a1B8JZZoAoJeYZAsCSsBKJe2vQsRnad/LPAdCWY0IUtC3ZjEgt6wpUeFX00qww
hUQeY8O/x+PsYmaNKvk2w0T5g/npg7g92yoq8+BJvrgzdA3WvyvIpc1dypEOZ9gB
HrUXRWUkfVQ7FnqowBDFu6fiEIgSL4uRZQY9ctjpL4a3D/3n/1gAuerLXNCqxgTm
Ebv6fSC/Njy1fIdMwD/fQlRFIWfQuZbqYMKkicYHrAStsFkY0CvF/q9g489iVoSv
gSd1g8oCcVJb1KEjCXGYNrxFLVxydvkvHEu+QeLLYVAU0g43MYiKypoyFUp+uVUD
oP88kr/CVXkfju7ukToZX94XZQNCX2vnDOLLBkThAt1nYPLGij5NQ/w6jh3wP2qn
ZO+7BjXNVc7bjVs8ElKtKyWTd+HlaQk55xccM4INyAXiydM8ZBVCPbdALI29e0YL
VSVnOBDH1+u4cNMnkayBebp/MtRY/ifY5SxW1aWIWNod3GT/EUQFXN6G8dtHG17H
hOKbJaPDWOgKznD01QdMzoTSWGNbrO/TSzMFmT4sscIGeU4JvDitkkec9MGML4K2
xvaGIEIr1Yl3JpdkgeqYLJ3gWbCo16nTQDQw18vPBssEokslLxl2NDqRfBMQR2q5
WSLWKo3v4sLWUPiOdxdMcn7+q1Fdvs/aevPPLlPYO1XwU6ahc/IrDtL56PMQ4DK/
R4uvnnr4WL6mwjzg5wtLcyb7IxY2oFyfcrZqwIH7SsjsxFSYIU9EzTRqoBBpQZXw
+hDhMFZGpG2c5Elbnc8Y1/f2YH9O7eagbTnimSZhNGIhVbNrzOmkftDVXcYcH7jc
8izO0U5fMkvQS0vlZ0FcKZYWPCmHix/bwgF5HyuJlwhlOKHf9CKlZJKqUl51UePq
LRM8HrTrMYdCElbl7owyuSKebfJfInYSJtLIceqVQrlQHyQQfVSBsB77Ree5Ku9K
eObI4W7uLtpJwLKACcP7+qk47bJeqG4gAP4pD15jx5BW8jfbPGeASqN+B1LXIg/p
FwfF6MtSFdimmb1k8SBOXC9YZXEfUL99Wo+bR61PCnIqHA3lzRk8hsBPZyukEZEd
gtkUhV7iOKKH62Ra4qp2Zw0OVm74tl1nOxxv/C2xnGy1Au3yPUMeR0V9IjF8DOXJ
yR94c4iPFQnLf9XhHcBnDtqyJN79zPEanRb4XarP6Is6t0l7LaKshudVgo5WG8K6
5/Q7EzfoPPCqhmrLSN8eKfzrN+jFAxYiROFqIiHKAefR7J7cZ09fpre3hFjMf07u
tGYHXCbpsbocPI2ciVaNcmz0/BRXLoGKgRUVtxQ/JobHHarNf2zdSvdu12d+d/Fc
Bqv57PFTq6P0gqJEaI6Z3nhrWN4r8CYXI7DgFLGYbqpnereXiUU4s9xau7ryH8G5
zOEEvtJK1vUlF1X035AULl90uWRCTa5J/98805vsZlc3uMR130ZWSGeNSNOkSVzZ
vr87YRUypZgrn+/X6jCBE2TQ2yN3kivEtkcDUzfcHu6skpwlkvOgF5bGpuoPo9um
9kU27gDy25hDPLOEtTazsm+CPhEWbBEt/FNfr4hiWxN2Xm89A6OuD8ufVo/FsIJu
N5v8UqrWMlEmuGeO91ZeaHrXWn7P3ZBP+1Ya7g+Et5SY84NDOOv7BiO2vXJByKOW
Uw5XhtihA0GaHvc6JkSrntxhhq6PI85T3nyA/uY9KBAsvi35Cr3sgfq41JGsa+QF
UW9TvOLFxStHuXHCSMPP0ojsnqOBTvSvRJ3zdQhbIdrxqNx+lUT6D+LVmn3LOmZZ
GTo64osCkJBgUJ+1jbYlykgZttMRABIOPyFr8U2cgktombxpMvZfy7NaYxWD1FH2
+6lDE+xe6X+40GalQZUu2v7vSaY1BTmycHO9rLUxAjDG81eeuhE2HApKHZJ/WTim
eMfeHIMmi80lk+wEAcI+2J729tALvtbJz3OfRyJbF3Jd57BQCNUNGjA7Ngkr47t/
w1QvJY+i8gWmU5hqy85PayMk6mFvk1lpEsBKsezBav7bNWVO81GO6pGHaM2aMXaZ
aJ6anLvN9B+UuzfEKpUsM3i49i9nK58o2/nEOAyhz1Itrf7dyXabPCy6bTzn6ISb
IZyiaqLk2gZ2fFSaWO3A0DqnUhXfaeJfXxMZGTzzvkK4VeoQLNMKqNwdtWiF4LJB
Nso3jplynUBYj3X0I3kIzxg72iix38oJlBhAQDtMM1PVpskWtgAd3vjCD7TroJbp
HYxSMmQ3WTsuPJalAJ6YVT8sRa43HAt0N0bEGrgf1s1CGayFRBt/XFcSNN9PbKt5
aEBOaPOeZvLcT33mGAMFByXeIh71yGqelM7Bwdhmi/4dA+HcuUo3P4mnskdLJvaG
FSEIqSsxwlzAwzQHJDSCEuO6/yPnTnvneU9nkALvvWlkZltjHPqiPlenhmIbcBpB
iIiceGw0n5U0aql1DDl/bRZZtwYY21yH4LvZwddLBtTeOd4sRrkLzjzZmaq0qP/I
bNUY4g08gP9H8CBRPk9JOPpVP2RDnOMBoXjTbrOv8jlzZdHiEKU1eEgMhmGe5Muu
SFSX4h9C4vAqJkgOUx0Nvo4LMJhoeMStqMVALRM5E7luX4xfcsvP2V8UDCt3fBf+
xGNhlTnZYIWSl7XRzQLbL3EHvJIhbHDShhOYVocFFtxrxJrTNEYsk3yQG5KQJ4ca
zo+Ij/JOsvAW8e6pobX5HP6bqtL6cShbPpIMsYxKGuH/O4lCWp6nLCnEdzhhwTjQ
hCvWLjpHxYGjMniZtfpA4o2wM6WxMYsgqXUds6PXCuGGpaQ9cjOLNHwEqLZYFBp/
u4q6eZq2yqShGJGe12ljZ0Me3njgtMciJmga2aLVEX62wJeiXtTAVMbKa7rthttq
xWTBS/+wcZuSVB5wTcJ3V/a2fTw5rp9Zn6dlJTmVUt35WIgl4NwGppGkIdSZZAAw
5belcYllgHpVgMORNOQW4drQ+1q/mVfpgTs4NJ9LYGXBFGZvgAwgqwLf/8r+IO4A
r2it4fypCrJZw4ngoRXL5oiOcfQN+8yn8JlyKplfI47DuUzCDGgpkmPEArDEL7av
bWJrclrDAoqAxL5kQU5vt1OjBXas4KStGP9SmtbZpAk4hdCRcCBHKU4MxqZeL0X4
9Nr8hjE4tnz8ZDJs703aRDtQSV7LBLKSJauF6ogFLVoG8AFHx6RAL8U1LouXVMVO
JrcN5UTW0JdgfDiwLOl52aSNpn0aDFpqLyjsaonNSB44xZprkxC1RoAt0X6QzrNB
WADnaL6oBYAN1nOB1UJRCcFZaabDgHMiCcbBvGIrOIcZxJTVfSYJZc59Qv1AX8xv
22oWyXTnP8KiIyFzEMz6fajff3KC10/Tuw74u/DOTrUMid1xmLY7YVqgrrD5RrOi
MUy7LL89aPzQMXLMB1YodRO26hUyBP+R8boZxG42XWvNQORPeeaCSX8C/OdfhZll
KGUKyE60h8CcRZIbMZLKRyGLNJXWMYBdrSxg6xGJfABP2dn7agokwbB/SMEzFaDB
cGUC4Ir15v1O0kpFSlwOh0y7I2+PU1ZsMvZzhYyppfjoGe/9kPh2l6IiBZJYabiU
8a8LsP+s59HLWKJPmuJf1y9oijv7TkzsCGbILs4kBPwdtErAWgPfPjirwbd7R7FP
trU2RxYeIC+TWrkXcoVsIdsoU1EmDbXsOWnWxtlCgm2Fx1/oVKk2KoilBoEp27JV
rp2rTJ4mvySpeNxLViIlwZy5UZJCLiqNyR0Ppl5zuHAeE7x1Th3mUj6hm9sJRvm8
cIlAvDK/8hquvnxA6iyVnKvFbEPLq8sMb8CPis8Rvtw9XI5HPy8tmdjT6/vdhKSU
DDTqgnxSR0bKkmL7ZsepoFq1z042dgEg/ThapvoAJxsQrL/zsea9LA1rg+6CID6y
ZWXU/XvyAm+Ulv0lutgKx4y03npqlmxzTeKz3DjSaV0SthGDEVzm+Fxyq8HKNeIw
2t4lsUpR+3uDNSdwWlDqxE8ArvutdrUGwDdBiSPOJPz0MpoYUpfqKC5KoQB8JnFN
Z4U9viiqP4SYRwu0z8QkFQzU7F+WXq64BKhldAN3ZfCZneeyUrZZSN7cXzlu1ycg
AQyRoSEBYdYkbbsTXrzMBk4ylYJrw9Gn/wmpitxAQDpe6Fx8FZg/XgYOFL3kQYwt
ULJ5faa2uPlPHNd0AWS7A67ElAQGGf0LFi62B8M1xHNBCf/eN1lgJsECNEVy9P33
mZMBDKr95UHYqlyfWE8T+Giypbon6GRryBoRTMUas6yQJSc2EcGAYrcnUAmXRBKJ
1cTP7BlUYgC3xFMpZsonu/jCpWdto+rhVTLMyMegIJ1Mt8xGSdeutBGD1slTKdx7
lv4XToIVhr3oHr/sFl5U0wObJFAwgIJ1jTxF/JW5VlavjSzcU9YgLx0Y1+HHKRYC
Eh08SSaHCVg59W7QJAim3VeGfNQBoU+gWUkCVJ2nRoHyJknJHgOZDNosPtHUNEOd
4zKua+dOzmVJiTaDpTIJg3ohlRFiD1QqLoPRgn51sndE4rqR4tQnDMWPXQCW3FAX
wX2u+R452sxVS5uIbuoh3t8JDye8zvt9am//ChYLXqNvWOO51jnJg8Q7oYwbdph1
muAofFc4d/doYuMNIOHGfqOIClv/1CSdUaA2zQ06u5lSpmqp5NyaXjVqrtUp8w1t
qv71Y5Vg/s050JyJ7wyPy1LTj81QdGA14GlN2p7Vi0sGia2tYBdBNdKK5LrcJH7V
xbIaIxs0fvgmDgEE9Np6uTKweIYBIwvBA0sRoGb+V/k4iWLUi7H6my3qHvHbW55z
JHkh/+SxFvmHuMPsWRfXmzO48y2qXyvqbZMGQUb284F1ofHzhkcMqZYDYFhN6w9x
AjpBvTmU2JxKGGpJOQIaql3+W8t7aTjW0J7KAsD7RQh/7+z/8kFmMmXMo4nHYsia
vpVClfYmlMBRV894rL4/TK0AP44ergnDQf9inqWo4qZEfjuwP9wHtqqekt4/o7BM
q9VFI/amBhbtdsaDJhwE9SXsV8roPzjAUsunB8B7kQxl3w/eOxBsbA+sPQCtYuQG
o9DsKSTFqTNkzTPIa+TKo5RsiwxF6IpfweMMDEU8EHfdGWJrkqNDvl69FpohsZZd
6y8hows3sLhB3gPZoAvnC3RcCg/IyPhuDwge3yrsOLRBuBWPppNmUwU1aLmoJuhc
o45khunZC/8c2e9ytcmdWPMvAvUM7kbRg798k6K5VIh/4GqCRvkekp8uMVKFpYm4
XPC4hLi3mhfspOkuV7J5niVImV1huocw0b7kgu8aR2fm60IuG7PeAQAPea4XjnhV
luv9KxDYP3HpA1mbqFdDmX8W483DI1iPGOWPQTNPLOReFcfQdxZbnKJZJgzLmlFT
IfIN49vQ8XF8e8VDyx/p4YVTH1XZNq39tW7Lgpf/kKrqQgQqJcn/d7+Sab6guHfl
PRRV8a/tjzrO4xpnichbrUAkjd1LRFokjzGwK92Bp/5D4+P+eSiEB/cedPc5bU0g
acOg43Lhz6WWf8yjbGOYUNnREHq0b6Y6lIqWajpiAfb6M7htCHK3FP6nM34nHcX9
znIRX9RnKNwfwoprRv2E0h1MuqfSwDOkSf/Uhm6JKO161SArGihkJCtT7kn19gNO
Dyx5Dr8+6nIwvhWuZgg0ABnGMuVIJPHdUccIOrQFMHkxaJf1+hFz9WHdbkyuR+3R
gu+vV8cdbXIQwYF2Vdlbyw/bnlXVZh1Ek/Trmk1vQvL9wRHYWZsCWvLtwtPQbJgt
jiqu3fRNPhVyIDGIqh2URC6q4iTy4kCAPXR3XTfAvOgdy7Vc1fReJwhDe9MBPU6c
Quy4iBHgAkKakGQ8uqSB6pVfLak/lpexNWJnrdLcqpaQqJ6L1Yf3H34+OQkzjB9i
fC9cXXPElo9SK0uHlJFr16uI4c2sDoxeQ1cmyJEgYz3lflIHUgVrQcTMTJFF/QE5
DpeS0YHI412ynoUEosizLapcOnr4PHs3fXRh3PBgI0esHj21mJwVwtElqY8cn96o
SOufO/kXWssTQGJjf+fZWQDLwt4LIzP2VK7Xk2SaP5BvZj4VXF8Dv8/UPvKp644y
KiOaNG90+nKp4hzepvT2az0O2FOeTVOAVJW4stDfzG0MnyadKSUTyQxus7dWG4VX
NOSsIUTrTcw39HqBw7Ga6yrnaaY9J337RJAPnZ5u2INsaeHpJfx9QnzFOR6VVJWK
TSDvJnoljmSirdHnbDM0tpQHzJ+DbacL6BeuPxizksU5ebwYBQsTrpsS+8+ejRR9
pURa86oBfqdhfYFYVQxeyfbeO4N34ajE6PGJXUrTEKXuRv9FJ+6KPXw8hHYVFOsE
8KexdDm5iCR0WJW1FHCNTrYLXY5U0SkWkZoZp0V9YBdGa1Fztqj4bnlJuDA1iodl
Cr/kFF2TA5wqNb/kvDeqbyFqWUrVe3BhHF/pIhgw4IDjYvz+A7CJPw7RlPGItIoi
Kn5YqsCFJlW0h4Th63NOaTOLM4XT1QTj4Yo3MSqF9EcDy1zSJnCRnp933hETkSCO
QXUxAG10H4tcpXCuiU/gqPbhW7RBetsu/p0e+URI0mza+TqYBvNNyaOrUzciUIxM
Qkm15Xp9N0lDLZKSGcTFY9ZmwBwEOFk4wmX4dp8UFymaNI4Qp5IO/WTMs7ygTM2F
i9W4gDEDDDGHcMW+TDPZxShsK4Q9klH+b9CcQOvlRpM5jWcpwUCypdN8wGwXA9pW
OPCU0rZ7qvFHPiOanm8RI7DzOefBZ/qQboigWwV4mwp55NK1cPKWSUHonuFCXTpJ
5FIWOUdl65G2dch+qY3eu1ZQCA8mbpxcXlicHCThB9fxRmz4clH78uOOXAYjrRXw
WgDpra1AhoUV3/06gDuKHYsvAlpSKFci07bJ0DPpnXgkdRipL2WpRvuR0sF3zn76
R6TVS7r+ytJoTZNMmHA+YFF8blQ6SaA0tph2V5acG/0O9eDEDaW80euAeAROlXex
96rpyF8GbqWMxhFdXIjBV722wC1erIshlRdCd+qwSam0E1obkheGWtAk2oSNDOYo
rcmbE6Qocu3LaaymUYRHR/GsWIDCo7lnYhPVFJCpkhMqsRiW3DPVq950VgMeDjQR
3sLOWEL2QDRKUP99+Jui7A0Keb+BpPMLoYktix9Xt6BnfnhiScHQtQjYLA/qy+Sx
mdhN5au6oVYVnqeh0SDFwCDZB+3ejx2oQtYT0kkqjKIuOTS0XCn7iAo03CY+sok6
sisj5sXu+htM8qyNhZMZZv5dOpXrGwpOg8wUBN3yTG+7sks+homF1Yw9+5lvUogB
dbbFzIUke7gmhALgD+JbxOMeoYHxgP3N7yD5Q8IXg5+nSBhZd2pCoEKgJICtVllk
TdLdJZoSwzXk6kAMpqhUqXCymPz64r0qNzAwlglXz0tXzUaZ458d9gO5Tv9YjA3h
dB8ZbBJD6aYlOQH87J6ZaGR0jeBNKf6kOH/FJxO7G3bGCT6Xuhl3/H1sU5TVyjzi
TQqs726pi+XYPQnaVkthciEn2nq9U7mKf7fmdMCesRcwnvQ0FRWjYPMKdPpOHYwa
cNt+YuTMEGl6tsPLTtwet8ViV35yrEv+M/PaLfGt+iXz7iSz0gIuVsAJJRK8IVWU
yP9MTgXQdm8ev6BImZCxIMW2s9UF0kym7qUkk5241NxrjASt+GSwiUxi7hVwRzx5
u2ofUTSj8EyIc87QsW3onLTwqn9ttjFTjSd5Xv1AoQkOs1lLoPuqJnpxZ+Bge7hM
GAfUXKxSNsN7xugzN4a4jKbSAm1O63fkZIGJ5q5/aGF4lTUdKtBYzBzvhBxRDaIw
e0JbJK7B2pxf+IZdXBUVNYwRr2jo12CjUDtjX0p477RfB/NgP0s98cifwiLURXMu
TBE+oHlBOG5JhJWjU2rUlB2Yol5aw8dlDcGODF9YjNciK01FDx3B5nmwgwb4H94F
aPteqd9NazGiCESormuvyqY1jUZ93yoGSwvln3ChUrF89ncteuVkhvp0ub4i9MvB
8EYntAcIHtCxbpK1Zns96Q+VcYT78I/+9cQ0P4i/yVCY5lYZ8jTiGKt8kTOeGtQK
OJEs7/3d0hFXly/lZ/zPoYtgMR1brDOjtg1jMZO8LBbBHzMA9zcFyiDifOlepNJA
77p0SLr7lSH0gsGi7TkzRlSeWUWYcfhtc5tE7V/TifrNSpnRqFyuLcPV95VEawsa
k3c6HqUfdb3e2TLoPj5u60C6KQoDPOaPAnwnB2sNpt1XQ/p0cpLYvVOIZIjhruav
twcwG3P09cbJrKuHbxpgjoTiFEzwTAAFHgoB94UxiraG8tOhFvEwkt+jW/kgkN21
Xn801dZJhtdnwGW98sEB5UjXqy8z3+kerVJxi0pt2HUqiTwb3ZXqjUdTJRNdbIg/
SoQ0VuWqCCMm1tZkg1T+qtwMSEBJTm9c6M0E2HlEZZKdwStIZhoHgGJXRRaCsrt7
AmnKCLMMkaoKiLUnEU82XHuxPqyJqtgN0xm1OH2Tn6sT2QeGwYkgJJZZufpHFwtc
y8q7MadDyDzkkO5AMFM52eSqwFe3cSw8SFWQJVlD5sw0tOB++NQBmn8FGgOVNavk
0pKB+XSxZDfsTEjKoyUqmkpUILNYJ90V8QYRR4k9LZKfFYH94D3BlX3jluxXaBEx
n6UcJj+Ti7s8EHGH2Fdxnxp61tiUiNxj+QjUmGngyAbSOELvoLXZKAXvTITHz577
fLAuS29nLzRRpSpxdw2nSMSQjIgX8kQulxQbUEXeYYAWNxHztVJ0+Mg6Ygn44h5a
t6eIM5L9YjcSyPTToewQJ7/hUL/MQNRfcA57IkmjZ1LTU+hhS+3z1YgaVixOABDQ
+Z1/Gm6kKVw/a6H5tkzK8OXtG+4OFRZs2j0vTFbIs42o4x3ptNZVQ2h+dahPdT7o
XlgcHDPjZaiQjCoKNgvB8sL6AjdKwFpw2sr/8Q/C/0eA5+zPc99vtnrxhyJYjGrt
jyPxBGtZkl3ebL8ghZhZFE9KboVZlG5mr2MkCbq4WA9h3dqVYB44pLo1mRTXvVS+
t4h1mf2ktSE85bi86sh/8bd1ygxemhgMHMMGcm1adioqztH8NYAJg90+u7rzJ47t
yR2fJehIh4G9R2I1C63LruhrgQsyYSZ8fCaFk6ChaLmJ6Fl5K7WY3PGy7L5zxMxz
Um7JhWhHA7Oze9j+QhMwHM3AifHGefJg9mC5TsiBFks9eOlsj+jtjBGGdmvGCQ77
iDks1JP3VVLY2lRMLiVfnqeTJFV3hLaNjhbE2UqPM8lJa1dBuOSsumOAezTMJL1R
nGSRx+vAA5X7qWVoloqHFOnhepdVS15SA7OGM/7UTlUH601vgKosWco7y1GucAWQ
HTHq/p0WAhEbHzSgOociGh10r3DCGGQDZXtAxAy9v1S+FKExEOnBxCmjGWbJxIol
mzhXMTsdqFmhUrriRg4ilQopUXnuTG88kIvMPJBIKsJg8nv4EOiEw0wcUjw3etPl
1a81v6Yoq5+kJRz4ZhW+KqshjUkPrJHqIhpLZ1xMSaT5MApUO80Y5919U7g8qfOe
AOmfF0vJuy30n0xOOVakej7mjFVYD5mhMU+N3a6aamRgWf+CRm/QTkVvg6zQ0mzi
EWCbvtYO40B0Mb4J0XU5NuOuLYJGL6oJ83jnsYz9hc3P6MYdRq7SQMgFCacaR1VD
q3edoCdt12WxeY9A0lJ7YHfDm4w6u2297izdFnUANjqaqo12HpwLikiM2IXJpz3O
Oldc8KpbBLG5qQtCqXx49w6SfPIDFKgyXWUsSHkOdNs/mOo6BhO9eC7rXaydMGKV
EWX4f2z2dQpzwLWAHoNmSbxl0gS2GwEMZQ5bB3x/PBSudBjXxMZ1zYPqeJnxqvZ1
laIeRxTB09rTj4r4lq3w+X1omY+zpetw5Fev54LnyhFKxZxR7uf2hs9oJkrz4yW1
8EalwcF+usEZER8jwChe7L7+mut1Ke5Y54KT/NacJgV299x/NMaaQo8Qn8xojdJB
OgUbTSeWg9Sgsy78oqAz/nipAlyS4cpIU+WA6Wqna3xtIWtMw0QM6QYHfPW0iSBp
tD1QZSdVCX8LpERSQNCwnPLeGuMzFV2H4oXfDa8FwnDsT0RzLubcFQkJEcbR6rP6
2C1o3hfOigcRVFk1c23Z86sJ/GNLA6CtAOFliLRlX3zPBoJb3ky6tgvgcFqUGXoV
2CQoyhA4XqWmY0R9HWPL+6deY28dP63Sm0TKRCLtHKmXdmwhFc+5kO7x+eQ2xDU7
kRpQaZJ23Cl4q1Zn5vU1hNbbUVv4udsbACkr+g9mX0dizUpGiKG8XTE2+UiW65J4
RBglIXdwATHo/hZGmKGVr7hmkCL1l2pMjkUoF8e45vAVN6UeDfYpcZ9SA3uNR4z7
JWimWHTNeMqJuZTlqOA0nlokK50CJ3vjtIMh16iCYvIyl0abADZMBbDxJHBSoN0f
g+gqJShpsQ3SXOJD7zwrhXBPQ6lvXL1ydR2tgfp/oQIu+qaIQodkLdt4i5U5VXdj
431kCUK2tURHclLzNIVTLEcc10V2DDd6VdPg96b1y19IYpFopTDba7D4tnLQOi3Y
0UD5AJWXuSGjObMu1E0qwywL/lwdn2uYaeZSyViKs9S0SehlOm7pkAwXJRDTrW/E
ZCEkTS2gzWf6aGBGv1HwFWvQGqoU5cWq1mo8IRF3JxYeru1mPXvVDKPsC0ax6Bkg
CGvPWFXOsgJXGzrrRliACId9I/ELdoD1x0K3iM7XZhVuboWzWMxPmQVG0BMs2lyZ
yUeCPrflHOLinZUlfYPF5JuRUrrETD6VqTAv41UwxCmY9/LTwwVo/Jz022GaHWZB
H1Q4rkhL/H/6woDK1M41Codr7pqMhcC8KM9DVkuj0XI61JIFWJa+YpKeBGUMsNzV
oWOvrUxfdxAg5Bx5NPwcl5A5PXpM4t4mNtdqR7bp6Iaj8GNwqXP3m7mn1OUe32em
INguxeR6LC0vIRDqmpjRhk4ZrFHB4iyjCruZQDeBYDbXDd5D1glplHl4jSLfWinI
NXMh5HUK10Pi0L7LdUSqUnim/fEkxHi2gx8JUmjy1JPZV7viGxc3GF6g3V7FW+a/
CONVoBl7Fq8wcVixG2Le/6cZbojMr3A3V6Fyw2dDmc6N2shG6hcjxa8GQnZw19Oa
iU2Ov7NTXaTublOnJle8B4HIA+LQW90m8pfApCUVNbA32V2GVRxExPb7omxDz/k/
aBiyrrfEq59ys5lcqKq22dDFL9HVXMskU5WBcNzVtE7YJb4CdG1lrNdsT4ysCexm
+69XbclrycpwVu2Xh9aEb6wgdUPvjRfaQyhpodnKL36OHb/xiYNZmmvtPkPc+AsM
70dTcG3O1CoHUuXn7IQVQh7xNHEeWOLTshEm/RazRzzqAeiRMBHYR42hR5Kp4SBO
VX25uIzHnFyPU9Z51bqgnnevNMlWca0MWrNPvcjl0qgvhwfRS9ny4dlaWhqdLqzi
ws3J+gpl9mXqIWDvgyV1sKtFr+iMEyj6NkIhYn5znn/lZtNnQqI+ZKvcisFo2Iz1
fHryxtao/0A2CvfQHeTG4wQdJIbWePxADKnFYmi6zlNe2b1NqUJwyBi3WeXwvwB7
2h5NwPdRjXL90B01D0sqHBymcUn3vHgzWjFx0dn00dJSpZm6C9cjGS+UDTBEAqnH
ZbwITTVGxY6PWvJn0fJONxMdjBpHEyEvlqwz9viDBqBmcQOIQYtkAnn/Oy2ijXwr
fEieqmDFEKwAMfamgH65MNHgeIBMTASUudkuWa/W7IBQm7oZm6xCuez6wMOPiGbb
OU547iFlAYd1yRXP83ERzl6zF/SXn8H5WwwZfKlEYMGZP8wuyDzWcBrX8XuF2AEI
uLQaHlRPfRasfiB9yitc6LdcR18iBaTd8lUkdporYIBdAn2lexYAW46GUvQUAvxm
AUvB0NvLR3SyakzP0UmKdlgiNvD2a3WdByt1Of6Wj2EjvfAaZfD9nSTEaEOZgkz5
sFx4N5XB15BKgTueTXv74xy7NiwjeBVYkWJ8fabITd+iYiYPuc7RZPbXaHkkvlDn
9DV/NaE9aF3Zzuv7wn5PvncKexH7DGSCW1VZoTkXVgMW4YMJVjoMmR0ynHdi0X7w
qR4USfgTmkUGO+CdQFPKqejE2hFgWbxYQ4XDH1iaXmZalZV9AC3cx2pkDGDtgyso
fjs9DGcggC2B6VcLNr6r9iREw70vHwA1uSkVZTsu6nxF8fxkP35LcHgwhBN4Imu2
13TJJ3GYQHDf6aQU0qaq/nrv58/hnY243HljxyRMjTYSRDv99SVqqeRVvC5IcBkv
xThyAOVu8B0rNacAA6PxTDvOyecBTmrPfeA+zlAhR4nmZ3U3WWlc0TGOk8AbCRGx
+YKccUYJNyfG3eGOHdaK2K1jxaKo4Q1E01TAiua0ikSobOE5izfzBq/di8DLAsty
6vi6JZ8ET9ym36CUSGtcG2Ei9ZaTGNNxO325vCCKlLhw8x5W1X/ddaTvuB0MQvgm
extfDU7EjHxc7APAibYVVU6Mot6t0wVTIdSnvfycI2Bs9+rdLrA3KWYAMXMTdktm
jjIDVFnSiLZJmaOnt9gk80wUXgd5Z7GtRyWXZ78Ge7gqibAgfvaO9HEbdRemPI7j
uD/hXaw7m8xKL0mgeKSPHldQIS5chaw6h8GTDDmhYeNjWjdowuBMqlj/D1U86A/T
nFTfmYYwHvGNTIBTt4YD57fyo+imfwotcg25lAtpEsEmHPJDj9hYNU6V2MoYVZO2
lxjBM4QugansJh8+DBrZeFQVb5QO3tky+F2l66HZUW2Wx8rPyK6j6i6etGMZyPQV
6tO2aQ+BDi0PAJ4vZQqDTEPcvTptoFGxI9Nv8xNs48NEP1d68zl83yN9CKMPSuEg
AumIbtnUfTowxCM9BNOEpYXHGCDd9am7mDGFeNXrx1U84yNlfQho9tEyRzY4vB3h
Z3o7wY3C31G4dBUo1VzsxJ7L1Hf7KzFAoRHA5i+Uf5f23ddd1uTgBUAbV01PKl/r
TSPGVVMokZaHdY0yhPn8F256KUwsfgKK9kyP2V0DqjYT869ZngiYhyEXz0o3Cxxu
H4yZ7DlyQQ9g90ktFgvRLYMCAuJFIk0qALSZ5CnrYVa+0nYdcafWVMapcoXWKKSE
tkziKVH3GHiYlQQcmfmA4E98LKjP9SLL4yuRSBnWWTlhQKyDal38AgNdrQW4Kcd4
BL/x90jXGG7BJnuTZBs1MqMM0MjKol+g2B6Yi1HLIetv1YxISZOJsTWGL2jeA5aB
G+gvybGEzeOI7UzOnjVL0rviXeOi4uKfMQyxbBdqfDflnb17bAEP7eVB4tCQO1ir
amevga0GA0OJsaGTFcv7fQeqwFgoeErS/hSJA6zc/b2C/q6t4ujBAlv4msQqmz9I
TOH3Wjaby8oAfg0WgvAq2pyq6v5IRgxPV561OivLbmQxgGf38ZGbE/qjbcKg05fi
Cz31oh1yOc0eAqIVv6XkdDZ2bnUWhtXFOHZUMMQcn6SgwzJCKuYzlJDV2ibD6ByL
8mipTqzXWnf01qNdzquLIivtb32HiNTkLvpfKbDki0FP5tz/I00oTQFmtSmjYBrr
hpsr0p0SBY3uyqIx8LhAvSVER2ojb4fQIAd0tFOOM0Jt9SlSK70lHbfoDm1UTguw
cyg+0N7UdjxTLdo6mr95pKq6gt9yyKDZPE9kPeJclgAHbsfKvM/AVdtCoHZnzkiW
eVCRfUQ3gZ9bHM8HbSGWhbCnAlVQ1wDJZ/oGIeDabN9YTglHO2NJ0y3EnPZxB8y4
8OhLwuByUcf0WjINpj/Jm/a+NTyol/5NoJ1P6KJPsFzsUvYC/HVhS2nYs8Wc+WEU
iOKDeV4xXq7Fu6EpXDNcZUKGH4vc68UtLOnHCsErYmqmymajHafJ4kOIHvlWkwUY
SUYfaqjy5AkNKG9510MVQ12iN8YbWlW6UBsypZTCGT3BCOxwlpaxaOP6gtUFc9G0
UiIi8D8vzaZYtrjaCHgLbF4rOFzWBTdWePrRe37wzpcG+594Bkv6X3OJ9m6GPN6N
PTIlUR3MTi41Slr1u39B/ucYTskW+Ni/6Px6qfnwG6+26tP52JlWRF64WfmqOBDD
JWw0JidrlI3RmFVPP0osFPRu5r2HYVmi8gJ/UyORHO5pbEQI06JKzedGYlbPT6au
33LPOSIPk+Jge3/cwWb74BpD0zFi2QfdpHX8nPVDyot0Kgp7cOb8t7ErPtCjiAqI
FzkCQ2MFZUKpOY/MDgq+rc/oAz5RyOwyCJbCYxOhUr5von9tz8uTxN7iroreXEaT
WJ3V0O1u3dCKMSK+kOs9MYuFk6Hi6T0Fp6BJxHRhWeIX6TJ5Gi568iW8BO+shRNW
Vbjfz+rmi0AM3GwfVLULH/lYzJWKXpX2ey27aIWk03ccTWn/UUvjg1VxUXNg6Ba9
ev+danmM2cNvsIK5sRxOwuxHZsqd310YVTqvpI1QSua73JPw+ZX11HnPmVWmZ+iJ
UmiY1q0loKSFzbSizdA2fcTZy3vtbWIC/hBSpkYbNCL6dQ3txHf41jWn2iOH8ZX+
x55ULfvl4SEJO9JdEwrUprb3No0lBI9JwAGmAtaGNGXsvru/K5z/j0Cgz7ap1+YG
hNamFuL4+j7DrhloY1DTEDLmD80Wna+BD4oOEt+BFhSod8jTlFCyFZ0gNksvpvRg
mIKcypeTnaXBZR97Ot7LSOvrnnZHJMAbo1BwVa5aRll5vQjZuNhlzqnBOzpc/ZGN
fe3gppQDv0rysm2vSt7aZjzL6Zjn1MdZrxrlhS2LFpXToZ5+yZQfLwb1TCdspuqf
NwPEvR71Hq8OB5Zo8JrDBr4MKbb2DkHKQeVM49RSDdy8qUZvPridHgz4WMf2n85q
EteQqziAN2H27FvGoSyic0iZsc7EHk2Os6O7yDkh3ocZ1Un6Cr/N3LrbpqtPQ70m
tzg2/XxgCqcyulZU7VdAeKgb53sA9SYmvhHOArnNF17J32ucNzs62Gfe4TnN5hdZ
EqFsJdPf+NH6iwLaOO+FjUFwTLoRSpFvfJ/1Xm35yl5TJ45JMr7TtuVBoIRAFGKG
WQHZnTz3IIXrpHjZMdAjqnl5UHVJyyYPClC5hS2hvOaNLGyx/x/++MLBuAoVSaXC
EIq78nY0BAXQctGQBhpBoEK584X2oQjUqnf94UCY4bdunlO7M5jGtHmx70c+c+jH
arkocaYmtlEvgoZfXYf5EvAADAy9tyoD9jaa9oPt86/Pvy76xH79+kuvDbSNxd8V
0L1RNSC2xxrI9DqSq/ZCnqXVLAwY7diGoxFa3/IhYU75I8tWG1JVTR45kbD8g8xE
f12yb0UU6KTUdyWdIHkWy+hN/f9ftHkOP79v5KnX+G4Xchg+PKnSbDcs2gz05mDB
/tDg2n1GgNysuZ9OnoyzmdMjwruok0BuFsNEmCEI1dxB1uTagxu+KEyKtmjaB7DL
KmQ1bqfH+mYXRanRgbC+lkZ5/9oXakMnBWueAPtwMp5OFbk2pCvUy7vnxndDGgRS
tsz5NtpD5UM6ypmq/dk8LtcHgNc8uo4b870ld2BbyejODRhK4f6Zq7nwGnVksQA0
1bqxmxR+cg0wiFqUhqn+hX8VRw5XJuPHb6okOXXkFA0hsXjLSkiLXawAlhyzTRTi
+SAP+O2wQT73374r8xWr50mvHAWzEtuXZYj818AdjYqgVR0CFHZBB3tdisvHT4m9
63qeKyjdfwgCpDm+eaSr9KOvvqXhz1N66qy2ohy6/AHj2cPnV9/EUDrw+JbSq0o0
t7B2KFdAAGEQKJYqK0s0+//6Th7iyZRzOTwvPT3HfQKVc3J0stSELIHiGbVBHSkP
9rV0ZRuQPOzE2Rr00LPxtJRtvYoVpC+5MCVEho6HnmXGvbLDIuayLH0fa1a6nWxq
h1cxrAPsvNVDANgAymtPtkd7Og9CDTkyB8dKaYa48ODb/qJq1sAMX6Zhc4zZNeKP
1AoDivMLpCGjxOhu0pGO9MZmpDYSdo0/Fij8FhgkX7zGo76qAztnoOCXCcRJyDgY
KOOz3PM0ViZHVIB9HbgH076+Dlpaq6v6Jdaz1Z+7lCXxyuHRJhoRNRkqdPaxgWym
QGBLShsMxQTRrP+9XNw5dsa0TQTic9jn3QU8SSJFo3ljUoBm9DUNb3yyyYuFQZ/R
fEd2OtX3OZaFbqj1GzoWqniHrMZ7zW6Rew9XEqZyX0NdFW3gAKuyIKc0hu+8o5wI
LgTIfzXz+w1FOmLv6T8+kw==
`protect end_protected