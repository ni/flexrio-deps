`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 50560 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
HdytKcppDjja7VfYQkCqvOxoF0fjBeVs/iYvAit7WLQGO+lqiGOlk+KMcvcL4iiq
wFvza9trDNurAir0xEnfshNnOl1MzuRTE2I97lGJMV7tMkUrN3WIoPBolEBF9A2u
MuhPODdQYigIxiuvh1CvQ2QxPquCS1+Aw20vmY257/2QbiWuOVNla5XSI6aIL1XZ
ZAM4Us6+0eryHzzPegePJr3O941r35SupnXGffpGkb5vas7ol56BdaHm+mUV+S8V
QgnDt9bOOP8/+4SepLXxeLj8GuTDD4pf2sqziuUGNdhgNRqObbfwAHnR3trtqTyi
Q84MBPCGbJj+LQSg7i30IxDpvJojRoqmerAl1/s9mi5TeqRKIrb0nSAGkMI5NC2q
4FAUmuKx7/IWLafVkj9RZFH/LwGdJHq+QcIwFPHZqfZFdh8bjFexLqXnFbihCRma
985ltLqBHhbwR7VaDt7m/za3P+JjpOUZkFcRnSOrr83A+3pmJPzZZyXgP+Qhv3wc
BK9OgjOsJb8OiAsPgvByjZP4yXc0Ry3RchrrXeR48EPFdo7w11oPEc6Lq8Y95+lr
JmRmFQzxGMwm1Kj21L4kT4LvdzhVcUlr9gyktn968XIm1D/7rSY+vBcniQSGrEay
Hv+whFVvy1e/Tkg97UWqdZw4PRUTOxuPNNHw6JOm0J5EkcZ7nmftt4Io/zjjGCez
nP7YWGFVeng8udHHIKXuUa6Y95+8x38bn863A0U7Bj6U6az4QYFWlD7BRLE9aOIY
ZG2bHLd7qU8/FEkdSTA6Cp3ofhAVZsSUfpy+wuY5+PyD+qTLHOZNR/2cSNKbdsCV
2xVdFF20K9otCxjS86rZV/jmpnAYMSaF8VEY3GE4+GhdyROGSnGQwgN2GM7yqU4O
QKGtB9PXxufxSpQQ1JRGvGu1cqw1Qr6W8ir11LrzS9qKUPLMb6hfUe73V3GGiGHR
xgvFjyJh80PCv7yxiRqN/I1bSGS/MnxIBs5ekZWhc+DNEuehS023IM8UlrClRBeG
Ke782qqAhk2d4pU1FpV5OEi36wCjuVqydvMLnfB8FhAH/h8va49UOIJ8GEq/SbpF
toMwyOC7/+S4hyQsD1ZvXmTAihmcNYQq97AYcto20qMe76iqbfj+Gta5b+Lc0Dj0
p3hTfHQF1f6Lw9Ixtntv69fhz0ah0Zu4qTMV0pL/Jp0HY5NutJNoWND8ebTvtZeO
xhJgU1uHTUeT8+NhxJ8L4o28h14/RKw4xu3BfzzPX0SCfI5TaK/ZfDQTfXWoSNow
B+kqNAy0oZoEp4dqntikqH04OixCMkN1ZAMfaar3n69j8Eu17NsdgnO+Fp1cLQ05
bBHQpIQx1A7RRLun1EHzGDyCxJDbz2U+ekpu2fD1fG79v7MdHyZUu8BIbncK0XHj
EGiv+Y5nRcltK3UOkr+Fv86WS5tBy6SfE/w9/LFs27/as3Iaq55P1ofchKwBjDeJ
/FK8gXwrX5Sq7M+c8awQy5COXLntllG8aZOyAzdPExo0v5qyMMkDmqzrUZP02NDA
hmkHgh2KoIUIUEBI81Yv6bfj41OyOa8yeSIKNTKNyYNzUilEPWQcnLscNkdOEeiQ
yu8fYpxO7MaPNZ5G7Q07/wy7297jw0CQIGVBj6nUPqpFyg0jbRKctjD9NDsthxkg
tzdnYrx9V4e59ej2s4vmcgSvKUFmBZ6yxkyMRUn87o07QdnEDbf7orFJq2dnU+aM
aJbpoQGcMZvsDblkB0UE/ZJcXgbXfQ+apUzCFTYjosaKKYaMYFoSlpqnkMG6GZMs
eX4CcKP9VeLetF8+//QNQQAs3PX8v1AZ+Hls5FfBGDKcmaF8Aqu/N2DJRmUpwMcO
Ha0L1O23hJ0hbR/Tt3VS83w7JYPqJblnrCn2lneITzgxSO4HJsbvXub94D5e2Avf
vfFyqwvnsySXOY1uT8RqwQzNzpFhssSsN9OmIoOBtuYHtquX5YqY1l/mEqrGcjue
qzKfcuARXuno+lLLoWu8lbLK8E1jgnPA/B9LJ7AgFtQmU5DCfPrMx+amPGK3Yhnw
7O8g8Ll0gk2matKw8c9Sj1+/qfkaWej7NOI9GpoBF88PsIGz59x7iqn3qxjfY1mB
7jBGWj8FnzsUCx9wlhuhW4WjUschp1Gm7tJq0+IddXY0JATW/LWJthig9Yw8XEUl
l6v/QcYXUUIuvHWDR2QUATwtLXob0dxL0cfkIQDdP7WUgJYDSp/26SjcgPQNU8qo
MycWc563l3QIT7zvMJCyh1j2S4wa77VHke9po9CyN/VaXkFSnyEHTkoojtzTXsWc
tR4OHvCjsjP1eTLR33f50HywU173fhhkM1yEsVwWR5xZawckAlZpAyxJKrEtDdeO
9l3EI6mQd6AZXXn7g+euzlvZtzmGC/6+2ZBzCBEMVFYMAzfLYYGiHvWx7fRSnQmV
vWAL0SbkWWqfO3a64WXt0OqwpYd4n04KKH/vJkgv2m104mHG9vcRbUgY57/3QcTK
5oRAWZyBC3cL2pIOnzakTX6HV4bwV+w+pnlVucr3uh2F1Rm2IGzFeq7FfEd4+hNs
HDfQ8KwYo+KgVXAc8GEY8Umr2BOm5T3Lsajdk5FLp8Lhq6/cXw7t24yeqZAY/kd7
7/prs1OoeTSbJTy1tGGoTBYPePiOFtmwlh9IALkT06C+2oTgQarJRXAbq+0wBTI0
FKNixtPHU99HnKVObpv6ldadIAnFwbF102PEyrFl5k8KmdcCrQ3QHOz3UzluxBnt
eP0nkKqwa1cDMg6NZhWNssh2GsX+L27/cfsr3ra9QnPlL05GhnLKpV8H986U0TMp
ddDCKUCj6uwAOMQ1AL3b+TeLjBZvoNhAp6U7qreXUA0tl5LIigK4WdxL3fg4kwiS
wN0e7brTiKjHaER/Lm4jt1zvp/4aU3jEvMlUB4+IJ93d6PRtpmMB06JshksWfDDC
bgLgLIddkj/4ClQV/6NUhvj/alW3x+hVsnOtqoY0iwIzGqsrTk6uf/xGEdwegDcs
Cp1LJpdP87K2A7x/ZCXEQ+V88v9oofeI5YJIE1tIuiprw48dBGXkP51yodquLbwW
pzRZazbbF7DcpRFxZlOacis0igxCJgC4Feex+4R3cyTjtkgnJAioZB9GR6dRnwvc
4hf+1X0M3ebzfBJknMGFl+3Dr1jRU2WBZP0igYrP2FIUkOIfSFWWx2Ad4n0ZiyE7
31a+acwMmNW7yDOOV9W540m6fBpzziTwMVILwL6a4k+wbn6D+ObO3JZHQWxeU3qN
fqFe0DCpob4bKszDX3sF4KArV/OGMcBTRg79ge8cqIx/vlBWekPM/C1++8rDbkvd
IYTsUQyyrDXUSxDog6lVjt7nDnMXYvK1KJKgdpaX3dXKFiQ5usyBwgyeNcSZQa99
S6PxiEZe1i4o6SG/Cdci5nku/8uqhG/ed0KzY99bpSRUKXZxcorpHqitWaSKdkpB
JgTM9epNGz0ODHJHqF+6dKH3lJpXNk4o5eFTW4tEXBpO3Y6l1Ld8KrKWpTJLMqM0
GGlI/qibSJMnl8+hMNjEKHHJ0+XSu058yTOyK/2NOQzKOBTxta/iMPl9HJmpzDql
o0oSjjgVcXRjBFSGM+hpUGC20dBe1+2MVPEceBnVNvmJntr3ZtlcKJqE1a5hHC7/
sJ4gyOeIfNXz0OGkKarX5iUWrYK+n/3Juvn+YLtvXpWgrDo9w8rpJDLTYhSlArTG
SVYdxeDwuL8oMmcGtjAIoZJCHJczgCqR29TlJcS7NbY0qlZ4hMgvYEXH/5BpzZ0c
fbwMBmLadu+V1KhJUXH+4FQCzu7c4csKYyzpNyvB8tkqdW0Jp8kzbya1cjuOixPk
cKYZ9oX4PlKn8oMJbH0AvIM/7mW83QeohRS2l1YOQCoVc8yyH0Q83HJQ2UsVvp64
tbcsGSgsr1ndW7XvKRNqR14E+n8CFTIx6ZLi+ibE0fhjHJ3dKV74WB8hlgJmAOYK
SoaAtkAFmAMYtw/sMLm/4GtGYQ2w4hYFolLHrhcOxwXoSXARp9kKG3rq8z3K7X39
R2VH7ZN0ZKGc3je6ZKHJeoTEaszQJS60Iks3Kx4u8Rn9+IQcHRAt1G7bowW7C2y0
mCLE11zVCG1nc9apZtVMyTPmBQ5W8VUHBbZ/cxW5T2hyzHPlUVHKZWRfUweLQVPr
O3sBuxXGs7swXgAW51MLr21KrCcOypaqCYNGXmklzTmUJAZNBMwr+/KKFLQjG6Qh
a9/gAYuA/L2XADzg7+LRdXIO6RSkobL4OCCYb/uGjkfjEA1P2ZwgQf/rgOBQMuvg
Yr5KE+M5WvZhgHXxWc81bAetazxX9krA9Pf7Hg2xZEjjXTvFYtMynCGQ3hx13Pfn
piO8Q3rHd+gLmX8xnS7Q+ZsQAaru8RdDBwKJAxIu/81HpC04W9C2itJXeEeny3Im
p4CaxAZrIwQ4sQ3VywcebuohncuVZ321cZI5ePW0jrmFLGzhfF8R6RdXpNdHrs4r
9KKlGGq8tp4FKXrK22GR3Zb2MIdXNkfuyOZfe1BTbzX+2peBpEluWvkUg4l3DXiJ
RP1osM7Bw7ALK5QVXSObOETXMmsuSA7NcoaxKwlsluhkMf9O2XHlHL4Q4GIDkO8l
DARGcROEnDAYLaAkoO19N6OCsW1DTDK7ky2MJJCYkbazs3VFGOJLhhHgWFV3bzil
6njylaPa9rK07TMlA2+Au5w6loiq0qJLn6fNo8Yv7KO5ATbJ8RnfiHEm2wfx3LnI
1m/8qOEJomgY13+AqaIgx55BBirwJ3WiNPxAx1I95OOFulNcjthZO5+lgIIljtig
OSvBZiVuFbOuMnrcK9vZ9w3lsZE2G3jHPr532vSgMJz1Hauzj4uYBhNXEyxSPyOg
HRtFCOEVVi4h8/vaq/jqCaqxwKLsMZCrnnuDMQpgA2mzDgH8WHhgHdN6yBP8UwHE
nd94IVwF9VRcm/czZ9yGgltMz/H2MKzle9k4XF7BIMU+uO3Y/E2QbVfZH0TOtRfM
fDtHieLFBejZhcomUFD0aFj2lPqaIj4vvcjnQm4QRCAg+fa7mDQNWKo/U8o5THSA
TSB3D6rwLU+Xy6VRggPKB/lQZvprzatUL5AesK29AkfomfBEGwEhXiysM5txlryH
pa2feSZRa6I1P7KNkSyeOLRUeQrl3jI8nUkEnvNnQ6/z4kESIqOVrAf83ndUIjBz
ac+jp6PEJ4xeFkx4AGumhQkrjgB+NKRistvkERj8hqBHF9zPf70NXCARYzuofiKp
9gJRu/3QfU5YTmIj+LypbMG+0UgGvxtE3Za3MPLqctkl9pLoXqQoSRhjRdrlbk3v
ibf7z5JzdT236L3n6jAFSvnyT6HTGpUjo+S8Eh5XWxLjdlz2pEfDYMEi+NhThm4E
EQixj6i7bJfNOzWDH1Czeh6qNfZSJt+iycquKdMhNAIzAc7ZtDyephGzm0kUw6f+
vLvZ6oTrVtaepqK6beWQdUNRLwqP95BzSvoU6m4UWUD9i+TRFNrPxRbREh/8uEPx
CcYSoHT4eNDITwy3ONQ2di0JnejDeVrBHqmIqfDgGPkJkVXvEe/DubTBSm0WFGU2
LYoIKHgUIGzSslIP2JmroDPwcu0WyWcPh5gFlXy+7pA5imIFMm5d7zo1hz9nI/BM
8FYTwaqsbM0QY/tjI1n2mXrnetqq/lZ8qK2bqiRujcSkE3L2CC3G3J0uskvwuz7k
skDLTfemtcP5d5IegtXfExyPxnCARMYtHah/LNecTeWZZmWCBnaqu6jCzGkN8Dlq
rOSWRL1pv98SGWEok/t5yWpMkIbr43cs4PlaeXTziwFxlSmaEo7E1FB87xXiydk9
Q+ZSZuFiCnAPuitKGG4I0abVnM2spKEG6KWzhmHUntd6KcauaYAu/JpkVFZ5M33T
Mpf28P2UPuoiQQRofyNdqWf+uTzQy6GCIK7pVAiAf9CmPffyjzt8dWL/FGzwLA5i
+oP/1bQo11lcwVZSZIZe6r0PmlSDeDqGmWf1rFgngwRQhORjYAQXNvzzj2URWqB5
j9jcvPiL+z00R1mu1cUjw+IW9brlCJlPU6TW8pNF8PMH5X0QAKp/putq+Z6FQP7y
AVBAYU3gToHPAQKWvlcVBuwSh7HZpUmKQA6b/H7IFquwjzRT8mbCPJF2iLsDM2Yv
Skib4GIWrTgdAXY9jF5gsAua31iGXEedl6cWM/MpE/6lplK1eNHbl/ZD3f8uSZaD
PcrtqcCxoeCRBC90XlhIwlq2DRc6Ezj2GodZr75mVZJvYS+CKJD2FAsuujkyvukk
OdBp5SEtdo+t/SDtxDehSyX8JSl2T4dI19fjFed14AyqLDU+a+SIQtVVfEhRP7NE
Yf9mGoLZcG735Y8tbdV/ClmjVODEImCWyjBMtd002OrkqlxViBwRkbdQNaaksCSn
ibogtOcYK98BV15G5IjcAqbOGvR1YH/vYGeQGnxHJ36o6pT5xalKZ4pR7Hw4bTqx
ZrSkkCXxo3pFZpjQtuhh+u33loVMDKQ25Emdw5LxcPM8sl2kpIrqZXR7NiYsEQ3H
HBmBYMnjTyYKHpbEgZB5JA1oeT8ahvpyqOuxRn9sByu5Q1T0dtGU0jYpDkQPnbRr
AQtR9LYLU8eiFXDse2o+HY5SL2jdJckBPzKMktvcaI2MS/jX0+auBsozWjp1cV3c
nwnewu7N2I6v2T7UtbqQbhTR2GEk/nMHSwD9ewsEtBJniuLITFwbu9ApjcFZ2cBi
r7E38Sy92+uCpTiovhP3D/jCfCKjDHGDkGmJX41A8d1kNKX1DYBmTSMZpIJw/ndW
/y8GJDI2yo/DjpRlzByD6ikQCNzHUFjaRdv+slg5lPNeF2ZFOdWTOib/6P58yi6k
AB7Y7eagRuF0gSZf9FQyz5dGEZpS5+zeEGF0MOIksi7fHyh5OpBOTR1Yzw2YDGi5
hFduxqBnjA+ON1hg8wdxsaBA1nbbHZkwLRLDMffY7aYUpTXih5MEWXgsXHuJ2a9C
TdUCajKGZ1oQNSqn3rTMm4keHU+5MHjgmWDGVUgYkkqCrFHzVwKzBG76/ukzsD71
R91QhXEDxYjoBlbDKgOW7JQiNnd+s6gigXF8fJ0jPwt3/YS5l7FgXMR8TmyoI+9Y
tjUsiqiEATWz5mhdrcm4UJsAQI3UuhlYTdJM4NDOeDd0vG3zy34JLQ8OjgFiSMdO
g6LwLPGRqa+Lo0KpuqBXC4v2/QEnoLQnW3Y3+hV5BB1/JTv6btwcdmHGvT8BujGV
o8FY/y5pQdLGwsseOh/JtpP1YnvaFLhTnjMj/jzWllJcgS/6cq2VjFC4hG2/aC2g
GFSUhTGVwoC8Y/mEVryFcp24j4IJ352MLDSrmpc9xDbKRZUCckX/hYsqpDwvckHi
y768idoNQMSzCXJPAnvcewBJTAlVfbNQFUItiK/5GJktyDQ2JEevIiVQtCSmqzAS
lkzgh2GUUJW8GrjdiksTEThgIoR26GCNkWjexofP8F/cuAlI94XyJTfvFhNdlYYK
Gq8LyT5bGa+ddW7p8dXNg2Dj723y/WfbjwOdWxv9YsAfbIhvOcHEVJcSDbGJrca5
DZ05HTxB1rp20fBzCv9LpreYRaS4QHy1qLbgj+nS8erVFgNhHqZJ22JVTWzuYL6Y
mt1T1T1JjLtpfbKWPyWNGk6Er7DhcWFwiUDweITpmdi7a9OL5C4VK3WqIO5vGw7i
mUTkIx3ACPFtO42MJGgVCnH0axekWJhpNAMgMPP9hPQVA53HLNHVesJtIU/mXfRC
paY92ybZFxpvB/FH5GLbpdKur+ps8ZHs2gvaI0bvZz/g3V/MMzzAXJpr68VOMgJm
DD8lZyrNE4s5+l/YicmMIc38sr6AWOS/4y4x/NV8ClkvpLVUnEFnlYWODYFETlrF
YkmqS/WqoyyKleMwsn6zqgr9Tv3oKCx4UYuwLJb0LgDem2yNrlzlpKkWgEykAKMl
2dfzg6sADzjLrjpaZcL2yO61d0ywWOOuk56YGNXq1MA3lWkIwE2tWSCSQRey/PbL
lvZF4ni6F4R0zrNjuucNMh2vG7znITVlTKq3Uw6aORUd20kS3eFTcCnM40i/tMpR
As38mO7B3/10qarPDseLlIO4yJkNvMildPNSKuCB8Ujarpldl2pqMYYjc4B7F8ux
T/1MDyaCkcq/hjrOIDJXks3hzRMXLw5nHV3yhwYF5SN3fL1xF5D56BzP1GulEYes
uqem3VX6JYBVp9ZaK/3hNSkDtClVPCAaxwmvTX/7u5G2AWbXKpbE35HJS/WZH/dC
0/BaoBH0AS+A/NMO+26xXqgjo/BE+xXfNqJ3UxtSabRWG8s7YPOkLdNFtNMCh6f7
0Ml8vZcXGvC9m8VI1QIV+qYtsfrcTjhmeiJ5ppbt5CzmIcdWm3Hs2U/EQ2MD77iK
vrZvG3kQNmwR7ESAcqsq5acb7rKMe+/jHQNGq0UuawXPfOkENuRTf5+/h8faqTR8
hofwqSHXc6lNoC+L/1puoOElSpFQilHgKpf6tmqoDGzZrWLNIIdgd1aHioZIS43+
wWgBWuPP/2PPBPJoyVK35eflhXVpo3sUyiOBscWx3krp5iFpfOfvD5H6MjiM7cNu
737RHvF15dzMkFQ42z9txR/vKn0h3igu8PzXFk+7/H2JfsseSPWiAmfWyx8iZFuz
fvmFFBnf+nfkdVOPUwgS0XYY8TnzPEpRS7yozQLz9lIcIPRyGbI1o4gEYJj05HUM
jWXdYmyYJkB8wXCl3asLoamAaxxlXJFtMDZGBwsVbtHyMYjEf+k+B9erynsYar9k
j4GddNziRy/Hv/tYFOjOi3Xy1brHf4TgApVP406jUmjEIl+p/sstsCnglKDIZ/Hz
QPAMqAwgTE74sW58wCSwOHvzZgj2yYnsYx8hbbDzhjvFMoekvahnMn+OEosgpsgE
yxvC/I32Sx8NhLq5VkGD7YdJIFGniq4HOLX+fZMSlwYP12eUNL0sOuqMsapr71ZL
e3W0+SbEVztNjBTht3UMSD4iNFkRpgfrbud78AQrkgLJK9wp7XB0ZcODYtTHRNw0
F4ZVz3qwzkuczapklqUz80iSYiMFGU8hX/QLI3Hm35DNAI/slIKarAzcF4U7cuoM
uKSehPD2ylfuTAvj7Qn7sbcwFVAAuZyVE3TsvP06Fr0aKbLG2VuD83/jG5oy4lvI
nN56KEy2+Kd3HOf7Nh6BmHnBYQIxhSIgN7AfM5W2yMXNJhb35LZWbyjPI2aanisC
bW7UaLtOeJkW9PXzNNZQ4rWGqAhnWtjfNNP4fSRtKKYmBBHt6sCg3KRmyikeFMCV
CgyxUaZXbsxmFHdv0AgdNpCC4B3WayKRSZUdIKEMFMgKZJGX6KFoKqLPJRa3PA3z
RYrEiyQ8dQX5YgFE1+VnWpajCYbCrc3GJwrVh2ojOp/6UjB+Ioh5r+I3X7Y5t6Te
JnfZWlTabJ33ZFCcQTPZpG+oaKbIu3ihwflp/Py7r7Ve2B50TP+XBT9CSU/Og0gZ
1gSmAo9tzk6YqJw1KteRm2LE1yJR4+rEKCjdA2hqhJhRhOgeoxzjcKW12xAqAMM/
jUMjfd4cMNOuH1hCrzh2PLEWBPZQVa3koXeXB03ETLHCnoFUHCGkEbDZsD/pFC3g
nKDpYsHEcz1isahK8p8qj+yPOHD3ioI2EIbHNl6uj0zWiU08oljqyusrjB2kcGyT
ScYDzAYuQ9uGL0gjiaslV1qkoEFCbsSD//UAinMhCquuTCHoipYn6TfvRsk94Vv5
iJog/bBsSbPw+fGsydJHvWuFtZn2QIxM8bmGBqL7LXBLsn/NvQ8ngKnNln/+mqjU
xUtb6+/nri9TfOcbzqJ5Io0ARsyjwQJRtIg0lLu3RBDgIfHk+khpe3mayrDw920j
En9NgRWwlnkRkYl0uqs0Vk7yMBHTQT/xU1LxW5nJKMZmrtfkWB6n0EQ1huUPGIfH
5mtpnU769xborexC3cwVGqhzCPWCThsbneyM5s2TkayM6mo7vbRAjnFRaQ8EMA0E
fpz44Ur6k1wAMn0Lnqpf5WVsGJO9RITzN30uG4K/0Xkvro6sgQaMV9xfsAdwdl1B
UwwRfo+3F+vJJBEP1oMZhmBX94LLCHSfFt/GX/x+H7hSygfA1BscoTSdZ+iE4F+4
+OJs2OEmQGWDOOLs3i4SVS0mvMXZyCs+a5mqiSRdlbKnv7TQPCDD1zfvwti6afqQ
5S38iH3lf6Utebp3PMyEWfBHaxGE3e7UYYX9ETOqvq86RFVCxcifYy4FBfCDvQ4c
lttPwL2MALh12ZK9+FmHGwPFxyi3M9DV58H3xZT28RY3FjA2x9datzpHmDXYb3mf
PGEc1GXgqRL6EGpWL9fZ4nG009jZZVd/cfKo+9CG+qGVDGC/bBkHBhiugfVJ9dHs
7MMjJZ/wy2/j9c2Fj+VwY1c99WILyf1vuwkMTFRGe0l6zG1GZ2VzAZm+QqbrLwZ4
7T7NLzYqh/yMCz5QTxG+VQsvDd7BykH82UN1O/1yh0zOT2YM0nBQZtEqWX1MipWc
fvK7k6dhHtrgZaQJDr3e4lJ4JyEXzIFHbHZHYjz5iD4CU1MUKKy8Ra3u2Zq1PGUb
gtJlJtZUJnexOL72wB+aAKAh1lxwMnGh/LQbjh36HbV0GJPIKZlx8uFUbcOcbvdz
G1NcbhS0n1Kogdxgzgdm/kQEpkDyMGaOOvz2705KQiLlE1FXBE6kk7yEww7dx4rw
kOOOJ/Y92bc766u/TxBvr9GHXCELxR6mGKyg6qJxv+FK3pk0bWOghaeZiN2JJuYu
UwYbZvPyu3Yiidn7n6kjWWIxiI6jwEZeTqt+wCOnvZPg5cwQtHNTotTlBlwPXgvY
wzCkdtQZpmzQk53/nDY3msQh+nBQ1lcY+gCvWqw64Q68W2O6+1855NN5Bt3fHdrw
bg0Z152CzfgzHDOZuXH6BIqnR8sb6X6KXwXz9kDCgffNF1WFUFWCSgB2nTJKuaVU
5E9B/JDOzI3qL9cRJG2hKQ/wI80dko7vEi9RM+OS2zSSvFVCGBIDmKfTcqBn7dVU
M69JQc9YBwhDaK5NKSgk7kvm+QsvpFBvDlPz13UM+Y6vcpM6XYNT49oe85C48kwH
bOkQWBoB7qQ8vlUa3aMa5JMN7eLhz+YUiU4c+T82/XzAmGIKuep4lyZ1dYJz/yVJ
q+sJzrQyVvVXXsyI7fOfSEnT3zgFygqnWllQDy7J0FQCAXkklxdktYJLpor2mq0P
COWRyZquTEHsHYcpMczGUhYqP0Lw+KJVH7ApNpY14sQ0LJN4/3q/HACfuxIyHsUv
yCi0agFZKvp8WI3pqyY22Wa3lP+RVIbCqqEZj7pWA1rNeCxr6aeNVnDLAobtDRM/
qt72OlSQz4pRohozqYmDmvQiZ/WhMxPvyNXqE0Y6yAY+EtB+bBUBdQHoFoqonfv8
pkNWlRdUkOKb4/KovF0v0yiWLFD9KscpyQXvEAEX3NSC/LHJfRF/wxNzjXLa2t09
IgFuQG2gB8m7yNanw7CwRSrOv0bBhX8qmuCvvXxabqQLN4F0wDTtJ1KO0nLsNk1g
oKK3SpwFsBHbWE0fSrP/+T0nMYxB4QF2m0RieEgvVoD/M2coY3+1SPeaoAJganhr
88uBDcz9/ervh81CnPSdsWm4EnZSZigKnBdeQm6TpjYK2nW4DYnvX2r59QVIk0a9
xbvWaOpZVuettrI7xYPX9uB90AvjS5z6hW7aMK5N9ItvEzUBZ0IN3XwHaLULmrEm
y9FFev6c0jkdDoPRAQAlh9zsFECyERFI2WPPIUwtQXHdOIdOqevt8suu+MkVbp0u
pBkYFit/IZwDO64mMu68f0L5RWxZvcBS6I/ag41IABkLLIZf5wqu0Qe9HXnsUZAe
wxQZHPl3ANBRal+3G8NpOHXUPXwY56rpJBOAKEATWeCcxhKvNgg5sEObQOKrWhjO
0A8Spo5xdJa2BdQXX6EwzZ0jrhKgwSer/uPMj6d6q5LQtAeHi40PC55eQRyK0aHp
S+wZCBqVmkzP1sXCd0tGMFMFEtVJAvcYMYMle0TJDf/ryi+CCE+1jqHVcbRCU6t/
Zi2bSWWTgP5VPwu4gmohR3dXyyAAnHInLVgX8IOgnLjTTJBIxPhJKc3Rh1pZVO6V
PcyxxTjzcdl807KYKzOfaJ9Fh7Y9EN2hNvnWgLiOe7kTAhfJngeXly3UnE1OCAvY
q30KXSVEtpBaNMMTK/oIuDELbdNPNRM9OPXFx383mp2FgWQ+a9CWPcOkg6d7Wg0p
KY1yDkUKQZsDhWh/BuqDtzXPnTwKKp8b3VTUJUt1QbFPKl5CDvAsc3aQBC8ZTF5n
gVvX9+IjlWxspFVhuwQ0gmg2kn2+sNy/NQewolHh0UrDcwNjA1vxUSmJOQa1YCwd
skcKc5p36Mzg5ubT4iEeleDPAIm/dwuqD8ayM7dv2LLa2yllVzi+BPJcNDnkLnju
8eWX+fOmQpxZIivWiaeHXTG9y8dxeo/Fg0xcztCknlRkZCNMdon13JCS2gCzT7xz
AhyQwq2QkeCIkfv2GGThxg6Wjvci4lCdYwiNxje4xBrJ8mrrQzB4uGMdH3G058ml
XK+HjEDVmzYow2w1OhiWGWWNM0fjyZULBGmKGwRR4xI4lKtnQMXsJr79rOPbJyrT
09qv3E7Bc/bcA6ZqfacFyy9+zxHZdiS+yH9zYfkM09wifsPxK/BmUtqj3d8FU3HN
09P6EXHaFzEhjvb+oQIWHanbyIXMJyivDTX+z8IM7i2xvLN9Ebm/P+KRefGAkQ6M
6G4CnGyLyl/hvFdz5c7eMbjvcDGMVNYcQTcsl/nHt4RBNqT5atXGSgKSB60pxeMa
6M8w5cYCfALbPT0RvOJsL0OMOZeIN542YUgb15o2AnOnZO/h8rSbcnk/8972b1ya
tAkXYQrkTN7Jwlx6LSm+PJNOs1tjOSjlS1iilRO+Cl42KMdPL6/fmI0c67mx09Px
MA281k+OLYYL8wk8CY6m+1PSL8hGIkAgkhnFcqGi2oPn0Brl2TKUaHB33g6Bimvh
73BHZOzIfrXlAkhIqthGZ4WTh+yz8TdPqMRBOwSaBFMQxd7/H388tHnC/TZVSwXP
0bMQy14TxpGSF7fC0qjnRS5hb+eFtMnxNJjmRkCyDelSVZIq97nuNE/i7RP21b2u
jjgAmY0hznTCujjRDjcAYLrgRz8hhOmzP57AIolIpBtGs613ULZ9ublv8xSUJThL
KNhB0SnwOprYkAI+wR3RCImh8n1KzJ9eyjQvu+4tnccf61S5U/WgP7sHvGlmtOJb
tQKLLBbPwhhSzWT3V9XCbHXDJ0JxCgOgB2iOPtqGkK2+zpgGnd6apT6Yk0ZMMfOl
CustlJ8Fl1A585roA3GJ6FSkL11An6/z2cwZ0MRGJ618No+BCD+T8fyagL98rZam
SfPocMdufK6rWyicJ+YGaiOwyvTNyPpuJpXtt6gGDaTk1xESKu4UmNG1pwJlGaFr
NH+2pPaD6XQUn7E0HbaCbxKlSa7Ig3B22D9IYzOYOJxjy6MmalNgHQdhDxCZzYLF
lw5tOBfBGwFo3eIEr8KJ2oBLiU9pgLwVF0cE4VruY4FCeyWAwRODI/AmJ8y1mHgR
V1Ds6DrLwAQrlpdd+OQAML5qTTe3AjMlKLDo6IJH2Jbytb2dWMgavj0t1Cg3Lmmb
JpfOERHVyWABg7f4XUbFYuRmlCfd0vlbZMLaE3wM4Kb6HR8LlGWAldMpuiUxA4f1
Sj3whROIXNgff3iotOdsHhU7tDmC8uiAkqo29OlgecRVw4mGL88W6iNGsG4EIyie
I8bwKZjasLFz9DkLJndzN0pvmmrMa5uU+3o81TzxAtRN4HSaLWigE7Gf3VfXAvoM
IBiW9sg1ltTu4d3iP6bBvP932/T/R+FGuFLu8BgLD/I8Jc+PGeV5twpPh1eVC1wC
KtWny1OR2HiV1BbMMkcqSeaTfCHt3v6GkT8gsusSvv6sF8rA9U74isUqvhx1qwn+
bawEhzVyPppjdKqQRrQLScLN+qkrPe6ISaRXWSu1vupdt1wbL4GQLgEZ20fXyRQB
ez0riU5aHxu7ypgE4QNiQUMmGWoozcSvuzF9Akv6uqvVcaA4lXX6ebc2x2Jcsdj1
FYN8Nvu/sEsGKp/jscwoFDbnHLv0eKZAswqghEHq9egTvx60bKMIvfd7ro9Ml4Iy
8SvOUWHCsg0Va3EZ7WcsqjZfS1uzhVWx1FHeHo3OrPCKm8Ny0DsO0KjjirurC/M7
WF4EhMC5NtfsCAhPxtVohlOXUQnPcH59Kd+KQ7H824MZFrQfa9BAtjltgbBks6dS
DRGdqOvIEl9Cfn9KsyOa0HbSjYbhXDfuxiV7TV+zvque9PrQiIzSNxSrfOunvC8x
VYxcWsKKr2Pf+ZQ/oPUsJdQ+e7yY5SMrPpL506XwXLjpab2g4DJL6ATTJ65EZToZ
G4EKoMcPMFgOhLIiFKwDQorDVHnEh1PG8OK2ixvr/9o1+oe4Y4rQt1frwQ3MGKBK
Wm+3jRnqcAHj8EuVmTr0JLoCljNe2wSBmE3rsWuryjvM6IeeKbxaJ9nvV+/JVYtk
XFX8Sur5/hGojumTIGm5KbcU7zysLlDlNZ1OW4EjZn4r8lnolVN2s8hHRQIf93e2
QmoY+noUad4jyhdRJLgcCnsMXnEBsCxU5sULQq2mROYSKh3SvC1w8kYsKSuwRGQv
+hvLKhnw830KdMeTwNaKgSqHpfp/666071cdpwYDh+Cy6YrDULGqVMuQgGUAA1Vk
k/HMh1mt94hHXvj3y8BgWwX+3ydq/pXbM1+tU1BCPNNj+zDznohMIWlVDAcX+Ivm
hK/jdHTXDdVbYNg4tomQERX9vK5MEnFuQFIjg/aDfaUdUbB/4Uy/czbB8IhyK1xE
7UW2vhDLlxhHI/oAnOl6Vy8JXxWhZAV/MzY4WbpEm0w9i8RdBS5+Wm5q968GTAMa
3NIdG9k+6zK/TT/5TTUz1JHr6LJrVnkHsb6EHbjf9ge73IZuRNPFpkfmw4yJpPVv
0LoRsB6Ax5VeZaDB7vbneB/SlPqe1WUO8IB9xld7eVp6RCG+ue9l3eaw/QPgcm/Y
aSJtSgpFwL1F0h7BmADpbGFC6RvdY3218XeLPgzgA+5L/AlYHVm49dkUsbergztt
oB8B9pq/J1g4HOSfcCOUC0W5bt2QcRhlXiLBv5AduRngYWc7oIszhQ8WHIZ3548B
qn79S8KSzCQONwSMBlhNwuISeHfagDFfPWwBELgyOunkrLAm/ZK8AQsdzgOYl+p6
576zr23n7jfNhn/FcouZIqbN9B7R5xmVrZjG81AJ2XEGl2S/Lzy5F2BU6SMFKJBL
glj0JYbsxYVL9ZGVfqO9gPY22wCS9C5/AVz0HHhTTL2dhpgaBVuow4VaVyb+liB9
G66NTiDzP2MbeDWtVAJ/Ox8AiaWdqjtI4tTfSfqr6olpVyaD7tMvfgRnXZewWoPw
cMsCMURQB0JhYrBOphvxYaPVC5zwHeFnZE9bC24bK/5LtGTsa75Ilfo3eBCAwM8W
UWtOvBbifmxhw2aZzLSYf+/GJuGrgzmzSrZCoqOkg8FEYt7UjQ74taoOEjggQMDv
DJSUYpF1EftfcyetcKfgLr+cUjXJAba8v5oZmzCWxDuSLZTs1t1OLaUguh0F/f7s
BgY4zawLkgld1Txbc9qW+L7sAcgzSUlvd7Jd1IL70XDN5GFOJdAaIFuaYOyCVJ7N
v26W7Yf7ymwByG8Vt98IMsQFotejhvWHY30NMv3jyYeNAxNnDvoClOOUhtzmNUvN
sJOcLvDMcMUd2qo1uhh9pyMMm8k6lS8H1/EVPfapVQE+7CJprFR/LNyFVHQJEyLy
KtQgRa8w/TIOWao/MU6eScLtlUpjlh6fQiOVXCe0nyidrgPLNbKC/aVjZFR6jJrE
uFhQXvwSQOlmoVX+r/OZ+qpZbbmKq+pEHRgrhKUVILWB0Yp71anOPa4Gmi1VLXAX
o5XmZ5i+zfHF/yRzNbEbgnscPRz32WXProthaWp8HETq6PGwkOAGZVCYJZ7hqIqH
l3NcaKV/djY/pSfUGUWyOFDKvf1NJ33nkiC/s9YPwQKR5nJ5ubfueRRY41avCX99
tpQJ9zx1McJOtnrvUsHASMxNEig9y9vKXGaFS3AVuQWiMKwIH12oxwNxiFdVjQAO
/tWDm6GN16lB3T30aPJiheNBbQJDWtjk1P+cE4IN0PxFFr5T1vph8BIeb70hjBiz
No20xRYfrLElg1GZ/2MH0Vn610F9s45x2uriPXjnSF4XjFqU9Rj0DgWvLTbzUj+v
AZPXJKQF7bl5Siavi69czWJe77VeU8Fk68OrR/qpNQMqnKU3r7QKDQHDAbzvfjJj
dTBtvDfbcQMFj66ufINNM4FLqqt/T+++mOLFc0rJA+FGALbd79PX3SP779KewZUB
1pGTK6w7HQRisjj2tMT4qVO4RN7Kcj7XDTGy2zNZYQDB+C+gRhghm1gUiiR2a0AE
1DKAzx9JUN+mOMPPSlqYLmBC+Z5RVEhWRACpmFN7E2QyLWEazBpGH8C90FfIEaMu
7RZHWOKeURwbb+wbX8Mz7+DvlI78Su6LNCWTs6fPpl3cj921lXsvGO4SZbSpKNmE
rq/viUz21Lshnx9G/KDGWdJhLU/h86OEO4ujmN0I97/k9P5FyUDi5h1sUnuGUwmu
JP2pmvy2al+N41tx5F7QHR1xAGA6HuwPfdpb1rY8Qk0fFZbrSmInz5c2W2TmM4iV
u2xqjv5b0//23kuXrUFCGsuDeunyIYHfJpG17g+mSvM1RIAwrKF6iMyEsr5mTQ7i
NwhjPeqvkQ7b5Pr6fsM6DI5xXaDFbA5X2DeD1XYe8LdTJk8hmDXI5ySyDdGfb+F4
JPkQkH3sExvf9+eSJKIAPi/Nk3BJByx3pUPpykbqNY696snjkbu3w9TT+QkNnoIY
WOPeCVXWyEj8dt/bC+rNFZS5PqEv+oRwYapAPcSLXRmtbzYv1lAnFxmVXeDaPBdi
6heSHSuy8XnDaafmjcp1X1YzAx2gjq5dl3NgKUHDbBp0cLc6Hr9uo8nwGWqeIDAY
ydvo3gJGeEcm94Rkiv4VMu4anaJzeVyAiCgK7yfi53V9CS++i2f2mvfz4dGVHJTu
wlCjFD+OUWNlTp9PID06zG/AevDzReblHO9aM+nK+RwfIUFKH4kef5Ks02w9yZDX
pTHpc+d+JwAKzTnR6OtTWYuoiTOBJCcyReVWc7e8eVEqvEYZ0qyrdrqJMsZ28ATY
tKJAMDL9GnldeuLCZvmGzrF5htFafZYoOCgYFJCiH9UKtRXfY9du8ba5sxci8CHG
p104GJPkv/D9QOhiwfU2G9r0ePjKXtZkWccM5OrVSvuQMG1WQJspMT2vQ8ogisMp
n6DVpGtmNf9nTR+oh4dbR6IwSdA4pt2x3k9Su+EwhjFbRokxf1nKTjhJ843Q9jVg
Wouj4n39hqWYHo6H142fJQ083DTWKg/cUk68K/cFA6w+m7on7dt6HDJHWS1ZaKhj
acrQXYrgVedIm7sNzsXFAQ3OM0oNgeGekxqCu0Cne8c2wbVRWWlqDw+drnBXN3Ov
F05KFA0XkzmFa9ZL2JMWKTGsEryxwK6dSOAwVL67Gkb+KSdvv/1mOcZfZkryTzQD
QjBVnybk2S26QxUVIATOJ4BI5n/FDXjWaj+1LZ9gvhaHubwYmNOfaYoQ9FaHsG8g
l1AsmbKMaqsWvjVaWnJnJPGlTCC+1dmeE2oIFXjLJ6yr23HZzQT6Zj4JgWqOlni3
B7tlUV4W6or7An/KwLpNBHeMy4enHDY5U9ZPuLG3VMFC8XmiknWFzykkiB5+2lVa
FZIRbN4lDThCrzwbVI6Ko/8uNggBmmB04FefJ3lXTsGCuv8l0OLxxqm/91zeiTgM
GL3MXtOPJniJUpw+NAshXwT/svCdWA+ttYIYotI9RWfpk7iPX9IJZtpM2pP98e0I
EVx+IIE8mEQwq5dqwG8GtC3XKMhDMIUzWzDJarc6hBUiRIcG+kK+3JEa4GdgkY0d
eqDqe0eR0yI8nzII+lawIcq/2WIFCRNq49UgGvgV00k3bCsVPK2Y31NbxMFe+i+J
dJTXLaurSedYp4BOUd9JCp1DRIMKNGDOKpPqQn1ZY/rVyia5aI5CeqJvfMHHYhGN
KVNVIcx75x57baF6eGKaiSSgvchcibKDFCIpmGVpl87CQFbxDlmRDo+SzwuLk/h+
29ECyFEbCmKQ4BasKeyVjujwfhsz70R/QEV99h4AZ9s6tgPngWTLmjs+Xil1sUtn
STmEGUYs8cIa8SEhiHz2io2i8TTlOVlgVX8RrUkfy+7Y+V/29n1RDfDCnwRp3CGH
j+RnZYOK7P7IQ8mIcGtPHr40t8iLVzbi1obx10mrr5ovQfffZvQRs64e3dsxHrRN
ZAWZWbKtST7cDinxt8oe6CPlzO/WxjQ5B1CCkyqOU/ucknTuH80McVjqo+YtR8/C
T2yoSlRKrQ7QYUPrkG4JSCXLeRRUFm4k0MXDXzdn8wxd7Fmn83blAeRyD6qE2Sug
n9wSK3oB+EaUrknaGKrYH/S//wnJg/88IZdZ16R6Z7RhFp+/7sueVAhfDnKcTHxU
QjoJPk0+KM6U05UGP8YYObydKHwpxQcSAt98RTbC6LjMgdmdnalupTh8skLxOMbl
o8oR7Lg3zJ6YhPNWkUzIj7BEjVHmMbgl62zuKw9kTitS1RdN69NDNoQReKS/5jJr
j8JKRu0mOPWlEJLZZi2V77dQ0BQuDRnGQ/8sNlyZwVLCqeNRP1PsWUKsqs+yEw40
1+4YL1nQOFQUIFsty83gG8DXup+sX9bDiwRygv1MLegOGCBE/A+JIFELrFBTd2AF
dqt1AVF/K89KLz6KGKUg5T0cRkC0QA9e3/5+RfgABUds/MSnoD9I6CNvPzZvEDxt
ssVyRU3lDONmlztgv2mZ3eUaXW2FcJVJaNC/n5iuy4Ax/ATNyFrNWIiR/Ek5EaO7
jaaoGqr6s2h9IWMB0qWeT/TdCuzquJUEkZw1PR/63AYYlSu2APJ2BSaXKZAa1j3h
M+lEuhGRLvTyC5BKgyLm0yOTRN2aFEfZxhyAIdhAOT0129UeX6k6YPX7r52Abz9L
PuDWJasqRtXYmk/8uR9JFkWbFLIDCnTI/euAT12Eur2BZenOOaVz+BU0klNPhd2i
34L48dwqQZjToXduZBmySZw9IdjaM8mUW7mN1c0KJ7P7eA0xvHLIfaBFayRhVZUU
Utqrv27EE4h0SDkUDHE8YvWyu0JNsgtaxMOPLRooOm42lfzi/yaYM8WszrcFh1SH
28ttmWwhC+Su9+9gUMQpDLmNervneT8+ExHw+G+9L0OrIlP/z9vuESLls2J2DcEI
6VEBuAQ75U/pKrxMRAK0/8xbPFb5wAsQd6UF+Arw8TBpZ75KT33FNuYVe+fJWqiZ
4izCCWXdHM0tB5nVSUEvOraiQ/qONrG9Q0Hm2ojd/wkXYvHzmVMyfdUn4Afe85lj
CEVBYKeFWzrjgrQfkQYZmYCNG4j4gTVZ2J1agNxfOI15OmeBb0ugTW3siVjUvLBl
B4W9iBXLg69SNdG+/LzBM0n0yer19/j2UM27B6eF9hD0KVH5Blx42Db/idgOaL6w
IDpEV5ZBTQANve20enAyyGQFe0wN0X/9uZDuTWd2QnKKAa9YNUX6dcTAQcPhpHFI
pmz6n7Im322/u4RWtfZjWPghtDNJ5sAl6o1Fixnph4gVFhV/MU5AKWneqJs3r+0A
iKFWGYt3qgd0fedFLcYiuyxJLPCGtQQ/RgsB23rFSWjGWpGMXs6/0Cu/6O8XQ9ly
TZk53j+O3iWP1uVrTupKzYLtmoPqh1/x9Ed+8oAPKni0Awfh+OzmUsiWVR0Y1l31
Y0GSBGGzfBfhv1XlKBEsdb7cDWZex3FPp22fEpWel+8eqSOWTXFLFv+C3Tk+UDVe
mtEWl8azzMorb/eZYhW6FT1zJ5+ocXhh20G9x9Y23kDLFwx8XIuvL2wSWYRorVBF
WUnjtkvSA96LCtUAZI+2zANPfrxuItcXpZjnLo0JPP1z/t4Ok1xlDgVUVhPggfrd
uOgTTfvNu8kQlh3xRIsJ/jf7hcdXVk5usO9AbgV+rKgOhCvBKXLAwlaSoO8BsQOj
Zza7umfe8gDWMNAUGw/4NPXTA5g3qV7Cx6cDOViXSpphm79iJxkSAgyDtoo505nk
XdiWMswE21fUVEbYMCHqR3Z232MjN+1APAnXnorUoTrZWQ+FPgwjZ1AzrVzztkaI
FsMtHj//dVoz7fCS914Qc9CdjU59+iJOPO9X/cZOA3qTtz1PTHpU2gwgULCIeTq9
3QFPIOenXpp1G8PUpAAUEzLEZkPiE434kCk2a2ik0wvxGgVts40rqFnp57i9ftd3
UDwYrbdN17OpFk20l2w466IfgqjZUEHaZ6rrutM+AyQpdR+WzipkK8jODKf05igW
t5H5G/DIG5tY1uiOJPVutmuKCke+XycpvI6VU/eSnX0h5Kjq3HimkJr09VgOK56G
y1AoAo8SrTJhRz7cqb0dhU6X2k4lTUA2Nrg68CGXzoLYiD3Y9wCclgMgCIuMBs+q
QAqQ9ta7otnTQxVcVGHZvO0l2R5PQlQcB4ojh/e+7WAPSn7S25JzGo4Cd1VgPTxb
eFs6iTQP2yh19QrXoEFruaad5guIv+0xTxJlahy5U1wmiULUI8mpoVpVLo09YymT
LlcwfEoQ7OSW5uVb1JJOET+CaSuLDbIL2RrD/8ZKcUYE/HzFz5MBHE/d2PAP17f6
B8chX6zzSubFst4V6V5EVQ5Y61LT+yyiR3MqehcrgOIfWV/mfJ+Eh4caScB3tS5C
QZy4FsyWlaqObQiDiQKwPmSXqYXI8MkA6rayNLVTScFkLwcJfvQ5PFg8OcyrJL3b
eIHmIZjIQ6oalpwbdcFd+aSiw/EG0u79fHrescKXk1eBbVmswz82bROYc+Mw8gy1
w2LjZgqSjZH7EqfokbjSg61z4uRYpOApguCw8PvaZ+Gtu8Obva7O9DzG5P0PY5vZ
CfoaVG22ZWR22cjvRJ2tdX8Vp1A/Uyd7GML0ZuWry5VJETtACy4VEAhiX6/eg0qh
wnL7ZkZ9ln//sHp35MqATDmVC+yelBAfZausSwNOHiAtkyDtdm46QIkAx4asTUgX
iGbyyFE/LlTfSlAC4kC6wTxqwDEQppLP1WrsU/db/1hKGVx6B9F8LtiJjYba/daU
m7B9C/WWg/RkcZB2r7fUCxALYR1jSJ6uxykObGrMgPt90fKvvtjYhRQ1vQGbh+7S
2nUHE2fBC3C7bD0JUdGvHA43u/W76xzgkIm031jYFRpF3ldkpb+jl2xUO5h6i8zI
nQN5U9stnOnuXjRCij0OJFVS61cQ6cnc4Yrqk/7gYZXjVKLJq8xal5N7RMPpLPAz
sxOOUMjaqczDJTvgPwJlhrAGGsK5+qXleUkZEyvjJDxSSQh6tVlDV52e1d5MtDC3
CURnvrJ1ene3AFPZCA6u59RjDplyoKVXQs2w1w7giRjLwdEl0o3eYG1zdqI9E0ep
PhjH9S3QKQOdb2lmvHn2I03lpUTCToPazxSBal2IXBtxRTyjA9AwuYpVm/SI385e
lHmAy90D9SUZH/eCFy1XV5FwyAA/8IRR+xrlsV/NXZI4mNIt8bc6e//z5XoVbtu5
BJ9N8BVwCpQCIHc5XkPmMKFxpZDIjaoq9ZeT6F5XRMbvtR925pbuzupH6GKPFZ5z
FvcqNrLxQc3T6+N0OrUfBB/RPev6CoiSY1wGChN5WPY5QVSb0OhZl2neU40sCaf+
grzF4oWavzgsu2U5GrP66rtMdu2U0RoCJg3wCt7ny6I7jbVYwKbaXeYFirwyO8nZ
gco9BlEuCalPtA7yjY294eLUiIoWgDIEf8Ik8WuP6hs2u+wldL55YZ/ow6CZMj4u
2dXMNoQQAfuYJOF+ZkKTBEFiecm+V5vZ28Ty38owrnX1481sZi7N/SmGGKyaJJBq
b2H5Wu9FfHwUvT8K3sM1ZR2H1AUXDUM/zAMKkMNp9OlOT0TAD84ozz/v/6sBAHLh
HvInIR8CncMUEyAFX/eQrQ/hnSgHflol44LDHEdlVygsJhaGV3HTbZuYKH7Shj4n
BzBpxSizCRRfHCxJXz1ix5hGgV7VmjmmthF8zSs6E8YnbHajxOxIL3cLcHlWXLaC
k0SMhpjnQ98d1kWhfA/HCj0S73h1aiGRZNrjwEtejQ/IxNZvL7UydJUd04YVkGfZ
pAcs7fYtvxJyAMIpcnclWgCM0enEKGXL2lS6L11xbPoqFqr29X20IsOTEuFUac+r
L7R7lnYCX3Ah86FcMVtr38qrKxYnxCiui7MDqbNXmjGwqd/tNmxyDI+/rNznAoDv
84BqSjxUTy/mBf2hdY8kwmI18lol6p8WQ3Y5PYm9ChDa/aWf+vJmA5PhgHSBWwOY
+jjiS/gYmmcFqlIUzb5cUmw9NBJVYrcvECtu+pKqbOFiRnFqBNlxGLjqbWMbq5ZJ
mqSuKAzywhJKhrmp4v4BZWAN0cQ4hGUygpk+MDfl2peXS1yXsKj6tCavTrv84w3E
q8+iZVRp4NRczdb9ft+f06U5Gdi0fFB/744fBlD9QykGf8237WKCwln2JX3vUc40
VzkdT04vGrncT2tZ68mvwKjmj9SZpou7GikWz0DcX0uKHBY0iTvKG4fETDcNq7Tj
E/5yK9fH3JHnV5tUACux+kcoH9KMRA/xXYKLNseoTy2obF8/4frUL8XTcRYsQvI/
bReeZRsZ3PB2sDFmu/DktB6E2PmiodH2RmiubJR1osKLUoiv/lt6XUla1HBXo0lX
qNOhprfCGjvi9BlsaNXGWyoDBI1sRKXnG9rwTeu+YJbbBo16MuWkNhY3IszSwo9Q
KjtySjX0e3pXipfGopnd7LZ07ejhfiVx70dX1EtCB3jUlnuSkM+IRbvWlmFplhz0
0p2L0Ab9DuTVgsaJ98O2UFDlAOckHXmX5TH6GXJkMEqfEypr4dv7a58bEdE6UQ6u
0mjP/73zA5ao9THh8MrvWjJ/ifiMig9AQKcwMh99t6Zp+K0o2Ya77iJUTnOjfBRn
Hs9QANcbjVAIy4HjyjD6jXSeF/n3oR42UJzdorB1dJDaiINNZHLiwIugY3GgQJNR
p63HneQANo3mdKaUZU4AGbYcEaszY8OqppdWQa6pqc90LIKCchZsbDxleIHtrX43
FP3ZanHTWa7pq7SZ2DKtMo1F3hYC6BTaDhd1EesYT2slcOX+LQtxey1UD2gzPfL+
HCJwDZjQt72Wf0X7kQA/VSQsCz3wQ/ewGoeytY3gz8oh7lJH+B45NeSNfOz6UKQz
jcMq9kkhg3fYOdghFEytb0UW681LSGL1reQ+QIf6o8UY2K9lmSSGw6tFSHQ6Yicy
8aLZTs8F+zS9qIKtnM/BP8xMqGRNPIJNFZcDxj2slQ1SrZNd5eOyGAJOTih0+U59
Fv+PVGFauBT6WN6EvdFrUKWg9p9TCVjlyqkum+g1Z+nhnRHVxPAnPF3dYSBnFkpt
cYNWhk5pKjHY6iHLnxXA29YjXitOlwRiD7LouD94UxKQ6Jse/iZGMfWUREZhIgU/
L16X6MXX3iXzcOOeDuovFNl9qOZ85mck5GGGIG9QFFv7GwKLTL3ko2Ev1yTjYb4k
Zu3UVWk1WIYiS7bOYaQ7MLlVVNoCc20PgwROofxbRrXMdz9AsNiQortAAeAn/04w
BJXKC787tfcFhbdpx8QzLcZV2CyI2HigLFqYLNyuF4A7OqgP4px5yllZpWJKqpwz
9Vrj50dVq8LHWtPWkkesRS11itgHrhnNvMHptvVMXaskGGIIWwfPvKC+U0n7uQ3E
9ZdVsiLaWGXDRk9Qdj5sEYoB69fex7xAl3yoez5mQmS0+oh9GgDN7hhnsezJt79f
muP5N8m1/TQTqSvViETe8qyKV7z+bMeEH0YWkY4UPU1smBKHIPUNHu4V/InJGBtA
NA1Nfm130QWSDpX6JTeKuXv3pGkByfZVgTEl/CNVrPCrpcSioNAhy5qpcbrJr8f5
8zrzvedp0n8zvsX9KNPXBncCCrNIBiXwXt2AornljlE28ZJI16BGhZkDZXUJCUiX
y4lZZwDGDuT0oPCbS33swWf+l+7/Knf6pl0wiwyLVSSyKjE6LNNKgX/bEakGmpgP
VJ20mMB0xsc/7QEukqIR/uj8/pm53wkEF19UUrkXEdZNnDjeWrOj4RhTp5ZIv1LZ
js/GCMhYbLbQODLWZuOQs84mFpQWxfyDlyJqsM1My2YQDPysiVmsnWhLkfMSqjtD
KS9sjcEjPcdD32DBi/5Zd6F5FTsQzptkMb2sHZaScU8bvIQ2tueCLIdjijLIytOW
CbxTXNcomaF/ISwC85OGJZKpACgLBPfyV1AoJmd8KB/LKhpgp5yPAPqzL2IIk1Td
4NA0CLiE5mkX+V93NiEBR/2r8rsSgUI0XixjY/o14DNRUbjQgc5DPl69dOx4Gdv4
95TIhiGAu0544WcVcLlgIW0KlezHdMbBydjU8G4jqxrGhanXek+/vWryc3/q7wtS
x/3TxRRuNVb6tDVCUM37FfrCWmFMZSDX5ORszVcRZSBUnMVGjXdGZMcnuEOzkkgg
ez8AMFEiDY682fhV4GIQ7Lejw/IXriEESp2lwJRn2EXUXXH9PjCGJsORnLoqDn1O
/bFptM5e9zw7+CXHII5pahQ5JnIshhDcXk1+DM1scK5OPKYuvI8tqBnwDBRh1nHU
tcj6ZcaW90uSz5PhwN+AxfwoPMYwhkSl0NzqFjbnauQSjXs9e+fdzDCFzgFMN9/h
tGYaZNMCgHexCbR99yR1Yl05iKHVA2AdgcunIIkwGvLFjervxhw618OtKFF5FZUd
ab4p1FTdHNuFw+zkSFfgV3mhdJIkCxGC9jIEfcuaYpV9v6kmFOoYWuv8/yIx+BpO
7l4Y+GVDGAgEhcvoBWI4/A9oo8q79/TtmruJCL8GaORrEwqsROa8YPBR7WsJ1Or5
Qoum3K6QM8AAEsde/tqnkGHblgSW2FqDPgY15/aLxnu/iFAoiSUUYuODCGkB0Ivj
U/FMsjoUrMrU7l7aHXO7FtEYxvcVhNermbD8YBOrP5Db9aE5TLWpoPExiGRPrqQs
kciM4fyZpL21CHYqG3RdSZ5OezUuVkkbzVWswpmXPDfQsKY/61v9BOselHXt0BXR
Vf9L00v40vPbvhwlJqEixdWr4nrNrgodDU63AXnGzXZSVYNQAKlVmffaT/wP7Y2c
WeuipruDR7Xx7eKrCaObuVNPKLBXhccXkkpBkU8ayWi9CIonCpXt7q0lDAtc6Xm0
+oVDC8vsu9Ct1ZPAqmKqOI7oJH8YP5NQrsXbXkt7tOl/WakhxYrNqot6enuG6LPx
FG26dp9ewgM9U3fsvW7vk0DC5vbrKsV0BVptroCBd3ywfAc4GfiMr6VJbRpcotcr
vjNO31PLt4uJMaoZzdj50l7gqEXo9K6kL/WFb1xH5FgfiDCarRzh0FaxPndwh8sx
2RcoLVDBRsa2rCTv92FrV4FUqJwKTxtRdnNuyKY12uUPVvQk3k2oUG9+X5aGO7gW
aszbsssmf2HF/H3Xqc03SBmqQvl3noX6hC4TDPnsWYD8bTkm1LszEhkHF3VVr7TT
UI0A2zYipuxnD+Qzbn7bdgjv0MjR10QCr99BbDdb+x2zeyKNL0ntGjMrv0ktzd1t
tTB134WmBSjH67avkOXWaWQyYe2FQThCdGIk5KsObWyX9NdbofWjiw9Y1SgYDm6A
BWyivcBRGhbntQacdDN6uHMUsEAbJm2I9MAp8bmNPrTDNm/QZ9sEXfKiWboPyEXb
NLQLVVXXsvluVfB7uMklsef00u2zGCXplY2poaaeRMwE+ZmModwcO/VnRtuE+VLk
SF/NMxB8NPN8EEVQ60WPzOv2Q/ca7bj/2Mc1K6bG2KkHQikFZlQjYX4I416x9LDl
Vjbq6Hob+FIyoA+d8w+zX5gCFlwFzH9ZPxOkXkMbiUOsaXPYOr4UN56sQ3lVPG0d
Fzntd/4uf8NbcLZ1y+yXldyK6zZtUjYZLPplRSh5sALyPjIcRXht6sCBA57KP1rl
EXQ17f4sLraskiUELr7yVlwvfrn3EZmd9qxaSdNKYkMqnz3fsEm7DzyFPE86w/t4
tZ2rNDM37E4lHrepy5yvGHRnFXbdgPpFTkWj5CVrZr1mtgULw/fG5DuII8IxcElQ
z3K4Zo5L0hUZTS1sTrJWZVsO6AwzsSi28+RFsm5P9bFs+qZlMkN40DBXfu1fe2/r
SlQW9ByjU691ODqLSues/KaWrGIf1F9J7OuxL/PHO6Oej/ouA0umVCg+qM8/BOWt
c5yubzRg/iQ1ZTUfwE/7oieBmZTpOx7H1opByZRXEVqwuXosVwcVjnNdEiXhcu7D
Mue1ytzjnAzWpdCXHlXHbu2ZCWQPtZiTO8maoWz3nWVN87H/BmmVXLY8c0WPdMP/
wOBkpZIwvVgcbmucc17Q9a8s88Y+eOc8xHE4p4x8NcKxllqZczLQmg3qI4KsEGqG
DgneL+cQCVR9e20Szn+JgiGS1TtNZSYSXAOcryzyLKFv0DpaLyqp9r+Q6nYd3NiP
4Pbi2Qa4xb+bIhKHpblnEzk5UH1avRsGkagKCjP0TC/YW3yzj30KMs6z1yJgQ9gW
7s7RpoNcx8SQhOFU5ZUA4XMBCQxPxZpxTzxk1wwVXOSV2MX6849BmS1tU0Yuf+dy
huUWU1pV9cpV8fGkVojq9ciftJRqoHdfeLiyYY8nILgRl/CkRzm/8IFMoV6DY2OF
DQp0U3OHi3pYJHN6naiF+k2MsZ9FpffDRcUlobJgXTAybHAJz4ZWYDyGKn48GGT5
IFpjinxIc0rY+2Afva97wMTr13O64ghwNOzrXECeIvblyx3DACtvSXRGFZsG8pm8
uc2F+pxQvXwMgAagpkrLypkFUbFKPLYf8/Ttlx1+BWc8nh19gLiNKmg0kd85pKrZ
yEjuGCVgmNXOibOJA/vRWSg8QZKWvBbexUSfiRPK5Qt6x2Dm8p35z4rlMOXvmaTx
nBnvRvJEjtccIU10JZ/jOXEbrqxRDmXhMLkgRcXRI2yMuTYE4K3LpNkRYwPVi367
lQXPdB++wUkZ2yATKddUm8n8AWnYSXNSCgGYVdQoMUbWaro+DW2tOn2LUBjYGhl+
7i476yAzd/quiFrvDEvQPiOdmCurg+MMAcwuke0sCjozDJOysn7h4qHJsQBQsppR
0E5ST5xzoIrmdhzWZkW/+tmsq+t9dWV44gCvlrevqQyaWasG0gWGQvwUo/UviDr8
wNDZ2TpjxiTP/pqtZC2nMb9mbgxNM19GUUvnd4J7Ga0RLEf6aNldF09NXIl1RknZ
nYOnTyo0mxm/Y/3C33frQ6GKT8xC+cQSQzBnVNBOBsvPPtgA+Hc9RIkwv92yRZpw
5n9bUS6tXZjogOBtA7Ff7ILc5Sm09YMLyoICWWvSpjsgnOYRKv/plyVkQI7EqWVb
v1oysXTw8BVHttMCmUMuGLKHiwVmqj6M6NiezfLAYFANnHRChivKqnBry8afWHRG
iEzIiAiNVW+8/ENajkOxtUEDRGhmwGJWeJCUtuTn8mVZoNZGIViZ4TJNL1ws5G83
DvlL6kjZKb9TPK5Dmy9XJ2VsyBZ/l0cRXhTm0x9le6OqWzNzlVWkqcaL8LMhHBOg
0VO5IoAdFrpkx3biR2+Be4G2ebTgRPQ2zupYd8dpt82ZBeyBLQIkhCW4uu+eOLmO
4UXVr11xgBQVcgJ84J8OLvtv8ZGpHVOcqZvpst3OzrDR/kAHXHVQpg1Z7y2IpGhl
BRUUSzb6zDbZL1JpQDtBwt6mGKMHSoFWLDqCRFk1rsGpSjN/XYvw21koQ1dNndCR
DzZZk6fjCKDxcSV/W+/buxz7PJ6TlekjILJLegg9ugfZY4g+io3F3/pmnnrz2mjN
siiRGfKx7Hp3sld8E/3AiEKaMtrk/LNWgqlFo/ago1QV83ANoExL6AxlZFPW73DL
YJiLfbxFJRsJ9GotKYaX5owINvkqEp8DljuykrNohMcZxRvDxKqDbHxtAsbcXP4n
1eGkC8k1h8/C+3h5zXE/Buh8jxnC8w9ojwwSS/gFOal1ztkT9nUp093NYk4/j66X
iFQGR8rqWYliiEQU8Fp+zZ/UTyH6HIJhB9PKA1XXgFZSwQ0nWUJU93RATPJWQ5re
I340+YHuVyunSWVsmWwd4miFPhOtukc8SnVRaGrqNnA4NiIjLc1A10ya1tHS1RQ9
duMgfFLTfZwZTExtNza5waYeOR+TcFN7/xYBwqV0RGGkk5uZuTEbjEAcU/E2wpPE
gEuL13e84ReaWNPgf6MQ4VlFwnxAXmE04W+9sH0r42vnJbsx0dC/RTYT2B7t5vvT
zL1jknh+Ntqk5D5WHwEDOnLy0suWmc7tj5hGd9dUBw4BuhyrFaiD//19ghjOU5wP
BppkojXqsDJVBDf2CsmOn9M9+fey0Buau8ISK6VGuGF/cdiWG0un64VPY46X6Jkh
HnlQQtH/6hMY9/xO0rBv1F+Q+AdOYcaBG8v4mmuqxwCde+M3x/ktgHct3a64+o3P
kPdg4cb3uWTX9y96hWGIp+0PfAJOTj4pITIdTaThrcGn/AwB1d6XV8jDqidW+FDn
KrjS62mcblbqmoAPik67uXoBmql1UjijWI7DWg+0UFmGLvuIjpOAGmf7iJmL0ClY
iPLjDizhNCzxlh8A+JkmHgpEJ2RBA491NhC61hqamlOSkUHZBemlh1K9AomQx5DT
Y6xk8nJxSMYHgS6GzwY2H16gOrb0UnqQo5uoJPRrXdwrwW46reI5r5kCii/DcDJy
wMVP63JaKJX9vINgD6xEdzAfXiQCcY+s8mFUNvjRufUZ1cMSwy9FXqeEQOO8k1aH
f4xdm0N1jGT2T/A/JVoXPPS04HYl4hI3hI52koDHKsvmNxWp1XFPUG8rOU+/+Mi0
ll7wBWHx2v/wIApB35APlQLzojkys+IyIOtPIOe09qy+DJWmPLMcBQideUZ3dYox
HG5HuyKk93nugOXDjMGpBPhD2UXbQzdczAz83RhIkVFOExnRrPsP+qZFC9O29Juz
owWXg6n88ttWFXHG+OrtO08R3Ezu0xbxC0ErUecPKZmWPBJ52Y/C/4n68agQriWf
oE3IEOHDFzPid1dB0da5SGgSnrKAGwfSwRCpOPB2GxXuqINjxAaJhIzd3Pxq04Y6
TzIBVqeqvZPnK0/rlngwaY4jt2CmJNPrtT/XDHNFGlRbgLAnVWQvc6jNpCJC0+W+
kLgQkUj/CP3h4mWGNRiq7qYTtZbeSuY+MXNFIvt6sJtJtLu8YGoxTKESvWgzO+8G
mLQ83NxyPmgSVQqrTa07itLdGQyg8IeblTS1Jnk6oncQdGf1XqX6Axf6fS3xyxDz
7Gr2XzgmhnT/D0amqII4PhNfZ1dgvIt0sOK96RHBfl06JyMYfYGZVN41z6FNdzi6
tFN37KGZU1Omm0cGN5dqFxfKduka5zhnVz9oTVzCfCaSdQEMdIf83SazQqQ58PkL
ZYd9z1Y0ZTQErDenSXB25551SrKyQ+vPeBrBT7V+7srb4X8lFRZdCHWNYBafS1ft
SPBvM9TALHx62dGSB9LisuQ2iGysr68faWasoR5rDcZpCGPF2M/YC2a3AcExRzD6
RAvzttF3s6Mhwq32PT8cK/XEudPOwJ/1cXwnMx1F1ahZKVdRwAUfl0cVOyiJ5WDO
WuMTLdleGp+ftrnKSTavGmS5tbn4E0XQzWv7sPYmFKk4ud2OoHgoouOqbmp6M/TQ
rqVQEfY3tZZ7kZYUqUo3o0Y6G0CvfRFmLXNmlykLhhfSzstjmKfrkub5wyd0cJ3n
arnIomJqj8togXnsaeH0y0T5W47achzOCWokM0iArNQ3+UMV7ajRFp9Wh68I1qQO
mB0zWh1fDxcYEQi9EBpD//9vIYLvyDRBApACEL6B2KTP2SjmOL7xdmRqqiPmfS6w
kQU8Qg7h+6Z/YHKpHwjGu1ZXZSjz1PtY9qO/1Dj0H0R8q+YAdTgaPxkRj+WuZ3xU
ywRMqr/13RG3kwXGskk9CGDDS9K1wvUktT8p5JsnO3c3sXqEAfdk7xeTSfvQgJRJ
K+bjARyBr8mE5r2KYNGpZn3gG2wTEm/+4OG6yk5eHgi+qIyHPdEG7Cokf3RVkwD6
2t4DJOPrdoWhSZluXmEoksThlti2miFhOEStHDoUYVk1zQT1AoLO+q9u98HmsKjC
woDF8yvPfxrMbaJ+sbkCXvJR96jM+qAIxXT4PY/86vSFUKZNufChojtWKexgNlwD
jVGOEWg0gPU7cdtIMp8jpvnJnt066YtlxSq8MsyzOUjZ1Q8wPCHwUphQeblWOTC0
nrO2YtKFMPZsQASjn61gwNc4pLK8l41eJg51iglcVKoqzTuEFc0XfMDCJuR4lLs8
uhTtIecMstlonJ94trLNXkyMsRWEX2udlBDg55j6L86LzjRoCopNjoKY0IVTt6tG
tKFhQyVr6J0vJcPstS0Y9yBDqtkpVvC7EGojOWNdANw/nn1YnhzJTp3YjnTKz3AE
kJkr+sqZI5J0jw523/nrD7bT6uZ63QrdAjGqB0BCGdAYEzyLMrDisfxZJETAy88A
jSznV1HrVjq4lz0+o9VQQAYW8sLJirLADKoWm3WwrcGgCweTIJagidO8h5rMpSPH
OeJIUrV2Yds8gsF0vVh4rVz3pMK4lDtBPOAm4uq2glnEJXSvKAijm8dgdt+KgVNo
hpGxZTD+r1kEJg30e1n59ac5PKKOdU3r/kAYnfssrETGxhmMytwlPmlIckGXBN4g
0UGV9Kzn7zasPCAgrd+isNrL06EXlfVM0XbEUwP+oYLn1lF/Fej7cAISvTq15lcK
Nf8Naa/zxhYqEIHXO3XrkU/NJJQ80xfAURsGLkMKDFe3vCvzNVfZ8eA6euISi4I6
jeV9xnuxINSf89HPsj7NN+uDkMVg7Xbn+ykou2uwUy/O54QbywVEpwfk97Zv5I9O
jgcHiFksykhCOEhfo0qC5FX1KOI/2d4U0vrlYpXVmDOQnwiUPLDRGXBzzck24P9a
yiFp7tJ0gyB+xisSrecJh+TYpitUaOTengPi+lGG+q2KATLFDKzwtyJ61BnqM3A5
Zc7zB4QlOj2vS41DJ/kuoPFhFFEb8VUKHRWx+l10LcfMcPqf6t9hhX3TQvJRxo3I
CIMvzKtyzzRjTW5iQKi/zGbWTwf0HfnTkfm9mQo/YQSVZTPIHkvdmNeCSVbU6Qr0
nPjX26LQ74zXEvpY/bJj8AsLIF7b7aEEfqSlZhIMsjhIdnb5CMx/NVJvniI9RInT
4DCS+T8TEtkAJJKcRncXjA1qPkFZrlB97oKbaRp4cNUVSkpPpA6XvpSRoKEf85We
1vMW2+1KxhcWFt5XlcRgnDfPylLi70ykveEt2tetpD9TnxcZIYNos1Vs0RcMxneO
Xwey1GLirGLT1oex/C+j229JG/66AeJPMaR3DZQr7rJoPuuI7MUwnRDqr9AihhL9
ovcdcTBPrPS4wVK2/i1vahcTyWXPifNL/I5GmpfbJEPCkZpuT1WstKGRRkBgcF9b
8nE6AWQF2NVzpdm4iuU3YYww9+knSG/uJDhEQLV8Fl4Re0RcSeNFGCFzU6WSWH5b
zoyUHaGmBbzHDxEYEvnIVf5y8+1Je5EmUp0ye+sRitj8jvForwrohWOgmt9neJae
3WgshATt8QcKIEQLPB9LhoXyENyMXnjS2eTgfs5d9FzDyh9De2FGlzqp9uKLto3j
8YMs+re2F62xyx3Fp7nau0PBFdx/xJx032gQ16u4w4I9EvnzVWy9vrgJ9cUagntV
cxaiN0is3RCQmRLG1tZbJysNT5Zi9JHoBr7j+YjtbDWSysXff4JdPnOn98S50nsN
z0RpfYMuIp8riqhxvBeNlHN6QEvjhdzVacAsFGOWhCF1mLGlNgxhMHfYq30mkJl2
vybpIzFH4updHVRTqExEWkr7ETjx9l4YW5DHu/EJVgUIXwIE9pkFlnKv+U1nQA8w
KmUn1QtfGRPbIZqBIhIbpm8B6uGuHUrjPw8ZMopHvlWNycf8RO/Nz/AeHLQmOPNg
Fy80PdHsWS8k05tsLVMSelZNhdbuhR6WOxr9KwBWfmduKPRU6VjCBXNkGWh19n9p
YYd020+0hY0iKdj3YZhm+MeSN0RCYCKsZpyNIABX2BnUGw9Wse2xDKYSNvedy1XS
AVlYCABL9uKruZCK9mmndiJbttXA6EN7vpPUNVdVPwf6L/Ydz2oH8FekUVNgd7rL
iUk3CYc7NTofHhRSIoeqRw4e6ffiwVdq+KoFBK2f/SobW9a5V9//omXcQ1poOwT6
5f9KNpaSPwXLa8TESODAGd3BznSkV4LDF5tgzkyM24mcEimq0sMmnLBn1BoTUhNa
sbUpTqNmcGqfC8MRMCEARMbdjIwlYa/L8RFuHBT2nMMSwK1R2Dd5xoXL0LkZXBTJ
Ns0QAdAdd3LvNw2hw5jEKSlOYzjgtHwulT7pL3vYeYg0A4KWzmObB6lvFDzBs1rM
CXQgbmxDeuvmyBIGemPNFGMGlAybNBur+IbbRpaO1IRzvMnbrCie6B+Jt2oil+KW
40wqARje3RVt0Pu27i+2YLifFfnpjDWR9cbhXMM/m48LBsszbb3sdvsxDF5oGQyD
5Czk78riAtGucvvibVLbGKHgzf6PDRrIy2rlYAG67p8Uz0ubNL8SHJnnlJmh7c+O
qe6OaYzyAph3Orc2+WuxE2S+xBhb1ObZ4sEG816ErHG3MU91wo56hU0fcv9apAM+
6j6zVOt5RFnlO723CqX5C5XgvwVecEzWdWoUknSEq4OSbDYNw9dVJPAJd4KU2cqo
0ge/3TXQIoinE9ZFPlvzsK4WCo0NfWwB1Ew1KgyBHj9/XsZRF/V1CLcW+2sP8/Kk
IA9Qn4S7C4nx2t0DSqDnBVYje3okOqLDULlnzbbyyUkKfXoT4IBQZjEIUUnySag6
7Ecbi38YOv/fDoEHo5HS/Ffu2O6ViXulT69ykiw70WeX2tWzQHogR5dcXo6ak+RA
RVkjnC3uJt69eTYzgyviGUgWKj/q84nbelqNYzYZXsPaGRfb14HN7xn7bv/UEMdx
quJrDy9T05cj4776pE/SEs08wgWnNbOkVzGaueLIE6xluhMCNeVGsZyF4A44A22a
E6n+bByfM1qyUkHK9NocpwCF/sP1wEg4dQRaTA8v810Ur7mFPMJ88U88BWT5DxwS
Uz/mV1mLky9UZnvrHXA6/6CLgRON0jAGNFEzkaAkY9f21I+BDx0aqeoAILrz/bJr
9NEmGlwSkoqm2hvBvjZK8PvQtdNgmr8MeH/0MjTCCRAthzNR/A/2+NJcpuYQtLdc
0Ikp6A7oR0k2zPfRZN7xONsIf8xlK+mFqYMoIxJxfVQgr0pw7EOsStB1o4jdfMFu
4E+TjxOj/UM2kim+KFHUIlTBWwE7ARn2sU6VQjEUSlU+Wj/PdWf9SlnUr2vchXAd
QybE0O5tLtmi+z9iQtuR5cUTpzXtsbS/65Z+uPbDSPu03WdEvX+tenWOZxaOU4ex
lqkmvNdd2nyy1xfkCXI0ur5zZHAm8RA3jsqQXkOkI5hpKmVV8dPdIn6SWPKMo08q
XGzY3icwtSG40AI3Qo1us6fFC2lHUNSJX2lhuTIwchVlF8WBeJzGJhAFLm/gyIx6
Kb9sBK2h4TwT0+EpmRYanuFJdByLujjXfMP3gIz9PE9XZE39ApyVbELUQJXiiZ+m
7b8ko3Gk9Fcfah8UhvsPxnHEXljj6F4M0CyVdSzRlrcyVt2faNVnFk+gejeXBzEx
cCyaeHbPGpEOc0UnMMTlJxy9uPvkYxmGVoB4/FfKiKlHKPl21b3RZCakvROnpfYN
BOHvy/Uw4A1YC1XSNuC6rEGhTaA8lNi9d/tbx6xpy7pzqb5PU4dUWVCCHj0KzCsB
4chnbd2+2RpOXBsP7sQrqKouh2sZmAoPcZYDf9voWmA7cMonBU6Jvnc+aIEW/n1q
KY/ald7hOntNuDo4qnqlAink1zBWMgMWVDicyMPP4mIOjIy1UkIkspnk6dOedhar
iRSXz/BwmkQo1vuvpiGCA3S7WimOIMgxZhaT6ROOBJckXSZOAqFWoIM2hAHEiYvo
P0uSu4pmHWsp+FI0DqfOg3kIkwpihDuLHldI9NRJg0LGDsu+J/6XDFq7kX40X4Sh
PGIJ6aOfC5OWt/9jeRrwdDE+1qaHzbABNhkjzVmOpJU8n3qzcFNKd5pspjoNP5Db
EPBlMwjMTgkzPmXnqXzT+goPaD9ockhVi02fnL7DVCXEMFWqLWWcsJhzIYOSQFrr
gwi7dCCRX3UgpwgNJvi7il6lAvOeBqoklPCK6U6DCCN62TD9qabcBNV3qZdI3KxT
hWaz9kJ7M8c2XTQZgKOHKaJ9afgOIsVNel2p5samHP+MP3IE/K+0MYYn7ps5QC9M
3LkgMu8wD/W7fnaNj51ZkLd5L9yhhr6dVztXQb+tpNIGLAJtFHi+RCvuxbkTfvZJ
S48gc/QCIG21cPMVzDLQoQRHOY+oHY80bsHhc/L/tt1NBy9uDMnJ+ReWPKHi20fR
r9zzPJSS0UY3Io0b/ORgnjD99sLYYts3O/jnDHn6yTondyk4aN3Qe7hhIrYh292F
sU/zCS1SeFofHO108bkTd6TTX6g/vQhFy4LxbRcEXDnjJ9K6I0mHK94ShJWuhdCA
zO4jFXBBkWNYX40L710T+TTsTfIegSfMLduKkLT6dFo3S8qUAy/supF2bu4rdPts
0R7rI4kQat7MTzekqo17JhZHOg6kWHTHqDjEGWUkfjamocxfasAAlU0W5Eh77dV2
1syLTglXs5jBfjsZLvkMGkojScYS4rBdV1eLGNJR86Fjkk30hiwxS/2UZ8b+bOvD
KPlLDH9bFyTVgEMFh55Xkz+MMYly3GxauPFvyXnZLjtrLAWD9S81ujzA+4SbhVRn
I2TdcCyfj3wvT1rWQOeVW4n7dpK8Lzc+xCbHGlHximetF0y22rmR95sSpz2ta+6w
lniCY01Ec5ocAvksD5gbzDu1lCkd0tXRcomhsPk9rMAZz8nCK+jTTXHYPLaSFQ6z
o7+4pMpDSJjGmLxH1PawSP/9PGZpIgK1IlHNb/7qjKkSoJfHA2O5v2xBlUC0uLfq
ZOU5oY5ZPg6qpoRSmfNb6k+Bkp4lmNsQmzOcxsloz9omQEUMDiijUbV7efxYZVpP
/3D6YtVfZWka1Pd3rHqy3TeBZbasUu9jUEB96tWBupXhlb9qRDl8H8LV0VfD0ZkT
e6FeX+T1fnULoLkBwr/DfzOeBEDkmbzYBvwM5b7c58vWxDbpLltyACG7C5/Meof8
ucGyHibBE+J9La9R5kd0MD5Gu8kVGttB8plfQBXt+3pGExECmKTrGRvMDqdCH8se
nodWmi4JLyPkA4fkdBx0PKq5Or51YEDFE3mMz2Vc1Ri9viy1Kf5RmqVg1gw2Ic7J
DLzw906ImgtUD/Oq/Tg0CB3wm+Ktt+E2OACfaTrUYq02PhThPLgclgd5cFBU0TxL
R9G8JmVaqMYGKI9yk3nUdqpQqEKK5pX+HhOzwO0bv2hhz5go03v9vWqJfI5xESJK
aCRAQ/Yz1lxuuzCvorMn4spKdJR1uII/wl3ubqGyC2DVXVf3XyDVoCOBGOr3DOCn
fHbStqdy+3SaE5g4PIZG9VygYW8stz/fHdCRAHF0v3uJbELyOfrtS5M3HX6frfxQ
bwyB1b8SgbFTXa+XoVAISg1An2wWWWLNANWzRIGergNksO8PFuOLtDkgKyJnyiwh
JZFdZNtX3Sd86xBCI/FLPKLuW8l2d6nsFabMQeHbYLc5v5RfhgmdOH96gC6CONMQ
HX1de5pgOV7bZ4Y+BAZehYDwfGDQQks3fFzARRsgGxSIETfut7Vg/J8uMLokgCaF
GoOWp1wDWNOp0UudmldG0yOb3xPl8ogc5BRp1C1XxXSLkb3D/6dMCotPcegn0fIV
6L9sWOuqbpVdVuvJy1T+eJ4FoCoEoGNlf89pyHqCp0hhmpUYaftp4uY9/VZ8xTO/
VVwxWN+mAoIZAaYTPSvHzL1/iQxr9QhAwBq/wGlbeg57zn0UV8+gstWllo2CCLUW
KdZo6rbzODCbJvrpbHWVIhLtt0qgypGnm7/T2bkokdOGOs64ntVEBouQXny4dTkN
FOmOaKEM/4sqoDYhXBGHu7v8c0IXKo/frR9AGTPxiy1tujQ8wRg69oJ31HY4oxp8
SEEGSXNm2CsZL7ACLbS+41S0tXei3YQzMkQtjFl4i5Pf9ipTtlB5GnzZNZkZhK2k
HCK6MLuGS7vyfbK8XXvjCZpiGtdrJquf/Nf6GOOyUBFY/xBYe7vZSpj2m6gxUJQ5
3F0RsrMbo1HxYTDBkGbLNtVb05ICUmMfYcfm/GZBH5k7VrAcF593myRdhpLn43BX
m1wsuj7isLq5ZzSC8scHl3KTmlDGNAhfIvP3rdBT2/YE62JU+UrzL21xqf/LFiw1
4An5GNlAVHhYZyBbbW/YqbS3s8JxnLo0JMgJS59Y/9SdtvMBbJof7nV5+xEy5Iur
/cVfa5G1L4kUvziAx+11lM0z3DW+gFKX90ZDhvIAC4V4yfwMDFHNOTpYxq8pKDDq
SplTfyFnWFRQtqhLN+RVWZxrhN+Ck7kVnuBEyQ5uTbnHPQQLJEjhMJBomWEt3MDZ
s+IjkzqseBHyypaxjRVXRz79ue6AmmVtyujXXUW2sAQ+T+B5E0aVQM1v+0KeHEuv
ZTRimqwxIzuR4i2RZ90yxoDr5DlOPG3Z0DllVFIp8ippUtbgGtpT3ry+tu4gXKYu
3jULfGW0Nesekj0gbS21R2ZipA5W3x/78VAKvKeKvxK694VWeb25ifcPg8hRw7wv
q8Qwika+wbpeYoOpxhVhw96FuXPYnbMj3ZzTBrwovKDnh3qWgOPq6/dsqCdRg6r6
wlGrrK6ssY7NLF3FYzY7r+SbeJkKaHyq8sU2aKU+A+Bx7Bnlq9Ghe1eus9EM7gPw
M9h9OsSo6NP3vecR5E7Wt6RAHnYq0bNJEoOWTJt9OaAtYWh+y8izDubQ7qA3WBpM
HmmRlEo40zbMuWu12x57kyUfqqbV7TLBr3SaDQa0mStryToBdu8AIP0ZJAb7Qpf8
rbHiH3ZrrJD0Vk8utzQPLTpHQQUNTj6I1ZMwwY5v974NGbss2yxEddZJo+8nZ4JP
PC8o08ZfwmDg5vz4B4ODNUa6W7S056dOGKBICv1XIcDgwAyceM2t8ucMjuVQt+BT
v9yIX+klTxWOIBdIoxT6qxEEXYZQcS9R6WQ0VoR8eRCwRtShtYZV3DYB5YmnqFGe
oHFB1eu0mfMqDDLYPUg3beJPgGMYB7cAZ9eo0OHPAOngox/8/nodKufxXfZkb2Ia
4uPOofanZG55TGxU7HQbvNPEOEkhfO+o8f+TB6L6rxIkWKeDGt3v9IBpwR66n1Rg
oSCUOGyZXvvAPctNJ6annmAN8qrE4DMY4Fn0nVprjE5KVeLHV2ABsoo2ciXkGyU/
upwaV3C8Z/6KtcvCAZKQHxJTjQH3CUdY0gm+E6So9i2PCXSdURJHi9DkgK60AyO8
ubGFoBD/9Xjy4Emst7UiWdDVRxLnXzfDbTGwmLUpvMylGKW5w/FMXgNRIVu4OJYw
6CYqAVufa+19HLlzuSf87lRF8BkAatiUKdE8PB6FkA2KGJfoytlYZeYSufOzimqL
v2SL19OgdbXU2vr98me2TrQwpIYJPxeyEYOvBcbCJX0IPehBwmcxktHU8HVJbaiY
YcZ/QEg/PAmrmSU4U6DqYM7xSi0LX2PLOzkg0JABBA46UTQWt5GtyS3mXc474297
cHRlujuAz86bkeh7GFgNER32tUYK+gb/7KMcYd1RQ3+alGv9SR28t/a2JTEsNlU6
GFX+1jtZ1d/Q3BZFcr4AXYw8SSKgBtA33wIyt925go3rIVC29wVYmG8LzT6lU7Nc
CSz3TqAW5xIT25MFeALBhbIqFFVzuwOwOFtQkYRu7zotmUdxDX7oLWBfqXeQoISV
aaT+qfxwYIuS4eGFnJelpWzV9jGnV+h6XF2UeRfx3FEGES3pUugiODV7g90bainG
uhJLYqfuLZQF8bwTmaxevhUMOtYzsZBLXL914D6u4Pn4kNuNaNdAwXymCgin0fWj
ubJcB3YPpZyoedLG9e0g7KqCEm9jQFCqsG5JGWogybTNTaRSYUZWQKMDerP53u8c
m2YlbetQG9DdfPgbrksyr1VQBveoJKDV/8i3NI/UjlRymnMwdLoTtFDQfJ44cdpj
TlKrRzVhPdcpOHA6yz3WAYicEmtEUZjKZbz+6YgCs3Tcj4JaYKBn36K88a0TiLcT
nQB2EDx+LTK+qm1+VcU6RysqDVDrF5pM6ev6bWOxMPBI5tj+Oo0gSyipp1tm9wwF
zIaowo16mgGlGe6mvQ5nzcTgzNkXbau9EFNf/X7YgH8ViP7szUPH9ZbYXSGgOGdM
tak6atdseEiXkMc6qciHmYoA3GO/EF9Dxtfd5nVePVDhpCd69NYK92zsLWjUIgy5
amspfZQw2XtSopAlUeeJKDCeCgUWUL6+LYTSgi5ktVkNDBXD2VtDQqqldy/XQpPk
c2ywQ31YdItPENT5slEq1bYz4xR9qqmytiMHlMsEVrM1a9fSX1jhziloUm/AzDuK
mqTOp/NisX+OqR3Be67PZIKgKGtr72Qm7JlTezilUmYlNJDMiqd22CrbFFZESpTA
duiJiZicWZy8wPfaGXjQ5jn9gjbbZfRkzc/8c+9DQyiyvwBATDPdD6AWe28zKK7K
eQ+56JKECEO7C7CxdDEsN/heqO7jVotdcM7A9hxe8OnAEi3Gn51Ub1PUEJUJCGUX
1ElLolRAu5VJkw3ZAk0n0ff1ccihPHameGJBePIMjqguY9YrY6r8VZYk1rBlmbVS
QR6TUTmttabS0C5baq8KO2ThM+Uk5fN2v8tyjssiRkqdUELjNvo5FAmj+UC+EnuZ
RKRn8gtpwEVSqdNnFdxFlqt9ueWGKEINpOhJZNj8l+tMmmYCPUDLswAFDmERom7w
nqiqI102ff1/6UJ7+ElSIM8encRjWWCvk6zFwy5U9kAtLJY1PaVNPcrvxY1dCzEd
6LDADNyEWJw1hhqdwqfr74o+W4LhFfuTxiMQP6jUm60rnTBLXCNmfc7LeOPbCjMx
ydPJHYcpew+YfdfHRo7opxyLrFHcaxvhl5rNoIrs3lV7sdJ0KHlV2Nv9LZFQlYO4
PogwLQE/h5dPOJoqQtjk9WsdkGoTb0fSNg9HtgTK7vbUkkJLApvtW8NhS8lk1GBE
QXmGjLa6V4MUe+XSoFyTMEYm+gl0pI6Wx2+g0IVrfQJOpkUCdSTjDuK9Cl8SxedU
2B9NqEh8cD9LA7KAR0wsm2+uyPMFBkuMfA/sOpV9/7vOSLZ6JJR51VArXjFIGqpf
00J+VkqnqzYR7ONjh1WBj0Klc3XaoZ6SNjbi0ykMD3W8QWf24KRgYDuzlkJUXMEj
l6Acqeg2zek5O8fSjt2XUNhoLDYQlLFeoEw5qXbdAvSiHyZTSrfLwIk148GgLrnP
WgBLnBMjhn8FWKI4bJQoldLgp+tEgthZgmPJbRCk8lpck0UwU+gNyxpYr8gLFLUy
DoM+R7QFbsA8HSIFrxh4MRHO2H2X9bCHZJOnhPiNofS/72sd98EdbJD0N30I5QG5
9Dy1UHr4JrdnQAdgZqco/cWlLKit+hxdsVCL3hx94QJn7YNi6O9D6HVmUpl0IRdY
glWgjWx/Gx4rt3Y4b4Cz18mQA9JQLjXc57tqGFNn4oBOPuY/IOqtBaCotuDKJdBY
LdxDd84hKZgWvkw6C1p9HthK5XQP3ThbZLXqfP+x6gpWGuugYcRpXypZ9EDUP9Ec
30wQ/wzgyVdTzw2KaRpx/AMryIhQhfmXkTYI7wzo2atD8F521srGd6CciZ+yeEci
gAQqkPVinxHt2s8VTDfIiwcUbRwMZtkmllDw9QxQjjfcoY7np8WE3+CIUY017Dli
EZ9ZagmmJjXh7itC6CDUNOxFBEytTvGTJFC6bssLYs92D2pFipZzSUL2Q2OjSx8S
f3uSS1LwP+/RId13IY34QBiKSc3P9HCES2+0YJKT1srZQOg47ufP588Xa6j/jNKM
7gTg0y2n0gE6vEETnabNcf1iTPQLuPzgS88L7bsWYwlo+PhbUhzrGu263yfuuZZ3
a3Z06JiJGhaOe+fyDp7caWLOs+7ltEa3k9x1S/Wcl/TEiNZ6Lnyt9Qb/TuxZHHrq
ZoLOsGsd7bgN5LMCBwSZPhvC5Ocz1Ll0jQGVD3Oihw/9fdBQejVYhMqskiZT+Ao4
sBt5HrJKumKHdGbjrwYj1xapLWP7gsUS2a9z+WGJclnNE3merYn0zegLV1tYdINO
+hmeb2e7WzK/D+Nxuu8qoURaZLzRRpGUrADhcPAQJUoE1yJEMtDH4IJQbKcq5Eyy
mKVzSLh0VjDXPm2twcHoRpxnbzWjdfvaN1hobT4MHbrDd1+xqmIybkxpLdPbKFOY
L+evtAi7KsZoHFpkK59XbS9OHkXhFyIPZPYp+247w8fnPatJBj58mVSqqAeDc7QC
g1nBP2/eGek7qh0UZsgzOdUGj4CfWlXS58ayjIXmeFOzAXVBBkDEeeE6H7/sBKVP
S4/3FRF9LkY5YjOT3ly9EVchigHQubBaN48yRFXng3hB0P/FEtJwR7p8zFacKaHE
4kysTihihdipr5xU/EGJYQyWp/YH3F96TnX2Pm+g+8BEwoWLJuJzYDlhPXUPS8Wl
df8l4j4vYJNrJQRt2iLexPbDTSDhbPJSEMn7iN0E9yiqKkdqIGGnlMpBmrG8gwZO
MQmdTSdBPVpNk15Gn4HuIBvafKsSdnjDYmsyoKAAuV6wDrnwoq8/zGr7XMnkOJ26
9gDr6jQLqj6h33C7YVbQwzAhYi8Nz2LeDdNwmG19eCZR61uExJa+xGo2emvC3I+A
HMBgz+6M8bCBDF1VimkPB6xW1XbMLzQSudwtJcXDfumZW5HZgwJLD99Ke9N7VIYk
wdDwitcBnISJY6/9z/mgrYd0afVOtsmY4/vOM7AKByJxnUvVhYQj/Qm7N9Ti127K
ceiqvLKklaXh3Fbwk5o/cvpUTNAmpDuQoGW4OqgwuCbYmUUn/axxo9FBxeS/zZsd
KHy7xXvFMJEHxGOTWi7v99EIl7kVXGCVKw3Vgy3bxBcIihUe2aEZWWTjIH9ZUU2d
7u5HwUQk9YqZvmYk2iTXj5yXEJ8es+PGrT6En1Nw9ZKtDejh6nzPRqEJVgRDDoP3
3Xp0mLmzOncsb1v1Rj/RArSG0EZmLnE+QDvAVmoo8cFAlm9U3T6Obx2rlxXku5rf
LDU7683REJEzl39zMldx0G+6r2wQGGYFDUbIJU1ajfwlkVesLK+2aWJ8AUgNLZSH
AognIkopbvJtzycbdosBU8RHN+At86irhDeG4qN56MQf2Ok6njc78HWs/3s3V9cY
Zl1R8gEKLhHETYsxg41KvsK2VIK4Tx0l1W+GKqKzda0svjhJ7YgokGR+FeYarMcQ
qwSoFL9DeVptAy33EUkw5xkYqfziCqDg46gVF/wA52iqooGClzdYmxKqlRymgIA/
fD7eIET872sUPTWtDj2V4YJs6p83S+eW6FTCRRqzhzqUThY5Gx9pmJInaLixpUtl
zXINxk8c+xn/tOax+u2UUL/d5muCmE/NN1/vzkOAol1ArziDBkHl2TXBhs6LDvZz
QGjKYCv1AY96zmvDS5rVHaAzJkDM00MAiRrsM79bDyENbbTVRJFWeGMNMcPX5yxc
7F6gHghlDGVFtPlL0YrHh5LmSsNCldpyRxEDmeXHd3pdGxIOrMAarAgaLFGroTGf
Up4kyJMHq/3yvgqO5+ISKYbzjFKAgHNgNmEnRhSZgpH9EvKUciY+U8Y8vPvo6gxB
nyxQRXeZdXCSAcwNAa8M0BW6vNoYQfIR4XWJ45VsIjhWJrrkVXPzAHryqph7lcKF
rOrQl3e16eVQx3GPgOEHKEuhoBZDYMUGUnCYQIUmJ5PqASdIEM0KwmF0Sge0+YP6
bVzCmvo+xDlg0L/R/WFVP3ZotjgwMmTkAsK00vPmYBp5MfNkF63BEY9IIIwADab8
JN2doNvgoLtJgdgg64eTPWr24eesH4PfyRRc5zBNeE3qZFGvKPf80J7867lElEyd
WdcTO5E7yafLe6Nk19COBO6yi2BEu5nGg2KlWmyavAoyK8yITf+czTwIQQ6r1Qyp
8vRBpi0bF+j+XzfVcCGtOPBJTBcOiJwKgT72+MYJL9b8X3YfrFqjcVI+2SOtmWNE
TIS0pscyDIvdIi49qY1aFvRrc0Vd6sOEXgqgghhKEHwsR7WByydWJak0o0/ZRvqR
KLVyEPCUWJ56FqJ3EfXXrw7K0od+Wfl2FQggawncf4iZGXQKqK80VVHi1mstJXpx
T175h+YacFBb09HfgZFrRsJrZjW77BNBSdztCEli6Nc4emT096qqfyVXwU0KsEFp
Kavw+pRwxex88cp30gjcSIimqhIdLFxqGiuTHxp+FNqrF8s2jeGObgGQ88yb1+hz
Oelpt+zqB4bfjJu7Ux7S6nH45DHqB4D/Fgbf7gOjveghSzP+m2otylHBCMadp/ws
pVONbiOhTDmvcsxBscvU78nObRKx/+026wwchWrOoI9lqDRiItceQBXAwn4ZYx+Q
fXcNMl8WcLA43v+IsQQh3R34Fdj1TIQfDf9Nh1r1wTZG5jUM0aOhg7p+5+5l50in
gK7VHWP26RcRlvu6QU4W4e1CLxmo7quzNxhAg2HlxoPL0gWh6KNO0R8eYsCroeLK
jTOfb6Pk5P//ZZ0+pblZkupzKYI8oBsov5HK+bvepEEkzaFIQN2EfH+vshPe7UJB
nhRwcoziZVuadRlJ2Z9KSeXZt+e/HpW5XV6PKT99eeezZGQst2vWEzJ15YPMFmbS
KFPLeJbghVZQiM932vPfA6vLQmURVJZ2TcPv20L4p521ihoEacu8Pzn6FvYdJOv4
DSPgvq0momLBNF/tW/9wXlZ63EeNxbIT1ioy7ZKlPrNHkqaY0shXYRnGzJwhcoGP
iB0RbL0dTnwi4HJjAj2+3yFdZDhDgKxx6aiApZiE68ls7I+i9+BLvFPm3mKJBwuP
BAYcVLuTyt2v1MeU17rFxZRiEcy1b/FSYjaiVEMmSTtWSUQbfE+YgtT1aam2j6jx
BOvshrzpLDjJFLeFtVhn+clZ7xlabUhD9fGKksEdd0+Sdeuor2SS7kvPbdK33oSL
akhwbTcLHUHHrLBDxZKG2gnwThw7560gODrrHyR7ox6dVhpUJf2j2Srjs50WYe0G
hrTFXMpYwmsmwTEXo2dpkT2NapceNffbU5amwsHax1gz1jB+FlT9xAgZxRrSG1R8
UfvS6bjllglPqwqcMplPrCQQ7yLze/Lf7KQ+gcTr/WjdOTP3WFCJxhYdwa8ykxt9
SQU1tM+dnDc5aRchIr+5oe9/C1JhRUaSDhYiKYEfdaMQJZCezWuFp2HkuWh+Blml
Tsetk2mI8CDhzzriUprCBJid6TR9iF47H4UqrREt24jGXYGuHpnwLDobhV7DTv3G
cuTGe58vHW8DA3RJ/meSpqH8w8btHOZz5M5aXotRdHiu3HF10IhDfqrTTwwyvtDN
yu6WeRpzxSOVsuy8QoWqKQ8KjJ41TNfDbsjL44iV5eM4uHQ7vWm9D6oZfc7GMCtu
wQQxYPMI/RriMKJnIp3VtYF6KS3SnO3EH0e3yvyauP099exKcGn8BZz5HqPhjgTv
VXzbohqBUtjGl8UkWVpZJUdnMQN2FFrzGMtkJXIOOw47HGExD6SfbvcRSppWUubH
wg9pE4XU1X3ujmQO3iQOxlqZRA5PC4eaRrlu0c/8u5fNxwyRMqlr/n2X/gMwv0Tq
r6Oy3eXIJcq5ajJrYUMtOfmjAIgZlFD3DJ+2oZHN4cYhP/LABNf0W6SQnrnUHBmy
9CutRxpGeqgLPgO7QUIUwtEgvJpZu9QBoixRDx4bKbTHHJd6vXIYoXl6LwR2ZMB9
1ZgSxU4tJlGW+fpXLKDpMwTciiIzVAPCHBX/iZ6rXo9qksodOTUizCYazmN3Xbib
hpU8lzaZ06l4iqSKJJb/JlUE8LxNo74kSCyJBkI0YlNKlVw15Sdm96Gwpg0FhXfm
oHTnj+fvwEP0M5svzB+JLOzJpe/05ZDfzVXDkVaqawwz+h4Mcuwnwjkb8fygEdW2
Jx1FxTDj5gftzoIwTdstHw9dTF7/w/4lqSh4YFX+oRlLAnHOB5ma3mf38EFGF2hs
hgOb2vJ5zBao/5Ok/p1UxOAPLTXvIodEGdRc2Hf0AOAWXva9ZlOyFKg+IUbzXFDb
OjePfc9Zm2XfVZQMfCKbhBZrlyoxvDg84l5oIcPc1EEhF6WqH7oD6yvSa7e13LaS
XOZG0fH+XuW+9Nv4Osv4w2IppidOt1n4pPTD4erEdSan0fNno2tOWJufTSZXr/Kk
uSTbMz/oMc7F+KtNrVDWN5N1OtDHhIFHjSmROgqbBXuYMttv2O/MWlO5Dl7NNe+w
wC3sZqh08ZOg0Wh+GO8VB6sWQBH8wDX70/5n46OpqnkP/u0TPbBfx8KzNFrUAycG
Vesc5smGnKN44W+KUNRNDd91O7OmbBfqQ/FMzDZC5ybSqIOOGnTQyV94nJFXlQIr
VafLONWh74fpz6yH9NwhaPaFHxfko7a+Y3x4CS4MW81oYOjGu+aSEUDsdZL4iOZv
1HdTeoKYYOx1r+6g9aTh8VChLp9c8BSgaBjP4X7SjVW+qix5sZhyk8lvZRrkA+kM
ImkElC+L/YhsFMPLpXD4MTn9P7huIK7srkg6x8xFNdHd63qhmrE0va7d4O3YuzvC
KhBeA+6ENngPrRFHtFX2IO9fCUprBXfw0pN1CA5oByrrRBCGChvPO51qMiuzxoa0
XBP2Q8glt2DUEpPB3S22kP023n/hGbWb9wnQRB2/CACGF0kYmSSpOw8rjFTYAYHt
vwgdNd4+ftNjwiRdeb2bMwuRS9WAGF01r/JCxNY8lFLPuc+1ZkA0X5BaOEFm/XCT
prFmz+3ct62t7IhctAiNgnsuPeA3/28sb93qj7kK1zLyxlKGD7+JIQR1lDG0ED1z
n7NGzKRSJG0K1sjqZphqYct/ZqYxjoXrU+FlQekAU+GbfLGFaCBg6ogb4HebPHtC
3LHi3XKnWOSDAnjxn1riFXepjnSOCk01y4C5HsncXQhFLhpLrH3nx9xZnUte2lPm
jxw6RLSyROwWtd+lyTHNNLuRmyQwW88YkGU1SyuPww9nOTV6oB1jpiupMNt7rt8G
oogCALnKIrOr+sI6VgP++CyowUD30e6Wb5dNwdn+eKTlLDKp3TSDWSQ3kqTVk89Q
wEWZRzv0LYilP5CuEIeSC/L1bAE8jr5/cyfT/qP9dcESfnf/kC0IV/8uhqeKkfzB
cF63aV3w4r4G1wJRoS37NvtH1D8uQldvjoQgQlslW9RD4kUbQEWvt8q6tdry6na0
OydOSaJNPB9uChtBfTh9+Ib00d3vtSWBQq1oETCOi7QQUPd0TH72vSePCR238Uzl
Y03AtD3rNw2cPWoYzMuD+YsCSadHG4wM2Dy0/jxDzD8co6m70dfj5RrrF7J1WkDx
LhDTyOxpkf+OrlYvJgQo30bGbdnDByz1WlaDtNHia1PGNfONRc+XPBQm7TDQvU0S
gq1glN8CBkT2SbOzwAa8nGNGxPcu+9D8zb4bhz7hQt/eoCeOr/yRCMzKCzFNKNVO
QrUvBiPSdHx0YaT2waGFcEK/r9sHIjG4Nol6T+80htv/BblfkngChbYIrAbnUned
s2oGDf4Dx07sVt8wTGw42eGaOm1POxTyfI7cj/vt7InPz0TEk53ZqWnUs9Vlmyb2
FzZfiL92DtPKI9zQt/lbAbfmSCFtFhNeFYpCkwBrzmLbzSrxvQ+80qUQJFVEClfg
sZJVlLCiGrTKTCrKJWiH0MZHrtrlTu0kLh5YRvlhgTnieFaTFHlwhLDrnD7HoxLs
5dEAQlT4FC+mUAVArwKz0oZSUrL/bFA2m9IOTFVOy0U5P4Sm8A7F+C8cK1ql4+tj
dZ8iLE40NZkaPWQaWmOCA9nh/08O1arAGIXb8oAP+4+v6MmRE2NvV+ko2GqZuNxK
lSZm4CaHF0rKJdllNFqJ/Y/ajxFwQN1bHXtaKbuCd6v3QuO7XH8h5/Ja6sWOp4hC
CydYh1XA6/8K5TS3h4KeUW24RK+oi91EWeQMwSZ9UruE+8P8I8btyWWgoulVNmrv
JqpweLs4L3zemSUvWb0/y/LycjAgo+6FV4wuT4aEVYSeTfjL1HarhoZBEUsaplmg
6TUVMSOG7X/JmKtK/W0gezKAE02PEqw3G2F0xA17I6Gs9E0n63sj5Fa1s5Sa1lQD
AcJuVax/1hjkxI3A8RXIqiZnn5IJIs1rhrXkC13ERp723zRYmFhsEnqzkofAuceI
9DcTEKCdkV7HZ/q79rx6NzPyN9kn40xlqcaJ3jhAPEUSmFdpaHz7K4PhY06uNahs
48OqLQjrzd6tx+Onq9HbSiVSpVDgZKXlA9hF6Kb1XuUFoGwIKtaBUJXirUf2+Gnn
auQGMSnDrvmcmYrNHl8bSLT+fPxUpjNC6Ak/XAxeCOl4oUCcJ8VljcuzV9fsNyLg
MjM8QsgDVjItOr80l5FhmSGF1HYwZAquQ3Sjqbv0kF71Q1KJXrPEfJPguynXW2R3
4Wj2017MeUQmgwOhUjlK5s7bK1LvLnEsGvMQMoJ2kdHrmd9mpAKzR3J9xlcwJI7F
rL8kIZOWlVfc+LF67GwE160ieS0UkIDRQMTKIr3WBUi/uGtae3qJNKU/E31TsUxt
5eu/2QJ6PRzftCe6PcChCuiAPXVUW6F1b9U+SgkMjnBEhQLebVQGCswzD2lRil3z
w/lORmZ8lxGMtW+GllAsrumASc0XMOrPsl28NUzFfJGhI1z4TD9II8xATQFnJnFu
MeK/SXtn+AumgkqT0CncTrTHBmpwoMLbedDeWJq5bA/+2DotdQKD2+S5wOZYlPGc
s+K2vH72kMqwPBcjKBHnFshUxhVFkTYkTa2/+Za8Yn85TZn6tV+QT3VQDuFOpzjK
ImBhM+g0e1kX+gFAM1hz58v+4NMuYe0LemNXQ+V9nRKYitblQS2PEoUdQ7/25z/9
KWdSl2EAOp8b4R0aAhYsMGFE/JYQaNm8oEi7EG+WQSC6B7/Qbmdg+pMhmYyz5e1r
n2orNoogIH/owYk9uza42icT0piuWHmoSy142GUIga/8erbujcJpZlPn4ywk5JpR
wuslh/T5ZYeRqM/n+MgtSlYJ5I/kwS6okOdV3eKHWYM72FGh9v4klMfpDTibLmVE
bCgemD+clfQZgNW7MYDUgKQN+meBq+XDoRqsLfTegzujjfpJoLDv0m/dyrQCfggB
srZ2os5dFAegkGakgMOTKkf9El4ZLqeIottJGKjAnU7b1Nics+PsvQfgkroJxmbe
bGvY8v7l2Fh9Vbyjxg9sbDJjlSejn0jyDihse8FW+cQLDnxJCz6K+u3hYXd1rbwL
YKQ8PWWOL8yAtq1ULBEPEfbcDHy3WYfcZX1+eJAPglzqt4Rgx23gv2xPVht956/O
tKPQc8O8a9vqURb/si6Qy7pXvLTeJ4o7l97d6gRWAr45+Us3kEd8NNP+NljHwj0Z
pKBUJWRJug6kIbdSse02R4vvBjS3fQf3szspVTt4LCfYhrY9EbXwCi1KmsADEk/t
wa+lXd3sMaHfvOTgfZlbfmOWQv7jUFA6JFEUwGF69dzbF271TkRjFChuqqgGlZf0
9KHI8rg6+A8v8fEKPvNUMD8v5riHxfFxI3lcWcvY7j4xhvNK4rlZExyrlqyPLHB7
2AXYxnE2DH5oeW2LWZ3DURjT8OydHA3xbrkepH84dnCKaxR4i6lNrZTjfLHcAYUS
23erUjaV5jXpNEMYCHJHV3iWH5/QUUY9VgVD9srkVMT8AyOKwYN4+RQebvYPwRGn
e7VZZvuzxZIcxCbE0EKqKGNIQUaexD+w5KyYYJ5Wtnh5GOihFN2hJ8Ptm9hTfDQg
6tmq8M8dn/tWbG1kR4yaZ03OPI1lmOkDH6h2Sf4gWEcOXKQXu0751OjTAP4FWh2J
yyIRwAkqJfvOE1mDHsGXYQw7XM8Y9kf6RiwnedR6I1ZsWbezatmc9Gn6Xjyr5xbE
ys5NicQ2Q1qzEP0lSed8ObN1YomL4x8z0EF9PFyluggne6gcG4Vd8lVnAfzg4t0m
ndsDnAB6h+7W7JZTQZw//n2Wxo8pYB5Vu32/tQWNNS/Jsanl8RcsJObfxH05Tw32
dLbJe7tXb89tTZy98GxEO2bqVMv4zZW1EnSyc8cdqifFoVOlT38gOLGW1RdMV/vg
hglSStv5RS9QjedQLjEHAr6ieFOO5vcEJDdpm4AMyNCExf20LREoE3l6TvzoZ0p2
qh2yHn2xIR5nLNNUS6G4ZUUac1I1YSk2s/y2dKv7ZHwD7KzAjgCGf8Kh5HfM8PP5
UZf6nVUJyTCdAcdV0ipNvp6qAj3ho+8cfn5tsqNBYxopZnnB9A0Qm9ucvyfEd+Ti
POgII41tBLttUoUjX0mmvZvgtzLLEB9sA1dZhYvut1eZ/x84uOlSlNVZQ2+lVZWs
Hb9k6ucTVPt/gbiX1RLN4glPnH9qiFOz6rQwhqRzywuYT1KL0FKfqZhwO8IllWZd
3XZeSQs6YS9UrPECWxfNZFefGAHpozp09zjzsQN3rGvDlMee3fOaJlbRzUnkjz3w
YsZ4KE/27ip2ouBJqwFegeS8j5MHaQbavBsNsuH6TPdoUFMQ0/WrBEA4dI2bmzYg
OQ4x1Op9vSHIWcL+CvF1W6giNSkNi+og/K+H+Re5CnH9Ujd415ZrUxa/8QIhPxsV
/h2/6OgBok3GOaej8PNt7ms3bY1+ymenjeOFEyd3wVezLa5Nz9c9VuBajIffWRG0
/fFbC1DwDaCtfka/qftsKj0tyd+4LGuBqSWEa8NaMwvc+DumglTjOXqJMxVj/mJu
W2M/4aFivWR0/JhXHmwAOsRMs30OnML2Ctb/VZq2RCrSVC94qt/eOdR185zQo7xu
T7eLUC5I4XAjqc5wHrcFs4Qif6cJ2dboIMEYRbDAhJSR1e6wkOmGoK9ksRiNMlKz
f1qyKMVi23vq1MHkEGnSkGvdtc75rUHmdo+VZQ78lhTDQWcPfEDP/7gBHtL3bity
rU49J4vVLLIwEpuTysWNURBWjhYXBzBlPbJoZRvOc19PQbBUiFykgPksStRRSvYr
bSfh/ZSkaYzNLgWSuYbG6jp2qMD2krbrDgArM5aWSIjhuQcoNr5yfxx33Iwk+xWf
IaIC7319eMSEkZBOZPIre+KKCoyyvJtfM262+y4+klz8SGTydiJyeFqz2dk4KRhC
iK3fJsIpETmSbseyQEEdLOk5pcMkBM0GQglhtQOtmmKOFFWBWQJHB8cLIJMtl8QX
n3vt/lgmMXMASGPtFcBxEl92UlVAefTbWQcmEy/HhUF/VeFUM0js2Wa1SgbGbNvJ
rAxOxALNXnr8hGrUfyUM8xJWKoIvTPlbP8Q87iLLN/OdnegbgEZyVQtGUt1qAA3s
NJRM+CElapEU09tmy5DO6/qdrQVG7kJgv/7oWygFazKFY9qZhkpt63pnv020heUk
jgwsrP2bPeUeREi18FLGkmjvUR00S1Deg3Dt2DerMRQxUdISTXT51MURN3MvX7Gi
NuFbwA2H74EjNOKvYAzNCaSWeOtawiiLkHwl/YcIjZ/4meXIrpyRRA1G2rsQuo8g
gi5n6pT0cWzFQWCme+pV8S+91kz00/XuDdQ36DJzuyje+dIAHLi1c5T/loSg4K//
VBY7iKr4zb6Dflxg9LPdzoNW8iQfqOKhvJdrRM418sgS6h0cf3VaSi1cM/PtDTWY
6KRIcgaGOyJLdtYOKA+1ACkb/3xHYhhNoP9jvY+2vkaiRQAAy7saYtvDKRT+ImSD
bT7nIRWJwPaCqfVTiXbLBocxlKO38Z7yBdsVWH4s7il4iomPgzYv2ZcwfN631pq1
qATJaUUNVRj3RP64+iYc9/vNGufQEXDidF3D1jmt18w/37TLyKo1i5GVktXFSQaZ
VeHATDVV9WVE9iJWiOZxSGtTa/JVciYR9qJnBiidqhWopYN5jkILvkvNJBxqBS6r
CYmYk8CFjX4L/BpeMq/AEVeUc8zZO2iAKxIN7bNvJlzXTcO8BZ+5bxohu9XKrGRv
EMzlE+D+EEnGmk+fL9C71KL4a3Lppdwoj06cTMm2+8eLDDTljj160cA83sXlS2fX
9hafm4hQHTrZhyWZWZCkUESMQPbcakU2EGSQyLPhMKIPw+uXn4lxZ1HXD4YOykue
vtvx7t5THXk4DY8NWh2g20T0yBzAn9n9zlX0lMK4gq94OE/uIIltOqQRmjUVG9ZF
2UOJ/JSBy5PG02tCV/FqY9gejjLJOj2KMUhUgm/OTgLLpGRyqonsdZGjxO6+WUmf
xzoD/p6NQ20KU2KY7YhGuROpteCwcXbgbOAkiMBw3adgWFVBaOA6xVoiSg3dXX/7
rrfZontDu+11Rbd7MK0cx0XK07FarG/XEnET4bO4+8+zTcw7f4fQF+slhZSU8Mo/
KcExJtP9KsEGlhBU3nyitPxvKZdEP4g4GDk+fAqn37XjimkuRVxHeJTsRghNLBf8
uRyKuH5dp6RACMn5xZdcn2+UucF5lqveq1r2CIcswDtEfnTMU+3vGma0rrYofIL9
TQBeWpV53ml5eP57bXkeFr6IH79eyDBoKX42oucEUQn1goEYWHioeU8BJII9EyIq
GBlS1VGjxDyMuouxO/3j9DY+u6S5itbmMXGq9ct+6nRUBOBjPpPbbPyrc14Zyu6C
GTcrZwGsnSbDWqvX/6tpMRq4OLpohXRVot0nYYeLMr45lPMitRRIT/cy2UKrmKKd
5pIBFdGv+ZgCLSjWHwyOkUEy5prlZBPVzB0oEPCpeKLiYhUrnYnNqQBK8fHkxxcy
Rl6/4gsfqDqub0PvGU2BRfoGEH57AOI+zi66FXTIF/vjdKUp9XxF0BAJwwq5Hr5A
oYZVY8QSasxvxJ6zHzEsGeEwOpuNEprcXGe7bKh3n5OF1TXXkqyTIj4TrETjQc9B
1t1lBcxoZG9FnI1GUdnoTtJAQ3hz3+fLLq0l8P2ywVCQR+VMoBx2FM8UKepLyFhs
n2bK+rDCQYotKnpe0aFYVP83r1REfJozF8nPsZX/ZSx9AETMQuBlpbSiOVTjdElY
a4J6F1nP4ubTIgIW9xzhBJc4zxfYHLGcwCt3GKgRCE86gH6Wos8YSIpU1WUWmBoX
iiB9tqOBFU472jY98XZf+JjAXxTUqczEyRSwVcKVI3u4EglRb1TW1JarFt1onMVd
9JiCFHAFtZsYGjyw73eulXBMxCny1G9+IFXe4ZVRg+oBPveFPurB7gethBM7XvpB
ByDmxCnWY/dVJiV9Q2a/CLPeiAZ0EWWWW7i5t9dpQZX1XWROKEdTFvxFGdiX2gTv
zFV/uaNG5CwL3y6nzMb5KVkF3ndIrm6nuuexj+VDOxffqszFEFbCtdY0p5c4DRhI
7lWpFUgwRw+EHV96rjmMr7EuUpEDH7C+1qqTU/PJD8nBa9ZhonEUPzv9miiCT0L2
MCdLRzyFiMfUCjLtD9wDN5wSym4yvMS+ztFgavnz0661SJxSSOxzPMguylNZmS3T
PiRS0xqq3cK23UOSS2wG0E9c2lBe93540w2zG4FjZ94N1v4QHCQEMC3mKiw508Xk
e0FlrV0IplXz8Mh/v58LjjR3KG/xYK9Mrgs27uAJe35lTUgoDk2Vr4CVCbnG7OBN
tVJ+jqslRd+vx0E7ztnZOm+XCQCsEN0ok2rx4DrGd9eLHZxY0mRTrObKH50NyBcv
zI3UtUhR/A/PHLYW+h56OGGDdspqJOdH2+Oq6bZk6jZnjmLJfX3FAqlJsS5j68tk
vA+dWP3pH41DXSf7ztI8/DZYl0uZ0yJWiZJMJP8K0ToZ9UieqGAiUCyPvfp49F8W
aFuhkBIZG+f83NEgBH2OgZMVDZIHtN5UH7LegOhdZ+hbaf173J+R1EN2krFLN+Uz
5JKAbB3gZxZRCKJ7hJVU7t0f9YIlDUqTK8lLUA9ana4ThgGk5+s32m3GcWQnLiVl
dKtUbVfYj2B3990uw6ge6VGmGUdx8SbwjmRsCYVOWVFe3BA+sELguSmpKOmWzrnU
WIT58cpaVMCnMbbN8JpDPzyeNxatEJ5DZVZu1Z16OUvuLq0eo95DRIcrw3IzmtFo
yCMqiQrHl6P5Rn2JmJotFuTxOHwzN0fC8xfaCYZj0rx8zUxXPba7dOV5ymTC65N+
YaAGoFaPX+bdEwir5LT789hQqpbaKzS/WXnzWyCYlamL/G8TMKhidXlhmZdhwo11
cwIOW33HnNUiuRVKQRlo87vDQZ6YtFLaaKW8Zt3o56QgWISs/5dtPj324It0nak6
OqLqbMXVKbzJEzCnQDWPbKWQxbMiP0phWktwvqZ+4ZhsxTb1rO/BYySp9cOk6XoT
b0TSAgefHfy7oGjnOcto/wFd3/AiSuHaMu6QHM0rFOpkwccsqiio5SuYf6pRiE8j
S2tMQHjf56HZbnYca8YZQeL+UCI+VONpF6Bg9WcF9Yj/pTcdFkFPaB5XFpEygm58
c6ZH03MV/2r9zj6FKybDvfSHMeXLi1h80Ua0D2FGMCYmL3pvkX8CvZ/OZ/sgBeoY
plP2FxMx1nTs+mcHt9Eir/uVGZQppTP47lJ/56vAu7jTi+Yk6itWsi/OFPPlpwYd
yyNxZJKVfHehNfT0zjN7QFTt2W9LPimPR45PezEEzJAJQgkOWF6mpFFtMt6vC36q
lhZ2NTMZamxwFWu+qj5AUqjP2Cb1y3O2RXNhO1Ct2TpUI5QXz9lzOj85Ss8wZXo8
70gr207CtpPMCdnKvDhLzuRNXUs6TP5tzk9ZopbV1wPsB6lgBEAvp/OzFyu65k4x
ZEfX7yl8VpvUVGlI+8V09X0w/iQcfoevXcQdhNi5xkX/84Z1N75P+4+PSyn2paDK
wWezRkBkzwz0ETxQUgjEChToLnkjMcXudievslKjLc7akj/rHZzQPcvlNtp4HddL
6ZV776FCNTq68W4bNFBj6ApV645/coskhxl5qDpS8zsv+uzE8CGZQDX7dUPYZimy
l37e0YLkJhPyXamdb/sXhtk+RssFK6ZTRp/17aJU/jfZQDY+AvFyzIzkPXLhViu7
IGY/wvXvs4ntFQsBPB203HfFAgV2nmmayyGgMer6C5Ug3O03vUpSrScHkHRgIDp0
02NyRHb3dsFp32Tb1fWpKfeNNByne5FREp2gKymgF55MHJxXufo+YNhJWn1T2zVq
9j+7Dh9QUIj9swi3p7i9SOZbE9sVCws0qId0qgcAkrU5RqxZYIkv1p2HibzLpY13
q/6dl4vF/DiNmD4zH39KkwgEJ3TeEid/V4ZBnqq7i8et6mPFb6THz3q/7BMBDjMB
4b2yx/FewHV1b/Xnhs0eWGT4SLj84OaY/n086f0kQkiiBshUI+LxhoNvxftjYsfh
Wf7N4M68Em3HrF1+g/Uatcf7oeMqMW1fmSzc4y+EaSsfL1reLpHp018MltuCEAtv
h1qnQqTQLuyf3+HQFTseNO49T3UkXQGfpszItlqo0waqM0vnubuCwKknetLfGC6t
rCS0583qSO0jFMFosFUiBYTDRu0SETYBjtL1nHva2+ZPDMycJbfFpBV48Q1VjbPq
TUP7ehyK8W5a9PtXx0YNZ8TAjIATu06HkfVmSMWjqxTJPGk7PkdKwb2ezGeqa7GW
vp4VxCckFXM37eISGhY2kQWvTr3MsszfWoGgHz8k2Kby21ECTkfHOoxzQf10aB5z
nQ7Y7xew9wCr1gW3JBI1ArEErNhkDrxTWoYjCFlt19aBNg/2pi+YiA4hMog6cs2f
lhPsLnvoYzKIbNixoIQmmAO/CMhIib1DabwFaACQQXf0zs3OyGfL/W1ELxZZaQDf
PL7p0ZpAkf7XpIalkfF4fa3OMzkgQqdeIOEZXcv5t3oUSPmBiYGRHGzlLFFJZvtd
akABedJrmnEk5F5QARpJXai3MhFvOqNBhe+4dbjiVD4GLbr8zJwOxkYhz5dNKKWq
t6ifROTQanN/r1ceoyi3HmQgsUCQKvZr2I+rumYbvTegbaBT0aADUSncAQTyhOXF
yZxTvlrNxKgiY8Kc/N0xfVCcfVAigvz2VIeVPa5WwsFTteVjJYzhy2fSzcxllg4p
+3JVgGBJQxRNujGosoPSvM8iSvikIq4MSfVGFENvU2Uy79TN6AZmXDTVLnEjsIX3
egabjMdXNzHmUkbVs3rXiIunVwjNTafRwVBijQj1YpXPF//dpBUpyfkdhRXTHIA1
Gq7iVY9tMcYrEEtFCX7Yp32hnKmLhU+ge/1D4fhdQDBxYSl+d/TbyViKdRWBNd+F
EYlzJFkQIFCeHI4YBCZqmB+RaN8gKy6+bT3WWaKaiXTJKQRePaYht4a0xxDGx7IZ
PP2jm+3ZflLbNg0GxEQiAkWJhZ02/4k/yDPFeX6QJGYJJz8jNQq8AXoNZojB8k5o
boR4bVwEwSot5kw16wjGDyrqIyu3uYFxps/B0oJ6dUGWvqlq7z9FupYac8clcgTu
HaO09HIDLMd89UVVxKTrgfLa+/Vx0bhg+gItRO4DFItF5Iuk5nchFnXMpJgGbXOT
MMMtN6elsS4gNiNHSmaz3FEgyn2SpCkI+qCI1tIUR7UNBQbdd11xpXzFcWjtEpnV
EYcNEJsBOrhqP0MvZanZCMoAfRnJccNcTQgktcBpjeirY0sI+cMg7BidA7oh9ee3
0pu1z9ObXmhJs2kse8b/pBHGtpvPcoWKixRUTcMJKxJ/l2g6qKI3CMzVSPQMqiSY
pD13CF9VA+SeAcqqxFuqgxfCOAK2sMgNHdUjXHwScb7tJT+34h3/aqI4uAAttlvH
vndYoABV3p+NNNlSO9LfFqDA8y5gqyLC6hpo+0d+x02PaL3JFhpis7Uw4eH7CNY8
EkqYpnn2KWhfLQHJBYaRv52lqYg96MXpSnJ2JOXDPNZiFTAYerBIfQX/5k7IEVU0
HUfDimJXdcKHHpikvlfVlumlDU3YkLahkySV60ODXHgIhZOXAqKvLa4bTHRBt0ie
EMartIzYBW6x/JndESCNAG+ltykDjEotL8Pt2xgP96zvOPAzzt7k//7LT3CUp8T5
zzONahqfzxM3ZuJrGsYPDooNPzKpHj/nJ2Qax0oY98WD2mSQrWIyzT4R/CxGoRdW
V/NMpGEPw1yO06NuZXhagASaTE7myCUGVg1Qdc07Mg7Y8YRq16OopucNtvf0wWnm
dpHDxUrsUJFN1BZi3uyuka0Rpsdjr9jZ8oGMVzF/uUp/zlpNeCm+JAK382bNAZvV
3n/kdBDFSPYr/xNGeue0Hq6BtivSZX2wqCMPgz+yEW/+m6tgEevORAjbCG66e/ds
NSFzAk7OHkr+u3dkKmnlFKbQOoZ5IbppDqtXXvMzdD6Crr22dhJRF867IdL75uD3
zIDHFF1VkH/rvcRXMuGKql5xK9GPR6I2OxJsh6CDqM1xnw+KASqwqhFzZ1fBvhb5
ROTRS97oT7PvFrmQV/Xk1zFJid5vbs6Y04CxA7l5HRPAYEcNSI07ST6WsM1fUg81
SRfxiT1z06Ux+cPEXnH7Rwu8W4firAy0280GoyzwdywsXgAvMjqBjOYhxrrTv4Gz
9dczR+iYJugP5uQkgROKI38GZrVg4xdIfTXU9SO8VDGImnvVyHpLPtcGyBQDC4ag
KL5scxOsDtA4IXUFdNq+AoY63jUsTwhzeWFKKbUhWUQ3jnuk3YOvc/vjwT0b2ECK
+dUEPiT03A0PhOjvjmbm/6FjmoTglQiNjZbKjfmHwfQF+BQVZHRaEXcOdRQw5QPa
zss3TOn2zcHnnjFnbi4kdwEPgLFBJfHxQM/UBBUf1s1vrR8jHESx4oVx29EJb0o0
f+nnbsBH0SGOQSWjnMYrCYCHQk0maqMnz5SKYN8BJZk3u41N4rDMCXRbgaBxdRTj
kRZdzZlAqpfgdgFin3fhABR6kYXizfhu156oP5z5GzZQLQknqE9qJAzLp5ExKlyK
nmCLwDmjwaW/qKLGz6nAn4En+PI4GLPe8J9tVhpLavZrbRk+u2wjY0HeJ9xIA2RA
80oMKCM66zB5BF5FwV3C9ETNAskgpfgaZ4aC5qFNjisnw56OSMrHL+YT6/OsO5ZP
uk3BWTeFpnO+Wd7bqLaOee3eiYzw6bs5rshdiGGYr/T0DzjNZrbPHlvD79tHRHHj
GQvs5+9+1QJq+Utp3HGXf+q2tAjMVCt7EYLF/vU1h85s+OXA2OIjzo0cd1XRf4H+
a7uYSW/RVWBvmm8qPux339zWu74Fd3aQg4AWH7AAXZi54VYlp8VnZgwNnROm0YdI
knNlSMnYEr2ZaXzbr9jkibMG1jUihB9+6/KLugJCZOUI0HWs+qJ4zoUNeGenFnR0
iwsr/txioPASTBWmvAe0vs8X62902bSLc/2iLXj3JexLyl5Gh/DT9ZezEFRqZ8d1
5mFZMETnscXW2RkIGnlBDdp3uyMHCIIoHTlQ74TYZo6Rb9VjVT79PHC3itJEXTs1
3lmwRRgjE106Vw6koSzle1yZHgmaIuagRJ2luU92a6E7wgrml8ehBd+DrTIS8n+d
LQaMLnD933I65Iq1c9F/rRuvX1Kdj2PXEe58Ua7axbFI8EpsteSgrCGhbL3CCtJ+
kyb2a1jk+2n4P+315KJyFgslf/MaOzGf2n4oENZoa5W0PrN+/5k0Ih+d7z14yYz+
iBJm0nqcEA13FqbNe8CamClT4MQj8xZYZ+3Jfr69dwAqpxhHTAsBJzzaEbn5EpF0
ON2WZIfdxKihOY/74ShhfMohfe4Cu/nTDfm/B3Jr+PreXmEBXwJgNqYR8t1weGkY
1zyhedJba7lhknYNrgtkGlHp7DjjpkpH+3dNFEP7yng+R/Awd8OjLzOfOt9eYmCT
PHmedR+C7xKG7euZFwQ+PeFJe+JCkgv+fJ3tQWPtcJcIvodsg72Detuox2N8zmCN
xrQVJnA8pQFarn2iXp+d6Wgz4l9NDH5LiQY4+EwgzY3MJ1Hbju06b0J+u5vo1y8A
Ld9UFRydGkGzI/6BCyIMfq/FQIAyv0CtzSwTvN70qthmwCvvLYVlU1WEc3v31T7H
mn7ppdUly+TF9Lb2X39ttjAbAeC7/cxha3K4U/i/eDs1vFZ908NsXK2tqBs4tuVk
lb6DFN7b8KDNByaqG12OOYPFwOBLhWTJp1vJjmU4yvcwbQSssLYx65XkhplPcpj6
oS75E2mrUcs7nBI2AKdedAhBnUZEw4V/6guy6rJQDPA+cKxfAqo7iUe86ItgrN7C
180uH2+W+VcGT1KH7QLx0+glmYL2vt1ZL7lYgfuF6zFMdr9/v1hAIzFgzY+ivdk8
Q8dkf9Zu8m7ieF6IDMTfAhW1oECCgiRruX/KaNVBp0+qnOrKnEIXbDh1NfeF9FrP
TvGKk4ouwXCU3MHFrO8iQPWIFIA2woldfXncdMGAfFHx4O5DpuiZvVoYFZqhhh+N
/QQclmdm5lnuDa8+cl3CM9VVyw+HwOAiMBdbpDW1Eo87Ftt8DkxxTtj9UkG64xS3
ysPqxuNu2dzviPEaHlIYlYTFJLFvijaSHzIfeYdOiqGPZqYdn0Byhlugo6BSIFR2
Ndkoc2yybtAkB59+LSa/wZwEzU1voZcJPytbK4uFVDzZK4iXi5jk5jTZXmiE3wB1
f55/8ijfQ0l6B6Nl9p27QpuFMXsm2mp10V3eNVh4AvRo+Aio+GfvLJbiGIEdvA05
9iScmhRE3+al+nvmYUB1dr0VVm9ADsvuSEf8u2HoIuYk8R3I1e9zk3qUB1IJGueb
c25Nuc0zZ14gJc4dqoEBFlDkaIopascbkY6b/caryWifBbmGnnZMDEABmoOVAthI
UNLgJskHqSKLDEI/b98WqTIN2M1+8NvxNKXSecXXBvFtl4zl599imExFCrzCoswM
lrPFz0UyPtv5A+gMFO2LLEJqMru0mJfwxvVOz/kmQZOSve1XHfZnjUlDkBaZDVPP
SL1lukRK5hzPGTGmPyDTI48K+e9el/SdUxYBE4CQWKm1PbIDlkVbcVX3gKR5eiPy
zBPrhQmXhFJomlaP1mxSBehGQ2N4eH5is2OBnehKq9O1W+FQyycVfZDNO9McSpqJ
XgIfIH5hiFV4+paAxUB64XnAGfais3rPESdcuXQvtGM0XndDEFc1WCKDJyXXLJrP
lHgeD1tZSceLNuh+jVse4KDsQmesB/T7JWk8fXAczQaghX3gHfJxzbDyE6mebuqe
fvW4BgiYvfqbcZIJ4y9oq5MwhYY7qBurBLEat4rKhZyyzn3QmtXBJRC+SphkRAn2
A//noZWqGPtX5++vFq2vx3pArGZlqA17FkBhNjrPg78JQ0z8vUaHtuXjftnUyhO1
mZ5oxUSyoPpb31RXWAHNMId1oGRh7Rmilbij1t5Nh7DZhhF25ty3e+Bzyr1B6XAA
0W/4dtOUpzBwq9DqlTMpE/Nl1nFKC4xJEqbOc5fyxdzJkXEGHpd80XyBtaxiQcWS
j881lFC35JvCKh2O8uKn2Xqi7w4rsx+vky8kUUxAjvzLRc/Kd+UpUnNQZg5tGX8J
YzXRVx222gUW2E/wOkUFw8zznkqQlAmPi7ZJIsKz3E9kjd+LujhgmYxewJdVdO/9
31XCqdSAFPqkSlbZXUDfawcvCCpYODDHmdgs2C1WK89P7b3UARuoV6yGO62ZGnKb
QGaNwEhEGiljteEtla2/SErjx4EX3TAUMQ6yLDPLyaCmZtJZNZ+SnBQMNmEh8FLW
ChStlP2xdpi6NRuF2l3VfwoP602W3Wwq7hBJlB4FAAO5omC6uY+TegBxw2dSANd0
QbvLwGirJRZNJnndFwOpiJLx5Nez+TxOpqs70/F3M6Z+r61g44WJdtAGQM5ilP3o
YptqU9leCw+vHAQCZC51x0y5PuAPpbTLJ4HBkixiwypO+OjvOzCrh9nw1mpdJ/aZ
8wuD/d/RjNXpZGm1Rdp60SMArMkU67pLK4fuTCIykRLiio/fXS6xFqhgDtbUGGkb
6zZ4cbDtcrwn6yA/zJVi3NrgVFcfJDOwSG3l9KDoa70z70gqNvh1ChvyDjtw3H5a
iJAn0tPth7QKpr+YsKStIDSZSqdKDJogovN2DidcUHQQO0peqth3T6faoknKvaO2
7EVMxHwnchvaAH6N2zhWonp1ThosHKNJRRw3jsAyc6ODOy70+ZRteGst18eRF7WD
u8eFpziKcGBPyBjXNAp2KzaoRYdbxfhORAWqF5fkZpsBaQJl4/21jWFzCCvDEGjZ
ORhZpSWutQVf7I57g9m3odXmy2O5iuGKy6FJBBV1zq7oqLfJI8skT/qbvQ7nL4X6
W3y7i5ZGqsoYc0ZkxXLtkzWwwzvSRkZdWJ9kX9HbVo2uQS/pK5lmpKb/Udbuyb1X
Qff4UqzV7oRA5U1jpBGsdaKKSFuCteCkyfmQvScHVW5MS3k7qoRIVypdO9/jIz3r
Z1eOczbzSa+UbshV56v8qeihLWX242b4p+GqjHmiDX+6BHeQ3HuwtFcbhc1QQlV7
+TcsBwLgAxN1tPzCrHYCtbhwp6tW3G5PdLsNkEknLYFAswqqnxOyTNR5G9O1a4Ct
Z1Tgmnnf/7bH5lQ+jcZTgDd1D9GOYO0WNWBJA6uTk3V9LiNNc9zQ2o6lflfIcVzk
nyTcuGyAK5e02Yo9v53NKvu8/GnH5sMdqT9S32EGhjmOnw+N455Nqj1jVsCy9ImK
Sb31xXrww1RNnPFY95PGquN7u1xm4/Vn//CtKl8rOTpcGR3/roCrS5E3trdOSH/N
VAJp7AC0mUew4RO/cFP2mN6m4H+tUjWzxp7tPKufRLYSW9p+yLGNlVxcHrWCJD7b
XuzkrLE6h+3knRgpPAv1hqXisqGQhYZ/HNr+aIvOBjn16ARbqDyeum9Bi0wWUum+
UguOJKmOX0OlBD9e0Ul33RPQU9tmkcZL8Vbms4SQolw6diE1UZ98FFGmXN2wtPWd
DROmADXLV7h4wlb4azksWy0UPQ1OEa7oesGxS7f1pMW6SodWraIepXoqols5Fntn
6nY7Z7uZtS55yev6qdmTr/SSNjo/FnGecRJXoS9A+d8RwteG9uS4IBSdJo2+mwwO
uVJkk3nIVFDYiobAblCfb/N72AmACnfn7CfDyS81r2rnd3Cpdcij8JGlsCeUBkQJ
g9kG4Ts7LApIhKh+DX/m4IdnPCtB6I3LDqRo2EA0seYGRfAKTpzK9UJtE4rEf4II
/zyhd8qflMZxL43kje85EaLSXd3TArZB0tTb0HgYpFsQAsty+g5U3/Jlg/7MMi7r
BuWsTCg2HhwLXryj9rukF7RKyrWwhoWEmHUskjXHuGikz6gi9OLMM5wQzxLWFOqY
tl+gDJDsQX34gyhlxZ5jnAKyz8RXuyunkyuQcF7AEMRPlKuewz+HegHRnCbpQYYe
LeS7IB7zMDIw0T2bcc1quKd8Ae9s5YY9/a0X8p0FQhZvDY2jWKcD565jvCc1b73D
2jph2FkCT9LV7FyiVSNFfCHJBUPC6yh1Ngoy0xMV/xxGgfd8Wp4f16FWYSfEz/k7
XRRMyINXxdvI5qnuYbbCjAAq6iSdZ1CRMyvV7nxihkSTyYlNhSK3e0/IUDRTa/ND
fJd6F7ZlHKR5VBhVSAqK0dlLMQsySadQMOmQK/jL0MySZzhQJ09LLlY3OA94b23i
KxXDSCA3Y+YgbmaVJhoL5w/H35kSFYREUOfhOZKlSSuDJSRTYib3BWmRKJuWvtq2
Usjz+vKz8IruS+5Q4VKnRa+8K0E+kCXQuTdYhAoWsuhoDrZvPjyp30KsrX4cMm1P
CfouHp2tnwiQLqxfXpsXDj6cmKQUcG+y+EUg3djmwImC0uy3/ohAsFEC5CL693zs
ezjAYbl/WwvFF52L6ewI3FRJh01WsnGG7Sqj2ORYUr1MSPw+h+YKCmVOaC/GdVg+
iqwDsP9Aj/kXHVyRgdcYmAst6uKorLMdwup3UDCCHIOUb+/rq4jsBU3/umEqmH17
s8JEN38P3xUtQr0wcQfqtbc2nF8gOiCLekzX9an9vw4WzvOpCP6WxPANunMbCnaB
wUy6yKQvKoFq4nIgQNUfuACCByWSa/AMCiyYJP/V/kEwkIrLxBDwYMfWv+wWlA18
cwYSarLTI+bQ8t3+R7oVCpV/AVnLcDpXjpv9E4kZP0Yu2MfDSz0c7wgRZm3B6LpK
Jvm2qLwVDiB/c2lgtMJJ/UTrvuAXI5ZHD+JVCB42xVRnWYV/kH8YwFHfKs/P7FFQ
eHuknXGgwTgeGJAzrf85lg2ZBzFRwYyfkbLnFUR4VpwnABI43+QsKQGLgOgZBckz
mTpJOhVH1RBe+paSzR0MM+hzNLN7j5+dpsUXio5gjsgihfSe4NaJkAce/qojYNRh
E1DOA5c3YlwQN74lFYxXDxk+pmhDbw4FE9eClDJnNxsd2LqadK+FTkJS8Rq/TlPd
aoD5IxVOo8yGz3c8CFYP6wlZxkJJOROK18aLVfoqAYU1CNERLpjPbu81Qs7sEkA0
YY36LJ/LAaWJzovF9Rz9Jo0QD5R+HlIMfEZEtfX6jhCIt9qPWvcaY9EuDejrumPB
KjDLum3C1187Eq6pYITDXxGlzmdaL01fggsFJgcVB7VbFhQ7gRIfFGIaiBiLVQVx
7Q5ttgfmG8l57sY558/KocMUeQmYP8dSEmmMp+Fik2fXjJntmPNKa1z7vSx/dICI
IC+BrYpPMCGg57aWZRSB/AWo53xNz9fSt1GEq+neg/U2jUxawNmrHprsC7BMrR/G
vKn9OxaPqpdJocPkSXl06dyUpWo3WvfPt0RV/AOsTiGD3UEIItxXem1/h6ngDtIf
t4/dBaWhxP/ZVac2WqKcyPouEJ3+nsvGS40DEWYzcITmvjqcaP53SV3fDdSWDcak
Sspak7g9oG4CDR/BnbivjqIoGrZS4dbM7W9EhBQ1b4h6ooSr+joS5j14ku5fRrZ2
2ux1TWRstwojDUacEVwvvrHLDHHQY2yhxh6/as1/cTlnAZIEEyEVfIEokC5fnh86
zrxcg/DoerCKCfC/vL26B00MZeQ702rMRfKMHnIxfSnwUEQ/Lb4L/HVgjLDa49GA
oL4VeNiNto0cN4o+QZljDLfLx1kJ7jLL6m2UXHJ9det8EDjFQlNKzo+4agKzeK87
6NKlQ6/PVbQ7tj38PD5g6JwLgxwP6T7/uG+a7yacNyHuYsUThj4U+mMBAkXaolwj
ZJVAU+n4vuHAvoYY75fw25lKDIycD1JM13X8gfbH1QO5woJOCxr63rpHSkAufuUX
R4OAZ+1MCCmvmEvJ2tlMCt8xVlEJz6ETPt13f2CgY8GUG6t2kSKs9Zl4EyMqAk/F
yKqJkin3wxZQbfMSeqf0fubwZWOVxJ31wuQqJO9OXAjjuj+35CxQcXGBChHnbg6E
drfi4T7EVkKsGJ2vlY2sW5OfUy36JCmOhzffbOWNkSUa1yQzn1D2qxVQk91rypdJ
FRjnvAlang7AEISlzzNXxVCoSLmKObK0KxJwlfaHFFnu/EPyTcNd364rZ3sTQbeC
rkx3NSJKZgqeM3dn5mw139xl9eBzumOPk/rLOQCgGi/cJCc7CW5+/7hzQXfwLiyf
L0yPTMh5pZPOAhEKBdFVla1FhVawpE/zk3zSXml5QCCcrlpIJlMCCLrkekGI5IPa
O7QvLmJvdkZgxMcUGwbCHFO4sNhlPWGHNrKAZPAqyHJBUG7DivMxPJ7LQAUZI6+t
+eG/88I9UCYf8auP96+TD2zsH2tyu9rF7zKLriwPNS65jIf1W/nAEN4c1iQPWggQ
icSSYgouOOSs/nG96pwmTcPYWb/RakchiMdKEtAX9Vl0820B4OjPsKKklFqNCvSu
icXtvnIj7XVvvOT9G2yBurerV1NCrkVVRpy9WEQbtR4eJFGERPzWTCS97k+YWFPt
oG9up/r+H5LkN/kSjG/gjpNZ4y6VdAPfEwHrUMiyIrq7IdcFFzILOnAkbwEmkfZU
iEpP0QACmCA4p2HvlfxQRSgUuyozi7LAjIX48ccDhS7IOetUJv/gOPaSeBAQ9o6L
AKYcN/SwZzJivJ0kGJSYMM8mnMV74IWxA17oq/ESTYp2SZvDxJJiDAzIx02Mn5MH
oNq2PJKGQhpCBILF+NZbCBa3jlRD1c2II/ahgwiLu9/UO/2ZGNTyxxZPd93Bi+Nl
59o4FucZYqpRwyQLYWkgWf5OYfYW+UwzmVTwgOWM5ekY4UIgQlq91pgDZ+N3ujqo
PS/UIkMZq4DwQKDyqaNp67olfaQzwdd4AC6i5jOjMnu6dPKtv5W6XciXo0/ScM8Z
v3ZUDkpFwPzeOsfDXTxfGzAEHFW5/clPJ9UDOImVi3cgM8KlNAqNrb9RibxypFus
/RTWc9yiC5jH1E4bWzJc6Ez9V2H0q+muO4uwAuMDFrY0gl39AHBEgsrRkD4chaGi
JyiDry6/Bh80Fjy7nnQVrnX07KxzhdrnKgvRKa4PHn+uYySq5/exOl/h5WATGFul
aZM5hgYag9qB3okIWmy15Kk42ZeriDLBv4i9kJRrGLzYh59Nd5c9ezSDc0k+1nsA
weZa4hIkgiy0mpFoaJVXBfNKlEc0aYOKbk5OpIejrhhP6uIUBWa2I3RiWWQ8yBQv
RNdDV1BzAGc43pvz7/qoUHkSOQ+9vDBcntwfDCGGLyG7VBDl3FnnxpXCwT7IrDAK
FkNeTvC5wIQfsr15bI94ThW5LFFTfRXtSRws3olMRoqbVfAzeEtCd9m94mYyi7t4
FnqKKyP1H8RoxywCSTlfKBwuhbzRycp2JNIdBlulL3BeDef2nw2cm3UdKl4VgrFZ
r8reEFwJ9NjVP0sQ6aPipM3nqyvrIeJ1NCUxDqZtlVQILVTMxSUiodG2N+ETleBp
gRRiIe9L2SkdE1o2ZQBXszA3xF+MV6FE7i/EXPznvBuK3RfgTwtkqUZmwfaju8g3
Y3iYG6CPtbVfceOkKGcu9MElCyCOe1Jw7fjhS5sXJdvXzEzGBOnHNZj+42qp9HBw
wzyANIwNzSVCbCGFvjG6Ht4uajadzeuWNCVP+s0SYPGnZxP4AGIG6YAR/mU1NzRr
wOwG+KDZxSBz/P7LAN5x5oH0B+5Tx3q6vF0uQL8/KfOz8OiFpxSanKzDWEFp+Joa
aCwG5qbj1dXFojyy2Kfj8fxTMw8thk56kwKiZyqcFEighc0G80Fh9bogArm4iRuY
i0qMfrZdvCHzF7PaYKWko6Ug3y9jGpEv+UfKy+F4GbuYGxRb1uDIwc9DkpJ9dhiM
o1Ci3VpXUncxkcIB85jVBNSFdDmN+ocrsyAmb67Tpex/WtrrTrOwIdOcNaipUNBL
xGY+zJMshlFfy1ji+uBsRqqpVYX4e2zf0o1FEiSL6OSPCNC4/ScCER6EBNMoTD9d
IoDVKMTIoLOAHO1WH13eE15Qfj0ujdNx203X8/ikQ7P07w5zBSgubdJqmJAQZ2mC
LhsBjSoCX04sIwB3lTYMW6FzeKynG5R1rEuctvCa5oU++LaEtdn/JO26l9rB92tF
xnu+mzukok9WqkxouWDUvgS0wJVIHGMMDliluTf11yhRwBcCdRUuPxUPSp4Sx5nW
FzJbiXu1g3Y/HTiSNWJr05YsOg6QAVD34cw22+uYbYyH/XosOCANJndnxigfm7e9
tIZKZULzvvR/gKsPgL/FPjadV/4ySGbJzmUQ9OkmBvZw3S8vWbOmoAK+Hinxd3R2
FOSztPbJBnLRMXk9m6J4i9YIYyG/DnSwH5XsMMibj1TkFsjPE4ThT0yFhzRlzx9W
qsXKx+MJM7gXsdDsdQ9l1M87Jw0EnUyNUPaW2Nn1L3Ti87m4murxSbXL93xtjEVR
M1YhAJI7GBvC+mqkgEaOdh0mhBWhNrAZQny9SyAxwnxMURAvl1rUygV6W165q8zF
QuzLoFnniQuRKBP8eLUchlX5hGob4Z9FwdKejMP4SxpzFQPneVjqNDLujnR8yafm
vq6YYv88zlhC/86lpDXwWlT3wjyz9RekF8vM1VkmHkzQ9FBwTOuP4Je+fj08RfER
PVP8fnzjsDAK6WaxhqdNb69a0c8Xt5VcMmbzLOKrqOhTnf6cLWENTilRt7L0FLvY
VoFggG3poqXYzU0wMqqkN9GzO0NyEzcyoPUB1pl7Hk6BL8kP6GGgDv6qGqOylCe6
o8LoMlyHX8hvpRTpYDyf4t74toY2w7r+O8199WEIFoUO+gUoL3GOSgnbUvFhoFmA
TYXX12HFYAKb66h/kxpV5OVJK5qhg006OMvTSXKadI9coReP+8YbFCPeD9S+bu7V
Gtbwuou6q1IdGlMEPl9dTcy+yZ3NZljfr55a2WdDz6z+bCm0Gfev6Psh2iSej/Bu
W2URKxmtbqwidPFf2UUJcxSea8QkDQnhw+zhMkqcoHViviqucuTizTPGr30pt01L
Pr4vFS39Ruythh3ii7uGQPS7/dJenQe9ArHG2jdeBeEpEoyt++nx+FuHWgEFuQif
pysepkDmHG4W/3RSQRPR1WWbV49aoUUkaiC/ZJ3+rgXzw8wTNr+Kx3FdZ9LOMzJN
t0GjgyWzfZ/6C0a8qM9d8Imw3hdU9QtmoAsGTClS/LGfq2d0z2JuBKRiyUIT+chr
iSRBLuxJCjM/dAOfM74kpXJ7Y331UIBTFdM0SZP2rL3CWKObhzQr/f+SXgAcZ1gb
E7tYaSfHlsFnawsPSD8p0CiUhP9u4nT9HYc4QYk8VG/ME86OkWoDjcClqMdUUCXR
NdtTQw8cXn0H/6hsvuUNSL4h91Jj6cAg0JYB9DEz6z0fbHz8st7Uu+m31m6iXBkP
1nOpB3sHEVzYQnILZeTQWwMETX7jqUe0hBlhCdlVvvaw/K1eOjramJtEGxF6gNEF
wACI+VFRq3mkJG59N/OCF58F/OpOw2H97hiXq72+h40yLOkFg1gxAz4P0NMQBQ2j
Stoyq4QHM4K7fPa2eAo5uKgi+yEUbWgPgxogMOpH1M4SJs3xysGq2/MHyEKyY+6C
sQvPQcY8lDJoOhx7Vt0JQeqSjgWJpL8ZXrwQEJgIK0fncLo0oLuQ7vgnAFzCY85X
aolK82pxBeUUrAApe3u0K+meNY84B1AFBQGY97XVr29WL6vjVg/Q4sQq938OUKdM
gQQ3F0jEpBn7X86eW6hys5aNYmIG4zwiXi24EdPhNmOkglJVH6UkPpQ34ki7Ldx0
6F/Rvp+ae8kb9+cstAdlTRYmC4vX/PBlli5huyBqRTe0WAHSUxyE7j20it4YVlWE
1+VkJAItGt1rmc/n00aQewKKm/KnffH3h4duuK+ilAr574u6xQDzgoLog36fPQ4N
qcHYZAoE5fRzas3Y1BVnZCuRZIbE6pG3JsFcY11ERKeNYaGt7pKo2ZJ/TUO8Pw1S
wH/7lCCr0v5Zu4Yr94bGmtS4mebYjyTk2pKiCY5TGldjdwrfX/5Ti8STG9TgoyKM
ELBXF13s36rLH8d7CafuYdilltYDPNLtu21sOlPtqkyDnu64dUZlIg2OsSa6TV3G
Ns5I879uc2dBeNfjwEAdSO117AQMxHC3/OwFSjuydjVnQOFSMhKU6JI1UgZ/+wxV
EBRy+oPLDZd0reOS4tXUS2DZuc/Slkb7BMqmMEJwiEQ8JUql2euI5aPtaJNRwpEp
3LV4s4Pp4mA6zw/RG+0s+TEzZMgCon+Pa9bNIhNLWahb0RSOQJGHK3+TSpiKLpmw
AkIzrC6dBGJJ3DEZBo2wexiwaA26j40mEEDkS3N9Snw7ACw5rPM4ZNrhl+WTnJFE
fbQPbOPyC+NbJ8TEwB0ZwX+SMAshiX7jM61x88fwp4uM7EsLGOCTdmyp9VbcZbsQ
a3Nh7/nwJFX6gaoYC7UB6U7Kh15zqa/lLzJUrwgRkmybSFsMlRBCopqAXg32gsHe
5syZZGgUU040rktyg5nK4h917fFVmCwphIe7q4wda9YbgfffYYEqP9fcLbgFmaER
74YdExT2580zE6BTBWVv3gTL5QCbVzAZZDmVWqHCQsA+lZKJT0b0jWVRAOVbQ/UD
kwFpBVi6Fpd/VnXzBZwZPOtXG8J2bWNa4ZV2X2zk6Ie0qJIzJjM7iY32qYmXIBVT
v9QCtgUBUxChSkljEVPffrO+MQhiY+kvmayaV9E3iBgborhBSLvpVAljgQWG6oyE
omm2AJD/mhhM89yrP++RBw==
`protect end_protected