`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11040 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhEl66vkmqNIpUVBO9a3D9esLFRfj9mQtc9u6h3NyKbnJ
5dMumn4FqlKv/kXo65d/L+dhWed6n7H4GAkPTS5C8kybYoonfuYMCf74LWmp/KJD
qrbSEynfd53lB4wLbv2Q3SCd7WRTKNhzMep+i72UWQGg5KytWy7luwcynT3nieAf
fM7JlIRXilpcNdxTsE6TEiSRHS6kXuFPSVGzfyqEtspa9gviAUVUHuHW6Ud4C2Gi
5jAOUNesowlYoSr1WyfmmC/BXxwvYNQTb8SUEPPAQHXFzujf8kNi/WD64BHq7l5F
pG923aWmGanrDRX5PELqsvkkF0P7kLqFAzlHlluHT/50juKWuyyYzt490s26UuZr
8YCYNxJFwwPtnmf9QD1vbz2WbP/B6Zi6DYHypex2cTOkbl2MPKHOKvsS6ZonMwEJ
kU7kvcf6bScRofVZUlbHdeMFsQQgbhN2xY3gsoDL7ReyGIeUxKL43o2qQebc48yw
2MeegtvFIQd5BQLL0X1xOAzYN9XaEXEn2ngoAQ47WAFSqdrGbyCwZOrqVJyinjpe
IUZzsSJbOXqYJfS9b2CiHWVs14MKGN+sBh9Vp+SN02hkUWHaMpD+XiGU/ZIIICML
w37Lphj/M3JwA6dN+fcZsnwQsqb5i0mxoKwsofl9w8BNspaLyoy4KESdUZBKYuF7
J8B2w/lVQjmna9k7rWoNyABlhxVlnlkqIRzBYJMwEWrN7ayGwnbKnDwTxU/egLGA
tpphekAJ9BhND9RqYpVqiZK6pFd3s/3rOW12JR/+w6DTNE1wxa8cP5zvgyzb03M/
SdbnUIjyF1daqPYdq8TzJc8k8CYU82fUbJXvAD8nA66fXXCfaT72Z3QGlWWh1CiC
ABXXH4rJTiEcVShUxpGNldZyjdlp2okWYB6ywNZ4gAQNYLEYua9CnurdsXFryCt8
qUB4dVlt3HfKspqfS41AMkgrOAJjTWsQzbyQO39+eG086Ve5bS7wE/7+9rvMMD3T
QCw1/M+/YvSwLjHfCeFSJSa6jvDLzePgkxVq6RXev1xZF4H0Z0lcbaHxbJ49rnI8
npRkYcDEsPGvZ21PguSUMBIyp3K4IYlwhel85jeLUjzR2MqWUN4ZAPRmjz1WHHgZ
8KpW/oCaGagURPPCdbXig87q1YfFXujgwXo0F6/MEmJgSqh1qOn8X8N7KWgBb+SO
73IlVrbCunmVc2QkrezbdYK/VS6AvwVj1MFWTXqRKOn224Tc3J4c/LNOFFtqUYsQ
ibRPZZZ68LZoPBMK0xn7qqkwHqTyJHYbJNbm1dO1AAofCmRkZGQYHWNtX+1rSAPA
OENCQjGiMrr9nczzzoIcjTw6ox5KNvSOrYjKn1ROHhO+DQ7GqOLh/ENR2G/bDjyc
iUkm3Drj6toDjMmpuEdhjZ8BA1xgTCqfUAina3ZPwECSGCWuBcBudepB4L+XoZhy
we/rWE1nvrNdzFP+07AhSU1a4XVRd7tpxiku1Xt9l28oTn6ZD1k5iI3U2flob/qo
i76PK/YbeMGPw2Tt2chvFIceXwF2+ICdYXbM5kddaiY1qe1nZDOsnHKmS28z+v73
OLxQT71F+jPAxod2jMuViYnCUNHS8yl/2Okg8RqwIMI80debu9PEF4fxyp6sVRm+
DsqH5JtembdcyGZhdPcnGbelA7+O/VMff+mU1+r5DM4T4Ab6UNrfc+jbjYmejenp
Mie+/NI9vak6t4mtQJgOwR06dMDH/m1b1qnLZlN4Virya7wnuBU1FoMISHJNSHhF
P4kYG1Qo44YO3uwq+u59hI/NU1bAIFyHDPaGblg5ea3vW0Y3Qclq06N4iG5YZfjP
ATjss7ledpJ11+8GOuZTM0Xuu7VrQAqp5VfUrgQIhrhtbnmYV0Ya2nZdEggh/fsI
urOg44QQIsh6zd9M2t6d01MDXMKosoBhGTF3TlnVvAZF+2Hm8AZFY9lDYfIi3sdE
I4OUkTMvlW0h8BWr84SHTIy/JZ3E6BeOLlvLuYZ3Cmxljod2BB2Kc6KxNeLe02BB
U/i0n6SPMVFGeEXLiTeqEc/pObKZUux4PMIDRbjWw3InlNRtg5cgZrNdHb1vD2EN
N7563e2B/LGDJ3I0itre8iA/gSmyNAolK5nPEQZVnbFrjPUbJujnTwhd9s8SJaVG
Z6sby+dUX51xjJuc3swunT1lLbyjVVq8XnZulH9G6NYNWpRc43QfnZZ70LgLMNGZ
nLr7X+IOwqjxgq0uudus06MQ+FKziXazLaoVKwXEIzw0oytBGqFVlGWtuoWicbBE
n4UaxXc5mUVTGX1+7G+ns5jnYGX7IuEJpcfKpUbmhv1/3qrhGigP+XK4kbmdRmXL
lgvW7HxGhBB2Dpp1xl5uAHFwyWjYFT33YTMFT2i4tDLwn/ZtmhCCV5DF4+TkTn0c
GizdUMKLji0CSwa9SbOtuOymz/JrIFCB5FGPVooGWVkS2aRfmT6Ko81Myo2iqThv
HF8hUWZbY87Cr/YBFsnOqwdHH77G5isOOeHXPyovpBYgx4v742K0oZO8ybxeaEud
UZgzswwU9NAcVQq3z+y6QY15q0Z0UOHcOf/j/jkp0jLcJMW2WKl/joP22dkyI6fW
a1yfN35F2faI8nc35NGQsH6iFDyMTxcEl6KX8Z7pYdB2+SuIzE7wbRgDyUq68Co6
70qGVgdHLh+g2en8/7jUEPK10J+eyOel7dHXLpwfSRCgXGSSEOfP8iu68BUdVYM0
Gy+bMma0+NRv+s01A3LJ3QWimVsM3YSfE4FS9W9lX8n2TqZWLtPfSMEWZ98AW7g4
NHeYz0yqpYQgAkfIzxed4SXPsTA0Q9Y3BRb9hrYLSgMFLsj5hWvkr5xiPrGxmBch
jGoYjiB7KS9HuR2JIaQvWTgM8v1vnVInGp5/V/wFtJW4TQBJhgareYFnTpQMPFCh
+h5neMZ0KrhAMP5U6n2/Q15usFJgujUv3pOp0IDs+pr9L2k2TzXYYLXTV7KCdk1C
CbMZ/SaDLpWhCMtCvGVQ3Xciavyu22dIF0g93+tOCi2PVKNy1xLuXliIW2UE1JCq
an5JSlGejCmzHG99Ku7EH1yXRl8HlMkQ0LuTq2A4DiEcM2N1qInjctCF2pDGYcuj
tYOaOe8oF1VL091eo9a0ECmOJ9E4V2adrgFx7TswPHztmez0ZnSdNUEbT3ZYBPeo
e9/zKbn+NKwMKipT2vvjD6G8x9e8AFyhXTZwG0+nY45ZYGlr8PsI5ywNIHVYTW5o
zPFIPyfz+LfoOQkFPJRB9/Sup+V3HI/Y/7CGXhQ9E5T9x5vS2msLGhJARlPclKPE
FQN2CSGNDLKRbsj6lqDVVncW1P6dRMUI3pJrKX64G2TYB+yZmUWC4/on2pGhRlXh
7hS7ZGA/vafwd/ba9AstPogtp+gNCBPy/U5RilSRTran8oCIFYjV650IpEFv9ybh
QBicQYhEJH+mVLj7sNL/jbWpH13HpE1zXWhygjCujkc3yDoaIxJccb40eZPYnCey
FinTvyCKGz1i86wfvz21ajriNqgsgofWZkSEVlrW48z9qtp/2xCX/vgzqUT3Tx0I
EqdefOMwOJWb5kzkksPzyqsTX2Xa2QB0N3x5j8ByOwgwCEZv/K1mDh4U/VjEvIWL
d9hp1Tuh+WgBnlDN6jdyM16P4XXGdM/L9qCusVuN21mEoWQKkFwAhVNcg5mDH3VZ
qmfXS/LuWn/GVF1OXTy39lPgB54e+/8yPGMUd+G5LzZtNpDQT6YLUQpI3KhqZs6n
kFYCyBnbMjNXoG+B8Hbgu+3VdrT2qJ/gF6eGx2zhvdPUJVgv4q8z44n8cXAjZqGA
j2JCih6SQqX2MEgBpsrSUma1oF9ZYNClAUuiPSuCgVVmXjcJzyiF6c8w3sLv67zH
PGbZ+udc/reQDrr1b0cNmcDj7q326jK/GAHdHf7pAvIt2AHEBKmm3rUZG6Jwnp1d
3SJRCJ41fB7qQ3Et7OjaI/4ybgRQM7rrxUm0mTcsJ0SrvAxxVUEcXkc3LCai4/pd
zdP6hZmS2r42FBRSLCV73aQXRPhGGFi6Cl3txU2q4NY4JSIuhWRagTYOvNBIvkeG
dhisKnTFqK8DSZlIshO2DNxVvMn7I6NamW4UAtd3uD4+W+q/WjN0UtX1Hg9Y7cDc
Bi18HqRO29lGqAloVhnefZgUxeITeI+szKlNXnGLSZGDSFMggZfcHg6PA2Oz0Zvy
aFDZeFCLg1bKpejPTACF4QGvGK/6MkdFoeLzh86KFRVnKGzfTl98O0WwvZiI8C0d
s+mDeKvobvYpqHhQHxg3KKyCs4JOqZ9tvx3cOdfzmO054HkW0WPvR8CNRGeqe2gi
pUIaWjUigwEac+MBm15dI4rPmSH6SmKiazvVzZ2Lr8FDWbCit+0h7+XenedNZ3Vq
+byD0MRXWmxXG7LOtyLRA6ESzfaxcDvS/hMzwfHobY51ilystSqo8G8bqMLkEZfM
5h/MJDOsU3RSQbDscclNyiuPc0qsLspaZqzb8D8KSP+gYS3bnws+Tqihtg6ejihz
cZMsWiBX8qDt6erowKtzLLHMMI8Fm2mebkQdTghLPpH9/NA3DkmbLEks2+gbMZn2
lp34IMgHpCLT10Zk4fuy8W8zFooNlJfZgQ7a/4z3F4bH3oyM3aNI2eAhOhKxN3TO
VR7FOWzufNR6kOO7NLgrMMaRiSC7y6o+QugP8JCxqF7I33TLS1WmC59YlKrXkxiO
owXlPipt9M7Noy7hvi4De2RL0n/JT01SBGyjvcfDNZ4sHlLZQu3DHbXg+jsfg1lj
8pZ7lpifny4OpjTN5t9E29ur0nLd7Nz38Q5FPr07p0l1KQls3DKLqD7RnXzJgqNT
G0+iYYUqOb3vqcpQmzVJ/v7qfE7Hy+vVjntXbbzi4fL5QdGX8Vz/KYJGqUodVx7Q
ZYawq6H+F5EYEiaTFI2e07NmOvN5vakk0PNyyWE1BO8EugTS8FQT5bShAlA4RRD1
fdkHGTgq+gGIY+BB7ZBCzqZPBBuF3bwgFlLEW9KZ22i1wHfLKr3Pz7D3Fr7a1Shy
Z/h5RNfkL1uFof/QXaG4vcSt4Ow2l2l2vDT/TO1U/i6joQMfQx7ZbYLT8KCPvPEI
KftQsCQasUXRxM6Lv0CS4yzYEnizwzKSStqfCoGAXueNy/JZpESTksQ5849HA/Cp
ZrYGq/PHQ2LMGeLeiLrYUQLFpi1/FImnOQhfxZ15KbSoEPDtqBWRxSUKh3vQ/uVf
Udah5rOCVYFTEmo8dYgjxSa+X858y3SbcnKCJbRQns48kYNQxRB1bbL/HSvYyaga
Wk+NFoFc+FM7/st2i7i72SvHILrXvaEoalRXqNV+pFaie5mMsNz4dHWSkf98q+sY
w/QjXNSLcVKKkYmPBc7N/ihjqqQyaob+dM6Lum7rVnjS3x3orKJ3pUin8RsbyHYH
KqBM4bjjFZX1RoOK0/saXwBnlqsuOSj17N4bh11Eh7i9oJ2X56koYFJBVNPlMpt2
nkcZ1zn8TvjJLoU6FZkHs8G6TZvTz9T4vm33kGNz3KC/5LcCGGYezd/KuvqcWkNS
E97AhqEQ/ZWrgVMxPIjUCXq8FWHdCCQUAL4jFFHlEViJQzZ3C7BsyPacv7vnxqg9
txGIKy5brwr06ntnd3EHkrN/WVSdb/v3nlmyEwClNsZl21/6uZS6lT6N3p55KXG2
dBUWxa0jxRItZcBKD2BAYcsnrCRDOH6HQtC5suE+higX859mZWVtdW9YnFVPaHQJ
gYqP77riOf70PQs+XiB/tAjGFFsbO60S5/u7rsq5P107vx3kIBXEULF8HkC/XqqD
6EOuJp/DbfA88U22+aPDwWrudMKMFYnIueweRgbk1O2Vw4u1I33htqtyzI9PXs0V
HPpSgsdHp/aNas/rOoZq73XeQQVYTbzaVuf0zwH6bWHYMJhogy4qzyEic8TQlwbr
oqq3renWxBvbtTMF7Afblh6UVN9kAXwOvJ+vHPAF41UmKPinxpxePFixky/7Nex4
zZHUGEEEF2nbULxKAXuEDTuHyUqgLXCHt04Z/MjCwuov9s7HBfsqwXo3pES2yr4p
eRyIDRfp5p4txBZPBhGcZkjnazTA30GpSfULs7fi+ShgrFCoVwTs7L1vvvEDKeeK
+xPVW5BueXBZ/pUEDa1/HiCVBTcBhn97N02RxQDmiqykZGaP7ZEHL+gnXH8jgrqQ
D5Ajl83y2eLI4JpAPSHj3ZG1qgI964i3m+uEDPqBYIFkPpBTZeX54+JCupRuaKhd
0FwsT7BkchP8Mr9ow4zeuxnN1O+3Clxv9X6uD9DnVVSp713AwKHDI7S3NnZmz4bW
21rBXpzXWJtBwtt57f4mM6lXAdMA+ADA3GUuxmQnymSWDc4FcHb7jxo9vpYAsbaN
WYdKqrsnv1Zg3GqjGzwBSKgZydXasdv+GTQlF1Lj2OiruOVDevZY2/FM0q1+dnqo
ggUspkT8UtZKttMZr9meu2pax5Uc86Unf7s4PRVN2qnjj+MxjhEbGhaKQK7yLdje
DgsSDSPWYB+07z0/piojBpkZT0S27F8kKYVQvi/Ch06LRkLLRvg2rI3ojGdJs9ww
DLkGBzlNHZ9mKPhY+XHRGLTejWBhfBS+lMXEFzQemuvK2+yi0mTdoOBqMiWgCMcU
6Hc5d/A+0wxcGBYZzgB8rSXjKV6W9xrAvi95TudqzCxn9knz9vIzEP2hLwMB3qTY
tt3IzHY0mApcP4X5aI7kdCY0jCcGu3w8hw2tOiWipSsJsJqzEnA/m6G5QEhDWAMa
ocH0vNbBxoho4sr4VE3vkw/zPuvIhFDan4Du/2JsZkykZLyMfy3cZrg+FiJBd12o
UB2HA7UZdU0KXRNlhFMSg44rCeqROZzLd8fdNHRMgynowDWyQjJRj44chFrpJAzS
km3gLHrRcct9c2ycOwZ3AVPzSWZNqj+A4tZxp02d4L5x4OLhBLrMpz/dSn2DrzSo
YEr2vyZSR9Bhqdt94BNLCf2/4DXyRy7SjK/wkOuk3zMagH5g276Z39D0zISTwdQN
Tuwx5CYy9Uk3UOOucuX9zrD2aPS19nRLmO80rab+YACHS9HUNI6Ax8K7ilqzfrNV
rp+CXnStx545f0LQ67lAkpy0c9cJ5cve7KjWr7sMqpF6yXRNrY2QHa7l5tQ14Ods
tmYXLEet4bkEiLPPc2G3I1SJKAZgs6Po0/PkVrKFtrtClPauxpNghxV4zc6MKAQi
wXBf+7X1SoFXdTpjYGB73cUZKWa4ekh16y4PzJlM8LGAO++rmNp0l5pC8ZXZsnTs
u7ZnXYbmtcqSU/CBNblxcHX9RfH92J5zi5xINFvR7lvQiy8NZLFdndrvL1gPLVGj
EHQvlXFKPWaJZ9/BnlHqGjoEcy5lyMofaJAubtmGAOk59ETmfUIU7sONlmHjoLll
NlAwsLa/DmM7S8GYuQJS5eHUuMDnAHAKFYOn8yeONpf/Aj5zAwyrfzsVTiiiOcfH
ts/MxqB88QBFS890+Nqwgv9t57nOvJmfhAyvOjJKGt8z5R/qiT/gTU8u1/bxTPX5
wQyciNW0GRQmhwNRKV0JIbx9oHKlt7tezWb9kqqP4uC530b84GavjvwbtEDQ2sw9
h+oPoXn49gDj6KB41A6VSPF7cTDpBx8QGcfCu3+IRiSgJyMFYh/bdgRflj4FB9Qx
iCUfx0ljYFdl5cldXWD6f3HadtHYIvUkA2tu7XAtX+IECotvOP9HjYqB4fWFPRiE
oUgIG307n/NSubMHY+Kj/qaNkJfVuhDgEP/rkPkAtHXNKRJZ07gkL7MtJFKedONw
vamJNPVQP3XFIzCh9VK0UL0ICtUYVZOg5wPVbTToIOHLe8iOm6/x/fQt2s0mkK7z
/CggrEFFTEytEi7uOgFZQhTrKGLSGyqjmT1VwThs147A4E9OSWVsdXYKY36qTjNQ
b8R5wzyH/gS9HQbsOFxP0hF9OTPhV+Luuq9QlVxT9xJ22AnBPp63bpDzQhIp8sbT
mbWqrEeRh30C/YLMpoWdSgnQjytM6WVOs5WscfiegDK3uQ9+veGjvmv9thGzm5MB
Wz764LhTbTIzxxhLw93UF+xLDikcL7RTaYKfozrMmyD/vBAuGdPk77Utfuz0fUOP
xRcVOzvn2yfNjwuh7hVWyoaTTHQkEWzbRYmO/u0GM5y23pLaPR89gjbbWILd7DKz
KF4GeOLup2+RuePw1zTy4Cfgb6cTouW9UqDFqVT20lbTr6C7t+dZOvLkYUd9FWkH
kW5Ej9DlYOhy/wmEFTD68vhI6mNlDSGgn3eJWqW0S9XNI+yJv55XhS9eLeDCv566
CkaLuywkr1XqP7gKbt4VloXZHC9/76KMokCcLApBJ1pyXxn8ZvVSkqeDg0dTJ2OW
1CBJopDpC06q4sTt5HC6euN8EpokbVU76Ed847//zD/SPnmEO8sN5kg47qJvb7eW
p07IanYoHNp4XfozX1z7MUbB2Vc13XTIW75Tr8TuQZnYVrupf2RO7MMG+4Sg859e
0W4Lwqr8Ig65s3hemZXr6QH6b87g6v6qqEpZYxwU7cqxFPg3VIGW/UGVYXLwLNRC
V+6UE87J1doVUXTdb5UCP8tJ4Sjx/0Pmv0GheYk+qVc3FYi8Zo4euFpXlBlYyAhJ
+HpG/1Yf4KFcDVaiMeA+KQSXNfLj97eV3GTSGt1pDC+Zrtt3M2Cr4fHHEK99svoE
55tLBvt1w1su4JajthDHFYDccpFEK+nuDoUJ9PS2q/7pefvdDtSrm8dmcqefsQK4
VabJJS7jieSCxXnJm0aYZjdglwbkcc2s2RLW1UiseF/yOGFoyuAh7qcdwiQ/MfYn
GQ+usnJmY89fzSzaDpzlT7SrZ3pCyRnpNBFkWKsGGLVt7y3T8bmuD+bJtfOo3zsY
ldgvLeZUfswjJLvDpYOjmTuFwv0+7m6HLoyuFRvJ9/8WSgWV7jxJ96YT2OJvBx3/
RG04qVZpgrOHthYSjlqv6avOXT9wibl1VGqK9M9Gp5iHw8IeesWGH14b1p8YUMFc
2RHtzrY9XGe2AiWJlUDFk0sjowihTq4/J+EOHMCLQ6KItEYz+bRZLcN3yZJyVzRR
6NguWEjU/UfT5bLsovwxEt11/gM6Eesqv/C5JOr3l55Rc8EbTjZuSZZ4Q69ggE+B
+wgYVyLCdUDRBBpyvkCmnBdA9Gk4lH+rNAvhU49G0SsXViQqKJ4AfWj9oE5NYVCq
eUucYB3hK2LOCmJoMhTr0hq1l5II0/V7lOcDOkxS7PwgbP1KToY2XQBGfMqRe8TQ
zG4qWvGNg8MZfZNZuj2H4+TD15uLHs7WIHl6g0/NQVa/qqfZdupibTZYkSNkNoDm
bFYmIsjSIIljOOQ+ZMr29YCW8Pd2X1GnceOzpLEn/IZUa+EwExOsjEqiA9j4iqpl
b33k9gIXqv2e2hH7Akv5bOqsZvsOgtE5Z8ISiTCwudG9kUQgfbNoN+CAfs8c6evp
7F+9yiyJ31BrzABJdAyaUki609UWauG6E8bNV2TFGRkpFVP7KPCe+mbi5fCWuFts
XMnjCti7iBnw339gTKlBZrYHhxLePeH39I/HRFoV1ISDTanYvgUr5yiWEcZglaIL
UgoWsBiUyfIThSZJoAQ7OwaHPAUatm1gOHLTKLvihzEMyKbAkbNAUpKU0rqfWq2F
NIAdujK+nf66B0BjFCyrUEGU0VPpoq1e4GFoxXUW0RcPDweadFoXQWnWmiYRzx8O
T8h9QnmK+WNhau28A90BmyZBKxqbePFByUZ5XVwKBXUB8DZ/49GlBVH+oiTap/tQ
KeOyGE6RzuPhgzpWhl4kkq+42MTkkS0Gdz7HANQgyfxH1AzpmpG2K0Gzc9x0Svvy
cz81JIgKkVR4A1/356Or+t5AsG77HEenJkR5WhgrVRGMuS+5D3hQT2bIpp6haG8z
b1qjCUyePtDitcg7fBpyHwagLm/6T/kKrVivjBQdwQ5KFodRhYQZwrMErH55Ruqe
6J0gK5peRnxMryoEXa9RajD6jNHi+qGRq+bLAC3r+Wuuv1gkb7frPwtvvvtbaOdC
CLzTIPdEmV43oKlozZ57fYowb1wA4LNbDuLPNQvBOMrSqooKcfLFDQmIbMFL+YwW
QGbtHFjLZAJM6ex+NNO+tAqCTDrK9mtqf5jCeJKIhm6XNad3zjf77pck1h1adhZe
jBSkfzvu5VBywSQlU3ldM7ml3bTOBenfz1nhqcBYDzVzZZv4fo2DSKOv7gDDs9dX
s7k6GtKINQN0m0kVACv7Rt00YJFQIaUWC5+MbbpuLaoHR3FwCNzvec+5HKXzwY94
Oq1gOmwI2fCvAhLyGPF9lTY0xrhjgpfZOZCutwki/ZfAMi5FjIvJSRBbexjoySJu
JEVXYltHOGuKeWHzJDLovTs8+0HHf6RepK4SSeXSGi8+Vux2K1n1E8O8KYC1/H8W
QQEnV9sQFkDCbcKsGHcnRTi0nT1ZrGur/ydAgq37ICjbPbbSZFU6ePoOu3ZuTSI+
zrv9yMKhnUrMg0Of10MrW3FqLRc2LHPZjSqDGwaA4cmwZhAxk5dIY4BhYhAMMasK
SoQ4pOg94D4CfSy5mxeFpJm0AMbU0k7tWnrOXEjML57NeJRsCIqfrQFZFqqfO1gX
vwszpg3/TL545ExQz3c9jxg+HuIYMNx3UqZC5g3mgFOfAIfoNcJ4lOVBuyJ77Gyq
W7rhMigxj9c/TESWxINbyJvesjzqOzMjpok0RzYcKXS89qLgcdvIPKj9HBwctran
2sO1+76fuwmOGDSbrGw3Br8/4LvCr7JrgImyCFLMlUxY750ZiizXuadvuuPyVRHz
8T7SPrnFa2mLtoIkhP8dGMxs68DndZOhpxTXbcdEtd3ICVKWeqx+RYvRbk2vDZ2v
hhnUOAmM4JSxevMXTRHywMQ3EB/fePPGiFSDSkHmzCLiJmklHSiwC2SXqki0WLog
9g5pRwEo9H5ncaKIHDkN7SNzhSu0dNHRz2IGFdKRd6fhqJMO+KjOiflpRU6KqR9l
r36W922qHGTCvuiuln9MHVKgaPic3yOgAuNXMTqUmvhlMkQkNE6veVQQyLJwpmcm
FoHysgzuiMWWIOJeK7JofmzP+/uzcYvk0lXCIvFhrLprdYE4n3Y1DUolEYbHFB1C
Vzz+Ly3UyQit94Af5E4EdwQ5KuBZba8mrgabeV0JGMhscy1o98ln/axyUWbxK/rw
1McD4oZ4LdnQCZzuPFLe4ZYG4ZrPkWK5uygh2+NSmq9fLV/vfTnPUCGM3CL4NeSk
XzOTSfCWyTUpxl97jrPuQ6smlikfNvZSocvhZ3WdL46M/DgF8EZnQtVds2NVl16X
14o+sWMnkvsFjU/XEYSBix7eqrEqm3oI/lH/7oultMk+WITZo+CO88JnWJ/RtF8W
VM+l+1I1YS+KsSUYz5b7wmvhMslb4GOjSnVO9hMhP6h0ef2uclCR6MzGl+45BWwm
fouRUgRxs08TgT66YSofruVDNyhj9C6X5/pTEQyrPGSpOQSOwchyUynYXcMC7H9U
+ZT7J/fzrXPJwXJWj7CSXzsMg1wOfiTzlvcRSwl+hePW8G/PkFTo9Hsf78mBaNB7
6aOE3zgypbtFnhZohgO/aIKJDY/cuM5W16Av3Yijg8RSZDwuOr9HOYYGezzSjJXm
tl3uMPdmG5TGI8yyeL7FWhwOO4laxO1BIy6YQxa6VqJF4Z3yUbIUjWSxMO6HaX1o
O0jbedtrVtVyE7lsmM3fE+9PnZI4Bm9Zu6WcIA8mTysV0EAVf4TW/qR6QSYVuxUV
JzjNylfo6PzkuodMvcIEHygphggvCegETHcm0ZVcQJ0FAO6V/0Xba+uNwrdq6Pv2
jHUa+RWCfwotEgKxOdvC0NBMHGasjAzlV5aYE/si4tZKGkuCqjKZSR+Gk1ILo+Uk
AZzq1SO39Amlfsa9Xd++Me8IwyJRqxYpnszROU49lGSFm4Q3E8QlsPvPnRP/K6a+
wnr84/Fx5vyfq5d2oOw031lmIlHKC3iKgeJss9tMynkjcsS60fCj1eQs7vZwcJW2
t3jesWy2cZ7/IucTipsV4It+3S4IUO3GnTKaxYlcTjQm1qCMpIt3LEYZ2iYk/U2z
Oa+wp9ExCsCw1cREi4ItlHnKNnWnNYVRKcgtna60ziIbCperFFd0XbaszCwvgqXZ
PJ2UXU29rbLYpPcgMbU+zptn8QHwwvqtjgtBgFxhXQwIolpAeSwpERgq+Ysn5jmW
GhIPvLjYgSwQ/KbRYDYiONbwIGA9AILUYV+/bDHl7jYyNGJaDv3dWHnQ4E/pGtfv
cXHVr2sLhRj1U48W0w6hgPLLCUchL/FOTlMx6R3FTxnCxp8LkgRHMLUdgvYCyO3W
Dv1w5JaQwV1PnMuiTAViPbGMgive2dtY3rx+CM5GwIIn7G4FOANWbKaCED8SJhik
T6KyTjXC+JkJ6PAPX6AAk7ClAlmy266ynTIyDJwp/jFVagE88mnHBe32wBgaO2Hi
zbTpeF4t3qhc2bejrLcGV3gYHVxiSmMtRqavQv95paMZHhaKgnWHDrslUaWCaDlb
SuhmOPsrNMEhNu7WXqtK7LTqHaDO0FV0Bq3gBjSG4baBi1HXAIlzvIW3GQ6ZWAQe
13COOpSNF9rqcB/+cRjNbRtuHW8Z3HToeDg/OMsg0VJKtPVTDeYD/Dj0xIry4gGB
o2d0WUsladp0RB/SFsWs7zK/1Kbl5lGqLTmGsWexpG7XDoTuhRwKdDT/ewk79gwc
v0qF73wIjPoVSiqkOQfso7C1MRmfUp6nQXZcSiHlqQ0Pfcq8wDnS0v+znA7LOjFs
EkdrQoebtThmeRQ03X3iReEU+c2lPE+NeFwEULPnCOuIGfXRp3MK34CNE3+dal1Z
wzUk1wxPJJmVuS9rXxoXDMnbWs1yazsQbUEHe8JS7tNgdOtkXyaWERt6i2Qf7q4p
Co2jzyB0FebkIIb0nvDE9+am3wGlbmtvREsZZLM1MkpGG45lsLWkGBs2qqGil0B+
xVgBCyo5OGQRbyzGSAtT3xy7FpGEQiqVIJuHHZkAdXYXHI1wKqqWunIGhJwgd0pM
4EbjRiQo823i5mFz4gWUodx5o/0D6qDRIE3xBHjvD2YypChZ5BFVHs5QQVSupdSO
NGGvbscUqsK3W54DPONffkzQ7lKfiW3TuK6b4jZkSORE4xlsLtF4ndZZIxhXRPTz
ieDylWBoh+EaN0eWaA/oD3rLKztYQcrOwc85D8iWg1JbewZhEIR5leCLfECV/aeO
Hr7OlRqaZDT5MKLPUF+AUmvcWC3i7CCtnrv2ZxkuVUi/rCXGbEGjMeOSSiuziAra
9tYuAiK3MZKGNXJ0kZinDdVMzoqJKW+wrqKZTG+Yw/Ay4OJ0RAWJSfppbdrF+SEL
y1e6JGz72CzBqFZ91VY1e7kAzjp32EBKhxGDYGSEyHzT7rfI/AVHfNZE8TiVKE4X
CukBPclVxHk8KicH/DdMd7QwOJwgEYjtrmr4xSXp2uhIC3ryPsLYwpJVewB/L1i9
TP+02qff4DCpwZgYvoVFHYfbona9J/h1J8fLDjMTUhIdqQTQUsgR6A1h07Yjevls
gC+ttiUBD6hCj/kSH9eqKWWT2Hkf52Ibo1n1yfRwXj8UgHblxTZdTjI/PS1kSB9c
VppYXqAuytzaL+1dl+OQIU+yuBVS5uKubsRATc821YozvZbOmXuZUM4nMTPm0KAY
ShHdXIjyHKQxsHMZscOlQvJ0byXytrPVKE0GBSwR2gNAZLkXu4YJi9qoKNMtxwbg
J1L6MqETmTjr7Rpm6erzXnIOCoeMdW6ccW4Vn7od627G5U4yowXs4CL40uUHPDat
AyZr/3GnOZwP/gI0y+ylWee3K6pnKtRoLCrl09viuO7w9iLC4QFQb3mmo3VZtsBp
WnQS0M3XTVo8ypKPqjlAbWdEbMEE0A/mHrS7b2lDC9ofyFqp2inbxqSoibKCC/ei
BpS9L8UOjSHoCT9rXEJLAazzXMihT4Z/H+pl76EBwikAIjk71Qss53gTe5zQyaBy
fzcISES5aqAw8qDmSHg26ltMP8GuUKuMt12uig45ueyNHnIdqyxc/E1DPQwZvNp+
pYI5wZHNC0FJBHr1Qu5F+FJE5MTe3NIC7N9BsxQP2TpjSCFa11fsrRY/TNL/xFC8
6QixraFlXFkOC+mklU/A4z/Mh90usXYcZ9B0/mi+Nas96ZNPPYEI8qSMpXq67poc
oZfMwHgvZ6WiK2/9Tcine0vAWIqr6b9cVo4uwxy0RUzoRiMK+UNeybY/ruD2+FUM
BdQleWKUm5pUMam1Q1q/tKJQ/PtIlPJOMpZVwU+DllgfyyzpnPeVm9SB1Q+rZYA0
uVhN443u7JaL5KaGqaY/yzf48E1+SKf+/wnf7ud6bh64M/xOBl02baQMc+2212tJ
2zTYPNISx9tQMcCdbOfDIGvBsJzBmjGDsBerIhb5HkCeH6NJHPL3vWCsla4XyYT7
85yHcAlUbFBqpPaqm5pj8oWkXJuTzohKG9XxVmLGWaR1aUUjBgAObsAt9o5SRwKt
K4pCwMQIK5PGWf7/97mFXFt2PL4f2iFxPzUZGsFK5xKAJZWDKxVITcAPE9m+Ks1Y
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11040 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/T97rZhQva68T7JOm4bkq25
b4BW57ADAHEm2yg/Vzsfl3PNZ0qsJqYKXh6pVrKzRkedl/wD+idrAnrENlDLqBw3
ekNML55I7W3YDV6oivCFYwBlfm1UZEUiSnYGKUktxe58n7oqZT8NryCi/gTw+ins
qApO0E4vaFu+RXM2fCbWpHBW7TPweGNzioUvTYNzmgvfPjTjlBw39GMHxwcFvCrN
2obtgamVyUG4dYn5uBCt0jW8+9yQLUL5/2x56S51+3zkA/8HUS0f6lLMrbpvdR4i
foBp+aY/Mk+TzH+W73RrOKJ3uPpWcdGVufvG2nqF+f5EBX7X1L+DQfa87lH0pfCv
dC6vsvj5c2iZJYf9nMSfygJLMrRiaOPBBYKoiQ1j0e1bTgqleeU59M3w3hwd0D9W
9iwz2PhWT+kTYLlCpajHb4Ciq8oABqqEA3nEHiggA2T98P/C1RT9yLsinjOiRSj+
FjUmN1UEh3/XppTtz9Z1xZikoPBrPH1Ejf8mfuzSkCpdTuUsvnEAalQZoEfJNb26
Lt94qdeTQosI/h8dn6vrluwezu4nK6S7bNEQRo0+chXXm4kVC9rMlAIzBm0EIako
3ZEUlpwjXC5YxU2sxTQjR8LXLOkX2Uw7Y3IGQY9CXtobfRKwY0BQzHjCBoIk/480
ZStpPrLx95upC/sJixuwDoc5gEO0Sfic+nCvy7oM3+UwPhu5jcgcwF2COxKmwKiY
QQkM3DEd/6jOfFpttJZs2w55K7Xk7itUIPL9EvdRVMvMaAmPU93PMEE9+7I2C3WP
vgaHHG0tkUNEuQQbDK6zza64VE0M+eiEu+CbCI4QpEOHO8CAnY9K8915ICz+x6zT
67LONHd3cZILKsC0U1Xm2SWcx23xS9WUMG890h5biI1gjEo3eoLhEl+109k1xaH2
IaldlWgniLZ2HXxR2Uc/36Z0agR69FkK1GWPMRq54CCacPl5sN55UL2MfnfENTuk
FRfnMNC83Fa4umTbVtWhCRMDaPp1pFJU1asogul8p89zZlfH//8iC4M+lCiK4/U+
FFuTzFmEkPJDaST4cqfFtPd35t0Tm3OIpHMzsdWMe35wF/dE7tRsba5xXR7oHDWA
PgDi4iec4D36YyTH1/+mBV72rVL4d30khyWYU2PZIBqCw2jWZdbSyuDoiDFGH81E
Ngsba3mz5qrJgZLq0co5V/c6YwzqROxnqRY+Gnp5v/5DfmJkrzQAj99428/+APV2
wVeLdTJ0YlN+mLXSv2CYfqUOQN/AVFsFi61D2siC8usqXjwuIT905cJKh4PqGvxb
I2COeluDOOuWi0G02TxIMj9AU5gEW3HsPVSWQ9NtsqfaXBtSFfp9eOOdbtYrkXeM
Z9vHorIZQ5YhK+KCky0qJMWTp6X7tcMH8jYIxaFluy1+ChsGnTV3a0o+V0wxyozJ
Wsk9LdaIsK1vIHd48337BYyv2be9+iFyRwlagO6ZXyjqa6Y0AUrO7lkN1LFDD0cX
WAzCh5nfNnO0Kg/vaipTyTmqebhLhQjcHuHcVIY3O4sOhEx7B6f1wM8RPRKOX5lt
O2/FJ4aUdXfERdHkVpl/PEN0NgQtRs5ulc832mbxwLvKWHWvYAbOPyskEmzzEOGS
UKJsmdydPPO8o4bK7if9g1btDc7eypZSqBHKy9WfY3HfzJDPuzH9697CP6Je+Sua
V5646h0KqSDQfgfL1UUeWeaWBYR1lS+C3J1TG//vR5cP9bGbchpAVcD+mUJVnAfz
UHGAQ2E4dLY74/+KyoQ5KQd8MCMu9IM6ExH3OSF6yQiLeHpYFvHUVnt/uXblwOWi
5D31kwsTj0yozzqV4Ae/5YwDMneLYRXLZavZuJHtKnxia1fsYNr9QXcBygJjE+A8
+R7nRuyNXhY96QyqfZWD2JR7UY7fN/x3lHYdjaLOkar8gr4WErPwaq+5tuCSHxbe
ChtzUrN/seB5ByYyg7fKJkfS+hUNZPWhLq6LcCdbsVhHhFLsw6qQaWDHLJS3Ghm7
eDa0xzkQExkViR5lwBtRRn2+HyfJaOaaytpKCgvvwAGS+1kz1QAsrq4ZBedNS6Xh
bnhr3tYIH+vqr3Qr1JW4Y4L7KWijOWR8owanCQQAMstyAdWQiP+BjhRk/eUy7vg8
IywIjyY0dkFWpc9eO/SqeBfO/kT3KiA0jKxhyJo2qiynwpSvh28Ke55xmDpoBcNI
l8F9V49I9OwmEU1zOR5nxfwLwLZ2tQdovWvRT5/RqZrrKyibad92+mMqoonbyA9O
dSRfpimpggskKSPH+93Y+sKojQNmjp2PS1a/GqhVcl8P57HbPRSPT4WCVZ64J3eI
9OfvQsDkiS/twDT7Wy9liXS/7KaFP9Tme7u88WZlG1D2U/qG26W+6QPTO5rB3UPv
fVlX0P6L3/MaMttFqlQkqeN+XI2SHjTbT6TeuR95ZMWlAZb+wlY/3RjcGTakymy/
WvI4C+KDpKqbU/l8ta9OVfjmwH2/zKcG63q8d/oTR7PcZoSh1Gd9ZFFndhUH6usZ
4bkIPrWmknvpXwSb4Sxv6SyCVdzDiDOBqswKmygUdCvDWRO0INfZXmC11rWIRHZa
d588lKo95xW5O7oOkmRGN1Vwjdqq1ptrEvxwpgxypthIq3flPA9LdApMprhkq5rm
XjYX/FW/u45DGYE17sR6K3CoHDizIg+y5GHPYV7Y5Npyz+h6VydJ4+H5GmO50QRU
mhQE3esv50uCexrw35RjDD+vbfy3aAH1WcaRaVwfcmS6wmwB1mZsaWTmnr0whT9Q
HchoN/SXwrPJdeAry/bK6RSr4i41WOpSXFLPFYttJAy5ikiTKgRb0F7D6xbgbLhF
pjMQz3UpJK2m8kpKaotOlF+i4ggD/ZmThvERvnhafWmNSFS9ujrfW7G8ccWQctqq
NfOZnchmCpHHeZKHZrezOxbYsv8PCaOLpJkj3cMtTYdZsoPWsNVq7KSlaMx9DeL0
2fV39vM79SL6dW4eqEokk3Y4M/hIUd692Edbn1yVVCa/B15ixm2mOu7Flg/kJThf
J4u78Cd6Huo6ULURu6SxrUqRXnqqFiDGr6nlYiwHPrYkYFJ6lXLtXY/VSatAC7y9
bxFSF+n7QElzArqhd9QXzVsWYpA1DAGmBsdZ4LsZzjeHykdDQ9S26nyoB2MfgROK
mdcT69EsoI4MNOcB+MvVnMbCjZRiJ93UXyPlSE7YIlAnW5+YFEXfofYVGGDMJt5J
FvUTzu6uDZIOtl0lSf9W0fctfvBc3/F6UogUStUg1EhD0IOn9tjQh8eo2uyTgfx+
tKpYdQUIOXynS+9LM6u6+YUam5AocTSRBLrIRxf4RpVlgKR3f2JI37pzj3n7i+HM
PQiswgzG/H5ottKtyAmL2emk9bCEu7Kjaxajf1YZusplN21RNCIrxcI/nSO859Wa
/KEN4n0M8kcZPt3pLuN0RdmW10rkrGWZSz2YXEil3Lk5Viu0hOW+hSG0mknc18Xt
zkOINndPg4UxK9dfX5HASXabcpOktj3jYPIxuUXl7BjcvBmHvTIH7Aq5arLFJf7g
XSqaEBOJTxQuwD5w3wUImeyaG8IJEPeXIBRyKaN/eNuWRUCTGO+XAoLpsh/7jnJv
O1mZPcNC/7bSnTroUIn8S+4KnaRDSNskD8Dyv/iL0Rpmuk/r2VN2w+baPP3vbd2f
pP7a0ta1WMndpreTVk2MzbJrtHZMJPVwfZW3/0pVNNRUzWcOWA14u4RViDFHNbOE
goJT4fU74OTVUNh69XBbuF4zw+06A8GqSR5J32jOP0jGIKXoOi4g5/31+5PhkxSX
Npn+mzeULshlikf6DDBsZTUCnRE6DHpP5Xqmb35b5MnrtNJmmRsnhsq0E0tsUTdj
Tjxr1F05rGzgliJdofjW9h/ioJW8laFwwVQi9bPwePqB8FiaArl0ic1Hk/kHVGk1
12l6aCpsatmDdCLSa5cuvKT272ZayNLm1dqgLCpIicC8C/VijNlUYLsuITmkU6DX
c/3O1ySNwAkPMYZGm86E3cA8ZBy1LKLxJ7rYKhvwfj7B9cxa4pl2TDP388deiOIj
ULAf7T4zNXh5lm7cUy5xlhBaCY0RYqjeuO107JtqQpueERVKaaAaFbNHlcALkop3
l9hcgABjH12wCefUHDlV06ZiLMKKZ+uZ4cc3yZG2mRFHfYoh72HoCSODaWu79vKv
3Sx4CamIu1LfTB4G8p/rSWy5vXSS1dlPKEMkle+yU382yk5hDyML/iqDcNjK+Goz
cwZ49KPRjIAdivWWMgJ49dgqxqMAbuEcxDAAFp/cekF87OPWL1tkA6WBDxanNEMO
ps8fe1eGwHAyHiksGBoxqWkAqkRsPWyLDgl7020R6tZmPjrZvi9mEjOs6t2OtYEf
P2OXEt5ruDf9PUPg/pGLsHI2pM9AKAh/em3OVpPKJdZQ0ocaWbaskLqKbFBsRM6j
nhCrGJVFCLlV/JINf6NujXHGdurg4gLFmN8w55nPLScyro6/2SMzbL7lqX595BKA
7lNsqv4bU9JmLSKxE0U8cR0gmSFZF8vgV5owbnEzQ9fJdPHoWFx7qPIa0H4DO48C
GfkztzHizuRdoJU5R5ueoSBpOlyL2w0UVt7B6GSnNT3VBR+TCZpxx1fTkArA7syY
4s82sY7wJD/aRjHN2VDJFQAdMqH81LbUhxgiaYVXukopFQXrEv1Dku0FPkcpPnzF
GPdM91Y5TBwG6nZgKWWe5P7epP6p2JQisnTSMhC/YWU/nAdq3xP5PmJjpRc0NNSf
AcF0Y0HbipstbzCtx1I4ABuuE4eWZmODwip8Qsh+OqsOiIywPOaFwEdvJzQrSC0A
UPWueL/I/ivJIHVAoepsCocnwdDvPQbeSZG3S6a89qJjRtU5yC5PrhV4aApK/ayz
ZCZWBN77OKLwVyn5Gipecavl1O3eZMvUYKmkRu7pMJVadSJ+kMUD7SzaRrSU/9gl
oIdPJBV8Y4Zm+AauxpRtLxPMhhtgw/K3RNLRbxT9LXWK0RioBkYQX6iL81SzhKu6
ZOF+/Sqh1/PT5jvWxzo2jUep36NagYuqFSDvcJl+lHqRrbCzWUfHrMH25dH4EhO3
QEWR2SaMm9xO5ZOsyFwZRLCsWxOVzo0/vpmSWCMi+vvaQPHS/Yvs5hy7BHKTFgUt
6qvSPg/63kbSIsQPznn67pv/e6dmXyHebhUqnmdY4VVxqAzKIFy5y4GHQq6xFcPS
CjA4PH6re3Yo1HpmJwp8G0CFWBc1C0d9DiA2XnPJkS708E7E+xyfe8WkOAlf7YIt
DI2KsSz9pX6DTBw5gfUXlmzrg8qG7gNp1jhUUY0aL3buEihsd2JS9hcDg1qh2/6D
E1wkFxwhRmV67gvpTC5fSZsgVYGcYfKUofyLTU1MxIWykRoY59if1+sIGMZZQlPI
4nrM6hjPbqa6UtsIOD6l2WREyQ94DLGP0GLaSEgEXHHNDqxHq1LWtJ4HDu51/iqT
Ynb3vR5RIzyAaKbgWOZ6HmTZ06OC0nD0LV5ezN7LxS5g/mEiQr/RhKmyzug9ra7p
1mrzb3XNWvmeChFMFLp2TlztnMX0EUXaLCHgC9gvRrlmwaQW4Q8QPvm2D3vql7U7
nf9qkiyevBu8vWLCUIF0hBNKTOdNRcqANAIlk4zhMkfKdmkMq/Zb0XJh+7HEqNIi
20P69yKxPBwa7ReKMSLTFBBkn3sb9ggh4YS/ZAkuMuoOrYq8R1/6RZ9ASjdZVq/8
aHaEWBIHYVxFGp6gBY4luOnifUTNnUWUbW7/bQ5hPv2QUzjgCJ6MEYsfWLoKQz2x
nwKYNAQ39d9aj6Fz4sQepxLbcI2FUSYsxlwYRUtlfLsK/GjJCxbcY0jHxzXZdnUb
ALE1vknxu1lDruIUZ8V/c8zzYCSSizB/KMQ2S4KBnmRh27N6MggycW5BRNGskuMp
8/l2T5sX0RalEAep10bXl8PsZW1ZJFZ3Ft7vmJjICvdjOT0isLF58k6JjY4rCELh
BXQN1dSeu/wz3mspMawmk0gLuX09CfARiyImngVZ6DA7h1JVaUCORMMXhjqsSwTk
yCY2SaYZqXdTKAgdvYpvWwHMXStDDivB4+vXWOGSYeTw4Z/EfuwUGb2JNqbrd2I+
Y/h8MM+8veCb0WHnavrKL19Egd9Sna1JgZpPC3HJJbY1fvW+68TZH/0lekdUVAQb
43NVbBBFdy0b94E2Aw3TNgc16pMskHoselw3CP0RYJTvjqgJZgKFU8xpSeUf9EiS
UUCACOAgVGEa9N+M0xmsNcMYoRK1fvZSWmAUEogxxikAe3bEdnD9aFumPXzOlgIc
JH4iUuQGBMdXvM+QmVia/cUVfW+qrZUJ4rPBbaa5gMKo6cSEhCaX1En2CHyG0/x3
IlGbU+6LZygHd4jXEDm18hEhQq+Yk0LTf5vbNvrb48YA9BGpJ0asAwtCN9tDi2AD
BtlZ86T2nysEpxgRLM5N2lsWzrHMk9a+YiAhJm0KzVzFu4rfK3Z1iWP9agWP2jOK
L6n0DvOgBm/JqHJ5rEeHVvEUn4SXvEsEv8RegyUo4LSEWyLn6eZKPLb6tqNIWvSr
/617+Z3d0imfdnNmYtVyNlGKHmrvfceMpt8v/HjVAvm0n8hOKmqXJDpPxyAua2Lf
ivjd3DrOvyK0Ot9+uWhqBAtBqsvDeqns4FozKAs6HMZ5A6VvhvtYlL7cRwaBPRbw
gAlyc89RCrqpt3i0XtVsZjcS6xQzhLR/akl0fs4xhkW6bGiEQB3f598XBHUoUsK6
AxphvtGMYK30j1uui1nBKrZU7ZVP6a6NAchoJifymtzyFdTK4nFQfAGudShLliUC
hjI95nGj+k+ek6NYY+wlBkyh2gOIx7uM+yD/fPGgvAXfdQS5bGmJOW6xMtJnNyQ4
LJqs8cLjyuNWtPLRY7DZqeOGPbYc9gldYJT6GyeXpVAVJsSTRqdhuQj9IpIV5UEw
e+AF7+bgjRM78WMLKQ6603kVvb/7c9SJOJj5gy2g5ytUsY9lL2V9619K7hjnGuco
O86Fb3teRncS3JSWDdzqPiNWMwBk3N93+c2vTlscSlsGuJB0afMSmogGOJ9GuBBo
9Ov1Ur3MqIydoHCgZaThQqUSY37+nYQIMGc/8zMMvvdbBVtuNdXP/9nIKz1HA/+8
pzgBG6nropfSG9tz5VFQlUaAJtnWb4K1kE2Hqu/eKtmqLj90WFKIXvYb1A+PB1k5
hr+wBMceD1VObT5o9QA5X3EPYYpLZU8RbTidfbpFIB1uLI6nFCGGiG1zVbax9HOR
meO3oSJUjC59aT2WJ/PJxfkdLRfiHn0ywIYPFH2tbqKpXK68vWbA4sWkbbE/oGLP
wcEX13QLxUsaVnVeBBACbOO2XqUCYDT7BCKBqyOEhMJnuCBlAhB8qjkQQeAhcaRP
PDEK6dmZf1kmjzxK7bFimLaajbGLJa5EVP6GPOoGCo4dx/3IbsArd9CkKoSLdkjQ
KZh5cTrFWtf6Kz0N27spQuVNttrZaOJhfQv9QHDceOxpAYeu7igvvUMKvCEf7CnX
WLZ8IMsaoZiwoG+CVneboy5DER4G1MG423n8hh2tJTfwJMDHiWV8egN/VSAN2gft
A91dsHqJvXhh0REvlKM7oUoSKyfmhGeHmG/QxLqik6FPwZTxxCl30x7N+ZpxzN7A
OAvVI2mpSjHwDXIQfEgECuPhdDA59Qfsy2pwHjS8mLQLA4nQnQU3lYefy66ERiAS
whzoTFVhpoE4gegp0ZSgzQuoShgdXDXlces1RxzWbOyOly0J7TjKc001TddvxRyG
YGErQ05Ke/bkImmqDU/ss+oIL80nbsKytIRp8w66gI1HN1Sp9cPMm1Udmi0Tz1fa
x+P/CLH611ibnhyE0bIYbzfwyWMPpotZR6dT3hP9q3QQd5nxZ4xjx8bOadigbWGc
TZV0LDn66HIQHgW+wi9GfYUxwH1YYOtU3IL8cpDH5FUbiPlgfeyQaL44TwVurWo1
+mTFUbSua5uBhwUEfHmdYTV6sNeu00Gs/44DLmToAEQ03oerwLWpCBu/xCf3exVD
Mp5wIYAJKENNVtzku+aFQ+SMJ4hZpnsl68/eZT9ezqDNoU4cXEiQuF9uJcCl2rEc
MW7Fa11Pmbbp/2hHbCglMTqb0A0ilhlzCDDTw3yCvS1AOadcg6rppuFH7jNur9MM
cxKSGLXNTGfLGKbGTScewjfkVGILj2HkkcMMtUgkKvlcHELUBi28h0RlByse1ScS
Diqbox1yrmzeyFJWGg2f2WXXkz8AcFRIRlsUpiufjjkMgmP4qgirAv+OqdIeow41
duedgIwRnzc4/xtMEsPaGpz9m8b1bnFrXnklsKukZ0Z6eFXTnfYIZQESKAZE/viw
g1pL7VS8LyxSIqmq3RVm2LCbpOO7FrtMfiiq4LM/n+ctJbYCK2frlYR37pdBkMWd
4e3k9duQmoGZGgTjo7hsu23gGlXR0dQzSrjyMjdbjP0vqDzSgLnwkQluA/hGMzaN
CK1qvmh6Iz45YvJAZ6dqUzZpt9mr4R8U/eRtlKPLVePyWGaSXwKEKo66803MdIEf
XJZCRBN+dMhTRzzf8K+MfaiZhBCjnAV9k9zAoxjjoriWtAWMitZA7xksMO1N6dLy
S4xHADgxh5qGhrAHBnx2bWx9F6XC0AcKczKfNs3y5N8g8S0lka7ThYtXOk0Se8rM
aQJ6z/6soOt07D/qgACWFYDsvVZvO2D6+sO//EbRjJa296kLCw5pKbs8/6FgwREw
WkKKRYv+4Ce9rZ9VW+hf198msO4lkEIVOFzLQuzm09EOgzttu5oD8iRrl6oALZm6
Ija+kQuZlKjfIcvprPimzy8d1GonoHzWepWlNUp+FugbvBEBBstCyiz3RnKOMOXy
H905Tajx2Ye3XZU79kMaZ1urUrLI56eWbczh21rMP1+N6p6tKG6UhTkMY61nZ3n+
QLDMcP7Q6JBMZHBSTvVTXOdpQtp5IBoypf1ZK3G7D83oXG1LSCAbZs0R7Kzf8t0D
KO5wjNv4s8Wt8yYsAVcze8JiJ0Au1jgfkKVN38Bb7j8S4d09J7N6Sw95AU1T26+0
Gosygvp4jCXBiapYTxIQYowUc0NQfhxPyS0mFZnnvkydK2KlKMnHCqguCcxHXwTe
2FbiesKtWEtFsZRg32QbimV5X+4jpEmyH6oRO4N/ducdKxJXfvWBw3H5qaRIBasF
Pc+Gbfpm1a6HQI0xyxpbdW/lVARaIwat0avLkhDQMeeQ7uM4/l/Uthb4X3vZNv0p
N8hopX72Lg9DEM5uENJHRjRkwKF4xMdS6Mf7gwO6vftM3Er7NXbACPOh2mtmJn7c
fb975TzmtymE+XbZLPPbrA3GkjYas+OAn+g5GOTcQ+pE4lkNq1J5s7AApN7LuMwi
nrKRXyH8fJoI+VJvdZqC8cSUEC/x+sKzaaeLKmHOQUSFZg5ABQeylGftlN1U5OxK
LOXpw/6Lb/SkPifdJ3tij2LdUn+1D8Hy3KbPeqk6nmfmPVls/EJP7w7ZsA57U4B4
9TG8NpPUXlwsP1rv39Rwkf7VaPX8W2qWmXazRq2Ygk4hLTjY8J/3IB+sNzg16R4n
QEYjYiHebsIxLqkPy97mkGdBHLLfi51fRs4Dhe0ml+smjl4z9PMnlv+6vt8TdldH
RggB8Sb+IlOwni/oL0iqtxKuh5eMPZa+w3mztGGR8o6d/OmjaM/bdeWziVtVH1it
SKYDQP5e6hUcHqA1QKRiz79cOVqr+RBEExVzh4bFiEF1+6GZDzia/l+nLmfpPXYf
omZ633tbFwiGOzwInT1PTtSNf9hXtCAHN066OG2f2JnOxnwSCBccKbq13r2Kizvt
X1qaVbNTiAOLWOmVXoCcozkNRAHVnuel9W5FQXCvHObQXK8HSgSwXqMU27R/+OWv
QbLLISTValYeklr9d7AkF2+37Jx6adFSRuYqZ1QzNhwEVj7EbfI4xx+U+Dvns83a
1QA3+l0yKzi32/DDWfia7I/WOuQf8l2lg4lfJ1hTD+Vn5yAM7KjxQIblK3nGxm4W
bK7xwUkEH44g7IdwFDRYAMGkAeXKpjIxOvNAQxNuN4ju1RZXcDzu5XYh1cjpIEEu
Dw7+AxIjQYNZvjuv7fOO6ekTTMo7e4TwlBRxoWLH2B5TXL0NV1Ux/OcYuXh0y+S7
6kxtmdqIETxkFj176KlPQoLIBR2OnwL1c68xTVpTiLVeglfDNXSrmI6wg6qcylIr
876g1SJfQP/0l5KNH42tGE0lIRoqAAZxiGKQ3FANXz8MERbSNCV5Phzi+2dBelQg
To1jVTe0rYv6mX4BvkbUarW1xcvG0DHeqM95YH5wJpolnYOtshPNB70RFPOxk8/5
NCG2f7+rWlHdbutduF6KkgJwd0tnBbLQyfhQjtZFR9pQTrD885lMdBhRATKmb6g4
b90JNBhu7Vy0gK446SCI2hSD+slHJeAZZfxercam4tBZQ1vLGxkKKaIHRXD8T34X
CXFjsCvUxXGAsr5482nDie8CPHQTIsuwnT966JXCP3K2ooF+lWo4d9HAm8KAyCeu
Ql+hrzhe2eG08yCWFXllI39zSekQvsafAoordB7zPKjR9bnFxd2YgiGgoJIAbVuD
w7g51gAabtfsBRhKIYD5Xgo02IrmW2KwPKe1fRyKmEO/H9hI+C109MQeWg4NnGAj
v7iw9uhqddkCzhCwBZlTz/xd9nJnXCdWIAhBqR9JWEHoxzTYcvTpM+AlV6dW713/
jHlMNA8XD+Ge8LiIFE66vh88CJe21OTqUGla0LhbPGqpsMpFovXW20cpoNlOq/vI
eb4Rul39NhGltlM/Ecxc/D8c01bcGyZ02Z/s4T2EJoPL9U+8aLxYo3D8A4LJ8p/B
bR1FnjChZJ8yPENK//kF8bFwGKZF0bXnR699kwtC3iTFtFS4QxJnhuPBz+cCxVaz
FoNIfXjDmbF3D988zHjZQZQE5p6LJjAcJMGOqY9mSX2Il1iSEM/1WTN8yp4+dxh6
0q9zZrfHReVscyFvHzxB/v+TjFeRGzJbRe4dpjMU09EGTvFsU/8QFQcu2G4PMs51
e0/B8M6yvXTrFPLtPfUuO4LC2O6pXVS3JWm9Wz/xPHrnUrM7c5MN9RVg4tOXZdr5
q3Z018R0pOnDzR5pMnhdirRYzf6WldvwqTEIwCVVq5REms88aj70u4wAcfewjOzM
AuMrRjgFkeBH+j11/TzL1EmI9tW7SlVNHnH8KxSYroY3qsQeBgYhThjhanKCerDX
R9v9izlqsp1Deg6621KdbpEoPHsNLeqPwH8aCom0xDzmRH3bNT3eNhbRjEzJFFpv
7RR/wNRdWnls3KuSQNM1QxzI4OPsPUIkY0XhEQt/cVvfuSqUeHxsNhty1oJhu9Ow
cS/VALT1/1gdffvW6n7nH00SgH3YvNUrZvMt3g9gQ0ay0tflpUpSCcbUEeWGjCAO
EBu7dgqJE9d6/cQnJshHsEiD6YI8iWYndk9z/OTMlbPj5GwP/JLPvifa8oj+GIMm
rpTyoyxGl5WWpsA5fIC4pogNtn+z5BG97zhPOduyooyl0TcO/bIBikkAxc4Wl9FD
qTzrmX3l8GHuUeDY/NCgEid77vX979EzLS83cJKZapXvh30qyGsgBaoSo9CHUTbK
HatHal14BYPgxV2Nh+oP3UA/PMoDST2rXfPvaCiPH9cZCbmdWUGWusMLmiQBxvQP
pUObVnAJjwp1oVQC/T93ljhUpoRRi8dkrr/R2vb/67FVIwE4xaFBX4ulM5RPRYKu
q9K4iSly10pcKP1BN5mOySmlKTgC/8Xb9joYGxTYcODXCknDmYIFKJdASvaddSMA
UFI5SVWAHssC14KVdrpjLwPu+IylkQNSrmdoqu4LW61hSUnKR0UoXWcUtETHRElf
pd9vwPDZAkaaFg/UU1ssNpx8qCzmmMlPlUYWTSXuHNo3B19Y/vBijmjKgmTzl0HN
qGb7IcBTMWSBvpdreWuQpndw+q5coYiwr7peewRgh4g+5Wbzz6XD1zgBecjD3n7V
jLK6mzwfmR6hGZsBr1wT+IWS0gKuRnLrQD2m7thk9Me2XuIA/sh1hJLjIV3n1wa9
cGJmM9OOJPZQyneokL7h7MCVnoeyhGWIq+xM4T7VQPuX9nQSMUeMNrOJyC4aoYlB
HzZwm/8GMY7vpMORzaoGfUtZ83OaWh7wnIUcSYDP0O1Nz80YCJv7On5hug/zBmKJ
KTCYl+bX+cPyIOBs8nBHYBOyFDBQIprIvnmeB2ZjyFajvnYu1+H/sZpeg//oTI0u
YWuDwngrG4StwuS8Ickk/+pPYGFw82f3O19AqHIfUAkUJOPQ8qdSkXi19elOTDF8
Gpq9aOItChf4Y1W17cDOoHPeYtDE1Qiena20XehSceFygdtr89ccvfQu7pKJ7U0A
FR6Awyhr33JhJvssyim5K6KYyd1G+r5bfcBeJWq1dmurs9bozX6wi0iMX3pRgJiR
WpmJ6noXxSFnwAHCRLQXPziwEcEO3ud7HjRhgL3V5o9P6Gt1XscT/IfX9cgP7Kjl
u5o24jvjtHktiseux3649uApwfqWXoJUnHXEK8Tx6TkhYL5l5TAbc0uMvkD/6sB6
5WZXyF2xFc8KhCfnA7kyNxVnT84DQC8Qlwh8XBhz6VTcJohshw/1SBzlKcZjSOe1
gn5d2MJNvbInt0SSnzdtNdHdLb2UXHzGDmMjMZ/3n4Fgz2k9OHXRhx4mfHdU8C7f
gs2skaTT6tEfNMxtj/w65q/89s7iQBEXf+kQ6Bf95LreJ+/1EFI3jHHXJSyJ0mAo
s9CJ19FYJjRlpBOhOYd/tRNG/6HQPpJ6AMgFnf176pGz0kl/4k79Hv+o6yjvopoZ
Yihfy0tQL/A3qYlKMS8xXP0WAqA33clqtyRYH/5ZW1jbBBhpnCg8EtIk9cEhDujl
nyZP4875rSUXGfb/MPyuDa5B18D9+KexHdIk8DyN/4rW+fuNf3vUxAesM7o73s/m
P1QD0W/KOzY8gPBEIT2PFrD6OIBRsoBsmAhlO0Q4Viho+H4lmLkK3X9Lg+5TfyKx
9BtZHzVyUzdP2ueRGJ8QFjims9M0gHvu2cvNN3AYrlz3Tbf4b/MXqme5Gxx5BF/M
OF/fKezagAmZD8K867h1GsXzHF9MlrzyZmbaHzVE6jzaTloPCJbaIgAcskIY9fQW
O74M6ZNdrfJ5xP9bzci+QkP5l/wJ/QhYJ2AX6fqMnQsJp6kwkMVUHW8IPksiL08y
CcMXVxHbp+H31DdpJ9uU1U1IREOkAOsPefuAXsSAZ0HT/3POdv4SN4UTGJCnLKx1
1kFJzXAcmWuOWqQ6mmfjUgzdAnwAnZyZBPLF+LIGy9R2ZiSXgxjltxLsJ0+H01wo
aaK1mxUPmboC4lDy6WtZ7tIocQXPRADphB5P65opALKpq3jyttKnvcNRFeKPtKxC
6jqqnXA3gqA7WxFwVzRCFtTB8RYRdaartgodBHALNo2OR5Ts/gNR0bqStXH2oB42
8WazSxU8oCWUxzWN6jHcb+Hu3s3Q2OooAqkYefrLjnYWIWvbCekkawAQBkoVfgqQ
3TmOhpM3h4LM/Zr/tz/3HjCRWm33ynv4NkWOGoT/hYG/wnXmCrlHCyYwiZpY55M0
NTwR6NnAKpnMrhE+d5CZZvjk3K/5r31LxMWSJm6GAuVSMANGAQ0j7/akLGaPMBmG
0Yk67vkzFju0sq5D5n69LKVt3T6Yi/bV2IVyl77bz5hW3l9kDyCz1P/p2DTpKrOb
pU11oErx9ma/kkRR+xp9aSm6LwVafw26l/ULjzhKsKNvQj+4Z9kPGV2e1CdIsC3J
P5KGsbudw5YmOzXpGanh9PurzDMw5lvP8iTGe8lcv3E/7j+Ty7ndQ9xBXS1dw0yD
sIXaVD8L3BmhEf7zv4VJ2ZTvY68TtJJmn/zYj14+Cs6ckkNT67wNuh3Rgi69RQcT
95VXkz4r9cvXueR5rwCtWisqdNkaFamleiLphJbr9sfI2I/bttleCk5Hx8/M3jmz
RlRjmtd1Y7L8VwNY845W7WWxMKh8LAve+7BuA6tZvoJ9zHQ6PPPqwF+Rgd5BcmR1
B891ovhhNmr9qYdRni6Vh2vkBsbKypm4ssO353i6uQwSm4Iyh9TGGGGaalIQ4THc
KvxJ4CTiU31UoIIYQvZTQjMTYcUEpcYzEKKT2BOVPh4mzA4UIbgehGAJy4b0algn
8C5I0cL3cb/ifYGSzLmqaqBilDL/wNcIrNikYug8yQYHzL3FGBJSU98tLwC24cNw
nPWiBiAtkmb488nV2kFjyOTgyEigHE5eOvpRCnmFvAiTFg07HN1D3mQxQq+MSFy8
XRrOEVaMp7rvurK0bUQKc02C9lVqTGjJNgzuVqOhLb89tCqX2Uh+3oRbVEYPsfWQ
UYlmtlc0NAefr4qKTCaoqyaLE9tUN0ZfFbEH+q4zxeQJDSXzT3ImdX9G7PU3AScN
NjdD+hEmIcde/Il4SsrzmImFawXwDEb7yxPD21fUypBvzIUhhOsYKw5hBUVWCo22
plOLbDyrE3GYPUY+0qFbXPbVgeLufIm9lGRZVp73WDDFWxM90kLk1iyOZ3q31NQ5
KCESM0zf13S9qATXFMZEWpTZuiAE4wRO2AUnzaIIR91iiIGumtPc4yNeSLkq4WhO
>>>>>>> main
`protect end_protected