`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 20704 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
TDkIdcJUWDKCGvmrQYRemGd9HBdDWURfz87+Ro1TgtsikWG3zrH3kN/gYSp2yIOt
JJ9NG7VWdk1VXj01DRkQT0ZxGFWRPjmTOCc7HoKUVge9/E/XouzQHet+cWBm36uG
4DVGLxW+XXRfLrecKtQs7iBHydDF/oo607KfbeZ7pBHOTS8lNNqh1rzwheO3jTDo
PmcgSEqnFnuoUfike74siOS18kC2bk6frMcNHDuDV5bqcQY6vgjVy/weus7EzNL6
PPYxXHYwAZyQUU3dSsV3loRnCnLMkCV2blr/YsS5N4hLftW+7wB2nJXNxjOey/4i
qKMPtM5MXlu79EMnrRY1S6LOnaxoyOFK187ArNpv4EHiTh0OBkvlb6IPio12IiPw
bbqIZ4i3LbiwBmfSHgOTfGcnyj/be7FFv3SBeQMx3q5XNBSV64S+KqyW+jbNkCoE
Kto7knVeqZHTrIS/0BgRvSdzcywtUcPLLxxrfXlxR3eD7MM1qY2/1XeFjJvHKUCQ
SfB5vwR46gNBIfzUN00UlKbAqiB8il3b9pcfQqpau8WavtCKiyII00XiZB6tBW/q
K/0TCQoprMGs188M+xwFE9M1SGxF+tK4CH5uDLmNgT/0nNl+ffs9ej1sn6P3hy26
qZHgcmEGfmFFmsR+YzCBjrJhPhyDswi2BIJHwVtq1admT4PANa1IaifQI3P/P8ab
ndsdj8VUHwDLPGzi9LvgKyYHfWZcxg/DvWwhYMA0/Qf0Oo2XxHRmZCmW03c2AmYH
wWEEAU6i9qpPP0ivgQu7pX6UBvYkSPRCUs959AOpOO3yvppn6+SePadaXg7NRgd/
MiSHfG7xVVJA/7AqhD/53C1Dr+r8q7JfIVIJI2UWXtuOfFKknN18NR/J47D5XEWN
o4QLG21gj992jaoWufmcQvgwG/1iYd8XPxniIqtjk7XcIryQEHgc0J/wU7GLLtv/
4fv66iVyR6j0cue13nbg3/cxh8PJx8DxsjrVYpNI4IbHW4vanc9EY6Bsj5Mjyhd5
eqQ0+j9kzEH0KHXrsMqGO5g2qx4+n2w4g/k05X3okDmdDKTYvftRR57ifyC7EvRS
v3kuBSNR21jU8jcT4QWast+czCa41oUty7i5aMgFI1CUOaYusrsaw9Z239G7M2rU
f9o5JeDUTeqH35zvblEDhHncEP8qpcEuWyrXoQ9tWilVsHLtJyRggayVAQcLkLaL
0KuiXG10a0rtEAOiFmSzqbcSLkdNaSC1enHEu71ow6qdu0AEw690GAJYrja6Upu0
GrnhMKK9syi9IKWdpoRckT/ERA9eAAY4AuSepCBSdkcguJIPQvekMA8c3mHOuGY6
9crPvGmzlqf3In0109PzWFO1obbZCKJLM3JJ0aS++F4Mz0kmw0CFiMINDItG1Qg7
j6btPPdTX/qdxYstU1lHowXAiIejoiRGT6UjEOe8y/DqmNNET+q65lHP2bPx4oBy
HJ6m210dx8cQFypSr1YKmCGmfhAwRqisAVIboJTySXjvQAErk83k9Pm5+fS+nf8+
OI58qwM9OGfAm4I7Ylh3Yky0NtRNSUuzesHWVP/zIap3xqhh8SpZxgqO1WKU9/Xm
G5hVOdgzRLnmZ9W5vZnWTQ+vnZcpGHvvXLkTjQtkU2aVpFQm3FY/+JqUXPQ3avFJ
rZfmtlJqXMSc0XYQzBuywOeU9bfd71ulsxtbKBQg5XdObr6RpOd741Q1b89czjeM
5RetqHz9pUT3gqY9STyPqI9wvMD+ADDddKS64NzSNbQrC6yO7Zt0E2h25IhH7NUD
Pk+JX0ShvlawPibI7TLLzf8/HpnAQpvoT4SuzwVvJf87ZDuaYiMWLTAZMxodOk+u
4Vn5srD9nbWP+r1V8vFSIaDfO8CEwQGHDPV/39ltmnKJlE4l0DP3DPnlDwYNdTGQ
3qHrQPSLew+JmZQInV51JxLXsXwCsIzLt/tRE6TRACbPJWKMmEoefT0pO6mfm4as
ucWdJfpy+HjWCnPacDsYQoLIYtVadT8wCJPwNNOwkgaHIhwu15HnKRr4u3eAO3G7
ocNeIh1yY4G/SL+KJa/Gms40Xneg67AfSYfSlFsXsBQqko+ATahgdYZuVRyc8Yrf
nMn923ET3m3x0nNRdv/a+pr7gS4+FOhaF2Maz2ri+LxGbRrl8MqH6GqtF+EKi7M1
YKBwsE8JAdee9hRS7yrt/4rjEX9/6Q9lEtfe3LBxbV2/DOLT+CGvav2vt6mG6tW2
a9n9QkZBAq3U91LydFiDq2DfNBtyLpMNa8VHCaWifT7sUNdffgEeLZdCBM5NNhUt
5t2AP6YkMjo8n0o4mpTgWYMyTUUshOMeSRkTVMLF6Dp5i9Nx4yVyJwiG/uxUCTZ4
tQ54FITvbH5dyUyXHcjHeMmC5M4HH+gQTYz633HLX/HP5g4pS50UUKklnlg6B4v+
JfDOKsNvHkkFZYP5s+FQBwkBSwW7HgPSw0GyPz2WAmNfyXeJtwgVVbDIOSNd8SZl
j5GlESnLJqOM+nFzKd9VI2x+o4J55m7pimNRI64ZFvaScWRv/S4gpl953h623Do9
5BpnrSWVt3MWzo/DrwVR8RfQcxrbLOeX4JbPnRtnXPYRrtpcG1aI/mwKs4swWH0W
RAkrJnNMwS9vJmKcOrFjSOxeNM9sZS4VDoU84MybzdmO1QVE+ziWIDB/xxZkPAN9
5cyf7HmUtknhMs3RG1Sr6skmmIBESirUl4ePX9f1H25dtaDf71D2gs1Z6Qfj2/QC
HK0qbZhwXzkKXG1VxMBl9CHlR+2eLdoY3z2mRWpRbFgqvQs/gALC5gOz+/DsWV4z
fBJm5Ix7XHbcMbCitC3XuAUsfvge7y/qyBnXAjJK0c+10ktTQLdHu3NMHmlmlZm6
kcTw8GV7VbpzHrcbZt7REXAJWXiZfcybngymhuPp6N1qnMu4czU8OYAwYNYM/NHe
noZO7sdRrU4xfI2z8HDKpcR47VBVoH9cyMyfNu1z7gKbYRhWDJMcrNEt0AR7rMwr
BBIF966/mVIll/8jy6PAbejs9PGeiUKuQaQK69aLEq7zpvxfTy3km+29q3b2PVKR
EEVfjcbYyWuX6F/iQQYJhjIjvq8jlztb/KNnossu26RnVuJLCK/OLK//B+KB09iC
3RtRwGWIFJpRPC1+HsH9k6QrrDQBuOT6Hvk1t8Ysk+QzMvrmqLQgvTDmMK7v8YJ7
HY8jjOCiXSr4ZlPZcU0xDlp3xbvvBlOKAW/A6+fur79EArYZ+YZVuY3kxes9MRia
f5lQM0l4Nud9E3j764LZtcZZFvJ5bf1w/HltlXNXgPCxzbtPKrnEyQtct50AbEX6
6lIXjJO6jUcThy6h69Bn3SFTW9Oy7oK7H1PyK3PtmWGqpIpCemrfs0eWpe4y8ykb
5XKcKWsgizSa4pfhPREch8YlnbYYvO8jD0P3ZZBxj7pQcYNNzmLy4Ymh82a7vgOw
q1IxnKrJ0zAXDj7WTKoLQBbDuf9RYKGg5aqaqnBpXqSCyQ0kCXX3gJ4zdD36Q2Hd
Kv2ode+g5uhUtIlEI6n3ZbjDuST2O5t6+iDB1XyPG5n+r/nD8MTbazPpgSgpP+CM
SSC2bKcflL3e3uChHg3dtbKBvMXrGB8HUxOlAAQyJ20C7CBT8mMX9pMdkJjQLoqq
lQe/xqQ/4GvzNI8dMwQ9686/Ccbeg7mFzsi9qy0La4kU41XGC9PkcSTvE2Bysl4Z
FRhXlb81ABSMHZ5xV2Aq3SlXMERhdLmKySsGIbYj+u2C9IJBbt3hG1rA4pvWRxSu
aO9jTXPo0qemEQnjgCKFmZIBJKLwiREDrmULFBPhrUY/A4PMcgqaO3Xh4hxJ338F
wMCcvJ+CbMd15x01+EzPB6DDil2L7euxKVMhRQ6Sdovu/Z0gLQudSMUbr82tJvzK
5cO4SD9EY1jIEytp9HaPlLAMKLREf2HvY5QBlyZi3MY+UnktNAKZ64+3lbTa3pbD
akWWNNcCuySuBgO9/2XNYYA5A6FHVGbM4ijZEtaiNiPUAZlomJ2vQCVMqzhqpIty
QB5iNrTJMnQYzFvLXD7xGv7rHIAlZti3EZdJYnMykvhW/9odOQxk92nrTqOee83l
gPOwP7MMXezBZw/uDCxiCfgp8zZBIUBDTvroE1TrBWSODrPjNP6JmBmXydKHbMvO
cwaSXNa80zW03kRWls+ybD2W4EnrVDimCms6LMSSGf91dlPyEWYlOutE1mH+lmDF
n8z7sS4L98UQhgSOv7CWNoXIhOzI02UbyzIooZgpeIu57g3WrcoVZkmQKcSoNiv6
DduorLkFUNrNGq4X6vM1la4b5FU10WrJDaBMYhj04El9NFJmbFXoajPKuniOnINb
oDgIWiiQV2nz9XM76QnsHuYztj42vDDKsxC4hFHwIdjXik8JejlaC70SRrQlJxvq
P1DnE18HcLhCPpoywbEzA/nH18n4SB+z0TvrTdTI+knjEYKoh92EXcoxCYd9m9Dq
AzTFVMlyu69k3e/vL4GNhLYbv7j231HIX1mc8zAxdIHQyb2Ezk8ZCOXSUIWNfTT9
4zVXCs8SgMK5UJNRXOKWFnW8oCqcdtyHRGqqcevYstKtUGMvFNedWXMq1AQDvdy5
rghv5Fj6zHG03Pb/BcAxxn430hZra2+QjFRhNhc6h0aIVZr5K8RE+Mm3vmU1OFeU
rDexasipN7vsugJoITXfKQKDdk3wcwRS208fbcteZQQxUhYcn58tM4oQ+0hi1HzS
8J6GTaUbLytI3tMO7NC7R+jgjLNBwXM5H6u3IX0vrBACRgUiujhrkINLVyQDGdKI
WMLLa5GL6P4+ZNGE0Qc0comCzJqyqjhYLJI/CWR8C0U0aRn0SysFvoT/mKhLhfrR
MOI0tVicwnXXJ3vsS6PbKzwrgzhpVZ0v6oltrZb1CdcffrvwgcxVOsIYRP4IoW30
zLgxtf84yMsLGrX10cP9ouvDN62uZ1spkE8GjH+b1bSER5CLTu36fT5gFGZa43pH
AQKRXMm/6bejPCT7U4iU4hBM6r/E03J8PMIVhGWwM7WG2jF4blMt0UuXfW8Ct5a6
Qgv26q4SzZhukp4SlPD9c9d8lwdUa7u8iZ7QqRBUssuAPzR3jkgEMVgOExveYNGd
bmDcozEI59U0aMIfBc8/2FrFerMu9CQ5Vfy50ZXO/VFSjN3IuvvvatxsSzzBgXJg
48wSOFFfWzvpCfZRlykc3wO28jKahKh5z6veMKm1EfowlRf2cYQh5m8b0mL2anYh
wLWZl33lADVWub6Fl8UbhKjuekEN2yrn/9rNZ+PrFKPM+J2wrGgUSyBjtZhpnFNH
yFfAxeasdfnSN4YshZnaYtiSQerNYlY2TiDobyF89p0HtUD9BvdpEQZ+YtWElIRv
drKbPCwQZBZ3R/kM15jdpEup9tenal+eZFvInRlAgmQPLS9lYkSddJvlMWUEkrlc
kUpUhUKBXJSGGbCVqthrkK/VOFagd7kBcDqbR3YdcnzVu1A3JFZCMUyEWQ1qFqrG
Kuz6UXvjX8RE+hpI7WevFjKUCesQ8cvLRQeoY8k97w6UH9lQZF2m7yjEZwD1rYKD
LmvjK8Jbn4lldASryLJ8kCxargWLqoDTUEx9S2O55LXGtoOGpmNY9wsqW00pCh/E
SA5V52YU/EiQ45XbHq1p5O8yXmKZXMJw7Ij9u4cvGaSO2ze+16lffwiiiy3ME2Zm
1oUN1gD3uS72/RwdauSQEduLPg26INlxDYkNeFNSOGvxBpFA08CgCDs8x2bjpNFU
TlIAMAONpQy/nRECqEdgNC2PItdgi8esB9GIs9DA7NiTBSKZWK2tzKXISVJRrWxU
Nh8vhEHA71NzMzthg63vLsVeHUr5jgZ8pjX20xmN6NVGIQm7peeYbV44rBAktf34
6mJKf9vT4VN+MWGeOqKak6zCUE8Ru6+dS906bqxeXzrLSN00bTvFCF80ySqDELqk
HoQ8dtJBy5RGyEnSLD6pFtAmeSaOkCKk65NHi6FFYu8lYnm1IMTMBRHoQtWnpssc
c6AhQy95g0Ym5lvL+vzOu//5xrrf2x9kTns0Szr9arxGFo4PrULBJo/Dkzo9+zrU
cHyfTItc6t5tDUv3aREhPjpcakOm0YRU9cl1EHMF4875yjdwtwskvAZTSHFoISra
b/6Rm+yHm0rZ5HK9tFyQJOTjyxCrTdqxgt/6iVRY1HnpNcBVqihbRVP46cqrHh4X
rc74Ex7bAUvX/BqKcZi/4EaB8q9SYLPngldHrlHef452ImK9zUhUDzb6w2aYv+aw
G+O/fcSsaWHJpvQpDp2MvDxR5D856uY7zF4beq8H3Dt0xvXZ0HX+yzt1iCtAgRQY
RBHLW4LjoUOwU7wGuvRaAcakexbN0I6d0cvMzs/iPWLiMNsh9FHkQVvrpkg1dNz6
/CLAmB0r8vZppSbGw/dQeVeUP7o7wMTQaitzcJmdK/g5/xOL/cTDMSlfxVpmEpCl
XT1tWptiPC9SkjQ4I/r9WiCiLaiLA/PsTN9mXKIBx4jtFC5OX/J47qGdPUI8U+pM
Lq3AORxDo2bur+9OSU9Kyohv52Hz9tzvF8BOomGEbXug40xlH0cbDURpgDe8eN0Q
dW7Gkn9XkrPS40W1fl04eXQX7D2dWOqOyMjJJkspSCmcecw51dE2+b4ciSSWt+rr
5cw+qGS5hLDDp0CU7FYfyc32JQjuO/mJpqAu5erA/5vIRx34VgQK9dqzvQoQQLpP
q/KpHDLkLQEF/Eu5t/lyI6erCrTdkVDfjVBPrjUM39KhL5y6fb2g7IPH+/Ntn0dC
2PIjbnOGnZ9tzZCxNKFEJA4VM5f4TbLDVxRqntDnEKHBOaAKumlZda6YREgf43y4
2GfyV9CUl9inr5lkGzwj5AQ9HnW28E1uKhbc+4Wvarfk91kCrxSVKpXVzBUhlFXp
eCyVAXAYL8nzRNmk3v3KHhlZmibj/Y7iUYCuBckaUow5PXmR929ssydMrTzbU3k/
4Bs/X790p+LPMJ2aiOiKF4wk9NPp2ZCGHW6InNE1mxXH8O7pCj4d62kFGkpe4kHv
H+ldWt9MHxwEnyr60qImEqFcwkZmcezGNvJREGQMtS5hj3oUOzfH2xtZNLlMGQFi
fw1g7iCsOXeSoS8R/9TWW+drdL9UPmtXRYpjOeltYygfaAiiSFhGNO8C1MOggMzm
l10ZBhW6U0Ecr9PLifCtDiKhmqUSvId3i33WhcGaaD1LAPTubLWBEt57fxv/oHSM
23LdUDXmUj2yD0Ke8a0rF4ijHKJYr3lF9bWdR2dcCtJArsMwKSMMdsRwQp3lJXz5
5BEfABd2nRdHBbLBbHVPI/7qAR39Dmr6HFSsfFUtcCVNHRv8ROSEb0bFDauFPrYM
jGCKeLyCFORVaubbMBKtZKJHh0ULI9F3adNVoJy2YQYDmY4IdLGa4qKm9zo4Xve4
hL3Neocx/Lzf1opFNvHxAMMiFF47JW4fpNtp19e+sjK/OpWDhN7TmzS7FGIbu+98
SUvta7Wsz1wuHF/MTkYvTIoxohXyKPWRZXFlGE2tVf7pFfUjEcIw2DJc+p5nbEEg
EVWm6SypDWFoCXrsF5ZwBSWfclE2o6+q78fMB4RPC+Vg8SSqLr97vkDKvqeHLmZp
WV+WoUOE/41wdhTGwTTwSsN/y5yFVdBztdJ8PO8g/HULuTI5o5V8evDy6+DQ7UFi
sim4Zz0w/l9jpN+TUhv2mLdktz4CApQ8NrCKx95Ys93NmkMasle0IqsLOqpNcsma
/xqnpmiBrUsCc7Q5fR0MxkjYBCXLe/LM2f0/o0utOEEelfaMObW48jlxXSCOgicO
+nijF3IIXGBUg4Wn+Z46Hn2AnF2cdQNtnbZbdhu0drYF/LG+tDxBXwWA3+FTtCXk
TVfQvjEFMIi5gHiJuUP5e8orgmoLYe8Pbj87+cNaIfN8r3r68hApAsGMJ1fmu1E8
i61XTe/lvtDw/L+tHKFh9WBawCYmn9COdJoZHU3x0CufLEeCV8AZgRpXIPHNCmsU
6qEKJqtpAfkW56g2BTldJA2KTvh+rlPANSRCAxHXgmY3SbyEE7hz5gvFjEJD0hoa
n6YPflVdcHNsLDNmqzme4/lW69ca1nNw36O1glkD1ili0+ac7PJmnRHYZIBAdX2+
rRQyzjtZLOv/q20+UqgAYIjmyXrSW7hMhVBPBGysIjTR49f43SpzZlmhMeA54dES
XnfiWKtkjNRqjtkFv2TkghAV8UDXZeG9JchIEC1CQX3wE0NVC78tdQmYif8K2N6j
puDzeVkNkZkc8esBRZQ6mvq5vW7aaTyIRYZu4/WylcruNnq6avqG9toP2YblmfLz
DOkZH+BoLV/JRxT7mSDx+ifZ3gRcAIiAGbjBv7/dh2XMLFqGx5lXh4gK3XsGndUd
MDKdyTqgsfOGjTXrdNePodkzJajwlKvLKApeMOVYFPkdSOnY7A8OrMb29QsuT4kJ
ZeeUmCmrVcYyt3BWjwSVOONv8IMEogLOL44R8f9FSP48kGGHzuuGbKpeQc2ugJzn
IGxPMtKcDcWScXu/OkCCH8D2p7fxS0jbk/FFL4FqKHggp1yb83H7amL3YlxV+VwD
dqo1u4EI9u7Zjis2G1gkuuVVqVC6GFxt/q9bFwrMPkhkn6vSurnn+opXotGQgdQw
Q7f3m9VeLGW24RJv407FDSv9YWPVVNoEgWNmveg6Dv7aqgFSFDt1BvYIruq8Az7J
aPz26XosHYo2KXNMngSU0HlpcMJ8Kx0Tj/F4XrcuQiah8ETJjjHIDnZwiBhaXXCW
B+Gj3JIj5Fj1HoT7rfNA835P1N4/cbhS+iGkExGtT3bMNpqAEyB4aqpzh1NFrqnT
Xs0YYyhaLKB664skffvI7ldHiWaCKNbg2V8HvpOiNFHb+12X3LuQ+CbzSLIzk4Yu
BOPwB3MrARketdnDEdppus7J6yXYRjaFlNeb/HfAkeVvAMS5uLhRKQQXtSAy0Sha
ss1fuUSczzhxKHZKN5HyIIXv+shW0fzZ1Ta51WtP+cq7EIMk0Diy+h2auKq+9xOc
a31pkdLeaCMq2DMyzHHZG3e2l3mA9FBDkFnGSbmvIrVXH0tAj9kOO29IXLcRZD5h
7mBuCDBeP819RkUyNHrTDfcVq5pwElm+CcfSXyva57NREgp4B2KWc96j4GbeparX
1tDUQnoDTOis5O5TyjwVUYp3uhZGCGVRY0spD2lGoJr/1Kvvzt5AwqIlEE8/l4bV
/uBqgwOACpvIsAHlwWmp6d9KofCTC0HoLQDgxL3i5+xrfAcyFC4Phr0yLxtlwNjW
YU4oXa6UHjK+gDpvJxc33dlTqzmCqUGVazn8h7erl4iWfgHZJfBcrumzTNToUjPV
iIf88G9/woIwxJ3Athjh43pjHwZaVgU07zmuAyzFbbcr2wBPxyq27pHLEd5quuGd
M682a+kDFvuWk8lvapUf2mn83I/McRQQyT17KR1+ZfGDxaWy8YbXIHz+pOiyWErJ
/dOuAzQtJ9dhQVa/t8jWOs+lI8ETqid1EfXWDw0gTutEk+dwInVphTT/3ai8XR66
SaHfALjef7g+i6zLKCnX19ImxgZqTmE3eR/IPRdRlmrnY+eBtWPOUwoRGkmqss/i
mXiNhkRNH1wYfcw951eTz8uqieRq1AxdpmbcvofwEcRZT6eaxzTe8aC1mSKIIlHy
IGaFXppotgDi07kYHxubwMLVjIeCfnqZpgJ3qxO1KDMjnZ+AsTBZyd3lY034stH6
Ei/hFyuHz2+SqFpaMvokSINyvMN5mKw7Xcw6ZV3FK6te28WecmsIBYYAFNdEKaF2
af3968kd52nAA+H07Dadqt4nOWEVtWMpe69Akm1O1EmOR3hMkJbPVpawawuxSgcx
KCANT7SEa5chcNEIAp7cB9KRuJxruo7Yhbi1e1cxUUSlRu5PzmTCROK8mq9C90SQ
RpWftxTcF3632tyqL5XSWjDL9u6tMxHYbKAL1nEC8xbO+tEhFwRxMZdbQQCu4U0N
zS0n3D/PIvPbS9qsKTd8l5688R8kZwJQnNm9AU821CXcO2xuIqYrGueYwEfgTNW8
l5CItRmS3/aBYKYvj4vfkXh9vyab2RUa9xDiFexJVErTAb3q9Gm3hBPR92OVL8p4
ZCNMJwfFWQ482Thn4DMU45Yxhiz7qCz8dLFn0qy4wuta8Z3bUj1srApO9nHrMycy
wL7zY+7bx88gKac222wLcnlw1qjtcbSE692cOC8DBXP8Jtr78aRDCZ8urEL1oOlS
s9R5LSGwO3Ym2lsjV6PQlciV9zZsZf058My3A52x6EefbOqOpKVabaNVgXXypPav
FNlX4u3u3ih5tPdjHAdQ46aV1qkLbQbk+PEQRrNm6rSsyI8Ndz2FQjuxsvXxJGqc
ggKHGpTmc2kEWSTJN/fWmMGPE3rHes11Sk4vx2nWKvz0QiQXqVl6MukKYZGICMzx
LLQVkiH4MDM2QqvyOBsLW0P9PAC35yHJtBLLGXHL6NEQJQv1VkrHK0d+LHppk/+g
Vk9tVDL4F2nLV/cy1HeY3UzemQhtQrvzFWyMdq5mkd0t/Z0KRqiATSHxgwuF4I3n
RuX4VbpokmbSUQ6K6sJqDQc1bXWQCv7HPO0abQ3slf67AKFJccrTUoXDBSmPbf9j
VdD19Eu2wAMxBFVNh+JBksa4nzHehQ6UYQDwb9/TYxT5snX5mPzu7YOzgNz+7NDD
7TQLUpTtng5t+oGseirm7UfPjdgpkhYvYzeVqHSzqxjio89wsupyf/ibBKX3Vv4S
t/ATZ5sdGxn9cdW7jdm4skQX1K5S850hWNn9wZUHJ4SHycE512wHK2iTyKVe78W2
CTtBZd4cHtLSHdNImryZeg2yL6a9zgYTt/LiTFr+esK48fzD6DU09hOc/nn/7x8T
CbAJkbI8e1mJX34Zco1565ILpFropPfIio1yoYf4k1NVth5bnQTfZ+AxHsYv0grw
ytby8kimlnST3qm53rA+G7aScGIZxsjpieYJD2Y2g6sgpbDoC0YRSI/3y0Mxe2+J
5vwSqKnqBKfaQ3oLHsCRCi4iB2Fzw34cQKzDR3nfnoE6ENv0arbz8TWVSOYn+B3Q
UnzbG0lywfui7cMKoCUxJosBhFl0zeR+WRqljoTcmzE4N2VmM1t/44YFy3AUEKIU
qO4szNkrE8bKnRbnq7E2UDtlzq1jaHdqI7prWG5gwVDtepKKyJr5MsthYkoelmi/
EB891RkSGKufRi45WdffF5PPt9EKlzyeBZj/J343l0hE1lwJekL4561ctfLs4pDH
8ldhIuSt1Xkh4IVgMgyMBtLmBBOjl08tO/+zO4wiVGu/8IdSrIBU6fdfae5qqopu
vHxSn9gHuR6l6u1pI4lXwUz7e1ixjYXH7emsM4umOc+0SpBx9Zy+BKNwW8Pi8HVS
sAIdL1dPpaobooexLTiTPLCYtzVAghtKMXceJzGw8IX9COq2PJZOD9m1bgYIgta4
XsbyLjvfl+yQd3YfmQfEAdnOD9UNwaAh+IePhVliiRUBrlVYzc7YSYzWFAoQJ0Tt
okDBh3JUfvcPWZlj7CJ3fbJxle8Wp0kApkp0WzZkYII+rUIpay8+owj5koiV5HEt
agskE805IARcKrB2ZiVa4pF6ndl4dz+D/EEf309kjcJuewfdtttBVhF+yOLSd/4P
fKxUgVqy7yASewXrKYjOXtSOpGaME7W7+U7dqr3xN2D9eNn1HDUvCfFxpUj2qup+
6Ftd7vvdPh8ELCdHRBYYxECfVCRUkYz0KX5oW22PDG0nzpLSyEMyiTBZqSEsqTMA
IuyCzXEqF8qEtYfOSUZCqcs+o2l0bjiaS1uwI5Zt1YtTw4YQ/7hhDObLCNr1R9ib
DbSFunFuqxD5lV1kKQ4YoiaFMTUeAS9jxQ/2eAUXcRcOoW/DUw2Xg3mYMgrUMJMZ
KsEHMCEfZRECIQazegObL41tAw7zKrYMu+vijQYizTiGuM82w72IAbl2yfkjrG08
GYH6dRkjYk7yjjq9R2TozZdG9ibM/QdcoglvXedDydFBjLxxxrpw8PCLy1X/HiGp
AeFjY4RzTFzKhyfSwDC1ArEgxPmaLtlI3SqFxG98k6ceWxGzjG9uAm+1XA4BPljO
Txc4miP6y2VPbI9BGgBzQN8ACjXQsN7PCxYH03qJcWxrpz1HNYCGmmTu7wpP0KkR
qfy6ekNX3r9OdhBNhQeN+GM2P4leaZ0wJBl/Qr9ZZq9sVnytumTjqgWxkNPwUgrE
YmYrjj+HZfEK1YPywZQw+TFBUqSRt+KTomEqRdxDctmqmDL4Nnv3UTgQv1QtZFP9
Cn8FHS0o8qlkyXOACOPzvnqfAnU1B4F3kW7kjDs99kq4OLejXvNFBpymf0TMpoIE
UPoXRj9sWRyTyU2ePhd1ab51mQVd4uPlAx4zyno9tEMAzWxpjUbvtFwrFsUlYi+H
3b5QoXO+AZBYbUGmP0qmwtM79/PSD8A3LfXzFzLAhnp4SPQUX4BNOAs3sKYUOOXQ
nI2tGij16JSsXdjUAbJcousjvt5DpWaLM3LD57m6MhfMwp9QvSGPHzJabO/iCMWd
f1NLwHul3SyHQeHbCqoh9TQzJzoY1gU6hWpzBrVND8ZZbt9kBeP0Ph40DzSnkgAA
PfCoZE/mz9J+tLshWA9CH+LnZRavMtuagZScBlNfra4Xc1HTCMig3fNPcWSNxJYM
VZn8yvQQZVNudvMmrJpTWdgAz+ynLMmOFm+LrbUH5F2Sdos/GDCS82FbQeJE5y/g
MAH4oF9v1VFco3PsvNkpHJFfJZDtLMZBcATAJHEOvydM7/pTFdTkstSdCl9rpoWM
ni0jywH00lP6M5mzeiAWvBnTQjpqRUyhIo87n/YFj9V72bc4Yy5GI0FjOhEQ4C42
djJp4yUcmaBgN8SxVRJaY5njZKiBtgeYGFRvYmeN59P/9ZcVGzzZkSAxL/cDHuCW
EYVs2JFRWydXZfmDnDp0SBvu4/s9HdkcLF1urkMIaSFR7MTaY0ix52eXche7KtLj
lWYLg0qWqpHl1j8tMaGIA89iUJRV12xdGtFmR3V865COyDzrcOi6YKEGDNUr6V+m
22L2+SHcGXfyPSELorm/ZCvvkS2ExADYbZntY4AdoHbGKawq6/gd5JsBuDOYbRCa
VtPvu6aMmTf23V5d2YIo58q45o30PfQ8JLzMOXnI0mCsgffrr5B51cePxPUdyj8G
dW7l3yy4BDpga+BgczLr1ICu2Y7H2tbUuR2h3UM9zVU9gqNM5bcFsNUVtWNg7wxF
G6VZ3Y2NvHN6ZEIN0rAGae+MZkv81TotzOV04K3gHt5bc3AYr/Zfed3IAh92KLj4
N8QHkL0FlU+NCz5kBrc8mUp+2JJg7ydJstSchg0QCV2OUD9Pdxlpr9QI4FqUECOI
o30BhSI3dNTRDJ47q5eVjDjjGjKlwJpVUUN48H8luY6MRSBqgMu2YN8SJ2xccpbY
IaVgtWvvihfRpszPxUDns1FvKNGOGJrW0NgwjZqZfB6UO8Pu8XQKEFvUBJJyFUT7
BA7JJ23IoDRb0WdNoK69MTyyyzkgwaTqLPYIbdl9XWcr1euS6bH+aqsz2mLznPot
x+3Ulkeglgrvry3pIPINO4amjjm0TJdSbSz/BEjopqsXYsg1toVUOjVASNOHzfDe
jEKnL5q/Rasm67Qkqm1psLRsEwRzEk4ZF5sf+Ur635fBJv0hiLlQ0tm5k0XN41GQ
T3EFtvYLGiWOHOc/s/mNm1L5xq6F+HqSeDM2x6gpWFlGdoMi52GSbNpetHVP2LVh
a+KYWHd3iCQpmVzRxt4/Qh6nKQBLl2CYhj6/X9NBD3+jmtt1TEkH1HmmR2Bz91gy
tfomkdolulzLMJnf5PC89auvAFCBLLS5A0mBh6Hf+N7I5+pSjoB6iwSXFodP/saW
3RFg1tFWOCXQn2ndA3uYqJKUw/LUm5qIgh3rHAiFtBaVHtxwc+dBdxLS3gY38rVT
aqYseOKN5rp3U57i2e70Vg/N9SnQDt3maaE5RlY8LZ9HFjCiKQw4biqctGqbw97g
SmBlNvQIjjOz+8BREFM2C0WXwWC66XVlQEuZjId1s7vuNZgRV+xll8kgdwUlVaxP
6SLcgVTv5GATltkih2/RntL3JblRmVVyb/o3kaEXDdl8uh6N1jQP989Bqs2HYaAf
s5MmWDmmQT7fg7iInNsAoxuqwMetZs6e1SDpCqCvbr+1NjCpjkzzyQnXdkt6XdW7
P87SQOUccF88uO7jY38GZOgUPnvET72YiY6nUanslDXSGsX7HQVhpc3EiWTLJBRj
P0kBcqbd9t/ycQL1dj5D/uXL6niBNP5GrW5SCbW9vWfabdS8wMTjd36TMWlZXmGA
kKU78HX3VIzpNzIxLpSbViyjSLFPNhwlQABKu7YwcmzuecqwXvKJ+tzkoMZ4yBqW
MVTDnNGSJxN+tPfj81lXuGznFJZjdHGvZGTyDIf37UJ842jtXEP+HF+gFHx493f1
XRH/Vd8KwTBKomGhd3E6/T+Q9A1arCUwqbisXQ+hloKUWojD5bgSQe4s0fpEZOwl
IBOXxk53J8EdySFz58H8/zjhIvIr5qzWN4HB5Zj2BWiWu0byWcw/gVKXp1zEcQd5
J1zPckmdW7T133wAaUwrqIalhmtPxa9b8he2r5spSVGF2PuSo9QcyYXWLjn58ftt
H31OV4IY0ea5tUeP4ItGBs97qUxWYlRr4hWy2jLOeBHsxgsZO/QIjNbxVu4Wls47
ynfEosiqIpiy6xVXkjQE0gUp3ynd+QxE+PBwoTVschovpP2aJvsu5zC38PfzovX7
OcC/+rbbPNXM/fibDDGfAyncCuDADznXrAhySgdPdio+BTEI17tVIqkVMA+RHgX7
x4VxCdG2CwmZtAVruPMj7RAZZKzKua80ToJi8XhZRxfQj9gSeuuWxxxoD/0WGV7r
ZlHYSulD8+yWo7K3LtLH3BNExJrNHOybl6aPO+tmT/5ugq+EvWqQadVu4jVwKIBp
M2+oP2/Ry02J2MEHq1wxNX2oON4CEjLys88lsK15ge2OHS0io9YiR5MZ1CeTXPm3
k0TJ7iTVTs1zYZxQIbHf2GppZUv5jU3trgH3C0By+vCxYHQfcck4dktUoN7vXPoe
F5SMRPGZ2e07l7rN76FJsEBDzdyhk94Ns91rJ2G6rhSFvRLjNJKsPUBDpS1DOlTZ
tsUrA1u29s6S9XJoITQG3xE9YYI2aEh1kC9X5peGiwROAPRJ5cfqcuNQ1gejjr8C
P7XEz0bNNFJx7CPfEO7xctldZXOF4HCa6dPvphuiuUdByA9NJRHW2gfztZm60RHE
9hlqYY/dEQeBQvdrHuIL1ET2n+HqSjhwlJZ4bbyir69BX9ZoOom7fd4JU+72jWq4
2HDNM9sYNSR/hvuxbAhajbUSjvCZxqbWkvsTdbPyq3g2o+7Q8LpEk2TNB7jUtBXa
mJo4WbPizL8RkGUX6X5C6UAq8TIStQ6yB7DVQuodOnRpXmkOzcZvmYSz/+/zIwRo
lWZE9OcjOwfH88N2ut+EY70mI6rMHdbkXcojgeMiJC8e3fYuw5gC6XtoTeGhzcGo
XvwflQkpbA7jg+Vl+nIQKpVUJeTiogcGfQtbhMfUGQRfWZye62OGw8oMUCp/83/b
Ebk0VfxPrq1OT8zTfHDT2/w8KHaFlK1qHGS9N9Eg+8vBXUNWuFH0HxEnmJNADOJR
wVV2MfQ5Ogk+iyvpzYRqsvsGd6k3+mTq/2GPFOvEn73bh4BJ5vLZC7zMBfuYk9wk
pM7D3lG2BPjBQZhuSqc2or7jVu3owWA0WKw/GdVPw2aRoQdjJvtf0hfT2BpV914+
Zjyg++1wk+idi2mHizmOCOBXOVMH8SN2N+mIO5bpOOi1FTrGVo9JgpS3AbxdQICU
Fs7i1dKcYRq+Y0M3IbwacKpdaIk9sMisRlX0D4ffSuEpRmDh0UGPuAnmZn5sCc7G
GazPrJqQBfGviLLw8GOUQaHQcxxxuzzqgS8CCOkUVRIXoy0/seRx6rbX/+yDXknU
hZVZQCmfDIKeRBqmgWPNlHTau2qXkw4fjrkkbHvuyIVcvMIF7okITGTyEtoYI0Ce
mgVe3ZSZ9YEc3jJm8OQKQns4OpBW2tF9JnekYuQPuQUvbCDAaJ5Gq308549xVHpY
kCn1gcZ5ps2Ml7CYCDEyJZYQVGLenN3pa1wsSLgbLqpkp4XSJE+wIV5AmWGxaWg4
JiVQYGnlhWY/QzktbVX5Zfhhobkmj0WdtzzTbNRO/rvcWLHwjaOOljWwVEsUuaxs
+M/OzpQFgeTABKVWq/mh0u9T4Mo7sr0Hr0szmYBGVfpP/AAbITiDunECh3nC3Wrh
Et4SJ73bU2iLb2zQfgG5fXJ/1YXiMsKROkRDpU4YXwuCd/QQPkiThfPgDWzCnBZG
tMqjw63q+eD0SABVcQEnkk1gx5FexIsaeH+9NGW2u41/ipGjN8rmcSRMFpmaSGX5
1isIo/onHcoHxEkOtZzTPcRgM87LhzM35H7Od/bk2yCRenmpFxqkmSdFihsNItg3
AMhbfjZtba2m/9qCHv1THgS1hfLUx1zr0vlMpb9Wcfj1Qc28xzXLwZqCBTfBrrx+
C3xOqgs7Q6dk+5gkSGiDp+mKNV6HVGcWDNWZL++SdhBucxMrIdpIDHVL/ZZq6/UC
t3ppWrwdka3+MdSlwkE7rUNp0AfgFr5nAF2fFgqv+1HSA6Vm5PjqlagonwUonEkd
e7mp4JN0o/29GyWPyLr2E96oSYQloP5I/19s3ORJdwSLmcBsnOGexJUbvTWTzZC1
KGyHARYpdJM/NCNfRDMTLc8/vOWTBU/IU6F/hcmUMnGymHklHLWpBECUdoeIG1Ji
EfUX7c83b6IQusNpJ2nn4N37taI5Sa6EU0EjUNB2lokTtDh1yZp8wTQ1+bvioHLl
5QeKxZR1PaKbkbduFejG4S4h9agJi+FrGHsqpPFMNMvZ+KuxbVrCnK+V8Z6HrCZs
w5anVD2yzp4Bw8IkEbaXDvaqm6V9zmmm8bsDnx31ZYrcDd9BYJuKYyWJAC89qI5B
4hFvnUS6WSsXPnpYMRK8wMI5RBIg0Zk71H3m1LY2TNNFyR+jLN41DZZvmnUrTPLV
zq9GCmv93MxJIEgDKemsIV8p/dUdrbVDQwsRdtyXwK+hTvmuj1ttrPJBqcYafc7U
eJ7b1qpVd1d0LsscxdC0AHTH0Ymf8uIXWnz0b9V8N9SUA3oQoMpLrje6vEbALAOc
8VeMLPk7D+3tMnED8YeyMK3YmFrpIPolWG0I9At+4mU1w9Aomb7NwpioGDvJERvs
PIbBpGbdUIJ9X0i2Wnx+FuOic74rrbQ3iVWQpo6ATpT6EU4pZJife3GRrHSHwyzA
DZcA8YuDC/AY1WIC35G+a+IKpCE1fdo1Jn3YC7LkXHYzZGrq/HqWVcKiYGdcA3/i
L/sOS5DsoDuGxwc/qwpSn2jVhJC5WmGbuOuh7VXWMYpZwZTkcy8jBUGTbbKie7I8
71jVkV9YCgqaOIfg6Az+QAoItiFVSFE5aTI60T8lgdyHM3ykiJI/I3TM30UrNO/r
21fT9WesPMAY8DPHFjmOLY0yxY7dsxJTtB5i/rbPvFpU5sazJ4TgNLkVa6YqjpjX
QyB57zd8Q0rHftQeBAK+cOZu1ZHRt2pu++hzgnYZmckwR8eONvtMVe0w3wczBhyN
0LVXhoDBO3007gue2lIlT9G8VIbP9Fcefnq5MOGYqQo6xf5mS+hDWzMWmnFmV+jm
Kz5nMJBJG0LzYxlvsXJQa3YwXc+tlY7jRKcGU9h+c7/ahSRvBR8jgnJAe9BINIgd
cZOPvfdQ6ZEwHqkyvpAx2jGFgg8Wjwp04QemAc1KkstvhZkayrSgqcUZDiv/n/7l
2wvC1nNz9Cm+2s0xw1MzTkAieySnsJ679QqyqWpVuIZbv+qWjy5TUHOLa2N6p5eN
CYEKsMBqKevMlz/ONtjEaDcAj02Y3WmT9AK14WOR9Or5UpjfVWQbyM+Y5QH4+VND
oiHmSfNJEBg7J3visFa1XIDbkxleIO6zNuOvhMl3V49yI8xpsxjf0N4CvFoXqigg
3LFubOjhdnNS6B7X1nnJzJcAsz9QSTpk31j9bgj+ZZLWkDa4RUBeOlNeAh+a3DV6
AIBVtuHPNjRj3V1D07kxp8GbW0gJdkLHa9KIp2U+ZU5pw7Xaq6Hn7rTTwAJ4IrXZ
LKBT2subbWjFxcm2oRxoDXDcfGd8jrGmDVm7rCk7EMJB1FSBIkRFzWprlqMNJcBz
uqyFsSLc+zkNRh8dreval1YZOB8rO8CY6I+80eYjfTEY6aybFSGApB2Km/YghIIB
U5fyMYDGXgL583O4rfAqR7iT0gV3ZxiNU3xtKpoiT3S8Pgfl1QQodL+VajdbYMrb
al7kbwVjqV5/1Mt8RZ8AtWpk8ZwmhpUS4axc1wY2wjifPvnVSqheFWIt7LlttMJ6
AayigiuLIXpievam5Aaf5UiHns8TB245S6JFfns3LATWXpQJzZmf8Khy+GHWYi9F
DV07Oa18I8H1PyAl9FEZXux3Zc+q5w3liXOYSRKlsnlvf79v27x1vfW7Yxe4WVT4
4jFsekifIY2I5ySl2yrnmPyT7c0yzP72/zL04kUcfht+XsuEiA0Mb/xg87aay4OO
FztaihvH59nEF8Md8a2SGo+dFyvwd6w8wLZQyfGB3v4CcI/fpn8yi9myWFHkEE45
bMFD8kZ2DIUBlaD/QwfaYQKJB3ovnwUvkRYO35/s/xcmvVyfo6bWeHF0rq8ztjho
qAQw6sZjz0Ms+bEr0I2EJ01d+QYwOkn8CBkaGHyElVJhHjjsok2mreswat4jiJHx
0n0JF/TC1YU4HHy3wGkGEeI9WIV6wSFPdjgjiqikPrvRL3imaNgate83KoDsbJaE
AdAjo2x/iFSzMQmKbmcV7m0VC7zd1WMz/3Bw+Olrx+H0bT2IiA6iNVjYAS/xsY29
gjfMmPhwxLgiYU0FiBgGru3w1ilL8wUsJ1IwwIZVcN2ty3dWHa6lSlgKVxCrcURH
Symoz1DDItYzMAzbB1igDYrirApkZTFHZKZVLFdzDO/wCCJiJ1l+VdeBT/dEPJ/d
RtjZ20kCi1NST/8C9umE+8ZlmO9jQl0/Xz4FQQ4ZSyGcdt+DqQDawkc+lz9f9pIh
1xQigalEy2RsLmldE2YnuV+qJu7X+d0j5MRvXG3zdNomfjG3TTm17wt6nCS+G9f2
TPheiUO5EXg/mDm4wiCGMaG8120gtJZWMnOqiorwc8h0a8BA2nQ0UnwlauWtg9ED
xkynhNA+gw0OubQC3gKbQmYi80ZsSrK+GeXHR/aQOSp5rf7yVhFDAA45LqKDLOD4
dtin9YFJGGty0kH/7mh2sxkxO4m3cYSpCkc9TDvqpI962phKoRSmVZMDDGOqP5cl
Aycozxg06xyWHUereLPjM56we8EJeJ0cKD1xeFLfSviGUXAmqjxJGRN5ZpIywvb7
WcRRJihlR1GFkcb36zf9hrpdCk1jj2FEIy8S+bbjvriHzZb1mhdO5A+HFrZ/JM5n
BW1g0MOQpK8wgc+QFc0tdOhBBd0kyEDZ6QygS6tsir6dO8cBoMzmq116yWKIc7io
F/LDHmQfvJh1LBvOjtAOjlxJdtWqmC050wXsQA2+ZMCAow3/elNenfd8aEdygxSe
qMftJ5A9ZOy8z+83QCgHQcdMfYDNpZWGJhEJ7nfEnJ8TML8/8K0Vw+hTWWLItnsF
GDfk5JOzyjpYm7f+piLY4Hb/GX2fY0FdmjrMnfgJ4YHjK+T9qMab+wwgE6vS5zRr
oqCxlFkT/p4FUbSBLfb2Ua0TLoB0X2KVVPX6eFHCzhtSC21krqhXFciwLxIEBWoP
teT2vqYSzu8SBuH3NvEMu8BRSUm1j+2ypnmi5Srm/1wH6vYZJICV1dby6n3hhp/R
E6QhD7WXRNsYvPth7Xng0adMv/pEFdI0XuAyGg0KXNy7T7BmpR0RK3QNyW+Rp/PN
+cEtISJRfSy0m0nrtUWkwfWeBI+PUQXb2H9l3Ufmw8mJsdk2x30l3rE+qP8s7InF
eFEbwBFhdqkxh+9AonA6EgAHiPnKT6XXGbPdJU4kogFDeC3e4zUV0KazP+0AMWaQ
YVjZhCHEEBwKtqSCnbOoh/Lct2szeYGZdZwd1pEhkH+Pu0e0IrSGrUjiTAJBS2RM
B2EmDjrwTQhVJFQMGAjLlgUZhPYKeNB8UQ/BpUeto7HE8ZWT7s6QKiU3KeIN+v3+
qNVXdcQPRM+eWw4yklay/qYeVt1FKhcViuX0NsBJueUciDfCYEKGW8t2/gYooPXl
8wS2j6QxHcwfCZKLuKtpWWCyfmjMXI0bwRy8bCQUAuNqCq+X0O7CBHCzlqPfqymE
fuoeUc2cM7iSqptYA1AID63kuwIiV/Ly3FsohMY0P3e2WFgUsIVOGbCKTLZhN7oM
yAvHEp2aa/AQxXsrWxAR9We9vvIQcKLJjeqYqJzO481+U6FDzRCmefR9jZ4lYQ00
7YHqHxVI/hczmBGQ0UZ4fhibeygZlCsSJvwQqQitv/chiiQeKFjmYsZJ4nJ+Hdd2
pE8rj6IOWUuS1nH+7ci54hDTUPY2OU4+ux2Zbu0FZrcjJW1BDP8gJqObcNrMyMQ2
rLebqQDqAl0uUveMOE9HR01+beKgl57igadtrir+Fnt71HV4MtNhmDHyEYLYpmF5
mgvP8NpFvS5l6/gq2HV7R3UBGaJ8QMVhOZMhjs9e9LKObPgZJ4AJcBCEm/UIQEyp
3OV0Y7fye2PszPvf8/+6V2PfEzxFbD5O57Dhy/t01x26b5FIZwjwowUPWGs0DrVn
3kTVnrf+1d6UR33TyG87O4bt6UtJf4sSQOIckeYXU6lbGHWm3+96b6hLtOs1d0la
6R9bGuOUSey8SzBqQrNmGl8S1C53FtjqgynbYo9UfWzMGtSDpdGbOUwnBV8hCQKY
U3E3TNfYOxZw+ovhvYoScL77v1cJinj5/j9iIDuH9hch5jXjWILcQ+IjhBlyZcLZ
ypbsC7oWIIjAi+QrLjyQk9EW7yps15IFm0a6pB50TpyvTJ7gPjyGXjjKrTClNTw5
EVxk7aDli08UaZ3RRq69jLNbcdebGIACf15KablaAP8OOqis4HFqekqFU7PU8VLK
ctXKaWqE3U3xzDaodDFZPR01zr1yQddhKngkvcn/TNkUlja6Z5VVg+43z3u+z81e
HPzdoNuO7QmXcPSDEMYIyVliAvjUWlRS5198dUd0I1eqU4fzLiGS23hSV5j44XQF
KaR4j97FBE5PH88L0HircqzkowWCAMzYfItqUgRzGzZIQUdeU0RupNHgEaQoIMi1
g55iRyaKdg3v0EfDIl3Fwx//No7qjpLuiHKoaNs5NabPpJsbU0azmjCMAlezGFCd
IHm5uyopFOWD+GcjCX+ojDf0jZPLoDrh1H6n4zOcrjkfh3Wooo7Ss7TRbr3X5B57
OLRFsDhoVZiUo8Iv6muiWHuHjnvxYg7dWm/0ioUgIWqOjhttgtrFFDPur8fCWsvY
3DJ2C4Ssrl3q+DDiIh01xbDbkELzCa4N7sqY1YdhQKF2GbjhoKY/t26JG20Aucow
o80imqHQEx2+Vi42NNigHDVdHWA/REb713wpKR9gRlHc45VyqhfTeB3Zsl7N8hRA
UlX6r4Wu6i8M3uDRvyI76qpvb0yMFKp3pY1SbsM3IIn+6ahiCGe0qMC0JkmP15nn
kbK98/o1tAQqu3WJ7HZleKLaa8ghgqknq6WFxpSDDiL4i+3dzgp0gWvnNXp3a/R/
iXUULQpMYatC19s8tDTqJptHQZL455Lazory3VUeIHR9b7XMK1J3cV8GqBRmit7e
BPO5opjMrp34X3vaJq4Mx6xPIAmBtZISUQrF4WD/IA7YlNxGC/e9iW0IqoiTY760
HkF1vAyuyPtrczCVNciqy8FYGvep0+cfy710xciQqTexSsnsgqa0LpHM9V2mqw9n
/ITH9posHVS50po5yh2ECls1m52GLEBTeQuXc5xxUptfspy4txay2E6ezPokjLUN
29dTTJGQq1rxvy1DTbu9OF+G+9UjFs2Y7ljv2nqKj3nkEWkgKG7eRQRPzU1/DRC9
WiF+CuLPje/bMUMSnSP1cj9/ygcM/FQ0DlAMnVau3SK9smgvbrUvHzal3sQqP+co
NlqlIYx53qQpcnFrUOAzYvMi2mQUK83YVR045U+6G9WS7+G48nzILN4hyOBJ7L7Y
4Aed/vO3rW87UbrkDuX6mWtPd9gaG41Hx8WzArlRBi3jeLfudnSLFA/rc0ozGMw1
hJEf6K0E4SWSpLPyqLjzPfWBigK0c7U2ab3UN6T0SMkhu7Uz384s3nH628dzW1Fs
MGw4ZDY7ggABIS72oKzUIqrRL7aq9S6cvo8KpULFp4ww02rCILMv84eq7dDjF85x
5SHvwWn3l7Td9LJcp1HeB8/HCtrerkhfDdZEGcFfqjhLN71THta4BhLDfZhBwy5r
C0jY6+mFyL+xsLvpJG9NN40aEC6WJfdworg+rv8oGjSUANwA9q0bQd8/KZgVTpI0
pKHrck/jlLwM2NQKoxe5Pz3MmuFUo0juw58+12esr9eeKTahxZbgizlpNQGk1XSV
Oi/bWfMFCxDa//Gj6QFZOkKTbmOeMiM7jKbu/2qHQgOtD0AFgfHvKBkzM+2QZnOw
bwgNTkSwJMFRXviZHEYIJD3+lkrSazzHwLwFvp5r7ZM+qgNdR3GTW4XFMLsv682t
BDcLe3eNAv5YLe6s7V6JsOJTEa62WVCbH5RwCDSW0l4kTM1mErQHiGQUq0Ma4nCo
FY0QAUIK9W0CAsWBX9iqhAJ+edNDaRiiWlANPz5FVvC5zsiBqs+Ebdg2uuHTog+S
0aQ+B9ZLDV6/JFI3J7L9THWqxNi4Fb3WRmS0qOvko64wNdWRhKHNz8uRH9EzKBCZ
X82Ie3IAaz1G4QWHz8i3U94X2W342r52C+t85lYdoF3ub/pB6Qyzw43Vrkq3E7Ag
se7F3YeXvp2kBTdRAKMDX2/gEVv17LTO3aODJxk3UOE5dk1ZE7RTyuIVB+DMS6hc
SOVXB/xnYetAVJzGQEPiZVQ9ee4cUW9NRx2PbiC3qnxanRbU5tHgKjssTwRwTj1C
qKHEPv7Vz4tRypsl1sLOwb71D89JYDsKlxDo3ak6Xhq/y5buMjDOqPsy6nLmPnSW
O8YFyY2vEMmg2p2U00SW1+rUQKLVuH5L4BZe6IZa53TGmcVbmjRNKoOspMDgUO3L
jPvWSrB0biB6MMXFeEhpmxQYB651VjnbkYprWFkcPujcRAOzMPYoi4xHsPvX+DRt
cn46tpMYiH0OOa1B91mbEFGrpFOP3qPLmQEIno/lAUDAbNz7H59Be5rIEMtSoLfW
4UyytDTHNMwhB/vWCbHr9qgEnyHkzNL7V7CSyNjcpweQuoVEyMOM1rrakxNexk/E
rMr7AfYBA6glxbbyrElkCHsU7tq/cJLiIEL6xkGhUSGbk9fhrSF81+955jbTAH7A
b8HnrBk1aTwNqqe5ZGxnw1HK0eQCilPufns8BOYFy5n+kKPIsuTXTVynZcTfVDvX
55jxB39lGyhucZMNpP6gp3H3105h7LoM2MvFQ+J/yeJABPOtphkNFqddhFS5cbzJ
Gn+Q7opzmvDqChzK537YL1mAe+1xzETw7zbHNBXtvbrBKrKz82MWhg5IbCtPeMzk
NXjflCOLu4tZ56Nj3qMnfkCvm1wwFrfCCCCOYhuEFMdNrep/BzcQaRqKqyOjbp9o
zgayraU4rDNwnGoqleaEFFRygdwIMLrpQXJuOcn7EmWX/oAIQQcOwMMryw+ST5lH
vvyGaqTYVvoac3OvhzElmviFGAcHjPek1iUOpM7nrWvJlITKcqICDGA8PM5DIK38
3y56KxLZE6UtRyYYyzeWu4eGwlkZZEDEIVhTuWN+JtmeW2j+IISmlGoOoqehiBFi
p0m8JA/p8GmpZJ2BsSBxWSz/ablMSLsz0H1I5DOc1wg2wPqJNopxJ4DSOhcAWjj9
neLtPmljK9/f1pJ7S8TJdgvdHgmAFITxZzBHMQOm+xUrvHzHb9ZqPKze4S+9tKcq
Z+Ak+RAtB1amMUSGHf1ssB+H1dSiS03pUIMtoJTeUuwjIcfiQfbQb8jA1o3NhjdB
yifIa788+R6IAAPNp3CpozNp3K/yj0P3Vjr2u6DzhSRh+qYku1O/874LmDEIbBEH
iM40FFMxrWSEEusTJZwhU/x3LjmRJRxcAq/Wwr33waAeNYcRg7VEe6kY0P63ahxI
UTAQgMfQIMyESJStSGil2raSNSMdRX5ZStNJVPit//sKjnzB9FGcvxSEG3wXOR7T
bIZHm8wZzEek6DcD6ekOxVKQyvsZxB/gLquglu6mELHPjuTonLJINYpppbMYfRN8
cwKelRydFpMF8C5DCHRaCugky9BYBOD2kVigQqYp/UFzjNmJuKvXwmDRPAErmCUA
52+BUJ3VPQ3giyd8gYpndbtlVUS/R1totHrYeNoDUmR/JF5Txo2N5a7/dO4G6Pkg
KEpm1RfVbmNCpJplVmYgkDdkiUFbeYXXLWcOVDFgVo07hOpA7XDmJjDTSDElDDPy
y5eTXOHDuHHw3/PmsYq9v9R4IdYukF6/DOglPTZZMiTxbypne55vtbaY6U27HjEU
+N3AkCEHrR0gBTaRScFK8JyN0BBmOEM+N90WIZmB45frxYI78akMtYHKZr+rTfgD
lC8QWrwFjpEXt5z9v5bswFJ7QHI/Qjk3YvgYwRQh+qvbsyfIQarQpFNNlG5HeIQm
UxUZjGGPNCILeJ+0qzDw9Y4LyDW5UBiN93zk9K3nCWnF6V1aYxxF0D75IUa+ruvq
M7ORy9kkrcxaX2ut+eJeJ8qu7WdCaisvyMER8L1r6Fd8crJcYWW1eZCXP3Q7gvyh
n6b6vxQQGzs5/fNXP8zHAKuQl9w4gLUMzZqEj40z1dVh3JZc5sgVA4TooECYGXHG
0UkSbGDe4DFhRoE/MpWGtkd3dN8Ma5vPdyaejAPTWjSxsTAqyANW6RuETL2Be2eN
hzZISsHm1uyX0PxCna27jppqV78a3abIDyCzqqBYL3KCH7z6dT1JV7U1BSbkm0ej
DIW257tse7EEEszZGwTBpvCqKpz+JDOSc4p5vMX75ifd7hKnJzPr4cxnwgHk/nAK
QjdeveqSLYho3BcV87k2JVeRgfATVHP4DtFx68sojpAN5LCqYk8Ln8ZIM3zPA/vU
V+qki+hIXVvacJnZbvmjSP2LDy6BKuaGfxgyviRYGSgOW4Rxq8MAmSdmSALtDL0s
QyrFmJrEzeTq865D79Y64PaL7bxVvt+c9Z70lTyH3a9wt16dHKeksSt0TTUNxn+Y
ffTfqm2eeNV4MgrDDMEPswRRb6fGLqF+5WMNGG8dWdNorLWR/VwntubHxcJdbV9l
IluES2Ln5KKEmPE3pwq9/BPVQEE7pxHEzbWZv388bMOoME1QqeIcGkWOyLN6JkLs
KL4u1vst6tE8Bw9NPapsM4rYuf8bFrmie9EAt9yhHTbF3DMIpb/EQLbR7fczu4on
f/0AP6A0SYnAwWGlYxHPD4Fw4IOgd+0M9n0xXdWjYdSwm4XNb0RY0hEImySy2GkJ
7RggUv036ZZ7kr/kj/p0PDcrGVc4Dh375XaaJQYT1Tp0k9cksgpjfXm3OpTe0ADY
iXJV16PzKL/P1G9oYPE3GFv7NW0PL5sxu8mQWVeHvgComjX83JB6K8L6gLXD+dkE
I7MRO/a1ueEvTbYh+EbtnZH2d0dGj3QsyOf/gyzzlgzs5y4cJcPcueZTZ/LOLHGL
Kfid3W1VEAlRb2T2baarpOOYpXuINNO0O/udxckgG3hA94AV38vPSFqqYH5LsJ3L
5591qZfJocVWFhS6hz9fAo+k5XKdd0yKVgXOxJpaVhKExCY3bbluBU/93azTPgso
kTpFBPv5I395iB3pD2FPy87pmYL97oUc637Q0Jom4ubAgGUNd+agjMugaczzqrT8
+GB16IfB6jzDrLnvpyuJDw3tqUV+IzlFx/AG6waSGDooymaLyuszujzogu/sk7n2
bS5JM8KdQ5bJZA3+7JTqz8QaHQVlKPk0jWH8NzfAPYfGS/myFqC8d4vy9+anWbWA
m2ARst1dDcQwYtxT3JyT9O4kmrhwzwr9/Z4Q3DAoylru9yLrCs+MMSKvhfL9z5zz
LjYy8JdXsFqp6YzdPAEU/TpQEyVx/xVNrRZsRhHj0X5oxMx0ov1U1fgsBSDHgVov
4Dp9wprCR76fK7cE9LH+JbQzLvp01P+NIPC1A6I8cM1FsGARA2IHtxVigGhKiGmD
UChTHTY3tp0RxhTHkE97g26u+J+smTrZMqPjDKb27Sp1OMGiTnNmK24lYl2kR3ur
wSVlwuwUZldo4ld+BeWU/lWUZH/eNOo5Rhf4ss8Lw+mRtkSBEszVw6lD4nD91YU4
goJ8TzRsLq1YMAu3rnLptbD6gjJ3RIj9OTyTPy+Lfj4Nrdx++D16TzQHeiisYh3Q
4DQCreS1Gl+PuZuNCZ1fO0IYHAStEFrzwuExEq771SgscMvdM7boNK9lPL/DtY4D
gYq1RsvCw0JgBYco3fFBhYMsQdXeeg6EcghKkb6vrUVLYnPVSvqmzNhrMVCOMGyI
Uq9AbvhXkU3NIkiiFnuasPt0VJkrFOVAcwX+KR+mvnga6nVM7LSat4B1xKGWCwEN
/RWkrdDevoXzw+4Z4xe1TCcp1T3hAtZw6V82+jBdYxPTnapNwBV/qpNQgDMgwLvW
3gmp2/uNVztZRgyfgB12hSaXkElxfplFH2RXrwcagv3VkZjQbRugFVwqhsKp3Mg9
vmMGnEmmK/A5UOAi31qngFNZ7bEwDeHGz5b3mozKVDIup1VfxvsR7Os3iIUfvazB
qVCE2M2lskUiFhqa7CH8kGGL+Ca+qoLi37T82dUaTyWDRvBxVs8jnTnH2sETZvU/
oAPC0sQgQNRcG8uOjwfVbvomDRv9zf357rp7mF/cKzpxc8JB4T693OWOod5I1fwR
2Fd9CWJ+xe50mDDD6h2ueuTrkjX9rvvZK8h7uuozr5LwVX7JYud+L5rCZ2Kk/ia0
ThUWD0q4zskBCiR+WE6akxw7cJKuxmPdTC79yblTUPTBNr+FhksvMm11fxY5iVrv
0nm6Wxb+VCo6eqnuYf9ZA5dg76bOdOc9ZP+bfqwoQpfWg5kHTjLHe9MMk8YwXnRN
T3ixWIjzTGRRiI8/N+sxbSCMzxyOxv6hnx5ipGPa7H6WbYpU4O7SuRJTExOatyYF
KhV7cIqLnfvNE5GAM5d/SiTgMSFTxNwJxzKx2rr6ezMxTRbP+I0WueYj9PRfArGs
3bWn9IH0d2UPcxOxvRfdyL4QJIU3auQ4YBWnqkydwF1U384KBFxT4DzEUQx2Vd87
1H8DE3X6zGVsew94INfTDpIialvdZQYwFeHCa7XzpdhbEhHTaFvUfZhtJD7eLiWH
vN7hEGYN6q5BbxqrYew1hg==
`protect end_protected