`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6496 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
HdytKcppDjja7VfYQkCqvAEIqi+uuSb2hcCuUIrVDosQwAplNJ3u2F2raKAeZqBu
iYfzozxnEf0S72sp37g+dCpYPgU5EON8ICqPk33GpFJH6qk44ogGf+UaaqgC/Pdh
7aVWI2Qa3GKLGN4AYgu+07XLDZJFmkcS2IN8AVUipF+s6b5mhvv9K5ukTU042+NE
t5/1yYS8gUCEBra6QY+jST7OZlapsA8abhS/z9GB9ns6J+j+/YITqV0m9yG77Yv8
0AjlWMcvaLioijRwdSkz+w8VVZ2nFY5WjF/TnXdRly0tNC6q2He5EcCBX3qqOv7h
kJiRDXIk5cke6Wm8t1H8gsb8PPDbBVB+ugK6b2iVFZ+T4ckkVM7WXDF3SprKl/Cq
ny7C0OUTRagabVQu5REdU7Mwx4f3d1Kr3wMXUAHMAlVF6+dl7tiqeIdV78XbKEQn
C8fw3WBE2ZnpQi3cp6OWH3lbjHu7PmKgknGEsmZMEz+STI/g5HqXAc2+DQUppcdK
+JkciveqQp0iWbfqHvQDZYEIFPOkijjSi4kyRPr5UBIldKT3LrwxNRdByA3fIDkv
ocqEMVAb2s9fdC9nwXZ6/gJb1dX8ih3Fsz6ah6y2JjB+jul9+IYsKPyJlktr0EwT
wV9eMBuQuoKuXlSA9FE9KCI1XyJ2W3sYunE6OM1aVMkezWH+2OMBv3fEaKoIL1sW
YoRiW7otTIRbae8msxLiDoOR1EW7mRavQqPdW6lgkfCqg7ENvXhbCnyjHY0s6l5z
sTmz3n6uZ295eChc8jA0SniE7ZxnvtZ4x4Dgx38FUsyOY3Opd1nsuIYsv5G8uWWg
ki5STeTGcJ6UJk+mgwLgAPYCRvaBJH64QMQWG2KCyC5vXhLPLlDBZG8Rtp6WaGh5
Nl/QO5755vwGWcog43qgl9gLRd/D9XDqRsQLqqDLbliByUdfY5eAoCH5ANYrhK29
dQ7cwPUnYFlZyTzrSDKLeM9Db97u7UZOlWkFmjaE/3PaR/Vx1fMSTRzXU7zlx8Wb
9hHY79Ohc1pM/xDNtm6mEdYiieuBVVzGArTsA+LKaYe4HMBeNbpto5Sj5NIwrWGW
Du54jZHgSrjHrmZKGoOiqNGFSbtcj+fmDPzGYHWqa/ESZjWArZx2sO2IhQ1jj2DD
Fuqqqw/d/xWoMZltrItbg6vWFDHNK4zofZlJ5QZMfEBDUS02937ZnIrLiBwzwZyb
XlocTFzv7RhxkjnVtBqkHSIXhmrJgIMuH/BJtXmCN8BzZNgIiVOBWxihnSRYr2so
EZV2dAcm8zXHYDbIgP26I2f3HCaJWuEiS8V3+0JKfV2N4p73ghn5GTU1aFZlvWLh
IP9CTNu+RCI8nXUKUMGPPDnHvR9ehuaY5IOJR3GOMD0BpVOkZoLZ6esQ9BmLnPtd
9gRmU/IacVUjcJiZyHkXXEQ85hH6nxTMfLrQwEUZhHO7pUQlk9tAVQAgvMhNBYy1
TzVGpZWw2Qh/PSNraIRbfQGtCodtHkWGhHA3N4wpI/ADeG1fidSxS+sDX+eeKTCI
zaHLdPU/H+75UuGoYuSvCY+KJvNkyyJuOk0aZoF586uBqvN4LxBoK1i87CNYbUpc
C2QGqURoHsMSyPSCxbHGeT4wNUJaI9BdAdFUvrQ21UoqEzAOyR4bV8JZSIvNsYdt
awfmWWgGWfENpcY7kHW2S3vsmkm2np684bLSnbadISsVWhHCGJZoZsbPkeCDakPd
ZIYa9kgd359Ctx7cxNvyyfhNsvX2magZADFbheE79hEp2x7TYQbPl15czwvD+ewi
zOq1IjkcQIbRf8vxuHRtn0lPgfv1Yh0xzm5LKO+oo8xqihF2jr5I1CWFHL7ecj7c
GkBeuAEx+6wghjqlqE1by9XeRodoXMkJfny6C18B03nA+zS1kMQqeL0yJJHLwiP7
CfYu6vfhpEWK9XkFM0v6FFqh+Am4vSvOFvCHYoQdxBqDVLqscsFro5C2nfUapMXF
vyY3O4FApKT/GO9jFzZYjLwa9vAvcLaCX8XWE0MRlfil0xzdx2nHCOI24kJOA2We
/kyl4MY2S2MwUXAZFv+FFSDgjnlQsi8Z91Ka23oIEV+NKkiU03tdrboGrMRQDMow
0cEhbuEJ80VkV0LzvpDhHTM6QHc8pYF3x8Hn5JbhLvbaAH5ALx4XAfC7/MyJ2Dl7
aQYGSMj9NzOinvaetF2dxVJ6tcqw+fT3CtbcJBHCYGo9Jhq5R/7AUnnWnbVZUbcX
W4+NYxBIFalzkVWn+1y5hLyefq9J7EZGtch7Q3+P/Sul69sNDAvLk5D/D9C/2F/E
DJqctS5C+OiwbWbUwzQYIfpZ/SVliQqPfUy5ZCKeG+vZgu7JoSUgpCQnkiGTsXOR
ECOwgecnLmB2DDlMPUExympUlSTCcGKbm00YcpdK6RXDd9xdWK847KBOq0/YSB9T
Kjwb8uUWVnOFToMTJdSh5Y5KA8vCXI4+gTR9FQptZ8pLS6HOu2ApcxnT/K6L1tts
2Vrn/DwWJh4HbqjtHwu6+JQACQf9v+KbK+L1k/oY1BEZkEbd9ypbrhyd65f9CSjO
zu/41WVZ0JbXfn+PQ7LpxaS2G1Hhyn1mfKZtvIsVAQP864KTBc0tTZsZ8z/ZjD86
yx+A9CubSKfGcc4iXqjqR44f9MaIeqAh5AHH+8xDz+ZrcWvmMJVSzNp8C5Us4Knw
+dU8s/naxjr0qmssb3Cg19wTxPcKdgHYPKwaWgyhcxnjwNfQaZhap9vby+rr5k4q
v0tbKNDzgy4nMDkJDbk9asa4MB0339WtbZdloQxukrrW9tdjolvFASVHaCFf78Yq
qp8vfbzNf8E+bq1eqO49ZDkT1gouOy0WwYOTuaHNAYkPieErb5qQZtn8RWEXTKzl
KR6cB1mr2DBH/fxc1A2csArT9ub9i+LPWMpWk+umC3HPyyB0dEgiEdwF0mHiaJT3
Dsg6Qqctvot3LSkrundLIiRolMfg96fUnOGTpv7YszvM3TOo1Bxiowq71Lo/UHIl
kxrrVm4veTA0ABQDvVsclrG4J381jefLDQRYSHZb2OOWivg3XLLy/VA1zENoqFTt
3XIdzhGMNAENUnpgf4GWdDfeFgWCwP6tIn+jQ59QGmEcWljMvZMuq52lHc2FPZhm
eAmOPuMG0PY/bunOONZqGBeIH1dpMQgWEQGTXrUitzZ4xah6n3I05Cz7bNskbIo6
9cN596ji0NKU6LuZtLAy0CUxEOtjqiL5hJuVECu8ft/ZHz3Z9PXiKc8wci/q14nT
GY/pdiEXUo+Zg4W8Thhp4AYaU5vhdJGwpSxaOj89MGrRLC1VBZsufmXOqiV0NZO1
63Q1G2DlUj9KL9viajXm7/wE4+my0LnCoLC7VaXNhTByHkLnSxozStbaorVYkLMG
DHQM1kNrnrOjqKXoCnzdinkG+scEVga8mooWEsckQwu9Iq0SyrdJsGJzlyWVjpqc
QPKa4Z45WNV++GOhhuYhcxIEV89SDFA7flLf2XqAvCb94mAxmOpzB1jE9HSkaeET
R+cEWJmH05Q/GdLrHmk48crLRwSXCoFI+KBFjbv+b4njYTX+RzYSAPS7p2KvFPIS
9nSCToH7SVhv9znsUAfB3jpcN7nsZKCWFDUNcaTzVYJU11GD4G8Y9Gln2WkSsdVG
O/6DKSs5Pixtial9W8zMniG6Sw/b5Zin56Iq360qGfTNRz0+6EZMBQqku/Z1eXRK
+1HYzuSZKwdBzZmmPB2PcHER84Cm3Sv3u7sFXBk/mSYn/A8HLzlpBFjb4sOSJbNv
D0fyeXs2xoubsDW4mO4KL4yvkJZJR3Xx+Wv8k0VeCkrZ0dz1/xidovi8tH/SVf1F
ePg5K6ufQdq1IqgF2kwh2B9vaA6p4m1ELtth5kIKE7FlTkluEAU/8eNyKijEuFHx
u9mBCJYW2pOtetek6YlEIbi9z6VRmxZdulPhR+DptW9ErcAYF5x9wXR8BhdYapGP
Wq9Iw44XI/ejvXr+3rPrPK1d2ikjhw8zl5MG598NLbR6KXaFjSZM+4v+Q8yHGLJE
L9XXJCNqL5V3CZLJiiPQP2Lf99MFauhBt+2UK/e2xBW2jons0PUFLjXy5+A71nBh
IBcVUobZN+DWhUk/ccMThApi9h+M8jioq0LzhqJZnj37/pbQSyvFIwu/7nSxo+JV
QIjQ3u4VYaoL3cyT6m6p5JT7wUfE0wdQ+yxlMa/TD/FymspJUlatxNsID7usCJT+
pLqvev0MYgDzxvpNU0X1HIZfl8r3vL8BYQwYRk/fckimbVLfpXnQrmMT2VyagSyE
IZW0gbstwt52a1akpY7cI5R3inigwXVejs3R1q99aZUWiaWS8rci8ERYaEaC73rp
iENeyiKIZvfeUjXcVX1XFDYS/LxBhIUyClo4IkokMrGk4UScFSaWfdGKtFAba1q4
emaxBFQLGY7LiTjir0BDxWKn5BncS4IWmgjVyjdZy0TpVo/TGW0nOCz/fHqonviH
bq+WwGvKuqHOYK8rWw9r2T7ozYVjhAh6AChwhMgapimVaBJFcZYh0sMaRXW9Nq14
f5+pT+1uDW6vAYByvxeo45Ied/Wijt5ELZJbgJnbe4jerOykFpyu3fkhl3Jxy5IT
D1ZrExrFP/sjZ4lxQpsocC+aIeJsK+zDaagpZj3Ro12Z7uSxrSgN1uO8J7Ono557
kgvn7gvX6vuXS78zZA8HDeOedOSB8yZIEQNluAcvrSxKRythzxlvHx4AdUu2sfCH
JYcqK4MSQ/PoOfuev48Iod6JMamkIKKkEuNAJJpNV0H4tC5fA4Y3sTFJequBwFG8
a+8Krf2MnB9u2Uyi8kTulpZKIOGXJPe0fWGN+5gQacnsNc0Qcz22lHyJenLiq/8D
gejzjNmOy1AOqtDuZCESKBAM6qEsINoQxK4Z6cWfyQjW1qsFnEpocJd7zO1AFJOe
ZxA8MKWNXo0952EDZjnA56M7Qihv3+iMcHtR17Y/NPYsCM4pA74rTCO0ULpmi8jn
WJ3ePjDnBLFPNTT9DSo0kgVoinLz/9NvQKW4Y/MMpxA8zYg8QHX0vKDtcUgwgboW
1v6lAQC9oqkuu6IBuBrdvVniJm6vmsNpycnV7D801phgLKoiZ/WxHuueVnj1I4zg
Pwu5E3qtvcT/49HX6QC8vyv+ptidIZGIk6GSJi+einy1DmpAZDNWDDWhdeP7WRVx
FqoKvuTDGJMULuRcDZ0UZBFgU1bBI8jWTMxmyKV9Sj4c0MgQA7Fn+e8r/6kLI0pe
lchwrnVi99W1ivYHA8w1HnraePAtmiod7Xpa50ikWBPVzOMHwrufymqd+n2RVwSx
hGTRt9ocvlqd7oDCUKo2cYgcTnHKYeLAuuFRgNLZ5aWcGMt/mZ+aRThTfW3JeAKW
lMmT8lP291EqZjoB4kErEiHne+hGoJR1yJj9XEJ8pqHL4JkZYztDihgUHpshYSj9
/CyW1c+1WdDmHZP8IWGVg5GUUy2GGTSJWHPMF7PuzMLg1ONEl///f9IaUCGstwIF
AO0HSo7PzC/JbW0fwDOZNO6qxN/AjHdHucJ+veYhfw+o/JfTKE+d2AghXTmajH87
S0OnUPJp6BdNxNmH1FcBuXbUN3EUJ48vFiz/0vcPqeX/m+FxzZ9yVmYF0TGjMGjM
YGrCic3HffLjSTxNnuw0XOmljSgH6e7fx/NpkeurF6n7L6zisbPcVCLC2xZW2yLw
MkLM8lusiD6mq3n2UKMNQpiqZIj2ocOWjHZYBND7VhvCIq2l4rweqlViVz/7m0q2
443haZWmF+BI0mwQKflbramFJpHbtjUi9J4A3btBYvmvqvBhgNBMAzVpUHTSbQxA
WeFBqJQSEcgSfK+nOCFaSwr7cKLOhtDOF+OsHl+pXvkZ5e0Vy+raVyHRIa4/aleE
lmBrDq+0TOcyflV8mMFjIetKBQVDsZPDDtDuUa2MFBUTXlKD8CWl5w2L2v7mvaky
8taD1wk6nxCDX4584Zutoq5oi/UMDQ8/cEFXWnslrQ7mwdyNh+WInyT7wOpBAsAo
RlHNkynDFZ4n/FttRiMgkpdUcu7bPTttfF8FZsr7ECw61U42+zp0OGYsTSLjwVw4
52H0ZiYnOF46u2jJAnnoSQA/Z1ay1FTh3UDKjbvRPVqEBiIWSDRE3L9FEVETOdVT
yUMVFH0vkQIMEM3rlFEav1Ha8KWaIsA4vkS1MmkPDWUMM6UnQB/l7ucM2vt2wyPX
odDQjM024A7kDksg8YVPqdWU9aYoBGLK/3UnnOBH7USNewsZqQdiXrJGW4bqYKGl
9jae8T/9u5w7viiuOhjJ2I7X1q94mOr9q4Ku2pjT8bsvWKaJ0LtYiBNkXn6oPaj5
Rzgj7gQ8UngXgK85Ycr3L1sAbbr5ji8DzeYWvkTb/LB5BZf2fbbqw3UYqNVzA6p/
hQ8TqRdPhAPNStgEdyqG2oNQAEFlj+3IBoNBUS2Mlz97kWVuYbMDO10Nmsp8sXRF
uJPUiBWPp5oe7t8fwqvxaI65n/1Qn0kwXyxvYFxFa890M0HCcagMcHue7xNvZRAw
L3zktEv4RW4NqYrNoBOSo+6gm1GbHJqX/pCxTxQjUtDAtDMoVVEN0alhlF9lDGrN
g5WUxl8xqF0+AR8507tIQPSw5qBqMzwSfv5PiDNJIGdqC4CiRk9WZ/fSPuRp1qR8
t+JAkBYR27QNB1bQe2jcKDKxVoLRDu6ju6UJz0WWJe0bctpsFl6JpbK/otY9G98D
YGf7tqBCY4G5VqZ6jFipapPThIL2z4MoU7B6sIU9uXfT2SQd9i8Dg+2gCH+WJwvC
jMZTsMvIqIxC4bn+icJQChno3L6YQpn/R53KZ++byBy3ClnI4Xh3SZZwO9qhSvh+
/pORReZ+EViuJ8qJdSvjvinyY8Mm3pcQEeKwLngwSgpSXuvkg/TQTaTwn4JLnWjk
p8INV4YETUJj6ROE+eH3qyh9zH9m3GMyeTJhsHRB6S3M5t1fe0qa0Pjxu3E40uPM
ZrwsQXrPHSE3/1ty51r70g/yFz28ggWnDizbgD0hOoDsxsVB5vHF2ev7lChAScLI
/hHQ4pFe+4RUFhjtGd7Ygdx0SxdrdqfICW1oiz1wU8mQmFpzurS+KkKdlCxYR0Mt
pyGCc3xXIWE3LADhmFcPfd+2e28uc0FMSnq1BBVWUsaVwBjt+zAe+AUsMJ+1wsoU
20l9+MEzr4h3VMGVy4jeBhMwLvy9hbVP9t5TwOUeDqKkAtBARSSGoEM69MCivoyi
N7PHHpsFru5Xd1BWY+jFJiFws9h8Jz+Z/HLdapV6CBEK+H7tsxoXYWO7SxbP8HTi
FHwu+bvc+w9x4v/H5CtdLRFT+rhncRGBOckPdi+vee61S+wZdmXNH4XpKa7IiSy7
3EtXknwsZJuEc9aky4wujYbC/pZlYi5pl/SRD9nw9gkw/ID1hhvFHVK8UG+X7b9L
Pn48TF2WrJ7W0IYPORDo7MZQN/66DtcEeDAwzUa6vvBUdk77DZFyQpl4E86sLIBM
LO+SJhFtx6FHDMuC+ElPTHZJOXd3iAC1ADPPUtfnDSKZSfylbtL5ymX3Lw27CZRA
6mng+88ZWZEx0qhff9N+8AGv8UcK8mqf1A7cScQDccpCnLHIUWUWP0GQHRhfklEP
wgNWew006ke/7F2rKDV7wEC1J+QP9QmQeUJcnvu+E39rY2CKGd1RsChvXtasw0YQ
ku2WBJEPiOXvh6zcZuzo8N2HYRav+70iRw2CKMBdlJdPzKO0Zk3oBvMza9hiZCK6
eJLppaFp6nHAijAiQHk8l8J1gt7lTMVd6G87iy0zJEfsJu5ri6kdx0jqD9EKx9IV
Sk1ChYGOssVoLBs0BJ+SW1NGw6hijTA/d9i7eB4ozqGFRWRCnJlr4QtfuHUfFV0F
V5AV96XOejTDhiWD67RYm7kh1HWdPgRaXH+QV0PgBeoOf8iw2dZ+pY0EIJpAlAMF
QA8LfGB913Z/unD1hjbRQ+n2NYEcflh/bQr72iyhq58HzaqkhNvhEY7xpwyviulw
2+nU/y0/wQwAJFuNcG0Mk1fhoPvKF2c3c5lgIvUuNNo3mVUiKugzWIexMTMeJ95w
/JhmdLHFokvxVjlIU6rvGc2XenhLS3yzBm6r/rCyEuSDkvg2UBsStkJxTRx+54bq
59a5ezV0sZHhFARYAK96+JszjV4fiQMVghPXaoc94pXkQIHsx2IkgDQaoSID6HZP
8tfQRwv3ImH0rvMmtDZ/isYCJCDEc7uRS/KosqgkXIBISS4YIldrW/LMzofwOIPj
xgNTinkGmb3Eb9Og8hRLVLK1pAMEhEPq8Lgk4SMtlhnjPdvzVaJ+RVsrhVGpO7UA
RS0wO/0FIVRJrPDKem8APaUdGQGCVos+URAq1JPZB7TL1fvZv8uJnFQ2szYtqGVQ
DeSF0tj/EXMllJ/38hkMmBUN4c3nJTqbGq1oSOVGjGDCKMq2CK2bBs/XsU8C/V5v
nlJnukfHe2YBXpX283w10sHsazhlLFWKssEb6jjrshiwBHVzb7yhrO9DH6JWRO2d
iJI9ZWXLbdEGUCpjXR1O9w==
`protect end_protected