`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10368 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
Z6yALt3nnSw9nTnZfQBUNTnR+I06uKzP8QjuhVpw7LlhOWjoSrezuqVoEH+XZ9n/
mNfxk58Vj/bVHk47c4RMisGBYsnfah2k25kdf6g+MsUhv0m6lAUNhYzhwFpOuk/0
SJ8wXX/7aCYioJvCiA0Wh1RUJatHIKnu4N0hgadtqRVmwG5stx37oUo3vPic8onk
3TB6MIFMUhcIP/IehZjdIskfM6EWUcZgUkBRX+0EIslMG0l73MWtNs1aC8U12idg
70UsGDICL0mPXx62gkynO8oC4OaJ/fuhop9LGZLzlQCMle10GDSqKFHESeugLR44
sIYbWebo9H+y2asxqOO+z2W5QuO2uPw1lInDIuuBno2Od1OO1tzwLCO8UjXZv826
RC6knkFdmt3XO8n63N4CN66LECRFp9TzPyjWz/so0F18A446BF6+nDPjguUcM6Lz
RSrXh8aM6EBBa5DEiU7DvWYAL6EL+WjoI3K88+pv7ev70gnH7KGuyhzA7JHxnpGm
j9y6IS0lZsHKzi8rJjIJlCYn1Qh/0OqP4SsUsLh6lvaeXiQV3gebdhrIS4wRnkfO
2vmfUF9wrswVa6s2lLcxFByeUEB1XG5I5tV0dkSzFbG56T+cjkhjKF8FAz9DEcla
NEH7M3J25tRR/aUj5weRJpuqa4rEMZ4Rgu1K2c61Npnsg904SMdUR59uoOh20okm
AhaYzp6mb0Qte2q3PMQNjISeal/9OUd2HYpZKKhU1Pdi5vgA1Okhi0EcJanA0PlW
cQi6zlDJsO6PgFvJFvbXIHDP/kR4MNe6ebwMwkQXGEjDPeGAi6gUs4AWlApkAlpv
UE57/8iEdmIC5NEtZOURpKR2yJyvQqoA5A65Gg1ZD150mUo2DgvFiucmyxRqSQXa
erjTK72dZhWlPk9eHHRXMQmuaLN/FaREeuAit9Cd8r7LfqIMEaUHOVTfh3V01fD3
3ZHpf6/elF9iXD31NMjDQDIX2ZW5Gmv/lnZwIyBvHOlE24F9jg+KNURsTKmL8qxl
q+/3KEyAd+GtdoMiIlA1BiWhmjmZPHQdaki3vdd7auuM/bAEgKpXeQJwwWMPtvGL
qyNajj1NXbng2d//NR3ZJvrWV4+8fGjxsoXztHEwEKbGLgL9Gcr37Iacm3PMZeNw
BCJe5vjDYG9ys7U4epT++4n0VAGieYSZdg61U6wReQtkWCAv2JkecCG2rx0XyyLW
nTKHjNzp58ZUTHVz7SzasoEqk2feJ4XFDESGQj5HsmsBzWVecrClkwOmBTSlvwK4
dlfp9BfwRZkv0xS/XPTKHLAe+Oa4zN/qwYZlOwCRYzxh0xAFHN2i9Je2LZAQq2lw
NJnRAvTe8vbmGocRKHnv83KLJNf5yKSjCUFcf7IqhyZU1hnT1h63mH4fO0QwywZo
8rPUqPncdjBQEE1xLwws9Ao5iBHc/5+bp7cPqyl27Vc6OmdVv68ew4m16vB4H8BD
URgkeZXE/DNz8NdQIbaApSPfBvOYRmBdRiwDLRzyz6QFwbUIiAxuMq16kZdPgwHe
JkD+VZEfnReyJRY1dDQbh96HQHqjtaYJFsbQ3g85IwIRfDHwb8jnGR/5BKyz8VhT
c8FJkEcwBk1+4kMq7bfWnzRl1oBm6sERiWsLNqC180P0Ol9vYremYWEqTOBAkJsM
2MhsLXRys2dEw2Q9Q9PNwdzPZFtYfZXET4s8h6NUTdjaJ+fhIxIy1H3MtTESXA9/
4u6cVKmfi1YRG32TYRtmHahAte9ApGa4TzCO646QFU+4gBKIbPJen0/V4og09JPC
W1P4gvG0ApnHS4n3dKNz8LJ0DxxENZU2iMZC7SqMVxKApx6UnellkPL9hH79v10N
R7Y9xke29sj7kEBr2ItWIqdZCDtYHjWtfuLzBQLutd6p6/8/cD5gmiD2m2ebIZEY
Be+5hpEUrlOkJysdyGoW3gtBwBhkhhwCi3cPBUB7Z3SXOLDAY+yJ4YHHUVl8UcvJ
O/OX162hbuWFyT6SuLVjPq6Kt8FmXdCM8ohwKKLIECm+vFff6lSlGsOVgylm/MX9
mCd55Eo3TUwj8f8lv3YSTTCx1Q7s+/WfU6SV/11TwYMJKmyjVt0kXOHPckFiMT3m
zAXEiUG8lb9dtVVjtM6lHc/dTLLGtpvRNjoOaqdiwaLnW6lqAYNmm2s3EStSsoMh
d/C1j7iN0QGXpBuPvltelxuznwfYMNZ4h8g8QwM64tSyJO4p3083j/4BTt4O1WHo
2F9ed9BNOb1ib4vhxKFciGjctZx5am7+tW2Z3jbDiUlIhVhLGkXE80buHgAaqk+v
3hGgpFwJomq1QwptzBHpU00LOgNegydsfaHUSY7XCB6OyyOnkgzGxMv1TPTDTv6D
8oLBvmTX1K/jCNKqvsk0WlMwPg1XaV+0R3Eq87uxZivnLNtIBssXRaSIDv5vb29/
RK2RRK1W4DVfVTaSM05KRUtfOgUNOTVNA0IRHQe9RQ3CxQv2aow7R+OYN9+SovFA
Og3QX7sWNdrzj6RoFHE9aNZZgvZJLyZ6XtVDD2mCf/nzIW3Omqy2bs/ZvxdjKSXM
hAAfppKDUtrKwzRdndlFNveluMSsF/j9ijM8fZqLje9phThSPpRfEwsszrtqJLUx
y9v7RVEbWloyHlROzQL1dz0FnmJMuVcZMlOEYGwrl7peB/qunPj6o3i3kNomVH6Z
CzphmyoXljMGqY2WSjDi17Ayq7BVVoB3OaT/kMCU9GojgR+F9gb2/cH/000+mRwS
2PuQnCTegdGmGfUfA6oLdcamzdicmOUNqFY59RQgne3lfTzVIOKctONMuCpbA8GC
fX+9oF1Grj48z6hVztbJ1XYo0xqCzawb0Z9fiJcsnxGQ2hGTbYJY568ESRyRpWX7
d9k2Ise5M3cDBetZUFwklsUwNpt2ML2ri3RzuSUXq1SnfYqgZ0+exA9xtkYeqOLE
/pg0EuCypaiuU9/eTejVw5dthtXcpeRt1903mGSivQQQp4Jqzv0AbrEkFkY8E4C/
f3GoZYUuXLG36w2sJyweUj4fkB7z/HfL3q40nVRZZuuu7ffhWryHA0wIRiBdw4ok
Nc9n67mb9drRcGJ7qQB42/TSQsiii4H5Qii5QavW3/zhgbi4O/H9RZCBBxZktfhG
2Jpirh9I/uECjxVM4CVOD1JhfG/8dJgweaMRL9eJnKSlsMFwWmaXAMxJ03yGWwxf
NNsAWlT4esWp4S62vmshB3xHwDkNSQDG9gJVEMjINnnpNCr5bxHbFlmCoc3SN7l1
BVBNWeSGlTA9ZbzZcToPSHorgQQX14duNL8PTSGzqD2ozq6q036tiOjWy1BLDiB+
2YLeLh1HeVfamBYJCyMJsSHe5WO4CdDcZweCouO381Bo2S/HF9LtceYh0Ha0ut/g
UV0bSjG+rFx+opW7j/KwRqN1GKLeh+zH2OXyN8ZVS4HrfNoYYSxUcaAlalJ6p16c
JsUYn2iq1bdhgH61OgjyG7kviqdwEFF/5jqAgE+76Q8EuffLPazEm0hKBZL3YNzL
LKyIZu9OvNicvpSHJqaBAHb3FVht77F9mYejINVm26yoe3tarFFGy+2t/zOs3NF4
sUwrglX7Os+uDHZl5mUIOTeDkgrYX0fqUOKorvD8w9egP4v16f+5il8AirjfX6Fp
7XvFVZZQZZ9A8KRX4o2sG40MRwMT20RfEmaFKDBHcPxtV1zw+eAT/XgyTNNDgGxr
Fjg3aW6S6WEq/Qp3/r7IwqvgVsyJZxlqy/KO0DOM/4bVUIaX8SQRnalSfamQjYcL
49bgj2DuKRahSj7kwUMvIgQTbLN7mquca7iIkiXkDNNrn1Ui+S9ARFejaNzK6Yrk
ui5vavI0+Sd37w2yqcppIaMA6GNgNX64H46xiHFm6yNyH6NdpsN8Epx2MYIZu17A
vcfLoHqLVy0Zj/YMcLaEloRA2/vvKQ7HDXZbTr0OYlCSJ2KbeP5F3I84UMMUCptb
t1GI+/wu6xWcTM1ZUG3iuczCcGyU3//VdPhSVIIXCl/2vyRInvpyXHfQTAjEUNYc
9djuNLx2KMVnwG6TWt65af93PdmUAFohT9b2OOtQBnE04lERnbxajcxR+9fFjqLe
tafhv0HKetJl3Ae2tDZzKQsASgrlaoV5Sn8XAt6x+jMrIgjj1ZjEK2LgYf3Td1pQ
K8ZXpY5Qzo7vcJuBzdifgJkRIgbVlCJ7a/9XdnWZhsG8gORH9SU/Xnvw10b/vsWw
VDMehv/wkW1OenZ3E0VbT9SFNPSk0V1IN//MvQ8uXvUXmkZA7We/6zWKcSVuW0Iq
bS7RIO+Rv5a3QQQ+8cNfsRZ8dmBOW4plrEI8VPIUQNKIEsoPduI7Ev3/oj9jSm8k
TspjFR9+GxJx5gKrtEBehpXI6MF1gCf+gp3CfmfikSmRFLa07OeYv11ELGL/OHR8
4hZ4seMJ2RP0A56Oq39Xef0Cndf/2bJ40xA+akLN3eAw+YLpwqo2kBjJotu/Afnh
JRv63zmw3OShfXl2nSUR+zvBWNmrdmcsIiBTM++QVfX7nwYzPQcSWMg4hA6S/mBT
c7qbIV/FjhO7tzPiy53tONHaVCXLKkBCA+Z1/agygFDnAyTVuaRzA5wHqwCRhPGY
dV/GzPMY6+160zTCNST4YQA7fwp+UlTX0D7aKlzHSIIs3UtaxiY7q0OKGd+pfpCx
DZ5o8ofyloWhJ8joq97Kyg49N0VeWksIYBrML/igWwhp0druCbgU8mf0i8UPC81I
edHQZW4/aHA8AX3WPu7wfW3PiLVJPZX8EFiWhLvkEkaMHKEggMJk4ocYYsd1OCXN
5YbMxzFek77X610h9yM8etZ5b/pKyA0ABG5YGxWy2633RVpuDyKXMeptGMJVkmWX
TudopQ6NtrT9Kv9/eHHkfloFwknwHGPlkkKWhVTS29RUaRn69OV3vCqW0GGQlkhM
+UJLKHxbJkARb+fR5+2EqY5KUsF9Jcoko8Rt/XtKEK8nZzYxGaFBvcjmBQl/jvzT
z7EkOWoC/TnB0fkBLmfeAMlAeonYeW8fxRmWaEei/SJb5ihV2+CIpWh3EWrInLVG
IYWGqz382BcE1IiqN4+PtIqErqUho97vH+V3mTpdewEgxqrccArPuH5LVg9/A6vW
6u/NnAziL2JmUBXVCJAYW2kz4ADGJK5YJVVZRqMdVp8s8wAv/B+iKlzPP92w6IlR
5kaU/ByOdj5yW1qEB/CLYElGXB0V2F4Gmuqnpwd2zNntDo6l/ul01VFKaxz7PBsD
EIOCzAEQoZxIWIk8+tMMqTgqdf1LqlbZFoUmbKPU+ZS1rLWiZGlSqUiI29wNxH61
CNO0pkmbsrydDJyWzPq3XzEjSVRuv03YtbPF3ptEdYHysCQp6jLocBnNTxHxA9X0
wS7XHApaF+aj5Dnx46zdtrUlMesk734u8ji136aroMb/0VF5VV+SDIhhHL1diYG4
Vb3gGzyE1cYekmzy2K81N52/0A6zogNvbTitkYFYpIK0LGDsPnh3Ejb8JimOyMw4
BgWeGg9VuOKZR+G5NdGfwFyDy8tABFJhE8XIBxrKI3xKvTpPflFcv6IbLNaGUSaV
cZ8qUzqDFZx9CWK4YQqY7y5HwnJhyRxMS2ZOUQrLtXNmrInXjk8xAOUUdb97i4/0
a6ZFTIrpvJbyIYC4DFGV3yTmfiSU9D9W6to587gsZRGcY/Sx0Gm47klm7u1pzg41
l0YnbEPfJiA/jm7TKXTgLa19Ilt4PGNYvzG+gFtmkkFOR5chMvrrb9LlKB0FM0Bl
9rRi1/z9I+IYEsCvm5BrWNmb9D9ivVnQjJWvZBHrvD3LPxOkr5lLlSyXydav4NlE
Ub5YUvAjDTvviGSEWODPq6liIr9lTXFK5DlGHbagaKl83FqcJkkXZ2TnBuRDvlGP
g09mKGbbORR+ivcPeFtevqlHMMEZjgo2J/0EDF+wO8599QqsY4m6WzGcgHQfDh+r
U7DRChjHRgzNRpF7Lx7scn54j0zNbzGZxVddUqhW24a1BPnTv4XNJJo61+vwpCKc
sE12IhAVUxYhfp20AP7wTLy37Y8ArnvtPAjjmS7M1bo+FX9EEmfCsdC2UgW1K/ji
yj4/87slWm4LpaTAyRIlPI0PAy7XOlkVUoW+X7We0HM4oHPE5BSelF+BoRptPLyG
ngmakFC58ZHBZIirAgpdJJvb8Z6ACaADh0fZYhsjtUWiuXgHCtHbFw0zekDc2Vjk
cnAWAWT45a5OxXBQYMH71tJ7gtbVo9NjkuyjPTJOU9ccXCXITOtfs8H2/6aDyOwj
O3QtTcvFjYE2iWkOsJHdz69nDvR8P4e8762kyvLOy3eohjDTUX7BQBT/v3OZXRjl
APsIty4ayGVhbPVkBoDtegFeH/iS//dsmWMlOXCo6ATKt0ybhpo5KdVPlvpchJgI
e+qkexVkueQ+An71gqAljWnRIRl0463YxYGNC9ywlerPzrBf/89a3akSXk+MJok4
v5yjjD2kPGnTyGNBf1tTHTV3vJ2vSy9GbJqqwU9LaRiUjJxnUg/S1rkRa/3+Crzc
kJV6Pcd+686gHtuA6/r8vZ9eDNiX0ivlRtQfx7F90NulF+ewUijVtQJfzsLNHBQp
VrupbI9lI5tUm9LZRiSjv2TI6Dw1+UFT9IYncYb5uz0OY67xGJfZ+Kp+rSn8bcQI
YIOOi/qGCLRWTkn11uutkwAWWioyzmUJ3pnDgIePVSbFTtevqYtyDbfTEZyUA0Ce
p6ai0hbdmCfihOnbhIPZwgHR9XQXvjcWnLycurvPkwUJyCRe/nP/EA+xKy17wTu0
sSkCCXHgZdfheufm7ZOsGMwEZ/6ntgRh2MmtlzmzS4quN7fVe6gQp725orVGkIBe
P+59hN6l7+diXj5Nop+kPaw1MZvdDzBsilIyF3eqN2hYaM6OP3QdefhyFvSbxe3E
0+DDlVdOlEs89Q9P1Xg77cvWOE+SYZwnpzSksTnAu1Mh9TedKJpv08ijQ1jSn0Td
Nztx/xU9WrAIRrk2WZHEIL+Zl+0muBuRE4H0SdpM9o34+8kNK+hs5gdub47xf5vS
2muxexSRq6Z7zYLiaUIfYPeopiianyg0AP6QXOH8QIeuYoj9QRvZjHFVLMALzxu2
mGivczmpZTbkuUo7QQJ26QlBi9eSP4iWKGP/WJMUq5li8UpF/+twpffFNMisuOIP
ltl0E0PwEGvN2RKWahRQhcL8h/nyCnLvZjtQugd4csYGBieeESotSpU6u/wjKqUz
Y8KHaNMlZqTmNBJqE/p+x+LBaqtV7mg4x3c75cjPjI/CjyjaRAiwpcG8ciyibu0A
wydAyapfSrGpvN3L+hhYQyTulDw+WWYlntvJqCh1Wkla5OqJcEg0kuhor18NVHbG
//A3N7ogc11swfmKuFpjqLMETbRMFGrVbF8CZT2jFPGl9HDbWXf4DkJSC4Kdw+c2
jitCiEVPrrPJG8FN8IjytXpnVH1dclEdLEuqiCanePXkbYqI45b46bOfSE6Rml0y
DOwxzPURJ03FeEYEI/Ob4maPdnhn5uvRNyQizEFC6ehM8SRe8BW0yFcf3X9r2z+u
sjl/jhM/rMAkpNLbVgBySqsZpqdbX3VEimFxGBPgyzQHucHDlovR+ATa6Nf667GV
ZA3D/FVfNnLjSTqZ6HsOm+0GhZSOuQatQglbAKKccLyTFFfURBJgmSx5XvVHOjg7
oTbF1oW7XpbodNZ85jsEND2Kat6tsMsAJOZf0CpWmKzG5AHJ38A+Wm30lurTgk+3
EwlgKLxQqGs/dSa2gqis10TepvTqdHNf3vm9HenhqVHbw8k/OKbGQiM3owhQXfvo
isxdm7wO6MxtL7htlWkpuCaOipOY50Sd1Q3s0wOH6BLjtFq7buJPK4Yl9jFdbjuV
wtJfq6jOcIeUbKslsDT9xQMPEPvfDJUFERdfXCCdG0mNTxBsOivWgjn6PdVd0TTk
IJ8y8t1C4LVm+NP8pI8s/Koqo4J/Gmo+U4xQpFYYQT56sNkEX+CvK89HtIKBhnwi
x5q87Kx6Hwl82sCCw9UgDGjR69QyqBrGPGCa2YJWKWbFd72eGmTfxI4XQhfPuGDx
WvOTfDzimLkY9hBkNAGr8F65iyuiqurbDcR6ND2CL6QhE4WTbAysziDfN7xob/qG
xEMr8f/9x/88695IQ2Myxes3wesLoeof4JHnnjTzeR93C+rYoDZ/Oay6+ukMeyKR
hhtgggpbTNiiXF1CQa7mVwsLSQaNzK9v1p2BP0tkBhiNFB0xgT5KfyUZi+Jl4VvM
33BZxJCS9lqeUCaYGeSJLjpmvIOFWxft6ZoOvUzJoukCaQnDqSRZn0i5udQPrc48
lOHurhiOLxRj0mNz3u/y1/LodUCgS5ryTepJPkShblw+dxyTYq19AFzK+UmKN/m9
O5q1g2xOC7GKpKrZt7yPEG/OjwppmY+09OsEA0pUZEaWDYlBBXP/q8ePcCF/ntMq
3B4Hv7RTN0CBVBrim8Vbr40pkPD01bE8WQsORybxq0YNhy+VG3uxYwW9DkmIFvUP
JTgdAGydDJcm/o8RTbcLQoxiIfKTwn/tDussD6QnmPp531MJT57uqL2eh+5CcsGs
HL/5/uXklk9jkJh0We/MsukzTssZ4vRoJFUWw5GPMM16lK1l+i80zX09XLzUs0ia
NpIwfeF/WLJWAQEcI36U/D7wDe7DSZl0qdp3pkYdoEoEbT5uOHVVAc9iAv0eGTnk
+YUSj1cD+LG1KJ3qFR+2VYxCOxaCaWj5/O806dMG8qssjEjvEeBiK9X+dSJMxgav
EHiYORHCQl/7d4cU/aBsnluOEas5ZgJkFuJuvlCnODLVK37YtKGrmQVDR/VbX53I
2qkmt1AOLPxZ1YfeslRp8ay+uWqjqjvIRSEMNoi4su3qwbT8JoEzLoQisKho/JDx
o/fkwqqat9L7WWHjprnpNqrj0qbKUd5E4l+PbpcpGN6BQPi+8cEvU3ma33RcJYFP
RTenk0nuU7Gvps+KZFkI1eQd1t/7mdpkjpFdfnB6OwiOAfvoPrFMqNR28KP2sB9p
yNwQ+B1XWoiK0Pb2vbaEgtesr2ArTlqibqa+4Huav0giJQSyuGoKK1SuCJAtIJkz
4aVVmgX7EshSLe5x29gB5PQBXrIrISYK7XHrdTXIifR1OejE4tpArnNsmvjVtizo
K6zXpR6LU6+K412c96uq68ThH4mvKKJ+5MCaIxrijU8HXlHLWczsMIxz8EsJrkjc
VNLGdMMadQjloaZR/QlxiQjnROozGLTAdA2daXAZqtNQr4GcCzmYxo7J0HzQ3v51
ZKWNl9RyVek4DcV5kh4bf1AaaBq0zkiQ+ng6htkKgRk1X6yHV+ErVTGnU/l2Y6bp
kQIgbBjMxL5mjoUxcDakme+2IYTvATQHe2WvJlnhhin7hDZnWZGE8SDpOhQ4yHGL
S+hClB8q2AUMoX5vzw2u3CZwJEMHZcef4C63HQruTbwJQy8FpAkOD7bX0uJQD61e
mRujVhjfLqwcF72skhLIBR0TM4eHkAeQLvsSFk8Hv55cP0IK7kv3gJGISfu6n8ZG
nb6Gr0TqB9WzWOoe6dLXMx24jiZqKgnbID0ySlL61x6JZT0IOoDT05qX0UbFihhN
nORSmoPHSWqb5kChWMM1/iufftgF3b69E6xw3oWThOOlPUpdQcCTn+abIqukYGlk
2vMbi+f7NuPgfR8zDzyIqBWvLBPaQr5HBBbAyZpRCa+Z27DhJFeDbaKvrDI2Gc+A
UXQQM7Slw8teshqougWf1XzT9if408GCHnHgAhHAd0uLX1145ANTz82wQmJiK5fD
z1xXw7DgOMM4NduquSVxI7r0BS7TDky9Nj5DpDjehEGxOUZgyI8+4sezCFcX3VZb
3uMsiMpmsM/rgv4XFo9ivzw+kmMZbHylo0ujnjGjnn8pdmkGnhwACtU9uskhLUF7
c4zOaYThELCwwTCPm92FRMYfuSfRBBq4cgFbZ7p8NmfkCPvzdq/0HVzaMipJawCw
oQTdhl3LaBz7PTCqWIPgGMz0FZkSgIqbORNrllRHmfxOSBLqIrEpLrZwfrrAomSv
fHAI9mYA+LB8l/A96eBJxJUxfiB+/6ruvQMqn20l2f1w2zIvlDT62rFTbZwuZV/u
veKkpWBKGtZJIka5zIr37C4S8n98G+TLVibdYN4taNVJs17+EcYRwjvbKbbHD1NR
Ek+GR1Jr1YaYXySC9b2lsxthfSBmy1QR6Wvd1l3p2zY2MXZoGFPOuxXFKBdSFWUK
7JZsrZx4D6RMFDJr9sI8bkTtDzQD04yGSGZ3CcanqoXKOrw8ys0fiEwhtIhnQaCo
lTTC9l7yF5BYVkbeAZEA8y4wR8v+nZjOY5aAiDnzPWmnln2p9fq5LRNEueklaT/s
mv3jYs3d651T7O1Vu+UwNzPX+9xq7p0cw5bEr5a0yv/FrDrTkEo6nondyw996B1y
dMa0W2qouwO6E1AjE+ognEDJyRGt+QQB4P2IkhKPuuny9oHocMdu9/GWL8XZe+L7
4sGYVbpM7GG3QRCyGwGWltSCvbchrKC0btAIpBUdjA//SezIllD40y6CI6Wxdsxk
C1DKoVSufnhoExVZED78mWmY5ltyq4mMrSTbKJi3aZMnZ77YMU/H2RNoSfnrbjq+
ObA+tNZlGFo6Foqnzs9sNPQo5SDRvNzKmYpVh7kfxm0J8Xy9qvMUc59GknFkd6Em
wVXAlTlVR5jGBVRte7jggLOCFPkpXFKYmR3fShO5cUIgIvpjDD0BlDYKLb87oKmV
g1aMwOLxwdMo96BC4SngGCMsOCwKAvQaoQCmeX3gltbxGra0S6UMHk2rlfzsZ3yt
zhm6r6dBxqJ8jZa6GCwBTupYuOGQMVPxE7N1ivQf6Cs/aHOmWOg52wXEZi1RGiLu
6O8KELTaePdT3o47hy9ynDffYbz1EANVSyP1iOZLPz3xZ8LmEOi8K3nKsV4ggY1j
3uwDhYc6hNwMzMjaedb/OqAMwA+Xq6oA2J7evL5TM9tLbGL8W1dxswC001SYEiWO
68+kszz6pqQLOh6r/2jGeCVzX9C8f1QjyLtZKUgWfUUW10Hu+e3dqywdjILsC9S5
dY1g+5SguPTLKueDK/fUk1qhoTkga+QbjPqiLzhJfRhFlaGDNlaDFEDghc88aprz
SEgnF/inNq9qPNSKL/hQbk2Cgi2YIjNGEgoeB1F4tJPANhHI8YMy0EVQFIpDDDo7
PSjbfzd6Hg4idjKd8LWjCoJU8JVDw595Zb2pZ4rWPVceuVA/ac8ONKR0hRwr3A7A
kO8D9nXxehLyYlsU4P00GwD+dw5NbNiJ73yzKOQ/r/pURNPe75gCb9aMpnyZkgH3
zfcPDey42ihI16nW7s9VOIsLM4kGKQhmNttaAwgBSJDr9VyBN3qaNX8bQu9zAedc
+eDJazMWEk6mFVvoTA/kqlhUNtF2gug4lGOeIrWtKY/unbVdYW+ukfSb089HT66k
6JyyDP1AWzjvgqIkujeUAUNq8wQZn2cfYzrWrGHuSB+4uCJketTjpnRw3OL0isZa
74stTjnFj8GSYC2QeVBBBW2v3omjlCIwTG7fkP9svOxtWWrmXXC6DgGGvh1Op2gM
kYtvL4ac7m6pE1rYUWRl75f9hJKKKsGiEwSAlOW9tIhrq1wtLLr4n8zUMABjpMDY
9ZgVsgPKfFcxu5W+EA+NHwaErI7BWa6k++92wDDdb0zdtv4ereweffJEXi0L7fcW
BvVvpnLNw5By1EYUEEvX/ze/rMza7yAGPov7WR6h77IyAUksnhDyj+1R1xlcq6Wz
PRTk9Aqsvx+CarJzhFA4c1V4BeXtd407aqaONsqHLyrwRcDvewI5GlTGoqMF0TQv
5QupqrGoEpQIDHzbxuDe7oqCKwxv9l5cZv/TB3lZf9msEUQMvl9DqjNtoTgcqflB
Vo/pDq0Q9KkaRfb4scBskEFQjLacGYFLlO8NxEpO5iCWJMkMQbGZQsPJXxFLEJNb
FtSo/bqdipL1Uvsc989gkn0uITPlfmJTpQ+Nq+IqpMhH2OzQG34EYh+HrbXcRbnp
DSXSoQhn/rmTyacjH5OCXgPtBL9d3AhY8Nsspz8JLbmji3XR0YQMbGJeP1TW8vN3
ImcXmZPbAUJibcJSBUwSZxI5BV8NsRTwspfd2piCofk9VmFR6o6ztfqRqDTjU6oF
dtHfz+uzRJaILk8qmcHeEgV41gdBjuyUXASzafJlYzDjijE7CVB4PAbDeu0ea6qt
9khO9w+qhBgD5A5D2xaCim4bUcet9X12Nm0bwJkBCYRHjp8UumpX+hMobeGRaRPF
fxqUio0G0kPEbUuOef4FIbq6MUaEI/ZRtcdVMCUohHqQTkzTgNe7UlZC4KQxfavt
wMEKG7JlsHfbkdetAy2VmvU7ou9ezO7KZIK+IJJMfY6KPIdbQQNHpppoQPstXCe6
hdRCpmr27rwqJI06g+xLiOpTI0GJ8xHMDcufidnnvI5IQ8Pt4tpZ1FYsF3uAQRuQ
vtnR4w8M7bcGXpFKBnoE1kRfy0O15vLpnJBZU//E5fwTrmUQBzFhYQKZHQtZ+Qq7
R/hhNL/z0vvX0PVAcZDd4oIHSdSffa/W+w2nHxh8wR5QA6SbtRrMoqW8asC0kdFA
Ymxz6rTotNK+mTiH2UcBhsPeXyeadLCmJLTKlHV+wmild4MAQKys56BjoSiTbs6c
eTiZxD1Q2EcfWwnF84+hmMzDISiBT2MS5jg9hxSoELEzLACAjXDRxjD3nA0Tv4Gf
ecViUpXfD0ATsAyL8JJuNJqFhd7liHkeKFPzEUjdb72ccaCmOpcKXkideaPiSVX5
DbiLwjE+COoFa3noSr/OK/TMx80akITSda+87ecXQWfh/m3Re6YD0J6rEuSXeDCG
QwL7VUCMOL/VrOU3p46TwhfsiSa7OU2DtakfE3qHUGQ9THXzsImdJavIGE9nj0CA
IBGGVyX7kdn8yvsLHNn/zeqapdAllrUXxsgKAcvNNH5kh4ws20sBoHhpir+IEfO1
lLk8k+8g2NUdTSovyL5QVDbS6LCQcK5mfsDR+Yojug8L5Q3C1Ip0vV4tBFkBWJ4o
7sCHfh3/3PjWauhelyGEdwt87zm0QzEw9KKWn+0Nn1Eq1B3d7IUP1YP3bNz7k/6A
bplhTEO/8Q8/QP8pgd5CEwS5eRVJHwGEsaT78U4calMiNM1F58jfKh6CJihoDJPg
rK55LzRsYYUkmW+6sN4Aaeu/Ap486lW9o2Lph8uGxsLPDR6j7OHUpHYaiPClc8kP
t8FZxyrvJA1OPFIUf0h/U2SJlfAk8DrxywydkzTZhyx6IDjamOXX47dZYyeJdcs4
WkAYRtJev+CX1FUcszhZx0DdyhP9MlWKWVdB6v9vXeLllFQyJLDv7YO3665Pz1OA
GXbuiuRu+NBpevyNtk+siyhShljCkVQPrHMj6pwTQhl7LjjP0aA0kfUfNitVhXJo
6lbPGKtof93ZW5kOWOBOEjBaDdynv5mzx99KRnglFqjWe0MEqKxwfDE+vDMRw9XG
oaikIUZC/PiW9f35uFNSlt91xCKvE25Iu45T9sV4fqmd7tSa5czkS4w3jPenVtCM
kZJIW80pNHWme/wOru0Fy7s3fg7Fg1QN/d0eYh9Ax48Snjo6upefvIPMZVwiGrT7
E88HYQRppnSidVsx7HwHPkG7tAJYekJVqjibsVA7oMYAjJxo2r7F0Q9Z7vB0l8XF
`protect end_protected