`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4128 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
qdq7wRaiR9k2mYjxjSYnpyexiOQyecCnxuKl5BCBbm6qmGcm4x0L25b0Rjhjs0Jn
VIHwnQu5N8AlHWAvrqFXo87WcExzmZSqDjQWmVORLtlIY80L8jSj5FLwu4KLHATk
9U7IAHCHb3cypV9OIYDyIiIkT6rkftjJs7dCF50x6nY43yew8BqUyhu2A7cfJeSV
R8ZVtcBa1ey8pp1R/W5BxA8tpaHf72ab0aD0Az7AEUQ5kizKOD2NKW7SgUqfe3eo
5uMXVuwudbhN4eSNlO2oCLlNI4ESpaj2j/9lSeEZeOikErZxfkxRFXofoKSltDTS
CAvtOuYQA77G5qnl0F3sejoTMQyFivh2I3WJOLr4hic0/lM8EAQu6qQ38L+lZbmR
AjzMfe5WL9MPPo0bcTzcQROP7W01LEsVav86ASS1/Ocnrcze1cYeRHRTECbrxU0F
+uxno90HEETai1r5DKpYHqq+gsF+CEvNY5DNTbNrrxLnu+6uMoVDngGoTtQYwpe8
UMapHBnNBakPs+CYZ77Bc8UUOqRVhc9x/ZPIqQnYpwihflVbRWd+suARFojVIljN
zTcdsqK5XTzM1kr/1lQMsTik92hbtJCAO6oth/iLnoAzSM64cTlbUkTpVijcsnoD
cK0E/QaTZnLf5bs0RAYmMTdjhFI+ksAFiNvTg18LEKZXQhOgodqDimFg/g8+iuH1
TiBA0f3+hg/6vyRQyvpAmUIlTgJSfBOTEOUDbNGJTLl+8AQl2Tu1BWsPkOrgRCwq
5uWzJY1G4SNDj+fAXzwbUXkVeXg4TqTtAVurTWQKY0iRXqq52kGN1Asi3CzvWFOo
DpXvU8Tc5UUM7UVmwsbbuyFYlHGRFg4Dr5crX7rK7zrHfCBX7XnnkJE1OrbxFPrQ
+LKmp25LFuGMhioB9e/XILtTjIw4acl/McCQIP3sCQkWwaAQa09HF5CoKLtjVOQK
CD6G4Kv/tcD9N7enxa0bEgLyND1Y9NN/1rrlyZyRsqP4lKrVVyBm6tG4sMmRDSup
NHU1usP+vWbbXZK49nwaOxDIGMY1lXbeDXUBp41VFgadAkhXibAPMCRI1ZmDG7um
itCeb+mrvCAHm/fEIpUSNeonDQFbfIxQA1vuUVzeq6splvXw7NulZ7j1DvNFHTiI
/efT4ezyBjYeREsum5ijdQ/PIb6sO0Sh7Jc3ouG5XXjuSOqvKbAsgaQQMPutSn7B
5WF6sDjysNt9TjHEe/07RafqVcrjqzBkAdwB67Z/Px6McPXUJ7fiwK+q6TBtL1U9
kU9bRMmzunEJpSUB0IQSIr90Pd937IwIUAjYRdrCEXE1su+JeXQw3M77CdMuTxcF
inPh2eitCV6ONaSok2EaEufqtimMjGs2Fv9vG8GpSlxwogpLViGJfoc8tzNUIsgI
9vlReyGgGfvC5aXoryCc0UE9uMBXfCd22QJlqvoWn0K2sMx6XBSxDezwTKWGt5sh
t4Rom4Pc37ub0mKa+z1lLaQDX65pgLhCFydQz+WAraGTP7ewOFYxnj9WVoRUJQeW
vMOlQuqbVDaQFv9ZyVnKpPS7B6AbJwtwVPKtbpQ9zQo1hXvZHvGjtxVD3LOskAzU
+nEYB/WxGoJ6noquqbgKz+FAF/TPZ6yybfavvIWJqC53PhyBbSJqt7rEYjPjXmeM
E2dxjCjiLgPMFgJPXrqiXPZ0qC09uHPeMraQPEYailD8hT2mKUHyOJwNDpKr8VTs
NwTCJYIE1c7J9+MOcL1nMYlZJhcNe1dxn1Kw+SImfLvXyXDkdopZCeLYggmNX/uz
JroXI7wSxjrqo+SPDOB1BUydJqDrMBYlixfz7DsyT9y6fmqVQZxJRwlnG5zvr8kH
qWoYrbmP8olysOxxWmv6OCFvkfT0Vl7+ixfsmPM11PwsCN5CiCBoLtcNKbL6yE4V
A4S7vU4qZuNxbUMXHnFxCJ5eNkGnrDrEmQJRz4WuSWsXkQk4Ozygd1kArAQiZ/sV
qhj0rzxzCDWt1fgF+tR5DJOHf8r4WNgpZVst9v1qCKPZ2VVGRc+wf4Sasjz8lAdS
6j1p6MbM1ad52fdVlRpZdelMtf1bOrnzt9SKoZuNmuuyMwdrANvLPQoF+Q3npVcb
OLXAZZ3nmAJWu7VRMOKiKOcrdMNYnYuIuScPdy4YRnQ4CZmsqE91I7EA33r4tHt8
ty9nbDST9BVDjbTztI51GyzJ4CxOKHq+Hhe88DRJpwpbJKW0Pi9Z8a1dErFr8ERZ
5CeEY2P4DHlDYSuG9vFQ1GZ5tqJZxwttRnScUfUtmcrVXFU+NTHQVlmNT2zfP3Uj
+AP4rIi4zfoquNxiQ77PF1+URIjgPy0qu1JU6Pz07is2o1Gzlyk3k4ob6xxe15F1
cXaPXY3EwRVh1rX8zWItErwxhnXf1vE/r5fc3ieUMiCMt6vJRbg3P7LrL/JCkjsj
V3YEubiexSgkUs7dvMCmrJ6m58Egxg9zQdMhvifnpkz+ee3EU1Oa53SEFTfN7wGP
7mxG0bZcvuvU8S/KF0/c5C3GstFKZHHXGBqy7tOrf+J9EkQec1blaDzetWR+YpD3
rewQUPKBJ4Gp6E23bGw8zMjpJvELB738JYHjfTP4VsPygkZ5o5q+J8WS5QZSNIIC
Lq5mEDw4BVaG7pJPkFbpJDtNM/MATzCxzzs27n8DSEtaXeAz9OGosB6NZhgh05DO
1NWsv6Zu4c00EYqSV+bhO0z94sEtGm+ifNvjXcrvKnLaWKv49nitvwMEXH7grLlo
fMOMBaEJEQG0BCk4OesEitClaNV2awgauTygqw+F49XShAAWsMoCgKMZxYCigGPq
C+TqlM7Ib/RN2yYZyQYANdrFMdboCSYMK7bVxansy0Dg0OTwvFP/Dd3ZBFthbQKc
gYuclTh0VgrPv9OdvK/yMnrvupY3zqB9BdUf7UbiI8VE45INiASpo9IyhURiRkti
RYFwPpQ62Gd2/jCd9Pg7l+jLMzLMLpFzaxDmtnF8UM9AFMIw0R49FzRt7GtHHVRU
MXyOObgZl7/PiMgCdKQNwgjjCWejmvf36ffikQHOPVTqraXkw2RYN2Ww8z2h+Eyz
laxflhVAxQHJ0FqBTcLZhHwdhEL/9MBz/XBnvoJPv+BkfG0DhOMFCrn0bYQWLzu1
Jn1nq6oKJ7Tf9dP6IjGkx/fzzSp8l9w4bDaLxGCR9UeFM4rg1TFygV9GenDXHE9I
BkFi91sefo6kihs5OZcFCpFAzbblKHvu9v60Mb4JAKdLXsfRskKnNd98HfdiwKoe
99oDXWMitE7nKOSeFjjCNXF1yc4X4MAMjMKCbaBlCuSUvxirf1b3m09Q7GqLJrpm
hBcKoEvajJYq7esv/Pij+OFuahdxa53EF0iOh5FwEptlP7pciK6DhuqeEL8hRe34
ZgvJu4C+PHmKsizonCi8gOeOQHGefn28WJW3Ip3aUux+h/4SSBpH0gHKYEJzucDs
bfmDMPgNjDpvd2b7Tpu0gtuABmBq7KO2IY8MHWBBq7Z773K1uXKmHwY8L7yZUior
XM4sZGO8XNfZ7JwdkstmybN8aPW2/476z6DRBzo7Ro5aaiVGjNd3OCUrcs23x5sU
kyQWbi1WnCLlpoZA5Da2GfFCppFhEwbGoHSHBdywAPyYRr3HVvNvjNctjFNPP3Dc
XcvKKh7CBOG9t+iiCRjTENcvn5Fpm27Vv2V6c6I/kLjVExBi/OmPjWIfGi1V0bSJ
2mNGzzxXj9xC6kCSOU9Otq7IVj9ONQ4oHg6Kv3p8D9h46neOVfs+0aRP8Et98qby
ztO90zGuDhYZ7IeBuNtmHOl4O62mLH36ybWEGWUL9PSCbInqFx2Uib7v29Hpxwk7
/i9On4hR5ql+zHzlkO+2EdryKi+RUYXMrnYMk+u0U56DsvCAyXGXpcPva1V2hNCn
z49qVtQfKzyY6b8SagSQHLI7P3KZRbPqTmqhcgcmcsvKTHdycfNCGx1HOKIVemNt
DTvmGiTiF9lDORGZTgweSq5StX2QI4DpjKtj8whx8gzTh8/rXO+ju0r706IauIVC
Dd+HyxWTyuSb/qr9ZIjb4fVbAfDVm5g7av6StevNYcPNnpRYROjYITprqFd+edoL
yprBLFE0zn0gP7QxQzIf/U7/VTMcfq3i4hq8ABBM9CevCTMDw3uQATR0cxXa95Gn
wAYeNXkwmpVv0Vdc5Wr/YlXHljmWCCZSNvzkUXgawnvdTNRTsJNkm/aJTj3K1SxK
Lu2hamP8IQXHB3370lXk+BfnkRuBKNvICMF12qzwX2VtgwGhO8hqZnQDF/IRXElx
w53NjjL7bOXM7ORf880WMfDgD0w/9Rkg976dx+sMgTKZOJWG8Pup/SD/608tgBeW
PIzXJvRNlIl+w9HHBUEIeIdWYXHZ6u1eTP/6OoDSsuQmjYRWv80uWGJ10HoGeda7
blPv1xJdBOY/Z34FS/Ty3votauYypAGyKTGnM68uP1CWwwaMzLBKvqvDxJvPuDqC
N/QfOKwkZsc0cg6la9PSbnpjcaw1NHC98T1Ct4398N9CWQQpozfZ3wDLP0sfdPTr
Gfh52pmGQulcisC2LgbbAROxupQDXaPDT7aevdWtjE7bkRY7WNndno8TzU5n+WQb
zt3aKG1EsJvmq+CKyDOx81a4XTSoCKRoPn1EliPW6IjY6v8V/K/+hJx2OcffCNgI
747aE8BtpTrvGA3KcSMniZXJxOQXI2gXveoDND73ILr30Asvl7OBcuGxsZWJXl5z
inBecB5btKJciy1kErZiJuf3INZnjGXfc7YDEarBtH1Eeio3ggQjEJDCbuwb6yxj
vVjz8mVyDMtdYAjgX5GFL1rf1UAwjrZ1LQgUM88k3AabyNynfnqHwBZ1GQGDSZ/o
DENqJo/Fs5O8+Yeb2cOShTQ/Z2WgyeLJ3iC25J4Jah50gkptlOVnEcooMhpgwtWW
sQXUATaFKOlFPAVZxUAb5NX0CusoUjL7ul72iPrqxH3AoNLYSerU8KrO34x4JK46
b+XYAIKzVYWDijJA7EgJ0UswGi/nWkkPG+jFE0evldt0WvN1tAoMilQQNBpc53B0
YC2UiHpwArqJ4gnWgS66eN+HubuMlZc0xe8zQAQRVkE1pB9aLe6ahjRwimCeAOJt
yRoKnkrvt26mAreFoT5lGyTzewI0vsAiRs725KN6su3Ss2Qp/qRKW4du1e8wnAFt
UUZNzjxsWSiq7P5/5ZpR5c+3MJoFxLlxNfF88oCElYOXGh4gRgBhVDklgBQFNYv6
1HoDTF0Z6VJF0eG6CgXvgtEIAptsjvyI8sfLndFP39G8ZL+powq4I/iOeDXhQv5y
kkQRDfkP/qtzSmK78fXfMmFl/gYnuebVCCf/BoWbz1sN/cSPhsdkPc4Jlk1sayqx
`protect end_protected