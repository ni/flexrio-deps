`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8672 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
VKWNRQF+vfUNEEp7apOJOYgs1Rrm24OlWOC+vFutdsklM+YBl5WhuAV6ZvuwLlUO
nGqob4+r/9jp4EDhUouAmLmi/F38Au6YTV4A0/Cr/PjaCK+BWv7i5kbUlOxAKIJO
QnCJ3Gy+9WUQrXwQS3uR50dzdFlY3QZVm0D+3BBIslX4HrRMUuha7+dTmJdYlFPG
sUtBUMpl1icrGuucyh5TD/Rjt7lSWBaut/C5LvLFt4ubbeCZk1sITl9I38WqknTe
rY5LPZJJBX6RIsDfa7ctV09WFKewNuPP+EivinDJ35ddZnIpLAkAHngTRN62kSQW
ULVD8vgWNAVR/XjkE037mECXkm4yFdys+W+sL5r5kiT6ZyHG1hv5d9JtZDT4KJnH
pwQUHINfMQ7iEx8A2qT0DrsuQTohgLW9eESI1j7ETZs+hsNeZFUzGO+f43V3JnNx
63LNbgn2ZzA43LsuIJ1hnm9gTt2X4KjB3TCXR46mtSchjq/3lEVivJx7agb2YnaT
4DbP+CBgAVHkFFNkxF139MDwV5OsXbyh2/DzaC+VQzV6QRXH/U3QFIMuxESMAN9w
U1lZhZhZOF4f4au7L0rq9kXijHwu+ksMkIR3XZtBQaC4iLW922OMuYvlmri40+va
I5UKYeoz9ffcFLcoPUQs4M2sVBlXgiX9UFAAHFT+UlvPf8MR8QMOecMoFiVjXHDj
zKnwMzw15HYQ3lHSMkVzt/7OLBBIGijP1mvEACKi7JBgFlnEMNruLSC/1dWo3JhN
41fSqIX3mqL6WjRTFSyAl2yLNt1PyrEUk6fC07+sS0/hYxyeE8lCWOkO4F6khjS6
GQ7epeGnB1NWAAHSJRo43KH+IDfoS/MeRAQKlwhMGFC2MyoNiANzpJF1e3a3XFAV
RDSx+Ok1IddUzD+RKcAyOA5u457zjXl3cVY57hBVwTLc14NdlPVqVsX7phgbfi+D
qQdmlAuarNhJ8t4dvnAGod6vH2XTPHmc5X/c4wlkup70qXEeT0nu02PusMH355HA
kTFvB76INd8C27/0LB1s2sZ2A3x4v8RyEcae9RgBtoAXjLaFRIVBZIfgtzj7bt/U
QOx+wgZiiiaKJRE5XMYHSjD40O+/tTZZwfirOWoH+BeopRq4NS1iCtGhiMi4OnoM
/i6JCbkr9Kr214OGgNaC0dd6PlviqkhRydPCJCDTUoDBU1Vdg/qt553zMOYzpTmz
ojmc9nlQYmBKe0bdJW5vjJzTGlrooDPcl+u7cK1/wy+XaILyJ+XDCKXToh4N8Jk6
cxSSfXhNe6slyZy1Znrhb91zrbjMn1yp3Z/jdzwGFd65IcsHJwkjJL9nbyCSYQLZ
d56sSc6B2HP8nmALben8Gwo6vXODqj+zv20rjQF47gcYTiyZQl/NHvnScHWPkho9
QAId8p7siyTFA5LdVVuiivk6BK0m2qFdhSQA8uM+L9pKwYjDhWRWNGyu6lldDIno
zUB8xE5NqEaOyRGsbMX1yWrjMZnwkgJxLD3HcluG+WS4AB8O5snSzORqhPxPGJcz
Q1OOZ+4EkVZISL7X0hToGq6Vp47o1fUlwqnCWft8MhjYZlpbC2OKQVz6gpht9s9l
bYvKUgcoBMKfK8YNa6p5yJymUz5Dfq5sNy9L9COcF5DCPkc9yi61c6epRXwJ0FwW
c3Sl+B1R9HibEq1mPs4e/hEPyvApBrN9xpPDfCddl8wfGohkVEGgRcLT0jqVHE7W
wsx11+dJ9nbLCdO3ex8S1Q7k0HX/bxf9mpsTUUZCvnmOwzDjb2nabnpECa/VczaD
095Zc6w5e0W4emXVBvWMnQP2yofiYwGgLlXTaiXPBagLHdeHl54aSqxxyByLxj7T
JpRnhgA5aDwWPqCK+6+rbjJG4G8HJxhHKUPeObSDtI+19NcPgDr3qwx0L4GkUFg0
OzWoO0MLFNAnetvv0eBx0RhxaoGdSxWBywWq0vx76RgoFM8p6Kc8D5ttPLaQEXn1
5nrSf2cuBM+oe1S0MHyYFpTNtT8Ucu6BjuPyMXAzPHGTx1WRWGt/EjBuoAhGiQ3/
oISedlR6/3Q5agRle6DMZRn/TUX2rlQ+/s/+7fBcpmhzTR9tMeSrqhZEPjylOd97
mJyl/rZrk4u8TtGta3LZjgczAF8YFmFFOBlGraVHBvLuMKnp/q3aztb1EeXiCpLP
Xv01z7y1hOTY3FPsm3IamDxhQp8B6zAkOVE7Vc2GuJ71UFVnEQCGyngzdXZW0lhx
n62cznBMn/X7iBVkcKeGeIWLzoZj53D3wPPSfKEj+WKCu1Fdc66c0qV/kF7aUjYl
TowdxCbSH0mWm4GnMY670hWLwD1rUJuU4e1oEfOl9hHHicjsP93dNSW8Pmjq/XNe
2AiPcI5q9SejL8cBqNMBZg70hWq01g7eu2TsFqe2FvANoT2hutwGTcGDEGFgM1im
m4hb8cNFuMkvim3+xprvUDVrwmW3ss1dCOaVk6vp8QafZS+arcdSTyCCRWXYI6UV
qD6I0vYL/SOvDmNDEx6/Cgs+IqXLjckZKfu82wLb68ijKKcHGK68L5CiErIfQ8bc
ya/C/DQaSjMCS9C6eviAbMYj5WRvgUDC0QJs4kMWkStqe24FokE3QjCnsr/sqgSo
X1E0qTnnK0Y9W1XcXAlQYIzWTaGcJ4MUhoY2mMc6U+5ho1b0pRDC/I3VNfTlWFur
RQWtk20fqLrjCjXsbyKs+4ab+3o/amwwr9hjVUIK2AjlOEHQD0H6wC+hBfUwXlOb
RJzcYhPoIPwwZA/1TCVVsJBKTqNmq8lDl7abCkX2p6cb82e4uFu4gvvvTsT3kwlq
cln6hBJcwHY/TbpwgOuTIWQjPtjoffIX5N++FBnbATWN/2rYy/lPKUAPd/4sdZUd
NnMUq7fKvG/T6Q8Hv5OTaSJqcDmsxPdRV+82+3QVDyDEg9sXHqU+H4+i+XXyN6cX
UBX1THqwRr0TODlMmUtmybA4Eahpz7xkiqV7Am3RDOPrQ8m7ro4jp+jhNritrfuf
nq6GfHoX2qEjIWQjvK8+Fn8FQb9Mv/lX3pAglia//winpBTdESvYX4eWyzMg35q5
fyOHhZac79GypPTajbC/jio/izj8wW6272Kd7crkYdMZaofmBMdgvkEVUTJVBneQ
A8uNna/CLnRBlXg9qh2bgAV5ytQEssfCMTRO2WrgNaGM1wHEEEuL6RkiTMY63hrh
9z+RfzMf/uyL5qqYvc84NE2rCcPLeLlqMMJzXawpU9+ykNM3v2mzFnq4L2sFCuGp
olU9jIZ1OPGUgnpcbIlR/mRwRc+kWD/Wh1JMNkj3Na0fdGbvVwDkoWJAEZZA8h/7
gd0kl99g0mhVjXcyNYIxwTZv+E/fzc+VLcSZIfMO09hiOKkoclTYcihTHrXJlyu4
cTMQ40bb9t5obb0xN8RKizsw5U5RsnFtGEiqiO3UHQyl/1IQMkJ+IOrN4Jm8N4sp
oi4vP6daqlqElgmE1j7YjDsdRzR4u0kJYFDH8si7MTea8fRssXj5n9x/nXWRA8Z+
ORkYo7F5BLjgofHCzMG9CGhqU2iUmbxT8Lv3hhE9moooShVmk3ahrPMiJwdfLBau
L4quDPGDq3eMlSoMNeZohb/IESaK5sDG2xdqKQChxRri9ExJWjuYmPAsgKYOaR1N
f6PINK7rwcZtL1PcqhB9N+kIu1qwvDuo5eXnzKBqVeMhVAhuY08Vm/aXamO/q4PA
OWEWdWBCqqbH2F21QPzcADHHiRU1cRb51E7oFqncyC1LXXSmz9D6uecn+Z5w9bYU
JJ4lU/WXm8eE1yGWFfbJA5BQ/YEAGEkeEpkgyQMeHTyFTHJPYG5kO4m+rKqGZqhx
D7vfUaw1sYchu1eVO/+4xrHVkXiO27z63PRf4i/E9xPgWy10e0lZnhtZ0+UKiBqp
8TDfcitsShgAzpJtYHvW6fx+V0TDn5yKguHke2lsLPbClBirLxwnew0HLIXKri3v
OJSNPU3JUo9mtrCcmfLsEXgAAUxiZxjWsLY30iXxSOEwU/VaRVfoO+LPARZclxE2
MPLjyHdSkXF/K4jfDjQGlLkV7nu+tNDZ8eLaQlb6YCNGUQw8XY2zFmDIeMQIeYas
x6R1Qwx42k0Rkj2SFI9kxoOpNP715/BWaL7CxzTBr5Lm4kvGMUs3P2kpwqifsBSn
ONWOnFwt8O9l5/72ZOn2EAv740JWKmCuyPmhvcihJDxbDq9GrSEnuiZBP/91U7A4
AUUU+kY8uEBc39yiyQjHgmtEtCeuvec/Coh6Oe2IDu8clPCo/KpJppSG3v/Q3aVt
Ak9VcDe7iKOitlFd42HfpJdZfm+fy1D9EOwPFTlHjt1Fxsztz+kYAQZls/wWREJM
aZy3RYerotYXnqDuOkw76s0FTC/shp4SmzurZOrxRI1t05a/YKIccgE+9VIwlVO0
WEeFtBvRHINLBgohGp61TAYCQRG+yGvivxmEmo2bbZxkrglq7s1VtYAYA+1HpCA1
LeaWBbW/gzoemFhjIBZIzOUhn3mGbqMNQg7qzfSydLbrisoZI/+7sLMn6nB/Tdqq
aOt/CLmNt+UPbjd1P19jMujr+8HOLw/YnafQBVKEYupJVd++PECGyd+ZBecYpoIK
uZsq9NcHyzp3CwmsQvYnbFeTkgZe9XdPUKvUkPWHNB+tu9kNWLrXDHXxCru/d9zA
ySEhN6llGBVfCK8QbVnVjaUFl8jlxK2uZz4c39aVoVy3Dl94iM9RGP3/WQ5WxJ9+
OBzCkHdDjyb9yOAce3taLJ11YU2MUioo1APbegIScWNHg3TeZta4/sRxnlW828jk
eAXoOPiyDa27L9s6UiinkpCksLXmkgyFxzf2USPByqY/IfTwONTHXolA/MlVgTYl
W5co7Ol1WrBP1PewMPW1UQ3rflP/VG2SN5Ox23uUlZ/6RLPQJABiQAPrdeHasiIo
W4RWCxFS4F+P7J/As3VfgICbrJM5Ny6dY1yeZ/l6oc3Y61fyHkPeTXjtiD8fe5Yo
5thFgYwpoyvL03EJBR5XOV5M2QqycvzCT6JhDo3A/94ijFI/BZgsH0JbQRQ4scfQ
p+shGlOwHVSuEoV/MGjNzLod2G+Zeyo1osfhNb2giZxbK1B86ZBvm8zAZkchl/4V
v/Sbt9TeajcK/LptZVk4XApZzVBeaYZsJ/shE996MtCE6VXU3xrxigfQHcqVMwNU
5fkLnEh18S01k/4b5OrKcGWt418MtKPrfLyIhoOUkwo0IpluCAih/QrkWuB4vr+V
/r9drshjsDMPKGXrwEmjHyV3TXPqOByjE7WYFkcTQ0FB8tAH72rJUfX4waAv10uW
2CiAL8OOXAY8jCh87nwjtg3+N3shC+HABPWK+l/CLgtgkl2CEUB/C96UQJcSJ5s0
ZiLUu2wrzcdUsSYo6kaOtP/W4W7tQMzvXTnShFsTl07Mi+HpkFjHyWNzQDAiF1C+
X5m+KN1Uw74aZ/pbbmXhhdDx3wqswTa/RXGs+9Yeg7wSYoWbYDeoU1mq66K0DbJS
+m+QWdAkNGg22haiJ/GqdBIs4fTYbTTTGk7YOnfdrN76ua84DzYtPmW2S06xT4A6
FZkKtn9H/4eOA+v/t7XZ55lqydDnhyOi6D/zGPRMYMaT6p9PjFUM99CD2nTfi9qL
gJUiRdVBDmSO83LB9rfEea4CToo9qeGEfLMzjAIlwSzP/NUosrXh3vKEvXUkISg6
wOSHO5VYxGoA6QQeIaLs1Wl/srx7b9RfandeBZ0WFbGr4m6J8rAFdQLC7FsEKeU5
t2So6jhQnoG4aMOXJyVMbFx/BGseANhLFsmngdZR0V+Tinvk7sYB1l0FrQIgtitb
uLMVWT++nwC6ioPQFOuyqouTrAbbIeFtRTLWygF/hmtihCUBc2E/pz4iSawDRZdJ
SCRODkhptxmpPuoOW7OzV4YPvD0GWC8p1HIPRywA8FShPb9JDUQW4ALpY6gxi7ab
jaI+w1C0/1W2N+qrEkTmE34WmPGxCIZ61HXnOAQLV2O9v04oelJNYBf8U3X/3Ys7
YRElK2Trxto43ck+10HBBI3lKfRdZf0FtL3jF4CDQNCyv668x2CnHM37qFkiI8gM
qL5AZySGLrivTwMXN3F8k3MTHePOse5dErAcbpRNJKuooncLBeAC+QN8lM+dietk
VI5H36kyCdpFJBd5Y57KEtvVi4XsyroNUZszqtVYZGbS4LE559FFsP3JoE5W8XAc
YKn03FHNB48j3VBZH5xd6ONrdGEfv/ogBZKvyiqWa8yK9vFApa4m65Y8k05w7XOQ
5HgEXt8S+U5y2iZaXNgmHqBjGrpkcYrv0dJFXvIVXsSurPao8LzNX4Bc+zojOyDJ
i92wbSlL5dkSRWXNkUk/zYC/D8BG1NbDoIXolJxtp9DfQaKA3eiWAmyA4x9hu41p
lj+QC4YvkhLxE7Dg6R6LN/DeRxcgSJ4WBovuS1kumLQjYALa+L4Ip/A1FPAFjb8F
T8mskvxqYfoVs2/QAt/reHpWghr8RNcEmE46CgAm4ZWsP9RUbmkStRdwGXEr10ws
03xutV3Cht0Y2fTSLxgDpZIudW6Z7KqA730Pyxl+/dcNCGrMcMqfB12IR10JXsjS
kD4zCS5/0RX6dgHgpWb6mcBLzjnUHMK8i56qiQPHlQ5JU4p2xD2r90JaghIg9XN5
oy28tuZj+e2njXQmjp8924HheNx6OTSe4hJnuQtOQ9KN2Nu43ygNGT2ricyL9cXD
IwOh7eb6JPoOBG61q7RimRXJVn8RqjWwPlEN6BKf6Vij1HSmnH0i4MTdZPJyWlN4
cJpza0UUa2Qy56BXdZXHpcZbU5ovfbWMYcv1j2Uz5xLD4DFf1uEzeBdKuDK8U/o9
KFYrGBCqsP//sGBn/qlm2xFgPUP1hMqHVPbZxwg2+EESbtR7huioxlAc4XAJBHaX
0Cf26xO5Wn6Ig7B6KkCjbJo1F4ShracqzQoEFp9PLbmCt4V3V+ASclmld9wGWAZe
Gd3vz4ZPsq9IPbqAO8LcjEjZPAypWoaRIm7vqHZ9sYlBK1YqkSoFvtOnSYSXlDtb
UqeZXkqLGAZbQpQ+joBKcqQDfjZ0FavrIuGT54HUvf0YjPWAw4nR7WitCMJQd7IG
d2Z4FRPF18YEMqfuqVsNNg95PmaINC5ax2G2qDniD/BTp9wwaMsMvr8Jxk3FDIRi
i0du/q+cHQII7smmwDmM6NWGxTBwGONW7lTHW9pR19rQlsdoNOzQJJ8XAg/OT+um
WhK/xYJ6xQBW2CPq+pwK9Ok8znGqOTMMZ12jAvZxfugELP+83d/hJtyc/sxBRZ6Z
0faoRLWth/1MAElXYVRqSBrj6V+E9F6K0rsZn0Vjac8N+JcUCY93y6rNER7TzqCP
DQhcitpoICsfk4306Xpy/kNNF5yHoihF4iVwJZ6L7MfH5xjYgY76PuA8t8M5ZklM
z/fjl+AQ8ujP2AkBeDnDzNkNJ12z2XYgP0sVDjWFL5LWnFrwLckq49NP5YpERIae
DJ4Uojl8M54aywXaLtwP12u2zTSqra5qaP0dqokoShlQumzI0V/H8Xg1kT6IIqwi
9CV81F7B25Xx30SIWrSdJJEnjfvofxi5ibm9MdZrapqNscsOAAnS3PX+TxhSRDJ+
7/UoqcEe77qj9KES1JpSYyDL8cocVE9yHYMnQW5A1i4KmV48eXbFJmi9ZUqjF1pW
Hx5rPPmxvY4HNbvYS8Zzu6t6cddTtfRmNywLNRVpFaQId4CxIEk9etZpeTb7kqWU
6MF9zirgCVyOBu8TZrV+4YuVQxZvLA3mRrxez/ps4EvR85FPx7Vbl+PjIe36DeSa
yZyomh/8BTeazBF9OBZqpYlzgGt1/HfR6RBwkKFS75EDYMOUCNykTraVLbm8crYG
HOKLGQax7e9LBHR1fqlG/7OGd8J8M+Ns4UeVdWD91yq7lFOWZZGPugCIvuxWjCR+
XaReOMBMYzckAp96Czjh7rp371l0a3hejbYnjacDLmwGw5q5dXqw8TJ4If1Ai2fw
UxJV2xPAz6K+C1TBWG4ewRRuDjyugz4rgW4c4CCQOPw+6opr45RfBEH4m858VZCD
CusHcl9415oylBCey7JX65W/TyLlcfPkwppiDruAzYNF43uC0riGTbeJoGLDS/ZK
5kFvxuP1NfHuWuT1dvDemygSdlbSIToz05bTJQRj0yUfDuxcNvd+W+0EZ7yV9Opc
qnYjponNabbwLJvD5RDCOFCOoDLLByKE16ERU+eSvMunzwD4vZo6blfTRlVCDReJ
mVjLCim8eriMixLVEROdqdY5zh8Mpj3TfELMHmfmXC4IBHGkRBN6GUMNhjlVJqI1
gQQmmMoKR9H311dKva49ayeLezb0fDK+E+uA+YC1fTN1WyfHLNDnZJQC6yjG6opL
J6n9plcIo3YdC7gZFUA1jVONZGhlYSv886Edk65yNH7ob6AyRvd0OlD+WKGolBhq
BRSyVMEdQG/165tYbjMIUvQHx2Os90MkFuqCtM7qGKZk9QGC+cSNMSq8gXze49IN
APIKBm/yVHg6+RA7vjeL/1aQjDNMakKwJGPPwLaKQBGZSIuJfA8mjSHC9NjY1mqs
ZLjlc+O5l/lgpRNahLeWa9KA9ojcc5yh7giwROcOgGSNPaB7QAc4/52AXEILGltZ
ZpbbsOQkn+qU20Q7kjB90bCjVTShbsOGk3LKZ3BPl+Cnmn1ELPI2Jr7ZWR05NuOi
vkugRJBAI7ld/mXAFmmdWW12blINNL5+vvuNnIQb2k5XNAoTTxKy7hwOEQUuB14k
etNJxInLQFoj+kKnDujAU6GkHRnOkWJTqq2i8sW98FrwGsdZttRm/n5Q+QH7Qv1n
cMUL2YwVPVRYu4Af09wZ1p8aphG105EtT40fiXmET7g4v+GoftrTNLEXFSW0QQvx
4zA2sy0s4g3Xqq3Cxbh+b9QkVKzL3nY6TwSg02FTfAwF7anwaCJRzI5VYFIm8bHS
Moa2wbZt4vnVsq+pKx12RtnX9EZmeyYz1owMnZyApY4Rw+xSzVHp6dN004Pr4tKI
Yx/QdELhFfo7kBM0FULjNt46zfV1RnfBCcFgMsNbcPmtodPVbot4ZOgV9LlWueuq
RZqzrgxuVfi3cUYOIgmiiSoz/KTwKhLNOfE0bjyCWrNWO9Lzp3vFnIyeiEihHvlL
ecYmmnWeyE3C2Ob17i+0hSKsV57+AzlmioMsI6tLUZ7a+z0dJFAWX8YGP9n8y1BT
8oO0LUGzyhv/SP0WcOuQW0kzjT5/SNl3WJG45wzocMlU1Uh3Sa42qfCpYer+uS0A
txE7oTWwr+xeQqmT3pZr5xRNrCS0haV9/ohaCSb9RYk2lnSGeQlyPaVsaJBTPz0h
5SORm0EXN4CUyElaHe5WWd115r/h4kKvNke8Xt0KSJ34BKojXS3adpI3hT5zZFLx
MK0yfBum1rkIxe873oRmYgMhN6CNl5L6tMt2FNCU4QOJUuc2YI4rqkDG9wFzfyBT
wnevW/Kqn96MhvhM2YFfPXLXlI7p9o0CD03r8FNrniWdny6zjjnTtVHS/xc99qpR
IGam60uCH4yWI4z4Cr+14sPmFhHeUZO3rmQgA0ZKfmcS5BAK1EazfE6FHbeea0eG
zL9khavpCBeX+abcURUE/4HY5guGrfRtIA2CeAN6jeBF/X9o2RczzpWQQzbf3Vwo
GwH0E6MbWqgqxF7LXzkBHmoUaQmu7GOERTkOpstMqjPF6U9+CTtEOSHDqJiV+9Ok
I0hcr8dBTU4OhvMRnouH9hZB2Uz9IbOYPfQvWZnICkFMpwfGrJoa3AYq6s6xh1K4
mukmuDv3M8PCoxDqdt4y6pMt/3Jt4zQfLMgPBJZRaEDc43SuwhE/9Opry35x3jAn
I5YlkA0lCZgaOhv5NB/xhoiGnEOSuyf3AOgejS3S5fSrJu+IQ7MU+PXaR7hKQ8A2
DV15hJXroKxYBHc6/fNux5fwHwsGtzIXlaXUJYrBLhMUh9/q89ke/BAhVI5VrCJs
JVEPFLzHdH+0LtUovG8UFwdUklIGSCIYcpeR63fnk8ezjQdtVMEoXEJwZHJCs2m1
3ZZ4MmlJgY/vWmQt1gqlGfRelYYrPuxhLzhlG206sO14OflbUaP/cX2YZTytWM+q
l8sMu/tHU8g5T/9IhSFH3swW7gFAHWDMDewglz+zDhLSmBl5bx34YJrKYHs9WnB2
eHjO7TiQAdBQKsHoqjDnxg5bcueJk+e3j/2vd4M0MGAjJSXZBpvPTHTUKruzz/oO
RUpbQZ8rvDVS4AxJkiFMCMMN/UHEoAvi79Ew6kms73w9PoEYqtXFza/e8BhiCvk6
RbYw/rtzgx1HA5rLl3+5X9RnzTInvWHsqsEpapi+Wl/2umTLa2Mon82XBsN/0IFl
lxnA5clblVkmm4A7BicwdDkOgoQQ34D+Zk4QEdTvk3Plre6VL+kOiEdocFpUIo8w
IiRYl5YTIyye7tsQ9ew03C1ZGmBpuoJxltUcQHFVZ6dgN6fRImfXCg0OsIJAd8hW
8ytgFl/qPLzgayGHv/gfzX2GCSsFz/tjqUZ8hYRcC+u/NlHN2jcJxy5DOld9pK0c
DJgI0lKhsua7DXm4NaCNPnoRie/oXD5krw1j1FSLbIfPMBms2qO0+v5c/oNBpfd1
Y2IuEYFvRuDDxlgFwdFiwUR7sGBJmppdAhO4EHL45ejKppM3EpgGzlrGw+4N0WUq
lfSfX0u0TEuD/Dh2zFWaSm601S9YC4UMrVzzqMLKDFS5XJbVUMlPOWHOmRXfzc1j
t7msMbv+rQlF9DMgXVbyGzia4BkIfD2jejFXVS7Iyn5hRg08MPg5lQjbodNbB52G
gZcKfq+L1q6h7yPgId23gDneaxjsT7oQdQrlTGhuCfkdxvScVmJDQYzZEk9wm86Z
P7NbexLOH05BRdSJZlNTPlEYGf7noVvWGOWXNY/43mT/pDO99buLKlChjvXbRbLA
sEuCF/mnCpxoQKH1VfeZmmFNUh3oDrMiwdMKQgxqfyAfddn5WxAM3fsx8kCAZbZP
tA8vmMr7T5XgrOvHGf6S/a1EnSDODqUU2G65TFUgactqxFZdcU8cSUsOih2qh0Dz
14q+naTkOoIIY7F4G33etp7jRfo2sscwRv+bDFktQN1CTMjtHG5DEYm8DyIE7vfS
OpJxj6o7fQCqOdNKxCJOv4dRjz6soTTuNrWPGX/M8bsNdtun0RTxxe0bRY2Fp4NJ
CWdOBz3OpBtLHS0OWjvslMYZc8utqzVKt/zPNf0+PPA/vrztYCHce3Fmj90GjT7k
T3Etztacb9Hmb85X0dmd31bosFtSf552SQO0cSVupz+56sTXXu+2pH7D+0Eu9XI0
IdqySyne+kfL6RmeVaYjRzo+cc1iMk63Wb8ZoZIdp42Qw/DTncCUgBW9ERdYeKZn
SHmVW6YRLBp1b1qF9H9zaspSbCQ/TmktMLtS+2W++3U=
`protect end_protected