`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 20320 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
/vEkqJfyK/81z5lf9X8oFQrc17ufBsoVkZNSa5830gYBGpa0JVZw6Ld11Sw7yIQ7
XnBIWZtjdJCNIrrR175aO/tqOJ9qcO3VCsvjlMutuE0sGmm0ILJAAS3RwpFuBYJw
liFujoo7pdZSOsjNdsxFhDayvNFQC5Ictg5IMNk5ebFVCa7IeEgX3wEDNJG8DNDJ
64Zwizjk18aruLOUF38B19TL934Tb2ToS6uHe+ZutS3J0On/PXvQb7iyCwa4yka5
LKFAIZdI2CM97Bp6faVYurifPa/fNXA8ryx87wTRYG7vCR4T7lw7dfxiQ0SWlHMS
odgaf8OppLr1oDE3ZI6kC0eWvaCQyFkzM4acLcAiVQi0dr+//TtSSQPOkKkgq/J6
RA7S77bjAJi7KiE9EGtUWUuX+P0ZF2iMapRTyg3w5Itt/PXHXdURCPrTVUbuAWo9
II3YpGKznjX+dxOUn+teH19bqFXZoA6Ox/JJoQPNPHzBr6vvcElNVvxER9gi3jUg
B/mJeLTQeWOea41K+k/FtIRLKp4WZnQSqs/036zzawsVBBOzWNxWfw4JGcCldDhs
yzOpkG25yM5QeOlwDXBALmBOIk2NDgOvsk35n2ue9230ul3Q5/ud6/3l/QnxL4hd
GaTcrmNGcusDGpwBOxaxpLBB7MMAd1UcxN9A6pDjc6bFqPJbl9oolumTp4XqaAyd
/BOM1BCu+8XHFQrQSzwVSPuTt0krjhV2RiF+X9aX2bJd8DzlLAy6mOYXFkq/D+rH
XyUu+aB9v7DDj/NQMfw38R4gpOEuCMeN6PKW7it6m+IHqXgbs2MFZYnn9gWiYazA
T0MYacyB7LQ8QqNuaaf/5Nm0E4Yh2n0sjv3WmDIJjjkkwBpccUzJFKqgcQA7v1o0
YktwVTxaJagj/aUfCKq+0kUZT2FZ2TipptazBL0chejWwYslu1jJbCy4ACp4ny3Z
GE6nbhRxn8TsZ8tZoJMTbbbqCO5n9MO07RUC3lHDSteMDjJKaIzFwR3Wy/u+4xxI
8frkGSUZTudop71hkgcOgqeqNCx8shWQU9h9QRoDYAdbOJeqgKYIa1LOTzBdvnlX
kMQa7CnqXzfx5b97HVVX0lTwEb+25ZXJfEBtdg7zv8A0YiRIhHt4fOkKca0T54C6
5FLp84LZFoFjrSXdFqMRhe2/6bcrVd6cNC8/PsC+Adt69sho0fRC303+O+DlJpVa
R1UZib2GHnYqZovXTC7Rzl9mDHbkpQEQTAQJVYrjqCcP872j0m8u0xfZFjikmf1m
9UvFaC9cYwRJSn9ISW33xJVBrsrkogJ1sQSDnj/vp5CVG4GS1UghZgXlZMLFGVVc
RdHQCuqcVKd7M1ztdDzxAAsZtRyQVKBSYR+OsAv3/kiSFwcyW7lNnmgNl6lkTwAI
SyzpQRq0Bobywz5fbw8jQQz0c4GpOmlFs5T38DGKMuC9H6BBNToCwaQcrheucUY9
eS5Iwocq5ImfJ8+Ad6NXtJnN78RXjcOLSXA6dkhLUiyhpN8zg0TfZpCwTlgDXJYP
WAy8KqzJWCnllcKhfr2Qiu7kL5JQq2+gOzSnQZX1L92sBU/l2WLEBocueGQIHFLr
2M2tXM/1NAze5dn9Ct5J6FYz1dEHp+Bm2zdeaRkWBOoQ0AqVjeegW5SYd0lN/qzR
oqBkzn0ZJ+j6R0wBqiKigTxhJibaPvztCkKdNB5QczG4RvUJymNAFIRDztb10Hgi
uJ48cGLzrunlKbXgs6BQFBRoW/YxxgW5LVs6tgJoMDNbXkJ5ZduqGFzenwq/cH1m
mzbmRY08yCk5SDI/+vaqsSE1WMRh+sN6AH5be+zizPM40bhBqt52sbnsGTCKqUwS
s2puBgPfIBAQNoZGc0BlQ5BqXeYQ8n+k2ksv1VX8ZhZcMU8ithGZO+d0+r+GEQVX
g4tGnh5VbYc2LRsDvozAifYSgegoz6uHt2G6uOEwrTqgjl82mAQRTRwl0MRDUVQI
5FFoD/kfG8mqnwK0Sw3eRViwnuCrq1jJYIsu2Ap5GrncL6Ywlz8IReRijNuFsmHG
rYRIVwZG79i0ysl+Tz56jtQkFIkWTTRZjE86B1SN5xcFSupBLcHctYSUv4gUrD7E
+FxXjn+hLfvcdNSnkh+05AyvMwrzIS8D3OLYvku1275gISNNafB/dRujv/zK7nmY
9UDbTOuRthRwPBmYdp1Ui61yPgoDXt9x3g75DTL0yVKZvhneVeHgeJgn1ntWiwMl
6PJhgPnMuMLT12awkS02VmQoCn3uUvUJmyAM8M+wz9EpSmDgXFFzrEPMUXE08s6t
vmVK/098TE0boiPNfw+TJPckuN9YlVbo8daepCthHHvffU5KWjFYBD4oUYbLPodj
uXpGXj4dd7QpSg1aUgo1xkzLcbPKnKGGpzTryJwOU7y0O9pp2CsrRL4iILrwa34H
mamj9av2q1Arb0q2d3Z0AnhmwWWqu5Nk+e9n8BONkCNZ72z1sxVCrSibStntx95n
1ytu1BzVNKJWlsC0FRRHtfKyLgXKFGmbS81PpFt9J2FiBom4pYVgSCX81+WXujav
+2iuFkpybU+QuYFACnfEe0L/u5JEQqUOVc9hn+f/ze/1M/srXwqlrPcTlbmfhwMu
PI2hylvfC86UpJXWHXrErUXdd4ola9dHcixh5N0u3bRK0LkRJ568BFfR9z5Xbu7j
gEh4/SngMmCwgTQc82FE/yRUv8Gv1+mc4CSd0QmzgcYl8reevwNJ3vM1l2Tp724o
ht9+yJFMBDxRRDTTJcNQH3zW5wHiYNTPNxzMx4tZYHi5/h5a/MH80vUz5pGovkys
D36omU8PF7A3+LxNmENpKFpGFOHMePjao7m5auRVizgUcWPlDXeWTK1B2627CdH9
aQOJc4QJNprJIOI2Jy4WUI8vzeb3qajXgTloKegQe9ubWJjqhOKlYG0k0emITXJP
YyoFzOgM4mkl1LindazaQfnDANA8PIGMYKVxgu4vF84ovIWwZlNvLG6MAK/pCVC6
HjLXrVocTfv+tb4iN42shxqBRi3/y65DxmxOxg2nOmscU91RmG2uLSt52/Ztofd5
M1Cjdn7OY8jchhg6CzKIEjCbYs2HEbdnnPSnk+B+TPFufa5/sAD8S/L0T+/QchC3
+eCKS3l/pEf6ftBXTB8nsgrzqEL7JmnzIU3GzA5A09RjHXJJOmlfkxlkJWk55407
C1+FTy4cVq1B6l8565GLnkWj3zwG1OIUSNz5+H2NBOf61DzyJlIoq6lLkfBdHMvy
JK9LCpoup/2EXG5xEVWvxFRo7r1cImUcJcLmZaPpySGMwM40DSBG/jAqPDkakIWg
Ggf/+FSGMhyhTzWw9//R/ewJjomJQQq0LRyD1lSWbNt2ugQlkalM71uxwePd5IUP
PkzSgTKF2CpH9ahfUaNYhkPdHjD3sopWTTPyXu9MfJ0wAs2Mhsdcovh2RbpPcXUp
uqILIe8BbFOZVFoeXpOm0BP89S2ewNm+iHwouUS9XtfbyvmHLl7bTcc17mckWD6Q
TN4itDf8ln92KA1O5q6JwHrZN4noaIMCtsP+VZZ3sD3a/XuB9ImVaB5XJLZdPSFu
6aFcsp6fI5eNKBUEEoW8rMvLujIZH+5VyN13L01LSZ/XSPq6dF4+1Dghw0lFxyrZ
DTODT5DfgM234s4hvv5KbR54KlsRV31FnopMGUQkckHGtb3I6j4cAOeSgbKk4yOW
bMCdd0U8LsGsT7Sy/HYPbmTi95WjhECLBpBi6DhIvsZb9/vCIK0EMz5AT5odRzAG
aLCjVE63Dl+W3k9obKfb0mMfRbYfJNcgnt/xf8QZGiMeCjsggjLVsbdSqhmnK7FI
SwZ+28VGjFI+sbL8mY9TGkVTliH6gpvPfmDnIHkp5ysr6ENnQDaL9mvxCidwgZ+x
ivJjRPl0LZSelGgWm8uiafDkwz+2SRDLm/ZW8gVCogQdusq8JB+bA+LTw7HrMQUl
w1jkr4GQUVOUleNnaJnTRFrQjsUcp4qL5IJaYi65KAoi6WgssWdIXyKm05Mmm/I+
Psies3rUWkv3IVqA8cok+6LaSs6UWTHvsOyBUXgLxGRUd5EBziQGGPQxV1qlvtiu
wYAHddnC4SK5r0EgqI1OMA2aFXCmFSrsMtunaI29jp1siScr34mOC/1piTYjINj+
t7p+qXeBuQj/FLsCp4xQlgrH5cgLL9bLs24NJRF9kzfC+qm2xwFJu7TLANO3c8V6
qws6YIRo7xIgntYk4stesReOmvxCWCghROf/W80LSdCTXgPCVXW9sA/6GVvsF2Z6
Hr4DLkm8kuVMYnRmIL1zldjPYIRGAsEdZua1XUuHCbaFoX5MKFgNM14VNHk7TCyH
W2Ey9Nw+9XjLOBDsdIOlBlwxncJ0Jdt+v1Vl/EnWAS6wrxDIfPPonUoEU6u8slDT
wvuSx5/TPTkMwXfuJBt8j9Dj4OpJKWJc06nEMzjxa+5aykrljPHTEo9uCBzgacKi
6eKWTziDal9aEzdnKVU46UEoYBj2OVSjTCiDYve7vUbaduLI44seQdM/Kbz1dZCJ
w+NILb9uwVIQ29/W6ggeIrKjSHhh4l9g31eBnqJDImfH/R4O6RAfbQrPN8AMBmYh
TkAUQkjVcATGke0MsnRQd5M6d1Q254n7Fu7pZsOPpTz3tTlw/B/q2U+teWVoILXo
+OKAOcePM3BlNvhz9Iq58Dux751aCaK071id/H466KkgtApSb8g/jfulH6TElHGg
eBDZMBrK+W9EbnJzKW/pFFbAtpt3picepDk/9ttdIzCl3PBS4STGc3KknlqchV0/
9l1O41CU/oBqAQBiqAPBpjR9ELUPFiZmw7pOIgvUUns7uWND0oT2Dckx3bWZU+6U
kxjxUsMqtOsEHrC/Z67ap1vQm4YgGcO+Xx7PNrdq7yPC1ZkQh093OnD/TqaeiiAW
LuXQZmdOz9PYpXhx6TJswGilTKn/nbx3EfzWaOXIPrtLZafvLg33kq/aarRR1vBN
eh2fRce4/fYtEhcHzQMlG7MwhMeArtUgzvVqwZN4/e/xM85NoJBSCe/WOcKnyYLU
vMEQfGPd04cCy3ubJ3QYaoTGRb9+4fIYTMMk05x/csGDbpbP2HIpvU9wnh29zDRk
9PLOu8u06i47OX414ML+khVYqoCS2bex6qejYW/q2rpf1rVGtwowNLeFFZrNLuQg
zIcvILFV7S3AVC9fkLz4PY0ciRNqrotYs5MGBj0EbJZC2HSAOVbIuKIzc2ACzMip
WafNeSMvUSSN2WAxWF0TqMOj6OYT/J5PUsA5nnQUMBg019NXcQIr/ZkcbcIp9J8R
KBmCd4M/z8yr/RZpUtzqrM6a8Gw6y43pavPadZDHOh75SPO4vtj36JnXsv7EdiGK
qs216Sx06ImGLx+b3092qx7NUDadhHPl9XmAKUVUFWIYgF5nBz54vTBNUTjoZs89
Pzpo7jGfdBkL0cMmcQ5irekV0TBOnVnF47OUKuxlFc0ViI6DoNgfPDaLxPqbORk7
niUUsniW8w0LEG/oWSLmWDIsBmwWMCZjtA2Do9IymyQLApoGyx63VTnVy9wm//il
08b2cd4KQEnW2dD9b+BpB0adIQv0weo/OzH4HhYDzqi7GsqlxMaMDdsm/zKnIniI
e3rAjgonKL1rk/tL7vu6iYHwvfmw86pJJD8cdhZqYOJhFwfG1KJgT9z3ERpdsrVf
k/BqHqPo7YfEK40/8PUIfwWtG9/SXbAcRsJsRS4V8m/IEshSiYLJokbKABCEH6vh
JOL71tdfFS7UC5bkdxkD6W0IILV+HN3kaJ+MdsU+kxH8Fth0S0jazglTv4zEs9I4
EyhSMiclcrQxKOnfRZ7B83ygWjC2SV/HOfghAx7aie0f8LPWKDar6qMgycAge02C
+RMOvwgKGwTK8ULs5aAE7h3V2d+ly8Ws3Qzq/RH05xFsZG6/QobLiTx7aoTCGsU3
hJnh8t1TgYj6MN+ud9r97zCHOKSwXBdc/enb7m67COs6mBhDZMcvq/COevvZ0yqs
t+e6tq5+reaIYem8IxoxPu807i5+kuMk+8yW1OnimhAVhlOdABwh4SpYNu1kb96e
qghekS/AqD1rwQDzR4xbfdOZ9MdAUSRjYJZSA9nVXlxdFhZZUpOQ1FDCJ7UkFgFE
DUoVF2xLOigLIzjTFHik37kcGFtSyefRjMPctTvbFPV1OtFOriQrcK6HYbXG8dXl
KgM2kxxBdmc6FWrVHI77UVAqMJIy1b+mEi94jH99/AVNALYjpDij6yR5A7oNNTMy
Wb28y55UtTCPBVbp7keh944FfogjSIOEV37nzbG+GlN66lI5+GzXhuQoJsNI4a2E
qe07zoOfVB2lNDwAfeQ1NP55QABjrLbPTv2a0Jx+JZ8ISGBfdrfzg1KI95tK/FFz
p1Q6VcaUu59WJ1VVdJQKDZ+BvEE985euMsY/pTUQk+9BeeQ8VgQjaf6XcwwTIUnd
puUf1WbQij8z87iHK1r1jDo5xEKR85hrkqSlKKyZ5sEONGFrV4XB/l4kyNHRwcdn
eqzEe9/GibTbQOPTxVE73fV12mnqt2cI/9m3c5tD2m2qzsjeTsgpIGFuGbWYHTzb
A3qFlTD4+u4VnhWe5lJ7bjDoBqzkv6NBsHQq+izfSATuAd3fpM/NKRT5k2ZmejmJ
ZqbJX03IPR/3HfQXz61UC6gvv6xXP68/G12/V7mMtjiOYskn5ErZCVP/L9p7RySM
MaoPtDB+C2UKqwKAsdme264RL3BINph6vqn3DOoTyudEL7NV6vFYivzjsGIhO3qg
miqV0sTsgFCSoAETsPgllt9DqotwlMxecK5RDXIvpt84OCYGTsvMGTeqaoF34sqa
H1N7O4Ic7N8ixQh81UT68AG2v5y0nyQ8/sfu0/bS5LjSpCM/Z7RtbKxLRiCAX8ES
G/HOnz1DuY2TcR7ddEWYXDi2rPjXtv8UBe8mqb8wbkmshUxkrHMy/OFHikq/pGlf
0S3KXlFXTtJ6rCObcVQjhD/F/bHloPtFEapBH5br0jQbzrp/jz5AWZNyZV7Ds700
Pd7UcJCM2A8JE3YrOia5fDAVKPctEWyBB2Wa1yL18eKiQXPSr+SD/9bGQr8vGmj6
iGU+0V7QNcA+pz2faUuXHqankflgA5P86T9b5N97UWW5vaNQgDwzwf3ymchU/tE5
yKLsq8+9KVczf+XKV4j9eEPWUhjfNcC9BAkhNqRkiB2yKKAitn0k2PcuG8DM/810
7qvBF/wF1hxxfJczISxXh7H0cnWqckGMGxJjFA4mzjDbOhRhC28hyEGDhqkNW2cv
dFrfyzgXGyhWCOOsB/Dde0GKJ1J0/4tpXyWKoUZqUV1CYB1lKjLUanwB7hPX0iwc
L1JnW1l8DqAs2XAwWBLUkEoDSXgzweBhpjGCptj13D6Z1Jq399Ki7Ei1oV82zzXF
rzOJ4qLmVg58wDVYylCqAdj6oCU5zdN1KldYSziuoOpRaR3uc5UzeJR5escPtxcb
4Bxz9fE7NnSjlkK/RUT+ahpYQcMugQSaFmTJaT56HdrC8n+1b9tpc6AGmWDleG8E
N0ZqcyxA4mqR8mpmDNjTCqrAIs7TXhieeqItnru+PDrPRhQkkgRvSzdSCMWhVlsw
zS/K/g7IuXkbs7NVA7J4PrAcQXMJauTVjRoJKFMKRThhgSuLEaDmMiA03+ugR7DF
kh47/b65ii+DVxVPjG+x6FbKevoU20DFhZJvrNvNfFOwq++GL+tPSrT90SqfKqw9
uUj6BSxwRcJXJNEPV6sm8bhUN7AayscWlR66O8sjPVECar/uE97AexMolmBfrR5Z
sr1b2xsi641YqCABPYXs8oWhAvw+U6tiGxGEaB8MNE5cKCxFsUydOLWZCXBNsKPt
vTKOguJ0e0KhOnOP/vnKUINPnig1pf5VIoeWeFjhQSIHKCQDuQ3td3U5Luffi4Ws
tS5L7kwfmy6TfDdRGNyi5PCmrAx9oPJixSrZIoGHSqWeOnR4iXiwD0Iq/dWQXqCv
YLWcerXbWMIqTFNzxO3wpUJNH4/DVTuGCcAKq6f90LwJY7QKTtNAak47E2i2fvM6
NoKMzxOtGpRcWWQOXvjZ5Jdk3MDIav1qLnNpGSs754J0tVeCL7j63ioQ52NTKank
WUk3+CUW8lHDI7Qj69lqfBOj6NYKTPhHnGzdgLMC9KK5hvS7BOAcI79I7zP1wshz
j/5gqADFtw13ipFPDKnFiM2rLrFTZNL1Pyba9mwUYLA25dFUPHrk04mUSyIbqQQf
7d+EmeT7IgcHx4SarJIhAu54bsgJYVQrQ/PBZLWf1ZekpmQFuGtgltpJydtKN2hu
ON/hOFuRYyZLx0ch3MjCyOpjCnk1j1ZNv1g4kZjbyMaE0lhUsSjmJVZOI0x7xmd6
6i5h2GKdWQedb+79+j4B8d5rpdlDkEIAniu4vJOqT/aKI3ank1DWaKkI9TLcGrox
rHWD7IqAsHBPKUq8KHPdDimIko7CM0ymIQuWCwhvr/3ObGcYrXOrp5issEz2JxiT
gBOmZk07JcGrE0l3RrYrxhZ14l6kUaSoM7vOoo5oyRpjLkJ01PPrjtlmCUexWbSF
EhwfBmmQoUpz4kZxWt9WQe5uy6XvrnbHRJsb8ybMoSJxyX2nmVxG6Uvq7/f11tsq
TFHH+wxQrkjagtmSsc9TwbPlNcY+K9pvcLDRicuA0Z5JTunDxkBwuwZ4JxqshmMr
6g2GsOws5ABLND4Qg87scbv+Nq8XZf94C1NKQhnYiQCEayVhTLttstYtfkV9dUHm
yFTdewfJqOgDoSirhptrdJ7/GS5MJAibbRa/h1g7pWpj3pFziiLvKaJleumUzUlN
tKX+SgfIUPgvzHyHF2w7L0jkSzye8W7+OVgVrMcRAVYxCJmueTRVkBoNGlVTCTY3
4ttz/yKylWXLso0qwA/LO0TKPZA5zCSTlFg/t3wggDCB5VvKnLNoHTXd6jOxLHxp
y/7uNopGJPvbraxnsOJvXO6pgkneLdV9/VC5FdGW5OasSk9NDYfoOjC/S2uhugJ1
86NdD3ATOgpodkBRiu0rErgU6F29D6AZSd/aBdeykKi+I1+OQdmGkf0w1Xa9q3Jx
geuG2guNpgBc13UjSYJYmmonPDySbLsWJgtkl5sh11GziyCISb3BiFNv9IsBCBD9
8Q3lkSX/acDBlypX1foUV+ReUaICRzHzvyh58JTiFUbNU/GJ4ABYJjDhUkuCBamt
Hib6vdUqfTdj0nKdzSGKxqcVmIZOnEw5/pBSO5vrf/ad5i0XBlbJAt4BXukK07S8
6d5dozR5pyQOEQi8tMiKDwwPRUB6Er5fHL3kriykCr8Sfte/Fa0p/3/cMYNf4aCI
qD7iyVsYiCfl1vQgC4GnnWFl5fEsRkgqjV72VkAe5JmBa/5EnYPqF6jCC0Q1bv1O
sMh/EHI8khm/CX9vVqPAUEV68NqpEzAsvle3uyCLakYA0PyA5YMGjV+3dSANs9Hy
QKdJLZpiWHZ0QMZk+isnCzUHCTIkT62wFvfbjEur3ho0avxm2BzzQ3LBu6hvKKJE
NaUtZPm/97Ba9bcagJHZTxufvn1g/PTYTrQCDygUq4K7gXW5p3y6jkdZeC1YYW1n
3tb04muwkkXpa7RWOM6RnoiP3VksUNEleSfM8TQ/r57uc8CcD6sGi4nGR0/s/QuI
BIy+qPpyFxWK6sARvOIvqw10Y8/8s56Gyu4GrizfZZFhx38DxvwmOa9vPv+2vTS3
fIE0RkSiS0VL+5IgubjBOAyclRnQCYZ6Jj4Xpbi5kilPXYUtdvMnsIKB/pkWNhGH
qlCTFpPaj7r9nOF92aiT/x4HTmEePymt2CVr13G0hJTsKqgbkNDiLELeIiqgdc+/
DaC8n3dCLp4+auq6mySQPBaF/Ndg9MBVZK/H16jfv3pxuq5jyGtuiEYZMc9uUjWv
9iYzVNzCeptCSKWXoHc0/pWRyf3sbULH75dkKr2INKn9m3szzaU65b1bzPic0a/T
AJ5Yeaq09zLtqgcBQnAu+3v/GKVGRvsWPmg3kc6s3Km+NbOJgv9YRcs7ccq5j1Kr
TkPenWL9328lc0L39plZ2yBE2Sypz2kQsnyA/tbP3bLijeISWyY7hq1SqKUlyZy9
1EsXCHwD1S2marOTX+JOULDdL7ZX/DYz2hl1Uqgps3/18o5JEWadg1M5WpiE+jMW
poIwDWgk5LJUa4hca28y7kVjrWDw4Y9GFhubwmL/644M67R69uLA4PWn4S3d171P
6Mzg4HfrPeL5DKKthGiq8qKtEZmzXAtiahrks5/eQMm1Hc3RsTBflfSwTLUOP99Y
3MYoekCdRh2+TLK7b7yF3Ua+GCMWOoEkAYdTbkTfHzUfO59I3aoOHkYs4Up7Q+6u
z2d/WKOwHkPpiIVvDGK0qRPcYdOQYzzjfrThjGt1Q8YobScUzL30l4JXZf4bxqNi
dQxmd5Jo/KbrsF3hUzVBiPegQrGc/3yVlN4CQLAg8N2jsX/RQ89iSOM+mUiczTBn
0Mz28EhfmHMOYePAp8MybPjVb7mBIhNM67vRKpTbhfKhpi4zvNfEEntZTobYo8Gq
G28rHhe+upCekgrPTvXVS0ALwV94+pOlXGOFaWAEaQINJYg+pcaCdvcMH/lgBn9e
J6XSSBVRg20nB75gshqKQnj5MUCFqNEj7mNmSFaQVYT8KiUTkcbPmNjpQwSVmL79
5qVRHAEQTaJ74gc430K4B7X9fT4NUUKK+sVj+E7zY1icsThp+/bv+bua2gNPJK3v
8SBLPyFXIBbBMHUlim0fHoqaUBavkoAqBJE6YCga9BpnUt7/7Dic86BOxGt2mxks
GXrtj8ZZ/SWlfS/RGhtLN1YYU5FY8SqdPwZ8+TXpGCQwJTeSi1JIPufCLvdCNNe1
LW26xM/2PbDgLNwAMCphJxaFcZve4SFu4yNLCigXQP0pk9A4ufIThdE+iZhswA+Q
MH8f4uHnLEAY+dWhY7tugilm4oKBYatwcc4dBtZh2G6gXXqc9jJ75m2rCnxtJxby
j/Mza/qUDgh02qMJa+DQETwIM4pXGaIeZb4GnzlWfx2zMXxzX9BRvK+SZAG8WIxf
TQleydH/coPys+BBtd9BVu5Ue0coanxYIJ0eOGBwzI+hNUuKgs9hDvOh0VXwamr/
9R6wZxUnE2zqlWXYEcO8BuuZrXdgh+pkoxa3Uu1OADWZIvKsnIFXhJ9bFxsnXTOs
ITiuYE9/leyUr0MVEwmXv1TThkG+z71Ikcqsr0op2ZIVPglJ8QzhgShjxoXfRn0z
T07rffKxRqrNGPCYoThVSrmDVZh8qq/edy7wj5OIivHXiZZ179bPegjGkE3WNVoY
ygUTxqE3Ae8HzxKGYdfADyi21/z8EbI7ALo5FcB3SSCCkW27h8tqJompDkFD2jom
FozAhTUMYQnh8C++T5B8NTBbkBWVGn71K9zL8yyJ4MzjkUILd+uehtF23MzvSEx5
Mz+0UpRRN6UmB5lpqC5frMqeValvCaK84NVQ2Q2L42emA+7XlGNuH+pBeZmBPDsn
nUrg3miYIIbiLvBYkAMKaDnBKhDP/vfA8xUlUPI3de7v+sLaDYlFgqEY9WzdIUrY
YHkweE0s0ihMR2+KhXcklPUdEtM0nBGax1/ZLF+Pw8M5I1G5yYd+Q8WTKRWty55f
S/SxmcqUR9jIvjs5Kb7eCO/NE7OuapM6wCiUxdx8j9AngEL/rNJlEWgV8VYoJtay
ZnAId8lUtbKlLfUItAtbRZqbyvR/H+1WP2/dtAFwClANOsA9yiJWHXseY27a3GXC
lMLmgMcR4tQI/YW1t64nDbiLHcmMyP+bdmL6H2KiqS8cQXHUu7JlGeuWVfkPJQOn
x9ou7+m+3N5jsS4d42lyiSR1WeALBw9gKQ42U5q6qkH+cQYfH/r5RuZb/oOwS2/U
vJIHh1SmZ63xbZyI/ycYrEeiYzEmlABeoT22z57RbSl5MuOD4SgXpqKXE1dFmvtL
GCJnEqDQyxSN0DWoZ/aB1HwZX76ZOhfRCbpeBFAIVbL1M1E9BzsMowlfuMP9t4Ae
OcH1bX+InY9LJKHJjm909y9mnSaONlHRWAc3X+/SuhIO9yFrVpLz+Hb9w9vcWguc
7PJ6+56jczrCS0w5SS9vFZS5Nb/rUVM8pPJprXLfjmQaHWrFxoY7iFRxGTJYGIBj
Rg9CtMwV20xdcdPDcdjW153Wmaw9FgIoY6wKWqapXJTS2QZVvJB9PXXp1ARGiIND
bGzs0Jm/4RnCnG5fLYa2Jn2zcTiE4+5ZtyHtYEdHBqkx7X44TqqHpr4iBvOrG2mx
Y04rJtk6Ca+nOAwjMoRWkQT4mFXR1qWyWwVrTOk8xMoK2SjzdgxPPzh01Bvf9dbP
ptwklkbhcx/ldNAuzaLBYyT5L9WR2L2sCfTnqUvHzEfPvKK9oEVeYUQ2QRbgRBRd
nfNp7EV+hVqnLiDQfQH8MZ7LnqB0GJrJOx8hfoKQ1rFcI2HXy5XbNN4cs0FdWWk2
kvXJB6tvuJW7pzgUJ/INJbW/FOwE6MQbVmb3rCkkHSg/sFnnlErin7/XwlP/2Qys
ujHic6QAfwllVtztywMKOBkMAritFbBKWdfEcppti0iMR9XgqvsrZVhB9Qcb0g5z
jwpk5wHy5bxEeCAfwtSgSREZsFZikMGhPazMNMsKVDysa86a/3PWZ5982qVUHPZA
tNjYeamCxUELGAOPbgy6rSbyJ+BWzurKf/dEOB0Ny48NeUfM2vsTtUGS4Sjsapqx
vMj1rmrTyDMIAO512XMFjSgqPaNgDH48Yf1+QZmmoac6aTwlx+6vCKsO49HzNetj
l4sHmOcg6rqjzTE4DCfJc2vnMs1BJAu2v7J+yAeVE/EwekvJf2RPPTKWLMDVAlFP
B3UtCJ1Pl0v+hrM9fQK3H/oTuNQZwbp3JSHeYd7g0d9dhJnZfOJSdsNJUP05mgdW
fF5xI9L+RztqKnv1VW3WVK6UrBhbEPAUxDd8oa+Q3Rf7llwJqmeIf/za4HAqUMFY
mNaXdXc+HaatBO32M/qjjFxaNMDfuaWfvc137D45OgkBKIYW2VLUt6Ouc2AxM42q
vSCUs8nJrKiq3RJxOltWAWPKpTsZKbsu/X+1+lqezXZEPf7WBx8xB7D06lUNYRN9
2LuSZJnzw0D1Vq/9P1z8mJ9UjiRg+VgnpiE/sa8+ZwgOnMTAyUqKdgf7RNQWAyx/
rwflCYKl85guiALU8IUPgge1gqeOyZExTsXGr+czPkRGOok71h4tLMYJ9NjyMt3q
0yeBqHzp+ViQsLkdqHemoJcdJt9Q0RUq6H1amvAiE+WLvL+LsQa6xUKAnVqfrZUE
LSsCKOxbKJvmsKxdQOoA1h7vQadhI+QsYvJBmTfEBNtR3mpGSFx6cWwnoR0I2fT7
WqCGTeME1Zs4FkaTGKxZshoyUmtgHJpUGbhSUYRzob5GFLRLEcaSAlrRVxqBAiYm
0j0U6+S0Px5wDhgNRd9cXq3JUo5WPvzoCUVcUA8yC2GDThmDzZkHZvAwXj1sTOnA
zoxtaLAEEHf5KXhcDf4o8igzUCh4+JT3LuNMqyEDFyeYKGBaYERZvE7kPar6gl7f
47w04QAfFJpKbzLayxEF0NBg45DMSSumPAscgyCAv7IOTXp63BNTIMrztdMqnZUh
CAShwPheuvE0vXk2FEsOX4S+A0dO2TSomfGwWHdj7evCg4at2gO+ecvKQzPvvocV
RLCC2L8X3TZ0K5/SWSYWUrcRcAQPzVHPQKE6mROqm7bRrqMQDf7UhEzrmqcQ7yvr
f3+UDKvasqIqECypPpfojLII4/nA8HLtYCZvbaFTKNEG0QqSYVjp7xqfyvEbFrnz
gOr384svpUhXpP7ATa04a4OddrkfgTKX2w6Bb9I1hzahZhFNP5kftQHvH/v1TTny
lQOeG1lC4iY78EBKR8dJB3pyCpcLRoZdYhkpyaxrPqZxLXTnGWMB3hzJRE/GdfE7
jdgZMmxsiRfwQUZrS3EDG7anTdEnxFQ44cMJjBPEpTG0KPJEAaRbO1vV+E8zPXWI
CqPyavAgkDq6k7wSsZgXRg/WVhmi8g92/O/oj9EyZqn124brVHuThaUhtFlITy5Y
z5xk+PPmLnbVr+WYHtxz/zlaM0CPaWqO2vO5yCJOTSh14OSqPMgSFjLkCQqoH5kD
9VFuYwHdurCUIARTkY0SBrJscyAG2bQK+IyQt6AbEXqjf0+NkJQxwcrU3m4J8HeP
eJlTkfe/6lkgneKIXjah96zkUsmzev4xjuacY2wanTEj4QnFhvvaBt8ITZeb6ecc
SV8uyurdfTNKAoRewHdtcQDBJWO+/APHQ8387ECjlHzETHJtp5eXJIWgFvlSreUe
vkcbYSwBuNfvXcZto1+S66tzX3KHKK62p7N7oPM5QF4pScgmiWg0I0USWNSgr1cW
qO4NkOmRn50VCAiK7g6SrQsp8xFV/dc2nx2BEjuq25fvEaOqxsrz15V4fYm/i9zA
T6cD48f3nH+AdMJ8zPEH1JQioxxEmp+gXJrgPalLnfswvJdgurcRBk+zXib8rAMs
qr0KJ7vpFAelHX1njGXEI0mfpXh2Fb61V1ju7Qz0IYUGPrQyfEW5feEYBP6vhA7v
/PSDn3IoPDsQnv472WpwGXHMoxMDeOjPB+/vo4Q89ZzP28Mly3io3GQC2XhjwzGD
j5sOreIS2ld9f7Q4KCHwzXly2GsLfwfDoQV1Ryhkb9E730s8ga7pZNq4hc3FfTxg
E6GxB7rWYpu+ltaGL9QVmk34L46ys3mZY7sTkLRjuGB6iM8Lck7QtbJTmS2Xb7n9
X6v/apPB4B/vOZOsSIpvamGsJljh7Z8dbY3Xj0nBhhoGxqffmp4BiGmI7lcZJJm7
4CrAuLuBwd57w6nsjUpAHmAttbozuDCttZVbiQbaReHZjiEKBnJpsTN8Ebf5Zhgq
MGWgjBqZi0fQlT0Rkii9BEK80PKx8LdcIgWaeLGIuMTpXsM4OqtOhIWruXdLhqRT
xaDU8gUKpgFlJNALzd+WetUyKI2nkEvuNs+NsYBJJT4F0vtGFWd7sFz6ynUd7OEO
Po+GBNe3RfFVtCBtuJ8865qrCX3eeyj6e42UMR1T4CRbYvWEtut1TtU8VPjGzZVp
ktm/duUH7MLrpoQgdfmgtzIQZsj//gQdeI2dRU+Vpaz21uU26+5kqtpwpoycJZUX
0rgguPbQ/3ofJSK1j7OwURjbAW2gTYfcXMcTVt+clvP7DP3dTdwXTr/8YgRkUnCQ
7fqb3ysHY2AXMbm/b0mDV5Eb7dgf+H5UBRSzeTY2SVfMob5OOYiBjQqW8NQaN5bq
njwt6vaVsv/Gsab8yect/OcCRs388c7kBwIca+9a5EtVGR9BOhmdmrsKNkzfHZo6
BoSPEkV9eviYi83/KswlKbXJf+CXJL2aUAJaGx3OGYI9bvQQQCXITFUcrQpxbY0G
88h9fE2jdXCf0skpV8PIk7X+8dd4WTC03NpMB3Rs+wlDkpcAyBm81ZRmFapk+y7A
fbtehfBR/q1+eXdUdzcyilzDGBzXRW8oTbyKqtyw86OB64WBoP0e+9MjHcj4aCNB
R+/VMnwWekfffH8osNwgf0kYy4fjxShTm+vdvQ3tOQRLhHtVbCPoFVpw/2wNKCWY
Dh9IPrB/aR5oWKsJh9DjaCOysHIxgcHI19JdvUYF89ezChpNSvbSiJ7ubrECJV3k
RUG2pAtay6RToz6hvWjFFR33+Oc4AVRcBGE4ndY0nSZmemGNpo6N9zz1XaZsiUsh
HWXRV+wQCuqEpjXJ8jw/a4HoBRTnwZNgJSX6e8m+tFXdGDfIKf43jqJpq2ydfDnc
TUWOtqW8dk2c9lXhwVw8SOSGyD7nK7qQJ02Tg0PmcMl5NFcqpzp8k6ycsThVNpdA
OzAbZlwvWLTX/mLJiEVfqVU2PjW6OPNDkTpZjcXwHYMNWCWuAGvNVxaCMRH0+bu1
Pky70gNXybdxeCuj6xn3DDayzCN5qvzANSsHC7YPzhOAqt0Mno8kvTTvr5HQQsLq
mGDrdsKI90DLETIN3BKgRmNH1FQANnZHYkfQrjIWiFpP28wl8Nq1zm2DkKEoFq+6
8zKrhbDXzmxm14wYP+8dfx2oMUVott34orvmn3TbzXDlxKwnVja3RMLDip9q9Xcl
nv2vpsWp+tzyJlT2AmV6XptPiox/v9HQo15jdAxjhnPqKgcmZdxy+D41qSIkhh3y
Z4WfOGI2JYo0iNhJG7az3VEUBX1c3upb4QTzAClKhkYeX//Of9XbwzsUGS0L+ye+
x75jAMhWO0NCNskUp8YG3t1Hk8teaT1Y3AyS18X9B2BcYzeRU9PFKVjuLVlg/XhK
MkiLe50C41X9koqv0gm/6a398B9hSxyB6S3MHxTub9XcX4cp2oGUYpwic5bUqwIe
Cq1EySbl60AArQyTiGTNqIdzSeBcIlr5QTq7DsSsmjpCLgcsY0qaCvJmq3XhhxX3
FKR6A9zhv05f4qOIiHF62HxFpuJ91Zz8e8yLHGvn0po39p10vGTR3MnOPA5zBLSM
DxVE19iJrQ513Vh/Bm9pYOJK+gaWmoyDGDkDAhfBTethr+BJDEdUdCMs2jN8NLe6
kaotsdg6+fi41APJN+v34SUdI/Yjz3WxWRsOEceesGerYhTO1Xg6fLeubFxhZm3R
bJ5XXFbXZF9RRjZLxVcHNWAlrSuryXCfCe4tN3LuAm6gtXT8UKKc8q5+bozU4RBj
/9gfjlJTZfMEHrdPPoVPpRyGBc+vkyH6JB74q3C3A2Egd618JN4nHAXr1OBSr5Li
51wg6KNMqE4AhKv3M48z1mvO3g8BNV0Gt0B/RZpvRpTJx7WEe2gAbbfDavXmw9DJ
3oC1Hpm/WPJplJwI2T7gM8GMXatK+KaKk09sraW32SRSf4hcJ6U/OoD0MwxNgF7+
B0mM+RTL+dVGscpmSOdaOezuvMM1wFqYwnmWHL7A/uiocjjRZ8QmTNNWn9UD+SjE
ZSfd6Oav2mQp90jo3tDUozcz8/39BU6s5hBZ3D8hCeGcafx/XCPlK49xAz6jBLps
cejCnPnkFDpqNUQ7dGA7xqqFyEIt8vu5rfYQi/vMU3YSGdpTru694TgXhTAdh8nX
ti5XfbrlI+d/KIZHNp4RTgizrDw+IklR9/U4AxRbCzKSXbve48jH3Jd87F043dM6
8FasAsgcGUTcAoIRZZf+Jl1zTFNZc6wsKDEJUEl9dtwylfaJO3vs3rYQoQeygJ2i
p3NEcqref3xs00o9hviwOaercTate81ZLT3L6B0lX067UH/2vYfmOlSJT9oIlUDL
2fAiIZ6DfiDfnbGBRVOxQLmhg2YUhJv7feSZYAguvbxnK35eoD/vb2B7XgZY4Ckn
PYSlGys9Bh/NWWZt5Ie543p+ODAbxWsHL+6FzweJko6f6MmAs/HkR36dtxTbR5ow
p+F1ikYGUnZwIvIwHVmMtz1Exp8A+TiAYqbk+5vWo7hPIi0D11ghI3wmJj+2Yc2j
qu7DUoknAE9dV2vDSntkCNPi7LFvrEWaP9tAu5RvuZTOZZDusSq+HPTxTJhayPX1
7pH3dMyojpUcOSx1BHWtd08NqjUVeR+FdnoqeeGyImHpfbu/ahtrDXys3JMBsfby
wnQR8A3XxM9d1KmU0Wq53/ALPjRsVGBAr9mFBFKSwfYjsBKBVWNO+8BKDOTX/0zb
hi7wg8xdAJF3u1fsZ7j9dHkiZu4fI1kgzoFmK07aoAZT7H558SiPMUSPcgpbCDol
VoVHijZVwDK0WZZhYFbXnw+mxpMAahLL6DC+f1K1Yg8wI7r6Dl/0nUq0gEdMEgKD
rT1cpkzHEA5Bp1JU3hG2LFNScvQ83NNX7ukhDhsUx5CYAqFTYEbgF7c8p5g3ajA1
hA1+96yZGLMgcysx7BOtrGLfPIlcU6hIT8tcBciK8pDS5iL13SEVth6GVqVuped3
ivcnMrShvVsP/TIMxtqMdN8W5bKK3cRc5bdAFmbRPihsFDe0FWezK9SVhr4XDzPO
UVy1T+4I8uHPU9pIpx275clnsZLvQbfcj5Yeqlji9syMz8PsT0q2h9F6E4j+M3IS
io8M+62cx1nfd/wtvptep7hwKk3Pt2Z6MSmqjspp6X9Ueqw+HmUmYrIJaEpTaOuB
GlSgohEa79Rjwr//K28PicBIfwppqUVrWfgllc1zg8y4dl2eUIGNG7gg0hkDHqFf
Sl/Tfo45p3nAKSxxfrbwOoTYU+h6/SUnyCxatQv1TolpY+RPrGNFn24BT2Umpefh
CZx3RHVO3q+VrFsxSY/ssEMywm8bHFAJX7n/TkLK0iEkUjzV0RiiAiuGrCKaZHxk
VH6z+J+gMm01YYXNpC03Ly+4XAeVYrMhe2wGT0EjOmAICuvsYKjKjaDx76BqjrQP
PJF2HxdpTq6OONzWClAkxlgGjyL40n1AqWa7uYg5SSlC1/LL/vGutpSs4VLyUZUU
eqZ1qw36rRzIGs89ITJCotSM0UJsR5ez01EuJ+jjljgPxC+5U6Dy3V9Paiu9obMc
j5wupg1ixR1I2IZFx+yX3zhk4D2XEQ0wE6a+M0lDyh68iyqfd9ukDRBxq8IxjAqX
jhVsIlr72DGlZ6BSZUL/urUQTTZr8aQsBFdKkMdRcp4RbFvnkf6qe6xwlSq3GdYL
XeWClq1wMAWEdwnjV4wtU2vnhM+0VjD3Au89aOZxTQr7zWd3NZSWR0pvXb9uNzaP
I517MYPTiIaDonw5o9oIXdV/ib0H2YYiiU55R9OOnhDzKEklSs/xoKE8qx7RwR3S
jlMp+UP2BQ6bHWtIP/U+9OqbCs2b6rdge/0dXwrIKKKMC1LbmCtPp0tQc9Sutgc8
0p2C6rirUDhwqgnbSjeeHT1zljE9EazvxacvR2WtUezXU3AeZ1R2u1ANfbvldUr7
j3sW8JolPSo8O0dxNskN9Cw+PjF2LSpac2kOnv7gBeEsM5uKBFgt/JMJ6No+2IaQ
vbojuzcSvSkDV1s/esuI76d0vSMJ1Cds1f4eT2W1p31V/UX4O8i1gdkiipBpgJqw
JdZETXjlLyINeVBHvBecQy90QqfgEKAZUI17qaKATWDFsj142lXhPnAOyef0DcbD
flt7O3GCd/QrQRGooSQpMlxBAxlDja84D5ZLCy7UwU7BNLSPCAexJ89h3ESS+8Fv
8DrdtkQ57+quApZr5LS7+HxZRPP1ogVOGKxmDPW0hOCDLj6HQjlJgtTYPtgHGiBL
bf4tJp5Bvj25SjeUhC9KEHWQ9+IuUY1PYSUtUl8hGNzefFED8XuRbKEUDsht8EHY
Xd6W5ZTOGjRiKDXn/VEFvZN1Lyc4NHb6EwuuPSg5TBg4Au6Hgy/13WGBe/8xRjNy
WeYvbEPfWB7HJXikLvk2cf9Ez3A4+aPHgoiiYD6t3/Wo4G693mTz1ibjbvFbtSb8
ibaxxeTjf64lg7e8xBYwSrNxvRz8MK7bqdoWeGrMo85gR5vafNU8DkPYHJHmH2W5
Tps9pYJaZh/7MVAFdjPsQ8seGd6m338tQiteZNVGxEKnWCrXoPMw6CQCffdCJiFa
1fIVV07xjVp6qzRHYLXBuXT8C2dHAR2IkQ0nq8zloQGg/OtBOpL7zydSdbwvQbMv
/cy4zb9UrRy8D5ufJjQFOKTceXwtDXOeF5CiTite+KkKBvEE+mMNCnDtVdbNIlbB
ZSoY+qTWfA9MSxpan9w1i6gF1s0yjSucE816OgcB2MP+hfYt1YN7tU/C52+X/PSd
02Dcd/q7cKNKz+2cl4InYrhE1fgywLmCRxkY2/ZpnpQYRL9MzY1YmA8retYwDzHC
qKPxaSYiY9gfsfMqZhc+MgrLijrr3JHdPfGilcsoncQNixt0r44PZ5+wKyDePmg4
/4r9OJoJ3jYi7erK5FKNTY1KlI8IXCmy75XKHdoZf8KKYnuEPfLL+9OPb/sZ81jl
Uo5ynpmw0YvXPZGSLKJay7+nW4QGdDbV1611lL4aF9UCIU1X7XGWIipc9cLbN95N
4Sf2xVkjlRXJv9WylH9Om8RYWrmRgXGnoIy9KSxFsewNhPeDQNHATGXFZ5NfznZz
krFHtkwI6ZiHf+ivdv2OMrolxz5/6go8SEID3MbhPVwOpQWZWGsWwBjFQrk4gFXq
XUvsruQUIHkjqN3FvBu6HXjy4p1pXM17nBX08YqEgK+WhiEu0yt9OmZKwiNyn59O
nen/K3iUwI5k+9IsVNNYNPhgdv+T34BtLUJnfIIEM7sGV0CkmrKpAlploo71SLv+
8zL5XzpNOC3m8DQf4yRdciEe4RtzRXbTyH4hb8AcW5jZoOKxuG6Ss7F+zVprtAFu
UlE9+qGqZonK5iPOMJljvcTew6WqNpDbUv6O2SaEYWgl1iwAPnirPexW0K7kiQRt
JfVSiH66YB2Buh4fw7HVNvbsG7BM3eDxsRFlyxMHRs9pKp74rh/fmthkD11YxSYN
ARor8T6HK/Qmv0QPLaE/tzLNBXD9669am0bcf8OaCNWHo9UoVCm9jqDp2JsRkfdU
SCMcqtVWpNpPdbqq9cXRcT5ibNlwU7D4v6TfS/uqZAiPH7mBnwGkpMuCvfcX93AE
DE1zbLXFP5VC7zlHAaCAEGn37uzU9en8mQwZSmVKAdovm2NUmrxUEHsmvHYE0t5+
oYhbGoDxDy1E4EIAoFzsxlKnHY5D3nRx+ZhIMXbdExam5rQDHRETJnUoxkNIhMKo
g8nL8u049gFDKRG5mP9md2MGnLhf3ksGMEMZCyAHj4143YwbfK3KqHxxA1SBOQmP
RvhGiA9R6G3QeTIlBJzDj+IZ7WwlRIhM/WoB4BwXxap1imBg+HEB15mzMEEChyoW
fPgiHUqeeiHhm+rvmWEEt82aWtIl6QqFicJVgcQAykMSdIH9yjRKEaUMcfdfuUTk
sFg2en92rdTnc+zQ6QQHnMxhppKnMdTtsQ+OiQ6iR3Fj9sw9LlLX7Hk1wOxeyd8D
wRiQhrfPRmzpBeLCdRr+Fo48UFQQErAqNeVmlTrOtY7rQ1mzPbXtyedbbgwPUMx9
8EhUs3Wz9xOE9obfd2pXiuXes8Bjk+vTFlR16apQEXJ/UI5UtPizYrPrMS1o0c75
TB04SglLLU2f/8dIWf+4zuLcrGvCddIHJ8ZVM85HxQpHJMJsc+PY0WMvf1BA1ZNv
bb5S9SLBAeSzGun52wcSZfYvntdYkMkI4K+c9UAd0lEkntYt5HfZvNzxrjkOyu/x
OfkZA0O+BGUjoLwjvDE4BVErqXnBggFmtSCjqhR00zuX2HNryR6WKbpjlf7Bb0Lm
Ckwk1vhWBRd/PHa8mGClRHo6YkioKj6d24xQFtTl6ika5JtAfDA7jXjE5WN/mHX8
RgGvE+3hpBS0cO48RlkRso7+JTs4MuTAfS1AgrKrKDLd1ozSmq/wYDUrQpwCbJoE
UNgWGQxaLqRZQ/KCZhTMeas+jx5SfyB88VxsMn3CDG+k6mS3M3/htfPg6SFftdAY
uRuQXb0P1+KF+7ie6dzNlKe3qpPrAtcfZTJY+Vn9njwSOKgU6A28HexV/6p4AyiP
G7W0HrY//nR236z1rPBixxed/JCF5JxErhsVz0rwPeCALGcZ8q+OP/DDWUCPbb4b
ZQOgOeOA4AlUNeRhOW7Yqz98SFYXEaOJttH38xzwGazHINx0KzIULHgwJaz6wGip
w2EjTyxDPzqu0XeP5HMSNKGEHOEiSkB4MlI/3DwTUGM50GU3omb7KwjjUsY/hh6e
U02mcgQnKziVtKmQxXp0uLRal7a+rdKgb5B0umo0d+RTHDIUA4wn6WKDsfpGNYFw
hXB6hZ3H3GU8GUReed3XakOAOmR2/5dW++XWLHzeDYWWbc+zT4Ooy8eHyPQlC8ix
tJiDVTuN9ZDfOmu23TQvV5d/WsasJy1urI92x6WZscKU+2bRFZ3Qc+4qDIKw0I3w
dGgIA/oU2PG/fU2/ZEPz6IUzG7TXOUnEeuVVKc+kHMhbigqRkTmzDxcyiOJltUcH
G/NNpmx6i/IAwo3AF3qOrga/6N3CWwvS5071IWy1JXdjAQdQi/LwJkQZxJNfjWx6
KSblN7WVLLavioSHYs8qPM+JieNxTZOgPu/gEUYARdqmbWRigXJtCr47//BXBiGp
V3UpT+5/svyV0O5UQaq729efgHwxCFSdHgpr+Yr0fYFjANmi2L3198UNy1sBLFmT
T3PylyAQNaON5Z98+UFnve5ehZAE+z7BgI5obic8ECQ+c9gQAVg2J4jCPpRSYKGA
D+EA0XXS/f0OPh4QdJOeEKjmgnyXNORQbVKed+1SAQOhng8TE3JABfOZ3k/gt3ak
CvcXwv95Rlfdd0ew4z0O3M0sOVThm0gb5UagmRH40HucfXdSctWVUX//WT6AXk7q
wPKwLWS8mE3OlPD/K0npZUtzC0UGbv6mAbeBH1jxBiZ7M5+NNdr2qT0eNkmHiIIi
176DjkcQZ+sISY/H/QZBIv55mcUVi7Qoux5VWKKlqdptR3kVYLbeJJNalyXRMcJ6
E6XsFpxB7FeLiBJnA9RlazdkEc5qUpelaC9+kVvBB23jJb9YKqulejid9tKBi1gt
CT8ZBCKhDzr0szJ73JRRrH2zW6CXTklRDQsheniMHbZrpFG6dxotQ94bL+YlkOEs
G7RRtrHXH5Zl2wtQID8Y8PK92SgbRDU3IGjKHikJvQDoM9fBhwxjaZTykbGGrr8K
B4vEGyj8gFS0eOJr3cL28im3YTHzGC8Pz9jUF9m9ePOgcK50Q6G80te0CRhsidkd
lq/IVKfXiXoAxztDd4IbkfKWDP8hdhLlkAY11l6jSIX8Efm9z0kTNeZisHCE2PKx
RncOTPnvrojzuZkgLznRKSeUGBwzQLV+OjA15GeuuHGXQrEQgWUDjUVu2H/diINI
Qqoco3a11kdVEGNm3kvYDi2AZgiqsl29zCjzpKUT5zABramMeeQHSelttmL+HtyD
+hbfENVlTFGp5d8NiKkFiD72fpzPC5o17FnC7hVvS2DG0DW3XOx4wRhd+ptibhKZ
QXyUOBtvi3wEjLduE/DP5wdYsODW92GWGdkMmknwX9er1ll1yaTXl0oqD59hPF6o
AzbFbPmLuSB21BXsfDteQdAoIeQnBc5ncczCmndnwPvf6Z9UOuggNItxWZbqWoXh
otws2CvnzQup0X7/oc4s0xESuazIMN/YmXL8L09ZC+GNfDNPUY69sPV0Fc9KSPAb
C7+aCfWAIKBafFWmGtDQSp0nZ8c7AmidBdrQEfyFIaPHwH6Orzc1rHiEwJq7jSDh
RoiYjIcWKeQ445dwFkNLTdYj5kIb/gQyjlPWOlIy8tijH/a8MJEW1pPUMPP8mwXz
IAFQMGlWUTUSa30z9EmeZZijYHsWLLtq2IepbijbUnxq3B4HYXRO/QDmYSusTklj
YjXeSVg2uNKiQAOytLgw8OtfPVfI4VXr2xhWLe/UxLyvcmREH9KYHZTRainReB+V
ivbJ3OJJY5Spo+xBcCupLUHLjSyJaH6iKwoKIojOSMPMK4x6BGoGK2/PMRABSdS8
3kB6xYHLYlvhRiCShK5M1nkNrX4GQcT2N9pRRse0gNsp8gvwxxaO28koagMN3+Fi
uoq4GSQRN8lPAQI85tdPundY1o1+1yp/MptH9Ng2/EyUiWJzeP1s+moXfBVloC06
H5ZF2oU2S6XYvejO3fVYBlVtw0H7E6wIqd8sVTz4hhRsVldCgvZ8vN8BxUgICJGg
atsxC5p7jJQasvk1r+zasavVxKS7UqdWSaxIioZSM+63yIkSGabiBWgPOCE2I/B7
jtNV22x6y5tmeejpiBX5u6AgjBeCCFI0Cxi42zUMszxl4oaMdRKDGuSb9gcLo4x0
+AbSeptYkCyRwHyOxW/GdO7SD3HbvgIoBVeFkLa3hpN5lZQEnz0nVctMcQpqYqdu
EUiFT+VOALT2n9TnX5tluX/y1qMHuLnERPjp09HrGj6tDkbMmDQjglYqxJbctCZi
y9ImXOgepBNm5jM70w8Qz+wi/hY+wSI3+ZOblYGo6ZqI1/J2IJfEbXFUvlGHnMBy
M6qQAAwNNxT+KgAFCb0GsF1TfWDwoZIxUtTjm+8ywjCrMOApc427IDFnoPOtyTbe
O+Veg1Z7U3uCCJfoMNeGJDwU/sO2PXQW7BS73950VlwkOGq2IO6TfeEm7IW6bb8A
yccXf8zJp1x4OEQADnDkwhGbG5YpIFFwwDeFsbZQrS2AlwPfQz4gCRNnxN974bIl
hTHxWy8fb/J20XyGuxYYcxFMIO+EWzFJJWAgJfm8MKM0A5Q4zXJSi/zGs7yboONS
YVG46gipuaskm0Q6ib9td5EUInUEG2SzmTwk66djLTep98doG67Uv9ot4WlSyvWG
vX71+UYiBBw2FHG+XjD0es7TAqKyvraV/CwekeZ3JNWMt+o7R9i8frf6nfunauU7
JzPrxmXApgAmCezYtFfoTVyVQVFN3gl8MG+ZNI4EXOunkZe3Z1DVftp0kTvCeOm7
q/TIknLKWjJBGBBKTObiVT5Sec1wTz7MPN/HrgOcsHOV96hLU00wGHqrAUyOJGsk
F8zVWZDfmt/1a2KwOwoZacilQacbTfJl2DPnxFlJYF6yuqZDy83OB5pcMhkxRqXp
zZDIAnoMR2veAscKcqr57aJZ6LoJDSVMhQV09poF72Nob4xhoXR4qcprcHmjjRvI
V4nDA6h3wrRRIH69PCQHi3rXUJqHaVinLHwTUwE+wYP7XbNfdljZZZd9KslbraUJ
FONe9hLcjg7mGKqHRcgt+STWwTQ++3y2uUNuxbQ6pGk19x7UXQl68EyM86vWOrv+
pCI/Bkfr8acdbZIPz7nR+z8v1DXFA51sTu1wvNInk1GSctd24x2jW0VhAZjctp/B
qOTKIt1hZR32wuUP15We8BMlFmv1Gw+AJsWoNUqtYSfhjKs5Vf3YmcIH4gwZ2SuC
mWBkH9b3ERx8MxvYxNcOBIDZaYYhJp6vlqkUMlUKc7etA02dMRnqzHdkoFweL0Ya
1sNKElJ6Xmv29U7YcurJBuvF80W3bnnl1C/hRp8NHyie41xZjGZJ5W9LuFrNL2lu
/WPQvcwH3LDZGxGdqfCky9X8PWSfZihhgSByC1bc/m/SLJFV8jIBjobLy2ipDSI1
xiCRMhfo1SLJXmSr/w2BECzBIZE4BjTVGiIyN0svg1IZuxPvs/pVZNahIjnBzgqW
OdmsbuDjh2YZLySjyLssNMHlJn/HWWVAt/ztbQNczv7b67LVaKpTSACBk61HZHtp
jo0Lonon/hdXuRvKJJYstQAgW0aip5iQYiwDC4UubNdufModbJ8lNzdaP0fEQ9Ky
uKeY+FzNA0xpRMfE9cfoM5TgxNQHtkbM9pEHNb+R0ch3TN6AFJTu1B/X8PvDnz8e
0psCq6s3tZYZY8QwxQTXl43Vwx8YKC3q84eWmt3D0As7dLei9jFC9Xc/hoKl07MI
wyu/vSV97syOpmkUTHxv+nUbqBt2FheGh1/JlDipWQ/uwIFYw1J+UvNM54t0Asqk
5BdWilYLGOgLgYckEe4JaLrONaE6vlstIZ77QCyhGPKWJI1kAiYbpKY34GFVpjgU
HAxiOHLIawmUIEQvQsy3S90SZp4vZ1zQtz8OPVm7V1K8sNR/Q8CtS7G+c6dT+ojf
7C2ojzQSOp+E/YSopHyQEQCMdEITrjsrt6Vt0YTmrHj66oADRU40mhJ+9oKGtaKB
VrpMFe9pW3P97zz8iyjRwIGgtuvkE21wVBfG9LpU3Ea15VmB1lvJIK4INORvSdnv
7LmS7NZ2au9jBqmvVlDL3wCYJKMsqRnY++tLziy1axyO7uy/wjLQ7hmigVwtvA7y
i6KXJs1IK2xMtAQ4F2vl/xMlWNBDCWZ4ZwGDodO3sQZwmgz4QMcKgyxpT2/d+FBG
FKJk2QiXjZixXvFd+ELZFxf1jKvYD0SdI+ngEaRPGKvGyk6ue9/lsh41DA+9Vc3n
f/RD5MH+jDb67x5cqOJL5Sr4xs8Z4gUFwm7xTKYysJscb9BSq4qNJxL/HU5mRZbo
QRgWSMnMRfAZopOLXIdJepTv3yw5ivvP775pUy7mqktfA+PmKS3UCIKXJnNVw0Bb
vCiZzM2g3hOy0BDvJtri0uHlFSrIvFdhhsZwtaRZkkcjmVj310lE7oQyUnaKZ+tp
8FrexDBUJdaOn8eXitRl9Xs8cNFQFdBCr4qoROUoXL7wRwfnkugF+HvBjecmleRp
HjXIXl++Q9XTs/7pjTcGY6kLT/VqJshGe1n2jsX7xamZnySpbbRnBKXjPEArQ9eS
p6AkCFwrqr/uDVb32dCK0pseaFCXFvcz3xaqmONTf3ts4BKXQk7p08FIEBeSsJP9
DgSHO8RgJlzlrI/AUvSU0A7PJRgwJ7PajP6qDb88TteNJwv5pIKVUAbp8IrSVYWI
EeJce0zxlg8oJpKydIX/yMrMCF1rcl7VndgPcjBXsfC1hEcfzi+KQFs7MyO8Ikxm
uSRUGerkDV8Q1O38g27/2C/trdo8LH3IjF95MtIniMTuLyOFLq2Cr0JPKSMKSS0d
vQxLoMhpIa+fsGO8dcOstRgvS99ISc1xB5YKv1xs4vG0cFmxt9Zr6QVnMul7niOH
e+Q+/eJdnTdf86MSi02by256FE6rudLxT1iOpqqFk8gZ4VQmDK2vsRTnsWNNSweX
QAUxPyezd2ExZE/4aNGRc/KJ5nAb7zywBKEYdUF2LaVaOKabmVS1V4jUHVxK11kz
j9Vnp/tzqhrLvSc5PrQRc8DCq25M40EuzWFQp+nZ2SLlxAnumQz2jfu/DJNn1MQu
hUxa43R6oTQBjzOI/W8TICQvfr2ZscbQfm45ZE8mx0FfMCCt2zWFVxqENOHd/Fsv
zTL7zJWP1nIstfhpJEsUiMsrGIJZlCwNKzFB9wIpsDYekLnIdLJ3rEQvCtSaVq72
kAtdN957ggwixzNUjjREo12VX1HgYN2eLS2Ay+EDiSiqSWSzofCBm68v7nrFMkuh
YI+QbJMMdbFvPEuW2kQLVg==
`protect end_protected