`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15696 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
kXyB7gH0o3qEH5aFixO3viKxTSl1kV0FgZ90Jct6sdvegHDaLU326pnrIuVvcikZ
Yk6jpUwVIcZv+7UVh9mYAXNMBH/SP5RHslGJECTJyKI0OU01M6b24qqN9O7Zbjw9
n318oLVCc2NfUY6epmCm/22zB3/e2e9WgXQTmQPTnlZPsUqaK2+Kn31u1Dc8Rb/f
q8H+CR+WlbKyJinDCe4NUsq0Hs35WLh4KzukIYtqTvmejBlrPj9JfMo8dS30qZjV
HCdI/rdVvgdILxWTM9hmNPUMEEHvx3/4HalRpi0cJRSJNxGB+VOYgHDEhPAy7Dk8
LmWNzrrPRaclDCX63XEOUiFcddQY6Aimf7z5eN0lspsGD7gCZUVsbJErn5/+fft+
zbmj6Drr0xLkbN8mmNORaiA8+NH56TVNqXYdHGAJyzPvn2nSqej/8ZoR8NOh6lG/
40jSQTYyE+TTEhmBRP0qBc3r5O0+8sGHBE5keyRoQY1IruqyOSdmknhM/vnxUAVS
WDEUXsdyLAw8TFQGBHHR8jaJZ7QG980yizB2UxLOytHq56cb0L71SE8yLP6wygRF
4ARdraZIXJOCu48vUzYiOwNHUzMjrJDEK+Xtb/GNqH9KLVzZJJZUZTFjescQKuYJ
e/eSBrKfMreGZn6y74G3z2FpSn709ZRLKtQtInZoHwn0SjAZyRuGhkraJ7rhGNKf
m4vdcLOPzwsVmwOsAlqQpO7LqguLvpRv5iV8HSvS269dpKRfnlZQXRnmGTuYk4cD
sw3eVbX3zrDb3MN2zgdSJr1m3x70u8fGgFDWNm8/JyRm+9A+3yzJ3xUQYyWtp/Rs
Q0bR4d3j11v2F4zUZqnyGVJW2502fIgiJ49rSi9lb2BzuZ9oG1kZFZDys1an4t5P
HYb/s4C4wG1hQnIjIRAvfk0A9lG6EZEerlnhsmeqQJ29ZEip0GmMAGrrtvwPFsyv
/HRt0SxeJnU9R9qfYpYpeFOxsB+/B9but56RsIaB5vnfTMVnnY9ujk7NQsMkkXJJ
d1K/LIUOus7FtUfzA4N/Z4bWsxg403nItBjDVrXfZxRTepTOuZhiU1yFl7xR4fgW
zFx4I6B8hi1IYk3RgBbwqPP2oAfsgWCnWWf0Y2kfFbr7U000UaaNzs1XeE5iqPVh
n5VNpZclKal+qXOTen7gjGLTN5IFDINHu3l4yJH0tgnz23wmWikZwjFUCWT9Qphn
NggBCCIKEx1I8rRXWsx4Vd7CM53uqXGx9KtZQAGRVFWcBFgMi/pBy+BR0iaTGmCI
3DIm36ew5IV9RRUWWcEmLC7QifnIz/hbLvZLn7rig+30/hpYetNmpruvqprLG4l4
Rn5vunvBt0xpk/61X0WZxyM8X3r3xXVmrTz7dpZm2oAKa+Ug4jBjz/Vy+9jnoyJM
60eGmkwJGUfYdSUeGCw8xdNeejSlN+/P4LSXLDD0qPR5Sae0JftoQsByu+0WSjXu
vm5B8lOTHpoK7iupcAVH6asCxMWmytnSwR7BysGzCp0lPqSxlPmq/S3pEcm4+JG9
X2+HCDJSqbnfvvptNFu67d0vFBNMOp/fogg6ueEIC/PtwETBHGJF2DxcncmDlLjK
bv1aQSNn1L6D4JZ7b2YU+CUA3rYVNV0NkTJ7wWHM+2OVY5LCO7f15tRb0ODQGOPV
1WcCN+0rmwPb8A28F/YdR48AXyne7mZEhG2BI12OMbGNTeuZGce2vf/5dh4BydOt
twIZenNHcGp5YlYOugRiTaeNCfqAqEt0Bc7Fx20doluNgh8p/71uiEiRbsFNHs49
VKuqSAfe7fupgntbgCbGJV47M1zYZGmIdAmV1wh7VXMubO8Qkz8SNjEnejdIs7tu
6hLy6slnc4sLmujUu8/+SFDfTZL0V+0l/AHnAz2yGD7NWJWC6Dut7DR6qANUR9Z6
Nd0zaScTq5N9IBie+40xUz3OxPnQnSMB1O2mSnxg+XJM0KfBP6mwDESUn75NNDGf
oL/Uvy+qw0hDd8U3lNdCCvK7Z4N7Jm9fT1YpsV/CjcSFuhNQjGv1KIcUmf+ElI+/
L/Y3e1lBF9zspI/xcWOj1mU2whqZJjsAEMfMUk5ie9H9+Evd15xqOjcUrTVa9Cbt
4T6WkEBBKmzk9WSVmx+fy3TEhnCvAb4OrSkt86esCruHBJLlzBKvzR/CkgHmQglk
iVHsDOyVSpEYMT0k0TOu/zNeLVdfdoZCxVgQCZY+RbpDYhuQGX4Re5Dfe7iHxtQr
R+zE5Sdbep0t4gHYrFdBYC9oAd96AFSDINscRAcEivkUX9R/ln2BKKHfU8r7Yjca
LdwSd0j5gl1sT1PHGVKTo1DmmVxTrETFtFvbFK62tsa5ZYimfH4BUzePPn5oXyt5
ybGZ3EJwPYOCAJKXMOTzVHI8E2BtPQyJTmbDs1tLAENOvnuEYrBuTXR9/h5I1gBd
0jXy9fn4ZOzhtaXsgBkg197Iyfe+GzpUwG/9+/WVqMWwsYeKcnTyO0PSblWKrYGP
GLmc2ReoddITCyeiNnpMTLnM86agj1fuFUyMHPNY52xv8MhEoqDltA2pJ0/vmO0O
Kbg8ZVBgXz0bTI80svi7SeTPmVNZGgQHnRV7s+Vi4oSGanvDinG6QpNLYUjO7bk3
OZOKxn16Ow6K1KCtstBOEefyel4E3Aklzvov+3Jn30/SxsB+YuFYV1OsdW8clGSw
ME4pvpzhpRn4m/rubBf/2rbXqD4LJmMbZm8HTCQ81T0s8GnSsG+FdN/gZ+SY3Urg
RZAj1ouK/t7dL4JIqnzKDDqrKelPFYZ9gOxze8OH41tQh5IzK18UG4wgQxL1Akir
q4uf7afpzTR8js8kpX4Wf0h2X/W9K2t2RoEYHvqQbQSYxJj63Et31rs0U8st0PH1
pnMz6q/O6EGauyZrTtlP33GG0gYadQolDJNIMPgE6mTO0ZbosUYEzDxr7MlVR+0F
i8pKACrz8WMeI7lIY4Btxnwy9PAzl+JpDvitBo+1Q/VJy1oM8QVqvs6eqC4jhi4C
ZFt4r0RDAQv9b85UK2mpI51hmadyT5g+cK+dAbuGv6iGzDxG6Cw/qbGp76PAzbxa
wO26Nz/ZJy1zbXj3e+K5/RQF6OjP6YLvrEhLH1pz1dfucD6h1huY7V7adjz7FddJ
y8+MMVxgVc/hIlNfcnKU5xoZqodUH9y//QHe+ckssWdwTWdQhmbWBXOoCbUYl6td
yoYeGiwai73gA+R/0gdAV9lXI5n4Na5nKrH+ZimPZxP8PMYs5g44pV5RsOSAcanV
SH4TQLtRP/tQiIxJfSn3O0mVQaO4bjuM3lLgjtZ7y6/ZG92KG0us+DT2LSpVL7OH
CF389BAS62mIXo9jE3jr4n5Ay3ILMS4ogpRxBQKYApaok+T9FAquzsjeAAx4oRVj
wmdIjoGae4tI7F+/bj4Yp2odYQtngrGHFdXT4/l9pEkn+Mk1Qi8BHqw6dz+O/umx
JKzP7X+iUpS5JNui5n8oWk9x9cKGg5BdaQ5Q/vR0q9AuUnsbKH2Ck5StItVHlAJ4
tP8bHFh9qXL2tfxcmtDh1xbIwXjbotHx4s1NejuYg4eBNY0zKeg2VwSTBorVK34t
H345rJVZiyfMG3ZrX1z6IwDMlqNpACtGqoh7C2oPoPIS48Bnsl2Dqw575mKp6Gov
USDVcxi2SK5gUGCLJe5S7O7RqeJzlmTUNfW5TJ9WSNpR2T3ITK3oMsbIUa9dDY9N
nsteT6P60a+s3z5KsGIdBjv5scMIs1jod2/5Q1u7Z3NziImASoI1e+WhkntgY2PB
MJw3D+w9gPkwwj6Ys3M6Eh9HJ2PpEUYGLFarU5UutNOImwt+LjSmbdoXiC1TF269
n64ngbkLeak1NlKGrOwMvyvhX1ik6CXr5cJDgmRm2K6khH0eOlVz7JvV5xHiV89W
FfDT5ajViz139tYb4+dPxWQG76qlk25EMy8dVrwomUtkkH633Jp0W1qUQKCkueAK
YrKZTsLOCmTOGaWHBOg8tnGuRD++pLaDZ0pcCIa0UyrLqjyUw6/dExLzLtqRruE5
O91+53pmah7ALmj7r6NewWLjAmvXC5tZeQmHIuBHKMtDGa2kP/ohIy58KdIfHp7q
wMTlDimS6nM5O/71F5QSu787Zs4ZdAQxlIruGWxpXGjAxyoUBdMKoI52fvVaRoo0
jENTW+3OLknhlkCDQxh6QrYYns4AOo8HJqKsuOXyKsOMey3tWaAQoEX91rUxXlsy
KndnmOgHlWJNqH6m/BnwPGvDymNTICvqkwkE8wASrUFP26m1ErBzQVErbXL6fsAF
CF7FtbflhFvhNkpOGAhOjZvbTiNs7JzZsQqCcWzXgwKpVF8W3JStv4pBqZV6NDxc
aWUIni+FsCaMWtDgy0LV3YcM+9QBaKpA/ufxsSQ2Duh9bSXxGtqEPrfQCYq4VzW6
0SwAWKSYplVs1tLlNSlOl1hPt6g02wJ4dgvSjtFlFEW3omHPuuBKkYa7MacEZctn
u/k2Osx3sNfaOP8S8U+w98DRF6y2+elxIw54gjHgt1wMfFuJJ25tnm4PFeUi52Y2
DhO7/jOD75RDa6Hwt3qTx5b9xrqEL7Gv25OxsmEFQLOs3HmzDGgZ9FNEjkdZNnuJ
i/vElvyK/QDZTH7RAkZv6AWybNJsF4m70yuAy4c+yM3M43gbE2lZWSPNSb3ApL1V
nHLWDTiRTpYjZaKIpQ7mkwxPiUNnqRjHBrMIj6HEuVBrjMr7wxik8mqz6VF3whWF
PKRklyikrTkfIngMfdbQa/ZUNzFkRLVh8485bUNOc/hYskhWu1zNeArXsRsSGWKL
3jF/bUUiUUZRjyj+8Qe8AGHnEOVd4YQ2OB23tN4O23PixsFgjyjTdC5+RTYo6kcU
DVMSeHkxEaJhnDTG8EITH6zFuIpV+cI4ol1pw0/fqyByQQLtlqze6EYDbJlC9IbW
8Xy/P0HiJNU0z87w1QsYudya5ZLOms523/S/5zO/rPLzOHUXOPUkm76BumBjzZrm
t2uQgoZAg2B/ZwRVDPfRfuuZo3Au6QLWp525lYE1GmOBaLIzIRHickiADVnJ33L7
cPCVScWeOmDhdYpVBb9oj6QIlAiMdT/8AG6F3+r3vZjTXgrCE1tUIi/BUUHVzioA
4GB1FvrpbASsgdYUGkTu8bBfsAr+TPWnH/DK7Ru6Lyf1XAOdzILj4qHLdaH0P1R+
Qf4zadUfs4S+4+tKkSSjswgA2Ir2Gk+i29IrSvfSxrU4JHBpWBGpetFGhBW89uzC
QSA76nJgw2AxdoZWIAnYrV6njD2OTttAcyklTeGdOX1/lz/cab2T5NRaXHUOL5RF
CHZG1PP3afHybHuhiSHFvxHluPFs2E0XPkJdal8y78WqBPEgJJFo/CztHkk9NJjX
z13R7VCtIK1K8AlV34M/CDHQChgksfwXWnC6n5dJK2EMQRSJGf4vJGguEKTemi0x
Gyp4LZ2JA4etI6bFtYF7N+1AIltxh84cCbE48NlYDMDVcCT+ySvlyu2mB7P3BC1a
wNmmpXxpxSd80IkZh0kDQWpKxRhiCD+vqdF/elRkqzc973cu73MLu14Ue7UIXsy6
zd6/9Lono6srw2bwSbIlxHYEkAeR8CPr/B0Ul5CVX0qpc8RzdAnEv2TDS8ZCwhqT
Oq4Au6tE3SOCFEQgq2oBoN6qC3ssWfh12PEidTXxDr9dvYZgmI3j0bZRJLR9zEqt
Zh5/ej+TUHxfScpfXTWhD4jpSXBQGDicqFWhSTsFhzC2Fpt7NNbl2J0hqIGMs2pf
/0P230h4wj4nefZ3ZHliwiodDsiOMZBGtBuv8SaMDNdhAZM/GtaUKb1kbU+aBKm3
Rj2NQjzSlmJOKEYhDs/h+K85e5Bqhs2RAGuSk+ivVT6o6Jl93CTHxPpdhLs75hM9
Upzrjyh62QsqpwbbkiyNGPjUfIscKj+HrqOT7mawd4W5cb6jZhz0V569ZsDsFUT+
5ekAVouLPZtAD9mw/5MYYa5+Zqc0WPSpiw24rOSiwWTWxblDIW3uVj03W6XfJMVd
cnzVgVP/Dcp8TnfdYvWisqqs5jHLI2BEAuWUoMefDJ98bvygED4mWA+/3PJcoyJs
9YDwi6DQ1argSIDvlPyNCQy9o4IRizUr/0Fp49YwLUUVuD84XMfDGHLDvms/MuuN
GM3O79jjo4IORrUw3isjYQRg01UrzkqSyX21aRIS6FJIvHND2g9k9WlIcFnR3Y2K
j49ThxDLFO5XtM62OfY05e6xzjw5z2kqSKDj+6HcVVmGNKSmSSmzbA5hH6U94rS6
zPjnddYGubm5NogidwR724YvB+TvuN6+cnwxSoUXpk5mE34FCYgSNiThCvqZh5u3
/GPZ7Uc2AHO/5jXd2Apr8Ery3S95WPtG/Fi4QqpGnNXATTggXtsbXosxMd/V/a1z
vYGIhhXkYtpUYzEWfw9vMACE+AJDzCqIgYGWnJFGa331lED2hM5W0hnMOstB18C7
9Fmx86hs5UfI33V9xoiZS6RKfoaYSXZBCAE7GVvOmoF+YSvXN3rGbKyINNnkT4NJ
5p1il6GYWSsVV3dCkFeNLjPINyEYqi3TUFHgwZTZU2NEb0Gno/Ft0AqLw61lTZaM
PXoVbgJLUen8kN0i3MzDKP2k31GILfQyQ70+5Icu69NUcQFRLsQvGciWBIdtuQ8s
VqjYleDFbbWuSZ+rAP5ywrWosqoB/7yvXLIigabPFmE7fjjhj/xSg12pYQ68ucYH
pjEoq1irPCaokwyPhrEp5NcajekC1rUgfqputmHa67uZcJ74fiqMimEHw9D24PRj
Vm9up3BvvS5p6oDSepQxGfipTgJWgqWf2HGvehXBIO+yVZT15UC/DdBTIt4KPNW8
9Hx8WJboWKiFBeDuWpnAvPzH2AyxgURRcpR1lshXGO+3YHQ6JfGiZH/9mKnpmTM0
skWD/U/cs6MBgnsWn7B4RUQ+T8CWQXEr7y+3wH0BpQ3dguxT0uHfV63prEWh+M4d
iJlkmR34Su+OxObtjmz5bHvbEoG5u4Pz0HvnKyDTef6emQ37ApQgjcxosQMOt73r
xWoiRCAsofgKV7mHJj7YrttWWILo83FWEu8Fy1ERetgCrE6tA1oxNfbiCxTtFgmT
88wnhZUIkzqgY6hCgzzYCMCvogjktYyWr1TZXc0kyng0kOMiS+3CaAwRFOXzuCOw
8eWmi4s/Y5ORiZiOP8QDLxmdpHXDfGy2TyTQ96gQPb/h8ORf5RfsFMj43rW0TIRl
79SMA8DUBNRbyFOUg2t6l2ItSM/4wl4VeotW9fqYaijrCiFNw3vez7GeG8P/T696
+8dk0fYoMryMPMiaG9wcWwv8Ksstb6eZIi7C4ZW7Fs5Pwx2PanK8XWCai2xBo1C6
2+Khowyh41e+Zi66WzPl+qx+3p0Tstkvb6TS1pAtnYAzlKpbCWpOj++WZ65I8ZvD
OmavTurb4bdgmvDZ9l5C8R5/I7i8fzyvupU3nMV678PBLrLxNnesDM6RigBB/b01
cdNz43GMek+34Qa4YXzVHILiOCE0YzZHsOj4oy6NTzmfvKlcZsSkjcmXwPqdRk2f
IPqe42YNrQvXg2E7H4l1ZbY40MTU90JzKbPMBw9dtqB4oVPykJifR+1yfBeM8jW7
Whej9KlKCZ/EGMVrCqLWnKy9hLCiY5wHmlkyOGMxp4EN7KmNHlLmpMWniJ798X3T
+CTP1ciaszaXnLLzp0lK6EIvDPuuF8NuHOlQmT6k7IF4/Z5w71L+Rgcx9a0jTa7L
kZ9apnq+bRgg7dWLg60Kdll7t+iL8hWThPGoqgoX4OkaLPs6X8ycKjhC9VR4DOuU
Q8Ky7qPdq1TO/WUP2Ejg9y5CHsKlMOkpEv9ZWzvllFx+ycmUkyiEK5Wq2iP2fH89
xr5LUFQ8H2S3O7rMoQUS1fc1PWNWRYk8RYf1NcuXQxg/z6XixFO7tNwa8S7VQOc2
CrF91qZCVVr/APKi23cPkwreh6F8oZyBQmvEgWEdObwP7/kVEnnudFdMZk9qYesX
7gVAIkFaAm+7lTWhK42xfMjEHaahQAY+bu9/wBqF5+DyynZ88svOLoqn466i/cpy
2XZehsInlnjMuTfybV5AXLpV0JXqAZD+unhaMDSTfbFvpKP/7i+XX/Ilkndd4F09
lhCmz8WvZuNxusCBwb+TmYU9lSXi+LuljupdrVFZ94g0d3/CMDFpcXFDYUS/xBD1
RtoP2LBmgLT3pxlysaD31dqAZN5IPdPLwox3XSWJCEsM6GdLBpNtqwanfsQAseu1
BjNYrqsQ/07ItKkO7pSzSohSW1kxhYZLACREukWAmvSRTDcmYfvP3OGeles25Ok+
gFbNNF2Tyqjky+s3Jy1YXCoh+KzGgS8iV91b5B4tK5sjNHvvz9XRJ8ngOBuXlcYo
ftmJT+31EbvZhqbYX6AtoCo4+TXm7ArAt1Ato5lR6/pjjHZXUXhG39IWYkjJb7FX
YLtkVq7gbeqH3KspLUNorJ35mGoOzPAGzPauqhzeaobAgrmiEsPD4l0pNR2tL0Kk
Si/52PlttShYuH45jCh3o+vz14FXbNCsClVq7cMdtzTLvfQFobl0pftrH//H0hrR
XRaaSPPLaMt0jdK+0Jl1tXyMOyQouDtUPGZjngFrQ48OVLqLutOfEPZ6PcKAi20Z
PPRcEfZVYEvhh8Qybu5wpxP0yBzJDg257s2bCwQxVshytNWTLsuwXrRQjhf5aqgt
o109QRPkjG5wZ5lfuSTj121vXkK/votDe4HWfCZ70QrRr0mjoyrIvUs/Ex6zdvTE
ZO67y10Faxy1YFyGXn6lBH5hkYykW+UWyPBNpRJrN9nXn6U+z51vOCzsVbaNujUu
DbbmDwU1FVTwwzSIv54Pv1MD+wqbe34vB8CDT2uPmAbW99yjkqlaXV521r9O7WQD
QmbFr1DakZ0cC+r7P3DDhGQmecq0yEDHcfA6PsBh9FTJRkEtiZu47mFIF8R3Erq5
pMz4lXptFVfVRmPs7cS9+FLSm3QdHsXF7tehgDB40N7q6QRUWD8/oEDK/du8UJbS
DZDlFiQ1do7Etq19A9ltn72JBl1AQUPAXRjgyrsHQjbbMZo3YoxkNQZP1fWqCGAl
0bDVTHMIfqHoR5ZlCXYDDIrMgGUfYz8OlFVvPHu/yVJdPfqz9vVqOT3srMkv6FaJ
WxuLymjvj12J6oq52k57huhkqNU6y6DPgg8thsZvoxvqzwCCJrgu8clyxRXKUAEX
nWmFarxpw0OcIUpJrOkNbDe/S2GpjiZLRzAvssgOyHdftAZTPiOUMiNn/umMqDeX
8LkRQDNcPcd7f05IKdcDecrDFawL0njx8EcaOa0kstLNQIoaelM/ececl69u52cd
Si27uMkKtKUh8F9cx9kgnVyTMvuWO129dRQQb4w249Cd1VDWbZOKLKjW8LTRgfdL
ZelEosWhTlvMT3jIyu/QaPZIZSniDuF2KWNBWNPv/mzUtO4VOqWyg3NsluSS07yT
PYvQSl4D1wUAu4CynWH1q6JSgFkNvdFVBTTt2nSp1gVgNwdx4hJUgGm1Ey9n2G3M
httFlwQ8wzF/nDoE1IZZCgiLQGG2j6QRqB3wcGeMIZhQuYbvHKxBYPosK5cdSvtM
BM64djORLozmM2hyy7aivXfdBo23iYZRIMRYsPWMf/ifah5v20rbcQQZf4FA50lg
PbAqtnSjcX/+dsNBtZwdRMd6sPywizqDRn9Oz7ZwbHqYM+1dGah2qz+WkNonUX9o
B8G6dT3VFAXi4ThwjtGWFbm3ll/RIJOS6exXuBTY5DtDHaxZzlos1xc5iCPt7gl6
6S0u8l/W07Yn5FkDBbwkbtyCKX/7wZ7I3Bb5Vppz8mEt7YznwgfI1y/7JzgLRGeU
bb+XHkxCqlc9BQCSIK3Gek7S3vcbMEtK+xh9/tKvHIdZRGnZh3J82dUDlgpgwdTY
NyOGk5O9H/twnjQX0DquuIVJaPW5wjsw7syEdjmh8VxfYFlERocTtYXtfKkmno6P
bRyyO0aU8WfVD/mKKK2dPzoV9dFwEkaDnfG+jPzOZusCx3iYoWN1wyITA+L8LRe2
ZHgwEhIYaotSnturJadkRFVD/6SYkyvwEDQ7ZvcfVqcBsB/f2Ih79XXIdjHGbU+s
A/XQ60eLm5Ps9nUkkDYtk/yXke5cAZKijE9uODPTAFZexzr2t4ozD/5NF8aO11tl
t2MM28Tuz3Jw/aDIvCON+2+Vy/fzaA1A7NF/tRakNgY3uhagWFzK05EKGzx2cXXk
l9HUbWMd4nG3B/aFDomWCadvmNFrZWYksZWAdTrtJq0gJzlmGkZkxkraCzGzVAJx
Zh06aOajoC7HbbmE+XZp19cfuVyHWX5DGdC2FgDUAWXMmpsE8NlZ4HLsHt1Q/9Ro
sD7Uclf+jrP2D2TrdhZSxRwhJakLOEycJzlHKJWXxscW53gdThbk2C/g2tJil794
ZsUSPZ3kLaBlEexBJh0NQ/AV1l2OprdUvBdBr1xILbA4Vrnzu7rNkjt38aB4OOaj
odmFKPP8Y9HWbERsfFMPsA2IIteJc/y8UVra6DaoxQNh4wAileGEZwGqew23QYPR
4j0giO934j/iOzZvcOzQCq11Hq4mNqEDmzzdqyo/GcI3CZRTq9XYopMluUySYKR6
tnuKVCpeaKS5J2EfS7svSFAd4mMKLZTlyI2pgy+vuBOsMe+BU751j6h06U6qkFur
M7U0xzxb0penhu+4wLS+uYV0Z8Dt6wjujU1Y3kQe0XeE1VrwyjFAfu3eCMRwjGQR
uKfLt5LrSVHnby566hGcYKHCNaq+zJ0H5nloh9zLQIEAaaOlBjr/Bt+VP3DkB6vP
IzqJzc9iftCOn2EgldhoWI6fQdwiwyXtabG1g/+WkT3L0H4/SAH1L+9tkJAjmo0U
WbAgdvnHoWcBQ575cYr5TL2ew9AciKv0Xd2GLR7AaUNl5NgFb2aZrXlws4GwenK/
Y/2BA+PEE5unV1/+5hDN31X0YFQhGw/KUK8AoIFpvqcZS/gCvvTnJhIDGlrGstEK
97j+EWhgJUElUmEAuhSQFiZwHBfR/vzWlmO9U3PtHctwUDmdgLxPbTvR156hIZMM
sh4RfBsjuusYm1u9ddFZ7WL6qITv2eS4ZDNWJabp+k0FzT9iytnuxhi08qlImeNW
c5pOvqKwncozzsfwinyHjdD9ragASM3qEhEf+Mc8oeXA9ZeZ0yuwOg9WaiE1Krha
1PqWrlafxSW7lLfaJUPQwKuPWkrAZE5HmBFijPdJI64hMvr82Ta4pxBfDJ6fCPXy
CgD5gRu3EnZcrZSpVfv1yR4PaohfkMCjNHhdJrZFzVT2UL62uba/Gd2q/bKehlHo
jRoFWxW8GTcXfL3hwfqCHCagmbeXL2GKgnemlWDJ0ig+vXVx92uL3PZBgK18aunt
lqkTOWnV1y3zZBAG7m1CtoCLoFkvZlOb6aALK3Gbb7ViDk5L9QhVNlG2mIawuAwn
lNC5QC/TzO/bI1TujgqEtD3nMsOZdmyLTGSjDCtb1ZOvfiYWfHnjLQhRLkrvJgZB
IQdeM6ZCTw8p1lgmxg+/gtJhC4/tAgtbl5b5sgJRaLyt6vZCdT2C94oNZyMcdlxb
NEOuCzYMkqbWdlr3aFxqqcDT3zlT3/iRuTecDwpK6h6eQKIODv24JE/KSsEpSngY
ZpqCOg8B3X+VRo110SWfNBXxmsznmk8fnzp72CMofFZ4W8yQ1Irdm/adR/RzuKka
Sr4N1AJaxWUbQUjSk08gotTSePUy1u0F5yF7tCYMilSTqT6tUOXLSON4uB9ervxU
VuvOuiqO3w4Rc7q4t1lcJbQLC8nG6l1Gm8Ht/fqrMuvSNixDnNjeckz4ofIbFCoP
RHae7PBY7miJxIcIy6s0XjTxHO5fmOjGIEXN20nGBd7AIWZUNlG11YEqCjXtZu7y
DzNnEIFHD0Et0HnaJ0rol0a8gg1rRu5Ql+RXkNafc7kq4ScbJnNXm8YAvDHIBU//
qUu5wZPp9AnRZAJSjze3bKeL6muk62kJ6uo0+jF6OiJLEaMeX4GPKuB1sUCgI5xK
+P4jfVJ8nuTZfucNfsjS5LVeGin66fWUFvu8Zu1aOVGaZU4N8HirMj2xoHQkKgrx
eggqYVjAmDe4DUp/FsCaTrI7ZTL/DF6z0zA7cZ8KOgqfsFa6GK6OpWEg3A+PUyig
LifBRRFNzqX9s6WsgrIKm6xcS0oNjZEGMtEOLm5CQ6ud91c44vqYgHS7W7yWcacZ
b1fXqLHP6RzHHuD63ogpjluOECG+fgBRZ0wyMO+NRlGXwrWsTAckPq3+ZWLW0aJe
nc0oOdN9/ywfopAib6eQmrS06PggTTHudtAMw12dbEayYewG5gaXBPOAzt/6VYlc
+VeRpPSQDTZmv5W9HSmr/gcYB0vNkhoerBEDx7VgO3N1giKW2gApXnMmW2OVRTxN
oYXKxxPr3s0fr/F4eoib4hFNArwJJXEqUEj0Zz2XRlNRazSAhmXRfEFpeveSd/T/
5mqH8vNTOG/aDKZQQETcCZMvlwo2vxTiWWk9HXunfcRfWzkMvgWlrAJB9WYHVbkZ
bhqRi/EVlH9ZsCnduSVPQZbh8wWfbqYnIG+Fa2uW1UQjgo8mcBGwfD/da5PRpFrh
EMLf4EFcsP5qowZy3PuUXR4e6JBHJqKk/E6dtXlclBmmi1A5SKMOWZl9H7kfJY/Y
laUfdIYhXuE9gWnAaDX/uVPqZW2Ae67+wWAj0fSMnqWDb7I6gdmdW/EC4BODlZZ+
3oSbjO8E5xGSY9wZQpxIY8Q5y1/hn1d+cjTn1G3rhI3At4GsI8AXjHZHijQty5yN
dSJ+M/fV/ZYJaRaWmRX+WOWXU0+JBU9/aEzKqghnrzONZ21rDIoxgVFieRAFVNjB
KazU2sIMiQqJbmPAfp2vgR7lS+4bqr2Zo4Vz0+6PEzaVhVrwuLm39XfJub69tYON
rVXpFZC6z2QxJYY2EeKhWXfN9IOU2wRoxztExq8Oubd7he7IF9374U40A4ei3J8G
cqsgVcLnH7nef4vGk0HQUSfo8yc0OWj5F67ct/qsbxpH0s8WICRLYBp7jNrWdfGY
zXvIPVT/sAsQcu6jC0B/acmqDwWOVHnfMuPjFL4z9AmuueF/Gbjp8apdYwudLNSO
iljS16SLCTb9+JJaKYdQ1IA7ydcb9sVdkxB4TtoLIA5FkbSjjdh2PJXULd9BqfaO
DAlzgn0gCKflyXCAggbMzszoTKd0asayC4llug4uQdOEw1U7iX3AV9U1a151s4+q
qpkEg8zAZZd4q/YtNrovcdflGmNIldxsPqNOLHXiyGqhbB8QroqFvsMK8oL1Mzug
2F1r2LXvgRyW+7XMxq71x5+Thr0eWM6ww3yI1bdqVZfL8cdJ7Z40HytDZ7rvkpt9
BzsmKnbPSDML9o736gQfHqnimEorJFsipJU0nXhQtovM4bfhlmr2YiyzdHutri13
u4p4kEmrncjjSQMXv3Vb0svr6r+wjl3+NkzJEGEaLOfJzm/KMBW+qG180N/lVRLT
UJdBP2PArYBdrUtLCBSwq7ncMLig8WJYDabwQHwl/9/yHwdG/ZIcQZGXeDILIzVA
4LP56ZYHaqSIMvTsZA8TLHjjPUZhm2d56/YvbpqMWmA5NuNXMnGwh+ZhED3h8WkC
SzZV6jDnrCH22xh+hA6p3TLdd3YebLaRstvC9Wc1pRbmuSdc5wkbBdOb5STdddCC
FPIrr+GcOgfJv5eFB4hh2CfdBFYBrhdr0xLea+4cvap/yKH7rHfufhqGCVNZ4cmd
rmINRBmSVQdqFPniyMYc5lQkNatPFXXivwf7S9smNwqqUp5pq+XHIV8pes9XD4CL
sGwBpAHuJLlZ35zI6PJ5Ti6SxEgAmMXeJYHZpELsmVfcXT7dmoWtpLBAICCE5NUT
Y/rMe3+lkSU/bNpqz2GqZmoTQX7IkUA8laVyQy6MpuhbsdbhUbxrzVD65cTTeHhC
TFWEnQkQ5hYCp/jcwIddIRN9T/IlLfvywEfqUw39lAvuRh2kkwE131XMIAmcAE57
14vqruFoUeluA85DMcvmbz6sWnPSPgCrPgBAGSu8JCCyh03oxUGo2bCQdP8Gdclr
hqtkIsvn+4WMH9r9MNBFftpNQdZ2MD0rgFOJjXJIFsjnWR/mw9jRaX+LzyhC1qu0
wV1JacfCKwsMTmnlnnROU99U36rZ6KL8dRwZTpuM1jhnb6OD5921ah09p8+aHtrm
IDyMtPwg7KUZSj9XfUX7WbeCHn/NYyxJ/k82R5tx2YYRZsqjrgcLwCgY/qXmdcsu
lfbKbdiObPec11wFmmM+G6CP3WgmFpjnA0jUEuGY+FeQLI8JLDkqDzXyA8vsSVFh
Z3qMcRQ5yqqjWhAOztofSx1ezKKpwirQV2o3mWj9D9LhM5hp5vWHYqby6dG1IpTu
JK67kzywMadFR7prx3AbaLc0VPe1Q+s418nrSfdInf3shisbG7bspJcVczPhdKig
NRmq6K39M0ZQqm1hNlm5FrxyQBfulzuH/miEp6V7QpvVGa2yihrlimzr0RJw88gG
ZhrB4Z++MGEqGEMw1JK3JGCxeiXpgRveWxBWJEIScqRIz9p2zcFjt4Izs3V++rzD
0JDRMQHJRfv4FI5SAIxFyM8erCQK7UuztbfHyrN2tD2vz27rapNyxr9BJrcoPlgw
0XlRN1xPw8ibHH8TG6SqSn/SkBZQDatTxDx3M26pXgLePVXF+nAfEbLG82gFqFgt
Vw9Y6XVGVfQMLw96EdlX/bXzy+4rQGR2jJckNMAlCY8dSoZWx1450aRhB077a46o
TJGX2ZW0iDJCk36j4ajSLAj0I4/xr/ZAXc5tRI6Ebc6Kon8ofxXsf3OwvOR/NLBf
3QnQ9B2DA3H54f2CxL965iHmhYJV1gFAB9xBjyePNdeqFyqHTq/L6u8UN+0QIHqG
F8LX3VUn8iQul9oS99WFMivU8+JhkrNXExhZzOt8MnmdD+4xIkPE8oqrtTXfVC4z
Be1tX2RgXqMYhgugdCP0tqrvBWg85WjpnBnRKnPwj73VLcBxQyTEQSfASsI9ZrRN
0zgRxgR8Okx2qjr1L1Y8EgzZitpWCKlCs+0jMCIzTL9iFVS35deHxHpdnWzV7IEw
1WtEKZ+Tah6o3khrab1R5Srfl1Y9g1LGt+2HIqpU65G6kv8F1xDIDmwh7TVYkQfZ
C/MAKZQvP3iDNyrvoT2VT4cs+U4/FzADD6mV2uVqAsPXnuBG+hI9BrV0AkhcE1fk
OQ1iU87cNQ/tcxw2aCvfL7U02Df2Y6fiRIcm4kklhZ1Vt45Qg8jMAdUAYj7IvKMQ
n3T7h47EQdWgLFDipg5UmA3taiCciKr4fOwrvW7ogSWw3k9J2epyip6qWGihAMmd
fGgc2Ec5XB+O4i9Y0YI5fqk7sypH/kCcK84Z1893pXcIKvxrA+HNgds9MWJR8mFI
LdZd1LzEJF31Z3NhYX1RFz+w5bdd+IsUlv/whu53IN0DPxl0KzsaVooOTwFafv1A
VjgLnwkvekMNgBSA60rWQP3yy1HcnsLdGJaIP4qT+gx0+baWZiWqWMuJucd/SNFG
2sei3NX7StsBluQ3z3F/wiuF8ejhCkvoXd4bfALWG72IXC600nFbUnmI6/XmahRS
EakGuZkCjbsOfPl8k99X+pKZrnfyUWL/hdg5n27qy89zddLzhGVSBU/r8Wq4OzVT
X00juD3KhbK7j2aKsnwcHERnLlxlO/CxSAZlhhiUA5sC/ES5Gpi2Ln2K5r3CnmW7
pMCDU54kX1nSQwqZaKWNdteL8U0LAP1aLl1vZQ5qlE5mlODyP81a+hLgtbNez+nm
y7Gi7AlMx+t8zVsRAHcEB0nQfN7DXH/EqwmHqeL4Edq6agKBOj9njWilA87CAdGG
9YvoUt3fET/UzxAarAK7w5Ju0rwvgvjAsjZlU0rDP1x/uPLZwtVEpAAEKZzRLTje
8jhfq94pf6QHv1eV/kh4k3rFh2I6e27f7StrN+8fl5hZmgwh44Few4/RkR7yxaMk
3tcDbvex/XSktrfWmeyJezuWN9vzmSM6UWTUcFdEaPaprgKjkXwQmz+fPpk3ETnr
sKvn0VnqwgOUzE4BoBkhrv+HGKytfFvsW/6z2WN+6wnqDbhx5UYyHHJ4PxsTOZQE
BaXjtVRX8Ia5tlGwozKdx1tX7i/rF2TOa0dyf3c+H5/vKZfAwjE6A96ncHnEnMEF
apnzyNvBrSlZU8tyfdRPtejAZeT2E60GrOhE+bn59ptgyi9vqOkFU/F5KBih7TCw
WqKtV3Tr+nwwlY+BdkqerhEXbyA4eMuZWE7lmoxPJCe0Pjw7sFc1serFoggXLOOi
dFR2341akVJMl0GgHlKyTP0hF+kEQL39ubBpVHxXZf6f9VjL8GvTEQ/3FGz248Pf
Rm2GR9Wg8nntPBePB0mY6X0drm/UEut0WkVonhVeWFyrmjP8MYRF3/cxXAPbYZUR
NJxhJxt28hh8NyWiXlT2KIqMUaH53PcIDpihg4OY6E+XJN9exMS3veqwpdGzZ8Mo
14Mx6qsrYfIHYx+Kw2qONKuwMJiFKG6hiO7K67heE+5DbABkhUsSBzY5SBrNNYQ6
h1bjcSxIkS3nlhkmRzQKZcDou7SEPOz2sG3D06UQXMujyGRB3Z90bUvSr7MeG7Zr
AAwSwabVjMD46/QrEGciK+xcTbFMJciD2RdkoOhOzakTIMTx0Pzdjjoax0/hPM4K
G8cCeUw6Ey2DHBgZbWNhD7FUoS9s+Y1xQonOS6PV+pVaqeljINNd0apM+IDgBEpR
3/aTerblfoI+LLvcSARP1gM8sdycrU6//vwmvNYKYd4hF36cT+JpBCOALU3ULJ0A
AmIk0zDS/+0U+DCHkNUTlj89oALECNFYoflioe6j1bW5ueyyysw6jVyDTxOhIqtN
d3OajvgVx69HuDnnQjqoeoAoXR0sxq0fnQEqTeybRB+SDNYesSJjBwbVO5SjG799
4M0Dooo/ygbxN6htKeSms7tDtMxw27BoFAGwQ7KHXKRHkoVKeHc8sA70kR4TpaJi
4Z1oJFFkXQeDo4YbMG/JDbBmsXtmpxbuSJtyU5/ls1JTGdRJ1SwCbDmAfbZk/xfQ
F3V0o+buKxZlaGM9m0GNahtwHucUYh6iLoAEhWatOm8ZyF0lZNpTJWxWQAJ3TwkE
3PvMvbxkYtCebXEahtsI/MNCHuDthLTwYmacJkOAofsd+A8q2sagGMe/LEvM9a63
B9lmfPXYNoxGaVC+7MPIHjk+VXEWRILsRDCjjCImUTksAt5x+h5pAh6L2gzfP4Eu
vDQMnajKttx6qzBMeqJf5LUDvStllpSysEDpXFCrCOs2jL2dKh5WGds2iIbNfmsZ
9ZxQCk9DFGafck83af0LMT0GJ+AHSDO0ekU7TY0kdYFh/SH0qibqj7w7sszjhuI7
vU4k5vAsYcBamvgDJeQtn/2jXThGtYlzzKkchBIQNe5kgOGAayCcJPK6MNA5JVjg
WBqjVcK4G+0lpYd5FzjE5EfGUap6Wft7YU8WGIa6v9spqoYQ1X/+bbJFar4nbBc4
7iLKV9IOKo3U1VXFLBk0RLrf3UXoIUQIvRsAZp8xpQPe7UYU7AMtHF62vtvPmwQn
dYcYIoj4zpKEsjc7/vq2mRMBzPr40tGNsU2ZDty3vvYQYhDj4rYWiu3I0ul37gX5
Watnhi0G8wKp5m2nPqewQaV73padvydJLknJn89AziJsV5LBm9TzUfrulKGsNs7t
R/s+cszdBs18fWxdiYKmbzL5QT4RSLYPt+1BwJJVAkuA7BMo7jUNbrhQ8jyOKn/B
lGaF2GN297/0CjjQkt8gJzd6FKzMlqPsfptX28uf+jQA27gZue+mZbLFiaZgoYLD
MKkTojHIS4VYT1CA917+NDis37MeF1SZMMO0jG1jlM3cSDr/CQtNAfKaQTTqEc1B
VN698Hftby0gUunfA88sySlhwu5+DnGeqY+Q0qydnc8V59Yipcg1U0Roa/wWLUYz
PGGN9rX0O6RKNsKASGeNoovDNT85GSUWtsbCeP26Xam2aHcD1wkSKNXtv2VrQ00t
FeF5xV9gCjI3OGAY468QkI/dyUnZL4lVsiPzurtBNa7Ad7kisgeGiituFgmUO3hn
6jPJNgoD1nday1vu2f6pgzgdcgFkcS/dqDlQdD7CZUpsqRz0aQai0/UAbVG2pOYp
z3Wg14uC4pupZW5AgeKsOPjqE/Wymvg/+3HBhWyOn6/XdUvAlBMsBjh51LoZF6Y4
irEW9BdC5pJ+uH0vWgxh3ef6+N7ie79oEANaEikPGwj0K1V+IhGBSVKY9nqD8Ro/
o0+5JqMHuokvwvri6MzHdNzIabU31T3uiJhAcsJcAmiknpQzXZ+kf00uDHQ+K4kT
IRJ0RQ8Z8TAxJdsUOgPw7rLNNVzsq5oq61QJwCTnIo5prS2Q9IapO8k4VMPfDSq1
61fe+S3ZgxVLFq6ROz9oZp/hVPqvbhelSdAv/xr1+3yy2tu386FHrZtuOXPkHcr5
e6bVgFiFqwGURfxBDC2R+lNgrtoKqT7uoTUq++8sPBCIjoxvOGrQgJokkvmG9TWi
123h+JvLszqiW/syKBHP/91EFb46Qqf0zVDmfHLTRmDP+awMaTFpbWo8P2mKclkL
XJ3/ksCAWioM+4hnFqRs3+jK0YNnjUJPWB+j9G5ibLw6+nVEIrfcgL9SzSq1krqZ
ni04eMjI52LBmJrJgukHBBSpXCQ3cdjQ3dX2/H2u2TZwaPbZHbVvudi4nkKyDHL4
bSfeFt8lmFuYWK1KpFMSQ2kONWplh8hu4PKx+NDOwsiw/OVzwKxdth18akqadzD5
8DkyE05jRykM1HBwB8rdd/RgRJ8IysNBjIicuCv2QhsKeaTOJj1GWvu1GtZ97g5e
tzxlektnmyJg4XfrC5IAM7eCoj0XYUuOAB+KoDIsCc9SPhEwYwhJJQU2/QX882Il
Ph3uufhJdxZEYK/0ZhMzQD5qBDX/MnN6SfhC668ZL+lTCkM2J9f7o+ictfIhvD3L
69g3QgpN1HLs426QV3nz/bPa17+/SLaTNvXumDPbX6TiG2KIAIQN3irKCzpdq6Nr
KB+Osfc2ffRyzBTlpDx66wLPJFocPr7d3yABLVTULIM1dlVSD0E4+VjdRMe9bxuU
pa5sFgP4ohjfB/TRI/pZlQn7z3WQIS1+2/PenyDTQJHGA+krPg9H6p9r4xa+SLr/
ie61oazdoDvXzQyvzMq1Rb5RQrRcE7RjFt+rYm7/7eSoYkhG3t+pl3y4PYp3PM7t
kd1ExUssu6upb1hY9ol54ig1zHsF56SW+xbpUwwistXLTs39uLsgRyWbQPW6rQDb
9taQipTjcBdzQVgMvgHbCI1wmgXCvWmW0R1lUBkCmxD30cRuGH7nhO8YviPGnyP7
HeysOE0J3NZhegnmec2KiqZXuR/+pOiWvYDGHLFziOzfduzQxueD6MEoUAEeSkuV
U7fn+xk4Vl54LBjRMfB/tkwWsxF/dWcfHZEbqKJzBiJkUe+qZzBoGHmWTpWK3rGm
Kb0BxSNq4752zg++UTTY1Jd4X7rgKBqOEkqVZTjG/9j/Vq20zWFXnAUnv2VOJUZj
d1/fV0mFl3QJvIcLXdPwYPfPvExrV6YYJYwgX/gJrC8XaVsR4CFtu+LeNrwXsG+Y
jOJhpb1/D38mvGgJs8PC1wCCwoe5CBPA0dDKlVLdlKQuRPFZKaFdYdW+Q5IzXnsY
kC78oByi4ct3v5ufYLtfGUAWNDs9lMA1H1RFOeK0vmuZ/yuUhq2HpRH5VOAw6a3f
EqFYGWDewY76932QSf0kgB1BGiX8/TEbiuN8w8IXbPat2HnZBZN0Ze9kpEzMLyFN
Biv3vxH7v50MkX9kH6l/0sYfScYzF5vI05JglQYHLcvKiUzq9sYc7zGbj9op3kAA
4Kl/JDwxxdWIFSWeklpn5MJn48fT1j7jwPRGxguEyGKlQpnq/U54ZS62wlWezmil
IwfayidR93eZaIOHYckkYcr4308IOVdeBqTAnLPRbPz0DwPvrZAmKw6jgWw90r+9
n0AWPhgIDd1lZWc8rEYH/u7ICwK8yO1yLJQ2r46qknTGibUFii9dsI5bcZWt43Mn
JK46oGVh4ILni1du9gB6OFfn87NNBoLyEYk+WQDU/UL5WKn+UlzrfBWrA03KX+pX
T3rIkC7taHIzCxcFUCYEIkYBwpccy6PNk1yhD5DU+abQ/4ae9QEou5MgUzX9ROPI
crsFO/i17HfvBSWRcPgdjynecfLjxksdGVr2zvoWzhyQACBJSMSe2xOF3m04vxI1
98lCVm64NjYVEi5p8NeDUnbLlOkdh3msLoV2k912ukvosSQqhrLUjFWTPP/zDiIP
mTM78d2xBTgIrsMY4OG2+L6VcE3m4XVhDbJ3elSzEuKKplZqGZ7Gradvkii7GEfG
Jh7odacpNBgIARLbswebm3osGuhp6/WbXfke2pVTvdW93CHrMX6RqkACuwHXlJ11
+Cpb/iMyAN6CPiiGEby/FYbPRAONAYacIzyaq35RFQMx3LKQ1QqclmpbsudvSgY9
4CLNWzuNWNKWScnbXa5gwe+iVPHX6eN6mfcqiEqEKyuSjbeTcEsnSYOIxSgnOXe6
ccdo5ECfdF7vAFSAM/qgI/QMjTQf7/AhgcccLpMP7FtrOe3jt7hMayxQZP8ByKwh
IXpoqdl3ukRR9eYRRAIVzkGlYyEJo7xRhKZYBqCyJ14zCXxLckwkCzKP0tAKXYyo
lb6U53uakyy86SeAcB+XlAJ+SQVDoGOJh16zlOCBBbZZcekildQbtYsXru8qokS8
`protect end_protected