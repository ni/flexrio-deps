`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Jm2uGAVYfY7w9Y5qKstopObZuZAEY3b/Io3MSEcWLhjjnKulVhCBBYAEQrAzzGsT
vMbffkdZgjdXQUg8jOLJXSHZ0Dgbnob2vlppjZs3bgyHCF7MoJ35E+LOsaLimUA7
hlqStcK49hR1hdeBPr/OwfT3UeVrRtQyq0eJXQ1UksinX1G9Pz3/CmcGfTZ/C72x
p9icpt0bkY4/1I4GBvNCsA6FFKH947JqH27OPACiQQRW/K7JToQn+1uhWr3LA1od
lbVrWu8PdZi7zW9gK3jiW5GaPjwbYQGqeGFs3bTKBILjb7sYHxfxw7eDLVMAIu5D
W+OTIN4JiHiE1gCnNEvkSQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="pm+c2fYA/4JT1uhlJGVUubML8hZi8lME4xPobg/m8uM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
nBaXksR//iZ9fraC7WMJWWSrjqRXHxmM1Y0+KKN3b10NElDzVNMlR76DLrcnamFd
2n7uzsxWqhhJR5LBl98SXO3Y90J6BMbw+OBG/MFM/zUulxh2Si5YK5G9GCrG9gvZ
5JomxuZFDu9CzlWGTuRUt6FsE4Lr6sOL1P+hraQDpMk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="M8TXDiNa0BVMX1P60yIvW2WA9jKGGy8GtbuPknDnC9I="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 41760 )
`protect data_block
/5TNZvs8Nu0G+mfp7M8H+iVAGG3Mh5DYZ0Gn3rRNhV8b5CcJKgjQajrRoGl/gSxp
rBAhtT8Vd5eelHgtvBjpvFBA/EBUrRH6CG6pqRt9r2qUDt4UernbZbxC3BC14KYF
uTWOLC/d5Ruad8g2qo0MpJxorLz9qfFc5+vRHE+ydtDTaE7CLuuo8ONg151j/LoJ
i00Fx0WzkETbnl5kZuNOiym6xolLputMYJlA/8IDX8y/4AZAtE7p+UKzYiyX3B8v
VtGbh+morusTWOJj/JgzXD0EgxeubO22lPRyBDqVv7/HNyQ+624ynYIgADj4IAhk
pgvbn0yiSL8c0HuOVlcB/hy5brQ5/fR7e8ajbT6NpqSBI1a9ldrAI8KNJrZ9jIPE
GKRbqqfOfx9f+va9kItxU0oKam2X0H8UUdAYWXlMRrm50zE5iYRkQ27IF1gpQVeZ
fJ9/81f3tL+atxYndnAOE6JYm/hpbkb/0oaJTMVZkt1/uPojjdFwGuoyXIipubG+
AzQDEBLMjbknFW33+vQJdTPx76DxgVTibWHY9mWmO6Wfi30zknYKCOR+MnwnTIfi
e9t0ym5AjBnn8S2a5mt6NMkTwzlqRUoSsXWPV/rcsvC/dEG+bN5Nr2V4g2QEfwg2
e+Y0CWS4Wz1nT2F/Hoqat8pDN+fFWZbV30rT5bc/S9gYVTq29Qe3iMhRJ472UM5J
aDHVizH/N3Qvukhq8QjitXPPMsxsOURgAr4AS1kIdKzyqeruOkDQwBazbUWOpKXq
UepNCCqax1Sasb5duirw3oR2NBUsB1WdGq2vjgZsqh5t3WyKzVldWgrqFffp/NHm
mE1OcgOP6A7WCl1SB3NmFQskjf1+HcEC/kBTHF+UNKZNBWLJEQScHiBOy2nk+HZC
7ziI1RQMAPoUbpPrqaj7s0pozkRZROYybXCAqjgjrYIZBFU1hulPk02JMvD9IHwF
ttyBlfMnijjnm9r0vcU8lABSU0d5omzw4mCzr+zOsR+dRSIzDWGQQD+hJiFWqIUe
2JE+O30WoKwmQgLX42vx37K/Z/X2Bj1C6LJ4ZAPDE9AG2ZpuarAbREXZa3bsJ9GI
nauY10qdVbhqSszjf/sWaalEV03BJrbVyN831/CJxJ4oeRKEAGwoGkVa/z3aM50O
jNT8qjo9D2DUzRDkBjbdMJlTGp7O4CpNny41ImZEeGHibu4VOwmhUhQR41wH5dkz
Q9XEhVL2V6+xURkPVnFlNxVTb+MQAgbugK277CVW6Su0fysgcdYojJLP3u3y6ETw
Yhbi2bIjT40UKJETrS0q1IYs38X3kf2uaKP/11pq/SwBJ+gtmDCECHbAeKWEhbyJ
KfVcmDG75ikUOiy97brA0FSdqtZPGp/PGBaYyumCbljHv40vpNgmpp6jOrRcziDX
bdkKp+Xf0gLG6AlfSAzrrh++t9YvD7SOMOqy0zaS/BZ4cYYMhwmAc6CEDqO1YoD1
+gD5X7H3MH+S9JqbyqQYocrm/O5+P5T/vtcEda7jayzqQDcAChBjQLve53swmVH4
/GXHTER/BnTzDmzNV6n+6Nq906fItd4V3kGPnMbUxJ3IrDVxk0JC31iSuSbeAA9Z
3CH77R0qECHuxYUkciUxKtmeo7CiCSFL3vmFAAYlEaBrqqnWz4PEEYPj7+eaoXZY
zKgA77gvoLKy1pew6g/rHGFqIhg22w+/FdYqE9ajLt8OLzY35TGTuVe/bjJiH+mo
IjUNGIdzCCSN/bgaxdS7qXFJtfF4hj0pOPoZGVXyNqP3CtZGcXuvUVGK09vlXikb
H/fjAiKPFcX/0xpEsTzbBRe5EZ6fO9U5B4R+yvs4rvyEjQsHFWOCfxD5OI6IxfHs
XUJTvZdg+TyAIX8RHGxgk1ndTi9ds/albW1Sm9aFpVY6whj58xZaqctKtHn60SHP
VA84oWllhlKOZ1vrzAghaULcGEZTO3BDSm+Y1j7U3sGnzk4QldM2GRJHKQCD8nEk
sogknZBgGNGz91lYFYSFhwGLmaZ+eIpb0opr8TrLhLu9HHm1y7Wx6rdMK3z2YaiM
TPXumm4EljLpjG3iRPCRA4LuLSRvM5rFUgvt1XCQdopMzTWF4Bei2T/K8ebqEnBY
pfy8MyDPK65hylSrJlorsND/jAwMdMkJC5e/ROHohraWWJ38vR13o735hoGKgGrf
W80puJAE0FOaC6LKCWmsSz76YXkpULTdPEF+7tpS8aab3ugYAChf863hHHP7Y/eg
daISFcEyJ0tcxnGdbICCOAk2FhOYFW/10nc+TMeer/oytb4VF+Uhp1Jq3tC0U01e
jn7GaOQdSRG5jCbCfesmjiMUxIRjrz3NtedkCc7hXyp2IKHx8uLQm0WhLwV/g+2M
sHB6PDFHeGxEckQOOMVYZ5CVoLbCPn36hhbLfI0M5cEzqpgIUu6p4jGD+3onwIZb
oCASnZw5fUNSL+P0aA1QexMJN6Q8lPFNrNF4MlAn35/MttUsHsCa97A5kTAayNuZ
B0DOg/sfc28WjiWg92/ZGTg0Lp4t8X0Ugq8toFGeCm//HZ61mwupQNoY9gi+cntc
KgDUhKcCrcZyFjjtdK0w9tyqRHc/NYksK77qXJNA32A+HD/ph/LS3wtb476RXvMA
uEA8S3QJswFqKPR8DeC5Qk1o8DoXaGjqIOagu6qHpuyUoErD6jgNUyKd+4xPCaSv
StMRFq+6zZntKRUSBC/6nHQFSFUdZis1NOscP+Am6G/NCYrICYFd9TZI9VO0NcWE
ccg12SSJI3zR7tnovV1Q7ElCtw+sOJl+m5ZvluW9B/QK9EzpQDZtBcZJRH8FtQa3
wt45ftdd1WIsUjLxk7H6R6F/hfyuxkC8vSAWgp3vChFKsSw0H3k39rlx9h4iapz8
AGsgK7fIX4h74X598nXKOClmU2zEVxbl6vegM4r4YkUwmfuBHR2QiIilU7tDRoMX
nnyUr1uMkaq1ri+Hy1FbxPQJ4HeTHmn50UGXEf/7J20k3moJ7VZdPySQHWv71GRD
4g2gSXCRgOFURf34oQRfXp0TLEOcbkYqOa1tLmFer3EvT+Qn+zTRpHDjbmp1cOwK
HXBbkZk5eqIzJTbpxPq/lq8W2uaRwUz8xTE19a+iu1gGBbhLfr8io3tgwLBLX2So
troASpjkGB8fq4M0fq9uqoXa/TFmpycaMCYkuMDfveNpCgvXW6RY0bo3alZZZlzc
XswhGDW7IvyxaKXLGFfLrFjCmTsGCe/Tcrg1Pn1bY5QmhO81QcRfHNJ1YthlSDcg
LqYxWuv5py+wwE5bEBWv2dHUZ7u1xzByxx7AXMRbCnQ6ssCeikFv+RNTbyCoPOBG
/4RaSaWyVXputmNlx+Vs8aNGfQomyBOVlmAqtE/GyX2Hef8MiEUS6e4EzZ3whz8w
3oreevdEc93RZTJ12Hd0vtE4j64ceC5IOhbQ9O6tgkX0JfDGj16IebTD/bPwR8vf
Bnnm+KszMkP7m5bGiNSz20aX/ZgYmBYlPXt/2YLlktMNa+q2WrmbQ+ipfnfjyJVc
EphPrQ5KZSEJBcIiNMS82r5Trdzzn9sTnzZ8uPq0d7qWA4KB7x1xQYGi+4O8Hlrh
FiioyWokAIHo4Xq+SLL2effRXTnLH12QvtIaW3BmviNIJtwDiN6y2IQwPF/VGyn6
xjXUrM/GgOF7Jnc/KCHIDclJWo6tsoNIaaPWNULaDJiTd6QhyMduVsKnkpcQUAna
6KsRxTwIBY2ECjpLVhJqu2Y0bd+1n6JOgLFK5CRlAsZ+YGj18/glZmqvNSu8lQKD
aECsjokbh1t2eLaOC1ulqb0OGNPOFMq+gmoI8x/sn2C3s2EXhNYJkWw8Xw7fQFiV
vR3wUOdqcM1k0isfrsSHKWvzrXuI8svVbMGYij8CSa/ZS1zYb80vkyYT4EEc81hh
18kMqlczEqh1cnIWDdQZf8AbfUopTqkLlGftKRnSHGBqx6lmnnbRoofexmdZCEj7
oZo4Nv+81xH9lKVAscDhPG10oarZ4/CtxsV9gfwShmUTOK3HkO5tzI9Bj1xQlohU
PkKG21a4qksEiPS/KhcsO4WeEXP7WHW2uR6TRRBm+2S6hAgi6T0cyr9O7IN7M44E
7/0T5xnUawbBnF0QFaTtMK6PJe4vZRw0ffodqM7nCzgsL/Cg4SfXUsTbiUceqLNi
CmQb+pMH3gGlVvE48pFUmEaiVnN77ERkS5Te0d0291nHtcGvCOX4HVLts3mUkhMX
ObU0H2A+bwBcJkDePkQLc0yMT2KpKwo/KBHdgfVPDrF+QJI9jrmE4EmzK/qVMxkW
lBTNZVQBwWd0eOHW3h0fzPJIg2tyeiG1QL72B3phZQYlscLezBE4/q2/PKMdlS8S
T01y+nOj82v6fkDsbDaRBGktFtefG7qxEJb3wsRmYnnLNQP2bQhMoaTssBg/u8EO
KTg/BYkdn9KxI/UZd4FqDMBUwQtNrME6XGP1JPb61xt/F9ctUM6TF2Y67xg4Vh4C
uEQ0LBrYjDmgoGq9Rz0Flcv8nsN2pXbrRi2e1kWAJVLRM6fsnkDxwtvhrrSL5No1
Iq9xFpg9HsTEAsbSY8Ft+EVaFbEVsJHKaNEsofeQuBb09ggI2/fOtu7/w8J7rt5E
dTorGh+kQNPCWgbTeAkkHVgH1Prq8+VmMwVqBcsjR1QA0L+8FVyj5ob7Yh+ClLxt
KghWTpwY828wMcEqtDKsb92eynKPghXCUfizOVqMGknqqeLxXqODZqBEjALo90f3
WTsF1e7crtf1uKOFFSbAQSXZob9Y0PtWQ5dm0BhGlnDsqjHFyYZmFGiEmwxuD4D0
UObP08rkJY08/MDGCCvrSozHdiZxSKPcrOJYnMXY6S8I0FL+RMER/ddWmt83KTTc
JW3hJoyW1I0nBFIRWavzvXYZEt6yj17wK1vCjDCglU4ElyCTawZcjTGY8kfkrzx9
ShuOfnreKe2wxRziZBpMCs/8LagI3+lL6HRrG5fnidGsP1mc8iohg7Bn+ITXvQV/
pKtbF2IAJ6QLB23hixlwgS0Zk0OB25LDD9p1zaTZOG6vKgR0cxe+pNe7JmAa/YtK
1xKuMJY9cfz6ZO3mcQS4l5cG7utdXsKE1YzsEshsSOt8hRDGX3D5qSCUyqE8z49z
MscxWDLTx+OAWZtSTxRZNuoukJ5ovQQVZ5LH0Co0ZAo6s/DNa0OE3FyTtwvOvcit
BBo15Pk+3ZI1FOFTe13219nvQOO4e0voUOJed5bOU2cVcPVFI42GfjpKSwEYLzqA
pFyDCKGIE9OSFQjo7fz9hu6L8VFbQ8Fq9+UC+6iw5TQxfo/uSc3arXnJaBlaabz1
tnJxkoMjSED64eH+YH9m+/6LebcBdw0/ej1KWp0QdMqAGtTrOMAU0zOQlYdLSxNR
Y8x9Gxvd380wmxzn/yOQUP1hAm9dFzP0HB4Y5CwIn62ZqZK0DpUBavKat/DgXPfx
zwDgGKrsuxbidFGiA/jpbm5cJ+5OSJoEENWfeDXBzgWpuSuDvHYsfNUncBJuFpJK
MYGP7rhl0i5P8QXTcQ6W0mzRPthxUw8tGiE38tGzXN90VZbUH2tbNiTy1X8QSsdF
iAYp/eHPhYRuQInhU6HPfsqoomQFwxsfde3tVFsQTPofVwCfCEvKCaMV9N0KaitK
66Ejmpji2tikBjjWpaqjq3JYhH2fvuK/hD0xMXfESS0zP0rGSGYC3ErXR9yWNKVl
LobxzYRIM7BfbKChtR+/LHfTWXORe7fNwkIOW4WS2FNHoYGCwvr+ZmVswGyB85r1
Z2jWKtG0MoPmgLR96mwYNubK161tgZljZMS+613fa2LptTW2B8r8LgTtOo/WioCQ
IURxgmRC5FXPIqDNKDxPPx4nOYuLlXB+YQ/H7IDjYQype4Ckd4+aKDlJa/6bN0Dg
jtI7NqXUofU2Vs9KH8eVQpT8668MK1I37U24hvpWHrioM8yV6TlMhcCyHgal81Lc
3zPW0J+ruqS1JlJs/RWYqgRgbqlOumLsyIcNbQOf571kDK5peUihxUIDa2ipGgmg
j5YTXFacv5q39NGTo+LfbYkpHdS5JMSJrrRMxWFKSn2oPmNKUv0/wMfgCbln2Hrp
cGxKYu6+jBn/KFT1UqSZcL2wYi0tfS3+sWOm/DibsO6RQ2iF46Fy4pTc4v9oxxc/
7F5ILAiczmJ//DUsa/zBD730Mzswfj7kRf67tpIRm0VFreK9TCxrEArpWY3+EjLr
F6+wVUsjYfzU2uwVyHOfInytbo/WSqmYPlrEtwu1t/nQSZp6P3fF5770nz5wtFez
SYQkMDCvV8OcSef6EDHTiU0GouEO4JwcjGdHcE3ijjqk8IhzIvYY54AdLWkQo+fU
XjrBJzkk7ch2SLDefDjEj0y+nHA9vGPLZnqPRb1rd98AeiefZBwddqUC+/A5Xhnm
a/91EyxKBdJYXqCcGlZ/HqA0VRsAKcbe1hqp+mxbk3rqGzPTLG6zQtmRNZDx/CDg
cYaBC1QWpbqpQbAr5amGAF8GdxyC9rvvh8D0QiQKIN4FQ9mB7i0jqLmDYJM9Lkk+
70vQCNCxOm9zScWGRl0oTl14+H0Mvq7IqlwUVIfVOH0ApTfAgRPj7ncrzXTBApou
Tbj5f2gN9cQfjLfTYyPkfmXKgIATXb9ooTBiX0vGvsRpvAWHEdz4/Ezg3tvPJqvs
8MTTPR+Z3OC0mqUtqLLGFM1dSinbf/TOGqCa+ShIam+co3DP7v79Ey6/vySaL5hG
anrpplJsWO32nnZtFnvFvI6WwoDGRxORXGspIo6MbdwTZ68b5x0vomGb4uvdlQOK
YnNxbz8keCh5JqjsoOqQ+KZVW/EWNdzDBbOhqPm3fqxRp1KSRzDl0YZpu1Zzr5wq
6/vEAl6b/k5wdZ2Jxb+TJrgNpyr8/G555SPL+nGZFqU7nlOOUvcBYMQJ77EvFneC
6U94LPTdmwOZFkJVaKC3z0YPighfnFSnhayIiTngEyi5j86M8WVAOyF9yDbFHl4j
9Coupx4jDpC1rTiqxDoXLGE9LZa2vjaetMnUJnr/GY09tsfVczVX4IlozvNtSQHD
+17pZL7z1h63XvGptg0bg6xpeFSV6REurRo872VRlO3MA0SW5/Ifpz4HmzfJDhou
CHyPF6bMSY3QM3ZCWwFJEBhxmclcsFeDIgXzLo4/jtMuSczpZQywyao6t2BEbDPi
ZUQncYI2LBo93BVwGGmvF6T9daeARL1NRASVkAI++KdLcOzX3rmcVjxD4mUkrfl1
60FV6BjbSB/aXolZhoqAai2WghSEpiWO3GEbK6y7GrLqq9StYDqhi8V0Hnzg50lN
wZ6uYvPei0IPt5Y+IaKra8HEUpte8Lh5sFCeohmjLo/OcHyxVd2hqJjkpXFf0Ps/
O5ylbwrQy1W7smBlaYC5zRJSNTWt2cJlHIxpWSfNrosZ5j17UwhrbYreO1h1b5Tj
jSPP6bSblVlwACwl5uS17VlVEDbejUfwC7uth+6rUjK6KcI6cmZIuXP2F5kt1Ehe
l2ophc06ZmYc0kmQoHG9ww3tDrN6ewZxJGALZmLSR5w67qQlrdTHZxE7zait+AtQ
1K1lRwKRNa0FpPmBTmOtgv/JJe6mG6csXZzTB4/Y7JcsR6mbpJiSOkmI8lsV4Qcs
wGQSxxlICauIFs5yZfxAgycGvgAWOL6ed+xjEPKjcWiUvSrAVsby2XUZSBypq5EA
EGe4kpxZMkJ2F4Kow8GquYJ7vlqy/0iEN90XeGVwQu959g5uVQRvFAsCUkJ6de5D
YCXjV8o+tP3pAzIytkk+cJU2zOzR97RlZDebPXahv7+e3XjTLsopJ5gSykedgfgY
OoGWQ8Y5AukndN5z2UGBCSF5Z4NkmS9EdcJ4AWaeonEJ5nXljyX2XNSmYHmel02f
etFb65M2UeNQx3JDyA0RUFeD7HvuupMKDxp3vIXu6ubHjIKAKWp1v7Nj6Q2CjOs1
OyXLnAnxyNnnb+kfi5EXCF8d8/lhhktnqE8TJ11vL72laOko4ktl5IlP6vXAfH49
L9hjL8v1xDFsL97y6RB/fWydXcVVSKTkL9n7IPFibPLZw1XVyTbxPWn8vp0wADb/
Yq4QGDLOBDxlVrqlNIA975lkV5WibH4x8rIx1+yDeOMlwFqZ3B5cCsm11I292h++
T3RfHnFOaQVzjKbmZWkXHAeN6UJvTvV8hCCVnGf1A0nLWmS4j++KCBDTZPJnPjqE
YvsIm/+MbtE4yViuDuo94QG9T6fudV2+4OxeozOeB/cVxKlwGG7WNg1ceJUW2007
anhH9JFkP4wFMv/QRO2r6N7pQv8F8jCLA3n4cea5bqx7Q/ojbOg8/BgmoRxl9fSp
rMYUuOcVYljXesE67QNJ1FrDCEU2H+9P9cZ8SMzx2Tr2/v1AWRRwmOG7MaWLtBjD
hrP1ljeO7PHwzFUtDmu1dw4MOPyYmw9wbo9PFmQjAq0qcxtM+063XxXb43T3/AiX
uDTIFMZnF5boLcEPYvmu+i6CadctXlVM334w+QKD0TTeXZ2OwZIAXthLRvREOMJE
oCAWu5W/Qm0NHSXCZEXFYvf5k+FWI8C3s59jeeZ3AC4mDDS6GBI8/zyBKK0jXrrl
VPPSISQ5dO9o/f1vhaVrA3flCtr7PpeyYtdmJz4P63AN/GvFOTqYES2veeuK2P60
3aRGdRuC08KwDDV3gFqMWejbOqqEEeG6MEOMDws8vXjHH9eDUc5xVZ+uax4k4TRW
CEuQHxSpm+B8R9uGt7JPhdtDC5GPIoMfjjWYz/dPmAetpqi4cgCvB10IUg5pLJrI
5FBw0qhEWuOG8XM+Ec+QgnKvOO0CqXQpJdkNQsJlfOerO34fEdSSHi0vFq/SEv3O
45ZX703A7lekQJKn2GzeU8DazPX8tgWvBbsg294m5McC6lB5P6ME9A9yj2gBJaIB
bGqlg9BUEGPOZ2Zwrr3u17N/MOe3t2S9TO2mwv/n+spoRHPNDXdolE2aM/AppkRp
pQ3jTYRmODcc7Lhynbke9Jvr1PmNN5kQGUQAHZgN4dUofD+lAmNqr8wmkQJLOT01
J9jkKBY9JSwjqFdTECQnbfkDXRn+iJdHRnnBz3JkqdRiriO61Ipd8weAna+kbViL
dlwsKHx2ZHKGVxRi/R/X5n5QQb6/mIIy78wMsfi4eRGqmxHf6syx68nnJf6oLg5C
WH/Vijx9xBEREpysVvbFij2DVJ4HqR+JhCEJHqLk5cRvZOvWUk2dfbTdHnFGoG+E
sZzxSxKmf5AGsdlR92R3iP0zd/vaDj0Z3ZU2U5lYasVZua5/ugIme72iiydajniP
WOlpZ/IfULKeWx+eVz8ZbitZZQbNIcMdKQvnFyLnYLYTZfK1uxy+rBWOvU33JefH
kpr34f+Wi/DetY5RG5FEax34/dstN5vNjJp/KPdFf8DZHDTG8EawJUfWqn3IL+zd
rXyRdwdBkY2DANYKzjrrlSNjr0hmNhj4b+AMu4hGp7g8TShqzEerp4rHwDOoMYUP
Tg2KR1QTyyujShQuVWJgsOGGyUCLHo1gCmZWSfPeTvp5o0Tb4hkVgIT2tQBq9BRM
++87y3ooh2UxBjz/qmXU4dOUNGEhcDMNRuZ5EYw8Hry0r4YQuBK4NbZxcBfZp1OA
4gCQpD1jjCNvvFcXvL/aEO9S+h3SpveNWMq3XI+NMF2wavW8Yk4h7OSiGLO50VNe
5qJWhKPfvABr7DzBegWSEmISIYdrEbdKEQ29oDK4oSnrOilUkfTteGeyixagIb3X
epna7uOvxJj/UrDwl2S1zfXm7cOdGSdCPQgzczfgIfZz3JeFEsX+WT24mi58UxWH
AeWd4VdkyQsq0fE1rzXHwrgjcVxpioohLSPt4CrDsdPnu4eIRLzn6quKaq0jqqj/
L11mUAtPQgtD6Vavms/CC6PWLtRJzsmHJMdIa9kfgon035x2aOy2hu9jnPb5YQdV
6E1BRIzYGhQGiLJUsVcjO733d0/7g4JXCXcQC4kAfwfPOVYDzPzMb/iAZP/Fgk5u
hDCeaLml/EsjMAWnsJjZGQD6K32prrFZHwmwsvwLodoQ3UpaY/9LGLQ5Yu/qDoW6
sEKenhLpaeQXxFzHQK4y12/LzRDcQ5dKa9gfiduySlgS7TX5NobOfkgraBSnzWgH
XtU6VJtLHkJiAbFcVr3wA+jIo6yFynk0QiA5WflnqJ6kuQ1vXZ3YVwVvbVNDGqas
IqYbcRvvWbOcgV7ySIoYQQrGKakgOwXs+HdtLIpSJQSFQ7vsTVAz4SYQ0qwE1tFq
61ZeZTw6HxDT20fPclecxII3GNFu5yqdOg/iPDpjvLIWF0qA3F8hO0MaxaQQLl34
IqMm/lAhFs017Mcwhh9PeEPa1dwJ1MUNtItGeMKtTVZ4Toa1damjCmedh4iKMt3P
/YZvd48QZiQR5uHKcrIH1Y9T7Q6pKs0H0sxq/8VyUCHJGrP11oKx4O6Jxs3CHNDN
wpYjddBv0pwIJIheZlALvX6dwDWEiEMt7l/dSBIZV2Q7cZHF+Aso1wi3kadb4aZh
kuQAiMoS2uIwm/HEPF/rxPtsQ7uivLM6HV6sXriImfgOoQl67a2xVSu26Vr1ADwY
VzEh2lcX+nsfv4LmJGmiw23Ml6AiE0BAl2FyYUhpvk/9D7zHa2LRJ99TSdqnY2OS
DjDygx7R/rLD381II5eFBvVtpB2XjWiLdq8sKOVKskjk/lCCyf6Yji/ZFAgLNBeB
aHzkLleNa3ax0WNH9+bm+DB215XtJqtSD3fgumEEMq7hi0C1+wPyVKkaS+XvCMdx
qXs7VS5kE9WqukTVU14gaF8/uUBLEAS6LRMfoWg2eRXk6Z9qvQqLwucfhAKC/tYU
HkAc62yBzZuONy1evRYQ0/wYlYble9JFRFz5/HA2T4TCx4z6jL+ZiW3vCLEk08zv
q5WyzX96jULYgO6vCdoteOvYJsPYTtAoPWj6bk6ao8VnuNlAT4AILXK8jCwLimtv
sSI2PYZTqAxLMutVO2eEXZsBQcanzgLaDI1Ha1DNp/nYRtF/L8aaUOVGWTxGjcJb
s4tcWG0n/1kC3Qx8+ZL8j3Be9hlNkqwagtqv06uAJNukAmr7C6irdoOqLa2oWHZ+
40RisUNhXgfvt6/CUugOGMCXs/VVV2GPy9xwfXKKurK8HOtdGdP15YL0/KfJTNgs
CJLmamCuQz5R3F3CXxbew8vNJ+kIXJyWns11BiGFWAKrKH7g2nATTdH+/29AlhAx
73ffl2hpy1tNANwmrhQCeXJ1a8l7/HVJzDuVjt9IfsYdkWFMP+Wpo5sHzxFddfGO
otsJQVPq6nMAOqMjVrG4tC3I53/SIy5BKxo8L1vqgX3GCTfAvH6dOF/4Twl2NFTn
d3hWxfMfdCEZ5V+oOyH+5cobz/AaGhN0fziPCal0IPTQjPQkyHKuctW15RWlomNs
iwF5SwBTtfMUBmYPR6nnvsUA9qGQkdD9YQ+fR/by27U3orFVhmqRtkx85cK3TN6c
RntNYvXE4eXom+StjAtX8UP0ZELaHowLHHFxYX6OUFHm7ZjBOwfTvAJTvq0YQriB
yv2YwGEZvzxbYOWXxwSoVkQD31M3iQhwzz8sBkivsWqOZAPhnpd6KE0sRjKNovjN
Sy5zexCyD5et8oTqH87VHlrFZO7vgFwbA3meJr9HbW0ec0A8WU236Vp6NMOKZcad
+z2VDC62hH7npV0JFgO3blDp7Pu9K404gHwvPYuCbgI5INlwCsrdOvwhVjAfOD7x
q+P3CWS1Lywg1lCLtHDGCkFqOOa473hRhQKpLxpBPsrnBrTD5jntxy09AzZRHT37
yGC/ydnkWJ6JgchSmuwUSRPFbkL9HSMzDznQzoZHmAODWm84SNHfiBqlObl6L956
GbuRu/UYt6PjjUEoNoAY9m/JsKzJusfKmrLS9ooFV1j3D9BnrdDWE+hR1Da31pHN
B8vXs7mpd8mtcJjCikRVWM+q+OF115vk8nXy53VaooSgXZSA7a1/l5QmI6vVDqmC
WhIZXNp1mkhCyqnnoD7xKmBfVfHQbl+cwLFdXdDaSLKhfkLlHThYSsrX/hpdndP8
YDHZJ7IOdNfISKE5T+1BTNQ3deMUAqrOQuzjRJy5aUh5s7i1lpl3AVJb1NchgcMt
ILKy0eQbIaEKQE/JhjZ6ZP1c/5heXMZVc+agi3/rmEA1nIMa/0MWtRG/ZYCQeJH8
tJv/Zr4DYLU5XywsQm2P4AxPgtewAtfMafrSEMZpRWCNE2WKwWXC+az90Rv5nXCK
6JAlYsPZ8cDlthAPz2JpykoKd8TkWQadNlebapJDdbzpeMIzIhEQkJBcptJZPJWm
NRL0/n1jCzIGGFABIK5THPvm5fwaxhsQnOzZWrDSPaFh7n6VW57VqWBKLkZInpPc
+o2Rm3ipgTCqSEVRgCYYhRm3gWLxr5jadPKDyZphiSLk7MIi21spsbpyS4kphY5G
+qJvqm5SbXvp/5TZ+cYfgiyLN9RPc6xBY9UI/umy0EonaxU+70VWg8CGLVHcMp1D
cc2uRCjBN5fztoC86I5Kce5GapRfsHUasHA7wgoldHAJV3ExeosghglWldYF55YR
rsEGdk3ISCSFQswt5nHoU4LKXSGL8MZoj2FQF19QJpxW+XjSEpctmeyvHGr/jwru
czsWGB1HvnEuMY0GVxBRc8S/MhhEBJ+KCfk5roCMW+/K8VF+wLc6FWXdWWaKEm5C
y2H81wQgWSbhQUsMMh5FOEDb6eyp/QurPLDseM/I0COAbUsN23YGHNPWGVL6Hf6Z
nJJJQk5F5+0GW4W2djbK6Sju7jttnPFtXxZSxhvNEY1RVC6hhMSoVGaNsvsjQdHY
vpcnMkSok+iBqNmrq+fY6JPYPNt6V/sutXlQRFhb5zdc+rR0nuM9d1llmrf37+xa
q5fwpbaW00F0fpgPZy4lzHPcVvZeAMukB3NiCzImhPFZE0kBS2enVQ8ehvM7Ed4S
gjqG8hCJR3T+6CejICwB9hurdzRtxBbw4gCsbu426nDbnq3PV4ieL7RKgtOrFSmB
Zw+jhNq6aaxIoemghxyJCDtM8HXeEmSqX5H7MIgqJro0VHbeK9ch9mfiIa+ABPuh
N3Sq8JrXSWowHWRebNDwm5t7ttM3zKSTLbIRx8Fsr6aipMcmJgiOt5kIAA5GoFJ3
KR+KnTPr5cQVMEcn3CujglMRkVr7hUQfPPznJIk9kOOzBM0YIIzzVX0HohuSrooV
xc4b2Te9QGKRKawP24UrdJ+IDZ/Wn2RbEZ9YirRiWvAbT06nEuGyZLKPDbKlhaOk
rum/be0NNe6/6us5YvJ0/VwlTYMD5dfa4w6NsRolvqZJqr10Gvs8owwTgolEF0RA
f/ad7wjW0hbo9u9CSM5q0Fvzsv+zQz6l58QVlO8SyMNH1tSgs6ElZ+gjw+EMl4sJ
UzgakctgfGgRKv4yaKT4H9vKXrunsEvi4EkZyi+CMCpXMMDXcfvnAOnWn2vX8O6r
pw4fDjO1EdQpI8bf9ntMsU5Uty80YRpuPm0r3ZI+/gaKRcieFaCRPiyrzcmEscNM
oDfCnzVn0/ZtNb6sRih+apIaAzCLcv/7PsJwaxLDF1E89GDPyCe1nczHbTdZVSxe
K1j8BtAYf6sA6H6I8xTye3Hfz0yZirYuUBpvRiWI9Wzw3aBmjTJA0qo3+vzNvbQ6
WsFg0dzxHXhafeg3wQ70XkNAEf81Jbikyj4zjFK/5LYzesT+n5CpdlHBGqHhR88y
KGig9fbijODz/jXgiA/b8f84UeUUJYViRlq1sdBXSSmPC8Nfio3qxuKy0vRJNiLS
ZDrBaBOtZTYXQrnBwYNhEZvrSnqPrFGaI+25NMv51cI0IQo2a6kHvfI5gRM3QZif
TYkg8q1DQyCRzq4/sg+w1yZ5h/UwNOnVod/C7TWzoFArty1bMQruUDOkQrT/F5Sr
H/a3YLcWvipPrOkm9vvrR0gJQrTmPdsT73NNSxxpnOogjWiFwCpHEfRdxPYUF4GJ
HIfGmpOIT973Auve2GDx4+COCGNf5CrYYmwQAcxU4BSyfXvQKCTvl5hGElxRI27J
cAMl2zZrbhuuOu/fCeUSueodADbN1uFScfzZe0FxwVd19zBiG95UynBkTsikUZIO
o7SH7ZO2+JpF4LxaBkqjqr8I7Vlv56WITV46Y1AKem0wsSW4JaaChtu767DxMlbr
wu8tPi0A+Xqan+cFlY0ri7U2SvZz6QbOuch8sY8LjrfIGtuxpDx7OAY8Jsnvts2k
96UTABd+dGIOkqw6AraaX10weHrDBDFUDGM36XFITJODL4DgLIFXQFx5pHJBr6pD
k5LQeEr1seaD3DMVEka08dzn7vG+XYGPWR/O7GZwM3iI/nBI23B0hab+0XaCK/Mw
AxfawqScVCBJfVpXyrZe9Y6EkSNAQlCMj8lNnTleQS1+pN8ZKe1iLrKPoh55PGXP
WoapgxPItHSg06x6aobbP/aFq38tr2KtUUogPiZ3keCVZNs0YnRJXGaqEJM0b4x+
EUrlJG928xpYOvPMMm3LgaSTf0ofBRpvUThycA76Iglqmlmym8mEye5M/saCwW5Q
5LKGVE86RxExW+mifLBQ6X9y/xOugM7CWYYBBvZGq1W+kXspqLaMu1U0Br5WlPny
dBLRRUpQGXFlQuI5fLNE9OzASd8hkxFJMqiucE4wG0KWTdciAe7h0JpIIFeuB+2m
qg03pkFLxgY3n9lf/Ecs211JbAUm0bVl7nW12Q1VI0qBv5eKlnfQA3Vt/Ydfs4qS
4RZpkEV7cE1/orn4JqOwZmqTpJmAP+m0B07VcecHADxzjZDpra57/4PTrZ6EhKwe
0nKfBknW9BUAI3Wcl+GgHW/MNuMLi6hcxxJumfdhJFSKpnwaZs43b7teS2Iuc0h1
cL9CdDoH2Ggg+aPIjEV/csFNOjsWyV5qTjeRE4Q6RldANO2q1Vz3xdz11UGr1qvF
aPf53fngZzJowvo/y8i43LfNClObgZhPijw2ZPdOwed+e0zEThTIx0TgUD2xqCOt
3V16emNApLrQq8w3TgDLaRbkJUM8XyxWutlwVe1OykYqkr1bLv7Tt1pWFPlRSrsw
z6myUAmY9J67kP8rm3MZX+194lTeUvfKRu2E2IMFiaGWlFihzuhBLgJCtjhc0/9/
EaR3+EGE7dYMUpWedVVc0zokNE1uVMPUEUmZAOWNINumxWqr8PtMJov+h5W+whAA
sn6KvusxEzvrb85B0DEbXD4S+UvZ67vfji42ZIjN7idzsOgnu49FymfQX8Wfc15Y
1asMcZ0CF1i8teQPmHK2ufGYbeKh6Gl4JGm7Ix4yOz11jEr5Py5yNf6FoaDWzhpQ
VXw8kz+amUiRRRnvPX0FN+i5yV7T9KOuaBx4471aac6K7IOMIRDDPMoL+I69VutH
ShTG1aAwn2N0jrUZDRjCwQB8F7geVL4k13dWmBYkLrUZJxpJtg0HBhDsSqSIRs6k
+bq21rP6VJxx2ULrFFyWMyHVj35nD2NySB7B5Y4GhdOHQINjutWzoxAXUeevoko6
GdOEKq/SeCC8Zl4aEWXT0Z803hxrsnYgkm7nn79CfKjmcXmskSDRMDx2rjai9fQk
5mC2haJ3+VLYuEu+7qTBEmr66eVA6dN7J6xNYxL7zylNN8VcKWFhs3IA8Ybi4oXX
C+OA86ZVsSQh5CbiQh1AICC+0Kq6IqimFkShkR18RzdaxalMkpaVOz29xDYb6jYK
5+3Ns4ljqoN1uGfOJo+zoZIAzoM+XGYWjIzQdB+5QCpdyxz4KGlYGj5wyHEo6xIw
ltdW92ZrXPM6oxN747Zh8MKdRFiiYOcRLwx+8fAuu7Kzj0kLrDcwEZdBK2E/CyBQ
hY+M6d9NH6Vr6XPBc4m1H/mvvYkEUAVOG6KIzDTeiL6mnSp+tBqqx3/B5tXca6Oy
pgXPDSFWX9z33O6eF/umeCV0/PO6wXQQFsh7+pUHeViaKvp0hDkVYBQkOKL4Mmad
lfHz0NGWtkjZKcV8YQu/jlwDA3ZeNzyV6v8e4vTVUx/s/Z7gfz2Z3ByTcicSMRG6
2ice6rEYk2B35icJbhziekG0Px7YOOtRItZqmXK7kQ7ZONkb4bK35RopjxK/jtdt
s1x5UnYiJhs8ln72mcIWCBFvQCmq+Kf5ODtOJMk8J/w8ccowvpp/yRHiTo4EuseE
K5cKwjPjQmA78GmX4mpVidDCDMo4vFZeKv41abq1DSEuUNL6a2MLQ9NWBPwdocyY
bLXBOQSWzbWfaOMh3kZkFns8EJphlFn7+IHFygC0wevenwD3xbzRYJPN3+LxQiNX
kMU3ku6SKGWE+C4zfse5B1xV1zNdITfiLp0AAmOWOvcRUUE9JiTnncRHaJKAQceb
0BxOqK6u64sc9Pq+irW+Xm+gEreghCqDu3BWrP3vlZxuXCd8aWZoVG5Tbsre3rg7
81YOHnYWtU302LpuFPWPbvosDUo1YwB8ONYA1Fufjn4nIRHuPRi0BKv4+CgJd3Jn
OF07udH7ToLL3NJCF2ZhUgOUXsGa6NQW/1Lg3rH+b7VaERMdrgduZlgZiyF4QXXn
aaneXd6kwIKw5YOuZS2sdcjOosfRHIj4gyQueXS3AcD0Vw9c3VGgq2gF4aMDr3wJ
1Sj8CzF7nhUJttjVU0qjBujUXRklWHkZeGIZDN7deQO72CYz/jPy6PrQwy1YKGej
1DborL+ai5u4QHRkiMYYgMYs2iswdlPidCPZCFjKEAf2j6bVX2cUT4QB59p84y8v
VFX7GAFJcIrDv6psI+VxPJOYU/8qD8BcnuqM8ryaPVi5tCr6TuE3abEnIiPuCVZA
M3hDzxA07jS21+OiK+RSRVp12Z/RJzNs5yYNTbi6KU7V1Bm3Gn++GhbiE+1K+BhR
3ELoHp+WfZ3qkDKd3tCTxOygmhZmDtNnPvZYo8ksycuIgZ7yF2JT+lcoukJaE+Zp
8gipdMRbGaNrE3PVyzRqWKj15i54mD9GptKSFvaIjcTuez/JxE4iXg+F9p6SEgV0
u0mrHO4btGFmCsY7VAsJRvXKRSw1KgQDUiPirVjl6IZmuDjebJxd50q/02BjTTX0
3oOK/LfwRyvgPBS3Vg4Vt5FLzj70buJxJoLGI8IpKiZKnQIC7RirVMalGJGsxG7/
FI+u3XT0IrqQ9sxWtotS8WT+nrYBBcYVOKbHUusQht+lIaHYI0ZjF/u8nfHQLz3I
vAqOfjjhYE3UJuaIWDGkggsTIC0z9OYtzMGV3LGmuYP1NDLj2YCmYlogU/AZ9qhD
4BnA51A3yTlOuX7VXax6+w2PAx1Q5cfXXaqF0hIXeZkG8irsz8gN4rAcawdlQMbF
/cirsUHbs2bZs7MeAATo127d0X1y5tcWlhSX24PRQui0qO+T5FLAlfNVdyrURP2b
v/+4vjf6Wn/8ntNeLrTNWrMMOtOaBcJr+fxhPfmkWoePoNnd9j0TcSzxnwvnz+TZ
CrbMDhL62pAbCc/YfC7LCfpELDGOpO6djPhTbzCd5WbFcWGGi7HD4XvRrYqSRmM7
0EGIZGk1S0Tf7MB74c1JqiOsEXn5QFiUfG44fvYXVcer5bI6RKGWH0/n15R8Uh+R
LOnpE1s5j2xsEZVyI48CucTNMsYaMSjhhyyAy/JCCfIvOhGG0vbWi9NNfmL98TS4
ExvgsEMG9Rcf70xZ2xfg/myrROjpwcdEM3bCK9u5iE/dKgqs57EF6gnKqvW+OZg3
aIzcne9iS+uCvuk9k68NZA4B70EsSBSZ+BiTYrFuffnlat+JWjIzPPil3lng5/Nq
H7bcoXvI9VAhSUDJ+isdpznv3T0GU385bUBsqI/O2BdjjhsXZQ8BC0U+z6Pgy3Di
F+1obYRp2SWdWnRA8WOIMQKu80oNyquzOGZ6Oiz556zEjEjC1tUFP9n6S6nsi1Lm
oZ4cQkw5t47d8ucMa/b1vRN/cXaniMZ5qktHQ1TdpeU3R0opTCVoUbPnVQdwZN4L
Nlw4U5GqoVlH3/XkHwRMHEpI9sByOQhrSfwQ+1CmwP0s1W3NVrjIdjpy4ErZnRN/
0zMOlSpmo3r1Y5v27DqTevfCjai7VyaqQMMrumnh2bL8Zfds2vBfJ5RK0miI2aXn
H97yRXyNEWefISAb4S0C3FZGx5oR2SSt5TfltZr36IPOcZCEkI3JEDYoyRzU4tug
OsEBkpuwJ8N7PNmu9HxrC/stJ2wfQDuh2MUVZT9qgSUoymLN6jwgllhnt3m993yW
1U/+8jZwPidQssi64ydTyslp7W1S9+VyQie6Afqfjf5RsVMLb07Xi8LcRJZ+jz0W
xH4OB6BBsDED58/LhvZMJU0e9RqsnwbuPynuMJeJQk0I7liPTyghs4gaYfCcG+pv
4ErLjFzRH448Uoxsx5/hPwngkhyXwJL4IEhrm9867VQXS5Qh0XVo4SqCzGghPaff
qyIfYRR81vywIWz6BOPbL/EHbiXFNjNZxMwd/2/rq0kzrG9YlBu41yW8zSrMueQP
7ZGoQ6jakixFNAKergkyuEhDfIpCJoaE5OVS8TujKI86C11gGwK2EBcUG+9FUqi2
w8xefqQwZG6oEAEGhcc8eLcat40c/j11sVDIdGmy0ilgFjJ4QQJ/5o/aERiuypAl
7xUR9mkKI4lLEa586ZY+wOtUOS9hwW0nzty6YxtyL/YsI6UulQ9QNvijg1ubVitt
PfTx49JawWylxKCXAuUbqlgcpWBRxwiXo2hxgvVMZq+/8HsADgQetHl0oCbiBw1D
ScmUhz2jGn4K51PXbTjQ6NvS+dAfFwcsoAXIw2mwHPXOEmpgdIoF689CLfClgke1
yUmzrUs7n7pEfrJIFCBBNlmE52ZSoLm+1Fft9x6/EVk6o7d/Pv1RbnYnKLIkVUhI
6oK11TL8oIGXdJAEO/7rT3kmT9XJQvgc7DHy8BNDIljMschiojjXK6mUrxZg/5gf
f13N1XSF2+/k/hNHrfQFngUtjll/i50jqtQBEFyuCffSx5vnEog+ppGgDfMF4eAo
gqkq5+5voJW6w6gzUqtoEu9HGo1+T+ddAZRb4RkouOr4ceQ9265jGy+/e6jiOWcw
L4WuETvg4YnKQWEJWp7LiDpbsQZDUdPdhWW7lIdekQdSLeQusqMU3sK/3STPEZI0
VKW3z+CroB4fiAI6/0GNYkrFOcXHnPwe/g+211NAOPgo0R5jZO6qhgT4NzlLHnCz
6drD2qa2mfs8EVBjgPv6mALOFt2fxrDbibx7h3DT4UMeNC1nLajZPtBHcWDbrZBX
joXMfdEcKOAM3ln/49TsUqdpJTt/Ivsjyl7DsAI16Uttu1cMC+FErwa48MqQ+aiX
J2hXLvkC+W6yg1iTsylMvKFFPs8TOsGqOdha3yN4AiIupW1y5Ivb+71hl4ynZGws
R/5n0neRAZv/aboskUoUXqENsa/Vssw0CV7m0Oz7Pss6k9+vioN36YTy43+BNjWQ
jf62IzY+AXicfeuTeopWnz0HLkkSZcvvwuy8VYIk7IE3SYlBGYmB7BYrMwaIG/X8
1v+XuCrjReUyY/6arqJi4zQ5xbn34+HAB6IY328JhlrsfWB3kE9UDvTOFuSsQaMY
xWLsoYW93woKEsVljHuQWudCdnCg07ZxEAsPLKu+9hOPu/UrQfrxaWi67Au7oEGc
ky53+gNRLSR+cBYEyOiB9oW4/cegxKcQaibklVPSQZnPxfI1bdNA3AIsXGVa+DAo
hqhoCIKfsIHDWtj9coAI4yVK1qZMDjjN/X1dAorK2oS/RerUSGj1cz0YnSq1ey+6
i+JbhfPTa5INzvGPySNQIDFMqWaNhc7ow4LiEVyLX9+8QT+qRFjgDYNDbltt2Q/M
PNBK20H/DnCP87sUZKpBKoUmeBPuUDUHSMgIWocotE3PnfbsRRg4kvxQzO5LWLJY
2iwK3zJW5e8KbjQy7t/A81L1giaJUJNGiu7gvegm+8vTrn1vH5kY2/2aqzs/kxJr
tfyF4N/JnsRJU2Gv4JvKiFAOsZYdWmx01zu8LrECRYkq/0xvP9l0rmYj1/isa5hD
32U5SLwf7i1jBTz/Lr2TremOYIIvsH2vJWft1K6Cd0/4WZeRSR7E+ogIFmSNmsqR
+AHoYcr8eAeTW+J211DiO7MVVpy4VmbvabJWf/A81sBeEbjPapP/Hy48H+nTAc2l
5/XHhQhIf0rGvs1kRHjwv+m1LLDV/xHzadTzBwhlForSA/S19+P2pkFgyMuNKz4n
POkZqOAoyGMl5+G4Z5S+bN1s+zI7OawkAJTS5IrFJ2FWWiawAtrBVuDAAT51JFA9
K/r3jI0w8XucPbD0mom7J4Kxk1SlnSewCkwwEm/FpSDGjPcWR6kpsnJaQ4iTpsWJ
2RX7L6yqdTjxE0Pc/Ia5Pwr2IrA5jPNhYNnEZdDh9t7TMwzqwkehhUUPN8OBB34M
rxrClR9plZa++yPltbD9LtAtuad2fnGJ+z3+7g9/YA503Uo5DWBcmzlQTDicVlpq
g8kMJ9T9pgiK4QqKbF14TWKQa6RQiyYNvpDG2Rxjkd6wp5UTrVWaKPQqI70/CYk7
Nl9fb83nyGslde8mRfFUJBfkJRev9NX7T8EpWJYjvOhZ/qTOZHQ052cF6Bf7kPIA
QbPSVzyefTG6tPQHTkY+QzOtolEjeuvr1rhx9FrWqqUV4H7STxof5SSS3tce8Ox8
AiZFdCJ1QcwSxmK0n+nFkOnSfEOfTjih6m5ROMeyKn1GmU/lNBbPDVPvYh+nRm/O
1I/wI0UrNIIiM9+audWKqC4r5+1tV2stU5/Lao2RR5iWvdKVeqUrY1OotNhsUA71
nGiAH/uFHt0EkEJUZZuiPvHCUYB2dZkJlRJDaIed5mAPz4FOnr7+OGOnuvig16Sa
kJ+Ld1kHyB3qTTyrpr2pgLwRf6mnRKDoxwFq7Q4ZiHjnCg/IgbUrzVWiFQxK+1Uw
TsneO3JwmAtmLzr9Pmeb2zZwvZDhJQU8tMv5zZbfmOUVEl5WEf+Mheacuha6VUuE
af0nppg77xHLpENvkv2CmWW+a8YDi7nkDwnvLTU3qyysFXuI2BUyAPHgZBXUKjdC
O+yG6c2exOUD07oPwbB//MuxCZlC7S9SlnvyL2qP63vdy417KQ43rVFb9uIOX5hh
hlkuwS4jAeMoMj5r7Ug9ReAqNBCfF6b4Qe+rNW+/08LyR/31Za41ecnSw0hT3uRq
c9+s+M04Uz69r4gwH3Pan90aGmEyhR0gTPuXmy0+cep7Dx29kkX61s+5MDsMaGJS
1xk6bevFUcg/vAhlPk4nDzRBD0FIyLCgY+uBwZ4iQjnGfHqTSikZJbZ35OQy6ACk
xHX4CrnLaD/PqpGRxTb9GoaZUGOFhjbBIoykSBYAiFUJYyVG2g/EXKRnsdaO6uqx
jLfXR6jnxqozkp31+DS8o5SE9hI5hqhq539babp2XiaZGn4Q84XOnuVL5G3BaX8f
wxHrdiqwo/R+dA83PN1X+/Q+B/FoTDOsgeXUuF347F5Z3lOXC5gPshQbxcp35qO4
/yfwkKr6LTuKgNnNPvIeELwBuW5M2Wyq6TXJkJ7pz5AG7m8eKXoYaF2M+mLxrI67
Tk/4GnTTWHmt9Q+GrvNFvFahu7seBE3fnGmt9whfZ+fsCIlSMAtfVfdT7mz3UnFR
TarqezrGraDz7CUaxjxbTBgIGPg24wMxQfY54HI17dJOb7rPV3kkUbaBUo5OD3zk
cQ4DwBFAiL075TRAgAjGUMlvfhvrd0k1UHjYTRQRTqnZrKwuJO0sjx4F7Pk3JcxO
EIt8qK6qgIe71JxYKaLxtB1JEDpxQ8FQi2QWw/EpnsHG9pzUVbskyUEHzxukfP5R
pqP3FmvYniL0P15BtilVS1WK0reAt9sIvEx5r+2yhZGJh67BzodratLLAjkhPqv9
GgHVAiHhO2ckgdeN2LBNoilhAj1DJFdCB6jNnrEYY1JpEhjTp8GrKT9l3SdIwwSo
oFM6POoqJjWm5E3FfkCWnN0HbjR6ey0R+kTgcVOUJ3aWI197AE2+x+pbuWN8Hc0D
KSZWuLBkTDzCw+VOaYh+1/dA4kAjHOsJwsDMHB4JMt5DkS5mKEIA3B5J4X3LahR8
zA/GbhoHTv0pbDfVmKFdUhARhQhfPskLLrNIhSpp+ych7BQszLmwG6bRPa3xeAG7
r039hK7gYB3zQZTo5121LC9J6aiPokghHfZ5ggs0VJfHuaJ4G4uFHJ6zZg9AmHn6
601rJD4qSw7mJU2wXCgjj3ruDJ4unKkOknqzoirkXcuE5n6zzqr20EI7HOREh+Ax
3XOexMHDefl9EED+tfk1sLrev/VlP+Bp8hnWHiVXLMwYvjgtVHeZeGvtzLHfGui/
4oWbYR4ma5P3Bv4nGuaeawPIggBp/P3iYUhe2wu4khmOvtQNqTj207+kTmvcpoGq
RrefSW0Gcbr9OcjLLRaMrMwlqVmXi3J10rIVvGwQvmgjcx2cyQqUNffNjrUpi4YB
5fnm/5FRs6ZEp8RrWgQZbpbUnyjpkq/rsFYSaQ+pBU6mkac3KNRAwyeqUfJrYXDN
jdCaceHECtLx/Gh+TToyom1XzEmk9+/7kA/KsN54t9HJCpDMQ+51X9iwDGhm1bq0
wwQxBePY++PtNPNaykEAF+g115txttQcU+U1zEY4o/Cze6U1Z25jIbd1DLrWHSOl
swQGVp7JZKsdtbeP6mnzx2Z/VlU6oVgEfFtBfZuar5OLq4Bejnmv/T3AzfciuX8o
aVlVOwkCF+NhNf1g0urDjUEjBetSkGRqfPYw7xQfsBR7vjrMdP25bb0Ussn2Iezl
OKmI4oUsO7DDvHGN8gpleRPi4TiRBxKx0+SK3iDZPedDmYcDKHsjUsZBA2vfvZ7t
BKcS3qDOLVwN4HCgxIFGdU4b/HjVFIR9hYKAYmxuiE0q7J7xq0cLEBkwCSxTeQtj
Hv58joZkovyzBg6p0mvL4usnlb4tApOy6GPLOTMN0G/Cefp+knwCpw2OM7uTM96H
0aS3fECs4aVNPLFgUKN9G1IXwVRDtmXUo+BV2muZZy0wIQqvENopNujv2E6J0kOO
WXI6lKwlU+y5IrT0LIJ6G9JDNce9lpKdoD0C7VU2UJRtLiTDlqNzAvYhnxU1s2fV
P1BgGqZ9LFw60WNUWQJ+62Me28W1qizTzJU21flh1y4YZobvaVw2Iqj0e5wMWmV/
y3czZuFm9ub293ZrTXL6KPeAigMvzpMd1rRF6gJmr5X5GF81NKPrTXMWf3QHqolg
pR82Ftv9JreNYzzy4VMyyBIwCJ3PQHGDHTQaa8UYX3iuBaWv3zNaHoKg2/yjvyDh
Y4ePHL+TwyV4RL6KgprYtCHNXZUZD4l5o6D9dJpWEcvhqSZWPvyfACT/wuWKGu09
O20F1iuaWHtB8t7nLMXrfIxyGhbePUxgUmZc6/1Yw1dRIq0XHnT3wLHYtcJptIQF
Qk9PHuOs71Fr/4eKG5M0im4Jf0/IVKxB31Jykrdhbe3HbYHQzgV/S5TnyckoFz9+
xyNHEDxP147DYdsJc4iRfK5e7qOPy8FoI4Ee2IfaGcGMk/dBTgoyQyaNnGusZYOZ
/tlp2Y9DurcE/YC0Tjz0jmifTwfm5QuUvhR+rzvtHcys+V5rko50nWQbxP4D0jmi
AqdxDYgODomKXxb4JXpZ4dA3HohAA3p86MRSouE3ncq/r+tkCmwPKQqU5IKBOo0r
K5Wfz0HRvX9MNsVAFnLnFi676Vx+2evrLQ2KIsl+YO4OmxKrxcuu+7CX6WyvzfuO
Fai+lyJ2R+clmsCXvXfN172e+saJMwhVDdZEX0PF+tdO9pxqOWIXwjyKNt9ws9DI
GJ+8b59enUA6JDS+lmXFqpyHugp1tSoBF+uBMcALSUrv2AjKoB23xbrwsOhVp46S
S8muIS0gqFq2KR0zk9bpwJUrGUf8uGt1UKCfxgEuPrhoYOy05bFMHruZBN1+epf9
ikhhH9tCfXiVTKqCS3+o3JVYsqV4D85Xj3IJqCAYPFSAws7gBJee1lHSLic2N278
qVTOtRr1bCkeD1E44zdHAr+WYXruClKKqvq741VXmzL2dS8TGh5THTiWGv9KGfrM
8a5NwGyxe0tLocAEHPxMX0G0oRTszOPdbeygSJ2vsv521qPMGG+yQFDuqMGtuz+k
JJR0G5KfEMwBW8lCl1BCEJ19TbxdyiWAU0eCqhpxiMaRZbpl7a6c7WUQ7e52eIKw
zmFwRtaBRcqA9RAQRO6WN8qKcbJX59iCOlhW2/B9EkGH2gumpxsbHVZPvI/oaoPU
awS9zphz0vNtav81FvPR1tTWpzzs02KExhvtMBajK/ocWfxlUbQuLguth1j8kbmk
J5I+E5U9vOMGTZJrlQXqd+XaKD+swlRnB+/ePBVSPx84U1+yFXkE/WVrMWKOpSm4
SMtd46qRc2AIGg9rUjslhX53FNfGFAns9G01tkrfSao8EJ8WN2vaYa5SY9sCI+6k
eH23TABSgAnPuLl13+UltVYkzlrI9J/v2YP7NqSupzIV+z13eS7rlTnBmSWYGKS4
48x3Pq4MUz+vjk3OmKupipcIx/WRa+X6G0JwE5N1GcqJ4ZvDae5nerpoCgAoxtQ5
ZGtVR2vE/X/cIfWQCbjqIMRcTu68yarvA3dMX4AduhymCB97IKI9CEq/GLU8cCLQ
8sSCibfHjbdc2qE1qJNbLDlXLfZkVRso73Zm8b3vGfN1MB2Kniw8CfcOwp6MDVTm
7mkzE2iMEfDoQeH9CtkzKN1C6ReSctrS+mT1QUOSk20xriTF7N6MLZjPQVA85par
hGDWdcFGH9l2pxZ7MwH98ZLkqYAIkUd7NCAshqwzqx6SbulFhdepOG9WE13YZyYn
5PutI4aGlj5SSB+VMHHD0CYsDhbJiF5MxT1tFCnvpETqpklfVNLcKayW9Mr5DnLc
sdfIJhOGNs+eiSrEYwDSeaI0gvQ3DudW+jlcpDLKSWnylim5FJCxNaVkkMq/CUgc
GaVTmBBE+iFMYYm92bkpvQZq0R1MYbcnVLIikDMQ6ZdJxGCgr8BdozdSt7OKJaaj
EqP8ezeLoc/xnuZZYqtB204+/rHZXDrdytycqHGWZUrNgvQ+js/go6LbPj1QThR7
znh/02ryfU6V318/lMENKumo74XAofPvD7yLSriZCvIHunTrbhnJu1f61ptyfsyh
G5k127bwcsI5M4R5GT9gvmevWrkG6/vljq1ZyepuQfPLVIHgtvGFRbBWGGS2GQsd
tRsSvSfnTOSK+eUZXS7crakmrH9ElAHuy3ysnKnL7DCBN7J7LCjo4jqFdGylEC8H
mkXw6Xot/uHLHa5jE0X0Ry73LL4fm2IKXD6/QJJVTnrrO8WjNj5L8XtrrvUrW26U
2mApDjNWUw30uYXCTi3lc2nX6hyykh3hk8CyW8LchxHwNHLh391Cc6RHpUSI0Wwc
gkAx2YHNO9N12C4YTNcBuyX8nb6INwY9gQ9yFgmGAw/eJ8+BNHYJZjoUdN91bQev
ja2gkX13ScM9j/jDeQa8nKOGldUd4Son+syZshIU7fPfy6x6VlUzZo3wPopPskEe
LxZknjnJHTzgKaUnYtd3CW/Jvppge6dUR+1f8/Vom1GKmaDbAev/ZAKdnajpWhnl
yNyfJhokuMR/qmDtuSWZ+Au1VGyJ2FKIoQkOJiSsBHQL8H7c+yQoRqcaJooOsgNT
QRWcluYS7jMSpRfTwVMs6xRWfdwcxq9lzxurQMHsSs0pUr2D1XevRhrycrsC/KOc
/eIsfHO72DZutOEmoPbZ17aNU8FPERU6Ikph57jQD7QBvXbWJg8ZvOIKCaEM3Ivw
mwt9BeZg+nWCFb3LqXxnuf7OBMw2Sr183cFDVVBMM+HAcPizPAEVy3QDuPRBGjxe
WlgIKtosvkZZkoizmJozUJHMSqck07tIcHZWiQQHaZ2Q9mDxdxBCrMHepfqZqN0r
Od+0O+qbNZ2ESpsX6MyVDuPAZyDOeMfC8SNT7Tf44h2eK0ZSi7RFW+0CLjCiR2tA
rFcY3Wxtf3dz/f2soHNG1D3c2/kBER4dTaeJSwm0BEconKV7nc9WeXQWg9es9aDJ
pqsY3eAVMQr5aH0sDeySWddoqYHswhr31SICgSmZXCd1dRTtX3PxzLsZFdwS63mG
4n3tllnXrWiisQbANax3nfp1jYY3b1mAMe2Ok1KOcjznNozH1KINk6khgOpEVeU+
FRnJxqfbFQFgkXXmQQD8cWQN+Zlfn+EjWWCas/jD1FRWqgFn1SbJWZAwcoLK9dzs
VySAwZ5IxlWONaOXm7arMj5vD4m/M/PN8y0I1uRZDK9Ci5svp/HnMWCcqe/dlNl3
DHYMXOY48sYAIXsJKiK9aXjPvFYah0APWM/va8nTly3sM241VOfSChAAhrzHLXpG
fhp9IiL3Z8EHaIdF6y2tFvs7V+oyFBGR3ea61Rd2lJiVd8/WZURYg0djIYJF/wQj
YgZ3bT86NHR6kJEULPdnzmoBkRysfUs7DiC3owrKAm00kzsR7DmP8bjp2E7wxPYh
UntyJznQ0bFEBrHkqgMx5eedCZJBKM1Mn8UDYz8oaGOZhwoRaGfFyLHPmhwQ8Deo
OPLNAIlhgEi1rSqBwVXEl6YGoJ3J6IrOpsEfSLsNNPvA5fGVxQLMMSZawBxRxDns
IKF2W8s8cnAvqIW0lh18ljmlX94OzaRolpS/F+8vW4g15Zhiv4kHYlNHvVD1xZbT
SgD75xLpFpDPwyvHRWmHMF/evShPMfaKQJ0aGgFbhGKLdv8PREIuxhg0jKdCunkF
3YJNp2NPUl3OIAy5L33jWvOumw6BjJmLpx/mwYfR5fiu/oUr0ZsurPNBfj0fZIDd
S0Qf1ssKzeW/Kal7fv+ROvnwlazbmld48aFeDnVPSnyWg8DtnoVI/gnyN4YYaT7b
irVZwJcT1pdEOU6VJbalVnA+Hnk8uKHlmyXgrefnKke7qHmOF3yjGiAWTvqlpi/N
zpWOAQnoOkXRQtd7DcBE19Oq9sLGuo6ClR0IFFPoLpwG0tqd1JVBFbY/yjjroWn5
9Z1LW0hUA+dLVfanSl5mS2Xk4Pypcfs1SLqWVK+SnjssVqqRj2t1JVg6G3QCf3Ee
jo85MGhux1XxSiH9kV1T7z52kn2BK2MdzhsgQyFOwf3sMRsnqrV9rtQOkVzfPB65
fhhcdZbBpkbGmxn2Pu60tQlLhgEm+GO7UyzOmYJFSBmOJUepDg7JCYvYU6P27NlW
TMcAVNM/MR2vNuNZBZXuXoFSUKE54y6FUJejNsASj5543Zu2VZTjTRp1l/Se2WF3
bE+Qf41rYUOr4xQ9EfiCZJbn4vBPNGPpxMJyIHrsmtUifhw26sTeDeHzs8ywUBCV
a/3XOCCTjRTCvhMTIshJlcbX6MSeBIJBFoKJ035J14/PrP5A3K1JpSDRNKFnMAyq
bpVdsagXP63d3eHDW2QY3b2Uz3wKyaR4xhnUtCLnid/1hAwHv/wXdJM/pIrXReTk
Jy4jAeDQqBIDzXBHSLa9urQqTHUmY2DcIbDQ3Vo0Cstcy5xcYOf4I/zX8D+aSHRH
M0+Wqhg4brstkBjJWzMi8f+Sp7oWh5QLsFW78lpYZIjbs0MWryKMatHjikC8Af3a
JtJrhyebZsXFMX05Wgm5nyczmeAZ27B9c+8L168irORyraS4vSAXT4yPamEmnvAr
sVlX30J69o80VMcIKSa11v9WrHBsXNwNWoJ6erlxoyfxhTelPwaprlfAqdF3EVNW
HkIOROyQl/98gGBU4ZNB/r83zrAJl659tJD9UwVPPG8FjRtedr59YDr7doTlu8Nu
vFa6PNLKhosTsNTEb4fn0QeKHWTOf31kvcENVD7yb1NSgVkbN+qQPqkcJgeDkAYk
ruxmvcOf0HwRA436qEG4B3xoyA2EHDwJGsc3LHq5X3fuySuy1QKZ22GOnli3YSb0
z6DoQI7nuuXGT+dlNF7XAfOg2DaRyTtvLGVS0jPopO0dLjLGTBg9/Kd77ya+Epfm
zxgB9q4U7mYKOkwXURK1Eix+Nr/WUmo0jJXEANPGD8TGt0JPNKGDJG8MwgaRdphn
ncksHuHE/v6ER2tFPuq6PBTbRu01Sa+NACrxuvBAoEtqy/27D4r2cCevevWLQpMQ
I7PP0lGg+LfU6+acxVxVET/UdlA6LvM/XS2UJthax4CyuSlueEaHu0pAk3D3tnEP
uN2jxoKUQDGovO37e+nWEK17Nh0vj43gK+PqnX0FfjVMklweKVgeW2v5EQq2mkuW
eww/AmaOlQQJ9Ldirc11vUqvQvY50D5N7Fqte8SqTxVoxZshAVYHQW6xpfiB19z1
AXW6ich3YGyPDJUmGaaqmR6JPwBArNi7H7/kuU0iYGcUPzLSUZ1K9TBDIZoZgzhl
OISoV+Wy1UNOpLWyr13qbDjx6Rby9FroAt2RQMOMi2G/30QV322AJY0+ptgeDdzV
lN4drlzYcrH1EokSLVFXI050/UnT3YPrKza668QwNw8i4u2jnbcDKr+7t69AjzI1
FU3DIMp5b7XZRXO5r6vCilhgsJnTJ98WoOsxWvD+0+IxCbmBnjFc5TFRP7qCse0r
84HjyyO+Q5sfI18mikRkzEj7sSsI9mJqA22U8ZJ5T+6M/Vycou4Ca8OMR9ji/3ZH
aH5uedG+Jo3i8AvdsEaGfGNrVNPtr28rp+4VA1U3kR67VGA4BztCQl+QkUykcAv+
zYzX7r205rZ/eHZgO9qq081qNEKgFVjFaX5pD/1dfJnBpwNBPePQcLYCSFEfQfp8
v2+6+AMqoJQQ7uS1vYQ99ievs3uEHDhmr7emwzgBL//cZPX976HSgBpOwW3L/B07
K40xeD+OlE7lsmw5NyyoAPbjH3qdT09v36WgxVNO6z+Un9BDNRGU0+plXUkWHs1w
ccqsQc1UzkGscOB88uWG1V6ZCsaKL0OJ12YUmsopkrFpg+cMzoqs39SRdJN8I2pP
Kl5Qmiu09lko+pcOyDr1n2M2bhGpMhl4GeDs2yRyJUmPeAxJg2ygiTN58AumTU3d
dq+yIAododnc4G9wEDozvF5mmYIi5fviHMm2EBLNx9CAzZCowcn3xayocfe0yGZa
m4SnkNeh/FAAG2US480RIOR+07gx12/2baOt3DlLLUAjEa78IyH7ER4EKSF/BwJz
nk+3s02bDf76OPexA0MQ3RQ0FMlSNh07uh7Pk8ygjeIBY/nC1akwnGnZvA4OGjBh
FOWzhcviXFr3gdF/jgld6TIRRfpWHb5OH/AZ/k87y9Q/35pUg3VeSrggJAjOqJ0e
7/GCb+dcnnd+Eqn7Rv4dRAv10DxKhpv/IPjBTct6vC7WdstHsvezXfl36Tb0/wL3
/cVj4Q+dXrrEN71nOiDEiR+uXnoQPG6LA8+tV+3D5qbOpGqQTfeEAZLgJ1sU5aAH
TrJdiFp+1J4BiXqQFpFOBdgh3TMmLVQSsExKzsXQoha6wdz9sciW8WWlS5faJlgN
PiMMkPxB3byaf/9XbXHV2rAWZ1NMTfGzD6Y8+6sNqSxwJhaRIkpCCizkt03ky/hs
/XsDvFeoCGo+BLqWy/gPU+D4keu8EYDCKUvC2ekQSlgEskBs6TGHIEQz2wfGWJBr
Tk9aySAtIgpX5no1n7Eo1ZrCpHjD+4hVMhgA3cStSI9GUSu0mhEPDC3o7h9Fbf2q
GGukTs0tIKWSxTaP3GJqWHAB33IdWK8gxhgJOdNzRN+2rkfZPBt2wyNTRJoZNzcs
jsZMxl61Co/sD/F5b97atnJDiuGl2zo8Yy71wRDxSpN5OAXWjLCM6tAPYPJJFmUH
NkUvDh4zQPpuAea4wv2dF2w9w/+EszGbEkE9Gt6pdBtwcjF0s1foqR1miGFn0peq
rvdH/VGSL+GjE+uLqtcBKNFgDWw9KRcoqq4mP4bK40aOtYOg/TtjRAZz43UvWSJC
7rnuDtrIBCswq/TGaGlBymRneTGLW1UPmkTinnWd+uKDQhHS6RYx65Nzgyr7gSLa
u18O8vPGoXqqXw+D4NPZ1oTUHMATlZRVdqlHuYiunuwOm9V6SFWJr8v+IqwPdXGh
hFTG+kLm5LCo88C6AVdvDOlSu1Z/95IYacuwACfwa/zGmJInSx8tYbO1NZ+IIJ/k
OYJFIPJZURYUeFszWP/WzLtXc575RMl+zWhTCKTMa2UTQNbUWjb94tuDfRJjlyiZ
N977vwO1zHTSCDeJueukXblU5XErFFYL7AsV/I+j5Zd2UnGopwdWUfy4KoBOiI9b
bBSh8cHVkaI4vMbCUDdb6RduD+qdQhjAVzu3Qd1n5Zs6Hs2xmye5Q/yVTSUv0R31
f8afVZrs4pNKRWfBUo5sCdtw1Nfq3iDiXHRNunayeTCnyaqf5KaQFN/2PqYqYYmF
0wT71RCbIQaYPGi6U+I/Ip5pce+YLFeiGwUW5ogwMyjbKp16XXy2ASmNWoq9DpbM
ImnOHYuUAPFoGLBxJSu7479mqXvE+zmLGpgn1LNtVdJG1f8dwkTLF/TsSJn6SjLb
UsCmHf3G1djWWPSwtQTom4OqpgKjen84iV9WrbQ/OJd98O/rRjH/nGNWStRR7ptC
c62LSvyedjZD+57J8OTtK934PQc/aLBkAydMnthnb63kcemPKpfzAqiV3S8gYxX2
0jOJgueuHVxOuVxvZUgqHcUUUpmsx2J9IGJQI3CbhKbzCtyzWc9RUhKqBoMYC+MR
sp7B5PgTxnF3GBkOCW1O1ia5cBH9WReT8UKD/l8S0iIuNPefGH1xLCBzboVpnLEr
p4RAglHMN6MZzyrxyvW11lXsNuf4AQCZKuYIsqpke6U2PfkRrvlon7buqlNiAP65
TIBDKaXJo2YGA+mfHpQn4Yv0RQVE4fZd8fJHE6UMl2EpCnlK8pP+VtfxSLwp6dql
UxJTI7XqjPiwFJgPH8aZVGARNem6A5vi3F63vRP4NEBjXve0yKetKK9cZII+pcVZ
3NsfgJL7svvPIkqlePwdXDh4HG+xsFAn8W2YYE/0KBgOGevQ7euHXUNIbMNVZPc2
6P4ceXVTtjqyb431dAZc+FI0YHDxMc5RG52WocFJomjmyx2jtw5x2JasZ44DqqC8
49ofLj10Hnq5ODl80MLW5MeD2MmC9ShskcAj37qfHVuwPPD7wyIPLFgc10kgls7j
Qi+rXL+wS6n10cwUS3CN8HstnOAXfJt+4P0w2n1nUgkAc3ulVxuLOb1M2s9/RFFf
fdHT1nsyiv/P8JZPfnDF4fR8TuSxC552OuHcP0aPNS2uFMCUZGQyNIhd/V0yp8Y8
gTEStbXe9MqUAPMR3FZuw48B3w53mF7jAQ+D+Hlt1H6o1L3+kOMtZJSuwgGEfVZC
WZZyaQ1tKyQvMzUNyrbBpUPrsOq0uj+Ddb7U8aRVT7R8MQSlVNRGk7N19NPMNgr0
r1dINFtY9gQZbSQNfx+7rcd0o5p5QdvYIMVv0GhDjLFP1wKVh9wMebo5at/lF8b3
89g1erRrCJRujl+Aqq6ei/j6cT6GU3ofo+VA861/M0Q9gkhoZ/dbgJBc3dMzIrIF
3Dxw/ZXtiMiTmRWKgXUUjgsiFUQOcaqJmzPYxQ62n8ksS4UiMNAQDuaBUqQOYVtg
kf3Hk37oFyCI9NhbJwZo5qr2mI9R002nQ787ugwMPAWy17vQzX1Dv+EMyReU1uyb
+oHv3n3hCt69q2N8crFzUG3yxSbwM+3ov0PKEoxqB01+FgbdrVKs3W8T7hQKmFwL
i/+JPh+NXqfxMXUTPKaYluplU/9W8OsEuAmH+mvxq3KABDr8+0FM95HtKSaB4zUn
IfO6OoPNgG3ryBNAyw8k6zQnIcRHSfCiJQLaHyltgkt5QA1+urgmnrVQn6Ih6myi
FmillocYoJErDM9vMbFFwAQcfktQWwkPePbqZLHLczucw/RbYEJsbsuHxdyzcD4l
cCs6Lo6SaJPaPhjzVPcSKWEmOuwV007wmPNeB2P3PzKCpB/Fm5Muqa6ITJIk/wzW
+MsPLyzyWP+8LfNgUdVcfzvJ3N/lXHWNir2IwOPXLsZ1tnWUq++C4DCObD7ka2OD
5AXAXRmkWW1dDznqisoyapXcVf+4APCaFplug83RQijH7MjdfEIBOnj4AIQNxq91
TVaLDozjKOjDZFKPUMuTl1ZF4MJwSNUbOOrD9bKIyIF2XquIQLynL1zidAPmDPFx
6Fdvx5x+NkWxJKlBHj5IsVpAk1qTD68I7NycToP4Su3ZuYUgGk/DqMITnCDe7uGg
JxxjJ8LFKR2lqGkod0JYLU+rKOuXgHgWzc0kfcGq1vH3QE3L8bouFfqyxSpUwxD0
mh3qinoKfRGVxBzMgb+Lt3mScTeoYFqXFB/eFuX0FhBVJ56DNUlgixGWhB1bTkVj
HfEsigtAATHDsCVkGhhyoZbXSu1aYBmYYTnLSWVSxmMuD6KCD4QGMQvybn0x20Cp
ipMnyWEHXEiMDms61iITA3h8yr0Ima3BZ8SrTFXfDN+ZkaC0CRhgSBa6gQueBtj7
e1X/sF2f4OaCdSeCnPwXrIcY4x9+syXTLjbF5yTAIFAQYzwxRau39fz1DrKJNzid
nW8jgJC9fqZGu9KhLrq2LmJ9c++AZwDs407as1znnwscZ3KUrJXXIE1cPNl/9PZS
OLUAs8IvdQOVrkQR+sY02To6Vk7u3QQfMJVT/E8MsQ2n8TArl2Skclq14Po17K1B
XjoAYzHRHwoAwAxDNoYRWg+80MKegu8VGDoOj0PjgDQ/eYHKlMPJObTSnjxl2ABr
8ERF6CCaYf0wCK9FedkOFQTp2D7XNFCNs3bY5Io/8As/Tsi9XAUdXkqivIPT7DgC
YyWiJOtuNAGNAjA5PaRSMtgyll34GkbjjW/T7NFiN0HXB9hXFah32qQQPmYOxN3P
xdsSJbiO1Dk8ICySMlgxkF3uAmvWddHhSVc9m32fLGY8j2bGrdyOrSmMM4Te6olh
TvrF56/8Fl8oAspEwdbrSyBCqe9F4dPc6nWsCaQKgKPUz0CTBC/G9f4MKFsRp/oi
eTg1NNIr8j8NTwf/8ijsF2kVtJK+TnA1t++MZhNUi2HUiOGg8j0PKhws+1iLSCF/
7dziTVnJ0T42hUE1z5secSWVJAsVY2X5M68mTwAz8rUCha4V/X8ZL+/gzaOIWunD
veskRm2rLiYocXjCIS/E1TYdrRpIoBypJDrQuN1/x4EJyyyBAFqe9hQ+9mhiBQ3f
MHPJhpHg+tYSNv8VxVNcoBjX9+8FhRQzJa4Q9xM0KUDO9o8Alax5NKjg7HwG98yo
6CEIzaOwQS0awE5WWzZOm1rYQZ/IcNdZR6pJII+OK1QTQsbltfj6AKQ/ofomrmgL
+NeX7R/7OnG6ugDJduN0pyzg5MbON8IhfwCUx0ZTZC+J4t+CWjaTbvbCNfIkW9qN
M5MZvlAu01PYYIP9kZaCzccvk7ImwcWhxho1ScO32rRtcPotNnzSLnlUlj3Sq+p6
EBppHM3vT+7q3OmuSWnvn2L0pNkLKivh3q2H5DEh9bme8valnN5CI10KyJUP0FKw
I9wxCDsaWEtlvld3S2wSbOKk2zfbun46YSncGl0+ae1VZH5GZ/jNbAIEiFIuu6UB
11kVDDzKu+DwMCO/SjrBUKgeRi1pConhx/TISEGBr6yhVbNOen/SDhplMeP8huiP
GNpczcYfGA4civTcLDPz3sjppZXE+XPsnpFb+fbWSXJbOCunTs47qDihaEoou92o
lDSIG2x18BAP1Gcs7mv+2Tr0tYCHDM8A4WcXSsitM8BxIwJn1r/GPbYe+j0Prp9I
ZUvEYChsH0N4xuNedaBPSm6RvmICEmeuNgIvI1NRG8Su6oh8FfJ86tIg4Mqi5nFE
u5gbpLOuN+YOnV7z7FU5lb7MSjEMJ5iaJwvlZV0bqFcbK/iZM0v2w0nPP7THKuEt
RMAJhSAXR2xhO70n6z/9rvYAPKYAgjcMQtj7/wAnAl5y0iaY7Ok32WWkKfUQtfeW
goKlFx5I24oldkezEJgFhN+H7maie6S1NBkOwoSc6VqFJAnLKkWudzbgoMcKHksc
DZqBykNKm6FapZplj6mmeEnTzkuo102IQwZ+8beN9YUPDtmIqKDxevHEfyKTwDTZ
qRNNIRyTEJF8tVYaViAIesMDcpiq6BTFYV9mAIDaqkXs6IEm+PwDiVB3TTFTWDWs
dKn+q/1X+Gr8zVTcgVEdLTfrQnewCiy2IAPjv9/rrpXo7slL7r7r+gGgFCLzvj3n
Co7AEDfi7aQvNXikGU0yey17Pc9MXn+b0lwd5tYrkUUkEtGAw3gvfDCuYoAjhZrI
wdJ0Uc4u5zdkD60TL+ektFR8r5eU++4n63C3IVc0xTDtfWrbiL87UrjlXfEe0tE1
UloZbVEU3h6ujSrgMupugybDOb68pvhYTMWaGhD3RM1dUsKfB6NP5X+wNSwrtTph
SdabEMkrnUhkT3YbcbqwriDzkGEuOdfnEMfqvc/IJAtvCOAjmk4qQEe95y0jobKw
sERlhgeT6TYCCXzrugEzuOXt9A61CYVngpAV/4cjP4YRBCSFO2LCaM6PIq1r5iPk
K2jlvC1xPWzP9FCthlJmexowoeMy8wSCYJ9r2lpaNwpRy97QggIbGIIPhV+uLFZQ
jf2omlfm8MMacI/v2J3znxGXm3WT6Rx4MNmtOw4K0hBKoH6lLAkggJJnAu5NdDFN
SHxfNMsTTkSjo5naEaVwhXiqDH0Fp4v/ZbErjpBD/xOBdmRsikNKNlm/Zx5vFtL7
eyOU6auKxKr1MjXssby4sAu6sTw6lJTd02OJlwngOMuj3l9G7w+uOBd3r2CGDo37
UzBDx/mDhlK+uIscYYgbqXoTTkncIkYhR0aQw3UuLoAsyuU5KKa9rrwGAZUugXxm
S1NNSyHwTyG0tvybyjDuVnSm15cIV+V03LjHGQABvuT7MtoFc6WqInW9GBWxHSGn
Lr31vfuaSDWlyzUFhW6Glr/0gpkbM+mhHfIp852oLOhfYgXgEyD67PKcPsvMxgAE
8H8w0ycNSsi1AfppgvyK4DQeOfXQR8T3g9pcMTka0TbRRU+SptAHae38l/DSZeLP
Uhgny7WPMKCNRK37KX2LB7gIov1CekWLL/iP4cT38iUh6yVabAmh6jBChyMc212c
6Iw8cdPqycmvtbv5FbdvQ04o0OB+0iT8PtsFcq6qK+L/Ud8xeQnnibtVmNysUSuI
YiaYDYkpefy7huLFk3fwVQapKSBeNeZuSoSXIlEK1dOEOZEDrOyBzKIfDad/nJoI
u6pY5TmIs6IG2IKBTFN+YjgTYP/HjAx5YwTtEoo8tUShsrtI9pBk3raOWbg01c61
/itmsmPSiH8jWvrWxl9rgWoxRtTtcKeqN8/53x7uFg0uc0Hz4QQwYjrCcsf5P/pc
7K0X8y07BmF2zCIodZ+/Ll2zSPYkUKKo2twForAOSG3eHF6SSnEibvjrdANXUIS2
qzwU6mfUyh/y9/6slZ4nPHhcFhIkGJ3DwF2inJawNxWq+EkHY8swyV+gVQnQiGLn
0RcUFAtWESvLWFyCnEAuIg+0eWthgJCvJf/Z7p9hBh7NduJM8nEI7DZ3lQXzKOEL
k/fM7HauokpM8ksQWlaQDvjbPfEkkHgQoU3CXHgzgHXs7xEugdV+SS5Igxj+OAeo
1uXJdqSUnvWkPVLn36s9t/ngwF/ag89l/Ilz6g2xOkQobWADBLkeAnF47tCgzPb0
kckR2kyQk6Q8t34UDECE4RUHSsebpbnkRtAUErDMOgEviBQM5jw0FEAo4SOyLn56
AtNaT1I+zv90h+yDb2z3iPrMWxrp7HpMPrHNtoMqL7d0lQdLrowXXMPX5iBsmW6C
klzsvKnwBgKxVAvxfarsM81Vrl2iwWlu0P1Dhn5xd7UyTHsjghc0kbz8KOEYF7PW
d4d3I1kby8I9CgJoIfcOSh/LKKaGXtnesbFNbIlIGZSpI7YWYP+FxwHdzzUFn/1y
Nn8rw+HNAMbfSzO0E9XLtieOe7kcJElSoQ5X7jv9SexRc9VRwybaToFZT1ovUnAh
bW0gk8WfkQj4gku95aF89gThZDQL/BxKtthfY+kxYEKXYAvxrKI8/4DZjjyclP1n
FhQd7yzRKFUwInJxKOGZYVrq5gDEwqHhyiQZwIV7CK5T/LYlwmArB9vz+hgfNBDw
rho0tyIaGDEFeVaSXamonJhSOy545lXk1Ch2dVk/hnLDSHrLG1+FP5nPQWZiYBhE
oUNcyW51yrSK4GrcvAbOOGYCB5I8AUYe+W1hQH7pVlCAx7hQfDCyKglvAOC7jpOA
yWvwbReBlcJT8UDjfzMLbnu5uFbIbNCZVSgC9I2dTE7tEKcnkZ/vTM6dPfVjzNbZ
eREHiEVRy2lC7PD/yy/XD4TBHaA/jhDFruQp83S2vw8K7n8oEqGAPIn1xS0MiU64
ofu633STwoB3EdhP2ysNLhmNcNYSeYR3t9Eg+x4WI0QKv1ioevdEiRhZfOJSPLXR
zIp+CpZoLP2UDT8JIj+IifP96Bc2Bt10U7iuMw4qYcCATLdVN8haEjZ2KD76xHsv
9ol/rLLrhqZv7K7t9fKwgb35M/BSdNhQpYZbF0a1mJNBt8oMBfbHhOuCiaxpss0s
iaFCthjehiaw2gFwfa9IWVgFm1BsLt+OTjVpBUlwivM14+9aO7HBDomF4FVf0CNs
mFk9Kl/Xs95k5Hs99O3tqdT2TkADA61CRmMLVhRhXPe7IGkQZHad4uhPSkKMWVua
XSkGVctgOyWLjZ09o7utB/NoMdMzsBSV+gECTb1ePWgdfc3x8exs+JL/z+Wk8PUR
6w18m9dpGhlOkMY8eYdb/l9/QutxBshVu1RaSqM8nFwWHl1NPMK6hcVTcM89dSFV
s5q1J/fBFs0b51fRMUDpErCcb7kruYcpuBBkogE5spThktYrA9O7ZrG0nwFtXg//
L0v9B0/iEMOOzPPSPJWGtHulZVCYkwMPcHaAjCEXs2qvZ9xgwMvnU6qMAI2QovtC
lQZabrYssaLdCB5zqmEBfVwRzt6hvVWmQLtjfFwD0Cao2X+fRunnX/GEq84daiXG
cloYJOPc/5ZydIrdt+7ZvnvbwGHqydHR5h2WQAggnYgyKIy46KXwHOnUTOEZCB3C
u3i2IsUx8q+lJ4vAKXDicgfgkNcM0YGGRH+WFkx7rAy/eVJ9DxGsZvETjhBOdssU
GBIKd/Oc0zEKWu0gmIKVXUqUTqHpqlGqTNit2tVE9lREtb7uNOZ6URTXhEzhJzfd
CQIRoZLsAT53Cz7EyA0/dkaEbeX6WNq8Sm5PczUsf/qIBIx3S2LdnbmIXufPfzZw
0o0hgGrG6U0f0DyQVzHe7QTrs6nn1zk6bgm+C4TTcQdrU1fiqOr0AvqwC7Tt3zCl
1j461kBDNn5dy6o69cJNuoqomK+7VZVSqFCjg2w4VnZwpAQJomJDqJ2z0aUGDv6g
uA9diR1u8pPnJ3DFQxXS5QMy7dO91OPYsvjcP1Z2k8vUSQOdxPP+JO2SnaUjJw0R
2MjW50QmDMQplRhtSAlClTTwPJmm7pV8xAAAxuk10QRYdQvGDt3jmjSvJ7blpnwV
4KsLNusAp/wAFqvOuHYfe+jq8poZ52CUwdgEslqYsAm6RFj3RdpvYlQ6Afc/0ubt
it3CJsiwpwtKNyUSgmsY8bUoeowXohsswhY0JcXx7WY0CuN5c1fgnlwJBnOsRM0m
5NDOgmLbr9mYuqFKRh2xnrACPGRL/JSxaGW906jj0JPcMvB6slRnoX1gLBCahEdU
CaF5mZX0u9FUvKSMAXA3Jvm7bJQSbxYLVCZtugMgRoDASEggCpqeZ3l19LSAbxHq
0OxPoQ6imhGXSGdR6HT9qUfcN6FItVKfZK7I7Wyn1iSTjuqAZaa291OyY6OQozR/
2WMPpW1hOiLVfj4fwpuGTh88iu5PI/J12I4ScbH3wf+Ftzoi+OFNAo4PG0Npcbnj
xcuUha2NCIIUN0+7QDc9G2O+E5ijPZXOuYmJjAms7GM0Xx0sFautcWFBF8BBTZHD
k2aWMIrBhF8ppIla89lw8HJCsYEA8k/5ucjtPC6LvmGSnSBzW3PD4XCOEJz+Mx80
wHNpi1eSXaSLa2ZuxyIcQVSVKmpR4sjwKrXnmYfDTJiREqukU9UIFYpjgq+O0Wlz
pLLQfixLlcsvnXG7Oodvyur/SV8NslwlXQKfh4CV5wUGjjUtQnsTdwadYsBcmPcc
0LJokio5upvEfnp7XTmrOkSLRolzQu3pan0m0eA61YaCckUgf70o0TXdkbu7TETL
4twHbjhaQ2XEbvmLPEj66dJzTNgrMn22JHUkJ2r4pWqtw/BxPXc/LqVGnctoZfVG
6+yF3M7p8JIvXo5ZBMe5GfKsLUihuKqbinyl+Y2Z1SSuU3zJzJlzybKKsP7+Jaoj
w6gsRrjBAikksF/UQnndbAd/ndrhugEp6+u9yroTqo8sSB23YDj0RdKCFyyCIFmh
e4mhnwBoKi3aZmHUQHLDW4MsHU7FsD0s5SShXLjNZv61T+z3mkEwTgAxljOeqSaQ
o8SxeMY+PRm/2fjXPQg4pHVdLPdbm6BNTzV7kxqN6jkfCAiSFKwIqp0Ec/QH5wOz
AW8vU62RqbUvc9whIDy/jc56Czy4G6YXJ0mW3SwDiE4E1Sxdk1b8pgk2LIFqMTWe
WEkIB4uWlrHtOjxTUvyDeyWHgRYpy/4lsqn7yk60C1RVhs2zp5iLaOjkZdBglncM
Oub4tb+uzvAVGlHds+4qEWb0a7K//3zr5hiVBe+YeIfXDLLmagZboCpxlFLkKmTY
zmalMBBQCj4DZrmVdD/34XmhAYGiXZr+E3PoPddHU7sHtY6cpEXrQsRA2Do1L+nh
e5+QByfpg5F1IDjshFKHrs+ReT02QJB9e9fSURYuRi91GawJ+UUrZUMp1kjTpthY
S/+y/VVKRTdJ+/8zWGmn/cFZghrxRqCOOuTsl8E80W1AxuMPpjm8w3FikGBtfjn5
l+d3jDvWLW6kwSuLl44/RThGQud2illlCcp+M3RPVCL1U2fVGSwQZ1B75+tCN9BZ
WK4WjPzoD8w2QSoCeFJjNlg9ZPMyz8gN//MmVyL1cNqUjvUTplCVM9mqJM4hPO0H
5h4cKHgqfG24OaGuCBKc8LWe2ivcZyGX7x6qHL3i/A3wF+NpSDLBILbf4sbXNimq
tGa/nOiGwxGjdSB4t9OXC5VCXS0lU2lW4ia9kLXDERp0hDlZIp2gwQSKGkPA2GG8
G8tYh84pkfmkUUHoFzWOqs8ZPjx4nQjVgCj74nHaz7q5UB8ZVIJrAPIwvkopgILU
6ZgKHo4JyqoniBHpumz92kkft7UCKFkmsQgichWa1VevXCCrFbm5+n6hPyhniO46
NBtTQf9jJD8Yf7tpBqL51zVuFRgtSmKDqsLGEcAhhfQohIA8gDsBEpy2wR+dDvjv
SK+pl8iCayucIIujlInGDwK6XveRuonImW0hBVRYxdQpBmzi+H2jbxvhwfHAHvEi
UXT7n4DLPRJZff8N1FGWLJ8N2yuY5w4QpCBqyE0Pwbj/yLVWPuf7tDAyPx7l0lox
W/txenMk06t13QY8nU+oiosJdha1PvgPJlfwpwf1lHz4H4BLqanSSpvyglWIMWif
EDH6YdAvlwVqt4F5ndYcCMEhV828qMK0lclSZF+Ox2fePoj9gBBxaBh7KFHAnzks
fWi3KvfzHpuBB8Szp57uA/HOezQp1nJT+xj7TqRXbVPqDO8SfeSFeI3a/QRJcARo
btMu03FnUg/QLviaFXTOxbBYtbKwRGpmk3Yp81ITZPhZC8ulTKT43EoAxarrFhu0
9f5Xz7vVVjXkdk27fzqjIp3mIquSlGARZxAjHaeopc0v9kiUITFSIa/ebz99uTpf
G5uiM1Qb6naNVkE2BBMIsYPQv5+IoL6npYgaggsKArJZofV+C+MA+VxZu6nYzhjg
K3jCvStThGcb4me01wAwZqbpDBrBI3UroY7JgoCoqzghvs9l/W45rZMytlLPPPe5
MpjZzptVPqycX6ZQSL4EMK/hZGquYrz3ZDGoWyuHSooBobuG1M8/A448GoagUe17
6xcnsV4JA30DpXtaJHGAybtb8iZc+bqBEy0fP3X+5dGG1QVsh08bw+YNp+WaZZ8F
t1eyUpYCDP6dUpU02oI8shO7PNXQpIC9QOaB7FunS9WGJcuHuBNpR50Aqx3hOaNe
75X9BkqFQ2f2+fhJUaCZykR31v4lMwz9Tj+qaM1FwhsER5srE4C8KlKL/NPHfo0N
Hlc+mB/kIjsyWxV6j6o5LI3CGBeIpRQLIX5dbNDbQ5Uhazp4WkGINUkieSeCWO/F
jk52WAC7Yro95p+NDIMY0btwhA3LP4Qfr8RoKyY85a+iWCfLIuvAzsMB7yiWM0bN
CyCx+67ui3obBqdWimf3zFfPIMAphaVlw4rN1x7+ALI2T0kvu6xHi5WnNO3nLUp2
RuFEhV3uc1h1fFSumo7ZwJ2u3LsjZ0eVWeOKFrneoe9o28H8BKaGPNC/v66+6BSK
fM2M9jssuMQ6ekrw3JajGCFeI4oSoq/mhX/RCsz00i6LQk6dVIe9ChQUq90T/1Y/
8l6howvN6S3NPHos7fooUJS8NrV2nBLOmhrnmceQgXQvJSCha2CfgfbsQqt1308X
l98UUzPyU698LpuWNGgYXdFOGSHgGD+lph06FckODAlXBIKZ6C4NZ9CeXikr6y3v
fAy3Cu8w8KvV4C2tkRKFdulo75WvwRXbUra8wRLu5ZM1GfQh+oYKGXZb879x6WrI
epZGas+mO17jfrnXRzDICHfQ4Sh9jr+DW1wFUB46HhM7zCYTXkw6MDl8W8KElDyI
KsqOp6lof6d1AFQckURnjCe79U0r3+gaH5U15g/9Uc3cy3oQDUrxUxHjNakiC8UZ
y2lZiWMoupvQLOAdw3RY4qrnubHAf/iksr6WExZwIQeF7KHFhkcbIu7fRtYc1M+Q
L5h/x5gNAN5/wxb0pXfJbDeMI7rNT/Z2SZi8BLg0jIykDp2aVK7N5G1D+giggQ51
M6dyuBTrlo0vOmsHHrmgILM6x3xUmeeIau41CTnMr8t6oPPGvbIInRE5qdIOGSsr
GFZbW/fgbfB38T19gsg/2w3KgxWbK+NVhSsTQz6wXSKRpuxF8uU6omysqtYZ+RlN
b5yFp2gbokvu2/8VNG0ifT/wdZosb+r9xvlHgdilVZBTLDBSnEUrEgdDdOtLhWDu
cNnTxMqiG2H/gjALl2Ipb7qLljwx/7Ra1xFalsLLhfa2zVqmbkxTaBHZAQvMPZ/L
+Q/m+O8vgx8Wr77YWTpzo7+I1/UI0iv37v24pvZS+wJErgzNb0sxyow7HS2QzXWL
/LpeEbX1pl387vTn31t3a2vOSEo8MZZXbJf3RRH4Cz5UWB9fLTc9VEw4leEoMwlK
cU1jB9pzDVIhXHSH8TGhXqhMbbDPxuW2q4gWWNaRpF65gOs8kyoSQr9umzUcER5H
CEPpqWMrqPtbE55l1za7gAD4hfJTmRJqBd10ypmblY4TYfH0Mq1qNF3LBCEM7Ziy
ovneHUeuULEM6Qbgw8P1E5O+L3RFIU1kr2jZHRLaLasSkZyP+SRR7Fa1T6SulFlG
h3eUbX0FFEwAaN/Ordp9xxC1donnB2bdb8WdXXjVstCa8bF7/t/nUXBv1n+dNxb4
rpnkSrWYAzBUOsaTjC/iN9rjkmhu+8ZWIzv+vZe9gHJ5RV0KSVRwwJro/O0fkcTA
vGYEwif0Cb03YxVJDiIMHz8t6miwalPJWaMe8y0+eYpcTajs7+NedljnKEryhRRv
RKlTHhpxgBoeXn0Gidhtbc0gHft/O/QQqCmxSUhTIjur+D2iVbcV1uq0TQSy3fmx
C1DhoPITPiQLdHnaOKVAjiTd/mSP9xKgsdeF2gOioYa2vE/bwAV8AKBgvnzDQsXO
fQVL6eAZUmWZUQT4z7GeGoDAiPcstJeDEWxtQLCBXRncyHCx/zFyAkP1XutwZHs2
u6/AzmdgrCdHBt2pKCrj1urPx2JrAa1sx1QUtBdwdjmv21NfDMr/7LeFQpmBDrEy
5xq44KQ0swszgQ6SoAhKJ03h53cgUiUFYKKUhe/WqmnA2TAcpAASD7WKlbvewxd3
SNLQTvpWuSLmw/pnZDIeKg0hD+O67m2likaQaud2GrNGVfsge+lLGrEbKqZYNQy5
/kAGzAl9PEp5GGJ4ZmyFYpPNepZOUwgVJoDUHzXtsEp6+cZVOOyiP/tZDpCx9T5e
crETkctgCtDNCa2ApArUa1EUQ7zQWYZETez8g/AjrNnd+GAQmYuf1+g7VEUZe1F4
qfmGiNPNSlZKd8VRQlh0nCWd4MICOYEkX1KjOqH2o9iTwdkHv8gHS2ynohZZ0DXB
7eChmqrIzaSC0XZoqtq8CeTVqB34BRfSWt2GsWWn1fJKJeJAq27liGx3BDLE7WZK
Xqu1AuoukssEgQ+sUh7HIHTKiL/J8v6MaI3Ay1/jbOBKm/tst/G9e43bTc06kPOX
8gfNVAuk1jgR+rEGuXzJXzNpoT/Rubft7c5ayvOZv0lpnxWyBRGeEu98IKfZeOX6
Ih3kZnv5CPw129049XmpEeY4L1MNNnopwQJ4JH4A8Hxu7ADgxZshf3VFV0SBAZpw
dc1F1qkE3mbBirDzQ+d/sBenqZ3jnXgj9tgr/7aotRFW5rRyk20vU4wL4iDnw+01
eIEe+E2QUdJBHYIFWEyXpR/grGHGRPXh8NBheioZEXEuUi3uTcX446AHFNBdZvWz
ead8zMv2/SI9YAbrJMXyAePp3S5uL2exHs826LtXIcCFlxNUV44cEr7RirH21Qhb
tDIln6mP1qxSwgwP5aujsb6CGNH2OaE5YXlGGWkyLIujgMNmeqsM5edF8hb3Bf1E
442BNPQS9RE7Dcj/bUTMLLXItAYmF1OHZRQmkcBo0KoNgBACXCLSsjV2xRghFQ4j
B/4mqC9Tp6HzdefzL0rW3sTFdZfWK+lcejVhi9I/hQXMPtgjIcucTEAPHlC78mLQ
rEX3t762uu9ZQa1zS3JbiShDZ4J/hgk3LXvTJOwm6DalcTCNDAbnhfb9y3ScMWtD
aPFovXxCyXP9TUe1V/d2PXyY4/wDV7mE7a673uL697R6U9yXw+BdKNySrtJZ7hUK
v8LlcZVl4hjACHHkGEhLBbVtNMj38Uv3PBhWlh1nQoEQ5cvJAxMA682OMyjOEp2s
rzY2H+kmO5zW3sc0ALHpQO4kNCndQFdTJ2bSo6EbesCtFSWrI1yiLf4vDK97n7uG
r3qm/3HbdC4bz7FmZ8wsfuiVMpeqNCP65P0wy6K8l8usczbz4xyuokzlDxGYzUqA
NCYwoDkI/zEr4x9X4zGXW7QIq8W0/s79DLCJovnjHZNvntw9EiMYwjV56z+nf3Rl
vwI+UcLud3gRUk6Yq0rR+4HaYy7SetYwWSXqIJej7Ah/KHP9UcKh/+DPse2SpQIK
GHYsNnJ+GcByfgcQfQINNLtsFpj4m4gZVaiq/mxyiNd/bxn3nQpirYNeacDhZjn0
gZBDE5YhBYNdWM5OiwdCkMKF9ArtJbNtZk9U0JVf9m3kDl4FxsCbW7WBYwjKkWl5
YkJpdXqcDwmej6A+Y5pJ2mtOM9AIU/UiC+tsWV9d5uFRogL/TI1gO4GtJeOZVesy
EzG8hf/aTvuZTKTiL/BKVL5xveW6oIWBh6213BMwf1hScwVDnbyrZtaaB2spN9oM
5kLhYLQjZwc0LEYuGY8GW/olebhvquMVRn9wx7clXeZNR4Zjb2SXuvn7HpXzGQ/j
koygNf9cUhlzpyfZMMj3HDrISj4Xp4ofmZJAaoUr9KOdn6A+CHaRCtQZw5w6vTGY
YrbZILVY85rP8overtZJSrMqV9QyifqY1+H5sa86ogCFmm43nfbZ2VotfGHoLgZ0
P7vbrjXYw4xZAFmzdbduCr51MX+yB97qe8ddtelcacGsaU2Ahhzc7jp0ogyoiI2G
mtjDyCcV8EGC0UFy6jMGxgiqDQ8cBGlX7SKakgWbVRvBai2WYY70tLEu+lzwseSu
wEY6g1XM1J5/Z6LONenfpRyLznKJrhPDMrobf2pO3gGKBbXSnnAI2Bv5Xa1ZOEuN
/QZLZ67w1CmiiYeo1q8rRGQVhzMe6ZyLyyyJc4yz8VTW5HgVEZtitbnaLpFzfhxh
inX3gHuQRrHsivfLqad3EAF5kY6gxsjCFKA7v/kJToZ8f5BvvK9z93l7lGBTQfPz
aELUnOc3st0j6vzlkRFvnJrNhgk5iAj6PAU85glLsq2/7aIOZQkp2aS1WK7JVvvX
hTyX8p1fmI7q4a8tjVjPrYcPLOXObY0x9PdowZPvUceAb3z/eQK8uzS2jEGTaq//
0QjuhqDr4FyuPtaxv8VplJbUBN31vcSFU9eUU/7GaB6gaMOku6ay8Ri9WuJl3bQN
6cj+3KGybGUBKZyeJn5q0fadanp16NYT2va5WQLhLCrM88LzoIIAXjDhk+D5g90X
ny0fTs1r4n06/lEXO97yokctQgDHupTT6icYPgLViMuwXx14rvmTPfcKWow9tfS/
Cze3cCBjZp3EOwxMdmKc8MdjUOLdXs/uMmh4M1hDdmGHBspmvAOx9lxVxdrlNJy2
DzSmnPmWRTNOunzkWmos5EFquP+0ZgRPDUKya8WdFfBD+AC6zigbB12DFwC+bo6B
rDrcUB02GdjDjeBTHLZUFpMnTk00GQNIpaCky3oqsnZ+HYkKheKS7453A/f1Z6o0
o0jMMli0YHLT7k2C9zHO4if1kqUWz1hg1uXtsxlSlf+ADW0MmNW7umFSIFjd4I4C
HY4+/2alpv9vTWs5nVQg/fvEXLgRNOpla+q5uiLeY+NfpK/LfG/AhFsIcHiQiSYG
kVrdni2ydfO+0cxqiG3O6MpjoRpkr5wSu2RhAYlFSCnmtmJeV0GArm30YoEUn1uT
UlHG4hXIyi/Y+h1AKgctTHu9x/lGky7a7g7wHEr1sjmUbUH01MmRp9Rz4EUtStM2
aFO+KwkY9q5nehe6HkMcrTbiETTwlFRkMMh0RCeNPAfvQN+bLtu9RbOXEQUF8SM6
rRYk+0W7+bXwjaJM3EPWMWPz+xVmYaK5/y/42OCJWBERHb7G6oWgDTkvUgBa9eIh
FXA77dcIfFYmuk/MFyoOYSUlqP8sOKg54LRc1rpgxl8OgUETxYB3UI46QdTocdKw
XQWLIELGFFmDYsncxKG4NhvglQwEOOoL3qANB4E0ONn5SBQrBcAfVrkT+zS05WrF
NvK/DQ2Wn3KEIGOlHPz0z+kc+rp/+/tYXOH3h0Lm0xTYNSs0ShszgPlMLC7rYiY/
FjPJ3sKZG5OMh0wZFFfmUmhrMn6Mk8/vlo2EnzO4NViWvPAkYykGa1Q46fCuZP9q
ZOchukILFgO03i4g1O3l16MaW1nuH3YIwwyoov+VZ6HA5ccqvr85U0GE98IZniyJ
BQvwjjNxOCOhlsdrujF/1Ay42QQeixJ3OjwDZEq7SDxW1FRP9DY4hWXUa8Ueziqt
QfYEYojBjWJ8W2UwCCVHzH5S3yMhrFWJyGpjL8ImAbn2DMulYy66Il2VRZomeKkq
vMxcnj4WIix32WRr56ZcMMbrZeG7r8v863ciaURCp8P+W/A0diTfKNQlP03dr7NV
bKb6KJJrWUGb2nPERW064FJfT4tDmzhJnjHunXLr8TLuxWF/mnf1rqx8CloCuux3
CQpEglwvkXdYnsY9dJnjOf901zzIbWwnSYNR6BE3iHmowvBlXHBjZJmxEQWWyRHj
Rh4pF03scEJay4wk+TzL+7mWZ9yVl8oE3IrNTwT5vdy4ApVLZ+wJRSt684ZgzGVx
LjcvgTKR+Xq60icBQHqUVL8V3ZKR04fivj7+51QdGSOr5HYOtm/mJxQ1NG1cZ/8J
4f1hbiM/R5M/XF1CREQAaZ4Bl3lMUrhrmprrEg9TzO2JxxgGZGNFINaKUTPYQFmB
ylXENe6iljoLOL1JZvP+c7SZSjOlKpsmS6dUuQYwpLxFr6u8GPvRdElZuhjbRoFy
eBYJgbCbKk6MaSyJ5BU5Z25ZidR/iGiPp0Fsdw053QEmVsIYGkOme+tdJ7NThW7Z
+ofb/2wL7TPbj7a6MrPBRmWGj834Sq3QlZrsrukItDUbG45TTbW3ZGb7GlU7fO3e
N+tNZkSYZO+SV29i57LO8jur2i9asSnGVZJApMD1MZekUq0NjPEuXViAK4ib3V+C
CiRtTdqCwg5k9FlNgox2H2U7iJMmWFqBqjRhNUY5CD9Q8Q+q0wx/1cC3i7MTJEda
rcpYwsBwrwaPKIYaEBFG9wd6D4t+6pWlF/s/STGqgDgZO5pfcHNOoLSvaMTmZXp8
zQlyL1AlEhFjziXhuuIdzi9tFaCkdgcGuEBjWDEmGV8PHSFKyh+TD8Dwpskex2Qz
B5hwQ4ROD066LzCb56fR79peB4xvKlSIlSxuOzT0v5ime5I/v/vBRYouGhyR9GdV
9nKzT0jFP6c/R7gIx7ulgWRsLXAG+2vflhowkht6ERy7ayYav6a04pz+tUTJGtGF
MIOVEo+mXNnG2BTR4ca+xSixpX7uqiEM0eYa4NRgKchAmBif6AiiKTgjNYupRi1s
uMM9x/Mk9cOrym9U2slE/ZL4dz6wVbUK2GN39XG0esb6LAytvwYaoPa+nNXk4lx7
2CfIW5hPqjlaZ4u7IGRJS1skCR5t6bqaS8fS+uc1aBfgSrOaeBD55mhQXYERxx1F
Fjha1ndzqkUfk52lJhlXtS5ThKnAdkE16Ubw4eGVbPpFgHur/zwWtt0vOaa2p7ro
eci28DwL6EvDMyR0mR1IskEMV8a7olVuic/nIDzworKhwpOveFo4THBGY+Id8VtR
OTg9QtQMVck5+3XhZyctLysShaA4dR23B3qvHmOJtkGwPmKooDcczxP5wgMZ1OP9
OjW6D0W0HutkBzA6bLhNBsRuontnzgvYY6xdT6G7s+JiO2IbIWRay+K2BgzO2XHZ
WByHxKd7QMhYzgqOGfsuQ1WLnFxsgmz9wX171S+D8bhmSPwxZs9Nbkye8YVZQtrr
P24nBGGn+mFa9Ni/XpCnKy8gqZufxEdYu9xcB6ZOD16D6ilKG2YQkWDZayzNoXbM
t3sUvK0UixeuPQHzWPzuyZfT77ctSWf3A5cItgb5lcQhYuo/2Np3XVzaz4dXF81u
b5ZuZPNQ0xQ4+1cx28Z+EIHnIaa7QKDQYSLe/tH/tEim8+YHhSvy1xI6c+0nIQYZ
LkKW7gXXzXeawMInF5ouUEMVuHde6kyG1DzsYlRygfM79+YS56b5q4SxP/Qb97+j
aFdxDIW4BIGJ4M7yCg8/xiJTY0V0X2uCxTCB5CQSRfLCKwEp3T4/qgzDlKuwhPMk
jCLcdWo1umFVdii5/O7opkxR4JzMdHjiK7hidZpHZ+DQii8iZFVdI/e4yRgDCPEL
wYIevH8gj5au4o2ldwFuWJh/yHcsXdWcgWRfpB5kjupuQYensgTzXMoPBZRY0rmc
T39xFu0dGRGn+b41ob6ey3ID+4oMBapXD4HsdVgvKfJBtw3ivO2chj6hyFZzpa7t
FJvcER+OHBM6RnaDBmsJR3sy5wExkSkwsWcyQxQoCwT8EFnrWtYZv+g7aEmR4hB4
T1BNQMrVBgjMfQl/SePZUIqFPSpUJ2ATGgldRfzh3Q+pZYSY1lu3o3NLRGFgPF8L
TYmd3R0W9LJiTzX2rNrAmyLaZ45Gxs/rwEbK3eOAbY8XPxPfqzPKpZE3xEUIMuZW
2J3ifQ0dJTFQaUsAt6NYcUCa6mD62Ze8C1hz0D26vuyYWYd77H8AMmT5sNhEC5fv
yxSFCWKBTUsd/J2d4CxFdzGjACE+SBbaY/JBlHU4UgyVH6R5XatnbmXaW9Sd9UAe
rrpa5BZ319uliND2hIfntO7UHoji7VxXsuV0dYF2fvA5tW4je4cLRcq+bU0dhCZR
+lrGaHoiOwNWjRaMmLhVnzm2h5RTpj0M+R8wK/pF31BB1u2qB4jeONU3jNfDoqNd
tHuAHyXyMfFAvISWfHa+wxtq4hv/GKcBFxd25xON02hpBuybUhNOy4VAEhAkjlXP
7JX+Z3zgLJhVH0ayNaHsawuxGY8rGqv8Z7b1AFYw2Id+1SMhfdHE6dOcQdWe8gpa
FdWf0wVVCya6BWAikRzgj0jnUzkWe5jJ25JoMY/G0n6rHkfPAIUeHyjzQErx0gMU
H7ZM6T780VvNYRY/rAqmX/Ke3b0vBAhUAzDNvuMB8T8Wz7bb0X79wyy73ShX0rhO
3TBCY/ezipft9A7bMjfGn2hw9rB5e5baykKyhpevdrwM3XD9LeeMnhgmrJdhhjzv
HyOtRLqK64vG7Cg5ewy6MIfBghEWbkbkYfv8elCpmyApBfO7O4tpr7agB7o2ez2d
0nJsIe2L3diU3Hqb+NHiKYFxvtZv39y6XxYucHX0hLixUG2/VjTIw0BFpSE4YgS4
Y4ytKsNBmcMDhvsLqUZyfDlL0U8Ml1Ibd0ynyYYhQwSsInyotxHtLtm4d5A5DO0P
naXjOh/Sp7tnbzLeB13NeA3r1nTM+kOLXx90tsHR5BzG6u8rKdkSC8M9nV/M3/tO
I0H/lh538bTn5ty9/CqcgSQfUU5xlHk4jXSOcDurUF4tAEOiIjxOlkceeDFg0kEE
XAD7MswpWVhadEXIq9/yiiAF1B3b/gp37YXDNP9kcbxpDt1IqxBhLU31ILGyBB3V
DTwfd92/VGpPBAyf8vmVusMfdlnLftR9knN7P8kRP1nEkgq1rg5zxjgb2Jqm1hKX
Ybm6K3rMScKCH0vzQXIiR5cgB9tQhQbLrh1Ocnnw2enHLsRAnQ+zTR+vvdDjyAf4
F2f73CiW95qk8XElHUu7ontJ7w0yS39iGhcR4qpWQ5eNVLNODJ8Ek5Z9dAR+kbm2
i4JNh1uHYFpU3lc07rXDyVOyJ9Ei3aykuBvG2+dzTjHuTJfekRkUhAV337I/ogTz
bl5OuUuFI19ikzsHdGNkKGAKzYRQWVNmGx6VzsWujMs71PtIUTzbO7EIpXyPAbRl
Im8djzGalnZhrWxZGtnuxKP1X3Y7DmBLFd98fRnBdO4+G5QfNVnilgnzWqzCoDoC
iUSIuRpCpo2BxtbfaACOr80NGblX4QorVdB6JNntTaDDJT6WRL+N2a5NTLn8lYNy
TCOCF6HBqG8HZTC6540lO1eER+UOprBdFt7/bcUYzNLN4JtAZMar8bRwH6JUYMbN
39tznxUsIrZ78vUe5gEsltJwVrKSgKtjuPzlGIUyk+/wJ16nCBmJ4eA1aE4p+jDs
rIsfq9AGfrsMX9MdG+9X9/CzOG5djCVpngERhRX+hTy+xhHSNRbmVCjIORSpPPaf
Qec6dyi+TMXJERJ/gMqR2vu3nfSQvRso+y7ATocvHh00HbKhQ3QDHNnBwXE/xOSt
HogU4i5byf6sQCw7oYuT3nwSVsSZzOSKr+yPz2rW2VmXdbkYhM84ks2BjDhTPBA3
vH5lPGhkt/YlkNBH/GBxXBgTDs+1/OlWVvDE6cATJT1s1FkQyLtBhX4F+qDHx3V7
O9/F1kvyjWgqlFw1HfTRSm83Nl13MLPuujYfzzwDOqiv/BKI8NZ3SZ6KzWYuovFs
a91jAzRBO2oDr58KvlHfc0j8HB74C7jvCIfAxQncb+H9GV//7rPfTVZJ/9mCI8Bm
6kHkW/eOppRw2IdVo9R2rZipEG6ELfldj4na7/ikiRi3ZrB9BjfhXTUAooyNhDCD
omHUPe51nr57vNcV4+j4/D/tbu7cEABtSHUYMTS4OZrJbGxnjAxIrDAWZgiTUyUr
oqfhScuTEI2doEr7ivHIMMRgtGQP6toTecR6h2aAmrdDH+4tzzQHG3dzXvA6w8hY
iye52Pw9CKhHUm3DcD1oS7Tb+FUIBElh3mOfYOWKz0MW/B6LZYMdRu0REFlCqwEb
spxPaGeB5IsGhwdFrc3pgCoEnmTK3KHnrayeWhKfxOuSulTJBe/7fzg1V+Q8MIgr
e9da47S/IlpzATcTonnBozy1t7CYaC1Vo/rT1xiVW9EtWeyKPW6Iys7aEo7knafp
KbwdK191+Z4AEaX3pm1HvWDaaqDnMTjAMwNMybkxT5LSu2FpgWBoOQ2ywcCh1NH8
6FO7JnldWEwpDN89LYwEulK/rHgaBilO2w2iAuvdlPGrlC2r0bh2tYV9wuub3ZmQ
+n7ta5WcnBLMonv7On5E2CxqDn0ZsLyQZmhdEijEim8LmHFAsRoctKcypV2H0BlA
/nlD+IXIfXNIDUaoaAi/PvW4ly8uNqTaZOSzew8u7GNMFQ7ABLNQm9vSAi21jlwW
443fWU6nt4fBDQe8M76pZCnv4LPVMmZsio9nJeecGUehkQieiptSds8SE8BVkqxK
kNRnsLXcz2PWaVG8c/7wGWnfECeU1uj2uYzPNPemMonXXDZJ9A5U+BlgxFvdZYn/
QZti1iDdCWLqj5xWRgQczIGS0B9OfrcIJCVAp8E8aAnikVo32lqUlEd76OsJCQbS
l1tEe1NDh+2Z0HcYY3RMNGVk8mauz4wE/8rCXZOd2WE9gIkJi2nozx1fD8EhyRMj
/Y/8f7mtiY7rGoDqmh4pD33tv7CLCJItbYFlcKqEZ5qivWxAqrkdBmbRTDAOT0Wh
5MnXnxRMSNMY+bQ/Zay19z0iC16GEPhqwHs75Ixtxd2xsNFPExFa8KPeULuwHd7d
kMFQ062Es9spZefsjxBqHxKSws6cXZvCCLfRvvQT3B0c43NwS0UzFrwgXRoFBinc
l91yLAJhca+UY3aek/Sw57riu7/F3x9bkp0JIevCz9/bHPOmTVRxclQbbtvs80NH
DIHs56ummxscsjh3Uq8yTCQ1DKKKZ8eMoksstPjqEIpRNTDLGqIyrlU/nIAKCsNM
hfKD5Bp6AtkP4ZorvyKnS6IWcat7a9x3jYFLK8JOt2faASrFAtv20uJwWMzHZZHh
97utfNqQIUAjgKI+CxFPlMoJxCNhDPZH+/OSw2Ne/GRXS9G7soAB3PUdLBDGNLNX
uYLNIpRT565bJ/GB6EL6yanXDEJ+4mJEib+UCaePc+vCn6jfQvGyfjKExNMXc+MP
8swen8E8G72YmgUT0RVzHuopiHcX+JVCIADkpZwMRYboCkiGsKRZsFjTTDNau/LU
7VJZZffAb2YkdY90qqtBl9rPC/6n4VuKuu07M2Xmykof4NfBKXqqwH58gK3n5l7x
MKkJBLcQc4bDtjMPU0ZlxCzJp7tPZKHyIV+xI8wZKWEKtkgOqtf/dJtlwoldYEUR
nrex6htXNKEA+4rV05PX/jQx1FpbEGRRr9TJAhBaNAe6kvcbFZkFqdFmVn+apih5
suVp8T0lKciIDoivQLHtUjvVXWRHBaPr2LAmUmoQwqL7lj5iJssM5y6Q5gsJsqM8
dNvc/HPNtgFGqS8wo2TOM6xyJbofIlxBseDDwc6t+GQidTFRyP0USEKzNAAAXb3C
YKdfOsBdIiqJLk2Fik/k+qkQ8M1KUrrsYsp/ds1uvJCh/cNGHrPgnRX8QMsBYB6k
CB5ntBkKny39qy1eQsA4+DSBpyh1xSP6+jmHZk7/4SH4WCk2snSnNI2xC3Nnz+zO
JqPl/L8MLjKyKd3R35pcFtaNtCrpyWlqhY0jVj7sKJ08iXmX19MZuvwhRNrQHjDl
wuuFia1GADXZbqNkX3tAnLnZ6fHzHDD5NgO63MkbSKJqyvJ1B/2RDIfNY0O9y2Q/
f2p6L17qYYvyr5waGSn3nZ+wypdGssjexl6fehRannQhB2US5ytWc41nL2/ZetoP
tJKUFn+6tR6CpQkTNSkiwj2qa1HpHCToltAFOzYpPit7QnwNg/q0/VTIbsupPlUg
DfZJtfkpfjY7iPt79E9pXQPCjemL7WsALkha5HrQliUNMyohQKuNFZRHFC3kcy4u
xZpfZjqvGRxyNMc2yXfrXLxJj8IB5Udcl4pBvuogC3DN5ThZdaGZBnU5wuZoneal
MNgUYdr9KKiccEgZpJoBRzbf8Q+eX93lBe6yPA7Tk7by+b+Zfx60URDbT2O/fa/g
E8M57/HD1yu1RXOx3Kb2Hz+q+KDkj4PMqi3Cr51kWyyGiLxKYFBT9pFipgqOLUyL
hFz3yOs2cTjOopeu/qWHDGTEY29/egJG3TtRBl0Mcl+fzoYUQnb5gKvWLkn0DMmD
fzODVUoDgezxUbS2EKiM0SsQYQrVI4TNZYUJvNEM92XFWy16paMYircFKk/1Ka73
T6DMcJ+zgNy70uiYqsOLZxTiR8pVZrj5zHAY4IhBp5riuj9VYMjmMoN+fu1wzxDn
pCKK2Qck8QA6dZghjfyHyxgkVZrJdl78vUOcGyU6k29fVmU4kklooZadA6GEBh3e
4o1VUbbJA45ybIJQuEBm+uJjlMgXgECmJ7OO4LjZVRha35Ueo9weEhjJtd+raBUE
lu/CL9ODABCgC+W/+MJdMvMmEYA7XS0An5kuzqXIZOJ2b04Syk40SrljrlIfRpAw
Rmpy3X6iL7A8h/N1757z1U3seD6eu37yF81AzvnWXd54qXXo7mnkK/OoIix4BKbz
SkkVqatW4LTC2C0or/OrrOW0Bk80Fu9ipQQ83qv92FOjDU4C5MRbGDVgS0DP+cu9
gT6RouLkHBrTNYPwzeVAq50PHlHCDasLG6VGcy+SywAVJLbgwHszXsMTVhc+qAdk
lobs8unqBxYI8UmaLcc8W3EWZhRvhTs69FrT8Ta+j1waPDpghknSo5j65fIgqzmJ
Cd1kOMH1P8spkQLZ/SzCM+qiWZ+dxsxADc++iRnCsTyP7HLJSkFwR2hGAp31FqL8
UAkloTlc6VooY9aTUD/8t7U/w+CIBOzyNp6E64mDNENx/cg5DgkdgZvnonugvfE+
B6aGr38hszO+ghONTvwYaabxqD5qK6i0khboBcqBgT2vtdUmmLGP8tH19OfXcfig
5A8rKzoS+kfrWbMMc6GBLygxvh0lluRc+rdlrbIFeb0MGtiUV/6otBs/S8aYyuFp
rv4/06gXA9J8CZHGfAObW32+fLB1tOEMr/LMhBImSvu634Sx/Ay/a2rIqmZUY2sc
VVQfYkAXKoh1IUTjXv03jSsEfHYK41DpNGC/+wy8aD2mD/kLtkcJyPbIZooRcivG
GQP9mQBLTiRpzV+wql4WudNdJudklpPyZCSR0WmC6gTBCtEEslwzpQaXLltjMIM9
z4jVaYKefr42zZ6A7JVqIyvC4Jcy9kgMpDN3kLpYAzkDJ9gz7eZWTJ0sf9Sx7bnG
q5+EVsiV9VQVsJ7rZ4ZD2YO9lyLLJrK53IIVsS5Px+X/W7HAmExXGqwZYeaaHB4v
MOXjl77Tggxv0xzLFNSC2WqAN0d0FDckQ25vlw6OXfoo/uxTK+QEFAEwiOWKZgQ3
9j71x+tkrYQ/0fB7qvrENuyM/NAN3r043nHJO62EmfEGC9ydeHu2dOYdgOkVKUp4
g3/AG0ayWItOogRD1g9UhcECU6BXYhMK6QN9738cinREr3VtadMkHZZFXdQ+N8FH
lrJakoLjG0M4/QyxV5unlaYgMZ+TLDc50UNHzXkBwlYLyzF9NmZ/j8NNoKFBYNIv
DvBZTPOW+7FSxhfJvAjUfjuRCxPYrRYIjSDu/LsADQJozCNqth0n9NK7ggWMomlH
Mgm7O20tjt9TirleLBCm0zagCoh6HTx9XxzWg92T+uRdidftZxnpCuXDv2onFjE3
HGrKPFt/O/la5FO0enCP3yByP4WH86ETe9CfbHnsxk11tV37bnKbrbTk65Zbfkx5
1Be+XNxG+/7X+B81iQg+u9yyzKfK+jRgALnCmoNU2Nujr9kNxu5MhZKEEpUwt34U
taBGcww7ghF1B8pmWEH2rxB2jETQuoV2Z4itRKfZWLmJxq1i+H3SvFSveIWa7Zp0
vk8FI+D+XxRyQjHHNOqL/jgjoy1KWRlk3WgU4Rw2B7u1VJ3u4+3kR7rWB63C/erO
HoyLRhBfaW+sIaYCYH+pBrYBzCRZhQaMTk1sd7JllB+nJlvCyO/CZ0NTajBKLE7n
7E0tcHtZiViSYJqnA2N5ce2jggiRq+fQIhLHGlDS5jYPndkQV1APMu2S5rVZsvh3
HG9fuFk1u1Qmeq5kUZr9ZqylQOAZwH8hfpNvpEQEQ+WKKAuRRObEQ3FtGL/KJVKu
/C12a/4mAO5EQIx5igwzGi+z8evRCAhuD4vFhD0lFuEn10StI2gHMe+9UHg/4yx4
xIr44Uuu5X6DHKx5P4l9ldxbwco0efyDP0PSqjuoHil0CyCqYNcpJ4SMN45nyZor
hdW1YorBchou6ONkuTTDskh1S9Ok/Cro2wSkKDQoL45BaZg18yEqvazbR4Bh+clW
fK4WXZGXoHl+phXfQxeeIQx+srjlAbkpcAtozOk4lEFMnnWUFYDzWeTmvCcwP5gU
L9Zetv40FGRiYUQNC822zPvy7+LyRqOaM9u9BTseyqdLCfU4zsHELqOSr6bhqucb
ctxRakoAgvPn4+gEvs15Xu43aDvYK3bIBd496SgwREOhti4AR/M1vjqwNe/MQ5c5
FydtuRpL2Fsc0KRcBncRogJoRxeFkW+CKqBxZ/ZlsgShe0juN2l/gm+uyCAJroFG
UwlE1MDH37JAKXjNvq9yHNt4YWg9q932AdfZgD4IWeDVbUJhfpc/qcywTUqmUQFI
1BTp70y2XoToJ7Em4HaS+Y0nYszjgzYliqWl/IHQdjGWbIPq/qsMO1SyTZdTntqm
ZbjkxGo1+aJqm+W7y92BOwWn/bykVBQ7V+SoV0XSwLWY/KpKHr1ARMQkWvQjROfm
8d6oM0aO8P/7Ggnb+7A8kZB1MGIV3PUsF7ZjXUBfRKGXEdIf642nt+zCW1D4KsVS
V7QOdbqHqgSuei5jz7rZK4UZdDT8PJ5f8S9Lpw9+aZ+ySZlhCiV4yEEFDMbMEoVJ
dWrDQ+R6yJ0YrBKDFlP17cBcxpLVSXRahZmKmVv2CQZc+YIBOBMojrVOMkPR1qRY
RpLz1/SNvI89FGxs2uRUt1E/jhr+4yvzG6huUJxx0DRaycY96K0mMK+vQ5qE4TV0
8gd5ukI2GoH0Gp1lRqH94cMhAgsvWMHD64k+t7i6NRV5d/SBlqxaSr6dCg1IMLmi
X1h99KiUQmXHbrVjsxW7pvES6AqjgzOOGL5IEmcx5IlwduVSicEeLmGsdJ8cyJYz
Gvn1UO44A+gKxihQVNATG37cfRb9wHmQsEhqgAtJaRYSY7CEelrlPRnn0Hel5CSU
STqM9ti9fFcgKbg/ZdCd8klfcYHbVnAUXDc+WdzQYKieRjzwlOHCf7Ebw9t2X79u
ggz1Ybm4j4hQhmvVW8yqhY3M0QsEgM1Kf+yn9x0aa7oC93U4NjYVvRhixzXt/Q+X
aDkgHziRIKbqw5n4oDvSn75L9zeyCowLQyl5NzkuHrN3KhW8aim3Q7jM/Mua3HiQ
YIUWtAEMCp5jykGQk2wZtuhFniYuBfQdETqo6wLAQmTR+3v09G1aZObhyWq5iFgQ
hqal0fM9kGQ7e2Ts3H+DHuz0PRrTZa0ZFMJXuMlL3F/t5Y75HS62w9Vr8n6P8abs
6wLzf083Rlf6zOZTvoqg3forvGDZLq/rd+6msqYdWBk22r9H9PhK1lVWqCT2aDTB
TIhe73Yretxx/fYrHdCwB8ElXd2KwSx5rVpvhVjnk9d5pkfKKtEsLzj4COCfGuVI
o6IJqQcVuvR8uywJWmnefGYfFnOrjLG0DJhxnoubrJ9yT9eU3/Udq4ER3HplQ4iK
9FcZd9BqUkW/at2Qzqz1eRgu357H4kbA1f/qeZubCXQYudTV6NzkrPStYocK3e3P
`protect end_protected