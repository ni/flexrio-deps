`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2864 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmWdo24EC1SLhDeUV9o12ewQ
ulXp2xSZ5P2RSggIKJUy/bzIIxK4ghZo//iC2nkgQCyMSEPdofNGJOO8PcTtBRdd
xDISyRQFTfMHP38fsNekuOOsx5yW90oWFHKdzzOqoogMpZFfCs3Zeq88pLCo1bhN
XaQTZlkA1hLk7f8raFzYwYmJOcVf7++klg1sMbBNz6jHNt2BANcVU+gLKgEYw27g
ADicSi1VuQL1zGQpZsLwRhQTIvKm8+aHvq68Jlc1ijpGP1deF2sSbj2z/PFoJXhF
iwmsWPQ2fm4j1iBoeYstWNgn4hIKMLscmpiAuURttZKIHjBlRqMDKlgjQ7jfomxa
lnIa/dKVuIGPBAfsIvkvyyYFp88NXTSE23FuqmVxw4PkDryOb5ReRnsojH4sv34K
DwbZRr1x6ogJc1Ougm+JcJiv6DF6lyFJQN9chrGpSvmN+SwTbCVPBIE0FbN8BUFj
h5yrqfTSENxwzUj2M3GebBQqrw/luK1enU2YIXc0O9OlEkvAPIk7k+RMeytHCWeD
KGwBbjMtd2EpMxHCKJX2wQfcX5wUMYz53uJqLWmYOJVvQTWrvWMMMULVbCIdxdlY
yZx2cQ1XxGqeGQYtErQ20fagkaeqgrwreTHI3GhEfwLGGIuO55JMhRLZ3wJr4X3g
iZObV6QiPJimU+KD8hGnWGvdbDeeidb6123xBq8iYDw+vUTnalAmIh4VrtyCSW46
GfmRqK6W+TzPAeND+Lyovnn9rvFUnah5BqlrxcSVtMCuU82BfxG5OC3CLFZ77Mbo
yJ0E24cio618pgPbrfI/2jC3PsVpb70c0QXKwMDfCBABzPNI1Ns2LKOzJSOm/bcR
1mdYMyb8Q9UVZmO3v/9QCEdhdjtU+w365i6AVZv9XtA5mbhbhCWSZdhvMeYR1Hh+
9QlArwDxNspO8w3UBzXp+xF7hzrEQsYE1I6Edo1kfm13oqtEK6TMUTRK8HHsaffN
aly05+rnqcgUd15A0CpUMLLL+GbyP7CWCOKNtNBhZk/JMWrEtnJYknxehne/XLTB
GUXx8Dd+KXL008fjhJgF4KBnbeAv4qyvVpYlyk121npeTQH/5l4Fpe62+I1DvrUC
lbaRj8UcqjhMZHp098Ahh7LEsYA0wbhQV1oDqJHTyv5tRSnETPSTttq3NWVLzqN9
dpfU7KJSJLLJbPltZPNo+VAaQeeAKqBvz1SDVVI+l4v1GIvzFxfgSY4li9LjziaJ
ZTy1/xaez3jFsYu5Av+My638JxUfCrDQowclW8dPnSb0fYFj7bBszggWSieT0FoK
Bs/ZE5MdTaWFzTr2TxFQZYhiYnMOZchgTpaM3+9FV4X4dA+55Br1jUAqmC8He2HH
XPanwBhwaI3ryiPPYwu6JvtAAsqdLzNkYgvySTdhKTw0TNy5Dv0jvw0CyToDA9W1
niomCbbBwkmB6qOHpzd/k5Z5YcP8NuhkUdtMnC4wAjwsp+fugPpunoPGa+P/y3Va
F+BWjbVT6nbPxGjseo1fqvPfoC3FfKFtO2lkvcePrJxsOIcEN3Hm1ptFyNvGDiBh
5WFSlr2hOTbF3cwcXPyTLv7kLAarkGCsU6rvRVnKuhV9T60Sk6sPVNpKCWPfIsZk
PQKeu05kTadkVinIlC9dUuRUB8nuBqr9w6oB75BfU1ywXfosxm7emDZS3fYKtdCv
9c4B5CxN0cPJfKZIO61CFswYK0hCzBqSYoorN7jCFe+to4AY0lwExBitBqsBOr3C
uoBS2eANT67dFqJBLDc/iR8bptH9I+qVgjr6MKbYk17ty8WOQnvQ0pSTuGB0Lk+B
ntJ3o89+n6gr7UEANlJtgB63sDp0+jrZyA91lCdnmRp0GWiO2IrWosPMiSGQf1Le
XYkApjlZyf7CvoBFWyPMl0NVlQqTw3v9v9ockMHC9Ubwfb9pGtmG6MDl1nWvHmeV
CtzpTrpjmpOK90ktH+cWsdZi3zJPlwmmReeXSl6GSrJ6xOQev5wyO8a/65D2CRvX
TAbB9OEr7YIVpG5uNvHWGU+KdwJxmojINmTGkOQjxJ4aYFrA18c48NpelgIMlqwh
XlBczykXxAGPpO0Npg9U1bIVO23cGH3iw4g4fnahPGv0vmmL1/3a2aCWFP236Jjt
7ERay0dyY5NsHE1KRfikljaLm0hofVI/wPt0dtfAOJJjfd0rsAbx9oTratihDpAL
kcW385tSgVGBKWWnq9VFIhHaZnvhIXFN6zbBZ6FU4LuHMfnXYXQON+mZQs78Umx9
dCBNxOAeCDG0GinqOlCzeApimg25YRNGnPBs0NOA6E5TUDz/zL6hrB1b5QuKUX6L
Iz269LKDCEIWpSSXPYiYxC6a3+QiWBetIPffZr9rcKGfKJWjIwmKuPt3gVvyVtwJ
48unaQv2ZI24y7rUaqIkiUquQrhgOx2FQY9XETeSH1CcGSY0Bf2Jnm+34TKH3oui
J3tAWYADG7yeniO0k5zP6v+Y3pGNyIKbXdv/2Lfk9haQ7ym53l2fS7UQCmFxsVGd
HQkull9E1IJTI6LhWytacWAgMm4xpaOHF4KuvJvUY654GKtUE18t336P1jLIqnRO
wt6HFUHd/x4Y4Xp0Ox4mhg6eCGPeU37cB2cSS+DsvRpy17Q+G65Ra/YanjRcx5F6
x+FKEZ5pKxQN9OOSgFZr0/bS2zy/SGUTL5/h9M1l7OUMLcdIXhrXRKRb+U5ySGQo
W2GHfQmttjnTI9Rwit3xq28u9SCW039b+zuqXIDj2F5dVmFSWnFMLiFJg7JmgnL/
vpZZYrHiNAoN8eoWCI0m5/cEsL6qHRmaXF+9qH/Z8kMwPDiEVmrX1YehkX7i4Uyx
SKMxiEtPBJVTptuJ4lytGkCclD3vvtPvQo3d0sGL9EgO6GQ4Pzz4uq4S9pmf7Woc
8EaJEc6UE0OXdhUoKIemV5w/n7NbBCKvtYg6N9pbUOhtx0abAjYnzWRDyEx8vGwS
m1qjGtCMfQ/dKh1C2mDXWMT6f9TvkYE/ey7wwGeFWJn51kLfQ1ieNsLM4E/6FKvm
Sw6S4XQr8M5byP2WXxtHwPA4s5JAKnUS4iVovJFCQmMt2BYBBMOvmITl/dexYh5E
yY6Ih3/NGZ/s3EsDVzlKAow4klIauWwI/C38jTKDUo+Ihxem/1En/ZnjU+6SX3/1
H9CtKwuiRcoltYx1VEdeDhosz/pXKMg/Cv5J5Zu0n+EUUfsu+1QoJEN+2kHn+QZa
ACsY6vzxutIjGKLQKGEfpsKzNXtc+DvD7oxgRVUU0gvTdpTf5VSXitunSzQZSuUW
Hlte70YyTIPzXgWlf3+IL02Y9bTa55u3CxX2FMFBnLsy03yvpPUHwMIIyPAgvFOh
4aT8/yXo4BR5Sffyp1K6dvseIRi7D61D4tyxIlq92wNl/UXgPuYSNSc0y/aJZRF1
3bEiqMilZwPwl3cGxmQ0YxgWRQSy7YCjMmXNDompxmEc9uDBqBPD12McCrVmh/UR
wm7ZUwfC6Z7UTFyf2R2U0BgylG5JW/e/6UO3P0nlgM9wz2vl5o9Qg6beDIa5iuJW
gzPI6WFN6JjRe1aKQ0sg92EM682d87csJ2QqxsmaMzNPJj09Q2yQpY6DFIKuYehk
m/GDGjcIDv9nFcwZhyN1AslEjgm4O7Yu90Y0ulztIe/mBljCApR20rGHkGrhqNvM
bAWMQyWvP93E7/ilrqKVlzfg3EjMEV5FYMLwhBCy42U=
`protect end_protected