`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
hVdJHWSfELCmA4ds+csnOQAALbB3ps7EiTSHEDd//nts1r+JQrRE4d3bDPRJpiX2
Sl8d+xAK9BIi4i+3ruAzYvB6kuD7r+gs02Jsvd/1kn7JYK4xBxCjtdDFjVHOTEl1
sSh1oNiYUwLuwR1yKfP+xBhqxD2Dv6pCKhH1NdGilpJQ6cvivGkSunAu0tzP76T0
4x1pB179E7uIeRplfHWX03KzEBF+eVtfgXVp2W1BGjfAe43y1pCvNYZOh1+TY62g
EgAFgbo7pAujZxZy/YSiZjUr2mGp7o83qMXyusx8+rQ41D3X6rxfuP0RiId2pOpC
6oq5Dfkx04a1dk4s8w8cVg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="Sm9DkM+kBxuxXCFA+l3fFkxuSWV4xqRc4Nn7Ji3ukao="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
m2emGBqRy4AuduN4dffN8194qYvc9UXRqiQc56IrQYMiIVQPyh59I8SYabcDdspI
7AFHnvKD5YaF6tQfxWm+mlcmMEk2Y//aUjxeiGGs+RkKgbHitJF/K7nqg1dmKvDg
a/GaBCq4Bqh0EehlN4ntP5HxM4qcvSfh5m/Coe3drc4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uG91daMWA1mGkhgP3oZKMYye3UAomMWgG80HuuXg2E0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 55056 )
`protect data_block
c9NqBF2D1wSep1rW7utzHsk2j40aow1MnrccxUTvKej2Q1cyeDDbgAml4eTSXI8z
QYgCADtWi7S8BeChdv4B2VxKcS7CMq/DaQrOy1MKTfQzfAlK0iubmlTkljLy0Rwd
qPJokL5dgHaoxHhpf4hHttDM3f1hu1GG25HPeYhj81LuF6RVYMO83bdFtH/uYsPZ
fgV2jtztlbmKjf8VP47+Cf2Hemnv4BkE1/YOOIoFyBI+h3tk97AbqZHgKpnBF4Ou
sEUxYpZAwftPPWzRG+nltaOybw6GhtRork349W6s4OstDPtnWosPsLmgaakoijrb
F2ebDQdmX/hbitwVNHlRh/REYnwu0RsIypp3dcrdO9A/tBxTfvonn8Bq60McmBmN
WDZTUwgum0zOzTxxNrbFAm9xt9TgDZ1YL4FppQsdzVDnKbBwrNR7ioMhnN6pfgn5
ISjW9MTukG3ga/Go/xyOMPIcgnwtCbegi2zuUXIJLlrXw2OeVhzY9Yt2R2P21gsy
iCnosTCC7bLmhnH443WphRX6QpcHFwrHkIjiSsfBntr8eUAm+ZSxLou4nccPKMOt
6aGxsbVhU+GW/bVlclngXp8OlnzpaJEhLTIc7ZE9SZdZS0GLOcBGnNme55VJ2XIv
AWowXvsplm71WuHYZU0PVSw0ZwsjsN21j6H+wCAfTOJhT4OMtUW16emSYo1G39/G
Wn6OQlWIuFwUTkAp6KbWfYFYJZZQG+vG1TV6v6MmbMPq0MPPO2zB/oYBA36peJpR
sc9aJXFNYX0cc/SHqm9FVFtOmcRD35ZXhn1CvoiJCrFHMFDL6DrzxrCXAdh93Xq/
vS5+zwRfOXeYZFsf2ESoveOuO8amuy67PhLQ9Xm8hJDusdK0ebY6yuXeS4cm2YLt
McXgZcowj7mCe0nVDoYBPxfLIpFX5COQC8qUbDfXMrKNSgXR8+PY6T7dtw8WRcD5
nNSLn6HjtGsYlHSM/p3YDioH7Nd811mL30B0HFbQbNf3rw7BYOt5idCUklst02pj
Uh88zG6dvv0eakm2BhzxKpFVvICQK6KIcb7nRBU8cISi39bA9Wbeogyo9A7biqc1
J5B0Wwn0KD9Zvt4O5jxiJ6gVr9uELJiNrfazhP5xlJGsVRXl2kRvxgIU5EIlzfgR
r9hfv1CmSgVdGLOHu615QCd2yftPz35PL5JgTeEX2bWzYW+EgQmsd51g/uqG+AJ4
9YTNkfez72IePpvuRwrtWG5XUckK1LVmhbSKAvehv8rXsfhH9GU7q1ZcVRoqjFPj
KOS1VQZDRyxNYdc2P3EK8ivmknhriA1ta2HkmlfwNZPU9hNYXjl02tZud1owCm/p
NwvKRQ4rHclNpLeElGutxXMnJDWgy28DgBNYP3zkwoaBDH594TdUz9Q56SgUE0nE
uRuaCuHmduesGwu8BZwifVn2hf8I8DGepi5D3d+KJg867I1xtbpZDqiNwpp1B/PP
cVvANo2uPufqgMVIjR0H5/A8iH2G4WYmdSWp2bRx+iRtekvoG1vxlp4abgw3/J5R
TysP0V8sJbb3DSJdpT/40kCdflkYW7Z/DwwD2ATi9uur/b9pvVSRlKqKatYhDDqJ
sFmIyr9NMeQButiGril1EwpkxQy01/Qme1vbuIB28WyF55v8yCVRQ5PC7IeYVukx
HpdatRP8kEFBGEbkz3zQRmBRD3QYUjmLT9AW8ICpC2GyN1OqqoEeI4CuENi1A4zX
i+DRMmc1/kILmdvdQzk797gOUtYL7Qgkv2bpx2jqSI4zzzJAYWPJTw282Gufzhxq
EcnNYKJkwRGwR2bqXofLOQMdLACC+ZfBy77cLFDNoXZdZ/gxbMmFGjGmly/jqn+p
R+4WaMPOUghxp2KzqsmKXekPQEzQKj3WsfU+afYQFV//LnjVg/tyRkLpepWP/NOl
QmsxD+8Wq3k/7OZJRrKlp3WYXzhYC5t00RmXVpgBtcVvHsj293VF/fIKRwkHXdXq
N/mA1QyKgTuSGo4xsh02JT28G5Jcy8I+AlsNbr9+s/r99Frrc6T7yeWv4P9l6bXX
037Uf0kOzbiWjCb8d9xrHT+cee+4ZSRaS3nUwawfZa8xJpd9sqQ0ldvr1R6zObdl
zoKpys9XYGWwvIL1OZQ6ZRLGUfcQd7jHPxWsGTji6oITatTQ1eCnFlEzUd27AM4j
9bfiM5qxxjIY3CUHCNt1WcBouFId87i2s/O2ZREosgPZVkMO+jEeR8RuM/trvl4H
fOlQkvH0B/zDRTIjut07GQarYJizV9IIm9nzXVNg1ji6Ey+xfw753LGjrHErwQqv
jMTFdmBBTX2hEDrPBChjI/vdPpgymOoYn6Uzq7Wid/dgKKvCRti4Hwh2dx3DjXWh
xYUREZGqkqh+YsWIBrfETNHjogAmNPykPdRd12u7M+mx6MpPdlgEoZBy/q2cPs71
/oWwuPF+GIpU2BPugG41pLzsKtSVWp81/JKL27Z+jrKEuWVYiNccAyo0GWL+Zvkn
u583G2uoYXzb+N5UzZHh3GiwHebwZEgZaI3r4F+JZ4UwhyiPqFJNjWBmAuAKdMxA
DplGFXFPKP9Ert8D9dhwmgJv4jhv9ragXqUN5HEYNj5gxmgv4XEcil738P9eJ2cz
TY4mvBjkhYiDSScIOot7W5x2VlTZDzFNos4HHsylo5i1jdetDZVmtEMlVCgov90o
BSVGGCTZUu4xuGl7zddEAXKrFHJkmoZTgHqBePkf/2H9KMvO5IwaFgKZRguQhFWq
12LaFXYuWJHOsEcUYd/RP+/11VnBLbJn2mi3yeieR20CSSwSlLREUmE4jKk2h7Mh
h7dqbNafu3bwxb0HJAPmKIGZuthVFCjplkh0hutDAjtvE7IVtC3UIMsGNDzNt5Pj
2PRaTpR36EKRgQ++e6WnDEUNapzZ9WnhnZaDh/O4MqvoO7WAHZdPtQIYbARUaq2b
z6SKw0f5OivxFemZn4QcWsyik6NEGz2tKUfUbbpinGOGrUsHSE74vKTIEFtU4QAm
tn3T8Q/2RoWqxkAYFXWDK2kIA7e250I3Ors0aq39lH46lIGcUb9CELMhxv9Zy0b8
SOlOmx/ogvGdqjtuWWi1e747ULJDsdYPH+WswkQ80ghFh0FPaufr8biT01WjdZEG
vdDzaC/hcMJsZx8GNdhfeaNpj/MCjKduxhWrKpFh2G/hBd/Fcr9pgaP1saX9+i4M
W7/UgeDzwqvSUkwYD32b41bTbCQpCLbvOKeaE2HNLBeShcl65aVnyCU9S74kLIt2
+wv1ZiA0PeQTF6Q2vb2ITIYAKJnNlXQrF8bx8IGVi3Lbp9KtBk9rTt8Hd4ZVS+fx
gzntIdbcYc52EtrNThKOCOEC0yor5o3AGa2ckZF9oIKNrBe7koX5JkaDvcTpQksD
Pj9gV45v08wZdNkMI42WUuoELOBzrHbE+1JGpHKHWAeobwiuSWqO+ICXFrqyFxi/
+D53jMRtvdGgAv+C3Ic+CxoNIjGD5BixJbl4+64DRZJBK/KHd0Mqu55zgAYXIM1K
MoRgXPN4ZfU0EHBu9/aYdkOVD0LvBgKB34JFg5fV6QnFAjuncH36Z+2c5h7bS0NV
o9TqxUdDsDMW0yTGiiQxtHHgol1EQKn2WzRWyy1V5nG6WPWH0XUxTAKiYOuKhrvT
A4wLV/DDom47xOwS1kVsl2i9Biz9F91K1VsN7VVplNdD/iD64setJbsSN8yxf9my
ov05v34zylTTCUPoxNR4xiY7t6utUzb628TgXpcp/p3M+hZJOrEvWIHIs8tkUpOv
cTALMeCJgDDIu1eb11x2o6u1QpX396ywRUq+lpwJllikCZ071hP7/jiGZhIGeYPx
51sbM52AUy3Il9J7yI7NoiwNFotpg+YQJ5z6TmnZZNidlFPIhgCCPL9Jijl4qB2H
Ad6+TL/dqQ1ZhkKZ5Tj0iEoNNnVXY5q4wGuDhAj92L68S7eaj6yUxi24UXk2p/Kf
cXXeFdZDlx/DSNXNg9nCsMkdySBfp4FLf2eSbss6cXIWEG/HcuBELacrYr3YcRoM
d0zypxay2cUZylBeRRaaAhSDbuJKsgjv7bBMWlCsuVR/PbQrXhpwHfROPoUusgLQ
RF71EjNxfDu1vFVwnAslWrKL6eB8bavUm2WxHfdZRjW3moy9SI7FPOb99V+pgxHQ
Z1ykfEDYvf/m19p9arhDkOmkch9walZ/zTMcVN9jOuJimeuvoLqSuMsI7rMACB1a
/nCG+ud1v/zMGDKit87l4ANUFlbaQdi7yRgzI0GGMDy9ySiRjuXZoA/3OW8GO5eW
QUcs9XnUi5GHldWohl0APEqTPkgmuOSgzClXWI01sGC+JzP0JwyNPXJZHIWsj+tf
pjN6ocfD7cEi2SMbd6S3Yd3GfO7vdCIcppI/ZvLzlsfb/tUXMwkvSo1Frme2kj6e
o2ktzN8jnOc1SezAfURgXfjB9EaqenD0d4buy0ZPyBJPa2yEpqAqoQ4OLxN59qGz
6LnhmnK6kPw19DkFT8IgZfCFMttIBSkS7h484A7E6IwN81f5G0Bo+BZEksx+1pWz
uDL1cEhjq1P8F2QFk/ILL9SXkJBF+gAXRiwnlnStXMjlN918FeTTwrqFtyqrkADk
o2EPXqFxgw6gbiO/Hfsn+3yZhGaU1w2aLxexXFNITls0vI1RFR7mERDkFjxtABK0
lGE+ARMIla/BtTbCGYaHjitBACLkEsoynIZDmxAA/WOCSuY1FryqgjdmZX6s5XJ1
7JuT90tI42Nylz7Q0gzQ7ddXcro5g+Y14n7D8c8oPyvOBs4tvg4o1FojpKmn+EC3
Kvlur7BC0n6E+v4ySxdDzBdQLEDpfu/MOzNe7XLTmZuJ5k1TP1DfmqzBxrs9vB0H
+B8DbNvS9GHPoONjy0XMAP5Jh97OAIznQsDjMCS4YO3xLa8CJw7IfwtNcTJhSabX
HPnKvNsOPWmBAYaL/5bJ+j9rBs1RQESybbbfBjPpedb2eWjhomOU2rUN5LWUR7S9
PICSnA+2+5MQadC8NTSoJSIilbEMWjwLPRqDhKcfKxMikiYGNQWDWDNVK45medbS
q1FL/Y3JU9V2K1KVN9M2ZmA24BA3f8q6tu1UMgy61Vh0mzvzl/ZduflnvNwVtcq6
1zxhY+N7aCnRN6oz3dz2vzQbt6RDoJrPWuNOu/6XVSUF0586+kaqyVO+kyaQr/5j
Z7QQmpRdHjPgws1kXOa4+Q8QJNrYMkQgA3k+1+He1utRETjxfUBlP/04m0qJ8lor
8gBHSx9bnmK6l0fz9kElKBPn9IDyyiIM0S7k8eRdsgjpNQITNZi+acRtlYABBdlU
u284KA+5o+eJVb6kIoi0e1I61cARopA3BZH2Apd+ifGcNzal6y0TjusKWbaNuqHF
m8dv1XoLXJa8TrqMN1EPKhCwJ/EKudLl6lH2U+fULTrr6lDbWSkepqEbxbQzQv70
0lwOdXDOJ105osZJbCI7XRHpAL+jgMh8rfal41CzARzrSQDBsu4QyquJOg5q+RaM
fIBmXN+9G4b0oltuITUM2HNhHqsYT0AUkLP+kyFq6XCNI6BwgrNQCgj0fpDT3ueN
fHl3xt0YE4DuGpxDRKmt84mnLP4+PT7Dz4UaozKcLjG+2ThVWyGNVDIaDjvNMlRJ
D1pb7eVpgtsA5BO/Qnm/+cm9gy52dARtZ/bIpYEE7n1wlAFSQClqlsk08BUdOOqO
gQfAtFFAyi9/tVvLF7Mc6oBHe9Xkrk8/Oiy8UVtIz4djd2o8lVo+Wc8CL9cPeIBB
kZ/JQmdimZHIDedaMQajgic/duO9skBMLN0IV7crtEsCHFS35QcGZeowK01IHCrS
Kb65c+idr7zv9VrGLF62GxTYNslHz9qfB7U77SfzthJvhR3Z1FvA94Mjdg76evtO
S8465mUmXexlIl7B+snblVnpDLZiSkFEtPtgae5CCNsoZR5wv4UKsNuIwkw4W2jV
QzlDz0cCUqEjM9yMQ4+3q2EYAmp/km1AMTDirfXACbrJVoSwkTimCvR+Omn6MwBp
wIsthpeJirzj8mFmzV98rui/X8Ioiaf2Bz4gLDmW/BlYBALIwqmPTH0XcxscEo2n
qP64q95vfd/s+zEbNmL6qhLBmoo/W1BdIjxZw5g46Li4vL8z5AMWPWCXN4bTtrWK
OCosStPMlQSRH1hArOh42kbIlI0Ncz5HzzUf5rV3A66T0Tz4/jEc1YUoF4l89PdV
pKlvqDTgYqEpOQM7SIjrkenimuVX/OK2Yh1zasy7t9tt5NMehS0+lsc8KOr09cfH
wi/Sd4MNOJuwZ6xIrDC619eewEn0petilBc93PSVU7oJ7VH72GwvStQn1MtNzRdy
VBfbj0jdzcfzpV7BauPFQO29rSTjpwLmdf4xYMkwUU9WiCBIEqg84OE1Jr+bFVhm
qCiX8JKRkxRzMKoQ8wp3edeUL2FsIyYMY52sjpK53WEbjZEBI7y7O5Fx6Z1sjJz7
IPWZqqgMIizBgzkEnKANkTzRgZAB2F5NM3zDuQTnrVkSeYZnMqr+EHYREHo78uTw
wonRGKkwsUjPqInnTfjm3dPyuOP8HpBTads7mZnPq4RW9ADNnXrajwwqS19R6MAg
qj4HMEqSEJW1xVCVDoqv46rMxIPaUG/ezCwaqck0PmX/nMWISm6BWbIf3b4jeg31
tcwElcUt6Wrj9SLmC+KoSe3lh5xl/PeA0FlUC/UntPxTYGJLtRYMrda1w0SfXCbB
zHweV0koiiyM3PEcYgkxvIAQKBstzyKxQMyyX/RsthnPmv5JD40WVZkVksJZP9Vm
QIjFzbsmPad1+GGm9cYexZOCBOlvOGy6WZhWtBf2DmTo4edCebYr2nAkal2RqarA
lgsf4ze67OJ2hnr90eE3yFcxrAaUjKDhmJ4azZd++1amb+wcEqrdS45Qo+aalz3g
9Oi0oU7Hjr9ULZm9XzClXklpYGybhmJotmSgJz4CUFIXYl7FTQW/9eYsO+z3M8UG
L81yzrrnozO7fwFFxmBsFrZ4XyptTrRbtiwEFSsLo2eagjzQhidjaaevkISTNULL
ZBRI8g7WcmYkf7OFHDpHxplWsYEjnx1zABJeLC94aYQ8HPiVXwSRmyMyWy8WjgK9
Qn1i2aoSyDE1b2YYlyLenkr9eLH8PhqzKmpVU6m63IeOZTQjdNmmTL7PJ1c8WPLN
cGLx7qCT780hu/Q89GmHqnbW1+AALqKPiZ2KNeN1mAtTtxUxjmeOfgpmTSY9XUcO
5aikEX7hYGOpNEQXxboLa89ZemwgPvrGQ6JSxlJXDU3ShJjv7YJ8g+03JlIoOdhn
UaT7Cnl3+RrTxRLQEDp/+QH4cQerLmxiFFRjvi91qkCFMzah8QUWMbB8Q0q7wWzR
mbeYYGx/g8vQeTvqcyvhS59JjecHCRI8wsEWoRLjl3dSC/vb2mCtqQr7kumWVaYP
RDkOihWxrK+sKprt2ohciCWQzeiib8aBFX+iQGpvhzfh7R9vDq/FyVIsfnCZOtex
sOfFvOrTL/my3rPvKDP1UTS1DkPC9/1jb8D68sopr9hFL4p2gSGIUUK3LlhftjBp
JbdaICo8qUF4YEyRMt9dYCXFZ4kgQplXyyy5U4rwUXQPZt8+T2aOrm72ZvI/JtYg
eLfWXiBaYLeX8F/CgaBXsbG4v3cO3S2BvGxlELG4SofXTEKroEf68DoTFiWL1oTu
sOEqV2nCTq/DK/5IkiuzOv+v8pTQRX3Tvo13k96GaqlbtUrKnXMM6LTCbo0GGzmh
gSwJn3CoSNMm3jMhfC231fIqqeCI5BwXwB3b5uJh1/XlzN1A5oRxTHI8YLdTBEii
2IwEABwL+TlZcA+dqK8HSmsGMzB4m57ySU43IzrR/viGZDXYPPNZOdP0913wb7FR
czbPWeVWUJesBeKa6Jg0JluBm68WARqSk2vxkPtjix2NrB748/TYQjmumvCCd76Q
dhrymHdYUFXlGGcy0QOTw73qvY5frz0IHTIIYh08hkY+Eg50MVR8UQWdZ2LTxldc
YPnpdJ23kpsIWN2XwR2aLC8PcNhyZ8Y6D33NZOAVclWw3PI0eQTZBt4LCfaWvCZ9
4oqZl/H8adwLu5yTH+IaQ838U+QGT23hMksZCycl89HRsiFGHal3R36R//hRJZkX
OzmF3NBiXzmUQhMkv8SuUD8viaqw6UB9Kd4j1PI+UdCyTArPL+B8Kv+joGeqgPj3
X89xdo0zWgavUxHjwb70MgfPIq6vrnUvYhvr5kbdGXFQ8SHbT7kUaufY0h/k3i5w
ytSJYFMl3B2/Rp96PYdDETpjJ8gHQ4T3PAqVe6RV2PJ+t0mLvJ61OjsxEgmZjwjL
ZkrrOEbqwZT7ApgOJqxYH7XcBkoiQ2zP5eTyjBd6UbuKVKIJEjpaKodyLYrGH5og
cdjdqe/DoSCEzddojyGhSzoqQFnwAfwv6dfOAIYO/H0woC483yAULQI9XaKRpvXF
l1PJj4QU8EFc/EveABrvNTFxpbX6zOEGr+7XGJcxob0Ma5XOR0Gk2+1nCyBXR/aB
V5HGo/OZafoZwKiILnQkiHTVgOl3R9syx9JTPx73mqrlnC5F8UBaL9Gbmi+AcrXX
4+y0Rd9KlXZ/wosVA6G8k5ugu/as7sdxoGd23wDXKm4WdnJLRZmJa1E8l92nAUH8
0kbWPRVqMKmKWEzV252QrdYOlCbbZR8TSBRXo5PHPCVA/Z3H8AbGwpvjbRALpO65
Kb9qsCe/SlZZO/6+RderHpmvXFpgQ7e0K0kujDIJItc9BCMjldyO2+Jy3Sstwto0
adgvNqt14y+iBy412k/tixiFcGEogof7NZJb/DUbV2UXggmMUZ/ma6Ojz0PQJbuy
M757Vd4Mv40gL9sIoX56yxRiQlCl7wL8F0VXKnkQ9cCqOFghap9uhEs08wd8rdhA
fUuUuhpQsqGzy8myLCjKmaaEKuXoE++TWyoYiiJwk+Hy2ZWv1K3ZuOUD5GzLG+NA
/X1ppg2tgmkP/oKZl9nn7BMxrejkdiNUY+U/zYpvNMfvNdVx+P1C1iVfJV4KeJq3
joqRDKjRh1hD2NTYsPnbIk6Lwo5IvxLBdLyWPKnPqN8fqvMst6x+CNfe3TJyH1cB
nsoPD0NCT+9uYHFaWtuGdJ13SVboLDwD/yNImw4NGzcGlV+n8kiHp2FAJtEjtfWM
MN8Kap0zvv1MDhf4MA4VS8xnHzNcnkW+dXlsakz9qd+xdDaMCKxinl7FcHMuQRa3
PLT12t4z1caK8Onr3idq6Ie21pd0a/a4Spe2xMUPn420QuFYiE4F0jImNQsRoVa7
JuCKU59yrOBJZRJCzBKOdFPG0MiqlFP1zket7GnFM4U5GA6TUT2zPRAlCzj3/wbi
YNY3mOkjcjYW+kQTFI3YKp1QVnBHUgxih7pGOOpcaQcyEAZ5Mn3/caaP5te+NH1P
ByAn2TJ84Kjm/c87zUacvGOAMvVD5CmXctOYO1Afy3vVLhD15jBzkgtD248aDERn
c6PVwt7kh0MlmDDYHRzRtuNbb7WepjE9xusGEifNoBVeckhICNdrsHoYCu5em86M
5SnYZ4mAerLQFyr7fUETcVFLKjo6Vo3VolHOC1LthNPNrJ5jbuTez/kfKMlN+Sdt
xCKHFMQ3rnXKgJLRY/O4IDic0LRaRPNdihzeUzJljj3hAfR8iwjL/tHRqC+WgXu9
11wjoC6PZhTT2HGH3assHIPoJxcZxnbCs6Q/1qGtOBSrF7bk5EHIGJOyuLeXWpDV
/GB68tJOG4wwD2Fxn/e69whChrHcD5QdSECcGbnHPMHZNl1SFZKvlqhYfMcslLYS
eBxrlYNwfxiBLZXVZPJTAQsdm7lnX1hYv4WydyL4BW+5ByFEolAMVPqKO+o1l8pZ
Y702S00yBSjiEj/FpJLAmnpZHbPuN3RE1FqHAtNsLiAfPofHSvTSeuWvNdQ47Jok
kel24eSbKWWmsd2lb4byIv+w1H1GhVRunKMRUtNzVkeMKC+zIQVBjSXj1FDdI0qY
3evz09YeFqArUhpKh1FJb69V1WOn2ums4gFDj1TU/cKul4cICl9jDyIDuE4AQT2l
THJm/yOyMz0FL0qQREcCGA1mmFoOGnARgh9TvtTrrBcMThPd2OPXnj5K3luPm+l9
DDm420pK6zzzJEmXKfZGLGhtgcsBwJoSWHyKsm+v9eQdqWLdXOfDda7rCLFWII+P
YVDhtj3pKuUG1mLEV7FHVlHI+/idPabPwxxPJXJIH0s5UNCpi6oOJ9YP1y4vssPN
7cdJR+SiscRVyNz7izKVJgJ8D1+bGCTJ9rA8NanxqKT3GIEOs8hIdNuX2ShV4V0c
lfVXwDIDQvhlf3O8f12YG5RK6ibvMmSV0WG2mg9w9S5tvRRjsX+gKJeN/G+1jxiY
i6XHuaBvLRsql0idGgAOH3W2A8jQ/FYoCIsWeIyMAMADWInSkHlKLRdrU245qL3U
ddCr/HkmFJZNCoQYZed8DckaO5lTIL0bSGSjkMn+nKq9s6nqjM3sgkdE5ZvXk0is
IUdDd3wuKlOQNtroQpdq6lIM3VRmoqujBNevODINq7JDw17IS+op1zWm/0qb8mb4
sBOR1JAfqLR4pPy0spry3qA8OGOrxHT40cc7uaH5o27RFohR9agum7lPFk/cjLFb
ugzNXJLLxVCAQUtjQmKzxRDfuoUMTUyQyYBWVgL2C9lerZHWfsyCtuUgXMRR5NWn
apOaTF77bjnaHLapb8cnUkOiFGQ/UboT4Su9T889YrY6/OHV5kIgxN1kG8wSMZVw
h4WXwnDEq2tqBGhx0D9Y5DWS5RzsuQl+12zUxgyp8jbX8r01w+gMBJ6iOJpdl3vN
5A+2P3x5vD4u4lLweakjdbKtxi8C0PTBXUvKl2XVnzGPoqc4k5/0HMmj8YxpyVPs
jr1FnNTn8eeLl00fGewqYKQa0eLN8h1eBt5Fh8WU8jnK9QTSkClpoy5vhT9kQs2e
j9rRrotmMVyNDaqIjU4CJnQlmn9Vbsj9CBYSVQq/z62vH8CkmM2CHNcrivSHOsok
RMcze1SGcqbI7MzjFgOzsNyjUXxMoAuUaL4nlBG0vD1if5m++pExLpPHjLHoA1/s
1BEY5zYmkMuvmGWxM2WYI4m8Lhi47VkFpgeIlTovIwnVAwdxy9MWB7PnePabfVb4
BUlA+pvNJIEn95xzcvY+SeF6mLxTD8pIdSX6qfEZZMJxuvCSe75g0z1riihfiWvi
6FW1sSsgNmohKoCi5uXp20odAfxxdL1I74fxeeB2RjAKs1fe0dGdXiwdng9XpKS8
3cot/ezoMq8eD6SIKKKv9mvEcOv0eV0l8JjOEhuIHQr8lQ6JmPR+s1UBTAielQPY
t5iaA4Qequmf0EpdIhDkhyTtszyBtken+o5OoT9FQJumcHXwUp99axC/lLfM42Yj
MG8c/cFpkiUUS++F0bHJpp9nKVZbknl++tuuaZKumExwTJp7O3d96lQNEZDTDUfS
IGrhQ9wYqZFKSvdLmPC9MJ3LGlp+YbUr5s6ecNps0+tSdMM76N3HiND5lduCizXU
IxhafDwSCPeRIgTWP6dV+v8G9bhyfBC3c7yL0T6xYg2kkJPd/fLUDZBuPX9lBzGj
+TIT4WhlL7GKAzSPO7SLJER+pxB7c4DRGbKBr/iE0Y1+jMoEX0ksaJes11PNW/4+
cHHCsM6F8SMf1/tBjyHyzCXneqcM0m6MCezXr1M/GOAagFvqi+Hp0s96+h2YCyj7
s7T2bbpEplqRUq4rJkS4qEpeMowvT5snvcsRxOfkV3IozCWwTlVlg7doTZmcN2FW
gZHbjdtfk/9W7GY+qw8PiTPpnRendsQokgfwIrYYK2TTI9fjZxV/uos9png+p6ah
jakBMrolNPSh5m6QRMLoaVtY8QVUyZi4NNziXkQ5DyMNVU/3o3nxAfqW0436L/TF
/IAj76ZZeGstmfpDO8ZuSzcoDsN/VVgj9Y08yRyQDHKZLfvH14nYA0u6cNaz5LSm
asKzMiMkSXwXNuvcmOlReHW5O2GXVtuowrQylMxw9gYZNWxEpvChN1YmybkP5j87
dSSLbA3mkeNjoA3DAiBi3xhlMPvd8KG4kpcs2KJeEpynimF1kW79c04yQzGY9oBw
1AZh7WdVWsEXp39rVo46AXAGNnxubql6obXBDzDbZuW3UgqUcPtZgQQSb4Kmr2KD
lM9HY335X0JZHSDrCYhJ3S60srvbwbFD7f3ah57n803BNzQ5a0Kw4aiB5jPQxhti
EQMLx5b571xuuZ6uAbT4KRJ53HsTnZLqDirTpEhuo/c8YQAtIJlLTOrrneNaCL2C
VkpXjbFF4BPU57Lp0BTYT0iBb2fQN6YDptQ3pVr/LWYwprtA2dFyCR8Z3SqZuc7s
hVjPsMJ3rsbMyoPJlYONdhMEQfTmtN4anyq/Jpq82aXr4FJc0IAnr3glhQP3WqKJ
z8V1/BVdy9ZP6tEXutaRRZkHI9tQQFLJFR2fCzPvdBa6nmybLFrCmD4jSIsoOlwp
LrLKG3VetsPr9iuMKksQJp9b6DG80d1ZINZDu9iOcEjwXgEZUdWMITMVXD361nyQ
lLVUOzTliq+7MenTUw0fpdOVTVmQlvRnzJDzrq+tMqn7fjxOvOtwPdkbdVErPvhk
vJRNeYGbeb7M11bD2han/Xa46NwWAf/Q9Vc9FY5i6qj488h7jAnUmRCZb4tis1Kp
bLszsNgcwycEvNqklSsnvOqQ/bWekWpOmwEW5db9lPuzpcuxgFlvgyDH8WopO2oL
dalGmtsrFnqnqxCVoKcvtQ19eN7LKyooOfcLcM5j+kulDW9DKnp1GQBpvDG1LtQL
OgNca+uXifuxYojMiVT/gGznJssyykMzuYogcsNkLS3+hmU2P3QisiVsTpJZjfl7
tyQImYmjNSGBIbNyqk0DTQ1KK+BmIRPn8/FjCH3zh2DeyL3ZPgBNareOqdpITHA2
faUSeyuEoAv3z1FW2THhdK5FNDAAy3wgkIq75FwUWt/mdeZGcaZTf/BLKb7XXNVt
kWjUUFZ5EkS9kP50XK75MN6E+qUlbSr5ouXCpbd21FRwZUfSIkjsoKZsbFpV8mTt
nbtG89ttFR+ZNxTuT+2/s3CdbYtHfUNDRFl/KQ6ELD2L6k0lUo8c0RVSLej4g/GE
s6U3fV3a6AXYb9c/K2ndHCRvFb7y6Sbppt+lW2PV598Vl3CoE0JK7XwBDxw6ecih
ju/Y4OGeLsCkctbzwtuT3CPH+d1vMJsi56cCFBzAcc5VpBkP9TecipYm0WIUl6mp
uMyp8e2VfINdYi0t7mUgTf6DehhAbI+aPbs4Re4lXR01UE/BRgq24Pst8lKfBwKd
Y5W92lJ6Uly6CihyGhqhe1f+evjOZRg8Uy+YH9+OkWAJZa79x5HKRMF4b7Z2E4Ly
YEVkB5ScUpgh6gdrTRnRAmXBcaE/R5Wx09PmVy8MQTgYmcxnTByH/8yaJyinmSAv
/dKmhko0NqKcBXHSlXBWP7Im4IEyssmo5+fGjDaqy4MbDNW8XIpU6cIUOmQiw8mG
exBNeiDrddLqLZOs67U6U6DnutpPAVCtH1JyZwJsRLHNuWt+W9B72viuZ9gcOHL/
BLVUa4skGtBhvBc5vyQ4IzJ98W/FZ9aDJhAjbTJ9Vf1iW8u+0dfxA82f3EgKUVUD
k8f4gF24j47MwFwlTX57sTyktEZ/jppPnVY5pHMXmt4yOH2qimML0QKq5UA9ruwY
/W4zYW2lqGH2z0h8hnk4ypBiaCoAp9+MO6m8MF0/rKvKa3GEQaO4ACn1xH+/5eZV
UXgBYS/9lHB9LHE8Fiop8ZjTh4Q6xbBq7YFa/6Jx8uYVSRBmCTzIIU3X27Njrlo5
sCwE03o04hejwC1LYn63/zHvFDNaaTMcRAAi/vSpdLnNAJZokM2rr7nSDEryhYoZ
q/E4gCJYiym2+IMvzPhviUcX9bTfwMc+vL+/p/AZngMYduuf3Dnuf8pUwNYmr696
rIalqCLpn5QapO/Cz/GfUYmFJNiOp75FMi7IqLXmEzKvrk4M8jWUxk97vzg+A96f
oAi2W2EcPYbDr5vrR1L1pzurhvvoAxAe0Vc3MKeLYsqeqYYVOAaUmx3m/o0R/kz0
QBcnmK2vw9hdC+HkNBP6Tp2cJSvdNG0nRWdgGyv5re6FLwu9nITiSA1CSlqJxFBS
0PNHX/QzGGwCi2sfbqjaYgRgEQ1SYqHvUeAq87AiTrOVQGkR3MYd4tLxJZRvwlvV
S1+5GFjxfwN3b5nReo79aSX/C3LH8EUg0GzYYvpI1hSOb3gQPtGm01FyO1hA9ZiL
ErfOk0es7l9uqFBbyIfqtnGwzYREPhUVqsA+AMv8rzJaR7vsieEiZSNRUZIa1Dh5
O4f0ifCDH0iNzhGJjm0CkdBdZgmuQC+VhMQwAdxPkcZG+3dW/zCTj3AKERpUV9DP
ToYWRRLyNUl7zZ8vP661h+FYQdwajAt34j5Bi1Tf4pQDNfCngi6uOnsBACBwQXTh
oy5NDxZOgf3FoYwYCHHp/6bZkyn7kqVWUzo/Q8mc2haFRRopyukvJAVsqHK7I3Ht
ZV+8+6lN1jlKRDBHSk0xKmNKnd4hGfkb74T3QHGF1B/nCrKkp0PyvDdHWZN36eMt
SoX7sE9tg2lGNT+lkKNokgGXTC8agsorN5pXLCIaVxVetSMiwNsOYYmeQZmAptlA
2rBcBnKZnO/GCnQ5IEaIBrlHIoYW8hxmRbspnwhfVMsLFHROwgbeWkE7iTbVDfQO
mI47kZlhJBaOHN3cSJHpFAgjdWgrepF42mh2UhyvA/rPtQsBRtwRrPLH4uE90xlP
qvMSxOeg9pjk8v/YOqZJdoR1xvJtFNeqsTJVpfjw67Uo7zHEFKoeTzRZYe6z+KlJ
svMr8XcClnEpN5lt7FdlE3WJO9PtzY0fEGIPS3XNJ1kFsuWskddiC9ZeHGtMBy5e
VdFjEBIpiYgDEixnQXkAZOrBGU+fpNJqn4fcHO7zZ5Zpg+6+T1x6fiRaZ5i//Te2
mXRwqRq67IGsDXvl7J1FRTysGIEi3pgHDerbwzMKyZ93hO0uDBwsk27Qw28Yd4/4
T2z+CTu6ffv2ZksDxAy/NuLwrQL+R4xD6UWpC6SeecAepnZT3GrAjFRqLNXiOXfy
5STH8lLVUhUgyoiU9Nx8OM38M7ANVAMkofE6PT6ydKNwBOcsYy2HwS0kaYbbPxgm
qhm0NHXU+t8K9h1YG2amIsIVFvwpNVcnahjAjU1+d4DbiLYXNcT0vomY8BrsX90n
2ehDPr41s51lnt8hqYLw8vzbylmBGsMOWaVSuHkWejR+dfVkrETR7n10yywBpk2e
9wLlQvlVSTWjjXjS+ft4pWAdBDm4pqJDgkACsPAZVmls+ZaQ0t2Wp+1aGrRQmSO6
0NvKFy15jqG5jWP30apGtLIjoaZLGjKBGfQqF0CMrjfJExVPKJXl6mKEC7DU3ZC5
xJFXXXXJwmj0t5Sx8dbEWQcCtVG1Zg3Tb8ZD96e+FcQlCFRmeizOnfqzcMiC+RIV
sBi8G4pQ0xpG0kggHyHoaqAO4kTfiRTlmu870YtyNKeaCzTXX9j1dORormwvdYia
vf3ICF8yL7DzjNgEmYE6ibZPIZuDo90KArJi5SmtuNqzZJJrr8naTDI5twO7d/5U
X9ltpwZSyKE2mFn4YLQB4Z2cHnlqTXmZcKVIQFBQsXU+vTI24dhbn2GDK7Tr+L/f
RIXgF0TIM2x/Ne/5b75tkBAv4rYpudN1p7138NznUYwL2JCkdEYXjevj9qVDGVTy
53C204bdmmDXvlxyX8XrxGAeTETYAMQJByqz2k4MPsoqDuVtnX6pxBcytGAvyDfB
B3obbzpFBlu+VijsGvjPRisdYG4d1xCELH/RAk2EmSaDD8+LWD0rwZL+xLTDv5Qx
4H1ZjT7xBK2E9NqLr5DUBuKdl/1rviTsC7ujyTTTdh2+2zIVVkG5+slUo+b97x9G
28sVvZSBgnW+wskH5yhxZgKgQLCCWqHA4E7Hmo2ME1LFZrzKSUepTjELT4Dz5Fhm
LKWHLiVCmd2vbTfVAacVkDmoL4YZCbOgGHqOBt/ogx1YU+zOIl1VrCVVOv+gQQMu
wPPVu2hQbqFArGVoAScBRgePKYuhsY+3xhb0wNhUgqPNzmWNeX6oauBW+g/WUFAC
lzuO8BXwITy+jaiUS1AzlV0psplaz4Jbc3pjjbervDIwaZ4b0fcbaC+7AnFq8puk
JFjaR92mtsUAVsoD1+13PXFkz/lvZQQz7jOC2vdJQXcvKfmaTLsWcORaBe9MNkpF
DM21nE69xDW1MNTfsQb+QWbY09Vn6GPk7AKXTLQ8SOwPBsiG0M+7NpmISrrE7pQv
ZxiNhBtfD2vef7EclHBLARTDDG7dp0O2jWneGhKhH0F1S/JxYU9NlZ88Mbp1SufO
jAWNp3JfRfIF0FmgNLV2J8Py8aV3TIegfpkCFXho07kjcC9+R7jbopJQFyUm6ZHH
fux7AWoPNlHhFFmPXBrVSu3+EUHnVjWHzhOeiJM9JKRQKAmiuY4nQ58AcLIpQWIh
/H1kWuvZEq7rPXq/tpPxaSHyJbITDWvNnoYE5vwEQralS8FoWdo0qDNmbKI0SLDo
JwkW6HTcwSztkMjdLewqVG2gfDEz5YJkCGdWeQmDCM7E9D+QiKVMoIO00h1tWIhl
j3Stv6Zucyrtrhoav4sA+n5+geualK6wUmjOjxClT4CSW7p5WKsKuMsxUCqntpcz
oFRqIouKvjp9f2Krq1BMdTdE1HvUXlg9Y872WurNl4MYfLKCBlm8zMgXIdmWtUow
dTb33VwErBUxOS2mYv5DPdimXeIyix/Yt2ksv7W0CC9Safn2M0pXGCD3xZECVgrx
dRK+VRXsXmv9/bqT8FL6dSnxw8AqOUK3zBv45LE4U1fqLTjmLjYwr/0G4x/y05ew
7D5BpKBd9uTwBkSVDMMuX0JsnmgE3jO2Lk4KD7SI5ZY4keRxey4qAV/bfaLrRG2y
XyE/F/AJW1PkCDRvz4Ztvj4qsDFWuD8O5pTZhuLKMuqOLj8UXGwwje3j+uXZ+ZAz
RyKYq2tmNtCUyId/igVCLHRwOOpvC9+yk7xPd6120r6YebyRfakSA0eY76jLi2mx
L7pqcFfGidWHAOIXwDnygtH+mHb0O/lfdigcLtq8/Jt8XifJPpoTbrLPVPWZNFJB
riA0eH0zIGJdb2xNHWGHllB880178gVVH8aDayvczwMvPEK9kf5ldTnValtUXLb3
+CJaPoJIsMJPvzwjjvoIzkOXGeUVOgahykEDfXJBeeoKvNQFq0B3Ikyoud0hfbAx
3anizaiuIMMTGVVS2EXA5WfPaVLOClcIsBMh6cgHVol2w2gpS1bvNwNcEDcwwje9
bza71b2V0MRpeC9BS8X8MX0GoydXIHOrWeKv3dCGLFktX7m9dbqCHVMFUAZ/apnM
iKePI2QyhpqkCCUQivbLD/jXDNwMz77g4XmHpKhAdtBKutB3FmRdjQjjh4V8Ue84
X7Yj8jdULkLjie7ukq+oiDByaJgPTPZ/8J9D8uZRBoe/nRhdMQA7AW9iU12KvD5t
TvhnAlbx2n3s+7U20DD5tIvxJBjwNjDPeeV2v+4B/sprlc84VX0qccErfcHiaBaY
4wMWnVOY+TvR+KxSVHbjqIyie9JLUUF/MtcGEeu3ss4qUkemTgS+QgKhIcpwqPgU
OfbiLQiXYMIUTFzro+GMjM/B8g+Ij0FjPBZvxeIAvPYQeX1lYYFnrH1pdeeerPTJ
3qkeBxm05gR9ik7DhgUzKewmv2UJDWofxgyVACdkAFJ7JKpcQIvxFVgw6tDALr3h
DYjz/mFKzVWtYEVw08uCobsBdxtwYuaEL/U9H+0/9G4ywodNI31Rk8KBgLobsB31
ug/hZY4Rt3V/9WYY9cNYC13LPZNvLi1lyYM9/Srie4xTeSrCzFeie/xYxCMzTf/4
EuzOx3nZPL/xfqsSNcQOQ0v+OUrk77V+JC0nlmYAduJty7tYeynUtlRf2oVpMbkr
5nk/ri1Ta1FnHQcufxGhckPaPz6/lb4w5zkEdGu40dagDOi4oaA8jCK/klEhxVe5
UxzhHkUIc3UCxX2IXPot3GG3jGcKQqeJ7QGATf3GYznUOfIRtljZodfzoHncwOIW
yqygh+FiQfRrpYek2kwZMG4Rvh7yd9PamgiSwC1MvT9+yk2obnlh/cXVoO03e5HV
1ia9ONk3CxV/iG1SOYc42Q0F7WCXktKdZU0WyffLstc2xGuyOZ9iTedgTQLtni4H
CPf/oLudUEl2dhCrdJJCp4UKRfecq5N+BYJEVGN7Dp1tQs/bsC7V9jEeZlacN7yM
wBJrKRCVI5n/euwG+rjOYtZr8jxW3PtY3WaFNrd0n2Wl9UNXbkHbb5A9jWz7Rtsx
h6DL+Bd+MUXPbWGiHmueaC+kC914zZSy/hygPQi4Oigxf5n4q0m1Megg0qNuWEsv
g/mSVX/RxFPa7gcpxirZoxbaX/WTZL0aBQ9R+/2aE9i3I+Ebg0QpCJzox23PXqYM
3YBPbX8lI2NZs5mF5QzC1mxarJ5DvODahgcMqLuLRH2isyE01GtFg8VdmMAP4JGB
KPuXCftHDEupWHScgHc8+BjXKzmKyml/r35RNDmx4721d4qjWPPQlBa3Ozxh+j0Z
3WMwoSVaQ/b76WWCXNa6w/NNpZB2graTrURReEa+H9HJStYFHL8rgwX1Xjdjv0GP
NCpCKNTXw7kgU1ILPDMCSr2xtakTEMOGRQDC3Kqnlggem9QMhy6AzoUPOAWvhmPA
TKmIuU+EKNdDhDrqKYuEn8vekkZNuq/b2C5Ihz1lvDxIkUWX+qM/OKK/zfv8g9dM
bYy2NtrxHwJsf48YMnm+BDfXtYk0mp98kFwbyIFWhBroN5DtpIXKd3zjdI2pnW/q
gDAF1+7ptLJUV0xetC6a+fMUMlLep1JGBe6iOSN4Q8ELWrjnN+EkYKh1c8jcLf6u
ZPsSvQeXM+sbySArDxAYGzuQFUwimAE0vG+hIpdNc1sq5P7CZqqE59KltoJZQTtS
iR5MAGx+OPiKlJtfGd6PuLva7bzhxUidJYleOXGdTC9Sw3YvU5oksAwZDmRoGj0b
aXWK6PdetB2yguBnmInNYvNXZrxq2+n4DMkfHIcob1pWkJaNiz2DOwV3Dz/pTtom
xjWalVi2kZpHlpH5l37ivGwGnu+7p2CuMjlLndiG7gCT0rtto4AvVYUB+jWqB1ZD
vpPkgizENL/IcIrsTytlXu2T/b6drIrlqzA1Kv6IPHsftEpdgaCjZ0UmGXhQWnK1
EnTWvpVxurPRUj4DlEfeg7zyVEfAYiXtPRQZzBCbSpocpRKpuEvno+i5U8idaxVG
7nQDVK9/YxHtlmr+DoDOuEBjgazy5N8CNdw0qc8I5A7dTgCqONsQDYE14b3oTnl9
Qzq1Qr/ShjNMYOIpsMds5D+bK4DrqexNoCZQ8DBWrNe3ugBeW15fgZAEYMbCPTCp
Xwv1PnoC4dPAByLKDUeDG+PeKHbxU0mVlCKPEzMKu91dHHn1cslBuepJI9LHE1Jx
2nNaYriY+9dlwYVxfq+urBohJ+G4LNBTzm5OZTYrI7pHa+rMck5Xc6hl92tCF94M
slGLXo2tik7EFYjLwoMGdvGMg/EXuZdNdfX2a+myNJTZeLSeilcwax6Eqm5Zk6yX
OXfLFKLz2v4CTrisJCqBKXE1okBrepeMFQIalcLImfNXCJfO/+aALvc3Afs1vBs6
ilkkXEZXwM3FNKKyZ8mAXOr/9CCxQ+gRhXBnPqgdAZUGit+b8wvDXvVE58St9K9A
PTuFNsVGS1Jv39aF/fbBp+xg54wgbphwFqKB2gB35V3LJKEVMMng+QzSXP90Rema
AcXJVpKE7m00EEI+KXz5nZA4GwkGsZtggJWXh5ZgaDj7ZMYw5IIh4+xIRFAtbUdt
ZXcQhz50ECkmDQraXQdVKBCRN+jvVqLEhj7GhAuJ6DeT+ppbll/EkUsTzMC9PMkS
GKOi/B57ahDqz88CCEeK3oK8A8VocAnGbiLKKXnaMtFvqHvjhilH1LLeVHHH0ywH
gAtSMWpfYohyFoI6n/uchbZmH6OpTaCVpaL8vLQSetUPiV5imQ1Hohs7ipKhsKQ7
wgcuqk6kmRfMmJeCZ+fBFG7LpyW6HWiRDhn4Thb/vPlw8hLpAgwybas79QjvkMfT
jsEF1IM+saaiNsOqvJw2X7Rp68wgr61JPTQqxRqErDCWwquml6uh/3vbfD+3PGM0
VJ6YCa2K3SWZroTOUq76vCVXQwLsKkyjJo1vXfZKR2xyULxfnbugjsSCYiUSVxsB
MHtJ+jFLMds+y0U22mFZAfa0xrxsWe+Gt2VkspLgtyVnp10hZ8rpGq0RZhxWMjR3
urMjqUFwaLxfhwSoNc0Inx4SnmnxH6Q1GFzeqFTuRLPWKLCvI3F4A6QoO//i7spR
CTtiIG6yTL+u7vx6yj8AHeepEzvC8QggAjeRIAOT4sFYnmaVA5xI2eqdQLUczyN9
j2YUOwPEUgd3Spyzxcz0jTyTiogFUSfEuxq9DMdhiGg25x++aVF2fiQYkmyegm4e
EkPm1GJ4J7qBIxbEUpZ8f73+Fqq30QNHdsnfVZG2Zjg+Yv3nDibSzA+Y5xPGvGyj
/Y/mNS4E9SmV3NarOJpveE+kHjk8irtORQROE5Uz4T4ddgD/xjH9PzW0qvbPg7FC
iokTMwzoTWfzAON6LEhtkI7CUyDNCPCdvHFk8IpB4I/gM5dhJsSI85gk83tLzrJy
R8+UjbaWhZIVuuVHnG/BxX0BXni1TBNal2b1fAjXv36fK6b2sextoUFNOTztopSM
Hr97o8qfZLbuGFIB3WO5Ou8cO7Qb1Cy3NdSkxpqPNRY6efK1GK0CI8alDj4CXgvy
Clsy70ZuJuwqhQ6YAmysCLer9dcYmmd6u3GTmNZm+JqwfvIS9q/HM8eLJLbKQrVT
VLwxcSHlhUzvTl1xHeqhzazI4gONJN24gixnyqTeiW/Wl+37KzwL3bNt6AG1yeQV
82Bp7WA3Axk5f8MgCJQZt/Yd6u9rEQThLtt/wClvBXMqaMR/USFqPzGr66Rfg2qx
zXnmogJepBfA2Djcx5rE3HbjSFJGM3jnV2b3XpCaUrQUyUGk/4m+effUzlWgyRp1
NT1DfxYVnusU4A8od/wMKTj3KHGesEl1Bi2WroOn4nfDeni2bnb+9+f5v85vPiyD
qWma8r0RFvVqBUJtGxeinS9W4R++tyYOJCY3+7mwgquNeVf74GC0Mbw8DFenxgeq
3VYYiU72RlKbCelE+nRuUq/mqQK6y5FGZDs5HQbP2Qy2LCLgzHZRLb+AV6H9dba+
/ZcLW5VVjrCmseb6Oc9HOTTinPV5w0b51LxrT42tIJv5HmmCCx4brDGsmWo0ryk6
f8ndSmJgV+I8xxF4YyT6K3QsFdsRlPBrKp89ayENsEtHc8O1aBQMiiqTYBq+y6Ht
zvXfApv/xKC8BgJSkzgaOY8hI6Y1Xgr95fK9wP0jCttsfdL5ub583OFJJFaZZSdv
1gAQ9qnIpEH76CI/+2kezlHlZGouWzPogNoPTP1l9vZl8K6Ejt7rooWW0YX9K2tI
i9YWB40TCGuDk2J9HzJ0LqN9OIQj1MfhOwhc9fsgwCOBW1vYXS3GY7pAm9TGdhoe
Huz1KtpAJEjvjy0676VY6cRMrcyptrzUu/NEBZK5noLdk+oPRGpmx6ys1urkliOp
mdzWbPVIedgmhRcYFuteeYrajaAKLUjRCiyytffMzzqnNPnbwG/SaHSY0V4U2Rtj
wDrJvS8mgM2i9iAN0yhl6L80U2cqv/yZWl36HrfJOoEPVCvJf2mlB6BqeTGBU6yj
gXKwUrX3Qw2TGDI6fq78SHehJiXPHuXuR8KUDW4Iq+ZHFU4+Osray+w1o5CaS5SN
v6Xsq6oVCwASwaBhunyLKToZ8QJupsGPIJaSVlMCgfpv4UdL1meAZdZtaq1Q0y7l
kCHoFy9hzxYNi3kQ6kAa1AHeOy1mQQW19v6bFkPkRyozRKkNki5kHEEE4F+Wkivs
6EIQs3AljR6HrSMS1ZtVdEs6jC4ci1tewMz9+HuJLdY3T8cJHWMVsSKkn7qjCbFI
N/kuD56KriDFCk9p65YB1p3Q4jLpyIQL5EmkxKgcgsbHnjpz2Di7rnMVrQWbBfjg
97HYJ5rpjH+jwtKODbQzHHCgN8QAs+cY40g2lAUbQugaZcv+B2cN2GnA87uZj4bT
koBX+WF6LoqdnQ2Tq7A5c28TR83oqsUaulsKEpSQe9GnSmOxxaJh7J/Z6otLSEtF
zly5jsD7jXiUAyjCKv6oyeTuGDBuH/+UbkCChHVUgw/nAmtekXpuMX6KpgV+JEYI
L9eeMEsrLfo0Ic30ryHgbTQ5ad91OnniHpSwRgmBlpZxinyYf5Vw70n2BCaNSfS/
btkyCpSYFq6uYWvY8X5AizxqzalJ1YiGDHsvJB0XtNTG7tN0I02C/gOkAnvEDo2J
rrdJdx9+XI73/sfAAJ2KRQhulsMCj21nd8oMfNRGdahURQ61NiPpjbpekC4U9GHQ
jz/LC9LeXb+66/ayi1iYiqatdVevWjPJTM0jZvOhY06cuSLZMYR16SCUmVLI4DDy
10bdjBEJ/QO/fdxZAcCj8RPQZF4bpMi6Y4rZqITxHdiqfYMBOYkfFFtkgtBBhmjb
nyajk9uNdpLINeOeccr36Lt0zRe10JLGFAd/mlx+kQO3N35bXUcjvNVtrh9U1CHQ
5Z7w20QIJB/mnKfMgsaNnS+MTMBGVhDISthEoX+CfP7owSQ96pbc2Rsdaj8kGXSL
6hj6YZWzj6b6VNtL7JHog3GkcJ4mTib3kLHS+71c2rLB/sirsBC8q+QQs7hUL72a
/POsE9KQktQhjuRbxUmhhNzpEBCbnOYmcF2jvPePw+5vuwIjIHpsWnbM8YGxSGMw
QE29wq/jOmyb110Ixr/B2GGKxzYsO3W3m3oojwrBqQb0XI9zMn1rPTMc9ttS78A9
Ugm6wQhPekBlQETEgUAAR70PHgsf9aA2RNmNhdWfzEb9b4lRh6PUletkgYWzlLoJ
tDUmVB3rmFhEylORquteZ5iJTpm6dFZBt/ji0/lGTBjsgf0hYuU4Bk0j3PXJzdV6
0ult34Eieg3kl4S4cGjn95WyiAH1a935t2YuTLcotuBaBr3Mr4pw9sJE3dWOjrot
BCmVXgaOEHZsKKT0o9UqZ6oJ5bXGzLk3YcvDo/KRFDKiuJh5C5scLwj1IH7r+z33
vhCp02FUhvPWHlpAEfKAqXEEAERzF9L7iB+RJ8Vbrfcti9vK1EifIX4mpm3MF40h
rFToDRmpeK3gx3AkrmcqiBafpZLCPnELnzzAJTnJElrYte5evCvJoLNUP/aFb4rC
V8KX+5vdJoqwK9avjoM5X4RHfjz7PbrTJPx1PugXs92dsBTmSu15LpXY+dzAAhez
YgnfXhu8fjVKg3ksELlbw1S4UtytNcePbhWhIVR48ig41VDHKuhkGgv3qkPu8Orq
9AB4pid6MPKcH6z4dgcrzdpFmfL26g8k16o37nNQ1JLh7ol8aoujOVyzHtTBGao2
J0pOcRo+1qdoz/jGmh4ZzTvKinL+h8Fkq+twp3s/ZD/oUp4IVy4wMvWQb7Kau1S5
W5dwpbGkc9WE4PVaI/yvxOuayYsDbKtHf3TNP3bAZ1EW4NkVwo2BSiZ0ql5Lz/tI
ZL11cyE/xqxn+/Y3FvJ2Ksjf5liEByQ6gNltbABVRWIlMdqCa5D9OGGbXMVazTmp
OLYjkQVBUFLbJXCC8o7XOxAs1BBQKqcaczKV7S7NhKURt/ujH6PqAw1ZGg0pTmTQ
YwWsiDSIiT3J4JCh4Dp6gCakgvh5wJjj2oayAXfyEeci9oL/Qa8bPh6CXeDxKLRc
xPeDOdaOWaQYgx0JYJWjArukK9OiGDVIpGHKBhRnW+3Qo9sdcY0mfw6puB3Ttb6A
yUfQJSDKY2BfcxsEhnqLyVOxkE7A2h+LKIOG71xMAsLSq9lxdYuDjiGhtjKKHJbx
QKDZXoqK5Uw031NIhxJ7lZhdMv/21RxxnReBd3lJgwo6QsQ1E2O+mQPFFA1Jzy9e
CgeM4+94k1SPvFogK+KWonxByfoqwibeXpnazlKo+Hv/gqQEDQ4JCdNpD4JA6qk/
7HKtpr2MVCmoViqt5CSWl1KlTwoLBHeR/1A3ktGtWZkACWR7RjrBZ8+dV3tSle/0
UWt+L2Zrm1Kdxi1Lwbj1XTbjDVtnYDtbvToIyR9hiFN9itzevEbqBzNbvGqGMhHM
gEldQFgTFMXpn6I1AOfdWW95SawiiSOUTP404dTKzb6hSCoNXoVu6Xtc+67yVtFl
iiuNLIWeqrTVCFgfWx+xSndAF4qUqNVgUSkXmwRpiIb51wYDeSrq7nl+X0j/dT3I
7Hl0QhknIMEOx53hdnlpwUz06ErTRfVF6zg4etVl4hD0ba//ugRDT4XIQsXjYxfA
TfjHAnK1WFWXWOQi/Ou/rvnPoIkEBqDuvczxYIUPbGn3u+RJ/dkI8aDQf5hYccQz
f7a9C3Be6flO7Nu1FLogNhu3U6YcREMxbvoFR80UEG1kAUOYRrVIft1l2SXdVG6G
OWsk42n81Fbg6M87rcjvZyEPyU2CWuubBfPeXOXvrgxwAABSqWQb7gTvJ/Y3H/+K
pcSNN9ZCrYeCP5k4sehqekNx7zt66o5wAdoGaGOy7u7slOwBnr2KzbXjYJXNyHic
FTIQyCTDyZX+IwfTTp5N7ZNqyBXK5vdC9prTqBz31UlPHhzqS2Q8N6yDkr43ZiKS
8RmjZND3RhxlmAtM8rUo/uYv+pCeixcQ6PR3IGbVCq173dU2cJ6oG0Oupi6zaTP8
wwIH23siYX6H05vNtjUguaAtheigAWjGb+3t+lWZQNyRa+gCJEJ+Xnv1szh3b1hY
tXW9yr2LmLBozYt6ZdlJoEm2s9qLYObNGfYfxn48tGC3hCzYm0DjIHm1cfZ69LR8
s/W+H655WpVG/dtXMT6B28HXymJmyHWynFwSMnmWvRj08yJqTdWloUf9UFrBeH3x
3dLP8DpfVCVlrXfeRkxyX6dsu1reG3hYIKCtNRcU8vic3WGcmIhYVx9qKwOJ8Xq4
B4tTbBPNndA6SdRyd42sEhiv4giv/JKqlT6mMOhAZhNL2V7VQ4AHfPW/yu5CKqVN
Pg3uALHPPTUnq/2Ma/JLcf0/YrCC16RBrjSvhaswVhRwY4VGaDwKE+HRQ0uaXiqx
+rwqEhkyC+U/gxjw8VbYPMLiFzUQyeV9fyVHEcNs25uUOCz8qL6Nj1rViYbxr+V/
b+3jP9D/26sstA/9WeBCnvTb8Pi11u8ZooEena7Qc7M/ZkV7KriNrkux7cLg5c0A
+d/fjYrsNKtZqoMmzOSIHAOBfq/lWR0TKj71/o0qgHyD3y7r8ZYrBUz5V1r9+7GW
0tnJUl+T8nHhKXoRfuRrK70FCPo8GKYRlezETsDuakN7y866tvyO0YyiHnpZgCUx
gSQFrV5gwzLxWrTl9FnJvn3rLeuVWrX14LJsPrW5f8e0PixYNaJa2PadGk7TnJPQ
UdNvfL7eLg3Mv1a6P5kMjqcAD2pu6DJlpAV2LPP1PRmrwWZIfmfwbRB4/cgQxF4p
q3ALuInWQvSlzjEcT2L2/b/wJdJpzJFF/EMLDMWSqAQqkRzlGpL/kfFCg08gYHeP
evQf0xtnmLNbregvBXaFj3aVbUILtLnA82FifLZ3b9HwPUusJfSmJ4HessOeTdWa
3EwA1ia7p5wy133iM6A90RKXk8cJ8Mecm0JI12/M1Hepe99ODmk5zXgr1veS6us0
RklQE633xunOQpCiwc4Ink74wG6jnjG2zsIkOcauQHyxyTR6P/cmQofIeE1kVINs
vOuIRP+/buWicJXNTRYrfnUeuJPkcbmOkSZ++pAiZd/8nDEEmU6YSxg7zlcLVRZW
y5P0xIYyfY9LChqols8ym0qMT9W+HjX9P/u7EYmn80w+GmKH51hYlmPZS7CQbw6b
Pvm0NtUFAJC0BlOlwk3uJhCvaDNE3TFPL/q+xYPDbOv1st7sG+BgbPDio0SaVEk7
rWy708KmiuAqBNhtdBbfN5nyT4CtWeLoM1FhEDvlFmhTj4eqvVEq0P4GygMGfSkT
t6X20BdAfaufwJrAntWYIxiFyfgpj5Gu4yhq22B8cQPNe2z0468VSrVlPF6a+QUz
Dm5sHL4K1wnOiL+xVMH9PAuOhNxS/ZutRJ/iE9Dt3kiZsoHMDEEPoPnl2E9sH1JG
UE1rG6HwwGbFmtGNsW3VUZZaORA+tTFGxSLHBWtTc0+WM4OpMMzp4jFaCZ6T4+HJ
dhsp9Ao8zX+j7aUXXLiP5xQCNuLru/4hYGPmutgzXxPTpPrtrx+jakWQCs6GidQD
PZQckhnjvsXsosIVNlrntBjNpGYJ2LAl6W+cH0QcjcpDDKld6bw4EZ7ovLFImsAq
RWc8amc+ApTKXi+N2Qx8w4+Wzbfi7zERI9W3mkcMcJ1XQZBLMzXjZwesFQNd/rz9
L4DMnx4/VOZktVKiLB60IRxkz1CUsifl+kBdnnLJLQP+SLW203LD3luBV1h/lOb+
MQQwAxgDjlppH73wC2btZojycOE97hyUsyp+nLkY8N35NwqpqLQsI2sj2eSJ9h8y
lmZI9GbzQ8LuCuA7r1HGxBhTA3/sYFGZ5hNJk5kpPmDGbsoRYf3dmdTqECYBDLxV
QKWHSMRjyty2NysU+Zi2Z1U3IzYLA7vNjXjW9nfTTjnhuVJHyybdrLg2N6bHvfUR
36QYhg+ynlQhX2oGSpWH3iCO9qx6Qy1AP/oIrW4Mr6nrgXLmdzbvphAuTB7FNd3x
gey9MUB5CAW1i8HitEz0QJRLC6GhsK9wQXzFDoPIkbraWWv0xa5xDynZfFY4qIuc
D8B16WQguFgDlgnT7fb/Nwj6fYyaKXhvMASruM2j+IGoR4p5eEhffo3H6fmftLxx
3/PiYFmPIJGQtOO4NPDM/fylqafOF7FQ4nNzpXN+Bjd0aNgdZyy1ln1JYgnem/WU
aTM+TNPwFCsST/JFRvIEtxXPPv7sdivJzbQlMUsaBXCyS/yKckwx6pwyLpXdxn95
hCz5ohOQYP5iMrlsRBeu9ROAtqZ5s1Nll4jRhae4lKKTi2CmMiJpPxkyRBjaEBGo
mkAeQLLnntaNDkcNJvMYnRVv1ch/aXVLPTcIECkX3l4fYfCk4vY1Z1kqkiBodY70
pqIvOQnLoecOBhCmC0X6Qu3AXhtoTaRB6QXdQnr3u4Y9N1Ifev/WEmNBMLqy0tCV
uZ2vqaI//PGRBU/O3B0/uPbmXKQd10ZEM8FQePO0Vjan5dFtu7da4aLv+/IXERJh
zwbydUejdj4A5thVdg/fM4hJNdECWC+OGGSJageUA6yo3D0kD8K5WQC6JuWyb0bh
ZSnC/uei23KMHIbEUTWpmMchLT+CvrnadR4GQud0z3h/Cv8bfpmGZB4N+XnOJa6a
QJeZTcmRwUEh3684/81gaPH5tW81r6Rl0ci7towLQdBO05i6i4SIqw//2BZITDpV
LvKQWCHzMZnqDH+Ce4Inc3BHCFsWLI1zwP620bNvFxH76m/97jmcZEIrVB068bop
iBYHB2AMt5VfvObBrjVfMsjkcXnrWDkh/y0dxZ/+KumYsxWvPqXvEiPrjz4EZnB3
9UxRuvPxBfLXaQZcjjZygswb+XGok/q5v0cQuqkSEDbOtyy5616vMWpJ5D+BspTj
f9Lt9KvsllhMIkv2CcyfKDWYZFuCUb1CqbELriYyMofNkXMH88K42Gr+5XHWOm8+
k9OOCPs0g6qWpOeqsiesGbKDzuyQWWF/ucrGOpnSiKsqD3LPiAsV+TGs5J+ufx//
sKx5SUY/SPr5+hPegDlYcnBLEPZ56YOc35J5CVd9hfvIwwhqwuZ551uMzndclO5S
qj4L//JU702jtHhPJcAQUe9pUKSI0mkoD/JOc9wdsmlpQvD1rQ0T5CHFoCZPAWEf
kY3T3sRLmQd296siwFG/cxILf8l0mJt1YFUQGFuWh9I1UiJQtcdqhP/oUlGto6Dx
Pi3f6gtfVTio+fbEQ22Ul81wxU1AR12eayCw2jUbHxbgHdIBG/vvB7neVDi21jXl
SarD2xQtS2rTwo5PvhXbjlXdQwuGk3hvLE6tc3SOXUDlKRgXK/9pBT+n54hfRqkh
PyIWT47eRUpIH34a2jkjh1IelXW+i1QHLLmBcScMPwOy/6ZQ2036KTWI6almtzHY
UY60Xs98Q05z29Y0hepPLbKEwEwnEsiosDtPgPhmYAdVkeQtKo4BwNUKl9eXZRdp
oCDeDMe2CKXDme0qBNB7/T/ufnjCky9IaWmXtXlUKeKpynfXisEAqggMF6xJQZz/
GwysmHRDmR0RU9ek18mrTPsWFRazbU87jJiaaDuLmhg5JHM5f4ztr3EnFxX+LUwL
3cgmYC/xeg1HUn7KRQoFSMeCX+hqOQg7ZCWS04xf4IuhxOHoJQ+RY6z7ZHBsB20B
XBuURpvFLykSH84WgtyzcBB64kWU3jOfw3gwyyfH9W0rwJTsI7vyUmO6ulysg87C
0E32INt4ukKJDM7a8yZdG/D1YkvpdhxWcSkQrpTwZxjDCBZXXAkU5qrE4bKIaHvX
cHqzshiwTOOa/dCX5Or3yRSTxCy4cvzXze7RN949FV2GIDhouyUHO9Qpx6YoXewd
ytNWNq24jHyj5PA64Uy/KyDj0qTtqYfxWXiyN3n6+ehjCDT1eWcEPvAwZpDjZi1j
DP0lzIRrfcjGWd2poHQhcbKd0xiT2t/i1xp9qkBbsvAo3VIiRGpXW1sxlP0MDoZW
rgO9ga2Je3iORw8F1EQ6s4F1MPpYrEg5ilovTW3bcdZk1gp97jlwyJm96xOkyduP
/J4x2zs3J92OeXVD89PC5T0v174UeSZoncj2SsSuP5B1CH/tFyfOTy14tMltmgkP
sY1ODceeFZntUPYmuEGO0sKO/eaTvWkzMLwzmTm6mNr4J4OEe3jUniGI6ArCiDi6
BQb4/RMU7u4mozeg563ftO9JUWb8YWTqicfJwvewBB4xIZMbQczsPdj4eYLnztK0
eBLMKoH7GGm9rYcX+yHMBHG7UFbKzzM/YCs8pZ1uLVsLaUb4Y2fASj9tvTOd02M4
0UcWt+A2MidYzVjpl19LVndSDlCiK83aWReB+eyulDd1GoNe8clXm6GDukR/9E7R
PLdHojX+NbBL3tgV3aNdTYqWFZbLOUjdt7uc/tfwlxwMJgA7lwNo8dvY1yYsphGy
/gugdDIeMjFzChYzNOQwYfYlVjdzFdGm0aDLnpycYDuUFXk79s/UVeVzjFlOR9WV
slL7tQr4pKWDCSOTBIYkQJgeE1rsysS02b9qwnVBPBYYW43KwUk1qVSkOG1z7bfv
XFC2vpDDNH9p6sbyZxklbkwKef34W0Msepm786R1wkuOiSzgvtnCZy3RQgTpJ1Kc
2YdZZqvvsmEjhphWBT+Ql281O6JRtHnJ9ReVDOnvTbeA3yrYgtZrUTkcbb3giLYe
fNIfMt1dPl20a1pTHB2gvgkjTdS7YEItpSmZq8vtVqyf3kySgIGvWCGMPTYo1FF1
1c9oc5ozSMWO7ebhpE04pG21DylwpjiGM05Yd6rMfpbepEWj1guZD90q2dM1FKX5
eO2JcOuQh1dTC/1f+vhrbRLx0D/saWe3DATivei3ccoh+VA4HpG2bw3QsrXmHO2E
ZIOSkVQfXZ4UBY6XmfbsjzXU5i6eNjwXMnpDxACmtBA8sFQu54tJR74wg01LR/Nr
2NPOC+U4YqjT/XGBGUxSS8vOrKcbotQydrC4uDeWN+fqFmum04ss/wLG95XJszC9
gC4bI1yQfMtC83IWWgX/cTC3FGm4oIZzeYnZGxknlzeiq7dW1Sc9oZoXDXkXkgEy
dZPW2q/or7BLBS2rtdFkiAUoF69eR10kFkYi4t/ZWXm5wgaF9wuQd5ZZ/DyFDJbn
9G+4FU548aYGV5cXDqu6Xcl7pNi/1StXjSn/bopToR5VCfDHQsv3/akRuh3XpRta
6LD0MbtGbZUANubZeaeA5YVzI+HVUVUq4ZZGtz8bVArg/jvXg8iCx6lEJiAqDRQg
4AMkBOKsqNZFR6bd6PBBZuSosthTwRu4dqIgcW4FroEUiVvr218pAgwU0N371b74
v2MCSh6XFZkFk3rDjIi71Um0Udk8pungZnKcSrAcw3GSfPj1qpUfDA39egqstxoH
K+7eHxlPRCOY0F9ctpclXp6Q85MXNk6OqWqlDSWcZLyRl+xsA25VvGbreSOh2ygg
52SITZ1pH5+1OYec00OBa7N2TSevh2MnqPEYXcV59OrwjLtpeZnljZfHthJP2F/Y
VbxvZgP/5j+5I2Tlkk9sycSVivBjnwBvfBrIswhIRkAZIq36fQ5jbXoiLBbB0MyO
b0PnWE09zv0LWgOQGxDJBi+ML9RJZv24LQ/1W8AEZKAdYZ/AVPCyOYDEBnNH/iDX
xnQ2pgosHb4hGGyOS7SnkqeW68GAn5ItDUKVBN4zEbNh9Nq5/3csfBY38tU25zDv
M5mlrUrv4grPTPuBZeGgFQr6zjXPR+D77KU6q0mSfPIClluFRlqDEpQo20heWnjI
nApSwe5OCTO0eIbMkAsC+e7DZs6msaRiMC0KCXXSnfGTq3e8bJJ5hNMlii6XNroa
oDD8FKj8HoaUYYqJvQ785cnE67k2b07kkxKCs7adGf2q9Cihx2EJpv820P0jcPsq
jczjyQ7Kj8+7GznmIBGFpHQ9WDoFZXFNcu9lEbd+6KvhQf2E/cZXc1D+MEDscb+D
7de6yZ3sM+3J5FpaedqKdHSMH1Ci21MEhGUm6WVzx3clwWfQE2EuIamxgmGfMbsw
5gaEbiq9YObKFlPOH4ZDqD6FPU3D+CzUECu+sG0xI4oJvHge/9XZmOHyrb8nJ0U7
UUkoOg7hWvCIoa6ZFFU44NzY08ftaik3RWAgaCgzJ2ey+rL2xRxTGg6qg5uXvxYX
EvLuPPqOn7DRiAW+N2YXSSYPGw2xNCOPEQ//J9lGGAaY7gZ/x6hsbiDMt5cN5F/x
SU9j6tZL2vTd1l8T7Te+GeE9hW+oKu+r35rveFkvT9OkHRr9h35JVn8Hsya90N8d
uiX7hpJ0fElPt8hVQWO0+vCPbF3ZCWVBjMZQCc/pyh7x9Fh8DSL4Nx5NIfZVjX2P
5937qQZLQVBEPLFf4kKgbnphqbF1BBFPX/ZFMRpwcIolVMQhC7YOD2sj9hyumEdq
B4wni5bqtzo+rvWV37i0X+Hr4G74/UGtPcTPyizMNQgUw23w5ZWNmDerFVXkNBxO
2uWwIwdD4F5ZThRDLq9bCvgqe5OcQrgAYW5vpcsXiipSNGkYTkw39CST/9Vbae0a
woEd2ut2V/0utWctfzp4ZOlL/H8kiXvLwewfl+MH2LeacBi3FUTUr6br9yhbh0Cr
N/dVB2aQlklolySwM9erLD/CZbpIxNkfbT2IsK1kL521KpPSej25wexr+0+/VLcw
cYSf1GIoRkkk0cM7QscGYnveQEb86N0RXdHEmO9WfWjtGcl0jYssJ4qnEnSRpR8j
gqik2ezHirKjtJHqt9Fle8wys0QnFGHuVBJ/qv4hqZWN4SZi6TAWqeejjcWD2Bb6
EJLwy2JMYqmCEZODaFaZafdD6DgvHJoo7LAiV3Ivt6/PKzZMzudZm5v2dVtmeWwp
Ryp2sPuiKd1/o92Wiz+77nIWsdCgMWQZeuo1cREUAK4TgWNNI1ziFvcHyWKfChMJ
qoAtWzuiV/CySsu2XS052u3nNWMfy8bQeiusgyYUlDzwPjB8SH1fvUB7rw9IEoEb
E8X9w9zA2IBMbKOCPnNBKKUgsOBjhjQAdOeX6fZ+rinfLtU99P/k77oZBSNfM4pf
/047BwtJ2YhgkPTBHT8l78k1BckaUeACfn938L81D+MiYe/2o/0D7dqZoCWBsNgF
7bkp/GgGuzu7SmFLlIto+4Iej4/n6/+TdVTeatLWzr2PC+PTNsQwBW8xCcR+zLOo
AwNZemgf3tjX8NjOwTTxu+H5YMQhNz2N3Og3bltQqfNFucSknS+bO19qAK+DRieL
PnkLCLikntvqwLxvOZnaK6C7V7IwTX7cHa0XzHKY8r54Oa0LH5M0LZAEaIEU6KS8
jvRUaLl0PlZy8NoiMrvZL+iX9JZjAPUrA/rOWeTBRWx+PGHt/wyyr8q02rGe2JM8
YBGKeRMDRFPRcEhQB2/Kv9YwV0W2PHbl2PDh7u18kAdHEOPRu9wl0bdkNZCeqfa4
6opud9KQIqUgTg9kJjjCatQR/7IUutbWp9zKapdsWxzK9tc4o/Uixg833ISlbk9K
WK9OvlInHy/cU0NQk/wxYqqB+mp5M4kZaZJT0GL4w/aAIjtlvsGQVxEeCApsOfIl
3mOLg2YXKIwbyM/T8CLfc6TUUZQBfwmscsM6ZyQLfjR1btpS7h6htEFSdYorF9wT
Rg8kPeZiE3WBGgAqh+qf542TbCBYzc9j2xAT6FShJ1TBlCVwiei11Q/G7Ffl51KY
WWzjpnamtzbQ81pIjE0SkjVRPH8lB3Ci6g/yxD87uWxhj6aECgFGEFfmr/ngkPSz
mD7jjVUvpbqgBad+Ra4liaIkl4eole6orOnOc5EsVBN+qs08/HkuNLynrVdYn4ZJ
p4zGYWImFK80C9NEe3azpib7kf3hrHonHJ6Hc4G6hCaSsRhYfzQ4RoX+SJHMVABD
6KNm3oavdCI5UbG1xwe8uQcghPp3r+kh7NS1A/k0UQ5SSCTWem1P4Gramut/kiJZ
AGcd+gqw6DBNnIzysY6dVDE80ZiMKJn8BTqyMYKbO+hmQgWUC9I8GiBivafJHw3+
+6bCMUpJpr7VrLD/BIqVi9NYv7jz9lZsPAgf5lDM7Xn1VnpYponmLOSNV6NKlwkK
KObhixV5G2GBJmbREwcO0rNEz6jjrFJQhzm/NfARFiP9ffS/FXckc8rTluwHwgUw
1wf7ohOZ+XqJ/GEtYUecPLq/zuhKfYLxZCTrPO3izv5USgl3ymQC0FFpCtrdyqd4
snBTT4PrTB6syhI/LWx6GgYYfcusWzyEJEqcom9Er0R8NcensP/wfN8fPZLzK+ES
4G9QSqpu4cTLgiJAsrV3bIyxMXNQkRwl5aRTI/4yUYtVhZPnjCo9C92IXtPQaQVb
lRcJOSp8KE4EfX23FNej9Kl5cwm4o2+3xtOjPi2EBqnmdt2qON98f9ahIeiRErOc
9bQDuBAXxoOw9lhWjOjwuwuNtQc7cYbsX2xj24Sl5QAeIG6H2m9pCquVxY4wEhPz
OBsZJGLGZM5eUUEW9NbHN1PuSh8y6w57MjXaHGdKRNFu2taX3o1WJl/zb5Kb9gh4
ytZMxTIxK1hnW6/uyk0rDew6tD/TJGNm6uVS5f+srYHaW7Vb+oUii1oYavb1G1qx
qySpKWRgmg02Ap+34DcdeBEVyxDu8HaW3YXMMPtXGOdd+mBvAZYLqFt8bXyODyWt
2kQjvv92VoyzOMTFPi91MAwCLeozRWV2ONCOC7Soo6HmUoX9Sua4WkHbTz/Z5dZv
vnmu3gYpSqn34pEAcrhgGPoQSKtC5QnmYlzKO/SE0tCB/UXjeZ9Z1QljqDRrfU9F
VivVregC7R5MTysxx5hQVMnYLggPI+Qm+QPmprNBClSkKXWaGnA16pNPi+ncJzPZ
WQswD7YlTrw2JkMd8HK3siJG6Mq6m2hkSnEGDPhXvvVTwKsWDgbZ2vD7YEH/HbCh
JR9p4zTDunFSmUWawiQg5cRaWXSq5rqm6Xd5iUPaD1pBJQ4xA20phUUp+FG2/1OV
HTwtSuNXs00cU9h+Znx+T8LQVtiyicznOPV0pUuJuTvi6G3nLYi+IsOoJiABeLrp
Bbr4opEMpL8VFwvp4tRaF1COMItCnZS4AliNUZkQqsJkcP7xrGfiZ4kPADiNefSs
UGjRrfmVk9fekKVw8Ym9SJ26yUX+vVjs1pK4yiqF5aMeyZvyDIy9wjBerXZsF5bF
GmzAaFZ+/J8F7k5vcr1rNPmr/FrI6roX87dSUiWa65cgDenwLDbFL+W5SpZXRxzB
GAUyvWQXV8txX7GQ/L+2qnElM7223ePRzHhjyFLqOOT4ljWotL7U580cVmQe9YeU
IQfOAlF+vUovTil7ddTh5XGEiomAj2LmWqTdYZD9uuA2JFKl5TeDi2SmnG9ejud3
m95h0kWX3f9kTE4vNEnMCoaL7wr54oTnE6weWcUbotTtHXmPfnkEB6hybq6MypWV
Uewj19kyFjI8Zk73Li//WaggZxEZ3yjXXROEb5zdof4gPW69NhmO8gt8D1FcL8UE
qd7RrA6sSDWfoNxVsqW1uDgDQXGLoY/W56NVpM5iDLMx74U37ixT+/GZ3PuZlmIW
jBc3bviFcVujBvarJorAt/IwRSNjVMmPSG6+GAuloa0dsmzoll3u8+4fa9pgqMiA
MtBESJ3C5j68j2cNywHqxaRKWQob8zBtjrZGT5rn7jdEfbf5s2QddW+xjHK5Yc6P
VIaWTk/VXYjH1bLeMhgOu2+l5MpJWV9Vfx+VdMHG/raeQ6+/AJOrW28bdRKwP9TH
5uf2dYA55Q6bt4+zhUPhcYtiXHKDu1n7IzR0cGMRbkJU7mFwYjxzyLTSDkPn8ud4
pMhSSux85m9xstDwl0Q+crIYsLtFuggOdQKVh904vDy9uud7u27j4T73QKuIH4Tq
bTfRWvRhkzq3nhAxjv6XXsPzUyIBhIEAIbk4kRqtSCeRt0/CrKFaNibTEp/7kGMX
5f8OFjuIdjslqiO8Xyo9FIS18PgSaMujcPzdULlVhlrGm8BorhlhhgLFtaFwYeXE
O1Ij5KEbvdzJGYnkZzkQmChJlihPk9yWgxfJozE6qXqEj5W/zx1kA02z492NE6Z3
zbRbI1ZzizojzLhxsbh1+nJC78WXbZP+AkEHlTC+0ZPifZLYdlzyNDMAEGA/XEW5
yMvV6hntQQMJjw/voFAd1GQCHzPIO2XtXRdiLNs6WqexZ43SHheF3fSImJiVQEfP
bvlpAX8QwkCD/lHDiKeiUEt9cguFMd0PYDQQkhdZic93EW8g71TckiNNnico2siz
aqU49x5nuGUc5lFDRyU66z45KzLp8F9r5p7/sPwjrGxjvf1yvh2fVMXUcFe+L4RH
J8Nj6oSbJTAf7uce5L9x829SJ8D00RF4VqcWpsBxieauNlEgaU1iNhwI51EV2RK2
nNO+zvbcNGrsERgBZDmfl5vAH/c4OlxFq/wXwM2eW0i2xBAraiH3R5HXQmgVN4sI
VQGK89olOLgwuO3pvoS79e8u9l0KDQ+AK+xr9TN0DmjWvmUMDujGmSAMyNqWdW+x
jNboYdwEyq6wypncLS+YGPlbmhBqCI6gSnbTYkTjsLaaStPanypycmXuvOYb603U
YAUGcQL9Xl/syhnvkQ04IhD9KiEJAAIUja9eiNLFHaMgoCH9DZcZfQCtoNv+Td2y
3FDJ4evMIMWC7d0CbEM3iHD2BsTVyhp3HtK7bqkHzSUfvF7wYr4AB8wzkH91eDHq
3ZUSNpDct8BU9J3ju2IcoWkk2/OotRmwi0tvH/hKWRKTdIvYgd7NdeBYK5a4uRX5
/1b/pOfFF0X+ox7fwhn2WYXkjddTHBb/Zj2V4vMv2+HOX8lQWXmbkfk0MxVguHJs
PTiP53gSe0st6av6KkhP5wOKT68or/zJWDkcvQEt3mpGCVN2MKaLJK4zf5KzLdDT
aDYcOuXOFOyhtIXbX0CT+L7/FNei4wi0IBnDFaO8qAqRAoYZP93i1j8I57D2sywq
Ys3vQOv8ks8y8JlDo/vC2OtoNICt65r0KmJT86A9F9ETT2SdQKBPv+8SPp5kOXp8
prsj+uPUHgdgaWszAfQcaQB6QMCtzfcEum+M9Lc+U2REevcZiTV/uZ2+h8E9T1rY
FV7jU4XS9ki12et6KscRFIYvEfjqOeJpncZi9HweANAZmAC86uqv7/a3LNg8mH7H
ktytBphsnqaKxWK2NTZz1egGYmNvBFwvLUZCZ1mdWxKdbmtL7LMcsmcFuvmhoCGp
FDm8n+B8QEN5LKhTRAcbWHcF4eYjcMB4LI1GhntvUlAG4Q47uuFhw+3HWMWUmkSr
NC8DHgh/6oYCpfdyLEOVeerOUmtx/V09lGj/NFlQ7qUm3huLeNp/IlTy4GTxJgfR
YFAUl3wyNc4C2BJny27ZNgEKTVY4JIWwrm7jHYzLwVGB6/ycJ4EOpv47Eq4W894m
7x9BxOeggMC7pwgZx32Sf7MPGr5cxQnq+0laizIBmNYjn9tQ1fNB25+DgUEJ1CE8
fhY1ZeTty8G5nGBp0Z5dxykbNQ/XP5RrzmPUkvJOtjAFfh8uajgmxD43YWqwC/jd
b8FV9D+G7ENcUOER3LQ4WxOvWN5PG6USAuhHzZ9PNn665D9qMFH1dHHPPGahYB+I
duHnEXFR1VVVtB5Vl1ihQEsRQXcCbVcwydcxfC4IWfwuWWCFYwsSQrWfYVD2ivOl
BAaiEiGMJ7aGS9pssMipfsaG5fSqEUfJRhBj4eAZhbMRjn6h0knCKK56pIDe273l
uBSsoyqFqhv4rTSkZ3j9tU61o+mUepLFxsRHfWrFEeAHmxCqcy+7h44u2p48UR07
wGyk7CPXjeOf7e88BsVyK1UvnNIJlCzSkoTXgrhV20JxDpl4D0xFUpaDGfW2KYZD
HSSguhKa1SEI1HZqpekuHWeirdx/hAvL91rjCxUU71+5nR1hLSypngfVpAiUDPX0
GRoVE5Yx90bhLne2yEf9Bnsa590sGxTgicM2u3kCR9EJbOQWfiYvEzIATEdSVqcw
tHu9H6QyzQwstjewzaHhSnC7HOIjFJMTht6JgZnKGSislvYRRWW3hQRr6Umj1/xU
2DIWsH9h2gEP7F3xDa2CGiFjsdqrmqgBvkLhfQcvvjhi0lbo5trAWrVX0aAPGW+M
grZvEnhV0uvHpUlxw0i0YgWy5EESXgEMN7XyqObyhfGR7+KAJMEFpialIwW72KMF
GAK80FQyZShLhL1hTiSWYbRZIf+Anispkeh9gAa2NN5Twqh76RP7IJiu2wFEDAr5
V+WYwjKPwtRrfZNDY2W62b8p3MHUbA4E9W08oyE/m/i0TV2332c+4HgDqHx4pyiN
D8cC/hVxy5nE0k4zHAFL/lRztO5/W8ORVVqseW5h6dFRny6fwQa0YLJEhLjh15QP
ocIb6rD5Z0vcIDgejH+xqpu8FFXSxO8eYh2tVDe0cxA/OwZy0kJ1ZgjzGcHRzEw8
3aiy0dAcQmV/C4bxIimwcaFd9ioQgHq47HuTkrZEQX1TrQqORaum3Fp7RT16A5X6
YBq81QYTg3qTy9HBQRgdNCwA5RHRcfC756ib2qPtwJdbklW0wAdW1MOEZv2eV2yV
IknBnQbJ4vQdPF/XtWiUlH748ne/ggVC0oSlZU91cmJe2TiIvunQp4CY+XsY2Si1
4a1fq6QSAdLwU3YIxVVtBeUpRq4rHRSsMw/kVCbVU3TgMrJnQhebQD53gx6qPHLd
gObx5/l/yB0Zj767Uy0x/aBaX5CEm/z6LOBJtMa02l04u3DWJW0OPvfG2vd+99Wk
KaHy1Ng5gat6C0qR+d7wrCIiNoES2hwfSrSJug2+HOYJ/SoFkNzvkEk03wBc6KG1
61LU7vU/hjc88StzY9Uv8x8lxX13w7SW+i9TeYGzX99yRWRnPqvsD3+gFK0iNeiF
cIC3vTyrkSZUlZ4C1o92upuh6DCwo+MWs0W8QeG/A3t8VUK59TKMOTxVIaAz3QvC
IujGqdZOOiGPiEG+kkx4SUMYwCB+5F+A4X2nyV43xgpiqv6FJaw7/97MP2J9un9g
v+8qyY3VXdgkaGn0TZskUDXstTUJ21rj6jLAuid8pDVrWAq6zyRp0dA+2GaZMBKP
6Nw/ACrMBdTwy4zerOTsPjjMAfyTVxpMg1gDA/NBxTkbwiGX2BpF2eBcQQIkRwl3
1QxtC0qWAUYGpTBOn1vz1WjT0qbTWPXTVLjvmGrcxmug+jDrBcR4MbUBGPUUVWD5
lYZi/oXpie9h9UAJUA2e2btJJl4IjmF8I6j7AyHnBLdTnxGqUdMeG4yvRH+lg+Tc
tJ6ADFbXzv9KD2W21vPKBvKb7FJ6INWWTw2Xb/uuom7srKcirxpqSiNhSsQONFhz
RVQEZ3pyN55kNmnwE0fjriKt8JSAcSthFpGnhLjS917iRKsDmcT0uJtQudRwQ6H8
YdlSFzN2I7GWmXIov7kn2Mde7SbCzAKRH/OactVBIgmfb6RIoqEfNyjFF0m42kt1
P601nmLXGIBynFwtvsSnrwOXnryLs+WAivcvCKh43Lj8JSwsC88wlNzlscvH1K1n
Nk/gWqa5Yg9rD3BUdi9hOS/W2T0QIBK2aemBeCK8bd8UeGEqYCGZ0KQFpATjx1SN
6uDAVG4ZYP6oVvBX8qYEHIX8lR+GCYbl4C+cL8y4ln0sX60gaJkllSP8+gU9OX3j
M2ox9lRZ/JiYUJk5qKOaGxKEqJ9k17xM87SFWtyNJyAMiPfWuJTF9jiEDWwTMjyk
prJtFAxaGl/tvHNRakbBpfsCNcUbJhv+tbqV2kMhhQMK0QzTGozrFsnc7YtY6yPX
N13jbNuNbPfhUdJA6bxuZj/vI0Lc3GlmOqx0TUDzsCRPxXcgJmN4c5j+L6v+0+Ih
z0F49JX/mUAmt5giRU+r9BCOlM8CtbDc22VU83cHBg8OMsfCwqVnrsT2jHZBP1h2
MI7QoHOrq8BHqQqq6nqqG8XEsWsGYNW2FMxbbo/cKaB7hfWRevWKrzQaCQp/PRKo
YNx5P28zd8Oi18ggdx5shDIlAIpqZasP1Z1E6u6U0mvCgn9CLU6SInh3aSudcQXN
MVRfsbhNMr8KGIw9/oCbIukCsimUHkzRpW0AWqkdm32EDrZaBZcUwCTv9c9mreF8
WFDIjtZ8j/2ILEWWXtRD0MJ0sgWyWnYEom0CClwUnoWLF4G0xlxM4TikFsfxNseR
/kOy46aeXxUWF5KHCK7ef06n/5qJIKMR711vGy7Vo+jbneypZ5mJYGgRbtQmh4hg
ZqFBQB5BBLAQQvyOeA9QjtgGwOVwPo/GHiPH1qr6OFY/e3HZ+F25K5Lv/+MXPXRi
Ri/HWlfKAcOkfPoI318OYQNOfVyzmnwEVeGZdAW2Si/LFcZ8Z02Jn9TuHfQZFAHF
Lnm3AJoonmezoK6qxiwYiS/MPIOSAo0KznDHfSXA925ktczBNU8bhNwZ6KPXjQbm
oOw/nMr7KyS48WMK+WkLeG5M9cC0zRnFBMy8nYP5c9+mNwbtAaAspY582TdWfi/S
LfxYiBrEXAfbx9c4jq24jSSizf1SEsNZklXrimvOx/Pr2Mqp+OeFi69sE0rKB3I2
a02svVTJCE+HEPSYiPHr599zKJyKA65IdGqSrHVx3TL1zrv0yeEjWB/UOdncgHwC
T6504LaVvLKUoALAk/Jn49MibdGVwHgbRMst/FDf1ShialljwGCl2fhE4Q+665fy
/fPBzd4bobp1qu1APUlv9RMS5LSKYfrDLKZ5PPRzrwf7ziNU1k0yCzhsVf9hsIhY
JRymN8kNsSOvOP2UzTNQVybCP3QJIEtRbN8vU0oUjV8tOZMA//I74v+RndYaGK4R
SziXT8rfXxb0Z82R8/kglAZlvtcy1JwE5oZioJb1UDMezagen4djCsdiWgWX9pyq
OJTO7Wzu/RRh2KPTix5ZT9EYnv57AKVcVJ4J0iLSzFvCJnekdwpIfLT/5L0T/8gf
26eft721sYHGZOwdnfzuPuRwTQmaz9eLUoep/UCZIy4ZkLD9H8t06sHQCvvWM4yY
Obsd81Y9dv40KCIeDA6vQg+VNmGGBSZJTuqF3vdS4WFxudKo5Ig0Ck9yCdLSR3UH
2rMosL1bWdePy+dJb/BcQozxeO6WgB09KxhIEjLeJyp2zMht7GG0wUQbgfV1NAtI
+GVtPm2DvZU28LAMUkLFSn28mJ8Fm5E+zVyclLqtNZYfRzTPyw7sV2moavrLARWF
oAx4cXkHgyJvHwJLZM/FzIY50sPSUqPZ6qbafMhGdavGXYSx6//XBa+tk7zp0kq5
A62WblsW8WKp9vPjI83Bnw/X6YJ/4HVcANl3wu4PaDjZ/Z6fS8JooquCWlRF+Sk4
X+sELRPLmN3Lrn3pTJw8cHr+blWJifCsIPxOmtwp+MS5gw1z3Yie3vgSPYzOBHtM
v5axjdHBVYr7dFmNyTf3MMB3ajV6UNn0o/nSR92RVtQOV7yh69Pl0IAFqylH61TA
8q7+Sb1wHF5Z2K8ZaiJFvtBPElyv2D6JAZFsujz63Rihwoz2finM0UAlYzmBWoJe
sadoMKNEqseTsSx8B5qg+8PfH2NKR1Ox8HO678PI8nxZBLEfRZfTOJY+Xzyr0oWR
o88C4XmYj7tgURWi20MRrcdXSmGaLlIAcOUsTExgrOIMKKq9I7T8oIZSPaZwu3ak
eqbY+nqyhkuFGNImpjsDKsir0hYrgDKFO7IrmDjaMwRzrQcTE4VxKcd3aZrpNseh
dvsafqIUV5+psb8HDH2v1Sm6d0vnWtou81qhCdlGqhjlL6aikAAJqjmZo6L0D5Zp
uNu1jwNes40XZdqL6Bq8pTIJvDpblPZX8eP+BVkIU3VofXNUZbEzpPTe1v1SyQes
+ob9WAtdIcAselKwJ9OtDcKnKOLHA3lJKtLhP4CuGxWsowckmVndK66xwOdYuBgn
2sIVGxb2UFbp0YFSGUCPDoizigCjeXbVDTjqOfoDA69cc38BD8Cd/cnrhJP06UBZ
LZucG1DQd3dzgo5lCjNobuAf0/VxzLXWXj+maesqe5WewTaP8vPGYIyCXO8Ju4Yi
1ftRtkG0IE/xKRQ/Bnlx/VhqJVeWGScBGhDgYgbm13TlC++KuWdp1sogaKMrvyWF
QygY5HTLm5TBQpveXlsTIBhPHYRzfM3xO+jLEfrOm9GPjHLvE5iGh6DRIz7n2+P9
i4R7XOf2Cl2SXdoEk4zzV4CJ5wB3DQGyaJ3Gfme0QCZ2JU1EfMwjfBG4pOxPtfF4
f+M+ACqJGwVvzAUuEPDZbngrxqFfHaC4sr+QvcL1UTWpCMQ9OyM5LoeQucaOaRf1
9P3UsyKAq70k20pI+8SgXF+hTWTopUehCSK4EDdNRn3TxTE6e8OoURzEA1V9ERTp
geAfm67W9cSZNX+GXrf7bobl9m5HT8ZdokVXTYixXsnMYTp1sfofa28hmo5iY8wH
CuK2wHV3ezdKr/3SmKaQREHoU2mkPuGo4GlD09QNCYlbpezh+pHzyhUWMR7NZfam
WUzGDOOPqxHyrDvm2WteWGvFeyKXAykJNet88qB5Ylk2vhLZpPfp4wXUUdGU7jPR
PsDRl0QqxhT+va8IX0p0Z/TJsa/H0ePCLABHK71Fzjnxgd6cs0HpU/1XazJH5eem
AQp9R3jZS220GweUVW5kAJdBQgvxtrbs3x1wNPOaHda5bBYk1Y6YA6XMgDAMTRoF
xHwr93tNwGvsM4eO2rYNz5Hsd46svYKqcAgbXaC/QkNJheBdb4qEOU8hPH9hqQAq
tpruox80Tpso0O1dUgvywR2vW8Q+hLXlxU5YpJ+4Dx+MPDAbCwe6+p4PiOwcCAVU
2qT/AQImXlpmTcLL9aIve/d5SzkCklVzebPsqgbuEGyokuxo97tmHzg1Y3ibPuYw
7OvYs4c4kh8r9OMUd6vKVh27PV5wFa+qYLylA/G3B4iQMgk2mPveNm7y/SDjVDFJ
KjTDntVLBsXB09skjHcIG3qwbRni/a7pE81oG9KRiZ40mbcmZl6oU8Y4DZDZWm2h
GGoUlBcRj1rsryn+4HfNmE1IGMsIJIR9zGFsOpDfjdt4LUJHsOG0RoPu7/jvj8mX
ifGgYsHCue39IBb3yyyX5qcmxqYQPEQcUY/cylNxHIhz6LJgOwrU4UWCVBVFi/qT
8HTDHm3nyBHQEm6h16oASaiHI1UjvfmJKumpJiaA+Nh1pOh5UPTza0lzC9IblYzK
G96K821qWsxxkLoJCaAefSsa59yB4/J3Oi8GMyE9Ez2fSQp1lLzkRtQ39ce3Q2kr
P7PpVzynaXmBi20+JjxLdsfGF8QtqnzJsV3ggmKwi/RTWdWSZQfJOW160lkojtPP
nhbbqXHmU1C+FgeXT1BkHifiQQ5jC+XGjXzXgSMkgsllNVHGvDQvZ5DiRVHAeeR0
wSwb8G9Mf4vVrXDWGlOhw/yidfPFvEr+KQ0itJzKHc+OewR2fdkbRtRYxDpBMXky
gFEMcb/P++e2b5IuIHKdunwNHq3MGMoTJ9IK0SHSkD3Ijd2AvwJjbM03aVFBdYzS
w5+dU53yaRZHmK5kmOClBoSeNe762GJK6Wq7qj2FYle9hTvCFCeYdeVYYyBEQWtk
JQ3lGLSAulDmw1NkrN9O0VmaFxhcYgGy/OrUtb50mZkDOvus5OIMBg5mlYWedoKc
tnSZvc/CahwOc/hXARm12THezDKvox4TGaiEZ/m0abBxWK7vDOWSCtuyfnbzhOuL
Aqbn+rQH/rNcXnFtkhDKMclaVpEO2ZtNB/6EeIHL3DQHUsgSVw+1RO1vh28+zJIM
yG/5MzGVE+1oam8hOhLjV9YNYTTOxRVP1qgonStZh6dUOUwYLhpvrQ+nCVjx2e2I
ND0fNctiQxrzKR2S1sozisSMOqmdgfVGyOPVotTwb7xfrk5TLuRve2C8FuvJt6CC
fjYUoXq6E5bz8P5mtSwSsFF42/qbArUWreTvpLlw+4RPOmBmlb+j2jJKz9BoFPgG
SRGbgm7N81TQqZ62PCl0k19mO/sw5jfLqic2p5dYkQ/n8AvvNt67rF4DfgFSTq6S
OntkQ4Cx6uhj1hQOwBrO4OaxaKKjn8iiVYjG/lvM1eu02kuqgbIRDlLFfpulLaif
6x8cnVJh2BFh47taBvbzwsvcuUZOVt36POj+AzdcRsbVJEubYPvpuwnwmBR+rx0p
+hfW2Sx7w9JhOpOTzzdH/W1XQy1cd9mQqQYEPoexoTV/0cV4ZzsRbxBjRFMx25At
bsoIYdZoUI7xClZTmf6hE0NRk3LkG2zEyaZL7wGJdm3JD/zN5M6GRz4vjXRVLamp
u1VAxcZEKcJ8KiehtQ/aurjJ3mZBwB9r8Gu90S28tO9Ok4nTmHe7KTnCZzM4U6aa
5KQbYx3cJh2ArYcjmchc/NcpmR58NjJVHIdxwKMI2k0bigFbl51LwZ23CpbCA6dB
V+znzg8zP92BLuuNg9zu6EvgvxsoNyVlAuHDmcGX5dulW8T0wIWjn6uCd2XfsyYN
TIdDt9EaquhIGbrFBBgQpPnl1fZcas4DNxr7iyLcuoBmzFTC5vebB+B3Quz2MK4H
VGOkwSxYU/NFL21A6ii9GGU2knjlOVEkY69r04WrtTeKt7hjuknVQt5RPDrbyoqL
CNVNBbGydCa9Xv4zTyfEFMV7GotOJzmyPdlylFqeZUaYv1oOWKR6kugNnoxRgIRK
CRjSeEmO/yP2eaVvGowG6Hp87fkdqEWeEayPFIde7QZo42/5nllcCCDvg1SyGvrO
XQzneOD4EYGx9T3kDjADGNQOgiPB22hkgPPyh7ok2snHqk8FbqX0KtVrS2q7QOmE
G4HKhlqkzL3habYGhjqPertIXU08egdh7gic2+1P4UOHnjPFrRiQl8GVOJk8SXYO
+/bO7EINMLTlrm7RROQij8qBhJ+8jEsBdwSU2kUdc+BFl8ABAAkoMm+hkMQmVnVy
BsAE8hRIbMFdWoXMqXtE/tPWT4XwX6EQYtQ/79DPnBGUd4VpyNwkd0OrzoIFiwFA
YA53q5TEUTJwPQbamJW9ug3aHzntd8A2PN1tBtHJbhUng9a1RMnGJ3Bjc0R6Ph0z
84Y39T+0lJ+tV6V0K9vdUDHSJwrp39qLXYTpSj+V3nbcbOqjdUKszyBh9q/RwHpU
+XjBOF9foVq889saKWHU5L/XHvmSbCLPABTUBnA0/quYx9vlhhMZLt9QSHET+5Ey
NBHO4pmb3nSzPxT7KJxLftL4CkOLrri/2/DDPd+7RAz4UG3Q9/X5NeLSMJGzrNp2
rv+E+rPkhXUx2+bOeCTNKZaNOvM58x/+FWP0geWdTZuw+fj7gU5zfOl4I2DdDe7q
VnWTnoe9eLMg6Yq+8qOyNI6Hgur8FlWL6z5KW7AxW/lOhMEf9ur6IPhoN5yFVzJ+
mLIv52UyY54vEOYifczbBUdfNcAdnZhFY7zT/Zq1DxpQsOANR1m7pkAWtlanZDIC
k/jpEc0fTDB02NvWqjE7a6OwhXA7bHOSeXQDlTsg35pIJq8O6lcTSIg+C6XSgGum
uAWtYUjVV0qhxs4Zwian+effPkYu86PgbQgAb44yxXd+qnYEvOl4X+lGUJLCNgod
P4PRdxwbFLjz/BS3IE8uI9IYnULy/HJxWniLs9my57oWp7clxN35dLor4XKzYZeC
E+87aBwY2trDEXWHPylVGA0H24iEX67ZV+hfj6fa9yU1PTALeQrI9ymmTC7CeNx2
q7A1HZXyzt/hOvGBRKGKCUlBl6mE7WsguQ/efpI7fzyPvJOYJkPMorLzKUQFrSLO
vv3iEI06ON131j/rtDIzmShMB2w/W/KX6co3xaW8Z26fpcgMKwh9RzOv5gxDZO4W
ckVj6O6c9CuBhomHhS80LFXpmXZSLlqeMFGvypa39KC0g2YHT/2SqIl6EWDJPxGb
bUHdjnObV3bCtsNtRDirPuv3MkoXJ+xV63DuFwpjjhXZ9FHjuAsfAVrzHG6ElJLO
9OJNmHjovGwfiP6MHDp6syqj6xpiUgab9jZO4pqTL70lQ9wPsNTIKqQ9FdcTjRYh
pTk2nOF+Irzjd59kKP8qd5+WKwd6kPSJQYtHXbmfLoMkpIF73J8e7IHIIBiMZ91g
wXbHsxlEav+H+8/EpoAYKhs8CUX4l8ZaDYIEF7BaPnGTDsz8J3eTpH8qT/rCV4rv
7x7rsf69Qu4RALTKMlKDa5yuWTfu0tr2wKF04K2sDPr76YllJAz1UDjYNCT9PYbg
TMCMar+us6BolxBDFRHYRD418GIUNkjOOmNB7SytVTEeIT6MGAaZ3fUXHF90GQF8
I1K4FeIRPxl4T5fUKrkVV9jnYskx/g0e0jy/z96uGSIequK1y8h/1/nE9hMy5q8w
fTcWdI0mNVHZYZ40CrqnHbG8LKn9OZmOrn2YYDppbI5xrQxNHjm/nOCPvRZbeQ6D
lbA6WUvbpwDRtupyHd2+OPLIdt0u2zCYxD2125U7ZF5+DZRKV4Rba0IoXalVR/L6
jGuk4tgJ7Ttm6q1n2RP0p0tvWGtCruB2GG6Sj017FR5GIOJTmSwuviyNJqUJyurt
XcJeftvj80Be+vpxi1Xf2fR2N0VZZLEwz4wP2OYB4b/rMOQRU4zg7j9m7CSUGedi
EpviF/CxaPhdbRlFYm75gH56dCBHwiwsUSICrimbVC6YGTyhxWZg2GlOO5/kk9bo
cc1vOh2xCOvEhc6jwaGVmmxJuuWqPwhNGPnzBq4H4gs2/ikksP10DcN3BpnKyvrw
TGzXIBbaRjxCOSyS61GAH4SxIFO2RxXcUTlIMShLnQGVCzI9twvMy9vTVkwMYjVp
xBa3qlBXAD5fT1RxH5vNIN7EZAVnmUbW2fU+OgH58SgONTh+b9qepYRu0WdG62M3
QJx/y51hHkDg6r93KclkTJGvYDQil6tGFuoXwsOCB7Y5U+dmPQHq1jneexqTlbrJ
KnQ0meuk1FAjrisKO3Z7twyM1+mQZNjnBnNfy4NXIga3qM0+ElwyJeXirWN8Qyta
5nK0+VN9aY2n289m86KPHV5WVDvxjOgpV9h3UFPXKFqZZj/7iLldNXi5IwXis2Q4
7H6QCpKlWeFa81KsV+XgbGSmr80DJMOEYiiVSqfnaN1wglwm8CBOicEiO7c+Lif/
yvsB9cseO/yD3Z+20nKKaQZYeXMjr1ysnxk7Ww14cwaqFjKMb86IQeNReKi7u7rz
Tycs+YtGWhnOiyRtFp/W85L/ak2ls35eZ5eX82+Wwzwl2iGw5451/riiXVxpZtC3
9IzvWpWNa6KbQANKzf03gR8eRoAG275+1oEDyZmRbwsEnvTRd+6lPrqRZ59p012z
9Y4Het8IRYAtAnThUpdp2goE/+zG7a7xIFdz/O9RHlV6cr+N6LdvpgbS2WNAWBWz
8xwaY7AEsR89xU+R5eHDHLdp4qUbWqilpVRSeyuxJN42qub3UH37Z3ZQOoaCZ7nL
eHGgL3sZQrgbsZIgW6wNcnn4S1GJZ/mLwc8solwO5QrobViFayKWAF45vsdtY8XR
3YWoZfxeM++B/TciB0gIEHNwNtSjxgHFzugv9o/psGtavndcJr6hwQ8pnNS13qGU
B5e6kH/+kbzrX8g0BBoyewIiN7KDZLD5HZBexD01dElqeg2BIX1/S90mvVAQ09jm
KD/GXQjniFhB9oDcPAXnbyS7pvgVXuKOj4W2LJ/dauerTX+Km8ZDOVdmta+fHtnx
RDSaVg1FFJ7pqoSHyMKRAyOyYPL9RYAH4KtMxEeJRUEnqyH+FdV5gwVyjE7w+4ze
ylMhm6VNxD6mOf2tDRUxoS8xOnfSF2JFrKbCXbnJ+JkqlM/9l+Y0AreyTZzTw1l1
vnpw8jdyxb+Opafbdvm2vaixWppQnWnA3DT0n8goFYgyLZ8bcxu7Lo5tLIAw39Fr
+fApORTCDgTbo7RvA4TIHEL4vc0oFROqIL2/ie6mYtYQIB6uODoHJrhChdh4xtu1
vCjor/Iz1QsL4DsQtJrMDnBqqqCuWEnATZBXP05XyXlLfbwMqj+xEo+h63wuwbwu
SOz8XPLfBuKOp6lnxhWPkZ8QpHcSLkl6u5WnL058pwRZYe1zuRPnlWYtROCvtWJt
1H7czSqfOYvFoQC6KKmxqmXwC0ZgI6zrIOtrNIe/XxC5f1kUZTa9wXELvAifeTyH
wtxDQET3EOM3Vh8CNQz9U5KVswVCd6i7lNJ4gHgfxyr6wHNHdOI4OGw0d0PkFVnR
2BV784FvExeypG5T4Tf3hvLkLAYGQSyZ9mxGVn1WNpGTNEJ9BEloYtRRT/5Dciae
0Wb6rl3qx7Rbip0+bdO9qZb6vHgi2t90L8jp3tKC9HSib0HauLlJggWMsYcW1kck
aVzT4xn0iBdvbfgbq33frg7WjljVoAddxcmAu1WkvGDKL3E/25IsRQeG5WUb7+fD
fgScRuRHf3SG56bwZHLQ088eVt3x2q7qRs2r+U/c45Edm10AgLqQ11CVK1DWJfRv
YOk3LpNAzBNaVN4NxZTHSZMsXn1W3o/V4N1klIcm9cyLV784SMs59Kcj8nwN6Yby
wBC+h1ndruECfl9I/mKdYg2mISZixumVwCimV0/KwX24zn+5nRA1gTzy9BWmHlQV
vPgaEdR9YwBrf781FTIrV+CanWjGEPKxodNOGnpeIfV0ONp8JRcPM7mfOn93S6ff
qOb7vtKoy8MNBItWCZRl4gAlA343NaE3X+r+EVlUYskazNGdbV0zEF5ZSvtcrY7r
eJal3QQpWwZ1SJl1Vr9rOROlNmcWrYY3YAIYOibfEfkdrdUdu2iT6d6sXq5hqOot
PnpSQ+kD4fOPkwnFiVsuTyx94TrloO1WiisGx6I1pN8v/GkSgMMNyy80hv7crqI8
VajZqmQgEultPBm9YwMqgzCHL9j8vZeUQv2yT2/SFJULHoA2SWHKiHXFS+6CrIA2
veVhblVUB0apBZf9JkVGpXNN2e5Eo4AJDdRGPvmst8Paz4TMsMAj21Bb5kABMfjD
oGqNg0rg1r5GlFnbUmA+xuq6zIz9IOj8tLEVP5LKy+VDL6S2lur20/dvkhdEy6vZ
SFrxpu1F8zLqEbFP4y7A6juSo7X1pAeOdw8HMRobHyjC68jfn4G7xVZsalTATL1z
cOCNZCarSIauN45zhmkErMeVr1JRlxAqDaOiUU8VpU5QIpMaNoO5BPcmkIhUwwil
uclodotEgRQFPo1rY6B63N6d6dQ/h6prv9m5v1gHY8SQZUD+J2WqWYvfUBPy2Jag
dSNLGBy1wBPXwt9qoaWmUZcC2ZNTww6pEtF3dUP8bHQ8p+a/ipg/pIrfjFb8PRnf
TRySl06P9J6EkFaRUcz/Hb6E8eJz71hXJe4ILpQ7mgmARfTRZ73hxO8AeFzS2LGb
RM/JoAMK0Tb6PeC/BHW1iGqgKscXzs7NC1MLivO6g6UxigWnKCaTQkbencG6A3I2
j6uFD+1FNefKH6qLajVY8IQrf/fA+TBEAreez7KXxlzE5TGHEwzDY2RYaRsB9N6I
bzy/gitrwcFGscd1zbr5Udpn7DgX+BmJNZEzQoK9Tu8mkcqFk7HSfyYjkhhvHnQx
QES1o98aRsAHHe5d3vjbsqjWtwJzdlOZoGgYNPe8nAjrs3CRIWq467am6E4KCZPF
UV8U1tAmHw18UusW3eqdtM9AGKIWdQWPaKHGLgKJD0H5EXbtH5ZmTYPQhVnUqPKJ
xzYzPYkHnGsEzpflJLWBfvn85UINt6jdO4f9D56l5Zto3C7lFV3DfqH6o//gU6kG
LFVWwNzUsMTFazQ9hSNO6j2tzb1hK1VWycaUoQoSyNPGs9Z0qkG2iVAM90sNh2NU
dIhmAu90ea/NULCkB0vOVLkpFq7WgO/YU9gVjC+D1JveDBYZ5Fx7Uz4UZJdZ9UHY
cixP8z/zLhBplzbvZuFR//u3xqqhabs3mEIOMbW6LrD3MkdpRBY52ZbgVeg8ysv3
jiIOIPzJFi6J1TybdJ/zlEUxWsY6ZEi4ojgyItLyrNDJvH12OfmdvuZS98KFmdPK
108D9EUzDolTUPceBJB7lLuxFt9Z1N/m4gLY1HaxMgZIKE8bXH7GIUIpPqAmljbR
3bDn71Ss1/4mVaTJ/m9VeAgCyNQmGBhYmovZyjMlE1S+g/4HBFTaPef6lCtNu95l
/RKbDVdLcEzHiRnFN80lGdEEN1QGRDQWL0M6GhAD2QErbWMXGQjJoXjw2I4ysH5y
g96vkDUV45M7+m14GYrG6PsttsmuIW3uSjxDYBOSdN3IcGiiazUMmJHPEC2j+QIp
DTJl9cLpqZINXWj9+CW/dvFkTqcJvVh1/tGfRKMEx/d8tuKSwmlZFfTTdIHTOCDl
CU/0V5o9FnWvvYWnVPBds1InmzpFK5suTI8uUDw2QkBeX01GNszZkHK7A4YrYipI
EUJBOFoTSgyXHhjRJe58tnoSzsy44gcp/l9Vgl1eWanA4vvxaArT29fvku2DjBGH
82+g3hhyvljYqM8wZn/P9evzHVKkWyYOtKyAjwYhOVCr6PHy42Nyoz0oFFMyyuN6
jBOBOJNZG22e2ZlNLmG+xrZophVbSVN8UZNuM8ApKTmV79oOa38veBGaLGqkvtMI
3abudYnG2Hy4Xd9BffDrROOcwmeeYBRFEBaYZT/JOPnxXA+obpTsLwCccuE+EkHg
DDzq8EeUGsgb4PMC0mNty3/mkIbp1hwBDe+YF1/Nv9O+ng4SxotLsXZq4c8MpRUJ
Yr4uGdf37sEBr2Cq3Du5DMK1eyT5EWN/wkW4ugEz/7MytTPauZA+W6z60IR4aaaq
J7bu9K/fl09IEhu139WB9ixG2JMsy0Q/vh3u5vPaVX75/wAcWc752gsdOHt9z3T0
ZcHE066W5K/2tzCUoTagazdodRKjwddVv/00S4ctnx+6GgV4rkz8FvxgCOpBP0nm
bmf38kA3+wlY2rBo6s4pOLFt1khOYo8sjRNeHM0Tu+YqMNpHTmKzEuMAQ52p5+V4
uBqS7OtPzszruaEiMounxE4wV0CtdfUGkhKAI9eYNzx+XX/anmZt6vFRNTm4pric
x0U6LSzQnTDmx2Do6hDMTLMto9nwnrl4uy0a2RuW7LTnkNYyM51oQkrFMPCm9Y30
p3Vo/eHzOZtC2JD9NXoG2H6pAac/AEYduoZbG3U6QHH92CJDIvyC1I4Q4NS+wi4v
BoWRiCpiC5RmZB855JPWwwrmovtAWLJzURBTAkdEdTtm4lAc9OsBdCtZhht3UxqU
bTZSBL2stTFVK93LLAnUOrzBhfCdeP6r5Xdkl3s5PFBF94wG9Og1kkkz3ZuP5+pz
iU72fPWgUFReM85RKu+PZ5WN2wbeThHbPRexOlfhBcNlFXm9Aqv3bgsXYfb4dEv7
rdKwSfNsOkCcOq3osnuaILrw84pwt2ktpg5z5UzXlEAZlIUArztcSCI5LTim+azG
QvCxR4q6niZmI3j+4DlPwylOdRh3J+73krR2X2vhXYpbiLb0BJA1I1cCrmMwWNEi
M/ZssCiJVZUuyAHObz2E8VucqxpqNxAgbq7iybx/ppQAowrQxJ37akLVugAlNK5O
Op/HsfjGW3IM8vNYhC2BE5sPCTAsKrTaimX+lMUz023IL9GP2SpQMetWSQbUpDJL
kiezi2pnNIddav2jzk+3Mcs0dfifXkllqiLoQnoD3fRs5k2LLv5VXK37FkV60oNP
ZORM0NQUU0P1CRQ0kSo+fezIsfXWk/ZSFXYcdvZwQa5wUlO5oizvfPVt1WjBGW9E
0c3IPRy6JQa6hvAiQXx4JIgsplWsWZ1x+vdxSQWDm7aoRRuUz+oR9IAYywc+2D/h
Tn/1dNCk6nkc1IGaZEAVasychujBqN4xwqAREB3KfvbLHgwJ6Wa4yQGO3m9dBKjJ
AdPwXrFpwFDxD7Q/akT+gkbwrgTfP4aCkzX3FqRktydQEB9XmCkv5Je9R1ps3M7q
ySb0ZDwGNb1LohwN5ZNQSxLQno0RViyNeuL1gWrJ+98mV3JC5NORYB5TKH1uJsDN
bd6LBsqiUktLj6EEuRxjRIOH0qYQYUD7VsylyrznAtLfmNG81XmoyXrATwLaBB1E
5ZbwjRwB4Tlegxg8u5e8/urNDH7wvHOmm2kXt48fDRYl/OQJig7ENjgLfaqUxh32
KFcehK15tUwF18keSHOzA0xLd96UUtqIdcpSeomFCwCo72RfC0rcd8HmTjStUcZg
nhLsjIAxM/iR+j5nQ3BZWHd7tsE2D68HtVU/TL08V714cQFBDumGo9w3EcwdzBBm
mXEXrDBbkNWMMV4pKvUf85RGYnCY1f/Z3701Kun6y8I/UaWeAHK+Uf/0bjcWTCYw
CBX2BzGsM96/ABHna6sY4MZ6qK/+pBDVjQPfcky8t3YT4CXg2dsjzXWfsK93BTaA
stuJU4osxx5yqhvgYLHbKC9dWDKLkSV3etpaGqYrI44uS5vrNRdSJmbeNcY5rN8M
LtHlGP33j7QyfnEw5FUqOQyDLPROM/Tlj+xkwydI8MCLt0D9rSKIR8wGsdI5/JVP
miujnH8/MydQF08uNeAn8xnySsegmtcLWsiWlWBtx9SxMD1s3QjucaJrkQ9+Nm57
V0WB5TH+HTBTmHPOrH06D/opqKXT+UnQ8x30QdTOqKdmmadV3NSs4T1NbJeJKiNf
C1emlXBEawGEN12KajnctAlnigRc8rBAA1QAd34bjToNtKFCWyiGdyjZwoCLzvi4
glLO+xlT6S0bj4qJLAcd4QptgTYH6iWUys6HWnP52YDL9/OjtXYwNcE6VgEZZ//f
rrV3tBeZAhabM6CHoy1f5d1pUC6TBQ80d2koumZZHtaostO23waabp2Z2WBe11MJ
M9BVgaQGngmGqFnq1zQQb+pneyIIAw94pNinkyOkBw3HF+SStPSGMQe7NVwFLKCi
73pzfsJC/NMf4dsGbQKmcgWKn069ifi1NuFsULZFRtg/UMvBt5mtDWj8AM9FJFbs
0EcvIOAA5s4pxwI4GdmatfudKt4T5pJvQTAr8d3H+jT9b4O63BJZddaSzbI4z45s
TbariHlURrb2k0nq79b2G2FyHwQXqWddGb7vk0+GGAmL2Xof48DSxG2UWJsPyaML
csQeSGWzDXo5Or7dlCML7rWsbjmXywU0rXnt/Joc9Uq2ZmNe5hDhROCvZSHGBqRh
BHdBHtYBw3ertCUFPPfosl7wpdyN6AsGciH0J0zbTBkL/iQKe1ajpv38IP1jTbAA
Z9C1ttHCfy6ovoVYxDLmV2IsqG/UsFa2loRdb98u0gp48M02Am9yqsWKp+6l5XG9
LhoQHd9//Ucdqap5NWk0HQHHY1Kc3hDsDvVvaWgdwxiNfO+150XGymNDNY8zQgDT
s3DrT4fJ9yBO0EeiwY8wXU0d/OxMZUX0fh9K335PsBNLBq3YtComrNE3Oj7bit0D
zKfDIqCPXe+4gztNuqi/qmJia34iwcctD05eCpoBbxky1RJvpf+ov/PGahHZ6+Lt
dt/7mVAexlgQwAOm6rXaqDM98z9revqhnKBDLrw5m54HnqMZnWmckD824yWXlm2k
UXrOEmMl0EM3ebPiY5sqCyTTuh8pdZTkgjau3zTsa+FuWf5S4jQwJ9ElpkA5pNjC
cePHvFYOHBNFlDomFjY5iWEahbReIH802ubxFR5q1bUgFXx1Nx2hpn2PwrEIQOCu
sLQZukoedKLquTByqR3ULSqwapf8jLoewWEQZyOohrC1j8OBvgifc2qxCHpbg4dQ
Yhz3X0yUyPFv560ZfY73CVEobfvRO71nrRepwYFrUy0DtZ216j737wSZQAxv8VE/
9OJ8AO+ZZpamyndwW+DvOy49z3zUz8y+b8Trxy9u4r/a5KC5mweiL0c5QuH4aSwL
YGmlTa5pODE3GS3iBPXKAckKJUcZYCDtGyUau9FDK+5JsglJrW/aXG8CUCGtaEkC
ucUD2xEnunnQ8a5NsF84wq+oyX2D6Ij4u1SCk+I2nCYqE7Yfv9Cq0heGMzeW7ttO
k4xLFtTXr+dnj10KAv9Dk8JIJ0InyWi1h+kAR2OSsMxON5JJkAUnrbiVa3IskiE1
GQPhRJcXNzka9vOpHUeTercBX5d+VPQuBcNeMTaQ0n8kJK+4Tp4nWhkU+e7vjbCX
yRd6OsCfqAAjsrPrDKwlzWB4vOkgZkkNiJ9OcP9ZxK2EsCCd++Clorf8X8g5ow93
biJToHwgsdLhidQ5e96tx7Bwsiu6p6urapV78aVpFc9yUaRoCDlPkZc7nD/0y01N
F0w9QFdkvN6xGMnuWBECBvYJVmzPFeUJXUfWY7KO6uIEnEEpujdsTaFS3P4tVYt6
rYH+loWTCs9KQMJK57jltdq4of2dS9exMpx9MRuv9QdJP1YKSWy+GEKLSZ2wvlrS
sTr+KEz0E1R9CUvpB8Y2/4b2KML4tGarZLL94fSQvNE65K30m9+kyYNCXVhjltkl
3BuKTa95Ki1qo3StMrriwBQqCb5rxh75CbY64+1TBlCmcrsFeRx9nklmGVmcoJTs
Ap/jgQ5KLpajraFWKcdHe6gq5SUEXFtkVR3yHBiOqj56PSNP+z6Jo9ze6WwIskYo
ttHVxctV/W0IDJT98q5+uZcurVnLDdM1qlsgBgXDDYtLZv17E4ACC/ogZqGi4hfC
A7lkXMJXno/MIay9mBXShdlvjr934rw0UqmzRSyb4XzLMg8hRm3pDml+U+Kg4O7I
NOJ72G1GC1zSKDMYf7Zuyw7ntGh132aBRjK5iA4eb0nto4TbAVhYpo3xK1XDFdYW
0hDqaR2rDZbQ6XE80Bxqcjd2BdamwMVGeL5L/kq7X4E6a6rBNXWGJRYO5OhFSlpF
/JOjt23L96fU/SkZrLJ83ECwBfMcZv2GsrezZZRujG3vU0I5gtMMG+jJEeVIYM5Z
B4TnREi3nltKgi97GWzvUwc+PbA3K35mjHU5zGnHxRAzlaYNom8qhryT6VZWKIfI
tztY4uqEIN5PyW/zmykwWkh8tq55/98xc3Q1Cm/Zrj48VKzebJcY9pqvEejw0JYU
dzXKmNzTF/FjDRdMNumjorKFjHyRf8qSxBqCcRkzTLI/f/DbkMGExFpww8pe9h1D
HcoebcwWXcQO1Tk2Y41asXevN9pcvMB889jgQihq4juLm/MwWlLfV6htJaB+1tGB
1IM882G+PLCQkGj7bkB7wYoqvYT5QnEaRanJnDbY8Kgu68v+NbWEH1si6WP1c5Wz
rbDwedXdi18oXyPFvY/HFDDSHpB47IeWbKv9467S+aniwVNncbhX2rTnyERi11jQ
rkxUD7smdplX/pubhI50wm56hiejY5B22F4WHezK2LIkYoKXLgG3kj+YHkZnk62+
1xL/Kw0KDWljyr54y2yjn5Aja4+DmmEnRxdUWZbosOzhErTQXXgoVjA9U5kUIx+9
eFPE2RnNfM58W5p0FFwANACFu4Iq9VE933XW7QDXr2srZZpR2I8Gpo25jDsyFf7I
WKrMSs+uW/IwUH6NdrdyDa7ksKJ9fJ8h5ZxW8Y4p6hZygThAFiSu7P3/rvb9YBzP
u3t3bu6edMBiA0CMaZfUfurU0dCRxlEDu66HDt6JlMPOA6fHjJYNE1XI/oriJMgn
rQmftHSbHkmD4L/R6x7aHI1rsAWO4wNx9MvM8DuBFyfwVNb0SImWmaZW97DD0yct
6bAyg9vCvuQASViP+op46Lis5afcIjnT7mycb5n3zm8rQ8oirSyMNEo5hy1ZEAEf
cXwb2/dIKYLZ477TYKaO9OrbyuMUkOqU7XfJUaoOzfWrDs1qYjV+9i5gqMB0crEc
6NjAQ+FJr0G8DWmOa/tkweDOig/fn98S2IOo0Q9NFjD/Mt8k0sJ3xq6BCbPOJMcJ
Zh75GT49Z2WGJ49Anq8NKaUIxu3QBeDZ2RpaVDgssEzGb1HStjhe/5OhuAQBpyLA
fDKRTKx8yKV44Pz4I0zrd40PIKLLWPH5/TaEJ8rNh5T+RLjhhUu4ebvmLvHsfcyB
aibMK/tMJH6BknNM6d5XkD0oCU1VIpNTpzC/lAPndugKv4EYCs6u1wcFbX95DQkG
a/xWLJFCi8GakqWnmhcsN9h2N4BcrtTHm/QHZRCsUYHlSFQ7s7wUMlotK0kIk5BS
QIx1d8AugxYq4HaLda09/EC8O84QYzGGKLu9iZ7Opv3w/+MyR06Huann2sitDP27
uYal+3TZ9wRojxKHm6i/cGqNNxj/YTpzldrZITo/6pRAwRjnNsD9imLzEO9GGSq9
XsnxITCYgh79EHgmiRHe4Q6m10fZ1CUfQG81qLnSLXfV/iMrH16J7CiBfMKgzXTp
AB13zto6sHyhMUyDApmYM0vO2Ldz/bpJcoRdT103eO8t0hTX1oCFPKyBKMlFcO1i
wKXOO+eiq+QrT56xZKn6ACeisc72D/H+8ZSqfPsSoF9CnoBy6BepJrQk8QMAtAMV
gCoRccNHD5tdwmogtKmEApoW7eiwPTTNf7xcxUWbExxyyEH/TGFrvaLFCInCCet0
9VTISNPK7Mm9J1oYAHaF6T2x0/JK6SHZNKPcg1uhZx12khRSJ5WZmxxQNDNNJhhU
WtmRL9EnsX3iMke8rGJ0OdpcJk8FD4f+o7+WGKVKLpM7XxWFcM9GfkpkftLJUZ8I
MpUprknFBE8OVXGrifmD4+KkVVpOtAmVT5sEGXqNYD3mxjEJ2/SrYLuggvmhD1PN
ekaMJvxMh3O8o7B0esPrnQ8wkg1RnWjiP3ppToC2iwcTGWBIBXBLWFZIk26vR2g+
xWFE7QWmXafkRhbrjLXJewpLGDRjZb3p0yo9N7czbKnX8kWmrVm/dcKX8RaLXRTm
rYk45eQ5sZPlafyxBq59ffgxdla3KIz75ED/3xdvKqTdII295MBVu7wrpEReeB/l
/o075DmXdm6ISUpAR6GlvPc7Uhhdxe8Hnu3AgvGmVEl9LnxEFWeAnTeu3NqHNyO0
2ZcBCj6yzGIl7OXEF6orVXsq0pQNe2mor3fSqJcmGTup6k8ZsbTIOZ8dYS+VCSTd
dlw3zTJiOAXZtL21Blq66wTPGyCKZnXN+aZy5qfCWWs0U4l6HWgyXNKsLchRgKcx
HmGatXkukLg2v7h3NGtz9Utn6t3oD2dWNJfaTvEAJB58r14ClarFqn0CLHsMBGRb
4lp1VvTuaxrJqgpWyRp9AWfBf2/MmYnIZNJMwLtr04jCr6wCJe1isR6aHMt0jSLQ
+V4gqRjLoiJznsxRrm8moYZRXhyHG1gWgKPW6zH2PtfPGq7BNHkLC6AxwBZIEvOa
uNNvzckk+1/AVu2e4dF4x+dEaMYyKrlRZrTcslOS/NgamQu/2ti4zIksvGOWEq5U
QrKAOfQNksEuA5PIq9sdA0Quqdvn0Ya7fBS33QyCyfUdfQa79KHJFRDHUDwenPFA
OinoFmzznCDm1W7U1urGPdCd9J29xOpNMC99N4dQqow5iUfOo0Dd7Lwz0eRnqGF6
BL2DAzPmb7y0o68sp0PG+UPrNGL9mlqW/zltG14RVosrqUn90RMvCAfL8fOSnIhD
OyNirQ4Z1S44pwYryCvOrm4stx1+rjhwlwp6vgfruhiXt0nuZehQmpJq8Kl37sC1
5KloCR0Su8c9o01WItLmXCKOIKNP35dZAolVIP+d8Bg7BiIV8/hAhOsueau1ow9C
ZuC9ZqB5lBZqdWZcXMOfHGjtUeJvw9E1y+3l74lU9ju2CNRrg5sQBKHCXMfvYXLN
USQqsDpFH7P0HQ2MHU2LU1SJnkBmGrVT2G182tx0TgrcVDGReVR7jxsohsEghfsn
vlYL5+4fOSK25SZr1Xs/+EloerUwIGYjYVCajFHTY7uXbuLpLftnIfvOGJZz02t3
JLqIg48IaxzzDqePHTuBgkUvqG0hcZxv8k8XZNtVBJv7BfXCynU/PV8NYsxxYX3E
Pm+fBKYkKeiDQ0q8jwtusMRiru8+RS1nikzrMbRIEOefplfwb8sw/3SpVGk/pY5i
0fjREkwyXPiPhlDybkBHHZgU/yRdHXfm4R4hz7bXxnc2Hwv7UW7i/DGeAo7Y/efB
hymVfOTBrpWCiTYCBRhY5IxVpOD8+Vmx/yxb3/DLp7cjbzM5HaRueGA1dJ4P6QLJ
FsH5FZAiAN77foyx0ENRv84z8N+KSqT/IzIqf+bg7jGaDzqLyn81N6Tft3ALlApT
CbWcuwfnSFq5UJZ04V3Pvfn7Gxg6YHW2eqPg6xk14shMGMNxLFrrmxAw9LzNxJMf
KhyLbKLkp55OBCXqTKunS/u4PX9wKxts0tEunCghHHzblewy6VllZyB2zviWPHsr
BgXTrZRbfYEHGW/vpciTyGXuE86tDyQy1cxaiUqYjCLC2TuFkgnh0RfCqbSDOsfP
uUNlwx85sBNzmYlUcWmjFRrltHHElbxHknV+CJFMqylOR+w/U4zcOJCyFcV0FMxS
mcBSgFYxkmj6qB/WoGwKfNK3gbiZ75pAcnPy6REVqCHEAfTcVzqv7Cnaz6Obxubm
+uvMG16yHtqNiarhgXrbmt2PsTLoGn8AowQeAiRdcXPV1/rsAdPBnwQN1CE5vAd3
Y8vDoLsPI8TfLvvzocRW2D+eZBHb5tNzUOTRm2UjZS6342O6TZpyCrHmmw1luLdp
qU+FnUuoBO1mfAbBDNOuyPSbj/4fzeodA5okP8oNGmqup8oEau+Lxil1QM2ky1n7
R1x2ybcj/CuY4vfXg2+77FuMaj04ZjfvQQDPs+zegiKfBTHYne40n4LOxBVAoPK3
ER4C5yPmvOzMXsqjRp2gRu3nhPPeE72nNWg+PxQgxBHcYDMNhPYAJhczUxfmzytb
3rdqjV/ZP/Ut7nWutkNMq5n2/cm/4jyQomb8xGPgu4gVQhEhArwB5xdKAFJb+z9x
2BlOfDxXAszmQi0jCIKHvVJIxXiN6rpNsjjzNRom54G5q+fhhV36s4rXyLhXtKkE
bqXvCfaov11ythyHaFumyN4sNtlCrx0qFbBINrPZhcajmG9YNlPeU8/M5fmfocyJ
PeJqD12MAcGGCeQl1RXIadYfEc7FJLp+r3GePU8SNyE9amlJb3A/SuIsIdAqQkup
H2Kfdei0tbvyzmq+kIDLl2U7Lj7XU6SoTagdbsOXpFnYjP6ilK5HzOOARdbjmNiD
AGhSZ4a9pXOf5E4TRZTGqQYekuvexR5ZqrMjwsNbj7aEFSrgBBeMTpUAQFaRKJhS
ZcQjMsSIjUFoOkM6OOJb1A9KhVNybaQjs574cWdTGgbTQt0jYNpoVkjbwZDoF+lU
itYtfQb0oy/i6ESx7rVHdQjgE9OeQAc6cQ+HKz50T6Uqw/vDRDiSz6757vV/QZbR
HyO+y99FRmAnuZIm46kuy2Phig1GieS4l3LwRO0oZZhUypA42PEaQ5rEAF8XaGjg
NFK3BD7XGwE098fYJx4kVWd0MRzS5vUyChEtUKejBDvt/jV4zhCgUq5K+3zBbYWo
vjXmFmOBbw7YrXhJa6BO1QFWmviy452FnLYxyEcpxu6qDQV4BAo2Zn1PSCparmqg
QpX3o+aEoK8Th8lsb03vMFpvJG/FBhVLlseNzsQEjtgg9QBbjkyAtAFR1fIX4vVm
wTDqQL6CcRFcPyq94I/ml4p3WNAMOhe3tPPy+t+soFmMw5a4zDuuEniT9u9OtM9K
DqhxrdCOB6vEcUtpo+bsruO1AlSFtE/cjW2Yq3xb/6skAFjx28B5A7utwH0+IEcy
mUPe4P8xgRWbwXqa+D8FRLI6EQfjarU3A8DEVr4RP/W4lhprxmy/PD5267Bp8c8y
8uibv3GeE8sf5Rim1M3gTW6WXycBRGH85f1I/8la+d7L4b5K0bOiyesp48KqsG3H
2UTnGD34q7yjY5Lah+aTfpI1GCIbodaRyF1iT8ZWdwiUg30JvSIPwVWHZozYvkdQ
HGKxVz5Q45w9HtKdBUi1O/1ChS0MkNw2gYtB3f/9wqBqSC5NO/qm+OzyZcJ4WyFf
bRUc+voWtfcnAfpODecZnwKZwqhRci1jWm8Jmx95svVhFcMRb6HB6tDeLKCPWV7S
gXX5gPZH9ehQ9ToVATdYWm0/RLmrCp+FVUMSc3KIUYQ460oAPkikWbgBnQGxVMXG
wWY+J6qB2GVrsl3eXs5jbB9BpaQ2Mhcn9Q7uOpIBrYvfE5XwFohqu/JJ3E4+T/oF
MkaAGmaOns9cBfFw7MrtravjBAUC79T20nX1KbOM3E5hcGQLmWt27WfrnE7n81Ee
wg8csAuveDsL22omJ4oA/IGoFrKuK8jagIqdVwwWk2gWP0QBsQx0MRO4cQCjjI95
5B4lgQl3R41KqxWRrB4SYM+Eca9s6iD2khUrtoP8EAUaQ3ZsCQIqgYvw9CGeuY1C
WQya404Hn2+4TqJI+MKYIxG5+fOXbUH7mDw6hubtOf+QOPZF/qmIwc6MdlEIMUw0
BQQ5ZW2Ap69ZoSLKs2HVIPDoiojvGi4ILwv/RI0fpC8+QTqT0Bk4fXdgN538rkxX
TNaV/oL/NafWmsgjKX5soL4qQBmo8Dwn81omK2fCYmVM1LH+ZrSm6PigebQPNO4I
HW7FY61+PbGRGxXJeCLx3xPBVy5Qn+4DSwLPzRAT1Sh5xpyrnvarAqUIW6mFZaBy
9G1Y69ItE/X/NHqdTvzH0Tfp2EODuNmoYxRxmapb3K8hhVRW41fNcHdJGhRy1r/c
Vi+HdGEkkYpdEs01d7P+KAZ1fYHmPnT/ryr2ugjPDwNQkA19yFxN6DouaAThkmqL
HCWaHbbb1u5RGRc7Uq8sUVDAK4pYIwfrQkLM2L70p0ehgo6q7bBL+PHKHP6XsgOo
vgTnNdgOLZrTyAtKcuqZgxkUlC4MeYwKDn6VJETTQoSb247O42GmFADB+LEjTO+y
oU4N0hScXr3suHvQVU0WRs+IVM5jVcxD62ipZ7iEGqRfljM91JnFboMHuATJJiUY
u05HuadrYW19bOu57J4D4f3+a4S+MToK6xhka4dkWy+iuqGGJEuvkxGWTFramLDU
gJaYwGgIvlTwJAyaEy7skvrvtMcr4OP3XPldIfB7UFy9B8PLU3ZucNcNnovUnir8
SFfPKTdXC4hq3u/TIMpeJX1knozTmZM+MWvNCElnKcWHUpvGGxMnMeVn6Japv6nk
sMx4G1SVpQYoVLp9FX5Ch2yh6xKruHRVBSm+6j+JXkKX7Y7kLsmyAPbLto035z9V
0/u9BTRMzPHYk7G274l+7h1c/QoxawZwJYaSMlCI1bMbLqj7jCETv8A74laYiacU
3mjk+k2cJ8WgNJl2S2ont/uX8BtgHe0bqIz1nGQks4+oMjHYsRn3rhB47ifWlTXe
Qh6E+8PAMbMCLwDdqQTb2bdYQbEqCGcG9aLnEw2iWlcWufpyBH3XOpeTzKv7uljL
ycecGKIsAXMg1YBbzlfy2WMQTAN5B+IEaexpYUfIVeO5dzp2PmNVkdrSaNoW8yzk
XzLXdNyrxecghFgxa82GOWQ2TW9bPoDfiqB7EuRq5oY5CTIAvJhAL2RlG5nvG8Az
BkcOtG0WJXY3kmU1feOmG9MBtSv2p/ttt7Kzu5YXFXvZpMhXC0WLu49NJXSxStEi
DBjRZBzV6OPpJ2cwirQSm/LWY8xch67TQOtO114w8f0KPL/r3GrvZZId9ibqzKbL
KnTKvqDzWwhFwg9GDXfG6Jvi7pq+pjET2yaH/kiv1Tui8ftlJrGFAdKrHJZANFKg
XvyVpeXR99pHaFmZEjvv1dUoKUiUL3wuH4n433mRDwEZ7Ne6xCV1h2xRdvvkpFvQ
Ln9plXlptmVeURh2gnHWnDOds67o3+2xFuoMhIggjhSL3ul9EO2Z3aj7VI6CCtaQ
lWa/fuOzjUPNdD+JAI7ehmCLucb4N9nSBAq2phxXwBJ1cvB0gi/+HSBqvGN1S53O
7+b1xXhTe+kk1BBfeX2FktFTSQt1kYzdklncajmWt6dnnx77Fx01sBejiiR5sltC
TqV7hAespdEhIInrrxSSqoEf/OSLfXcbtccS+HgRAEwQBvpSJQB6dOcNmeCaJTYv
zEMCXGc2DCTGQSG6Bpfa3IQLfiR+8KuRwvi0akrnMBztkAOwVPH8VYl8zPTrHQDa
1VR6V2GXHPetbguM8lCTdGZPwKVfCl6u7kKBKHP4Mzks3dC9n40TKxD9/VaDkbc4
ag+S6Dz8fYPjM9ZZAx665KbTG6QYT34XZvx1MZ0QSi3MPKTsR5CL1X9xUtaftTIY
Y5rqzwRFSIl7UBbVIfeJrrssGA3xD5hH/f8S3EcDRYZzIYAkGLU1NxEU6jNdUtP8
hhelmr7EDt0wgcZXzS0AUxw10Ioehkmlsnv312g0RFRz29+eOjcFWHCqYVvm9F6Y
uhUenGa3xDWpl058icFkD9YuFX/v7YjdfW9GIl2U+KuXqRZkL+ihAprtDdWHdWCx
du9CG1s09j42hVB2ReDPZFFemmSlmrJLj6/vpHJdABNwM1N1pUOVUYOKx9iTvVqY
k9ZA6EkiX3w4RUg44Lqf3rLb0FUpguB0Vb8pe6mWYIyQEpQtTT/eaV+w0Foghp6R
S5BgfoIeVYWg+wXzKhG3zHLmL7Fs4LIBqRzWZ20zrorGRVgvyIElxBQKOjP2gLAl
/W/jikmAvNnI9EJVsPRJp0kOLgoR0JsURBPHev8k+B25lPIDd94VIgrkf2kjCA7n
gAVJsyhM21UwGQXFZz7ixNEvIWACp6vh7m0HifDvzaTQOfShn+Zej4+PMtqyeCGV
D8aMrHSNmUHIkRwk2GyF80UPxR2osr8YW44Tvy+Q7jq+WoCaKT3t1AJDsQdnkjsM
tfMhmucBjL7bNo9TSJQcocnRimo+nNqjxI8XAYBj3zJV2XnAmJ3stBnqwfA8TPTK
Y+0PiZEWsuRijX2Zwtf1rbkqVHuOdNjEK9PvAsQueuaE+pUh5eKWFqfQivEe+GoE
yZiPT/xne1I65VtRRm9FgX6ik+XVLEY7mfIWc0EODiXeD++1Rt63yCVjXMvJUdk6
Bt8qqT/pDLEQniZg3TNIMb7x3O3xzTTRzbdYwxS76H7pMGOSM+0Z3SbFL/I7+gDt
zCtcGYVe5/75K6AyJGM46EW3/BTq85qTy7xRkr9GvHwZvbqIj1LLMPvWZq96xNEB
qf6zL+8kzSwlV43OoNrpgCe/TVHiSQwHxdxiMkhVu9TRtxqaliTtGZw09eGFbrps
SQ9pTA0sg9/epKyQQdmhmZPdJQhc2BdG+Yvn/Oh0yzCg5VxKvuKZodWZ7w0MOkR8
U8FrYZacCT1arpqFE3VmxFNzGeJFVIhAaf5ogSnCHO4g80mCmuK46F6dXHxhCly8
IASSZ4fY2Vx9S7ZbQjZvBy1JO1+HuFgwb5TzqPCpzQL9kEX2j5aLo/ZMtUWXJhtf
I2T7YkZlXxbft3wEZ42Nz4rLoNH6Hi4U7/KY1rJcxsy08o8ab05q7PSWFQtrXJMS
MWgRxJI1csSG4x797RaRGxYNK5CTRVAf8LSkhJgw4IqNIfrr6KXb0Q8SRxBJ5nC7
oQ83oKse91ydzLWgL/2lRRSPVkTjkenNzVb1va47GdHXD7RV3gyJo2+PCDfp7cS7
uh+Eapl4SBgwOvagXVhArFqox7vE+pFRrTxf1JevNUWT+t1OIlZRPtP7Xqx1I2s9
XOs6qHg1OTH5+ONa0mECzLNKJBFPyEvSYBur4qss2s8/5hW2nmzXBIg0yrK+MU+C
XB2NHa/FrGkwhWj5U29Coo02Oa2Z0TkUoN/RffdZRHv9fqYDC8j378vA0GIFa0uV
r9ZSCbR0BIOXLOky7RHz7udRs1Ffz73rf1kdz3XB03SaqKw6fKEUzsfTAaVdF3wd
Cfm5d4rrmdDtyUArBCxLQRhnCSIzIVitfIRj9O3hHKIWY4ikXVInC0MNn6lBOWHD
nmLWQ1fCPQBI5WNFx0yKArgwXXdZu9z921KYmUJGfV4qAvA2syq5Ora2yl4FZkyc
F6kSm09WhGk96Nna48GR/Otgd+DfTEleuVIohr7vSCDKAIwhJXHNseqLG/0JSnKW
X1gL/pJ7R2Ml3kALYzmnEzE7/xeiuJD4sHa2AfiUJC4+iw5Jt2dbDNj0EG9Q1/ux
LNT/ELi6x2+CW3s1su5hlPdEAu/kR0QEhGtfSmkvcCUOUPtJkQLZguDdAFfDPwEn
T0Jpa9W7XsMCcP/4CVSno9DQeSsB5InzkiOZCA/ljFleEpDl7Jmmnc10cFWCEjrH
YTjD+knhuWIbb7/bA3q43iyHKFMU6HLEGOgz1plOFvuRmvDOOLWs8w2ieX6B2btw
Dp4/32f/BP76P0fJYK1dU1U/1hLZK46+WlP+K/H3ff5wpXu23btZ9rVNp9GT41nk
5EChsgO0pc9xXQvkMEC/XrqrfqXQW0zzj6Djy4LP/RMGI71f5J4VBZ3JZFEMpfBy
G9PtfO56bW995DpKD/BYuZEpRVFn1N1vdqfHJa1tO43/8nMb7pN9AVhFncdUEKwR
KJnX8mtEBA9M9nMus1nS8lh+Qsbpw/SoKphtmsaa1uFYzOzDNJFtN33Z/e3PqrOT
agVz+LdemTTpINGAVglN7oFIcS12HqridPXRCxwtLqb9/StNO0VuBrQ++2v3q1Sa
kJ/LMD/HrqtGauyqaXLGJ8p7loY50GVQ3GISBhQbO0bjsS9jL2hPoYa5kvg6LqTW
gi0YwhmuXHPJkFp0kQ0jPLCAeA4pIHamCW+UIMp9Ih8/RAj71g+AjyrGBPxTb17a
c7eWUJg1CGne9/yOjeA2DHMymb5SmASV71wRfh2mwWEQoHkgwZv8rqxIfpH2SX3a
5c3kcUHdBRDKl2XQK8A6EsPo5EZ4VGcN5rbW5/8ijuBjp5yxwOTrhcCvET364wpz
lQwI9+mbQOdBafnU6m/ohjknFIh+UPOJjYhvj0CZ+6WT2wOyS3xA6I0QKCn/DoHh
lodMgPE6zjuvqlzaCr+FqlgCeyYr3tNBY3ZbLXYrsRcQFNO4ALaRgxO1SixGQlLA
1zaG3SH8vpb1dfmIH4HL/9aHTNCwt+Kjhf6DW/WaXh4iirkJBPTYGysNFPyuSYCf
nEJllODgY66SDPkbEj9WoydTFqokBmw2gepf5JVi2p5Zq+3j+TZMOJETj1LzXdiF
6fcF3rHbGIUWczQHO+sTHMzbR/X0rsDR4U1gAuA2fMrNL4tqoeZfWVURswn+KiAy
0I198cT8fw9WM0IuendZ2L+00wd3ZwZMyoXemHDAdxTnv3wcKx1l5Up0lQRyM9Rb
EbaqgI4KX31D5rNsF2NQZWp/OVze+ZQ1RWTyp653fH6L/315mBtkaf1s1/6u+8sT
rDCrWS5Hdi3nuCC8Q36Wjdb6e87BJYYDILMldrnFuvbOoLOwOYoP+m7FDav+tnta
uhF9k4R/LPRp1Hn6WtFcRZ98iCLrKFVodQ6tP42d7CUbwLly4aOqPy4ostsramtn
BPSSGRen1Dl5G2S5GhMAH9ePbX8GUJNvcXO9x+V84M07nWoWqLAwEcjulSRxnBdG
+9X1URez7eJI3kxsjmMDMNlMX+VKFt6XDABNcfFh4RR2bNy/0Y0Nh5yXMSziSODF
LhW3rTw/hiKS2EomyUlXWyVIRi6kdd3rul80QAEjkUK2Vn9JWOClWbOAEdD1kLud
+GSu0P/GuYFZ6UkiJsExIjdcZTXA/TGNknMEAmrlI5n2LneGB7K1WWIABiWZkcio
3k2kyIyMgxkyH/jx7Y3THp2sCRjTC2njKYVh0TRj6WMNKquivus8JL8BNCt4F+Mg
uoq2YiiYThlpMU4OTL8j73PsdNYUkYkEt7R/wMozQ4J/M9kNo5KCleaqQZg349Vv
FRjT4lUMISRTCNJZ/69w6d+ZI59hlFMqXsaXfpVrGOGMHIzzUKsGR1P/tCcQX8KO
lDbCkLxuWjkL+7IUmkWu1ZRFfzpjoIGIEQdP2wD+1iRUfeZ7Ulw1u3TWjtW2fZd1
ApTJq53CuM64gkASdI8UqYBfEqBi8YhPMrq+/VyyvjUgUeH4W1H5Vi11gHnlzNsJ
8XrMBHtShmYfGVCF3NtBlrm4Yq3AJ98ajitWOjkPzOyczsOM9xrCVohOHiIqMRYp
6WiNwZy9IZ/y7aRoYYEwY2Z3UyETdIMbVcP+a7VMCDxU6waaNGSTcPCgNiWONS2s
WymEPfY2uhd5N8NQFVCcY4OaIWnQ3F2d4rp47mgqRyS9GLvaTYhHNnj4qE25IgVJ
S6vUTxat+2hid/uxi9RTLQ7ssYX+hWSrn1GnfshHPHpRDGmRlkuxgepkH/RL7RME
3/CVLYiHQXTul+RL1qZMhg6SJaokX0JBE5kHcU2AyDmhBNCSQXY8x5o4W6SLEtNH
qAMldROYpBGVZ7kxFt/VMn/289SvVzUk09YxI4lVkAYn1PukXwcFhRvr/zMq9C33
jL7vGQHgbeuu4rZaKys6qlnCeIpiWHDsVPm4h6F1b8xYRhmrYbVZMs/nAJw+GaNu
g7ikqTLZWQjHdInMt9u+H7n34Y8SPaYT3Eo+g4E2uE0za59ADOQCOk/B749W82lA
FVYONrkEdqDQb6iofYkCOozCPJgKuLGWNegE/1sDYZYgh3bNowlPJqA5kASLjqoB
PAw+6GGlof1+68AXpH8YR//KCUUGls1sFKIk8tO6sCVgXo//imulBIx8/r/fbV/7
RP9iH9ryabSwPi0jH5X7t0AYD6jeVeMjpkkuhEfUrCrzdn7t5fs+v2NcBkh8o6hH
apojn+GXk2dsQItoXMBstX+wnvZHN3k3nVrEPlQqOwVU6vwtEBDBEuO0TG3iafpP
0e7Uq+CSkRSq3r/pM6LoCS9glpLaBAmSMOM+mb/tnPsd4OnbAe1hSFRK9x2rjiMU
zrCyUv71pb0mpMR7RhmYQ1tHVdcQcTMjVy+subU+mfYwdu1ndrUjrATPU9ZogRWT
EwXKIhiZnuaXEyYf+qVvtOb5/FZTUgX2gbhWa5742FEx+AFOS0m8gAMbZsdxKTao
0sOnt8q/hJvyNq8yJWIwz3vB0bmFgaSZNRsGfuSDKW+SS2qUrp2gx9amAFF36u24
D5dfck39gp3KObUE1mvN2vXUBP9KI7D44EQ9qFA7Rbx1xFwPrtO9xo4/T1jBIGJ/
gv2QuTcireFiM7AbQ8r87RC8e7DGZlOaFzlp390NlYmDSGj2wZcPpgovkKsv9ZJF
OPCu06RBY//0sN4C1btbjKG3t5wvy2pRjDRyasRrcUyFnuHj0fX8UoqhYuey3yIl
SIBq/NwS81Ckz3tLqLQ3fHGnY0mYfS1IHQ0r0U/D2SZ7/WK6siLmmfeRnSHw/hxW
dUx2lChnyKD6dM1mfOVlK6YGIsBK+Rjb7+TPO8PzxdFUn/o5UFmlytYA6jVv9yjM
et4IKqaKwszeefnxz3/55zkepb0n2Uc2AfRds5NC8uxY73GBzwUrvUmhVwjgtAeG
sPXuipIu+VjQGBuDfsphS6xXFlpuqhVJlB6E6qBDXP4pZiIeTs8TJHWZ2nP+IcJE
gnKcoCTPGp206f7WPGSebZcCP/Cr5LPrhc1qwot0cXQMlELnM7wBM0vIsxMXHSs9
HB2W/hWTstzh4L+U6Oz+CNTl8XllibI7YsPvd99NCQoBF4LEv3CUssuhMB2VkBwJ
1+Ha82o9FnCOwZ8MDRLOF6ClfdQYMUVFyiO069ujuDVQsZCKBV/zupk6fA1F8Y7j
yiQLbbJbQoFe17OQ9eifB+yi2hpQrluzkopF/JAEXwshJ6bjRUBmvA/VFtXZI6kV
xFqISpepyMYeY6U4SrN05Jul8m3m/TfkaEQZoz/rhWQpGG9d7TPbSNP9u0lba5m9
ELCCgUEPVpjLUA5b4fkmduiLVK+FZWK4QoSdCQqu8zhQZOxrQtgM8sFRie62VgGG
srKnSMSQGrgmi+gR2aD1RPwpNUcCowL2CzS1IpxlSpotm9XLPzTu2YGqgM4lwJvf
juaR2OwLk8bX7eTgA5o+waj2IgWFBGrpOEy0KxCneUQkwvdlrXebGrNVpJWVfSL6
nCfiboVFfQm23NtVfi6c8eoWlIqF0LfGyrPzNaHGNXulZXpJwXU3iw9YvjDkxANe
bcmWt1Sy3QrAjfU8VWxegD3HMf4pge3LvwYRnMJgfesBl0/hbsHNefPQei8GBrHW
3myv9qH7MdzExCxobilHpqootMyF525o4i6NrUGjyngtPkv3gkqWLckg89bnCHPJ
ECYL1M5gD9G35EFodmI4WRfJdXqk++jI8lRy7KSHS1ByHtpXxbYFgYvRTj9pr+QI
wXRyb6Ib+ZC5p4vidmKRZv4/X+UkyDxDa5pVVJMyKuzKRZGFhsdP3KynNx7lhSY5
cdLQ9KaqcVRt7z1+X0NOQ1z2w1I01OUXYB5cxF0mjjdf8GyRHdltQNTPID7ZKngC
/EyWODjsVJ9nUQgzAQeM8i6eDIE8/XLs3d5mh27Pyw3NACudYjSvGXhsM7eGlaSP
acpFG2ugvPiBk+TNR/nXKr49QrnCWK9cqc8e4uJnoBR6CTOT82RaCqrYgayhDMos
nO8zX9WzRuTG2M9QZZDvDh+Pj6bYLdYaEGsn6HCEtmalv+IKtcQp0T6oWxaq3xa6
43dlYS4tOWhVxWRQIj0ealMhzowXlOfxiYfB6hS0fsypfxWJN1oy0iPIGcHjnSgS
O+YbzXUeChCCU2yPFBprovyEZLFgyp0I880YD1dmy7FXlP8/0xyo/iGQFF7tIHUq
EVduN1mbySYQY1z5+rVOwZQvoIa2DLSMW2fns18AKaNgdYC4d/j79VxisTzV4mS3
Xw3vasx7yhGsCsKjFNZ66dggQqwj+3SAysO032yfashA96EFKFJAZX8rdp3gC1t2
/9fUdtTUg2k0NGgAYbZnEs9M+B32x5Ac8Q7LmyTI34omAiiBPiq+7QYonNCeYssU
oPXpL36/4CRExmFNLR4OcrsTkM99XBxkTBv24QwdyKZeiHTw0yfpiNGh/3ZGpgAM
Qz7ZbEw1OKUoby5i7BPd/2pJ+p+fBNPF1r3+92Riu0Z68dZu6OwZg08NTd/6uu6U
C1hxZuV2A5BC0nUbUYfDQR1YZuz6ianydMf9BACz9qxiMl5Z+QY2AkhVl7sfVFEE
iFuKaHgDSSnPN8CyaA4q/SzJiQz9XgERU2N6Nm9U9jOJ4rfP5pZa/oYLFHSIPWVI
SDatCzxD0Nnj6nZ+laRNcmbfNNIvbCFeqY37EYosQ/38ogrIjcpv3sEEqmVG5uHv
p5FkL57zwWd2aAMROa7mM0Tgo+Yd79lgc9iixw5hc1D8/lpaTl7xwzzJNz3pbVHl
fFWDwvrqaHab/HvmrA4iMm69ZkNuh1cNqTTJarjFrJqD9+JRHYD9bEqrV+wElf5n
Rt+vyeqL6C6b0O2wfMlOiloWANWJOJSby0S9J76VTZYFK6WuF1F4+UOHqVv3zyjN
v2lj664NHPBN3xGctzEQaG77Jkv0boLSsEK1HNqZWijHfuBs3OIRXN03jsqm6bU8
PULkTknSDVDm9gGBVBkpH/L/lmv9Yc8GW1PvvKU8uzbvoCvhYVo0x2B98eU2av/i
KvQxu85URlRG53hjWfRJXXrKg0bIbZgAdRmvbYZxS7zrYwBX0rKeW5+WPnjClQJh
TaSeFql7uJKGR+Ei242bp1TlSxB/MY9XxoNfGMf2gvmcwKDGK2KhuWbEAbORlM7F
CI4gQ7RSsX2U842k3Zp8Wuab2D5o34fOgf+kiVSRK9fmPpg45qPNVPiqwGgEnjX8
GKiND0kXImhCiuNmXBCYgJkn8XpOSoIhrvex3RZVBk3g+SvV8mqVWN4L+n4UUuIl
Vu7nFOjVv+CbWYajde9kOaQ/6NbNlpx2sE5ZRG09N0rQ5eH46OKmPdjrjbYIO9Af
mGREgSYraG2rtnJdSB/6zh3mJHW8d43XKwRZeQwWSyP0yJw37OthxKLLx1pQQrVZ
q29KqszYZPWdABDrNSk+zFubN99beiB4l65qKgslMX+FgmLlvBMzCTyoJZcH6RRB
L14kZi6omh3ts0MQIYuL9soNjKNHvhU4e8/RPFXOMv9EVOnJpb0UItDxGVgYTLoD
G3D5ILZhe/2Z9v+DjThNmdH+JDlmkiU18vXDhXWnj/eWwA4EBA2nkgbk0k6GPUm3
apSO483OY1jhOGHZk6XDJZQk5vsjKhmpDRdlXNcPif+KH1JOtI4CmnI4NXlu4qnv
3RCUTEgjumiwLt2QPcSUB8LmbFfgK4fEcxvhb2fJJeS205ZD6WvC8hmh8P2OxSNv
9qWu6d9g89l86ybUT9buK4SBJLvU4zaeJNSS7cdTnQI74tH9A8li7+ReGfco50pd
5gwjmqv1/RBF7fKtQVUYJ8cyfjxz042r6iAoBjJhAzJOjO7g6XjYiEKAC+2wyGoT
m7pofRVunwkAbX5ngsiwi4N+V3S9ty9vOd+dITOl1GDsCCmfe3SUdOgamCGT5xy/
xtc8lMUy6enamjNItgAvffZj8XNTDrHyPXnQEwj9YD4AnGVniKySpKgiSOqu+B7P
RxCjvaIh1q79a0e1gsXzJvfBZU9rKUCUntMf1lPlu1npYUud7e6Is7M4cvMpJbm5
LYlBt+/QLWSqxau1PEx6J5xo4Qn/fcdblbeRJjVtlb/NPSNpzJ3d1ntL35rzGEVE
pBAP3rnsL5ORbW9M9/t118WJmHlnB8phhOQjVWVrzE/dfmGlbSgaPGb2Bw6LnOTt
liFHrLVRV3VVibpc1yW+7ddM/wTyGf4Qm3ehNJT8RXwubeVgkdkweylffoxXvCHN
GPa8hArKkYZcdsCgGIRoP2JrGdyyeubs4qe8DsrEKlpNLpt5sGdFOfHWdf3KH29O
+QXhdM8b2/XVNKQZku3IyQmYBzkxKw7VTdBE5FxfBpfxsuMmLd82dtY7dNbwG3Be
4C9d5GDMooFSwNuAL/Lv9I5Eh5aeG/jf7KzHd+IYhYdNQ4HYNGPYF3ljtW5Rmo1E
2CrK1UKDymtqa543ZHXNk6UN32V5i5JUpZ5z8s1bHWsJha2OqKDYhBx5w/kHtbuE
g/p6Sb2Znj+uZOqmHWv//J/0iTSq5hU2aAdGmGRrMbzzfyqybH27Vk+fAnpqEODX
fJtiU0lhrVkmhjn8lQQdqv49RGOYea9IMjtBshzWHZOLFouHQAsablZB8Re0Pgev
B3BdO5BPwNDQDnPlEh6qtkFXGVvrgVWX69LpgBHQcikZstdEQT/DLf5gXH3p4ixq
5K0gINVc997BUj6B7QbQVOJc8yMHd0C2ma8QWOm+yAKLZD82fL14riTXi++KZ9MG
dyxwyDLv0sC9/AX99EAKNO8L010BWzRUy948Da+niAaKN1NWgyRz/KObG4fJQVW7
PtlOFQIPvpdZil6l6Z0IJfrU6eaC2//amMpxFTG4fI+v8bZWjereVpPilzIpd6/g
ENn1PhzQpcr59SBmau7r0a8hGh97E54FspJsTNAYH8Fy3HKSiA0LBqW4reovCIr2
tGHbMLFOmWN+h4xMdyzIJgMdR69MuxN+2usQeAuOZ8JiHYo+vkrSv4enZT4YtGKL
5Y4tBUmZ1UQwkVeewrxk/8Jj53AlDebOt4LJwCnIXpkVxvHSwkE8stwgyHXSgP0K
/OGnf2uNoDQqF+syDvDu0ONoWFBvpihYHqI5I7ujP1RQevYYb+4znI/KoBh0CC7A
Av5p9j1jiv9gAWZHRPnADFVbx1Lrde2egovsZjAHE8rnqXPLP0IgOJQ2237E0i5a
+/1DQhhu+VKZeNjQ3xBJUrjnyv0S0py/VdXEhq5CYFm02v+J4IEPC8XxJ8SJoQbl
8AXEAEi0yyYHrfWIau42BatPnz9C8Xu7JG3XfqpZzfIYIJBtcjOZuygT5PjbXx5w
ZiMWa/swFNSeXYgGWoFVP1EyEmBJ0HyQFsk2xMha2Ywk+u3t+GD3IZGKwmGEP7dH
qjGxLm4OL6U4P4mN3jAIssi6YljCjBYEjYVUskZikNyBIh1i4PCm7YN6teFG1wxq
hpENZ+fYc8yqR/AbAvbpmJlR8cZ/EPzOCAcPOT3QZP73wuSFFArSynPSr7Za3Y9g
wIjFkb3Vp3drSOHlkHITWTRRVpFHVMfTuC90+WcpiN0bsSHMoHfOpmcTqbcrKzrm
UNEPdvv7jQF8Ez1SIvm4gHMIEZux1D21jRRWqAAsSJTzpTwxuqYOpFPQiuS4u5wh
oDyCLTiP5gMsyJbqAfYw2FgJaBhVuQbVWrFNSrjPvofk6DoHjZkaXKC9rfh3WNVn
0fXbdSljmdz62l5uly2axQSznzp5H5u803km/M3M6IML0sIjbqkDH+bqyAUDi3k1
Pq0y5rNW96N5BQHHjz+BHLr5A5Iezox8pF++/62geUIG2TKkM6pY9qyshJyklsZf
/WVf2AVmP9MGGpcvnQ/Ra9jAZqqh7VH7uOXCFNutJIwT2MgWFJTDXJx4OeEhNSxe
e57ayIbntNmYTflhdJmL+ntQHuEWBFdBzNQN2eq7sWLgR9bWehPMkF6ZeD5bSEiS
4ZFDxXwYaNVSgeiMEaUrEa5UmucLnp/+o8J5p7EFi496rkkTZf9SMy7D450jeiYn
UBOMhqKpI0D6GzHQjOGXhGQQcjXe26Z5wGEuSDQ4LDBVbcZs0vV2GiF7rGiEssse
yNt6WiZg5olTB4gWrc1q5quZnyoVvxnXD/H4BV+0MpdRPVlGLsc4kCLYpcUS/Evv
woQKvRt9z6szRuQ/PAFWMINkU+mqLS7FAfd1tNKr+KpaIVfn3U6tfYFbJp/61xC/
yWwmCdGOROpy/B8UHXhedkNEiGQzy6LtCo8VNnCnA7HnNW/niZ24Cfd1hvrdLN+A
lbSX5zdvJzgXXC8sJVZWH+YRS5WlZ321GNSkRG9nef3G+3wWZ5gJoD0DVe8EaxjH
AquvX4O7TXd7yDYP0ibHzu/lHejKuRPKEDDVcgAtPpnu2AuDHYtYqSVzr3eeEm/L
U7K8uXzsXvlUyeBByqTFiaScJ1nir2tMfA7s8vDQWhjIeEEhwjx5J9852jA5kaTu
4mnNo+OaMPI1IAt2W7rJuO2T5noIuVeGoQeIRJVeGRr6uvO38UUdlkwEiTqY2kS8
1edaoXhfVkNJT/jmeCh5dtekcQaNOzevjzjZcTmlxc+sSQzztOAr78fIIhhqbvaQ
H5H9YDjMsTEw2JwN+xcw6pnkRn0Sr4DWLK80cOddmIoxiusVJoIeXPrDHq63n6rK
amxS6yfnhDxweE6q0nygDg72yeiF65GUBA37TgAMBWxnwpiFwyEjxAgC5242vcI6
P6f0qo0XkFQqoXYKXh1RNZULx7Tl+puBJWwZyhNGrkuaYdtFPcny3lbzfoNdnji3
xupjf4TyAxi/ywmEi69WMvaEl+lJsdUD0aEheQrN1EENpWlraZQGt8RoJBXWjIhE
Hx+8G0BIfOcf993rZGyENY5PUw13VbIblTna+43sfw+eORsgm5kJjFbgMhbYOXY3
X/ZBV2iXAua4ctLzZHnJisd18SJK4RX2yipj9mZQ70TGfrWcaXCtR4c6FqCf5z4p
epIKjX1DSyNhoeOJYCxHM1dTqFPPMKXBCNqTdtfGM8pcfsFaAwEwzGkjRApzMKqE
DJF6qzQqRh3YrO0HwxliV6HMWlVSsEolQY7tNlAKnYsHe+jfTRAjvO0GypXRJCCy
/DpHWIOi/QiLOzhqReVRGPBIfR9XFcXiJwNDk8Pdzqi8me9FRX8s/CIQ9rf669Wf
U6D9W56bBesj3edGyG1uLRPDn3h6H22wfJEvjw1W5RT8p/v/mpWsa0EZIOobI8Aw
qe7DwEjkNv99gNHzuTTJse07g/Vz2kUAQJYNmlSYfKW2yBrS0reQvG6wxTdX+3RW
fTd3qV3hEfBMDSKAGt8at5KH+pTtQ0C/w58Ns99rjhX7Jk+0zhnVgqID8EPMO4c1
x0/XGaQJSeitipvgW1LKHq8Hi3pmp2KWDXi9t06SLAmqZO0EkPg1f7hUtEiRmHNT
uE1Lulk48n18QZivIxoWH27xkU8N+Dv7KKXF4Ba5+nHAMcfjupgoEFzkh+PeSRqg
+2p9+AzS+3LbVJbItKFoPIal0zS2kOwXQAgMQO8MV/kLc6k7DP3IFY8wJlXqtKnh
Gp2Ni8cMFqKNuKiZxPxOdxzjVPpruLhxCVgJtZ87aMCA4zCppVIZRUQPRRAFO73W
G6Psj0ZRZZkL/R+gFVJZiL7cHGsFmGmrv0rylUrDvm8Ek+PoOnkNZALN9UU+Wrp+
LYljBlw68DalWbmudwH9Lk9g6TPCnDLg7s8FHtcTlrViMQtoSL3d+yMzYMhLqolV
NhXRHKrgwbhDCKcpg1MsAw9+pTMwiae0EmdCbU7iy1kALzyoN59JgiasjSdOcFhR
BI5bCDjjkRL8uvEGnJY7Xjj7lB9jsrMFIA93fm1oDs76LZQvovDcWx+NOmQTwRaN
1sj8DmI6FSY09OqdsC3mZkMjIjeCwwAJTo35eDXfC+JQhBPoMG8wY6Yp7BAEFGlW
5x1MO6BfL1EOKlSzbVBIvvZvCwxDz1sk5tVB09eAKfVZ0Xn0PJybXgD9gMLd6mSt
KoiAoFjceP8vgCk1WEfq8jnGD6my/eob+M8atLRxErQRxwlKsZzVcB/BT1f+CuWH
LEiI7m5mOHNkM9CopPWX50v1JW3w2ozLcoFwzTJ+IzazNq+QcmyrhvX4Fr2/oPoE
ENaYLrOzYwXR9bEkAY3WmWHBgKS0telhdFarBfgRDuCizl3MjSCfOzqMdx7GB380
`protect end_protected