`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3792 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
wcmpwSk7Xh2DEFViwcIwodbbDLmZ7V8Ty/vbMb+w9eH4srpA+IXKl2anIFkEV710
RxmiAy+V7M4e12UY2XF2CEVO9hpct/RAr/q1T3Yb26Say27qMG8Ro/oFD2zC4pXs
ADWesRj2ZUE/rdXo9CRb3Z/qKVvKYZf45oaHpO0WegaegP6an16Q2m0TTVeatoJs
0+Sk9Otv6qaOe08hEmxszEYzQajP0SnL2XQx3Am3wpZc/34CKCgutEEqdyS3wXby
FLQ6RGjsSRTp79YxgB1a7vqbpZ/knOAhDisNr2oNgu1+EQtp2rH2skl7BW5Tpj8J
0Nes8N26ECjyn/hja9d7O+RTkAweIDF89/MGV5xeaf8ksVrShivDlSE6zTVJ1upN
6KgQyrGcTPStPGGJCEDYU07M4+wH4h5NlUAjZ/fTRX3cVMt/g9fuCXKFhYEQ6rPC
NaaKLLqQRghGhLHHqtouPkYCoWc5M1HpvKWvOLo5MT+Wgx6vQRT94qo45JRYFLFK
U35FlwUB8EF0PmN54Z/4FHTrFjbSoBf4AGWY6gZsR4ulps4GSjp9cin9EhHQe7Lu
uVY5lMqyIvCmGp9Oalo7HN3PQjm/GdaOc1Q4Ie+fA2rvWvoaHKD+tcfJ+KBDEnZz
b3KYQVHiIpt5Kefh6/sgKG2xuxgYQ1EL2HPmBKF9G6c+1uznHbonpVi6+sZP4PaO
G6wANZFnQXn5LeS33naY3HAHR8r0GsXdOHW61pCgFsAm/+QivX7YMjBXg0lmN/RR
1eXQpuE9jqxGPKXhlAQmTgckH0BMoWeXkVhlJcd7EanHND7mGNbBcNvyZvGSpsJR
sH5MlmLyNWPBdtk4kmm6Zxam7J5yIaOQF4Zf3X150JhLrGVSVOX+nF4VekuYGJ07
1Xv/J6mqiemUWILlwdM9WRA+nXdzPmbTD57CekL6RwdXkz+gIP5D6Jj2IFyatBD7
6vJopS4FHQh78xQkk5ERPVLUP/O2kMmu60/5heJGJ9IuC6CvR0durUifpO5HnTcg
FJjgY0rQ4CUdwgpbf2AseWzpwW6Vwlruf6lueyz/i+57ng5gQSa8C47ifMySedM2
Kp+Satx6Uk98jRDfvnyOos9+R++JCPCEbPaUZWURv8+d4z7YCXJqL9ELa2jY9ztm
GMEYcyIq5d9/jQbvA9icUv3K454zaRURhHt6uZUCA7vL0TF6hrT2nJN7qFhAaUPc
wryvIMfUXOAp92hx4GlYdy1uIcvspwnP2daY8IydfrXORa8zXF9QLN0bD0H5/aAy
onW+G8PTxKkqC7g69mcAa+f3T9h7MSb0zGUz9G14h71MGb6l2GK8HTIMPeV2UGFN
+bGefMWOEo8UioyDMwdYl8HQ0yl5u3pldmUPHyCjaLqTicE5llX+/MEHiSJBc/1N
q9LGuGnaOe5UmZW3GSjh6kXEMLM+6nr94l6uQ9lnHla8vfwbGK3Gvm6sBhQHBkjF
RvMF8G45Bj/I2xdOkQ2FoG1JIC37YQ3BN4+KKpby4Fe/zkDBIGH24OkktV+KTNT7
ppsmGwSnOadU0Aq1UyGE6BAWBcaMsTYpv9eWS8HCmEoy4Y3jbRuxvKb23IwcCPlL
X0EugwE9u/arv7lfw2JOSbnTn10NpM4YY8+Aet23G6CwenwNI/pq/whGJfA3xEFn
Z6WtH3F67nMEM/jxPfSodrOy+6D4RuWK2y2VVO45CBHkn68ZsbQSOPTM7bnUhrRx
SywQaQZkHK9g3gJeJHDdjbbFlMu5SgN99E4UIwwWh5GmxTl3RcoukwEs/lOghm34
J6EfcQV/WNSGqdhklWyfy01PK1ZeOMuo+BeSYud4+zwODYYG4TpCi4ERr4IxExGy
4orbSR8U3UcwYxSXyn2ig1LNjcRpiciYEKgkNwZe5nKLQ7DKo+ELENH8p4MnI4vg
4l690brd6phg1dnspcDN5mdPF+EgqrAYFDemvT/BakltT9czeBi1saBZFKwd+iPL
PpNAd2TGow09ElfWmJHLcui06bKf3c/fL5dA3/1avU9jpH2OthJG3MTzS/v380TE
5PSLLBQZb1LNAk+KZjOw9jS7Uw73HQ+IL2FQKQ2RV4+BOg2m5w2BUU4n3JmWUR8f
84eblI0E2LLAOAEwKvq4db72FgPdCWoTkp+OzXxMWvv1YniHo1/LfBUOS7z4UWMq
YrofU8ANEf00xJiQaKaz47ancQ3/5neEvWwBx1eiH6Y8qCppIEKMgg0GwdnTGDGd
q2JvHAHGpBrw5WpHFPv9E7hJwkuBBlqxfiNKmO6AlpyrlrEZ4rD9vqhi0w3Bt7XM
BWSfL9tnTPm7sisoB0Qrt+nIb/VHfPrfoC17kxrZb+ksfdK1BJd27o+8entbdwpO
yvwv5J3der4/4q9p7DA2frzf0np6FfOVJAPeQHZXyvgv3Qspw5ls58rHLug7Ae+4
FTWmHQnqxK0J1YyRLXprgRf6WDN8uR6RMap+5fWy1iDU6iYqnsVj4W/mkU7GVcfR
lBiOL7bDWOro43g2nDa/dWsGOWfXv2NgiQJ85mvam0TZyAkJom/ztlqEw7JeBLoM
qyyv6Ae9yFdvLtPOQSmmfOnnF80imDznT/tS71QVivayziNNjSiFvOUoPIm1a4GG
aEFjQq2c0Rsdj+INonMCsqoDSWH+/zhD0QfOpPM9B9vuQuB9lAmtmrQfRsWSokTJ
O27AW6CI5jntK3zuH2VKhSw0x8o/aIf3UjGnJyc8SIddgRi/pfFYFzFKwSHUKq7T
5V8k5sfC2Q6fEhHVE8Sv8OzqowGDSEEyDjqfE330ZjPdmTEU86oNV0x/8n5gj3Ch
TdpiPLZJcGl5N/SANoDHLoPaW8Bl4kGoh7MazOW22kAowNJofKfHjesT9hGf6EP1
8tKnFdJgo72gQFvYryRcqXN8MBNschuYETwKEjU4K2Oxgq4I9LiVPS69A9bj5If4
qxjH6xidV0djTOijwuqZilpF/UgwK08H2iC09Se9cGXyQePo91NLdRXxxKM5XzNF
lQP/Q8IrO8Xdvk21C8Non5nSAAcqM5r46N4eludx62bexA9lucSpHy2q3VvOHBB3
ju3/aDb923SBM+FsybhU1UQih7WE5wJYcmeBrGBMxZcci+kTvQEuOslOwsl5rcVh
vai6y5wvs8HC32w7WzfuantqG6AfswSW9SSeUF+zMLrYcsONI/E79zBThAAiJanP
YfzuC9odA8HWZNvGmrfqPCPu/V2cTp/p2R6oc5+aolOrMqBAaAsEkeIM7oKmyJJd
q2GVMV9ixXyVgQJdsUGSqEYM8UfYjCwPAqAHO9LOIHN6vCAmvO6npVRB2Kbe+7fA
Dhcxpa9XC2VhXqCKJ9mTCz9ec7oCvdzBV31NrC0Yz7YDQXuD6h81vefS7ZhhMnxK
JN1bPnWQxhkn/X3sUH5qTRhduzsfVSL3z1AZfFC9zkVldJO/ilTzB/yeXmhGvcBt
IV3u7kTrc1Ijk80Q6cS51ziz0lUbRYi+kUiUvD8vroa8QKzf+K46o+PxwBD2FQRu
XEDGE1iJRilv1SRrY9cjfr1SBXoTYgqO3/SK+vggonNIeGn8o81PvNmlQf8YHpFb
I+jOf9heQbxapiw1Q5op7mf20LPo/YMWVz1XH4DkWcwDj+qKXGmjuZjcukC7ZXrp
B/KnLc7p27zGI3zD6u8H7RdI8X1yld2OF/pwRp2M4bp2g07l7ltsvvnexR3dTnBL
Xk0dszLRa8JbZGQlBTWVvA458l93G+4ac8KkRF1d1O6RJUuo9OvLwlh3Pxhwla7E
jLCxA2wWB5GGvgtMG8OC5JFreLuNogwOwH0JEj6nntHhfIN1+C6VGdjXQME3bCpM
QEc4BPaeDopOcHyHB3XomEcZV/zy6pJAMnOcdcaDoLl3lbI4cZUmjBrWC4hRgnwD
jK9KAwM3uQ8qI3A7oU9KW0duN8xr+I3lIoIcp9U4lAZ3WnqaSoYCDkKKVpdM4VZR
PVjM14knzjKbNN+/bwWunrpEiOIwbSqmkn3DkqvllhgQbmqb6VCi/RTKAebkkqE9
S3WetQnDDWPlyfWkiXlJAmH7T02BG9gTWDyS+NcsuhCjyfgrZxWGJYhsGjcUsuAW
81eIh1WGG095JLOYJBBKDboSqqY0qZd6AaYngIX/+4SKYmbz73VfH7EvEvBiVVP+
D0YWZTEBMYE7z+bRPFigAtfVZd8SCTfoZdlfnf1HbRnKsah6f0QyP4IyMPqOmue7
JTQJjMlQEhPAbTN4DfxdBOjkVfRcDJBmnJcL3F1jCnpiWWrybVUy0MEs0oecFYzF
9Oc8WgijxiBru3sfITNEKgGotdLpD9MMxBFkCJV8bHOJvq7BF7OOrNhcye38xdFR
EKQTSNNbs3069xwALH/fbd9kEdvzvQEK1wI7GP6Nmi3BwP+pxOVeB6AEewbK/Lvz
3fl3I+GKqAP1JAeAi2tC8mugPyHl12PbtvuUsxxgeSpr71hd7xKHRRzoUVJejfdZ
tGYq1iSqKzWuCsNsntAzQFiYJCMOJ9VpIJuzeP8uM/id9LCcpVUT8XFpUq7t+R9J
I2ysYA6FjGbDFbYtaONyJ+6YN5ceB9SrIYHnjkDMN6JnUEFeb+WW/SMhDN+JyoQW
r4Y1ayJg72q4e1XG6UQjtHAmawR/KQZgUsZMsZM5+9ZZ1vcY+NhlBF0FHgUAuLXf
CusKbVH0NPKtNotUfh4p0IM6+cZf64Mx2i7W3rkVnF4LphuDHBuTGAxd3P3fOgQ+
QfqJf+Jn/GgSdQCGndA6+ZHKsvAW3VayamIj1MkM5oiM2VHUTu9ryHJXRc4hE9fq
zlaM8XaNxTsK8//7QvT/yIyQbUCpbSnUiFCVwJJhG9B7DoR9+HUceEgWRdrkgS/j
TbqoCzAPR617WYiVIqN2UR84mA/w0LpfmhSYePFjWQ5vbslPRhktRtuLVyBW1HNh
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3792 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
yLhC3vSw3ZQMJzW1WqPsUZZMpXHRp9hznpGVOhvQrnSuNmQBCpOhSAqUafBGCJ0B
VK3bckqRdGw2ahCIEA1R/5l1iMSnIZK8YzIUyYwgnvdubJ9cQwhJERQKORaZPDg3
p4xBlVaZNyl28Ph76sBprO03R6nAJKyNhOJSWteA2kkHLtA8OdokEMxUOVfinI/3
DrNtkWaO1TiPBXmA75Ed9MQBYwb3GySXF8aYmN1Qi12FfHEmKdImwPvNfJCobKs6
paYV/mUqJlQbJemcbPRm6q7ALphXZE5YMDTgfNYriiQzmQIwupu3fw2mLswU//aB
mTUpZc2TWIwbXOloh7X0woQwUkRhDQ+jo/YAGlZ0vjqXhIpBCtedJ4kmpUdPLCTi
6T9BboLBu3no6MDokXxMPh0RMcrGWqMUqHVqbyWIt9Wb8hlyPgOXjAuvsRYm5RHR
6pFzFqPrwHfVzW40U7TxNHM0t2FOuk9poOGEqQDy7h7b/utmglqj41lIMDTWrQm7
clX4NB31ngi77DeCegfp4aw03XsNAIiPToH8xuMIqdJ16Bja/fmhV58XxYzb9yL/
4yUCgG4qGUHxjlT1/uIwv5Qd13ol8ux2nkQ2vFgaTaT4aD/6KoOWYNE/shxAMgbK
uem3KErc5FQvzaxC7N4q9oaZAqrKsj1N6mIC53O9bmwY8n5t7Hl/9IoiFejnQKbl
A2XdjkLBxrRnvObxZhR8qT3RvFnLwYdDvy4+ufnuvUVrODq6q1jFElE+NUXtwIlh
V9arZknfsBvt/aY8T8+nsPeOWhMqKonhibrGc5hGph423A1XcsBerDzP2yrIwicZ
KEznkyC5d6jaOHtQPRPEKOqYASBtu8WgjucLnK0gg4EIdtRDU4xXm1tmfvfrjuC4
mkYSdS7WktjZxoiMpYftviOe/RQrs9GK4lPVyzceLVmgcZbFweECmTZH7HFoCkkj
QTrqCuDYLZSK2Z1SU+z9VsqqecKllRwHRm8L+FTfAOsIk0XD9IJTUjjKrIpQ+111
IcQhNrT7EW0FWWg+yFXb7M/r2ziEJYYUKZnmpzcMbxyJIvQdIF0WFW8pJ2C3bd46
hwiTdgTQ8miSxWWQ2NBD3vdusuPyVaLYp4U38x63c1iDxEeYf0ZTefaYqVap0YJ6
Y2oC77vco85skOQpqFiHRG6PFBMY4bml4KI+KqJWuQr9VSvX2pvc89uNoSkadeK+
eBSiMReXMAoweuwqcJqI+oaFpEsFVgPS3mrad4tSD5SBl3yVLTEtoBAx+5GLeav6
1AkidiTOgSj5qFPLWbctHUI8SKCgaiCYCforBSsDwlaUpCfXBlwFVQQbFHqJPFEU
Nqg/uaJQXsrZMMgP/YDD62n8VuBI8x30DK+ffXYQ4S6kY8+f7Lpnw0g44li8T78N
hqzuMVKkWv4+CwHfQzaissfq3fX7oQLq5uxguD2Te8AqU3g0L8mPJrIdPrqmsDLP
7JTyQffH1tmEQETr3YsfKClOIisd53A3SGShJJL0UXLLbxCtEAtoCHBBLWOgZpfQ
YZ9xqvHm4ecF7LfMLCwK7hJE8BVMVnmaC3LGWqFf7vXF1e7LW2VQWNiC/0uly0cw
KxyZYJiGUBl4LeL4kp0ywOa4JnRpRuhC/QUk0c6tw29le4s+gjpayG76lC9x1gGE
Yar3X2QGW9dL4Oj918OVC/UkQr8cHN8losQIsaW/GW6hjwLjpqKbGkIZItRxuJRD
40hLZVEiYwyiZWZbBe7zNvXAckevNGr3wgPQjgUS6XXpcIGiNgCsPxsWyIWcxAp1
fBYAZseWZpQshyJCY/m///+Gv+3045wIju7M7bo20IK1Q5aEsdPYtKHszaiQ0r36
TDVCN4YEoaIjF0DiI3T817XmR8Z2x2mUwQdfKjLr3/B5XWc/PrA8gpylnXpypaPi
wOhPgTChuMx32CDXLt4uwfAU44wZ0ILykfI8mGdOWNyY673F71JDzvVqZGM+ABFL
Idi90Wirpg6x4a1bS4V/0sUI2N8P69FCQ8fWcAPs481Px/EIevae0dp0kYi9+u57
FVdlZ+LkzuWDVxlF7wnmL7YPnz0ju24Plw1pNAIQpd2C+VhHScCr3li5zB2b6sIa
kQ9hM8MOldduLpwo7Hm0b5thzlC9mazS/bUTFtd12wprCi9WY0Ej9PMLB+p15YOE
wOVtN30gzpq4MdJzu5nywrOQ5uuxP1FgBQbEF9/DCDD8v3xXV9J8KPaYZS22lVmI
ql6CTEW7GeQFk9eKabRz/vWDMH2SD9QQjxuKl+EoqCoxjFRsi3Fbbc2OzbFx+Yf9
aAZ4xJbe4Yv3fpoVndZlUYk08xGBdkvgg3yITHV8xce3dJC9f+3ZmMADYyaqD+iI
PClUpj4SaHHdRpYcWDuWPLM7KHK51wwlnoWqgJAZpM7y5v8rNiQGLwaomv822kp0
3U4eY5nqMb/9uPjXfN9wfpnKdq11SwrxlBFRcQ2x+TY37qvUrqxnhqr3uxwSewUA
LU1VKvGIGyt60rtiyLGcUmN6pA1Wm7vvhJimF1thyOdhK+DXQFO4YVqLrvc9onkS
V7xid1gRv4rscRVYbB6uggl8bBWYYVgh1qDpmMGSrkX7mz6IWWBROH3bLjy5rRSC
gmEaeaOXLDpShJ8uD3ufx+/apWvxW2oqJyTFRX8ErPusyOFSY9ueZ0Fv6Yoljke1
aaCgVEKFyXmN8jEmZ0jpMFjJINoY7VJJqohvtGaqXVxHNiOnuBtxN+IZEcylnwqT
5GRJVkJ2MmbkXb5B8ayZwm2cUMoABP8n1fwpZDigA8M9o8wD9L0FM/fOWXBJ5zN/
gEZFsfrKlGvp6Xu2HTc9RLnnh7xSqq3Hx51LhYSD8/N7f7znpeOHLHL07wsGjATD
8FWzxYPqFQGoxHwViSDug+gbkipYDB8cXjHuinO1XZ6rE8H/wzwmWxVoizY7U4dY
bzcX38BUPTlvlJHCuBhqTHAU5HPQs6BOYPC7fiRB6DJi8mgp9Pp4RY9GBY9bwAuD
v9zdgmTbqSc1GrsIx3k9Y8N86ShM2oditjoEo7vXmvvmPwyPYa3JED6CqhLHhZLS
Q/n0jscctaFmsmmvoQ6o9RoA24P1m0dYRAaPz464v1YOlGH6T407u2MLHZFS/Bzs
owBUeY2IMR0pbpgM3tv15WwKduZg3W846YhgU/di61Mo2uC5GK0tmlfJ2oIZGQcz
jhKRl5dPmFX6wYdGm+VuCPLFWQLNehIjeOWs9zfiK8VgZ5NQDzc1oKzTzAk9RK9X
qzRycSPq64bJXdb3sLX8gjNSVdpAARZ9Nr0zuT5HDSR66KFIBOaGucSYKYzJ8Et9
Hz/mW0HmoiOl+QdiyDS4T8ccSVzOJ42MioyA4YMtA3A8EvMLeNhPoWkhtk2157yz
iDG9i+3EHVXZX6stpVorbYmzayL1xKKhc5Xk4zv+l1nIUpJ6hd1/CQrH4bOjI1eE
tIjNHdW6Oqsq715S9A/ionJnzniZCq97/JuEzyEdEa9TgmD/HBLRsvW/Y3gQJocF
uih0D8NIIqFQB6ziwnuDOUSwE3DQYS7JHsgBtqkz0anCb9tKjDayOkzUDQJ3CV6n
ku5SXlwODhmu3t9wPtBeOa1VhmjPbk9QvMxBLRwVeXr0/jGq+wBxxke28gThSIkA
JZ3lXBJC7hoOpxcPwfP+P+KW2A38bDZVATc8gDFlTe8lE/BEZBWTqLtkmlAb1uI3
FekM7vvQjEu5CvmT5bV468TxSdPNa+vl3fTYL6//vNEnzlJ7X/nFnAOIt3Dr57o2
JEsqNVycOFK9ZEoablegPHi0aS8H1A/dhsFQFDpmEmufDd8M16EaSsyrpjuvJRsv
Rhj+5TguUsJNC6hnvd9sGkg2tD/oJdhHkjqt21UjONix8WgRrfhtNBfZ6ejwFwqN
bAjr+htiQeHgC/ar7eTAF5QJOL4qVOUNYOk360X2GpkrmzCE5ZHRyPSQVu7uCi5l
UjYXbavgN4a1HGAr6tjS60sniLB+XIjVdffn2cBNL4WfLo3CERn5KJMijaQ3frRC
tmWA7DSYXzKCic/lM2lX5R3FPL5wzhqxbT5huTXCvxfTnWKCV2qpSei9i8puK+1K
LYyRfy++khGHL+WWjmVK+zpGsf/7sPNDrTc63zQNzVbxnh+wIp/SQ737EuKFrIgk
YcVOppX0q9vUURsZawIWjZW1DOC0eQeY/stAAKyyTtWZi+mud+VSRVxStf7QwLCd
pwBudPW0cq2hMDFYoKJJTRoTh81/YEj16BGlofCrZ94fwtmYWT5lqQ7/CL3z261v
lf+jinvnG3VfA4iGZ2nakGLeTA335DYO09mnAvhYENJCDHKfAsKYE8Tn1Zp/GpPu
bHrNez3CA7iG12fZVAUxS4oREGnFljYaEa7YKT/E34awTuERIi+k/N4a8g3gkbnn
BmJ2QDkWY0Y75b3NBY4jZbRQ477d4e/FwDCYndDNR1epIA8ZdTIvPYIekrQcUB+l
Bs78tKhlTFi93tusDYHFwhGadyeeWLdiN+z0wNbd2cOH84LgF+NY2vzwYxzLqXR9
cTAnFob7T0Jl6L3Mztiw96oGbPaZvcKN5Uk/+GkW7CcmvmywETDphh9Q/tKv3pDD
rT06DQJA/tJhXqLeWrYwBCFUbtGr3vC0eLUslQbCh5nwop7Qn/DBWEfDQQuEo4H/
Xj8A7ONBtLEmcjcY0hWmzEgZw4bydJFeFOwdQKzY1Ci+5sKzZ9fidPn+xQ4wbcK0
9srf/XbWR2ofkjuB3qPZGRtCgLs4Cx2aTlpzUys2gc8rl5QgJZX8t9N56iOtVv3j
n9UTAyq6HClZCbyfUOFg/NFbZqTJHriFHSvyRPbyRoPIVurATd23aY0IYfNI/svt
fiZpuWBkwX+GCDUHjyVivH5W1mI96CoDyYDJGg0F5WrpKcpA17LpLjvLg1sCBBYm
>>>>>>> main
`protect end_protected