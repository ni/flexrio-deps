`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 34752 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
EmxAgecO7UDIr+OXKjjkXABqalBXxig/8b5H9JahKJZ8xg+aG7DHwCQSQ9Hj4UHL
PXVEDKTBhOS5YJAmfJ2iDDCo4bIyfa1I7zu9YEVO7WvfATymbHLBGUAIb9IC7vsV
QvjdEcG0mGPyLdG8b38X8VTwqMIGxPE+6U/yO4k1eOm6PCviNB5+Adf+wfd16R3N
Yk9CDpoku/P3HwLxyZ6vxw0J3Vtj4pYX3IT41UQcUwRglFCdrNgTG6nSbbWa0XeL
k1kdCGjcHtgpm7UszvpHy/DkLzgH7QLPx5YfkEE8qvjXRRl2sLrdQL6c+cfSZeDC
ZleTTE6Q2jIJ9QAW/djmw55sT8Jn4fxpNw/7zgiq4rzxr4BOPOHV7WddDHKt21Ov
ZRN3l5J5zPkhc0KrBapN0DwN5MB34wZxAJJidgfi7JQNe4iXdI0mJbCttJFmneX+
rKDfg8SC5yQR2oS/r9+rwvcA/4vG4kLbUfuC4Je/QFWTcIO9tgoMBHM5+80wbFYQ
7/NNOCznea27hFKXha5h5aU8LMbvX1bPF+uuYPP+Tgnhp1z8pvz7crrjg+0L/wZu
x/jsFqoBqhnQg/g3/FZQisGb82PMkXRhqZWED4G+nQW1I4X6pKWz7frioiiXmAll
4HXUNsm5u9byJhHN8jHrCzoJoFPuaNcBI0EPBjPSdL6ve/u4JsrwD0fZwDKGgXvw
KoxQGGpXMWyJu103ru8D9MNrJ30VViTfN9fGD/5O9dVfNVujnEOsqRaxOVaSgD1T
05uy+f78zHgm4oCoEhhp/GZomIP647oMl9h4anVz4/WFca1noAHoxuEsIEcqiXhf
7LSPRYGLSgYQ+Khen69kHP4Nesj5suxrwondlfCr22ouWYzcYAjPJYzdKzR5jdOs
vE5aSMTZ5sT5DUAXm7ol0kDdVMkF1XqDGPiv/6wEFmkNrDL4amuwqAJ8GUcYMcor
yFLsBn+MKgmT/j9imsQjFW+6dLo2ieXHRszWZYZt5GW5hpt0ksRqvHsXZ701cv75
wqmJWN3opAEHxll8cM9rWlayg4HYRpNwibgGsIprYGkDgzMsZ3wovGaMLgtEN+GN
S/y2GIqeqhHq0YUur69qqmpBdvw92AuPtu/1KU3eGmLUbND8ZP0ZfZEztlSTVfHD
fLdnaHunstLRnP0vfC3KirjxshMuzdzDJDszXV0nK1GsHhLVlAhUmxsA9FvgmsFI
o/AmDggWtgjNnJ/ZYlZmT1LZbHTPmB9Ou0Hzbz1Oih74KVvrfoMhVA9K1glaxD/r
tLynSmLbeSKNuxp6jTy3lnda9/kMM0BT0iYObiOr6QdkP9aGqigGOnN8jkh2Bz4s
eNzUvMyisTMs/ROEbHRmMdvGgrwlBOl4dSXD707GTzI6hxl/wX3YXXkPjUEuzwSX
OicSPAEu6RTmjRIjDp6HD42fz+x9zDZX4yI6Hah/775zzHt+0qB3q6OiYtkdrUyy
q9Ic4LdZbGy2EoTu/Kjx2mLWZGShny3YBvbOkS3HhHdac7SnGR6JCdyVUER4QjXo
gNYAGkRtkPiAoI2RYCq3dvyoduc3sVZLkGoNP/TesCTTd3dN8HAtGdH0BAbo1LpX
5/234MrA3NTfJM7cB/NzU69BhJp5tKaFnWx3ngYhraqXWjVgDBQ3T3wnb31aEeHa
Ibh67m2ssqgf87BV1eW+13ES/55gFs0VuLtxV1ru6TUMRqMzELaXpTxTjtODFMmm
GvlKNcKo+zkVb/JtvqoNKG37lJyOA52agIQF5hSjhxvy2v3+LLEs+Fj7y1PoY0g5
v94Li/xJTlNmJqp1Nq06YHoSA2PLLY/oz3b8dpJFXTVFIjCJZ2f0HUDgYSbkaQ+E
5QuJ0+WOMs57jEFTAPt4+Ircwjy7xdMYVrqoRcdynYOGNV7T0XGG7G3kLZJBG3bZ
XTLc3l6/VPPrhZVgbqrNVY2ewVzsSLx9RXjwXIZaaih1Ax5HTBUkQBUdjpus/UjA
lIwvm87/ZTxzogLjUJssVQqtaTRiz/XBwNzRjTHI89hf+HVz1zoi7n9RF3OU380z
TZ7a/Jrkxhnb3awIxdaj7qCZRwZWol8VLbhwbBmcyvy4jrKqKepK8BxRpNpCEfzd
XfYYWh2WaRQfKixV2WWq2CtmSh4xvkqTPZm5Eu/uLHKLecRQXEJSLCcTMQ03VRIr
dKY30Q+z/YOK01VNM+C9w3TgnQItqwOSgSF/Y1ugZUEaUhPJcp9Vw3jSMhcvTeAN
PrYsithc624+hbpfYhZivPop6aNxpyW7M2s8F4kuVhndQRNvniMtAjnov+6mZoG/
JnKt3TbldxEXdcVxL0Y5cR/jK+Bb2wcKeRHJCFcUAdHx7xc2RoiBvZBNABAnwvvj
lWj+ypngEqoij8C2e/U8B4ZUhE6FXYWnesMTmdCcrG6iKECzilGF43QXvA8k2w0T
XkDCJWMWGZfED+3ChTrDOxGN4qz3KRE5PfjxeuQsqXCMZ4vJ/N1w7NIhFuauphMe
zd9Mu5hWOdohl8MZnB0MPzsGiUx0x2KxIqqZWHuYOLN7tnaVQ2kgzBQmFwAedKUq
iWuPI9lIkKPTyQUBTjGtcG66gF5JNHG6GNa0gA+IS6WiPa0TCVar0Qigoe6yjmzW
OelifIv3+iIMEuIljqWHAGvKciyPxSxW6LeSoCLY6CxqUcE9HDyKOYyTctNUiCNn
V8UbRqzYTVKPrOym7TbGhB0SEWJE0+AjPz1kzSL/vuX/gVN1SiDAiwYyNx0ki6vL
XB8M/CYG5D0wlXID7SbzWE6OXIY03eYI8HAbjdBmH+5ScU2ty50Q3diSIsf8zF+1
8GWIUEo5nISVBjlcqUEF9tqLCHOFURXxHsTVb8k3IpfFMKOr4InLxBIHhKXnGVFa
uDBJBpZdIfcAjssS/iOacDnNUsTMFII03LzjmRb7UavWRq8ibqs+HrD6duzab4AR
ivKJR3q64SmeL5Gu3kQYQCeaTJ9D6OIP3xQuIgRLM2hy0dDqcaYKy7b+OpO8TYze
WDWlw8LVasiXWJQSQ+LwRw4V41wYzzeMUnd4rpE+Vwglzixalx2QkoH//vG+xWFA
ZXr3ldgXArucrudh2blOO2Z25npbmZkfmnsMLJRnY5yn9/a9HBknxdNyh05c8fAl
s7xb9gsf3+5C2Py5MSaCHvyD8DcVhmsKbuUK6XqOXTiXfU9NkuMuKnLGvJ+354q7
DErvix9o1UnbQcZgL+P39sVaHHGpjzBythVPJoT97H6ODNtSwNCM7z3BJZNdf40b
AoKDJr9QgYrJchxf+RyxuUGFbjdp0KxozhkT5MSQjZfNvXeyOVsEelvgLPChxbYO
CVHm04NfxKCBqoe4dDyiXa9pjZpQ/iKHP4xNWbHW2okxn07pPRDr63KpZRwBJ8Zt
zxpSZC+lCmpyPVoFKOltDuCTOhyUGQX0sfovMX3yIyfPpU4LWl2vqQ5a9ZWN8yLZ
ucb/Q9p3TKloowK5UMHWpGi8fj+3m7UckCTScpnNmNknIjQJNNMDm8Gxp+WwZiP5
v8WlHlzQutCEkFwTuDiSJfIGMMn4fMRZI5uoU0vczSqRdLKZWdFyoMsqi6IQA0Rv
gRGy0ItiROd4Y40hydP58aDmDge9dLgfzKerpVS/uiiJF1Mt7Xsgd/NjlEOXkxmv
hKFRsRkWKr0c7YAklLn89HrknrlOTRxC5oIVePEQOxi99eRU5pOYlwaSTv2B0aHw
ErI7pKo2xqXTUJYGQEKhW0anIB4uonUCAVr1W/xROozjXmPmnr0Qgvd9LI+ua9Nj
kilzFo5f5vvZfF1BMqeYBAN5ao2Xiam8gCy2e0krsK9ULV8voEr/nZzv+2ZW5zsJ
vXrcukBYy+TVaQ9WfEDQbrYJcYUkSx5T5L2n61X+Ot66Wf0aqACCsGWShScyYCrO
AFGX8Ei7t93+aTslAU0il2sHrcIBsotFsZUiGcxLsh0uKSQ/ux5yPXdvnRBYm8NB
H4gn0wQWBmhDEuDSvCysL80D8h+/elsh4Kspvr4b6yTCudKmdms5LRbqFhk0MBRP
03E6X37VPapSSE3MDf2ZxYxasI9GdRaZ73O8Opmnuj9yHtY6QmABen8y8Z/nvva8
wQ3LmKBzhfc+9Zann70LakgTxXNsOk6oWpER1XrW9HXf5oN40RsD8flFEoBzsXgu
ZVp8xJXz5NarJ/pnU6XvM0mQPdoMZoMTzHZEBtFAgJ+b3CM9ykWQHF/J9txZAf8B
Vc56BmVD8c9E1UmBoCYEV5tYydpmAK3BF7UXixoWyMuZiLhxzjGmLwes4JKvYOex
3dRrKh2fNaTDpRT7YNWIf35tR9ug+q9qUt4tyWzQ64wWohGpRZ+b1vfp/LDBDuyW
xKNehGM6qzMduvsjW2NN8FVjGv0hv0ZFmohSfF6rMR642jFp4R+hUBaddIL00Yma
gIZ3HHbfce6gPh7TyerugO5/MmKMN+wG09Zwmn8eVfsLjhTxJzJaJ3wGEJr+xOjt
1E4a+Ga9bAGEOTuJleFvFHzOIYhoEkSIPsk4fzbI/PWpuTWx5Z6peBwYmTcxBN0T
/d921oxNAyhzHiiOFXYR9LDxweHhP1z8y8coF8HAcNRML4Bch0FrhHfhrveIyGjT
QzWuV5G4njS2LdMTedQF67+zAO5N+rW36QoGTPefjuqNSLhQCJ5aEix2Wy5/I4lb
FSEByQhkAWd/Q19hB+N/EUIanSeK5vhu+6vZMcx5Gf7F8PY91Lk2VrLDacVQcL98
AnQZX9Z5Wb6vYowfIIcb+GaPs8IulvPZjGcViK2vMZnK6n2cFDaVPrbJFzGMpfS+
M68Dj26vUUGfJwEUxHPxgBneF9gEKYdV27sRu8toy1DKkjh2TG7wIA+it7fJGHR5
w9xg0tR1VcHYfETpqTgbvbImS/tfdmG3wHbcznFILF6t0nmMFrQY1GOQLWSS1it1
vYU8lXeQb5t+ARWLer3kS/T0m/K7eKItQu5K3kQhVVoo42ylpy2pJBxy+Jv8DqbT
IvNCUBOLs3/xhqxicTX6beJrqx1nSN8qhzImg3ppw5YIKcfBcrNG+PiiXVKX9jZ8
AI2TKYWg3dtpF5onASp+sqTfo+Z/3Bo0csniBee7FFTadh9+S3wvVAGhri2tXeuA
iFZetob/9jK4q3WgAHsZ8rpKC9kDrbnrzpWgGdeeBba7OUKj07ucp7tBCsgSX+aH
y4qxJgjYUQKwwPMk6nDaY3LEXpZ3LlVVw7ejGetyMSEeApwKUgzjPn66FgSQ0NcP
a6QTpY69R79iZoLMkEH/wA1YQG9970eb5mTZMW8mXImc2g1QaMpvtbQcezgrRAts
vbIPS8VzKDE56PMH9+eOh84lA0mWWgE/j06g4ujqwif/pZRbgTUpSzYFlU5XzTQM
K4QkCR8h+yFQKtxRq7pnadp3d67QuK7VOKDj6kAF3JVIXEFCGsvwew0IYPeIpw2u
6IQrKcH6y2XOdUoJa/DWMLx+rNhixcD6X3uMGkmb69O/+3zEDaT6zXKw9ZfRlYid
3JYfQZiESTdaVlJTLuYxCeP9L9+socxrsh/IFSSMAPqWM1yg5M7EMN7s0eNn8TK+
+f+e4eVOAuAzulFn57O5LiNdkfp2ZwsDam43FsRi2eU7qRTsLa6oHgmqgHwkze2p
qNmLXMLt1fdryZAZKLdyGDWo3iUoeAHaLhkdtDsQvDlb6vvlgNyW0aE7aosdh907
SEFfdCMsE2oINNLKrQxjEQ43zmPsFREHDSvIw8ZhrDXA1wfrFVPQQzAzKaSPYsU4
yMLOX0/wwc9A+pMajNIilHKmAaYJkSedLnmVnfwma0SrMIL2aCNQScP/IuC0OBua
JapEGDP6/l4eVPnhWNILQWztm8c4sG/ffellDR/bKItkdPdLn/UrUhk9uQ2Vt/aG
3oM0DY5Ha0g77/KsQn5K0Ham8SWzLSnSDLsCAYgnpjivc7VXlZG/Lw03vL9vBbj3
x/GRSdqAUZnNDg4sS4o1iHuYPITF3BeKhYD/KpUo8fkCQ7T6mKBrlUejG5l30swR
BDdRCyqonZmnRKCE2/hcrX+AGAZnTYgxLCl0Z1XGkyX+ODWK0qI+boVIO4MOembo
ueGoXwdV/TolmVrN4WCDXgNvvwH+z6bE2ycBCYHUFwM6f7c5kMmWB1LlyxLfrSYu
BXT1JrlkV8B4hG5MoNHPmfadQPzeNhect2cC8acmL9HCb54aInoSBhPOr87+akQI
Q4fwIcfuoSaHu9HBq/0Pn+2Z3VvGpPPtiiA7sB5QqlKhCGIi2JB4YO2hKaFHEipu
9VQFgokDWSpFBpIUZQQby6pP2PLdINDzxMN3wjPLM83q57D/1WDt+hQuVLVqkyH8
oZUPQHbwZ5e17OK4+dKrlQNxgkW0DX06QW/vi8/G7XmKDhJN0dCwLtTPvT+dSxBe
YOZLPWRMSb6p2f2us+eQ7g9G0FTDIKiB6g2SQ0G0eW6v57mCPb29yiEwJlDtoq2k
5Sw4ozhZGs3oswc77Z+fH2jkdJgOw666Cnq17dnN+KUNpJBEzpwmzKbrNMzeW7XQ
z4gQwMODo9lVhk374fF13r3ydbN7PQNpR05Fcg0rJo2rjynHK6bH/v/4ZYK3YiqX
17BzkEJIcMW2jqkFRNZ6XqiEQ71ZrjEnIMxZiLZLbMxndPqO4xRO7fj0ZiQWz8lM
VmVlEi4ck5OOcIFhllZN6JsQsFcFnLh7anXLbCYEkYp3FidXREA5IfBOe0XITqEV
wQZ2aklDN9BuubnmkUOwJnKKccNSmtD9DraBY/XwQMb8SZ7cCXpywXtWyhQJOSoK
VUtbV2nTSFER/XwxvUAtXYVI/0Skvc0gjr4qK6XnK8+PvxfmzamHKplfVOpyB7/d
8SyH0cy3KL0qoMiOPTEymxS3vdEXu4JxTPXt0SVr56ntrwmqps0nwwI7onzCy3dt
UAU7nnykwQ08uWAFy6nrrb2whu6UtQG+RvuUJFPBV8G8Nk3vccWLtk6CGLjjkezH
wgl1agu2AHa3qY0SJdTOiQNI0jk98cTnHuN4vhg7heh21bjjNBGHP8noX/mz7S26
0mMV52ynDVjVz12mtbj9jGAOq5Z6drJoZf5ccbBryc9vzDuc53twSaBXbu0jICuP
QYhJ/CIxGObtJ7TkIa0N4328KRVlFFpFSxzznYgjkFvaJ9kh6rax0tAumqok+Ut0
qhPf/iTCaV5Lisn5+ryaMfqQ4UmkDdJexGHehZbLoJoP30XvtasBEgYiUqr7qC/0
NpoIXm5L5NPG6+6uzRfuBs0BIAzfu8GAQYRvYtqGRjCuVJ1YngmxTOQo5DDu8i5k
LCwA8oSHeTjfarG0sqWlSQgrKMDqzfSzTrvwroj/LstL3btWcUKktT+TALRj5rE1
yXa9ClYR+plQg/nbReyASGbJckgdMSbIBGVF8WP4OQPIsV8tSnjfAuB2eGTae93r
Uh38PHN3i1T7VuJ0Ubrnp87FOQsn9YjPcw4CObKVh/lNVcIxZDr0b4WythLK66oc
/RBXklBGxWkRcmISXSTBo/V8uNmF1y+y5h91hSxpQSUGPR7sghJY4ic1zMiVqc5B
04TZNx/F7cjnHVFpT2RZmQ8TKaDCHwZJjoNGjZUdz2XcaS6qkOY4ffnbvdsfSRRn
7/fMVNEhVSjx3dgAvzTa5sRxisSVBRGb2eJ1lhUCJOmReXyXtgwJAo+5e/kPlNbo
+P3OnzFHjWoQ0KGcd1J8RbEPbpvvwhmoYPgCj+4iHHXOGGtfHRERRyuK927lbrds
MCCNjqXayaQr7qFewJqyqzimEdBFEuaQaDqfGEikcLvCU4/dpAjONQHgAEmuzDa+
2FAQgrlxYH/zFAIHKKKVbJZB71c97t6KIpTcPX9h0sRgdkD67fSVzSzA3m0CaR2N
W1PWciWRPEIdwSokvgGb/qr4iJOMs8PJagORvV6fBPQv8Pdre/nr6bc232VQfHE4
37nMRLth/6Xoz0mVaFt9RwKycHIZOx3vFoTn4wlYD4DN3uWmIe+Ilct2/tJCcnah
Syx374i8SAwPdkgSY6cHPAfQGKTIqq8GYndU5dbaOQEn3TPljtK7exo0h9DtOhRQ
XBZT/YL9HKMm1k0BdXliHnBadGbwNMp8QQSok31PclsCMyKltePUT+SZ3e6af9xi
g1lkpWtb+RzKwHFqRybXQAzwheel+vKiHBA2WdhxZKni3CXAe7q3qDlVCRUNweX5
ydE3q6gr1PEiHKfR7BzzhiJC7urGOACpVBIw126M8VRFoVWkGvOYE3pyepLYEGtR
kcHy4LZSL+k/ppo1a2otj2u53atxziqN0ze0nD3GSjjKNf3PtVghXaJ1q8R+/Y0M
FujimmNFckADKErvrq7r7fU5b7IxiosVcV0Mj3Efiug5tVcnFRbf/09PkzcTIq/1
srxMweGVj/bY1wj9r9+NuJx5jQYLODXYFu5vfpQr26rjMf8NGNP42RyQaC/VeFfA
VMMHFlYbSHO7IadhDGHcQ8mY6mxmPTIOAQDQ93XJB6f2QSTlEqN5Wyc0ewXqktr0
YMtLaPllvY7TZF0iazsgo1yMtZ2p6arGLzmvnrwLHBc2TEH4ZYrJbtAq7wlAqDek
WcGf7FTjI+QbkmFuX5ic+IpWgL/e9JTgrqdCg+2nXjIYgymzfrxJRKke30w0XApp
AaSpyxkAJyE/vV9lFsN+u5jl7t9dudQZsylOQM6E0tjzhVa908n836i/4txNImbK
NrOSFlSwr597dfOHBtyUoYDxWvyJtGAwqCuOaIPmWSXxyYxt2Cd5+1kKwgb9i5uY
vqHPDe5sB+4HIMy6DsiBYgUUTko8umOoOoKO8WwSiU28QpZF8Bh4e9G659CkzezV
QupduCD2uiJpJZGgig1RJTvcsLAOeRvnzCB2Zix1dCbC575354KH+wHnaoZoVdCU
IB+HN68CCwvBKa3Nsz2TRhotg/hAwrtwFrIprFfe1FQ0YbXy6M+eud8uQ3u0QMah
Tm7UqD6dWkkrScCcg4uNAFK4JVqDkzM0WO80imavoYe1l7Gk0VIRaNfas63kCeC5
9iP8v0qGozBnceg3bYkA6sRiO2gstR5yLJYmXi0Ng2wol1AvHObxh46ualBgpkpd
deytcc2w6jkP1KYVyrIn3YrZCP7v+PxyFUU+7jhfHXfStPE1RLKLVa8MjngQgtds
nWjYLmGLHeqjfzIj7LbvehZGjeSGfY4mkXmm41wGqJpu/XRa55YvEGpLFv/2eee6
DpwSAEBklQinxcxGfGBEkuB67j4NSwa6ayEhKG0PmBPAzih03KXGuj+JDAgU84zn
ZRi9kafvUuAjesadYI/1nn1apDBuTYu35kVnp5I0tubY4bHBYV120Gqi8BPilGaB
Xnx8hq9kZ1RjF8ABKFOV9IkYvAd4AeMNx8Wlfi0BtXqd0Zr0fLom2Fivkd7Lwa7m
bgaupHUvzFoUJ2kvEdy4lQckKmHPI+Udz/mLzciOvqY3neSYiZp1HRm5Bx9QsfB4
kvPd/EizIXQhKmVZbChYvCrFD+IwKuQl4GzND4rkfybqL0MFtB/sX4i6ztOc52Yu
pLqGYMT2+ITFwupv2/2qglBLn9pn2qAU7owBCQFszglgrHKlRdzCc7kS9KyfwiQn
mOMNk/0cU6FUDCROSKgp3vkmEALz3Fr8DPHHcsp0RVRbwZBUAPmrx93i4XGV1Vpx
t2y+EnUdF8T6t0Esoxx1I5pl9Dozv9Nc+8ucW4WTvdVz44IRgBDZxXlnmfqW5L/r
Pn+3gbLreUzYYnGOH/cl3vVvX5i5aS7GyX5AepWLnE8mS49fQIE5jnB3m5huTEzh
/peJTjxzqzOslX2EiRW0yp7pvpIzzRA4+PGoq68gK5t3thRb3l3+tdk3fIQnrhox
Jnv58J52s+EeV2pHc05HoHftoT4rRb0chTAeMq2pl1dkaVk+WcuC4CnUPOATdfz4
MruYCqOPUeLdEBXhipvMcHPOEiU/RY16XmK28AvR0Yi90pKwZQeioHrbSfy1N0VN
XrNfxru9QisPNyHn7Hgc4UcAGixqtbqOM1ZSueW/1OP5iRX86OORgZMF/uge/uaI
EOVzW75dg1xTcfXYiVvEU+ZaxkTkMQk1Bl5BM0izvNGMSN4mHuGwfofkDiy/IrGY
VdAgMEJ+VZJOeRggaw0zxJ/IitZ5JKOnnx2UP2QU2evATA0sDK6ghud/dAljoqNj
7zC9FIn0JSblxIh2slMAY50jndcVK1PmY6NUZzobUWrToTFdc8yveiUSvtkg5jNv
dlv7O8scc5Euu/9JgFVsHHcsBiiUr57IrtR3MJCEsS/DrjxTypLhci+f1jYhIVzo
8yrew4AdTQmSlahgYJigVllDZhlW52sjmYRY2MenenlyYAKNrDX0mj8tiVW+ubI7
E6m2T28UhqdRySVQgp5MGw06AnpjoXF7tTETQELPNmNpzqKZOQKsX90RajCh483Y
XWkJfzuh5nDP5S6C6pcGg6l66COpua+EygRznmsiJCoG39QvHhC5V4YVX62e7c2V
gHXU3Hwayi8zBI9uHgKxnK9QquRA85yHZKlqbrpcMIiYfaz69CRyxAVPeU9SCroa
BkqWO8gbcZTYYs+8BeMhw7AqYgQmlc8z1UsE8C5/Ok2ovh7vAxFJF1x20MaJdU9C
nFZW+SrCrJ/5mYwjK0NycBm/JudeeuVjn95Wugdb6wg3sz8IXu5ShGliHzmfK7b3
1DBzD6/tA0j3khXOQRW/2TSua+Z9AzE+Wp+IkfDLVisbeW4im9goPs+Rt15Uou78
K2zNS/iIM2VaJXt8Eu0GdkGnT6Bd385KmiLvnM3w5PFtHUFN+HCmPyjJ8KpgtxIE
rBuj96zFkecvuFnOMptCd1Ue9cOa+BAunYgYXNm/3R7U8KdA/cJVuZKXgwFySZat
slKhbCFJgzmos5EMwJZ89X5SfYJ7PVMjwT0eI2aYkMpvXAH9n0gCTk/KiPWpUlZp
/LrTMvMJftzQsBkGVMKg0SNfJmseFBE6E8SNHyVtrljYm/zALH9hu6AWq7+Zej7k
lvYFj50s7BonkrpzbIcxvc4EyMRoQB0fEIWkkOz0wddqoPFI4FRgWvqHN0WNrP68
60R+7WV8yl2A3iH7uFZSjzBz6865DdASUA5YO1mK7XHCV8l+vhJEjS1n6Mh67wMx
fhG5nxWNGZ964wWiTf/rIUgLTLiYw/R1htGVza5PU+N3Li8MNiiQ9oMIfH72VN4e
WRF/RlnuU5QV4/JV7n9o3VdSO6un5Ly9DOrERyk0N3K9BzaaMreG5v6wg9lRORVe
dAG6SCcpcHks1u/t7YDyxiM4/Pvb2ZnM7Xbk15QC+QaeSBlMVRmoZ+y7YnW1SQB5
4LWg8+QZUWVrzuBMR870dv55Vwr1ycQDTSZQuG0kBkOxTkBBEY0lt8mR7MneZBax
axRYN+qbOSjMBhUFTd0NR9X1kPEQNIH8/yxQX3/Dv3HPXUUW/LBG61X0aa5PNkFn
qUFLwfYkdb4Mqkf7SOOJnhYdLMRLo72MTyfZCX9rntvofdcviyrtg63prc8mdvKb
xfPIrVM5V53tZcoAI5vQEJcMN5bH6ybJ5YrnAJl28M9zOn0QIHiGxtsAxf9vY88V
Kt9+yNPYdrrmjiJryU/dgH1gxBnIzGkxNGv5VyQz95P5j+xHm1tFrhYiIzu797P6
rnup0L1L/cMfiG6OurxPrAmXVkiXhBhk04QFYUIyic1U2Zb0chCXmzIGM54EZsVm
LcNjzpSSoiepMW/n3fbdk9dZcspA2tzB6/6XGc6udXxXy0anS2CBLvZRXVfKhdsh
ZZpamm54LZ9iCxyCtNbgAOErOwnbisZtpruoeQ4p1+rUuP4AcscjrBaFrHnLPa7a
TVyGgbVkoQEnGu7/lI/VjjtCAK9dETexxLILF81N25Dl2q8f4wN+pTohUM8hUaFE
ENU+ABtPWctkrLJzNzbZyw083dKiMiC+ScfgkGOEVRgJI77bjWYi4wZYJQeAffBc
MV0Ft/6M1xmaD5Ybm+nWTfrL+WBKrYnw5deV44Rhb6GolBK4slTDvSxDmVERLGN/
ZRBdHbO/38i7iHPhDRXeprfqbV33F9mjBwbgtrqVsPnP0sotWx/1fjSR7qGFUof6
qKSP4WIJ6TGTLA5h6cpBkMGHk+HMIOdCZEInNgUmmBXcaPPjU0iRgE4IHQlbGvD7
NcvAhYS11p2LuRFaMvsAqsBo7n5ORRFIRxG0GnFMwSeoXwvzDvrO29K5n4tANT9B
1dDIBcwt9IKGCBNx8WmqUmXSjq8M8X4e0w4CfdxQgaU50vsDADvh7EWBuUBKF0ca
RAzllY/szbGUQbiavJsE9lmGjpM07kz26+Tj1ZEbET+7EYkZ6q3Prg7MNQCy2AlY
2BOUovCKMghM/fRWeoeof8SThAACi+BDgukSBuN5R7EsnbRVL40E+nFL3Wia9KM0
s0VU+azGmeX31cr5Tj9jAlvz7rGvSreyskadiHr/KtH6EfPPGs5TfHe+dJ5X0zIX
DwDD3qoqb0FakfTVMYrogTSjcivjCmquIpQtiuucSUqcrWWIVZ2qvuEOavuLj+S1
9wKfzktGjPWlWOPix7hrxI6VrWKECSrSHm1+3KIULz6mQ92LM/n0mdcMJD5BEt66
cmEVDhnirDO9epE7jq/jeW1+oLh/WcTyfpstcP1he2eUJQQTBWK8zd6RBQ5BXp7j
U1RIzSSkKNpsdb6jeyRcM2+QkW+B0nbqq+12NHf16JdgRphVFtdDyKzjpCeAEdR4
yw77w581TzFl++nKSVNBxPM4iWo6iIKVmzz6v1/u/l152OlUFylq6bD89vFz7xLt
L23QJ8JgPU306Bjyhxb5S3PhPv0M74r9AEn7k2zKZaFSmdXDlgrcxzlMuFSZZVTh
fnTtObDsgh0O1BvE1T6iaou85R/DhTeWBA7fL2N7lCZVP+mPh2lO9sG1N5Q4nqkt
vTyCKaWtcsNDloMqbrh9V0YTqKLM7s8EFiKcgqGevLciezUEaEmNCnLp+Zm+UMhB
57UKm6Ss3MA05RzGkcKzrOo6h1zyysN57XGXRojTmFsaGk/o4FMAytBa2K8hYIqZ
EiBv8kzstnWgcAAnxcok94oM0RnQBofWoGSp2Tc9olT7sRXtmgW8ROVb9ASgf9WU
Q1Bjv9rkfmxgIXioK0Vq59TZImxdcAIY+DGVNzUZ/IZabmd1wxtclH4hJWtEY9Dd
qFVwHLryjJW1BsMXqttn4QcPPTz4uXtrTww4YVu6hrmKJSO95M4yPI4PmbL1gRQl
mUt0gQqWhtWMIalM6XB43k7r1xGiriFL1Ap5htHGPuUaMjepve7EHPb9j0zyiw4a
CgyOGh4keh+6m4KtyOtysRT6kQJ8qyEWCP7XWOcEHT8hGX1g6Q9KSF/sHRCVrRtl
st11b9y2h1bQ/6x9GzjF39KBpasPxluL3yrFd6yeB2IHBdcUoppm86AdICXWu34z
KovhyJe0bVo2AJui6+XrtVeKI8YzNEpDYjm+B0EHbb2TJphoF7+eXobq6UrhcMPV
18hScIVkE7uLfTs/1N23QniaeNVMHbwz2u93Na+uuNM+qEmwdPLLLaFD9ZejOwGS
SXdYvCVujlZ6xioDLlpggYK8axZrIvArN4xJX/Ry/63a6vX2OHHA9eB4wJU+oO6H
CTVZyrjD2ZaxDJyvI/ZGV2TBAXlYtoplYY+vX6JrUkHnjAB5REoQdQ0Y7oMRf+FD
GfzBOEWKbbMVUiQc6thUPIj7jr1zigCNsVkcDIWgTs3bmL0W5/Za8Aa+Fkyxcc5U
fyN+mq1YmmNpZVIhBkiMAUp62AB/qhD15+emmY+6mbRWGQystqtBA/qy2LyHUXVC
1lszTGgCVfJi0x96/QsPwtMYNnixPQ0UQEN6nJdWi0hOCSXwjPam3MU0YWeC7vDM
z5BiPOpuR5DwX1Dx5fIg152jTx/99WM/VQ3F9HnaDM8B8fvCXj2QWxAk4wHyCwWp
O7CkG5Ii/RTb7SOg5Jnr3trXWauneW9OV6CdFR0Gxp9nrUqjf4Tn7B3515l+p4Rq
ywFExN4B+kzvlKycQEduw5wbTXoNSFUwk/fmxorKqYagVdB/5ZJfzxh7gKkLUojN
1LXFfYVfmWALYcpOpv3RqN7rv9VwIxhTm0oR7kQUuZIYPO6SWh1okBA+iasO5Zka
hxyZFfSyGBkgkKr+hocBGEkchK2LukJFAExG2stH5cEedKNlPnL6/oriPIMgx58g
Da9LPEPSsh1WR6lDNXW6aevPIQqpjwgjf2bkE/a6fYFybWuD3WYWOnsH0n5fdcex
M4qypGLHk24jpt/TjIATG3Sja7uQFVrlZC6gRG3F1RcLcSpz2OZ1MOQLT/p2r2ii
ounUe/nbMqvQnbNFIvBf3mP5FZcfy0/GlJSYIbFSEjNrHI4jQ0d56fVEjCVBuDzg
icNIzoNi0+iUH8a2I5Bshl5Drm2VvepeF9l/gnpKgpsaDUVo7bFdhL+b2Lqa2ct+
RFCE8WE2MgBOgoLiRK3Nm5+g0i+YBMwmclWAoegIG98mzFl7qEQWlQxGoDRX6BSr
BCOQyFkbAp+N7rqzjzwCZRqe9jLuD3LA/Jp4oClI7wA23L5j4xyPSMQ5tK6Zpm9Q
1LVG4X2fUBBWihHe40ZHK6MpwLwZul+LWNryaaJggqxR9KF+45PuvKItj2807qea
3TULulzwJfSRXqu0Jp/CzqeSe2ADWMJWSHoBexuDM1JgaatbnqaNss+qSQysj5cA
bVvJqFig5jyPtUU9gVVFFoQi7xq99MTNybgXYHojYniruwhedAnHVrVtPSlut0fO
5TIAg9hK0O24zd3mXBa414Rcv3K8niIjM6EwoM4OXzEFtk7nBD0Lv+busWL62Jj0
eY5yAIg+pETvv7G3eMqABlE9wWlX0s68VzLTzKu0cZSv8xitdI4hiNaZELAUcQlH
vN8VJo8VfyahmYFfSFdiYnT5tQmzgC/ipcI3Aqk/NEhqsMtALTY15deaYt+R2YYR
BXwQkHurd2xKUGsc4XTMwxtvO8RtWLD06syJjMKkGXexQODrXtS+/5vyTXyh7omE
L+uIXkTIeROnK5hhU7V6+/LcYv1hQE5PGFJQ9ZkKtr+l0yr2dkv0oljNn0cOArHY
Np5GbYl8Cr4O0FDkDz4s5+QSbehRgzFt2Rmpo7FdKX+QP39L8ilWWLhA8OuWZx8G
f3cHJqdaBtef6zIgH+6HekSXcfKhwb9KHdS+TCvAhPqMrfK4VEYMtnjlaGTTCNa+
Vme90WOpKDyuTYL+BH2Z6cTtse1yQloLZ0x4pxdktxzZtm5Z9M4uuCecKDlDRgWs
B3AFb7d+D4yeRpjqv4qFIEidBEdg5K2pkdZOJjw5RxxQ68BBN47eZtl0Wa+kcgQL
WdYPCdMIbQlLOsGH964xj0+VVPp1P43QRNrXyPZ3RSaDLLxBCm4lTFVriWXVr7ff
5pdX/Sv5zpQvUBa4pKSx9eNjarcfzxR/KpKN+cOuDN89CyOku6zrWThskEy1RL1t
Eg/iX+fPd3RbrECDpaxhC/qDocJWIhRbfIswReb+neRUggmIDsLepSZstBJ9A7HJ
xoztuyMA/xS78Wol0subBeK467B3PTZShmnrcm5ZnjJIOcgXcmNB+WZwfJLOcILz
VDUKD57+IgweDjyVzlQaHP6MeNGLZJgxmzIEkdfwddY/gtSBGIft9LZSGxx5b8vD
8Skm375fJW0bipjzOe8WxHAy07rsiMThu1U9tji7qKnbuLKtVyxpMdIVhoUtItTs
9YVvDa/8ttXfNra++TC7i5ovaqQcQqpoPYWXoa12ymD3n+vn1I8JFtHkCAWBHBNi
/zztD772OkAOUaMI1DuZtTso8mEzxvp75RVONXHpk6oTmFLXbDZUHYrTnQRpYrRA
w89yTI4x9hDYseoboF8C5xfpc6ZWhfCUa4GVnT4Nq+sLSUUHV6Pg7EJo/LMuhBc1
NRe4RRGfpg0IgZEt6XLbvHHtJkE4tUAZcGIe34DgTlokMEApOLXawSnfhycr80WI
koHotH6IepDnZbu/xLa6slD+Jn6gxO69bzDnXbw/vE0kNh8PDAIuck3e0wgnSz60
eIVmgRM2cfSvmR/BnUeWsvHS5gVNAVLHULyPfDS0p4IK8klTgh2nyMxnOzs5F6pF
LpJz43mWKXMkEAEfJAvPsCCB9iAN4T1B5Xuz8SPkf5bK4Y+o4IlM7/04rSbdrhGa
qkWJ8O6BOtvF+VfnwrTEk4FgUc4HYTOgY5DG9/6YYNbndDKwiFVdhn38ZdowT8HB
u86oooBV26Ft1jAnfHgsYfugLrcAPyeVLLD5/cLE9DnEcIKnK/cz9Jo9Y7MQ89tF
oC4d98a+4JFRpr0kGArKv7NLoM1pi2WuiZmt7Z4RGE1PRcX4iILlWf3hphZ6vEAV
0LoAIgRL+Kw3ryshwKsG9MkKCMdfiy1kkityVxs3W2nMvaL2/hRIKzWNoLGcLtwk
C49WbO+udoYhJp07aHBMPn4VOuW7AC4QbJ5VrrrqP3eqw3/sZFqIv/BfyAfkyxnD
8eK7fEn0zql7v0atcr8GHyjPQ1f+d6VaWLhQ+28SPLLQVsaBmRtfOqX0u3b2+ecV
7fC1xukpVvaPmnwH76gqPLWaQlseEs79rPS7b6JRqU1a5nGIpIux9N2d3cBVO1oO
HtLSIEYePNY4FwJqxsp6EDkbSHOttFXHlLScot8VcfstMs8blKQR+HUftuhFydhI
wtskNiIGGXrbg6UCwTJbWrmJYy13WYlOo937Y1y5oIIzEAmZEZvaVWYk4l6Dc8WC
2xFJcTDffqQIRJscjlKknAFrpECw+6nA7fr+xEYPlUH7KnfVXBEpWRyBeo+omepw
f6u93vM+IeawRg3FvLhijAfTSiNpiPWvpR4J1dTRglHpCm0iOrDvQyfnS9bJXdDA
pWw/RbwtGZrEsdfulOCLP1azwKbgxx4VdM+ieelUaFFbXTyf670f/VR35ppMiajW
fqFe5e8mv6KbM5CJBLUb4MY547fehUQ2PDDkp+blLI8Q85HQNJB1/NUEtXBZ0W96
CHEzgpmSzsNCb8imKVmNVYh8nEPtHoKp5XUn1ZgCpiolMKOfBr36KTc2LKtIqoRG
x9L68V6hydKmmf1CQRCn88KRecnwCpjeQ2LzGqXp02TktzkJpAOuR/8DkVC5Jtfc
IpOT1O5YidKQ5G/rzrz21EpAuU2e2C/zSbcKTPchMrPe3CQzRijtMAmo6OX+J7Ez
Ju3/vml+ZMR69PMpKNNQMOYTO38LUdrtwJf816kVNOaDTqFFk1tMH570PGCvlJph
lUDg8tYmPd+ga2hR9qZBHIPE3BV2QZ8wuSXj2YFYWt3zMLW9AH2IltkHep7YurBh
aq7lzUzdgEw+RpW3HOVC+teoFsEKrbiWdyBPAs8G+f8/ZqEezIodXfOJyRv9DaJ2
2JoGKgJ9HQMMAMl3Bp9ZBzxSKxZZ3hx7IxuOvNVKVlxG0i2H/TSm/4an4bPxegka
JSLRtQNJ3fy23xn5qFevRo/QCqW5vdBpddxtJ5usy9ouABQB0w30/qdOWS0EU865
jU57fgQjZ05PwVe837cj4FadmvPtAuJ9mUftRo8qH8reHGnXmjHnVPOgf4DIF85/
QmyZKfCjHJUKz2VjFovlA3uRTjIjsCr4Sm3tzeZNILd0TWJWS3nK7bFFfYT7V95I
/6zGBZBTZECewYP5f1Xpl7PeO1s/s2k2WcUXVdbVRdgDcAsmg8Nr8HsUUu1fW/KH
PxH/d5MnKIVY0xajuPkN4rrWbIvy1sTelRJtOQpXlGa52bb8mvSuU3DrV2z//duS
P9rRAUUtvWj04YalF9m9JYhrfQIVL7cchTOQayNcRs/C7jEVvWBtv0bxn2jPOjF1
W+at8Ygw6D6ieVV6sueRtnSM1QZF2eDiYBuKLrKduea9aJUHUUoFbxO6J9/KK7cu
WuPCn4i/nd0V7xRyZXC+ywxsC0/LYVFSekNNSFYk1HCNPtmQ5oKQ8E7YxQMmgZJQ
zjOXHU955s22rmHp9Pl2nawqaNBnGZ0z7YFeOv8A9MQ1WDy/OiRWJ23IULyJIFGX
q4Emgu3PpoZGgCLauPwq+3SWYE1O+w/9GFJypCt1yQAY1hFxce/dsJAzqn3s//EN
uXEhMvCNz1lggi7DdYR4/+wdJtGIbeiW0rNC8YmRMxZy53Ny/M84l7bm5rJUSEuR
JrKjoGNb5OyIBpyeEE8S563L7fgceX92hy9peqTNt0mKbTJ/OJiOlSc1fQ9/jZT9
9/M/KNOD5WEAN9HXcc9A2zJp184pTE8J0gK8pJQEqTWhIAy6TMWFDCf7vf9T+Ok9
X9DFyPy+mkV7iT9qNQN1FvVmWjKpcsbmBoHRc++13cNvSsB2hpwLXqY7OcYlGiUA
QaPXIuxxXJy6hle2EV/DQf8ulnwIMG+b9JMJUi1H6xSxrulSQHaDPP73hAKOHjUI
RTACP6AZEwP593tilBvTCe84Li25SFZ+hH9VY6g1U6LTclD8qKYoYuyYPt7tVKQC
ZAVGh6wXojxHc+2HKrIxvB+Jl5U9JGAtdHgAVkkRggkjcQfn8UbT23SwhqhxEYXw
L/Btkc/PbvmibYFFmBax9neEneT3h11ok6NmznBcnz/TRdrcr5eACmNljk7pHKOT
m811jCHGIkZn1bZiJ1EVriepSNg+VIg9WfTNO9h9LsyGPBgssANZ++Pqvf19wa9j
kOHmW27O6nNPAkt01C1sHocBZlfWq1QdHs86b3yfqCG1uQr0tszNFccSg6geIAf6
WoGox/0iX55wx5GX8e51RkGHE3gHvFaDA/Yt7N/X9PTb+g8gtYAfXwpvO69t4mys
sYdfmidzTtIREr0segntmptwI9SPNTLCO3AAw4xanpvxmiaQYruIs34qWh3Pg2Mm
OsDMdHoCkosos8xBSeSJqAut0La1cVvXmw91osR6CwXiqQy2MdA5fK9Rfmj9B28b
YZC5EZg/YWjRvmf0oaHbGMt+7HTJcUFPRtH8nvrmJ00ez9LvXW+Emq5yAAwZV/Dj
MAD+gxvsxnysBBKKvtQsFFlnlQCI+xZKmR1DWvJBdmsnFj7IIl+dCzWVyUkAt4fi
WmzN0DLo3dUxkjgCDvGFLNVaXGnJoogUAEWClMS5PfW0XjiLViEx+tZohLXVZAMg
+UWEzaYsAgUnAx8q1ylu67Q2VB4pRz0O2ScqWs8lJ2qOE0EULzW4rjmXw5BekH0d
lPa+ngye2ToychMcfArH2YTxC8Ek/uKaAOLoqLMbERmOrC049QOIYgcMQYW4EfK9
5GsYqDrHa9/Dg7iQIQ8HNFXNZGiy0gBhPJVI7EiGwTAGX0UUL1nm4lAmDfZ6X/jw
5KpJLbkxvSu+dH7lanJT8uQzR/L6h5qvq7EuCdTaK5Fcp4Bv7xRmihO51Ke3OVme
0IHwRg1K40VF+YoYipKEj6Fbduxq7sWv9MW3Dh9Pe5nf6vlX6Vf3rhGb821N5G0I
DEf2LbCDPN9a/P0XtO4Nu+FItbtazCH2e/P6J2998A/eqjXmOuTFue/UReW2WMjz
cKmxV9/ofeS7Y69faFYSDNeeyBIjc0XI/4oGO/13QRQyGSh+F08NFKzF7Hi4eUMP
WRJZR61ZlyCt33wog5uqEMkPjJ8MEGSDxzl15BNtitZapwwD6YJ6tTXV5BgRfmYY
dGk9Fty7E0YDizPsGwJuTeEeiM4iPaYVTF8YswCowFo9WKIEU+PfNXNQzHNHt6my
1xHT3IujuoqiSfHVYkxXhYOlgawr0HS02dJ+rTRtBeZk3bnaP1mSbHaMy5lHd7FD
AZd9SnQnTgqWF2LMLhQBob+V0ep7tQfsx24lOipvhDyB14zT7mYkEWoIf7tH7AOZ
DOOcWWBPSB2ckWi+BicKN4OuqY0boZejzV3g4HbV1+l7X8+JAwAyKfhcmP7ppnr8
AA+3XcCK2o6Vwnh9quw0lpTvLAjjN5xOEukbRXOx5imufkQhrwi+DUgwogXE8p7L
gaGPZ2xQkqZac3cRilIIUMQ99J1SLxdQlJ/VawpSbdugpG05XtuhbAL3uz4flJTS
82A2YgGha1Qd7Sb1VODPDR6MbDWEth8re4dtXcwwIKUMeLWdIBcgpPs2czCBTXli
cyVASPiqcxS/3Z5I537VSx9aUPtNAM1c9k/CcDsAFNbGZMgBmlrhaTkcSGlg2003
pqfqi2SSAPlOwfUiUFwGkUHUUszw7xLP/BfJTtgRImT85axnPnQGXeSd+GhNxJqy
2zfdBB/iLN6OhtqbUfrtN8rO3Y225UxDnanRH/xxM4oXmebdvYX1Ram81KzTwFqJ
pTg5CHt/al5Ws6BllcaHHH2SpBRBnYZbtf79tkURFQpxXX+7p+eV6YQycO2Urfky
srHElrv18rbhirug+Vx2yPpA3rlBWPdYxfxzH6b8NHK6mqSe+rh9+BlJjeaoeW6Q
7btst7VBWJx3HtM2rtxqCgnIhMszb4vWvW7VJnZUQPnIRGsfsqIIFhASdFso0mLN
FOg3UlrV6bYfN5Ad+Dz48uRHbEkGECceG4OudZkYTsPPlx8WskeiosEHCvtiB31z
VpPxE+dJqT1QFPc0U6ZoRMBZKY+wcjw+Fw737M/wX+UE6OrQrURTIsYsOniUCRP7
Jin/T6Ba0BbDh7Vi0PayQGAFMXa0W66h1vYuBLv7VDfjX3nDSOYcZutguvoonMUr
VbB6CVUNAuNGSUimkH8loKITSkjnah00DRNTCws7K4DA9MfPNgPcX4ldXF8hmW7C
jqdRFo7rx8okZmhT3LFdfRiEAxxS81A2mZk4+Nb9Th1VeTfXMCUcHfiB17dUzs4s
fS4tCoxinklummjn3vPnb9CaE0hKTH3tvyD4kwv61qX7lEuml2CRR9aPdCSl6VCu
d0tYUZXnI3UL7FdWjvHOnuYy4oZSVW+9hpLcWNbfWNkXLbf/WeVtpTunAbyJFgD2
7h8ymGhNmoyNfXW1V7unw3/17bgHfjcnEhFpCqWXMu8SIwetYTWAYZTzUC/ufeqW
NOD1Dp0G+/1UeoKEv4p+9lTWhS+nZYDJh2jYYG6OVF1W2Zhcy0VZ9l4MVknE8WJl
LfaNB0L4jkLGzyE+NvH8j6r1BvPtp8cS977plJZCUv/YKw0wPG4Xc+R6IMUpgOSf
SMP5BmVmrrOHdhwf0qUpIYoDDA66QYR5kMxwHlK89wjvwb2fa0vlbKn0pm0GH270
DpPuoSXBuWTm/NZSgb9QoOUd0DYuobtJE4jhdek8sTki14B9nVDM2zdLH/xsMZ+J
p6zkLNsrShTRpllQrgLZmUDqUKN3gaLJlRV1YwdanK0Rah0dQaxoy3s1t4Lqu4q5
FvpjuTB1Q0lXb8pbjzZXOD1tHdkSl0Wp7WjkV+L9tYslGwivbCMriwcrv9EQVoIW
tANEyvzOvS1k79+b+M/7Oh2LnlZYPi0q2UNPHuCPNuADH3zbb/MLkoYk66GcGC8a
z0hXeKD2QdP1lrlZwB2biJ6uQkLfjb0fLzd4ePrwnxa6Y9tdNgKsUblWEIDqeF/c
7kJXkqnlWnGDUUHB6Blelbt1NMdo/CTwCxozu+2fYkjGQgXCY1YZuwm0wthl9Txd
diCVnh31z5+XZTGzyGIa/m6sJfT7jgJRhdUkPXS86WtzmIADq3KSrPOHYhsT16h5
mA1aWj8vj9VULoEUBYOl3EoJUucZSqzOcgTvYz3DOFKgqj4s+l20IBsp1So8syJb
peC4BDDEAgVQCxcWbaTpCAvuR7yEX3+lzvDWmRzIfWRaiTRVzGk9i4iKA7DyXivC
lGbS2QfROAT+6LqId1EAFpElACaaCnDYS5jT3dG3VxPnoNEVrfO/IPmBubS/N6DJ
KfdCc9XT/KpCRhY7BpbJEZynJvAzwp33CbnxqrUCrtoiYbmaFWVr6kee4mxkfbij
OkCHjgfeoGOw+WzkXnoIjMMFRe6EQymCAMg/r7D3jNK+mJC38WQH1ZOkpqp6M3QW
Lpmp1K+q3faVdPf0eAzpkivfgLsnrUI1nNZwEmyFGHDUzxih8pqSzV6AM8/FSrfv
9vcAlMBrjXZqTfk47vg41mieUusWgemUyF8ZGn0y3+Qmy9DKD6ntNu+IanRGjAP9
KWp+q1KfzYYiDgSfEnVlrxqp88y1OJBVUM7DfVPZTILAQBmlw1uEyaRdZlzYGbwK
v2IfMAt/HeXuGyRiia4TU9/m2oEbOMK3hnoR2ABHaHKMBKpxm3FUqyGSbeTvJhMn
G/2frXymqMb1dyduUBkcw+vA8Ui+yPwsQHay3Ql8E84AQHTtOPKjzkU0hZmOyRT3
RqX3FOFsxIaP+tiR7sEfybJrWlCUErSlYTocGRJoj687Jh3yBi4DjkM6Vn+DZc3q
P9AzMrNAxKjN+VgwUTTBPbgL0DiEVdxKy5mb7l5P2GahJ1cBdwF/Dqi9ibDRV8yP
FrzhdT5quJmX9XziyfmeJ13z0QR5Cz7uSRigWf3zkfhlKEfsyrsEZ69mF0NsTbOp
Tf0nqCnEqCgCkTK7gHHKOoKp0vLfKaFv//vep1vZld2nf427QUUtEbQvrdWnfaEc
y9Ljvx1qOzzLkl/S30z6zweJBP03xBbLVOfsoS/9YtzQXNyUoE33gR2hfhXdYPl+
Z9SbfzK5UCGU75D4DnOWblJSih3PJ1XfFDG+lYLOxj7MvFvocq4fGeDR7ZlONxSv
yrstVvXrT6b9C0uIQlCMm/F6lC5VC9DvCSHt0a/djOi6LgbOQl5tn0uZY1esJiq+
MgcA0otiCotIWuWe+hGzBLG6+VpjvGqeE0GF0WTibqgd7oYZlqy3HuLNftIGdSRY
xG0IwKRjrNg+GVzQH7bv5kg7iroP5OWyb08UvScnAO44lyEaL/9MwfkwRktYqwrz
+UTQAwSwFmeYmO8V5RfbxIWkgvX0N2DYMC8B1WdhWxssYBw7swtzRLLivbdo5nIt
Ud/xyuDZHbwVn6PFEZO2OVGBiWRniV9E2ENCuBFGjVkKgNqU7U0PlHqKFlR0025a
Y2B+QpArp6hVLV9P8m89nbZ1Hag5P4O9Pdb1SsYcfhceXwRUF5sNMdtV0TfHoZ14
vubX1QF3foIx9YrA4qog/5D+s81RACzgpmWnbD5h1+aBDZM6/NtslR0L1h4MWqD+
aZXh0+5SRLIrjPQZ+VI7HEfp49VXgdYQ10zKjoaxodCpt0Y96T+uIt62554+4Bu/
mMHY1lUE7ksLN7BPfImS/LiSIIVKV1liEgbi/CC5MNoiApCxv248/nn7vd1alji2
l+WCmqUtdQ9NiQCs4FpGr8u6Bot9ed1cL9HJOCiydOwm3vali0XjGMjKJjmdz9A2
qOitwq3fojLdP1dR6RUdrZGVSsVgU1YBU+PflIVDMiucmvSibteDHmR+4iEOMZ2U
EEVofKG1T9OecRNqL/UNrthrNTZydHVHXmQ3+g/APpuWfDSTKErCmykXuIoiWki3
ldQPuGtXhvyQZB69A15zQ2FYG8uuQqM/oPEauUAQ9HpgfhaJmpNoNRfelOzLk6Qz
cUnrb5A9GZ7fxoxu46q/MaS3uzk6SRTurTXW5XFzIFj5c/1n0laTrfvoiTVfareX
x/YO1p24bH2Fh5RXUjnHy6+LUsydPT7Lwg2zNqrd7JwaE40FUzGAiIT2i4zknTWg
K1Ji/LziuUxoK9x9PKkNSvrgMCuJadwZkV04i9SfpX51WnwoXlIN43qJwdPkUGsh
w8QBNfg9a3WAsc8MQ6sQZ3Xw9TSBmme2vGJJmc2qFIdFdUIRuTBCuDA5Js1wu0EK
KOTW4E+yhq3dQTN8quc/YSeKZSBJSBexaXPXP1RPDkisyiAfQrTG+g3kHoN6n5bG
DlozTTkYUilX8UpdTfodVXG4ZFJS2vwsWX4n+Sda+UsWvwWC8p79DRQysQ+aqNr4
PPvNRE6aH5tebnYnnma46zMoOFph2eyb+NCU/UPJOfLN4AJBHp3MpWqH6ae2YaUS
kCg2NAMiH/IEnUF6BM7ne1/IFhXNQXuoilhNrMek9JZddpqBTa/s78M3QwV9APqb
Vs2ZrZf/MmWzZwooqt/oB8zvFJM3tvL7Alqr4jgwKELAZ9ckkK1NniHpbf9ry+3+
3P0sX0JOv3q29QqOjp3e+CxnbUBBxERG49zUHz8fc92F6fjDEt1jUERtlqshieTZ
WhQ6Mv88VOXzgsSzY5aNEezBqIGBR1Rg9SJPLEJhe8s7wV/cYVheBfMtCWn5Y0hv
f1HjFBEwdXK5DvHjKljxBk2e9kyxphRmeF4afbVVBGkQhfDdMhTSKzcAJY0VWkjB
XlVv+pIxXNThvZNhdR9vRnsOB7HuXInWmiaTZDIU1NfHVFFzD2at6CToCRc5O+Fe
D7dHjzxTG6PtR1+ctHyGLWs0bc7eNUur6dbFHI5NgsP3eEqBq4z8280ouKKf4R0P
OBZ7qf4Q67RpzFXnjgVnxu57SVphoaC+LP8MPmsJCm9a4wQdUbP49y7zb2FZNJ9F
AC1qhckQfdWVxKvH7y4eywZOqWU6PnRPh6bgwq+RSYGMDjBYlTJcKq1jv7vJF/uB
IXM4J6SQ9Spcb/WckiSj0IGuvLv8SOBr8dux6Fhdwqcy7JeQ5qajUwxsTovB5v0I
OXgqIV2Fmt8n8sgEJYoCvEWkRpNEF/Xg2iZF2LY3+QQVuE9r+dsEFpMK0P53DltP
ExCg34PffMYu88ZIhx8hPs7PY5vTxib7FbnIdbOWUj1weXpKUqIU8BUeQScGe1if
LYgJ76TLIy6J1jMT6X1qnK/CeMOOoHBszQLlvaHDhlK7cj0K1Ayq6ZpIaYqTqEQj
ZSRPX5QN2tYkuz28PbeKdzkZ8T/AWDRPH3KZqbtBV5ZEYUgPCzJkYFgi2unHXMux
C/CZNfI5A2BnIvDYJA1R/yqouJy3uA4kUywh1uUAN6BLObZXhVbASxQG+IEvgdUB
09uTpUrD5VXp+r6KP22WO9b/LlLo2i2ySFtrH2GEye0+j8NjLU8KrHcKCvMWy9ww
hJwLblCAj5bhqmATTOuC/xA0+/JUEQcWizm5V0Nn4osThNFVGs3SBlH7lcIOIDuR
gs0GJKQ6ZkrAgWvYp7Zgfum5NBYvd+4ZFtk8OIZmXBAVTiadZAo30UEoDPzG3mxL
nky8DXOMilOWg8WtfHhyKtvXxnos9VSRtTRs5Bck44/Yb+QC6HTS0pm6qX2M56aF
jvaqLUzgObEMKmtQAi/eO+QPvJS3atSYABkQjM6p9IzlR29faiaar2UOFd17znFY
ycX99oWY5oaKu1zjTLc7MPqNI2x/4+601+DKkSIMF5ephTWwjd3qZBl+FGx1ppDT
DlpxwQsqEvOniUtn1SS0eLSePvevhilNbCEwH+f4i1kiD3OE1V5ex6dhJp93h+Qg
2xmcMcbPJeSqHbh1BYDJCvKuehdJKHdTH/FFuolA2h+VGFJJKAG9ZZ+bHmMI1Bhk
mzyZfQ5nNnAT9S4BPpik666e4Hn0J+/o0UID2PyZDEc0v9UKmH4gWOxJ0DPO17k2
XmQ0WQPKqeG39LQM7RdU7Lyf8MO4KfN8mYGgCw/N2pEPNkuQ/ZhfikrJC7aModl3
bmwnkAFFpVR+qoI2jYpwAY3NCg7OG8Pk7APM3+c9kBoIliOVziEf+rEoOhYAZ0gB
jg4/v4/qZViOciy9zMoOsd2eC7fckffJmazDDx0LiN/WoonjUFTsLq0YwK4PZVBg
RriMWBakw7L6ZbYjv3cnCRczM2hW1H7I7oIXo6sA5SuU5r+vUZEXCQNhE4OxTt0G
pevnswZkv+ipAlYDi6Yyl2aaw+iOsKjdKqg99MnAzk++kJKe7/AjGL0HVTQYz5Fj
113PSjTrZh7w8g2rLXvgDLE7bDXul65YlG6PrzJy8zzbmxTDgGdlIQAVbSqGBJsT
mzFgYhpWxY+8722KA8uIldEw1fLbBRZRHg7hylncqWt6/q1GLd7Fs2KyViBdLhTf
o2aiN/3KXiGh6BAreut9glijm2vrv1txm+iyrs0AfFeH4kBe/vFMDnkAFVsA/Zx2
ixbx7zO4VFgaJS7w8Uz5JPkZeUv81FqnCgKklLrFc/qkXQm+1LTEHTVMsJwP+CEd
XTGy7v52s+wQi49gX8dPwy+2gH67+kuUdHOuINmayuW4gtr/ZqO17LESH1tYXR/H
xr0hnSh6f3HgXPDV7bsUSS0MNuV9QAuj2CMkvGXDoByYujUsdnBHhVJruBfGpJRz
+h9ZMKL+cViC+BQSgf3H9a67Rd5Dk2fzM0wtw71CeqO51wsfnJ2lflXs8AdA3NSi
k726DOIB/llE0g1INc6ASeFBbCrwdK8QCIDHkdJlIXlxfyEeU7YUfqptmcCtxOqk
bkL1mEPuBjcabpQxzMN4wpKZ/1+dJh2tFbOZDHuZzn7f7/xvch1s7czhR/KSJUcs
od2D9scYduHA7YNey1X5VJRHXowKn0LlWwnk21C77OST0ZorH0DQh6UEiiEUMmU0
HwWklAOmvJvaodrwt6oA+bL0VFHvdpDekVXXqsq7y3Av94AdN4y1pBD/CpO7FniL
9aJ5pVl7TZ1p1Yuih4O9cPbhhCxov1cbtE+MV22VX2iczsgA9M7vMRnVi5pYO+bw
hZBQlflI3DiHj6iiMPMxYjKc3Al00y+HJ7WGRI2GzV9A3D7UQLwazHGABnsLVyLC
tEbzj3JVyp7fdf9Mbe1da3aMVx/cTaOkQcOm/hp/R3joln8zAc4cKFmg+YafyY7B
KbXLLvuofoSvUJ+il11bg8V2YhzSG31LJXxm6rmNhLnejx7Om6gHu/lcB4PBA40j
4MZQR2RXnjP/8rN5RFRyRbeTpNozD/NiGYLHfaQITO95tHeKxdHLh6/v4ZBhGcZD
7e9ma8SVsJmnogpyjewyfXwDSUrOCJEgL6e6pCCCoin+6vXN9Dz3iGE8E6fzWHF0
9xMACU0ByjfssC4/rN5hs92aqz2VS3TyWimXcvlYXWxCWqnN9PW8QXj54mpWvGTU
fwrY4kok5ZPSADsMgIRR4gvWxXrKaht2IEgllbOQCkRHJwVBbXUnZyBCR9YtDRUJ
qbIywtjcMqPIeIAFkpdPD6a3T2aagfFoUclMgdTEIV3HZ3iSZtxbsjsKzNsvbQfP
xPHAHi1hRSFtBGNrgX+UAk54d5RRCUTa1Nj9koA5wHYAO/opOiKlgsno+OYnkN7G
gbxaxpphT+tYwVSYRAvmLdEyvBrhXe+J3AsG7pvVjxejrgiCDo5VEO7p6ejuxeSL
3iJZoeINLYjInh+bA16QMwmjRPFW0JnOCSyIQxXdUea7dcZ0f/Lz4so8NGmKQSM8
vhBBWGI94DZAPDGkNyeirk+T6FZeOZSejD2C/EFmd7IlaipC+Zwr+b43IcPw16VU
sCZuzmhJ2/C4E318sTVDg1pCOPGQZ9APQ3CswzEGrRqmT6Q2kLhUw3/qI2P0cK0U
HsqQOoZ2/TcmZsuw4lH+cxA3yPlaOV0BhU77lX18dfKxa4ZfEgY0AyMbRQ4s9w60
KJb+CIKjIKZ7B8vxiEzf/DQAFXn7ztVaK7cgFY/A28dG48LJA/cT/ekIWwjgyjFa
FcpkS2tK/fWZICPLjxNgwCOf/JgVE29jREa0pfVQba5TjtjC+U3fC8fl34Pqlh71
FSRFRWBtSMqictYhmXCoEpkoLXIyT5KlGWneJA+xisx6k4Y2oajP3p6Bx0myd3ZC
L76d+xEvoWrooFLsMdOnkDELHR5D+2yhW6nwP2p9sD89FfaDFZd4jjYuYFJhWoQZ
vnlfj/xZN9DK512W3syHlIDaYGHpArzqSOmrfuSYmYmbI5RPCMmr7LIwMj4ShxOq
yvh0ymfohVHUdXkg1pOgcULpoe4JM+lXzwjox1vVK34tx/+8PxxKfbMk3h2a6KZ2
pMFrQ4PH6gOeXz4BHuU85HOnjJ4vtnX7fT3/dB/R+V5i0faFMHNtdopDf+jw0sIY
Tl/T+k0YoSe74KNPWRNI51PW4w5XB2Ff1/bGPcIlvXOr4FNAeyM8hQAAs81S0rtm
wvGWixQcmsAm69PmirW/7fxqhcHAKWqHFU9rO6H89YdGfUAMXowANDUSnF321bhC
le/1wz51UK6BRDcWuBCwqCQt2SC7BfZv8SxcOHuE1vIxfqJFYCiFAFiz68iTZ5La
VT4Y7uPMrtp0hPJb6iMEVQh7myNp5LJn7K62rgth+Wymi3ubNKMwxOEtkvoYLi6w
/m1lm+9msJ6yHQEB1Io1slVBHa1afuvqHISXi31nb4TufNshM9Z4byuPS4m0Pebj
n0aPxq5V2XiunT5QLK/H7PfbNJdQv463hqhu5bGoGySQwTnwrtOwbT7HheYUKG6A
y+HPMoQ0pYARS+OkWrw8x5TLrZ1IE0dIuWjd9QctYDIhclDl7WQSeS27InX/M+XO
ZK5XJcjxFoz8rV2YqbPONZ1Ztt5j0tv8qtqZvCc96uhpiyxtTBOIRroFj3I9sCw9
0ehMUWrASaVMbGekGHTzIj4dVzFTfUyN1ripbZih1E4V4k/0w+jNWUIXjDnH08Bq
PuVrQkB2MXaMV7LLqfG8COxUYYOseNNhPnXU694gxtAyBqmcO0QXFjdmnBur9Jwd
LuYV07/4Ho5Xktd6Pvzm7Golzsfj2kVXH1AaCB8i4bu7ApTEVeMshjD1TnZb4E5s
dN0K828dQLgJFmiva40sJOE6i+3mTx9vr+F26pOm8xHLpuMww63Gj/lH9cupWmUr
daga4tiM8WzxfCjNNKgobmJUOwsbSi+VS9yaKv84TRy8+nJATTXzmqkz3BecsnRR
1j47gz2JINjA0HRGKNeVq/MLba4A52yT5dVZa283wtSUmiWvkG1EmqumlMsGe6hg
l2e7X/rUQZmfMK6sIwdObDN/gdg7x3LMVWi3Zxyb344qfv2iZgEYF+JHhOQJh6Lp
T/P/TmGAluhKKf4eOhsBK1bUY8IfUvoO9FcFj4G6n8k22EQztL71aXYy+vj4agQy
NFmXrZAD2gVNrvA5DiDcTSlt6elPPA3JrqKoY22SABWeRNrUviXSNGoV9nYSghsc
6B2n+pgt3euG6O30XeiPsGDtuczdpkbvIZxy4C3L5qILIW3oI20vmSjXO2M0EJO1
yqymT2+HEJGPkUtDI0iQXGqJRftqC6eYeFEU1NwIjL/yoijyeWvLVBpFMSPLIsvR
sEm+K8QzCdOxQozximeNq22KbP6NoS/75i3O9j/IOgMYm4DrkQSoOIibtNX/vI0W
Ahv5kDw5H2v1y4GxqwQjAbrsil7+jGumhmdd4aIHQgMpMSiBjeHmglOxJiji6/M4
lpZ0nwKEtdhE6Oj81qTSci2/IlZ0Hm7yJjQo8NreuR1/yn97/FoB6g5VVh6tFaDa
cCcykM/bPOo5xOmK2Oz23j/iTkWfXrPUAePU0nEw1wOeZ/o1gExPxYn6EH7fR+Mp
ahAJ2AZLSzXsUCP+PbySpxIirIFOqIQVGU/s4eb5gSkyHtHlfzL3U9KbYl0FMe0R
8A8sU3PAyjwRFWvVX8QhIKTCRhAqNCc4QbPGA+of6T4ExkwkgVqOKQ9vA1Hr/qmO
FwLu5lA5Yv2MyILgLPQiHz9jmApl2csTwhDRWmNnoq+OmmHDJd235uIZEiBDyOJX
pKaj52MQGkc68ZAqGNeLhZCafc2fnKTEkgFeC058hs10blxlDbv+xF2n4/fP0Cul
K7Lwbuihtts79qj8GjV6y91nY/wC2o4n0LUgnuFKcQYU2meXn+wDU7wqcWUnGCGX
0PFRCCXPPq5MgNfPdExkLk6NoYemqIng1Ftse2Nt9Mr0S4jAIrVPO+aNf6ADBbyE
g8UxNFjKP5cwDc/IKvlPLIazFAMu1u6sk8GY61FkX2Te16/XzWfmgDNQaZN3Gtsd
ohLYqkFlKcWZC7UsyiuL1b+hGzOadxT2KGqQeJhCmLUWEzk+XOhzZNaZezRPDNlH
CBvKpvE+iLG7YsBIafjjjR7VFPglzkvI9lAPJAPu7zIwhUUfdhYupaxzlQde+8YQ
jLbOflivBGjrC7cpBEccMa0zNXLX6U1drYDTEUFURt4XU0+SDD2QYf/+4pX6BGMP
av6a15AvaE5+bDz1W7VJWqCskQZihS4TSBJ7aFcgEtkkl26axWPYJ1A5yRb1uhY1
VPaX6WapaC3/h+V2cWzjJfl4Wlc2yiuOhdHfPf4TtZX3crcgydScUXwSZFHJOVez
4U8/4WWoPtAQXtuYZfpoUj9runALHCOrceWFIJqdJkjY50mCg+apG5FvBpVCsDgE
KUBhZD0j3C0SD0d866VEPyWXkhIlNDEz0NtJ9wKHYDHYApuqVE4lVHhququ8eySi
MGwWa7/xmvnLK38+DZFf9rDttLLwmCagaYPfklhNHbn0qLbXCcYjKe85moCsYKMJ
7NcpDXrbydyOg2HtX4ungK7lPxgsyWNXlfdVaHoQE/JT9wB+nPLTeaVtBPr32qm0
vkZIoLBAMCyHbDI1X+B+d5UYGHjHgaDiDWQFu7B2/G4SHQSzlPJKTmMjrKBdsLmo
HkPhdXWUB04uDQSqNlYr5QvIgj1pMeS69GBsQiy0IYKzmy2VQcmzDzjDyvFyjxj0
CWqpXFn1/PpUK6YVsznTiNHAQQNtEkcWKyfJ5zOrWfvYheo+poeJ4s7G0SE4+HQ9
tDi8RGPdLuCDsaFCSD3JX/6qs/itWbEi1gL8Y9NVmKsQMBc3uIYI/NE2vgct+HdF
9RJGggpxJdg4kFr7XRnBDohfCFX+wB+QIjYtAm9uj8BJkSdVVPbqxVwlyZURJ2jb
jeEi10iC1pTa5CbByaGW7QRncL6kb+Kh1W1Bvb2HSEtFSV2d5x8GpFHNKyWtuqPL
dbhrecrYmGBZBlsrnesg+PguJjnz2TXwQyh1amMQVoKUZu73vDY7uemDEsE5g4BS
UBmAxhryx5fpO1ZPcZVzcvyAi9bvs2gdpPEK/bc+IHMW3x5sjDtJSNp7LiywE0VK
fB3rVyaKW4m6rlxhGwUtvorisq60Xx6JYRftZxC7tNg7Bks/WTA+PGUD7Gcy9omg
QuEVbQ9UcxbFUhIeDTMD1iQimYQwjAp0g07ttXFFtERGkQ8BtSStvlLlGDPVr0y3
qbeBbzm6D99+suGhFEyx5Be2BIdL6TLuHXQ9tNQ+ezuGbvNbgYL1ChXvFBRzjqjy
q0dhPmW4LFsiwnjIRFQLKbs/0BE0uQfmgBglz5jsefrHllAn1/igdgtclAcTlhwd
Ib8n3AYHJDLr7i/5avtpJM2PH9JHO7aX1PV8Q6RqMmkEhTIhYK9Gs6rK5ENypQyj
NZ4u+h76/Qv5UAjW8ykaP2di29RtBvULgzE4NyJAo1pt9ZB2lXfbH1munFGjvu5j
tprBwD2UNvIcHPfYbwGf1t5UOnmj7t56B1hkP+ugS/2OXlrfORFOlPuPkWB+I1W9
1QXJEw6KWYYBZfaxDR4TPB9y2eWrCbP0/SzpnGpWpZh5gU+sv0yVhNhom9YcJmeQ
BY1nE2XMdBpekJJTFOJz8rCaM3Oab8VZz0LGyNmuLk3u/lYaistNEKuyOooqjRSy
xdSHtFM612UVKlBW7tzxN/Hu0icEs93ZiRz/kqS5xcIkKeBSob32OKLkq3RVXRIp
FyUTy2CJKurcefcSCbmF37skGCeQr72qaTMs8HJJNxJ1/cOhupf1loPzQinxlf9F
AJolc0c9cpmoYrm/gkpzcjJjnlOwcGokOUNFfS/R4n/NJUOwkDPOM0n4EP7yziYw
yJ0X8oggO0rgR2QWte5Oo+Nh719T1u/G17SDSs7L83fpoNFxpQ8EoIb3zRM1rP56
hO4OEAsRowwRrQ7V0uE6zPqHcBLcrL3ozgbieAnsz1lE6jNlvtciCMJSLyxah7Pg
JTuHp2wqnJLSpSSweJ0GeBfWXHhFrJARSDV1SKr8uRGmZ/7wkbmwczHs+EA/WeMm
KlGdLQkCtcQXI4AIWc8wLu31sSLhUETCkSumkd67LmxJUSmcFN93F/MP4RE3p5+J
MqyPuEBWmM4h5gKe05aNcTnWaWljAaUSrRmbPUPUj6sd6KgvOmMm7HSIDUT87yA2
2aWDooyrmfUnUKm8I4reAB0KZjni4/SwUYScA8s3T730M8kie0QsHniBP9wZ2c5Z
5XWrtIWaOTWV7/DLGWxVr26/TvTNh7kIFTCzO+dejuGi4TQuRzNYphNxUIYxhyMu
L0rDJE9A2pWQql3jSmMr6iHw8/3aRhzJP2WBdTFgiPkrw3/myWd1Yo8DaG41Si2l
74Z588TAkuDqjn1Kim0KCLQ86MLlqkQV8lyvtXSIQeHKoMwDZuQJPcVIp5Gf7rz6
UX4CH1YoDRwQczB46B1uMWHAPvniYuASXIvpoHxqvbESifX//R+cs2RjvUfsUcQx
B79Vw9WwexGPUjsUgUT8mOXh3iytiYFkdfeou+G3FJ0UAaDvgvu9TCt81xJXSBGl
OMBWdY9z6zEfOuVaL0vsLKsXBPL7FuH19/eoKIjSHYQEoksZvKXGOtPdil60dOzb
/4RAtbyHVf04njvSkY3Ku5jhqFRQpkmiQXp8vXJWf35LWegoCto0rCYUZEO9h6Sh
7gglJ7L3ZjW6pxok73oIbjiz8Sh6UYXzYr9LoGyz/m1xR5M8bnXdvE6aWCAnHqNT
wTq1ayOUjpzrJCwX/KO8byG49l3VuRSThF2SIJPBzTk830bdfzFxcEF+Jos42PdG
7ww3+T/q/MtG80lvEhpzRbjwSLHJCC8KaxXrVGe1a5oEOwufJb/Zj9+HCQ1IIMXy
ZPFv2Bxvw73Dy/edXC9VHFJ1Jbx8/m+LsqgglvLP/X1J0UDt2FteRIv7zL8cfCcS
eFkEaDwlD/KiST+LGMpBGFvcgMkuEGnirYA9j5ECkGOBRZIpQpbZdRsTMgibgJx0
9/jqzjB4xf/SSP9zpqExzGFua5A7YPa9xBVbvUomjy/UW5tZLCfWhXSSN3wCP2BZ
XiGXP7r48VyH9tF9snJ1ieuypj7yTmOUYRhMX+bFLrualhcEI7PegPZ8NcDGpXiN
xy1iQAj5claPoKRZ/C/dpEFGWwtLePvphm6h3tTdPddTPMzY3DSxNvGBM9D9QxLc
8H1mmGXg1iznBixTppstSOsBTXD4OfmNeCkddPMLwLy7qxwsRCZWiiScgciNE3cT
uoH2GmawB8eqU1zn9lpJS0f29QiSPZi3CaVHLXMFJV+rJ2QXaluBGlv5tnpGmDaf
QH4Yg8k1MTJw8XSVixBXap7SoDMJY1RiRhOE3Io70f9yK1Mh1MEWL7QUhe9Gk0dE
UXw9QFwe8/v2gPinFQ74cVvQu7J60iujIOMLtnA0zS+itHRMYODr8cd4gl+xANnJ
nd6dccSQi8FqdIWldFS4FvZmUF5b+LkWzVbzGNbt2IQ2fscArSlKKE9ADDgtT25k
BvgVGJ8FbB7i4e5gVhQBPWhK3bnqEdPlPHA4Vj4bA897RJlACXFIqWSzvAu+H8nJ
By0+4bjRIIesreMY2dIwfZnUGlkJ4LJENr9GnChCPB0Ld4T54f0z1vcwG1ELFl4y
IKi2Hly0RZKhgvaf7ELbyCOJYRmzbhsEEs8jcnfcP1K7d5cpUizfA/vj1XAcHuZS
TF4uGRRNHqTvfPg6YyBkwpMkq0h0bjgjFYdEM0E5MUylfNjIPwoMEU8n41omQ+fQ
lv2hKXaNmMeOR8v3QQqLOoAx1lPxsyAvit3y6hdipDlRiudcnnA31fh2ObpT/go4
od6WNAUw35rtgKTJDkzLPDNCGy/4viOvq4JX34ZwZc2NRMUu+YakSXlBQA5b8ApY
gxxp0hL8OMhv6/C0XOtG0h3kFEFyI+aVY7GhZf7Rn+1NVDRZfF5jSqR1iNTCp1L8
kXWOJuocH+EoJUdH9OKdqKqeW+g60R6ggzk+uvtPPFSLN8FIHpI25tajTx2uS2fM
ELvq9WO6cH4ZuK62GckZ+pNUh3I0sxiVFmAc/5A/pASNPAJhLxTZexTaoTvElZ4W
DFR9udbsSju8Oip3uWWmIpt/X01xWYTcOdQgr2gC8J1xp0C/jNpP+l7XFXqWI9GB
Xlgwd40DHtEQWTlNIj+gMFqH95uSoGlKbGanLN3KtdMT9UhYwyTAGpw0zfXj3f3Q
PwPF3uUURiUhUH73TZiF0I1pkY+Bl3DbqhgZ9z09njx/PdqjI292uTZv2cr6zb2k
IiP8r0e1MtV3H8dahxzAhtllLjJUfrFpQOVgaeDO73hiJ5KCW67yVXldhFq5XhmD
AMz/iGYd9Ko8sxANUH6koum6pXl6OOgiqqXYEHI0wSsEh3vRyEitBUGrQL+vbPVl
yqlIIWQcLObhBNee6NdVmdUAWJmaxmK4U8iAlKuJvjW9oiJKIIjiHxzlBs6yDWqI
Kg57SCGXyrhkjkHcHyQorrKrBerbesplo+6qpy3VC0V0lmebPBh1B5njqqD7Nkr4
wj8ceTe25MVMjWSiOjZuXP8bVDFsBqFwXTHoVtOqg+u3pmfGvuscax8pHlOX0vay
s9BTIuaSHgefBOGek+nDjrlPsK5GUjVg9UuA5bR/nKo6JhKerKXEDQTH7GjUgmIS
JMIFXtB/7l+eKsMYSJ6WBan7Rgo6LM0cisekUSbrPC5Rl5c29qI9fpu5CF5MXsIo
9GG4YPIg6rB8hpDC+9iQmT7ObBdMnwmYJchGf11z1G7YYyJqGl+KVjlugKqgkIrk
BhEloWgeY5Kj5TsIxC8LsRro9s4ZYpWyIchUO0H9GHlDGnTY1Dzyz6YDbitQy85x
2dmeHxZ0fNNZ3MJL8XPUGsK9wbZe9MeKYkEsq/EJTKgC91ikUdijVzDJelLf6y0M
bQiNQQJYIwo7wmsfhuuqLd/xv2RjXlTxvYfi1za21hVqJjrWMvz7vgV1J3ek/Zwt
/1ZiJL2rTeeFo8wFEUGCx7xWqlGnC2iwSEIB2PlVKKNX+1tIxpv8dPbzFbcv8x8X
NfxFJrjQya4T1w72wb4wZzsMSa8YJR11Ouk0XPfuGsQRz1VnZD6U1E8RdGA+hcQj
xbThcnkIHiN3Yp/gJm+MpJWeuLiHnr1iDpWuIpB+7T6PXm6dwTqUgpBKq8tgqrfS
W9Q/LfmO8vVlK22K+DIroJ20ooZsMHdW9/VDxPJvERCZK0tOlVYz1BG3nie+mSeu
GOrP2SmqEWCfjV9/GZyaTzFob/9sgPY8SmOH0M0T70P3xR3uxu75j5W7f5O8j2mv
CbPnIrJ1ri13broJrQXR+3XseGI8Q9bYVtzWV1fkM9HCg+GlrzKWrk+Ctwa3MMy4
rJZPF3Qml3mNirFrAFP/xDB5g2QQfWlUv+UpG2a2FxNZFpBHWmr6bbPHul+5GXgB
q+RwPddcBIWnrHRGTyhDIB8ayHTbbkAjoV/2i3OE6RejUYVb1BvDPc90qW+mX5QN
3iBc7fT4+x+5gyNx9uJG2VxHGtnCy+gudOs7OxFKQJD2ZKjlnexxPI7o1+Ei3w8l
f41aNAsv6ekhKlJ6MPbCbSvUngGeHYaeNwroODTd8QbEch7xR0wabS+9EtLrfI2r
v9q0vIpB8Q+t9vm/EW6eBV37EakMUinA45iTCJOiUw4PQ2uCbvwEMqvSMOofX9kG
2tM+tjmgamGqW2vudSy8tPKgOYwdA1WZ1Wo0ggk6C1EzdZBs1Dg4KPgR4j7byh7l
y6E7ZOhuW6qEdhO7D5vmElK6QUdV3r6hd0zWU6U+57BvX+XeHimyTQWXcxXM7Qtk
KVdEqG5ZqSGe0jUXFUe0tKlWoe/eLFtkkjFdbkqeacpgtgyQzUzZyYTT6jdFaPqs
1Z2jygpO8XOmZ4tD96dBmYAo1jeYCOXDtOdoOd3njpmveWZIbd2QN06neDY/8CQg
TZ7jnZ1pMz/ccCiebPfVM4cBWd3EgykxW0KRFvsB/4l8W/zonm0agd8tTbjbR/BJ
XoUGayCnlsXMrTGK6vX7ECIckWR6L9s1oyik9cCdCgMofUZajL3Melufoa2Nv1sh
Efh/l/vgFu3CSlsyepZ/1FPQ/zFZaqpgi8jQibOXXkP0ZzyMD9To8KYwFrhFpUpD
sqQcN+ErlZH7RNxPpqyUO2NK5d2g/tm8WYf/MjOvwJubpju0DgPKFnHvtxbcAz56
yS86MlmCDTwsMVfyArfxGGczjVUztUgxbH1igh1HL+7mkN/h5OvBGdfX+S25zEI+
G6686zxEuHATX9zhbax0n3+BPeeOEM7nfVrNjYPvJXlkwXrCJQXzswJlsMmKI+Wh
DKwS2KbsOoCM+NFkuhLsKRE8DaLIz91AK0fSBvyGAiyF4c40QMfccEFHEsfnl4c+
CMX6OwKeBBXo6rwr6kFZlkd8GkB9trHyKJhgKiZvD2DxK3a/wN4887bRDRexeuAE
p+3GBQfu2pct3NA7Ag+omZtTru2K0r8jdW2aw7m1f9JC/6suUTHmPnNXSs6ZVaON
dq2dVTx25A6f5umfxQolbAuf2UdjVz8JWvMV0VnK4Ia/mEuGJJd/8GlTyOi86S/L
TyJ+HwoD1p52MGQDR8NV79b+mxzWmL13tFCcRh1SHyz3xDdAoEM+U/MA4V5s+SFb
qtAtoEe/bXQDdcmeu1dozh6SyAZJ8p/0Hm2smPeQEgqGVcqTlwL3SdxXr1AcVrya
VLt1D02xIOakJS3A3qKrZRstkQ46lGjslaVNat6gDtb6FmOpoqPu8Ua+yGF4D3Z8
In9+5Ftqk2qkTNqOTRDR1mrWNsBzDrEMRz0YtAb2h8GtQSfIJctwW3ZyhffgsonN
olLbJTOeaFV6T2NWoL5JKIrPNt8vCGS6Bks9+C8+vyB1n/XDpjxQSnoXLTfXCptO
v/jbrvP7dOwkqzx4U4tntWVRqSQJ2/EKXih/jscs5oMPPebQ1EJ/PLIcL60nOB87
c01ZZABR/NtwWt14RnYFJ+80pCSxRf5AibZ2NhBYI0PIzDocsRwYJrgDCVAO4BHF
xuyp6sNscqDVG640P/vZct+zI7mxVYOeG+g12GP6E6i2RsH8LZoWUWRNmT9XRDHb
jTyXSiWhYBLHNEr+NH1sz1uBLq1+3VTDi70Zl4Lg3lZLGFumZu190opjxqkAAZJP
tiFVk3lcJdpNwjJEvYuNknRpSgBg0DrLgR9ln19PCss9uwcGwHFSduyMnJ2bL3A8
r9TqIrJpAJwb0xl1H5/hKYuPH2etwRxRbfOPbtXKXlV0y1ssQjxD3pybBMPj9gvq
qmLx4oJE4IK3SYArJdiA1BiOP0eJnWx0ce4AyRSX/gUxshL2VEpwpLWCn5lY0vkk
JyeTgxKXEr02sQQ3PuH0XbFNY4eN0qR6BPAuQBIVYyjoQLpMqyRIYgfrtZnKYvhC
6DVTmOjByLxgQGb/we61jljE3tVkrs0VkDwcazO/EHU+PZLsRTrkw4ES3rCI3rOY
9JufMzNjj+OhI4SYeCS1mVVLtjHyNTM/8FltoBo10vr8DEb2crZrN5j09iSPVNQc
QkzYbXi4vcR0FJ7fZKuGQOpcYSGD5mFYdgdRZN2+IK/7b0AximfZr1mi3qwwFgES
WxzL2rRmmmFPk9PgvdS6+veaV75P8b0aebIkinR/nLst2c9VHJ49+xfYhYZDdRnf
lZatEd4yCEDaj4BS+nZLAeU519SIojBjs1Ep/B6DsMuuw4cXP3Rg0JI8jjqoZ/PD
YzE+g9a5J1Vqj+oycvDlaJwyc0i1qtRgC5Bl94xLBgsgUXz2a89be9QNp0hZXkvk
EqKzJ+mvQha0fcYg3y2y6ktFIqtueU3P3jdFP9IytRk5n3ksKr7qV6A7CyjYHZRt
BA1QfICR/H2apknaXWS3IXwYmNjxBiRQ4x7GGH/O4L+MMcx8St4GDjc9ih0cZxO4
l6/XatpnkINl+oEF5I6HA71rldaUnrDr2Unsbp0Dn8yYGQsFwCWVvvQUy4JfSIhe
PQmHvXchpyYSxsyXhY+Tvo0C7YfCWc2omiVK2EDbd8MPwQFMB3vybCvCj+vqXY1I
yHucK0KfhdHFj1r+07qiQjWRUgEFKf6OtPtt6kk5MdpW5Ji2VgO8g0ffKBb+K9Tt
HWtZ0ASs9kbb10aE1DPdo9zMnILg+NIe70etBA4mkhdXHoIDoIdLgguAyMlbI/aF
vr+1Eo3M+4VyAWfAf3r3EEXza7U30eB3qhgBU/BkWQ+CDipbSPDz/5W1q4PHydeH
p8CHQ6JpCqNSEyCpR2uGKkJu+6wvzUefuwG5D/d0o/wvM7q3jZkqB8xZFFXSvgIt
Ju0alAwkqssfEEfKVfzW0T2Tb7HqkBiOxLSpzj520kgeRdIDgzstFj7o2SFn+4tR
K8qTJAi6XazNBPVXT4e7zZO6CA5eW8N5Qjh7OtU7KNf5RxS/zTTNHzrhUxuL6PBX
HjOXAeH38oIgLCJykt5Etcad0yVMujx48Hx2DeuUWxVowQBMyms9DpIaP8qdLy6B
ZMn4KVlQ9h6lKdwP+8VoyUBLdiHnyVspzOtr0rx5kdxwdCmA6FHzgalS9I1sYm5g
hlaiV1XKQW4fsLJzp/C89CPug59XwdkpUeV8v860ETBQ3Bk7fHymKyImdMA8YCHd
wbBONCcLer0wwLjS1rXN7q9dH8SsiuGb0qr40QgWu3kYVjw30aZBxyeqCTOXxVqu
HVGHQWVzxWEpC0WVyd1rbJBEsRbJ5UD7MHsU1rtwiji0m2eR5Z+mgcZEqn5GUa6j
azgGPHXSBizarsYCRcZuE8Z+2hyaJgaIbofhYoG8kLLc0+Xir4QPiqOP3jGaRnXa
hE9okxlxXdI6DNrClFPYIKVFzpiiDLy1tM7PIucRbm7g1ptsD0OIDbGmYBJNSzd0
aCfCQ4Z0VWdDVw/IBVT4cEc/Mh5IFwz+lpWS6mGSEj47bsXenKxK43lXacTmfrz/
SwK1/7WE62EdYxeFOQAiAsafzdwIirq7fIPPPo9bGmle+McupWziBEKtYTNnFCxe
tHprK+NmsMOR2w/bthCRQtFyUjk/rqkpaDtvQxZC2xLbG7lnWOoYYj8PkAcGBHiJ
5Rt6mMkEsvO4MwSDY3/uSDu/6HnHmIA/0xTc45gM6I/QoOWUEWD7wwoDWbAOjhqU
gMBnn/SHcql4Q96DjMT7+rAaHNVCMLNK8wcwWFb1W2tA9kfygchqqTfarsjARj0r
xEaYADGIHkUE24UzErne85ieYKCYYct6+wDVy9ysXd98ExsEGuv46K+LLsqW4am1
k3ArC/XmXmI6vT3mlcCoCkCvQt/c8eAj3x2tiQmug6bBKgfg+kVek1DeYfH1wpvC
cq0MiKR5zhXHfc7oP9n4yUZ5NU0nWE78R1Bk74SgjO84QajRG13ULH/9ENNvgrLh
ugALuelZsEq/re+RTkCzWYV0Pv9CzzriqkAHAB3K9EdwMnLWiGqw7Js0/K2HbqOO
l0X77D94hb8UUwTryGSh6AvL4E2JMkpXJNrSNtHuiusAE5ZPEvlUjQlL4uL2FMAq
abbOskAVLXa+mDRmy067JOYT9bQ4hLxaUlcTl+U4zHEpOvFPVdAsyLPdIf5M3ZrQ
nM3RuSkro/6X6uO1h33H8VWps1yMrNCvz+0XQ2ZdMWAKNeyyv1mdsE//w/kjhoWa
J/oD4ahC9QTHIvXQeq+Bw/k0xALguEf1lrDrUdLdRptkRbpxfBTJPpYzKLV2/vj4
ibBl66tZwd89YRZlOLCJCGQhKi703VbplLREF/q7TV5QkNsyxTN2+7ED/ew3/49y
+H24IK0p4QRD8JZXCxGDbRRIclCprHbH9Q6OIeuKgpy/QwP+MMozBxfk9ZL52OFN
6//d/WNeFyRGyEVQ1Fd5udfmIwVqRH+fXceH10v+M6yhCWKFYkOGupjT8Kjg7pQb
c93CFbR/MaRgKWu8p5TUsXP+oRBnZDDrO23cxSn13qmcwAuB6A9DsxbsQW191ZRT
G0FYhvZWd5eaiVl2W3dp8aveAVTycFy+yBO1WA6we/ThmrTai9nj2NDPyDcaLkGQ
mkC0Gzda0lIPAGl9S8PrldfQJKNEo2DIpiDZ5odAF4t8JGehW12tEEkK/X4pViVX
eoxYRLL0Lgdhx6Vpf14h9Z8G+bX5kZgpCOBLFtGQ63SR+ZP4/zmjaRc7jhObe5Zm
cq8YhSaVBSIH6GV4PkTyF4F3zUrA+2n0XmC9qqYK4W0NpUmKbPhYw6lKuXnGpbBW
9Ce1L4aB2uLzsVTXLvB/DblU9mApyl3fddI7x6WsrUgmXwosXNPUAHtkbiHB+LRq
QN7NoqKDXdDZCIdJ3oC9OY/vYaAxU5Qie/umQgt2JKsuMV+9HlbjFr/JdZrx17q/
k9Zu5xwTUchIOPXIYiVYelPGERjLG3viGh3Knbr8CIl0wNj716GCgyQnxiSRArDa
Lltu9z46cM4XTreQ7B8zOf/CFoIxGzAiPCDxqsupRhNLZ0gkpUSok1+OAgG8z3vI
ffXp2i2dxiOJiwyaT6JvP6U8hDD+InmTd59VSk4lCHcXDQWycD+NjeGzu7/0F+TX
oafR0BmN74CXR7FTGnXwGMraHouW0JLSen71f1Hku+2Y5SzEdqPXxsis09X+kVSF
aRCy/D6mkrnV0QOQjtZoJo4APoBjXzbCYT1DQ5SQgxWWRdl5zmOSIX4TVZ5chf/7
6t/aHjEDv1xSfWtfmyYd7XYH9aa3GedBaCYhVrCL7SgN8z+52IQ722+ZvVfTuZmC
T0bGSRaiqsBlAnxkmdRg+3hPNb1H2WZTQ/MTnPyBXbQWP7N907wMjYWrIE7NfpuK
BHO/NPnI5QyJ1eYo5FiQXKdQzjp92VZXoCsvtvSipXoPUByyZVTbltDBKgln76iU
03OW9oG1sRdp1MVApvMJrku3zPp3RWWaZkPvKbEWqWAw8MZGiOWKfolvFvjqtsWu
n/I7D6+Y2RCwv7zgyEr0ygKkzO1ORmSHzP2BN84Xa8BXhQGmeYQBii0pzyXZpMD/
r9mRaiQvFAPYaNM6FtNDLqkGOOpwJ8ZH0rtgPmWO5kkSP5x1sJzBugPdvWFwv4BI
3HF6IokkecKZz9VD+O6pEyx9sDC/G7Bnmnysj+9PiXrRKM92L8tEu+sPqUM7M8Xu
+KXnMizjitnOG6owHun+A4B/fayVJKreEPs0nyySrwDUz8mH5wlwjQ1UT8k2R/ya
mBMB8WSVSenikgSeUvmnydyyaieDKUfPNQMYwg3ler8ZTRHBbAm4qtRKbQFl1x9U
ZxtraDZd+weAwdkO8kjh3wHi8JeK1o0n+2dbR25/IIVba7rWPBT0AV5onjc+gb92
dmpWGPtEVZnQR6lb4XNMIPiASL+lyud5zUJ8Qb4Cbltpq/UKEhmTMPnMnZrUrnxQ
L91p6A5/Yyz9Z1GZfwlhnpZ7EDRtKW0KEsVkQDEkwfYiOvcXryrO8XLeahFKFyGc
FZhuI/7/c9dZuV3U8A0IcWo+I4ldHQbnrTxjCB82Oe8Wj6DS+p7alrf1HjXFC9jp
jgXiRbv5tlnwjuyFrT4Zub3cBEJ5zAWz32BYsDNfepG7fBFuzRoIuMCSaopvo007
KF3d+Ush3pLNJrsqmbVr7JFPNoodCdPfQRKmfYpKJcOUIvnXj4irvmFUT0nBp7+T
pC1bdYnTOzxD9jU6Nrvsv6J/dSNXYn8hAYED/lv+vtim8YOZpagk86eyJIDtREle
eSsCVgTHLB3N0gnFFjYo4VlwHNvDpfGkJWma3TCdI8582itaUIWWYv9j0ciZVpaE
sF1XB2O5985Hchw5A9lfFpC4n5ZQ+EJLt/o5M4QIj5MoC2zxlKSWmaooE/nOlxu9
jXr8GexiOjCG4o+Vy8xfSBuq6aLWPmZxDcfwEBQRK16xG2oRIX+Qsl+TcFAPWYFj
O8E+sYCp/++omqtE9ujPwxuLRmLKWZahRbJwDyezSKINidaPjO34o5eoKSH+AuJD
gzW9RKb9HS9DzmEiglutNj7wQ+nsItDh5Tvh3MUnS5ZI89q3Ac9d6PbRGw16hmke
6TypDh42BXe441qlZXb4pOCDar8EuUye9pCw4pHbGeylSk5NU6b/0GUP6sX4xE/B
xtDZqTy9DAW03aEU3ZCrBRo5u2sw3/4L0eQYnbYCPdj1NNOME+GhOYfHcltKNUD7
bF8zhAZQ/arcsh1Ibm6hjqfWyR+oZM21GT9Li+lGjj4CLI5L+IsNSs91zqxGYP1v
mnVdavHVfV5op/WhqlUsgjDLeAOZeoFZCzrk8j99v0Sb6jFSEkgyKxApkEFTb79U
+C18ryzZuv4mCCMDT9XeZJ59kQwifG6xSzRH4S085m/hnRrQ2kq0OLlEZrlIFD+c
eGSlhga1dutz3kmfybL3vvw7nzlxuvqpXjjecQJ+dLSqSY/4kMSx55QdUNvzY3Bz
pcYHXCx1cozrNWeFRMq/NzhkJa1ehuDOSvDUuoEUdQSdPNOUpX35Ap2vkkazeOwo
FJLf9rGBH3xfmg6qIUvfHCFJZHDR846IWermo1p8ZU6sznXzuKGADAeM41btiy1k
3d+uJ3oOopH9i4WJG02zLxLGFJ7RvylJy1X/VMHvCcGzWlVkWesAqIP0ddoxAdNG
gWVZxm33UE605YFtLvjeaEJ+LlfFS8aM1R/jE9T/tjh/FfbwvFElfymDV255G81T
tzjjBaRLxQ/VgmW6Y5X+rLRz/dez+goZLFXn+dJuo/F7D9TvS9A7DraM8/ADIgu0
lJ+o6JJqQNPRpqxwSdL+OyoQy0sXB4JslcA+ZwpoxIX+WOFTZNqQ8R2p1BeDmyVZ
IbsNSg8axnWbdRn3zXvolNhmOVOSex58VhW8JVKAZ74ALLlwQT4YIMoetLi6xrsn
+lF51xNDmgJl9oLzekSO/qIqsF2ExQx4I1WiCMmMONszp/de92MmUEQm6hyIdHjg
POUTWSUj/lD7LfwpEIMXMJo+7yL1CzdLczIGka+JhdVKMgi3A7InD5c0AiL3psRM
mwOBfPGGbTt/jx4oM+SedbvolmAhtsJNevuuJzZFf1B8ogd8++8i6BRJ7QXquGtz
X97IvNax7MIpcqcCbJwNn57ftkz2NkT4LWIVVhcwG4LG9exhVUgRwxApc0qHQ458
XHVn6VJmlzVFAOIYKV964pGiKnN4wun+TuhRKxxTsSotOKwvhRIbVAcAh6/RGntN
Xumh6DWV+/L68YQxNl/abdyMK8LtLh4HA2oq0nl6M77jB4uEYEfc6IyWowQvznhG
Fz2sjpAjFu9wKROufv9oKqf3BZ5RH+YCMJdNaDaioUro9dwEf9h4fPS3epXpSjEk
ob1DdaADxT8JE71OgamRxjkzhD0cNOlOcmR9JzL/CV+RD0U+QiSJpNWaQTjPs+JM
V22l02sD8wHFO+G02s47zK6t6bR2V1ZlWYFTUwwMnBF/vXJkwpjNd2PX1HCJRZlX
juPa8Ysf44FXe3eV4sD4Qlb8Jf75qNuuFUp8Jnk8/Gw2ox3cQGXIs/Hsv/0+Tg9Z
SXVtn1Qc/dUBVpjiAtEltKq1tcUV8Dur2XciIx9YDvsVyvlC3/LpdfaMD2OLhhlR
+zjyG2bGtJwFiYKR3eh/Om1B+DYCNQHYfVIHBbm2NY/I9X4jiyzlWu2W7WGZGrhx
E/9G0LqsSszD4+d2dSBHcmvADvL/4y9bxW3ImG4rGth5nKXKzSikwlgfbQhVYYvE
1tk/s1zQh52sQH5UGDxFZ9wnHxplnLiKgOBqWpZngvoV10xviq3a+oMB/ACHiBx/
bABT/CPkThVzUQ7mFlfEnbAbUBL7GLl7MMBuMakJDurhbRltigP2rS47gJkJjqTc
qNW9KpZVgT3+D/9a6wEGD+7RirdsUSFA3DmIHkmlZt+F7Mch8Rlg9esrtFojvCpK
TPorUowVOQUWbWvx8MoeO0SMSmrXJVNpyGP230XPqjcNWQs913IJMgZ2xLX6EM6Z
T4vCuSIY4bMywXKK6DLapn/31U93UXiYR+s/cRVpB5FGc5MctQCCv1lXC4/85eOy
JDPiWuN640qyT163RM8KfaXUZEQLtHqTip5Oe8uo4psum/vnLPGA5tzvAuTD3Alo
iQEmHxTi97NVoPpgFDRnvEUCDojA7D3gSLKrsGScNQ1sWyghOdT0+m1zw/h1A8aT
qspx6pklSwmUPAYlvWe4OtlnQMxolhKiKY9Pyk6MDhEnWVACpjY6DcKFJnYi1NMr
m+4aQNnGAtko3206ev1qZEGoeD81zOyx/XQ2qefMkivkjRbrm1fg6L9G/Hxe5DGP
7zz0kD4vkYYDeCq6ccBAvfeGw7/AXXDLg68FVVvh+InhzLwxZWKoQH7GzxYrYIJZ
G4IucZkYLQsBgqjygNIhMd8NebP8mGYu2k71iHR5u5sAv5PwRlftXTBWd9OBvO3a
PQzPHmdJNXQX0lDw1TojCYyeAwCPPnUNBsx1MmrGYG5f+2b66zPTj5okh9vZmMTB
+uxyCsEZaz9XEsJL6TbqTyFXpuEH3IyvGWN2dtQAnfZ+IZ/eX0ph2ltz6OaevsOs
y4v59jedXBWeXyawDPZ1JpERkaAMay9IrtEEVVm2FqUw4Lkh8VmBukD0/PPWAStK
1F/naN5K26+aFYLkCoz3qppqkFj9GTCpAKFTLS/Gxh8eFCXUdni+TZObQh5wbMDU
mnsz2/oew13AWObTbN9pVj3bWq4VhnitUpUZMaWjZVbgkk1XHrukCkHN+nU06bHm
fZ7cSFQU7HH34B34XXXNgridrZF4pg/j8LS+uY/Ls/3PrTTo2arha44Xxgg2/I9L
s2Iba/mIRz1BTYoV2AssaAyFeBqmq47sWWEvOZJFuCCwvH8zh188IGUSR0WCKUKl
mpcoVINDoVFcpqDH8fF1e4QYB66oz1dYvCBU3DeNZNmcQ9tWx4ROLETx8Znqsc5R
3UeVJClW/OAmRjbZYJ9aM7N0f+neexg0KUIyG79qVdr4sxLGvpGKby4GDyp4M3TY
xmV4EfUECUHq9B2SMX4ZxDnSf159m2VcrwxbZun1wF6fqh9BaYVhDW6+iudICztP
2DE5682QUBJFtSheqpcUgLhB2VXN6AactPn8XQp9659prCdaeffnE4y/GHh0z4MR
QBpjCNnQ4bsfanncvUIj2JhCfwJOY6BDVxEZUbi92s4xUD2G1nq0s+zKTcdMKDHD
GDNb5qY8VT+Ii2h67Kc/vJ2CjQ9/0EBqKnc++ptXAergmoZ4IBtSRuiavaiSA+ku
VcWFdQnqMhpdHxsruC3zC3sChpenFE7JioCOKI6cMgY/KSqTbYLbYZWhCwSjAUo2
34mavRfndMSH5pdZVE45YJOIAeS+QEwsavqwqJGgAany7g9uxc4syhW7CiDjb6yC
Ob3ZHCHPLbiSryRrw4SoHHQGSzIjpLpSzt9n08tvp1NYAUMoBytxXlGZA78zkB8k
MHbMdfa5VVDehHVAIRTyXkxQxgtYVIO5itxlfeFPOlU/fWBTD+LY6zY3mmo6qa2a
JME9q0iCIl3RDcb2AR6VTMJ+k4Ud8++qPLIYxd7AaxR+FeJZsQ/cKIwlicMQbGEg
nR60fCkCpMAQ9FzqnVkdAD91Wigqu9peC5oJ44f7GGJEUJDrBYq+YG4t8pTiYCR6
bKgI2MG3jt2cR9mqgCLIPJvDhctytPyBXSYnk+/Kl1UZgONiD3ha81zpnRcbnypu
Cm9dK+9QmAEJJ7LVqOlznFK3AOEHaCY8nUhb7zQxFGU3VolhWL2s6HkjarYdnbU0
THarqeXFj1mTsQ2HGg6XoS3dEF1LDhWIr8s9dw2cXggLY/zQ6tJJ708XzTqrJ6pd
3xW959wuHH070xVpBYO97lOd2S1z0rGBRB6uBH4b5sTZ4lHejc1No3hFyjQwqK7B
JSWYtaNT5d45y96+Qrw8Q45XOt6RYGYtMtC0ssE8UPDZDPfJpF8ELsBnJi48Amvj
GSMQUhHDT4laXMvPPV83WT/OIjCUbkRrgmX8VzJmiQt/ElR/MSxWnI9keq3leEeb
jgGpU8NOKBaZrGdY8O0O7rKhLJar41tdEs/iA9VlDNMf6S1OhxtipeULbjTzsR9m
8EjiXDhz5RX9hAWD0HOfKQzUql4QeH9xKlGSDQ7k/BwMiqn7NXHWSzQzoWfckR0b
03xhC+g+dohhymIjgOQa/QsM2bZ8eilqcpGOmM7RAgTLiZJ98Cyr+OLhXEZyN2Jn
IWcZv+FQoi+WT1L+RvG4gLwUy7MEUm1J69GiyXpuIWHC/TeWDHbhKai08t86HtDp
1pfIPjDsvt+Aj1FsUi1QMzOlxDJrhVuG/UBWCPKCSxS4BMC1TMYIyLEYgAOj4cSr
qHOulN0k2NwVTybmvIcoRA0WoLSYKid2piHFN1mA/ORh+HI4IHh8J7JoqJjYV80P
`protect end_protected