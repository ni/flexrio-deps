`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 20320 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
DBGZtUPdvgnvgIFp6VMrQUDxmA4KAY86NUjqZUXeNDN3xeREYggpl1NeAq+adFQm
JFPQQogWULhLhFERIjxueqOnk++uBXEH3Dwxl5nSOBuA5a8kOHMANEb3FP3pnkFr
pzT9c3JY8oodGYDZ3aDpDApi3/7g1uY6jEELRO/rl2UB0wkgRV0CaHuY01WOV3hr
rpNYiT9+WLUiai+3CL/ji5Y7VXbMLPVq1bK9vYfOugK8v6W4US2i+Q4IGrFAKHlm
F+fGoBEUiFNDLN5Ipumj7nXGjmUJ3MJtxDh36Iz43QDnUxWybY/BZ2He88UdKCPT
g4Jqhp/caqiT65T13nIa7ETRtzkHcaIyWucSUczelX5NM/Xu3uKT1ykWtISeGCqK
qU5MSO8OHxdyhx214l4HPTqBt7PsLbQEDKMQOkTlm3zjAV7sNknQZtv6kxtpcG8k
fqXj9Ve4tjyDfnK0gLpHk5cfK+gRHRtVf6ma1IL9SZEmqKe8hwEImlQyc5LBNLWr
UPzpK0AOb50Girtb44zeUPtcz2VL7eJX9pSX5ZenLKLm+p71mYC6Co+rj51IrdOV
MHaAuk8XOeTFJYnCVneP7/YX0lU8OYu6zketJxUQZrBb31FPpun3W2pP46oV6QLk
v0kDUfHbeS2DJZ7cjMnK8CfmRlcZMG12DzMQ8XZ5Pt7cJlThBso7sjHU3mQwvpVm
PCdp7lVrq/hJab8EYSEsL3r+MFwbSwFisXIlQHjnik2PV/mk7NiGts8BjTv/Hw4W
0ECapl8LRPaef7WHCH4yoVAwT+jEEpixJLRcJUmTxoy0+oKujToPsbDU9drKHfj4
iTQ0Cb4LQPv/wmHusC4dnqzefa/3yuKAvO8tuyqhUfY1MohkQDzEjw9D5Rw+wj2p
MXANgJXJgZcPWbriUt4+Ny0d+s75VKOOyUI0Z7QY2Nek4UsMK5sjhn8CBdBRx+Vr
RstaT1ifOo/njJnfeTo2Zyws+LmQN4VPkue8dJG0dEubGLJGsJOXYf+VTJ3swY2K
ocoz8wk28mCb6lkSxfmBDyxVUMpIdgCqsClLnUECvdtLNSaUkQcOtb1qGeL41Je3
uUcBV11uHSvaACEyKzEZ4C/57ert68V3t4t75H5CDaiDUl5v1vRe21OzHTuw8+1t
NUJK65Bc/z9ELtXFFyAD9vvZh7V0uAnPEBNelzSOZR72hqbeSV/ycaCL2JBEcq5s
cabmZxUljs8stsQ3ryQAicKOLzdkxGmrg6g0CnIeOn+m9BM1t3zyRhNXH5TLsxZf
LHL2Fu2K3wHmNo+brBcuW7QBxqoTRuTdAQgcoTWa++cbTuLwqm2DN1PvFmc7PRuY
YEIatYQLGuZu9IWYj08yQb86KkT/RTGqZFRT0x64YjAZqLh1mdDDyAp8NQ6+IRRq
oOlCKId8JjWRf9O0OsKEiUo2ClS+b8aL9l++YNnxD1AaJBfeH4049YhVIJ4YpVCG
31QRhXQYoigLjW8VU5bogf/PUg/3ZShAEeu0nm55UK4v1VAO96BmMUuYp9MZnKa3
tefyj/TQu3c7VAKtPQ2iqQzU1/DFKjuaeV2Fp9SUUOd9jCk5+mBQ/tcUyVFE/HIp
L+520DylRAUwg/0ub5w7z1wfOuUGGwpIdccwxQYFuM8jOzuQ2AXVzor61RqmkegO
K3aKONX8EeMNZiV/yWxtEqo9XxNw+Q5oT9K1IHzhitiAACjqlxbarKg6ipA5sXeh
LcCqjVwH5BGhvhbKEPWkVnXwP5KWpt2bVPeL5CukJj7QUq2E2Cj2tTn1nL8Fq+ai
MKUEUPLFwBHzJosX+rQ+HvUudznkEdy0lNqE5UhfcX2xeijy9+VvqhvABRkHxYsD
5jOyxprHAX6GE6KcFp4osALGAOqJH1k9MFRkpr0KN345c6CbMlIL6ldf1Jowiw6L
6FqpH26+H+HwPSkymvFE525uDKx0S6ALxsVZVUZ14+alWjFIX8yhg6HjJg2dXnJo
bZOf9+SRgPpeqCqMeuUTXJB4w7BtnpRmD2LT9U2LGB0/qwakghmmkcbGRUao5U8g
LsRfU8Rk4TU+mxVcAhO3BaCpfan5L7Yyo6fkH6IivbhLqDbK39BsOuyoeirYvTFI
dPRJAIIHXDy2Q1pPVqi4OGtOYKdF+bYyoBEoxEvlsStY9bOKQ6I12vGuMq7aAY0x
ruz/Wd9ysrPDD1cU+BqyYY5TV1obrMjv3XXjo1HVgd4UwWtTWtWK95SsiTpisLq3
GNMqy+ZJa1TLfVBjWxOOiQU2BoTfp0lNfuqQMI2Iw1mQAg75C5UxSuKsxMIYuENa
Vtp83QnvhdqyGw3Tw+mXKYPLQa7HADpz8Nz5qjwDZ+yeQy/awsMnSPxVCqp/bdyF
r26ZK/7NDTsWZWsXAW1YK1+7PSKzS9Sbnhonj0VjcWi8PdVPspNM0sT3qsAZGrSF
7USDnt04W7w3wTV8/+apdBemgW2Y4S9UYCygrTcf9YRSe49BOEzdH2XMmuCrWcC9
ebZQA98wh1PzNtVWZxK3b3D+fLPtG7P+WzyKSz3aT5aCUzLXxuqKPehO9DnYz7JD
kNIIT55IEy1GgB8MMQseJEn+f4/yztipB9dTsZcdf66ha/1STk0/bTYPBz3TbmaH
/zRpebfth/wC+kPOdwZPUFofULkoNhQN/c6jN12N+xE7bD1KHac4B1BiwAIh7kS9
qQHTJ6LK0i4J7ncF4bumqTxeSpc5OI3CGJfwPqUw1Jqyi+Ugfepscy6MHy8ixBCi
xJCNHqEEeuJaxFCn/iiwFTA6gjKMfR3kecJa81n/EhzDEBhwIFNTN7lSi7sBVy2e
MLqin/3urxY4NF7c/OlxzZ2tbJCm/6tQiK12b49WuHS/+sZCU4KtNZrvoFAuWdOl
t8s2SMmPZizp8d9NWP301lsAeBaFbyCctPVrL3bf3DxFOx2LtOy0qR4jZE9YwQpl
pKPhksAfaPDthEcYkCBA2GnnoPlQwlXvQtxOVE9p+it76t8cCm3UCxNMMiSni6wk
bHXrn0N6nblkVY00Ve4VU9tF2MfXFvFCdIacRZ9PM8+SORRkclEilhkW6AFjI0BB
jhQo0ugIuL5+1uGKBCDJEV9Wo6pvdQBFU+/7ufAuPO2/YDK+q4aVMAZcgf9wzB41
1tKd0HlBVj3AovKCCfBpD2HYcFSmHm7tXoj478HrmT3qcUjtbavnI4C7y68xMxFs
qL31KfpmUsMHzgiQnf0zkYI3XCBzx7W6io6kRW2MhJPUnBh/SQSBkHkaS/6W7Xqz
SqxKqFdqxCGYqUhM+2iRT5wWI8RCfaMSGavBlOEKgnVkB2Egy7laWuxi05Xsx4yS
wtG6rqBu1OPWCtGACXZ5qmyWG6bBqofdyyr9mByXI6fLEvDE2X+c5OT0BXXZDE4v
KauWfQaoVYJ7fzDNQ3QCphZgELu1LjCaLbxWqOhS5jD3ouDQIRKS1rpv8WwKxvTm
0uOpdOVYbtxTB8MYJmc/l1GnMYVFrtR/IW0s2rS2ZxRoifMOSNB8lu1bPTRW0xPG
atQe4mAKXQpLlGVctYyBVse5MLd7A9kkdowOh0DMQxZHFLiEmtacwzLv/whAZ2qv
XHjQdhDMv7/OiAlDfYP4pl+HE/9+YUtlRIjknt6WNzhko9c6iDgwybTx1Y/RLbg0
4ib/AXFGR01gZiuuJ/4dz4/SA3PLsbIv3VRP2qMpVGC8ugxUrIwMlNR56tKaEl3S
iWQgBGwzSn9eizDWP9m1++eaM42R+XfzQuPTHGdH3mhd1BV2TikZRE0lDjhb0cjY
ArkPioIWgrWCp/Q9WQ7fcI0xSJKXmGPo4aBNTaZP5h+jSwy1om8ZzTt7f7vUl8Nf
UytS04HUVAbLUGP/pyp3w5jqSBS8xnpfqjVAN1aoJomUsT3QO0gKkA8GVMCLmUgH
aAFhcUpgMQgFBWxU8Zc/zv8I2z4MNVJCNJYrbkO4Njcx/bSz72s+qzPZ6OmYt5He
SDJKEJpvXjgp4kryR+73vcBlPIFo7HB+ATdltmoxBOzkGh/xHLlgqCfqn0unCaZV
KwsNyxNUGfdExRyTGO7pQUdBDbattoHgj/heYXb6C7lIFTkpFRlNvTtOHwneW7J6
14bHex/4Q1P/9ZuvHHyfCNubvILd0ycn1Q1mXkiJkuDvMh0SIZmmgeuv0sgzXu94
pdK1QE7l1VgvISAeBMMniSBlYR00lAvUpYomUsIJ6Fc7qeA8xj4C1LRKr3xxZTYM
fMsFbafnTJ+shW6EVD3JIQAz6b2ufoQyH6COm0uaMaW9T328A2S+r9Zqt+K9UA81
10x8FEhStvb6k6dggT3rT6rkM/zNbaa+DWNSI4HmsvZCdQr6akJc2d1Bs/CpwzP5
2PGI2vho25BACKMOUaMSR7JHb/D0bd3MBgzEzu08PPmLrjR0w2ylRDmeUB6IqpGT
gv+WsMmHf6vWTQGsu+3NqRlRpbm6SGY+hGmYkVFsAd7gV4M/1c/AApKoi8G+ToMa
lekiBVMEaMzlHJGMkeltn5hIuvDTgR729N5AeMK4hw967lbrQJUKZIO8qfc4QKE8
cIiJSj5CNfoY6BNcwVdXx3AJcjj3z7HM3giZBNsqaGhPyCmW1XP2i9mJHwFQtm0T
2toS+NEr1crBUAy7E6koFKHKMhaR0+ChqCwoaVnUw3J/lCrcACwmKUrVUcLeiILS
cSX4jRN7dG/rCSP8X3mPkFL4ofyzAewCksFrQwaZ4gdZZYB81+0Vq+mZ52l2EvVu
S/g2H1njpqcmkhK/mamwu1qIdhVgT0Gi94ohvR+NqeyGWCM1KjebyX1GbudXRnw1
+Xc6hQ9TpB3B57rI6t7gbDDUmBWwA8Roc1bc601V/uwcTmaMZvSaQEW4SgPA/bZD
PY+FhiObRbd6WOL2wNc1AMP8ULlXv8grQL88q1Rg8V2Bd2POZlsdDg0anzDeZ9Am
CeXjOBtgGJadEgk0ifJHaw1/5Kzx6NMgOCAdknLCFJyfaEL8dBT42j4MegCvtAar
lmUrBnjfrjeCtoMRVrteM45PWjPgrc9k1dn5UZadVjocfnSdtNE0lDfxNy30WLkz
qFZGqYRVh5Cghng3RtMALHWdajI3SolGc0r6JzW2LAoQJShuzvKQ0C4v/vv2KhRF
tUnxCk/ZNsaSrtUfw5mrEQzis613SaNCbmq6ow+wamoe2prEZ7d6IHIZyto/r4id
Q2ezljwWLDeI/x9wioL3h+Wvr0dBtydwvEzvbkQrb2ypVzaNJtlJUGa7dgSV783X
K98QmxsetwYdZR1Olbp1pKWgBmXVykVOUmNP0cG6Rdfy9EyT2E303dKZoyanC5Ky
ZJex6r+hp0I8xFhK/W0Dh1EG0bN+fuTn1/0QFMT8GXuvhBgfEMjCYJItQ6BZXiGx
FA3FUIV6aV6PBUE8oQuE7sftIfytNn+IiM5wDKEpMy79Bc3yfZMITkotOZ02x+9s
/F8L5+cB0XF8Ne7J5mXKctxX9gLNMLho9hVUnNZZjHLOovZBqyDNJG+aoJWXXhu+
hEqRt+RHCvZBGoNE3yo3PuWAY+D3jwYmQmJEd9XG9QwOg9Gzn504APY9zPBvK6oJ
pvvO5DPXBHS/USws1iuRznPFvC24cOtH9HsfCn2IrJqerldoS/egqepo/pi5aLMD
8/rZkEuAaYTvq7QwEvNhat7K57F6mMaVLQBoGMypvq+JGnocdH+vUTwyEHJ1LQG0
3rmRjFQd+8fgGjazzo4j8IK7YqkQM188lDaCWxma1+rYuaP0mPVyvB4gM4YdZeUo
t26aujcNAger4NqtWKgUr44HA0AHrKCpidrsz552gEP7WrJDkXsO3kSvC8bNMWK1
mmiJEVjnkWKn77FpvrI3KRqo0tO+0S3xBpG2s/qfMOviwRQoZPe407VMgvEdMf1C
vP+0QnH8FBJ/maWfVGnRYg40jpUst8E7LNx27n4JTiytkEoLoOHx54VWqop0MlX6
tw4X4vp7Su7iLOLFos/AplOPquj8biBmtjIoCL9B2jONwxV1zIjRZVt4bQ5YwyXK
zLDrqSY/RmTR4wiKOCBImbbDrDrvqGGe5ggSvJK8IL3T662GeJpTh/drGyMo0WYa
ZzjhQwBzS/ZdHXydxZAAFEHk1GHt/4jGSrezHfoKiWa2GQ37P0WbcGWwENtcJTEX
T4TknnufzC3OSJkL1myk5HAbUQ3xspkem0DU0KRfaduU9jsOGsLe1GnRZAoYF10v
bvffZQ959aIokqyIcumhCoxLLR3ARDVt1OqOz4NPNl22L3r1Wdz8SBqdpiiwdDQ1
M87PBHqbg01NtnUT6SsoplIslliEkWc5TbPOAcjyZ20jLkFlI1S3YQ3QF28gL+0a
jNEEPvqmb4nvtAxFJU5GGv8/owwchGnvZOqZKnZWy1wmezSWZ0LXa+tGoqt9k9Xs
NlBOt4E/aJNLJ21UU3FwZOlIs7RvGocO4M68tpaQvKaONbfDXpbOvY93H+MWrp9h
M8CDyKtfPvKQYZXTX6clwx2JLb9Avq09iz/phTstzO8zt3/HRZINf/tF+kOO+c3Z
IBXBCjKxFo/PSxmfEc6fYfE4FaECIQ5BATS8dXp3RLB1WOI1ZwgRrhIY4WUtMqj5
3WlSHwa8BJf/ErFTtzqoDJOJAPF7yiXWDtbH5fRv/4eTCPk4igH082fF9NPG/1YX
Qqv/tzB4/xusYYJDEsbku6QGEcq5OtKmA9jGh4iI6JRteB6V4oY3yhtgKypFE/jN
PBFAMy3Hd5P/aGU1u7dKkAOij31wTpe80pDIkm+fHBLi089mtFIL27UzoWxWmfWd
O/uqbx++2oQSRKzo0Fy9YEUhiE/gOyaUkDB4tXeRyFkt7CQ0ZjzNmqW++r4V5T8F
2NJkxpTeM1EKFHX/nHZhPwDgP/dm0BgH5aRR/zSWO/g/edxa0sksDAsJYxPPJGXq
Ls89Mmk8CDvKkkkxhHX3WF55KeEMGTLhNltLLAckGoAhJLLckvEnqGTXgqdfq/0y
RKujgAPOJuW8DCod3j9EuKFHd+fTwk00OTqWQ2wtLde4v728/rD5OV/sD8OjJv0k
ziVd/cGn72flX7QZoA3Suhma1gMJJ6AMSUQ2Ccvz4AIF5uvkU26ejUkskgwYu0ly
e2Q+wrqBL8uWQr6fl6RlXm7UmiEN2z01XVywHgJXY+BAOaHXG/hFLCFTAkkEnb/b
q0Y46UjYI5tSM2nwfQXIVUB4NBUClXKCqnBn+CV9srC324Y70IGCf0LCQmpr3yjX
9gHcFX6JBSfIz4MP2HRQ2kGYS9qt8ubW72qcrZwLQH7sRXDqXVBuQQrJxGUYaNzj
z8xOGvpCHXsbZRip3De31erZh8+Zpa9PK92WhIULOfM1zUcZzwoe1Ib9XOKzulSm
SKiUS5L43zGr7b9ubLiYwPJNNl1rY/KHJMOd4Xekjw83Voed4wIKgbOXUEtTnEmT
CrHbbb5Fdh/7Hf60qYI0audec8K8xTc99L/T9cgVOlbI4plkYLWOF+3O+/8Qu9Eq
DlGXVDf29wAN34J4wSryv006ro1sRXGaIePB/IU3aNAk4GB5j00j73JEIArKQ+RN
z8JBpdPPG0STeFIy6npmVwrcMTsz0GqeLeSxpu7fMjo7XtiXrh2xdKUPK8KyJj2o
S1SBI8EJOm4IGMrz6VRaqlCFeyG89UaTwlywI2GiowBw3u9GMoCQfsechcHOVfSm
YJX5b/tnx+58FK41kO7AgTJYkuSZfKNkZjCF1oAy8DxlVCq4fVl3uDF7qkW42ep+
oSanX6LNqQUy5TtxdKylbOgWwBzgDd2+nTEs8FnqOsri7ykNFre2J9yQi8Yla8Jl
k7MHBi7rnssYDFCsWhgE7wKvngI7TNQaAaUVioOAnSXyOhdldXCxpEqS2k09Pj+T
7gr7vOzajprBFQz2IWORTXT1g6XCvcm+lWdbOUegNblRoMehEly3eLcy6GGwzsS2
Ha+FHe2rG98/m54/99QY+4/xW+6DpS5VtroH04ZseRJKZLR1c2zd3cwgBhwvqW/Q
hyioKp+u23sw/Y7DKdIBrtVWnvkA6+PTPM/rANFTBafeOJwX3ZL22M6Y50GFzjcF
gl8IY2wLvelToA9ZWvq1Wt+BgulHKMDGkwFn1ufo16GL/K0hwkc1gRXpFhbrzXJc
Bc+OnIPyOzrrylD0CXLHufmDqT3KBFBpLI58LbL9DCo4LYIQqTakl1v2b0TCvLdV
+a6Gngg4DLlNjwFxMhGfxclpmzVhMJfDzgmxUOA5kdA8HMadmgASGBDcfUsVRG2B
EX8GCcdo1ZigyY+AjJjfyUN0qs9sVtm8TZiN3DyuQuEPnlRgrd3Ve0TpNSiDPbC3
MBvbImVUH5Os7ITVd7ZRGhQp1YJCQjOs6tLm9bK4WDd43B4bjj1skhDV1uwfLuYc
DXBRk8sSr+uDIQ2DscSeIQ7zZQ/OOKWD1cLiOADMFn9t5RTnLPR+RQvYqqsXdaH8
SthtdA5//fErY3/trQV1hq/7aChKD/YrU1b3P3XH79qZIdp5FvTS3MrxIbBKxydb
8RQMe3TgWdGCN3g248mFVj1K5Yg4dsoNlBLzskRSSW3XjQJmHO6/FTkfwYvAGaxK
49HOMnwCEp/uffd6uD8mDIkLieUQ2TfF5p8H8psvjx6pG3yokL21WuKz31HDNv7H
em3188rDr1wdpP06zWmWL0NYyokJDJOi0MCObpK7dfHSpsZK8wJCZ6wAqVoZiVIv
XojjR0zysIK4/pXesx0+oob//VHHn8QmpcNQdS4Q+j1GJbdfLIGSUocoPgcz9Ugd
jS9V8Te6TibJAG776Vf4fqH9CV8uH28PtqMbezlcLcU++gQLEqOkumjGfYjidj3C
RBOLC3BSExEpU33GrbHdcQkN9TQQNt1q/18qCdFL86WUTmvMinbBrvjUZYM6w6SY
bdKbMRUxZ7Vbi6bXAYe+c8a/Fh2oazY+1kt1CeonTmapRbzHXVqORdZ31Pc/Perp
QG+JKFQ4c2z/VvjyXyPIzRElBy+KVUjvtcHofMUJwizYiQcEKQgFUGgUvGGlv2FE
PjlHk6RwgjYVuJ/qLGh14GaoUENDqANT4+LnHRpiQpJ5aLYqumAsxCdncFtzIDow
PZlrQhnFuVdjHQpvhrdrkyZl8n3dvnQ5hAIOBX5c15BdPRvmBeUe533ao1cX8RCe
i59/1xHMJ7l+CoKUIgQixMjDgP5ONf5S32sRITDNeXbY6jkyYBXsXLQs3viiZSSm
OtvyWrAfBwuftNkeqlNJ/vRCipJ34a4xg+NI/7wyEcweT7Po2irOlm34RddBdDrq
Ul4PwD0DNYYZy4BkapCf9gq4lugM5FMVM5GyLVUuQy6KoI9y1q+uPBd7T5QhGd7k
4X0VnGJ2EWXgDtTIgJ8It49bleTBnHxY+sCxcDPYS2KID7sfPo/DLG/soG1Q2dJ8
owONHXBwIHW92cZnIpT67hc5nzb6Znjy+Yk8CI0auAIb3kC2mfUvNBs9jQPLfPzL
4PN/6v/nXGRpFSXo2/sv1dXMHsQPmZxwAYGIEYOWx1hkojBlBrQc3ILqEssgMpGO
8C5d+6RbD49geMepy5smFMeB/OYbV0qqeIqAaM7v0BwEbH9NobsPWjAhYGatwQ3s
tsOKP6Nz+2MM7GHTcbS4skButbErsazEl9AzPsARpunbIflNUUEi0kLsxMwlrNL2
eJYpBbQywDCH8Bvj49PSaCpH9/07X666Opy9hVCYeAfAzhHR+hwOv2lKdp6Y4ijk
/C1xW2pDXuQdJtnVcYEruVKdUG0R8SkpsQ1NTtFRUnEUwAwMbLvsNM/axFvbR3cJ
AwZ8VyMvrvbr1qapWUvKEzFm3W1mcUDP16dxMmTpNBtnnLibQqAhtzuI8AIFV9Im
JecWGzYBs7+xfaLfeOnx50+dSTNiN3XD84EbcBQkQTWFLQDQAqccB8Aa3CSxVRve
ls//r9bO1nW0TaksWAsgV/UWzfNMuAHCyOzAW7wBrM9Up/Cv19BqyVYe6o/oN1rd
vIeVhkRXOtA7rEIVTPC3y4/ub0yonc7QmS5bI/otL8b0G2nU/WLheKHY9ShNIwgI
7uuuYJRgzZak8VNQsn2+4vuU3ds7Vwc8RgMikYUCdyLcK29/JsapSrNI2gybOVaz
DgmMtjNMnvled3RQNp/A6587hAxrzHksClkNWAaBmbu80Usg2I9cSp/muyITn7SM
jUd1SlL7XzF3Q2rQwowK3gM+gXdEm6mAgYFjbKN4dEHZ3C9KtXc69LP0r+VPTV9F
yOGxXr/NNxWe94WoQWP+oywUb5jZL4d1MhnvI2+bAB77PydfDSRb+wCOnmoJTT6R
o/u0HGDTEzJuUJBv5Sx9HfYfKaV1BzZ86A3oy7xmn/z1Bnr0fXV3t2NyvjSWp5xb
CW1tofrqhD7DLRP/TxOvtFnf2ZHHfzV2Jup4wkinI7Nanf+rdheGfUjFAq/t848X
y9enSkklTWu6LelQQhHO0WO9NFp8ZYai00UoS6NiRDWUCGlg/CSaM67yEuEJhzNZ
15rpLFCnr+KjEVx06LLOADcf9jf9LEWyJijdCZaOhU0bftwBYAbUkl6NQGqAtJz5
OmXCAS1VBl6QT8oScu1oLQk8HEr97QCw/GI1UE1l4ENHQ4KAysSoM4F7xTQpYdbE
fhYDZ0W66SzpZGh2Rg+sThGS2W0+ZaAWPrKHeNKSR7L2XuiVYNldM0okJpg1wyCW
hp7WH60buYFrukbF/BxQe2W214RX5IgGyrGVkhRt4Eg/3wmSTm3DxR+h0Sw+Qm2V
tXfaAQnvdzaHNN4mi0LiFrCkIjZzQCnBRL4JubnaOnxHJv/lG+l5IRrG9mEsTtos
Wc8EfDczTVvGeqgzBRJHg6B2svQhjAwcNmMD/DHGhFsN6xwtc0SSEmwy6Vptc+TC
KKvFUyJiJCSTiVTyfVTL6SZlHnC7stnx9HdCGHiPjoPfPtznRBoVbquNG4SoGANB
V0VF+LSx4om7bwRLv2T5HUBvGXYo9Nkvb95BcSM2RKmvR92GoN+Sy0VGSXdOt0zb
25mmg7hvvlgxeQWA/7VgjzgoINiTnZ0Pt3s1JE3WbF94MQrZM0De91RPcm7i8tBR
DvBMcmQgRxozHPHbDUTSSqUh8YuoFvRVPwwPkWsAZxdZBBF/NZDzyIFAxO0SR9ma
s27yPL2dtWxOtBFjUuPmURsvprrkAiUm6crKOcWjxWNsfjsJTsDoa24PqLHVfOW4
PCrTzoyW63DF4wZ6Wgy0dASqzrhKUGRL27cqp+XHZAtn1UI1rmhCRpopF1e3bvz2
u1IEjLhQR+IMiSvgkuXWQRznR3fMlnOSBM1egRDQuhQByody0kiPRKmxepDOb8Hq
GBXQCRLUPitgkQ6xwqz8nWCfjsEdADf3lNMAGnC+iii1O54PWOHsmR7LvQjw23CF
Ag5TQyV1tYeLNlsQOqIf+FK3V7sG7ktl50U6EiOz+RiYS5F18WZEGH8Um8NvZpv/
h0yLgOrLoQe3mAB/xxeSz39QWh6rGck626Q9I+5Fir3vcTsOiaBb0S5M4riMdjgs
igSO+d59MqfVb1onLW1cyBd+NeCCZ3eOZmZ67NUSSqs8kWlpk/nQaGQpYEBvc6Su
yKomS6i1usGXmEqOQYDAYXYc3fE1+MZjiLCt5kDg3sSBKWJ1CSop/SMZlV7Va0Cp
vUBvDL6cH844tyCo9Afa+MWGkFiGA1/ZbyST9r2EtN8UMiuk1wpshvMVLlswFVoD
X9qSkRrd8MBnhD4aScg0+yNSeojBj02EOey7aRfG6JbYfXKGAVDn+C9d0CE7qrr/
p0705aqo7A2HLPcJ06T1zIzEu86Yf1qflLjKxf4A5H98jnxU9wGhi/KRDJxEC0Bn
XX6dPhKNobs7p8krYHcqatnZVWSqMDwFwbt6Mvn8Yr6JZDKH1q25KL7diasH23eV
i3aANTwx9IWHjzl9tj39K5b+RNGu+9k/0yCmobjrGnUDyamyYS8zt3mpjEVN8Fur
TAjK+Etwlaexl5NElYJwYt2Owp2l3UlD/Fu4CCfUuBd7uKgEazWsclRfJ+MpAY1/
EKqB7fTyHAR3hggPxw4WiPHVeVp12WxuN/46ozNS8nBenmwn35PJHNBW4VsawBxN
MjTOl4D8h8RAmQkZ1NgMiVF18aOtwBZc2nRpDC7Vj3242Ls3GnCam4WrKiArC7e+
VKMjBBsg3S4PFOxurDTozJUt2mW32wthkeAzAvBWkZhmxwkVUZuHJk/P60jz832c
/MPCStnBdwv/ZiboXa9/LTxm0AHK4ctX5pS2+lvFb4PW1KHxgNVwWZRmTzGhCkCs
YXM3IN1jj+tmcAHEQHAa9dDWCCnZsAVAymfP5vF2xVjGJOj7+NlXqkatvNolFf2M
9Okel/BHlWxWxE15y7cwyUAqJbIcQ/r/U7HK3IFFfwmtoUyIgXAOa5bgP80eNDHb
T8ki9amHQakUhP5UMdAU7CBNjdYoHxIpM/Umsjn91P7M81c0Sz8I16iGjmeb1N0v
Rf+GaJtqxoIwdsdExgPvW1Rw+Tj7xf8XuPu4kfbR6xEfgkS5pq4EDP0wX6crOwEZ
xk7Jf9Kqag5ls8F4o4s4BCwycCD0+FeD/3zivPE4KrOWT00rN+Y9vRpgkPxjpmpI
r0rLeJLWgnLdGxOPawJKFtwmgl9DJWmy42kR6vEiP4Nu/ZLrWEgC8eLiz+jECMd5
qAX7JsVeO2ard4Q3uUnveOH3do8KkGxAS8wYEMIOcvvxMXTCr59aB3n1AVOrjwHP
GFobNkkCwRzD7faNtsakTZayCdYaNW3CSb3Tw4KTV0pk6kbqwX4NAfhSTrCcsAXV
omeXDaZktvy/AmJB77pSPc3IO3AqL8c6CjnPFMc9jae5rCz99GPw0WVd9z6ujI3u
lGW4lQEhs7V7NWlF9gGWNp8sa51Fxsl8XmLP4fhe2HH+0R6DMtCeS/2yhltc4OfA
HXBy7521FdG4bnlFXpPzRHXC9ZoYGtWKPwA1iR/Xg1k81HjazSAI70KewETuF5aK
2/Coywh9y/WCWftbIcTtjF2IcilRtLeDbLYXeRZprPHynlU0juJWrSHi8Cd+71Pf
pmfcOdrrQoNBGJQc3qM+naWrjbPAWF6p4zCxZldGhAmVZzvm1u8QFIOrleMPY4SQ
mHuBrTMmWeUqYPyeBpioaVyv4iXjXL3VUzMCi6gOrxpAG9Z1Crx/Sh2UOb1Mtpfx
Yb1m980vfPxDvLsRVMH1Vqz73bN5xcO7Izn9W+lcmsLuBKKLeTrEfMe7L2gm/7R0
uAq8Aws0FvBhHtJiTA18O4+MYWv2f3nYlwDsdYtvBJ+ztt0lgJvREXRrVhI+ZflW
DfWxQ9/CExuZiEuKS3jY0O8nPiZ3VgWzeDxe0LiO/Qr007GrD4wRkuO6WYgE+5Hd
4yHGKmwNOdZUCUlPRfZOR001CYcCyghpGDvL5E6BUs7jk7p1xShkoHo/4hAgIreF
N8Z4BiYA+eXlk0RjXPrvQZmEPlYz7nH8oDyMbmbWrJi5akXr4tSOMiYovYRnlxTE
whcnbqzwS6Oum+2vtQdF5FjY7l0K9E7tm4l4P7bg6E0CK+V/H/wJnR3y3uMGOcYR
uGmRZYchg9OA8XEJITz0WneWJEWs9PtQua5OjGvxIkrf+Sy1tlvBMPNBOqM/T8v4
RpQjVi9SFoBEGsITixp+uAemmPTvxu6A0CHc81LQAZ4TqE5a1lLlbAEpMOoMjKOB
hnFgzQrKIjtZ0ErJzUoBaiKCUP+ye/2lkhTm4OSAx212hhOjFbdl37vwF8d6X++G
/TxjiD7nJCTEDLaLEC/ByNUiweOtaNBNrxU543Oo6MBL+oeL4oS445wEP1n/zjfB
9+09xqBVf/iV2rJwZGRn/t/uf1zO8NfJsI4DFV4Oh/LN4j19TxiG8ll/LXe9ivso
YGeqaDQ4pk2SeBS2hewFQ5+IgYV8w/LbPYWGqGHfQjh1w2dQJyXg15+toHAGNMIH
7ubG2uSw5XDdLUeezDA731zbMXjbD4EwWYIS9ngg5XCg3vAqxpZFV2KYvjd7hYbE
n0jAvMHnwNpWeA7bSPRMKMna/o9cPH2lJKigHASfFXcdVfCmTeKanZI+pXdhtRrz
CBn1bbPRrsE5xK4oF24+g2Su2lpdlrpIhOmd9LNO3Yc9cRC/6WzILS+YkRp7r7D6
uUWqJHs0LEbGzyiDr5CohCgxT48ssWoYOUefRI0M0mkcYUP1nLd5FwbsPNKgJNYC
suXYjkf7ajOgWKfQPyMLKpOkTLu46PWSgeRuq5rNJksPf+1JUs6VBnAN45347ZlT
p/LHlGiALL8iRaMVzoCAL/UY0/Fjl5fDw9W4FLQa6l7RPmD/WQ+cxy41wpQ6j9Cp
LqwnLzXAqEM+TuTDJVmrq5kRjPQvmgxPTtrc/WYQwzJIGxkoFuaxcwb3NYEkXfAs
Jh2vgTgZDa3mT9DpXSKAuv9FdW9UA7vxDmMrzeedANyM6xzTBQkHeugwp4acKK6m
lGmWYIDEli6HcQ5iIg7MhDvu6YLOMaOzSRYs5/wEehpc/Ajrh/8VGyfgEAZEA3ht
fS+hU320MfeyQHWazkhgo7825LTy7SHFfAhI7B/o6sXKqOWsf0riQzHO+yhSnJrK
I1bPEswwAEhAYlKxlMAqdYEc1zguoi1m+lcqzce5O1qLfDmIdbCZwiW+k5UZc/Pv
6PlmA0CsQVHzyXf8TUCOn1BjxoJvc1PJidwWQx92fgaUTzwmw6acfDv3HEGVrgZ6
pBmA8fL6b8/QrpVSEnhE5c4Mks8KIleV/ey+787AK2ZgxqTYj+ON6ddBHa7Z9eRi
+YtbnQnUXuAT6Ruj0Rm9V0/vS41kzJmmNLo9IJltWS8/jVhM3x0pX+hZmiZd+sw7
kqfXBcDH+f/tsvt+V+pMZIplr0ABFNN+nzdh+KF3kAmJHmcTXOGlReDqD5fDeYaD
T+J6io4f63rt0Zwn4UaDmwL38SQ2N3xIoY9xzH6913OFtO9/OYFF76PbOR2ffNZI
d5b9lMWana/ax+l8Aa15q7fpigaO2IKeHSsYHqj+rfOw1Y4AvYfAhVDMBPETBot/
Gza9RHcSZKSB3QNNaXwJKsjtInmer/rXVhDVCZiiR7/AIRqp1mVaGlWtV+zTH8f5
XC5RO+zYkXPVj60c2j2d06IeP/cLdL46T6KzIolMEbxdHw/c64LasieD8AGjN/mq
9FLciUGtlvG86XJEGXVVW1mieJHg5WNVO65SupmThdzd8ENlP2w8XC5xyFiKc8/6
Pcvf9/NbKzLd7iIk1k79rO8HIJd2+GBwzEUSu/ikrbV/aVb6oqSzsu7XeECE0/FA
CxDiNvkt3HLp8bIrjVNSCUEQ6Y8x7m70470nSZWczYZMp2aIUSnylK7nVrINIcWM
3X/eaBibX5ENKghmysydvVmLy5F5Sjtphmawck+xA7Z4qYe1Ul1n8A/4HfkUljvf
MVIb/X/TOGfAf4IRHECQf1b1GH8PZaZbQyPxwyBMQNP4NwcHpU7BqanuwrpmpXU9
jTRhMc64DOWE4UyyLyGbP8pj2YF3cXtxniO1zQo2U4JLI8pKaszCpEYXcw79SOv0
rahpZEkp2wJEsc+2We/tEskYaUxDV+ufqDyaHsTrrDI2OhXuRT0P2FKXsQfqhFDW
4L3jct0yMY80y7NwK9erkhSmtBXI+Esib3zlo0Oip0GV/o0/TYbTy4HngkTWd2GJ
x6w2v1Eat3WzH39OmMMz+A5luiTF+QkS1TmMDHkWqKOBT+OFMqtjdMo0DuR5qAJH
iqONb29T5x0tCDfQ588Z6rC+/igIBoWkvi4iMYkie09ugweCnNDDuz6flR/N2uZ/
XM0TPPoTOfclMEOb4CE3E2f9SZsatwR46wWMkNoe+rKcauWgAFc92kef5T7eFRcn
CjCl/OfbNArc3PNo0fNCsLtqddh9dgs+CjIJatzS6w7kD2266V8scnmq4Jd1f1nL
VAOu3z7uRNH2JnjTT8VuUAxDIv5Xbo6JJTRcRFc40uEstCeD84aEB1lNz2+anGau
Atpb992bzA0pJBAP3exoo53zrW44Mpm+leWkPHt7kIezVaDf2Qa7gtiakakO06fH
WTntl5oJK5I2RUxA6hxU4wQMkT22RTKW+o6kVL5VL4ByWTCNRESgnh0JgtCKB4V5
rjBuPok164oSf6CbIQJNQWvMRaK+b+S8c3Ni+oRmvtNwfW5sdno0UjVM/sqfXAzm
ACGhuG0soILwnpyFWcbjZnX7P7sJJQmqbL9YckCyPDtFaqYJTDFoY88KKqgKO+Qk
cFLeP3U9pRkaIMZ5KjkKbAoSMD3k3/kukPT0L7MGMzUQAfZjNNUUcZQysQozk/St
nfZXi2IDUBXjL5fEgVK8AfQWKWUi0JGar9DBdohxq8+UuFL8LCR3tDOxuBKozerV
yKpkXGMo5JvCFkgHaVpZW6iilQjg6MkrzmJjouLHQFuNVCAV4XK68jHc8ft7SWEH
zVZB90Pwq5ajQpZB7d2Hao0vr2yjk6ohQ6p/PXHmDNJbC52uoa6t9xYLVj/lNvzm
6AbCqTHhJ/euEdd4RID+wC6IkrIGRXyB4aBzPqNf21Q7eHJM4nmIwqjDoE/SM0V2
71L+QwyNPFNMkcnIpxThZK7vZwlI6I4HY++aO4rz+g5asf7yEe6vRrO4P+7R1NcS
2iu92mSU6fqFL0ZyNLEmbXD4btRhna+3TkNaua+aofgZ3jytFmABOBXAkv17XAxY
UM8kqFb+eeU3j1zclfeuCB87aps1JURz2qJSeKNTZJSC+42Qmz6dUBGfWPZLznXm
t9xkbDYnp5ZVatGksvRIRZr9SZKvm5RS5tIPcheuNBn7NqDkqM0qQDNATelTpvYV
AYTSj9ObLQ3Mcez5h47fAUtFw8n6T4dyI0ETw5OvZdJE0NIhdLfn+DK20C2KzbSj
h+dSq2edIkeZuiu7WObX8HTf6fqpsF6GTfLn3tCxgXp6rJCNzmdLK1OwO8K0qypr
3pStrzyEVt/lldqoAYcAV4oGlaXmACvatItnouFV0Wm/G4YBkr3v/PK/bF5AM3mV
yJ9DZQcpMT7V6/eNJJiUpZQN+z+lS3NWWbvlc8svFFneYzRDAWyygtrr2dCyns0g
f4rwkHMQITQydiEK3+9rJ+9oBRmZ+Y5LZ0qdtKHRqQ6jaQNaHcXlLCON+DNHOpvP
fp2UdYDruBh6iRLAKfGTZmqtJKfMUmLeBZ3lGa7gg8YKbGlTx3T0otsg8oVtM7Ku
8S637WbfjFDF0Hu2zSPsYe0mh5spKNMa/XPe+0jv7o/i+SNRYgVTB3yjAehZYcli
Ka1iNJv1djobLZ1F9KMscm5XXbEOds4iqLzwqIKgf5rWjPmZ3e6xq0vOp6Ol9Zdn
YOxeQAB9StUxbDFM2ozkQsq5SKRx8FWWOoB7Pwr518eSmxaXL1R+Uim9KystrWqn
ywr3TqLzwurSnHAZj60pQeNxnplRACcEJIHPjAHOZ8QfoI2ilGMYn1YA2T4aCI7n
lAa01NPmzNtXVLkbrsTg+0QPirX3EXUEWIyEY0Fka/Y7wMtzl47e0nv0PJHWutZw
DuB2yx7M3Hy1GRuw44i7dbzjEQzK26cCKxNKETYOVZpb2Y6iocGB2ziB5owx6jOG
XvgAB5a6JGFC/0kI80QXR8zZQ+Iy7oSLdszQXCVdrkkZiMfp4YXtLHAjF7cCvbU8
7aelUuDDq4AlheOE/S6ju+41yee2rE2PDeoKXQ7BBNhPcvN3lebdi/o9clEz/LWc
Pn/vyevmmyQzkwQqM/lnxhx+nN/2hVTx5cGqmDHc6B//o5eY/cUkWfWgFcUkZJR2
jo05FP6SiUmf026cYBcij0Gg6KfVyMaiaAGXl/wte/DBMb7qedkxffO7P9jbpbf8
eMDEMu17dUzPOGcOznnCmK71ii3ysrxtFvssROC0OgjMcYNe8gWjVTZqQNKidcNx
BjSfFU548xYRz44Qs/hHJh724J+NAmWUWeEsuN4w8reTjgYP5zmKs8CnqVv6mvDr
qyV8iJCpq027sDj96gP70maZglxG6P8A8w5PPNcr2dvAV/8pBsxp1bVrBcJOECY7
MyBdmqMpwRLwEiXCwKFPlkyQo05Oz952Pc0mr+kA2i7WA7liou6+p1xtsCwJABvP
5L56UCTXFzVtDIz8dI/lvCgvgrBX1DnlisyTC5pky7LxuYKqCNEnvpKk87mKbyAT
KK0iuYu3Yb5R4x3qarqhVfDoyjYB6VnMDVZCvUvJhrQ2CcHJLrahH8Su63VloqXz
O3GtirpR07v36KvCAsaGuyjihGJyiSmb6TlD3PxQmieCDQvh8q9xiflHaTygITDi
Kf++08UlxLYnk9Q8s1Ze8RHcW6jcyONQk6SDT5cI5Bgsd1FJVcwYro+7NSw6KZMx
L1rjiSPCNupSdrKHNn6HShSFioSe/z/7adr8gXVwhL8NbS9ozsVL4/RstYTYe5jk
OcboTLUenXN5n8QSb0kKnAQaBLKxhj51evLIj+9dFJTlgWnsk7AibIZOMPGB8k1J
yi+JVn6nTIN08ifqfUVPNnhmmP6i553mllwBnpOGluNF1UFHts5v3CRYc8JeRS7f
kcXicHEwmToH+2VZ57cTzmjScIHBlYB/bC08YPu9Zyzg4g6JO+M4Q7LqRj1OUNHW
gjWswXJRlmcMvjLYF+6O6zL9e23D/+h60BcvrfjADO1tg6hu2FG4g1o+eJB60QIA
tqsj4053tzQxV9vowSZOxpLAIYSX4gGtJmIoqpIm9cE7vUY2XQ3pfRS/yTN/TsYj
YzkXF7c+UeJyvxqUkAULHECa6ju9pYuqvEX87P3WHDXwztunUX5qq8uNnJYOSnvG
xwzzpGLQejass7rOuNLm/N39qP1g95tLZBw899Xz+4LKaUaHw5gbJBiKHgglZWA9
Zx633RuN89emuEr1cS7SA0/557sXDjEjzmGVvIstn8/EQQWy50SvcssVpBkNmknK
FOH6kOjhmcYDGOmcJYHVm/G2yQhTWEuFLcLeFLm1DP0BmMG4P7YINk5fG6E+du7A
Rw5X1QzU2xX2j+KwTznUdsRSw457HLvkbWMczFuJOSJzOlVVCqk2M4wvhAm+C8+0
/ci9FmZSI8FnoqISAJYFo9aXxSreqypTeJrecX6q2a8Tq9lWS1zu4GZklUiEybx5
vGlO8nB6riK66B8agGRakUHC2jSkaGgWNvEoLh3RsA5SrS/sJWCgzEu0vzg9R8hx
Wna4SNhMfO60aTnGRM4Joy5rjgh2Bn9ADkXbxXpZSbF7XyqmYDnOnJLu8k9nxya7
/osdtBk0ngkC8b/gTt9uF40sCJ53YjIsAdLSlohnauxsRWFjRBbhTLMc1M8eXa09
C/aj3lEmgb3cKrx0b2yK+A0fJPUF3AeF+R1WeTDcZPJXoaX1yfzHIvGQmjI30Muq
kfqIQRZEbgJJkUySDc1jy5rJU7ojQyq5ZyLZ0bXlQ2AUmoW4HkaThAERIT0b36s2
s3xyPn2+AlmUzVD9+6jWEaBcLzG+2kalEgqKlnrGawej18E/5MP5O4efkWEATe1a
KY2ei+r73lqnN9RwoO4MYnNOT610ZwVil9p+gEa6TXnCp86uU3jr+JkEKxetqOST
lDOw9ZqfoC0Ia6zHvg11iGhsl+EvNh5o0lj6+Gjre6ySKs7KN+eXDuN+vXiUBNt7
fWOWtLOFolRgjMXC0eNAy9zjy34tH4pk9Vtn66EJiObqRhnenEUbCCfAEWHZPdm4
ZIZ0FvKU8aAYNSoLuJPBlzR9ugH2YQg0VLNBl69hYrt3SQdKF45ymNJtpZbW/OLR
LX/5IVTfyf7kY9ErTW/ZZXtOzRMOymvhg8UJpnot1MJm8FiUgc95MwTy+DvKsw3P
Lz9EvUquk+NBMXgL822UTcS2+ZNqHn/LLEN1/H3RQ/EwbZm3+JWyS3LZRo2G43Wk
HuYiWJwfBaILzjy4jK7VkE70t6Ulx4wONnpEKqRJB5o6k5s9oTPe6PJ4meQHKzNT
VRuBk7OcB4s/En+KSfpRHb2E/fK/g66byB+K9k3X2S4+pN3JmaWQWnxRIGX1WQTM
fKQzoLhyZb1Z+gHp9q3JjNNx9EZJkgaJNEolYMoHsqHvZ1LqRiJXdDN0daz4aGkg
Ey7JiHw2WrTkAA2TWB7+bqTQzadlzOQ+BBwpqtBqqsvDCsyUVyo4/uXCC4EN8l//
4CqGPBAK67I2w9I3ZPbzpa3EVeLdgoXxu9NO5OMp5mJi94Wk6qE8O3AuKn+rdjMa
xyL4yj3KYmG1ImtnyWdY0K7k+oVrT6fu2zagaalqSWA29lDTT1dkRDL9jNuTo5E1
vg/qb/29Y32qw1AM+ZdGs+IdIfSn1pyb+wWBjmWxt1wLtstd6Vubxf5fFGH5oEGJ
QwB305YQKwQi0+AJlYnaH8w7T9QdzJJKIwoODuf+67MJq5MpFKGIzdkQgAPUMZHP
Z5Gnm0SBxWNy8OUzFVCzKhfuqQpBgOf4d1R2ilYRm7GQH39ukSCnoL8KOWN3s6bV
6v44RJCIpx1DdRCb5XNFwMITmnTKgASw2qP8drO7DnN+qUJAJuXhfhGkljhjiIE3
gfGzNKPfpUpWoicszhM+hsh2jP+eP0n9PWrA/Yb3aJMT6UmTkAJ40uNgpoyhWioq
eDtzjOIIMWtgmticvhQigZ9WO9fZ0D9+/0Q4t6p1lUFe0cx2PQo5yTB4GBYGbvWl
VCZNyR3nYO59cZjiUGR4lQSZfUDJRVmjdDsFM/RwQd606uZDNbuM1QXvxvRmw6Eh
aah9kdyhSVvLXjfjhwWyAzfKxCs9/4tDCtGat8HXZnZhAF2DiJjGJLSqcWFAXEqS
AtBuz2YtaUmxea89Z+y9D8PPr/Z2V/Gbezp7TzO4oZu8Cro2fz/kBoOqkeR4m+4P
owWElx+Zp+zBpPXI3F9Ylhbm9DN6eBoW68WdM4EhkBm1H0xw1ARqvFIC3TkslPyL
rug+8pNDnLldkzNqOM9V40ntDIHHj39CNHKxXSiMStaaeOyvJIaLTWiFXVgtc4yo
UhnmFSHvhJ6adsjUzJ+bSYUSV/8b2vDqkNiDcd0C/ohO0npbjbrQ2jkEP1/ZcdKh
LUp25Rp3Cmq/CHM9ONWNFm6m+xGn5cSL9aZ4EB2W3xWTJi5FLCKlySRAxfyr1DKE
nFVX0rwi6Uu8UbLCxY8IhtLkwimpEsGmZDL+jSU5T/3Qgtuq3foROtgW0kdmxIqh
6lrQs+ermyDjV7IVti6VTgQmlUeHX4F7BwBhCoBnj32lZ1807Mkxgb0cvklVzERY
i0CJUlTjqs2roT6fOkInfbrJ+wOh+lGmSL61cioY4hpB+KzYQ56+Op4eXbiCM65e
bSTKgxIXksRjBHZF1H2lPzlSUkQyMzjY8/fNlm7rvs19xMHSaZsEeyZL1g2qjiOd
4vraqDASSQ7CzojvQlbt22nCxmoJyqbBFuk8J/T2iEEiUpsVOG4/sx+SHujRw1pp
374Aw8ov35Dqp3kJAOvwtvHN0VdksVJMRRpDEQ7zoD4vQqpfWwHLkysg5WLPMznW
WjlzMEebnLbk39faz/4ori+IIAh+5RAvtY0qg8iaTF2ZTCrb75/i9GSuxbzz/XBL
0rnmBAkWAlecG+aKBu0yQNaNJUG1ofc8OfwpsbtWJm29jD7B1W2zGeH8YFI7ywaK
qFZUARA99H5nFwyohFNPA9iKxBHxKBMqUyCOqMXxDmzF0y3Z0cMkrzEzy0OxlxBl
JotOXATxxyXlWhJxV6qQJLyM70/xxM7Pyy5OrpcqjvWhYLCY+ak2BV6iI8uW1Mgi
tJJ56tVXTSNu1p8SboI2byn73IHStyDLqV5GKE6R4nhmF3YC0sj25nMWveBpBatN
xdjZOcP68mJ//uqeucvwfchCiBpVaROeb14ajeWuc1kH3cqv6/L2KJE7XEc2Yxbj
kdnt6Wg431KX10V4VDMd9WBDRc61BHhvw/0U+06DurVk7Az24WPq10C0ivRJhFRq
4xdsHddv0HQda7+N0ph8+u919Qw0TIcJixzFX8Q7Z4ZFr/q2XXYcy8XWgU12ocz4
9ZgYtnnN6KtPBT/SoqDSv8e3zYIftbzgrhXVJI54x5nc0VHwWq4ozYUP6vJ+aOpw
nRYEu93r35SyZ6YN62RfvrUqEdH3JJ7dbJ091NKVs2EL/YpWc5xbTJmrLgstDjq5
P7OjrRYnEIpQnCvNI+7sdKucM6AEdyj10nHPGHr3hEp/dvMZPJh/Jw5PvD11qHJ7
7E+r/GqdrHkLGpjs6peFm9AgX6sI9v41W/8hcZ65UnbQ2MMd8NhEO87j/QP/X9AY
ww3Q/2RGyHG0ubZKtfzucynWOJdFiF7abTHVbFS6MfmDqk59vmtChmmy/Mt3DXx5
/SORi5KKhgR7T35/y1uQ48tonq6JBYDWgGWbhFzRqi2J+gE5hTBHYQQfgrL+8nEX
SEZ5H5Mb7s//UYMKsLxRkwPhO53lVY4mNGMtzyVRjFQL9o9hXRRRBwktfkVlhBpN
ROR3S1zr+zMX9tB3vpJvUog1orAFJeDr1qAiJGo7SFQlLo5RKFXiySj7k8wRUJR8
/2fYAnAaLACgsunS8qsBufA2qeJvd8Li9A0uMtw1GiWnJsBx+lk/J60thZQXCcWM
zfLG9TRMiCsEfP74WlIfEBwC/C3vudz8roAfjMj0q1kaTFyIFRkUITjkSV3q9Ix2
n7bwavDdlQlVCaBCAeCtHV0hY64726yEYDTdcggVCsZhC/8+D7A/ZwsbDMtn8V4d
tSoupx6WQMUt8dpWyihBj6EZswC60+y0SL9e2cpUdP9xw1mTL7oT6cvTcRHa2yu5
egPUAlWZ9WKO8pRYHZA1GSTDkuLXNp3iVfSxXINSLV4AQaaguax7esVvJToWSmlC
jIxkkC52wT+twV/LwFN+FAsI2cs73L8O3zpVQVqRjo4tqT4llElzYKtqcpH7iKgc
1j2lFJ4umU7MigRlpRR5V9ZiOMOPtiMo4z2wxBKY9pHqWAbHzaD4nfPU6Snr1DJ7
bavK/rFKk42Mzpm9sooH77a5BFsD8T+7r5AT/tTes0rr8iBDIN+lG+x2/yIZRrJK
mXRTl4rD3FYCCKUipdRQboFkZ5uincFFV/T+L8/+zTF4SjTiO/P06coLudmGbJ+A
GyvsXwarXMAOqTDoHMEzupxky6cPQuTtCSFp7yJkNKmllV0j+IrAW2nL9Dm5BPHD
BucAf5DJGXZY8MXY5OV20G2gIjb0blXrfdo3o4A7PO+P5Bp5/gsLyeJZ2DRktBuo
8oyBmrQSMdK47i/e4nd2365nc79snUeEE8XKtsRWXhIkjVVd4ZBcCYAxfqmOgbkL
dy9yA9HcpdYJ31HybtbBckhjrWtKvO80BHXyfdHUaMaCgcmr2lHzPr4utvTwPRwY
Npz7+uezfWOaV2uqG4G0amOUn7e1H+h0PLUigM4QqOeDOR8ciI6I/n3OobxCaXBR
JtvecD9jA+Ya1dGDw+5To7iVvcEQ6h1TGesWupKE1fnlfqUWXiFWFY3ADCDO3dqS
Ue6mpeTejvv9+tmCENaEQ0p1ZWgp4DGphNfPLrpv1lRGeHVunzeXcQWHDOlQpCpJ
Q41Fn1G0CW1U05VOFUIvhQ6wN7TRgRGTluDgUzYziTDbrmqAz4+ZK3a0FXfDRgHp
OREVpg7mXJeRRiGObI/pdcMjHfm39mk9swRMvC7+DVj1J0OAJuemcb96tkicoMps
9P1TFnYpjtz1awIjl9sibUHozaMBk3ZR9qBvoX2rr55fO+N4lsP7+8pnqTTC7LNO
X1vJbqPIC12JWSTStLxXOZPNfO3kSbUK6B57kX+EraGaNGpKVrDPam/4j2byPZCw
z64Rt+xS+tKq6TKr5fT8NzhE4lbqGgnj8SGJs3SZbJaSsmpkf2IlVljcP0WFLVlD
9M/Yuc5vzrFZJBGrSC6JWQVofpbrLnDvxMvjupWLgckErdFdVCPuZcY7gMIE9KV6
5JKoMqG0/54UBvNlktadrCqLKV8IaUFVhe3F9Uk4v1lvMCuN9yWjCDrMhTDaC8pt
Xw0JGBHVjGMbJ4tW9j67zB/A2TnVGBRLSMuGlZvd/4GRqllgDMCQQcpV6sGUGNjc
yTOVj+ElNiLidJT+iEisIXDbHMIHvaE0gghJLItbc51PCUjpgs4mM3aFVa4h5tiF
g7fem1wfbrrg2B6CKX9tUkpc0SVFY5R009tVi9g7af/ll0dOZT1tcBi9Li37pT4d
/y02l/YCHT13n+ZgHJeCzFVVtQ6WWWq3Nlb+V++uV1JRVWu5ZgR2V3Z5DgXIL+oJ
joslJ20M8ePmbGv09dc7EQEOT8t5YRyRSlZzBCOtpygGloxwDGe6REPy92y+ha+I
HIb+J1s1dXj5pE7gt+UG3kQU2C+oOb174MqXvFIusJhnK0Yd4L07tAGYMxXa6TOk
tWoa2YElRUnm9XqfRKnJQqC1KrKfpPC95ppXBzCStWbteMPiN8lKuO+7TnOf880z
wVx270qtczCCmBUiv3MZPeSvkCu2qlsxePMat4wA9IzAILibnDZuJ9TrQoeYjqVs
SAJ6Ywi3RwZs5i/cFYhIbsB0g7IfpiHye+39T2jUfZskWg5RCarmh+5QgxgFUsRk
9jONythLOvsgVhnEU60ibf+m9myZSALq1xNCY+Ico3yjDRc63KeQEJYLnx7jcMUt
Bgtn9nRqvZHbaRDZdNrspCNpnDy3c3GdMs+n5O/MSVuqb79Ks3nXuwamer/1dWd+
qmEt6lQzuyJT9CLNrM01+xQeta+sZuUDOPR7WcDQ+2yoNRQWKQCy+PZjxPD1rRZ7
E0THw9m64Dg/A35bceoSVk5ZE+d02TeGPwO0oeTYxFRG7C89BkGiNf3Nmtpdec9P
foWVSj8aWQOXI/R6BYXzbS2tNdGGQDoEvg7L0y7zkkWNTSVpa3+u0Y52cRYOaOZP
ZQLAU+qYcX9kza/Vs1gFkHo2WoX4glqOFhGBNfe7ow0y/RXTBFSORDjLFh0Pyq/0
PhxxF9xJtNlnt3cvwChnQpm5I6EC7BMbmvpV/giYTUaRRcLbCQz6jOOeF8JMqqzr
/12+KHelUb1XVCRllFHk4x2I2VM+raauprJ4W5AmP3k/L1/a0OxWNFK5OKDPsGOP
A54H4hy6TOkKMGePH7qs7rgtKuiNeWzHMRRF7ErQiTJNLob7ucb++3o+MZLjxAwd
1wqKG7ibksXBb74p29Q6+2R8h1mY73hxq53X7qC+NELSDWagGvaPzWQVt5lr4L9r
fgaOf/zejk2ISwfO4St+4YllJzQsJt8SK3HLU5m93hddzKwdHtibzzU9OFdTM1h4
yYSaZhdO4EkDXWiUCjv7sHXe0dYdsAHjkgwL95wN4cjLyBoaI2DqsIuUAkW9VWmi
JtNjHv2IZqOyRFgcOIANRxxzLJ9dYxDKy8QTbHS4L2xmu/ZNCIiw9d13V3LVKAuM
c0rbCrqtuHWxa99jgBNnXY/JPq7FNhqtV+qhbvtvhUOerXN6aorO/xVp/k4stugP
BDllGlFWX0eZT3+KSoX9kACFafZChAU+8q2yq8wplOXpi3yXPP7/O6d8RdX7qmtC
eyIRFnZYsICXFRdiYpui5kCPED1BLMPtTAoEZ810ifGHhkvKJ8RBwwE59nnsrbWB
tzwnw1t+PKyBXm4ehE0ghIzn+Q+lE2cV8zS9pO4YkRBtHhkhn3aV1wqAppZmdcjj
dIFNwbuc97NXSv4djO2LiAWZYqEf/f+BGIYac5j3YjG3hzpZ0Xvs5I+/7OjHCMR1
CFfHVAfhvr60lzf2dAV9S1rQERHvzFfL6gtWIt7syiBm4lwAkbLoSg+bQ3KMCfUk
aLnsOArMqpRgJdWutxFQSC0VkR9p459DB6kiXC5cWEFkgR7n8wd3uIuFJ3KZrU7R
emX3pV7wxiFVUPcAwQxcUWVZ68CmUBA3xdxZ1k6SOXPUj1KvGbdkhHhg8LaeCmKi
yX+TMErxQxp7aoD6/HUp6ossnqeVkUHwVTA+ZzpnTwJ7SWwQtihu78Xd0W18d9jJ
eXzfHCeZY4sHAB5c6gYjZjnG4k00tsssNuqSqIeh+WIoJhoIQhEUN4vkpEYWaKMo
HWkIr2LLeylxJaHqyijukAytzIrsm3cSvCUTNSVfgrIZrMA30ssbpq4TaSpLQpMr
8/w+so6FYcEFLT4GrbHT8TiQlmmcjpZMJQGvIL4Kj8m3Oilix6EElyYiTSP2dgpv
xVD11Ct4ulKSoS0PlhgMvAKGZlvR1+KfUSEzT/09PcTdC+nJQh3lL11SfC/vi67k
iNSTQCgnH73LZUUuyhXkSMcFIddcdRWtQ4RqFNrAiq8DxkHSETK37dTzyOLzEff/
1YnmAVHbg2ALN4KAOlULL6HljwmEoYPy449i6vdZoJ+xs9MJsQhd+tLE8nPQk93P
AWBLBpxnTmYRWez9VEY/6miUa7JNVQvPQxyADR8bRyFqgtZPm/freX3EQIdWvc9e
IAM8MMZzqQeAgyhaeZyE0vQR3NnUJRdxI64DmstqoYJfUchvtz+KgbLxhj7ouKRx
qjLmGV90/eXu19lM/qYB1TlrwQLhfIXfFSoKjltvYPbqAQ+3+eDG9WjrMVdWo3dq
vEwb1TF3dQMRo/6bs9HUMdKvX6gfi/TTeGMtpKVRck0j0bsfD5WITBP8BkhiO9jK
SPPYy3VKvGkQ/5WiH9qbBRx0nCRU0NJzmRuNeKEwAOjHcjuPLp4zwbRusdS8vz7D
Wn8QKpAFWsd0xeJv3ozc3Q/NMYIpwshruO3MAE3K1XQ6tyhT3ck80BUOfKnj5QQe
BlLGZe7J7XpIgmMzfCa9MmKK4q/0VVYk+Bai1sRjwinL2IlGZHApa5D8wuhN8g3c
k3Lc1AJLCReDbYU3f6EyGifDOsPKp94NsXukHp9nV3sUNVTX+qAB2/Rn65bgz29i
gw1Uq4TBZL/NWeeGzD+fFXo9wuyLY7bclJyLUzs2E7stHigOVPyvcnCdbDpT1U4h
OcQrKE029vm+M2YHLrSg9g==
`protect end_protected