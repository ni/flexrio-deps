`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11328 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMWORzZC7bo0toZS2Zods6Xs
yljw+BvqICQb54hGe2JGpB4Fmds8pTWAT/RNPofvXQohkP/2DFIJtuO5yxgZbLn4
V/G080B/2LBGTq8XpLJ2zq34/QyHqsA/nn+ElpVfNFJL8OkCAkZzMX/KksCh/J3f
UYN8/epD+Mf6S0NvjWhYaxCLRqPFvQAW6fnd/ooG8KtLF7rb5GCdWVLQCVr/EE2p
CjnRDKQ9CX/rWHmEOXlgMUhudLcdxT7KSFUCDAVcUQoUgEqMcWuwTfAgMZNc4Br2
nGIjaOCqXQPe6/W8TzWI3DCoJSuSlUnN/UqkG7uHptYFHaU9ySQ+/IJoW1WtKv85
fBxQatM3ERomiV7kksT1wM8gtqIW0TA7w5otnjmT6mAG6TiTvSVKmrdFAXJOJoN8
BAJFHHXWpMwjAipSRaYv+6NBZJwRK5/h+2P/qBoDtJpRR7mjcWa6PzYlcIbB5Wu6
TEE1Aa2RsKz9YgqNYCYF+ddhgO62EVJAlbvFpodJXJrBONzhF4+NVbDtDzsbaA2u
hQoX3cjJukCIpMDkEr5isQVKLLkYJp+25QZ1m9uzAX/oUoENPJHskdanTb1RawvH
ymk1QuL4UiuPoDml5plWou0XPtIrrrPklzQ5nLzHHzk/TE0UoosdFElJqUjG/s+5
smB2YqG2It9+QOegfqIlFsizNhSovRE09/5Tix2wq/N9rXOCfQevwBs/sJIusGj3
X+il9n8m8cxjUmQCLrch/Twk6x9L9KgKciftlwUP/Mohn2WxvzYEhgHwglQqaT98
OnVJWlCjj4qHOxG2wijO6RcQ14PcIsdxuiHbfqVj3dCI8G6dtaPstdQGcZJlEjoE
YgV75uThqodfx5Hrc04WRg/dAHm8cEL1EZJmMfDlSHNbodjS0SjxFMLDJJL5rNO6
UaBi3t08woKdVdDtt60MIvdcXwBK3PUJ/BHnfjNobO51jLAxAtcEn2PAgZuBm0j/
Cja1Q1sRoKz+2Ob1MaVEMbLDD75AieUJj0oIMmK9g+iOXDsPe5s4BqIbVtLquY+y
zs7oa2sh8MZ3AfG8lfyOlJx5PHrAlGo6tdX4hF5rmZas+Mx1cuy759rmjNWtxUMk
VgksjDbC2IuVuH6m48bz7tfFhCHpvjeX+amD4GoRjSCriDpwIXX4qaOLh74Qa6Aq
hiOgqkjB63uZVAlkrUoUYPYRr1SLI7Y1g7/uNw8Sr0GTEPzVm9nk4MuS358tZmjb
p/TWM9Ah8A6pQPc7ro9jpcMgPcqIdUevTEXLlSeOSpgkHnrkwkIZWUq4sd+C7ltp
mGY/hI17dnFDUH2Gvw057iZsVjWUzIz/7F72Id7UlHlXHrKWpTn5nZevohOzJXrw
WozAcDqYMwwbsZRWGsZqPBKUvaZqd7BwcNlNOaeQgSWX0swn18DrlKGc9KEwBawI
pjS+7P8JtfUNvhIzu/1A9JcvKHzWwf0D7hz9OwbHXq+BQ+ghTAtRfNxmBVXxkQkv
zCvlXHmvsAkptKhtbtgxCULcq8fvWQvuXGDkLn8hQtJ+dTSriLZy6i9v2OuR9jiY
73wIk9T5mQKyj0DhjXHiIZr+l0InaH5S00SttgEHfb5mO4tmOyB2ADDeHIkvmwNI
/dC/b5VAchWr/+Q5tQNVfqcwMubJKCTejILEm27SisV9RiNgm/QxyztuLOoGZAo0
1o3c6/5zsAMGeKBBV8N4SZXgstCiEqB5pKXtVlVJAGhvlnht1vThQxLa9y9pSqeN
yQZmP4Nq3UukEpeWb2bCmkNE69WMfog+6w2/f960domxA/J+ofq244CQVhkk7dQ1
cpIBoP43coJQcK25muVSFRKut6Rw4FlzRw5RCEIjrAdNBpIVhEXGyBdT7JZI1sc2
9NVPTs5oozakHa3GpXT9a+27ADWC97DGeqn1Ck5Z7gR0ajXS/3FW2xlGa9dmUKjP
QfEsuqYbNXGxTaLYTPTMK3aTGrZNjNYojleexpPg+RYgeHQ3YHlkvGSndXy5dStM
QlaOuwptPrEwcRzvu3VTw2OMY1gbZY1jxWpiGt9DfASL/BrHqrlawKvVY6R3p9kR
2IaEiJpfy/MFu2DUGs3wd3/LFXCD5yVXOTjClAjFBrLuJpnr8SbDhzyn6R8Bu0bP
18x/ND3LAGSQbyN/mmtVvj60iJ2iwMDAVQPeQ/IBc1X1YaXmKOyfocZZmajWlZEi
li1w4Ke37/Hj2B3Fd5CTWZp7Daqb4i1UXb082QE+/MCejmmBXWV/P4bpbeT6MoeA
hM/tT7YYG3wfKoXHOuJ16NmALAQrqd0il5wi67wHAVf/NNpp8k/yfpK7lQ4R22Uk
CuuH/AlLMbq1uM9+A/GQHA2caApoFh/WOvYitPnAzyyekCoSPHMvd+cfdSbIDRR2
52K1f8/UaWWHtG9QYUGHikbfFHz2LLfGY4ctT4+/CI80bu75sDC/6sRJawm+69B2
W/HCLTri7Grn4eJXAIZSCUpclb6o4Dh9DSH/4cLVEy8QKiHJzkMTE29Is9ULFl+v
1mmhofhpFVVQQQx8oo5yEcF/2rpZTBMevAoo7IzToXVm6M1QsBJJ8S/UsIfE7Rpg
5jGm3SkorqT1/IdC9k/1ISq0OzZgB3iotPwy7EbeclHhJjrZ64LIOPMMp66T47Gg
sYbtpLQQhaAcShNqpqbj60bdAB7deJe+bdXjUseq7lvJy+gNgvsqLPwtxaufi5q5
BlicVg7qXuUDCLNQAxvPz6Hp3kvCGMAzSNlmBivHkFsjyZZjQkV6sW314n9euI3U
yBRjs5x9zPXP5lPEN3q54onhHoXZ9izOLT7RtvAxpF0+vOioX2LQgxKUrIjICq4A
9k8pFnUj436wS1YwPneMDOBcckNfelXkwBRNupReVaDThqIJwm75Gx2wencXip72
NyruuXNMX4aX91zp3A6C49W/vjT692G3ugA0bJ3nNk6IAM7PHAWASq1bDPyX9xix
+obVt4R9QA2mFhHOJ6yyyDqz7JP1E3xoAOMxRg6OkWCTjdeH/w4Dj2wn6Q5/SSth
yvILE25FFzDh39orf8ARZKD8WGhbK06RU2bMz4RMteJeLnwRuGv/J/a0KCYUJMxu
E0xk2VEb3BpAp7w6osIDC+iSYPlFN85QcJ8Y0y3oGh6LowdN8tUmsEcqVxZ6R2bg
yJAxMvTXjvcep1ma9IVWrbWJ5nf+tOwBy/T/FoDr39JV6W82xrDtqWUM/VvAs1dp
aOFn6f+Uopkh4C4ykK/7CJyMYe49FbqnqtJXd4eENElpGeZWbxd5aW0RsGQYYw9q
3ZePQAz1BbGp8UfViLby9fnoMstrTWGLWzsFeI24EOF5j7K1xMg1VkkyaGDUvNvR
igDDSamUcg7ITY7NKH0Nlmc/Po2blLm+4TP+XE8KyMdXbYOxfep0GFhn6djQyIEu
IJPViYgK/qdqGLuzzQuuNHOyA/mnWibWc3U4rAoJQCaF9aPN2TC9BKJDFeZE+gOW
/CDHPcD4fqjsY6LaJwMpLf4a0A/6JSOx0mh020nnO+5tCizuLxbua2tbm/Qt2qVc
634fRnpGCnvREoba37W3YfTzmKGoxljIvuN17U8BMZKPV1nETDhgrOYz8xkMlEf5
mkUXPvsO1tokdlsIP90lo5yVDp/UYyYA0xYVXTCebEPQE9QhLEToiCGag58Ie1tb
DnwULznXzX4Hz+O4vMt8a/2MKwRlonFvWc8xPumHdWf7J7DdE+8dqYW78lulDND3
kTcb1j7tgOBlRPjJy3mXdbzaPXKZkgkzTYxL+DblyHQi/TGxR1cJcOcXjK0ICIPT
ovP4AT7BHUh44hxoN8y140/fcK2GZnhSegBhGBEVh9vA2bvCY91uXavTCRUlMsGC
FNyU7g12yP1hI6BMtAScz3ufT/RujybkK5bEcfCLjt1kz9TeGKj0LpXqvZpRneBM
mhh1buQjsbo9bFC1kYMV5j+vFTnXy5MSzHOwsj9EJ8dFgf1ZMPJ7mNfbe6Td9ll6
rX9P6UH5ylyeZDD6oGVzlQrTpZbJZ58X2kV/W9FbSFU07khCW4GXurQ63eSUsgFA
gQowKaAXLZH7I1Jcf70tEbHKl3HTMYbXI61tESs8d2159ofGi7jUxsD3HpkWraQ3
B5CpeCQJIMUSBNORLYHHN1m2LpTIkNA3SKIMqv/Nk4p9rZqRUCDnm8+wpULqRlKb
OIBxxIUgqem/ImrS7ro8zFmNbSSrb3/h2nzboL2XIitIKQcjH5KqrFXJ0ys1ndW8
gVCWKcgx5rWLXNCt+S5tdQFkjiW4RjCFT7HSkIon3Zt9IZtXR6FHbjOZXPQnEjd4
SpUSsCMQ3Y/RXxYK6JMu1CO1K+ZUwM4QdyK74/AwMPwlc7wduR01l4+o1lVV9xMY
a/2NhSj7+inPbvdsFHKIJKSjH2paoDwUExZzHpb8MmwNfrURSECQiQ9J8jARqXV4
3rln+Op4NyU+ZxijRKC9ncZN06FGASw3NGlinE3d/CznABnLTvXxfDfTUgAqCPls
zNUWomxw4/lbQabLmUaCO5BW7WTfaZf5h/Wt24Fj6RKya3srEAxeB58nsuHW7vOk
RRCqxNCRscPEaABI58orNy2x2/lbqmf1QiWUcUD0IqgomjloeU9b/0Rp+Qa6c1i2
EcgyGOGKomOBJk28JJnpLN3Nr4ZsQp5Doh9lMULKgAbRmINoTqmBFjB9OQoZdZLB
/SHXAD1SaHA1R8m/e6Qd4AZ5ohxg+kI/nPt0sDCcCQXnpXR8+7s9Y6gC7ozrmXhw
8y2ZO/4A7pzi0MtXbA/cCBQs/5azlfcQYBtzt1AyizRTpPC3OlYxw2stCZD/j7t9
PFtjbkZPkKYE3QBgOtOCsjT0ABQhKYb5kHPSiH3dsPs40x+dDRRYoZoWGs/fMlWb
7+60GC1JeHfLQ/9tPm194BsfDgn5Stt/KFR24VE7d/7RusrrPl7vZWkXtx+Jrqqz
nU/kVpuLMYKKT+qojjdPaemWLEjghjMl6oVmBNrDSinu6BF4vD2jUdkXxjHMyZEX
OpdrhtxOcXS9rKTR2U+2fOYvqW2LcXo2foCBAhWfwlVqCTOwAlxJuBlFa/irZ/5B
COdwCYGbs7uPgbnZ4IzQp9ne+CcSyzhlNyWhecr8c/ThDrJxyGCrS0SK3+C6cc9S
U4JS2RUJUeliPdeNkAK6p5ToPXmYU4+XipU/IHXX9op1dbZmVfYhedoq8+BzaXYn
IxlHE/LLQ/cBlvoWdrz4bRCVN9yHEQqIUpAL5xPMhQEcwNhXTCMnmWAYh7P2Iq8p
j9My31tFEIk27Z7a/t/M4cZnEbI+WYpOymDKtYZ961MafahFejpntSb2DN0jEVKS
E7oXbo+UEodrzJLkNFu5wqvv9q1gVS1jjv2gcUqqVMhljuMLNIYDLQO6DnDPi7R4
SA2xInUsToaecYP3FEtl4EX1DWcgExOa/Ys6KCtdcVD0Ei2/7K7t9GlXEoV8GBE2
+qqs8nEaO7vvRjfQB01hygDV5YsJ12d7UAug2kklMYsJBN3NL4HSrn/C85Y9N0gE
hP0aobnC/pNRCG9VL6WcGVpne8VGNFi7AUBWzhb2IJPzYwtfI2+6KlLNOjEuwTTw
OzrClOuMueMyIFzn7zsFu2gGCgRC+ubiukLxnv/4H9/ZAkCev3vQ4bZF2qb3tYEH
h+OG6AN1cuPAh3IH2xq6C/KpRYgYl8bEpmw05liFe8skQyaY2R36R3DE0DwbbyyL
SXLZMwrgnGIid0zC/DRJRofA9HfkbaKJ/e12Is1oNvzD4tcNBBj3xDJC5jIYr1Cx
BgvwYISlklzadNU2pW31Qs1FXoBvV38mAmoqngx559iucf0d/bl6828hibVRUjw5
ConQfZrkJYdFa48FAQLT3ua08KOqE8hMd/+x98AXxk/+NiZRvK16UNl9lmD9rjbF
laFYQvN26rnQeWI3EZ0PDdGb6NLIevrV+BAVLQkK97QlGiLNTTR5r75GUa47z5z9
t/krQVyaDxFOksoePdPgC/yawkjch7lXoBjwniDncS825kSZS385sEKMOWex0d5H
Ct0ycj2e9boRCLzeRbeuvSMlWDQzu9F/HaQQNd254AS7SiVb2Pi6GTOgCnWPzjM0
C5uG/aezxqa9xi5PS19ayAjMCMEkn67891xKt/rGk4RaiNlDeKzXqc1DnGJGSeQA
icj7uaQr9WIj6vKTwMbNlCFyAu+Pnvd1bypvPpPzLq7RXsSDf6MUBF7w0mROX9Ij
ZVyfJJpS1v5M07H17yrArx0ATtmstC7mnvI5ys+imo2rUHLSOGvvJPa8/zq8cd+X
4mDFedFRLksSy6QXrhom+CyVh62xoP4KmpxQrRdLKz0XYMjh5F5398BfW/dWYcFT
H306hQAf5IfhLpg4Jk8tm40aFEVTphiqCNz0KCByOHwDq3341U8naw9XO6UwgTPE
Br44eT7/4Qy3HZvAnMq7ZuweploBDl/Frt6bTLXL6NkzGdiISspUi9nlv2dCpCt9
aU/ueam77dI/0E9MjUpuk4o1itM3/zANzvpiSe6IHq+IojDy6xmY348yB0eUvCva
xLGpPrWN/17AykTjE2qtRpH0to8/7prklS+Qz8Wkeff/AuUshGeuZ26hX/ISREOb
JaWhLke4zt010gdwn1xAxdlxttFXP4wCKuWkfV7GBUV0Q/TcViQbPbHNzL0Ovw4t
yyIB8h+p5W1/wCa9gcwVJqp4VOmkMptF19aSK8RjXKQCVQ9uIkIkUBzjC8TBZ9x9
ppElnB1tTY/CTtF3K3GF5Fg5M2QywqhWbcr0UdISuE9jzeOkf259BoiGJG6zABpg
9ZzP74YiMobfP0VD+8QTLhptZxpgXzNqFhj6Udr4Xu4abLFXCCnXpnZILKSaLbFb
0DK0V1HGsCtWIH6imZU49b6WWFh56UhUmy568mHUgpdVPZAZrRdni/hCPHhS27md
XNLS8Sw6DXJqNJrobza9NvxeHUSzFLPBUgPFLC6fearO3hncY/aJQB948wlQgEMy
2oHBI0XXlw3Tyb4drM2q17G1brMKvWQWzLMg9jxN5IS0kUwD6sMuMQKWGibRyHA7
zQkZhs2N/hnpKRO7wyZwAOnCzX7mYv6mpGe0yQ6EQVNc/9h1Im2VHA6Y0WZy/oZ7
1lxND3Oj/ed6+gwQewuuTROuf9bxclwndBFR5Gg3BPUQ/jsOA4OU4wyAKAoSCHpX
ddQb4+TBp3Q8BleWhdraNX4a2vtjOulHJ5BHmcQWFS1OvAlQ6nirv947fC7sfuft
Th2JPnd3kzTCv921rcx7G3BqjnAHKoKamoMFk3R776yobEXYBFjxrknNEm0em+y3
+6iWweJ8DHHvXOYj0cuMdw6c7mQYqlkWWIZ8Shh6Z50VuhJ/fkUjF4NGi92nnOSF
/ZvIOEGdGvUlKZhDY40Wdf65oOFSfYFv7BVQM/xVtjYDPiOZmVwgKOYX9X/ylXUv
QtP8e49P+WMY5SIiUeoioyCkAG7ctXyKQjqfRTh1Y5V0bmbTYDreeWQi7B63PYZW
18Df3BvuXPST63RzHna+P/8XDw3hBZlNWqs3sQQ3p/YELgJKw3KasV+E14It/1Py
z6BcoNWE65WykfR9oFGOEnRU4AjnVb4KN3sXGtO1HUeZbEyyXhdAxm6yOzgEdCAi
ZQ7LusvZPn867B+76NLiE7Jt17w3UWCcAcKaVK8fJ0KNsuo+Eg9jLMQzufxOEB8D
JM1oHeTYSZVmjMaA2XkcvkCGTFYBXRzOt3GsaQbInfjG2Pk3+IH7RlL+kzDU31gu
o/p9jQCQoeUx6j6jwhHqGx7Zd0egNB9Ibndqt7yo0acgTfqXk/93XBtjVMS/htw/
00j7zRpsUFCGCvlrxpy+jzgiQRJ5wD3JBjBOa+7C5+abfpPRSWauKIP6hgPy9BUB
IApmJyrdqjRZ3ASMldHcM6byhL0i1osOptOWnzBMD/TuHtzi/qDo90h571ePqvMi
mRVFWsZW6BRzCRD89o0h72LbsXoL2Mdqhh/YnysohHXIUXbb4VpmU/A4yI7wGaYN
mV3RQKZkAsXoPPsaNK7gRxDt65RRykl/Eb9MlOybV7ccjqVVbF9pznDoAupDMqvl
MUpT8Vl9RZEMK+23rmyVsAE0UkZbxrVR7ui3gCcZijE7KGZWpTU3tM09KxWhWBua
WfFPrs0OZK6p4FfBS0/RcqDArr6VMMlQ897PXZK886k+OOtA+cq9WftKhcpLPimy
m35ndUzGY0OX3iw020sBfLugFKPybyPgMwO3Vn0zm8ubm+4vk5wRYsxQgCmpkPsj
Vh+4yRZyvg9JxRVGpytVSZcQPOlbi3oM5ne84Efd+u6yMHcgZxgtPkpTG/YG6Bl8
BAAGwUkS6pZ9XXYit/eSw4OtAvpIG6Np8mJVEOzhmzWoSJcLpWn1/Mb5DuiBlfP6
3aeQhpX2l7pMiY4z7Ia296cvY9OVOdQ4CePGs+U2igQFECgKGqjLhibpBeOnLEsu
X6GRpALm3ve8zk3YDtlagnml+IBGX6MomUMz9IlWoNw33vWuAHDXeu7XKFNcK1oy
aJVgk0iD/AoaeMqaTOr03CD2qrnOxVRkdIBgQbdds33X9vDPizl7oyOL0lACPvKG
gsPi+537G7tEhmPZirC26qqAxj+LNRyZbmi+oruZkUSYag61Z46ZWVjn6GutSI+H
dxf77Uaj/YwEQ9EV+sI9N+4AD6FFjvhisbsOOjpijVoOX60ujNulh//6WkP66JeV
RdvnhYAYz7VjRgLu2OhBgALUiABkLcY//YB/xm+FMKNMsF1Sw6yljeb563mIpdUk
/NZXHSAcg0ozawhpdeLisksVr5H+5EJTH6tj8xzze1euKaX0cIKUXsBSeZS9PKJO
b8OvBC5/0/LUE+AQTzH9YflTXfn4H6ajFCBDZolId7hlI6kXPc4tIxJsPf2EEBk4
bfb3chUxNf0phYJ/5VitNw3eIoj4Xy3AcueiMyT6OQDNjNenyfpgGtBqKdYtyuxi
SjL8jA+n7n5m3q7b5gnYBX2Mtd5mW06sILvqGzXYf1i9Xb01sB4wG3HYZxQTCCZd
nQflRLIJ/JxhZXPTRdS412paNdKr9CzqIs1Rf4ZbJPpaSTeSBvey/tvZOjXDKjXA
uBTkMfYYNU8CRj+u1kzKmB7dAme4VY8hSWShQRD9kJT21BjeMKi8XvJlQCddG0Rx
gcXcV8JocgorTTjpSqVZzuM6MAPC+j/1c2wGYVlq7Vc5+K05jVaNuFXS8liNI/wk
vSO4PYDNmUeP7XxPBRQz5DnuFDNeNa2MC1aiQrTaFGIDqHv16DAYSyfjC53Uk6au
vX+IEJnaB19WWIqMMkrLkRpshQEYGdD+Qw/elNktF3kFxyQAjRTvxAvkjiyceiMS
biHxLhDD1LUn5beXFpQreaq+OrESlbLm4C37B/WFo/HMSQB4Q70OXJrjQzk1Jm+Y
UU16dmFAGYUsDFbTdvIJPYQTkj2xIM3KEwkzPhi2gpkvNQbYVehoNGjDeVMaRsTb
IFhony5D96AiEe5p44RftlKoMuVUYv4YpOKnrQIvlZeSizcgh41DUi8Xoi0Omcfw
+9y8mD6ZmqS6GyK864ET3QGIrpiZYNku0veQlmA29w1D+HJOzks/iYh0mL5wwfqo
q0rPUU938dyJH2MzfvpR+ZWBam6ZX6VtItOepqDjUNSZLDXM9ezX+6JCIfQmu1Ep
xKyt+mgV7J6yVG8gPgT0MKH1pPu5unxPnQZGKnuyBmMOmYNCrk4g1PmtQq1M27cQ
5XnMF33O6Z9EgEsvVcB3pC+jfDC8YVnkiv/S5udXWu9sS7ma738vI3tFC8NEw0PN
oG8/y5hFK+cH2y2erwRpXYQ067P6RKIOlJAjtdfxrNE8Cq2i0HbU+h9s8T4G479p
rCkvWIRp49I2hrGyFeK/hYq/bImgeRl5rRNruB7Nl+WdYH+N70AvPBrBipS+1TVv
unuMlVCF9aZhPwFD4PX92uNsnU6fwpvk/8TubYkrgFculT1yighGjG3+k8Bsf6H6
QIAARCSZfaaWBUlX8FbCt3zXEY42jE6pmBxtMS59wJhZxdhmLRJgO3PP6QBTfVHh
aFRu3r3haXozGESlX2LNIekKPT5QwRidCo6x2ctNIFJQQQOhvbJ2dptu4dFXOTNu
XYJFtrhKAl5J076uPKxTELVLzhiSL63XdnL5yKnd+Vjrliu13bIhz76PKjHTAXH4
qNftjRT/uxTZwZrBNajYiyIjV2H4RYgUh/ZoX0p0AD7pEM6NiBbt2JS3cBieRlO9
PyP+FxYPlD0uzjih/8uOa49dWUXhLAjjvh9yqr9iMrkYornvE6pBU2NSQ+PSExpX
nkg+os07ykNsGmIViv9NktQqkH0qHrZtPUUyWZpwPQYW2Dv+gxsPGNaCJez7Ai9K
WLzdeNcUit1DcVt2FyKFYVcRYFqXidsKHeXA4Svs+HmK2Url2M5Wh52ayawop9Xx
J1CUNrne3G5M9YqMsLvauoVgh/dgFw8Ll7zdIATD4bPTNAsOYXwxofyAe0SP49gP
kHvVfjRFWdCKgrqWohQ/sa4fHqN1t3YViLRFQFtb50hlVrMR48aDKXwGsYILk4VS
NRLcXeFwDAominaSzT5GbnKpX9Gf+BYRd/bAIs+lJJDYF4oPY9tUMDQtkBC6aoAq
srKBMRXPO2CPYfLjWNAmVFsQb1KwmZnS4fPrt926Gv5/OCqI5KnyczdhlCCpF1e/
9BRUtBgJsF6WyFX895SgWB9Nk+vF4NcKJPSYrSnlVCRzBMKk8ExDlVREJ2ShsRbB
AgFGyybyKZNbGjb/V/Wb64rSGxVfVoGcyPb7gHFU/SD0bJ6QwpMNlTjehv6W/QKB
5+H4wLL0HZWuvquNuGgS3tyfyFHJaTq3y/ghRZADF0WIG7yfrsNpX9i7TeyAnQVN
uG8QPlxasW6gzRcEfkr1UKbVvb/FE+PiS/AVY7Q1FC0rLUQZbl/CUu6fjKosGWAF
9umPE9wJNSxdlOloPyPP9e1wE32XWAEtlQRbPMPhOkRS14elZGX5KMY9oXPE5d81
8M5jRgfO8NecxyTktvwVQQy+MAmHswUHot4FOjlSQFthqcdWEENZkSdfO2qWwCm4
UMAko/a3AV8YAXMkFYCSt72sFDlZDFnfAG/oJczIwL9MJkfS7hM0SPAcYA2c2OBE
28H2u+habsiMGVcI/1S3+oY4sSvw1dMNVRR10U7EjtGzKJPhWJ+HQCcLKhXQLK47
8NHCIq9s/aNcN8TUrR0joayJta/ZuAqsLD+5GZfQ8WLzGmExw8Uh+ogqxJm2VAB2
eCCLFHedIzpI/VDfQkRJAceAG4iKtE/VQzZagM+OlWeKegYl6ssC/C4eqt0MWK4y
LbCFtGfIglHLxApsNrggYT8rvv998IXaxDnGmWbdLr4AiAlZZBZdtJGary5MON7c
pcqHVpDl2aaKKIlnwes92qgG/DhjktuHlWf7lrK9QkXKJzYFhTMrQ26OxqZ4H1Lv
ULV1ipr+kNLSgKE4FT25w2tSbee81TGGzvQt2MTCaNra9LRYg6VkYFtJHOEBKJRQ
GEoTB4gnSrdmOcEW3mb2ork45dW31DX2+Le8peyPJs6/20R0xIjoatBYabQJl2a0
e2kW7GlCql8AXtfaOjfgODOD9vocnC6D3Kxqakic/SwiC0BCx9+wSYr1ktTLVf+n
LV51FUcsu5BsJXd+PTCQxPfTUz0celp8w9TbweUcA4H2CgPz8EXpb+a+0NNehqQL
UYtCqXyt3qu5zycl26eoidxJkXH8JCMjFmxKea805+FbwehiAzZWLsfV+4PLBBlY
f0yITHMQW3d5u/Eio/lS02ulnfCjXRNmOmI3exaPI0QNsZZIEievJqNsKwqhQJu3
LiZ2zZVGGzxQ+CV85ssoOhCDQn1Ek7MpPmxLfcxzBA3TtRZ3afP0ZIpLcj+mw7P4
FFwACuCnGfdZj6UUimXk5D1bz3tKM56ftlKI723kaqFdnUn2EIC83a377eVqIXBF
Iup9IX4f0cgTl7+ZJpnnAJY+aiKsBjkuUQppklR40xyPoNccO7u9PxafuyCDiuff
6dGkg5tyKTfoHaCVGsPZT5o8DEfqvBZtr/W3OzzcMivghZupMlofQKoZ96587LGy
AuNmjswx0VzJgLMNPaO/Z3HHutLfVmerkgUZiI7pTmSwOw6hhvN7zDtb5Xe0ApgM
nEV8q+pbyCVkdPflJ/ZKfGtVUT7F3sXC+jKa36dCllhKPLS/F2okNneP+HYZYa13
oGG/BBTYq8qeQlwoknQ31C6dlGkNNWSgNK6bJY/Lr2c49P+5GAXs3NlCOTovIZT0
Lajb3qr65msmx7uUAr2ppdoQllrMpmgIHL2u6BQqp6ya78bTTYGgxfAGwOfZTIuQ
JTyPsxoqmZNLYrv4XpXFceXYBdcUyDeAIxAp4/F9H6BfhG+CE+ZTJqDhOtAw/nIR
J9NGmZtPPbWS1Eqy32/Ba+ZLyrbTVLlgCqzIi0it/qaPMhdqkdOlZZGM/BeR5j6E
0mjAy9s9Wv2OurSgOS4Pngd8PWqaRGXDdTzab1rmdqUUYSQDlWxnXTSzbGQcxOSD
qGFWZfAxSVAe9fBexDMmrGKDuC0bAS7Mhu12/3iu4s4QM0U9Xk4vOyajJ7Yd90IZ
S4wYWOUkRxWRGpIHVpraWu2Kg3HIKUB0cKjfoAtQyvCOIPaJ9oAwQ2Oin6mCXxqH
eE9uoWraZ/LpR41ITvD9/24APqgEUIFiMy3FsMtbBRGy7HPDS7ygDugaKyilU11D
VipjabmrgH5fQj76B5K5MFwOBj/5ZHtOXlBgI3Q6A6f48xe0G9n2RN+kjk+8CjyJ
/g9MRA+JgLEKPfam99v+iKebGzaayWDR46nMjRKxd3DTB+CjvP70GAT+hL8LA1J7
guW9PV9NSbmg8gjEO1HIOQq0fTFrRSB3VjL+ll34d2YXPvSCV8M+uc+zYULtqzAI
l+rquBwRauTfjhqkf0S7iVwpSOUvuu/Av5wYUllnlknvxrwazVnFNI3LQNEWNyvF
FgujH5Qpo76deuxFrDcxfqP3a7aGQ7oHzvFKXfFpkvkgx2zNg8S0K8TCTRuxVAOQ
AqCHiI0zLawn5y+pEMT/yFX/eshAdUKu/lJLbgqW85ELPO80XVozIZDiweU5mvGc
WOA6EFCpmM3Ahg8H8H5VJHSwNK5NW/Se8hZ+g2ihftKEM4ksZyVnwq2lgLgSqi1B
H+7L/SIZp0OeHKCkLwJMPNLSFssni/rdWP1bqnxd6hGa7srAALQ6NqkYXa9xRFsi
ho1xUQTanmOtt1+BzoeHj3OA6/9+NZWjP2MsjkrjL/87LU+2z8P7S/z1izDK97l0
b2d5Q/tWP9p6Qg3l+gNoDQ/CSFwvLq+PVv0fL8gkBMAXK2YDJkP8qIAk2kbsN31y
C3rj/yfdzognknS9yUkMiGJ1j48+2ORmdnljT0q73L25YmbQu+ld6MkM0ykCtsGU
Bcwbkr6N4fC90eZypV9Gr+b2TB45gVZqI3Tz71PXpAXzAqMZgeDHriYZt1y/NQEj
bEcvGs1YD1RirPJanVU0mKKWth/QIJhEYCj/z0PwC5CrnxCrch4i0nyroWDRB+qi
YS2TDNCd7tt0qvBiHFZd87ybBeFKpwLQqOr1Sh+Q4n/4+tvpHfGiARk+AGtcHI23
tAXtlCv83WXEdl3GOTJH5OC0aWqJYUjIiurzypZuC8AqyJqo1UzSJhmLYj+YgymT
VN1m9QwARRmeR2DSUfYBtnzrIlRNbyFsozGzLQtwwDGe9v5FhPvbTGJe/LcqXhYd
H9jC2K8HJXw6QD1JBNzkEnZMKOD4Ykm/EzbXSoE7ExcMVw8jT7N7I2wYwEgAaENk
xzT+nzXAMgigdw0blYPjce+t9qF6PoiubJq3ARetlEptnBjYJ6yZHvJrbE5q3XEm
lbTIKPd9ddqzawIAu8tBZm5x6xGH6MN+QEdcQWXSmHqJERVzYTzytx945/cU2j/h
0ryhMBkFOeKUS0gvbB3jrLe0oKa2i7bzJusnfDpg+o1uah/UzMUtp7zRiCUA7tDx
r2hUJLhfxspK/bzdAO3fpNGVGwKi1egMzMicQHbaMovBJfniBirklP93qOvEdd2H
58e9rZrIXpU4qWbphhihcRUBLGu4ovQ9EzZMBuVy7ojhnuI8R32TGPJPINxWeJr6
/b5RzvLNDqpZ0DyOjB744KMn/QSkqV+A1dZzLpspo9JN19DFAFJY4DO72MjnWELl
q4MlDAeQB9mG2AN0j5bH3CHs93+2W6+DRW3vblwExL3HRU1uPDnE1FYDN9Hum4k/
2MpDiFzYg9VM+WEu5e/LxlOYMOLCnl8nT1Ug5lJkWn5Felogi7WHSH7dQemv3Peg
IKmfSdLvOiUigxlmzC3j+jxO4Ud4jrk5S0a+u76veygsv4jQks2uWZTXlliAb7mb
AwL+hlPb+URw10cT154Hc9F6rn08ZkugN+MTISIn365ShwevfRW0xu06sHcZnbZh
88QcpkmVyfuTzsEG90x2WFAMhCPePtLGFPb7oy3oabZXf/yECC9fLH7Qn00DTLY/
7QlYRAzsdWDo1muYYDz8zIy37n2jgWMYl6ZEDae/Bk0KUt8/T3fLFjHOGOCHl/PA
TBjezRisk1Rcwc1SJNXbS9FhAB5Gn3D0NCxksiLjYQZF8wKVR01aWouZsn+ZGuTh
bWGw+DP7DOHqT5+wd5bpPcd7GCY8zFvqXP1hzY+2ewZRujmbA+nzEnDN5VSa7yxt
sWt33zTwFPPXwt0Fsuk9Nx7afHLiPpGIacoBbyHP2DmBY04lW80teN8BK8QlRr2d
PiSi/mp0bEt8of0MspxjDMxdhI2nMfPK0K3DRQ2pvSEXBqhCPjh+ZZNmX/vN/Hwm
j138G6FGmfux+3G6YNj4HHFNt8fSWKSFW1WiXSWT/FDWWYwirn23bzxVneVpCyLN
iQ+NQCm9+zJzSpeo8EOf7wHvGEbsvJjtTLD6qTo9mo11/Bimv9ScjPc6jVnIq/mq
`protect end_protected