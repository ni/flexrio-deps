`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5744 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
L2bRNdr1lLBT0eERw3vGlICEYF4XrVDvP9aT35NeiObEFQ5JxaUG8mriewy4yDGS
QZQXkpLz/XyzRh5y5PgvaRaxAi6OpjFLYpnuu+jSXszY1HBpJ4KejUoudvuK8/4D
1jB1Yipl8duKZGIJiK31an4p4L3m3SmB9xZ/sfLQvE6nTZ+bPDQF9FQKEGNoGsw2
XiSuhlptosCtV9EWRjWROg5S+kGWMfS0nZ6vB19N9tX1SpDi3KhTQAIXCdHFDBu1
2MJjBwN+o4q0us71Mk+73Ddgu6wPYS6/7kjCnCJ6uC6BZwRYVWiElwDrZh5WaRLe
vulPHfHesdEV+IaW8wLdPYekeuNQ2uKFsMo2pliHwTz7/LVjoIajf+/T/W6X4sMt
BA3Z6zH3lP4SGMnhjuwjgBpveyqvMPnIYDSSeKMVwlbRD8TjYy5eIYvd2FMd5o11
na5dxhKLr1fnpT+fJYd0iStm65bV9Tt88N0156YScNSzhjGIW8ha0MC6UF5bxpZ8
tIKCNX1SqOI0IMBTF2vvcFFJyl0/tSCDZpa6OwezoCNkDHVuElnAcJYrqF2o4je/
19rKcwrHT8PwT1LtxV7do0iUfkhQwielZ1SNeVYUlVjUnr8uV9BAE55wHjjuDj4h
Gn5VqkuqN8mKmhOoV3Dhn/swNiK8QEYk/OWS9e6p7p5MWuxXp8eZvHOban0PcTDk
Ku49/oyLwZvC8ms0vvC2fSRSxbxIFf/AwcO7PVenqtrDmd0tKaju1A5mp0eMAnoA
MwG0M+i3s1fJGA5dSuMxs/YnmoRvvKpo1bHOFnM7AbwvN+mANj5JRmEKIS5NT+Nv
ezkPwlYesPvoxoZ9DnGt7jaLFm/k6nCeUrlS8RQ1d5VeLYyRqDMV9nYCQEeFS/rz
uXCY0+ihu+OOn+hJZbW5OFvTZnwSziIdSmpPzj/1aiDTzoIO8HYYDPXxZASrArI/
t9UQnfrUgL+eEjiGd7seQdCF8nAc2p2Pp0LChudjtrOTGrUfMDD89ezOjzKERwOc
jHC/CYLWUwxSXFvcyEGq9y2ycem1Rhd8fjd9Z9GXcbMI/2f5FS+vkRfJd4GCfl53
yVEXrxSrQT8FvTBV0ja2jXTJMWZwLkIPbf9BgIY8YARiRsV77XElhLoInYofJ+ix
lBteytTzM3x6nomRjfTtKtueE0YgN0IhXJ19AZrLhdDlTWA0xtEzH+Zsb7aqQmUu
BKBbpSquPm3Bo3TqLDI2Gd1KFYDkGJz1gVpkJlPj/ljECGEf2p6L1WQ1U6HXSX5Z
s0v/SoeamV/RNg6v59+tTP5KTz6nqWEjcWaGiWKSl1U7qNIWa7iybGA6NW3gtAh+
adGLcTyHPadegCJMJ2CgbsZfos9FQxMZrOM4qBc7NpSt6/SyRO4G7txPDuqW6uUV
idDmjpTILEuAXUB8+MBUzZgfhycflryzbdN3lydLTMrCgw/YFhHjqyCHlOlOJQmn
pFc0Jcy/N/7jkcuTU5Ih0SJe9JqvQqqfqJMrZu/6DYFO4XmT6orlpMjuy/HOPrB7
z0txPjJ+oXqrEpSUynRoSKgYBhxQfy83RK5z2Snd6WCSsjGJwVHZTHnvMCkd79RY
bZAhgnGfLTICPkPSzAmQFyDg/cvKwzBRNVu/8evLuBtmu8v9YXxqx6cp1/NOhlK/
zL56SJc11B5arrhSnpLHgO3ZsnVJYmVR1cS0DMOXHEIJ9X089OKqxjhd9N3HD9QR
5FluuEaHe8yvwPwdrb9VrtTOgveIddw7ecwgmWToaXF1bHNxUM0pmS8u9w19Cf6g
xM4Bj9VGQYc7rA5Ww788gj0cLc7q8gjivSF+aCJqNKh8up3LIQfypDQJ3gerGsrV
YC1pAIN34+nV3xn5R0P5DJquYBpel5C3FZu6khSmaiwalHsVqENp9+GitgB60Ux2
fH2ZpspNJRE2ntpK4xdDe6fZWqWsPXY3WbvqcsHytV2rw3eye0d5ByLpJSTTEA/5
hJHnXfvs/J1khPpytM8qWJbX+JRNSzgIYK/EijclUzHH18qE9XQP3tWWrjCs+/cL
uDW/beBjCOujEFkYD4/5XJ3WNztJGVOtye0l6LOsUU/dibkHadanZIGXqI956ERm
aqoaqGJD/ea5aWrr0sDmlDVoqORrtaood9op+v0F+EM2j2WhhltzHBsJ64gpyVjL
ebZ2HWF5JE6l7RWqnzppbX3zBver3FevahG1v7qiXWiuvz6nlXOKfbdtA4KfQixd
8FPmtFw0sNBHNAYd8guki9umrH9DJQXkZmjFOJ9R6d4CWvo7JrmW6bAkbqAw+VRd
dpBrPgB/d4TXtHyu27Tdkj/IR2jMrKf4ls07cMVJM/xkD/kkutDBc3z1eA+0yAbN
lC38ll1jb9To5oSdP2zb+XzkBgJ3OEc6D5nu5FpJWN34FuUDYuY4QjZ/xNcJDYBI
0Adk5GNcCb5eaSUqIq+lytwnV4grRqnjQy0NlU4nbAnQQqnqcogucVZ+GFifbcYe
1TVeUE1aZh9TiWGjueOhvo6z98D/uQrg0czcLffWEC3Ot4u/yU1cCc8KV1egvQF6
DGuW180Fr/9hxydF+4hxanfhFktC8h0Y/luiQwZJ5Kyydwg+Us82J2oK71G2P3N6
wmcpOvNqaPA2WP6EHHtSVjVjNuzLPZNGpybq2TDdWmK4VGaYV4W2MCGtbeH1tCqb
JQhkVeGWYlcn4e5330Yyh7cyUKiZ/uCRuw5P06UDCwUNZxHxi/EwKfDBZvTTWvkL
Cdu+s38jkIuFpBpa43RmwD83nlez50JDzCJnsDcpQnOKP7TIfmUvdx5z7QvEv39S
XW4rgIAgMuUF+nLSgIKapLxHyC2JEfzpLMHUZnweO2LP4kh+83dbSOLn0uAeR85R
DpyxyraXHLbl1QekGIj5SemNWdhONKwasVSu3bE3j+cNUqB+/J1EL5xL0OAEBJ+r
/paCV2tId/WUsCeT/GQffgEMMzSfpwj8SA4/f5iZwscZjpeDFO0adTyElskKl5+a
AQhE2aX6D5RjnP4+zHgFCIZmel/z5ys6zn28oqMadLBQ9uR30YZNgOkMjg+7NPnU
7WHhOdPnduDZk6BmhM8WsCd/OvQ8N8eaZSQi+VqKe7Cd/rp4/9FACZ98pZfvSYGg
80aP0xrw8qoDL6htxgYlVmsQWe4AMvB5uSxQIOKIqhG9W7gXl9q81vjWYf1Gxf4B
C7Xql+O1rWioSnprJloFoOYuHxXYwvwNIo2ZWT7FoxPqfG7f9V4iLMi5D8EYGIOh
dHx8ARCrAo06YReWc/z/s3wg2pnt9/T1GTOudN9mnR4Jir/wgaxxzoZJj5JMiEy4
SSv4XL4J83lX2kCyiuUyuYM1DyT74KbJeVPhyrZOeegyuizB4BG5/JTDX6q4EyGq
P1A3PH6MhrIyTW0peREDMBJPmiQ/0REYX/WhKpATvkEqHXXMcMd04326C3LeKpet
+F/+0QYeSR4y02uW94xuUmMMAzjlFjQxd7TeybTY4OJtw+Wvcel7WBoovArwXdl8
s6wjWdfSfqfetZNbhs7TEi7I6QD6g9maqkpijBMl+cEchi8n3QwdvAXaweDZvkQr
5vH8q5EXyJHDEuIV9X+LN6XmVNjab9TCWcQDbmlFg+iZAnPukt6dzXcbvwnf45/I
VVYucjUIpfXw9TJyGBcEmSLaSPa0tF4RTljvF5QJvoM8vUMHG5QaBCMYUI9MindH
w8eO1eluRl07JDLU6zxXWRBOCq76xakMrOPdGX8Cjh6Ts+qGA9HB5UPO/+YKvQ5w
GTTFB1WxahLfjClf00rL/BojQdefchCTuIAGXz5Bi7EMbiG84KY1MuDjX6gH5iEo
3rr5VJ7K9z2NvYLObKgFBgU0AUZcqFxRVMBIMLA2oisSaNSBJvh8jNMczBqi0xcH
0C79wlIzdBAJqbnP42KiDgUmE7rUX36YnsDSM5bzs83Ov4ywxSGGB1JTA0S0m7B/
fK6//do1C6QpPZz3fEKYM5DNN12DA7qoKe/YO54NNRIq7g+Jvk49pvPhKhcn7XHx
bQUyFAHMZFL307Feldr32CWxj3891pPloF4/HIAtiGb/Nl5XMDyAU4IE88wUVElW
cFX2aB/YMyiA8UI5MgjdJEC3bcS2qhvdsZGipyHPjTgiZhSYvjyhrv8dUwsBSe5N
fyQrC7cN46pLG+mKkccqozgiKN+0hPiT4mBOgSCJSjH6tni4kqe0TuAqptNgbrPR
Z3+4mQMRqKhcStWH2e2E+ogeHGWV4zyGKejzyEjQf24Dps1Hxlp4cIzQ77wG7ViO
4p7atI+QZdf7cHSIyMxUtK9yFp03vjigJDYe98N6N3LtN49jWodMb9B5qt2sTDP0
tdMjXEMSekscWFV9Cq4gLpGxddfdeCROGqIxjHi9QHs/T1Fkbmn8ulGDftiIst71
umqIjy0Ns9c6h68OAvhno0WvdG+jwaUi98E3MAgC3JM9Zk1OhX+ecVaYjTQEBNQ+
getEeiig9z5bkY3CS7wKrQ9rL8kK8I+D/doaw0/0MOrca2fivFk3idWfua7IczLY
S9AoHg5+612374uBKBXhici5LOP5cYlGBjdR0PPZ3PELrPNRqw9mnENKdFn7puB5
e/QiTAgrUiWGTtYZ56gX72ZmnR272/reUa5w3PUv77kP2BUOA6iDnJyObmrkM+es
Od+jQ1db/Roxiovi5vE6ChOjPfXcrCHNtpteUCpvP8LG+GxzdPtmqXtN1fUOp/sz
vM6q53xeX2C7dN+uLIJjLwuwCHKrHVWOXHpF8DrtB5fLqb93AxRxEzFg21ntaEX+
eKRfHPOkZTwydkyXzIbkrQwq7sY2rcIRexNtm6Ay3Hz50vYrPdM2+bjZ0fAABAAD
hXsCzY7ZisROhEncIBE2GyOOkQyDv+koohJYp/qzXhcOuN56DCC3CEFgF1cr5mx9
XsG6fNAN4mYBzUWtVKbCeaJeYCns8kzUl+aXL+jbvqYKsWGzU4YoFHea2+Dc/C56
omuOn8m4WqKL3CTzELzbVZa3WuRdaxf9Ay2iltNQ15+lNBdv8MOW+I8bRMQ5hqVC
uheeCEnfQkEP0Zj4d0wr2MU/kyvzzLePS7RC7SdMMBUPHpFwx0pplcabV4Vf2CUN
+Rex+pv2i1POViH6lxMhEHjwYtzTndY1Q5wRVplVLVpxesKB1kY1oD7TbpLChWXe
KELfAXqgIyeqTpRbzK2olF6UBX6hOn1VUp0Q4r1745OegHGzV6xQ++Cp9v62BMpn
mWd2JutqOVEMqzBp8OGZ5OfEqoi2BwRYe4/IMxD21yR4HheIRCy2V+MRTSwjLeDY
yokVA4DlxTEcZ5wrpPoZDecT8r11H3jT66eXMaR/fX4Az9EGfmuv/II+5+hXLi0l
H4bM60YNOv0gyjaPnhP/C6vD3d/ThaEYeaZVDOI2S+M1YCg8XzxB+FDnrd69ln/I
SzzaEzb7BFhFKrbl/a1wuVL4xuhWm34jGm5/3hWhF/O2awLroFWbbFuLCwrwUT7Q
mH4bVzkoN1reX3I2OyMzVYEnjYs0DfnFeOLlJPiYukeRehSDIhwspI+z0W0dT7KN
G7T9WSlAhNJWu6ypXbsHYOsoV5ekh+8xTo+P0n7FT/jGyexdqVfEh9bHSS0Hjp4H
c2VLQFHgpUZpNgLFVOUGJS+Y2EisTeQ2EIz1jA1s8F913mucfltW4oMtGwfgrbw8
7WuvpmZZyomLQHB7usJP91wO9FZxO2CjMmkFfGl99YEmEsvfcFxVr/Atr/HsCnJO
7VpFoYW+5Bualk72ogm3CeteDt2c+d/1O9eXmZrW8IUFkjfiZqHh2tK5qwrkGfLR
H9Trc2zFqy2jewbHyF7E47yBoGIEeE2xf5vB5/GGMwpXragZ+Uoq+rhAWPv0vkoO
cXC+nFj8QeYWgqrA/Trt0MwfPC54qUfNEIvWzZ2vOi0mVzgncOBjg9sRby3LlLil
WIMnfza/+0bm+v/AY8RY9bxzIh2lO3TT0vc7o4uCisnSzqDx3QL5s7kSU/o6Cd4b
zAGAVOYhu+ndkw0G/sf06RXCN8TPk+XhY2VvljFss0GzINFHpSatA32qzHQwofrH
keLLIt43+p2L2IdDtKgflNLYPkxJ4bbZscjwDPy/uqUywGk8Xoc8oMuFSph2Rixz
FNGdGHYdIDG246PtkU8RCjD+qq3VXci6d8Lxij9Os5AkMlOZOYjanYn8FkD3l/zz
Napa2TvYIgZhtRlCvXTE0tA1FHjx04awewU2ZQAw3bj1KkieWxnoah8ZwbuLUHjE
Jsn/2BcT59apNT23TZveqaL/1rL7bhVV3YDdpAI3mAs+ql4ztN8ql6F8WultdIWM
NNjSzVr4l9RoO2rVBGSyYL+nzTEtGjeL4Aq3en7jA4UIKTwXr9uGeJIiqRc0dhlm
UTQdXvILuN4BRIFapL867GaoE3Ly0uH50qNbewXEzmHjsnAf8rWhyyFlj8TNzgP+
J4M5/D4W8mp3xhDGVahDW8WB61n8uYjRdPOlBFPnqC9f90v6GuycUQOtsf0wIUgM
GMk6hHBeOSKSM+jUEYS6vda8Lo4ifATrXuInF9eDjd361GjFL7OWmZKjdb3hy4QD
M94MbobW1NJFi1744On6atEJXDd6yFm43QHzU/yU+kzXis7Dv6itP4Gif1Cx57ia
AE4J1R7ykh0abd6WkUATdKuvIIsEVYdXv3yyprLrC4KrWqzEpz2I2F8cP7BsKhGd
Gfj+eKZh07Boc++mKWSiHAFMW8roxT5DYOQBbYF0hPJNoJ0LpmaMkq8EY3f7n9Gz
CYRtPDDyQLO6iuGDy0nLnpi75u+uSb8AYhkRPN/3AyTpu2XbYRtMeXpAkQN/18el
hEhK+sLN7NBJlm3/zSk/LRadnxpPbRSSbGuohvsLSmkaFieRB5UBno1vrAmkaoa2
awa0yQbi5cFSPqKymTR3qqniykNTlxeJTIk3pOYOtzhBxQRafcORBkh5RSpMBhpB
xxl/S87t13/969ImglraAHgxOk/0oqBZnJLaar0yq+LswY6MVbRFzp8+ZXAasvvb
bt9QnMFEcUqMeKEtvpnL3TqCDJsCx8y4TOIEeaaYGSgLIjmpzKguT0Uy+0qRggd+
wYAW2Tu6Gm3o4deY+J06pFzg03oVniMjGUl2f2PVe4e6IHauHC15OAvVQ5TYfR64
s8vcwmgWeLZfZ2THc0hpBlS+C/Ho905hv/VX5aDerwxngzJAu9wDKwosHdHGvsV/
HNtYyL+YrlKDfRwdcsITXlBtW1BYaPe6MfzV7wJVi6hVVGZhXvLkz6Xib8mg4WpP
cEYocZNdOe8pwH2ScCuSuv6sJYIxhpsLBvStUnre/P3KzibPDnDLatW7j+0hdZlH
B5mhtbxTC7SUZ2yOYU9Wf37z6Bj5oz1qAeXjF8uTrtb7SI2ssVdTm4LB/rJ7gVhc
AyxUf+LLwGq8VkMmZpwzpteC3I7sSbg90+F0/oFEHwuce5dQakEMrXtL5mpv/4TY
mr8bz2RHt1/9f1ZpNjrw89Ka5nY6pOP2wgB9yjzUKWc=
`protect end_protected