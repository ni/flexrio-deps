`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2128 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
CF3xqpHcS7h2Fdz4qp4osZlfFVP6txHRXqhrSWosH8aK0RbBOlMaFbYI1u3A8dWK
McCN3teMH0xQvkneHrKBdvzzxru2XGsBbRZ77yXAHWrAl7vhquMP5/ha4UEITbZr
UOC7c/JGFKbxJAIVYuFCxioEB6TeWUJ1ngFbdf+hbBRNWWUPi+hHQL+6Xo56KZLS
vrPXR2diE60p6RWgaxRLkUe/JhUN6MgRjOD3fFWtQzLw+3w8Jc7fvMl+/wp9G852
3+EYO+QgZDiU2DTCIUhC1ShZBGejRKUTfcfi7e026l7L65Pr49KX82vZLr/zVyVw
eYtAIQnY0oYY88bgcI5H3aTEv0psHD4wQqTtnHALsYFoczR3y7nUWYwr/vc5dq4K
IiZLejv902SlsnrzXtW6yGgMDozgrwL+uBHdbt5Qruok5cEBFE6OuLxs7m57g7++
/gM8Lwyvd0MeFS6/3B2NKhUUBcLLBn1W8WIkoU0znnFZdGJ0nZugumdKWviOGE9R
5znszshiZZ/dVET1FwIr+J4GCYC04rfLoh7SU4VJXCEwGzXA12wpBq5jdHolmfWm
vrFM+SfyOiRaflrUocTGBbG9khkDTEv8LWXIFRLU8R8VqjTs0xz3xaizg6EBiBu7
QH48oMtxivzhoN4snHxRPi68hLZZhTMVAXEDBW53ba8K/txQaw5PeVZ6mMx0LdAN
pvJ8j+k5PLNpG0wcVJkP/6wiPrWlY5rvyVe4u1gykE69DEC6gTW7yBJN6m1rfuwr
cKIogDFHR2eykvqyBQEtyac7RBGO4KyNuB4zFCKpzCcHR9ErY+bY3Hcv1nd5lFgR
KB5iu92m2+lzIO9s7aTgPE36mxKdW/UhA8dJRDEs4FBYODPYhWX9XhU7mbxz2o0n
WFhintD/xGkMKfrgJY1tRmitEzKklGEHyU0n5gWrExfzg4WOutsVpE27zs9uIPAg
twuyeAKtrNrQ0vpdzTCSCT365t6akkNvx5+nlMMk1XXVb09OKycQy5W63oEt+ynJ
kKNyK/we1LW6tQOseILcvn/ExlfTU0y7bmUvwBsScj2toNtcd+NJsSmRx2NMUjqB
CDx8AMA7JatgbFVzE1476uKKBYN/dJKgySam0J8uEqYGUPPkvndsJjh2S3SuI5Iv
MSfq2IRs/8bmVN+8qo7S7PiST4rGox7QHGij5Bf51/Hd1Y2S7w//c0VQus03HMsQ
IZ+pOwrrqmoLzFz3iFR181bre3GzqEcWlIF7gTakTEA+meZOy12TRoZxgCrhOro6
VGORPtKxR4uzKZ2/Mp5CbEsOk2IcXwBScjdXsn/PQwajO+PyZGLtxqhP4aRa67fR
QzZ64cdUv0Q2As1GcoVZ3ylfATcRdgHMFg1eGqdcoT/YYp/E282Svotq/gxGfx2p
YHx9qBFrIW/gffF8m2x4c0r8oLKxATI6HGkxrShaVSizctFpNY9l5DCZMtirsS6D
KrQ6LqSJidQD24pj6VW+IJWzddKvhHou7Fr92gz2U+qcfOd7Mt6aJvTcF1aR8QYo
xNg+38NZMCx4ScvrlnyRbB2LrZsnAqYOAUqbWO8iDSvD/hytgP3IpFqjsikrImGC
bd0xrfELUcwYlFY9uHrs7aB9tH2XWCXJL4oPnzmJEuEsp/mnWCKeXkj2uGIeAHhi
Upp9SpYW5HsNzE+hJtIBBr6s5uE4X6XC5h2fyWXHvHMqERGDv6JN7xNPLDgAgDfu
5qC9nIKzgY/O6FjyeRL/Nnl2hlo0Re7VooQViMVzYqiQgbtUG/L0xwqfDg8pwM06
Pb8ywVrAW+0Ric/eKjXFOR1Vqf1143OcMyHTrLRETdABrap10E9T1BlB26IR/KFs
UzwOp1K5Fs6akAR0uxjm3ns9Hry8oYnsRe4PGHbDwiVn1I5oFwdynmq/vtm/se/0
LGeMdAyVLdxhknEnS6zPVO8yBUQoY9no5gm5eBymI8T5bw9we+XLSWMIUnuHVEtK
jsaB6U+PHTbHWaLJcYevpBmlowIdR0sUtnYPk7L7PouHcOxbuUJNO0KEhkGkzI3Y
a1dqoQCfjvGHku/OSvDiw+1X5knmKDRfYS5DQBkbvCJOuut6xPcLHnj501FzfiJy
nSb0+fmHddO0Qwy5rW0B5TBzMf7V4V9UVwgeS7ZEUMC0ukEx6AVGSeKGAORCeN93
J/DlGiAjbD53JFUhqBlegs4nB2eNiOXL+Y5zhUBOblAz4A7JMcvi9WCere15bE3o
eCxAZIRtUbG+zcH8qgfrIwrTISFxbywJpSqB4bSKnxBDVmeve3jFIrSsdi7YVzTL
pe/ECmOqoEM2Rg/PHkkSikw0nBAiVM8U/JSvz5QyvF9qlsvQNixjOkKX1HBnS5jV
zpE/vGp9u6tqVWgH+aIMrKJpVQYZZ2EyRZrSD1nuUfEijclZP92hwUAQo2zTQufa
j3I9rzFnLg98NFU9g++9MpRgtDO6vNXQqpvRIVoykq1vuA5ZqCk8ruU3gyU7ag9d
T6ykgcnNL2QvuEacJ3iWeJN7mmIYvum/M3nvAoyafgIRZF+EDqFAdOhth0lM0izw
xpnGfN/hmujzvrTyclNNVazsKeOIif332iJb4nwzTqCexHVdMeZUOvEyycRSbqgI
ulB1s7Zqa6NN8wj+qhR4zvMO7Zqq0eDqxaBSQMPVnKnSSUj043RZe1mYDPDLna47
6TInuH0g5zfp/Y1HnxL45g==
`protect end_protected