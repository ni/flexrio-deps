`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 20704 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
ZIICkMu+S2rq/yOQyqhpupmJ1IlVmAI52F7eUhB0KOTPlwVodnCTwPAtM1OcGW8d
q4EsjI6rqg12iBPUAflA/HjuiY0C2eZXsfel59l3rWARlXuI9PB7w2P1ac6bACD9
TgpSzUc84tFTTtDnOZ9iE8QjGcJgEWBA3D0o/Mux3yC/6b5QjLEWs7Vwo/NlJ/84
TEeTHCn/LOgDLgQbg5nmfu8xmPKMwxWsC8txdvUKLVEjq21ALbkkj3RS+f+pOcpt
M9TmW91yR5FRo3iEZ+sJwD8d86JRPx1B8HnIzPaD19CRUbuO66TCFKbx84JZuAuW
cwQhI+Tek7cDgWGy8arVr1th9MY9rLkZ6CeUFkCxacpJ/WKJfB7xg05Ego0/qvVv
ixADyLQ6JjRytSooPiAEtAxgJcXyRFnc9oketIt9qcuDoOA9BTBOH114GTGJmBo4
q79Aa0Y8IlUN7v6OqVT9AoQMj5nUEeshTfnwMmHRBugPG92JVHGzNDDzjM+jzL5u
ZC5eaMeDMTqe5rvA7JtOii4h4+QHlq8pT54gnOr///VLrJAxrnhIWzqlUewh6Mfl
JiebF/Gxr8nyJn031vCmb+8k4qgsz0F5JK/HTxbAMq0OJXAjCX3zvH10x8fvWPnu
6s+T9k6FqcnpHGzNdn1Cdbabd1+qKRl0uWE6qgCraqX60wQ6tz8ttyFObwk7vjMq
jPIkYz16/jMbkfIP9pg97MAW8uz1RsPxxOquGx53ooj6Ae8YBTDKU/OxDWEGqMof
cf88Qgb5i6QaZV3ApaAXtUJcPCi++nEupuYBI8xtcNxVa4bOj8nxwdjx2/oRk7J2
PWCHVJ9hHiCAMUYLN4zZ20j2xgtTDlW6++08QrUR5frcrlMHcAyRncqqQ73yzs8W
LeQszkEEDEqW0yYx/NaaB5kbu0njhQctllve52C61Bn9A3YxudlNyU0gJO240yvN
XRV0FOylzSxuQycsHVe/TJpONXqFAQ3oI+GZhYWYvuIAyR9C/cjJerns9qPi/Alp
zJyOHDrtHoM+HXSVxXa70eZZTB7vuCSZEgAECfUdoLkZ1lja8eucfWDMrUBLwyEF
ymwjXVIEY7c64zCJJtTeIERwsSbPyWzC675V3ERW4u/ZA0CBXz8YhEvNOsaxZOpQ
K7SXwEpFxUl4RRNx80XDngqi/U3C1BzvkIqjHv9kI/9faUoD4d+t81QYtlWbHdqP
O/miRZD77vtEI9/aAwATIbp8Qte1PXrWsAFY423dQjxtUgqOkGaojaa/2smxujG+
ANXT86cDHHXj+W2lOHy1ndeYfvHRptKHkjV1j8u8PFfVFTr2KXV+4mmegtcLgJlV
s5KNPF49LFFA9FvHyBz3EbjvsMhHG70FB0kW9VrwVpt6E3qsL+wVQPqvZapyLHN6
ybVunYuGPopV/I2xYBG2iNBKOmCzTGFErCub5xAWF3CMn8aYa+rCjlWHsGvlV3IF
eP6swlkWtXT9GXgoXbUtLAl0e7E8wbNPYi7AkKkG8kc1TAKMfFItJDbANxuh38de
oo2Gzg8qtfk5aCzoOCB+veKShdgpeEa07Tx8MEgGm05wf5pfzT4wDaDrQDZh5Yra
HehiPUk3RV7CnbSOy+0D7LLqLmP3VIuv1IUhSarAmM0HWY06nHxeIwycYTh6PGor
mUHvFtDuG2RjkYoLM11/ve7q4uxGg+vvW1/rOp6d6fIQJy0/UnQtqyW2LqvY3Q8w
pa/AY7oFnEXIcTxj8L2Tpo7+PRw89U/msrBh0TCb04YAkmPfi5SAoJSGd/FscdEe
kjyzc7x/3Hh6xOIP0uTVMNGO9jc8KsYE1+FNYp5Pmjf8XM8lAkIAKAGeMyJne79w
ASyMw/3LnHG4NtFkJlyz64cnb7p0NQL6uJ4cjV3hISOd6tbT+tUokmk4BLHUvP8X
rYv3SdGwWwkMw66jh4y4ndM8eYMLkXQvUDPsUmuNlOihSAe6f44zb9VoVifk9Qi7
O2vZQNQSKHmOfcVrlR6u5Zlym4EdvgLmGlu0bqq9XHT+PQ39HUI5PwrrBb2qnUI6
gORjD90igo1bV7zdDRtmWsvaStJIXwTsY8v74/dWj3DAuQf7LRE/1mtmgMEUbLEK
TjGoZiA+4nGR5ndLpKliekzwcCmrxMpbBVHor/hFeMLwHqiK3zSQxdpp+GomeStU
NV7dbhDvmZ1lS+duFvuMA447peTCIr+nzy0tD+RbUXF5zDJVWMY49+L6Z98/dWFu
PcAR6JcvU1Wk0nFIRBruTUtIx/tRLb7A/qzZtyl5TRn/C2EM9BTPZXf9XiT1kYyA
E/M98+KmqXh+SwBXzalxvQT8mQYcMmjIua0t7n5EFCe9BJky6d5CSJqIGg+PeGTw
EEBnct7O1RjKDRtXZuUXOiCehw1gCTwXoqFYfuDHVesgV1uCu8r8UEJ6CxgCjFhH
OR0wGbzjvmTrwdTCVKr+jNS0q1zi5Eu6/5tCfjpwAcDWdk5jm71tlGSD5zgD4Yw3
n5LNa1PeSy6wEp+lsbgnj/B/jqt//2iEC+bg3a9a6J/oxuozcNOrGRwmkCaLZ/GQ
N69XE64xHPOOqKZ0JM5W8WXGpUQ8iA3Fscnxw6Z5QjNntIOS/yO1kcaMVfAGBpaf
u/eIqO1MXz9/1pDcYoVk+dIvLwNY7Os04YKNS2rXN+N++THQm+7mZcTcWEWgFU67
Y7/ejTssprUkhY/ijxD44wzOngtab9+kqiI23CXZy4zF+Y9JUeRi0OxTZ85lNKv3
4C4VBxBUmwSQ/H1qEIwEpA8Edrh5IJaC7jlSR2ZMBJvC7TVh0CXmDxSz7n259h8n
bqBaDp+qUejqGea84IEgVONxdd4B6kJn44IZRA1mnH/OF7eHTsRsLe9JVGlntPxe
pvmGjpMEJAAAW7wsQsTPFjMABLZQhPp7VvmwIzoir6oesLGYcdlwf5SwHZhYMKku
oTpmNgVntcbX3SBhPKmv/PvSqjFc9QIAlCye5AYp8/GDF0h0v927MvCdxFkiFbqd
lXpiNclleHUD+JyMkvD67mEY6cBJwtVax3dpI1QaEEQ5blmk8zHlSnzCAMQyZWc+
p+83t43YGrZ1rQDdo3QLEdBbCo11em+YBZOnXhxR7HEsDX6tyjS4MJ4/eBihkYL1
yLr6As88scJmOeWp7egd3I+BEYsLG9i8WNWmcqIILggwF9z53TAWexvan616rUKV
imklgShmHEKzCFPUwhALJA0szI3H0Z6f6v4ycDhIwX4lXAK/WrbniXUI8u2Mz2hS
rqkkped2A/Foekt3J4cnT1B7wUdES6C4/XfD9eHT6wCW5KFHH/D//SNhlt4E+jzt
+qlob/VSY/1gNNUyOq3HdVDsPcOeIM81kw+QG+2QKgyKjnOYSKBRYF/ZDL/tcNAJ
ZgYfTTGU5Bn/S01XaN1e9ePwvVLG7SN5unhdA1rZR5+0JABezlhIuSiyHrNmNWP3
Wk6KnC+pXCRKDnktJRN9D07oa3AYYhtgFV0nGYgzOays6Q2hcXiso9jEIIpkyXa9
r2qopSl+I75t9gX+CDp2505qgJqkleZQbYC6PfYHSvLOV9vciGArSFkidGALk4ph
JIrMulyVeWTUJQ258q7J0pMOLciqkb/9UMVv/3AGTiPoVQ8uGweEXHdCUT2hZPCN
yNZ/G0Qydy/6Q2msiqeWWLrcZr+bmLXokxInMP4C+L2CroYAI+6ldSATyg8q7Dco
NMq4lqZKk/BJC0+iXs8B0IrCELOUEiSpBjok7C9nMrY5hH8V78R8bAke5h6l0ymw
rCg8QETfnhe6XRtx6nfGKOQ5fVCXKUjyeWGTTIxAQrinXYGZ8ZPOOCxN5XFpzk24
RupLJfH5wi0tsvy7+qt680TjqT/73bVnuu5uRHAr7sUl5sgfKTwGZLEWsVZL/Ump
JYpiRTkjUxBi/OmslCKEK6xe+xmCK39cj0wVaah2bYjaxVatvTQ3CpIbNgsoZiHK
f0AmX4iIvTUGcGci4j6701qC0n0edbUJxAH0XAv7ntChphoGNLVYaaBjFpRrQA+z
DxW/+/b8j9gTMgiSxd31RWjB/9upNIQ/cT7PiKlxd1o5FoQUF0brig1t0oVc+jRK
uIZDFBMNDMlIuyrJL0ABrBawLQmsnF6y4hLcw9jeDNg+KuALZchMhAO/D+RoCUjC
2rrk61NdMgWuB1lQbRaKT8oZZXz3qBEcZWmNN1p53ixGxUjzH31aV4AIveGCTlGn
Mi7pPu5XzIYfvR1a+XfiCjSnnnUeyKYGtAXszAjE5th/t745bkDPQYtzXGkxmwua
w19Q4s8SbaXsnKrvk+OBVun5NsOexndZwCMKH8WmVvUkBICd755P72b/PBtgeaXd
Yr+BWNwC7gn0EvoFIFcS1NAAW5oRaD2d0S+h6GyN+BA+GIIPpbgRkR1lWID7V1ui
S28bksduRMRkSnMqtYZujxKwl+fYk2KPvKiwdVIbYdiRpCeHIAspzlVssmYgAopG
i4h5y4EIAgXZvp6oURXgzeNMOV6hYEESsCyotU2EPSi2QeDjz7ox4mkOXPh3a9t4
X/ESMKWOIzjYyYhZHOv29HBE6Om1kosURv7VPBerhozPjnLydNHG31EFFrm/ipeX
dKdljP/lJfHOuCzYkISZRZLcJXRn5uqHEweWGqipe8ymzYUw5h1/NrS274YEFlWh
lodNHaZbzW4Z4u6ZAlj1ylsxtMgo1l4+yHuxZqO9dvm76sCaErF+BKPtdqzwF8hX
oe7h9TAS6S6cknL3F3ZgnSZ1R/vsWnqdETbg/McgyfidqJt/H6g/ZYYuBsAMbENI
XIxyKcMILYZKY7sLf3ZsZ4EqnWK4gxcqS5KvpbrTaURiVMbm8oU/5L7FKMDgLkyT
uphF4LqGNbyuE1u1ImfwwJ1+EJw7MpCbaLg9c4xmPEB+ToAK7LOzDZ3Z6QtwTOaU
E0blIFkoGo5NvRBeJWcyS/TR7meDHRdEsN8jGXK7ZitS8xnX6wjn56MVx1xYnQfe
9Ch3Jalg2LBE/3PFUK3/B39y0/T3JWXFL8dAODE5Gu1PptVjY0A+dGFqYM02A2c4
AmyCFxWI/Vxu5TfPkBlQD6+OMZUQhEylYmK+JQlqOGA8FsK/gqz/Yx1KaRzPKes5
/dagKx98/4bupvvzCw9hPdvDqSg1RBXWOkCCY1ldHkLbiQ3ATBS5hjU2mpmnU1q+
fO+6vBTeOfYpO/Gif7DB+OTvkZPJaHiPlJmPGvxVzu4NqHKa+zw4kL/AtHjYjmey
976NMnYgA1VBfqhlu4wT59HfDMoSpU6YY6APoQ5HPyhqdcrsj7PaVI2AefUdY+oA
OFpPggvLyKpk4kcJGW9sr1tSnUQchV1BagtZtKXheK1Sly0T0vKhPg0YdTe5liXB
xGSF8rTInb23JhYvL9UYlxPRI2cRPFcWItERsjGEjtZEMbcRp7f2fWXYV7CJbOhE
L0jmHTFVaDCJ5bkiwqHg3XiNgBUTkl/gVC9O81v8czMgqW9fxTvj2cYfgwiVoogT
69hnCNuuuQTBomNHjgobHx9ajJClBxA5Tz3cDmGjArrHyWb7IOIz2ClzTe2EAHG2
FCNdAqaOdgpjxnaGqOSqNvglldq+34W7vFn4BQ1zN5xRC/DsWyO0//FVrxnr7Y64
Rip8zxMVHznLUTbER7JFA4Sj0Q+nj/eKQSukn6dTGB8QCyDuDuQQH5VnxjiTjkFm
BW7/w3ijnEmwDqHZLYJ2j2REfd9CZg3x21Nf6K811bia2IWfFMH2JnfYxF3F4zDP
U9fgzRdHPIYEfhAx2VxgQexLCUX4efCm+QMyx4mYOWaL4r/NOcJAg4sQXxWm3MMR
mQq1YX3OyE75SmFHECVOQxBuSLvn5xU/EpqWhpZ68rS3aZUaqjnLcbNuEaTwNiDx
8J3XD0vEEZglUoilt35JmkrQVPmeOHZkRNrJPERHJ7AHi7cGnFUd1VJggyTf/xFT
X9IWagQ9Z+yu/UafmI3lWgeCokj0U6ULHNgFOs7IjUE61EFl48LQdfrEfL3aC06/
qnjDXmtUfDZj6aRg2WRa9Vj2KusdkU3DUFi0JiynG3d/6R53M6xPY0QCMpffvgFK
bBKBHR3vt5NevN84ptoSG+hNQjcvJxaZHxY+V+h3midkk+YnYKa/NLr8sGHwR62a
XHHP+ZPd2m98uobrEzULVwP7+iwYScmjixcHy3Oaj3lyiKdoQKn508r8ZbfTaEc0
A3WDMM0t6Vur5Kb96ZNkS6fQTuY/pzN7o7BmYYdLASnPxmc1/kYfP66L+bvJ1XIH
IxhNMyP9TymkXm2fIFrP18x2WQV1mTG/4O1G0MMdVjFieguiQDzopJ+6X/kduTYA
qY5c0s3hIa2YruUea/Cm9wuU0iq7Z6kN/ZfIDXnUY2IMZlVS1hcdzteqd5DOlqOA
1yvoS4VY3+oY8v7gDz4spG4sky4lcX4Nievtn5hSJkDJChksrclJcAD3X0hiyGnX
6XGo8VUNc42+2dzKc+oWpvqDjeUvd3E0BtcbfK2p0uRHbOsVPN50F43xX6MuXL+4
0oSl4yYLLiIieC66rGrbnSat1uCbeHtm50seT3tqLImjPBzRhbgOJCd768xDKuYO
XFwGCY8/cgZXupR7LYkB2X49cu5gRWhh7gdhS1Wb12cMCzKz1L07A70dcFrUx7Cv
FF0A94y/TKBvoJ2FgMR5w+I2O9fn9M3+EST0UoGbkzZ5nM9BEY/u4AjKIWerJrxA
wJgo6mgnPquh6cRagiVQBngk4GQVxBH/or2oE+bvuDSM2J90qqM081Jl5Tj6wPOB
d+4NWKrgfXI7j5Pf48VXVOWjyPAf3zf3214NBDx5bQdlzTtImgni35kMjrRaqAMt
9lp14GDFZcatW301xr6mXxF903Eyqqfru0WfqHX72bcdaADl/026v9O58AUBZSkj
1R97TkBafacegzEPiLF95pmKRHvruXIOft+MxCJKn8qQpDf5BPJrXFiWLK0lWtAy
4yrxJ90+9EcgZ5EuXNpuTrH5cx137cu3QaGSlelrlraSHuoqb1pxaBjXxGNMHRMN
SEx6mtv9Cxc7JXbbI6lvT+AgzlsFLv/c7qegJbqkMdh0UDeGXcfDSyUh3sTj7L4S
MWeFri+nPHfCXxdf/HYc34KnBZ3W3mIZJC6OxuN2AQtOmsJl0yC3EEGGVPSHUc38
ismJYn4UQ+clOhqi/403nJc7AxYoMUMqTA4tZm9hGk+DvAar9hVLAWusSzeNA0i2
hOVnfFGOTppXRxPPlPMtonNFbqr7rT/rKnn+cYivGs5sYwebZUfmma2N/v+VrLJA
fdbEhb6/1jcefEiQNSHGsCcvRSDu4ht7HHl2Z0c5vDu9rFHVsbftKFPFRFb/mX5z
A3FqFALIxKu4BpN0ekoSHfdKMW1gF5qcPzuo+D1g6SJuYb2gAA/tJECwSegpjIK0
7qYPOFw3Lyp06gpTzYa1bvzNkwNuTjEn3NOShPU2mqGG4jHkCub2nWTJfwOSTgR9
iefK7I/ItdN2YKaFtxUay5ZS0h06ROMjTEZ+b54qkcx5O6LongYiIK3IAsTR/HO9
h+H1QN3JXWEfiDqcgJIuNXFXgtDnp7L1q+v/ntqNsV4q/LLlUD9/R2nN3Nv7TlsW
vB+zd8DwJfR7/zh05SPGghoB9oQjhg/juQMFTqvtdSSA6bBtvA3DvzupAHKt64ak
+RSB2GYkvITPt5+nayQL42cklKy2zQHoP04lEBXg9vWzURKyz7JxRX88tNwKItK3
qvw5kfGBPsRilaJ5eDiKj7UaKtZA7OPdz4Lel4rxxRysEGiDGcNL/IbrEfguLpQf
65MdC4Cxd5qZ6YJu3kCTlEASHiFOsaIc+LlGaYWREvcRs4/pYmbUc2a0FnCh4LG/
ZfdVvfTHABTYnhv5Bt/EeHFG2SIy24MX4T3dnaQLv6ZlmMjaL86tg4gHMNGVR/xs
FQI47lsHrhzC9HeuaLsUA+XIOzxuWkl+rDyvDHg1XY6qH4ACtWDeD7MPmuabZ/FW
51J5Azb+Kpzog3hh10avloyspExrOHD8vo2+YnLeRdjXbGG83LmYEYBN9i5gwjMA
WOtXzl5qvMhKQWX3Yc+I157T3pBEXt7/0Q4VCmnhVXgS8xvvrWPkg9oZnTogeMDg
aOD0HedZA6TG6AAmv3WWFf//ms/m0aRG9WoR2lWccB5xjF/nu+bYjujq4BdT0/Vt
nPSRwqSVHk1BP/wrAQjxkNv6JH1w965RjSMf3zcOVsBSPZ8p+l1PYt5rp9b/RDiN
LNoCiUGNQjRDvESfbOY90kXw3/AuyCUVmC6D0Zek5oZLl8vrsZ8MJuX6OyBBjOfZ
BHdBU9xgbYZiQ87yVXpya8NVx2QIj2wnt2H/+uw/oKRS5170Ar6WS8P37R0iuZuf
uFGdYpC2cSIwVUrAMaG50bvBdog1iLWbnroyShpM+m97zRTbImxRAQlLaNE3yucP
5QXT6BWwALPh2z0AEb+Gklz9TGOFtZz1za96LfzMGybi3gNAOApucNjsXqL+ZETz
TNR09DmUOr5dhbnwllDIPXrrDQSwNlXeP8aTeF0y4e4pnyycMmkz2HhZUWDKb4PI
rLr/hV/9J8XJXHKYmE4X5wXShnnYGVWCkmBitRJ7XeIqByOS/j+/pySE/4T9P2jT
htAVZ6Gzq3rbrJhJaMfC3semi1ow/LuHjRYQroFhL9nRHitlhQNPK/6QFzK5rObc
AzSDPZl2YUJKdu4o1FUPRo7dfKAEEcvH2QoqZMmlxl7yotmJhB1Oi28qBQZtpKFM
PujOfzOs9LrldgLq52jDfsndWPIAzR8Uyk8GIvg+pJkhDSwbBtKfc3Dsd1DZrwdf
LijDqyIyXo3t7d8bRfWOtnyc+xWsev0Cpjm+uD2+qNLPNv0RUTGH1nfVIhgFTyux
P+rZTqrMSo3bF4OXJ6nTo438SI60HCntIcdQLtrwWOeUpxD19cObV1/JzVHLZDOl
Zh+LCfLHWGqKiIb1869sLb4s3kxyB6OCy1awVqh9nQfhq/P81KYOpDntGPkdSDB2
3kiIlk9XsYrQpNSx2QkPLXJ5L94JAWqRER3qHXNuR2VTU+G/6WNf1P6uqznxukB9
cmjfGy4mG+Nc1QiSDuonxaDwdFRWL4WsPggGK+OnSIR+mL+jKzuVhobDGjprhvvy
vEjQV2GcU26VSr9zhxs1kG83mHctYuPeeR1CZlWdm1i8y/GIySJGDs4m6txaGYzr
7zLayJbJqfB4skWPIa3R30HBm+FkBmSLSzR4HTLSMR04vHttpag/m/9mZwQCVyJw
MAVGksV/p1Rqfq3kcQLIdoCusShEyigSZhCyJBm1R6juWgscKJhxVJFtY+XP05JE
GFszLVyNRZHpITx7v08SzQE6Uu/K77ZcNuMDplgDMokQvNx+AgccDEs2BCApoYL0
TNJFoGlebg7TZlSZJ3GvptVm1C0XXpp4Sk+V3sJ1vX9YFlal+PbccmFOIIKzouXm
+4u9CTsK3kpNkpaw/eTRmiKsMCMxo0vHyQqYQlSCA3joIjUXizR9SqoUfLCgUrCg
sRBwvusehO1JIJ+61RkZPnP73O9RYIt0SsA2m6NBCG4/hS8vX7e6QMxK1h8BFVol
OLp11wgXApzeUUMkVdxcVw1rXL9evk9rVDdS/BkA+OHHn9sWGLbkWSSk7jIVOaK6
1GDpeV7ZhrB0ntqf7hpSpf29hJ+d9gaxt/gI5c1QekWLuKUd6WBn6TO7Gssqq9Mx
Vr0hcD7XvaYkfx9NM97q4OUZdX7/UmAJEo4rJ6N2HGoSbnx47BDNXpSy2+T7Ovxz
jug3Fuxt9/Zx26dpVe1DMBfQRw6wxfEuQTnjdFlnFWdx/Pjdfu1ZAOhWNLVgLkrP
i/0foECk5r6mpoJ2JBat8OQvhg403OHoLYVNh6mXbkYuenXfcWkuBvZOxBcT417N
oCPZq4czBjPeYdwamSuUmbgJybWDM+HMne/r+5Ye5WEco8sCi+YydhvoeafoSn8a
JOvXxjaUrRd12B+9E63M46GSnd1MY1uJqcdcN4z6vJiYKt9Ce9lPa3ELxVPBZ0ix
+8FqXyQvRf47TIsS9tsvkaTsuYl3vsokACDbzRxVNX/HY5OXSwsOmD+uw0MwJHYA
169DXJ7VvIs1V456pHZ0t7p5yCFBC1dg+R0bjbl/tRymOshcQdKHTCuloCc1Nba0
V1yReHIHNDJEXlkKbOAIu+vtAZDu2Gw7qZytswPhgJ1y+x5l4+i+eEwycXtUm59Y
s6eWNI9xeibycJRdeuftni4GX/wST9GLZI6u7LihmTXu5f1rsrKpI23NQeFT6MAi
+Ypla1eeXVs9JMkBcVQx0wUxxhKXGSnfpIB7/+icPVoOFsduRc3lyR75pu+YVfm8
vwHcQUHo93VX6X0nY8pWeLxn3xgtzfu5TPkUkErD7ML9nXLujHdRzUiQzdKLrLrJ
0BaYn+AkTBsBAqJOjEnoPNgiim8X1Uj04idnNmMAOfjCq7gS5mWv0AvKUYmkmkjB
S+zZvgpFQBPEj4h3hMXTBiNBpen2ceiqFyPxmu3+NhUQ7xbd+T5+rreLygu+/FL/
8WlEYEB9F0S/XYwbT/n77hUAWutW/L2rnu21Gc4wZmUqK/YzS7gUoyX0pvkpiCih
GX4+fw5hIt0vzc1O5Fi/akQQoCJlia1GN/lR49FkKyZXHwfEZMdz+yfu2w74JuBa
d+54sNsEMDuTZ3pi5s+BNTdrpi6jzjD+HrNkittCa/sLWyyFpaOhayGiK/sWmOym
IKUtS8u1FWvOwGEB3LY9wGPDYlKBvwQNz6golxISEn+eP5l8ur5tdj9bjO5kxWWc
WhAMSoLn48WBUMKtbeZZ0u5E8zGspaZbZqKyJ/I+kIgKIKKnoh4iqHONPLtn0Y19
S/dR7FGM8OKVnJWZwrSw3igFONuoyBS/NA+AsEf+BBs67eSf5DdxFKkfacdAATL1
NeahQuQyB7B1ezW1GnW64oQMb7+KPgrJYYtXTAhzMoEEil78Ue4OFBtvCkUH0/KE
c8y3/qYI7I9Hy+uRvfPUeAFBae2KskNnRbGVjNPgbYo5gOBsA9P6i4dL/YfE7oPt
172+NT03ekswdW+n3pSZ09ZaU6QPR/DG5t5OfoqeRXwaC08ZXGgGOtMTetNaipru
KEqw4xgdB7oDT+BEe37GiRHCSqk8lMZ5cGqfNvNq80S3VQdP23FhDd7iSclzYfD/
8moDj/M65BWaoeNvcZzgWylMkqcq1zexvp5+zrn3NGbFG0+ydSQGmhytq/lDn/sl
C721Fs6qm1ue1OCi3yBPgoScZsqss07oobP9H0ew34zZY+nSYN6c/qKf/O6uuTyg
qO/WLjd9f75wdB5mdisrF0BNkIdwTya9VIWEF31WB1S+7aW+TagBtw2xCEwV1Oji
r6ACY9sPOHKXDxhCbq75t7VZvG22Oy8cK4vRbxB+WSnxnA/8f/cgfA5sipZMNa9o
E7bCySQlega7OuzXrU3jTxlWOW1aHqQ/B1EnF+BwqOTg0GAa4HMoGKEeoqOEbdg0
akaNMn6PoTte3/2LSpwP+oTAudB3BWxHRDPiDBDDVs2QNnOsoM5Szdb1E8nC9hAZ
hPhvXrPhUv1OtSUGPzLjol6XPfaw/f7yk/HXU69Ps5bHi8pvHDdRdAmbeIJ3/K+X
sksKCz4l6pWJoubexwgg7JaJtN34SH4gTZs0Vzq6UPwoJ81nFmwTWUyam/FxPUWM
McwbYkhb1k0krMOxdqnS1b/WW4TzaaMMawKUYSuAOdsekrnnTfUB9bKkM+v3zr7/
9w54a9+gJ7+XsESjAfaM41jswRFLjMdIx6XTR7Wts3BZebMJa6XjNhSrvZkJuJqB
9apj5uehsnYi4zjbbwmgewv4fqyG/YTNIGOZlYZ1UZP3J1AmJcUQeL0viYii+Ndq
RtsDGQJzblZRtpzp4s0SWILmPj4ywMgLgWoAx7m8rA8Tm76FAGJmp0yWnZBECMO7
PTqV8cskuBgjTVlemZkj/GVetPxqcFaSOlfhGjL88FL8wDHKtSnnZlZKgnGu8vfp
dUj1ZU3kcbxHlf5obHVNt2YkUWQfi7uRP/qlcCr96L0KvGxA40wCiaxjCyrFhRNg
Zw7fcnEQqPBjv63CUs8hFxKIuWvhH9BLX2r0eQIYklU+PF7y5ozC6z0qwUQiR87q
8TUO2DEfu0BUBxvDHkdr4IzE1UXaPieGv9h0JYPIMMAYi8wSUmN5Vd7Lvg0Dq6Hs
a9LKdSo9WRfZW0YNV0fmtD+hhz8xWVdQLp2lJ+Mc2p59sL+30NGwOHDq6TahU3lk
LQ60PItgqFgWk9zV01DJNQ563MgWWRcMLehSKIFaZX2A60xhiXonshcjzYLz7uYO
nsCG1ki5QJJu0ouFpZkjYweQ042hSL6rxf96dL7ZLfx39fTnNi/wqxz8eis84L9i
896DtMLqqYv39cmp+zpLTbQSqJmtKqwUJZiw6VFMYFqShOzLxVpdKF16O6rig81u
0TMmOzCZIAKcPA8xGmaap8JyDeauQtHXqkVWlxgADSRyzTQb8KQNZCVMoe0sYuvn
EU0SB8FYUyrDr9hJNkBWxoFGK30yTwinplXUMP9YFVtxPvVTnC7Z64a3VeXuZR+z
FlSlQ2TnNpPERAuIvY4S9EjMRz7FfPLDJzTXtTz/9G/QBZPf2nlGf+CHc77orzEm
/W4BehmQG6cHrxzCmUWB/cvJZKkC+ckx8YKsuA73Bty97DdgLsW9xmhil36DX9Fh
m8FIUrz0trP9EnQ5TD6572yWBVDVNMmYg9yDz92yNHfcpcn/0VF+pxGfx0NsPUxO
XHayIb51UILrANcNb3MW42diDBUcW2q6DkY/7aLFMx9mEI6K7/n1MxG53bwMHn2I
iL/CQZZgRSV0j2485PMJmEtAgbK8x8LQ8OZ5utjBariSAQB2bP8/YZEESHnuCiKi
YxZ36i7E6ZV5ZwEFPrI7smp4CuumFVKeB0Kx4iDKqTGwGkfgmcQpBAFACM6FKjHH
GdWy9JhS2sLYpeUqTY+ONHVy72ViTCaXE8Te8rv2Uq2HD35MwW7fJmCO1lC7efn4
o2CNg6YjGC3alhOwPfqp6ZVyZoO09Qe35rYrjpuOFcpeUQnflhG5fZzfVL2XrTYc
Yj1y5xcqZGjszhw0bXF+VX5XFQREpDnpYv1QN+BTTJ2yfEs/2nNEdzyOXKG8mSQ8
V/veyPROFCWwlicYWjK7wopbytcFi7TD9dEdMwdw3nv20z9Vz8Uzx0X1S33cZS7U
tdcAuNyy6uqxGE+10ZeTQ+iwZOJ7UV5mumhAjebtia2/jv/cMpVkNW6MvyoUHJb/
kmG0pDpiR/JRNqVr31WfihamDfwL/2weUQCS5m3qrhOuCOqil0dZ+BI0tWkQISOU
Fqq4QD9Qb9DojdRzALfIfX/f6KEBgZrGPFyRz7Weeau6LgnALlS2sNkRUmBcmYZv
NslXOSoTkAP9A7csgWU1FPaWDrFDX/UMFdgEzd256+fFtfDWf/fv4giC1MonYvrK
m2tLhypQlL3BB0iNkGhvmqfxOjjfrtNSvXS0pk555EcSNCsh/l2cscm8DcHqzrVF
vdWS/VSjYkI1jPDr3VTYLwiRnfzogPQQBaFrPA9aWHiXu/e8U/mEqmfTKQmLexXy
IE2RTvqtbnXXbL8gSLQc9UyyGZiuztmKKX4cRMnjxhz7VkCJ80S0Hbcz7jS4cJdK
ylW/PbPgqqYOUuRw6beNhsuGcbYhmOj+Wei5BS9iMJIur/BAwRaA+c6nX43qBM1z
BS4ZMe78CCCatxeUi8L12sD3NzuzwaOv0S+iMYJdlq66tOvDA4pvF3QCgf08eFdb
j/K5BhAHoE6bZA+vzQKmkeZxFUeHFrSQZR+7Wy1JwlFWEuX76ecvhO8wAePoqCWz
qay5QW44QXgf4YGwSuIQ7z3xi6Qx50mtEgnjUV2SMX2fL6nTtoDfyTxwSkUHAHXC
bgCEdLnCat7JFfRdiiPIOG+b4wec6krIGupknfrZPjQZxhtV+uP+nqxDLfbxs0GO
q6MH2uHPqqNjewghUuNX1gtlcPs8m1RtKXPCgV80VeLAViKxea84mIy8fmbyjg/f
ymUKnkX4itcwgnDEXgDM3Kbjw9LTC6BNo7PHTnGGj3Bt7K9iMHutLBjz4DzZgGHn
5J7njHT3d+qzsX8ByPDq+b9aHqPtq2xtG7LTyMdZTGvB7lC5yvzJx53uBH+5hebS
u/il4jSmANDZMI9d7OEdI/Ynu6r0BCiZHhMd1h660Qt1lUb2jYey+VI95uK1O1oI
1/Ix1fF7CHGpkYLOe7ElQOvPuwE1JTWo8S9OnrEUTYDCF9FcGTlTNznm2vBzFFPo
8aDzyUWoRH7cl2tKm3yhpJpxXc/Ur4buRcXU9v2BJx/AL0OPeRMqUizo6O74kQVf
B0grsI4GimjbMzeS2JIZsY4Sf387gYIm31x7yqraiFJfQXpXEnBCXFBCv7kFVq8m
1MeT/JqhDfnP+c6qGpwDGdBWNg2DmEarHerbxCH26HopPChQEZXNYuEIXaRzVDEA
rnYSaTqhCPin3Khd5Ccx3YBp/5iF2DFmSJoxnG3gpeZKKL41Y5IduvrnOyv/+qTg
IaznYEdHT67eLPHTaUviKF4dIG0ffPByzSOD6L36WR0rWBF7PUY9AYqOMO82jCbd
e9Mhff/eRFRyrdFx53pAuHKBlyHr7jnpdh1HvOtNxEOnvwbhxhXLTVrXmrx4kv8Y
dwZ95H8XE5cyR1fGm8rfhyVvpLqaWNLF/dv14XFQutGXRRkyBu1MYuGxeBIAful6
JtR5zk6a8MHhvu9A5ss45Wy/wHoYsHdvB7BIbnjL8Orr6kuk6Jddz1lZ8H4J6phW
tVOVJNvPhKYskogW8I4gjW3WqJj1lyziw+a4gAoFOgzWutQRnvoTQg85Rd1kT+P7
703yOoRtpqNyFJcf7M3LYJc14h0Z1D8MyBIzCZbkzyz3DCozc+JTmxIEgll5yG5/
0pRXAcdneFLojrC7Sd2oyQyM9GZJqm/N/Bv3Q1LsXNP0ewl0ExTs47MG9gzsizah
wM8t2l5wwNFb+AKIEFrCJSfEjgV6YHW+VHOss608a+5nur4jDjLK9kku7o3ToMN8
O8g57+s1RNKg5oAscFpq0KwgVKl26v/CeBlSHoeLVCwuWnN+xXsA5EWSSbhGb0Qt
c2k9kjzo5vfukz46NvR0H1qUjixaKgrwrtQ9ehOeKyQ59Ctzbci+EIiTw+ZU0Fl2
HfFuVd0hpWnCnUovM8GGGTWkC8ikDgI2Qv3x/gjthq7nVuuyVtWCCbSGfsn15Ylc
tvo232pqByiI9yofJbj3uau0f1zWo9pgaylaTYX9Gl/0AbKS6L5CuFVeFv26OkGn
mbM0IiYV7IAh+oCx/0ZXo71hIdl814VGHX/y1a60Px8x1wPOsfUEM5DqOGoLBhIr
JOau0Ed+gW3YzzKIXgqN6Epx8wbH64ZDRF6pckn7uOIiOCbBVgYXO6mY5dQpFfyf
BDkhj1HbOo2fybnAQbwSOck4+ZMvTGdKfb2hd3TuZi0rSRpGlE7FH0q8qLYa9qPm
a+WIyOy0Rc4F4qPojVXs7yv9kAo3fFXze2cHKZkgteMdyszTGTZrg+ktj74q8OOQ
f+zxn6vHv3PMS7vIvrO9PLofRTygVwqLvXPaxHRXhE+aJIk0SsvYCBoz+txMTd39
B5g56F5lFIITjNzy07iupDsDVq3CmqSMN3GT5fc5i9PzavbQNqhji92VDWno7dZ7
FozSfFx2wbyHDZhrp0vS4NxbE+1lzECgy+ic+Ap9Lh5TgQWR5n9R6rJbAI1yJDUb
A9IFk53dPXWE9WIOG0JMYYvLR9H9wO9VdCmMa2N0w2sGhI8Y6/mvXe53guRUHsxH
RYaIHlFVFrEo7o2b5n92g5u8JgiDTBAPgdCUdfwj8aF8cyziFMrdDtZEGsuein/l
oD1mHD55UTT2+f+qziWAzl1i+9XjGCR0UZ0KmB7jefkiXmXlI95Qpb5MoGt5Mbpa
+8yKQsyQy8bgaOq4dqZTzHJDZcnAA1GDsB7d5b4vs4xXuD3/nYyaRzmlDD26uyBb
xfmICiD73/T3RVNA1CatokActId5YEvd7vG7LgoWpI3ujea1jPlfqKZwwF2du7OI
Ya+On8ndftKYmeQuRaT3FArv5jG6JZJFE8NLl1VxUFLOKXsNNFy5n/l2xHkah/8/
9YI3wk59MB/jqAbzWqmohm0KSwGd39MazwIXifzVtpyss4pWfrt067D0RXVLqsLC
Kxq/GdYk9MfNvMQJHjF4ANKDLNkNAJnYe0emNUS/hgtP4JBFlgwBDJT6rmHefZf7
9OPpwIqJ+v/L0/1Ip0PUMYRGRj+HOay2yNzy2lQqmXh+mrLnXnbLjATvS62fUQ3/
6ZnE8SELGnNGMENN7nQeWtuRIc3B+KFEArrZBDlqSBtRogu8GnjYSpoVN4tZVKFa
kXBKFL9aUBB01e4czyB/lQaoUpXQKidc6AD/hz0t9DzgWSUbW6Cq/7rOXE5nz1Fd
6JfvrBnp+ow4X476rz4G0cX1G1GtYfx6ZlP9vScvY0fKOdHM8eKyXIM5ZWBxmQ7a
ap/NBcTDgcZTjeBH03DHhfCcHQltIN0T9XsNELNQeL1YPaMNIV0tABhD3PHt7xJx
eaTHEys7UtrQSXVdGz7359R5izqHJ/yB0D5w7AnFANd2LAIrVaHh/Q/+CkkwqvjK
pezGDwpeMESLLAJSjT0ocn/zBpGTuu5Rac87PX921JIFUo8iAudgEnUdmsEwMRS4
HadEQ2OrSmahf8iSBRNkafsFlWwGHY9to5bm676sB3Jt96VGEGQyoVLIgNID1OA4
Xjtu7cFRfJ7d3NKGdgBzyZ8drJ/qASidDmNZ1FPsejId3qt4B+tUTb6S6iMoAMBp
xKNQ+vtlsSg+18uporKRD8HhavhScQMyWS+gPsA4oQ6EBPQ+jX38ZCU4fMfp3otl
iWtNevPq38wULUyEa8kMXXo8TmCGwH8HGl7n9UFkgVejU7Dstm0/49PUjDAw8FPg
/MvDxMsuUVSdYo/aw2UGckBZ6tSsH7crG89el2N6RIhaNu9cL2/kBh5BEzbe6NGi
NM3u7GpHeEBpob+t/1suyjlllKgethWr+6KX2RKufj1Al+ebRINWMmDTk7SHXxxf
1JXYVge7g6wZx7W64vCgCADwUopDJixzJFFCJVTL2N038v0gB5IUSATnncV7cx/e
WSCfM/esojbXfxsl/rbzWajoq1URLfDijF6ekfuzfLPkg0IKdvw85CCRtwGW44ta
66RrmU4wnK53geoEBWW/y6Fv7HkU6LRhwnulpCnNDVBkgPgcPP18IcyBY8l8MZzB
dSDl1iPzDy0f/hXlhl9vKyIKBgaERwvSNMwx6NTlgtr3hvboNPDA0qS2mee2ez1G
fxlMtDFwkT/tDy9v4ACJ88tprmL86nY6mdzUbDI1YfMt+50vyBvgE09fuo8Ed/h9
0zSln2iN8VjX/Q0iRSIlDn4OK6foKS3Afwq+Pt6Ui2E6eFbBFWr5rBeAa2OD282J
0+NZfbDSs63A+Ma21CaAZs1tO/B0Y1C/GFLnK0Fm2KyxaJe3b4WyC0VFy3rjmynR
31y8SEdUq5VhpN5Nn5Ob/8Glfyc9RQyFdWm+3/7vv3QDkX3FreXgoNEP5JtBCmgc
x5m6ZDWvaLl6IN7B7X//CO7XVZgo5CTrIo1Sr6EvTSTpoODuvMFaffjIkSQpbqA4
JckqPtjfKC4Vz0u2VsEZJpLAKh0j3lPEgL6v1dWfFrl+03hh9BovMJq5csWIPSqb
usJspQzlFEdJZLAeKBsnJzo5oig5JhKNjh8fOfy992wCZT5gKKNpIoue0+oekKgP
ebwlYNvIAMCW7sZThGVeYnvLamJDN886/arz3LUacny26GAirDvKqiYc22w3EMg/
v1bWqPhb2fMWx9Fqdu8VYGwCLhu1+AvzT6qzQKvI6YKBcZ4m5Gl+4/64pEDJ1ur7
5qiCfeuo5NXBXFwvimJofJUxrCC0nbQXvj6DtwlDVp1gq5JXHigq3kJSAsACavZ9
Do63PCvrGUGRNMNYJKopyr5WebP4E3eK4e8S80Q645ShiibHZHUvlj4u09PR17X0
DZfn5Cn4qqsQYg8lF2TJDZKfNslL/oWJTrkaZ/qxTADP1pLn24530nkq0R3I6IEF
5xPiMvEoEGGwx6CLsktMFrRRreaFmcU5PxymbxoH2YIJKz9fNhBicuYY9ViEpwgK
ozlkKFW4slyz0g6B11J7Lnu7y5YE7NA8Z5HAaM4OOY3k0QjCjHDWllMc+SnW1pBB
XWcC4cmfLrrjPuJz5rdjs0hxTPMFaC03AV321Vr+yMzkvOGrn7Ug4a2lg5/kFFyM
Aa8xQSwgV62LUK+3fWI7p9Juw2yA4xQwkK5qBlRH9jtomApBRC6wIymVZ2XIRgCk
b3dWfes28VONCE9hWEvE2exH8oaOBozGRTLf+9PoUneS00r9/980UJ0UhLqOCtkY
IrpUODr1ysOZ2EHeK5YFBReDaleWIt298ovtI7ZCmImR+JVl3AYVG9gELmEpa5tD
u5hjt4uN42gx7NyMFpR8yo56bexg1hXEVpKtrf6Yp4mUgBOZOzFdW7T5NKr1bmzo
HoZeEAgs9ZKAp45Sjrnt3QAGLmdn7cHCdvB2AX8qTZyGjagSsnuciR8k2G05l14Z
lbfyJF0pXtv9o5Gq5+NhpNokfbuGNvAg35hEmuFyn6Bk/w/9ehlXH7s12TSDRDsu
KL75fBfA6W24bJdH+v5+SUKONjNyQM34JGLw/p4rJ10ktAQ4GdbdyK04HdtBU5w6
zcIyoJCuuR2Cf4ckx5Shy294GkviTv/zuEgF9a0/QMD2DCzOpAs4+B/42QNwemjo
jRrvccMxElLv6kxKDvWWcUhR+k79qYlh1jzbw/hpJBnpSGRTlZO+eo1gRcKSq2f7
aU+FriEljxDhdrrUxqNb/kbu8HDBh5tMNTOXxdeumwnUZmsidag2hwDe0Bd0SITt
A6Z+6uL5rKkNhya1SruNKzAJiF8EI7WA6LTAZ5cORfnuMmKE9fTOtpxKOh1jI2MV
2IRVSGfc/p48rGYwK/ayIcgLxkUoSO9hNbFy7dyebyD13tX3hYnuybkl22gpeiy9
8Pi+Nl90JD5lqv/plgVLocTrnPqG/uRLd6hbY7gKBVKRNSjQvFCt3UYjTTnaySRG
e0cODHPcmEV8WEy6PWdF9cPhTbk/tEfw1wR/U5VrFEJTLcvJJpwJzxFHqul+LWLS
8xojTtoTFVpCbxTra3TXGM1aB9ebDHVq1+rHMwtKUqHl+mkTg/FBmdD/Kw5RcfWy
zs8hypPAN3KCQPXKUempFa2OJpJB5w8HONb8k/bjy1NlQkmAJMfcDb1ckNUpZtjs
QskLSBUgRPxiyN4NHkjxuBs2/IEMdvzhfBolnqwcFMNraa+jZRx2jzMu552JvQX4
JHkXlzHMLkmkuFloo0EFW2KuscXpbbalj0QLm1yZkHgYT5+Wpa4uK74CbD8Ru6SX
I9t5C7V1B5M0Fzl7OOXN183yZcN5/XqMxA21a1rMPqr0XdRx49Ej3VPgrfcag4nM
h4WF/E0yAda5c8xix+DKOM4vuF4qElo67s+Uzi8Ce0GUFp7m3db/cr0GEa/TQ4ez
aJMkijF/1yomrOalZFDkjaZmFVZvb0baXHF8e3ofZt8BIp5ZKYHIy15w5g36qGfl
rseD6TEKB3e79N2nXr+sMV6z4qnhGbXJ8VEYPlf5Y5P06ViC8B9bqg9XLTNJKmch
SScrGi6jlOTYPVHlT7uY4ED21AExQTQHhbgbRDfOCXG0LKRZBA+LNSj6pKtSvYKE
Vh/9QnVzzk0eZspkTlFT1KawCbCCy3ZLIuVaqi9/w2fdriR0vRlBjmFtDRnZbjP/
lOjd9LrJMw0Vd8QBKX88pKnuHOWFRunv9mQ+WUwGdBaAVJx5h7hjMQy52TSgunFZ
YfFY48T8ZNCbqG08iH5eS75ztyJAzHIQuzb8OIcjg3KLfg2S7hZKLsvlxez+Ddld
HIX9TQxUIbefDMcQhkgLHZm9GsvKmK/mdaRRKPF1fJH/V3PGkk64J1KInhjQNs2w
gVUamoTOeP6sYODDmZuwtk0L9HVw5jcJrJZzLal3JCqJ20IUizRT7C1j5TeCe3Pb
AChBBaVVD1pAdopjUPhXhJlVetrRD0yvbIJzAmjAAnaVAzaUw1cshXi7BKFPpRTB
gV/yhjoJGaPIzRjVbcZF+KhKxiwYt1T6nm2e5mfLkB1gVMWYkTcV6KciKg8n/eAO
NdcaAyDVthAHhO5/sqlz+Swo38PMAxyDgrrDmsAYfpXTVQ+hpPmsi+JXlLpzNtxY
jnXm1eUHLtdHosOB/d5dRHv5E1NkOIuyHcw7WmfKY/jUE/m5XE+4Pzs+adfezGyp
IafNwJ79WjavRpXKpkLYqnsRkI/SmifjZUxHwjJb+ZNxtpSMhQOoN9zemzZFD/BU
9ybkwx+jN6Gt9QTuRE766INocqEGjYvVv504SykIE3Y0rNd6MhqETVHbVbVhebgW
ROAZavfjqcKLG++Grhy0b18nD3BEJhA+QHa4dXq4O67pMdX9UGW2huJ5mOB+OBf/
qam9WvvejI8FfhJNYu2KJnCp+37d5fmprpbMV1CtFQFworPpCvhMkSlRmcHcwhWT
DgHGK+oHwUI1O82Syje68nrVQ4Da0KsoPcOqx7kGRn6XLACbljLhAXUq+/8jSAVp
xK6xAEB7DUCOfYmJRfT1XJ960TbXpSVORsnY8nHg6oHcLSx2+x/teSTW7mfjhJtg
8yaVVy6UKqI1fexGQkQcnzV+bDWcZbA7KHBwa46/23S+shpCybIUxDiaXaf6LYWS
SKWL5LBMs5S3r8WaLpwmqEgDSUST+uIZSWJ87SuAJnXQBwCHwEgU19wAOg1tpbSj
Stqoz4gF7HL8+fKOp+rfSopfyUCd/9uiSowc4xINBKTE7clC/1ydBzlt9HqOiefB
C/qvwwtNoVqXoBojFUldWo4Lzx7ePFQn9kucTTtcVfxVeGI7xKZlBTKPYZFHS1kq
wpisMsHp6b1aqICCwb35VtouzyLUSN13hfOQbnSpf5RpSrLYJ1BbrrIyjtdvWIfZ
zD7RPuxwn4r0TIXk4uo2EyGQnV5hxqw/NoCwkVP6lyEKs3KIr9TpZJnRZZpj2o/O
Ue3S5ARQiIXm6JjqUpIuELtdWW59eZL/5RmBYqb1bmq3yW3IdyqDEW4wnDMDruP5
IkZUYESS2zy+u9oYmGGChRAQa4h/pxZin7TJiJ+GNq6aVeCCEp5xyCc/afMnzBqk
7GPmW1p7U3QH3mpCH+UUsBWHlpq6aLaTNjtKaDajW2hMTMJWL0JKIdN+ZOcIclPk
Xy3L6WALnEtI3vQ3v6ZpiIYykcDCmyIL3e8XZM5Wp3mqHu7ORnXsIgVT3YAuJkzv
aHZgnNbBgZP8F5xozfW/pQwci5BBkOhPbfLg/Bsfg6V7a7AdgCMb6sm9QuKfa+UY
FWPi1HUPbA2nw4taoMpk6i8TdoECK6vGwo5QzcDGBcQrv5cfzdhKYXFnahWr5khF
SY99ahNQLxZfOybR6UDg2CyoG7nNiikrHRJn3cnCRUg2TWP934oN13TkplIWWfEX
UOrWiEfpa+OXyCxzFQ8Cd9FBkFZjuI/B+ct1Gd8+8FCPhmbo8pEmG8wnvnAVNUkE
bY5W288saaXX6ANkogcH2fP4QWedFJIt7HRP0wNGK4fthF/8Ktc5gBl5ySXMPnxC
/ONYAKGRubzthhLl8o8Z2IWHrRTiCkvwUblJ9tze40UHhiF6fTqcXLg4eMOS1VM2
tIlV7g0PwQqkQK7F7pJSuloXBStSQGQQO/PrOq4erInOUvuazpbkTsdHGk90FJGC
Wrelhj4bEDCh4wK5pQwQsEaDPNg+BonNC4dNpR1gaetL+sIyusz6HfBd/8YXylX+
ljPv08boWWE8VWz5S3rhCr2dFL/91mXX0r7NkcqMyy89xJmkuxdilUzasAWxQmdD
kvck4cQFDDgjB6PuRJmzxNOR02TQLx/kOM4PSnp6aM9bX00kyU0DaQ8cbBuL01rU
A6/99ZadX0j5gKJ8KlfbnTLivJg9KqUOqxM026IqSeoj2ZbUQEy6vfcCCy0tKjnf
XmmEVl8nEq9Qp30UDlBv4gMRAWPbOy07uJhdxTmJGuEFFKQ2fxeYmTNDsZNKXYZz
WXIoZjWS0DDZnMxoNN+52tkutOtLhM/O9LzkXUbjUZqUY36Fc+B02DDCefWcK8xa
XqsLIR+W3l3EbR/pNihVWklxyZBTWdW6ElsHcCF1H2QdvkxD1JAKnnR8VTfaZUge
AO+MZK3hSKayGxov1Unuy9BPXsnlPHatOIRgiG5LjoLgFH3ieis/fjp9qQlEa1nQ
LvTWjtvQFaLj6JD+ruGZiBJIlv1gFIbSrmbtsi9brJ9hwXdHzYbQ/Tn2a5yYfi+4
lwJIU0GKHZ0Ixn+iKKwP5vcuVZVu5Udnz96sn5qKpu0Uw8MtX/R17AyX9bYOzBoA
OWBSG9dlY2KTvPJf4laf08/hrpb6uK+xMzewip8WiQBvUNq4O+H8nFrTANfDvSbG
GyEvxZY/mJENW7rWckQyyQZaVkxp2ixNGnrABa98fFah/lzt/mxif7at2R8RaEUc
9gLSGyLZ0rUVyRSSfxYPT3tKskCGXdiqBa683uGUfC5ng4d0qE3j1gRQbNcLryrz
GhUXornemEEl+hafoSsinSCanLzwZLO9fEMvPbynjGWm9lgo8CFcN80sWMiIcPaZ
M+DLpa/q9giRTvzhmNp95cqUkcCsrPLKSP30gCZFQv5QhDslfzS4P3PU3+sn4s6w
2yP/G6XbA5HnBXqAymvQ2KsRVsXvbqfQtkaZxO/nkpLF2LKkHeNbbmLjN1AqklOa
3Mb1nwsSyG6SaaBe8aixd+aSvqy3lKdq2jannRR4AH7Zg9Yp8MvuhnauduLw97jl
Vc6ETQqH5p7UYemDwfdi90wqlyyd44HP5ppDh+/FzduDZFnXyv9xsXIpQXigMZHi
SdFk9qVRheGGl+S024qQizTx1slgJ/HVbbeq07PFnHG57redBueXwU8wb24ERIsW
BVuLAGytEBJRNYx6ynq7npwXDHPL8Jg9K9979ucWlwcdPrPu3MxmvpdEgTsaPGio
RkOGXDb22KvD4y7cGwTIHfWPUVhaBbQkBT0nBFRM5xeW7HLHSSaM8RzPy/HO7P8H
nTYpbUISkLBne5KFmHpDiT4klUPOoPPP5WFfsdatU5jgrrL/OK/wdMPrikdl7jvJ
12l4+qyBgTacfFqW123ug061WuSMdGbVUCmeFN59urb73/AWL8SPo2pK0PgbsAAt
nVvIn43ZLQcwe/DfrNg+RnKc/8nobGjiQlpibcdoQIzs+yONZxwup4f1y/xxw7FP
iK9cbQYOXa43w8cxyzVHcEAXG3uf8Dw3gfNxmoERKdC0PsdWmL33JXyjrZ1Vh0Gh
AiYd4UrUFvGaarP8FKz2Efa4fvzcYHlqEakzff88J+s53NO4cpu8OiQKP/6Cbh+M
89cmZmUpLEZs3NJ/WFK007ri7fhRZAacXmJYQCdt1OUtzdtLO9ii3TmHTD7rFO9c
D4tfYCW69tMoTxxBkXInev7iokzPxf5TiAFeoLjQ7v0Dore1Bc2J8ECmtg2DvWAe
Vl3DXMaqQv9/1CBjA/b+UU1wMvscqTmBJNtFKIn5D6CA9h+F/vPZxMldhbPtmhoR
Yg9zwoy5t0letT0refSzs4grJuewRUYlMkr2DtG9+EAElZtuUwnjUHAupzOXi4nQ
bVo99UDLMBU67AulJdIscz3fQFSQ+UQugrrpdYXIunZu6txzVuGjAKh++QXrBIKG
JZoYSVk11wlmDaCXRNOBhtLc8oMWThMgsIuf8cnfOJ43iuOBTLBcY3TzyHJ1x68C
4lJWj+NzO3TBMPdr79+7fhOXyzEKOmnXy0YkdEBKTbN8z/fbmLIqH8W2hyi29jh7
zgo4CUY6B8LP3IRU8dCf49GmaPTgDJarGsZ6SuO//tIE5sCQDmNut35+VOH+x1+u
0O5fApdgzBq/FGmHo0xXvUQ5g5HrhuJQAHgcw7KSTC7K0OE8dhoGTqPEvFKsrzUq
XPx7WtM7JZCuuWUZrpZlc1uek6xaEC7YpdSze/qH6sFMxVM5B28gvX887q5sG/cW
GcdKJhLiF9vqP1AvfMx6bcRFd7Rj3BnrDVPUaBVTcYLWEo4n00P7sXlLuGFUiO47
5pQ7S5fnYEyTU06HvJx3nY/SNuOPmriUmmvq+H6Zdx2Nvgs51bThgLsyejyR7j7N
6kvz5c/ajee8Il9OtQ6G9nJQgvkG/He04QTRcMulPPHM0J6cte/776kLTTP+qQL7
dGM1955gp6HDl1HRtvyjcJH/xMY85ZS2JbeHF5dwz7pnzN32FypQ0TNsToaxJ/19
ypQuJC08+c/xeTCJUaamwLuLuvPmozH5O/SIcFdl2wqRS4Pbn5CHRdYptCVtQn5P
AM/kdAnlN5cV2ntCAqhVpRZxYhIEqmH00bYC8p2rGigsPN7g4onQIdUOEaYk20Lh
9o7mP+0g8x/1wLTmb6QRi0CC5VUdDnymHSinbXg1Q8MsLCsEC7WjkPAXc7/x4Xv/
WMCnfHsDod+/90TRdPNGckL9jYLqao9leS5o2OjY76nrkALYFJDhyGxcgkuYgFPm
n1r8WsHVgdNkZwIiR8qcZpVVoFEgVM+GFwvo9x659+yXT2nXRn8xZjWa5RVS5Gsg
r/tTVSTiWbOgROx2BAZviTdLASOMd0TUkAKBgc7e4iFj6AtsD9ZIeXoF/wEwtcCM
1LNS/iA4A4F4qbI/dr+zhkSYqOoDvu3t3kn5S4D+jzK96wWaHsXUypE7OqX1Lxbp
Blhl8PPeOp9h/7SMmWrTMY4+6ogIBhH0VpBoIA3LpA13BRr3yNsfutjmr1VciYkr
89ky2hsIIvs7zGL1KAoDeVJJCHUGHbgMEXVXaLsMVrO5p9O23gnDHvWk+kyNTYTg
WtWXAbHJbO6+UGRm6XvBcSa82BLyD8FfvenqdYZfLJSDa8U59PWe7oav7sa66IGh
Op3IDMOwegH7uyOW9WoFQZrxpU4EweFiq7lB7g4Dg4kRYkXNPP+Cy5wppH23y48T
ERwcwsz1KsmGtoXIiBk37PaDntPXOeeyGky2Shkbj3DaHYWoMduAq0gf6Ia7zMVc
MGIllS7yzxgLi9UJt2fV3cMAfoqbwMJCUMfH3OGzxRtjQ0mkksipjq6EXABLcbhO
d4oRCue33z0678V83GyyUFeldGbc4WQoBLg8f3sYpgBzpiaBoc5hMSvx5Z9pZOdd
gXxM2GhOpOjaEk3K1tq1gkUNbA2n6VuPuZUpt3g6OmzOEovSs0WC8KwL5QBUqpR+
gPGBgwxz1AFaNjoM5CdD3XgtmOIdXh8ZqtOs8SL7rfd0ktr531OW0Nr8SZrD7rgO
3kP6tYm+dwOJjOwxs1oGDYiSNNzO9Lria512fC0O+pG4O+WlYwMiyHeYayYxjnZz
B2yuXjzQJcqKBQn3q1LlEfdyHMaTMPl4qjrS1ug1vZUzaTVaVUnuEcp3fT4F47tS
nNE1RfKcUVAZkrDTbuw2CV6ECnX5ZN3skczOof1BzIAi6P8u/W1rSKceh3tiAiOs
NWNu5DrFigSdPEcriBfz/GVKFc2H1GxF4+UkONaLa5PgI/JgwEZbA0EmgFOQ72vV
jjHZIKJgJWCKiAYEcs+v1LlUgjNBKapSwKWwsxmJughkMuUd/rlPbc/up7tkvKVE
+oC2EzWdIlfEofE+vSlhVVTNZRv99EYisSyY1y4Dvs+FfvFrtfm/s/nUV4rX2f6l
C+1aNMpKYfXQYYQVGIt3D15IS5XtN+LtLxUYiFKU8jxYVbLAgyA3JR/ud12823NH
r9KQ9a7HwpEbKqz1fWlRyCAH0W1nyQE6jXKLE2GLQHuTY+ZtkO/4U2zJ30vF2lif
YftDiTlbXiOVoHSiRybJGVLcT6M8oUcNUench6PtV/qzHUXyctFNluqdi/3J8wPc
7o5HTRgGdodEmccNnG6H3fC5pJtZ1AxNcwCey2SK/B8W1D4AptCdj1a9/8NWJwyh
mP5iIkAQ34pGMDV1dtf4Iu0/OgOgdBzFLAeomddtb7E7545xfy+6te/titidCrGZ
u7VUZ2WIB2pb4aDZWGzq7hQ6Uie+2lrwyc/afiZDGSDGWIHtRQV3MSKjy7rCFQlY
OnjmqdGkkfg7v51SfujgJCXxQaXZTclF608Ek/yZKENMu3AQszU62nUREZg2IxD5
O8zWTVvzrawHzf1bys22eebnPN6mgxgYbTFH0VD/8sUX5x9YnLWPaamZU2JKOkqd
aMNlR93w94kJ5XWH+kOiZ7629ZskFDh8Fu/Gsbt8JVXVkAnbNFzBDDGo9eRXszch
ATHYtj7pLLPxbZMyvD1uop5QVldQf5C6E2BGa7Kg/FBmoTwUQqPs95d3kptabuZD
acqzZ1LQoiRk/h5zAwyXM7X8mZ3I0pC3XCSLuLIPS+S+iP0mQVvctl/EhC9x6/zf
gGd3wSgiau8DQOs9E338JuhmqHJdAi7yAw0Uc5uX83qOCmdH8xviF0z5L2e5tdOk
Xlr8gSkCgvwHBHfgrfabb4HWw0e0xXBcHumTxpVg6aXtxeH9MNMbEx5iGtVfVFYp
Pbfx0t3aleeuSs8DG52HOatdF8rqenY+SeCxda0HKlEOviFBezhEEjpO19U3SgTf
+q619b0hs2/Z2ur/l1t0cZnjezCA17itKbMYWtMXeu52fRcmSwSagiLdwxnu9vUj
nV+CKhnqFzGgQPdYo4oEu19bLBz3jzmvygW67UaASKKh6unSEsGrgRJPqqrDxu3g
ZSDo5qdMznap3zoglr2PgbdTUXhVTMX+5P+SERC3qnmNmA699P+Z4ytML53mS6SZ
/aHchotUJZV4hfWYLnjjnb9GefUuYREFeeskUZUEC7/HRWexO6I07gSi99fa7CfR
r6bzpgyqukUrwYxeVIQfaIIVoQdWyC37g/TiE643jg6wWGLr8BV9D6FwCZJaRzoZ
cHi+RcZDEyCagPIW2jbcq01XjXjXZDLJRXNGskO9QLdv4b3Y5NCXd91pRRDUTff0
wAZTVDqw/64RocOi+BsFFYsOQJmGFIvqzDMFQGfXwQH96E7En83InNB8i84DAvIR
8NCz2bxCK8Va71UXNBGNWhsRrq3+ScqiAHkHYT/wI9h8eJHzitIhM5hmMjJZxO04
wdSWDoutBMJBjlQknCygUPxU96SGR2KggYk57Z4n7mSClBPp+B6m6lfYrJmYlO3X
WhHe9lXJ4g7OsCf+Dm0Hm0aRk1I9XyAX3fEkPskg+BmV7z5sZWfV+RhynDZFwoua
8PBnojS7eLEYZ44skjUb6R8s2iBlVBzdWeOdAOVD7yE7Q3dibvpwOawCEiBW1UAk
cTqoT7zjqB4YO/4Qa+5s0A==
`protect end_protected