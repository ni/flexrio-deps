`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11232 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
DmI0zUXpjr6rtg9EJrlnT8oAkBeuE5Of2s0kai8/hOYkr1jSari2ptFCV9NaK2xW
zVcRZKwSe4xxHoJcuISIBOVv7HVGayLbcZxD87XL5I7pMgj/UTH9wF7AqH4gkDj3
NZRw5fmQfTRRnjRaLzjQdZ+Ix2TcZUFZeHxJ2VRZMPUQnYznq9Fb+ybVUPC5jXdp
VXiQL4xQyK3h04yL/XjUOTLM6HJu/Aj0omXedoUHsKCUzAguOiYQxchPdSuD5MMA
+T7CMEMBin3wfyhiqbSfxaqgEWjmNAcx5E/AzJzbGJ+4C6O+SiNRCgwWAefg0TEJ
JE5MPzG+s8ZWKDh3lE8Ih+Wij6lVK8o4PzDIJzGUBy1uUpZRALnRyY593zpzRu+7
VRGl9GrOcck5vwZVw3fD4D9Mo17dwUzHRyDoMzgkeckhGNRpGJkl0YW+UHV3ivYS
FpBcu6bGZuL1rgj3Zaw8iGIQUXvzHkEk20musawA/KlAjLYb0J3t9J2DPOM5G7xc
uplYfqPuGWjtb8hguuGgZD5u8VqcmuwZjJs9J8pzsyRDnTIlxrBbtNUMbodVoqN/
KPlfqvlKs1X/7yIfIsDgBqfR4C9x2cq5ACrIuvhMEVmadD05Uh1fDV6y3WiHDdiC
Pky0ZHhwoGkGZ8fR5tx7ZMQNHPRe7DKEwNXRMtkN7hPFWC4P/UG3UsQy9yy0+BCa
hFbieWZz/j6KaAxe13naD+Ca08nRRze0ARUNL9DAj5796fqBqwtl6HC+j8yo3Lpy
8d0AfHMYWlMqKi5YW0ORA/sEmzUMYJjLbgfID7FeY0tePMntliYS6tEQWeSaAEll
nod7cDKqCft9f0ZcdJR7Jd8UfV1EjewGeK/w+9+r8grPxNrfoSJdxb+6qHuPrP43
WEQEOxnqzes3JE3BLIBgEoOKIfOPlsAprF4tEoY67XGM7vWGchXQWLJCVSxTyNwf
laiml7N2OcwK7Ibh1XsTbPiMlzRjzYwiguORJzbbAZ5oGJ4ACeJut4bh9hFkgoTC
/2LMzwUIOlEbsRCg7yZdXbLP5piYp4SX4Nz+Cxyc1FXSjWopXL89Rm8o8Wx9i8jS
lh9IAZ9xoYEvfZt5zxuTnSXQtTEUPm6Ie7PZDEGdkW5mCWKFD7wbtn9P5Jqvu4ct
ndJF0G9JrVy8tozekLGbWaAP+GwhVC8x/cEab4aQfRErfdxzae191IpKvTW5aXu4
t6baVmKQcHCOWNnTajDwN1noGzsA6VBQathyY2QTR9nV7ejo0h/aGbrZjb0feuS2
QabIGmPRApmN+9hjoizCVfGvozkAfFJfr3gexqtWoKwawTzn1jc0Ji2xghyLKs4a
OjnsCHU5Coma6J82hwGJrGT3JwUiG2HtBxibsn//5YYjAlqu7a16zoQNPWUKhl4j
8Ovc3eixyuGfbJnNO5aOBV3zPrhIxaxUK2ipoem+hZ3QMO3qzsijr5KANrIbPKyz
tG4lID48TRtwQZGo5UoWzKsEv57oYGaDuAMxUAgqre9ZT1Dk+G4ZiBLHfglzt3jQ
FVENy3vHx5D+yZg0zCmsljVPbKvhuyRBAq94juGa8obfnhuIQiXp+dV+bnV1PqvW
mnpMNqM0Voua2mGXCNr61cZoo/sXIi38fOYwmnq3RjFvh13+NxLSgAdOHN5mMvaR
AzsOu+3AzsS9SlX9nAws9Iu1K4tB5p6mpGn/CajNWA/gyJsK6+BoxLVefe0TnJMI
32mLC1SD40WvVGV4k2PENkTACBPM+fiVmJsDB56lhQUVMtqAKqhK3nZaZzlv8FVA
3Z8DrJFc1xOFZ4XhxD/d8yGkTlF3SyjAqCVn5uAajBp9iqC4B69jz5XkVIRYtPFE
vIo5i9Uz9WSXVFNEKc8u97gULg5bmWGazyBJ+oz9bG6kD3bxdZhzX2yvL9kLlNk6
26NN/FcpBxZWGPSctD97euTP3qhbkg8KQ+hy1f/v8xr59510GWV+D0GbH6zKQ6B4
X3VYEqRIEE69AQLxO0yHqag/FEApaQcpO92VPioHy5HJ6offTme/PlyaoU3Ge7/n
zi8+SrBF7XbDTt4aHAzc+drAWD5bMYoK29lvDI593aXTzRRL0h7+0w9ql9UUQgib
NhY8yx4lgKmO6NrxNRTIG3zAPR4yC5mPbYlNk8suh7JxgHF1yjNgxBM+dckG+WF1
vubzBzEtiul4OBWaJSsQS56gNn3MBzDKeKFMNs+b2w8lhh1v2gTTOwn2eXKEFuyh
m1w2QTdkxZ80knY6r0OWwE3VRhtLkl9el2i+hWALOEis5iU00Z7KavRNKiC+X2Ko
rn4Am2TCfszHPqirvzbdtFO1m35dFHEGbieNlwKHMzbl7mBuGb/X1PB0abdoCAqt
JLDb/NcKFuU/8fr7Q8nqWY3pWzLcSNZIdLW2aa7IUjkTbSuoVown5dOQZauICaZM
mbtmtXNVCliu2NCwquQe+fQDb3ow6vdGgQHDZXaVOPQUQ9wS9CiyA2+Jf//mKxMm
/ZzKn/Euo57wnr/O942SW9qOEyrfULaaepoje15eehwtCJzzbquaiVA/tefy85bx
jD7La7Iu98T6P455gaM/aUPgTZsFHvOJqgIMtys8tOGTnHH1JAobR+cUDKszYNlK
Lj0Ayk7BfKyBvbue3IfsCHkz+ZMgVbFmEufvNnv+YtWiJKAsM8fRV1PJE07y532D
erIKnZVjblWTsyL0ldHytaARL9hGXX33BwloqPB2cir4GICsD+5SZuZi0MR4+W/1
rH6eYkfUQOOPyZo6JRAPIyzk9GAGxL+J1MWbke8aMwPRu484Gc4wgIdpu3xJP6qi
L/erLii3MVJoIOa5IJwL9LkRtrpqaoEcaHZVkfyqi/G0ypehqb/TDkgfQbRwTPWw
Me3PVsT9Mvlhy0zYDfzmoD5wC0Wb1vB4THpUYatcWvX6HAIGtWqVnZ23dy9YGZDx
tGSg1phTgJFsC5DulMbOXDmSy1QrokdMc6IxJ3HlYRH+p4xQCiIylQLzVOCyYE0+
IVX1VndaxKHkMzStebmS52kOwtbVpu3fYz4mgKzlGbLwHrNq9OgSME4RfM2kE8a1
ZrdRJu8X5NZcX6fXcI0pwepPNiAit4htqMkIOYJBBv+WJbVq0LtdZ39wetHEC6UZ
zENt8+cGyAeh7pQ7zS5ud9XOmg6AOKXVNo0JPMbpeOBeGplVuEkfWuEyv1XqqgqH
Xlvj2gM8ZeKk9Glo2yUqmuxImu2UGFmu0Vf6VHpKnVEFaXM+UNYasIGOuDmDSiz2
2BJpjFPsbXay5rKGRrRzq+tcMKR4Z1m+DfQ+mF4OF8mAPUDH7yUdRZHY+Wbcg5+z
v+bMmUVXXyehSx4Nd+AlqVSETaQ0dd5CXYz+4gkxJLkCfQvzDUQXmXlsI2M/SsVU
puFIXlY1VS08d9Ku+5o5lP7tlwx8O5luVK4KB0zcMnOBbz0RwsazLTTl2ynxkuSN
SKzk1Iq2Sz7NHDdS3PzOIvxPoEk5CfySWqpKERQ17+WrHQ15OH2IT+UOLbUkTOFg
spXpao1j0YqZSJzQlI3/9Tl0kJlcSOb46JthnHWzbBVqDfSwRtEDJKGMUQGbItI1
odLNoQuTIq2Vlx+MQ4VDqV3eR4LlVMIvgcFZnACI3b15ZvDvRcy3aVM2RUWOcyrC
t66DSzIsumEzZG19OQFr0UwiIzpCbpNqUcoDuYG3+AV0BQ01+oc9sl+i+Z9leTRx
O2E3vIwv3o1dMhHsiwSmmOI3C1MJ3HgqxNznsgS3RLdTnwJMV4DVUJf7HCD3roRp
8CRIeiwXlvzqZge2N72N/kJXmpjrrcQdx2p3dGpjU8JKv/Xf9yBi6WYFFWt6iMjS
TONrpaXBZswdWW8aqeFgwiOWYUId+CKQUC4ierY3/WTlohxmmvSdUyh0zRThn/Gy
lA/k3M8R3bbH89g+3q664+BczO0gyp2GtLP7gh0wAXk2VEXdiUmKkN3hmcWL603p
ru+U0LMDr7fpoof0LjuSkeG4mr4al0UV+/P9ir4INWwWvKMNs+zaUAq8hT80Hd9o
dr/0+NkLRyDCbz6YyI8UHEfEPbwnPI5eGWhHhmsXTONIYptLNlbPPCWPG4gpBeKy
X93bHrGbFkIWEmBC7r8/0htxhB/BOeRMkrEJ+JzkgKQdH/qSgrSkJRT9LDfN4vD/
yBTDd9gy1Zze8dweU11CwD2g8v523A++9UT1OBQRceu8INNiDO1ZqQHPzVQ/+HC3
wYhwz9ZL1W+is5RDMLU3r2rQ7ZqupBLvu7OJHpTqywhgxoSoHaEPGJ2wj1Y1D3nr
+6vK+HS3H6MRTr0PAOIEAFyYW+6UWdst0sNICVrq/pOLJTU6gixlShL62y2tfAig
r1pQVvdGJYOd2aUkGPPc4OCcenJqHGpJ1Gnm7ujouBMz9W5B0+hnPzil1blmuJq4
YAVPTfFv4IuNgUSUKvPHhmptLHApQJOnwuC6xKZpMJ4mprB0U/2BvJzC5K2uxAGF
42nR0peGhRvcUR9KJUzjUP2ytHqdQ99l/588WK06wBj3ItPoPjhJsSkDZZ/szyN1
9dRPrxOhf0YJvksO7zuFeAViAEMKLsCBIQMXsAxAlRF0Ip6TNeCSeTR+Owow7YnP
trgBdrU+Osw3uhJKOk3QtKMfZTc5lbPIaAEueG50OAbkH3WHNQuArSfHVnq7v2L0
64Ft8xbGGsBPQx2WAyW7ksbbcm0NCfcN944rylBe0BnJYXlIYCwUxBBqSAoBhCNI
2KvWrJ4dxUEnOfXUDr7dTkNGoNq3pyxYJY45a/41HM+I7c8hG6yjxSEFnvJBRpwT
dXpV23MWjbCZ2I0cOj/axyKlXtVGhzflEJne7q0P8o1TtN1dOJrEwXc/QY2aIJKq
oDCY+nVZAOiL1Awiq2JfEXPwX/ewsFeFT2ozSS6ahHTYkx6HZnMfcNleeZI7SOHU
xD828pNwq6BE/uPZSEkiq2OILMISuVKSjLtiQm6FHfd/u0cmFk36ejlpzmsH4BUW
1waW1gb3t6fUQpESyrRSjrKuLfLv2RZ+OlnRABLTJshoeSowkMlhB+9D1T7w3cj3
vXZAa8x2cHh6VFmr7oWcPYN2Tn/+CBea1e3Rjdyu2xE9W5UyXMqHIeRHNpichJAZ
9YYu7MPLiFSTNasgEkaUJ05NVQgxJQQt0l0KWpQ9kAlfgC/vgrytcaqaZEQxpA58
wMuNwZrJSZsQ1AsZUYvOqznhsbnp6ZVDlWEecJFwIKpnuHl4gpHEdRY6yCtlOkyG
JF+ZGnc02Idw1mtrsCPKY6sSIAYkRKSyxa5gYOEi5qiM4V28vOM1lmJhjKIuHFCz
75y4tYyN2IbTypijuMud5Yf1RhjJeueld0w2Hg7xiXS+R/t5VAb/bNDa/wai2rlA
EQzdlS7JFuRt8GCjQHr77huZMZarO0oU0PBelMr0dza/nXNhbdbfyFh9p1DGmQdc
dNjin8WW8/dethUnTz7wHPn/rwV+uuFgAZehD7HaKxaxa4rQezR/YMOAzMUlVOF9
U9fTr9B0Kl4zYYG6uN5poHgTBhUAfKo+cNz+b0s+32k7XrFvOeWXWqwzaKIF18XH
cYaFdRkhULyqY2NZvdmUMl9Hgnw3KUTWgmyT6ZNILI+Ci2hIH5s7D/yjbRGXoA8s
+WXWExZAGGZ9XRlDAYHHoEsEjsNg2FBOUbklx+zlkF9zemO+vRPksvZpVL4CztoD
rd1ypeSecb0Gi1Rcbq141PB9+LXkGrBKHe98nEHDNNE01swAq6BCM1SIn2YhI6dj
cbw+pNJnLm6+tAvZ7uGY31/3afpIoEOe94Ba/osB0CCxir7fvSNKw+iTQB14LePP
ed2brShs2M/1vO0TUgxWDP95cxIAzc5i4Z58tIa8jMUZe8i9xlJ6W2Aum4/TWXto
bPCayKUdVSQC5cggrkPx7NJmyZNihJ07sdUBfBtu2eXiWA9KSbHBJijNkgJ86J8v
2dQFtK+qeKut+ZNSkJ1IngHlrg6OwSvaWW+31hUa44LG/xfhbT7pmTvOBTqjTseL
XwQLxznwZiOtQrHgMVSq2+ZMgIEqYSvwSlV6nS/Gtubqyj7ts9adpDXIPUwsCJ7E
sp/qKK+8DoXiSqBduNyvTxTlAzsGhkBtWZ0hR+zoJEqtQLDO+WIsABJZ8gusHYc8
Ysv4QXxGD4MZvhhJoSVLQUpsfhHKONW8TztpnBUsXowkd/o1JiMZSFXufLh98LAc
iGBSa6AjNnR+2dykpEMQPvCAoFpAvwognvD4TX2VBjbMMqMv/Im7Ebw6Z1Ai1huU
RqHz3XFA/FStRtj/4jT8W4o+V/rD4p/uyZy0eKW88ZCjpeMZPvNMY9U2eRa2l/nn
BQ9pE40nlUtHw8wAIzwjtxEngTVkccBD2NakKYx0FQ8cAHXgP/9IBkrJBiBT9JDA
Rg7alIJD8XjX+DfgvFiN1XTfgKBjv8LEkjGyMwSzvCYUzZKbcVD1kNdcLFAV7zz/
jT1RSVPiTJCF7hjAn+iXXFUWR3iOn78tu3xbdp/d+u09VQBczB2sH/aVDyGNnPGC
yKmMoccHMR2ZuHOIlmXfY53ozismS9esl3xJGhh93CZ2nut/FMde//ARqtgcciRa
Cw6JZo8DhFkjMwepAK0OzJW4j5jITjftfB6fTL7UedMHP22/bmfawbWSIuXYX/7h
w4t2gexFZfxC+24eOMar28B021SO5LDv5XoUmRV6n4//MPAHk3pFYCbuyKpOSIKW
OU8Xd8GETMvxlzaFDCoeyMRcjxlOUc+eRCkDWiD2Wb1e07ilNgEniR1ycCiUz6xR
vlMXt0a/iiLOFWc3rZJmKNjAMFAY0edLJXXrCQn0+Oia7uB15OReBg12V+yLXERr
zTaZCFa+Rsg84b6NltJCxYXuEb91eL2rxupzY5oUK1k9R2XIeCJGcTAwq8LhmTIm
8fyDIUvQ2V2MDIt08ch2JcPZSML3doHgYjHr7dg/G5wURnl4ddJ+JiSzrRI0tPfx
tNyHCRrFTzRGPSdNiX9qbdIHNfkLGDYr3xgSJ6u6DCHX0Wk6CdzXoQBwPc0YR+7X
+l9DciY0Veorq2L6brBKGpYolsrhXXt1dlF7mFXj5UE61i0e8SXyAgVXvT1ETvtV
K/aPRdzMMn4vO8CWyUwRSNfdKuYTe+Y2O1segXp5+IN33kRUNtNErBUsYHt4NPDz
GH07G/z62hQg+PODjU2cLw/abG64/daQlCBGfcyPi6MnHArVIAlDO3arUgp02KFk
+5ulOUDXrJIH/PKcYoBS6RWloroTCWe8NNBqKb4N8anqHpzKLHjJiRCwp4UDQnz8
/pvjGZfALoUZJxbe+UKF34eIKs3t9nm02v3UmBU0cNgV9ByXOV70FvSBbICk1w1t
XIqWclgMH/fTjR+948y2nc5jhNwRtMTf7lC3EaCOQLUtaU0R7wd7JvbrWUBdvE0w
cns8TXWMfuqR2S4NyfiAHce71/agV0HdfvxoZ5G0RUQRWE4Z+BGGTRSTpebIgryT
Z7G4A82MRlRyeyx1U3M8sbUdd92gBHbPd7HSyQUUCmyzFeN7BoH6AaXkCCrF0Whk
3TEZKQKMkzBNkhsAozpfB7Jz4kcexJG5TdyqVbenDVoomhoPxgBQutIro0nlVHSI
h8OGTiWh4i9ElX4WQshHdHcdVpGOzlYnZHW8X3sFSyHCksKucsiuiFAXGyZIlKBH
q04tbF7LuQUwDLDb3maT38Vn9Zjpil4d4Whf1O0Uy4I75+2zHGMadYNgJ+SVJ3Dz
+CsOx2XmfHhHElccEXNgVLVggNvrkPOi82puwc0licYrIbAE33EbwhJHDIGLUGuY
FX2IzugxIpgDTqcMABk30lhXPBkc3NEsw7e1XzFGmogzUNOKRk+CSpKTbojgEaPS
vdV1lJQSyfhZHqznsPEfyeF3Gky4ETUuMvEMrMqX18Ny92/dlicLqGulEM1WxNgj
20PPmmHnWDQ3rOxbdFoa2AmAyoyAe3ZOGnRcbMSw1s2aBr/9H8CvQ5SEmDGD9X+Y
bD5PHciqmw8ahLWvMEXkezqSnx/2bxHtXYuI+XYV1QTrJ0QvmU9JzA+f1pYPE+NN
vSiY0dNGbz3QNtGrEbzHJRJYEAfBpI4hxLq+tcgJ4CD8qL16UnYnptpUVcafcDuz
pkKDspkzdwXDIDpxp1Pm5M9JIjjzJ33YCGjX3kl++z6piyP33ELRavU4brwB/2pU
Tf2OsCibTVU8gVyOxnSxNbSii3J3oTEnJXRYuABuW70f2jtv81q1wiHNncxFqZ01
zPEdEHt9Fj+Wss9Dj0KL+EBlOt/MgCLntKbjOD89S0tVLuyLJveXUCQd5wiOwXt1
RAlDy/6V+rM/LuOZcKZoyWULYqj+GmE6WawkFmX6RCW4ZaDcAu2gOz3E0EmVSv7d
zVa5MV6mgXudT8k7/dm6EiTiDpZSUj9dzdlPPxDe0w1DWwcqIVvIdW4uMT22/3n+
LHHiXEKKLD+GbRn608VHELSHVXjCVZ9ReBuB0ka3H+tWXWzRekWrBka4uV45p1AT
UjeRavOD82QcaJ13eJtmzCn8otX8odZG5We1Z7IQrq6QOWDsie7S1jfZEqSvv5/u
Ti3Bnv6ExxsZX4rJtotcVHfxIb4z59XA5UAk86JRgw1o+ypDo2v/VTkNhjD7+HZF
2ocIMftfXyXZ7XhfOeppoIjVotru2AzeJRoYrwXm0/wXTwC8vuZwtSzoXneJUPQG
lIjyFk4t0P3J21AzeSRpGoIgUwbV5/BKoz5W5qN4HF8CvhFGnFVluCVZAkDcMzma
xoPHZ6XslNlgQ+dV5lpRSNDlUOr7+3VGd0ldgxDJOtteS8CI8YNXGOteanUOZcjx
9RvrBcQCe8739J/MnRVshGIYwHN3URcZWOtotjEtnyV67mAuIH+l7Gygm/IWfcnw
Bv8u9yMi1UbCtTF0o7gJoTRuMF/wJ6TUezphDIZcC6lgw2BpjOcT1mk4ysCBOwgm
VHguHvu+lqe+0TJhCjOOQq3XuYOmCHK58d1O/JcZe0AVYtHp98uF0DbdxDTLHwxB
PsODE/sucXz0i3YMMsm3qg/dvRwMltu6bMgIhqPDs2JtHUnJDS3vhqPqpsvaFFYS
GYlYsFle23NkERMg3khp1dyAPpwnU5A3qri605/jfXZSYq9mtICLo6ij4y745kD4
zE9wGUxM1GavPIZyR2YbGzQqIyl9FnB2bUdLxsOwhxSprmAZQMxCvXVrv+SmSVjN
xJsI2a82bzo+MV8td2AFk7KJd/Fd1PfAjTLxy/Sgiq3Dc7UISju8pcXLJ7BND2IX
awfxUm55I7TS0PF0S0qx8Ueld6BDlThs+6jpJVi76QwsyCmx4eRXS4Ag8hXnqVKc
pl7ZGnILMfiutTB4kTOUAEnjeloxAN9BO3qqg+FESXctuQSaRiBpfVTjRE7V13Yw
dO4PFo0rSWdSP/218X1SithWS397Cuei6OGuVBXJDtsqpEojFJ8h+9oEDGEP9PR/
MAKmcdSllDiY2mmCP1De9st0r6ygwsZqipcCpNQ2zVU3PnIxMpYPKCw80/zRToSR
KIgG0JsTxht2SgDDhjc+6muRddeW3AwdwoGkzIvFmZ9olci5SI5OVZy3lefAgPuh
MxIBJLg8ieA4KXP/F/F4OzIVj2DbRRILq/wNYGxGra6WUwyyF9m64d8kApFNJd/P
2+XyNknoH8Jh3NSVBLQZQV0cZSZHKLaoB9GbW3b4UdxyAJid/GO1TENBit2ZYXEk
TqqVaUreGmGfj0zJFdfGQNjS8xtv9VD1mylSM1MKLi7W59POFxd8WNKhBxaGnOsX
9TDu9IyvF/vmSMNectFKTJ/XP5LT4TB3WbX2c5oBdQTNQY14fMJX1RUVXy6jxfQy
xQsGzWXlC2wTOdAXYhN48Vxu8AN3hfNpvFLbh/JryKkVfuI2gPxOnR/pIPqZmc6U
tpvgUdfrVMm3DiPtfoKMAHaPt+aQjmpSa8z4KRm19dA18S/ImD6awhIsaNAWCjJ4
EEeMBEDVCzxfqIAevrLG/IYryQJt3Vyq+S8jcJNAIncHORROZ4KofIsdypBhDC55
bXkt3P7Uoki9Q7qyEMREmxOIOsfFgVjKstFeN+Hzl6B8MQkD0IioivKYM5zGU568
32d5XZFF9OiwU5KNdn1KS3o0whBB8wg+n2/XIkf668+4lOVkbFnORKhBzH82BH+Y
LZPx8gvs4z6vnVJ/In7iwllf1n4va/+8WyvoUeFiC+Ey5rCp0oLlMrCF3ENOuOz8
GvktFDdW2KwKHR0wdyioe3oahycnxcXHXIvJmdn26KeaN8vaw1rEYtYvYB+T0t70
ia5/dkBvuEiU//QvOB8ridmUoZ6vT+C2HFUet1I4a2gdbjTS5HS+/+/5AnkQKSau
K5XD3iHVu1o5PS4r8NkQJfPpT/LfAnOCypUP8kD00B1eC1Ev7SkG/KzChzolpdYy
V8iYN6Qn9cFJVmdFk9ftdd6KbB+y/zScOtxADtD7eFndmVWJTv9LiGyGWJTg88MI
xpDY4uEwuniyS+urOKaPdnIqwvtr+75glnqXxA9x40ZIdOfQ7qRRoprNCHzaoVL2
IO/aJWF1x6zekMO7sLcUfjFI9XM6nQOD4GGQAuRAB39UT/K+yFmcKH1TypRtm1kP
0GKy+0RNTJwcQbJsksRRsVASFkUvKMVfN5PRb6B+vOHC+S30/dxC4EkcPT1ev+GC
+Zzvy9n8EQBtjllMVuqQtlTSO+b1lMQ6sb0f28YQvnDf35kkO/vXV8f+CUTW6NE6
9asJ6fUpLy2DKOGKv24UeejjrAsuHBKJSWhnNcVDYEvJprqV8823g/ebcAVGxnrH
1neK+gJMmrab0tCKi8k3xQGA8wuZtT0SusptaCPCsnG5aVqa3PjQPE6r8PW+B3eu
sGpo3gvkNlP0vbOHS7gTfLUTY8OCkzHj79NhFjp5/5yCq+t91iXke2RWSeeQfj1d
9c/UVPm8ppyp2JXTmHy0Y3qx247ONqn4bgUvBc3sXbbhpaT/MhdrzwQRsE66VA95
Br0NOt8zBurwr56o1WpFutWFN4Q6qo1oVTB8r3xfDjd6ZWtzOTjjUBA9LS+2ZQo9
29jArudvhM6s1J+vaDGtSpPC9FMUengK7fuvZUboa3mH9hCG8axglVnHtWj70aW/
N9jJf2KlwVIEHQ9gnouS4TC3wntxoO/hUd67hm0PYa4cKfEaD7XdPBbat+yIDnH2
Gz99DMd/KB+C/b8zua19kp3KcN+RamobWA8Pe4ginG7UCljxluuXBvPQo8E9Snwo
egrD8fyXTGgdx2TQllSkrCOVvdU279pv2tsUZZ25Pyn/f/Kf6BOmxilfIWud0Q5e
VbmeZcvxsDepoFf/wpKLsRr4/nbkuL2h3RUSBxONtUhh3j/sNxm//9fHBxIoDNOK
OViP5uZ1UpFi7PDr4E3KmfNnUdMD8NpQFgvdvCsLILnuaDFr2yBzDLaCReigPn5M
aOQrDOvxg5i1GH0yAn+6abl0PFU3uSEoiNIhHZHlzdIXQUVGsou2xLh9okjhIMJt
R2Ap4MT+M4OHFIi7kEIre+dH9cFCU5yMfwolA6Ic85ieNb1ZlHIg01yp0V1efcj9
ynAXpL2pq3SuJyJALkTWa2NRMlNrRiga+4AcOX+iuy1I6WUilaJoAyxYGac+jK52
lpVrJ/w1TgKLKqvfrHsnEgl7fanudjPSXCfIEJVi6fq12auF/cUm6WouSbHDrgox
tMdmnwuvU1OvQOp5ST20/KwsLZOOaQMz9lFqCGfBjFusL53QX67To6ELsEB90amX
g9sAIvWoWvCg4KUDq9H30aKUPuYwrBZTpxyY86nt13eC99J+NI1Mx+R0EVp+ruWI
ErE/Jj3n/GOILjLIT8zcn73PDVIe+CNUc4/PEPYfP+STp5oX6ICRSqB0t6l/qMuK
s9cl6yjw5SvxbXO1q0Xno2CHE/Y+mDiLcM+Kew36v+CF821XwN30mcPeeoffv5y5
3HyCV0ARB8DwS1YZHkHI8KrPCwu3YMehRbT7cAmQufyj3naJYx2m75Vo/cYLapaX
hQZ9iA6n17AwDwVCa/SY/mKuuRBcSBKTd2/KDva8XVK6H5TMHfblG1jerHnwXTrU
8CBnztgwPG6sHQCVxCJs9V1ZA34ikmjyya0RNxx9ERwRkbn72Ed3VINuUzFxwLcx
o0DmdmG7+u+Y9vdS0m3QcbAhqLx5lCLUuJ2FmTZxVhlAV+p+Rg2DDcUJq8cjlNUl
E3n7/qyWxfRsC/IqWHmWK9YZqykWkBxn53ap3EvNDD64QlPylLjVAjajMcPyTkFX
ZLvVBkw2ewGKxxr+d8gJvNIwSiQvxVsbhpS1ui43IAUedfBdzf8/RKgxcHMpSfqy
dVSLY5b1Nged9JQEz2ie4zH7FeK16Bp/KM7p7cKVdz4w+vMxxvM2DWg8fiyL/yfq
K03/xcluItEVFmjKEa+l09uqdzY85LWjLx8xvYP68Nhq5kGw7I39Y7mgXmC1TJx7
fj6pvIkx1S7IEVQS2SndTPafxAG8VmICBAIH7FYMP9KZbb/4PU+xuO60FFFlSH+0
Ad0e5AYtibO+mEYBlYvA8VkfeQg66fk8gamxLigHDJAQrny4SH7KwVkkEhwySTkO
ufL2b8/Tp6gfXP8dzql+cga8iJwf0pGgS8JgNLYWZOwx71mxMB00gmZDBJRCbL9d
OtSPy1ZgDwEkPQA2QqVn2J16T8EyDvhWpjMYAL/DpgnT98feaOXV9mpjUjdviUWs
7N4hzZtVrvFOcO1pVnIs+k2cmooN4mNozXCm545mLDvwNk9sLhyGSicxYAKWS3++
nBmGIuJYDYOcmOiIPi0amRL+rF9CBRF10ooUgG7I5qd3s2Ma3fC4t5ZIEkj8jjDX
MWVcizn53rZcwqPmdgtM0veMH1FzB3q/HCDfOsx37scCzebnCT2Ic0wkJE1lgEuB
JSMRh3eoVuSoUQfLSc0rsKyN0ibBxRBhDQtbDFCCfvRSnCYH/RVAnv1pq3C5vgKJ
PcLz1YmCXZffp6iamhym6iofJLCrsYDtj5JWskjCe/gm6JzwDyv1BgPGF95hCnNi
wC+BzLhjYiXNmDSsroDoisRpLF7OHWTyUS8n6fgNEUeiu+7fOGNLhjCjoWrAhEwt
zxUsRppYzhxUQuy27kvyfRmqV8eRW3PAnTft70D2nz0yTOGIsljhDDUZxTBoRv1k
BdA8CU1fJeCv/BWl4+hFHU1XiOzgd6Ni7R3yaKhktakx95HC3L2xFISeR97Z2bEA
hTM6E8zpRQVrdhHcXV0qNhjS7228GA7V1kHnjXyw6aX9XhmQCyz5zElfhQw3O0vT
rry5C5liOv9av7Egr+0RswEOxLVtTbeoNJm2pgX0dOxtDnfMAG+bcqQkl7dXrrah
Fnr31UbmJ7UZRheAZO4xOnkxBfuxlmIthcMBK+axPnhDNsE4gIdBylXdLstuzi+x
/5rBq2nLvRKX05aB+fEal6hYPJ03NVC4XhAgyXKG0kPYPTFkOIa1Xv3Iu+VgWEVd
TrUTD4tMta+jzXaqUnwFSf3tuv5WmGsExIls1HOCFFGfq1c2Xb0PwaNEK608CA2q
Rnt7sqNce8FkOmW0fFMI4HsxqXNpSx8VkLxOLeSUMPNbmBYcH+ASGyfRi+gYRUao
leZNwQjQr2riy+JfYbk3WRROrrvAZUX4ObIwKCRTlc7jgjTj9gRd4I9TUEqFw84R
kKpNiSXsGV3IY9ekGYYtYzqbZcIiBg5MMwxhRJtPjej/cyw5Dl3AaDobJoqW5el5
C0OIQoLtPC8+x1p04ehHoubZ4ofSpIvJdWMVU0XSHJzraaTkhMWorHrQgKBi/SXD
ENCMOXt/uinnFE4aHwRhG8Ha/OeWNuzkd32+AxLHkS/hFGjDAn1PmI6A14OwbGjG
LOt/dWpMH7nyMVfrKnBqc6MwuBrx7aZFlfS2wMu5i4tIfrq20Gs7W7uHh+gAjrJG
DpR6dqL6UGmGa77UjEo7G0GWdbZwvadfbwl/PO0J83c1onukQ8fb3nuTIHgy4hUc
6doaqvsx5rCxVOnftSyW2XgvAFbGVrg5Lo1fteIt11SK4zvPIAFVaPQhJlCHJNG9
iwFo1YYCch3FS1BggWlXlBDrVOTnhpkBUbiboCi45+QH/4id3stI0MqpHvjYmz+E
sOzy4/DbvD4+NlXjhj2xc+frTN3bVOdKnwZN2kZ4CO8auumIap5oL2AQsbkOfnfx
5fcstl/8aLZVCMbb2xuoY+9MBDtAmuyoi+/1RHx99odsdb+LHTDwgAoOZP53Wuu7
SRPBkwvo5FumEA+A1yVghnSoHXqQlUVco8AadTSdViUCWdqDIEL7EZ7ZzGZeUcua
+3iI7CT7Swah12CHwslMWO/4h62TxERdPNTlsZzpgK1ZW14GzdFJOYGTCNiti0p/
Jedc1OMft+dAD9ymlvpsLU8z/HGAvN9xhHoSApyh6NuIpNZnQM0a5CNooRKTh+RO
UNEzFONVo2N6+yMV8c/sKyQC/bt/TunITx3YNwQJkCo/eUjHYuQRpAk1C/p66A+M
7AU5wj1iLEHm0axVXFf2G8LVHqo0evD/rrthxAQYuZWfwTvdURM9xxtD1YGJkXzX
GDZNu/dUfVkl2hjVe/uE/S1+Au40tSj1DrgIFiHD2M+/cuxeCR5+8n4YAtNSvGyj
wok9l2xzjBRiZ5GAsou8pgcchphkHcz40ikvkDEnZhn9b6HlqcFzLcrxR8srua7d
fwF5QlD/u7pXyqZnW9b0ABTkdbv1jHqJUSYFjZP2vSgAhUFHQaBbRjloUMQXez2w
69bunZ9uwVaxsFBz/uTOuoM9s8dVsVLLs9ikfGAlBm3HS1xWKCSl4MyoibFG7lni
`protect end_protected