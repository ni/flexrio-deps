`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36704 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
iOS4T16637ogvUHHJHvO1HmsKLichBLC+2/sfbmxY8U3jfdyMosn2gBQ6C0ju6S8
tlNJwlOL9wJUkzptYblkdZktOe7/84dAc6v8XuhbsHuoq75aj+j0qASE2QLW4f3E
Foyds3OC1cIFGN59E33gytnDnLN68KiQ4NGW2AZCiNB9mD2SpZO+Wcpz0YXD+OM0
tPYFZzGqzyiebi0Abknlq0Ompf0GJP0LTwUU9Obva7lbZMD9OTwP5C8/8ZIbNeqi
KgdAFFC/jCLdDJBDAVsgUYhjSQTCvqrggsTjfvi3qCBhv6DTDIldeI005ZwnPc6W
uoOCvVlfjpiatsc8orBPR8Q4zztOqpz48KFMFfFODkaDGQH9NZe0pOwED804Runy
JkZdDrVhOi7kFMXH9vXRAYSSMu0kS3q7aWtDBaQWCpjL3k0Yka2zH5tpBGF5Dh+D
ZJ1upkaA87p9AC3TYuuXL30AdlvmNRH1zX0w/p2dmj+pOS4+rqczVo2oYOS2RFLN
99AqT6qRNRLVMiq1k10U7xc8BxU9+KkSgJxZ17/yKT/ryR/I4ilsAdl6HijKSbaP
MhuC1drmKd0nZLiQYxwDQ1feTNDn6l6jIcX+lY/QUKMjlEQeL0jF0clN/NfmxXkE
h38kTdZOiPtwdOw205ppqrkueK+qEtXaR3fq1FP3fEHx5NP94XR4eTnP7y5Wb/0l
WWEo08XeWQjjEPDs6VBs8AI4Jm/fNKHcTOrCbSQdihjZVBJhYhlxf8Ch+raax/XY
vL38W/Vtyti0Fyp1RqPCIfgLQDnb/g2Klubz54HCXK1kenU0S4BPksmznoba6MOl
ZsI06KTimV9bKVSkCI5RUCBUL8DFeiYxjfoxLsmNSLgvG3vr2urtrWuGpCo3PhDW
0ykIK9yY7/47LPT+OJRPHATDru4UcL8L57wCH7qBZ4mXsexcEuYI07haTTEeVFVo
lax+2kMfi7qtOnLI5Ta7naLf6QrlveoThzlxjOUT73I8b9xu7KPEmND88G5fSI0E
tFQeMzUgyQwqW34GQa0o1KHR0zlfXSnxZDjO+sJ8tZ8xF7A7q796sFbcVVyYJrut
6J1URxf/C/D0OX7HUa8Itqmb6G/rH0RS4VjInI9DwQI24AP0aZRAa8SSxScJ4zEU
5AwmcBdtYcApSlM4Y9p3goJOGZZ22UJ6OZaGl6ONIiCbbHrhZskjzi+etdsS+oi6
3cJr7Y4B4boUfVsqGChP44DWNiM2FFmShrTOLEyie3K/KVy13xatUvcIzM0OCQqp
pWz32l0clyORfoPNWpbfsxpeyy78p/aF0P8KGV0PRete4ywIkk47daG0y1iUNMFU
y1YVr3ScM8sdgtE+2oOjd6+yoZvBxpu09UkqFjkLZxV/EbYkNtbo24dusGmtaS/t
rLYTUwMqPwLgdKvndvtQwgrObCHcUtjzGHNeva0oGdPMVMQdGt1n02LV88kdzCZS
VuhHnjLIXYqNWhWjBnHtkoX3OCwn6edv2yG/W6ElWYeix2+DQn0ophkHJtzg3/kr
1R58geGCx1TaSo2otoaO/gB1BU6fuUr567nrB8MQK43+yICHk1fqfTQeZJDM13YG
VjT9Kbp3YFQ21bdRRqQQYH7Om8lsXCUSSj7lBfkREnYRJTOl91vdIcOOjjiFpcj7
N5Hm5JfBIwRZ4mRrGsjfTKWQOtYQYA6irEdu84zONXu17RWV/1O+uaA8UoarZqXb
JJta0asalxIskdOFivOZ+f98IHKSJeoeTRFfr8eJrVTh17B7v8WbTWLAY4jqDjSF
uRCXs7XbyMfo0B9By8azfEuxOYztdmExyH2LtQvhH3KlBcjLjR0isXlapIuq8P7U
EO3EPgeu0OjjNaluUJtnPmveywrOmrjJeM6hgIxxkTQHJJmiAjL4yasYA2TNXLPc
bz3kIEwJdvDSlTE5Fn0ZVlGl+E26Oyfh7hy7Yf/LrdWJMehnB5qjNdYlQmw+vFGt
NGjKjo8AkVr28eMpYDEogCDQmbOIWg2qbYyVSdhmZSq1rQCZbtJHvOip8+STO0Tt
ENPmAwtpMWhbzeahjtfbUIrhonLWY1JJvomYTdhY9QnmfG5EBVXWdjAXINhYfVpm
v+BgNq1Q0YQn9vCbxUGM8Bo3mGInKKhcfhB5OpeUtF/VD15hTj2u2DJ4yZq2QwEM
Lica5KgW2ykeNDTEJmrypaxTNxTM1NtoEKDZcWcD/+z2FnXGhsIWo9G6Awb+AXAh
URcrAJmY7nwF2LEulZKBcleNMO9GeriP6PuYStqPVfAYPOAKT2756H75J31bQAwe
ctaMrFVwGE9NrFpVFy/rlij7565Ef/lgJZ4rBBe3EynSxpDRw5oDF2z5rXKz3/gn
EwbI4h1Je7ZewV5hhaoaKGpxZiCrATQ4U4Rs6CDM7fT4FKE2rbEI3Cd9IYNmAKPY
v/Tte+ETCJ1p7IVYnSS+WbMd5Kcw4XunU0Q3P2FtC2qbyFK0dFxhJiGAy4yRW0ni
3o2yXqQk3J3I2KpUIil7Qp2XyTWqo/vAQed4siUF1FMurMcmsqAZ95yAt35yM44Z
KDVx7vAVZlVgYLW70CUw8REIVH0zlYUnbM0pjNKYHmZ+HzxUr20vz2BHZwz0yvTt
ufGaOjj1zg3pjiKSchP823RHuDwavG4meCIUbulykl2YJ2QAIxpDgQyT1+4aZJRH
YNNy8ErcuyY42veWP6KJEcEWQbtbfEoXW9U+s7QJ3PNBviWAW7Av0X0/x7yjcKgT
IRpvAqBDH7t26ZeVTtWaXVUrGIqvVcb+ug2VI+WDQ6stQVCsOBkjF/U3FNq2Pjwp
Ph+ouG+Ki/FqD13YNYSPbMdZxDdoSbDA4rOKN85LYlonRIh0rdnq4ayF8f5RWfBD
PAJ42/OMKairWuviNsu3+EaJj6gxtM/biZF5ccCw0BPw2VMCTVNcgWkABzF6rgz3
TsGvKsa+r/ApUSMUGYPmDa0VHC+vvzQ1lHLbrUwoyJ3GIelCVktY7SmfHVvWHrBn
GBN6YJ+3WQnN5O3jzljvc7lorCVdRshNIrLHXLFOZsgL3AnfiuHflbOqLWfiqVvL
xws8sWpkctqF4vFc49odEiAaKeBuBqwOD3O+ILh8Cki+DUkF1odVc/ZpdRfpP6R0
nPozB59Wb7YJa6W7N4SALbw3F12cq3yr9MxR5Ile2658oxqJUlmaJVglfSmYZLxt
HqGe3enUQSPpuzTXab/4s29SSO6eozqA0idBjeTvN8itGTQENyIRibYFMS9Axvt7
noZg29uc0DdvoThyT0tcAkHvZpn4RKXE9B+wOVXAQOWJHj3Oi/D0T6fLHQh3Hcrv
Jvy3/7RDmin2Jn9R2XtjdSNPb1O8iIEF57iPXaMmKQeCu43mHbaM0QvEP8XWREEt
NPSCLO6RBxvx13GblhNhHTIAZ0mYqsaoc2ZXeDvi92k66pUbVr+bCtDBt6w6kM0a
uoa8cUcioFjHYwHjq/eoTzu+oxjQCYqoc7jLR3pTkk7r8cPRkDasfyBHkBdMKVzV
Xtd3IFwc9T8fPjxCOKpbvaVqak6oofFzuiMT7RywX2Hdu4Yc69PMMlGv4OF2FSWv
gsNeCf61jUYCNIn5LuQxxUw8p218S+s8dHl795T8ENyroJRvP0eYEope8sCJvy7J
J1jmbTG96Rc7jd0y++CljHpey7pDtzEPusOvGCtiTrdt33iNjbcM6+CgE55AWhEq
2B4G7O9Qn/LmrO5F3e2WII9w7ucM9vlD+g0SIKPYJWJ1lIeLmtVKM3nNPfCmXGZs
5Cxm9jBYPEdZvugH/EJmk3sJH3e02Z7D4EkcW+S4SdgXnUNJbyrB9j6Ky3foqlAc
YS/bh72NOfN7/Is1D152O8PEkAeKhyO+HaouwKHBj7d5ypJMCtugzJq7FI2Zj/iO
Xr/1hcptzY2/xR/OPzz64WMvOFctsFQvkqMyLz9ljxQT0cM+WFweyuSOmxwlXYE/
qNWJEG2XXBQFvrCcJJmY8buEufsk3Adl/RfVyulFTUnqz22Rt/pqrG+bRsMyUgBk
KMiePYvLDZ3HnWmUBxIefw82T0ODyCUkvnhlGPGFj9Di5y3sWDremdI4uG2+gYIV
32FTE+LV7rOrFwaLrdQ7ReTDRrrQ7U8EjaZagx0np7WP3zAZlAKDBFf9VMsP12Mn
2P/k0sTzrZzFk5mcC8Uf+hEh/WmfIAgsvbYlfDbCv5nyN0Oyk9w6esUXOVnqqZZM
DSgStvWc9Tsqbnr2R+4gen0HN968UoAliCJ8pfG/R15QHM4nK6F7NdcrDmWMiAjd
sd+XEGucHMODpxYKHcd8SgE4R7Z82TCCUtp/gHox7zERxU6yaiLM3fuqUt6MPFV1
sug4Bpdu09dAFiU/MYQig7iG9xUf2VlCLg6hzOwgN5Ax00YQdi+f04mUmYXI+0RW
t4kRXUR47RFAVud1wMZi8V82iQYcm+i5nt2Ai9TtYtO4y09LMLwFhu7mwjPuFOmE
aJT9RVcEbxdCI9QXifneSJxJ2wG6MTkAUQ7ntxwirH3R1hUsN0dbgWWwpeDp2U3L
pwEM7tkvMLnfmSwcGIDds4R0u9EQa1/dHRbXvrNkegIlK86cMRaK1HkhN7CC3+Wk
cf1QT1wWKyln99Cuyg113vhA+1naAYhXAeFmK4g0ZXq9UeFPgO6x88DmDIBHw4m+
Yeqp4mH+Im4f4MO/0kQSSvqcup3rYBMk0Z4R4Vlq58IwXNF+EogtN/6r3FlwUQF6
4bbN5jh+iCTImLM6HHUF6Tna/ZPvdy3sfasEc6HJ1C7m/3Jl8/2uUlwqntt8g8Kp
agO6x6z4dDytydRoIDbmQpb7JwccNomlF9DA7vMy+md6GoE0ieLlhmeytpdNdnsJ
Bu4mcy72oyq08mJmW/JFjgx7X29XnNie3IalOkOHK/gHeIJL5tDwUgeqB0C/6ncO
mkLR7bBifTG98vXzwCD/aUlBDuNJGrcBo15ZXBYzOvGakunyzWJV4jCYgffKvUV6
URGfWIZGEiBgo92CKLRW87yESW9Q6B8FP++l2OftpEDQcZ21ArhAIvLxessM1H/U
2rUPjJ1EVFhyuAq7mMl4tXvijWIYL9dHjLEGFztYGW7D+C9fctf0FHWsbcdqekHq
eAj/RAFbKc5QibDiTgJIJJ/l9B+1VQZXxQeWTGyQarASEbMaUIP0ls7TMNFRZSoF
L/irkhwv0V0t1VDoJvIYfltuvpwbntgtrnYEjk5cmFapzewxsETHeypJnuOQ5LJI
BpahMg9jV2blFC4+iMNAPL+hcGTdMqfrvVSj1dzrMPNRfVaOVtJ9AeCA2SuvinM7
fOV/NLlRSLxAGFBG2yqib2IlrH3RLH778QOQ3UMhBBZwNdUDz49ikLpy3+zP03eE
PHGHe4c+hNAERjCwx6E9tRBvdni1gkdeiKneh9nBngF1xeBDbrglJaTbQbBFrd4Y
qqIdz0Vi8MV5RMwgmMiQVU89beUjpJJC1CBc0mHD5VNlZg1XJrIvr0jozhFt/O0D
ms8BLYbKr2YJ+iDaBhNxQtgYtmJmPZt4nQBFNd9W3HqW/QMdl5hop3Et23y7m3S7
hdpdI+Ri+x+91cgScvaMHmMOix/LW1OW3GbPSsWHAfGVS3JZwMlmEZ/ZR+0YaX8U
GsIvN5Mf9Dya8IVyFdDHk6TSWjpOUmkgJkwQRUusBr6Xdcb86s+7IOTxeMfRJv87
YhH7goDm/iN/89r18pyTT8nX5JwNCW09T84G1mbeW34ufne10YoozvIgQCv1X2vz
fAZ6dx4IjlVde8Lvs7Du8GAZKrDYe0npb07UYQ2kK473p6ZAjQoGw+4hZgOxvVoa
wNFzxC6uD2pRSkA2ALrA0GrXm4MWWq6y9WeTtbFYw+VpOeAnDgW3ACrwnSznNYYd
qhJgi4x8m9A64zfb5RYUA7xJBqHAB2iXCbVAEabiVS2wFjdh2XLOfsfPIlRlou2+
9E9bjMzGC+bo9dMbc79c4N5bHrk73OjW0uA/TSLfaNSzMkkMIBnrSQtC9fokKigh
LY3x6+yr90P69Ei4SAchHc7rG6wmMjKRTzDYeqJXVDfwkRpEAL3zFCPBLEVdiXfl
C8r0UpP5q7igqOh//puuyd+8pWU64GvH2PLxL+6xyUsw9X7wWpVe4+LE2xW1sAPM
MKOBMeUrRUjDARsRa8x70CQCGG6n1V874Jkt8kuQHfN4A+QxJwAbWB73cn2HkMQK
lUAPUSCjhrcSeCUKgG2xuN+ymbcLfMAoiQcU7z2nvIwZ++8CqPGkzGITW7EvLMes
Olzr/XKvkITidIv1FAa18zx9Mv1uxRyGNYDXtQaIIXFJbb4CCE5orDwKPa0pCAAV
uJgFqice2XCGpOHivg4C7E1VlqmCPpdPCuozJzPAJvZJlo41I1QO0tNncbA+lsEd
cfPlwGXY0FzmNwIZaqLKmwbWgFGW6ExXptIvelvpCswYwIDGaL3GcXLZBUMvErA4
h9wVCGbG5h4aM8wK3sWVG7OD/slW5VuLxaXikGhoE6dH0HQbpNalczULlzBn74al
0VnAGbxLXSZk3DT57oq648rDj8SffWsGxi0q3uCMaiUGxYGgCMcKIKDCjgfWIHOm
nOytiD7OBogvn8S26fcPI/j9u4JHzNNpNNoCOVJbT0vZpsqW101RWgopQi87Q7rP
4FAJfc/EhHBC9XF09Fkw6UXq/UZHBiFiq/OcJUlrt+eglR21UIyfSPqUrFhh1oJo
UB2U+88NthDT0QtWeYUV4mMHgUVtmri8HvTQxPiL0nTYSNYlPTOvbQQ+AtV1x5dy
PyFtNZLwfumW5eOqpnEfLaaFEVW4UVFH9aZSWlNAx/KsBlYWewTHNZ1bDheLCESG
0KM3qOZvC2nX543Cbp+jLDOGzsxSWl78eVlDZSPqMFsnbsUrKZXsPFOTEhoHRhGR
YRzVSUTOd11skNOwnOXmcKkkp+XRxBOvx/4O5SewFnHX469elupotxAiohrMxPzV
cF2mjfpU6zxqV56RV1AZBWdnUjPAPD70hDTnSiX9+CS024X1mF51eNovJ/CdYZ+J
8OJZv2TWVWurFnHVEu2ueUDMIAslR6NH1nryk+tjG2vlG21fSOmOpdiTZsKMRKVL
YyLnMe/FjNGXHslW5xyxYxxSmcageTOL6/MvwTKEfkiQ8n77uCKoX3e+2l7x5Zin
WsVl02g3RCwl5Sn7d9OATOce12SzhtRMW+WiY86qM1VF5x63mQE8q8eql5IyFv9T
LV5mqJr6PQQZXWFloFm+Go6/rp2jPLTPyu/9CcpdKYclr2GVndQAk4O6k/wf/rl+
SqhaqUmQ5TFtqo4WntJyPEXYdizVFa2MuBI95ArpcFvsuiejeZDaPKo5QNgnrNvg
8EmINYiC10PDtkkZnKeIPrUc9xyQi9Cny4NlhDihN6eUilYIX1b8GR0CWll6BLtF
5pJ3PHtiuAenih4Xzw3ZWpmMiwFeCu8nCoIJ+TZkx0QcZ9bhJ5NjD3g6vJdiR0jT
4AEtQcYLZBT/ftNdrXS36HS6K6F+W3ENPUsdP2E0tz53bvhDJlPSLl8mjvYWBtOR
s30X/PZYYUPI47OOWqdA+KZeR82xkUyIXg/LL+6oOK5yCyGHwGDl5g6UDJGAxruM
71jViiLd8Ty93bVJeN3K946KaLxXImWE/tPTJQThE8jHzbQQFcpwR5aHRumDeP4K
1YYh4Qb092Opatu1Y/Vi6VidJuozhj/kEFT9k0xuV3J6nlTCWGo7R1n9LPutK/gH
XiS11FdY2nwcy+xize1eIFlnMvVrUmw3kw+Ha2Phj2AWEWPnLi/9G/mWLyO3PB5j
CgEPC+uzo2aU1cLx1h5tj0fNpPrWf81dPx7Y1d+dhj6gWduOO6E0mKu7rJaXNLF0
t4kV0164N9yb5S9ndDprH/YyvNDfkt3W8LobE803b77S4K/KW7JX0fZwXAkJLzIT
7uvG+lTF7TRHxYY4ACubXnqPNsp02MV4BB+D4IdrqF6d1KoE7mbA6BdzHYHGOK4i
0AAfCxLKEAFf/3SpONJw9gb38VSx8hWSExkUqQB+MLC3620ADbvlrHxJlOTichia
GIrwyEV125yAkiFuT177+Wo7cOJXdatt21J3410Oq/rdGIHoAyetY+SRo0NFEyhO
ADQKiqoprrT/vNMrA3+Tmktfg1zE8G3F2o+b2HjFzyBX0oP4efdGX9viDVVONNBx
6oHz3Woq7wCbkkjOEiAhNeBRtIOs4cllNoiNkCNJhdqo3uiHPMalwVzSFLC83E8p
xRBaRy133kMKAeQDBa99SvrwMpoBrg2xTEtyvc2HTtQ1H/Q9+U1pUcsu6HAtKEMC
3IXTX46ypMugFXzPA6H1H8/M/zar7fP11ZZjxS2VMNgX5P7+jnTGLBIIyKj02UZn
MAyiI+a+6R1aGr8woKXZ61IsykHqDTztAdyOxErqTW0UprWtXVoYtPkReaa8g4g9
Dt6dw9+BK6+crbwo1vzf6TJ9853G1REUdVBA4QzbeAxfG6zciGPMvtjcFr96sIN0
Hd+cKuETI9t+Bm2jydiQlPcMYe5AAppxBQdzdP9XFijP7vQCfB5uMYXGjmNHSyAL
jgdEl001vqxqMrI8BApUf0kUHwHuilGG+SsC1HPfsiLEmGX8czJx9BGYE4ARXLIR
StGT4E6Olcddr0XokZXWGkuActYyzRik/XRLzaMug9TW2q6sr5CMLSpbnWkZvir9
ymaCYxlUkl190ujGGESWi6zCLiOC1sMeJ2bg4ySNWFvvnuZvRMP3hQoYJfRPnQ8n
/X2nSnM+wvsTWnfrfmH13CcqdHLotjiUKYbXdyYPER5WXiUylPUE6bCtGqIkG+FZ
clrTmFeUb6CNjZG+VVagHhUsodl6MXdLMIHuPIkFcjzIHBuXg6l5anIcLEIfQCat
PfYUUr8Uyi3KH+HVukRhNn6da4O7XC/nIbWs8yPwMDd/tkhtAOD1z/Lz7rw5rPtD
GctcQtx8eLbd4brdFOHB6Y0Ezx7g2h8fqAw45Gqoyj/OH1L7hCYov09Du+tFeOXV
cNJeNWdlzfwlDSW1O0rMTte9Ih8ywYPc8CHCZgKKwBHALkP/svL85llhe0GxsFzf
mVFF3pOMGRCRKh6GXJAgGoRZZZV2aJRhR9XMnNlQjU/7TAWhWnq3xj8kNU7FDULo
samw+dtCZziyms381TuYqN7qV5FnnO445IaZO8dXrtbbVrGNokwyBog0/UTEkQO2
3hghulpMoqTK/PNzc0ugInSjcJ4VZa27GcTTR5hAwZBcak//bfTCuhjtEqeu/NDl
NKUeDisny3hpJCGSy0A8OrWYiP1ohJUM7xwSM9Z/WY0SFd3hmLAQqDbAJwnIU9b4
eMWNIrf9k4TKlMRHcHbCKFRhrCbYWm24rdxuTRBMPoDCbfYyyf6D6715f4iMaMDK
YnBytseyjrmm1Cw9ZiFTNkDayM9Y3dqFcJNgaADSDM7pQy5p9E3oPbdrp0faKUgS
BrVNmu2G/04MCtacfnla2YNnI0ZX/425Nz+tDYnJXGOmvDh+nxCUEc2b0G0eG9ms
xjKcUbEgIqUjKJSm3d72qdJOaFWz5AkmcV4YEiz31nj31S7W+rc6AwiCdhG4CwTd
FriF/nv2O1fHAXz1o59yMpEO3IiL2nT9CLcynp89cNaM0dgwYe9tsmOzSiIB0zpx
/sUu2GpDdaJddSTHiPWhlH1Kc1gHMi8jorivQ3acdwyQ2Xk0z8vodQ7uFYZpma9o
spPDVgRFlLBD0D8YKI3AY5X/O4MAF03f1dkQx5raQBZJvGFMblPa3c1MtR7hzIZl
EL2D2yshVDRncsmAEpyAz1F6uTfKqgMbhRyuAZTbguJrW+iRVGhIMXOHn8tAicE/
FK8QP1NNB8f+zHWv/lqL8mphd0y/DpWTM9Ynu7Ovisd2KQ6TnO4YxTpp/q6XSvrN
5G3hAyDsBVUyBKXdvvP0+bXNvE67XsSy1yTmE2gEwdc2K/bhT6Ey6n/ZVQoEeHv2
TILa0saWdu+/dHYutLwOC562KMGvqWEufKffziG1Cb2rLMniBeVyAzlfSAR89qj9
yu5Qv7YMpybHdiHaG9TcyU3eow7al0LtlTM73clBMtxUX4B26zhgnLxzfJvfzdTc
TcR48j4kBlrxKTl4l2Xnzg7n/IhpCnPSbZ5RKgyoskCQDg0hORgCBonAalvAOH+Y
rugUMmER2Hf+XanYiML5HK1ADN8GEG7XnytOjHFAV+whLcnpZnQSwdn3tST/xlGw
mNI1VQ75e42Mx0s1ymDIT4lD8Akb9Hx5s3XVpa0+0X/Is+PnIs3N/6qNNN8L602M
nww13RUB5WBZvWnx6z1IndMK/f8m7gcP0VtW26LL93qdO9J2Hl0FVU762xf5i0QB
K0Zr8CTMKMKRAm6MSYpnZYbnrG1gplbDiAz5ck4hUzGtTsdcehnekklFcHRCIaz6
6Y/waj09rgyAMA8pDVaEAUqN858BPGy4UZYpzOkgisTxuxrhNAGm+PFau04Or2od
3T9ZQ4BviqfG1FDmj4u+kl0XIEZhm2H6DGvMdGdrmpfDwyETXlCPMuJ8RhFo34UU
z/wZWCbTfqnjlBnLcnN+t6QSjWS0Lju76wVoNj7KbNe4EPdmB8AgfasdorShYBv3
jhwtNn/Zlj2ZaMjejIhWktRHabLmgEPu7wpMR9hBBMLQwvcY/fIEpriUvD6l1/i8
VHZyi2LIWrVwLIXPybPYF6sx9hL+A6n6G5r523d6fs9XGiGOPcsotZGzdMFLn0sc
dD5zB4rUECdgv574gEhOJlEzdFVTTJdU5yLhdPAa4YyJXhzlxwL0IkzCN0oFboDA
aOayjKfFlMhR52UiLH3GPNJQcDLldbxdHuRoX1BTQKm0AzgQjz9/ffxi4TtuW5iE
EFSfVmqSoHOGGQx7/ZXk9ZbvUQ/+HLWHBFBduGu3YrbgMj8vRyeXvdHsWbTUoQTj
T2+5FJ9A8UOD3ZzWSGMeJR82quaR0EP4gfD9zEta7FcezHRBidTxcb2vBxSaRtj0
LYsDXXhnjMVAnCr7P1gNBT6SmIaip639p9DOfDMTOJfe8+2RcSeP1NuOVbXsSHQd
9Kp2jbJ2fFxD6VVt87waxJC5ioAwl8vCYFjAxkKNAYjQr94vwspp5eyNHDXfzn29
h7BQRFEtBFv8WN396b76y1GQ4pRLRtV0hHKwe/j5Z7FqFuUXJugPPw+7c8JVM0r6
yKtoTuiwdaOXEidcKUZAzk74sxpyko9KQPeGGBwak8EAJ/HlwqOEUJGoojQpCzBA
WS38WUXTIhcJI6cM1yL/xIVsypmALY9rD4RJ+uB4rRIdPS60RZw0hy+eAD4HJZVF
FVs3cprot5Lasea4gR/3tjphirW1arfDoxysDQyrYqlAZDK/oFuGtmCYY1Fggj21
BzMT/lHHE8CaXuxWiSVTR66Sg9h/mGjAYTcq4YtIpizqMV67Bap66Cb3HmTuWYeB
4xDLtIqsI6P3x3L5c91B+4G8QaxSzsQHnEVOLatcUKTx1zuV8dR8wdJFjv1su80t
gOXsAdkeklmV/HdybVIzg6Nvt4sD4V9f3mI6iVgvytQcbdMcpNvdAiHZocbrvrWu
wOOebehkB3IKOLOqUKdqoUiBukHDdD3c2CCzQgfve0SbhmKIEkn+rkNCjU6JwwYF
6CD2ACcVsBOubamiJL6Cz7IVaqQl0JkEQJwyxLVdym+BJaIztuPlMnhaCQpBOn8S
fRhwAoq13r5tOf0D1iJFlL6poF2nLCd+m9VznGTpHQUE2D1hk+rtKKM0M36fFY/V
v8XVIwrb53SRV3knNLM6/B1ldPYrZBPs37JI4XzN3FJ0x2q0RDYHV6BBcWsJiomW
VQkCNsIA/mHKUDkqRoYrSzPqip8bLAwn6QFtpmnHrSIoO+FdTftqFvbZ0aJdsKuy
ajeVfGnB4uDyvU31jzMe+iuYtYQchw9NWF1GLNVq8jMM9G4ZqwT59W+4qo+lpWB+
CYZfpE/mknnNjOU+eAdV8Glocy/67COUhlfCOm5o81eWkvUZyUxKhmzP3guvb+Ec
9PJQdoi1RdrVh0qLvtm1ipwUI5+eWKXT0m809QWkHxi0Qfy70i3VJezr9Qse/6Ae
WVAlzaWPoygEhsB0Q95aJv2/rFt/cnYcW48wo60vCuzVdFSCBAeXVYwUDtsGXEsQ
UXx4jdg2Z9PMV0KB/YJDZB8CEyEmLVFWnGp/NKofGDCCdCQ8hAxNRFotW3aUMbtk
znfLSI5L/xfY9LYznLtUSSBoMlQSKej42tgivp/1teUljgIu0xaxkAk+Z/Wf6JIK
dpNuACrQhk0CtQDAEo8LLHGeP3eX97S0dVIJkSsA8ScBZh+bSs1lR3KWL2gjFsqG
dUJ29PXzzLlAiJhrtJKMlBsaxb6VQ6J7tMN3zLwIN4ACOJStX0jO+87SB1kWEyWy
Y1K3Mel9sKYMABBTEB3S1rFcxNOqWY/s3vBI1VnNagIETkmaL3hNcGUPyoi6C7t8
yk5rAV+mwlTVG4H6j3RCPdQBC+R97NC98pZY+egRjgTy3bF3pc442fQFyTOFGgDL
LQvlfdDiQABaHDgy+Jmx/z+6WJQIhGoQkHOPPePowsS1RHlwpRo+0IZn0BeyrM7v
eWgP6jCJm+/hRuvGZuGcT1iKoiCOvLrQCwxV1HLGwHqFkj68EAs0K/Hz1IbrVJm1
G7ac9Tc/dO395YNzwBcdCqpMZsk6AXtd1B+Np4LGVzI10usLnBkOhXyT0Vf1zFBw
5rEECzAhplTh5Kj5Zdi/+YMY+KgizzXPqTm8LASZ9FwSOSTk5Kt+QdjF6ZtFzw/G
qVS4/xaS3t69S5TuzNaBEiBdnarfoR0V+Rsa0nf63W4UxiwJfpF8In2aUa8SQ8Au
gW0XLsg+IIW+fEEe/Xb5jT5vwFh4EDhELIpmjC//05X+9m+XzkiiwG50jzhhxDhk
qiuIJK6X+RedRdfZYk/KY+SeA7KeCspZfalrwWrJgV4acQhqWDlfQk2wdQ3lxyin
C0eAGXLpPOiGD2dvQCtCuKVakJ0QO0LELHQgD4Y3PRv7EqDmqQ9JTJNGSBMqkzir
F+D4B/RKdhMwuc9HoPoECCLWMMc9mKrT5+JTQFBFc60s5mIP/jLusUJyLzBs8F4Y
VdAEQgqxRplNQgyQwqihs4it4qxZU2XIwVgE9h1WfElG+ic5rhWKD17V4p17cvhX
ZMHqXEPS/vX588N6O42Wmh/TrM2yrr1rWYfO7GatTF/b2xxpppD2Sqtpz7pGbYlW
DYeUJm/lSkP80or3TN4BrHmoWoDIVUI7y0cGuxn0YB9VYJ7Vdym4Lv4m9LHPuBzh
i+D7ByMFRVKpdRmrEpjYv4G999LD8UT8v0RKOkRuh+EIzQdpHRs+ucpToPoLIrMK
A4s17+G2EcPIkBmQUZC7uLONx+46AMpM3KaY2YuF4Nu3Yh9ge0xq+ggavNoNAuqW
3qfoAy7rI2yXERDd54NNKxNWuZ+y3btjhED92kRe8Ti947dus6J+Ijh+Ltly6mJn
3n+PQLAVRsGOTsc6IXa1mNCIWdPNw2gWdKbkaVAJfM8rqe9wxhUsF1lYibQ/qV2+
hxrHwdSAtGAjI0Ypmlir3WqkNX7vGOrUadgNQy1GVGxkWNVj4dGQrRa3roVQOOmU
2Cxh1x4v271H4wcT3ryXe3XzBkIDxID6U32uMpVEbehDF2IL6bCfCBb6C9AMme9A
yp7FCboFLe2BiNEhsSnpcZ2Yu28Bkrs234dQFx1h2x56uDphAAlzUYbUAgdewxTU
zTC7QDsUH6bir6Ic4YqP0xSyN/TsueGRJiQehf9hNCGkNg0E9ypKeadJQw2mr3aA
XD5h2uQOt7U+Vwv1CaYjBw2ySWdPZvJXdzJQZm1MFvubXQ2eXc5UEVMo7bbnZV+f
hmt0jREL8OH/S0QfE7pWa7FoN7ImH+9kZJBvwSek5hQPRSIk2HJKhrUt4VIeOB9F
FxNwJehhe4VTYMv7ZYZZay3cCn6A8r0/y6QWXgaYNZiBxlDmZ8G3+Ul53c+ilxtf
91MQ1gU/U305H5mCAA8rrW2N8pmQJgtKbkDg6T2tVTmezTnpFBHso/5zmjtJOcEj
AlU7UnpVKE68Kr+5NZsS7e1scIP1WFdPlXDIv7fQOlnhdogTUAuXJQzdfakeXnij
t5SoxHbbYoOcenQgR9Xe/8QxvNHg64gk5kn2Zo4kuYwR+I87MhFbclH+Zk3gfBkG
chWw7zSaK9Aw3cyeid9dZx7gm7b6EXEOoBW3fi8aAngdQoMRySGnfLnGa7k3e+gT
TQ+ZkaKOz1C3yNngEwI6oUiSLZQkmQ77Mka+WOuPS2G+DEQgWoZPNHsjcJ99btoo
Tgms5aQHurMc/RqSODLB2CkbAVNk2VlAYngn4G91eLpVzuKdxBhZ4D8PyTxltaqS
1fEXLR3olfO1LFdmhqPGX1YHVDUm6eB8+nOgJl7VSYeSa6d1JaLZ3pBmcpsjgXvY
sv9ac+Alkx0p65oEiKSuFJGoYHDlA57uN5yrJMBJo3ZUkuuvGbW390Ic53lXTTa+
0nr8RrVWyCW04I7ZD0PPUDRGiPA3dKxcgdWp0d2LdCA69Bs7Q2RuVAEJm6ehqssS
XtGBv13/MQxr689q+0hidn6hRRXcybHzqpZbMi8CE5MYjvzDqqGAJnKOqOSzvQ6+
cDOQnEJtOkbJDn8In4dCeQi38VucYmkFkxwl4mjb4tuWjmBA/ZM+SIYT++zjC03O
+3iLnOH2E5EGagLIFWrE3qommJ0zEAlR0+tJVF87Q8wHKFcx1jxxrfpeB3Y1zsCS
W+JbNFJGVcIrEZAag2X17X77GQqoK3Ye+q2xCnOcWnVil/1cX+h9THmEvlsL1zrc
/aIyqqfSVfhAowpAhkBciL1rVbtPLx2hdG7ZHMrGs9icwhEYiBVPFp7XJfuyQjrL
XCpIcOWOmk+9TIrtV8gqvNXFaxr7LFuev5Zkouu6vhdpvabTVFYXawuS0bfzOu1i
PBN4whceA5/dd2qjhb45Lvn8FKBuW8oWnvo9Tbq5Sq56J32llI1Vo82UlfwT+M0+
p0sTXFcDx4vZid+SJJ6zc8Ls2JNIABCCIkAh5e5lq6VXY7TW9Te9noDPySmhLh5f
NyoK6V7D7/3/mwOLWJZjDEL6Gy2DXMhmx268RMClkHvVcAgw3ZkTWeOva13m8dPM
X6d+aw4/ZXehRxU4ZhPkVrYPlYdnGmLp+oLQjSHbgVaS9Y4NU2uMB4eYCNt8VU0u
o3eOhGcUkStE3qbdatulx1Unmo4nLekXwl0/mEW831JbhdznHisq7ahThlw7UwoT
RaoQBe6qaeyYPpQt1Z6MAWsXx0NlTjT2D5gPK/Ip8Kp0XDryPLsGQ6Fu9DTkjDzq
ZaMYMKC3cRkjxYAdZTBki3MdOZx57bPyLPHgkeDjTxdAYQ9sTmm4zrKganZFQf1o
EikBFBFtsPkDuSjKRVj3gxMc046CEAVw2Qiq2L1dUBNY1PYsZNGF79c+EBVRdut7
/NU58RzvfwC6zCG3ZvlBJAz2OMsvXatT/ma9Xe1twPU3zAHuxloVRxcFbAYkxJ0A
gBM8dPLz/rt8DPGP348DNaAxQykIvLmoSuUBmChCkpmmmuwtVnjf0AKpNazzZKQI
vAaTN1tA572PY9TobaSb+r5y/lP+xVeDnAt5yvprYiPQ7vYiicozjutLInbN0Yal
TpHd+QKB9EML8lM3q/UJexqXqNpj4+xh25YM8737oP4RwlcZVUIN/4cB1qFdRpp0
JrZlhn2GUdaC75oIzpmeKL1zxk9+q7hQ6ywANMdiC1Mx0WtrK1uY2Pf36+mgJqqR
CiXbR2hKGq4Sq++H2jkBIfubvi58bZ2Eu/NKpCpTnYRmxeFzJJaBKKw7hFP8PVdB
hBUYAWrINc1uCAp16/Wh1e2N77h1BDs7M+ENu2TH4BREAgmhnm9fkm03siPJaFg4
sEUIJzHgqAvS/MYd7ZgWwvuWpDGdIo+t44NBZ/diL7uoPyZuGFwwtyYumvDv+Byu
XoxnKkv7RSJaRWszWBiBoB+i/W3JY2WixP4mvw6YELUa4pFMECNNnV3gRz61bob4
f7XUknBfqiDqmCuWB6uFA3pJ9VuShJ8nU1ocRboRoK3/c3K1BgfXsQpL844qUMby
4GwxalRXOknAMArxlaj8VYipzzBwXnzOqxSoslhNPAEQYsvHzbiJaqGoAE3ghu3k
9ooT1jLy9PdrN9LkfY5P6tAZ2ajSAvarS0g8clNi3QRNQqB5T21hrbtLnUUVt+ez
KaCcHYZng+RhCq+TIuLvnYrKP5l4MxHVuuOpEDGFZr0NZGtiWFhqMsHlxDI63uBh
kChm6v8htvxzU//Q40Gm8eONg2sTJP9SOaswmLlgBji4jWA+uwwPskrs1s0mSmxO
Ab3OxVPu9v/nu8eBBg/j11NPAPUKB35XBngm1CEF+L6U9KBrTYROsalZnyKUBTH+
1hoK18mc8PncYQFSIIiYCo99qaqZix8ZqPA/pTLzv3Rdmaz0c4JcSjsX2LY6+GmE
7VE50IhqoOk2ZOdIOu0Irk+mN2P1ianiMV+SdaH/rMB2N32korvymuC8XZdMPmXY
6YeZ49pt49Z4gzc69GF58PUGwfP/D11rkoLiDeFCxXmbO+oj5fLGG443hIPPmsDJ
96hZj3FoG2QNjLIN/drlXcgUZVjFS+GwkErx7pEm1Krm+AFGA6Qt9Xq+2CITcUxR
v7sEAgQ45XW4rqZhZEQ6CZeldwnh8mpB9km8DAivreIq8A2hzYWoHNJOliZMfG56
Lqvucs89R+dCNPrp17U49Eh+4FjpFRy6nNVgjtBfQNdZrTdzb7itm+aoNo+GKXlQ
arx638RWpFkzeLA0BzOZ+OBbaBQ27KHhQIl3xKB0p64B8vH6N8w7+vkUHkOZ7NgU
5AQVoKbKLlVilqbsrZq+RHQqZQhI3DItswlKdBu0emFdoXOtqFtwufbus/7tAiRK
JwMi4Q50MM9vayL7e4jXYS10iybxucciQie/L/Cjhm/MApWgE4lQkcFZLpZ6/M4F
ovYNjGWj/TJCq/xnBmuxRHM1NhcsfU5+71sadxo17qvuh7aVFoLfJ1d8KnyiyAFC
k2u5hy4xnABYBqifOmBTgsW8V+QNUmpJzWZm2QZQF0pPrn7qsaY3I/Etc4NLiRMu
OVuMG9hZ6UXS6BacguH2nh0amclmGyFeixLEH7MK/pdtzy0nEBaiRP3Y+hhi8e4Z
OgSYBW5OTkZm+KOX7vlIIPMb26aDedWCCkyGgOYk+SQXFzXP34+5F39NgxNI25X7
yjmFHThvFvnwnpIpgIU4GO8oqCTzElAi869swaOCzAACXhKe5aZuwZon/jYHlLvS
i5kloaNTdRoW0Yih3iAuUfznH/7rsp9XkuDeQOZQ+elIsvs8vNRVS0IQNoZaW3AR
v6qssLfb2VoJYWfrgXA4wiKCDFwASKSKIkFWhZcK1PqGZ/h8i5PHMy0eN4AW1uYA
Ed7QAmV1PdQPW4ZpHqHb3gevR8bTRlxE6oW0CFKYqC+SGyc2w7cSw3eFF/EzcwD+
dUt0QoVJlmU6lH0fEx+FqAV92cqhGQus9+1dVUUY6vwnqbaY9K9ZBVhPRDyHxgMX
8mSbTGyluvzxy/+M5rWL1XQ9f+Y7UYF5wGch2kNScBXqdjJJXETHX6jxMcVw96J/
Zf7ickt6lY+FlPE3c9WGEWp9gR2PtuwI7/rC2iQI4fwKB4DMVgGNlJLQCvkN8YVo
6VKXeA7vRB7zkkmzpxl26LlnK4VptmJcODCL8D6zROupx29Wm+F2TA9aaqqorYkV
beXmcr1MvZEWb2K6bXwm6UukolYakE1tnL36PTD1vZw0snmBQF8kbkX9a5j+yv/3
K8FnBaVmLGESU9aXBhHjgSvcfJiqOuJ2m8RYQdqcsU+TFnsHpi9I34r1WCKHzXTH
gyOUTgSbBrAVg9pfox6AETbcDU2zqjUbZZpieKK7HjFgKQvoEFRJtp8VjlPcKRpD
WBqYXoYlEgroxQfKiNGe7C8ByFVBA2lCd+cskcnf4y1TRBKrNkDg+49ojfIFUJxl
vvGLrB2T/mpKSO4GZYeS5+Dk7Ze0WSkzjvoRy1Fdvt39RthS8JLdvE58Rg1FOniO
+tjEf+s9UPaE9wQOVvDejEU/nEoCHc5FL/OSFbI/3OIfDXq2cYZThlQxkt02fqi5
9V/7BCnjit68D0J7d2Px6AU+iOGpsn/gAzrxndluKEODfrz/gaBQ9N+MRzqNFFRu
ICJ/+qSDTTd88QondMmJPbwt4yNUcP0sbCJo+IrzLcMhbXOqZU0hBjAP9/DY8Emk
GTadBgUXsL+uEcJcVI6xt9SctYEckg/23OiDyHyK1G+G+biloVdqnaeLUw9rfArG
SZI49j7Np0uCirRPcUQhDqWeUdODxK87CpTMlM2zmG7eYbr5jQ1T+lXpeeWrJRsT
7I5hEJhVTFnquT360t1gQ+ftTYJqnqjXvdaCkfFYXCJNMxS9+nLLBUtW/lkXqsfx
oSoGMWuieBrYCQuu8Cu8bzJs8HznqhW0fOWBPSBcmfYpL99VV7kOVE6LWe4uVCvh
rOtcifTp2HSQ2W6yxrKuIuvEI8I2E4FTFnIfqlreJi3NsfR9HleY7+pDP4gyAuEL
jOnFHLmMPIxqztvKbRvShJ2wIEecYsigzNCj8u1OE6LkdH/nUiSatm5v/3tfs2Ip
nBdU7XoAZ86MsgCv0PIejFnXvfs28kvZKNLpLhB3aFe5LZW1RddmffeByBVT/Gqr
jMSeAgd5G0gMBvaOE0q8tqksXAI8aSOPrqdXMQwx7JiuEo8pRB0eK6NZPWmaDtxl
HkC4DXtOe0SMapVH+1VYxoQVbkL+REjarbVy3gY1UnJtVAd2WMIs7hWIdc0HXlmM
Fv8OdDM4SJqdYcI6cnUGnKpjhTTaBJVJ9xE+bDn6LOBACbpgUSVrPQV6/yrJ9s0+
REEu6iiO5Ge8lD/rPKZiJh4y4vOe8ky2FQ4Z0KXRyP19jguYSeS9iHkPM2tTUw/5
WyTdT4v0sDDZXx8L7FBYK5XAeKMs8AxY7XnIhPT8p8gj8hEoiXs3YBAnmjfyy4cb
takpGsTLI+Qj9a++v7OqrG7fjQ+f61w7YDQaXhZfJgsxfv3QNxRoeGcUY6BzogHS
Z4potASZUbIF5M2VtsSCJYySMu8oq/auASVquTVNJmwsm6HM/7z3Rpa5XS+VkYJg
jsOwzJ8qA8cRb2qHitYpTsBeuhcPkagHormlJ4vhl3zjRg6ZeMl8GWtK3rrDtLUO
rIakVRQ24De68c18h8r9snRqZzXDMRYpVUHi9AkFpI3Kq5TTtlg9i9JkqORU+l2L
0NR1bSJmlWlCTyoBPaJ89kqYoVMXTEAbwbjnquzVshT5pdjqh4UMxw1pRwwOJ3hg
htJAMYV/WVEpxWvFGHNSahrLGM5IT7RKcNyVx4RNK5bxMtgGeQkJgDmSmzmvudCS
HJB3CL4c76hNNKTveIZUaRTJ61AxSR+k5Sk9iN4E4uUjYTRotAcfXNJ+v9VV/Wr+
AN/1H7R4ULePn3LygmzTuxl31UQQd4t+2wCb5G0Wf/XVD1e0X0hKnsiKIfqtT0hM
qCXKfZmeZ4jlk6fhw3K4vMewNdSHar5p75bFUcM0B3FlDL/RJwa2zpd/9yUwYaH1
sLF6KP4Hbjbao9Ugi5uztQujir8rIjVwclxkT/5kxZz9CnT81xExd0MPMmy2FerO
BHD0ywu8w9K+XBotTIsWV+3+I9o+ZN5Mfcw8NEN1ooBtoojh0pCaXw1Sko17WkDV
sCGk7XEyM6Mo0W2B6w/HBk1TyZcYw6nnZ/B0/1EB+DX0hQZOacUPlm2KSgwGtTCi
Res4JY5VQjIZGyW6fO8ZcvuFPpM3KpT2RWNPYcDO+Yhugt6X/BX7EgcDao4OJS0h
QGfPtxjSp+Z+oOJMES9QS/6Mhq5YM3Jj1IWi2B2k230uZ8TIK6zQ7uVVdDqV5mbQ
9iMXIxsyp1Ir1mpKHZFXd9LivFGFFQ+J+rchWsKhj6aj5+pQRHUhk1DBPQ6IdCv3
okD/sBEylymmG/haGqXC9U73wW50YVzqW4nGYlIjiqIdxhfXPJTPzXHvDjLVvbKb
rt5vD1gzQLakXLdtXBq7jIuCi5ZB4awor9tf3WuJ/0BVxMTbeuuh6OBtJ6msAT6N
Qr1bVqDIlgtWv6M4NB61asmiHp9hPGd5FY7wSh6wEO4wIoexvRFbVjGD68XNgsDf
+ol87CTvAvlVI8bCPLL6vVhFUJMYy2E+NPi5wrWL6XLXdE6U+H1RTRVIBYtr0Mr9
LJVeaow8mDAd8eOSnzFudClnqxPyU+SPvAlKUBmlEqKj+5/n97FSPcYfzDYc4hY+
ivs3B4lLg/PI29APG7rlGsGaS/eD6dUZXVYkUS7dDLruW/lMLqOTHxrkZvVcTWzw
TB7lPIpfyv182t/dbfbtWqR5uCPlosdszLDoYztk3WZ3uFNpzO/K9CTlsiFCchU6
Q6KbRg8oRpGZ3Fd837y8IP3tYXroJeLtlLYJ5UIzoL1SBddsF6xgNxLoAwX1PYKV
to/rSJ4MYtCk9FQIZr/ZPop5B3cSyHOrMDCE69W43ObHvspsWXV8w3jNKgzbna5E
PiRLNTz4fnecqQSSxSdBLKcoSZI5y4fffD6QDnC764GufRbgPD9/t/9e5AbNwPLY
5W4T4YaSKHLJgeHFyroWm1VLIYnZcTkfPzXWmJNSOV4HpgzFe7/2AuzpkMzrQi3n
lQpJSnYvMjEMChReCnMg5Z6keapSnDXLiNv1zg4SnQ7JrD57z4k/qj1VQhHff+4Q
P0x/6bqT0TC2C2DUZhQfTIz4ElophHaNoX7jcqaMdZuDm01voO4aG53BHSwzVRf3
lv//eyH5WGYElyV4naaTvK36n+0cyjBgaCk4htxdqrM/5JA68NhpFZfcJNL052pd
ZrSazjPLU+8ZTaf7iBrULh/yA7fzIO8uXV4HDD3N/ivYt0P5oS6wad7Uv26jCExU
KtrTGV9oXUdChztyDkLRReAVf5yimkf59+RyUGa8mS1+ENB8ioOZAM+5Bund48OL
GiOtQ/YhqkrZX1R3P7J1tH7zpU9S+GCvafJlgMf8blpSHPDnFAHkbX83d3Yh4RlB
nrLqGKKzTW4zyWSIYsyWktXH24at7AqUVgh2vpqpkhy+dVWytlefUAvlWaGORiad
hR9RxHE9CFl9jCwJUyzJMbeyQl8pyg2PRj/crNksPDzwO8c2bTS/9HpPKgHQDiIt
1BDI7GaHBFngGC7Ozwh4fohg6b8MohDbJIaavrB8UsopPZLyaxOpmcLTxiFU+bis
zFUd0IijCNBj4QQMSSj/xw50Twg1/Dmo7wQtCZhWAEcvUn+6kxyBdie/ifLAyDAW
uZRk3ee8ikPDJ9eaQVgimY1/t8C8SkFLQDfIubWtHG42iePnMGlnDFLi694Y0cA9
0/nwbqHu8UESbjMOdgwuYz1hodsFre77gpBjkeTBid8RjSP/2oiuSV4p3fHIWrj5
5wRg0eAe0mK520QZGlu5OJqLswuQr8jv19GioJ2ihUe3lWQpWva5p/SFzuMeWImp
1SnjD0NdYtFB1t7BnOh+O07RKXRUhhFXhV/V7rcWmvsvuiqEmtnPXUQ2SG2d4jnp
xCcIUtL347FJTQlHtAyHzgH2gKyiuf9iirOAzCNr5kXK+tMJPpDb93fFt/1quPW1
v8EWEu5kwnhn2EqbQNlzx70MKexshhIVK7wyGcOqAyUK7JpXbgg1uT8ukHCrZYM2
54pT5hzTt9+4y0Uajskm/Bf9v0J0UabwnF2k+TvV0CgF739yhcNPhdfK9UYHkax6
TvBKtPNTlQomoONyr8xPRuaA/towypxpIN8LZBemfDq36OMUHPSVf7lk8agQUkie
L4K/ZeClKlL1dt3f5fgsN5GBSnRQCAMig6GnA1CH1DVIa7VDAFGF+cdmraEauOBf
ynsdoW00CvsY5h3SM44HugkZ4605oCJyFu6aX40eymP8M+bgBEx7v34WzjatyiE1
lyrzuR1nWujxhnc/8unJvzhzIaEBjQYk7U5YZOgh9YC+sG320fMO0sp5lBamDSQK
zAnC6gHQ8FQpOCKZuBEShvtRloi4SZRat0bKb8DE7Pmeebp2QRN9QEqr+90G3GhC
J7byhuTA1oGw3Rlz20MxLxxokgA1sn7aWKWd3pzy4NRLUQBYhfXiTI+LYnztyQfi
7hVGEHJ5Y5rORo/3QKV+gHL8PLcnU1banRbwM9Jg48bWFqBkgkrTiCNgyLef4seo
chMQ/e50/DSZZFwe8/qGKG4ZMs7cPh14q0Zaxzh3yC9TGlUwVDL3R377Rdtv3Rxu
9g+KMb1+233a4vWEdXUc/l5Pu/bVhGbdlpvQKXQKtRSCGqyAAO0QgsKCeBgcoE2T
iL1aCW3vOCTbJMatn86kwHgRncF9ohsKmcetyVI6irlJEiWFw6ULjOc3Ks0/+z5A
miIsuODiz/xAnChRDyN58IY1blGwqp0NznKj1p5bU3KYc0XI1cbMgDN6T+9PmhxK
QuUcoNoAH01uiZKjbCaQnH2LDoT+GzCgrot/Sge6crW7HfgaNwGrRWi8Kqzyrgby
4KdNa+1k6wHuV+CoQ9sjhnuT+DXOiKM2GckV6dbXMe9/Lpxse9N91Tes5OALRgFG
b8ZasfYD3TSk5utNWE7KyldFwT5UWF+cIZhwSHXc5D5dklu/yRCAZJpHatD9iPTg
SleUS53hf4ZZ2w1vZC+3RTEBXsARpa4Z1GcahouACvNiPfHjB8DtuYkLELDTfLGl
lOCk40/EfMC7ereVo9K/IjZcPxwtTtRjQh4C6GjLHn5w13eJPFj8W2f0iwM9TGTQ
Xt6wOqg5rjReQEs9wEcyX/37HQWG/Z2w2YkfetFIsgEYTkIoJOze7UP3jwwk5q5c
c1YKQpbVfzifbe0EWhFU3kaltNnlqxA+BQDn0Wpcopn1SLd0cJw+ZGAIyMcl1nlj
X8FsJmGmlPKy5Bs0QoUfeIDqeUZRBv2xqpgouYAkdiNmrIcx7bkSgfxdeqUDb2mf
9x5wcqPf/4j/SIJl3jxaEi9L6pf5NUOn7af2jbf6dbD1b+egXNsIDK41opY4SWT9
AOVg7798NYmJq7gD/gu5H5N/GBwfpsgxhz0M4TH2K8y27OezVQ8vfZCx/7i45AvL
iQ+HS4jfomv5sOsy5OREiJTdHVOLlJBUWWOYpFeW5IQ/rCMKkT67VRGffBvxm7z8
Ja5Fxox1awPl9AIzMb5OSbDJpexNBk9iZAr1izUZWDg/j2OQfd9IFV63m1OU8dHj
grWb1KYhlj4fwyDIVkuzD4MV+UCCXl53hF3dgdnv80u7pB+ptuRrqQrNQICiRYCb
a/ec12JwAriJftJHS1m1kBroZoESFicvOzEmcHzPDtaOHMHp5E36w0QgT24LNgF7
f/RQEqpcumABRzcOGhs7rj+JK3zzzqLwq/NhEHdzuOaOC2Gdw+FrjJBcc5HPCiXf
o63KubwW+r3F1PsuEhZneCgc0ceKZja6FlAyo9NX7PkQ5kQwh0YdfieXmAq5BqKA
eUOlzkobEx+2e1mDFQ4B+Dqq7uqGcyeE7BnmvxYutRUah503M2haBiNa1kdkCsNi
Vi8Dwoi4/iwYeOjG2lWwDIcp83ZewU+Hy7Juxlnci5iWeVV0NDktRry91pMcCyFA
n8eHQ4FpyCZsxEG45Yh0d4Xa92Z02cobasQThzA1S/MxWN5vK7D/AaYE+07okZZX
YTbqltpWHkivutuPv9MRQhnDX68IbSD6dhaBpq6IHWC0enI4fvMZFMX9s3Yr6BXP
VseU4nOQUbJ03Q854jOBVCYwUZQp6BIHpnazBxxOe0CwBiu8UyTTIIohRNJCwAhZ
RtITmeXC/5FdVaKdh/HAfcesMj8GLRDRip3TwCVyPN6YXMZgArCiZSUYeOybjixr
oYyDjMrd+p+mabcP4lxtb7PoztiPl3u74nod8N6i4dMkeT66SL88HYfClCBeDTUm
EHxwOygMhw3Kz+pGk48Zk9lUlE7ZgfViRrKnsj8CKccDfj/6XXMqfEmhcB2IQzMh
VPl6VBxmjLVXCFxQwTG4rYGN/E0wgL1I6qLh4IDt1K2V1EUiIyhZgwX0P+wWF8Oj
V5TXuFfUmqlDKdiCjIOqQ5tPKPFSDXKjeOBZqdniw60QCH+GL5vCGefcwa//IOFH
vZ2lROh/4sYyXaJy9l3QHli2RtzGI2xg4D0BTwZ8Nk3yCxUphK1N0h5Ki/Uxa2XS
1miwmgAahkXJ4zom/ciIepiU6jxs1qGc1RoEAbNmwjzFSQHNy1RSpiLxb8IJ0PnV
pJuDREnIZIPC7rRNyflLCwXJ1l1vFq3a39B5rY3g3jvNTw/UHmF/XGwTJx3P3uGn
eQCGPFewHUMqqT1Ci4/Zp1GH+bo7o19RQygqL4wfbhEupL4urY4KRrNlf7f0hakW
BQA0oDL7CHknOVS07OQbmWN8eKdfJwdCuXNvjFG/UdOB+MfkHz7LewTRjy+bpP7L
036mQwLGxIvMp/lILUt2DTIZkcLej9ULhSpJ5vM3t4WiklvVZjekiY6ElYqzB908
ZTabOnB0N9Jpr+9sgitwvpKAJG3xQpnKhR1HWv6imqBnPSDO0wh6KBnSz+r6ctdo
hskwgt5drUR99nmeMsLcJWKjl3qm5Zj0hrv+iqV378cuBa84mLSbCk9E/5xFh0uU
KU8vqPoveQCtk54WIlWcn7C+8WIwsMK8RzaAfaj464cyURsEDFDuVEOXBcSDkSp7
JNS5gyWE1NVhQNR7L7ZoCnmZVElXabEZ5J5//kke2ZGRA1RWv+RSTbarix8Wlnms
swXNleQ76DhvAqQxDFs8Ch4rLplSh6RlEpxGFUCLQgSMucsNbyaJawKimLlpUmZK
uQWp2IypvXhR/DynDKg/nYywOK6beGYteMvyGehC4dFHmJrVk99WPPK5DNc9XWE+
tyFjzPa88FvlCLHpZ1hJsTVuPzFt1SaEgOre8WVZwRY+myrr2rusrpjo1qsYkhvy
JxooeIEzWb+eNW2zmquszd3yHMZyGYDLFtmMLfj0CckTjwHZElhC06+jGpaYwBry
08y+vO+ozadLCquT9+W3U5Ajpoj71wbbzeRApFkKSPyCx3TpcnqXFWbvwBATaU64
etOIc1RqD9JRuxBNBPaORH9UxSBRU/37b/r0GsLkehgqeQgKGTGWDwaQ1q0QnCr/
3e89gq9xSJcfTCwJkM7ifxQsv8ga/WXYFLZxWBH2Tx9m/9CE1L8uwWq8FeY6c+Ng
4yLV3VHT4/0K2anH8qfS0CheeNOxnBBEdbuAIQt9IKcvV1xJJT5cmln72lXQeb7w
pVreDi5XCyV/7oPVr8Hib+Jq2YLhgPu2qPK5nAfPsITkKV+0wqkEXNbjnp31NwVM
XNNP58xxgfcnrH+C/ZDr07KR4aaXhAQTdBX+Dsm0dwKTvLE6nvWMelitB5940AA9
7PqhyQnrPa34UPOSmGVhozukL8uVVn4bNiE6txUenCTAsY37p1vrZCmwftpMaFn7
X7+T4fVxkI9ydvlZBm3GtO8VgZsjUfivS1Ez8xbALeivKsi2ALtO2JvKO+vivgPj
fcLAY1ws/EkOYeWUt6WZ2QJDHLonTkgPjUFCsJP7sZ/Dze94vOBba39eYx0iAp93
KI+PY0R83EM9ElCK9T4HoDg/q9k6yBbirc1DPrRKLio8ExXjF2IMyFmEavHEUk4f
IX3NxyLp0qo36mwRZxGVLZkVN0nCYDg2BhMCEcKNBorMRJGiulvtIRAiXP2fkTFc
bYzzYMvM+CuQXcehE5WzxJ/DqZHKwo6dbvaaOIHXiQYutkOtAfnhI983frFvmjIF
z55g6n0i1XIszHTzsDEEUXapIAAHqnb7BjR5CyuhmxFUr6E947CH2vhgclzQFzVs
5impyXlKKCjW/u1m/tqsP82XJ3f3THVoZ0FhsdZbXqEKWzTWrlC7ABrarTkGD8DP
Pa3jPusQSvH6+RX1qqKrehXdgraPWkqyS/jS6lYZrd4LLPO0dop2t/9PxViC9MDO
V/MYUuOorXLSVw0Z5CgwiOlYPHLNy7WFthDw7gjMTAG4YgTbmjaHtxe0eDumnELn
SS3mZJuaLf+i2flh3ghxgQitxumVElYl/CIELiTI6fGoR+9XLV49Ry2aktYaqVPp
3YkzACN2pW0OFZ25ldI8haKhTSs9MZMqavahA3HbMRflcMIZzctBG3iIWw2Q1R3u
djENjdBaR1pJ3HUtwgxpQKEe4QOjqPJTBooyclxA/Vuqkv0Cijouj5lo/y2FbXHN
6vpA5Pa+ltQNlrbacOxuCvM1Wqvfy5KJCUSjiKi63iEoaR5Yqs5XfOVLrBEofN+Q
xR+5pCXU2rlaqic10rrkTbiyWSMeGN/iZa3Vut9PuAEqy41CIAVXxUeQSNnVAe/Z
9pI0Ml5DV3B473kq7OkJBUpXVGuwx4w7uSFNaB3WksWy350Jiyu/Va8o4GbF3Ki4
iPizNg0VtQx8c/MX6z4y2x5d3ogIgWK2i+WAHIT/LifXSAJDU9J7JTW/eZsoZoHR
fCsT1e/OpMJtV0y0u1Zd/cR5ScjKQgu3hjKd7GQH07FQr8N5Q6HDfc54v7MfcY4O
HuttfP262zEP5onUIKXt9Vib0MdlKynsC0yIMkw/PjR/YQnfhmm3POkq5nsjDa9r
6dOGAI1Gom6OVxkGd+jYCwkNr7bgfXhQs95GhPYjdr6x9wp3d0F0M8HrAJ+Ix739
v9mq808vPwTnaJyhiLepRuZW4jycDF8pDPjSVEyPP0IYcoVB9hbsiwQfdRks4ABa
eyT0QkTO4AXkecN0EwzMAs8+JI/SxyN+v3jDZvMRzCv5eI5szqeao46rwUkPIgiq
Inx/nC9hTDlqDSh5vpuEVciCbE0WTgW7pX1o8XaqxdxgmUI3MWj+30xfp4ocz9+c
sLN3EUHeh40eOpDbGlZfutYCYsSDEoDklrBOrQkFNu/PLjWI62pmceoVDHcrGwx1
uThmKurYjg9Nhkq5VXGk0TlSe2THFdIg1XSfRZ9c0ogsq/1KjN2LzYZS+SFRufI+
RnviNgnJpvjqGV31ExSh6akZw8iiOEBgOCmm29240bDxo4GjnSC5bQIeZLlcNPDU
3ovExikivKBYrL35n/qwFoYIko26lbmIRbK1Dbpk1dNzaxsKPqs5gu0Ba0xQleY7
GrHouJJIdMvPl+rmKmXj57fhpIZeN1q3VdbBykIw0ppckrIxq/AeU5sL6KTjQUvc
WmY+7gj40/Y9mMpIYmx4b/uVXF/wpMSjiWUVe/V32eDxFup5gCqvV+xYmqHFbgDE
EVY3Rm+xO5Xu1GJyhCyCAti/8/+8KtwzmacxDcGTSKQFwEUMFdcGqszN0adNSp9U
aGDC4nBLcYggrt99GZHzHOelG38w8yMfxze/czioWUvxt3gzQ2w9Nlt+dngj9GAi
eAM60E77rpVJrHn1fKpzHhBIIfPoShk2a3MpK8viElVPClEOyK+nvGz48gBAbksF
Ny2k+Htkj2blkVblNcskKqAwRank6Ks4gAM4FgXrxpjT8m7Hj8aGtdVadc3NLuMn
LguA2nrdCzhVePASBZsEzwPTQxMZd4YjPSCjLR1YXzN/Oj89KKT0DGZnv5r5mQxW
Yggddb2CTdNmRp2Fk0H8Ke+VFTnTl7T1xk7qzeuB0kyK5hzszaNHWvNjDxsc4uyz
6hXGI2H+n7kCTuFa0DapOkT880teyKWOYrxwT3eQTuxv+XrOYCLxN205EwrCJiDy
4d9jJeNpi1j7lBlq1YpqdtqXTK9wfVzgnWkMfUf3qOwDoxP6wV1O+NVO59vKHAd+
TtiQjt+yMsgt0zs/eWsTXoRPZ9H0HfDOhe88BvdLT7IuJNGBBflKQH3QekmBkxTB
0nr75jGwYM7ycKGAMb4hH9C6wwz32vHxBcVd0InWomBtXEWj2eUxec+o+lq14TLj
9HtDzZDFEIDqLeB1lVssv1og+x6oixhBj9y6mrjhWzgMjm4GUNPaXH51Wnkw6pUJ
NdkmtgjukJlNLSaC39h70q+EVi0OTE9594ah8EI8rcu4q3iElfIZdpNl1u5fP5DN
xOcYTZzclSPN3CEE8HEX77O15BVdcgqP0wtqb7MOnMuVQ/5jexOVIlyFOnTuiwmz
hpUrlrJTDljaHBK3gzQ2haFxJaLnIqY/9uKsS9fNzE/lpr4hNlZhnpgOJyidfI3p
wHhwzJT7VJ9GuYw4ypiUFUnFE+urtPjl6OOODL7aOjRACeBBg8h1GsXie1i0Yprs
4cjnONceQBUtHErv7pYv4rgcEe6bM36jCSmMTezo9YnZQAYnxwy7jkVIuZ2gxmQE
qBA8ChCjtcwEtCt1TFxMXnCjxizXbjLnIBPRsUX9u6nyXt0JdDFNu3iBWFfa4R/q
9aeQ67gQkl4qMzekLSUPbtrpXUK3sVDx/EVAziXGHqhKbc5r38SmPUIjIuDea40T
Go8voDVMPtAYFoOAGHwLAQWkovJiJcvBEApooz8iwnsTI85T/cQnHTHj9NpLr1fz
NXRFdYA0pznQxSAIUmiiJBD/3EDjxL/9VfPfSARIqnMalxIjcEo1boa70/TDtA/n
UwezANShmvYFa6CP3DVMfYxF0RAY+P26cTKTEzcEYzIzbd1hz+KVrDJ3NQUWfelE
nWmNz+OQxZCH9ZVXpCVmN91C2LGT0gbFr1K15I60ApNu5QwDPlnsXuewieRyIyxe
Bkjs2HyZ9tl4vjfTJ2Q0XxK7c2EkxG6xIycnFLGK0nbo8SodzWhd/iNTWZESe0nO
LPhxxfIlB3yjwxdIXjRLnJfT6+CSIGplpXXLVFNn/3h4stfqGkrv+/v6ufTEGEgN
mVSvCm6Wn2jlpEbXG0Ydx1jARXfUv8iy3K7r2MeKJbiJGipd/xjIyrwVRZYrB5lv
LAXX858U9nFpL7X60ty8dFIG98xfiZxBqZDlzUBV89LDJLebCG6sHkyufAlajAT0
tq7WMV5fkba02OQ+6wJNqeiJpDns46XTDv8Zh5UAxHIgfaHGjrwNDTgBGTQqi+Y9
TAQ58t2GrmR0xjdO+p+OtVB/j/Jul1ynyPOUxyHZBLz9MG/ddxmf6IKIJ6rcYCdD
DlIfuaqvQLOg0mleN9lZAh7Y3uvXNkx0Yz4+hcv1c4xw6bn2j1UBSZZsSjELXPLr
UZ8uC9q2+SgI/CrzzjKD4ARfvMMnvhjwwgP35kYOznPCqUfR12fWkt31INOPoF4I
cMExQAb4+KruQYX8P14xgRAQpVk9KM1KZgTMosLrAFCGDbvnVBYIiyJSU0xGeUj2
C2uE/26xQw0owLNFL3Y6x2A4Gp3UOKPYCuQ64JoDnzwfzzTAjnRVfweVN9dZuLlf
tToQuRgzB3fCnOWF9MUikz0/9/p7U1XClp5xRFbJnlPrfTXWOdP3K10dq1wyjI4c
3wq+V23uT0Q79kcgb695IBIN3CGyggIDsGLSA6NujxFT/xr0rm1DrfUp/Xaj3BIe
MOKli9PSq3V2D/JLBrk9XBl8XUlJLwpPSen9BcSS395126AXrnRghQrGZiXUkml4
iscB4gYn0XV9gomlOKiQy8ujLyLg084eM+QDk2c16c5DnWuFyQMcZptt4YK7mwor
qJ305pxzYFiS9TiJza3i6EHp/xq5GTtA3QB5Vb5h7egOWiB7mG5KudZVTKOaljFw
bh+tz6K7sbx4SzHbuhiY8FoWlUIW2S6UqlmSvyySWP89YhL2WbHoCPbIJRFyY4ZY
Zubpo717T5R2+7+LnEBS/RnCGUoYZIoi2wuif7cEkDZEA1oLMDJcyfsYK7dLwZbH
9w55hG2yOVdlbqVO76HI9bZi6ulF1K5WGcIlr4PvYe0lAmUNQN/1V8Mqs1wX8Yqy
zYFJ8LBY6dMzV5OZZxdewbn7+cY2nkaKgcjmFAhXYA3XJQrmU92yfdS2mtO7qNtU
2TXaRV3gCDv/vQfpcA+XUOJljBJLZfxlAU6hHiJgR7uRpJb+bzm5bAmEIHc5GRdN
YBwNceUxVNMeXQ4NuLNEwurTYcoFWhj9BMdsRpQapgqBllRceJzpd+BGSIf7yBGO
sDQ7Lp2i0dstR2fBwEyZ2vOcdOcHOxHSOAlerAtRJeKmvc9934HCPFHgSG/oVTU9
2fdrK8wmrGQN/blUBgK9VpPAg/VLb5UzefVEku7KVSj95k3IYrZm3GEiwUkXtqrd
9rrzB61AV2xjCwLXqbPLA5cnqlX0dK3p6zcKNBQOHSJKF9zlPT7YTA1dJzNQ9Jfc
z/F2mQiZ0Y3qwnXGOmsCn84PYKvcy922n9kzSy9mhjQFNtCGfmWYzWQwrmkLa9mS
+3rMMOvD7aL3QbKYOYX6iNRE+D/N5Xsz3irtf9rhOYEqWB/Zf0XrzgOMURWNrnYM
73zf/pT1elBRr5V3xkbzaWOqEhg0Mt7bUpxJlBntlCJP/Du03QFpy4lzeyIaoPNP
q315X7Ja9p6Y8m279LrDW7LhHdhKgCtCKvmPxdQzSGfBcY9A3dh63rYDCYMaNf1C
tnBRPxQh5sF9pf5ACMbvOWP1eV0uTlDFQ3Xscy/1mnrGyyHHHo8GJCc6X/Plb5jB
zSkC6wwwV2Iuazi0YJXeXO7S9aFeOaP+ZW7NTIprASfJqwbVODp7b0y7uC0O3rej
C/2zDQRZBmrXzYZVLn5R+pDRBKYpobZiDXuBd+TzzU3YjaupuygNOW/pEaV38gV3
cSQebT06bOvAF+Ghau4TTSDWlKiEbi3xYEvjwrIGxVecu8ooufIlty+0Oy71ngKF
0M0Gj53iGav3xnVroz0bqOX7WjK32E3bZ67lB5qlCI+he9SbGZu9y1fQ0tGpZsHn
ct/3UINcohpP4s4a4Qt9syGZ57GgEvd11lUVZ6+VxDzcO4nhEKp2G60SN2Zg+Yl0
rNmSZ+Unn3Fjhw1SdtEB/pC0OJ21JPEkUUPRpYt+rShmNczsAMrAQlrSfa0RSKEY
fm15KOqP1FlmXWyB/d5CV0shshJa8/nqr0O4QTCyW0o4fNPqRsG5aKWDs4zFBBPp
uyKRhSz+Y01fPBo1b0X8K/YgCegopn+iXdFcg2X5E+Cj1iwRGaBPoBaD4NoQurCP
Es3+NjiEYQXa5O9yt7bFQk9TgxefdvbAJgR9n3ya/z+GBdE9SzF4InZ94NSg+bvl
gxPt2cDXNUIxeibEy1Af8cFSc87Ym70pgDhi6MCppW9O0BnBHUl8mIUgm1zqcL/9
EBbZTOD0LfQB5wTEUyswGp8E4rUIiu+Lmf4t0CzlXR4YAOgr8QnWCs5pc2t2v8DO
VtCsofRI/lji0F0XWEAIEoouZ8C1Woz8TIShRnugvtyrc8SSqUOE8xr/4c+0cA2P
cFvCkk367appBjhcBDGG8mhehpZigX1hBq8yFDmE7XQkKQMl1O+GGoVpba5h72by
8saFa0LcIBfch/wqh3PxRo4BOiXipsfze0GB9EQzD6+E7686Qi7Gf08h3AgqvlT/
s5F04kYKe+bL8gzemkK79GTJx0PFlsSvhQRKI3/sBwxaj55sGRo4j4+5nnRHm9Ke
7iZFw1l+0ZJdqgwEuBSDAhjYkbpEy7O5qwGEnWXEjSmrdFUx+tjNPkAMT4145oAG
OuvZVzOLRL8CkV1dKT1WIZGuD7kfcGjVMTfaEO6kCR81i6E65ChfHT+gidvIKv6U
+GuPLHIt1vgjItFynE6f7RO7gGve0i9k1RCUYbfl0QqbICRQYibPl451VhAvHAub
7ik6gFI2ekrflkB7RE+TXg1ofWVUiuTZ5ZtjFm9U+YU1Pb+2zPxX3pZEzYgiUD3J
8vdWBEE+zrDceHBeTTiOATiMn8pezzvB7b4vF68kkHeuANt/BJPDZfR67OWa+XCK
5csLP595CMO3FYIEixYFhDlxPYNDQcriY/PJdBkzYLisE3CFMyXtiQTkyT4cBYcl
X0b2YPBDQFiqG3zd5L9tMprVqnmWnN5l5G+b5LdYDhr5uOVFs1RMwe86M3WsnfCq
IKP7FjPMqfahgPz0sE1nf/GS6wlvUbgFy8MznnaVRKTvCfXANlmI3XnFG9TCnoIB
HR2UKOaqIDzVRDXxmMRPmK+lMrXuAQiN2jRJ5oxj9kXYZjvaVsssO6zTbIrmE3Cj
ozK6ESWsDWz5xcV0gUyrgIlBJUciGXdohEcgylilcaF6xJ8J61cKZlq5FKEoxoRg
DqsG4WXeDvU++v8JdNCJCN+YYFoHy8tE7klANYl9ewjOtUR6+4xrEduL5St9MQGz
r8VZiyQbef1f0i5DaRcZx8td53CH9brW7tqDGgAdt10ZoS5Iyt6cFT7Lbe9KdCCU
DFls7MmLj9jUExwmX++Bhk0z0i1aLB64wBJkWdcxl6xh4tgiKG0m0CAqjWi1JO6d
FenqJ0u1IQRp0WZW0VRuOPSa5+BKzYLH31bVF7g3TcdYc2reVnHTr3cs6YkYEtB9
JN87ZgfK+CVQJEXs80OU0quRUV1gk+5UCDd3Ng+lFKq9/l7+Z+kzrKcRdc9MXaff
PrsZY95XQt5NkCslRJwhGBoQeepDrHvDrgXT2FDcwJTMor74N0qnaeQQrRfcmcX1
rHeZ5H0Q42s59GEaJwDYcdBPGQgxYBlQjiEH203AfFKseRQvB1bH3VFxr7GdCVeR
NK1r/JOzfE3TfrS9PnvNonYidq3pUVqQxAkq/QyUzG/mKYRQSgaYZJww7oOfLJIF
4tLl9v3E30X/y8JwFIXe/JXpMNAILPUcov79o04t96E38NGBRQVuHdbDN4FDQaCW
AfmPCZ4frVZaveBLWLilFecO/oj0ZFuX9IMqhBPj2pBXiU0aJPaWu9kaXc538Wl6
mahv/If0/7E8plceahJsI+28hoA7lpc9PHmxp3zGFPF/wE5xuZYmzsbzP9FQvXhj
Ap5tVyAlD67dHyrOn02jS5DAR9U1KtBIO5TwoWAQWBcWN1JF8Ku4h2TQ1OL+QUVj
tSI0uAfQQXcMXT45HH6JPZHgasgQv5sfuXLuu2LGEKBS8b7Ve47Si2WsAbQ2FYtv
ngK/W4+ADHt6K+EtSwxbW4+Rz/eOccHOJdFmr+StNvBhIN08XIZKZcMpgW+U79Bv
4nNMMAYLdm9a/68kL2Z2YYMuLhKWyfYlbj+5t9jBFgGPRc8Tilsr974c95LelKh+
R64WlR6dlEvfL1UEH94WIV/JGYVna8YDK4Hc2PgFy3C10h/HhejK+LWKMuFV3X2J
X3Gtwd4pSfVBzomTuDkoUMGtAWjNRpo+z/g8cycphc/z5wJ/Kt6jaTpCw2LTm5h9
fmNrAQZ+nQRIu0kuaIKmCKnhzn1aPq77qDj6LbDHg5Q/YmeBX92gxfl5TlA6NWFT
5+DL4JfIxGPYzB1cltzr4VyJHe2TxRHcDVSLFUlQamBF63+jWrB5/PBjtF7OA3L8
F6sLmjxmUuMsLU1gZ7JE7sMqkDUSOzHirNDEGdWxgdd8N4quarOjHp2pxcTBG7t1
SQrdm+f1GFGmy3g8ogqRjPgWn3f8p+jTMcYGgUN3phjJ+2ggUWAJKlbQbIBW9pN5
yCNnezE/8hnqjxf1X66TDVXI2gF2KzXWvUotloQL567S67EDMSzivWfftlmbJ5WW
5C7orgYshYcoGXT9rq+OIFScjDhPOFBgaiLJZ8+g/Bz9+GhzNRIjV5wBKL1hFRbi
hZ7mORSy+n+lwEwjCZXrfOxUyaz2TTrq+38yRRB98nFjnszTwWXii2QetH+jqvZ/
vQHgjH1RIG4u8HcT3upjPxeX3RQb3HXb2dOcwOka2RvNB6p0OEUdPuWX9amwsUKu
CJU07gWCj88WCNDUPnO39Tg7aYcX/trpFUFIl2ZgAvLkXI+ddu5gZDLqrgplTdWk
ESdx/rOjIH6/u2dl6Wc2IFLbnzhS4ii4EC8lewV9tuYWFoX17Tu6rl44799FD2Hw
Ueh88yO0Y6nlN41NCVjC+Iy5JCnBgvbSrYW7TSoS6gVIPlVb2Eyfyo0b+AfDWFJs
MSjI6HWRKwlSQ7AX6t34bMl6tKgDHaTxCwuaIvH/6cUdDyzhiM75HvBtzRbObxMA
CGK2RlR3VMOs0Mkz4JvN6Zly2KFlETYfKciyOM/1/qm5mZZBOfoH47LosGavKI87
rlNYnQ7m/WAjAUFmO9/jzG6h1XQ2TVCA17pJZIgmmhEax6iL+2O6juwW2zf5Srp1
rD+D47NDyyH4xopB+l4NCrvW5/9PBfQJFAHLFdNJkthlYxw5AjLDmHMUsrUnXs7Z
i8uDrLxZuQCnSCuoLVrO8ZJ5CszKK1FCZI7gDFWiMYQOa3dNGGJHfN+SFJ5H8uW0
Mzd8G54AZdH4SDgmcsmKrFYdan7ZIRCZ9zcTOuRzu9XF/YedjVfGFzsQ8bKoLX2e
B1Q++jGJIAfbkbQmE10quR874QMOxjrrEMofXfD1VwR04H+qCCDMu3jNAlTOsnvW
JOJkRanuaqsmOGUgeYKTUu1QlKu7cz6nSZN59/EYc+UrZUL20/udybrJ9ykhDLcp
yAyny/j9uhFDxHC4G0jb8OakqgzsDjkq+bVoRIkHNOhhHNGKFKsQpCrG2qTjMt9T
qloyhj2v5BH55or7O9WT+hhTrkz1+BOr92JzxmTLsuG1sUxmMETwi/4uMgpSPAD2
lDPqdlOUewLPOHwTCCza3qLtzhL0FPSICKucC1SHW2ZVqqnBMsGQg18NTYMJoH+D
TR8ty4qk7rqzzQ89fOn0LiJR8+zsKzj9Mz5hQFhlShguL43ru25E8zigrKSvii66
V03ypdtuPofK4FDHwZsM6492HolOqh7z57R9FmrWlbiJYE92Vz1IrzNJByebYDwG
+W53kAbWKzk4UvTXbUu1AwPImBNrtmE0oxISCNT+L0l5/o31mlLVZZS4KnxBYWwv
kTGgsRz+ydGsEAffUbEWNtxlNS2r3EntVsuhDf5G0GOAcj/em94vUEa4BULJ1PyU
Mx2YDilmLfu4HQpLmPWLG02tgTPuZ4Lz1hLRWJXKsde1i8l1QCpvVaTz6OXHXHB2
p3Xhj5opXQvdv8icttFWmeBQpTyDxmP2YglMEOuWdVnHQQONumXN6Znq+eX7mFVI
NP2NR8M8lvvE487nIcPvEsLVoxh7GenzCm+Le3/whdOLeNzm79Xada5E71Vf+c76
XkuvxKAcn+rtDXrKqnQsXJ6c2yo9UAuF9keIkNyGQ0OijvwGis6a3a2zls/Wuo98
oAi7SmqSGdjtY9EGavHj+kqs2syA3kAnGb8Tu1fKhRrXfqu68GHgg7f2A9y4XseL
2qOhZv/qPL4A3ZymPTQvCeP639XeD2R4GueDLnZHiPhMYCiBTgGN9S9gI+DcsJhx
yWLABVHqTO/Z4tXECCFQnkpmpMe3aXX+ZDhMWoVH2cjHC5VZEVkQPNikhgd6x9/9
/PYVTUNE1wPe7OATLOqmyovHc3cfISh3SMBkc9tbveVIJv95f2AvD8CSmjmek+0/
A/26rDhB2Plrb85zLuyVsvT5fF7p8QRAjgnXs4PvItfnkxd3/uYjzshkw95cwNRN
v+OkBQI9C0empehWBXcK46ugdVcov3JmRFGqLGAIo6sFIIhZWq88VcVwDe+VErmV
bt7dbbJYn8tGEyWf/1wIrcISWyXURjhQGCtLinqSzRccwA6BvAkmptpgQFvmSPGr
rvUTYSDyqzwqyX6mtNY76MaZoGlI8puqIiEtZoSowBna6cBqyzPgyk/u0HHqroF/
G/s7OTFQ6xoS1nUgUNDwP7jLs3iQl0WSBlo/YTa9/II7Tozw+2NyC8uy9MAUVKtW
D78xjM1ic+cEgJfP1rB/UJT1m+REh9P1dIVENV6Oa//uWrVKQL/zGO1OiYGS8IqN
1jKsUio6/hNM6kgnjKxKv5ptotluZD0Xnvgz7c6FvYzcsQnrmQnaS8mpejnNvw6T
XT8ZCDh9Jrr4j97At8US3vJR38n2UoraMFmIoLq2ndFaLndytwR40I0LJkJJ0ON6
+Cy52dtuG87hLHwhZT4II5CowKcQtodYLZh03V9UO3YdO4XlnY/+2MeVM90lC5rB
g7p6jT9pFlgTioC4sxIA1EcfzJ0Fll4bfNyCvdLiq4McCxqPNp3oeerBXQyBI158
QkxDvSdRfihfXw/7Qd+c9Tdr09tqrNMGL/dWRPPYEkUxeiUKh+v7nWjtHVP8x0xT
BZeiOUl0EtobPAOOJqinKjbxslH+N71pFIZuGlSG/RdBqEP/lF/SAr+sWYo7AFWu
qu552OFgbwfxWIQeXFey3lRT5DtbCMKfTZeNw3rOac02cfUhyLGURSAjuAO8oLmD
ifKrT06jZBlGKQESLor5C1pk5a+bjTM+OgIPZGraLTkQdnLCYpwX8cPE35LClqKY
Olj5e6O8SzMbI1bo6sI82h7qfuH6yxVQY35UwVM8cL1a7qlVavubNR0R0lSkJ4/s
LPoRxq+OK5N/PsXVBs/So7NPHGRgAc6Vp73N4n8y2x4alm17JjUfm30/mQDHFBYm
mQdK/4ThTm1i/3rfWTWpa9f876z+v5fFq+6w0sZ6Eky4V1xZsRUVb402hubbxF2P
PerHS1+/vgqJHxTNV4ujI4NPbyiJIApZyhIdGj8rqocE4Fb3wSAbK8d5lhM4G2Ok
2fU3uVrYCFYpBt6NBKNqU0t2BNq9JA8K4EavuQIITmSbOBxTkAyCFBEW7eaJwmiV
Mk4ax09bHCHs1vjkyGni4ezKQG5DTMH6Ojd/6yw1hgpZFRyluEu2ZSIjIM0siY/+
k8/6InBLWkQNGrumvapnFfOq6AKbqo8/1HpEhDcYuaFabVqS3NH+JM5GkkMwDNVQ
5v9PXyj1k6cU+Drinl4UG0WrWoDMds8M+bfL3nVCTUDe8fYw0UIekXl/ZAbkpaA/
d9cl4aguABlJSR1rYvmcNFW7RiS9lfFF57EKCuOS96uy5ASCl+nPZdaL3IhNCY0H
DqYI9at6FB/MaV8p3p6n9o8k7DYddHDlIzYnnxUfZg424mR70QL/5+12XtwAYa3u
NNvUkuNnUgD37zIZKTkhwsmwnzaaGXDnjk1Bj90l+LnziIjh0RCGYS2fWwF8BxUj
UHwq7BtD2ZBl7Ea7hmhGwLkqZzKctXLLreNhKSUgcJmM1hyl4Fw4iiW43FCu+Y14
rdzRSIl56Gzla0QghsImjkDcwdhRnEIYjfW+fhqoKGMLeUrSN2rPfQrMgLyog3wP
Z1PBrC+6tR3EuyjC451q7ji/DyK8mk8wszXIDbrom2iVxThYNG1m1AcjR2jP23m8
nhH2IsHzdNIRzdNEDi2C2iJZuXQMy6/SSb/J42B5VRn78BtJAtDGCgpRLtTKPkcO
VJpEBQhkqqvTix7QOGStH6IAk25U9+xowRBe3aPrJy5FOTjXh/GZ1U21Bwm4LBFL
pJ2UsEJFT3bJh5XrZXizVRJRoWAwxPvkbkga8+ubTwvF4d8zBu0K4SbuH3gxn7WP
W/GBhUBqV29KpNJxEJ00Z0bfywzfK84a2EkCDFmZJsBkNxGSAxitG5cdOeTWrCdf
wUPMUTdh+7CNKXFy4QttZQZsIadzdfFUnDDODKzzSzjsT8eFOBKIDt+jNGYXs58o
iGONJz7JGQgG7PNNH8vGrwEMc1g+oCB+SbK/WlEdUZdltZVa4OUtPvxw3NoFIWTv
lcMapHXnGg0OoX8D1spa4KEFqwgegbQfejvU18d5mIGVXU5rHdj4VfYAFlSzpD4h
E36R3oATy+UhOkht2sVUGEecPFp82oyyMeYmTymSptiRNPFXnDwKRVzxB264gI/J
lM4bCFoJJB0eIE4wH57oMg9ISJmW2m8yoYtjeeSKJvc9yjrGKDHHlvuLIzy+EgHo
XU0Xu3TbBFLUaFfhF9EP2TensHEYIGYFJ5o9T56Rw0fVuFiyNA+HvsfPSu7M+nrU
WOyTY9MRo/fMH8yV+ky8nGZVVErVU3l2SPO6jWYNUxYeZCO5tYpqGnhsMADlHumX
1baiKau3D9KCDNEnPLY6AXIiulc6iw3+N44Ui8aijMIuXYHp0CrKfF+QzxHxG3CP
gAfpSXLnePJOMt10aDSDAcu3oX6vfve7wT/GdJ3V75FPYCtqJBA89/hEKW1m1j5O
nb+T07QQGyCeBZ0ptq2NBqIlMVhBA0K50X2Zxb8FhQTRVkYo+DyHTosm6NovHX3G
OWvWn6sR4/hXSadYjwiPlSvaks2GRplcjYsjrXlh+5cuNXFBAucxzPjqrg0u+SNR
1oDRaZ3BLO4ciKN0LS5SM4qEalZRxyJpTgV/JfUE/R6vqP4x/orojOkyh+Joy6ZD
R8Wp3dT0nAfDgojBxun22C2sD5DTBWPxEL8JQtpKvGmUdtkRYMkTVGXyFBYW1GqE
qw2bFYWxZXTyidis9PkcdmjJyneOXo1qtPVQuu8tqV1d+3lA2Yjk6tLGMhN7CmNR
4MU86Q6L14oQhfHTU3FWTUAaXJbsoWQtJnBGlvDQ+kSPF8+bv1b2VMQ2nXAWTm65
oiAlxCQk1ZIwQwJBz9tuFA7JHvcaNTUq5HAvjGp8q5dlVsFkqiv11HCra00gUIne
u0xTMa3nw2HUUUT1e0D4NFo99cde35V5MbC5pub3tv8Smh650KBJpIT9JSh3lzNx
jSFesyWGgekRDXolKyeO10dXx1Pt1Jgf4hMDtjRTJ9/nJet/jqS7azLI1y4zWTb7
KzZowDMTTHo5WGq80pIcruvyF77AD+SlfxkIz7xVK17uKJh9TYxOanWsGhP/b7Qw
OlEczJwiKyKujIvSYPI973J2WMROwyprmZJio3nWvNWVIODfklBb0ncfF+cCtExd
4Vh/KrEQS5ssaJem7aUIhsfTmbyQPHj3TkJQFg/MuCfQKSO74tChNnyJZiSbkDr0
cjMYIdW2xeQdOQp1UhuTZub3CK1oqMf2p8CtgNWQoBWIRvBOCUtG8MNVa7djICMf
Jxd3XoVtIJawIU8rxKi7qsvAToA6SwwUDnjaon+0aqPTAmCCA03Ihoa3zI6r3sRG
EmRUaK/DbUVJ9DW4GKKs9tjQm44VS1bnkBy2Ol4oKYEkfQQBKGSDgfrsfB5Iqfl5
Min48WIRFBwhFYlA0e3BQ/0bAuHhK/GVPK/Gt5qzdMGci5+cleNqu0advsBV0alK
PGrIE5pw9pA/2pQzVgoA3/OHEoA92P/cDzXNgV/7B7iJPrP9sFv8YmPK4SRDsrm8
vgjquhKCJLvGCPuzjNyJ0HErSLRy3EF11s0jyg6LllYXdEC4NKZwiOvmfr9ou0B1
wv+bO9BZZniTSq0w37TLAEA+H5EoPKlFxpsxcVypmafag6+Xmv33tAcKczmHkwf9
I9RMkQZFxeutZyQ7DiWip1TG0IaV0MfzqnsJhOmClEs3H923nyEBTaJ6mFFJBIst
HBQ11/h8MXcgOyfUPdO0uQkzjqiG+UZTWFkOM9O3WPkfXMSOT1cWXJsrmVWihtP8
GzmMCKu3btj5aHd16TDDDUzfngkgXFoEpB2KL6WNS386fftrGtSiiaO0oRIzncpn
4LMASOppSVmdQR06SjI1Ibiq6+mYJeVUxjTNfgUzCJvrrFhMRiHS0jb1jbGgKNgZ
GtQVkwJKIR4+THJXPVOAm1klyXWkdsV4P+RSWJIpJA5PoJwxT7mhAkAIPNog/tVC
N8fy0Id6pWjBh6P0dUX2lkEhxGGth2Zy6MNpXVHkJXqjm4gexXrDB04z5b37lgQg
OqXvVqbqN9nwFAIgTUKBPVfJqJjabzJ5HRUmFGxosKuxWSQEFiSIMgtDK/r1nYNk
lCScK+lBLkm2WPp0n8hvGzTGkbRVMarn/Dt5Tzz2GIGwkuCXBWea6PGJ26Idm5A7
oHuetCc2Y+lqstmAmBURxLPebt9fqpUPoqbBByR3g0yFW41E+PtKXIRnTIjJ+gS5
kc8/TNvIJl3+PS+8qYt610+ykZM79U1pmp7TGTTbw3OkB87ouLAyaO7CJMt+K428
Oovig118guean752BB4b3PZ4uNgRMrviN32cIbUG4kDwDv0NU23N+hFc1a+7Aj+h
HcTvntUmFUpezOBGKM36zuu2Hglw6L+2t2xSUoTH77N4gSMjP8FMNOnu/4AgaiDi
rtJf33HZmqvZRQOJyhancTleAK+lU5e8vK3NIYD6hafjVLrDwJ/Sx/idIUtFkizE
irFtsIuegBDTsRHM04LwphSEM85f0CzJBnufKoNI6P2CfE6EX1PCbN6fukEMZ7d4
ThtoVmcGaHJ1+Ccsvrz6Dk2YezMczvTyIVp0l3h1hG5Y2LlHkCV4YcQ0HWbB6AlC
5UkX1w7l7ylAUjbT9ugjVy9Uct7FGHpOvxqok51jsS5us8r4gxDMp38STvGa3Qus
NajTjajDpPz+Xs9YEVt6py91txpaDCOrgN76ZieyK/S/bVU+Z3c+y/lPhLfUIryK
wMpDWkwhZnDnsx1L/igfNXOoifffRZnC7hE5qshqtCcq4z2MAOumuHyM/EwexBaT
xh9u0gwwrCJmCkzLZY+ncSnBzL1iWQhrprtb+fUAUnZiLfU6GVpXOaYMiTuhFSQD
emMl+2BS5V0qfNuSPfvXqIcl8FRbyFy5WL7nV4QoJ8VRqF0RNjQQM0JO7rQlPyh0
hamdn6D2IJQxA8V5ROKAVV3qufKVnM5I3xcoT6thX+nR0kHtTmIbMvL0wNApbxzi
1G86CLDu0rFEMjHB/hn9E865EttOWRTQPRJ4HTqJ+JmkoMJaoo0a3EBaj0hguY5T
U/1S0nYQk36vn0hIo/EabxrZUKgDBl9aRWt+eCvLlQnMKKTxRrBgDGYQKim3SQcm
HQOD1hsJ/KXYwDSibsPS4LqCucP6vCwP/X5RgccWVLCGGaFVSzq3lkEk6IC/nEqU
FuvGbXfxVy+aZTuCOLB95qjQUVti1lb9kcLnNWB357I8L3V/yTPVf/waW6+C+zTI
oz0+sib8Hu90kbKjgj6sRWytI6iLN6VYd2SBMVVjeqiuBgi3NDkjotKL3PHxqAOs
9XtHdeinc6FrRwDa9ZmVv4JZCEigtnMwwrsAjB2xvL7wicfeFIFWvt0cq3RGSUnZ
EjckiT1B93Mk/eU9rp9Jlcq+Gpnc1KLsWQx5Nr3+W5SVymw8w/t1KKDfX21zAeCF
WfUiOmffxpmZYFpmDwxezOQHSyO151V4LABAFuS4nsCoOm14fSoElGJuM1aPSJFM
QU3eefsZKBFJcfy5vkMdSBhtVeFDr5Pl287edxKwpZaV+u2ogzBdk758igcJ2ZKc
tRANGsL90AuGmmkcli0Kk7DY/AY+AUNlr/uIDaixZoHBKa7E4nkVS+IBflawLmi+
UZMfyW2JuOfJ3TS6QyePKWrJdDX2FJZWAXGc7Z+PZGLS1WWkzL6SvB2zjH0w2Tsy
Hp0SbTicoqFAkm/whrUQIudpreFmCcVZk/ZsVdaIXqIke453YHNh8k0I0QmLOxkk
KIeC52+mJyjqw1faVq2Uxgp115xDPlJUlqpmZzbf7iJnOjd7rN3HmqDtqjSIs7OH
Hc59R4nCDdCvcSKdMkQv/iqZAtQrPZIXrYFARzH0YzJqgV5Hst0x8WJ2dsauWpNV
//LXpbKt0hUXEa6CiNNqxdqRUyXhJz3WnJPj7GULeOk5Ypu8QvJiaE2BcbtXTgiB
26C3bxm5ApUsJjE8XwN6SmZDUPauzob9tLsETjbseUIaIaWwSnaVfqcTYPbeNoid
vO4oHZulw8L1/WDDqn2Od6taxLEf6Y008yHS2s1SuHwka8suiYRzuey/umbah4oX
UfF3rpUy+qNftzk3wlk6RjAVCWvvJRWTgsWX9wIzG8yNT68Wc3I5X3xY62/JyPFC
AU1ZpOSZhndnx7hw/CvIfZ8qIpNqxFALb5uECwwSoe3WV+8eGUIr3jbuR799SwdD
BbC889df09DnIs3biMuwnGaOuo4JIBBmUxgUy83KcXJbCo6L5uIQFO8vC/jrbEzF
Yw1Gh1Kq8O3W3fj4lFWpRfZbG8oVEH6ywI/OKuCmL/3ZsXcjRjF+QC3AgDcpYof9
mZC3rO54pqpy/TOXhNd0IiWxydAMePtvdSAKGJfivpILQo31FKq4HkZoXXZgOw4D
2Z57W5H/6/sBHYHuqcxt+nDpnTbjZIgC8tRFNG97iDsGfqQd1br90GMTWcD3qcU/
u3OukLH+Un7KSa6U6F2JE0n+T2E0akaFwqtJPwl7oOFYmFrO8w63b6XuMda8riY4
jtx95va/ZMl/u6s4dCUIspJ1EY6c9EWpDRO+mYS65qNqHT7MhyZzVVyoahQJ7RF3
ymo8MwuQfAxvVPPTYLHrRSpnPvQRCc3Aw8viem5HiS3A9nK2wUh9YOVrIzzmRxi6
+4UlmDCQixLE9H/XvLbRyiWEY9iYdV0fwG/I8aL+GU5rPnlMnpWSnqyOEPLFbMH2
d5PDvLZUPXOyjuSzQm2WfgtWKaW4QyXHGOnz03cfT3TQ3WrAj/ibRIaIge1zyJuC
b4gv2XrjshVchpns+TL/66A/djuQYMu4uTmCUE9bhONbKv39Ff3ycIWWC9QhVMgQ
jxCz82OCn58rlLzOJASYdqamqHSf7JKVp5N2a6WqDR4IuV6NdutHasL37kxWXOvY
m0zm1QvF1Udf/1m/DF3tnAcnhSZPqQMFVnfgnTi2H6SJ3jO/gZ2fYhiSK+2WV6xn
HtEVQNVafUFOx/HraoPfJ52paz43r/r2vx7Rjb+yfDuUvoatwU4F595EdpEGeoSS
vALmAo7a80mUaRvTJHOfNCiARY6T3ansQxGoJCo/oObTr0ypaiNKJftsVQ93RUii
wdgHKnPKOssORK2+fhEG2CpposqF33XjuRtYK/ez2IvhNDHMQBJN0QzJn06q3twC
jCVqiRcJxA2fANpEGijrAQEqH/3fZy14SUiVgmVnR63hvEe08zAVT4oGZq0nIbZr
ZaEL97EYqrmlREwR+I9HLSosBD04NT02k2dcRholY8O12+jfSxW2KzSXF0ql8HEj
Kl0rQG7636/7Ii+O8nMfzN58O7lTBAEnh946tku6GlVX+JVxg+HMy0Ru7eo2uRd2
7I7QrcwDj7cXHp+N15FwNS9Cmy+blrQg4yjdePmHl6Z2DlRrmg8h8psLjbjqVhDH
nR8B2zc9l851Vzt5hx/28L5AELg17gE2YmR6FaMY2hzxzR9lbvceoKm8/nAAKJ5i
oDFcpQjPAq+kzJswyOR3qbq1Oi4qtllXs0IGMUcU1H8Snruie+QUR3iILbpN57c7
yCtIE8Y47qgANTB/oQvM7hD8wOQQAVeUASaOhTJ8rADxrgnV76JDuAwmfbGVvH/i
KDRjP2HJgUzY9R8lJWcZzvEBLo/a0aGkkdQAfHUozbh/YqWrqyKLstP/q2GdKZD0
mdHJdD9SmcRJBCUPc6X/gl8VAG7+pWM9BeQa/b0vz3I8S703QAqW2ZINVIyAmYrq
xgKSidxP28mxrW6E6u3D/YP65THi4RiurEUCQGajMiSKhgfbJABM7AcXdX5mDJg1
4fuONPnSJyNsqXFUt0DXdxjGOqwdGP6VeFEq3qinZJZgnNrKp/sIR3PO2UKw7dTU
UgpPjATYjejx7GWbVZCLWBNTJHo0hPt2hikEA3wEHV9ZyvEEmmB05kswR2mD+f96
5wifUV1xsLjQon4jqncmhwLoCVZfwyqVvSbhvcHvAn7aQMReD7XQ887eRn1UXnRJ
d3ezZnJ/85Y4KmX1YeDw7her7rhiZQ4kjgVE7tmtgXGdmqILjH1+OBe4nI2vSL2Q
SPrJPh6qPOyl7DpIr/CyD78o/A7+Pst2AWZO0fozeUNFloV1abtbgdmj6LPdW5kZ
IR4X1flnY1n0SMOIL2xz4qO81E0L7FbIyp+seeCgg90QZNwL52WjrGK3PNcpUTyh
Ot2+5jUyMmp1hFn6adAHuWSMcyHPCD0NzARNMAeK93oShFdK/Rno8vT0+HjU+Vfd
4JilwoGoegWHqpNFwEO4J9lW0t2pAbeBCI93d4hDbkWoofkWAMrPdThmwzxvzDXA
Fb5DhmlsN07XSJyMGvt5UpLhKHywEjrNbXiWj/fX0XHMkwNNgbWK5h8MgYy9T5eI
qLBvwvBgV+12/sRm24qNcsZUWm6UnN10u3Z23wmnQz4pnM0fxUcTydQCjeDseCaO
GBVccqIQ4VmxiT6kiR0bpmK+ESLki7IV7Ma5nFcAPsHnicUeH7tqSCJ9NU9YVfjV
8oWg1ljCNf7YY0gcdQDAIjbSOqBgOEk4hhPo1Iw6gt2U8oY8e9go1d9qPGuWuRWV
F2TU0byim4/wlRkZFxlM2X/2hfqUCd1dbPFc6LTJe1HzDizPXiCMtwNSqwWfNJyx
cS/jDfr5/08X4DnTRbtHMPx86yYCN9m8IFkUOr9/WebB1z/usmknDCKNsH2iLeMI
QNSmtw4UpQa9vJpSd31Ygfs1IPnu0yzRa/EFy4TOqctB1KSkiEp8SdnxYnIiyUmm
9m64IfQ0Oqc4XGyMQotk2OeHE0chV/xsb9y3kcePoyedxI3MNe7YEgfmCW2Qz31V
UhNAgB/PaEC3WwjUk7GOPZuZcmbIb+65fkyi0iGovfeAxNhjvn6Y7CYD/VZPDq6U
j1QcUes1Cxv9CFTRd8dY4Yhi7Ivl6GdA+JchQgEu5EESWxEBGXVHI1Os+sfPt5oY
ylHb2ICN71g5Z6tJSJHacTUD+G8rxlLWcuy0VnSvWOsGB9SSmXpm1XbsDieRAJwc
TYRu5FzOrvkfk/P6H3qbPAcNWIKJphJNlM+rv3UbVj5JklTSJF1bSxbd9w3CoI3g
7IO2u05rRIqGcosF7n94S5FiunL8xORtRaMfOStSodKUTyZTG3H49A3ebDFZSt17
0vmxpbUEcySfBLy4tWyXZZIXbXEvUiOTqpVmd1MIMe5coQCEfPsAqhmf8PFcWdXw
XXuFLFe/QJqgJCbjjSqQC8hfbCIzjWqaNfWKWk/s1aNd2RNKIzTvOr1nlBUXwvOt
g01Uwb+enw5TUXtmgYxLqVOrXdNNvEFF51A+B9slzlqidEdSVsH2WPr3HY9+zwll
EGB/KReeIBqUPR7tQAhty31u8gcb8woKS08Voc2ygLcFwyGDWT6AVzihcftwxunq
H9jaW5MZa4OeVrt1FsX9MFq9IGOntmcAQddhH9G7A8xDVa6U1Mgyp9GLJp/0X/lZ
5edObVIj1RO9GVQRbhij6R/guqOKzy3Gw+m69grhx6oerZ0TJNg6zzRUzz/VCp2r
NnqUvQOX9pxBhyy7Gz/6+x9V7sWPKSMN63JI40CV2TmiR2D0+sa9iINAk1SZ4Qvo
sx/59TgoTYLdslDYjgG3q3bsVGdBehckh9XXiqGHzquUaOozZEj1fU83Clebz/FP
i537jCYDHse/swxanFG2AtA21d6zPGrp8R2eyPQO8NajicqE+UCmUFU2R4Klb86k
62WXCZo2y2NvyWcQX1uY/fmEGHTlexBvTJjkGEV8CIxDUFQSPNIOZ4fcvbqHO9F6
OTlsJhuFvqyuZOKuhHaP/QzFEMaXBogjEFk40i+Tb53S/AkUvzLOcfO06fS2jbtY
JhfZMdvNJD3PnomqZtUQqOHrlp8LEjV3NMXd6tTgGBnIh7oHnXa4DbnzJYgMX0xp
mVv4ntBilCFR7ipzm5YmXjwQNfQDy+VjkVNeQg83567kB6T7yoGj4Aqrj7e1uMPE
qI6SgSC1Fe6N747Q1u6Dx3+Pib1qgfcApKvikjXPMMscK358r1np4Tja6NRFKvCK
V47/NQ3GuBGNKs7UGlc/MimkRwDmmJk8AsVsn9MYwhWDGyeiwJUGSNvsfYdR6+ve
9YVZjNV6QRpoHizHCaqxHANffvdCVbGiVxZZxheakq7r+OZq/DSNhu4e6exTd8jF
EcF0icKKYOJMcv1A+PL84oRTo5v8RvXWa4BJwb+DLQ2Y9mg4juidBT69g3rsPYQG
co1fIXMDRekUNQEpzbLoaR5wYSylO+4L6exrisNQOdDQHgM0qLJJ1ZyBXaPc+/K+
qaN8470Pg3L9GDLEM8lhh6IjHOy2q8yV42PBIucwXVr9mFQPvi/qXhgaCM63cM3j
lbVXfgzgIFJx3kvqoCTnkAZ9ZUlOxEsdFhCmQZs3h8ZIKECyBZsGLIZY9GXRCkoq
HeoMUVuqwf5jknqoIPYQb1vnhryAmUKOqX50E/H/P6s17IAUqGq/eAwywwPwD2bJ
D+gU1GfqurfbMiqIxYxIRhRzGr3g+EIjMgvKoSOTn523234/t5RP6NrCdc2Q4QE7
bU+mK3PAnouo9cA/Z3/jRFnPtbGfoaURmr+1OChDDfr/QBq+PHwemZAgeUhn3GyE
sGr22e/dpoloEutwjLI9ga4ssJyTXL9RgpE34UyJeJLPcBWJxaGp4PzclpmqHFVO
yT1oK7PF04XlVbD2TEJZZslNM3d6Ji9+A7pil1OrtPkTLVxKmNH37yqADe2rsUag
DNlHHsgzQvl+EGvXL7bf8a6RqHoFZLOMd2Vi5bGcf91AUAcsbylhxnMfmFg2iZlJ
wNsc5frael5OQj9ialVqgIRSqWI7mJTXgPrR76I4X+4uE18ClJgLRBxXRk7LoS1y
9hv2pWb11LR4Iseuyi5F90xPLlud1QrSv3YKzR1DDF/4txlrm5YUZFhxN7Obp88n
0f/94Axcg1R1PKo/r8MzR3kgy7tgy48RdzoxftB4KA57QofAbYeyGy8oPYQuTzuY
Nlb4Jo/6zpw6ADF8khEvIx8+DUwZ17oj9XtU7SPXZ1sleO+LsdqAl4A3d8ow3RMv
6uqxA3onvwRos8LCdJqm6/ACMo5KtxJo627sUC/WgJ6aqOlTanRv5zj9DiEBZZpn
MeRVzWd0uG+LBwLgPBHl6xlmTbD5Y38Ceg/NzeDUsctU+sRPayRj1zaHtviS3For
TFEXdgAGXUO22BzS4gDZ59rIQnxZHjzY7JkXR6NDnEZ+/JHrRYwcFbcsVgDH3Oi8
QTdH+91Yk+xvfkPDJL4DfTTm+i/VRRRkHsWAdaHL5R1KIVbrR27neloEvVEjriyw
2mQMxlLe/4zzD8JF+pzQjryKBIg7jXjPIJU1FcbuI26GG6W6zJA66kRZDhS5A7UD
++AQqdfGuLoJ7rmfHb6Ozet4Kus8uKgd0O9lL0jMhx2/0Dr+n5XCHF2N73m3Hv0f
45Z95tWuCe3wL4S+I/r6b0a4f3b5TRBt3EKCKAu+KbNy9GC21Kc2S6Wy7e2QP5vw
AWWfiU/Hk/885kTjonUPEcIQvGwQppbL5mY611tK//uTpCtvZRKeWvAon/1ntre2
cnfEpup43uzjaaKPxoqtNYIoDXVJ3l70O35qlpxc/HmuragEQSdEVm/RBzmv3CtD
d1vehMZbNImZ525VM0Wah0sg+bJ1MrSD3u2ObGmw/59znHgRwf4mciHtvGe5Q2Km
7kbpIcQu9oOw29p0zULjUAod7h3DZq3TJaESqEvrY29MeL2RzGFAk5H20aUJpAhc
0w3ThbcLGMXzgMiIRXa4ZKGEQWHjmlBT4wfPhNcbiCnbgcGcryJ0dnYjx+w9BcM4
z7EmkNljjLnSNGaaDm67LvoqAsKBENMH+uiR56JChYVMMyV7Qr0yvrZolhJO1o1W
GCIPKvB3WLLPc/o9GzZxKUs3HbsyD6flO/spMwyemFCQZZlteCHNLFdT/jchU9UI
oo4mngZSekLsE/hplQydXN4msXOvE7+fVJ/7ICsedmKjOlg5zzpqhOCLvMc8pMA4
OHC+MKCZ0JnBX//lKnfpZLv8xzhk7c4GEhWS7P+Pno80ahU+DghNZt9TUzaG4qD7
diqmjsxiAXZOHZFXLJl0YVjpP8R6vcUUwg+ZCdoTHcpqlHpdbzE2TrdcL5ik7MZE
DUXKbllHeptLGmrndhE0ywuxEMA+qOfnWp6rZ7mnGShuyXgh8PjNZhgrtTaNOXQL
4i+JREHYBU1jaKlTAAnqbt2l3fjRxlmtb0MxR10Cub4CnzGiHvcXsK5CSDefVbIA
b96RHu7FHD567R4CuarX+NPTCIkP+M6wyXuc/2uEJh6gjO41Lw2sHaevfgMJhN8N
AmXt0EVteuXsLWGxO3R1L4CNBSz37RjiOq7uJKM7ndg/K5sRSzvyqWSg7K0ZYGx6
cpLQ6BW53VY8l4OdEAiKyp/4mXMQU/IpWV06JSX/RQ3eUYoc6imtPNGcLf/NkSCZ
cXyecOGn6XnFbwx2F/r8lMmOY+D0g/fmsP3aV9oZc7oSX7wo/ssrGTpfQ95hkSU5
6kYLMNOTCJP4X2GBhn9dcva3amSX6QuxCBcR8lQvLuicdf3YguyaYUUBzEFKVUs1
TqWfHP8hESyRuO/A2lBzbl4syWqzjHMEm0p/sf0RlNvxh/p0oUOx+/x5gPJKCcZG
ElG7kPjJORW/OifujG0zMwhkmjewDVWZuq/yiM+lKj2ifTnTfzm3OLbscSQts7h5
ITteF8bGgiPJ6hk4HSBpIvHE+LO6aUNQnkMh3Tk+Tilfc2ZM0pc2NRddNQJzVflx
pRYAB+3vVG4wtTCBlPNmCPHctE8iqMhoYGU0Ielf9D0D8cSbYNhk9lFmQrHyZHMW
OuASvnazmzv8jbCffVNdWxPlvn2KN4KSy2F4y2i/nXkgn/awGDVH/lKqBpuLg3g4
Ai4CW5n679tLCGr/eWagMEbSuxWAv32yCZnrR6ROzYDmZI+GJsBAAA3c35VBohnX
1uLcA3qLgX7ArwWbX9M5IMqBnynee1x7UREb9nlkzikKUld+P3b4/MNnO+Yu7eWW
efOzX4F/7S2iZit7nqpXAq4oXZALtbN8ukXgn7t4jBEfxz7uedhVTO7M5KiLYTpP
73LcWJ3ai0+GxC+79ZTxKOehxmR9Q1N5s6ApdcWJJrI=
`protect end_protected