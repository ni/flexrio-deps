`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 41760 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
ZIICkMu+S2rq/yOQyqhpupJbVN0FZ8sKjNPKoTtHL3Vfe6952VbrvHsSHKDS1mqO
Q1KW1IXEqEtz821RWX4vTBbX4FoXLSzijLAmfUWUoPuZdvSEFgmWTOBcp03HumME
RyGAA8TPHaNLjnf3P/gnc5V94cndcOlhBx1gfjAjJnLALVEcEK/Mq672g30lNAnk
P4SANEgIxSZ06P31Vj82DrawfA3nmR8FSkQD5ZX01Kc2f41B82TgxZTgQPHzsgV1
Z3+a21al2rVkNTbg+LSw2gDQngeGcPUgIUiKNDO67PtGZaS8SBhtxTa3HH3lsfZY
k2ZmQ/+6FW8FD7SpZI5rA3G7OX+wRnRrq0BotZnVEwDjy7zVNkazZjKGztyXuhFq
Nq5hi+DiugoHe8SlsZS7LcPs0+DOw677iLV4BQk6Zqb1mPhPbqvXlywf2Bci1+qo
ni2xxTOzZJl06LsmRMr3K1C9wvwXe4UZpvGGv2nnlT7yiTFkJroibyL1sd9P6c8g
k+eFZtgZ0QlUGprSGVZa3lzmW7ZCBbribr1mZtjfZozwEzJH4odaZozkMLUy0lm/
dmM9Bq9kDK1erfvGddXaqiNmn5M/q7un7MBxFo/kUKHq+yU19TifXl00+TNKysPd
uOBNmj/9ic02Nmf7FFp6VfMp3Mp+GCYQ28UORuRzMJn7ma5LQrWnJwI4Flw5dowO
UBkwhvWhunku8+2ytrSdOwV3rEqj/0iHMiRES9qeuXZg4YuPldQm88O1AkT5kR7S
qCiWlbfazFye2MgcgIqzTzwPiKqyACev1R9J90mfcc/5QYsLXeJ9B8O/a1GHaA/3
OHSF8RO4BPx1YScnu6pG/gKGhSG5OOirwQGoXKfMqNrErMJdcexTJh8v0MBAYyjI
jAYhRgf8FcbTlKUrJr+8EVqwU7z7DPC4+f+NoWNmtP2p1asVoKU9CW7Bp7RxbRRs
AjOcbnIHE+6fO57Lei8q3D6lOnHBarJaoKFHBY5W1KC+qzJKnF+BA+jCXkS+Wicq
6Fb5+Yck9ZsL1D15n3LQrOgtfoTFCjS1mcNX3/U9ffLsLveJJ1gVlv0TE0fLfG21
QJrbxS9VnaJQmny+vyLRaPIeC/wJbdAEJp42R+AD7DFwBRvExQV3sUek718e8mfD
Dxci/+IZ1To0chEQOqtWk0kCMJ+FxwJMyKlurcNqWDfaUDg5YSJ+btuUUQXrSk4Y
4OzgnB3RSAIYwzHiwU3AgExgVcPZFK4Ne23rtG37YScW21f6FKYBbsAPsKK4Tqu6
U55asXDLcqcELrAWr7nwyKwRSuuI3aZ7bJOBto0fPK9s4aREm0qNsHVP8RutTT/v
IcqpD1XQl0VrH74gp1hS2w49paRfnH267sputc7ZrJJ8U/A+IRuf9I4wJtDrDQrG
EarNF6QXO5uj1nHlLLwxGfCkr5rHWMtuhs/8q8ytlhLDFUfz8ErfYc+RyBVFqbiK
/x0cCblbH2hNHUJFqZO/pAyjtnP4RMB32MKLZbmZsAD5ZBMR8npfice8sBjxvQmi
HaBGxB0PUat3DLvkAQjnimJgymHKPmPbSpgKcQsGrzls3yj+cUfi7Yr9/MHt5ouF
qEL2uauwmTkHnfvER1RC1XW0RO6JVz+eX6QRWs6YQutogKOflJ3uYaShHZtixL/y
KjZbj7tZxxdOzz5WJ3zJx5P+/YFmZ/JFT3aNbQiEHM+90Q5jY/XyrhSKaUDr0qLr
WAMDvOk0RGdEabM1jWuSE6h+++fNf+jwoSbXYgWFVumdWcjq+PDdkqhInhbRvF/u
pydvZHHLA3mBM8gViZ5Lv4Kqq7FgZtoh5W0x5RAsddFdatfzEme8di5bBB6vMQrr
VCr0vF3zjvfZI6V2lYBmu4nMK+3WwFg1LL6P8qK0hN+1q7bsaF7CXdo8E31YBgGm
/sREczprjw38xQg7YIEEsv8ItJ6uzobjxVIkOjJp8snfpD1x9JzpqrWyW0DQyM/Y
BhASMN2mke7qUct3rS/DUE/g4E+Pp8WJHITjp+G0ofCNyBEz3T5VCYTm8sCnutA4
0uXhTMlVM563LB9CO+WVl68rZBO2UOamNrzTcH88jwZvMT3q1XdJdMed4yPc+L8K
pB5WKdviqHcRdF7odSRxrDSJMNyGi8u3g7G/L4BqTRT2qzhq/Zbr9TfipQa4zZkt
3qudZBtTveqEhnWKwM43rtX4L9sjvKAbEjy+KDm0khn3C5aLBAS2CBqzESzk97UM
9XBYJY0Ye+F0ZHj4nNrUw4uexQT6Wn7NvSY4cj/YsCQIh5oa9oT95UKIc24zcIBZ
9hv33BhgeNaJSm5c/Aa7Aa3J0HSCxlhof6nz9pmIrKQt22HeBezIcl0gzrd0HrtL
wNVJLIm6nW4R1IgomjrxgRqdPy79AW9C1m7gBIyMreARPQsbAoHPJSq04CPVuAPR
aaJPcCxuS0s1h14X70dd47hHC8WD+0MaRSmfKXfbp8O41mkKlVzdgbyCXVUeHs63
0EAer5v4CM183e9HszC3zZOahID/rVX/67m/ki90srJa8ygqbH1GJEw4vmHHxgES
GUm6Wn1OQgJz1BW6WunbLEMKo0SxeLwzFbUpfFGJ/dv7glCXxyPYdf8csCtsLQ6T
bseXU3uMjadx8JhwjEbpHx+TFYaBgII3zK0Ga6U7oSeSaSQAui0qv0ixXJEPqUWb
Gws7FbYN/PeOoTCMR94jpN+a1GPMMDgszD5fEYLtHQTAorPcLCDVXd7V/3gpS3Si
WI1fvg7ZKT4n6LJ8pyy0VWSAmPZzydTKOkyLTxouB/IK0I4vXjzKL/s5vcc6oOXq
4JXd7z5XGcq89ZkLx/nHbfnhbLBWq0xyhTO9X4VbPshSa1cTRwzCQ1hkoTrr6LCj
pEDosO3ybj0xqF1EIHHeim/UX79k5TPzzugl2FXdUHMPX1aKpbvRvbbFLwTwTHj9
/H5IPADeee/7umy/I5kdp27awd0XYtpLc92OsERHE0/OXJ9GcvCDMFO276spZJfv
vCA4zABuLABg5G31LH4kLvwbuKji4vlg0iCqxTdZtzVftisEmNVEjh1kuZ/jjZ/t
khSl3JMtKVHpk6rTS8VQgUob1Uo6lCjy4pCQw30CGADtrkhU6QYemFegHBHmJQKN
vxwXeNYBVGpZq9DN95rLXqSnvwjZC0FY7W6pjRuSxiQeWUIrgdR6UstQQuvj4Ntk
iwhuX2rIjM0SRQrJlDWzYwAVoCS9jsdnXDESXVbnncHyGUdmN1/+siFJvCBlZ0yr
slVmFFr0y2FBEoTEbLOibuhkSBXQTkrjjL2hO4vXcUOhxVvLpYdJH45nq2pDz7YK
SXfiqkaEJzz1qVlMqWm5bJTc01nyTNd5UAe5QkejGGUmqzMBWBlMpDkVCe5bN0Gu
enoF6WQJdninQWgZkMLBbV0+h7moxBg3gj8XbrV7lPcu6i0ZVMr/CutFnIfb4etX
qk1598hcHDTBuo6OgPrmqfoKxkrzsuXdWk3S3XQPEUqHGfI7PYfCIhAOJ7vSWHKK
bRFBwuLHxm5yh7GfBuXLabikIQuvP/7Fo9rDAlFMrrJb3N+HTNCoeUztErgwaujs
rCZIpVa3oX95/XlLQ6dRUbClnLn2TGWE8hDTEsvKLP9tdRg9ghooUqZ/iQdnUmWB
ZmEOb4Pkxkli0sZGVeDrHgRYRPZjUED7o9Xc+LrDEhyA1psFz/7EbjhflVOopOJ7
QkyP5uhpf5pdx87zsHSUsVQoiYNcSRIrPU8L8PddFPTZCnKantNPPk2qBdyS5t8H
u5xABU+I7Zc+LV+HxmBdPo6lnXCSNmse3RPk8mMLVIxoCZhbTrGgPdruixMg4nDj
HeRkXfSXftu2KGeGUTwrB/7lrqXTdrVjWsgLYUETh5ZKnzgoV+8eciGHJkYa3DpE
e9TgJFOHGQbLxijCr3hffhHSggy6ZBv78T42BpsHESEOaxXeyXaLyzdwZXHrdVNY
0D+uycd63m4KoxCo0643jNqeuD7VcTTfjA4gvJ6NHzZiU7P2qDC/tm1tPDfK6y8G
9yepRoP/Z0qm6yrwp0scYt1Mfln5rHUU87aJXfrJBE1zthQOBBhyzcXz7DhXkO86
3Rg/oSxyhONFgGQN+6/AjvxpFlJDtBLAAQO+yAJx+Lcy6KcoRWj+lGP/EXtbXd/a
BWPNvgL6Jf1g5GaU1zg2OepLdAijjA6NtkXGr8jf0zIvQ2CM9WIKK1a8JhxqQ2/k
VGbPIFvZIpC0HbO+ux443+6qXVniT25eOcT5J4JryxDlKGtyRkTm9LZza47ooe74
vYeglz8eAXnOIN2EOKwiiEga/USB7YPqHgKDNC8C3HKufjNfb6/OUswziRdR0qGu
lT8TW9c/rQSVcKSt6AOIlqULfYoSbrXIrsIjl4sM5FZcApc4w0s/Tmf34t9I9ZE/
T469g5N6dnsSb4YPaWWJqHCk90h5jl1dKO3w5IDgy5N6RMCEG3NJSBQ2oQ8xTuvp
bV30z9HYN6vlekbUXrPlTnF2VqeyvWdf5OSzf37/iFnJ45DQOLisCdnj7EU4JZmw
2Lpew7g4qBlYVAft+Yvl6Y5ZN1Z2rItoYkMEUrqwhA+knWVgATWFgSaI+jUg3wXV
GqQt7K+b1zv4tubem7m13aVh6FpX3AJoPYIfxZe0rJ3K+WwR5lAxTlGjh+cZoJN3
X6yZn9/foBLkHhB+jIwVpVg8mJoyDTpgEA9YVF/1pWM0RB3QaV4x8zCKVjdZmtXH
nZotGT4cg0x2aZ3q2ThXO6ICE4S4hu1PeMkLZPwSdWKnraKJxlBnF+4kMLFXYT4c
uUi5PKWI/Jjo1cZvvaXHl7YwQBoxiihbuWLItYnVvY+DP9Fcu7HbR2d4GADPAgj4
CEGyH2+P1/1MwG2Fl3h/ToO3tHRi6sfHHPPArQTbVbxKBqtOmnypqcW3v/ukrVmo
QDvzJaLMxg9B3zEHSVxMN3ONtNrmAJVtaJCgYQtQ8eENzQKssfoXpvKHzbqJdYfA
1cDH2fw6t5VAUvcd6zxyVmODmx8oIYRkXBI231DEv33WAytXf4kPg6Pdc8bAQERW
sw/ImlWr28h3DqFr/+WraZi0tj42xNDq96CQiJUZZQyaMf32ZGT1Rvscnkt0uoCa
h34+033t6M//wsBxoPE0E6vdBS+XQ1ohMQvPVmCJApLgBu8RutsWN78RgSF82xfR
bW2zRx/7nR7Gfy9Ulr2pXJh6H3xGRJyZZ1rS1+QJaRm6i9Fka1cxLWVhdzljipV6
gPcZZjHs5O1AED0xufKAvW19V82AVxO/DiwTQmeYp5t39tO/w+57sE96sgsgFR0Q
6bGZnxHTlL2oWYLnRgixo/jaZuY1XhbgT7if+GicY8VmQtti5ukIEpduzbsTeokN
hh1QbFotuRyk+CmOAz4s+7IKUvJDNhfHjv5w2dbQKlRdScYZPhOZbs+sZBk2DyzJ
xPWajO8sQdwpxVTxIczr2wUU/VoaX9TMQESYIyvzj3CzJDjjB4R9Ec+hWxQmjc8w
7Wf2l53tN8sezNoJr8HVIG9NQn0VvJDHYxr0t81eGOEno3MMpCMdWHGvARjy8PtV
HhrxSTWYuBfFs+xCTNqYpR7U9bLozY3rYJYkJBfemexjZuAOizCOXqcY/nXliImC
P5xUQUWGEF+D/PDxh18w8GJqQ9pvOD5G6fi87sYvU8jqOIzqIMctOga3wYXnmYdF
0ihvyjOyIJxQZfDUwW50GVQGbbpJA/6z3euCXaVirTimMqHDmGEeT7nzJQxB1aG3
+JeJOb3TUS4y33Rzhw+3qKThIWH+4LPDETQnBua8dPZvFDXuHOAuDyKG9OHWcHas
KLINRfRwtqHaOM/57ZBGTjx3t65VMXv0cGvSRuiY0GOlHoZmmwop2D3jMvVD30KX
r+yZ8w5B6zwOsdK4KW/CN+HwQXpsLMwucWdOdW5i6xaL91N2e2our2y8kASLDwDJ
gvtvOHZ5NyM14rdxaIV+VUi6Bvs+qgGxmQCdRpqpWr7qBmfLN1cwQuFlb1nRltzT
gXXw4odIAua/5+OC+nZ9SIB/M9U1lW0TFhtWAAnQAIAqfr8LINKFcS7OwWr/KQxV
wAJA7rODSUn6R7Oib/9V/XmXvU9BKtuwIYQ/zxcqsTadXYTNMxAb/0lMI7m7/fnM
TvmSVg9OFukc2AMHQ5JSojib4aY55M7Fa23FD9eqkWF4zrldhBnYKQaYbOH7r0x2
+7HZDfcK5fb4WU67R0ES7ef6r+QMIqTcXwGoLA65dHaUVuMJmtinmE2ppv8JEFfk
vx1jiZieMpRAQ620ocskw7BHBVXQJh7fVbp/tMogfLc/a+jIjaB+KmghYx7LGzRE
KtYNyxHB2uKOBi8n3SxX49p/zPybWtmrnMC3Zx5oqXSMotADbthzOSXNqnzrw9uD
kXUPQrvKa44kM1efu9cHrOznSB8CktPFJYjxeCAeSxS3d8uJ4IcTcysAguuLJM0W
ELO2ZPmkaz6hWR9D6sus3bbPAaUepBCBORNCnaeopvBp4GDBcvoCScmzX8QByQcz
nll2jIGZjF/AgKrNDZHnpF/n4KhfALocfTWPixvhaih/BdUA786ObgijHjgzn+Gt
+L6C0WCDZf1kDZnDAGCmChPBnOREV4bBhTw96pCGdK1uYUHm7sH54O495pw6+58w
L29k3WebspTpG5xvRLJKqTMuajQfUiYvSZFHNNevqbS8ejxyjXuVRBHrd0SYleQH
npGT3mok/A+uA8vPS99mypkpQZJzgxShbyDwYndyfh6m/gTmwrKMcrobDEbScEYa
ed+1cQiCsboImGRhMKu0FLK42i+2vNGr16zpTBe3jQAdc9Ydk7HBK7ktLLreqdxL
oW5bVUQ1vpaUZAAqRP1+49G4jjxrtJqnXBLy7+wmioKZeQtUu4gwkTfVcq/t3CKC
VLoMbE5dGy+CE0eyVI1kKdw54K58m6qBpDBEjsvHreTy1rE6U1BofLcDsDjBhYYZ
VGLtYHMDA8rOfA8U6PhMtSJVHLapSv5hXPnORmMoTNx87MxbD/R6B1rGX//Y1Boh
CuTrVVtmBpqpuAjoJ78x+CnfrYZEMEmTaD0oN9TulK4aYJM4qUgiBOw7cvwPCkD8
PPEodA/pr3A3waV9XdNk/XJSwy3PS3vyv6QgCV2X/PvX7kEK8NtIG431xjzQBYSb
XWoGHBMQJ2E6pP5nSBEogH1+dhkBBdTdW/7B4H2zo3LCPBPbGIE4hP0vXj0BnzLf
m6Vx/DeeigIfucZTPj/9YNDHXrU09MRYe4GMmBZeBFlMansC8P6T7Ga9G39PbHiJ
veQ1P8tccAjFORNt1FlpYy4aT0NlRWTZh6sggC57ZJb6sF7ajTeBxh2QVZ/WXVaq
WWLyi92BcmzeqtR6GjTCWNPF2245F5gXC2Ru9FJmPSvVbhxXB4c3tGR/GIR3F201
Y0K56G7ynLkxM+AC5SvsWvHJceWA9rJAhJq/bHOWPoFAINnM9oInFXLZgmc8ykPv
XU7ql2bUw+5sBOaRBmgJSCsoh7VivUXzYvz1/RDIL3tpiRfa+e07M6jGgzmPnHgu
APJFaTZQ2pPLxHvRw0E5uY+kBOS/gDgDdom6+QvsnuijDu2YiQdCY5ZGH0+liOHD
3sLvCHTVhvrmqeR/XDbAkoTU27l7Fah76625tq+WMJGuKOHrFvnyqe5zsDgc9O3+
KsfJrWlB8zsK2S3RMXpt1kWO3XhIH4sIuqs340X/AvjhbdfyeX/gfd2LAHTlZccI
n4CHuulVO7xAHwVsTvlKvWGto+kw+7PX6K4Fj1FRoSV5N+aBxGqWA4aXAuVO32HT
MoE67WCLfyRWcQ0aoadzhn6/ltXI+lsY/MlaU1xT9lci3e/XprwDSW0LmlBtcp/v
+t/O9m9y1ZIaxKAaw6nL+rVxEjC2BIo+AvDOWNSwr5hMTJYZOBuCMQ+dAE3oBiBL
ia+W2+BCn9z4MI+GoxrRQvOsbPpr6aA7giWk/ocBo+yK10DP0ZeYUSRN6psSHGR+
JGbrAEoNEgCqhJ1F2Wg/6sGJpKTvz4QMct3/suBt9L984zYITaUeT0MFAVeeConL
gGHgjEiEHSYLnQxN2BO72+aCqPOXekDjU+UEkd+cosBrSKKxcpq0NvBEEw2oVH2r
c0hjAD8DsWIBUXwHiHx2NSpVGcyszfpxbT8qhg8U5mnvgXKuLspB27fPqLNMPuHB
NocfD9RizPmSgUST0NDvTsvzCKqon5VosJhSWhgtFV/TFtkK/pcwe5coW/yHLRUQ
1P7DKiPvO+0sqBFCdII0DbYtP8kov4Tvgd+8kpRZgdyAOh/hjsj6mQKuibHq2GCu
gL4q7rZyE0laZ0j2LJ3m3k/GdFQgrIKcL1kqdmLFAU2+HGn2ysNgq2OCNsBNxNUV
DF8rBaHcMgeaTp0Lzsmq+++FnQMqLRPjz02BeTv++p21y9OdQwd3flj85hlHmstB
z/euiNMOOayLOJBc4VCMSEVBw81p7I6anbDHyFJBphwXx2UReEgBMdj4s5qdDwUw
7RDljnyMgJQ5TTMAD7JrqN2Kg3gKYm6etScvtzRiCShFYYRt8JlLVBHaw/wAwofK
d9DTdUl4Plbry/5ok8Za2HwNRLAjTi/DyV0sL2JSxLbFl8fgqihMn+cszKl3SxPd
8/irb43Q89/OaQfIOEQoTu9Zh8+YjTHADtcw/c3CssTmv6z52c8SIpbP5aYHE7OF
n7MXJz3KdhXv+scJ6H/PVsrqBqEYgUwwzFXTLarHot9SEgs01n2xQ04qVdoDwqcq
5hRn5yqaX4U9j3n+jfVs8be3Rbgt/LU3O7iXThdgN7VrlrBbi5SQSBvI/Eij+1QF
oVqAuCdwWP9YMRYcf2b0DVwY4wPs6vtvk89p9hl6Dvua3+z5fBUEPMZkNhYdEIhI
VuzoGsMNV0Ij4YC0vbtg0Wp58NtRGhj20LQaN0BXRiLKlaXPIcLlJGnXh60BsHWe
x7dL6EbgCGB9zy3YDABW4yvvY9vpNK9eLvJ40E3dRcdHyCzFSTS3h5yHIIe3Q8ex
5HnWXJZBt+l5r5NM0Dsq3HVLDwASI7rzpG7fl3J9F5SkagYodL9yoCzVtBE0Adkd
aR8hd/L67BuTo2kAB5jBEurMUqJIFqKq76GNLYlFqNmOp5LJKja0HYGowLYoPqJO
CdGN7iZsSDbOv73ty0BgWiw3Pqa1GDLgOttocA1AhR+1uZQXxSx+T6YYX3HODS4H
naYznMfj8+lfBgd1+qaW3bGcK+c7bDdWmqSQwXlP6dE52g0Y+gqIU9TlaAXu3uer
niBk+yvPBJxqKJ5ZoS6wWfTKUYMLiB3ij85pNYsFN+VyCQBY6KgDMKHJ84sZ0WtP
r81LV1ZNUmeTJUuxaLbfursMFhkdDEnBU/1nDvO8nj22YYpxUOn8olAX/mkvv62g
oAfejLgEHJ/SiPtpar9CvhKVs4818cr9puVJDExcV5vwU3adDdCxznVZLdAiPkG/
3iqAh+tqysVRg76+RYDk0NXuhUmVPYd6IEEbYQDeo6252HMadMvgAFNv/8Yoo7Cy
um1NhKlAhh/8pwZ2YPjwV7sEbsrNFHFA3pN9Wh3Je+ItsrKd9AzKPbLONJ7t5eJw
JPU1ds9yBiyhgnvRADV4k3WGBm5OwjQTIZ4jNdfsoH8HPJB0Iwd9RscI9nFWi7oc
IxkmtJEVPa/W3VQH5YkcdBbd1q9HiYnsMACKD2A43MuSg2Wwka5J6rL7TQd6uSX7
1B3SUiADLE3q3mlO3zq5/zjieVIH3GaGiHOrMAEFpb0EJyGCOH+dWFX/wBDDL+dQ
2y6Qygk9VYr5BTKMJBxUy43zdgYxY1GH6imdSph9aXR2QAfAEFKp+cpP8gSzBPNq
8VpMlkZE4TjU1xUrmzglAOOp6qdEsKNPt9jH5q1D3g+lkFylcVpmlH0J2MuWMVnm
yQooOCkUGvvrwYX+Qz6Ike/KvhkerT5aEv1bQcxffKJ4d0yIYfWYuTm0SRSCNKks
D1sdxKmsgvQnKkkSkdSkLZE7U8XcqFppXqW10TlNl2qTmaoTlD2DVn4wXy6KYIlL
Uio8l6rCy3T0GezWYm3u7VEyoHTy6drhHZy6J+z25WGhhzFZ4NvCV6pGNAJs6Vwa
HaATSiw7rdTfgDF9pmUGcNZiuh4N7NmtlHn/BXo4qr/mX17COe5KFQY1Y/9pHrR5
ppCffIliM5cc7HNdmlswkImJ1GuNsGKChIbP7niabjGYlK1l6Jd0ajY4FTrJLyyw
YSyXcMd7Qw+7jLbOSMWRNlxsNvLDD+TxttYUg/JdKd7AEZuLzFkKTc8zgYcfmmPX
8q+JfhXpwbu3+YDxMr1KQT5Xm8ENnkcKj6CN9tKsbJ1W4EWgeqeVaneQcRqMk1Ft
LH8q8ScekThMIBcsD1YtHrMPt9/he1YEPikXRVdnG7QsPhDTcdGTk1CQum41PQDE
rNxPvoCysUrcMlwa7fS0XoOR+0FzC0/q/o0g/00GTsrjoZ+kyvpcPLFGePoNHVkj
MunLWOhMW6EYkk+CRJZg4DFNlVCA2n+XOpbgQ+CRyrcFEufvuTO95lRBTfXEz1Ij
RbHrrOOsYNTQDRmPYvQbhhm85xlStb05iz5yehuQLBtf5aQO1zyTRNZq+92ffv3g
mbdPWBmqAIYr8mr7S1uIgNDXt+RMXarEj3Bq3h5mCrIpuLZJEkFyvAmFAtTE9Zd/
al9AP2E/LwOpJhR3/bcUH7KjJjGFabIw7oyH6WljOJcNSuL/9PPm3X3XZ2RcEztz
GAWHiQluWsTdZzE4d/H5tQhYjdpGugTmTMZ/BIUXVW4aHHg8M6ZvASf0TBW7mLzp
H2rYxrAoUUlXRW3gfDzKfIrhBBXufe9JDAeqxvIsu2aXUWuWbxpRELJGIjDWk+B4
6Wq7Gd1XuYNoQVfjPOS60wl2tHx2NtZrzIvSbcOR2joua3fYvqh/urL5OTrnYOi7
izLEtsTMC1KpNsUgnvvw0pH7G6FfF8E0DGxN/Trrq7wGdaRZHx+kIwdvz2a35QKC
fBbrjGqfMrCmoXkwiQ2Ps6u7kMW0tKGjNcQF0bKRMiAYH1FnzBoD/rY3sMCd8AN1
wBp0SI3OIs/W/UKIEw7OyetKfcOx8DkaGr04bKH+3naYCpcxjvp3NB5R5fJVndMW
dJdiKtX2yYKaDxmlmhO6nfJSn3w2XnP7CnzEs6vZFJwucWMpAiBBfUusr3londYD
a0FIxGo+88k26pPNFb6G2aJCovCklIo72uaQ4rjKfyyE5EHNVKmLGG4PyhfJkV5T
aShdTS6nJglM50FqagE6XypuqMJyjGkXNJtYFMxBgTCCK1yYOeUXhjf3zUm3p05F
G5Aa537e9XzBPLJM9hNSJM1l9NvMuzoacjZavhqaynxyGalpjNOOc8XsohuuR00R
o8qGLb08vusHlvfVljoighLmh6Gqh3R9ggsTlO78It+vI2XzFFNdq6I/Drysb3vs
FqeZ1HERZPYTqcTpzoqM0LENRH20Md0mYOP4tgo6eQl92diG7k+V4gXeVe+NNf5x
eJW7idQwJeAmkEVsdj0fZiUG3kVwM9BR/6LL9olZJV3P74yPcIgG7kWV9p92l8z2
17QQgIeRHeZGM4mb85ImGaUGvG3I2A3ke5JTrpNp3gnA/CHwsHBPvrGALDuTQOYf
iBz95Qh7GVear1fGXL7qr1L5NGsBUKYwvyOcehK164I8+HQatWQawT5kKM8Tbglr
4dlLebHFkiup3ttYSPgWe1FYZEr5sjiX46w946xdk23nWjYYhELqWdFSm7Snj5BK
CNRfZ8aqKNFV/r9QQwLRXADrQiCfeInb9pVw8uvCus/hvsBdPtRNt3gNYLXJp5Bv
/ft8/AhjbRsbsFBm8/rQ2AtZ6oyM5veZk/8Sw4/EojfX5F3lYzdDbVMzp57c5fK9
0riW6QFO8CVMyYk66Sv2gpeBl+1uK3uG6MUQBNlsKbXZjVvflBvCy0qZKp6kMlqE
yReLRYsEayil18ZxFhzCa46ib74AS5dAo78OURtEIPAsAFAEYlrt2fCQdBQBv29x
CWMsFZkvjU5wKJBz5EO6v2vTd1CarM+ThVZOrtCPLgkNyFwLB2xuHZmZaXTnhid6
g25s8ImyakqVegzh7YHXk85jgvfejbMKBfP7Kcd3pnuE5pC+clAewxz4NszW1zkF
2gyduxzvL6p8YZ0IitSVJmgJByMVaEROQmvUWqapU3QXKYViTqcmLkFLYV4ttjFn
YSxeKymGQP3xsjWbdaC3LERYQ6oM2AYsvq5Yn89wnmSX3nJiExVcO6TucAc3m1qG
OSXaqVMSPvmxhuPnSK4L5O5ItF9DrSNvaNcbv6SDginZO4nvrwaeRiuO8s6/YnGO
BxV/1eCtRxf7062M65gIzQ/aU/+xHylS6FVuTSzEJPYmqER5Q5SWDDCz8i2a0Sa2
xRfYDvPY8Ak5196jdQgFYYB8WvYgdMVq5cYOACxFHat5zO8o+Wnx4UykWKT06DJk
2ICk4MmA05orkTksVxvb62PI1kq71fw7il9U5P+qP8eo82vAFmRVehL6HhvhRB4r
bBIzdZ7cU4LR08VFO1maiCw3vHKznGhnjS3ttfPufDv3uFi7177fsjf4lnAob5r/
Pow27sVzfapzgahZcqF+tSOLOpFnEmcExaz2oBO73ThXk48tUNEDruyV0vfCaZRL
PkDaXEAXBMOuje4UUSnqdhXIXjzp2GSaG5FYh9uiJW+o7y0IjFP112ng/FhLbGi0
mwI8RLG9CseoXhKWBQvHssj3oQ7XOW6hAHyzH5P/7conRkX02YWneGc2q/m2zNX+
ASlw8PS8Lq+8oFpSHYYSRC13ZW+CuvHUAslajEejLvHr5LFiRQyJpl0AiLnrx/yg
/0AqqGS9JfeCWTMRGJqm+wjW0g+oB1YjSz7A0f7x1rRjL+odUGJfMvuT4OjvUiTg
rjb96IVJb4DMNWPaiWTgWZOD4B5wVPkgnaP9JU+YCnzcVIO/SQlwCo49aOVYzPCN
cJeUIlbRWUHa3Yi/PEHUvqBWu2R06cb7bxmI8cTVcgSGukAIS0ZTMEiPxYfE21/Y
iGuiBMWkA/dVUXZSq7koaWteTxfwvNg+eJ2gemmTXelamlBiCurP7kiFGOeSsFAb
cBcNuensLalIzygECgYm/teGaixsLPI+YUrM2F8EjcJW/BtAw5VBg1F5BH/g+JU2
7UJQmouPnGRRFTZd5CCJgXMdsFsCgxXoyHh/V4TAPm5oqud1CNfgJsExVZV5BN1P
UsZdDQc1VpUmWW02XARbkFyBvluU+ywrAT+axU8qqiIzWFitoQUDtNgoGpYlaISn
QtkAEYqLaqeO5iaInIHflE3H3z3FdX3Izpl6dKZQcNAQS0zzQusfoX+iWfVnI5xD
8lj0mMVpR6Eh2c6jEbshrwIzEl3U2havAu8p9+oqWsE01v3x4v2KMOEkFC0JrfvK
QY3qNG7UcC5x5wy1ieBKxuTBLAR6kjyLLTj8R+ZQHa9urg7D7Caj0OgQyULHHmCR
HbkCIltKr0N5HL9EQRris64Nxpy0XsWQjqRXZi84a78U8KEqflUF+IJ+VzyxeACk
LUTm7HiuRrC9UH2rVu5/xhLVtaIDQWKFmPhfYnbM9/LYlOWOB7856ABhNBiUT+I8
OCQ0D0KwnJQmWf9ampX3nYMaEo3duMwDTCkDPJj3bTc/BV7QRV/651qBnXDhobtK
Zj9fVuK6wIbYDdfmxEJs8tSHVRmlppaUik6j5XzQbWOyag99337bjv2slMLdhL5k
HC3wk2wDDV1bIYWn/n5GOdvMlruoISdjXzkPOeQfHQD1cX5jOpAPIq1bNyrylLa4
ZpBTjQE2icjAjlS8ygrGJtksxBgH7bruGLHyf1RS2kyyfDl+a3OQNyceKqWD1UOY
3MpIiM1y0yRra+OsBWJpUqFmWnkTNWFOfM0aluWePovaN6IDJm0Lc/vI6vW1bIDm
RiIaVrK9DLvSoKCp+MtUM14DXfuUTtVOCDEBZbhfNna3g6kOi4BxlHwZGOx5KxLu
ahx4fzwfl8Cxyc7vvGjPpjZ60U0xOGbTeCvixNNP6/oEQ7oqTzfWBWkZ4aFnAHj3
3TRzJPX4ToNrkqUTWQjfs4+E5EkUoJQNGaab1vfwui8wTfPiJmlmHEKZsIjctF6Z
bUaKYfnvLRrZFxna/fbQut+iV3vTCLZbq+/D9tWAsApiLqa048uzz/V2II2WtteD
rewywDSboGEPruNPBiJB83XQX8u0zoMeq97a2kxY9EWf8IooSKs/0mWfkJPLoYsB
ec5kk4idc+FFTgIur933KkJ3yiZh+IXfn+4ll//KuxjBdONlQxsGP4M4LRvxA7Hg
EwzMTRdUq8l2ujgLaoQFIWOfMpdgU7g42kDKveT29RraYZ/+V0D6zH2JBDm+ZVZI
Klf8JoDCZi17GArxi/Jwj0xqbb6siBQay4fEbE2b60d1G7TVVtKwIv63DVTp0xZL
zBa9ehr7oaQNI4x+ujDt1dFFitZhxoWZrC4R9BSvnWNRNTtLUKRycRWnZ6tt9xw+
kAQOL2kxmUZBNV255ShwYxtJyoGr2/SQlTHjwlhsRzcqj8ViT4Y3fusdYEz9H8zE
/LyQRhZDjuDfXD1adl5VMHlo+xy0G+UZrm6USKGIv9C3pAQR1ddt1Te+Afs2bTRN
EimF4y9l9q1u5H/csHvcBW739u6iV2mM3ifOna1ZEWOzClyjIE6u+qFqVNx+pWtW
RtaCTjsK/HVRFjY04G+ws7cgI2oa2in+/aXTxsqDWfO60pXd7uaUY88MXloxlVPz
EbxEU4ocflKiLY9jC6DXdtTHAPC53TwxXUvQAKQ015Kj/I9cWdg5Xgxlivf51hnV
Z47KGMCsyq9MFheMtMSG3r0+uEYRHJ/zL8W1J/o/XHKXkPo0OjO5Z5JfjcFotmJ6
EvddxLE3slqHTtSoo8LKczMqErjsjtQ5zyaWgWZJOndUY7cuZlgS4N4n8cP29KNx
YbbOL9dn51FraXDrOpsNtrKFdTU9RajTRDcSviIdI7JrKJbF8sDSshDBlHZrVsmo
BlJxfHnXX2TzB+vbO8TwHSjKx1xOqdUM6h3tYK0CBbLL/BmD49RKQjPUQmkD6Dit
o3J8D8omkU+mQA7b3izUkicJB3X6YX0gQyNJi2Yltx1bnMMOTBE1mgDbd+mFdIiQ
lpYpj1tlC5gLh0GcjeI8AnduUGFYVKJn8GBS2kZkbObTYlZJfFXpd4Uup73HzwzF
P4SF/r+XerVk5ejuyirwIN2MNdQMD/96EEKITmNA0Bp5pCKdUcozvtB94qhx2SpN
dGzHdlOCy9mC/8GxZ8/pZ2lImxPpP98WOusB+TC2v9G2MLWW1pSVLniKh+XGEazX
vfLVIWHP3rMU5vaCXTcV62Jib2ALbGK8k7438pNVmhl+sExMWInjlwGzfQRzwKUw
Fx0paBgnQyevV8eBWcwVIgaXa5yMB8RYiU2FsvEDn4DV62OC52yAY8zVfoQa4yU6
Zq2tw33cO74truWNc4G+GHJuA1ol7r6GoLsnq6IM06IE1BT/HKjRx2ZBITv4/PmO
Ls+QoDuMrNqfhJ0EJ5EEHPVdj5Us7S6ViThWj6lF0egaJ8AILH+vr3p1TPAG9dAi
xb2cHshm+AVUPrXC86O8x5WS0Zu+bnt3yjIw39Qaz2/iJqiZigWSGAPs0WoGPf4I
N4elzarFl0XrJUHTqJk8A2g12hOKH3s8BbqavbzakIW/Fom2VDUwKLKyLV8cbBDc
1Xs6ERwW62SPmAT5TfM5YFb00bgo3uozDSZJca+sUtNaM+juttybLvuA7vPxDrr+
KQr4RwH/75DKEBr8j19WPeeM9Xa73VgK+THucEfI0qdUoRT8vahw14PdyR16vFAk
ss7JrTCM7PVb4b5MzDMhDKps8rFAgb7geFInItJs6N/ybw5rQ9Z3KbEctTIs8nbM
gH5MmN0FenGwhzHyM+vzhKax7xynSqKPu5foFCWDKJqUeWTC6MZeJ+F73wXiIXPg
ZI/PsnFZeswinWY2Iwcsjxo44HHibInjE37WGiYhXh+emlflKQpvB8izvRhoapSP
2hWdvKrV8tsrBmhRqLwk/RhC7LS1aOdQhh7XsdS+GalSLiPki3f6bUdGVnwgFxsW
XIj27/ZOLIe1aPN/rtmuOAumRI+g47ugh9Z7OtzE8Kdk4YLpwo8QPW3TIwkGV8bS
Vo4vhGBCleuQ1bF287cVtXvENaDTX/a5IgbqUedFuK7N8OP/GesFZJfjVJe50b8J
Oh5pLJXVBRdNnGcwHEAI+zNy+GCfQHVAVYPvW5CF1k6ur9gGJJOCpcsNFiCV4JHR
FYGCRNIyDaE/o5s55viOyHcIGeVNGG+ytcye9mDYF5OxxGh+1dljwtW5cuYxHxhG
7zreqOelEhq7dKm8Cib6ikjo24TbYaW4TiQ7TWdM//WRilFVjEVwXr7C3AnCvJ3E
l9gbJfGkZ4FzGPdZISNlIBA7FHz4gf2P1VDYhqNZC5E82AdiYMhZEmHgl8y6DZCn
YN0MKsBg1cVm87z3CV7my2pZsQFy49ik9i5pwCwXSmy+dVu+KOEAoB6N7Tn1J7fC
g6zia9bnasrKenZ1V6X44gcz51KFULmPH203OL519Fqz+XdDXZhUivFPwgqzgZyK
zv+AqKZSD4jIlWHzKfBEPXe4Kw+/a0FPdXOQNhyL4koEMPn6dalPNk4nKBXpnusn
HikkAllCkO4bkkIMaoNlxVVDccLkPE/t1KoEIWGmn9ckK6+oBQYm9pvLGtm53ko1
kXb1OBtt/kLe7Lxu5QuJlKpI5BC2SPbRERl4Scw8bICBA4kIoVHN3ydAd6aDCklF
r7rMcAEoo1iMt4lrM0vxDesV+DGejOe4u6RYv+17Tum94zRdd++qJIUUEzMThsT6
fYfWnUIoMklyiSKJa+IsaA4IgpnIjlQwDTYlZh7mrLEK9swv4ZToLR+bgC5+ocp7
KGGnVLSRD9iyROXRUd63FwQ7TuJDZ7mKknE5B4l4ikKU4BpMfdlxhfaI9z29AG3p
Hr47oNCFy344vR/oWSSlcZYv4HbYNP0Cagjl+yQnVoKbmSRRsxpVrG0ktUhuk3rG
uvQ1C8JUYVyAAEUSyO6/89/FA3PVPoMtMkvVdVq5pjgtDSsbLY5NGa9LddHOQ3dp
S7a8t6EE8zBbS8leBIUiyGzPbEZ5HJcFf1HWReBwXEbyDCpp/ZCZFtmDBdmeEpha
Ak6vW83YMCR64kwUQeiR7rCAIUYyTAAbqiCEVS7YEZXPjvCBTznuqPOlAEo6U53q
V6PnDU8aFLBBkpoFe9QgCJfxxq7ltz2EPussXf09dcbl5a87oMrszj2LC1TjQ0w4
GFhCbGyRIBP20n0S1ePBXGvzYKADbRaScbFvlE60aFi2yjx7QzZwmZg1/ATblJ2j
L8b16QUWEaYnEFkaKsr2/MCNwMFQ9XYWllyeOT/Bs2MyAfA/6bGqZGiqe521YPeB
FnMD7UvRUqaZS6V03rjY5jrwjtV93aILhuMNRHAIK9QN77bc4B01RJLnGsQ5g2td
J6got55vRFyKwmjY9ycAQm5tT/aIUjxG4oiSjCB5cT7URvmsb/AOtymHyMmdtIJ6
BONwQ/6qzHOixVFWWUF0a3swtoN/OgSvzTFN5B+Txml1mojzKERV+uzDOknbBFGT
NEqtqHom6AXi4bvZOBOCzlbB98gOhMeje5Kq/9v+lY9ExZEfJnIBqWziRfuMVhRT
MflelLjyCHwnC/GuGyITyilei+FtTBNL6lAtsiC0R0QdtP9/qBxYLNG4+sqKgxQg
bqFWm8kBc9xiK44AqwCF7O+/tiqc+ziqTmq8GCg26/CtDVIjGlj8Ob+OElrM6b6f
w5OymV8jTFExc1VAuN9h8hGzCGIn5XhFEazZMSv9j8pIrEmmkV2jTg7BpZAryPiy
Iw4Cjtc5SJY1K5KB9fBycpKjR4ugf52YoKzx9RCeRoVQDadx9PuICgn3AtoceP+0
ud0G6w+xz5rtjhPi1W2xPsoJO3VT9X4fA0Ls5SAm3+N4NlvS23rVBmSdNV9cIqCF
m0T0B/PM/h4UAoUo5f2V63RCEvzU8+gi8IS2QBCxBTM+TCHWD350px5ALl5W32tQ
kIWhrbVrBvhm8Z/VodPen+A3oAhzHVFwEDYYRD9rH+IUxqHpRfeV8uX8nSgEM0da
4Q8ZTArL+GlT1iNWPC20OxJOq2p0vjrmyKfAVAALoN/xE3x+Avi3KEXlqYzzdE9q
QRTV4D55GL2W0vnmLyCkWyVI9szJfoCcKUYghMNbnNWpVThaePgRV39/SrI01hyN
MIxWq3epxA04O8oV8kni4IXrxeQF8CGMzanzhe9DYIOYwr3wpTzt/Ue4DQGFhucr
bdvs1ZM4qU09/z1dy3K9QdyT0DoIsBuk/xgO+4nNwaQClSrHXxJhaBeGOEXQMEFs
HilWq+f50DOYhTqBurAcC/M1wrS+hky43b7CJkYGC7xVQcpuU/wJPAIH7ULKJyNC
1ZwwhV3BsUsY8qh9rEQjU7nr9Cduh1zJs40C1XZjXaM6q9JuRlyb3Sfh5xzde3zE
AVnvP0nnLHTgpMEmirkXbxeWTgtJueoP4IVpolaKahF88WzIR+IVG+9llvXntp4u
D1Wkt09VNaMdUjuyug30SwqOItN6b/XfsM5k/Arj3645ZCl0C433HJYsoFbO7kq7
myX97UO7NtXHTuqZIgriwp0oyfGv8IlsHPcUcZ7qUNlmdbRlxWKgGaaACdofHdoK
3JEoQcPf1/JnOdfvKhSr6IS5JXMTOt9GN7rZVWEO3vKjmE44idZUAKCXIDpGm7TW
Ma0+muifi+blXaTlY9iUC+tkuZw3DHXcf+Svp8SjQ2gDliSSJr4189SkNmU1y7c6
jMmg0UYf3LwsGwi8TxXBDyNDP6/aR1UCNNXC7aCk7fWu/NOO/OhYdTruPouY814S
1Fkyr8dZ0VVRN3I9ILUcuzbg6SoEMJh+rZCcVRrXZQVmoru9EUe7tHSoq2dW/ZV/
YIar5JGyQiZe7YCZFL4SWiLQxB8o2kd9PBo+P/XFpqx8JK9JlRO6fLnXyYS1DYbr
WfZtiKN6HN/c0zuXqneeAOAsVwEVhWxkNqpOIJdk0uTfeskXBvM/lG68YfKYhOpt
gKWlRCOEekpTPttZ7S15ZHOPKR02I8AUUEhR/Prk2dfiQfPjnyd3FMgKorN9didL
X4GrrALerbu0krXK9I/dwSmz1UqaBMDGrACTIQpZGLdksTayCQrQgAO6abAa4OZ6
BZnuO5uxoofVXdoYDx3WfCNL6hDklG/F138v94FP6/Inc6is3mPK8d/LzcHcSQoK
QVHRPm+6W8Ypzs0sK4kYcgg0n4M6ol5GhjNPnnp1Lwxwc5QW+x9tMJ7iFwQijCeN
R0Bo8wHJJBn/5lsftjfm9Hcob47uk6J5CMoXN1N8VKEWrNrndpI6DR81D/DwVQ6w
eYdbaTqRvSnsEkoBELVdti+fxlpDKMq4g0B/bISicCh4XJMoRmZwVnhdg+f2TUDB
i3RGWM5EB6xMfPZBEYHK3Hpx5E3bYA5PZSEZZ0ULj0Z61eQ7JVX/K//oC8Lt1fRR
k0v8uwOMQ6MeBntohsjYiY/QIvpn+gibbh7M12H+Xd71rzaKpYX3NbyscHsol3Xv
yXiQs6EIAkm1DkcnT7MPFg8ZyVqB6iTXBQpdFiwlCwvVVPanEe86WDsm33GKVjGx
vEhh0GPsY6NreC0Xpoc8Gtl/mLE2A2g3UdDxKmJgCC0ZQHsocqe5rJuPQ8O70Iun
mlgOyl9Cne5ykwnx2sWsIBIjtikoV9sDvzA+3kt8qlUFoKYy4b2duMZ+nZofVFIH
ONOBA09lluyrciEOKfrFT8Yn72m6L95I0W9N3Rz9/jhCkkGt5DF5uin+tHWPgzQL
aqZRfCsdruEcoaKye4T0uSIOFucvB6zMEuyN6lgpbXQL8adY4e2UW89LIPks+gbm
j8/ukVjoKZLFHsIjpf3D/AGKgMJZhXMkCEoGhntJZ1u3nQ/OKD43UHPhnpg63bfQ
hExLGpx0NyQp4jGD7VC0JIr01rWp9Xio6gieBaswsI8Lm2zEtxI8DKDrU5LjByxh
7TIaNUkGS4qICa1bwFkYmrwifL69H8zdDHGm2p8cZlACNK4xDMPetRns4F6gRW7d
hK4VSfpPHn1ktLYuSL35pDR7sx8B2Oc7d+mUI1m+SCS1Hi6RfJfNzNROHC8wfkly
ER2RBVWTKsYAr6ZzEOwM7Z3SqvOY1Y6qiGNxPB/xF1Wyh2t6zT4yiA1vtZ5AiKzO
HbwjqMF6RM+JkXMfsjrfX8+6l5dAd8LE047OfsakFvLX5C2QE4S4TWw0jp8TUt3u
h0iNb1x8a/+8c4BOiLyylNgqaDgOZAeYOksuPeSXZdVzQXTohkjUKDM5hCvA3Jmu
PS8wbaHU44GsuuMyRLsBwt1Gblp3EHYcGpKd8IZb0BkFkMTPxFO4WTcaFDnZxlKi
IGTR1Qv2dpesj0HF++HIq+vBCEOX6qkbJnsKH+6ErUvSslpIBbONJyr32eAQRO1f
NUJi14qpGzvQD2mqg8VGTI543oJHHMwGIfsEYcEE9mIMOuXK+g3wareNRADryd3N
VKNhGTmiEO+ygwFgul+4EShXc95LeGb+eV9rAt0v+MBMPPIbRAtBHfsZZQiBRlq8
pTzRpg/jJ7k465ZdDrACoSmjDhFz56ReURvfl5wNL8huxuHWp7Aw4CvAGf33wlgP
4VkFLByb9qKdtQIvscUeCixsXbRlWOSRBqjwVB61dGXxW9SIqLRzqaoll3F3dAjb
VT5+EbA/u4uqifnSZ/B5giun+pbulJOwl4brOKk/+RecSo7ddXhhTuqrdMM7yeyq
RrjASAQYX3SAKbY2tbQxJ+XJn88pkjwMMalFH7CYPKMrao9Fl+wkkqQQAUIqkWg0
ULCnE6fbKhgn1FtZRzmIyfIFRvxEWEbJORFx2BjudZwBpaTjesmbCBHDy8SWGca+
4VrNWnO1cyqXnPCQmZOkVDmRmAnpWb2OdPi8Cby2eJPaw9WH/7+pztumpXPhFfBQ
8k9UP1byVJid3ZTj6ZYabOf079pRq2HYe9GZ0S21l+xbtkZaB2ofwVubWmJ7pA85
bxfUSluCO/wuEbljLpzmMzIorDtsRhpYAfMDzJS8oORrZOCgOII4EsHVFb+eY+UQ
AHj/Q08N6U8ZkgJNa50xQ3e2JAiqgoX3gKMMLBzVwh9qDA4LcV+OCEH5LROzOBVh
eZElsnWq9aZ8aoyZm37zkoIky5iDqBRYjZ/lsD7VxkPJ1hNZSxVoh8/fdNXA6CIK
tkOhSoJsWFjK2knjuEQlrZ8fPV8+E7aY5NBNdeNQ5g/QIgao4JP0+DDRR61QIsoF
nJiFBIZG+nA8v1yYRJMU3Cw7UvcQvimRyJk3sa0mHdknjpFX17PEDASP24ebsyJR
jheCDblc8ZqKfkLpZKDa5PVHitspwvZdm9KDAh8jPCY+0/GuGpANCEJZfBeH1IMV
zjtGKZ5xuEPLPAej4kpekrN8WdFdFvxaH1+OcNuOqro1h/+0risBxAC/Fxs+aelT
EoXRbSQmj33Uew8F1CxBuUaWuV3C0isjfy4heTMEZzghMgD/mTZFcr/Q0J11mNjg
JcVFEIqiuVOE1Wt6ZhhCHPwMmSUV5Zu/bCOt/+uPi0cxtlEQ5M5aMAWxULr7qxYV
Cn2Ly2jTGKqVGYVv62q0rQ01wd33HfZq0q9v6TIP+6d43m/nd+I1cpJORUS11q4q
9HtqnkLc7klPCG4oYqrnfpQdpdWDHLkhUZb6UTLsr8LxSY0mY8XReEvES9t4YShL
fFLA0NVdbrWLNbeI/NSb+5d+2kgHr/0UP8hocNBAQEmbMemp8lWX5gIWAfBe0OSx
+zpPn86WbWR2lx2041L9TbDxoFtAbJtyyNWQo7PjxsXHg1xXniEHkEN0yWD+jb+Q
BjzbUhhH/LhL8OMsdHRdp9xABDib6rCHEZyyNW4TwpumoIM/FGuFVd3a1zL8OyI7
g5BLDke43w+YXck/YW+61Qdj6d1aJJzK2URxbVa8Pl73/MEJvLw5vcD9DjESYLoS
M7i8suWiWDiwSHaE1n4Hhq/BiJuD1dz5Oz4tcUwnMDETdrJJU5DkEehPiaQ9+T6R
/cT5hHty+E+Fv+GH9E6VtHf0OAcRYJVFfk3s+2szBhlNhQog5fl67Qh9jGJf+Ioc
kXUVCduaLMxsrdg55oPmP4rTgEEJ2I0abWZJ0exFrj2mequWm7/auA9nvTINIypJ
3L6WdB7YK3E2sIlzWrVpLa5fTeVYFAeEmBByLIxrvWHPIqJU+gGaMk5Zn6cB46hE
Me6/jIGctN6RXfSED0r7z/D5ZR+Ez6TInKv3qALCtqevJgP6M5ZmkNPCcHfs9LHM
Tgwr8essQAZGFML99BPTi1j5f7tTgwYuMs85lVAR6CNpddLPneo3PvoKtULTIY0G
/092wr66dfMtDq0p0yT32PVaM8pXNolWm0WW106alFOmk89kACznMKReSw9OwL7t
Z/oekhx4mHxxZpiNZlM8J/P2sPEvmTYZck+DCwpturB9j3/39T3GIWL1zbIROnti
mN1zqp2fl8B1RIo2wwWoTblHSk+auTPJeaOtjXTZlii4g7KdDRZq+nZhJGIFOYcx
MxFUXJq+PuLt8ctttaWPD4xZ8+H7IWGPguWO3FyqESM0L+ENGmVYgI0mUj5lnU4H
xkbl5wXDU1Vu56bTkyZD8oM/GMR0r5SaZeD7vdfqoxizuEzm52gaT+IynDuiuIcu
QjKOOUpnFbkO/VNH/qGi8n9XnNyTU4G74O7pr6TnkHhi9pVZzevbte+me0Ocw3h9
nzExDWQgS12Pnwvt8yOGPDxNQWRDNlTVpw7GfltAIopzXMNwkcdcQyK0euLIpZjx
mZvLa6F4qMh+wNaRuOOeYJKzvY7Vyqmcw21amHnhXuiOtHxxOLcdaZibPjq04lI6
r31/6s9qE8K7u6CE6eP4klz1P5fBF+tN92cPXISm0L5aGK92GodkO+v9zFS6USvt
uJJxs0AO/1iLwd4cUfdbCzGeDTKREMY0949rqJnT7Urs/vlyDP2bp4v8gqco4C4J
+xKCvZ2jPkjFeJVGrQ57aQ38BfoPHPCiKaqvAqkK5DkXWF3TaCCguwk2hAwwWibz
Ta2DNOaMrQnLK7V6UguYZCitCinitySh99cq2eTz1BByDZvOilxjsNgel35gqpPM
0X2drJfy1vbHbPynftRXfnnJ9NGDudORXaXm9P90bzV9k6lx68d7BMaXyj8PibvH
6CRAMuINMRjj21rR3YHXSi/tb4tOn4rEjq8zD/AGXhBSYNSUfmP5YeWLOC52B/Wb
06Q6ZJnGxVwpLB90viN1AoXJb90om32yjT+ATCwJVBDuzRwzPfgYiab8WeOBtIVf
yLR7PImBoBNU8zin+N+nnNITu6ddjHpp9/jZB2pdjtINyOeZdDG48dCXpAcI88bt
uVIx3092Ry5svahnBEXCzyOk/NdtEm0BiSiD7+P2mBwTy2T4LzeMa3FJyoUotir1
xKLXXCtgrP+oH19ptfDQy3Ki6RkyV8eyn0HfY4LNQhVNdiCDiV3BlhGWTfhaphJ5
ALoiiF8BMsEsQb0S4mOcSBRO+TTYdTRw6EEmcm3EnqtrEa8Icu/1wg1uIcjRS3PO
rOb/tWYDIkvQBk4VJY0HFsO2pTuCHzQUJ2PTXGdFkUu2SC3sAbyZG6YSE7x8i0kM
7zytWe9fldsxWSKPOd9mfaCoy+4Xvvs5cEu1qk5VdrUWace/1FxIbXx1LzUkfIEE
5m2B+Jlaq6N8YwuN5ws9JWbEYQpyloELN3/5Y8XlafvnfN3vNUuH5zrvhWDVEc5/
Xa+DgGINdcCjRPymcGdCXiFcfFLYZl+JQc8eFqKjyY3TVjpWEBegZGLzgaQ1Allt
w44KsBWqJwoMxEIk3cK9+14As1vqRfjaETLlknqOh6fPaGSYhoE6tm+/P6jgWJD/
cHBzU/pFxkXZmspabHSefjAvN818s/jKJ8wbAJCOWYhqQCDGUJz5ttQykmcEIcbm
4ZDG5+pqnbuvBdYRPVz2xdSIS9xzakhpT/r/ijhdDkfkD2aFjmo2efBXhVkQ47W+
KkftdeSikOOHg89ZxcxMXp0ZagaV0J9Ypoumgq8JKJZOXf0rmh/ob8oPvXraJPOe
o1pK7jW7IKet2VFgPMXrbRDK9ForPrizCh8q4D9WWWAVWfzDJAFW7vREpN1avbRo
vE82Odes3EBmVk6HMx1mnHbbIjFq9Kdp5NuEokKpLcKgo2LNUOSf8229YnTgTbwD
d5XqiVJoZlzdpAR6iPxIYqQMlHZ1NqHt1frI+fNMAQcrXxnMWM4O04IOiU5JvMjj
7/UHh0MoTCeNKTA7KCzxLt1PuUUGF+ISbF4N8OrLkB4TdpU/SISYEdh5LT9hLpjK
CarFC8dHhD69UcE4sqksViIOnGGbDs+0OVxA7fBi3wy2EMX1/fduqaWVv+YjJZUo
QXnUR9AZKAdIX+nS2x2g8kY0jKeX+S8Z1RVlqF7SwD5EFdwZx4kMQedu6Cf1BxvP
MScfTDYSeSYFP1KwGypk07BVdOcpvIBtVxvkNNHKfbVgvL5Lqk+/NH0tAxHVrkaS
7iSyJRxKynI3POkkEVuZbhK8AWqUC+MwdGN5xNHYWEXhGbVrOExBmmC6joAaxP4D
euZFgWxSBGXHJocVTeFG7TJ0dCnB0rX+ebmjW2AirifneNQd48Y0wb3yKHrBGHPL
+tSK57TQvkMyqAxfIrkTR2Q31ySO2ZUBWARcuQo306NQcjuE0L1VQ/xmOePANif6
iqfiY0yozTiVKWMTEWd3JpMJIMB+8TTgokJAFPuTO5DUK/n14rkN7T7v8dizf3s4
ASDjCyL5Sv3ASCVukKJWn2aOuRF5KtmFgA3O/tr+EnaHa821LohJFsskcbEGn78G
8K7QB3UsS/Ps/RmFD1QcXzfqM0M7QNfHt0BOLqYRjIneo5rGDCOB8IV5ZA/lxV8X
M+VJlNrpDAbSI39VxkUoKNX/Xc29tFLvqhCEGnbsztRs3UMBnf71dX0OMnNqiLQ+
OqnSAV1WuzdfHKKBq72RSWCHKkY7DqO4Y3MRKDHLGsg4ZZKnL3JeAYo8D2XZ2bFR
PY0xwLTJDU6q4FJAtyx7vPDh4jSw95anVezd6/XWlu6ittPrPlh5anPxnv0Wh0oh
BUh34OVr+o6Ey5BdBA+4Z0ivgsEgVI+8MitbY59Xo/pyfPuWRL92z/pdiOs70A8I
VsABXBF0igwrieIF3WJvwkdh0Ostcg3KRtyJim+FyVYJTi5WNRJI0iAPPDasngMn
faefY5u8JJm06ETE8YcHBq9zM7UvxK3o+av6pC02E4aEIB06/xpo6ZUPi/1+jfUL
RwqnJbxrUgKcJH2Br2skyLKRz0GT11Kp5kfNOkGsfFRcWFVwB8uR+ZQ5mbivayX8
sTh7MlYuBy1yZTGfPg3iSwQpnDcNBMFi3NcjzHjK9cfKjlpetW2YnsW7sEjX93En
IhlC+YK0mBE6IHAzg3BcO4Gz+q7NWu1f6qVCpJQDIt80lsEli8BPl9YpqpUlDj8/
IbU8L0dPYQW4IkHbMzrnLN+EmKMqnbKPF9O5Z172DPgzNDjjF6PiQprGTVY2XIQR
OMMQmK0hIL5yLa05IvWr27h2TbVfmZYf/jCfiwf3FoR8OyxuK84ivDswQ7bPtKzg
U1QaouhTp0w+FPuge05lwLXTWyaldowRTFzrJyi3m/VeK+hWwZOeZiEt3d8tSlbp
MhvqfMBrT/EJmb1kt8hBwSCohdMtsRFUHWSkFSgcNeQZaF7Zsxows7n8wFdDaNiV
4Vm2Ohp3M/bZbYqBnoE+j3fpSmk69fkDhrOliRPqc0ZMelEhnEUW47qflbDnDTSb
BOUats+0tmtZeV8fc8ndWmw3vvL+kIqawaeqo4A2UFsPxluFWNwJWZRRtqIlcWxA
HW0uqHg4P7sqRI2Zk1PyGYLiUm4SEW44NHUgNNuLtPftklM/AYXb2JVBaZXzQz6k
y/TaiQJFHB7reJbfUEEX/kjeITLV/e82gY8VVSXDsCYrlHSj8+ACR6duKoM4/tmZ
sNQ1q0pDcEaxUv0WD46XH0Q42mGYt2gAXkQ1EszSu1/kQUBmcVz2sPmeY/mac2kb
D8+gcIBH5xO/RPZd/Vx9FRmld22U+C7d2z9lRc3LUQ+eZo9uw1Et6rorbt2UDPg9
efd6/iGX6DVaIak1Ds7Z08ttaWVwK4Y22QL2Z1m/Nrf6so17+MO3U1P4DItt1NU/
tmiWQP4FTQ0XIIT4umQVZl+KWOht47olTAXdWraVOR36RStyEbAchTQThdn1lhqa
3MbG+qVmXlFtVeMt+zwvGcTRP9MfExQzk9KkoHtcedMiFxqPXqt5bWBBWI32chsP
XAofSHcTwJodLtG4J1eGTPsLVEP377Uc4w54lqMZZRs46cH4ppLsE105BMAfrj4K
oaR8tp+oH4IyPz5w+roTnKs0zGv/5s0n9k9j7cAhxe+8oVVFZObWQDJ3KI0KXeKi
Qp/75Wb7o18ikiT0ESuviDXJZ+QC95DDFD8FL92zea8rGNwHDUmjBdgq4ooXII/V
6V03NJlzMFuwoNAh5tI7eBEUtLBJygK9+3DuWVPamo5mK35r2qNYUQwdJJgqHTDo
P1yWZwlK4kzrmN4gg8stsLxKlow2agXWSrVqCjevRnkmW+JCqWxG8h1NqN04JruP
HHafpq22gUnfpaVRzG0Ykye/dkuzkYQTmfk0VMW0fFORv1dqbhEuObshoZM7k+Ve
r3qP0gd/vyyrMH5/SwNZDmKuKiXKIviopngW5NfFhGjkM6rnazoHy4p4LowvxLIM
CebkfeJLkzeEz26bRtXtq4opwjQsJoATyc+CTDq8woQHe2MFy+221d37KcwXkQUh
rLXHJn5PeqAyr9nhvttpaS8CBdFndM3NEHfwKwiSruwDkOxaalrLGEyBIknVZAft
jk+QNt93u226lB3MsUgdqWcv4tmCbP132Pues5zz3Det/H7AfYqkut8ubIVMyth/
5+QZ4PHYAVXF/9wfv4BT6FvCtjRPIIHNupsAm7VEueyeZkqiLyBYb80/5Cy2WL+G
WI/EVwzoswaryXmQpTv3KjqnbYqCGx7paOAAJ9Ek2Qkb3Snhszgus/sevl35YV2D
OtL/42PPky/PIUqVCuSOkWRM5EXbkwIoMrF/EIsfwlK+PfcbznqkqJ3O6LfZj5RV
/PeBZq6Fuamng18+C9PBnYbYmkf3n+KAh4dmxJ7RllM5bTnck8ffq13tTrhfvgh/
eV2xcozxcCgiejgakxpUn69r1VuordYGh0B+42dQG2VkZm1GQGbsWN16RXdDLEUL
WgW3YZ1+A14wGwiuUv/FLSRMoftaURof9lCQGO7SAmQB4fmb+VXVfaZBfH7bFLgZ
JIpFmom3cgdUcsMx9TjCS132r9c0ryBfByigB1vZgpUnH/w6WuwaW8DdKE2Urffm
FI21h6g1aHh6+cb25N++iagO4h/yuPNia5Wfms/0Bzg7MeoEQ8dbdFOa0Wlf7AuK
J5iI3YvJfffLZxZ0bc8fs3fI3T2crEQ9DRq6PLIjaSoIdmd1N8hP1GI3zPfSfJcn
wlzR4hYQZrp5XyJ53S2mPjDSjODkC9ZWRMMtKTnTJGEHcWYlA2YJSkzaNfNPzKd/
e9Lh4Dxva8iGAho022HUWmRVj/zJKco3zrmdYEfMNpM0MtLaBPYiI4bVMpcZ2h3e
UhU3L+Vfz18lA3VucGJL47Julnree9mIbyCW8ems+v5DLIL69YSo1O2fXl5tXmJb
RiUT+9cCmIefsNMAFsom/TgxQsj5oRPG7pqT4fskpR2ouHV1VgtTf3Yo9UOuSsnF
i6HSIQRE+p7pA9o3/YaEy0eRhhkpDh8jtp50AX4UsW941wIR1rdc1U0SPYPAzxRW
kaQxJosVeWFw+D5aamKJh659wovouuMpLeDXzQevblbYBiUV0gmlxLRchJdQsQHB
3WdjGTI0sShvEqGtqlxruexPMVd0kXeHhxYP07VX53D2K3Ob8I6QpWdcL0QZnGCV
fbmk/UMyowVP9kuxjs0800GLRMxOVE0drS0cCw54SSzByR+49peWo3u6TRpSs+g3
i2lJRt79SeS5qnkM2Ik4HxJd8IrMfg3l0gDd+OQ9FcV8+ntKoI/vrfjM0LF3OaJc
518rbZ10JI8VFsQoXgsDrEYn9cTZ1MFAeWk3GHYjrqOOjaG+UM9Y/wh/Jjry3hxZ
bvdRZ2uQ7K0rdwn7y13G050Tp/VSejg61/nw0SabJCR4wA8mCx3rWNN56MfRdBas
MZY2s/FXEe4+rrPaqGYznClHymXUeP78ep1nNRJCP7TIUyKJ1aIfy/69Zphpvqn5
4amOLvNB707D9tmIL/gc/VadMj7rpKF0HJ97HiopAv+TBhj+L7Id/5lMrkQU0FUh
b+PezfSmtwnaD0Kh2ZDB7I7N3t1o4eagfTAN4MVkV/1CYdooMKPwerVOMhU6yvGN
n6O3VPesRQnshCV4zixuxj3/g2reVF51lHlYLJoOvnplWYCX2mG1qN4ayUbzaB/L
tsQrwzvM4A70jGqavlZi5H0On3d8eqqk6qO1Dz3ytmuJQtcYbRfPHWKPNBT9jz59
dxjfWePAyqXpD4wAASAqL8Oz/Otu/71pIvaVzz31mqbfCwExlp/ZvT7xa/d99sO9
kUqbZqz9eA+zBG6QxbweecxS1Hh9nq6ZW8J/B9MvT6NJUTC/iZul/NAPTMW0jwUt
Mj4FiuCIhBnL3mN6ItJ2cuaCULHwSS4SFmyuN8uIClcwEDatfKgTqxFCAUj+LMq0
uaNAE6LPT20v+QGNqqK6fsH1nZxbl9dpXQoBN3daVTq8jQ7+SaMl/0Dle6hftUmE
CILW+hLhB6P4QueoasKBOeDH/HkuvMWLh59EK4LaXNfkF37zfz5/oyy5QizSNvUi
P9rgvaE7FdLjslUxZ1qdR0xqhgqiy3PHiiYRnmfU5DXYLUdWomLYCRlvBz4k/OWF
kKO/v2GfiYITDGZaOzyEgE+7r0VSAWe0XW1idz+MdLc1HpoTUeXA+VcHiHi/rCxz
YcsSPKncPOlIjiBE+BPsVHzcOBL5qJ9JP6sNXcbysY4k+cvfN2SGPfg8GRYH/klY
MTX5N4NPuy+eXpEzdFNxPVf20uzTxqhUFpAGNZuNfwHr+se6vIVPrhtH7FAPIWTY
M0ZALO7kdp8G71EDjm3SWTnWLZxjj/VaxkPGAYDa6hVbGxFV9zIvVBExSxSShUYP
5Oswsd0VdNXDvA9cGWIjpY7aPrrBydwhB4gRQ8GtBPBn/jqpmqRuQSQvVZlmbilU
7UsO1nlcTYzwA3W4fdEENx5dmer0ARaZpKaDCJAb17qYnCeOt8Hkxz8QHTnEBgHH
bQgS0gElCZarOROa6wjK0aAbfhsmTa9xQyfR9u9sLbFNbmNcjId3+pFWFRHYa4O8
++mYbmXxOnKp4fugrFFVAfYiOtuVDKyvBe1GHG+pKjCwuiOHZop3wXgBH10gv+02
lI8lOBzwhFNUa5qKk0HVM6U6Y5jWal7RJaHOgVYwLpwREbhVi+JHYVSTiWleOM9s
hyY2aZQWNXabLRtOQ9mXIdl2DWSnucj6S7ACwNUPDoZJaNu75JBZMlUfHMf71g8e
NErE/5KoeAUK+O/yEELurlagvDJAnyQ5lVCaXIsABXWWHmeLDC9NO6Y/8Ya9qlCm
5zi3ZT0kig4/Cl74OtJu9tR5lxq3M93i+IDa25jkx/VwACzDdZTtCU9JQgogbSTp
plWXwPQ7NBp6xeqp4YDr5jkeJmwzfRH9svA+YNr2EGLww+d+B2ef1gYfV1h6kotv
sBgG3EQs2EIQwdDCa82DkX4w6XHYNJsgnoybafJ7MPbSJ2G21bL06NGH2Idy33pJ
C2i+gYnwk2bc0NCVeuCrXf/sOzzebOEEC4ESo3GPtGizUGsu6Pul9zw4RUbtpUQ/
krMWUaKbxucSuVve6dhghvUJvNHFBa3PU3GTIqgy1Lxn98q5aAPIoMfkFR+l/QyD
ol+RweO//EN9P80bVimy22AUUDpH+e/XeZcfNpPHzBoS/nSG5uObHapNgLKElPyP
66hYFHVnxvm8XD4MpHX/PapHIIKP4OKngro/G9QAcCrcakbC8w0XmlY9NVm0J5pK
Pu96N18Vi07mmQbDq2iwyHXTC+/9FdlqR7tzxOdn3DaL79VsEnEG7Q0T9K65WaTR
myZY+7Y2kEGcbtUZz/iEfUOf8hoAhgeKZ23JIPSE4sxITjqKszgjcEdKZVSIQOU7
Wgy6JjrCweqWUYjKnNwMgZBC+/NZG/LglAkH2mEApmBgLQLpvDul6Pn71Ooa7IM8
zWWYsw+oTx4O/gVNA+6G2B/2KB770RdfdZhuKRyv4Jc5+UG89Y5AkcC7dzaJZNRL
RA6dg5U1UflHdI59J/4hn8RVQJ2YxGBvXSCfDdmtUwtlgoFqA8P+6p0E+JdpOPkL
qz8xUXlVzwrXTT3Fk+ZhtJ6BR5zIpsuI1WJKRjDNjWMzfLYOa8YlZoGOmLGIVQoc
6eSnZIvr9L7Fp56Awvu/G9LHOUxgg+Cah4rlTdlBhqYjvDC9BkwlQMPMmWiDbucn
aHHlejiwOP+9ECni4CaXIZ+rnOKbkZKlh415OKlrOJ2WZv/r3sfqxY1tZUR3diBb
U4J1GWh9vrMr7GmuSXHgp/chS/OBAom7VALPidSXfq3H4lBt4Uzd4GMhDcqsuWhu
pcVNDjDp5SSn9nwjQ6y2fSOrO2aS9IzhWNrZJE/GoEwLu34KKy4erWVqbfKZGL7u
MOJXTZbptSjX3ahjlxw2ezX0XqXNu2T8FRHLCbts+DBAHehDxxV+jfhLQxErF4WT
JP1UBKPlRPRRw5qPt43duv3nQdchvxRN/XZFuKTo4z6FpmAl3g9wIj7kcL6aIogk
PLpX1TUqch/UMZu39JPrBZF/2gXrVRkCtmtv+IMDHXAXnFGUJsQzV93bX0wYMYn7
Xf2/Vlqb4+CAwRrgd5rrXtkSeStZKdqYYLEHIlCCCayDjDzRr8W2LZEwOK2T0ugi
UBXARydI2qt5RgLH1/PHEMOqQVIlindyORbdOpihCfE8eVuIkLqjHXVf56JCEqc+
Ly3hJHebIUpWvaofg5yR+y1z+y+UI7o12pBwZvneYbdSJ8TaJd0U3zs2b71Wl+T9
C3x4J2AJMpP5QCDTD2oPXcc2uWrZ2MoAKpWdSVGNIaa41/OlbUKJYw5g0XJxINOZ
fUl0INb41AzbCE8loCFxyLM6jZ7gr2srvHx3wP+BaUMWzax7JbzBjPNOChERTiu2
ZLjd0wM2j1sABKZqlJ2Ok1bF8D5VjM0ssGG5Mg4nv3mZ0RvtROovy5zextjQ8ZMT
+ZWx3OeC15jd7cKHXpXqzq78xJd9ek4HQBZA+3MgSV0sVif3GYZKV9K2gyeATUJL
PxQQWkzaa3RVTkGte7Kcqwyeq+4LTdgfnPYMTExVXihqw19KmyWlowjejbEx050L
7OFdAGzfS6HpRx+OAkXaJHkcsEqohW2pHotYfbyBu+6fRFkRlwQ4YWZLNxQmrGva
F9GsT8QiJUX3xRHhhrSB3veysJD5aXAIfFqF2Aw1AFworuGAg1vmaZZ2bG19HCVo
IMOVXKzbwzu68vdVAycuwSSDZADPNE4/tJ9LfqX9SdbrpzOgOUGP+iSsR5D4Rk19
kNuGvnf6/Ki1bYg1Mr+7W08PR5ansDnmsXAjaIyoyVlQCNy6EXz5+/YYRdmUDYb7
0X5LKAmLCTrgOYvcWFU73XhVFA6dspMJJPvGxMu4aOH8fEhg/nKM9npnQkDdcq/z
SYNm8YuaFbpwxPG8lTmSIUz+D43c7oxHVg2A/628F3H7b7NaJSRhA20IvZnFAxKZ
Y3Sla1Tqs1bHsqIYGwRl7gb2OjaZ+tey71hKDAMMp85GfathHhos+uKwLlei++f1
eU1QfdSSgVEojRf2Qs+lbYN7IqiYSULZAouSgqh+uRk7V/LUnd2umkXipUm0HAq4
wv8rehuI5gUOSYniZ+DzfLWmr+UuFPvktbESpYryP5AbzAnnxt3Rzqa2sW2hwylS
+KVurPuC7fNPGTM2eGFuWKqMGec5eZ5QV7CSsCBp9AufFMcW3ZENhSh6lcHy0l/r
empwhl4d7YaXx3P8vD719U/u3UKeHg9HAt5DhWIUAPvSa3XK+mw2gWCdkWDWqoXc
45YSzP0cRMKX8FJlpAiQnG83jONWwMN89Ex3gJl3uOgr7ctrTc8WymLiYzVxD8Hm
N/bCn75BJ+hm8FNauts+R9I5cJ8DGadyZblddpLVSMjfDcJjKtBYpm1B1m8mE2nk
+mx32zXCzoGlacwSg3mvY/iNdgtaycMul4NBee+JtVUi+YLGVLHorcklZwqIKljU
KHEpMmqdQHso5Ms2yFOmitDWFcB1mOpx/Dhgjm85KfoCPE3mj8DdRthlXdPPzCVC
wyZXCqnyh3PP7PGhjKUVOk5WlbVSViRtltnzWPRwTyWEM7ruIFlM+GQ0+JzoEVWN
WtP73n7TFVGStPdYuHN3QEhgwDSnuGL3QRbWvZag3MfjFlLLRqlm2jVdPt3x9J/3
m9+5beJKFMpe8eI0R7wRoHWg9glXiOLiNSp6LRoTgL1hVVLWHWZpsWLCmSH0eD3h
CvfhzgLP8pVegXAJFdK0un0LKbLslbVMOk3jWz87/CAch5om2UGhnJJth9CJZU6f
QlTT3SuQf5FL2uMSdC4FrNJ8Nh8Id0KSgFxqK6ebK/0Iciw4BE6y5F17WfQ0+jGm
75LlvzAB0FNR9njwmX/LffygDzGRiPByQsXlK1K+GOtCaZk+QxZLtiDhlUrqQZVJ
IYXKvfM0XipDkx/tmT5Ii/phKNiy5cejUEUYbzRIa/bZvbRvwBI0dSsBeG4jbwzL
0tiTfuV1a8CsmhGRBlbQo9iNXyv3jLFjV/iVMQoTa+aYyOOUD+PJocB1+ZFHXWQT
b0HAKmOYcZmrOYyWJp4yDNCynvUZQDCFo7VrQpLk0vah+nLx7wsmMu/dsjmou+1f
P4J0I5MX4jc/XzIThOKtRZo6c+kRRglkGneqYvc3tpLcQ+fpDoJOGDvccH6leIJ4
Oz0QjoPZyCEZ5D+2c/71vJ2wWnrXx463gcTWg8yOOmbEbdXlQxIrqktmYu9iJbwX
yv1do/BfwRsP1PcXkLG2Wydu9Gx+vwPQrKMHiOCcuTbcjJe1A0ZKF95uNJReYnT/
XeWRcArmRf2GH5O4jseljynlGB7mtmg/UUYWpQlCE9YjQxx6fdNErclCTs2fJkxS
m5Ic/tRyF3CiqdN8ftXCHeYDsGcWDxMrcKhK7YSaRPzWq44+3AfN3h2vNo8+1kAR
/NsUzsa0gMLk9pnYDREk4K4yWKcPLXUgxovMtli3Z7TLrzCahhoOYgfEuz3AJhZy
EOkQVgX+l0PUhnohGtswaFioBEUcsYGsQ2t8Mw0HaNJgY4rf2OmMVnVjEHxQ96Oz
+GvEVHMlOCNjnUst1p3WpEujLCWRzt8u3OKB6t/LOBa4uhYAicWd7RUpcLALt4WT
yhWsqvbbFbNpdW+HCjXNwviHwMwgJ7fmp+qs48mSrgWsQqbggjRUUC04LkH41he4
YQVaC+2rS+WWuDNg0Vt7O8MTLq6k0SLM27+VrC6O0UqdIsSIFuv+SiKR0u9moSG5
YkfYCGB/ynVzgmkmJHGNMegVf+jbgJKVjpwGECiHHG5N5VcpYMs9gEaNut35I5Ey
Dm/MzThssbp2PsA0CjHeTCHzqrr0ub893Qkwuxv0MbrCRjTqoSOh4ty7CFJaNHU2
m1DpuVutG/yAF4MWSC4Eg0RXwVCczwWorfjCKZ4J+eBzTGRw4aYKUeKZ3s5NA/g+
yL5boAArXwzhv51OcfRDW8YQYpFFPgo2DUIq+ZNJLhtstR8uHZTUEejrcBQI/ERg
+YHFZr+B8KjQw4rFUPaEvWtPrvpP94xmaemhwfUS5tjqNdawWnst0EnXjf6MI1bh
zIDNh4rUL5lqpffn7EhjjA5E3+/l3K5GZ010VJcrn2TScD3LS1hjqQnLVaT57dNK
HHwWZQFnQGUqfkB8W0lFawpz8w6WnCOXddqn4oqcLahlzohFXJEm1hl1CJipXMuz
IpiEorDmLbCzCXA09aL7wp66W1nqiTXbc819dH4Ndk7m8ER6mjMB4ZpugwXTa+FJ
Di9CLT6sYl4aFS1mKUTjvCNky3eRuHu9ryXnzXGifMB6HTeJ1uk2ucdR0RW9I1v/
C8ftTAzerWuL78z70DewDg1drEiUqu7LRVPrc3uK5cT42Y8PfvYlB2ZK6qygbN1K
4CBfC2lxQQjmJ9mbbojmoMUSgfJVo/k5Wf+Ko0519T9mmqy3+9dqUhdEIKvDtf0h
RE2MarOTzrqcMsO3IbhKoshvKSmvXp5mlG3Up+Z6/8r/37qI3GokiV9rG5o6869e
cU9MC8bLD3t88a5izxDtCsUcrZ5b3I9/uApmUqh/+1SXVSKeMCKn0G2q51k/Asmw
QfwLzOdEtHOruXc9xTTvIzd6sAo/jQfY41CH92hTWRHBt1Nlk2CikUFR4xBprnLg
k+lslULpfT46e7MwBgh12/Cxf8Y+hyodoqP7k9thGpIBSYKDsxCEyObptSwGrrLj
6aSFnQdfxfQhFbrFiTeJHWkUvo/G4iZMTCaqhetszxH6XYMkhVXoLKWsEbXYdSBH
z4p2Gn/Yghp4WUOQFfjGt7zMJoauUDziVJTIuYfqKiwLbb2FYwsSRNxNL8b/iJms
enBNHIr+uNvwAUg6nJrnRw9Pobymc7/V3AXAoFHU9HyIxLwibk+fa+wVxdPk1yZq
xgLaG2nVGUfhjQo25zo3AlChO8FYTbfYQZiaYQh5ItycPwdvgrTIoAME2W5Hr8In
ch9t/xbm2IGzzSKcpv5mgewzhcKcTT3QQZGANyLo+C82CwfCYaRdx9tbWA+oY8Yy
LDOrABmv6g90pt2FwskJxD1xz5tg5SV44o4cR7nVBx0jbWftWsISQQbCqCV1pEdD
mT0N5vG3sByQv/wkIN8h4iFSR76s+s/CQxG+otrtiuVx3Xlq76t4WPXUiGkeVb/i
jcrkuuoM10k2HuS+dK0IKvUB55RK2D5fe95pvJ45hFGSXknq2z8iAsx+m+1l7eew
EyzkFhHN9rZWZrXmAa53+iSFAfpydCjRjAAtBYwKCSPpF55nTBxaYjg+/zGG7uzB
VYBs7n+iSqrBGTqv7Adj20GLWFtsDOF9gRaRnhYEJePeeN5AgiprpDcxtMIK5yWI
0pjNQ9LirR4SjLktgwA9wnyIT5DuOvJLuXGnh/HoUH/WIsRsByvPaVq63W5OR0kb
meA85zbJ3yWryAARhNCKBr4WoeEEgPwuyoo63AbmhYCUgb20sh99Ug5M241p69eV
4ajPfx1g/aJZyM36Psoe10eZGLulJKHW//fOSsCeOseGY4S7KK/btgeS8gnYoSnP
S4g5CA6k37x4X9Q4ALnwvXUHpcE4I2lIeNSe456dRpOV5OJEWn1mq6vz96feAYTF
o2fS5Jsr2LaYnJDX1jo8uOadAIBHkR5xdLnjOhvIB4Ztn9zbLxxOEMwZGNtAunxy
pM30GSc69+53qP2dVZ0O+8sK8YTdFkAnD1Gv12YEFbn1qpwVd1pbS4xvmyQMSMek
iwhB/9Lwv54TBpsVD3NeIdmWMNtAkM2pn6szBB9LS5B1zxvJBezW9Q3X6uhfXIe8
GbRhHa5/+jrpyA0txoKo8z5ymQSPk6HVTuMbsPggFdLXCNP1wCzeTxvEpMJf8YuW
x3zIOCnw1aYdqtwt/GJZTw/jlpjrlZpnlFdzU+FlBaiwRMirXw5KHF0bt1xPn6Vv
C7nxvFkZzu5KaMhE8fTUx/z/KOHukfKF+pDvuJBaOuOkcOzW2PwM1HYBgwWoi6+s
UOFHXz8qCtYG3K2YYdvw4xp/lM0mCZEo/emOTYsMR2UsXS81Wf9DG+3zSFt9QByf
XhJDDPj2Gyob6CmA/rHHxOfBQQ2dvf8MzCpI8GHjI5A84n5bQ1ownSWCoq0/xjQD
h+uDo4hKGIgJ8lImU06ByNRTt6pMXB/hq+lJGgYsm6PVTSB3IG2Tt/XHdWUVX7Gd
FNqN7rz2renEmjJ5BYUGOyth/H26HW944BmxE5caEW+2EclhLFEHehk8jnU8D0vS
WrtQfkurZ46NocYzvjwA76FuKMSw0z2TgtQ+0zlAlt1KPYbICdNsOicLZlaeCZWb
O9hC+uQsA3WpOqC2Zmy7YuIZzIzY/Azw6uOKaHYoMGhlGZPptqY27dcDbNFB0IIY
h0r50brtnzak0v+8E4gEUvgC0y79RR1zGrKCVW7gZQRrx9f5pZ8cmxI1HHM4L/wO
OMxnyINZMw9Lx9gJ4xQ1m+APud/zjTESD9xPRoln0rZlj0A+PtfeyiSD134fr+E/
rP+gP1EbcrT01eNa7D0eOCJGDkaesf8DEGV15DVa13B+GCZBdaC4AbXZqGA+KRb/
6lqOCaNK0enBA5mqjBI8ZuruduhOKBXNYY6MxFNyiuLd9LMLlY1ErhJ5HGHinWVr
VFYZtvTFu95Co1z7wqNVzwSO+XEQhIoYxPyImoyg4iX5GZZrbeVYDeCDd50OPQCa
fGUe7AUuHQhz73aNplDc+jS++FYVj18kLG5bEC5vLHtKd0Cl/j/jASgAEAZXKp+4
9L/0NFXJ9xNiKz1iG0XskXTzXks47iulztwQK7Ze+IUSdJHxO/S8C6mLlg9LmZzU
ecfHzWxAUCn3wYNzU6qWiLb/EJCAebXtwIMvyadFem4cwLGqPBFsbHMOBNkCp59Q
fjbEjZyHIMHeUyfd8i73+Pb1EDVMuJTTRHC1ybI0+3T2q5iN5n/oUiwEwT4pXuPF
spL4620gIzWAfKAfwbYPk7RtTKQlIG9wm1/txAAp5M8kAd1W0Vn7jEF4KFX6rW3D
7lxsvK5k81wwOoJkiAXdjcNbxiytoXXbXG2bOPHUpddIBJP8+AdfEiWxouuzyvXU
lBH/7Sub1efjkfylUPygmuKE29xi+5prsEPGAmSYnPocbYhLZO9hFxCbY8Xt0tmI
fU8RoU8eN7xnIeExSi67qJ3sozr8HocCDinQXXPcPwjDg8bdPfMsMBdlpu3PsXxB
nwfxF9rxnfzeC1sKNqZoD/5TQhFb0LnJC0CAg1kM2hdFE62lSr8gks+QcDJHjKPy
fpCvDqYmohYxl5/uBxx5D6QYi/7+xMD5DghlBaOMj86VOMhoMN3BohW/cJpQ9N2+
bL1WVBnUnIflxAaLQwio7/GjgrsUdqvpxXztNxA2kgTc5kzGtrQj/Srr0LBdVsuY
DT1OCVIYrlrDid4K4l5NlAx0pCMn+Y7FxBCQgbUi7R7DGlZ0oaDOoIxPCAmcOHf8
X6RI8C0auiAUBNEC4/ReM9xU9mhDFUD7udysR1b3GgIKMW14UBsGocvr483XCKac
oiW0x2Vz5l7By8d8nOhiYu5fpn4H25nDSYkyc39pwVcC4n2k5rCw/YyYN0yqctVj
d/J95q1Ia8/xrbyN0b5F8y5bJn9oUR0pz3ujRNYY0RjAcja7/YsZh9bKQYGvPqx4
8+YggR7fYuSjpoZHdE5glL8H2oFNX9iVIn/IREDH005SanrT+i3NgvHRouxWgSK6
a3Mvm86z4Woa+3rbox2IyKfoz654RzlDT/Wp9fKt42YfGPHPEIy1uz0EcUjiKXry
enEFEyJUGihWfYVfQ0I9icELvaSZqBIxTX01aG92IggXvRuA/VqvfkLCLaJn99bz
ZX1ZV/sWY+5dPEvncEwG2aEyimDBaOCZMsd7I1op8/4e4bdrFzG4IyP59fupw9fx
3qS2nMpHAaZaNliEfDAN50IEex3TrSDcrvEk/UGeNlGLRMgtvkf4tipKOFtgeAn7
3OYtth3vmAqJUhQuFRD6du+99B4MA/78g8gpUFtoOFlSZiO7kttxNBCZ6Jwjj1mr
ybYePV+nR1K7RunZbau9V0MDSaLLUye5DRynZTg/i0LkA+x84SlMQShdq1FbCD0Q
KSxtXiJu50/SL+vH+fQ7BixbOO/K6laQxWO4001ocz3ypDGy+seD961tGt2eHjz4
g5iiUt/mr2vZ19ohJ77WTvJN5jyPWcQflK0NV9rjj+vl/z759glRf9pDCT1Y0RHS
3NzpRKU1g/nCooaUf9ZSx4JkYtfty11oLoO73lHJ4yw37wJ1EizcVAGuuiINplOp
i0u8GONsFTBcBWatuWxun//mDuZyzbYsIxfYLwYzjudhb0327lijmlvWDpIKFLZk
QwEP0YIDqIoFcttavQBQNq1aSlDqUpWavd6aGOu0Ux3eS27XuMmIdToDSJFMjbki
WIZMmUWOLc06zDqx7RAbIXLZSo6J9EU13HeywoJYbjB+BA/ggv5jx1ivuUVos6sg
mOSFPLAeNL0YDCEGLKMyKr+3Dn3EdW7ozKQIUjM39TKaZvM3oIOlQ2kzZcOBz2e1
cHqKPECC8b+Z25JFqHii6X74dzrTqtq55N1vCwUSLUFOrwjIfBHVHTYaVizuo60h
EQ0KANBma3Pd0xvzUFb7kn8WEmhuuWPAEE/24tQ9A2ifEulZJV45m7zZFhaE/q1R
dP0T3p6cG9db48l6oUoXpJMHw1u1+z2E7zNv09iBKZPzzX/TXymXofTyDLt5HUlE
/5aKLAeoKUBv8Uf1qrFt2Ct/J4IjG2ODlkMsY2IQdRgA1PyxfTocIvLQRN3RHZwA
S5K/0IhFCEUfa2kW4dNy15mi8hcdiaIFE6u3RSf9bsb/TAde2QCYnsHN844EgalB
62v/tk+aq2+tb4aZCekxr7MmRMxjmC0NBUkR5dARsrEdyF13M40GHPcI0jWcnSzL
1mALIIrya973qo+LosJXTh1HR6VMj0aewtp0OOE+GueS5GDkJ2z/IVJREdOrJRrX
0kykZEiVxWQ6g99bRWtn5cQ2N+3nIWuWqprilwH4FuY3P3kh8wVgogLiBk8UxbpA
8QbUeMRHKW/tiQTAH0nioIXszyPgu1ydLrEyQEyaSvXzIDd7+02nkbm0LSswo781
sKa+GmHBFDyx3jjdNCCp6D2LgY5i7nqlIeXPr8y29Hkh3MxVsWPgL20R2ZhEUu8t
O74GZ3nuJyYeejFJMxb23ZBud/oHseDJs8Hn4aOf/yJLsIopaDkc9MsBqzyWf0eY
u+MAyEfSDnRA6KHJpKWaR2zW7IKsc4y6mv8kJ5PCqOyYnzQKFMoefKzYoV20eBsC
fbZqOm4B2CrotvklNIP+fTSu1FrTSH4Tk9+b9azfd0YwWdu52cU21N1KeylPrvr+
EOcdbOf4ZNCSnEx3vveSqh95TAis+gylvKCbfk0bb25giedWSNyqeOlI1zSu6omS
bnFNJkrdl8JgXs9MCl2NCwc+fP178vNXq5s6ATPmSpSYep+5jDL4sNKdaEXmplNs
ybgZ9ZRMhyCFZUwblfYBKfw+mIUJkCHHffbJSUcp6xmMHPRKJlthrOpmTcVPHOPA
ELNQqAxb5KkPjAp0Q7fpKI1mQb220eOrRNlUpGq6xNK0NCAnQQU3+Em8wsbzBBdM
+Kjs+sgPynyXIccCYkec3yTsI1tjv7RTLEJE7pgaNw7HmrNIv1TTDUeSQa6EgbQ8
U4opip/u8qsMb40/mSN1xWU37qp0y7yLg3nsBRt87zVZI5qvqO+9M+IfqscqymNa
9/sDkohWqy5iqMLGqRqta+e8aEH/wyi/unhotcsSBeQr3wuDHKHGBmcAbtCP7zZs
urj53A3hFSMJ57ahMpa+KWGXamQNC/aEtVwvTXvcIy5MkvgmVVXT2n/HCq0KKksf
tfdlDze4Nn9Jrc8Gaz+0G3bgrX5Jio44K1wfXK+xEn1Sz0H0GfxcBZegwq0qdwSe
o9H277emUhFf/xXgNqgphLog6sWeH6rBmTZxJ5N8OZ+PptRYTV52esq+FBuKItJt
TBDYK8nnGfkR54Nra83PxcQZhk4iHWcsXqaXZIRlcf3L1utEAL/1cUPOwu5UyX80
EzzJu3XNu/ZdCpBF+AQWOiOFLey6aHYHjAHMIVizFRCg9HCUtlWlStkGJDfp5bBm
q2HJB1Iu73Hk2DaUxFUXkUoY7B1KC+7SEhRXcP1zxcrKwqXr3MzN1c+W4/t8Kkfm
+WUhdaXZ7ZEpySNZ8PUhBgKIAQPRFFDAIGqKiLf2CBB2tkEqX/KSkwifzKrUfC5f
aOBW1pmKBF/fRRSHpaArI0OL9IUWJzNtw6zWba/lIOyUCARPvV59zKo4h8UcRIsN
8bt6+khzwoxzosLMV+OhGH9n7ZZTkC+5+umqH+AsC3rDKDFwuKYBGSm3+1ehboSL
qHRk+jYa0tUXG9dykkLGr5gbomsGbLzWpVaxbPLiDHkdOAXy/w2HxwX7/8dNqUez
3ajWozvXQeFErqNw6PB31xIOIASL8ZjZBUXF9XkvBQm/+k43Gtf4n+fHFVOSgyWa
1tmIdCLv3BVzdzbfEohBh6fHZWqIAwyr9lcDplJJqwvCTUu1Kocvl/jyViGqAMC2
Z9d1E8whSOrocAd3OM+XlrSfJ5wqvEZ027BmADW6Yr/pMnNKRyqbNidjqn1upc87
eXEd62ciRvNydotKXXiP+8VgdnAFUGic24O0Uk7zkH1KF3pmdO6a0oG+Z9XWXTD0
D/2Yg3WIXrZxElB+UdNBPdk3rIpMevwU7wfhfCsHzj8mFjcwwXHIBDwv1FEbCnVe
4Kjhlto3EITrsIYnpvHSeYki+VWp1RlFHye1zvLTpJyUWJvz5dlDrAJktmIOxU0l
AQmXizew7lU/OxwOTcc/VnZ2hqE+I8o3tlDDz9IZP7Q0/nP5iZarGmRSC/Kua0f7
CbWQr1eKDrTqooa4wyuEapcr0JGC8jMTC3Ru6KP7XVPmsSrfTgK2lXDSzAjkVofd
kpeu6ZgpA70DGz19nhZYSjM6nEu1vcPKwpQ3bwnXcpZaB3RTNNwhq9Koj84nUHCn
PR4JFO1/ICxQ+IoXrJMgq4CP0EXsajIjgJ3U28Fw4ZJfuniLuPD5pPmA72tN4xRY
f0rt2epExKEmj8Ac+ccvZnoDTqil3uSCK1XUUJ2skRpG6UcPJgNq4HHJ2Z7GAkHr
XGpuxL6l8ulmmSX7KnFnpezNlNYSH+9d/e6Yz/N3MLwH2lOwilfbvij9SQbiOc6j
+HuwrDmXV2O5O1x4UGkW5tF5kxcf6ANKYRORvGDVPT0Xyy9cH13zBNe5zkrertj6
noV7+lOcqljCvFx8lLFMfEqYkQHPdeTI92E/GpdFr8nDQvR2NnjzI7017/GIOu01
WtzrPQ713yP7ImoeNXaeevnIdealA0ASyu/HDd4GiZN/FGoH3bqsa9Ejb+0oGabj
NszO1cz8cKSgxZLqXFn6VpAaO2Mutef+w7Eoqyg8nLv+cbMuoxNfdJUdpEkTkd4n
NZ7naheFkUgx0Pz/p6p98NMYlAPQsE+iF6Tb2SzNjOlHT+E6I7iHO0zFqaN2GN0X
MZZaLQKKS62UMZcHT02KFej1xGaqrWYDdcP6fz7OBFFunJ5kv1e/c1sg8B2nEpVh
fWQSNDHiUPmFqOAS2itlHgTpx+2rKYCFMhGypL/V4OP3uCifDljN2LjiFEEZ6jvy
6xu1NHwY2sm5AFGxb5Rght6ENRfGyvANyG44AzsJxltJJNQidDyWPR36jaQ1RXOD
D2+IQ6W99TV0Ok4xy+GFYVOgAn5RNO5GFrBFhv9IOgvmJuSVOs/kJFuivLYyzD1m
P94Q1Jckd6oapnBRDiQoMqLImDhGQ1XxSU2Egj9vvsCt5f1s/WeRmYsgBlxjoap+
NcsTb77BiJHGq5n4posprGk6N0S6fD0TIqF4RlpkoUWyuk4kudHROxk04rNP3Zq+
JZ4LITrMoTDdXo0gkNMFvfjq16ONcpNgTsgTA3OV5k3YybWG+GGPiHnDfEr2BOHs
HaLXgP4uJV6jmwEI7yMD00d3uQd+e9exGECSFHTDLMSL+BYwrLqVbHpU/D5JVnlB
Bl/5stXgxBCr0FlvEJNDJeI9uOvChx09VIVdVP2jO/PpTv4PP/shfXw6z23iwIS9
+hGFtaNPCbn9nh6v2J6Axq5VuWWW6LpEKi8YPA6IXEtkH5ZmNATq3JpIupz8uSE0
+u04SOlysO/+XXzHbPmNuJXFtzlgs2h/04h8yVNrvvY2R2yDgPA7WOXaB+Zf4Hf9
b3baYnY58vJLmeDCkszIh0Df6lJQCGl2MpO5XqgXUdW280MvUmJWc1ISCsGtmirc
bI4ph4VwjgMfv5xGj/N2WqSQP58MTQO9zTx7LKa1celAYGaPILrwTu0djE2E8005
5sDoeyW2Gyxf/rhh2EqW8VFml3oybbOW+x8Qk850RWCdYNU6oUd/qJ/ZD3Utp1zW
NFcBEZ0IHbnHDRyf6Jjy1vLblqjXoIFgYlC4dwP03uFOYdhcuna31MIFzxcxVZI/
usOxC/7DwpjRTa/pI0uN1VKvxc8vN6bfiqDm1Wo4UCNhvBwmlSrIp3U/xOfRG9kQ
LVTAgv98TJi2YBn3efeUgyyYlRR51BV0W2bWQ9Vxy4Il1nxpwTOQjfWJToXO3/rP
Sxr1YRMIopfyDLMiLWcXYYL3VbYevCrVjZmSuXOXrodqV50xJIPO2IR/4J8yAWg+
eYsN46S2usTE9nKpKGUATXRD2ZNRBJLh1/1sCfO835g1ojKq4tuZiGO/O3+lgGhd
gPANdPLm7QqWKlGKRm5c8KCCqlCWV2cxgZ1SpWeJHZkU8+0KqUosnHYEmMxRBRdI
/GxBW3nKTJCnMDvwyEm82tvfwoPDu+Xg7Z//j8b68x16VZRkSiGCriGc9OrRq3DE
thiQXHf7e74ba8o0qMoW8igIYZJIAbbfak7Kg3qvyQicODD2wOVdzSPlDpIX5mgQ
dM7X1AsNtr/GGuiMRtPzP26cwaQw/3+uJirrmH8kja9EqRcmg0OkWHZEFi7ax8Ki
LwcVJkRlT8Ej/gMwyDEH3Gk80xXUWX2Mbvnq9Nhs7rBhW3XIAfiQvctra3DnQMc1
s4oCrHODY/Uk60kWY1y2g4xpEhwD02krpQgY23Hm0QdYqX3zQhwp4B5p2hxjDTPF
MlGyHdVuAXvsUbQbqPLecFXwvGibvkDMfT9MeVYIE+4+8Do7H2Rbb8fSyM1ZgqFf
aITYc/7+qK1pHSEMhi2CCnWJB8x2BsiAZBXt8GrfxTlslpg3m4zWy7OfMqJcTg38
hobteerRrIy+7jZMeXv89qAmnWwMnRt4OD217BRyL3SqsCRAL8O9pD1sLdpaU3as
12v03o5OM41gaYRizwFjYhZI5H/ybLnhibiaDbbsDICxOq23SRoRg+LfcSMra7wr
Omofof9AXMOSK+3K/GdjyPezyc5l22LKcihb/u6fTdblfStXNeZtmPAAvVFbxVik
HcWOCS3TBPhGk88GH8SVvHVGoD4AicrB+7NoGqWAX/o/OJJb+w9OeNwfhPvLshGN
5wMIWA7lP96DQErFl5EJwljH2K9WyWbucH7kKAkPLTJ4oOInAHh9B11pqD2kM+VQ
BT3PjZb4+C2ffWwLkBdITFwvhGECJQiX878cdFcgf1vBS5PPnEP9jNi5n2whMj3y
LoNOCjrPgmc+mM6zR2/zCse6V/CnL8Omvy3+OL223k48Xk0Ww87pA09gSa8DrQ2q
pADHreya0e5ozcKnL/3VfKZrfLABbXy0AAWuljyjcoeeU+z3l6mKkr9S5lY7Hvya
eiM448u4OcCaw3LRRYoMYYyajWdyW/oLrOPrgMVkCRw5OlIq3VQqIFFMVmmeA51P
qqHc9qb75wTq57O6RVwBaN0BnQ/WnEokhexmMyHdSYW+iMysPRJwNG/4Kzj2bFk2
SZoD+Z2ZzXaZ/ejngJAnNlGgvDjixr+eJ10CUGUbQCby9aCCEtPdvCxfi+4GkyIy
n1Nve94CuSIsZ37KCMAzcDkhdkGCShQKcHUHRdy8yIpbIgnKUFA88psIuVgw1qra
/8Aba1HPwp15HVk2gmsgxxNADlftq2XTQxUasIm8i19s6JI0RFTUCq2b118WJcAx
n51mU6/rIRjPOPjggkU1mPIe8+PfqkX5jdihw2mRCqYj4XwWNPepYq8IqgByOLS2
RthTjJfmoJdyUu9KWXPJ4MkJ9eDYHZApkhSZnIrn9z4bhsGFj8AJCWwyKrpHbcyP
3CtiMDrdy4EZV0yE+sk1+41G1mXr4LIsu0hmNAwFyiTeCqPxRWKr+nJYxBiNHeJX
Tb8Wtt9AD1ma5rqX+gon+ZUWia4ryJ6CvHI6/C3hzDjZFUJ/XzzcfmUo2bZmncBH
rtdp5vD7sapVAdquoum3hIYG9vCggdZcpVQ6XFpkNLhkTURTSGWriTxndjwnjAx3
Zc3cN5ZDoQW3+B5eOAJNiSiHy7FVwRTYzfimc/Ltj6gU598f0SaNfogfV3SFDMSH
JtDtvaJBCBp0panTNiJxyEuuxDheplU4FZmezZ80J26GMMyBMvSVrA10af0tbnCy
xCreWHt84d7JWalhucBlpHBIiOcmMC7Ot+zh2+PKCvQ0uQB4Wa9kOknD9B89Ba/p
L6yc7jODCzNsvzfdMsTtPPeir7+YUAh9KclJV4zLm57/s74HCmS/HNTsH3dsXpmU
3gBjjdJqgo21AQlqVyGwuBIMsq1T5r1ElA4246bsW9yWf7a8Iob5qFPnVvC31RtN
jfqHP0neDYT1X3snPsv55crrF+jPIDSq59Z79dbqXllIrIbtZYJZDYm3HQWF9Xsn
QHTwb70ictJempr1ZjJCaM5ZNA/La1sz6s/B17LUrb89xMZvuyreDVtfSFkqv1PI
/ukRiP80eqj3erTUP4q93vqbvPGYxgfgTVyjcvwrHZFPg5QUjPdq9fF0+aP9vNkP
LyMv1uHumePqk/4SJwnRNAUD7FEZtU7urHiMGYJYusDRCHka1jGP/T28fxCn3kT8
SlNIFlRHALziFsQf57FOK0xZoWya6s4TxB4M/Pd1SiyMlcDck8dzO2wtQTVP5Gqy
ziSmGx8XYosEnuK5ToqZDdellBAk0+rOKkkZFQd23IjCsbQe5iCdSW/JpbAPXLFH
K8FwWNWGYQDJDYNkiqqKsm+pTg/e7bhdcWuWac2jytePp4q7K/eEmi0FyBv0tSw6
aJ47AiUn8AWItKiaSlHplML4ullusAFuOjHSTFmIgCbFvioqMCwkXBeibBBYOZ6G
DOpGJVswwOMevylvXvTIIQKqx+IO2XZ2zsNKSbTQRgJ5irrdKrW2Hum/ddqfTonE
puvyO3IKwoDjJ+Ght3cYbIlqPuwvMMV1iL+1qCuAy2FkOfxdBx+KuH6HbIbAbjKf
SglO3RLi8PPi8VVDL+x9HJ27Nebhg9MD/BVmHB49wRW3vCRl2aqIXz5WdphSYnad
RrDeJfgoPdCAuJUPtJ92eZ3Exns8Tm4miZmAJor5TTCcoF/jszKb8FdSWTRJBs19
kaB1COUBPoWD6xScMDo549WNuZeGTHVUP4jV/09viBFuCPd/vS3NQO8XzI+qAy3S
d3W6eYSvONZYuAd/aq43Ee/olhUwbF36uCPXmsqoxX07GgSbNJWb7tcq+f6NQDQu
yDBU275ibHBgHX6UwxdH0AAvFAfJX6rBFb6F+li9XB3V7K+j3mGxBEVO0zyIpDM6
9gwM2UbEH+khwRFhKI26l1QjmZ1RFy5/AOPVf6pN0eN3jXzVJ3hVOfysjUtFWVOR
doa080f/S8Hfnv1XKL5hqHZnjiI2srMH/yc18tNNKzTkYxnuKZxe03TW8CBeW8Qx
ubPRQ+IQgFOz/WUy063wxmjGPEu+WaEDt6k7WTE2pB8w2BRmJgA00ec/jpNJ2K1z
Vg6yCeJs/hYpGfP4DlMOrENiGOtuf2+zyPfz+VkQdLTrqF/7WMwIwMMogz+g7tJ6
E/plz4cfq39wy+qqYRYLcMvsdu5fsY2BQp+h6zmstjgwDYwoReKJwSFZdkGE5kaA
gZsec+z8JpahirQlnLKEXfxsI3XIYu4VLSDNI+0L1hZeNY9jRumXBQ7BYssOlFCA
Wd/gcztcckxIc1SjI9Qq3qQICBKVo4AvVcmCKqxzct8ARtVNK4CGoRBzPedaFNqO
4ArX7qhzo/VAJb4URbHLwrU8H4CZ6Ieq49yEbdPFcv5fFDAZBAjp3ZqVRmktSHDr
WayR3o4CHJK/jH1Hz54qMvz7MVC2ClgG4uMa8JAV1ilvY+uWujTQKYb9W/RCfsaI
J2wWvckFPQFfbzGIZLOsnqh8cI3XgW56SYJ0NUDnDGwzIjBA+FyU84hpD7LhWEGI
v5g9wWX2KhDkZZOFshYC+CtbI3n8D5d45TnqsYNoVbZUJJ22OkrRC8mQK/9lFGVD
qRjA35W/mF4KgRF11zxOeweBrlPuqr+FcU0r3IB+sMONRksNKj3blO3eOFArZOXh
FTu15FloPA9bbLd6Lqc3CWqzBxW3Elt8LW2TF/aDgOzb7ppn0l+BTfZR/23CQCyQ
lMr+B35ttXNnDKFHN8os1SogxjbiPxHSjRnKjoao9cSAIjMCasBob5TIaSaeX6KP
YCC+hctxzbjML2FGpAS4Np5EtPsgUZUyDVSC0rpx+eBWhMA7QnIDPnqLiSwcMxSa
gZFB3r0vmsV5RgX1NybGz/gFk1ZnQy1FvDMPHx+y/chmDVzKQ8Qdd6gI1GCYXhyd
nhQcT/4g5OGsRS4HoblvfBP+M+xu6gVHAckHv8DzqSzPPNvCVvM/yobFQWXd2/SH
avP1suJb57CLRVNV+9jGejPh7Onw7y21GkNGfT6NJloFLbSw67gCCol2DcCBXqZQ
DgyrRNBStJsCWyq6g6m8A+z3YNaZDXI2LXQavgAXJR45P+HiMEP3/H6WQ6RNq6Ll
tkIrlNNFd0DZv9gIhX7ea5kJFkjOjnRLu9m797esFhC5f4nrF+CphF5uZqN35owt
+jAr/GqzgJKgMsLI+iJStOZOsO/adaseFUhfHkE9zXJY/Jl8lPQfSn0MgiiEXHcA
CltXtiqhg4gs8dVrzuGwr+gwxf7QSKva0yV7IVWxwYGMHnVcmC/n0modcOAkZlgN
n8+U+lEVPCJO3bUoElfR/Qu/dsXCHE0ZRwnq4HEtYXqhbTsPeWnZbA6tiHnEQLDl
K7I7nb3Z+0r9QMQfpr8F/zg788REKgt/pFhx+pELcmcOal+jfdAuiy+ahAZ49QJ1
Iug4vikf4hZ08Q6Jyv0fXdsGT3Y8f2T1dXIvqHmpS81Y2eZca0LpjBnhwjjXATkI
DRyc/aDMa3GcYAJunCu1I9L8ce0Y7qRnUv70OOuhDKZNMroc8JieuNR+m3B5eaSI
Em7/elvhhJHfjp3X77s/dxwR5puUXkqTBzljm137rahZAJVJMSipDSZ9bNm/E0i/
xybFsYuCYpc05Uj/zYQ5F0g5XkR07HYsBhAiZ5sR4mYTZCxauJA2Z5HAVMmNQDKh
SwJrArXkRW0OB/IKFXpRqT+bodp5YCso71ye1p4tW3850qU1Y9ISHCdopbtiZeo8
WL68aKeB+27vkfmNkokri84C09x39b/VwVAL3Kta6VYKKkiR3ftpyC0Rt0bIcP5/
UG0dp/cXZWrehKDxyjT4U6oIvhIgYfKRqYfVsnUMu4lNvWVWuB8tXhepb9Hj7jbK
v09fd8eNKY+WtngqcX2Xyw61eUSarucNj0UdVD2h7W3jl4mnlntYDgrxXD/sk1fs
/ZQoMnMpOVGlP5eI9hckP8pSqqa05glIV8fJ/gGUeH31swF1cAyeW+rxWd25M7iw
FtUYVzvK8egwGihwDNSbqdISQMsUQ/ki2PbsH/sciGNMKWC3A4eV5UF7eVGmZ0IP
DgBAxZH4TIzMCJtolP3lYWWztuYdwdDJ8DtBMBff+jCFKflgIg/7auQAgnz+yart
6VPe/mxunALVPBXoFo592dfZ/k9YHXwd+aiK7W4vuFGpVF4SqeqQ87CvZWwZa/Dj
aCwOtE10eNnhQUFCCkq68MPB0+0NbJxNtJlzwyzbgsNqUuGfKxAhYo++TmNykqo0
E97hT0uWHNZMmUPTWIsAKIuCfq2HSElGRQyCfxxiHBWXY18XpNQfLLS1i9OEQGb7
lzjSnBOIhE+zwvWettsH2Cb5EfP5Qsr2I7e0AXrZhsTq/rcNqsHz9a2AoE3L3l/0
QthMn6HqqTShc82KZDEoo4+DHJ07FWKAETOrlM/kn37EaKAQ2cLpRuHiK5TQd/p8
qXusU0Cdfl1tBVrdfaWvqftBz0yvHl08EJ5Dij1ggGO6po1RVo0DMwKmlHUiOY5H
QuNbZ2Giv26+ucQxJWVO2Oz3osHlgmmldovb+U3DgiwNCSsNy3wROvLVAhKGHlIf
FGhIZ+LEv3plWMfiEQn3+sXnmNF3X9XS04V29U9m8cB6vNhJNXJMQ+icQBHHiO5c
/M2o9p7v9IWtc4Y4uR+Cr0k0C3OXUAWE4ObAm/Ih7EwyyGiyJCVv0mp1RtpY91WX
m2EvRetNxcou05SUwnQMIUfpw+JSrJrsku3xAEK/jTKs9V1S3D7cKISqrO1yoIWF
yUrqUPspg0y86r8KZSkYyWAzPocc39CFVLc2IME8hP5+H1mtSbtEagzKPMUOXXkq
KrSyV0K2g2yBzhoKWm+wrzO4bln/Lz+LmBsETB9EVDJQJq3/e8elrKcfzzKuktxj
wJim1XBZ+E9rGpqhlNniM2R5bLFpcBcbkeGmjwv/+Slog26Io6iFtrKT3ABSSc+d
NFPkH6j9cZvW3Tbt9Hnr7ElHJHvKLSyXFHPbpiupNhO2WHAZJ+J36Mil1igVRvhQ
wDdltfhjmB2fiTLYLXz95UqjwJ2pQzSRPrHBFZ+vkZ0wBQQOttY78MxPJcrZ3QOE
ZSG4+y1XtFhsr2WjmkgfbomHkOin4cMDib7JvnXPjUDk+Ex7J/O98JZxUHr7Isu5
ezRaG8halJGPfbDPkAsjDoVUh09gzGWGsJNYKudnsDDZ63iOzfVd0lmZK6BN6RWv
Iefok4Temgzq0uvVpEQulaFuFpF08+1JnDIKJ7znybovW16Dkiz1ORegLjT92YMD
KToHmZhS0GHm0povxLBHbz/I7WZWGAFiQcMgUBwkw94ZrQv+45yofUBgKNqIpznx
BFXiTNYSfGaZvcR2ODaOb56KeA+WpcF6lmtXxmaTPAD904l7ub0B21EPbG9AUMfs
S3KKv/CtGSAgqb3H0G8iJ1/65aDw3tyxAmpRSbYBMuv/WKPc6yv05qgorFOBUy9l
mBEsVMHC6u3yZ9svmaQtev4JdYX9ryHKfpkqhVhdpN5XiDdydIl9+izEKprtaK2x
2U3MM9m/tsVXqPf4uD7PydH3FAcFN2YTzbdvNbGfv50w7Jle/m3/815S86KBm6ay
hi8mErBqTW8Ndh6mdLRN92PaIYhBG5daQUJU9lBsTFn5mlHo/Tz1LHAYnYLEC/E3
W6oEyixmI940TNThtqSU0NiABMVvUXBkxYUfSi8ICD8GNs5gCq134qbuCrzFOnMQ
m2P6HrhI1EGYSpSNnljA4xzJf6g3qQ+e4iCFIxezAdYsT9ruJ3ru9dE4YY1G+3MZ
lNyt8C6TlSsklbyB8uQw2tpnZXGVcUJ5pIm2K0ZS0R3pRQmS54+VdkjtBYf83biy
30jTUFlkN4Hk1xpWA/h6KCmDf4f2xu2hITxa7hS1z0RcM8qqh/2STJzqhO3U0vfE
o189GGLaPG4Rsteu4TNtiwAUdk5SPFCGRKmIzDp+KFb6gb+GQNvY1NS91EnCnwqP
i3932RBMuJsZCzpTxt1bvdxxjwDtfjN6jtBOU69qxaaQCL9AfwOVOWHbCkh167dO
5JpdMU17Tr/FFiyL9NY3aHWRidoaEnsZpsnXEp9nxIYx5ZmTaDkyuERLU/i6FgQC
ZPYHmQCn3GjgeM0HC+afNsGG7pfYHr9imhs1raFZ9fcudShzzEIt2wNVsmwiSZRW
GqWhE7ylWxjTfIPSH3Dz5Li0LcDVxHOma/rZl7GOBcSvtNTT2N9zS2srrvRxlwqm
sYD2FcoEiguAKOz9ep1Hcgk0+ebDlq39nINYl8/wDa5BP6T63ulh5/YYfwvOATGX
4kA//SZ76r5IFOxc3bmVCJjVft3OMTlWHQW0PoBS53ws+mljjtW3k/MzHghenqUH
iAwjECMrPwORHJTHgPPMOgczUTmj4X7oUzIjUrY32JfoNzxtl0tygy46XukWzczs
R6Q0+mYI9Xq/sQrB2aX+lBddU3FAqAB2+t7u9TTdg8+i5LYfq0MfpcpZwUokiIlO
r7OfFn1ABO4nDHq7mQ2+ohL0HnSAMh8Vs1qhXT3m70kBt02CgOfMclKXCmHXxaP/
O5pBsSILXjfimv1D2Z3KQN063VwR1iLYFaB3BHv4U1fzTP/LVFRRsng6uq2VGBs/
m40gz0nFJTdTTixli9ugaexh0P+3trSlHWzVK3GaFhSPM+0UjKGqapqog6+H3GTb
ta74vOyfXPWFxFSkIEWiLKSM1V0DpxaLUK2IeENCGDFix8ain0dDK0Ekt6OKzh1V
VPXXeH1f2rudXCvn4sh5Y/q3S9WaQUSZH7gPu2ATQ9eJ3bNimFyUSQw5BsbIq44j
wC7lJ7x7iNdSuEjF/DX8PfQlUT9fG4A0DdyT3MRLAXjPmmrtm6PgVFjXbpjamAt3
/ri2XZWT+mI3JKFcLmTofOtYKWLD6jENB/Vud4f5UUwdPJquX4yJQZr2SjdB9Y9n
AQ9ISwmftCjrVTLOaOO1YkZF7cDGa8NCxHa+n9gGHxEQDZ1gDRiMQupgOlThMDhM
JsG1Nnoyg4DvHiDUSJdCXUX224ZMA8I2f6kTaRRsGztrHE8ivLtXQa3geTLPu2k+
XV1ofAqDXPUJSiJZPTU1ehUqthUiDHOEp52chMWx1KIUBAqsH7yto1aMHAM9xpG5
KWx1KbZB7PQjLR20GNffNhW8VRGCF6M/haKM1kdtyDHqKY4GyGhEm7FQ5sXqDn5d
d+KI3PXa5Nu5kZ2U/ASq14E7ErTvJh35HlKcFW0mMDKHEF4WIbRGxIqszHMHgXzY
P/iTku34V6BUTnc6iBCrhP1HwY2i115hddmJEVA4dBvQC/YvCz62JcKb5sebAykb
YplwagKNC/opTYRZTzSfWJdkU2dXVMJvhhIhENIr3gK+QLLAnggET4lQRkExwpUn
kqbn7+ZeX/iDpG0HDIkQ/XwjfSh5nPbfy9hoG4ejjqpB1xnMnW+ODLQIReZeaN2L
Psi47wH0NtxuR3a1CKnsdM8NzWS2L1L4EY38XMas4c9WUR5bvEwjkzy3jlgR3iFn
oQIRB2uNJQgeaue3MVv9NLo5WS6zztuhe3WEUeCc/9Q65xlN5Pg4CGZ7uST3EkSz
K9T5OsaKkByUHhZsKxSxAMcvG8whYjEgu1PsswvcPhsvbnyX4n/lm2a0CtXL7iLG
nUPfbmNqxwZsys1cGtoU4C8rmrrHTUb5l/34LcKeiYG6TtHZqG3DNqAFH+XGukfJ
hfl+okXp8MwGoEDI7jj5cwe7Er/uydkfDvT4MkPoSUoT6wdD+BiGpEoSCCWtOQsa
ejBg8YlW7ufHuYckD2TuweT8V2EXJ3H6buNNsMDkaXuec0uxF2TeRJuusupfbUlv
2nKZ8l8jgaZNxcQG3MyhZrCb+Gb1vydWQ9tgPnd0x3mmx6LOx2FA8qX3cRGNEgvC
MXSgMnpUC6GzUdBRN5RAGpuKnFY+GPo21xmexxPEXMPWUXHd9214zqprUQetlyKS
Ndi/Hz0Xw296wdO6bSwuZZM9Wo0wOcnNSUYC0zjAt7rpalFGjt6A5+X0JEVzRhMk
jtQvF6NPIBwyhx8ULBF0ZX1ceR+/HBCc+NEoDLl1O6QyJASWU1Gg3XBP88ON3Y9h
SlrcP8WZMUUxLc8nglBtk9Z933wN0PPlJBnc5CN98MoFSjVgsCskteog+mYsbljf
QqYzxeBzwCzR/+oyJqLCiWn1Tf8MR1qgEtZXfoTrhGrjn4fZnfZttBgYnY+luCxF
WkSLtFpdnKw4F3R0SATgriQeGIpxNn003ArM6HtFjJVLl+d+6QjL7COBzslZt0C6
7pBVHvWWtmellaXS8SDa9T6niA9CetNgSOd2ml+aA81FLnfgg8IYUBdR6GTrrUNK
xglNB/dwVXkOlcRX8bxqdWvucl9bbdxHjcNC/PP5wlGsdHDrgaxAvwp0arXpNFVv
lyl4NytDzPWrvN07STEtOVRuNxu8rbWE7xqHC2lCKJMn9Ori9z2w4TtDhultulMZ
KXhZW9yuMISai0CM/cgdZfGY2eO3mpJvsM2BFNcHk5ByAADwKpnQ17zuoZC69yQd
mekTY4GpFbbp5Xs4JLG92XSq27e3C0jKefymmUTq35SLAUCvZV7gkqmQkh/ulayo
P3cfmLSPHsqEye27pWFwUF4MQHB/PN9rXSBrdZ3b3dM930Xi0uHGTfGPHUuRrOmI
/g8odljmr4omon4HLWAh13/vpj0mUgYZaWztsopxsNPuuCmROlxRZZ3ybEjsqFjx
STx0h8MpKckUHdiIEsTwbeWJCQMoILYRLXT7Pw6+4zKr/JTItmHLwJJvQdhjkNyL
P2LkqTUa6HQHgkP6dnjBEu5tq8D3F7LS8WUyYH1Ywwh9ki93oi90UZxf2979GlRR
VYk9oa/t/Y8oIYYA9AODkXRZ8e9VbdUoff+bDHfN29fHpTP/K/Re7a+per5Csea6
P6AbsOT55fluRah/bS7NImAN1VtIefoqEn2r0QA4dRkqql1KRMjllTnL02eyskap
+P6SystnIi16muTzVQGpV6/gEPSCf5pvGK3rELNweT/hzceF4rjmHIuPzJBSuIlf
9+CnPj4f+izu1ZygsFxYB5V5BKzqycAW74AW/Hs6XpUe4NRenZI82nxNOAN6jF8S
/EO8iDqd0sRZ63GwZ82wlA27uuyOXxxK4CwSSsE6fyyS4SnmUGYROqf2XKzjKlmZ
40+EFrvO1HYW334MzhanV/8wMasNhW3GsO1zU7ZA1Se3nwF995Oj4oxJiuHJnjLS
pZfLtXYqfucjUIgECE5IA/7nLmA1hD1s0Ejum6CmvGr6xahM2+90FmZAMgxdpcsw
LLMsQahLZPqsZovBo5Hwut87FE9NPd8oV9xieSiSTykcw77T2IowSB/ayUvF5iYW
hYrmM06ELkKVMtHCd0lLunsZD82PcuCzht/It6TShLs0DE3JjnEoarG1pWljoPdo
5nB99kPt1I6xD90G0cRL269iU9Cc7fgqm0NvaiP2Catk92yybl4lJvLnsVCnBGHx
iESvsB+nJLyRGYdZxIT0aVd5FPjVaz01/XhE1IIseD16MfdMzsh35awChGguGqKp
qy5AhRspcxfJ/9Esp4ZJq+1stYFoSrEozxiaN0mhyXyPecULd11NmrD33jjUMNdp
7O7VqYelrJ998OT4h+LDeVVEdxZHdY8O13ElTYggraBt0ExXNcgxTN7BbFDxvELC
AGPo9YKZadKWqgcmlURtOmpX6CU/yofygf6C5ZGMmvkI0ahCZBBvtC6O5ttdAhgi
HOTTuAOrlsX3f7XAiav0M/g4wJoURnZrVoMJLOMrYsBtSQDpmC4BFQCXoaXg4RLA
CE+cNxXU+QedExzQ4bWxTtQUV2tk6LfITkjmmKK+gyoJKXod2XHHGdjS0uIf/jtt
MGNB4eChF7bkDxnAbVdABsSRl2e2RVD1YPSgwnzWw1r3jgHSsJzIdv65g0cP65RB
K2PZYdbbyTHjGvZAIQyYQmuI+WmviafbFV/1QarPwvos5xZqZSO/9c7SvcoF8E+W
rdunmfCRiidh29++Yi+nzFRXFvsZDG1640FSSkgip2HAI9JrPoGln3W6LW6ANw59
ZGV93NRZV0s0GgFUUU/W+e21QM6WOezaRLmpbJvSlW9a6mpRde4mcB0SdkMsciPD
CNLBmtEghPqTW6wj9gByMyTDzUUcpFfrIMq8por2zdVhV9DqHUQth8PM9xwpIpoY
YF57GOGw0fMq81M73KXaLAOaAI+embXfi6YeajkzT6A75+6kjX6yn1bVdPriDrnA
jmaRZThpqJ7+2AG7HHq4pdF8WoqdDCosJiKsGNkQx8nSvc1U7QmurQfnW//WH4oT
OX9F7rEB1wMfsAYzsBLJpWmQtiNu3+wXgHFPXRU5pNJrKkoMsdtPUImNHcA5Tofn
Cex30Q5ZKZV8iRpymW2jeQFkeqeBu91JTJQVouRd1gjbtZ0HM9MgGgvoJCXdOOsJ
6+uliiqSwl+7QxXUc+sQfsy+cxCXPMvEi0xC2k7491jFqZj1GgFBDlV2iXpSMaqF
CfMbd/xvzQ4LoZeF8WRRa+My6/ITPJ+Y857E9V7oDlbtscRVHPyurxxhV5G5RoR/
FBF3eH9o86szoxwYR31EFiVkBZYauI5g2kyt0jxyobp+wc+ZgHiGGzSBqsy9MbOq
YbEN3L3OSRPApZ2ukcuDJ9qmF+fB0P0+xUAakPSnAmDHiq+gQlZpS+6WhYFxhXDI
IsS0tsJrFrdE/+BWocQUV//2GNWJ0D2unoL806IJGvvMZ5t97SFIKfPi+hHy05Ic
93Hzl308pLoMHCMJN7nGE+p5aawJPU9A/HfihpkACNm0NXVfjIwQzskYMuJ/drU8
EEPi96mUQqp3rk0Pp2sd+eIkcyNmwHB2ePCtT8J96pmE+1RTXpMw4MTuxFLoQ3mS
QZ25c+j1hMrZAEW5TYs1FuXixvMSxo12rXdsTmprYr/8UwG5fX33AOKnHTQGVSn7
0qVQQxPvRGYfALobjSe4Oj6Ysp3AA1Sfp5QoNncZSmYPIu8dsb0/o4HbEAx9a34M
4fBE9+Ap8oCH+/KSlKFjhcNEmEuUeF58QIf4/0PpqLbgY2UqO/RPOgGLT53xnHQs
u2iCUqZ5IZxcdHdO/+IzvUNuxFsr9hXZHVwdmfNCgODkUQdKEHVtYkrDI25/rIrT
3j5ONAk88ba7YCXs1W7kW5xwf86yDLHSwhaPmoObl9q2Jxsb0AffNklTXFwLF0dD
8KbsF5kba09Vhfxf6l+GqaU+5bKeefpx1z8kOqs2hnY7P3XytoSD4tWMfk/kt/Xg
JtVlm1/Uv0JpG7FJrW/iuGbyOyYfUnnCzKoPTK1pDD3YzC/U86LFF68qJixeJUwV
MVp41t7ItvU6ENU+knRO/Xq+Q7EZZqY6LcjtMckCscCYbSOcbcOgwUVuy38nCICE
oBNZ2UYXm4iNV9x48B1+/KKXo6+I0vxXEqn2TPa23zeKpdvY7cwA3Ifp7lo6tNBx
8pY2dl1eL5kE4XbrN+ReMIDQCWPv+wFdFn9+kZikoqOfQeRD/oPlR3VEMhmNUyN5
h7ok4/UgBcK3O5+f61qmBuNQhW9NgMU68pYkyqglECxnejjZzwLn1l4lGYgPQQB+
5eplLLlAH+7LVRQyZagnBnYmb8AFO9pGAMEXx77By/i+lsIXCSPu4biR0fGZomI4
gvbC71bWapd8wVt6UhsGh0XgwMo35UU/1AhlOakUB2qFOr0w+qHnPFMi4nq5iCa5
`protect end_protected