`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15664 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
ZIICkMu+S2rq/yOQyqhpuoEQW8xstUrtyHAjlB5CqWm5GOXMQzjvklJlEdpB2GAC
JyDme6h85Z4FdQWmRPLPFs2FqKQvakX5cWflFejpnP3ojWGu6nA5tvqVAvY01+bY
Xk/Yyk/0THkd3qROfztDU7BJEeU3FGM1QJSgyeY1PRypJaTHaH0COZ2CW0DyGumq
S8QvgB64DLntFrNn80nd4AZH+HNOOgxspsBe3Dk/RL6RaMlBThGfrgJeeBfykPKT
5rhUISP5fSfEASv0qpJ8JaEnHKhzKgzYGTbEjDckCenNOALN9p5lyUWrtSGHVzFW
bfehmMEw2ZApakzVU4UOy2UlCqKYcHY098FFYRonYF/Y+2O38LLEmJQ6NSlfVJFZ
+gzqqY/htTmaXkTykKrzsC4X+25WuBBBv+izvqd0iY0ZUd91D/2Odk7c8FtP+fMr
FvYU/0kjVgAL0TMCgxyM6VBxpAI3qDtLYzZLRyPjpOcjR4tkJ5TXpeVbnZ1+o3/f
ub+s16L7gwp2IHNaCIRr+3KApdkcIaf+Z/+qEw1yoU+IX7ffLjGq4+mxuRJOwW8j
zKrly63wpylV/X6Ta6bgvDdJ8v9nIt8ytOMrPQ3bCxRClqxs4XaNZpUGHNwUDICG
/4YE0De5gc1vtoQRdItNZnl12YGBr1AMNgbiSV9UJon4/xh3GjYHPjYDLOlJ/qKg
fv2hUGn/B9HXOGd/XcAPOHg269kCj3vRHcrRO7NvMgvBS0spROUVxeauvp/Pn41F
kqz8nfJc1NbjdCMCzzk7AvAf95nzW5HSvKBAjc0kPXq4OBZky+Y1porOiPPH8Zwd
eB5Mp5oJAUidAn/zIldjxOpUcnXwTIMSPxBb6lFxS9Kuo/3SwIlwX3eQqmCmuWnP
E/r4niTwFzwDJA//LHqejhTgAfXC7wJG4Et/kxWVr4ZQ5JIHKHuOcRlQ+qkzQrZZ
qO6WJwSIHjG+15QOobMtweahyHOeS/oggh/XqK3HAzlUpfHWSlK45U88DjTWyTJj
BnobDtkFd6pklUUp6ek7Zpsxz72zLp6vpAg9gZrowTrSEynKGTE5AIsxaOOYtdQi
DwSulzaR55+1JGIMqvNWSyVbUJKGNIBXNYZiQQeX+zUJpBIffMbCElQXWgKBCqFw
cEbTjAeffh6RdxojUusLlyRBE/2x2BULUV876bfxxA8g1XeyXOlA+nYX4ScT+eYF
JkJjwAzxI+IcPEqJl9bSkUfiL7WO5o5tum3mIlww8APseR1+n+VIt6M0DDXa3O0z
dQsCsU3vOAbkbKXeQkk59ghg0QugU2MM6BH9M8ScU5X1OBbzWxJIgLmWt3ivq5J1
0ynGso4M4WeN0JpvrN8U9QJ7bppT5RiiTICdCk/Utk9JPcuU4tmZ2CrdGxuojhHi
aCEqSIvHFhEvsNnHVWxkrD4X1yn/gx+Hu3B3usfojP8tX9yB6MkeXlx+1QnUTTLz
pJxUQvKVOGlkuVr+osHIVsHQ/e08fqvpBtPqKvNdbexK/KITabId1YJSvXBMAedz
xcX66bSLWDFu6gd7USdNBx0kv/GlVQDw5vPir21PLaKOGBQrtvnuHKV9WU+EjL6a
S5+rymoQJUkSXL8XRsqhcXRW/0naa5g77Fqk1Licl+A9abqG+4k8CXd7pl+PBMhj
qL1AkYETxcK/7d4HLGRrc59KMcIFse69WJOqZ+Qf5jXjzRGtkwDxyKrArCHA6FWs
G5+OVBCjrnUAiuZYie9TfwfkttYKRqsZJWDunutUYZkXqvImCT35jygYKYVpnEXl
xRO3H4nsVDe2XzGmpI0ILv1tVrpl52B4pEm2fl8MpmRHdJ/LI1IDqCp9Qwm3Pins
gMRm0/JzpMFHtlDu+lz8UY7yyU4e0k9Bj6f6NV3gBaXEp04hLx9Gr9dTbeoCVBGw
VlL64lRXYjvfqb1YiRajK02JhBoDmg5k0i1Y8PVWnnOS5qdrEft+CSMJ4lqxXOiH
+2/Di8MQdK5/NJkiFM6xM50rQT+iHV1IBDcl4gS7+qibDC/z8nCb75RGSyqmauQw
BrsB72kkl8YuVNLSEKgGN51EjzsuwNPnDU+kawUcCY+cXb3BPEZh4RVaa3Jn4a0S
47oDutUDWFDBGBJ8K3wY/nEUZyQlE1H3/0AHL0jdQivs1eE04rs1I712mbIVc68C
7tnoxuCeDjGBTVYMjUSbDye5E26niKIB8tkydn7Xbt8CCCD9/rCuzxepzTDMmovl
91LVvcVvrcCilwUBHxSghWW5e7HAKz1DK/ZCRQLuAMgYhDs1GHyQxpMho5aL7Ydg
9QyPy11sI0kAmIk1rWP2M5ACP6eHfJHJo0TafU081/ZCdg3GgeUFjO8gegEIaiAK
ITM208sigIwwxUv4gFRZ462C9Db4I7/L0eOI0Dpvhu9y921nk3QqQW3hvRPEPrJn
GWGp9m6BaIuYk4DfJ7qna3vkqzn7KxjcfXVURLDI2o91DQFTSIX9+XnYxz8z1Jkj
IMnqI5Wl9/IB8FGfZ3NVhVqnIUX4BzLRSFi/DQbOHphmC5Mg2g3Wb/qF6YzgiVPq
IJxHHXL/ExrlTK3qNbRZBUNGqH2PlV3fe0DzagqbQJK4PtoNJcWYozp94mG5gwYU
qHYJO7voEewN9D7VER/UlHgpeC0DuPYq/D4+RNy/BxiNp/Tk5NZ/A2GheM5on8TZ
KamuZ89LlSy4jvunbj+jbaLN9sz2miVNvwA4M3vd6BAbrZuVdePAAPfZcr6eMKDv
t1VfcBfgSwKjf/VxqXe+o9ux8Y5QMFEmLwW3rGVAF/egxVmwlE1lFY0bawe/oscE
TSze4255dsKrsMK306O6qS3oYr25ic2uialMPj4ycN7SHYKE/gx6eetNRP3+HJ5p
rhGUiE98Us/8nLRrtIXRhx75z5GNjiWWBXn5YJPcEuZSdE0EHDw4O2c0ymKA80ho
/NGQv7OPeAa0Vqrpa2G1/i/6y6dPVOMF+eaesHf6oOawZYpVSi97aZgGIsvoljZe
I8gJ0SpVD34UOwPpx3NGG7StahBYnpcatO6Euil/1eGh7E93iC2O8LVkl66uQim0
KmS0TqWKcVknx/ZrCxs+TjVeKQNfDSbGaTCmHh/hXDiLDWOyj3QUs8Zi57Xu50FM
tRQyc37CNuvroOMCFPOAfZTQVJQBbKyi0YTGbmZT8R8PGqjMzRkTyiG0SzEiB6SL
lV3jg2U0VsZvF7j91giO/z7P2sOe1khrWrzxiBcg/nWBlPi9XY9FH9FVk/yhXMQV
ZUrHtMdyfJe9eF9fTHCNytiJZ4g7/iLTFBQLMmm/iaRhEpU4gSkYQfpwVxcRbrAD
YJ89NRdQBfq6JQfRckg96MJteRWVazW0lxLlQxKMYWh/MweFbzPQRB/anbXQdLJX
c4LpgoFElo4Pj0pNvstJkeHrFsJadfhtFiy4UvpwnLLNnXYfQaPpApclz/F7CUaP
1ehoNmXC5jWkIwbF+WEc+c5aAU53ufKTja3/VrKcK8g8Fk4CBjeTtxB9awKaViFh
8O1NMv/EWnnDs31U/YuCmowKnfsBH7slTd0QrIV0ZI9eanapoMR9X3gw9Pg8hYY0
25ClTOfPy8w2TSfC4Ir2r+ziJQYD4TfSI1+QyIsMIG20Z2ca1jNXoeVflwmIDYvh
x3xDZGtyeo0F7CMUPBvc+9vh5DVTEsJUE13i5izpgSPTGfF28oVILPfdkzPI0KqR
VzKouwp+1/WVLoltznC16U/8NCk3izjwMzN1TTNcIAn7mtRUaQjAzWpChMpluX1o
KeKdMxa7oTbIwaV1mJ/Hdlj8MnB+659iZ8aCU4h+kjfMWi95wTZPyNC08xbUZIWu
mpjHrBcAutsWzyRN2/UyqSgljoh34vOUY2R9oVE3NcELQFjnVx5TGJhHNazS/j89
lmVnqAKPSQRbXExMrFnIERIiaMLSSrKr7az3noeLa0R96HUvD7nE7B4e3UzEpOEe
ZCGRmR13Eh0m9LfMvBpUTt1MRMGn9KqwmYmwBsUXg4PWmv7F4FogIrIvoEgKadHw
RAenF1YyLDhTp7MY/UwzyzCdqTSh0D/gwFDzOJ3eWE/kyCAfEc3TYtKU0WV9C7Jc
fXs0wxr5HQ70+5YdQHUD2+2GfAcja5aEU7/2oaix7ls/dAIyb6MLiFiCxbOjkJ0W
HgUGyd5bvrFk2AtznLQKR756ITjPR6M/z9jk+AiPeY66R7byAtS/Re9p+PuKkRIt
aTO+SaGxrsVymKNVHBg+5DKifuYMhIXaV4AZa/EpMMRNKrLEsRSyz+goVrgBPHOd
FM0FQOYlPaTmoTKhsMyR1i0uDfXg17La0HU+QGVltfxHgTLx6CjKx80N3HXvflOK
RM+PfH0kPBG5U4SYrvPOrwd5mbeRWthfsg/TIxd3fJ/Jx66TJTqnMMfMH+wXKyGB
/QxsEquYY6q4amcFre5fBZvQDZfS1qd2mLiAxHQyPSyAk58eXyG0APdy0hacoPzl
BMI/tW4JPHFloyk8tHHhc3LyH9fOO3/rAgjJGuNV6DqUQpMrDobGKVSPoqoo2+v2
/FqCXKQL22bPdhX8ymSDJSsqm7vW5AOAHqWW+FWPro5qA+egpK3JgWHgo+cspCF4
dWiE6l0RZrU61cz9NHdGF51duc9rK/YyaWLnebjmjwJCOtbJ8M9Z8OUuDrH16aF7
bH/fMPMmMDTJQ4UDKfeHD2Bls09ZWNMHi5hIb6i5oHCqIY3XleC87vtnHxKMZDEG
61Ru1t8AABVo/+Yh0AJoM9fSusxOfmZyLU+A9IsVdzrMjWD1Ul6NjtyqxETKOILy
ClTdq84mMu2NY8LCa5ePSQkGkR7FcmyOy/mdcWE731CudT4sjl6wHHcfnSbh6CQE
L1O5WKeMjI/w736hPSQRbxi0I0jozoCicfMxTKSV/X6/HfddREW3U/G5X0ul2pMG
e2pNG2g7FgHm5kyvI7UF89rSHl/HKWuThHzVV6XzAmFCvJuHhhakO16AEjyH+eHS
BCxCE2a5tW/dqkygsa3xiaSqEWOwZeLx+pCNox/adZM2VstOd5obhj8bv2oU8xVy
74BpOXQXfykPvLVxBROs5UAbjoWeu1hKGYlA0z1PTbqKSbxhtmW7bAxDaQZhlduR
/AxTTXez2V7iShWYwIKasDCjVIAl2rpwK3WxgEgHNyjZ2mh6bfCrCJFfURwTHtnA
UFO8/h5ZjnzEo/0zkG+Dmym97058Zdm+72otIKJUoZf2xCn0ctUO8ftyfuOlFAGR
J5KiSsiBe+0SjGajXt2e1CtXlVNw0cHOoA8e99vB73f2lrUPoFuztKEB4eSGsF98
sP/oeHF2jNR0M28JwpI6MnSM8qo3m5bXuCrByvLyIajuodm+LFTRxM9O4ND73MDC
EFKO3QoDzqkS7XT7jXuOg02kv1vXvm5J98HGh0YW8sqfkqjHe9ELnftwx+afTwYv
hsa+qefciOvw4gCFriB8SMVM9Q17cNiyf2XQMC/uOfsLGjGumbLsVgiKgnIiLwJ7
jHJez8O5xQwNqlqiwRI3liiZPU2Bqgk4MQEmgp/9C5Wpz6fKV0Mjf3IPMuA/cpCl
1RXKy4+e4KStYgJusoj887GbJs5phvBrubLOOkAsX3EGvD5MEoTSyEAHwwLn+fmi
PNl0qCSvTk4vT7to3oItwvy93wIgPBbawdNCuuioQq6wwvuDxYL1a3cniqm3HXEl
ISBXJCgH1SScuA92OIiMxjzSDAEAKjSJwtS5ejkg20xCHH5fp58WI/c6d4BiHOY1
ptRbHRBgnmk6UeXMuv1CkbCFXNEOc+Osr0/6wYmYvfBieJYy8+GkRVzXhkDlxW7r
iunq0I+ALDRd0IB3K/DxsUFMcQSQVzxy3zAhc974qRbHnpx1QFOI1L07IOk0h6N6
Fi7q3Tnoxx5KWC2bUr7hxlbrwpgRlW5kDXNPEtvMmqJ7/ATwCQHos+4LOSlSvgeT
eaIXxdLoBsIM03FumDJO+EBpn51iRrrbcKTl2jPnYfYpUnpi4KvPZxLwD3+cLzR0
gbntYJUuMK6ESw2NwCcSJA9bYfltcGAnLzo0b24tSZ7/Z4i/Lp8zGL8DiibOVnNw
bRCd4gqMnD7Zuqg6z88n/6FGpTDOZvywL2hzmiQ6MAYwMbi3wkGPgEputixqFtyr
EJsV5dEo1ryi63ps1Q2SjNKuh8PhFVl0EhmMe1aQUqv8RHdkBUBmwNHvrzxZmHaN
LVCPh+xU4ydpx3Guo3CHEXZbMqbk47SmT/hViMOUN8HEXGQc66IwTH+wdFx1ly0A
tZBh6L5d94McrB2FJDcvXXw1Q0029xZZzeQbvZfWUogmuaOqR3SuSym0HbwLk6lF
sgM7x5sNG0bGjc9Y0mkI/JUoDRC8i5GNu2XnlSLTE0WcCtyZkCCkMGN/YMzotx+o
mhtFz2RK0o3BnwuBUeuwh8fi42e3gqLERyRNHLnvyq3kC0ZnguITwtn9doA6T2H5
Y3rn/+8QLIqtsiT3mv/0UklYNtJWNrWWEEBqj9vXsC2ZSK9b8KBGao+1FOeThdcl
bFiyTVEQgdUTHW8TLrm9TdQLguDny9RvWA5cXg3R8mR4kZ7PwNTFAEDgys9juObj
KfDIw/3kynjmrRTuZrJEJEIDf6dir92eHB4AIGVtFVQK46r5KMf0L4yf6GOc8jFh
wum80WmLg1bSpKA/GSpRGUdrie3q2gE+ySRTgQ3RrbMhKGyMvyW2F/Jq5PySSPTq
fOUQXbjNGXZ8RqYEHpvJ1VBxifE6pZD+RhMiz5TcDjrnKOBysdXdbffk6c2AVwds
bKvkPHHls9DWcNvdjtM5ySn6MlUh9jhgFz2CKUNF89vjjDLyYiLxGhiFzPBR/eoD
v63Tqnsduqs8Hx3owlD/m2LW2p3dbPZQ69TeMSrLmn16+xd7C0HsgSIX555Wnoc0
Qxa7V+07KoncA1MSZZsnsqPqVHbyT/4uX6jrXt7xzQARzColuLALwAIMSjR+TgeZ
FwBT5HQOexDZERjFUwNAsXNBr8vHXXBuupybAWRo1q6NMmfsAaEbRvHowtReUxuw
e86KUIgvboXvq3AiCHmMoJnM2qmH5zNiRcNOCRB0UMhDAXpfASEO9h14ial9jRlv
jmDMSM6cMg+Xn36om1AzUzqNkUuPw6ExtdjxgqJY7YnMPeHDPgz1VadXI4mHWQPB
GYI+4PPjmictOwoh2nHRr6ddIPSnhmVHkDjSj7ZOyQwxPWbz3KEASMwZOXqq3SkN
ynYIuxUA26YFPnVed4bGE56Lm14LaJNpD80KnHvJqmDjeKnIwlbaeR9SQVQpIDh9
xjKXwo91i7JbURJdsqY1MknKnaleUlXEPp6TTm7cv0fFiRfO2GnKFwqGevMRMzvQ
vtJdMCDxula0x3XH3zwBRa6/sJ8xQz4lBCWDqthwh3NzQqFaVmcXX+VzT6LQcnYP
JWNRi1wJlkHJbiX4sBYBKVTx65qg6i/6BSY/SW/b5LJz6EqNaAesT2Nt/mmDnK+s
0nFWvJrNDFBQyhmDw74ka04hx/ibldAxWhC6DvPW2sOv9qTTJ0GCMq8ztkbIULl2
DDKq5cuWN6fYUIUUHjM/A5+ZrFW4d5Vc6hFe0+CdrWs62WKnDTUHDOsvXCQefXgN
SjinCJRnv5i9G6YCkLSWWtZx7eh4VGxgHZVvLPm3mAtAf5uigRQSLduAPUsPEP7F
77gsbxqAnfR4q5dbl3iHEyHsgrSW0vjSjy2bJyBCHvperE87WwhckXbrK14BT8/c
8/tbI58RnmON4v4tAA1YF8G++ISkFA9sg2aSRVNUq97W3h38mt/G07yCwt4peohZ
H+yKKN3TIsgd1MgPYAOAURCm3WY6Xg0zmumtfOjVfQoXbgI0Cyh5FDZgMa+pzNiq
fOeQ4nN+bQ/NsefMRq+QVW3ZEqm/LN+t8sTOW3kpWqbZ0aGG5AiwsDReSc7XnTLy
/7eDmQXxgd9BHG4/YjD8pMRQcS2GjvJeQZ7UORqfxIWelREOM1ErmEFEIzRgdM3O
9gunYwIXCTwMMNUuMj1ZVN5grWTJWeHISZNjPx+8swHiXwZq5Bx+KJM2Zp2SaPR4
vW9fCNhdLkYRaEh4rmwE1s1uX+CR20voCHlH7uaPeTHwkd6m5tdp+wfFQNieJWMW
/4xrHdu8wSTE67GS8eMk9KY/8+ymcTnVfwm4xYeFd7sL3O+vSh2ZMDTS30YyIlQf
bEuWpWg1dBdJ565jFVGtekn4s2aUHcUH33L14/Vm0ysE4POeCXheOe0Dkn9FNpqp
JZDpeo9YYO/xnPxsPt4+Zuw2xaaoTDlDfaCVbdphQOR8Dk3BmBTOLdl6ZpVowJLR
8K0puqzUH0GFwlSZ4RXfjlwdpWjI9T9FJjUqLeCjkZwyy+bdlgbV6DNsLabdh8lB
rHvv67jphbfXqhCxPTBLyoCoAIMvds3JdLSWV1IfglEMAqECDKpyjzLRohESRxPs
kYGzIA0uRAx9d2xcOKF13oV0nsi6R37tHXVi7WUlbT+6fhGHZgOf2KMuEbEKwsm+
HtwaDmBlY8L+Wp2h169W7iDSfws3ZfrZbWzWHWyV6T+OJIRjNjHvBVZh6uVvlCf8
jhUtEY39YdTuCAJnzLB2kGbszgx/Ura/A22AlOjjqpBHYIQeRfaiW226TLPlIG+7
dLhZ91riBUZtZUhW9F0SPszxYsO7/1X0G/9X2Sn0KJ0r+Vui0zRY8LNXBFOMfhmh
vzrq5UzueQr3hC1wTo/kxUcrSJpihfO0BJme/K344G+jJsWPKlNLNPLdIYjEA96R
ewteQOX4SyUwRHTQcXStREYVaKN7Lsj/yrEEWowWq2168Qa56z0qC3qALzGySu5P
6ssaX/76YklP/D4HqdCTW5NvmjGuWWgGV6nDh2SUOwriVBeJlc1j4evR3Mo0lIgq
uIYJLy7bZ2JUs6X+L46snpKYN1IMMlAg2Sl6wpHBSPBg84eI90I7VbyQj5rbn3ti
ahgNG/JvO+dyPvU/YhAcdzlPEjXWIKoFPRvHCExvDQuLDKXnjnqMV/nPXg/nAhS4
mjb56yU/1hvKNvReFM+z4mwF0nct+tWHcZVxq1lmX1hZSMAoGQkqhafdY0yLLARw
aA2z7w0mxxkbMikdCxNxKCZZRWDD5sy4YENcv2hZ+HmqfDmm0hvuSAqIOjP0LZhf
HqTzlxQKTAPqZqxryjJr08dZqvWvzGAVUXb2k8ZocfWR9HDKvuqP7O2utVYM1AaV
8fDdGzPcTPN0mQewbQxMsjvMeToYOUGhMaz0QDjEpFR1OcP7MNAvK+vCdBtkn34a
aDT/865vpZU9jB0nONCJLmdiKANlrY+z5Y52unTJFsoNr9IgpetUTp9V878IY1w+
LX+4X8nUMNPX57WNFJ96o4gd7alr9EaQLujLowgG6Ka4aScSkplFkkNCAKtoO2/w
T0F/M11UK/o1gfDgXC00ukket5Kdakx1SVXb7iepsJnexDgSF+tHe/M1pCe1cvf5
Vr9KH4o0is8vE9kCjsD3l4bKvH2ErSt2cN05IiQfJ6Mn5pOyZByDWlJsSwQo9IcU
5dVU4Twn5oNQ2VqdWRiOjRBGTWIwduhzTF7joJ9QK8puGwKSPJVgQLd4rpz+Mqgs
/Ix3WqJuMHErBnLjBkKFpb3PWWoOM8q60JpKInnK4WG/lJZcJQS0nyxr0FejBWTc
ZuihjSJJWGb84X5QeeYWJErdN01qXOrlQQO4a5QG4r8pjJSk5qU9+1WPsUuQkgKE
u4ag6KxXagHyBq++3sN0FwMUGqO3m36FwndixFnW/ue9SdbhF/Lyy1a/JWc745gZ
tNwTcVVQkWrto8kf6SQmzGWH7mozJNqppegHINkurD48XtM+gbo9/SdSVcaWGUob
HUyEmoW8Skr/tuv4QnV60P/I+DOjtggA21AI0HjL9ooYZKGa9rNBBtgG9Ezx+ZQe
t59csrGP259OIYHXEnKCb4k/6rlz37qgUk/EGQ0oUh9SbXETBBrVx/na3B4tZSTj
seGifGY63xlnstv1QUXw9SFLamerx92XnNverZ3jQxJAoR7wq3xEuBERXJ9rfk6k
JPrSpJ3PU7wPCVtppsrevqMzlFXrSoZQOxEd0yJiZ3HVHxny6QffqGpezy6qJGGC
ZLcZOfUMr3/kjcHvFXyHoR0ee0irLH/t5QldE0XugcnnHjgnbN0ZM4pIbeMVou71
SyoMl824jOeKm+UGbWSlAI2YPbaxeUbAZ80anouKsA8FGSWXwlcKePU2YIgd3fgC
Cg0DC05p8B2mSxXzDpvx5sR+QgUOldRefVyZr7jTK53tB4JBwkkn9dHO/r+0IqyY
10v8VpnVsNZTSxSJRx9XwMNHJNecbb/Dw/h//9TYeQKok/UA6hGfCEQRqWSL6yCb
daXr2JDRpLtNN/5BJoN7waMLPkN9TdHlXXu2bd9DvNuFnfVZGP/zrq8XMoTf40Kf
jSxE92bTnD1AMbgOTkRvu6HQ73dyV+rCo6FV7mRMXvCwlrECfuLiPi8QFv9W6frN
aQXgySMybRfz1rA4GgcLk/pxbQVubhcNQlIsuPMY/ydDfto2irXXV7gxtY0FGaxa
zEdKmY3qsu2Hvx/2jCGnfrIL/wVs0Vj7P8ivhI1doSWp/S8zhNHt6sNH1/0FNEZS
xNcR1NlVk6qKHFk/YDSKkmZj7fxDnS82O8IwE47JeEHDeEEOdxxarjaQ1Ii9PovM
rdvtZbQh7MJbgd3AAAhNnYq8UAz/fgnyze6mwf6I0IPxC8/cEB4xSiCkmJ8QhJ9D
Pq5Oc0YKKcCd72FbN0AXSaqL9T0MKytnFdZj/wH6EbCWxEfcBNDzuIftd00y/tYQ
SLhGlOTA9UHsRkqyfhJgEThsj/LTkSJrVAwdsl5FNemA8e25l2EMBf/qFOYPMoty
/KExLnu0WYBeOM5ECymhgcR/zqaeYLUK9c2oCixZZhy25fp8eDcvcMf189MHtdKZ
rxVptvKkt1wAsadJQ63gUJPVfvAXROtg7Fcxc9tPp+Mi/yT15t+78ZLs4GSS4ILj
FCRVcDozG+dqpZ5v9Q1VGOiDYf1T+eQoEuMJwjABmcYJbEPhNPV8Ecec28vVw7we
XabMT5v/dP8nCD1qXdlYIF1AlHPI/WJXtC1AQguLPqARrB5D8fHaEIwoFV0BomPH
Z4qUByQlJulthzImi0uejMZWpAhkhhVMaPu83GD43wREJrvbo98Rh7ySoaGM1IuZ
18n1JkrGxd+K3LL7G2XBBhAx3QaT8lkx127uiW5h3t1YvAe5kr0e/sfdfXxLrrRZ
mxGb5r/4x5tAUYG9dBqpE/bTtI/cxvNz3NudyAUIw7BAPB78XeBG85FpxWapDNQ2
MewSQ1/tvj7kijUV8T7iTxPIRCSWwrT5dXSezXd6vVXY1f6gfBjY2Xi4r73R55jU
zfVDHRxKNWfYOVkCJwtQ6czVRmtPR5e+USOmeJgtN403R111eAy51fUXnVFamZXc
opws57xwo780YGXehBiRnJ2tP4j0LB+iMfbbsPSYiuOk4VHz0hqum7E0Xk2XbB6g
rSYPG8hwYp+3h8S60+bf4a461giZwPDkpEKcWWAg9scL6e7COgB7xzgU1b/7kG1C
t/5vcqU5ss6S12cGOlEplnhyaQsGk0HLHac19ZJCoiHpjoqk40UT2WU1omDDDry3
ZUYRPPXIhTrPvVFSjPOBkRoetxmE8bTlfPhDMhK+JWtqj1XDFAANTSlwE/1chOJA
2OuJmm+BL6D/wJs5QKt2Q1iyVOZMXmhk9KygBya7N99hzqu+uRj5fas08JZzi4A4
L9WMsCxEngg17wOgYYtIubbOrh3T8hjyKRYzQghkmi+61MK3x37W2VCRWeXMoMii
SgtfCK0tziZu8C5kBXkOA4IP4+Rs+yCqrdDi2qwl9YaBdydhLa88cufRE+E5U5S9
rVjzLChZNpChRJP/4JVB9Bi2T/mVWw+cX/XiJjier4q4hyXEof9gWQieNjEUCVPW
tv6BAtFYw8JZKnxdxOi1/nNdppz3rQtklzj107/PekuBSHGpNfUFUqYZ/UGFlKnz
+ivRcIlswHOumZ2hcvAkQ6KnSmscNcn0C7Y6JQh0bRrzpNijtWwyJgUTmGv8S1q9
tXyLAcz2QGZ7ok8U52f9kOMw/kLy0Hgq6SOnG2p0YqMUcI8NY2MXqMooDfIIjf8r
/7TmHEISJ+oCE2rKAab1KwiiAIyM5RmarXn1b1nOuBOyYsXJ61AoydijTCXR8upH
kkjajAL8l9Pu2vHe84nDZxwFayZPivNzqXkPT9XWFeMEdk1uPUj5hgUEEaubIOfd
ldEOcmsNq+786AI2IS14O++HucYxj6PohHg/nWQgs7o8NBHWq5JpJF83rbVEz04w
DXhgKMrze6qREH/RKrxZSDFLMWLNTo7xjQW/4Y30RkooNJt1XUE8vqLHiX+Nj2cA
ogHmZNifNS7FshGm89lcFfREgr3CnYZJzL/2xQRNQKUcRCrND3iUiYuqBw9NHChv
yUROvl9+3Dzu+Ox9bKIjVHSJuBKYfqALYIFB1m8HsHQovhmXeVkB5hb84GCuTjoN
n/EcKMRz6qkWoTxyGwf9gbzj/SDq+hbMzxAFNhT0fiQTC1V2SiA1DDntuqIi37X5
C0UsTHp1gGox4cpTsBTOi2fhabyI3gxqX9+5nLAe4eD1Fx/cmE5FzM8aSkzzNJJo
96kEYnaMJ9vz3rytcQyC1BN+jEQBHpQNMVtmJTmuYjzAXRjaK2KRngGQ2SEA6NnJ
T3DPARVOb0B1714gE1bp6mLk/J4B4u8eGklDfdP/gX/a0EvkjD2dLmTywtRAlUUV
yFsy5kCdf22Jpou9lbnmiJL5K9LHJecU5/mPf8YSYh6+3ia1mEfXpk1XmXULP+zh
iin/KEJUfibxHo5r4JpJlPf8BCIeLnCEQVdwQMkrjtpkk+4RX8CcdBBaN/OAgbPw
/aEXCM7Hlfuvg2yAN50URB0j5VbIsMDb+QJOL6/ceBDWWRmWO55CgmKDHLjo3zdI
P8R5QLD3Wxdoud6iI4s33G7/lPZwR/OD5or1KiAiM5WsIRkgdqa2gnUbFJ3h5dT/
Ahnnx88thugOCCx8qTbha+ht9ITnrnS8gpzn2XSUki10hWShic6C9YYymeKZB2SD
XeqF1+cm7isgQIeR3o4l76kfa8ugJkt6KJM7l25NAYK4kpt9Di4UDI+LChzrpYQc
pvdwajO/qtkuV8C3ZPDHNpKZPV/bBUZNi+WfJd6Jx1I/E3MR2Cf4D7E7fZHLC22d
/PTmnxqYMxlCcBmvZjS0YPsAiH38Yo+l3BniupFdwpnfF/PqZ92kQB8pg+QEDtSk
oEO0zK5XntuVbMiwpkQ3uXMa5eayDo2Oid8q/xa+O+f+aFxT8ISZdAe1zKGA7oqo
EpqOaBvwkon7vhQv+ClwJ+wSflGHo6sdKzHWGvJD/8aUmXUayn9cLbLXTeR2FmFD
bEE+SJYX9HlZWe1AaPnyUEMgHuI++EkMr5YMtIduJ+3PmYvW97t1rpfLj9jqH4gv
zB+tFE5eeSGSnBPwt/imHYJuxu4n04IDYO/7lkWNhLky8CV4CIULf4bIZXHXdmZC
PzdjzWCcMTveTFJG4kSvUB7UMCFyIHUatxRZ1nR/MWpqlSU2mDMEBK8yD4o6A7w1
uP7XJulF0PVU0AUxJgqYgq5dwYX9LPQEk6OLNMKIw5LBGflrcjSVOTWZY839WjT4
d3CoCsd2P8ckgCSlPA82Z5GIn0vPt6Q6kWG7ZQPnetX1LVLg5RhKCceSv4zTdm5o
2mprHWMAHxepj4iw6KUdCmQNxKJUAwPLMJrHc7EwCVHukLv9vFEI7bNurd4bi0Wv
uCSPYuQh6TPKOVSPIhd5fdep1UFrCDW2oMsqjTdFWLDGTAo5iyKPqe08SCPkIjCU
BcU4sfSrCMl569A3NQNYt9y0BhlALwjo7HfkmHhUf5SQgRkmwDp947qDkbmzXYzJ
f/NKdehz6GflbtOGdmKZ8fu+itETbD8oWBbg2/H/djvOb7EpexGMt0rG5hYRnnvi
zTdLHh2uSFy/Vt4kj8nV+h5ZoAGIyv7tSpJ0rhmO7gpRfJToSEt0O8TlC+PdXjb6
f6nTPEUREquRh2cMfav1JxJU1H7B0OmD8RT1Ukbx9Y2aa1fhJTKAa6WX5vlPLw9s
tleGBrfEDgKgW5ymNChYGxdHAzFPWCLO0bYRV9+EGOxPfqi0an0n1/veCUbyp7xy
HkvWvQtYu0/bMyJluan/6m2GvYsDL04JFUZbfVv00qiGDUN2FqOb5K0SDnQwMb46
m2TISjPF3FVKvGxZSgnE9BQi4tM4/pW85h4TK7woNw5RpP+m3/tN800TtyD2k/9x
smyOa6nBI2oH2WCJYo5c0HGV5Iv8ZaHUTncCVCnzim9e5dVm0MhsuPF0ohqZ3rRA
GSkgGqwfdQ/I+JFqFtnEe1Gk6nxzhydPi4Fn9TUtYlABOxrQ/MycSK01WQ75pqMs
g+I5D3JKqcV19/0dQPIijEU2MFSPHriPAVqhn/FBtPVikD+lZxLZwu9fbVNxyiTf
ZBp6D/c2OMEyPZSR/0Wel1XmMbRy+QEYfbJDxqpFagK1o8yRRoT47W49C5DGmPbS
p8IJcYZoi5ZTpMJHLOiV+QkOg1ngUcT06Rz3K7tD8DHCKBJ7QuafkGMEbnsK+anK
H1thUx/FEgLBwVA1EDCtUnSZMlZj4w7Y7iVLlC96sahYiKPEqy0dP7f9YSxRcC5n
/ok6ifGO9n45SGSxu2bFqEc0Hr8EeYzqKA9ULRjlh/+4RdzHckuONloWke+70v0c
Tyv7+yHbGB2J4gV9irDbKZLwGV5IFNYSCg7yz60V4YQoL+QCjSSv9r2y4SlTbgPH
/mKJ7/vfFoa8/VI+xO2qr9Zv4GJ110GXO1/jY8Jg0Qsf3NorMXJVCeYUsBWeJg6v
fpF0AtksMaHETvoSjdsGUEpWEqYHoSIBlpRzlb0rfUYkkh61ehrO+goRpW5vMKgK
Y53otzt3Ho6m/QTvmRGV5x5YQIyqehsG5H+pmOqLEmtEBVgYRdbUGNxbs4c3xMZo
8LfnFIQVyS5PV/Lrvibxp/u2Nh45K7INN2phTenbRoeyNa4wpuYU65BydglK83+o
dnakkPXAhl7bYKYwAPs6OhP6C6DRk5PfdY+y1PqNGQ/uyn4uKbc0z8ftyGaRSygt
v8MJ6gBKc+z4s90b0AcDrBUzTh98JHLaOsFviwIlRca1B2epHcHUyk9tRqyuU5kj
68zlpTATYnJYRvEXCj++TnxOqIaLHEJDCCT7MviJWKrMVYCZ3LFu3zNYhPEOVEM8
dfLhaWIS0dWoJtd1LoU5gwJm9CUEKnQ9WbiwM+l+RBKZ/3XGqGUAx/PgASl7sJtA
6+nWQ96IHIjC749DCV3P1yaxaXl67iJ3Ox2680ZNLfHvoXlGcrQvruD4BKVz8Wd4
/W+7oLEyJs0qD741oF5jjGKYmr5W0slpV6tm5zDcbLhBZR1TztiLwpPT9Zn+yCLb
evlRalqve8GMt6vTh/AaJcEVXW0shBKk24ZsY6M0x8HwYQNE51iEuf+XT1CHlAcs
ylpY/5fyn/xZrqJrlk7AKSUSfWqBORAPYA11cV0hrykr69CY1jrTePgX/4tfEXsI
UfDNPscmFhvx27fdCuzZU3hJimR85ujzssFCh4l0SRuviooKYOXgsh6mf/YiAPBm
gs2pdFyqgmlrDoRh9Y1TY+cQguarC9wBOuzLP4pdhk9dqs6ws5nvABU0ijlvvgTg
nSANBCZQriegC0Ri/KaZxOBhgYc20/1VPYi7ub/pSY3kru9VaneJERNKQA3nYM0u
hJQ2ZPGvFYu83x13oIQoIfqMoNgMIVyOTmzutmS4heWdjceBK/M5fD9OYTRyARB4
oIbTFgNwAMzdeEniKVWLWUsq4YkPEJR0MhFMHIyHXQVaakIjZ9biGVow0CEWuSSd
Rt6Ie7c3qAY1eW0D64QflBbegcrgizN0ogEKse1RIKsGbXUQvwlhE3X+OO1ClcuX
vamOIsHJ+RSWCaLSTNFPpEw6CyHT7EkL9n5Wj/7tHRhpb3+fKKvXCYoNB8dEGrMt
Fuu7038JhC8LnFOXOgZH+Gw5QhUSsor3sDT9UyM/hwG03yRppDRcgsH17gsxQ12X
Wm1YHC45mcpI0tLCIT9PACND9dCQkuRqzxbpFO+YKQzTOML0njFCTMu9LFW9NDo6
9a75ckpWPYNZ4w0u5sO0sjT3TndovlcttvU7Hg28SKm6DUXvIXyi2i+KsAQenrKw
ZW9mFZ9Ei2KCds2yQQL9OElpTD62zvuds0IYE0krnJ47k92awkVRmMK0Oat9/Ot9
xtiGeb1xV+NXTOhm+TbGTWuUVvtwgzH9W96GDPKvYxHGQjfJYE9Wv3HS5Um3+E7Z
ZschO0v5Fsnn38BkUUm6OWMYPjv6LRJsbt4g5YQjxA97q+bvt968xF8X/JnHSu7q
6zEchHqOG3OZCQoC9AfAkb8fNZTEHlRFjPkAJoVErnuVIURc8pXqbgNP6lQMWqlB
yIpw9kSegjQmTufte70ZNTAx8FfaNDYqeV8Fvq9jtGXrAm23wsnPgDOYFaydnwF/
qo/ZH/8kZzl5mLkoh5bc27gutgdrR5M3806VPfiPblBt5eZyubWQF68jn3w4r0KO
VZ/LpBN7HYFsO2VLeUZxT31Uxpzcf87JHMY76nu5aB3AFajm9lzL0eEoKb0NyqHz
XE4GReA4Kw2VMnl5X9P5VEki6rB4CcIJERZSFLC9a/yGeBq1unCpHlaa4+kFP0xN
bAjr9VoxgJdnEzz4LJY4o2r0rU5ENJuBXGWwxBg0uRO0eod+OJ+Qu1ufukmas7nQ
LbSV0H3WUd43FIUfswl8r42EVJYTT3bHU0kd7vCdbsIcJs+i4iy7XlsLOiYVduwT
oMnv3Zsr8jFg6XgbQ51VYdJnrMJP7VpoHlTEVfNaGT5KNxQtyLBnFtJRz2FAgvX+
LcyyRcofnbNJL3NQe0lZWfdMTGXEoBbna3UTvAbbBIga4wZADFuRjtvK4A7xU8pJ
rcHkqKJWKMYUl+NorLxnIDKXgxk5lGb07uMxg3CpkbRvTguyp++TwjgwChBaPC+B
fs6ZOBXYyIBFCdmGbVHHa+K3LrZUhmXpBuHNMgeb8xwPB3V11U4HSkXpkZ8eLZrD
FfWOVcqzsX2corNx7Eep1wnteFu9hN7y2LdNZEyrCf7cgHj+EOiMnn+TqHRVlSsS
EFwcxY4yThON4+n2HgREgGJ3vSIbX1aZZGuKDFUNKYs4y2Fvt1nfN/lcA6Cv4jJL
0W7pCyJHQ4dipBClHgQnGP/TvRVUJyf0KR0MRBbDzWy+fDWAEFUU3hAIvPb1JmEb
yuYDLqpbL8woW5+6A84GixNJKUCyQcgR/rq/HAq15R4PIogX26olFnyQ9LspMP1B
bS6RDuuO7+qsQmIw2KxzglUDatzkwKJWopYjNKy+Cr5J2ImDpQHgwHCXlRK2gJQ1
S0bz6G5mEcRp2gWL2v3PqOiLHIImFuW1+f6wiprgr1n4nxWbuVTrENEXVxzyxNFQ
o8zWc1+xKoppQNyPjJf1tqAH+8x20u6U60VY8jflV91LjqhXrNjWdaxvTFgwE1vI
QwgYm7qc4TqLZZMjyzXSUh2KqTRreSpEZ+qp5CqKpThc0qcI4UZ+cmLJX9oUbdio
0IQQJzhgHA2gosmhxkhyuSsEAWRL7B7G6rO/QaDMFa1uiYyWC/ROgwpDTnLJ7Cwr
n6I1WYVDfQ7DfRgrsWfdm+bqnCb+/7ir64dz+r/XhPWAiTEinUBE25vMl4a2TWBC
yYGxswJP4WECxCe3/DMYxE3nF7M0xE24K9SK7cvyVNp/Ov80x0FBP54gHWOFPto0
fU9Vd8CRCJifCQ4eI5vrNUhSKQCmK2QFcMiHCrDCLuv66lGVCk3ld/Ggxx6DRpjN
JkN3YLeU1UokJH34qKYZQPTWZpd32poA4p9oRSJXapY9K1yPe9//Mh3cci8KvC/y
Plv4lpmJ09i2R8Ane7geju6bSmxUUWVMStQ2spczl618CFOdFvtqZOYNDqbuDz8K
q5A1lvMsl3IMDZ7FQmfWzQbf3ZPugSr0jAW5OvIMvAq5EQehkHflow3aCbgse5G2
mJs+J/7s3tBcEF1FqRjnkhNPyshT5DoWU9Mi8WiaGk71BZt+xIfQambTAD2DSqJQ
gjuQoVkYdEmsdMJQJmC7Zu2uM4GYAPjc0oWtvftEqNbb+uqCtqMU0u6/oJCvJoU0
n8nVkmKxbmqiLTxUThanvAc5Ku6NOL7y0A+xPskCFT5ScdFa2Y+oiMriTFdo03po
AMJ5Hcm4xz8RXd0+Hsw2lpOoV11Fl7z8dTHh+PbEPFF9hYbW0gXQvPSR+Z3SHneQ
cI8YQHqdN7HOEv07fI3Tceytp253f/a4qtakjjFDM1YwPrrZN+xWE0xYxYlx/Zt2
GACF7Np0T53i6OjPT0+k2UvhGWCNVlFegzrMfxfUdrWlIwdQ8j3WICfUR9l49JXD
ANHvSckeZDXDTaUgA9k5E7XGL/+VR5MCB/8Db5jTU9lxU8ezc62+zUtG5pdtUQAs
ibMtbSlZn3xSpZXeMwCVUyJPpl7wUTklYS0mhGg4FXY1b+MnfFYQH8e5iBHBtoa9
/CSfr6wH6ZG1mZ6SoFPxx3DBD0ZHas8tontlGxoAVjL+AKcUYGwwhBeyxSRhU9QD
IPMJz2gmwcIwQL+TobHO/IQVqyqS0qxv4i1Eok3kawvEpW9oJKwenNUSRkYWqX/A
airIlgk4aI9tejyr5jXNHVGa0cdP4YyspC0PNbieomiccKelHWxLxAskuBc3CgyH
vcQvebQ3aMvEQenUXjSA1f1/At8uwY+RF3w2elY6rTq5+rDk+tPNvplVrHvt1Vg2
GuVRZwRKGwLHnJJ7slfMPi+28J7aK8BHr+MV5UJaWtMdr1WyvZ35iwBlEFsyZcJA
ND8lpcZBm4ZOgOT6Oh4e+G/jB4Ncx6+qZEf/CrFtFIX5I6WBKfbm4/N51KvRXLkw
eX55spg9+aaG/Fl/5P2InZmsE48htl4P+61QOduT1Sl9/kLdrW80el54ii8EjMWm
E98B1MmiZ83F7kB6tYn4Md+Mmyv/zXaRsZg/R9RWKw3lHiYhvVtEFBFYpuHnegF9
qZ5sPrvlukFZwpgvT9O2Jcb4FEZXDKSgxjc1vJGbyQPuaH0oBzeqrGth+PqXSeIL
QCe+3KCaXSWVDuxJXq0OWA279TXbrkES0ZRUzX2iCx6ogUWmvJluX1SJqE2aXmcg
bQWcvuUCrR2a+B4dkn4pAX1w1gJKIZY80Ww6MfN+D0pSBz6/7TnXcOB8HAaTbv8M
XX40TYOL3pOwyFLnzRa+FZhrTYnqWLA7saFwcBZO+22IdUlmBbWw7a2UG5IP4uEd
5MMVe78p6jFMPur/C7nqvLeR/JfqEw/YA6TVMS8jxw26RtLA0PEWsffij4dZ1/op
54MK87Ut0YKomncCacuh6FdEmop0JVYGJI/iVXy5vNW8Ap5HTx0qSk3IRSbjpERt
vCtL0NQ7ngh5gHzq2Y/oZTOh8sz60ozFnWjhisihcYhDtE3GLEF/NiEJhmI9Ktf5
41NQk5gJnFn8Knt7dhhC9d8f67KOiugr4FL0DhMTiTtTRGaA5RXfyaInan1HV1Ni
iGZ03D/S1hn5rOIJRC+fKd+uSc1g/AO81D3y5d+lxXALCNREg6js1Rn0pU5pxjEl
+rmUlb2FpLYM+tzXhADs7qjM0cNqgqvvE1+hMeGBaVtEXl115HQoL59oCM+uj1nl
gPvq67wrZ4Vfe/wIIntmu9b6DSXvufcBpE2xd2sJkwLoGRCiYiSjJEtPNyeMP+rA
bwagwp7mp2ZIfIcAh8bPUTxOYTeP92sMUfaYEFkOMnQtfdKWicN6rMHZzt/FOoBn
vMz1ga3LV+CCF7KAVOOzD7HhmXikUAFaG/bXItM8mAxFPMoCFeVtJd5XgggP08J5
tDrOtJscNU3HsHWULyBlZnAJx65IQDVgaW53gkQY7jl5e4jYc0xDUxLwh7R63Npn
u+7Q8l/XrxQxjtBHUc3LWieqot1FQaGzD8K2Qthm7QHJ1r128sttwwGtDMNBIlGY
VQ3YuLkP2tv/ZzfGrZYKnB6ij6xXTJ4gZDxyPGHqVXvgayhU3mhVCMSDArmTEEv9
K1ZA0SRRobvKqJyRea4t8lTT5vZpKdYsuk4QYP6GdTGXtfQPv/L45fjwOYF23niX
wK5JfecIc3rNkzrclcEUgipdEiCcW8ba/7VN5fgVsdnyYKytE/+fbUPZ7ylLlyje
Z2mzTIdjNiActonBOqtTSHrZ9vCR9nCvRsyDqaYSpkBNT9/gpvQZrRu//Fv8tweR
2Z7cCSOlUJYICJZVOy3O73hnSrM6IUTJXK12R+HvRbgbbHby6A116qaftqJOVwxE
0rTIg1cTMLF1lvEBfRct3Kq+78qeSf7ybeZz5/oOi1byB2Lc563do3vCJi05TNNv
etUxdYmw6BwjWK1h0Ub7rbAQFH9E3E034ZSg1vFZf8bs5lg9ZqQV/6T9mF10Ppdi
h8cc2A6CfrRbdRy15G42YbJiMvH0Gem+YJQDiBXsDrAShGobm9pqUGjOC+ofqKaF
f0Mph+r1SJtKcaZurMoPiJIEXox4j7qewmsTqmaqmnVcrMET7n2B7B5JAciZ8oDE
W33H/71tjkPyvgVgwF/MCg4qMtdc8f9CcoWSKnquuHalI8r3sSnCC0wtuQhOyyAy
5cNCY8A1Cd/LX+Gs44BJBg==
`protect end_protected