`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36704 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
YKazAXTwZvVeXonKKI9l+wyioV3+AZWsapZxqCw1h+/K+KvI1JkJRM7ycMaiJ8Cr
X96ghURLJFwIHxr4wylS66Tx7uSkz50MPahbCaC+k7DDli7Moi4jxnsbZcUUtR/G
wtHD5OCStw1OR+9Of4pn8LBojxscv5DeA/UVHvvEPVcGIYcBlv0VfDamzaB7uYE9
RvZshfp11x0phtU05qqUdMYhTNj21e+Zta8CzXVcwi01LvkUbwRv6iLjEMwXYMfk
Q3aRfmyM/wwW08O2OihUMJr9NgdTdMGu3FO5i7bJJY+8ItCvq/MLNw448soCxGqJ
gJsaDdvSUchHAd5691z4lhrRxxBPqgyZLhk4gJ+8dOTLJG3gPtaNPcfSYBxV7Iqy
GT+CN4A2AU+6NLZw35yyCbbeuJ4CGPHqU72VoE9DwR/HCEM9bgAd1S/aEApJASFN
WqH9/vaTQPGLVThD4HbiL3JGFo9Tvc/QS9MbSdpfpbxlD2ust3alvzsPxURym8gC
W5waYZ5627drBvawrvZ4CXynFcaoiB4rHKeHi+y6RTzsvWL2Cv15j5kRas+1An75
eUPRS1g38gPEv1G+cbg4osa2AoY2FQZIYMcWa9sK4fXtKYGRckF4sgFey8pDfbol
s/6e8hPBs4HFk56n7P3rKLZ7tioRtczyvThI3TQRDWHMeJNv7/XzBc5HY6icrFRZ
/Y/kPTYGoaRL/RQxGilqA7toyF1m2UfMHCNHTCnwjys3kolosViAgDx0ReGzI8Wv
j9T0o6Y5BV0npdLMDYfNo6rtKnwq1sChRbFEqwaZfNVlVSwDuuCehXR03u+BLeKY
uQ5sduhBdeGGh8pLDZQLxk2why39pPBx66C3v2ztRu9gjWsq8kW68lDbOZrU/3VT
2S/Z5Fv/msnrxY52XeCp7OtWKL4n+GyDxttMUaae7+XXnoCzokETaE6XKB6GwKZI
by1hSC2dH1RYa3fTChA9Tkm/IVGO83WBHSa8ZCpt9lseps+fyg28yJ49lIL9rrWQ
XTGVKCAu/vVcQBke0XLasffGSqZYkV6bmfdSSp8KHz+rzlgAY/O7xuxhxlhzPo0G
SAi5z10MNQ7N2ca6mbjIygh3Pa9qP5yV0EO7BXwy5ToOJ5ADL4NAMFJcvSJffhSJ
pbhSZ1xM2HcTwu9x3lcSCjzgm9VrWSV43wyFikoOD2Gchozurjs026/LMMgs7hmR
Otabb6+1XFnFKpDEhK4ICbc4xJrAtKEYu3JTq34VesKiP2BGmQtYJzUepWWOGT7W
iu8jTDBOmYiaubeprGuME5I+moD7Y92IhyvRXurvD9SVL+348fCO/JBcrBd32UGH
LkdWMkDqDnXJOfPwWHEZDVdN6OKFDRMl/qR8cAQlJDLEFALM6f3R0N06plo+ngzW
m1YRJjzOF0fVAbQIXCC5ZEACveXuWARS3sTrJTzRcAh71QEgG+7vJhmVqoeaVv5e
yZIMxIGtn24lcbu0yMkZo4Q4zfgqcTNAh3XQbyQTlr1BULKkKKiNxnYi0WYS/TeG
+iEOfYHZlfv0HldVwGkn1GU/w+nGrtHCFBuvaSjeqcilDyogZg/wYDWTKYEuscK9
5PkpwOyS8Sbv0Tjb1b9c2kU7fCo4rTGZk/L7h7xKEoskZq/DE2IQ2wKzrLZdfXs/
8qJuWpFqG0KaiL2zhp9Frlmc/4u1rSBFaPw+9BgD9dfmOKMSrrEDHtkDQchDk6mL
t2VCce6wBd/wa4x/mcx7aHFvT0RMKzTkjkQTq6Ad+noZFcen+Aq0g+PkIcgxH/Lb
Hm/kpMbA7l+lglaLb2dxCwlBvJe/iMyxVtfgA6w2xxbYfNhDO9Wo06euBybCiMr+
2wmGyIF5wWjMgZM1jdFORW8w0sz7WL/o0QQPiO0fCtAu5a2n/RyIbUtZrJccSMUs
ruKihuaTq9zMhws3KGXrxzLSidpL7v8btnuin3FLM8PZll/GRulCMpDYXIjlKuw9
1Mw7cGuCGq3fy/aBBOuhuZBRJ23FAHYtTdh5iaVpxDlY328eAdStKlrIyZGRTPAT
RExhK26E7Q8wGWmHRtO0Ih9pKbkLvA9zTc7F2QCP79SjgKhbFDWHUKxuzyHVq0KH
vcDhR/t0ougFuapobP5ZMfheLSy+j8SC5TN4boJ9zCQSS8pgpd/uDMkAoPZmi5Tu
xY24Saz+MlPuE1ezQrn1cPwT8jVgJnUkhCp5LWiUf0Syyl7ujAdor9U39f+9owVA
TUGyeGxGhNQF5o/lQMheEuVvVfTjLRyl8mP2JSw/miuBW9xCf2/af8SZdSHACvfU
nNFsOUdaE+wElkd74ngTWHdio80LvUwPdOM5EtILcrtZAy4rkhjR26cJ2n+TtLLH
hiVyVfmfWEbE06IcO7vzr3tsVw23zckUDe31AG1HGf+vqXQe8RI8fx+S6AkcJVaI
fEgnxvF6BmMUIYUP6jIL9I+gmb+nAHIC9V/PHOEmGGftLTr72WwmU1Kf0c3CtqJb
J/9RqKbjxMfoyM34itHmp+KWwKPlfkZM/X7bZbbIy8JKfqKcqNzXOfTPIqlbBlJS
P/pE8yB0EYGXY5nqhjXJU+0vDFTueC4wYWxpwkEgp4R+6/gmjEea09u4DR7UnMFs
enGTyuxaPYdc9YcPtby7z4tLPKjquiayiK59Sx7K7QkTmJII5ZOnj4upr+WI0ksQ
esQZJo5U4W0/mYTA+JrSMtoSKJqj0wIX7biqnxFRzBeXPVGfySyhXp6RPqpRqijx
qpW8lyxOuFqaY96VwDsqwXDn0Fdi4PscoY031oxiaStC3+qVo0A6fNclyLcOyGGB
m/wCCPLKO5eiBMLeaoRYlTGccXyo9zOeOrd06Jli/7n8tb7S9Wg6ihz/SYhpdCPt
ng37o9vsO68DHRr3mRCELZrDwiSuVQLIBs3WIr4GBEwpczG6GqIkAI7C2zRWPoir
a34d2O+a/TRfZKq2BghzTeDsdhYAxyqF7ljxMTgb+dpoARlnX0z9ZOnEA35rfe3N
rSzz6FMp/TAoliYLw5mt1HX+cnmor7dWiH/WAyPfZWW6y54VT7XhYUMWZIxBhLOL
SVeMexIUneBTv9ZZC4TodKF1/kASjQ1iprYE4zOkA8q4YYhHUhV5WrokAn+b64vL
c3jdeRpiQlcgvT8OrSGOYBP/5nzU4yFrYg59K8NERMf9j4fYVP7oB69WY33gPTmL
Wpte2BrhlksGrpU1WdOxKRM9M7SbDM/fsr7ZrkHO6oT2J6YZO+P6cLylHkhe9CnZ
s0h2mQou9d37jYZXUUynM7Kw45cu2blbvsug7MUbxLYCF4LoHrAeQJVSFweSwW+O
Bx05fm4X/WIOnnuCKcc5VDqWr+IsfVG4LISuvuNLALX9wg+FRqXlAb5gxfGtc3j+
iRdSXOzFixzfd+kTlhe5o8vx1Dwg25BJI0BoPjsn/gRkMSbaZgPuEBu/HVVxX5AX
uTYQblhPTeUlMOe73Npu8NEjAaqbEUcVLPzlaBKDfYE+c2b/YQFp9PbPcpqYWTCy
yWGN13UzkhWHRzerJGhPVV9hTJemHNXavPDPsktp7BQu3j3BoEBHLxzZo8hefli0
QhzDe/7LEGrohF4Lv5kJCwkUMy/Q7+yA79N/IPLq/Pyj3DB+Vy9/m3Wv2QK6/E17
3XEuK5qzVnF/Uxfn8oyXDwHoMxnIJ4qRf8mb1oVArB5KgqS61fiJ3ZVVqkeGyBuw
5EXFQGnn5jTKf0jQeSji1PFIEnazD7uPwS2Z6LybNphhIQOFMkODGZ+aQ7VRXKgH
LZL1HZJe3qQZs2opD3BxRnjyFS26uINAoRgi5JDqjiyB0ifiMXpll7+LCdMLMeYx
mrpgweEoYLz6vovNyq/XEIzWzPJ/Qrgd6zlpSqJHpCrj5NcZdSZBT2rmFIY4l5wn
wSasmtHQW0m66y/drawGssj3T3qgVxCeA7GyAS9wPLfxAOcpMNfdZZtYguuAjUIl
XAS2fG0bpLGMl83yr52TC8bjv/CaBRPW7qCV6xm0G7BU0uj/LJZ1O769624CTkKy
WCp+aYVFP3BcqVZuyBqQxbA7itOTaaZIjueEonV+uhj3w51/36zQyADDTTMyKcYD
3bTaCuM9MRVWcy86Up94hnEqj0TlS/GrGSIEjGDD0TQtuh6hgR0mlVur4JBTjRkf
YHRUCxmpiUOd/HW/6k/fAcJmHP+fMn3HLlde8ldCCLLiWKyZ+A1yAkTDApBXlRG/
zokpCsm/x09y1UitG12uhH9qWz6nv61v8nKFNkiJp8HIRQMuAsBcQfZn705HFhJ/
vnJd7p5y00H9MhxIhsrgdpT6hDakVGZssEFPb25Ihup6DBbYYcCMAvVmi1oTztLz
BXaKdK3C+pYXWM+sPYBx/pt/z7Wp9GE/mcLH5hIQqoeD5axoaIMIXo1JcTznlPkl
okQWpZg0PiTHXQPsf2Xoxx6YYW9Yue+dfgvmXAPS2hroW+j93JKxx+gXBWn1kAiU
/gdpyBN3iUTxI0cmWIXOhnxYN4i2qNSqrass5PaB176I/fuiAx0EBnqu/F4HElfm
Zi6UBkW06eYNsi26C3j8coMRNlcnHoB35jLKCPbtiRhd/Yaz3dPlG1AVhrsNIvFQ
46cI/0XcDNxrlNQVH8P0Gqp6PiNaCy2Lq4PvzAA30RLJBABljvfCv5EUFd3CXb8C
/vXnmvdEwmo3WrvsNEtGU6+jjiWiDiZSnQl7z/QAyYomvhQn+/aZaRh0/A0xJLzo
i/PV5T/pJj8DiJQuNUXmcO0ikYsTDP2v1dF9t6jN5/eS37zWFWsS604mnHvtbKi3
HQnCCVdGUe9bhSb4AvFj0yIAr/pNAGAAx7QQsDP8cBGhOY4DdojjxDDdJmXdjHHR
cBvJYbcunTarqyk0VlRAeKB/MJOY8MEjkhMjYvKdPTgmrd39ooCiJCS9wMqwg76f
0LclH890pAatUUbxRIbuHXj+tiTdvhHOndNznCCe7Oe19VIQK48VMapoJSGuh1UT
/zig/NQWnYPczBtQrTyr9h3eFQ4t9hGHIej+mKBwLHrtrzgtMDpbd82Fr95YSHkJ
WNVk6B9pl35YUVR5b6PTVmbvSWCpu48e98SSBxymHFUhJsViHKlYWUIMQZdMOWsX
8M6UJiGXv6SjmT7UsYBprl1k3EhUZotHxYNGzc6tjTY0wGBtt4PR352ddbsvKmNy
xtAMIXlHTfkwuaCIbeqXOzlp+lsG/jLzXvzxOW+5Wth0Im4VWVVg3dnVsut1N9zp
pRN8iwcNqr5bI6FkHPMHB/K/v8ljXp9d0tRRiH2HI4aTIji+CsY0+zwsFXeZWMqy
IRoW0RgYK1c0YoOAJh4Lpt4aeb6OF7yt6qK41cRAtzJ7uX3OA2e3x0s3tO8bTATk
YmGeQL0//A7JOq2MbtjufwTEGC4t3FN+geMocT6kl72Us6WWeEgK4KdU9hifR9Y3
JdTgWTpYob1ORUSjpaL4/djIQ5K9D4p9nRBMolKr3XM6NItbpUVlLppdKkr01LWN
qRUf9KeRr8b7r4hnqFGKIOC5Owwm8f3jWcCb5zCKC0A/vVkKkaJJPuOd3gDt+huX
thM2EwP6+FiCHNMtOK5g1G2UHWImLzvdd+NxNJfbu/2KudgMBf/vJgbSOLzNe3WF
wnfBjniClRihrrfucW5BWy9gud+nv86iW5AhfMYQPFSqKz2C7HrNmlpLo1Si2366
fCKuyLbnhMpR/K0z6oPNT43259KZNlW80X3k3IBQjq1Itt/0+3xtbvYc2ZL/EkAR
d512NrGdJP9+qpx6elG5Z7SmFwdetldyRoejFyGLjm3mTYrhcj4MVNdBHi1U8yoX
J0Fico4Q6CVuPxoE3rGC7fu/9GgfTYky/2wpqyvEnUdgKnJ5mCRn0fKRtiQIeR6i
loAi63d0vTC6e8Jj2cGLtXR2WtCyy70icpGg0CFkj4K9pRj/Ew8g460QX95v3rUw
3Wz3hw9ibjq2IUYu0f8x6CYemG6ui+9iGxK6pV9y3PTID0EGU/8PfBwJ5i44ZvW3
JmIhkiZlBoMDW35KIxjHcHIEdnvzVOvCNZ0LG62fUHq1JiZWX1B5u8ndToB4ZeqE
Kk6TP4/AT3rmM6sWbwRhc22x+AdMxJ+pryI0t6quwdCmHW/r8OJ8u2Tv19wACa++
FqLURL+N9Jkc+Ai6P1YyydrzTp/59acyiiwltcFXYOB/ECnok5DUGQznEyQVE4OU
RpbgVhJ1u9SobZjTOLM82tKSwTAqoWysw234WAxAMlspVtizQhosRFgO/42X4iVQ
kIsPYFHqUFcaI8BGh7xaGSUr728h9Rs7FRHM5bWBj+LQeyUvCwOOGAHnNMfAjyp4
oueQuZrYIUBE6X7i+GPcqXusYJYB0bgXGlFYuvV4vXSzW+7C55g/subv0cUJCw2I
NIOsCNAVJtVugeMEFHC+aZar1CF6j4F2T6RDEYLB09cyyXUh3wFYY6X/1qwj4Tzv
fFYfV65/BdI4xL+Qz1VKkVXa7PCMzRH4dKBAmY9kSXrKDzPvgKi025Mr91o/zqTf
Ej7chueeOsEPJuHWzd0CJ3j+kCoRpk3Twm4OM+r+5ygYFelCW0X0BHgHsabpyH3Z
MIVugrsbApEtTMHL5/KnM08WdeSgeqeQDc3iUUVgCJIXRVC5+ZDN5p/V1YHqHnU9
vstVrZ9sKJDWSUhY8KsLS0zwXEmaZLeKocdOFcgPC7FQEjN6VVr5Sp7i9L9lZhW4
JzuKAqNNRfX4daK1uffYf3X+O5v0mly8IDbDJEq61Q5HTCMnkG9HRlJvxY42W2p2
NGn4kZKRFtFoWo1kzClo5Di7Fsfrh1tGjQ6GSntajjaWVZucnz2LdFqaGSKyvkqB
37rVKJQgv704H6rh3Wti7awjjOJ0QhtsJs15tKDI2wbkMLzRLBMnjt6acO+CntPD
X6EDjCy68JGNf6DGeagDg6OaRTvuvaYQ73Yor9F0dhdHlYoDWdEFb6ee9vP3vT+b
bQ2TuhbmOnzjTZxzYvM+JKdmXF27j2/QLT0hXP4Xpr9k0jdUfH+WqMa5BlPQub0H
UjVhNFzhZk2z92PE0qMpYN288lCbGJL8IjMM+/hH1GYTz96MGm2n7W43P93YAdk9
5vqHl61c+cN5XN1a3Kx7whSLXpyFwCUn1FJfyjStFc2UbrFivcJogKpaH7nu3kDF
UEcr++3n+uToHMzuuRQkVOvduxcoCQ1lvQxbvIIs6BORUMUI+b6heMC1HUiaM98a
hDqzwmKcw9wliJFk3i7GEVxa2kl9XJ9jDqOlC3yqcd/zi3bSJ66y1iC/ey7pjCrC
B64MmPQq37yRUdhHA2xgfmx3ozE8l2Z/tgT+UNLlClh/Af53MIMOqsfSPT5leJLt
ecPN1QACC9yf9tpFeBnwJYtyP1icdNZpEw9SXZl7cWrDTMWB4igmmWT9P3NtKjHt
mRkogZCgtq1/oUVrOGLn40M7s8VwkYQVHB4cR5o0wk0IVW8L7lPfqBMKYoGuBr0n
LnKihcPXA2+jQQkacP2Y79FYMx8Dzzem4swC4OwkdjuNreZ8n/dNNu3ksm5bDgBp
omIhcU+caQKUwJwzAeVNe1HiwIwbJ+pKIw2gYWKkwuZzFr08F0LCKvCFHnZhL3u9
L++LXU/ATDVWyIqUgdn1af5eUmnO4YDU7exFlo89HiLylQYCwp545GtqvrbNGeGN
Q7aVrN3bdoHpTIj85v0g71jtICZBPYRkkxkUTbHATFEpng/SEh/LB0r49NNo2FVf
5zELl5s4qqxyMBfxTgbEhSoecl1VeLEznc82fuV0H/+WdLK1j+CqhZztImTYzJft
7Xjxuu318w2+pBQGFyR9/jBUUROOSTY4xZowdMwCNBkrqN+7fw1ssrrqXztq5jFu
ldZNvTIq4xBHnfgC2+L5qC5Vv+XdD+WKYPCrx8oR4Lnp8EyXVKsaXWirEXCg2dsF
k2sOhghikbVprBEap9xFoBicwxAdt/jV15WjAWzRIVfNdWpisfald73nmWQX1cNu
SQcVfjcByu95NOg1ksmP5nRf2r0pIv6gXTb9Y44F4JAGB7pjTn9sa/6f4wo+zNoE
T0i6zYF1SEXy4J30uoO/ORb96e4GqsMTAsrs3xU1/Ln45SAXXQOWxGDMGMfNw+eS
sVacARVk8zdJ4KqYhUEqVh2D/15rLUDaBB1BIcUT1czvwTETbqnNw/gMikcD0ex3
TcSUefp4K9c4R+eew2Wb6INBhAm2aht+6Ms38LQu8OIqX05vuxFBIhhVPt+Myoah
ph2DnqeIEV73NNixynokY3veU0AdyBgtwnxHoo690Epblfblzos4YwlSJY5c+PKV
EAbxwDSmam7h0qUwXV5oWePQBsGyMFVGh18hBj25HynbndB3ozh1aLyvbviGOTGU
wJWGDs/ZqidZi+VO1ecKy+ll2AA13rwKfXBUKuNdn8qEOSfQX7cKzWlv9hFhzWTm
k28BO5SjZgJobRv+T8YRJ+q/GUfS6txvcJam/GHPMXboeSipbyDd5v2+2HAtrcJ4
OdOIotel61puA/h8JBLOiKjrq9BCQPlDl3VbwnhOrFrFbcLBhCDoj6XW92l38o+Z
UYWfNa5w9c6cJhSM9FHLy7+8ujUY+pAdHSrafpHAEO3mnZ2qGkwF6Tj9zKzpqJSI
x5481+pF+OVKBKLxCGezHdJudNpq1JRUmGwBc5yTX1e+rZ1soC04AKyi7yH2WxpI
IY5sWpwEiiXJrRLT1WJs2ZzdraD0s04MmKkRnY+R6FaCvDrPihxoJXJw06D04End
UIh/m1xDpae6m7f+S+MF33yr+4SfyUYJE046Qpv5/GXX+93Br3gjWpjSwHxTHpNv
M/7hrwTDt4L8gZksCxDMxg1KGI3Kx3124k1PETzffteGCxvJUlbby51NCkbLyH7m
yXc/+1NuPTBI13io1pFTzspyrnSEL2s4W8fH63lnQaxJSDpgpReV4t+uFQmSnd+U
KwWVoOh6tqgMba269lPRz9FcMxiPUZGijpzU3xnBRz1ryEHzkv88Afw1PV791+nn
m0vuMsvyxXTPP1KnG2GD+G2IT4zz/Do/MjlfxnTDoUCdFHztUAj+hHOhwo7a15+n
z+j5AdrTBPyI74WTNy7pw2T0+V2r/NgoU0KNgqmLaJHTnfh1U60fY9WJ0BRARK+C
VIkFgvw3QkBNSAXFHU1DV2pB3aMbWx/vfX3aKt/hbjBOVHGAYomndq35121Yewyk
76NZCktT0b2KMnkKJZ+lMlkkTK/9B5eHrEGLaJYn6jYgGlLWJ+LNjdXBEz+MRPXL
7QnPDxh9xuDMLZRMP2VnqX8jCeRQJoSwF/AInbjo4wrQWj0a0a+CjEJ0K1wGFJhv
zdzXB8fCOgAmKVWpoXYAeG3lB7Cg1guORy/8eZg+e0p5SDGu93yjpEWdhacALMAE
W+hLJtIPgLRm4kYcLequ42S9Kk3bsqKtHc5Q8ZD+VqHvnLtZHtH7p9KtkbqlJ8p2
Co2i92foAKpUMYkp0e3l845FZLGfZFIEEm+xV+sNN6OE/+ctNvn7pT1V9BpsHHth
sWiyiyoCJ9vxiATTzRD6Ew3PuH7SEwyHxI3ogcNVhQhRl9ggDXzHYwnEyPQugozc
lh76kwbFH3Z4XRt7Na8IVyzOdS4A1S3GxCd3Q7G1Ss2GC5oValBsZjDweuoA4Za9
glUPN0C6lAEEjamae11hgPtpGyU8FV7AXPZjrcFR9G8n9Eh9s5dNcyn5jc2dxTxJ
gXXSsDDulnW3GOmhJIrej8hwe/0pcXzbEZL8nnRxzymGo6+J34B1IUM8mG9XXYaL
5ZO2xqJiKVNl7eXeHYDG/X98kOCtfrT1vHB4Tyy/lPAacNYn1c+JeP0lCmF0dm0Z
umg+y4x23dsGKyVb4Gkg8MpbLmp1Whz/VWhKJ8+7Hg5k2L7citTfATs9KD53n/kI
j++NvPbYw9MyOLURSiyh3MlJFzn0DFVrMAUXyRyDbxeUQdkUeCjRW3zf9lDZf+Rm
USpQhLa0pVF87mXrmqtKu6zpxmdtJIC0mr9OLImbaCu/rcpLiySZCkWUDJeFQXga
M4+uovrIjrysGdm4/rnzcw7UamADrILWL4dIBn7glIAyqkqPnaydRRCm6GJDAS+u
PNDnW88/W66l+3B1jCnrr2gpiyiHyLaAEnCzE7EJaY3nv0vjL48IbNb3Uc5AdwAK
tR+wgzgPRiOe74loWa9JZiY8bnLjjtoRsQPzmTVPNDr7+LcrJiQe6KgacgiOSYnd
YPsz6H9mLGx00cc/2KnjAv1OcXNnv9iwZqCBD4+vFGhEB3MBy6xranWXbxoXdGTq
We9MqaM3tksih7be45veHk1ZD89PGPBF4PeXeL4CRqeXudv9R+8qlHIXcBpjWBNY
2o269ZfHUn+FrsOR6I9FA5r8jRxuz/II1ip9vuLNYjo9lKn7uYuImJcp0A5IQ2Py
YSqeNYXCTqCvHGkxS1DdVWNl6cGYUKB95mrMHfswkoglLRFJxmLDzAJ141AIQsG/
fU9Ab9p34mANIpjQQ01DCUp8COlm0SQlZSZPQ1C62xnduauk0Kb0AxFfrrWBuKQb
lMFarT5dz+2eVZx9PkPVuBNY1JRXpQMsDOb2UlTX5H0ndGZh2GzrJqGPw3kqt0ox
nAPa0GCpuKoI1uozU2GZ52UJGThE9AaGtqonM9kKyTJhoYGv75A0LEALv44R+L1n
e32bH3M3ggsZonspm/lrg54JeQGLB5UDbXzZam14+Mf9E/KAdxbnhCSyR3KPtig+
s4w87fjvoKcCSRvt78070jCjKMUhJlM5vcK7gbusoejMEth8CVsDX1K6yki6NSNb
p+FIQwU/wqU943IynnpbVVpHtercF9z40dlUVQ5VmoYt+lN11CThNHJbY/Xz3Bi3
ke75gxe8NNgdZ0RoEOrMxspzl/On27IdsdJ+641YNDG0NUQ7ePDHxAzPjNWyhI0T
1xnfFaIECGBN9dMI0WeKV6dRAkorw9Sb0SHB7N9BjvzZedJMWpnnRcTLClrGqovI
BVUWMfNCHXZjQGwfq7vX4FnEACqGSzd0tZvYas6cF/1jK4YEZiGimXUVzr/zI/vw
kp4jZgXmzeTUCFccCoelGWPccWRt8VYFtcD254AEAWVC+TSCc9HKhJfas8YUKzry
bZK7kIaYCp0XgN/eV/M7Wnw3T0KcEnHczPpo2B8h77uQXl7gLS9p6Gsdovk3Y9tn
BQl3MeknaDx46evUr99ZuSRsm9RihBlRm1O7tRdfK7y9hsEHfbG6ubqmo0bLoZPx
MHCemkQEkqw9LEeI6s4X5i9P5T2fKBfFmPOEFzHTeLf8C1M7cKUG4xwphRABchpk
4OwaEuAyba3IJRuPFQx/44mfSspnh076T6fRwuI9DYRmN3XA+4r7NEAUv5NsxMYQ
54gIDigA7L3b3LDMpC+2bn5Cc3c5pJKl/ZGjTw0CUTfWcCQ4AQk6ghXP/oMMPspw
dVhbvZdW50Dq68EdsFoJiCFq8h+5Ri12to1RaAHc9NyDALSODoysxvp99Kpdtk4K
szqKYMU6Fks7e1VNrqk39vBoXgZbo1HLWYcSDaZjjAc6oDJ5wW7bMt7kzB3a/Dbp
/FNk2X4M8zrYB32auGa6Na2PBDAg2HQ1JwA/9msuyFdLykzRr5zNIwPbzXh+jw1p
sAwNsLYxdfuoTkjOMh67a4tePhgjQrLsHVkSFwXcN9JY2lyZ7XfrJJoE7i5OgqYI
HNyHN29QJMkZwFbiPalG7OWAB2m0oYDf7QTTi/QPOATe++ik+VBfiYKda0cwqjhW
gBOM+N5lqekAchGVT+Zvpqaz240ZO3EWv4LcofRJWT4MrH6yF89k9a6fhBfPJYVt
S9mxE0W7RgvYnCEN/9wtUxThUZ2TiO8tqP0O0V7B4i0NFW9BH1z30aC1/+0vwAVn
PxIiFIE18ZGXcexh2wIuK6mMh1L2J1vA5UOLcK1oy3Jt4O2ZDI/gd99Lf30ePcT9
N4y+4iP89mfD0VCp3g2D2UHREtteaPks3icdWRT4ITTCr4Srxt8Rmd9uV8l+q1U6
4ntMN5wn/S1PrCD3LTR2Bg+LhJ3qMPAlu7s+/KU8N+hMLxPuLzWF7Esq/NHHhYM0
yrExFJrxNFMV6AOahpzOHQMrbLHxIQ831ek4e88+Cw5CUhunmn/jcsUojlUFdiop
irdapx3Fd/+WVIFwTlGsoG/C9onyRhzL2Du04WC/HYAfIpZcHNv4HuDbTFspIUfj
G9gBX8axH6k0M20H+L6wqbtZjPGAUYqtxZHtrnOUVZryqJmm53bIKdgDE2jh/hdB
ETtrSm01rncOgMTLE4OpZytQnN/FR2i7pWLaahHEOkoaXRBvPiIUEDqnI3EMLawr
WHpyZQQWhuM2fbx3Bv2bU5yJgWKcet+tXFyMfDfJ8okYnSJQbXQWbHD0qgv5/qyv
BBhgAnKsPHk1qRcKXK+pBqohO5uY9tIyimVsCtAHQp8vYSBvEt6xwl6TndjNt8Kt
x5f667Orp942HYH7blP/RIDQbD0hMKfcG1/+ruOHFNYsz6hNxlXnylukqPlIvwuO
B2OEgAHbneIt7T4JrD/q+SQ/OKNKTXA3UGrTEktvFPxy5vkWjJXfdglCB/CV778X
7PZ49iSl7KIQQo4OXLdbB5xoKQMFBZDS0hflHsvzdbNpyCQpl80khj5a6dGdGkYm
INXXGtBFRufMmVrjKKNxHorvxITv1Twq94y+ZIJsic1tEDRZV2mN481RuJbjdZ7J
+4liNZa2cB11Jptl8zMq9imV4FHQZ6ZweKCkG6vHA0RRAO9pkXAz8ZeMd/yuKOJy
9O3WebSdIpMTLqE6vn7jCHGpyK4ZYs9JSbt7RGYYHZGu9hLZwzCrvW8MiARN1uiB
68Hc3S6kGRTQixy1N5tKmiu4aAeQhtddu3uHlfNtrCfMufcTTOEFNIqMXG7bWdTy
FXsxTAE4Q30+N1UexXMI+Gg7y0322CTqYvTjZZG79ofg8cMwk2RzIY5X799Pqi+C
mCpTQuFnrf2D35RyAQNoSClBX6l3rnUreOmBM4dG1NA5itjkZ2hsRyc5z1EIHtqv
KhqqZyM4nocQ8UpfQlM8eb76qlq8B+QBATh1cwzYtvaiyp+LRl0XMbFh2+NiKUH8
eBIjqxtHo5b5/66e368vzxnpVTqmnn0nF2d5G0wsaXOSnGmRLekcWILWXhBaMUNN
aJXG+LFQCuXejG+3INREUAwEKpN2MVOw+o5aYfzcYfjn0E8E/S8y3erqd2KtDeRG
mN7vpXVw8oE55LyUJ8Kit9WXjVGZ65+PFsH9UFG5nv50hW7r1c6PA7ybmlNJAtmK
80++09MOMhIqFVJCU0jGPF0LVQQhbT5izNvmhxQcbnMBQW6WFg2ctffUFer2DbS+
qnL7ke+z+VEFawd4vuvsSIwmJDIBrrCQELAo6t3xixR2VH+LdC6rkXEeZbxgQHNH
+saI/Y5ZA3XFscZRAx2V0CnQ6gpMvLl7N7SWutxj4Pw1GEUkJQcfSYoHwwdbGkHy
1sxyWOesEpk3WRMfjr+qBPlcBK6KCJQU3L7LS/Wmm22Ao4GrfMW3U2MGiv3mET4J
UyjhTjS58PxvjKl6vjcbTdyDMzohvllB1piI2Q6KY+S40EyQUKFpanrwqczMSRf9
sNVRonPsVYfuzU5p8fyU1knHZz0V+jxQ+tTdyP4cg7CmV4b5uNfEVBgIjdDikc10
EMmTCTy2c04RQS/SgjrmfYkbtkb3mGpT4cPMRkzryWpJgm0k368obV4Wpxt2DuJC
o8I+YdYzdZV4lnddd59ArLb5NGz5P7NIFdwZucplMsc0QFyeYtZwasJ0EZaJFEmk
n28SDg9qf1s+9CBdTqpzhtrKXTL/53rkMMGogcVcYEgjcjk2dypCzJVzx/CAoghj
dgIj1yV9hULXP4EQflUUTTt9WQaBKhsGHk5yfB0fz8ZTdkxRa2H+YGniJarWRDE2
Us5+KwWZh02WzpL3PeYQAfDJhVoKjxIEoBN2VVhZG3rW6rEITITMUteHiRrAdFHw
N5ucUfewA2qG8hJAGtmLEbBXLZ1uA2AODyDtyfFeeTQzuHmoJBQ8lyW8t59tAj7v
BdmVlFh1apLdk5lJXYXl5hbWsg3VDftXaHIlOt98sjwmzSnYlPdBJXJjn9wUpLOf
ewK8fO+bwBJx0245aCWv92Gmxc6UZzst52NFL2MUgND1YyCChNck9qNRgvP4Buqr
IgjYr8VTG4EEuJ+A6iNhv3IXEmSDddT/ao46NcLDNjFlQNoRzJHmCWechjcnuZT+
RN4eJnN9OcuiXald5aaHjYrFGJfe8EdyjEkWX1zgafvTr7AYEEMco0WHP7nYRbWj
WZJPb3oDJG6XP13VtdXjZf2F3jPXfqbSj0WrsIkMWp4KUMYUI4fTZznx2Ghe+//s
liNQhUBwjhEc51bojPf0Q8K2t8HMKGFHUUkTpeI709NY/g9x7ysxA9pdRfn8Ssyf
AXXslEYsd5Km2LziCEDvw2qzRO3XjzwRjTCs++ZuiEJQFOSP9U/VShEdv/2xigwT
fqKOdSpq+m5pF7H58GctP+51Us5cPCcP6iAHJ6MhOHUhRwYSIjnbPTSWBNc6hDTL
2aomLxv2svsZ8ktPnHCA4d+oJUeJKOJP4SHVfM6ltijFI0rlWMVeg8b/qWNmEV8F
NCWRTs3+CdZ0WNCABssjK7ZIUxfmo5b4jOXW/JXGyIL594BE9B0JyVBOzFwyyoWG
sAMG5819Nt1FAiBRwZ+2yr3+t/oRQecskYaJCaR/wysAjL9elPxhyf3NhjN2+qYP
ilC7pEOoP3on0juysEMzGHsnbgGbFr+F1OOUhd74DFB/MWl0KWgDyF3Sv+3YRFkX
kYKBY4L8SQDme9IgXEfDGNiR5YrlWF6Gr6F0HELqn1zec/dRGrdKPsAeOEuecRJf
QrJ3SL/sogZkL6d7q2Yz5MibeDgxX1xb+HiOVImk47mxkLUapLjAGiTt/ccv67un
Zz4v5mCm8XncoKx6+yW6OA9a8tWGZt1WMe9FiDWeSXdMIKdcGEUQ1c+S8O0n24HE
3VA5RUg+V/tHo68Cn3WC7D2FBWmpa+cqI2EJYj5m7EVLhE/aGuP2J3qIGNMpr5W+
niaWmJ8hyYYnlCNvlexhBeIomjRuOtjNwYTd4ZYsayDZj9Z80A+mETd0zR6FUktq
zhCpgCB6J+7ShuPq9OMg4PDsYjeT2jzWuTBBWKGXYSVslEY+jpgieB/Hnm5OCE44
4JBn9Cet3wOsx5UTCDBBvwJ1KXLjVUsDD0pwAnGEnjuyjpiOGvagqewN+vwm4Bee
PouooCHpXpeuwKrbG8ho9A3z3YeQXs86+iQoWDj1gL20ZrNJ6rspSxXnz2gjEplS
cHmuP+5bICc9tqhBeyeDWtx4oAIK3EX+THdf0684uGg5LYeiuRjVwos5KfeZGKX7
CEFnITxRRuj3HbF2WNKssq0J4ktezXQoHjky6rSgQNiizLRO+ncgipWgrucUhlDo
g1MP5A10W+vK0erYI6TjIPEAtC2jwfXpLClMWzZjBT6PbEqJSLYm39ozEUz1mLK7
wGl9VSTsiXj1fIuX+Bd4zzhTsXiBHvoHoxCsxsWfy42LPiHPsebXz0dQ+06c6tU2
TL2GNZdcCGzAtgyz/PTQinCB7J5bbmOSjN/sPoKBQ/3llRd1poe7ds6PMklk8Zim
gP2/BQmQcqH+7svqDAY0qWw9ye1e0A1idKvTernS4Ho6u0ib7gsxNBn0eiQUvpcm
lmqfXawckF0OnNxyk3MrD87xKFicyMvHi8A9qxsRNfv/LG/uCmqLF/CM4FIKB0PW
sN37Rpq7fsxfwje9MWUxZiY70RBEEQhA3tMRHaxRZsWQnGR0o7Jt9pIqTGjTQOR0
4YgJju2ZZmiFVnU9TnPgMsb+s6FB3Q0fr1oNwrUjKtam6u2cD6gUymOr2ldfFr/P
sspXxRVwX3yNgQQWW3jiJvm56EoiossuKd6USdRwkkFedykggiwst6QE9ZfakTAg
+/gcDPiOHzYNmDUTPbTMzccGKvv8CU1M96ocIO9NqqDAjtRD2dO2eeYfCoreoAoY
ROVY9KWaOuPY+v8LBYUymooG96ZqDVdr76PUhnI72kXYFBK8ONgwfiFklLCMzR78
6Tb1NRZqqXiyfrpzTJ7hXXqsMcCk/N1SsOJueQdroSS+A/vQsvkWD0fS0PZrFJN6
T/MDiJF/r0nzOwcCWqbx6UvHPZ3vUjq0XE0DkqSAIJL1TGcmH3Ovz/8MPAZ8PvB4
pTfegpFzWRVq0DHdynW5iHwzxXQdFWvTb0GJmwEZcnUXOFOX9cstpGGguI0A7C2C
OL8yEHBTKfQUoTlzApaH3nN9IhlqvTeb6VEUjNy0LpZFi73mtkDJXWu+EAeJXmgx
QZpiJ1kVE7+mYdXPjH3XIU52jWZXTygHjo1/+teNOKxq4cr9IMlVRVUjrzsGOLZd
oLSfJQlIs7pjPwYPLn24hXtDvNPR0TXWPxc6JKO66UEqa27YLhULFgJfUZqMoebh
rlboY7XAQhwZSKR44blvJyipPos3pvw0SXc/Suh7UcMU9cFtFO6WOfqE5T4WID0a
GGiiWBrgHHQ7ffnijkiQN5dXi87T2/u74Ak3ry4dVUn+/D2NHOeQWPCDe4iNH/9y
OnbOD4KdwhXwraPv9bcjQSXVQHpJCrgf1UYQI6Lj79PxFkUmMVzKD39V6a/gKLAJ
z05c2RQ6pUIiap1c+2Hq1wdfoepzDnmn/gTP7r14z7cT5PrISAxmv9F5jm83QcJl
OhkKxpE0V3pXPhsfh3dPW5NuK2K4iXHNyUccVU3lM/N/hw//4814R2CO7EOOKi++
anPH0LSPM5PVYv3mo+Afvl4EoeF0o9VWxAbGissqe3IfKhqZbtnxarYv7COnkbOh
2rWA2e4/GCJA+SAtpxbhhXgMhLkGWcxiN696fyltJuPWrWTPxw8zf5VdmcQoLVX2
fxoArpdl0mmz6puMb3HYo27ANzuK3pdZPw3Ij0wiBWwJ3AsCqq1rkVUdH9Ecdjs8
SNayzPvVxScykS93e+3p0gJoFEzu0O/pPt5jbCOjw32R8BDF9AH5tLDFpw6Iu25e
U+/TxoBEol5f+PzxzpB6MD14IJ6I1r+IkEW4zxqWFkXLEqaWGwL7N0EIvE76QhJM
ZC9slJ+TdF0RMUd3IKNmBn+vSSdVMHJfE/vd5Vi9r5JXh9RDxIhGgbQLrddLbdFs
h5cZkMa76N1CLXN8vWlhoO+itdrn52MKBL1U30st3xvfYN2FArCTqFuR9M92fQcm
KUtch7AM4wTAqeQFH9M6z91cnqPU5mF6MZL8ljHhuEqqvw1iDnZKc8LDsEoa0JTR
caXXFtEctvLyFN7aDzUbAwq6yClzDTIBKfWrpxhv0vF0Wn4mlBd0fIdJwJVGD0WS
p3WW9HLqrBEnqb/ITRtNF0o7LMfu8y5udzrZB/4GwTTJD3GF+pvXJpXOJ8lrmxyy
pDNr1uqBFY0PIRPyQYwcnNUXAunD6CovDFfSL4djwQKVdK1FFxszVjdx7FaNyhwI
qED9O7yxGsizMTqwdHty5lEdMS6cP3ASRMi3OzB6+O2aBS10t+Zuly1qm/fsdvW+
aoO0KpPTHMk1UolZLMhuO+4GxsqiiuPLPhKPU0z2iCZ3XTlcgzJ+Vp/vaIlnSnGX
6c2MWaCHF7E9gS+9Hay8T2fa/K/gQz60T8xvFzvYTN6f1cHhO9MT+alchFPRPIwR
w0wYIrrPT2sXvvC5t0oVe8K87JfXSyLwHrYtp6uvTT0owICht/l9CTovQAfeaqGO
0Dn5q2CWjwgITIOsZpN/5IojE8Ld99Duf8TkHbYBsFJsLFk0XzSFQVHT8Ufn9zF9
SV0ElyYj5Z7A9su0VR9QZCJjPxc0wENEzMPCs++cTHUVxbqOXUmDi1GR7LHsZxKj
i2FojV/V/RavgsWrcG+Uq3hY+AO9uM3+CZgYLe9ClhK9DGOMcw1sIk6gwIc+TUyh
0VD7u5CrHed3vme1B2+5VmOOZ2j0l6yQjv/m/MP3lDIOl/NDZRN/4QQlLfyFZ8uc
UfAD846fQFiS8109iQ87LU7gHki2dcLdji5/psFMbB/86Y4XbBeROYK1ItImWjDf
vPPK5pi0SsIGVDBsxS1pHD3xG7ZvL78KDivgAPeonhTqBdfWvRlGmZpfKhquq3SS
baHiryG0+CMrsB4jniMdTNC9ZLHmYRARUE0JSLfkGZXr1Bq4UkC6XLJFlWBsApKB
GW4NOrrNd10XZdd29OLMKsBtFdXaP910nhc82y/nRw4cL4+AByB6pkdp7Jl4exNR
xNYo2QQDWq5wY6sQsW9uVQd7HJ6TIBUla8D32Lj4EQHCwCPySMB62Pm7a5x/9gA2
J3EMvp1JDFYDbSXHpUv00STbZyGagcdIzZ1D2SqFiVLtk97LGcoByD86OnGKR8sb
MW90LTzaeuxkSqyAPRZIcr6uFctfbU4qqQPckuGrjpQhOjDbugb0qYPUVNugc++i
vCWcW+Cq9335cfpLoRkpKwoJPT4Ku6hBFG4LVr74t2H8qN1yTAOFa96JZZdvzqh/
HZTxg0cd25FKkss0xI0g2VXLve3b3LXAmmCaWGCB+XVIdBCrztN3EY28YG6dxh9L
Sii7K/ZmD5YtEpvtEOPzSCDUhsrvkbetW9m/083Br6s4p7IEcj+4bsl9SzNoqPSQ
LwXxbxob8VVEESW2izPg/bqQ6SwM4RXdDsaP34S617cibz7t3CHoaMt8Bh+rocdq
bDQr8SzmBG28YGs3h0CIiZ0LFWA2LEWnWqBLw6vE7SIgH7J9/OxNWvYy4S7ZjHHF
KLd6zI77TnqX32pk39ydbJFL05Dok5Vt1OMOdDuTULV0UC316p8GcirsXn6G+/sr
MWj9ncLAsPAAWekB8oMMmvU5FLVft9NXTMippZOaAzCquSLFtbz3xySsAviWGE2Z
ZN7YWilPg6uR4zS4a81eAEqZc+8lWOa45h0RJk/Q9LLF8NKhScMKcEbD7j97Z7S0
MymUmLwxQ3lozggggN0yNE92N26P9a84rDbzU9zdt9Xr0b3VnXX+1z3rmVZyLRxl
uVCZnhChmCEBdZ+IPMcHlaz3sTw6v9jwannExV1GVEhFgojR95mpSo3FHIWm4ZCc
jf1+e3twP8/uiR8JiLY4fONL3r3BqnxYQy2/aSxeWIxbG9IqXlM8+hbbhitROPxF
wH6VQ0Eak4sNGAu23YmSbtFwJBc4x0U882JIE1yI2sUAveI16QfH25FXShlnmw+m
PQN7DvB8sL2M9FQ1S7YYlDTxMnWV9Tb+lIUbo055cZT0+gEHPXqpZGMs0RPY/knK
LDQnbOhHbGBB36NK8aj69CrvMVJSs2BLSX/cLySjJtKq9k9GtFMSFOnoLU+edM3k
F5fpfT0iEihfqEz9B51PHRMMwALWNp9aFwKEYXMs5j2l0Dl8fKjmH4k5dRyqHe4Y
qtfUksECfRYW6f65kxebprG0hANd3tpy8KMC0ikH/UTIavu8fTAbzesodoWgW24o
dk8iXNEv9zXT80na5XYV4jknwIWqP2EqdJe3xShGr/VfL6KZX6aNjPoF794On5qN
Pc/Nknun+R1SQbLaL3LTtGPcxgTCfjNWybRoEibkDdxivx97FRnaWTqxHmYv+N9s
Tx+13TP48nG6DnrtPVArkdQju9R53Q5z58DXJ8iXzKYkFu2RfccUnFnHmBJSbKYb
JaLqeqz8pW3b5/UCdU/XZ/2k1l5ZbwblGxfJkq45zW4vLyCuyRip0+BsVj532ggK
rYrPe2Sonc9CjrMyUJdpSYXsG+p/TWMx4bRqgywxCZh2vjUrL6wQAa+3H3d9jV4+
ZFZHs/kgRjY1MTdaz4qd8eFYf8+6xAlDym04bvz9k1CPq/a9KAsEpxHjtR/Ksmmg
Th/XRN80bp/95MVh33oMF4FYDmzuayi/tAQKFrZKl36rZ7uZUv13a9Jl7pbX4EaJ
fk4NTaNpks0U4BHSY7W6QSHZ/1LjW0UE/zGXO8ViPkMQMiwYxJ6kwbiAo8qeXL6n
6sSvk/CPQD0eaK96HANN3OGrwhjVH7HZM9Y8+mCgJhRLJY/b2C8lIWDbE8cPEZCA
lQ5uofGgmnlLTs2e7daiRx0L1Gmku7mRmLwOUP2oWtYr22fezd4Kt/EM8uuWlKvk
jd0MKnladDNSGojyaeAS8qw4um7JiOmMzIT2+3hL7tQ7f8gLFXS7Q6eX0wMEErHf
pVBThgWtFeRzpVdksQl8I0abIJQ8Q7N0gMhANKHPgBRf2tV4LIcOLXoEhDv9PQit
TcD8hHT3H9zcoL7rlCDAv8mFekkS+WT38IUopNO/gREGYHpCY449Gr3isYkuNVZW
rozxXUcKox1RQJJiCEiduV8INyUQHH6Crs65VZ6SKEBrEDw9lYnsuExDkrNL2RZT
daTddUIrBA8XbSsarklj4in6wPqr4dTmn2uXNrUUrv6ax1dGVS0eALPS5XEjXMbe
7OPU5cL+9b3kZPvIipLrxzEaLcNHHyanLHSAf7T74Sfdzq2VZMwLOoC1//ruSSI3
NZBLLIK/EqeDluu5BWlFGaLeAbeBA7/81V1gzuU4oo/1fdfZykznriA8gOCFFax9
j5Lq8UsI2IMtlajSSq+9xi0wPjeovNswGbAte/oGMxOsbiAOmQA3hRI2I4dziKxv
bRPAWeAYZeEEYBd1iDw26c274k8Vx/6Hxg8HB3QYqOVPGMp/pv4QXKzTfLEwcOFE
OgimoxOiyc1xMX3UGsPzpv+n5MAYq7/yOMOxBCU3C5zmKMvxqfATgUsCv8k70cDP
olb7MIKk6DoMeZtWfkNJl2S2wEpFtQgm1RzLEiWZ8obPFJVGsPKWLr787GKM3Z7c
rZGfPEd68PY2nVaZGypfIcoVzXT4huYTUBUeCpFf77N2wmr2eDyU9Nq+0iZHlrnZ
NnzzSsK8oM+CrnXDt1t6foJQxtwM0XgrbuOnpnH4s64WvKVdtqLCh/6FTQZzSg/3
H4kOGmcCx787JZVGijtWFVRw65SWwR9HOqsZ9RhkotnoWnCKFUZlGNEAgh7C6iJE
zJkqC7noLUi8cJ29Grf4TqEzSpj4BAaRyLCVH4mBwF8pdITBzYNYBhV3Cl180t+T
AlcJzF03Eh0yil3GwA3WqXHvvcDtXO9uFqtos25KY7Tl9OMsXtYWikuIjtUAfINF
ZMRLV/NL9Dj0JkhINrIA90fzHBqNT/s9rXpX8O3f6+Bv4L0O9cy3dShw1Y7SYzoG
NqUgvhTNdM36A/g1YSx3XLVQxs0uLCy0oYXmGmkj8KvFr0S7erv2cMNR2OEEoVX0
eAQh22K19oTyGsAES1MKCUzAODXGVFPSOtYTyblcMY6CWZ8hkBbnZkp5e1rAyU9u
NO5YZa8oOWpQi5QvXT05T/+LzIVkGCHHeHHB+dKl5eJempvYExJx8oTrr9aGEJsK
AolfKWmsCanU5wK+SuT74+jgSQqeb2vCwnR7jFmzR/7ujlu/tR5ETPrHWDZeJMEh
CQC8haTugQqGsJSSWrbl+J7veOeoordzt+BRgAHzVj8J2UnBEQ0QH6FmVmsDU01O
xFPMFthhONDLUgasBBdMokz7GFCqyVtwDxHOIMAI5VorRUrlYaleB+y1I7/Mo77t
o+e934cx4YcXwFRlhfdPXKJ60EY+G1dhxp1MZxv9xPAN23v99e07Khy6zBQ3kmoq
3VmwNGvzvJBAnTZKohn9jbE6GlO2esC1Ax/lmgvgwZ2hoxY7RoIPr5mCiY3719rR
2Ib8950iiiwrR1SbAPLqDj/t+9yDppjcf6H7ufsB1wrqg7s+zr0l79cykdTWDoXr
bkm/rWjeyeWAj7x+XXRagSchzrc0bSyNn/D8pF1nInhD11P9HaeNAfwBygbPNxeY
bzB4uFmqFrBC3kFNh1wm3tZ1/Ns6AYjIkemnbqn4UDgx/n/rkSxjsGXDoDyIax+1
Fud/P9dGTmLldOAzybRIHQtru+qkK4FlUNvfmhIbWQIjlopAKMSe0Ea6Tz1B07EI
LADEr4A++RUHJI6Bak67mtLctjyR3JIFsgsTDs8iO/ixsweFSAjjJbLR5CfzuGcU
ngBAZbbQZ/7Jn1f81WmT0lssSNqc1Oz8zCwuJmo2JyEzZyq0t8WhKmUjIAWNiYHI
6PouHpEluQb0LkSGudF/VejyMYke1YQZCkcQy1xmD9DbXg9O8dVfY6shJeD1x5+X
cNp6tRF57uam8TyOkp/5WL270JIolYNcsjyADKaq/7FMby+XtwAGe3tpgZyblUTi
Wb/GoVWP4Rjxg38lX9h8yPRAhH6Hk4nFq93VM6dEXG/6cWSXYM7a8yWyrXMehZt3
xSsSBx8NAbkBY/Chw6KM/asC2L8+UjKI8Zxh/4DALz4ooKkH2WF7lpmUiEq7GwY7
NAJR7X9f5WFPicTE36GfVEdECLgiNk4bc9c1bEt2IB7u3Y7J1fvzIsHm5KUcy8xS
pjrNT7dJV2Vc9bh421AiZwNJ5sfWaEm94GSr9nE9KvrnlmMMV5LP2JsPWeXbbWei
6z+xAiHzSwVxBe8SxhGeEon5i+IHlHM1IoYrCXUpmAqql6uzh1JVakNrY5tAafCv
VJ9/Dtm3GH/EBl3fDIkPh381sUlVC7NyQmR+2zyL+tduO1vW+1jVyz7IVGhxY2H/
mT8o1KdDMR7tRnzoRuBXmkagw5yT0OXVAOQY5epFFOe47RzEWJVvplfgTEaXoP62
OkmEWW3wKr7p85pa+A9VNKKOD6IJ6MNHvrvSNwHkfK+gfj354KrvnYlPR82pOK3r
Wwx5CVtdRfbnMt8zms9ucz8ebH6MQETRIX0kO8dmYyvN+dpj36B2TgCmsQfPgc4Q
uXmXbRrh8pVBvLX1Q/Wv9r3uzB99d+SsE7AXOOqpI9TpQ00Uu+6neCJEI7FUeFXH
R83I9guMxCpOH8PfZ4iNqOKLzwGtlLGrmKY6qDBu9Q/lQed1T7Spdg5yjHh2Vk/L
7trx5lJKfhOLNmdqaTXs5Yr0xWiWxkZQ/qW2mdJ1KCyG2BeLLibLvN5rO1DEuq+G
VVd/wet5LN4lW/8wjsWE7H47tYhKlks5Upo9K9E+6LsEEEKYBq/aLPos8JP5iyAr
2rFKCicF1ekYmyFmwX0lPp/j1Qzy7WvjUmSOojlg8wNkhCj1Voh6Tr6NShIJ2Xdt
Ytmvr0VflVt+XHZEs7GB2O3zMwyrQc1hIJAwaX7eebO25tYQKiiOSaRve26+Dtxy
6JZClYcLbwDBGE6GeO9ovYasu7R/WbqmWM1HlFjDKNzC1BwWTejIJc3YSjg6cBTv
RmEcp1tym2tTRfD+LHUakWwchGO8WUx/TyzBshiBuTonlWbfKRJFvxqo5hy0Cppt
vWIqwaEfA8tHm/uNmMLPsfoeKayzKdKO4o//oQDA0KR4l/f+n6F3qDjw3E56cRhc
ELPyo/dPyrE9LmdnRSj6zfSX3Rq2u1igqVqdsxTtev8p//bagjIegfpuL7QLFfkd
+Kybndr9V6L+0F5d46FvHTfDKc0Aa9KKzg0XPPeQVR+JJ5bmLBSup8kCky099Bna
2H/iZSWJNY8D1ASQ979mbKoWsDwDEzyI17ANMCcKsSTvO8ZMVxhAwjroP2yAx1LD
5jhJ1SqHNiEzg1m5VFg0FhuKd3T6SymE35NJyfOtiHLNtlacgaxx8k/wLvx/0Sht
c2Ri1vCbJcFvl8FL1QtnIuj2S4qepSzWFlluSg9ffQ5AkJhY7zWuxQCLuBtUuBPu
lUyxgPfW/zchsIJwz28rQ/MlMm1CKB5HbURgTidAUzKjrdsKxKds3QvKcGm+PnN0
t+nwKRCFSpDqalb0R5luavbyfhWwAgNdxV4p4jIdal7gGTRoOrJDAkE/E/fYgyTc
DtZt/EGj8cNKNXCmdqrFbq1QJt52FmBzlrE0XNE/fLPDN4OKJsQd2RmZKbdz5cud
SEadS/QWuSelgiCRJFxxrV6NXv1ctZG6HMEBdzscWDncCbQzyFkIjKkcp0YHpeCn
hTy3OcZ4VvKOJSn+L2ZbmVgA64dOZZqCcXLgho7t8tyd8j2pEwk2hIfrqZ6MNigx
kfLfsXot6foiua6cxLwNpllVCPdawxMpnaqw/v1gvLF7QINtnwozNdjVSS327eo7
sbHtel4+OiUh9yK93g3/lH+3zuwFj3vxZykXZbxTeJ+g7nNWYwI0lmvChi5gsCdi
izz9h1h00awGLwVgMNzzWTSFf4umTGONqw5fRc9Pw8uy3FRTEV6kVWtO0NUq4UaP
qPAxxyIt/NdihLvw6dfcM9pPxjzylWMNHE4fVt0mLFKP1GMUBBnv2QhJjfYsce0U
gu+4RmW60pXV7obDo77gXTSvdsULaNomxx5LexYD2ctZGfsB3t2uwKREhDEmlJCD
JmHGgtNrWRCD/jbS9TTmVU31AqCadtEqdSihoYIJNI7IZKmjrbQ/oxQHIBjG/NLQ
PPVuVKJkJXqVj5XmSHWVYC4aCHBbyaOfhIFDSxyA1Dkr4B/BHQOHkO77qAZrMNaH
oh2S9fy2vy54rKN8NQy8K/Gf2NoNoHaf6sawTlG5rJ0PvFwijUkxGq1naL+V07vk
wJo/dLxmDi6GkpbDmjvl7vBkdsQjDJm0lzDomIaotRgLC43GGfC04xYfCWT0buYB
HXUYbOL9ciBtQFElNkDD/Q7mn8UpnfLSqfWmW3SWBXC+t3taKJBuN2W5cUY/MUGN
Jflq4bLk5W8aH0jH7GiFPpIxqScF2enwETc3zdnjGKLAYJFzhROCmHrZIW8nJNbx
FL8BHtPOiQotz0jwtZzqi+porBrxv+8UMLWbfZhxnqcwEEdhX4ovUIcL5yXcuKha
GJdOrDDZgnesrhwOtZRgptSyaL1d7BsKBh5p2ScC67shMw+LvpLtWK5hB0egu73f
/EZqN5ikU0fWHrfmUEoJMweilTCYuACBe0ZbYYMcK7iA5npcIPntaQFlPeAjX61z
e/arftGe393hmEeYPQk8u4qb1ZmTONY2gaDFagYZypbgQGcvlL7go3vfhir2Qo+F
oMjrkOxqch2D3ppF663foA5ZXEx4Gt6K1YYsPu2+uUvZMXmUFrzy10gr22NbjteN
NEXjvnAnro9uTP0CvppNmmIwQAEt7Y7mKwlxlKGJqswAQpMFgisMj0GZ4ycE0Etv
N2XT+YiRiTWrp0FUOgIdgLJs4ghyYvr8rlvRyTTJOfK93GrpeD27l6VArRiDm6Ql
KZ2ggFpSxMXaOnberwoaI7NQk8rw2BG/oNl61R27H3vojlXkVNEOCn7HtGFiNkkZ
gTOkKny72d/eszt1l8QSAF01+D9W9xIrSdSL136HQQ8s0bq3gMLaVcScY/oDjNNT
sZAcIJfgRi+Fpamb0zCAwT7EmNq3Wz8SWV+XfZ1b7LKm9PVNhumHX7JPJ8qIlQMh
chTnkK2H6x6IxW7zjnU1kZeT2Hh5puBnqUMhzz6oI8OvhHFRp6YTcLxnNYvjGBEF
RIVVEg435JYdIG0rBk/tBMu1nnaQiDB73ojqwR4wBCwKkQKIABxWuKV4iHRGctFR
ZfUBPcskLNec2gFuyMTr6/M0Vl9QR5siYk0OgNxCZXxSC4uelLN4wiGmL5YnkWZV
VFLrPtxPiJz9nAZtpM3VIIKVMzV1oNv3Z+dlUclUPAU4b6oZs8j0+VLPaS5RCSAs
YX+fumzjWndTadQCGg3kD7hCsSCOeTiHu3c/eMRB+qiAvt98qTZMQKaEv5mtSwVk
Ucn44N08MrbsY8OnRGIxLd5zaQUz0z7MXfVVtIOyHlCv7METnhfqH0/4qsXAJQSo
uvJEPlbBePng9Xu7AwUhwyU7uf7hypf/IAFdWfll7I5hqGr6ebLX/s7SyCad97Aa
ibOlRdQe5aq07qrkVh5j9iQUSDkcr5uDBgiVboyQ5/X+EXa8y14l0iqgyjv/s2GS
2mZEz2ZoHLS7yawy4JCR1M+3qwbgV+OuvGUwGlafa/wom7G3LiIb1aC3ua0EWnKO
yKXpXlk54knxsxKW4a1K1VOBCtKsUgHkdhC8x8ltlzUKdBP1Dye2ARpH2uyNen1j
WJITb1mjsqbBdN4AQIyvvhaPOqEfcKwE/SlZ2XY82wr9ju4DiekxWAK/H6Gj9d5J
kXiQT/3lCTulDcHduxkqHpjit863srAzftcewlc07pRLfELqTxB3LzMs5CjazoZP
Qs6YE224DU+yoZiIrRFmkANgjYjJjxXXxoiT5S702X41QO2uqA1sNX73zpsu4t0X
hm3d1xles/9Ib6/6IbowTw7PuF7IOMp98WoYkK7jRsXldFybwcT/l4WMlirQJAiT
q/SAyY8yw7kSWPKRTz6pApJgbzp0YRU46O005fEff8bCm+2E7c753J1IpbHelY47
n4qg4nrhjAULHXtr3zpuAxb/YFDO7o1l1GQJ5jpqQYy/eBn3aV0wygo12wDrWNg7
wOjIO71Zmj+HmSmaXv+pkMAcyIx4uNs6R20ggflURNCny2t2Nw1en/2oTu5SU7JC
7Ty6jyxyRt69xu9wYTf2507eCS5Qdut4okpatYougM3isjMNc/VyEUaJKib7lLU8
WqGZ2RswuuM8tuoB8E0A/HC2lBp1m7Jhdp3V8nlXtOssALzZvPqAx3GQ+whissEe
3x00IgdXemnvAMczrTl0nL/Q5Wrt8bk3U/XMe4JDqymBTRu7ju/H/PsiuZVb8Arw
/UBiOZ6OCZ3OWvvxduM99vw3L5iV+TcpxwHtlKbzasQT/qkmIRJuQ6sA3rcnJekY
RYi7cShJ1Bc71bVOgUbMaHJ7toFrIehvVqPqsKt5iFTKVpD+oJN7vtyaGns+dSrr
16GKmyDbBOQnIKLb+12obCuI93yY/G+7CzvFCg2Qwpw/4uqtPR4MZkhLQqg6hj4E
q1rxDnrbHxyxqAkoDRighmRngfPS0950ugL7H998+BegUrOmZSO7F9w3b97ef7E6
8Ynr0tfm5KvLWwS4BR24zzBOMLnTaAgaMLMe+nJMKFifpB2FmRXlSaWQnmvA+VCm
09Gk8IkSPqNOspMhod9PTmdnp+pOd6/MKbf2/+DVJh59pxZUBS5tsJreL6d/YvUO
+nGiX5+IxGaVLhCwYaqAjtOWQrrhe27/JLPTjpPuEGlmE6Ab7n/n9YM3Hk05ZRcG
LNAEE8fRbr/cF12Y8zQGF60y8wCe0rxCLRbIpvIQ3T7h8jDcLSEl78NspuZwqI/A
zMby3SV8fIP7EcZ67RBVz+6mrEjbL3rvcujF7AOfTlMWMcTmYVM6iYEluaYxFZi3
SyzgLGGqJBARn/1SFf252a1VsptovId4BknMH85GZEb6xJ9mRdQTH9Rp+wKs/Px4
9C9hxRHKop5klI3QAdnFdTHvAljIE8mRVk3v6sDnxU7xQESpFgRmjO7B2Gb9lxGi
hWFJBzPEEmISwkC/5b3mpt0Xqms8WMaRAs1c4rcBnZ4bWzXz45iyFMwo/PqJFYJk
Gb9aU8qKInvhS+RsSrjtW9/0tSRmvvrghO4c2rRA2W7vFauTXl3qg5ilz4nzvIQt
uoVbbEiwsDmU1sjuwR+OclJoF66wDp/hpp2tf5JVE5Ult6y/QcSwTN1T+0ya563F
DNHagZo7igCeg8GWsDw/8qlX8y7M4qEABJ58MXiE/LU/5actDNbNQRLagW3jg2lN
pEmhsTz2IVQ48fxszcrkWfwjqvb9Ijjvrp4tjsLWp49w7yfCWaZvrVt1wuJnW64m
399YYlnH5PpeOYVAFhjZdQ3g0LvOLksQrDLmqZPZjE0H1fjfJcl5QL/LOX3Klz8S
Wwk2TLZbqQNj6ro0nXyOxZUUv/dJf+DaOK/nZB7MDur7xqOBI09eBMM/nZErbymP
0WmB8p9dyCyacY8kNw5GuIqEovqicN9QbXR5Qo+TQv0+huN9ZqeLJl6WpsrW/XTy
zZtNf652343qvAoo1R5oDtg3jctKJdM8FETTt9FXdG2PUzghRdQG/XVTCzIOviem
ho+JNa4HqlB25QK2prAx30U3hDE5EkVlRlx96gBlBzXlU5XPohCfw1L1SociXGLt
w9sIJV4vFWQuc/Qih+UQHN6V6M7RV6sK9Mgv8rHspjvQDKa6Wzq/ihXC4Sc+hF1T
cwOxbTIHvP1dSjhEWL90WoozXsQP3CW6t84Q1zhoIXqfwdnNxhNahRM8tTTkZu/r
n53aSpTHImLySBVvG0AogekrIX8q3U7Bdz6mTroCBLmWB3V6MqEhUo985qCqadIt
EqKfn9dLjH6Fl+Ofjhun/tby++7Vprdl7VqvxNJbkoQvZW4JYxFgyGiqZ8/tZtwM
vFzq9DI55/ChyuFxcEhUYlJaP00JxcdHVbwiB3X5RiCumNjRq2lRrFlQehRM/sxg
7fkGMOkDnBaiv/86DQZYNhi6b7HEjY8DpPc09mivvuBUeC7OXSGMfKYojkg5gO8d
tPDIqEx1UUyqbV0jI5ET1TD8Wxd/74rabEvL77A1K13WN2xLY9scDLP3fbDiSDKj
Fbg6XUyrTjQ0hIXHLUt8LJ8LxfjFn5aKNokKNQtWfofnFZw63sHjQoJ8VLtIjP/O
AsnRIijNygf7FDh70TZg1c915It1mkI7o09D4laPCIoewYBsRbpQEKl89etqx5Be
g+Cv/5V1EiC75OqPoASwprU+Gvab1YSXZH2SSKDDcBdnBgbXqCVzkTjfuXoov6ps
9FD8NklkudInVj5ziKgxry/HCHtm85ccWLZaccY/wycL31OrG7AdaI62mzcDUF8R
yCWfns2sl93hEVzmya0nFrsZ7upWdjSkJ2cDCVNP4Z8iIaSKOE21aPE4xpacXkP0
NI8nkw0Tbhefy884uV19V/8O5/DQS7dMWE49Ym77F0aOa4y4jf54VgWKtZXeA0Tp
hc+x95Fc8EaRO6fE19DaNaJC2i6vvBynvUI3Ta6KIdjLXdkUWNagGp1NcGVFcG/+
LEKSpOn4HyIhQDumV/0QKktrBsp/OYduiSz/C4OX4k6rKCwPfRgYi78Kx6YM9KSL
HtTgdvILCq4PGFHrOztGa5VlZ3rkX6RE0XUnk7gAKC25FeyxyAfoncPWnTQtG1PC
Tk00Owb/9KP++R0VgAFGiVs8pFMJpe7dWSdjcmkIMUAVHqLet7SlduH2wvnyiCAb
u05Wg7Z1vd9LO2mMbs2dU463WS4Su/o0Vx+HcTD+KnadhPOGBSRyX7jSHEJyisex
2Ys7Eb0vMYZiH0xPCA5/1cjh32KJWYIeqHcVtLAPVQsBrAw5CQ2AuFsM77ogr4go
jOerqfG5st88W4mAdF467hTf5WPXFC9xrBo1KVLOTGNSjERq4oqsxNRbgHO86Zfo
/JJ1jwDSxMtKrNi8d2sDpM/REbVcS4pe31jW1wCWbOF2OCbzNk59bVZZK+Nr8rES
dg+uZLAIq+phJi09HpeV3r6C+/4QVuHsbPHFrIh92UD6u61+9bbnbnGLBdtwJTuN
GE5tQT/M0eV/o/dz5AU7HGewZxB+4Dpsnqd7dZ4OISLQgUfquZjd6Mpb0G1Zd41X
nwl+K9KI7jbNBHBHWOBkCGVQfACEvNUhADZlufGeFOrLyOPN6ATjeyh1s2CPPmgn
tE6q7uPBTLCV8imf1uFUGFgU93Fo29t8Is99m2uh8qagBAxyF/scLoLjiReMc0Dc
b0tBhZoJfiUQyQDzCix88HDfTQnWBXd5rk8kk0tK3NwHmMEyJQAmSN+IBKmcQ4s3
IINxyxLyQLX6BLfqZaoek4lmjGQnL8BsuA/nBnCNRbKDLSi6DzLR/df5BwHfv9V9
3B0lzqLXfTzwbFZ5G2iBqid3jzkQvwmcSmPzQFdYB2nvzaGbrQp969GoTzlusoXW
tkcMEAZoiRTjFnVUqDtJQ1yID6YMA5NkAj7Q5C700NNl2Oz2K5ZiMHf6tq/ClWZR
5YeQI7lrEfFqkyNuwVJ9aTeBpBNvm/Oa7V2ZnLa6mOsClyt3HrAmVnAojDYO+Nk6
VbIWRIJWu1rzWkaIo8toe2SK9Z3Iws950zMRFkHoP2bLfi0zN2vBwHhmFOjBbbf0
wDtP/xUp+HqkIjWJTWOzOb2GLL6pf46X9Rqqyzx52yugbUGrnqjhLg8VBATMaBqy
PL4SkG8nABZUh0Q+UT74eHp1N0LyxIE0SOBCpZ+H+73B6YEsxpmBjwtVK5cRpQC8
J4gpxoDaBSoFkUurh6amWueju9N941QylNLPQgDCPLZmvZtQ/BZRfiP4mITF+AeM
iv6cIJp503lZlpZ2lNJWKk+rRRPh8PfiyMgbcpc+3uAPZeqzBtZJBNBXuNMKLpRj
STseWO2oMN4C0VHYVubIkzgzHlghUVTdipDzTfVyp9XbjqdOwULi25uqhi5xH5pt
S61jG+IqGH2hgdKyaFl96ZUGZ/cUKTgm6opg7wSZm14c7Wwy91eTsD8RNqUMwW+w
/ml8zDBnAlwv9rde8U4bhvg+PRZsSVbfhHmMVG3YSki2VzSLz/iyZXOHKUOl/qhp
Hl1YiFaiB56DvOEoJNfxoUnyvaBNFzuhHysnrtQkGTM6lfUdslC5Y/KXj3qDjKhk
wukFLKTBWzuTHN1b3sMCo70vsBiic5xPs/w2vW+DYh7wN2AB18K2GeWwdW/RB6cN
JPXxIKBM1TP4ZKEGb5PgtMC4uRDZ+vbEfyaAUvvTOuu7kdMWwwIrAfeVbgxIagFn
V/qhpegHD5mDtsQhDf6+pHcchPATXt1yLCCSOhPR2AtpMtBjMvgffrxH4WCbr8Zl
ak69ZOYGTSmkzZ+5jkWR6yIMktf0ElZOkoveuvz113SFghl3etHqiheoXu5WrHe/
X6whmpTktY47K+yobZPqS3p8xJcKwm+RVZ/B0QohjSFzsYc46jfMknl4v1pOySgV
A7GQe72tsOYaZI8aiUzO8PwZhUS0CCxcAk9LoJS36lvS2qfrFLfd/kLT1Kf1coUk
KJRtiCE+q5GDNXcNj9dcRmoFGlX1keHh1qCSvz1AGL887letfJ1BLGHlMfmthgv0
qn5WaGSdxAIVCmmp0Nvoa7D1MW79zCqzOP3NXts5+ZOx5iBsa1RTsZyimfo1hpEr
7EyMImFoJeDrtHvDSEK93Qnzsx4h0ga93m3ZwLpZ3rXbs3QJ2wchyX3Zz8ZSLA6O
F2PRgeBb1iiq2rNzdDubeHWeO9ys/JInaxVn6N3jR1mtRndxhUC++uc8JhGFgfip
dy23Ec7ZCmbcYrlKnF6GS3wcwEGs5TOUm9o3ksqj45f2GCa8Cuatuw2zfPHsiSFY
+OjclKogSiMNhr8sHeZQNdczW8GnkhYujbnmY+hPdMNjLDLSsRhqocf9JbDIlktK
bVWKXFgzrnkGwlepFIhyhgElCWlPOhRtSz+TGl/0QMVnkO2dVYh5Ix83Ld5dPa3l
sRtBpzqLUf3GMAS+3C76ervi8MYIfSGgyAW67BPddDE1oH8GpcstZj0md/5rmkfB
H/T1MSCLlVbX5KVuaw3biTMTmm87hrcfsfO41kif/5sSFULt5e37RrAAP+2nZuIr
lKhe8NrZvFV52L4Abr/oboJgh/UbUa1wpmI9N9o1n4M2uH2PxmKnit/HNfOMYLgP
EKGn/LI1g/+208NpFh0O5Gw47h/gMrbHFKVviFYWqePCgwbTQRL6YUDQESyWY39b
BBA7jkaKYm4XIIutCVjOt1vsNKu/cR+p8CAIJy3tH9k/tzldV7FTx3DjvF5K8NLZ
f1sXUuCWPZwkSGtSC4NRJNpJs3XsknimdgSNOBCApV1uYb4AeAoc4MWWgvSs6mQV
YGh5kR4IZB/6PKR6sr0DMuzKJ1WZ8zQ3qg2Ie++nTqODvppkF8X6YF8G+/GfHzHb
tm3wUpIT6vb+G2wT3SdUke+pg1SHnHSp28nHgwoiyC+eg/bNGCi2Pw/j4M4O4nd8
Vx/0KWKK6tiBjhGNVAYTgOiPBeh9Jt8mQA6riQhrW9l8ObPBtn0zcmuLSRaGZWzl
Q7kni+XDLQJ94WSk8AbkfAkihjsdgACnbiFNbp5iURwGvpChOpGrKze3x+mGRUWe
d7adfy+QGqINyN35CqqVGE0+kvpzQvUHILwgXwB/8S6RL4j9SDyoqa818y62LQ/f
iPc/ZNX9xi1DqeVlp5I3h7uiZ7tZuRTVnylZqEwjmdZvcG/VQIZGKsjgruqCPGqs
CYs8wg0ooNzfxb000G5OZ3kO1NKu9uwU2oKNi6Jb81k2+KelhbpP80/7yQBeO29L
Z6qiCLDaOWmLjjRYAujSyw1zTfJ8rfOTHXRJh5ebc810Jfdc74Ybu++Vd38R4oB9
lWkTTjgnpuLH75ChfM7qBEBT3B/ROK8NDSRlqg24tO2Ggnp4GH/034yWJ16B1kPQ
PS/PQ9FOoZWpgnu3m+dIo3ZByBXSz+DLpJoFFURaa2V6qkm8brHhYPqJFHB6JkFL
ESekS28UJRrSIHkyd2WoBew9kjytPnc6X/FBawSnBTfvK3epvahzaBytNMDiMcUE
AzppXpqIlrHpLJ0hZJMobnOxi+f5IEjftbuOgq3tG10Nm4kwnjVBEROC2QD5xCH2
DrTfb8GY07KCnuC83fi8EYQdni2MzCA2XknYtW/oy3vpwWi+dLhNSuWwyCeGa7v9
wdrZ5NUYCVec0Gos0W8SpdhnDFB3btJkC+URskksKM4gzw7ItG1WjpewfwEIXzB5
DNSlpeSMWmCtLYRfDuGTjx7+Rf5mOm9EdyMzURspXBinLuqHtnZx9boYurtLtxsb
+9MUFmpBqvxEBelgVGUpyy7opz0ZqKyWlLE08Hw9I6qoP7Jt2sPVax77yEwOhTOh
5xrskNsoxTxf1ZHMA1XnaBKUFdXC3dQ9vidXIuhncmTqeGMWi6QZsv1zFaLVj+mj
NebySwtqxwiu0sS/5vtHIOW/ZpLwvgRubUhcpO6WWtqVDV3T9YsDxYdlopsnd8Ig
/rJVwDbv8ZJ+Pv8UyR3QWQLVnao2srbFknQMR9BVEYn7uo8yPdIzX8/ehbMUhcJM
vpzR2Q55HmZ2Qs3b//GDr1I4BtaxKXdeKtt+Jjs/f++/lnIcFfPoWvfP5a/A6K9q
X9Ev/VEwBKog4SqysR7mN06q7/aQzk+PMgcjflHKUORtDOZcYpDoanQNQk+/nvdc
pNS6aQhXVL3Di2DZnndpXqdGDgyK5qMYma0E7P5hjEOX/CBOHfmLONeaofhX65sl
4ApVTkrVZ4bJ8Dnr0jkfA9hGCAGF5kNofKLoO0iODN4HMnnuBizkgbCcbT3FpiR0
G4tf8jnfxjF+kj0fATUNddg2e8SRGEBvdLV/E1cMoFT/sc06EEXwTglXaWPoCLqk
Fn1AoWGxftiPeFzIOtFH6PZscdvr83VGrPfVOiPs9rjlTNkFBkMaYrFMQ8KMlU0/
zy1+kcZnuuqmAb9gjJA4SVwUhikBAIWsMpjlC5ObI9hdIBRk1xm2OhXNwEkJHWJl
IcpywAcVZ2sdSQgvdMb230vYhlmdkJNddMxYauBFCg2xqhpCv8Ib/bk83SXkgXLA
R1TvTdfZgA/hFRAoWa9MU+DXSb+MiGIIrK2I8o31LwioOhiTn6ey1M2/7rno2umx
nmrfqPK2vcrzysytWucFseELxoEtqPzqDCTuRo+Unbhxa5nBJs8EU2ugVqQZGHWC
BBQfUxOI81qcqz/i69q6AgrZ8ewYAHMALiqWO+3uKmOOiD5tvv70V6WEkHqpLsdY
kPBRbm+02ZoHAZESXga4dyOc8ieylHkm30dnfK0hQBVAwvjCm/haQvpe7cG4lpgo
n2OyOsKvXzSJfuTv/XHAveC3JgUslsNRENS1iAwrjDmoZJykkeSqe3lqLOVtalJL
Pi2V8sh7uA4WsTHBYskcVOn5G2UOHXB9s1R+zroK/Tag3D3Lxc5mm7eKTlMKefiV
2hDUB4Of2fjQdvoQgurrP565j06Q0Bt3bzLu2ayYJpKQs1XbxqY0iuC1eZnjZCw2
LQQMTOKbyw1qbHWr7FryZuTwpvYy5283aTtRPsprRfTIFQ50OtTYl2tQ55GECnL3
vPrdpiZEYCzor88dgJKFO3E8SYLa5aPG5AxErpqnZRgFYzQCLqe2UWLQmhHgL0Sd
bmBXvhk7aUQU6zjhHUBhdMq70tt6WnFipfgolhhrttv9uoESTL/hqziKweAOoLrE
1BHQpkNQGTBGbyMGCx6YpSjPep90KXr3b2gv/M74w0XWKzp5v8iVihB2oi4wEDIY
HOW0lileWMiR/ihlMkSqAhH16fsVj2g2U/vI8KpNOmcNOc6OgrmVnDNbcgk7Q0fT
K/zwnc8njGcCDtGEoyL2XrMapJGA/7R6D5u0JKl2zA6pdfBOeFYXHehbCj61OV9e
ptshH/UJlb+Tfm+idcuv8LKqGKrau9rNnHTfdJr+sMOt2rGwV/0+j9QaOAbRENGt
4eriGu/aSAvXgMz0ED6a5G48JjP8xvOyYGXQiZ0CzclvY75HvBF+VmZc644a0f9X
3Mb/dr2OxXqov4slKgWPa1hoOJE9AZn+XYwU2jlRQlwAEOh70aHcjK9MUUBkSncN
6PbXofyGkoWhkRJzigTMDfo9fOKIIWYMNnnCF7JXzZgcb1T6hPAeYwlIqRMk78WD
aPy/vJdo3EU1OsZHg5U7RRkHFMH0kNXF3NJ++LU9Glct7m5odyQdgtgS8NRWjpv/
18bErcpI486akT1LWSirQ96FCjIccxLD+NmW6ko1Rdn1E0DBwMymBQIsEUXCRVeW
diSprwoXCSR1YBRl6TGjkv7bK8Y0OaHWkkj858F7pfD5xQTpRW/D38gABuR10By2
aPybeKkk//CAAzn/FfN1xzfir99xtnc3Oqe4cBX4oV4KMVw0tfTt7i/4n6Ez03X3
O3UxgotUN6HtA1jbuNr0/A/VCpNBDL11v9BK/vyJFlTJvcnXjzgwBI5pyy6zYDkT
xrkeU39ZNqR6wSROItaosYCIvkj1yqfce0T3931wXnASrSnZQsoWuvz9xusFNyaX
jbtTirWWoanSsnkEGzOiDD8MBUUf+hkz30SBrjRpoQMHkTRigC2iYBWqLZyBm2P4
GMk58lYy641WKCfUVK0gdSaWZgcII5AjCneS0MJXGc3/J5+L6oW2+pMha04i2req
I8DpSu28t06qAoM/0fYQ/+w27UvcP8rFJl+/JgyDcjI7QqWyIjpUYsodYqw8R7e0
5UjLv0u2Eb0LPvnnR1AIjSVKQ8vV8PAUD2tzmYD3XYGX5QJm4e+9haySSplXWXoG
cFyAisLaDb7+KAoEc2d3k68oumpQTu7Ght8FVnczOlOgGYF3owJItqjCPencRZC3
6dAbNtSdycg+SBie/3SWWqojYk/nJSJYPoUwc8aBGrZX8XDswWWvS5DUB250AJjs
NhMmejq6+8AeQswhzzCLIOHJt9clBUF225czCqWfQMQlLwfKoD4hpiZIR0TQ3wyI
S/24Q5T8VjiVp1Agka7UyRk/SLbXPm2YEhGQPxuBY/wMN0t1McQABezr9WgT7ffF
wKQg5LQVwPp3tE2R3NU8+gy57UD9yN2c8+3KbcDEIVqtAdiFu4wZezjpJ7Y0iIm6
hkS5Mch9L5G+vumAONpsmjX/a0CKfihcyVUl+aKOaRsjZtAsFzpoDHc4PWCd9zWI
I61YFsfuRFoybbKIK4mH4I2yReVsP1x9L5ty6Nb8qUIOHg/m84rB8jD5PpMX//KH
+zr32BvzztqJt2JcYVjco8j6ftdCu6Rq198othOxoC6xHM6uuoVKL1vXDES9jhDd
NwhKiS5ZNjGft/90ZHf8dNPTyOzpB6k5lf4HD9l3USydaMawYFkEPatKpcTXc5TT
d9PUS3+obONJDU9hRe/kDAbVEMbJO+k1Idh6So5QefvZUb5xe8bkefJLwCe/VxVZ
0KjB6qXk3xDfnCCp5oHDYnjjHmGZEhI1CUwks76b9Kpg8pkNQglFONEgv/6uGYfi
2mec+HuZKq2CqMjhb1nxVIRoQiGhBtVAWMpAJ5y+euLU4PZ1N8ps6JKGkHdUtHcE
Lk4w+qxtb447aOuqxkhc4JvUmO1U+Q9kZGZ9pJlF1kzQMfwxt5/krpDzI3g8sgTt
X2TkPEM4DeB/uaipVq/3uMZ+vr67ZGB+3oYV89z+XNNCA/mFbYPAshkccyngYGZA
P6V69v+9QtnTRUbL7NLMaEtqpjwcr7febuXDLnjjNtR1Aa2wdlSa2z9iCorNwtQ/
evHHrlp2rmbEoy32MVYOvVl6CuGroxwWtW38ODszT3tex9DobqHmx87+hItFCHxR
hpcK+MElH3S4O/2mUfvOXI8K2+itb7F8rvBN+0z7QEzFkmuDBOtWuic7nxPkIZOC
HYniqCx+FilwcIG/Vy1OWog/hgRBZVdoMXAf0TpkFeW2cBMHf5ATD72nOinyIbF+
qJmyMNwDV0XbE8Z/S5wFPPR16xkOz6wbrXTXqTJx7lTqoZiaMex3As/PD7br8DjJ
naevvF35yBBayBALscS2n4iBODBaopamsF199Y/EnUv2CXRkG/hnxd0NtJBV36ms
gaMe1Lh31Mp84lxQMs+SnCmbh06oiFjrcGaeOK4aXD891+mVBiPmaRgBGUUQH1Jn
oMvye2tGisHs7ALWh7LB9nZkCCHAjvkbuUi8+9jKjloH0Lg3oCi27GqysQsuWEFy
089L/JPGT+mN3g9LLyDsNPyUhy5ooYOAN3deW0M+gXRjwpK3MYVjjoagXQNpGhc6
4tVXKUX2VIwJnIWFF2FbmT/Pr9CaLWNOtjNA7YjvunbS1gMn1VyAHbkxCYHkbf8y
1vil6KeFAXoc76F3JOf/s3AVCKQ4OIukKWo6m0ZHexIVMB0e14eAbaPXSvhff3Po
purBnF0agVjCzk3X43Ofc2I7GdejXHVFEN7iEhm+MaGJjzyjh042fLlk+r4a1tFt
r4+060CXLszicxaHDzn6oPBsgh8PLu18YBoTZI4Jtg+MeoGLQgJI1pi+ynVxzBXQ
DjkjtnokNeYEz9X2H21fU/XYi5YyFep/nyUf4ti/mWvuw60l+PeeaFU6xR1snb2L
3JSXjSCOaBgGu2ywvFMTGj39IHPwN/WRgrJ6YCe5cggShFZ29aD4BBrrfN3Jpcbb
XM04Vfg+n6VsPGA0eihL0OMWJ7VPu4/bVcdINgrsQGdHLrqHDZ9qVMfdYtX4+zhH
uJeVVb+yrZjvdpv3jslYnyTXksGfMH3Q7Ae5WsXG0AFvqaJoAy/Ndnh0i9pm0Nek
o4uI3VlsRFvKQAERN+1LjWR6aSIvPT4v33Rhwkh4UpVJ9nnSPYMAxSsaNFqqq+H4
D/eXZyVI9nvn9rpaF42Bxh5NWag19fI6p0tJVLw3zDoA4DVR6zMKaW4BeVD9xFgb
TYzAohobAd7MHKj/JjC/DgoIknb6WqguUIyLw1JlkOV83yyKomR+v0bMWfmna9Db
61/8EWJbupzLswI5dURAZzVAzf/r9rSRGcHtqatsLnPJuzgoJjd+Im6lnzydrbUE
FcI21u8BHvQqaVJVJX2gryDg8F1iLS6uaFfcB2IFGZ+N37UedAlZ0zctCn/P4YAf
67YmUKjRNQg8bvBArgGkTbRed+bc0s/NE5MDpJm0MaXQdd1gYd5lZqsOVUL3+3D7
jskh3FO+5lp0YLsaHT/CZvmNwA9zE9zozbyXNn1g0m0Ro/y+N+llzvS2eokQeaN/
okbgJVETTgVLwPsL3suiqSboECEUNdz9jLp4oenvhN8x8Jf70sAPBO/CY160jScf
Xf0kksasSZ9R6G3t+HGEYEUvBtcZLxDoel0cP7TAvQ1KPYHJnaHFVcr5woKMwib6
LwP5ISqZfutHgo/aZHaRm9FC2KE+AGLwAKO9JhSpRwrfBTyNdOK+16BQ8DUVOL5E
t2bsm8d+jcq8I0fYIbpZqei7y03JQvs/rNuU/GnZFeZkSi4yix4X9XVqmPQrSJZh
8bP6KymV6PwQFEDKZBOtzOVGd1Kbt0w/PGkSGrA3+eKhov3TcMnKZ3VD3Hv7x0Dp
+vLFOyIn7xUeOF5F/zpcyhYD6JnYOVaS3T5IgVcPQhQWcGo53SSUpVVFifUCqA+S
g+6J0OvlA80JeXl9G5T1pveYMZo7+oVfqhcBiY4kcrEU9inTNDUkEDS+1whiwyzO
FZUoPcIes6atpuULuY6Qz5zhoZ1CRbQJD0/hSl4xW8owuafxHOS01+pWhrAvJ0hT
H0fHKn1kbKS9p1itn7cuH3x1POiMRTPOZMuX8aXg/JsXUSG3B9bRIjeR94jMIE6u
qat/nKVnrnr3yVcsPwGmgJRzhsodZB+1Iyt58dBGfkMg4kjgItX/Efalso0DqD9F
S1BatTUpYw60Ev6eQzNv7vjmpaTCd+UkNkIJC9ShDUvYAltg+KzEnzE28+QQXbuU
LAn4cmoHUuY+0bvU3BnQv+cAH4qCgvm+5dZPt2N8cXexb0g2gylEX/8xRTpqxjSc
p5O/VonNqB0j0/HSEg9NOqSDprffpwTwA49Afm9DUKMY/vF3zpua49nWi3DLoXd+
T0bwg7EMFt8gVxC9dbpre8jX8v/wlenb/PJnNjbMpbxpysdqEZmNMkBYzvRr4bqd
lkrOCfPCfOJa1ncr41WVKjQ6FYF1fwEhK0eEcQxom51I0GrDvg6h8AaNDNaKC+hf
jWq4yylCfo/5+p92Tq1CBfBNVR/3JQoOKEIQx8Yme+a9+wGE4ZSehhVBgO3Ec+sz
xFJSbuv3eXDG4DFwgOIIAheGNA+bdh2w6i7ZqVaYhwNTjX6WYka9/D5sAnV1FACG
G5I4WrJlbZz8qM/A0mva/FU/E/rCKJnJ+4kgSBA7sifj7d/S+xuSFeo4BLVx6ILu
9p2lOoFx2E3wmuTR+bUGBcInH3mgba2ajA63Ms4Lq1j33p9c6pmsxg3fyZTM4/Px
8prR37rClN+yKulWBRK5J2cR4DvNGMkTMQzyo4XKKg1sAarTTmNTpxbAcmk12YOO
upKDt0O0F3VAgnfFhJk3eTVT/5uT2t7mymOmfolO99riEBgl4HOHQp0NdTJYZr2h
YSPX7ZUZQX2Dfi/3DQ/+VuHAtNa3qqMsISJy+++AOZrT5AahbDAZ5JybIeJnRuoO
ECOtPE3BcXhfZ8tQFas7j67nudWzNunpZN6ZoyAiBXmrzMMK8heRnduwO0XJzvyE
+Rs4FYi+wyFZOYZfQWCCV3/ifR0Gc6DibRP7Sdf9oDQPTyY5NjAJHdwVSVWSuAx8
jwK4m5jWG5SYJ0PySgtnzoCDouzQPiLKY5rlMIsyNfc6vLKoRJjgz/gkZJvY/CEp
KMJEpn6LxOHgOxUoVSU16Icki/f0/bhdlTylP2xBusJEWYxCghU8y3OtDCxAj7E2
1o9Za7kPh7utJF5Q3/2NJbVNkJXbSD4QM2Rp8fh7xuwOG/u56yDiLSMGL+S5klWy
6sooM6yEm/DB0UJt9Akvk3t1gPtqazXlOfQ8HlElc8Ec8fgLyTm1jnsZWbMfEAMu
Ifp2BixNyaXMM/RtwOLItEBtd5Fm9UZBGW/QiaY647xfOQyBd8y1LbIDos/EYnQx
P07980hiSFG1adDE9fqKEgCyUdaxpVQuFUCt5akdFoIb8Rzs5SYmEUiGVjk6Yf28
3mBdACIES490GbQoxeKTJ1fuMrsbUprHp0r2NyLMe/JA2TIOHFe9LxaJGSIhuJ99
n5UA6TI4C0kGvjFcW1frRaSjgLdGYu/QNDUXN7XpX7Mj0oYRZoKJs9Vgfv7MUcrd
5Yj6edlscBZQIL0BG7qUvzhH+jzQUTYw0m//NL0Lukz1vYkpHBBTozpNLAh2vsdv
1P8+AVGN0VuMJzPQkWL6HcfQ0H4hq0+d7jmi01/wONuAiJUk4wWuuU3lxTRH8L0w
QJ3kbFwT3k0kA60/JNUxZ9kFUe9z1VYsgEW4VWf+CIp5dH/LT4QhQZT8EK9AFQnm
9CmaLvmB25avk3bg5dyNlpCMi7ZW88nOwrMVpheuOQmaJ/LxXfgcBzar/ny7etiW
QDM6BYXFQWc/7QM/H4/myP0Oxj2tZNlV96JZyZfMOjweA8OVpXoRsY/0nIIzOfhQ
uRRHQibh8n5gVD4b3z4+iaEuCaP11Vri60jckYA0VyPQ0WR+FeCf62JT8JQZrOE+
CzdniW8UvkeWBAiGm5ucrruvcGNYOgzselRRtqzpYkoHrZ2Wvpuj9bYoDYNAFohH
bLNgopOZesxQLNsEsnDHHtxT3RLYMPiYra/N2PhpM4muYZYrdzycyuRCWe9XlqMC
Wa+AG62nPVn01KnUJXSq3xwyRjHn+0RVxyfUgVd72auPKXG4UCNiRT7ozPWEO7PZ
Tg+p+eTxxUZidkuqaVUjp7I0r/xl5Br2cmC1SLMaYM/8DXNhxSxBtEug5sdiL5lF
iCMfpKXC/n/e56AXpadTWT0vtNmpVdpq9PNhHcyYHmbT6NbJjeSlQ6FmYQpkPNMi
mPVBDJnADNNc32kZTeW0qQp7nxMrNuQ9NTwgFsnEz20Wu/D8GDpdLB1nfPeoUQpd
KzZRJcTnG6IbRyMT283chUAK7d8dm1S3sSMmTYM/oFw49yerMd8K5v/hGDkIljoC
lSsO7cgan/sYvwFWH8QrdMP05m54IZr9iz40xnK6iW+fG5gaTIp3nIL018FS22Uf
Dk9pU5iBxw7tIasVbt/MR4zt/kiuOk4jQFBJYVqZu/BpWulalbMIfz7hVVTuQpw3
xzSysRZqdPS8u9Bu7qPbOOFtfP/EYIo8UsWbMd0iGHZkwnkEpj8qehgknLGHOq1k
AZwX3PzxGN9s09oHERk6pL+g6iocWiVdjzeQ9oeM4E27K/Na2B8NzxIC+JrLeA6N
amyKjugJrwWt0oh7l96ubS2u40Ikh5HFb8S75miQWqTNRR4xH/FlqFsRckcByoqw
n4Vfx/XLJ0I7TpwD7kig8lVLzTZdBPsN7YNGzAyQ7ZrW/chvzU6grJnsv6r49lwE
OzG63Vtlva0VbwxWPSKurLQM6S3mGERLgScVhHY7wWICu5xFiRlGNpR8pnCs0ycc
bMd86ZnPjULGJRPZiI1MSX6H8+NTdJf0fvs6MRy9tDVg+0aqEiIZABfXsq6H28Sv
lYoypY2J/8lisubchYXYM9j28P2RnESXtsduEtDVZfpl2BKIcaTFmdtl+F/y1jeT
6ekJ4xrfTna8xuuOz+RA2xGR2xPdOgX6kn5pyJaObFIXUUQzPv81hiXu2r79KlRV
2xBnuLKGG+iVcuJ/fkV3NXIAjsM8hraovCGqDV3rDSAESqdg/+NtOPvRlfWOuWZC
CssyJOKVGmWq8NsIsW26AYJJJwc+E4NDyfFNjPfgmapZq7jKmcQoA3m8rwbGZIS6
elg5SrJ+OD8Hx4cYLYM1b6JLuWUuYuj/AQzPNeGNs2kDXb043/Yp/Na9YnPh3rGe
KA4svPXz1VWvnA09C1y253vXP+n9LVy0w2PsazBIJucV6dshP/L2ouePMWKfo2+6
Ag4N3YYKupjj/oextho13F7QGuGfDaNq7/vDhwwwkL0jolY70LjvjKX+sEENB1Tf
zfyiuSgrKz1J/oWXgGxjoaXc5CWzIuDMiaFhRCWBDup2HG8iCv5Q+qCnJOzSaWMr
jSdy+3zSjqCAY0vx8p2l+sDVFhcvny5nIM0shPpmO02iSGi02/wjV3K5i5/AKFWq
xXvKVUQt40ls7N2bzsoICeKE1Fj1PiiSY8IpHo6LHBpBFZf0PpScw5ntE5JC1JVR
xdXPaS5rXE+Et8fDUVnAAgog4O8whZPcIwkBXnWsytK7AHg8EemKMgOGZ3l1op6J
awrYEWJHDPAS+hKzGykq7LTp5Iq/uAXBeNiht50FU2EJbQg1y2FUVroc06bQgMPv
QMQkZOKcy5K71rlO8m4kWWS2Szo8EXXvIo8jkIDKaIZiXiOnF4lDdmsjDQ2Kad+E
zTnogZmcccRCMhFoE/eWbPuyc8J9jMG3IymVDmXxFKJLZpX/VsPRbkMZ238u0mZf
OdZrASEqAvZhal92J39Wo1qdz99iah8+zXhsJcw8e6G+4Ods334hvgX/7TCoEOwn
9y5Px+sJvZWDqwtJxY8v4wmtkyfJFUnvaiArKe60RQVeTfSgpXMJ2wY/UdJkWQ/8
kRTWYuMI4kf06xniFiVg8vLus5M468zdqZi+DSUIfJCUGDhOqHvobLaMKUrV14ZA
oHQx0RddWK/xpQKbUdBPcS1dw+0KNs/Gh/lnZpJlHBL22r/TXxbzZCh79mnAVgr6
t3Z4fM0gbF1aDaEI4LhdSsCwPxRsG1tQnxo8YNxEhSGkjYtPjL8kUMgti3S1W3eg
UeR52zyfbuC84CjU5pHrg5+s5DYTubd3ppiXaHF7aRV/e5W8XLo3Y/hB+/RriHFA
WldA5XPYtxBynPLfv2Kb8Yl2ovuvO/EH3Hf8MvOETGVgehab+quOoGnU4pWzn9jP
NrekP/qyyfBwg1X00sDiWhAcJqkak5M1nHqhW6cENChCpdL66TPVXWsHwM2C5TXh
eaCKEXTa+Y/DF8zFFXeKvxZYCQLAk9c6S7WQTPMWKL2pnx3B1RxqKAhAQgSSCB8+
G+rwly3lX2sp1V/dLMYrIyqCWYAOQJLnJh0L3mqDajRzw2LEdA/JiqlLpQInueav
S5O4/ELnrFcmtU6ycvL4hgXQEY+mJ3mCXYoLS4swSaHr4EJJ9hxxnqPGJtJAyy65
DikDLU1ixLBOkkzIJAeF5mPNgDn95CzhuCEXbwuaRZpSHAMcGhg3cS29lyeK8o0I
uUrqoqzLJFOMsMN3Q3/OmVn15+EY+zutoG3qFssGv+p0XYJNOvzCfQduH9iCkiKX
rSWA1Bt1be7XtpCDOjv/lrYje04GPj7xjcJuTqPWh8nM8BzT8DKEfR8hywvl9/k4
orI1nSsaalpXo273dZE3foOrtSgC5l4cJoQH7joeDSLbNZ6QXEbtOYZbbTkh9VEF
pS1ENvzmYm52z+KxX+ommur1eTWjOIEUix9i8PFblMhWFwVG0zkXz0doCL8OB8Be
V7uR0glfwx/n47iTGPTmAj3l5KJrFvtoLadec87x1NTGgGNtuxHK4maRlNq5C1aU
JLCK/tNDaaqDBvWlX7GM4ddAHeVDx2E+EdKRm5QJyuD4f2IVkcyTxjCOgpON1AMy
VgLZ974oyRCnZUrRYTCdiNNmj1xijCNZCPd+reLEpwJDqytuCz2bmt62rcDo5oxm
dUzjhuwOKP2QDEKI795zL8caqJ/HqApWV+ylxpBof448s+lxuJYUXVvj7p2PiDo8
nEKHEIO8eZubIDr2P/Es/LewE6plz6fwnsDTMKn3FUrIqcqc/r0iYKseO8CCucwY
LANT89piSWlSK0DN1Y1DMxKIVorR1kMJhoWaTre8RLWa7btLWz5NQYdeiBpiw8OV
KIoQC7RrDj8RnQwxShJmiz+HjJtr8k57YbUWiuMms2LOjrCfl5Oe+SkFrFZG0v/w
M9BYDKVrci1lhuhk6kd+iAJZbP294C3eAgmC1OpZd5hTWF8Vkx2zesbQihyHKBpx
y1/UUGA1Cui6PXw12KkemNbTOhi+L4lf+cHT86zAeX8Z7s8tau14ucr9a2ZkRnQC
r5ScwPnHVGO90PLW56nWyewtOxQFEGTEerhlRl+qt2a1TJPaXQ5asus+QiCyNQQj
1NgQ42t1axlqzh70wZeHUEVjwmztEvV67bu0xVVUbNkiSYhnQG7nTPuwecLcLmVS
QdjaZrZ3/k7bnKV+OYCvTMEHAsRKztkWL+TtJX1M9ljwhK8c2INkUSvTXPDtuqDp
99T/jNdVpmNd/YL3w7wDiAZTNtedj8fKE/DK5UOZJNx6CapS0xU7JdbFtGVjWFgJ
L7gYja9F2nO4UkKx8rWTuwyaSmyWdzlbtb8csiybDoMFp+NvxVmtdgTIRreaYqUB
NZkjgMUwooERB6jBKWbBzsaEAIA1wvx2+XBd3xqfkiaFV3b3B1a9jNcefk/JVaB/
+1WWhFOHaNqjl2vD9/ZPiWB2o/hrlBefYS4MrTLUBzsHH2FfX0CVtviLouMDNp+k
hm4HHuEp6maYTCSm6tFpbNXxBSfZAvb6nCXGZb76PeZWcGJN6fUbfKlGYI8F6zH0
YG/5ic0U9GwHxRApTBgcnmVZJdxfAq+vNllf5+Kz9JLmkoTuGVOcidlDJzV/NKOV
uh42pwFow5SusWzI4Ys6rg4bD7bNr00m1PfJkejOlSSSFtXtt/x46qJVMe2XFmT7
9j6QA18p7WS/IyHyvq+pBKdEoGgQ0aVHOPyOIR+BXAlMT4nl681P1oVreYoWl9lq
00c+NYhlv1kFw/zfF4k3ieDNvintEtKmPmDixwhlNAQqMWTVQR6P2xyBld6a+sRz
gPliJCWUlHavS39SAHWw4IZXFxVhfS+ybP0FjxmXMfg0Pu4ALdPlmxmFQyEbRMVY
FToF8jLtUS9dF6rMT7oNuzQErCZOzW4LnF7R3SxgidZhDSPZ+C13b8e9RZpofVYG
gTapMPDkyDCH5XTYKEF0MhTCJiSZ/Kv3JdNoOsy59sX4tvSyJC+Xh8aUhvbyjUHm
0rLQJQlJkeVMTinD0jFgp3e12ttbS74Xpd+lT4nieUmlx7uGAVsNYmkU3pHM9bPc
ZhbsQBxMGd653474RhN+XVPbkuIN5sp+jDkNevDkRwZvrBg92G3oteKTut0OLhHO
FFJJHsY/hwxHdR+FVG9B0MBWfxmg+UV/IvZc29a5BCkPMsrN0FIHHc66hxRzxNZv
3kqTntcBeG+wU5h2GrFMXeGEPQjICUbbHgrvWybB6Ria9twrzSEgAHdBmArh5eS2
nspr4YRgK02AfdzVaYXV0OKhNHTRnxoKvmvJagGCXD6fvkaBymPxtWn2+GBLkrKd
cI6K85tfYUMF6jFmYg51Dl5gdWFvrMeRRsSmlP4AWsMICa3fZHPoTMtxUeT9p2tb
3yKZxi29RbwtMTCHkb3gS/U/kbOUDGOedhmDI7vfHIgI79oQzH6bViBM4ccvYfng
s2xWjwZXYHKcMUGJ7+Z5fqd3g0YELZLzRRy+IlaZb5rGw6lIDXvNzXv41NlaRwmL
zxKVAt+s1dPifo2ZZqgdE9yabJRTmUXcNC3hbXM3n0KUnnf2pGxNV0jTx+nRXDgZ
CPD0VVdbHtnq02BvM/GmdQS0VN2Zylj1Z0z8q+AIKCkFTA20JU/454GwpbQ6BWaq
Ot0rgv7/oM4h0INq3E/xnfUZ1dsB/bHVdxkQgtEDgRsBAnk2xgY03ln6kOmhU12V
8bBquxAoxA3Ylp2Ya/YGjvccP0Rucu6f8wR6dIESvjUv+TT0aWsBo+iFXDM2oFeN
q98AH46uZKA1m0zS/7M8FXw5h0WVOZJ/E3xtEe8on+W5CWDTVYsQHrNhV6ZkJ5xP
1HQfuOZz22kfqYi0MMB/wsn1xViBdQeBKVtb6E/le1+oMwh/rZTZ1CMETO8Qc4iN
b4DiiWEDsl4skwNV28QN5S2AmKT9R2HyotWUQ8mWSAUw5qhYyoivTX7hbZp7Xhgw
a4sZQRdelcX5vF6TZ1vDe1QjipREqKT+V8tAlhHFWXNKlLxTm+A/S292we5ZdjQW
FhjQayxmR0iaaCSW7dHkpbtciZjsGJFVKKVjK87HkGsGKQ84Q62D4i4im8mxo04O
sdJvyG2qD3xSLyi7SUdCQrnXNrT58ghfL4yRmZHxkk76RRnyLCkhd5QWJbvbWdAR
NDmyMW1dO27ZU9g5IXaztuO6JQosJcsN1YNSJHaj6CEMUzt2dp+DEUHUW/HphNjY
IR7vx3E/srXXfErgUpom6xZ+BMiZ1RhZqehmWnPNTFx4735hgty58G0B2aQ1cHRO
cbuhPwzm4BPvCwOpiOmQSb/6QoQZhgG7ES4MVA7RLqsax8qRHGNsmRl9AdDTchnY
rFDEhPyMf8FVUecC+0y0gkjCU0qnqP+9r451bguLzSteBbHFl3tRahFlVOMThLIL
3/uwpLLAc3gAhKfWRTXfPduj4nkgEPkiJkfL+wZMNujktfU3U1Kl+5hKFmdj6ZfQ
l66wSEEppsrBUpLwbTlA0eDsVxsHpPpjMAQQVjMq02IY/YXDKAWrHvF82HQOQfqU
gZrgp8/tY+1AEGICnt/9oLQHHRx6UJDHHXfW13tvkUrpmV/mhzX53EWJ5elxhLJl
3P6ysvx7O4ZE8Jqh7KX67HKFODurTC5VT31q8+e+XIhibD5pd1GVeJxGZDWolk8G
3l3TOJ1QbVJLqnanqxZLelFpoZ1euirgB6yDTIfdoKhm1a1Dr29O7J6R5sUBWmoH
6y+LZoI+SowdEiXQBTXfPy20kHwdZtl7BuZ77Y4Hln61Ct5zM7nLl8GTmPv/ie8L
fOrT+HOnLvZ6nI/SWSOdavj3V+EQAq423TeTaG7s11bw6XGM/37/EMu7HzMbuP2n
r4hD0jhjPxpLWkFUcmEamTVirLYJtwH/FkUXIfw13FB1L3HmniyIcN/uwgA63Z4M
onL+h2ZLEBJ7rMXkBOFdfvxpVPJ4+0AlxJ9Ek9k1txftjtB78YNcnw6yCFAjgkzl
sbFa0P6XNnCxGx0smcqEKYT2bM8udViHGlp/QtWHyzUkVvsGRQ8tVJQCGOXM3s8H
GMyqblVFwijs2dVlsXC+snIOarq2its4Q6wyXwPjmfd4N34N/wCFVeUoaDHCbuKJ
ZbsDqqpmaJRsb42nso9ApB+M2QWZS+hvGZZSG88zgKq8oTrtjYAkNctAUQ2txoHz
+COoeM/BrRM4q+bjYwrLwYlYhru3MoOMVefrOa53c7SfcbUf758lEGED8JMoKs/M
xL+Duwi/EJV67GI/FtA48DyKItTZRx8oZtYsB73m13VSTroGyf2PhfSlOxTfHams
RsrqIgI8eg6mWW28txHyqv038Ga+yuZPW2YTquTT8i8OC+n23djRUrtTYed+Xysg
C04afCjVasdClQMA2drQb50sfc6Gs9cHioJjimgAMHVRrIZzTwDQvJcWzkWx62h0
2gpIeEScAmrqut3K280C+7KRWdeVTVDuge8CfPquIbUnlZ2+wl0Ry6jGiNV/qa71
UovlMqJXzJs13AbWZc52UqM09LIOh6VEM+6hl7Ve3Ma1+Ah7OPajui+w9N8WyDtu
jRPZK1gUHkMW9QiEq4aZDlgVGBpkM3NMaMPo4Pn3tFYP50KQufEAYuYIXqaiF/Xo
zjed5iKKx2GGBJGCQaH5DSYiGx7q/L2KQYbw9pXi7StNH1pFFND/pbuYf8YJZa8M
vPjwbaQ1g4eFQD52iA8vVLsE7oZPNb6t28D6AHB9IQFCKZnxsxsoTxn5ecSoQQqM
NXqzpurHFde94/PSqrYNNTP5DhYFzwBHn9UfRxcvs4kEZBh6FCfv/v2UmnXGJhMt
lL0sFlFbzw3UiPZdwoXZXmXcxq2DQBBAunssNvPLVV/knIAW9yoEf2CMx40gk/qN
x2j90WdM13DpG/mGi27XwnIAQK6X9cs/Kke7Pik2gZgA25mKLyf86unqFP3m1Nan
5Tk+c1dpuHaa5/i7Bdmjml+52LpOD/e0/DCGB8Q3q2NLhUwBTpHZjrNxsMwRixID
e3YQJ1i+jK8z4gMB3XO6ibslntAhb1/Al+TL6s4CpdJviyrZ3hzGEBmSpMnMhNLi
jx65wg11t/DsplsiuVQxz0t85jUv6vHPcKLxzY/KG6qVl4j8QdCsaZrguBO4XR1U
+37yEaiKfpm9tjm5jkCI+l9f+T4tvjsXhDyY9E9rZUkQ8RnIILfJ2fhH+a0FUODB
2r6D+ZXaBrbePpE34W9UfMXdFw9OWSHxhd3i3NXwW0NhSccXcu1PgUQo0svjIEyJ
JCwk6iWUsQ6rN8zMLuXF9MhEdxw7kiuKj7BYTYBTyFgyNy8Mynvu1Eb/uwNj59N4
LBATBOoM4nscHIe60LOxvogEqQCHY9s1EyVzg86rvXifoFxFTwrWIQQIWmgwVLMK
hdcvxv1bGMOyzzkQP+xF8xkLS07Czqjl0tdx2d2T1mdW0Qv/EqNRss0yIoqJT/m3
XiPs8g2gtyEvgS1vQlH/PSVMpNZX5DTxRcoOEEg7/M6lqAUmtgX7gLsgUYknRJQ3
TlSiX5ISuY7yDntrn0Gxzwz8WLX7J40cDK4FgKh5ATqBwrDkSTKjPJg7hdFEMmba
F+lxbUmzhVtYveIWi88RIRnDEwmq/AJ+sy3WqKh6su3pqJEzYDYwFGKNe8gaX9rg
IwJidnrHQabONlw65mjIDhfLz5FJ2DMzNv0IGOLtNiUd88J4O/iEQVCWbFusL5bE
oRRQtnJPXImoaN7EEmjDzXmKAl4/eskcHSA6RW5CROvDziA64sfowENVNFbQRWvO
fRXuvqBR08K8mpLVXTSryoz2QVyFPLNhyTi3wHQfe5wFQ2uLXWTR1PpXkvrAM81Q
/GmE6ieYX9+MmdjUomvE4TviYAe4DgIbeEcSmcBRRxfa+sFhLjl8UeBTGebr55Yw
MIQIhtI8D0nsuteBLF+HVVBjHxUwwJKVLdKHrtDqvC1zawOCgegM3mpUs1/pJ3xA
7akQrmifbyQUrosfEo2vyCV+/whstEBpbntY3mKLrKivoaE9WOo0d9Rgo0OQydyP
ZYarO8sETedr6jQuaXYlD68JsQxrJ3o2LCkXyfPpzstAxEom425f9WDR/UCWn522
fUlPnKIaQKCmWog/aGTcdQIpFV2C2SNSpkKdZ/oklZ+///Tlh3Du0PnwFDZT8tW8
f0Dcww8FOFariB4bZMPsOde8llwhDG03aXKjHP9jANEQqL2yDy/kbIq5oJS6x5ws
Tq7jEC24P9D9j4RW30YhnSuNhtQEtT+kjcwGuxhRsqc9J/t77TGeiayMP18SHB0S
/ckVoErQGMH/2Epr6xm6Fow44SJTRlewQgD1c18T3Tc=
`protect end_protected