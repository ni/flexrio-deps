`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12160 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
dnVBOIGMhMFpJZXzCENQ2C4zQeA7ThBtRChFyTpiOgJKNq6vcOeLPzEpmpIMYSUY
tv3KHMo9Pq0cEyDnP8TYFz+VKc8b1NG3smxW/gEYwBngSFRXzB1cF+ZPIuKcfuzX
yuk6jFksVDkvPAQAfD8+hHCdin+VQCiiq6UE0jve6uxK7H67i005+dh+mf5LmzZW
LVIfLBfmKIbsBwUSuhm2iDj+m8rLOyjeGEDeF/FJTrCHOaDjcws1mnDRd7px53mK
4Ot8wBhUS6cHQqbbrbTvBopSkJefvLxP8k1IKs2cXcdA1UT9tW8tsLgVGMUijtdJ
9cxu3igY1bnX+SkCyYIc8KwPSElGX6NZADTZI7zkdZbwnZg3wNHySkL7Tzi8/NXT
QJE+zcZXOa2JSrg2PkGKP35/o0tJY3vsaBCdRioMXN0RGQL87uLERSvqV2S6TQFL
W33cueSJ5bHiFzj9xj4sdQc7K0+nn1jds1BVIcOfCbyhCk4sOuh3B9NKUD3kted8
Y1r+lICkwrycg1Py3xozSKSXnCsdFItnS77F5ebsMqXJQGAzS1bJqY5RDQ4cFpYB
RxOOxVtPcx2QttBXjsHm0cNW9oMT3z5bQakXIK+82ahBbdxdiBCsEfHOhNcLozhj
j46oQ4EvkGXAPWb5lzwwDBXoS//LDaRxOD4dNSgj9fvE/GRGJVUxhB9jOk5Y1CuC
+IcXBVFTR1oXs0TUCMwkUC65W46iwkSzhQph1Ols2FZjnPrX6rgiIMG1IV0gb17l
T3z+YOB+YX2k31Zc4Q0+RdCtKU8Wdp/sL8ajTuRyP+Wa9fXpnRTVSvdMue/nXuP0
/ZLYopMf2O3d6x/oHlc3S1g5GqWZoa5UnSFnavp6ZlcK5Yd3En9gIvCNprqKjG2O
evVuQe6gd66qViIy63PDMRO2CJKahTBB+UGExGGc3MGxTIrb548DzypFV82UkXnO
vvF9LIRuGxss8z6+6n2MEVFxCeBIJFFAmc2dQ7ap6fk3b9n5copVNPAJQisrLIiA
sgzKdma133n5OPEB7MMmY86G/9oxfsR+sZu44JFkxew20L7V65aCh6Vtoi0dbuPa
MMQ0ZGW1czYXEijfqnum24owiOG67+gJbbg0BfRA/oefUe55Wddg0tBlBUpGctvS
l7Gytcfb4pf8ce2UoFYu/YkJHHCs1vTS+Irosbxdgyu9M2pDODsynH9BZvxmG9zr
BzNBUxMafMRbzepqEym1Rs9TXybwa1sd9eeNrljgvtmQzCdJ1bFX44Zx5ac1MJ+P
LD3a6QbXsFGWNLX+eDlbhn7OEsmKfxKVrrY40pAmQBE5yKkNZttmJk+EtT4JX4XQ
45FyOrgziR2afdH9vmJYwF5C8f7nSA1TvR2aZzoDY0dVUT7ZOTmwHF1t9BCEVIXB
bwk+c3Lmm3Pm1UHaSPqcA3teKDZry7MsyPWQ02DJwm+wzr3VAhPITdT7lY5b6/gC
c5rU/KPqKOj+veJaPSxsS/ZIW0C5fZpxlrIK1yJdb4H4VcvTSXvt4XJc7WoFYg1T
HsZ797WRVi9agFUip/tGc6I02GP3kPMe1K5JaqUQHUObUYV6wp7jf56MRWN6Neba
ylaSqMSI7TuKvQQXplI6gsfXm3v5aYoRJfRL6RV3D4gN22TdWD+6b6L0Kfh8aIGe
HU03LIbxwuPkBaxiasMuIcIQJtwX4DIh2YupHuvPJs0h5c3hqsx/m5j/p1hVedIS
6PQ/kOn1yAJzuWg4WyOP7ltBcXyvmN2opQBc4eLhgPsH95q4LzwKJSlAIe5V7Hv7
qTG9WSU/rSrlw4rcsSSS5YC/HNSxw+bD5qCIlKHia2mKayHWmX/4QrBRhlZwk3Nb
YYsJ4N98OQxNuQ7GNGLbZ4BmmIie0q77wfeo3pgh20YdeyVZ8eapgD9iSFOc8iQn
NdCFplgqphnkupX7D/1lZuYy8nmXdCAGSC6fqiFJfmK1RW0wkCP1hPdEFqT9XxMg
VbAXzLobEtw+brHFiPdg1/+CDVHC20ruUYm/kD2v2edSn1n1y5Eg0Jvw0j/iXJMD
6I55Pb95vfgxWiPo3b8MickOLJt4Hnv5TJJoKIS1kVvewVttD9IJCn+J9+gCc8HS
p8ITqWD9lKuO7SQIrxTJqPmUa1H4G0cJMxn/Bm//u0BRkHNZeWkOY7IVSTuaGe0+
oiFv2U0f6MfO8JKP8J+Vg9yXxhhx6PVitXBki3HsiEOT2QoaLxn2Vzkr79Lgx+Uh
6Py84n5lGzmsgFaTspH3vtl3dcjLV+WvA2RLj9ryw1ADziWcYLSopOOFfNBRUEKa
2jM4toBEoR/Uy6HY/O3KhCvYUgi2X34MZpeGlFrnWii2NSVQClYRnlw1S8qhfWD7
s6ucRMrINe/ozLvhiwDUCV4AG9pwafe08+UwL5j8TyBXylbAJMBPsSuMOrH5nj/y
ANhDADXMZBhHt9ipjRQVQ5Q9I3G9LWVjCZUPmDLG1uOm0LrsPQ38BhcaQ2qq/s5w
ku47ON7eCpWv0/5GCil9ZEJNbqwwrqbD5V/LLshAvsqhZ9cV5K+sHMQF+D22XtAY
uOKO8HAi6SBgOP26bzarp1w4efwzk+6Rpm5yx6rnG5gsSlth6rtxQ+CAk9S7nvrD
TEjQtCtj9X+rDuSpOLaX1tEegoADU9Q3CS7aTiEkCZvpyO+K5cUJwYbjU5ku91Xu
uaCtcMU6QL/wYG0YB7ZV03o1JDYrnjrmdeQEGf82b4+Fs+uamxXmPeivl00YxBpu
W2jmN9Kxzct1liE+nPkiggR3agL8qILpTNdjpdRwWQypVQqAF9awmTUILGQwAzEo
8fwLXnUPfHe1NFRQg8v9XkmCMLdMESUTt37/LwOfM8+bwZWl+ix+tPizj5ob0kyy
JAqQ9d1JKzfNLQz0D4pkxc/cDkCP97t5lTTS65cnwVlN+4zqDh9PPtwTLDy6Iiid
CztMEeknU6cGLe9w32kLGlDo0CexuVxGqhirNc6xZ5k9xsYJjqXL5ncioBostKCm
YkMIWyY3QQyq9DujAnO4fpAkFsXy0++//uTg4xLC5uF5wnc0bD+asLthh0XP6xY6
8XX6m9mSWww1tC6/Cdnb6sFcTI5NP9Z2nhVFjep1aL/7YiKZk9csrZokjeakFLVV
C0r3PZf6QROBGzzrXilzPoNehDmywDa01xQhBQXkHGQqI68UA9P2SiA8IDPUGqtf
lc58j9PW2CAF5SWDIaklZQg4e8IRchPqKzfDqClwfSsJITZZutn9hW0lAsUfDxB/
1bKuxrgGwUvCACz5KBVy/1sIPvZ6oHIlxOYO63yV3eNOFZayhyYyFMGyS7Lmjkai
gx7irOQdbRYGjf5lpB+1VX2PB5RVvwRz0yBYsNPQxdOmht5W54nNi24CuuP2z2NJ
xPJFSm5/LG0ahPaiO9WHdHQo9uKWKpO1GWdpkfLMTWVm+Rl4lJW0JPmAkDPGh8av
uKog57F4e79H9vgwUfIZHJyi+pZ6/INqtnULIr84eq6hqutl+ztGmYFDhXB/XAr5
ax4re96fUa05I95A21S/h3vkvPkif2v7dHFFkG5Ez/11bSjg8/iGP6jIG4eYWhed
e802s8JcfcIy3tg7PrLhdZsJ1geW6alkUzc6cD2jUIEb7oLevNXzvzbbqRlcJvWg
xZiPQ3poQFmUUMMyVSs5Un4LHPFRRWk/65UCKaR6YvN1lecc8hZZ+ZvBzM4omP9k
UJeAi8mZZVguIbhuWR+NRp2ql807lqUtr5IobZJ7wTsBY+iogch7t8XyHa660a7y
RXJTct28oRmgfCeReCGtDPGw0SVYy5cN6vI94C5PyvvO+kh+GM9Gm3gFz5j1u3gM
65hldGT6tF7APtFwmDklX7YLMixCneys1lfRzj1cIJKn4AgfSps5eUdH0p8JstT+
Mtw2XfRB7HyRrZkx8f2t+gDpaHQOHewYV2XlmdU/T18hxQOKW6ZGLE7KO9WZ/YuZ
29/JeU/xepgHVcgkUaN0uSHUh22D2kHdl12VE91sNY3JxHn5/zpirfBaFLzpPZr2
0dKiL1ileRq/wGhLwZBRPaCrK6WdHl8BOVCXyqu/RgXpEz6jrHcxesysZv7mL/Ed
eL69/haXAQOZKpvCajjxe/C2quztblPyxrK6x6o2KMllRGK9BBUsMjjdsYrte8v+
7EZggMRlzhk9ubXzNSGUIEg9kiJTongkfVwHQipV+UUnAuOII+L3AGJ3pDOD70Qr
WpGeQma1NCRbBVgn8dts5qYa/6z/6Nunxc2X67/AmxSgI0apL+aPYThkqE4sukdK
z/4atPnl5/zRgUH7soMHHHTHVpO3K5cnPWEOMBYqSs4EokJH1OsJH9MTHfFXuwFL
KAWgZzjGjrQ3HURlYCy9khJMIZtsKcou2f0msIVUDtyjPZ1Qbw0L4XyJHIY+J9tW
0PG6D8P1ceF3I70RKMFiRcG54doMJ9HxGTHod0CrJ6+I7rF8UFP9bVeXhTLJHuIZ
8rZL0DrKARrMctGCeI8gFfXA146WUcKrWzAzIgMcV5hcUwBktO9sryon+YlV92UL
3KnErsKvB70qpfkzw/oHRWjDQc/LfFfM+TtpWQqPXw+RiJu9WyBKe8guFXh2kcRE
MjafLD/a3CsjgGvaGbkwRCdAhdLwHGEqgaaNmWfwGJJsdYJkhPml6+dNy6KzGomi
IktugE/MQfbeItXARnVzmxfmntO/QngyHYQFsrmPlaiGLYWvN3dbM7AqctU1QL0P
8ZJh3YSDhRj4+PVNyEFtkeWLOtyorPJPaTIq7phbM9jkB/UlsrHYKyYnJn8Y8TFS
RHgs0ZlnZGdBLJD8dA9fd7k9LwoyLggJROxBTx12F85TqdwUqEHHsJZwrCcTKa+e
QDH70hhnMETflCaLqKjlGW12PR3STSIlPY3jpPPh5DXB/9NZZT1LUSNmYNKNsDbd
FjVF307iKzbnMJ9rlBBcoy/Zi9k+1diRRtd1RuDedTxNcQLjJMzieH3QoxCDxIHM
bE/+MhjXOYgH34BGyOi1Qgax6dOdPaLjWU1KRxatJUIUeJ8mQV2mey9f73yvOLPN
YfKcmidGl+Ez6SfGoGme37pLf/wLIWXyAdlBtrN4r9N/XWMeYzh6p8mEF4zlXFYV
oAqqy4jcHMrqlTrJ8ZzWpWkyC4FPnvAbxBVTJSJHdeGLimacNZhrXpH79jFMU3ZW
NTJiCoSkciBRe5A/Z38fZu+W/Zw9wcdhESJrl6F6gMb2B3qE3Q8HWlAUaM0uS9lG
u4bkTnBJy2qh/mw/jnwfzcoiAu7wfh2sbMEhnsxth18qn9vs9ZQDlmlI12L+KQhd
Iv2OuxCTW2I1wmnHlnJhcPzMUc54vJ6nvlUdWFgDFz4tL9VvUJUTdos4kcpX3h7w
DOiL2AkJ0gv2uD1bl/1tM5J/3YpUHHfq0ZhkKnwB5gpPKmdzLphRO4WhfjqrR2mD
/HyTsbdqQXVdFEcqpasE6I0Opo5BlNgTZA0wjY50Q5vfKY2lhfO6asK545ZgQTFv
rwCh+yfCEMW/hzoH273N8egYUH5nXzXo2eALJZttAgMuCXA4lshG3/xTKpPubxCE
EdiSSAh/x7z7KbzKHUZ7lcsgpSD/2fJ6bFshodRJTEewO/iLm8dYB13ZfXkzJSPN
kB+M/kI7qUQWpl64QtkKFSj1b/VE8ePrd7g8ph8W0AE9YUPc9nHVWCrE88MHsNDe
znxICaOzoZX4GqvFe9X0nNdHjisnbNdhFdSjG2C8st1nElGN80OnGTG+HcCC99Yy
KOajjCjNJzB/e6JLpTBPdMpo7waq1iclUCFE0XgjV+cRPFzNQ602acHHfwMlk+y9
K01LGkIp2J0S0oiqAL2qa+ZBQl+waDhoWSAdRP4noNLtqwuZzams50dl55+edqSr
QSng4Id2nJBeT6WMToWc/m3Z0mhlol+JE+5QE+c3K/M0rm8oN5qck6B+LkMU8cZa
DpNt7jPgiPe9tODipOWkiFLupOP5N4lKu+yBpyoMHbi4890Bo4F7ZwKpGwMU+jme
gpkKtnLe4U05VyAps+DhskHdqw6ojWbuBQ/FQNtbB+PC4YeRm864LXWB6+NHILua
5tBEFMPgBcubwAvSo7Q32cQiV2uHAEoiXd98GJpc0J/dD0nJg3tAn4Qdi5LqxznE
d/p9YMx8P1o6/SbG6S/rRUhbixwDV8y0eIrfft10pNNaG22KU2T6KuM4aM+U3RuS
g6egAaS9mWeqdmrewEYZo0vKZIrRg3qFy/QT1ZfuDY3x67h2OdrJAnz++to9mIhC
DeLkCCNrkIuU6mzCs5cNA7o8+KORjhxo+wm6agN7odMvG4M3yuxvzn5narU+T5Th
xRWo7KipOC4zDlBbAx3U954Zhi32yLpS8shOphuZdEz6FHoDyUVWFPsruJ5C2IG8
GtIwuiFxnBuesUmZmrbVDpti9RwtZWv9LdNsKJQBD+yYh42h9g1DcioIbWfzUOt0
RvHe4GaMfPDxe5HGWR2EaLpcYzhtKuRTnAIVatT7TLv3gyTMSGkKT9GJ7VU7+PD3
1gn1vfj3loAKhWTqsvjPuxCff9TNPRmEW+81qwyqGhDjsxbYDMFgimV366+V+Pve
IO5UzJVlbyy4U6P3FF1+Al2HiZpTfu/ktxqFV9pM3FeqniCws0134iRP4SGq4AWr
ek9lOxJIKdQX5l+dvI2j8qlOf+XxzZ6r1Zzt/aQMPShqwfhZRYocszKPhGvca649
amSregUG8fXIFKzQtTtafCqKIKGmvd7bfiubmmqXPe3PWG3IjdhcHsQm+wWTDPSR
ZCivxB6L0upLHnwXIMXr3DSSPCotDQcl3Eo/JLczPhgMzmPTDyZzQeOq9NpA8YvE
hrAfEJBJnD81hK99pVmXK5eSKs1z6uRwsqbAHagOHtqhsBp6iT09FrhhTgriZ8xR
TeS6CXdVIBpqwdOeKLU0nBqv3CeNbsVw8nJfe6PQ4s9Qo4XOID84FGh63DCsFIiX
frRujkF9oBy3jd/b9MJSBV0UGZWhpt5ppw9a+cuFWkU3n7CjSSaKPQ5x/17UY3Xo
v+xaCz1Gu/VdLvUO8RlWLvHj641Cv7iJPKkdbfVigyT1AjbNzRJXMehn2U/Rcf9n
i3kiwqDVq1YSgoYYwmsOtmsdPbhj6IIneffkAfoAiH62/3lPa/wu3whU3znFoVNU
+PIAPe9XvjlqLo9jF5KrORUrUE6TMsCpJuAR4/RLVrI2KOM7Ox7RYyaiCCOK5dRE
HIyR2EmxxcoOprNyqQR4FE06+3EA8lZP/16W1lBzxGtsC39c1NC4YztIJFz7w+pT
O50L07yQwWDms0HZ5QzFK3vljR4DXCnOHA3mnwdws0bnWNMkQ7jMo8XCRc5oeFYO
TxYwP5Ux5ZK+b3SqUGOhQIBcbROYsbr3e3/eh3t6qB5u0QOsz1yIAawj+he42dyi
OXLyMq2dRKVYp3jgQTHH8jwNzMtTCElaf9r1cOI91kw22RwX3/tzdVVVcvDk8sZ4
TrRVpsJBZkgOvzTiGHiKcs74HxBwdr4d+LaN/K1Pg9IjjF6v1fremeARopo4/5Ox
yuIInQWcYHNSoqIEhN85+jTist1sMs82gpp1P8TO4S6K1znANbzuQYAFEZsrBoEE
izDAGdUO36T3hieKnSa53E3+g5dpSDlbb9HVs7D10axAnxvivlm+Y4Yh9sN1pfGr
93NXupjbU8+QpGn2iTzWJB3mdA7gG5Sbwa9u+PE/1H37Zhl3RKQHs1/VI8KjBpIr
zTaIXnW6GyL95BrvUnW5zCKBnbgsMH8EIdf2Vf9YeFZPdaY5vuhuVO+/E2CNTU88
Ehf+YHk6iJUYDBkIEafJxjtYDqfIgdX22D8ADx2Bi7bAbZsib03mrlp1cULuvufi
m9Ep/pdbakQanH1IuH5ytEPO0ihMq7R5O6QglWVrgg2+bl7EcVCe/8p9ZnffpWUa
O98w6ax0knsj/sH569Gj/RfmyavGjocW/oJ7c5MKM58Yq8mtIcdJZqJIvwxKqyN+
KoTbw/iYcoPuvl0e6hz9IjEklHicu9niB976jxzzvH7PpWnYpSUzQx2S4+W0NPtJ
p1De7DuZJ6tUp72DWbfYRv11vyxr8ttfoWRggrJtxmDMR+Gwnf+3DGg7IgQubXsB
Woo+1BSCP3XLtkSi5jHutu96SeLoEw1h+lDzwxf/s/J5B8M6r6TmqR7RfyDpOTlJ
X9UEp3I9eLgZ0g94QLzYVseRn9jJ1jD5LbGKHxzLjy1lW1/K92kTT+E0d9hyYTk7
dpZULnNXNWcYgB9BGyeYrD6J9zOqLiV+WgN0/A14ApbvvvmaoHJCvq+uaoXhtfRH
6RZgyFW2ek+7rusVxFZXbOaMsFTNKXH6hX3b0XY4rK9RyX8uCovx6cFgwa9i0lm1
HBxnH0e6TK58QvODNqEavWUbat6G3wos6Qj/wWu8GWUvYMqukMR2RTk1YEgmyrba
BgJlpuF5T1ZNOb1DLce61gYDUERvgoWP0AlNvghlNkESvw5aNrezBdUNsCZWWpPb
SMoUANKdDhWWcXWWEWr1u2CGWBB9+OGtBykFMPIJqvJTKJPvdZxWD+pFp40x2CCc
I+3GbA0yPQODV+AYJdx4bcTESi9Z5kLeHaHNQOzIRFZrgsbca2BW0a8+CwQSAD6i
GR5Sk9aahcfFtYDfgjsHSJcK9tlnTXqEI5xuLqgtCgf2aRgfl4tcVX0LHYqpmdoa
G9DWdRZDTQHyuNTzKTz+rEbZ8sDMi0m2IpST86rVXhh3lc7tmfSpMBbq8+gSm/hw
bnjM2ZGqb8qZ7O7TygDryhf+ZMOk8DnEKNSnDQNTJMNy66huFrghJljnpqAIXmoF
S/842GPDAisA4HEMTi4MFmYt5I1/7B81AvBkfg/lpO4DpIa2oRVNtqy7AhOcSrfW
ZDLTELJ0FdJo0FqsrJWNBIqsjRh8sFg21H5SUFNPegUCumqEdGmkHe/GjRQe7GUd
ZlOtTmvQ7yaAlQYr186Q4vuRXdr7Ito6mH3As21RQD3VrZePQnjPxYpKXGcesfg0
y9lxU87RHvFNPiFT+wOjjlDe5omcTX8jSRA3UC34a6brKa4k/kx7R0LrFiq1HxTh
KvCsquXDvk/MTdCCavRkP5w4PlYoFTbM26Oz1Y8ZzysvZ+QixPcp0Dnjq9+N/3tf
dmpTybN8W8VJDKOuLePjLOaX+95mp6Nv4NsawYtLR8qVBTrIWHIzlmDbqipFxfmJ
nW8iySikRFUG90mFrEfm2odoZCfNRbJt9qFP5JxfstBqAKbKeUSmmCqqvpg225Qh
+ic/6CNyUY3jBSYGOOzq/w4fVCWsLORS2wC+Qpt+RwdYoblbtEtbL/FWvAl87fmx
nguhxcLndREq5eeaVhwCLV0SUZc2LUi/Mtc7lbmlC+0bDpNkatMpzHIbMHUyktY+
5BYrxIeP9B0CMJF1moqUZ8ulV6RCMaLJZKbyYtIMNTjqpy3vzQd/M63Ezz5qOdjH
0/gsEp9rtheVFBHiZ0G0FLaKL38lLfVL46Z6YoEfA7FYqL5ckvvpV4TVO2iSLIU2
dSzxU3jhUY64JhIWCDXNKEL0CCsUeBdcnAeybnas+9uEoRQQ+48ahop2dVpxfp33
fdfQ9T8QTdZvrUt3la0GMgWt3P1fWu6pHXAtt66KIoBNHuCPz1dgVOEpdiLha3Bl
FCwv0n/GAAgykP9urQvBhC68WAYIEK5wOHk2kSsMwADuVhh4O6E+sJpiyV8w1YIu
eGlMt494Zz6q6fy811iOhCXNU2c++JAYn5mAuRIr9i8Fx0Zgokzr9qyQmaT3Prpn
nmUAxq4qKkAu4atmXr/zRhfVdpwmWlRgGc0jPDO1PGuRCtxYdmsvch0xEqtBCEmc
YW48d+HgnF8ESecUZWIUyLvrOBLMRYxBdn0ANdgzry35T3YrmMCfhybRxgXGndtz
5h9iOoxQEe9u9bTq/jyoY+/mPbyt81m3qcqvCcS9rVGMi/68auxApA6Vvcxk8q4f
mElXox+cpMKGgSdsUCwDaqJJPMv41QTzlNgSKWAxZUiwe3+dtkbuAV/X6ij0vwy4
mUvQrqSic2OMu+KnLGIR6djnnqW/aVE/dSJdmu6XDziGwBbvFjrDFwzwYliN4fgU
RiyI93QGyZEa2fCBMM13L0JD3+VQjgQ78z6nu1JN6ZVc041kRFz8zFFCUcf60sfi
TB8G9fFLbsQjqzk6Hy4+Ugb06hGoI3I4fZ3usLWuPtrSaY0bGxy645JmJzUyAgpL
+Qvs6XOP4tJtUCv0YbLB2viw3Xlig2RiUwBjB5VlxcjMx3o925qgI+1anNgaLMDV
VGZgJvPa0S2gK9cYwTL5XMAxWObFD6hs/yChPaCu2o2zHq8xIuk0AVMaWKtinKnS
9Wkg7GGacKgnU+p0RJFCt41gb4y/r1zuW3Ppkgr/Syo1sJEhHQDylx4Gt0I0ZsCG
Wt2rLNWWbbGVsyheNWNLrizL1D9o4QxHpp0FKGEVx629wkp7RaOBUBdDIWtt32R5
Tnmxi9QWHEaB/Z9YmRNz0YML83wWgz6+nlczfRal83I/WSFoi3WDT5D59ZEKPfBT
3p7WKXThHmPFvnKedx7RoMwWgGTBx7wEkCbZiwvb7kf6xvORqk1Ral0sgCVCQw3p
KwXVJXBzrB1wIxHeBfJfTx6iVL7fH3fTdZRwWe4IXRVP0t7x/9w3CQTI0hSywYC9
INz/IVG86ch/zWa2j4PbQj+1JBVz5t44sEQ9YvkrWM0c5KUmECLkwun+Y2M6z6Ec
bdI8DSKxh/UhBVo9gHKWLBcdI8OqSMmhKGIqE8UyonzdnGFsm4yG2FdLT7bnIEmO
iuJNOZNnOmXpENsdegN5P5QgQbp17jXe3g4NfM9xhH7M6beX900eSNFuAH4DF2qM
4EDqRB3M7iDMS7J7VcrkMOzT2r3Vazehc/9e8b+bJzjrJyqO8+LYCPWVGiFIlEaq
PPNzVmud1afgvsJwh/t4VPOVaDCLs3PSE4chj8NDBnoEHgEX6DZNxbaj8DOBQ4PX
HJABjaKrKlnBZN9xAV1UmhCHAqjxEJu758X/Upj+czA3TXkmc0mBewXng0t9V+NM
GMQEEgGbRZoL9JNdAwi1O+1u0y+PKzdbHrc4jRWrTqu7vCkZ4V+aOZlFdCBN4i7P
JuZe2GhLgC0385xo53r2TsTSS8uJgT048sYMXxkpRyYnRADL0Iqdwb8fNw7PfBTm
HMLKgtvzCesHCA7fHvIoRNctK8rOFFBarKHdp90XIl+LDfrMvdLRYFp4s5D6Tecf
3fDQkAy/yXMKaMD7Bakjst69zAV4DPWGS1qkxfiqAsBb+hv0zeLTPKNtqqQzLPyH
JRfFpGvlcudJnKKKA5vthPtoinc3VbOzCWWxlFSe6xeDD5Yv+NDVJv3Hizg3kAVH
Zt3SuSgbeqhDlX6a26GEWTbF8M33HQNy4cG+/VLzESZWFS7MFNjIQrdFHKXIzNp0
funQ3n8owHAlGX8PHv4tUY/4JBAdn60aK123oZMitMq/rAtLUgTqjXBDrjy8yPcZ
7tMX1HAfKZt5uYdUmzhth44f1oO/ef0G0/BLyX163rCpsoAMX4H4sw1oo1oBO1+S
RDFzBV7DV8FG/oZZbYuUFr3jrAmTS4vQmDEGiSqxv3SNJ6+wy4uYjP81PLdA0Zq5
z+Bv+bczOQkCEK8wWdulC0ApF11h0u/3QzYnETN1c9hDa4kiVL6MEzl0WkeN3hrs
bE5+OfU8xB1Qj8zpWvAsf/gAkAQTKoO75Iyd++gWYoPL8JNv4uWCjSALT1oYcuK8
zcYd2FF0OjIKUpHqch4yh3DxidbW430m5SEACADfk6WBslLnMb8c5M8j5eIV8xB/
FAHhan701eBoTQ42OXPYLK5kec40Fq02SXrCfkwG4qmnmp7H1F2hMaCMDRBlWfL4
7gKoNeA9SLZzTS9delN+jWKusKClwtHZnrvRbc0bC19W7GolvcYMLkqNPe14upJb
86Gn/bRThkI24V/RFlBed200I/eCWgQUnO8rl62QZNj4cQ376OanKKCu6BFQYDmf
fcI3XVPzkDRM75uB6t3RGgSY8NogWH9wdHs8qYOim7zxff/rdyu9rTe8zivTD9RH
iBsfWrjSRmapsXMG8VTI4lJLmcmu1XCT4btEhk+TGXPM5y6YnOSU5T6OtgKV3qLD
MmKgG6AjShaUSEa6u/4wUC49xmIAd4E/wGp8wfP3D3R8gstAWVjXaiuXM2vqbwVT
Br8WerLNWqZw96TNur/p6Ks8Qw/ttVzecdmgv/qjSb7mRad84ueMzYqkMd38TNwa
lMSmQcIcn122KpJWfvLMJxuiNMFFhlQhkUNriBYmzqBA4/oUsC2zF5o7iijTvmeY
+BMYm47mfJhhJc0PFL1yfLuNHYRaa7u4Nsa/66uiWwkmyKQHe4IssICsLxCYB01I
AoVSp91XYnWfnidrwS2ZeP5kEYfAZH3Hu5M9TmHIm5GWjPwmgtWU4RZkfKwlGhAn
zLbP0oAXvEnzqD+Gg3L/uxM5wpbrwEJQbQ7aBn6cSh29yjKlxsLkH8l8Z/njcQIv
Ga7ygsnksJlI26tKb9sFrB1t5LZX+CZcwnRaZTunP8FuUD8Wbd3I7Lzf01cOH+Kv
LWkKh+jn/fSFoJyhaiE9qJHiGG+NkpxZzIt1M5Z6dqYwtYOh+biqQp8GGvnm25GD
AS8YWX/FrqzSv4iIRcHju5SwZOT7PaSq3jUkHUz2njgBpymJVVybZoTtKEPF0etx
gB/86uK/METTlP8pJxk2F7/AfKlfE7fIX3QK3FUBhr3m6tkn50T/2CfDSCxBQ6PR
Da4t09i/ORs/jz3qxkuPcK1mzeynIRH9mzvDGhIntMd3LEXmpeIEerBm4gdD/N2z
CDUn6YgY95z4YlLTPuuwGNA6P9Dt2bCamM7ACDE6S0T9IEe0Fcsf6TsyOaP0nXg7
zuuPZ/tJbCawvM/32jFlgBu30bPVvggV8Pyniy+2656yWs9AQ4jl+IOi2MyTEn1z
J8E1R+qomxJ2jWW5nE17Uh4cO3ThyZmYKSQ0f1wLP4s4fy8pRw79agdHL15GnfEm
bdalt3jZ/giZt5rDOWpf/RDHABanlZvVtoL4PFMBTUpouetrW0i3T3mvF4PS962a
1CV6T0Xoh9fnk7TIEKs6gVT2W+5iXETdo84Af9UoncVuf7k8x5xcc4uqET0D3Ej7
gHSdk14vnCIBlc0dd3Y6vJHSTnGyny6It6ROBdw/Itl7F4UnhbpYYrwKSbDlEtOD
UBailH21D8rI+666dwQQQCFc4J+DyMz8vX7zdoMwBNYktZ7LjLcrOecDZqZwnMhe
n2Cd489qLE/bqvWYB7uQhnRDFRYnl2ui40MCX4bS2hNQGr1fQ3h2/kNK5T+2epKg
wzvXdgeDrM01PbgbLsssCMcU4e0P9QEWxFRj1jy7KVnqyXqJ45l2dwzUwOO3mSSd
WNVT5ZXotYs4N4l6ahYg8lfUMYRbq35H+0gGIfrZ377qYUN9gcLtuXhAF/nC05Nu
itl9a+0aamSX7QBZcySCpivU9nm9SEeKlNgkh4/MLVhSvYOLXHpfOBibHRHhFzfO
bPksboO9q96a0AHm4WIiltaPGD1598im6KdtfoZmV7JtcTV6D493WtCEpuAM0vzN
anxHuqQ3OiD5GHdr62lIpz97jOi19Cbkn4O2eIbG/8pTJ2cm78cFotXS0pnA+ioe
0XWxUZgj7+ASon8ydk9WmpT6ayaHsEDoEGl27vS4qaampHVZUAJHb2Zpr4cIGLvo
ZCT4fQWpEmYCn1d5FvEx0wJJyYrNUxho5GowJLZt1P/NOe3AURQcOwyvn/l+WuuU
wVFHimpAuQFlmggEnGuKi+obrdbwTSmPUNuFkVhkLMoF0Zv0Zov5fanuJuxM3i9C
nM8gjg0TDu8SA562aaYnoJ8cEej4WtJyLtSKNl44u8ipApgXa4odGpfXNKaAbwVK
GM202uJa7EwY+Dd8xG8G3LYRTV/knHH35pJF8fr2UQaIIXCMZOXI0seFsfO4UdUt
YugdB3aOa+Zh4qozMgWsjV+oguzAQhErlX7qPjB35T4esqGwJlPX1iU+vhTmABWW
S7FWUfdihMuAGns0K+yIO2dMpRn8t674PbeLt3hm+lSAeJGKT5GkGgBN7cGo7KMT
6UY59qHk5cDuY4kDRCBl9gcfAOfoiZswR0PRM5xIJcTlxM19guIub8Swr+G77OVk
QD9qY9u04o86BssST5X9zvll0QEJYOa0lcwPmcj0rMTubownEWKpgWJ2YHLDEGAj
E9i1noochgQysPjbau95GaGqIjNeqddn6qcQUZamjJ1xF85GI0onHTGD8Ew1fESC
vme2FEnmh284BQe4of/mVLVU4/e17pZdqzloBwTHMaLNS+xeXohfjewAL/Fb0CSe
oXSjDTozdBksPRYxadrgwewwGydtw+JOt/1jZ+bPGH0+VInZIeNIWJ99/DMTsT8C
AssctZjGUD2AVRPZ3y+2jyWtUBZD33dZjPimBrep7CsGmF7iD/FsyZyUz583/bvK
FLKSkv5rnAmNu+M9z9X4zWDfWzOFeLCALac24gnA2kUxj4UOCSuAi4e62XuwQLqi
IWuoe/V9SDBdP74a7vkXNwQvZ0wUEMWUybqc7O1qQLXcb2s6ZpWZ35/f/zTejBMg
VzvwbBRGc+3izNvLixnZBAtFcZ5En/UyNYMynCoI48TSTLMgJRdKMdbSTQZEnmnY
BBrV/HUjdLlRTMflFK+PIZ4p6fKkpDEYo9trlJT2Ce5zLVvdj1shvC4Itcn9rpOm
b8SO8BW0iPqyfZ6WWLgKMiedM8MygHoZARuo7/+AInvOYz8xrXR7bXAXE+ppxKHD
krXO3JLqDpstID73Ge7sjwFKjKbR7tlML+RaL762GMY9ExwU81HYr27G+WK1OILq
M38pihVHP5WN5ALdGPEoTEGp2dU7BWp/eukoBWmtnJOhRKhoiRHjJDdkIl8sExE5
7UK3/tWdi3c2D82KP7+2K44WyQGMBaj6y8wH/ZdbxUQgWqwJW/Za8DTmFaLCd/Tb
VhDYIjIhOi5mjN0htacDEJkxjRNcSOrQpJq7C1MMGNmJzgjurJDblY2ksySEcH/G
Psal0DyG+JPvETnyhuN6wmk5NF9ONcZzCPhPCKUfa+De28iZzNdYMKi1NADeXIJg
oC9VLxSrKEPE74HHIrmIMtvhlBmVFCq/pmPq9Lhpij1++VZWZoAJXgO78vpZcBWx
dh6vjRFEg+Sg6KjBTqXQkfo5fHFeW/n9Lb/4Cfdk2ukdeek+9lNhB7uzMgHxrAtY
Y1Uap706sWPfb7222kLcEa3ZELvbEm6tzKm9O5fGHIzLYUA6Z1C8FKdQYMtlR3SS
Ej6SMTl9YrFdaRDvqI8v3EGCu5R2PYg/xQMI386Ndju1gUvWvQW7W0xDyONFV3eo
vEoRxdq2BI4pH/hadLuFea+uOiPv1qP4MR9TeLUtSCbBPYGdHYpz8KUstWajqSlO
Kkb2d92Jrqa10+XG+Tc9zLGA5TEV19Z7H0g4gnP2xBOZgDdiXqEHfavuAtrTn8JD
BnK3w2cAqsbK9+O020vKuPGh4YzwNHwY5EAxnnuz2jDHT1bQs8Mk+885AXHnJJNr
ab8Iz088QVoRVuMbYA0r27UQXob/lX+Ah8f5kxPNjW5W+2FRM/U6B9T3slbn6gdQ
rQ/c4oyDTfylNZ8KjWJhNP5gOEMW9vvzq9sOOJfnGtOWX8BqmTDZXqjM/hxOoqz6
HBNCm+yyYLFlUiptO1JSGi9bS90TlcMmkp+TaDZOtda2dgjJwjJMHvRjeswMk5aL
0CxRj/Gevm9EK4QfXbokga6ZkBySj1pf71kU8VDS/GbzcnBRUQMJ0NzhQhK6zTfd
0ewOpXsIhmQ1b6k7JsRh0N2wySGY8HaYiqBKVDg0+/dzAYgRyeE1rjz9KvR5SN4o
i7IEg6pRzHosb2hs0Kr9EQkW1Czo6kb8hWtfgcDdvyROP1P+6zNJCUrlmWh0gCcu
OgN/sM9PJaWX6zmHe8iwjShyoPS9omyrVqSsGEjSAJqWxz3pi6RToeok8CWX0zRA
Ck/SQUqcCoXCFos8t+qwKQ==
`protect end_protected