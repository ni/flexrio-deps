`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 55056 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
hRRAlfE1xLfeNfywbrz10MNI53HD2kbyzTp8JdAFOC7FCdNDGaMvbFM2gHQv3hkP
1x3wJcYukr7SlTatsV9T+nnH3r0FrcEMZqp4KEA4DXgADC4HUyZtS7roaTeqPP47
j9Dp7TT0ozHb2ExCc10JttwV660UeKg/6waJnwfdXKJrsmbkuLAgBMCnnVrGgAZA
r1CSZN6+GDk3QO8Nbtw1ETahzlFAI75P9xuW324g6U436PC2oNGOotwwe80pLzLc
QQNS9uIbf0NLxXQe+9YzqXn4HrUYE8q0L/+I7WZ1IyyI8xKfco4MYikNK6DjHeNV
CnNmtkF+P8errC4aHJ+lhA8hf8yySw+ALsVbFDvcyM0hedYXPAPInpO23MAuNk43
ToHpjv/UHSVfJwvyC4mzwB718jrtaBVEihQa+BcqpdopswzvdRhMNlBD9E0ovZPx
IYsdFW6jYvE4IXiD6/Aw5nF+/8LeVjQkl4VMPZCmTQ4HpEPAhTjXFlAaW6hj+L40
bHUjBRet1xUfbsfTULQ5O2cewH1z0WJ17TIT1WZ5HAevpmUwKTlwdkcMTHi+bvW4
7LMQtgDu++oEfxYqzL3dJGzPA1Cua4zFsUvomKVoJF1qLC59vn234PM7d5co55V0
0h0pblmi1PDNhVGpniND+LzWUrWMR4CUmUhQVxajze0Dx7ykywGGTj/h4QA3G/+C
kegZmG3xv4qUVh75XXuWf6oQH6nZnNWzEEmUUuazwHdszceYQPhpM9uPXV8tsGIo
BXb6N2gVjq03duH3NXRWK7AvroU7ER2u6qz3CVX/7+0bQi873B+P9BF2PD6UvV7I
5nZ62DrEy/oI8oaB0nC4GMl4lswA5qY+asuT80OvCh2lXvL4ZvkJAHpavlIwzdQ1
I1GWK2g24lE2Rkd1kgkn2lXPEGbibP3Gk3A5+EsjRA8e/IZPHZaOA9rMtVAMf9Ez
HqSNSC8IS1klRJs5Y9lG8jBrxATPfi4/KE+MSgcnvNgRqx5fHjDajYDupqcxpaW6
0mpD1d++Mt+2AsyU/BHC5v6Zy6wEeSC+lM+ryYckcp1752F7RIx8wLhioQgDSscF
oNTsyZ/Kxtps/TVUZGtZAvhe+CJpmunwWvUp39IcrEDqD+aMrAt9LQ5V9ICgnWAK
6UeMUrs53eKpwrRY4ZMwGlKFn+oQ37VoB3nJiRWrmIIUWclLrSU47PvepO+vazwn
kY7YSrDjbnY0OxgOrAMbBSd+paYzkXaOP8O0glCU8ycyio2BOduLDwkpVEqXITLs
PbuN081bWfRlYsUFBuOlIOezMoeDalp9JFi7oTuDBV4lqd6ofxsA9Dtm1oV6aeC8
hPHkdzBSWe2PnfNxhi7SXiI/Z7j6bAhp7k/aaLOvY0yB0dYqkYK3LgMjAX5x+Etq
15cUCO+oSXNt18LawhfHueV5e1fwArFmal00byIx7VtCMbg7B1P4CiYIqj95iOZJ
/huXZb0P3Ii0S7EKSOoQ5WrrJoPjqWZcIXT1bo6D5d19iYS6mgfcD/0OUO8izpAk
iivW5SnmI5Za4aOUaVVOdkgyrJjTg59O/4iaWRhdYpKj7h+MeN8WNIN5TTgT9v3x
EOw+Ig1kjObzUfF6HLV2JhsvNvkjJZu+hOY/VZoXb5sgtSWSzhfJieNu2I+wuNwN
M71KO9Yo8zy50ivp2JqLUrNphrKXAWNyEmbsRdcEYgCUDxwVOy51yRPMEdQ+CcAa
Qkxi+CzhQ5LmSr/KjbJt351mvTmphffO2Do6fAez7ogq2xkPRWbXa/HLrvPhWhrS
FuR4XB+433ytBPzh0WjtBBMmdbE4LMAlQUg4Y29pUEfxnTG2Q244ro1ym0Uxj0Vu
H5Ll2DPPM7ET0Edh58qcqUTDhKFoYYAH2CfLwlHhtbONr1SsCyzXwzDfYp5BBSEu
AJECFoOSvAWLZOS3hSWlnMNvN0LbAo6b/99AyeHRaJ1ISicq8p45SkS9eRDNZea0
xPAnPeMrrUPUAO7BmJF46LvLs3QOgdYIH1dxxijVox262csQzy/ap23I1yEvmgC+
HyfyG+FsjK6L37tjGRAkIQKm3/s/9VFrebSVPYcV6Kf/gH9GlWcj4cQt7HmtoE71
60o6VjsOFoaXI3d+gwW/WBGIQ1dnafbLb/rMM4XB2vqLxuerYBGOUtrE6Obni6Mb
L/oOMwX4DP24aYgCgXSJR8Xks3I/k4BzbbN+cTqMG8auTqNR9yFAMGGbYG9MciJU
l/uNsyAJzfsPyFZcgqc29rmA06UK+Rxji2KfYhzlQY4YinT+/J9cRdevVxD+m0uX
KbGrIAlaFMtpcv2cBzk7na1RqE1PjGjeE19vC7jMoXHgSbVoFkCTrqvTy0KYgzD6
nVMgscLKrbLpMm7PNl8PFoTAdqsDgATO0EerAIoUd7ibgoPHN6o0iLowkrOL6jbu
M4mQprEYyyMnwamMs8cQD39RDfYCZ4TF7edWaoieHRTH7HHmrlzsgoBfn25okr8x
m/ZFFafDG19n+VFwWCQRytqsGuRRxo2gkdjqf2LX6e7xDN5yeoD1GXKwHr8CAI+S
vKm6VDobAf5xgJZKxqxz9qRgWr1b9yeru8fnYrR2FdZuy4nE1jWMadF0JB4oSMuN
LzY97aPPK68OWezqEKcd9Ejjmq5iQvvhE2yzF9I9+8iHCmPx8wSe+zVYoRn4B+wI
Zlh5DFaVrrk0D05iqaFOdB12Ry+K2jyrWjbWoWo6EOfhTIEAQyGIAmfb90VBGSti
QngcUmQnpsIwp5pvEuheAZrSU4dT3w7JuHzdLu+icADGqoiEob2JQwoaz27Mk77r
Z0ei95qeRkRQ9S15xpSv8csYZ3DcXgaEPIlbFFDZ5QyoErBLJA7bYAb0mOHXI54n
aXxd9jjQfMN18yvfiFycAvRrDiJOO3b/bGA+RSQlyisCO95iyX1KwnAkVLuXYN2j
52brpSefC/xm/PCBgrKKcxm/oUVhOqnKSXHy6Bqy/hHsib50XF8Q0b3XmeXZepQM
j/e/b2PfLiOkM1dWdp3HwJVo5YBedKt04SCF2lLo2hSh31ZIZw22SyBj7lfzMfer
05DuGwdjZCCfgRQaWgz/dJFqKsq1+kBQp/ZAfNJWjPaGgnpbW0VsxZOZRLmGG9NS
JaqZ4YYCdQnOOZHrmrpU2FhK85yUgM3h+Zi2hNcQmFaa54+83sTKHKFc7/UwwAUW
wfbvAi/au8XdZ2BM6g2hiL6psPCFJDRb7QeKqnGD9xWgEHOveB7IcixBX046PR51
Mwp2O1XALdnuLVM/TJg8WKbMpl7UN55hGbjZm5dE5Jc3Y57IuT2Vfn8aPIYHvMbg
+ZDtg0H4ggmWUzghydl9R9z6YMJbKHnEJPQFIOg9zXPL8vaKNDS91oDC67TN0jCz
O1tqU9aNSk3YMpo4p5eN68Yd/KAiD/6+v10LVsK8j0zP41FYBPQCXlsmk4oeqhsw
4wtAZhmcJ0wctUxe3n0ZFMuIJtHngWeoHrBhYwNBYJlYtExRQqkjPicSmpk/L5WB
KEqj3/jDeRUW/WUj33TiwO+vVFEcsOcNbSJmAbLEaLgFyCwbZfDZHecizQ1AVeGG
77Ox7TPdcrhBIzJlZyBAnauxCXXolsAsHlWqi+8bA/PFcKi9vQWSoKoDWWIjhiIM
rJUgINljkTI3OvNqE+vUTy1JANOs5+0iA28kwE4GBXaq0iGPBqFIKvfIkq4V9iu2
GknFJ1xIQYVXtUaC02nBPlEvOABJMauc9UuVX7Ng0Qaw8IVoxewq9YfAWXoya0kH
jr1y4tGXAxBtEm8kzXepQKp/HiiIUrlGugO60yy9AIcJziLJrJgq9rqDIM6gC4OJ
8Yvfb9ZFaeekQVamYjF3iO3PHNBMkJOTUt0jJNEoP27wGWLLx0kQ7TcXK+9+6ixw
7PZwVbeKUlPn72iUHsvvVIkUKvlWL/KZreQAtcqxVTWvvUbyUkhR11ChfaIZuJbK
5Fa6SvZhnOaK+xl73jovMqIXXs3ak7MvxEQl/EAEsxeCB1IY6TFSVtU1aAELRjO2
853uukriPby4hVUur+5oWgMzybx8zLraeQA5F6Q+K1fRpIX56jq11bx/6NnHxNK5
5R3JLVDy6nIoze11D6nb91xzQO+GvhLB1+fkTZogoQsnmuL9aKyi9JYJGlEzIjXc
yuxPzRrpSMM+q8V5QT5RbhVGZjNA6VuuWbw+EUvkndqqlSXPvbzbV1+NtpbO17gb
oRQxRzNKsU7Yc6MogCTFfKIddWvaZfHFX8alnhcqAHZJWPl6p2Q7jqSGzRxwlCHH
G8HGPnqpxkpiUwgTyxDZNgHu5g1s6X7IJDkcOGnUWDwnCz5qSFdqFbb6S6t0v4UZ
KV6OaoHUYeHNmkdQH/t4K5oGEQtdvykxpWUu5WZ3gEY03F3Ta6NVlohtTlMZ7wao
PLp2UMAGlMzYoIlOApltfuRueSlwxJjN2UrrQuvMIvu7O6WVzn9NRZFey8/MSW2q
d3Bn4vWq5YxyRIYRCacavNd2jnAcGnFCGYtnMxmugYtGA7fGb8dypPXw50kyh4tx
zYCFX2Q3TuKmk6n2lHXLy9a8UfzEYXnRKlt0Wr/vOaRFHd7HZQ1u2j3g/DFMfnsD
Y4+fgG/q+36O3tugJgVKGwLB034GLfg/+RpRoA+MQ9lAF+4+wqtTQUNkouiht77t
r9KqxmVFCd53NFPz7w7QVn6TjShqyNYT0c6uGWrFwUGl9rKQfRFBgenr1wVUH6K8
IU//LdinN5wXvvxUbUkfTXLFxBe4iG2AUcRJl6ZVJrFZolyofpyf0uSLHFImE6D6
Q/z8QYFMfZuum73/y814doCTYYAKZqDSyaSKdDApQ5DaUhHXCKDwt9LtN7o7BH7K
+1A8hg7LlCP+UOn9eEBFJATyrHjE6G1K1quKTgb5j6sPpApdza1ozczI1F04I9Ce
VuGCJzm6SNF/p5OLCQbt7y+ZHAD/waVXebWEN0DcUrgUqnT6IzI451mOpt2jgtbj
Gc2NFbZMzOtDOKw8vRXncwMyRbMy1KSAA0RA2QqCgxMnWsPtWrOKq2X5lCvLq9TM
g4KPod+QHJz7EdqPcGwee/hb3lpI01CNHdI1w1Eo59wxHYVLRUWxhloFDh8NIKW1
wcxcQTcY4bjI20FJ+z7yjPIl1N00MWmSTtRDtjbLOQOan57UlQBJeCMAYhG27k/M
WaDbFNCHrWA/bv4w9VMn0Y7y9S0H70fVspNI2VtAJfIHJxwuAfVDUM4j3emKpQXP
PrOIU0wlg8VcmMTsrIy3DXAiUzmdSNFuwob2wBldd2dDgZLukLUDLaGkMPOPHasZ
jw1/YM5uZxF1bl1Alb5xzOJ0LGW0eZwxTfEwVKw5nfHtaKbcoHLdQXael5cqfQs0
xLkDTq9jaYv56GETOabl2KlmIZBhv9GvSrElMr+6kOBPGDsWws7yDbfQ04oPmeNK
f4nnbNc/YBkiNJEbrJ0rtVyvy524FET4+yaDvB3WY/pQ3PYbU5FrqcbOEtVN44rA
5b3cHhz7ygJBZ4D70cNpWimtCGAXMsJgDf8buGEOlBWtoeqN7JXU7XFZQQEA4wBW
szcO4kp1Lk2NubbQfmmfkRlzTHhm42Do/tHUk4OyFCkqppiAbAD338Js0C7s50eC
ZxZRITbU4liwKrQ+t3ar3FARLFdHeWpHrN+6GcmeB/zft6bNWFghLr9G2ecjnDXP
3eKbSuBfj3h4r7xOc8tsn5zcbvwM5rdEqtV+/vpw3bWCeUFp3UXQSfTH8+Sb5dNs
txDQCOM3HZfo/TyuLlu2lRIx/rCwBfBvKFyEvhg4RmbEQY3o8NEXSaYzarGKnN2T
at6OLxJxds/fQq4HuQnnt7Jh8mP8e/tkjL6aeDpaPxNIVw8ZSqhY1kDk7UBPtnPE
NG7ZF8wOsUOYHBubrCyKZ9CrxFTw+5uZq6jCZ6clhkKh950+44kPZ0KDOebRP7DU
hvqPOLCXpGt2Ksd3xW2wyGrKQefusKt6xsaODkdFNzJVhgincTyTRjJ+M7X2pTK8
VP0xTGEJ6Yl/7VFwf6IhB37PRULhQKb8/bG9WyqEkuFxWHIbvzNymWICif3/oXak
pXzkP2h7TUZ24YB13IHo9h5XDWmPUmMGkznr+iND2jiT8AHQ0OohNWtBRHfd5S1u
qkBwYm1pgcpLtMitgjpnSkMa+S9HbkB5tyl/biaCMqgMk6XvlLpe+Kzq+c407uDw
P1AgeerpweC8IvwT3XvPGDTCAtQFFpRW0w+LnysPcmjZKcXqKTFjvxqEkkXudNAF
6r3QwJclfjFfT5d57HE1pDXh19Or0dBRQKcG9OykMyUsUIedf4OzwXmO99brGwpY
vvQJ0TrDQ5AMH+TNBbhhcWWNwvcD0ncLrgHAyxdas5SsicdFuqWvQAL/WpVAQDMC
5jgCSFf620KJ8chZj8VkdjmAswUiTZsvfmn3U3VbO+Bqb3OlXl3brUqPMTe/Fx1T
XfNTAPiOJdvAw/mWPKhBYkwdz+mmC7gKjCteU2RHrjLBn+UDKX9Jr83Pa3Zanhbe
abeOzva9Nt9zdvR5Gqk7nfPUz/ZA8mHb+RbtZ+KSnf7Ov4qMlkytOqG+MbhuGjFy
MTLMg9VQ+wfO4bH/FDa6U7uS7WrHD3TGh3rx7yXYrozpY/KI1ruaMcNig3RhNuR0
Li9YhmytFzfw+L+EupudN8SJHJEf+O/h9z7IOy47Md/qMYDIFJ+A5KcuRB0Opd+L
h7Wu2KFjSZzqkPcSLOCd4QQE6iKw51JVMepZc66+DBKvBue+zTEOgetHc2VzvzV+
EjKQStzMwi1nW8oDah/M9viNGGf8cEZbBa7cZDxdX6wkBrQ0qVy+tuOYiX84Q7rG
yES8I8N2MkAGwjUJQwvFDK5YL0fKAweW+oVqGBZX5GdVVMyHJHrvFZX0ljqYu/25
ShKCaz0zLm0OuLwL+MHYIvIZ12vm3oRKwdPETNJDNHkKtRYfxQaMkzNrm8BYtJyo
Ar/l5GGLlbQx13rc7LvhEzz8NayvcBTz0lwL1tSSGd1XFh8ZocMAEv14gh8v1Ds1
xsLhFRg/lPwojaTswvJyz49G4kelFa7NzhZN07P9SiGVdwhGuSWYEFByu3DlumuK
4Mru/OoRNJqJ22qu2WGdsOEAkmKxq0w1HFpMjeVTKTDrHehkuNtoq6aQXf91sYfl
l/AugWE+eVd6P4vw9BtGA7RF2RulAS4wx1hQEegRocFoOZIHYKckIqVr2RZTVRGr
mNPoQLG4zYxz2yqr+hc+feot/GBEXKRCLr0Pu9zp9lto7c5sMrHYzN24XCLsYJp4
a6CMjZPoVp4EgrmZ1TsWtuZzkurEeE6LmGmw5LgZhlEoQoBW1CBYx9c9oIV8KGuG
PiYMAvXxynKlVCu2ka21cXoUCkhF++oz3JrPJ/4KdJkvsGlV7+Y/IbDc0SQkqH1a
q65yOW1rAs7hqyrNdCnpbucYW/kl/125nAAbM8zJ7J7D8kDGqj62QclrzbH6D3WD
zLa+6gcEo99fwq9PVxZo4NM8TJ4WMe5pI4G5YbwmCvoIvisAtH/h8+xAvF9FPvM6
66VznEl61E2XkHxg8qfxBIuWpoacJ0dr8809KhEghBOxPO6o1nwGrm1tuSFIjAlg
XnMAIJYo7vyJgd/lOP2cXe2buqolNQ/Gbyz9xkS/vnf3cIglSw61422768oLeD7G
LTOwt61tBg72fDskDoX/e3kTzvGmSrV8pgi4CRLH7sJvYFb/0TUnlXZk/01nHMW5
FlhVeRzDCv1VC5LRx1yaOoOy2UwTEnTl1lZzQMER7dAg8Nf0LxGfzfA0VRsWmwoj
G1uaQ+c4y3ykSe5sN23xAkCFeWK3S7Qew/rcP7BQFIGgDkOjfEH8J0LqTWihKkDZ
Ed0oyfuNVS8HsYmc/mmEcV2CeP43G4dfokl4gdkvZ70KAjesCzIgcrU+OszwFnvV
ddrmUBwNDmMNhyJ7tz+Gof5sxZoY3zlnv40w0zrxlbwmS/DqyC4EfSJw+Ct0gTIw
4toYWQ1HpB7vaaRLSZWoDeL4rWkG+xQVfdxkDuKpcQ9nI2FvGRqJ15He2mFPcjPP
vmiLTjJKVOrgaPaUbvYWSNMzfrQeuujeNTCN7ZNFAPkRpqOwKKCuphgy16VN5XgA
ZgJ4CP5cA5Vvhx8yZxHIJRdOFkar3olLCPndyF+iVjoOuedeQB0cVJY3G4gTZJP9
l7WvSswp8QxT6624H7M5jiFdlLYmX6cG75rgL3EEQRXn8qaS12nUybkMdwq0APSW
qyr7RvvQz8tVcOdVI+najP1ya9Vg9dyxSAs3JyeZrNc7jn2ABRBKQMzMns2nNF82
6y5YDF9zS1dVExdQHNe9Yfy++vsjcABkbsdggEJ6tyut25q5QDMOxfedM7FD2W78
lZRWiIRzZo0A4oBZWzNYiQKiDkBOtZ5x5vOujLYsOCC8DCX4IZA9gWpULEDVckqe
795chaQVcbAEhQq5gY+ims3oJIGReoy745sdTRh8dZcTUCj0z+LxTQ0FaSdZT1lE
FhHWk2lAR61bPzBkTqWDgvmn6wLbOoCvSSuVVCuXHI4IEN+KLJrZYfErCH3iUyCC
VOrOz+th53CaW2CmROPtzWruODKitj1ichOsiTmfWLDJmYfgbgbqBcHRuOQGtSyj
XjiCugUICPIdS5I2n98obXDkvAI9vjzw0lxUBo/cAmNu+tbvPDMrID/qNTMSBTwp
ofgYsiON1/HX6vd1fcbhpp4ipmdpLPupwrcBtG5TB/faGxKNhVvWPhx2KWub3CXY
DYm6hWChJ20Z+Pz5IF33A/4PKt9opmuhgYpSbUxtvdHH/6c8B8N1upsDNRtKgcyA
pxC0p2WxbSnjTT3rXL/jYvcW0rZQCKRRH0W/zsqv2BYUxOWyDmTkeNJv9BRDlGmy
N24oTk5QRIKRWnuFTFbJo2ZUKmYTOs5biL19p4GwXouaJmrJ2TmdgSaPR+pXAUb8
ODYWQGl6N9sAsld9Qm8eMET6c2FJQRrtozXML0T8+OyCUkTxWa451iKxRy73lq6x
ZEgNkGCmvu1t1eKXZL3tCGkT4XaHifXSNh/MH4Vh7gdwB2ofkkFU/4+GY1cU0d+6
ITREAHNfk35fKzaETDtynkDB3Tg1Y5sWZoKBQ6MvqlpQGFyqcLfdEJUJ17vvPy6j
guIBegLNu6k72V4/x9WSQX9/j6neuc8kfrbUtwqpfK94HtxKEmIvE2/YsqWiLVKr
lw/jwnQfTulX12w52gtTvim5OBRCIXYwAB+1eYr6cS25dRHy/nnC0an62QynAOgj
Vn0+7FtgBL2zQ+8sy9k4Kvd2d2xLTdZBM+srKxgfBMp6cBHHh2CjRKpv98f35FAU
McV5POk1uL4/9L6ZwyEDE7zeeq0GA9JiL45KL0Vl4c8/MeNsKGhvOFqpeTHWLNYS
zcYMFkGxrebbTnqhxv5xaBv81ADhi5ukr1ZzKJNivO4Pbe/l+fZnOSrs0P9GZCGg
rj40bcxsqDB+tKusM2KWtDAyWA2TSU5sT3wQX8et8uNIR8a8lyllpC6ktJF5Ovc/
zkWCJ/4/GNktKdoW3vG3jsCbUz+6p19eZOFlYIbBQgZBeZZx4DvEE9rSnR2TMoRh
c6MYgSomQBGR/9KKS52gKx0We7CU4UrSXGV9tTK/n5WpKmXtIDI5eiSeo01sSjcD
NYd0TcDbMpBECYJGDYBskDzdgkE3QOux/zApdyoYSKyGCg6ayarL+SJRCxvmht+R
nRcGNp20T9P5kJma3L8HoUgv1H/aW7JmMw8pzyjPaOzPOuBXa5azcP79NT41rPAX
d3wMUoDmRs5/4YbEEnnxvevLurQNaL2TpbwdXuP/hpWZptO8fLBWOvv2rxUKYAVm
aie94CefHVGDGQb9ddtSUMrNVBzELNDytfxHQ3TfSqWEBSnWulPuxHliRKEY35R3
FU3oqwP4p3TzJ11CrEmQA78A7SxPDMsGUM9EC40Rs2VS83QO9jYa45CFgxzUkih9
CrIPBvi0kO3oJDnHwmo7X/IU4Kh9cHuhbIxtZq+SIdsKdeyO51Ood5Z6mi0/grba
Qc2SSijHJLoeFJV983rQ4XITppaHJk2MbhKqX+hJa+YquQ71vdenIj/gdkz2Y3O9
Wz/gSXXJR8iLZ1JGm18QbQr1GKB/NQ/27x/+4mmlt8OIBFs/BxdDLCMXcjtp5LDd
dz+ZiIhUIqfwsK30rpifh0HINuQY0OfHDr7L96KSaTkWE2f4OLeDGPb0VqfyIqzO
n4mhO7z0ava2+wCvVA00wAsPCMoOeVHYzamllYNUsuxWuvveTeFWDzAwu5GDlCZd
aPVwulUAVO48HKFbi9PfcwAQJ6+Zhl7SQcwsSeC/oq/Oue3vy9c32beXQAFH64eY
0wep4GO1SqNpTnEtAf55gWaHrgmnl3+eyS9ZZXGBgOQNzk+0xbEuNXnL4Xo3Pi4T
HmqXP5LaWKmCevK/Ipmz1ILt1wfKKxmiTsuHYlR0UnnsO35ulN08uHD0DX3JIuVI
1PqgA3UhRDiRFf9mjZ3gZYMPvGdCQ5a31CoAIes9UXQlaEwvAsxRwnoSKNIQClvC
y+D0rTPr9zusBG4Dsu8DJ9Xo8I8UCXeM8fo/lCZvy3H3Z0HNFhhohxyFJTpQQzLR
dnNfUYhUp08Wobu90OaizvKx/XT6SnCe6XtkIKE9TF/oX5revXl2lssGfd0RWDW+
QT1yu56gxvlPtoVPNJmALgiAaiB/6xLKpw/T7KACc0CKKijURp+vsSVoDwDYUCCn
sgVkYJyq7MPra1ROixyCdVvd8WAm/TQtBRmvciBmjovChSg+p89WisVAuIvA6oPM
D5SwfLMU+mEwNEYUD6gEAypRPAWbFMD1f5iqt+pzeCMVrFvea/w558C3KIqOz0vu
8OwTtsJtUqgcqIoGRvoCy6lQ67xlMZdkLU5p+NM6XInXVZqcuU/rNS8S38kaNhhT
EbX1RF8ig38jTatYNuOpww3e/5qaurk8ffkXCQSXhM8zMQD+FVgbUDwzZLjMKOsb
CRciERiwFENXbS5nVFeSlRjrJddUO13ZX53/siBgfNYNMrsBRtJNNLB2s236LeiW
WKgJUeKrdLyEh3d36EDS5uRNiGhS5GljbL1GHc+2ZbCAyqtfwT01YVpOXY5A1Z34
NbAn97ml9tnQveHAxVTo5Af3SvEzdEPWJ/aFJiSTYgQOjQBQoQe+vm5uGSlRsNTc
gytfP3dzi6Om6OdKCeaZ9xXk/n49STvGHInd9ukLQvgHBmkp9GcG+8ZvZ9MY+Muh
3iaoJoXYSBVFnOsAWpEStWL2y5ZtL+JSEC7J2wlpOESgTA1O8q4w0ntu95JdwlKJ
QVsubtglm7zQltH8yxjEwOaiaBfzQCabfABTE9+LE4zTpdiqCn09KYn56THjnOLa
U/wutECwVSvrCNz9aOpcmoZdKVtgWL7YuPYWQlMdWh53QlyvDuna23NPRKSn1nTu
omEHv03BYHA/GbORZCWi/Z0M3sgDNv3OmyCJ2Dka6ucNtKj6Mm6j6Id7RTkY8u8p
w8Z4vxwWu/e13bzEBhUh/GtJ2OuGVIwj1aZL/GCFoJB4GO8M/34RDJXV8QyDaQpN
EPuUC3g88e7OkD9gb3p93zLggwoBaxkTRrt5+9oGarka8xLdoBlrfwC9KM+uyIWY
5kBuXA5k2kzZFvXGnxZv4obUepVm+QjM6HluCme7j3sY9dIkz6vm4rEVKIupQthD
mvHYwj1N4UmKl9ox+9iI3vB9VM65lHKVTHquoLR7WaA9sY9u4dbjo14vy/lNOLQv
dmZFWz8lpn1JKmpN8h5DOeD41w/VcuuykILXYbQqIecpHHLkcDAOapIJx8cv0gi+
X9Oj5K9q/FeYRlacmkTRN4Me1PL9UTmXo9Vm7Zp/VbsIjGoht4zF2CE0QWbEL9kl
GX540yV/P5cbnXe1/vX7HOp2GdXTXeKpWrURrL6zAkvDNPopoTbWfEz6jxQr24PO
XK7D7vqXQtFlU34IREVGbErvIGwr9x5CBTmJ8z5wPeonbmdkHPEF5crHGxXzImpm
hmsze4u1jWcgucHqKV2hzhxdOHMhGs/AYS+iodCJ2XBt9Fo2bh+Ag+r/WHiscEK5
RXlSXRm/nOgDt5K/JOSTRlfdxdIGfmQ5h/ELb17rIUfNuNUlZks11Wkkkt1HbFA8
LSxCMFtvzJJJIhZEC0M3+IEeKUA3gEI0J887Ac1dVXWxbVF7pgXAJh7clSxH+eJD
CGDggkN9P/4q4CdqTa7p81c3yX4z/oStFEHKJiEiMyC2Tz0st9agYV2EKxNJaQmG
LXEkdG63RsZJI4Yipx3eknH5rSuZGSup/doSnCiJ1CoH6i5v/d7RkEH6RcgmvTLz
2Hn4N5GUEg/49niEv12ulEgC10cxhOwj4GfGpXw0TkbVrYcjWNcvQMqQIYgbQWpf
ttnsXZHcnBeAvQ/sEHC/XzLJJ4bk/9fOAx9F0hJRiVJ6WVtma/wrAevwyKfqytVT
zkpit5DNgsumoP1+eLdCJ9Wk8+K782z8teCWnlSee+Em/8pOKYa+zfED6/o02Eti
HBj7BYGuvVs5iY/dNV0EUDEl3Cb3G1UCKAo7afc+pzVTdpglNPrEOcCvmic467Kv
nmGTv5LZ1Et1yzz/3UT0q72ITVxxL14SkNCUK2fkzo42Eq5hp5W+qbaa/dpECt3u
f3g2+Vm24ubq6E6t7tUXFE1qqo1/CrYEPhwaJg1UtIKxyy0o4yyGBFXsM/JO+thr
MY6pm6LvoC4MWq16RQTKts0s3gaEFG6kuoMgHOgezcCJntyEzSrKeBx4fGcnVw/M
0JkmYJqAYRWiozIQrGm4WNRqGwJpMVrV2cN0kY6yTsgGk6lQXVuIK3IbgqP2wZ0J
Cak/DfCLPk24CNswaFJU+d3D7krEqtpMCNN1eFFvgK9hANfyVGDwYzrRiKaIw5+H
TszVd6roJ7d6nZLqmOOLezC77sq9beYJUh485UQbVZKf5z4cWIsK+hAIyHKHXG+g
GePrH73y0gfrFcHIl9NOzcyTTOmgDCKiHuh1dpcYvV0jiL+UHjaGwJwsIPlzH35w
t7Pd28yVwdW6kE44mq+Ic5IW9DcCPPVafglmzfihzej0IKBWPrr1w3itycbW7f4R
293wtuqTc3+m9Zaz7ccftfxr8JUWBOEMeSiEaExIfpa7tBrV3cPB5HrWrXeFJCMS
VTfSdP97ZFcFPBhsjPah5vfskwcYw2h4Ld10w/7vX4JMgDej3umrIFkX/krQzj+b
i1GLENYVfkdD6oF+rvra9/mx5wyz4VEutllnHRflBkyY+PsVJorBsBXhi4PdAivj
U6LxHiMr3/txxn7m8PQ6B2wrcdNHK/dchNVO14IeCg7iTyfiHqjEMAREYrgo/pLh
sqZLjKkS2kiYR5+16jXjQkp1nl3IDw+fphGnAOeWKl9x83Y2fV3FcvTKzWA61jd5
+7udTtv2W6iB8pfviWrOd14DwpiLkin9wc126biRk9ury+4HfQFNxGDeC8eKCXsu
waFsZaD8++U5dlznqDXw89+X7fzL9jdsnW3qx2ynhICQXjwAJo5XnsJfmaxwUC6i
7kpnzx26Ga4OCsVI8SFb39IPbzj+BgCpqrsNITXydUtyEJ+Db40pkJpYXUcjGQ59
BFHHB0fYooue9+uyiGeErkIEmmHe6V0/HFIixHtl1uVviOxm2DCGCOViUjsMt61a
Z/1UzJDMxIGUSEqeupeOOkAbQD1SSg0aG9GwJo+zJsiYHKgVKEKhPBLziLcRQHQD
nM4+T5Vac37fl9uGYb6PWhJr9AUhRvR9ZNeTmrV14z2im5VPAJ3Vi3dmB2rpCUtx
llmW1fpYD/cXW2JIuuaYgJKB9D0jsmtja3ydTsfz2YzX2kjkCvc/oe30Qkfhz7eV
o3j+bTIeP9PnuZRq5I/SRoN9gIgx7OVFulbsvTLwyZ4gan3LVxSJm6IP8LiYAr5U
hnZnRbWO2ZBzugXsfc/lpavGv7t37tFxHWrc8cRtyVJK3seDhSBD/oYqLFFEM+es
OrQ3mF0h5zFYJUotXy8y9aWv/K7V0J30/o6oK67AaOwJk5H8PMNr5ozR4hnRtm6k
YjI7S3PhxUcM5L1+VrxYk/5u+BdCn+EonYt/dXiTKcvJRnlyqsg9Xe+i1bsHjj5p
3lllO/XcbmY2rAf7EGAmf01PcYX2josuQVV4R+gnnriuNiWSKSELv04ZCcV9KChr
8duHMl6/StbJbTfgUxpMn0Cfq3cCwcsptCmWXeFjNMKF7aqs6kR61sXEf61lz3wI
E4zfKOFtGyBczCioqW/BP/YzDYOxuCYfV9i092kMysesBUP/6y4k3CqKiQbNUjlE
Ssh1yB/jaUqNfBaeRGSXpBUYkHxKlS95cXZP2KcmuXl6jiCFmvtRj6WmxZ1Fwqkc
awgejsSK5k6PJwZ1gDBrApuyz/YuRZuKLsrKopoXyp0zH5sQDZl7Oj6JrBNPy/xj
ZCRs0555KiHPHUC/g8/ojeeMbWoZouIfCI8TeXAkT47Af5KUsucESPq1T4Wnk0t3
8/l6SV33mqBulf2uP2v8SatvpPrq1GvV7sU2hOgbbBNL3DnYQJREbcDdLES0Z1RP
hTATjcF/r7c1D+vZPhX34y6iUpJbVqxB+qHwCPR481F//bQ0ELKTsGEzV2iQ3qoi
GyUF4t5H50GUVdG07wq8WsjVOynqsMqNc44CuWLipIV0Evvxt2W5HGP7Vo5jjR8o
mKhtjby1BKNhGYzmZYGdia51CI2wtTatYBN67vTjOmpBn9PFicbJpMo5tP1Xom8a
bzPDX5bFQhClwWgZdA1gZiKFJZUiZVnU7lXdrXvTJk0vINPfKMzXfARDH58AMrz7
3jvKFhCpzfQoQS1oobWjEO0pR223z1ZiuRS0IPIxOTLHKhimUFeVDmU/Shfoi6cc
SM/zQxV854k/WT/bomSFab9FCzcbV6cMf0XJjq5U11+Y+IEpdObkSXgqNsyQi05T
LzwWQQTS4SAgdYBB/v7CWUu6CplMZHycJ4h9+K0aq+R1Vlw28MzTsxzJzuWdJNGp
0vjc5Co8d5eruHhwNn3g4NubeQl/XpUMlCBcczML4zsLjvkfDwQ+JhHQuEseQBQe
XnEPNQD2g+2ovlAYKKPIzZp4+4ZaVLUnJrRJ8NEU6wN5qKQssZ6Lfx2vu09Bw+68
dTwZQG28CyAtw4sSqGJ2OtVx4GRk52C5R7oMmbdSKyn01sLP6f4GJa7BR7B1wSew
YR05GvIHPQATD26DmAJdNgGQ/AVc2HukqjUN198Ot+2U6ou2FOn46k7yeDYRM9zb
WvF0tUULgwFH1mpY9LS21deeHTd2Fzyo/637MBBbt7+pFhIqE/QD0kB6GAW0tP+P
mGPTjQYIqRJm+LHZ+ILDO7JQxjGd579GGCsiG7ffGctJ+3Ny5qLjY4WLeb1uUqzd
sgP7PD2UGFXnSVH8CddpQzWZlHprni0w2RcuR2av/vT+gdM7hL4jpnbrEAgjywS2
12+F4rhhWfeETfiiTYXgOJiKE/F7b02E7fIcOvhK1UOcC/d2YuhmYENkv73lsUSz
vwnJARELc+K59hvheF8qsIoYCtWljyli7wqK30CUT/tubUxeDM85sLbOh97zNm4I
4t4M5ejsDel9FOU3SZx+2Pfwv2mmCwvPkjCWtN9svEWNwKBt8JieKkE+MU6dG4P2
pC+ea8eDcSc1N8lZRlkipsdlkLaAzYVNl08t7OaHaBUZinI8CuHwqO34uqSLpDty
MdJGOlUEL69rasOOJAG30h1UBjLV+ByKVELjBBK8cp8M4+6R5uMGn9biNCyBbEcD
YtLJGIzE8O4yXfWWgYcAIMlKQtlD20kP2gr51LtRMqH1FPwZGZ/c9ECTA4Lwk260
NmH9MzYyRD077oSe3wl+OOom5HgdiNzqHPmy3MSO4NPmU+cuy7jrMXsU44a1dbMY
cY+QX+iMZmOA19nOsKgV0/N+vO4oTGu47sQoH0RqnoaiuRxlQW8VxiiwGZF9PK/u
63xlUhxKjbpACccaXsvx3InZ8icY9iImqNHtaVALgeepgHPJrAcllukE49HuYVWI
g6U/lJuVDSGVGIymbGoSfOUHyrCetWruOWWAKwoJF3Jher09Tel2RVLADZT6LK4k
nThTgrKwQsUm2csyELUIFdiizj5VS3r3HLOb3OQJ6QOpeT9dIB5qztQG/q314Neb
bas/jK2R2nWvKfF8jxbt1BhjyZP/DAlWNTPASSUGJKACWZroiFC41VGxrXuJkb0y
ZXN9B5/n2x8dA436bW+8hT8uYnCE+eCBgaJaq3q2jC7dtA1btGnHZ7eFAFPgs/cQ
Tom6D1ZXi5cVp35MTRs+yOAu9CJw1H8xf68ZplIf5/zu9Rc8oPGTwXulKpCuLk/V
QgqhGziUUnqKYpIUaZt9k9zLpIrCNEUCpxhfUd9++27AmTYqvBaCGBwWnMAL6gIY
IjbVa0TPAk697FEkRlCG6x18qW8DkdsROBB47Xe8l6hO+EwiU7tJNMrH4IO2NA7/
DcUmRgiSdip2tabd5Tl3yETekAGd9eciGDJUOovvsUxTMB1Epd+4nt764HgfE69Z
tHW4+YV2SrkLGn26vt7vAvl7w6NQ5FdUzop1IGh2tlZCGdWPy6svX97g2TR/wDoI
imsqWk40/4d8MfCff08IayhbDWyRZrAJq8xJijC1kWbyrXJOfH9z+jgKqqYxw0tF
W23986/quNzTncREERbyNsqmVnHHTOSt41D197BFFnkcWefF2t3Xix7s+ttC0zeB
CHAlowHbvUSrsdZLlb1FTPnU04KcubvKgT5HynDnXSaj+CxeIrMK2IUQp3hgmbB7
Fcyh/IdzSDcZE01nK2q7pfD1lKfN2qMZ3gsolF154feNlz/f/6LV4JQedUZy2hij
q2RgDC7sBwj2uXID6bAhZESO5j5j8JlFH42yg8jC+Kme5c2x4Q7lfqwdHyY2A//w
lsldyGFvguONRK3dPa4cW91+846PuHSR7PmzYTnweaeeMS8ujMREAWC7drlIEQMd
bBguIYNZJKurEbZtrRXayAAAvkONWQYYln6RIdreKSTYfJN8lX+zzfMHWNe3nKrJ
9ARX632ccv+n9js+Lzzroa46k9XrpO5NziZewoeC9jXkaY6/qcb3ljWGbBX6bzXV
9hUMUpOtEB2AbkoW0A9SpjseIoITGaOC3SonXjfqubzAnriVKoD/udf3IsvswymL
9V34abpVUucrnbRYi/DQY2TdDfY52mqQD1P0awB4EbNNdXjZyfVvs/tDEbTIe9J4
EJup65L7gIUehUEdPLvbgVvIob7GcHYdURIYwSHwWLYfNaaU+6vjju35rml9BGhi
uhpfejGPOMRqr7e3QibMuRzRoeCgbY8PpeKAuLLDZjhL6EXOgZA235hz+OhM4Jny
yQjRuMi/HKCQRS/ImluXIb3Zh49bSmayX/4ISkuNLilqJRqRMi+L4N5w5SSikn+G
+sYZjqgfHf7ZAXTxHDH1RXCOWIRn1WvoxmXJow8lrqQJw6xXYwTz+YfpAduVD098
BbOf3s9RdDX9CJf7t+foh/iyhqiT/RMi5X+ds4M+RrIGmiBfC7nfv6j/t4TR6tVE
thZLZ21UyW2S+pO2vLfCMk5gSjt8lQqtgqoe1vQkq3MRJRZoQC+f9p9TM71JJVpS
8B+WQ1BZkB/kPh19fcKESZWmP4e4GP4oxIY0yJ+uL9KGl3ooCvCZZik0x3eDhgNJ
tYW35VDaQLG+UFvivSgSRAbbnSPQa1gfo6ETSfDancCxQv+ouRR0rE6vsihXo8xf
UZR+dbfmKr4gZ9PpsfTAahtGU0pSIv1wMeq1gleYQvcSUnJUpCXd2LVDN1+z2URx
WfJQY+lOGLmemFVBqKC+pupGHNKrhS2WsWwTtNoK5O/58+53yDt7TYKnB7WCO0uI
acWD0HKouXzYkK5tg7zrgtGJcw29Pg0TQik7u2h++FLDVet3ZfvbUCC9CT0Fk+2T
L2vBBToutxmZFS/wUQDXgxxuxwUUHGpSXkU/c8qjCOjDKoxRhdLgFp0WhLhbY10+
484x/DvzCBeXwevolhElM4NfY+A1tuqjspG4a1h/4MHcG/6dttpRlrV/eTOkhLhR
tLdCSk/4fi32jW6bKRo9HdATGGxEsTVrrA+zIYL5L0O2tPn7coemkZ05IoHngvoq
dRQfP7cfsfXihmOKO6A+8BPxIOTpQZcc4as5HbyFliZ507WBakl00sXUjuz+it/F
W1rDhcUH6mCnON0Z88zk5GCZqBviP7h35zRYVzM20nrPPUOw6R/KcnnjAMeMKT/I
nZO920v1Yh0H7f2h0rrbxrRzQ4M7Z5eF8Emi+LktJSYqL9TD3hUeKuyTl7LNEpux
MesvlSnjME61PwfjuPl11v6RXeahjL9YxcsKH0DmmUvKstAasP5T8UlozmXDX2di
/V9jCVO5ltpKS4EJxxuyyWI/asDz9A1WQ8DDJgx9s7Egh444TZMU18c6/cCqaUc1
Izpd+EHWzWrLn2rjIAyZne5pkReF2YKMWCCOa3Oc5j0tkUI3qtH339TzwutDZztt
HGnaWyWArZ/OOQXWS5tHTj5PGT0IAOu8lyHLrhGfL+rQSL3o/U93tALt/UHkqkK2
KS5Pgzkpwwgst1BJfpORz/d4TzCGe2s3Wop+HIJyCHvuk44MmmDQyy5zChnLwE36
bY5qXUYv5DOLJTuTHqdiGwVNKX7jmPpSVDNtgWZHkwH5cE+XOZ3n+/+08OAB09d+
VlNJStqH+5EeBJL4+SxC+zHjNP1Br3+goYfPysx+ZqHx+ZqBRF70R7I9fRNVEEN/
TzWgmPFL1lmv+ZYA0zl4kkA4zMB2HTBIBayy7BNPxhEjB00RBeEnDtmt+mAnRrwH
kdNnQ4UbZBCZozHwExcEky6xmPwLqVy6hqOnOATVWe/+aIlU9YQMTRvcUxZAJO4Q
LsH391NeImsi+mDagEsBGx0RPbhVLYMoaZWW5eQlspcQwh9fCD7h8jUMiV4H1ZH4
fBgWVuJbQbR7Upqgkf0+2+P2Zgl+nvoYG4niOeg5CyK2ySjSQJjtXd/wp7iqXjJH
G/I/85/XKwSSqQvlm87845ttVGCNNklgUWPQwH6ywgrZGwarMXlOZzmodZd0cmUB
TR+hlrUmiRX3YzFrV21VzWJswoR6AJByygk4F7ycIM9EmFEISzCF3Xn8/UPD9QK4
uYAUEEmga7gwXLimWg0F0fRNbE/i8zzbgm/b6LqueGdeLMel5oM2Uk0JKnU+qLqY
SFKgK0se6zCxQxl61e0BWXM73nXrLVE0ohfdBP+0NYHUcTDFSuRR76k1qkSzxQfA
vQ4Use2KNGZ7Y0xN9OtgxcMNACs/+LNlqsI1Ld1B1dZ9Whb1B0ARuYEPh8TrOjkA
y2WPS9sqWNUnfehM/4Bsk0vm/E3d9oBmckcDcM+ygxQbQCWD/xQNURslBBHJnYRc
Tk0/WVeXG+3eZ1nspsqksdTCRijITykDFXN6d20KoOiJo7Laui0tGqVY9K5BSJfj
s00Pfwgi59G3OsopqPgElJRz3ww3pMHawZ/udHnaAnVSgoNf86USwy14yc1zmBcn
BTmbsztYW5myaxq7RdaGNuRU62SeJtXbsY3NIvgkQWos0mdHSNg9O+TIbaJ3it3t
VULDX83CK3p4mS+HFGt8pv+YgZ5RDJHBieKSCylWA4nJdbe7f3AVILNt6fVaFJiO
HAcb2JVgVahDKJVJ8xIs6BZjLhgvnNFJULK8LsILjwq9JF1wphNVjWIOTnDMMLWa
7SGekUHsR3hsCd2tBDeKIE0jFHvglt3nTcM2XucKNWrTEjNWh61SQGhFgNjx+f1z
X4Cu4SA176IWFkzf/ZiYWFuk/3JtSi2mvPY/RJ+PIBgpeurB56egoS8rsk2yBUve
8Jv69Owz7ShFGVz+Lb17KMKUR8b1vi9ZUljPTO88gbtvgk6BKSAralbyRW7zfRgb
ojJH4XsMmil++WYLgBbL0v7QA2FfOWIeCBwVFu8GZaj4Y7dvj43Owk9sKGekxvIM
pINJ18NM8G3fBOXd5hw1qPfCMRiaS3USI88G1UB/J30gZNYs2LZYC9EXPngU8wVu
i/eVUXnBSSVAIJ+tbREj1JTC1fEVRC0efn8iLzzSjY4TkMFFcz0HrHecOzHCi2ws
CfyAeei8wASE89ptGNGrCJ6NWMuOuUqcJyP+9hDrxSeQqbASkp8xHga3bK/dCjin
vQz4fQ+Ja97v7YGw2Re6bLfDpLfifDox4Nt1plVJuVQLl9DVwbxZ8dOZ1R5+n+jd
1o9X8EMyQLQvBkqYvmSWI9teok0HVF8kPTq+ntVFwgHoLJWstpyKYmkhtoucb/c0
AuUDbCBrjU8tLU/URM8fUgdVFrvL3e4F5SC6XRNRCao4adR6QDIkyw19GTcCvQOU
q2tvHOEccuf0pRwgI7qnWKUU1PVHYml7L0Yi94dgtVfzO1IwOJynC42xClg7q9io
BevRsaDzmEORDi0n7PeYLzeLkaazqTpfscxfNexULOYzGDfqA1yr9KSdW/z55xxd
/4qx3tK/+nx0GapD8Em09zwlKuQ2i4ccl143uNNBf+dkIyKZfiHvyC3Hfgcba6DW
kCZVaUrzh3oDypsP8Rl1/q/r2I1zLCKXuAJna/fxdz26lzzosYdWWpY68QHifJFN
K9umIKn0ThVCTidHJSPpK9hBKgan2D94Cr+108jzUbZzry9ybuHDUy5je/Mb6Cgr
xCF1sBoSb1lvLMh88ZE2+TOTvriuLt+q2Pzp4ig5MqjIu5MfyDudDvnZ6BPHPyP7
TflvvO4Pxr4UJbTlUIGAf0x5FAvElkLMwgjsQD0soMvcRt9Ln/r1At21tvP4Xo25
eSttxs7wSOPnFXYS2oLqEyDHrIgO5No4tph9ATW39WiDX3kdNirLF5zot47CVcBS
KpkeZB7ve7faak+lx9EKNPLY0B3YehjDTCedG91fwQZv41cm8QqeUcO7RgqO2gch
iin1z8xiw6Zos3btzDJTKsGyVn9gOj2BB3cS+fnB/YPrkB77BY9HJ6eSHHIUyygY
idcA3xNd0d2hJdA2rGcxigAF7pgB+zmhTiAOfObFok/sZaccVGmUpcpW+u0/f+Jp
7TOkfyCCPxUALtwE2ipVc4RJjEVjZ3b+WZAt0dF8tw+v1GXgm/A0WwZEfQ39yguU
sD2GvegiX5fWV5F4OPXXkPPNYBOFAkTgyYAYcDSTY5QnsArRIRGQuNoFSgDh/HrX
AcHAZVT9jKMeevMTQYC7MdGR8Os4bvcIw/rqTBDo64JElbp1A0+hNQPPSi4WjXNa
OWZ9JAVwVCPH0fO8DsmEoUbUFwTx6mexmpdnSL+mm0IbrJ50ZYnTjgqftxx+hj34
RF9/yGA0Jagoof0XhwA6TT9yT1HXbLpBN376aKvbhFHUWo/HVz9bwH/u+qYVlPFR
ix9K5MiYi5blOh6oBg9FEbaOTZGQZ+klyJwZLYcIoSvOC2J701zf2JQcxFsKeKZy
GfCk/OZrLzWzs6pp91QIcjp/SNvZORz79Y8tC6lSkShTLxj4rKz5kDluevo7mHIO
fM4T4UbEqyJsmu0zLVUN5XpvDYg/Yt70BcAcgdHewSJr8Fz2R7FqmbLKp+VMpaIK
jCbSWRz93+DKpzofuFYv/y8LdoiWa+Rt+k8PcZniR44CxsLaqnaDJDGZ+L2xPHCM
Ic9myeeG6fOPdfPcRBbByUpiBxvdqcAp8SVOj58BchdAbE5FLRFL6OZQCco1Czb8
mDCu/ZhUK42TGbetv9jXhOR1aYS7rD3e+5lvIeGFTnR4Tba0XQ+9xeGX6fer87fQ
VPtY21MtOfDJR2phV3YIJp/lG/SQntGOTzv2PF619K+XkHrsrOKwsXyzOgWdCuLq
ZiPSAXEW+l1AvoTEOQvWiG1d317vhhU24cN3L+GDqhbfynm6qpOzSPujwk5nR4oE
PpizvQc/H9uiKjn8cQstFjRyDuZ3+zFHswgAAeoPRxCSEjUPomrKx+Y2JBypyvBn
9Ir76tYRKuVu4PjcalndYObiHLwDGxqdlV5wk21rEsajO4K1uDBNQtQoUrl+MVks
k4zNntKeWljpGdEGcoEq3Axz0B+GEEymyjvov4zSmKa5RYSL4bHFMhqHk2PD+cyk
6lZScacBoO80vSjxCb6/xe0l2R208stFspom9QLR4EruH6NtDuvGz0nEnQte62J0
sePeTrrru/6ddHX88aK88EjICikITrLK8NWCijv1UY8VoBFPMqW1i3fZDQKgx4Lt
kN2toi4PXEZTL5y7wNoyZghydtrGaKAzZX69VPzdT+GW+8KZnFeGfVFmfivhEdec
R9bqGBBOhOAKDEf++IMit5UwVBsdAkh2TCbpHGWzPVqubtdNkkn9agzuAoY3HHzS
zZwx772lFG/048inhb6+FXU1ogdaLEizP1nLOPE+APTVN19+5Z2AgcZE1uUZob6m
QsgkRCmv3z5izF46uaf9HTLz8sn65Qspyh/IRMJ6z7jwHE4PMSMpUsPRFisvdYqp
FDm/RBNoOfbDCnaF2170UVbi1Gov9Vtx14f0xt12PWP6QMH+4f6zIM7HTZimO9Za
EF/4c8XhUAde9WWuM95BQm3IRQBQ6NCurr/wou9/Rz5gJ4PNB0+cL5OkgV90yXE8
An6WqJ6k4XaWxsjoMe/82a9zvKBD36gSLeSMRQJKmNqKhrck5arPXFJEitrsdMW3
Y4xCw8tTWgsNLt51Zh0hh3EyzliCe4xKOheyhz6QGnIiHlLFBWiyB8+XGCRmDBEE
+Ta1ZPdI5Eq06yAk1EASx97uEKAhduQfAgrF5khbLRHvuHuwZOoz+mSJ/JxH2/Cg
ZrvJ4hBfYYK7H9AVMRwiOQwgvB1ATTD71jRB6OqXFT+jSGltVdCFe76Q03dgw/Dx
a5m97dlvKUCAs6b42gzmWTOfF002DvaHguw4yKpIBfIyDa+UCxkocljKbm++iqCQ
L9hvQo4iIvcQ7r6B14THklyBZ4Aai27GHhkUvBhqA1VhR+bDsJQQKVN4yAeCBubq
rHdvt6C29NU4jkWlCF/cSOaKQ9/r7XLCXtQCsCzcCf6sFbtMl6SvyDWhpO0lLTNY
yWb/oXzchd0Sq1DKuBE9AKgDKo6tyPD/ymvQ8zTZb8auCMISUfCS4Sof2X3b42Ct
q1/9JY0QG/dU/Y9ZXgyNXeIzWUa+vQYHgiBz7kRFCdxDLa88JKq+uL0HhWhm6713
HAeL2b3V4eUkMshVNosct79DYWWFq+f/Y5JdTDfCol/TwXiLRHaD1xxFrJ8UQkR+
UaT2nem8f+Ukr24MspAow3WFY5h3Dt3WOc79sLb5u2rY9SyzBpmuzssyAoOfcvIS
j619Wq8OlQUgl4UjdxvhxPfC3nE9VmN52QRYzmdOgzZfcRNmYRv9lVEBGoMzR+JF
WkSjqfjgxPKSCzrMiARsuQDdpZKvi4w8rSy4HZtPJkndA9mgPwQkbVRfaiJz3j9J
O1mg4nvqAcuw69/47U8bxtv1EKbIqAGiZYWm+Y46wVbbgSSTeK5Upf6FmfdytnLa
DzgUnPLfYRsnteSbk33KWCAlI6Hi2gSyWx1IamgKFVszoSXBR9i2m46wlXDw725N
gdBhw9FNiKr5gwMrY2eV0kIgmOuXXDkdIipsuSd75FeknX4GYyn1OUXbK7Aovtfs
pJ6XT93ECa4vWFo+cqbrtXH2UmiLLhp964cukxDdix1cjYyc3Txn9To4G/KNr0Qj
sTJhzs2fpjUSHqGkt4xpKvSH1Mw1pWyrOpdpyFOL2ECixV3ndhuw7VFKaDSJYWiO
TKUjQ7tnavqjRR4lxfz9YBZhX/OKIn4smdKkYL5NsUrun+NihKsBmmXI7fRZUoV8
MuroroFJPBY8U0ednNaomDpuXkXgyTWzGnZKDDXoDPlf2YrjLr9/G573NkFEaO4R
L8dHM31/Pr/BmZW5ZvpnpgkxPQh7ftBn2PrmxqeQkwhlRtNuRXvdvzNqR5ToBxlp
eT2E4ikouXiJ6CUFFe4d2qaIqE38aySZKx62O5aB0+I37mQ2bmSmSQrwtUC5a2P+
6j2CDS+qRtJnZ3lzsUpOQb1/0nVR9BmKL7InjhrKFVXsxXHKCmnIpQjMZ7NXFpa/
8eURafDdvXvI+j8lUv9HhR4HFeQ0j9zYxJ1tE8r2/eQhHd1TqATICDQIVkyeD6jZ
9OGij94ULjZ4WjIN/iIcWEPsPIwQPn7JN9FSc+tHyM+QckjiXcpBPobQnpj7+Ftf
oD8CXKsDD83vpDn2YmKhfeTvhpiVEwqlPQIsz86i3I3dbms9qgVvQ4O3yduWzBhS
zGcG3QQs+Y8+ZLHM/9Pcqy0U/3A0lj/pfCDZFUz0FmUQKfi3Et1L3l96ooOl6fV6
/aT65BQ7lEL+2771h6A1P6ZZynZ1Yfx/wEr1sR4s5huR0uakbMd4DTgl0ByPR/f0
Ewyok4nw+Ze8XeHdfFcM/NeNXo4D+721BoiVl4p4UgnGsur8RLp4TBKydfRqZLvm
LcFj0BAocdd8Xc3B+unK8qAvka+2QpQO/UgjuoSUdaMbaGkNwch3RISF7UlUd8YT
IgaPynhYzqP0y+7Ko4npKCNClMo6TOr2CGdXs5OJUK4rmZDHtwmqAEjuFiKDtMt3
y4Xuv4Yu/Jhk0wK+ATtGwejltKppUTyNaTbnbSU4mPDSJgX/JhvVv0Rubpm9LuXH
l2/0KsvH4QPRBKx3frnVd/T7J5h4pPA8LuaPt1ieRKyuFDFYu9+HbiNxUTyKPBGR
Fugpk1GKRnDPK+OWuE2H8wUnCir2yIrgtlYdH9HgV5ECcUuqwloU42XrKyvY4cT0
o5L9+OpSaQttfCZzx4iE6rS66V2Tf+1/Z8maVHhf9K1OP7ogajNiUcAhkMIj0hmo
bmx1gXgpyYKA8fodERHL+jNOSQYqVYCYAuQL4ehCLLg3xD/yIS43yKrUc551Rq1S
+PbFOl3tyD82QzXdWmNPRvrGJEvQn5/2dIyhc5yByOINdpvmH5n/2WTc+jdF/zGD
hlrOwUOfoLz0+8sgnbDc6pzFbFxkvw8cjUzo2/Xpa2sotQYsouWm335ExazafFrk
sp2k7uLEaSCtQ5LXO/n/XPJT/PVa2xedaYN+FcDtSAXuUomx/lNZp0ZU5BVdikiY
iQv+ItHzGsimSMdJdInHV3aEub/W0Rr69ZGvZ/RtEmDRU/dzAvSSnIxNexsdK3rz
AO+3tebhaLM+97cvDG9NM/LYG9q4JdFtdVJBJEHZ033C+urb7RJbyYddKPZGiPBa
G0Xqe6EwXi1WfSTxeWBycrTtvAJbALKzOiyRB9p4En//QPNjNoaOrB/YkA30R6Kd
I3N7imkVsvQBxDNdekloeQTYFMpeRuUnIFq01nikVdM/GVJXK+OIDpsCddKW/OcT
pZr6QHd/0HQeGLFUV/DZME0612830Nqzkk2cCN/k48zcylY3njDIepN68fzqOvVn
xlMeoWGL/VvG9ZRs98NAsb/YyO7KeN1yAJ+p3zY06CPanbwV+alnKPqcllF65pg+
Q10eQpHF0GAtoLGKfzvL79I1FgaDZsV8c9nisqAWzJEEPXpEqKiBfNlYmRpaFcf+
Vtn0+0ehPvXewKk0/hHjG+XKyCDqOGJ5S6gB8UMjEnZz9rmL3qKpJAW4Hn6TVLjJ
EYBNCQevc4TadezzfthhC1oJsPlnDo8FliuRNOp8LV6WBu0Bkdi3piMub9rkVEB3
jPpNNNWgUK3++hV1c9eMIesikbsNOgubDnCNP2SJRn5sEh6DB79pihdXwvJGOd1q
DD358oBLWW3L5STQU5xuu4lMM6lDNBiNvehIxAzJnVL6nPvzgEGu29OBQvR83mzc
1OLl5iX4M+v62gryMF0CuUFE+7f28jpxcCOljwYYvx6Ibha1b+uju2FoLnNXFwM/
Nh0HQqF4xXdyktV7xkMYwVc3esxwhFcCWBJqI+UM6QbqZ6/xUhB+/le1QGleDo6B
/8wHER1nWOu+DWm2ceJ4f7PdYU5ThaVueVCrVzkm4ygO1OGBCa7XhIWlZn2YvJC4
CAIH5ZjpJ3m5GVw1rzkOLSFAJiqXkiqbx8E3qnze1Cv3oBQWUZw0PPuvFB7Rzhoc
aBXYDi0KHNFNFl4QRXORfHEMC0BiBBCXcKXQKG/78IcOyGkDdVGtV3ubGiqySB74
/o6PkJqueUC/MlUOh9HAmeeiP+hdYAzFMI+7ra8S1f0zkTeOLDyJs0iynwInJ3GI
XQc4F4LXlwl0h3x+ZDcEpbRzMI6oClIWSK2+qyQF2n4y51VKxYyC5AGSA+Etugx9
TZSYPGyTWOTB1v8khbHhzm9uMvpb3kDIO/6m1vbZGjC028FJnfQxmz+o6/wzIS1R
Ow8zMrsUf2L1c0Xc4NHJKbx+dA/uQ/oipYCwme5nFx+39iVNWXZQV22sAKvfFI8b
qWEceNiuZ4hKmISSukL2P7p8zTzTeyq6PtSvczYna4ebyfPzyrh5LYSYCR/i/ngm
aT/h51kcPsCy+I/tCILRdCzYokJMMsvgRbkszS+zlSp8dHzZNPRkTYFKdDm0TIgm
pbt9yG2kvwxCpF+NeOoV3qdKmZJj9nJ2L8ozo83stBW/sP1Dtqch97LeF5uy+hRQ
w6iGQ2tcDeHXE97eLr7uh9sdyKwim2ZlbAbv2IQLgIaTO9YreBVCqZNucoD0hl5S
DpTuh3Lgfltx0Hailr9sSmSw/5HrNLuAKMeSiT4o7I2WdmmLHRdaPSP05OqynF2y
CNsMVib5pPvwGhCmNxpmsv5FQSazGpY59TxLBXPKImgT4Urh8muhyrMAT4eB1kLc
cc4AkmRmXouGqAw3EHtIv1nIGoavGnQPbYSwmcUretZ4+QGAkj2KzHBBhxzrDJXr
47DCLBE2+gmoPUJGVpjNpR84pF8YvoqmuIxIS+FOtEJS8BYhwaQCTehlPpASD/uK
PnQtEshJUMplUEmD/+Y6+Xq7KtlBlh5HZVaJw/QASKqZ8Q5PX8bE7oefezQuUFuV
J43I2J3za13+9UQBXn+2QrWodpNphu9nnOq7Seo/N0Jr6hCq59G9NabY16HPcIIh
dKrgXvpiqRhm6oKgihurytwAaxgQkRvBSrkDfql2FbxLY5zNPDpkH+oeud7N++0G
R+Q9MKgQ7g0Vp8pdkckwzb95GK633os3fU2sM7gL1SkOElpURG21GkLTNk8AwkWy
lT5ahIBC/GToU7Wb9lZtOvxHgYuf6fohnLbb7S0RVlShJFfjl0jqawz9H+6cFKYx
7l3rpFgVkAVoRiEI3i5p6iXtenVUhcEw1gHjof3tQfj2RILOMSB1yANxS+ngSpWi
ocPZhEA/F9XlWipcHHS6+d3nc/yFyzBnSHFa1gDZhe5lFsJjiSLZ46Wp/btjA1e1
HezrU7X6Dzw9wxsEQftrzy4NlD/vRCNECQyYUl1djWD/+T/UBYaOCKMNKQf3zP4I
9bB+++KwzgU4h6dgFVifNVsKRfyxKVQJG9nPBEIOLI4GWn9503F1qtyGrNyBn5/F
NAX1p/ehcJQ91o0f2iQNRm5/252BrLZ5If6ZDWHfPDoJpKL+TZmWbPfFwVHvljsU
T7/T8upC1Db9tJnmNnBQGOrmtuEem786p23tcQO7H1VN8jxKJG2UqLauGShZC4Sv
8DX7BS0r6xXes5n4OucXUXUdBGwEVppyxTCUdgbDMTkqd/xknsvYIYBwcbhBg3L2
8ooWBp+0yrj5pBJYmQGOA8iu9iVknJd6VFgxflJcvjypHHQIi8ZckV4vu06b/iJN
2LS5B8oQydCA/v5P0S5i4zuaT/+8KnHdF7O12H+1CZu7qw0O8wE2ioJ7L6+kNEA3
BijouuAO/PBAtWCKbticyfQgWR0+N17/LvIsG5iIbQyB/p9lYSRFVRwns7fTffmF
SVrjk9eCXVw2AGCgBSPLsDOwnUwZX+pfOU5XHQhfgLancZJt9FXOmDhy+pp4HzIk
rzD2mRH0FU9HLCEJRrEUyCa6mNijG2DFNozWfjY6u7JLHTggY64Qfq8PwzyPKvuf
EcGAMtk8bpFOaK/eGNmAuOxZSfPNz4MNKr4nNdpqtP9wHIg98bzA+93A8RLBUTYw
AJax58oO8CQJxbQS5P6pDE1XBde3eniehP/ZpaFh4vfMvIW3vPeAjX19X6g3YDD5
kTlhWW8dFDLdonenF+9/yda4o4tLo/U23NtVdgDck9ZeqcA2ce4LnRhxTkQjm1L0
A8IuuJksu2NNJLBqz/MoKcG9WI2oEWEJkNrRDmzX6a9itML/DVtfqGx8gbrfKlVn
Nfdh4jHY43RjffDhQpSCIei5nn6fDLBlMFkAE01LfZL802yghbELUzEt25RKDa0b
ydjC11GMqUgEjEU6IYQCw6QBiYBUy00HeML7Vf++c8v3k7Zz2n6EEs/ekL99yaHA
tsZtQaeorkIEeZM/So2zZc7ceSsxvTmrZt3qoGpJE9rj5V2O/Bpck0KozKfqOjLW
HVjoUWtkt8OhLJvC7pi2tH+rsxPSA44Bda7arWnFaEy9cm/ES6uVjy7zU8+XqpA8
vpuUE/SsP/iTV8PYPNIPqaNmH98h+D+Z/g25OZHZT6jZhoIP/ytWjKI4N6/DYitN
zr/v+YF/ZCgCmDa7zkabY4rsLY7YnyEaiQ3kJdQW/65dYU5YhMKFT4od3LJVK2TN
BH0ul1z/4vUlpyNHRNLb5FDc+nwSD5pswDoVN3DyJcePGHYXxSfdBJjjvS2ncpUr
TWnqmmR9C04NFqeyTmu27GSV3HwIMRj6no1qpMusWFizEu6mrEe0M7boxDNJRlBB
JSpQ/f1BCYFgyMo5sfusuPXArppewNxwArUhjYkhsTtxtLoTrUFayZqHwIN5xJms
m5XvUltejZgUEsyFApKAJFOGRJDw65zkqhrMgVYaJGjLn55r5rBkSXnHbYVTaHWc
sHxd/mQrPoPlrWXfXu9P9P7efZ9IAgRhIMRlOVJTb3wUBTKBqs5H8OvpvXotMVB4
63juoWJRNHeS1AZch7y+BBnGYvUrJkVKR6vKWpiusNXpdQp8yUfbhiyvaLuE3Yd9
D1jEccAPx80FXK0z5KY7Z158FCVFUI+pLU9xlT39yyy+lt+jgWUpUB1ZiwKFzTob
g5aeV/OuP+IreJ4E1p4mhky3BWv5iCX5U+yk06IUaMguyVwVX6G6BsWNK3k6q0J9
eAqhPIcuFjVEPz3xg6pmrLTY3WOVYhnoEnj8W8osB4wgxw+axFybQbN531GSLyLo
KNun6YBvSBRZ0wG68PJWfrg9qn4cHUomUCX0bLLl8ebIV2eg+dNXftmBhux/8BpT
kRYUoqSncrNrLPs1XOICQUzuzQcMq2kM/LjIzWG08EH2oNU2Jo9XOC1kHsQmz59r
YsPCv/t4dLzR5/v/DytUPqJBahqBIO+LiTzlViyqMLL9+4kWZPqkNskkhoKoMkFc
pTVxSLW6alidkwYm9Rgs5m2aChF0ia9l2p8QjlnNN24CHy7cmONKatEliTE6zxCE
h7E8S0h7PovESnHXcDdL+2XHXb8M/EKxB5IOQvWMrHzhrT9uFhz3KH/hg8wHCNMQ
bK0Bn+pcT5bC8BbE0jvJflum9jr75MWMO9eyi0BVxx1SbrTymZ8kYCNjEnr7zgxZ
9Rd4dG+vubttHzSbGtV1Cba70Xg4vdpH3jyg4XfBbd/gQ3MkfuYIBGADZ5tLoUP1
+nln0tKP+iv5q64Bqxkaqig7mzH+e68lDaKSaeWV+dOewX0AKLxyBD+p2sU8zNAd
GRc66qzw22rYrGn84a0rLaF/kYb+y+6ntTz+kp83wkYq//ut9YX4PmDAoSysUsJ3
1yQ1r5ktT11HElIak6lGhyA4K7slN+AHsE84z/mbOwzzbrbO8HpC9biMlqEz1igx
pJrxKLjiOXkBKUrj32zYQwYBeeMIy+ssMRV8IkDW5jIcpFogDpa5UyUXHJAhMiTo
jy0yu4FdJDljjaSVfVMG/unHN+5nXaN52vR+4nr+M1cr6E4g85SAfcZcuEmi+Ljf
xhJg5ePThi0p3v7B1Hqcp6Dh1RYC0nYMUBfEGYnISfdUMzDaaafLS9pl5bUKBFWo
8ezpaA7+zOZdUnbMjOeJE5EEuqUOWrXOVg08lzVyO8p85RTo+TenSglAYCwCv+Ja
n62Zy8CmXrUaH0Hq56430OeUHSgKEqaiEDEmrJuxqRlyLDM06RH8aSzHndNH07qv
eyTpjo7Qf/nX3VGfF16jap1Nw3e9GBc9ZnAySNdTpyy4Dp3N2cGXWxUx04mK6QL/
utis2Vgf3klIpyazgC4KToG8EsDlxX9TLtD2QfaDiNp3nBfvJrWmssJTnzFQko/E
cp8PbxFtwXqjpic0os73jiE3b4rKq8BCT+haHZ4Ul9CS0Lp56iDfTnSRdwrW10j4
UIo2mjnrtxdc6JSPbOHy0RLv5msNTr9UhWM3FZWmEsoLqIRkmtRs50bYNgqYV82A
r9jAx2RI2BVjJJ4NsRAMs6i6XgbQu8pZvEV2NMivP1cUzsbS8x13MwcdleZgphAE
FDOmV9n45ICH4rqKopC6R05tLpDxeqiTmRJvVystpo/z+7h5THgL6Veln14Ur35B
ycZjQ4VJjoD0Vgba2m+MpWvLqiVtCq+bJHmhZ202HUwMx7JHUEiUH8Jp9adpuQCR
+H4an+UZWPBGVIqproxmfE0SrfeAKX2XGMVQTA4kvMdwUZudtseQd2fIxRwjVEgu
N/03UlKJEj+zNIpoUrA8Utj3RvFt0ozIKtR3m4H9RT36bZqHiO9jELLxwfV34aww
z1MeLVghyKqx1B6JVIc9DJbywrQeLY11h0sMJVB34OHvM4dq59hhEygf0PITPSfA
CQZoLU50D516r40bjUWd/QPontf3bBkgzBUW5hU4zE+OfDwH9mK2h1XnHZlgKvdc
xDZilcuUhZ9BFbKAzABiknxMR9nbQbHDOMPQxLpcNcGVtmQ/pDmwJ6FBNj/XMAHj
SRCfI/77ecKt8HqEXpH6WDARZIf6jDtx+5oAqhHRV2uHvD41DlUy1nl1mtOyD/Ph
ClsuTbngbzPHBQj0LYnOMZmPwLpOOi7a9ZWFlXUmPdFKPdQvIiy/NeczH7hOcJu8
m+8jzkp2eeLM4KQC00FExpvBwV535Lm/oxlSMtBlLvMJ+c2RDSJtKC5BrzLVnRjG
oz30ZHehRSBJg9ZAyYwz9qtPQtrVTv3EqPBvYbn62FmJwhOWjdGXGVGFehpNHEAU
44lJdKHcCOPEJR/lU5E3I8y7VINpgdYEYiDJtkEDXTkbPomDYI+KEq4PIoNhmDeo
u8PAQS0luFxDOmWpQ1+26/SYObyqF51wMKflxxDf8fiM41v/LnmwFZu19blLDeE3
XgKNWV9ZmVEj32S1f9VyM3CNR1R2P1j7edg/MlFtbOjV1Lwqp4ONVC8gab+/YHKl
+1VZyLs8NBuryIQ7KhqamCZPqo1ThYYWJaxuQ8av7zpVGrsTOGXddxW7PEcwphWX
Xbya8Gk1KUHelk/LgMGH73otaMzDdsvVD+DM6hEQhLgZPJ6iarGSe/q3nZYdTFBl
eDijl6iRckAYdxDENjniISHJ9EMjzawMefvttirjMmY6GePb9KCOtQlE+3oX6YXF
abLpDcVALtE0xXT3IKE3gWj1kDHITvwLz2Uac2a8FbhkQcTsdasswq1LnF/GXi/C
pDVr3I4d9/7nXHjVnLXw5d1e9BfWtbhFRBVAzEfCGUvCrt408hTw/ck7C1fL45yQ
da83EiGyB+GhGGCPryCUca3Gg9ft3LomgJopxyMaWv/QZL6ueENUveHFJrobbo8h
xrrmWzfmribuMAjIgfPEKeUVLoJVoviOD2zKlpuzewefzq/5xipJtwm+113kTzIe
vWmCYd73gdR6P7pl3YN9ZAWyWC2YU0bujB+ghrVBSnmLhp50np1EdH6mAUP55q07
ii1ocRsepGCPCx8R9c0z5J79OSw844krz3ZHz7F4sVBHb2K96QdmW257OB3VCz0x
sMs4d6b3FTCmtWxLxE4qbLdfKCMLybVwBUmQkMVoitScD7s8ozVso2gQbHLF0udp
LVxlQnL1s8C8q21RN/SkD+a2mjlUgjrrC0MHchoTVpbuU57EgXTYUWxLtLC8UOXY
J6G/QAX3gWmocqscDBY6etiY1TQR6KxeWmFno74yqSdI3vjTpFWGijtxcfHdKWss
mgD9Ihwy/6TyldTKTzTg4uBxwoUaOtA16rY8UQxdjTOUSiL2eBi+SfR1RLe4X1Rx
aQnwEynD+1wjJjvS/5dqlihhIawzmmTrwuXI0KBwmZyjaOSnsrm/Ca6DdIxXVtZg
JinaGO3w0E18pb2c7EYjqj00oFa6XI+22ce029K4elZp76T5KCO5xZCKhb9q8Y6A
d0mem4P0IrZwPJv9rknPY+flAW/PAiGVzxyJL3r7TuU3vSzWPZzC3MS7LGCK4Dud
YrOZhRQCQ+GJhMXJMF9w9nz5fU8U1+hylpMnzgOhTPRoaPLXpGyTiTyXz27u/qYD
Cn80JB30ohVnUJrg9RLnyuel8AGvGhi+x/t5lqEVEbpyLyvo7+mf3pQEUx71XlF1
KytD3UC/njll2a5T4Iz3Brk/98PO24KMZz1BbLBwbtOtKthM6LcYEv1Oi7OkcAbp
4UJadvNIgg5uCIqul+8E0FPMAkWGmyTE29Esm68xI0QHD7LkccTYFe0da7QjgCAn
MiZHKaOqeslW1R8dq34e2EzBWerPZ9mRChNqq4FJ9cmf9NA1VoG3D8c70EmK37+o
J5c6lTZ+gXAhLViaTD0MgzlxSQ+RSIfaqJmZQTTrgSwbiH6zUj26+17ob50wAezk
8x8utrN9fGv/x+cNSvukeoGYV1SOLWd1pMRTypZ87L/blIFwGufQSO2QPLnFzUXC
QSJDYo+Az7ZuWtSXnvkfK6eVCeS4jOtgtEukrgzn6mVlX5RSt44vaD5OyvcojsRF
kmo9tIwWzGAiAfJm4XN4ccTP7siWQBX8Q/90MzWcG46S5MxIrz5Tzh9s0xxGSWrn
uLnpQLP0N7gChVD0yKoBhX9Gx6Q1/Zrol1Mz3zmPgu4cgzotVFyjl//ihedDqIps
+7xLLgnCjZWbfGgbJB0z+ShvJBtX56W0+Kp64Sd8Di7guv8WvvknazPg2qXX28Dz
jNIWCRYnPPUfA4hJTQnsViPxw9CsnghZJflL5J7pue1gu1o8Amg6/XdpYdQf+kLN
Lh6hXtjFLLxFPJU2dPvIpX48vvP/1a+Wt3rq+vQVuYB26wH8L986NOkgtLJRcHaV
a7AYw3cZHD38kMPtOpGwUhxAbhauwx28RqqH7q79uzGGQmQebJspUwfpTgacKLsx
HqUC3iJAjxpOqckoitK3KnlnH65xk46ZQ31J6JJOOLwpv7pMWEcQXkjrRM64Si0Y
KA29tLEaTqbn87Deusd53rK0OAyHyWevoHPTejeoWWoK5RUNFKHHSV6SuWzCyMgZ
clOFNUtvzZ1RwODXwGwlPXQGU9uDlgQvXzN118I1sUiXpAlLuNK3G8BGWXGld+mp
BoSMm03FQXUHnFLIBfYwvCHAqzsCnf1CdZRNq3xBDoowDRZrIC46DoJro8WgLO2b
VSyp4odXyUEaAgcvjHR4Q+VEBN29Rwgp/xxTRjtTLmPRy2di8UulMPgnFViDucVd
YbYUmxh7Ls/+fbZIY5JJx+iby9dKCXcImcVPBJq//PocoTMKUz0kOMJaukddPtx6
Rn9agKinW+uXMj5AhJAikVwivr9W/psibqmv1NDhxv2zZkXuiiSJPe9z17Eno33E
m+jgjIx57htXKOauTYM/mr5LthFOtmtIrmWs65WnIXMw6ahmKUox3EM0SKoUsQNS
YcP0oRv8WNb7zM9dm4YGffjYwSmDB3T+2Wn8KzUJBZ5VOzMyNGJyxCkpB0V03KzO
TklgVmGdrHOx+d0bFSlpqwJfLXVc70MpQCmC4QLhtFZ1+DxsafNI2Ql8qV+fhGdf
2XhVCca+IZjWHLtvr4SWrTrALrN4+vVxBwKdkFK1sc3763EdKxLJzc1DiujSMuqz
0m/jkk2g8bZ1aJLjGym5yA4FJmsdsoR4yFOp8QLQCeOKMmizdw05sguNl5lm9CZL
5AH1Xpi22hEE8N5c1Wr9tp5EfJIgeIV+7qJ6LVgbKuNfy+4ARycmD9BwnSq/DtLf
vbU8Xqv/4gIDnDD38AMQJyj/9kEFC1mSF7r5Ivqxs1Hv14nHowp1nxrEsD7CTrpK
okQzkwQLMbFHfo8wdZ6LmVPhEmlikGc1UgxKDNuqTLaJloStwHHUCMCH8XI9fOSR
84j+Rvvpg0pTW6iNXpDC8KXCk6FDW3AHptnOpC0ANwXyT1Qschn3IYi2wPFFJW02
zpAAyEQq+v3r6Vn2Hbw3p9Jt1o37byhqGRYDnpSkFgDNZ2v+0o+Dz3a3c0Q8E645
Kzojrlg3wVjtSmQfY6bMuafOkY15vdg1vcTkj+GnSHAc0YrgNgJivENvJ27UFPYH
9p8gxgTjXEaolE3exr14IW8WKJx5XXuHHH0OO5/0fLXUH3ntmGgZBFURAYHSMdOh
d3E02TFIPS2+ENE4oxDHplmrbmNz2oSIN/ZhQ5Li18voys6d2p/qZppIEsQaZwZY
dxv7p7oYUS3lxzIvMU2BEGSdULorOkvGkZvMYZ3gBA0VhFQbUpB/cIDyRjr/gdDP
u1ixmXNypcnEN9EER7vO9dDyZR0kXaq+AOWVbrGs32WZwx9G9t8piBH4n2zOwGgH
6BdwghLEFrjPt50K1Q43Uf5VFuw7ohC/Kd5hlDC+FGlIL/H6EF7KMAdOSZLc6t6A
jqSBhjZ8/4zTtEDmD2lBXkwD3zqwoUx/+Z79+xfAE6PlKGiHh42vcY78BnRRPBO9
1vtm67E1FvY/yXBOekst/a3GsV2alyl64lZsGmsLDM0+O1iKsufsSOMReoSTvn1I
joJYDRQnnal1Oz7L+ZHlZ2e9769kCGx5czeg9f6VuSDN9sDXubz0ZDI9Y6xfMeuE
Z540KrHd5XPpRjns9qer/k7COjYRNH3SHjpgNBISsLl5nV4J6ccIMNOjOEqgL7SS
sDFHBz/RwGOSqBhdU7qU9w6XOUN3hd9OiUW4+22MA56SzC8R/B6MUOE46Vf4vvnP
S0LaHIpQLIxn9ju6cdhgb4EL1K/1uUBpsGV9mbax4VBHJGYGUSoXAl69/szXvKJE
FWUKKpsIICxqSBU3kSII1LUtgcx3TDMcgYwxHHlM2E3XYJ9OPkCgxoCc+HhHJLWy
TraLDi+NjAuPEjbddj/eMJvcnkKQcOYlK7megqN51vzN17wq6BlLGXkW99iZgydy
6tpgbxLBXK6dD5VaqBRlCQZGszgtkar9jOL0vXYpChW/c0RLx+BXmbVwWbbKvJyL
KQji+RZ4ozEiwp2ydB/qStgY1JKs/jlQuCLX0NeSo49Q5yD7LL/5AM/arbEYqUOU
FdE5MwSS5Kn7mRfnm62ikngxEO6FQHVwXXyoBkwRXMe2z4UwJXWV33NpbxUB9VRj
CRb5LIXFD15cSDgWWdE2l3fz5hcYL7VtCpeZxMVWT4y2heOFAKXmQgVUzPu0R3jK
lPqfk/icM09d48OTzFeuXSBdm7F3HxHYrSPNXcNA4H3ImKE3TMpN4xQb8bZT0GQU
/a/jMROjn/35SAuyfVggO1AlwA/+VHj5mU5l7vwtJQaYM4LeowsfeP2P0twbcGxn
Ws4ofkbhGTbtcE7XuddwZHNy0mS3+Bv0oNP2GDiVFNswNsFw2U2iuBubIcXvhwIp
vwWJO8Yo+cl7wUtaPTWteHh9ipTBzaPAQbNc4n1HWuQ/6Rm342itlrn1tpyPHrm4
iju+UVMspxFrbEalWzHtAbLKkfv76LfmUVgHfY0onDKQbQChaO0wxzXij7hCVYKI
I+m6rI25NY6jHnFmkVivHPhHCLUdjXsxbH3Z74EZB+K4x6xRRiC3Ga9eLY9Cj2Ya
c/fPCGGUNztA1KB+bAP04Fv9sN7ZzR8C77mUBaV3nfe9irUmxWCfaILjDIQ5SDEH
fRj7UsvcJVJ9jL4xeDe5haHfDrD0rpGV3M5KRvScjNPZP7UsnbXFI9AzxerphyhA
WMUi7uT5WVXS++OLo8labLSwpBEIGgoL0U3Gc/n4DPkIsk/W02eJXuMj0IZ2b48R
SA69kInSN8XRwUvpMQDe3HJfWyaeDNCPwNEotA2ctZ6Vkj6rFNv6W7eizPEIX/2z
WgogguUxz7Ebc/Q9ZFVKjEILyJpypbxsW8S3sT4UM5c2BtmAXViePsmFxcXMjhkK
K0wMhj5hnYSJn4XcYPWB50RQFc0mgmFlZ8jourC0VFs7v6lingoZ0c4E6vkh+4IR
T40a3njHRSkAYFsyb1PO6n1DRCaUeSX6khULLbcNNGgSEWlUjddR9ZdETUJJWlep
0vCnUmQtACPIHeVqP046hsQgpro4jiC+c8PDiqzNlFL4cYM/bGWH2lQ1c6stOI8d
8fUhhmaKk2IxWDJXHkknY0Crz1ywG0Rzl1JbV2gFdp8tK7Q/UCVC5Sv/OTijOqNo
ZkY5SbSt/o7xM3Hd0a+pZjNugsyBx7SGwaQ0qBOlfDI8m7jQyoL0Rgge+li/yauD
9WTK/4NLlq2duDOMamU27q+ygCKj27sMh84uBXbagQm25cED0Els9Pl67gwjbN7x
mxl251K38/3YISsX24oLpzwblogZNzs8FwYlnjxGBRqbRtN6igXe7HUGvKxhaYeZ
UMMHF8JMSDGSraKxrnHKrLlx1MZujkFjj9m2YN+JRelrqsR5Qd7qXx46W9ZItMmQ
7HQrb+9MyCv90ahLy3Cd/5QXsno5pU8E9ysifFf7HEZfh1DxZhYr0shTtwv0YQYj
Sf6vwebxD/vgcpvMdEWoLwtxpuXdOnpDju0I3XtaYbs792DTjK917C2YzMMeCYSA
1fqmI2m/uh7IUCFxurygAE9BMftmdCmr5Hgk+EDGqAPUkeeBB8BLYMzk65L5YN3h
yTGgGuNvOjtm28dGuuSYoR6DU1gum/9UVAEj25NpdlM2hBGBU6uvCwPqe6FBCy2r
qYmf7SbLeBvvjCr4zif7/iSv+PFEBb5nc/EFRNVYs02+Jh9DnoTpXXEb2NAfGZdx
4apKyrznzkhP8ZcXjQu7WNrf9TiHELQNjWFZ4nDXtGg3TzgjqXOqHhoOPhTeNyCQ
3KPLi47pou2FdS//nmXdRHPwEjeIGQn+slTI2hEEruS9fY4Y8UwJgCFJw5RLSFC8
R07v8FH56EbcG/61vZ1jp3oSSDoKK/PY0Rxud6Az+Vb/s25zPaDm4VWPhQe4LPa8
3m2yeL0ykqPRazUG5Esf8emLT9Eq+eb49Izw6Jl6/8AxZIcR9Hd88xX5OnLF4ELi
JoNXTtQBmtbPhvaPROON2WzytrKxNK03z1cW/dY1DAmPBKElfpc13e7yfKsX469M
h3cr6/v5TUakL39WTPOOLFgi+EOHT7ttWfYv9ZVBSoan9ufdMMQ73FnLTaq9g/Qg
xRX0411BAlGh+D7cBAoEWlq2QEGk33ZOxAsCxGbwy1KJtmh8F1tMeJAq5deyisV9
B/CvTxMeRkxGbJtPBcCL2CbymcqMRhm5krvcZdS9/O41l1o0dcTT2tQqDQj1szq7
7zroNKQHHAwrdeSZedF0sru++NwjlT07fWSXlc6xQzQ1e2rCZ4I4Ah+M7V3oj4hY
j9YxwxBUosZr3cBl4MewA5MzhIhEoVaPnVS02wBubpNSyIsi+bheW3lJPQ9Me8OQ
ZOgqVmRDo7ue5ZODcGIVIKx2eTbaoXatgTuSzg2Onji7mNkfO8Exc9BMlIaFZrHY
+biUz6VpvrCX4091uZCRmCVjZZeYQwAasxRvkBv8q312ZTAd6BvspGtc11UDCzKw
X/+CayANVTv1XjvNst5Lr4sjOGgfjlxsWgTaJp8D1j+vTqyDDBmnMZXs8EBBAPfX
mnwS/CcKFTcUXpXVPVtkVSAZvzlCpl5sg9UC5GOaQheIrHOhr6PTOhHLIizPJhzb
28oEu/v5D0b8CikhTHLWQyLiWioJ3aH+oycWcbELgq7yWORPb+xL11ltYTC1meyM
iuDZuwZGpZjxRIpVuQwPHXYjYz1TnfQXdCOUyNVtvWBXa22sKh3WxNy2K8z2Ch/x
Cmx4Atdh7liVXMS2Trtc1EbjnpUupxL7pRnfiulZNdembZkhSNCWcKSeP/ZOzbsr
ZexYnDQOF7ikvMfS0rblAoVst6l02iW7LsHRnz6UZCOIKrmKb0P39zrg1IK+DiiD
mgw1acf39p8Beqw9VgeBW/0ZGA9IVLVYEhXs+hyjytDNi3L1RfQUtKzkXlgV3BTV
Pi4sKhMGtB4VGsspUSPNJEo6HWXvGIQ59rBgvowNyWu6Mk3i9lTesYIRDKr9YL+G
05ERPWrsEgrOIbepK/yYf+L3j0PUTp1xNY2mpuOu3tA2qXbS4luS+VS5OkBWcDEB
PPLgi2h15oQ2zJDN5KqPTjmvfbL8UyL47fGy+OTJroeBtFoWU21VUz5V8V8gELWa
MDgkiXPRsJBUXUf2YYMZo7c6GpH2swH0t786mNc6QUTb4i90Ryvm39HFxHTBl1SZ
GJIiTxkVpO7O3j3vtcaPz1fwYr+OGzdhop3NTgLlxlPN60gGk6XwslR5UmBTTE/R
3Yq7xPgmjUVPgBstQcr6gwWU23QKEuKZJqgVETi9qBJMAMx9SNwlsK/1rjFuweXf
8OG/I+bXy63oetKAdkgUYM+VxFzyiF+aFLBxhNoijFbz5LWbV1u83cYGxauAV2ql
2fHrWPA4V7oSK5WJfDo9owY2lK9Q7gFGKUw5pbr37p8gcf4gst4KOrjzAeLA2Nbd
f8z54XyrBq+kJNLw8Iv4Wbs4i1F5F9bGy2f4/1IXpWjvJz+gXYQm5y1M2q3Qtcci
oF9HldJifTxUQrDosg7OAx2v0P999QiUIA/3Bf/rzjeSHBZzK6baVnnxoTr5/vso
1FxOL6OA5jjo7OSTfu866JZ2yNh8kNWNKC2onFYV3rQsWwttm0kZH/xSkGhaV6c1
pRWtdzd1CfdveUazJjdTLZmATLN67Gtd41PKBvUgdLloFyp7P5T5pdckJD/kK7ol
0iBWemK/ogVA7lOR2qXjpsc0/MJq1q9zmgbQRlwruSqhUE0jQQCY34NUmV+q48bF
XT0l/26qmpX58ryox9l1iiMTrQqBnJTshQdGiqIAmItiaOZI1s0NWczfKzeJ02fI
vRrc4wfmknWuKWXdv9er/KAvZ8u8WwghZgE4UqEM65Q7SmoLFbfDwvhaEvvAJwuA
nX/B2LSepIZRlUb5wwhTWBacKsftDwXNqt8V6JWKz5NJzu0d3xKm4yBHMkAsjDbE
CGyjxdlQ9ohXY5ZgupoYIG6vh5BRcvXRWA8IvoIsHzwb1Rl/5qaY4oUN6v66v3rW
Lt+pe2CHv93IUwxU1pJTfy5FJ/LNY/xPmG/wn52hhLv4f4YKVmxVF/duVIwL6jmz
DmVqoGftdPZ0ZV8qnaWqLg9OBiA2wa+LqKhJu0xRZco5/UeWwmvnTO5DMTZDGgzO
BOawygM5lKnAMk/VpCf+5lKX4OWGn6Qc7bI7IXuacvwJavLfTPL/xDPxTtZCUiaV
85koiH+N98PkTh5TR72JhyTZnv0m6lKe0f+cwn0uoPaioAq2d6mn5Inbol5HkDMq
dKcx1022+7zxgTpUE/6u1R2MWfsJMJnYjmQjNstJ0rnh9v8lqMy0h9vk5AynTqsh
h4RVq0oEJ3vkrvUwESOzmZg8990inja5ZeDlPhasscxftraobEd2XHMAOA1v+LFX
Udpzesw2PKXB5HpmBjqgl1wJTYdOqAxzhbdkX4b2ZCRmn0Sah4pJK0WlBcT99E63
Slbo+IOr+rea0opKE/rMLjOJuliiqhacp47rU2h6Py+1n/7xlW7PCX1SPbb5iqCn
pyC4carKyx9LNvFzYwH/djsNZV2ZuGYEA9NdzzxV8Kqr73RkmlLD2ArvA0m7IOb0
Djfas7p60Wm3/rgallrTwhe8c0D2yhreo2FW3urzhrGtZ9MqS2UKW6clsFFUz7yS
4ruJPgGdSXo54/Vn6dIGT11XfnSgAjhtWxeekcrFJHw1S1jjUFVkufQUsFoKIo62
rsO3uoMHUHa/SonxhoChx1kaiEHek5yO6+YbSzHM2emujIWnRhdKllbu9Wyalcve
jToh5gENDvdgIarXn0nWaqXKBCjWoc4jDqVaKTzjYyk2MeTzrAnlNM50DsIy1PYB
Msuq4c2Bg/G2R7wzy4WOGn5/9MCcSme9fqhEqr+eAKWkbyyvj9YhxBgOu9uPpcrH
EqBavt4EKRO3cySY98mG1Ooyi7UoRInIt9ZmuYedBu/J76yuW5XCDZqLfByf7eam
6uYdwlVSCv4UGnF+XPwqr4zNzRDoTP7gkLegl91JIuMXpBowF8ZTKZs26uGj8UFa
1/qoq5mMU0EBx/UoSft6GvA9PLJDtWDF1uVYfVPsq3rI23gmEMhw5QPY2XP+0Ifi
jH4kQnf4nPzveiwwpO0J3ZXD/BdrxFAa3rnHYuRioCncLfbt5etxAAoLWwjPsaL6
JzMs8ilNKyEhKznYyhmV3CzBm3T6kIBdZkTjO218h2x3OEFRfei3SqeDOB2iAFYR
s65Z8Dx0AEwGVH9n8cKjIt2QTrW9Zek7iAwEvLplPsBOkvT10Rr5i23LxhHOnYct
sha8FDur6/RjvuuuEiM/fcog3IG2dc51848+OV2NXbtdxtixtRQhl2zWEwXPdWtT
XvqZuNpesqkXdV6ybPSMLOyf4gAfEqcEguyvrGsJtcN9YHvOGCFd2YvicqadLz9K
ksUdd5JJYBaZdSndxHj5NflwUUfHfUe7HH0VVr2RiCJ+E39xybiHOxgA5MfkwEfT
mlFfEqWXBEktoyrWDzGpEX5EhrcpGL5GO2AzwebACUzXGj7MP9m2lJ9OW3RWYDYV
95urHPI/CgdcuDAVBvDvQhwPVVmwQSm3iTUw5PvDwREf+Op50tsnDOdMnnxg6RJB
/ZOcwE0YAH6MayNjTRsJuANeMD/XloIk3vIE+FBDaB7muINKGmElqv8pyWRtAhgj
iHVBmFc82uQ+B5S5F8CTKATA4JGaVQA78lVjwyuYYv6u6BHztb9KaV75D1wGrg0J
Fwcd1Kr6adQjI4T6ZL9Qr5Euq8YptP+Y6dvuKnj+LJqJqgtoyspkWEONuGyWXAFE
5KGZ+AX2H+WQrp/67rzZtYBzVRJ+fZWOxgiZoO58VaPCNddd4YyejgkdCgNgWLWY
KY6SlGnN41+T7mvhUPgrxaelgGvnBqUz13JaqV6ms00hOXzfot98HMGylSIGSRiH
3fEERM/LUUVlr++9rNQkcBRdAcjdPYJy//BwukEsoctzLLnWb5VUpWJ7dSp+/qV2
0Du4YMqleptCiV1p7FIgTOs5V3URLSlkexhlnnk95HibOEh1UlkOX+0BVrxlZwBL
POoWI71V6HXidoFrfisMp6UphpPVceuyzuwnkcS68y80YOMltX/If/ZWumVwSG5L
r3kOH97HX1PvBahzTgak3uFTAglnJqvDQye00xlctrHAiAkioL+iB9yZL7ZaRyL0
GHMbhIfLEDwYWJ1fGbimekZtLwS1IdMd8vgxTf9zj0Bnbwur7Ly/C1tGafYgM1O2
uuDPlLaAXcmoPj4th8exS+BM9MG/rYISqGK7KNSaneigjRct8PrOM32EjJwIBP/M
eCbSwVvrg+wcy3YekXe4+29SXImDyQEcMKuHcdoLSrqbhnfepZQEPUaQs/qyv72N
dNIpexxpTKwZf9LDgWKIuOtAUzilABx3dcaVZ1tHdzmLnTIb8/gju2PtJBdr1uGW
76pvQp28aRQvYPhP/hiNYRhLzxXwZX5nbpd2yuGABtQL+S1XI1KIHxYO0YaxuQhj
bvkHFeFa4B8rim5E44/o1zlyA9ztLjcUg0CMFjZsfSY09f13ziuGRtWLkhwTIRBN
Av+W72gL6EbvPT+DQFVQt+8+Ovxvo7MFY+bKo5NFqtpyUb3Qi5rmNC60Blu360r6
OYjCLM/S1JjOiy6kpT3dhdE1vx4ZjTXWukBisgsVZ3oooFGB+8OAc7B5s0sU+bkn
zNJtZOb6cL+cEGZKplgxeFMmzuf8z8S+JjG+AG2TG73O2AYdx18i2NLxBsKzH7br
UfH9yWBR0bShuHzQp7NoaBtw1hgsrm6ZZDcQ2zCXvisbpaW9jKBkhd+aKRAC1hHt
C9H+G+yMkyQJBtf1ko92eJIGEF35YiSAexFH4xElbnKJmqW5jjTX+X8M1JRCM+M8
rLrv1zaziLsPdxtd7J+yXxHt3vum8FVTttU4w+cVXFdISS8J84jZtpXVCV9z81VY
1fu8yNI3IpYtw8X/HBNNI50sYmdTJbO1pHfS51uUqq6WVSV/CgKS0Aaagih7wvVc
CAuMhwLJ7gtLrWePLdDylp+4DW3yQ662ZtpC14mnVfHT0NsIOUPWQhuYuOZV+T2m
v+juoyO0mXkk+IFTtXi2KRIcbswBBpE4msHOSHb6pGCb6OFX0QTaXCtxoUrXDpTd
BakCm3m2gTk+b6vZSLvjjRKN7gNY6gkYOJoFx5pcA0gVYvJ3tB7OOujYZNjxU4eg
mfR/kj/qrY36QwHfLFwVqFJVLflA5R1eZPoFfC0xg+jFBxWXk1hYOpQ40zgPO80A
SQX4C2YK78xbsxHyikj7eiT35sQQtVuyAtFDXGO4U7tSS08lj+2hEeMRtgJnThSt
S5pZdKxf9m7lNaCDdCNUhLT6HYOqDhvOMtSurMXbApGcIkl0A87/C/Qio42O3Jfb
JoQzMihDJ1pFxFzX57mYGZS99w1N8A7Rou3c96rLsp2zpPqMRs7UZDC5fvd5C0Vc
kC3MUf4IVlDVu6wjuus5BKF5jPZ9nYDxfvfirxfPL1hDM6QoI/6IQ5XxyWy+uJfR
/aZ3XBosprRsoSQM1HPno2CuqDRtZOA9Tu6EYTNfrpD8HcAl3DgeR8D5C485UEy/
rLoRuQByE5KLdd/Vaea1BIaff6pDu08IYGI7PXjCCuc0+PNO3nrT4Hzitar6qkGC
YaCnNBmeVVIgn83q8twics/ub6qACSOUJm2PVoo1FeGeLbIH7SvmfaZYbCOxK0/T
eXYzdeD2CalgSrmpViSa9Ky/8667CZlDvcfKFlHHmhZeaqg5hlU+ER2KXwvSCTZm
7nwz/xJVNfk7EoMy7qVnAgwYIlu74FX7p5zfx4wBfzyCXd4Hx0BcPFAuK87iVQ21
zcILG1qhPAFForFxqXOxWQrbHRooANgKRdmhiF+WoR/cUCFMhFitxlU5oVDUz8pd
HlhXSUOas8vatoGL+xMAossCFfd96v3gEXB6Mgaw2Ak9MHz3LAJfhOzJZnfZ4G9H
BRZPRAmkeAabLldZWx/vG6if9ud0GwOL0Ij7WzY5dgdUAhrwVmvwIN5qF3kMhH3w
tkqJRZBdhZ/aHJFC9grcdeFUszaovt7z1RhINXLU9TATBA9MOVvP4OvdV52qkVQ0
0JQvh1Kif0p7vEVvvscRnWwsWhvi8JcLszDaIyR/YbLmiJzINQMvF9knR1XoexsQ
kUA2R28XXreqXeD2qYd9Vt8I5ilEo8RpuYI7NHDJdwPclX0YetFsG9e+uN19BOl9
SNbhBOnVg3puMBKMbJ5Ye2ZAcgE9JU2fRK3ju7cAYjWifGz7UJxcAP1IYrZBMQEk
8ljJMm+lLbhG9b89t/v6KG67D+C0BHBBTKGw1LV6mZVgqHMKn66TH/siXnzP6osj
AQAbdCdw0uh2w1+2oTACCcMR005btACeR1R5jNpWJ3/U+WqWzPyjA1xxC3wuW7pj
VdylRrPbJXUfZ/khAoC1IKNxj2hg9AWGof/1KoNeJwALaSubVUrpGfdTEPZfXIGA
jNRYcsB2BSH0wtU/A4s7hjHL2XGV9AVOESWcA25r8qty6+0E8z9W4WFHb8jrWXuY
zAdiV5Ulx22JuH9BY+uNAx25DHEIi+jrElGszafvoHga9TuURcrC+Ct9kjA11Z5C
KnCt6DeYeMBI0wjKIhFd2EUvRybpCNPDaA3XSENia/FUiTE9sZ/K32AnJ1djaiA7
3+8MmAUni1cc1wINVyam14YrKPaH0d8YnfM88ZgA8v/f29MeFRlD6Bsh0TFO+AZc
7HI17uzrVU6z14+AxK7+cjDT0aXLj1zEsaf+sDGtCT5LbRNUxRO9uk7wbbwHlJPv
R2iIsT/YwiD0/7AoE+uinHlR5BN0koaXiVsanrx+bHWuh9y7rL++sc2/4xEAupjk
n4ybrEwnsS4/QpGKlu8RahTdAxv8onxlJMEi+LOQkDe6knUcZMpHNnLQgAusaooW
Mi5A6Scuur+xZDO+f3KXwju2dTKZPLtOxrGxlwVSipQ0VUhZmgenv3kFs/G9wkHt
Fe1IFe6AvHppgC85ox6dLXph3p53sv3D8on7HAjEv0HX9cxwbQR9xVCqoWLfo/kE
7B8ffNBeE8MZ1eXo7QRHkCW5N9Zb8rwU99i64/HrvtC9wBMk+BWJ4a3cLOdqedpv
1R/Gjz1DRj70LbyEeL5Yf+vlAuDZp5OZhQphacSGqzyPZsKsxjDU1+eZDYv9qvBd
ktWhHiWBYGjtPlrzlSBZQnC2m177EoAL+G3yjfI9PP0e+7cnQyznxIPGBDayaYC8
Uco9sy+7Lp+mQFJxd9x3o9VHJuMLAtGphhuf3KLNTLI0L7BVBnK7ky+8659phnLw
pDoKFtieC6BS2sohg9V4zSttwTOuvseH8nvfIMCQTrzfXVvqkJftqYrWLkYdbwpX
db5554vq8TrXTRza+KGwbILs1QVEkW6cl9I2htqHnPbKK/QPZztHW8YGfFba1Ixp
w4Z0SzPnhwQg3kmlR7WJdUSKcpYCymdaT2ra2y4jucr7jVaHnhqyX7rL/WV/6ZTQ
dc4vmUvxWXCmM9Sc0J3LyRoQdDcEiWQy3E5o/6yfBNQkkS1SO2sgNhoKsVfDu8Ul
YrPR2VG/qeLVWUDjBxn3fuCHtfSbq+8J9muInyk/g4aBGC5732wsr/6e8C/su592
U5GAu/dEdhxsDdEWYgenX3ik1eTxGk0BEik+ja5WXooYA6S6eJttW6MHu1SWX546
Y9tJJzIOYWYWVmA6HKlXIRCaw+UyKQY6rfvhNLBcWhsP/80f4bbQZ5BgBRntXzXg
GacMAV1biny/wquMv5VrGzFy7abqSvOS77t+C+Vr+VfVMHgn3CCSX9OpG687rIHZ
Xt4DDatptyzpfcqdH3qnKtvfdpTEqrPJeAcmpFecdqbswZTF7oOWSuwFtak3PIBm
mkoG9t4y0L2DZifCL4AQ2uJIvaZB5Znot+0P2n3xnglDbHkg12oALcITzz4Mhb0j
W/rhRZqhG81k0CoP9RrxaQoHJ3nQODXfykL0K5Y7RpNR0DWmbYa8H53i0CvS0vIA
Ni0ywobik1bGkLo9TP76BIIocwQ4+lhbxz+vR1QiF/GuaOcy4wDe4ggkS/KENEFp
0pWoAEHPBgvXcj4aaaCVNQdAI2d/AqXRLvnZwyP3qZ4ctiXSFhl9VKPZMeQIxObK
xtCJo6DU1U4XlKGfyc0RTYH+Nmbh1+IYZVIjdOsM3JZglVv8GTqJFl20ZZaJeYSR
Tlgw/GF0ixEbBzoorBe8npnHMAyCwcG1ov1YDCyHeOoQoYczdgG4BP1k7ijMQaBd
XiaHTDFeyZIScFNL2O5RJ7sXRas+NUiE9jAnCsImObOhkxC6UU1a4qcZsq3+UJ7z
kTpbHTkMYMSVTPRmL/ETCFcURo4d+NZKYvwa5IJ5G+0uFVaEYnVCdAZmk/iI418T
z1hBRGtKZqyLfUqH+lzjbOWZJX4jLIm+FPC6gfyvgMJLTL7IbTh3s/K9VxMVwfQt
oRqWD7qA8+ujrKwHtAj+jWhS+QdrMnl4x++Cd/gbRhsFBHJufYdqcpKVSOu9LFvV
CXTvy58xZ+jFpL45UfIMWVGKZUxI2yS662u1zBVUuJHlGC2NglT2qZigic6u1YUB
I51XQpE6/W7gNZbd3xJpaljO6lG45jTGCuLJzcYI2uUAk0mZF5eLglsYW2ZBFCRn
JpLY1yODWsZcwGNmK1W5hcLjLWAI+hAOOolHT9KQV5TO193LEazQTfZIHKHNDUvx
wtIrMbE4uwxr4VvBfAOlzNg6wXgLS8JFzYCy4qsaw7JRvp0tKX1Nq1Ibhppq+GBd
Ezfml4zfIOmL0DsbzH+fadFykmoUpXBk41JNqs2GEiVbIWyEwyYAkgnGX+q+xYa/
Mg44/mcEqA1FRcM5Hsb0W9IUPYh/wfg26vqWNPathf+aTovbawOR5RkVjHvJaFDW
45J/wdIMfANHXRLgtOoplEq+zhx7ae//X8kADWHlAy9EGdSSX0Xf09K9/WrRW4/4
mYN0MY1PjwBs501Qk1vXDY3Sfqi828ZtO6ZhyEjAheHsaYokZS4wVtiq8c7u3YTb
bzfjFZVSKXJ/JOW+X+K7zKHGRtn8cm8cKtRRW02IewE/eIfvduNHEDOFpQzj4VqP
qaf9YZtvfLvJGerVZ231dflbL+HKfhnIIswQTOt3GaSMeN7CKZpOpsZvhc/45JVa
xbLwJAintBpeINsQ82nj858VCZSrY0LR5tu1fkeGtsObmdVKhzU6AJ0APcZTmkmV
uaFpYfiD8II395NF/5A7FJexfGx12EwilHFt/ZPP03d7/uKwnoZSJzjZ4It6zIV/
lUocfNFrhEpt6erNEEqVEJLzfpIFviA8TcGMp+wfbAYo8Ily/BjX4nMrsnQlmjup
9vWy2aPIXiTxtKll3sCp5gCFotEiZq/sI6beeEXQ1elMON0aB9wasnEvPyxKh5jj
TjGUZIP6s/SlC+aP02yGVtkTM8FiwxBNNp87FrB76LvM5h0/ybKWeCypqKm+cQAj
uxfrnuOw9ELOjEp0xPlYWPKfMxAeund/ziAMMltHpdXhRsf3n93SUnleO71NXkVi
CkGShbNYh/pKodFf8R0XNkZY8efTknjG0RSOSz3/1ya3X7jPORFLQSHlg/NqA4VO
DBcX3wuwPxi/rTQKJ1/On2SxL7NChDBGRxzFujxHoQruPzHTuTWCyNpxo6VSjlPp
geFMSK6Bd+suvxw0jpyPYo9lellGdJHdcr64RnLX4+vAN+ToB8O3XSFQ+VpZFOK5
BV8T6xUxbv0gebbqXTSsqfbHF4or3IvGg8PwZhl1hoKYAW5290uFKRQO1DwQzO2P
hxQRM74NWDabC/w0IrAxK9F7I+WPz0ovRKht0ejxVZAthHU56FzrG6jwnPQDgHoj
euyQKQlFENi/sMQsPlbaUAXahJL1UZURrDYFVRCT1sIkwm3Trv/EBW6aV+ZLO7nU
DmREfMnz8CQP6jdWqRje1i+o/GdI4XKAnTUoyqwU2CmvMD0PXctDgdlIUXjveoIl
9KXILUZXBSH7DI25Ctum9sQyWuKDFB2c1D2MiqUmYLDMijEkit9yavqpKRffkzOb
DT1vxcQfi7/lAbQt0F1jugkQlvg01Z3oRR5ceY3kSQf4ZimJAJgaJ6wbV6rp3wrM
Qpnbnk5d7HQWN4P6M7CtZvQ4jwHdz734/GwNmcQyBPA511WwsibfJlNDOaEK6YDP
ikS2WyjMNKiIEXlPR0OuE1OnQrZaPfhVjzTRaIdYqa9x1RTGYaqrAregIRH7VhNr
31VH4iggWfU2jT/tVivW6HW6CER9UM8ptba6WRDjibrdsM4b7hnl2sT7hUOmDdwU
josZ2rIY4kVn9TRm9omuTK1cdlNyctrTgMvFdaGXXLZMLi/HTZUFHqOGrfcEgxM0
QulUc0LBf17QL1+e+DW3OJ7Hf2LeWbNmM+MNuTEs7vGNiimRsvNcAla/IEauSqx9
Xow1HJp9waoBeWt7PZCgNeiTaQ7D90NIGRxHH6/Nx16kJ4tPAV8A7lCX6L4wCx+X
owb/Df79/yp+HdPOFEZr5FeF+G6BRdsvzCjJmmR05LNjOmAjlVzcQ0FibaWHVNuT
JnwrbMej0b69VmgUtgDfBE9xooIgz/MHE3xad4AZQyz8ifksSV2Eo882WhVyW4C6
aqpK/xGgJuXTy+VtQPArgCuSs6YsC0W2U34hFEkrxGg5cAuVI8gJP4hPLmwE+kKR
gmrsuAACbicMi4ezL2NT/hKhcx/xmR+1BiHayUd4vM5tyCAujOLs2xEDorPhxyHm
2t8uJfONrSOWffrpl7XpkevZ7SER4QZ5wVLQyaP9voBoKk+Ze710PsAGEutAgYWz
IPFOBNDCUQCOpYLYIk413ZapEvHPhZqXKScYICK/QqCE8eNqFhU7q8bzbtcTMkNN
0T0CCFgMFYc13Npaj/+0JLwwD6R8S+pWTaI7BJHRtvXjwAfwMhYCwXmd0tZ+iLGU
BSZkgu1URJwrGIDNk2jbHINt4bG8SezRSMTWkspbQvFp3gQK8u2rUxFCbuMq9z60
wwfuQH5C3PCz+XX6zMH2bZH2O79ijVLGkNdZkG2KpMT/JlkVi0Noo8A5Vl2bM8V3
zJpmbvYfB4BBzi+/8xdgoG4i680lxP8ToewOTfcvRok1zsEJj8eHZ1X36HguqTLg
28FVUSPR2+KWrySp4CBgr45oT4X6ilkAKOsUP+S5AonVCRLzqyhlOamFrSlmPIiJ
l9+//Q6qQLkQiupQdozJQcp2UCYQhQYUitGusQ3ZzuMNwR/PtQ/95ffEfQIULCfs
0AE2uZ3m1kfG6GW+OPL06dAmJPvfpsDwqhiLQeApcNprZgzwZwnSEku4eDPiOAay
di1AzSOpymai5ejjKM4VF9Cv80wLhGKHUQkXJTz/OvELNsIF7ajTXv4jWzF9mrdQ
1qi90bw8omQgXtY2Ra3expL/Lis/tNC/9qsqI+5CsTlo17pa3orNGOnelq+tlQ1Y
0buzDoI0wUPMGD7Q21y7R8dT/CHcUV1XqIOZLClP70E8uu2G0gyMH07ERzkH4ZmQ
Td0MX4XjTsFwyopzEL23oOkLz9Zfquh3GaKfa6BD3tdedI7COttnswmK6ICrv0j/
vB4oQIdRUhf3bQl6JGSGEnRneQV2I+ss7qgMYbuXpgQmSM7vdFB3ot+8MinMpJsf
xV3G8LyGQ6c199a6j0EmaPLd75pgnGjXFx6sh+XIbeGqdPIl1Hfm/kkf0tyXzofZ
31mJWwbglK1Tm8SOsYQTBIF21bRCmjG/ltFcG2g7bAqki6bCPlmhfR8Ex6Xg/aV8
xdf1NM6PbUIGuXbRz0FY83yf9y7xWqpu5wCyM3Xxm8DiyiqSDs2/YckCsuP07oqt
94gmTo193i54x/BlFdrM2QFUrFYeO+0fiuQECAoMOY8DxXWbnoaC7LKLMf21GA1W
AQKoBX7q67Q/yHLEgk1shLuDwmygcg1jSidvGLqOyhZ7uM06+w88zqjfmj0P12uv
0/I6Htf4i+dqJQhWPcg1UoilwWmTLQuAblbs1DgvQGo+uSqUhPdXl9ByoLR/TjRx
5HkxfU/Df8WXX/3erG+UDFa/ePFmbqUQTqLcr/Um4n7a8YzwFYWVjs7wWsq19jvp
8rs9U5iMmOgHmVjKJi+ecu0lP6ASmvQmoaxzQkWFnVEk9lFTPz2Ar1IwOilptLM8
usgNLUJK78/aIYqVxvf93D1UrG+m6WbUSAQzWa0c0gJrRv4JbqfzrXhgsZ7EBUc8
1sh9hVLaFNKlhhxdyyKSFCj/+hB1RI6nO4TfkXDGnF0xYnSEJyZ7sLHIwSIooyWz
CtXXpuYU2YHs4pts11DWlDBcJGCP5xB6w3T5LLflBNPD7l5VPEv4u1CFR3hKCo4r
zNx4hEKd2nbb4UKesM/9SK2q8kFBQq6aF3K3jv0lAGrM/d+4UTzARxhJBrzDLLRP
q7n8OAvJ9J87R5jrJyHQntHsCZXxZsMHwxlWZSJlO7N8Qr3kbk2b32mgVJQbYlW2
ebnUuytWKwnSH4E3PIpQJWPf8JSibE09nHBoR5yRU1F9abrprxhIl0/H/zfFnjwI
ySOxVQeFPoN8k0fhEdUm0x1E6gconfxvIDrZKSfUD2CPTpw51/es72O8oJ1e/Rsa
SXmEUDxCVgcE9NScNB0bTrYfmCPuNw9aDU6OUWMj+TiXpnguLyZdr7p/jGnyv2dd
ORU3OvrHlgJ3V+b0ybkhFebR7aDkoDFnu9D1tyNIvVuSiwQu1nRPTOrwT1ObhDLq
IAu4ncUbVkw/t3LCnMq8kl8u21+GCITXtJXd4BjmHvnPRtONkBxopgHFFNFGpY0w
Qnqxm0GO6x7GpAlaCLRV4U01QbPY9aBOGDdI8yFxu9+WgVxzJbTtfsWguwStQwjf
clCLGwwwhTxTZ3A8tecTZ1xgR+pxwPoiFBUwtcjkCT4HGisKd9Jhnf/7wUR9jwJ6
7YbvIGiB32Sjn9OA1Lh/uDndE4BjjLOyLOuXMugy4U/sptgYRMmR/qzb/8/OrbJq
mAZ/EiaemuktQtIGOQlKvkBCEvZUWikxVFLI4KrzWQj3S/8YU1HHikPBJjh4p0BR
7pQZ9X849Wet3P9B5nlDFuIrBVharLaE3dWK2ssviC9J+KZ1lUw2CzmI08q9iAVg
aWjE5j0jo3Sb1PyuODeWkM4tjVsA4+5nwZTX9C5TuDCziE4dN9GNceTIAELKS/66
nz3A+UIbfkbgt1UfI0KXlTsWVgY0jP9Sh4TWln255amewoN+srqOw84Awjz4EDFG
yhWIMwrC1NLnTpzFhMd6Zz8UYsQTannZJiUU8ozWfMB/mvlXHf/I1DBvCCINjyBS
lfrz0VG2WHmXm+prcLi92RYlA9wIB/ZLUYAQIJstYEVK/z5YDWP0zgBc60zrFRoE
pL+M19wpZLCxN+A4m4e24pt7JlCbH87a6ZaKGb/o55Crl8tGtgTd5YxTKZXVoYMU
Xbr+8XTSXLhz2DA3D4fRq0M0yXAIzg0Jyo/kpVpEe0xPXpZiqmfU/sRpKlPu0caM
wtfWaxrEcD5ls2ahyEE7j+1TkYHul1sUqzHXqrEs5E8bXBnWLsnn4uXfOLGdSkRc
/b2fDdTJ2GWNQGHXtjWtI0+6sHSGTRPt6vaQcokyq2dsvs+QujxNcmzeUGavpw8p
Rr9fIhB7UuucVidDKh/CxCpIo5ZVCFRR+IiaZCcGdYiEpKdFg0HP5RQQmK7jpN/b
r8agEbwOnegUNVkPSaiVwKTgjeIGcWGHTxw12GimUDRTj2Adih7Dd1H3qu0jVn9S
iwOIzfqc931cgMShgGg+b9gdNitO3GRk9fZ32MIjY14ZLfiL1uor1FgVQXw27Qrm
p2EFedQgA2pB7X81PkxTKW0hjuiV67xdrrVo7ADgXb7f++70rmbILVlf3KGQTZTl
Rb66YsSDv1qf5Uq0ax7yo0EAtqSWW7i2S7JNwJ1utcbfnMmS7UqcUcURnudWCMlV
LDx/wAVZj6LK5zVV+W1pbOCq2ItSa60kNf+/q15wf/iy2GIjTdU3/SRnBsJwdlep
ulCuvE0epo5TAiip11pfD+Zn7q5R7chdRqxqo6tqnWlYBS8YSMSe9seJhwF6hreL
fmWv8AdpAcXPdyZeFo6ZZiFVXeXtunMeh7EMCD5eV4Tqa4Kt0IrcqjgMTyIlQLR0
dHf61HIzhDuSV5bqb/MS3N1KHNaO5hI6FGMMZMEhTl4JIjSrItVzTssbWmzkChwH
X2KpotVk+IgjWy0oQnVinH4iBaFoI8DTpuXSpcAysV9Aj9SNKJzIzDpKmvyAen+i
InQTC7V3L9NIBrPqyfWBKmXq8gLsWFQrD3ma/wLd7euaLIWGASHyT8uV29j5h1Bf
HjTnkIg1uHkjUI8vXfDI2a1ksoRLvV9whdKUhPFJa3CjQV1y8ytCtu2gD08hyHpM
uyAoNbR0Esxc6H4wvQ3qFMUBxamWhrOVgNuS+x63NNzn5sErWN3JveKKwEkM3sYX
e7Th8C4JRk9FOJ1INzAHqSeVMW6OuiM2M3w1MwbqJ/5ZMvd+g8bYHJL8dlKYhFoE
SJCkj1Jua8n70HrsDE216oBMW/2ly2EiXuc1FyOONo6R8ih60KXOycDmqgPdBf+G
AzhlHfmNUrTZO+6zkNXAONhPYcCCtjmyVJIsmVNJrjOm9cJ59wNxVimg3r8+zYZA
PEtRZl9OvwSmkupTlJgrk5WivZeysAeiGeT/jxkx8bwpJqnxvujZP+sn39oC9z5m
CPj/32yXWcD+HQa38fkOdygNFEFTNnQY3AJhzeP4GVL4wDXsRjNuyPEwuiXzGMr5
vA6AdBeQGQSwtNCgJTHSRkbvk1XCtXKIQGPhXvbdH6+aHqC9v+BHyNl/91fSE0Zl
EioIPlvVSQm6Cw2R9ASq7C9yZF0a3830Hbk8sqP9PF2PwTQ3f8ypREB39DMGz3dO
zda7kZJAyd6RUi3f1iq3j75+ByfPOxNuf4f6jWKbUw2nAxueaUMt32YHsllJJDLy
ezjgKZ4YPbBJEf2BGJVaZbRgQiGyTD5Y/SlJe6Rip2euRmg7j1q4sWrU9t3QE+KU
Q5E+AHtf2AotoMyuV2iWLrxg0/mW+7dUkLcDLDzVt7CMRKYmvxWe95X5EW6OF0hn
hyAdOlOx40f3cht0xSWJLDseOolcbUqKhCx0Bi3kMMdddH9rIszm8JPe5XyXnCVz
GqRypTIiEnZsEcV1igDPmnIyJClGrWMrxlTfNplxcQoNQb4zp/Y4E6fojy5Syel+
VLYpkkMB4gYKl7Dqi0DjwCnIHUkXYGhN9UBnJ0kEs9OJ8xMIhqHAIsK+bnMFi4w9
gl3U7/KyRDNX7LpL42sGeVPubQTdA6FoUGxKMkN8XWJnW9kHZrlxqReY4Uica4yf
BSYX/zX7j6J5T03/A7eF32Z35JV0gSslCx/0gzgWKJ/dn++CBcv8uneb0Uygk1EC
U0mplU/RKecDP1c/YBD6ofyERlTD/JgdbVI2D+IvSeF+YGjLmpVbYpXQ4Dq3otMD
EuvCILNIHk7cLj4ex0Xy/SaC6rFLsg89cjC5P/xAQECPVYD2MpLE1gT1vzjpbW8/
iBRhciiPpRCfPJXjQwqlKpnYbdj78B+FlkDJTSinwyz/txxTLS5Y9ueRcPt59Hk1
RTcXNBGVEcATB0Esk9IEoagPe5DrdHrhAGiTI/H7ITGWPfT4HE/FfK8kH8vfZZVx
mbu246wkn2ldGUXn14K9Mlp3etv6IA9j0bjHJE69qwCgQK5DyMXRIZjzQkvfZbp5
38Ce9SEUGXDfKdVBzjTbV3G4IfneRhFj4A4B2YY3rhKTVU8Lp4PD0WJb9uquhyOs
Kb+eZOZNJAGgMVAa16pMGplMlSxMBgx+R8JPkZ/GX+z1EytxOnyG8hcF3rcsRQc5
WGSaeK/muZU2ZMGg4XlNzHD8gCikFEAmN4y+79sGfHQAh/5t8gzsN2nujWExj3Oa
k0V8zFiwuaS59K9onnQWIvsXQAtrQumdhF2vkrNybotergS3YhmUKWKmjn0SK8H+
M2+oTBKtpRybmhZDU9lfq5Xib5bwG0HBhWULe9+Kyu/ngZPjwVXV2gR88JsAOIr1
DQIvsaGgsQnxuG99nh/bspWv5bWK6vI6cT0h+Qi+arozglraJruA6SoY5tSOusSN
ZxjjXMNvMZhlgHHeUHZjXoMjXSVAKkaUGbTx/pF9y71SVcg4ViId0QN+HluZHdbf
l7U07XXc0NnFWH3C56al5doWLUsofN6NqFBxoUs5BKD3k24paCpczZ2luC+x7cDd
kknhTpONpatqB1WKBJ/6O69nA3UqU9XZf1noGQFz1Fy/mQk7ETvalm2NYpVVXuXS
5EdVh1D7ParChZcxvBDtYaC+a4iyzND+iCdIdJiAap/NT+c7o3xo3M5pOQrWPEQA
8ovP4MuCGwJrScO5t0YOJ9vLCaMKHFLwX0n2Znm/Nf5p/pM2/ADzudgaUCoO55VH
2iGyvkGDJ2ZTJDtlQKPkNpmS8y6soPLej0iCDzfQpmaGJGsteivGn7WkpP+T8cf0
m02Q4VZpPPob1CNQEV+uOpKUm+U6bWtdQIW2heRySRRQo8n1SYyY2m/WA/4Rr1PP
iK4dhTAJz2pnKqyclbDqisGqB0D0rdIqnXbg4wsqXjkP4Vo7oyIhcMAw7Ru62gKQ
5PPiZmmdiAJuUZVxXPRam92r5pSK465SonJ+Im+9fV4NaiRPuBHJi8dQlNNXSDwL
/YudiNQM2xdODw+7bPEoKiQBYQtCS8Ib8pQdIrEhmECsG909YNPL5avaG9V2upQW
3HiFcx8FoQmA1ouJIByIqNGzMxLd7M4FWWSHRMpABypxf3rl31a4N5iBQyCA0ccF
+uRwHJbbp57PYgaO2hg7C0gdB0oRYL+H7JK5Ux/r6/9UlJhLXiP+P6asDTs3sHtC
nP6YJ3CjBVFFtxT/qqSiegoAVacvHJo37j7AitTgDEtR8YR4IKMexMIiBxDiHPtW
NehSXXhOqg5rIpNuzF4Ihqt6xULGENX11iPnKLo4X0s7GcrhXXCk5LwSUm1ludjK
ELdtfSSKLKZ+JV6aGSMO+cUPP96IEQKHt3ZQAwkOunh710UAA5Hcag5rTDq+CtMh
3ZOYlUYmNuQH8ubjU/G0Ytk6+rhMRNHn1fNvPXJ9g4owTWneq2etvyMMGgVWXA1p
SZPSEGRQ8d8qmGfIhOB5LOv+D9AT/Q6zZxYxGRE55Zd+/QZV1pf62HtUQvxfgp1H
itK3r4ymCe5vRHLNuUdE4oxMciofqnZKI45zoS2OdSo+VyStxa/i9hvAb2uuPGkR
kGcqXRL0Dnw8gyJxLGIDgijgkr5WG9muO3v5jh6dQg3oM2EVMKarEhgpwdgNqqRr
EfurueAbbIZ5fPSgnkScFPllfnlmKAXSHABV++BdRluiH1I7T0xstw1gNGvtS11k
vISegY8Sgkn6INbV3zC/5bhUuKcjul3hu/cI89TtGuoBEHSDAAITgRq6zSd42wtr
7oscIrOmGSvt9yQmHUipxf5ye/ZTz0rI8rbXIjRHUhs+p611TKxBwbBo1F/vV8Nv
NdppOL/lZvrbKPbuUWRwuoMEgpza80dfJmLOCkE4HsyZDKoJY6UhsLv6TcuUcgU1
5bYmxZx2P2Xx6LGNa7Gp75gbfMShm0sFTDhjLWI1U3Z2J4M6ARh511ajJYN4zB7k
R3XuKno5q/5yfS5AMAcWsiS0pjXA1WszNM+hTr/ljM2h3WD73uF3DGSc/cua4IeP
aNxGixwZFMnkkQMTHy/BeC1/2ENoBZyeb373ZylGBBqkpubanMz1n+3ZOCDCY+JY
kSqXTjZJ2C5AO3HkK99TsafgMvz77JuyRe3QmWXzVpihCq9vnNkI2R7ifGfEPDQH
Om03i5kO9dPcavqZTVzotTORQUVj3ZO0cphwwVePOq3j9fKTu9uVH2eYMTZWQaPH
8L5kNht1AX6p0KidIDZurCrDe7nVCcrCfNv9IazEUtIWVE7zVWpKB4YnbPbwx17z
6nGEh+5V+465osTkMOvRKEcFWqxjzohlQInYNpb2eKyYyESHkWCT0+dykAR3e8B4
pIyTAeGdZIPyYcqrgbOBKpXCNlEnrbSHWtI0LGX8zYrvHRH+5ng+V4qaoFm0Jml7
chIEbAoJ7FJQxDxEibuVobXeHV1N4idWrDNPZt10+2WQHJml2nFgm56WiWoNVolz
0WdZYlavjRCkSk8ovkZrl4bwEm2NOrjfiP0aeIifCWWb8lUpn0ttbjrCqwUFLODi
dvFDNP8twwb1k3A84yjBke4398UXQWk6tUCK/DyuVwoyOc+a+1WHhEBnnnJ+W+79
yAFq/Zahj+3cmtMY085ITwScOml7O1S6o+RdtSP42mgAaeCSzlYP+xibHGNmxz2g
s28c8YfWxjM7+nDcF1Gi1pVTDU2gi2+545cGRT2r0ez/o7v2ckYhrA1V3fr34n3g
xe9Uu16SaC7wd37Imx/t+5xZrPtXPqiUrZA+Zg6qRaISSqO1hUSt0IZK/3b0sdEW
xamRiR4Fc1p6TKJtjrGlsBLW9KhXbhC8Klfc/dlC7begXtnKAAWXp31zFj5uySLU
SGltqcYagc/7dCQa+4ERtmDPQ9d/hnQhGMfoCPP99Qrzlrm9eMd2HmZdP6JgItd+
ssb5Ng/6J8wPvilRWtdt8Ysqy7Gn6fL+RNb0ZOaqM/Jiedrv0roH9h9S3wVUQhxb
ZZfzxwnaDHpm74eBoZG0gIYOAPueHKFPeMWFGdI1Nposz8PVVMqRekDprzBI0K9X
WG9xoFSgIYnUWlFUTjUeypY9rsDRr6hKtzRmTvRjFpUvLVmebY+tkE2DWzO/Ykyf
9U+PF94SvsUSg0YkUUrr9iYqaeGMJeOF7e/rScnKJzIK5cNGtsCrzEZT8Nkti+rj
WcBylJop1m2Ay1keH8bD/VuUgYnVvmzrnROyeuH1isiUNVJVxNcFVsiwcN54kuDC
4mZo29XZLazW97V84lWpFs9UV1O8U+8NZQGuMdEEq0YZhuJ1i1louMVcc5uuecfG
sgoXw1cj5og7oqrN5yaCc9zNqImHAKDvq9+zu8yoElXzukBE7JHrrknGlCuZ27h1
BJpXCZHRqWFSBzbG1pwGajH1xN1RkW9H4CWmzlZaS1cHMe/LUxttg8Vt2XEM1EUz
Qba5YStw4NloVejzhdWUwkN4VrCjIzX2zAV7rt/Vqpo8wgKDbxwShPo8ozzAO3zZ
UxZJYMWQgvdnane6jeu7ps3ML734VCxLYwl6cN7+4SBjo3mr14OWjOkef1yXjDZr
393UWRfE+X6YTsPqmR/rFtU74Zgts66vdjXuqR6iapxYW2iRNZE9l51Hm5WURJs3
Vrlw5f3PgFxgF4jwwclW8ctulj3HSWkxNBOXosSOLndFhTC+06yzhhaXjJsTbdNV
TT9a8WuEy4krA59e+VS1F0HXQ2tWlSpF8BTtB2IHrnZxcG9Yj8IP+TIl2iHomGLk
VaelpsezjVTFYLRNxKs+cltK6JyMujhq9HCckERjqn9uGypMl57xYr7h95Raj4Of
xr1YBz8ua8G0hDhFoupFfIg7ihpFpYLyOqdJfBRhOopsXLs0xDNuphK9q0HsC9yz
jxIeQsqy4Kzzp1cFrzAvol3XSxvV1N32MoWC5eN1HiIsbe+/kXEI9j8k86gWksz8
UaXCXaybRJFBhMf8uZsaSS+3VpJgfWH5oJ0+h6vDYhjERnkMGMplIhZnMtVhmzQa
b0hzdDUd//WeAb0QqFfBro7SMPmdWF7I2ie3TDj+ROtHlPnG8tq5bPY1ObT8JS3R
y/aVRp7D7x0OmjZiE2kx3rqWwVJzClqmi8wEFnGdq2CljOb/fLOK8nW3OJWjbXNx
5In2NpOJvFeaNMKFfbk8h3+L/CBxh7oTtMfdSLTLFimHp2M0rTH5pM37eV/x4nyo
uRTuWG9yavqijfPTJzobxIXfi0r+o9h2AMjPhqYGz308dnKBzxpoHyn8JtF5e4Ab
J7UmzJy2rC+5CdqXiFTcgA2sQPFnc9/NNbCij6m2BoWdv1OqiOZ6q2EmJQZcvvXl
pluJ9CaUUNukxZkgAp10vF7KiaxS9YN19ekbk5Z0FFQB5Oaf+YUkLSgSNqdR8xrt
4W+Fgsp1PoumVd0XMvUPcMe6inFq2qB5Z/HnLX8WVzXAna5M6Qk36KyTowbm/AZI
KXt1lv27VrCgEN9YJznXXF3Z5xJzK29RO+uj8nWjRng+PwWqIrZyWfIuuAUoP6Nm
bDkso2PWDVGqR7A8LHMG4k/boJsl8lqZg3ms8czZsXmRBiqewRo+GeeVaEkieFfx
hfhPKO+5s3wUeODV32ITo6ktK7ZwQBAf3PuktV6fX5h4jIxMrOdvlOyq1+TZSAVW
g3SVvboJugRiHQDcBitNtsuTNAZpGr7QMgHX1aU7hR2DKwF9ZEDLlIfXR7R/04YI
/oELYCZ0vdph/E0hTl8GzjZQwk/4wd+USUfpJ3jP96SQgnPfIEbhTfiZNCwCAyVr
3PEQaAYvw8VBXAiS5EqyYKpMttQpSaBrKdg7ioevccUA6cl9jAqqFFZ1WOEkGTvh
zuaJJPq4PlHmd1XrF0ELVgHTuop+zz+sjZGhJ9kJG863k7KaBhy+4ZPk+DPZYFn2
C3oFHZX31ZvWvl9+JoAz23sFVp7Q0pESOf2ru6RF+wsVduVYOclOsl3GL1uKB9Rk
GvN4tyQpGA6VMKBxi1TFifHv7iK+543EXmdrTYVaR8neNU1LKLpAAfDSMjQlF+Cx
wNqozVuRVK5fbgh+3AfKw1UwCywYXnnLn4sVJUJSJ3m9k4TT/1UgUdTf/9e7Ex2F
zltVIP94kXlsaIOVQXMwti5SEvjbmWqp6YmeEEvoC8W0XvC0XvgvUN/3dUIE6ptZ
ExHVQDzIPX06y4v54je941HUij67O37WLDdzek+B6kURIxA3ZO+NKP4usWRcejr9
ag2BoGVLKT7/8KiVXeoGZnhuIQaOdwxD06tWeArkdS48RQhENd+MJx0DDcXn6zUX
8LG85NXR1ZYm9MtS6CSY5lap65w6qZaBUu8wPEM0Dm8djiNj2wW51t5NV+JVWnJY
1dl1ZiuVuFBNpOi85dcFqmnaczCZx6pyu1ltcuX008ZzzWOM/b6XK2qzNXoNds6r
mX5rieEPc64dp5/8A6iUlj0riaGOWRc2amVSSE9bPfH0+98yVPa/4QfXWQ76HNxd
a92D+qBRWU0DIUSC3DWpTXsEdNkvv8iORt3wDpD1sYCuU/Q0a5fV/ejSaa/OsvyN
bJ8dLqnzpnNWQKCosoHii8GtJSkQnr+XcGfpZGrqhco+L2aaFbEF7BxF+wOtXcBH
MdknsM4WXSucDrJc+4eSgLDCkpNwDkLn/lwwdDNC3TE3r3dA3hu1YMArVTifhXlw
o2tr9VVjylUbsMziuBTE8R94oAScdz8rKupPZF8RR8D2PPw9D0BHx0eDo6yF0y99
z/mhkKSZhzhMsnGtI9MmDAf9H9cBEMDe7UToUWbON6WJCPaFGA2IH31xWY3zOx3y
5s0sC5Glx+EPBqAfFedGyzDZ3yaL5J3j6Gv+LOQQKBYmwAvuHuxA8OeJOIObS1L4
pEvxXum0VT1PULEwfAo8yYy+lgkCwU2SCyO+KLxZqE9Nb9oKHVi4Jtlrqs9Y1taK
8eM93jtrUN+LgKHVSDEwGWovdfphrQyTgi6QurYgav3p2kgmGuT6HjWBKnP/BH4H
jp0heNIubATGExnr1zKsPznAdukGCmRNd/pMSswMd7athKtEGfOEQ3ekIWa8Hbnu
D/Rhbxh660+ORlwCyeVRp0iFe20rg26GiGtAAAvHgQNHs8uTJW27ElldRmN0akHs
bfhhhM/WoWyBUpC89scm8VuVXUFWdbnIjcWNtbFA+/7BvSvvG0Ro8wASYldftFuP
g5Mk7iI+FYguizWUSpKAm+p8b0Xr4XX+41UwqLqNF9l7q7M6GBg/j+hyo9P/u3jj
9t6USZ0LbfCKeavRNRa5OCHL5/w+n85x2NbCFxjClwv6J0wKDJ7fpvCoCU5sbwDz
0SIz3TpA+yhREQyZFsyDSeoBQ0n0uDi0sOZ/PNuUzUrS+c2iYIvr/fTw/p4ABeoQ
paR14furqrjV75CwDw4ggzTklICWsRUOMkBX6ICAx66B/7XLnCZNquliAp9ndE8i
hqRIsw/QdAeqJ3mRzMhNHygSOVFU4KJFiQ/Ns/eShWoPALFDw3r3O0kps91Ypwn3
oSMYlWNEE/YZ6W6Z78qqma4ir22ZYvZHr+GJndAlaw5on6wr0r3Zo0MX0TtsZZAE
5opZig9r6L2chgAuQK0jThqGNRJsbeO85UuU6UVbDlN0NTNsS4owvxN7gX4Qksk3
UoA/PZ0NmAJLWMbCszzBNt0GBXpyMRsYSSXf/ht0CtANxM7NV9pUehxu1vjFI2CB
HgZGyCSWiSlg15Bbb2yrUdcYH/eI9hHl1a7mlDSEB9Y3azYRBpD1eHlaq1GgOgYj
wURvIAOa5ouoBZdn8KTK7z8K9bH0VtdVAo9K6lMrSvajCvX+stcgqwpR8hToLk85
AiulWBIIhReu2AX/T/RU5rW+YlDjZ1nuzR+RQRpRqO5z/lOf37u+iqTYq4pFXg4s
S5qK48tyvIPdS9xOXKu348HSfbwWNn417ohRtVSL5pKzbu4ZD+Sn7ES5mVI3O33V
ridjow9kXhEmHYZjVg0HaHZ538p/UcQKVmfx5gAIVxpj+gDg6OdRnKt6Q/hEdxEf
3E3YdNudTAxEGQ7pyc93ekF9aU/SJdRm6Rs0ibnH2ZvzBdixZm4NHYaZmKYPU51w
PmWDzi19BTIylIXdLCr3cOQNpvdLM3MVyuCImoNAXlANziCeOPVqQL1E47H0yzpc
gVtYwTLccWamArSt/0sR9LjICg8EllHIIkr0Vna99LvOdzh8ymK9GkJxlA+8yKTv
NBieJ16VxQrAE4C+OqaqIUtiPbWa56TvavRPuXYMgIT8c5WinxvM9hUhOAw+i8zq
kGKfgQwX3mu89JPP0iHvZlLiKAZqpaB7eHh4F2ejJXDYmJBjRy9CufVQYEcngddH
3PtE7d/uX4tWuc+Ew1RkvmLFuHLLi76C93fILDCe6EJ1awc6Q90U/7+/yvwNvp3a
S3Lnm/ULRBJoBD6+h4DASGU4yCfflj867ssD1FFEaVb0c9ZvLvvY8pr0ZLUQ9ZK+
uU5oFUlQmHO2oXXRBOEskSKSvKUNCBbICgX0piW3K+oADUEjSSYX/nqL5JpUn0CH
zKfPYuVuTQfZkSlRuS8XiQ0rE0sAmncbjodc+Y+ZMIgC8tpoQnpkUWX4tgsUmRie
5Wfv6K1AUsPiE45ABv2pwZoBNMeuRTYWuJgsd7DRN1+W2Kr5TSLw0JGbPBJ9SAet
UNm71sLCsrFxl5nc16PY3bV34GzzzVvjMJokDbJhwDtiEVlZaP39cFpLA2klkAzR
cPS9FkGBlvjNLHELJ+vjiP/oYMkS7YVOQ/iIMPsgqHa4rKfOzgwcnoGlwzRr5Md8
M+gyJ8Hr45CCOxfm04paQu8PU5Nyie1BWLuSyUHfyinxBfLIzr+8gQhVSFWirMHB
8PdmWsILH7dJKPqJy3IyitFRojM/XWxyJ9K+yunUeL9YSJmKn5H8ukxlcxi1WQQq
v7bA+dM3fpZ2jqyWJEfhq5puS9LAgyVDeHTIzioixz0BAH+cuYVNihZwLkF/YTCV
w3gT0ca6wahe9b9sbekdpDrHqKQN813+BhVp8+1Rn+EpaIU2SZKrqIiv69uIRStM
38ynrPZy9DdYE8uZQfsEAJqFJp5gXr/e0ZK9FTb6kreHS/p3X98ezw8IdoKAAdZ8
3opuscKG+ae33S7/FZzoarF6aH5qv8RqWCQmcn6EJ6HYrI7UpQc9bsvIgONjzMue
EN0FVDHVX9JuS8K3RIOshARbevz6aXt8rbUlYJu9oug3tX+dvvnmYnoIhzf1h6TP
o1WMBHzMFQpkqkLDXsZNsf4sU6yFTeUdFyCm5yh+Ffl3z9eYzd3lOQd2Q8PpRsm9
/fSd4bIeD2GBi9jQ06OFjO+WnBh4FWVTve1u2u0/Q93RPiAQCC9TsvqmBIHXoCb/
Z2Fzm4Cg5DvkmQ9aqMZss9e6lPRebFcYZ9wM5LAP3+QxbzgTgbAyFel+aj25i9E9
V/RW0zJO5uxCzt4dycDdYRcUelbxlhRm1xZ69ka7MDh3ZcCnSe0x1zZd1AsNQxgb
ZFih8qtlx6JmR0i3B32YzqUQA4uAJyU7E3XDYyLHwQes9a9e9Xk8BmOL7z8GEB4u
akImr9btL+Np/+F2m+KbyyxJEhaNlGFQSvbHa7AgMZWTsKXQGoD90wCF61M0rtls
hAK1lOEVLcX1/LNk1ky/TpAoNt4yoJ1f7P45Pm8ZUTaJ7euDz4vt5h1cUrTdyJAL
aC88sQ3MB2shvUl0feB8UdtWI1DMqaoRSOMBMPAE67LAcIKPq8tlUts9q0Vks7Cs
Yuh3wvgCFzU0kfkT56kTAy16vNA3KMSvhnWVgYO08UhtD8WpE5ZlGMethH3C9iEH
n7gaJ3CBBcXwQ5S2w029E0Y9wEqwQ0x5Ks+gOPfodstuPTD1GFIko+EBlYS+BGcm
gRx2bninOsxW1hPAsm5ReacVSO0HSXITfIbcHNWaY4c1PQ8dVGfZeoUg7v+6xILZ
qw+SDVZv67xrhhtjfFKJs91k4+hdYPWrxsw8NBerx8GgMBkkfX+yzLoyJt+U34XI
4UoOn8dy7UUSqGJ6ofRSQ3UPHK8hVsv+c1FEO+BGrzj71szrFcobeC6J7CvrZcbe
pPgqcSiwo9pNNy6887xh9VBaFrI3RRhIuZTFe0uDCdniaADmuPo0IDLSwVAggVoX
fcSku1mpDHZkbKCG7qrGbMJgItJVUFxyh0IrkYYCV09N8m0osCCiYbyIvvC/BIt6
EdXL//p3TnShpp6SUXHuOdTO/mfBl+mnkby1TvhlPIJlGC7yx72c+KWMry5myQzN
6JNfN64XzapjUKvv3THyrX/71e9D7rYY/3R7Qwb6pyrWxIWcYmYKpcoyiy3qZOSJ
fkLX4XRKCnZoI/b7c4yd6VvQIhm31bm4yJclPLMTQTc2Tkj4lwbUoE18bHlrouW3
6i9oNw2gjfzncSb2eVm9JSzy3mBFSI9p71xc7x95i2u1Ivb/KvvMw3BtH+DMjotL
+xmMz997x+7Wb0w8/1iKaWZ3qYFCQ7u5/ln34eMrFahLVqKBRADGQPWL84kvqPjc
n9YMfut5tyKpoqw47s8m+Eqe0sTyvAkmLC/OtEqTAUrgexNghDkt14UKRh+bR27g
ai368dP9R0kxQ5p16fAUgZTm3H8qQbUIP3Ds0JPoyk6+tFI4O8OclzUTiNPnYHNP
dVP0XzWYPUU4kbQR1AExCGNbWBkyu+nLXZqnFXgj2HPFeoYDIwpUMOVURYOJpu4L
EEyWgW/nVQeucSp+qELnV6/QH1ccf3/xeWnT6DdN99g7KBvJ9lLUByTLnn7GnEWH
92/+vE9Szuw6zn1hweGYKmhvNYqv6v1csKFj2Bwkv7LZ6wK3ybRTcBnmSzkucbJH
ptR9Wh4MIRxTX35EFnIepY/+zYD5RibrLlMM983Jvlc1667h0eT++QrCr0WrmNCX
wcpoVYML1hGjuVfu6G9bQTXlkx2FOcLc3JQlfDFzNTimvyEc6NS27sXqFGQ7vyKS
C24Db7hSpn8uSZaLSe2pyhhD9Kzf1HIrFGl4VqlNPEmLg7VgQDXXp7bD3ysK/OS8
GLvxTYUXpeGtXcazL+O5Nwl7cLZqG+b5sMtz6b/N3T0zZtevXj5Z03S2V5D6EKrL
XoOcps5p1PgqnBcIIK7Bmjtis3EfJ1UrvcYBHKuPRkCVTuLS7yd5wpi4FPE/SOdE
phPJ0KS9dPpfafxarrIzozE0djclka67Bt0hyzsA7RmuSQuY/0BXzRVLxK+vO4AI
EHuXf1tbVR1NbkoW42NFOR1UfTMl1gH4wKpNaGLJA8i9ZaNoBQtZOSLaagQOlrhs
vNScxFSmUh0JdVdtZuu3d1W1PirpUsRabyg7xe1OarcJ9Ni79u06NoYLO+94j/N/
ApddnOSfuuY6BLzmbY8bMFe6fmpwV9euZKe60Sp0JifWmod3gmLtMRzktnVlbHSR
CWWz7C79eZM9KZR0uOSP5/hJ1L58bukZtc1nCStJ4w68J9YbeA6Vw0zW9KIOA4vN
/MMtGJjF4Xiw0kkVr9mb/yYO1BRLgYd3l7nuhs43mGpMuf5aG9MpYaYtd1vE6rYX
m6v54dQ/kc4D9f6EfNwRr+xTjafdqOaro5hXKJrueRKvCLgOTYqkLVhDSlSUpuTD
K13pyk7reTx6n5lQAsVIzdGXtxBeDvlNUN/mgvMh72J7slYn3Q/igWpXa6XNBuuW
hNB2qF0WkaxgEUxPX2gYVFvox1YxfgJzfKGd01Dx4IXCnV1c0PEBomf9F9HV/qko
Xw9Qub8OxUrGSYvxnie/eDvTKsfGWZNggPS8rpGolSP76l/2qoGzF2Hkn9Hen/kq
xSdHlRMoVqZD/PG0YbMixqjqqwCL/mdWs86CqhxR9TvhM7oRzrl1q7RaWg/ndKi4
ylme+dDBx5vMI2Lh2ep26QkvbFV17nc0V7BN3td6g8qxJdNxD79YBixeMFW7BssW
tn/mpixS6nZhqxYU/fEnzfBxbYUbP/2U0xqAxCAD687Wlv+iiJ2W/dStM8ybHyN2
muFuRPlhTz4l+OjN3WBNAEr+H4csEUJoWjuDF6n/q3Y0vXSBzBG8MO5k94/v7LGk
ONHXaY60E7rGYbPdSc59hpjAzANIAZ9ZTZ4LVX9FQ2LCdonWqqPM7Ni3qMKborB8
1ZtJYMFvv5fR3byt55MKWJ0ZQOR0FN6Y8YKnUhEjt9mopwWnTO2IMMFANC/zEgjN
iXMOSX9N59XgVw3QML0DpfawY52TpCS9H8qMQIoz/ZO6v5V5T5vjMfbyoC1lOjRB
cyxiunycl1Fiat6TiVe3mSFgpP/r2FOYu0dW6NA+gTDJXPyGjmG6SzvyJSJmUpUO
da2BOPL7X0MP5ZuV3rwTcN4+zKG6HJM96YuzwUY/A87AU5rjYfYzJ89i2rZ8pfpt
KxgRSnmTTdSxXltzkYM6Io5fc7DlDNQ413zh3y7ZMTSqipGnR9cAmGCvsCTsgv53
1LMFJNcZm9VX12P6bNceYzWlNbKk6bXqL6p/qO4KlUSor8iXvdkzSDLwiQ6T2fcP
U6CRg7kDUkShpRbl3KCgVr8NdqHYJOv4o3KB8o8Cn6yXsIFIxr0lfnnkXWGc9WyT
xz1bDIpkQk9Y724GwbifWP2EMcQc2xzaDQ8jmp3DfD0UOWt0qYi0Gcx5uvFhxawt
vY+fO1+Lqxgz+MhaeuyJSau7BVjKIptu+mHe2623+Az2O/4w2Zjzto+qBhboM6vq
596dw1K4v+h2vQ0XFUJd6HFnYYja/q+oAjUlF2ClqHLbqAop7uiP1JEEf7zdopCm
iNu32zMIFCVGEMJDY/9MKYaEEVwwZP3/YXDnJFbtPdX33g3bx2tguRDWKOgSued8
6Xko9VyjXVcW0btt5RO3e4bLN98aDZDTYPtYhuGPsDSo6HRc+kllkOJ8XNVYYgS/
rTvkc2roE5zhmq+8Z7MEuF/gBEpBW462aQJCXdSbM09njPC4lXTGOb7kOxkllOHB
3Bwvt3omZabyHzIZXegWRs4hZktKfXZNoa7YjDIMnDdMJvkJCmGAWq1ILeIcLo3X
0kDDgHq9LIeeoLwTUsP8r5i66LO3g6H7hcNp3eEatXR0WpsnfUkeWeOj50Goct2w
+QjfyGn0QrGm28yp5H0fJFOPCKQ8d+RR011KNhA9qSSe4xSORCJoO4BILW4jH1RZ
vPRYnn4lto+nFq9v21STNiHy+DEst6afeaj8xaPBJLvaJpLASP49/hF4WnCbWMrI
ASeo8Y5ZYVuGUB/zstyPsSwK3iyhIS29+8VQI4ZTW2Rr4ioREjpGX6wjNH2AXRjR
nN4FkbP09587P87u8Fc1LUVGN8x+j8WExoM3VKrhM3xCnUT2Atq4UEnXS0TLPl9v
4e8YvLz+9rygv90ZXodoz9ZbkFQ9co61KcMMf2FbO+o3oJMD9tUzQ7WclivLd3Wp
1ZQzrxBGZQU4h34jPKjMoDXhnvLuEaY9gKo1mVwqY0WTnhhB4PklxQyJ5CjJ66Tk
us3O9VsYJBVSdbbgVKZFifQvjkNJFoyL1NsMsZbIE2ZnTJ19dCCXVbwiGwN0ciZK
ev9ah5mQvoSTUCRoUHPm1rwsa3skK/HHtNMPy3maYyuld1s2xuWDWJuGCrB8/7Pf
1q4qtbXXX5f0PigDkxBTPYnalhrqmr1oLNrY4uKl8E0EUmnTu179yoQdIcQSxwzG
Lwz6qqzCWr5WD11JcPc+Dzw7TZxO3ny3NpZ8tQen4Vx8WlXwu0nTH2+s1JQTrpTu
qkckY2lytVUn2vG6FsWzO770/Q5kVBGb5WmXPqz+6Z5I68eKcvx8o097KkJ9pKNP
Lvw5vPu262J2gVcBVffl2sBJSc0uLLrqjJfOSOxgKtYSUBJScDWuhUzaiuuPKo/w
+pibBaLFAG8l0Mc33l6lchdLwmNgOKP7vDNombUaAjYkp0YV0qU78mZgCT3KeAVZ
OZhslFzSeWejDL/YWrZNQbZbBZy098hqn+NolGg9ejD0HlAhNQqHkG/kE9Qiw5Lx
N/oIPDdKjxYrgNOkAKnMsLhzi6uJTQ3prj/Qx0e9CIgLLBpKV3PNXOXRxAqCegnY
wmhooZofbtDURQZslIwBCFUBzof7Y4ZsZOZejZwuVCod8oiSe9G6/jpXh/F7eEOT
bUWmMzYuy2a5wwyeDb3vcZqKbLYiSU6xszUZKYyaAYpBDyr9pwvdMvYf/QUVaTZ3
8sIg8NULOEw6ojGZDNZkwxCYHEAyGZhvTtJ20sz9qgJH7hGDx6w0gVXGlssmz1+Z
IwJA4m5IWkAyu9OKjZuPemQuRA0jUKEPEwP82eoB7MVNYtcpe3tLQCfy0qwgk32d
NJuEB89xPViVl/W8DD+PwJ4kcR2GgDCG2COQHqyPAFg+j+0itikyxYAl2w6kkZOZ
b8s0ADO87J+Tk08jIjHvrDhI1rOd6tmvCewG0pxvTs9a24YVv0BiOLuwHutUX8JB
9EkmNtlVoutazGtKAgyhfGcF2ZgIn4x52vkgZQAXFENz6gWcw+lPCFkopbp92C+t
qo0zI4FMbGaW3Bpjs+yGrelSPsr495KKgJ9eX6+4Z9uIYvCtOEpnQns4ynkRPg0m
955jsOM7u142l9My9MNPY4BZrCSKEYXP7Ni3b5+5YPaEMVJ7/qwLjLvaZuMGBMBD
/ECZlyhYzo9JwwexZjvJgbSf/GrJj+Et38xxiJuKJlAA0mhG2KACwcJcnWI+Z17N
z2ochN2tQWdF7il6XKMzpe5ZEwNKDVvRUDKwtMERuRqPMeVKUGKYHnXSBFtie/WV
K1OjKYGCBF0p6/4JHMhvuRkvuQlDGithAtbT0AL9mW1t0PBZ7oVVQ2+d2XxFbtIw
ySK74Ug2VAi7VhiqecKePJpXa1keSWglX/XMPVKcNHzmzLI8ipQHOma6xvxaJaFz
xos9zX7orvEu8WnT5B1Wps9vlApD9KmrIohMfuSxDXXTUa5gSngQL2OxZDlgpokb
juYY/FFD23lzp42Rtn9SVNpPSoVUgJgmRevWVBaaSUwNpL7avGS6hpgfz1nzJt17
We0g1KXwEiP+OvNQ857/jCTcvbg6D5GAgETam5Uob2OceB754IcCb3y14KrU2/jo
hvaD/XMAaW0i78irYo6KEN3sygUCLKSdMUpGz1+j9AmptAcmdpbyrJ1S0nbgnepa
j62f83SBieBfMkjI9Ssavhim/sFo9zf7tbZt4RCp6J+GuQmwuAWZ+MG/bwkS3HnE
M1whK05c58lNhvmS0SQ0nDh6vnbGLu5Q7fasAbxPcGKjG+JpbrRtx98j0aLQe4V+
/hJh3e4O3CFFJ940JIXBLHce8OXCJaSkUtOgfWnwP5EI4VCCS9MO5lw4ZV/CA7Hx
qxu3Gj8sfryPRVZkGAz+jE548ok25ZOAY5NGaZ/XNW/c7S0CAt1ESck194l8BJ4z
aLi2qb7DMy0wQZ10ii+6yWYOt2oyHKIpAeiCrsj6aXWHcuaRAWs3gnG+UVswDLcz
Tp9f4dqgyx8qyhKF+AvCLeLfjHDkfQu/OSLS+XpZH0He4Hq95vetuap18T7lqEcf
ZNcbvXNmMK7NKH18nBqRzbG83OzM5odWXp6faS2Ru9exDgjVDPUBYMmRO8SOcGK6
Cm1GbVAalOqV212UDBCDS/mrjBOgJx2ZUiKrldGcLmhhLSNJxx8xe76y2hy/S9Gm
iNRgLUHMealLtuROrCzJcZSMBJUaDWUN6z21FtMbDLH/v2VdMn3w0TntZS2z6lOY
NgN5Kw3lT1KGvENcrA9i7ax2gvF+0ejWiXlBUWAvQwAirHZlsi9lz20R0Ly1Kqgy
Eri9Ibuhn8MPg1bje9HjOIFJyuhBt+7ns3g0gNdF9X+ZCOX7+uInNdUEc/NkLEAi
lTzYeEmXh1/ySLsK9nIsM1WKfSXUS5Acx9vLPjwpc+01nB1yjUfKVIfZigBrZFd8
Z8aumQ5MOQRhNBelAVut45MikFkrX82FTNJ1Mzt0AKmNyoDvuBGjthcv7L1rRw/w
72ZtB/Y3QeEqs6OuhBFPqYm6RAc6tvwXbNeXKtvnJw/A6rn55O+reiLRtRCieE6g
TQXAX6nvnYEA0LybzDz6wlKh6J0y0LYPO/QyAOeeDPLsETr52CyAuvX4qQOVgFud
UF8dg/sDhGH1wL5O2bgl0RAXm7Hy2UGsB1tQhsT2ssMOHqAMatE2VQrhM89HbpwI
8qBEVPyQme25N34UFPpc4DyOptJZFwxBQZJb6dG9/nw5ZR1kfMW2Cx69zcmrrsn2
WkLdQ7h+vQ4c6ygAW6npHx5W5ogof5x6hOqHlC/bXjTURmqs0WM8HDytj5caFPFY
UK0Ax9DzxwpEyzWGzWZgv2h8lkhYZP72WVXiQlgovHK+2/rRW3fslGPdLrcWLLMl
Y+TZQuRl/vEe4PPy9SPqnS+53PNakvqj2aw6GUGZ1I4s1VV/KvAwMlY33x+S/AWs
RpI3duEWhELQ+NXmoxmmv/rUOthz4USryDnrKSHQCb+iBjZFE+KuZ03l4LJfl5Ch
d4j0dvwmPxh9tOdZN0TRTYS/MnpBvVZS8Y960F4bl/2BJ9rzAQLUaUVe8RhZ/+1U
0LJ37scZx75W2X+0S2Wv0twIyD6Puxip2PByI205vw4ToWipXbF2elav9+xXYLoh
fzdnGzP3ofAW2uVX2CPI9j4GYsXf7szjmce7UWYuvXdAKmA86nUnwupjP4TBWgGm
RLCedj9bk1n4EN80iH+cbOUTlRRiWscpU18gXO5vynhIo+eW/gERtD6dmccXgBAj
7liaebyQeFLv1KUWDpbe3mKVfScjgE0Amced33A/K0R1TtDq9KNphDEUZTZN9oYu
pms+KsqsdEmJpcGPGzNYho3P/Lmpuw58jj58sZoZH27d1UxVaisYorrR8/ZRx5cF
SX7H5QbrkHvqUO6KjWvQqvdxNXEAob5o0KmTLkzotGiQncmUI+6+i9ZwKo4PwJaf
+cudUJ3iER/5sIAIvM6x4X2c8no+4rJIghP6UX4pNrOAj8CE5tayrWf6ib4133gK
9dOeU000iA0grCNq0lBMN3u68hrFWQyf0WfO3Y0jH+22064dBNrgeWtPgxtSDE7g
K4gB2k0Pn1KoR596xGyqtWsRuZ41IkE5d/Xq8v/jqu1kUjQWqfbivkFzcf25n0jj
4kxc+I5uZtv+ZcddWq8gyJ5TkWjS8Q5cjbQZt7TE4R0uDRGuHznz9BMZhR60EH3q
YqBoduNj8/RUu2q0Bk9b2TO/EOsxyv0DCzzBxnTorRJibVJRf5nkul7jV7pG7YiW
7PZLHPiWWxYuGjKADL9f+RGLnrBzWNGddPFNySMxhkptRX7Jlpu/DRgxtHXHPF+b
qeSVLEl+DokWvQ9dABGO6AJQ6EOxQsNEz+7fKr1GqEMY/iCW1JmnpMlOUr2G88yM
DtCdm0w/dJlcqE71qE4qAOwfuQH125ORKUAQAnINkC2bMbUsQVwGv1vQFdKO4clW
HGwXuyuP43o4VplhWU3AmF1Wde6XQkHuMowpfSF69bpsCQo376zpv8Hv7qO9Pgup
LlyxioTwkw3zSpvIZEBOU87sunSkyPRJ3i9/+k0da3acI1F/ggrDBF3VFpSw9N0y
amLKX8+6dMY9sH4sMe6zSdbmcrRo58dHFa4M182vQTpFHY+xhJUVzc1A+0LS2ycI
2Xonx/NqpZ1Aou1Dd2vkj+1CHH0Z6erWnQcGink4cYTrlTvAyNcPtW7c1EJ+IJGJ
CklH0vvJKmv2wJDO6nW/t1UOoZ3zzt/KxCA5nh+iKzR2yVEagkXew8/E/RJl33Re
xCPIJBytWJivBIVo1YTtJNPIzfw9Ld0xVuepMmlls9hUPYAwII7iN/bMQwExkr72
YOJc9Tomc9EuyHE6a8kRs2mSCzKo8/mdGBojZF1in8hL5O3s8B5C5Tw9Xb3yIEFV
GtR0It2og8kqmqp2UjID7EzVDMdFGuBOFb6CT01B0JDC5WrApij8/EDlL4HikcPa
SC2TM3GUGqboaVE8xMTSDfosQlebITwbo752QenvtnES7JxxeeEIwsOYTnAttyw6
DNWIOZJ93ziZE8bIVd/BljuM7DdMAFiHu/vdHKAui3C1Z/1smFEECvS0Q60eVSpQ
+EWbL4sPby1CxdsKzcnFxXlh8376Y4iw7nFOz/Ruom3FsUPXWhd/vh/Edptzv59Y
HmCay3JkU/FF3XuNouvcOOOK1qYsGj7h0FlZ47Fo/kJymPxldZGwteSeWZibTZgS
/oM0taqXnq1MFKUZcpNhABp6T1NoolZRTvgZ+9L9gclS/CGY4JDXdLxm6vuPemod
JLyqZ+io1S+DK+c9FjthLz5sfCeFF5Llrh63yh72OASX662egLCHGTa4bmTvfxBK
dPH0uRkJPRBCSC28WYQP6OYqoeZ50+wlnuMWzgJ4EHNaxsk914Ef0QAXT6yTsfTd
FWgGSWgB5VHc1WOHft/b6TzVsR5Wagfpx4iYrwcgMq7FXwC5UBe2suzpzhp8HF9F
IlP4FPOSTFDl73CMosA1b2+O+hxqzCEm1Mcj5tM4D9SxL5gDwdkOFucp5xst0C0E
jHdp5O8P7WkU2IbFWSEyz0WyZQtiZwRTtC5XlfHbp99Hzw04iDVkEcSuneemmzIU
/5soL+lk79dB1qqm/b+3SFULcFHNlW8L9kzTlvychz0VPlx/G5S9SJnHn9QJQQVl
0ADwfSijMp+CVZ5J0t5jfzV2FWTQouTgfoqrNg0S57BD3HPhxrjv222QJvFpHWP4
Ep/cMNJqaNKh5zzy2yNcSIWOKhCcX9w+J4n0s0mzU6LzJt3c4i8SYFm0k4PVeVBu
B3BUeCaF31smzr+NqB25ZHpk6YEYKFwm7ErcPBdQgf53lUf/T+yFhbxNb2WSrd6R
3pZ7ByLeum6vqJSokBqkCnyg+dbkGuIFOSVYz4F2v5vQ7x1/YN0hPO8ccU32qqMV
JDLhjLFZgFEJxCeMhqaMv4xr4K+rCaj5U4p6JgW+CFJOJw+fZaPARvm2mDmFgjFC
zp94Aq0M/5iHNTybQTT2mTLxN6iaf9kEepAG1h/Z0pVW/Asvii5AdK1yr/YQDaqo
X3WuShxlVvPpeuRtRXf+gq480xEC7c9rpGx5vZ38wtPnRjTEU/mNdVsGykLAjbz9
/BhTg4KzZmn083P/8ckamRSx07HtO9s703U5X8zv67AuiQ585gfqyOqk8UNQ7+sE
R9OZgX5aKbH19TjOOrw5FsNJ90R2X+RsLdo2G7pmZuFL5sfViNPfYg6YNqtQKlMk
GCFQSrrljgOMJ07QxqiCaAtlkmi+/ioowI6nNJEx85rHW+KgteF5SgZUJoEsdB+S
1fS/6xL7Yq7L5X4qWbzVGpVaZZtD8W8+sVyP2YKvDvCUTQ+xbMp13zIhxRmiNH+w
QGFPYr5m8q7sNOpoJjF/FBLMyc/m83cze3Hegj5nYxM1zH4EXW42pEHvALIulxnc
cqNqdkfG9NqOYcV140n0numrUUenaP3qoK+V411jEagihOR7ubQpiWbQD5Anuu+g
JtYRDpXcWl4JA1D8glK0yXilFn5zvagDgu9j2hmSC57zE79NlmWjWBPxBxA/Kd1x
u/2qsuWWgF6RqhKJS99EHY8wDHQSPyWDfyDVvDkWnjKSxWIXvqa/5JAZeWuFSPp6
5Otf298yQ1GPV+YEcwmjd/2Rzejz1f36JT8fXj5lND83NZ3jQSbNRoXrin6CDwim
EWLPVTuKTFLdyqBqDhO6E2FO5Mf3+rPrKGl0sy50U27c/b5Gb6w6hd6xVR+EXDtr
sURLQk7PIpYLlx+1Ig9usLaRnuhtTd4OzvuuXdIZkWUTzy9jhMune7oJTa1ff6kE
xYoZuIMIoxDhRLV+X2EosBBE0QkuFkQn5ljW2YEAdL1Th+wbHMEe09K+ofoSZbhy
IbKzxRNue3CRhGwYXHKa0FMd/DcaSBP1fxYuu+IGpHE2A/6C9U1fayYZC+MlpDJf
wepdFta7YaKBPcSR92XQp1NtudmPicnldD3S4GWMXSM18MKUjiWESttckGR6c1s3
TLPyhI+g13OMU1RMX2jG9t1ga+f/P4RPhQVdfZlIpMEDVqSZGUioIfbEfoayuVFl
RX+W+zHsqgj+wACbwbemAz551Csl2aTBhZFz+CSkztGMuCbXXLQhS/LGuQ6jDkSa
/WMfgMs+P1CRpif9olkPS4clxGBKTxs1S1QoL6MMQ8ekSWPr2+3h8rZVHmH9sObh
jRD+WVHbhg2+cWYI7I43DuIDKfGQxYerglz4Hh6qq/LUv08BkrjZBhVnly4LE89n
a4CAjB1UQIs4qmeJSn4C95x89+kCqUn9OV+BhwwwMzqvvI+32Vq3PYYGz4hKt9dn
efF2gdgx8ZUv7RYITlhJjiwpoD2aeD9EdjrwFOeEeE7AVh+/zjUFMU1rWlFq9vp3
gmTfVIf9J5gdE0qM86mQZwfC0XJ3r41Nm4fAW3f7jXTd4sX0piEr+nG5g+bey646
dkTrHnzJM3HfCHpsCMcJ9dKKh/qBUxwMiEhvJ7La2FYYa3LHElizO9H3Jv+PnhGw
A3WAXUBPMa9MF10Cr+h1Oao6mmuhqDGbUWSH45+Xx/+8QnAPK+C6AoHRUNOGvYit
kq2by8nRPCUEvv5RqHZJoYRW5v2rcdh4c1NOz1QxbPSKBsHvwMMm3ht9RV7AzyJv
ck9pD/hNe1OFxaJ1iMt42YkbKcRvz4R4wB4Dmh1PGeU08NetTdm984qeeUMXh2GQ
TWnUl8vUQSQZg6lP3rEgwqZiV4MjZqThxsBJwx9wNmppNG/NwlQIQcdBsjawltuL
+qYZsLNSKHCZAwj9DZv5a5mki3R6GBviDgZs0jquoXGCNjv6fGJ/LcpxIxwU++ug
FzLcjGTZZhoFaVKyhz10u8/K4IA1EsXu38ohaEQBIRUWT1wvxvmuTzn7ByjMTNOU
8SgnTVY4Ar9qdw2lly29w6VM6YdLwzhODoTdjaPiQ8/sMHUbi7PtTciHqQz+SPKo
D+hhKTt/oe8pLXwN1fwV53+vEdQEi0hYdswFEtNol3U7DCIqH4AsoUizile+ktFJ
qCeO892wPa8mrvRNrkPs0rz81kf6OS5baD1IMj4Kuc9b1xJKHU2RyIm66nPWwYlT
ix296JqptU8aN33J20HaF/+0PQMJJiNBNDJe4sYwWtMYH+8qtGOs7UDauHMSACXT
`protect end_protected