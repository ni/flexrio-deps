`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10128 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRvp3o8+RItkxKTewZIo7szZvdGo/iNhFVQmsqdn5BB31
cLW9sNftAlHSmSNstmtMZziDkGpEWj/qbYc+f9wig4uq9EXrBfNEyUvvMTUgJmlu
wq0dHooBeVzee+K/lnMtmvNJRU3O75miwXyRtJpvji7+wjy9MOpHSJiATyw+Uyy+
fvdx/fQ382uqT4uwFMNksJ8R+8CdjYkfbcBivo/eALRWAXp0xWuaF7OJS3uaOgjv
Ozjkmgp4O83XxuRZ66lgINh1fi8UMpiBkPSlDer5P4LoZE2UVKo3z25InU8Rclq9
9A1whhdhi0cBraRnnaG6bXIGfIAr5+DXhk++rIRAVxcrFQzaeJG2Et0U2SE9M8Ku
kfFEx63+mSJ64H09Xs+ZJKIdJYfpzyIcSPz0p2eg+5xJd2mUk+xNvXuzO6akeZ6h
S0Qq8VFgRT6gpuA5NQnMPUAUIGx0VXFP2kE6uxMj2rZyeHXzbWbWf6OhVQ/K9m9Y
KmbUAfslmwi+uULBp2ZRZDT0rq0CoetubIrIBy90VMnlWnwnZefo21laStIdczXJ
FqrMGsP2koiQHv9INxIzNZxk+1ImoVgdc7lncb0LxlDtM6HYL/UUqVzOOINwdle2
7ssuZ48s/HIl6ZJbvwttPWBJYY2k7JtAgjas+nTvDfBMim+c2G0mbW9hPPmbNUq2
tUHJRRXgHp7GnOm7I2hu2h9WndRQDlLcXNSJVcKsLM67e1LuFDf8soL1eHy8alnW
MjWjAbZ5Ve/0aS+lBnWoDrF68Q/i1RfKCAeo0FDx+j+vr+rP50rsBgoYYc6K7qiI
CJ0k2WlgIsyxwVlfpp6+jWL8HtiXD5BHQWC35ffGmTjmjYPCBQOxFaVzLFmNii96
hqu52jEyHILc/5zbc6n2ls107pGdtpNTyC2clBKDSbaoFgd4Lb9g9Gj8G2C2Fd5Y
KqbYIbrXorTSWq7rl0ZZTim/vMJPgMTEu57etXZND0h/VfnxvL/9ifpZm3hs5ipE
6uIupx72vrOistARKqSzRAbu71Dxhn2XTAPAEgQSrHrS2f8FJRu5xDXteYPJwlz/
WXC/Df765gxJ2bO+XY0oCxeS4Oi+iCbvMW/znKP2si4FKHp1ZtlNYRxuPMClBJC7
DAQRWJ+i9gah7R7aP+uI9ihHMwnDOKrgRR3jHej7DEoV1ZaeQgRUa5IbO4pggs/l
dgeXYWz9E6lk3re6Z2WecpCpr1KXqFxXds3FxGRVgr47gH0QUj2Qswu/SPRszK+z
7fx96fM2dmUBfN8N1LdCbrPE03DY8V7lJ+6FFbcpYh+gsyuM49ff/2WzKmpy5pO8
B2qJ3bfYvQyxWiYw/dExnXxJatzMsUBUKCvJorFVsKQ3hy8OlfTFDRnH/1clVmil
JOhLyGEsgfm20mJR8FVWR35IHzVoxuX/34FewpZehdmYNRHt7vpIHx6YXm2wDpDC
WvrV09sblAW9iDEffYucN1yMVTIYugiHTAWU6giXf9qz+6Sm7kXLq03M/HOusm5h
xr9rJuOeoGIW3U473JI4yoKSQ38aCPGj/cly0vrsQzt2U1MYQF0cwmLgwJjKZSbT
n1hH3VzslqzkWzy3Yujr36sp64/mTL0yRiNnMdfb1ZWkorvz2MMaaSH68dl891Ah
aDJv3+/Q0azoR1KFKd0pN2ANhFKfQh4dZLw+I/wubA2DHaGifLr10tnoP2tWXDkw
qVMiXDyUE4NAqayyz77VaVUs15K4+Tb3ZnXJE6eFClNF5kzumVWvgya35fV2ZJrP
rcD8TWM1N9tTARWBUVKLY7ejFKDDOsDTCpp3MWLPsa738XNkeqPSe4xu+SFhjLGg
NqCqzZmMoEIobnMh3U9o7FP5g/9MdmJNDKxF2HNk5ha93kBIAUnKRdX0VH8qDJLa
wUmhc1uSsI3n7JILaRrFcP3aE8xmNu9gQae2QCHOTn0Kue2QTubYbZFFVbtqBvP3
yDdb7YsaHUNj4QZbBN3GmxC6BH/qeYueZsQXmyoU5GXg+bXCnpjywSx8Mf/Dixrd
BF+A7uNKUjBu5rQ2sUXQRdY5AK6WKHE+AzMhEmoTvghYU9sEqOPj1UTNbTTbTVGJ
WA54DiDF6yYoGIGSmxWlfapJv4klHPaEEJo2yJcgJCpPycpxBIFS6vBx3+0iO4E8
3ZODQ/eYFYfwa3g288fTIfwODphNtKT3FJTgpSUv+M8T6ifw4YegwbYGsoEr5dvH
SK7+fHmlxivSOrAIbekD+3yIbdPYytWn258Xd/jYma3X1je2YYg6JrNNqztCV3/L
6h7AsS28aQ8OMOiZPzI7ONCyNKwsaTn1rj1WFNQ6WPU1g7miemkc0WZq0Q8DBSQh
1EuZtUEAoOKPuSgV83hYOBicrMTCf9fzgNtFZjIz2qQnePnjuWVCRH/byk8psrau
1kIlgG7Zw9s3FyZavUUHsxspL++08OP3YSE32EDdcMx/jY6vQkUY5SiFmYkVXu4q
GuF0wPF9FItrwJcZjVxsSZyPY3mRI25eTTbiBtzAIO7c4OLq6raitV6Idm7oipav
O2kOEpZ8fw7allwkPpxO5lrHRJlyQ0HDvfqtnhtbsz3l3jMlXKgi5q2z7/gWPgyR
GGESICC1wUxEkvK67c314au3jedTVPOd+CZu9515rfzT8U3o4VamB62eD2IQYNhB
xYGEv81HzkS7Mq+74EkxU6ciReUab5+j33Eg7QDdBLSfKR7XCYYDTSakQ7gVHhv8
PJuOr5BocLLXrW0TcaJo6MIbioXflKN/vuLrYcCUpICHkZ2ixhF45Y6pCeArUEXS
Atd3aq6KplV77B3BPHpSLXjxME4phLAtGJlKTVJlTJRBbpj8MKNIxAN7dKuXYr1o
t6WCgFvbWq/673IJLLXJSUVXKXjPu2EjvllqZaPcCzt9RQG09vOqyXf3dNzlrY3F
lSuLPj1wgTYGyVwwmgAZP6MFsezly8ZYc8p7A89xYSnxNqNu8dOL+4vx4Gx+jMfd
uAnEenRsUd/Fp86MAlJehc4dN4w9HH5nzdwgFn4KvY5UEBZkhXHlVB8nCevIsdL8
fIUwareSqK0x0pGVkzKwn9owpPCNNs84CEuriLu31JtoXtEe47RPTklFk/vd214C
TLuiL2hDK7VFqqwm9KjWXeocIGQAjLEdLkXIH0Nb8eB7LHqYr55e1LSyk4EbaDsE
aOPcDYav38FBJd1qDa1E5a5BSFgECRZstMQVqsg+jLogleEIB6sji6gMIKMQ79IH
ct0/KuaXwFTvZKpMTJX7grCCzHMmvl/b18vjNvRgP8tM86DwqBRWKk1J3DsGr37y
1dqE5OPaU25I2zQMHSdKwgCdXK1Q5cia3gOqQAnWl9dj8KUkEiMdRnlbgeB0sQax
YqmP5iqRqA+UMPu4/NBixEsY8rLut3ArmMc/YCoF/yccF/0jaJen8zp5izU5F0mm
O8bWN8paR57gztaaNPuo0L9MOmMNfnF22lUar4wYlMbeKosP4Pnv1h35v8Dc/fTn
U9ULG2YBdVBZAQVWB4Tp6/nQGsM3Xjg2aqYBpY5L1mLR6xyNslAcNe5XsZ7V7Mh0
fhLaxp/76ndZsKo1v7JJOYy+i/S/uXnf6quq6XG7/8nKaoaijj5O1WwpLBdckGWV
O5l05GIe7V+rqzSo3vJXQeKmG9+LfaN8xyUNWY0MfvaFubzXSOA42T3GCMe60pnG
qyKqa4S8tCtpzOGOpysPWdQPogjAfu1yQ2RkbXeCjUJ9WGmdeKobo3AjZKP02y8n
9ajPfI/3p47GRFTOkTAbmkuGVFQPE0wvsOPdlz1DplvGcC7ppdNq+LfVW5A6bYpb
8MIOLnpAu/9c2RNoqCLkqlkUMcEpxFvwWK8GO6k7Il3l3XOriyck5mL5qQYqt6rH
xs1sUhqLQoR38f/9P0gGNGve8THncmoNZDHi2V1R8Pg2zqKG5512RPWzQRWHwY1X
atjDUsC1zyEMmvzHA4GilVe0Q118qTk9d0Csq7VEBbH8LVqZYcJHTJhFQzg7oL0B
DYb0RtX9OTfkjjkKu0yZFASCNBljYZB1wHF8gaBKmeooEkiMVPCZSyi8Crz+vAa1
K1Hr3tqRVcquGGovI1cIQZXMhV+VCKWO7ePzLGXsn0LiOM7gl0lFyES8hmMzxsUn
BgjtzVS42ZE+I16SHLyROu93uTBmRxZgyqHs4csdgoUk5ZOMC+XE1h65qp/TPlvD
ZX5H7pz1ad0HBIDqOYYM/sLxj8pPJ9xeuJ0hkKGXJVIXewyvgW7zCeOCCb3L+MsP
AvrtrXpkziGxCdMJLlTua12O5AMyp22RTGsmlpEtNHNrmCHbKcGKqttiBGXfpCwZ
7FBc6R3eM0i/eiOAOSW1ztlQIinxfELJHtV6FDvCVrIasAvWbocNTGovAmNfBP/z
VENyGbXexPBCdrOw6bz4zVElesibr9zN7LP73efk+z7MMKN8kDHqOEmAJsyqRGY5
NJNspuyCOB2TPgqIzIiC1H7cLfYq/C5/VkGVDNGVPwrrrvrNRSQkMoL6/AVxLqWX
LJ3AEmf6yhDi155+r5gUorHXnIHHbumd945hgkUYE/89K2rW8Zwk9NoPGGlSVOd8
5DtBBe7BDuTaRJczTvL1x9DLND0gwo/JNTGxYdqlW847LUCzuhfhQaAXF/OmJ2DA
dq6skUySqioEsIPCC6XWQfrnkmCGRJHp+sEFg7EAGHW1EkqWMg19j51VsI4Ow1wa
04E20DqCgSWbSCMgArvWDrh8OGYObcIh6p4b4jR2KKln69bf26/NOI1zpDbZbO1Z
CHAFNHkYUtCM6mPhT+Lfn21DSZPA9lQ2CRKYePVS6dhURJBMXdsLtfNbBl0AxEsx
s9PHGp8MREF8+uPrvKToV+a88nqQHIeEgOoSXDzvbnaR0i3Q95FgSlUyXKp7umOi
gkSOQD44ltdd+YiMLyGjKjdPc9UNrZ4V8uIJrMgv0wlZB393sv8udEi4MmYLK/d8
c6gP9zvgLNso8KZhMg0M1F0FCypP43h+fd8sDM1Quzi2NEwDHKT1MLGS4wWzKPFT
Qy5eJqLG5wn8lj0/uuiRhvG4mHPL0C+P2aU4r4tV3ja+Wo7zBoYrcacIlddf7wIu
ECIZGYXY9Egx0k9AwCn4UhpRHmyBU8sUxjJGT5VcKd2TJRsOgiOqzTH5GBU91xSB
MrZofO0wODkAuJzkFV1x0/4Yxc2aQcOlsqLpwj4/zcRkTiRW0OJu+i+/1vl0RdMG
j+uh3m0o8l5zsYFj3n8CHb5oJEAAMRad+PnqTOO5RjnQ5I8aZbRjp9U9hhwzTK3e
ZSn7rJHt/o9DyEgiNmM9Dxa6jMcrSaxl/qenTS1PoJMGOhSLJm9R5fB8HrUCRWDb
XBKWvpMk8p25PG271E7+giIYN8OHEnLikt/zCxJkAtjIeTfu51cQ0N5G9rVosKww
cktqL8W0yJ5L0Al+5RnrMfepgBcO4cgMdKGf/YvZnlNQ7+rsnEJiL8kX4YDHD/wx
oUJ2Lk//4GwrTeS1dbf6vBuuhFaYJpuPlDf/QGKIr0XQJMevp1Z+RTV74/m/d8jD
c5jYrbqbRhv0wQ2RlrtODNEwDjeikzSyGTUwnaB6Y5jAILk+BQLElsosGMOiUgZb
ofOGglRwQwrlNYAYkp6x/LJVlOnwd6BY/Ijd0OK5wZMQw6OeMH/XWrIyVdgfIknz
0CGbsu8GPf0ZV3+ihmcOQ9aLuzIjLV6Cs8NhizD32gzvx7aJfnRGpUz6RN/J5KKL
Avs5T7b5sP1dZ4Negt3LI+yRSuon/VcnfKbkbhPd2YXUTzpfKemOtJCs4bAdtW8d
Zl5PeoRbBn0/ARcAvQCx40YmOPl/mgT933QmUdu/Q29N/UZv6ZzbyFu9FJ+aIZJ1
fwtSS0LfKHTYuodYBBXWDgnwAw1PDetdiknDhdUDF48Z2kLUrQe9zJLqka30lDFR
EnraBdLtC37cXDrkaFA9zSLG7bE+cfM8qGoXMSoHtFHDui8pnqPHPdMpK3SWbkRM
bbXLnh1Bn9dVm7EbgJ2gfHr6UfwQNHcrmohC/IX9b1CO0udTe47eC8uWIsUwabFt
nVQI8/BGkDsnvmgVma/AHfa2RmIvWkbXSd5fwkCqfcFSUERQtuZ+LlHBilj9/dll
AAAdkCNRTUJ7q3nSX7YmD0+EL0tY/9dsSWmFfM/zUI3WV+6ewstpJQqgzq0GyLzC
jVnpHkpBvFb8iGpxX4d5nSWCSJFSJXVC0QLcGfJBVbGKpgz2GG3RKRB1UdD4nhkO
qKvL73C0Ya0WVV6z8GuJchtXlvOArtFqexrlJfajDFtIXuZgIlRYb97Mma3ON6Db
njGNtqiY7Bh6ggdx/qTv6LsLCRk+SWnVMaczJAEs8ObtvRzDNmdk70q2ED2LY2Jh
YwnPlVhzGq87P2It4mwX8mn7ICO1obkn1O6uBCgmqSqu9sPPQ7qFMWTNdK02GD2u
T+jopzE88YI7wq9oON4qdv0j3eF0GG2cwbP443XDqj4HAUSsNSD6K5F8O2vrYj8U
QvF5zwRwgcKJ/WQKBz9LkaNrhWMmaGYM97ewLAmfEXo/4p6HWWr0hORaYZ5fNotz
dJSkiX1c+jZcXp1PalxO57x3Yw2+M0cRKSjUTwr13zLFnj+49q89ATLnuGxxKZ3a
rAQCYtuUEMXYvzweVZN+lox/C1TU9SJUBUGdQOCXV6z0fjZHO73Q8iTRLVWzwZ90
yvCOKQqOs5rBZ3Rh+0q52neVBN1KBA8br245eoHHVcnAJd7wRMQRN3Row954CgEE
NO7iwBjr1nxQ1KsaHhHsNS0vvPQaR3TOVBz3upTzVMfa9ITHvTzf14J7baOnTk1a
GnvesDOXVTYl3NuicSTleCtv2NxFxrR7l/+VDse2qoZNbEeBEvDXFbDCsKnRP0VQ
n2/OFSbZmcMNhPQoTEb8r6gCXw+Xc1pEVWAgclPNHAbAUgmNPCvlUFEdFAfjWDTR
P07jTdK/wu5AgCPATADP5iWLYBSLb1Jmunyci8mcTSGPX0G59AHzbN8azBQZztLb
S8SP0uA34ghV2QCvROF8mQco3geEdgfxlhgfSGpLv9paaBz5J4cUs+xSCqJGebO0
azlk0L71MffFRyG/GdbVIQGAHm5yIXNbv7qrsheH316Bfy2/miSjpWPy5sbZAyOu
t1koOo60G3fldV7N0mYO9t8guo5sf6puxHOyeLR7qj2yWLZ1WxVI/HP9RUlLMW96
w/xxb5QPtyuyf5r1WCKuR4DuINfFsWw3U+yp+vBouMKuVnSEBz0USmPPLSn0m1FZ
l5IilA2bKvBO4d2XVlfp1vKOdhlGSttkKgc0AJOvvFGjlmGdwohP18FLkBSjGa6Z
QcGl4OwKiyoUz04oDS0XT4e3op1j1Zk719N5d6gYVByodH/EaYSFpuidU5N4oH0C
yPQRv9S+KLeQD6UtPig2Ahb8Wgd1K486Yxw9V3iV4mXY95TNVvk2KGn9V+KXK/J0
9JVM08Izo4v7QIoNcdQqZ99tIQHEaSUOfV9ZT2PlxIgfxHE86bCJn8FN7oikuVeb
iHTtR8Xv/gol8Kjr20wgCl+VzaGGkiKzHS1bXVLoX+RJ7xWYLcuJ2T/PtWiFw96v
jzQI9zw4cAM6irKrB+c00qbd3/NYzSfIGKaH+HUpPH/8vdVr/dEWL7PblSZycQG4
28Bba4j4KbyfuuO/dlcD9Eurln71XrFtYTPF4vMwqCFfUFt2KyPi2cb6SwMjsn+d
3Rk9gsq96umHYT1LVCBLlpvLJ8DWPb9tZnYVbu1PVAC1ogxOxFxt8PwdVoooFMf9
sDzhxnRy64UjSO3O2Nv3ka6fA/wTg3V+J1RMqhU0mIBgsyBfDkcFNwZIjeQk0avr
Wyfr7a+/HySjjyUhmoZDFvrpyxkgfqdtL6hK4CRFGUZt76KFX9NXIYq7z8DUliZ8
K/tMawYd8bMMYh6nmVt/HI9Fiat0M631XxTmMK3MObdY6LpxxOgloGs61dKVsAhZ
U5fpjci/6+dTleQn07xIeS0SjX0k5dAJSBoVnfq0RVunQrU6bxDIfxWMyVMwE82O
sgsHWqYCOGlYxjfzqoD0Un6eLoLwUPeYv3xtlnOpM/VBuxiqer/4IWZJ4VlzlMml
gnBntauj2b2auj7INQomVSJ5B8HvKjV6RtCHZa7M0JucJYJpIQ1/hQZUd/2QKOvE
VR+52KEDsQMT3F0HYi2ERiUX/rFPZ81WOFoIvu5t0ZGhT82k1h1pPNKzwRjCe+4L
PoIHFrq4VcGRbDE7+np4rYpZ5zWlLQFpPC5v4V3AY5t5ANv1a49evnA1scL04GRL
id1StBkA91iSvXGE8mEfHSTzmpjRK1L8D2V8wfoV4d77H4pUFEgiXnEtxrSfm7n4
ioB6fCRol0sd6c8Y/yoE1M5azmX2tmBRvhkxPrp534ikV4LCHA8yohPG41W3ljVT
taHNsYVYp/ro8uKpphSXLhWMAfArokMOIfboCnUhduw80LzkBM9oLNo7a77izYn8
sxYG9mPIZTGijg4rFJ5hTXAmq+xCv80z3PKLEA/5+Q6ogozYqyT6dl4RUnqb/f3o
79EOGj7r21SL2TFbDHEbbAWNHmicWBV+Wiwspng3bpN8S9KYuVCESm6ejxtD7mGe
GqvbNUkS/21c5Fi6nOvAyhCyecgoBelVTWRrt9RtCjFnmW3WIrTsbvSVfSvTotHP
XmBPtQ/0jKQHkLh/aOqfo0zNTUbdnySGf4b2+VsJwQ8dZPAQIDqQeJ+4nLGzDZf+
q7ni4OEpgoaJ1jZVs5WslIsPbljKWyGbOW7ycD0/9UP9Vo8FMAu2EL6x4Y+F8wzk
T8DngwwGUssC4KPrG7GoBxOevdhLRwt0RY0PPTvoYJnnQK7EVGAuF3iVoPAkL3Zk
WwxiDxg5rTvX+875E0ylD+hD1e9p11X400/Ibs2a/qQ+EdH9p3WFy5+SHXGJne8e
fwwNM3FLJs+9MXXk++R9qVLolL1sawC4CbcTx4YsnlysrAKYNSscbsQCAEtHN6Xs
nSmfuO8YYtdsjJQ5zaTM/oMyWmF01pFzwQeF8ivQ/Nc4Od15b242byFOm1o8X+Xh
9kUU/luIbYaZQY+ia7xxSGzt7Rv+JHIQ7rJjCWGRrTUXmEPzucFP3EVg8CxrektI
hdRxON26BC3DRjs8AoDJy/KXuhrCoJsfQbVacY9Us0gmYHDXrSHf+K/53TgkONFk
lNRQFLvormcWY+NO47WS8DyWSKAvO4M1m/XIu1Oy1f96wbymQQzPd2moESoW+KVO
yvQEbZ8wWeMta9FVCk83jhK8o4Aum8b8l9uKu2P0a68QzLtYR9LAWI7gg/5T0Uws
TtPW3GIVaS13d6Z4NRr35wL8C39Zsjp2BYrdIvSaPmv1mm8uqctWJIb0zpflVCax
HI7Obvn7WQ1QW1YREpL9BlGCymzFqV6UGC7qZP8l0IoCFTT2WBQZJMwSprR9w+9r
I9Mdn/M1xlswEgniS1zzjunAT2RnstSXoys5qsC2wmoIy5AzZc2OispSWYnhgZ2H
OQdpF8EnmEvpon1AygDKBsmCzClZmX16i/TBOXx3RbsJ3ifAAIjG9JKtatdeXKDc
r22lytE5dUoPCi+gl3ddBSVRY5TKTNV+05tSpFdriuhiM82pkjnhl8V+USLvq1L8
+8rq/Op1jrYdylSBUxML8L24wxuVGfbvK3fIde1pqT8wGuFGoj5Xod/BSMyK9Jly
sKwHYUbXT+qIWJVBqt1lISSLL20VqoQ+0/qdUayjSAcpNEJxgTEDWmZORcvhXPRN
ju9yZ1EUx3rH8yMvjGkRftILC1i0HqrsLQg2WuUHdPP6mCHR/FOCMwU652KSWfs/
dGH/9A+Zz94vnCFJGv6pFFAh0Ui6EZpLPRdlLS1U0HlAQCyhwxE65BT0Jbs+xiO+
5oXtLj3dHrh9Y6fA+Mf33y96psjqrH7xTEK+orjYjTQ/BGO8Bi609fh3Ztb2jJin
2D/MyoZZnasSHFLw2KIc3F5TJTtxHO67l/GWDEhlGr0GPaYrnlp7PimGSui7nkqs
EXO66fZxW4GI8koXfOwo/Ng2FUiKtvZLd8Xi0jJgjOduZ0ZMBQTzodIIvfsQpXQL
omt2n7bNpRRHT+kMI81DknOawuQPMGM106mqoceGzEx+9sFBg/fLrBekT7gv2iIV
wCQeu7+j4IfNpX50sIuxzF24MGluV7Kf8iqlOHQ8S1InArrz8V4EaeIX/Sdz7ED7
Z57GwEGUgEoYXXoZeem8Df/OoC5HZGrJMo4na4dwmSeKImXOdSHzt0OpLvQhf9rx
OKXGApE0vcQQxWDtZtnyg1WQNHLw5CUOTyDEtyhmh1604MT5FdFzjTEfJCtG1igB
keZoVgeinccjYX/WiNqzBOWVy6+wL8qyacVzYJMj81qOJtFaZ+I5P8D8znJ0dIAl
XwTQHcI4HbE81sObKDC9urmCmbpo9C/zGKrI09Cp+Kik9OjUzuG2pXxtBbGOJZmR
/tTXJ06RgebL8nvrWD5mV9dhIupH6noIPIYA9MNbRAKObSae4NYMgwuo4Uz53XCR
BH3gGETvk7N76VsodPmHCEhDsiqyW1kf6B5YWXPzuADCnhGg8mMkm/OEFtcydNk7
EIwcnXTGk0Gh9NKijx97+ETQy+isBBQvOTjDi7+B7yhTpTPCRIQStUUlAaxfCTSv
eY20om08DU6nDQhBo5p1bb8mIH83KsND/K5Q2YIc79e0LN8NUPOtX1UJ0Hym6gs5
Rv4XEqMerBq+vi4o944ycYi7JFPFgHdhJYH0BCT24Ft9snsEpUs4j5v0oIxQNL3L
XDP5NkJQ3ueOf1jaDfHKDVCBWzeNSTHefmjKzD9bz7bsR92wfH4GAz4LoSyrhB6E
YGyy9CDeR4Bhd1O1IxEMobsG8/Ee5S8hNZPuDt1/ssB0xeljKfKJF0WkYFYIAKhv
+sUFCc0u6G3gtO2fd/FkFAJpW4eLRGnvyZwtO4nk9lhjyypBboJx1zKKK2x1xQa+
MNsYqZIdx82R9O1EMNxmfKlxuhK2aLVgGumXL/O8BbuAzzSG68KtJS+4P+KmVD1s
lm0eRX6nABNHsMI9j/EhcYbzEXF9qgPRtSg0wyurxCPcVdzb/t8JTA9dhx0Tnj0e
i68n6FrA15UrbdsMKaFO2FB29tfMs7k0liWXCAjou/nH+nyJxotg2wPBQO07EGQN
n0NPJnTdn1ERgHtkxmmzDVTwYp1QMY4JVf9FZQ3/shrKv7VCzCJJVqibsqRfV8cV
k7Y7igqRf3Nn3LQPoFMR3NhFtnxA8DYaOGz8mDUhWxNGRWqtCUjjc92mFzi7huJC
qRS59IzK4DA/+2JGj7XyV/lEzgzDSq5JALEnl991XWk8HZcsVHophyJK0qXkaSu8
Nkh+BQbtxjG8BzstAM9Vasohi7DABZob7e1W7gGp6enCpbe6s5fJNeVPWp2mlr5V
9cxr3UDwGvo5WciymTlKXfpNTOnGa7Y3e8I2NvvQrsfJUsGnL+IeJlAY6OZz/KH1
GiQpJwjS+ad23O/+xx2Ayl3/YaecMaz3mFKvDZtUv0oJwdwB+TrnUZ+lq/EN7m+W
lMRFou7jpxpNAvT/qz3jE0Pc9IvZF+QCq7Idv1MLtHCtLNXtKbSasun6x8PhDplb
1YhTRN2FNvpRqhLTIKWcFiBCbJO0xDtLnWS78fm/SbQQ9A0sswWytz95Rc5cdvXh
9koeFZB9SAWcnb0ASWdD5YTle7CrgN4NelqBe5q6vhI6n5bxpKp4a9j0wEiTgh4x
EE3HU4/3LzUpjNFznL4Z+6J4kt4GzB66BgXXSUbvmP2zSqb+i3Cfa1YGDC6Om0lk
p3uNGRp3DCbzquwMcKboYGM4haWKiX6ZgmJIzQaJZp9weF4NcVG9zmG28PaLCfbV
jw3HqjUiqO3bLFxglXlRZVOd+1EJ2iWjAykuKJnml5hvYgLO1DDO1J/aj0Cwn+WS
Lxhz0eEKJOz5p8RbPhYY2Jyk7MnaUGMMYdEW2PYxEg4R9zH/D9Vyeryo4i9lq+yw
3U7vCR4VY4tTKY+GFageJioozK+jZb1Qj8Eftt/+Z9LnJhOG/G5GMS+dh+qp69X4
EDMasnVmh8Qbfz0mDHBshoysBzsccyOVpWuCwIeD8GNcnVQ75PkCPZYrFVT0JE/k
MgmRQ4fGSMv8lix5ZQTDNcRH24q8PBJeg1ca82hYUkBDOUSWyXnaxxgYSrTlYi2H
HGh9CuunTcvsV9zMLWcvD/pifIFeLjA7pPh1Ny9F20k3jY+SCL8UuRu6CNjlTnvU
4v2VB3clxclyr07sZm07dFZFBI+Q7YWTLZHdVX9bXPNLt53+CFpaFjXxv7dnJYrM
HDsssfbwp+VGDTS9sL/AgHbFQGhvzv90FeDJxz9a2+iq91goIObe8qJ4VBDwDLxI
ywVHmd6h2Ij4V0dCyO5MZEjyUEuiJqNO7TlXuTlyEtqeQ8xvKaqTazIODV5lgfyX
184oO6cdwaRKvuvQ20OK6AlhYwgfX9cJkBk50PcwuNuJW4ttBv9A7xKEQko4qoZ4
DRVYbkUqlwbdnBkgmNk6fzjOyw4WXl5GBm6WufWvrlf40Z+hP5hX1USHOZmhv2Ys
MqeTl3nGjGe4cYyPwT0a4vdGm3KHdOmUPkVyP3SSdpVoGv32Y/WyXIThV728DkpM
zQU33YmBCTFAxsQk3mOY+V6VqrCzRIzc/fUcZpopB+3326AFVdzVvQ+j+BSerNT2
SufM419C2cCkjFLKvXlJ8aUucWNt5pXxMOLjYV8N0Ajs7ZWMfr7zgd5Kci32gMvM
+WBqcE0PDKEI5yOx9MOrx/5A8nqyPusGCRAluApefB8cra5c8F+X+pxcx4UzVBFq
yyD9gkAUcHLlsSL4lAsQe+TEXkm6xd399IrM6f6EQxPdVmhBsgIDOfYR4yUgMoPT
7YiQbHk30MoWJGO2XPi2igPwhFyXRiCPibQnU7iGReAUNby/Tgt/A0JXjoFeM7Rb
sBKiwWrH2MXTn5cvzVjkFUNwFxYHMAJ4i9ZOJOOiGUF169xp6C5c9Ws5Gikpy6sa
lhAbLltsVZtCE9Em8JxBvgvvHU288FDgCHl84oORJ0vtife1IwjTze0tYB7EI4DF
rHL5Z40W19nt1UZ2NLefOGZDU//PSObdr0dfYMguDbVbOQ3Ewneql+6jxYlgHq92
qZDYnZPcPEdogUI0HdKcPVgGYzJ1+IiZxttD+ED0Cb7+/oIfUJfYWHsHqpvUjSWp
GpJd9xfsx9AxEQjbcL9F2DvhHjLK12ubBHWrXbyRybVn+z9snzCPbCz85XqVErbg
GYrGXaLe9MDIu160suCAtdtCDT9tbN+u0GELj94QWQ6ezlsl0OUFvHfCEXkIGOG2
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10128 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
/GMbQK29Y+AAYqzOrLs1adJXUyNzEKX18xw111ld7mUZWMUdPGS39zmQM7G1RKq0
22ZVOx6Hx2AxnYRsAMu01eiqz7k/94ewuafYUyTU6lZ52yaqwf/Vn1DVp5H/+2vf
4baviWfDyB9l65lbR7tyR97+iEQzsJb0FRMZniU8pd3zkxKYApigrnf6K9Z0jOOV
uRNm7ePQOrcvofGZG7pXR5tiiFDMgdoBUTU7Kh7BDnCJKprza8bLBTzFCtzWxa7v
nWZi3ZMJah9bk0zUgA+umkI44zPG/rAZtcM0gE1H2LjpPtNx7e5nqGOODxphbEK0
Qo9oi69yf677ccU3l8AvvnynVrj77tXGlLvgo85IZgabMfTAqdczkHcE/aW7Gvgf
Fz0/KY17F/f+JIAQPRI7dNy51fpmJOMcZRIx4TfgwAR8ROhsJWoOBPsXrY/I/drw
fIyoEgys+h+DeFWGYqBzqogBcA7kQje0KeesGi6H3FLayo32tQ4y1JHe34aWZBvP
uF8XTXTQWrQSPFUB71wMVbAjvMElV4ROWFjuJrGFq8jOyf8ClbX3UEuUaUN3Z134
2Uqu8RGGMrKwve4TAiHR0CzfTPkMuqe7WMdeRiUMuBPNkLwAac5/26PRI8hKBhzz
Nr1aIc+dTZYVVixlaUd/5oNsWeombytfk31gTlcXj6I5e1vYJFUNc+ufMYkJA8g6
3kHpp46UjHG6fGVSlZLNVP/pZrDEI+HmACigJeOlITAp/UWwXgkE/sknFLUdoUwR
r+gnE0rqWbgsL1BN45mDsNaawJ5yprifenvRzWCPjlYI2TGujea6i0oUETIUONWm
P6MJmR7uO+pxrL5elPgt3CWlV5evT/GvR57LQiXHRERYWc+/0sXnovn4hMcg5pU7
Y37cg0gQxXDf9k/cq5x/jpKz47JINw551aYF3rbCo8cVMnQjqqfk5HjJ3/YuCUp9
5sl62tu9kT5J9BQKHqzCktHsE/gaXX+QdijHssbhkeeLvPfX9reLE+IGm/xfpvcR
JYgZEpGoT4kxOpLZcErdZi8iwqOtq7yX84t/tApGdQ/u7bRDMNdIwP4k6oF+DhuM
vXX0drDhR1EjrFn+xiY/TcEvfegExTao/s3KUFIySRLMlR1U4fZ63XBsLuaHu7uw
EGMdo2sKB3Rx6ks07IXP1/hRskw+zUglSjJpFj9DkcAvUIQLjPjwhbEL1Oiclh4a
kAYhuZCt0UaY1lZTEY0GQEO5oLJ4DcR7E23Fx8rkHqQq3s507XgpZBk8rqW5avDz
MJxsxjPW0QH90gZxYBQFcmU2ifOACSVJ6you9weRQDEvmrn1fM7NPW9RP1UM1/3g
X25op1HH10K/RpiRYG1/J6CML4L9HNmIUUEPaF0jnLwGb0RojpvWRg1WHpGzW7I8
1Xgw6Esa9SiEzhtyzfMNDBsbPnfPTpoH2aYVajRTOsUzT/rDeBX7eXdiWosaZ7Up
MSfXcJIAxGp00CX1wzNIaYSD0e5chvx7B5EHbPdm+kdHYsyvpajyrwLoPHhCs8GV
mc6KfgSjibcq+0Y1K6Ry1UeRZpbxE96x0U9LdHjCop4yfIE/ho9Sy6i3inidIE0Y
j+4cbe5+ajckKgLqkVGAQnrGTK1J8Y0+GlSmk/Zm8d2R93l8kkufclQjdLKq/Hy/
g6oryf34i2c9QTuI0XhWsG128am8TwQvjIfYOAGASst+QnQjij/+mNYkfiW8o5kO
Rot25U5O0DjIHSGN/IMGhzjeTbHd7v2BdWRzbu5n7o77freoGHgeQSreFoJQonUi
6mQQ85S1rQLGIV9887lJ3HAi+YaWROkYTLXK/ZebEHG0sVcpuLCUMJ9mfn5xQYRN
/jAEUB72eDj3YQDC0kWWQe76ker7ePVZ1+oVPIQMjI+rVwURuOt9tCWwuxG/h97h
j9HatkbQtwl13H8lYMLzfrc1Ieo/pdwRXMaAYtTkFTeexZwt9dOua1eWuATrla6I
+zsE52sxQi7C5d1tc2H8WarhVUqkat5EIV1b+w1KKjuOX6tzKx5hze31HqqkQErU
VqHR3MJNa1bBmHVKOqpLs0EUFy8ZNKflbES+BHLS9gXby89PFlaUGwRb0tAAs7pa
zUUW9jY57cpUTGBKzU/ahdDzyFTyn19HmlOSWrt1SCBhiIa7WZpqwmA7D2fIiQkG
CZDWeP/SdVntBQZ11NpHuLGGUSVBUbn9nMHWEhJrnaC3nuHslyHaQ20G8oAU0abx
/q+EExXVAcRnHFKo/oLa6KPRue+xKdEYI9AzVbdMo3/B02uzNcIwIb0n7VtvSPKI
4IoJtjdD134kArzpEt2eX4tmPv/NcaMsmH6LieENYEJL3V29etsiXWYsnzCBLeTR
DJ68ZRwdbqb8J4mBEvs6DH4qw8LEBlAqK4wx30D/KnljOJQ2UYPTX4cxBpG+D6C1
b2FWo/rqO5f+8z515/P4MR/kS3WXSjhT5suzlYJei1oaDPUWHClOPD43ywdNX1gh
XlCxMQDA70lnTXa+G28hdV/fw9vCWyIwD4e3RCub+8jby/6o/csQrHwR0jSz4wg7
d9wAOCYwbFy/03O3wJlM0/tfW+YrLQfO1VUqoycnjY7nI8ZgccrZzzruJuf7gnSW
hIMgXLRQE9NXMjsfUIVGMSf/UVxeyWWJECeEkD1hyG6JfRRUXnusHUKscnugOu+N
OlghPPjCH8OoAu8opWpyMNlA/OpYZv5E3xa1EovlQASut5UOf7sIpSZF3VzkSEWr
vaIP8dA34Pdy25o55xXM2TCukLXUOTKNm1BdryFNx1Tqs/YiJxNoS9Vek5D3b0Sg
4KpKiNAg7kLGEaEQ//rKq1EfyM+J71OgKqnXgRFg0tsUtnpmnAMbJq4GrrPPqyUR
PONfNBQUETJkPzcxFGUGOcr7I/9cDNTl5cfkihlLp8q8yhBVcNmSkGaZJgqlG8cA
dGy5hjLv+vyByaMbAR3M8fajcQnPbOoCijURiQ6dt7gLch9SdSiSzizbPOWCxDF9
WmIkg6hlQG3yfe94wWYC9Sb/qh1cZMhPZ5pToqO/KDRVFRgCbC5B4unL3zkNm/pg
ENIpuEX9xtUvcQX8EI/ODMrHMWmIX6dPChrnBmOilb/6T5+u+49AWueXBvPxAXJw
AiDot/u+p8jhpfZBY4HVLBihaHznNROq5P9OUpgX/44J4mFqXGiz2uwBC4VNH65a
k994LNCQhqQ8ZNtCPdrjwRc4asl7AL/wpWNH9I6NCOQRxpzDEtklSffDXxqC+UQJ
ONsaowF7Lg00oN3vNU8Ic0iEDTYgK26FpY4UcH9/hwMzE8lEqCJz9N7193Z+iKvw
J8vc5fUSK/LBlShIhqSCr0+I71tD+5lSNjQlM4nHoRkaO7rGIy0TKOGkPMuNRG4c
uGVoti86B0zM2bH7sa3qauypRbXMP09mm+g23f+DKGYQ5auft/JkXxnE6kliKoon
OnkMm87Gp9AKQOGcPLwPw2VvbILIlsRiEhYUO78hFSHsZTUmaqSO2CKfaEwNxJhP
SEKewu8j5/MSIII/13YPvXfZuOj7+X70F3GWzPb1AWvyQL/if7kfaCZYQs1FHctt
RKzVyrhO9IbeAc2VXdGO5gq1r7NBx3UgyGvskSRyJjppHOtACQ6w8ULtO6LqbDuJ
ZsAaKUDl2TNID2BIQftXzMgjFoE0We3L17xHfDC452I5z57xdO21VAGTPJ2wuCsA
C+INOf7hwE6Ab8E7SGEctnCd4LomOjpnw/g8EuvKNdfUm4mbzkG9O/FLti9Krzrp
M4CtUQQiGDuQeN0M3Isz7s76sYzZACq8T3ZsqIT1pmzrUIzxhPg+ClFq3CRlmq0U
SBVSMISeP+VshH65pdf0w2sDu+DKlslX4e/LQxfHbJ7v+XsJSDy+wtQOszveRbQ8
Rg+IgmGomPqdY3jjAatEa4zxzxyyW5nseiiHLDTQ2WZ/mxOP/trw64+mePZIxN6F
egeWGi8fCjgCIYZ5B36NIBs0W8lp03aQJlYUf79bC9sEQpF6qBHrbMbPrAQUauWL
+dNy+7R4+TJsiTHBQJFjkSvqknhn36QGlAUrY2JwDSX+8yaoHaJ7vaZl5jDXthIh
fGZbgmPt4eBbPjf029vVwjxwuu+zolznhgG/9EKp5JaBVfP9jHyiN5DAq3fbcsw4
cfWWv+WbAtfCs1/5UZvK3rMRMtz71i0ZA8kP7KAusgJ0pKdoQuaHbcSv+21e7dgd
wB8h7hlRh80rKxFw4XvcUWt3VEDUOPXxWwYcUR/ss2+oyaHYx58VsBF679Y45m88
IKz2bAY+sTmlDRMKOGbjMBb0DqgB5JegOQptJoZM2WzCVMiq2y5wl9CyHvY7t+hz
Qz6IA1EuhKOlFb6huXTjEp7dYXJD9DwIX2rEB5LJtT7pMmu7RHcIqtYPGLFMtOJE
mEWm3YEAiFhCSNvq7wsmdmhIJTb2rFnAGT2Vr3C++poA33/xb/Saa56jkdQlb5Fx
nZonWjE4f4RMoLPptnWswRrfp7nAAbjv7lZp+2JPu+R3ah/+zKpKWJkYlKCOoTOy
Oc/3MwGrov1JOPJKFwMB+rmSX+wEj7aqvn3ztJ+bB8JnMMfqRjDPNZjSBpiSb4U3
bi4T2BstDDAXlxiTmLDO2fqfu8yB1unUG97PKaryJ+uFfFhupoJRDs4a+1j/umGK
SARU6oOc94KcBH7uOc/8nECpA9p2xbecr90M68HmcTitkIVeUT+vZEwoHvaF6UbC
Z4NZ4VCAmQ041bWxSB8tW/h6n7hKEM+8msts59nSv9ZJgNzwKsuVMJT68wVwbGM1
KXNTN+zacbhL2RYqLIz5sgeK30Oaej3whI2ecKfcYTHDbauNiBhzfCTVjAxNMHFx
SXgFBGaygtTpZfeILtaPFMfXkM9iVnhCLyPc8LD5nk775z6SYVAKIwffW6IWAYR0
iDMbmvADuPVBfuAsig07MKYnxwoVD3k21EbgvpAdMowZUqrkGNSQ8lhJicTicIkL
AqefPNtPSA2SNVf/JNQeD3yDdziXuvczDPm7gmVFAiSlg07gpJhSHU/TZbfSviIr
4rkjBfc3Pk/X9cWcD0UuAhzLdHp7O0GmtFQJjfybXMa8d9hqcTRM15T+7GUcfsNV
6d6JlesGo0HE2fi3XF3yx5PHg9sXsFAfquL5YaTsg4b+lrSaVuuAMf2E0ajNGxeT
GW20ZSPjor5Iv2cJXLU4eNrjlvM7h4QkmAObApfcMKnKh6z/rmUe8R2H4Stdh5Kv
BUglFneeQl7Z4c4TcSK5qAaC3uBtG/E2ZjZF0wjTNqAi0USctZnumG8qdXgEXm60
M3tFvX+BmGxYNueorUwHYBvCy4lIQJKuNx4xhpj0iy6rDnNVkwVrB1Ni3kPZn21w
DB6vodDVrSVBHMaaXMUGa2DAFtPMvDe37xP6I2on8cwgfmZGEqYhd9Hv7DAMju6B
9/AZC+enyjBvsJa0AaI4sfi9rup6HE29Y6W1yFWhbe9375FGhbrakVKCLhA5LGF1
1djdCB+Y4BGcXGcODowzheLC5kRR5+NiHAcufCRdZp5AMRDtKRzTqxYKQ5PHbZha
6bzIAXoVsxFV6j2Pj5OvHV++ZRQrJV0EGaiTCgxKiFBQ9DJ1smBEdmuUkviZ6hvH
5CUSYLvxal+Yw9VNgDY0nd2d5gL6dH9y8ju74F2pJYh4Axn9JrIaxyLs7Bg/wWD9
iUI7+YeLFYATqJD5hhUo2uoDDHiUU7zOJHTfJueh37DbIx+IGYqzTtrEnKoAB2Gj
G/2OzxkjvqXOCMVpLlFkNaKBFec4wXcZf9m9zWzYw++6rDFjzHPjbmqbBnf0JLCj
U24uK8JvFIlxRkhXinWU/omcsZk7mCSZycF2c+oOms8MJxACfzEC/Ewqdy+OxXzQ
bkqqb8veAovh4sBglUI8Se+smcqMvinV/9XHsJzogNLX5yR+cgCXZWh7YuSHuRHd
nVvzakTk5HjBDTMmJ52wpVrQRQ80TTL3U7vob0b9NAfEgrNXVlRZt8fW6BAcGEuH
uWUd63FCjwqpjGWcUsIVGUhPGpwFsdQBqebmamR3LBo5d1Ef+6sklSQkIyoFvkHn
z87fEYo+LSgpfytYaozE5Ktab7/sLZ5yeRiEX2R8Jzlv68bm6Ja+Wa68bwv9iu9S
/v5QzmF80vLhHBRUH80wijIctkBAejQScS/J6ENUhyytJahyKIIbA9Uw1/bMwSBM
6SILK7Pya5GwQdhTbZMXg2MpeHpA96/b1gS9MmKfy2qidLdJ0dRgGS69Pg4ZfiW2
266GnJb8nOK/gMR1a9ePd4wEKYVW7kE9byVMcz3p5jiXb3xfdajUTFOY8BvloGFO
cc/47zQEsFskQ3XMIOCY5wS6Wo3f2SUzU7db4zsQ/J/a/kktH/DNkUXHpv6ejhY+
Qy9hZV86hskyTVz/uytlCGBVuR/wHlY6PGctkHRnxuPciErCKsFRufdmJ/sRmPR/
cAF+FkJCNQV7y2szZ5qlxNj0eFRLDnVETBfRdKlwYCGEPS25vr6PJHjHdjxllxDI
C+d2rbywbeZnjxnP/vA7XL74vgJulAZwAwUiwvTZ2TcJPkZInOHN2UqJ9GmLmunk
QfCYvdTO/gZlKI4zkCDpWhb9fGA+nU4faGq2BYwbNiANHGzOIT2RFEDdxwZP8jhA
+7Q0rgPHP57cLIimGg0L192QEBCRXzTP9k3u9NZ8SU/+55deZGLuZYVg+MxInHXV
qCz56l8n42p1Ot26d/A3Dp3tC9lyTp/ip4SFuheV3VqXb+YiuFNPb5XmGyzbKMmQ
MksDRMbrEF43GnUaVtfz4ML54hI+f7g5AsQFHRTs+vcl0j0G4oPPC5JUkT/8RGLd
qub9Q6M/kVOxqmh5TwDY0oNICmoXFFHBA6ZQbGNKGijzw8yIUqqE3m6C75FpcG1s
CzCCczNMS/vHGN4dYneOlDyfcKG8I+9piZWvs+1g4KxFrRDjpPcOPE1UskXU7Ahz
X1r7j99ebXiJBs70lajVnvZ2/KAB3S4qQAw2RC9+n4CP2izaNKhAA3jL3PG3CeUB
US8yr2uYqCkiDTYeRGgSg7LtD69dCgnfyHj4IisXyr8pNVXb37U5gfhc4tvP5ELo
fYKxL3zz667huGUXukFxFlm+t5bFyt1gZlc6jqptZg7rQfDSUUgmvQ8N8hisPriz
7i4l0dfGGwEuhDsFoT1g9DRD+xnSOXKK1ee+xC2HVHcDbod8q9JKuVtHe8gq0F76
IHabWRAUeDjmbDL1R7nWl2oTe6YUka5SyBW1S4sMrBueQ4YeYg2iGt6lxCIn4cSV
hO1eQl3y+2qyWwt/qwLl+hjySdQHBdA7rEiWmzVc3J1F9cV/ol4QA/g1w2zY8uls
YiaE+j9F8iLWHkih91ij7bhLMK8rWaXukWfkWUnnbYTNSefpETGiYGgQWnZfAlH5
1ijxKnSRDkT7CA2KNOZhKbWp+I899h6r/TVyWNzFxzOJqkccxTkj44WcoOpeG1/J
+gI3TCFhhIXhDk8laWNEG3wTY9KFo1kQWQ62kAyKh+Mp0AxX58ZjXg8ay5gdqUKd
CrNxVjbcMZBifR0tqLd8exulkdI1bwjo2FKdgFpCKwELl0P9OEmAC4XVUirMYO3a
bXiDDytDWKqVqpB+tQzo3CLmUVRvxUOi+a0h5RdShY0Fk89ZTVuhBNz8CTRV3vSC
jvd29as2Gw3feFXOY2RCRWIJw2L/FF7nbyX1BvlPY6uBbVNUuGWG8lcRsdzSxt0u
QbRnhevS5Xhbkh+eHI94K4lCl1nAbrkXmTk9QCZlGjwNdzzskZ4w5PmyraeAcnY4
Dg1O93yVNb8JFwzZVEmBpgCBADKrZnfhzSKBffGJHGWmMUkRz9eRrril7dWgdR8O
+6wzYglSk7xGfV7f7ZObM/hzzWuNSOmzXLDTLwF/WQimclQLePMOBu25Cb6Kwve0
R10POlATHKNaxnXL7sO9rR1Jw5HWkCYT7sAC5lSsaxpEdjjYK6M9zR8mxAsiW0V8
a+0CeU0OeoTeQDODENCnnLFwVAN+US0QFVxK61PCSPe3JSkZ9zLLgzfRFUdkJTfj
zdDIXVbCK63/MN0kp9DGz0nGJsDiK6skwsjyHw9LD4HySDAAYHb7uKV+ioEbuRow
L2rFNtL5SbDTzLh8K7iSmwdwK/aF8w8NShTKIdX9mVMTL6FzyLaRXMp6zUe7FCTx
A/q702OoRUFPD1xl7oyJ0BHp7iujVOB4XjVPv84KVVce3Io8LiAJOtp93A7X41Kr
u+P0WxBlhiuGny+mKdV/G2JBLu4DqLJNpgwNjpjPn0cOCpmlglYxTnpk9WamZXSA
+aVRWg+bexnRvVlhtDPLtFkqGNd8yobFITEqI+eoPPBJs0nKghKlVFNLNwr52Jdq
TxGXpotk81PMusqW8oVMfi8HTIvmtVMJ0PhxCblB0wxBdPer2ynghd4CzPkZnTMz
+a7I5s4YyeKa9f3Rz7m5FAaaVJCOpoUulhdiwVGEL2c0secI5Ky/X4ny5q3X++4S
nbmrRqsTzpRGi+5KR0DMTZlgHRvJh/mPyoNp8xJVzOKL841weUYlGBRjWTBs9Ylq
x5eNxLvCRDb1OiHFMsT1c9AAb3/8yrA5DXkLM2C1fyjDc8lqJRyaFAF9YPlY0fMQ
P0EkZNzEG3e1+Q5bblKLQ77m2fStcGs/Zj90V0gYShM7XclNIu/nCVrbKmZ50bO/
aZYGm2Wf3SP+XX5CMvVhMdPaVFSIX14VyFI2byiOf684j8GflTeD9mnBCdyQduwi
ghcacFNT/EM/7WixmYYf5khIFYMPs7BYuim0KT+3X4dLNXUhSjd8UkKqk39/ZjSu
PNoZk6mOpYNpJB4HUZMNY3+wg0XVaqGHATyuBpO7BJdp+GvCktel0/gaRA3yeMFe
Pj6B+ndXzrEKdjuhUv+o9e4ygvJhX+gh1ZupRKpWIJYvpZvEVwO7/fUpkt+Emswn
yAfWFLaSeQ23DZCBpruBNXv74O8MOO/bY+blx7VorUg0f2tW67EZQOY+WF7kfHzi
MziTdbT4zuY61cJLi82uzzLAPr+JxmYf/ol67M+92yplzi9pbk4BrZbDj/09QBvI
V6CToV3yKIunTzPlF8Unq2T3Veu84I78Pd8PwpYLzok7DNx2SjcjJfGNpE0/JbCM
MoOeDJs4TQuTVf018c/GKpye8xDcd0Hs45rS2xJHoFIXhgqpbQLwXw2VHq6uaVbL
c/QEbiDnz8IoI/Ocyn1DNGCAWsSd9ejk0T9q2N6VbWguqYZaBTB1FrlaBLD3IL4C
iZNHoHJNTzeR4Zf3IE4sXF9k3FXZdKRkU+a0Q9ecHspSKXPw2wGvMyapa1cb8gyl
tbyAVYDTbKfpUMIrEMmnNi5Z4FxolhKWQVw/jWnyRIhg/L2C9x6ph+DrbNF1PayI
lOaN7q4eKKfD4HBiv/acI266vfn5aoKmP6+EFU2tdF4ALHOGTu2JOYCj368ikfSO
vdMskvnd+USTGNPSOS0tcl7h/9SeCOmqUSQiswbtxdVTBqNl7lWItxR2q8NpDAE5
vWk/0arc6Eb/Q2NDmtYmiElheGWqH+nea83DiNe771rmjEVuQ9HCC26NEPBx9dTT
HDwGmX3OEHozXogAc/rUc+8dKmjWmFk/OPg/PR/XdEfz8RPskbyWrTDqq56VNSR5
/iQ+aty0Ww7/xNJUvVoroaY95OguZDm4CCTRKL4CSm3al6YTQWV+f9lFkKTNr9bS
RoWHCX71EIpBNh0X7h2MTWK2v7FV7nPqou2iGFLqueyGb5Qr5jHasWT9Lp6+e9Q7
UQ04dHO8rhc7kpAWFqYmrLorV5rmSOzODyuTkmSIoLpSvLLEh5PLgIRIxFi9Y0vG
Tq1IUzYGRXdR9DvX3EFVCPUrIdApnxLdBihIarJLqpxy6g9te2EBAfjM0slnjVML
yP6WhEHVnt1IlFYWC96E+dFbFuhOAf9HRKdU8zcBC77mXPY4ddcrEuSN9WDMuIuz
/Uap0D1WKOhot+WAMTsdKXJG2RsAk6QbTzRJ/ixkYadGfNp826R/W9113m84EQ/N
k/jeOg0WaAZxtAGFgqk5SU4FwFdkCuW11EEUkKktnAk0xTjNeDgBoWR1Tkuxhze7
3kN0jKuQXjtHxtFaKOWbcRgrzq65vCXqf98BBl4zO/trhqgakPDYu68VDOgZL8Ex
wODcLBm6uk69KIos53pjQdZVPuNdRtLnxLFWYgw4ba+1/NalFde5XvjI/MmCReM7
FfuTjRFlesavZvU5oLp2hOEZIfaJyzUzKhuA/SiI2LNnqmUzxtrQcBG/XjhYFvKz
K8IztVEzaYYhQBvZQX7ATgVng2Vqt7zkQW8794QSi6oXAWb0n4wViriAdjx8JSKb
5C9AJmLPZ/nyci4JTNuX4HHQQzDmfDm+qHWXG6XpP2Wk+PTIY2Y5iEgLqmnYMxDs
xQISTqBq57Ikn4H8iwmqO28cwTeIGJ7Z+TPATavZt2sWGNoR/dOISl8EANqrtfC7
EcLH6YbJsbgVuN8nieLfE+UNiFEt2mRE5S/cq1f/i0VwmVrP4oWwdVKcRmTKXq6T
sf1UcXPDwYL1PjqwWr1tXyOAsUVR7mh+iQC7NCwtSrKAnh2t16P2FDgjDauxCeiJ
WtMGO5RGuX7rj/K57BRK2FYAdFuHib/Hzs2edLrYODKltIPv89xsm/1IPVddNRrk
NnqfLvoOzSy73DBJgcEIICsXpiPYFIcwL7yhROLjGzqOtrz0QlTOZ8k4DxJowkgZ
zjRerBzix93PzchaYtm2JmNINd933+1LujKfQkCz1cyVCQANNGExJgfdyAPjZ7mo
w1A9lsgyeAOTHzYR3j5CQgfK+S5NUVEMjYAVE5INIXRPTCrcNLsU76esrG9x/wF6
xSma0DcE0zVYw1siNhlaI8nfmYsxaOMuNQ6IoqaNdhj9hVltSjekmBsagPnHI3x1
cML09Dwy5kr8z2S5jAwpgP9OSiIKRsO9dGxzYzgWLDEBl3qYnNaijqo+jevfs4JC
uBVtL+BmJXzVSgdPllyOFctyjs+QiOa6OM8ikJv1H6nGx9teygQJKH+Z9dcHIPW+
pMkXwad3gDNqxBut1J02jCVvJFBoGHOtiX2yk1S7PAsCxABepS4X5pvrZ0WXzhNF
Qo1MpMDzcyNtOOOlRYkVkoEgNmREnjI6aTCxeVG6b6I1bwBA+cqwfz3Lm1qmxM64
uiuNwixSwixib2t4bx0JsdgKBlpNCVSYooPe3fZYg/Ox14Rg1INt/rjCioC0Tvfa
CCO2P+v0fg1VBoGUE67J19s+KegGa29Qe3RnvBVgWTye179KYdvWUR3fdMko3v+7
yJM9Jts0W0c000Yo3/Hza65F++NKL1kwjHp2b6ygJ2qo/eQGwwtVeQzqeeWXho8O
AjaRGAGskABGD12MAld7xKr3Xg2SxplGHampbvn13r/EQsLxT4WWTihcBzVBEhp6
aZfWmhROsARt3K66Wyq8PYERIefICQST6PT8qyizdJxLHgafqdI9hS39apk3FaKd
ypNNzDWFmXjY2orr4sQ6QjO6JbXWOfr0pe7yDEYQohQUe2K3Hcmf4EwRANzbe76V
v9rjNwtC2Zzq11mg6j3X8FhwTfdHf3hhy+W02uiLhg6knZTXUWeeExIpEPmf4XB8
gQXorbpOjEyH1uMxfNrAHiilMeUi1Gvf9MQto7EuA49QMbpmBtvtoP8OnMm8udsO
ON8YQQBr0v3Z34QrHAl7avKp8uXqi5LtHcQcoIlxjudBiHaClvsPDVbJDJXSq7GG
xSSikb6qbHcqWt1Cg2t2sXpYD2wM/xJ7NHrFqjZnJZZJRMsqdUApun6b7FuwvjtB
e2P8uM0Weq0vAFcSVF8K/DFmG3zzwVekDWpGvO6pE4+lCEZwKzTiFnVgMhv+N/iP
Li8FfsNIW2fS+qp0cSUgkje/HW+Qgxe2aTGNAkh4jRB79f5YtVCbEDKyOTZL2MwG
glmvLtuRyT3DhmUYSkrOXp6o0gJUN+wUwjT7CohIuA2Ss8t1mcEO+6WQaGodp/0X
lLHs5l6CPIS6yXoWYlB6EOK4E9z+DV5hJhfMi+PKDRoXBelszmZ7Kd2CuhSI3D3M
DZSSR80ecSj5GaUXktWW8W3izCUYFXj5Dzu7RBQ4ZbYeH37k4RXdH1R/20jKjlKt
3+iXd37jjcQBmCvKcAl2wuj8+YN3eA68BY90bSzm+6A57jO5P8GHO0tv6AehgHzP
Nn2HtXKfXZqtUGqAc5PgEKiPKiMj598JSpmgYXhAWVmTgoBxd7QmNp5DDpzCG6xw
kf0ftiRmuhoO7GWjzZpQKIg0amf97DWxUtCQK6B4J1hhHR6Gt+vMPac902fb61s5
+pVQCfrvSVObul6TDRSq5RqEuh9wg1Ondi2Zz3GBDNw/e/FXr4qlULit8Ha36abq
KopA6ljsVPNVkBCAOlu5fjL6nqTv9XMQR91jZi4Er8kjS0NfXs3Qtl4gX9P9WbQR
OxrMsy04x6n2HikfaXyeDuSKkwJSTJhK5QrgAk2MGO3Ou0Tx21N1/38gh+wPeCOS
62hhVntLkz/ITnJw08y6xNqWKBaPvTur9+gZu9b6DSV/b8aNMXAuyDIM33dnTsYQ
i5/tSjuSVq9h1Di7ARh/0QyDN6RFKRoztxb11becAMZJxtAWKR5yNDkjX81PxZUZ
BXC+ixSD7FcE4P8R9gGC0o0ihP3cSUidwh4/PaldO9OSVmmbFY+Yis7RPuAl4NXL
ZTQTehsFiXJjgELnGGwNrR1N8BuGELKjHi5NoY9k4QRlc32ORQy4/P+FZY9/HBpi
aY4LHWrYZ5rXjVCkpICFUQepUNg38tGjFyB6QbxjmlyFvLUBEJparo7T0v2sXnXE
z0Y70FTY9SX99DZY/eHOrXpnNzoiMKDGhGB1eIXpfHTYdH5lhSx1TwUCwRb2Y3Bk
OJnswtdHFmNuQWfKgo73A27CRNrhgRhurHfNTpsu1II09WwuCakAA4N68b5/51b/
xWysBhv7f7Zsp2sgiKexq0wk3ct+jlXMoQgfvNSL6VkBoJ6cptjZMaj2QqxNVxy5
6D1UqZz2OeQ/jdvrMa/Dv4dbeR2jI/CmX1gdtU4NqdpO4/Rc+XztVEIGYzaA6pfN
Ec/kcunE9KC49jFYvbbnqzxQWBXzdJP5ELQHmMa3M/F/reqse911faI7zzwhCy20
Q7y2BhpjOJ2vgomUMwFS66iTEYlHdw6nA9LcyR0i5QeS3t4ji8nFaYdwUhvjc66x
az5qyfx3UU5wLfyiapi4e1YoIblOBl+p/njrGya8rVUPd+TKmrG/z8rV1auNfee7
vrumUGmbrKp20Dpzc2kCWV5KFO7G7tFkjZrav86wXBs7iHQig/K9h/t2poEZ5BGF
>>>>>>> main
`protect end_protected