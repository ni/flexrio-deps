`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 43504 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
093PKSQTlIpLKOLa9A382RrHnn9NN2HzKYpA1RVc+G2TQFlO6eEgyAaqIQ+BDPlD
HClqKi3GGfzc1lrBkPONZU9l00qotx6lX8A2/6IMkn0gBn3o+EoPrgg+3GxxYfQD
OrkVBZl2+bSoUc2Y63XoAIP3uoqMIL9mHQV4zgnv1exvBbtxo0CPzwWhqEEUTyFX
7CXtx9Svv9YVxCy1iAFhRekDdsgdbttjaBo6Eyevj0erL4k1GYEr1dCFrw2oMofE
vHKvh0UzRqnUH61rRJDkBHU5SYrngwLN2D3neoOgT5JQ7xGdMwb1APvDRAkkEd8H
g6BkKa7mPTYxarQ2aqQYOp0VcWb531jZ5Hri1DE2LqrDyPc8m3AUKC3zCk5gmOLn
ZyQ97bXh3eh/K24Oe2q+bSxIy3vaQ93O5PVC+L+oSx5NmjNFEUHIk+Y/GJwVhbvO
CZ+Qms6QS/G1auzUfNpulrOCq2Uctz2KlKR6wmcqlyLvwXkC4jqXFouUXIhlh/Wp
jFFtnIhDN+h6qO4OqAVLv94ESjEgJ6jwuiDBHGfdea7UgGv2tJjVsByIZBVuiHuX
CmxMLR6dZb04A0oeKB6C4pUQA/wlHcqOOBTZyGbTdaPBGi+FpydlDTwdYtLhD9jd
29XhwVDaBuasrGbl6DopzzoDocs9F4FN6yWALzFW6ZhU7Z/lYoMWwn5DJBedN+vC
wciDFXGLnNWiNr9/9eTY3TOxxUkM10CVVUeuLCkjy6gZxBMvZskh8uKEkvA1ouey
bqjnLztI+lvvtYVUs5Izz7e9xG+gAKd06Eg0Vyzgr43e6KNvE/ehb+ZKaZQj7Pak
4OfP9EZmR0fuNUdjPqaUgLbkvFoHQFOhfPvTw4a8VEflthg+crbz/wHXqNVNRZn8
R75m7eoUBMNa5lOjxmt0bT0Tjy1wGN1uLiXrKw1Ei+62HYrkZlM7IK6946cGnuDB
TeGWYB1BDIAQW7ImI6pX63PwtFD46KCFz8BIuNxP2En3oN3XyhvIRxzXB7SxxyZz
rWaXhPQa3dDN4vuENHyFzQGFPmI2xrjx78uVovskz3wBNOGIWswQ2l5SoTNps8Jd
e4i4jnjudjjRSpFOhtiehSZvfNz6yAppbLqLxd6vdHvcVb+MqdN2ASzxKUiAy5+V
vx1JUzuGWCkJdfeYK03mq7gvjHvU8MibKLH8apbya8lEYV3qMcupNgPxQTC8t3Vx
kpIYUDUbr43F15NiRJTsBFQgkQ8frpHkz8RSx8fGZBRcWTX1i/ygGlwmR9AgCd2H
Cv5kLpUqYc2OLEi2VuQeGMM/i+7GIwjbrX7fC9FADbFISJrb+qXETJFL+rtwcNsa
E4crpqfY3IDodhOb9qb8gDrok2N0DScy0AiLAcrcKSae3HlMtCsRtdYQS5DSXWdU
0bOrFPX+f6Rcmu5VXPXLdwZptGgXtAfeIsUlmT05DTo1yNJzVVLclAWgZGMsYHxe
3tCS8mfQzYs8LO4/szyDkt0TcJPp5/m5a/UdXgiqZB5PlQynngg7JRDsmDVgqEW3
TaTVqFwE1LYYMow2WCl1vTqR1eMw544s+3ht67POEyt42Zj4FI/LAjoWQnDT/DIo
fWjA+mRamV0ew5lCG4RrlgEtAd15lI60yiAXizxGhkYa6guGSxMnqFyMyolMl7V3
CT4qMCYmTVwd2hCHrrCF4ULM24O1Sb/RcOPD2+qa7LkRjYcfpgupZVm5H0D0h/uS
pSv4MACesgEI9f0ANxdR81JZPvbJE1LmPjx08k3be/TJDkhhejh1DgnLoW+Co1Zw
yAlzupZqxbiH8xjlnlwpbjKP86yrwZWcgi2IjZQmHe36pmvh8DmUJ1hoWBFQFF+6
MiSLWmvXwBIW2VOi6eQvTdTzznrv40zYPuFuV6lvxJll419BxlHDg04B2HE7Yc0R
BVebw+bYN4Do9X83d4QHXPSGJ+slA3A+0noT2RrLJhmTa6ZfNmqLoJETPrkB7jO4
+N4cUB5VEant5k+jzVgSTmcbjkj5SAiZRYJNI5xtltJ8aiXx7bCc/R5P2ro1syvb
JHSTr9PN5Lvljwz6fnsn8Jy6kWh5s52WC4Vg1dnynJst/3VRDxvDH/plAlGGyYd/
Ef61d0IwzxHYgELK8DmlkDSZua1Xa7EBqvieib1jY34/BjlCCIWZobqCG8m6alGA
z+rs7bhlvrUM53knwKUpP2uooRZC1saWIz036Zic1u/StvDsbKJSZnmQFY5cJ2ZB
fEOwgQpmuoe2xkSGGPLl4WRDmFULntrRCU89AWpFu7UwILry1/mLPBcujWn/kKsl
znVh+1ANmsD95wI2Zf/tsy1WFEgQ9RbDpAM6m3+FtcONxvcmFxxpIgkGji+/7CM/
JsIuF1zJSeypWl++RxoTB0c0PaVSG3AdFo0kVbBZ0Z25vbLBJ1y+71Ri/3vniYqb
nRSGg5czINUmSBw6vAjKBUeVjcCcNa6TiW6T+vtbk29ePZnFIfrlx06k+PF03uTY
3z18w/FIldu6dzBeyQxmr7yllhtcyJjRznBmcnZ3TM6JQz+46BSIyvve+GuRFiGz
kyvo7rMYad40gW2kMfWJIQI81Qx90DttecfpBF2i5E4HizJFqq+j+z+lRk74e6DF
ywwajfysyGYjJQbHR1N0IbtURiQhOnyEP0GgvUq0RUHM/nc2eU9NdnAk6QB8VDOV
wCRwVrDq8vq/u2x1ADGCCkwbipGRa7JT2uoIAxzQe5dGYSvfo2i9uP6sLyCB+MzN
7gBdzSXSZTAkVCMLYV6joa0INfVMp9gfa/830sRqnIn6dIL2i7MiTpGraBF37gde
jPyEdwGjv8Yx1IrbMijdQorf80UuVeWIyIrcfVFF7EUwYW2gWAFBCr13XEapTrPR
GqPm2yvso3mbbsNXzuZk9C9kf4evDgBVoriA4FThi62p/RL8YlJb9+7pMi7qGaVW
IftgiNVvuXXqP6yQubYMSeRqu76PBdf9ZVE4umyMDvBnmP9neJDCbR9hZTuv50PL
BM/cjqPLu8e7USKknT82nplb/rJZB8DOkPz/1xfrCHuHczOmNcfwNs8Yt4z/u3rY
4EEDMLi4ynTRyW5e3LgeCmMGNwVKbIWdfGVs5UlCe5p2zHjnEuqeOO8CYRYdIMqb
R7YDmJQoUk+rLopiYRJO7uWj7M4CLsvZ74hBVG2RlIQvj9IpIpYNJKzS/kZPuimK
l2opG9oT3z1cAm6wI47Jg/cKh7XPI/LIEnHyQVX3zwOv/x3xWE/+IYNBS9lcS4it
P163mgutlMs5eejYbs9CWxAlsuaN9fGbowXXa/tJNxZbpJCgVkdZTM/0M1q3p2lU
QPpwK129psTEJKLVjp6PuTwVCLAES0zzidqOBOUoYPWFlPy6zVvVJ4AbwsBpzUtk
W5l2gLlQOEZU0Xz+eHJb0Eka+fxH/EQebI49O+C0QKjlqMPpRp9/Z9AhmtHAGbq0
pRBLdE2sbNkue4yqpp1/S+G9d25JJ8uWMHuOgBk7SendYuZ14eASNUSgF/HpOCgu
91gKp59uUTSERnomtT9kfPX0dn/Ktgdc/VsXY6Zp5nNT8XMnv736hC8HL1yR1+rN
8Mwiv+orSw7P6YUBGVSmBlLe9i+4q5zy2TZq5r3wSF3atbEcJyyL259bf711a/gL
RjYBMEqzfQgxTUTeHO+EDT4Aw/LLak5ffUiJR7c1G5MyrGd6rNR9W7ECZahznPY1
948gydxCc5Cd/Hw3PB93mUxR5MQvCcjgqkHRvmXT1TttX8YGr2oP+7Fx5Umd9Mi8
q+batFHm1ME2DV0rd3caZs05Wx5crusGTPF8DPG73PELXsFzCj9blOFR1zc9NCFp
WCnSy47ENsEqNntDMXXH4yK80Oa+BHk7bVAalvMn6rGMsRAbOKxyi047zNklLc83
uldHLNvvb4FPnPgi37frthXFqQ6lM3jfJSq7gHtVK9Mz8heimk+mx8bfyuwxD5N+
TRNpeeVwhyVnr2Fn8o50mlXtpJC49sQ/On5RsEVG5FeH9VgxbE98nObX2njChFAP
w3zkU+LJMHKAC/dmu3yf+I8BVZP21HsO7pqPZ4KMEpTmrX6EHdkFcdvHT4aAvkPY
Y9gcKwrr/r643SwTf3TDuYQgBkM3WGgI5RIXVn16R5O1ERI1wKYcBleSv7vb57py
cKwh78jLwWvnEqLZihDPI2jlqrGwnwGEbEr9NkNeGzRwFed0a33RB9h2Kp5xmT+D
Bvx3KAA5PJZxTgXpJzT6I4vw+2b/x8Xvpi5jAk7Ir5NavydnKy3nCXZQOdM1d3Ou
geiKhDdcOvAOXpfRASHmEazOHVnZe/pgaZgsbD6VupO7AthnphcyzvW9LKsENWjS
CkoandBxV5beObb9GbsdjtUUbWrgZAr1LvJfcaA6XggKXwqpT2fWdPhW8qSZcAox
NS4ZseX+MsPehLtI5/+TitK/lCwl8p1W3TMjFw1RYHI/C39ODj7s6+vdSOTbZuvI
kBIaC0mpZSj/d7GnD451XRSEJJHmsX0Yu6+PdxC0fQ9Fxd8dveQRMFcXrG1eYTAs
WPSkKq8NU9lkhuFiPaqYsdfodacIL4w37D3uu4zmy21XWBFuE6OcrZFWs1+tBxO3
OroGO9iP4dA0Pv2ccFqJ8GvUruUXurIBIQ1mX8T8G10NnO3iJQGZAGw3m+B73X3Q
o2itawbSCnCyLPc488Safa4R0Yf2f9kf9t9HlZXvJsrSpsoxzJvKQ4GTmqHTiLox
haCiINSpwin4UeqlofYTgtKtKivHxk3I+JN8q0LWLsceFLvYy2OqrNyjGn1clHHp
1a5w1/Um185wtWVATVHVH7gaD2yT5m/zfBQV5O4Z733lMDtO/nCcxLa4l1DvL2Gf
LGrSqg18kO3YL9FK4Ph2SVLqQSwzvlaRejk6wRxsDNEeUhwLrLiCuUsGXPLUy3Pb
YuyiwEFI+j7wsYoJblHGRP2UW28fOKFw4QceGwxIag5TISKoMvyKRZ26erc4jb/4
cbNRRIU0tZirLN2QDY+SyAji3BT6nCUVLTiOXIyoJ8ZtK+dFDxUo44NJphcORLmJ
pGej5dzQ+ISp78aLZspaRcOMjFRnm8dkRCmn/opygAmnb1NHxJFf5DzlNP9C+uih
vxbhTGFqtf/eHtEgzaDbcSyleSfBP74OJ/dE3+uc+FIii+cM8bgE09AUEC/fILtT
YyL3on4A9pGe1ONViUKECTauu6hWBGASY7WRKmb4uK1AnVKRJTmgWBTLQxOrQ8ck
o1LVzybKbssnaXlSc/k83LSUKXABVpsI3sZBTX1ArF2kvnbN/bCRlp+ufyUttzzg
pTEE1MbJBLGSR+e9b2wyfj9UhDWMa92nPpVuPB0gMuCdKSSyxlk6iSSx1oNtJ6Wt
CuUDvGOsJcuIUBYV/Uwf4sR02s/3vOxa73wbV77jFo9V0NwtUNlWCtTwyAztXFbR
UsJ1fHd0Wp5pQgpX/WKTzYRYnGAu4gepiItWnCqw9hwqfcK2FQMt03FB3O9o7Evs
lpPhK/Nwf5mO4YMQ1R6AGsm6HpE6+ch2oqzuubExEUlycJq97lxOYGYB0joTKki+
8siBMBBwJXNM9oCIQqGHhnd0NJUHpWZL6QtU2NFY56hv6aIGyfliH9G9Oagi+57X
addTAlTlwhP+qvdKjXHC1bU2De6zwosMldtnzMtxzcavkI/cjuwiLojaKUAd+uYi
jU6P5ZpcSYFeR3C/LYKEECY08W4mnTYofrSO2gwxaWcdOkeEPtmPkBAOg1LhBnZG
vUPEMP3Upku3TpoAfNjSpu8shaVP5VK6quKvCDD7HV7Uq/MTLy5/WfTNt8m6rwFi
JR54DqwXlztOOP3bP3JvI6ki/DO1Zk/8UebuVA3G80om17+vb6SrJV49wdgrBRhH
gROeL8slIdcHmP+EiErMzOBK1zQ81nQ7P45Dek2/5mB9ilCJ3uXGHCUUkFs9zuSP
kTRkViMbIIdSN6ET0G/LpcjpmsIyi0mjGvS35AT2yEyCph3ONtjY6iZvXTmaMoVw
BLotB5s4JURIkyNSJF8FJK8fc4Gduv+6xJL5yDEaFiTugdOrpI/uElPNI+Xp0QDt
gqOMNCTjxXMLbgdxWtP74ntVgJEpYFqYSyvO4IRNSmLP0HPffVWWN3jQOmy6SVxM
oHj7DD4mBkju7J8+CCijbNdwqYUZNujQBO/b+bBicwB0KoeJc7E6n81CTjUFtAmm
1vWO5Jv0A4oGuVfVwReNxL6poC+reqpbSv9c/4yDcFNJgRnhVACOHgHU0TEO8LRm
FfwLXY6X9Uy3ibh1Rmo8Eebn3eeeyso+Bb1HHBgIUEodtZ58z1k0d0Xejvb5JZv0
/QHwqCf4o9/FlEPHah3XLcAoG8NqVmFspfeqIdGL/SYwtmQGF84IQoUEfY3s9X1f
99rQ92snTRKpLKknDLTi10uGRTfEjpRiNCQ481zKA+tgj+c71xtWIo7FCULcM1+y
FgULKEg7k6tUloIwNr9TSYR3lHE/HLLLv0uRvamQT8eo7ysnzrGsJE4GBSesrRst
VDNaiWBYcybSWu6dFu8RRT0ywNoIZR+7p7QE9AGXVqpXUve95NNoiOXN9/zY2FRL
Bwe9aBHhNw547KlDEnacG5u9XhLP6EuNjYKhyKd88E5iW2tG+gtFl545RnSokSBO
kIojioHYXm4WfbRxAm1fBAp+x71yHkiAwzMKzqT3HC0Xj63UX/8T8BneVfB1lVDL
WBDP7ziqmzOGdBak28uRwu3FXIARE4g6DTLqgOUJZoOwRpWsnMZR4+c2QD+oL5jd
60PJ6rSA5LHMpSJ9SlT+CccFsbQhd+jPMzZGEJO0roa4wddk7DoNiaDaU1UufStW
xqq4X+nw4RrdjnNacsY2GMPFbDW2/U0Q67+Q1KztDsBUlZ2a5DpxQDAOXcQ/E2gu
zdqGPvE7N18MrOTBnS+U8HT3Q2V1TuM6UjSY8t9RaEHXxtilnz6L01C0sDLRo/oC
7td4QiK/s4tgjL/Tyy8rBt/yyMzVso5Tc5uBLAE+X7GzD1RnOw9NgOx+hX/a0b2g
dZ9JlZguYQlPfd49NhlNPQTFM9LOvq75WdN4ZBXQCC6bywnB35aTZAtLhhje+rOS
cvECeVPW2WMm5Mgrh00deCZwUwTmPAqc0hhrmgvRBkOMeVQO/A0R9eu/ajASHWLW
C23P0pv8vLDoGpWLNRGblhhLqiPerGpOymJszen8yFP2hG22tYZ21hT/gbuaasXd
NrprSc/bxW0vLLntib++yD5umldgmuEaDgM0rpn+vVHe+ALhb1Aii9eqUr3VICCY
oJZ1YbVc48TmvJIenTdludAdFbk9R0kUMyTou+2GgeH4/+e8LjAcGK+jX207tnT/
TlsD4c2aoccBABzTd5tFh3S4mFWAcGFZAXdgDLhSLCJGGQ+qM1oltg1eIA5qCjQ4
nb7pvtIaAfnxHwYFmky8WG/AZhUnDKuhPshFXZXOy3ZLKVarfgVoHzXanfz4+HlH
B3ZC3kUq3BB44aAwGQdJAiigcs/cLtU9hlCTgiOEMaBKAyR2wP362QA1QB1+O75k
FtRN63C8B4iRY2lXIO9gYzWctvo9vyAjJdutxYX/+GYBebHR3YtAk5wkwttcKdxi
4FbLPV+r8GAlo6S9DxOdyACB5S2luso2uriu4NZxkCZGT4XlPvp8y1CJegtqP70t
y0Ti/dWKwPzZaL5P/xwTGCLD+5Owd1242OPtRycX4UGI9OK3Sz40EVhLGl+xTNNl
Sxdkz3w1lI8+fxO89Kqnpitp6b/hmuHWiBII+zc92peYwb0NCfzfR2uq41aL4QcV
zmtW5S6tvcxYqFf71jMfUWLWTeW8khCpdBEg/xPi7ySVyinopa9qBPVyPfOOs7mL
iVKPohnVrk3jfw0bsUsCqHgkUSL++5SFhOMgKp0ZXv3j7/JOrXLwaC3o4E1K+Xce
TKC5wYeQp2mngw0IshDyv2yCo0fkkyYARRSApWiYz4Uw/Yfp9L3edghkZFWjQaKV
0N22sKtorrTuDuEnoRAatt25sA6QyqJtfaiGMmS2TASdV7v4yGS4FFrMPfzudF3c
l5EEuw/UeFj6Fc0ttw6WRQq5zA0/vcLA2ZWtivjYhL0KD85W6ms8xIxhWLKqyxgZ
CeKgT/7754IhGSLmsvPFyGqa879fm2lxGn92mz71EwC11RkrtuKyoG9Dnurl4H8u
IlRClUpofJT7IoS+DpLwx1b8c+Sh9rKU1oXK4OB3bvtSHmFrtPJ/u4DoN524+wwL
4oiq+6OGD+GikI65c93TdCb3SJJDrLjKBL8gNLrhzu18blU9LoueA81wRzr8gy9M
n6vU6oLYec7fUz+hNTL797G4lg1me+svUURA970mUxxeFPh6dyZ7knWpMT6HiEFl
w4BIRbHeqh7KSQ8KgO8b4drV2O3q2Pn1y5/Svw5FgNT+2yHQGdwmxuDGWcj0dcKN
8jYNZ0ndApxG/ELsKfvgyUZenle9chUflMFG/z35LFGbB6BuT0z4moENywHJ4Quo
WRSaZrO6+dcUhuK9xKdXgudp0BwRBWd3XGAZ5ayudHfDXW3FQzvnbPn3zIBvZ3Ed
XPnjK36fkQq0WjYsm2lBTN9CRTpYJp98ycmo9vVz0VV1TzPyIet8+5RZgug1F129
AaETCRz4GTnJMocQjauALjt2Q3bdKLno4KBRciI3Mji1+HH9O89C14tUBu9cuYss
sPjng9gy8EmsSJ/2EgdogYaa+dAEGo2iOYlwG3EWMxc0XERNa23W6JAVOeb9qpLf
6ySSe/ZIwQQRYn9uij/zSvOSwjyHl7j2OeIjAb+RZuwVNCNi9VkfWZO1V6KyNrT+
zHM9OiadmyCaxBQR4M+13QGUW/PRYGWQYstQOI4oD2uS8/VMbn6hJGfouPPDPpUP
ENPW24nuIkjdLLb+/40/nk+C4J7nKQJjnPItF+SnPkxXJKuJ2fpJ9EymUaPfliDy
4wgdsxtq9JFygaw8f0LaDf73l87sEHduKR5Ua7O8rbVpyP3KeVvpGB7WDtMnwZ8L
Jtliwk47MkQK3UKxIJ9w952RiogumTEwCno/+zCwhglm+zSvmTSr2JdZk9qeVGcf
dwSdeo/rLJNsIf1ArsLuu6U2iUInx2EWepDCoeMiY29xb35SS5HiP+ZKkqrMk6HH
i33kbJEPFi9MQgWwcu+fEnAbYR+cXILML9sdZ2hUS/ucSl2+evEuhMZI+wfmq4KH
Aur+O8wGCVWgNj/LoMnCHHV+eo8W6S6ByvQbWuz8kfx84AiykkMyAACCYesgHMxG
4Qgs1v0sncQjBPSaWkwFrfrfm0setZF7zGW+PyU35U3CEzZqpT2tCDMliZ30jS5L
xtD9WtTmN6ThJ1vJdu4HWnzuX9uk8VH8eAW5oI6Yz5fTvQXy6JjYViObPrNav8CA
cdrgtvXP4t7ecOIUp+6zHMd+3SB/QJ9xNdeNktCHk8BAbIxWCnPmIYRdsoNaX8KQ
rh35/eVPaFo0oinXVG4IaSBQAXUg7bAbPDH7DoWJCDGikhY0i4ahGpWpng0VbkBN
tCLPUft69Fy4jEh/cjd6vt5Jk4RWRJXTLofhy0yjK9zevW52NOEwSVoI5ePbGXIi
7UHAMnFh5hKuXBYodMNqDXJAchKF1TJDHwmAhaoeBjyVhckUe97XAq6gx1e0I3Os
cxD+V/hB0Dwg8WNs7t/lPmEw+vGePlMMio3jkD54IIYgNxQY/6rYafO1CCrp1KVE
N0F1MBKDvK/tGFQt7/yr8/8jdWisSadxiY+xy78e9Xt8IeA0ghZVSOG8uKyK89+K
mfADGoTgPmMEtkvR4b9Us4fVNxgBASiXhuKwVrVrgQ48p7za/ckvgjffm4UgyJ/f
2AtrevtQauVl2bx86EuBXQz05MPMd0r1PsR4O0a86boYX7XX8Nl2rJPRfqaqXDbZ
mVMuExD0cFBN639faXz7lSKq/DIlc+pAGU9cChAf10TvqUoqVyu/Uzk3Eokx4eWh
Q4dtyPNsls7/Al42RfJIhwOTJOhalpGQJ7wL3qUvGvJLAGOsRVkMuf1cL9cFaA+d
2+MSKjPBr4EGOLK7EM1nobjq/Ia3zPrrRCJ4zcSwDNKhbP6tKpwnS0qlyEBhwdzk
AuQZQ1dVmdBYDr3M+XMQZ6X3WxOVlDKZu9vHfBWHKKISMJEDuDjhrGdbKgr0RBVR
mcxs+fnTJnBpXNHbMxYaQxAD6/jTrJsI63nmD9KRXLwrZ/QYwVWPv/vHkcV/nWJt
S2ZjNSUQ98JwfsqrHfgxf+a/9CozY1p15VQXbnOLbmfbLiFfF5Um4NRp0y7YJmGw
ctkrgtxr0fwh5KL7bZro7NfIF+LCX7D+v0Ibgg423H3EZ/Gs5YTPTnNKyY8YUIMO
W68hfNezCB8vMNDgmDm1FHFgzAE8fe4FxBfM8TSDds1zeUgUUzXWrWjOKumJBEyx
f4sO1a+4oF1EKiYAG4pJaNL5TrHonZ3IYuGn/EXc9HBy4rVoqgUEwp//HkiTaJnN
ScOy8wbAc+mrglSiWboXQE+MDgLqOPfg5QoJo3rTv4v80RN/Zhe2cpVGJ1STAsSr
yfzbDJn/dzE62E0egT1xIMmRpmx+yGFh7V9YK82ZM6n5RGJJkjClPO4+T/1VVCtz
X1PJcaQfbWrCQka+nQr36LR4yoM/8F6GqmKCA1vb4KmvVhNGB0CE9/WAXi2HLlXp
ZtlgAomR0pGOXI7W7IpQozYZ79fV7Llu9HZthAc4UN/t2vR1KTyjGASgmnGzplLB
x6kEhwPAPHTasfqLmgkknrXZzAfVOQbwo+syi/AT8+A/h3GMlOHJzv3d9OZDqXHH
uLE+t7bPAmBYAUHe97prr143vGYgkSfuWHhUeMK555xWeGuCaXQw/hfy3cRhrpS6
V3TCfHZ/jVCbRnAYm51SXKV0JTg0GhEPnJ34Zuc0aKXhkvg7e0WKqalC7+91Qtn2
cVf9sgGILL0hgzIhX+Pf2oURIzQUS9LqTSQaXScPHNRw+zofzI9o77EHLv6bhiJD
MIrlpD6rmUOQkkrZ3QwMvIfYVxRcaV22twqDfxibOghw0QthZQCxb/Yx2lrdpb7g
s+0aUXvuxyZl9Q7RLPi44SkkSTPhFknoG0TLhg61MBxMHrNblnzJ8MyZ0uTmWJW+
L8Nd1waRR07I8XbMB4hs+bewSakjzKFOSCjGjogQsdNTYpjctUcX2sEN0ygCD20S
Okb79RQ2zJJRd0gGbdmOgSJ9u9UWqhTsbaQBdjrlKNGdfff6sTnmWyQ3gwzYAw1i
7Jrgfg1Kv6RfiR2Aq3tTMbGWudi8zJOWFjumFlCp4LEpCAX2nujCpdlKEvwoEFCB
9UASmFLFP1JdbX4rrQGIRYryOkLKSjlzf7LybS9v/cITzZk0s439r/KQdtVIZoTl
neFGKEfxVzHlagPJkhlnYLz3x7lSuLq91bu4d6PWPkSkYkedO5zAbum9cFFkGl2W
N7NSrDtp/Gtj0TLSoPrvUMOsplEX9IsSBemgYuxdXVgjgm3sXR7NY0u1EXV2S96+
qJQ4QMvl4CsZLVpNM53wV/QzLmMqxzfesD8RhFFSk8uEaRN8rQOHMEHNrI4vIoYe
SB1TU8Ne2cuxa3oQTqpnHzMMuDpHCvWinPBW0DWVa+AZTtLofLxvS+NEx1zj47+3
TKZ533lP1xAdUj+42YxlDzVOP5+n99RYR/5O48eANGVncMYHDjU0OnE2lZpye9Et
Ui4zLjREWYMZwaeomQ9X7ctiqaOTsYA5vAt21q1CEL+hgfC3AmNovP2IViws85kg
xJ0xgoQf/tTpRlel+cQzEDquV51F4Dxr3PswNlR1bIBMvvXcUTc2CzHfUt2stypE
ir4zPNKbQRGCV+868qG+KWt1pFDmU7VlJQH1OZjPU64SRJ1af06W3zHybb78qk1W
FSxl0H7yCTqtc1iAHFy7rZSFgm2IC+nNxn1Nd28q179yLVFpyf8AuTI5vciMybI9
s1Rpe/2MJeuw4ICK+HWFqm5m4QpFga8Hi6fBQeAiLXfbGRPE9gE3WmZvYAzSe4mr
vLrVYGomnVPsHNSPU4llRRE5+twqH0QzjRzZKm1qKnPAfBNMqoVXG4wlbK+//nq+
bpgpWUF4RQBdZGY/tJbmKWVMIM0fGVDRsp0oN35VTG/K+xSDMDWS7a4p+ckqAvqX
Upi1JYcsyvkVbh9mupKDt7BFJdg3VvNBiT9KqOk/c+0ZNGKXZ5iyBDI+c1IWKier
yXsK2tkE4hhKD7yjteNV7vBMWYSTpPaUjOEG5DT5m+IqRD/2N/FG3WIR3e05M/8a
wplV8i7UjwsAKegE9TA4JstDMvx0HjE1n2sR1SfqCW0vz6lN7zqQk5LeyuGI0+KM
D63xB3y0d4ZGO/qy/ZLpIYdTarcXj7fdrGprrpIkgK0iuRRFaM/6HTSFzhOGxBvO
7JLIkZC3bEY38MTc8AfRe+b8ee4c8XJYLEKFmhQFaVwZ64wM2KnVmwx2H0dPQxv9
QEAthPwewCaGZIpHRxzqIVYD6ASfvuLmHIMlQyqsqm61rVjFlgtLzHTzKrm+gNNq
OONJ1DcYDSpuy7XDVbIOVh5kvM2qM0TJ6PcM+i9LGchFyxPKBMtI4vKRaF4NcGhX
oDMpLflfuZozM7ILIcTWEDMMZbv7H+bAwoAj5zBBHn+7c6qko3t8YXE44tLhUEo1
RRxO1SVkfvXCbG53W1QFpjCkou79omMkUfNtTHVpr8KHhkD4wK0AqgC9AAnfUnwr
j0t5lPtP+1iJPjIcADEzbNC3vM/njsxAhqe4kcDy57Nk6YYdGiErR2I2Bmtw96vo
DPFHFatqnX8baiE8NNyk8dzmgbZ93y9hjzql2b+PREy1Rx0DUgSFSRwXaRtMJW1b
DElVWCG+nywIj96lie64dF0pepUHVegCxYCiOwGn13xv0SrZgG2y6M56aDJ7fVMg
uNKoygaTM7t4iZIHYblvLpnHdVsRy0jX+T0nN2YkbJqgo0NiM1zMwiBPsQkeXbWx
7FzG34jcXEIBkKpaG/FJfcrxRoWUN5GnOF3qXHJVR7o6QuFgPUFZ1WMoyHRudTTA
LLrqeOTaWVwahK+hoPsGu12LKRg1KULhpfJhaEYnTk/8PuIRulpmIVdAt92JT66l
EDi3KFV2FoGDz+lESVaVqkTQiLWRDIJrL7SvKRe55i/g2AeWJri1VmCrwONhSq34
IT2bUc5YM+iy3r6rYbb76bMY5juqJodhyEBvNQnxdrHrrw0J1ZqBqiDE1o9A3AXm
6ExmTVf0rDYKRTpY7maAF+lwA+/TueX2emZ5iUfI5Zad1oGB/9Ir6gAGgXtngn9F
WZH+2aII2788wWUI4gIuuENk6/ZLaphE093gpcuYIp1btGjdreTE1DZWdVGU3IDB
j+du6ikWgvduWsvTCsE9hgSTzlfeES2STdDc8dQeVWRiG6ieXMbLfvnn0RUS0eSd
HAZPRH5+4Le9cCRjExXTBLyamQnIdXhJ4D7ljp6j8x7lUObTuGUtyaDcVBOp2csx
NCQiJv6e2USHrVRo3RFcC93++gf8B6Rr8V+2IVWKc0SlbPI1xAVZkrQl6AUEv2Zi
tmvEbjXFr6EB6On/DrwYdhRa8rbrXg7omz2o3aI9/96poh6rT0vKjmYgSHEp/XHn
mqn2tP9aHi8/2qQUWtpn/9OpE6pzlaaqSH/tUiYYuWUiHC5wFSV9JvOxMJqlCxr+
D9M9SxhAQVHHKyocCKOepu4ei0ubmKadPuOsdgoh2c+KUyiP7lUzpSkPxhR4+Nxt
aadb0M4FUH2Msl5GMhpLT/T7trWI24e/ZhvewGgrC6SyjAZ4dvLIGugl3R7C4BH7
08yGPbEsGK7ZHXlzfaumlz6mvlb3pcNawQ/w+jNCiN8o027D8lMpqSgN1t2N0X7U
JbCWZZyQm9WbzB9foTggZ6ARaUmAEIxVoXHe/Wz6xJ4gMdtCMCR2ld49Sn+I/N2m
KoRr4ng0dM1of8coF8CHJ8Afz2X3eH9p6iAXzW/bpD/CVmpLxC+W6VhQmq46k7qU
sCloOieWMmj6kjfkS79vsxwCshpwcLAh/Z6XVNmvm9jzVzl/qkfO8Gvq63oOYx//
NBERChwl2ncAyP8oXGrNVWKY8OnIO0XO3BL+4n8AKrBzWs4q8/zsTQtg64DRacey
cuVVc8GnEjVZVvPas3UumVU3LqCUQAbXm8KFxQLut1fZzktmfyD1zMcxwgRB0fgQ
T/N9qss7vzPKXo/9XXVya25C3P13WstCSGcLrM86yezr1mUAWc3rAmZ0J4f685iv
qS3LqVLedbLOanL/2mxuRo8W6YGcrCfpD/QZqh/B0sltkP8NO2R6jOjVcfxV3VjE
A8420QvJPJEx2O2SMJMQWyQLsKDrdyD97pAHHNTKZ4uBZadYMWR/+S8qJ9NIUx0e
QlF3Ul4GetpXCtkxs8i/71LZZOo/N79hBuZvqd8dHO+yHeosCOhlTi0p04r1QMWp
YpV64/1ppeyK6pJuNmp6pXyWwl21QjIhWV00B5fvWE+c8vQjE1eL2HSYHW/qeH0h
uEh6P0eGGCiPK0AQxVTlRDhVdnf4i2Oapt4nbJOkXzmiOI8xFJVcdOExRqEog0XY
4qA/H/RfJCQnq9bGZCbmaveDBeo+4YmE2M76ZJnUDRDopC74eckXcPQqna9zpRJh
aSEiPnAxVLgYCNfug7joFo14YCdXs4iQLfwadREr6Kmf0SIqV5MJ0Xp4fD8FckSR
LSbNViJUn+ciOK1yjYFMTs0B/tghwv7vy5OyMPXHQ2GBVJgjTRa6Y5fxB1w/hEEW
wM+sfsCP40oD6FWxmXi5lrLFDxfhCOgjeqfG3knSVgm/eFJWCbJDhorw1gwCtfON
VuBjVQCn/uareRZCYZfgypTrcClgHcrBkkJIhUgqDJijYtH0FxiNn4ZweB5zlO7G
H5mjoyaaSBnLp3OEMG6a9htO3UfWYEkKOAZxkmQk1OuqU4cfOuRshA1nwmQI/X6M
oUsPDX0cU0gECULfylnqqrwD3ZO1+UuJNzZERbqCZlAMB/foggGEYfyn2MZBezHx
NY4lgftnCmCYSD9QXwlZ3czx8P12FRU748guxVyyk8bBjWevW4NDp8B4KZkfqOVd
7LXOQ7Bn0QH/qdpHgJiqT7jYR0Ibx8LpHHJwzmHrvJRFnN2IoZnf0sqoG8nvk8p2
TDz/8hpa1rWcLvtNTmxg7/PSS21QK31RNA9xtoe9AIzJXyVdWhSBie80QWA9NTIo
rSOR6OBlPFJW+U67p5YYe0qD3tjXFzpr0v5wdV7BJe3THsLrHsXXam1cJ7dqjFY1
hasNPFiylBRBUBpjrEy7hDIi8nhJ+Uqf1XmvqjvzWlV/9EBq6s1YswYeQUP8rmsC
x/0TH0mmOhrL0W3XUBTxMWUGj5k0tDVWFeqW8NPTFfugLQkiBFcAEN2K/TxtQ60r
org7RlVzR4E1BdTXyEGXJwAPNxE9Cd3bPZtDKq2mHbyg61pscHAejRR8fRbQ2LjK
plgUp9nDU3DrPOD6vUzTzR+rl8y0UwbaE5nlSZQKE/+LFVxv7p70CGMrmCoj6sPl
CmXGEjHxfKZVUOcJ05ZiVcd8uIc+rqm/ozPkiqHBenWmKts+gH8tqoX32Bwdx44M
Ce2dtlFzyt1FgZYJihRg89l4kn7MbQR/JuX0HFYdspVRydS96BHOtjVpurVzqkGX
5QvWO0F/xqxwVHtSYFBAK1JJrpLXJOh/T/GSjlidQXY7KXKYDgaAR+VB6GzWeV+O
FmR+kKiaPPoSKdWJh6pwU3KQkFak2WVLkCDosPRMW4X8O7mVwXI/xDPufbjZJ4HA
GWpnrRoEEmEi28cehKzkgYnwHSIMCQ3n+94mS5i9laTUGP7K8glRXWhwVl8dFyPB
mPHS2GSLeDzms5jx0ju6f+v+vOAxjsvmJ7gPqCszMZAEESlnUgQcIkCPmRvrmVxf
686fCUl4oX/BZ3G7CNyimQERHfcG9+NNbswyDr1KYTtUsZWhPED4SAQuDDKw+/OR
OsMpc4GVZYcXRfIIkRgLueMAKqtk2VCEhvJndr1zlWftLbOGxt4VGWqlEdaPk9QT
7tlWu8bHRxMQaCJzjAKx0GR1SRupVYs8wXeJ3N/7uXO287YTftfHDRmSqm4LEYMh
w6tEL4O7MQKAdIO4KB1AV1CpPR232+O/mte/taFhVIh3ILpc8MQbqRnY4PDvK9co
+UlmdbYKTK2/y23Ve+96EJmXA+Cdq8d6X+ayQxhoFYdU3+eiYSqGLUe/kSuHAk/y
ITXeWoJcYhBchVXcL1bjkXwHcKhICUGLpmSAn/1xdtZVgWSG5RVts0UgP3GwGmgO
CyDM1ltk+ot3SFhhGzQMYZmu3bF7hBaRkO1MXz6kxf362XhINbvXZPmop8+lixv0
aesGJ7w3NhvotdpR1TDPkw1wfPaJibDvfVrVoZdTlOGnFaY5A9deWekKaiUrG2BQ
8/vPAm9Ce1oq8qcCXChCRwotmZNMgmEeSiRgmbc1TxIQL63Ih243+wePIwJxyzU9
GUCdMG/lzZQ1Fn1BVtmwLMHI1TTyXnJbSOmle/En6fapQVqOnIthGHa9YVwyidmj
CW47eajU1j5LVkgzdMylYw79i5fitgksgHhVLR5RqMJTeZfeoxdq6vzanuqZPgMn
oIQJInhOCSzoxG+uAzyNXXw2QGLoI1q1hScW1J3E3T1UZDw2Kn/vwJkiqimx0dFx
q0Wa1OJrf0hgNPlVgW7yEvlvvwY8rDDedemdeDF1QDDc3u3aMj024kN5ieCdF6YO
ssVRLvZfzggn/2qflISF9vByTdvpb27xyJvth9gVfXinXEKjJK+LjOYk4Nvmy6u8
Qysf+BCEu2k4eI+1mFkdVrxXcmujXizevpGm5zHvb8ne5PwckhJwxgpq0op0kq+2
s/+FFeLwDJVf6ZTiXQhXOTrn2d2HoFeLLFhXYq52LYvOw+3YRawilf7nF90i1/dV
K1XVHUjoPkLr9dub2ad31O5AkENOvUkB9k1qMaPlu43ByhjDrLrJqFmCpq0UlRpr
le+K0wqNG3S2wfSPdwg6I4Mjg2uOB9RbTTqbbyjOgCNV+r2idRhfCLxMq+KPTUCo
TAS0UebfDwyGRufkvONHrAmLaciwsnRl3Ih3ZkY5UHyhdNCyX18fQUURe7yXGra0
7aj+DrhXYho8pO7wmAFymj3ZUBE1xeKbiGFCJttbp32pkHIu+Zwe00Oik3e7Lqeg
HJlJ+4nCpThKF0DpB9qehcn8aqFQugP4ILNzZJY416u6VEuqCpLIy6jo5QGFSPj0
0H/Oci1v8Z3C5PuPzzJR4CgZalhWA6bD8BXa2cTO140SGVHO9aFbRm6YyswsWI1H
1SKliBZsZUtbc8mEBYh3TzbQuZ1gLmglpS5ki1e7yJrAM4oVV8GlDPMb8P4oZlJE
AMfQvyAR6KzEgmOmnsPABNotIQFz+/SVOLpcdhUOGyPwSI8uTPFBbBif1bxx7VHF
7rG8cL4MnGduGfex3NEnzV/LVUHehE6+scQd/63tXGTYzTv0jhjdUjtzLAnSUATO
3DRpPfwvg8X8UCxSyFpasyKoyNtCmVG16lrJmx+bsi+X5/8XXWfWzwu3BLMRiaKN
x+LuE6IEEYGj7ryZt1ju1oQANtxjBVtudPK2QHHn4PZC4U0K6dBtGpLv/qGPUL6i
WLN/nDmRN8kJfbtnyqPLBRXYAZ0COiOdvsgkBjeHxNesidp6r4ei59YLNcUt2YkS
1yY1Wnvd8xJA37XkihL+sdaImFfUFkJT4v1/HvU0cZvyOacXi1bs3UgPaUhttNK3
F4fYkJI99OR3EJDfyu+AUNGTjrTCrcXQuBdVsk3coO2U3MkKK45H8C0Ryj6q0yxz
tjg0Q6DAnAaEP7mJSUep929Xew7Nuo8Zh00evvmjN/5ptjMnYcAi0bPLD3LrRdZo
DROTE3Ax0OBmn6bV5/WClq3NpXZiImJXzN7bX2NCa1diFEKFijrSxOz63hMe90mQ
rOFCT+ulmC1D8K+V4TiwRYzWMevdv/bCeQjSi0KMwUBTWDm11UXDI5m0eMc1mohZ
Fsw8JLDi3BcmZ7/KNV61W6wcwVcSYN2cM7Q2Hlhuffg8NrjpdXYR0/r3yUiS9Yt3
FQhK5uqKouI52Vp66plZYr6vzMNTJMThtzIfljgvvB9v3SMV/GKeP5rDuCQvFvDJ
i/xh1F4eDovAUzX0mu8KtCmK02mCdGyxtTdsxE6rwgr4gv3oUGp4jg/DnInhe93E
pCo8fVPhE5+yYxKkIW8NX8d4HKIDjHGk/yQrmDv6kcE8tX+zULSOt1cyrA3CWtKY
P5Yp4cEYlJLsCgMZms241oIsiNY4naa2Q1mmGym4d6VzetZxRIevR5YZm6/hBEpV
EjSnUTo3/QZNriS/EuTVOitUIbeQs2xuMSKjNi3NBaN15QD4REIjYF+Nqyb5cYhQ
vImAuJTUMlm8MoD20Me/aVSxE9/JLJFCOxVtheBcUOwl/KSFJ0kZkgsOj5vK2CMn
svJDD4KvFsVfc32Qwh8Yu2hCsS81PQTWwl9cfR/33FAKtVrmg9TYkglsKlbgLDxd
0kFfQnzz2Kfwe3ZuRX88awrYQDboVzNjJcnDCK0Hg3jmkHThRwTENYl9rzNPopPb
B766VEXQGHxr2j04be2h1D6euprRn7JwSq5LXndijouYyELKvjG3CfJaYC16DGIP
WjR1w9cuYMDsTAQRzZ7oXR/ZeQ6W3y0O0wScec7Zk0QCvsBwHSMqDncofwD2vHnJ
ej18kgP6ddbEDljCgdcigRRaCtN2PLNk3gklszskEvx8YYQdJFm9K6syLSCtbx6T
O/CRYFNYKv+XGKjeJVRrNk5e7YDLogT7dRDWU7BOFA56SG1wWKD6oy0UN2NDv/Jx
v2TxGis7tGOAbYSIVtO08fSzz3Ycrnm1VUZ03RnqPz+oJFHsBcxlGcHtkXVtRx0Y
oPM76Wmb1gZAVJbjYDynFk7GWp0LM0Pw0BLeJZvbdBMuiwxdfh5k6O5/cI/DWUpS
gxujsd8+/RdHz3FfXoyUp3DSmdTVaaC6cN3ZUXbFfrTmQy5eNnd3ty286Wrv7I0W
lv3vJ62Mg0zqcZdbolKnQBDKMC6as7a/E4c74X6c2rKPgzRJk4Lymdu4XxZBYTyR
rMplcJhDTDkyqjg6o5Ek2G3tXMRV2iLZbrqKg3NUenfE5rx3AkwBQ0j02m6OqFap
dRGBI7rAd3yPu5OlUHnhvNiJBwZ/tj2ZZ1L7WpuOoTxO8enmfSSetLDBIqK/Z3+R
cS6zHwAZU+8zcz9aexTEN1/3zeOVzu6C1/pnHNE1FBP3lvBawUxC88VAqtLDfPj5
zgmj3nz27Ur47OFbKCyVWT/PkyWniA722axy8n3On8cw1VwzxbqTuiZ2MU2L5vnq
nbBtVMIUeYNsOAP9N1I7CJyiZ3zyeze552MYRVa3AcXCj5V20f7i5E9tszRQt1ye
VuEJFM4J7PSJ4YzTlZS+DnR6u63dhhmKSh3j7pV4JnAhLCvddJjfmxGtaZoCsfnm
g/K9Awyj2lKOq49KO9hrnAY7HYUv1gprdo4yhU/BpkmtP9wk32goxd/sqUJ0k2sX
lJzeDVGR0gxdB00EQ2LUQbJhDaJeNlpUr9BWDX3xu3ea05F42Ez1BLdAMloISEaf
KTspdu1CJrBid10ZepORHxvMaDMYaYSNjiuT5z/NPzNDU0HjWZs5GSp5iGEZ6EBb
BVN71eM/0C/1bcMIUODpHlVXQE/9FfMZ+9hqBALTt0XhTk2txQPyPQhTm9qtBh3V
bQZCvCzy/hFp+oO/UzT9q3avJ/hKge0vxQZmm3IM8A6FtCouzwa8VIgVQYdUD9iX
8TEUT+Xa7aW/7jwrsascuwvX+Ijmfer6tYstWH04KpntQrmOo1e7O6wtXcQiYPXy
KjzeuCUXZyJo+hV5tzlzceG6fRPJ42oHKOszdGbl9uXOjYsV/sjm0LmS+7iXpfO+
/ZHkNx+rS10W8yKPqoojBEB1gcQMpIRzH95++JQlrmKC/Ipr61zu1KPxj/f4zLrm
WntdKxT9fRzAyJ2dNkFbtG323h0wPX5eUq/Ms5SYWTTK24DuOrU3Walwh9Ic2rh8
wH+CgAw95IERbUoXv9/VOgChp4tyXUgXyRU8k7n27grJdIqHUozeKrXDZz4r1mAo
P2brSAtE/04cBrHiE4m9cQWLy+1SyWhqe+e2Gnr1/M2JQ/3oc2j53yTYZpEuG7yj
bcHXJkN+OxMOTazjEu66OHwQyd6L8z628p3EtK5kS9e8v7VYHxFqQT4B5q1hRFid
ZcUvAigAuf+/3zzr6dqwGBuia2Di8SXn7XqjC9m+O4+soLcW8Ve77sjCDfdVL1S/
tZbI5Sd/avZOEKzN0gEtUKkC64smFeO6gJcq8BJGUnO+0Ib1S+H6HJw8GPCOhvB3
p8zZV4hpjx2s6IXj2QyneGmu3VMODPELWoig1VoVvYr8GJcL8DsiCywem4JHHOLc
y5005S9iC3H0Y1ZlFwSXoBQh1ve6TKdcSskzCeW6J3NHjZC9yeojUGrpmwp2RAHb
xdwFSXJ8aykAoj6qLfO3TudYAsQqZH3ACQg5ayg84nsAgPvSlPhGwlCyhmGytFgh
9ATnALTn3ws2bzxCt3y2qou+cuoYXpKhTvVHCZ4rWpDgWR5e1Ka+j/GEvXAyn+Fz
N3MwpUjQ7coNOtFyUxxgNyCS807NNh7ljfYuEf+1sosndj3x1fOQzdlpvdJjlova
MPU9fZAMiSD5POlonzNZ5zdwPcrSrpHYTEXk0pnDa6p6HUokzpfD6R0i2KAx8Nt8
2gJGW7nPocuyEhkcYnDM/4858fYpWYcvdGDxr5VggsVsy0v0hEd5GBL1zSzHkq4h
k5lj27hhMfryLrXyelU+8Z6zMo2B3BXzq1d/gUy2kBBupVs+w7ZSgN70aXbJMKMY
0j95epuDrJB+Jv+9E7kpN+6nqhOx1nP1m3YvEgqSBh0SNS8ikCSSX5m91fzOHKQk
Z9VN45rS3aKBkj2qAnez3sjDchim9THwnUlBfDFat2J5tvuDYP1LvR3RR8Y6NZDI
LmI9x0TMb+hJoA+c5zfdyJ1Cpne2OTQsPjIZzzyYW7yfl993qEW74NqpkSuwE8jV
mpeLqeNwdiovkuB6XtfOJtuk8E99wjehm1R9W4gsCVaG9nM7Ic81IwjneIJ9Bo15
lLU1XvolJ0gWoWH1C3xVFdINN5Qa5VcNJWfSkSlt5ZEsnDD7qmc/PBU/NFc0TKEx
arzmjgrPo0c3ghJU5cD0cRkokdxVUzml5deAoiwawfQLCdL4SsV54CU990Qpbn2l
yg2Qws5OsVhv/xr5n/U/lVGR/IuEKdqigSWWIGfbc/W2EG/N7eMTGAA5ulcHSqKX
8QPjJdT/HSzUsAysHhgB97qiBnxjs+L1+ztPR3oL80NDfnVUTwl21IYlv3xmUvVk
rZDDwictG38OftSQJgX+wl2bpfMMD1LaBcmn59kKNXAOa7KJS8705R7zf1pDBsZR
gFg+GYPYhn/Q22qLmlVmDcINdWyUwcRMYjunesGfGsRhpCVolUPjAILRuScEMQKQ
gHowh61JRc5kZqlmM902I3aHPIA6J5iF48bq1fNptUvyVMDIZryqlRgSNL9aCYt0
op74iGF5zv+n3S7QUdRcS3l9hpO3NlGKRSkJnMFaQ1aPkp+1FaARP1ezmoorXx1j
GqHTKwtSD3WeUZ0DUe93/H1HwsqR1aEUZCYGEJDDSRvqMQBkCz8yMtyV6h7qYic+
8ZDYiGMlN4h7LoO8VvAf0H2ttQcj535mpN9drSmpJTtUoBVX+6c5CO/JbSNKTbHt
i0ZdqfvQnSKsKVtz5pXSa+c00uA9iV2zViGN5DSrjzBQHDzz9FWyxTp4AG/FLtcj
PcjSnaGzhYHb6RroksYdraiocn51qsiltHGsgTGU0JFSAU1IYMz+LLoffd81vka/
uMV8H/uhl9ZI16p1egWEeWXXX5kStcasJOK02espmRS9LG27gsK2aHpO2Z8jdetR
my7mr24VVXU7ZaLO4m/E80hxdFcyrr6z9KVfV99swHW5s+HeLRyKQ8Y4Es0E3ySm
EoxrcEY/vQj8vuod5Jrn5yagwobzy7nlCmIRgEBgrBSP5FJSmImLo3ovngU1E7md
DmgS388rMu7Q2bgBXHsGe1e15ugD3KUTq5bo0O27G1ShYg2vRr47OnA1pP+TQn+H
nzzwbqP6Ooy6WwNimXmpTyMw6TubA+I8epU07VyQ0KCCvEwAMy7lV4r3ODBMJRzl
wQ6+W7kvbXMuYUnRFmo+Wxpu2G5xzDeVmz9gNUdolJFvW0Nvr+ASt2WV0LqAtUav
CbBqdbxMjzL7qnXpVeYK/2uRdI3TID195a4Dtu2CsEnH6BonQG+VKeBSstrLb/W0
u0lfDx8lNHLqBSJmeCOE5rPlDMH5YkupQo0Tm/M4r1UkDwgI+P+ztiCfuidht1do
X8lqzsPsPoQEMOjeITyXswW2UH/Md4Q5bzLB4MY0K19Iv+P2tkpt5M8weXq6+Y36
hZXFf48aKyZ2scd+NPo/roQmbjXCvjf2pK5rXXfRuFz+C+fglsTAWxNPaaTV2N06
6dVw+AJpkwWqpWyxSQr87nKBBVjSqrjHOoQl8QGFGffhMPT3I81MWnZ1DtXfmHih
5qdL7/TEBb9F96w2fdoIyIIcv6Jbv0IFIXqv1gdTGlRyJitqXGUPhJxWxtXZGnOy
s3mMFaJwtLIJhj6cxx1jhI9TmKUtvG5qUCc0Ck8gqTpTb94/Sy7Hv+yG8+7dQNgF
CzQmNFO0TbiZ9sKtlESCXZCxgGIDVEvaeGk4TKJcanz1sKru1p8J41QP2k8tzxhU
oItE+nUNvDKyEXd61zRFWxNlR+ZTm1tBaEpLkq/If/zaNWSwQovPGUkdJHJWrWhd
w9cDzkm/Kq3vgicxVPICJZxU9KxR7KYB/HzsinnwSJW4rwoqxPF3d7tk8NhrbCTX
TJy1yhEfTQvVPHybEvnTzxXCLjyvs0LZsaxuhsLEw9ZyO12fRDrFxzvaj5R7I+6y
tMUce2slzNB5Sjz3j3hWPHsjT3rJALREOIZmlJbWSzeG08+qvsrRkUYsKgBkUCyk
Oy5a1t5RiIIeJSOpWFX/XriOQDlclzSwAqclPj6kEs36TYl1kG4kF5228yj+ltgR
8oQK9AxavQMIkNgHFV9Ws21uZk6VLqGzNpAmXa38W+k81q1AR2YlJMevtusXrkrA
xB7sT3O2SMVMsdP+cl2FPR1km2xPLF08zOosD7Ay3cMbwZYwURNR23nUECLbUGne
C9syp/HJBHWKrUW+6NHqB76LspmRDLUK/TK3kowhrAk7Fshmt+KoV7gWk68zOihZ
SsIA1LYXGhsZzUDQSDrfNCrhzE+toRdZ2f1kHAQbhGI8a0j9e67tgXrwyiaxd50p
3i54LvGPJG0VODPp07rLWabCV1l73U2V+9R6ZaXIziCREL1J+YsCRT4+lnSrR0jH
4Xe36p74AHNVcADGiSgoq2M8s+dtAokJynafFfsNarUX8WSIGoFXH4doYGb+g33H
C5zydGwC2m6mf3tQipgia38zcv+nXShGj0eRQb6lTeAN1+km1ySoruM3PLQbI57j
qYEyue9xJhSf15r0xPwRE+CVMorWw0jKz9exdR+/Chl7voDYQ4UbHkC6jMPcUYzo
+rzbCZixm6/xdpG2+AkLE93wnfwebTtNhJXMJ603Ow7+A4DXFRmRkdTTWtwyASOn
AKxQww0BI36im32PgcP8H9O8vR6OWnTQWwKECO+AmqAqqYBzNSWaiG/bN0/S3YzZ
ksU5BhmV9uRSmFa47xOD2GPCe50fgbJ3suK3BUeI0C97dLaLALVlxzvQNPcK+LMg
F+V2UETr4D9w4mXYcJJGL001tRjFDIV/7XclTyOZFYlqH2g1XVsGKAUAZKFXXtqV
pmPyP6YZ6hT/640kiw41x3qH/pWKuWD5r+QOjBogwF/fT9MH+kCgv5Xiwe8tGM9W
iIzkCsQMbDYADQpQY3aB8BLnKfP/QhbT3aPWqs01do3sjcyq5F5UBRetqP6Y3YUL
SazvT01690MgCwy8QAPltoV/OcfqhXSgUQvX2zPUlz1NaAOhDnZVNFYVk19a38pO
5k5HutbRAYCSJkbNwFPpMBJ5ws4Ljipd4PPUXVdoin7bU8ARpqE0W1NgjNjgLbiQ
mUKO6UqCr3xcAaoH+vypQoBB35vAw9IGTjfAWRx1BaWTEDZ1fWXlNd/KoblgUM9r
frEnyOQ0irshG/UjKW/FPS6RyDVQWQLmp+m41GSZPeSMllPOuJUONEE29ryX3edA
CNufEeEabxbgoq0Pw6dEv5B/v+iEykUfqJ++Ps2TkVQ5FpuaV+RRqwODTsOOCCB4
wg5pj7qU9ROWS+qZY1rdhWoAxn7o7wY4FL8pa5D3PmTbeLRuEbJXR5TXyI+DWyQU
iF/WUWB0my0rMAj3FQI22aIaLnkskX++DLYDpxBTOvV0inWkqTJLJLjDU6UVl0Fe
tdfH9/BhWMc/IO2KhyhAtY2wK32/QI1a9tDEkm7gnNp5NgtAUgwbD6VCHwQOMZbq
lkJY7EjfhVuN69Oy5jNcsnd+j5+xMS4N1NglWYcWMqDScMhYwbSe2rMBX4i8iGOp
mRaiTV2UrH6HkyTsSZ17gmjdcHDm56GfXNyeSwd+P8QcqasLugdoYwwKlTc3tC/o
ilGHNT6Yd5IKUfD24DUwMWwZhSpJ5gAXif0dqzUN8qBFG2D+y1MsJJD8FN23WOXW
Ev3hac9TkRy6WZiAQ02fb29O6H9xnQwTWjfnWS6T0lqae+ynIynJ+uMwjbrhAt2N
j9WSKGZoUBXUIzcQPzuzAZLNcczNzGe7jJ4MPelglMY8byhk7XGpgElSjMz2nw8v
QtQP1k1cEghVZaboqP7FpahNdnhLR6LIGyDB5IJqPTgTVSGisgX64Pt+LY0V/lSe
aVYyTI2AbN+ZI3OURumG0dMiyPeS2KKc0FhOdDfyrskWgnAalRecbPp7TJQmqz3h
90I6AkMVxKcIniJGxqFDWttic/qS1a28uYIrKqjJu0Vij1IBtrjCtqvdVTcY9eXw
HD/fE4R+fRuOK0yLfesebQu3KJJS+IN7jWQ1eFYZbLpdsWcc2h7Qj/rMq4OieuwJ
wIKnmlix/O/KriJYAw/QdhxmoE2B4apcJ6We20Xkx+dtP/sEws+Kudoh8NVS8/R2
1eLnqv9bE0WydX6izMhjmEfoB7+3fXESzpbdsa4o944aLXOxWhCuVpQQYx943ehp
1zUXSWgZyGJV4KF0TGbFSNvYwCB5xFxLUpqg08/AKP7fUCfTkEyCJbppMLgyfpKb
y8FcFHTbB8rAomiabCzHygtcE2jAcM+iDNAwEpgBxEXP06BCvl/i9TqSSi3S5sqa
PoD75a4kdlFVe9XXB9GWRLfW36ncdTXMXu4r46Q/HQ13+sRK/eD8MUszM+HKmF11
Sz6V8oQARqxWMu2fTbZfp/DZykE8HqolwlLhBCkLjGMTJoyknh0BoQm1vBsFu5CG
b3QE2nejL4HSgxpmVVyFbTLT57rYpdZk+UrHL036KV5X5smlxBY4XQMpEsiFleeJ
U17lDPocuJ68qz4Cx6PStStfIcEsVcdoJtucsLX46X4/o5Qx9wVssYPgBfoI9o3k
4qQE4pISwsv7o6+QBJOdQ1nLAW5zhKPWUwQH7noeyWJtC0qmRB2zmImaHwM47q81
9W0cIMNjdb9ftYoIrAc2lvkQEwj6Oe6jmDPAgARo0KzuTPie6vz63aH1XhT0l21K
kdd22hB5jcOznHH0O0Bh/BHs16eN7KPYjIH+YaN0YvzDkZnh606Pq/FVJgfqoG/i
MaDA4olB5PoHS7Po2zUOmZKj5poDnTQAgGCdzjuaASK1gp2ss6u3Q36J5jRulI6b
yYTxSZLUjcOzvw6vTIP7jCPgH6qMnU8yQnKO/FDEj0L/JenGejthYOlGw7hsI71f
4pl3wMd3zFXhI5PRSnFyU+9QFbcbG11SJfFY7YdCncpLicSEfbpywdix+0GdOROZ
h91k97DXY8PeHBSk03ro0Y1JKxuB1umzxrwAc3Ag/Dv+ie4Y5lr2RVCEFqwRuGgn
by4SsOUzU2OZCb+r/oEhjXiznYoCBTHdfs0pk3aA2fu8v0Ysu97VaPQ1C7bSoA2g
F0ONx/tLll12C0mgCRv96qQldDEM7F6YCcfnInXqketa92QRvcw9rALfODP72BmD
tdr4/bUS0dPuS9vn8VkBH7bcqmYcmxvNiDG0TmWUIXsQLmJiB0MRSyDMJIiZu8hv
CA6lxbZUKvyjnUSGijKrJHxhTH+prY/4V8O703ga4Offeu6fp7ta9uXzVh1AeCRw
4vNm0QoXEMiNGQjQO+vzPusGaemxxzqh7xOisqE12mno5ERgViQZTHV6l/oJFEbR
2V1RweT8bY8QhTJwxvMJOUWylYpjE5roA7Tn5t54p+nTUvXhGmv+NQfQKLpN8MVs
jP3b6+ORPGXYeB37XkyFQmhApyBOIkULOFzMC1i3HLdCClQFqrALmJeszqlLa5BG
a8kIfAEMJTsSueZdtbTiIgdvn+O0X7XgYzBD8BNl8SB4tMpGuGai1d+i8M0nVcNb
V1IZbpmuezgA0pjAz5NcNVdxw5/hOVf2QaoK+OIuQ0R8tQqCTkSyAXdewrm7iFps
WrMDcgXqwLuujB9dtFiAusMgmdyC9KA1nqB56ZKKfYaaASruah45dgMrhRAs9VmI
/BLomyKL0xd8e0anTSKf4O0kHVfJy/p4tXMd4eHrr4Qgcy49mG0cZP9p/82fEsFq
3C9Yn13nOihEaCOv1oqOZZ5K/KJl/VKCv6ggV8C/GkyYygy9mqqeBLY3Q1sWZW0Y
zz4SJNJ2aTFYVNJy3rQc6+ktRYSpQLS/kb7dqhVuvLStzAoTVr0FKjQMNfEYfBdJ
NtYTrcFCPqvd5hxIIUa0eOAR1GCNCK1pUuhN/cfgyG0OyF9RWQObYo3N2nQJiYfq
gBTaBqVyc1hcG2ckXi7x3bryppwuE+Z8Lb7cA20JhIGEXvLVa32kJsQ+6Ew7Ff9a
IyNajK4km4C3YISmPclklGd++hshg0M2z8lz3QgRh7kqC9LRvqvSNEbJYRJVENYw
+a2XWSq3MdnrpKDqFzb3oiK9NseejzBNySd6DMcp4Fhh0s+ntkUhjbNwh0IX8ryo
fWf19Zbsw56DKs+mmcCLRLrMfqMY66paKlySHzfdVMd2rnhVb7BGKPeVlAZvUIDS
JiWjQ+5NTwktXQKXktmPVALfAQrRQLuJWFYfRXAab7Jgc37cDoSbwybEFYDN4+XB
x+4KWs6+tA0xvv8p0w3vEIKxVl6atVpG1/dCgDe5hLUqWXMkicObUfwb7jit5cVw
tNtaIHNS32v8e5mWF2UBlQysmRpIa0jAFobiNgeyouPLNz804GIpXOsl9KIN+u4S
EMSNdlKGne/lmWnzhd21ayrqqjPTvSYBhBj3eT2i68gFAYKstAX2S/pzGu4UY8X/
6b2P8T64eFHZsmfPdux7hLcCAHq9NqrJxGMTt9AgqAeF5EPcmXYHcoXfEl9WXbNg
26PL7WAK8RfgnXD8phLjjWKze7Eg2NCrzi4W5kXHGRUbb4fHpiEP4liugkFqJpAT
3T35dSoeS8eT3njr1z29nS1pLbNsgwBRFkpC/7zD9LRkNbxO3A5tinSdGhQ80Vu5
DHhwevjyhKAu5F0NiqRyf2Vn1+pwAkB+hAH/ChBv5E2zITiGSV4TnLdW4kczIBFT
011PkeNaVZClQxn1A8D5CcwEnNCETj3ihop+KG38raOyqMrgLopxY1KKEizFhJ2T
KQfenbbWdEuFOFKmoSfup8sr8AiSZceKjkvTq/e/MotUrnYw3/uVJgX2Mo6o+u8f
vlqUdxZlWSeRpaakMJ2/qNbpWl2ZA4M8GyPz7fNcLQzM4/4cqN20SqfpEx2qJJRL
qpFveSZoxCUbya9O69PVZNMDvatr+rCAP9xyqzRUAb6mEMh3bqT76qpuUVXUlGdv
092rIh/SS7K22cPofxzPmMb/yJxDDKOgjY7oqKa4YM2xoYJjnAz7kc+2d/sDMNyL
jiUxkwnA0YO+aB4nwSgnALKiPYlk6Y8+jBflGZCl6HVDfXPNCzuw1ZMbul74kPnO
CFl2/qG4+ypLMCd8394PUv8nrPQwEWe8T1ktDyUsngH9omBbLDJoaGOqpmHjcQGj
3/ZYrIHWNnFX8XhcCg11WodMb2OdvdrGyYGeyVRT5/zkQsCFcL4GE3aNajQZaVFr
C6NBtWzKBF545DSC6w+RL8MY+3MD9cJtAJvCvOqkgaJ5ljvkoADxR4ybeCanfAt3
sJby3Imz22HZLtwK1eA7zW5wbH4qO+t+o2C4KVhG9JSkB2D6S4riEQpkPLmOXcZj
q1qx3WPY2PZtDYd5DeBt28EhhPuCxD+u8a8aWXKCQuOXU93JIpL4zibzjmtyxORt
xga/Z5TwOwlR6+qnYdKM9qPOq2IQp/Cb5iald9VrG+SBT2eTFJFhcOQjilYZ1eTa
R5KoyUP3/sTx6N4S2W8bqIdn94L+D+w+P05RoZe+zJLJ+dIGhvMmMBbKQrLL6akg
HMLJ8ibe7BJgeQT2dQ+DzlnP4tjuwoaf6KnSaI+QvBdKvq5vPm3V0ZTpnWzL+KkT
dVowOdnd4nCkGR0jWBeid9Wev+Am6uFHBPFB5+/RjtqzxSlaoT/iosN/0FxGDj4u
I1vsLPjkx2HiksjpMbSMOXi226s0MIH9JM+K1TM1WzcpklBblSx85Ah3y5JtjMGa
/nMrdJXawKJQbuzGcRkNwqx8ohboTwq/h938ppOtoJJD7q06xFU949FEtkjmtRzw
gwjjwlahNjtuBqj2ZWc/Xpizs8vtfWJciPLsoRa54bjURAIZjlLYwOBOibmIe+xH
EFLP0EKUoVyJFiczVXgrRRREws53B8o18Cu8+90LUYAp9InUdE/XL/xPPFfC5INx
K7jX90Grk8y/V2Ir2jHHqjAKBjU/lm5t5TM+s9by/QdVa5QMAEQt8bdyjr/mz0Vz
VJK+6iNFn695BwXJGY4px4WS94pKqGGu5mTxj6IKEv4OGfVfZSqL0/EKcf3NvD/s
lEJ50C4U80meyLZ4QlqJo7XZGvxjsluysG9F9og81c8h1XYoDvyDdHXUG2jDwVZx
diFCyql64n3JUIwbCegdb5wVjaigtBFEXSJ0m/i1flWQtL0SEHdlMbuEh2ZwuGNh
Csma7KjZ6p7c3O4YgfQ3J4XBMf+Hplb+rcWVDZuT1IqODO2eh6wk42YPmVrOEQnE
huu+dRvUl+wbqTtS1zwWmS+zQP9oNUZhi3qzLsQG40/j+4f16nNmtG4P3PJFaJvd
8wTDMEFbmQosaI0z8mck6ISCwuNsojgRQCGpYXwXkDfXmvBzjpkGMMHz60IJQNvL
/zRVao+/i3/25lTxkSgZiaOG2nl9Ii3Wj4750Wq594Rqdlirbi+B4Oq8pJqIU2y5
mZT8wjOfUrUbp/ojpm5gXluF/6MAOW7T2BLfKIn2MCJgdJzvZT96g8R8K2GwX18L
49w2PFlqkIM6uwUeo6UoNNpz2cYesZS7wltDmwH9cjJrlhaITL4KcjPxldiuwAX4
de7kppj9KXkEy5Q55Bp2bWYKd4gokzyVtgVOAUjCemNpg3ESxdMGsRjLYt4E/sZx
/sWqp+JpyEiZ3yINniWG68PZtuMXkLXsAoCT7a0ZgqlZSbI/JPPCiV8B2gP9zeOD
2e5WRw/p564uDc+n6DKjQc3+c9PSRwta3Tm1VcaYmsnaLB5FyjKFdRVfthZGBVHi
lGLwpODrTw7m4JWNtHSWd3VvUESMnl2lFRqW5T2+OnNbAXJGu5cwobOMFpfnNBIw
7QAX5h7KyOIQ5C/vdASFgSOZ5Bc56jpcZsr945o06aQD0+beilR38Ax5KS0Di2lO
uQsLaUQsoghu5WFRkvB5nvKAD2TCki6VzZ7BGG2eCnoiuWCEnKyocIvmkl0wQuDC
4gM5y9O1XrP3s3w5nO75rQcBzywfjpaxO5ThcfX8Ovnpu5w1rhS9i6JAxIdRzWh1
btG0quvXhnPm6re/pJSb5yvfNfv/9KuwxMF/Px4i2EpCtj5Lte0fCnrgYEgUmHZj
OR9BsrA0kb7NhvEjjP2FuCP17n5DrHaGNP/L8C13SrBkGxGFak6fznSmU45Dr51e
iVG3rMFRjDchRWfFfB9Y/SHKf80i0GJwA+WX/tTbYyB2BUmAG2MMWMRsN3rk9TZ+
9WCbaO663LO+lj4O/dE/W/jqId6uwI9REgYwNPK+10OnmmXRMAifseCQDu0ITk+M
Ub8RMO4LuhZ5OBse5eYDv7XNPss4oYeeHL4Fx+IGTpUUtRkUKpLv+xNlaf7Ze01J
5eQHp1zWLmnSZjptk+f8epN20A3QmSw4AmAvlVDSUUKDewO4/dC3xpH01kMqcDG5
4neJOY/lpqMadVZ5/FGLBOaUasyAFoO5iJINxJd2UNIylvlSjN7FYXP9l9Av3iDt
A5HwnCWkZ7e0woRgVrSTGaGJy0AXdYhYhS+qWoXMIwJhMkZ5Cmtq60XInPC+LETA
4aFJOmVvc4p1q1XuqKOkivsVJY8gjwZmz8HSLmy5UPWoVCB9GXCwKn4q3CABAzzb
pQcSZPOqOrlh/79aBEJHzfKsfyyN9Q3+Py8Sd9BpfvTExhUQ3ShZxM77S3X5kFIw
WWTKr5j33r6G9nAIQNMwXuDlk4EK6MroSgPaSnzYUZZApoOosdsY7EbVyYMQl7/E
iX1c3ZPWHI24WA+bFCNdWaY6x1N7JPq5tBfm4E43WckCfheMDHJFwBnGg3cqd/tX
HjDS7TgLBq6ayUhUYajTeFCx/mwkGQJ1+w/4J+lk3ngS/TTkEVnmZhOiphNsShVK
qWfWf/LupwcX6yO9BqALwt5idrB1JiVJaXdnsvPo4qCU2zx+/DO3/WB4/66eEXSq
uLN7GOZT1EbtpoclIqq3vC/QY1kUqjl/31cq8qQjVVvDHeKvwhdhWTxya0KKoLP4
gH4mBAs6Bk9G/zlwvuqtJevosLum3KPL11UKDwBdQNh6duk+MNk6gSexu0fMtD28
bCwA6UEC7JYChWxpM+f5XX8N00LrW6v0NfQq9DUKCeWNFtz4IgfZDeUD3wO056nr
Co97/4W9xo1X/fpozkQR0tjvFslyQTltolfkeGLBVmHei5GqjuGyOtAJWNkMQpD2
mVWaKK1LqtstoUI6KRBzyteY///0gwvJz3rSixa31TBILfOJvrMklkwk/kh9meie
NZPoaHZry5vyu2d4P09YGb+AxKb2wzE/ghBAUwjlsskM9SChbqKVJI/UtBN+3okV
XPUzqTw238bN2Eh6/r/FXUssbpu/vAlahVKQD/hya4zz7Av0J3EK6+zhX7ybHy0Y
5E2ynpMlRtvTQGk0++EdGpu67chAxxIN7swcW8HDPoU6/h5F0ZRZs2oqKCodYeGC
4JIfdGRGoMoZNG8Oavwk0VeX3mS6CJvifHqYHO95oUHRJp3Cu+W+IPhVTs0j9IuJ
s7IOddYhuN+UMLgPsf8EY2JpNF7CnaYQoJOliHVnbkh4njZwvUSPjgalHTLLTWS3
8ouCI+eU4cCWw8fRytQPetYhovFyR3zVVrshbCh2GQenZu6PmeMIOirZHDvMuR1N
aHuFlrw0IwPE/hlqJTSp/Q5Z4o5ThjP9/YNsqjPd0C1tFUAX4tr1EVDizXM6ak0D
20Fqan57e9xfIMiqBn0QBUQ18TOAtObgiE8jtzX881K78//g3iisSZ0C3yR+bDHe
jOEVq/HvCGy2SOWJi/OR5f2kBi2CjnpVUPnWva7XRtS5iBcTvF/GNchS+CTBD5Xx
7mn6p/XaUqILXGfqpbrMHU0PebOBtUYraYOTo0ANKxmwF5xMAvuqv3CtUWqzKpmw
M7EIAmgXDlBuY/VEVUo0PpvdWOIAAHPzYNhkLjP/ZSLLTA3vg8IPsSmCi+KqdENz
2itocv0vlW/EvddmUV2V+wJZtJ55e8fuSAedJAgbBG2yylkrNTdzC27UhfG4mqBQ
S7RW/VbVyOMuoq+LTwgyZhBSf5gqDPDt+yLaZc4WfxH82LM8EGMYhtkTOtJC/B0U
XoIBXJgdSSMasE7v9m+4LAEAtZYb6JpJSxFC7fKNzM8W/9OxNjFITQ3A7joi5pYl
y1cwrmerRqgd8fzn9W+karJMT1YQSGgIbmMrWO8ZtJHMbSRQ6LSvZp/FRg2tSr4A
16/oWNLOB5tsaGdfcltP/IeIKeBdcuaXTcKiYGK4VzQCtlyZg2+79u0gsYHk2BLq
wMmh8xh9li9nq76RdzQWmznbUszRgRbirnitGP4mJ5tKpjoLJVt2WpXhozRNRQaI
u+RDz8DWe5p/xEUq5zb7DireGynTbNm1qitiMHJdmIjz8xtgkGLZ7UybBxmzzBTL
wwRi8wkBQVCAeJvHVMRdPsqHqEfG08nHZYItr5vfmG9eNcVBTxa8ynm3X4EI5lSr
96lv++w/JuIobj+4hr1KzSX7QAtjkfdENezNFhc1Sciv3ZgqTNsRokTEAb7N6Rvi
q4rkEVXC0vx5E3adJNrFhgp9xQ93D/kvy2oOlucDM9SDVywIm8PKb2yzy8SwIzl1
hfoIbYoEzsJgfp97t0X6RdEZF/gz03ZPIE5uovGlHp+RuM01FLte0mbx15SuQEl2
XRyY3l9ezrnP/eeNz6oDqnjidOauni6aJ9WNZmIeCMr0a91tpD2QWM23W4CG8TTE
sOkjhdt1VMNUf3P0w91b9tX+F5OFE6o0FqZmt0PheQTx4MZ9wyLF3T5j7M4LiQnH
aEj5YU4Y0rJ9ZJROi3lbwfqflLyqAGyTtXP7R2KDCYWkE1DmvjYalBi+Lj9IxN3r
NGAi3B0Rol8SaKnxt4VaHQtXZmutKXhCOj19n9ehDZLwQOWbEzFDNnCBr8q9+lLP
qoJtFKUbF+h4RCSPIQQ5L/Ks4EiLUsdvjlB6hyPYw1NPDO2A7QVxo+MWnkgkqe9y
S8hqjRbgksDuJneu3zpKvLmtuW1SxxupfyJzWNx1/1+xfQqeFIalgxB9uvUJcwiJ
l5WGe9llnD01GfxxKWU8dajmMOosExmyasSuBO9GryPph4X+GEk+BfLpX7P/vAMA
tCbS0ImPn0Je61uuJWbKcg/xB1SIjOaqxINg5CAT4F5cGHJY8rskYPyGw66bE3Nl
/cDGBYB1ge8AUBAKGJtza+ylIxkJAY/phuaH8HW3F1KUWxSYGHHayBE1kwWGzaSD
qjgBg8kS7qesRcWw8xGLKBC8pCIYTlcy3qzPfhLuKBsV8epVeaWp/WjdOaDWNMWf
PVySvDFDKNih+9KIOk2XQayP3APC0EUeTVPbEkFoUW9Sp2Ic8ykl41VW/WDvwxSU
xdbAa0vf5PEvSirCtWzW2CzKRyCVtjMXjwS9NYxSYV0KgG8rH1/qj0Dj5yECUSbR
XxaLWJ612xwO7nwf3j4MHSkRHFUe5iCC7/g0/Y/EdLS6Vuc0uBPcZ3PC1Xj79i+c
L3bAA7PUGKBWCwMy8NhCHEI1o6x2w+m6UPr8LQMjvnwIWKtOD/u6+uYGJWWXV6ze
cGP+UdDUNvFHuzpGcjLSwcy8k7/hYWZxEY0jOI41jSdoLF4Hr0RRb1VHVozil9gp
h9/dwPrep2W14ccNYsxmzdnasvHC9ZT80IhWtnhGWzc6KSzvocDsGGv41neMn9FS
oxToaYECb8yZHkA48eNKGeXsnoEuMWKXpQftQiu9G5qMcGrhdar1WUcJxG8MFfqy
R8Gr1+DZo3mrqw13oyIQU50mX6RDy/uuR4YuYbVr2CZX27GOdZ8Oqp2oEW+6hEv8
/DLINGcmt0iMze0G/uKdzbWg5lwibNuCge8z8hXo4ojPNCIbRNLlGidx4zZuulJb
luIKMAnY+7k0Xkxw+kOuSuqYwMTbVbHogXpm8X89Ps9udNklEiigmXUuOphI1WMj
5dMFwi00Omyt/6FA1shkABjiPR2RFU1lB9E3KvnfOFV9F6BwITeiE/K4pNbgUOnB
OSp8ncvcFhTa/7zt0DIllFtXSoVLE0F7uLRw2V+d0JDkeJse6YTelnIyH1LBVP7z
TugCDy5ybeiuu4JZtkP2NQfq+Pi1wGifJlXAECdHs8H7poT6R/HKT+1YAlge6j11
IjviQsa5wy/x4GVkWq2ColXBB9Xlc3y5qslMX5s1NhgoiSKh0mZqYVbGUxK0QB3h
I6eub8/vmM+36yEmNP6zU6MOOpfbyVeqruYOhifiU+yg3aMUcqK8zpUOgZHWMHf9
fxBn/6al0In30h9s+qBY/OqIhafcZUtUT3zAf8MHIwApNCzrNGcXV14H+76xMyVd
x28EVKIJxodNHL2goWwtblIlmkEftETG8R7RWlkTKw6560OLLY91ZjioOeJ9HHDm
JRYaeE1WDQcdwuiAu0mtPgKYUtI67yLFKwBsfQodU4YNRAU7xzUv/sgfIG7O5eT7
7XYERSsnJQoi8SFaby+VqOcSdJRo66XsUTdgjKytpPCmZGGY/QjkqOPQ33P8H8Gc
yxmRe3XAdvCdQpS9aomd2ygkkPBnC+NvjPnZpvRpoS2aDE8JG4kXDuahBFGonSVO
19kgTout2EsJFZNHKdWTDqERclVDhuUyhwPWXMFkxhoD2eh0IKstQZT/bGkSk2PX
va9M9iXVGnhjIceMuLYJfyrKQZl5ya/sCPiJABkI+KmnU76Gb3Iybj6H2UMYum/w
kU54NeboucRqEm1fEjUn6KPjcuQCNU8hPbDqcZ+WU3eB3oM37ZHzFN2uKfuigG3N
KserO/cDFgCw9GE203oSDONBYEFVYhTcfojz4iI0xLZSg36KDMZsn8bbPYrdAd1f
VmoZukr153Befd6YXZs8fx2OBwZJ4a9HcU7Oj92x7JougXIkv8sf36Eq0J0ezxbX
yOogm/viHIx4BIzSFvKfaxiZw931/uhW8KOkv18UeLhS0l9dAVp7nqWq98majVp8
IKO4rBEw5giuBGXiKbvcUY3lMbFSx0m1Dq7DPr0a0cuGyeGDH4USL2G07BUDq2Ai
NLr9pJ2qJ+9SI4AI8TB6FMHrOp9F5aJYWP6KtTY/InhRdQ7jCMQlVsDwIW86qxWC
TIGcbim+7azKeKM4ipNYfhd9Rdf9wbMBkAHuX0YkoKFM5Cso3IHaLRJj28Y+Ha30
xGU4EPYUpFcJC8MU4Fr5LiSq2P3XaQYhbHIRnjdrlrSv/yNXE5pMojf5ckO5+wqt
KQjwXGVAqgW9sebj7SBuLbMTEgTJFhpZNyFIYNMZvPdWX06Qz6cQVe7s9g+ULJsm
fHk5Gt0nhbbgbUhyPj2nR4asm5SLW9j/tSIs4wlk0H7fBv3v9ZCX2TEjFeYIzqqG
YsH9IUiu82EVIob+uOIXqOLRa0cHZYzsiMJcdNiqxy5RnKISYhSmta1Bz8p+Jo20
Au9VmgTwFEoYPESyJHXjudLeEdyWcmDgSdnmg4oPTpEZpbznHL+rMR59P27ypU90
lRx612hncF7otqKzSbBLGuE2u3Zsw7GQnAUCMs4J/OEdeGMkZynLBiotpYkoaek4
J9YTcOqzXWYg5JQvANPxf1eqCiItws9Pi8A4iNN1TkUQNMDi9qXM0t/1qD7u5Eeg
6xx4EvWMYnw4jxwJjrac3d5pwwTj14XT5sRA5QC7iOi1gmJRujDeN+DBW27Swwd4
JMnTDJZJgy6QhUBjZOGYxcLxh472cb/o3UITjHmR+4r3EfH2FhPr5wZMxBG270TJ
SOB1blworDSmANAP8m3Mr1DE38Y8ujlecrExC0BhDe9ejZROo588KB4G08fJKOrr
J7VULTa00OpJV06lZLtNJxkqDQ+l26jVRsZSLFQFxmql1kJPs2cLb6ZqZkvlbO+L
rlzvEMmLl5c332u/qdbIs8x2Dnc3EeBl5P9KudT0wbOn+nhZo3jYDmmA7CAEv6yu
ZtM/38s2KUrJrxtfMdg7WVKHDcCfqTlFXXdeO2g9sF4id86Mk5fe25PV6b81+HIR
rsD2NTVd1mpkaBU9nQ0/f3Nw8z0CMFtcQQn90bSQ6glnvZCKOHpnXBoxEo2Ol2jU
NkcFd1TmGDB8MpvfT1emReNlGFlyng2lVjMxJuekZbLuzOO1AQxK5w1akylqIeFV
Xz2m0OYO4YXh1nyHSeVuopbzRQktPDYAoo6skZAMbUSzK6OwkqUEG3jqUEMPs14y
n7B/Jt1EhU2conWsqdVei5Ha9iBWKvb9olNwD5FMJmIPpZRAvgGrsyH1KT/H7eMD
Rg1FK7My4U4sjCWjsPVwQX9q2AiOWCI4opk+UcbXSgTPfp+Bqh5kqMX3fkNLJDUx
8cXfrbW2bBR1YeZvi8dYF1igrvYK0ROGM7kU1IVLB6CIWF/QQelMUyge13CdPN2K
HaOHbex8DfFYJLzxhnfc9aDXYY2QmRcVGwRShrLCc6dz5/zOaJLKZMH6SQrLiBH7
geaiAZKsznJVPyMXkGl+Iec35fq6CR/pHMDo+6LIMYRum1OCVgf5l0Vzmm/rG7UT
d8ixVHC/D6djnT2lZBKMWZk0QU4hmeSgqeC4+LgKtXEiWbB0BtjQfPWyI29o5c9m
EtFC0oVa5LRoM4n4cGhvp6fjco23nGNCrIykqNtI4ZpVjk/1z6o56RtOqCTn/NhI
uSlnQyu89Mf/Z9NUcx3Ak/MrIwIjsgka+bUi/uLNHCRvLRWYYg1Ef+qyeagN5QRc
80TJDrtwu44fMY4YASQqyjAjlPP7F8TI56fTvsskn+Fw049SZ/gvvhErGU8uyuTP
/s/yTq1MvM0tG5Hqo0XjGP71Gvffgt8DkSxSQVOrkIONOG4uZgq6mtO1Pq7jmb1j
kTf1zJ3TO8J+qf/C7ebperOFMc/G2ss1f0wfB/aqspu7Z5nYvvFCvTrdlLuR2ipF
/ZhzDAUG1WISSs2vLH/Q4ObBC5z7Vb7OVhA7lMScpYv4MUCtxeCIKjJhQ5OL//eJ
V6jkSDV6+mFi06Uu23nsf+KhjKCDHE1duIT76qcYALQFtyKL/08ZCZBHKvgNLFlS
3v5nQZAu3Xn/hQwnHGEUPAiGbap307Oye2qVjb9UvBW8+RR96SJxnA1DDpOPV/Hw
58tRxVajJy/ZW+cxBN1f0R0AYwWAZKQbH2AnOteD2TG4jT+WgEl3SgLeJd7/69af
Z7SF7/MRzzq9SCcl7m9srxSct8NkQL2INNjvb01BS2XVJeWJP51nsNFBK8Vx9hho
kfm+RJkabZGTAbCW977N4yXmdkT1DndYp9pa57SvPfQykl8mvnMppx9VtYlfQqZX
REYSNRvZIeoVE/f0AN4YXIkPNtbWfY7tIw56EmiQy/u6Lid7NvfDDfAu4tTSk+cK
X5JGg+aHkwRW0e5V+6kVUVTYXlOV5FoupbEthx73sHy1IkC0BeDHxBPP3G1NkB19
wFZEYwfOnso0U0ifHn00Rk7HYH27U+0kcMyDnLYhxCbs42MoxDCC2bauDo7TwjC5
FPbd3u+PNlWXQlL84Q3E6OngfgCUwBJpJeKid5LbKPoDd0a9NfAhuKHX3ReaOuaq
RnouVgFBwjGzj8gJX12wGDjTb0FSHeVoAvBQuEZolFNLhyBcDGon3v9eBQbWg1y1
ijnoFiLlhdr292JI9y4sT5WrbfntmF5wKUFIJCDPQdqdPx095Ho2v3Z2NNSF+t7E
F+Wwff48fdjy+jA3Sy2PH/a3wKF6U4gXyd1FiMSjII8E1aqtaNav9ubTjbsIPGQt
B7eejm1mIvBHO8ZJUJNhlwdOpz3fJ8R1NkfNHse5v/73iBhDCWXqT0zdoBbYFGPJ
g7Mc8IcpTj6JoT5ughglt6gACjAVJQbb+9s4datIExCGVB3Il3f/+8vBs/oZOTbp
5U9AxcQWFt2oFjFwAE2XxPk1jL5lh9Vq1P0bc1CEsNnJXb1JgDsFOzg0viGQ6ilw
XWpo/qvvRCvD/OOIMZI2vaBttZq8HemaG3zCpfFcWncNHJWdVt3t4S26/rzGPjTr
itljDPz6Fiz3Ulr22XvkbM/IpFeewBPLVPFhiMs1ug9EREoqlOdcoEXDFcm2aBb/
JSssn/OcNMuR9B9Xg9RHZ4ZoX0x3HQL5EqcpdNzp360iCJIlFjSKbGzDAmpouLUm
r+jTErNzg6IND8aOMLTZgbk2RwfrM88NIg0HTgPg/pydjrrXoXfM1LsMXDWulNB/
Of0LtY8SFF4PEIGt9/NEqqFq7HKss4jVrbouh4ry7TSy8JWD8AF8WhQ/5AtOa3xR
vcsV1NuKq0FmScyiILBAvpes01oq7smDOuLLRbKmVXVadJP4atl855fgbfnpFLnK
ocg7hhKD7d0ow/PZDfvCNpGE3S/6glRsBU6yIk5epVtKyLs9XaqoZF9KkM3vE5zo
nInvjhPhY+SERtrEnU5jvbI3m+9JpTMcRXKCy1nIi8u/3FaeBossjWnXHYsWwOFf
QQZpy8uGShakjd3C0HEs3ju2hIJGruquXe1+anBEMHmK0awvXfsT28HUykMQoR62
zfywiKlKgc3Anq87e1Srux3QAaLqtsJ+IbZrkfgaoo1MrAhV6Tx5bom7O6ubF5c6
gRaMCjlf7Jz7wv9veV3o/i0q0JamtTB/i8N7v0jR2wfgc5oCwkf4vi2cC3qmQHIX
RLJ68zBl2uLE9n+1phk4LQro25+v9bsubSMb3f9irFIk0iTOgrPq5gdDhrsL9NjF
TLyIr1BNnEM/hoP8GEBJqWDym6dHK8104wdf1K3SnRkiKcFd5vyy2n+vmXfxxeMr
0bTlMmCYuywYzGeywtgTW6fhMLPOxhBJGEqfvz/j/KMCS4PCXwOa8JQfslK25pEl
AUrYvgNIPdAJpjVVNAYJOdB6n3qGytqdhFmr4hG/xDRRVXe/xHSy69J7othR8Veo
wZSCzeTZglvIXYmWCm7SOeqMo5GnURL55O0u6xMyc3w8vNy/E+DMuOgOxnHO46DD
ubMELmJrl2Ek53r+QGJVexLPicwNYEjtIF2TDSVagSHjtWfnFmiAeq9Cdw0byq/8
NAaJN9Dqxn8sTS4qn7e28R2dBgPzu92yD6scg2jmRcoeuRqEwCuqz6aAIafxOes/
o5fnCUIPq9hA5BDuUDRVWHC+/5ZHW3KFo4pk10mwq2ylD83dBGAR9SgAPxUyPyXG
31/iyl6wNHoiGodtaSM73FfNLvFNn1T6HkXasK2FYw1FeMFEnJqGAXtPisXTZing
vkV3O9Ik/IehlRAHraiJPpJNpc28OkboISysaEd7hyEiubEhgIxw4uV+sxpR9Tad
WjcCALCMhUjaXzU3EWkVusPSNuai02RrZckir6L6c+B+bc06OvMnsbbT6WX2sc7e
9yaWFkDvz/5EVWejOapBtsmfsUB6mJtgFqB5vj5BR4sLGFttvbi5IeAbsgLazKZ8
wjsVp2j2uOScTLZKY+LyrFZToJRXIYZjPLsoSGrcSyleEwK7lgOVq3e84ZLVahLR
mvfqG5AyxLXj9tgwUmbgWIyH2zma9ZZchiAH4qEmS6KKGcA+G9EqmBazzXCpsTNc
jFB+pjOUcz+9Rfgc5qn+OSResw3euVAmBzPW/D0S/ll27pxKHgvKi9X58lEhlyG/
zmveRtqG3OPGnUKssQHpCDvJtryojHstVu0ynpodP1cgctJXlzeMWt2sSZBblGkJ
KsUaacWXhiOh2U79/TSL4EgKnG1Lo/otYrPn440i3uVy6gUEYUXQsUNd5npomDmp
SVhmdDYxwO1jBVmzdLrOJnpifD7sIzjlIAOt0QS3iW/K3VKKDJ0RcUr+5b5pA5t5
WDCjn4ITwD4AuLfcEMi12LOzKCZnhEThEoeqQqF1U7RleUWULV3CZuRA8kjIEWgQ
M3kMsG8K5A9N5QqB12tljEXgUR3r34gHAAyvTaDvJDUWr8jW/o5TrsKIH3bx6ojU
2+alIC2hkKDfUCXQqDUBB9BX4qfKBNC8nThJny0wEte/q2n9jTcsQ6fsXjqJODP6
lu8wZieNQZzcPQ6RcgMr1K19WuDIAxlbUF9LUphE9vd5rjrVBWoOPvsIZ2bPo1xG
FTpvqHRcPXekMGFvrE+0y/6Vhcf52IfTkZCOAtrdr41Lvqf+w5/cfSB1U5Yr/o/M
A3mj5s5V72Zq/8F7fzogKwFmuptuiq5/iRKV4gETlVXRk50+hDSbiuK1L6hlR4bR
IHl/KwUs6iAlUzqJ0w/YzJyCyajo1aESFu8z80bTrLZGsJJzHWrQR8be6LeZ2tz4
OWxV0RaCk8n28NZ9RjBZ+GOOM6TlTUidQaBqk4a7Q4p6SL991wOh7jTZsNxRiqb7
ZZeJ5Em9EpOyQmje66LUQnjBn7MHGZ/vHLUEpAxbuTy9VBrzr5qv7KWv7HMzgz5W
wIoW5mIdGClC0Kpted16kgElue7oi6/li6hgYsDpZ75KWlcxbufFiMi4tyG63N14
zehITEoiYiSXdITd3PkP9mBEoUgjuAWU/3uy1YX/wO4whLtWXaABK9Nru91UldXx
O7d5Yv3sua8Tyirm3IuM8G/ppaO1cASX3F1AnMsq+PKAoobaKETyO9ckyE80ywiD
TwebQ8YIGFjLRFH/ach0aibnIgLVo6QqSWSmITi199usZIozCrZ77AMwujhX2QW+
G2QlsFrG/WSleIrHPsPrvbZ3s3VkAoGH7OM+Y5i/CtwBmGxK/Q/E1zW7aUd8wy2i
4sb78Y4/cJydS3wp1dTeN2tHFj1Fz4lFNNqdPFpUm9DOhCjybzIqyJ3wI9SnuoK/
SxREQfpdwUTro2oqq2bZBykv9xzXJeYe51mIz44SD4VwKwp7i2d/SpdsX2yw5SED
1bdu9Sssg6tCRDTpCsNeJdle2BsZvJeUxsgZd5YiOXgXLX60Kp++P2Ooo/SQUzie
7/1+5KXC6czKUZOO0M0IjbCvrT2QfETQ14l5XGYckkOV3GVFn4GQIXu7GbjOoMPm
5xpEXNTFZFGglpgn3n6I2sVjJsTKTgZiRXxxGXFiWsNqBE1Yf7wt9JxbmJDWD/PD
ettQ1EMg4M6h7WEZh5kV/vnZdATyHen1p7pAOB/tvnrQ5dWJI+/ZOEC1DD/Hy180
Z2mKsL5bxIIvRX8pla7BeF27w1++7fCRSGhVka3AX7clWh+526zXdq3YxAuVUzAv
lgQI0+Db/IKzElUL8ZD2V92aupD2jI7NIuXU9q2hDociv7PSkKykBLjLuqZhtKgH
Tsh6ML6rzqK3zH5+gZ1+61ZNNFQfrRt+nfqY8TFoqp6uA3Xf+UUCsD6WrjilA19m
XOtTvZ7hDlFPC8jj1aEK2vh4r6NbCR1mo590h7cFC+odhslGlsW8Y7Nb2Sx/khAQ
IBF1tUqhJPtljGwqEVowEzMyDr+v2xNELOz0z5VxzVJuUfEwFDaUjR5v2Hrn5G+P
Nh2UuYgElrIuLUl/I/glse2PtTjfVAtm/GJCBubRZ+srC2ki7NlXBguGfoFRUE79
FqGFjXrGb6hFjf04VYAfO49rTYo0wPd2Lk46XwZ0xaXfV4PUQIgNOOCkdrFuU2Pw
JObSXIUs0p1GiaOP01c+X9L+gt2W4y84ZLPly8mblDPNm/onQ6COktpVa6fQTXnZ
qFG2xnbmq1GeCPOju42N73DOAVMoEAZhRAJKIaW8LA0E3oTlBDrHrZLxlwX+IW6P
8aPQYqZNLqJP7apo2t7PIZcjquEt8HFk5psoJXq0lec9Hnjd/lp8C10L2epwfC3m
N49j3GmKcLBysNaDcS3Va0AHR1Zw5nLTshf/KwgW3HQD2f+Q8dWU5bIloFxBIJ0U
4/1FqcSGH6daB9UzO/L4tN7txtMSlnh//6Ebn1M0JsnHznh0ZtwiTYnNAMO2HraC
j/QIDvJ0tt1hQME+CUlXfAc+zRjoS+cP2rSRdQbpQALsTnz3Usm71612XiJqu6Ff
y3wcopaIKykOUZdWDnnpOq51swBo2tiRKurMU3P/NMt1OFwIbXgQQwH+KhpSap7m
AFGv0SdCcCa/tpRU6iIAGRIezCM5pc+iqLv3iy9lwIdVwpPXV5YDiyGWbedQiOoC
sJfVXMnFAQDWGpZmdFem2g7i3N4yjAEdk0V3hi7orgihyF31SDM7J7iC+3z/nX/k
S7U/HJL28R8z7ax6ROAXrFHF2ATZ02T/oSLoj4/M2EPFfo2s7kbZgexAHBRgf9pK
UgO0T9T9z3BWJntB1cMUcgIZX1RjvoXuFAFYcopZU/eDw4S3TKVDN9+om5TJGTEz
Pdwggf1YKhErfXnwzN4tD53uxDe0J2R7I7wkNZT4dMAqRafwnKPTZSHJ0T1+GQQr
KSSO85aO9Y7fHdb6Dz9ezLgu7FjPq3c9p0Jz0UHa5ojZJFN38ELxQy84Zx/TBoYJ
5oP1/qF9ynyHmriVTG8NL2gF9GzGioR2r2dlcGDbpIVYSzmfmahYySPH25iJj2iu
eXECfMqBG4ddTjk938tl5KwiCm51zytkvDb8rFL5VueaMrlCu1Ms7RqCrgu/pwTQ
iYczVOy7LrfTdMpw23Jumfg2VFTK8wBrusEJHFkCafZv9tvq6txb4oSvnfxjrLWo
EPqU+c/e9mRXop9xNmQJcJel1VBCOQ9Q9m56C/CDNoMqRplWBImuU+BgmxpEzGK7
8GGv1ussNh/o1e0RLODcMjUpFAzC1Xyk13GATdcJ4OAx7yq7z3/gmM8cO6tA85n1
bYUS2j5ecPblXTlfQZY5Bvyki9UJ1Q+tLA6bn6M4EbPt89mAQz5mw9X4naWd6tOv
TWPWpirvSXwbnG9plFjZPWnQfMkzTzFrpbQsYYyiQuKyr/SfkeDmuDZuZeXsxKI9
eY2V6h4Ev8XiKGzJN6pWDP7Ht/O6w4hdRijTBTqJo7TkB0csUNOq05kztm0Q/zA0
NbfklavVKxGiI+wgWAbJzpOTuoL2a+S0CMJhvvfbGCSw0G/CLD4/xuaPdd2r5E+2
4bQWZkoBL/i+RDxYPqWN/sH5fbBQXV0ZhpMmeJc0YnLWklCG55EX69uGWYwtKo49
XGK/CtsF0cLkJfC3fxPwqEHInpDeqA01MuzivhBPOxzDMllLEG5TvnpEI6MD45yS
ou3GdloVg18LbXyDWOwtsbmX4OwpSt7l7iK4QaxJdIvrhKfyxAQhaAruzCrIYr/i
sRAlm1yD2OijjKcTU6jHqQYB2KW2aneNUzDr95VlxLAV23Gobr4BK3dDImqykr4B
QP9XbWP04jYWPgiuh3F6bfnUIFVOrOrCPkrY4f+o6d1xA0nzvjlLiwKPGVvd2qDE
AVOKw085dy18Bl3kE0UU3qH83IXAJo5WFt2O2GxzW7GFP0lwR5fQhAVVD+DXvOAb
6yCQ/4iH6HPLpPzrTQ02pTAkD+pNgHCfZcooBa1y/o0nrqpmMrEPAMph1UAKabmM
MT7uW5lurFoDA5N8qq6PYE27CguyBQEjK8Dzt59Td83jXmKpOyv/ZCZajipj/xw5
nD6mY9IqCZdUmrSUA2Eb9utlxpCM2zb0GqRG9sFlJyKVi9QVkosB0R0FOoo+rIw8
XOv5Y0EaOohGh+8mRE/kqAMTZwhcbDJmQ7sBx3w27cfbxG0PvF6isZDgG/VsTSuW
pqDHZLgytTScOxw6Q/N3e02cl6bM/X09L/UrGLvIE3q3+Z+A4CIKgHq7XiO6L79z
WG3zDYp62HTcqhgR+l5Viel6yR8g/wqAPdVB67CzYI2de3CWXG+TrF3kN+UHWt/m
CuFcYBelgo47EEhsG9UvsKgXBNNYAMOda4EV104Jbbi6uUmpp1e+Gns5/QGdaaim
hWo8Tkxgi0xPhyTcYkz4qFkKuFjcDiNLj7fDeP2fke6TsHt2jEMxCueM/fj/gORu
00+U4owU0LI3pZYhcqYXE4PY+iMWuM+3XPAqsYwwjB54IXVJ9fPF1ThZqY19Q/pr
l76OFnvaq+liKDpon4wFn4rpbwmzmsIqGGAjWGI4FEJgfCbg9mhzS2axyBZaVWJY
eI3G5viE5p4adHcaj/mvh+femnwIgku5lOqKfQRBFRv2vF16UAtCBd6YiuH9Bc9T
awkklpypk+UksRn0kbD/oz9MQrm+8/VceT48+6ZFbDTPfu42Y1lvrfvRo/1CCZWa
gioHAyu/hkKoeJSn2u19Zj4niOINdNCrM3NidxYBNqAnX4l/WpXJtIaEcgOsZ9lI
J1e5toEOwSRhIaSYNr+R4uyoP6U42n+KmB3YzkPGSl7fWchl0+CDLtTR5QDgOZ58
hmtMOhkW+K1/m8WFeI7jWC3FUeYu+w5vCHnivVC/8s7I2zsFeeUdM+0NCOY4kkvo
YYCUFRPuui/6tX4/Mz33oobR7VgotfM67dgY3qx/uDQ3/yzZFfpnd75cZRe2lNSn
D53UBGWOn91tb1pce04NPMWcWp6F0ovYnVociInxIxMCyuPnITeDYyj7sW2LScOC
KDWvUfluLeB1YdzsX4+u088kMMylfZGkH3iEMIVaC6yMdMsWFw5AL3TZZXKKPHHt
2jdJ4tTGAPmdewu1ZpvJrpgfVdvWRUEBp+2Dl6cOpAz7k9xpYTYsCLrll97mnhw6
ppd5r/vMw18ILaoEeZ3xd7bOiWjFj7vcUVhMIX1X73FBwgisqpDQkvnLdZSzfUbG
wwq757s6J5mtOM6O9tf/6nuIch2DmMN8cGrozT5R1d5ycubJHH/WLG/dhXK7SgdQ
gKO/bh2Q7G9Io7oUswnL7xACHX+fG716wnhtD2bzJwaePfL+9bB+JKjq3KR8mRgI
/Ql18Ji+W8duf71gYM7cR1JgFdJ6Gmc/jX74NNWd0JUtL3Ib0O4/eHfGE3Ik15KY
woG1uKUcllFpsOk1xYvNSir+LRhrzbvepJAC5DEomG80WYHosJjzODE7/WdJTGAl
9lZ+idOuUdMfFh/ldVCggNGU5hEcwd+DwdgaLatLLPzsKKICH91bh0dCXu3U4tTI
BGAeDfvV2K5+Xc0rN2AtLkxjAwmIhAKLu23Cgyf+Sz3N9xdHy46c9rQZ7chqPrvT
b1EXgKAOESKJr1+/qSd7by340a3xsCQT2IDh6s0tJfBre++DNhN/PxiYalC5rGdA
dgXN3fxTrdbttEB1+I8Ckh5d/HJzUhKvLiArbEya2pHrtWAiUlKd7tovf9fpGpba
fswwsPQqVz6r0/150t9LPmHmzKD84/P9fZkuEEDyMvCvnh2NI1+Yv9qPKrAUzcWx
adt4NQURvI+S3t8wYlTP3rfNhPwJb6rDSio6C2hCi9ouNqw1yoZ7q/sKnszywIH0
YItkvKwi6TAtKt8pXc+FbxbDSNviK/54f6jImZGz7+xK8pH7xOM5h1W+5byZokUk
MAuX8tXfcLhNAtN0m3zgkV7VDdhuY5jIJTDgJVFGTZR0YYjNHDmp+eJnDdCjv9ZH
z6zQnTZfrZaAX/R8QIzM+QDirNkFMWcsqBvYI2GsXAV21jL7RFymPwkfJFuoLG6p
MOciBnAB3jJR3QvqIQbwAvmrM1FyLGzIjX0BByB08JFRJXEY4HoJZrfmden9IuIU
feYcnqnVwIi03yJvmY/z9TIU98lkGiKXoyAaKxuXy+ZzYo7/o7a6JsIgs9CS2Tih
2BW0/CFbCgkxACod2vj4cEQQTuaaNv3RAGhb2XmeS6deRyB7i0xsqGMxW7xy5rPs
KiE0DvYo/H6mzVlDpDuIKbMAKQ/ZOwfoiXJn7muOkpop4gE9lj1Pfgfai7XAv8bG
chiR8ydVlS9le/qOD4NDXsGKZnxxJCfDEs9ZGOxDTea9cd3PFPA/CW/Il7zhzX4s
IxDJkB1GEQGcQZpesVwddj+jrt4FEBh3bWiTtYaWKphe61DjXsalCSLm+nmFEmrw
hzb6xM9Je7aKOSdJwnkfy5+ohUTk5F2Q6Ioj4TD+L/7WaKMPYoHsBSVpjmvo/1Em
v8TTqpYiZD0Y7ZyjtrRyz3XZc5sxD6sRHjj93FJ2uuhXSGNEDkBjNxbw0UMf/Sp3
vphd+3mn+hf7kpe4NJQr+KpDVzyaHEewhMJBdLfJxj7CojGA31W+dOUz572sbS1J
Li9Hs8lBa5fSvRbZ5uc5Op6u7GhOwX3bAAAbkGkccD1uL9+606x8TvD0swZomMAl
UKI9lrYtzcjb8wyQrIQRnh1ECF2aAbJv1OOVqJqrxqvPAk0TqX4C7CseD8ECjQtk
IvhCK9Fre0+oFU5sYM3iRa9flRuxVOqTMvDffo8yjFiGsVnyuAWuHXjLQIztGV2T
4plFfpW/HK37F72GBWY4DhR+Ds2MLVemwGsl9KByiI45eJTUjzmTUcebZe6d7RG5
88ps8keRttNRZ0Gqm5dCL/CWrG/V6Eu08XfZ0MhsaDIAJ3qyT4et/g8X1ZgE4ji/
3Hf3M719mtD1gafHTEVRGdZzR1FW0PfWPp4ZmIQdl9lmyMBDPsceR4/SWiJJND6Y
s3DSyrMNXrX5F1tORRH0VQ3XWR5nAqRW02pHXW1wk6xwIsnneDejgOGLhZxRqCUV
IHjAcYOsHClXZt4dr9ZSxabulyRe0D6mjxaexc+/iN8FG7SvKA4ncnf4CJcra09z
koA5ViyUE2v+PeLtCHAbmPvaIYD5ZqWZI/JfbXUcL//FU1QmE/UFtgZ8VaXRkyMw
OBNLODfh0EMUHJUzz1rqYdPUw01yUB4HLYQiF8Tbn/YLHL72zDKCtB5qm3+SGgY5
0T8unUmKeTyZWGIA10o3if2YkB32bcy3D7ELurl/XStrnc02ds3b2Z5zYxumajpZ
jOGzpuJUauEKE+oYY/qoFc4sh8WRPP6LG0OQBAE6OS1tT+WgJoZABU4fUCCIXb3Q
4ZJVemIQzSJA+PffYucudu558R0JGA8Wy7QFz7PlUNlFUrrv2EQVhiOGPz2M7Dop
lP+yZMrCKuAUaU6ZGaa6GF1YxRtZ5CDU95hzPzT+zIRaA7s8MT3uyDKNvuFcwhuo
ux9KbuKhBrrKRfUynhmQYkfwak9+StzhcZK07KI9BDRvL4EjwW3Kk5XTALa3Uhok
DWQW74J2ihL74MmPCr94jkfIsR49a+/jzfhVmzEYqVQNGUo25BO+6BkgLrRifxhT
phr+wUMC9zA8Vxbx1cYME9R6EvnrtpeYDKWMJmciJYmuZKCTmbEfyHrOphVCnQMt
EYfMpGJiTfPa//Kg7DRrUYHe5I1746q8hUBCZeWMgzdJCxMZDJPwLDxt3XySdYNM
jkuyYSsiImRLFQlj0MzXwyz9u0eTfLHRI5dzf8i1Dhnj9yhOSH7TMu+4K9q0f2n9
e68UaIrUcjTCyP3T4IYUSKUs+9NKiShznC8kyQ+ghVxxajFUsaeWZ/VIBICpBCHU
m5NJtF8lSrsFmP4BV5zFf/T0CztG5widb0KELME90YaXsg03+zOrMYc+JPslP2FR
ZSLxvbylGVgisfR9DHsQ3brFtrqWzvON5z1gYImBodLapCZaGlscoc0jROIz8A5l
VQRwzpftNY/OmOJxiYBNU0J69unkLDTFLinnCAIANr6zGCmI97mnH3Iv9ZW0uj57
v5V0T/AjyZ1BEqUReN1uLbkK4yqHt9YUgvNQ+fObtAMsyfAincW67zqQ1Zyk8ycp
IUBSQVpfAhEoXNyaqmfAGed9FKPvMaT92yqfpmo4xNyxRkmBIoSDudwkW/+FZuZR
7BlqCxa/iwm1glYvgWUDIjhqrcA4qom2tIbl/JmwXH/qRBCxPTwN3z8YA2Te3Uui
PgVA4d4aQEcm9HSM3JJB0tksAZU1xknnmptFlU2brj5KR12y3z+6YEFsv1jP/Tna
TIDKMxi84MQRrFh+ZJZLoVULH7MNzOnxjjg2Kgv3+dzgOGvmWIMvJWD2yIEY3AYZ
88y9zqPK2r07QTfAwEQ7+d6hNm7vCg91r/RFUsTv3QqNfL/UdH/MyTKoKT8uPN8I
7NvvtjSY1ONBsEtDNjRsI3M1sGvosXNHDORDdX3VdfS1wVwEm94QUPhgYjanBoUY
82LelNQ3PCysngXBPwYP7mB7LEXLnXng4eF0LfmK3NYXN86TUyaClxgJ3pdrl8G7
eL9v8KaIJS4wrvc2MCC0IqmOyUfi5KZrzv42tyDNMARkTMaR7Y4tSmQaC6XhVWcV
gj32iKoFKQJj+/s0uOQlh49LLmFkes70+w/6nZA+RqX5O0Of1tvpD7+acr4qVPUf
yjx5ux0yLOx0XAeXDhlidoGrNb3mKnF9kCpzqnxM34RUg9eZeIbougiMHrSnWgUc
8KFkIFm5EfH5fAFcnl4EouYZJbWMpZzeF5MxM/dGdbd0CVfPtsO/tduyipQmyE5c
p7qvcbGONvgW8vBuMLWAJ0VeLX+9QhNbxVsAs8y9s4xin9qQxASvwidbrbp20lav
4QomPFvMk2zgCxro7ceLZ7E0KwD+zOjmvV73bIujeBaapjfX6RzbFTObUC3/b+QY
PH1hsxEnA0SrsKmA+VgdDVS19unOZeSbrtyLDY6sMXi8727n/bt685NZL1UDF7H2
EahnIEM/VDzDX44zy0HE5rUfkgAfyNFJ2ZSOICIReMU5cASRjfiankzWGKOSZX3E
8R5tIhP9FW77SvRaAGCJOiYEa0PY4ll1e/8NyEHTiVlJ6bjHgprEiyi3PVzq3HRU
DuN/zHZKkeF7foKLiJdqPWkY2IKKhmbkw42+YIpmGk7KKGMeJw8xoSTKmhbTj4PE
6msNTM/kHWv1nmpwYid7f2knwlqMujT7xhq4kSgpfbzpz502if1k//oGhQ3ef2Zc
1sk3Q0xwMEoamkMXERkzY8ebaorqxyGLlErPBtfwvZ/GWLGrEowoh4wlnzFfNui4
BClB5OoGFM3oIdjA+0RiOwyf+iSnGTBf1I6xjm/qn+LOoWv2zMdwENK6vyg+4Y/U
nfV1Iybz5jrfWawgY4QxQm8LCOq0nGuuV4uayGJCYdgoXdgC2X7Yr7BmsO0KUBrt
LeYUPTbBx6oAtmH9NzJhMJrOh3hxC7z5UfM756RuISHSDVPuH/RdI0E+A9KEErjf
sfqb95+n0tnYM0nx2QPtJSqRJTahDvmDljVOHlk24dqPsRpOTkisZqXulPzYOFx6
QV26m6bsw/Vf5qKyODk/xkdhT/jPxTviPf+KcB6PQaoGm6bhp7CQcIX4f7+qHaPA
TetIg0sZK6KF0yjBhPLyvrEqruRVT8+3d0RzwtSx2/CPs0/iNk9uZlCbWvbhnDk2
QX58TaD+d0oKIuVTmZeLNSWF4MGUOTBhSww2UzmAQclHzxjfppvDgSQTeol6RJxv
YOulMJ6ZZOYWpZEf+r8TaALgGQQvRhfto1EtNf74eM5CCZ2h6suLcHhXWua+wbQt
QqfXLOtVMs7nsoPXzk3eT4c7BGhZocw/byZLKkyGj0NDq3OeRvA3qrWNY86Fs5ob
GKa/C0sbAxu4yhbqMcVAo9Yy/Rrk7YjWQmxh1rIbrp5vT0THVECqUBp7Sh81kbKV
ISvyZy04Dj3HQuj18virDRhoxHz0MBTCrUMdxKDEXirs5PWc7ynJTrA8GkoJ+jHF
m9OTFTNdAv4FBZsOrdh5OVrYYMQyTol6Ni0BJY9v2+2ik4Z45E2oXTDajxv+87qI
RwFGsiUOVJYLrp0SYBHojSmTcOklccR2e4Dbea+IlEWSuGW/ni6XLmPWq8FTdbtz
Sq8NOpCfWxIhuz/sA30Rg6XysOlKpAc+6hOcPtfekA/xOE8LfGyLXCur+q8kS5EN
wx2OCv2KJRSI4/Dyl3VmMe2T0TtqF6MlDVByB2jtAFFYSyUFJncGlmM66Te/2ZHM
KgtJHIGgZOSAEgvZgBFAUVmBDH5a0bP9uKYlhxZinILak1q9AA8Q87K0H2tT1p2f
fdtwdusfkEgKN8YlnpHiqUMot3BEO0Yt0+lTmrqhsxzicWKIO4nLSC6mQNfenaDo
mSirtujDQV8tvpHGZw4LntXsFuF+z2ijg0VTBaA0Zufx6/muDPEIWLMdtHBqr7sM
ytWk+Uj2gtOY8//6HIREBUgdDino0PZ1nnU2VurqUovJsKy7GuoWrPONneduOOlA
ld8CpZcLhkNUBmckfUpyrlcm9flqNdpzgJFCawGlKr0+Tln7irPhqqg2W0EVjrF6
lL82BSYKZ8p+OXTSNR1cwWEGlMqkDof6kcNyLtRfSnTe/7pdiNtGxzSy4+3qu3WJ
qcdCiEn+9Xi8tIdsHfI8r8J7LCPLxYFI5sNJIC+pgRj27sfXuC4pw3UnTmHDE9Pd
cCQGs6l4nalLGf6Mw3r7C4wMjeH/xY4BZ/WiPF+wnieYbzmD1lo35Y+JMJ42zsA5
phEQxtGUbuccJcrdIrNqmOi5VDlaNzBamQRRqE79dTppof6y2cjQruqHbPSXHBgT
irDyT2yWaDB8jhqRU2VuF3s0cY0QafXHOOzIBe8GV0O+g+59pNaXNBRzlZv6oVxd
VH0F46KCSrMLPVIhmp6m8BmNPe9Pgz//QND5ppWv+kxar4a8XrCmhUnpkqTrurYP
x4s1xCA0VDmiowJWHUJq/Gpco5Vw11iLBQGOOomF8QQ/6qvxxXTE4wcVUFMc/2Gq
XbSUFThf5DRJo6mywEG3Mx2V8F/VPu5zAY632lCvEvzkVxdI1EQrwo+NLrwFCJQP
NUK28UJjB3Tw2iU4auSy6FMLm0ZJ1Idxc3ncUBQFX0mGapXFRE4DsKUfEFtSkt11
z3rIn1xQyNngb8r5rZudo6JcIWYHBsy3gMlI6Afm4usshcconEWZBkDmocmfp5XT
ji/LrVl4nmXHEKM8ffzSfwnHyBlp64Ny97JyjT+39r49fQxOR7rPCP88BIUnau56
A7FkWcdJiwtfqP+54FyAZxehU1dN8zOgjAjtTNUDFPpYX/Nnk9HSqDFOAEMqyfgh
B8sAFkpRZntLuPy+9eHLYyWun7CDizh5eJRUYFMbeJGBV30oSCHSuJFzpBr5oKWv
TWICcAU5ZzQYVnOTXIPNUcya5lA0H9XOmnH9P2NepGH1NuhFNcVIcaCBr9kr3Nnm
pQzERuzg72d4yXtDBZwdQe9/BuVDkHH5bE3ID7mx3S3eiLmL+Mu224UZq8fu57Do
c0GRpQdO7eYvqIdRK/0+GTQe4Rj4Y639oJ5DlgaOTHv6pFgWn/b2KVvnuxTyhS1L
5m5jezbmigWRzFPQ5n4XtARl+QeoW4gg9AEDeYwzla6IWJqUyeiFl3HWMG1KKB2I
08BJ6ijeAwTXu2tinjpRUlmZ3ubdUWDOCBdRReFXDKsFsNTagH0HOx0byCqa0QPL
jkTYrIzxYDTHmW1ZyBYkSEv8SGV1RIMIr9iW6SwZ8bovQvrcNTIjZrQQHB750Sp6
+1RUvw38DG7OrdpkONfGe0QrmXfxbYWBQPqU/pxO6IQk7FZQRujX0FxL89lV6AYq
wCvAp3DG8qXTkkFHMuxqWTj04yy8DyOsbksh+jLgvMGOA3oxmcYadQaNKqpENgzl
/qxeyLZbC/XWh6Bjx5nhku9QWcw8bH69O99mRtto8wScdJeei8a3vaHDtLq8XTec
KR+S5wW02ysz1BH8ZGV/KD0oIBP2UuQ3hIk5ewZW2ihQo2duGDOzDAThyKvuGaJI
5DzLNr+u33NP+GYlosf1+weGcOrc1MEl7MY+Jh6eq7sAzx/t8cC14JgH2ECKzk5c
1lf8eR5NEUQbEs+MZjOsApT5IHpDBlLk+VQENm5yX9HhOCa33SG6dz17o579X0bg
dzFKGKZtSvf14tf4GELPxhdhmCbG347J/n62iVwbvHnlzfoYknEoWscEARaVwvcq
NPbEkipg96o0akN1aU1NwTmUsgJFcAg3GdmYZPzseKJhJ7itjBS37DSu2GxqAiMc
rwvUf2bBnMiRgtjp84gv13UtZ24wlH4T0hy5hG2UJdTM0Nx592fAh/KvEmBUHF6Q
ywOjWAS1mdsRTmfjlp4UrgfyrtDpsVKxFM0BfAI1HNaeT/n0vfCJqPIfkSTG7KC3
+pcaQFLUQvNfs26oefIyMvzcPnKsgvmi3QxlLXhHKM4WokT9re6w8h6T+O24oGn6
PjiH0nqOqrS4K1FnQ8r9MS9MA/AvKb7v9vBnbwPTXwhFuYXt3ymbbCCfin665+Ej
oYGPB2TzTojHKOEdB9Me5uShQt1ffJSWNR9a5MgclGcLs+8yXeB9ALnyM3y7Y4hv
Nnh/IyHTVi9i5bL0wDvBRFy9By+TCJGlndiB6hqL6Avv3oUDCbXwbPQn/8NJQv+s
J0/z+wGiv46JCWb8GYd89vCrV7x2roXXj3pUNHd+HwdW+OZp5qF4pnWa1W2bgBrP
LerKv6QGgTPSHgWXEqtP9krZE0XmYeV2v4p+vA13JX32RdvOgl/qANOJXYDGRupR
ZURVlrwrdDGIeq6UR08uZcI+qWYmrNUUkNPHZX3uX+ROx0eJ8xxiXHxscsguLmBW
bXE5q+YU4ZlrT/TnKEO2GOrrzu7kUrLtDdr9AgIlfNbwDyhyLmomsETu8zFGK8rP
wQmE+r63pEzB3PWEVZrpjEQCHLpPzgFOepj3UUTF22kaKAGAzlCGXSpwaFRscDXQ
ohQL68J1GhJ4qc9iEk0j7YFNO3xag44+5gQa64NSy634HLStd5lKaaizUxbgJ5gm
DyF1rn/ZCuvD0ICwLwTy6mnrgecEjjVVMi99B+8EkV/R7EpLCyl45dsrqRbE7DDu
f8ga/BOX2MSZ8wGVQIj2hmuErS/W9Xj41+6A2fnD1mVqXFNktl7mVN5gSIJJldty
te99biFLIZzoZbaDQocxZi4k2VgZ0ijCIGrgfiVMT61B65wvoZ5q7AkzVFWcx7W+
pFBPsHiS11QpoESqiUU3d8uzRlnWDkGhm8RWYLCs1cwKeEq6vhvu70kTxFOv4sBk
Z69e6LeVd1FxZLzkMUumc/YaQFw/oB4xA0EXNm7KVkscjCK1RyjQT4Z4lGjV+b1L
gDjt4uy73ePC8FgZpxxwhIo+FlEb823MZUrZFPfZDae0jFxo3jYS9OVaN+2AjS/L
+EsTIVqPkryUJB4ttu+I/RuFbpfbTBPCoadVZKzWweA7EpkyyTwagyrARiu+3TrS
Vsn4bu9I7PwGO0L5ePX0YNl/weKJzx8SvMvzhgg++BO2aX7nMKpVlP1PwPxsa1bq
XZivBSOIwTBcqor58TGv8WRpJ9RYRKi4KUI1R4+z1pCn+a+bJ62OwzQXB1nH1hHv
kgcrlVd3N/PtAwVmfGMJp4tn+HwmJsCl70Gxg+AYCPLpRO6JkZzo3Yh8JGMAkx8i
QnH5gNxHHcRR/t73it2YTqkXavthwr8q7P7tCF3sxKq9/77RdxKRfk0yPGhmCKVo
FTai5JZ9JMXQbFSwS4I7+eOQiVlE4i72AdWqNtL8h8uK4IXLWJbKj3dwk9dq28xZ
VH9weI1qJEqrDlDjWsHF14fNX/79zHazoJnSV52E2lz9+AtxeUxuONcLaSagzhsX
OZaNiBw9w54HeJaZs0Xa6Z0RoA7AWAONfL74dvhHXhnLNWY2PiSshBoUP2zvWt4r
u5WPrvDcN5ks4ICd3SrlicFJjfmvVZqRQ2t90qJ2+oK1c4qWPkGLC/0q1PTZ7PSJ
2wLGrghw5ZlXLjFjaJG6kEA+PVVGnfn6n5/pg21KEgPWyMBFQ1i+T1PLfOPyJ5Q8
ti4bVQpSdVu9pnEAtIJpv2qeHM8H4ZygqlVmKjAlumleukGigCFMXxal1AJukWlc
ZW5JaPcDEspjXH9AqkJ9VUxt8KP3FRXfjpgiv2bDh99Ozm2UXjQ+AtjicCSfIu5I
96DfkxzbqCnIPC2U54XPoMyZ1I1GLsKt6Kv6Kh4Pe7n8QcRpusdPfCYNfPPDXFYS
vphBziGkwdU5RRAGJCVHIxWmOStaovQFV0XaHwuj+u45ynuJjvvfkpYxgKAHfhfg
b++dfsRLkoARJNurqnqATUiujibM/WQ7BxReplPhH5SVfVZZl4ePSK0oX57O97vb
cKmgR2B2X4PR5j/jx0FqdeGS/3iG4EGd4HC5ABz/+q/dCg3e3sqsILvw7kHgCw+y
I8zslkKO8ok1r1N+KklOz5uRrucngShefnlaNQZ7gZ8y5l+VXoaYRuJ9YLYo4Rqg
Nm+X9/ABuYiCZzWM2nzTTfD3d+RMqHLiPEZTei48KTBEfdlB++hxenqautmOYqhp
qXlJMHmHcjuTTAPi/u7h/95RipPmhRtQEc34CqS/6tkoGOCTMqYiUPKDgaWDB7bF
17ztw85Jdag+2l5J+4Rd5Nyg0kFbo7h+Sp1leFCi+X261NCwVR9RgzE9iar3x6Cm
EKjyxClfX1w8NJIOU2qmeJ5KT7ur5fi+e1zQ7pvkgL9PdM9fWPJ7GCFo42/chfDN
8PnGj2zBFYBuUbJUqsRBeccoFCQYW97hwj9P71kWQdIuf0pdzCwQ9w0QC9ZVJLSv
I7wg989E3kwN22jJ/vbYLITf83oajH2Pc9v69wBZmR5x21Pi34zwbiiM86RMFPjw
ITb9FWVKNwduPm98BInIhdtw2d39x4GdqqW8wXtPWBKck4y6JzG39hPoDt5LvfgK
syVocU/pQkvM4pkjl60D6Dt1t5SU1l3IVquNleGkaZjgM3oxgZMDoFqXYOP9CSuS
SjixYMO5H9dhfbJxV5rKtFQZdRmvtXvbgFj+mBsKNGCBH4Zgql0us3J19Yg/FsGN
qT4bQ5QDba3mkx9t8pG+YdSNiUAMt58cMi7CEXPt3TYwPSOtE9iYj4STvbZZhNlm
xiTzEBtOuBuh+FPSI4OQYdRLAZZADxeENE5t0rBRUrenIIkb6Tk9ToX6AZB6cw4V
KL3WJF4VZOkiWBZAr4JXv5NNftVmjBrB+ByYeg+TiByPragGGGrzpjcgppZruLWo
/u/Y7NV1IhID7+pYafgWtSfeXu3gtMeEIhtyHnbsHcFpaOzyWSGZ+nR96DFJMGI9
Jr19Yipuu3oJMIwyXlN/i2fR7Z0h/XVmEdQ4IgzKHJXnoEhNHXPd1iGrOe2NoM88
3GZJxAcYrvl3KNkVUBhMci5CjcwI/upcgIK72VroR5gpYhS1uTjPukovfzFFNI39
MCXgHB8E6TRAldKi5WHsFkP+NUPAdmryi7DtNdU1oswvPG4rQZYt9Q8QC3ewpw+y
gCzN/6x8xf8X29smlXYyzLv7/ZQQ1Jh+oEGx71w+iEHihuVu0010jf3J3TdWBOkn
tirHy9pk5H1KGS6cuzFt5zba0rR1gEcCn9JbdkS55VKWJ2F6DmvlqxvNvqul4b4q
1xaD/0m3PPC9eTYKg1zKX6TO3LAxeAys2pQV2PfvrpMzBmC37oB8uhajfasog9pW
c5K1pdz8U/5rOUMxJCoh+5WOH5wkkpMHN+kaqSMMVpzSRYVak1clnleDCcMwcXug
CQY+DF2KcniwspDqY86aehvpCpzPiqaS4hrxxgQCMqh9uNS88UAPlZHkCVvu+Ecv
4z2c4G3ytf6lFQrBTTlR5c8gV8e6FgMegPjPAjm9hym4Sq1bFfAWHTiawkyOweZm
1Ic+Bhn58vRYF6seiXdoAS0s2tAZropUvdR2PZbk5h7VlJyB0Erz7UKmXTRf4ier
ZoaM1FwWBgA7ccwPBmmAsB4z4hs5oFEuY9HF92OJb1cn7dqJoFtDdGIGSC6c6ImU
8jT20OJgzDXjF/Fc+7kfEhdsF2c/idrFbzqM1HNhqZOvZLLRYk8HdrvWA1UYgWAY
CTHWnCSJME7dMOccQUQOMldjLdbwyN2t2fTAzhWLAWboPHBJoIACu/GqnjoWuHLF
VFMqOiUb3UjLqhvOuefwi9gOesa1ygcPfCrxcyBBM5xC0Bq92H1d+T4BLKZBaCOw
aqRc5XTEFXXnHU3nBVj8T8vlkfqrRH78CHfkDO/h48Wuzxx0gaj5U+TpQqIUbsCb
1TdLDt7v2ImaO5fapXQTGyOJHl/B9MpXJzgsy6E6cuZdghwSwrf/mtpFPY09lavj
nBNSAKHc9oaheVkSAELYMGNxynQOfkuUsfLUzZkF4gKlBf4XhQJw8NzjyZpiCLPp
xXf7BgtTLSw2diGnJpONBT7k+PvMfaMqRBO1V9jGEqHkvHIAkAX57SpIYFPhvvdz
sH8lK1DMd/8lqvXaBzGbKblAnFW8kS0gkEBilFd/c1zYXsD7PAxPx2Xhcw+GVBUd
6Axa8JPnf2xlf4TmMkxguTeAHY2tLaLWCwVabkM4CPwqGpmL5mpjeNXiDOGRteVa
fY6cC0OhF+nnEHIirz6jVYht/yv0a6soq/PJmEpnk9rS35bhsNrKbLVgoKzAOQLx
jcA03AUuiSFU5QoPiWdvapwFXNyVASDY2H6greJi92YthBg6cP/+jZqybop5cr+F
39EjM4mJ2ccGDB+xhEgkyzFV403C0hYv0XwqzpYbLumF+DmsjLiEgGbecOUA28a4
FLsFq70nKCKATR8XzLSQ7PX0jTzMxtq0dM+E5RqYpH7ohU+vFfKUh7sFkZnNforc
e8P+qebQ/S1jdF1tW8ZoIFGXQamzcYsRxqrU0rvlFGxTauMYWsVDFPD+GLJ/7XgC
EZWFYGiFFcRvgkZPRyguAs2oeTng33xjCheP6TIWlWNFXjK3fH31KoNtSt66yD1Z
F9R0lEKrvaajPBwkt2ZU5ehcCvOetk1qVspTMVINuzGyp9w4UOK2/GZAnJEXYB9z
DEoV4MqO+3/HTi0pobYB2xIz8Amn/mVcBig6cmdGDJBuzvqG4x/5QKPQALL09/55
S152ZTz53vfMrl5R8OObhXE2KRDlHWbnUBGiPojF+Mh6+TZKPC1CK7wq8ZTM/sm9
GGxHplbb4/yEGE7wnYOCvD8Ao3bjfacU7elLLhsDRw9XW/fVYRFOxnRyjjid0j0q
rA3LmfX4i1yFRjO+TaeCnWfmUxVeoPTmBz+uunF0lPIdmRFIc5nOstITPna0/Zrz
ImSaZu1E8RArlmIRD0m/CSFqK8kj3YE9w7qaLk+gXre/AW2EGRzPcamKZ97B3shD
2dialfkZ+AzxUQe/uqI7YzNFEnTVUeALWInOgl7qxsajmEK1Y6vSzyIlzX42zmE0
2ZuVvUsQWZY4nrEGYr7BvRN9JMtXV5ih54VvcH4xVwPuUt4n9HGV4625rap9WQJf
K60AWNxOJD+xiXmMJZcGI//eAWxgb5OV7MBM+NXBBU71TpAmXwIx8eUnE/7RSElo
nh8gLSfGxLKCsZlWx1QOiumwbagL/iqrUaDYdKQ+HXjlPmmaLbb+PcJAR/xsWoNX
9L9nXd/9Jm7eWjocoGWzjGpvG8Av+0hkfcgxnqVvU2YxZpAMCVL28+WcVyewi1Dx
CYFjvz9vc66HCSw/I/v9aKYDENLhNEpIfmuJUpks0S9vW0QKHuXyjLJId/RLxISp
Fy3lJjPXp+oLLnLHE9a5DgW4GC04NU19bWs3PW18F21mFqeDie2ws5lhrSefaZ6L
oWZNWnfI5ZnoQn6vkK60zRRckSFM9tPLvf8icAJWJ56MgPsBdzrAcL2Nwwkg4LNg
S7UEGA1ERjgG8WNRW8LL3P9gR7WAQd/W84JNy5bYhmFHwwTKRHhIxbIZRAL8IZLD
kE5f9kSFbSV9fjQHH1/GwCuf/4M//QBMK/RjISziveXN/fQROVxoo6tPJvauubfj
gOMFOmXjT5XtR/aSqnksjr7TPfaEy28SrkHUoXKjyTmspuu/cAt+cGzHDqczmLWm
pfhvpTkRFIJH6B1DU4sbidAkddUDvL+TRU/m1L1CYZziIo9j5yxenC+x5AegtfwR
xzbzV61qtWPd2YaKPpvhEAsd7Re7G+EnQvLFHMYF81zFZRtyewObmOT3fc1Nh3rV
mTPowe0j75ZCqqy/KCGFD3Qg9qmTxVkzkakFyDfidBqR15JSONpHSW4xizz5lMlU
mR4gTKavA6huqrVHWooD75VGAZt117Bw3u5sqhsl6ib7qgv2fvowf8VQKXjxNN2M
V6TzP51sDMuA3SwX/BhJNg==
`protect end_protected