`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2096 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
e8zJV2MtbGrDSF9eZJaPGQohIljMsihRDU4pqONRWfwcCcc/8TH9BLucbo6H+Xkz
f6sfnWiRkbnY6lOjQe3eq6yojE2wnysHFzsDAOX3M2NN08YBtr6jz0hRD4VY7qka
8uY5I573LAfriU8gp6vDXiBuCMJZZYbbo7GtyXZSpksamIfmfK5/OZgkjQnJSdIn
23EuUCvw9FL3MATYknK8w9vqRi2LfMzIwEpexWriZapWLR2B3T9ct+3KYbelx1uS
Rq/PgPd4zjATEKIRzfZaYgdQwGAI0gt0AxfObAEQnbl3uZgske5LHFdLBZXAmD14
YMVj9VvvJTAklWjkDlbttBjHEYH2lcAPxi71yTnxIA8sPRcTxnnZwTUnp2uJMmFH
nP098BC9n3IjbPa8nMJehffCHS9mMdhxmhwXs+xtNRTYc1OCPIOaNGBaem1o/1i1
F3GvLbsQyPRI/dxIcCFmPqPD+MjrUiwFvop5kkY0ilF4AufIaUy/L4FwCOGyHS1u
hG2TjnEZV705U/PXmb+dwyRMF2XARM6GZ3G8bLu7VE5H3rHyit3MO5N+8DqqAdbs
j3vxxO5APCdBIdMaNQa+rAJqFkEXhGKxT6pu6GWBfVohAyPIkoerE+plYfTg2jDO
2OBswebQCDfwGXda2ffBi+/axqVRhY+KJJO/3Pl/E8f5UnfTYmYIQEqFMF9eBBRa
9T0Nh0XPpzU9jU3OtPbvtqQUtQkRrg+oSjdkkXGTh7g143U4bR1skD0wnoWk0V4n
I6rHeuqCy+uUkCZmEyvWpHVpOmELCVtajVxCARecYiL3S8s7tw86ibaurg14S2dI
8fcREQxNfOsiE+iWV2B0hPKm+AiB2N0q/hzsBQfDhzaXScPngMHop1vYa8nB7/s0
VTnkip7SUhQcUnDBPdVP5gYHBiYYuBiqRtOVAu1ZQlWIBtbxU6pBnhe+BIpWhFFb
W6oZnLuiIAVH1WnToaHXIjW3jM58Gn3KP5DFUtJcF51KrMjay3zYBh0iOZgGmLgR
HDfRw9WDRI75/JqW537abKeIUNZ6ARi9koV78YKas6uaCrJdciVLWvj7SuNslaP+
u7p5xUo5kvyYn+f/00S8b3r5559eZvkGuS51rNX0QzSUaLwLx8OCcKeau/VGnWnt
mmxyAxVLUneFI/qQ2NXKS74gI6uLBbiQpS2LbXzp0FCBBB+AzR0ZeaqgUrElOVW3
H9ZIOhnRtHDrSAlERIAyrqxpUfa3nXFCfcKsRbFp4iOWsRc9XxTnRNnunWlrCJUu
50ZrUKckwdu5HZVosNixY6PSSc/Y7YDhBUvMbUqmp1yj0NwaYSiIMNKjDMvda7i3
AGuZ8Srqvp3zuD120VdC4M2lcZKdvmA6rFIu7/Es+KvsL0t4X0lM4Op+ytI7PFmF
aOxSB1StmPoc5iGzvYSvQzJVzB43AuX7OKCEles1Y8uip0TMp7q8O5h3kAUgBMcL
FuOYXwrj8eth6lwrDN7aDDSuw7xT2RNM12lGrDbwjJ4i1MSu4MPn5YXocJjGJZMB
mGDGzNqlL5KQ0M4xdjiK4a0H29cLnellgCoan/D2dm58NNLg+N/QYs5vAXTLhJfo
RZMpDbOeQnV/DEUof3ioOU5O9wdZ1wYFQgULy4ilH0YC1eCZ/XGUfzZ+DHCz2iAZ
KUyuQJM4Oc6EelYRp0eJZ0uCTjXzwuIAwSKRcFiPbHE4Ipndz1aEHjQXarSx3lWL
PQtFo3XIBd1fYiBZ061ArLFDH1yJOvTRbjPtANTJLXIkTKEkrHevYUFKvyMAtC2I
YNVybLIL44a3gMiCdAyUMxaDYhe7OcyLrh19fxNKwE6izWA74IuSKafbDHqpLZuc
1ZDEsbCUluatU+QNTwKeurOkTN6kKiFlADBa4n2+Tywzd0uwT3c6XV0DWMZvu+0H
Xjuz281w41bvn0kQQeztjmfPnPo/htl57TCPk6yHygIXB5FzoIk6AyEV0QsDOh6E
oHBJziG8vJLEXFfppFYoRPRSY2mBz+CHRVDtTX7/F8sH5TMLyKCdv2G0gyKPeeK1
oInbh0/SZPcICF92bvZcnKqFemdz03UG60iSMca01Y33RIJ7bZkJ5SykOMPB+na8
4OiPdVpVPG7xgEUeyHHXYq/F0XJ48Sq1lnB+K/ylbxivsTSPmlEh3iE/8AcNLLG/
+PJ1P8g+X87Trt4H0hxt8MPpfxqANfxxw8bRMIbY2EM8AoAluk6oBqbtJ0q1LbsZ
vXQtP7ReHL1Z2a6d7yWlBmy+4C/nf01FwGQwferE5DUq67w1MY97xTA6AxIqBZNY
8dQXUp240mJ8iSzeIV9SyTNVsFWC/iB85CUc1x3BUL5OQuxfgjaueQ4T3Tpw94wA
Tpe1z5rD54zBMxyjO+5I2mS7oZwOj6tN0I88Wup56F02v4Xaa9gNdv67WXMch21D
WTHsNIbcYPQmT9H1P3LaKFY0dq19UhguSecG/iH/zwpzqXOg31ABIK/Jw6gXc2sQ
Mp0B3k6DuZFBlD9kR8SsACDjnTe4GUWW/ACX9LyTYKceTwHk7w4UTeDTKJzxSVrf
5q+5AVIYSVURcCeaCy7fYtNX8R2W6aA6apfeE8XhVTbq4PfRcSYpO7D1Z9OPKsHU
fPs8CihNxNTuHsSxprBN1SYyI7UlymqfXIuSNcbAjQ8=
`protect end_protected