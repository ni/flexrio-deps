`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7824 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0gQgIG1mJzulW1XOK5NnZR8
C8XqDUtXW7uOWTnSVqbIbgsO7PF67C7p9H/VUn4QFVt5nhI9PIKDU8u37MA9VZFA
8KZaPmkWUk7o4AMXwb5vK/ytZuS7UKPJIKWf9lseheF4TtlmXX6meVY+xqodvP/N
Uo2dkB//BxBPrO972TmvGgh9dwr64LmZiVRPJdCcbRjKsdLFB8G7MZLcQ7woHCQ4
snAGFDfHakTfDcR/elxuaeiuKSMpz+s5wLfxhagxYwhQdw5KAJRwYPw2VfVuMl4U
A81QfIUGp8LZ2gXREYX1dE2WQszAD6mv0KlHEN+IfLPAEmsgtAUjFvROI6DFcsEi
LXU1Pd8aXGysaVkT2poPnoUnAfZFSy6WOuEoy9kKuqXgA0XCXztYvBr6vzSJw1+V
P2NQJN6ht2ekFCKXrzl8bMA/mOVi5Mv9SiR3qICGQvT+X0mbCkjCyhKWxn+qPHJM
QI4WYbxX+B3LDySMqb8daMhu+44HsDBfYoRup7F2PB68AHltnmnQia/ckVTyAgYP
ToK73MrBCMj7S1C8BH1Lt/SZyOy/ok9KpPw+4UfqAVG6OSZG6FAdXWOWXnwnbgGD
hBwvlwWBVnPZ2M2WP8+PrZvoIswQb8IkcWYEMeTTEMDhs0GjrtwBnIvSnv6ut/vJ
VXvROJwcinjctKbu+HxO/widRmwMzRoDuUjI2ucuZcEXTAYkY6cXqQQmdM75jT8f
BBmHJJdTSxO92puIK8WTlMrY7B6UTbQ016GOS2dDOjP/ycpmlNTrCK8UTNVU9ecn
aRlOAFehyfDQ0KydcsrvOQBFT1eopx395LlX8Lq9HwKs3mb3w6LHscrCX89976Bv
a/w5iVhW1XCgNqn1cHPgxQak6lrzBzgUz4ABmSc9DdU2BHHkVBZioOOpD9xC3YK5
OaNFmNH5HLEp9Hdx+TiCHbzY19PXjnHHCB3Ic1GJNuqct9yxOmKH1RtxGKWj5htO
OxUry9HzBVO/qUi2+Ie7xUgwLUDVd49h7WtsKV2e7iOk0g3X6y/nbKHNjoXnxsRJ
uU0tx8NpNxwRvS4TvwF6iftC6LBtc1XKi1U75eBGm6s7tvtZBt2nj9ewTzc7OwK7
RDo6Yww8XFAaEWrb+tcK2B6jJ9YcL5/tAwFKLc/hwuro9qpeaBknO7PBVhmaYO1e
QgTXAlT3qV8ZhFhH4F7Q/Z/sfVfCgXOuzr9FVzVFJ2p8EZavXUKn4tZpQlO+kBnE
StlSXau8Q9yfPq9KSU4Pxb9xQ4wPhKkoIUAtJEvOuNFkv9iFeXXcjuH0xpNm2xfV
bEZG8dxRAxdEaXIUtTtOi6V4otWLBE8nrh8o3BD2NMw+PIYgeitZO4RRc3jRxkFg
U8Wp57an+QGst/dmqj5qLCSV2VpnXEqhoiBZ33LJNihvrT04wHfdiDrx+muzhXo4
3KW75odIDR9uPMvrr6TM3FKYcxJBkptpMYS/BAyYRgBn0Qjj4khSX7yFlKI3swP8
2wMqKqAucTwSfy2sOG+q7+v7Yo/tAqyMNE057k3J0OAFj3LaeSTVZHJj/e2ZwKa9
KAybZarW3Uqu98+9GAX72NXvAidWGL54EE8i1feiA3+zdYGFF5onRSCxHPP9WVJJ
bW33Jgf934YM+HB2cCYicmWcYCcoWo+Hcl7wHZ+RkIqtMrSXZ2oTE/+mDJ2QNnVk
Hu3Y595QfPs27tbFN1v2zoVmePoOamQukUlSoOpGfFKX8hJhCl1GpPhSSE9lfGSC
h6AgA+MY6XWDrEYrz3s2aa2705U4zUk76FUoIg+3VUwg+cuPvLbA5D+lL/Kzi2+s
Wg73uQxjrYfa/Uzh/kozInVKmFXoTXdmOQj/PrTybYh75CVSMT2eJhcRu6RZEDDM
pkp3qp7S5DNCOYhZyoXQaneKENr/lTZ42eFFDLw10nNauj79Q2Hb3EilcqfbI2rd
oDZcsbgxm3RAI867U7R1id5xOQyZtLbZffMfEDU1uqWRs3pngPoaz9u/l/i2/Jjs
IYkGkik5c++AVgl48dX2FFwKQEETF3vJXgx7j1vD+eJLUouvDQtcRBeSUIb8uUuB
CY95M1yLvjggmJSVq9BG7aCaOwQdGqDFWtKCRLhOppdeNoKRiF/Hr9zCzDcvgOHb
E6aB17IsD4zFB7m507NshyctkuJns7cSg3DTfswv9hxRdoYnCqy2S2IXqS31a0vA
S3ElAC88/wupntsQpyGvNCDSErk4lz3VqZSFLCZqwuP0WAPcejn3Oinc2707NTWD
T7a0nE2dSAoA/QMbO802XpEJXznJuHqeXRX8j8Pvw+liqpWf+gbob0VxKx62C0Lb
jq+7OyOaWhQpZAhkiCw01CBMRZbqnRkwRIj/HomOcMM3DXcQQt5Dy/lzjfU+9s0U
rwWg1v4RGONBCKmsCN3Bp4xX12Vr2QbH8vxs7Pq7SeYnNVPi4UhlMD8i4o7SYFmm
6pA4NzrFkUagdw+ZY8+V5hxQ12oCq1coaDgobdAjQLfdZ0fEB6SX5XmLDm0t99fQ
QcxylRMHgms1+v3CFTFlKfl5jxWW82KNvrjgKwHB4UlN6xDfi+e/sCAGbdbklqh9
D9a34c8cXs4sXlpiKDzo8UwmqPnqURUphGsI9kyfQFaaesa14r20QhrBqgaH4P2y
9zuJcrhg6gnmgUBBEYcqhb0+pn/SO/C4qETC48DagVACXzWG4em0KBSjlo1MNecM
3KqzQM0Hb+GOwzEzD0bxeAJekFcBKbgKX4dDZikpDAAgDh4OyC0tSDviDK/thrl0
bSgwGXdUdqzlnNkobx3bk0wlX3zZjhRNzQJ1dxjzrc0yJ8D1CCiKVwCXqjntUl6h
SOIlC7Zzec0krcDjiI0cdKeunTpjs6BG98nTRUAH/vmtjZaUR8h/QVTgoh6awPF2
C1/Gm/w1pzZvj7Ewnq7jkdwkQE+hU6BS8LxC3EZjON0ZJjRAhT7F9K1raYhOMwT6
rjKMGjmPkCQfYZKrsULeQERBJiQ6f7gsiYj7+j6sYHHnNjyr52aMcSD2+NHGZeQb
knU37MNKLz7myHawk7nzl5Unsq14zpiHiGAecvY0RWf8pCYzgIXV1M+JmTgx39Rq
80h/zeI+AsSblvFBKUqifkqh760+VQrX5SpzyLB2kcb/7jgGXcgYU+ZLFZB7bB3G
hwl2iR5X4ooJbw2uam+1YN/fTTxbdOPVP0upzoszEkElFDPIcjtrcfjhJzH+c50o
BTd5AuB0gsGNKOZMdVLZ422EZDAvxaO8dSZcWFFDKgjURrVG8sbWaCW5Gknx4h/W
iny8zpKS+ALYDyTTkdF+BtvO6VBbpZnTw09UTy09qf+6KC3pYmj4DkvQEhlJoHp8
xvfgY4vql45QViEN2b+sEHX5Moes5iETmYxJiHMzuYboMn6W1ZVOUcAumoFdsNlP
eIz3XsyzMwWHbcP60uib5eelL+e9ZOcvzys3qIaTv3tGAQpmbGFCbLhDwP6W++XA
bzd/ZUyl5ERAPHN7aI8L2qp9SejXBZpCP1bnXgnySmj5N37LYfif8ZFQEFmvfUyo
fJnMdcng4E5mzIXvJ6BVYSQQD9IJGujVqKh8nAf3jfQWtFSHfyO6IfnOL/K9cSzp
ovftvFKsywMyCEyMz7QpFffEWsQUe+UofdWrddC6QnGYXG78vjBwz8yQIJU5Owcu
T2rf+YcSOQQ8EpL/m0ysVpKjp972ZRtaq2txtGLVfU47nV0MezRYApkgg5TvZKyu
5H+Tbt4K96N9SD7AkQWu434XS+BbcBCm93EVc6oqilGpctSZl/zw5YqTLmg59ERa
8UhGNhsmNd55sqby5DL4hCPEHSPIY0b3MbSMhRjmf9PyIYOtu04xKXHh2KrGwYQk
4/ODGpZpKRn5HIZsKHLBPRvPilFkHCVETnsqwyi46PEd27TYJiUbYAg+iMZQ8hrq
43ecMEEXSpBqXUe47cvQ6VUa69c3SUyu8CnTacq0pOQ6f6ZVITD8G3QGF4rkf0Uw
Sa2ZoNwmH1LGyUgvfozJWz4yAzQ0Fod5Ff4vPyxkVX9tjTrCLTuE2x8g8QB8UJ5F
vWXSkCOHiNbMMbdRDF++yqdnoDZZloHCg9mmkFqV0UzFIjMX3fBgXAUewioUvt4J
dFE5YF+Kd7oj81Rn4RBfxOJNaCqX63tkQsqnpaLcT1KhS1mCW0Av5EVaZmie7hGJ
v1YuETLoNbQdKlMe+t/jqYzfb8E1ztrUyxpklkNGjvg32Xh6lpMhTdvQbxVCgInX
EBM7TqqHEAdjerq/rxIkwCk2EfMaBNblxNxYDbyEiNCA5T9FZYWni/jNw7Ngb5Mm
2HfGypilmdP43Wo629Da9qKZXRwjHh55DQe28+7+wzUen/IVQ4CII+iVhYaxZIU2
oSz3pVkhJJbJH2xBTumpyhhEhtoExheiudcyxjYCmGJ0TK2uPZ8gOMVojRRslav9
A6pdm1mGgwftjuyP9wM2Z0IHUaUsl7mKsv8TuBJuzcHfYOhEOIf+OS6e2UTCCOOc
R68d67eJ6rV7LXiZjX6mgJJrA9iy2A/XwqL1JUprF0tsF6qDhOh6DNrSM0+06C+y
pokK2BdD85R0z1hq5SwkwJGgX+IA2mhUTqbwmalpOrHIEPROyFvwJGy1+jRPJY8w
tayDZc+d9COMcjDtnvLLGSwUJU6hIt+sN7SvcAb8CNIlb9jLHD42fNu18AiSTEC3
anqWBNY9Stmq04liXjFkvduj71ps9VJxxsBNmrx6RvdRuFbCgYE7YL1t7TLAXbdc
W9AQKk9GjnISsgCLdLYB2YbXG5/i24XdMRROJYKL6pIIc/kzJewBsyaopeTkVhKk
kIeMiBZUYc3F3Xq3jTojCcFh1awdabDrw9bE7CQ2Py+Be4YGNtIPZ0UjKsW2ZfpZ
nCSILDtFzCC+KM1AZzFLx2PmzHJe2ZretBzdIKFl7tvv7yOL9dXI4V95H38LE/Oo
9t4sRGBXTPQNiVvvjL65hyGi+QSnloPx3yTLYSSFI2n4x06nQZBHoL0yDYz4XTMw
joo54vytgV7KL7nHjsCiT5ouVhqPVu7yeXsQkOfe2ZYhG2wLgBqUVSd88BVbe9Bi
FWa2QJZQR7GFxmYGqASPQnJoiSEf6pA9IyJamLJNDmKRjyBqiL0azqKbKrblwFbe
z+cGftGkIK7JcsJsUlTr7PPBl4SaiyzFzN6MFq4YHwFOitIW5dC8OSKhqnssMugJ
NoshN49L3yf41XC1LBN1djrL6dTGboD74k4Nx4cWcX4rbBw0qHwFfJmQAsWpmrKM
t5ASUoLuix2ggwElHoTYXuuEITJSqzABWFYaAU7yczK6cSklJBYVqAAVtZ4t6l3r
Nj4uXHy8AP2jGXeLcHh1Y9PfGpXyu2yoNpYRvIuEWiHT1VdIfI5kvV3P+K2sjUTE
vrkeJKcPCHDjaTmZ3QimCFqFizJqsajfBANFCjz79R73bBbkihNhSce+qNeXlTPh
OmrW1GGchp0qyfWlyULDTARhUdk+AoDgVUeCfFXPR7qlEqYatcfG4fDulQ/LypIs
uB6i5OnLl580Cdcczf/X3Umhh/5Q6ZJbClzsy+0+13nyr9pRmjG/KU1FaQdix6SJ
PPG7AWon7+ZwBU8PvYRWGhwDExdNZzpfJVa0TNKg7JNnA9zI5yS2rTPT4mYw0fo7
nfywrm1dKQIjJDF+IZM7Tb/rmzovsPnwxvNV5XqYNz67ReC1fQDO59W3HMamKqLI
hM3d8eOVRh63Xsvo17S1h4SafFbOWAu+SipGWCvi7aBaflcKyaE12floBSW0x6ON
F2X/JctivYt8KVX6sT4F2/OvjVCAIK5ixOhVEn050BaabgseEPxe84EY5mRR6yyx
t0xaI95vxkmUF5g4nI0oeLp89HZV7kL4UAaQDyeG+oGao/Cb0GFzU8/GDGwqXyF9
AmLeImX7N8bbiwsuZLMn+Age+A4f9s/3pOSFb4CoMSWP18tBrluTGzloBqBM1HGK
z5uzVUx9Jcv5yAdO9zz/z1e9UAhYKOMWPJ8mQdrnpU+lJNkgBZkfh2NfAK7Ma4ai
/Fz5X63UBvmVq5nV+WQiCr3Xc6h8+Rwip2SwE1Mo/0zBbHcWAmgpgdyj6OuqSV4g
8CyT615spEqfi0mgUvjQWuq8qvxSraW7pKl8KpbeIN0YQ0XEyjztXBzv9Hsd5A0u
znup1oV9ncmg7dP8aNo0dwvj+d2qf+mqxUSC0g21UCq4jHBY8XHQdFuNpPQjQagm
eFre2HHmLSuomj+CqRtqCUXy0XcBbK3t7ecfnCoQifhkoLo2uYeI5LGdD03lOBeQ
4WbI1GVuSF9Ydw+OgAYLWNWXq4B1TC4dp8zYJ7gHWOMpBqRSYfLU0JNtjVp5gOwQ
msL8M9YdlMR+CcPKH9Spr3dg/TTFs2Xwve1lewlfc1jtLZHnViYLbwuZXcnMqLxi
55Qiy+m2xdmio92trmSx5iP8T3Eoyy3ZwoS0BP4ukj5JnXhytlIhbyiIx46DXVuU
qHKOyEvII4F2KG1Q1dmbpy6Wt7KUubT8ooKfZAuZm8A5vrDWJmb+373EnfHjvQaF
R7xl62z8pIyaMXhK/ogNuBPzZIUlBn1KN3Uy/qLRfopNQUPZPXcgu0+HnOVodojW
ovPC4XiDMbLX1s9fVjK53LrzaO4VKIFJgp9Nm2OPiZW2mgEmao+WyEVkvTh4Ob8X
eCbn85WdrKZQA8ZQJrElV9sZvdP9OiIhYTdz8QdfzkYvgYAqhzovzASXR4rWwah7
rZHBsfE79zy3FLluW3jQkokc0zxyg5mmP106690MhCjRdR9XY9XvPYpZznbsaH3N
M8q6jDEuRjeZuZAJONIzOnHTSyQWbKZI/DU6h9RDEQXk5Gg4knuirwRVAqetkiml
UOi3cQgYK3qk4rjVNGispizQUZ2W/a685HEZvo0mHT0rueh13/ri2DDDV4yBjRA5
NSng3BVsggHt+EzfFsDPwtKuecFyn8aSqkW8gBz90aYzcbGVX0fFfpryArmfdbHU
F3oy5o5nYPVPcE6qJkI02v89c6UEuriIoKt9v6jaeFgxc9nncMJt/bItFmbtduMn
0ilXB2aWI3+SRfziF7zR11zodexAQtOu2dkbs8PAcm9KIRvhNnKs2xYWabYcSubG
ejlyzmXwqct9uS2hXv40RNi6XTDgzAF5pOPvrBit5gIhdNcArNhYGkDeKP9b3RDi
i11UmjaU4GixqMz/tjN15fcIdNHa5uoHeP5cSFALDrBNT7vgFIBNQGgaFcDKOfGq
2bmKhYoIjmfqSaLmKp0GDQGW+gA42O4gt+4cVVLhn9x183UBdrsou7SuJT70/9Sj
r/0m3DTahUWz1HIk23IRNO7yaIgK2dEnkEWUkf2jnFnxPZrh/7Q5CZfUdolHwHpG
2BYIZO5SZz1L9E1siP/WTsMW7X1INOAiMEcH84ZUBZuFCPlUwNyMdmuXS74yCDYW
pkR3wxv7PguP0z+QS/xJMVvxa6eh9FcFiH3pVzyqTcv7h9DxZdt3ebX8yrFrX5jv
2OEJTCOusqNoA6oCAxTkO7EWtckMhdhbiVPisOyy6GL5UCbkCOyUr1tT63h2L4E2
3kpkaTOLg2oMGWDRahK5uW/4nGvHOKlmi5O6+8/+J+ZVIx6FtGbFgJyrHuaRI1hu
YrOSHhEOB0Sex59VCkQGXXdw9bT8L+7av3daXLow2H4xocZ7ZN/Mlt2bCb92rlsh
HF0NaDWqIBsvJWhghM5DN3s3OcgnDijj1SlmHCR0p4IacSSefcslI2LFoYSX8AA1
rwdZNf9ZUd3kjvt6sVe/J95b+xEDNTR2JmvMHmZCvHHOJUMeyDBmBRtGZu93YT2V
SyoHgybSEnv4uzqOKRaTeT2l1xyOTiav2zBlHG4nvRBXfswin83JD8uVVbrsYUXf
/JWIEVoViEUYqGl/1Zew+aVGVl+JuTAxn7G7eREKEo51RPji+7zn/c4N++Zjf7bh
miCyJ6w9GWDD9qlZvZ0HyGPiJ/foi6RfrNq3zC/pBnh3oJvMP8oxPvu8PBhH4m6v
pNM9bXtGWy7NxObXhzxYmhClk5z0sfFJ8bJc4z9vDlDUi6qmt4SM4UI9Xgjimw1T
dNTqj1GzM+vMXVE1VLCMhOd3sqj+kUmZwu8ckRdyRN+qPKw7E03FuaFHY0yZeHmU
Ps3Y74ty80T4t4qkTJaEUe8mrbnnFC/APe5J+GQwtR/8qGXRr90XrXok/yKJBeD6
CcRlwySSi8KUIn4lXOq64Lpg9BkiMtFeaA7KHoTDXQ0NW1Mv99t74xZds4fjNc+h
k+OEqetbqCHPsG0cqahfk4dESoP44vIwNYMULgftBkDZ7fhHpmPLrxPL7d16gDtl
Kng528mvV8Nunv6k4B2R5+la1LQ7yJ4jiOWh2He6eilBmM8hDnFuseJHvR9LYGGS
qom6ih5o5PVjLEwWYXdIEOnLNKSWX8OnNPRwUKfEmbAwo5SDgOQWn9aF05VJg6aO
QiiJcVHw/NWvedFDA8cDN6GX+WLCH0bVc1g5SXZUv9kVT+ufh4UWTnhSCj6cyok1
Y8tTu3gMzWROkxobsUPeS5CMyPagqxnOlpXx0Mex5eHvaGYPJURYIVDus1Ro5U0W
HiqSif0LLwoNOymbNGPW9dfZcxZzKH4CzJ2R/SsYmsg2pbDDaxbFDWzRS5/XkFCR
Os5WRxWmd0aV0N8M2OyH56HiAOXrUDm8rxlvpxRu+VZ1ZxZZILzRNFkTRu5lngCz
GHwOo/iVJ6WoCnhgWPmrVgzS7rvUhi9rLSKgshrafOIAWK2mPFHNZKeJuIq0PJD5
0g67EaNpv9W/1WQ7o/Oop4ym6yzKJE+QMlnuB3S/dHMNQxgi7fvZYjJMBsgcrSCL
5ruoBOGRUkZbeeuB4WSYc8vL3O+Yh4UmZV7L95RZEvbluxMyQ32pwWQ+X26Tg1y2
LhwoGaVUAHj5bt9jkHvF7Uyut09Oif+jX2B34VYat4aIHsI+Wojiyq9BHxzgB+X+
BLvLc+MnWRg+F0T9KURx1E9gmqkRaU5fcNHIdPJOfafGoljQnrEz+rN7KCC/PuNL
uKpvF2EHRn3NIukL7FF8DjfIpaaaAJ1t+qccM89wNedWnvL2QCTsV8eoqYnUBoIL
PLx1R4zUTpaOf1jV3yLZMv4Vm1VZnN5PjiL3cGtke/rEY6/a7jh6IEqwWMX0ZcwC
Lv6yrEN2E1DgEGvW3MSUgCs8ysNfdJvaudK1kirhmHnGU+ZU95ft0+J9GtR5CGyz
xH5FaPmDJT9P+klSoHoutRFMCbwDMfss8QXxPKrqRWSbhV/5t2xw4t/puPAFvz0w
zIMxH6WEjQh575qYC2u1LuB1J2bjQ6ogsYCLu3aJWcuspZil7b6Kdt5wSm8gVYkl
WeAJQvyOKQ0WYEA0NxkaV1IqONNbjERjZA9S/FQ2MaaHwIzUXKDBMw8aVldHOY1P
Yj5J4WyjnBbWWNohIVyoa2qAaJJS3Z7cjuGqXx7iGJG0O0pko3O/aq3HwR4y5+Gs
R9TYcGxELw820wvVNV92WPXPIHVwBGq2X+5lCB3oCrgpUlpQEtxUIJumuJn17xOF
bPs2xw69WuLYKNFgVjRuZ7eEXcEmnm6splds2u7boi0Md8i6wsAKp8G+Yg30Iufg
fdfNg+coJiKAtEVCCJYV+2iww0/v+uJyRGw19kAlbkSaz6+jaea4MZUWDLKt5B1F
4+BcHKA8SRdP8Yt6hI6AlzEAs0gXpx9T8CXuYApf4l4yB8+6tVtJql992+ePWyV4
fDfK5k0qVB5ujE9pSLuFokt2wsucaCc5b79p3Esk/vGJZr1+Ny6GuzMe8nMWphTq
/6BQeAVvIYmrbVjUQd2i10G45mAY22Zg4O58p3m/I2r2AF4IhKHr6eRYjILC1zw7
M+qVbMp1YhjqIzBah1dqV8CnZYBE0K7cpEzez1+31wknPJxLOLxe29S+n30MwsoT
rOKd/5cW/1HxSkSVm/Fl1Ay0txYqKimUxTVW6JHH5GvUSy9jRttZK3FfW6Mw0kO5
p1DWhtIUqXODFcIZNHh3PupNNIIbSkja1miwi91m1lET1oofOqPU1oBVdyHAOpKG
iRLJNO9iyJwgFcomH5+NaxJMMaMKV76/eO07nLFkZfz50mq6NS/uBZpiku2f9Gvz
/7uDDQ/vlz+2ojUJlcIrdCr91+4XJI4ftxlZF//mu7Ri6JT165qJqoXNzL/yIn4b
qpVNIlXh2HE47Phgy02oO4f1K0QKfgIA9TH6OQrT8VP3oCFjrtNHUEle4gycvJV/
AfLBXe3mPbO6ATaKbC/nfXPzOfI7MUf56bvznWzfbO3P4VBO02+G0Gz8csHdjg0z
`protect end_protected