`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 43504 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
u6n3zq+imfgUTXW1Q5t5Cp+ZBwoXgs0ONrt+a69r8W2+DVVKd5Y0rNS4DSjoPx0A
Ulzdz1kdB4F3Gh3NUsnYH9SL4yenSHgmNDWMnNnO2IRi8VtZKXFlhd2zbMyg+IjI
Glgvr99wsp9KkWQ0FQogJEn/Fypn1Q57mSuAgK8+pxFTGjhCU/n7lsZOsTdXpIi8
FxuAkMXPL6+7t6Ofv86PLzhKcOt2Qu3m5HU2RWOJJ0PuM9+939t43aNtJoFMUEh3
uNZ/BBxL28eT9Hc1NbuaX/Ua3eOZhQJqvSTSAQBPUMYpwzBbA9A9CIDEEP4tn6FS
+HLAapqKH7g7jN3wiTXaQF8SgYv5/oBkxN/BQ5WOzxnJm5s+1A1Hz5I4pvpXpRlq
2uY8uEN/bLjj6OR1BB5sq/4L4boSjSWpPnOyFKH3cnXx3tVq0VZkN6XY0kWlqGav
s4G7XGAsbttzUP5WgJzEteqbKN7KrUVbHCjt19x3j+imd1Nb7rV/4pLZEVtxmeY+
1BafaeWkupT9ilcgK7YEIg8aDKrvGviisAulBEVa5KSzuQUsBggIopHbu9/yYC4e
6Nq5mbaeDL4Tmhc1GiamOuCeRFR5dNuQqdN20EhKMBrOy8ew6Ev6d07FB6DSIOml
Bvc/ZH9QDFfi+XlsJClfMGyp9RyeMHRuiVE7sQal0FJCkSHP2dBFnGBBTJjtJadY
rDKMYrMVGOAimkPVp0nIh2fInjKlkU5hFNZZouJmo86tW8FCvhEapd5PldhRuliT
AWWCiJNZ+J6N4AhW+IfjV4orpP8uF6FdiYO7iC8KiUjHIigMSwf/YAB1ElUb/JE4
80d5Nso+jlMhAZkkHdtOEGVCV7z5UHHlLFrTYhhz7nHAFL8KeJI5OPstoFgJgqXx
pBVgpK21Dw+/IiyRIS7i0c+iSOhflZBebvZbPWmvunOXR8cV6DVLTK6d3up2Kz6K
JqL4jcYe/SR8LHsKt0IqEVEomUlfbQyV749pgMImqFBU0eCibz1MCno5hJglTxFQ
EwvNdOkFFf5molzf21lbubtaVohvYS5vyxR1jxp2gfAPfj5VC3JNo9THZiQavbwO
HYtsyNIXSbOB7wjgkeD/BNxdzRREX3Sf8/xVBEI7JSvjdFfj3eD2BkCGl5Mq3C62
Y4yumLV/SRhVcj3xfIzPvdLSmoz0vKlfDCeYijKqhumixbCzhUrN3Jkmn0dbArBw
Z6uKGYpn5sff5PIuODD7frCuDt3sCkr15xrB5C4hVhpj3oFSnAHAfCPr4Qvu2uvP
xnzEO3nA7KwyC4iLFp2no7CLRdEWa5SYNiB7fHxfeWho2bIORzrvvBIyevLt5waW
OhTfn53Nc6Wq5I7kSmMu3Z+VSQscrhpH7NleaPb2nQX10XAzVCOQee/N8HUxMArU
aLWxheenNfB1jKY4pNVZiqkOHBmkn386AcgrZ21zu9sCqlMoeFAsu0NUJZVZ9Uqf
KH0YbP0M6jqm9k33OYMeHms+81rudM2dRTx7UJXFRUrMrTa6vCKbx0sc9BfR9fRT
PcpHPGElP0TFPKVP6j11p/Fi99dALlXKRiVxlw7fgoq9BiHi4J7GVFt9Et5orp3m
L2QumLL/+56vi7yWnVqI3XhxD5pUS+1HKr49n0r2WfecKWCwEhBzojlREdkuF+4a
vdjf9dLFGoXMheDoM+71EtzCkRqKPt/PybjwiYYDnaiqg6o5E3ps/ugDWGm143h2
+Qt61T90/13ZrDKAU7iXXe3OlsavkjI0hD9Y8rvjtwIvZPWnnJcArcmmbR6nphC2
gs/vB+2s9l0k0UP5VmBWjuJEaa1ZXzjPipJU2XPgDdxvUI85vbgn/bPXI94hJFPj
mwS2Y/wL3gpVX7kQc+Tveoo78ViWaFgL4O1WKuBrEaBcGqKkHaK3CiK9m8whNAqY
pYlG6STF5/GQmUqbW/qn/ljTfhqgT1Aay99Vx+wERuUsDbAgP4N+U2yeD0s6ruzj
4on+WwC8gfzzKc5dqQiPpue7VXY13p2QfRh1+RZpnG7PXj45MK9Yodb7cOKNkbCQ
tmX5SMdQFO3IfB7G/v4v1IoLBxmhxW2ULw1ZO0azwK6wYk0pOe6oDjxTcswuXkUf
h84Eo3HWouEua6HWOCmHUw9z/DVPLl5Fh/lo5G8BVFV9RCPpsH23AovpRmjDZkQQ
bDeTh79OkjMnD3NYTEZKXDgzVngA//6CxU94HoeIj5JBrup/JoiyVxCE2LiMwwhD
lRSe4oDNvsS9bTPPzaQUXD6JfmBWmmvdmm74t96m08bgk3+9iqLDcdKHTmgAgZJD
Ls9B2vqWJvoNkqDSLbxyiZmyb+oTGD45XjmN5WVKW9nss6SqMShi4HTYiOG0UGoO
/kP9iM/Ck/8/MRX/cXFuSzfOmlKGaUWirIHupX5SWWUSf93H/FTzrSxuxO5ATxP7
5ovyL6lPzO4H+rAzLgACsdkICg1IZLISbsCFuBLhz+bNAr1fox0jTcPePMy19wkF
d5IsQrIs7L5Q2LiQ17+MUsPQqJfZ/DF82QzjcYRBhOVg43nwFIpM5lwMZxzVqJMz
KmxaAK5uMAJFCBhly05HCPcPn4ASHiUHQvaiwJHC7PwuWNcPK9j++W5VjA5WbqSM
f6GzvbgiIyw8xDQXGK2TYVTrbzGOnI5pNMEJ4HewT41uJep4A308K//R5LGEOjmr
a/QfScD7Atk/aNl0dGSajAcjilVZor8QOCr5leMyxsOzQF4LyCTm+eGz3qHVCSV/
ymS13Oe4XOvtD+illfbtozNdEyj8agbJBhddw5FJRvsei7RK3NXQ123sV7s7ptUG
A1Jx2DBzcCJ2I+W963jvRnuCcgbPLaoT+8hi18pgDEjdeTMfcYnxsrB/eLLsMPsj
goo7G/KG7WCGcXGea4Xt+K5nWX1FWl/oijDCTGyqcnO65ZbhXcM8L+ZTyMfnFHlA
/FUEyMf91uK4EhLIw5503Z5Tjdtql5GWBUjt8pXTYGf0ShgycLtMmTMh2Qf/Zf/b
mHhTfTWS3txyX9X7AkzoRLPHEUX4MR0aFFwFeyFbyS9yOM7hHehzNUdW3Q+N9JBN
9mOZMtcpVN8DPqn3XGPKVC/RtzCW5yGpmKXzQgc9ekyB0rYLsZA9nZCilPkQiNCK
QciViV6kvlBD215DHCbOzYuZjVtLGDZ/qjdUTN9RWtONI8OaeoyIzhnF0zIYlnZN
P/Vf6EeVNz/Mb/iBL3VnyzBnHXRjvn49xN6o8d6JDZ/1vg+1zr/Vmkv3a+RFi1g4
I/Oy+gWUt/i9x0VfFKDxGk/NXO47SiG6Gw58vON10cSHK57BjvrEFcKBjNnj9dds
Wv/vX8qHU8wOJifx2zVmmL0Z0H3aWhvhRW5/s7LqAJ2F5AUhEnRtyjcQIjdeAjLc
lLA2QxuSJFi5VXQsDCFOl7WPUkV2FpoMfOTkOjnx1WNsXsPOPA2ZZqIOM+EDdbts
NsN2MuX2HuLNBiPoj8vUz/jq+YGXQWWk++2wIHGDo/oGRviR1H7gl6rkGHHtzQKV
f2S/HUBoh/dnhP0CK7GXcvPDwW57J3ydS6MR0yC+WhhdNeAq9oMyYzPvn57PYeLv
kG2iEEWn1OQ2dvKRX+Vkt7QyT7V8K0hiCkuRpx99tnCZXQ++x0ksZx7DE4VEGMFT
IkK6/IAZeeumFs9G40/mV5N9Spx70rrSTe3ZUC9v2EsVNz6KID4p+itMDpr1Rj/6
9BY4IYikqlExN3MFEBcnHSbX+Wr04CX4JNjZT/ySdYetTMj/uOihpXR8hNaHmLk+
rMTagnoiA9EmyS6ImA4Dt2PT+uUNp5z3VG1jyhPU61p03IYvUVnNe1CXTd299EnB
7Rn5UOX4EFgcEAxmcjcowhHjwLGh1M01TxkoxXrS5+jvcOar88FasCiMmPpn7jZD
1O0c3KY56y1crvzzVmfYA2tDrrO0gsVtKF8DqVnpIveL7r/fF86Xle/LgtIPvVEo
0BfaO28HdKt52yqkf9vFzxgoeFpdIA2zjr9fGbFKw/81/omR1h8cZG0zWKYl6NKx
E2AmIB0hY8Fsx5hFKClFA2llfD6x+06SRCkmvm6HWfxv/RqWrKY7VCh1Nqgd2xQm
+cHayjJJSFFbAtboloyFDPq+zqYJJmbWYpo7aNlWP9BFdxtw8G9HSddIVd4nQsVq
GKCBZWwO93dIbhMX3sxGvbFBXXf0J6El1Ind6CvOajkPbeJ6neQfEAIQUSoGu+EH
Gid94/SxMldTEwHICuyYQe/nUOwm0cNTKQAVTwdd9K81SDnX8ocqvSaTBh6/ZBAL
//b8jHtq6TaKiQEscY093ZSpeHkeGLZhk0DTI153+rEcJ8aPz0E1P8x+D35VSgt/
RdlbvgZyXQvReiL0UCynPusilviZmy22ZySk4K4qcSrt8u/RzZ0Vi4kBvb1dtq3y
sV8OB2+VhBtY/Maf76da/k5Gij3ZRdwTULCSJw9K8xNGo8v/Z7pz/yZth7r1NpvG
bWhhVu+VwSAQQ9KYB7e8arYkwtTs/Gt5ra56vOQ62G1YSm6CKZP5hEtw/2XN3AMC
3Fa3P9V6e7Dqur6MGT1sfimX36gSgfT38KWJO0LNDDMNCTGJgoWmH9BnbZmJTMe9
E7Cs7McHDNF+X7EC2a3d+vs4vq9ReqPS70tpfVK8xscrmJGBrgqxGYl6F/ll9elR
ZLJFLYhUTeUqtdAOQmz0Twr3SCRP8y3rvnmOa4HzdYq4yebKWFpoN4vodKq3v+gB
X2f9C9fLwCZhfH3/OBEncWjplP/GQJs7ZBoHCneY/3oDKm2T+ZxNZAlBjLboz3DB
VjLRgw4RL1lwxxnsniAMOZfQwTpFzILythl7pCEtiSsXi5K2ln/X2ZrCWWbuj5lL
RbJVIoSSwl7yXVXENXiQGkcnFX3FC0ix/kA9d1AGwOT2ruV81lkPTqxnZQkEDpqB
wqgXUIq5EsQa8gUmlFDjfEZJMYRvVObbf8MsGWUJ14lBesVoEtJWTKB2gNsl9ZMd
YIbpqtQuSmuAJLfKbaVqivAJrYnQhr0+WWXXqKArQj3QR0FkvQLg5+aYHmJZq6+A
uj0hrCBOykynqWm2K0OBKqJJT91xwZP+0a1zHCrqZZ3rnyH6VRDwGY5Hr5l0C59h
UyyLH+3+RkL3CHwRn1X8UBUlbYYo7bpDl/Z14dw88oiNktAjaiENBzMIq8XKOUvN
63KDRYWG9YULsV/95d+1JVNiUBA5XLp6nndJvPLFN9wBazZntqDDjn+fzR29w/NA
O/z0LfT7paHgQbc61ZQy2/AMNqFh8n1tKMFUM4W3hP8dNq+RUiqZa2TrpcFrJz49
gON0rTYZGvS+/SrLSK34MvpcTJgzxOOf5PqXoIF7WHzW6S+C6ZZQl0OAMftKR/t8
ennmVkJJO0GtRtCHopcjY+dwQB5ooDN/Iu3l5V4I5YinUxsWQiHXswKKl7TJiUMr
2LpNrdjB0WXwOPjpAtFI1rFsKcJdLAawS4h6Fi578++TH4OkVrdK49QGI3Nlpv0a
vEbAfMitws39iX2urihyRpmYZ1ChF67GpRPlRYovvUmylWREgYDcHHks6w99vukn
29hxnmRPZPJ5DDgVae6QNhPr+2uTtUSmSSU+5im7CcSEXb7RgydDPSj8XldmYmHR
eJLL+0wSTcLTEvKrt4JlaUEL1lAn24uR+q1o42FVrgZv67YuRAYepxP6LRHAmOHz
A3ZV/ItoF6BSkkEIgyFh+v+3zfudkinD4+oqxeye3qrGQs1q6quxt2ieg1wyvsB/
VOmabnKd1C72Vzda5cdzBuCs7Lk9F1SNJmAmN7qxZta47SJXpfNKyI7nIPhmQ+xh
FejR5c3x5ZOzJnb7NfRm7EHz7RwPsQiOZYCiE2KR44H42+rWuqJEpfH1xfqv6pjm
gCXg21ogt9NVTgZfpmo4PWXsPzvyHmsN9FvKwVMkUvsWyQI/kQ1b6E1Err4urYn2
XuVXQJa9XX6zJjJ8jZ+1qPO+Zfw68Oexy8IJMoXPa3TgY6Dcr7bSmOjGGKJ0ed55
jap4p8i6W4fpzKFezCfmt1RhuRida5jG0qpLgcQw4SrhdV7z4PQvfgCOgcTYqOwu
kMFgaSdcDE/9UqHHvObzjrKs47nW6H+2UAvzBa+zO29EsnwqFGGiZAY8Nfsw/dC+
ugihAYJ7R1LWJT5fzucveoWu8/LaawzKerdO6U5/YgeE8rKlH0T26XLT31xi55WC
YBf+iwbEu+/SgsBY03nruvD+Fbm9mngnoR/MiZPguj7Zov9EIJ/iJETlDPZE0M8n
eIlUVI5oFHeEE9j6X5JnMeeIDVAMvzQmoCV4x0bXEnRYg/NKBFCOWv2jhrUZJot3
QtTra99Y1fU2a9GmazlLcqc96ntvBQDnNdC5QsWCfFGc9HyBXdwYzjGZKudgZyw6
3yydMK2Zpj1TfKDxNjoDtYEtXOtoyMXl34iOQFK1TjIOR51XlqWZZEtFpSZK0fnX
JEo7HS/YFxCM8g6NsTG+ecTAFYdqjxpyKRTtpwV9qJrHRRBpDD3ocEMLuNUsu20b
8sUWAkNo4JkyoQ+SbqOuLM+FdYVtQgJTQWHyCUjj+hdVYGtNTXo+pVmXMhtA/ICg
ei6jziXaw8inkKUYITLTZg8xSgbLECrAm/+52pMHVGGX9jDSg6bCDR8seHowPZZN
mVlQIObvLgb7KWnBaYvCef+i4RSV6x0c+5S7DbVTowabEtnnDtqd0NhIXc5kjoeY
5yROo3h3mevsCBpaw/KvEw/8FGBA04Mbob9kUtIHozvg9aapRJJX7+4a19GxdI9U
AjnNVCa3ZqKpo3U8eUxMDDj3jrU0uxxtVuGQF2NP3EOMC3ohDuJu7knqBZFvinFO
UElvYpTGwIUFSpyULe8MykR+A1ImQ1YjTgIF/4xv6yLhsDKXiEnbHvWFkpxFqzxE
3WRJkFgZVzQHnNNr1lW7ljKpIyXRjC3FwHH1ZB8xVIKrKLv6feVxys9WVF1CAP3F
FqG5R+ZryzQYxJGa8oNcfbTK54J8Y/k97PEhv7lepbI6CGf8HAnXueMiUwK66T/X
ZRywzB1MHdck5ukyD3Y7Y6R/N+gnCi5kfEYWk2IfSfxVS3XPPiaHb2Uz+/1CDyci
y0YMQxvNd+04SS73i5Wo3OVFCnRfYv+srkwA01EweT7PlehON3jCZUslQvohKKj0
w3r5kLQ2Dkw/vcVigNcCtN+GZ++5LGZwbSeJQrrmxsU8yJ2nu7XhjhYu/6oT3Uc6
cUXEc+Gb2TwNVuYQvCLe5S8H7c28RH6wNTZWrvKdrzp+7ky8BIxYGfK96xu0d+Vt
sh4KJZx6gZosonOCp9x2graN33GOVjWIvoyGU6AmsiasaYh/yrvZrGSXSiBj2AAl
yhOlOejP1eKjvzU6W2lu+qujlbZsjkG6u0y4dda6t324N6pv/TZJKsRzrh2wYlBs
4Wz2bWPsPR2Q971te5UfLKqPW4UhcfFTD66G/pb+utKZTp39s8LslhB6zjfukDtC
Al78GwQ7yCjwlZtH4TlObyRFnAuYSLxHKSC3+7iZ0YkvAqWzl98M6vRrlITlEHPy
3s4IywqEop5860rKO/J5fDN+o4muMA7+6BoST4nc07dduhFBZvljVKK5JDiqM3+x
4rqA0sDt9Sl0Tl752Oby8htCKTf22Weh0HaGOWi+gYcCFa4Hciss+WNvZ0yK8EIL
hTm0zf0J10+gDc6mPlMhJCt/dzAn3FSYJ1WLf8eSIdU970Tq3BnMv5KqKreuXvB1
T9ZsKmfYAenBvakbosMT0oCCRv2hVKqteKMzSjKAbTw7Wd1ivbz1Wu/Gc2mmDa4o
oe2PJHt5de0Pjsdq9dfQN4+kZx/S0ZwOoGfU6/690+Zo2cFoV5b+dta066/6a5+B
8KUZS1AJa9brdpWH+npVzjbSxmBt28ylTEDRccUau2jRuvQBzHK4q/LzhQQPI+Q4
kgWYcC6fsnfBaFDu51kkGnPZubXIqOOAHpPEelZqUv3YFHHhL/bYuhXGY0aTZi/9
nYkgtmHEbvZ5yeNjh1fOEVPhGq7Xne5hUSB2hi4bJCLXAbIysuQns2Q3QAV+mjLg
6d7f+P+GDX+r2McxzxqY+N9N/nk7iX7RMQMGp104wqCB+R5t8ce1UUOVPfHIn4ko
PTSc+cW4PKFwB1/8MGYPJC2arcmdPjF5LtCVtHFvis03GUxSH7aoiipRi1jvbIfs
dUrhn073mt6dT9oNP8fYmt+IAClF2AlrH4RPtyLxUOnvuxfNEWtGMsRmI+qfTjKW
YrIB41n61lo7SIJ2/910+jy9urVs4b3G4j7ZGbbjMlImgKaSW4cY5JvtzRnL0NdS
y76PsvT7ri/YK9sPEtp008rUKfl1RhlbPwxfisc2AtKD48gM8HuQF9f7jIH5af09
rUZ7tp6Y6aqvAGcvIdLxfAlJP8y7+TZtb+i6M+33a8Dgnj/mOTOPum7aVkwQwIKB
u0TOJgpMOSF2+kdaIGZXk4GEITTzNu0e6i8ClCkGWIyJbiC46vnSlVodEk76rrcf
y77WPHBQhdyoiL4W/Abo88uHrPAxR6pNf/q7g2mnlTd6MNHlk+JXN4s+X8LiOWHE
pdl5LZRelSfrRKPHOjIzybwhImtrvuLejID4Io1u/1rwgKyznrWHMoaUasu14PrF
nRyMIyWRIfknorakXsulL8Ikqi4EeZnH9+FT5tDYdYg2jz435hXpo08+hgBlRpjJ
vED33QJnYeoLG1+ftg85dXhAjgw5F21mj6pz8Lv6Ppp9813tHNJ9sGCeW5Js/iKS
xDRfCvqMEP6M8zfwHJDbvFmV/ZI11dQnZPUkQ3FDf/ifJvJTP3/bUh7QbWD8vXAm
tjrRhc/u2o1bu3eg5U4D2gHjeTuXH3UV1peWRx0HcqgEUsIWIWf8q1tgo5s5TAS9
0v3eIsL9zuQ6/fIxsIQV2d2UgLjAk6FwcxgiqG3EVhhssGm8XvNmkohCYCgks+IR
wtFgnPyDkr2ux0VrOlrsg7lw5iVXs+Tk5I/xGFZwAhKUlaOQ7M9poQo87HHHp3N6
kfVv8wJM58hkiwa7cUQ46kLY/SPPSQjGSqx4wWRHLwwVFtytmAvIYpwWz+tvZ2/T
dFELZuJ588nvVzYW4nrxfyR4G4nh4pWi+Fi0tNsc0ruwfDa5foODgExKNngHPD7e
M7rKcTTLOM4+EWlYCdiDwMP3HCjW7hXxuIbVeWPnXzH/l/ErWTID7VFa/MXas8K/
/Vz8bn0in5zEwF4S3ejqn+7iAWAeQC/u93g0wFWcpYV5YiMC6zhf1yEhMWLY8j8M
rvBwbIWV1lUEycZ/QgpHERP9tIQtPJuyoZ5E5LEpOIAwKNq2W9GT3fIARcI68dgy
wqRo5s0+YfeCQb2KO16iAj3uw6Io2b8XPhOf3D+N+lrhDVT6hlycFpTiOTU2XJrJ
a0V/GL/iRMe7BLGuuxSvRH8vJ61p/KFv11HNLE02jwEde0pQBZYj4nynmlwehsyz
/qol1YZARmw7PLb98i+USxWElcCAhJJN3FTIHZPgiCiiXWC4uQVLM/IPLTtQO1FD
hfmITNSXxcUTC5VVrV1WLIJlkXLHteK1L5OjGb/a5deUQs0mNo0BgbESjYOE6Fg6
zbKwnOpR7g71aFeuTgKpdIdaepRtd5YkSNFqEY4DnHvj8MYmzIBx+DukEvevxcXa
2pt9BBrPCWWDBjdFxW3/IByNb/K/zdlLS0pI0TyDrJzo9mks79oricLQPBrTRQsc
OiSEFyf+9LO9DtnKPIMzb6T/ajMF6Uj1NFgOX2pemM5vds1rew70dtEBniTNxxC5
h/ugMgnRp9pCDK8MI5KcPC2x5pk0Ifj9i6bS6m6ET6fVRYwDCKOvsw2itlFCv6td
D+tAPMqWsUFwNCXfo+FLd8dJ35Tj2cVVId5P/bkg72EmtTz810hnAuU4Cw802wMZ
WbF5jtK4065kEkvCqgComfjSFmpGvXyhCt0+bbIAnwdWXQke6IWKpJR4An1mVKUJ
hgFvdFxbEsuxOEnmUhsSL4sosXQYIohgQud6q7hGVR6Y5HUJKeZjcgni8g06aZB7
M0Tnd2YQgaPl3oYJzbmSCjXU9BBG91epgVBEpgq45cmf47nW6jmfs9GniTdsegJb
1TZWxDAb/99Rjr+AdQgn6PrAPyRa+vApFihGUOicwBO2mBfVBfQXzYELcdWqGF//
4SX84s1bxtzgoP94uCslc+Ix7x67UfmS6fEVSmLU6woiWSLfv0FwhcK4OWr8zk56
l2ZJlyYl4Cra4W8x33Pld5fWyCmxWpEaGrWYsPPdKUvXi6k4opNGlA9lSa/rMQY4
a51fCe2ao8VSoxHvgzojPPB79yZs41rJ0Nbd+yKcCYBcEPBwTpyy6gYc3FSwN/6B
tUZ1G96a+Kq0R5B5qMcLE3l1WN2GDrBelpLZVONFrmDoaQiaWAq3Iy9AnmQ5tiJw
SLYTaof/AvEeho6aopWEa1chabVDumeS40SEbObBE14FmH0DtPtgDUVP0dg7mUQF
A10vzSP1XuJICxKdS1o2+v6/E6QuUQUGW07JjUkzRf8dyaHplzXR37hAfQcDyMTp
X4EUrzvcIJBSrOLjQQLwOdFgycjGkrwUZJf7ANayL/2fcCz60rk53377LELXP0xc
6URgt/QtuUX19/Gk+DL7vtljGD4RHj/BPFrShtKj9Qr7kgdPMu+nhbVyV2Ix1d7W
fDJ4v712qcs8H7DKMbsKZ0S9H31PBuq0NJw0EnCNNI0XuLGzHbnsy11zGyPBUJnQ
S62XN/NmkBh0J1blRT1UG3hrkC2FBy1DAG0aWIH/80B4lw8RJeCY8xXu3bnEv1Zp
QoIZbCfv6gp7jLsuycV+8K8f3fGPLaxy3ZVYsnMz+QQFJRIIgQRQQFPmdZJsC6yg
QsbLdgDMnFXVpkdc1DATRH2WMdxO0ansFIVKYqlktCcO6iIwdI/jTG47BOViKdiI
pxxDiFZQyeToMusT6II5vQDGeBBhxbUxh6rFbN0gUPxPMmYYd+lgRpR606e+PSB0
dEYWw3wdQubioaqiU0uq+eFKJJY3jFsIBGPRREG5t+k/UrpDZIjhq9/ePlI+7GQ7
clEOSMv3oZ8Eor74mActn2gS/j9ql4Cpf5Et5AI6YWevKYLwjv6DOq5/T0MjPiN4
fFaITHFzjXhM1W9FJueEsa5elaxPaPA2D4Zpyf3jeswA0NDmrXynu2EmzD/p8hnj
dXppIlfwvViG4b8wJVN66OoHRRQgHWdmnvZFUXlAQgt8UdUFWX60ix1i0QTxCIdh
m6H3cd87i48o6ZLW+3fRatSpv8FyP8ne4cZBZ1i3QCtKT22WCTksqm9HFQhTsI3D
KJx2HEyNqGBFVVRN+w192tLQhmJEeUQwA6FBz6inaG1m+c2huFI+BelydnH9S9uZ
XuGJH7ycYYYZprtdPYUuLAX+sSnT3fo9Q55OWGWhR/Ugsv+t1PCqXiOn3+8vI7gZ
bR5KPM8NvhHg9kSDJ6DASo05yLIb7oeFioUHpx00i534jYve7q/wSHynO5kksIQI
GZ7wn/1iDmsKeAg0H96oLWOFy2F6XsNqN9lApRkol2/wMWf2IMaOUYaDPrX+BSw3
vTnV5zgJ9e1zkmduKtbeORhlOQqY0zqE+I+2hSarVJzNgyzqpNF+wCMBfx7oeN+G
6LpNa3izBQm1fUEv+g8Mn/xOuMInW/7flc7fo9w/KLGWnGIGGXuhEGh9S6eTCW5X
IyuBxTQCLtHB94ayT6a9iUwtD9IlQgAk7yTRWMYfwO4GJmjn9VSADNsOMPFgDTsR
3I4FmIVbqTYopNcWcjnjZ0Xy/ADFXNdHKp4/d2NjXuvnfIJWWCC0jzOMSpXvsnZ2
CMmf1XtptCxrQp+tDMOuMWCoQATntoznz9sPlp+Yj2I9Ipkhs+B1AHzHY95BchGn
2NGFj6pJgbXAChDCbDyFLhRH1Fa87nx8bj+YZQSJndMUDnkAe34J1b5cdUqsWqt8
Pkw23MwKGFG+/OXL7wL+u04/olMORlcoj2EY2cOKmq+5Hee+ItHUdy5gLeviNgTk
4C0k0nM8GfOoAYkTir2Ma8f8J4bthGX/XcPjEUFg9fZYJIFuBI12zqkNrjRjyxsT
lHVE/z/di0aqujXVuNzFCyoDPtP/RF0IXbpy1Zv9cKXe4i6dsHYEwPA+lBizV+2A
3oGLwkyEZAbEeYiLBTfoJV5Le7pwAGOGhXUyVZVN1/7VRYqJp2lkqZEM08sOGr2D
uT6XcajYFfNlrbHlX/2NqAPIyFnrcoXCrK8jLziwC63lsjH1rv++Z4xruL16VjRF
rYNwgPg0889DHVtLuP2vrSeNsSKk7+B3xi+aCkp4cN/ip7UU15aWegesS1z7mTtF
IETtHOrD6yUGtIM/iLpwBgwLT212uorTNkgP1uy6n7u4pj0AO8kO6IP2WuQ6Pkzc
PeHUndp+z+S+C8pUu/i9GqkKaDPKyECOcBtYRpSTlvBncR18ePd++IvDfuUvfpsE
iKpd5Ld/edWMrKEQ5gIxJoKqy66/Xasg4Eu71tmeWRDkdyQ6SGTng5fknhIIMzA8
qRkrLthyDK6E6gIABmstcKj7YCkiTnPqms4Msu1TXK4EccpF5zwEEB/IISwoMHYq
3HE5lHTLQWd7oRrpCdWvGH2B6YswP3u+cJKYn95UeEzDJPMyz8aYpr6B6znwU9lE
ntiVAUdtfi9o5FuqybPZmAtrIAjLWn0ZzBEONOnCT3eqUNfJT2oQhvdoRwXQ14x1
0/119boitcV4RRfUDqGUX7XDy2GrCTUPPyZj4CrxMsJuJppAGX9E0vEbOat0Y11G
vCRNGdkl6xRrKvJcJxaCURLxXJpCrfgOosZ6qRPP9kazH6KxbM/a1Grdw/q5YCkz
xkJcAKeqEh/yVTx3Ugsp1d2Ue3PgAr2STQx/8ycUodmzBU82TLq42lyGm1ChIGyz
h5z9gcbd2d4XQtIOoiLbDbIcYiKAPNoo7YKd33HFe73cIZJGeaNRYryEbo8fNUTY
rBXjTFX64dMthqkXRw9sT5YB3z/DCoybPNlYH3S4pwhb6xWwHvrugdVRKVrG8CjK
prO2YgIxNpLQcFB4XhAgZlNslEYM6FtveoHVeXPTPyAm9z+vno7vBNfaW/tRa9+r
cqLO68bUudLQpADHpHuLkGzJJa84R5OIz15+OtImtkSbwF7Q0TPbqIyqgauOAJY0
OMa1NSClKEIgbFwuW1/3+FQBhC4ZtqNGtbtQhURF8BKvz8mzQjuEzLc+sko+kSh5
+a2Ko3KXdUbkdVxC9jzzIgeeonzoArqfDymXTctjtPEscfHCg3fbDHhpH+267N5J
ZJh/1gZARfva4VCLKYaVkVnxeNOqzUNmshHM2MS23p6E8qLYHORoa7+KbP097ocr
NSNls4wu/F4umyY1FQoteIQDzuSbe5MPQWMxpiPg9PSALHJll7CoqQRh2QefH+VM
y8qv/5ntip1aOoJnOem9xJsQpNosV3WrCneyz+ZPR76XHzCbia9/2dwiv58X9xcR
k3bGuHy/Dl5d8U6t8JwiuaBAU4LGV8BH779bO7V6H/RKujg8z8lrUoHDRQEPqZrg
q5NYbduzPc2AuXU9ndDRkUsyO6+rezZHu0C2vREXer8hD6qKAsNuKwh/rW+BqutT
i/FY4V2Y1Ts00l8w/jKNwY/hXSvXPS339dZVBxZi/dhKt2p27YDHleq2WOYMYBGI
kFi91YxibjbRiRff/aPTbyK/XqPf+OuGvU7kT+iDLJnacRHWlPrhxqrTJLxbSe25
87Ztf30tMeW5hvMPXgz4Q9/3odwwB5nRtVDIhM0wvQ3uBXmCkPYrlG5kCeHOPtnx
Xh3B0Rtkda2shdKlIEvEklH4LiXv1n4lzV9wB3akm04IR4NAPRYwX8GzQr7HfeBf
alWxJO9e7FjLj7DZbuHzBPhLUtplLcopDtPobhk6Udns/kTAznIpzsK9OuzOTZbW
aa8cdRxVMQT6R37sXNkdfjP4O7bwcN7oxh6rcmt6zfk+yZCY2iBnki4aOag61V5Y
FjOfxrUPJmb5nJRjMpGILVv5TzPUq3oxXh0VYEpl0Dvpz+FRWSsolgQs7nNSfwpi
J9hbru/GmJzQytACq76XINFJiATx9olgA+DdkqKBOpFtn/UExZ+vY3HVB5NnJgph
Ir3oFQALYaxgn3AOAQH7CInbnk9VfkP/UyHj72jSAhqRGvZ9O8dFwcW9dLyeLTd5
U76F1Hd/eC9KVznsXQ6Hc30dST+9scZJ7MboDDtuMpVksL5IETagVUTiMFYo0/+m
UdGOkz5EHTurk9uDfNR5vN9nZs8VkzBJnE3SSNlKj8GURIF5a5Ti0gE0cEgWmvnh
g5Cv/Qq73VEmNPNCudMi86y9yVO8jr+7BFMJMgrZsrpC4yURtp1+u5Cn5JDssNto
OWZ4ispqFI+pGXV9OalcXChxOHYfT0vD4hMcv3szFaFvEpi5gK6z5Kh46zQsRbHv
CrWwiFZvXoXzuywB8BDH5R47uPbgxUrtb6ioeqhq033yqNmU8oItB30wepqoZ5ll
TYIgO1G/jr//wqDCJuzMwxtpPcn1HPtGZ8InFdoi/ijdn8OYsekye1ZEOLN2v0Ku
rSGa9RRug40baM8aksKEDasrfKY90xGnc0WeB9nOpr/tHdUFOf+cD43Ex8BRbvB4
Jfvc2Puui/hqRyzWpPka8cC1EdCeo0LpYC+mHzNAAHccTS2k2wZIFr2ip3XDJX73
kpt24hx0ZceTJxk8S+zRoKN9pg6TtvHJFdyXohZ4vMiIsQupyCMh8m37Am4r9wMP
AGL02s9IKtceZ/Yy/FGdlrhn9v5iPw1LFVOTREI9X4EhfJgEvfDz5+zIdDGUsZ//
N3bHai/bQDC24OrSJ02P8D2v0+fJO1PCyQWpSwnP/6wve7gLulpgXDWELXIx7Kvv
jpraigaxCqZtAFOH8rb4tIL84tpsCwP4xxBMQXFrulD1V13gOSmkql+QMY88h/CE
bz8lkpnMcc73SJuUA2cXLGLh0LjrP0vz7EMpkJor3qlMy0Wu69uWHOTViAl08KAR
j4kqMLZzToP/onRJ6P5oKHIVqZiftQJyETJTmiLlrIatvxJiNG4jesvPNLSn/xuv
Gi5NG2uzeQlvOoaBHsj39YyLU3VsWU1WXWlXF/QYudcnsXtJO49uDl882FFc4t6g
uvHVxSHKrSScBQ5nBWGasnUxSlInYG59DxfcjW22wBwjKUq6vVkETj0VmHa7MOpy
HevC2g7KjRJ7lY9RG1guhaEyjHW+m8tv2XqT4EIy70JXlK+sOs6W9J9s7cvdmTO5
cmMER6hHpT3etxB/btYw4VbHrERMTBQvn6V6CMEc36cuDzKTaSE5aaNN6Xd52f0H
hlyJi11LC43Di6/7WUZFdC/foToCnHbjR0R441I/VR0980q2BMrNaDJIPSkHmWph
+2UkfkIdpdf+Pk7bR8TqMQXDtU3vXRZGqF8rYTodi2cdwG5CBO+1/KBiYE9IKLnN
+g69VrJlN9jUtOoe+5hG3WPXllWxes8cXe/b7jDWpejz8ZNcwyLBzRhkyWWeedwn
B3OKnCHQ57DHZXRN/zG7Inn/ZmS3AUXaOkyZw6v1NvYJEuW0Dng0QRSyLT7/3AQQ
AwE9v3UuwyXw9nt18ck3z2B8P19uEg15z8rz90JfO2g0Y2AMvUCMLUj5SSFY/gEM
aGEtTbXj3rT0zLX7X2iEkRkrP43zU0RnTZKeWVaigrP9OGOenIAgqtSU7sOiINpD
ADLv4yFHnryxExngAtZexwyq7YHkkhKj8BCPysAysWiY/3h9QXaCoTw5EMn899Hj
CBEqhGGanvm3+Rn50EVEDaA/WRRpEOAIrRWPnicZ6z7mhhz8/aWhsN4rXbSQsc8U
WRO6RFFeRuwgueJclbB/CVjLTFCLS+xtfCOQGmqBSAEyxfB7Us1ERoPPgcSrei08
HuaGcthvxO/7Ac1wxWTK43E9wSMGTdio19OBtCi1ZAuR28ga7n28jc4GhKK18bvt
+eBStqFVvTuM37jG3alvvlZywgTuq37DQG7BCabiJ5/SxhkFByiQErpRwUPCTxi2
GZE3ZDk8/puZWoHg4QnO/b1gRfA8iYXXvytt74Vt7XYXkwvMX/PZ4UMMBsDDjQv1
lDYmt3EAlL/ceWfSgi9MTEv+sG29/gbx50z6UyDDkoq8hbun7Kct0ruX0KfFG4X9
e6G4VCaw++UmO/c/CKvR25HdhWDsyMCbofv6UuODcWrL4wYc61pFyDL8VtmoxRmQ
awA8lKQdLhlRUg5wGjQq++asm6PBxtBhngvz6/jKwU65K/Mt3HpuDfOMad2nNrcp
QIZkwh1UhyVBjC4qM8Eg636+6WfU6bbZpon5tlNKBPe5jozFE9SZZDpk1ApVEAGF
dFC2MjMwvylo4GOyeO6EIOaUtK3b4ygUe0g8SIJxZ0qEjvFJLX3d15xaU8RmzPTh
c7hVzkAZqBcds73FClOyTzGYjzglbhd1tGlwa31Bz+rF+msUkU7+caQNGgYMe2K4
3+s4U1+SkOqwCxVAo0d/daTVKjb2bkTkkyVfPfcYZyKdu4SPyiyxoyIZwVU67z8x
hbfZ2V3k9OIjAXbGNY4sBK8PApgwG8zzJ+YEnqjtH6YntCU2MDEqGWAd8r6f8d9W
Ssn/V7e5JohRK6FXUu+af4mhSJXK0r3xxTp9YRX3/vQ2SjMjY8Y3reOs7R2dRtT5
dpq9ETkZHfoM2a7KJkR+Gu9L3Ay9hmRb+C2rNaT1D6DXz2diBgoYaQOx/nY939Ez
ytEU4lbFbOpQdZw3YyVHeqXJjyiW0fWl8V2j1HwlHiTPRhK38svl442vlbN9Um6E
SKAPQgc6zxmknpc01qH4TRVLVdnWhOZRvm7P4uCda2VTC71mgtmmauAUf68Dq4Hd
l41/c0Q+GTLp1YSkC6qP3hBEEJ9x4tWO0T2XwaashNGak5gcc1afp3K9PjS+Td8Z
Wk7W0kxTXLv++DUjRU8O6mCEWaCrrxLKgtWceal8Xa2DxK9SrcxYFqj0FKKGOUW1
8y3emwjnjJPNaeeFDMynSbQ5uoxfQnHsDimBJKamj7jawgDkHXxTIsPff9us7V6r
+bY9Y9v4gwTOquxNlnpnF4iw4yBFSBaV72k6wHnROI/9wvU6b5aup7+ioCc9xIee
T+iwMnXeX3hTyYLjh5BbYa6IxBHdRMw3eXxVvTIz7//7sTjIgR36iOTaq186KxEO
TTiiJZhuROOuPlQC18A3EpH0Ne27jBGe7svHHMvjKf9+yqXdfvpgR5oGDZ/X/Cam
TxrPSmh4tlUn/nL2/iU4gLf5D8+GgRTGxuHVoaWr8IRvKexGSCQMQ13l3NJMXRLH
IwCfBmWGaih+SC0HsbYQSP7LEV6FsKl7eNN0U/hWGz79PfnjdfmS9gc3D4syO0s6
FGkO30RpOZ0FvSmmFMrjOfG4v9p5ALjKtHa63fCdCLT2juT9T1qHZlIYExo2GCTv
PyWiPK26wj9OYZrtPGBcs437WD6GX8AvI22DCi0RC/8tBy08LQ+p12CzQOprve2U
r0WXEZMGmWk65wA2OJhEor4NbZqlQu/nkQkLBCeNDOkbejBUtcGyqharBHizKDPs
tqzmN+3jBY+OfLtyF1oL6V2ZdfeGpByn+cb1sszEjDgCgMdvP8AgDBm3nyYIAh27
dJlRCK4Lni7lRlMPdpBfIpy6mrSeN5n5Hjf2vmEc4DKVvzpZMp7DDziKHjpYNYJS
uIWH4XKUIrFx6U8yvF39lLZEwylIdRN/dVR9Sqc2Ggk+DNC7ms5wQW6wgJudbaT8
gIHVLc/f8XFBeOGQGGzJZmob5F4OHKzNqiWyIhwp4+u1PSI5tDDlWqhdsNOXXn5U
BDz9nkR+X6hMJkbzp450ooyjXYEE5vRAmp9hZEQsfXtnbnMEl+F8mJymf0C9WLfm
cRh6D8ezgjs97C2k1RXiPArmrQ2ncEs98p2J9h4vO+nuKRmBcLI19rDPXjkavLH8
rgu6MluJh+hCUBOakPqsd+FpaubX5IdsS9a8g9jxpupYzkfziyk1dictkcZ7tU4P
Cvht183R/P7fl8AnnJTptVJYOqw8zASjelpBSBteOvDlFDmDSV3dt7NVT8d71avx
gAkCvkK1aGXSlSt4K8HSvWVR0liyP9hMbj4sCNAbOSAAE32cnkASiCLsDout7FzA
S6AhJiO5Ae1pNAbwCrHyXG9vlIJTAFCi4yCuHuTaIYhLm19KaABFae9IwMGJHRrI
ENjP8SlghqOMnpC3E2l4lsAC39CJJsf68bHN3aLRofnRz0XSz55SK4bRX1bdJ5Gv
Z5ZqX/BMKCLNM9gvUJWjBWiKZpdd/8839yQ+5MbRy/NKP9gmbKi7cyS75hcpyApA
W3KcufNSmkLWkFJqZ3j9m69snLJcnKH2ICJy8efNw0tbcOhajSZcmbcrHAsS04OX
xBkMyKgqnjuPyIIVb40+MN1vVrz13eY4p2+9JLWAOvoH/QERIk7/nKgmHOtzguSe
+oylrgZozO4P6pLIV0jwOkSADsmA328g7K448Wn12TQDTSimVBGlxSSdRtaEVXvF
XBFNnjeZnE7izTy/sapE3sxvMgASnKSzQviq8vrJV1yDYWGeaxAcIEFDgPtNackC
6wpYSt18G3FBOs/ThRYmtlBSLtPOgdI3akKRsj48K1ti/NyKqvMYLoZiQAONBINs
VGDzoj3UrbQqtRPIFDd3JPxz3/PakzbiblJgajJsabhhlgTmYkcdiRAuqNuNKCCv
Vy9DX96qpovYnjedtUUzEkNLenjs3nQLPgFtwUIz1oJ6H8k6b0Vk5TegjrOlrPs2
jhbgl987wcj6NlxzKBx+P8+aBkRiN63jz3Z84mI+kEfg1l8ygJbBmgUia/qcXij0
XzitWiVX9B1ZtFJWtmfjwauOUsCqLHIS0fNB8sP2Ltqk3DTN4z7gOQtoPzrLejcY
jZNpKdzLpqrqoQ+j1X8OeXepgHoNhSi7D/aHq/sX0AzSKiHOhAxmCn9D9hbhLMjQ
7mLlMObgPPvdfcnrfNuZVPdy951fd+vO/RZuqZNrx9D7Pl4PyxCzMkkSwueL84aP
ZPv7UgV2AxtsShkE0wOzEusGN7XqUPZg3lhRS25gzf5KIM2Dyx0dIgwZaw2ScvIB
IXrxAZirUcpEEjtDaa9X9/unKPIIGftmA1YBn6jQbccsjwPk2vH+xjfTCJ/CRTaH
ViEVFtpxMgExYtNTqd3nIz+qRVCC3Q9authtuO4Dp/0nji1iSEPNJI55XwuziVwV
6XztPYA2FJqh4LdLfi9+jDNNxdFL5QE1Et8wY1CoSwmshfiOme/ljyN2/v6ZLNge
ilesWBllNd5Xa2Qpfk1SfCRC+uuiwv39/ZdYSIm0blPGEuNZv0fvi+SgvncEI/yV
EaWovR1g+QmJajyAglaNT/J1t8Ppq6Ng4Ve3AmgdK0W7kKFR4ORNhiVQH4gWvTOZ
fRic65xWQCojFLRIgbrZcM91VTfWs7hNgcP87R6gy8RS3UT7RatvXh/+d8wEdzCY
3sEWVLW11YuTLi+2d8NzpsntHmUZXB7GdWNh29OCqYsbAlwkDNMgziAx93cFKV4z
YGH17W8vj8T/j65N9Qt3p7YSsAJAyfZwWE8V5Pc6RkUQ2efkZ8Ghj5IntD+uZQws
k09ReemiHL0ezcEzIrRI7+2Th/Eo6FjBnPtPFn20R8h8yAkTDX90kduY9lzqkiJR
6qd94eZk7q2yj+K8qWqBL+Ive33E22/zPed+YhYhYvp94ZyRkCZdHdFHihapBt0K
xbu/9qGssUl44YUImfSCQhxBEtM4w06zxvy6xghZPZI1z/UBPapixw7z5wBgMP4G
7GaNrH6X3Ul4A38IBFSCVK+assXK0JipFE2lloxgILiegT4cXL883jRE8rIMkQ7l
PUINYslTe9wiAtxPPT2Ef7L/VUEs2Ou1PE5JjheUogZN1dif/0nSn9Y/Y2zcmtUO
Btug4nWtY9TvhZdvvxpKeNnvOc67Mz5Gs3pqnsVOnz5l37Cv2MK6loTSKZYdFYSh
mJRFPQJ3hbONZl4MNKR2ZjIdcD/txBtLpqnZOXRkJ7chFytIKreUU8sUkkQxscAE
QdwtTPopEvXeDzPF1CQKM/LPsGReccdJXogxLEvsD/Wa+xKtE1ShSzA0zmC9uCHL
LY7LYnV+9rB0O1lOwWa2mSXUsJs46YeCol4+9GVusA+vHscsA26D37znViU4phAj
LhJujxnFJl4scodlLoENa4Ug1dfrudJvlN1sgcxCMmsbZKuEVx2Dce4FcNrNcsKY
mQkepjERJdWpKTAYGHbKh+y9hZ/rSPrKQ8d3t+v07Ve87MY0oJTrd/oeALfzuZ8t
vzK1P81ixGrq/8WnAidnRFypXqidlXJObW0Pm5ozBv195X2XGYPpw0t6769N1GRx
DTqyZrpFlosb2gs7oF5HliNaB/dYBP8HTtXTQVm4JbsQBHAr3xQMRgO4SAMil6RG
YFSRBMLJT+0EbnOE5vPneZb6fb5pWxp0z+Y/3zluZvGx7jlirI8iS18DGVsGMkiz
HUUwyy/RqTR8wbGkf1hVWC16rXH64FRwqHoif/u1pRFICgskPDf/bpNwlrpxsuxV
F/nkBBKlX2VNs9OF1+7JYztl4SoeSaUYiQKW9ervQW4TkgJpgXX+isaehUbL1lk/
S7n5DGQxlT46Y9U1XQgraEFpg5R2qWRaEmDXUSjLU4DZ6/em7ynQi6WUJfY5SWbi
NpJXERuXOsyoQsMbNQbvpEkQJqgzlsDn4AZ1QYEbzZSLxmIsblzy4aL/3HI/tafh
XancOHiqUZdwPgJ4p6TigFPmN3jXaIwNQINmsyTZeveI5xt5kvM8RrUgqC++01vV
Ek+p4anVpYoBOUxZp+MGasSuSA0uuLY/Zxga/3uIBSm8aICz7kXFUkq7YEvKAI9C
qcfS2qlBwsyJ8Dw2deoUzp58qPEkDCfkmZJpyi8DHjqDrBlKp+SgAftTkQn+EQe8
E93VjoSDJ7tpERew9ZZSbuwkOU3jb3CYaEDqFYYCHYFaQBSYei6+Cch2Oa1dAU4j
6uOzT2dgSAmvFl2pCKrNajhFclj4m+O+erXqcLLqB/8HxujdCvd777XM9yVfCqqB
zlYQv09OrBJPZNKkhjxN5TRFZOfyLdSjas89Zs/y7R0ukxQZDIjnJ3cTT8ZfECgR
xbJzVsYmmloKay1A6gINzX2WZ1F3nqskf3Ka6hbH9gfEK+MXguU4nTnzTGvLvHN7
ih2ItuZqMqEGle7sDemBuEp1nkjcM7iBh31DORA5oug5My6KKaykTrTv/E0R0J/Z
44qgPQ2/8k16i7JZqdEWwYWY73s0wDZLU4K//gdV/9ETjLn2rwActjMTeouYCUME
WFil4wN8LZLjdinU39UfvQb2aLodMpySda8XawqqHrbSKghqOqobvB2hhi5TG1j+
5WUtx+634Bv0WY3i4s5v/nf5MRnUrryUADZBRR/ZzUKq9sTlz41H4NSzGKosI7aF
dxepBnRS2UylAX2RyCWY5Tx6enyP+fi+bZXh9+BRgCoa1M2xoMOErRSuvH+2+7wD
OS/17u7bG3LvlN5TCGLl6FvPgwOSDBQ6ygf9I90UktNllXZGeb9svE998ge49RGn
Z5zMOXxgkhHc88YQTMwuGwwXm5Ch6xKpPQuXW/4bDWICW5eiGWEaT226eTEiAl0V
Ll67m+dMLDjE0IRZuJKXZ0XVjocaTaCxl8k5h516oZxP5q5M82q35VrClJfxZ7O6
8rcdDQ/k9kdSc3UGSoD268y/cpFa4D4iTDe7PDH0p8ks4VCTctFkHRVkXgDvjWQI
5o6oSAXNIobKYuUFk2sReKaer4PdEoQhIWyXJsUTnAOsUb83MZ4z+wuBn/emTvu/
s+oFoqkLO/ZncvQSpYUxLIpO6ezvQOA1XWapga9+bOiQh4ED83im2JNUdRDubtRK
pHqzmEipSdqJhRrAL5pDR44USSWvWmW/0YTgCFNUkK5MvOaDIJMyK3lYPg0yS/fX
veu0Y58Q1qn9vMNrRJSypmlr302m2wFjlyVMI3b7hyiOJ8foMQ7QTxE4oxPwqWDG
+VWcggMQCYZnlR/Rxs9qlIVkblSVd5P2/RMyC3Jt2z7RUPzeF7eLx57ldZsWMqhC
bPvJCaci5kasApo3x+nfFtNQKsZ1Odaxn7M4xGkl1Q86jwmqvFW2/PgUW5ts0LpC
0rcOQLz40OzUEHFrCSZBB5scPr6JtYp7+nTP1hTmNQgsUekRtRs7PjxwkKePLLlD
lgrP4fMs7UpO5BLwctCeVA0gp+qkZOU6c9XUBL+g4kb5aet9CZoAJStAG6FaDSZA
J1lT45c5ppbWvAbt0CHiiqr+Q2gMoeoyDn6nAQ/BKr7GZyBJKxqHecyng7S5IAiw
s3g7pNSy93TEIfsTMH35iEnze3uE2JfO2gPJXnlGjBXRrhJitX/zjj+LHQZ6CktC
3rN/BEZhwAbJfijaYUY+JxmaGYgYjrypcg5fIunWlntSri1gamVsFOJGhh1yqdkg
l5iFhdgFjkbjZJdGMIZ+4N7/ndJhsbKW1Iglohjus+H4nvW1VkH7LjqYg5dtR10f
U6tQMvhdxs6sqhcurB4aNS8YuUCaSWHGzdvYoZxfuKHXmzv1GaAZc+vVO58zFv87
eYOl6ECL2bQYqbi7wqasdwt7X1gHbqjUSu8hw+taiQSsY7pabTqoGqrZJEs04+5g
VuxM93ORXcRkFzWfcANpLaLtb89BortXQMIr0X8vo4LT7y53xzxhNMRPAt4oVGZy
r1Wtt/EtZLn4C3u8HYGotO68EeZqC5JrlY6UjnsedP4n5IzaqR2HllHKCMOi9t/b
fNGQxncm4GzuSbFxt6MYpl+X6hM4BZAbBuhUDtnYisR+uxywSjVN1TmpEfK2b4Zq
/KORfHhV/FkBB3bxBnWogsXKGV7lVfe+k0Lc1yWxlzkwg8p1qQR9aONSa8z25JiR
Bk0MMoGqo7JROq603c3nMYAKncsoSfgnufEcodmetCu4My7gZB2h84T57u3Ak1ad
7aOguQb3ChDD/ZIePBaccgIXykvM0wP1FzjPuD/NGm2YqbQDrd799FD9Pc7mhQsm
SiprKZDs0ZudLtNzxVXg15PdS9q5hhTfyM+3ePM3+IA+u11ZuVpfgcWtS7bsWuSS
VsZ+yGGst7kuK3Va4HG17a0+MjnLHw0TlSj8mObjqPxg0otWo9LsMWZabg+9d6aD
W0AFoQMkA8REMV5jfTV5y4Kd00Hu3+FRt+l0tqm0msKGrtRD3hbH5JnPbvjw15xx
xj/E+kZgiRqZ5J+qFmPnj66s/ZL8fYkZnyMg/I+iR/t61CdS0IA5oxv3k7VBghtA
kZ/nifcM2Nu187q1Y3zTpmorpb5J/P26+Mt02WyU/92eoRfIVY7+brruUuskQ66u
3hLXwwowmoSAsMwfugd5Uid2GNQWe3MxjWNzAl2MnvHaSdHueAAs5RRzPIDi5JYX
wgaY8b8q4cC88/6wc672eilg4qJEYKMSqIuCUdbBtAIG2nseMnRI2+RnyU/LljCU
+h8Slt/Mbjl4eeerFtW5ek1QIBA16ynmYp3aSmEWLq/+iNpSK450P6WnUHLrbG52
M2C5zLvKkCCS+xEo+kYccluparoz1PALppf1iLgSQp6RzDs1epYBygoKDe2jEkt3
sxUNTDSun3lfTiQB508xwHpnrWEJqa/+oV+y0qt8BNIaJA7Lz0lmM6c/J2fAn+ke
/iNrtdGjsewmBkU3zPw4ek+cBqyHkWB3rSc/7eXAAolT0gV6HUchaVWltgN0O5cF
RiTyMiP/pGt+BqrKMTA0SFtzHdbzWVIDVo5T7csIsURtJ7aRzmZz8oW+e+o2rWmn
jWLYjghdQ1ZLhM4qwdkO93dBo+NOv0ZakNLleij62splsOjAg4ktTxy+gFDfth7y
m4H46M9lj3mhEfLVrbTpmN0T5B1/DYuSsw7UVr2Bs4qjYdQTaXLF1/SI8oEjwzPS
ZJCYONntzYbW1w/OpV8EPqJ+xO4QvzcZfooOXeiSiI6u5w5U1sr34Hbw0SOI3A58
ALVZk/MYmk4NEXvmSt/3FMpsR0HjKJMRAeQO8fw8aOseTNhtJe+8ectyAKArr/Lv
qJ1XLK1qaRSu2+0WZNse7o/cziJjNRjxBcCdeO+Qr8r+cTlqyTRqAIeCz0S6/JRP
9g1CpIDipE1QKVzYjkdPUJ6x7P3djNHMzBTQBvlz8fq4HpvFI9N4hhp+YxAlsimV
aLyQ3b3eQGuk8URgecPmyp36c7BrUl09bvw9gNwf2NU5iYLMiLfNJo+Dv8N2wVjS
shpKdAjtQfTmdY23P8yGkXK8qqkB9qXhCuQ23cUvdWUdxmisgmzZkxz0s4tqG/IS
Oc8KnAy+DsKSmYG6Rp4rYCCslM0VGOpQryUkwyyqF5DUYHtOfDiWn872a+6Q70Lh
BG9Rm+SqTkvYnJZOttYGDnAvZl26Z0C4cZwnZsO9XuGGeUFuJNfgd+6aHOHRnD1U
2P2f2BMjChEyy4ClJis+TSUAWoe4Tm4VefQ1+7FMAM7W/pHGFVRlOZ9yQFZf5uQm
Xpq6JJQPhg/d32mCBislO9awx7MWKfRqDWJwT3qINWkXkfo9HqGuspnXTpjTq49t
kEuBKLP22JF5n1AkQmi/PedFEC2NLg5LMnzBSJUy0ga0C6Z1UK0kge2PeyhsNs/s
jmnEBXyH1oFjwA0h7Kd8G8VUznOfk8LKA0rGy8jSrSj4sSNxKh4cfS2uUTT2+qu9
JnEMVIiaI8zrpR+DBG//9vFU8yUZbEX6c7rFs2cjdIUzeeVrSPGSQweDL3BlucI9
Cu5kM54HktIstAsCrm1DXzE2/vQCCOM9yo77eBeK1/+e7BjAFwQzcXRDbaqYtiv8
I0Fm49kzAFBJNQsnDWIOuc3r7AV6/YKKeVcOPl1MtBOG8Muh65NCPETiYDNLeHNU
MY10SkgXx/JyiEr1LArWX5dcu3rMWk41zDKGuR4T+O6RaQrAKgxzc8695RCFaV+O
CPhbf6IgqWB2l9Yw6D9t0RBdm9lOix99SHy6lkoL1/uW3omr6Gc2XPZV6jLUQo42
ecO8Lvgd44ZStdjS+qGp+03RB1JC1OO5RtQpo51H/fG9mBR6mFTUL/hYB3scv6Gj
jfiikmZYSqjzN7TZYdqUKvQPKq+mfHPSq+xB2RIXtsy0gEqQevdMdmCsiQLXeawr
wVuyBYOoALVJr/RF/9i3Eq6YgDFn2fFnHma2UISEsXdGXGBxr6p/oxq8SMqAujbV
T6dBcakxTSkfLqIPyiNVVWC9IxP+KQaorHmpl/mlT0V343FAMlSzYtxMkcXKfBhP
RJ/shzrvnMexryuGoXUX03rZBWDCnkj8V/z3XKQ3Sp7pwQ9YOP/Qiq8z/BJoUh+u
xq5POtrIWxqwybsW+Qc/Ys5B4MYbBUerG16IT/bomcXwJOuUoGsPi5PDzcNp4z7X
bp5nDQkVfb2MgQQVHilURI51W+e4h30bcX0TjFCeOKX9E+9RWizavRZfjg2HiHQN
LgI3pP7i6eVdSkgm5qGyqX8mImEKBmsN2crUpUL3qf6ktZreDHj6Ms6CLAPHFl21
4xTH7sz3SwFBLDgbxFKnMsld+q0LpIFYk56B8ft1tRyQ1cbLtGvG3NqbmpdjsHBR
teGq1UeqkQlkZA2lF71fiqtkqpO7dFzjNqwJvQoG8P/EHZhBXX3Y/TG2SuBBoPth
IsvF96pF+M7x426huTFsUyts64VNdKHAhUs7LhaCrctuQO87wDyOZIYSIRrDsIij
I8oT367CSqgoiN8506HQtdott7xQOei9qDw2tthN4IXXylVcZFApB7SQLxk7sLHx
AwO6mMBV19FmnCKurioL7b3Ryxy7lhCVmDgfzNR2/g0k/aJz914VeGi3M/CqCmEj
8MecLc+22klaJ/JPsPEeJ+ZcpYTaGjbIm5YgFGFKMULzmO3mZ8U3lzm+OaWsGRzA
9GJflVlwnVQzmaT+yyAVrqjfVtDz0pbiMiSRlC73p1uV5jNJjxAUz6ChmSAtrsvC
eoUd2VDm1SQ38WLbxcwSynEDAnx6KKtKHDpmx4DVG6GwmataNl6X2pfHrh051w/i
bATHsXOixmreEQkVnYcOgFkYZCZDR23QtY+0f2k8TiyjdWSlQge6NnJBSlxKdeM8
4xWbEl/zRB60L0eyUbiR6coni4aEFCKxg+7QVMbqc3zEiNNPROJSEo++pDjg4Chu
Jct0Kmf7LlK/46Y927QQgB5mVEz3EQVWdC2GFGVxwuNVnTJx8m6IuNqGP2sJ9Ugp
qRE9gXWvL6PCXys1JxVjBKWQRyHTJ+aXyWTJ5+tJ4ExYAuoEuw7W692Ij/yI1GCc
SYCY2nqzBtTC+OS2toemn5uzRFm555p3HWmSPqDDec2Aw7RfrsPuxj5mqIZG/9HB
ee8+swiQkPZHUC627PNsri7JCC+dW1C1Nw01ceXwr355QQf8AyZfF35nWMfL3ROz
+zZvhiP6rB6OU1tuA1JVDKPCZKrOUWrk58mGwfZex9Zf0og7f5MAsdMzK0lf6HLM
vT/7H9LOirG+radrkQx8gasjfxPkIq1n+9gIufb3MqU7gQStl4mcMM6FcQRmW+XK
ZPiUCQPQhjMVVldDMZ2V4Igm1MtzRAoU/HZ4R3uQ4XsmL3Oa+Zm2210PNY2hJXXn
zTu0BrcRb2KOeUsYMm5DwIYCJkOGn56cENlIxRSg3spDNH0UEquh9GK3GH7kR0Ue
/S5hVC/QxEm5jhSsFxd2YxjIygMgkE7cx1OWjL9rFHAELTOzsEdqvkshdX570CDM
9DZyywLLGR6ElmcLHmRhAKUVxVi2Rb2gfZdtrx456P55zxDZfhwAfgJ0c/fInflp
CmHSOGFH2Uw5rAilLJHoi1DTP/qVBz07avQKEowxkXwjpQvjIpS2U/yBRIvLddzL
rQt3yOgOHl43N07hsni8y9BSa1D3kmDwGlyU9jGWGX0mfeVpbRqrh0LCDJDHZJTi
S0GWmXNCQU1fo88mJIlOzV1wCSX4QyYkv2fQJpV4pCI/vRWtPcrAXWQiE+GrHKSJ
fwJcSBi5G9HPE8NsxZboj860WgicZ2XApf4dqqwo3Z/eE/nFGi8NWCQQ2/6p8BbV
YnanV/yiD4T0hfU4JgVSW1MNPRSqXr/kpVDyBIcDmQ71ge3LAFPpdmbb2sAtRZM4
ViOwTGzDFwEPldwLHMLTyI6sKcn0UcgHsyTGO11RbuofoSjiueT4kHVLenocRgEe
QFgOGaMMUqcfrsjg2NbbtHm0SaGsCsa9X+jhy6/SolcfYeCmX0clQivR4MLVPdwz
5xDXTZkFNAVB92G0CW5Aidk3jiUUT5vQxFvopX+PnIzv4ZFE7oWuBAKe7GmbFFdA
MUv/j8yjqbQgtp6PgRzFqV6Lj4JYyv0kOl2bwtfFgrUYXxOzcycDOP5xJB9YIptu
CVMqQztJCJ2447MSOQ0ex5qKjAa0vb4QQ9F4NSOXpJGfbPKGZnpRj38o6ap21QHL
ZoWsy5tGF2RWB6+PCp+XgwXUQnE6zdX6PKid+AwVJENFdbfdEJrbftzmZGPSR08t
l5lhUvU+ebqR6Fkd7CefsVCUDyw/hGS1OOyxDkUNPS7Zhc5o0JPd+zQWqV+ZE2mI
415h2Xd62q18JD5AVoEoYW9y3uc1RiW/cVhNfpZ1kMxr5RFjk99ZQPiJC0KZlSnT
8wf8GSg47wDhkCJasu9Ceb1z8KssfqLbnvW6Bqqbl/U8GBb3E7Oj3qI4kJKt7VaD
biPcefJDWxNTekZZ93N0v2X9717QmYY4/l1JB2BegFsPcNRe6BZuE6Xini64mHRs
k8nSkznG9mrWOl3IFdXOKClm2waCqIrttiNeE9p0R4zoZb1HgSzCeuVokbaFNZwx
BFmt4w5ptSrZlGyhc+oz7804acFNApnWBEffTT6N65QLxT5lqDWET09LVI+yX4q3
9qox4SY9B1JJOfvFgVZNeVVu5L+Vn+tTrXAjWnCT45EVAsZKJoZlWTZsGcNEdI/4
YsNevtRZLjXsaniQ+hkxB2QWInZ2tTRsuk1FKGl+nNUUrITEjj/Zqz1qp4o/3Ouf
7mYEYgOkqIdo16BARVYRPaqE9YKxpHJ4TiTQjFUWrzCtW+hzrObz2u97WFmetjy4
iwchn1+udxEonqZQNc8mlRW+45mIQ+NqjizBKZU//nT3Pv/V0+XaD95gAHGMCjGj
zGk1sduiD2yxB+LaP/wfuZu1Lu6ILxA1ub4sHwSe4F+kfLg4hGrQeckE2ks/u2CQ
Z1yVD+dYVDjJw9R/pE3u7YyIkZKEJK4LQNVRRoQP/sjt7ksVnG2vcvAtjCzsQxtL
pVWjisYJ8JNesdDq9dku6HOsA4d8IGsp70EeS+teBAHiLx6iekwLVuXE5CqhgY6k
2kOi0bKudLHoxDO4OxVVzqJ6SPy/GRRGuUOMuKbdR3GSCyq/EAQ4Mhp8YGIVaO1I
CIyOO1NqG6krOFT/RMlHCx0UrChEXhS55+i+ZBwAqbKkUvJ8S0oWua71Ke+j6vm3
zNVNO1kv25ih5HarOa1oTjans/wphKWEh9ueiQ5ViW6u0zeMcpbdmvuXV5MbIHuL
Zla/ZBHaBo7KiqrmIL9DJz/qCmzUqUM+2BhxYYtHUmCz/ZctlE0odWAXQeqaBTh2
Hd3387zdZuDUGuFddd6blqy819BTzxXLCXWxTcQMUD+FPDU3smYddgEqiGUTbAPZ
fRgTx5rrshIVGqEZ7ZLsqfCc/5sneok53omVR8HyAQEVAnjMqINMnLs46u1Cz/iB
CSGBZf3Kh08Ir5lkq4i11GouCNuh1nby2fbiNKaJqa8VTNq5+gmme8vGNyVi53h+
xWPh827/wHdAfkVxeH9cDRrvZd0QZ3TaFG5/WJi52HT7f7VcWS8jZWkZs6JW14Yf
eC1cyUWX2YoUfeK5vuEaM7PjxTm4v8nhnigboN4p6vq27IZ7PxjdcQwf64YmOzry
n70JMEW5Vt4OcHF9teovNWFuNp29PPAEm96/2BLLvejFAKMj9bs7amx5rsKQTMrW
pZeAvFm/lPXxCFwnnuyFrjlOmzeRg7iTmEhO1SbvAAiUpCfvtwsLkQtexRQXdjRb
ZTptwnCeERGofaTsg7wiuyno9w39VMWwTbkQCKIuPDQCQhbiLHrv7P0qC5uMI+jf
8KlLm17BbiRPBy523/kkvJV/is8FLY5QNikAKvCCGO27XFUsq5IL8/hVspIvlRNL
kZfwPSdfXBINjE2yW21TH4GROqVFid0W+/8b6U3ioKR+hBKgieGA6oFEQnoXcJhJ
qz5KHqFPTI0gunFjtFaoyiPFWryhxcsT/7DOLt9jSkj6L48nlnjBSqrP1eusWH0O
tYVJvd785LguYdRjwhyqVqs+5blnQniLnlT7G6bodRyBu3oPlCJ1Ek5aTXzYytjo
fO0WZVAnnIlFSv3bphdE36ecqIFm3K2VoWJJnsQOSTBjedHTnHq3DH8gOhAuMMLk
bsxFxk1ownTHxH7gJsAz6wanGIGSOQpEcnQhOvIkFC624GVpmqouBRaee+pZb2zz
X4lGt4f0HYIaNOj2qkHWkMutdqq7dg9HYv5y794eJ/+YMWrbbvxgL4hh9LeHTED0
t2dsrpjgxwuMZm62TNq+OSefa/U2HfCeoHlW/dUw1+InrycFtCKXnQ3c6CuQJf/H
oK8+k8omL/os/ZFgFR5+veThPTevHqDvw+/BOGq5NtyeKwRXgWjp0A3D8ClCGCSS
+7K5CBYnVSytWu1wS9G0gRPRIIeBKkhiZe1i699F2hbn0J+zarTlTvwEP8PoZdrA
JUy00zLrz0tYZOkpgQfozudN1HTU6CcdUFtnhvGs+WzQ19kRsRvWkHNIbN9MYxVe
s1y1I7Txr6lqJrWocH48LkLAaIAwhUlg861gX/a70BHyUEYqFNhaof5zvcBidraT
IgtM+59YI3x7GjSHOjIWA2nX6IHfL/jk+aASyhvFBYnstmty3u2BQZrn7NR8KVt9
KZ3syQfNqdjnFzvVjiQCeYgVci5mGWAwBDbITvRhU4xgak2JfN/mranVYHeBISya
NOtE/F+WSs7Srs0YrDDCSEI0mIbGuzIbUzXmikBa4Pqab5YW1LDWYGYfch7FYvcC
fkiSYzfVucb5s2nGsOjcp2lwj11Mu/bXjq/ssVdq/MKQ61x0/yFglxd51FVTBruc
lFlWTYSpbNTmQLL7uLdtkAsIe0noXSUBxINQML1IhtmcwZtMXb+HkOOGMDi0Z9mv
oy/odch87xNq3/E5IRFgcKPMHcPRdPgF71Rt2Vpfk004OKk+3WwcrIIE46v8scXZ
CRtpnu++dCYRRCRDbFTOIsrkCfdgiLIywLcfmLD95g5IP+fek22DDHPT1PdHwJLO
+Rv77d0CeeNVDN06bFmVZ85ibIE2wtbEJ1P2kRNRPUP5tCY34q7rGCbBAv9NxZmj
KFHbaHIBEO+E2E5Jw+tyNII8IUvBqHaBEt6vx2TJmHa3qgug7yOk1uyFGc02z7uN
DZmcKXGAJ9oGgUFp1U1yXXxW+PzPBnfeV5qJV/nOpMHEsBUFGatzjN4PvafaYXo/
EgNb38HAdjNlp1J4m8HgCyVBdBuoK16D62GxSLOUF6w3nDyazPRPafWOC09IueWL
qHbsHpHtFwgUBebpee/D8LndVU8tyyT6Rq+pucOB0B50TbtXOYOC4b0iWCKDRS27
ptFJyuXkcGKdj+/m4qYI/0shFAMYO2SVfkkTPviGX8pXSBsbDHvzZXL7i3bWHdLz
lKKl0DCbJ7zpbN14X9t5Ff3viVTk69gdDYUtYWE/UI/vMkZmkPKCKktVJ4KvzeJ8
xQMT7H9mXrqQtIh+x1ItdwS9eKDIJWzg6hlyUD6C30RpvzbXQiW8Q/kcveaoF14o
s2Zd+tRBHEiVs1Oqn4hw0TaMx05Yov/gy/gVfnR2q7Lwm/AcIO6QzTCOP8RFRv+B
y6Phsb+tcKEPjMhC5cVyzEW3+FAqxWbNQXkFL7TOks6W8Fat2r5vWZRQjtP99kd/
Vo/eRakSgcIVfR5sbPYpDgX//Fail4l11xda0mLeYtwz2cisxIftCbnJ6ZLlf08J
vMpcpkOisrnKBF6+T1HTnRCZvF77PHeZl2OUzrq3znTyGftdZsjbvaK6yVxa9Z2J
1HihUXXTNcA6BkXakZKgRnkPobFib+/akZGP3GqaZ3iDNmsZn+7U8qV6FNBG/k37
W7e6ai7ASMr3rzwvmOFnOWN/aHtQSdfq487o+BamI9jB6N+/ve4IYtDa2ytUbxAq
zLCczT+POxWZPgILOiIwAAtn7a1kKM1GFnmqmv2sh1S68D6BknJMGtN1Gmp+PhQm
9HtTLHoXiRG8Ooz5uNY57YkrRWS25AA5auh3Dq91F6UJkwe76tGnp/DEbf72qMt2
+v+MD2nEzp7xbJNuRhDNqvjwURf3w7XCLDVnBwdYWn7U9XMEX1lrd8ftjBNZOtc5
QI9BbLCdL7HNHOcH5PkmnTpW+HWKvZH7ijUdXoCxrBD163MvA76UdF0NLiSgv0MY
WyDtF6kbpQWRPWoCVXX0idzDIp4Rol5+1TtTmXIVnbDWJgUBxOBP2cV9dJLbcZzD
1Qw3oTz7khbhMjgms0eWVLOrZbId6FIWsmQsVqbj+q64pJ0ntoCQ2TZl2hGRgoJr
dPZ3R1qEQm1SzzMSh5UZzS4LN8Om12xSXDLxr0/Bn4aqFfZ5verdWYtMvdG1OApC
/566bRsqi0vWINWmiRvB9qPA6/XcHEaYyyE3AhMHqtnzkY3JMK6ahCXOOqCU0Ke5
iXwjQVn9qfI9fe7VGXFd34kpkf4NnTmVEGzdHTHb/7PLgrKkO4tC7Cf5cflefALD
3eu+L0kksAMcTvr0BA15uFn+ZJ46XmtKwWBwIYwKsM+Gx1juvGiljM3FEjTTvlh9
sIYohdzpy98z9V8h1qkp8lY6o0TOk6FO2XHyIfHomq3I2cZyqgh+OR4MIKMERaNv
LPozj0EX3yQlBMKqed2UgXMLWnmAFE2i5g4YFXYUKd3QYL7STra0SmG/1WAP61cc
YTQuYB2HJqdv07pWubL6KBvbTfZstTWxkK+evwQldn29oTvyTafG4bfrm5bf9rSD
Jd1eYsj1Fkb2zhKFfcEIZSnPwXJMunIu21STqnkYYJQm2WXGCku+MZuHxRthOKaT
W//6zNk/nEAC8ZFuEtc2O+QRvIWfnl4m3wXPJ08yepy8XXO+8lZTCnRjSZ6j5Oc+
+/K6efLf+vsRAfk4o9ihVPijhH2xdeLzPBtso9+VzvJkhOnlMbv7JsntmGQoSvTh
bdsEKKaOuXmz3r3x2jfQ9Mpie+VtaclI7OBQqOXBG5wSzrcgFKqqr0HBkbAZYKk3
cXuRngN1nrMYENbNsIUKDeywnHT0rseQUqH/RKea4k3fy7pvDjK6PvswmQI6y5Oa
bD3g00FqLuCiA9QKT8murDx3e09cpOCBx6xi+juC1srsvCFrWS2EgDb8FMe4J3e0
vlJkWE7nhMrJBy5CilKZPEjTfFUBBKKwj1p6r3DWpgO4ULW9nLje/Lyz6xkWH2zx
gIDvC252WUQCRgfMSyC/XHIdb/9Jjc2x3Lu4ZoxlnoxC9j0S19aqLqzKEseZuJYj
Ax9qQpmHa8IuoSXmAhWa8EpCgb0yneybpxMw/1cWVamGDv0osWWLAOn1OOt7TV/R
FHYUoEKi5m4Fg08XaA+n2XSlQB1SXlui8KVcrO05amptLv3tRKNneFzI0lNuX1T8
rK+6Yh8cG3j7pFBHQBECssleV/hTo3KBerhoM1KmO0b7wtXJpBxKBxIlhpAEgoS6
GRTV0y+wdJ+3DMaKYK3Cs5LBtDk2CMjCR7zqTZqt/fWMo6uuwdUMi3fh2kkYTsL9
2311APZxeoFV5iTR0Z5zIXHA7YeudMlBiG9lLBsq4Ty97g8/1D2oBEgXwTewQ0iB
vNDjiKOjGCSmMhBQJWqlZZqmWEVpCOIMJFnlbF2SujZxAPPy21xB3Thowap4y9xW
0asH2tHNHZ6Acxe4AVM/8eievJqiEHhUGdSzKqN6V6Xfnjr/6ntNjtIb5KShlH22
kPH4MdnFKExFjY/FlLvV4C+ib/v+O10QJuxI4mvSfAfMghMP+Iujsva9AeP711x6
+4QFyrOJQfMTsJCmRcEGKdfYKTbOJ2ZTdVRHxHDAY1gi+xXQ/chlQK6by1Yj9q/L
K28R78v0eQVj6T93nfVU+olGpFIuLoweAdbV2OtPKVz40jlHaStXT799IaGqA8bo
uEyYQpCOqqSkrEjfcbsHwm0ijRNMcnST+sBGg46W56PavkwIYMXcD7u1Q2Q4uRll
K3qzaqqnc/NHuzCnwo29itQF36X48PM88yLrfY1MRzdq+i/KAAvTLnTPs+5co8a6
V92bTbdP81xRarEnWsFTsweya6O0kiIlHXOhJktNLt3HmxA8OlvpNqjiJmUP8zsD
qBk+Qa9nFz2lOlHw/piIkGiTAU9ftPyg1klSQIJYZkY2KAkORWI1bRwvalyrzuJO
xyFAdhu73qx1nuGx5g2wtid9US0JnIeOIfk48HqzQE4839H0Bo7HrcWxy8wmkr1R
ukvIeUWa60udPa0K9Wp79xY9y0kNyHv40Jmfk13AFw+4D0mvi4o3xS1S68NdmOXn
XeehgsgOeb6wK+ewu1SmDYF5Cphclo5qEsmvgHyNuIqDNbdCA/uj9ROqSrJBtyMj
xp9JXepi2uPUa2q9057rRHUPHv3FCBlzq741PpjIBENMkfHwkFb+dQ8FlohHTRxZ
oULauykXo0hPNwhKhwVUDCLuQomuOI+r3Am9MZaqR6zxS4qxaib3bVbmri5MXssH
9zK7GBsKxoscY5GgnavLZV7ZyriHSltG9tdpWxAsPB6VgTohVqs/CfVwe9qmatL6
VRO2WkN9HIip9p5ZWuzw0xMsm3vXFLBdP7oeAYmpi6ocWV+u+NWIMafS0FHAxuYz
WKmrdqHuh+4XT3w0/y4SQrMu8ZBW4ol6UgOqY+ngxo9P2wRLlwTB8kNyHh58Hr11
twgSmodgK7U/jOgeNX6W6QdnzsBxzjowQKc84PvamY3g0ZJlrCP8mZfDxi70M9bp
nOY5bTf3oYR/WXZZOs53eSHKq4MCzBhL17JRlxkj2oeGsHUlR77ECF8KO0kL6C4Q
Ze1peFBJEg2vTeyuihGzmmfTcdiHaf3txjm9DJQW6at1qiQXd2kTKvAjN+kKxquJ
Yn94Mu693HvlivrtgwPQP0iL1z5v5qSwlplIjXL748Hv61A0dBC3ivapgBC4nVTG
WgMmlnFBLcAiHJu8kvqMLfDEZ0Hjnk5tt6MngXUuHGEokSvaC2cF8bN1eEpod8Pm
DYpOzjxhTw9zoXSlOWi1bVaNcv5Z9aQBQ8C+f3pknLfH/5U9Kh5yHxb7VCPB1Mvw
5UNMoVuMNxY50O/5GeoRqDnQPDzuV0rcel9zh5J+uT7HYhYQPgVgRVDtICzUPKLN
g0OUNrFQX5UTCMKIFxZmZHtP7FdexBorR6q/NvtIuj6WyiVjP2QcDrV/RnBmCnwj
WsiOtzJsa235Kx1GxGmcwczl55e0syrJzGyxAZ9/6HM6kOjHgg0n58+DzS2EjAO+
OQyyUc0Ofpkj5oxKj4Qj9ZHd7z1rS8FNYJpLG4JGK8XfCUhkhoCwI4H9ae4SpqM+
uwQjhtXNe9+cEpB9YxsiD24wFHaGce6IsoRUbaYGfyODzDhLnWVzfuYKJGCA1LVy
eDy1oSH/W8bOKiGO2fIFTN6+jAcfcbxIW9vc5XX8z64pxVh0ISDn75yQ2twEdZEU
CNi+sY91ThYdoJz7MU8t5BuP9TAxsEwxgJoFA15Onqhubi2/ZSmZX9b/5ffX3p+U
LoEqzzpuOVtLkWkMoTtk1I9YKnW4NPSg9VQPljUuvBGUgp38O9Xyh96XcdMsDcQ0
NDkcRWVHKMnCOvWBVMLJSjmhrxJZM4CcPNUYvgd5zNfd/hsbra+JjURepSgqUDQj
9szbI4v3Wc3NDM2L7vgpo5FQ0Ud4tIca+rI0wZc/oPCs8Yu3y+8XFzK/Mweuvkja
/BrfIZoxfgn4I3pF5IJnFDwVHZ/cskGVazV/qZ7NzAYomaxvxdPT7Uz6/DhI+r53
sLM3Oo4WN2b+7oPW4/8/6qVKaFipAhdOcZvQ3sOimPZov3xarTcwMdpyhraGyWD+
QH+Rz43BVJsoOQKMYLScVFcjdVbVXTjoiHc5+wUIKGgPErd1t5k9eOGe6rCXYA/P
msEqtxfAsuN2uvTD+iJZxy63JbEhTS7YubWImP2XeoSpiTfHJ+3XqLiXEHGucmC5
miKRETAS4qn/U55DyN9u76TmGfjGPCcVIF3wwC49UoneOcGVL88Q0PGASLWeyTDS
lSlafwGeG5hZur2vaoSc3foJgPxcvQvwaJvb8pV2C9OQOuXUVQJZxkZK25b4jMim
paLgfhsaFXmqtbONmdGeH0rqIPnWdSnMp7rDOsYlfucfxo48Ge1DT4aKLiSr3pHF
D48zl3Zs1kTd4Tzm5U762mP91lVX56ufM/jaw3LAt94CoKEVDJuTTHe3gpLJYHIr
tBqvcbM5E4BVhcRvpvA/XInb12R2zuBHj1NV4ohT0jQCRFreoCtDSLunOOVbpkJ2
wVL2Rg+az8QVjyGPu75Sy8mwQoQM7MNS56h/amJ1L0H5+mrmP9N0ox3uvq1/eVU1
KPjA4/j4g4aDkRPP/clnoN3kL6JPLu7OL3/3AcBlDsBC1muYmwV+OjxvhUPWVFj8
8MGrfUVqq+9IpWdGjJmC11ywFp2B5gD4yfmEZKpxTxHNEG0lPhYszPEWtf+RrCs/
jsHOOPzLEPUfSYjfL4TW/9p2QohiMM+MpJbB7Y8gFSOCbCu6U/Nhn8+4fwtmCUgh
VCLe+D0/AdV9HxEVUoky8mCnYKBnOKfkRGyDAkfHqN7hbXAwI5xZ5iPqrp6tZgIP
Ls2CDUp7hH55QDWZIfeNSk2tlmQ5Jjg3x3jmLDbGXxoDj8BPTU9+hJs6kFthn237
omnXj5nfECTOM5L/O65Ock0NibArulZ6KeEre1Bjf0tEgCr1gm73mh8Z2vINW85r
S2kNgqvNJPp8D0E+az7ISpn1Y35t2mJCur0aZwbO9f9O1G/H5EyI3Uxqd1Z+B5L3
X+cHHhcWW48fXfG3S0Dl3dVXJFXiawNkwsa4g3hRot74xHsNDITGowA5L61fcLcA
5/fDs76LqDHIuwSZ6kt8s/arYFrpbykBK5lKKzAoxNtEizlQQWHwnTIyJM3eQYy9
lIQ+vr46zh9hwQZAdhGRA53ydpx6RKB5lylcQiDm5Dafh6q781CTCf/VtiLTxLiG
0kBGzCIGXN5K2wXzUmK0cCMjXtoCVeWqG0YnYKbKL4sQqnlvV8Hqr48siIMy7AJM
/CsNBTlbRo7QxvFFYcQiHI0HeYZAj4t/EibwKMzYTJbZ8WlAuuyNJI2oaAlnCw8E
8QuNQVcvory8SIr8O4nUy8u/hgpJVBXYrSsmH2Jo2Sh6kA6Vhgaf21ihaepdcrA1
jaCfcT/ziwTPzVn3ZXzOCmFBaDCUk26DK8mCk8HWCbIjllzEEcN7mEawp5yf/YBE
+LW6CHH/djPmDPVM1lrIqhx98+I6ucp29Qy54ukEuS8fajq4E4F7/rtUuhKjAwF4
r20cg73PKvl2l3F30mji7VVP0+UeAIyaYrnIf8QdFYoE2wnGexNuL5tl24sQwLdi
fpuEt3uRKJ4mOc7einAWicwSJwSjIjVe8HnXKPMY+5U4VetoIQUs3mcIVav6G8W8
v/TKCRB3clYIkvTR6gZFg/42yGy+52rrvKxbio+LBVcmmZM7ZX119d9gWkmb75wI
J3uZ2Xy9Q7xoo87lA/wISmVH9aSK0aX+yPSMuPdxj9b0sOuSMmTtjXxb/4T1ogtJ
TXGDkr6EYeLnvvTk0QaMf7EeZJv8bZiifrnz2aAr45BbS4hi5NVd4XXdKhiYSjL4
cJipUeruaQjr3+gxojH4FmiVvJVHH1tIRZb2sQgepkc6tss2Pq5fd8+d08jwRobN
+igc929TdnpvKxX0yJuQ9v0KJGHUnOeUQlGoKe6354YQ1aAsAfZ58cnP49gzDJbp
XWQ30R2AcUwP7zX+mSXpwwOx8bSMwc/Bcfon1jS+BBQXcvFHGjL2pReizrBZq5WE
SLFbeDl933qFJPffvH91F/lH1A7E4IFPk3dce6/7grqA5PaACV8aXRIUi4KBubgx
sJy/NKN1Ic/DUmYkPqqcU8JXMpInBljlesU6C6b1NPR5pSjKmi/SLJ7BVpFIqWSG
C50azsgLAz69QwnsQjzTsvE6H6p9B7NNubTKbTGAoosyN1dYkg8NVYNbrAu+AZOI
L5VTVJFK0uiDMl/YHeyTW+maabWLD5XgbaedFjInMdg5Djg3RCNOsVcz4V5zllMU
39ZdUTWXCz3F+2dRTUFw+rlh6yUA30H5wSt3ChKF8uUtjXrl+ntnGIbFJY+vNXbY
pJ7f9clPmqvdF3nLt4toUMfTMMrsed8UD/BGIPbM9c3Hx6Vuw+3SiiOlJpCXYTWi
zcITmySP/IEb2YX+Cuu+UZ/pNKUPLQLsyxjmYHp4OwQ5dB7ZEf1pN8Jqdw8MVVPD
0kKde2q0i6uKt12yZVAglrWT1Q2OvAvsHaprcDKkbd9Cf/etBb8on3mX+A8ZI/Hw
aB9rJR5cnFQjV9IZKKMmrG/Zz+wepc6bJMeLff1LyjnTGsbvzyS0NFW+ZTl2u38K
G4WpotThiFFisd4GEo1Nov9ombmV+fg9wgjVvikApTVE8W2TFrLhDZxOXUG+BOjW
stC0OJi/af+Uxa7rXYETUFZYnU1meqW9Ff71IBz+l/larz1oFcBEnaHQKpi/MYcF
HTBVoy+kJS7aGItWgVpfgSYqkTQE5O8r0p64mDBzt3gf5+DSDqbdYvXsqDjiAkCQ
VQzAduFPhjzyLqea+DlPeRnTWXqSv0E0ioRqQHOSdHAqeg0VDtLi+I4KusE2VBit
bRPqLZpjZkXu9qkk+sAXsDgcrXsK/gliMC7W3RtooATRQhzZOwkH0Qpuasb0zZ14
4CS+uZ8DO9+PlqjXodIM2pLC2Qdbkir9bmiTKmVXhF0Jx9p7xmYVCzLLz7LzFUsT
Jx8/OZIuFpsuZEzD+rvWC8qqeeniu0gAcedEdgvhCJYnhDhvz42UYFiCG8X4V0M2
Pbc6PA5FA68KPSUvG/qCs5xtfGNazpaNohTOobMuXTebjJibR6EaL50OymoZ8cXs
KUPDBf7oztItj6YBMDRk0dVl/xqFZkOs4+gVJKmHkO3kLQylAmzLOky02S2UB8DM
mTEi0JJ5PPAYvNrCvy/U3WTR6jnYT22ulEuH0lwhVUtdlG1NA0tQjd4sAqUl4VSB
4neW+jVMnnEvL9iWg4bsNUuoS2yT5jyCaLbcdOOCD9q3t6fgKJhtyFjwMNUxUyhx
BC/b5COjsu+XSL+TMOwi6Nfh30KfpZ+1p8DXzt1UDbjGsLCRmoh7zkR5iPPUR3r0
pkOEwJKKqKz/uxrVbmpQTBeViyVeX9rNANLiDa2ntdBkG2ta+leB84WYoS6L8rCJ
v8kbR14Su+VHhS5n+NEhThijaqeUr+mnANQTEgX9BJP6x67q6AXApGEP7V9YJU0O
d4JVB2pEaaiO3OGCfwggLYfn6RO9VVLQYZj0GrJAwCfvAfX4YP2yq9xd4YIToyuJ
Khuo2qvKV7TKRxcbr6UFxigzIPcpEJzXujaxR4USeXkCAcN4/8FSqyqkvxWlJYh/
1RkZ1vPka+/COaJpZ+tmYgNtEE7tJs/6yrapbdTpRma2KBDw9i6Nxq0bNW7EXQWh
kMzvinaSRi/3hSyJOkUxBuDgfZNjY4+c5RODPn8xNWDiRNtjYlS6S3ZhlG/itzef
N+I7bOkVQxd4CQMRnG3uAgiafZcLXoGrzahjSJK/kREIjx6Ngn03wGzEvL3GtkjR
CczTKFVa7theJH0hbnekO7CSolxuKkkdNcfa1/6GdFX7C+mHiJ4DDhoik8qSjZFA
EaokS0WA1c8ULbt7+rDheOS32cLahlNoaQCyPOi22OmyWctQGiMbyTdWo0REXj40
2pFN7NkSGW8/e+uHt+OT1rO6nOda2MW4vvBAY0dxDpsbc9b0jgLAfdOBUFeFlYpz
63QKqNbCsA+SsL7/B6SkN+Cq2NCn+OT6HmXgVMNZRsWgCibzq0tvHCcKN++VDNgi
1jBHQ36OC5loxZtm8/XjLkNN+WaftOAiz1VxaxccqeJcs0/HU4fKTSmmq8hcJDYj
1oxyOc1KqMsIYE/ydM+SiAJO+HadmPW9gcvTKVfGU0CgO2s2igqbEH0ROaUuB5Kp
RU7AQtNGD2N4Dkd0YbVSdn90OYOGTq7LWFjTvVF2FHsRfFqu8l4Mnqsv6D1MtpWT
Do8YjiQhZ2fXlPFjinqHVC63yFwMHnMHwnB9IhaNTHcq7PhaHQ5HW5vBzSssdQgP
xIygs9gMgU4HrniDu5v8LuYpLwU/pGvFoQXtw6v1h36UFrOM/ix+1XnCNpxPOTnw
8lIii/zdAZYPZ13eSjUeUeFs9uHTeNL6BBrw8AHgDBmeK6wPZKYJC5HOfnHavHj5
brcUaMDV8ZuFsjbZ9PsramGmsxSIB2BKCitaW//CncaB8AL/jRTj2fr/ozi3CsZk
hgxQDzUx6sZtGEJWQ0yMXbaJvCl1XQ67uT+qre3RkzojlFTEir/jahl7XQwZSpcN
YNJ6mWH6NLEWmSZ7icZCqCC1VZhWorE9LIoiPCLV+830I+1CZn2VmAGJ50ixlYSm
nrldWnDatG1jYE+rO3IvoKtTWEemuVfXVtyU7FaYb0rGwXyc/9s9EGtSkEWacYSu
Wv2yEJ1SJr6yIxvW7vYdLzHCPSz1iEbDiCrC763eKAHfFdIMAP7L9s/+taGQedBs
6YFqOnMNi09FkY1vLavu1JTpCBN7sjJibeDwSSujI8s8X3vjI+dGUhdZLfwTG9M/
R39HgMuS3VtV6LEgpp9b7vQTBSQI87iu/VG6sKawG86l9JJ2I2jdFvuwZikL0wWm
qSLdoRPCMv/JjP3/IoqD7CN+7ZGqQ7UrLF0VUCbnweCVMrIwMKK5TJjzJwcXUnLA
K5/kNPYml3SVahL4D/Md8CYWNsFoFygge+siQ4V42gPT9i5Z9g/M6UoaGVCp6f7N
DEZ7O+EMelEavwgDL08IC3yMEc/p0a5OsngL+SYgu9SKiFAVLQuaE3iOOik552wl
csdGP3DVraiXMwYepjdZo1CxheBH0TqDQnn03Ub4NyJA6EmGRkv89QBA09oqX5Nf
fXupQn2jQrJ827AJRFgmeBwCXn1Fq456teYgpsPjb1uKekw+6XrYrxBFrNxgS/RL
bVajzzMEHYMV4cKisr3YfwM4EZ59vnvWpzb1KBlvkfP8QKnkslfrpdxUzLdreAHy
mGI+RaDlFs5B+x4m8lwQyxBOXShMFKgr3+2dQwTjpF0YOE06WTtcxhvoDS30adwG
0cvo7WVD1j3ZlDcv6gxJltGQBbQRvBxSR6+wfWtKyj/rtChq0pzL39/HdJ2ogwHP
rZ6PhAvUYnjTLziMJrw10Ynpn/CEbvsotRuVubkMVT8+xZ5kEjrLsxYISUfCtrfL
hIqXz/Drg8uv679nOmqSuxI8fVoWAcDkV3YYqrVEMmCwp5Yek8RdWCgslG2T3gk+
GpupD1lqJi1GjqBbueuL5uuZB0tFnJCbOeo4UUOmV89SI4Oj/Zi7NPzl9/n5yq4O
gpqqu61+IpvgqO6a9jjK82YfJCqwAtzPOsfxDTZ799IScdzLP4F2H0XFSXszXIr+
2F7qG9fpyolIpsFWGiFC2ubNAcSs6PPL7Skg2oun0iAB+cqThzT/4pYSm5kQqaxL
WGpvdIdsGc9dfePa7wVDIVmEy8Tv7sxJjishA5p+UeHd+9xhQOdY+Qn1zZbmZolr
nSOfFFiy/0JB1KOrUOK5dC1fDKfoYj3+nSuE/PBZ7KBjOiehIs4WkO3dCjAdiOvN
VjyccPVNRphfPbMeadg1ELe0n0HpHvg8pF5+KaLjhygL5KQVhZob/XVh/CiIfG7e
4D1XADeasdTL2ULWDwYhBoLkxhVpMjJIptU+5LapaF59kZQa3jlGyuoWHAs2Ttuu
+ry244O9zcFcuk4oMaxJhtJjVyWwB4Njd/oca9ldRdXcgcF1tuThfLABjVLa1E5A
YfglOmRNBgRO0r7YjEortzOrW0hN8iVZiahKdiz9Z+xovLK6ww+UNSQW7DrRKhyi
JLbPSGDl8+d5ubruYbP9P+I4UlxHSks2HTfoD2AnzhaK+9FhYayS/tCrarxZ2WM/
OSwRQeH1dCql1KvBwNJzGKYA4FplfSjO2T2zSxMEbSKHvRmebo2wloA0bInweVmG
wkqfOduezca8U3mh0cSl7djjCZasLLFy5zDiuJ/8TgCTwN+Oe4eAUAzfTjGp0/NM
OqaaPTVW0KfNNPwXaM4hkW1PQ/iqef0bM0ToAetX6XSc+/LZy9isEZ0GQKpbGxKj
qjL6JlfnPp3O0HZrfMh6hCOFrRzCcUygmNzbSz3yzgBTiXfHAhbsuDvl5P+gNqjk
e9lLc1ku+NS9Wk3Y6zdWwXmBL4LfO4astWvimtsY0f0QyV/Kdio83A1+QIqHlhFC
QuQCgXk7XxFHJL/29APalPsSzMVf/15IkmyGLCQfuXBfBz5C86R9IO7C6l4VdvLW
eS610ADEhtQagTDr4IUkLtabjU+ihxiMH3M+i9dT6+gPmFYztVKyRD5IvtJ3B86J
er5epolbi/hp0IvXeROzoNR2GefYdnGiW5XG8lvV0mKAkXtJE55RnOqyUtnAhQSR
Sz3DTsQnigv6cY3QSPRLCEerBx0TyHoBFppIBxeHb6Bs5c1jBCV8N1Ja8s/Tj+5g
b0Q4JhAuSPjvyh8TVqEpXMe3+J/+dJ1kQSXEmtci6xi7LsDAOCYWDZpw+ikNd8Mg
DFCwNjZoxDMFvup7WjEWewrOT4/Zbg2L1iwbDaXNm7v8/Ulx+nd73ys9PTLoKxBb
FGfdn6t8ipALeEq8w9gPAY5Sa4G9k7whEbrWpFkUsdd6bt3iQMWLKmv9kBZQxIL7
iD1plxjIz4xcfOmVde4uALHuYadtHFV4DfFqeFTC0JOMphLQ+X/TZchYHKH86I7o
X80C5MpcbzLWHuaoDgcIrCIVhYcMUpMfJkfsGa+dfT1iEy9c6gHtvSORekLbsJML
Osku89EyYF507QZl2Zxk94seRNptn8AqJ7ZNk3nQAFu9V15HkPhJiWwz+xt9BZLm
jSDZY+9GtEg+YrnoFsPr8GZ1vea9B/sap0ehObUKGkMpv84PX655gD0+h0uHdYTn
I0sCTkutsRHyK4ld/WlNTPOSHXNrJvKf1w1qWiLx+e6fWSXcUt9JKlctF852eoQo
JcqLCeKA1/W7Up2/+ryqstoDHw2eadLFoCZeRJTnDeJVPxmHyzvY9U+b1EaGpMor
DznxlJSa+DuA+Y5kpBzGJkUaXjznHMFJX50K6SIEh05AZwtwNG6jgWbE3lTkjN5Q
ypapK01JH8yOD/HQqaGc6MZXmliUZ3HhbJ6toIZv5AwFZADVsg0xUJrQNqL4B2j1
5EcakNbmL1xM+1s9q6N9NPd3B3MTti51U6aCiyets81V9fxg1GD9CyQBHgn7/ibK
hix/lvcgKHNwPZn/xb9p/FnaPwRrcDqRA01mTtw3ILrHNjbC2nybFsrRlYFaCZIl
qxoZU2++/L3YxoV/BEEGcPHaWdPN7OcgjAvjj2uu5ypfqJ1Eo5lUrp+d8F1Vmm+c
8j16aAlR+XsiD4Ca7mcK0WU0Lysw6zJWMTkODDCdsRRApJFHInozCMiYcqCUr9um
xiMk4BLcpewcpSnmzJsv6rz2pOVcjKNl4p/OmzkHrzh21ameoeKI1XivvSkTZqCr
E4rafuzVstZ90+PeiI7xyHYj2lHVPMth3Hk+G8/towJ+gR4wE08UzlMgDZuyDlOR
j/IL8hyoIqiBYAukB+UEjlFeA5Vgp7oSJH5G0CudlUB+LWK4zq/Vzx8kFkgwzECt
OLXRWPdzqIto5ks6l9aRPpcdjOVCxMqPnW89124ESgh43LhXPEiNKpR6l6Ir95TY
gGdR+hazID98A5OEwEYnbw50t2PvaR3asg7ky8Mlk3iAlz98O8ifTXmAMuwg0Yd2
6mFoQd+a3NolNvHewMZjE9QWKY5f+d17hQB6j58tLMBu4aX9Emrv8TbdXyYqdARS
jaoq8GiC0U51EKgvvifZti7Tg0DMz5VjCW+/ACQj9DKkqqxNGR4n4N/BeQQdN0GD
U6m0pTvEFy/f2fXn0exxMwfLB7MmQxM7+2MJzC0qaHpqS5/ed4lMPYyEMI5JjEaX
0oVj1sx1U+EjAh63TnsHz/IoBM0D14YtxxhG4P3q5PzCujFn3hkXTSYfcLydq5uR
9syPrh//xWIJXN3pN0IBQib+1yXxcig4Q5brrieHXNFlC0LiAKkSjK07cBcfuoc8
V5Mlqnu27iXWMB+XtiyBy4KCDHGPSkWuVf2ewMJLT73aQjntso7Bx6pGvvX83QCe
gKo9E9SoJBj5zXUik9CRFNtPorcf6+r5JfP4v/xrAxjAtCPKYW9JmeY1dN5/0AOG
ARL8gaRcS97zoOujql7m++Dv+Ad4jcHAk9NVA1qAjURTt85GtvFr2c65Negra3yc
3w0GUFsaSKfw1uKa280BxUMvIxpwy7a1YNrMG9Au+YkU4uULzhqpWsxCpPBO9AEa
EPQ6PZzhMP4cI9qLgHHWmJVlKoWjCyO6kTMmToChJCEeouNUPcWYYIwRzr+ICTOS
XJ8KjTRA13OdynC0/1FPsowIOEQyB9HK9xjXVbkMvH3jI8S+uAkHbP8a+u8/PT2E
xSZFihmHtkv7rfmdh7BnPfKNlsOtE3YifXQcCnAd2NSPhGDo9hYvqrCBdCs41IuR
4sTAB9hwCcexCEothOzTRbjkb7W1pX0r7blUtSXKdopw0CPw2O1UGLYlTfwm0rF2
ury7qUy8zxFJWJoBaATDJLa9LeM8Sq/B8wyiG6a4NXdYb8bZMpwgMw2Cbm+vzE+p
QEvXDS35iRx8j32M42Q4kZP0NkTv4gDrAcsZBiyP42+/IGI7uoMgbQh9dID1rsbj
uGL2Y19nzyAMtaiRlofINJWGDfB+fcAx4KScCgoiswySgK5hslLsOULuVCEJnll+
AMJNGOdCNBWlhfBex+COtBODByDDeM99FcxwRjZFWjrrBcMIov+p1pL+fR3a1QM6
K2bHRYRKDKyn1GqcWjaqQLLl8ju1ErMyEVCB+l9kuCd33oq7jbohXlNCX7P/4G6e
tg7RX3yt9DhepU3IDLXR09ZRxfqYXt877qHFdwCxCXU2ysEpV5/Jc0lvDrLphUa3
qHxxiAFQjBjwrv+ENihMZITyVzimRadexRnKtXhaLPpQjawyGY5OEke2xKWdbgM+
B/zyWU5tiAFwZgHHFhdTN98qEuXuL89gHfT3p4rbUOI7kxcd+Nc1ZhfzX/Fb2v1U
RF1T4vtAjHuC686m3cEMn01aGNGF1VEaxkVNWq5Kn4H19WgyXYpuskdPtFkaURuU
WwgkoNqGf/ucMdISapYaXH2+Dt/q/kUVx1FAL67C3VHJY7fF7/IVx+QaeKsUjVw8
cXV6GqSKeO/RX7RpKLxBx7sfy2cBFDUhrRpR+h7r7eqzPNQjpJ+fKp0hQtpqz+7k
9j+rsxIAFzypPLwSrLpr1eRfYMM9P8/ZAcsyEg9N2IA9fE+1Nvr0xr0FYng9O8+e
ICdT+veAK/iReCTsAtF2IGQsu9QCZhI8UEwCStlgLOqstHUC4yGrugz8oYhAUJuJ
9bhS0NhMEypg6Pv/4AJcihqWZckRI+d5MKfrb0D+Jmim7GoZPDA6q8XWLRIaqEDE
tPDuQl1nEF6aNYtE4MLZfQE/mGe66B2SF51f2pXDujnnKYtVXkujBJlS61IwOY6V
60SM5FB6I/zJy8PQ9Uo2T6e5Cckn8gEuZBVkaPEUzKrI6bdEYQ2vr2rITNqh3eTg
Ls8uHCo/qAhfcOYwYylXZsh6SsbO1kKrPdZcEz4CF93shZjBy+d/tncQ6xq7WmYd
WTNdiSnKYefmX/bqxsRZ/xJy669birU87pH1pj/H27jACOlmWb+794EsPYtrx86D
yucZi2ozFTJbjdyudNwDt0SvK2EEEn3bLk1aXk7KL7MQti3tIeWalbtq+URofA4T
/I4eoFjyCIPuyvhxIl9dipHbXd0zzcT3FNn2WNj84uE+gqoNUVQ/NHuOHW8Gq1uC
A4h9+xs2tsOHs7ltvOBBA/tdztTU9Y2bf+v7EuVUJ6IEo3sLh0tiYefYk3UugoBP
jMB0ihPlxtFQemR1N3BOnqxz/8YQxQv57O20fNbDKzVUfhhuehpIAvSDZKKW3mnP
Sghb6OO/PsF4B+1Wg4oBh/WNeD594HwvcT47zcfin2RCtQhGoTuNhGMk6dbrw/sk
PeyZcbEjyYgKwKnoGben3e0pE9ihNpmROrpn9tyXaV5K5ER0evBWcbkKDDPQhFdd
JxclgniWRd13LglMeJ4LkB3R9No0EUKeHoppnIfRbltx2Uszl8FmXk+KPjMsGFMP
lweyG8ZA+W9w5BPHhZCgtGQJ/uvpWZIXlzGfDePcGBOp3fCWKLiLA3xVKXWlhj0o
9HVoupwamPA8qd/OYhS4jiRLZWRtCYxD6OtmbKcf0ehLfmCNPmYbukcMx7YtZne5
aPuG5mpjpxBXNijQYbkvyadLLw1wTAM8dkODhbgtWTkodZXx1YdCH30WmesiV80r
3V1Jg0VTmrxc4t0fJ8dBVoZcDArYONZfADJ/Ek2suDtiArMd+S71ERIGNIIz3mUq
g+sVNAdEIxZbMEV3AYI2MFJbD6TX7gLE985ViHIyTzxDSTp2T5LVM1zJJPcQfUjH
xNhqYmN7CXoEfMuEA9ilqCim4gNepJh/W8H5kLUBdEIv7nVcAWgux7EjvpGP7sCG
y/gHMz7Ccc8+dJv/Clr8GoyVhXpRRfxWCCSsEVtC39bQ3PSnPytYz2NBGTmCaW4x
3vhgpbaz0UdOmWBHlNV6CQ3qAHmPrN5bzuGrwPuM3XA5pI8b/KN1/HQvf3yh4Sg0
uoLfSLYsPO4V//h72sZXQ8ARkzMgrcG7s365DfpYzbeOa0YrKf8gzpCqbvuRORjX
pl5pRuoYUKk1lEagR2Yc8J4WEkIv0ZSWXOW/6FPLn7wo60qKAOX+/glpOlylZcTG
bnbNUZziWfWM1ShTPGHyrkCcVRkk7w184maLLlxtVvc+9A2Ph7fQfG8SHVpDo0Rz
R1Wv8oYUG4oEkmdgtsBO8HoWkQc4/GAB93Z8nbo2kz2AMDz3b0KDMMz/1f3Fpx9h
UZLOq0lG736ykey2dmS4FXsAMizBJlK94dDeCWG3+AJXFwOJ6aHO72JfcxgV1zll
r+fReXN0zbeqejsDdrVS9WtsxV6SDA2lyGi0O54swyhR+AHyoPhy3yhwu1gIpjv6
jhNGWPbZSLl6eooPt3j9q7C0fEshizyYzP1WRvgHi0wm7Gy35xMpWnCW7trcxgEb
kncjj48EJXen/VTalJTsbCqVGne+gURIwgFXa2XNOfRRHhjSOVFKBgKYG7pMnxQU
t0G9R1fy8D4SQpwfX6EmTRgKh8CM/12hLzuqvs0U8RBt8759GAObF6YMM0ych64x
63zHHGL0WohET4prnhEIigQaLpb/N46yV9ttyoon85YrN2uqQ3lM850Sr1/ygiKN
DB0H2CrFXkdMBSgDB4Hnjgpj8uNsvjQJa8cKVwepEHP1e3Y324D+Fkfurc2SAV/t
36N/IRF3iLw+lOJO3pLCXJCiBvCI4OnpCdavJOw0pGZQRC2SnEn+DOXNzuOXSyur
93R8+1C35TFO0VvGQubIJ/14lz9SSEp2p6R6zmUJ98/W3ThfUV4oFE3OjymMczSK
go5ZFU4SFdJ0JZUJpuBzcWUxuJBEI77JhDW3w1R0b2eD1G0SbZRdjFMy0Zm2J+Fk
LXL/hajyQuH7dYz6htJtu2dn2gX1PiFizSk8JAhhzoN0+26cCgMyWGC55f9kOwS3
zTUGdDE4SwvmaFbQZbFvPT4EFSmG/hepbKZxmgVn+HsDq6v1iYh4osBc/w0ai6zX
V8XMXTdVoj3d9vgtLdDiPjreve82DA+RE8ydL6yKUnZFKqxZBZgcRU5zg5RdTOhb
BHzRto/doexUTfQPWTrNaYnT/zJGr1C+UpnQZY9L/7Iv1jKPDE8Rlg9zrAiu+laZ
YJbEw+6b8CZ4A1X4W+g51gWUngsPCu/Hmu+Rn9HSIoX1UdGDH362hBDJLBtZg41V
dU9YIhw/CpuXdP2ZbmRfhK9xvUipRinGrGrVSgxYU9Eg3y7NdWSguvOgd6N6YW5w
aUEhfpQBZNgLrO41aHTVlnv+8cJI+gemJx/m17j3i+1/BnSS5tFLBKDfB7cldaew
Tl3d4WCBfCMpMMyFb3g+HO1cM1aPbG7hL5pmKJlK8oF1/XaInaew/fcGsBLsBU4i
jXV8KQn5SKoSGBh7WypyrL7sSz8yUcq9buiCl+t54oZJ1aK5OljE0OxPqz/FCUu6
1qlco2NmVdzXOTcYl7zRk6R7cx5gJ0neOjBjlUInHuB154+j7t2/PoPqzHlCqh+K
ZTeHW2zcCJOOZg5dtIW6++uo9DrhixVZvlve4nqyc+UIT/rxr0rAfY7yWzsHlqvD
nFJPH5UMo1S+DYqYjLQ3fA6TXOWUqjlNpx00lAGtjVmqT6NuSK9MdI5Kyp5iL04v
8w+GYxp2SGuh4uOY3keHU/boSzfb6m464PTYrpW6WPZfwhz3j+nziIfWPWeaeTXj
a/UKEfzFRU6BXPQMeWInwbZ5mq9mcYxPMsPYdQtKX0HXNPvRuG9AVfO5qAXJBoWA
68qCHpIdpm1P2Rf5jLD4SdnXtW2V44AwJHVg7+D0S/oLAtIWxtvQxybVaLyiEdUD
YEQ7Y/sawSfQYz3BUsxDY73pMlaVfMLo+0k+fgU1BHgIMDp3haRAuQFa0886xRHn
MhHqwLi/m06x43NoSoDjHxhwY1op0ES/MgLFA5wlgSRUI4ntt+uTKtb5EdBgjnWd
54dE1EOQDnfnBdV6zcm9zDKv5woNt3AwBIiRCOWfD68srY6lVIrai7IBEUv29DZl
9WX1CdhpniFcU9rRjT3Xm0UTxSaFgUblUCjUD+Q86TgJtVvZcKSXVp8OVtd3aaxO
UuvxetwpmmyvaA/5YKPdOGke40zXNDgMEFzmV52fWxvLybLoDHFupQlqxZyNbpT3
jeNmAbsqeQ/ebW+tguMte8Lx09yFUrek7Arh1vWrr3atwwS/nsrSt4WCckWU+kqy
OIZWpe2ssytqjdZFFgT0vK5lcZzx5U6eEDxRQ7j0MeqYxPNJv6URVdDUIvhsDLkQ
NdHvh+9UPsPCelfZcNB5eWr0Mha5FpeBP/UHwmtfSqoZsks8HcAB0GgegHFwBJ4U
8HyfORbJ9U/JwGh95+QyOagczHIkwNWOgWo2eGOvGrzA2GbXpW7Ph+3Mq3o56KOu
izXcJ1tT5xTuPNY05u6yXfZEEDXeUf01TnK1dHtycYa3CuQBAX4Q6x8GNqX3in+U
OnvQIyVMdXt96ZzE98so/jj/4+7j6geFEdwzMJ+ExJQtSNGBdSL3gQTnXUwsHSc/
bJEWiowVTQlbdu/xE4FCOJ8H+FV9GReFlKkf70dVs+/AaGeE+RHdkmkNVkCyQTL+
l2PqBm0mACW92LxIzSA7tmSdoCGyfys3rw+AK1RPPXvfaQLjf8KODkCbz4oUdrZa
g2e37rq6ARlzaDGrN05AUfUtmdArVNKtJ7HTfJhVry+THYLQumHh7Yj7xYrjZVC1
v9tHpzsfTD35t1Yn18+UmIPeU4v6M3E//zRcoWJkfbwCGx4o9+H2WwVV+sN7fShA
EuP4dczFfWthl5oB57wbvCDk2nzcE8CHJaN0StEH7VX+WIFcSMHIxGp6abseGQl1
7ZJIwMaOOSZ6KgBbtiviFCps3wP2o1eH/l+jc/wR277dUKG+ArOXx+PogfeCVoSN
9R2mbjP2RpqQB4uP/Jri4YrVvlT8bsxw6n2U0rsq946v2JTnAmjkqLH5xnmcuoiJ
hYdXY7HLwGu1Y/KMkdWorOimbH2yvf27ciz1bWEqk+dwn5iLzIErJ0LRG2RhTfDJ
5BvbQ6Lt4wNFbHL049PHXo8EaZXpuLtmYz9hEp5eorjdFF9j4zRKSlbJTEMwwBd7
dE4YlzQit3WiQVAfa6hLf02y0Ep0qToMgri48PGJcJsaW8g1K3LsR/JxYSRSoFa8
Mg1cTnubj2DJVWbgTRdaknlmmkqFYJqtS83OVL2pAlc0WWWeC0sHOW6TRwHIlaXL
TkPQkVP7AO51befLhJO+I/FSsDsI7PfGCSI+/NkyV3gJflq05ndHAe7Jb2IwXHo6
IRCjQZHXi3+GGQCghRltnIe5qNFJ12M9gl5OTYmHp/AR513sgv8lvYDwvyvb4QBE
Kz5+uJabh7gWchQCiTu2etn1dmheZULMejtjlvB7UJdoIbtK01UHg3y7BlkkK6b9
G9N6HLnkAqiySQ0K/KsTwwAMkY8yFbVofAPouxJ99DNJGlurN1yYi6wf98UlIoWg
FJlAGUy4M2YzB2X3eiYLcmrlhyEDZuvEMOy3xftdUne2oI3+EsAVPdi2UA8mWwkZ
YEgdj3keCoqhgUWhQuB3RCEwQMPePI3fETsVTo0fSsI4V4F1k1frFTPbWSQSd0vB
nWTI5ciL/1cqUGdz5QLNuCW9MU0FYft0BtTtnOjaOy4EoNAs8xInge03HS2xofTt
VqHV9aQwvft6Ov7WYcr9kWMjkocUmz5wC1ntfo7cDIT3wQ+iwTaX0F2z2YdUi4Za
MRa5LOyUA4hrSkkI4OZNtPo+E/VkEvNsI7bgSp6cqlXKOyEuLntNy4TGpFill7wE
OHefL8YknT4lluXujdo5z2ztUNCq8iloiujMXC3e/EFF9mhyDiou8DXf+LrZAWRw
sWnEff70t9mq9443nGfsDMA6b8RakePC+69SciG84KjPIsjiVD7bRTWTeySF/fbw
WvwZuFTfLWPWzIJCnuV0gY+pF9s0NAvnmQYR7T0oN3p89FrihGAPiMfroiaSDoHa
PTsWe2JkeCX3d+S8941hyXyXTDFrYQbD64p8IAX7mYEMd/QtDo0mwJhCzbtrkzRV
uCL8+0yvcvYdBedilvMP9CsL/bSHRwcFxThs030Z3c9Ax8imCBddrTGTwuLaG+Js
0ZnDe2PN3tPqTG8UhP/zIHYit/jCj730D25fWUY7Mubzd4BjbtJDsRX0RS4kVifn
1ZVJO3qvA5iFvigTmgRJwv+YoZsXn1ZAK0q04/0uub4+sfKxg1BizDR597QEKTC1
SHNpOfXKtAZGz3AkqFHo72SU9iKFnoYVklYIM6nyxfQv/jmbGs4jkbtU62XQVkng
Dzcd8Gv9shIAl4Zg7VUkF5Ah+GaBrQ2TvUw8uFkKivAGTmfi1APbdaykEbAtka1I
MIfGzL8yynsYT4O+blXKwP5LkYJP1qFERqJxCB6DycsrkhO/yoG3BIlw19FHusIr
5SVzHOAWRJWH0CDyAg8KsTyDXQksc0Qgam2HBD+q9ExcAenlfe1wJFBTXEXJuZlA
Dl0CNn5NG4cswjoZoZht2tbrggvmoZ5mcPd1tJSX+WVpK+JRmYwI9EEekFPHln9u
v3n2uTeNBSDyL4vB4WlKq0hg8kWRQYaUc9UOvtpGFUVfkMTGo6RWBALQZG87bBX1
4tX/MHbEl0l5rxYtO9UmXl5XRIQezd/h893x/ONZGUMVVUwxfeKjVvcW2TuQjNmo
KVxfHmYm411l1lf0ee9KguETUoYzSS9Hjxhbz9DuGvdFIBImEiPIEjiqQPmvckeK
JwVIaYMxPboxqBXkNOjjMbHc0rGLexpr3AaZPJmSV/zpFX3gIeVWNeHuA3CWWL6a
ybtw36x0xJq7slAXrSTPv1cn9v/06JL9q+pfu5wf88ayGL79ZFx58KpEmb2I8sWW
8PNYqm3hOwnTP83KW9ih8sqSYJfFxZ4cIAD+Q+I/dl4nSpC5U7MZ92iD2FwoED04
iOT6U51PywctYluiChpZfKH8R93sipGkvyaMd/u9+R+1hP7hnt/9ehBoS8EBZ2LZ
C2ewnWL6cfpk8IdCy41onyymzSHxK+3TfbYuaOL6p4A9gqA89BCSaw1BdVUocr6k
BYHO260GlsINLe+mq8ojPe5+nxYcjvM+Oa7bVCmjAG1dXb0TLKwWRisQpKoEM0b7
l0/Ru5ATaM/1fDj9FOGXln3v/DHDJy5a1spoJovtLR4+6KNrCVCZVcKL5O4nqt+A
UgqCJhDdiNwKQEdsAA4TLoXOpreZ76BBmRjukSAHydP1PT/ONLSSDYpSbtbuyErP
wIO+zI3ErUm8D7idvihQG81mwlpnP6fSuh1cLrhbbd1FeIRy/peNgO/tJ4Cq2YnH
qvQkH4OZe1xx+qhE+RhOIPuxahUwtY8PjoCz+FQiIIe0xKe9hrVQH84ZP3d/DQNW
H+h0AQbwuT0Ty+KADXOJeP3kfi4zwiob8jarrCklXzTvXPHx2kVN1YEBnv0AZLXb
mA0gDqVlNaFXTEMKotaLzSfVK76KKYdPvwfYv4jrh9pQGUnO4g716Db9kVOg2m1y
9UR+C+FPnLYnwARzh7MgUnAVMM6o9Nea24ggAvTZx+XNKn1P2571aniOHfHWQ5jR
/GSoz6kDMstZ2tcuZHRl17CfvkqNvvKYAJjct2UWMx5lR4NZomddJAqdAEcF+HFt
6kSdy/EcxkiSKfkhispZjDAnNu2mzyY/M831gtSwGMSu61MBHSmGO+Q/ugsMad6t
mSCql80UVjuxw5SC94qK0uWaxgkvyR03RgFtgx+6tJBSF7FXzbT/S9x5RHXgB/EY
VsB1aJyDfqdkSkcNeYqksdTrSqqCRzJhswg16d0oTDneRgT0mP6eSYIgcOe8Qmbn
pfk98eHe1hnK4PG1Txh/MPkS8EcUJlLwrSrDsbOrtEfSToIk3Yxhs0hMnqYKsRt7
rktVvmGsB9Ntw1ckug7V3ev3GM1TD64f3RAzWz0Q1PVOGMg5Ycr1Fb7vWefRYfP+
INzalmvL1OwryhK+DBrccLBbVT5VJ0XV8HhDYpNdepPWY90KeT7BQHf5ES0ZmeWr
5VcUTdLv1DjMFkloO9H+WbJVfvxEg63Ftc+mQdgWdAWsZuxKSP0ahn91aWq47HAh
6nhpusMcvlO6Lt01L5HOZTcQuPH0ztVobkXauRQ+jAAotoe0TuHALIwr+oCkBx0S
YY46ZK16iPQsXiQ9hl1SW7xc60H33SOB0aUi2qCGygBt4oFGC4EoRKgMSUa84X6I
QIlJYQna1YAhbwYNZ+1d53tE4MSKpP151BqmRwNKpnHNYzCS+mS2BMDob4zQVA8n
ebv4x6l7Sni8XSg29SU/rAKeFpMRb+NrKMxMyggmJwWx/qf/pv4Wv0FkHR1NudK9
sORRaeuHWmd9ValkAfDSqhE3LpDxcIMUucr6P4KrRMu6z+jbdo5Hw6nqjKYr3E0o
hJbccNGTWl7OwncK56s1nrqchsZ2rv707a0p0jmpAYuLh+ufMEeIfLEn7bKaQNXF
KqOCq/kIQfK2oIHLNg0PgdM8h8f2i7MIpfeQaeIEhVzTUb8SAay4h3twb8PQR2Ch
9tG1nXMtdXIRsO6lx3HGyii1k3lGOCaF6miNJBNlUvfFlf9unRNe3WSYD3scb0Wc
QK8aXmDgslgpfqYYTcRgJNh9tDQhC7jJ95ICuzWC3PCs4Rjysq1ktNFunel2ScqF
0iK4P6Arl9HEOii1XMV8HLhe74CAutoivkup5yVtmCTXnXe4X3XtqTkeGSxZWYts
pMKwW3slRVnKKBKUuEekErMMkJ5fJOYVBHInVNrMTR+QETXQd0xmdWLKPxhyjEwi
bQ0m8y91vAFlJYRgTQmgzuN5SFsysiW95mCOYrgl2eDkLYoU5dberGVhACEeE2V6
d0u3VLTugIH93PK+Xk5aZT+IzV4ESzGYHSJ+6bWzSMOx64/HgTQ6ZJCiTT0o/6Lv
Zdx9vdEV2cZfb29TEkORqQd8GEnwU9JnBwr23L8cau6TfkDnOM6A9Ppw2xlpd/R2
CtUVYTdBPbD4epiqGCauxOi8ww7W9CHWNScxncf/BIGWj6QuufZ5Fy5R2ed24CAt
fZjDhwXUY9HYabuKAsdqWOfoqAjQyxE9UfUUMyEs4Tzp1M4zAiSw7wWW6RYM+tqX
VNArg1uOoaSsPQfNvuOBxuIcSjBKH11jyOEndp7WMMN6cK9is5txatL9X5vDti1K
FKkTMjanrFlYfqvSEoKXnCjPpY/fo6Fj+r5mblW7Q6hujQ1PmVGrkliAh07WgSqt
bcHMPW6lqygb/8Ho+J5vM8jWO7djhABgUe4euAh4LDOSm9X//L+JL9lrFCP58L+u
EppfOb+E7gZLY+vcOsKIGpqTvWhUAbH689x47Wq0uVnz0Xs2gtmzRh81MV6hYk2N
ZmeNZnaHg7c6U6b7yDlWxOkr/vk+lEdDmgXhwZpkpinIDPQF0fF/9rKLEh+pSOVc
svN8hbeFZxR1rSd3SGA6Po7bxmDv2Ge+qz4lJmXKcgW4F/wg+FwLfQ382mnjIrdf
o8Kor9ebSyzqxVXxNZvYnur1j3YnpvwlUTH1jc/dZMefcuccSEay6Z60isT87P2u
gXyQtKpQzeZfTFI4z09xz3vatGYoS+firL3lwfpKtlWe8go+Fgq9Maw1KTgalFrj
QoHGG8kdoKA9lwk1p4BYykEdJ6+Ho9cWHENEdgkBCIkhP30uOAEbDthtZl4XmLLD
OROJpRAYwplpqkj1arUjxuBdMMzn7G0oePdaGa2ya4joxUztO5nptn4YoxoPAcqa
I9N4IglRHnDwQQ4qyTWyN9JHf19EpUpqUIfGPfaIQHGcFXp7dig267ExoJTJ0r0h
HSQmVlIAWD5KFMW6bPIFgjOfTcQDyv/GCLDcnAEWChyG790JiMNz+hsxxp0s7BBE
s8VoTrZIEaHh0zMy5SLsdwtjryiJAgU7tPg+PELfYUtZZ0MOZZvB7eL0NZLXQY9T
uUfD4uT4lMGCBXhTTo8ccRHr3LK6LYelr5vnFilKEqyVbCGmg8E8Z3jSIlKdAivZ
PXmNbX5SF+PSGyoFOwNhTnNuJ9frO2lK5J4gH2czr2tAvfDabp4vUXDi81SGk5FP
nBcxgtG7GECZC7oVWf4AsgJJtrRrxsB69YzAaf+JKkWqGAFYRvTWtl2GpBx06BDy
RuVPYf3rapKmz4w/+IMKt+AzRBZPpukVgf1SDp1FGDiXjYpys4oDdQ0Yf0QwGSid
uph7hsEPlRDZhR86dnky5h32yxSPJTjFMwcx7E2RB3Ur+pI4kqEP/fnnX8ztxsDS
SNdHhMJblLhuzYOV+uyYc6GYb8hXqAeW9VMyj+aoVmIMQzkXzpxEAANhvnDuClxX
CR9QLwHj6QNj3egfN4CTSY59tooofRzSBsZ1ASgzQki0STTey4dvny5FbmxwNwqV
/kSN4f8qFGKGfprYXLZz2Xi/gS0IS7lip4YBCrrruHbQ0IwhtFPkLAdprxkkAxZe
Rnq7TID84/tUXShAcI+NxTqhy/JjnFijeSRqLYQd2EHg8W6TDSPjvanRcNU3t5T5
X1asvWqcSnYOi5pK6XKJ/xBkglmcGhwi+NRhtRD6+CfLMs5tmSZfR5zykDkr1sHM
FLG6DYbQ8Palu3rPA5M/4XtPfahatErcbif/Sdc+f+dvyp7srAbEwy/ZIjb++BVN
ezvtkCMqgY71jDjJzk5J4RY0zqHO9wP8exBRUvVApjaHixazLyasVHt6+uISgH9F
cfsTqOQ94sKePKOJnT6t1pwJmJvDhAWN+nqvdeMWUvl4OqkbEI9U1z55d1Ztv8cu
cfKaBvoLEnP7b4xemhsqTXhWSa5vur44ORIjZ3bWms/yg9F6jO1j6GDd1bhgrvFC
MJWqy6sTNcX+owyuYLLZJUNiJS0yRgHlVMjBAvXzYsxj2Cf1QU9Sk6sjTLw9tdkf
FZm6d3wgc3D44GzoLEbAXvWxdAyoA2UleE30p32quhtk23CFBtb9Pjli/8iSBVFz
IXGhdyQRBAL2aIfwuNdwbRnhB5rE1hCEmiStkJrcebxaPZqWHnlVL0jmWr8G96E4
IBshoZ4/e3GcGxjQe8wcGHTJXvREHYuNsOQZNuFrmH7gs4VkJR4r6QNBEeBWARTZ
lqt6266HiWo73ImUj8h+ANi8aePIJdr1sl/6NZQGIHytnimF6Ba8Ip5fP/Xw8PAT
H8smGB9NVdBL6WV0DQUmD+y+Q4yg1Ly/pL/BfNlAKWALkwGSA0YxRlkBnhJ7ao3h
ThrtkZDGMfg7/HAUKUDzynkzgJXr6JWd6bGZe5X89dq6ciEShzcArElfdoPvPi2/
sLK0LWfo2qjFc0bwu6iWb/ykskVImbSoUSNJmrpjWDDHVrlyPD+66ZMGOUco9PnN
rQeUEcXIRdXMBcsSz+MvoPkXw6Fr7/YHPVKu9G+FydM2XByd1kdpPVZx/BaBoPbw
t3vwKRBCeuif38zctFZZ/z1NMfwgLiaHPh1CQ75F4Qq1J4yAeO7+7RvNUtSRunFt
QHKJEqAQ3cnjwu2cyo9riii/VeCjlNr4Qq4ZUVVZY+ws9XoYMHEN7OuIhWCMfNed
cnqZx8rqMVlotTNMT/gH5lSrXsIALhXIzX8/o5YQ6ujL8xyKtiIA91XWvFairptv
JwImy1BrhTMuSkbRJKbqs3T5L/syyvzKxIzHNwspLS1FeUduJ6+3Ku2f1LdzjKOw
MN7J6msi1ZX9DlXWO2mEQe81LjhufhMVs7pkpRcJG6crxuBrZCL2KABOEmEhJLus
JxFX/ByO/Pto5Hj0zUqvszmaX/1oQEjHBpA3lQMVzXz76uOR0sKHyFvtXlnJAlOr
QVUT6Vovha/4BlhmrFFahnuLsJhjp02RTbeoLLOl8qzAKHz6+ivkvBYL5TWTpix6
wq4Ed7qqYL7y+W9mkaRaQY1MWN2DO+rGsVF8ttnTZGc8F1qZu+N/iCxYdWAvmk4U
a29eEh0ZchePglHOts37qo+xJpt/jfGhdWPJ+s5G+dqR2duolNMug59R0+i0Lsyv
+3oDFxcDOgVNKpQFGJV0RiXRaf/R97mLwwBK7MoqCWMqUvfcA/ejPsKZvC9kLN/3
QDpfhL85IHpbjSUC08dzCXyXixnsGfsRxdx6/XXnz5F77wagvZCnNFdQ+XKFBPjl
bmOskFIeYDrNs/EKACxFWJEenh9yH2GY6dE7Q8Btj87J38rmde9RV8qtToPlVqot
SZTwDX+PM+TfTxr51bkhfN/YCPQdVVfy+GFn5Fx8WEEf6+K5ORD6FRgsTYo2NEhC
GjUcaYcfTDIGpGkyZw95jJ8UefscDkysJ1CIVilfHF2qV103cSEZqywSDdTLHb+5
IsE11q87W4dnFOq3ZlHdAOXkd6bg7x4aH1uD0CAVp2ufsEtQqGOFUJue1uSShzmN
c79F3R63wH1Yn51Jf4RsnZs7lKzl9+oPkXHpDandzXGAQy4JpVUOs6xc1g/MSFQn
4cinVqNpIJkJAO2021Xk/QPPD24l0DOBupxnpuycz/14GcsBblSP+J/q8XDd4B6Z
6ePGH9mZ2sUbj17eE2lKlhwwI/vAGbggw0G4xjvp+HhRnNhogFPSMZbMAyilysvn
gq3lIseDrPYSHLMrO6UPtLQPFT2qhiEj7jl37wFHJgjDdqqGX82FM/DMzNpOl1Oj
Eq4IBwm0WdLLRM57KYjyW4z5LNqCChnW+O3dhf4Kr1S2M8Tp4GckfQbDZqpEWalS
sEH5pUNVrB7QZd3iAxmwJ3IjWT51NuHA2s50R7/vzjh7cxfwcpvs6SASJy3z//yH
Ygb0D/F0wYwzvba5kPptvqLMDJAQicyGNEcg9kiB4zsMaAMfs97tLZKaWFezV3vW
gDiszPpxxv7mldsc0SqjIfA2Pe3CYUGfS2hECFl0vwvrBhkqo+M5JUy6mdgHBf8D
SscV+npkHfiErZnQZJQF5e+CFdVoPoHJZnSEB89W5rKY4JhdL9P/13aRBLtrcSva
AckD/quAwd4NmJyrGg6wO+NN0tMpWUd98KqKdKyRIkvWyRNP97qdoSDz84hJ6w+9
2BIvK62IWZYgTOW6dBRzLd3reJ32AmtcqtiqUL4GivninkZcBAQmwfSNYPv9I+/K
yQz4H1VDp8Xz3KfpofCTiNVAEeJvRtMJOcIiquMlQNVxbwLRp+TSLL0/1Umq1ZMZ
RLOHTvlsyBLX/Kcbc2uIBFs3dgHiYKNS/uqIgcb+mNoDf+Kopt3jFxU6Kza4zeKE
MZZNuYrUSkSLQ6wnhaL1o87CMzTC2NxRsgXw4sZo7Chb6PuaejZWGpy9YXjXcoqr
cnybqeA9/n3EK8j8U6C+m9wtFoAO08HSeifOsSkUuh6N1ZS7VCqPF7KC/8W1/8pd
mq5zEH4mVnsCemZ7cIWILpV6DpnjfJZiRL/cNgowqFr3IAUqqB79Ejs6FuPbm3jY
olj5+nmE1aqOfqWBNTwRxbsOJFPIt4dLFP3qFxISkrYlETvwmSVD2X0albHXQmRH
rLWUtMsTzz89GQAUrvMwACcNernWcDRTf0S010oXV5y8Uwz+3nFzzUX7I3A3Kjpv
f38fTRTDJIwTzJ/HyARdgjSuMtUEzpgDXhB6/FXFjdOcz7ev9ayYfpVpq4k7Be5V
vFerQEfBr08L09+qjKKDu97HHUpZ6fp57/i6/eCWU28dAiiXqn9CsSNktXGbRIwH
fww2bo1luKbvAnZiBVvGtQ==
`protect end_protected