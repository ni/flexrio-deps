`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14608 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0gQgIG1mJzulW1XOK5NnZR8
C8XqDUtXW7uOWTnSVqbIblwOHrDC/GFb3kYl7b/cVSQLjXPskjGSeGtgjRvW8Fwq
viNejN0e1mebiHGAGvQK+ksnDZtnvi8HJ8ZAyZ35py84adBhmbRyhxY9aOXihvyP
Hfuzbm+QD41P/moG1qupRR805KWeVALCTpHjLe5cIkGqdoCqriUHMQabEgR3henU
G4+FrdWIvvtJD2c6qEDNWKKKEnIEYK1+qL/8VF3AuXksEAzPJb5VGoZxH2pCwSZs
fAn5fNLtu/R5ZaKBIcNCcwZk5ucprAo/09qdGOYGidjz3WS0Gzl3tu2IiqLpJ565
CqnZ0siaYsIGy5lzHOLFgqZU624Q0RePr7DK7nti4LyyfY4chcjUT4sBNf53pG7t
Vj2x02ERX+rtnVIHTX1AldVRXU95J5SbLE/FYrbuuq1iQbTPB96pU8s/xQEAkcgR
U3gvxowN/XsUx9s/71u+CiMWYhFfsrr5g39ciPxwDEa+oixSeB13VwwN7lJGA3LU
uXGUKfBsGFONWaA5RzdvS4nmXqJCvqJE5q34tRvFXqHw7A0BJbDRKjUDGF5p8A/m
nuCDbDbRCPSlBKuQ37JY+ghIddmUJTaDwWA8O0ufH1KAx2Hrh6rTjfX1uyeL5y5N
qJKlFvd3mVTDboExAdU8GWEZwRhh1rZIGxK69tKpYoSgzaQJkGWkdkcqeLssgyuO
30I3GymxWfC5kNh7reTh4Ow6IhhcZBSD0RKD6HoxHZh1uYo6JzxaVnuhuOY/QEDr
/VnK72lilui/UlLc7+XeOsxnC6xgApDQcE+2uA/PkcqR+92bGND2zmv4kQew/huZ
m5RuKYEqX8mtbDBsSmap3XGf5SvbfBzf0OUZTsKIqexqj7vHO/6rMR9HuLbTxOFN
pQBTic3sU9OM0cBMa5EDbQ65B5THDkl4dy8FkiTpuIaxxDHrT39RMq51jBtgVPD0
7TMxfcp4X3fvmTOVc+ZVx3lCJdwH45wY6XQlnCNJm9mGHHzor55bt6APkmALMYlw
WWTHR6hGDSje7aUG8zxSgrpnjDDhDHVtr83GS8OzcV1Cc3+tBdiogf6q7MtKpKoe
40l9pHBOvYECkPdwYhIhcm6KsqYNuXHpFzjbXwKNL0fnLEwKcfh9uy39hICrrr2u
iQhZbQ6B8gZfkJnsGmqQzbVyveMUj0W3XcrdaDX7pY///qgepnBtfa3k0rBABySb
EmIXWHYMD5koAO0cC+pW5elaOPNXgahV5hIxsFNe7IBNIn8wi+9aThvf/IhloRuO
ttcvQeTc85Ac6+q3jNlSo/Vp7oKyPcCRimhUqJdfTWEgRsFBPesib0SaeTlyNNeo
4kFRqtpxYTeJ5Byf/zsSigTI7wqPEy0LKHhP/NHGAPHctaYnLPnOOKGgbhNhM1Dz
f3soFUrHabmm+Pn2x3ElehnPcTK+uTMIQulBWki/lZYTJX58FLCyiG3SZ/ynx908
MsFkUIDc9Zg5X2u2fnaH0xpOa7wXALTu2/W93AHxW9RplvY8KqWjSbQncNUE7Txx
kInTN+bToxXFKgSbcPBYABFyX95jfT5Ph3ftqCDBgR8XnlvoxLny3EWywjXSn+hd
sxTHodmXNBw4o5JxQzwhnFlR5DzxUu3IsNp4Sg66ObFJXOPDpKUk8K6t7SpQu9tk
qgYRV9qkT+OQc6yvCixLPIHMDAecTJqPlRnaNI2MuBc05jM3+Q6dj8SejBRr9sED
+xiD/TsCQAo4wxuS/r2zN3GTBhX3Z8GqdyGJdHLJU31VvU35NP4qSrqV17J0uLNW
yhNM0mBlBHI8H49nQheiwB9J+rO+07jAU8/uAAeju4oRodFkTMrtcdOy6sMykDyS
gd+nKAoAYe2AMwH6R4JuCTdk8tOvJilx3l2bVcQdGdUKli6pSwgCUCbzMYYqk1NM
7N8NEeD2370EhvfIYPfACTsTGz6WyHtPYw7X7k+UQM+vufWwlS9mkePFX31HuRS2
upaI9l6KocVio2u0To9F4xNFsucZ7owm3ricqJ564VmYvKaSEecEx8AUu6+AYJD8
6JXRFEJ4dCS9ve/peUmon8M/b4ydPcHqNGP/qll25Wl44TnkA3Syxe6L8a3NAuoj
VqObpe95Mq7Pp8Xejp3UTGcqscCiVKCMb/F+YNMek6CV2HbQ/Adbmyid0tvHQYa+
uTciZ+Uj402jb9OrzGfqh4dSuIKbdYaumW6JiBu7TMgtusGoip9zns0fIeGtx/j9
5pJJ2x+c5wWSF49Y7jAU53/s6+3ntP2WVdXOycVK5lVYud2YACFknnQIUTHiin/T
BO4Wf5Gb7JJIAyn0VCPfB3Sxkhb5xza8/Ga38u1cuR15qiM0YdjozuMCJ3bUe1TC
QLvBCkEdmk34aLtnyMUdlHinxXCdypNbBA3kZILOJyTwCVsW1VnbWI2pyJLLYatv
QH7I0q3T6mu2BXw17ObEvT0xWx4Mu1YoXFgPLcE/7Xd9s1k0h1N3+ysZaBhuhSBn
8mm3tgjlnW53uwqQ9t7KHdHBO6fzYDlbND3z6cLj/3EYU8hwbgmKabAJA3YLvWn8
OopGe+vPNTSODgJhfHeBZzx1Amdzx2qqvmkHkk3QWDbNYwNngali4Sf/8tvZXnF3
MuZPMDYUg3hoFQ2TTfg+Ly0B8mmgpGfwk5STCF7FnLLWI9Ax3CHqEEz9HrBTmfFg
R88ID7dKaYGShqTizWYfPjJVl+i91Neaj0QFsSIJ1WksLnn0AdHBjSCQ5Xl8UuY2
JpkerPOOtRscy580N/UHTbJXWclAqpwCPMoBJJjtGb6QbQFvcjp7daEzacYUgZvi
oDLCIx/f+zmJxh2lxXjArsYJWDw9Yzu0SB57gAKt555i+B9HZbWLf5GG+VvIzAtO
ZDPDKDgTROZTL5nar/LYtNUyl0HUPH7ZOAah7jo91yk78v6SXcCkg7PLZWiO48zs
H1nrAilSMP0CBHJNryXqAzkWDenqqYrExE07FSvt7gcMxZQtVACKewRK8QGJyhID
F1eCDAIWMXfQLwpWw+QaBnxsmR818FQ2hUIBDu6hM6Z3wSLGhjaablIwBjd7Fiiu
2/7eodKc/TKsALNiRrHclsz07Vlrgig5BNaNRX2mKgL0N/SbkFf199uAi9520c5H
V3mD3x9YaVsElNhli4L5xNXWhJ7afH3S57FJJG0ZYgKwtDE75XAYPy5ygM2k2XtF
56xThkBuz09OrRNvqLk/vbXUEjM96T22FE2I+levuRidGmIQS+C50uU6EAXDFfMz
iXS3t2J5RDIwvUIXNvtOiDaWmJvt0cnlaXVh9Nv43P3ZVgDBP4HSlvKrnNX1fxFf
ZjEt/DTsRkG0dE84UV0ptHm+p9rzNwAdrjVyx2tZZB9PH/voZ06u1U5hlgOaHT6p
SiSLXqEBN0bok3BSM9aDT0rEw3mlWTECW1IhyQ70UJ/Td8Xb7PpFAqlhnZ33FJ+r
MW9Co6aySj1xq1G1uNEljBRf7RK79144YcDoiu6DxWzwkD6legWv5J4MLP92dVlk
MbhSRUzSbAW70yETRt0ZzM4Mvvmafvj4vmBYftl8UCGckGQlOcufiCjSjbpccRwQ
ssqv+I3MgKsHGmON+gbbpotGNx2mlZC0B9N8rOvhTS3jz03aD5vwtOF9M/m38jae
TPogIhODMKI8/ewvzW0ma78cqg8LOEN5o5FMXeiKgmt0UNEqeqIPnAP3T4TuuiOS
nWFzhci9AisH897/k134jFECvklYzXWpF9t9+Ezv4690yX9Lt9NY7YuTMNXkDeMM
1tg2+PwYjSwYrVRe9nzVI18MjqSxCpFDAobTsWTiqsVgVafohq/uEqwq6rcObXqo
WUqrXx0LIBTRzh2afg3hLTHFtn6WIWsnqFdWdiNTGAyWh+rSnBVJH5HC64Rkw1mU
TabkzHYMShB/wmWqYZMhCBOMi+efzmpNZ4ZjRtAmmZtDOLC2ha6p9zOH4mDLfXQa
gnBmQO9tKD9H75Re1CPKJhn29DuBKeCvt2/WIkIyD6SNX5ZffrLCd2edddVgQTr4
syH0W5AkWJxNrVS5Ks2FUCfQxyYVi0izgG/yBiQGjKjBq+JLYI2Il6RzAN58JHd+
RUndRazmha5+hVaHVF3GYRdkJyfpVgKSIQCg5dZSRzo15O9MAQd5L8xHeL/hTPHV
pEyvXl4C2Ihkee/aEjsbuzfam3UXssecpES2mM5ficmXUxRknCkiN57gXQAvnaR9
AZ7Es9LTe2NbA4J7YBmqc3yTV6fXQGkAt4kb4eQaAOFLEayE5qLI6O2Anlfc2+UX
wozl+ozWNAoKuvPyIyMcEonylZ0v76qSWV5vGR3weMIc7UVGN3RthUzr3JPzN8mh
WTJFOMQ397S0kl8QwkQf0TyvPGd7XwwwuuRI9lx3EaNsAvKtUbB0h/Y+O2FK6xxa
Q2Wy2bfP1M9reTYQeiwHPZwcVvedXL44XKKRj3O4IKPyW9P+PPU0dHMKBfd++GIS
PMBPMsUuSZJgjPJofqVm1/0nBa90627mP8TIo3xCwe6PTy9K2V+P5TQYP7uqLoGk
4rzSEDykw26GHtvwkHbrwiuwU2ItRSUI9yBf/TP+QBQUWw0YGpXDfeqi8Ju9Jhsz
rd2xGUO1ogNkKu1mNCzS+6A4pLi152Nc7F0QLon4vHR5aWztxnm04XvGpqNIthgF
B4FtlMeU3qH6jj1AhMxgRyeSiFGvHoYQUGVK6eyA1mECJXHRenshltDBxw6+hdJC
x+vd7JRVaInKBMxgu+JmxICjD60aHrnFdTUdfYS/GKLRQ6RMHQkq76o0gYB3GDSm
Lia2rf+OG2lufKX76MsVx3fT5sKqLyr0MWgXMWCPmJ7v76GZT4gpBjXFMRFzmrEP
ZAHhoJBtsr79kg7qQsNdX5PQXExI2CcNU5iiEKXDT4XMm9Wbs7G1aeQy4XA1bDsa
GmJxfEOTgEdszk5dEZumyb0A/+lalWQxzUEfub+8FVL/Q7+dUK+8jkdhBHE2lgRV
YKxqoyu3ZiWLgqq5FqwRB/QJbjXmnbTfCragmRQxTiV1Nh1fIJ+K0R89EXRtnJB8
lGSR+DVnZ28c5VNWQgT/H61BqrIlMHbirTyYxK2UvpZG6BZBRl7FrFthE7R9yVHQ
I0H1f/EN8bb2MZ5mjg75UrxvciIr7hbMyg6gE1kArUIG3sT5X5Ys7XZqM9lXZttI
PPjN4X0mmRgE/YEdm4Fia64Rj/ac3K4ZHYjJbIp+f9MoUo+vATjmd22N/9LA6MwI
L4W++wtykbFSphU8z3zkySjapQ/iRiA+47pCyW78rj1+Id8qnyv6w1fqsvGoLyvd
Yny3p3OtNd/+MXsP6FxsT4wX933c9nYAq2aV6QPnph49RIqaQlqU3ZoMSrV/xxVF
FAkxlDx1hWVPm/2wUKMTo7X/EVfDcST8OHmDWLio746wDw9CKWNgaJ8/Y34Efxdo
KMu9vs5Vs6DoIIBvEGuxafTBAcbWEcSfIGtlbsW0OO3FMQ/wwQEobj0kHmvPLFIW
8ynLdyt1J39hghVvmglvEZCeh1KiDWZr2GYt5yLOLbEsvHr+vwRpi5L7ITu2jb+6
l03s0gQ1EBkG4PEgn0K8l3vV2BTvoPh+kVnLOQgWpOq0FAehUnp3CKAdbBhVa26A
VIS8XDTRryxkKe8URl747fnXZOvZ1NpkGZ8lL0LX/EzCgCfJDFdSI/tgL+N7WlEm
rhW2Iv6BNMEPhe4ZhnLDHMAwjhWyjNw6BUS0ma06SbALqTZIR8vXt4sk2uP9v52d
R7ZDpavIWI+KoHhkaBJPqAAdf4bzV8SKaYwMfcNrhG/nwDRLqFwPMjl+JQKGqzPE
ViPVf8qO32tX263Dm0FZt4u+Ve5WOtPdO1bmWwyleptH3mbFH3g3CnMJwf02aybN
nvHBzCtemY54BXP9LAAS+5H/UggtroSIH/+PTxheIrx2LUOQmz7Oru505/vuQa32
e6cFjI2I3izRpYvrItF9lOJgDe0faA227wzDUpfyqjsmW228H/BbJEwr3g3QQdn4
uA/oq/+n110NEpmKMa/CHietI/D2CJuS83jt+bPxDVIMH4Zopd8EuB5825UhRqlj
qmuVaKJyV1cLTMlLYqcYuQeV5QV2w6aLHj2f+DjEzFdG1AzW2PPS9+FmMpbkxURX
L77BWOHxvH+0n/0bG5Td6UWdUItE9EB2P33HMEEgDuMKhpl3wpcCKK1bOY8udFQp
Xx3Ko4SqNIjyjNSQ+cYalO79mmzvV7m8IoNiXJmP1Ezq9u0eD8RsyJXkCEDzq9Wq
fQej5tfvn/1e5lQRWzuwrzDSlvg64T4VjXFX+yb8CWGVK8dxC5eQfZWshHvxie4p
9tT9R0J3oGpcKtCI08+6ZLPnRDNEC5DWGXNjGpsRdXEnD5zfU+S62KKb50ZFFkRe
UtYBkPRvcCnrgAx4ptDoKOZ9B2iHjqLakzNs2MdTKnSMnwIuZJmlP6oXVrzXEe5H
bhRmZENv+zwLwh8WtyYKL1ivWAgHKlUH1mUPxGx6rg0X9jec+E6E0+1cMv2dQ+z1
/U4MGJ6QBkOnwMJdGgVrs1/NLNPyjVxQZKpzxjsdquvcJkOoLhhHQUJAVCEmKzPc
YcgKfmm3dSuYkNXmCkZZcr4I/gy9FIM7DwCdo7z6gRGo77/TU7fIUE9sZZcpYlJs
ppo/946VAxL/fWDOHLA9iH0G9UtQibSrqV8Io757vL8i8HVbXEBknySwupUc3gSn
duvASv5GfPF/nFhJcp6TAkD0zTI0rfS7HLdx9ChYRA+oxAdhRjrZ/fpRcRloLucU
AOs642pdmXgRUWMH4wLERsuR37ixM0Q8hJwQtwMrOUZUtQc1GC/dhqssBuEwMbBY
cCNHOpVLtr7mNr9xbdzbovraxANpYCBCPxAqLHXnGvsaxIHWX810mypE772rKd9U
RjhcCrBD0WFLcbHkPjP/ipCUyl+dIRp2OWx+j/syIFjJwR275clsH1Pa2MyhTF5p
4hz/xPgTZzWFo9e+3w8IKABDF5CFvqXI4LU5yGss0OQudR9eId7DIeMy+JZ7+uZ2
ekVAZT9SOs/kHl4SlQFYxUbm8vCiLwPvPl4hhSPHAxtylT5tP4UseBuwrn+52lje
MHz71jMPVjeQRnp+2YqfX2fyCqXhkx94R5+7zJ4jmIorRoD/9FcuFAPFuBT89LDB
tLldTeCMtF7+OQbXTl/0R4Pjpw1vJsediwD+6RdIj5uTDJf/quH8x+69sVGgzFuy
vFC/QS96hZZWGFr3mYM5zAXh718adOUz5L5pK0Ce1aTW55OzxHwwqUsxd1geLQa4
aFzJ4b/KzCMxtFugxPRMuO04ZFeqdJvhsnPv6TH/rl/QVO9pLDv96wVkhRbtozDF
AxDrHDc6ILtW9eV1CdepSJc5Kcmo4My4sozI8ww2sdypmg0FJMwiKM03THjpuaOs
aYKdhbNp0FPQSE79Fz6a/Lki4bvUqGftyYFP7S8pO8h8n932l7nlk41HqNw68ptp
hhmlzrPiTiTUe3sNt9ZOQE2VlHZVNcmogGge9zMDjyCXZjFn2R4KLLPR4q3J/n/X
MjdyD3chZyabR8cEVKgQ+p4A75mje9ClfqFYiShMNxQoAvLZkl6Fnt6R6aIWBpiO
cfM68pRWRC9vNmQI4PO5+SdnVbKyvPmKPRXmknxwbj3tdEo/7kuudoL/wn3ZSUlO
XA+ZLXGyN8Dv9ZD/Jb1rkh1d+1YGG40YBTdSfOAhp8U4J7i3tVCdUiu/CJKbscAN
wqsbA9wJqqaL9n4irpPYHbWmL7AW1vaW/f9R6dKLh2VeXCNv4u04BGVzTEtGl5xU
KtC0DNVsXCuOjSgOoMtOD1Ucw+l7u7PS3qzHJSuZRwLOm8fXCLPzkGOHQQex61jE
f7FzPR+ufNrm4t13EYPtApbgrMKgdV6Jq7HULve+sNbIMi3/1HusUG1LUriLRQi5
f8ySOJswVBv0aOQ7q+WwyGxBYB8cns0byh3MVPcsNyZDNzlTgsIRFDnMXtVRC/4o
VNtAtzAm1RvoMahHCWn3WQOg1YXPCrCIKlaCIPFwMPvedxX1KFzQ4r6UT6fn8bZi
SpxyVroEvptHHPjwM8MNPcE+q7Ce6ahZr6SExL2eefXMJvtPcCzkKKRmcLoQZQnI
B1wADD+NWnf/xONHz4Bt+RGIkE8lbXpZRYoTXdcdoMPgd+Lb1Y2GG8gpVyibJ7IY
xCzDY48Tm8GUi9RAqeA9vTKmUpOl934/4HCcncaIWZ7o6fQBPUzh5TvzZa4fsoF8
azbT1qMSuA/pjLYp1yp+QD1Toacmvj0ow/w9IzR8+L9L5cUt/1PB5qxtgs7xNmzL
1Q4gw7KIcl/c30GYNrlwt/b5o+c+L4Hl/LLXQo99f//7zFD+U/j1r8WD5YDdgCpS
HtA7emmQCbXob/PhlJCMaFZ2wUwBc4nzNRnn/2TX2tmeWaAHCqdvkBAV94LxThGD
TePq5vVdEO3gKgQ02AFFhNOZ7n09Cm+Zb6xOn5eldnPwMJ27dBRiPnfh3eUdvUJc
nrHM4RZi+tD/CRieFlCrAdF4iW7dFJ12UoiuqeRGUYpKUVlhPhYp8TS2LWR+WSwa
4G04FxJgtB4IL8vdI9nViBNOLw6ftMYtYLMaxXM+DEwFoQXmkRw4FYm/AsmmD+Xr
IADyUIUl+vYh/6SucBUBPpw6DMXiIwKpINvfNYrUmFRBVJzuwvIaYKL2nxWVxyQv
GGjawao08bNfWDMPTqYM6zNhymc+rUTsAwV7IXXuDtu0k1EzKUkBDaLXkobItKAs
akCg5Rz61SrXXa9pRkDUb1zDmxFFjqhRkisE/bHwMnHFKgn+TbYJM1hOLwd8y2hP
YBVWc0TcNXfF9cLqJ00e+jv8ZzOd7xD/r1Mf9MUljSSC7inZYUEGdIxeHDfk/eC0
zCJOiUr82B8zMDWoeeA1uEz5qWh8wisG8IqGI9pD/BHKpy9PszMJ9TF2nz02JLza
jr57xK0VLM7t90bI2NZzlp0MmyO7ppZNlP4p1vHcW5tPovj35ZVQPEXrSFwZa7RT
W0slJ+1zkOwLUotpYRyJurKTaGXN6LkiPVofYYGyegM6Dew+rOtd8Cz73Em+WyvT
GFva49WEIV2hSvupJMTIZCx/AAjSXywpH6pchehAUtxKx4hpwxwRgPrxpO3EMVgP
FyozU91zNVktld4t4w05wI8f3cSZCgz3HS3QD9CP3zq/iDCBlB+qVSVd0fXrFaRx
EdabcYvuBHeQspBKpdj6RnWcT1U7SeNIdhwYWtli+G03AC1lmRtrViXrh0aOEy3l
QxzNy5fcc7/n1DTOw8tZmIGYucwt+a8meLIEioACuddZFQCb2DzyaOuxSAJ8xc+r
7nnymwSUmxVoopFIYJF6itw6ULlNLjrPVln0QqGq+C1BaYnGAVVbEgz3T6hMu+Yh
ch/HK2IL75wh9L+nF7IJV5mTXVpH5Btz8XgzTf0SXrAxR8++PcRhUrJqdJRkMJo+
1NEJYpPxp3MqjRdHZLuF3jlfuds8m3cUwSKFl0cw8XTc+PBvr5pRV+YfyVfG4bye
ht4FCK5EY+QzplIpaO8Jl++Il8ukW6So9Iq1IyDz8JFOJKQFJjzLuk4pTn6AJ3pK
Nkoism+4bZIvZHI2/g85NJjXomArk2dRh8H4UCqKivjEcbx/04LLwpaLAzTnXeG/
a7EzLMkob4jRihC5AXSNOZaISA7yTTBUk0w+aoEeauO89y0xfwMK7SDkDrzeYoQA
gDGr8pAgjVWnVqWOKjyIptGfSV4lvddSpjeskfnb3Ri7MrGDdsLW9p3bPybW9eSF
AL+2ge4/498eqaoL6caKZHMS7222+zofzs9P6UYTkN/kw0MBmf6lfh4qM/DtTFOe
cj1ZkV12AF8xQY7Zm42MwD0vF9WkZ+R1z+52dLvcEU/VPNlw7IROyTMY3wHz2+B5
m1ObNKpwlWo/rOo6/MFIOP184fXMpIDO1tyCkvytCAJpc3W1Y7/Q0Dg1Elsx0Xby
vZBZw1m/EhHENZpyuCS9Hz0J2r/m6S0iq5O7bCjZyWtEvBIxpKFXTyaaeyc1wlhs
KaY2gs34m59U7b2q6pvx5Mm6PShIRKo/6Fr/gGmiD0UcS4mPKlbuA8e1JeRwj18G
vK8rWZp+KcBhpEKt86e03YIRoV9n+oMmDU079kmn9ciKOyEUDUmaCiFYk/KTuC0p
h+HmN2afLRVsGE5pWAYPTwxto/kGhAQ8HJMm1xefsv/bF1ponsky2ULwWRPooSMA
GhZAYM4UTnML4EhIZNw3PFDlaP9JnXZ4KL1fFQ4oSn2dzpUZkwuFkOpGR/RUD/Cz
AC+2+fiHDxta/tm2brNTYqqOgVopVPRfgZ3MPoFKO2qpBvfTZ5+Awa+3IPVMcB+f
ReZBZBC6hmqn955rVsvFmyasSFtcA7py/Kv+RoKHq0Z9t8gSNHh1jzWEkqn6vzTO
Gimro/6qo93f0S0sCEjPKmEf2eP2G94DxwUEHx7nF8sMch8jg+GTQCwGC4Mt0U7h
DtyZ0x3cMVMLGQiA/hEeCB7mMoo5vzgK3wk4CKh5tzv272wjeVyYQOnYuAnxNJlL
GWA9QghOnf+WoscmeKSeoUY5suy2TeiWJf84bk5Po8Fba7bb5KTtJQqkUTqyA6JO
ZIYZkC3ayRuPehoy9FEs6muIZRWZqYkm/4gsl0eZj3BIqwxNF0sWeh4y335LH5sB
N77e6eyho0QkTc4XRRxPHUeKRTWhcHxHc1P1l2NtGPrRJYPJ1ArLtbX5PjFX5r46
ydZLcn+YEFRjF2mqbnHb0a+fOna+/xZX63mlDGypMJDWi5bHcPQtSZoyQtCulwYl
LTOD++Ybnp/Lu2bEz1RM9BhYwTz12CHQYiVqSo6rhZSZ+42H61JNnKGhCcZBPBNl
+LBNkLBx9IPxTWJH2jXvADToVOdACDgVD2A46WFVaBVGKiX3kXR0dCjVJazgNrd6
KRlc66hdselmg2eR1eEivGqvnTQ/RV4fK3jSyZEOBCRDVSctky5jCSFZpP7Pdbie
yXibdnZ9tHWnd9N08WD6JKFTEoerMI491va3f4nsi46PgY+XA1SptLf15MKHKZpm
LuzidXJ1QcoMx4RCXX2JiWk9LazYZ4TpuyZUF0+cnx1UwpNVXG0G/BYuFN5jqIex
hyMZVID5sGjoUH/UMISiIRFcFoUloXlhuSj7j7gnOSxz5I/Of7E6YGXf7hW0zoh0
0YirJZaZa5HFTFTDH1vkRTqaijQo4SmMO55VtGmDnzmjGGENbZoqT1sbWAWMl7Ut
CBzC3JsCgU6dD23Xt1H1lYifCRrb4+S1XoNnp5E+TyJREOkPYxffEhX5VzNS/9lr
lfm2PzCAkFZoNJxfIVgMOie+iswL5B1bg7UFJjCCkY3+ecMGSq2c0wOdlOgNpNUx
Zi7w9H1bKP4y34s3q3bX5AAb+Ag2bYC/zIs5dkSB4Nb2ckR4tPziQP2FTCxkiI86
EeWxMqpnwss5QxUKXL/iN8O8Q4Bd0DtAMcFfAwA+E0ZfLf3+SZqxFsOs+CutM0BH
wi8JTWy29vrqrDO6kFtsORjaYPkNeulwVvtN5cL8xQ6OmUcNMYuJgQtWdzq/DGpo
0GfFJ9iAMdXZz6repnSbdHsxWmfuXYGxbR/cYzF+pGpjOgTUDBqHbNqT+v+HPV/C
gSPfIN8piKJ9cirGHids5Jz75YLAbdJqkINHun7DJwXNybfRQjrma1j6o4spSJP0
7wQYZkL6K84sbIMPTL2hqnhqvZl9YAxZE6xlmsSCBLXDNPCY6C49/dUQGgIOymz6
fngQ/VUDHKltVwBA8axEwGwyCtjo1ieCWiPZg61IeakOK1o4ly1ER3s766XUstY4
wcgrfvG6f9T3Yvs/ZKKEQ4Cu60BSPVPnuZYzS8TTiOnIWQUF+cemndCPZE5lT2nR
WK7CZrNxktjelA314csEOSUiG5jKFjaKkPEdoL7bVaqsKB/7H4hYInRV+h5W+DMH
vZOeHFMKLQICBHJ7Wq0fQQ5fRuF0s5YOQker/Oh/tgjg/W1a6IU/WWmauhh8Y0pw
gZaYP7bWaTy2hwRiVmZkr1FIb6Bl+rAaVSCxpk6d/L07N6N4Ts+zcrT4A0z/B53f
y9J6YK337/YRqFLav2WGL3ai8hIlOTl3hnZ7BXWdLcp3UydAxxYsDA3sLk1jh9zp
YdkPnKLuFj0mt446qGoGU11tMuBQkV4nLXKZhceTj7yWXFvPiG0jeoZp0kRK83Mx
dg7tYYRc/XyL9HXqTddyujZMGp7IEzWCQ78eZERUeKcqryHoakV1motGeCmIDY2y
eS77C00D8IstFS7zfMU7Lu7py83jOgf8nmR653hSLCxA6I6irk1gcfeqfW258lJG
bimiIa5Zph0FYRAJiQQfyKJ4W0pZoMYgQb5Q2K7Cf4TMxw2IdFeJm8XvZLPu20j4
y4rBoiVsKEEOXIBw1KnelPU+DMswxITCyZ3H+Ul53LRqsDcWVuvOctxw9tPQjZX3
DhQcyhFvn6DlJRoA9QprorgaDYe6ezFVbZR5ZaPsfwnKQppYyf9fIYUX0YkyRKMk
pYg+pQvnvRvlxtGRHIm1THdCnLdjAIGp7UZvRQGcqbf07MtjpognmROdHWc+f6Yb
N+bVPebZZMXs7AiPulWKD5Hqyh3aT/A/XcOfmHrYEVvi9uP9FVHR0rB2NO+06Qbc
wfarSMvjEFlCiNdnkZFDszLVBYpHaP72Do+UiIjverftyR2i17D9jKHqb7ZIOw42
rGO2w+CYB8TE2+x5se+EV3JTjMo1jZjjuqUNe4mezXa8zMbfYM8DY4Ivaz8pGkbZ
dO0sav3lOjE8YidHqZ+afRo+t79mNA3gUpY4SCu8cDJsW9fKf8E7fE7OTVfecUkC
wbpH63BzHSBC7beLiDx8e2WL1q7YI+IBb2B30Uu4L9K0xdCvU8vWLVmuGzlZrsxj
j0ZS8iczRtY7XfDHc9qeCdrjvz0v/f8AiK+7I2qNxq1h/ox+qDLDb/oLdiML0kaX
/btZw6AqJNi04dfowIJBsUHSvsbx3A9qnKVvpfpJfzpNE0Y/j6shpz2eeSy6Vgn7
IOrqtqkjUwJU9vKh1VmKib3L4IkSnYByUUkfeuvR3K/2mPwFKT4J/bkJlFUepki2
m1r+J5qHw8eZh8UvVpUVwiEVuTryFet7zl/WriEjmlP0aZrt79yb9RZKP74gdgiN
cbKNJkCJVeIA4+53V/ec3aFFOpeBAh/zqg4ZsVSVfuIKQoIIUzBstXXuPwlSbirx
i6l/scwgQ+yz9+sI6lJCWdiRZWjswizR//JB3neFAnzLTKzscxWcW7vNIkjYDOwM
+lxwAEJ5311xd9kt+HbOQYxsGUPlGYPmdHWRTi4tcVjW+3iYL9J/AVe9maknYPgV
4f5Kxuu9Q2lNnQedhD81xyCSxGGLhPYN3Za3SO7Pv+qZPUlH7Hn7BcTUmVa1KdpE
C7GPEREmSIE9+YlzfmMF95KmctumD677KI28PQMihqIdc6NAfA5hFckZFbtqdc/M
JWHtuf6KbGSN8GfQvGvplDiMi7Jap8tEzmo4l6B+DgzcFYmWtY8419t5iw20moPG
p0fQOw071pV3kI2bRKqAr9266h/UYe8iNlrZ2XS0qsVIZL0o5z1TqOvLa++WbzB+
lAhmQ7FPQPXzAqby2MzgOH5XCAlkhysGL1APFzoxzhHlN6uqO7G2IX4/CnXW2F+H
Bh6/3KXX4CDFaM18Ehh0rpn/l+SUfp/VWZ7Sdrrr9QZIdUc7jn5oOGlpUdedgndp
1ddYNdFWpmiOp4J8SE/6ZIV27DsHVZxQOHDUyEPGhNzSkKuQyXqxgm/A+jf8aaGy
c387Jke7mZAehsiWZ0A1mF2ddk8moeb5oYA8xgkg/KXVmXz5ydVJW6g0HqamPFuq
/FRHwoY0thHog0VuHcdqW0uAuMgSd3VprV3vUXjVC4G+dtArOBk+TaAGMU6NOIBb
8MmuRe4n4hZkkxog9o5UTkF8ac1eiYYikd+iBo4l8Nf/2xOGyWiMmmCVKocvWWf3
Fg3/mhTPlGbbzWYtU+kNYTDIRz522Cm8LqUJyykyEt091XWmfYk0qyugciC4Be0o
+liUnNXs2qu/TEfRL/cxWkvWD5RqBHF1Ys/R3EHGKZ/aef9H16sGGE12LvI+NJm9
duhwMbZcjS8LzKKySFZv6NWiZ0cp6f7o1Gv9KTklG//lBDjcmxEq7ohWX+uw4xa8
NfOHR4MHUOm+fNDfWVba3lNhEct/nFGjqiSbTy+aBRN7Vo8Ygbb8t2f0JFPyEQdE
8/zLxD5umO1JSCni+yuqE7HnKv5OSIzXwBJMykSJTgfegVerD7/NgpXNKDCWQpIi
9YAD+1x05JlSCrLGOLtxd6HHNXlclyrnA7je5rGD4oh8YJwaXqBoMzHNVWounCqg
zmtmY/QzmheAsfFdN8dqVztY+Z7szD2XTbel3L9F6AJ5IJGh7xZs1qGpucbTHtM4
jdCX4tMe3EBGJEMmXjKzJUmSXJB13dS/H1gbVRdpA6l6b95E9k1nR0lxnG3bwCkp
XL6O2pjuBk3MHwkNX7lg+yd4fKWwDDUmK/isIc4ggToP2P+b04JsUAvLfe55OdLr
q3lQzZ9Fmpb6gtqjOztl+oIIN9I5uHhK0pc9DxftCIhoi00DrlCZJRnB2m8tSd0W
Ngxfzz1hLXxpT4aYDi/ZuBgcycfhCi7BZLxLpir0b5aWbZIOW8xa7lYtqexAYTg5
o4YoL+BI7ZQMF0AYEm9hrSxwDQz2xX5fUtdApGVMgn5ShzV/lRE/aR5awxHV0EDO
wEB7D0ij+uW2HZq2irbpVoPtm9uw9pzwUjnvlrRl0QaWLBs1UemOlVMhLpifDAyw
oNrvdbEWdX/MBT7xTh6aSzFFyIjmHPtJq+GB06c3Aw7NvsxK3J09rg6E7MRrKu7/
tbtV2M513JdjI6kGEEukBWKyw1eQAGDooJWLsKPcCQYaHP0mMCy0BchiCwA7MsMj
e5Y6GhJlWc7cjQlwqC5j4dIYm5JXqzaO9bTWKZHRlZQT+WtbRgKlseHoUWwtvu/p
16jxYrRqkhZYx+fKQ2PxIGKhM9qf2bLDbViBeiHKxI80VXf7amv+ak74TDzHm1b+
Fn4ZGS1VNWs5rMflJfALB0j4Ggg94XsIdNlOdCcU9DyQg6ec51oAyRC6KPn6mnCg
Vt58xLuAMdzb1Jxc7HF/qraVSZBRzI057JXQthAHCydAXhv3Zh1oORGLPv6A5egL
d+YzUsCFgvudzmrX/IU4LV/fZnqaUpgXExd2svK7LhFjZc8SINmEbf0nOYuQHpft
rz9ivjwsRSGcJF7Zw5KlhcgxSEojGszcyjoWyXKu/9dgFhAgGLZGnzDSr87xFLzd
FQOfgv2J7VsvQ8zwmYe8bfhIBYS92anFXYbe9r0t285uanRGTMoNse1HxBfddpSj
BKMuf9CK6STe2UDXnnglJ8HtBb1RR12kqxmMYFixCmSbjC70rUJzzNyR0b60ns6y
R731SWYGY4TLo3Kd8/ud7gSwMEvUD1lVroES31C8ROAp3Ds32uAgRojf2UkYwepy
nHgTy/z3JWBKn5GiU4X0/TJp20S/utMP1Mr/VGu4laAwssp8oywJ7dX0T5xdU5JK
kBO2y3vOQh0uQ83zbsyQXkPF5xLZCtCeV0GV0YsEWxh2TkjNBMgds1j/MGkbpNpz
uRUyRLhtYeynb3NUdq2+VQsg7u3boQPvR9uTkdG/V254RqMaNrazDmIxkkOPSeVk
sQluBAAaLAXaKYjAIIZZQNPsRQ3m4MmmhcMU2CEJWGbYPQA8IUvbb5+lm+V0hEbJ
b6KOmjf6rbxk7U7oT6ufOY3cEbLjcZUHqGJbHwCmlCdFpM9RWnDTNY8w3U8RLpMT
rRDS2rzNQzFsRLUs53R6phjC1OrC64DumthPFZ+ugbLnQy1FqaPslhT8UznBKL5N
s2vDMJILxUs24vMZkb/j9v3sgCzJFd87Zk8Iuetc69wgH5fih4al76qw5WKnUn9+
YV8eydXqbO0cEHDX+ajWx2IX06gqnbSWSKFAJVgcx2GbakgVAo02DMNN5q7rCt2+
H/zzDmgW4jCjKqUOrLXMXu7bEiL9/jRnPwb7LFh41err/A1wYT+0ZWcO9v1V6hQl
/1cLFsAiz/TcqTI0okPdxz26He5u94T8McYKmSowDn9C9ZeYXh8WHxKXrV2sCa5p
UuJZms7aofdNDdAssYYL5E2bYor0nBgbTzcuB6DTrNrptc6VOSyIKffuvvz4Yi2p
NOk1D5ST+0yk5GCVwyl5aBSRV3opGqRekDQf7R16gcD80szmpvFV+13JUlnVIwoc
YjV8JA3DcMTMR7/AOXWuyY72a9Ign7MhMTdjNjo1gjmqeXSiteM12zVm5FekuSyZ
34e+bnPB59KOGDZ9ntH3GCXCbAriAFzRui0sX4XlUxhruXks9TchYaDRo92ywaJv
/xzSEX9hIvcIfR7WM9TU2mFt/Ek6mwQS/iFiJA9AAbnL8dm1m1ceaYiW/EZD1tnh
scuHUtu5Hzg1sIOQibnspY77UMDOBCQ0xuUxfBdrpzBx6/n198P6b3HOFA6v+d4m
cpIjA6m9Eaieh2a8q5IzbHop9naJiy98WX0XWYX3UhVn00ryUKMqVn9MU0qDXANc
eK89CRb3hULYviK99lu+YMRlwywis2G3lUUs5kh7JcJTPvstshM8YDz24ev9gu0I
Vxubk2UXIeqd8xCShXL451ZNBZkwoPxdfxPtVqUJ4CaODKQo6fh68INC3zr4m2k9
pGNdC4DaM9DBLrzqFnrHDXyshxPmH4Bmdhdm9IpM0aOaFb46Z8Gzc4R/dsAY1OPi
7AtcXUYHK9dUfXVkow3vL/4SMbMS1cSm7i2zlfSzXrLJZtkv10Iw1MA14m/RZO1U
FWmqpdIaL3eRgCf7awQm+lZ2yxJtGX18uA8SY/iddjMuauZwrNup21IW/RI+S2Mq
t9VixTqU/c61uPy1d/EZvLJKMSZscBj/sKtDY7KyP7Rntos3T/JWOKSoDVbMZUT0
1naOwCjEXEgGysT22YM2SzuCvHB/eRo0HlZ2RAm7bR2YcP8TMKThrzG42j6Y9q6X
OsnBuafWlqrCJTj7zzwNyK+hkxvw0ASoITctAq11djRT/RbcWs7tWcg/OVXCGic6
vtCo8ATc2ZUAZrUn0mY4JgtNfmr16OMkNpIX/tZ5VJhEdv0xtzZzCBg1WAQy8x/I
IqShhtBsJvKBIvu/wq0V+hIhDkE5/o6bdYSyHC2W5Re0MyIB5W8FboPzwiCcrNav
m5tY68spKHycw9gtLaHCnQKi0ieoZSpeOAfvAwESrcmzYGRARL2288YGqadsdBpS
GOp+ojQCO37GjvSgyRJT8E/+b0MdxCPLCbz4eHT2WgzhN8Clv6nKX9MKfjQog4Db
M3eqmdbzYld4EuKgIe+ceeBk0Apvq05S0nHhfG4GEF5NYlF4afFlldizZVyFcmK9
SAW2E9yTK99KAwgzSpCCh0nmdBQn/zpJNh2gdPHMGi4hcSMRxDRBg210RdCL70Jr
hZCXduv/lRaZI9Bm0GJUfCyYpaf6wNs5OgdntPnNpSwHnNZPGj279/qC6mbZa5/t
mNeM+CL/DypBHt5yriQWGtG8jnbIJl7ENDpovx284DYd72zBvOAi13ANkxmlxQRb
AHara1jttckvehSms2S7dPSV2LI+lZHYnz8KCnRRBcxtrfdxlKpwHWOjU5BaexBl
lOMi9Jp8z1ZtUmUANKoxvXpFo/s71aWQ2J2nfvINOqNritSWkJF+mKnRa03ucRQb
QWoJ77IOpfPkgdlPEXi99o8+DTEIrx7Vcmi8mxfekmtHI0zqF9O5WeQ28cylBS7l
RpMP4ju8jf3cB0zgE+MYVsP93K33mZ5zZxJriN3GhuAtAXVS1H1kJP61Mjhr2UCx
GjJjZWnVtbb9fFgcCzwtceTUpRbATrm4VKP83oT/ziKv+D5i1/NnXQO1DLKO45b2
J4SUh+qlYeuPZ64jGx42J03yQ06f6sdVoCdlT7CAx80UZMShfbnnQzdBGXYGEfbF
I5Z67MpXOBaqcMkE9RqxUjANty3PJUsAJ7/1I6lyX/QOLTQO5HduVK8m7a/SKrju
Q5D0lAWwjq8v4sgRY/7p/77F7eA9IkLYhYAXv757SolwgTkg//eaVr8F22zDfMnV
cSGnIcsPhHCH/3AGy7ji+T+/7pSBJFgggZ1FURtbkaztutC4lLp1VDKcKDXy+FjR
UIBS9g6iHOdgzwyaVAjKuDcyZ263dQA8sekh4QeQGAUk1oZ47YFY50Xs3wB+YdDZ
idwW+SJMRHJsV9h+3NOk59+NR3vwugXp0merGVHhk72JvF9swldLZc0WobeTKrvl
D7rynKsExwJ2uinEk9rM0SJ3nqyhpJKgFdR8JAI+VB+fC5JfXUR8+oVF3qLft5J9
K5epVAhL0gYO0EHcjkQo9UWTzcbAhg8pROmsk8AheVNcSkioyH+0nrXpupVh3ihh
kMj8xM1CWwK2ZDWvU4nOw67FPZmuMdnsrFaGJmWkn7sYvDoSP9fwxZmzkpr2k/f5
CrRQzXABeL/RyQy1tvH7yc7IrG7Vq0cRl0dmx2g8dfFabePvC4Dayw4qOayijOLA
CWINy/Z3pS9mA6IqvZRoIfidLCRGJIVz8Zk7EoUPXYqPxmpNYl4XA/fgjon7Qtjl
snkjvFjKFi28krHRRJRO3EAAt+bOSWpjbQIys+rL0/Dck99OTndWZcTsNar8vzot
Zzdb3bfLwHkU4SJXO425tyTYKJhHyWefEhZLGviJfcpXZ7ZQW7Zecyu0h9gvSViW
RR/I6mjYUzfHRbOGGlex/Tk21X9XAY3NyMVI1WogCQRhulanMDVhoGnnL4bjAaja
OLSjmmL2iOUzkKC47Rs3ykhcL9hTmY/7jbeBdJHIcg01pRwKP/BuQq0q6FnKqeKj
qQZZpbpysWiRc6VnlL/RLUMnWQsaC2iIKeeU8pf8YvHFoePwsPtyBMnKqoMDFjy6
G9GLikB8NVm6B2sA87vWvgzyOO6z00PJZGRy6GkLVAN/ubVMLCQ9ezNrW5Qyj1WF
M/uOWC/JFVRijBLBocOJaeu3XT5bXjiqAKKPG1ateaIwZoD5A8KioO8s8X4wmjiO
qH29uF5JU8H4FSZSQS5kEreoVpMqxvSTo4sMFNG/9xnYdj+ul1IhlMNsb0nM4kzw
vifgNuth52lgAWZbcCrFX4zhl9k/v117ZMmD8CPeIst/GZtUXXy0v8PcDaqo8b+Z
/ye5SMXJQB1QhG2E3j68E+c2lmkPfFcr8OsS/awDYo6BlUenjJM71JrJ22CBrb1A
+4p2+C8CK5xkGaJ2xPdYFA==
`protect end_protected