`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 50560 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
Ju3IpcJpVj/VshHyynUPTG7kN5gTlvLnmXIUJKrchuL0/Z6hL7adSW3gqI5E1HeS
ECumD+lVTq25Le0QK27XVhbhwrdkI+NOg3SleKn0ZbnYcw6wTFeZYlHzZsdbHdqB
PcrEqfQQfZ1pQuJWTy7DapaQFulUB3aC1bFGk8G1H2tw8pFb4DJ7m+ZOWEg37r8i
kuKlJHzIaDeR778lii3MlZOM0/PyCKl2PbU/3WKBT6qrt7Ack6m09NMl0sIX/MjO
ewSvO6ZiM6jdiHUJt9T5bXRiB1MoRjxm66B65sTrcd+p+N3rfmxwo56fK+AuMLNw
LbyqrNZd7n9dDhr38vF5IkdyfUS/VeVzuItlFQB2Z+zf5x5NILRhPMf7v8Fa7Xah
kXAxOrEcaoYg8r8+AvP+CHJraVKObm0mbBGmclz7zTLw9riTi02vnaYI/YpvoF8G
JFdx8RFyVGRLn5KsjT72D3Arq/en+0y89rTMOwnLAQn8IJa8aNfjiH9jszVKE+/o
IVe2yuiXwwABjKnQpxolh3hTwaAl5+R3fUHJrv/CNI0iGk7OBFnscbKD1zTuKeKF
0jjavdDw1DFp2unV1W3yqhR4BgyKQdzkwLWhcSvcftA6Q5D6KrS4tGCq5lmKSd8l
QC9pMmJIeywi23dr62QMNz8qf6KeslwSg4whshcKLhMWTTPHpZokIdjSK4Di62V9
GsL/a6Ap6mPj9On6yrhO3GMv2WjZNyHGcKarmlecV7x1QRDHVaeZ9iogy/Ifdck/
j6+DBzAjnSgNDkFttDrg9/zdxfkm6ihptq6qBh4E0tsYwnjZu62/D8pX9qU1YaUy
6bzjj0+2iUCXuSGuX/QrkKzGsP41VbxPQjwwf8cyIC2S1k1cu16wk0dDbTheUVhk
KuXIb+4lyaiHtyHJo7O4AAzJZ4mCqEd6ZZJLkC354V4F7vTP/lx6DufckwRENzLP
9kM13fhzS3ciGVECUECJz3H9fHlGK7lF4SXME0f+nrjpOXsJWieyWzQh+ls5dGP0
6s491xW4s+S4JI+lAiBGL8AuLxYkFoPDQBWPCpconNPRI2xqwOLwE1RX5wYanTND
TluGZPkad3ZiizVN5+fX1RIz2nxvdyonxxluTcLCkGwMw6BpSVYtXaO+9oYXYOD0
/rm2n76m9V2QEot1m7gZI4Nwv1dNFqsrhBRHcUGYWtywXKK4vD3PmyYlPcfWTHt5
JyVN0yCMfen1vN8X9iZDD45oImjweC4eVvYzjFVs37pu++2hXjyfITM3NTzXAfkw
1xOE9vURpgpXdLUw057t/0C7G3oDAdkd6i6F94b38+VGcT5h0ceEcCvszRCzY1ox
ms2z4cjIZU314T+CZDV9RTU4emkJ4XXoh2uZY74o0mr9I/RQ/S9ZziCk3UZXcioG
czPeWmYaFx9yPhb4uYBp7nNh6nprVMXHLl/vKc+x0NDQyt8/Tzv/huAx3gInz2+b
WHcuM5DSYu7FU51SisP5jYINSa2N2iT3i+NVwr7+3mQqnF7SQdgmJoSJEZ4F1whQ
A7kzdXGClj+ay8rtzcPibqxF4IXLOJjF7K8P8wpbRgswqSaFC6D9IEN51zAgngwY
5laZ7JSlmAibpesgDlxgYDUMvmRM9YFkG3cOe7zxBiBG1CKZat4vGCUJerR9AeJX
rUfCYmLwsPepbnF9KlomB93q6inTlJE8cNAXAXtNtHW+LkqptNtd8LSxDwbFnUtS
BrQ39hVAruRZJK03XI+skXs0I4O5fAHr6H7jPNCUy0H5WbqeQk2SDt7xLwiSsI3B
WGz68eQH2tQWUccFuD8ZGQL3O577POi1XvHqcwPZxPceGnaLLC9ydA1avx7kjJh1
+7IwBeiMGhSTg6JHd9etCHVokKj2dKj49dFXwEOU4HdRUStIZYz02NfTi2nwuYlL
Ig6EF/+WtNxZdknpxCPSMpCw2krWtS3+vblbyGKTLtEi/RW8mGP3gMDFYLxEJ1Go
VfosKxoRMofu75l2Tg7oHRKQEMDKz1TP5Nj6FUIv4s8faq3ez7nJMR4E9M+fu3zT
TIf9qigixzyGuVe7DCqHIMfmP2lHJE3KSCaQK99PQ4QkP2E0VHwTroS9PkuHz51u
CdkamsVkdV5AlBkBZnzTRDoFjhohEJkXNzEmQy8MDYo6xmFMqyEOrB54lxYj4apA
pj+x7ODjw9Q6jC6NPZFkFiyjc5Pb8cQ3sitf9waNq0ZOK1FT9V8oZmjvA4KlWFgW
33zvPbkXaL12SPA73/MCNkzrag+IT7aicoNROlkCER3LqE/EcY3coTSIdvIvVvOE
QbFyMl7Jje8Da7jhMju3n4IJRCuanRUhAxmJQCjItZyQrtXym3CBq2PErPkUOK2z
JIzz939LNTJqPcC/uYaQA0uun9sEAhA3nks5Vm0/w15wJ7i7i9C3rH7Amt2g1HBs
zpwidv//WnlZnRtMrsfseh0lcYrA/HhcXVAdxSi3wmkCf1jpUcyIzWXaftCoyjj0
wQjL06QUjNVP5rBjohQloe7CQVTOl2tTAQPAZ4idxMDT2xC5nK4b4MOFR6pR56P6
reeDq4od95hD+ofEROFUlUn9pWfUEJUYCYleaosyMMa4FZO6Anqr7NnWleCkAuPI
pDjOLoafdCop4XswUzACNzyffaIqxAdf2rxAlWXmaeZqFn2t9uY6OmVp/DcTyEe/
wOon3upIkHq440rMtc08XY+g0L0tEnMagl34xs9/o7jjvXvdZPqIiirYWgNl3/rf
cEXtwoWNH6vW5JM4FrilOtzdS90mSJbPpe8y+eyFF8K0RVaCaXFdbzElbSp13BOe
iLwFM1wvAnH/jg4SS+eMMtiR2ByxaMP9896ooCHvTHuqHTuM2xIVa/jLUPSIxamm
vk1KSZbHYBed+UwrQGzlGoetsJ4KBP/jEU7tkj7ikqh5dGlNqNoPTjg+NLQZlJWr
4VZxzUd0gVJecjAMF/4TnXCSzCzJPMJck1s758gI12ZIBSswRV0sCMcdMqXu+sK1
Q6MijgxSv6MJwaugyohb/rwNv2W4BzcEG87eAUs10WyQGUbyhczOZLzJyWrFMk9O
Y1jndIc2dimqix3KItM5Y1+HV36t/kf6sfsecMn3TVXN/Eth4sTpDnK5DiGG/hDR
p7VoBiaR4k7bZGB+5PIZfXFk/4g2c6gk2CBeZis80e7xncjLdpLR8qPRifijimYJ
uaSHSQyt88Q+01DfHVqvY9ctjTOwYeBDm/waPbT/gzK1cLCncZvLw1vF84bJNn4K
JNVJP7L2dWcP+4ps+7K+D6tbj6X7RXgKGa6TSh4m+Bmpelsed+e2aayABQxN08/u
vVBiTDLEZ8LZ/ai62M7s8e1YF92NdsaDphWtVoVKZ6ww2iOw4vrDASRvy/nyjfpq
RCb/1Jr2ZEqRJ0yOShm+14iy4MEUMSKGPpBX1ordge+wdlpa6KByIeI6yeB3t2gQ
z47kjDGgBzNmOvQwrLemhCiUvjwoT0oPZ1Kfsmg4QdxYBR+Vbn6/cC+eqcAvCANU
vK0Z5XdHvuVe9Z8AI5K9LOkErDWSpIcs6NRoIsY5bFLHgkMwuyNCV0Eta94fEJjf
FX8vQX12qf1rnK851HV4y+L3aJz3SrE0s+ltA8l00pokRkULoAb4/tsqxUpXj532
+cm2s45asdkZGIx/CCMzxxnpTCyecIvzlG6bTo9uKMPL+nj4f/NSwAfkXOIpxsbH
xkAtlShfmpynF7GrJWk4+NJdSFEiB3jPpvN22H9UgwmbA+uLLxTGNpCQ4yNb6SY8
AbyX0Dp77G50EYvTnQFyocEjGB2xcuocw1K/GCQGJmKPYYXIScNZDRKEaaNT9Qva
QYsilggogcpt7k4gYIDUGI97qQVhGdInp96GoUt3lXjHP2PuKTTCBQnWv8e+9lCl
tZGyWiobvakycPmXjE8ougJS8Iy6tehD9cFosFITZMzzMVq63DwmQ3cGGKtk7eyh
tEjPJehx+yyUyBaOUiBqTof02s3WJLiSJc68aPNkyw4V54ILiGRAIhgpnVmL7foE
C/Li4QSSI516HAafi9MkVDC4/QVx7TTbCuIC18QxqWWKLwtipVY0k64VcnNtjHA1
0OCh71KCNWpUh6taIK/QiU4YINkfJZlmex6UpOLh5pK3wOG8Xn9WJTwsMDuUxkua
EeswFFLMdC1K8q2Dcj4tmHvnuDl8/6S2kSp+qwX2XqMPWpxsr4PHxcO356bfq7uv
l9gjiP6qQ57sT6Di4pFz65hJjBMXUP6PSY7OEQs6AmbV1QiMRGb68Vh9Rf+7Mpu3
mk43ZoKolDwcrM0+PquIa6H17XIe+HTTKaAxXUpYQD3FLf1bDu5zy+yNuJsVgmQZ
dbEVfCKAW9gBEd3CmN7MX3EuUazyxBloGmC+bQ7mu2SUGeLV+9457lTUnKLRlLXy
hJJgr5YwirLjWYE6prTszr65BRPsV6W+hbLQGSXKcZ8BHa3p6N66yY8CBO0czYP+
qGH1oLVSzfVX52udttafBfOxr8MbHI3VidIEA8KmWBehfeEz0qx9qlSjYoEtcDWc
+ILIFmN5qm2ofZW43+fLb8Qc+o5fpwL8PJqU1zkXPrANB1lGAxNzV+HGbaYkMy/z
c0KOEVR0yQ389oPpvJfBWE1joxNdHxEBgulZ+giRsd/48favcjjjJWgQuFTyVKXs
AAhB1Zup2uO06S19nc0WHlSPhSc1I6yEP8PC2guM3sFoLiSBNumf2U8Spogm2A3o
iEMPpxeIOxQD5ytjYfYEFkR2AO9UBDSewzgFeeAwqrn9hxCvpOdjgdQfmEQMV1T2
jz16FKsd7WtZg3OBtk1vNDrNEP3AF6sr2Ce+Xl+O1WH2UeYjySra3JKKDAodpJNG
sVtATomoSjrcA6ZKEQM6qcxA0L7HaS7RfRWws43uOh0MMmKFwRi7iydYuEXnBEZk
/9q4hcTKTdAazoEfrACRPj6QwjdIjyilDiqGULhDOaXoDb2TbNDT+cUR6/IzzuZ5
hs5e0B6mojI4EY52rTMacraUGmlg/mpxuBkzLokLqiGdlV692Oe5NHUjmSsJwWo3
Z4tBZK/1Sc75VmWpt+BQUd0xPjfGDizJu287ub3QkrkdkYptRXHnaG0QeyNztf3G
dVwvkAdlQwY6PUa4xSURkHmvKWB0AVjpDCYNpIRCEMDkX2U7DGguZQXiIMvKn8zs
P1wUrAY+EGGDiDrBMYlyJyn57EgHcghrttnUR09dSaAhDZjDdj6dzpKcoHA1JHJN
8vfic3tfxxAmx2MPbqCpa2eHCMrBz1cvAdHBWpzQV6hxz6kABskN5X6X3ktg+sHy
9R+UwvZuZiT7ExWWUulvUPjNf1uVVBbPwkHpjK/lAtxewSsJ68sXwgZtXksOTvW3
guSNw5EdFEjJ6EUxhf1qshMixFqVa+PnAMPVCxuV+TIEiYnnuktlfeXoX4pFiWP+
MJ/Tj/uCtigHjEPvQM1IMuMkwXZ1Ng61juW+dEeJkwC2B4I6vtBmgZGEQAsaqqhv
3eVRwV6gXOTPAlO69wQf4bOp42fDkkLLVDIhC2oxoOJdb7T/b/uelEiSIezyMI+N
QGlwf5Stlpcmp5ScImNBqnB8lCpk9EJUqziTrFnztyjCguTWskFvI+g+cvPetHf/
VY14/wgS2DHO/8DHot+Ewor1GUP4Z75qbcP99RXXAoVXZYd82J0ebbSoTfOjovQr
s4U1IYE2aB9g5DsHVWbwUxeNUztu3XreREZwcVn0jCvEC2RAhXJdl2aKGfaxkeX8
NBRlhDfzK1fLFh3Ht421ELmGoJ/Tz8h1JIcywaC1NtCsttYj9u9jwCiJyFp2LoIV
63fPnj+NaTxkP66agHbbVNqWg1kZhI5r2NG4QoWse4FHY5en0N6aR7ABAVjZ4h6i
PAoy+pFUhCL6vpDRcDTlU6XlBYmbIHN7B7taoA1WAGIuUDtb5LDAF1UxiB7clLqM
Rp+B5oRa6fOtpFw7TSpAG59iwUKH3aZnP2oqeiI3Iv7zZigaWFw3EZ/QFMLTosp4
itQBq+PxCsAH1SZTaBbNUmRa7tNQef/V9s7XbMum0z8UnVQ5mo0RKbj5CYCcJGr8
V/mx3N/p89sMDFRDqVGD8MFhm88TS3uCit5q9orJFxfDIngsp2wxRRSVETG2AjJI
pEsydFSPkJ860B4da22JaOFqIH9DkCi9CqMPrpoxLCCFU71aYxYhLBtAVj0OIPHE
H+7Tvahmt91hq5NcyWLW41RHo8k06mCcqcWnWSKlQUzonz8Uxox59UkpCf2WvJJj
0IXpqyQmBkhKI9eVXzbGwMQyom6nyshFQJH20raS5aDynDOky3IcUvTkNiIM/gJ8
a8pvj6Ki1l+ogVHQpP6BHYdARQDUdDrfARWOmXr3niOeJqZuDAJ1049Z6RVu2DWg
w73+oB/qR574zo0/CK7vqHrQUq+JklfzgGrku+qVcmOEhuwjr9nZc1lFZpEGF3Rg
cuYrbEd8g5P8WZf3Ou7kDdM2n5POLw38QrZkk85cFqWelF62RIJYFXUYXsIKQ3QW
FNRDb3rs6BlXaNMpKLlEiTMmj1caluEd8GfpTnQsRTBmgctb5V3RSl4FDY6ATo2n
RkwgWLt2tSyp15Ub1vd99+efaaHLY9x8xyeV0u3pYg/qezxyTYRQg5iVtHMIQJxc
Mkc1GD8Fh5WU+2opMGCGD36pstsq/vUEYnNwtaNwIZ044XdVqSJlGrlpNs+o+b1n
WPMrpGKtHy3L0jde4Vuuae5PO26KMv/oNykRxLaRh8wqlqHXR+FP+jctmUSIuedU
DG0U3lsKDzMipg1hmybcvpfWRSXN18igXTtxvqd3BThvSEvyccMPasYXYTt+jq2G
sJZpyfrvE3XP5zhzESe1RcwvOHq5oiK16ZTsf7JMW/dbWkm53rwlPszMWgRemNNl
Okim+oUlMP0c5fIhMNHeAve10fmXrse43cfuEIDx4uDNT3G+oSuJn7Bfn320vQww
k3jRgkO7G4/8Ik9SipgdSFgICRSArIRBBqglPnG8TkJzXpmLBjsxgVZClj1NhijY
lMEO0v7e8aPqSqrtlIzaoeoZLfV15di49+5/1rpDs4o87QTeVpatmEXJVV9lp3WO
UyBpU6oQ5Qn/EzfDcOhX0xZEnWJNC0w0n7EsErLDTUt3x0lKDDMAZHdBJ1gM84xR
sY7hp8hUo7zvlwPBDPabaphY2HRv4Wdowq9rIWYuXrrFWHa8ir89ozA4/PwkVFWM
EB+mDIEFncNSN0FNBZ2pe7u/b8R6cKbo4GpNYoo+O6WvhDLSXLtzEPneGE7OVksh
wbtBtNYXLZCybkzf/YRSjxIXnfwGO8RlsM+AJ+lwVp0H/W+HGWjPC3MYc3LLKCd0
LnBmxhQezAZw92+68pTg/pdiPvwG3KENtOCy/lJWZRoL03diWRWI3odNNhOmxA4Y
NZcTOoHiXV/IYxp5czX0Uy8QKVdrOlD3frAAEGMLRLVf+QK4v4BvFZFRKmaf1loQ
x4yORx/hBlFAgkZdXeKOYDCCqbA8p6mkuVutVKGfrw6TSkRf2BDfT8HENYdEo8PL
/1+1URbwjQB4tvikNhFQCE6lDfWZVY0yfSvTgEzHC/2+AZ6pbTHIrR50rZrl0gQT
UyMOoDP95oRvnRh5gdRRH+vnAaI3jB2TwZmK1Qc6OZyikp6qlwFQj2JEWncIrVV2
aHdRFDfY0ZoC3ahGohuCX6pas5Ba4fStdKIYqT1ObhlVG5EaObfcQPmEWMFKHsqy
4/3Wj6FZXWhDIDDp4sb44qBQcE2O17Rt+Ks/lkFSWDLQ19AXc02MdcOvfM+YzRAN
DaRzbMsWsQGR2dKG3C0W0FLqfa5avCPmzElrQe6SX0wS2/9p0Y29xXCQ1z7Rrbt4
7U9QXOu95BQH2M+vGIRbaSBFqQ6gXkATYPNsNBSjs5vamlmcNKeIG7AEYPr9MFbU
rbLysVJ+iRjkNrB+3NNwP19RqvEtu5JYp43E4aqKYcrcNkDXqhnGIt66BH2VJkRZ
Hx7ed12Gp/i3yl2InfCg2qN0jl9TRSEO5xYdwxm8Yp5iBwBCxThXX0M+pLm9HUm8
hM4RfJCD1H7H4Wph0lE9SGStOvwC9wy6a5e3P8Ikya9ADdmkC3fDUeEzNzfqs+qw
ko6h2k+NonPy3ROIN4L4eaO9CHdlAvjnAAq6otujiffPgkotCEFn0fIj7rpok3ER
j4UARYbytPnsKkTH4ZqkwR+UJihkO8G6PrXthzIB2R014ZCcVIgaNuyuPXjbhc1x
SQn0pFg+Vegx1P8zrBVeiKB1nAS1CV50qHk3yUns535e4K6dnxXQ+Q+vXK7lXb0u
Jm8LqYclVMDoVVxk2B5UmnOefCl8JLv9MfZgTIXVw7m/zdbLHk25YTMZQOoKqTAT
R1R2Kx2WD0+jEvNEOSiFdXZ151y5vvxL+B9iaGBVeWNkWqN0fb7C6WMvDzF8uoA4
fKJ5PF3p2uVhqmDDjal+9RPyBeP9b6Qwblp3/t85jusdy5HXedL2+IrO7Nan1FUA
8prCWcXi3kQ7q2gLrhQV32b5IJltq7/BlZaY5RftSchrdz/RFXAZETzzY6ZSDL9p
jzvriJGREtu78e7Jv1hy8/jtI6Q4iZzzTciqF+p2WcB7nJxOT6F4Ai+bY5DacC3x
kkaOWQT3GmK6BXJCIUg1/CDS/1kfE4OyJlxvOAsns+ahG+Vnc2xwY5UGmlc+PefL
EfKQRo8UWUASXehRipV39WjO2bgIDrOHbguAQK7TE7WBnYHYIAYZKp0O1CVbHD8S
FeNxbfUsMPta41KTvnjSRPEKzOeF1J2tiPV4vaiP8BxEvz1hIEIK2qyopzz9ii9v
/6OTq6XKXuu+5kqQ5FmSKBNf/gCT7eydTpJFueu7htTP+b6UBTk6xpelGzbTp5PE
J7AEW6yfIhqOZBuZeA3bAJHZFh92/l/KPmQsMNTCRDnU7J3nSSKUKnx2A0A7U3V2
9Hi79Lg+srjHWn8A69pfyXUNsXis7lDwVjRiETosoEg681gk3CaeTuxeghpE1+1q
FqymrDwUy5LlGUGs88H3hAxclLWM/ga/hpbGmBNpAjEmwmu8vTDqS0PZLJR6OJ6Y
46G5z4MTdTZ3wzGUHs/9noLlqzem+B+sBix7SCFdqsCCSNAt489rIsC8hbZ6xwiI
WyKOJCPi3qzefNsaSc3x43rKEUIt8+mn9XpCFpv8NLn7jdNGNDbJysOI/48ymfUv
8gQYmNpyDylLTIm3jhRyOwLw5hzOgZrqKhw33+QRrTGp8bXOwyKjF+JuxV53JyUs
MMt20Z6MuZLd8Ju60VYea0Pn6WBPixSTankhUDoDY4GdrMI9fMuDX0Hm7iJgzYS8
2ed0/vdM6w9XXTcxxDjiNI8EUMdZ00mrGWV+Xuym7YSZ2+96Cg4PaDLccFo7NtcU
mO9oFr0deFXYchqSGPDsj8SYcbLtyaL2qrmfoE4Cf8HcqxZF1aQ1IDtCrzLtcDwG
EOGCfyTBxHENpjUtrGI1QbFu8xeoE23I7zDFmEe9Z7PVvnKxTXVZFZychGYevXY2
4AKnQkJyqP6Y0QkxGsn68tEhmQIZAF8B5PkkGa4CyujUYC04KsRX8Cp9Fgs7azmd
gkaRVeHwbryRdQG//Sqm9JJvDhNBiSnSwt7MDJyTJZuuColeAuwhS0Vy42vLezo2
EsRK9NDpBSnr5kgbzzmyYzm3RbbBMKzDSAmV8kDaVLeDy+XUeCOR5UcEFQ4UpiGc
9jVEH4ZcT/HPBc8Mu1HZB8ic2zHXjOnNp8rVLHsa+ZQe2c1280T/KwCQGryFHrAI
F+iox9hw43ursmz+KTI21NsQMRZ3L2JM0Imq59z1yNAi9gRlheUSbpK+gz7HBoNq
nYToKJ0IhTW5mKV/BPtIyqqueI4BR4vDhNjW3B6sPWtDyyPptbBEZvDUHbJUQNZx
YdCBNblOAdWsN3nCKVjlMLw5WoJqgoNX+uun82S9bVvF67PONS89DR9SG+pweDqv
w91S9RHM6D/7YGmsiN41VT29N+8ajX9UmBGNHnkUP3zQiCLnq5GbfF+zCOcHX8DW
6/+QWpxAaok1Y1RVXSxrQ1S2ykKf+T+wiZA7Pr66EfdmbW7aDCYEFcOtsHSnv4zF
fNPEtuo7qch8dvkKsv1MaJaiBgzRd0I70OKks53Ik3Uwl3J9BPCbXxu2LSBak8TN
R4+l54TdjqQn8Kuz8GxZOpr2CVWqTjipWzxmuwFLISuv9vc9raTIfrCmk1MuAS4z
ShpfL7d4Y0tkLu8IJBhplWkby9cHPboTNZ+N3mZQjSJgh5KKhqytkJK0LKwOw3NR
vHJ4yx9cpqdJXAiE0fNBTgFs30jf6qOENMUEIfoGqTKVevOIPAlj1S3xNTJn4K7c
OL23pFwiKrraRmpWTHksLEa1TH1tVF5w9vZ8R3n7cYuGdVYcifOrMP/lbn3DvlxW
n/tKXDsPgIW9qywXse/Fp/dGfr0/ns49BKPTiYjhYlaSOBljG+j47HVM/6J3lbAd
LOxH0Lrq1hX7JReTDp5ccdcCN0oFmPs4SoYLdelbHZnCpuTkTdti6qtMS4Xu7RH+
PZ5G/P+IrjGTzLfP2e6O0chgMgQCV9uujPAOH6esbRkxQfs9UUbeY5wsP4L5TFUa
UDVjYdVlnBAH/01Ma3BoIZ9VvYY4aeC6i08h0Q6ysa1JbzxtI7Z4kGpLvorJbHOI
2J4HTK/hUsFSFZvvANBV+nWobv92FCIbYiV8+SVrwVmfr1Mk85meFYpSFIavBggw
uxDkkbi+epQELroej3VyCnQdO2cQlL80GK6BBEgQ42wikmtAbPrLfloQrPwR+GmL
rUy31bV8B7vpwZxFela94VtKs2MBF/eYe9tJeyTStuHWwm/jChM6dhr747ZLZ+8H
XQwNe/9rG6SPHwz2BlLCLP22zSWLmHdE67WVvjShUHNfXh4XuOkkLRJGqDVJO1wq
z8o5QKwjTY6mwKop/6CROzHFwti4z8AGln1CCeMD8BDTaEuo9palgg4b1z/ZfbpV
uHoy4gR+UZErNUC1GWf6GxKWj7M4IYVzNTJZ/M2Fsr4EoabkeFIoG/Peo6EoENwk
waVbsjgKMLH3zY+T21NPzWPtucbavqsw8m1SkjYg9VY4pl7kmu5yS/neUGol49Yx
IOQTEhbr85YkVsXlpnHEUQziEuRPGBg9SjNLn+ZFCGmleqp8KsAueyU51hfnMdl9
cstyfd9WFBZiQkybFCFMXbrq69dVSAC/GjfqRAN+/QJ7X1vJTGkISYZgoTczp8L9
56MPIZnzNHvCyvuPbqIGAc47O5P7HW3vXwOIlXVnACk/OfYOuU+N4aRkOE4qPHIn
PXdZ1PrS9s50h2W6BFHGmBM385mjbECojhXaxQ83nluTF5qfdDs76XnQw/PEIJGj
z19f4HemQBjA999iwIgxVIXSDQsN8EiFsUajPnesYAbkkWmK8/LiEkYCIfUmxQ0E
27ddCT8qIZYHC9de8qYxIP9KxmQCjRB+q0TV52EVp7FoDr88vvBfu7GRITDXclkH
ZPt55JkdLffL9m9RbTP2tO4KD1bBkUliEBjB4rIFMYAoZQQSVOFkG80hyzA59MWB
wlPzj1HE4kNHK17TEQjISi+MaEGvStvsZ5gCHd1GwOb5LCvbfftDQifgz7eqqzdM
0h68l6NgeBVEO5TaOzIZjrwnbrn+Pap9dCcUhmI4C0GvUBMQjKpIrSitO6J21Blr
3RElDuo2nDX8BSOrM6W2aok6xINJW4YMchF/Yv6aY0RaBZKfHV017gVGkKzj70B8
rrrXG8wD6AEhZDzf+hb2W5FoDHI1tGuqYjQHQUmtHK//kieFB8CZGqgTh6/G1WHC
tJsS7/spJXqLTgd5yaEowibMeQ4Cmh92AD080jRImpjoOY+8zBgUa5d6whRC7kHx
illadvjYXXQkpFdwxfeQD7j1bJONhmtAbYuORwNwh9OCd5gdxYEnXQDpu/h6Pf3x
UbUuQS9o7UJSkzx5akgCbwUMYns2sKZTOaDqnwIvAQolKtAPZwLITweXV7+z2dmd
xkhGbDvCM2dQHwc0d4+jWFSsSAwp6HKQe8D5QAOIlsehzPCcndqZWAKBaVxkQJM+
CrW6Pf62BnTfjOTgbkRhMFFQycI8Ur96Q/3toXMq4Brw3M1ULJ7KVNdqf2z8xu3A
UKtv37oGnNDHhas9AkNKg72u3HAHkq79OmkLfwN23SYbbePO+3T3mKPrLBDlV5Kz
RjPSqU7uL5fqSuKVj3xTk6oLKSnKjdVy99czAeT9B21vNkTSH0JYrYva4EtUFcfa
E+X87yJ3HbkBuywMCCtCaQJW17X0J0OhHrb8vd5CE0j0GAfRqmkv0igmXkwDYPEN
URhSttgkePy6SvQxSsV0tRNJgawM/rl8oQoxjdpq5eLlKN59k7fdsEfWuRb3REKV
EIx+mpBuINjlKxXHIO2T5DBqJNIlw0+v3OfD80KK2pJlY7z6Nt2nPVVFwSF0EOFZ
JZ6t5TrzZqhMo8S8AzSDwOaRtYURmrTSa9/2W/HTBhpS/9V4TEsh6sMZ19xYM3eB
KNwm9EfGjyKiEpBplnnFrCNZj+CUOjgSh6QgpbmEqDtfFdMU0IBFZSv5En1FeVWP
+id4Yvaun0ldMpnWBgqVwaOSaXJ0c/aULZoyzTulQt1HZFdeBERldg0X8vh/gv9J
qj1xZfN5ElGHx/Lz682CsHJ13NMz8V9u6QvGJmf6HryluaS4lHYhVj3SgROf9nO3
KIr1dygFbob6+pW81dCGlK8f4agMKQFXkNkhLeBT/NmlExHWepOkd+eQsyHXxSOE
1Sz9oE927Bw+GpOq9fgohQaqlkq+Li72lH0aEHhGxD8J9gy0OXs1NFIRy008IfMc
VzD6eCXYGxwweLFqeESs1EpnDBPZabinigFGC/WPL6rLGA4SOblPXHNI9Wf2T1dH
SrebzdpUlBa4WjXrU+AFij40Qdzu4icJV/uLa9T7s3VFvC+kt9po8EpvkMvmxOY8
7IzgbKIuzMV1ix6iZ91EtvwKTKsyb1S5HfnbhKrkJKStoAsv/SQrKjq9bsl+3H+7
Hk/rzoTrLAjEYdKfPXKpxGEPNTwWRAkK9J+0WkLAL8CJT702SqRwHudwp9OKF8t2
SbVxaYNILeydynU3q+t9W/4LgFtvBrZ7qhzscrLRd+LLG+g7qgrzDPwWhEoiug12
IS0v7jzR8KlBAqQRZqwcOtWuRZOcgOgR7iJNv1ztG7TMba6YHXazCB6H50NvnDDI
nnTQgsZnFs6TWJE4AHVWmHq4BBJIBk6HBpsaHYbL6J14Hm/zbP3SpYpu3yn0OHSs
fvxeH9STGOpwNsjWuQ5xVMbOjXT4xez8rS0gGjLN8QOMeEmwuHhZWNXy5de2NGVk
/dzukhrkObYzBdNObGNsVeOCnvkyHd2v8CLMnrnXPzJkyhpoojJ4a6WNneSdWGL/
bokML1NuLywGCpJJ0VTJCwre7tt6icPqZnjYY6UlxAH+hjqtufAjl0ABYSmzBX4R
JXUggB645SGLna9g/6tNLFr+KfyJ4h8wjetaNixCYr4gYlY6uk/NQ3AvoCnnEaS+
ezfWLXcOlaT1DCtOzPpO0jTMgmuraZeIvwHlYr45GG1QtGWZMKWGu58sflIbAs8V
/wTMGQi5wOZcAag1N1RT2BSg3xOLPBusYr3In160YFQAdhoWPHk6BXwQ95uShweg
ryeP1Zg3RItUBpbyye/WxoEYtSVEKEFsakkdwrkqJrIv0xZCnkQp/CYYWXpf47r0
2ypOKdgKEiYoV6NybedULwREHuJ3G/oov5tVJVsqZQrMCHg8Nt4lvFlrkFTryCn8
xjX1Mr/fSwu6VUrlqQlQxnz2fkQF0oO+877gYJ61bdcdHY2qpj/Aq2JqSGumT1uI
ZaGspPVNYRpwWSHaRQ9W/VB27kc+kWnExuklx0/x+ROrtjt1QFirS6ecxFY2GK5i
5jXc8c+1v2Mq7HVa03sSqsDTTwex4jwE8R/oic8dTrigbVjRCBCq8Tvn0iy7CSFB
7WPxvSnT1LLm2ef6FWHh4TX8eqHzz7mBtG1DPTvSJVC7Fg3m48ZrxUBAzoPzD2+r
nWgGOLkj76Tv9Hcf+ttjgcE3ceJ7TWY8kVGJnTS5/FUK7ny0Gy9exUnauS4J9AYk
plIDxgu9F42vPfmYjEDKkBnQo5Dh4AN/iswxlf+05y01AiMa74pVfi3vf9TgdH3b
UzMy5NSf3JM4IZ76fWJkdsD6cqRDKycAwMMzCuVCVHWs7J1q5vG8pdNZ20Rymc/s
zMHOBRGMo5PIdUctMqPDsWrH4FriobZCwvf5qjcLfv8fM1QjiSdf2e9qWM3xgwzu
8T6Jh1x7MUI9x5WyU+ZX2TK2D0Tvom7Ux/L+MH+a1Y2A0mHJSE/lulXTcJGdb6vW
+2q9pL/PK7KiQOngEIxXQeeKD+PsNQ+tXfWDkji15Nj0k81hRVCOkIKA1sHb9N8r
6JFNWtMdH51e5ZdDRFO5AycMFPnFlOHKJ2fjTLy2FNfrMSg9ZFTFKLIzbRwyxKSw
kilBIWVliQ45DHhWYvWm37joLYVdYOdbGTe9jRDd8BnvnCuLT8q1ecaAz0CqGaWM
XOxAuhV22t4AgSaDMYqMP6dMa6yYWsgSobYOY+yZ4qFWYbzos54xyx3OyGm4w12j
ErKZOFUrhhZHlEQ4FWs8x89dPCRsNfTftPCHdwXrTNomMjLY8+JZ8JtA6XyyqQKh
lFRHPbsSfRJlDiYUVQesYDSVLGxiWolkUtg6R/WsMvJlZXznPR3722XzDHaaGMzi
x2BWYJJ7XGRdn/h2bnL/B5miyEpTavfw6/gmCC8EiVovsUtv/zczEjyAkn9X+m1q
WBQIulaW7IkpcQlKuKUU5wt3g9yHvu5hQiCaQ4rbydZH/wsPop1k/OGna5nQmdmJ
m52teZdgQJPubPx9W3kzSAmwjsh9dSrJ6YsVxDzw0ZRx7B87gSvO6vkeKi1k4TJv
x5GDT7OfLaKM+K5qTjP1KuDVgBmOdhQZG824do/Pywt+qQyvrWlochiqTozUkqsa
r2XOIJj5m1yjL0PgF3Igo8Bzgo7ASJhTCTgcOyPGOY7K4yncYikrYYlOQjEn4gbv
7oM14kZ7FNWqQYpwteop7hLYHC6PpHmceoDruIemQI74Zaf2raOLMLQTgZC338XE
RHGcvYkszL1syNJpYnXXM4ISbkY4aZ4Rlx4jPOjyQvBKva3pWy+DJxAGoAASiJHE
i+VImA6pT30b17NppC16N1FW7E+tuJDw+lDqQl6QHLUUBplnJb324gQAlgRBSqIQ
H1kCd7rxKlBC/08Mcmfpq+sKEH4alF776wO7IVoTXKrGc+ARoH7+1plEWB+O8MMM
oEHVp+TdpeRebH6aIlcPKFNKkrlLPWSMC10uuvOQusSt4fuK8f0CTej5nCN1N38n
zo0xzWLF801vRa25ngQVluzORJSVeJyvyP9rPBF5IB+UeaKzEXrWrEI+lzzfsbnJ
UGP78SkHI34b001H21xbbWjKlEiOcSQx+c8hpEeNzxnazDqNQFg7pws5aY9Ce76x
Eoycqsxx+sPr9BbEO5dDkH+KXArgLm28GaPFBSUiNMHE0kOLzMD04y3Dq2JDu6DR
mCpr/bzKwtFs8ZhSAHy7yi97GKazgfNjkDiCmh53pqvYF+cNFglxbx/bI4uF7c3o
Yl/UmX2dG1GlK1z0pUI+w79BpmZMVWHuPeSbPQ1zhiWZ1f1/dn/h6czdouIZL1sT
0IHO0f41JMCaJ7VsmdyMLLyzy368l6Ch8tLReyDk1fpU6dA0MZ5XVay8OoyVpwIX
RSSfqoRUza6+0f8AG+3Ap2cfxcsi7wkxSJ7IT0woiSwGZmm5lJr53qgQ5jDAcqYQ
86mkJS3vXkBPU8WIdrZBoDsd4ztQu7hB25y4T3QerGe9WIMpsmKcIIlgi0sxpDQN
adae9+rSg6qLi0/WyB9A3PKR7q5OxxkgSWnAQIyJ3D7uRHuCBQlP6tbhZKm9CzWk
jvcvDM1WrZjP+x5RPjsv5JZOr+rij+RvxUlSzF17AC/l/oFsnfTm1LbYB1h6jNb6
J83/oJ77vIpNBEvE5oPI1WScTxnXzQbb5LN/ilk+BHNh7EA6nQ2gQhMDGWlayM2s
T9ouYDylyCCdwP9xkRYy+5SovfLqBSXFxST86bV3ihfw3LQn3Eaj29uSs+7pVcgP
+6P2nX2eOlBBVD9vMEYEXaiAUTLfCNDZPIUfyPSRYwA1F6vOJXW7FurAT84lVhch
jvHgEMjAf7T/pKjl6PaJcyj5Z583VLAVO4tvl4Rz9skAuiPTN51eIa47hixWNdpY
DnMw0bh3N8vyW0TfBMupKK6cVSi/d0SVDKQEeEhqK42LwoCkA5Eh1opt8qoyHE+d
aabgNPbHEuSr4H12woIkqQ8sqqsJrhejH179kCC6gf7lv8RWKQZjAdHFaeyilKs9
iIN03NjsqauNOKJONTosT9iuaSsOJ3kFQn3Dh2kxu6H88QxQQSxkabqe+9ShQzPe
jHbg9kNSFk6es7683E/Uf4qlCcWNHquJAlR67gblKH0MYoTbF4TIDwqUwwM7KSzC
iU7pHdUn3NkUA1nL6S2BlawJgoIGRzNQMQFN4UbDV9jaoWbS/bYYuGVOlLWI78ek
Ct0O5W3ZhKpUWygNlcH0wrtK/ZhTeHTdB/ZBuMLTVHslNpM/pJLMySVrc2og2bwx
W59pKAnkbiOvQo4vAW+zQyA4LRCnLTptTej0w2bPg3jMkpgBDHIvvaSNWxpeHvCC
z4ZxhD02waS4WZdnb+Vhe4TH8W1K5pUPH/76DB5+mA3ZTcUKyhm2MKXKXAkrYQN2
ZSi9SROf1wARvU+Te0UvRu9XiBDMeoAMXddiYjat03IWCdPomniQOxhaUkYn18yd
tI6vYi1ruOTSzcQAMfpST5vEByJib9KOirRr5XQsikXxnrtreBap4ByANCaf3R8u
FfUCPygn7ZLRIkjEuWb+Gnut8Z/VVUY70EXbRMw09G84TLyV6PKipqkqIQN5tGfu
HljcECXsNXizJ7SwSZdt+mK//jcAcbhRweFeA7nwt89dO+TV02xLWOdF86QOYU92
2uUcBGcta2Lu7QOXFqHA7zXTuQuOwBKvOySlfhqs6cppmNh6lIQ+TzW8Fx6OJ9Hf
usXZrZx2anE4KVDsVMgINcPXLFtDT3Os778s1REvghoV+hmDtsKGWlwrhHwR3frT
UsrdzJ2bo20mp0Rf8JUe0ZtC2tUBQfuILFAKSHAYXprA6/XNjOzxzRnNWKguz5pl
cEiDvAwaJil4o+FDtY1vcbuJA7Vuz1b7RBjOaFjCnh0YczpzINWKGNwcq+tIt2pf
yyo8BBvf6w82a0y5z28zzWzw1HEd9vH8qgC+xqm52RF/VuGiRhON8uLOnnyGB5VL
S9Tzeq6L6C/UOmEhyPlvqfqNxtCePgLD2rV3HIXHXyB/HsCDEyz3S3jdAkHVH6sh
NHoJTpgTbCVkqg0Es0KLI91Ll9s/EH+xH2+ayDJybbwGz9VbN8cERwbwIgvXhbV2
wIqdsis3Ef3W/ormYze6UQ7mYts4jxU6IE2uUGpniLDDHLV91pPY+yfayph0p9OQ
DHr6tkMXBSi2XVTrkBAQgdDKOnwTXWcffh2H4ng0t94lBfqdG0LKJkxLPWvi95fl
wboH0vWd+vwifmw1i+3p4eq23+5Q1LcNsvYWVcblZb2RIJLsbFvNH1OmFlbDrEXD
+Ge0likOm/cFD6UqSpqSxHZJfy5h872Uim4OJxMhpAT4jTkU0ngP5hdqokV7x5V+
Q0YVttRVilSaxEkIWXFm2oHtR8KVVi7n3TQEGnH1eEhy+SRWCOEHDgTBU9vLLPXN
8KmEN5rHiQtA5ZoZE9xeY2oQC7Ugv7CDM3/uIZVSOogjENf/qZCsRa9zlNhq4IcT
2GcqG4tpsVfKSnTe12+kwrdu7Jm/FNbEqN1b0orSm/tuiwsvVxXCESPwFuzl5gOG
UNpIACzq0uGblf0vvVxqAoLn7gqBqf4g7yHOj2EUsGHLGBb0gVsU36GSmbEU1qam
h3Rqn093UTa9cBhQQIS3ZNeto8YJT3xAheQJlG8eH2qpjn79ADPiyBnt2qWhPKFE
rC5GWGg0fhWTNug6+1wQJXb0t0Xcg5AHPwG6oRBKD1O53wL7QMeFUEFX5Qk2cIHm
bPRnaY/NqHzD1HpnKPqD7QEjXN9ncsYdbYBaKdE+A000HLbHOR43a81mXe+wF25e
vCr0dwkgaO22eONhCxJztd7HC0ICQo0pMC5qXPh6hIaD03gq6WfMu0wvweI9Nwfq
DbVpUGvqymN0KJQLtnZrZ/irrkx5hANyjamCGcOFlKAlLxTp5eNSoyJ+93ujUEaY
Bzm0JD8avOZmAglVfGzGzY+sB2Ybj7zJJQqs0bJY+1yGeWuISybOQ76GYAJYC6Uw
Ldh/ZFu2fwGavtyiYjL5uNZy7r/QplUEdJqxRfHJYq9lQ83ATEPue4PZ+96C7i+t
KV3i9oUI8OJxnk5RDVfX6DS599OHjZb+UPsUPFjSSoAZAFvtwCF78dlta6NvOywz
ToWFVAW59xbkOsCJTiO4nNJrmesdTNLxEVcK+nnxW0I4Sc24BsauGs+Lu2a38sdf
MuMuH/QFlZUgI/m5b1O/u3zT2TjEBAqjscm+4lRnchJ3J6tB7xk0qvUBcdPclaqg
Tsdoi+VP07k5BhGthPlf4jjNsmwEz2Pw3Xw4URy6Y6bKG9eZ6Yky8LGkPodRr0N5
YDVyN3H1Rsf7rxNFWAsfB5nLGnM6vyI/yjQAhuLG5WfCn6ZXiSXu5EGBor8ygV3A
DidlITgvR9/sZwf7V0fgjmWq0PN/8IKIh9n4EH5Z+jnYfczXmqrmpWwjUfuVurRi
vn1ixPXEIfUbjOj3bqm94saX4b8dS12l1wNzWnKyP3KjYe3Kwmu1NWQccpsrBmVa
zZXi+lL/zL/uxkyBenn4v/Qe5DH6sbXGeUlSwTJeKmbY4UI4oKIMaRgxgnZElaQG
8TdrTJ4YpVdY3d/ailUBE6QZ9oQ/PtLw47vq3ucnKRtYD4LFk65Cu/oGKO5rtiBR
1HWfJFN3FgJfjfJSFgAVF96EqA0qhwc6gN5wOrrJEbpPPlHgATgFZa+0fFuL95L2
Hf7y8Ft5r63Z6ojprLrxgALbLLyv3EOiFWcPwAJceTxuLrc+sPeEFiZo9t/9VUay
A1Q5xFGgB1tJws2O//nVuMCGItasr+sHSL90o/xWki+gMzIiCrrDHtHaUK1r5T7w
1Ehb0Yf4KZ1Y3pJf5ctN4D2nKFa1XNCYeQbZcEFw1y/vLuwrMpSDpH4fkdliwayN
avZfAANoNEtIamyxGSST553ColBdqa5Ur9G7wflBxiMLHljq28abDX3eEGKgsbvK
k/xurTUdGoaj6AmbDZZiPWJKrkMad6wnGP6zkqsK56glFgZLuLMaJ+3yCoCn5AS3
cpdfNgFeiMp6GnN7Xrb8C3IT32DAh7rqNpGvmdLTwuFkbER085nImuMxEYD9VISO
UmzY5fDSguJtQ45s7aCK+r++0df4uzw6GaIWkAgMWqoIH3jNLzVmkD/R3UtNSCYh
CiNplkMUqYgzfPmq5ghLB72lS5flCO5RsV5tcSm3eDPXw/ixzayioQHBb7wTsEaC
6iZmP6mQie4JzFGEL3KOC9hvQDegzjNWjRa2k0ZYVp1/EOtSAs5A15p0Yo2V9x3L
oM3vC2TaO3GvcSc3KGKHYB9FtxDrAmDSMOXW8AwVWmHQfZxaY+4KWwebRT2/VB9G
ZSqkwhbRj7Ah6MggngDzCi6IyIHMFGzKYURfDZtB0khJ9FBIwuUYdWHuEGaE2pXT
W3W4WBtGusMWypjFNYOX0HoSLR75NZa8dOW6iBEs4VmAu92+/CST6fffUT1oioVu
2D2pTb2Ctu2nKz4ejwzKM5rF2n0fif54IMTMcSRqnEC0bqxXXvMCm03+/Q41FRVX
fUpBYCCsUtbo2nm+hnAjd+T4E1y15noydh2663iYfzR1S+WQfRt4fpTyQNgTh9zU
wk+Z70kvp4CjpFcezsx/u5L/MHgXEpXlbJQcBndBDPr08gW90PL95l+3WuJe99ZV
g9OIMbE/ihoUYfNwhHRPyYUNsJm7UjwljzJj4gvMv2gIK/daswdEQ7bRQODlL86i
qEs42OyO8MIEg/prAg0krMiTowQhS+Z3N1wqYt43qO23hZPEbqZbwPZlEkodnr3j
aXMHhQB3jCubpbQfBBGlMpcNsXUDpPjQTwuRKlOuZR1gr2D3u2rOc9xnsVgxvIxt
qXk/gj+q+0GLWVnFTeDjYhJrxDtAiLVT7dvPr9Ees8ZDrlYhfBTEeE1OGvY3gsxs
y/NG8rRHQ5Ke+dSVMAhdo+NlOJCSF7psRfxdRTuMNt8HWvwsxcWHfIJjazEwk/0A
sMYkLvsdIMuA1lDAmo85fqOY0mfdG7Bu38om/DHmHNzqBLBboJbjVVgFhtzGDwTj
1ncNh3i77erdaDfTPHy5E6j0MaOviC/mdasvx6RprAq6tu6ym5JSDhQo5q/jMFZW
lG8U1iL6y8C357GH3VtaPDeHwel6zqjeZGzJJg9VwtbtQcOJTEzpJW4xFAC3pPwA
S7cOEF6ilhS3p1WCpD+BsEDnDVdhfkN44V7+4osht/suF8inL6iFaN2yjHYr5WP5
qakwOIbq7uzx8CXUG4aiabAzZPSFfdcGi+sjzmNDOI2/SImlF1hRkbPQzkCwCjcE
KWg7/GWi6KAkzN7VsvG80oMQgWDhC1K3yb99nM5XGie/YY2xqKTLqLi1Tz062FSw
nvOYXdxmsRd2hQ0Rba7NxpEbFLiube4txWOvx2x540Juq1h55zhCIw8DGzT0RVOG
jniNewu7DH/ZPCjfw6nv70Tk/+DnYBBg1RI6XjYXFCytahXwrbwfemlF6AZDRsV/
tJOoHcQMkABy2zvG/YnDglkyutcW8PHH9zgkGnpMW/MmdQ0vyuSithRsuagKMIhC
cKjJjgL1KBdaBPv+10YZzoz+vbaAuFJMEOZ+hQWZM+GSRn4Db2z9SKexK6op+JTm
HFyG9MLd7HO+r5ulSiobWNrWapw7JwBAVd5CiY4511Fkx14yxY4y21jON+oe9mmR
MyRchadwW4mhgt9YJDwwMOUEI9YzwJfKRlv+2qGODyvCXa4n1R5b23aRC+N0v08E
OOPyjUrusqwokIfGopG7Z2BnJVe8LJ3gTC2TPEXjGZ+R/WGTU+OgIcOtDyaIVEO6
idqgnvoE3Zb1BeQV9omTAvPHwQiEfDLh18/NPnyxUODujXg+63gbzWbib9jc6+3B
bWxEqVw/WqLf8VTG85Xs+Fk25zCzyRvELWYehDpDxgYjNpm8nmkhMyNyoLENnGpA
TdEx3TfXpvhkKXMBYdod4GqsIGfYdy3xyXe8maXDidjzHGfvwNWZ91C0akBn+41G
e2di9dqhrLabxgJb5lWBJoMC47pxSWsJce2sabKC80PtBBAL8m6JXquotWcBzJGl
1qvUnya3prlVSJRt90yhiyORo8rgSUlS/XRE+syX0gyK8WrXapKiHppIuRU7XHK8
MP0KnVMvfSy4N8ZzOe2VAwYLL8VvOy6AJJ2pkvIzJ/2LJKKWAzS+oiyOoc4wcghY
ObX35ryyxyPW7pi79pZ6dqZg6Tcn/fabP8QolDkNb4m5/eLjGD5Ha6eavjfG3Xxi
6HRAD/Qgpla/kEeY/w0ujN98IIzU6YKCDuxMHn6+ceeLT5NUxiIRkqvlzwLLZ+IN
Sw8n9erV61+RxpYr3wOFGqSReXNWgWk0/xvu/fnAC6x3RAEueTG6f9NhCgWIrrVJ
AcS6/OGJ/OUbj9+TRQ41AbIr9DRfp8hluIvBhlH4IY10KWxRmG1La2WTvorVYENP
bWg41WD2KI9LXIKztVR0g55/l7KSrFT2gXvT+PhE5ytg5FnE2jFzTyfWr7XLaggR
Fkb+APl55e4KQQEBPfdMCHqQwLGJEXAQIO9x9hdrD7HoRMZoeCcfZ6ihuqeIRXhF
1Ve5NJfLkInAHm8fFEf3lr3wbKp5Aa1rYU0rQtK5OF07A4U6zJQcnoe1VVPN0Jxx
0aQy3DGoc1cuMMnEALuy8gIciVrO6LuRb1XHCxlj81RhgNN4A4aVh18VyRCFMTRL
L3qR+2kJH9v4gmwFLJTCTEjh6n1MQki8BoMttGaYVQhsS3Cv12pUZyj6sRB8gucu
nKBlS6xQnsQREBVor/A2HzewIRj2HfQQ1bC5GjXYlgXvfdXWFblAopaxhTocCTdi
1B8yrEyrPEBuURDgYsSft0D4IsN43cqaIhAkB/PVi0/vLHGMZyp1nbRydaobhds4
FliEZzBRudt1aS/Pkfmw2+624LANk0y9pLEsX6d6F8Rg+U7U6C09zgvQff+aBlDj
WsIxE4mBdYUYggmijqUqZWhpT8kiCS2UTSCHWTKThll/VbQatNPUf8smhMuQHaxs
dmqxIACv3lq49Xq6Sd40jnMG0etTJkwmQGscMDmgEeElHwAZu73UU9fZqPq0uA3r
HOH4mPONcWlcJS52OanXzzS7rSJlF3nn1ti1Cr0J8BXlGa6pT5OQjATfNvHn7jeM
sFFK5+E1S1txMvu/5jJRhfsDNQJ7e7p3uLD2ArbgyvyADQelTSQA5+h6gJEtAOMl
QHJfShJ/+y5YcDsuHSZLKnoQXYlPkWsgEp+4nvtupSeOjru8WTUr8HSVT0cadamL
tisHeH9tv29EYEqWqmnYjkyaMqQuWca8dF+JOmfKLmGPR6udswSYTdAcyjzVaiIn
TXVJJ1QAKUFk/dIRC/4AjwXqOZoZLtSbO5DROUMKqAeGqkhu27+fjUtdY9cyJpsN
19O8uh6jEcKPtOURIEK54FqFcY9WTQK8OTYA+YQnVNCa3XOjIZrLYJr84EOnUvt3
rFAg3iSqoAKwADtaGF17/7WJY7j/8nQnyk6k4356RubtyuCb9WDPNnFzzCED5h07
AEO4UrZAfj7sFvYWLTHo7PdBxkm8hzZlVgcU71FYfoD5gjEa0twJgj+J7huEJneE
4ytzkWeff0Zd0EfbcU7q/ky6eaqFvSHzstIauPKqL5hhQ9ZsAnv67G8GhaOzrNBu
A/Hss66cVOp4WGNfPkQ6H/YdBtqsWgza7Jx29/K7DqrOH8zCYwh2XpntJ0YmsU67
HmBsALyoBVU+o0NiLtntjPH+XrZlO1GlH23H+O2qfyBPA/PelptSNKOMXmreB/pD
bTH4l8ABgo6Nkm4DPHHztZwCa/tq/scz/tdIHW6/jXohxD9KvBWDfBLMzuLkaKmF
r9rbvaoMmkWOxGwXiBg4WE1zsO7VB6MLVP/M0nGMKVT3Kg5G7CG8krg82WYKGL80
3Dn57nHakFWyqZG5ZyQ2EItsUlS3CDMplIrWRqQQLg2j4UFbe+6WjJTfbNwXAD5C
iVUYynIkyDlR+nd+L2viGGH8uuxxeVErYWJMVz1MCvLqAE2Il8v5w69eIMpmhmlh
0gtedlCkZDHLJWoy4kOYr4BUHE2OE96MAWR+VyjKBlu+mw86NvCXg1uVXRg960E+
gYNbsCtGkhHjtuTc9m0EtnBzqKVAzSbANmcHGL9T9OToRxS+oaIPfyyT8gamJgRX
HEtieEsywn7e6f1s2g9P5R1JMuIAKlWn7I8vVWVL2wDNUOj+aoheVn55eaQzl0/H
HAtVR1mxxdoOw5b6lzGhhK8HLHfY60KC3ILcQklNa1oOBRQjNxo+2elOrzSI4HMV
OkJoLH82IHDG04GhmPQQkjurMfs1ekzINCL4sRriT7QxNTjgzJf7P2Xrd4i2O+LH
g+bZaHfBr71oniNOzJn7ApZM6wV+eWcURkGcIX/hcRbT7ApFCFDfVlIEvheGiY+X
+xO4ersduhT4m/5P4Ri3vUeEb37WY5KNzEY+T3bNSYUJXbZQOOyCKZbLnZUS8Jxo
Rp2D1Nckstpkd27MwM3fka2mrVMKvsi+RpzN2YttBGJyei+QzAIFbDenkYDV+7Bs
mAmTNm+YAZkBNzLidHdbuELCjqVJoIMoygKtLeMKWu4ew0q7DSsc5FHKVFP+hR5g
Eqq5dUW0Xt0lVVA5gC+vpH8yYbx4ZoD4FNw18NJScguQGnctiR6oeBJSf5kdXSka
/nitCUJdx96XFgpiS/GywZvsburRHqRI3gBSNfoFvPAr3miQHoC+VclwhqvPgym9
9c/ofUPl2i+qPOh24rLpqrD3h9KcM9+/NMWbBnUK17tnWyQcHu28npcIhZ3AaTnJ
k8LRy6X4UoDDBWBe0fPQ2F5wTP26XU2D0cRnGZeXeA/sCdkcgVscPOqSJBidIWZI
O3IbSAljwgzwB9mnqWSk6Mkxn/T2XK7Dzu3iJGxVYdgqylqzQ1cJH1ih+2E2k37O
RV52mSztURnegUPsx18HC5LoGOqGN4sT6kOys1QW7D6OAPG8KUY5FIJAQxvaEz1F
NhALF0WMawbe2dvCZrQD9wiWBdHr+toXPvF8LE6HAAh1ffpFhAQzs2Vj/RDEaelk
oxSY0ELHNvYIh2dSHJ8LnNJMnh6yQnD3jm7H7Z8NP2AM2q5/xkXkIbKyJMwso05I
al1dQDc8D/NSvaj+3TJ1qy+d1eTDZg37HzH+Z5HqCvBdRr+ioTcjd+yj7rgzoagg
DySSafVJYakIb9OnxiBxX8sF2x4s2NswRVdbVyrJyTa0tWwkpx61qcAVGVJgfmmi
56HUgl19KC5rWwYfo8g2LFYhU4TIi+IFBRiew6tKCeN4A6mdUkCHm1CwOCPWs9iG
yVDctLSrCQwz9c2VqFMoU36QfCpfZx7IDC82uYVBc5NELpboGVUAnPgTpRG08PoV
no3s89Uts8OAvLfyAKLqrk1IqLOpdFCTF5Sjm6xpI5StDRtz/rLLPN1KV14gXYt3
rOfjxn8+cLQofSe6CMijlKHiHlMVocJ2jdC1AwrkmCAQpUHgYhDL0TEyPK3K5AMw
bFS0C7dS8VZt8sv5guWpri//kbyUI4EOZdg1G3iz/tU27mf4JHj2Rsqy6eUyDYIa
IfVSgSSnB+/4LlsTokb74XN7pk/x2qikNIsESY0eyxaLmtEOj1TJ4e+pUsvBfybI
d7YtwJgcS0IlGINSyKe58jJDiJG0ebVJ+CnAjuWeZSRzhu1hPMnQuUCOMqvZAITV
l0tcZb5V+6zOPDLgvzlwkSQIVMR97g2Vw8CvSN3Fzz/PnJ5aid7gTHTIJ0wijm74
FTCLcS+jHCNj5MnAlcS87obQ2sATFo15iW6O5Rt3ItlegBa5bhg7rAW2Gk+3xdVw
9iIRezOTFrmxZVc0K8eBFmhLLe2RPZoUsUnKwJ9uEASqL0TiBwuMr/TQnJ6wBjWY
ZXPLjcHjhMJGwEvoJkHDw/4ixu+gi47cgkFVFYjuqV2PF3G4h6QghVlB+8ufVXJv
Qvl+5M/1if+rQr3w6x3CDG1OqGt5aNhvJbsdeHToMvRQSxgqXsTC3PwAiyOeABq4
Luj/2JC2xOFXIk4OoqiuIxlMmtl1axzBiaHlspgZk8bzjuUKeAADvxLq5ZpTUzh/
r6eesaN+fFhtrbDkAyWCofvbXFoNbNj5UMa3cre+1cQDcYK8FhbeKetaSC649Lvm
wO0kmx69U5QZtsN9zcIThpPCLYjTA6ir+J4T9oHJsdySlRjqUr1Y/nY2EqNb48vy
LdBotNtDRMv+c5Tg7qZgydcSuX4UBoyGxY3EpsvXRAcPHz/5OmAk2KQD2thtjJgm
EcnzWSfQUcoKoVQVahnnnlhHCvVVx8yWwAshVsIXW4zC9Ld2j0dpuQmPRTR1i1Pj
2ZhsZrUAhuwj1IgoekohFVZU/rKXAWtMYGe6GxzFeKRdd5h6pZ0+L/MjrL6RgHt+
5q39CoEE8E1CjceQE3wG52+uTfUZXwEBtMAtU9ekoZok8su4iyXFiz0qQpv9qc6m
JoP6H1BzBLYh/ITf+Se1wOXOrYeBGfGxanFwGxB3XFa76yzx6H5lMu2x1oo5ngbl
3ioAgvOyQrq9auB15AOMKilEOP69zHz/5Vx8cpBBnIBLCtXS6ZjKNua7nmMRqITi
O/Bcuny1afh+c5XTIA/kkWhctHa5EowB18DvQEkKBDYD2e9q2b9X4g8TSZiIhze0
grEps5LCUyCUVp+xtURbHSsYncj7J1lx7rhCIAJLA/JM84G9MRgAINEVq9h8tjdL
6xKu2e/wfAArp0wt6tRala4ruXrjeUlDONkNJcLMZy67YFoFvA729j3eaxJh73J/
8VCMNSnQ8nSBT7V+zjDy9MieUmER7AGnq+LMoUkh2ZWvW9vHEVA1prtGaOb/dhxA
kI51IdqEYqM9zzHx1+2mDJ3j8W2PHMUdgppCD7asUFCt5Dg1iQCy/K4kd0dmXmPO
lYSuglicmiFzihS1fI39LMI9hdVAJzTuWsYz5tDE3NWuayoKce2yEQMTyvIzVbWo
oGV4FtyvyZjdvee+xIzxZyODAiCc4ps+nAUlqyTNxtehT8P7+zGZKDpKQ9VB8QPx
fEiWKUxRO0ybv6P38DGZYOCNHtb457PtllvFjib9wGKSbW8iQwYV1vY0mXUygeCG
+I34mEWzMIKl5DN2GDxaNXQIUlc3vshhipOSxvQSKXzyp8hJdhSx9ro55nb/u8Qc
GceMA8ZnJVW4NzrNyrB874+cgI3jk+WlMF5W/WYgaH5X0K5MBh99rDKClNGp15cE
MLmIgHcUvbkfbP9CSZRNVtIcL5qZ26cUv8blWAuOOY7TiJDk95KUmvhTqPPNbxdi
x6n+ZtrLy0HgUUTvi/6yzrq7aROqh7nBOjElmSulYsuKTsjiZAuCfj75VSES5rUH
HLCIbvmNxT+aG6Ve5xcFjDlGkBlTYoxrahxJ7jiG96f0p+kI48fa4RD3xUfSnAxC
UXvD2lqHHotB4EikWGvcIRLnKmMvnrMHO0DPkQicriRmknD/NlH+AhYqJTb3c3em
MNxG2e2cIZDLMbFR48jw+/2eiZjMDZvMJacjIvHVStc3SxwT+OmLQoi5E5ajd1dL
IztP7CNT5j+YFdD3iGlrrPs1CSonzKFjl/1GteaBYlxS8a4F4iqEMqMBPp9FSAoW
FChnqwz7YOBWY7hiFusJyy2BqKxzBj3mr4SEGl7qMHOF8KGTp+U31zP+USjKLaE7
vFFcp+WfjYWJgfhgiZKqmRvS/L1X7gZ2KG87ZdbWFPVuuUxLrj+QBdQ9qgxlIEqH
diFO8eMRpi9WG7LOCxGRgTd2AhdCTtTwRMPk700MqNTbVryrfAlTS+Zj7Zghtm+H
U2HuDGUs7AQQ9rHM9reAuepO0ZD4tfX8zR3LtuIlH0Wk6BnY432q3w3UeSu3T278
TM4a4abpXJ3YoF6M849H5UBy0g1AYgXLsZrE16ZwCvX+0O5+vB5t2Q1gNJpCuZyc
/L9INH3wfLGhdKTkAGvB83e2A/nHAkD0+4IuP35EVjdemJ6AYkTSUVahMZc9OuqS
csSOrxv9UaINf4mecYpGqtvThaX+9MAJLpSdoMkqjuzeBTMzyB6N8iXDX9JwVeia
JCirHTL3llQnMC38Nqr6IBd/k2duQUQCXoEu6iZFCn3yxSkIuSYU4L3046Bdut5P
z5DfNOy9LViu8APe8YH7jCYYQKnlkYDS2k93FIzuz9Lupyk9eyhPokQ/Sm7P4KyC
/D8k8GuqTfrAkZAlKRc7Kmypf0ihZvtML8J0Fn5+tA++hWKymkYWhzEpSo6ega3O
0FzmpPYz7LOmBVxjo3BPptzS+w6hY+prJX3kljiB3d8qjg7fU9vvG384IkjMnQv+
VaFrNNNsxlb6b/gelKY3VIM39hroVVKb2AzuQVrpWCb9TOGFwylEHMrRWfQlBOLn
sQlq+/+cq8B90MfeX/Gy1kPAK+aatdmHIGLnnV5TRw1hW4wA8WHOL979jJM2qRON
29rAcfhVEB3sYWwASRjDaBY82uno3awqiPM6g0dOvmwCZNeRmlmknN4MRWZ4yz/F
6UQPiJd2HobIPaqy0/o8SMcTTRy7XMn+inEnfanKEueprFdRj624tLo7boZd4SKa
5KSaCGLm+i50DQsN4JBc2QOYWdeRbbjR75fFclObWYmtmijlwIP/e7Y/+2eHYD6P
jO4KCoOLo/ZdE4gS53mpmik8fYFErF2ohkMyZ59tVOAN40ljrDW16rwfYmwwl668
vafiYYJlZKqBd5/Xw/CHt6OnisjaUqRLvvOJJUFinUqPj8ojNdSMUbKuxr9fDXJi
b8cc51Frv8qspLZ9VJ+1Og9TRiMFTIUIxSW3D5rCgZFiiE30z7PjHdygjbK3TwSO
6GPLxXfFlTB7dzRsCutxtRvsvcDGvFQpiXLg+ad6RO6MI9sK3cd7mghU8hJck7Lj
yvOVWQHJtEdUg1E6IIgTowdruXvKPNrsSqLhcc9hRD3Ke0iC/qyJLy/xpZ/LMH2B
glY9i/Z2hfHDzSTkZSSIg7ajybWy5JhNEwwrhqdM1wFTnQ99R9UrIUfVt2yegTxA
fqxRjK6V9EOCUHpZxs2L6jw+7kM80fbWGn/jsT+z+VkiBuE14cQML2FaNbC3ou3C
5VCF9KXV4s4g/lSbh70MdmKXiDU6zQlzqt/OcQEaMmfS/qX/rZCsI2ueITLjCiod
eUB9gu+KBIRUsN/XB+1iAflxATmQnkg0fidHmhr7LXsjBC/9ewrp2jfHQbRtFJf+
H7pHxAfRRNUW0A6bhddMFd2at48+2k9vycLtYRmGHBm6FD/PNdWZ0TUTEaju4GSO
NEAEDwXm+idW/kIGjkSBFI/noNcvEMoEJttuQpfUA6f7OsVXFtD3ITrNMwq6VuCI
BpZraIzxb3ybYDaoEnefZ5Bg6/D3Q9D/STDybum20W9xzX3+39nm/60++nuCPxr9
ZGVjyWkQGQ6qE93YZerHR1OtQy3BVkSLbyMbr+NkuEsSzdgrEmPTrlb9lgk0QD7K
Y4J3TFqbYd6XMRNmU7DDRS2Zg7xYI0R2aaUK/7sns0Se9Lr8gRQVqwuXq6mNb8pZ
FusFYAZNf9RthkzGwSD7i5P8d1lFUNMtWBClJM2vbSzzh3hTd7L5SgCWD4ckhDnb
LNYcUPQ8aespA9BX96eCWEjOgm0FxEV3e7GJCiXGCESEXRf2Kk+RW4om2cic3Vha
gjLyloQNAl3n05piiCmg8yXdDd2w1hmbViwoHmRt0DWXWG2olDmA41oLKNf4gAlq
8a6jKSV09YqLowKCLpyWaMrJBaTzhLb4keQhiqIz9ScK9tN3VNVh+NO39hyUo6Rd
WmdtRpAke/2KqwyhwhWm1sClH0WnqfHtT7nNZ8Y4PatdwQR39EbAbrouphXKQndn
7EjqxoWVSAaUsqSx3sxP8xXGilGsrpJalq4tFKe4zMrxiNTrh84bBsTDfXQhMNGK
pYzKw80BZMXiUd6M3RUgYDBgt85R0oUSenijBBTo3o9OuTmAQnixb/wTQj0FfEJ5
5MqSxqt+7zOgHJ6BAcMle8ag919qR1kt0jQ7TFkwf5I90Cg+hk49OtUwhC39Jz1W
HwzQckjSJvb7BgseURGWvRudoc3qjdWJw9xTQXwFARHeVTMF3RUXEF+rqZ7jJ8sm
CZn/jsaoIIcB+Do1qkC9aoPUqiZNvxOBZUsdlv5N8DNrvaxv6Iv/G/5JOZhdZRpO
YhI2jBOvwdMakNx4/vucj9C0gdX/enHW+aI9Y6kLnelxDCJBEjk2F7o1rMv7nAjS
xm+eiy5T2w5A0S43ZuYXiet8Mma/Ya2Hi7a/aRy5TccQyq2mQz9LyqqPaNfwM39C
a4UJJU/ph2jc13MK/6URDf4gRIVmugMPZLQgjUZUdIcpQy5bxDRO2LwVfoTz5J/j
Jy1CRhAOya4u4Yu8/d8GsclqGHggtoztW4SRQ5D9aEeqc82RMvDGWeKWNTr5zphr
0ExEWnbpwn44JZGEvxMa3ZVP+kiNVYlw5ThqIw59hLes+qfl8OOSjIEapcsOW9PW
0i01dW8Aw/urUI1j1iVXn/I6+3fHEW8P9U05d9zpBhec6ZkMEEsreM+EwPfz6C6K
aFmqJ85bCXgmZ7329f/He82rQPI0ptMvVZx+IJntRjH8D3oH9nIlqygqDHV3Y+aV
c0S+/kLemfD4UcWW5/G/6PR3U3G66wxVmGZcbzM1hYXTSZlE/s6hhGq7ftUSDers
wBl9ZK/M9PxIBdrZ0Rtmqx/b7gV2vHKSDdAzUV86HQsERqvxmK/C2mnAdmiGDRuC
va5fKc62xXwSatUZC8B87u8CUIuNCngOlFjyzMJoFWyLneSYG91oF6QkMMcJvdYv
pY+EMhSKiHasZji8jMzzeTn+KZ2U1f/k5k4sdZwG0MQaOBYWeC6ndkIc7WWoS8yl
V8gM4hlsbGOCu7tDXkvVMCKzyRbiVSEcMbdRw+RhO+p/vZq5yPAB+UomXmfx+I4C
uR6qgjlZfbRzMO+X3Jd+i9JpVnviGFlvHh2s2ghNX7Dp10498CTNGa9rj2w3lhcL
C82rql/OFTopTd8CmlMcL6hiY9L02cf55dA1Cgib8WOvKMMB7Kj4SrstWizr3pQ0
veHvXWIWnqPiZB8/doXhqgNAOgctbMQ3Zu2ImpyLB48m02kYcc1EEovKROnhZWzA
x967w1+e7vRw4Y7N34W/6GtwfEkYaog8g9gEMjf/hnrT8wh3eXVgtXVezdeR/+rF
bUh03OgGF1wL/HD8MRrLXADoq9mH4NF/2ZGp8Pfbttf4yTkOKkCGmco+DOk8D8Lw
F544vpGTaVxBUwvD/BKrQA1Hu3d0ylZHylqI+SlADnxDncX3vDoRID/7S5idRRd6
iC2HiIIb0+5/8Y6qbxNVUSeuwUPbNY1z2Y524kXuvp9iQyTHAZ2GNYOpFQlncGyc
2+EiqGlmDfcIL+sZqwHVRHbDvTym1Yb0iqQNVlOrU+C7tso76/8NkR4uHeTU7jE0
UwcuzWPbmlzhfHWk96ih015BwT/6Z33tTyyl783AZ2b6qlW8F6Vm2RYRZAszxMxx
F/9W2ONdHrRlpyq2Id2/B+t7T5tJauuTy2wcgqUay7IjIFtCuMaosGgH7lHhJmEf
zF4fnvSkb8lHbyj2yCBa8p4zW0F6Ew89kTvc2UwWgtdHP49oT+zjer5y73LVZEpq
0TqgLvMeiQjbCL6ZiFcfhg/Sg0WBkywRmkct00V+negr/6b05Mq3H82L3QNbfdU5
QtNOOT2SttDl0agAYWlMVRA+R0n2O/+pqLVTep0hotiWyxiBCMcqisi/24lq1e2M
mYWa0l+LHa7jzMYdpR72HRtbexrl3l5Nfv42CJx8FYQeMxyj4O6yuzUL6EvOkBOF
/5H6oHQQZwikMimehKGiPTD/MtWEOqnhZ7Swl9wjAn7ZTXhnMZcG962d4/C8cVLo
eLIMbCUTh3l/HOQHmm0LwRBZwdOMDsxL/3KVe6vVgRt4pOoVYRxpXjKx4cCqNfFJ
TTXvD9UZErog28EnVE2nOhYxyBZOxcxSKis/YmKzlB1OWRXV9/P4Xd0m9XBJfNh5
Eyv9fTWLUclN6hwwXArkGGElzIe+ww/2hF3h6ORH28SpCIINEj9EOc9U+Cc3JrjM
ckW75EdrmFLmIb74MribxVEwYARSoR3Aqr26stEwW0RS/fgm8qOOcYsKYuiSpkrB
6W4q/lcWHnciMS6hMLCVgJAHFVIesAfj570oLsWbbwgCgYbmLk5cNJ0+Xi/7SVav
iXyHRajj9JQVQ0FjaCDRvt+lLzQZo0T48wjvcw6R56J0KSaa81D2QpoIdaQxHEuJ
0rjTBNGpGCisbubt7QVymsxRNaMKRr24hZHMRllHAmY/SRr7q1hE/wyUzoPXuELc
cCA+1VkT3W+qEMgISzBrBKGXMLcRHAbM2lyWKzoSD9Fy6d6xW9gIWLwhoHPjPNWk
/zu8+rSfhYS9LNR/Z/6roufJR+jVFsrDaTO7JThvLIb4wOY4J5/u1qxFohQbrhWg
g3Dq9bQTXExWli7+I8n/M3H2hCO2XcYe6NMYtARfEDsixUyhXB3sUxy+FeT6sRBA
RygGnkQ8k2gZF7f+rb7lxs1dnEoNcnmiFWnvRKSoi4hSLXpbbvRavEBcauYgRk6Y
2WGBWmrnift1UJ+pES3gtqGuNxsMD7vwmZOcgA2Xh+U4r4ZRgXlJWuJN0kbzdhkf
KIL1Tk8NBdKPrAVv42XjvP5YLzTFH+nTL6YxZ5WM9n0wDHLJX0gj8Q6+1AkE+S6u
wfCjCHNTyBMtVl4DPIk3U5oKE/umKF0Op1W551m7FqgZ5vkn1iPIDW8C6Oexgqn4
1APDRk13q8Vg40l5nWKQLBxGm/nTXh4hHfMweUNIV9adPakAdrun9KF54HArACXB
sMzuAz88BgluyaVbD90bzCb4jX1EU4wC8A+Zk6EdeyZybQRC7R13wEFzSaylMw5J
PySNJZBbKv/sbocYrxnflX2luGZ1b3jbVdqtU8huZ9qamZ9Sg17GmRc8pyP/mI8m
f/jkhm/io8c5QqGHJdy6X86FQV8teuX2fi3jTyxXuBK/IdTxyEO3oxv9voFGReQg
qzNZ/pZzj/hqVgd1AYaK+fn+YbRwYusHigVREQeX6bCZHuSmi8ACgPJOn33FcHEw
E+30O0w3wno1ZzKYia7rg696QWi4JK582m+g6qzqa5w4/M6WQeCzhGXDN8AIwEjI
ieGYNliRP9ugaHv/hxZxy8z74qK+ip6efBIYeCFOiijydMfIkgEb7eYEV1fUA21N
xZboX2nRJEJP9cLwlitVos8MDnHiouenbWikwZyY6a5CugpGZQoXCHnBMPVfoM+m
5rWqMMGSHW8fTuYccinsW34HlIxpiLaY1RkiGTl8xa4BrCZuZSnm4nKLsDsgSeuv
gfHPyWz6XLW4EcWQ2NglZhAYbenPiImu5tQcwDvGW2vKQCO3WLR4vtEfEv1XeU53
WXygyKuXTmBp8FiTfHMHgBqwK79OcKBNsGbcPc9nsxKo6om3bXIuVl/bZ61f6f+y
ddNhOobMsE0ulUci0XJ3LMVTszZ3FOk160A+kNQUgZ3sT8CWLmHe4hgab8npgLcX
9OdH+I7h+2LlHka5HKRMgtEEhvnew6L4TJv9JHeAlJQxR9fWZc8/+efXdu5IyosR
6YlyqI8NpLynXJsCDPXrzdSwpXMOFz24DShAupkSX38uro/aE4RQIcIQClh80zKC
NybPFC2Cmz5avTmN3N1tXioW6kx8Uk4ZG1JSAefku89Bi0+awneLcz/jMfLkhlIM
kM4GATlJxmDQda0PzP0atjFgGzd+KGwb5S/BhPr07j/HMuEx6LyOOZdW7LW+ECnO
rfR464r3XFa8Gjvi8WUxe/VevpK8jOD2ob1bILSmRdWyicvMxdLXznevGOqAZucF
fyJl6JkZ8iwPX4fAFHah/RcuIAH/jWRXlFtNn8URC1/VyMBXrqnsVhx7IV99mQwF
gf31AiMul3L/2PyfyELwrHLnc/5SXyOB+z9oJZG+xdDUsIWot8K0ueozDfpoSTv4
fUs9+hd8TuTFNfH/jWp+vGwUzoq0IKyN0TB/ivo2Wb8z788YcCVnTIadYYfVfgt2
O/zinccS5SrTto9U83v7XcuUnUNa6+3ys66pJ8Gm8qH24uUf7m6u3mE4gAtN4Xsm
6pJHYj9H06U9UtCHtDJlpmIx7CMsWC2Kitl4XIQVnIIQ9rClX2JiKZe/0NFxXf0X
RAfO60rWn16aDUnY/if7vfJP6d+9KtFSBa//St77Uu9ZfckuolLtAPJw1DtOeSOL
zAVxmScUP4hEsmmPQAfBkLpNXrUtaKFIwZxFQYeI2I2Wj/ZH6pkcux8If/eRF0YX
Yu4UCKjm60ylLCgf56FCy4gm9eKlAC85k3D4fA/mjHLnr1QjvW+pKx/OmxiPm4cc
Ne6rAUkoVyTOTmxDZSxq+N3D7Itjj8S4xZCowe0kg/Y14hxGbb7SD8vBFxDgAIE5
D6cjkii9fVYPZXttrwQi5QnpAPKd9G2k/e6YEW6r/d/LT4XpaOSu7NwNkMlNLcvm
TkaN6CVkdA6J4WQiZ13NTetyzkc1HB5XGTxToVrzR1qeo2idnSqpLpAw9oloUHeF
y5Ha0FgB6k6+8e+6DpgUbUaMggwG5W3B6EyOSh2udNWnI7bv2jGR2aBXWaqRy+zZ
+sbDnJ70K+3fz2HYHmp7ktKogqrub1FUM/bSOh29f8/fw3ysnOHFmHO62gIlQbtH
SwOL1kQMNAJ4UbrYPr0Xp9Gx5BqgcLCh80G8E0nZUcimFat64WBJ4f8fYUy3Raoe
7qPX8FxGw+dliZ1FtyawPzTRwnbZXHPy6i1GC08QKnNq3oF85BDwtue6GZTdxzHv
YuAys1YbdiBGmcS16rYTVKenQETWJMxzRuQRcL7x4wwjPonclYWYyUifJSgiRIwZ
rwNKeUG+6jcwiJp3rqK4HHG2XfDbQSI4GP5XKsxYVESTlb5hpjfnusOeMi2k9Tt5
bCZynGpg46IW3MrJ7OF1X4NjEg/Ripx9ikAoFOIVX0ThykZMaR6ZxAaL3Gvz9VDh
qt8oStImxPBxJhYxWaQNoLlLCleWCgAIPSQ4/+bLVZUBkiLqtbsFfyMbKYF31YNA
1d1UeeUbtss9QN8cqMFeYNXYKlhh4ANSvCHoInlWiIc/6CeC9AoMocghYx6D7PdI
XVdp3lxQADE34cvX1hDzr3rPp+JpU9YQLV1i+aI9tn2lyxRTxExnB2tUYHykSWTS
FXZyduNJU7zdmVwQ4Fr31v0omWgNpyfRAGYBLMUpkRz4FgP40SbKvh4ZI5axQr/w
XsRm3xurWhkVIGJ9lxVDEvx2qZeD/VpUT16IXbRCBSyqaawi1aDWqjEVL4R0R6z1
pthYQlAywJuSXOesa2m08CjJzS3VFk54oTl+JRsXBGV/UFpjI/q2ky9t5mpgNihE
9MoDNkQwn0USBS5KyZSYeUjz2zVOI20X0avdyKpjSnA0XatCT5Hu4bWWOyvEjT09
DZJArOyllVjGmdlHEZjgqh7FSPa5app8osi6iWc3oEX2N1ynoxShiBaDky3audRW
K2Kgy30JKims7aQordyUAiHBTPM0DvrH7FiGa3vypsvgQA0pIQGBgyOKnpU/pvvu
bLPVXBNdkaosTJHQeaYYIl69/uk1x1ID40U8iO1DoVtDup0ozyuGolJdIss9lT/E
+Ta6TpiKnzfm0K+qdCDG7QKFUGzLG9dYvHOOdrkJss1n802zWefesHQI0jWjwANB
Usk5Sl9nvBez+dWwqZkOx/AfowypaHh0htwfdwCGvwygjU/bqErhIUT+C10rIj3K
oBKzv4syc9ZTj0aY96sPcgSHbl0Ji1RR3R8yxU9ryM6sSTTmSmZir306lDdTRNjU
B8hqNByECkVXwBmXpurInho1GRlug/F8Didlneu2+2Dt0YNnSh6r+f9zydH5qdnt
O/d3p0333cMJcW7oUP6WiIWLEPyEw8V7OOmlst/BrMM3tgWXsRpP2+UNlcUgcMfa
cdTm19WhBer+zRkph3d/0rAm/PXiZxjxGR1xv51cOU4QXQCS90cq1wnHutPNzn/d
t2Nf7D8d7/hNQYHxFTxQYIcF1ATagDYMvc+qw1BpHNITERkkMlbQzk3RW16tQ79b
vtLx23KBgJF5qKG15BSeEDMEqDRXNy0aBl5a1B6BkThCGZdOH9XzZtH8+6rQVYSR
GWKU+b+Sgcq33mjGJG1Di3sLhk9S0Dfay5XC7qwoTjJCEpaD110fp7yXc/wGiBQu
EJj3lEITZWmY2EBJs3+6nsJjnFl/VRdBk8W7ogre5CVhcZNd/iV4+aXg08GwPHYo
kOKKKejhCLjghYEoLBq92VfTek3EQtDgKC5+24C+X0lLsXRw5h+UhjPRZK+ksy06
Or9SpHGJWtyqN57+jhjqEHqTdh9KZDMJDJoJrVlIa1wnedUSgX+kfUK9nUZbdOC7
Y0JR/f0N4m0m8tHdjOJDYO5z7fErKOEiWdXUSgndkYhxZocST5cOB4CWIIXowvoo
DSO0HCeCqOkrHZOc6Jh6BgFi7GcVadIoEoJBpjWrn1DUNKkJTGVaJjSRLSSTIVf7
KaZpqLgSig5KhxjzV6h353zFuvvOs9kviVHn64pqG5UZcoQshNqS/G18E65xed01
Tg7q3nMkmVRyuNqE3k0jEjX8fLeN+D2PKwg1fwhhsQfkBYq7dvTD4TCeYiNmt280
KhK3tz8W7NM9otxVWdpFXa75yExsmLRLSnxZTRyFOIeeApECeVQe+rYNOLlLFiOP
u25pP1gh4MxX4pLv9UuAACqjkMomY+LIoFw3/0ojbLpNKMFF+B/FJibeGtrXMppf
kv6uJ8r6x510b/557vOvOgq4p0KOzSIy6yr+/qwd/t+IdPoiMEUFn9e0LHospkHr
iE4n2mNC7EBJIRLIj/kvkyaKOk0sN+Qs7IHBsX7QQj5jY8Cm+W8LriM4ur3omOXJ
XBGpwpV/unEbLNrVApIdNN9L3rkjVpNigyAdj5XiFnpdBwJ5nt4IyMX40XfFOsUD
vRBCiSTPtelaQLisIi/k2JW5yNiIioCizQNxGvMVC/bulea0uTVCayp00zsEkDAm
AP54AQKDLZ6LCZwF3MnMlGo+714+teQQE6e1Oxua3opka2aVFMAgOkl1yB1HX8ps
gY9sUE3g/oUwbCjbTqMHeXdiL+xhhPxkBmof0HQIUyB5KWZ9C21mD1gKnYUf53Xm
bu/RQN5o1x4FnG5Ql+RzRF2Nwbj23HmKAQEm8VXLhvj5eNggOSmEb2cf0IE4LkhK
/WiPdPdxeffEl5fwhWOWehHOM6skMWxk+md8C64U5P4Sl9yNZL+q7NJu1mvvBsF3
gC0RfyfLDDFSp/+Fm7eOLcvftK83p+qFX9QWT8Fmj1v0qQFjUTC2Fmtbfgd0DbZl
rYdJih/hnLJRyYQGf4dyvOvnlBK90cimF2HqOai5sxjPtt5FU07LAb2BllsugV4J
s8MWhczVI3cWOqjpnEIpQRK+1GQo+o7RLME5SidpPPFmZgS1gpj2Xr2lG0US8sFG
ka7t0H6noQSbHMNkSrarpRzoDDNg3lvW6FAeMbUTCmUGqlMSajHGaZlz3fiomMUp
C2V5uyFdZa79krsQ8QfdS7fiSjyIK9qH5bfFHP+4F8BoePPBrWF2eA5LA1uTNz2J
ObgwVPP6LR0MqcU/NPxET/6pX5i2k4D7vquLdu+bs5QtviDnmV0JFHbMPAft2g0A
clcnY50TnuCvSXi5Sn+bKSRID9x5OmDv80Ef6SWXgKpqozmfOUH0TWeKP0+nc3dl
gojpbgjdynOfxZPPj05FQVs0NYezJHGNHyH5zcY8HAPeACA7tBHcpTabT95hJuTU
r/OkYm9Gh0krwEZms+blQ7YE2PaUWQxWZH8bZD37caFFu6zcGwdvnj80OyQWHzBj
FwTFTp8m7kINQbBfsAHfI8hg0v+iNvaRE72txslxReaQCLbbzhWgFhNhvymmVaQ6
/HS0nI82ZDhSxvUjgSNnNx/sBsjxg8FzQULwUIxiIbtTNVSaLIt1WM4ZQ9C4O3NS
ust+fORYRLGSLRFYTO5YACLXkspxtrC1o+ajC711zLT0C6eT/5IstKohkHbicBtV
fQGIbFyuCevLBHwYLUSgPQ0tS2QyjGVYFKXYddgYCl3ID7tr7d6E/GgShiom2iBo
F3TO7fwfbOK3D8GobkPCxIhkQOHXG6f4uR1ZnrNYp1J6MJouo12s1EAZi7Xuc+Ih
LD3PIJv5ct2wIEV51Z8YievhrgYKVMWWCJ/adXXphlG5EK414ag3DM7ocnEheoV6
eAVrZ4yRkmhoBHYocsn5MYMZ1OwOF2ukBntA6d6x1iGeHts85taGmUDNehb8xZ1B
Oxs+Wnbj6bddDejFcFMgrJzMVJe/XRhYX5V8xcHeThy7nRjij1dozQtA8Adj//bE
MA2dJe0vUEuFwi2C8bygyT7VI3AlSk2/8hWjfmyBann4EM1rNZw17WqKzNQYYKRv
meL55nlSbIfNDOpyoXhh5NwF+Agm40jUUcRw+0D/cfxqHdvClgSr8bkm+BZO/vb/
N3LnbU1aDaMsVByZXxdFZuFFjz4cV4DQm5SEpLxPJTWY/seV7CEQKoVh16q1aVOt
xWe0vdQNG2nlogkZGvbIcihewUtTqdeK/X9m0KIHgma8riPjWA4LbMKdQLzRVJo1
70oRR+orjcPNsQiYCMTbuLFZETbyWcUJCV8+Ias7ao6XAWw93L71Y1sn3SsYzazZ
Ek7fJlf55xrFPFVP5sipMhmZn1lbgz2+hlZ4XxGUwad5Kh70wqI8lJdq9slusTyJ
BQyH4jOdW4hE/bU3e1ARSCgIjDBsdnVlfkPuVTF6/Kfw0rpElkVAgZrOvCshNoUu
5zoX4i8IZi5PkTKQZcf0EFbcPkPVXFNI22VDs8iRBcqzXjGyIovb9LxmgCTl37QT
6TqEvUr2vkwbqs92Lg6WaRr7JGPzXGiSeg+fpftcOmU7913cbLaTZ7DJ+KBvHyJG
lPkQIGay1GlU1PqWHDLso1CGhic77o91tlpPbOrWjTzRJIn3EVCIbPnGhpTOkqFS
cNEMCwyyqXqPYSUAh3smCagCjRdole+aSj4wn1nNs2nPJF3BhqxaJSkkUYCPJBWa
DUFNp31Y4JVjKFLCI5YXE6mY1dvE7+ugQOlem9rsE9qkU+Oz2MGX/SUWJI0ROmog
OrQutlO5qvo7sYrNqPh8gWwfb6f+n857mDNDRmL/RUbH6qfCMMNBGijsG9P/bK9F
8x6aX7QvGwFe536fp4OhNaIBy2u8+myO7wupiKd2M+9o2pLWxHt7QwzsJwlIH/M5
E0CQsSPWH6qsdrc9Bcs07k1cPa+sg2LygO2zMi9UQMGAZ/SkwGTguMYER5QIpqUJ
CvMZoUu4jbu+d3Prk+YOyQl4U3CmZwCi2sNY2rDATIB+NcF8U9fD5Du4nET9huss
Wmo2gEjEK/UdbIidH1GbMvVHy5R/SuaFWA5gjGL6b6ujA6b/rwo5j4XAdh6jyUDf
8vi+2/wuv2/pQ0toJzs5knKHRFQQu3nSk20edFnISl7ry+22YKjGDodYwqQ+gBz5
FogBpKbvnNUedjogZNmKApD4KsEXgpjCNfstefYy1IltRlJnbP8hDgjtl2mQcsPm
iyt9dj+JB4/FSPJjyEGc9ScBR0wDBxC/PhPaipfAE79ipvHKrIZ40mxGzm1MYJXA
idR7ds8rNPtz4z3ro4GTQn1AgbRF/S+YzDaI6str8AVv7a6lnDAnxa/M1kMox9ht
za5lTQ00ay8p3L5BQhNvJo3WjzNe3VoU2e8ZARPhJBR/eXyHvPVhxdVBiuUhzNyf
alUsDCIoWVGGiEBiJMqdyK3bIStz90DkoXPibxfpet0Z1n8PWFExhfAjlW0Svmks
yD1nGfMbesIBMJrpNkf8I+S7BnZTflfSTJQB9u/kSZTaOKAGRsS2ZPz76y+mqoz9
TLnTXL1mnGp65tRDkwDoWGV0SEF4TFVoUKAlJ9K0tXm9jqCzSMKV97x4O7h3TMfL
Z118PzaiwLfFMG6OWuSnsnDU8LdCxbwfz2DMUSMblSdG6AUsDaRQrBpEEOPHCx6D
5UjRDxbyCFYw4gC2SN7Fb8LksteplJvdtg9fXereVcac3xB7qrNyAM4+g8Sv1XE5
b3/m6uYgbn5JQPZj73stG616qQmTv/Q8f79wktG+FMYAYiKwoY6/kEQcMy2vn7St
D1QpYYAzceVDXWZv0AxCsMXufIjAhhEvbI5CCJ1rySGh5SANk51Y/bmzvbVUhK1f
CS+Clh77sR0+8amHOiBzleNOdDh/3z9lM5uMSHx3LE7xfDj1VCKMP3zkUmxfS8/v
Oyu3wcjaSZ9mUOuHKpCXRhTvK2Bzbc4IJyMLRPKwISIhaiTykmAB0d0B0R974dSD
osDGka89X0HY82VmULThN79yuKvXKlQsI/TWJBSocdJr/i+i8KPWK7Ho4Iebxc3A
NSFjxs+s/7FCYRKGUNfCLSz5al/c/Foja0yvgvtb3d78S6ePQ/qCrNTpeAOkmavj
Qnk3fzHc5+8hTigG3Pgk5N5MQ1Ko4OHjwvD1hoStdxz4+vei2iw6F/5vmPegUV6p
qJ3zE2bXe2Ui6nd1/EGq2Y3Jb7z92WOhRGC7/KweqMSKcEBq9UQlM8Xldir3Ia6g
QQuCERX+vBKW3s9sspPZxo84pKsbAhG9/AAe5y4ns/vijCsZztaHiMvs6qaoQqnd
Trkv7G2NJJTuxuSvDaLLCxUzbwkBkfAF2PjC3vkRlRXu/C0j66ii5ibqfbVDairB
jzqK0NfpOprfPQRpy/CSk4QnS+BWSVrIFCsJo+qIDTAYyrksFOkRN2+ljciwXWQY
tI00KGg66SYj4SN9PCo1LiYq0+DTyc++aKCDI65bxD9GK4k0r+Y9SPRMbbIene4G
yM75eo9H0vfKBL/rxizp8yqZOlJRWuDfeb8t5gDcjoFpfT5IjXF9BzD3Tj+TPtTY
jR/9TwbX9TAyHBbnS4qXl/wGH5ngHIva8uqMlIBzWT629v1AdVuICXkWmqeC6QdZ
LNSL42xnHj17iu7BQKLSt8Uy03XqNfIoYA4JVuVz8r0pdLguSwNUN/wbtRmv/5ul
r/A3X0Q8AIfALWHa5hB7J9isBbBXqPv+bHZG+/7cxgR5/MD4ufReGWjCP2c1OFJG
Heu9OLa36OuWvIvt9Cbef39qbOwYb3ljJuQST+EXT7iWmMr6oxQAszSi5XyDJP4G
tl785GEF2jjpCRQTFoWteZKFUknYnQPwBvEHjnZ7vSrvckoinlE10wgtHlP8D+Oq
QT7YppTpigy72esi5NnfNQljo6rUmydcbrvpUINij7qE4Cgz2y3K6PR+94pwu79/
wTYmO18+yo7NEepAuEal3f/OEgQB++MvB5tk96yhFsaRSa3KAnXMy2KWlort6YCd
xMwIJAQa5xEHfaRT9NaYSrZL1FykLZ7WvRyIMWbm2Mz9cLddp5wNNd0jJfkKcMXv
C7BaEHvFkvkJHOW/EcxMCGOtqkXbfzuCEB6A4x/mXszjf9JrUOTdlOJyNFYnzQZX
ky68BWrxnFrX1lb8ifH3BVxVD5RaUWDSokV1YW5TUzQPKsO21ktdetSOLWa5gRD3
bpJnaiuO4+tKCrrYL2Njd81D7IHBW98R30HipL0AYWT75dpKfplsF9ISoF5lrEwl
gGrFiXj7+kGZT6FdU5A+Zt8SzuPnX3S0FoeU6wNr8jolojKKnVhJtNMEavNGIFth
sJAYefUwUoH4O8tH3+nemXYg9RiDJjLBejKf7vwgCdzIu8NORjBtPGvjs2UJl+wi
sEQyxyQjDeEXGPI4jBQXgTjaR0i+k2UGRWsyC1RZN0hOR0fRN9imHBzCFRRMngmN
KPbnMCA597riiJByVAFIzIg6g/XcsxzVYqsl1TEKuAR5uGBDiG2VFmfzHwaDquKr
Ayi8/5uYPAu2Je4RgONuCRWLL7UFuVwZ3pn33j4rvU5hBkYA+kiZ2J97ksx7A5mD
jEHHwIds4G5Hp2Od9quLvs1ZsKAUbQkkuCb+eTbwmsLypjh732bQJwWRRKsZZsvC
xMXv0w/cnkKdJ2r/N6eTUXOY30FkFTtd7oxjnBl6XBCFcnBbYdvzfyT3NfaGFQIb
fSS4NgaUG3auoyr13xy4Bdyg9WpGi89292OnKZ8aYz4nX9734KoTHL5c8DgqjfD2
o9FVDsX/iLJCvrRolW9RUTe7SF83tC1QfEc5tXwFl8bh89u70Yg0PTu/xr6VMjJq
gi+As0TXTcm9Eu13QVwJhv9CIYLEIqFsDp6muxiHsrTrQ+4A4M4JQ/nTojzuJ7cx
RKNIyvWfjmx2vIfyPN7Vhs8VSMPL4RPA/M4/NiZAmhyjZjFYmHFqeSPnHhWGBNPz
KKSPpGEe1gH29H9udwQ37w+F5g090FiygsVeooAhDvveVMN7ariLriJG6ZLBjtbS
3ZPosvcSR+8i49nIm6BLnaEBqtjFIOBK+U76l7+1Obibr7U+zLGBWuFUfsNy/q5D
UAIOQRhVD4LxvJTEsQ00Q1v2oYQliwvh4iAL49/KAGqIMN89GM7T6Cie3reQgPq2
LbFlbxe1dwZGK7tck85846TnrKfeFFqABpmmjWKKW83Ra5tp9OTOpMPV9w8dFDk2
gO87iLCmaHSWjvMXHaTumD/RYUBodFZXjCdA0kJH5QW24Qx5xDraQ5i2lh3BfInC
Xa53gvutNtEqDZD+HaHFgYw0uWOYKg11Qqb7TjhR1h9W6ofZu0OeK7C3qoR+s552
k/rMlvldQq5ZS7GtFKPEVkpAiRyy0wHjfK8QlfC12d1SXUCxq26znkebZv6KkbHP
n8ArDDcqGIpE4cI1/pNrDN61R0GGIkmdGEkh8upXc/szRZA/upmkVtKX9qhNW5+b
+Zh/KmIHrhqCaf6nXMKp/wJy2Xs0DsMPr+SzJeOnfleFMgZVFGFWFmgfg7dF/Jmw
SJZSy6W8eDvI0SoXibg9yC7uQBLdOvMyiY1Y5KSFlM9ij/6Sfcid7OQ2C19cpQKg
xn98XULC6jsYYRQxQbU/ZZODfsc16JfX4V+WulK436HTqAQ7+OIRJiLkW4LRvixc
AzYShybQo5oOii8vuCnLms8Vexu9z6EZPGAn3MXs+rh6Y6usombPpotTc+2kuaO+
SUUkKJkrm/xEVyGlw3vO2yzUYNue1zyQoJd380Ho0VCnt0mjaLZD4bePpMjyFrsK
rYoncag3Winv3f56TgZNn45lHfLlAPwxTppO0SgxuBvLNz+m1DhxTXRd70YJ/OY8
N//A6MMKZGH0S1lc8yjvO7PZcEnw35wU2Fdv8LQHHZALFGKvY1k7mJ1rZQhTdDXT
z/fKIvFr1ndaLGQ+Ycjr+vwC5gFMzVqoqCGh+JaHp3WfReom6LX3uGE6eMxeck0o
PpouPESv+F+zAEOm8O2cNYRo/J/59kf9Sep7AjS18LAtUSSkDIrZBJhvJT5BUNdP
sNo6ruwTj/e7PFF+yIUHAX3vfcYRRWJ1Uq9Aemr/HN+bq9RmGSi9eINUZjKI/L9p
qOEgC5Ctp+qNgmKN3j1VOuf5DcRoxhUKmiayHRKZ8td4v6/kTnzLelzCbUbA7cs1
PrCHen8RmW5eq0S10saR8qjXt9xiBSMpKG4ZENNFbgz/IMYhSqqo7PFIJxcDKLe6
ewa+n5AyQ5M82CClXGMHuU1NfNAX/oOPdFUCGMUp9ilaadSboEZw2HFcxwrosHhC
7jdice7jzFg7r23w4sUj/IutO/Qp8vqZSI5GqY2Gp8My9SS5CvAHcD1xpVXsE5lS
hKVapuBCcSAu/27snnUxDPbsNoOMiXoYqn+bliImErbFYQbIn4/7DUvuM0Lz98zM
MESUg1uqoDqLKue7bM4ydcMRZ2Q9AA8uQt39clLdorltoWZEEQyuAhv1iaJ+k6r6
t6gP8PUneRe/eWg9/Iu/dmdnOpgzduIAuSkjnLzdyj5GvlIJNidNwAHMRW7yBaZ2
3KFA5xqvIP+pK1b8VIVmA+e8qRgw8AYydHq9Io5BXHpMjKZ2vHWJuYh34Bd9FqPR
0et1PNPqmAX7X/YsLxvzLaZer80zyfDY85jTd7v7Rb71+PpjWPWHXW9eNjn3aNIo
iJB1aaQ6clv2nKvRkgfp3N4HGMLCcx82szPwd3+xfWnMo+NR0dK/ZZBoN6j6B2P5
/DPHg4eavENcLpRkR7Upoypeua4i6bxO8KHGzz2iCQ7W624a/Bw3147pMMRJYfvS
36LIqYr8wusckJ6Ntjq4SejbI7eOk7OwjLZOb3AZQ3gGHBSGr+OCUUOlsAwMRYHf
t1qvhfe9LaURmhox7bvRB8vuflfj4OdE0igdhfb/rGbJvU0kvvWxLtHf34gIsfch
Km/yPjMEjD0w0Puva3dz7Zm7KCwcq0tZZ5CSQ+XvkyUmOOc1RfhEt39RHKtdtvrr
XbfN1nFco3lU0WgRQyWCq7+bh5Qr0whkNRnRDr4Ec1ECwfQiXh/8hmD4c0go5ZDa
XcPK+HejEMYJ3jDFsGq2BJz7CYmzX3VfMj0GN1qHUTRJz7krXUV9FRW2BbGaI46u
1QzcVSkEdHjE1LP4bCzehU73aOepIgFcfm5U/XeufYhTU6GZJ0b9MHhTRXfK9IUy
1BwghM46ZVAW99Y02efKsTVluad+n9YA+Pwm7hagFziNVYN/VIPIV/xJ6kvx2XGc
RmNKFSh5B8+zMhQ/HUjZIBfDD0bgYeKH+chO+Zc6jDl6qCawtXWfPWXFON9guJhO
VYp3sMXQ3IW6ji9Gc22otcchy52soYV6qxO2d6az0CUovjBWf40pfMjGSW8sFl9Q
kn9urr1r7r7b/PtdXoCKUnEdZIjbkihUPpwJGB9FvUUca4ievUybC7775AImjfNJ
J6bpBk8P0+p2EzxvzPsNRx/YNtWc8bnRj2CFb/gUv3Ixhk/ByBgiy5qb2V2m+3BO
pk3B+jCwXl/GYIqeaAzTz/smW/dqaqzgC061lp/mXpQ/MB7OWReVcQm08PSuynk/
C7Mhlu6GRtilBzLK/EzfyFgz+UFqryrkfoAIjPn9mKfUBR8Zi6w6f4BjjA+CRK6R
Nn0bXFoAIBfYrf9KD3AC0lAbI9jHv1jp1HI1vxHlYZVLi2w8w6wjprd3IuAzmNKd
BNmQOl43U1k2n3uVWanYf+QmiLj3c7H/9kIbJOpV60qdgz9c/0vtOz5SrXwou9f2
bzQC9xhv7yyr6epniUJXK87BF7cHYRoFn7+pF7KZ6jZ4//HlTMQ6+0WpLwER/uC4
CkJJvVfiFLCdqFX/77PZyokkVarBzlgVAqSbzr9gfnK6ZTsw4RBb8xmfrutPykiC
JvIXdHbv7DVjs6YnQq4C6aqO0Os92dFEr2AbhkqRJ72Uy+x9QFRAO+gchTaOwfWb
qQldyv/OHHI+dPaiE6jnt7k4RmC0xWuD5KP+TydocTMg9fHf/bBGZysX1OoyA5rs
eiJaegjsg6G8tTUpjUfR5faUeGB4UXZk7/223OJuEHOGivD2PYQsi5iMxXg0g8nX
KN4N3wsaHcruaZDkTzuwL2Mzv99NPmPw6xJOxKiOqsBnfevJzBXH8uw8d4KX2OPi
h5aFxib4I5uMa6IGaWupmu9005cuHLM4rF5r90Whr02pAOLKHoak++sPE9Me+zWk
rVhYtz7SPIuxNIe5Vrtzkp3t8hYa29+ZoeKqg8oGoZglKZ8uFrZnoezjkJTmhIx/
5uCFEp+L+7NYlCmxL+OIuVX/uAcqnmSKyOgeKTN4l1cuKe9Guwgh7twmCBL9nJwj
EHpytVgTovpyatPzXF+rpe9A0MrCTptaJHf8dLM7lLA3yD8fvm5bgKbcKQ3SltH/
EZw5v0XjM89eOU5GPVkOEkACtOELrMN0DCRqp8mdhh/sIm2X39NZ2GJgV476GA31
oScMTmuy2CHNcf6gwt33tGYZRG57TlT8JXuz4tYRTaYnOEwHxAqlM7oB2NxmAbaa
9ro72IApHa20ORYNUMeYTVqOjEwCw1ULLcKPD12EQOcMYsQRSriUuBo6SYkb3tH0
bKzLY9TrCn/nbbo7WYSIpECGik9Nua4hVLNokl82P0Pms1ersJp9XRJXGTo28Dq4
VMAC8q1isdCCgNE8mXgdK39/9gvNxdHgKbvRlOKHmZbXG32sn4IwnJeBXGxuf6Hr
PA80612EjDVnKfv6RdZMmLrEv8eXrOJyN35AFK0xHhrlU7/wifY0EHXfCrYllTeC
75r/3B/w91q80YT3mgHEZv6lK6T36AtJyryEcTzDkVo4aqLK8u4B9MSRlcMjdL2I
RiZ/JkMLRcyqxZDRAlXtRopGzfClKg4HLYWxh7oP9n09wqXtJTN5bwdx4wOdADbo
cB96Ffd3SKKKQ59gb9uDbuBBZa0cgY8ldwUzH0k3LPGgKiHMQ0P9ZXXmNNNwhdD3
Y3kMqGYMEXOBU4VJhWrxSFu4Q1wpWA8KavEnQVRamyxRhezCCKTkeAnMvCJ9iRz+
7KYiAPXlthcyi3Ml+94tJMPP536Dqd3SkfAaznPMpkhpEZbIx7hk+3f8F3+ykSW8
KWJO09/Yc0GteCXYhuX16ndqpEnPdcylQ1IwYKBtVGWFdhdQZZtqym/ZFKcm8QLn
mH2i+BgnJ/SjwRlV0MSl29m18v0I2JpCcw9l7e2QJXppI4f3tbIaqZLCOgD8TSF/
Msj9144gxFY+NTgbGeoNzKRDSv5z6kSz+1Q6zWneDvmFyoDr1jAW9lsy8fivKpcg
qSt2ZPHOmghjHbvcs2ck/Z9UmXD6/r3o5uD+BKY1Pp4dMQoaSFtPECxkaG3v2Sk7
82Si3wTo/fSZXmZkZqX02Jro5qmOUrDKQ3truaBsBAX/EX7DYvhTXutmzrKlCbhp
AjEV4CzHB+nFn+fLo0kcP4tXZ2xjTbB7GPuGtcelAzQMGI72xzR4vouNGykiiENw
Tvds1nxEKbu/wAlXn70cRspk+qShl71cG5AvKfB4Ryb1vJKfO8MOUNcmUgQFW1f/
AZiEjdLqsDYmCz6n9zOLgWC+hA1m2704yw0QO+CIyyE8vgjdk+q5van/7+N2Yqly
6vO89YRFCM+ZADd8oFLWh9JZXWEY6t1FOT39CJrdP+0mRqgzw54PZ+yiuQVuTduO
9XTpCrPkZvQKuGkon/feX++Cyy8OfTyOKMg2uqRfswVmPkmXyh8xD10vDm6f8dfl
nJ4Jq034Z+cxVVCxNrZU/IVO3MG96v4fXuZZ9easWyQ9BF6uUgTXFaodnqk2h/Wy
uuJyv/O1VzzvIqsrlgRGH7Lj3s8O7Ppbrbgfy+6qVSezrBzokjv2zlUDgR9Pujo4
M6Mb8cbXPlLzwb4ZLWOBPhc5tO3cqyKEgLSNxHsHiN/+Jhs6KyJEWasn0MQ5jQ6K
VrRGD4kix9v+IPv+NCYzzm87SaAO2bELxOU8suoYiWJ7HI3VVm73kpD2CR3ycdnO
Y3wf2E74I3le3hG5g56DiQBSDvLdR4p8HEmgIkhOvr6Y8YNJs8lmxXrYFuhalquv
PBnzkPxtYgRALc3YLZxrtBRlgu7SJQcjBvMjclptYdcYbREDs1x+Y9HhK08M/Krp
16Pa5t69jk5C56YY8SgkF7Nd6p6JiZqxta+ky7A1nyD+UUNx+uSHIXRDu1AKSqjw
2qyZUrbL3hzGqHhBN4l887lr7e71Dofg1qFGIzBcaRyU9LbViOyTRGDeSL4oBhof
MMG1iOPj4cO2MbUmcNEER/o6UAUfzy9teR5rtzBCyhFaBdg4ihXDZTfaqb1sO2uf
IoEQ80kt29DkTC8HTRnKh3Y7oAoFJ45KtNF/G+6xbwgPhicwYfE3V0MnDB3RR4Xc
SZwBR6NTd0R520kkdVhAxxeICj+PGSHCjmrfLFH5q8JgI/fpHX0rUDiLBH2hFb6i
Zrf2OXyB+FfxHG8F0PSOtMMwIaDnk0PdOW305aZX4HaJqyYo2J8HHDW6hoQV4iEf
Jaz5Az8AqvnwAXt/hwQhxaGEbfOQdUNE7JU8Z4VyHTmFMAQLTC6bymtb/1sPrPkr
oK9CXtkL2G65ROGrGh2xL7IgXFzo6Um1aRVdvqr512NTleoUKZcuj0jf93HU6SqK
W/Vg8D4yQkcHUCp6kngitJFUQmUJ/a6rsaC9M4xf5da/8fcQF/2ztk2QQtpXgVB8
S7Ic/bZWaYcyJ66j697bQa/rO3plubM+aYFJ/BfCTkXA+jiT+8Hh1cXEQfaM22G9
vhEzc21c6s/T0hgWNx9OPa24tGpU/OpfDXBl8xFng7xEguCViX6UUQkoy1n96dt/
n1kdfMwQHuWJ2X/luCk/aOI4+SVhswwrR9sjtO3sjAZ1AahKc6+cJTFj+SnakcSc
xm9T2CRktO4mNGq5ySwYIwu1mIAfIb/weIzCJ+3O36iKUZENGpaMRp+z6UfHtFDW
W3agafpOPsirJdN8+70t0HfTb9hhYDIOkaZ/3HZX539HXUnV7irxXY1H/GRZ+ZgR
n/zvc/puHLroNfmLLKOmSPMHCTV1L8p6oupT/S8yLWCokIpwF6NtG9S8rSATii8Y
UELgTlyeFAKmuz8QRfqqQHR9/cJROCmK7Igktg4LBpiDYcInRQsshVOq3G6NBoz4
Xxw+48bRLWs5K7F95FlY37qJCQxpZGk3TrLDODNiW98O3PcwsvvdkvSM6ndAZaeh
M0vBckKDu2bimKrAXZNVRz1Iy0JsGWROff/UDujL/QzoXJyYe3WT8lACvfJ2jRXT
UDCbgjMIGL71qvy/+gdVVAzjVl5b0k0l1rOdX+33Z6y8L8omtApAbkMJdBjOzTnV
HzFmK8sZoQKzeegl9qdCbUgMAnVcQzGdFjjUSsvZF0JqckPuukK0oX2i51UC0tAX
FXRYn0iXguYNdfSB3LzeXzgTHvz+zBPFuXfUBUvme5E6wahl2QKNybyDuQH5UGua
xcUjZpb4WjbaHCGpseq//+1ljOcZjjBtUHbpn9p87XWrUPo1IERPGenvdPruCO0v
nvUe0gyR/tu43JHGiXszYcjGxk9tgu3ISpUIHpripaoqeKqGIM20ZA3DrULocdxY
ol/HP8BGvYJbaLKnfpUPNcpUsIeer0TnMpWhBVYu1cKGIS1VUN0SoH5QOZLRS2Gm
k2SFOB2rZkX5+q7SH5yXtNFeGTRcgC6LdyDGoEvrkb4NcumSuFVYltVi/z8a12KW
u0f4bE5kTQQAOCJbKjt7BA8k2dtO9EMhAz+Ko7SDldJWU5sC86B4XPuxSZiQmTZA
qgjW5hrGNY+zW1AvXifCzF12yzXpAFANj3aw7YZqUD9Keqb7We8IKph0/9ggP2kK
wVToLmHHe5t6SAGUPpJ2at610Ebc3YcmPhBp4cTQRYKXgAU7J62Q8CUMtOysNYEv
Z63AS5ewh40VP8LnIp0eNjP/D5tGq8Oz+lDHyrxCgxzYT4qQFSDD20wB1cigo8RB
w6tdqUWl5SeGAaSUql2LQzEIPhey3phUj4NfgmQKx20ZJ0yJgUIi6yAHwh4yC0ZR
PPMdd0gbbajJOhnIygVWtoe7l33Isy+JiTHOtWJWDOO87Nk/djkFWDoG1Fwk8aRA
Q95aBfJihBt3YuOY4xN95ixfOUmuZfuWBDJAN8yNHuXpu18pyehKQWRUA9mRaxFl
uqz1+on8ib2Kc1qERENeXxLKl2ETX5J0+h+BqZpFsDX5z+NIfUUh0EQ94LaCG3k1
2btO1Hu7YyOPMhdxUxVN0cojeIVn7MnrbumT6mTpK1yZ86iVjEoIvY9+6VnntjXX
AwjqS2R3yUBAZTgPAz8Sn5u+R165mDIOgq/xZBJEbbq5dfkkPeoScdV41wACIm8/
dGGvHo/P7rCnCEfzbVeRixZvcndzfRdE7iYhMv5LyvLmy3vXQlR7wd9LnWBFSBEo
Xl3EnujJtD8xDHFUVg+WCEL1JINWoyrbUyso97xxIRjOayA+6cK+RWWg4OyX3Zia
DMPRFFK3ndA6fAHL5Y6E+81yFHgfm5BgxsaaSFFfLDXi1hESP7xjaButGIIrHCI6
NXIjDRBZYSSMrJxRCkzljvj6C0EVn5Er+I5mgVK+QLPXCNG4Zh+2deg8oMLlJV98
k3Vk8JKs20p26G/GnMOHtpJt7yxVtec0SOLQZZ5hpLsD4RZMLBn7auJujqt2Bs2W
9nBDTk5SQcr4v4j4HpTVT59wVEpXoxEcdcPIc4Ox5I9YzyDZ01G1i2OjZrdORJaI
1BUQTiyJvqQvzMIjTcnKBE74cQWln8ZGPhtZ6oGKp5jSzKi8HJd8zMD9KcTJiRFr
8lxDaZ9DxsBIC1xJ3jJvFR+6hKEW1CYNgeYDY2/PDZVli+87FLxYIQEyb0QFmP7+
7jV59gvvpqkdQShjRYjZcO/BMzcwZSk/Hnl8te1vogxLre1bTYptB04jqBuDm5oL
4fJb/0lOhd3CHxzR+0dSx/oQDGBhSESDr6QNhYYHmTEUD7UdavsNvscDwZnWGWkT
BtEOhC5olSgsMIwgDT5DK6BpGmdntZPGW4Bk2/801a9jPbqtP1n6HINqkOIcVMnH
3QstnE8S1DjJSYgjJVkJ4L5wO+9HYGJwZu9aziW3vSzzosMUfeS4DCCkvvDSpMLb
XGVs+HJD/ARL38RBoknf8LToBGmCQhg2qxlVzL8aed0slMCaq+YTjZ2W3PSYg2jQ
/hUwMc9+FoNz6tje12qPCWV5Fr+ntkBBTXuJ9Z82W/zz3Fov8EpfFdnIEL1+LEFS
zVALzsXcrIByA8vGrCLVtX9Wf3KS+C8Xo02FdeciDyt28FwLZc8xz6x8UzvKXSHR
gl0kKSm/efvRzKW50NorOoybGuHBYjyNxjI37dBPSJZOuTJFRrA2dtR8iHYeAlf4
SOOlej84HxsTrCb+l7K+pW06ELq9hN5SNkuipeSU8zH8h4fQtx0v0bkflRE7ot3U
JJCVklxsKTPzGIPAxyj5TNTBksvoDNnuFwOP7XXOa0B8n1hVBeWSS6kurj9P2944
X3ZChZSSfWtkdnPwuoXc1EzIW1M4rq2XRc3n2ZVnAiLTPyC5FWaxMC2ynCdZrYOb
Atv7c8htm2jlqI0XG7A55W+3B1m7vLlMYOSGL39mW4dDwhMybukVefUTHxo6y2aq
REtYaaBAidbbTU5NcWQWHjlxS4wUAX8ZUICzAYXp2btO+tqO38EBUcvk/MrSqAVL
mVwYuc9tvCBE6+/Fomb+Di7/XtODLTdftSAh5Tw/hcybLH44RdkSHX4t4cY3lwEf
Z7FMtjxDbAOd5E1Z9p3JrRJSATpambzB3IyQDlmmeb+s+ZXqsiuILdjn42YwZPMj
BiPlCc97nDxlQ6b1FZM/kvgdtEGrggdAGjnygD0i6TZ7OnHO4XNuQLAM3RdQkv4z
Rm8zceyoQC77pM+xdnIE0yTjIowq0GsTppz8rniKsgpeJ+iSiss+j5zPvpzBoRcD
zGs72NdmY0ABq6h0SPZLZfZUGTr13kNnCSy9rmuSvuG22Vfu+gzaZY0opiV7Q788
4vlNdRymqeKpwcAMKLV8r5w+wy17Qg5Mny8egxfUdSQZq2BSzBcS3KJygoOY2WJd
wt3+5IrKE2Gv2nKZiK27eeMLwqoHWD6hlqMEZbWWdt5yaqYKh3HydIeVKD7cwXaf
1c5MK8GlyNfKVYY+8nir2nbto0oe511yKz3YFZaZDZrJnqbs0P3zskBIaiHqgfFx
LVE38TzItKFGJdgqve6tVqikGuGX90ndvvFpv24+pfqouheThbjXVHxxMAJcF5ln
XKWsrTaUkEuNMRYszeEWbFNYXxS61+0ed7sbjc2+DPIuTrEGE0PwgMPO8DZ0U1TQ
lVGflKu/LYpdmMoA5kUqP5jcUmjGQmAZG1oe8gH50N9lRmbBVjviZ8CTT4D2/cD6
SES7jrEspTECyKwyPn9kIZFG3N4figbM6KrzQQClDiov8nTXlXELHnN64PFC9FqW
/E+bI5kHHzGNp1UyRRjlUG/Y1E8iqHbrfB08f1lOg9wt4us0WS0zHlqTW9/vNR+o
u8eALtKXH3HOKuaCRGrFShZh0r7dYeBQdfWHptHtZvxLYCmFeHy0rT3sd80qa1qJ
CfxqMWsP9O93boRihMfNPk/UPKvQtdG7JycT+kHfAWq4Dz9kdwLJ3/Zr0Zruq0OL
J4WTRd1NZsPaL/CrzYw/GRiqqD+suIqRTb2W2moen1OEd7242i6rVcGpiLt7gB/G
oLEac3pKJIErRYQuHxk4P8fKgsWNYGAwVmlulb1Av4pV33grp4TcjTZNO1QJaPpe
XUPyjv0hWqgVzSXjLxYPzMQjJZfaXx/CediQ/3sKEIqvnbM7rMulhHDb1o02PiOC
46W5LkSewGUVErZ6MmBqOT5GMn1xuoQ7NPoiF+s/KT+ktHLd4C4C217UvrRIFkuC
WY3YwEyXPErafrCbx2GdJdyjqlGN/wNje/tebcHRqbrBUIpEyLEqYCerY4bLWzYb
1qo9z6u2Bx5yxaNfsQ/Mw1d26F7Vc3zWBvJ1wyErwaZne90jz6pzdow1GG2HGvYt
/O24G0iXTvL0LcPvgZYni/vKuJPEJdpLroqoLgX652MUyuvb3UdjNjAc5Z/0g5nL
Ze3fPYWouOeUQ2/cFvXqhDqxsIZcuAxY3OF7KTvSBwWw6ju60yWMT0/5I3++kGwv
+dcMbPbjuDPMSNbTP6KYFmYJPlKBlqGxCJoijPcd9fF356m1grKiJ1tAMbP8VDn5
HxLzIqXROi4sw2hpyetT9pO/r8bkd+Npo/pmtrXt+kofsn8ci4YQzEO0AX1xIMlf
UUwxx8z9pW/qUn0GAuVjGfFQWC+xE+rsyQ33aC6bj6tDplH5104I4f6CXfoChJRf
d7g0L24JmynYJsFIZ+5rq4itMzRrTndT31P4XmK3Ji/X7Oz01tS+eVUTMbBixu0O
AcGXMnvaQXqj/lEE9dn2ZQYIRlOsXFBh3iRGm5FN5NamdAgmlEqETdzzUAVlfrwC
czEIbPhplUktScvdmULfn0kcwk/0P6HH1LP1Nhq8969TEImdKmTXGix97ETO8xHF
MC9uH3s3gI1jo5ccDYC+n4j451vpzft4t4Z+4bxO9p3JKO1hJ3FD+SrXEdZrvuG3
EpmtT8YLM+4+IrpNiHb9BBevQPEhOOA3dq52UPTfAv9PSy4SKYFRRxpBOWjuUc1Z
7MhMHSS3bnmvO9gErxeuj7BULQdS5/d4yPVpRLaggCQXOZ19nCRuU/uqe3oB26Al
hKt9WtIdscjFcOKf5PPqjIJNG+fsY3DzZBL5Qul9BFTYE94WmF2oa0UwiOAfvuh3
Fn4+uRoRpvRXMwL7XICOCgcSrVl1RrImBJQj+5QFdq4mIqbS9PVBzqhAjUbLZ9EF
6O79HfcKohkk5j0TFBXoDJXZ3PlKvPD+6bnIeQQwMIcdbHYqLnIS7Psg8Iz0LRmI
zjxtLQS1l9c+PywT3GzisUkltfcGKo9D2OOVnail0Wb5GucOQPJ1gL9qCi1kssq0
ui3kwB4l3D/xIsEETXKQVedBPzOs60F26Nsky/0zT2O5JTTI1SkKMEVbCqow7DT5
0CadbaatuXiMvA6ByMOz0qbI8MzW//zTW46LDpymsLOD4MDwD2fY5NMp4vWqYRIo
Qqta+052Zb4hxUZeow/sBTLz5NG62vOUu2gpAJ0A7gHx/IqsTEypm+l4ANKSQYGL
ReMAws4mugiTpePLB4yzePTefaum3QZfqFHA303t72ceeiI52bCp/7FwiiRqnQK6
CdakAib8MdWg4Tt15bmsf2WYSKY0HcH3DZ7JVyLpDmDPdRTtrqHWel7cUAC4jYPe
ohea2pdMjYSWRqLRyEKn8Ko/vuJr7zkus4q/YgynwIMUSigfAn30VuZ8JoaoGJ7r
/cKujz4rYr9zBdpcPSicKfwdp1fZXXlpJGifmyUVDTbF16WGNsK/7JKLUl3FEbnt
Tjti8NecmXDuCKUfbjc+v7jzOzArg7Za7J0qtqTY/WM1VNck6ynz6FJ92KPm+8gl
CkTDpZb1DyDkCl4QsN/pihkXYORhdqJuffb1oY8efU61xPdQGVPJgqd8sA3/k7en
G9ay7G2fJKihsmQJ5+YcyBwDvyLT51Tr5j3HjbX0e+w2ebxGX3Glh7TmwfceT7yn
OrkHsQxJ5l1tT/ysioJ0ShVOzbDohdLlBqhgBdGMJx3X5Gtv6QOZGCOW5yi2mzXY
mudeyb1Bpfxz13OzJnWR+8v1AFyt6sv2hgXf2oBKYvlOusbpcMf+Q9KR0EajFF+M
W/isj8hdEmQKaXNLv2WK8RO2DBjIhmS/Ujs495/ICzXfXe4xN30LmOI63X3R46aW
aMRDdv/B7oMzO1xv5HW9hSih7Uz+1lRrGc+Mp5gBpkET3M/HBlzL8wEReWod0wTx
pn+UfEI7cGGFztWtxCac4/b7fWyS9/wbio3bJjHP7w8TZOYxFTzDQFS5tAbJ+LDe
3jhvGyIqJlE1QWX5uwvHUFTUm4FQcNMKhlfei2UJr8gsxvOmSZk3lT1uuBBh97Pa
cnkEACEScMBdMNW6Yr+d8nMz/NaSRHuRRZ5uefp3ntt6emMUiBfVvaM62r+ZWqNd
HQgxXPJXN0olgzuPqNbmeC9pgJC6fLPh++ynhE1CC37uwfnsJa4pBKO36LM2mg9g
OXyS+rYFBQaAFCBdOD+zQU1t7xZGeOxQGAk/93Egt5EXoXre9Hi8ivnJQLLlaKtc
8Ntqcj/TxfUx8zHQZqTmpzK5MTqGyc5ULQsbjTR6qQ9DQQsN0svwXIuqEB5X+OiB
HDSjtMi5HS+usdHJCU2Sdqchoc66N6orPSiVdR4GamExJn+mvk4/l9PuX+B4W9so
i/H+GEMX1BDMeLkS0U36M1xjMPQEhE9cj+ubkY6XvfiP52kDKQMbHJWEQrZ0lluO
qD5YyiRPgngbpWkikvysSWeileSVU+5dAnadRcOyo5+pTTLBzwd27WkmzXin1pOs
CsZryqp4F6IcruXza1FWVw/2k15VEOGLn/I/olUhm5cjbusk3/kQNy0T0QVgdi3o
15bA1L+YIG8NvpWGCENXBviHBQLwCiCN90YfYQ9EDk8VM4CHuAuxQ3aojCJG90+d
eohpJvr51XqN49ZxGSAxx64RFZZZCCAjofT3FFmanDXhoNO3qKyx2lhcEmOfArUu
FddL+Jz14L4EX3ZRQ1aOVzv28l4Wt6P94u8lrZ6Zcqhdw0Tmw/0ynxV3qthzGD/e
cs5o70kRVV1MHFQ2oB22LfUUbWpXLUDTqsXkwKi4OHAwda5h/6gw4xkF/he7iU2Z
F89Dkg4rEpYfbFNtTUcUFqxJukXR2SUpwejmuIcw+68j6xafv30NBoPqlN1rSfiP
XY1ScQGMqXXRfhzQMIF1135XvGgwOORqMj3hf2hHGf1BOCiSscN3V9GalyfYgbXT
84CvrCyELzZIQ8+NOfjeCxoSolFT45MTRFv1Z/j51Q3T2fgcbqLjJj7jY5aDRVl1
0pv8msQapNzGkik+ZIaaSZK5w88RHqh0ZDINYNqFaAyXOMC1lfjY+YRcx3oFue+4
+/NLMOXnm/Clcl9N7eseNb24UEZqG/fcpNhqJMglcEP6duebhqwFeqY9dh8PkIk9
/RUkSV66yPEx4zRUd94dZr21Vxdj4FV0rKjNggvE71a/mRJ9l/O3WN2LmkMXJ69w
xMfWmLGfsB+x95/QqpBmMO3ETX6vJQMvHX3zX/otfyd3I/E2TN6XASDkqC5cz0m3
N7NDOaS2LSG3adhggsoj+Mp/SCeQxbott+K7Nz4/KR3hqhH0+D0VXiNXyLYHv86s
R9p0bw6IOBqg704Yus8k3t0V1wZ7+EiC5zBxj5Xx8FRdgxs3XP4YnBqWlMCs3PE4
hI8ocXlf7dFQq/EsDxfaptukhFIM5elZ59i03OkuOIc9mdB/CM6AvoDoXNwDb2Vj
2OGmBsqaZRV51LQhzmRlgWzP5Sp0JlXzZ5bOTHQQuJOS3CQXVUXvVeIkoa3BV/oa
p7fnMEkV4w1NUiWyyPjUqM6VaDHQiWflOTMrZM8zY4Ztm5DJmkN86f0VQT71ym9l
tnFQyevlMtMveTeWCX96Frvp59wlYAuYS7MpI+arOY9+1dQ8OgFYyN1STv85LpWH
jJ9+8NxKa2YBZkR7yj+r8Mj+/z2Su+zopngBx7cGABiq0uRT7hVQ2Sd0NeDeVJ9Q
t1RsQaSE6F9Uy8tTJnOJO1fN1B5/VAEwso+IphNRXfAUdpHo4pWHhDO31AVCAVK7
eXnTamhhNuLA/0mV++H0KSRGzo/neOUruRX9eI09SNBpNksr6ZEY9F2fObfwPaL6
uBZINJ0WfLX2YcV0lA7qJ8zaeEghKkyeDFH0DdhIQkJktmfyvnwqZhjCn6oD4frG
86oSl5/kpNZbPQ1M3L63e6mgHB2PBkfXYCXQUszIHpNeNM7TlwQs9T9EupByDXPN
L0wJ5d2C09cpokBrYJAn0lIJ1QSTwHDuUwkkbWmt04vwWAUfItOa8pSvxLitcmaA
v12M7VNEV028HTxKD4C0lfS4nsGbvZAjl/CLb0FGNA7vMq5vW3TDGQ9g/jEWRycH
9cU2KBsU2JIb9XXVvkMfTpX+8kO2eyNr6iPa1JZ4d2PNuN6d+WPG+IuKj5oC2hle
4RsA5GPVPxh2IfaTQqTht4lvWSldOx6uJkipVqDHXVPXskQoZrik07EH3J14nqOV
TXXBXvOwZEgvz/ELi17hDWhM7XUZaNtFScH3wy4g3E9lVuzPtVx5Ib+K+kjB+dAK
yZYTzRZsuKRIqCLLfr69RcYMNzfC/n3ygW7xaj9bk05Y+PZ226AcKfNhbM3GhhXG
4QvVmmJsOtCcmPHxPq8ryPuslwFsSLgrMguwwGBdHyVcERt9jBshKmND0VL5zjpA
JtRhIQo0LeWuGGz10bBYIJrEuQqd1RhDm1mmJcnDVoC4/b13b9m9vk5Ncy/p3g1E
lu2NbUt78lD0hD1qJXlx+zs0pkIBeKd3JLciAv9f7HxrLTmfSUOGWLjptiuJnvk3
J5sPSDkTiIBY088NDyU9UppCgdDDnOLSeNv8T9uoO2a9pCaTUj1dn6/EmAQDIGtf
uVQOKMj22S2ql/n1pt2T+1u90wWIG03nZQQuXueFmtOzoq314azzQH5g5J70MPnm
zxt28awFhgo7+XljApdYHb6PNZpSIoyYQfLJ/gNGuBf9RYAFZGfm6XbV8lCJGd+k
wFQeimES6vQiMhXSCgwvsX7v/+zYW6E9eZPXVgABVVg+A7q4Q0U8WVrN0IMlKuAV
bUo5rQept7bA7/RzY4fIgENQSQQgD4QI81/gowMDLgCh35uoQ2omKUxJuebaR9qy
TktFsFbIPvqwetAvAArpO2Dj6m1bLKtjFRJihVuyWvB9unAPXBFiOFe6kWByWiRu
C468IiHYZHHgKq7GzA9IkU0dJURV6UL8trBxIfpkmpEbpS1ihLf01F1zy54KhMux
vEtwOD/oSLDJcNzkYMmTphrB/FvLOYZp6wjmfLt3/iT2ByECBEWXOyX89f7BImv2
PtZDkg2pUGzxBRsywX1mE6T3togNNyzmTvlO5E2QFPo+LCIsw6QbyU4bSGSgiGWb
afEJKPosnvbHvzUirR7iUzPdVws/Iz4DMFC+FCpLfkYRjezik93T97NgZsfaj3B2
TpyxJyEvU1vv2lAmeTISPX55x5fMns4NPpqcxyFw5QED0lse97TINZpe/k+tkcNH
FaRxz2Bl0nri1I/rAd8rKWHOLOBMTBwRKvc1GYmFFlSMgSD2dk13n6OrIB7WCjcn
MX+6a+8qu4iKA4hiQNGADoQAtd6Z+WIqRYEHxKHOTld6tTWHZfgvFZzBlW2DTOgv
Veq0pOpuOsZWWMEk+ZBMhHLUVvYoXPsiOLjwQhyBdw5IC/jDBQAYMoj5Po21iTZl
Q+8uashhwoZR3SD4mEhVAeQ7UOJfPkMQlI+w6gU+2S6lec5+sRhyAcvIZjw/y5IM
bsp8HnRttJG55m90+lSmT91+uxoG6KD0CaKIfoOOfBn83kFroFDZmufAObYXJkPU
DfOwmzIQp5GcL6KetWLpZPZXOrVFLtZF/X20V7059su8rLU+84BFoSaz5T1O7M0a
mjUoa7dwyY+3kVc3x1UkLtvEREEtQfK+JtYwCuQOt+xyNy/GcUEcb64gzhcguwtj
Fgvgln/qVHDkl4oDd4rwwvkLnjsqdovCNXnFceh6hT8iTPGjIje5ekhrY6DkBljM
/4XvODyVtCP7OpI+YYRvkpunrLfTtOIfzpQ2IdR9AYTkDTc4CXeRR2x291oMu7od
RHVZlbQ9xnHszYRE7IPXnKL/i8S+VbRG9sFkB9WRQ3elUaszQsSkaHCRjya+rgsm
0cbk7PqxrUgx/Z5Ufx+65jzX2oSibaiven6pDpDSFUGLqpacD4/KFrC6oEXV4uu3
a2moZ6s3Eb1F3fyBBmZ3Us96XMM9J8MOqvQDzHjLoi10g3gHtjWFHRa8V5J5BsSA
KVES4DZ/+hZf0elhcL2HnYl8UsD5gmKWnlzgYk8miR/e8/JLyrZrUTvdvHgkq8xx
aT3N7sYkd+gpF8JBXvjsV4fkPPLXptYyVaEacz/J2ZAQdFxpEMmPF7Cwm9YOow78
uuZmMRejSN8M3IsntH4iR+JBfiIyG5He5wBNXqKHY+5HBdfl3rqRW1MRkYgDoKHf
HiJ1NWFjtHv53Us7r26YeO+OftcdckeXajyS+z7tR10tFzVtTI1EtBSmrB1bnVMC
qkfvOwWwymESRLbpWzkLlc8MixID05rPG3bGUpAluhKw/gelZDMDLu3YOD1z6HE6
2lb/uIfzoxOYu2MRbBo2WhughjTEE2RlKBXvOuo7KA3bHkm6qjbEWIwPXWrJmBHN
+S2cj+EH6W0vurYO5LKFREAzC8lMnB9FHsZptZuKs68byqf6TJCH8liZUvHookAd
M4shNuPm2VVGEn5Gw6cTEMHNPRsAUwIUEFBvTaZtd2qr4PiHox6X4HUht9g0lmpG
SXyNBbYKxCG0hRS4Vw2QzoSDbwzRPS3Vvttbx4F/hp+RFPvDBAzqnvdkEDQdKQw5
sjSIM/S1fmQm/8VTD4DtbOtf7U9H33VXFlt2HbI5owc9Pj0gcIR6KXd/1EqHfqmJ
ef3Pij8KYB/DjucE8Y43w42eXtDxS4tfR6X9/K5nvXUbSCQp0UrfY3VMDU3/6g1l
EQ03JBHgdq2FupQNfHZvWKbTsFYvVOp+rnIXnB/nDuBTmMZxifwOSZSAgZy8fqJp
vS/WLnW6Rkbh0Z3Do0EfUZrr01lRCQysIj3auH+2Ql6znSHRBMe1jJAUUmjYJSTu
8bj4SjE95LUVft2mI4r1JIBytJfyJ3sooke537vsMxlt8aMECqjcDesf3VsqHIc6
KwFZ3bax0DK0P/mJa2HETbgcPiCehghve9do5Lqmgwg1AICGWePz2Q6aQXTdQ/eL
SmCh4kC9CcamZJWU4L6R1pyhVqDwiHhOX9Q0/vO8uXjq21G51RDNcUscmHQ1t+AW
1IDU4LOOuCqFUj0vuwE8NKt9IEkOJcevbj1UQPsxWd5vxUSFxhFx/XZDnhpH45gs
3P6gKDLbXUjpemU6O/GKrpnzf919CIkDxPcINdPT7Rr2vSb4zwjQRiOXrBD65ONy
711xAUo7U85MP4r4pjWd0M5QqETT94G9igXWQpH/yxvXsyzyy1k5QPk/hajQubsT
s51pRSKsA2cSxtMD05fI2DElDjzV+iVxn8nk2A5211/SHJWZ0+9n25Re//gI481A
JEcVYvldnUwAtFDxDz9fdM555h4SoO37mkk6jXZQbv9QwPQexLt1Vx36Y7CC8jiU
nB8zF897Y+lVbLPwMDOgNRDzhgEyMn4GIMDhRBs/p6/p6HAIN6QrQKjWMpva0l3S
NX06ZyM3CnSMsD8Euz3fDTGC7pJHBce0Atq1i7Lx6i6Zdl+ulhhoDhwc61jTqCYP
8jbWPzkjVxxAWnNns5ti577avjXCq866NRGlHSyBogGj+aEHIwMCJh3/pA1q9vuU
Z7ER//k7F8bHoRlogjcxm0iY8CEnvOV3LM4/sudcNA6qlz/989aOF4G8il3uNISX
y4UNFcj/9TjWNi7bcLeh06gjAgUv7mC1kZnFcQY7LzPd94wUKdg3iVkDfo3uQxbl
NQB7yLWwxJZgutjDdI3AMuz8SiXkHpDPoGa7ppTJCfCZX13ns5e7R0kPPUmEA8N0
0S2KQFQNC6jEVntG6vyS8Zey5dpUEn9TH0KiOofukeShTR1HOodH46xuQLKrrQNZ
M5QOrFuu+ZnJQDp/xvbhmlycGlrobAk8YA27oW86j0Jc046HUVXoaCxUjQFNz033
/2UGBdeVlWc2rnn/m+hAfujZMUwZBFoJJudwwsXJV4iAp6kz6mnV0mQYJgX+TOW/
qMIVcPRhyupVulHMb3gO153r5J4UQL62UlkG8CU/6pU2jIYz5of+KCrxUydy/At1
IyFK8t5geVaAYQS6iBKuGMzayJFy0HIsLFzvEm4Xp25M9iDuucOf6rTG0510/Mld
QLCJ7IvpY+PdQKZfEgIEL/vQdUHOE5Cp7liygn9SoPoHw2qQmMyDDrDLC69CMzPl
m4a5LUsBnZA7SFl3T4dAlzZhWMovipzshOd+1XgOudtxkUvcaxHyHBIEgpq15gCK
MGEqN/DkGWgKeWlx3lP7ySVtODLmqv0iuV+UUWE+ClizTlYfKeFpmS5fTgRkfoZm
sg7CdfhXyA50cCayP5ZIGFRUZJr/92FOz7v+dr3H+UHn2EMYcIb7smqNy/sJfGLp
GuH+SQB77EbwbS2GiCKjSNBDSFKssvuJW0ULL+sJTJ7MumwqS3tASnz9FFwQ1eCH
zToVaD2hGb2pup0F4SeDGeKn6SdMyplg7i5qi7WvIg4HBiyVv/EFdSFBVs+3wHs0
xaR7sUJ3W+fCvWoQuMp7wfOB4uZS3wsDP8s6YDjmMA2LwJP2UtcwY0R/VBKmSxvu
9K1Wna4sbkKuu/F4JQr8oRqBZToaZ2OTVFlBDZf3s1HJMdZhiqzOAnN+sFNN/qf9
ea4mWgtUd3IQ5Lvt15yZa94pRaqJ6aS6C/IhjzqpWF8gaVStKezkuiUJqaLdXj7A
2MXfmJhAtOZW3xpQysCY8voglDOXxQfL9jpAqb1j7j8rKdtPcLvNvUHcftjLWf2B
Plqh7mpoB+Kkkp140azvINjyOnaq8Z+FGQssr3L7DTrwbzaMbwoLCfVxNwvY4ts1
ceqP3MT+Ql+Eo6BCkNL5hhRyV+B7731ES3tbyQIGks4Si4xqmOw1UQzDeppY1b91
Sushzhxt8wK4HSQXzUWfxd18KrkdUoG43N/XPwuWQw28ooKujCNsuIhDNUu3EALf
HoGvErFj9Y827gZgkvOayoJqEdgaF5TG/p4RiGSeDN6CCymLtTS0RUqKZoaWYsHW
BMUe+e0I8VGrh32ShxQtSbDEPbzBFJHeooHi4KLDsB1kQ0R/7efljzlPZKhCTAck
juAeibzZgGwH8SzME6ZY5aVwL1DGHXJnHinUBlm5TyOnEFVu5pyph4/DcPaF+uGn
TarJmB5Okz9g24YZwjtn0A4UfXbk8GrUS1gzTYTRzABy1iYvaSls0qJbxmILMzFy
K95thZ6JLAjfsl1NTqrxi58ab4VPz0W6BUOS3SN8PtnM6Dmf2kHc1nkwOMDpVfSz
66xzg02BxLNY2e0FPCSMcVy+ziGoU8ln7tRT7Kj68AK/FNEV7jyYhwq+hkpf8vFE
kWDeKhms6VD3p1Z8W1v4c48C5gro52yEJbxOe49SmkKD9o7aA+PctnsS065gfBdO
Lgq8a/lv6x6d1SXxswmCCcfiDfFPAn8loY/CLDAnMd+lvGypm8AEDCMIwtL4+CYq
wLVNDr+VOrcBbCK4gkudZwys+d/qWYqMqSuyoIuPwVLyWv5x3SN70H/tCc7Wxy23
c5QgbxHr4wD63HqIAF3CxmZVDoMo/pKGIBBRLqnJN5EVDoOpNOTqjs9KCl7M5PZ3
VM9WoeMxX5meHTJPoAcXpPNTLddHo9856N94E12+RP8Jsq1XrBzD5I+qvoArQ38J
QX9F/iMtNPfoJPBmNE670upI4pymwlESfIIwRqgdjLDtSQwNygQ7HIYH2S7yj0Eh
N7PTcZChhTcLMjFN2IxKqBQExYO9Wu0Yvico4YcIqDDbE12OGYJaUoZePG269gia
FGM+Unn0zpoht1ymkBHygqstPrP0MiSAA6Ii8/tjY6VHE5Rvk81gFVarYCeSaH+O
TrTc+lp0vE9cFU/qSdYNTFfqR3r00OVbgpGZMVtColO1KaUkRMUigxjMONPaOLe+
qvUCKtEf0co3TelHl2PsHr07E4ONik2bfP1e2Us6jYABjDZiwea3YwqagA+aQ9XY
6MOz6KIwfRELK0ZwrxtG2oosP5Kk9U1nTgRYbk397nfOr+M0dR+xJZ3P9gjgL8K+
m3VT3DsqNJc4v5Hl4WnKguH01XATmuU0y+j2uqXyr3fd+VsjHUgwU6/6ruB6w2uO
Ks0FzQ7z+8PITx+3p7EwaxQkSrrDsxdGeBxIdPH7IpU1nG0gBb733Uwfv49GG13E
UbxJ9x4SX8gww6/jvt9IRcX9Sm9R4tXxQ7RsKsDDMq60VuoO77Kvfn2MzR6b4oym
hBFhuoroZt/d404aDJPQdYdGuN2Af1Tp3LCgAOO9t24cjAxok78MLSZXvNHxgAw9
w4NLHticAZ754fcNCYNQVyACz9jq24mKe+/giDNesF/RXt8fA4FHfxNKf2ey2cqZ
LCsoUC3OiOn8jea5jPt9XwExmll2ErLutmE60Mg7d7FRxtSWrPvWq9XyRCRkLPCb
6CDokJW1lR0dC77bLXJFQtHmd94j6VLXFsSvKyDLv3EqKL4/JHQS/+7zCLdvR/fc
dLtG8v74pDdFN8YgTiXk+7r6gwyEDvsKt807VjJMiHJEZA3B9QUVgiZeD3E3NQBv
m48V1i4s5zofSqtBnPjFaPP2jnlYz24glRfVfkFggD0FUTLUIVfuMQHyHnEjRF9X
Ebuhac9qDfeMSHzGs6YZlORWArbse9MPjXcd/JO8TGkyM6Nr9rNa1mRBiXL7xnlY
b3/asv0WrGNTS8Q0Gihkt3LLRXv6ot7AqwuOw0tX/g3UYrYYT6LZYy8+Fg1kD2uZ
TECa483teSHkqSQ+i+mDczOxjzhlYxAPitvQZqBghUGJI0wlux27jMqM9hqGFdTw
0DkUI28JRsjL4Lhsx5iHZ/tPg5MKN1/WgVJPXclLOAxBL4KAmWtJCYMasNF+jZir
5wkSZaTeEdzYJXVRFoq8UCWBFjHJpAfINV+RruZxMyUkpEbmoBdjTfbtFqZ8/9+g
WcT7tkr+1E3Em2RSRTypNKD/+KEUgyA5ETmpgxBNrzGRifPoBysOLQDfIX0PDIWK
jirY6HiwGhF1rs4bKrSn43JQLeysrUiSllIioHhp+FhBoRfi5YkAOq92fQEDpeX0
bnzVOyiMrlM9OiFU2Bovyy8eVdoBFi5j1X4s8o0ZJSFzkHMa5If96+ml38mvu2kN
LgUw3wn1RcQtye0tCBFhQv0N7idy53Lu1LqCL4RWEeKisK+nl0Gsu71Bgtm5Hq1V
Ilw1Bku8DnVFm/3B560JkR4nGfZU19E0JQFO/fJl2dU4gxdxsmzcYN6m4RSE5FaZ
1yfiC731uT5eYJWZXDS6Ea8B5z7KYm+Y2Kroyln1KNuWCqJVYZTf7L3FjyJYBoFc
VjbLn7300vtwtiQHwENfHmY8AEmXZExuVdX7p54aybm8yGAOtckpqHEjcPS/5OH5
axMt/feiM++Yh9wyCHlPRI116RAt9PD8NLI1jxprk387/5gZXjqkhPdicnWFWFiT
M637sNoLx5YMMpqJBQ12R7Q25bjREN9ppt0nAJWHuBrKGrqWchVqmINQd9bRMoIQ
dMA1G9J+clJPhq325ef+pum+U8asHySdlb5pH1Hyc/eQU9maKZk0BadBVoZ8X/D7
FFQPPK4LEHqMUFCvxqlYTjEuuoJy8Pp10/1yqoDHF8NvAZ5pAbOzTn2srvpt2PnR
/MXNe1XIAviRnWTnngp9x5h9ytPYGjK7ZAAZ98qiAPkVE9zFlV0s7Zkf1KjogRmF
FhfpKFBd6fApIRkLOA+O5oE99McMcJx/+JodJkb6w+tvqHHwgTLW2dByGB1czA6J
uD9hlVCfLKS/YHwcxcO2cW9hVzT24gikhs4GSOQ3unuA5VxE+SAUHgqdFOiuIifk
r9s5Ekss6lJQHSWGjzqegz31/wrlI8+X/4s1jy6Jkng/BL4FfaXWZUjo1L3AyXuC
2Srkdr1w3jhAf9YtlDVyG4yzmQ0hgX6HxE54NtmwBbpmdePQSm4bxB6G+82WqYmg
v2Ptwyuox/+NkKj2kl0lZ52Hz+Kgh4dalHX7vXsxvAF6FggW3F7fa4vtIfK1lJpk
qSI3R3vsSKsWUY7o45rNVhQtBCjiTmx8AmImWba8+4WSg2bhj5RoMZb01RmI7LAv
opSoow/wiRTMl0oUEJLjFcthJJ+6/sqT90WudHCVZkZziZ64rb3u8+VR+HDeHdDC
LxT8WzC9exJVGhaOmLfUEKhT87wXFJH2ZfgRa6Zk5JVuwPSh/PLiRas8VWHbpZRd
Zqtiw8FVUMixEQsYfZc4Q6Fe6ZkLrrLVgdtOJcTrP4fhbRg/N2xafdIm8c6MAwxT
dtyR7vzKkGvxEODKzOlFbPewcYzF/hH5EdL7NfI0xT9ZrgnkJg7eo7Jy6o8Rv6u2
bIcXvpIOQX/WejaZW6NzO5DHbJqdQfQHFNkd6qgAaXaGRM63DXP0Oa1KX1oJmDUR
xmtqnQ0plOltEwr2h7AMFUrYNC3EiF63ZxhzUGbaXRa2MGIq99katyBGjvtPYWwW
KvjHzOfcgBZXj8PKGl9AtiX9msNhDNkuePPPm+WBjTT5krXtjjZJMOEA+cK4JsHG
BreGn/v8xaGurNn4lstBipx61Fk7F9Ar15vEGMBzmAf1xVOTEroer/X6hEQluyth
tOAlTY6pNeq1Bk+uynNauTxOhk+oGdNjfiIoEzHxqiqs7XX+JCsRHVvdRG2EYemE
QDbRF4bpJp/j0pE/Ejgsz3w5BoZ7UbRtKN5TxEV0/qBBTG17/Q9KVFrhWquip/ih
QnGwFl4vgf6aAXBnpWxsOSLw/dANjH2dn4fqy95SWuf80G/cpBkCogRkpYEw0+Si
8axH2rgE8+tWIJ31bAp9s9nCs8jVI9tjXjCHQVfmSUM60exurROoI67vdihcSrPB
T0DZfeYaQlFOHxMWftXUPvGIYzhxfn4VzlzN35zBsrC/nZ3wvMPgIVK5PStKTTdO
O79NlYG+SmE46NsuJx+GEQrlb4EH300KdT1/wMocYNRLHW2F4hhXAF8fczvf5bJg
Y19hH2lGyVIbU50bk0805irEWLJicK7A6hpdtznghYzjNBw7/cDX1woYlRqkpFD8
mh0tqsBAzi8rrS3r+C0y7+jQAa6uwR5cQMAjuaghZpPYhmGTuXwyee0EUgnfsXQE
QhmDd1AZ9V3gjjxv4cwhBLD9WKnk7XMV2crEKgi0D0O1FNKn4jlri/gi2nnvGILf
ppuWAqWNCtuMomQcRKd9en0Vy/3gyPXE5TOYu7Com2xgjMoWxScEqfCt49IqcKY1
EvTJvaWe/qjnLL1RDVABqXL8xiBp2avtSKysffpTnVZWWvjbmq5WQmMlWKUV1WqL
RY4526D6nIXuzVV+uoEwi6cIYEeVJHxMY47VolaNMfWtN4sSJNA4Nw9p96x0SmHV
Th2adPQhhBvFPFY20KAsCOaC4i3zOr1n9E2P651l8MT12Qgi8gSX+af8x7+tApDF
wJMjIWNiMwdHEPhJcaGvqQCjoDjSelCIBEGNRinQ18xXPcvPOY2KVSwtE5W864XH
uQ/XcAchnKpMsVZ+Q8aqJbvlXimOt5LelY8RgP5PtY7IDztp8OYVyTYIX1jjJk9E
BPO/KhfX73ANcNk4n+cpF8jMG285lkHaiZvfbwLrFJwd/mwe60GDqbIZ4FKBkb3w
wYSqaas82YzsgCc3pY5PXFLqRrhOoH2JamSRiFZfBERVi1e1bsH+T27yEScbjlgp
RQ0e96dvViI36Qw3vdZktn7vJmRmE1tgeDb5qS/LrTuZGVtCa8S3Z410V8Vx8XZQ
acNY9tzRcE17zunYna2kksiJDK25tsik67rOiqdtdsXHsULqoBqKqSIReIYT+PTk
hR1Zj6fZNpBdw+3zdFlmuRTIXS7k7Q/e1Pl27I5hZrOFcLxJkcOlAuwQn/y6AteH
Ul262f42hrXQErh4Yxi8zfB572Pib+SwLjjVuA6jZFB69mJ/WxijTAK5HTm+YJj5
6uJ7nSan1KEyoN5EjSWy6YO/RHMakRGAc+F5djKmOlIGTbLc+bA8gWtywUmCvo9+
uEFhrPzb3ia41lpirg6yfsoRkAa/L7+9DAb95OtYzkXsr18Te9RG+r4ET5sp0HFd
ljg5k4VLAZBCmzku/FtimpW0yXxy1CnvO1+2rxyxRAz2bZ2WtwS0Vul1we9tFAC0
ivVKrx9o283Fed8timQ70UGt2/TRjgVBqP7mZQQdCzzkFokMGEVQ/8QnSMOw2cjW
7wMIIcT/mT7B7iFasqDfUPQV2A7JxuBOiTQ6REai/2EvOrtiQd+Mg6bK+ifdWmBb
jGQUEmU12BkocBFG4J0oBNmqYMA7aK25KXNAQUqu/mx5P+MFy9AImiJjxXDor3Hs
APf4dO8cdGj3RB6YN64F8ZQyT/J1jUbrpAkxzAx003DHA42REeRWDLslw5VMAL6U
sjnbpgkCzVOuI9oS5aiSjjpRUexFRNWUCi5rnmQFRsjTuxOUIXvBfNvQ+h4wwfCp
1XEBOocQTrMNy3JLdH5wnIisFfhvwJ7pglgsgzsEre+wK2+b8oi7n6OKVY0bf9Oy
/d1IrPHvv5dYVqt3F18rrZHFDexUdQwRpbLQ70VYpWASycFo1Q0VF8ck5tIlUjoL
UxLKFuaOrS/XiwPoalWtPBuztyfNrvROCX8f7mkUjXLelsy9MNvzFHLe1qY+h36O
KyyyS8xUsuseq0v2kO97Ffl7l+xZ/5Yw24NY5Iq/DrWhUcKvgi7WGGBNyDkpfW5k
ducowcg9oi5/25sfL9E/Pd8X9ads5vLYhzbMxdJ8BsEvvmj/zK+/mK4wLR1Vh7S4
fih1Au26rpkgB069Pu1H/MpzoS6QWJUo67YHK6lAEfD/QQU6fPcCIOZ5hPB+96gJ
i/IBP0ytbFj+dlip/+luyV1KZ299FU9P3ZD9vVDMN1BIDjw8tRFbxhQJ7c1i4VSw
TDdRg4fGNYBXD7jrFFjvdBA0jy32GDWTiaDM2V/2gy04y6evVzLJXdx+pNXpYsy3
WyKfcZHb7nyzLlM4nJhjv6iRVCPQ2ULgpfcwNbPg+YQ2Og/KkdbVn44/wT13l/pL
SdSH6aRko9DdDEdSbvOUSpIrpv60WSS2tZdp1IN3asp7PEF2jTnwE9E5WB0L2eQu
lh0L8BsAZTjQNmB5Mw/K0+wmVGzdD8TB6rFcbAtvzhx5VZ2eAmo77fiM6IHIlKd5
Wis6YliVPR67Q7rn3dHsQdJEC7tw1ryc/QzmKz9HFGPn3qr+Acd+B37JdTGnkAVi
2ZqeR820ezREYdyX3AAPyYKN6WhhZ/oUv9A6CzPI3f3j9tAvVOXqS03/bz8nn2ix
xSYizNIWyYR3kWqUiR8nx/atEVA3D+HP4YpISswg3l3l+Me0y+84NQHXyUoHqpQS
7evgLiEbezTqaDJ3pHUWSrc8akQt7J0MavvgIo/zoDYQLQwdRFtEYar8Fly+Q+/R
6fSebMe+zHJsN63nE1xGPg==
`protect end_protected