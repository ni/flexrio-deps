`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 34752 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
gjQxfoUVC1+c91Q8h6upBt6MO40asmyzYjt6VzGWHBbwm7lJ9Lhol80B+zuKYBmN
mcYXsC6GTMui+6I97KVF5Gvt4jM9DzHYcXhJYGKlSZ1LFuAbBoP70HctjPVDs1uU
K8OsbS55VyhEjKn15xiIvtXli8aGjXHeX/rfWqMfS42YUCbSyppgEsJODINwwOzz
1qRUUw2/jptV19c5D/Bb6RJm+DD1WPAcwpMfK9yt4tt5yY7aldrWUkuXKybQ3RoV
uy4U+pYfr3W/CkV2CFVLeksjTXHWQavgyk9MpfadikRr7Bbvpb8mmj9vgqfXNirU
FuwWU4CEB7Lj3xKCC5lz0AOsenn427PLgbpm5lFI7Vt8g1d76B01xjieSo9wQdsY
fy6xg7fPnBWhH93HJKW6laKa7uA5pPRIFnR8N6neQujORfa0mBLgPXva1p8X6n3F
/+uOR7CUBSJ4KycOaVs2y6PesbVc+Mc/+abM5Ivjh2XgJGj37Qvi8HySFfyPHwoo
WPADf4Ef0cA42gysrKU+GWwuP9gjduAkuSAig6wvduq4gofglrqhCENzBUIUINIC
o+mzymAtmg9Ko/NRgEPqqsY3E9e1i6Qo6DfY6J9LuZQXm1pRpxnE9atrhsZH4kt1
0bZWTNGYQoLyPNODFhj3SLHkQFax4M+lcTkhmqK2lJ3xiYTrJJMnLwoUGAXIRPOj
Kj9v7LYuadDGcgUpJ9jzYBj7ZfYLOUL7YWM5SJm7lhn4tmA3VcK+GvDBSz24MpfG
f4PhCJZ8DrEfGU5v7xN5ipIER3iQ7tOvfJBG5bUyl32B7JzdThiGHekpIPeSjuUe
g1A+cJr1k5o9HJYsZsG3taOo1C4mhKm0OIMqk/RUxPsyEx9KavytSFtfYr/oBboF
WiOsYQEmy27k2ClZnkTfsfzpO2F4b40zXoS12vf7DxNJP5iTkUGmuSenvyb7/sF+
eo0fT4R7D9RMLmd2PdevrdOMQPwVIB5IhL7tnmtgjtDHKCjOlBBP24O8ii9k/ACC
VyQTPB2eNfAceYUYdbipcU6zdaf9ehrubSxW8UC1Hd5f7CSUQmufGMYdrJ4lEm5G
kaU6Q16ed7oIM9zrWmZJHxPFiieynBGT+A/ONRlCU30htDxDA2d7llF+RSXRkUIM
KonFXSkysG5mV016JFZujiUHUXv3e+5vBFakIhwnyZYQwKvScohCxaQytdyPv+Nv
MgraL7UKXwqgACIRibVLm53JsJ2WlIyYvzMrTRzbso1d+mMGDilwVdzEZOyNVq4L
JqTDJjcsHCkNvQMLd8i3jYBiRqhO63ZyBF7ooOoicRK+Tq/afsRh9E3Ve1VDZjIx
ucli7ybR59rvIt5odT7GHyWfCyHtI8t/OEVo2GXfqurws09cHaziaL+cqDyEPGUR
51/VtiXiwSWss0XCdCeYOKm29bBzJlv56+65ql4E4hDvC2N7DVXCAxC3N7WX7V+i
9gs2YZ7dnCzKRR8t3JNQaB8daJfglY7FkPOkLF7M4qSjlHTu6LQyKPQrgB9Hub8h
fbTCWcftgFLkoUyIhkM7hjSaVUJ+xVkaG/V04pq+iD9HLNo9PM0I+19N7RWmqznG
7rifboZdc4fuOyB/aUoSVquMD+lZjKPo6juEaOm1eJhCLRHYTW4XqzjVZ5A5bvX+
H3aY13f7pbId7d7a2Yuvb2Ynz5dzhc6oAfQyCtJACIxkxcz9ZSinZN3YPKJTyS20
4DRTI4bVpbdVxNy6dIT0jA61pdiV//VNVYdIFYscUBz9x52MZ0ylwIGjncSLHPDa
zddfnpeNm8xgV/ouyE4JWZhumf23Vw+yUZ4taV+Wyld20gDlvIRmIoYw7lsTlJdc
mL7YQjWcqQR4cNvAlLtoLDJoItReMMnK+jdmrUSatayVDhNsuouQ8Y5/VOZkqUWv
rnb6ZATUsHFdSlD37LvGWtt6G9au17eX7jjWYGbUC0ZdyvpxI4tDmy3ti48/AayN
/aBxl+uPnzz7HBFHMeKzoGXaF+7Rd5gLuI03GS7Oh78P2Q9gopgIx9JPN/FVCBuG
4gLn/xUV1DVnXY/hs3Yf/Q8TEN6ixazwMCDLFL8yB47ucqKB9b2yrGLBXij2JG4i
IWFqP4s+JQ0Ckmmg7358n969/rgfXV+1P1VG5bwoUcyIRyedB50klNKVZfhRtBPB
M2shAFoCfK0+r2OuHA6Z996ZuljfvWGilLmflIBipEDPZgHoKPblnOPUW3oBD98y
pNUAx+ompypga3tUfVYqEkuiOFoEemjQ2TWahAC3bVEV0n0jz4j4LXmuVdeutJWW
N5l21cB2d0vIIDvNcITCT3k1NhNH8mJS0eq6hH/WtagDn/bA1qpDd2RgB13CXh6r
NJ3FGC1VLyqaYnqSmWdiXjGxP/2dyg8Gic4MtaHgqlCkSLhmUm4hZfOJG7zF9obv
3vf3hIWjRyZgx+bya/NKlowUy3ZH2hCLPgtbfLxEpwBvqEKYklBRs673/K4T7LG5
Qa1Bz3sMCPKmsMxiUtNPBf26y2VlnyTJCh+gZK9BbqJrw6lJmoYkpqGigjyESOYp
P7HuEmKRoA7JNshvbuMab9c/I9CFLPsP5iFtbYjn+6zT/BCACxU+hohr0rv2JT//
cFiorKuAn/idap+GiCzieK6OUdnUBPVfoOBblpJfHGrczLjsFz19BPjvy5dE8aX1
W/UJ+q6dN7asKRSoN/XEPLaf4zKHf4Nt/bEWBwVjGAwzs9KLwaUEVt27HyYhfIOq
FBGKht+4upzVIErZwB4Ftbb57xuO7IYUnCm3NbVyVhZAtUl09c1Ykp2eI4CsoV/z
4sAOHSGvRUyldNzFRxSrQur1B71o2lNhcaPpy4D7DU27jutDdlTdVhcQPv0Tz+SG
nLh5F+K9lZJO9NxzLqfqGe/t/zO8kHHVHoLhJetrGtJDPm5ybdJn8uFTu5GfazpZ
HjDTHoAvlBhhVLKmBtgHUjOv20AyxibkpbFWegFnSV8EfriuaSavq2HSSMLVT+ic
MtPyuxtUgVM25uTua1rIwTShOMAD9hkfeinq6BAGu/IBZchzRBW3dFl1eedgVGod
TIHHDK7cI2+RnN/bbWgZtMN3qDb3t+uIx+iuKMBke5zNElSB+JreyLzvkZniW6SY
jOspbdYKvzjsQ9kk3pt4G4+7cN4VnqrhLWj4YwkaNAV7J6wt9PnAqcjDGZNURiV6
jHI29x+/sL6G/8PNeFn7qg/w2LEkNZZs0/gnePNgsAmONHB8DIdlCAfw8/4To67F
dX7RNORsOkQr/0g2x4LY3aXBjTULGnfqvm6OFbYP7i8Eeks5lRQbtRkqiAK4winF
esegeIskshJISFNnpQ+Rcb16RKFzz3IexPhfuRPLkQQVkKxujo8Tnfo6VS04hJGx
LjGRwVMB96tMYBkwFtZhBESMbaGJQhKSDPtG696nt8QbtzmY2JLnszxCRCnjdQiX
LmD9VKyKohpa1Fu/V46LoA6+CXhaGcw/SCTsuYYBp/8kJMIJP05QhcTN+baEI0qA
EjCvw+3cEvcg6auA9FVYZDvgnpftHpiYzPyH9ylFNm6b6dRSZDRvYsiBcsOyjmQp
+KS9GrHG/Z/ansVxltR+dn99Ug0YtAhQdDYLHsxyuhxiA6geEbySd2I/JDCDsCl1
tnuE7gGMzu/CyUZ20kY7O3gMtiBH1VAl/wA2pvn7BswN4V2UO/KvOmcDyXezmb0t
UxREvNQTf9du2DPQrB3zDwIohaf/Mb9MtSfoHsKAbT8yHfVgW9DcjCWLFJRH20tl
ib4aWYORZjBEMm79TQwnXnT/2dne135NbtuCl3T2YB46vAtvLniaiegCTEdeJ3ej
sGVXB060JC16z9aoaZ9PrdA5B9nPWslcRqaossT/6yXGGZB4WkmeoGyrrlvOATzw
T2Y71mCCkpWp3sgC6gvp8IXnJvmN6fCA3WDwi73tqMxv9o0KcZsw707L03PRRE1l
jCqQUeCr+HJryMD5a0ex7Yh7qn2MMsz70Y5WyAg2QL4hZgO0TCkXN1KV/StvJK3M
YeFDq+YJBUM2/pdOqIpv5Cr2J5ueWKKNTwTAwMODvKEdxQ2Bb2iVG45QuVk5zntC
1wxlWkyedh+2Q7rlGyRQs8dtyn4qMK9Uu6WO0c+QPxdMtrdSCCRyfSBq41orRZ0R
bvwmgFZsiTYulaQGYegploNoI4fa2kUizwgynyf9Kwc5Q48iZ0UWWHovLMIR5vEO
673pvDYU+2M5GtbdOKQcGfPenlh2pyP7vMmcjUNs4Q9oKx335FuNfGHZNOIDyELB
Z1hkq0pdVM/cHhhUbT6slDmj6bccuGMXwdTpSjh+r+UYFJKcSls4HYxLTP0QPjCP
J+aZmvAIeIvPHv3RBoLebBkQ+8WuhnKUuFpuw4T9maWgatsBTQvP7A1LyZV3zOHk
sy9vnUwEALivicBXPPepN8PEy/qEAAAHmBBzfTQ5iGsKGIvnc8sxA0DvfxfCP5Ry
41k/b0MSbrLGAMSXacIrL5lWZgqy+cOX3+jYyJ0/ZLI3Jc9sza38G9/GQI2ctOBv
b5DjKPEHSFPUB9h//UDdJZU5iVw3gNn2IM77o/mpqN/HA8qtyau1e4Nd8rpxuzQV
CX+o2J5IImYQJ+I0Dki754w6RjZAZ3SODGH6Dfs7g8KpwpQ9co7VuKL3x1DM+eJu
v45/tMcxavIeyK6m9RMYt3rJjG8gz2OvdS23jN9Y1CsS/uCJRe3gohslS6A1yMoT
ZtBB4Xdo1zxBaQ18//jQNJSlBor+yqyTu3w8Vpgot8zhxNzI6ZWhznPiqNKZ1HZ5
68YxiEPapzWCCAKkh2Pa+PXSNLIKPhq+1BZfSqHM/UcLRY6ZPVohWkn5N7MIx59/
zxV8rm3WM+dvzfA/UDMKLhJoIfbLdR/qALOaHSvo7wN4ezl95s5Y0QpA8VU2/7q8
zS9SlykVF+sq1zkGA/Vx9ajwNoK3AX3hYjTGf3OPLgwxdnlRiRE9CIrgCS4NpoUm
shG0YmI7/iNVIBAj1j16X4qwTKOVc5rGRHvPqQs13y08Uu6Xe27pDZGrGp4U4bsb
NnnyA0syKn4Cu1GMBl0PSw4tIAXepvKUTfU6eCPwh9dl2E/BcrmPzGwQ/9yUNhyw
kap154aZsCphToIkxrQjaLwFh18EZBxMPLhHB1tm2jQACCZGwh8A2mz9JLUBJbfO
/gAMnO49MwTdC9MelmGXbiIBxqX4I/hnHOlLp1PY+F1HTWKiqnte8ZVGNLwgRNFv
h6OhyMYG1si6vEBvIiSB4oTiL1SC4Ra9PS5eZJmDD9VcsoEdW99ogXXjBZlwSZBD
k8SMny6h0hPvb1jGbj0CWNFuaW4Xcn+DuuHuuObCGW9H445GwbkT7soOW6AdunU+
Tp919E5Ol0s6A5BmKkimdFqVYhQPWMd5hTEzuefezbuIy+waQKcgZIeO24JF9fsS
hnFQUs9Grusw8fYrhtlT0doT/t6+ewbuoxu4wcVIuju8nu7OptkjFY8eyB9zumf6
NM324EEP8p4/8Rxtv5Gg9gECobCxGhUgNtj3YX1q1CRSxbePfgPzv9nL41Txs6mI
BWvDVr0HFcdXbnNeDss9qx1ingEwT5tCZArV/jfYOyUGp13Sr84VyPJOrrNqRC9A
a+uD+NL+61AGNeldguldXSka4pEoM7JKZYenOrsMWLz9eSqXjtWJ1FeI6QBmwYBN
f3ANCiNh+I+NgNlG6ru8qwGGLREabEK4aVZgcyUjVBBmn1ZvxSOMxspgd/y879S7
v0BjBVSlw6s0MGIDvyuj2FZoeZuR+UxBuhUTYlyNDgLtwqqVcV2ilwzBuvFarigF
P79z1yrXIRatfMmc2aRywdHNsV0ChioOlguSfbydElpLNKK+3+xMZSmo8YtVwi6/
mltacA7xEDoVOosU5H1TA7PC5Tw3vKZiJj/nN3dV6GcIe0qh05EuYx57miyQ1kKg
vfo8vIRS98IzqjXL+N1xQE6Gwhy8DFPXWi6Ys5U95zx3jT50Qyea+s4qmbpSlJ6D
kPQAZCaODYDbtb7HMm2vZPKSJ0gBg36GSEwkvOwa4UX5DVfnoX5dZ/5ehj7DDRDo
mVnKcuvFmqPY9bR4TOFtzfRL7fcc72DKkjC9oNQeetzmjWyG0/uaHP6kK/Rtq3GZ
/OB1Or0rnCbkhch+PVyMDqwb1QNrolgEnBzs0ZSn5hnPSgGnq4Io4hYx9K8RpQ8r
qAnXEbwVdOlq2tDv+uhA3DUV/3mCVwzkiNp7547fFWOAolVS3A5eXR1nXdBm2HZ1
msCNy/bp3brEIaaqMt5gxifN13ZhH4zXlWNyxhFslVLHp4CCPFEbsQGDhVVrlUBy
CXkOa49Rsnrj4CT6X/MD2UvFIaxQNG0WrQk4THw1ZmBkc65pEVmFFT7f8HzJj1gB
2Reakh/Jkmmy1j+G+KyqRdN+uwUTUW5oI+bRtrN5lCAEQq8z7bR5FCKRYvLRsb3u
H2Ia7rEDDR3z0vqBVkIxhHnaH+MTeX5F3UV2tuDZW/ZnErVJV3V+a8Rxci8b3ZMF
zKc2svHUKHXXhUpe0CP0B51HHtHuV6bcYw3f4Tda13iqSiOtK1VogOfJnuG4R9W0
DLU5G4zvT3T34oboO4Q/cdFsURw0OUnW680Or3o/akvvKJaMCIX2xGmQQm92MTM/
1dViNZhfRDqz+baTwkN4Cm6sv93FgiZ1KcytipsoY/cQf11gH9rDmzb/d8qG0Z5y
XDRXA6IQOYjs4o+riwat6wIdOy24L6LKrYh+R6U06C0CZbkEikQTlE6O4sRMoS3M
KSIiqcwynSV11+ll0mH43Reip7DLWRKAvdUyK0+//lu3PZOtBDuN/YHh++lnwb4d
jPKUw3G9+q6zi2PhbijhUMgbieSdQyq1PoiCJ49qnfjQ+34A9woUfvoBRBYVfjN6
o5dZzfKFcqNS2P/XQC+1LRO5R2zV2DhOXPPCsuYkOI/Ycab2giC1ZjgYtMjFeqHf
2j3IDFpp10ocBLwcTibM5iLPZa24OCpIbBja4hryNW6H1WVMOrDsC7eXuBY8X68G
D57W7PRUr93/JK642AuAF+r5PIaEvTb7LyLne2DSLAqyhJ3QHuhjAqSLxQteKikc
2nQ94WUjguwQX7hb2sxACcsS2Bj/7QiYYLb9v1K5PgI2KeCtxAU9sHCslAM5+54H
QBYBu7r9YTtyJLeUmAqvIsyFXPN8y+QovVTU78M25c/fgTXVn4sosymBhogySX57
pDqpc8vieN+NkVufuHVWmt3dfPJNSBivjwcNGZ8hzDQxvKYYCRqmbvnkxaiFQtfp
dvEPt3pALnyVfNpkhR58yUe5pFYrBelzGa+bbV7c3GBymmlWRcWRvLRdCfEsBEUS
AzkIDx399xNMLm8ZIk28BpsJ8jrNx9o6XupDgkvh1X9kS8zVkSeuEO20SqGfAObk
G6kwQhf1gVayMdPcnuSf9+UOq7Xbj9XOV82f7bEEuGPtvGHRyS17MHznarVrJiOO
aT+aPjwrYzeoPT6f8E0p9JqJMQB7Nut7HH7RfxghaICmiaaSOHQ+50bhlee6Au1Z
JZdRTa+Zqa/jBguxXgJF7FoKO6PujU40IVMblIlfT6HAHf4iYvchYFwGaMbzpR4w
nPoLEyc5asjqD4Pot//oBvVg6GrowokUDEQzn2g/NKVlxST6y0fw5cGyXKAPCDVw
OCa5zjGbj/b0twQD2lPan77NIbjxsk6NcRAgpISb3dtZRm+sLZWnuMGDoQkcOdkp
9iEs5aCAXbnOwjFCdmq1ricX/75BlLd4JQhN3BQtBTNhRecVY+EcESjO5mWFK7ui
rF5USxheYkRfaQIqBovzsJBuuzON6RWZcuONoJCtjVKh4Ag94v5DCdKnISWe8bWi
NNlcz+J9BnLovfV71gX81kOHmfn6XMldWIOrh73BQb6LdG9HKZE+VsovI0Y9YZ2z
tRTQq/sN89t/yy8yjyqtLkMtkrqaV0Ys/geQg2SScFkAf4QS3Ap5ICZLitW6qo+h
HQxL/MAdUY2CteeEsQbP3wDGhhhVoK1Rnma6mECIklvy+5Y0YdjWtcLU2TyxQ+cg
xpfTEoXTdKRAUS/CCQmyPRpFATxjAv+5LpcLhvKsejL8S3iblrMMHFLsDP7fGBQj
yGoMx7w+Ma9vtIHvra9WySgkRCOkPs+7VUeZ3sId7gcs1fVtkHY3Hy+gPC187EmD
fcQkhQJWUD5EuJX+y3nFr7RIWa6nKSNmg8TxAgnLNasVpJIt614GTzapuD/6OxLD
G/HczSGM57NhAg0+jxO1so3+vXYEKKCugZ6fUNi4u8lSEYad7eoBtt+DWQgrxfT7
xEOoBytOvt8Q2Kc1vidnSk99jbBL/umbjO9y5/aGLhTuwI7Q1P3c0skyhfcFyS8J
nUGuMpUfjl4qEav9YM/+utbfB9fopEfjK+pfUHjkiOMG3DB1r2enosZNlzV3YgRg
7c5qB0Bjkde7raQ+PI6SFV64zY9qj/je+RfqPK6qFYRsDrhOLL5VeZ0Jmk6VTsdC
37skkJlCRrbVdNTdd8SXr783EgcyaIaWKr0ILYgiNzw2LCJLd1e48bxgaiI2kGlU
7MNuyzdMANxMjXnBgQx9aaKZMks1Y/OoE+okuw7D0yoy28Vvm9QBltbYo/uAgQNT
B4XBArTkN8Fu4pFkti2WEg+gHrFRmtZvIn4uJc7G7xa+KmG1YvgVFUpGfKF7ZXMB
0lFun/HZlSjqpk4PFmhYqvq4xHIY3EnnHA4Kcct85VhbJ1437zgOQ4aqRhOn5g0/
YdYQO4q+r9zU4qv5FPvrLrnYIWM5Ghigen/wD/NVVR4KAt7TgePRmQcFB5pMUuav
VYsWJIlKPpasSQvRZtkHmTemmwZaQW4F9lh0052bGcPRiDBm8RJ8iEMqw6LjCxoD
kHSOPxuQLpu7CwgDz3UZiHQIJFdLvCDt/W+4e3DSOfLLxVs1UXGv6sIMVBc6y6xY
e71AhZ+mELF4LsCatcOWLBOcC9OxnZcrOoT5q4LfUoRckCzil25ndVHwjUuJdJCZ
Tsg6c/38229CuyiqRjRisyNYyflftRIQuGnPcDPO6AuJD3bWjqai5Jpc/H4enDXn
BuR6W6R7UwwIUcUGTrXso1DHnc5zJjlrt3nWjnZX3qXLiChDo/xvT/POpXCXHhO/
HRBeuZFGNLG+8toSMV18YSnsX7FgFr1VRaJw6LyB3/fq4uxWULfqefIH93rSiznq
wuOq8Mo1eKihVrAhe7xy/tFb3wHdsFERJQ6fPS4OCTcnbL/O8zZhLP+TfL+6AJpH
2IE9y9XyuiK3WhAlgyU5maYTUS5qh5NQwjZ5tMJqA5GKGwrvYbX8ZxDdGw52tmlf
VflnlwAdEtuF41+qg2o2JQodkz8yatCZS91cEClLMG9FDrHKKnYAGrfJvSsYBeec
2GmzLfbAFgNck5hoI6nIm1p0GJoGUwyoHIuAIhnsp0lFUJd91FrNR7DZvW+ail20
Ermxi8ehVf8ATVBQ065+lCcXwDK5nfnbLTtwHluS5ojn3oiXWUWBOGsytyT0SU0t
S4rocAoktCl/ULWbmtcPIp9bswTXQcgiQ88S2g1BZFLchnFFYK078YQ3D0kgxceC
ZBYB8SSfZKsMrU/dNQBLOeYxO+1sy5jOGWaDe75TTGXtRNshYomc6PPa/sZy4i7S
SdJ++jkY7JOLS/zvYoQOzIToxd2I1Lh7DPsqhstgmCPQgr9aoU14fLFxV2YPL9B/
nqlW3aAfZqctuTD6IHwp6pJU+Zq9V9giEgxEVGsLuD6RKOi4VcSp14EiwyW6LR6z
cjUKHbJ+jAf/rLqVs7ARs89Yj5gzICAjYex8rqPrWFxKswSPHs9mpQKkHUSVc2HW
aPGfP8wCcEtnMVD67vkVxbbZEnod7qLuWKY658cOgTQSev4TyqAZfLT8YgiptAeY
r20YD72lnvrCYXY/CxWg9h0BmJVsVLUjHwYfhgV/bqehM5z9zdWlhhh0rQS6BNrJ
NM6T88cwIssuo9s7wwbY7h3VSlQ9MI0R03kuFCXRY6J/u7cCiQISJBgyzrzl/IoL
B9X655nVMI9/H4hoU2FUd1DPlhzHM94+KEAfIu1WQ4uzW5epmu/ajdfsSIWnicKT
I0u2FKMxogvFAEuyq4s79I3CSrdN+1NbuZVv19lDv4QiOajw+lTKrt+wl+9c9Vqq
l53aBWBvEiFWqd2zOe8mG0wS88sqmBYZi3unrLqIrCr+mOnPOUcrPbEkiCNx27Fm
XcXCeqoIlmpoITzTe+YZGulddkSGy5fESB+yGFL4jq4LWhJY4HxPGMaJSdnayvL1
Iteqkic2L4GWup5Te3BlbcPhV7+2FKRObSFISFNQFR2PluBhBZx+kzmw6+X5b7v8
CRRizq4J3XDjeLMext/c64JnE32PXijy+XkRJy2otnU4HwecbvhQerqo9Kk7gzx7
BuiEODwphRJrm05Xd0eawDCIYOw9BmznHsYjsaSfZtHp+JTX3Hz+dIO4fDCqp4Is
rIsWdKZRZ7iRZThrCxMXHx8vQvAnUWEN4dkiQvj8K9xXx/P2EfYRcqPLN7veDj6N
G6YHfD+wOr7o6ZxUnKopAMAXcDExqCK6qFhA9oK1gg0wiFJi2caEvw6ovnXdWPwZ
vt/v+zaIoiHXjLQNPb3GiMA6BMX6uAt6FryUhj6VswjgfCB/vyjxMj3eCSAmn8aX
odcKfSUKvO+Ml0jekzGJBaTuu+guDEZmL4Z09myB5NeAeRj0y5L+PDeD5poatZi/
9Ym81hdExMHT9Cao3w3KHtW1IklVsSKsWNCWmPikog/12BEVQ0gvPolKYBrrbwAH
7BojMrWGPrRwDfmGl5mL1ayUUZrg9kJsDMs2v2kaPtJrHxdZvu4fTdwCiEd6UKl5
XZmSjkOgF+DMDvpvKEm8WBTZjBLP8iEaT+jSLPjaGoATumP92hqEya96obtA9sks
thpjUPjwnsYIGjJ3sOkTj9whQPaYP1IOZj6wg/3pLrYz2bQfdRTSD2nINQz6vrTb
YvD+5WklZjhqUnos5tY182pgaeLGwlvivdIVpF4RMCPS4I/2tbiQ7yB3om4bCzjK
yFDzdU1y8gKTUsuCqvCnN+pW1U/JAP/W8lLlWDcXj2jJGpvSN5OaoehQej5kqaT/
01Pg8CCBb7S+vlcMCnsyB7QmutU6toQ8bTa2UU97PGQPRGeKfMY2udrbhRXJQ1zD
k+vCZx9cy1cJY4Kjws9EMXdZu1G096npG0TKN7BHe8mU3xBYzx8BCHMQ7KqRxRbH
3rDkjmf0QweDKn2JUq7yZTjz1hlfkFykexS9KSOMqqxrqGEtMVhCgyaNhLLtmyp0
PggQttNKX7Z+fGQlL0BloByjkIAfRp/r7iVuF+gOxoGBb14zSF99AvVsqCit3AWd
azovZ836apIYe1/q5sU1KtTiBIxv122HCNjGxKWyLIHbq1V95FDzO+I19G7R1sVU
xCBXUgEjfQ2CDqmWiB9Yjdqx3We/UE+mMUf3+p0QKMskRJX/StNS51YXi4/TJiX5
TIYnIbqHDqTMklrpELxR6awDlvEhEXTElfxg+g9JFjGoTwOrCm+bvxPRhiXW0cC9
w33Y1c1sPtu5IkjyA7KE1m4VAYYwPV5nmMWwx0jk1h3I5+E7z2YVBCnhAAu0DVr1
VY9npe2t4rD+Dv4nP6oYu8nbM0X4Cvek8uvMnMP9ndQVdYSJAFWbAe5YVZrxC1FR
gNyxDZpbpW16YHb4JQb9bqxQcAoQk3lfTWXB0WbX4FvI5BBkGDnTSy8U7kcFlIpT
aNljyNLvJfbN22wG+ByHyu5Xy/DH9feC+zFldbmbj/IEu7VJUJ/vrddorYdmyfdN
GOHRHH7aT1kh0HKAgew813jgF7H8vbGgbutwgaHHIG+i2gzVRvsBpyedgmayuyc4
kG4B9lNIZ5fzX01PVR+GzEb7ObFrZM2DLcuORIMENA+QEz1sG4R4PHCnaW1jV9Yc
3/s2KhyAK6Z8DDZJJddnrFpTZbVv8igdZZBsFoquiqIbhmtEyRCVGAVsheSHTauU
zuo02UdW8l/EYiCohmxVVKzGvPKlXoMpBcz6/RK/r0QNmOur7yHbZRGAH6UD0OJc
HmoZTe45TbFYnDtP//3zmq/+K7nav0cHu74kxry1LUBoH0W+YyCm0ls/thr7Ms7o
rlQUS9QNeYHFKqkjJ8Eq+0j3+gKqvBlTsf9u4lzBBfSRnZ72Jv7AMF8U33YTZdva
ImzzrkZWVKhY0R/IVLlYzgM4+K3NFODmu+TMU8VerBlK4MbMuBno3aUt8CVTl0l7
OrErNFFrGv2MjNB83psnI4472F5vDZeMKdpWommhF27/d2wVoPuYTBsNkhmVH7yY
6t8Hxqr3a6eYfWw5owUScD0/Q/LTrHxbMohccscXL7KvAYCWtg06Br2W7BBrrimT
mGcORMbRYSLi4KoVtAKGTUclgpP5J8Skfyx3LfuQBIj3C7huD4m2CGXNtQIc5xyK
QzViUMHpCQVjdwJG1SGrHfQJhwGhP+KRV704KrFfz41Cee37RNrSb8ZaFUoEarVC
gh7+QoSlxKqMFsepBjBwcN6C8WE7B5t/EbCMd8bFlAHTcyVH2N0UAzTqRjzcw8d9
hVk97Hwtni7Zjm/O/3TKSOMMfz1bB+sfbn4sncnLiXviishwY12Kk2/iM2pYK6SD
xtuIOfbsLyUWivBHl3SJX8EXd4waZQ+fagZ6YgSW2BJX23ufmXnZReutJb0CQtLp
yVObt5xRFTBPO+STw8gC9SulW8Fmbq1zjrIY+AKrJYE/WYuKoqYIOquITC+yI9BD
zZdzBD0rvAmjv2QDySgb/yNhPBf11fbKAwX5JNgWd8vG7XpP84Sg2z2nNzNk5gIZ
+ZOlKDHFvlr4ZvmgQn+v+ViWiwQesFoB1lv8VGBeGnT52XPD3gngjwupJqx2wb91
pwwC6KCPk4pxQFbrUxvsT1HUm8rUv1lflRvoK6BeXWowp0qHRSdM4iZYIE34Znzs
AW8t6nxJ+mSG2T9R9WPJCVCwSqij8zrxP3O/stWLLHJjoDSCtxIannuwQXd5S9Di
c3DoNGIbJlNRTKpyxSJRoU7Vl7h73NyWnt9ZT/80o5jB38FhuXdY+2WoGUMzH4Ty
clZyY59TfRe/ePdymDIwgAfrBG47fxwI4TmUtW9DNZXMSOC1rHIDoiodQ8kLY6DQ
PEXyXD8Ph3N3/EzrITPiG5Udie9ww9EUrR7oUmJ5G+xGvUd/HSUo1w8Tvt0HZL96
/w6osR1G0xglDZ+i27/jyNG7KYjVaquUn61DIxXrpS1QoJaWbaIDUWa0PjTUxLRE
lVMaIMZcLFiuQ3x9qSLE2WMyyLIIEAKGgq9wlVul3bPsWwkTE1AU+bnY2brINWyl
i4gZbTOqpPpb+4PiMhMC2JK3sbE+7PF6mdiG4WQs4o8gC4Ta5l/OHkrvmYqnFsGY
Twr2SvSM7iUJWTOinwtqzjGZbnaCFDoodSYz9VL1K1M/bY3JPO4eh/HQwUUbDWhu
Nc9T/BhbI/bpFI5dTLzcTmGtGm76bvq7CUKTQkXykRJod8ahAMWkrD5uvwXD/8Go
PGCKPThxy3b4vjVGPLy8cU3BJ7Dezmah7zu6zN8XkcVR89d8S6z6EMwuG+AMW2Qb
c7OARQ7g3SXAMxEhBLTWBcKFjFZtXvFuqSJhqRuWDBFEg/wM74aA3KsIT1l+/O+A
w8FHhas1EgvemTDrJCZbiX28P2NeB1LTV/lA+WfLfjuNtwoCsXwoCu7PPrY9tisj
ZZESYvY7hRpMf/bga3oThow2Q1KKAHYsJrAvYXYFRF7xGjsCQHiqfGRBhz5dTu11
YTYqjdGCbEBgMrDf0QqqtPaBbNQyPG54eHDCdwL1auArpm4SYjTKxDd6CvVicCQk
uJY7WEPc2kzPL/X1qWlJ8Pb3dQ1rP1G6v6mNjvTfDQ8qJ1SkUcD8f5PIq1yasYRY
aEaHGHKd75s07LqEjbOi/8uLn+vLo6Jm4HqP3ZezwNT4jADA6O2d8d2R4DpPjzcW
tsD0VJq44xHkY3TZ8OEO02vkv3jK7CIC8TikPWyV3Y+iKQDFZbHIzU+LrEO+Qha9
eJCUSlGyVhhKtPN9yUlEhBBcFPQnyKvWYMv8aQELPrEp7xc7htTu4c3YVj9qmChd
c2uU3KQJDubb2C2SfWGqghOtS3yxPkIc/0Teel11P/KyXI5eSyIfmzx4mWyKMMyi
QPaJxiy8vtPhTWjhEcBZAYxdNaZtqTDlq5aU6i9TDzaP2qtTJvm/G16sRk+fPv7Y
czRgGV7LkS3OwYhGM0CyNol6qvfPNBX7/colzx78eIAcq9dG7woWHaxGumDLWEJY
OanE3YwFvakY3SObMrNPrEqOlb5SLU7bThDMfxteQh55pVKcsBcgC7eKrFC9ipd1
eHSm49pVgOWACXS16PbCRJAmAoEg4e5gu0RgJjCDFafV7k45rI+D8WH4GmRw5Ia4
foYZRJSTCBNilhbjuBtflU2lh/pbEQY8TEng6RXu4s9y68hTWabGdzSZAXaAcva8
j2lg+Sws+30CdpAiOOYfnIcDEdYKKDuOK7IVqog8CLEJ0NcUQvTFxranA+AnXeZC
NLs/N/GU56839r+WK+IZbX1m//0VPGEJceRIomdb9FBG56yAmq+Z8S++Nven8xCI
GLGNYUQNpRMidKWfTRhos5a/ejOQiG0pghVgf1i22TZ/TahDjlkVIGfg9nOrsIWE
AuMJWKh7voEpEB2jBRfXjAylk3ahe0smlzEw3Vc/zm+rfoFLotsrLnHA0sD73G5G
c/vSOq9/w8DAhNJW/FOBEwkhZks4AxOg/bW1VGL/FzRtQe5mtIX3ymBeZIZdLJi5
cNiVLyIDXOD5dcswB4eSDCf3WzjUrKmnQVzcqCJqUPDCHxeH+3Ma7Cj0ROmojltp
0Ui6PQom41g2vyBHbPpM4y2Ei6NHGd9A9C36peyiFJ81Sj9b8xgWPZayUQYYSF4n
toKVgPLyWfjQtQadqR/sHeq9OJp5nCGNM/x5TCcjTtebF+WsP0LqhyiT3LC3WT6y
G6RxejaYhyRQ0HymdgPMfZw5gjTD902X/9I00DynFYNyLmOEu9fL/Q+Ygf05vWkk
XI6F0S57Z917PlAtyTYA66hS5TGumSYFHmtYywD7sRi+BXJ343tmseVwsT3eN5FF
rkRk9+sz/DUUCcNtF+XWObmkl61cPaQF7zCqdAxaP7ZF5tKkTM+27a+MmWcot1Ka
P+j7Le9Hlraz4G2o7C8tCxiGM2GJEVyvPlGQwbk7MLxaCcZc6lSDqGczHSZYUHgf
094tQKp3tBehsPm2ZVEVUBcXF8UrLVe7PFFVAZXpx6cSKXNbvdmUC1s1p0LwGVCj
Qtvu/Ot7ctxq7yjF8x53jZnehtXfCK/bjiEcOXkKgr6xrRSBruiNiGBnhsJBveD5
LREJbiVl7wEcx+8ICMGM0GQHExO1B26NDNWrnoEQbezbgy8bK+KZseRWYgSNvjSV
e/U0Wf7mDxuUvghE/D/lNcpX1g9Qp7jM1Wa1xBHxzLqQCoDCKCoxJDc5QMUR8ys1
vvVSTh2rpyczXk8vguWCjmFGcA0bsFTbLf4N2740VPrVoRZs6PfwXqG1UmrhifZI
AKuR0bfwP/xYeCBDr733yjmv1q/IpRmmZLGhwerrMUee3RJ12mqx4R9JJSCrPcGx
4hEaQS3R4jmexW9RbvmGh1Ed6qnOZYNbDHGSn/wdNZ3QiVWtlBJjlOqd/awR4ylC
hCJWUzCMHGn+YFl52WRdNTmX9q2HCyFVXZYAnmGcWG/hnAnLqgTSfhwPzri6iheg
hqSy+7scYmRRVOSf97noZFAjS6QxSJK4QiDEfgQO7VvDid8Sod0TUizyGM0uME7c
nW8NAoKFu5hiycXQ5TBzgtrmymHUr5Smt+VPdSAdWxc8ZNxu687HQzMYaXQkb327
RkfrFcQr0CF9XZm9vsksyaL+gzBX7P2Nswd+kX8kzzki4M5sL8P/bakzuOufJSyB
SYqQZNW0N/FEeECgKmBg4fVn/19/MYBtKBLWPC1jNcgLbVBrpP486bpdDZY9kH2x
yQO9rBKFFnFOSe8cpbAsLTiMd7fafCdwFePMzo8N5dBTFlycnege6T79nfVBCDui
Z9VRQk9tp7JDopk5LE5HUstlmd6nZ2lS1rSAEuZHnsShu/blJQSnT8NivjGxNt9j
Qs1NY/17/LJX9Md8NbmP+doiOy+ajLGmlaQHORzGxOEaxgMQDi0fHnzOtwLmtZlg
e8R8xpyRqsqcRat2XbOLmWVeoXYTRpM77qkBUeYbXtRFYnwImix/rWNsInhihNUW
a8pAWUtH6dK+0fAso5mK2tn2l/XWpSX4ZSM7ZXRlQOo9BAoqtCW73+behF4ZaiZD
/u2tLYPamB/SGPYk8hh5PNX/DOnTDLM9NIl7YP4xbanMRddrGnCfn7iBA+1kBeIo
Am4O19bij7oUiEbninSgLxQMSgzEkmPcdgtfv/p0QgAZC8MtbLHSXUgDfFdsv1bO
tF9BxjmcHkSbAl6FbYrGGiHGurTs9Um3bM8tdSi+4Fy0h+cu4XQ5aNL+3KhwwOcI
4h2Rf5RgM/XDLA3Q1cwkZqT5+xh2199OOZF/zzv0BzsUhM7vNdQinAltAiTcQxLM
m4xyB9dGswydnUwvMzX0w6+2Ads6Xrq2b+8I9wnUnLEroDE53CFRqqc5cDqz99iR
vs9e6FC4lyjps4Y1hTwVgVghJldBhnoHBNbbYBj9Z2gqrEGJXEjS757ZIxi2JQRV
BC6BNLZpMkNpKUZCJgdT1VXy81S9MMGl+Jk3iZOyPvGgr7+YPzJBgN5oIFB42Ndr
AVePxbEfcNNvp/1HDDx2mAEYKcFJ+sufhh7oIos5P3vusW274uxOPLs4syO9IT+M
vUGG2PXWDozBUXSxqZ48UclKBmdMelMfTR7Q0YZnr++DTS7FvbkJ5lWz9jYtDv+c
rbqlNnBDNzn+OupqX3SimfpQA7CU0IcnWzCJD/aJSH7B6sEw1gy09O4kGqelftgE
DJqr4JtONjBJy8ZwFSQQVyN8akH+N+otwPwB7/Qx1JbVRdU3PRu6bgAXitn4tSsH
gAUtTB2e8E+m180HnU9lilufqBCys6dRL/eZAzqtBAFf4AjLlfNrtOXsxbErsnzu
SBBm4OPHeGUM4pUszUI3cX02KpM0kFBJKdtZl+5ImZtVrqOjs2NzOODCFoY43pg6
M62RUvUDmGrdfM2ezf4BeQkKmUilZyWUPr6Hyp1TgymvgfOVv6mU1Xnt4lNya19z
nxdP8XsiH6T/TuLzqe2QYqoDdulZp9jUXH9e8Pl+LSeShA/7j9Fl9NsHMYCnxaFA
GXYBzKVyouGJPtZ1OQR/L9BVQJWjfqFmX5RR697AbrAEe99Nj8zHPno2yu3M/IBH
WXKosh2dU0acFOe2efaXIFMfdQJ73b4EZyQJ39+hSSIpqegljnT5oaXhpI9Wl9m2
Kd/rY4B+OXulwqW8a1w+B+b1SHtoh1qsItIpBw2svH1Zp7cImCdrfVM6smRmMUAW
CsEYoeisH3NRdJDmtr1d1/oiOjvsBLyFBsdYEQRWPLERPXdUckopSKU8w2uQxq2o
eNL2T0zUPXdswtVwS93TophtE+kzV3Tk0JTEeeJHzXVxSgnzetNNaenxKrvuw4Ik
0o+9x/34hS5VZQuWZRWSwLQwCWfkL05y8TMCEFbn24u3bdBszdPHtkGCgJPK7vjl
aaa4+SntK5oIXBOiDY6VkJGJpm7JHHaU6riZkFpwme0T2g5jfmhNDH1bwBi6+zt+
5v+Qj3wCgSo641yCCwgPvFbgTEEM2zNAjsAEB1Vdjy3+I21encb8v3m0x19P4tPP
05d6hg6fuiJ5a54TX3A1si6hpmwsCouVNrHIQqf4dUK/C6XzJGDBioExOT4BX725
I9gujwWWJowV4SV7XlrfwfjNniUmBhcN3ICj13Nsh8LUS9KH0WPXHv41Ymbz6Zrf
1a6OUm8BBRdeY9qN/pcHvRur26V7P6WMM+0yVZZhDZnoj4pJYe5QCPAn4p8yJN36
73j7DA1QB7uLlrHaG741GaGuadLqAvcEbDgPppFNc6kizM5akDPc4W9yq/KxhD0P
dpWSmaYn0xd5qs/HkFLJIyRCzMHIzhqAzovwlPOzcd9xptHsrwpf5/yJ6W/94R4I
XpqXdZXVtltSwV5aEQUP727wQOZXI+aohAS1LxOKzXojHX6Z7u1/2+FYjWjZGzTG
oYlRqNkjRTqlyEd1czYSzEW4NYacTsOoxeudRpO2++bGbKXFfXx9m+xuX3/xHHD4
NE7mFCOCeYuK2rFJG7Vg+m8TXtSpYxkuwpcaQBr8TMezkhNbS3KhntNnuG4g1LbX
TBxJlrzIwgk9u/yQ72J0aNlF3YROnmbI4qrdx41zMbyvq5cxtKKKXKPeFaUpnUom
1bGtjLjzyuWgYonxUscmMMt9sQgINuyICKgZmXA7EoH0kQzvitg2C1fl6YXwN+Og
foBn4eb9nSNWnsWTLlcXfYMdQBeMWT/Dy3eit6VOOzFt2Vagv9bIjSYmymEBN15h
1llSnYMNXJIA2aMa8uAnijygzYPjvP4djM1IlnSZcOpHOFtBwQiPLpr3trzQvZZ1
v+SDYZfXOqqhzHLtXFJ2BtDKhImA/sdO/pQpJ2nTL7U970OtCgN8a9laNCgzfCLe
aTjmQS3hSl6WOeHsLbti4Apn9Y5d82MsDj189B4X12A3/Rhna0OpfNuZptB8V0l+
Vtcfxzv7IcchLRgT5x6t8shZDJLYmfmmzVvAyLKfhiZ5ZFx4vlARIG4bDyl/sE45
cXVtQtkGSfG+Ly6SgS2WMUDKj2dIXbjoQtdP7Ifryx7qvgFAIFQu2frwu4SXZcHT
Ols9V+0FmUvVWwXvafvUqqNIascqL8Cvyk3Laqpu6J64kJV27HAjVUrKjFl173Kg
YsRI/jXuFIpQXhfgrSQlMRRsQi5w0ccXjn8EvRgXVkeOOY1EiCwCQmHqH6OvOBl5
KK8k7zF/U7T+JhrlvZNG4jjBJinq3vSWHhE3u0LLgb08PTHKU9c8AN0GtVE4j5kp
CNgp+w1aSA84JXR/1ha/58IkXPdiYLm+tSL+N3w2cKgdhygjLt/fqSpHW5k/tiqh
KOdQTrylb6S+G/eROhynWHLHnC1ERsuAnV3uvIGIkPs224Q3d6DhcnLMyEQ1AeS5
iKLam5sZJkY2ahg/AQT6yDAMuThjx0TcGaR02BI3ZdAwbMUALAn9R0DzWEh0RPpJ
kPOTNB5UipLMGrIuEAA6wLAegpuB5e1qMBENp54C+5hsmdp/41cVidXo1kvVqtlm
yGulSbhxx3n+7OtvbJRyEylRTp/cUeN93oyd9qxZdRmpJIAJkzMDwRplhuqZK65H
yfATsZDoY0NTDlCrXTZb3fzTdEr7MTLbBc5PNE3t982L5P5qFtzZwFKOP5AF+vG6
4ptNZ8W4UdXvaNocv54RpuQ6ICZXae+hbM/fXLvzXmNqVynJn30O2RUdTTCYDSsO
N8m5bw6nA3iiNUVJlQHVg0LAmyS9tlh3BSbJk+tP4cxPEcVclfcrHTKBfQ2S9kQ0
2/BZqpD5gdiR8Ni4POzapt92Lhw1zkSdlujxJXnSxx2G414YgpY5+hzGkrggRvsu
QYBpwr3LBhAPDaXWvbwTnv642uplOMYER/sG9RMqQPgBF+HjsUIS0BpVD9aXfBl4
Xw7fUOLFOjQZmG9PCsC9q62GIiG4RoKBptn5yEmmTKVGp2/1BOSZT+xAMrkI+lf6
Q2IDcPhAkmaJ/FbG18sN6AkdnVG1R2njeMjX9RqNXpsrcc8yYIW/3COvEn1sadXv
z4lhkKklSUZTOMX7cJwqXD7h7uogMOMrH6lVn9vPAba8T/6SRYptiBH3TChdXGB2
gGN/Mb17SN5BDylrp+/0A8wXMjO1q1iR6wNUBtNlGagbo7sXZu8RFHBvsoHiLpoW
fFRQlDbXZgAgQMB+W+AyMe2bNvJaiUZELodPvB+BX/m642rQLuRjnlS8LW3KXf89
t2zq+9n5BCmiUwdRvB5kblR97hIq+pcrCAcmHraJ4PWIRV0wnKy2U+d4ak3AbDBk
2i9qoHBDf//IuUOg0nnKGc/mBH+fLvNSey+GpPQcuP2ppxHdi6b2P/YV3/2XtBxv
cuDyGk6dRwFJFKfB05k5nNOVunbbYRbuKwwNS9n5aivpwFU3WwIAMqbT2higbP0M
3yyjTXbIYDNWn5A17HfQuPIlquTBas421ku9yhGpqNS1SeodCxMndqc0Bmgo9Gyr
hOdvggwg5FmNnSyUV99T2LtBlQCINHJgsHMB9HftqFgLGgoXmD/ftqdQlphNpT2T
0kz1U92DhV4LWeSTqm1A+NaXsnj08U7Fqc4Lf2YYcKYWT7+ynFDgOpTW0ThougAw
CAQ1BqfvTGxUXx2/CBwR0eacWXxJe1eEDAPFLbFXcWeiBzO3f944ONbnZAfeFXLr
qDHxK+yjMJ2anGKgcdHo6wgEJVy12D4SZ/SMpjh4dZBgfKCPDGvVUYzwV9M7yOoE
mPWB6Zo/OpJU/UrJfza7sRuHjDCmugrRWw6OeuidKfd1//cwQUT3r5FeyWQOGfRA
ZzmnMLzwJQDNEmCkAHVmzGQQMtQJ7OovexZUvQQVl1AlEYHYmDJ8nKKJIfUmtwqf
Un9kcKzii4M+NGVNvxbpdEkfu5P0z0tuWy1jU+oj8xL3XmToa5zCufn3oKK/KFZL
+qisE6oj/8AmJni7lNaIwlgLI70BYP/GdL2SzWgJV6AMRH5m65BVeGTAdsQ0XAHX
iJSnmHoFiC0CRMGbgcGRfB0Fx/6HtHrYPuiD8ehEWLsJjS5j7DHgnvhAKG9d5+id
u8tCpA4AkG1kcQy5RlsP7W6QvDCP6I88T76v+dDk+bR6E6CuFdhgGI3CeSzbrbDi
2lt/u/aaL7qfSBaEJ5i1tOumgVF4dXtV5x/Mldtd4ExVylVBG/zYDW868gOeEIBv
nn1zCBQtDmWF+yW8cK5dvYugrDLtkkLO0DpFtMdR4sOvoSYbpMuRJei7CVsWbTLt
aYXF3GB1j6W4Rvh3/nF3Jhpb9D1rvHNrev8nA5aGzm12pzAekf7N0NpREypk2WP4
drFLFyuZnb7tkH/xXb+7FtLMaCQ8skCxBztwQsGpoK+gcIqf43O3O9wMerrw/kP7
UBMTO7YkAkY10HDfAL2l/8svX/2w1qI3rBF6tmXYp0EDNoyba//ZRMmYFqMNGBrD
omy3KeZijrP9UAdsM+wpF3jS2cM447fhEHqHKC6Dzk/qkuV00yEpPxw7dhLB7GUQ
86R55K06OjDvNO0bBFcnZN+xP72n0d1gfz58TaoqVV6l2IlwlsxF0pUyQgwn4khK
/23CR1uLUInYEPhpUrZI/eaXSFaaH+78GL4GneLAozr5DCO3v8eZo84FX1LLQnRf
uR3gKlEIuIlvft+EM52ACVku/U6voTAOx6WFpZGzONMnJOIHXvCp6rCKeGXWe9eH
2xINqxp9Cr8W/H6aT8W437X0ajDv4fD+UwlBIqt7ShnhPF3wwDpY7M34y+w4GCsw
pCycEqSU5AoFIQcoSwPH+8AexsHmLHpUljUyelqiIsFPhfOs/y2W/3jRLbCNdcrr
nW4iqBqZDQgkhR370Irw/xt8uTwo2RkUcGyZPJzlyVYQ1vsuB2kjQyshX7FW8Rhe
2AV6X/GwkbQUBVNXbrik3h5Nhqka7MfObuohQD/Kq5Iwwsn1mljN1mxtvcbck4hM
HLeIyyNh+xSjnqCK1WTRXxZtMEuYNtjTYH2NtD4C7oeKzF8b0UJwJ47/GURl1of5
NdsfzQKf8VvNrGJEi7unlrmEOHl3hhqL9Cuh5Iy19bjEcSB58k2a3WRxDY0fnk6b
v2OV/skb2o0ZBepXdWmsVJDJ4Up7ZPi19dNHvV1GcsHG91O3JSZ/VSSUqgsSCZE3
Wj9j+2CTyMISDGjkvz3ALfNdsRqswImo74eza8ozaOrfmCMPwBOF+faRfKiFgghf
Z+9TYtnuKwPZcRK7Idm0MkIl5CUVCDMBMwfpM44DKj887fCuPW5/M6zHnno01ls3
jBuBD8zVHFQiiBW6rXu4xLBfXssj2N7xD8snL4mDAP++2fLsPgUEu0wzpzoxVr/5
Uepr3FyFXGXF9BqFtfcz7kLDvEpkGqf9XbKcy9C+UZ9BAvB2ubnjt84tJKftDrz/
KiJhC9Z/5r0EwWkUQOHYVEh0Nr58CUxsCesW8c93mFY1W2HBi3RSXyPxen6/CrSX
TGyG9e99463Q82vZVVvhPFRe9RHQlXJGNBcoOECdLopR0/vhUxQQr9iLmZffiFeR
1oIOdbbIVApujddU0YlVii7Gog6SAmWDIEA25/pmK9XjMd7vRjwPohYcNr2rVrPI
xlJSxDin7Bxv/AXBnRb1dwfLc7V5YoxP5XFsWhR3DnQlPnhl44qRM0c0L0BxubqA
d5vrD7SyZOhsWSEjbKBPeKXZJVXHUUcyiVDZ1KYqqk1ZiBovD9HeslkbKbsiAV76
bGkPxRIFMRQk0xTLG6zdUtKUCpeF9R34fuCUWoe+VCFE+nEk9xsrRMJtH39thkQZ
qTSvx10AWaa83eMh7+jP9KnOGDms65/WH0QFURb6wJvedy2LtEOCGVpwhCfiRioW
nTX29t26AHkXpz7LYUGmz4T0ct/3hhbCa/uw07OR8qcL3aZkPAtovrT0mh5UIpu4
22N9cVW7O5rQ0c1/rJ2IVm/vkud72yt9LnyrwuzRu2D94q9tfGgv4epEvqBvKAS3
toQyl6r4W4crHrmYdICDGSoYbvKx2FpWE2EfkMUKyorytGRVo3H1aXBSKBhVhp6W
id8Sc7DGtXg83EbxdCUq8MPCRH7rVqLhuc1+qtYj5C5lh/1Hqj15CM6trQjqkl8x
jUusjGB4NXE3X+mL5wWce06BYZBs7IkabxHvGSZLpOu54uH3sGojDEJMxcMd3ZRK
l06ZBwP8JJJiOb7afbnd2cBwwB+cE07ivvIHIn8oRTKuJWs4IHC+9wVNV3HM3+Do
6EQpTYNSuXR2UarB47gebGENlaSvP3DfUog/2YyRV4YVjtFeAwPeroeLgJy/jtzI
IZ7ENEhMBN3rKv/gUpehxB62C3EXUfS7V19b+yyFpcpqWLKSdkRkLdta0s3DCgsw
kFiNDC6t4UwtlsLwUvcf30ZbhfQo6GW8RcSTUp4fz3rVXZa17lC/xnft5drMGcEy
MV6NUvOJKgRVXX8XD2CLUqxzMVE603M+ag4H4+4TPrPYzFPiZKyVICsvjNc/CFTy
fct/f/5mg2A4iIu+rv5fVNBSsaOzqQ+IOYG9e2xG/iLJ5Ni8YwnbqW33LIkiiqv8
BNHt/EIPM33vqCsJ5BaFFNviOJR1vJwoKzpWqBDlhRi4Aw5iM+9gKTUCILzcK8Sf
+oa+ovQvoysY2qLNyYbbv8LodXg0m8P1sf41gvrs80yY3rRWXVuDn6LQ03bDW+Cc
b0oHdlhvSuzQuVnrXsRpZF107X1AwXQbJv+XTcJAVitU6mWJFzAmH6kstNIJndqi
7Y1VHLbSOwixWLjJng9lUvPGCdGtHeqFh8hluvGNDewCMB/jDFHMsMTQQ7eRlaE4
zLrj3jVFg2lJhRmCn0ncuvLy/vAVddYPY8y9CYTuCsdMXfjVY7AphgZM4yv3qj2x
Y5OtQwo4cJEr48Ws4xspg+cKnVbBash1MzswlaOm8QHfJxt6mJFUZ78DoJ1fWh/L
hOx0iA1i6SzW4BDE/98LFkGr+xUCe5/jXeWOrgp+V2rpN8uVbDf+ByJvUyAyhqgw
tAlPrX1id+roVWFYVAIWvUqr/B2JARHT4081nrxL5lCzUAbZPshVCVxoCUcMhl/A
ple9CK7IIV3r0gxGSvr7BT47mqCAH+uaSOOeO/D1vtNwlaZ+ZMDTI7eHHwHzlqKM
k1pgvuNNRj45awFZrRzbJx5pAhjBFCKRDbOX42/RgYVe7ebj8ePM7wWJPlx1XQSU
lFBzZbgN/vARZK/zoI6VCCQD42bWS9XfzSMAfGof8Ivn/fRGUd1mCEJSAiRikweD
N6bUlOAmUMEoDD6XthhKIhvh8SE6Ixv1Ov1LvdQ7WVzBCgitI1JJwgK9lVXVJd35
s2o0aVwjnKkqaoDqJ88je4rIfKmS3ecnvFqyNnN243CfyrkYyYgtLUwmoLeHCT9H
0TO+lQC5hNr17NciYBLCoa0+OhOzZ5jp/8dW+G2T3WtypubA5uV3DYqkCxkxX2sE
6K11VMD8DqzYw+Zld6HZfH01uuZ1KRqIk5CdKL5d828IBqR8XhjnO/KJgjzn66g1
zklPOAfZ0ieO0LoyhaCcPkk/Hov3OkhrgKJcFdobyEsDn6KsTxScMARaJPxBIE4+
fQLvpNGGWc0UOyaoMnP70t3MO7yHcyJuzOMZty6Q9jZhsSTnNv7vKxdKVl8h+ENL
YChZ6+eedT3DocTxenAidL/SwFRZbKjSwRIfTji85mfwFvi1DY7q4QuhBY0+iIcO
mTms7RdHyflY7a/t6/BXKZYkCvHjHD0QhmTnsKMGMsp524C9YL4r37gP1FQ3PhK5
WD8x4Gwj9Wnw3dl3i8on/Nrdq9XxY9fEEJh0TVmCqF2Kiap4VBOh8iRlFwvQ14R7
v6QxYh8hx3OksYY6cdekFfotAkYXc3wgM6Aj3v2Y1Bdfr6ARQDeBp4Ma8s1HPYSG
dHqrtVEFgZ9q+ijPc+Ss1pjyxI7B42Cvjhpim1K15ZItZhk8upnGb0ioABKg1B1p
Uxk+evL+LYAjE3it32UASEKDOcNJwoKbNyAF1xMTreTdOZacD9n5s6UJOpmf9erP
WS2MdQmKfIMdfV6Tpe65e3qhVguuUwZIlqjVoZxacp+1NiuhDXk8neNsM/oSYFx8
WnmOTADk2t7X9V8vA7btnzl7MPTQPd5SHHUVb3tfdGjDK93XglLIG8WYPnWD7luX
VL1g9746j2fP1De9iOnpkhgOZD/IIqi7mBcxyfXkPZfYJkP8GgE0+vmjX6KG51sW
TgKyuOpRstrV8R0zNK1oqEmHCUrBa/Yay8x6NLBEPp794gFmUTvQbraElpPmd8vT
GZmNfF5s1jYUnobvYxpikO19yjjz5xjEjs+kc0rmvfYfyxEvOXI42rYwMTb1MJua
XooCwrHkrdy82NC89Ysn0Qvh0BJFdl4dUktd5J3qn9at8pe5RYufzV0w2JNnblTj
y98QRJzJR/DlPRScSDT/ssOMSybLvYPaL6JwsUOqR1ME0gFF0LD5zGe6wdABDZ/u
aXz1N3YtfciGZ/YpvkMVbgWgFS4F5tEKCT7hkSE0gs1bNQvb2O+UmZZ5v74gkHMs
f47eGrkpxB9BHk2prd8Ahj79e7n2lRpxRr2yvLcDPzjo+Ij/A+3u6uSu5qVu5wH3
4JRv3Qoom2xyi5FNaeV1mo+oyrr+BjVAPz78Sg6hbRkMfNhKFrhC9vj1VHb7Ttos
lINCcxKGAMPTDv9zwxOU4y5su7G/51Ts4MBUfvr8qqZ606dZ0uW53Xce7bwR1vql
i46Exn6uUcijhbu8ieRbdWDZAwBT4ZxK7r+ATjgTQ43WfFmDVPB70DKZ1H5wy1dD
urAelhc0PeVrV+j44BvePEuDsMa3EierJJRjXRbrDgSZQsiy+aVUdhcMTsPGMKPf
uk6iBqEEPShx6YmTyQw4uTWVw8pPaVC5uyMKJDOLCk3gW50UWKgDGy9N9+9J8+68
TIqvAhrjx6bsWzZutGZ/h0LxdttFKOLtlGKV57NoLbPWrS8U9KyaP+nHp7/I0PZf
nVnBBnhHQSQOlUjf8W8EwwmrlIOvyeGsQVKxvetUVUrNonRjI5kJuLDpr79uH7by
6VMmY2cyYr6T/r/eECQlokcYJQIamvcLJ+7PhS/x/kwcD3GDax1w28P4UQqi7UM/
zkytaSFO2Gs90GO+bLdkEkm+5+FqbYPLzEkrNjEYwkCVZmqLnCwXJUOjm8dG0m6s
yD+G+aGqBk7tBhP+zkv9SdmvQmFF3DwkeZcBf4MCLalZmMahwg7AfCz7/CIi21AF
zNX8vfnmFRYk/dwZ8WSTHfGs7iXi1EdRu3LcDLr6CPMP6d/XYRAMeBiTWTyyFd2n
6pQK/2TxzUQz1gsy6+a/N0L7javv9RKVY9F4EGXohaXOfj8p7E1DvpZSxcpYGVwL
DnDFfJiCM8aiHobe/iBgody1y/l1+9WAA711wclp/qyibjf+kRXCdfheyLc56B4U
UrTcLyisbTHwUisazyzIp2LW2wjprxLJtQXNZ3G+rivfvLmaU8cCkJ55aGGrA8EC
aoca9ujok4zAmtQHeqqVYWykOiaZ29/okelg7rSZ4JT46mrT22uo8vfZyklVw9qd
3n0d+KlSe5y/ydexCxBu6OzwcE/PPytkF/8GL2BcpRqLhe+9BLr58NpERzR/7eOE
88shZurNspd4W3AS0HqVIxdRFLc8tmo5y1szCAMB2oUJPdIm0qaR3saNZL3KhpKP
mjzZpjT4pRoV0RsFPCGcC34HSKKBUDRDC9pCHyCxI6lJA1vh20vbsKbqviWvE4RK
jRIdk3E4nYrv3JLx/eR5kQ2izyvl0JYRf7sXj/u3famJKwPb+d3H/E6SfjZ38JNl
I9aV/W0ef54jUz5ohj5VbeG/dnKyd1oEKTOCqOPiytNMP17u2TMgjw1MIdbND0eQ
d3xWTIro98FzenswW+RvK/9zooovsL0zRQxf6EyOWxkqGqBB0JXDyezjyJENdeGr
Y2QLM5pvPCIIEXagJXY2sWkbSG3NaAwaZgz4XJOUXEvMdS2vySyhakmamZ22p8NL
uc1IWN8iwWYWR1QA9F0PQwHlMqHwgvvRpRHsxM8m1YrwkgaQSfwIFokrVQtee71e
uYBOQNIgpwCWrrjv7nbbQ0iaK5vxW0tOEynX9ZEJVOPooxAqtXCr9bsGTwpRbjZi
5gjqHuZsfmS3K0dToY8Y8wa8IWyXRZsrZ/N3kckVYcTGHs2Ah6lxMSNuafDZB0zN
LZaaJpTUfR7UuPQADNHGLIRCadYWaWY/iZUsEFB7Wwnhy7Ey5FfB7mw5DLUHv9W+
9DmbaEBrbueum0Zg/VAHIZgW7QakF2zFn/f4k5GiDNK+Ah0DUV+WH8UdsOpE77xo
rWbqq/3zH8drA2cHeUbeBpSXJMd+Gre2kVcOnwdLDvBRXdES4hH/MVtbXwlwLkCB
43MZAk/4+QsRVbULTdfnqsyall9t1Ad6W0wdTSFm/6laqg8YXUmLIspppY0HY+9Q
aZbZmbxOsguitxwSXgJ1yKpGUwr62wxcj48K/u9aT0ooLo2jPcxDLr5khfHueUal
8FkfT8SzB63jiqwYlzXEBBWMBStwNKde5kwZysiIt+ulZym9X+PRuSFEat0FYuOh
q4eDSAirW6TAvljikOAzrgkTvhl/92DP6NvArh7nzVypylyPwlu5VTaBQLziKbFm
W8dzeyY+HbP21NCtv1xduXklIFGKCWhVBt/KYMXir/JtIC5m98R59qWQjhidpxdh
zpIukkLCPWspRU8BpPUcD8/sTf1xnva1slCSdbTzhVWswK3Llpu32T6s1pAmzvir
gieIU4JmLJsMN/Uk+XQAZ2dfo1AtSZ8tZ+E+M/v4HG4kSGGDq0WYrh48Si/2Tm0X
IwbX97pIG3agcQyeXBoYNqbEQhqCD94TEACil41uVoO1LOYI+FgFmu7z1AbqFUdn
V4upzTERfhOYvjhkB8Qwq/uwek7pmX6KfGbHuN6m4CB+/CkSZZUg3CK0FY5ryI4R
3rE+AyYYY2QPB8ly4JoF5CoRB9SHaq8ujyNqe7VfOSWVjU8+SonNKcFJl60rdktH
uQ7EeTV7YRW3kQOhv5yWRy0ONSwp2c7NA89ewygtSJIDNf71ob5N2uAokGfqx8fa
Vxa76RdUDvf0yli5wER1tShtGOJzb6hJiQ2678RO2kXwwQkaGxCn2+gmf61avhSH
XKr9a/QiBYUCwGe/DH0u6UL5AI/zYnP6RtnL+0cDDIUT5MZoeQaEp3BNJPRrPZrR
/HXtQZq8uvT/r76jVIvL0QywvkPziJIAhaYdrQ0VaPXcGvtuy2rPlWaDvroHy6yX
I6CIEGfbB2F5kQtYegEkafKvZ5h+1PyKxALLremmGpIp7ZKZB7So40/wkxXtIcO9
ocjr2Mt7/sBFv4CTot5b9oiPz5k2m9wvtE4i2bMtocDjTDCNpiK62pM/DX5CUBvq
AER9dwMgMQgg7gzcPK4IPjkXkEHNkmdOC8hXlE1zJywoC5LYXJEmIJwamrs/gCgJ
1yohG6UamV/cspwst2cs489CFsJfNFwpbY7hjjWTDgSSrcvaWpKHm5kQPGWSXVvb
FAAKfOo0ZVav8eQTHQCizUuTgpIZQR8iPiWcDx5I+R5o/0BNcHyUiemue8qVv9B4
oaWI1yFOYcHv2cQEuAos2DT93tjF7PQd59WVlWXSnRQppWy2bcNOydndE+us+Dqr
Q0M1hutOTXUru5hnTdFk4kz7tnzejrZoPkXoMiaI7GOFj8BXT1xWq5n4R6CLa+Bb
QSzd81DTDAvB0qbSzuYsL47Z8iXM3AxpmVxrwOr30CpPI56jksttZpaZuFCgynCw
J3sUuenENmeoNNnwvdZRMxtqPY55BQmx2x27Ui6EyFSw257Rwwho6kS8voME6wQi
I/IROCU4KlP96Ku7x+5dM07lQGT8KpO9qV2+UmGwoSj+yIK2XAP9vK3kuh6gMklO
nHN8TGEokjyYbDOSZg1HVvYsw/8YnMPF5DDD2xaBq2Gi/Spe78pT+ISbn0wsEz5o
sCpEbqmHnfDSQV9KHtSpNnYQLG3dcnOmElhet2oDlhbnkS0l+ED8yOzRvWi2kUcI
7BoCFcphjgoRqa7QVjXZocHsVBtnCpIwNLXYxo4v1dF6jG3luein2CuZ0yiC7Qgd
jg55jNqokL8/OYSdQcP5p7izco+uuSw0ySM69dCR8m78sFEKPYGdyEKjpMDqPGks
TKjxECL7ZECe46o0MZq23hdqTr/Zl7IO33Do3hHplmI0/Zrg5BhAfIFmRrypHNxc
AA57Hof5eheocP80EEFzPzMFAC6qIKIkpgpPCGegJo9nTZqxqpagK5OflI6FdEsM
AhLK6oLoLlzkqS3O1yW/q284DiyNbdPwZkcom7M6Kezr5DHFDdAcujn0g2SKznhH
S8Sp5CailAyoDa8C+CnoYEJgoyP6oHqw+QULtcOwcljGNqK/aP9v7ICC3UaSuJvJ
zlyVpgR/pu3RF6JPq+8yIYRHJBbjdGKTX1CCxZ0oo+mPWv/LL0M/4V1GmbjBdLVC
sohjuLooDekiF1m/Mjk5Et3LEqRvAWGNgZPX5/Ehy7/QZjyESxEoajMmtzZi7z01
rgwXH+Q6gYGs3ORphE5LzrTqYRlPybqz4SZrojbKRMsn3IWiQ63AYYDOHBxq5Bzc
9cL39jr6WqtKixV1R7B+wq+XCh2Uji3ts7sn6FinZo1WyLa35ISjncbIWuxhZckL
BRvnWTbe+Mo/LEdTjNepV4FtnO8DIBOvVDF0PLXOlRVAiN46Dbfui6QklEUZ/6AH
s25SNs4floScyc75EfnsclxPNhxuBV048bmPHGKBOAl79M9DPUmmX8DcQCFyqkCq
EHUaiRwEvPPaIzXpphlgBUWtKLAUWBn02Fu8ypPw/PNzA0WNxqnuXm4dpduGGUr4
R6BBaSYHpC2cL6c9y4feW6HVhYFJjlF6bjfwtgEG1dITFuMpVBY/dGjYksFMvuM0
picsTJrbN5sEKlRTbLvmh7VucPXTeHBR71+xUNGJFTewklmxE8VnoNdLcqQCG3PW
DA4fQlfEV1n8MYk8A9hrs1R8fQ0IBAEPlwKj4UNkhVOddAhuVz01plbmiU7t7r+2
nwBLmr0abztpn6+UP3nY3Quj+BLP9DNU2TzqaBapyfFJ5o/Zfa6U5b9bntsIoGu7
sKHhX6iSo1CDAXPquJ0ast9vZ0V120S5/9kGK7W9uWgbMuD0/Kn2m/QYy2KdkcDT
jZDr8dNfB/B5TMKnbtbj+OMVnGlkA3E/AgooBbiAl3poG/R8bc16IzXBkzvj+u+m
pnMILMUAudO6ecTmMyII4pnqM9TgmNBgZ/rGdYH7Uw8Ajfp71f766q02FfN0wZ2P
up6iUjIUiSq0IWpyEJKL0J30FAG0l91XxEB9F1+4yNG+f14/SDMajv3rVX/Y0me+
89aY02YVOQXzcDdQaUEYTRR36/hs1OwF0JlC5ImGvqU2XAlSnw6hoiG5+QAABkFX
4/daPOYddnO02foD9aVSf7OhvN76v4YuCaXAmOfI+qhEDnLChCYb+Gmfr63ryANt
DMjxJ8jjBCDOMzreQfceFEl2TSm93aKe6jQs699oToIIARTlhVh/dssqqTgZ2xjb
kh8KVVfAzJZ0XF7CGp1WrumLWFvJSPBuBTfLl2uVeTJxb9c4UTCPScfGCLuXqr8T
Kw2ad3HqIkQQLJk5R3tPYZTZWXZI9wDQgzgDHOjQTZcHaXzTaddKVwJ+9DUVQMHr
ASFbwbs2Cj/vXt5RSc1LY1/x/PmJOefKryaXBkAauUxCRCJHDwnLYYLLtnBWDu69
lLv8p2S1KaIS/F2qkE0cLXoNoCRB9xV5ZfOJ9RPghkWRqcqmlsAQFIKQpFh28qs8
rkw3xOMLqATjfBQaRkMy1Cgo9QHC0K7FRCeOP/nJD6F2kkKomI0NYDTdtVgdYFK6
cwyWREYRib++gPQ8+ftMYoWB2xo/fmLLnEjhWd8FH/LNftk5PJ3P2RRU1ksDKfyG
sg1UOUPd46O11Z749pzvjMtZrU3PgY3msaSVD3WhYWq7NtTTJME510iB12lXb0ta
feDsSkgwYE8zPH2vagI1u5y12+3a0JXNadUnQiYQjcP/X3lknEzx65ntJlq+YPaZ
kN4Tv8VaMvGGHl9pQdKo1nvrwPZuT/tzkvTkfaObeDpbEddJrGx1KIQHMbfJe4mv
V097q0rJVhes87SnGhrzv0XLCO6+Upt3+TCgeWpKtDfy3Ge6+WyFDXuU60z07IRz
8Q35KMZdIenYPBrsD0FXK5aLR57OzXucg5jTwO4uIW4hlkEThgkIesAlSrES5fj3
ERRg85yYoNIbkh3JRFgFdVBbIaHh2m33JOjKrG/nBrOi7bC/xSSYtB8v3Kyx0rT3
izVJnxKhuY59Ogth2CfNidRKZEqm5i+fV19sbEPhjuyDdE7WNBb/fjSwDnf0xN9b
npAo1GjRJQLgH+w1vnHfHuDYKzJmg5IWH8cVUC5IEtWuE0UpSwzJ/qrZVEvhdc0h
4DQOqHeRrZ2JiQNgv9eIB3ZcO5mhT+SxX99VzW95/ahUkTEkKWeLKaAKksg7nem6
zZ5D6cDsHg5+42cdevNrQbzL/1hWG8q7Marg6VbWHEcvJclDMq+Bc5OdIFSw+IJ+
szK92pXrb+B3ElppFF418pglxn3073DKLiFgBbwKtZAxmD9+6liDOo5JVfIem628
vOClOebKFiGkM5Z9hpcaxtBZ6zWV75W//K2k8D2jQvVkm7g8FCciNO+JI+M0CR93
Aww7hOBUR8sVGZfrrwDTnZzEapBOg76SSBFdUeFGw0KND9gsXZhgahCNK7INSUcC
dL9/bZ5PihKmHeR2yUG5Qi2/oPLIWtb3NMmHxG9EFnHMAwUkuNoJTGyb2cYFBKHu
IH3z29rf1d2jkaVIwAYDZR5adnoJrd7OogeCa/RhN9UG1oCVUfKLqCbUixyTuPSG
SRysBBdP7eNj+VRWbxirFSc/ufporsmbHjmOYHLpK0fhSJp8qwp8zNn/nErGwLF0
AxTBzGju/qoUCqKBTZo+2zFeYcOY3zkEEhYDIy15KeaNO2co0Ob6F9aatCB8GKwR
ARVg+23UZVaEOXxBHItx4kIuYGSNbJY0oLURu1pX6J+KFZac4qPjWZIwoC2AvAPU
Ce+mOHhhoDd88G7STErg7A1ByGTZhX2xfxWmaOGUU90dZ9b8WEhh9TjWDixNxzj0
49IkYzLJ6zQd79XgWVpB/gj/R3ELGnQ229mnFHVAtuirTYrupncuDdCMC6WJRCgu
nBOTMkjOXdykaHS2URdnHKVQL0ldnxr2zgtuQ/BPOaOcjZpud0oePH4TEL7PzhUu
8M58We4wPl+DVueiEKx0gQruMID7Y2cdAcBZERZba6/OOpCxU9Uav81fTFa6cXRN
m9sulOm48X+AvnChoGTAeNejiiO/RYNQ+UhL94cIWVYy/LRKsk4Pdg1htxYRXBWp
ktH3r+Exhj4N6RY49X35qKumdzEhP4J66YPZ61xL9br/7cvDy04RqZ0lu1T7eAFz
R216mQEo5gmWPRXN8WGQQOek/spZSzpCuKFXin/Nx/UwqBnP8+2u2AyA7W1On5ja
k2+1eSkLcRTZpDyMT7iDy7dEAN2W8o+5e6ykKXmQIxI8pjlhCfhb4SXLHDgKnEDv
J+LTu4fVK0W7nzYM1FJ0k3D/2wshPLHOBOHnFr0MMwKUM9EFJjLBS+Yq8aRupicM
fadaHmqBr2LaT4amhJQhMktL11GbdgEyPym5psbDYVTRZXOkTVsXfPShAg/DJcnQ
OfA1f6+/TSzESd2okKdLbkUfIDZajFHVf/cCdfie1xBr5b2qrv3Ao1vaKTl3wdQj
a1Z6L1SV4mV+rGHYLkZlAILId9tv6uwGL7clAu7TNaBLgL5YEf9Hc8C5BQeUbpN4
CtGKZNVBpPgNZiwlip+4e0Ch5CH1/PF4INY/Lz33zJebK7erug9cwT5x6uhTPNpL
UiJ6F6WVN2SFlR4aMKA4y+v8ajkaePmJsQgfd8xtzyXe0k/+ozsXnJH2vMweRxLW
rZf/u0NYwI49gPoOklEIOuyI1qggFIhaYCNquGNJ6KrV5g+WIDieLACOTx4WxD/6
ZgSaJKJXPT/e2gsN+VqhtSs84HhF8jbGGfUe9X9CqNPnt5AdWNQg2+BYhnEdAk2L
B9oG3iiROG1fssW1epHuLL/ll9NG7OZ1LS58ndm0HauBNvBwcyQ1srFnb30Bs5Z1
XhedMrfnkU5jFVKkvewiUqVGe+aVaIFf+rse7WWrgX8cMuDQ2bbzJ2/TVTeYkD7/
yFScISmy3nXlsUb9k2KPK1RZWiSumRNKeByBRAYbJs1ye1VHuyVGgObdObTSOkrz
A4BrtTziRNZ0YIkRB/oQd3GS3X+XykfoTbURW+/vK7zgzBACRh88EAPv60La3Yre
eN8Y9WMmYM1OagBPCXz/5F2hoY/gooq2qN4aqvxVwWWrDtpVt/7laOKE2sJw2OTy
NhnRqqRSN7/1aFlOZHmRdwRfDDSK17IOBVkJgrzFbEFJNyYtQEx642/ljtIbATvE
FDBQydePKESNza4U2Pi8ljMxepAtz/jtQHF4aJJtj6TdwFsj17gIvKRYPM+QlJSi
xk/enaSjoy8aPv03/Zj6iaQKzKfJWCYijN06Czl3CAqagYvqWjRKbykCJNOIkBSL
oCoxssCNcRfhxjhrIh02fhI8WqGhdTr+E4XentbSBoZmHuaHdsKfnSSyjYTEXG5e
K5zacHEw5PgIGpL+fyubKoKyqQYfiq5turKMtZ7Y9Si+L+9OUEuVCf0j3zJorgiu
hV3+lKcmowgI4Qe7+R14jSdeVU16Wq3AEG7Fmrl2rNrMzY527rSOsXIBwLU4FQ0A
gR7dyBER1PxhlD0DMemYCkFzpbtEiD9Qgd7YUdZyIECXKtqRdTTHTWFIsm4AKGs4
imqb93hUq9HxD2QFkKjS8NqIjqfBLwJhCjMImy1cri7uO1hZCa0vOpcpcuNKJM4U
BYLr2G1BSP2YeRv0tV55lDmBKL4oQBG69E/nscX3qxMLQtTwQLDRC5KmZrKGyGA+
X8IoX1pShSkIc4SAy7aGmsDhFsd9VOKVeGMTRi6l6/4tL1G6kCz+Bnx9Kc+YtyL0
OFPW7rSYbQUJxlJJ1PeUjp0DZS69+Js3EKO2VeDQgtFUDyjKwQHsdB0hh4yjwqvZ
CPYpU+gPWuRLGQh3FXVBgeOBYnWxS9B6uoZipsmtJecBnqbafewTeOam8lyyCfwZ
uDgV53NV/Bc3rEZi8VuVFm4rxarfgCoZJNByd123oSraED9wrKZgMPBMXJ7EE28V
/UvsNTuWkpMaFfmz2+w/mGW3XYWRgw/Fgr+NmbUmpelz1DWAzuyfEd0MWj5f89+i
PyWknT3sVn8mGlK3Gaa7M1rnjMmDoQ5FUe13PHMwspUV5T2ihsMJl5uBJI5dBi90
NSn4kssX28VDDJ3to19/+JupTzQLq9V4qykyIdXkUXAWYHb3NSlumPFKv0QOANe/
rHrgxVAPlGkwi3lSbdrpVnS1Ggb/VkNwPNlrQoXvH6SO/KqTm6vFrLAZwQpLvIZY
YobDDYVN+h1I5T/z0tcvZkWlbkRjcHz3I05bqrEGCwdEzmU4C2n/aAphrRVMEX/2
JTZR3LVTCRL4sj//dGeUi/mU3m6zYyLcY4DZ6pBOkMEZh0TgTb9TWi0Orzs6mQyQ
Tc4hSH/E18uMSmkx2g55MgddkJR5f4Vk9iLbWURR3e0aDxxkTjwN/AgceIY6p6by
59cgHuFELE/BjqXMb8oNNcTD53sRlKx+fcBTENx3vB+aYILTjWc3J2Vycl8XDmRl
cvQROFVPTa8X1u5FPkmzttAQ85IPfSkkrE97uNC9HERxwJukw5kkVl81S9NaFKZL
j3GTwcKD1WRdRV71H5CpDp2utDYJ2YIxnf7GQVOkJuufwXQMj2OiABudeEjJ1Lhq
/UsvMLq2gZ+8FvYVz8n+yiPkoG6/Tphjh94l6+SAb1Wqo63NNbeG+qF/fZHXCnd4
gCQpxbynQ5VVVo5Itb0pYX3qylSUYErmt8Gjxukufd3TZommzOYr/prZyJs5JH2K
/t6d+2E87vCuet0bL9fsVIlgLJIE/tsST7/WEK4XHeBH8oMwWxGJjwL4GKdYv7lC
qhN3N+jSD2fHUvHbw7zbwVxKwNEsGmV+fqTodUqgjy49H+IW1WS0OFqQKg73eHXH
ruykLXFqUg3pLMlbnmLUf8VyFDs4wkSudESKFf2c5tmnEPuCOFKc0CvL5H1mUZGP
hrRqPSsNTPhKHJ4lMgJQ4Bnm/yW8ffz7e7WZANAxO0ygX1uWlqUzdJJdktj7AthG
SHj3JMzNq3ST3bLZDK9xGXXwOD55soCnmGW8O//PIAGGVHdyJ6vH0L6ybiDEdorl
osD3g37fxrLmZ3WyfQAjhF6t5IG7HlyQ/mgGTxXa/IbyBRCc5O7fvYQC+jKscmHM
jTfTZ/tPe7l4oaHUs3MW25k1N4QJSV7ARzM9ZY5JEeclZIsRHtbP+1af0VKaR0QN
UQNejr3KyVqSyJlM+6kSNeLLZyxjwdDi0FdGxqkdaLg/+DYl5C8yCCLTnWNle/H+
c7H+Yk3+NVVHOvh6xHhRoR/AHU4VhhXVeztC9qDTv3qqMdzObzBbjfGug6tMIU+J
+eGwZG/ZGTI0CMCM6mqpo5cclGfs4NhruRn2PZf0Z5IkUGKOrwTwyzeZWwH1GVsw
xGRoF7TKocKgYN1UpUQy9a+cc4vvz6pVs+h0o/g/JxZrfr0Wr6TSimZrq5AmNMtP
R1glzd/SZDOMbu1KxKHrUMuaXVfVsZBZLW+yHDaFuNfYRo66WFamPzzH07Dus0Xg
PsmrIagdaYURJjooryXnI+QVrLX0g2eZ01AOs28Am5dq9Pv+f15RM94IaIQJQ2/e
bZniu7pMo02BPub8ZAchqT/lDc5qkPr2r8P2jPqGM9J2i0mrxWrmPkJ0mXy+KDKL
Z46NbF2cL6lEOKYQ7zUmhn57Q9Rwj7EMRR5TF38HrlYI8K1GjHXejXyPGVsgWhRY
1KDM53ez2FxS0QFCdoHnikwzyhsrU/QXgpH5kYTiraIatYIhynCMxiZJy3KmjEd6
s49Gu8ME8SI31TpN9FbqC4EyohTqUMj+oLrnk7X/TumRKnVOfyRx6l8VebGdfaYD
GdoFpCX0It9UVSGKc35ZfyHURkJfr7DOFe5PjZjtCoVSqFTer7oNm7h6geiuEMpL
4414380oqO6INbU5gKyvTaPpbc43ZvDljU1a0l9+Pw4975wOltruKZvu2qgkctaW
TTaUjzHTlj7NMPEl8/MM3i8Q4MeCMUlk/KiMoDlPivdLfoDCCUpOUpr6BfKJhHne
Nc3zRsfi5dDX52e8oC0uLhDYOlUtxC50EcLQ/y3nqrVL9LKHpeuvvQdNsV7VdJZa
09Reh+djO4ivghuPQnGAJaqFK5aYyYkuVXy1axHP141R0r8tcbvwI70RwnGfD3rx
1vV8jJ0T+xqVYAPClK4+MKn3wquvMsw6wDNbjssdqmoj/MEsIQKwbbWWH0Mivt1p
+BU6u+VkP+6Gb3gIsnAQDZztLra/SMkWQcP4944Bkx4EC9DQW5WCVSF6QrGTxWw+
0FlCjacbB7QXbUtGY2IzPwuiRtBXangEvFMvIq7TA1p3Z9W2/cN15KBTGBrlS4BB
fxg+7skYTAhrbH46ZysnWUfXPeWTAgfvSi9OR/vxbpISYIq+FL0sNJ7IfamYyRHZ
Vf1YTnj6isFrPqpF8JY8zTW9cpqhxjTtrTWcBUVzBqCE+uoCZkE771DJf3Q9zory
kdJ7FmOAuR6Kmtl4+zrZhA/hXHoWURr+5g0jd32jFB/aZRvBf1Z3pwUI96ZnOldK
rnD5YMZfghNHkCkJfemgzI6JCuVb69ccbev/f8UxhIk+HUZxqFg+XrEjdf3+Uikk
VynMdlNn2axhhx3eWmqMS5XCZiQmpqXrAX/5LEO8XTHm1Saf66torKjcCMKs6Lio
uT5EPjVvfj7XNwEowWIVzaSbB/aBdtg0QXs6vamWPKM0ajRLrUTKnwrNrF0Zx5qA
FHtLxbayK6sUOux60T9XLVGCYpJpy39iZ90FfpQYAqjc8yricqSeJUrDnFYIpXqD
Qzp6rta+9lbFZeYLU+CBshCPsoPSwP4tOiAS2AQdAlS9EjJWOja8UUxcEjIbqfzN
YruJEGDn7rf1LFvMzPPCRNKZjZW86Qs1QXnBnjVxfIxNuBl5qmh4HpBlHXDCfkor
dx3Qv+pECe+SWWQmxeJ/YC7vdp0M0e3zM26fdKoJRUWys9G5tiPJ73wmLOZUxvhB
rZxhARrlmpNjJAcetYFKE60W0cEG5B7Ftqn2CWlRJnvyZc1J10dQgZMR3shRzNY6
/kgJUT8qjiZ6GXExCyRZw1fVMO4N2zBQn4b0BBh8r5NtRM/8bgDrDohde5G8zRk2
S0mMZ449/rZURUOAVsIbY966fvLD2VAL1WW3RSQW9qXI5O/wQbVLRl6GehC0h1L7
aV3QjU5p6LM7FpUIBTuSJ2S347DY8We2PHf0S0kcKe317SJMR6hZOJajzX7ulCNq
7DvglGPDrVMpHs4z7JCP2HeP0qRrhE327FbJtuwtUXe21s7nAHEZd9aSnUDPqXOR
IYA9Vmme7PPa9bwFhICdXtHErJRQUXIt6qBqWOQizAj0aBDnfueSrWCCUYUsjrCx
F30rm3/mKfb1S8WSiSX393wKN/4SwweSR5tMgxpzHVMe6l73ojsTU/BP2cQUbPvl
rhKiyIjOAjyvEJxiAVdl4hm50guE3QAfun4rZocMdKefFxD6QUgNEm21ps5L3xza
7Uv+YsBwF21MDa4UCcY9SQ312n+TSDLnb+GjjtTElkuOK2WbyoLB4vu0tnyRwXax
PPHE1nDubejcg/I3jk/LGnJbGCHwKSpNRcdrPX+fVZ6ij9RBXciWRXhR8+C62pYM
L0tpKPj39yoZGcDFnf4aATI0yb7aNJF0WYeSbomdG/5BAA/0JwK/q6ioaU8eoUdb
YHG8fHEAa4y7a4vlZqdLLPQjl60rLV7MGWCPKP8lYtRofOOZQsd0m/O34Lpv4kAs
4k+hkeqJuH+zuidmkI8rSCHI21rmOw1H14q1oIJDvqr+9CvzsJMxPkgbMQguCC6p
u/foWbFJGkFjdahkWUQfIj1ef8GgOk8o1nvYyd9W++SfhaRCVN/HEIRGYVWOUb9M
TJ4E1rJRxfFFxY7CqJSeaHdYeBVimQ2xMvezxvx89ibONNtDS/R2ub7vy+Lvs7FB
Wm9DhN2JorGL7PzWe56QcNeriiY/MeoNV2wBPAGtjGQRpXrSp4YkcgrFz9mLlOgG
ulsQkSeinSoVeLOMmi2kfNFdiM1iz1jJZvuc2RMMZ/YbUu0sqYargFvFqMFu4O0Z
KQ67HNQ6/j5OFwdoZjYtl7Jw9Ls10OVx8B1puVqNvIdIZadvF+VpEEjO+cFBcBr0
KxyDSbohhw9tvB7byeQyQf6mHxuM/EUPaEzJnh0NEy2Q9DGisMSsdfU8ryToRgTy
HGFpkNsF7TIU52IN7nTee383Pp4irHHfMWCUW7JTrRWKlBRm1CfmIAh2XEtf8NCQ
m1YxOYTAJqj0emhWiBYCEjDSfXhSWuHF7IRGasiDO7FdqQUFFImFq6jXwjdO1wuq
BLAIl73qq2BNJu9Xae7fe59bXv/wd75DbFF1CmSVkrrObiIj/eENMhLWWGkRn5Jq
HmASGchFuOjS/RYwi0jGnDX9TgoRG9tnJlVlcxnEwW6wSzhM1TE7x/yaPNn6kn0a
cHDRT43/l7zKc2TyRzjZVO4A3qpsbQ0w4Rzw3yB+BezHbc68jOXeDcqZK4GQjIH5
RTa4BQ3C5G1CafXa3fEv08AWp39K2R09yiVjMxymsJh0+MoQH9hq/ja+NYCAHetN
6LLAprP2GzdIzkbl7E1bvrHCPTd/w8vVy/qctGau30XabvjXfin34C75j1iLynED
tniLyru+YWyn2rs+ITugUIdjI7K1naSMt5hhKp5Y4OQkiOkkfDy51yb7nx2VtDWI
E2Oge2W2cV1NLZ+bfeiazcm4soRI84AoLEL7ed2wUi5lGeJLq9ltOM5qavYSrI4m
ScykbqJpgtamxBVm869XVaANGeioJmt4/UlnynZIdKgQeefu8II8gT5ufrjM2VKP
wn1R53C0jLadgJdnFLF9CePKFAdcrC4eLll6dB1t7+451Mu7Oo6ZU+H7usocU8iR
AUDssawlxTQrfPTrb6600WNvWhpCFJcbEiUajXz5B4oAcWyLiHhzxpifqzK/Z3V8
kl0ELakC0MgYTuMOqD2lzvtFAqDZUGCdmGB9N0UxttPpJcjzZe0eyzO+3iY26v7a
GTZF+m20C1OQU+KjG9Ml/wAPQMWX9Ujl91IY33vndVoT3CWOHNBuByDOnD0X98AL
eF/pqm10t9GM3WXB/+5TsuHTG/Qe4w3FLYSoSNcOWP+69KjT8eIRtNli5eXiAk3a
etv5WI/98KOyOIqn1oCQ0//XxZk6ACjJLaTZrGG+V9KqMW4VTiGGyQw+lGXnZs+e
ox1ih+bgNo7afvCT733cSbEOBOrxc12wSFPPIK29AW6Jr65zI4p5/8tIXf49kqQy
pflmceXh80EE/kJjXyu6noqAI+B0Ts5lePU6gC2ymZUPRElCY28Y/AWReRXt6Wig
BrpOfRFnBfDTZZ3apDu6klGm+byz/R7teC32Ph8IEXmlO19DtJdTRpMnub732YCH
hKMBEpvfc6XP4u19V+AhArxSEIdht/O9rgKQDd76w51TDNQFdxcmcAC8QWjZHux4
ZHjBjmo1U1PJVidl+jXG2QwT88ov/Re8Zpp2hnSUS9Noxxs530BBKPcRaQkA05gf
0loLqxQVx1++kOYjwFW0AbUXPoM76IEU6OJbWEILhTqKUhmnLBzuSlv2X+4fGjZY
Aa8I23wrLa3sL6vSRkPAi0m5CSFojFJZ8dFqoackg4EegPS3D613DpcxWcnCQm8i
Diq2LxFA+tIvNL046WtL/StUNyhZaAgWYxu0A33LS7MpIwzn/lneN4Y6nO+NeSEJ
xmOpA0+NT7RTk2cMGJnQ1Ckb4BxYfi46Gx80qRzbjQY5lWvKalKmqjK2TOMs9mR9
taqTNBxdbdLYxV/1sVTdCRTaRFsMYfvpdKCkws09ftsfum8BXpbMCWRDYvaCLM+V
znJGvDtL8OQp4EVWCTNq3JCllQFta+eutsS+kvvM7blpOstiZw1GYENtAVZ/MaOA
b76vDcKrK4TrvAVua0h/2AsqCSQjpHTCWYf+si3C4zQjzuHCK72lIgAq3BA93P2H
5LgfSGnKghy1ebeIYp7WdyUquvUjj1MqoztxByjvx9IoF/7o7O1ffH9pVA3wNQMo
sa5aPsL27C+Cn4EXQ/dzbmvxdBOws8FLPxVuP2SflCXhQzfu88Cu6O21ze+LhUp/
68rhkGQDvVeO7URezRz5eRkD6BAxAHWPuT1/7cqOKjdvE4zJ3//1orhHfqHhF75N
GZ5JqmO8pgYWAVhHtdmItFlxQGe5Y227d40Vmg15a50XrXkwepY9yffZMF6uRcoo
CigS65kpLK3zdQVU+UpVg8UQ67hAALCe563ZBawIy6dqXf8M7AsRusXSxuHopstJ
lb6Yq8acdM5RKC0BZJavO/5rF7uZCd+xD2BYJ1ujOsTMGpaU0dzgg7Sdgsm5/E5I
gmG7f5yMlD2xam6Knui1f9y6Nf8RXXoCPJjE6kmV1w8HdcpoRK6ayAzNyfjdvSf6
i+sD87U2euXBsc4UowDkemD8W8c9gYsxgHX7XwVQgiclvjhVoDtkEso0Q0i3vrZr
/3lgCN04r0hvJ0D3/Lrd0fsWJ/TR9L4KM4I2vD9lWTMeSUw1nKlJdk0ecP/fd9Zt
vrcqZXqmEtLiXwUtcbtmZv1ciOH8fNGazyIs60wHlgHRKX4wd8gp5DpDBVDUulGF
zQNtfsnT6GAVSVNKApt5ETI7OZkOTXWOHUTSQSz1Etrop0lFLRNdlHK+RLIKxEsP
HgWcmF6wTGSNk8Qm6sKDu46lomEanFZ/nVwiOrgdD7XsgzRIJuO/dD2TBdRMf/cr
ki+ehAfy93uoZf89MswD6KjpIh0xCo0Qe7KVmbOPxsehX9C+pGBfd+XfsHiZiW4t
rPTPRRovZZYOGUSTGXCRP5puHmAUIt8j2dr758DxGjIRS+1cyK093BWF3oIMahHw
ybFtiKN1dkD5E+3/pnmNLsvgjKCUvuSwdUq4kmoK8DW1/jqlgzleqgqNhO0y3Zn9
o9hD7okQpnC9nmx7e0uTq9Aek0NbsM/pgabNfXRAzO6oh7CFq3GeuzDTuFdnjs5G
rcyWdGnQOvswSyHlZI++g70dQACRJuuRcG+dNrnDeoU9LfX4Q6cAIQ282Wpb984f
XSeP3QRq6Pe+Mgt7+pFo5LZ7LrI21m78LspNdIHVFRldRSptJLF+Crjp5E2m+Xdm
v/I1cVyAGoju4e02a946I2tws4IJAAD9i5e64+cf8Mve05pO8AZLsIP+p89e+0G5
8omx/eeOZ4W+x0x9TD1pqeHj1xZnMiyqU9+JiBS8xz9yxC6q4tksY5iJ1sZwnJiE
MRE7DVz4d2YHYa8Pd92WGiav+yaAr+R5MR0ACv2zaWf3CkQCwu0ccqILciOita8B
hEcJpVv/yUPfOXV71Ttagd9la6Kl7uwXDX4l+y83Xc72MRV72urno9qKqZXSv5BN
qg3frgC6tulJ4/eqhL6yFpVjFJlwaIi4qWzP9Ut0HCuAT+K3+eTn0T+kF80n/Agz
1VecRONLM+Ss7ghX61Rkkkkj1fLWze1pEAtLem0PYyDiX6aPodW/oEMOohi/JR/g
T0PYCKimwWPiM+avaVafxco8V1okeghEIwX+TPVItyZB8GoIrMYv9iv/hevh1sxo
ROny85KdHJbEoN0rztUIaN4TP4K+E1y/uoIjajtI9yjke0Yoce74VDVyayHRiCD0
4XdtppIqHZEb/DsjF9rMao+gV6Ef3qZkzjNEaHjgTDGot7bVgiqgtPgNngpj002/
/0DcPX9NWniOMwc/CpQ6+IIqw9D3T/nQiShQaonGifjTlYPsFo2s8HsUorUFkErO
+dRX/d+DpYpjcTR++2MoC+OpQijWqrsnBmVH5vrPhyjuJlsNbGaQXZGFWcgwJTOW
7LRGREb4Aluh5Cp6BTIKAQDhzDYqF4/NP62rkvmv/63RPkuSGu2G0pxKUaSE+jAR
uLqmY+SeHvHlyIdmiJLd2rLNhCkOh7uJGU4Kg7NAjzCG9foQ5DSEKJLtfZ1bk7BF
jDR/3ZPdRT34Cr93IWdXHCt5/A01uI4mumWHXlnw+nbtfp6IbL8Dq3Nn4dmq3UD+
OAEjP0leIxexIho9r/MfQug/ZlHokoYx2xJXmEMroQidmEwXYXOFIZQWQ2nAw2xn
5s3hGh0sw6DFNV8aBTlNHR19k4WjoQI9bosBbEbI/XEPJOI4NSJjqEJfNUZqdGPK
TDZCOM1TJeFCoKomD1FOK3W1eWlaDyaVbeLgPy4lYC5+Zv+Zew7beBxee0tfuLFZ
iPxGrVIsIrPCvZecZgiYYSnQqFnRy4IVxQyFTcq2HE6S9Y/UUCyF3EqxqIh9cqYp
xK8Xe255t+zR0uPIB4xs3amXlt/1qXQ+Lt2gC6A27n1P02aqsnVrfPJStU3Ks3+i
4RPCIN/T23R79A+XKwv+8JhDl6ljIr66LmBAGr5tozlifz3CpulIVkBFDBJvica4
q8imuUWkY3rtTbD1DLI++5qVoVoI0/DvOwj/RbjI6eNWEkqGfkGdygae3W9KSMdi
OY8c7JrI1pctWibsQZflPUWv8L70E/+0Ax1ARc2XgB/t+trl94K9DQbCqYQQxhEI
DPt0YlUyIBlE2xJAHZRag0DB3sFzUaRJOZa/WzCq4XjBWcPpV7ozDRsnTFVOAako
lmHs/ML8IGWzWM6WllIraVGXCcpv0LRswVdObVDfaJZxcbj38ETDzFNIxq7C/Dik
9BbY/WWKoubPgmwRAnOt57h/WY8HhDfbU5irCkkWpth4ZRhMhV6eSRWOQHQl/ax6
zLgizCxYW/DHMiGPy+zKQHXlhmqycb/Qxz/eitMJoIyLj4uvGcPDsMm0uFa1h1OL
uh00EbqrBIinpNm5IEe1VOXd3Ot/98ECqx7UOnGUJ4FOMmXxELFUn4LfhPSQ9aYI
0cIwrzsGGQ+xTDphlG25WyW5gOrhLhgW45Up2hRdWh523xbhtU0TYaR1nUfKbITI
38vd5yShxNbeuhr8kyCJxyfDEvrOm8uxM89dOLdATEf54Zz7kEwKAZnOlo6nTXjd
4kxhUBhpBuiO/fHSDGJ4cQ2BNN49GyhSSPo80R8CKAy3DLGpzLfdE2PIht/6vQin
qcfegzHsPHU0KaWtb5VfHEkSf33QHm3PLI7IEHm7Fdjwncs519Eo1r7g0fYHD2Zo
Dx13rhIZc94wNCo/m6kYXsvaEl+I6A/TjIlaXYqdyu1Rxy2HnM7LanHC9Gl2Z0z7
aoi95jK2PD28DYeJvNGQNmNTJtmXjpZVNtse7QrYeWOTb9N270HJkIB0kPwRn34R
SQp86rjr8QrLm9nqlWFo0+aLdblrqKImv3TNpplTFFzz5vClVntgv50eyaqWnlTh
Dp/R7e8ZrETJtOAfRdSMRNNG6f1xgQJrpTDloAhaZV2lzChlJWbJYaliP7DElIcH
iieURGAAC0puGtP7s8/bmRCN4EUt/d98dCZ/i5MJK8Tlx6pJl2wMZ+WV02PETBiB
QohAc84YgPJGQj6DwWBOHP2HQePDIf61zcirlFdlkzYDGLrNdFfLWlGWVP8niAdz
5aUWg195a3A7y63ZqmkaYj5mByMxAarBKzbN9BSPo8zbakjSwBsWleVGGpIPUEEJ
LSgpf1X7j54wJq1baOSbJ81BhdX/g7nwvK0o8BB8QsIhLa1n4mP2vwVGrX8Yx9kl
W4ctWddrLTOX2WzHBiwY6FffEWTf7moXXblBHwf1rZFL5ozz5GKRW0ZDVbzPSMWr
f6LId1y+Oo1bHgk90rGWyM0lxKY+PtQBamIugaWT/qjbsu2RLTvo2FZjSvhNkN6H
8rKv77YNh23U4FlBGK+zIrh9mq/4F/qlpo3GH3klY63NxWVy6TZz7lpIWCJGs80R
DqV52wzUIsbUapM9PtWxu949AdOGxNph+mBUq/bR/Cxd0Jb9AEdjyzVlJ8exiRvf
yyJHQUNDPyKQXvgbGgJ+hlvFNXbxDmErJZz3GAbsE4xusMdzrMFxpdHE3NH4Tjoi
TAVKVpnbCUK1gOFZp0+Et8bhRd1eV01LEnUMPwBYaCsUQccRL+MVaKW9UiPOyNR8
zwFSeaZEUA+G7AIIX141eizfQhxYRcIdjxdm+Q4RDxdRwyfAtIt+xTRnSXQ4i5dw
qELGMudeMIFYXiBxnqN89JAmDhI3ABaesrqL1YHNNkfRpAjcAT7qTtUmJXg4nnUb
Mk/bAb6sziikUlwk1VQdpcUiImmhw8FLJYEDNCX0PzPnb6izAZVde0GXInOCZChS
OiQeqSQwdtup4S2dF3/lZEkinvyZsFa4lvB1TLV+NnIRYsptmxbQBSBDd0lB7h2G
ZbUikANZRxvpbP+LfuKDvkjYSuhoSz5YybrZPwTwkwzvJfH/908GraxoZfyNWN+f
957eDUAo41vwJtGhlYVG+PVmIJiGS8CPa/QYR3oVxXCq0o4xSciY50M+1l6OJ31o
twahPa5RtUi2CKJ3czMbwYwpyaLU7olaHgrB6eNOgy5Nr6VTSIihy1tMO49ygA4F
4HhdcwKHpFDnPf7B2jh86jlCWmuoHte3modQyaWyYG5393qKyXVO75bVfSj1ggOE
cmRAgFgXD6Ah2QIx2lzDopfFqWhX4o47xhc8vc3WrzE4AZAO5B4BjjvCV2jKWyrs
I83hruuBY7rrZgP00KJWRpWZLX+XmRtwd7I54oU4UYNy25g4rThjcRZxDA+eDSLq
Z4l2qgAgQAk6M0ycG6UbY0ObrXf7mjpcyC2rAmAVzr47AdSIg1jN4waFLrGATcXf
3WeXFLVvsaKR6J5F0M1f5QAK4QXUMkiwrol6ZD652CYh+0oaFhsUbstscjyM0cvn
3ybqKI+D3Inw8qDmHqifhzNePGTXsz3J4cfhCbuqaRJvd8Ye/IEQlL85WaaUsXPX
mMDSvwgEL9juY9x3BmGCI1znRLr1eCEKfDMSeNbHyG1ThBlEIeJoow6NLrzWAe/L
3uejO00UFrIF0nUjhbw+TwO5EPKPyDZVJKy49TJaB4p4SPCgHCTuvqY3dRVj98Ot
Yu9GrsvEio4RJNgicq6wtQnf+2wUs7GmoinCirEZIxa/UOO6M/FSHzq+fsmkwKit
qFmAyu7vwisXG8AjFHwP5LsrET1saTcb8yGeBkxYHwr3QkG+VhNL9xKdUBV06TV7
ZBhvfGYqV7zmA/hcgMTvZd9BXL8uadGXQZyFpKeyx67DGEM7x2dfRyA2YB6/I4oM
KonLGGe5ktkZIXKg6QmGe1FaUxxgLtpi0YSOPpFTt7QUH3YIBtsG2uRV40tOcSzX
w+kyyJHmL3QRPsfkan0URd1owi/CZTQbOrONuajhufoU5x39tsFuGStZIl9g11ff
3b02Mvj+Fd3gcM0kljFPdR12cpooTpcoBh6XoMTp4X3/qPULcLvKPR+9iVak8s2U
6iSQqlTOD0izc1MBSp7rWJvLcltOUwTJ2dn6NYz8TFwm++xRDIF/mCe0ak6+tGer
xwdPfvaUaqJtHuDkAomdpOL6XuqSwgKjAABHiLoW9COKGewdHkw5doc+rUszfTdQ
1S0i3qsPaD/wadYwdrzvbmS7oNIOoyPb4LJZ5LsHK2qOkYOBpXl9PbZmXzwXPJTl
fXspH62yo2ihBLFEndRRXCaa4YsoNwZgRb4AhvpLz6C7AUdvIcIy5zPsrSQdsFsO
S/UKE7xueHXYu4JUMjvEWCU1DVMj3cgwqFiuKWKjwNLdQPQSRdgtxYBL+rHVIdX5
BRGoEKOfJJZ6MX9F25q26ijlzyHzXQidMalMuLkl5vWnBLlZ3ycnBIxuylbkwD2F
u+3nCq4xX5pMb/3jdHi5mVQQ+ByPhljDrzgm4zZsuXRs7TLUsgwR5ojLpEh5L0iK
AZPE9pfNxKzsEziPMkB9tBTuCAwPm5ouqg+OhcLuKovb46s7a3L4+qzY3rNpNdUO
cQv5rtLqlBEgG+nfgikyQ6BxqMb8DP11yA2hDhD5eCD9un94X1I3UeZqvl3xJXyb
+9D2qlyalCVS8TIBBiNE+l6v9tkfU/RP/UCsx9iFXLKYmhRQRJ48fBwOcZNcmUTw
cz9nuHQGjf9Og8abf0vbL1XF2uVtat1ax6nbfdtIORkVyeGXQPfmpy3GFQucDxRv
`protect end_protected