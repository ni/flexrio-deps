`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 21376 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMWORzZC7bo0toZS2Zods6Xs
yljw+BvqICQb54hGe2JGpCy7VfzPucQWBxxbAs+GRahg9412xiERyTvngZg3x2MG
UakpXLdTL/MtFAq4zNxNHDI7EWcR7qfLYYM8QIuaFrPnTqGIdgdVlYdCVfFjsDh4
H+7lqeTW2wXKegY5f23ckp35FGUVvE8/Wb730o/aWqYkB5D+IOWPRxc9Mnj9rpI6
D+IXGZ7ZnfYk00/5gCfaTP0DIPzpY7DLUXSj55DhMTDp3QMn8/cVRYAOLwbH/v7Q
AA0P0ozKxFlVP9Ld2O6gvs9rQxLY5CLZzEnc2Tix1x+mxg5j08OIcogJ0B2J4F9O
a3Sh5qtIYd8xeQ59oLL3IQlXQhrAGT6YnIRyqNBM/1d6Qf6uYvFpMUtvcfwjy3dP
XuXS9YguY/PeIyhDd5A/CorQ5AjNaK+Kf0r1c3uIGnsredK9BVtGwN72UPXkrWdy
cNXXjw7t12q0qVkZxCnziwx6fQIToX/WauHDBuxGQXS8v4acbQn81C88568cmGQ/
L6A0qHl12Uz8guBxBUfB0ejr+D3K1nWkiwJ4L0PyP+xw2mdu5/vbkX8f1HHkTLgq
r5VyRu4jZFPMHNxrngkuBPSo+4Is3bsFo6mOAIq9Bgtdc96VpXav9oGkV7aWXpp5
M8d4pUJSPO3mJxSOA25LKHRApGl9Gdbbt7Ud+3nFUB4o6WEQzaymUOTaS3pR8SYr
zGqlI+xwVqzGM/YkmIsKp4ybkEYdLd0cPMRt1552YL86XkmWh44K3FzV/6nmKd7Z
+fLLvUeiEC4cF4TVFRmc5k1F99Z5hVWbgyQ00niiqJWuIdEtZJfKuiliteR1xfWa
8wPKBkV+TYIW15Q7t/jM+Rix7LVrgXuPsmAu5QVoL3xHEYNVspNnGkYf7uc4B4Jn
f+vkyfuo+fW+3l89gG0pK8Nqa+MxxUhTVGnVsCUGzV0jwKV2mBt9FZdwA1tO0SK6
6J4yJ/gbIs/fHfm91zytSZ4J/fA7H6WP85HoRhacTzt0DEtf69ZPDEWL/1HqToKa
5H8JAfx5kIuB5BV9lB59IBQJOipnpUHLoTPkL3g0ju+8gUmhgozwDIkPvv4XMkLr
eQr/QHfHc1HEpJY/ByvFxVGXJdqOLHjYfDAXXZMjnPNE22UQMg4ZUyHfFQpgddW1
KeI211DA+5HAXbnQQ02PGCQei+sfG6gRTi7xfBDq4xc5i611/2ajwHW2LoMddfOO
PhiMzAhvelmBZcr5Vg2NMzzxRv1fuU0l4j4d9hiyM17WxlgORrdoaMbngkWknxP2
bHzsdpuK4Gr1mTuwyt+A69e3tQgjFIJXnEScveITNftI5YN0Hv/8DxThY9Ao95kv
f7TQ7vlO1YqmcV/QL/ozT9C26jnQcz7BETTX1eSmk/mLp1tH+nz+dzTiD392hmBw
CSGwy0xZQRGAkpLmg5sSvPKWb+y5WZ8STOPY/DAKzSCn4A0tYvskMGAswoE965EV
f4oiikGhLHQDhc7QoTrdzQL4SWPoFgJ2oHSfouO44xYKuA77CFbEleOWaZpvxft7
MP2anR+4srWZrl8W1FT3uUUS5EL89U4LCtUnUgVpzbbRcBHr/FFlBZPtwpQf/8Ze
FQSPjhoq+AJGi3828LyqdBe7aMSYRCAILML15eD4GEXaq8w1rwkAHxHfIBckd3vO
1tHZEKeFu0Z+ClqZOZtaAj0fBDopuTQibxkLiSIISOu8VincmdSAg5C3EyTK8P3S
8GOOOqFiSAIXcps/VP3cQauprEy/HRBFYpaajZAEaGZ7klSCu4yzi3kuEQ5xs5lk
QoJs2hqA97OkJy7jT63JpcqVTh4j7a7wDTjxs8cjY7Dci7G8hEE75ww4y3c73F1f
+GoMvazKbqhff7FFldPwkjoCdzYIYq7WlU7piaPYFGYrfvsq33D55r4bM47Dqakn
dDWEIuLtDY9fqvtg0swD98ySCk5au/Bu+HDyqLFIdqJqrWkaFz8Aly6t6H+di2wg
gTkWdBvFZCXj/Mg8AgYoyg8Pi/ctp2eolWBBIeEfuEwWxIKesftCd3t8SW9DiCmD
xxiegVNL/w90I+RoSKfDnPTac0dNe5ubn//u4FvpsugH/rEQ7cRUG7eUQn7WkwZN
tRS8nD1WcgR7cr5u8vDV/4auVaywv+Ctkvi83ZihrGWi1EhSImyvDieQZ05bz8mM
GjlJ/OF9M6fLAV4DDf+vwh+ZGh2YN6O2Ux+hEdszp4YUjwiDIyk+Qj4kviOoWqWO
f6ghS0LfwM4Zu/HSyrozfZQrS7HL9EWloV64cPFhVc1dUyBhTvWxvdNjTajldZ4L
l1piHupuIh6JsjtTTqxkvdj6N1zTridIvhnssHW08ckNFoIpeDkeLO5c32TTXmZG
jJmgaMaTIMI5aTQlNsBWstDq+QiaqUTAgiBbi96dceCR0H3a/ipU/fYOo1grzLSg
g6lsL2X3donMENxRufPUdczuRgKt+1E5ZXCVmvmVGcs+M9aKtt/1ohLzm+FCm/nZ
s6TTVun1NGxfMc9cmPPKslGC60W9CJYqaMBSc0VS4BGjGPlDestPdK5+QJYh0lO3
HajiHi3hSDO8X/qPDrAzD/PGc+nM3wBqoCKi8umuRsZnApGTsiEN5fOscuEIKkOG
w/kX1t3KmEcgDaSU2M9imjl57JaBr03S9ZPXJ2mz8Of88dMHfmLNKjxm8WmeCH+j
u2JfN5KN2drGX//2WOrsyaeRBX41cqrzREQv+Csuq/eJCzubO2ufbzYyPKTjgSUG
a4t5gV6D/ZoaqIGi0q9x73cb8PkYszf0h+5CfvO1JGKrS4W8tRJKGzTUJd3GBx2k
2sRQ8cBmjqj1zBshiqTtgsXnmm1AwgT9lKWXA90kEIwOUu0SNlUVczIICX/hkIHi
mgYMSTJuJJPxl2dB1QvMgPyBtU3iG9Yympg4hMb9QraZUrBYLs6C+aBr0BUXIW59
ImefM+IgD3b15KC4lyiYIVg09oYA6F5KDHbcr2/W4i0ssyoEByYmhlq7rZ8blG3e
jESOTfREGujEq6QIbVIsb1kVb4PlQVmVFPjYEUe1i864VlnVzpRXdClZxSTyRmir
K+MhYpVMCfE8CYC1o39RZ0v52Sr5+M8pQ/1Y2Za1vMfE2u0b4WqWiE5Z+dQrfuYL
Ov4ZalFFQg1Zjc1AZGJSV0bHjD1Y2V8SONMQZFcfUiBRQgVpWIusAM3bI17ERbVT
tN20g0sSKuIaWzn3PQzd/YBe0YGWGc1m9NOHQKuFg1oaPFe3HJg4nGlLdKawW2XL
qizkA30/MkwxOZuRKYUpSral5F7FXwfmLlfdB8sPg61KtD3/MJW1uMikuWYSPQqp
/ivwS/l99cg2bfJ8wnXu6AjAn7AyuJZ+mFJbc1nvC9WfCyyksa+WztD5K3iOyrg6
IMp5oG2JDD4QFE3aT9AUP11fuO2pC3K5mCHoCS68hCELQ8UirZ3AWrzvbtAwdcYn
QdSyistjhgSOmbT4As4m6hr5ukg6eu3x5EvjbAyg/S5JIVKrJ21dFIzUpK+XnwJr
PJivQ/tJvT/DBCizyTMFdNLteF0E41mmLOn92ING/H1pvxEozDZ2XIlT26ZAfQig
Dw4XLQwYkq+zwjD1JpzYrcDQhfkrU977y7S6OwMnhJ1AatUjzRJFrWkzorECTCXh
XCIkJDXitOQtZ9FKQuS22gCmHNqiDR0UcZzRmn0gD7hbdovYp/SPJh3WL9qjA2Pc
gcqrxH4IoYVunZCPKu+XxZAuVdRmTAVA8YQZOL5Xpo7T2RyDS6jWjtTiD53+Jrdj
Pxos3RkpfWXKK+Y/kNHpMNifesnEYipefipLvfCnISjlByitufqhWFf8AgGMQm3m
VNQd+LBr8a+cFZtHz9I/u9VSF9p822szeAmfkP0XOJ96OdO3uBO+/8pRU64beUs+
o5nAv6xs30DZdTnM6Tba1UyPcLYdUj8kzkI1ISF4e0NieTV4qvytayWNTfAT9vsk
J8s060F9LN2iRnWuGNe6RQ4t7MPqNLBY/Euyx9PoMHyg2cBbDHVhPpu9UyJjTXov
zqKScohZPOyLKnp+fHaFTluUgR/Pfm4aSZ3ARCBuKPbu4JrPxQL7eT+f5i/KeON8
EYqStdq02h03vEofhDtzyrXX1sn7kyQuFkj1Hfa+TQzbNLdVRPkCaZ1zmiS0Xif+
eAxeD2QvN9Er8HBWnD+vD4FBPcWDdkHgP8EPsXuesTRF++AxlxeVdE4wmFPa43+k
H85ugIv/TYCqXA/i6vse3iqiClvSPpVa8hHWQRJ7vWq3bsxqKG6Vak+lrNzyJmwb
laq5RxeEVf225BpZEpBSiNYRDaxHxybrK6yjkiuhSr6hq1I4mFu33fH5yvp5kmVZ
rjTXUhTZ9D2fLIiu0d4/QxiDxO//5JnkwH3ukIv9X58O7WZ9Jfk5PkyqOqc8oKam
AZJ7GUa9RAwZGskcQ1ER43ogNU9d9ArAIDwNWYOKEHu2ipIoyG/xKMcsNUCqjP3y
uXZPdNe6YUvUdaE+RUA32F4w3xrThjVHp52zToyKprbwRRtWPwIkIxuweWQphixc
yHuocQln6Tbj6S3IZ21Cj0r34DKPCuF41ns0CNEMWsHnIcd4+qm6PU1tkuskCs3T
AejwW+evhHRRRbXqjGExaTcY7B8tnW7BjK8lcb3YPf3Ar3IyO8EmwYw3CBKwNEjG
BRGF7qjCiJCDBOdAwLJclbDkRzK5zKif6B0J8vdItGhFykiTDZRh+vC79VmZaYNg
Sgyh6J4MUF+PHFD1zeZjWBosDlgqTrwAKuWO1GceftnuptavjTte33DcvBgq3dEs
thRUJ7h2rVRKEIBko3rS5hZvxMEND0FMHA7y0wV0KGVeS5wuGjNfNNkhlvoFFqWE
PyW1WZR+JNzMiJCSs309R+MsoTkQzEVlTyvB3BzqqGDp6xb1+W6Mq4a0XDMzSj2i
+yLccnxpX7tawebLmZpvvjrkdVdOirirIoK1ofz14jjjmIe+uYALfgN8XlT4Cgwq
85TaxLe+vWnDCbGaP4ZEoS2qFetadc0U+N/IauG7/M5WfyuEPh5pCZ92t8Rw3+QC
s/WxYbiSU7eHRP1wTZ5vwfEr3bopNwG0HAckQQ+K8CGLgJZCMaqBIVvtv65XsiQ9
vS4d2/Z8p6nAEjWImZfeOkdTpz23/QH6rR/tAixHeDJdavCjLrkt0ZyrcXBXccea
6i0gqIywT4kJ5i6g38+bKiS99EKyhFm6rGSwfFBLJEICH7cZlO8q1Wz1rom4Ho0S
6GJfsfDpNPy7N4vR3D0A8KUIXexH3rhyeTfpThLhzJgrcch/CpF99co50tRajR/E
/FVL+Qd0XcIF7sW6PuW/cz2wIte8zo7JxOAlmb/jcdIXM+JPXy52Pw88iXcI70xp
Jp4Uo73FiPlg0glRVcRYH9SwItNcAmiQ66+R+quTsFtOWRDm4A2Idb+skL6/fRwA
0BM2sYVP/hTM0M8El/OkL8rON+4GjJtXhACYQfrMLvXLrVc1DzMLNo9MVpSjdkS4
LNbSf/3TjWfEdfc3N+AITCR4UzqCQ9nINf3al8NknvfEk9uxlmGVJ3OHWWPByHTj
WYl1dlBFm74LnF6L27lvxute/VgyfTTADABEnuL+D3EH4FaF8j7j2tPaHZjhByLu
rSv8TLni4pCwb+FkAGLloqf6vDNTXrnAP0scu+PDxkjp7dRaLF9NT6Tq9OlSB8JE
ITbH10rXJ/j3z7G68Sl02lRCN1BtAK/y6O07jmKnmdiHmNSiISCxFR/FKRiAg2sI
/V1KG3A0TjxehuRyNvkTb81wqHsKdVGuns373MuB9vjlygzIUYz6Bn6WZWt7MM23
gPkAnAc4KdAPp+3SyWoxYfouk3cNQr/vx9uhrj8LYiaI4oq2KWNL0eT1zBjKGNuz
fGKcCeOn6riG4aYaNsmmkBaHzJesiCSiAuXbRmlmFX1okPRPoQVQw0zxTLrhZNGc
i7s6GNN35xxwicyrMyMEb0+WZJvXzhYeoP8QAQkliSbnmaQlmQYNo2f5yBT61M5O
yJTfrdpKbCQXp7WOiTdUTqYIt0myMzMZKu1izh4OHgItf3ynBKL2dkuUWcG+dOWo
zrPz0DFDrk3uU1pDcZ9apzeAPqYwvRnLptR6Pmbuv7UNMZW0zdLMPY7nQkRI82ud
lQaVgDp29EywN82cFIhMuEE9ckEH5KnKtrarj0Bvl8jIx8ULEvGs3Bp/23Zk/aq4
iupFFlnX9Pl3T0eA01YwXXrpRxgA3thgWRx83P8MTOqDebs7YljZua6WKs4bL9hC
SpxoQDIG09VnRIcRkwobQZYicoEtYne+J2YpNgcX5q2qNDmEOPpULdiTM1aJKZSw
YxMAJplyJk6SeT2BMztZ3+xSUzFekrrdMysOmX9C820RdV3ue3SQ5d5diq5hbCz7
RhFw25ngN+ZTnwVRoZHxVooJtRyqT3oMbILw6wr8xfJS84k4axdK0tXw5kRotrP7
LrvkLPNBNmYsx7KHmNBedJt/MpkjbuSVOvG8y3IWuHOiSpfu+irgG1wM9/7ubvyW
94cZPNVGyhGvWvc1Bzy6KovnIp8e60PGz3B20ofHH7Y0QzH1sbSoiwxRnouBIr0D
Fz2I7sGW7TC0q/twBJhwMqFB5hzIQudwHCCxVFqMYy/3DhIB577uIna2OKIWxWpU
6BVkRTxhaIC1l1dzR+UGDmbcwiEgMf+dJHsgHp/RcccLyK6VH507Vzax4nSqqIGU
RB8SsVJyseglTJEBB94RYk2ZEXPRQnpmYutW99sdPPBNgrhd17RPPWX4vY9HPOJt
Xm50jrpu1iY9uC5LmHBqErz5pv8gMf4CIJ6XgN+G3B/0nIjvNsPkSjkdCypl2vR/
mkNY9YbjGEK79Xau6gkkRcsPUIpUrlyJ10dUoFQKfh3PLn/vIaxnqsGGolJUiWXO
2pMQa0O87Mi1dfSXrLHPRXrpKeNY7iJ+OEQRTqje7idkUSIxIrtUxcNp+iYSWGer
4jFQlkXQGmAUsh3bfkWiwYffJhzzQeoeSI538WRYzRzld8vOx0ElGIFhOFc1+cQ3
DDYGsZB+xxHxOl507DZpjmckbfFh/IAoMOddjT/hEHvGY6F6Kf3hpfJlELMG2EJw
MGGk/Wyn9v9OABpEB8kcaXuQwRlzQPXEQDBiKZDW2luhBKBoyLaClKB+VOvmZPsa
JH5LrwyIBj9ZqHbWzNrBwq7YghWO6EoW8Dw5aWLWpaOr9FXUhVrqu7dW4sgpky4t
HvGn+rnBwaeA2tERDEq6wbqvOtgkdqmddVofY6qp7ZTA6Zm5d6YBgSNOn5X5kion
qv7BjkKpzp3CLLYTlcU98dQgtPPzVJw2lg9/fO1dnd750mf36yAwqQ4TKBhUOWvk
hUDGQxfrJuIMuadgrqJu/REB/2iHGupl9dkfnotlXOeZfVZteC4X+cnKHO9cRCYZ
sX00ZsMokjNmkoPpp8CTO465mIr9fM682vNWgoMDMetQVCrh/ifhmdQBiJOkG0T0
Kpd/neEPdUHAQPrp3fKPiDrzY/RXzNRNaxF7a+Qg+KEwt3Vp3mdvoF+ezkYA5ySa
nUOfuKD/VYGaoSG0JdRxtqlGPP8gK1vY3HSm3xMpVLEkU9C0EQHf4VNzbEHMUVVP
1FIwIWppib9ZDe8mm2BKYchKQYioSAhHpA4TIte8BYtxi7yMzuhamwwls85isLPt
EZbV3oHD64RrXV2NoJ/1+Ofiv1d9QHNQDo4fTXrJsEV8235D6ky1uCGXoi6P9iCL
DGW4nQmyr0era3WMg3eguFM9WPU++K+W+Ml9IBZ+8p79NmVk+RoUcOOdc6u07kgA
nIhceQlfY3ocj41sU2YY6vaDiTAQCDOg2NTSdnPqFMU7B62i5AWbU3smldt4cDnk
yacccF35WJoN//T4XUuug9YnqjUo7NzmPCtNY3MlS1Ti0E5iLb2tuC6iXxk0JrJ5
YlmSIzyyRINsnDcnuQ18CZm9Oqg+aaIB1JbYuGd1zHPuZd4EvrciWrCGw4hchPHh
sjpq9+BV7C8iBnCEVTo7x0Y43aGkzvHeaVlnVWowWBOrh6UWJ2vmFqLWMCDKxJ7u
IDw2NcQWf3b56PjaXdTY+c8GAJ48aVN4A2NBvCE1PvqHy9JrWDntx8/0O182epBG
N6UBUmLDr+IIvQfPtGKdysf9QisGUYa6SSbk/bMOkowxOgf1dM2PqcSQYGZYDJx5
POXuaWG28KwNvOA0Po6/j9h21dT4i3xlwINxFxyfF8hRRL/y52+CY862G2I4Sixv
oyRv73T9beQTILOZ6Z+LYQfFxoHBUumPXz8Q41VmMVlHkeKuKqKlEgJ6GJIbHiX0
i0lkGSTEqKW1SxLGHT4odvfRmjOQoyMxhUVtBWRkI8PQF7vyb5rqLHSOO9iudMya
V4buv04W6TcRBVIslgur7q8gwBQcNoQCuj1QpWAexrcBRTEjVy6+i911ezieSWx8
Qy4FDmaQqEMne+ZWirxmxZWGMQrt27nnCKD5679mhydA+CvlV5bBG8EpussdFbHv
opY/mvTetGqdypOW/rCSLKPp42/9vrRCikCD32ztXH7Wgca0grgYVL1RXuOqZvKh
GlogT6Ac9eZqG9LfJ3sNRJeyf4x4+hTEphuMKwP6SMT2d+GeMylKKW6XfpTz+8tf
YJ3FazKKIRoRnbHFHqGSxhz14QND9K3jyda/0Yog0VPYFiIHtXC/fedWp5xWwdoV
vl43w6C2I1x7rUh5Jaobi5YNTJk/CDnys7TvKRFUyykjmO+Bi0+eYub/EqpziYOa
KHd9iZ8xT8q7PzaJkP2rhy2XnappiIryJ3UT9irxXIDmFvfFyFOMiDv0topiUHLg
YjOEF3uMirQyTDZo9t3RteFVGA5Lb7z5BwmJ0OxMO8c128dlX480RxZQvvTtCen9
pwaRL0yqbof/ssaGInsRWAtou7F0erqja352uTOzof0nBPytO8UYQbWtZAWnVWPz
ZTtBwvFsVICD06vhiHgm1Kr6qjsXk3PLkjFNwTuZIdvI8evkwawu+U9t05jEKB5c
8f2DUmlDFAuzqwpVnMkbxkgC16p+gALZQkDknpwjzigIERY/VoRfr7Joo2rjyaIv
K0vTYPCnHQx7UlVmLRCA9t3pf5/L4JD7xVt4ODnVITSdqx3Eq3P2ZsUB8Oij0c3f
+0L0ZfbGf2uYTA6U+gNsz9sg+beMblEfGuWBcKgjx4Rjc7wKE97IHW4iz16UKemj
Dlby3scmeaq7yJxLXJOOOLPQQUoqv446yY7VSPyqwEJn/l4II336tTTUU15NT/MC
WfkgXfAm6oqhpCcVyExJTB87xkqVNGQE9gyY9kuo+zdb6IJZkQJfDzK72oUtpftj
Pq0GXVbKm3OgPCFK6k40MTZdc3b7fQL1XTpqRsyFnpy+6JChvgYInyhyq29DPDNg
zwRxKpVHBGGNTbXs/Ws2tzpxm9kHbDA27wDSFEvdIULS8a/T+msaEnBeBYRAXVMK
/Wb1yXEgFu183OdYeQdC3AChlKdt9W7yOharQvQhDX1JysdJu3+3RTLLOccXC6rb
4sL1s6WpaV3qaIZoR50NBEFIRfkj+hEHplypNdf9FttaCzCyK4JIG10W+W2SSCvb
4sOKYZ7TG6Gu413c4yU32Pl/V+p2TPvmWyFK0u0T+ZXhEW2kfSz0emWnKVwfhfq3
jLDCilU59moe4MlO8eFm2+cS+kjLc82dmIwoqbA6PvkQLb9TyNZQPLfdu+wfIaP7
vOIahXeghIbRAy0mtoOd4i3/NBhXNC3qQgFzFlTO64NfPeISqEOdXly0U0rPQmxy
vg3W55ZeCsvD4qlqkq1NZ7LC6nkmv/CtlOHQst3H3FIrFozIoAFmzcWmNVhB4/G9
3BG2kxp34e9cKzE1287EzFyzwSodAgKnLbccyRAMy897gC6ll9XmithG1Fj4KRad
v37opNBgHlB7U+yoFbl+yto4Ss+1KQM/eRg7W33coOWpxBm4vPXDv7VQLfuc6uT/
BNVMoDk0STayOMMjauGY+7sHMdR9RP/nTi4rraxbWSHP039vb2TCAyalbdQSuDu3
3SIyAauWNEwEqsnK3v6sMBsRnJ1Me4XodgHaAM+E3aGJXI34i1sbQGDQN9l9yY/5
5xU7FwIfAFxwYmxL6+q0QVxa08ZS+sHCzZd50xnEpJJgIKudMpVcFWbYwAJsOQ2Z
8pv6j6qL9r3R4ETtcG1v+zfQO5bgqpsF4VuL1ftQRwH+C2WAC/Yk/lISfUwooSlj
pF9BUqlAhZ6zh/HDcthZBuKd9geESMuvHJ9eMHSp9+aPI76WfBdj5SMyLakjbpXg
PRt/uziF0HPuIQOwDyHNs9XbYve1w8INzWID45M/peqEYgf1Pyb8hg7c6TdJdIRm
ktz4eYruCqRxCjRtiawj0AfWEUxWmZ8S8PzmMNxJzxafVYzp4GzIdKUnPbnVxx+A
30vncTWGKgnSTc6q1+MuZiIFEHXJDdD34IoBJPkMpoe7jYh6WHA2Q7XovhsvGiva
hrGYgwCyLzzzYXF0yN9SfTGnVXOLA/Pu3T2JfG4HX5YMuVgbh+++LopEyOxKHbsM
bH/we5UDOw4+v39mC9EbbHFvMS/1iEPad6XP4Zy5iQNyzNc9CLubVOjQS8CiFKuq
+P7OtzImimEqJqvHGLr+6T9uhhK6PF5lznmT1IVVwqmIT3dD+142CP5FxxLi5iy2
Ql0bNeS3x6lYwQW8kp5TM6RwBf7QV0Dzw7mf5mYkBRGTRT5y0Pmdu3uzt4uXERLK
6PKAPoYv2XbaH4mTNhREcAtm8RjSDMnbj3EFBOPvid67Ved4LDVHUs6Tz5QQj5+d
VWxpfN7aZ49SFLQwJ2sMWXTbhr4Qj90x7Nr8j0MKAv5ouSCBvHC1HxMEmY0WVu3C
CQkWxOg24I/wO5AqRfA4dBUpjVsd+lZExy7ol45dDr5P9CtqKgPR52qeMtQeI/sy
M5JfAkFXNlmWEKCcCoiPuiTTpUO0uv2rOo7C6UQygsb/ns83A6ficJnCHIsho+VN
GGzVAYiOHEznxMNOH5W/188sPo5kSNV5z/X6yXb5njGzADCmTW97CWc6SuLTGJi4
7jTzcOh1JtUMoxUBl32ecZ+HewXSNky7NyltVAc8a1oGL8A7vpNz9ig7h5ZXrgz5
WrzdtfSJ2WbGQlFQ/Q0YflgjTAYUmO1upT5Tgm/TeWDaLN+OKN3Qr6I64d42HFgR
5cP8he03a/EMdBSULYhYp28y4jd3Zu9e00qnmvYDNdsEv4KE6b7qRQXhm6orbX2b
lBXrlCuNDQLJA4eQs5x33WwDkRuiZoBevjDX+p9AAoPUbdDIjhKKS7JftaBSHSQU
gzH4GCRRIOt3cKLo/7O4qRa8JEFj1mU9ausKgDonfH1PbnT75VVNbg3Zlf9wgQhw
FgIeGPumPYU7NRYy72+TISb1KtvpdzGKm0FU15ue/X8tn+2H/g0pu8cW0qkg9ryS
s2KyOLS+Jy8eNBrfgRgbpmfUpG5n7A5WS30D2DhuP5m+dH35s8ErAqG+9AKlkdKg
T4EyAosm/zZbAhJNFk5K8K+l/N+LLS4J4zeLpkdgN+NhZ8fMik2/9AL8EgFCNqV3
j8mt83coaVvl6j8neBJnt1lkJUi/bDRt+wTzb6hi56Hpumz4NfUkIbM22ooOO8Mh
yg4/CA/pceenvhhyI/iQMHJ43aE6lnnrIw7rnLrdhXwPKJcfC957SvBJh18H4Q1v
p/oNkXHLyk/I3h1zFZ15uJ3lTrP2OjZlOO6wlVFsF1P2ab0SCyOdegamn9+h8EU6
QCzs6XuBW/d0K64a4XbYLaH1vMivmIkSDd8j/ska7CfBPO/tKeYfwKnmnp+JEBBE
UJ7LoTFCZz1FTJvkMnTV7KrHiAD8614bdyD7Rf+umZzxtWFZUlsgqZPQszlxUAqx
MxB6PK22WwOUxRePCF6BpfA/VbZ9K0Jjzs8zjZBZ+eyrS27DDMLMzlR+cdVi1cdu
Qx7Z8ZZr5/YKJ9btC4TYYqBkmQcLuORRCQPv2YTvj7CCu0PxXmGlj0yauL2IDQKa
9SI00Zh3H47JN2gCA5tUsUvEGl+MGjA3jzA3D8e5zktwEtad8X+AiTeGhxcWpXEc
d9S2uvzchvGiA0V25TKIU5i5AhX+3CIb7wmzBnpGqeL7hgJSYp/H48W0b9kqZNti
gqrjRbbe5gxu9ZnWwqC8D5l57X+fIEa6onQTDcTQj4bVktodckXEFXlBq/nKs2yd
VefxIhNNEGRQPs8k4jBm73eDnbaOY6pHUQzvmvwdjoMI6226r1yyUrOPU6GVw0d1
idYaWuuFs2/ouJmjrF01OcIcoiSShTaBCD9Zvb6EGqhZFPq1XHfLv4UJVTNMPODt
vneGvUlWa24HCXMCxeEkVL22bJ3o7h6Bm8tZ4Bybjjl42JhuMxwIwN3wfIS1SSem
mm3MSQ8O/Oq6EbyzPm9ZU6e3J1vhHtIangf6b8flgZNeLoDPNN25BQJKvOQM/9yZ
AWjDMeV7lzB5xv76eY0RmwG+QcwF89Akkr+g+KPTgER6zzouDQCOvmpKuztkgBds
vVwkhNiOrSrRQFqphsgZQ8y5XxOQV/ePv1LPYymDNuTuflQIv5dL3PYyfHj5ZzpL
CZGEpnZVmfI+J5k8SMYar7S9wUWcXb0/tQ7sBID2n8MK163AlX3YenQiL5eKqjRG
5vVTsrg0Su1fTKOdXJ+k08+XZ1i3oxpa4kIJFKfrJZVG8MFUNsnEMXyTFpYWoBXp
NKAW2pCdjXMNvGX50H79JUdz1Fv+mwP9tYIoEb/UeD+ZvtJp7y0T6MAgzG7O9R9l
dVCCPqumzXqMhIy8EbOiuIaYbonRxiHqn6HLWuDj3Jfoz0OqAgb8h/TqggKiCFkv
4LXzbuxC/560lmeZGtrU7lsTKTl6IFZEJSovRNgT5t2o4nMrZer6m4Pb8U6bIZZG
tfeCybbzLAhHVZldnsY0r/aqii1k081vOzlmwxQTwGIekHk7//XMVwHF9FVA9jh+
OXdUHTJ8yxeXte8URAlKOaauuDXzlPU8QF3pANelqb//WFdaSEmHElTNd7Q3TZoP
oUCGuTf0P8ffoHKCci1zRimvrb7DujNiLZCj5dMAY6nnwAu95vMF1NwPSdXBc1f7
scd4p5gnsemC1us1Skbxe85nvGYZtz7Sq5RCeZDfpaRms3LkHGgszoMVULi3FA2s
Kas27BWHFgsD02MzSik6+gwvmWcxOVzinYN0GvxKzOLbiA6YMxS0b+gnUZi1JXDx
Sc52iw3ChopfWrUOue33K+q5P+DttQ/MiN9nhQKFCqdBM2tFNAVDOx7xIRlXXO07
3JL4s2XSSMnZ3OQnEPi/419ty6o7QWrRrEhT0tml4Z8Y0E2cDCc+Fa208QC2HMJ6
T+ENQh6Zk2hTMgcSd18cvZdlmqiUGpvYFyB0lZR7Ygt2RgqKDqIF0Dv0+GDBCtaH
KJLTLQBwwgjtLahs2k9S//ocFTxQB+cGn4yW7xxTZNCOb3dCA9Xh6E+ip9TrHAm6
TeRrhddRgUopWdU2GgMxvJr2r2mwXlsa8RTGULxlmwhSL4/O9l17vVUKPSIrSCHm
tyWDEZCtdZeaWx9UzfDS7ZJLrRSKq4eB9W7MDitYoHBjVRRSZ2E4sWGSYqc0R6Dd
GeGbCyqY1TZaqvXuoSpg1ixSBV/n9Hf0LYER2tX+RqvMgBuEuzdI5f8yPvxDajMl
By71lrxkPp4PAiRNp6T0e7GJPLlSkKqSbF2wx7CT/Hx6tx4IMbFNVu+HgO5AyCBB
gfNhtxe9tu8jPbIBbqw6Oz8t+R/CpuL9d45o8FAsFIQVrzsOoRooVk60DnNzaxZV
EGlNhQuEBRjCEHlVurszkGQgCNSU2M074Lgvz8TS5/VVYNH6fMvuGyNlR9L1Iuze
eBsgqTwwA4t+hRHaGjAYCEsPabL+YJX9kZMNdExqRaOL3zdBFjjm0iwis6MV22ks
DCU7WJszLgbU+eCsrJEcKne55Op3DCW2PR4qq65QVBnq0khQVxYfjiEjOnEd7rln
eYEb9dlyQxjBIXMB9396Hq35VOUnDNU6Qen+NBQpUIHrrlaqWc3ChPiHq//GS4Tg
9MrS9Jl2rkmBHyQip1cdRQijKE3GA9EV22XonXmBo3/dnrdmel1gQzC5T+k77VBs
J0nxzuw4ohtjjP6At46yvMQek+ip7TrEu7FV1O9mOcC2FrCadCmOy9ePjoJ3Ubh3
RVcTjv73l0pKd/3f7bpBENZB0PsSWd07ClgCIzR85pa8GABcOwFHl4y0I/l0EFFq
soVH7AmYFh6L7ilDcOjMdsiTfgktzOTt3w3EI8a/5Eh+LqXOJR5+z09z14G+CPAV
zvkgP616xV0NVEtiXlXAsdBT7D1NyZFWdf+38yLNllWFLoRh3RTD8mvJgN1kqUkO
BxDmsQSpsIjQQA0A9T3UewUKCXvajr1b5r9zMySkbGYmS4tei3NZyD7TEE21xRWi
jad0zGccHe1LXt8+7xYCN0CGwSaV7T9omcw8DVYHLnCFtd+JAsNHFc3n3g5nNBFr
k8a4oPiYJYQJ9kRYdDSae+XePmK1wC+6VAx9mVSZ8+mgnDdb3N40ySqerKwLAWXW
cr9uRdPEfOAKrVoMXXFsxUxYQr3wNiS5RJabtBctX4QTa4C4pl/TDKInevJ4R0fs
yocD3tsiWurM/dp+uo//I63Pu9ektzAefTQf5N/EvY+yGo92/7+KHbmcaRc9q52n
/4ip0ojVA09Ns1ot6vmt5xz2c3U3QqXz8VCQ02mH+F8AdRPcVXSvYMIX9erMmE/m
9vMmJ/yVFbmABVzcY3958XNI7I101tHuHmUSrnpXN3OaAx2wc5Fyok6Y1cLxNsmX
FOpIbyHVjhYub4uhSSG+XNQnXI54EVOhi90mqXBEdaq377os1FCSDTyLO28scrDP
DtsE8hERNfWspihUZSuG4Zti+qzcU6N9urUWIivJmtbAB0UoRgM+4cbd2u52E/Ff
lIOMJU5l+c/zP5xv7xqWHnGg3kxb76S/Zure8m1CImVcPlVQlHU+MmxmtncBnxe3
lc+2pwKDktuIlaUYuMxEfL7kVyQUwFhtyxn6qHveccaJC/99MG+JSJ2qE79iBNRT
n0XXnGo2H5MWX6lkNnMWq2XikVUopoRAIxvlQvtjq3gixtiQPHzRGrvFmo0wBVU4
cFiNZdKuOq/a1QDqOAZmrjWcQ7EcR27g7vPNB0/JH6TDgSWeUdDuxV3Guh/+LWHH
UVf/0eXyKESOSnt8N1fROQLyCZvC21Bf9dmDlabSCcPjPlGwKVBb9guHiygczlkb
qBvMB0NCRv8dwogAyrkKarNUFb67qlLc76qWlaqyxulAa1ZfbUWp0lgaR3G2i25r
cKMWw6Qlfe53E/2vJAoc7tdAO7A3i9YtUKVyvTmSx0ZSw60WCWrJ3DAv7Qp1Lr5g
zYKz0tOePLGaZrLDkt7uwcbaPbEirRU+3Af+gXDASSKNQ3xSMVNjGrFVDelhr96x
4CVUwRE0ynlnGHmhWDhQ/YgHGqpTELEk/rAbGuHxUgWWKKoVpbbTd92vDe2ZNGBS
GcLUppW2Y0DihHHCGKJlWkm2Hf98c+WHWT7FexECThPHD/aSex6ya89rcS5YN5h3
1fDIjsIPAZZC+zX0JyxIV6dBsj8WtecZeSAqa2iUWQSoXhUlp1a5E0zvsqRv38Xq
WjulhikpJoD0WA5m+yPYItirpwVwfKEC/dkMXy8BhOsR2UTGdVTHSBWrYC1oL4/4
y/vfsAMqW3GtGJzjxsXhvyJxcuu5ftXIZ0wF1DgZRN3W7d+mL4PnN3a5QW8z4col
LDyt/EGWT7Jbcrp2FZY7aptwubdpWnKo9d3ZnGFxmnsq28TxnhubZQy3deAW3E5O
Kcv7UinfhXKATz54tfWpnEhcidtwkbdRpSmxDkvnhZ39xs5QWbSAAYVLyKqWB7fR
Azz32BdZVfWo8KOfRXZNYSeWEadwMFkZSjlWt1whq7t/fYjovnx2UaF5fAF1M90f
6cwF4B3iJgRWzPSO6IFJnLJMq0526hYPJMIxc1q5HqtBLHNw5LRdeDryc2h7Eeqi
OKuE31BvhyEviuqb4d5KJsnhq1Uho0dpKx6HSOifWgeCT9iL519H8v09Ofikm/eu
+yH2GSKmsQa+ieu+UlNEMzBUw06NBsSABid+efvfe6ahHK9tgcmkzB00VjKsCVMO
Ct4tnQSk5j6b0OzDr51G6G4M9CswCv7/xUUNmdANns1l82YXJcn1WstZ1m+ebE69
STRcb1IYDbKOClWSEW/OZnw8ZC5AiiBusMzCfSga6FE796Kf17uk2em464XsnOPi
Yath3AG+G0dwEPVWflQojWDP6wGFr63XyU8v2TqKKuIsKQW5DwQROjz41pm1sQOd
gwj1y1KtNWyOPgLjqnmD3XQ6URPFHVwQMUs1yABiRbHkDle8ses86v7+bn9/Ez94
/HXKf5YLLWwE0oLeEhfTgpyIlD5/EdDeAwjfsbEounHP/+bvV0iv6jFn2vFfREo5
WPZgIOqm5SspwTELSZsgfnC2DcJzFe4+QwE1AKsei88H3c4GWEY2NvfIoGW7ooMb
ZH3pax7y9dp1EU0jpJfSFfwBaffsQGnh6Tu+zSE4N52MU10MB7tw1d6BjNmYd+vt
1QJ8eevpO7XJ+b7ts/Zx60Kz7/7w+SduRr6MgwGB1aQgchVXiw2pko3WZA3OZ9Ld
In1Ot6NigCJB9sYDCDiVpf3Kl5WQPW87eJRstcecynVVAmy0lt4RIg30w1rtjWMx
jYtWvFzbg9cTqDBIdAt44CwSFcLPg2uBzI9vK5phjjYpHrLdQZjk8Fn4aKhrQc2z
bxFm1dqeCCZSNwvM5M9r+ty83WYvG4UIuBdb0D+cZ9izDY+IeEsnYGqEaMWH8vb0
FfjFmYLjtqJeZTAmnIE1noPUZGN8XQM+eSwXefIgWLymm6reWUrsXt8xliXa5vHJ
CxWZ/9MFJjiKZDyNSiEDrXsRbO3jeYuOUP2nlrDpQ/ZCQrLMsVtv46Y5ZWhkn8hZ
Jj9ggD+3Xpa3xTW15wIX5aefnP/0ENOvuOaY0rYXUCgcr63GUmb4qEVX4sogSxQt
T9NF9Zaj1bI9+SyZqSvz0CHmhXSuR7N6sPrwV11rSiExKsGLO43TvdUxBvxWNm2e
yOUW5T/58I0SYimPvv1iCXHAY7t1LrzR08kWXyKXWepRHimmBXCFL3pYd/ZxYqET
ilGBEN/1j600i1PkFQEfluiIs1peFCSIXvZgND44yYTVKi60bJDniUNq4bxV1K+q
GWvSnvDOXnzd00SeTAaKZr8BtchQ3dr9N2UV/14hKh++314P21D8sCh6MuCGZENU
IpzHGHAjiXOd+IMrf4tQU4DM6Y3twmTbEI9xYP42n8QX+bKad0ebBB02/e6WB6Uq
a2/LkTPLXXvDsGVvzZGr2YWAcLRX4bx0J/R93mtbqrscSl0Lt57cRWp+pgBeGJ6N
wCr/Kqysj6rQRHqEx62M6bxWK1jTrfaoimWjB46CRCT8DfqYIM44saIzsuESWxTC
76IzeU6TQQKOCf+AfYiIKRfLGN51w4AftvNmUM1fm/EVIAoOvh2Ol8/w5TPe8Gt5
HGg7IMVcyE4H8uq0vLbQI3b/kSBFIe4fpP4KSuPa3rm+12MrpJimgLABV74vf+8D
r5hbl2HJDcB05XI3EIwlTvcx9mkT36pWboGsJpuVr1K/+Lh9NS9OdjneInq3pY7u
d7mRL13okZxBhWic8ALU1Jf+OYEdygDiykeEpEjKV2QEQrTyXsccCGx5aJHflX2E
O7zKqeQ6JlxAq5mWFIyX0Qg+zcoqM5N4EkheLFnN0k2qZS+SldYDhyEy6fQiliP8
AbyUpZFZZ0DfuJTbQEM0rIT5t+o2C5Enr8uO95wXn80jbPIkYg3Y6hSAEhoXFmuF
RB4Jdn5/+cGZxkhVVGPxScigIfs3On2QJwSIbyaMCQBcvYdUPP+tXH/iZVbMR7Ks
+vW+rSalWT8iVbMnQeMxdiqsvQ6jQeZCvA9Nk+L+cBw6I9WKKSbxJDmaDZpXQmx3
3f79WyMiecHHp4Cp/J6X3ssjtCeJnfBc1vdCrtdUJKoV2yW+H5sCHob3wW4OYrQS
JJPgqBgG0AbChTLRd7LGUdTUQu2ufixBITbGlYPEnoDGx94fidWKmRxL2kz3Fdcn
Jj6KVEBEjreYVZ6q0qIrMUapXy9MKX02ryTmRHcUDqHqR23P6luounaJqR44jpW+
NeFWFxNpqknLtYY9jlbXy/elOuk1UvRLc9QL/vviWCfMu27431uELmQuvHfloySh
i52+SaLyDT1MmldufEBI9RHxNAHg1Ipfik6iic/JnCECcHiLqKpH+bNj2GZQ11id
iacK/M2IjVJihn6ijPpCRV01KzB7sEcFXjxwy4xoxQWEoNKsFejLSHwrxtYoGqnl
Aq+6o1zcDiOP3e2ccNktDZgkSNsDbet47S49RKY7mxOPQYT35PeYrvjclMnyTg+i
hgSEpXfycaU6tWm3Xn1bVeFtXOjNrbsRsiMXxp2BKeDty8qdAOXL6J0s2i49YpTQ
YeVyvOc3pJw4SnUxC9dn4c8UDizttjfq6q2vjVwNSDFgVbCgw/VLIP5drcfuphyB
R6HgzzOTjjje5QdpxJwRxwJPyxDAVQelueKoX4AvoxCvqHzq8ON4dlS3ieKK+Cwv
SMNh2RGqIeaajQQML/s+RHOoo2mM0zmH225yMM40zVrFVcyBQvKRmbTJ/fdOZJ5J
IlXWxOVK466obKgRRNk1GKTocdZRPTtWzRYzmJrzEfKj8a/H/BxPwoLSqslUx1MZ
EaMOD64kgzeZJzbd0Rc8ll/IoGdYCbyXAE58qMbWI+8aRn/jToADqFd/9gpCoiXR
PRKJjuUM/vGOm0VvX3jn3DJaubu8W4WBvFv86OIhCgFOUsSDmv/F4z/w0vUHC8eO
ryoi9BOvF2k9z/Jfk76sOd3tDLx1pqrFWk3RE67ko23HEYKfl/l10V4Tv4fw1/4j
bdCWapc1lIoGN9XB4r0LCUnP94BYMeuiCXHWIvlTpniaQO+7QVuBlnzKIFg3t9l1
99ixLhRYGWo39ez30mVjddlYO3rBngPLIh3WfSBr8tJpXQX6jEuHR5DC4QvFhFv+
7gbPmQxsooIy4HcLDHjCq3bhNcjeYHlCYyp0bz2tKfnRgSwdKuJJCg85m6obcoxa
KnJGdn30nOB+P76YTESVWTmDSxoRjSvjQPk+t8PCOvPyBWB3JOm8MHT6ml++iXCp
fLRTe9FniSCwEVXH4rMNpKZa6PsxcZijMH+WrUpwJNJnCjx4UZ+3+qGCrqplGDrs
a4cPVSP2nLPBhVccB7UHmW2aDLlJJjVA5vHwzEC9P+8Dd26ode+18R4Nuv49HGLd
3ytLsg0L+ftclj8spbbi6lfS/6s7rb/41K9epBISspx7k/pgYBYJLlp5PtBw3fKn
clTbI1F75CE6bmCRmEFNq8xM0/m1H+z5nKg3nQqseiN0R0fb/N+XgD83pquG50kM
riyx+EYQeQig+FgbSNE6SS7cAnwZy4d7VKxKMi5zidV1IJt+FefHJwITm4oh7YQz
CTANNFX1mBqrn66ZUfZWyIdt5qJSXiHUiz2vgn8cebj/bbjlFoPJ+5yaHBah+G9V
lUnRCHcTAnafAeJvv6IUwrzMOGAvRfi//xbQ/hCBXIA1uNW+5XuuvB5x8mkcjyMJ
F0oQKjCTlDDa8taJlmKTUPC4ehM2rywXnarsa/FP0qBd3a+eo+6plLfR1Ce7eOu8
mSOAt45F8I6j8FZT4Jnzzy5WreIeNxInQxr980V7iZ2D+xoF3gwKhfLDRU2PbLpZ
odf5PaL5Yc+EeGgRqLgBBx6cVKDNBjnSfawVeUyyP9DcsEqFrExmYvz+o73X0RKo
jDWb2TCOkVStxd4hlDdzAQSjvuV4B8QxAb9cE74ta0eE6t1jl+EEXjn9jlao1Mwi
NDloAnPmYpipzUch3mbArA73YXFcHN6jKOXjRkCRniXZ2nd4UNw6qcbCDZkUGRTk
lSL/ayM15ZNMoZ7ZXvEns4xAw/xgd6NiVfKxSrIWW04vzfGs539U6kWGMDqYoB10
rA00ohUySRw3cTynXbRkWhwNMywY7Mvaiqd191AtIYSzDvptbVk0kP46P4LsGs2v
E8E4koWwHtTfHClsnWkFQrVeHw4G/d98zK3GPMOpj6KIJcu9XqvPP1ys16o75iMx
YnGEhunfWoYD76pDuvUDkCcLxY9DAfortMxjMcl7L2i1sw2Tgp1pi6eRpZxsAZ1V
wntlStIq1aojcrj6zKeK8PAHZsgzs0BOsB2gxJvG3Q0dj1D3YZi9hp+MES/Bo5xY
kkB674UWsjEmOQ09whvBlntxlsNVXJ0DHGboGXn4hZUi9MpBPu6ryWz8wSG97+Zm
DNyyUJxUj8NXxl7oEPIOWLAHJ9wEq9GRX7ZszaAgTZuJCdSo+OhtaB1IGemVEfbm
vyFAH5WSo/t4KnZmc8JjFcpnEoM0p67h/KsavsWekoQgAEEJwF4FrE7M0YHPYfoc
EtMHXe0JFHc5j8TrmBERmBDjJvo/TlrI65nzMBlDoQBYqUGr3GhwFfpPkN6DsuDL
GD77ItKklb5Rjf4RzHk5OSOrm8bg58au2XTrVJu+3eo9UwayKS3APIUTFLf7oOG/
t5SG9mUrXMWpm5+8dDw8TQ/ahyJc/kSfGmNhCzj9miZb5R2bUjLIaooaWDBJOOCv
Ff9CoH17/oCAoZ2lpdXMTQC4Yu2UIjYyueau2C6D1VlftWzxboPrO5gUQ0tsVEJ/
5aIlmCue+JIOjt4vc/kv6F0NKd9rF6M3ZVVYrYGcOR2GjlnJ9xaTtnPLMJAzkYl0
cdpZ4BUwcRy9vZnKxmHIcCpMeAtqPY53keKUnhOogyEQ2JDaGWi1uYbWOcfAoTIW
xwdOWMkQZRb9ErHGW+p8nPn67Fnd3Xbs1wtYrp+/n1w8/Yri+sv8eaqfHNM1pSYs
UO/jwiRk5lsyfafM3rRAXzGbLKROUk998FkCGPNzEXMb9o6SLgyr6XkT8isliASw
NKjyjXLzAC/V4I/Bvm17M8e2VymDKHtj4anovjHjSoFVn2IlDRdulWgFeT9Q3sIy
QSxjEsh9mw41DtfQ34M7hwEAHROufEpnOx2ETXG/oTgkmYGiE28DdzToEjOm9BX7
skWb9Xo3VUCJFsnwGmdd4YfD8ZgS49bVyhb/eil7izo2gGkQG7Zm2KlnEySAJiFQ
RtZDJZxiK2HhRyCM0xy3/YfUtw1KAQ1aWGvsJ2p2Lmks0kYl+g0GEgGBbRlgr2r5
TlVB9OENcpBwFeoefraUYerpTtYQ8p0x+Hxkyn7rQ+sYp502jJbGIEOeyYStG0Ps
2kGZ/O8dT4qjhw0j9EV2/xpoIODYsrcTbEF1Y2KuF4WPuqv7rt/6Q0bDtDAGs5gp
WDN5106dv1Hc5rwKZsfnM4etazXUz1T2p86WDIjqK9O9Kyen+EaqbXPPLbO/EBu5
4lNAa3BLqAGVGzqBnnLOM+XWzWxukRjrpPIF295YOIR65Gb28s8MUqw6pBBo/3NK
AigHxIrCm3t2jydIxkwK1wSuk/RcGJ4vfBBZZqUBFe8PrE5hqxiqpsExkwMIuJ73
zqJ+E0R/+oOCrUB9Tq5k+Hdp0xXBwqjbvbTiR4R/DPsAiozKqi5D9pah1fjvJRw7
+qR+u0D+6MmIk8V7sSdK5PgoVrzv/3nHngCsVU8uALBvFugiALHRg1SHXyLFr0Tp
oUFwEZGvT1SpjoFUquavEScpyBC3eVsVIWUuKTN5bfj28CiFvduiEFR1sdHHs3Pu
bdz8H7WBnhdeoTDq7RfBEXiEXjlHq7JySMQB/54E5sba46fRhk2gsF61ZZbwSm6B
EMHiuo+K+0dHflpBHl2gS2edTdkaonxHUOCY/HKCCkWJv+qmOsaO4c6UKEWgumEi
8Bjs8DubmBmM9VxbJBlDgYnhJ6FHZP3M2KrL3GA/e1CioCnSKo0HiFDBKbYsDtyH
SQI//p5US1oQRqAwwbPCGonTBZAfxJ2yJE5nPDrmN4k7llFP1MQB/XU+RYbLhnoW
uA1+FMs+jOw4yj1HTvzMh1K83FOOvHG39pe8tqbMsIamWyMuHAAWTJDzbJE5+9i8
glN5kkoiYKq0pDNQ9Dklmw3WgZVYoeXpE++nmssX5ZuSKWRvtW+dkFNTjzkAgDVn
+gR/mDh5omaUDMOSR8cs5FAQnFdZIOc8UBFU9u3AF4HkIADl4cJtrRcByPddXaYj
4Tw5WYVUELKxgzD0ZzyKtJNvX8fyI6d2Ke2IYak+UiO/Hsr+dC+A+Rbn8cuiM/Y6
F2Y/bRu12F072thuPwFShF4y95wCCUjUCklCHn0V39ixX16UtN98mz7JvlSfniTL
Ps1bB5nYI4S+3bTET9uB8AEXjpsBbNfSHTzG1eN5OopWWnSCiqFMkVKJzW49/q97
BaM0eV5rWnY2Wnod6n8SXnaHlEiHRVSTY0M7y/IFq7T/pG6TLuvWxXP608gHOhsf
pXI4mLbwbxlc5VIIl75ZrrzV9ba0CMlmMzczd4bnQ1qQ1MST0+n/UAW5cA4DijTW
EwiLu7QVCQrgm1vE5eRu4qqEJnv62Gsl3FiKwxwn4PM32EAhqatJF3Vxcs6duvSU
2LvXhpamfPhekIRCABYi7Jk+K05JLHK28Pogav8Bfu1oSOubKHeo7aIARm2Y1UsK
Pf2v8z3Viwyl1ds7zt0ivbnudCGYpfRntPquXXEGUIDzdg91GHQLzojKwshwYo2f
FZfYmCFgs8SHV6ZDoPJyhstLB/FyN4335PYZQe7XsJDAPd7PtNkM0GjWt4pz7oqw
R3pdPEP3eTkeNSSQbD6KBA/oSaUT6ERBDLPcpTnUQQJGT0yMEq3wuSfE1aeGY+j0
p68/u7tRmk/CH6M+qMLExZKb2IY0o5lPNUT6HwesOgrYUSvpScHuZ9WzA8op2MS+
SSM8hTm4I6dsX0qsb55qKuqEZOl1duy4g1vDrss0EaH+QQ5+YW2SlNO29jnUExmH
o9QBL/1Lxgc3qN6kEZTrlsR9HmcWKpaxsw+nY5UrVU+O2HI3yLz6fqq7BipNMAoB
RRIDULj/cpOq6xahjwAIFwpoVUC9JF+j3+n3Fs4jAWOIEPIv6GiIwDsmzPomCcap
psshsf7m0Z6iXjxaMEO/HH0cJJBn4sqN8NJ33vdyD9BdJDi73fldINmSJRBPzwUB
0/0sefxYHc873RCd/bd06smXmUVUeSwjYrdPd1cyXViRbcvWtkTjgMyUVlArp7aV
d3bQ+kiM8f/bAXjcyW3tCjN5dZYJG2Oxbfi+rE7RmbkJ0y9OaOGE+T1d8Q7zieSo
OM1OfqLuAs8bnw8YcsdEfR8JDZL+6h11W8gPVDclZqyhYeGe3qxTpS290c9PJbBh
EBlCX8sy0koqsg+Mui1MnBlYZ1H4Uf/C0F8E5W+0Fqh2kYv320jpHIlisvq7AI1n
ANed8pCQBhwF64yIA8XC1uccGBkYQN2HEbTLkceamxrgAiik/RuB2h8OQ3dnSs9Q
hHgbt4HFK6ex3TaWk4g9bxek72w6hJUp8mCI57Ro1EeLeImqEe/XCRJfncS5prSL
yQSQp/808TS8PPNxYCToFs3+IahpUp4Ya+Vfh3V3bugE8/UQTQFydjRdlY5y/e2A
TYyajmmkZAHp7ue8XAPUIt7CY2b6KWP49y8to0MylH06c7kOBUPCDPW6rGunlOti
IZOxNGD3G8rEDE5siAWEEeGVW5m45N7rc+F4khhQQVxdqVXXxb/P8nRr2gEamUdG
ibTe2JHo2TsjnQQeLPhDRh8CVDeBPnea+TtGGVVaZi6HzLtghZrNsiixojt75Ds2
GS0bFTXpHdtOpurodauhuRDcP8EwBmEVtgB6vOnrNW6Vw9fvjDaY48cQ2WbBWgkA
QqgvkTU253Weq5G9MwZCY8L6U2OfPVSCCpwgD63PrrTJR27NPYbR7OVRGQYWkFge
rdBAaUugXKYwo6pH4zGHT71Q2a0GyyXo+poDUExu+aCTSe2BkPK9gz4Pm1qORl05
UcT1tRXWVWAuR2X145Nrr4RNTinK7JZ+UtdOmk6MrpUCmSWfNucI4jG0gB8+qn0b
LUNGZfM6hOgjKoBK2NHGjaTXWGFCrOCdAONXrut1RKkn1sLx4t077CoGvCxq7663
25ccwyJAA1qEAZ8rdwQWko2ZLQgdAgkkQ/HTNApPGEEUY7u3GPUwTPSuZbUO7WlB
Ll5Zl1OHpzSpR8sfLeGPxSJSd91QrFE3FOKQGFyKzmJKa+7JeULBV3rKp1XuBnRN
rqSyAMEZ0n7ZaFj1HtRwJhzr1G1ee8uHfPPTeNa2Ubq3MjPUQTXL18QkiZv4Vgp9
YDA1AP2LpARHGH6WrLCzUOJmpnFEJzDClDF9+s6LgS6mTyMuxnOELVapHK/DAUd3
NbvT4ZqwDlsdI7UCKEJqC2UKCQDLLiSLya5AVNjnHhpViDeFrij0nZTZSsXXIwc/
FK+c3BcBi/uQf4WZ/Xo9gLcRFpdA4ighFj7pY7rxmqth9BhPdCJQ8phh4OTPOrFe
//NZBanTc63FG9vQ9AOq7b8KnqSpBvyE0tWURT9SFGqJ58uAjzSBXZdiEaAOTKjH
wXW6SUdLy805IFE/r0NpSvxaqq3JpS1k5fQjFINDZMTdsLE+jAZtblmTKZFIxW61
rOLhagCGyGrZOmJk0MNhSjGRX2l16F0B5CeOID/o49nL0wJMeMeUEpmMp0k/lt+A
kmmhjn3RXdfMAWko94WHUT46iPRQrfytye3ED/JSmrsvKl5JogeEXiqUBTRVyJkE
fZDyTpm/rbCnEBP7/YZ2JqciZgesKYCbhMYtyvyNUUSaQd26dTgPxwI3OZJkSbId
OVkXR1DjzbxjndjjLR8NB/5zTcfHnh8vaPlFHJ8z/lDz3yPGV/uyTNZNidXnjum9
dwTAZbINGE2Uzfw9QpHj4+6F4xPlebbx6f+ImHLK7TT9KGzGqRy8skmDcK9aAtlC
7i7mQOqMRE6LvqNKuCHd0kA88ANNZkt2Pa8DltdDRtAJa8aqFFdjXzB6GfYWvla3
T6qLfo3leGAICM7Y0fkzzhNbjQQGntE99YWnwvU8ubILmILu2Ac7K31Jfxdp3XkO
umlJNdrdTEuP1XcK+gGUH8Qfd+WyxvP9xoLPN8P/aSxa9gMGrkzQrJtHYvUBoHqM
rx5WTwoBWNAKmUa4qTmDCJ4uk+2FS2CQTXTR3ydJizkfcOnDkANZNTnVznXjPoVR
c8wiBhv+NtkwQ5iB/Jyo6WgoZanE7e2HeTdBgoaMgWbsMmWArqVQvKBBnpqVdeH5
3S2cBCgtzMkz/lZzXSqCiMHNKAxZU2i3vQQT7VNhnRj/kD6Usfup1Vox0RCWaADa
Dpy6/9/bDhLwQ3YHxwcCcQ4NVWbKZQHu3caa55rrAazFFhhVWYroPV3hXHN8IgKq
bLBwfGiEL0r93XEGiAW0f1y4yGpXiDzsOR0jxBmYU9lCNI+gqy27O3eZhMnAtI2s
p98F/rFlafybOzTZUo3R4HFGQFnHz2zkMdY7cHSzVy35kptQuV62ecfHPY3mw1OH
21BClBPnLAFn/aYZay8beWVxE37Z/zVCwUHKOsLrBQ61tfkA5rYv0cdYbn2z6e9V
mfpnAVsZ/lY3/Uv+5Ql22Ek3orCm0oRezySu4xTpo+jUMuwdZ7l71CYm/Z9xQf59
GccB+A53hU+khL9Ybf0P2hMYqMxBiwUE5vp1HkR5BI7mEP9CEJ3/Z9/1I5GkBbxu
T7KwM6PIDnnMJJFGGbgkg7JwrCuQY0j9B8ySAL07tioXSBdjovS9VytNIHaYh7s6
qmSzFXHwi/9f4dV0vrxq/TOz6/hcSkb9b+EnrTyn+TiWM6ba4TZTXFSQd7u4q6VD
oSDrqo5s8jKVrYtVbzKRUhLx7SGhfj4ByZZiACSMrUIHkZblhJCE/B22U3/sjlhT
45Rn7lXOJ7zKcV+d8+rjsIMh+YLzc0BNiYPPY8mRgXfu0c1yOpn9HoeTsqqLKkaT
T81uyFjSxj3CasR7wkZwU4EPF5N8zh4uCoyfzlWw5yW/sRdh+uRBPu60P45G/MDB
uOFGuqGC1rXSCdVGp39I5+3WWMkE3EiTXNlCPNpoYthJL58j65jm2eyz9XsQkAB9
EGFvJiacgm4UyibuJwMvHInrHXl2+nhDKBBse3QVLCg9qoGuTtmV/hJC55fJMwCM
ZecLglxvHyBs8LTDGeM0fNER27D3aZKWMIjMhMTFe9VPUh0ZcBK+mRC7onshMwAq
quxm2wn9EsO46noK4XKCoV6MEOGFn6jNR1JLKFlaOQ99Y3BaG55mMabYFCyMfxNP
BWY8Y2s3kqW8E9SmQu6b00VUZazQCCarQMePHyhE/cOgk1Y4MxCyDdoxzUmB0LGT
ZKkU76OQRPo2dvAccL82YUSnWX8VM2xWFFVosdy1zHw5FMZC5JsUpRnW7invp/2I
u+hv3F8aKbp4dZb1OvD9vxdf2zbfBQLOw5ZFQO1mpwY0EAyTWS+QZfi4orf6AJUI
6gxY675sOwUvU4Pgli8BkKUK1FTpfL1bOl6BcKIJdRSEKl1EsZiPjta3b4/HkAMH
GFHKLVmgEa6mJFX22s0dKtGME7xFpc6ino7m2HM6F0wGIzHovGHXseWev4hjjPfB
c2DL+mJ47PW/r/RPdbi8JuuPPyhVs+NfW5Zuypu/IdPF2mzRoxuT5G0cyWuJM3c5
uRo3lCK62ZBvlBqP1lJAV1Ht2ejQ7tm0Ogo9XDTG0eCTHfbNgMTcj6L+M/PJfxbp
sFZ2Wp1Ck6/bGn/bv/nzvkeJrqn5e0BaHzIY9DVMAUdr8HDu0RQH9kY1EEA4Kx12
cydbU4KZbFWJwo/I/XoSiBqmdPdhaBZCc8JBVU61KbSGGHZTQpEMmb5/DjfR3vG6
sQHcS4aqUaW9JVBPlB9LDGjxn78wnU8U2W9X34Tlh06HopSDyO6yAE5gkxMbjZpU
kSi/DOVkxPhN8o5GoHg1TCCt7BC5krcwvC4HSEZtTtJ5lqUzShaGk7FQ2yMSzVsU
2h3pUmaNb83gdGaj1Hcbwk2XYjUxWuwBwj2tz6ZDTe2dpTPfKhS/nzgtuo8nSKtO
kjyYK8etFJyIcrNsj5QLSVaItpoRjSunBgeyit1cdzx7d6XxSx+0yYxoP5f4X53A
WYIcgKIir4jDs5zjfjnqqGzTjkHkqulXXOXqq3P0j1OKZhlU1PNzKGFSJVMOc9sO
ImOZqxGm3vfJtVIBKTc7Pq8XeaWXzwbd6LaeVFgWSvnn6LaKOKTOaKtBtwRrgyd/
m5KOZhtmipy/uzibkodtQLI98BgjFVTjLPTKTe+E64YfixJxNkWb5hBkyhTJStiE
RxixMj8X4i1K2YgGnMHw4WpU85vlynGF7Og6huemP/kO7XXxpk/rI5lVQ3UD7o1Q
VKbtakTj3vdiJAjF8ZQ5gIAAclImddvbZkddkrU3mXb1EGaZsmJvl97vYkADeIoT
RLkKUptTvlmvXqPS24FdvLbX7pr0PzD6O2VTMbZvg++0xQZvRXLJ2kx/2OLNuu1C
S6fdkXXw/egphGhE+UiFiQOZLUgyyxqH9QSDBYnxLg9pd0Yzkh1Uft3VqOOLuYWs
+bT0KwOLFLLuq+jWWzV7/hJLildvwnfYZnf4zeHo9QqVHyZWvkqK9xaPKn0L8oZj
cJ5ZJIuVx9TOfkQ2yY6949wP3JIDgB+kyJTRqpJV0ITWLqm1sA+JlAtHcyu4GB0Y
ng+y+1ASExA1UEUlZHkNDLkDmwa6EBP7zKUjoN3ZghB7u7ssmzYCYMBU9IKOSJmY
p1tboumVRQx3O14KqrxJ/hxeInT4mBi4YBudCP8wmvQMFKZXwwlAb2NokI13dqcF
9RUe5zPBQQbh+yLu+POoLsMnWAzeD4bP0ZRzTGX69o/XXV5o1s8gqo+69JEOY6Ca
06T9NHqqq36U62OdXm2mED9G0T4pyFsiRncFuBvwh+hAhKDA0fo24sI9ulYz5Ux+
2Uu3UKHWiluhtwG9n/4/rqmFWD9j2jJMZ13MZoJXxqTUVxS7w5Kgt0RtrnOzAcuY
SE8ld3JlvshTKme/kDE/wZ40z9gGn3wSBsO8mXEw11zIy0yojeUPCVPUhZe1RIvb
T1XzbXhXf/QO1a619s/D/AoK3wtuHsnskBdA/BAR0jhUVWrbnz+kjHRGYIkqH2x7
n7ze/8uoXb58GyEhfg006LL/zcSd6/hdSDrLzoc7MN3qX5WjHddmbzCqq6oskUZu
EmUQyHcZY4VCtX8QQodU3EJnmCdgiOmSXDwy/K9czY+809MMaJr3J1ueAgYpYd05
fL+przgsvQbEZsEynFkrAw==
`protect end_protected