`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10368 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
Ju3IpcJpVj/VshHyynUPTG7kN5gTlvLnmXIUJKrchuK1OxzQ4c0/CUTLSKUrnTxt
0LhiTpma2HaYPPVNOkjQMTMj242ulu3p/xKN8H7YUDr+9lA6ZMKLuujzF8b6y5So
cTn09VI3m/piOWs9O+vVuKJt1OI14cJD8WqdsJ2XaUThLdD5JKYy7N4GKWNbUNj4
YYErfiLQt0LWRAdtHXpCft0AgEPhW8MV8P9gCNLbmRRLvtBF0vC3Q6tNfFtMjTEP
+vyyoiIXvEJlCfV3MGHScG1tx621l+ECYCg8qXRG6eDMkugEdEcatqwUlf8EvDsQ
HAWmpneUWiRFZ5wf5ZKDTu0rG1IswE88rVN68MGvDIN0ZYrOcoP8gEC2Yt2iQu5d
FIjOBmxugzprAJpNz/0GAADZWakuVtSLbpKEVXH2R9R6xmnOSZ56KKbJ1Mzbcm5A
fZdWWM1pEAp3jKyr1UZN4r37VE5yMIEm1MpoK2JToqvp+HN5yG03vLHuLgRwK1ab
9QEQIVhTw7qFSVM46RIRCBrdUBEtbhRlS0W97a3z8LYDyzfRCEu54KlIDtbyGKPi
vdcMmbsp3O9nVaw2B03axV7vdXJNfMR5WHl//cuwIBMFl/ctZ6FzAWnrWvIDKbPm
AQttH5jFljfWY0lBn+R3ay5dOBQabjvtdrKPr37exWNw+0Xz8TIxRB9FZLTTHya1
EYAfLk1pGy1vIHtQKSl5YGA6oi4iDWfVtQ2rKCyAoOhlwBoU2VxYCL6/T7ZmuN+d
R7yIb9tHmKhPXkDibvtQXivI3maiA0qO1I0fPFbcBDKOM8o0VB/sOzA6NzCZNCbY
zhP+kDDLm3Wk0i00go1AL8ZVHCjDTM8Il7mU8z3ZH0dsuyXMYKzjJio6w3AWO3BE
mBebdNa4v/xvVWzu89zs5lBAZ3SCOkBqtloXeYqmIR7LVBzn9LScl+sru/xBJq2S
KQ3lVk5VPwgZbJhi3WklpQao3unNiO32wownI+uBxA8vdNdcD7B0bOAmmGYqIOdv
kSRlPs0mAmDRWYEGP4OG8czT337PW4+iVO8mknnd8y9HYuXODCDwEuFVM+LAo2VH
CmmrRuY1GlgITggeuo2VaFH7TbZZsVacqfX6yiNUZ9oI609YAAgBMM0hZx3fjYQB
boRVnBPMdosnDqK89l84+xUE5idpJtf/v8J+jEoZxJOroFg9PiB0DeogckBIjlFD
NALiNebYIukeWwd2CoNzTCA8HD+2ymLpd4GVrTJfZqipzyC1PPDOUf/glS+/WO6r
KDLQ9bb9vUQ0kWsqBC1wTRTraLnreqznVaIW7QJ9m/DSiI+bO7gGY1YUO2oTc5gy
TL+84zvyRdoZqzN4MpjlYJgMp16RxAuQKoqhsgxXTMKXpe1lnCAwbhZCYtzigm0G
C9lrroNWQGnsW7B7D+v2E6XZtv6yMRj3bimzHdQYslYpeUb97Pe+XUdsF97iA4bq
xo94DFbF1+whThrChgbv3ol0wY4piKjJ03zMNWfgOAYxSGz5Bs/FKs8bv2IxQtbK
lS/YYrHpJUftAXmFp20ncGB/8Ee3Dtg0YxeQ61yDYR6a9ObQOh74S40FTAvynTmh
UosBozEvkSFcrUwvIB5Zhsd8wYMm3QzAjTP7GezSqwOhbmUwXjWgwAGlc8FS/Bzo
t0fMZCVuC8XpAQ/Wao7Y3GFwcoqlFn6fHfHPSwVzcijC0JUOEm1DY2TctyOxGWQx
xaFF/2m8axgSBIY54qv02QNXcp1z2AN78WM0LZVLw8RwUUHQEVJ389iUJ0OziyVt
+uK2g1Fhv860QWkUyB2VjyXUYvWRuZINN9o+9DobOvVwNgLMksbN/n6imwbc+O5U
O9NtZ77Uvq6KdcxSsVGEMRR7RdYS+GjRC9ccSHv7UFAFM/xaCmHybj0yX7OdaJ4t
7ved2InF8RRXyAJqYFLVpmpwiAAOcz1dx/SV8IsgrI6k0NlGlQ9sRyZgw9TkI0oB
WASScLBv4Dna02eAHY4ZGGkYUCzQSx8Tv+x8meqA83JPoYd7TJpY3ogG67oOXzOF
nArnyMfjHhu6s+T/yOhgf7erRKNqssLEcZCergPuz0JJBa7nG/GnDR4+nxLxkrrC
swsw1UjAhNU6ePnSJMhJnhDatZWnq6EUV+B4FiPa/oB8vdTFhBiHeI7kXlNUMuh0
r+D3FuVXrjDL7cV86XJxGaMNR/+WTHDt4ut+rDA+yfgRYskr6AvCCBRLQJ8lIQg+
MDRk5uZsqMbCj1kGZVwqAvkxHjbXx9UK0HPkaU+4Oy9dubxKXU/DTqzCD5b5xnLj
5xuZ/QNVL+DtlcRMvXclCVALhLwuPr08cNfiWSEE5CM8P4rmoM+WkluxvKh+6GcQ
ZMIt6HAVJXDEAqjD4j4lwqVU4QgAbnO8ui18JcBO9kAPvDI7mISWC6Vmst6GluNk
jtnx7MtD4erQakHKtTv6QJaXBCV9pmzB+r4jJZ+53jrMw7xf0wJqMfre2Vd0Ychq
6rVlqR0AHmDcKoWhZPvi85GCLqLCpvXzLyGWT4hJ8BJY1U0aNSjj07f0NIv2GuS1
BmxGEU4jOYtflHYK5u93EEirqpq0CdlTi6duPrw9iQWOkHaW+bOQbdyhXSgxtNBZ
Rz2FyKA8kcWuhaSRsGNzZRIkXOBYxPwOV5v09+3UingayOYbXZgenmZOYCx9cauR
kcIH6fb8+5vfBnkZ8ekiO35sOYWIz/Fr/TYEDT+6B8zbtnEBDdFkuKqsvYVUV7Zk
ez89MStxRe+VIvk1Nw+Hvx4fSAYP8f0zNWepulVPuNHLDoKWSmbCes9GqshDeFW+
a8le4ERDBL8KdX94fiPdljRjlkYQf6Z001l41h73NJ35lyRap+qkznH1nHJDzN2d
8eNX3BrCsH63muU3fGffCmawHa/OC+1iPoi0OKwy3hAU+h9VnzpQMCQNl3PBEeVh
kk+/oJrrFwKQYJnPUIaPxqZ2nGnd9P44oB1vem7HwO8MDJ1YUkCBVxXUxMH6fuRd
7WrkHtsSzHWZbaSyUl+3KWdK+6EjLmrdJtnZFXdPgxOXwzTS45/jZaxADWV3+2Qk
bf9JI5YFCqCzCxFZ/WnYArG6/+mjQ7Y+uj/C8OsO7ezyzsqKauiCARuSYsyUz5wY
sCyvn9wQMWa+lPBrJvIYjMfMTRtjC+bd2MhQCLUUzfj8rFpcHLs8ABlJCOtWvuTA
jQ6KeQ/Xp+rqs1dxZIAjhpGoybXNvq/AyXfYxDDa9qBO8hADWgBDSgHp38Nw7iK5
zPAg6UJpguB6/Pi5qEUS7MCttc5UVilq8YT9KmxLzkVpiRrNtzNyrsNn4ZHBtw5r
2pfzcSVByi337jzJiOMS0fRAK3xUj66Kmyky8Yap8aJ8JCP0u2f1a0/Xa3iE0Dzl
YtvtwP4h3ip5GEfIy7yBfwroEMbUbDQY1uXv20ecUGb+YxL4rA+aqh4dMEcmBSVR
XLkuWZtRjQgPn5fdV7LS+kEEySgTk+2NKw6ZBhKoDX8+VCsz4t6xd7uvUV5Pf7QY
N+/rlahtYJOXZfLmjhf85wnEXdtPrwAM39MghxTmFcIcrHnHHawl46UpBIo6yYID
BXtH4eTEB6PSGZEvhcsJr1Uj+NyvBNLx4sZi0Xh03YuajJBWOJLvMqSemtgZwQMG
egBHZzPJUIaFavdE/N5JhnBcTOL5dYEffdKbP3FVVI3WgRXwhCl+taqLjPd9IFNI
2gBLmyKwUna6oQ+NZ8X3LkwBMPWxJvDZX86XUyFnWtbDAsYx0IcagDsNVdVNYNoh
X/TKCtmnLo7BWGJVBRd5J6IljHvmRz3uwZxdboJAXdxZYpLztMPm3AkqbDdYfgsp
dA4jWJvwVy/+BqrVoYdZxoARrUQDunbM6Un9TbX4J3OiyRumS4mjsZw/kyQDUE5K
MsGZPBaroer+ZJRytoTy8SiCZSAzkZCEtZjiiYNDWo40gkxFzWzQmrdxWwylkwXD
kdSgCYATryTj1NSp9e+DSdfYMLbqjqJpepvPoWR+zAUu+NA1IxAuugKaq3JNLWrB
oWa/hQmzwg4vPoWm583BhF1kK/Mnz8DqAg5YSve8riisReiUvCxpUTTMFNK0ZemZ
C73HVU0TUMgFDrqT69iMosnOqe2Z1Nxwasxnn8BZ/YWQfGkY8QxeafG8s0zreInd
+X3W/F9eMSXEI0BKKxRmaTIquUji553EZM1OdOOsIre59WGtVbHxwfijBqb54Y2q
PXBC0Vbv2rwyCpymOPHQxICKMOqWZ6Gxu3REMhTr+s8AtLj+b9orIBQqBaqGDL3B
Qjobe6tBCYqffmN5tZNFt5IA0tk/O7dLfdwh1hNAoitHKPsBsdNFQNBCJZiRn/ZV
dG/G113SIOLNNRhZ4loEcBPv1HR3QQV9LF6MLqmudw8bq6zNty1FrGFkuiJYs+dN
98or5tnriVCC1gNlSesdhvA9Y6cKVEO6nZRK+pNIbyw4EI77zRO+3dVfGqnGNWEo
LSBK0PwOxrZT+XPUOeb1zHUsshgcrmn5X9eXptCQxya8BjO6PlBfe5zpdRDolXm2
qcJxj4Hd9Q/WLFkQBJAokN798SG9Py4UUMnaRAQbTNmUgGzqpAQUMufTfSxjNcV0
Hl91nIXLjgLMpD8hlI1D4Xs30g3IE432wt06tk4Y9GQ/9JEgFSkQxw8vFyfR4C37
zKHA9msdq6g68n3lu3ycqn8NHkj/RDREBJgPVmsehyDZMb6ARcxYgv6E9MObDSTe
wrnIHHV7Pq0TG+ZAZNp6EGpVUmmmNRH+g4KfsHaNkhe/vIwh9BNV6cDbZGa7rvlt
Y3uQiqSVFCfHjCC+5tjzxRbCOovnMBeQaqq/mg9z44/Cec8EDomoKStwa4kQ9/8O
FCzx4SNFr2QHk4Riuf6WD7C8OSPfppKVKRRo0JPwYMnwJUc01nH0KQ9wcrziuVgX
yGyihXkVpSuDux04I5tyxyjSODJX/ThAhPmwu+9WBlhaTPm+1R1sq/67Mhl7tT8y
anjphKEHeUSVGVWUJ8XxXnpkLo633sCSMFV5+jW/biPExFR5mTYAbWqrUCuxutgQ
q9imQcI4fjuXy7hjEEgSDqSqUZnhUClPuFwAYKziivgrCBjZZxfQiurxSOoTO94F
VwYN8t4fS1CXQP3OhnzEKyzPh+OmthKNKImDxScgzgBGWg05PIYRyEhtkkk/DwS4
sVQVqseKhJoXEBzHK9dX4q4H8hh1x92N9RTLdhS2IbwWclzEfWlV9JEEF7jcNWOX
jIVe4UBgEO3oiEIiiNhCOvXLG04w/dY/oKqd0ZCQd7iyOguBfvFH3u+W/O0n+bxp
v+hqtpZEYAMEUjb0Lu71YWz8OzzUGkV+vkDuGqYEZvcwn3pD4fJ1+9EHJlJDzmjQ
PqrkmWltTV/SKv8is8qOjTsR3GXNCbsi0X51VWEpmZ4sXlpUspp1MtcTHrXw2Dl1
OCMfjwH5dpZzGwAc9rARQ5xQ7nCUJrSsgGy4Rs0qKhADdCNHF7DPHnWrd1qOXjEp
Iako1GgegB0tny6gTPVVqMbXl3bdfKndzpYqZU7TPmJkILLBpxvvmVLzfGy+e57V
Reu0FN74RlHu1FlVToI2F3DrZ8vY+I5S/3jZ/H37PSHYfYoaekjUwpEdYmzYRjX/
kaRg2qEo1Rthp+cEqvoGYKMn9c3qJPAlz1AYk104wKBXgyuH/MlxPRyWwbXZzrpP
nPLmDOcLbVE7JlbCd7pcy7q97sa+J3zMG5uc0aNMIk/DpaMUmS24he3aGJ9Bur2S
jCYVnDHg1KWrVeoBnNHXiBULC3zZX9hrwKhM/8uz/wIIa/NOBEftTeBeMt2Uf2Fi
pnEtNRDMV3xEpap8RFpzxutVuuYcrEk0/8XNBG1opY1eygni2KPznmmV+TlhTMYb
dAUfLYfPVHCC64swjNNzW65AasfpdeD+7mKE2Y4zJy7gJGsiZNTg9gr7T1zq8Tsg
uNn+rXN2mu0koS9eeUqMvl20QLwnDj2mjtwa4n8edbnbxZUNwAQ090g7RZ/mkbaw
D7ypuNVT+Sh9IgL+VvagYlGWv3zHvDMbdzWWd6p2mnaxqDlFNVArwApONoTg544t
IJiW2Vk1x/eP8/RHAEGlmK7MHgswKOFH/w/JYHP8INZ4BicKOVWST4aQsDVRDY2F
vRl8lTbT9MeR6pujopbuF1j886ivkSof2ukLh+A+pJJC0tg0QjS6hTKrHV3ZKvVX
4hcwefvcOyBa27pwG08FDFOS5lXpQw2j8WxDU/JcCKRpH518gDSIQeuMrfyYSSYU
tZBG3a6XOZxnpriUD0Pv45/3lWvXWV5MV0Akg+932CzQXNSUsR78Wjs3/Z5g6H50
HTgefwMC2+0xa7mYE9qliISUPm8Ve2e3LYiaBowaYrfSyxDsb8fZ7KBZxANdQ2fC
87vq8pMt4sfLyfjijDDMPcFdVxvFT31LjOj/zVLjU6hsm1XQOCp6x7CSpbcmp612
7E5Wl7IyABEfXblTwtpa8jkvceCq3N0PD8VwIosJ0Vk7NIgmnSZMx8PZ63o2exyH
/soVhTGteTnWo9MymFjpWpe8rF0gcj4noYXaVTZn3VIxsArAfodauuIeEyHydbB9
hs/H6TlZfzwRH8iL8Rcwj+2570U4NomhAU644/HJJzZVGQbM/iX4Bs1QN2ltMCaR
ELc0p5dYUTiFdzrpYf8wb/Zh7+EVWT2wqD//76fO5R/jeFfkUUV+v3kQLQS3aRNW
yoRqvk2K2P6EKPxChqGfFppy/1lv+TR51doPK6kZLK59cmb0qOcnRj5ZbRDGCxIQ
ZzLSMaBwCo1BAD80G3emdeOR300YqYeAx3Xp79ve379gQ+1dCpvaABwg9VIGL1Vz
OHGmqPWbaYnZywIQ/twmMicr/y0yTOYlugJ2iQqW57ugl21ybCf9YTIwO+ByNNeN
mbzfzAtyk9zzE/KqSnQUEzJj/awUaCIQncf1FXgZmVUsN5+wEKWZY/hMsgIFEKo7
O6FxsOrzLFACr+Mxo9caC6Quj3VXLu5z1X8k6LUBQTxWGRXGE7B1WGRJqySbwFnw
pe2+RR/zBh8hnwMXoOs29KP/is2eCM+NanCUZAv4v3/vx4oJwGVJDVg/nsaGq34I
belOPvrdak8s+64Dvd7b+ZHmSGQTrDhKmFWCNNWdU6I90jePG47ki7B7JE2WhcBn
w+RB2X7P/AzBMhn6hO9yqAH6TER80TRMLKKG2NiCLmPS44rR3IvAMUbP65iHkg/z
lBM+9RVVgvwX38WYJWpc5OY3mpYGgiwNT3qfbnb9o20l4RvFA7X6UjwSTpXD3yuC
gzX05jNFxuLnHaCL6VbouF0MYkivZWUvjdEBey25AXkV70x/WBRHhrIn1XLe2po9
Wxn4RcGfs+XQQbVE6nSc/RF62I+bhkvxyaBuBubv8PEcaasRTU1nfCDg+ab+u7Zw
B6z7fs30dApv0GyXtZ9pNQWG9iwE9SZdGaS2STO9ebDHUUuVYeKalW3JY9/o//X8
jwMtJtTwAKtCrSyoIEolh8BCV0oGkiWb/mskawHazo6+37gpWgAHOuHdSl/Mubf8
X/AuNCMrLG3IW2dabTI3xvN6FGPkmPwaFrexyL3eeDix9bc9xhbJYbiW28pjtTdV
jEMmc/L2MypI5Ga5FPFJwNhn1JlQN3VP5VBOzB9N5ylMhwQJJK3SrLLhGvKIIEcD
d+3EPpXGogJvXSj7eSa8rzizL6KZzKAUXsjAQzpg7FpnyLv2RzMkVQ2N0S7N6a6u
poyufQqK4HvlipBU4cAmoUEoIEOg/kH9J2JE4h7m0qhIjjJTHoTuekFYC9SEGpn1
V6XQsJxLKiL5ja9gNOW5VJGxkY1YMvSB1DJzG+0DZMcA7WzoLDCHpVIfhAoGTzOF
yybkUmxGylDJfioB8wsGE2mUwdlAv42LtQHxXBdB0qPAujlSmhDo+QOjSVPKAN+p
XkyS6902r4O3WvWyVaqFD7IJU4qoBs3zSLoFp+L6LtJe6ug2HP+nS6yMk00H1YT9
kFGuU0z3nDZPL1upi6hHKjq9uoMhZDaFO9A+sSEPitinTPCj65BKnRBfuO9+0me3
vFibUPlkqTFSBQ++we4zyCoex9Ox/0mNWPgUkKeoNWCtjT0VpyOvGGi2YZAV5mwo
vpPv1sA4TcN/aG4IEm661lLyg+53IBlxoU7wPvp43lyLc5EB/YUZ+IfrFNXKBOck
Pfcs1SCWJ+CLmPEJPPfGlaSuVKdWIEUqHot0ZIb9Nuih2zAt0us1hItt/uhWpFtF
0vf7GhRqGVqFbXpedo+S+Y7tiovrpw9q70XahpDEAJr/u66b8Mfi1znNquJx4Z1T
82eqGd7Fnb/MXBvJaj79STVju0n2lI6Ao/2XcCIIMM+9afRV2KMQ5VBl+qIv9lOy
+Pu2dlOhFI9iRRWQJX55XnjtcyY6h2iJZ17PVloGilyPmv8x8dNRqLMNkv4hrCCy
Q5wNiiGETlsaajnmpY1fI2wFbmh407pBRuUULolW837bdnyxsVSj96m0YHSThii2
GhdQBbMYl2Yx8DT6f+RpMeb9W41uBrCI5ZwuOwv1r3irqiKln1WhBTCmo7p21D+k
2t7fMNFfAUQi5q4q7Xv/xJ+aG9l3x0zjRH5yyUemyPDHb9otckfRKEq6esLYQ5bS
QmhDDtDrijX2B/30UALJKHanFGuSbwofbxYtAlxPDKefFap4yxoOoHE/htoHFzJF
6yd5cCaeXfyjafasYHuAtXs0BMxnxGkkKelH2dr1c4gswQRjiKMwqvWcWVksDZB5
asvYbOoLfJUAJ5zGQkj1nlvXoyTAkszZSsxL/mywFcPOkvM/Je4AM7DL188okog0
9RqF+y5W6cdw2xnxUNStigFZXlivQWyGrcjrYNgS3qMhxeWL/BPsN3eTxiYgu8If
VUoDUvvO1H5DwCWK9SVrSRSs2Fkr4oSbPw/Zicfn9QW/RtR52DASTGMH0hBpwLkc
T7ttVlQNSKt10MaLtfJrXIYuTV6MIxUXH4AOOwlNsGcdNLKmvlmw+cm6VKc/JqJj
/6E9UBDQ/XDJIyvkx5ZAZvDnq8u6R4VMdtOp5oMApwL4S/pXDSkJm6Au6vwvovsC
gc9xOkbADS5EBD1yAhlm6xc9cFWPu69dXAQxsdeyrdo88gdvTh9Z3LpzflqeIYRr
PG7ovfRZEGZdgvb/SRwNqasjubrmwAi5yS+hXFmtnKowkmRz0yK5IEYJM//vqKxS
7NOXxh5SzC+lXUk8AAhfwXbN1PyY5U5i2fawKFf70v3UwwOxPcg/HsJzg4FltQ7w
ngSBOH0kJwxSit27OfXsYYX80GplKlcib/Tv6HMjmHyUkrefhgdOOnrIKaqRotW7
FVOUBQkQBP20ZPvAtAHVEmnlqczGM09qhr35LGcBCGzElgyJz0m07UZwqj4YOqz3
jr6NFUQ169dHR80Y8iLpoi3Fwnv76JtqDF7/nbfMHqfPkFynLr8353vF5kS1ii4X
gFsBb3HZyN89y5gAQdBh2N2V3T9fXvwuqWeuBFIUA4UnHUfKkB1qNkKwQWVINeXq
iN00Ozwq4ho44+7NXqjMwP5CgVt4ICnmPbNr7AEzo5mpwf2DoZv1M16rDnf68mI8
3TbtIFLwnrhWdOhkwmM5fFZ4ri5RWAtKrjPQdBsDfcSLQFg3UBdY0DYFRqBTp4p8
vWBS5GwXWVKlpL2teQ7LMlF+g0/01xUfR4oy3+pgPUxWmfcmD+5/N33kwfhvHVck
JEIU0gGY1n+UwBnkUW/MRNLzJ4tDDcf5wIKBkiO+L3Mg2AO3NTHnrddXq119yHOv
kwgKq93reNzKm5/6kAmCOc30/3stwpXB7KVdiUYoDbKRI/2XWmZedDlbcx7uiuH0
dbmzXR43Lna43qD0sMUlQMpRtvSv66AbyXTNKmyijQQhgdKjPzebpOzVq3EwvPEh
bMM+Y5LCnRt6dhm9ypFqsdZg5eXKbdckDuygYny62omOnIrtBzhini2p0c8G44fv
45bpaMm9ZtwUpuv0WKpyz7UU+RC32v133BLXSZ82ZexFVozyb4LBKeEyAV1rxop4
nfDewdOEmr+XvJkUpUrKOVG0uL9JV+Ygt0m4BJWsVkVMrQx7ncM3BFt6eqOp2RcN
pf/Pn93sslwXereKL9rCCtiwalOzfj9kboIdT8SAr/quO9+i1p+nKkrpxCdXVD47
AK0BWVK0qVxGvtRGEw/vaHM+6GKRAAh7FDSr2KTxDdyaSmZW+05ZG5ux8vsF/xVP
utrSRQa3T8Na61atTxed//t9VuPTmxbW38DxLwXVvEqhwd3wm7xzToPK24phGLmq
95EHAbiGLVl0O3yrN94m1+Um2es/Em/ksvur3KKJfhWuYBHbRD8EU5aRajCxVt1B
/He1JILawvVPyCs4Xv/hOx22TISM6asPpOGKMsqZXc3S7cCQZUe7sei4KlUXaUtw
kV9w+B4JcnE57W0Osxg61QFoWNRI+gWK8FLm4XQkis7ECYZHnGGLKDNMUTmcoDYq
h3t0uaW8kdSWCdwmgq2xh9L/egt/RgUwnTCsJCylgC+XGjT8z+CU55B7vM42KSbi
xt9AVDrWGcfFVuZo0KsLtw/5W9gvfJ9hhlqAd41u5/Z9ZfI+9b2wIM8OHR4ssocK
2y512zVuMjnSqGdSXtye3OnNbXo7haQJro29l8k4FOCCS0Viys/vrqb68/4e//5B
GrXgEEg2YqzAdcA6uDH7B/nZ7pHuAez7vNB6UtA2OcLASSt+bvM/A4Nuk6N6iwsK
RItvUZCuKc1LA6EDUvdFC+wRmOpo+nJmDJZZtNvJQ9IhgYPlXjOSXqOJJSufwJiy
va+vKvypMrID7Msp0bZrLfxd35EGLsctjJWZ0TEq7RrDFmngp2mB5Nbt1mBbtU1M
CQ4K3E8uETYO4veJJnIZim4dH33+EmxTfSY8Ywew21v37hy61zdBsJGJsAXzOspZ
t1rYR6Slcy2kNrpUnQVYogbjdX4L6RAl3Q5Dh0c4hG66pLG8ICkOI+J69p7MRVDz
lrmYD2ufPmjfvVQ3p+BZPgkofJOADCk2gpQD2MDDwD3jDgJSLLTV5s/INPhXfuD6
xBrUQvV7EnGMa6/aIdFvpT5EZDWNgGjrVOdoyVs7VxNbz+QF9Vwz8/bNz12P19ww
8XKYD9Ftta7YWu6anjedjkftKskJwZjYCmf4KbhB1h39K3fDlWhkUADFLdcFuF/G
m8SBN02NlFGU9SWd4c5J0oibpoFdHML0p+jFM1QHX0h8qtE9H3sIWLaSx5uNEoaH
tkgFMFDRpVozXqOlGyyjGYdeC+UVuSzjbRPPh04+3cMGLL4EbWO4sgjgLRoK+31Q
WWY/gqUPpTN7ThbPqUdcRqav5lS+pFL50cQiJ6s2kwebTPPS2AUfkskT2NS4SB1S
E7E6FXwLzpJnitr38dzCvRyAQXSNpwOSK2S/qay1n81xyAa/wqKksAzqMXt6q8jf
fNhQSO7gRZq1oTIeOVtMg9Ft7UxupAnmnoErqD/Y/Iej1jegsUWg5/MbTL6aiaLl
z7thiQmlt98qAv6Axb0hH435jV0E0HQxWlJ46uChHCQNYeulZSY4lqSM/lvlQwIp
+nsPSlOT9E/2lxHEy/IiqpiL9tmCk5b6+IDzkTlrSFuqUDO2v/mVWXqI82nTYWjy
rq7ruhx/3hDmMdhGJSZu27XicpcDRj8w2DSW90sjguwYZKS7amcxgmZKIy0rdEPu
gpC6DfBjbFz6ST/OFWf56v1WArZ3I2UMMZK6FDlKj5HlPqw1HBWnzrvWd0tJQKOr
mZ73oeuxzpNhj9wDJcRilco1yFLIpknl/x11Set/XA/CZRer+LRpVWbjX7G8m4Xt
78DYM7AdQZijXH1dLS6ptkRPg6Y3qOMpk528Mf5ytFKCxhoT2LqzBfq63LlXBrH0
hd5BrLlae2n2/xgq2o3pwLuiLQX7WnsGRvS3HQNW+h+Lgq/OPtF8HwVhkVaSRnzT
yXW+tLjmErNXculYyKq2h60GV9QMIcJAJrkE4Iw1m50P7RA3YdHwkhPoZMGMIEh9
OJy+RhB5h3blNyGNKvL8yfNG0Pgwh1IVAJ04P/WhE8buLy5VwaEOFD8TtUXd+1pQ
0Ulh+o/U/sevVvhCREDvq9uwn10ZoEwjBL8zAmI1Z3aP2k2S3hXf83adJLD7lNPr
fa1ibvDRHZWKNyts4np3wXytwDfttQfwptbmkEOVHrY2aUnlqoQIEsInktI0xxxq
xrK284oUyAc6jKCk2TW+znYwVUJa2/m7Ur3+/7yfJyIN6TxlKytJqPRaDuiu2tiL
HKb8Ylo3Yj8Udj/aXvH2aRjzqx8xhdruzsNh5iuow9EnGqfLhTZ9qKv8HVyaaO2o
Mlsoc5KoGf8JVJQ1Zu4oMt7Tp3GMkW/6qe/GbAdk2R5dHZfIMb5JF6XnwF43zHEK
8bA7F1FGc6fbU9+wz/NPhDyjKvewcHABuy1R4a20npr7rWppafWTH9S1nbThLTj4
1USEH6gToK/wPNhBG/G+g0ISuV02SaIN/E5kek7mYQXQdaleY1cEQMxAkZ3ylR38
VQDbHh9H8MNGAe6b4YAMKLHZHKcAIezZ1ib9q9ViN86lXEJxEMd2tUY1qy1kvXVo
oTtf47Ja+rUuAR9ZaYN/DI5IOKa4UdZzrDWn0CIy1L9PI33ZmSXoQIIe2+50EPzo
SEkAZEW1zaz5u5s+DglZyaRrZHgoIUW79zhXfrzsru9kjXG7m+RCRTJsQEVE5q7n
hZp5Pfz7W2No6no55TJ/u1ishxFuHbEjxcHXoQ5YJRt94wxAoCSqbHvIVuegWDuy
OGh2imqsfIyqzv5IqYx2sY05dIw6F4S4snN+XyHtU5fAbntqvAOa9+IwZwlgV+Kg
VWmBI8a41OpKYV1K50Xtl88y0t7utzizdn6CVksM6Y4h2ViVlAHg50JN6YJAXDAO
fjsZCt/D072jkFhgLaWjJMCrRdHRQ9mv6uqxBoKIZqFOskgBoh7yfrrH97Gec667
qsqLu44xtWJodFn/JRhNmgF9Rb3+8aRPHhtevoaHUSGYbwubXpUFOoOAtpBVOzbE
VH16pGb4tgyQW6qI8W4oaAtymVnilfF5vvcyDsxIpyg4++ANc/DiQ7BwpFzTXtcj
X/Vav2kGCV9yNe4UKebw+D5Y4dJSs+ehUfFx6yvBEgFcf2yYM8E/3Us6AoWbly8k
LRNZnLtapNH7BU6FlX4w4CfU7b9NK8gj0BaHRr0c3xan8ZATzsil9f0JO1JboPUB
hJBX3/KwT7pFjhTuoEkXI1fgqYJvKPBaRxTcRKl4JYN+DMkMueY0s4m5odDkAYYI
ojLKA5jluYHw2yY0mFCCTfNNJno6qEqAUrO4Yh75gzCk6amZlLVxLj+JvY888E9b
/dDex8IKU1Z+1ECteowTglGnwnpRpZaxGyXzvn3l8YO+DYRhc4hwRaIeXfHZ1MF/
WcehFiyackZy4tBAXS+h6AdTgeyC8ROatZpGBuiY6OqVsUUY4fOR+lZ3Ekxe57jx
vasYKLzIm6Wj06/HV4YdmcZScN7W6AkR9jGe4330rDYvOlWxhzwU9JSrV/L4juBg
+hvB3WUdKNfw3NT5jf1t/dhzKmAsIhA7Cw2VyFFWKm/I5kz0CU6GRQm8fTrTcWKS
y1Dxq1p8D4u8ENma6QrbApMBFMV6WzNtXjyuHO/jTfVmCSJ5/eAqVdR8XZzsnNKx
`protect end_protected