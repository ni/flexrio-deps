`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5040 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
DmI0zUXpjr6rtg9EJrlnT0jTVkJqOK0vjVIVF8haM8e7zeIxOZKy3nGk1GjfMRzx
D1iXhBnZsKh75oVfDXoeE/b+ev5MAqibR65ghaABhu98NBZbkkZvIQQap80NrFFh
lRWKqFC7+a8RbfRKbJpzGSJh58Ww5q6OgGaNEw2WG2Mscf6dZWLg0R6W0L77lWBk
3Gmdbcy8QYGbxXCVOeM68C3d5u7fBHAFJHfZs29f1gVfQwpc/hs4kIrSED8w4M7g
EUNyMKCyjzcSkkEQI9+6EKwVFCkQjoqr0C9qWDrE0v3GqSL6KRynXU4QiQKR6mTm
y/EzLaj4auOx3b30I1bwwfvvv9MThZ+YfVrI5ddFmZTW42MFm8zHQoWWz5MmrRWb
wytPKwTWZcFgP8gqjrZW8tTG70mJMptnHa3X/sbWUqHuhaA3PSLYS8/PEkZjxPkS
w3cjpSpy4NMk4uBqoubZsB6D/OOx7gV6EP0pTzKzRISJT70Ngu4Upvmaia0r3Y8J
p2u9S5lPqFXLTq4Hwvag0yfJRhLjUjsWcaMiJmh5eMfscn4BYMhhZPaZx4GEedsM
8izd8ut0qO2+3E5kmQqlv5debjsfgQKDwbzTnefSlLtO9B0YdQPADny+IWWU5zRC
5l4gbhugYZv8IY1HpCHf/2tllPiy/WsmCQnnsDnStvRIwc7lkmUN1FWEs3dPG0Xj
IiDz8ZU++feepndFc1bIYl1EXXiF9Fqp4R3LhWZgk6ZvsqyQkg3Lkd66s9SjlXg0
lvUX82Ij4qjdsx5l3J5kgwTQXjS71hDbBgn5EmBKhFxbWbs8OWX/Hp5oaLg60v0H
BPeWFxZnkl/jcWl194YRQlEMfG2fU162INC0NZcvEjP4EELZVZcJJMpIeUFGXmoQ
X952VNDqmcGKMJcP++u9LAmc+ftBr9tpEgwQFMEKDZ9J40k75twrrzxeAmXQFT1m
RM11DAFdx/RUcBwZB7sPLDTHE/eM2Sbku52PxxcnA9zVveoUntjQB73qFLcOkm/K
iQCez+9BSFiI3CcK3ASAemlNjzb8i2MSAZzSo8Gx0ib9/q27PLq+8AqVk9uRcpAH
pi08s7hRZ3gcB7who3tUXe301a1pZ7Se9JPFzt4Agi/01dRWNyGnoH/MwL855z39
q0ZC8XJNnhahEgtY+n13C6v/taDxmA4Q4lrkCfnGP/i5LLiuk3ksAYZchbpWrC4v
rpn4feHUBigVOuJMjmkAO6S8VcfmZlPoABTPk3K8t5xSEFNzIOkUcwjZqO2KO3PZ
U/51YWZ/oPud9bXZiLjJ+fq408uDCyEACoino4rgWXypZkZC6Zo6gWlJI/unzg+I
79pnWq++azCOQB/897365T4zADzsJ/OkjBDi9n8LMBRtx0TpJ5p0gs3jiHCKZIcD
XtcNSa50f70qGZ2dq9qJsktF4sa8kDCUaMzF+ACkqaXBPr3KTH+mosRW/RMKus8+
x8iO4IuM5PE/37aBcrZouYaxGNQBMFs0UQkTC7sqDcP8uvvz+fvMKdXEgSwxiezh
4nK5AzzIA/YVqjcCoIWOmrGO/vDSWBEXiHAv11XB3G3OAEkoD1a0eUuNgZIitRjw
7hgSGqv1pLgYqD4IB4jByzBBE/ceFV6KUhlQQmYEkxHCyxpO+81/wnKlHpqT0JE4
KuwR+AWOzmJTER5BcoGzrgzDURg93BX/hxvpR+fLyn6MTnDW5UIEuYfszJEsvo5Q
iAyAnT5w/8wx3NUAHUXrJJ1kMurncJwNpcrEcJ8p27ZQ2inWGJEHrt+FI6G/+KJB
/vcuD9XFJHCZuPAt3o5r7VxXuyn5xfIenC0P8yuEXYc1sSABQEJ6fsTMeN+V/jyp
4BzfHEl50uwPCBLK35TkiVvFBR3JJQOxH6CBpP+iTGWcad0uOjeA7nx7bcIWW6Jx
Ztb3ea+kxftNKIFuQRX2hJJdBmZEAMkvIgvIG8Nl6RJWmBrDXELzOVH17JrTAo01
2tkLO2vemLeZZkS+0OBXzPfb2yUy4+5+5ytLzHjRJAw1xCSfSv26DWQGS/684qvc
XLuk13N9g82+8tjp2zoyH+tBoVf7BLYLJYp9D3aaNRX6wn+OTynO+o44fJuH5w01
KIRUZ4UiNoDLKf1bjsGi7u94Is/qPEcGy6MNpKqHfA93HzrmRATxbpPWiw+DpLnE
p68IYIHYUjKuTi4n58nxdNm4c2nohP0TEWTl9S+mPToO/9gX3CuMP/4mk1t8q2QN
LSIlE97u8isM+kANfyKN2Wu5quaTB3j2ORXIKwtWEoXSHjq0tqKCFxyrZAYLh7Nh
Y5uQrDRhyrESWhJb6RtyPX4RqFH7w3cUE2qdUvBr0MlMNHhmETAleGkxwRFbwI2e
cAHM3TSulE5rA/9sB6RveY7xJDathL3gXzRV8A6g2znRjlCwSBITE9PffRucYg/H
WxVK+GKGmSuxTW4kx5Tpdb4T/KK47nlbrUoED8H5hCf3iDsLCV6IUMZWsjVUuQF5
q5vMcND2NcTce31f2MUOwKaONsntmnEOn61dfiVeD8zHqh33KAFxgBOkG5525iaq
Zikvviz9tFJpK5qkUiKZmMLnTHIQNBbdXv5kN7w8+Z/KVaTf7p4Uw8ZsMvk7GBZB
bXsU4pQfJTCCF1Q1Ms4bK6x3oSFFkA80pkynrBdUTnP62Tw7l6h6EkRyymeJkCpd
n7n6q5OzH6z0H2g9sDqlXYyjnisAOBL0qsRnuY1FC/7vfpxa1HL1kp5PgShKHslK
XzVQ50Egwm8tlDP6HNXrlj2ghPwlL/aji5YlHL1y8WCgetVtEbXt2mTBoKonwIZZ
7W9SocAzBUixYaLgzMUzYErlDBVtE8qt4JExFivnYQBkZAGXuuwEYs3RUxneLhAP
6cDw6bvY9xxgAzQ2ogDqC/+bWGukVQ/R21ea520FtnD3Q5oJNEyAc9m7rPczaZ8C
+wFtlnOupWuEMTzu3nHxR+71/fD5AfinSK1q70BYFAej6K1dsB1aCDCMTnmhChzO
L+ameIQGCOWH7r2m1D9oMxwVz8hd00u2vSNz1TFP3alkr5zntBV3OEY3/BCcN7SW
Xjeoajt21C2+N/5qsuZek59yUGTpuZnodfebGIMTdmoxkQSmz6RslhuXzWXV44GM
XNenSfsFaG+oiG/W7HCtbBihPYE3N+FslqSiYpT06Qkr1fCdmbmKUgQHj2h7AzUK
vrMExz5g/aOw1dpEMU/ERLELTX1iw6irZjnbmv5xTjflxWp88fffuWUyRqHNlyX2
IZr4xtvGtBBMVz4i81F5JehKCbIbzPxf8KUpSicEuzS777qFU+xUhS/ZWmoLaW9p
YdwvcW4flR6BjmFoebV0UPHQBaCdP2tpZksQSNMh1NOb6MJR/oZPaBWPtmVvYOqH
ym2WLd+y1nOe1eLeQYZgz5vWza3L4Qgk7h0WXshheCzaCglrw270E1ZVhav6s/CA
TL02BXLd9BN54vg68AL/7CeYw6HuE97i5uQHJT0R/o1MKpGx423nv9XaqMR9bMeh
QiqfZjKP8kII8GKQNjzWZJ0itiEKjn0aBgNYmxO+BjyJ0YF9RQNMZnda/OSPiJqP
KjTIMTai0VD0oFolcR9j5qNPPcCmB4bR/iT1QGlrnaTBHbbfV9dRh4o5DjdOxJuy
GqijuLPsgiN70Lc99FOzWRTrPv3q3FswJQDPpLFou48Of6qTBWBdSD5PmsxEKC0M
d/xJn+YI7dmPpIQh/2IF6gBnxZtlpLwYPGMwj+hi3JW620nAM/e62KOkC8sT7+RP
sez1wqc1qT6Ff2N/K57lX8RYY40nRyow4WFb4d/Ouk3SNe9Uk2UVVZmfcBEU+BRq
fPyYoITYT+J8EOXyVCR59Fxk6z6+4iY4pFZNt2I5UCW95A74Rb/JKLYo3MgbQazJ
+uAvFi31WBvpnp4NIlHXgITiiIq8K52ZbC6wBc/bsQvniFP/e1lq/rWmWysPlYiO
rAvaeTsdeYWyAesneySQ2yEAFv1d7ewXS1zUL4MfeQQwPN6knXS8L+zxubnaAd2x
Gy4dCWNCPkuD5bgveekFrhmc/Kz4dg+/FiqgD+KcvrgY8LKKsjA3gjrPKe2LHYOH
it/dGgfzOus2XzgsIL8P54DB4NQ+HqCr24LbPAOzxNgRz4xxOVKtuHwDkoG1lJd1
9Bwf+qCkYzgwrG3wTPvWm4gfgTkUks/Y75qXdjH0rtbtXORQScUKXGxAjtiVyfTX
qvpVotxn83pAH0+j7ngDkVkY+SlsWoF2vm25LLMWTOk048/1dhTUG8Qooy0Wow4u
IqQG/dU7h1h7v16CvIHpqVX9mU0htZDJ6kw8IkMUufVnyrIHnEtDX+GPiLJdN4ij
NOBzN0wFWcAizuFtFs7crKi8uKIukk9cjXnhHsv9rDCl7qiF3iOVcYiKCXi+21rB
Ns6v75yyX8B2PN+4iiR/QA9s2+8ffr4ILV2gO5FJQpul8WlyePkBVKgHu1aYlJpk
jE74iWZUc0xywf9eSscNqzIu2aC+l4G6+nS0gXnbIfgweOyW/vnKQ0vG9fSKzGFy
j1ZbQSub59IuqYS3yFQlEt+Tw5ambwjCHw1XEfxPD5rtK3P35G5G9MPq4+2CAEWG
DmKZHdvMneHU3/mH4nfieu4N8DWfcILeeZHM5WvTPIJS4TKFA2eqKXGW08bXk1rK
uJEaNWGqdZzSnwMnXHpSgpMiDFozS0tb+hTZIknXhKMlCas4TFZqqzNl0j/A/1U7
np7oAzLgM8zOAw+gph9w7ilUPSMJtqCShXw36VMfE1b2qbmugrFfOP5qco3usHSb
zn95t/SqryX3aqBpwekKair514SBM6qOeEVLRsYIZJvrNx+c1GD5tIN104HPLmYq
GoSaBbRlrs8RgdC8wURcwUA1+o/EQIa/10ytbIiZvw9vyvl6yiM7jc1CfqhW6HWr
zsJLagXNBsRJGwL1qE74jz9Ip6Fbc1aHLrRVvZKvbWLPtklFIFuz5XBo+QVhK8ov
5MCTYRBo+SF73gnH8phaP5VEDAe4oMKKknw24/zuh7vI0Eqxp7ZYAqaydSiBBsCO
IOjz0GxYSYg1aGIWEeZyXY4ScI1UxjyPS/A8ZxB5qPSF+A0n3qI9wMcBEYN9YAMq
2/bx6AtpRt9h4EfyykTHhUmPgBT/26vwMd9hpsxSB6Yd5tZQJMI0gUWcczwaM+hk
LqJA3OACmOCaE7LFrTzp2hpih20lGDU/vPn7GQzAVpO84WAii73SIEXi0DfPa5ba
jobP80OHF1RxG+iLabyfcPgpxg+el/q7S6M3yaM9o5IDyH1wMeletyhbkGlpbpQO
SX0gXGlWvzLdkeZqS7sAkoo0zAeQFRBteQyWK9QSwEPLhaXrJE0xVD4XhLjnF8i1
QIPA5iXYRGFOagaO6Ncp4Fy52Rlfw8jd0UwlPzDeGfj/8BXnB5+RWR/P23hX4qc3
i8IQvKzyR0xzSOThGiZIIv7VSJJkvAj4PUWwl5P353JAPsE3evnl655QiQEQdejo
GcfujLSM//vzELBCVy4Wr3pr7Q0kOkuqY0JoWKkYRSr7lKZbOGm9LrJa9aHI7+EF
1rDXNcGMLe8IJpsZ2ZxaL2qxn/Va57qyzFPsqJPrCUaYdhv4ulRt1LwfUb5xoMJ6
GZ4nEwgJCVkkkA1KnG2l2SSzEM6ooRg2vgFWLpGKnGIiNOLqKAzLok8suAgaaKpD
K8+hPHe/NesxOsq1s74HQeO75OZlYbd5KxQqdetpYrMdncSbGCLI5D4V01fDCqpU
5AauXyV/H89Sg8sMtlOCO4PMLqTidfU9IpsuTJ3s/EINocqt1dXdH0/blULd5wLr
voBb9IhGMXGVAWk3k/3c5uB3TNfPj2CCAlz+atLswTQaW2E1XUbO0So7riPJgL9G
RenSkqmw+woJDybQrbJZ5stJVjna5L0Gvg4LD1iDifk+5Vk6uZQVQznfbQSf72NS
Tr7gQkvEomdIKdhusVZN+Ik9fIhxN5DjX6foohMGRRYXDqf4TMJvVZxKxQKVJ4HQ
SjcrYdY2pWkcMsrVaLnNNhmsG4S68XseOOgZwGGhbuw2kwrs+kGfLJKYVVSeG7G7
IlC5TaO7DM/2zAoN0Ro9WG2Rz82UH2gbSYidOICWkTT1EcLuK/e30W5zybdK0l62
+7yetD4/x/Us3M3Uvc3s6XXhUQgslY0V3bSxIUP+LBFgTPKOqqhdqyxS+w+6yqhE
BewKCxYiccV+p8bkwO0Fqe0rFnCHgFdi4ae5a8PBiPQxbZljNTsr9OdQsWqwlrBL
m2D7YmbGyenCcVY+kfX80bNAuQZcc0J9tAXf+yh4Xutp9lS7VYZ8EXjeW2S2xcje
GVtZ3+ZIuLtxW96lU8xJZhACtoa7CGwgfPMhdyZd4V2JdnEAFbG+T0dLc2yUNPP2
juhaeqkpub+qAvkD0Ef0xoROHVW9zdnUXSSeG4q4FlsnxCT+2KEhKeBzHevTtaQ9
Q5rPWoLQXSY3Y7EVrb0ouV7frEqugY52jYTSj0Ew2nrPCeaF0C5Vnc5kQyGtqHsd
eAcnjQIXLpO5A3K8obfRwA388MkIfC42TKf4LgoYNL/8TArOnnABdKOryqKM4RLp
`protect end_protected