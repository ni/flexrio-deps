`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2688 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
oechCC4pIyia/5VZUUxROmFZfxTBqhEpEiYOuNbt6yyACBr3BiXrm00BSZuREeAi
VsEfDgXyC9aS66MrIacEP68UvXMtm8Otnn1UuKLy+MSF4Bd53fxr5VkXzxlfjy6B
JRjXquMKN4IN5JqV3kXClzXG9aubmiVuce/gcEDoqcDpeUAoZDYw90KvDTcZcnWA
sX3CSiUiAOfYWAr9l97K/Bv7f0xKNBDBWryXN+spDCr9r8vmtw6Mb7/ADPQ9jMrk
uXNr/H8xcL/SRt6duySNyI2aAJHZHjRj60XRPk/97v13c4n6ihJ3TzV2tZ8t4g2n
Q7VOE6jqMK3JgwB/iQW/G+KebVDT3mi3iiXGDkSmsSQqkeEiYenz9e0exJ8i+jzL
kkmz537CIJ7axAEYsRAj8c6d5G6rXF8X75DI/mMG/H55vauI44z7Rh8kFLo3tSv9
7R/GwMA4yKUB1blNjT+bHtJOV04R3sk0GqKjIzUdjZI28pEndMQr1EKWGFrWywJ7
X7L9GGVjYduGXZd7H7mNtCv/JyBF9Sj+jatrtmy9RdY+S54GUEJDOrWIwfSWNxt3
YxMIwHH707Ts0cKnLiTnfe+5xqHn3sJIKyt/qagUMnpTkhC9V0THG0nJyRiMI8xF
Gv/zCMqybBheIypDa0voC0ezRS9HRUqPiMt2Cpsr6S0Vc1f19eNecEcoMk7NwPdM
UPz/Ll9jpgGhUnfxTcWmkwlIwAQ9Yq7ldiuh/46e3+nK7n9zcbjB/MJY04Dnb/J9
C/s7KlqUmAv2mXb5sPTU6Fsy7AVyhHaRsVdtiqXBGkBkuVHr1Itl3sUjQwhhyZD2
Ar3D6uL60Q35YfJz38w3vma5K7g2g66lyfiLmAKhOl6mz/osvAAmnQZBUC19J9OP
2pEmKg8RzDOiraXymE6T8KGN20B3hvdaNT/sJjC0YkuyjUiXbCvgEZi97eu62HNi
IT1sQYpCetOYPlZh7YdFlV75O9lg1EWC9e7W5A1BLCQ1Dl2YPeTnpYk/ch/B+Fws
kSt9lt8ZWpuNcmqA24EgGNwP0p3xDBLpRUlyVtMxXH3S7JJ57ujRAUz9Rdgsxb5K
IgDTAO/DZYu183ZISz2d2NBBC6BPg7cN/aopgDeGvEllFHqbxXpsKyEJmH19zviW
2apxnDAKM3ilfOpWpkXKpBq2UzbHy2AdO//w66XgClc2sfU7syuae3fUfUlktQ51
mOIWQJN7ZFUxpioGP89bBHnhK6yOkk8xniU9nm56AdONLG0HqrzENQlel5ku7OV3
jSxNuRBq3EABdWrcr989P+AYfiDPYWt0Vd8L1eha/KYfdDfrWQSOCKXWaWVJZ0Ip
TGxfyflRhVnCWt+7kI8zBxpwng0hzw8uxlZZd9z78/7gDGVMfEIWEjBh/H7M9pcU
WGWEfbo1xzPwcn7hDmX/GWpB+EzXaTnUp5zwA++ZWZRPIwwT47uCzS2uUZ8VAgyE
eWl/nm9U5GO/Ypj95nQ/VtyGqlMtfY5TQM11pQRB9if5BgST4B2ZK7XOvqS6K3Cu
NBjkgC8RXoocCa3VSP2JGZ95eweLwV79NeO1PRU6ovV31WFtaEKaaRgiRCm0JuUc
hdHJHSk1eFlQC4Y7C959gdBTz2NCO8adjS5uonil9pJsV3ez/5wlt8I5PjTcyVsl
WeAeAs11Sb8AWA6/e3LHFzYuVFHArVqW64YuK5srCOvH3i9OAWwQFtLxNsG4LEtO
UA89v876RQALFkyfeo27g877PBsAzwV/H4QNaUozlQNxPYs6LNa5cPEO07dCZIPb
ecJG3F2flxId23Jn9TZomPdIT9mxNoeVVVP8u7XLGtAccB4mlFqZRKETpUUrpNPd
9fOPbNTq2as9vxOTSEY1ix/OqHaB4vyifZjlt9/hxziGHp+7/XOUVyySMbPJeIzb
THmB+H4JmYJVomSSMY2HxuZ7zR60J6lcyt0BKWtDT1spbMozBrEO8NohShtE3Ged
dinTy+KUdditbAv/wcLQACp0ma47W6LdsxU9le7UtnK7Z+LWrJ5YfQlnAhLbSVOj
2Se0DYd4cSB8XpeM/kVRrzH23yD4hj66uG7dEKGMKCNu5eyoI6OFE7PxVCVEXUHd
h29wWi6KIn7Y4fel+3MOFD5iDbQ/eP0P8N1vV3Fuv3KcRr5M2NPlKxYvo0TtDFeu
iZ1U6a/YOGU6ZtEA2vZ31SXKkbqRohwYXERcBmsi2iMXy+zB2IHoPpd/IBBz89iO
qsGpZxLkgd/Iuugdj/nSgboGPDHboLbhn8QYcYdiNxSxkGfBB84ZcMPbnQ44mGMp
uCZCw2D03BE8nsf0bNrTPT4DN8/J/4EImFyMaoUOXbg/z33HtDisd35P9JfaeP/T
yPOCBiKi+gMG6NfTdXSfzKjjHu92j4ke3FdIo2aMtL0rQp8oj9kLuAsFtRyjByLL
FLbuig7KLI9wc1n2Ndg+Zdc0JqPrVp1CLzDc/xG4EqNW5r6TOmfA0pHSqDNbaqhX
y4dsMXB7XXN1Un3oQvll0aFcYydmFiGmn8j+YkjWJU2xxL+gliQrge86Gpm+toTb
B+So+t5s8Z3/LMF5uxPIALlK6aGVs6bYV/mAdWXSOIBGWtL9gvEez38iW06uyaXZ
y4IRT4kJyCSFOskop0pxXK/62UfNZEp/pCdGgzUWUo4gwjg2USJ/f31gYqqwBkSu
cVpJgNyrQ+EBE61mmadoX2sCn+2u3QsOXKUszMozq4g0uYyuHwvrY4l8ZGLqyOfk
aNJRw6/3TaS7WIG7ETZwfE6C/CQnhPz2DG3VqRYwWGJrGH+PIG+rcK36jmwZj+GN
qy0pMXfwVA8tn6pa9MzMXTaUkyjuVFkmLSAkouHoAdH5U2B8YBYL8be4jYodsebV
aLm+vD7YcyI6qE4xBM3KB2jxoZRBBhnArqFJsYIev94tT0pHl+kcH+yDzrrG3UJj
gjBGcpWgcKkXjlx7I2CXcF+aaoPs0QGh842ilfPdoIZzlL8kZ4f9ynPpw3Nl9NkZ
YfiXv6KolirJtOdWqFrWyCYW1zQDjac2IXwWPe4evkSgDNiH1p9ZK1+iOKQGxvxY
gf+QGKsbuDNZdBUAAbxZbuVlOtM4tU+HItdpMnt9cNtMVITIJICtP/1b1GAWpvwC
t1A66U/hrhi1YCLoL1o1jYxM92U+8E1S8nPXzo7n2jIKdu3SHIA75m6Yk2TAmLsz
z8AV+asCs3jU3ZHPZmhpmIzRHy9/mMu6ojIBMq0FGbhz2QdK3xATu0+bNWjhg6wk
ZY6lBlweU6FBRHMAx5G0vFOye/Qj+cSvYFKvpjE7q7+h0Kvnkpo/uVVfpGHlKDae
30hLX/BaR20cDZjdWD+MFn7zT4t9oJME1N4WuJi36vbnAhM00IoJ446Ako0HvyCh
FzgxEq1ry4GsA3G3HqHfLmACbiq+cxWTmrh8vhu3ZLRvAbL9+P6cf9CfgEHPehKG
`protect end_protected