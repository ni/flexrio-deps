`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15696 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
MvRQqf28vVzASKXcuYPav6UZkdjBaVquNNzFkAKlpsgQ32RZwq4ZwY68lN74WzTg
6kVBH3mLaEHy+9DVVY5I+IlF7Er6a2Ad4FsQIwzSnDYkR8o4PtwH8tSUEL9Xcqt2
jp5RogmWUndJYEt2tS+blGvQurr+q8KF4RMMup+tv5XgKs+yAWP6/B5VJpY4prZ4
JSn14j10pWh7+DXIe0jlOwRSzNuBTlEKP5D1FlCyfaNAIuwzi68iCuRv12CMjmcz
J/OPlV3MVVntf0vLHV+ioxECj03paXsh+sdgmw9DEBSnSA5vSS1nJ4i5NrWVCgiJ
HekB1SKfGnLqUUmuF3tWP6t5saPwwe+202fY5NN4SaJS6m+09dvHg9IK68vOMjSp
j4t8bO2WruMyfZmNGt5g3ufrlBRzON313muCRE4LUK4gsNyBLNDICmC7lQIKavxM
eHcwmtXQ9tQyd18LqtG/bHF/YxbeQg9ayA31RqS/p9Jlh0nDI9z2l0uPuSAfW0Rz
yOl5NQ2Q6bqKMG3JI5xyliGnGHKb4plmM1FGeyaE64jOwJgFQQRuzzKS7SA/6RlR
DC20wfij0w6PIjp65UQ0V3G9C+LVva+NF5lRBy5ewS9mHnR81/APQ7ulEKjQ0Q3Z
DDC9OwwAQVs1D+WV2VpGX88ToXD6j041kYhghCZUhtPPKtNICd4h3ZPWbehoObMP
No82T/v8L/0b7n7ybYGgRHOwK4ktXjLDh/qV5yxqRuFqxhgn0QFFSvyoN2l20Cm7
hrDHnngYE1nSJdl7MoLgnx3SsOfVkkoq/CfULxqvpAWqFcYu27ya3ACEfUqIE2Ls
8JVnvP7/lSOvfJalquJztZhao3aw1bA6qlMgAgG9B5JDkqBolD/m2gNVj7zdcDpd
fyYWSjc5gkFB3pDVsdz27wiqXA4u1qFysvOM9k2gdDfmh9SKXnGyx+CefdRD8N8j
6lqE1d9M4dWGJh/iwJyVXC6TnTNA88cE/KzKWZNIIeun+EQ8NSj0dz9afGe7VoeI
BRXqzKlmkYbsHTJPG+woyN4Ojt4vb11zZxAm94eHYwPznxbXMgO2EroySF1vSPYw
kV0uIfAdHliGflOpbkWud8Q5oB5AEg/H2UGkEBU+8NG/4DyTB7JaIcmz8oDQAOEV
BFGwgy8RD4f4pXgTs3kwGqFsxmWtRl9AoJmKN/U5+eZSbYsdDa6Ksvh4s/C7PLR7
8Qnjq440/KeFJKU13j6rDK3ZO/GMlnYjaQeYDuAwPOYRKGKthOWV0cywIzh5CW4P
wLYm1JnrU408jV8yxNVOy6hF0EnTMisCeVsqAUJWMLj/Blh/Dr/+z7lVUJ9r9t75
bucDnszQ6fPqt3OY/2wsflJnqM+wwRIDX5ljP4dRfrhNd/bJ5IHqiNnEIURMFagx
A6gRQO2AmIJLLQE3hMMkuq1yGeddon1ux7yq6bkd9Xt93l1gZPWNsh3FtavRPjAS
tD8itp6jStMSTOgTD2Nl3g9pmcxWfkuGHqIaskLnD2wkWHu/vd5VXn9kmEgmj1nI
BNsHXIl2FWCnlWrAsGbfKX4s6Z+qQi6/Uq28EWFhFyZxBNtBgKOUeaTrmTA4Kc3a
9edZftvkOTcD4IlCIVsdUGoGfw2ExU38wHUNFPUl13GkRk1AXphe02WcoOD5aHy1
4o5tlpmXmRsy8GK74t96Bh/WdU+jJuoC5Q/HJ9quRX2ieYoYwm8GbzlYpBMBk2an
gcouTcnR7dMgJPU44Uff4RTcUWJii/ZZN0Yho/XwMGq1mmPJkEBBDwDloPWWKkHW
kbHbWNyvMlbrMisO7oJL6pTx4Y/NgwnMROQzBhWGM40TMu7f6wGYGqur2Mkrqj+5
QQolnETqoVXC96YAzBiJxRKUw75gWYNx+5N2X8I5IDBwCxKqNYXmV2xf088HhucD
BL8O/XkTVPxKHnWrJLXeA4fNRO/jgH+t3VfN3HHsXLOh5mNBFg0te7YfxdUf1MoB
rnQd/X26z7cToqAlcCM0z9JF7oyKpWZb9L6Ofbd/lgaWqWjH0Af3PP7baBBMWHOJ
3KH9w5act5BWL6pA/Fa6dKZjnedKQedB3MRSFsAk98gDKfJ21bN3wqnLipDGq4vA
3diKjEFNKYVjTPCAsFosVu5qzUr9ytp52DoxzYDpo0E6GxOa+QUirL5peuvV1CFa
+Rkf/JdDUBdLiCb4oyQ2agih//B6Iyvld9W+L6DIqU/cQ3wDpLeyUJHObtOTTCLv
wA7yppEYDJtLL6rv+R0gklWMi87wUQ8s1fEPV5BOZTaNqvN/9sIN+Smzxm2182Ii
lvepjALBxhEHg0tM8di0cFLprkstMSB8fTkT7YnlZXZU8W23EVx8lz+V0pRjb5H0
TIDkL08dsLscjyEHmUdZlhMljgHxW0kN1Q2ngCvr+D9H7c1In0tXyGq5xkQbOUBe
5pViZ4exOyVc3OWv+jRXkrGgLyG09RVtjbHAzIVvhctdS/gRnkBwoK+VCj22vrk9
zfeyvBvAzLHQ+25M2SF70cuD882pwFcVWZDKe8VF4qIdO61L2osoe91quLW7JRW5
ATB3NUB4QfAZK0nDIDF+iOodkYVD7zk4J4Dw6c9hvi8dYZVXVGfa0gjkT7FGKmiL
SKNRuXwZO7eKvQVAlaM3PEMAMBJ6jwreGjJknJ0TlXAZOh2JRhVkte808h/d4i6Q
wxgrzeovwsZ77fqPaEzPabXtJMQCOnkyQBR4MZ2y4THEjht4oKk+HdJAvcNxjMp5
Vlh6wswYGhqvYrKtOVStXKQBewjWflcakZmrN0Eb4BMW3efbML3XD/xg1a9XK8AO
iQtf1ju0kB/GAV0h6dK0+i6OZGOe6TGNobf9lVRG1XJvOSHmoKjDY54Du7CkFRs8
ytSBbthM06S/u18QsgOUPBghWCEVga5UZbw20dHFNmP2svaLydJIm2gUKiYRz1ZA
L3u5SWeBMSCDwQ15xduxbAOnQOrHu5pKr4C4XQhFQVC7X1ZFWk6HtB2fCA9aVA4m
QJdyV49uu6fWMN53ZHKYJmJSGruCRwr0KVudXYljx5DIvtt8vKPuTGwbe1SX6MYh
Sv5GK8b90ZCsMyhf1UyQDyLOsnv2U52OZvS9jnCXCvWyCg8mysRJCpvUDhYmlk5/
G9aYxjP82j/ODheDZXO/0xT4hODpcjM8f4tdBkQlVzztkOLPflmR9ng9uXYpC/6t
RcigNFPfgFL+nieO0erQJnfZRhMWm6+XCYxw/FlOVr1qdOnjMADcRdhgZKuwypHZ
lX8X8VPTGeaTMInVeyHhBXzLJWE2PJiFQXhS4oOrkVpKRiZY/JfA0K/YWumpuYde
OTcVRz1TkI+gxLkIlUAJiq0yqcMcgsYp+xeGO+2JdcjH0QNcqcclkfoJ90eM+Dlu
WUKqboS4+uCfbr3Px47bJOi8UCqJCiTY5a+6bSCmeo9Xn991EiJSjxYSTP/mOgnu
PNR8TfyzzquE3CQ/fHHoXsVeYI7nFlBENCudaHzYMIgJrOAc1mYANYQPLlt5e6JS
jtnbaZF0/4Eu/ZS9Ma4STYuWepH7BhvIDT2DJvtpV2HOioyE34EJR+B93/LArQ5T
AeqM3SMtUXlrMas7S4BLkbI3TOonw1Xe8CG/+iA/fLCCHWh1SF3NqjOjNAag2jV+
HwgPnf/nWn1tQb2LWYjm4MreYl7+Rl+sRtcAQoen0N6AYxw6/mPMfzgKmDNKRvcb
cs2g9FNtN5ZLVVTCtgQvEQKzOkqaidVzgaWHJmXNu9Sh0TSk+4j1koZ1HnTWMnLk
QnH/ZTgyc98Ak6JqBN+r5PwIm7YWoypO0e+bTls8teqk1+yT1ysIOsbIEI7EzxjZ
1n50ZjM46w0es7O+CeivQL5zp0mOieTb0GSv2sj3jqKunycfQgssaro0zbG9kUp+
0qDSV4XcTmlZlZ3lk3cCmW6uRJF4B686Dr9dpqjzlplNyIQmDMf3waQ1cK9ejZna
7SMvSZBQf35WfGcqH+OAbXIf8+P+oYmt+AwwdsM8WcjvX1Rj4Il+IcihVM2PHyWI
9K7KQizRdaXr51Fm8dhXjrOlTq3eJDf0kza+F2D8DdPAf3gEvzURlRq7hInNFScq
qM6ZbvapIyw9mu4WUvX0M9zpTOOXZM+gBR549JQhGuXfQmW3uCB0uB0YadA5g6eg
fvGirE16hLRkFjnLWKGYMOl+6TqBtQumRAcM5ER+BNokZ3UcVqVpimUEK5oYPtSk
EYTNHvc+D6Aym6t9oVRBshsmBobL4A721XnR66FVf91Yq3NCmYX6hZjlzqbDwdn+
+TjOxgqoV2YwjFuk4s7L2ZxcNqwuJgrc9gj4v7idGgPZaUYoLnUE6ENzlYLYpu4Y
KRqUA7Btz/MhVf6xeJWqg3uNTUnGQkhQYGOJVpzP70q/dgYPYxfjVksQkux7aHna
cfWBhQj6isA+AATY6PFL1yQEc78of6uoUmLMzsbzhjL2aW/23HuSdSikjfmTxEqs
uOp94edlTeitnG36nthW13WRULM0SGqJH8uSxnE6lTpCPb3LEWa+FhgCF1jgeHau
4HZrOWS7i+Fbn3Y77kKA0vVdigzFa7zdSmewtj25jH7RYRIjZ9k6OafSn5xi32wy
dsiVbpzxGJF6XDCnnjjB77NSSoCHH1PwjijX7dG8Pp/EyfDB9gEqOcQVenoNPHI0
B4Pt7BMpf/mw0zuHgdEyeFV07mbc+rDjxQQtq4/KaSLqyMfgSPqT87L0Xhxzk3s8
4Am7zre1Ukj5DRRdVZ5nele/ut12a3l3Pjrruoso5u2Bsxx+2RJDO6YEywBNgfm/
JPw1MTN/Q5+l4BLNOwNTftCMA7qaNWCV+iWxh8x9cbqvl/9Gb3fGapeVMyOOXWnT
QJBU4esTiFHPUxpzJWVHiILkweIxivrW3F2XhWi8lon85TL/j1waqoai/WHnjFMm
7ry6jFISU+/84elB3qmMHcU47hI527uCvPElzPIhg5oXKVrwSJoFDTJmGysvoQRZ
XtYBfFrwaUW6M3hTeQ9DThGp8suhZXlqIwE4hNJNSbUbeFThRgtdOeyLUL0+zWDS
seFn1jOUjUaFo2zZUVxZLBCIKHv74K0k5kB1H/yzSyagsR+eDHmfbpCb3cnfmXCI
QOHH8l//bxHgy1/wW1ybSK8wpH4kr/HnwmnPrEfzolbEkL0UaTpqz0aMRGSTHN/7
35f80nR5sAmGd11y3vlj0suIUUxNQif2ReWYD8fp8rM0hvOTrzi4eFmKyzFNGWtC
X37g2JgGq02QJwSprQTao5QoI4JTg96jaWDuaqPC6Nlpah+bmaaU9+l7eNl5/44U
IHXJfo4N3MxLayxKAVIsKjFc9Cq3ejByuX2j8PStfY/9oNRmaD4NJaRb5mIVbzgq
hJpd+10pfhEKS3JTr3P378VuRgxHO/RZWXIlfX07hBueRZF9Goa/IquUeL4w1XkH
qz9xluyWrFI+A7Tzl4YUgRhNXC48o3ooLJKXkuGz/mHohIZ2TP/7ttHHuHDlMsOm
b5oEnrkg0ylzFKasgcZw/EZFi9sR7n24Uih+D/GCyD+7WFZ6I/zPoWus7G6Fy8Uo
58IURO/kKRLcsymDbV1BrFdv5+9zzW4AoGIBF8mEwdxTAEt5Tg0z57iM0k0iP/aS
Ky9JKnZytXGQFBNxLxXfPHagYrKzwuNKlNmC+XphoP0hE9hBVahQH3OpxgQevIVe
2F8T1nHRwMd754u+fXoGAIDtZNS4z1AQOzzBwoJRg08+vj8LY5uT6l573rnJ9cBp
Y1qXbzLCVE+W16iXinMhxNyxD0fJoREjewt/PLF+t71VaJsV0vYe78groCKPegMS
ckHRb9dHZyUBqVrn24w8JWWtSVsbU/4hB02WwinY7IED4PQh4sGpyVaJbdoomrCS
ZYxWSsTq0UoMLeTHIbY2T8fKqtXXyqJP9lnET2dSwGAY6JyzdXN6bxUPKyu2wftn
Kwl5AbmmVxoP45JGKVyvKEzEUolAXjLmpFKkkej71TCwfdNFJRmRdm2uNN2HuFHz
BJr5K/i5ad0WA/Rv91CuuscNBm6RprBiWDFQ7oKbeBP3aLtZIs7vr7CmZiJPn0T+
ydvu23hWFMErSzGk0R8VvBmY5KVxPzAAEbejQrZ2PyVmECJ5tKnyYnYNRTQUnNIn
9VfNLX899Pf9J4q0ZjDa+a6vHlfiogF0oo9zoHnlk+5Ja++fk4feO/lFCcdNClKZ
Wa6L00m76bgFqYdd6l5zLJxBegpdLy8F8AxzUsP8fiAGQZJQ8FeQFV+i0YhHIyNM
OAR/+sn+N4fa8j0D7Jmk8/XDeNQcXn9CyS5i1wE1qWk/1sH72wptKkh2ka+AuKzp
3vzeJ+OmcHJ6Gd1Es9E7rrfoe6OH/rg4t5DH7cxePqrTaJi81osMD3Ldu/tALCpU
5JH5FnDQ3ITCW28jg0Lp2jMN3VKsvma5Bs1joMs/gl8p05mS/MUYLe1Z7207Ksnp
Ee8fsmnkZ+oZTsRB+sRWRA2BmxyCbttV+rVjLkbtyA4nZ95U/Ip3CP14k/kV9HUQ
mYm5yxu9JzVe3kEvu2shAPoR8cPvJo0ot5e/FZtSHuRBBVg3gBXHiJ96OBjPoHZp
pN9gitvPaJrFnbHXrQ+U2xe8JJxHxE47C3LQVirLFmCV0keuh8p89LwCb2KpTHCx
/rql0UbQhxnZmi848TrtntYz6MTsIQMZt6IBcxl4lwOpgMBaBeBYLbr3JlMc0AfJ
aFlg+/qWX4FsiVONtn636lOOcUY6hPjOUNkNdzT3qUVBgkG3g6/LFfoj1iYmRrPm
FvxrNmbpY53kmhIiJTrbNaxQCUKgMLYbp7BqDwhybx6xq8QO+4q/62PbRRbr6hGJ
I6i6fXwwL7ZaGAb1iiL8JpkjOGSuNIq8HTFZlgKXbQBIS+vwpmiKb8hmqgh1klVC
NNvJ3hKdqiV75mHJ8juGSnvW5UoZwSRfHakUB65gfJDw6jrOL2PjOJN7OwBwMje0
pUMdkaPyED1FBa9nWbfxM4lOu64Z+LUyaOBMlKtH+Uc61EwlEmqjmNamVIn8K+nF
6zqsZb5qCL6bOdi7ywFgxbdDy0AOyMs/RGJWXUGY/qkd1iRxOHPGk0qkRawjq/Za
ikjjLqnQUpw8JX++nHHI/By0a6VRsZlkpya5IJ96CUgI1qdNKeyUEbPhV94nxFXg
IUPraOveANhTEFoAa89BNfFHRzNi7xD6H8kyiahMf0iksf5haooUjmu1FQwI1Wz6
mqMFwGDIZBtjTIvZn12ExlQjWglE22I9ZrRdgdiPdiLnqTZoOw+tLhzDRujltExP
D5bVLiPy6iEjPo+NspCbZ+FB6K+5yLuRrdimmEiZl697u5sl6hFYj0H5YC+h+0za
9dj1hy63HQ4rW3ILCgWENe/bplVSshM4wxoXBzk4eqxGQBsov4DgsjndKIQCz3sB
3+omkDHZTiv9imvwZE699a4jfZm5fnhe5drPuK1D1DXfqkzpsFCiETcauGXeS34M
7xGC/SVI//r/Y9x3aCbb/z+PkuWwMHU/R5B3P7RyqzGwc7DJNquI5OQGwmWowl4g
20MBoWvcU2EBRTsp3zkznNNrUxF9WLZYUl949EETvTOXcgnvwYo/Rkenf6Mv/0dD
ykuMfWLDlPdYmP32in+RdAXr+AnUUSIzoPPXBu2JIvA4yn7z6+VH6Yxwe5nABvgF
1PRdVIBkNhBnA2d/huESEXlbrBls+1sAkJOXyJJEIA4O46tCzeCpSEGp85lWOMW6
muz5KwjGsVYVmxUee5vXXYU+Jvf/rvL7p0gxkmxLO28a08mLuoHW/3YDYOAHWY0j
k4mZ7ojYUzuSRzxgl/T87jSze61/BUUkxZ3F+RlJNWHsEh5FUCshsAntRer15l3a
O9hGzDKploExtL3UXwh9nwp+PdmY6qUb0cixYoaHNGaBNtcTjUQZhTCubJXq3KSW
vkfuHo36/jysW/bRPR66JvOdNq4RTTQX9h/HxH5hM2L0DuNGC9ra49n/hvO0+z7s
scRkGiszxO2YmMp9/E4rROB+PBwvWACOjPUfi57Yd4utNRNuNz717EJP3AB525Mw
dp1VPngVKSX8Vwara6607dadb4PkaxJE8SEyqsWxeFV0/KFXC58QeEW/A7j0yLOa
SAeTWmjWTzEpJKlC6+toZgeOYFfmG3GfMqF59+F8ohkBL69eFn2TL8Xn5nkZSjR6
wDJjDBmMtSWUGSV8Z9eprW0TuWhAMqNxvVA8mHEtD6TC+dCJkMA0tZfJLDILBQjD
rhZgY2Wxyap18sXghtZqrkFW4AJETz4ZbQngUrjmDpR/2WIF/cJBh+5Pmg0xQZnJ
lqLUnMqWLHzDIsaWMfHweA1/vDoT/uBPJSedquOV73Hm0SC5MRP22GnmmP9uB04k
o7GKm5KluP2w4JHPciTUifLiTZU2jUwg74fFpQ1afU2iY8o3Ng9WAmQDlGKr9+E8
/EH4DlMXlpq+6jrhGRMCChowTFcRTX65yb7BBzt+g8JNV6rCBg0x4UPkL3V73jNR
qdsYR0cDw/Hhmn82tglsCXAs+z/O3HClO06zGR1dcKvg92UIenWOe4q74NlfKhPx
RASSzpXjZlZ81t62xbt1yQ4PB2QAjg/O8GuT21rnV3ucpYz2XO8Q1pW+N6nJD0WZ
SBOkGd0trYDvyi9HN7rDcLB9yjDAF+dXzZT8p0wo1arivuiWBv4gzD0DElrsiiM5
rxkpx6F8MbYy1n8uYAYphkAatsN8M0921WhjfN0mum+AxvGs6OXCmy0AvdvE8b4X
2jLFMGXVG9MYh+XqVdngtCyj4uc+Pnc7gbcrUqoTLKDZS4h/OwLMzleqIMZP3eFg
6Jji58JmDhnAw741uU/m/xulvRJRvAGeHbnO2HAZjYCAGkp6N5xl9RgtQHA4Wyna
ibefofMBcfQYENDydOtBSnxZdpeNWCVt0DYX1FhtvvFl+3o2TmAojJny11p85g67
5kBMGeSF7Lbvgn4ZG+nidGFAP9ZmxTWSXRVeGLvIUDC/C7CQcgqMRsXdmX4Yajyy
7hDI1vZcZYJZpV0Ao3ZZMdDqNhz4uAP/lSadJkeC6X6p2yxA3s+hAu+PONVdPAIi
tpa9Ls1UTPiubRbUxR7a4Jn3FyvVWvoZLXhEQQmvL2K6K2tdk/SeH1l0MUflyoWe
BMVMCnbYO7mTdAcIPgmAm9Bdjq3FJNUU/O6z+DBOIqgtlax2C9Bnkzb9MQ2NOnw1
c9ZXq74ejWqTC9o5PXAjj7GkZZkpvb4wCYSPOm+47ztMHegRDYQHomIV8EE9qlRD
XLciVCq5VKgAOJaXbgtLamWyXO1nn1v1haGYxHO/NssL3Z5JyHq1QufQMF4dy5zr
MCEmeRqnsY7DxvPb8b940tzqrmnSEcaegYep2+MO7DFkUMlallo3sH7vpE6aWiL4
herOtYdAtlcABKFKUrZiR7VaCvc8/J0IPgHX6L+Q5X8ZmU+zP3BGprbPNqGjD/dD
1I4Ir7M5N2B5LNBEZO04aS/1pL8sxUHuj5CA6swxKpfArLD8E9TVWlkvV14Orzii
UsPtphWsRSnC7u+7vhaDbdcD47EPAe9VOfbRGJQOBGF4E3QLHMJt1Q9vV9zx+wl4
kMm7mxyluSf/kRJR6scMoCjaJo8yw5lta7nzCbb6+mLnUuAEYBirSOSzokgvOQa/
Lwmsj/ncbJVL0hruZfH70LdAWjrCrSY9U90To94CXIjxvjSbWDS2GFuVpIgQWHq/
jNrO0kOqpObV1vFZBqrPpUcdE5v6AJgkTa1a5tHTTN+uoGJCYqZGqBEFUY9rm5lB
sCtk+HEe6k5uvZp2I/CVFafLMlSZ/KJ7YzY4KHOqOFmqvzMgninLP7IJ2buTcCGe
yALv8SIzAQGVXwPKsI8dDd/YiK/WAwX+PKS7QqnAK6jlIH/DSD2X2Kt7rGFB4i1C
b5z0hWq1cU/WqIV1HmJc2RvmGUm9OEnx0iKx2B3SMrJDE8lDBaFdiobHKFMNjPhf
JJzZsYx61fx9XXoV4hNCTQbDBNyEHdkrXdBpum9/gxiRxNrk16qnkaMD/kplotNJ
0+HNUjM3FRXRoGMytiWKfEm48kU99Lwddjn1JW93yEZrCza5qmN5aQQixcgKp/j2
ScMi7SWHEyPP2gBcHY1wrIvM/CB18ZkFxeT4SKP6Eo8/WHOLJXISNk4iilKww5qp
bxFas262Kg4THTgBKvV09fHJuZS21wHz3ljUon2MzdYX3s0f2ZO8UrQgsHWBKvzA
4OOwuqsj/ZfwWxmSvIscGAMKFshVDE4tuBRApGQAi0CVqiP+YFbWK0ftiXyfwBSb
JoUs+3GplXzyZop2ibPENGsxAmcKE81JPiGc4kh0EeQd1SRpH5RlnlL757ipFpp5
hSYkB9GVA2D2K6ldOHVz79JzrJphaaOrC+2MH5dpoagX85LCBVQhcshZ5oegGxW+
3IkeCAzYjFmxbBM6mUK0uiAY/MQ5LtHJ9aVbIZ7WAvo/R6+dEkKNuDGwrj4rYSGI
8iyb89vN+fNw6Qj/ynq7stt7et3XFs5hC5PbEF0yzV9qrt3zC5QOf90HO7WA6YT1
NqAae8HEPgDBbyEhwauI2nRob7Ad8AfQTgbYRTX5ZPaXgCS77kIn1eeodrkkFmKQ
9yw2cN6AA55lqH7kpJ4nGb1Q2VbpCxxfJQGyyRhMFU+EHedlZRGd6qNe57Nw4ZMX
/u+W25kto1CMF+5oHe2h7pk8qgmg2CP55hOlVghXv7moc3EyigPKVYnhhZH8Tm7r
wLBIAY5QtKOKUyLyX3YcCbjbcTdJJAL0vVtc8cSeo5XpElxElTq9m8t8/0YGfWug
EnnXb13DVCo3XEXMoA0dBX0Ddy4aV7SgkEneeSmg7NzrGsVLeRj99jtwuufUeVaY
mwuCPyx5xTfqX9ZHtC6cL3qDbS8rEUvgu845SmE4p7qhPc3j8Mzrbt5p4jBTFsvh
yUn8BRKABcZ1/WgQ0jFzI/tl7nXp2Y+AxlSfnhsdy20uHuwGvxkdWNELpYr4Cn89
+mtzzUUXjlhBSEYzaxu3//hEVs5EfehVbmHnEzXfSmvd9v/tZbpibj5u1KObUtq0
eSkTJtlvQoVYR9zs5GcImIuGREyOrjRFcPsQPAJwJWqEac9GptgaahP2IpVeUwwI
qmEGVzhOSuY+cauaZ2WIWbW4cMhxfMTlTUQduShZAigM2AomvWdYqd0gN/NFeXx1
TtKYPl7D0ObYkdwly8aKBryblycLWywXPUvz93XXepor9KxImhMaOj+5LEfexDSQ
vRz3KMyHA6OzwbUNvpdue+5WyQk5j++6izX9hxYpIa/inRJNWzl7qI7E4t1C+K0r
jCuaYmy88b3pX3XavOu5Xh0/tTD4VnLnCRfy+kDdJpd9pEaegRM7ztz65gC7+XrV
O1j/11IshboIIKOYlpz7Se8RNZSXSjVemLk7l3G/sKwBQv1qdLKCMrmD5/o3CZYY
oIkw0W36c9JLqkIA89xnkMEcimcb++2omzU8J1fIyGKCioOhvM253W92NMNglArf
To4G7Mdo9bNP9tYyotTbOpGvvjIAL+GWjKMbhS62ueA0PCuiQmg6GI1zfGUfPgsK
6md6whAxtnj90zB+R18KLp9lhzNYLuq05ejHqAykuC0owmEc2RWgG9QkFPQJACQ3
ixBFVQvo6teBOC9i6fz75Ty1x0xI50N1IaZ9D7xPqmw4+1ELjSBRUoeQiSMCsBRD
Si9lxN6S4ZYxOffizOGE96Yzyw782tz8tM+1HrarG0vnaV4HgLw+/ITdvyOCXeDU
iAFjsfkdzrTfadzoMztj/jWAVpe1gATkv3/1zmPOmkxy64vRsn9+YEVBvhiRGdZ9
VcSOe/X7NRuu9O9zGYE67+KcMKfESFYM0tBAQY5mq/0NmS5r15zq+1yESghKtDBR
ZM5EizgMsQQqZVtFaV+SRBGXFiaGSvxQFcXEEgOGFaevsUBiFSQItGCl3cwnuwAJ
APZuZ0QNdXZd2AdWF7jdiyTJ0QdOvOCMzywBnXCdeb0TQIKEWCiT6AN8Z2SNYJQH
hvmK3cvsWbPMsS5bV9MkZo3qxWcfXNt50kn7ck4939dyWEbriQn306LOHPaV3vxG
f/a2gQk0iXzMYiyocN7QtQfrexQTrwnCGab2I3Y2H9Ve+tSloh/6OjmCZT7jCEk0
EVk3ma8cAmKOuTyOthKPah2NiPK+XjipDIdqcl/AjMGXTzjrOdgAt/Vwfcohc44V
w1/SMR9Osf7EkmvmmoK7a29Mx/msKZC2szbgZ4mkjJNN1BHYleIjBYxTvjrs0X3G
tT7s7vDG5k18s/0yr0PZ9IesCJrFsEud+ngOi6QqgAzoB0tfHL13QLR+OaNV7zil
Se3lk41wcroc2TRwrfePiO/2mM2FnsYCODYYBRmi6ZLv0g4Fua7qAluaZzzx2LeZ
PMeuQKhu8/qE/6eH/cRaLvkbpQJQxLV+bFLXln6NJyz8oiS3h+kogQg21AWLqAI9
leuj9FM0/TPCCdPCC6xT5N1uDmdTxVja6v48EFunrbq9nFNyjjIY1arj+D/31bc1
Fdz9HSsO9ndTfhcLson5odaSPTCxwRKPtbbIKUPrI1ocrj18KOfDev2y3dOoBeik
SSoSTQZYjYVRTxtHJ1cTg8+FWb/O+SUVVnIcU/q22GTqyAYEaiYS/p69V2ixd2yV
1C08idwXkY+FTPp7PKsAFIsQrgOUUftVZUVHK+cM34Bx+hqzeiirpkI6+dl9GHNk
vQhm5zks2jY46m4vwXYaNoeU3fJ6Rufip/lyNCRFH4eaUl/HbCR74yLQNKEWMElM
ThFmDRWEPrPWfcFnGLIKAb9jCGC2E0l4FFbhNtXbX92FQA0Q5xyn5TyhRXYYjVLh
QhQJMVqanoXspsDX5+FzS1cQ0/roO88KnUjhLQ5E2LlRKbSHda1hVM5c95YoJjYr
Zogv6mhYQ2+2TN9m0Jc7kbpIve4WSq+Y4iSM3T2gaf6gqOsReL3Wh3U2Lk+Vo4oj
bU7b3qxExa0f2lami522uCHkWk8uVwZJ9Qs5Q/YhRkXVt92WSUD5RsCIrOJOLF5V
Aj1mB3QNdbfUc8FxpcZ/nH8CuCszpbNFeNHVFoluxMVruBB4pRzT5XCTC3rAsQaj
hUXZJl+FbPk4ue6/ZrCjtC75Ro02ZHuZzGVn1aPA/TMn40uIDhMcryzma8QDZnOG
D4XlozKlXbhsYvFjrXLGfgaQGlOreT+jvGV2J4+pM1KuW16IJggKPdBetLHfSGeW
8usHr/QLnHgaQfSu2VK6sAQrVuynoReFXFWEt4a3UxQKAow4t69yZRTHLdjSKET/
ztOfwgQRRBNy3cKgKj8253Q22CGo6BKGo6SNwfnxxn3ro8SquZaPMvCBlRyQK0Ny
Kpmk5nYig9UZ1wC/liSsr6uv7IyeiHihVqI8PMIz/kpinpZCFP8HuXsiPRUHQ/8h
8aOXRyOF6qUxI3K2SKbpONTTNh5dhAwnDE9U/Ry1dY453CwkzUYhp6UYad43WOin
ThNtDoIj4Jyk0ImjGYZM12cuWiwlphLmJBKNu5zivb85FpTLcU5dWYG6vWgHZ499
huKOB0Vm3y5bOHM0iifY5PsgDt8/9EqneTh6tEYy7e7qCxGia//Hao8czf6XvlJT
z+5IeUPywR3qahS2pcRtgpb2uX0Az11SDVzkRQC6lnmBXsfUfBKNegVbuvq/trUq
Vx91AN8XBh4cVnwG1y+Na7YFphaCRL9ql53sQalcnY70L21+xj9O1j1/Ez69akvZ
JWe9Gd/f0twmU3XyWjrdzUMpP/p+WciS0IyLCZLaNCnZeRqy7QiPbMvJi7h7prXl
forMH7uP0yeal+PGRwhcrQU6p8oWtpx7Piqzb+rOP5BT3wHfIKKTVlflfW+1E9Lt
9HnTlXulpZzgTQKFIqITF0B2OWkeBnj2pvm8QXzSKVMfV/eWJP6oHUEmZ26TvTCU
6V3HpmXlFVu7WwY8jReMmOMUlaAJ5r2lISFTcBrzflDEbImy+MVCzkXGFjAo6r5c
3tgsktC1LAD4ubc+LA8EEzG6Np8FMKiUxood+FiFHVDU9GXB80QiuiWiOyTr4LT4
jMee+NsAX1/XWWFSY6hw/b5SWVHubDZ2Bnwi/yDPVRiWNp157DIomNLrzkRK4e3m
zygkuZibuWdR7fo0zK1HuUQnkeFBi3Dlwt7UI5KHmAxREY7CcChomJqElXbVxUSr
e/ZPi3TvSBUNOWq6ZqNYgrAe5YPgHuU7Zv00T9nYqm+jky6jtYgsu0A1t6NtmVrr
XcnJk9EZMNxXpQFgY1m6jNyWurEVXwjY+HPXfz2K990CEzqtYdEEoRSE5h4SgWmB
F/2Rkrxf4/19ZX2sY8lW/Y6kxEyuIG+bQi7CtnRQT2sn4puIoVtLJo3PDjTNwRDS
cvyCkS6jruZig8dx3NLQ8LiyIIzgkHl5sfW5Brfk+J58VgzswO3/YlNRadQHkFEP
yKDJ40WCOVcoAby1wPBY7xYK3D/EqQ+Xr1YuVkgBfQowgmLrvJmpRO5BlPCxOV8a
sIB8Hm4UIIjBN88AaXn0KEWdYMJ8HwUYBxCHobn6I2Xqzfb5yjbqsRGmuLHxgm1L
M8rIiuRmIyiApVNesctLo6Lc/FONZ3mAekxCtxHpHp/rSV0n7sP0opcxcWHAKGF4
c1l8qbCeFGknkPcmi/S7xwaszTTQ0W/WK3aShPlkmadlVMaSubWVK0662NvMSzPL
mKhLfKPsbMAogR2NkJzapfZ7LnV3uIPKWq2EKNHdQf4AzaylkMejD9+qkbX9AGf3
Syfln3uRsJ7A9vEPz58cd2gV5nkD20QMkgYmxDa5h12xkQd6qG1GvS9l9W+bN4Lx
49YM29vyiBT35n9QkBOf6tWMlvOWBTcMbrW9ALlU19vg3suOpHafB7aYLzeSLaZ+
G7nbs4Yt5aJ2jGvvOj7Ph+hz8zIoOy6TIuGLA020/q5oeb7KbSFA2k0vZrPr0tkw
tPlfVeoee4kQ08T5Lh+7WM0TfXRm8j08WKN8CtT7oPJJ+1JI6kpLkh9AGw2HSlPK
/mZwsE2ouUavx44HcF0wYg+yINOhQLuCh7sakU0i4XQpJwKJQMJQVNXfpvujFKX4
scHNwq1xjlBdX9nMQZh1w9zdAJd2CWRBT20p3bNQvDiV7KEifWUKiGAcpLH6XT9k
Fa3hsK2hPvjiHaBlF9JVYqf4JzrN5ZPVBdhp0mFejgAJal/1TSCvOQ4M3XR6RAkn
BIRX0F2mI4jp1GRyOCKkEMAB2dZGHcXAc4NkpAcbrchMQXORnssmDRW36vUtFXBm
/JdR8kGEFNUrRdvawDFuw2Lv2pRb8m9ilhPgGANHKQHGzAfBM9AHOVXDruft3aAp
V+ECapwLnAkbhjJJAaFA/mQZS7EM67K2r8RasGKIz4qeGtJR7UZSArQCidzu47mn
Kot9FTeBwjEehoaONjmlZU9dJXa277CN5jQp8jSCx1HQJGgX0C9m736/g2MioVOp
wCwQe1hhis4/0n8MibuVeMK6zVbdSuUVgKyEed7YtIxbC4kztXv1Ypa6W94TrBj/
AZPL+VRMyJ2om0lHTcNs+WglgEa0CsX3cxKp/HVoiojWOrQ7RWeCVzdcpVftDA5j
2bz+k/4hLM9V8XOtrkQFdPBB+SE+jjbOZGL1QHLuK0l6MA5ypY1O55q8YEEliri8
Qq5O1b5jf2B///ovSprOpleC5aXXZN6Kx1r4gq8S43ZJD6qVrgPaL7exAzRVg/Hd
qhi/M2qS2LJgUnIAXpPjdgKO9f9VHcICwx34afaQeoBGAJprWWiJo1jo++QfhfvO
ST4D3p3+izh/iZXBixgt+OQhyu7+6QeYqzSwPfJvAZsAIKQye3qPisSHa27lfznU
u9A1+M0TO+Czk4VHJsmodLwv3eAs3XCSs7vnzpgQK6gXq8uKYMhjCaenyyDFJSY8
8qKNa0AuJju7RbbkIZuYepTQ+yq4twOiD1DuqOiEFm8id+7BEDUaXOBIH1JOMpuT
WxOelPOSSvGfbQnQOaWCCEY2dWxacFCYNE3y9pSCjFzNS27DqVGPs3wjbXd/1Scb
Os8Mp2tvKDFpyqltuQcdrMh2f4KMeeZXFHzhPpagnlQIpx5FcC7lsHPOmc/aH2VZ
lNpcFXSEytD9oOp/KwrUXzY7YIUh5BRt7cvWQGh8qhne5Lx1u8l9ABg0q5jA6eqo
U0gJeH6aUBYC/+5B53nvxfbgi3feFR/Vl+9LCcwA8pgQjXMpsimcZCzTXQ9EFUvN
rYtDdFQRy+u2YfrIzq+6SMqmNVcuQeo4NbzkbcTckW8SRCjTomkUmFP6Lm5r8djM
HZpNFjLxmAYfYlPHnf4xlRDvlbFPp/rsG8TtxIx8f4KyueCicQUu9WX4ztC9gQuH
lwCD8LKcszuPUak+RFv4KB3Z5OKmuK3yLzFFLQw6qLG3eTzNTOFeUGGy0MfgcaSu
bAsAnszQDvc8EjMYPp10UvzMMymBWwrx+/uPItXKy8CMIVBbsmzEbLkXncDCmGOj
4tQzlymWSkgVvY4bqAYfWRl/yVvRnn72cH/4FMCEFEJ5nkSMQbA0HTL0z6M1bnmo
Y9Gz1sZQpr7u/n4UlEuFiGQ906BS7hvA7aaYh1S43JxMfiioMmTiwrwber60ViVv
IoEQRTAQO31qn0sbC8aDvkyKIVK6/pffhWZjSg2I1JZrc7bx4CNWP+zh/HOWAjhl
wJaTrxPHqH9cu92M/obICvh8pTlGvOwsxySp6SydWdpbi1HcHzRamjxrikl/tD9g
JxqyMvcXGsDT1JiBJmyWpGFMWJPHg66x+TI41IYSM27RA1Hhxu20MQxA0z8XW/gF
KjQ5o+UNAB6DtquyLDeTCQMyMR2Jn4NelnlMNBTmiJZwuTHcKE5ce/PKhm/0otcJ
++SRV2+fT1dg3JZFfXMzmHvhTa5GaErlElfGUzqaJe8wH277AqwMWmkajfSqwF9l
P4ImMTjiwyHM6f6RQd9zAUQCgWVvpNRYdDnwG5fc0G0P5lfgk4lE4OIZyrQKXCO+
de0BKcNxKMPLJ96OAig/65vtsvhW9FIxwOfagwrFv2N6mVrduDToXG5PCA4uYx4c
MSWqZHtbADPKY0tagXcv6Yfrg1LvZyRsCu+gWoCNva35atRE7nXDEw+z7EElc6ml
XX48JztOKVE5SzQ3ga7kV1yd4lTOgJU7vYAEQkNXWLK+/V4pUReRS+OJhpm60SKI
LAIZf4BAujr0uKUsZVkypuBGXjUUCKRZn9QSAk1O0TvSV4HjP2g3xEvvkaeUHmdy
CbSCiZDCdlShRLnBIZJutW4Bskof1Pz6yqry4H+iZHf+OFfHfJruIdOaXP01n94P
IgUdbjksggN+np8BkboWzgnRbZEMef7VfK9LlnwTK32uZtBN1pH/vRkM7FnXC74G
DVSbJq7jFn4E/FP7zEpJbvIFKiHHlzPSe38Y1b3FhUlvd4QAXO26EKPoKZZUPek1
sm3ey36jFQEEMqHPU7oA4pPiwVrH4j3Ck0ku2AeivmkvxZglL6lX1ngYL3GAEGOX
cbupyst7x/jKBKPBO4+Skkd8X8kFMnboQCf7d884zQniZt+PUkkxQw9mRdRzQgKf
vFXTdMFv20OaBVZPCvYlgjTxzD+SaPw/0XCHeAXE47tD19QS0XVNZ5ZJ8xP5nExx
i7kUMEEZBeoj8CWexTDLSFX3fQx0gv3Ielk2wF7+QnkezDIXN8+OQX15oFIunNVE
IWmZFbKsswOhUHAXT5aXUyMbFdSAR88Lu5Rtz4IBRbR+LxxeGoGJ7flFeHN6bRP1
TXZG7dRmaLCew6mVrJ3XBve51mDoaKkoebIkmj4i51FJafwm2VDCzug23Edx7647
FshhjXkyvSL3nfbvdSSHNueNXlJWn3U0SJYQicz5lQwGuE6xPBfwZ55lgGC2mMUv
EjhWpMhDo4X6q8ax1xSKpn2VGzsmnuflPT5cUqwgNRiTGGjoOTo9E4g0HL0vl/qa
PL+afHTlVbh708zFigaxtod+8bgRRDPsAoIx3s3HaXwOfKQ83cKPGqJ1b7LdyP3B
e2NCqiVJbznoENh9GCMBd2iw5TvgIXE7/MaGuWt8QLo52u+GTzQMXQqoyay2orTE
mQoJemmQFzM/dMyfbq0L/aT246fz6dU49xQ8WWnJyGyZLCByW1CE47XF4Z8IbDmZ
o58jwkOvi/ELTaeZ7yUWKpWbXXhY+lOtMubfZUC0aOCEbxD4Y2GFeXTt8k5DiQ/r
4Cead3JGCPmmMgRLNUv0vzDkcTk6iIn6cNryUa9t3ZD9McYjVJ0yTi+AagfaQO4n
Ct/A3GYu9AAb3SdBcIbafm//eRRGUYpUHABACmJnZ8I187cWPp45irdQkVKyhTHl
FEWAQ6bEMvWBiGDTZHMCHjhz903uxeaRg2ZaoHMHLwYxlSDL6oqGWNnk8GIzpOtb
SyJzAGrM042rRi5aA9jXTm97eEXVfeXzFXJVpEMjCTB9MqjyTvkK3kNJ6jhpKGfs
BMGeRwPt62XYNQTDZnB9okA19/Eukxp3BtqJEzbkUNlh3MJoVpRCOUjwA5AfnDtA
4RHsH93N69dTYkCK5cK1yTVLtndgNx1GCnViEyPf4dHHZaDUxsCYhY4RdpROniEY
M6GUBnr/BJvk386cbAg83mSb4wxIJXGPgzSH6tw+EuBrxANGytNo+2IDI2n2a1GJ
FGDtJWPkq5Ubi4G4ktCQkf7RFDtMpITCyZZdeANnCzkBczqEwQJsOiU01NpUrqi/
2DV4708Al7+15x+SI+dCGQ1QDYBEQ+JLW3ufRcjohOPZqH1zlaOGmfmPm2B7DtV4
IvW260E692V76pB5Z9nXsySFqyamYViN+7GD1B5BrTxbhYJrT+DClbyomRxqXeUt
LU0NbJqjs8jQOvQvePyErz0o/oVJUD7IzTqPB1bfOyR71UObQY1h++jBIU2RMaUG
8Qf7agEwZufDO0A+SSQhArsGjLyAkEsPPbVYZkrwwvEW5pxWZrhRcKDadoH0Z6He
an5yZUmBGbca4hGcGOKX1DS9oZ+a61e8IbcQ7hgXhvawUkoyXjb6YULlufSV6N/Q
24Sd0jGgxiDNhF2MrxCJlUDPWSPYMs4JK4A9GZ/1yBWgPsSKVURCuDQX4GXLm+qT
27/CLQ9IxXX2HtqCtbx31KM1wHhDchZGLrGgvBbAVA64UA7R47z+o+Co2u+VhEHq
dbrGZcu4BW8OuWzW3wQXb1CE1E5IfwB/oh6TZO9/V/atfN9LyMXqyJwssA7qIOUs
xGoYl8imgibxto99+66jhJzT18NIfQsYAj2TOH91aKQxlPhqmJlIjdbiyZjE+Hh8
Te6sW/dKWbPVw8Y0jXyjhHsNOtoGfKv6XgoPDdIcKxhmTl3owf/TLSo6qti9Iedw
O8VZbohlv5ZdaSMPlcHzd1HbHsGAgUgDk2Wo5dHytpRT3OHP6N2byRCmng1PBHhS
3mdeGM9wPb8ZWSROnETHfx/8thwZrd+S7+mJIr+rOz4DAXXf7FK3psDGTlXBlum2
xWJOq8PCsbHobi9EYlr5mVj/2sa/jNxhc/d0awtX2juWD8NUO/obFsJO3DuUi3ZE
qPZgnghFaDoMc3kBcaC6/Q0UxvXwhsnNMA+9aW70Y6+Q3bBt0y4FBdCcnVZYO4oC
AfPjz9JS8KLlz7W2LqFqUeRkeNG68aXYbgrpTn1Bn7CRtGM/rTpS7c3PGGsDXZKx
69q7NNfHNRFCiffThki6WdpjU5aGbZVp9blmqdG1Ue3kD5fQFc3T0CE9rIw3cw3Q
HNnt65zYrbFab5eqvhJH00KqbpcHJUEfJeO/JqZ6nVA1gZDAoHiM/fG97Bbx2q+a
uc3uHdRjUYEGWhAwmWUcZCuF1SUXHFiQoslOSS+/c5EvSQ55gwHQ+w8wGSPDtahV
leF/XY369I6rWzMFWTia0sPBonUWD6P/bZFCIMAM49h9meVbcytYjOKQSoV6kyrM
7yaiYp5QvPWhzOOCCJMm5Ytwdr0vKebxbfoy9+tPTOq77a/UPlzlGL3UirDVdCc/
THZFAW+89Mi56dZA/5EU6fSPfEU4apvcpnFtpN0rv6ymtKl1OcwNIKEDbLVL6/id
ga+48/FfED+vtmI48WRn2w8oDFPMSuWkh3xIBDGcFmL6Ag7Zw4KqcUl1Z6DKqowh
YfPcy6BrXGkThVziV1o78fCpEOllNj/t/iJacB0OcGIVhkV1Sd69uevxQ7j9bOuf
ftWzXNcHZP4PPXoxtsXKr1elYZZ8VzxXAxgDVIb7GO9JX4Nu9Qa9yOQHnoHntrPS
ZqQlXIwzj5vY9ORhBCrSF2G3/x58sDOLjlr3hNNqu2kIFI5n/PJC7OmTUvyaZRlh
H2p4YBOtN6vVzwy6y07mSKvGsBn3rL96q5gmUWzwBAdsfZmsBIfDITbHMGRthEb3
TThwqocVuSAA2n3T3TCFgG877iseFoX6wpWaFct2/RVqRgjK5C1vofuMfNbhsmZ0
IbCy1P60+neAoUjvpW63MN173EaVJ4H9yBDJVxotVqHdUmxPG2XdzVeDM9QxA8rB
rgOhCbHHDXpQ43uQpeRXsyj0i/J21Tu0cIABEKSvdUByRKlxjCuc5pjTpHIBHvjo
XTlltqBK1asI5llLZdq2VJ3MYi4wWav9g7a5ke3kIT/YAejaf7jt4xYYgaTiKxmp
08NEHkDJbyyar2/Xq/KHZawFGsa9JxUwmhArcChm199CsLh8eqJ4s954xVAmk0Pa
W4u4bG6UeswyDjQxSaEa0qZKb2t1O1L4wtTCrJmHvXTTSWBYGR70KnmNcyGIl8pE
`protect end_protected