`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2992 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
2n+M/KhW/CoPvt8soGKLVvPxiuvBMvQY4p6CW207NGGHimpWqg+LjuukwhvBiJkf
juDlTOabsps5YiyLeU8unOu8fOWahdE52AslfwO8ljumUARiqTVQjLrhdyQNfzyE
yRTlRf4ynP3wwr+AGQU9hoZxtRPmHsgReNLg6gGii9FizH/RMCzLTQj6dyvpGv6s
GsjtbOGd6OHhU78mCMvdeC3chYi0RB4Jd6vQpuMFOyTtS2mE3sdiQYf2zFrN6Cij
DpD/pyI+kwm2jLWcagATSdEZqq771ChVXMIEmPXYyWD1dT4w+ZygRw1k2GwmA8JA
g5dTuZljEoZ6P1AyYEpyJYy9el/8kDhaRM/NYrmys208ltcmFX6iHwCj1+FV7BiK
Zc0sYn8beMr7qQzI4JhUl27fP+mMfcFHI96Q6TO26wfVnfBCCRErUuMS2yX9tZbc
GGG/u9r/SJe7OSzsaY8fh4uOVxTrM4kzqxrDbo907TW6Md+qBaZlFejJjRcp4HmZ
+A1uATbvmq8TnllYMhLPYgZMUAJEGQO9yC/xGoTHdeSvzHCdxLasO3X/oAXwD8is
sNpTiKORwtSyywA3KTpl4vOLXGX+gTxY4iYffBHJ3X4Bv0ErYx5S34FxrMUXPvjt
dk23hytHFVwl41TpZFOVboO3mcpIeMhSlfFo3qLyacsNeOoRcEp8lWLu1hc5VWE1
sWivS7+C+XwGDEtzMXUuzhIlqq8beC5RQZcaBsfFSKK5GIXkPZl63PXLTRhWKin/
Y//Rbma0gAuZV6plRmc/MXE/parLPjUllkpRtx943Es/OHh/LhG6ch7y2fxkgn9g
Q33j4kcdHC/JW9VmVqfXKjE8I6c5XRT4ESWTUYE7+P2E/KXDz6JBgz68rPP8HKGf
p5yQS/Id6GeBaRSgtqC/oXMwGhW73CW/qsj9GL0zI2RdZ19hX5DNYG/mTZE4osWB
Bv0L+rsAPJDpm8Aa3TQ6Jzc+R4bLNsDBsn23ncm1KxAid3ISP2VDdFM35TyZKt0p
jOFwS3cXJJWZ5CIOEFdXlBmN9zg+K2rBzxk4Dfgq3Pp1sDvCZcL9LjNhTYx+048S
vv0twefhOddEl0/8qFwUxDMCNeGdh2QaMeS2zbcJJYT/Nqr3Hq0oEtwMLAQxS6SY
C9byIExzxMS68qAlIKFksLCqqy/088tqVuzMiFG0txggnV8LY6f/yZN+fxSrzaZj
n29xx6uwmF0toZX2g4APlI1hZr+PcfapQALJCV+bS8jm/dCdPEL6Wpw3XlNnIUXV
N6Jfr9MxGi/Lmeuy/Eu8rYAvr3rkXBKpZYpJeMUZb0KfIjLuewnq/1akxy5ZuZn4
lslSFGIUj+omhjRY2J56CM/+bWxn+9eDcX3G3dRG242u3VkgnhzUEzXQqpQYCnGA
0uV3CxdGMiLrU/eYYidx3AVamGjoVehR1dB5cqA0ctEweGkOIP9zMng0fxmoCmW7
HofrQ3+BIyQuvq7rrogtujnIHiRBY9VZ3Wx1EDXd6c46W22NQBdvvTOC8Pgz5hlD
VNk43EBcUrRovadlrwPxS3awpNRMZF7y/ICgwyyedLY/1IHbplJDjqiBd20Muznb
ffWI/IRVV/Qd8hvKLVXX+GU9yVPOEqMvBl/t1uqpIszM+0ewGsI7imjUSU7lvJme
F+gEgZXSAb9tGQMvJEz7E5RZpQXhzg13ozsLZDInRyzsCrUH3XjH8xDlkLEY+kTL
97qH3RRIVoq2IzZ1CpXF5faBvojqvPv0Wvg174F2LBilix6+KzzOTg6YCgoXWG/M
s9dOZpja/Mvc8HdhrkgrgbJDxD0gu8eE3t4GZOylTSSA7tHDSbP8eIfYOpyv8wFi
WH/UhBUasEW3hoC8eK88IYAJ6HX7gU6nLobuYunMrxx5/eG4xYbX2By/qfO4UZS/
f2bcxXwmKA0OXeKoHt7xoPB7fqfyuufZy7dldO9X+mh6YDBDW/RBQvO3F5TKaVeg
n4qYvED52Azh71Wza4NIPz0qILNHW0BReTez3TTxa/7qU16FlnH4bFC+IaTi2x2r
yZh+N/U0ix/StUEYpocn15lNP7ty7ySrrX/rwjYoltnv6dSmAbpGNCFdzpVDWx2E
zrrPe4EQ8U/s6/axNrGlPgKc2fR+wZSpML//uEKWZ27n7lP5G+a/DGyiZSEGihR9
ug+gUEvDZqrCA6a2kWrGD7/UFKwQ8Inux0U5Mfc4l74dxuUELxZ7Snr9bgQ9nZ18
Tw0X0GRNlJ1WPQqlZzH9x/cXRIuamR0SEo+w5UUhEmPNDxQfMNa88VFfz4Bh8nAE
W8tTC3ToCvHQwSY1mQSb+rj9bXSygevNiSEscIGIVoQa36q9VPhTCEHLMJgdgUA6
Lvp/vAcAgVAg+7A3wG8qOQIKBg3oM8wp12r2jEXIbejgx2LXRP/XCG6Q/YcdQgNk
Tv3+XjQBhssVw7NV5UGNrlhWkQO02tzjKWNm0mzJ2BIgn9BJgo52xSIr6Qpv9WRn
HZnRgrcbFvzCTuw9gcLrVssSzoOwm5TXVS3jMvBdB6l1Hj3ncMRCmuMuTd3QJddY
qpHv1viMfXiirihcWLOP9xNUQWTHBtbJJYgfHIuVb1gRz7iq69KopKQSv2LBiTB2
xkULQDNdATDaV9YDTM5DN0lano9aLBCa1wS8IiwiPAwiZmnn1MIPyIluur7L6Jex
l6HnaD83sNigJmiOtJGGXIdlT9BES2mBCZlG+J/z00h6TJeDx/tbhneV6TqceH8p
5mmYCl0SPDKl0gX0SBygB3/Zw8+KZLPZPqAkuihZiiLRBTfVMMnIJJmHd64Nvg7W
so3G/0LixX8oq1jd9/AQpF6GvwSp3f4i3rtGEJdUkvYKGEKVCpmWuNWWYeKOrMVU
sEeluH/rzQHiQwjn9mpFFAufdgXMR6JEqdzSkIUm7by7evDMpmGUVKTIVictmi+F
dgycMOEr2FAdjIeAAqDbxtgDLcddX0r+EvFlXxdxopGyywG5aWfp2p9GdgREwqiu
SVpYFjiefGEofNEGBavAsryDzT/E7EAR8vYapcpb8DYkEv5a9OIOO8AHE1xfYwID
nHRHcR0iaoyWCiZeLo1Ad1XR2vykyMlBvYfqmJCh3zUDkuhoNWOUPtrnxzYifsot
35is2evZHdwqX2GmIOfJgHejswhZ9gp34Mk3FrBah40k4EMVD5H+9MpRYPHUnKT4
vL6NxiTIwWmAOH3zWNTXfqwpXgRrmXOoeWwV192XGp1GM0ae8C+BPgReYkUkGkbf
3oo9OZHcrRTzHQeUgh/wAaUhQd6uwNsLPCEIcJtHDNIepG6I1wxyyTHQOwy5hOLt
lN8KEMREx7T6NI2ovWNjcMqfT/rYnrw2lRpNtNYiJzjvO4mc5Dhbp8VJLIMQA18M
tBIpLk1wx56rcvELy/u1p6LvNgWj/iCPFs9osxdTlFqq+Kph325FF/QQhRNI+8PD
OdEJBjFAkSgg44gBP3FSvXaI5bgx0QGWMx1DpDsVBuR8n+F+zENpkEZsM0fJD8oV
n2fZHop4Oba0RoFJvazlQC8N9QjTJ9j/RYKC5AoxH9AA4wjAgCamjjo13vt/vIIW
8TtN7A8s7sx9sRUShgJUagcbLN1cSMVqdjDaYefAecgAg6bwDtvh62ErXyAw86Hg
Pf++NusAenKMESHYm2rCewk8TmnosdQ1NdIulPML7mayG3ig8YZSszux2CCyIHHF
OlVnhtJm1dpnQXi9H40wp5Vypz6wxIeXV0rsKSp5GNI5kdaUeiKGqXvw8Di/2nSB
gCz8MC7BomhLpGpWhfgGVFikRBZ1gpTdxugCvs2XaDQC96lo8lrBJApAN0iDly1H
gewg5sdSvFQY76XqClagkw==
`protect end_protected