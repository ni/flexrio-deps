`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6656 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
sD5jeIt/NS2+ECTgxO9JluMuufYAgWfmumrUMOoySDmwJHU8OjrXB5ZY8nXXCdF6
P+G9nB9uU9SgWTFAuzd8rTHqmZrdRIJHKFJWgnrjpGEwSPT7UeMcEh+iQhlrliIS
QsLEfbEmuzDBduk5yJiNYY4CtwgQIxilQm4Xqn0dmtd+lp0liBLqInw3N3fsMLee
Ls5cW4qhIZO6DBr3+hJwMrVHMPXGapVCs+6H2X/lRIcAM45Lnc3DSyGhBZfBGQO+
hK/AGhHr0+VoKm5w0NM7FILoGllnFZ6WlWFnJwxwmeMl5XpJMwmOnO+Nm7cQVEa3
0EwLuSwsLxBepvjQOkpKUmHxxFQ4OiC+35052SxVDnk0HdIYZ9vb7Ao+QODmgEFR
0Rjcuv8LXaZgezeHx86LlDFJT1UaKOetiv4T4zPAWwsgeqgldee+alx7tBfAeTA6
wFBck2vCYf41731yVK2aJaE5MdbY9oXZiZ6rJezvek82W+IX6Tl7lW45pY8V22lH
inDoH4v/VxXhv96A1BatKfqabOCAiyPMLgfotV/f0v3E7xZ/cli94qVA6fe8bKWx
q8D1+DR5wxEPzvO/apuPL//l9RsUNqyO9smfCz8DkylmPyQCGhcvi78gekx4UgJR
CS4HcGEhtU1l8klw9miwxEhPBu/IJZcKNLFyXzvYQfsQKb9JptmzCOX+iYUWXU2q
OBBGe6piX3VpONL0Kcm5zV3JSZZay/UW/JihMepFw4JtSKGWbkHnsAbOXRil54Ee
SAfvFlWAuZNLra70zNewQOCQviSb10UOYqgYNAHqkTm73y68Mskw/Kyv/mdH3cqg
t5aaPz7DSxBXcs98+bgxhUwSYkn8s3AzBOpTe4C85bwTMVlBsIH9EvBAJkwlwD81
0sI1BlOP5VATCHqwVk8f/DVFhSAEjpZg7BnEupCDjLsHCXKI1IoGaaNfljjMCMdl
397gf8HhUNxhXwIsSYCNNlsUMqYdgT3l2AcvFibTaoAUJ1P64gju5yEcoeZes4oj
oMg/T6rQ3JvHjb/8p3pdKJ25Rl6aO/nGb0WB/YNQ1DfitYbkAqs2TEJ918eNDNWw
6MgJkRkBD2Rkko4AQYBZwW1K1RfEOAJ1sVc2cz9fr6VriIFXjl9bhouVYKQyWJwt
M31GoPGcoMe4IvfbyA1AOqd6MOJjF+33fhzz+JyUmueEp1yAygQoiqrzPb7WjUL7
iIhh5Gcn5BqP53KkNvGMqmVqUBQx4kYcKWTCBXonmQ+CfvCMRs7ULqqXv2Sz2D4B
ZMBEPYshZZgAMscKUzx/a+UnG7+Y0f7u8A389OIAXLZaQIOi4+Gon7U9bHyNvE3O
mUN38NRVpXTklJh3tV70lfuF1f8eOy6LoAVwBuNEONsd2HrvzqJNiClHm9pnZlQZ
MwF/VoawY62P9iUTYpC/R285FvA5BxYrEkLWs6lNXG/Q6I74L3DKo14xzvvxUFm4
GsKUdlkp/7Z4Bls91yJBvzlNHZUbc+gyE2XwRSPk1N7m4+LdvEUr/8if3FIFgOY/
WTg5hQ4Xcvz1/UeXU4beh1V8tu2z2xlvhFMS8/YS2SoNipVPvfuss9eSlXnGoLDf
SIQb8XBTSG5JR0qz0AUVTSWcS4toqM/HGtSTXXmI8wYiH4NfYN1nORVpMNtYEsiq
8I0eUJh3qKrRpWjUSxAsGDSaCjCh3WN0fgtVHDIKLTwCIXgoUlJ3z3tEbjZh92v0
H8ORjC6AwfPTyjFaUZjsSp/EqDypXe/21guODe36oG/QMvP+RzoSOXYQtvJsgkO8
o97tH7at4i/d1KqNDVEzF+wGYwB95rgOnU8fJIqsGlEUWQT5QrYg0u7lTo3IN9/W
1BuNdziSkyJTxQVu+Kj6I9g+gG0kQiHRsNScF0W2DD9/ivrrwrY0m/0KIyRe7Iqq
75hlpxZF/d6juVISzbDhwN6Xv+v/YpjCqeZb+YcxmAcZ/1uikJm5wZ/Oju7RuWOV
ZDDEf2Kp5JlzlEruCsYmZQMC073WcoBDDIWHmww3rAnrbWhd7DmdLm4LyBC+d4h5
xUvk/gMZru8Cu2n75vkoTvLXWs6hmQ0IRz7nLJexREw7L3jAxWEVKYz85YEmBspF
naQKOHoMFRyw4qVfrXeolAqW0xnqpzqzTAEsqhhka+hthpGmw9oKGGbqJJcGE2Rk
/b6YNbnDQLepwFigbjXd6YU6wdXwqcxVyWoGwQHYTmYxvWvAhrfK1+qUe6h7yt5h
OqAtQKVusxdlSYtSgZmUpTj/kAnvZmtXNBB+yDD1txUxrwYFe19/Jb9Klabccrny
tunVvP+LJAzntzLvf9OptFlWA3tdFw5SyFXd9qMI/Io7f5vTEURlh5HjkhT0yvmX
IHQJzStjnakoMYrIgR8Bmq2vU7R9G3K55rYct89xc1d8qxAoZzdr7ZNURZASseoo
HOXK91wPsdlgfWxZY63Kgflf4LZ1VlCaFfwPQFpq3yTQhq9955BabCPOz6MedcYx
yX6/fPKd952Y8p50wHsqYpCrmO0CckYUvvOu8iVJK/ufw2p/HTUtMfUe2wIw8O/+
IxG+EuSPjXf1hietsHB6H0mA7NuTzWW7rVraMD6zDflrKAqRj8Wlf9ycLP8PT/9r
Yvierm/YYWfOUNEmXzgaSSACaj/OvUwih7MTxhwcAnpx6i1xUwFxQvMrG7hDBDVY
ae86+bWZJ4ryaynpP9BQfSeKr9RfxCnA4qB5NcLITjhCTG61DkpukPKzmTWMNg5b
jCA0regNX/I1J7Ul0cBjR5TBg6sGMiw0CBLV+qD648j5xdLJEi+JacQS5sdQLbAn
o4WGVu6R5QOYDg3YIRF5mPhd00XXnARIL4leT7RkuJuCet1KjZha0DOlf9DmuXAi
DnzfevZxHxto/H5cuXvzUoKU0+NULTRlF4QOb6U5xcgr8w5AxLpu9jsoBxE1YmTE
IPSTQyLu+vokLmTm4uwShzx41qZ5otO6H4h1bDodD7Chztuxq60rRSUiOqrBQOc9
jpYOzFdzaz/lTmv27n7qtXW5cY9w0sDdlALxpKgm+UKbgXZlM9V8nRJWvv0wRpaR
NK4RvWVZ24eVQuA+wsPb4wC4mXyuQHkxQkNZS8FKgQXEKgtOU102km/yka0M59Vd
XmO0dBbsqBQhzUk3n319pfMcGAGSdIQ6ATAejRHBLyJCIBdvBLImPQJ2r8AAB/Wf
EezmPKiFDy6rgVB5IIETK202qI2Ri5er4N6facxGEv+CTYFsWg4VlhD/rCW/o1Yn
PuDLVlbDoQ6xRMCHVH49NDcqmkbFotfuaxOgQEYxgbc6FPY3nK1vfPOlMQWdEwmY
HAM0nYufyOE01G68wQHctJTLWxtfdtLq0WL0OEeKVUuk73KkARv/wxmYZDQW1++j
IB5yNe/BMMayieBV1OK4+oFY+vXKzO/UMLiHT783A3uEKPJuNtcRgM+ZAG0o/Scn
GUNkII22JABB/NbNlSYOewu6BrPCbVArZv4kheSWDVstaI+ehFeuCAIPgif2u+KT
KBtaMIj0fgNuCKv1Ag3NbOPR82qZftXaHgXJYiDQ38dTrYFcP2TejWUffffbk7s1
6zmUg7ghYp9T2l9M6cuh8uZDmg8UvQFool6ZSuWwj8YOx+0abT9Iss0O1SQenjfy
OUbmOIxyttVkirFJXJkKE1xbrOtQImCedkERwwV46zx4RqG0Krqfu6h0H7TxnWZT
ZkhpQ+T+f1HIOhB5GiEP7bpsvJz9lYPhgZqzTzqD6XWIQFdILu8BTSGcnd0j3lcf
GvPrMbGujD+97Nzm4dSEpb/TbGtQlrOr1XNT4qmVsww2aQGYaHA36fRCRs36iPa7
OzYnSZXdvpA5NActZFSrMd+9puosFRJqTTMbVlnVB6odKU58oukYxjJrErxRB4VR
Uu2wku0BNvrrCqe9KvJ+hIuNwRJz3y6kWF0W7yQA1N6J8a7n+mzUqLwDqMoKfbSA
fFbk6+sWdnqHvirwZNvsDZV0uaBqEg03hErZ6wzO8Sh39brzn4zsHDYEDTrYwYqp
XNE/OMq5+7jGGFIjcZOCy73bEA5QNSKY9cN+Jdr2y0nWnduElK3rxO3LxQhgGGaL
TUqjS+baGkCPM+ZIMptIW0XmZlSVQVfwKStN2bPrT3KUPwoS3mvpyu0gZ4mIBnfp
GTGofFrVF2YIydf00ya/wxB0oZ6YIlfOo4YeI6cn1gsuAK3kUZuh0TH8IFj7eeSC
0XOaxtrkU6fiqnqneHXIG8TRPSMQIewLv2qIsnC9JYXB7xA7AZ4qyt3tK76Db0J2
x1/5XUycd/sdDY8Hzzhv/H698+k+6wlVOiFEBBgrP0tF4T0AGEk8uW55cW8DAJ4n
E8G1hzKoYmvB8eZbJo8fJDoxXNm+IiZp1tzTWMJHXM0I0VvTCPzLKeZIepijcK79
rcgy0xUlfn0VmideXyC90MQ2NZ+vpomXkpmxSgCo+dWkOI0g70zkWlhKF1PEhXRO
iiGvL3YOcfNOBkSuVJDdJuNVBTChKIddVLBH8wL/uDQZHKw+8ZEqSrXpbgWzGht9
tdZAGr3OO0yvhaQNgvtA91MVHEaBZF3LNFmgGnWBnw9ATbbLfdlqM7iEPymaEd2Q
Cyt1rfdylQnRAaoXBl/O4uHfOT+U+xWRBkNUbo8c72NbPxXp88OrYt11FYrCIAS1
JjusOpFSleruJ7O1betPnK3H3VjQBER1JIL3rvEgl2AX9F/v2YG23qxP79O1ZyBI
ZTlzqaYds4gpH2GAVVYwaemPwNyTuFdKgBy9Mj6eG7HmBIXyGWH8CcRQv4dO4RyX
UfQVB8LjK0nmvE8p923n+f5TCcttEu5xWWsdCpS9DhgKqr5F/HVUGCxZGd0/W3l2
GEEyjqQpbpW3JQN/Y/Q+ZqLEkoeSMEppN7uZ6MC3iOC5abjNVJlSZXCniacPoYmt
Lk5IGJk4dn9dcPEv6MF9LeArRIAL9ztyu81WlDO38gUR+QWwtbmI4EpNDyDZWpwx
DRC+EjvEF1bnvKmcGmNT693H5Y11D++L65IHFEOr6MuoZrXx+13gEg+en5zp5sxA
loQJRAzYXxzIU887wiV/L9AuuFK9Weu4Y4J24wl9W+CGEoj9JR/CQXPGkmptvK8W
E9gQtHyUR0SelFeqTTXnBw/qlt4/wbHnXClXDcdU2CUaUYeD9KE5Fe9WLISi1Qhh
MeznTyhpoNh5+EfiHjKAkebRiuuAgBkbxd9pFTmmWal7PZMh8SlMv85MR5v3oVnA
pxtnu0CvYhHLVeUNV8vOKRlTnVUHhZ3n+Vw/toMUv3GUFS82RF5MM9WeJfi5icZ2
zDlTy2+sZ5sRZ02sNtjWCzub1/nLUN5ivCi8soejFharyqM6pobICmzS4/IPIaBD
Kwzmtt32PmIg0A1nwV2IWFxW5L4rcMt2PdWnrhY/I0qP9Z3b1NCUZoo1sq3V5HUm
deCGzb12g6vsoFmwuQPD7BuVjsRwINBsMLqBjx7OGOgTc+EcU3rr40LpTepRlGVj
sqXQ1uz36EZ7D52ZnML5LiIhqsRDQX00UbsW5dziZqBLizWnz1SKxTh9i9n3hvxl
412J/z1uUJ9cfDphq6wzKfqmtWBn15LFi/U1/cEf4VabCNfx9yQqchpWWJ5W8sT5
yI4gc6P+2hwxLbbcmcOmX/iFyKiXYs4nEKeq8oF3VTecM+IhW/fy62RiWs99a79E
Z/ySD/v5VwgW52tt6kldJ+iLY/wir3qq0zftoLF+H46FdjN4wMKe+MH0BwnM4Sfu
1LbOsxbpOZbS/d81OL/W1Y8NswvGEMZ2ptn9uJHInH6pZRQsleYb4yXK1tn7dWbB
JsubYf1gEZN4zWtBAdI3S8G8qI+KqpGBi/pVxPhGdZmL3Eka3Y+1GRC4dIB60gUe
JAmiscY01mDMqbtbA+vub7sSJNsA9LvJwmAuByZ0O/g8rABV9qCykMSsbvCkaawK
iitwH037/MfDW3ahGsJNAHW11nL+DJJ4nyKMCwdpjbfNc5ad4tIX8vNJR2zddN/U
8WerKN6eSTvrR1QHSOieJw1q+4LTZHQtaHPOzWB9hWn1HY5nyitl/DqShHNrXcUF
r17N6B8p/PHGcQQVw/Ja4UAizw6n3LwMKo4cQtPuQHGzrnVJvcBIaYLfUln2aoR9
302ypN4ehVldhv1SoBhiF55+OkHQrpNipDmeBwgs4VAEs5foHsh8QOs2zaL5vUJS
OkHfH19qkphhUJfW2DHYsGkHURfaGZZeS6c+UANTpv6NUfHzkuEhJJk72QdUN5Pw
Ln6NtFHIqMAOogeiiKmX3+d9m4e0RkhLCzqaabc8GdjF+dNd0CQTShZecK0BQjKb
tlF2+0tSxON4B4+g6dE5PXWCPEKM0al5QLuBHtkQgbjHKUVjxFmN8DywB7B1irWH
R9IOCJ8qJtuWJFdYZ4KFb6a+RiqjI0jYwQXqVXSLep1bb8d0kgBCfG4GDMBIxxP3
gvaDo3tvCS/ZaQpQsBPKS4C4IFMI662VRxFPDTtbSz+a9JbZIZNyHbH86BbHI0/y
V3jIWVc39TIm1m7YbCGLOEL+jvHvdEROgfEWMuYj99qoTgRG8kwv9bHPaxQ7LGXp
GkUzHpe/y81wSvspHm58rUBNub0aKinRdYEgtH5KlFktP1XsblF6jlME45qoWMnf
0sJKMOTnZtcpPHHB/Qozq9ytqGPONyX2Gi9kqwW15FIgKH5tvASQClWBJBGYEgRe
x5Xdnzd+y4FfQ35OPUq0ZTvtDnvuG4QTb0qnP8Oc7UbqC6snnfNeK9tzf9Yxem3h
F7N4O9/ebj5rt2yIU1yC4pJPDzo4HaXMtLZgS/f7gywJ1L7LXk3gUauvUyFz20Dl
PXmUM1ZHwfbaS/ZgMvPWstj6h9I3uuMwaJymuzyMNR6cqGblDVCVFAATrcYs7fu7
hsTuhcBroERSglTQug49hUROVROVKT0bKE/iBxQ9K2CllaQriM7Vl3Es8uzgkp2U
vlBf7477FYBsnjPzhIlfqqAhZjH8I8zosRS2LO6B4AMte6FxnvmrsmeGGWMCHKdI
8/70NPF9C9SCdTuWLv0pmMoNe2365/sSQQXpoz++iMDoZywupJ9slTYohSqGK/Km
AhUVIHABoN9NuZ6071ZNnM9nUrWDWWiE8pCmy6b/oqv0dI5JOAIeTar1ddPCgMAX
Lc8P+g9xG1NdKs9MjlsEz5NPmubZJ62aquW8zciNpFdmrF92cS5PI8oU5FsATcGT
YceVGfak4EPnwjfJ0ftrSmMn+hJIiWyW33kvJi8qNAYqTx38PO9ugvAucDUmpL15
Rf5yrjabPFrXL7E6SYUgrCbXPUxfEvcCmEzsqzBpO1l168xaepFbTmonAm3dF47F
eTy8zU83zGLhnFJz0NoEeA8kABIsbBk2pX5g6H7i6/SxadbXEWMgDvDjQ3RPzhNH
NmHV08htgri237nYIGcKHtA2u8eRQfQK2t5FW6AL+KxCBwmQMjqfQBBVaE+74yBe
teiwdWUEV3RIMI9twKWFrzXxoZNGRNrrfsZZBAvh7HcYB1DHIEMunmHhWf7nBIiS
RYTm56xI6/Dm2e/zpcMD80gePVnLs/37xmMwgh/9ThG4ZfN6CZHNHdPq1XNJh82j
+a+qPBZ4/yVY6XAMuwSd2KJ33e/Ex31heyNQSr3/xqMK6kdFtTVyoqcgUTx3r+D2
prsCP3q56/lzZb/U2qymhJK4gJuIx/VnmO4oq2HEzK1U6Mp2HDynaxNFBIJMtdOT
6m0Uqlgr1VxcbJZ9tuBDNu2ty9EvlrpiqfTfSYppEYTuU4k0hlmg8LKk/evidpgi
IeJdOgODYqVxRbOE7yCwBfkeB+0br+9Eb7TPEhka1dAF/rccsPEzV6++acCG2ggv
hmDwqQW7hoGdX3RRDf7WQdLGfQhtWEj5JbiBTp29euZvw3v7xLWqt2pCKi45vSe2
AXKRxfnKGzFfimsZp2JUZk+Ru2ZL2kEcL6TMRh9zcDPnt4RYEskhvZ38i/1uJPpf
imne6ODiXhsYIxvFUygk23O7XaiBV0Gjfcp++rhvTZZJyQOfayKto5udJ6UEd98q
rBVLUMUlot9FIhxxLhehSAlH3uHfkWWSF80jGCDgy60GfcFODPql/PUcruGs3yCW
ETxLvelr4wbcRHGjN2zbi/EQ83oQofMrrghN0v8A/QOPE/tUK8aXQqOQIP0f1/Pt
g4LYrKst80TXuHUl0ve6op19MpuzGNowT1wRjonV2NG5bcf2FoNNoGB05oZEKIs2
riKxZ2lKTyIvt9SrrNGRX6QzNXRem60U9HGxZ4Fa9bN0V2EOFRy9EdnQZCl8RLWt
RZIKsK5s9s3EdrpEGaDTwH13b8hK35YUSbufqRNzUPTtp8/IbNczuJgpxsW0hOG9
Q22dPdCgect+BFB5HY2jZG9/wTStWxFWsn8EfO7Oz7rNm4w5ENuDWI2I44ZErgEM
GodHiKa4wSiOi4mSXa+QQjKw/pPWwRRLr8B9Xp+Af89ilwdU7ADoEhWxF1wwK9v9
ZjX/ezGSalqixqukUPXpCn+ATVgDhr4poqyHsy0iJCqsSSeim7eFofjBAazBc3SG
icxNk8/pFd4oAdaW5ILHkZsH5VAqnqrcnSpRyJ4oYWaO5+uJwrF1EPfcCFILgBy3
qXsqMSP/UFYx2i3+qPverHKDrciSMR+GzD7DkZaqg7a58kAb/AZActSMTs7P/Z9U
JPuYKk07iYGUjym5/pwfm/VibIEkuZ2hlP9L+miM6PM=
`protect end_protected