`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8496 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
TDkIdcJUWDKCGvmrQYRemHc8P+xeEMS6bKuiqBVNXMwJytRe0fEYE9v9/pOg3Ysl
0fDtMv8alkGrbO3PMY7ImBuIkzNf3Y/W4gsF62OrvL1P19WqwgZSmkYgY3EsTOi7
yR9UzSU+1Yl8B87OGIazsdKlgqigpPSMlXkGRvk0PVUcUuTO+2NFAO+34uR+tsVF
dh0+utS7kvL17H91pVYt78Htd6SMYvpQyiD46AXGMpHBKY4TOuEG5MYAIHDx+F5p
pVGhOP7cnO2+xOepR7rT7q1y0Jdd74mKD6TGry7j7du4w1hUwmRiSreB2mo+hqpX
b+pYiEBCPslS+bO7Rka2/8lgxBej6eDmMi+wDV3YimeTznJ3G8zzPg0UPHM2KqS8
jzcOd0fdSQpNOo5nyWDCwe8hKskn6kNCmp02xdRq11msvIDhtl/7ltksVABrjmIA
fBqtoR3roX1FH2SRq7nJuVvQjVTEQ7KJ/o82BU1TURS02xh3zGzTul7VVA2jEGnR
vIlROLZh9x4/TuzlsWhvsEZE3nuTFws248VI+fl3XMKsQdDiFgGZnrnmxZABq05N
kw3k8CR9v2Xm7JyrIgd/ZRWff2sfB1+ByAMKuWJgf94CvxKhUP7SNxPobVdGRD9O
FDPzDIgJzhwbQPdDdfsdx6fOA6kYCit0y3GNCcv5doTArK7x+DpVAkW0CCQSRDUB
pCopZBj4HPWW52cl5/vGgDFpg2lCezjagAY/A2snn6kZdFfX+JS6VJPLzVqmxjfC
MvCnmiIDKceGGO2e6QZ+PfXeyk6VG/HR3r4Hx0axUHsDuveC9Zu4SSt+QP+GhEDD
IUJZvOz7bzmAGsGo4nqq+3whrrXFxTZSqK5UEIiJFsaQ9zAY+SFzhxePxKmF+C4N
7UHCQlA1QaFFRfIKOlswnAPD5lbfq+jOn02ptOQ4zlwX7r0JRO7c/z1ltBxZ9O0q
cwEBvhvpcp2ECAucCkA8nc7BlS0da4/AJ3SMdI5pLHLDgNSXhV1EXOSUTiDZGFdr
aQ+7fw0FSLq1KfxNn4Cot+P/vuHW0r639SOXZYmeklXZ2iQ0qQnhV215KbmjBssN
PuRT2hQd8vlu3yTFc2Zoi71EEq/V54k7urRFf16rVS/j+Qx1eUlYvdx5wMOO2eSg
jv/CXLkQ6TF7Eujqu/3lahL6sSKl7rAWF2QUq+vijj2dje3+WmQ5rej3w1vzEK8D
NnFamU0bn4hVDTCZWvfo4Jhhyypwzdl2J5i/1umCte+5YZQYZX4hGi7nT/xLryo8
Aj+joo/8GAsFVFHYw2hpow+KBdIyE6gN7WSx6MTxMgDv6gshbsO4uo8Zh6XZIMCK
1YmLRS9CAzZxYihdrGgItARGjxCv9SA1/88q2brOa5wgJdNBCdKEY/nnUXYs8aw/
aSuDck44lnG2zo0jl4hNk7ZumFFSTX8PMYjX6QeZd/TK6mj1P3OmlgVV9eYE6mPz
9I3qWeh9b/dYlCOP7JT7+KTL62MNV+jlYwSjzUDIrBcszW0v4b0AKiU2+jq4ZNZT
ZbiJ7mOtDtxF7PVaSamWKHF/O8N6h37wfCeXf1VOKmvmXpsgmWNt4aNVCMe6f8fn
uku05besYRs3iOwzZnXq+c5+blYHnoSiP/HtM0NFOyMtsj33PUepFFzG52UXfFOv
ruze622nbVrE6SQYDGhAdV73cLSyUTaiQmwU+lHqrN2ismwx08DEbzLuY9ylrUhu
dDF8znpDWAHTv2ElNzjNRMRgzNCaCxHgt7JnkImjaaxFxKOHs7ofU5+eU0154SnJ
v8GFyrNMa2C1fIKMWYQ0O96WhK2rlh2ccB1hvT6upTlh1pwtU1a/6Qk4c6rAoqZv
KG5wc+zm8H23LlGrA1WzvdIXHy94Vgyd4aar63RftfnzW75BhZREuEEqtjNzLgaV
6ZPJKm7oEY9+jY0AQZRAafmsN1AcDXcZu40N3v7rlh8a2c3cArJM3FrUpGb53QeY
z0Awwf2oN+78AEXuTjh+KEEghC6bCuSTT24URXxt+BGoqwRKPoEc9yQatXlK6+Hz
Ew2j4AA+P5kadHg+mkDZOBvd70GOVNvlRuuzgdIPVOjbUbiwbVJ7zXo1bq/9tXwx
Kn3463bLQqgQRT2KnIxBcDt4+mGGNvHV3cwXrZ4PbBtMgdmnsqJ52QVemKHOhF16
AK9e5l/euIB1x6fdpmn/ECoYKrbmW4aKe9buCBBLzh7zanaIeO8trwVZvLMIXECx
2Fz/DXjNItxtdRLcqstAktM3sX27TYM2inBPjso4D0jLhjjO7/QUJnq8EqV4SseX
60/8XDL7fsWWfZVM4BKdF1AE/Y1UsowCUIYx2KT67oiGBC52vpgOYDCftY5NYqm7
lDI9Bs9ZMDSjk5l3bAzsvm7eXy9HMcNeTEHocwX25TUT0KL92MAKMDlJ6F4Fh5w2
Ac/EwRxfonM9sJ6Uy4l00aPtqN77mQ6e22nx5D+Gkt5tnty6vmk+ANqYZuDGnuwN
L/Fxzb2z2guJA7aGwL9kOTB8OnRdCzVjqRuOaBfxMWxH408ZELO6j8xbLKDQ5kT+
pZJ9aYYXLt1i3pewu1LIPlVJ3lRHG26dpip8TL7dcCslwOnI2wGPSF6/1m13upUz
z44ICc8+yxiha3r0b9UbZVGzW6E9zxOyFQxSeZ91U54EW5H1juejNW8G4MkySq0D
h0JdZ1LPrtEIPw+AJ9+s6w1V+3AmhIXhIZ2yjICEP5h3POGoXgtFHAqWpWKnf5MY
OuM5whZVBbhpUFVj7FALkaldZne9cZytrSSngDWKHmuIMH7xh+0I4SR4qqSJCc61
PdXkHgcTUzbCQARi416C4YEecPThkA9YY9lF4kLwvZi2jPdiQeTKprD2g8aktMa+
+uzmF3mQVRr0rZPbACQg5LUJ2Jgq/PnG8wCHMOdmKfexskMJ4Txaw2SYg4whbp3y
hbkKIMAg2bIzegP3nf13sDcAK18AWuSSyIaWUzyHigWs2TreVgYJBDD4WebhjEQa
CCI3kPUPkkzKq5uxeP9lYBGQn5Pf2Es0D+fktgaQzqA7Ubj21AXkjpSE4vQZy8z8
FklZutX6FR2MdOfbUUgWprOESwUbLT3iRB4TrlGZ/aU9fBLW2F/lqkvU378g3c1N
5KUTQpqnoG2+1MK3T48yS951zALenykv69GAzDr6QpfaIRf66bFvBrll4Iir8r8V
tFwg2HFGJZWfekYKhxFoVYqv6q0dxuuqmOT3VDqq3Za+oJdsjCs2HK50nwNwrQs3
kF/rApKe95upWogbdxf1ADCHGfdg3zdGd/AONLpwd7xML0GytNV69tyAS+3hwG1B
OtM9QJsu8mR8JrtK4zRPLwtr9bXXsTjztE5tUWc9snHXan0ae9Y9VBgea2skWA6H
pfbh9YUtHHOfMb83ZxHU1qV96qq7VK4FxYZ5BjGL1OvqeN/43O1kLuSyTshW7kww
Tq9+f8oG4tGuusDuSzkYiCBLNm5wFNZ7r4mx9jvei73+31cSANxaDlYWToAD8hob
fQ8pNSPdMZp3Kk9ugQCY70/x9LB/JOoZdaoWJGj9ApC4RvvCV2uugfH8uu9AoW0y
a+z9V7ORSu/uZbKIjRo27NnK8jnUmyDi38/IUiP2L9K3bwo4o++csiX44YMfZ195
jss7lpiQEB7/ZKzwgqhcv4M8aCw36/hqPp9KzlMxTYms+H8u+fu7XijcmYjrjl2a
73rhY2VfINy8eDJQtkSYCpZ3YXHelHgVfom56KVhwIdEcoQq0kk2w2SBNofJewmv
7HWXnBJsjux0K41UYZhYaVyPe3qjxuWQtp4K46XRh5c2v2g6hXpNSj7ZLhCYmaYj
vwIyz65vZMXwtBFPWU57Oqt5DLtUkxrLqly08RiF1dh801zgGCLmOt9ZY3N9YEqQ
7scSvbVensHpna/IstOWlnc4wYJgmEEZ1C0pZ3s3tOoQsLD0lmLib6R9GGmju+x9
ccPw3tNTXiNcG83L5MXto4ns/Aqz0AZ2ekguT/vlBmNyXQQB8BKfPLgqb7+4bZ0Y
eGZDjD2Uukjo43KDXD4RWAQbNUXWHo3CgOHRk8NS4P+axM5jRP6fS6OsXWnKF+jJ
v3Po9r55ZyUk8Vcf3hvRIzkYtN/Tk/lUiEWDZYa/u2nlbGH1dJTHSdY041vHpoJG
zaBQAeTkgqwgqNQbbVxAQijkQCoG6AkYwm8xJ02RIEamy+m5yBZyLS8PutqwG3Hq
W8+FfLoj55EerDx3U0GWrwnqbq4hAs1/jeUW3Svdz1y2enLQA7KJwFtnPqMuDBe4
LJAFKHY66PAw2M8Bq3C0DZHjCoXSnHmPgE0dq8Bh/jZz88ohr94Mn+0jEH0jo2De
iQ4u11t+l4fNkN/fBwtv/vtHP/2bl/8+yksmQs3UXj57t+cZpuuOzfPMvF1qrD+k
8maAzxt7g/hkuLnk+knNtMPyQdsR4YhpW/eKn88r8ODNOjIhTFVHewEQOUzJJrfc
xezbBhrqZ4KLOOmSEa6i6ALl5jorsoM2K/oeAJzhcPG+LziEGdqV/GF4cLX7Jfe2
iTpsm9qUCJXnBuSPg3Xi9mhgFAzt/ikuOsTpetg4leG4cmL+lxLLYUVxptKRZwNT
exsmXjOUHdeqSmtEtWcv1dPQvuhvdc77V1Q8w73kp37zZHMr5WFIDKfoFwHwotEV
nmnmlX9axZOycl9vfA+FuIgLA3fdhCW1b5RJki3viFSz3sljHohnWgiej/qu3p0c
5ijNe6RDGKveeb+czDe/Bj5iGH58MNgr89BXVOcXqECKSa+vGVEn/KjXAxtkMOLS
6BLHSiSVyjPxCis2P5HH19MS1EcpgWV6scFPsfJNfo3SH0MzoejrhYgaDbNSxfrX
tROBmAYuoEzZyiKxtBVNzWlq5vB0Q8LmknMhmKjm0vQYJ5IvVCKc3S6/FYFrRow7
/EZlsnNKD6I/kDEJcVQRnhHZOW++ovgPhrlu/hbVGX38mfLUHlEcKex+O/PZKnq7
zAnYhFCPkTDs3dgk0EKAD6ZjDrH19eeAik3Yi3erRGI0ZGFT1mMXSC8FZgS3jP+u
MIXcW6O1ETKFlskOz2RtYOa65l15b0duY0zpYmSjAQd8VkucUe05n0HrUM6W+tV5
PS/du4vwRCcdnxT+TlIEfwTU/bbiHWqIVi468fVaWmv+AsoBCF9SqlJvV1wyr1Ki
dYo921NJxl3wQBRyAdccclUR81GVt0MppuFTs4SV+InDKttB68a6rdG0GojU8cxF
Q5WN5NY4vDX5114m76Xke8gU72yDl73YyhjEgkx/DGj31tjDi9UR0V/fVRRF8aAp
JYKJtdl/hxDYUqXA0ukeTIQLahyDnVs2MA4dsMoXapPl2nKsimIxISNBLve6Lze3
3d8ppVyX0UmCnGZgOrbaEKUpw5CxGGPnP+TUqn4ylzdqnwbel5MgEsAMK8ing1CR
O1XR3UT6osV6Key3ERbUOs7PbyL4CcrwdbmsU+EkWuv8u8xp+h1VxvHq/CrP+2N2
p/CFrN6lcUHtDdl5+0J1DUImzzGG5zA/NXQBaIGJn/8IXteQcgZ+/yvnufYRgpTZ
yDFy/CW488sycSJD5uLzNpWhx365HkSC2WUjUyNKA/Gk/YnDbgYEU5vGe7J62e2/
LHhsNxvfFw5tRA7m6hzYNwRumMRApUIiaCUiVUFEvWb6Qd7arRskgAEpaG+GaOEt
pvAemj898qfel5ZHvcR75vcp0DHAlxQ6VRD9THvVr3nhg+TuNKCHgS3qSGqVEZ15
lqQEojzou7+warGoW4CHzs3912coQ70oT2rGnhvqGYH2ixX1D8e+t4eD/kXYz2ZA
w8CZWYI4jlEvkKvq9kMCI3KTETHYztDggDG+9DmRD+1Ta7z2KZhjsA1H78+7nGub
UPOiTTYamVrcoe6HTV1zeltJB9zycACVhyFsEE47W3Wm/bD+fNw2JLUXSDpd7TIf
D/g06qdX9w3BYB2I35fRdo6lJTqXX3BQ036uzB0QWBviQiQH/UHJp6PCniOHSJOA
igirr5/AQ9Qlgwhap4tZf4BXCTPDmm5fSjj5hw9BoHFAAXS31zxpHY71LkpMqF7C
HJpU5YQYmXMN+w4648fQmDHPHzV0wPYslah7m8mk4p1FYoW+z9i+eGTEoMiwRAvB
RaP0jG0D9srLLBRmUKgusQ7uv6P8yC6R2EWWGMTbdxgjHEI4URql6Zlx9uO7fuAn
cJhulTFXxSk4Ga1t3u90SKkG9eOQlO/zzJZRZthZePn4k8sYYpZ9+QxsmAodGaF9
tpHC8joNnyU8GRKAX51fMQt0FmAMx411fTO9b2k0Umicivn06ewhU4UmPniPllLt
RiVbuNb69dvhs1vQebnlwttfmaHZc2rs1fCQPDK4vqvy7+fvy3Xk77azrulkJUzq
XtUQv7b/RVVpJVQOyulg+yQgONhZEJPMSWOTI83k9Gm2c5vo1MsgDRu8Qye7MvNF
2EIlc35UREfVxvseSnhv14VtSLl5z0c+8/GMOjOcfj6cDWlT5ALaZUyysa/EvTp4
y2BlLniS4bwqDv3eSYRXuk+fZbIfV9blWbBRq0T9TC/OVbEn0hOlvDaSoD5TudYp
SPTMEBCjMG0TJZTqE+PLDADM/ivWDUjtkBLlfkHNhhX5FUDW2F7t/WOUJObrdHSr
qhMI+TwOK0vSgQ+YleGXiuUt2E0reIHlUn75+7Cb259i4QopoN/Ycav93cC+XXTq
O0lHCRUvNr5yifj6UiwOrtbUMhEJNl1QoqvZaFIUCFeuXmFbSgiFjr1icbUGz+na
+MYEvFFfkyWnmAI+VEdm7EgE0nHV0abXOqWN82h2UM9F/x5q4ZNhAv9hymqrVILA
wd3iNPOvz9cW/eoqbf35lC5Il14jzLvLEr4OeFMtsqE6hPOqHQJq3IgPfzJrs3BQ
Ng3JUNI2h8+Yrgs5Je2S6+qX2j8f3ep7wi8E0Y+F5IXgBW6RzruAcQ37yalYzcAK
rr3goPE8Wf6mz/V+gidExHVLwg69fmxFAfWPCyL8QKv3mpYI/FUK2TXV1RHAcOxY
hfErJXAQ2rEqQ+ImZKXJdwDz01aXiLHsJEMCXMX8eAiuIdQk+QuYrUob5sEg1tw1
qEvLZ2pvQdNIlk6csmKOTyKRI5p/r1I+pw6/usSosKviOPG1q+UEbRiIegjk/MNs
n56MB44brPze85X1e+TTRsclWaLGeHwGXloHUu+GLvvH69oMCoimKfmEPxBEPYzb
SFR6wT1oTCbPrQi55m3Fpt3hfvRuMjw5i3ABKZXlj0fr0tkIE1VNtKivrtKx3CPp
8LcQ8jex4pUGTp8iVbKiXrN+PUCCl2n9a5ZC/PEd88xmfdCjdfjggqcP812QZ633
RQwi8jjgx6QXvKQKMJoxXOLg9wouIA7xfigkDmKK6+VTq7c8nCYqPN8vgp8IrW3f
3Rz8MQKl3LHU64g3Z190oNGcPl3/R/wRSPJjLUlBBhiYKM5thzW42bB1jWGnYN9B
LFCZ20QAcVUxZoWQo+jhFvmIMsrCyQgn327YLh85h+Hc/yt5z35tceVUm1XYZl0l
KCJ0HyKHUG/nEP2y+77nBnvSG5Q3KhcUr2n+NjuRfYw3xdDaYNvVrp5djGx19xxm
hPWAb/RAQOwrTyY5znL1Dz2+6kxCQi79dkjcgQKceo8US5hfrTi0y4d6OUTICR0S
mKX8P295/klHZCwVHFrjL+ztcB/HeAoIc0h+VfSuyOqfCnhlZptronFZJIzNRvgH
0oxzqDbruWGj+805ecGx5qi4Bq7KnncL0unEPgOmJklClufzz4jM08CyFTWzmQeI
AI6CFpbLYsG1ax+Gdqqc/703Ue7a2UXPe4Xsqo7BIgQU13pASVJan8DH4Zb1M/8Q
hVayFedSKWiB5fB57zGLccBR6Ocf79j0k0R72HrMAMjy5OdOo4OkwBCAFYSU24YZ
yz0oQeSD4r6MYQgp5D6QShEXdY928I7B/5bXBYNMIpVLH66/Pj/atKaQlxxx914N
rh3i2bPkRptOnAdYVnw9e6wG9gyuIjzPi2xC5L/UtaCp13HLgP1abBezEpvcUwLv
HKPyEZ5cKJsBfookiXJAxF8qxEQATdOXX6wcGovLBPxdRLOaomPowOXw9DI7Uev+
DpariaJ/Ane4peu2xaM7fEvSmdMyHTlYDVx0kUBt9i6HO2Cevv2OgGs+TTTj9Fxr
fT6J3iQsK/AqTUIlrILMLe0SbEHO56bICmbAp3TrXzHe7A+pvhQbsGRycb22emd6
GsH4/8CNgOUS3KAIOqaRBgnVNqPMUjEicZTFZjSVGyP3CMBbytTqCVXx/gWWjZjA
f+hKKMdMsxafVjppweeK4ZBCoGPI/OplTvno9NDK9laxDhcRA6Pw6Y9iVpYtkCuz
S0jWiQGMUNIv4R/zQfYmQDZ6WYicjmuw+N6WwbGl0UQySne5jWpm8KyWrycPm+XL
ekHKOqb2M2o2S5w21pKdH3H54mLkj7mGUcOS3qMCNHLOCk1qbC7mJ1ymC2L7fd4h
2AGYznZlHx66uC8VgiSl6tCiZhF8B1ZQC6RsqMKncPn9kFSo0ZEFOfnG5RZv9tLp
loWZ6HtVyG3a9kN9dD090uz5M+naHdvrFISmukgpVac6PY3dCeWG9H9VLWTb0l1+
mFlWj/Z/vAmmKOn37wT52idoB/3UwEZSk4fSVlOn5hbuw7fTMG/HtKm4ZZRiOi1e
jrsg5GfEttk2wPBHb0x1QKPA9+QdIA9shMzB3NqgPq/3yYWtmZENjE659Xv6TA1q
LQq+nzpK+QXIBZ0lzsJhGuTgpFRakx4wh53GP2sUX8xoqEQp1fQ8u0uZT9MY+WOc
+SagYiAyUjWU0AXMb1llEfy46LY4oHmxmE/5qNE69Qgyr1PigHlHedzMIZtMXykZ
fCLl4mDzYq2V57Rw8meAVzrSCkgUXj3tVEVMt3mXI5TkRfdC7DMZ2lf+L15o9dOF
xQ6zLjr6JZqvtSgSWLyhw+v6kGQh5G4+YbyuITBNqc5hlurs4hkpnR8X2H0q8IZo
QdeJmMmu2FrnRamSozTrnsvDKKk/kQK3SZBlVYXyF8NZelgorALBD+OlJXeUwrsz
ImhLXuJAOB/grbQtEMYWT9HyW5R2LvC+y5BOCAuHlPKebr67qrpX7jDat81ydWll
Kdsf+GU/ic5ATnUeex/8wY7brwOF1ANrI8Phft1MeMlLMC2ACwkvMdL9MWEbrHP4
YdgSWsQpJdBpPW1J3ve0/gsvnfnu1Zz5uiM79gllfZBQivMwBZGGA1/HqRW6KxE8
8EGJUAbQs7zElON9J3hvXMkXKRQx/LT52XL8g1n1NLPB+Jv4DsMC5gsWnUyKaJVm
1vr47QgvuaVZIdhP4sYNuxyWQIhnotsw2zC6TK/diNzMVYUCb0v7U3wyp4gsfFvr
P5Qryg04n2JNanMPjPVeiJ9W6LUIJwm/Lt03tZusFJr7E3mN2o41ZBHJCDOJPiR8
Gux2JkHZ0lTZn29VW/MFQik4VVZdi6OfoPCgur91bt4gq0yjbcr9FKNSmSlF2GUS
6kCIXi0JvAp+05Fg5MyingfspGAWtAKbz2a5Pq4zBScxTcaAvcP0NWDFHqRux9Ri
Iw7ek4JeAhLZgcqfCzpG2Zmbr+ClWhrDMOlu68SbdqXYP2Rn9kMRCDp2hiEhyCsA
8ou1vS3OLMrfLzODZImQDPNRJKvGvlD0QJcAnA38oV4r6AFizWDg1jc7I2IDBe1u
wiF5uMjn6zI59gQl0Fn62C2XgX8Jsw/X4jatwalqwoX+Gf1YBSlZA+Ajh1AvPMll
Ntun7hkF+rtydRo/Nk9lNjBvd3qXnYG56cXc4Idl9a+YZoQNz8LGXgONwU4a/Jkd
mW5EXuMBp0NUj2TOkOZx2b5A6VVAIHuFUrdSeVytipl0XDyY5AWsDssTASL2Tfzr
yFskADi6aMfhZgZyyV6YXy6phHM2eHD/b0NLVuXH+OxWKZSV/6sN4GFhrThHXhGN
X7khV6npHzvh9FzvmR3sF2WQa2jsjjFHZd0Nt81rRy+jgjE9TgUdwwq55XQmPHQ+
6r7RRFr1P7SJnCRml3v6gt4zKFf68Xf9U/Puq3U+bGq/uILlp22WL86j0xlhwMVn
mMdNUDgXaaeIflxRDMcsAT+aBXle7bM5LGnIVgOafJhnTU2M051l5wuMh7XSxsVn
9qX4bUoh9lZAPbTthCgsLq9Y+UFEWxx6AalP4aa+u77/K+XcHbk57xJJa0lxFd9v
6krHdh14yv5eVqGesb14T0xIul7eP8QESitQHhmCxCSrDdsmOEs/HowvH4HTwMPa
mZ/mU8Ait+SZ+Eh2UCsuzWi5vvYXioactc9tXyHASSy+TIRyFtXA+FkR6llBS2t/
JRFehY0W8T8bhdAysUJoZJmDznz3nfVokL2XH9eLUf4xngMCyjTJLcNPrRPxugAE
lQg8zYbTQ6CcYGK20/QwbRkib2ynS24vLdb8tvMwinTfrqpuZpl+2sXSxHCyGjJv
r2W+vjl4T45ciR1U0ghogTZTIXAGSeKKCVAb5KdMIOTAN8SPLby94X5eZsb04QII
11FjO1npgw5J6KEkXEs/oqmZ94l0l9fWSk/WB1zKtp9M0d4/djjmfpz5HsPZgg1C
0oq1wx82Rc4YWf/xvD5WvJUZAc6yLKNAMoISrltshFsc2TbwvwgHL4id1bI1Wsd8
hh3+1RNruJN5M24kbNHDsdSQE9svSeXbPHuEdSpKL0gVlXr3znZsv3o5vPBvTc2F
9pzQfCHIEzS0k4/PB7AQq7qtpYjyBcO1kx6gh7NHY/tQCkEKd1bZy8CgQ46FhmMw
fIZcxfRqaXOzhBaGlEy3Vg3dHsl0jbgbnCswAftdzbh5hUtIsSB2OG6ewa+PFlyb
g8MlHiVlQKZsdvoGfQziYdOoYuZQ+KvtZjj4o7aWt+LAEOo0NYKCivqB46FJ3AQm
GA0PyekVswfd5N58611z6d/y2AhX7mjoGOSzuywkorN466jJ/w0N3O4ZihrKgoUA
uzHJl+zHpL6Nyzky5QZJizveM/Pjv4+r3fiCjLQY6hNpkVD9SG6EvEFZneCw1k8U
QnLld1hYG5bbwxLJYleMcIsVYmUoHGq0JV6igxFCevRVVIEjCp7r8DheoTTAJnEX
LDPILk1g7JDZJyEslqjpzloIMk1fUYd2hpAFnrOn7p+EXfY5YjfAqyRzjjJJPvpG
`protect end_protected