`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1952 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
OyGGrfLtuV/iB6oXYN0vYDeZB+mjqTtsvTCs5yNhxaehj8Q7vEVKt+5ZG5umdfhe
lvP50cxD4soRm3FQ1tQIpcA6x7XqY1W470mNS1zSgeJiSlZ5XS9dYyOgVj8Ri5T3
8uEHwoGf2knpvdA3hcoLM4aeaZOlW4XjipvuSnpf2kRKFMpLWyMu7eSLdCsSgAiq
qAUoQsAkXUfOJocJqJp7jR2S+j/c9We2oo4A4zI5J54DoNLoQvceXZ+wQq6OE9lE
7s2sdV8SjdMLnVec44a1LjRu/WrxaLAZxDLckpvFzKQ+0NjFc9pfGJKQKxjmk8xv
aj8hpBbjop4hGv1BWH22Jt/veniZ8o1fLRW9R8iLQzB+JmIGzi0n9DhsGW1MabtB
MqE6m7jj2G8tnjNz8lyMyBX2r1Utoh2tkhJQfy6At1ueqM+VjcSbm3xHESMstNaB
/aCrF67yWpodyPg2/aJs6Gjuyz30K0j8gBmJEf780FhGlOIjsTrBTc3i926a1zf3
Kyg9yBeX6Dj6l4mVOKYwwhslHc2tKPbmZ8GNFLenlL9JdSuFwIpQnCDEm2r4qkLM
L1F1mrZ0fl++SpJaptA02sgBdwUyRGiseNf1LIeuEqidYf627tLPJyAHTVIXxa46
lce4oAhDZke3eV9UQ1s/2O+a7ngMF4iJAjBRZWmQ35opTzA7wLePOQu8ntpzO5dG
mutD3CCHXLVVhb7JZ27rBOWNTQDAcDI9Rhaenu7WnPJPZqVvVFjwjnH2pjPmCjlK
zgHUQBUpoiiFS5YlU/G9ozw4uWiMMADPo9TBn8aRsFZ5yGdKQ/wknhJNCbu6otKe
u8V0L/ichgHHhIqtt+zCER/rlngdjBegIdfLUc5QjjKYLU9/euxeh1rVGPdw1WT2
asBHcJca+2q8CBPspGqzoCr+lv0pCehcP4QgmwKP2quwJRs7XnerHusTouqCaRNn
f5AgKB8YCRBbNphcMnhG48OwBbSJo6O60wcK0QimB2+R3r50B6SE9j63RskWadJa
cFi8VlU5FrinzsZY6uS51LnAaC2wU4YLyFGERvHWO+mDRHK827m5+B/5ki0mIK9f
hYokclPE2E8KbxyqbLdtCZap0fkgB2YPA2yl0sw9TI1lgN13V+I+6R+COsTHRz56
eKg2mPLJDW8RZWI1aj90lO+evF2GFgZxBsudsvRzQovkUeeeiUPlKf02TYqDHLk2
sgnAeS8yVGDst7O7ckU31HlRCQUbZWimIk0bwOF1G3iHKFiXtQA0xnUyylnSsvcZ
TW7dtTDsuSGE6zD4HbOZI/TlihId5554GSapn8LTJ603SprWsFKM30BBvHkn13qm
2fKN3QFSJ81Ca3lGHTHG/B26gajTH6RdY4VUYVyubawdSYKynCURnQz/LZ6dii1f
NIKbEk4q+4eg/ZdjN6o6xsg/PEljS37p8BuAbKCTCnkroUco004DeNRRTvlpIErX
Q7bsJ/C0pOcI6JeFrrrKgQeNGwr5oaoKjeIR4A2prGJQquQc3m2krCIRxJo6t3b3
VrV/SkshUm4cJp+hZ5jqdSJeLLCBmmzoWIjPFd7rAjZn+iOpNYeukcubV48gDJ6u
GwL7R3DFtZgVKLMDqQOLhq+9K7zZHQxX3GJYzhU9veLLG5YMlhc6cnu9OBEkqOwO
Bz+8atr1bb/hqeJSTWfKlHs1bHzUvaUidUlxxVUCnIxlRdXeFyv0e9XlVqIfEmMC
FHf9qMrstdzPnT5T4wlYRZUqL3kUhaSp98+ZvMuE8CGQ19OtqPB3AS4OJZgY0PSu
BVOf7wgLVtJsA+LKrD0n3v9Cd6422MqYUfdsy/29Xzp5okrI7jLeNaIiWj93yDHS
MopF3SiR+yrF4KFZMTL9Ju8xvkAeUaevUdiItFQFQpB5wv2ohRxbesYMdcBgg3yp
KcY8ueY/NOi5PNDBsXuaIE83ovfS7ckf/ABLdB4QDruHs2SrCBCcqm9s3Pss/lUV
iOI6m48+8KIP0w66eScerox2r+tj/h9CowJ7nztI2JguD1+31XVQDz9YY5ardv23
bw2aaj2mhx2/rKzgvm9hPubVjoxwISwLZm2jbB9tZ3BGZTEonF0fJGf0IVLqxwhA
zCzP/uyxEZFwtCsk+UK/oH71hgQNtjpLgn50or+Bg5w91+PqxVanxEY4P+cu1MY8
Whwi5BiZWoPnimwn14xadLXrj5jAHt1/els8ns+m1zTQ+UgqxrkBu2YfN5WpWeA7
txubuQMV0JEj/3sWW/4DEb/N7NHrRVA8EI/sZTPrM6DrSAtvvCYl6HlCFY4VaCMi
qSFMRPRCSVhvWs5tW8FNbAk2hvzeDEo5tJ9vNMr2FqzcLMvMx2JCIZghD2S5yJ8D
VknLfgc1gd/ncXm4y3D0QYlmCASZTkOiAT5X/Hjcw3W+bNb/uQqbC1EkJYjHldxW
Pb+y6L/S2fjS0Jc9xUdxm8nqWlSR3VFeI7QiR0sSQ04=
`protect end_protected