`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7824 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4sSkgcOrtFFGmnZEnVbxgx
+l/NC0KUoptgPj67g1Rb68BgpBHvUOHuD0YjAAf2WUHck1/K7oUZJmK+Ydp0p59K
Ad8aFAIXS7b3JVggm7gykqomP5aA8ZOqFxjqCBG/69XilUS815/GFZhbClYPLFkH
Kt+am4fBaazd+DwHQ9b3ZFcLTt1EKd5mwu+oYd1/hVOYOE5iIi0PsX0G57lplZ13
5eCeaV4ZYvR4fHo1EH0LUvg6nUFwHfZiPgcS8gUUAYafZ7pV497I0GPdOFb4CKej
r9h1TuHGMdcF0DxRi1nr26UDsbx7L8i1w16aL1b4pZfncT9foKlPCFsWy8yHti4q
/WgJfBoCWZ1bpL9SrWCWp0NAZm+Hwkk71hi1zElUQVFcyd7HinIhe+V0vqv5OyMS
FqXo6B+o/TFdIjEuVQC/b1LzzqCPN+CO54lWSrUUv+grzVJ6iE31nYoSvXvD4ArM
QuT8bH+N1RMwVhPfVGR/MJaPzAVphVII74C0LzxA7vHhDpHoMYW5vJoOj7IH2En9
o4LY+/l8YUx6Itvk2QQccxgj0dkn67sZ6QeqRn5bv8Se+xcEXOODzzXU6nzu9LU4
qpUlf9L3/Ybi6B2LWkeTpjJ47BmuS7OwUkaFB/twpsEFuiEeUWgGctwRXHyuVQ7H
MrsjVI+1fZaOgMia7L66IGZ2sY0ijPP1XATux7RNpGyXdQ1bVXTfdoXrdUAAF6EA
7e/WTWLLRR+W3y0Yb3D8M/WEzG/uwYzhchJSD4A+jLEilimiM5F7I5AvZZLRX70Y
3Uu3b5sOg1Ick9VOpU4CemY2Iqsk0ZWYStkaIb39jtWBWNqg5Ugm8uyDSLkpvKXc
W1kZcEhFIZrmWtriY41pWYnPREVgoRbW5348TxK0f8ZXKb2wPDokCNM0NY0NzYbw
YuLBxE5eZ8UMa9FqjIXj4HQ3lj3ZoY88tgQEZo5QC3NT5iMdqv9PAnDXRVqcrMy1
/4CRUeuJOTzPli5mnx0u0jPnY5bMc8VQNPinC/YeTcECxKMWkOM63L8euvq7NIUV
6bSzi+0BdluUv2mHewQ7lu4LyrfMXpap0vUG5HI5zs3SV4AvjmPtnCoTk7VJ3D0w
Z3hfISnlsTauOJ9TwS5oVnj89IUmmuebWm5OVYrKiHARZ6jgQ66m5zYErnRkY0q7
Aa/Bmy6uRXr+guGxGLgr2X/bOZfvcl3Ee7wx8S3e6WpAG5bJBYcZ4R6ae24gpKdl
urN6dajfErL8+f7dikHZJccbp0aocqFICKuJb5lBEOCtZ8QKSiJ84KuUErDokzl7
d517Kp5PJI7EzC41FqmJbuK3RHkNJ9dSRlMC65c/EhnpyCO1zm4pefkXJZHCU5FG
b6ZxVE/cQGp4GMpI6+O91P6sOQXVkV1cFl9bGjatrgAtTBgR2lkOVZw8O8pUWaZx
+oWgNYWyWMwx8CYr9Gl41qPs5h1d+kJjwZ9bDHyOMs2ctyvhT3KR0Lda+QdoGXW/
v7t+6Poec0f1wbG07dAAqBj7pGsCX42qChF5Wpk8lhmM2jlQnbeM6oFcfyIVS7+b
XwhzA0dUIxqMueQmXP/Ibxzb62lBxNaKuwZ13yexQwWNdhBUdTncXL462VyN65ua
gHLeG9l5pAos+kxk7/LnowWMXiuDuPKfJHA9/aO6ykxyLDsRkh/NuA/k1xjVCp+A
pz5m6srDYxvCRPSH5I8K9HIE92uemGemp+9qnyh8DEL/k+UV09YdR16z6w4yvpV/
vlfYpIes24H0t4dIeVkTgNye+d/K/zYbpjj27O5i3bnWBz4SU+DWZFnKqfpGY43A
i/+rcXDPeBM61934NF9kVI4OaoOpiUnJNG86kymWyx7FgfByknDT5xbPNcfEAcB/
0RmMIjY0HgDuZKR4NPDxF01WMpm/VpAJW0YP+l+n2d0OtdIzECniBnTxoQuHZB6T
cAd0KZ2ikwzhehGepI5bTrH7fgi9xBDytmE2KzCpNi0qqPvRmnftM4sC5hjWFUxO
4ZOSs1kICvMvL27gPNzh2a9vRTPcUpNnc4hpuDfMaXhjI27xiIIuC9nFWkz3fRSB
NOVE6lu76SDuNzJVb4OPrFQnzBA/sgJHRyWIRp1SsAamEi/WtnlD0p3q7lB/lO8a
QPufMn7Qsrw7bNXC6wc2odRFmikjbbfP19Qr1vWnhwperu5GB/dE53Pfty8tFEAq
pvgn4qcASbY3v0AoomL0juS5HdB7SgrqEovE3gDCk2X4c0p4qqR2Tkxn1mCYRAet
O4+IBz6bUnQMvH7dujZQckO7DbXb135KLM1QrHkMwf3GWZqbVUDlNPaR5A+p8BXy
FOSJmrVewwFkghhQ0ZbHy3PZ32wM8wx7ljKQoc/UrKAw9ll4rzwNxINUo5pkAyp1
QZH+SHS4FoXZBb9dj7x5/Yb3RhusnB3iIz1FyWx2R3UsHB5E/Ew51LOuWl8pfTBx
In2LdrNkWexJetiQzPjACZFIPNC9VmYhMMo2pKvzBNleD41Ygor5vlIzbSLyQPYb
Mqk0yh39RYmdTPRNYwoww2R7XJTKvYWCrPT8eaVhWsLqprz6vP0583O+/gW89BAh
AEng33KDnvTH4xJr+9vZb9jqn4YFsKqm8IU13bDrgz8VB1+tO1jygjyawoK9HroH
FmHYnwIrYs31b+0yOiJUoGKfWr8jezNZIsukoJTBp9c740938W9BtxLGbQE1Ppv6
J7sVihBr/USIxz9hITc+hzx0LFGDH24VnFqYpxyC/fGtZgW7hWbcblqk4VqvgG41
8uQyoJ940mNsai00jCMFluZcFP0Erq4MoVWA0W8tA/SUmeoGYQ9EngRYtH/oFBaF
rThCa7dE+5sDESaIvE9mDHIMAb0uz24SylW+IHQw2YafhQkUqx+cY6E/N6wWLEbq
/AYv+qbN3t16Wr9NnNlsAG+/EfC6ZnCIOhHcFfxStPVGftzZF2Zk/R3BSENZ6Xly
6ZCwfGA3ATCZOUMuw5yvfNbeIYpOJioLSkGCKIeWB7VWj7VJPSXnmkQby80aeLg7
Nui1ORY/+i4WiUWapVPQNsmM+7Sr0B4yoD1V7GOfzWkkOZX4a1xbxlI1kV6fcTya
4fpgW1yOAcXy3aN3YykXWSOJ5NcHGZi5HWQYE/CG4hqpaDCotxJFDyoqvbtAJxKa
sDZoyG4pVjI6UzQqKXQphNi3EniOnQpKpIV6G0gJvJxLZHA3giK9qm5JweY/Zuj/
Ee3XUQ2OtGCoHrr7GAR2dFLjDU1/fing73iVhYsU4FgR8owzmvO1SxvnNfklrFfL
sGijeTgEkWpOWFxZmEhB6HtfTA55ZuBMchonRyF5I5YrjUPv9/rI+iiHPGEtqE9x
eJdBOrGTDGRtnGde8IUzD7TL/8vgzNKlaE2FNbW0Fm5iFAup7dPqKAVQsTRMy4y4
XXoTFuKikw8N2hhfu+wqoS92sjkDqU1/TyKP4p/vtcde6pPDdVTWdE63MH2dAoHr
2QleXlSxjMgH5tlCDocZbU7oah2sSva7aqY8DAxDfVVdF1lIwLgmhLSItvWkHJl6
aWnT/S0x+QIOyNVxQsJ1rnZFycUhe8j5YU+tMqaMymY8FIBLqugwSt8DVCaAgt/F
Lspw5bO83k/KYBXGRrUmv9/0Yn/LWzJIIqwhutRic88YngUZ6gkZmE3TDc4opqOo
TZujrEC4RqGsLgqyRutTguFSerMbK37TAKXfod2oiE3H77vVXj9amoZGQ00x06im
BYB3bU1DWXpWpyQasSqOgAwX7LYHJNvvBc0fLqZXk5c3qYld3QY0KUlq8N+dZrUs
e6p4fIvp0HrQugNGlzoe7E5DE9nNqbyCMA0XH/YBXZmz3KzBq++4F75TFQKVb6sA
u/EUD5Hcx0dYwDhW6IBGHXobYZdgvre1XakdEAux9GHvEK2+EMnG7J+O4Qs6Hbk3
AfyqcEALZFWGt+xR86DIIdDg/R342Ng1qldYgm4DyIVvwb1W5dJTKlOUvvuoyuvU
MLU7/+4FMcVifH11/sCloqL9einxsd2C8LHFriSZQ9LZfBfJfJ2jbQ97pSik5m19
OrRFPj5vl73jCOpe2qrceNjc0h/W02r6jI4DV01qeYaJphEwwHoW7Y1hPDExmLa+
evB5W0yuLJ2y2CWEiNoI6FBVHUMnc1RnWMjQKvj3t0pcoYOmvERPsEhzGAU7gCH0
u5rCJRvIVHidOZ/HQx9GtDKYY7Bh6fNIilItQ5maalVvT80V+K1eTinqY55tW70W
VM0jjGpf2auc9XQuAYz6HlFPYCgcCtLziCyVf/zwCI/gkPtUQn6GzjTL0qm38etr
X127GoqDgAtWjeot2aHMVTGqrdw/yRCnN8ASahL/7Wb0WL4IT4JAAuNErG/Y2npG
G8veeuhAQE4vKaAjIYLzH4b2QImKo9UHmTMuuKtRDHfU69qbatZ3TuSaAmqF8K5D
uzQQGbJSsJvUJn9mnAKgMkI0EXB+e7ihQe3aYOOCblllAzExef6BS+eLB7kPzOAW
7oSkqh5Zq6T/gaZEiqv+HKjmpPIPCoTl3W5KxMULUG3zkXqe1xT2oyclzOn4bp9f
VYurcAkDviy+wXKVwjjw4niil8cRgkPqY/fNQu194b4qM8r9BhhbNwUas22iHDXc
1g1WjQ9uw8BJPmZfqrtpWJqTSHoCBX3pgxXyDLxnOtGeoC+49y9w3+J6DlWZf4Qg
IPjaFC5pOiUvQTEf6X57xTZDElsGkpHmOuAVCGtMm9cPDuHfCplLWHg7OwPhiJHt
i5RCHq6znaeRyl8pBvytRwN1MH23odQV0IZ8IOilvyak49AR98OBKqgoUMn3hjap
IGm5OgaJoFyUcJ7TdPH8z4F6OAIbrS3Mhu67C/SIJzaVuB8q8x8jVRdD589F7aH+
3oaSIadJEEQ4ElBI/kkuFMeXEP9bOsq5EM5d7MfQkaKDyx2qIgnNsSMFsSFibGoK
t5qGQyCFuOYahU3xpesi37/KqIGnX9mWyY/5hnNkTXkhihlD4R9zxVJ6EdF22Ugn
IzRIssj3aHfznzYLfg9H0+30joBCOXSwV+f4/NqnYoO+zH4xMge45Ux6wKn6JzQc
0jbApvSMWVaMtRvlA5uJdrWqRA+jk32OeY35GPRC46TugXjx8SshoWr086rkSHSc
UR2I7fKv7YC4Xfvar5vfe9Z5n/WEJcOwDUQJ/DGFgbSMs/mJaLvOPk0vOBFdVmDj
Td7rjwaZb4q5Iekk/fdusARxdYmt5Uts+EIeIkeyrVbFPbNhG+aEfaVqw3hd2ZwF
Es8dgvEmKtS4vHyKjqiAWRweh7uSBpAodkQo6RzIla50DK003C2Hcjxj0y1KsWVC
ArnhJ9PZgTfnBH0UJqFFIEjdxWblvi/1navUBBhODG5qdfiV/b7Tqg7qvOiZKIgT
zueAG2iTzG92iRcOhJI+E172Jh/MErZ3Oo46li6VrqWc6ZJq+FLhEhsaPy/VWCUj
sCQQwjfaObz1zKotBqQ9watKBFlTTKOaXo372lThLdhb1KF+/KS8YvLW3WiFfNB4
KtMi5cnjS+OsF0g+h+htartRp5bgRgIdUIv7N3utuALcJ1e+IomGu1m1F0zA7946
OiVgAmfsbY77kZBTqkiQNLGp3LSpWJUtNywBoPDgbTfPcDmquILeE6+mqTeDaqwo
vHokyTGuLhgpP4MriBQAVBAR6Rz41+x1eOliXG2SmEwsVd9gaI67R/IU6vS7D5ua
plfCwLtfGYTojNjkFXtvFwnqO/DUfKx06624RqGa2du7gtpN96ePx9bIbRA4tPR0
FFAXPHZFJFoyRrjN2l/RG8OrAaWt1yepQFmALnZhT2XdE7IKjOuyTWNIoh3HoRNf
sKT6vPFFaRNojtNj+FqUBW3VA1dBpaLWjN8ogi7tSKF5lHkomo+pETTvjMznnEfM
rLWS+gGSc/wcZcIJUH53IHT7KXZwVajg1ZH3kY+usOijybbfeS9Ses9cQ4VQ6Mrm
etz/eyDqAgVFgYGH9fPxaKES6ZUM078MBMSFs4hfOf+BbBeJtlENlrZNqReIiBnb
/zXc/IIag8ufiiGNfMp9mcAuRhPeV7jsNXio9zZIJyi2BfHNsxGcK1aqglpn+kut
6I9HPqvvZpMGTlH961g8SIKjmGBbev/lqgQundryePw0XjLdAYB/5VHSZsIHuFAs
SUwngmTKmQrsrxx8Z+3/zzcYQIUcWR3WeFTjIf/k8zXyZbCU6vFQ9mBzxtMXP/sG
MUZALu78r3Dy6qj0/MIlJwE6uWwEZ2cQn2Tk0Sk2hmF7qCIe+BvfOSPQmca/B8Rq
pWPh9si2rARiKnM+mmxPm+VSovudyrhFE2/Y4sRcOqo0zwDjuBPqBSh+1RmjNDwh
zK/rMI8KSw+BYoQGZqoD1PJYrKKoZb69ejMv+A4jaWucdSZIEi2ZIfNbjZ15s35r
rFV2QCFxyMPQ/SzMIyrIoEBbabKhA5/TIprLjO4VEYKtJOBpo0Uv3PZyq8Gzx4Yz
VHU5ztUbbl9mvMU2lBrOlyR1Yzhf3oXiXGKP05FyzHKkJ/02DHeJepX2yBtNOksv
MzQyQp/zE5MMMPDhYktseNtWAyKl2GdGpa3xljx9SGvkHEFWhbXLcR/4vlJZ4u7P
hC+Nlk1Dy24305O9OPyj34Lbuhi7DOsjDqr5MczIGZU/wQPaw35DRU4UJRpWZjjy
jTg/qOfyStN6IyzDWmzWzLO5y7LDxUkAZ4YC1sVAHUge/NwGavDQYqlLNBn7Hq1J
VtDeSeJYhcrudXR1fop/21JcrxBJZ5y5l+SYvf3NWKccu0/Fco/6GoFeWuVkRQnD
yHMJagXCcz4UP94PGOKqy2jXpYsEWK5waskR4cV9Ix5gPv7N/IK1/sR7E64Itp3P
7nrmOkOKQwJEUx8cA4hQ63M+cj/zr4D/z48wezbDNuhxJvWP5a6N/MGEryu0eb75
FWbsb0CrnZIRv1A9+LR/cZHmWcj+gVPvUjmxl/vAqx9LfzWGTDzlM+isKo4PVI4p
vVuixZqedrC9ZG3Qs3fsPDja0Y3Jy83uEiMepxtmb67pbJp0IX2QU7/WUoxY1w/a
W6MW26DtpkGIn2Dpd14497khViXcnTLZuNQvGyMyOq0RxMg9gXMHSUT8ceNKwmbv
xg+nUP0fP23uWogFbLexXwYcNAtA2PZdmceeFD5WTIevINXHGlBPQQ2zJ+NjlRF7
qfKEc5x1WBI3guuW/cW7XdBHr2FxEukqQa8ORnlvrqGs7/C2d7owWZ82MtU7gXR/
mfmmY2nSpBzulxligFbPsQtSQb4bmNWUarkC6AoMuV0dKpLvWuH/WW/Hj/OOxdNe
I8uNH1Lk+2hz5Yc0RYgJfnyygDiVXgl058c6q/dt/PTBJd3YKRa6EzylTLCdvrw9
iKGqPnU3FSRIm7K0h0tCbYIepALDM2xah70yR1NUldJwBd8f6I23PaB26PuHfZgO
7m+kG2uyEY87gy3uBaJscja5pjK+gwo4SF5gD2kh8ajHYhMN5OqVxPbaomS+PhpR
AW315gd+mbsXYEz+YpoSFMdS93tQkt789t7qHqPl/D4sBltgM17rGKCiYPIJzn19
SKtukjI8nTZX9JdUB1n7rUcaWfvfm+BiR2A/lX9SwXY38Jws2IlYpuWU3eIJhlZa
tNiiegl6CmhfBJnfINCX4vI5urQJaSjSEHfuS8DRaao7QU9WRgfsXyWRba8Ltkrx
pLVcpqZfE6mIoOGa4ougRTxWem4ac4zE6zW39ZRXjtq3/nilDrZ/2xuUwArYChSg
aicjyDqXI8G7ezbgsuSzrVaoDVI08kRlMT7MrtqYBRTr5RWwEllIO+gQTQvnuAge
NCF15mk3Ea40iZEjccIwtqdOFWiM3B2L09joNQEOmtG4ovi1vYpc2/ptTzj/alnU
vROzLPARkSl2wsGxZLrcWg84H9As1hZwJfLT/U+DOaqfciVGIBeDO1PGHsFDGjz9
Uyu3SPXbv4Cq9BYOdg6nN9PTR/JCBuPrZ/IueF9zj4xw99kk6GnxDfLt72QUq8z4
eLDtE2may8nH5y3RV2bfT5s+mHFxf0B2BbvPG8FICQLdh8YRQ6t33gMQt3VVWlaX
MPbNtt3ERulPs1E/KScfJ0qkCbS8WZIVaJhWgDELMoSPUBjwfHbpfZXiKGK9pOWV
7ZfzKjQVRt8JHAAM8eC4gA8D6Cta/wXZcIU6ikQ9S0hngl1pdBgcEND7/zL1wC5Z
nhy/H6I7B+rOpKGgNWgTBASd4hyt2OCjMI0Ow9p01D5m8bQkiczODY/t+2QQdh/z
Fh0p8wY0zygS7lNgneNvvjFsS0nnmXqPxrFFhZyKR3bOj5Mf5iT2tqOax3ZCevwO
d5a09X5cP7xJJM5H0GcqaEFRpI+cx+p6CHZgt5FlWWZzOS42Wdn54aPpG+wSK6KB
CCSUPqWJycN2wXtznTF5D+0cfuOjhep5kHJAohu0wvqVGUtuspdQ6D+fSuPGXvMX
k2fOHKdRard4nu8t/0VvhFQC9nFIr290/Jx49eSbvW4FzC4q/xe9Meix7sZOJdG2
Og2hnm7V9ZoxSwwi3rLfYueUGuJOikGCE3Ap1zA73ufAZDvWbIDsXCB5o7jtZnGY
BxhfjAHn6xxkYYPEqYkOOckCZnqMiXnktGDjGIhCpsxs/6dAspyfw+6aW29B6Osq
38bYdzanhmf2O/kTD/BXedwkO2h/gbLiwvYX5SQu/FOzkaV62q4oryBzsZs++LZS
SMUmmFeQ7vdGXScp2kk8FK7W291Ntt5ULltPnhv2rw9ax5qS4MKyL4xyD0vOCOgg
7lPdWr1mT9Wi7ba3v2HxLDXqkIlrjBJ2j2Nkpgd4YXjrTKzKvtahlILNxkJlBc67
s4mpHn55Z/0SB/Ue77nBeJOkiovdpbr5A2NSGjPUmQIK4mDXZu7yGxI+Mt7v02Nu
TqNmwHaqOleOtuDhjZ6B2ZFfBpeuTBfwKGY4Jz4keWTr2jJygmHoiQBPsFVqejmI
+9PBU1Jx7A58urXm/D9/FRYw03tH/8d7TiBQVyxvOmfaBTp5m5mSPMga2ghe6I0W
bldJPygvH5Xzgxm+vBUupiHrEETTQY6bIShs2xDGrkVOSjhvv7XO+tFvr4PmSlVm
ggqcEQKu+pAYaWgtIywZQcm2FlziDnSGCI4R1xXAKlM1ySW4ehmgrsNA9qArg3vB
3hEP0ltZzVbT7thlXqzfJghw2DTPLCIcK+vjrSbHlI/BoY/Ag4CCfHqmtQy9vqWr
Cg1tajBkqdYpMcMhqKs+GXSn+GojHoKi3d2P3kxw8PRWCzYn6CtLFB6EHLSIoSTy
GLykfTJyU4uEiZsZQfrR1Pn1XhNVRS25KIXsCdxkTIX2VCiyAaZxSkPHwmIQdt0E
wvf47vkHDcpK/ZabVWEMf4FDSpsyJU9mRr/ZzCQADbINDzzZ4/jEttUPLkcT/TeU
6XYgrWd/BI0QZBH/iTI7lrEo7OczR0jG+MoDlcfymnbsNdRdLKKVgkjrJtUEUu9E
cDfRBCNmPFEo5ic7T8V9ZXcY755yOdvD197UPMf6wZjoSj0oEBTN+ApinAJ0wnnh
PpnSoLgcE2VOr43wXdedPXzDGVtaUun4XvmS7wrRDevqvLvWA9q2nwitkuPT2u9T
yHTPmv8fprWcrstG/Vqt/0+rH750eADBQoPh5NQNH2CkpLJbx66uVbkpiYvfJrFk
bJ+YBdBq/p8M14kZoSwnkUbxNfHYfUP8Cp9NQGUFRrKM6PrzbPoK1iBWwX0yNZ8k
//ijtMOT2529q59CmHhtZSfrEB/S6nocQXqVWP7YgDbHSN5Ve4gxhE1ZiJXTAHhq
jBGF5EPZy9Ufc1U7IyJvrTJNBZsnRPZ4jO3ttEhkMwwTYDkzBO2/9o39AvvKMLee
dIXeH/4nM0jB+OJecf3ZSrL/hGWJvBE1iRxo/WmFt9MxHaY+5iJoDXlfZfRBYTOK
dVYc0FTsGsONs/yeeAuYgnCLju+Ktk7a+3DodHy3AXAOeBpDSbyS8/E0TiLstEp0
bpVPu/rj7WgKlZOV+tn0WsTYIb3goPcqmRAVaNa50ule4UTGRpidIzfUmYF2bOpe
cBiT/+dCrtaTNrE2etE99t4b/5XsfBLGfE6xAQeB+XS7zpccE1/myWseoTGHgt/J
j1lK2Er3Zfh4vwxzBu6lrPLcV8I4NnmFYNyyBirraC+2uLMKN13dtWFhAYpDE1JJ
ruLahAqsSuxZuE7nj9GyMMPXWQEnIH2eYn6a7PDHmiBtq33QLGdpFSeOY3BiTGdo
umhxMNZ/188g/6aWD1227z7/DxfP3RbdZjU/oh3LlO3B4PGYl4ujL0DgeuEefALa
`protect end_protected