`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10368 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
Ju3IpcJpVj/VshHyynUPTG7kN5gTlvLnmXIUJKrchuK1OxzQ4c0/CUTLSKUrnTxt
0LhiTpma2HaYPPVNOkjQMTMj242ulu3p/xKN8H7YUDr+9lA6ZMKLuujzF8b6y5So
cTn09VI3m/piOWs9O+vVuKJt1OI14cJD8WqdsJ2XaUThLdD5JKYy7N4GKWNbUNj4
YYErfiLQt0LWRAdtHXpCft0AgEPhW8MV8P9gCNLbmRRLvtBF0vC3Q6tNfFtMjTEP
+vyyoiIXvEJlCfV3MGHScG1tx621l+ECYCg8qXRG6eDMkugEdEcatqwUlf8EvDsQ
HAWmpneUWiRFZ5wf5ZKDTu0rG1IswE88rVN68MGvDIN0ZYrOcoP8gEC2Yt2iQu5d
FIjOBmxugzprAJpNz/0GAADZWakuVtSLbpKEVXH2R9R6xmnOSZ56KKbJ1Mzbcm5A
fZdWWM1pEAp3jKyr1UZN4r37VE5yMIEm1MpoK2JToqvp+HN5yG03vLHuLgRwK1ab
9QEQIVhTw7qFSVM46RIRCBrdUBEtbhRlS0W97a3z8LYDyzfRCEu54KlIDtbyGKPi
vdcMmbsp3O9nVaw2B03axV7vdXJNfMR5WHl//cuwIBMFl/ctZ6FzAWnrWvIDKbPm
AQttH5jFljfWY0lBn+R3ay5dOBQabjvtdrKPr37exWNw+0Xz8TIxRB9FZLTTHya1
EYAfLk1pGy1vIHtQKSl5YGA6oi4iDWfVtQ2rKCyAoOhlwBoU2VxYCL6/T7ZmuN+d
R7yIb9tHmKhPXkDibvtQXivI3maiA0qO1I0fPFbcBDKOM8o0VB/sOzA6NzCZNCbY
zhP+kDDLm3Wk0i00go1AL8ZVHCjDTM8Il7mU8z3ZH0dsuyXMYKzjJio6w3AWO3BE
mBebdNa4v/xvVWzu89zs5lBAZ3SCOkBqtloXeYqmIR7LVBzn9LScl+sru/xBJq2S
KQ3lVk5VPwgZbJhi3WklpQao3unNiO32wownI+uBxA8vdNdcD7B0bOAmmGYqIOdv
kSRlPs0mAmDRWYEGP4OG8czT337PW4+iVO8mknnd8y9HYuXODCDwEuFVM+LAo2VH
CmmrRuY1GlgITggeuo2VaFH7TbZZsVacqfX6yiNUZ9oI609YAAgBMM0hZx3fjYQB
boRVnBPMdosnDqK89l84+xUE5idpJtf/v8J+jEoZxJOroFg9PiB0DeogckBIjlFD
NALiNebYIukeWwd2CoNzTCA8HD+2ymLpd4GVrTJfZqipzyC1PPDOUf/glS+/WO6r
KDLQ9bb9vUQ0kWsqBC1wTRTraLnreqznVaIW7QJ9m/DSiI+bO7gGY1YUO2oTc5gy
TL+84zvyRdoZqzN4MpjlYJgMp16RxAuQKoqhsgxXTMKXpe1lnCAwbhZCYtzigm0G
C9lrroNWQGnsW7B7D+v2E6XZtv6yMRj3bimzHdQYslYpeUb97Pe+XUdsF97iA4bq
xo94DFbF1+whThrChgbv3ol0wY4piKjJ03zMNWfgOAYxSGz5Bs/FKs8bv2IxQtbK
lS/YYrHpJUftAXmFp20ncGB/8Ee3Dtg0YxeQ61yDYR6a9ObQOh74S40FTAvynTmh
UosBozEvkSFcrUwvIB5Zhsd8wYMm3QzAjTP7GezSqwOhbmUwXjWgwAGlc8FS/Bzo
t0fMZCVuC8XpAQ/Wao7Y3GFwcoqlFn6fHfHPSwVzcijC0JUOEm1DY2TctyOxGWQx
xaFF/2m8axgSBIY54qv02QNXcp1z2AN78WM0LZVLw8RwUUHQEVJ389iUJ0OziyVt
+uK2g1Fhv860QWkUyB2VjyXUYvWRuZINN9o+9DobOvVwNgLMksbN/n6imwbc+O5U
O9NtZ77Uvq6KdcxSsVGEMRR7RdYS+GjRC9ccSHv7UFAFM/xaCmHybj0yX7OdaJ4t
7ved2InF8RRXyAJqYFLVpmpwiAAOcz1dx/SV8IsgrI6k0NlGlQ9sRyZgw9TkI0oB
WASScLBv4Dna02eAHY4ZGGkYUCzQSx8Tv+x8meqA83JPoYd7TJpY3ogG67oOXzOF
nArnyMfjHhu6s+T/yOhgf7erRKNqssLEcZCergPuz0JJBa7nG/GnDR4+nxLxkrrC
swsw1UjAhNU6ePnSJMhJnhDatZWnq6EUV+B4FiPa/oB8vdTFhBiHeI7kXlNUMuh0
r+D3FuVXrjDL7cV86XJxGaMNR/+WTHDt4ut+rDA+yfgRYskr6AvCCBRLQJ8lIQg+
MDRk5uZsqMbCj1kGZVwqAvkxHjbXx9UK0HPkaU+4Oy9dubxKXU/DTqzCD5b5xnLj
5xuZ/QNVL+DtlcRMvXclCVALhLwuPr08cNfiWSEE5CM8P4rmoM+WkluxvKh+6GcQ
ZMIt6HAVJXDEAqjD4j4lwqVU4QgAbnO8ui18JcBO9kAPvDI7mISWC6Vmst6GluNk
jtnx7MtD4erQakHKtTv6QJaXBCV9pmzB+r4jJZ+53jrMw7xf0wJqMfre2Vd0Ychq
6rVlqR0AHmDcKoWhZPvi85GCLqLCpvXzLyGWT4hJ8BJY1U0aNSjj07f0NIv2GuS1
BmxGEU4jOYtflHYK5u93EEirqpq0CdlTi6duPrw9iQWOkHaW+bOQbdyhXSgxtNBZ
Rz2FyKA8kcWuhaSRsGNzZRIkXOBYxPwOV5v09+3UingayOYbXZgenmZOYCx9cauR
kcIH6fb8+5vfBnkZ8ekiO35sOYWIz/Fr/TYEDT+6B8zbtnEBDdFkuKqsvYVUV7Zk
ez89MStxRe+VIvk1Nw+Hvx4fSAYP8f0zNWepulVPuNHLDoKWSmbCes9GqshDeFW+
a8le4ERDBL8KdX94fiPdljRjlkYQf6Z001l41h73NJ35lyRap+qkznH1nHJDzN2d
8eNX3BrCsH63muU3fGffCmawHa/OC+1iPoi0OKwy3hAU+h9VnzpQMCQNl3PBEeVh
kk+/oJrrFwKQYJnPUIaPxqZ2nGnd9P44oB1vem7HwO8MDJ1YUkCBVxXUxMH6fuRd
7WrkHtsSzHWZbaSyUl+3KWdK+6EjLmrdJtnZFXdPgxOXwzTS45/jZaxADWV3+2Qk
bf9JI5YFCqCzCxFZ/WnYArG6/+mjQ7Y+uj/C8OsO7ezyzsqKauiCARuSYsyUz5wY
sCyvn9wQMWa+lPBrJvIYjMfMTRtjC+bd2MhQCLUUzfj8rFpcHLs8ABlJCOtWvuTA
jQ6KeQ/Xp+rqs1dxZIAjhpGoybXNvq/AyXfYxDDa9qBO8hADWgBDSgHp38Nw7iK5
zPAg6UJpguB6/Pi5qEUS7MCttc5UVilq8YT9KmxLzkVpiRrNtzNyrsNn4ZHBtw5r
2pfzcSVByi337jzJiOMS0fRAK3xUj66Kmyky8Yap8aJ8JCP0u2f1a0/Xa3iE0Dzl
YtvtwP4h3ip5GEfIy7yBfwroEMbUbDQY1uXv20ecUGb+YxL4rA+aqh4dMEcmBSVR
XLkuWZtRjQgPn5fdV7LS+kEEySgTk+2NKw6ZBhKoDX8+VCsz4t6xd7uvUV5Pf7QY
N+/rlahtYJOXZfLmjhf85wnEXdtPrwAM39MghxTmFcIcrHnHHawl46UpBIo6yYID
BXtH4eTEB6PSGZEvhcsJr1Uj+NyvBNLx4sZi0Xh03YuajJBWOJLvMqSemtgZwQMG
egBHZzPJUIaFavdE/N5JhnBcTOL5dYEffdKbP3FVVI3WgRXwhCl+taqLjPd9IFNI
2gBLmyKwUna6oQ+NZ8X3LkwBMPWxJvDZX86XUyFnWtbDAsYx0IcagDsNVdVNYNoh
X/TKCtmnLo7BWGJVBRd5J6IljHvmRz3uwZxdboJAXdxZYpLztMPm3AkqbDdYfgsp
dA4jWJvwVy/+BqrVoYdZxoARrUQDunbM6Un9TbX4J3OiyRumS4mjsZw/kyQDUE5K
MsGZPBaroer+ZJRytoTy8SiCZSAzkZCEtZjiiYNDWo40gkxFzWzQmrdxWwylkwXD
kdSgCYATryTj1NSp9e+DSdfYMLbqjqJpepvPoWR+zAUu+NA1IxAuugKaq3JNLWrB
oWa/hQmzwg4vPoWm583BhF1kK/Mnz8DqAg5YSve8riisReiUvCxpUTTMFNK0ZemZ
C73HVU0TUMgFDrqT69iMosnOqe2Z1Nxwasxnn8BZ/YWQfGkY8QxeafG8s0zreInd
+X3W/F9eMSXEI0BKKxRmaTIquUji553EZM1OdOOsIre59WGtVbHxwfijBqb54Y2q
PXBC0Vbv2rwyCpymOPHQxICKMOqWZ6Gxu3REMhTr+s8AtLj+b9orIBQqBaqGDL3B
Qjobe6tBCYqffmN5tZNFt5IA0tk/O7dLfdwh1hNAoitHKPsBsdNFQNBCJZiRn/ZV
dG/G113SIOLNNRhZ4loEcBPv1HR3QQV9LF6MLqmudw8bq6zNty1FrGFkuiJYs+dN
98or5tnriVCC1gNlSesdhvA9Y6cKVEO6nZRK+pNIbyw4EI77zRO+3dVfGqnGNWEo
LSBK0PwOxrZT+XPUOeb1zHUsshgcrmn5X9eXptCQxya8BjO6PlBfe5zpdRDolXm2
qcJxj4Hd9Q/WLFkQBJAokN798SG9Py4UUMnaRAQbTNmUgGzqpAQUMufTfSxjNcV0
Hl91nIXLjgLMpD8hlI1D4Xs30g3IE432wt06tk4Y9GQ/9JEgFSkQxw8vFyfR4C37
zKHA9msdq6g68n3lu3ycqn8NHkj/RDREBJgPVmsehyDZMb6ARcxYgv6E9MObDSTe
wrnIHHV7Pq0TG+ZAZNp6EGpVUmmmNRH+g4KfsHaNkhe/vIwh9BNV6cDbZGa7rvlt
Y3uQiqSVFCfHjCC+5tjzxRbCOovnMBeQaqq/mg9z44/Cec8EDomoKStwa4kQ9/8O
FCzx4SNFr2QHk4Riuf6WD7C8OSPfppKVKRRo0JPwYMnwJUc01nH0KQ9wcrziuVgX
yGyihXkVpSuDux04I5tyxyjSODJX/ThAhPmwu+9WBlhaTPm+1R1sq/67Mhl7tT8y
anjphKEHeUSVGVWUJ8XxXnpkLo633sCSMFV5+jW/biPExFR5mTYAbWqrUCuxutgQ
q9imQcI4fjuXy7hjEEgSDqSqUZnhUClPuFwAYKziivgrCBjZZxfQiurxSOoTO94F
VwYN8t4fS1CXQP3OhnzEKyzPh+OmthKNKImDxScgzgBGWg05PIYRyEhtkkk/DwS4
sVQVqseKhJoXEBzHK9dX4q4H8hh1x92N9RTLdhS2IbwWclzEfWlV9JEEF7jcNWOX
jIVe4UBgEO3oiEIiiNhCOvXLG04w/dY/oKqd0ZCQd7iyOguBfvFH3u+W/O0n+bxp
v+hqtpZEYAMEUjb0Lu71YWz8OzzUGkV+vkDuGqYEZvcwn3pD4fJ1+9EHJlJDzmjQ
PqrkmWltTV/SKv8is8qOjTsR3GXNCbsi0X51VWEpmZ4sXlpUspp1MtcTHrXw2Dl1
OCMfjwH5dpZzGwAc9rARQ5xQ7nCUJrSsgGy4Rs0qKhADdCNHF7DPHnWrd1qOXjEp
Iako1GgegB0tny6gTPVVqMbXl3bdfKndzpYqZU7TPmJkILLBpxvvmVLzfGy+e57V
Reu0FN74RlHu1FlVToI2F3DrZ8vY+I5S/3jZ/H37PSHYfYoaekjUwpEdYmzYRjX/
kaRg2qEo1Rthp+cEqvoGYKMn9c3qJPAlz1AYk104wKBXgyuH/MlxPRyWwbXZzrpP
nPLmDOcLbVE7JlbCd7pcy7q97sa+J3zMG5uc0aNMIk/DpaMUmS24he3aGJ9Bur2S
jCYVnDHg1KWrVeoBnNHXiBULC3zZX9hrwKhM/8uz/wIIa/NOBEftTeBeMt2Uf2Fi
pnEtNRDMV3xEpap8RFpzxutVuuYcrEk0/8XNBG1opY1eygni2KPznmmV+TlhTMYb
dAUfLYfPVHCC64swjNNzW65AasfpdeD+7mKE2Y4zJy7gJGsiZNTg9gr7T1zq8Tsg
uNn+rXN2mu0koS9eeUqMvl20QLwnDj2mjtwa4n8edbnbxZUNwAQ090g7RZ/mkbaw
D7ypuNVT+Sh9IgL+VvagYlGWv3zHvDMbdzWWd6p2mnaxqDlFNVArwApONoTg544t
IJiW2Vk1x/eP8/RHAEGlmK7MHgswKOFH/w/JYHP8INZ4BicKOVWST4aQsDVRDY2F
vRl8lTbT9MeR6pujopbuF1j886ivkSof2ukLh+A+pJJC0tg0QjS6hTKrHV3ZKvVX
4hcwefvcOyBa27pwG08FDFOS5lXpQw2j8WxDU/JcCKRpH518gDSIQeuMrfyYSSYU
tZBG3a6XOZxnpriUD0Pv45/3lWvXWV5MV0Akg+932CzQXNSUsR78Wjs3/Z5g6H50
HTgefwMC2+0xa7mYE9qliISUPm8Ve2e3LYiaBowaYrfSyxDsb8fZ7KBZxANdQ2fC
87vq8pMt4sfLyfjijDDMPcFdVxvFT31LjOj/zVLjU6hsm1XQOCp6x7CSpbcmp612
7E5Wl7IyABEfXblTwtpa8jkvceCq3N0PD8VwIosJ0Vk7NIgmnSZMx8PZ63o2exyH
/soVhTGteTnWo9MymFjpWpe8rF0gcj4noYXaVTZn3VIxsArAfodauuIeEyHydbB9
hs/H6TlZfzwRH8iL8Rcwj+2570U4NomhAU644/HJJzZVGQbM/iX4Bs1QN2ltMCaR
ELc0p5dYUTiFdzrpYf8wb/Zh7+EVWT2wqD//76fO5R/jeFfkUUV+v3kQLQS3aRNW
yoRqvk2K2P6EKPxChqGfFppy/1lv+TR51doPK6kZLK59cmb0qOcnRj5ZbRDGCxIQ
ZzLSMaBwCo1BAD80G3emdeOR300YqYeAx3Xp79ve379gQ+1dCpvaABwg9VIGL1Vz
OHGmqPWbaYnZywIQ/twmMicr/y0yTOYlugJ2iQqW57ugl21ybCf9YTIwO+ByNNeN
mbzfzAtyk9zzE/KqSnQUEzJj/awUaCIQncf1FXgZmVUsN5+wEKWZY/hMsgIFEKo7
O6FxsOrzLFACr+Mxo9caC6Quj3VXLu5z1X8k6LUBQTxWGRXGE7B1WGRJqySbwFnw
pe2+RR/zBh8hnwMXoOs29KP/is2eCM+NanCUZAv4v3/vx4oJwGVJDVg/nsaGq34I
belOPvrdak8s+64Dvd7b+ZHmSGQTrDhKmFWCNNWdU6I90jePG47ki7B7JE2WhcBn
w+RB2X7P/AzBMhn6hO9yqAH6TER80TRMLKKG2NiCLmPS44rR3IvAMUbP65iHkg/z
lBM+9RVVgvwX38WYJWpc5OY3mpYGgiwNT3qfbnb9o20l4RvFA7X6UjwSTpXD3yuC
gzX05jNFxuLnHaCL6VbouF0MYkivZWUvjdEBey25AXkV70x/WBRHhrIn1XLe2po9
Wxn4RcGfs+XQQbVE6nSc/RF62I+bhkvxyaBuBubv8PEcaasRTU1nfCDg+ab+u7Zw
B6z7fs30dApv0GyXtZ9pNQWG9iwE9SZdGaS2STO9ebDHUUuVYeKalW3JY9/o//X8
jwMtJtTwAKtCrSyoIEolh8BCV0oGkiWb/mskawHazo6+37gpWgAHOuHdSl/Mubf8
X/AuNCMrLG3IW2dabTI3xvN6FGPkmPwaFrexyL3eeDix9bc9xhbJYbiW28pjtTdV
jEMmc/L2MypI5Ga5FPFJwNhn1JlQN3VP5VBOzB9N5ylMhwQJJK3SrLLhGvKIIEcD
d+3EPpXGogJvXSj7eSa8rzizL6KZzKAUXsjAQzpg7FpnyLv2RzMkVQ2N0S7N6a6u
poyufQqK4HvlipBU4cAmoUEoIEOg/kH9J2JE4h7m0qhIjjJTHoTuekFYC9SEGpn1
V6XQsJxLKiL5ja9gNOW5VJGxkY1YMvSB1DJzG+0DZMcA7WzoLDCHpVIfhAoGTzOF
yybkUmxGylDJfioB8wsGE2mUwdlAv42LtQHxXBdB0qPAujlSmhDo+QOjSVPKAN+p
XkyS6902r4O3WvWyVaqFD7IJU4qoBs3zSLoFp+L6LtJe6ug2HP+nS6yMk00H1YT9
kFGuU0z3nDZPL1upi6hHKjq9uoMhZDaFO9A+sSEPitinTPCj65BKnRBfuO9+0me3
vFibUPlkqTFSBQ++we4zyCoex9Ox/0mNWPgUkKeoNWCtjT0VpyOvGGi2YZAV5mwo
vpPv1sA4TcN/aG4IEm661lLyg+53IBlxoU7wPvp43lyLc5EB/YUZ+IfrFNXKBOck
Pfcs1SCWJ+CLmPEJPPfGlaSuVKdWIEUqHot0ZIb9Nuih2zAt0us1hItt/uhWpFtF
0vf7GhRqGVqFbXpedo+S+Y7tiovrpw9q70XahpDEAJr/u66b8Mfi1znNquJx4Z1T
82eqGd7Fnb/MXBvJaj79STVju0n2lI6Ao/2XcCIIMM+9afRV2KMQ5VBl+qIv9lOy
+Pu2dlOhFI9iRRWQJX55XnjtcyY6h2iJZ17PVloGilyPmv8x8dNRqLMNkv4hrCCy
Q5wNiiGETlsaajnmpY1fI2wFbmh407pBRuUULolW837bdnyxsVSj96m0YHSThii2
GhdQBbMYl2Yx8DT6f+RpMeb9W41uBrCI5ZwuOwv1r3irqiKln1WhBTCmo7p21D+k
2t7fMNFfAUQi5q4q7Xv/xJ+aG9l3x0zjRH5yyUemyPDHb9otckfRKEq6esLYQ5bS
QmhDDtDrijX2B/30UALJKHanFGuSbwofbxYtAlxPDKefFap4yxoOoHE/htoHFzJF
6yd5cCaeXfyjafasYHuAtXs0BMxnxGkkKelH2dr1c4gswQRjiKMwqvWcWVksDZB5
asvYbOoLfJUAJ5zGQkj1nlvXoyTAkszZSsxL/mywFcPOkvM/Je4AM7DL188okog0
9RqF+y5W6cdw2xnxUNStigFZXlivQWyGrcjrYNgS3qMhxeWL/BPsN3eTxiYgu8If
VUoDUvvO1H5DwCWK9SVrSRSs2Fkr4oSbPw/Zicfn9QW/RtR52DASTGMH0hBpwLkc
T7ttVlQNSKt10MaLtfJrXIYuTV6MIxUXH4AOOwlNsGcdNLKmvlmw+cm6VKc/JqJj
/6E9UBDQ/XDJIyvkx5ZAZvDnq8u6R4VMdtOp5oMApwL4S/pXDSkJm6Au6vwvovsC
gc9xOkbADS5EBD1yAhlm6xc9cFWPu69dXAQxsdeyrdo88gdvTh9Z3LpzflqeIYRr
PG7ovfRZEGZdgvb/SRwNqasjubrmwAi5yS+hXFmtnKowkmRz0yK5IEYJM//vqKxS
7NOXxh5SzC+lXUk8AAhfwXbN1PyY5U5i2fawKFf70v3UwwOxPcg/HsJzg4FltQ7w
ngSBOH0kJwxSit27OfXsYYX80GplKlcib/Tv6HMjmHyUkrefhgdOOnrIKaqRotW7
FVOUBQkQBP20ZPvAtAHVEmnlqczGM09qhr35LGcBCGzElgyJz0m07UZwqj4YOqz3
jr6NFUQ169dHR80Y8iLpoi3Fwnv76JtqDF7/nbfMHqfPkFynLr8353vF5kS1ii4X
gFsBb3HZyN89y5gAQdBh2N2V3T9fXvwuqWeuBFIUA4UnHUfKkB1qNkKwQWVINeXq
iN00Ozwq4ho44+7NXqjMwP5CgVt4ICnmPbNr7AEzo5mpwf2DoZv1M16rDnf68mI8
3TbtIFLwnrhWdOhkwmM5fFZ4ri5RWAtKrjPQdBsDfcSLQFg3UBdY0DYFRqBTp4p8
vWBS5GwXWVKlpL2teQ7LMlF+g0/01xUfR4oy3+pgPUxWmfcmD+5/N33kwfhvHVck
JEIU0gGY1n+UwBnkUW/MRNLzJ4tDDcf5wIKBkiO+L3Mg2AO3NTHnrddXq119yHOv
kwgKq93reNzKm5/6kAmCOc30/3stwpXB7KVdiUYoDbKRI/2XWmZedDlbcx7uiuH0
dbmzXR43Lna43qD0sMUlQMpRtvSv66AbyXTNKmyijQQhgdKjPzebpOzVq3EwvPEh
bMM+Y5LCnRt6dhm9ypFqsdZg5eXKbdckDuygYny62omOnIrtBzhini2p0c8G44fv
45bpaMm9ZtwUpuv0WKpyz7UU+RC32v133BLXSZ82ZexFVozyb4LBKeEyAV1rxop4
nfDewdOEmr+XvJkUpUrKOVG0uL9JV+Ygt0m4BJWsVkVMrQx7ncM3BFt6eqOp2RcN
pf/Pn93sslwXereKL9rCCtiwalOzfj9kboIdT8SAr/quO9+i1p+nKkrpxCdXVD47
AK0BWVK0qVxGvtRGEw/vaHM+6GKRAAh7FDSr2KTxDdyaSmZW+05ZG5ux8vsF/xVP
utrSRQa3T8Na61atTxed//t9VuPTmxbW38DxLwXVvEqhwd3wm7xzToPK24phGLmq
95EHAbiGLVl0O3yrN94m1+Um2es/Em/ksvur3KKJfhWuYBHbRD8EU5aRajCxVt1B
/He1JILawvVPyCs4Xv/hOx22TISM6asPpOGKMsqZXc3S7cCQZUe7sei4KlUXaUtw
kV9w+B4JcnE57W0Osxg61QFoWNRI+gWK8FLm4XQkis7ECYZHnGGLKDNMUTmcoDYq
h3t0uaW8kdSWCdwmgq2xh9L/egt/RgUwnTCsJCylgC+XGjT8z+CU55B7vM42KSbi
xt9AVDrWGcfFVuZo0KsLtw/5W9gvfJ9hhlqAd41u5/Z9ZfI+9b2wIM8OHR4ssocK
2y512zVuMjnSqGdSXtye3OnNbXo7haQJro29l8k4FOCCS0Viys/vrqb68/4e//5B
GrXgEEg2YqzAdcA6uDH7B/nZ7pHuAez7vNB6UtA2OcLASSt+bvM/A4Nuk6N6iwsK
RItvUZCuKc1LA6EDUvdFC+wRmOpo+nJmDJZZtNvJQ9IhgYPlXjOSXqOJJSufwJiy
va+vKvypMrID7Msp0bZrLfxd35EGLsctjJWZ0TEq7RrDFmngp2mB5Nbt1mBbtU1M
CQ4K3E8uETYO4veJJnIZim4dH33+EmxTfSY8Ywew21v37hy61zdBsJGJsAXzOspZ
t1rYR6Slcy2kNrpUnQVYogbjdX4L6RAl3Q5Dh0c4hG66pLG8ICkOI+J69p7MRVDz
lrmYD2ufPmjfvVQ3p+BZPgkofJOADCk2gpQD2MDDwD3jDgJSLLTV5s/INPhXfuD6
xBrUQvV7EnGMa6/aIdFvpT5EZDWNgGjrVOdoyVs7VxNbz+QF9Vwz8/bNz12P19ww
8XKYD9Ftta7YWu6anjedjkftKskJwZjYCmf4KbhB1h39K3fDlWhkUADFLdcFuF/G
m8SBN02NlFGU9SWd4c5J0oibpoFdHML0p+jFM1QHX0h8qtE9H3sIWLaSx5uNEoaH
tkgFMFDRpVozXqOlGyyjGYdeC+UVuSzjbRPPh04+3cMGLL4EbWO4sgjgLRoK+31Q
WWY/gqUPpTN7ThbPqUdcRqav5lS+pFL50cQiJ6s2kwebTPPS2AUfkskT2NS4SB1S
E7E6FXwLzpJnitr38dzCvRyAQXSNpwOSK2S/qay1n81xyAa/wqKksAzqMXt6q8jf
fNhQSO7gRZq1oTIeOVtMg9Ft7UxupAnmnoErqD/Y/Iej1jegsUWg5/MbTL6aiaLl
z7thiQmlt98qAv6Axb0hH435jV0E0HQxWlJ46uChHCQNYeulZSY4lqSM/lvlQwIp
+nsPSlOT9E/2lxHEy/IiqpiL9tmCk5b6+IDzkTlrSFuqUDO2v/mVWXqI82nTYWjy
rq7ruhx/3hDmMdhGJSZu27XicpcDRj8w2DSW90sjguwYZKS7amcxgmZKIy0rdEPu
gpC6DfBjbFz6ST/OFWf56v1WArZ3I2UMMZK6FDlKj5HlPqw1HBWnzrvWd0tJQKOr
mZ73oeuxzpNhj9wDJcRilco1yFLIpknl/x11Set/XA/CZRer+LRpVWbjX7G8m4Xt
78DYM7AdQZijXH1dLS6ptkRPg6Y3qOMpk528Mf5ytFKCxhoT2LqzBfq63LlXBrH0
hd5BrLlae2n2/xgq2o3pwLuiLQX7WnsGRvS3HQNW+h+Lgq/OPtF8HwVhkVaSRnzT
yXW+tLjmErNXculYyKq2h60GV9QMIcJAJrkE4Iw1m50P7RA3YdHwkhPoZMGMIEh9
OJy+RhB5h3blNyGNKvL8yfNG0Pgwh1IVAJ04P/WhE8buLy5VwaEOFD8TtUXd+1pQ
0Ulh+o/U/sevVvhCREDvq9uwn10ZoEwjBL8zAmI1Z3aP2k2S3hXf83adJLD7lNPr
fa1ibvDRHZWKNyts4np3wXytwDfttQfwptbmkEOVHrY2aUnlqoQIEsInktI0xxxq
xrK284oUyAc6jKCk2TW+znYwVUJa2/m7Ur3+/7yfJyIN6TxlKytJqPRaDuiu2tiL
HKb8Ylo3Yj8Udj/aXvH2aRjzqx8xhdruzsNh5iuow9EnGqfLhTZ9qKv8HVyaaO2o
Mlsoc5KoGf8JVJQ1Zu4oMt7Tp3GMkW/6qe/GbAdk2R5dHZfIMb5JF6XnwF43zHEK
8bA7F1FGc6fbU9+wz/NPhDyjKvewcHABuy1R4a20npr7rWppafWTH9S1nbThLTj4
1USEH6gToK/wPNhBG/G+g0ISuV02SaIN/E5kek7mYQXQdaleY1cEQMxAkZ3ylR38
VQDbHh9H8MNGAe6b4YAMKLHZHKcAIezZ1ib9q9ViN86lXEJxEMd2tUY1qy1kvXVo
oTtf47Ja+rUuAR9ZaYN/DI5IOKa4UdZzrDWn0CIy1L9PI33ZmSXoQIIe2+50EPzo
SEkAZEW1zaz5u5s+DglZyaRrZHgoIUW79zhXfrzsru9kjXG7m+RCRTJsQEVE5q7n
hZp5Pfz7W2No6no55TJ/u1ishxFuHbEjxcHXoQ5YJRt94wxAoCSqbHvIVuegWDuy
OGh2imqsfIyqzv5IqYx2sY05dIw6F4S4snN+XyHtU5fAbntqvAOa9+IwZwlgV+Kg
VWmBI8a41OpKYV1K50Xtl88y0t7utzizdn6CVksM6Y4h2ViVlAHg50JN6YJAXDAO
fjsZCt/D072jkFhgLaWjJMCrRdHRQ9mv6uqxBoKIZqFOskgBoh7yfrrH97Gec667
qsqLu44xtWJodFn/JRhNmgF9Rb3+8aRPHhtevoaHUSGYbwubXpUFOoOAtpBVOzbE
VH16pGb4tgyQW6qI8W4oaAtymVnilfF5vvcyDsxIpyg4++ANc/DiQ7BwpFzTXtcj
X/Vav2kGCV9yNe4UKebw+D5Y4dJSs+ehUfFx6yvBEgFcf2yYM8E/3Us6AoWbly8k
LRNZnLtapNH7BU6FlX4w4CfU7b9NK8gj0BaHRr0c3xan8ZATzsil9f0JO1JboPUB
hJBX3/KwT7pFjhTuoEkXI1fgqYJvKPBaRxTcRKl4JYN+DMkMueY0s4m5odDkAYYI
ojLKA5jluYHw2yY0mFCCTfNNJno6qEqAUrO4Yh75gzCk6amZlLVxLj+JvY888E9b
/dDex8IKU1Z+1ECteowTglGnwnpRpZaxGyXzvn3l8YO+DYRhc4hwRaIeXfHZ1MF/
WcehFiyackZy4tBAXS+h6AdTgeyC8ROatZpGBuiY6OqVsUUY4fOR+lZ3Ekxe57jx
vasYKLzIm6Wj06/HV4YdmcZScN7W6AkR9jGe4330rDYvOlWxhzwU9JSrV/L4juBg
+hvB3WUdKNfw3NT5jf1t/dhzKmAsIhA7Cw2VyFFWKm/I5kz0CU6GRQm8fTrTcWKS
y1Dxq1p8D4u8ENma6QrbApMBFMV6WzNtXjyuHO/jTfVmCSJ5/eAqVdR8XZzsnNKx
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10368 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
lmOQgIOM5jiJrGbWpsW/8m6AI0QamD6tHhrixTgFXzdakMbLX+M7684Hzgt7Ms7N
xNR/q4QkFoLmNHs3AqXRbReBSxa9+eZpfUsFT2L21BOpzmE/a++xw/Cztd/YHoUH
JqzN5NKhdZj1NUQpLvY2/5VldPQ4SCNRseG60R+owrskMaDjWKf4s5GeBaqMY10f
Q5yMrRKORlqQNjDzNLieuA/6cCXL0gM9P4BW7TFst2SmseI1BGiNfcAbBTQu+WBG
8btgp/3drss/6rQjZ72NHhBpl9KsKV3MMzh6rhlz6fGguOA7MRZBnW1hDy03hlC+
x+j3UYaHo8fKINMMOaQ0AObRPjjef98LVpDL6q2kC2+Yyptw8U2AqLPW0AKqTRV7
pq+WWepjV3ZQ04pkruB8sICSnEWNziQbTqMFSIWsZ7SMb3m8hZlfa9SbkXRMo3xT
jcxSo1NYSKgw891Qi50kF8utwhkfWj+C2+3ztMv107G54tN4ObIXWokthzzTdl/i
mhLYF9PBkhxLVSxcH9QQsMLRjnSFdJkHM/YvRfWnwo8DItGwClzroXFRjZ5UWJJe
zIrXJHijyRfAEcQWsx6PyFZNEm6eM5VdahS9fGuU4e5VORmISKnE+75fT34svpYZ
NlUwVqvGkSXbmnPrvxDzvruF4J5fEH+srPoZs0tYgCIe1BcR71YB9PG8EDzhohNk
ahY8asLN8RAbGDJ6yIOAEijkSTj6p3lUMkCrAS9SLu3B6uxI0PrDUzv5Dh7izZUQ
WhpfzAoQk3U8WIIioupocFMMjo1a6pEUzQD+CbkltR0uub3/QOmdNNbDPrjt8wB5
uM2adMNDXeV3pk5SKE80E0nzGQzT+RaN6eaKG3tLwqsmTM9+JuqgKo4N7M8dggkM
rZ2tD8/5AFENANV6dbPJM7pP8tAean7WxBOL551oUGL1wJKOT066o8s+971SExMj
Q0JdbtL0LErN2TY2p6fTuspl9gS7NhTef6wlkTn2Ucgq8Xi4TwvQ4LbHm50fwPla
Jk9crju5iaR/COvOEXQFWOr2DSjXrWF1w473sYcij0d5w8Cd4hJjIyShDS9PHuqD
WJh17o0g8bKQaps0DUmyp2EHxaW1uLKKnhGt3OriVy8DwHZ7Q5w0vZlzzNtAsT2C
IU6aEG6RKUV4CiyegtjCzmlXmH98OI51ykfTkKaJWcFeCDCMozWF/pILSfWXbx/M
qN6uQwhJLrNV8y61tcq/iLDzwodUiM+Bch2kTbSfKz+ahmlox78dgaApgwS5rfgj
SJ3c5YXfropJtMQH11Vuep9g4NWY9EPf4Wqyvvpf3GfftWhc9BfpJSOcp3g1HcY9
br2L1LDqi+/b2+V0OPLtXh0btEGzEabTaeKwGK6rsF9tV3+UeWbH4hztY0XpghKd
2H7NODyvjJC5AhI5CDXoN1F7o2K/1jrC4hp13KYBGk2v1kA/nuVjMJkvcsO0iRpl
Ns8nJmPc9jwC9Nw9uhQslTEyjSTSisZJ9GaVCys25dVbv3uTdGSKY0xKXFu9cNCl
kDxacN2cPRJqiGoOXiNsnxG2QUKi6cnzolTLgjRx7fUx0mmP+bjEMm39rG8fBjDL
vn7fYq4T6aI4JqFkFGvHF4skey1a2xsE87LozvpZoQbqQbZF2Nstc5COCpW9fF34
msG45EIyoonvjWlP86UnM94yWsVz+0i8UfRLUmiDEJf/rNbpoiStQT5baebjxDs1
Wfn0C4Hos8xxKC7fctypiW1zaxRHHQhnqosgoxLmTuCT9VifhGyc1iAOinRpFh5G
wybakCWyyfWjffWg3ZS79BwLHSvhCAFAvBys/iQUmncXKS5h+5pDAm9nrmPRGbDR
TmBNeJTIc3o2mI+bhb8XMj0pFCxouRPvFmvY7jFK6xmFLUBKwAUJQLge3bcGT7JU
Jj5Cpd9wJhBLNY3v8NmR46e/IZ5Mf+RjqbHJ1TOmZRTKzBlMCRfbo7V8Si6NRQfq
1NwVCEMT6DQnSkMQsYFlCjNWpzdNXi7A35dlmVI6H9k00roorLc2HpFQDmwBGvsQ
2g5ffKuaHGmYWNtuNt1qTi5bNDMd7V9p8ty1s1CByxuOBGecpnr3kv4QJLooaI0b
NRy0WdLToNHJU1Q3omaRkmie2qfwEKBV+Kmqskh55v3Rm39F2zx815jX+gM5m1T7
ShrmM/wTWkZYAsnxvgLVrAOXr5zOp8RjY+jWz0D1ZcxhQfl1AX3aQwg/eXtnugPv
SdtbzaL7XsyabK01ddKOKbmOONHrSOonwm+3yqKRCqmmcYe1OMQTLWXDVGqWs4kI
5NbNmkFC9t/BaUXjD28inJxDNprFUrtVnYM5uApu7oEil2tWGOIsRGUV4ajuerN3
kQ2pMZe5NbeyHhXo1LDDfUTRuyBrn3+DWIvqCzkhgs/aju1/0U+qZB8Zpj9F2rbT
SAkf06cR0224Nr81M10DxZ09PruDxO/xJ9Fr8xS0QNgitUX0Wlo6m5ZxN977i3hO
sZID1hWctMtReVSjN6j5r/NTDoyOPTABpVmrcQ71brhYO6IhPy2yL2pxNb41odKL
Xq1eJMC+o0Zno5gDhuWTYENoAbygzrt510QhFDy60GY6oOfrp8y9Z2t4jNEd4pjH
qPosXfKm1jze8hAOYcYtlLVKPaJezPKzy1//JtocSLpwn4Nj7ABmL6Pp/7hJXM8G
pnAb6GO1o0CHdBkmNylx8W2KfbDu0aGMk2NKBbsKwmTpvenPQpXTGfFH+MSMlEag
WTHDafXT2AQPF3uSg9ttpS/sfWnSQrqGkwmINbpuID7Ffc+k5D2jipG6Z6r4kHsz
Vei3eMtd/3vxlxGBQ11Z7XiiE7K1eJ/tcRMaRWaby6Vs3J9Nvq78g7iRpmsGROEU
eoaflEyNeepyNJC35ThWei1SFPG0ky8ISB2UlwQQA+hDRaiFXbCCufR8mkSQW/3R
f6ARTN5JjrRGSQLJelDCxuYkPQaJvtdtug5UytKQd2UwzouzT7FoMF0mNhgXX4O0
Vi4F/SEoGwDDONlPqXcoaaIoVfvmwxQrzk40pn5m4oOV6Cs5TnfwdZUXAW40lNxT
HRAXrJAbUMX9bd05G+pQaeYUTxCn7vzHQ2JQ2bOeyjxE0Roehc+iNMV7KXn604y7
BdEJS+kv47YsoH+Z1UvDPg6kPXY5lyEsknz2ghHfMIsbBYkLco2XI+MNq4DxELm/
ogaDe8lwsoB2orcQeJZY1HCpWbZL2Jt0mE36V3y/t5g5mT4HFwbXImivI1fuGByR
+c2kN8qNi52UtiUgCZ/LGKYH5+5VuLFdr3sOrTmSulvHwGMbI7CAC3FxizFE4TAr
3hWaT+aqglxtgsLX5t6MQzRPtCMOnYTfQyjYpjkuut8pHhlmiWz28jfQ0yo4kZeH
Qwz1oONAGobn4NyRTt8l9oOHm6wbAp0OmMsnzfOO1G1KKf5ydegklLodQ1vsVlfx
oDivq1W3nMImK1GwuyajwFEaJXwrmIfIp58iGgr4R5p+6Pu/1GMU3XfnuNHJbKE3
Ge6g/rSiuvgo06WJpwkNT6+auXxSDDM9mwi/snNMMLOMBG2DAg64rIjkpdBjhdjY
faaRg8m53ZFu4mOuk6uzkmEzeaBa/6hQMjXNrJACjF08v/65yIZwD9tmlGhRfDIl
gQTPZXoesWdXD0y9Z8+3JDL2graQUDpBDD6BXIMIzWNxyGUK6JUHuRsLWOZvopBF
GSNI9AV36fb9a1yR+nRHHoFjtD31KdDVVkI7jtlDPfacP/M/otilujntOrXBpqO6
Xwq6zrpnjM6D4TQMF+FgstoBPRDhHpT5FqTlAqc3vRlAjZuODOuQMlVDJCkQXEEd
E8whd1HkL+sAG1L+XJq/f/vZkKwl3IKTQYhKcgiqCsgFAG6cw+VeOBPf/txZeovT
Yge7LbcTc+fbhVe4+chbSvoDgFRl91iW4x7M2TTUj5bkSxtv3XQWZxnhr176vtwo
BCgwQWBpe92wddiEggdCVhQpaWJbhebptcXsRBsa/h/12PMf6QwayNCbHF/jGFA/
qzJrV3sbb/cGzZ84Og9kbu0sdpO1tp3J47wn4L9pF4lemh91x6WIEHJpT8qGHcFn
iAHONwkAMd7VDXIufdT0NCec+LvTIdpBQSlMSypJNAkxDwL71+mCdTyKp6CNXPon
dc5TDoexGEB47oYxtuoSxkGnWS03d884uqm2mjCQ6t7pns+QYKR8L8zo5PyK9wNc
g0eoXik3/63+RSBQuHAVqwYjYVheNvS4VkstjE2Hd1idz0HuZGS3/xcJ80VEWC/p
JXJMwDckowKsaoA+uhSoqRXq+OPa8AyMfVz6kFApg2Q7uBo/NOi1lJJbNIIiTCcU
y9oxg6P52ulH6nqhr2XFqeAr6yAIkSxuRR2hjYZJ44iZ9H8eV/6SdcdVe4Dz70oS
pX0cmHn6jWGua+bbVoKNyYUqP0IWwPkfmgYiRaeEqQAoBNX00/n3xlvRXLYa3XBy
m5j+duTbiMg9wtri9NFa3umvWSvKBIK0uCfcDVKUY0UklUtSU6FLqy6ZcZMixN51
3I3Wj31i1/LlebvCFte3cNLIjjAMCKCfpeDLB8886RdWmsErDHHnIO+RPMPPClRT
2RQCIYwBX/CZyZGkwyE3bxq88TTMvZAvK9npusXetuMr5TCkyK8T/aNvyHz450pD
3mA76cPnCPP3m6xXg1+qFLhwyTzEVdXOiaPOi6khlWqUfbt/BecvasMHQ8pYDyxv
r2LyYT+Ufmg/a9MbN3qNVcsTEuu68ek6wEYCBi9msyKFcGCs6Zt/dUZJZOhvhknH
f3nIht9UTmU4NpLvSM4h/uoN89qidlj1G9PrvQKwVu3ODgB3XySqzxoZn3BdbDc1
RzYu/be5Kp+nMLFI4VeV6YCAlF8DlQAzn4RC0XtEj4ahnVVv15AmvUi6rgZjBZxZ
2VvwMMpIvf8KIOI8p4vBMgBgdoMjHyAxpm55RVnVjJC6TkSIxpmLQudrf+Q/hVJx
CfyJRykdMQh4VbeCkqeLjzy1oVYYkCk4IjYoUp7DSfo06fsxgNNVy4oUryGGRbyh
2BKbb2BZWtChVdRlgQFrmLhUFIRRlepKoWjjkKBlfWt6jUFBdEF64jsLxiz7U5/6
GlJvpOW5R82l0fv+AMDmztGgYgeSEFXib0FtERe5nZfKxNE+E3cd/+oqbu2OW8rk
ocp1LxVvmXWc4AqNzeYIX7prml1zI3+SH4eMt8kXvBAhyRPmLkyqhPmnBx4iUBSm
47+ITYtsy5REgDEjX3cXPjtfhw9s1j3C+iOd3ikA+ANXpwtkGfVqMl0sPyAZDDJq
nIkrUt802WIi8jYnDrlwvnezreXYKXHbMknqdvcstB5PV6zGkbNPyZBv3PPnfKL1
OMfnreYePOqODBGJCKfd98HimDnCqnKNOcDi5ziXiuzSsl3v2YKqqi+6/uO1K2V4
ZZbQe7axIOCCMY74ZanQbz+ueIs6lx0RBrZSYhVxgSis5fW4EK9nlN61UOAfK/gH
Dx4MBvKb3dfyWB4g56KTMMSSZrFQWe7ElaGZ5KDc45A908UKA7f0wOIn6SvTB4iC
3mKNM80wvUnWYt4MpJDzPjzkJ78EwTiXfJrfxE7tgqDabpDxVX/UnuNNSy1uN9Qx
E/NMO53QCVMIzqLN9G1curO+9QTzM4Cua6eEUWiLyq9rR/vM6ufoXvtmqEFaLbz4
s4xLjES7irqoepn+vOhU8svbyDmPodPTfJbmVaYgi+vQGXdAnSep9iOSpqZww6sM
30M9GVayHWz109+bLxgB/zN1RpSEnXKk5dPY6Y84Vxzj6ZP2Qkp7UpgbuQpKA+Aq
luQW0im8HNlfVJJi+iRBt0h6Lc7j6EQcCWEED5nwbpkADauZZvW9pjFDexD5CRBo
su5/SjQE2bFhesdqBhQ3uFC+fmalgdlO5EmbbzAPi/2sMmjGJ4Wfap9Ttl9J4Kpr
eJL9xmR5qYwfg8Bo8806lXBR1oBhubIB1ERaQbHKVSzBQp/QxvDrp2pmqvlW96xF
eQ3S2GYMOoUYW77bim3hEYzM+wQY+8vukfRH3ZMZ7K+apIB9h7FnTYvSVZr9dVPM
ETiq+NR9dhCZrojaTcS/1GbKlySary67EkZmMy3OfJW4V3l2s1/MKBx0m8cvjxZ6
POmnH9hToLvFZlx8FCFKOm0sj81+dNMj7WdGvHD8DznrsaIk8NbEzGJkOd7ret1T
H5tTX7zR33tzYht93ua+fzGy6QSaxiPoJrnqRmQdJHz2J+d1L8vVWxM0rwVkIG2z
phHAKEyi9zInqbpyZfPBWz4U4XYJuLUva0CXOGCvFHJEo7nPhFMxf/qyNaNuse7N
nT/5w+4/bJrjUYYq1rpcvsRGJvSMAsm8WxcvTUQObYOoGwjd1ypx5DuX+/cj04X8
F7Wy8+EGfeX7zqD8S20lRoyeL1v+Vv4DOlEluR/xH/3pn9ubPoxy/UL/EyY6DmNL
47HqBA39O0kG6k+FBY9w0VPn+E166CBVOU3hOpMu5QsH/yaYi747/KIEEVYwJ2wb
J9TbM0rxUpgfw7Iz7spMf+x+8WUlyH1ogwvaVxHtY/fXMRUZmTpMK0tN169kjA/E
vSb62FsRgcX2beJUTEyp1Yoy9mC7hYdMujezLP1dnzCOlpD1ZGLT+0C1Hgdcm+O7
ETO0VPZ70OeAUDjc+cK6pJi1tkOqf1spzP+1IpnEIB8uAz4LoaUoAkrZ56rm/K0D
CPvDO7Lg/0NgyQzryA6avamdWINo6seOLUNsZ4cXcjYcP+6A68fbnQWtYzk5HFF5
BUx9eRd3zvjDisb3Mx2fysfj2vVGQLiVrCYUof4M1GFiS0x5kURf/A/RX2SGjlaw
fPDC5JyGtxMfQU4oj+7PvcvxPmgH6xjKbH15OTyJigVei/gQHOz/JVZJYPVC8Cbp
IB3VhV1KWMaJu1drebnBstFvxH4fAnzgLRMoU45BCpKf7ZPVKlSk1YrJThyMZRaN
Fc11saLLLKGoh9aniZ9xvit6TE7RhoTH+bK7t3uG4l0AKaoEazBNoowZG4kCpPhu
GKr5GQok1h9o6DUPBBpxswG/Tdvh+0DTv2Ic+OM3cL0Aeg1cVSK86wIzmLDAbxVo
TV6onsCZ1qoq1uHUvI8WeDe7/6cIEuaJML76iPXNplNWZ0bIJwDPvsn5GVVRvhMs
SjTi2gKt3NWp9DaqIUsUwRFpuMmlx90eZo8939TY7TVFFoFJXX+TYtGGbZXFZneT
GVeGEveNSpsQ0KzXce7/yiEK8p4jYvUhIEI7eC+MsOdwiUYiGR5x8xKG2s/pK0VQ
Bju9i21FJJY21vR4O/OY15X8g2PY++8QircOtMUhkBGqlA6Ef9Fy+uvyWDErLxzv
Wf6wFsHTTkE8OTsfhuFTgFaW2dBikKQUbEJ/5wTT65JzUwVi0ojYmDWA1B595Hsa
wOCgYKf+0yV62MOmy0W8ywOjtBznUJiNCQiVLCGMmwjtn6muNo7Zmos5aCHxhejE
ESvrSI93fDfSqsclBa6I97blo6bb1F8JcW7IraWZOybdl6/isSh/jpzADdb4W6zw
K1+L2lOh5K9Fl1h4fAGbvtsNSC9EzB7eTUwgOQkharn24+dTme1/7Ye3eqdxWj/x
rb7tc8Yd0GAuyqMa3y9R2PSv2X4mL3SKV8rBKhuXdwOYRjGTevIrQaV0/ha8Efme
8uIaR5RnEWU/3wsslBmZAfTVGXIHDOfZOACfe0cWlxJ5oIFQRiiD8gSNFjaly6YA
TkBHOuTKgiHvaWfhCG93HgumUbpy7NFjJhQo4altAoQcehyScRYyyv3OThu3U4cv
kWjnLV5DsRF03orWMt/BVMPT9OhX+Odh0WCqyRHoQXFbeISwmxc+kPyURGsnO0Na
g41UHeu2cDUdG87nu2yk1WAFNfwPPax2ICpbv9ZeoeNLC8tWbdYuTbY/Ej5l6hD7
zuu1nz+1FQ8IHZi9MUubvy1HhO1iSocDMs+UXq8zTr3ntTMaciedZ9S+IGiCB3k+
W1CAKZk5YZjmyeBNpUylWprz0MdSW+/ksNskTBxZUcbVyJy/jM1JAba/QgeHtI2y
1Nbea55jdohEx1lPiOmniuRcE23IeY39AO9Y1qmP/CbjjxrjWhmDWOZJ9dLT0Cjq
pFKulst7hD8wMPJt/uYaoOVTRHg7+B//q5566SqI153ScWccsBNV0dGKC2I8IpSv
vboxu9QfPyJvdCdHzAf5hCxHMEJGTQea2GlS/D0MAN9McPuc7hIItpBR8qykeOUd
xQ0NYN3+jcUZUB1ZyK/6B0jne17veQmKm4HEGS/0zdpnm99R/ngqThjOlEwxcYiT
iea3mW0C+9P35VCVUwZ3Bovu1H27Ji0noHU/pNuW0q7gQjy8K1YNsWYYcxRAOciv
4598Sh6Sp1+QLzhwTDz8ARTjG3Nh0SSqkgxDg9BHEkHhclj041cUHAVNwb7ShoX1
zW6+oxyLP2SXvcXreheCneNaK6goLVpcUK1fMgebmF7uaDogBkvlSahrXiEpjthi
AmEl6slEW+fX8uYopf7NTS5+/pxE7LUnv/fexPwwXQw+dS57NxRRO8pVUAiiALXd
3/C04tk1y1yTq+xOFUSJd+P/Bvca3tzyp0MAwQaGhiBui3BXfTaR3eGEgu20Pkaf
xseeJXKypwswIbgJWWgXErs6BvivI48RgKVSbiDs+AnF37LZlSCG9DIMaojth9Kp
lVbq8zAh5lp2bGkE7M7l5d1W1pWVy3A2Yld0YL0D3HTsAwwL1qVgDBVRjftBvqD/
tLCrEv/8Op5vXge39oMLUMv48x55GY/37PvmabQZbUY69TJh5aWeSgW/2U0NrdNv
W4PPobJLzBAmL0gNGua/gOj8MaYV/E//MXQD3tvxKEWF5HbnlqbbW0+U056JEj9K
iOL1f6nXJG0eKJZ6iaVC1poBYa/PrwcPSa95WSnOv5ZIvFOuYnJsQ/N65/5mN4jk
YJgYv6dDlTZgE92IBhBkYAgNAjchN4ETE8Yo0xtJrIne3cPeiOtjQTEbGDsBPPnN
Nf715qom8YLgZzK1UcNRv36Y8gsqyGQv3p0GD5USrHKVEZRkvjnnKRmUJrw90wnz
GxTl31WqqtPtY/gjwwS79UxeINyejRzY0c3eNGA70wcQwc+ouB2k4tNgFgf5oP8i
2s0dVe4dLCXnfaKL3AgLIL9+FYcZyywhv4wWPWbBeWD5H1u+x3sK3WoGGSOZaZAN
6vL1+RaJ9stRn+fZj3QkWjEv0ANSi8qn7ItuhgLWGbpNlPUlh8+n6gBYNB9GDfWV
fbfljzDkkqkq35qCiH5nkpYwl15m4ltwVROlMtsmG7GN8OVT635xoN0cB/LiOW/6
9FG5pauHcxIKZZoLWn15emY2nFK6+dlQS+gMhmBEhitKyiznk6JrawnrC2BUjuvV
1aYDo5kxFtmtWqdwIdbFnitxuYtadDydmyjDRR5mrY+YVusABpNnIMn5QAKTbaEM
WhWmBCLtwk5U+/GqV9BMEUZrEPmxOVwfitL7O0quhF6tSoe+h5V6VBLU6/z0J/ay
bsmDxNO9cD3/xOxTse+JQCcU2sX5dl80RuSpWdGyvbbeRbm2vu3c2BcecAhz0QQD
QDoIkteU0us7Edug+6/65+Cppm019x8pJmvuOA4wtb8149MZUCeRByviU57DwKV5
uXWhSqj93SIOb17rn6r/RDDS+guFhylo0bFmNKn2nSo1tyE1UUtmkEfI3p0HMMU/
v6ubdqpuGjA/2SX02GQ0bHedin/Izx6KdggdNENwQdfWI8NCTQ94xlM8/3CID1x+
XHyvAMV8qUl1DOqCQQcWYqz5s/1sI4LbyGESGr3Rn5o9k+LQa35RajXJHbYazcgw
263wG+tclnABpr3yMXok4lHQmB3l7ZTsxbBAfFzt6XX924KMEWkS0TcoTkmNj0gw
m5KKbNAkxtCJRtP89yZWnRiSO94Nfg7Pt3H7uHRpa36XtCFsAL7x6xJ5ex/DwdsW
5EVxdmBjr12XhRbx3RKa8PEX3ab77AXfsNwDp9bCuTHxiyTz752/48GQBo2MZEBT
R66HSCEvk24lME65wHO6fPO8g/vLs1w8yNDv1/mvjsJTJGPCPYkuNRUdyYTuRCtc
n8m0N/9KY/sNLSiTkuTqOGsohJ2a+6vTYTOaxhuZfsjxje0wdza8dj2yNVJ9ntym
0KAMc8WTGv9OwmueR5Dd/fgYqQ+K31Rt10GAYdU8ZMvlZ5bShKyGJveSvG4gW6B2
UdN8fIuuDgEVPIK54dM4IZv3xRbfGhkdgs2vRFNYWULjRMFVgoCrxw/5SHta93eX
kcjdDp2q5nZ+1w6YmPyIWqvnawhpUULHeRP8He8aDnQUMbWlnFonc8YocVLSKZxP
WiuafI8nFV6FiDJF5NAtWsbOU8QrBqBlDOqb/J1K7uJ7/j2Rtk34+DVeQyzoJGu1
zLMUUON8mo580nIGqLD9edbJF87oiGD5YftyLzKQBaPHY5cZb3BHYbl/7Fxgtcxo
kyoPP93vOG0l+lorifgW19F5FcslPeXdPBAOfr6q1octX/qKXQiYuA4bXXjERyk7
QMkGhUyugcCw13dpBsqK5sDlQoOi4hKqP7c45CD7vffrPId+3QeZk7jdNmDDZSrq
RVQe96ZawPezeBqmZImNneDsBLAd+wcNwaK/RwM7eeOz7StskuVw3FfIsbfsgAFI
dIgV7/y0kRfHmYAnc/xINTuKPhOS/gvISAVjW5PvTpqutotAT9/GSKsuw6NyYKVq
JGW0j9i1JrqsvmmDfdSDKmUu6jpwtfZ3E+gXl+De4LaAHLnz2d5C9qdEmCAERBOc
EXdR4mqA5N6sz5BoGWJX2qFzEQN/L0qDwZn5o124hMwpDjjz7z1oddhzAcf6oaSQ
D9HdU3pNtTwY4DqgihTow8CSx4d6c78YuouUi1QJHvrvmyBNvI37dxAKq03PuXA4
Ezne7aRwLDfpCJKlWaAh1OBJxWJQhZwwGUrA//3QXtonuRHqpcUky9omP6RL8oVS
yn/uha0lCuSjl37Yaui5aQNNFkwvjHryBgEZHb52Hs6jUktMa4pmydgOId+5y9n4
CE5jB3oq5l5y0i94bansisJH3DcjkiucLvP1zaCV95KIDhjG4xJb7py19papbNMf
fptNu9nCKD9nhVr/fwvh5ItPDeckxAo0ZllA+yTeL6WupbbSdCaQhhG+LTAtDvT1
nurM0rzm8Bmv1CFoExQhf8i+U/UWsZEEkzZR4YXoIPjIroF2KM/B3nDfJKIDevtv
ALK5GWgAIpr0pWXFajyv5pH1g2vVPypv6nt3z5UCngr/7k2FkAlLGxx3IKnmiv6j
ZnC5IDOLRl+kn2WD3XuQ/MDZBy0aOmqbZwoFZokQH7TWKPFipEaBy3tg1kawuhzh
w3xZ5raySyY0QwSJxJkdQec3mKx+1xsruYWjQShKWIvEoTDH+QYoJjW8VjUq6Tjm
ropaZQvXdBXzfhPCAxHiika2zqKVHhD9OZPHKANkkLyfKVOSh4nfPE4fZQxcziYW
X1I0gAOivMs0AxmMum+LD6B1sDmCHirjQXcsRIQM9szkhbTdxLLClrmhUPXQpl/8
FUJpVGJvo9vpqvWt0OLk2t1XDbKfW19h8eO77pn9lTsuMXoS+Yo6xx5KUbnoi9mz
n5JT+yRXFp1DshPewMquetkN6hUkfkTFmQZq4C/qQxCXq3/jGo1hWS+S+W/SrNkW
wHyysVurpMXC9fMlXYXRwmHYWFAWijdJWlL4z8xl0XUUxOgT7ug1X7knLFre5OeX
QFhG6hNnoOuzf4OrBBNJSbmzB7Yx0VY777X68mI91TotLh5j8syHlGzjBRBrnqxN
+4S4usiDbUEaqGAkskGOz8Q6yJ5Qkp2adNq0G713jU6BQP/FW3bpsk3jqu6x83GN
hvCv5F1jVekOgFihmpjDh1nZpHUqp0DrLEVhwaAL3chAm4+5mlNImaGQH5zTUH0c
KGZKOBlZ1vJZfIBST4qLoVc6WMNSgNan8rog2/Y2B7p+ER21ekN6YAoAXDWpUcVZ
Y5RGNFO2buwn9+E4W5Xx/Jjj3aj6lITW/d+PPtjlT2sQSZCAw+zl+hRs3xHcXNnM
/Rdk4TVE2PVnC36j6Xnw8S7zu/P/4FQJyAQx5XSxw1DR8KoOdkLzdI5A0kg044I9
ntH154TIWV+BBsBP7tP34NyQO4ovTWnLUd2tHRubRKkFXGIi5aJzKEXqJ/NkvDAI
hUGvV7hXS45ZtUpyShUy9IXpaZCAKkBYw/gZ+I8uYucE6Z7C70yI7tnHWppFzVwU
dX5BIDypRnK1ueN8CkBaejo2vnk0J3RjL69vR16E7MV2O1VJ7KTkZo9VDaBlnwX1
njKwQqT8dv71DgC1MPVZSOgDSJg/iy/+Wcn32l+3CNRA9S3TYEout0LaAY07RVcw
1jrLoRh6eZOjkjFR5XoSZn7/qdgcgP9IXABwu6rmjEZqBLOJDYC7+9Z4RNk5OFw8
NHHvrmodpN3f+NPuVgNQwzvLHty8e8sXXBn9rw3P2RSBMchxeMeMr3tyMf3GLvGY
UbcuAIyNslOj4BopEFogHoJ6086vBjpubuO5KuOfC3J2Ydpk9I7qooEwLgrCPsSW
JOcn35eVngDOVqg8meqT3ifLbAS+poB0uFlLnEjP5s8mgkNMMlXnFJu+/DnkDqVC
/ZHRZd6sWo55urDt7/7aehCQdnAhPfXO1RiYR+0SqHAq0Nv8ooFMRjzO25Xwm32g
HL+1HodFoOQC6CVNmgKFaGntHtI7sY4YLeTmI8crk8IDIynfbQkYi9f5BPULW0TB
wsWIBIgiydqjnIB8DsaV+eTZSwjl/7sECLk+dq1qBSSQhhKtwJKAHIca8J5m/Jx9
zLZTxZNKFBm/sSByLjI4/VLaoAsbu+7Yz5ZWqFareUwcaufYGiPq9Oo2+GL7Vknw
PFK8zYmrbNxLApCfb1JmXFdEpyQrDA/zyVvPV+0UiU+qlCt1qXBB314cdw9C7SNq
y7t5+eBFz021YFpIhrdxe+tqj7dkzUmzd4X453EaZhIXlf4RzxygYs5p8HHK+ILs
WsatqEHbaNHHOna9h044BvRsUn8xBgJgCSaIxDFPJQQaqQZplmAbQr865MRhNLmJ
Y++FwTzYWIa0KWsR0xSKcQla8t6d9E/4HEabYDSEBvtHmMIKUW8GOmaD39vTw3c6
l1Ry6RcJPwLpKbl2dCMBzu10JSZRo+2srwuR+WeWF69U0Uw5is3zaXdpCYCfVXAy
z1hTGG2SSjpwERVcN/fKlumaAKwHTc8ZFZ62b8/pj1HbOCuJNgNaG4IHe7ntCnvz
kCqXEs64vdyZ8vVgs2lIHoKxjYVms8uXkwiXCDFCcdKyo53QGoURr7skMQ57T4ro
BMVDM7MkTj62hQeRvYT8JM2BPh/YYRfae2rfCbH2pROvjEG6UK1Cbk5ieyro+cSJ
yKHU4boiviQFyIfNyoemyejUPZd1RrmOuOhdTmYVjOHVKE4LpBlbgU1wb6pB/yoI
josh+i3FyNwd67qw5cfM0vmMNFu9ciJbCDcpqCERqrpENrC7wGeggpLVXyx+ix2T
6SwIgaU9w4VkZrSJ/t87suvz8+vQpzAM4B4PspJDjJG6ZabmmBrEGrI4WitYsClq
NalIClkXu7h8YSkmRmHFTx08V4gb8BnQbAmUFvxRbRNfCpn0f6y5LJS1LCt6FZ8Q
>>>>>>> main
`protect end_protected