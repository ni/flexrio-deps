`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8432 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMWORzZC7bo0toZS2Zods6Xs
yljw+BvqICQb54hGe2JGpCy7VfzPucQWBxxbAs+GRajeTM18BBDxG46Xr8Nx1Wvo
cRQgBp+22l9cAGE/vFqx/vQSAPQlMqK4YDPG74y6guGSY+a46gv2FMcJY/NZhtGb
4bk8j6mYnp9HQYcASLmXpINFo87zHzJCyYapXzcdM6yVd/L7VZO7FfwCur/4IFb8
us8l1ssSPkcPjEh9SXPO/dWQ/hZEyTMO3r4jm5U8wRLGV0aD0hNdnNA57RoKok//
MhrW7fVMm5C6uDeFl34HCASn358g8b2dpqHeietpkxkh2HGjCGoDJWysYYNbCR6O
7n0E9lJ6BbBx7Xob9cWUvG0tQDXE4QI+uMiGpC/IqO/IGVt8SML6ZXocWvqTrZyp
LmJTKN9JQQWRuemRqWaAK3i62H8pessH2gWTcU0RaJpvGM2Zncb+dynl+BrZBO8i
wEcw0TxXxdlt/sGrlKUcu3ePAXjR5ldUj3noD5e4JODPQBeyC6rHfpD3gVJEuyem
v5+Z8b2Ev7Sc4hxygm+GMy0UBhD31C4xprUQUtFbU4pPpjoK6PmL4HYN2IgNTX4k
gbtmHtPQT5QPaPFz1FVgcHm8dtGV2NGpqZpxkIBfiW8I517biEtkS02/qdP/jNiD
e7XRsId7/YJSty2QXJwq8ndGEVQyvXEbw5g/YDairUkqzgCngtsDFTJgkZ5Fooka
ZXGvddHzv1R5SOiAGxWxIwIG1C73hdu+bq+RSqAtj1OlaEalHQZGhnqZKA38wKtD
PGYTXOobJYcTzkyBj76aWc4IfH7ah7WKC2CIhHijon3/l9kYQ0ZZQnzM0crOcOEV
F6aBezfRiBuA9bdIukA50lagy2+IvbIrzn/aQa9VaAG95UYfW9xFZdz7qaavGhan
Cw10BYfRUli9AhWQ0xak2JV0sZyI/76w2B59XqfaYLlfRfwtB+vRbrZ3i/+R9kDZ
UAcLC4AuGG5rZQOfaQPI3TN+KMZ/zntz2ArNHdHrKgpd6l5m4iJV3nfjQiAFNkwX
4OXKC/4efAC62gczIv2q48WwpkpH00uVwLt64bm8d8ZcOKNKxJei7gfONdUVPBig
15MOLL6P2xe/n8z/3dkKkRaROsL43NTW1xM//4ahNQ5EG/uhkUxexqgKNRrY5iU2
jdEI7qxlj29GclfGa/jJLgsUroSVhXRFWEdvRxiBcWsYcohLkehF1eUVwvZNg4GB
g2p7oljCYsiOUae+RkgBJDnC6++ZW2dUbAFscKX0PFBEzziUJ3vvmnBVITJcFIRZ
CzwkKr2WZlvbNQQJ1kuYSn7mRyIYzLI7swdLo8fsysaE41tuRuHZ+/V1mrGsKYNp
X8ri/+uc5Dn2Z3Ftr4pKYpDHakOo0QZgFR3rFPsUo4iDjgav6c/bZOWPb/HL5JnO
rAid8mN4DUg7z/neyb+X0Ct+T/zkOQUc6fh3MQZaW3WqRwa1PUwa36uQRU/EnEN0
KT9ht1GpJfYMVM/tf5NoBHU/X4oIzvwK3BKz4wzjW2TugPjn0ZgVoy6or3FkVaN0
vr20dbjQByvVt71TDX6AOwxI53P6u9iMnWF4Yb3E+eazX9CW8wxoRy+QA/om5aqw
18ILbd3G7wocMWmOL8ADp1qc6SYni8N1EiX1qv6tXqbMrgLfHzizYaXBCuxm7jXO
pOQkKe3xcUjwWmsygn2e4onjcAYzPPO/kGcFVkpLH6Vx3MTVBr9FU2gAC/+OdMvs
y6N6bmiDYbfaviOkP4uf0W1HWN9RiFm0rjqq20HGyhTdEZUciUBtBu8rQJIF/fac
yEerkDbG368udKX0Z10LmhYdTSF7/6Xdt+FwBRMb1XlaH4ATLVbdKiVgnC0MQ3+L
qEBmb55q+dRNKlttQcRjPZ3tfNijW3tAi+a0vM/ym5PVtUfcgrEq0Z9OE307rnoU
71C45MFyywQOlc26ZhLiMuuCCGbo8tNq0B2wElw/O/vO3Hem7cf2yIeK1W9WyEne
gVupuRLzXT/QJDxcfy+kx+7os+llIFqvufhnuYqDjLGjbY4D5t3ej5qNAZLYFGTM
jxXn06BCHPiT8pHJE8I1Tyo4bDEUkwiB3IcGc7UBxs35LeRLGoyc03+W1moT60FH
ZjeKGa6LpjVPOoSf1ieOnrXisNiKZqFeCvTnPfFw9OumHCIESlsFOYoCx40e4wOd
N0KlHbh7vlbqEJEMsnP2ndClprqOZfN+pK9cTKsNcyqKdkENo7r2KI3B2APIpiL2
xl0ia5H9g8O5pOjvB912I8/y5VJTepx4DclHZbkY7j1+8HdOJPNNZz1WOJSGTShk
nkGmE8axnRuu69NiZUxqPfNVEqrMQwp7PSyOSHE18r/uKvBElcJmdX0KjGdMl0Z/
eOApjfP/4bkfLDVuibIkaP1GeM2e+lvt1OFJO6AqdGjK2KtydOw3oX3enUpoPuBp
KEHBBb2Vf1O7QwpwPZFFEfztR++6hp51ee8I4zP8vNr4XKjmQC1gZBYRSSMUhr+0
R1Iab1cyVNUdabQO48NccGMVDNFCtRNVBlrSH5+3eIaH06FAwcUubsqhYvFx1fDW
pQV11snHCDeFoO+FHChMbgD7zyYXnSl5ILti0G/T5gzRQV6mF0asBpZpjUTibVoh
q3fOuBaoG8MGurMcozGl/y0lzGm73gRT26vHqqFzuGBpjizvqPWQSqP92esp437U
Vj0iDnLrm2Okb0wcL/1bzsXu5//aWCsAAzFOpA3PAiyAIUIEOl7PEwhKz9GNcb/g
vyoqPBnJ4ZsgO0CywaUyCtYNaNYoInDF55G1sa3KwGmra6U3RHsuW54b4f1S+2Cw
5fKhz1VyqcoYlXyYoeZtvJ6xxbOYaTGjEZ/1k7xk6FQPUNYhJpAvlqepA3U5lZQb
Bs/stgdmWvG+uvWCrZN4QjhxRGSDvgvvkQLwLNYQmOaw97OLdZjPhnuHgzscWE38
T4J9qdXzvSZfG+Nv5L93q51awY4Cm65I3n089yHy5LdHqJvAjJ2DZLX4hLouHiqq
zeY34+D5y9HMuOykHSlkARkgRw76gCjnKn7c0OYjfNLTl5UsuuNuuSyXx6/WBzr+
rEtvszGewohbnR7GHIlLZ67AKrLXx5qqiRL53BXeBKNQrf0p24wTxNVkyozBDC57
I6hno+6EXQaqDBI6MTu7n4xicaC640qdln+KjryxFAGf5bP3zThh1OzAOJjF90ow
QUm5vUYIf5/FpaEWY4tg84j2pOCJON5bVrM+NdL7RoHAxrZuxb99SqibJXet7alV
LOlFwLEKdd8KABX2SvCwvzgP2Or9hN28c/MZ19N8fzQcbGFe0DTvAaKOjbJ+nniL
TdM9pdn+TGlEk7p56EaKtg2PbvLrrMXxsTy2k2pMtb30L84cPCdYSXrZ839is4OO
GE0N8ynjp+zU0F80yiSqkwU4EKWrbOKOo090PiP5zMO3thzQjlx8Job+JAH8xySi
YyoMDONQ2tNW45mtIB6QCcyYoSRCvvweQZRUYRnR3e6f86vUknYi53Xvz0STjKtE
5HDnc+z8R9eeOwARoBrkrLTvcCkO7wYF83LFJ7Pv0yiAX5irionF0qfifdC3B/GU
/tdQiRjM86jcUmLC7nmD4tvr4GplEYX4yALNPwIrjwuRhLmTHUwfzJLVf4CAKl/z
6XrBsqt/mbN2Wqy0vWeqp9bf/cqyxIcI9NgdyTvwgtzk/owricHejDsAWOQmbViS
jmFoWNoLWJqeG+RbSqzdHZNA24/o+fSnQaGldT7cny4lib038UxTvoTVLP3Hq2Tt
lU8NIWCTUJg4DHLVKbm9aiSPqDwW2R+Dq0qgLFdZjZ5r1Tt10AdKNOqgzIN7T7KN
WhQEYosgbJCzRekqH+W/4XPP0A9MKbEK4ohv3YWDH/H/QUtWmqpatD1aFEbUAc/l
GVw6acyMiiDok/AIJZWjR05s6zKZ5AkrlR7rQXQo5ic/ZYhqWWQCdv70r8eIfzzw
zlPY8e7AYBciiAODGTg18rA/pL3wAkspVSUV1IzU+cQGw00xJiHVJWRCcdBGO1UF
WxwTyoKHGAKDfjr1+hqLcpZgW+nvprsdXHm/PFmWmi6rAJlil16Axr563P8xNpwl
3IqkogKrdmeLKoAz5S/9o78S7aVAUp2JAwoYPrj+jkH7IypD/JUFcgz/No7DAFph
2GIOvdG0hrjgEptK4KF9RQ+GyTSemjMzcAJZB0lkCzoOrAkhJxkzxl4QBdfq4BMr
eNb4AJqMwdR9gl6clesb1Lf/UEztzKqNDOCG+/vzBSUrujh5JIYuX/Fw35bkk+gg
wgL8FHCUAibZaBrenF2X6hHSYILp6IsOkwM8rvichQ0SB6qLqipZ4kUpm1I0tGP+
R9a9lqyFBL86VALTE7uhA+uDx08/bMBzbpoU/zoJoM2QBGTR2Eng6lKI1eNoE+Du
Y+pG1Yt/ARtWesomGZ4GN7PwlzqLDuGMXsUhChWwhxvj3szWajKRAv7nbBMszoZ0
qrLTjUAXC4b8TQjB6J4IpxR4Y3yETaaD+LKyj7qBayuYYUhBVRJAI70JiCUkUjfX
JJ3RoaP9lGJ2E6QN/zUgutJZhhbWDmR/COVMFA89e3u4jGjT21kuoXvpcxZggJil
clmHrPSKLBWIadHU3V8D8QtYUxBwUoHUDCdSp29uwajimaOLSa00amNxirW0Zlc6
iwEEl6H79TreM6ADvnAhc8hMmvbVgIsO8gdDdnlqPhV+tTsaBMD4S7JbRq6ofquh
jMWZrQ/XudXLSo2ytXGHwGUQm3VEPn2WZOLu17zdleDDbUa1c0xDkOhYjVRMCHW1
N44rf2SDxGXHpDNMK3Dkt8Ymay4IwhCOjaeDN/XBI+1TBvmZbfbYpykMUWM1UNkC
LIXRKXek7KfrMvXp8DRwG60QJu4ebK8j4HctQyCMljih7ZRd/gB2MF4gttBppXfT
EPF8jIybFsag0bMz3KONGrxPZcOTqoh68hhYtVeBFFMPg/3Gh6s+H/RTL++ewEH2
NtGP4qwOcOuei+zzLovxdgYUyZeIQ97mmkUkpfHxC5ko0J0MBw2ristQLW0hLVcV
h+boMwR24XKmw+azSsu/yS4eTiRBnJyqudiagJr98sHL266o3de2vRjSUR1oJ8NN
WH8qtRYtBwU+C7RU8kAHr08Jx3AADAKPIDTCwrib5ZDmpgJ4OuAw2QeXtsP4aeJY
W6y7U0aW2GtP2M7TjBMur0erGMzcUDkq7vMwJJFD+hTV8nd950aB69SThFTzKDGW
4FcAxiUUGN5wnJgYFndDVHWqlH/hQ5DGbzO3ppSqT5tcmAnGmPeTB6EiHkVoB2iv
6ST/7Ud3zQ1sgLx9d8Ep3iwL0t6nEG545FAJD12UYv4/ZG+jxqLzQPwjGVgXX5Iv
C/gWNBdQ9r8FFjxd1gwvgL++5SGyNn9vhcGi9Xz/7ccfQGtx5YubnBuq7oOyyktQ
OTl6Tyw86r3Xejtnd7JGtJ1s/EMrPmfmc35WoKzDuOA9TOPyYbIXqzk5Wg13iaBN
IuYv8k9lerXnp5OprWfW378hqptCiiDJEvg1ONX/sLd6exo5RkIh/1cMYk6Sbo/B
MliG9MzbdkbHGppOItFZNDa2S/DEyqAIqlsOia97HKmbNiPXTVeS2ygcsc7boUoH
Vk6aV/1n1/O8cV7Dlx/8nN8LhYs7IOn5fUY/vP0gVFWoTIXWZ+lbOwQrtkYYwn20
F/MSxeq6YIb5OKUUCRlOJj9kVvgpJMz2OLJMrOOJjzY1GwUZHABhl/9KIOyVXtf1
NR8XO08jR4iVzGUIzFBgu3iK6Ng5x69LBWVdzklKxsC6NbRfWYx3AnY74NWCGa+1
6Z2FllkUeGfrZ5yT8y6e7xcVMfT5eyNnA/NsMJf5jUu8zURQ/amCoB4NXzCl/CGY
fe0sI3+jWxgiKSA/mzLAkETeK30V4LgZZUiYz++ViN29zittLvjLSkNxWXzly4R2
pcpt7Y8EPtxiF0TzUuyNrQ3A68SPSc6DudjJZZrpwKdjtR6vNn+W4BtMZCQFick6
j3QB5NN25tDqAwiF2b3YCaGv6Zcl+H8Pzfu4DOFs+zWAtIBWNYMx2iaalY5iUIeT
CqRtfaG8SQEv8w6L0367VwzCRAUcjeU5dtNVnhVgGnxsAogCmmHBVw/e4jfOREf3
JZYVFU/0B+W/FXYvsJZ2unp66cTmi9iKDlG/vYhcS9E+c2QQ+EaTIgC9tTWo8XWj
S1JOv7DGhVS6QhknJkXgIU0nSpb6OdDa9HUjnhGWL1fkv4E85QJ3mgAzjwcbGMdT
Dkglr/0Z/Ds+ySkqtyI/yOVeiXTAspB7q19DeKByTWnHzUsy2K2gPhvtvC5zm3Aj
lFHwiCY3tm1WhmMZBbGbkbGYKAOVgYSaYWHmhIoRRXoUbtcEBkTBp6iSSTB//tEn
DsKIwLBm4Xn9uW6MLFfyqMnETVVafD20bZSd7c3CR5U47+POxaQiCFiDaFIvOymY
qOEdjwBJ/ITqA9CN1TC+zfeI9iZoFbdgsF1DZ1ibpHkGgmi2YOX8aFP3MVquoZa8
fSTOMk07cp8UFKi3f5EmAX85cwn4C37UZyBIQG+zHaPNndOpUcrw/O6wPBkDsTNq
q3veNf/tyPX72xK2dp+fyR9isGbMoc102vA6dud+AdbX1eWV/uNNOErlTkWXRqHv
99BI5oL/HHAkcA1y49bTxz7455s9igehjm+6SrCkHwYWzl/YJl7b8TTIv2yNG/+v
YkYMHZEoDk0ffq+x+S2iHleK1kq5h3WLB1h8BCklj9//kcbGaqAAObzNEFtJEtWo
DvsVx7e/K/ZTEYgQabATq5F6S4gWGQxEfojQVved4HFQ7czW0W9MTTDywJt9lCcp
/pCvHlxOHO0TachsISzqGhwo+W5OiJMq5yy8EUixC5L9aJge0txThkt9QCnucRAi
e1T9L+osV/GneYiz+gr89gzX6TxUlsqLZtjnCU/YO1GjimAvpD65/aXX9HeHBHuk
v9BGRgpbRUnhG66NeNbW+yRWxiFot2Fxj5zK66kMWHko65bUBkk6v8cSITYyMUjS
qbxOq9YiDLcE7zbEyOiZJfHsJnBvwhG+wXmu2E7KeSD5VvO6VFIxX3LWKiKwTUhO
0KmAyMpqe9XonhKTI8xbABsqgxtoZf8XxfwoBr8AFHqowgK2rsGVr+TIK99temnU
V4n5UyKbzlnqOuOxyfvquPFK5zGLTifGYap1/pF1N2gKstjO/6HqFq7FfrXSTjJo
LAcFAM39g2NsWFzrMLh/fWjOdJsFMUlkUEKdbkuBFuloJLo9ufARyBatNt9XJsCt
su1+u2YcqRjj5y1/hVMWw12rG0Ow6X+Awx5AvXvDItaJPWDKOn8Uc72XJwpSSvjv
pcNpgMp6H68QaX6wlPeilfA4VU2DuqX5QqKvMMCmI6eeo0O7MeP37Kqcka4SdYxw
a3DX+b8x/12E9NoL8W6g6y6VPJtTm04geqCAgCCMXWZ8lPpsEXsJpXsUMDX5gcnS
bMOQIwJ11LLWhjywC5kCXL3x4vUaYZ2IJTT1G5FOf2Wv4Ckx2JQ8YBGlu8VfMcRj
BvBr0kLFRgUj1AJ8jyhODdUMHIz3WpFYkQTP/GU1NvlPT9nDZChmmXE9Uz+VybvU
9rzO1M3R+c4Qmish7oudyveUljxW9nhzd2h/8RdkAr7KsCIZRgD3rLkkmshDRwHb
NPpZz9PBcLAF+C09/TxvUIBUNfhpmylu6PIUkpMg8GpAxUG1MQO8XgnVlM863Azr
9aIM2dGe80J9yqqRDV21NYQf6AGdFqjn6SGhbd7EfNn43Yp65V35JZ5uvpGJSSr+
rSq1XG/uJlG7egZ/QZXb2SqxUN0IfuHXzrZKuSGizSBkRgQslLrhojJq/0jSS+9v
2KKDn/fb6qp0/m6XvIm5Rrq4dC7QB76s8k5n7e66vEIyP+Uv+PhIiOGEOa2LPCl9
nEbZs3h0sV+cn2LqMiMohUJRHLK42ouSCVEf8G6TjMipgC5345wNSHYsiAhcM7us
WPUT3uPsGsRiX2ukyufxhmp0RUNQDnz1NA3dOpPcxgocgXc2bFWUb46BlurL/Wzo
2x2sP2cwAOvwFpXW6kXYik77pNDIFkpgqNwLG8YIrR+ggiCzf6e8Kajf/bqHLsPl
Ssn6zfE4tk+YK5yDrKGMYl8xTBiX4YAW7j9RGl+ci2B630nynwKCj8TK+tyHjnho
eY6JS+i56tGDnBBzYbih+zNX/QzB6xmxN8kAjPXUskN4S7pp1BxpW0Q0r637LKnU
3pQj2dSUy7jtOn+TOCGm90IaVOwurXsmO6PtvsXia8iZxBua/Pnzv3og+LRMKIxZ
5kysDISVI857KWKuzVlyecWSbLutgYH6DGVs9YPz+B31w0lEavNJwQp9p8KU1xm0
ydS4T5lr/VDsQw3Wk5gyUYvB6NlXS+KlFrEonkaQxEli205c3MYZUITd7wbpicMn
v5K1rJD77oJoesPwAZKGUHeEZzXu4yI+HGOjO1Wv6Bay49VInmzuHAszdSXDMlx1
k+FmAH2aDpFK7bCvmAWkbvoTUZcD32qqn/28sIAAJeKWpIAOcqywwXCvzf80MLSq
ZcfxQesKCUFDAJ49LHjfuWU5KDJ4woBASWDHXyDusPCCKubVRUkBu1wmwrPGZj9V
bqGXhkffs5w6uw5v1sN0Z5ieTbpk6XzUG6BMufsDVT+VhsGeduUAB0Yb6ti0OAz8
FMtFTR31QTHDeYLyy7YHsvSxpH2UoqNH3YclrNWv6JCQoRh86M8TKQ3rdSAllh1A
AuYx6IOYRzKP1SAk2pK79SkpDRidHRK5H/onmdWIQoK3ys23bjTITwr/YTOXatXg
TbWLzKVSifpx0rMr7tIArKlHt4vIdvPloTodCgjiLn9OUbmIJqwWJCMwaQEclQQN
OPGSennb/KxiQFvph3t5+047B/P7GtiZq+A6TQBzGHoXQVaA6EbbyXVbONzTsiHd
0BfLtTdDrP0tkISM4qqzksB4Sg4BfsnnwaMNXDZEuh+kwcEihK10AxCneyjwOIN5
sZnHmvs1snn2Wi/voFZN37EQKhUVYP78CxAxZF/I2m6PU48/vm7A28ThcQlstAZI
QgZxEuV7grqRU4m+apsUpCeUGipWddbiO6jdKjEcLnQK7L+689ymleiO54gY2wIb
Qny+NUJToDhJan6B5wxlb1yYf4n3MpuN3ZcUKpzkX+Gunc/UbF+CmRQAatAk8KIR
wsCYBrrrLY7IKwbi+dU465/mfTt2yhUDPvA+b1hgdm26w9s2KpiWtAgLCnmmZ5F+
aITQ6x/zq+ePcPiEBQievaQU2FtG51+d2+dJ4Bs4yXJxChbr2pB7wWVfsNuD30ul
5H7IgHmMr7sI5OFc6Gq1hHF5b+6uA8h6ielqDZpyNDeII2e3TZx7ZkpuQD8MySjU
oYjRPejt17fOsBiD5u3JWpURPHF9epyzgcpxzTIiRxliuPLf4w1fHo6ckGt/0tjW
ZSeDxyhEjeP7xFod3qq5KsSW/WzY+SJKjsz00AZQXeCWYq/AFAedMPSpC5XO9YWo
+gZESUSU/7C1HVV+OcmTDa9CxueT5zcXRclKWqv8QbSm6v+7/eufj6OfN4T2Z5OD
kdYB2aHY/FEHzTt6XXhWV7zLsI0HcRw/2KP5INqt7MTcTO2z2givQUtReqP6+bto
4CSGSiyYJihYOONlr9QCM1qU7uX8+0GdMaz/4YumJxsLvz3CYOmIEdRqmA73Ximq
ey6Vv5tQZHMPZxvMPoaZak7YGfZEdWtOzU/9v1Qp6xXXEujgCl8K/qf1cWrlPO2d
oZsx0k/ilj0gweFm2D9ZpkpQ/3iOw0wbg2dbmih8DywEhEefZ4iOaEXXgiMqnlvt
i/AJyMNvlmz2D2fTklWIeLXkXUeH9pTBCilKBNLqkkd4Jj5HEE/gvaTV7+5hYRQ2
ls96h6DEbl9ExJnplLNIaO/eki6WeLgFJrfa6gvdig3hSbzbQoRjL/NC3Z4b5dv6
bIlgwGxaPE9FZb+KaWIB/suJMu23wmMAlHeDWCpx5kXSlYmAtpk78BWKCD9g4a8E
zz//tnafBigKiHbygl2nthgBibzIOIbNUVeQgbD+y5Ec5Pntjomn7Yd/5iNsb2wy
JEmvb5ySQGZq+UXxVcubQSeoquMJJw7hgC9/anOz/fCOaXFy0JpfQJ9zroG+pC1n
9FFASAttRQaoua092b8iisC3ZxhHNdmlZZx8ZO7wwujG25gzoXQlb5j4RXms8KDi
KHFRD/bKxyAOBE7pjujGSl9IUiREkBGLD7QVvXDCLT3rM+Jwcac8/5uB+ONhi/nF
3bBsJkaPOlrAeaJPCj/9PN1WRujLUKobAP+BQ4GwPvvqrJ+WhaxqrzHNtmGyc7lf
FWzoK5F/BM/xupI1bAEKPVPa17zLldO/hColDawmbwU7gT3S5GJWh3EIcNPgFu6L
ygLbpyj83GAkf2AcAjrMCfikObMfv8FvgcGAs3onWSUJf8NzZ2AlvIFXO99uQ3Ph
ZvyiPXcGxXw5ZKsWMcmKhQaPFaVGEg/UovM9vbT5Hxe0s8rgdAXiNPiiEG8okj16
aWsGZduY7mgpRir71eA8RAonCyY3gdrWJaruAkLIwHvEPD4rdkhVgIExg2foSM19
ODw67K3FPyrUrOoqGa0wZqYh2ai8u0OtXKtWdcO874WWXqWgKhhWzmBWG3albQRY
aMZWhJ+r7Sz9AAkG5A+MdhfN6HNf4gjd9CA7sSts1tWAAuVfFwo9PThD7YTxLDq1
g6MvGVYU31EBa+YNW9+HQg7wTm6O+zVTxtp9h6XjAV1OAzNquOrCaMlbMvnB6Zot
5X4ul4yvH2oUTvfGnxXCyLHN0oSm8UMr2e99tpHDa788rcsckDiMgpCK2v0FYJv9
yDHS0WICLBwJh6mMwImYERryBDxnP8YkWGuNU6r3XonZeKYnn08gUY9vgZduY/J1
qMkqL6sT+fOl4h0Qb29yWV7FwkCu0sSHkCmKjoZqi9zgze/Q60k9YrcikjjFg4M2
pDvy5E3jUfYouh0u5SXOOoIXOrWoKeQLn1ivdtAaVCnOsXU95PsTAqCoICMr+/sz
SixmvJZKRh7n78Ey6PztU1VMPNgNjjheO1XFg9inEdw=
`protect end_protected