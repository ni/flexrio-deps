`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1648 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
FTGcP7VlpSOhasofAJvqcHplzZKt3U/IyJoktXPAgJGL+beyEHy5SkXLq9yBYpsX
it5q3n120RVJJvxpkYDObRSSueHReLHs98XPGnBFhUMm6/oZG5oYUb167NIlaJPE
ZbPScsX1RAPr3ugIUkWTglm3SXsijKv9EjK704xCJaQwVYCFdsicdWGere9GBokg
Y0E+6Ae/GhRg+A3v3HqScNorTLSw2LxOdCk7WfHkHBxlc+Ie2lmFQcq8E4eQ+07B
3+qS0ZTZw4hMHpwf4cVARJGQ7Giv6Uh8VRNH9j4aJcXzPOECj/TnGIee+/rrrxZ3
OCOP9Q/fX02cSfyyirHkD0uA78h6ZYFcz2ZQR+84u1rC/6PF2oCsJTS5BkNCvEy9
GwTtxo8+ZYRHRs//Yfzq+vXoCQ36psL2iYD1Sp/6GB6XbNtuQTYubMRodF4LxyIZ
1rco0/6AOUmxCDkwYONAAM8aXNI7s2cIRQ6fNGUQZI/6kIwYC3NVpxdtc/F+x1sx
Yq3zNUoZ2gl0u3nRa+r/N3aku3XTinqkPkmxKAU7PLgMb/LeoMPY2CtjHsDw2F1l
uQC5IUuLORLfKvFyIJTV+DBd15kndKumNb0egJKuZlv6Th383vOInu6W9p3thHID
VMw5Gvx+Nx9pV9wdpl/Rtcwh9nLwKxPs34NNYcFdTZ1v5YlwGCDCcgkHFSsEi8yn
lvg+3s468kJySOhWiWK6/sDfD/wHI3h6gMHcJ17Ojbrw0ftjB9RkvCzS6XE7Cty+
4O6hSd4ar4lArPUkn+FnYJgor0zjgXH7OL50iuspx0u7+oe+lKvi5mY8rExuMQj5
vhFHSAGLGMU/4/j4CAHXFMW6tnjxjtgf21ItlzsXUuyst8S9+f947mpXsPicSOj6
LtlE6TAWtIEAzwgaxGRpHkUso4Zy2knVD/wWilTUA+XzXDqk2wYkst52ssNc92vj
MbklIDCy3zpUkd1lJmjY6luL/ShJESrW4lJmVqM1s4vQPkcrLf9J+XWB1K6qywYZ
vv6REPTNegx89wPPxj5a8pzUu/pL54yCY1+0bocAK7kiAqKBvxE5FniPjGCjZ//X
A/zHWYeRLq4O77zhVPO8Ljel7DJ9PDHx/hr+634Su9kvlAh/6YbO6mH7yYXN+arq
s0TOHPHcwy7RYi0pkWL1+A6OhcLVWXOBkk9q4VuSwh79qpALoiaFdLwd2fKyoFV4
qd6tRMSvyWbJNrZ0Crx/B0hf4UNtv/f2DEVpbsO528zf/VxOSwuhYH5CsdrlkkDT
QpGxUyZxyurHOZgLk7+nxNB3N0dssMrNaqJRKmKJyGS9jOOpqbVlcuUhzE8V9h2C
NJMMhJ66serzo174vgfyqf/lkLEoI11RZmgcsf+lzgb2dYvy7SR5ld/XFiiV27qd
013TFQiKFCFHUjpLAyND1h8pqACawa5UdBxCmZLTkvM9+fRPZBL/jZKUFBC9tMxB
t9xOIhnHqaU7DSJwzeAsFXCcK9cpAuoww2IAC5nDNK5vrDpx+1TrhlSb7jiGQ8wK
26JblnQfQSz01l3X9uBgBP0pdeSVMkFjM3+FF+qwZn8SjIE3mwvnb9gh7C+Lta/K
U6qW5cAf5DgPcX72k6z8rfTOaHmCfLl7pzPW4xnD+v2cMMEcd/lQ/ylBdRFTwzvL
jtG+lh62x0Ms0bqv6njr4qXBMp7WCq2UU3f2+3UgQDaaJks/iQUfcmOqISkFd6f8
TG/NTa/XTGW1RLaAg1oAOE7qxHVlnWuTtA93SuWU539EmlruUf3QmYNjM+Ew9Tb9
chxHURjmLvHmC+tGDD7HIzgAbnhNqKKklK3M0gKYqpXwcXFyj4yc8s7rfJUOuIkc
V4XfjmqLfbIp2I25Lv4ToB+d2SeoOkxxP4Tz0EFIDjztGcCrEmwk4vfxFpsLOwqk
7jtWNXYbDIj7fAOz5QLLi3HivymvGPfqViewtzjM2qBSTu1vWsK3DK8Li3hJyoIr
VKbB7HCyGUtxuKe+qCtI+bSp+U7tTBiY5z6Tx5MJFCYESzkTX/kSMC6aMYNLAcAx
2ta6buVz7AkD/VuELkkxkA==
`protect end_protected