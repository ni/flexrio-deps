`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
hVdJHWSfELCmA4ds+csnOQAALbB3ps7EiTSHEDd//nts1r+JQrRE4d3bDPRJpiX2
Sl8d+xAK9BIi4i+3ruAzYvB6kuD7r+gs02Jsvd/1kn7JYK4xBxCjtdDFjVHOTEl1
sSh1oNiYUwLuwR1yKfP+xBhqxD2Dv6pCKhH1NdGilpJQ6cvivGkSunAu0tzP76T0
4x1pB179E7uIeRplfHWX03KzEBF+eVtfgXVp2W1BGjfAe43y1pCvNYZOh1+TY62g
EgAFgbo7pAujZxZy/YSiZjUr2mGp7o83qMXyusx8+rQ41D3X6rxfuP0RiId2pOpC
6oq5Dfkx04a1dk4s8w8cVg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="Sm9DkM+kBxuxXCFA+l3fFkxuSWV4xqRc4Nn7Ji3ukao="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
m2emGBqRy4AuduN4dffN8194qYvc9UXRqiQc56IrQYMiIVQPyh59I8SYabcDdspI
7AFHnvKD5YaF6tQfxWm+mlcmMEk2Y//aUjxeiGGs+RkKgbHitJF/K7nqg1dmKvDg
a/GaBCq4Bqh0EehlN4ntP5HxM4qcvSfh5m/Coe3drc4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uG91daMWA1mGkhgP3oZKMYye3UAomMWgG80HuuXg2E0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 41760 )
`protect data_block
c9NqBF2D1wSep1rW7utzHsk2j40aow1MnrccxUTvKej2Q1cyeDDbgAml4eTSXI8z
QYgCADtWi7S8BeChdv4B2VxKcS7CMq/DaQrOy1MKTfQzfAlK0iubmlTkljLy0Rwd
qPJokL5dgHaoxHhpf4hHti9VRBMmMBDKHMEzZlgVa9/1noQ6rVPJobNavrn5LOMB
zNSlZ5tPXYu7VIsa18690NPw1EhhWQ37qNmAEdRu+biZ+A3PMUvwVihvHQZEg6VE
1bSdFF0MvmyGpPPHM0medhu61P/b2tSmRjzrkgv5rFJn6kOxNzpaAPWVml1fVRsz
amQKwZrGr2uRS4Tf2x52ucSXhgaVo7SqJRv3iB75jXRYmfbQC5B4knMWuN6FNktX
qdRAifZ6YBMLU597r0fzG9K8+sfGhgw52k11dxiFI/ppThyyYvoCilcLk9xk3Q9n
ly72Gc2Tm+S5BRwxKcHi9F8/50PZzcmmD0AOiBmdFKWUlVTC7SDwuiP6L+I3aW2z
CWa48xTg767SVT35JxIZWbrRzT3rBa48Fklb7NWrvgUB6xGNtptNnpuis8g/4ij3
26tophFmVlKNfKRQhop/4i78CCttRrgrQmWlbZzKtx73vw8fje8AMvYox4uwy1LS
9K3vVA7Wg5xpga75MCP5hecjiZu9xBfoXps16SgTlIC5Dh1xVcMTJIjr8CC9siVU
YSxKqguoD1FtdtoDgzgwNXOj1j1jN+dxowEvHMQc8CHrrOgJx4TPNDMvcwVnY2mJ
Mrj/ltpz9RDwPTliRGLaRXAqsX+lgV4/RYFmMRtcCD5TI7mx855cJ3DW71wykWLB
ynUaPMUd8IMJ9XA6P6qT3LPL2KLDo9fD+FE8gtRVPmTkoZxqm36VMbzmS1w/QBrc
pkMVw2HVfkzysOrg3BsXVftID3WP1OKIhALEYidCcZFfKRdYNcBdNx6oXBcI4mCo
12rGrjFcW/Uf+1YQY1QOLdk1d+p56Z913IcDOb2XElCxQfEhNTNGstA1MRWCJejb
6A9/kRobm6aH/top7bLiRPUOiFJNGyN2/5wiG+YsRlZUAmDAxHb2PrG9I3kbVmkr
Cv+XZidHLWrSYhA8N6GVGQKhHCUUI4hPSzmgOQ7Z7tMnHIR0KWm7p7SmV+YzSm2P
h9ZE6sq7tGIu9p5tNv5dvbK66Qp1h2oT9dHXhOqPG76I9ekKWvwE75lwOL7CBToO
Y7GS18c0COT22/43aLGnZ/4s4AgW+YVlXEreigYcj71CnIFaVgMnXYOiNpTYcaFK
Db51F0PBS2Swu7cRx7A9oZ9vhdpGFo+PWmIXk3UmyoZfU/Zo/YQyQwIjTrZS6lXl
6wpQAsaquPrWJkdMVoG/KkN7oqZlJcqnN7k+OjMgOLMgZQeIJ1GoqNakhLHBKca9
YVP7pwRpR+QdBM5e1j+zALAJfmYoi+Lwoimij286DTJfqejjikSDURTa4UmlBCgK
kanHn4Tskf0pjjwlLfB1wfH4EPC5G4b6gZakh4odl2OrznbNJH6Yu2CsEWnV7vQ/
CzW4bm3HRxyHOfUJ5koqgQ9irEyLlYi47OYIJNBMw42sQ4J4SwBwLuPWltgIOUck
b+YJMVmOPuNlPpMZvaJWyD3jpF043dJ0yvXv2Cj/OpyAYO667nKjZrQGPCFBRcJz
lHRUCegEc0CfwEKMuELJBdhDBdUl5zbPE+MxVGh6FWQwDdZQ4InkIvvKXCRCxJbB
IBKgFcs3caaIaGYEQFTruIzxwIY3Z5UZ0frScR2FRsSCsjYXsHE4EyuahPkNDpJJ
6hMdQDWEu5Sf/ga4mU3WpqNKWkaoErUqxDWyocMwLMvOMdrOQYL31i2TAw5RRxap
KhS/N0RGW8nDeRZutaG3LNjv0Di/GTfenk31wRrOJzp6DXIFPeVCAadC21EsrHYW
egugGNP+bJYAzL1SwzbDMkWa/lkzUHAYYlHmej1r4gT6eGx1cirglPzTuUUEHFeT
QGvrcN6EAy3Rw/VS5H5JNMiilI7xXtKA+AxnZZrgrbqX8tTtAGu5ZQowrNPwJ2S0
+d3XUgHa4r6BuiG3jiXZJXALIfDubFjBLjOJk2JEYfV+qw4CW1Gnu0cFfV1CXhCn
Pj6+qZ6WPNVaOfzsml8oLQJSurv/eYzoeNM5oqZuOuo9HD3frpK+EFo4b4vYzPXv
rUifUEsEnMgZ+LY+4ZCvHrtB+5MbdPyUmbEzWq9Z1Mfh20q3qMfa7FMRGWdDBxrs
Rm0zjtVSrakp0jCpqjfZkzx7YhEYbkvs81eDyITppjU47TghSKqcdZtgLgj41OTl
xms25d7OJHru+dUcFg6XUDKuGtjRNj+oRNBJD3F2TFuezEXvHxuvbhWVoCHH2Zp5
rIaBpHqc04ryOQ0M7qk7E5/bJPKJkWq03836K0iDlsBZhgFmuyPLsunvsYOGW1Ut
VkTcXqkw4MNW1KYxnU71CgFOiL0h/fF8QSA4iTd1Hcdbqz0Gx9naxqaq7XAnSg6/
+AQT37LIfrPSyTYPcNfwKIUPZLUYkflf7Dpo3NQe/2e4cSLgSn+6PpfcRZNMwMiN
oh/pE7RFZ58z3ihMcwSXD3VLQpujpxuM/wCHB+roa6YD6oSLcgFfF2ZFh4u/FNWs
bqPWiiUR1mUSCFU8ojrFknWA0TCYc3aAIZicslVQjwsXx7sKDuZc57IjchaWwPvB
Ccr48bI/BzJrLbqnL2LBlWtWRBJLKq//C4wSLEnsgd8WBhzzaCZMxTFmgEN/6mnT
vE6BUaJ8fHauXXgCLCxcSun5a4Dt2mK9oxUxJlw7rhwOqwfYrgcN7BIPyKKa6acR
3ebkfQ4k4BIudRadQDHbRCipWKnrQH87LELnqlcMnnvbb82uGVU8Z8h0MP6QNkDY
gZVKOMzNFvLrrt7j3Lk24xDRUKPUyaR68zzZpFOFe9nznvt8+ujG3rGi26GiUlda
ugjI1kzZeo1J2tGBRn/9Rv7kpLrFiB2jVY3EwDZB9JCvCp9v8XrHvLDsTabGup5y
SruRowJ6V4iLxn91gPFB8TmTAKqjojPpk8h8drZoF+4TQDKFhCYvtW3XtJD4j7qG
991VSxoaJQjPFil/sp39fmpDqEEqLw99aoXI5B6oMcMtsbsI8pv3aYO9u02uiwzv
yhX/fpvozq+VXNUrH6QrWLEukZzlYyauwBCTBbOt5Qn+grn3yu6Ld8TSU+AnsIHc
x5wfPiI9QtAkp1Mj3vPwSn7FdL1GUeN0SKZLstlvY2w18Ruh0zaas49AXJLAFf0w
7R9TOblxxTNRSiLSAN0ejcZBdYzJstikTr84X1A2iaQt7867U09TO9lahrxeX7D7
Ds8CLyIB0dDcKHZXirLAJ9YsOwskEbK4P0QsAV9DtVcm5lJ3ENuSD7zhmJu8p1Xv
KIXP5NxEFsJRpucIQW/i+/S+wpIv8Of2o6kifXcxHIwT+WqySJmYKW7fzn09roWE
zbSQg21vCozyHA34ffTDIcjq9gH6D4mvdExmXYaW+s1wUDfMQO0i0Tf+ARVkCHMC
i6e5SAtTRvxvg855FvYYqa1fAwnJgGDQo4jlcUn7XsxTr4yepZFNgD8pJYCGMQ+M
DgoybVZW89rWrWXT85TGtdH++o2qzz+/WE+5cGJMRzLeLjBSqKVwSbV4SPctU6sG
0KORfQ2kLLynD7R76Rs6V+tRSmY+bOtGRdAXXxaH6/jISPZ1ZSMUokV/Q0x3VsOM
fUNVj4KE1pN8h6NpiijD7iVJoBommOC/s3d61jtKA48hMdk8OnN77e+Lpfqmwrsk
ItL8zJ5l2nLEG/X83mK/Pya9yu/fmjSj1juLdvFQYCnmJj5QPFq0Luh337zFI/Rg
e9sLqFaZbnrR5J2o3iN4Rbwc+7U5T5AUJLzEYPUPGT2quRW1HOoE9dPWOrgyjPmb
wdaDV1zisI66Gnp+ExgZQimi0DfKIPXYq/Q6K/8w3PXhZYBu5gNi/7/Ow00kLGAC
+Z6CwSdblglNAWzDRf4lvgd7OqXHsLQ6EzTHyZKFjO/pDCTIDhWiU+MOV7xt0H5I
aDtRzLk/lFHc/NPwS0VRHBBkDGTlziMAabGoC0xPZ4w2hO/6yTmJgXKdfksysrio
vN1iZdV/B0ESCnNtd8wTD9ZOgiyRUMjTM4BTk/IX35qeDoxM9QuSdZusHvVI7A00
BKQv+T923Mrk/RwFt1foM9exnUJ41X/SSSPEq9cClujER2L/c/gq867x+x0cCFux
+ZZ6pQQ4/wMuvTkHB1W1yfc143RrHNYeudo/SmHzkOym82F0X9wbLrhwuG8HvxkV
/3IVf3Ni/n2NopgT6hFMGEJZMKoPJPWNrots0x4uKUXmXgjQLVaogTV/HWmRQMH4
eUxxG5q5ZI+mXc/l6GumFg8GODknR+CrweYBX1I6AkxAC0yuX5S3Bo5Z4uFps+cL
hol38dM04yz6Edl3VWmDk6ZzrH1DnSWX1gqNzh5AfEQkVW5QFOXQXiRg8dphAJd9
TfOh7sLHJtZjwwHgBrDYAReHv0qrzxmgvAlWCASCz/E/O/+EotglLSgtR0BM8ThO
t3eygdI1QNsiIgcpNRYRusdw6FgF6xC/eDMg8k3Gh2h/XlOv63XlJjlckzgmKGkj
DfTPIEO0C7+OHK9xBCPWn+FcPmA1lYgWu49x55DNgt11h/cjALbWB7+1/DzAAK+I
ZqiigatHhpgNZm6z8aXyn8KsOMAA/2w8k4Lo/oKhMawliNViPADHkyYrCce1P7Lb
9BpuSk4jpEb22WflSQCVk+Ie5pRr9xxmYPskc+sPGWoqH4zdyAmT/USSWD8MSCaY
iRHdDkREjpL4nb/5/rGXC6kv+armgqZJNcj2Kx9cTboCLk8Ng1lQGfy305rRDIH7
Tcgv4SezT0FBFnav2bBTnme2xjOJzZSAgySCwYohLKNZ6cLuFlgkA95xmqXQA2Xn
QrmVgbJ1bWBnhcnD5YuhY0HdtdpZhScv/JQHtpIQRWjkMb2wWIqTtZFNvQu4wabQ
ANKyVC2hkzvWROIeQCiPYZ1+xWE1gSz/KIwxQNv/YxrzSxbHkh5irIt1DLvbKMrX
7nYqGriwiKk5foNfKBXIalRD2mJoPFez0yBAeulByazKAX3wv+Pq7TPmWTPLOWcB
sG62zZUL4FGnmhUAp9ZAc1YifuoXcDntA8CjVZ1FUkXqEyOAwwhPpW8p0gazQ1/a
by0C1jl6YUaE/MPK+iRNmvaBcIrWHsNeIk0qRHFMvwGc+oCgKds1+K8NYpBTJHUN
xTXvSh3fSkdL+pflDQijT5pqIoIiaRulZic766lRVcfi5Mt5D64y+ArlNSbrcgL9
+CZ5PoK2He4lDy5k0+2Jiigd4hU7yLS7fQw9OJa3txW/vr350SjbI5kYQjVM/LbN
ZOgBFqN++M+3bdxA2UoVOp15fZQMPSkJLOM/6A0+eOZ0MIdN/V2YEDraN+x80qgw
eIwHfSGSSeHMXenqd8DA49GglW8n8mm6IfOuCsceTujrvobTCAPOcFIFDrTlkBwx
TAGRZfieAqo7bTv3WTCLZq40M1fYl7pu+46qd3OkoXBhrjrzyHXzFPGaQDcSGWiu
R0XAc0S+SyVmNxiuxZiJqJCBr/+EhpY5HL3t6kaIO2vlOXzwQ3j6HB5fPFdcEsJk
SnJjL3UhOBzUJY+7RBDe+sPAYhpITLNFu3oKw+I9OU7BAKuWHKQO3m0KI7u8IAl5
WHIUIHwnS08Fq5eM2WWSH8icaEalliHGv9TquPzmDq9M9zCaqCIGATBgHnopvrxx
t/7CIhP7hjS3Ubsu//uhDSnaZZ32qOwwHJZz2Z36YmtjaL93F7MIi0pS6+7qg92h
EuK/CIQGZj/YU6B7afcml0e+cJMqmuyUE4nMNyOq4dEHwsPJNR08kFyfbEalVN++
wqh9rAO8kWEHVTnBb+H8Jm4A3E8YhDm/rQBOkOeH+8gr5XlkFguf/EfRDUSpVzWf
fKRHDyLHmP9B6IT1TvvftOpz+Oh5YNjdM51QmKmnZqcV6H+itRpJoNyIXLejhWFI
MqcXciPUYKvPTRo+AFUVjrYquaWH33aRxk7eOR/ll2Ca20y5LfmQtKNITTl5b4qa
68ATqLYk9YuxEcbSnDLCDAeX0knzXWMd5NwZGz/S6nATU+0Ff/CFsjjwir2g8YJy
U6kc1U5Rq2vJ+TYrqGwvb+afnjbjT+UVP+RbdTrdzdz/T8Yq+mvu//svBlFstq7r
rnbZFCxRF+ig236sHSrKbYkJ7cWsuRJYpOQdZWyW8+0n5bKTjEmC16nOoFjK5T6y
7SvIwRzjoIbtcqGgd1UrT52KffLyrIcjfBhVdU3tJjjMhoJSSR+lAU2nfurSBe3r
Xqa7wKCs4RInO2VXLC4RJFCLjsuLvnafsfU8ruNSyhanumeKNmOsJ7VmRvmzpGKG
oQl3TgFdjoXB4GLIFvCazGDsG6ceO1KYXwfY8hMBV0CfnKTYPH8b3N9wwan/+QM9
t8c2hBna8ckUFCd2GgKU8EjVZAVbGEA5AKgNDeDxFH75lloftC++8ZQkAvWFRSl4
kBB16WQdtDCRADHOkYt4mz3pMAITL2FrqO91tYYN9ytVPSRLdXQb2NYVxBWZ2s/x
jIVnUNcgSB4AD76/wLDHhH6ixSPFQzSCq9yxGjpcvYDP8CStTg0ZF8YnneDDMREF
VciaeuVevt4F1sNKan+apvh0v7eVQEwRzOjDlN60l7up436JN4l7NCljV0lk1eVv
ZrEYdkIEu6UaNIC5hdeI9sYHCNf2vysCtOWdyYEpoUFBvpEWKgUjPZ3fxiSfn53F
3DAxzNFvkoQPqghdjMbuWxrv80xL1m+vMktzSMmwAQhOQO5+m0wVNajZsDQIoo1U
q0Ic51kAiKC1jY2K0V9zQo/iBhLR8D5nHDHifhBH//dQd7lQVRGdkuUWp2splrjS
RHU08GOl/mgJWKezzfdWuTB3kNP7c+G2pxke1rgFGgVnS1OxNklfsMwlKx1yUJVV
1GU+gUmQQeB9O+UpDyprTrjzmKqEkfvyncCqueu70qKWBzeyzFjM94d/Tp3lLgr1
ugV9gXZ5+UoUCkMORJm0oSbFwAkyScf2TLKv4ZwqGvJr1g3lHjQl0WSJPNejAueJ
nM3SbRepfrfNk1nTiFP66nxFQXem9EZlwb1rKgZwQ9srgWPYoXuy6t6OtabVGuum
b6b/feSM+g2rotulxyaaAxmoP5oRYkwdRMm2aPZ5c+9FRjZ1+xS8Z3A0d0X3weMr
DnZ/G889nZEbt1Emd3jqC/O2OI5nISHyWCG3qCBCCUbDzhmp4vmhJ6QGAT2pvPET
9m2+WGCZlhPr896jQrzJ9A2cmIMmC9Bl4V95WgtTF6Ru4+U+IykkMwgkcVrQPvcE
qNsbUrXVEs6HVqE0yexsA1ALQlLjZ3dob4XUA/pF2vtWWM/b1SpbrS0NQdNgsIyx
S2my68+zTjgS0uAEHRSnAfyCqlFiCDLkkN5NCZ2TdcMPazi+K/8xU6SPYsYsxeFA
Dtj5bchJpfEou3C09zLgBY0O0RoGNfjkA3tlQflSjyRe1tmJ2nDWCOEzv6NKHlAZ
lADFEGBedXDTIKAo/JiO4DTqLxpj8fTMdZQyucEDAHgGgR/K6LOhiRcxTYStsAVq
B43hgJu0x13NtlJ8OycDh4789WqvTOv2Sx0tUGzOgwT3FOC1WqpwXVbcHHWj5Wr7
GcHC0/NsBqDSaZieWSRGmjcenv2DMhgFzOsrfbC8LvTiZrDkLUF+uRh9bkBwsC0Q
EYqxP3NQhI+UG1DaELI0s7U9MvEtTbwW0kg6OxkXk7d/AyCrQDYk1HqgOyRLjEAq
m0BBSbB6/8lYIYK9NMPgFpn8JkDmzQpCFNv2CA4GdadAlVG/hwkuE7UGLd8QVkgi
BFDlhwJ4oGpPn5P7rKwyUfktbBq5nTDCKulY2gwAt4sAPW027KJGGewyhpFAYpUq
45XX1zg97bTHndhkgd5U38iHMa3p6wiyMwAtcoFaGtqT+ABle/erJmvLqvSMbKXw
IpOxfzbX3Zyrv+31mdveo8bPFTiLXNM2Cu2pcu3sdpMzkScI4w7qbV+FDVvgmMn9
2xaeouExCjV2SRkOkw1FiD9cJDkyj3fYs3Kuw88sEcvg9doaFxESp6Oo75zLg5Q7
O4h/yd6t2s/lteYaZ1V0yH6BFEtydHwWwhX7rgsnUT5ks8hucflakOasG8LLxHBA
wI4svCuKZgLIWzxecV2ir+lRP6X5uGDfeL4WOBwhDOEXFndWcWJ+wRwm6RjCdChL
R2bCQOT36qv1PkXb2pmphfyhqitTqQccnd+pP1Ix+UKuBmYP3/uUJXy/k6vGVji0
Yyq/Sjlvb23Ya6Y9yi4HazcbAG51LspkNukiE8V0mjuMg/N0V8ikWaRl/fTTpjnk
wRlAPG5f4fkG4Bs2pcE0VWZxa8ZbiwvoFVx054uh4wChskmptSbY36gQ6gz7Wq8t
StRyAMgHtdVdazmy6U9U5oO025PLnHmtC+Y95eJqdHVSEyc9f0msCNKLFTHthUz4
q0UppzejFgD9RN0c+dvxV44B5gtTM4YhNylzPkR6f2SmjSWItevKG/kTfnixAyas
wbiNSy/6wCnwN0l8L0iPgXGscjNO8w7/jrpHMmdJ1gSdlxUx2tU/eKVY+MKyOvqm
JZS/biUe6SQ4hl47//x8A9UcKfKDnQYaGJIbwIY/DqekOf/TEhuET/UtANcj36ho
Y51LMo0PzsaS8szWx58cg/XYfQ2Jh9bBXxlsfIegq/sf2vLUk1wLj4/lMDFafxzi
LdTeJg2vF+z+70nwdLkJ9rFrIgJEq0aACsZWYGBtuP0YpEIkSgAjE5HxQtvOB2ph
A2KaIjya8rcHDeEyJlEA1qqSj+YxJiPbve8vhtmivJPHIFqK5LHkA7KWMNIo7WKf
ukk1/XhBz6AMSLDBwFAwYDUV+IR+9Ll6w6Ew1OLQqaW9kfItgDzHDn/xJVy42i1C
ZmlVQvpo/qiBqzip1ecBacBmM4lS2vpjZ5eFhSbrViLez09IllOzoDeMaCrkbmQl
2iT24U0KlcUIzmiB54ku3qam96fUx2NKtOp8NvNFqCGt20baCFtsp5Nrn0S6eS6H
4emXMAubDp7MzCf/cmMYG8wBW5h+0mxVBZD1+9Q0B0v1QBIFde5ULQzzXc9aHnEk
H4zug7w0/LTCf4aC4Am/jAgRURtqY5hSwJxOCtUPhrwlK9fj2NDVxNB5rRtjx9up
Z1xN94VINaF5bBQEJQDaw6dw92vhQmK/8ELKSzjc4Y/J7sAyLBoYC1NRcDcWNktY
axRSnS+nDl6W5h+s4uNe500USSk25bw6IM/94OiFcKTHXl46E9j+Tdohf5CUzoZg
ICRSOS7Yn6yEqKrOZa8pwd3gMrB0/6MUSzBZe/+6jW3TcSRyjMNj/uars5QwKN+l
CwhhfdjNOxk7We8vmbaIu+JJ7gYdFpmVIi742YIA+EAao8FI8tkpvJZ7BnE0MZR7
l6WcYl3NR/qVxROVniArRyWi0RDH2jBurzziWSt3FBAR9VreFhOwSbwffnjeetrH
JB2Q462NRIlz2e3a4XG48pZXBnhIlgZJCgMaUgAdGNB4Jbh8rcwr2yshsWL2m5RL
3Dom4zPkSZquXWpdqX5GiqDfE7Gmq/iQ8izcxrrz29Dvmz9yAf77Y8uFTa8apIa+
LS+iEp+Rg/nLkN5wUNHzASe3Hbbw8M0c4B8Xl/QLQrBMNCtoeqwgypM4yzPwomSy
6IoMhxqT6WNawO3LdP8Ay6T530Es6jMKr+yW/zZYHaWdVhm7aaA0MLJJ1uzMZqwl
N2LkvFatu3oPsMuWCRe/ZXHWL2Vzh5zbaVTIR51EyTZ6IaJy54iqrbQN+6OF2vpd
4PFml+hGySb4+3NaHE+j4d0v8wKuBb8/Y55q9G8sJ6f/D0Ib8uzMkColWOg/yjfR
IhbRd9z9ClxrE787fg9tiRkCqEjRy3Y6hJmOT9PYGwd4kzGQ5hoh2IN3xa7ab3tv
TiPOYq6gBgis5lr5F2UVuDhZLf/hxYlm3yQpM1tq984Mfl9MzznxX7khbB2TDTG9
MJeWp8Kp7VqaQZ7IfEkJ2Cs9D+sIoq/iHipfUA0rPv1RlyetPGE9tET0CvDE8p1B
Vb2XDeDlnu0Xf1SaZ2MO69O+KJ9wraIX8WxwEZln+KlPltXuvOOoT11BXhunbqRK
xiYwq3Ztxxa91KQvh9SFQ0pi5rOzPcWg5xF78cqYDl3H40AuHdTOHvy491F57yN8
mgxrPNOKUIrJU4akjd/lmeIW+Mr9njsSAdvqReYkiAUaflvaeYaddkW0uz9wz2DV
F6jGCdkuwCzuHmOiksFmB6fq/DwDLVsL/5oIZHs/5op5T1heuk3de/Uq0vFxAzas
M8n8qj0zInenuMTe2PK5Sq+05p/REf1L3m1VG7dHFRUeuM3r9+EGBnalBp4RhiU0
LAlVQjtF5ci4GwvHvWOZvKjAdhafc/c+aPqF5B0m3nVOUDg86NXbuovwaR3faQJs
R1cyNcw6RhG0Cl7VmMfabc2m6XSSOdxugAGMZs02F8BsHiPN+esP9d01F8oiytnL
rH2+yJawAIPfjTzWdwvBGQjyhgp+zAyTvh6Wd17roMmNEdPqfM4+6lqO/JZ8kfIS
jPWNgI5qF6m6u80An+wLPdRwCxRcWbu2VxRcIA+gMmgFS3iu9S1KhtNu6rrgI9J8
uFhVDZ0Shf6yjYuknxFsg9QNSgjMKwbNLvO8LbUHR5+glwYSgfs5861bduApgUWg
m0rgyuEkexjX15oR0ICoYKnsvKVk93M9Ct1ay9Vnc9375uyhNlNE9qnBZ+xRhSUm
yM80RNylelUPVjWB+TdA/VVFqZ6ggFMAnaFPWVIX9vT5sqKJvQ3OSqC6Hf49awE+
eRgYsf4zkq1pH1dUrsymd4HUuuX+fZOa5SKco/gFQ+Qizm4QB9ZkqVw10tUnKpl7
nIYgysvRWcl7YZZJQ1Lc7Rw3A2qgA5mwnncNxZlEEOgWYA+3L7PVfxwb711L/OPU
CegB5pqZOLIy9kil/RvvglU5CI2gMtKfDLAMjgz8CgV4DBhJsTrHVPv2B+0LpFfT
/DNmE73hnVEBHptQ72V3tVcJgCIh98t7d2ApO/6iLnRvuoZPPzpfrbux+kDqVAO/
y9F7aPTYkgCY6tG3i7J3QMiD7WdLey/G9epq7brUFzGTwi0KL2dcxuBJ/1ZpXSfj
fvMvoCz332KNcR01ecMel0ZtDOZMSMrlDwBfeoYjNcPnjx3lv9GDOkD8peS6oPlr
087XzZMloV+r7X74UL1+z2y+7fpERJwE7fkjJYkXsTay7E+9vW7sIJtmAXG5Y2xH
8D9XSU+Qz67uf8udqcWWTukU1LolqUrqN/9KIOGzZPHrN83xZ5lEqtAIhttNOhs+
YEwIhMqhwoW81fbFK8viIqV9WfXiq3opjugEatk9kLXRJYq5w9AqeIeztP7+uQ0T
HkqbGxrzqwzpGWiYfX+Fc1mUYOsL1wDjnFoy/MKf79FxtxYlSJos72y9RRfin/99
az6XX+i74JOVcC6/Myk+/n/h/TtIfpKArqDLfGbUCPlTMoAJwusHSA5AGa7bFshv
pkjccsIgkKFpgFTuv7g+VQwlBapX3mqn84acsbl0ho8FDII6TJf6raL/fuqVG4gU
jhSdKdOHuJFC7LFeLr4WvwKAZoSwI6dfteTNwA7bV2lY5jE+6mxjwbJgAfqZy9D0
ZHo5EXgspPSampj2YZo2HGQL2bSNg7zoCO8UqMxLwukL9Pn3d+PqrmXVjKfhIzlI
0JO3oqPbTv5ZRO+IPayWvRIWvuFhVChY42mmqigdGJxryogrSo2RnEfX0fmGOu3X
DxqydO8aAsUkze3Ek/IUIx2cRWJLgnSvBe09QjAwsJdnxxChpcDBznSgcUdToD6j
FPN29p0vKARR3lMW/+rTb888zm4WeUMmDduYymcTzL+tlbv3oWAe1sq/fmBF9anZ
il3XBNaaWPQOvmxUZEzGc0u10YZxn6OWSOPhWAPKL4QoTHBIy9G9VMkeorDL7mrs
LDl9ZkbGubDbLSPUgd648J6czqHGOE3LSzd/vtrGU8Bd5TmQqXIYQaKkfFH0AzV3
5VTT3bcC8vRnDlDYkS2v9Z1aIvm9VWwYcJDIPlyzgXhC0TkFO+lyq97/gUcIsDrQ
1UY2qLeITArw3XLXSC+aZh6Pt8+yI7JwZF/2STcrzL5/Uziw6nhjegcSxG04yR3h
NzezNgB0Ay4X7UhVfvcKCV6r9oqMTvHuSAhL2DYz4ncLI5QCbjq3qmZa1wJe+1ys
it09MNYupWwH1n4s1OHeX7y88Gk9famCC61eXLcEN1u/aSxU2D2zrXdbcpRxR/Vk
/BVUwbhXSbg2K4/yKykOW/GW03KbjS3xDYeir+4T8IScwiqdHtBD+xkmw1sX2GcP
YChLDk3o+L7UD5gAYOJsC2gLboynm21MSv7L8P3soIIEFo1DgjTmlzazyzD5L5tN
Ko9pI3YH+ZjHO6ts3L/iy61HvEzlcuu/U/Gd1JW6Isn+tMBcEYDBKrjmReUXOlj0
PdBB2GwOVhDX+FlS5ng1gIJk0RKBoSP/ZbfPylhL/85JAySr6OvawGYcxAYpWMob
tHJd847W5lr+f6imMxRGHiPnvo0LYwTE6VbDr/1mhBDWN5PpkCxSX6If8+EHGHJP
MhdKFMQ8mhjUH9pjnwkZC5fRzwqHm8dSzKfGndlTeDVHBbJY56axbsLJi3B/UYQM
Dx9w3FsXXwH3m77hM4Wg6kzTCitapEdkBRQChgUp933NkN5tB3JPGYfSFU7tkmUe
i2lnJog3kcE7qjfO9gb6R4021jMI10kNOMbd+2Ac9Sz+UEBwbUQOyv2vLjPUQJmZ
dFyqUJC5qOEAW/ZISooyR2kUMViqWG5z5/2lbpsa3Q1dT+fG7YVGBI225ELe6q9O
38OEtBWN3or1TH+gLd0rOrAk/sjHvUAJPHGEHLIWupdk6Jx5bdgk2U3FADHzGYev
53en8FgBONXMVToS1GY8hfb78JsInPblsKDYvi5c9BeMJvxDA6VWFCqM20ZfXvDp
iV2MvDPdTfaRz2n3jJO4BlANPy6gqRt1kM6IqT8qhfEhSMzUX4nxY3QuVuxfGrwU
Fp3PJVzwFHIZmGbQD6Hr4x4ObTkLiL85PhTHKXvU1ejNXkIZNfC6hzTxfJF3oMWH
vqU9Kv1vQd+Wim4aV1athUVFQ/ajNSC1sz/ha2SSQJgaWdwYcUohRxTpfhaMlHg8
jZyR05fE9z44NBqEdH70Z7SKfagcaVD8WH2vLPPjUXfcOQ8vBBua0iDTYeFyDTek
pQvv2W/ylC1OqfV5BFuWwxCacwFnh717VZzqDd10pGEgLdcmAbbmiy8dW/ZNJegI
iJ03uVcXSNR24MpR3dr9WzhKQGFv6DPYLSLdWmTuljxcRcf3Oi1X6oapKzr7DoTN
TjMQS0EQ6BN3g1TsE7LQ84bqHpDUrGWEEImWjSal+NPbba6Omt8EXrsn4pc8BTSE
YDxhVzRQ9m1VvuOSs8L2vIOSmHqxZUCx85IeHqf7VP8XCVQExKG/Smy0bLllnXyM
3dUXYjoUiDlQEFmyET9GbdDXek1WG8HRvkaHxhAxmQPJ6bl3ApxaGNd/hqd0N9Dz
YGjausUJ5r+/PLUXF7em6OUg9YA3OTgihJL92zbR0wSsvFZSrEsrgX1xduxZIlPh
pgBmCz+tH64O3lpHtDvfmfLk6JLR1euMehCjl6+tyZXKFs5dQ6GGzM3H98M1SgZt
1/YTYnQ8NvECavp2TeA4uUPGq8pWpbmlCsdECnmeIp2gwvfFT/LpMp3fXuip9kpr
Ci42R1eBK+PVt0EcOySqV4ycWR+1nHvSzV13s+0+ANaj2cLaq95UNsMYTrun/Una
dxAa+Dqo5tiulp2/+38oPbrhTih1JItQdPsdsLcmVIqDmtwQ+HW5pXjHmz7K+tK/
Qnf/ZGtuc1wIDtLq8sAwdZSjGQvHR+r6Z+6T6GzRBYqBwM6raADjl2GZduQuG+2y
UmSddH8//QA53lbLUa7jILtp0XX5FG7EDQiDySxYhpM5wWPGs4LYbGpQ7IK8Wexy
TD66dwdOH8VLH1QWfBfJDvBUBVOwKGwjRM9QY3H/xzLGkYiBqreJri0HF/Ji3x+G
ZBti+kOKTb1aHdhanpsLPJE8G/eRvHMkHeJHFpJEDJ89TNU8uFzBM6+ieLFO4w48
FU1c5dLTQFNs1h9hmiicNLSWHO+iOcST3m8794VLmKXO7hMsruw7EtZLR9Up+c2K
7KpUuzm+USiMnLJX6c0z/r6w8LZv3ANR7+XZ5Xtqmm5qj9RRBm2/g1elN+MKyetz
tjQ+vGECfY2QB0n5zzGN9v13spoGtdOMGMp9Wkcbi2HUw/Iuwkrsm9n/LQZvbdNh
Ft99vbPBe5rjDw0bCIyYhclBsWKwPLMHRu+O58MeaAnvfzFFQKIION4LHvzJMOrP
eAp3EV6Vsf9iWYw35T7O+bAT0e8sPIBkf/Wmb56Fp0gWMBtYPK0s9aqVVisXkeOg
dSu3H77DJ9HnBlXXIZ2+U6i7Lq2LP4dWbH4rzezIPjUDI5hTEI0PqVP6EuyPQOru
FZsxV3C4vSI1t/ffNV3T7zDiJbK/EgU7Gqb6w2qgK0TVM4yL2Wd6lL2YLAH2GuQm
cJo9Ex//y0XMRuShiN/M8xk5j4Cgfnyem/MwHL+U/HQQL67l2G50AvbVOuQX26hp
9OqJlWAoxziuKZehoc9kxYuS5cfvQUHknYNvInspDrygonDNh4akFmw9bE4LsgDE
MvKyPEtbm69F1RwfOcBcfPvQyhim4puxOH82on68rjIQkLNAmmKhX3fZ2tw93WrF
gkhmm4nwIN84nXlTi/c6dDmRqFLt5j9MJFsBT3Ssleg8YNozn0MgeoZCm3e6LLaN
jGocmkpqxNJHdJIEiQCfhpAN3rVnu/xAatC+ehngcwzfgrL8/dRyfeRW1nU7Kejl
EDI0ZE3XVvT6zH4VLuPyh9kbgS8sO8rx0u9+ad2C1egoq7Zrk0YH+NLMDo7jYneo
+hcplr0wURCuNf9XWC3fgWBFc2s13r+2xCNDlyIBxRTV++S8UThunbi9cSZy9u24
DAefGyz8R3SQPyvZVtPBZhwKQexLc5WpkdQZnBuzif80m8Ct4fg6lkvz5Nmh5VLc
pfBUNZc6VUu4PvEdK+k9BtSMC2C+E3OfAa5jKn3AB/5yrzaqX3Nr4HWL4LXjdvpV
Xt1BW91T6U5hZCTlRDFjOEAvsCDGAv158x+jxg2kXQszemshP1mQoroSCuZH/7N9
gslvun+hWCPY2spJatVJH1F7sPYW/BjUcyBMOMhHCsQdWlfm5F7Rw3CrYib3Xsln
8B7Q2wAEB/LyWpVgOHyZ3UTqi5mqgSuY2FCtx1m5H/Lqhz7Y4UEtLB0OIN4r6Bzn
B78GL7bYm0zlJjoc+FWoKPxD0VFgv/RXk7UCAVGRv+kSn5X7lRobG331eFvqg/Zb
eN3AyXY0xLS2wYRdNnZPsyaPnfTj0KLpJmA8xRisa1lQZb/JeTtpW19ANdebiG8X
QQ+x1tD2E3Wfsy9l1bEE4c+c3mViz1blcOmoI87MfFZC+5RF8RwrPGmgPTFDUlTe
OjSKKaGX9iosvKMCsQjigJid6PLjUK4FMoKOx3m8au+aovJtOECoHV7o3ccyR0CG
KWM5LoIjbC4OBpgioVvMA4dR0AzvnDoG9/LGNdFV/x9Ds92YImPeLK/Asxo8QZiv
yT4bBwTw0mjkrRaejead40HcxokZUaMASEZ4KGqBOMm4Cp052Zwqdzj2Be5FhUYN
/yURH2BxYW0UrEjms/NJBBfRlch34rTeaGIPKofjiayjQt5DGFMU7P1PAspztV1s
R2DSEYLEu592XBW5cJ67O0KaGH/M8rxV+0/p47r0gzoq1pCIu11H9wvkFSPBconL
Fnvk0dY/kw8YMFXGwKrh0kHFmxf00T5hZFx/QAuvHJU3c79oESEMZr3onhTQS38i
Mvcc22FBPhrRH3ivLuVUMwPjOE/ujfwDKot+jx5ZicTBMzY4C6LwuZ3RrHr6h1hC
z0K4HZvYrqcp7dskJA73Oc8hYNcTAtv/yYbTlYF4+G4nxxwJQLlxivVi/sOYo7Qt
QGrc5czQyjAIYZ385B0gkmsnnkwVz4Pd4J3DkeKUUHzJWfvaN7Yjj5J8OVwTt3of
6POhNxUnMloqpe8kWW62z+J3FQ1+Tqk8t7cCvIuEVeA462rJtf32CAKJtRTqYDXS
2bIcbwmhZpgS8f+PGa3yCam4uPY6AgTTERo2qcxmw18dFwlOsnTTc9TAvw/aMAk7
lzh2iqN5fUegalAbtXLh3k0mjNFN/+VJ+OYOvoWplynFAeSp5Ohyk/IuRaiZKSCB
HLjzd4yHSyvcjXYmZA9Z9RgLFtlu3sS807GiqPhvF/Xu1tlWIWvsv/3jbv8ZsBtU
zFjid63OWHNFa4e7AOZe/P3wdI8iphA6F75ujQCRC7kjv1Z8zjBzO61Y6wPcshxL
TS1Hcjau7uBEHWq7I9b+re7bMEbfqHUxi1l1c9Ldcsh+/w7biBdRCncl4joXK+/s
OBnjd3izgKZPxunbGpGw5XaU6qTrJhlAIJCaJuj1EZOBRsDKVdByAp9wQ09+FPGS
IDYl1or/zP4U9iO2HQZOz5+H7SJHYh0PsohH7IImvR1TPrWU7+nNNkqiDMj4qD2a
lEVA1e+Otx5BrKoK2zd2fveUR0Rc+of/mOipIFnlD6UxAjqbQEpjg91UtYAvC6zM
vojZg3qU8XPNExzl1CjjKfGc16B5HZGElDhBiSdneVFz3MKs31GCU7QnSDqEibGb
j76eavg4zkq6dyE/M6M6a320vjNZ1crqgFq11zd+X4Zg7x/HlExdd9t4k50Uk9Ij
btiqWsmzw2DbQkcL+8giL/1d0h3Wnp79Wz41Z1nquFQrYWChmsJyYIHoPzfF4W77
uS3j1bdfNsMUv3aGkxkCYImkN3NsoRK/eJyV5Eexjm3JFg1TI6t3rBPWXMv71/Gf
k3a5emmeoLa+CZ9Yxb+1sT3eHZ7lyV4bj8KktBSw2mFF0paJ0WkzSsv8DbMyx0+S
aUkE4U9fynXdiypqhsZEOlzCKEijKc0K3dQeFp8Yrq2U0gu3Coq7ztqk8YfnrWgN
BW2dtexxxaB/WQ8IdQbmpIMVoRdFr73up179upaSbbsFCYM+IZuLjJTm9HkKoEmJ
Egejbc8FqAMZ0wmj0ocRI538sWOOc8svhJwaDZuTc+fGLwaZFCCo6CNnPJ1kIPtz
18U9izTZS1rHXSdfztn2gq7dSTgJJjQ9gQ5VQMVw+AFQItnQhNJ7VB6s2Zq+GE8W
eTpsu1X4ZAUBlcS+8T/J+VGYdx8r5VWSAOFAlxmdlSwrOLkA4mkc8x9Yk53bI5oA
R1vbTnr3gQnTTeOVmx1LRU2QxgLrbuO+qJkjKD6D9y8EEsPeXRQ2IWYbDfoOGUCB
bYkUBBrPJVjIGcOR7wjMlNlzXV3qaMnJN1Mm7YneIFjFelyOnueI4gy+JmdJAdTc
N7VTUHOqsecqRYJWnP7LGOIDSPejFJk9j1eg3gTM0bwfEu9Ouzepi+Kgm35EXa25
8/5VL7Ib/CkewF/sMq8hMmFOF9JnPkwJytD1+hD51XdL7Zu1W5TKcL/V+q/7ma/B
yOJzC4vLzbCeMB5/Yw+mF09mFCVJ7F9dkmzVffB0WH8YQlfcVDChWcMKSQSFMEaY
h358SzzRA2l17XbN2kimQr4JJBXrHKRu4bwq+CzhcEtdY+s7fJU8GV8G4hmg1+aA
kedKn+PTm6WH5wm3a96KFw5iVl+RGXp338W55FX2UhPK+9nBDExnwO+yDqR8RA5z
cjNzdTWJOcvAtmbFFQnV2f5iIn+izz3VbmAOFB5I7PrxU1En07nKpIpIEnX1s5ii
ZHk91iwE098p82Na8gpM1Q9oRQgUb07YWQMGx1ZHWPzc7RQtpesLNRV5mPPvc20Z
rzO/F+LkbidkKPkZbjZEutuP0luN48XY3gEDuWfQjofwLqgvGADrHguwcAg+0Bgz
gfWIRwu+BIQfRHhAnpqOBz2Jxeu/tOC+uUXKgO1irZ4ZTBeNGrbpGkFwVbKC5i+s
yNORfbkG0ZG74Fq0yH2y49sn25hCAyauSHLdpr2P11M9aPO2E5Mvj1G1WErEiq0G
g8ywDfoOuswqUqPBXlLENHLUJViNrhMzOy/cJTZUJ1HUe8gJiRvO30HQvI7hsHqF
r5VLU+vkSqQ3zN/vdQr9cQ6Rrdjg9gtLnfr3DbAOICVW3kRUYUQJkqPBlkLwgzP5
HB7HH2IKDC5YY7mX65nscdK42ZBa9CsmGvfrCiCLXEJ8k+hCaSQFCDEO8xu6M5OF
yMfHU9nSrLaLUErJBdGYiKI0d14wZaA+s3KiUJcFTXVk5ZBCGxVlvC/KHjduh1Yh
VUrBDUgOSMkg6MjYeER0C0cSiYGGoCganOxetsXN4S6hDN+YChrvGJa7tWBxDpim
+6vaU8Ukq+7ntGxSEcJ5iGXEq3d6WcMbHuv84AnEzLerjWxWejsMvxAL2q0rUOeX
nmRnoQ2WzY5/5UG47DxnWKviD5y9WHzLIxbfk+A+vzZ8F3B8+sp3K+Z7ZUxaIKMz
ubB4r64Lwc2bW4Q4hivTqNObPWRYk8EbhKbSgil+0Ng+hkXzeE3cQZYoDGcegux3
Yz5jXmLwUEuoOdzeLDuaOv5/mLU99/VEFE/Mo4c1M9/QCkVDduZZMFWsRVVbS8YJ
bQz1H+lPbk6ep7cKHRw1c4i/lROAxPOTL8UvgBDaTK4VxbF05RzjUS4ba9iBH3RQ
AFYGWWaSBjuZoZeOjRDh/I0zQNeYhVU+G7/PwgMBuHsMCms+diVjplgrGa8RC7Et
b85u1TVXSie0yEyTcibzZOq8xatMWBArGaycCgRigqnIVEps7bNW5eTz+J2Wt6ap
ZFndgBkK/7J31dv5M96MPlFHvslzAgalI/9ywYZicDlAdxsvAyNJotVVmU1JTgvv
sOqioD+THXco84GtI0vPdbdniYR+JA+BM22PLR2qqPTTvuorPF9C5pbqQDA0ON7Y
vGb8jG453cPk3ArFO9MVLqkrM3oX5/WqLTig0y7i0lzgfBUkSw5Bz9VsBJaD+yAt
UL7Kl/pjiq7SIK3d6ej1iGaUbH8ic8kioNKykdx/F3QUv1qK4wzdUXiou774ppvr
Vus9yGFJELOSfwP0a5qCLaMo+eXwU7EUiRJuBCMflHHISIOazh6nHGJufqqyun4s
OTpR7rEz8NMXKRpaNsygrUPx/rCP8Z4auYxTAOSUNdYJvo0c8dqG/NAoAGF+dxHR
FiDQ9FYDYZVySZeqvlB2GqCum+mbhqui8qfOTocqt0aEPhgIT05jsRK/OsWDyUZq
3pa3XUQP5R6B/Z4fuLAn3WJlguvKJ/aQ1DSDELE9nw5/hTSQEpr85/K1T1OvPXh/
K42p3JOVNPABH8bcy5y2X0FMDLLuVcIpzIaWK14Uq7HVDuA1REPvVLkDOJqcL910
U2W+1sm9jFgmRGN9dkelrkdhWD4YDAQUG5H/WKTfaRPU2mCLZLZ0BDz2pUROGBf6
Dvr7p3gCp0P3HDt0l9UmZuMG8RKBmr7n/xyYW3KwLGI/ugG2iCwfCKO2ez+dWtH8
r2XodSOl52C9RrniOjpzKAiwcpu0TYuLvxU3GXBXVC5B9xdP/RgpwK4ulqIcdLeC
dbBtFl/57yHKuFyQdCHimSBvQvQUNh5BIqcg53E9cRDeSpgF1X8yLLFLLf6g65iv
3VKDn2TrHm/7JNKJs3iUojU910HdzTAjNLxGAmAdF+Z+Sf0B9fxnpPLwWoyGfFJL
8wAIUwx8dQr198Hh8YeFGxRmxGEdoxzc58FwLR425GKrnUklYiBERV6eM3Col0cg
lREShA4ZzfA2znQPloUoMHGNARr7w6OM1mJiCXS0Ei/k2KjeJhSK1yRjU+8gvRMd
X6EQ2m4LcpJH9xCWf+yzlHG3xtpv63c/78iD5tCwGOFlqfR8jwNhdVVQaKM2QNw8
SE0QvLmUy64XQGeTT6wBCpqsMbY57q0KqvvZWaLqG0NuQpU+S8hEIOSnAKaiJ9HP
3TBOQ3aQD7bsZqechvEvhcZVRz0QqQcW2LSDnYGdYH7lJpHJO2GATzkplJdJYi7W
3YFnsk4gyBseqHIgX0MJ8gZrm3y+rZFdKEL4UtaV1jZhjYfjlx8pcDKTnMuXVA/0
40sK6u/3Ck/aL1Y0t2U+LQNK0j8d8s/JGNsg/LAJtfvHpdowL8jvs1GWVTKYEqho
L8jTHPT8RQNyrop5NDM1MTEm7q7/bWlortoU7P6NqmDP/ZwWOCUaD7v739XhabTE
nD2TgQYeueqi0Uv/HVhX1AEcDWyxTW+p3aeZQVSucmivj11yFLFXA2xOMq94IC7j
IePpQzopBWKqysg8YbdUovC9MTILWJ3R93tKfHESEOn/EXbv8U0zy0FmwV/qWws0
WF0R+Bu7t9zpRwG6N3bY7UcEbVyQXkeG4wwqxZmSEIDP/4oqZpbuRRmrvRNK0Avg
/faCLtfH6kCbVX6HIQL/W/CDmXfdaRkNNRcUrsFezgbGk6KREel0AMjZknII0/Yr
WEnhEC1hhQyhWbZbRDZoOhXXoWdkJ19Qv2wkKjm5Dy1L93NMFR5oKJIfEhsEkDQJ
PMs+a4clvS9rw1RWHquQZpgsECwRMwvVHK6Ncsqcl3+QDF/NxFaWwfzk6rWRHp1n
LLqSA/rsJW/hvppjzOr+AQqTJ1sXCbObXoUC95i2ojtC0gN4qnGNV6MAklFIkgOF
qh9GIpuGzAq4j6COgnG1MXCb35t8S7NTkhJZ/5KeQgqsKHqlsipst3NiYh4juc5J
pxlb531pmTsO9U+GtrtPpfK8DLiO2yF+t8/ZMtYFm8QBS1dLdW7NCqzg/Ldp+1el
607Gs/iSZ1RKWiAKcd4AYQHP0xQw6s2KdZHma/4XMueXl+lwbCehozmU/RKGrnMw
09kLhQ4F7Uni2o59Npx9Y9X/8rR88FUAY8WsaJ84kPYJJCDC2T84DPgjFYXtMdJV
64hRTOPv7UBiKQ2MdtFPONVKHk/6slJ2egkPlsBTMT+TnaJmWj6r7cpaB+TWBU32
vV3WJ2+C2wAwi0rPaglVh7P55IEX9TTONU1DbqxvfxjEE5yPBNaENqTlZQiXpv1v
RmEgfNzqQtFB4gTpM8+A8B4ECkVo9BLClNR9i+lEcG7XhlCjFcF3WNlJv6H0Lu5x
xRLML45nCyQAQm+huOLhKYbRHIE/UGI9AhKSc6kv8yNKexSiZYfrTGkObRkwiYBQ
twZSyhQ1WMmTHxQ1UYMJTV++YXz+nHd9n7KrfHjMxuX1pO5N0F53Ygd9Jb3sqWUl
nrPcQg8393ACr1ozePdn+dUPBtpvf4Uqd6X72TH2Qi1G+ppq3HjQGt2wmhoJ3tyy
9wAOU5H20u11OxbErlDw3jn8+JfIcvmR307NTrijQbEo74EbIm23K9UhkbTHQWgO
X5CNHQKmomy50ngTepGmZQA+y4OMcN9lLE/oN0jQSp/yj7tGz6lxRfjMFxv7ddB6
KwCHmrs7n5MXYMt9IXhv6imwEFeCTAuFwX11vRMkpUeEs5q0MrgZufYrcVpT9V0z
iex3j3mQPf1J39OR1GM0nfcfKzrF70pO82cpTw3s/DXgwqb/SlgLuv9MwquOSJaM
SPI60YsvlnfXhYUqWV4U+7TF0M+q7tJbSkHKRPmIro895UDcICjqW/3NVFqeqRp3
U59qQOh+U9FvGzbsOTpJ+mB8hLqNJPz7qG0pmG6560ntXWw5lWRvmonByoml3y53
URZ7VMsJd21lqiRCS/IYqV8cHsWRhb1dK308RaH6b9Tp7IGhME1j/MTwt7vfuusv
qXwhoGvkIlK7OIJFEzlpQF3rAM7PW35z4qkKeL7vAnlUQZrUP41nrNc46wX4tAUV
3yKJvVEfRn0HChfYzf1+2AOzIjI6LifdPG0iX6Tk7Vz9aLaTie6V9cg8btRG7exs
Yfwy31prSH8r/Tc/t1srhIbjwdt/PfxptqAGJDBadPINe8y6ikeyKtEYQryX7e8/
1gWlpywKTFkP6yQfFus448cagzxd09QdAXGm4hpIfIqIEcFiiTgqX3GubzalTwj9
2pq0Bz7r9WMPPjM9Ac5h7rlng0hE1qWE2FYlj4XvLvBUFIuSJx+DAFfkQpNIa0/m
hfvqT9MhqZAT6oiWEFgtEsL3ibHMWd+uOyWte3makKiSLSiNztvcnZJZ19+3jWN7
XcM/NnTB4kv3vzSIV44bEEk7Tutwjm5RQUkVBWsifB1c9mhvFjo7lQTEmBbaOr2F
DD69nAq1g8KXGv1xXgiUI8+rZssZxjKYP+r05sPiYtcHUoXhsW5dsOxKmXN6oAjO
/+Z9VaVDTLKB7EPXIvdOnbvpCFVOqN97g5D3JbdyituZrA3ZgF2cyUZIkvYtrEoQ
FxZWDFJb+6ET93oQAhsUTGF00zOc5bfF7p4jdAnZwLoAw0WjF92oJa9MHu/HtF9G
Vxl2xtABx/Veq+rvn/qcG0RgiHSP0cN4zCSfHW8E3up1AprAlzmxZTD3SDbShjb2
Gs5zBFT3rpTWnAYnYxDnaguvwxu6uS9bep0ySkAOLi89H4lJ69Vs5keax0n1IKnJ
ggMFspppc0CFh9FAtlHgi/iQAGtvmO0iB2ZB/ApQs1nYmTxy4WkLunjNNdajAO+b
0GYX9HBCWLoGK7iA3e9zBFErB6HVvxW8n4ICF5UsuVBam3jyIn1hRd5Md+Agfn0S
x+KGmJ+4Qr51ZqtIbMn32cdcso3XK1SAiUBGRUmzEO9qvx06wmC3miqupAoJgqG4
4n1z5wmnmBufBQ+F2rKvPqME+uBAu/g01IHxC2qgdfRcjRQt1YYVYpmF4b1xmINc
6JOf7dxRxfSUdflSnpT1d1bY8ugaWGNptJ2L19crNO718+6V8dFlT1aXkFWj8jEr
27GoZMQB7fQI1S/sXH2w8JHCxuwmdpBmlRYMjvnNcXCEshBOSTFdYFuOARCEU9Ll
AEVELSrXvzIefne5VfWU7aqi2+XCBtcSqPjnnyDO1OIVcOaK9h01sQgubwxoytBL
AUcZzPJDVvOlGukBTb5oIwvf1e590DT7XjZJO88KNrHgWGAn1UyPgGLmVcr2g+Xc
fllPTrvoREyJ+epxJaYf1R1tJFg17rVdm47x4YGNk9zrcKfzj7SK70l3akrbiD6/
WTeSQBeJgRkPywlYzs1EKgWIvtp/l9AD0DAY9pRID40SSFZokEa+4tBPYaJ4+GWS
CeZFkz0KNqePRXLzxDWe5n1HeCH/mclNdjCUVz+5BeerV02qWwdysNPdeUd1rUZJ
T9BJlssBeee92Xin29CVG4psyuwxFNcpRBfHPHDgUVpt3J7W+UVMrbx62IygA30E
jtIMRpODec7ZtTw65Wbd+5rXIcI8aWYzsR43sSXPlO72DCgzmqhiLlw2GK13e1Wr
KEqPiSBeS263d/9AzFaIcffVKiDlDqiUbiNLSk0Sxcaq+dfUahzhq29KwswLpiKh
YrZtmYc31XN9KmQXlhi+t1aI9FYLolmiVSohwIBbE3TCZFe48Xbv9Pj0hhS0yxR0
21a6zNh/jk1j4m6MeCylpw1QGHd6QjWRzq8dowWQInBdWeu+or0a2/6IKLl6xaaN
mREoyRwuf0er6tVYNASahtjzt99RrvbyWZ79agc3XI42Z5AY2z9jzKSh0fHa+6Kv
mqXkbmcKg+fm6FMQ7Bx36ar8l/2CXhMWWn5X/JuWSFu6qi9gY8r+LFqssY5O82St
WejCpbgG0bvRWWUGbRX57sXXphe/mWXiUicYoiMpfbYxqhJQBXjfK0XoP0MBQ7BI
HVd9r1+wYpX6ttDpedqcH0+Vm1UElQyxFCKH4NSNPAjg74tShlbzKbFli0DehwQJ
UuDnnVX+fv7JNl4oT0/kmlpGP6wb5897ukhOTh9QFGCFJmRSRxQAtpotqTk0Hz9W
Zv3mrnC0cw0Nf/TWRdhEnyKkNb/jJ8fK0+lyQWSjJJ7uA0VROAmdJobCDXrL+v35
zRsL47DYsXCOvsMtdbJwG1OQrOcgWnUV93+fN/uatWv0FOGU45wo4BLM/Zvn2sqd
rJEvZeLxrwc3o6f3xmDXS1g8VGcXzwQl3bFdgk44hWE/0JRQ6KC9zXE+ZylgxzXm
5tTR0lk1ln2MJKWdHTZcD+nwTrISE+5UK42GbS40Ur0CU0vAhliIRjyMVWhwiK5G
RP/meV0O8ua+9TBeZTytwgyXmrQkI/ZDWXrWn/dxc+s9buLaMsu/QBfpFZB9Qn0c
OwI9/Dp2Z9Tr/iWhmSKGUyoWgmrNDulH5WaMoTUbJpH9RR7LjdNvlkxh+8dnmnp8
VCWL6lalrkh6fd3Uk0Hq4JgvuKQcwb2HkSORp47IS3KeMhhL+4v2JhOUuEZykhvG
6mtEOyskOvHgbTr5BVuBVda7ZIAP50Z8wo/C/DQ10GViReYFU0iPkm46VdqySqGn
tXxWdbYaFoIn/zyHmib7DJEb1F2YglduOlAFaa89y3FZEdYJIu6MjpAkIMfAGSE9
GMrjEKDIn9Lr+qDTkrcyF3P/tLnqn8Vr75QEp/ermVI90wFGvYVejOr96GBdoAv9
Zc7sEipuCp7I+RdDZfcaJv/GPbs8sldib44M880KtjmWUcxkoMvRnGcdPO1oTmkh
scu0JNQQQQsvqf6iTvGSBqf71bvpzAv5QSDC8vfyN9RoZo0GFEcGckXzNHIMJ8R8
2uL1kFZM72DxxRfFuxu34BSzHxWAZKFcmOCK8mu4yk8JUimfOLNicx/9oFCfrCE/
lPqZBZGOPmTedIUFMMf6EmVprGKFd/8OpoS22nyRJChENV0hpqphVIlKR/3ODdf7
6+0tPwCvTp0cxMSrQxoxJOd9C7Sj9IaTeoV+z8NGG8xb+TnCsN/IAg86C6zE/lk8
CzclaRk/kEwjijueWjuuOEtL8QVldcpjUMGIgOyNBBq7gTyFKZy17mzenvpRsmmi
z4tHdo9wH2QAH4q0cm+jjx1qmwtcSDmZtLwrdgD2TuGr46FrBSPB2VKn7gyH+BHh
O7k3TE7WkH++aJeJ26wfeHq1MRwNSCEXwXGGVANQtpNoFrTeaOXOLzaMIPJYxoOX
PEix9/s/aZWnHJkBFlF8h7TFAVyaCxyPhty6oyRYGegzQN9f/3miZ87UbIbtgYpr
AYoX63t3dJvG71oRZf5/ofpiEHdbRqzJQl2sud2e93DXgQGecZdNs7VAEkAfdJ3j
rqMMN5Od/dJv8AROo9RpHtThIU4njrPUKL30Bxv7jgXICFzZYXv9rvD7SM3NaSBx
F6ExyjSVszWHQJKiJssIz1jPUah5LBjeOCV7qylf0cZNLQ+DroZP8TZwdZX2VM4N
wmqDc9Dr6AAEi9lVkmwPhpdSBYET+2GJVvJXARk6nnWykCF5ejuGgtzrbid7f1K0
VDf3b+zHdFgGkocevKKgjYCTVZDW5JJrz8ZzDgelkOqsFluhz+8BTyUGUsLE+5FX
CAJigH+GeCQVMWN7stO5sXGLQ2Qzi7hFWCT8tR0VlMw2JRnh9YFuLhU13n6SE06k
lUN2NOOFSaZxQqw4RkytXURkcPxIfJPsKnmK2d2/i/aanfoqedSumMu2eLfJuhgB
ENi4c+nqGvVHYt6W5FoiTCpGxNjV+XfKKHiqhKVkxnyyrBICbrscQ7cbEDxW/SXE
7/MzwHQpBfXZ2/AyEGnuv9Eq0x9j6QI3YaNurO2B9e/N5kCFqqkY2xXinqaQyda9
cefep2PYrLRvkWeN/LuSlQBF9OiFqavQOPMq8PvYbOLS7Xi8zfXdU10Smb5uf3Pp
wWzYYmUBPK7CVfruPTEvo1KvZLQRPKHHYoKsLhIQaYGuGTrzs3w9TRyVUZlkUFhW
+AUIu3mpP0V+tZCYUn/HJlqCX6g2pW8lT5hyQzU3MlTPp2FBbH/QNWzs1J16X+89
DvcntmSNooyumXElzFEMHiaCggiiY/0vcsW4+QcUGrmTI/U6HxjhQ8j/zubmhzsl
wQ+oBmyZ4ZkKo8oc+sCBKMWQ/eeSDLw5MXpFiKaNgf/A9yNQ0jCvvmPo+ywFh+Fl
CzoNbMJzGvhpzPGOCG4mH5ppi0Tu4GfuaBxq7DV99oGz+wwr4pBv0nIC4/6N9e/w
7AgXxj0oQDBRRRLlq/V1pyqwkoHYPJxeWwrnRVihskhjb4d9i6HxJRCjDu5TVDgv
D4/xUqEGT4BQqlJk9pVCzT1t9lvcgDZJ5GSiUuyfhTieCdQ4IYQpcOgxTVciLWUp
PsrpaKuiv9r4hZsmGD7JGMwm4w/Ukjr77BZcRhXld0TvDy/CktHWmjoLiCcBkbld
wdRNN4zAgaFxBDYr9Od9x0O8DjwtGpmN/LcPQaJosgRoCZkKGrzhdXzpne9C5iLj
tRzu5QaZTmGCbxMFSjydMvMJ9yCYf6kgjcBjUh5QWxgfqqrfuPOw8yJ0u/1S7KoA
SovVZvco6TjKPOl92kj7c6/2YVCogb6ThNO4/Ykg3lu/nZCczJV+W7KoMIyXEFfr
p6ndzsVdik2hPJ59s7lFbmv03vQZAEaGiM2OUglJdJTzpPkbtQQSgqllYHN3kttf
i951AN5CH5OVF6iqOY4hkLUgTHPMfrgR1VJYNvZw9akO2R8rGeazyNIS2jhbo6Ir
YqIUs9Orhrjx9SM7DrJ6+M/6TLtlRKqFL475caw84On18dMIggdhmuathyYjwiV1
a+tEHF5vWU+/zyh6LWdici0ioKwpJgg9rFBYHjngpPsHiZFao6UqIkJg3YUJa7da
oxUwIjZ3xljeeYWpVDUwnSDOVq0XZ1aHR2ZhA/WnaW7KTI0o/b5TsjmrjTO1sa2B
eVkH64q4MYJ3zDQtkf5DFg85qnlPFkwcQLPpcMnNCrqMlKr1lAnzr3cthSB1zlX+
bcjhBcjzXbLbSSk5I90BWbbfbBrzue8ZmJp1UypmQF3rq1/SLbKz5Dyi6HX4iB0G
A4altw7HOVDgCCLclQHwtLeVD4ZAyE0Tl6xOug+dBrd5WE97fiXG6qXqwWSkoJil
4WFrY0w4jq0Jw3ysffxadI2lOA0HJi2jGrahjbMSvrfKSHBHQ2YP7Dg1kwucrtV6
MYWKD5CqyxQhEucnzGXiqRQ5VfNEl58hNSRYZUARpPVwMjiTDDn7mTQ9Pe7Dilm8
AwMX79kn0nnUy9ppeSwMQJ2TI1LZuFGv9zStpxI7D5yAzSUM29fOMBEmBh2j8jO2
Xh8HGz2NUAabPlW7dlRHRDOhRYpz3st1lX4Uq4uu6VqF6rDVJ2jblt74izOVm19+
W8XMgUHQPLts/8FfHHuz28OnHzmBEY3m2gReQhy+PhqqK4I5p89VsJr25aBuuXBz
wmfUdSVnIzXpfX+mfN9FqHeCpUE6A/bTdGaBw0fhQYtXeklbtZRZh41dPp9Mga3K
HzJEr8CWiUiXcFIOF6CRtus3RxEqzuwS5txj21InA8qL9dNIC8l5jbjMba/5Ejqm
6jKq+bru9SRYmIiCK9fvmDW0CKH3i4QzH+X3efwUQ6J1OFMiIiUIGW1Tj1Qe3jwF
DY4XqCNT/O7v0jbk915CIWxDgsC6uYeOY/EFVd73Wdz3fn70iK7DtmT1/xY6RsGI
Sjbfa3GL5nNVche60HoRNqVXKTAlWCayar45taVrOIrDGHyGNuqZIRd7RBSMgE6m
19Qb/I3FJEwqAGIcqj79PCvdMEq/QP80CtDgHe0SWQ4AX1B3rl62vrLpB5zCgzeL
cH4UmfT41Z5Lf1WQ+1+mikj9UksZ73cVzeShhgGbl1iP+Ca5szlxFi3qTVklMFSL
zmxCyNkDbvFKh7fm48WNReOPzIGfg6rhB6hh1+UYvtxzG5m2Tv768S38iVUQYvZj
z1F1Mz7SvYjrjMYpyqHUXf5k7qAyfVsUTfQqtcX8PnRo7L+Cyj9Xszx8cpGlc1p8
xxJYZgbAjb2k0zJSCkJM8dskzsD9RM28zG7H3pXRd2pFhd5CDKkpKp6WF1sAkvZ/
kkFD+ISmz/b0DU+mSnssQX9d4gsiMOqpyBrFtJnynLipejMGgIcRwd1m1JhU+uDI
XM9/YLJXK7RkeZ5YLzwvaYGtUXYqhy8xtMPdWPRmU6flZHE/Lmge+tLBXFDseCBy
YJeMyHWCBPUobvHQdk9RwXX8zJyVsVCCTgx7GM1bwbBlNSqUFeoVIkbeOGIWVj+s
+FBtEMUXUPDb0QiJD4TgfcS86/6eaxvCDmJvpoHCarkB3XJKwCe4Jczb751ALd1a
bAlZhbzwex8E+MjFwaF/K4MuejifyBVYz0phknVRisM9tlVdBRR1g+FPc4858CoR
+n8GWpcsuZ3BMSHL3yMU44JJJxrmmw2v52Kzvc7wVnaV8L8oX5CJi8Hf9m98MpEk
8aUPem/zLjiw7VPLN8oYz0lrshxcBL0Fq0I5BG723/2dmZ6TjhgLRrNMQhxOO4oN
JtuFICy1GqaZKZ1zH5AKVKcOowiEe4SgQ1Z4I+47iTHIT8IKbR6JU8Xgqm5U9u5I
z/qty+GOqUw1NxdKUaJgbViNIW5Ld5SRltG7IqS+89DZs6tjYQm6xbKvMerThHEN
X+p3aqliz3hFRa/76O/rBudGeSB3k3GgNXVDynmT6My3sQkqA02rw27Xf54zlO40
wLlr/oyUTetcLJIvSUi2IghKQgH8oorcpEO8YJtRmKzCaJkGB8O5g5LbN2XO48tx
rDop+3p+yAtVmzBbOEwSqYsOZi6cZTOIT4dB969P8o5P9dRIv6KpZkgho80TbSvk
kxMon/c4SVQZv1c70VZTIWaMaJnOyYYdXanXXxW8U2kqyTcTSfzh0TbWZApPTrlO
qKcuAW3iDzyTL7coSbTdrvYSIW7mphwJLfmv8VbG6q08SHhGhFDhAjyI7GZ3jPWf
/qybyvpY+oIlBjc4V76ksGhgwDE6fwe2e48FCyevjZ66VqliCx1sSObJq5cr8cm3
/x8fpJYn6yPGmMt/PuKiB3JFSFmXUfErtcxyHuyDT9cAEMmpC/AX3das246OoCvH
ZFxaxBxmSdexHJR8uliP3a+zNDNYREyY7zl/gNiph4GFmZRa9n1r1u32wWfPSfTp
5aSkOCs5QcQ3lJGzmg5ADZZWk4NAtFI8BMw0o0NLM/Qm0t161RgEMDGL75UBu4Fd
tVKIxFp15AsP5I23iVO3KQxHnodYpE9PLhyeZw/MCopII24ibIi5B7tlJyePA7Fg
/lx1fMD396aAFUo3jEiFjCQdwR/mieLYSDxT90VuO1NxNaKr6h4a3rlq39F431vz
Sq1keUgmtMDtV6fr+K7U96H5fBohjTu/h8Q9pGyO5I81/FGoMVP7MbKLcgGLdYTr
pGIM7oqmw35pCCBUZ7hXEp8PYDpVisDzYTkZlpxyrtPV+SaPIYClcWZYo7OT1FAK
VvMONjLSNGX5ZNDQ6eRo0C7g/603eyByO/nKLZjHhCLNl+wuStc5YZefYzPHPj1k
HoPPSEQ6LvsmmootBr50RJvi3nuEX/ZvVUt3nj3Z3+OkemjYGHBL6uNC36QGm93R
k+/chf73LiGiRREeVsRdaJxGQ71nCGqFnO8BuQqQb2+ScAIur9b76jEOn71VEAT3
BFeKQLgKCMwmZyjVFl2MgrfUmr2d3qWnCRbatloq5FJ5YxYiB4ADoXijP9vUsApT
tpQazqA14QrvBRw4Knr/IyGk4hTv0bqgdBo2S8I6f1PHPFILZGbRmr3fODVXdrUQ
g12p47pDlKnAW550uoyA+nHRoEzBxosZU0+VSoZyFRbA2qSfNoXe+eqN0b6Z6+tQ
2CQ3NgY6fZDKqUOFIIwWVjd4sbzzfUj9RaAByzP1KdTceUAf94NN+HyLbV/9/4yB
/52qXJPSMeZFYSyU/BiQjLVYzhJsih5TgKlUka+0YfDo2EjDnFttVwZoklGRXVJB
cmArRCzmfCT2oY1UyPi4hKzQOoV+jBQ8pyeBmB560CoruO/MBNxudAjp1XpqSD3S
ggdXQ/f48zxB99EeUPFbWSBNVHY5ePucXW8/AsXZX/8bJTm6ZSSdga7irUa2s9/+
eUaY57hsBR98ePp0G1uwj1nlBveUWdCFSIEY94FRHO/NxIicOKXEfjLf+nVr0+Wt
73en9Wy23OPlXKQy1wSW337LJT113+F+KH7QE1sLnn/YXwM+eyoYM7xivIBdawz7
ChbD5AWrrpGfYkRFcUZwe8SBoKhmToQsA7KDrnb3PVoKA0uHCgbpQcgc2r4PUYgW
wVgm0/o+U6ZR7KdAKJ5VDDc0qiUI1FPC0CK1/pj78KoOR8pzz/NUCOv0oz3sjK/e
nDocw55Cm0JH0R4dDXgtMVGPVELrZaHh0hBWu3T0kPyFBur2IwNXL5HHxXy2u0Um
0h9G4Rnn7AIzHdlq0qo86VJeBBh4SyqB1FMW7jMVSIabhvaf0mrKLy5vJbhBI7t1
jjNFi/kuHiY9ui4Cnes2ZoLo4e+N4nE/rQMScSzAdhpP7lUni0fAUpPK909AXFlg
Riq5llwBm9qQPdAiF8IytkpDQn8L/TOJNF83gKbIl07cUSZBXkO6BC7w7yqw+j5Q
L3sTF4Uzs/wU/Kn5fAbNbBXoM6kscXUVUXRzYhN7aYmwfprf7D3tJ0mK8Hi3XEuJ
ed6gjrCpGiF14XKjPSoLiGC82ZJ8rK8aBD58potxKk2t9dhAqzLiN3kLOLVLA7os
VGOUQIUjugjz/pc9KTWKmJOkUUW/5Zr7bYSlLLzFEjsU5LeAR/SL7QO67PDZJLmF
ZbLCtWbVluhY2/2JpPiXbHzZ3PxeKSh4F0a5fqpn+ApFDx5rWY9J9oLczeFCm25m
xS5vICfzARlaUZ2jmCcrd12ugDuaAzeJgzOhUUc33Q7NU2MNS9MXIRcw+DUJBvqm
uQAIxCBfAsDBiFd5Xrt8aVJSXXjLm4hni3+We/LxAZTBjU8Za+OsEScgfyk961Dz
UjBsJvRQU8NLzOlkohLFnyhBdCx5HD5ToSDDBapr5exJSSMCj8ow0s/12DVps9sd
fP/tUEztLslMjd9DdcKamqWFtnE3RWpusULkLINef2qjRAcprCRoSMoo+X1B68Qo
Jvu6DapPNpGqfNNXf2201MLj6d41s64v51hsS7zZseEME20sA/VYaSoFXUOEM1e0
gzlpnlOgGGJtewKtAHxyFS2syvJ6TWFX5UQU1kY6q/wejucNpo2uSjMu68xvdYkO
C6zPNoRvGmae7NJ4vb6IJWqdX/k3rft/5jpl0HGvJLJXmsMvQtYnnZFzGf3LGlb/
h3Kv+YVTD9NpjnUi4qWS7lEIGqReUKlPM5x+mnNOWhGm3Ht5omMlxERg/Z7L4BWd
dxx/iyc/kKnJjgoOXlNk+I03/gOf+BlKj82UT+0uFQgRESPTM2WmF014/kBJ5fdU
lYRqJ8NQUwivZdQrWaUS4LOypKWBeM2+jIFt/8VjsQG//iqW2YL7BHzmfMzxQiWX
maT7XBLiNTAidWTCyeahr2gEcJzf2MscQOkeTXj0gKdyD6qAOnkfhj5C8Eu1qf8p
u6Iud0G4763snuY9DVnekX61sa+eKR5TDRjqHIQQSWuLSJTmhynLiHpQBpxsrJZd
7OsF9wAJk95k814z+l65gmn+cgR/joG3v1XWLwtn/pe+e52ZAdMzElktFHBkM9Wc
i3xmUgYtdjlXukhscp24FM3CHAgbw5CntdLqDZ1mzjU3/Iy1g1vHxxHmL+dyWmOG
FMCTBtiRvDvVmQE7NfYWCR8L+Qhfk8mMwyDH3Jxsw9lt081Es5WLtTS79VJkKx1L
0WBlj/lXeSvW55nJDCQjf11clw5DYoo7n253ACaUMj/zBR0nc4Jutu7yXuwy2XjX
pn5exmzMQt+ZRKOTfwM228pJB+B6HDM5FcL+GG5Z89BJ+lehetOjBBaBoSWUxQQ9
MwWmidUt6rqMa3tfmbflQA9Bn/W8oGxPfwE8/iFGxvrwGR4uXpttYaN7+rg/zq7Q
w99xSbsGt4q4YdTg6WIf+SYFeMOIzsBQDQ9P7+DfaaeHN4DJN1ptZ9bcPqI1zVKt
xXFoJ0j+50jKRJyb18fWhNySbmOrf0sIiMe6roa6aruHvm4UvgghMS5MBHyK55Dk
Px/1f7Vq7x1T4F14x+yT2wfCCw5L/hyU00U/vEe4kSttk8N8CDqLxvjCUVjFsnt+
o6dAUl7vBEq+qT0nuEweVoYYejtuvj47Wi+1WApvWRxekcpC/8BYjE4kbxi26qMi
nvnoEAqciJtVRPA8TnrU+sXni8bpvGBZ1OeiygPmi2esSRKDqxnPbkd+sslBoEV8
n7Cr+HqxwmT8N2gSSAL7XAGLofKC7/BO+827NY0RHZAV8xj5l5oihDG0B7NKxecL
rUSHfOjYSvAYTh7b/HijfRjx2lqm+ALc8M8e5SZ0pclQC5QB/yUpfbVSWZRymNmf
zeRg3rQUxiJRzuolg+vZx/gniR0ycPrThYlhZtt4ZU90qvFRwSho1bIfwhbtuMIZ
Nbpe4i5sNHwEGtdUIpohZKOKAZ2LorDIWkAklKqrIyzZBkArDm84+jfNn/qy0wUZ
G1r+K9+CBK97O8uAMeBZgC+mI/GIVhxNn0jRf6loYI2pNXl+8Zo7UQlNOQcDWwez
qd5ys2UXAZei8YsDZ1Gvj4O/bzoxHnBLYOgCNAIzC3lUc194q8oTgDTB5Ij0OntI
vuINxiIuC2ARf86DGAUspDgQV9SA1kZE1uAd5DwA2aXO9VswDZ9pHqg78F473T3o
4U5ymg1f3HrZkkZPIOnmt9TeBc3cnCqH1j5rmi4yrnoDKhgLlBGHHtfrI8k0fHU+
tHWJeBdt4AV56A/5OjAokAe7jAqAHhSBw9W5GdFB8f+KswugA6Bl9tY5glT9NuBb
Eo9EhJWVyO8x2mDvnfSoToeXncH9C7sC3gOYbnKKyrmjMK69TKw0dpKdjyC6mOTe
s+zvZ9TmcTnmdUPkn141gBpXfNyyse9f3YAuNM1ixdM9YX7AggmwyRhchwJbomOC
q+lH8L/pphCq+qHcPTWnXbj8uL2hqRSeX+78PnPQjSp8qUxli7/cPoJdWrFCsnqo
ZLB4sLrQ4QMy74UDfrRaC8DCZDK34Nt/6QuvfHBkQgBT3cz/AQmw4IKmlSKgzrIW
rl0ZJ+LScUs0bz7+P80i3kVOkx9R1/UC9yoTa8S3coYo8iyVfV/kkHxvrnt3rKxI
YcAk+Cr2LAsGVTbHTeJ4JM9xZmDGAoMk9tunG/x3KGzLVbocWKKehTHbC9re5/lo
E2hfAVkMgJ+Vq8aeQkfcQgfKOkQeiCj2eRKM+FBVJzEh5pfpL/qiZMYaW2apv+cS
4VHC3CzIEj6QEqdaHauy2VXTX23A+MQ4BxtETS+vsKJG81oJbia/h03hpv5nur1g
R56HwHTCjuD05DOFQlA56bgQbafNim0l8n25fvUDS5fMzx8Jvy82fdAZ7pVE5r/n
Nq4fp3ix4AynF5uz+R4sxCzkGTddOTOFMQDatK5eeLhQJXiPWDzJj7rs4is3c14d
MeNrjzKKfFqt/hQzLHa++jlNGz63exU3Zdyr/J5/iXSq+kQ00f3l0L9E3fnNALNr
wP6rWMx1ztJotEqdmx/RNWuzAktiA/lfyRwKEKt/Y9UxkDsadg9/iQZNvQlCOElf
3yfPf8bx2nAGr8sWNWeM+DYQVSFd0f5MO/1Q9Zvz5WqlI4VSfwO4kZaDqaP/Otnk
x50tbVcXH0YtvgC+tHsuoXpFst9u91jQsjo5fQY9vlcDTODN/TVvlvNS1E8nwTaj
knsyz2UVhv+rkta9GpnXJsRfyvSw4rnj+5XAixFJyDnMYt0wFl6vAypL3UQU/LE9
a1T+DINR3NwWMrjkigbKZIFAT/BcdM8blsFU8w24OE19fpNgfzWnKP3l/W6gW6uR
ySZZLcu25wqBKOtabW6bZhipwBdXZNYJT2N/X4Db/uXtUPg7Dh43vJmG/DpYyNE0
L7kaTWivEIEm3pny/XsYq7ycwvNQ82YMWE31oylS6fdPqGcJhj7A14zdEvlLxect
z+VPmeH9Atw5pVYu+sVGg8FAJqC1Jpwgdd5mIY8eXMSoCxWXOlxvBMXacKIqt3jw
2DuItQffYI/tRfqp5Jq4KBE+qDsBl930SUT7VgH5lndZgPY+/H1SUU8RRrfPdujh
Sy4I5+8jlfyd1WcytXnVZNq9Abcd/NU1fWwHqjBLa2ekni7UCIocsYaaJlhVuA5x
xAKRcnWcHZpo2ieiELPHXMT56o7AeDp4vUlrCDVmQqnFNGcwdyvaNt3Kv+gc1KD1
tUh+a2Qx3Mu9tNJwlFAhQ7HcBAAe9THUiZnA8o67DB6kidLeYLcXAlkVuAOuMrGA
7Z3YNx7Nds7Idaz2xbcxzimPPmYGmczV/9QZDpkasqpWbahxwb3aBVfpVjae41y9
niSBCsuPeE/ruu0fcXdxpR1q7UIP6vO+BqTx/ijHM1x/w8Dod2BAsy6EgbrYVjxr
JCsChpKS8XgU9WN3PBgjR/ivUa8bFIzYb71VWucGJvZml+vaT2bf+ZlhXLVkAz+B
V8ozafrd8B/f2yUW8rCYnJ7pyqcvDFxPffvdrLn/5ZMzzJxgleDHGDY7VKA8QshT
nW+ygDNDBP0TlA523q0RL2LtmZ1TZnsBGdY2UBPlUgYj2fSpSDhMIw0fp5a0o0Hs
Vg33akuf1gqaUqC3DXM3g954rByKg0zR1kUawb1imOD9w7KYFOqVWBSK3n40hxRv
5E6Ay8c7ZlyFsV5AR4k9jegzktjDPaHK2Y25MzH5i56KPyWhJyhDtXsk9cddAwP6
7eCPws2SBhBhlhjjYD/Mg6tMXVy7WAFIew2y9QAI4EiuyeU+/u/KV481ea2DDN6r
NT8vUxq4ObpcylTwDvXCPt3Xpqza99hGskMOm07UlnThjKcj02o2x90b3x+qPOlO
GsykPai+p3V9deUKCdmnVyxrtvVgky3nSGd1tsYv34w5rXdX4pAaAKbXFrAZsSyp
qEoykk1wxLUngQuvCZ5C1cA3NBozMkO//XN2ZObcyoY3eY4MqZuMeaCLF0UZjeaZ
mpaZ8IgOk1VMpUIvtRUFRtYduyxUz+PE+EquXlBWl51Rk2vng2DLxgQ0WESM0ui8
UpsaZuxzMtO9e1Dw+Fl99kb2uac7eDWQnTv2V8FG6DJYhkg0tZhKmWRPecuG8QRr
+EybY+YEuHpaPhHsq4zOr3VMz6vmV4RykzWc9k1hZLP5VC1brrimEQHVlS9j3apl
Rvh7PQKYPPPCvL3hO8GzaHxqgQEYk2aSBGzQrIctxRKWzx7E8cZOub/y3ivFUejg
L4RDsxAQArgtem97APcbkLugvi0tgyTKYI4uczwbxigCA3qAElfiYJ9IpfgfMYjZ
Xs5coq56NWyn0yaNZgICQkE0bgKFsWPmh4YF9Oin5xujS312ZmB2R3kIbVOZ51gu
TT/SdcBahkuXyXgxbXWAOAq/6EWh76IXQ/j/SkAiuUkcNdGxkXMEgnD3ShutthIP
KK9hZPAvCAHL2jVDrgr71YVv+fegt55WSuEVNkiqVfEkgz+PCcLWPp42Ow6OoL8B
XhSJ4CbFt4vZpaXM5TT3coV2rJg0pF1AUqTyQUpbzLTpSmiz2rkHkVVz9Uy69WM1
/OGcrbZBh+tsOq6er8E4aEz+7A815zbeUGI6GveOej/dZQAeh3qevEi6QEzgUm4Y
2myWE7jX5P3EG7UPcEmWrZhWbwzGyDTode/uOSep2rqv2tmrW+WNVifvGBII4o8F
SdvICLp5022RkfPDjmUbPVMorxn2P0EW+fKDO7Ni0elH5FGPg9B8kT2fCQLl3G4g
s+JN3VL1U3LsCzXT/dUS6vcyb9yUM84X8Q3beOS00n+AD/pvC0cudP2TzSk+Pa40
Zq6K+jVhjo6FdkFfLV1UnWqrGp2hxdko+3PKwW9RfQmOEtoxX+bL1KYznwojhFGu
LeV1iwWEyqxUW1U5FZ17a8iQnxrIeOoGt/zhoWcJ0kAg9K99rk9FO1L6EGqbHZpc
M6I4wHDqYWfxwsWl6s10GfauluYBNNJJLigvGoi+OYCK2ewVj2baUlsC91AKjvJT
DcJvTp6XA6qRInW909JiHJ2QniuCb6p7ITWpY5KfRMq5dq4GieuLSw+8ePhGeLjO
dS7C2pQRSJwZ+3q+0rCjy7jw/EfxJ1dS/HZpuYdciLgadkOxbsOvK3uKZx1yw36j
KTsnol/FEcinj5BbYiLm2qybBq5YYXDrB1tnePSzh6rotoirbvnsvZqt6NBsJSfg
qwDnRl6rhUTo7iPS8x8Bt3vuKRu3bZXCFwmI431UIQIiB0N3WN6EeAw/dTaJ7NET
nrTbt7f+judlw4SwFtNN5G2RkUZ9FBFwTBlELy7Z9Lkn4o8GS5fztIxThdJZLJls
vOvRZnYqfYuZvauB9yyOVKDy0Ak+1aNep6Iho5WADLPOxYcAnxzW+Mvhj9QZRfPN
uiT549/6nmSshlxlPKpbjwUFPTXJW562JhPSWSs/BUNCJB+0XROnHc0cdZ39nN/L
4jPUre/ik7tHi4S6KNAsVBn0v8uIOA5OZTJbUQQkR0/b6Hqi5vyn8p0xq/j1MJc/
WxFXySFSRTydkYn+gRFSHDUXEXuWtGEF2Ww2d82ef7hwqThu8MCKvSlvJYKbBP8Q
YahYU9XIc66Obyxzq8koBCouxQMbHMeu7wskPEG8zTODYtILXYJ0J9izCS1kMvhf
nNXuT/X/jER9xr2RmcWeZg0ceSjZR/H6zsRkoVuFDvEkwZskAREWZvEOljwWfo13
LAKesP3nxl/4KElLXjWJrQ1gep+YYhZU3pGYrCWR5nua3d/BKjDVEd2DIj4Dcg2D
Zge3+0f7tG6BpB+0QSw6SwLzCRuf9BxOXqSEQK7iKGHFUPPEdys1ch060AVBJfOT
/si8D5ZJ9XINFf4+nK98JaZpcvMf+MveT8e28R9siWGRr31vSvwKaI/LmLJMjm+H
078Lz+xETlYT9Ip4RKFofQ/gPinnAnfdrTucV6yWG5JNEoSk49OXZttXwk+OjlQU
rQtOlVZfAfH7Us3b3j3PevUfc3wak0k3BgMW01hxMoj8VtG4HKry7PgmJ6bPM6s5
Tr1e0o9e2p6rubUjf83p2JOMshwqjIFfAcAf7//U4R+hSKqm/b4RXpqFgKEbjtdb
WilDmaDL6+eKC6BhurZUtzywliNOzD1jrxsFxamDggyfeSUi2plcVXSltgeG4MKR
Ws5URAquB9MBZJjPrJ5Mhh+VKO0/77fvrcWSfESbt851g0xuWnL2PYKy+ubhxlPG
3U5W+NwaaYsbzJ3lbKied5aJCEf5L0n+zHbzatcxoUVdUWx95bC+pk3wDR6dfkxd
81Sy+fmWwyAI6ZRrUt8AGr8F+FlFOvG/SWtnruDhs0oMnqImh0ECMl6coTQx+gfM
guG83y9uoUVvxp1nMtZ+Kg8n8KL6tgUo4Hxk5fTpsFTZje/n0M3IgFMhLWoXSJmB
g0syWXpcywloF8kLROFk/jBUAjTA5QTP8gy3G7eK8c9aDhEbAh16YGjrbVyDkjOO
l/C/AI+8RwdG91rOPxXGreK/gb4Qdm+QOGMPEFJfwJP3BE+k+3FBITvMlr/hu/PQ
Jj1Tn18WPgTELRg9WrhJL/3SJjQK5RMfZz8PKUL+PCM5kvfvzEqFgu6zudVQ7Kjw
WE+Tp5kJUeNoORJ5xzS38F5Hc2HNJoHfxTLNTLaDO07pABcil/PKAhnGMc0b/B1D
XPT+NR4BWurR8IUROuQaap3tIRomziyuVCBr0s7jd2wnDMyKkP4dTbHqHc1w9L8O
CZk5oNhRCOTfTGaNJjLWWE/dgzUjRBA9E5p4Sdf+2lNaCN0AC2C2I+u2evX9/Xyc
MwRxJAJP8hlx+7N1LOuJSkhxyfzqtzJrhgcf/HplKCnpzHM2PrWIFHZbUhnBYJGx
MTzlrUYNg55AkAWxiIeopRsEB5KhMGw9Nx8BuMyn722FY3O5yKnBeoQts8xOnyd0
VzQ00X2PaWcpbiAlbyJCZFTFXFwA1QO16y+k/XQ42a1HvOzo3eoWW7u/cvkdklmE
YDwRdCZHT0hd9DMmdpN7bmbc2/JjvhawNYGyoMUrb1tEH5nGepQShW+HpbSyfBMw
bgWQFMwUz58La0cDN2GXzmACbEF6S3dx2rgWdGk7mZOhNAUkKl6e0762D5BR+SEE
TMwEqLPorxrEnPMeY2ZocmLidA9cqQl+y+T7SbrQltLbZZIOZMR6L31FO+nSq2yy
sw9Rxx6iHSinJh40DL0AY0VJR8KnopnE9Zc2IjkxzK5DIW4y3KM/l9nDo5S4xT1j
s+oWm8nAEG7dTzWuet4QdkgD7X3Jq6ByRfDIZUEv3b5tmjMjbaSDBhFltbAcML56
f6z3C07wbzQev+Xxxf99lLtu82MFMY1qlcPUA+I6uq3/5O9kbblz2YvLEVez6J0g
dB0RUcMAQf4cJwE9SA1zd1HTf2lR0GjUZ9WOd07O/OFyym4Hp1zHtsWdOpAftE8g
rN7ZKYTngb4a/xc+LVw2uKgoD3Wh1y9EGs+E3Hsc5xbL9yrowxEUbJg+CG5Ckt1x
YX6FvKJRylWtMc2aKzBZaJcoE44PdV5Y9EWM9gDbDopCsem3OsaXqnlC1b7ZWWXg
kqOr01n0p8NLWafWPOwl1Z4DnOaY4X8qPhr4gnk5kr5UE/NtOZNkAQa+lYpLmxSd
3H0Pf4JjEm6uIqH3d0nWbMIn4ERnjFpv7YAx74Kz25CoVmDCbDC8GQKv4LNPbvUG
sbcu14ui+OxZT4PUjwLgE0CPm9xlm4seT3CGOkj+A2oVk39jbzQi3QzVjK2N4tRK
zTyAybUdyB4WCgsAQ0CZN+SaV+SOMAxNztuIiB+QiC8Ew4N3e/2+QY4ucwR4flWq
hKLr2NKiiT1PmmlMFH4ynymRSZ06RdzgxFXvD6XazB8aHzf54QOTyDfFenqYWvh5
Y2Jd/HxXD5B79ogw0ru8B5ovSdfnUXEl0blQGqdywRj2BQLfhs+MkJ/PWzUWLLT2
tCu8s7QC+VejbnyzwRH+eQTpwVjk67lgTcVMeE4b/goSty0SQ0SA5c8e+cPxdD7s
u2n/tpkljQNblZs/lysgVBqC1DUZtBzW9CDKBTyXlR7sU44PfuDX3pZrT0HaxQQs
Wg0CMvcGaEEqhawnivO2k9N+/J7xwHR9Mt2KbtjXQ23siT3/aLkghTE/okMgbFLd
Oc+swHlFPVv6To9fcudvESFMXN43It9nDzqb7lp7OdW5r190uYcmFA3pfO59+vHW
8cAZK2JP2CHAo65FMZ3vnVxZS71EnJbZfG9TtuN2eqesz58ao//ukwLM7tMA0YxO
koeY6sxtFelGp1cPBGROpIebX7Jp2Q2pfgExJgFaA57U/C9s+ocK/oY1vuJNKBBD
FPFrxsaX5cyyawwCC+3HvXU4n1UwVphos2pJR5e8Xw1xwiE2AjQqmKpp1UKWPP/6
e/ok+F19tNHmGacNxg8bZEmt9W6xcpeKVKNH4c5jqUYl432CknZOVzP4hBZ1PJ1p
10fP6+V1OKzlzQCLiD78gSR+bVNpi06Nspu8wbqvVk1Wz9sL6ImXHjNABhStws5B
a5X3R5bmA2F9ee/iAlFG4I5r2xIGu+8urZsHJOLvvo5kZmc8c1EKX/eZaQDurqdp
MN0W747zWJ8saqK0GGLlS2Q2/epuFBIz4Ui/Y5sGTnGgBfLCFwL2FYEByS/fwGAg
EeBfxjTTvVTZx4YV1K+IPrC8c1jMxZiY83DFyBZ8TX/1p97CvyYgQ6ZAc3g2bOKT
ceNhzHWfP3ALzoJgFRuvt9Eyh2THpj0QJHQG9FYrlkrW9ijOkLpnv5RCDl51KIlL
bliF3Qp9dLwacmRz1069ijTN1CjnoZfzpJW2taATSyYtUvO22vInBUK/JoHc5ixz
PojgPtzw+AKtVmk6JSWJmcrdgoeyT06g8YwdMBDWpiI4S/5iKmUI+cpm3jDjzcV/
khvbBxEkmrOslHzFZXtM1ch4oYMaSOA6GAmH9wHPJAuR+4N9IHAhbqGHTGqbNRBk
+a1F7HxL8MKubMnGhlae/rlq2iSDN+WjP6TU0FcmtngpKKhTUPWoRuPxmMMsBmNL
C4eN26PH5TnxX4aJ/m8RnkV8ZUMQuA+cw0r48MBJuN8g+AcpHJz4V5LUiNfWjhMu
vo5FPuKjRZNqMGcYLrOkJN4pcYL4EKYjIq1KplJXkSqeKhxyE7qNXADKoHF1SnX8
9/tZwF09kqrFepE5Jvf95rNkiMBh7/8q/s//V9are1Nmfi9Wz+pD8IXN8ik3ZWNg
Y8xHV/EIuc0qF3v3goSIwnzwRXDX5GMaIgqEUNjQ2fjCFIBf3QT9AKUjEdZ64CtQ
D6q1L8HMqfu7pqd7g+wv3czO/qRS2e+TLv/q646FKPsLsgxr73l93S/V/X6Ute+R
4U/LD/c2WfqFR7JtcrCnjM2qFRr0HjLCsGdWCVVaUIfWtHJYDtpdQ1M4Q9TG77XE
MkIdOddBLfDaaB0zG7mtgWVnbidF14jg4DNgQOMk7zm+M4Mja8dxDtTWvZN9LQuI
29Ka7biA43Xpi6Q4472Gh0HRSvT1hV7/aVYaFgtbNVUUJont/IimAf/3Mq6qAPmx
dge36PiuJUADTgiy8pBSwrZtYGUIJmU1KistL6PEjGDY+NqhKe4yrRY6QRjYdNGv
EA48EXOSG+Ulx16D349m079dlZ8i6xJvzGULCLug5G82ZUG4Vp8OpbguM8W5RsPq
6y3HWZJJOhbiipa4EYz1Ct9tal0ZsFoq4+V6uTH6XSlVQPDEL+tAyLrvHSVK3OAy
dd57l+HuCTLIz9CMQM56jzsaSXftOqsjs5PozO9C1QhdEFDprbc6cvhzREQNflBU
iIBYXcdaRxyoqJgF3YWaT02IGTjsvUbm+ZBb++EynlehiOf7EEjdsxNQovYDqVFn
bWwbWeGFn2emSI2OP3vK06YY6F2RZQXU8AFjIdSZJh8W/FXFxMvl6Rde77uVZqHg
uPCnxZTF9rc2xl2f98yrLj12z4weKZ571YBK/D3VM3RpQswCrohvH2XoRu9Q2Srs
4Q3W+/QKnG/JwJBeFNWaKmZQJXzkf46i2U9dzR0Z+/Mhdvr7cE3z5LK1cfk8B0PL
Cc26fmoCGGwIEuDUNwd0NhOkj8l4miv7NxJSgYVAc5VbNHESFp0uBtC5REpeG6hB
Cep4TKV6JhiWvnt3vu/cHLe3icTZ3+zPe9TOn102PMIEP/JhWvO2jVaSjDtsduvu
b4zWuRuNfd7xnlpCE8UxoEqBHqQz/nh240FqiTqbO4YKFFDzXz4TAl29ja2R1DhW
0VWyuNS7FzbUDU80u2DY0bUsNRSq+bHIcbwY/Det7jEil15YyKWTut03CvqE9et9
h96yMv2D+keGr9r0uWVpsMZsMweDvTZt2Gxe0bYL/QHBHRFnt/SWH483/I7lNnET
0hiMtk/lxCDnY7PNZV8MsxTFVnPv2DMv79ALHLMMHRIGtSdLZfzHVW68r65gQJN1
LTX5FEpf3FTHq6Ud/HuVIK6Kn0pnKJ8u78um2MbZoIPi5EUNk731t+8qSKAjIwRB
D2Z8oPU6CgWDJqWPVMBeKo+4/ufe7ZzePvBWw7Nrz5ifP9d9vYLY+uFrUT7UuMEJ
FZchzXdlrlykPKrQevlubAkjGVnGDSGgchlUjk18caKE2A8k7uGIzGyprr1zejH+
/4kx9kM6cUnz86wZT/Y209V9oa1Uh4up5aDHVsTZ6ZxB9J/+/psz0++ZOVXDJgKO
RaU5SpaAQob+L3pEyFwuoBggvWYwEt6u83l0P6c1icU9gjZjuNL95+wWNzmP0Aox
Y9fkBGFfbGcO2bUa447GJRiCIEWQIbAcelCUtXK4l6Jeuv2dHvNWrZI7KQEovM4a
JHeXx2SjaqW8m7H2CNmFh2ka3bmA66iq2CrgMs4RyEJkDdSTX2PSclGzeadIvHKR
w1Wp7gkz9/KLUvDXM1yRCk8bkY5KR0RpdEJe1GeiX7qyG3ZNW0we9k/+enUfaShZ
VeXxyaY/2+XJAcYYE9dHbIP4VmbggkR44i03jTWTO8A6pxxtatwqbp/o8zAn7/sE
GqGEZAulgyr+XRnMpWgIuPMONHYeL2cIKB/eC+GObZK2jaIhV3ezjpQLjNR790YU
6uItVY/cCagK+Cqeo4ysD/cIKPLAqWjyGEm0R2XI8+xqQcBQB5dX4hV6hYpPC0EN
lRe8WKElsew1RXmfDc8kHZ6s8Vef72lBJYbakccKiLlggf58OTUikXhPJPE46k3W
vZ/tpMZ8W4xeTZup5zvCLbKVDPgjIFGzcTKOeTayndlljVo5w91ThCwZNJkL3PJ9
DSm9ESxWIsxMtKi7hoyh5niBS+grcIKu+jHpB2TQn+KandbQwAxOEALvIO/o0iZW
qiu6PKvUru5xlFxC1BULCKUZj4b5TsyaCI0XeGg0YY52YDQ29a4jNhargop3d91R
IYzjFzk+6MjgE2btqSS5IbxcSAsHXDm1XWvo+kKvLDUmtEcePzz+MKwBLDROC0Lr
tJIKU/eQXtRC/bqcUufnzBU3dya6arFqMGxXFsPrW58noefv08CKnZlbIEFwjP8f
CnP01QqEomod+wzREj7ZWrI3oCL1efXAmwRy+ttJK1goZu6LddxNMjP3JsVeGIaM
9dkOgBnRsfrmLxZAaHdzuo22+d4/i0wdJjmPeaWkJSt90I8r5AuHdDPAPv5+Lsyk
0T2+5gl2q9B9QnM+qzSWdSxClB33bG7Q5eN+H5favaB83zoezbn0NpFoWqD/tVK5
xNfpbghtx810Og19eZdjeEb7mV4+zovfm/mFEBKnwy9+AkzETl1h8n0hp0LzoIrf
jfsyLvCOGaQz3tKlt/Am7OVmB4OaRpPsDp9adpbwdQBjl6KoFZJ/LJqkkCjqZkkB
R6G7zuo52zeUA68CiW8hNffdoAAJt5d/MaxdpX99+gkFrMBZpW1yGuoKtCBk7ZWt
bFIapt2Xv81J8pIZ1h7X8u7FyovKyrguPPX99tDksixxgOBvUeECb2bhtGIrSm+h
xFo4FLC+UYOUHLQ5ole6SrE3Vza1X3LzuFl6RJWHdtpSLlBbnwHHbKEqW6LA6n8D
q9k2F0EwG0tMJSgdOSbn3USzfRs+44wq8ucUHY1fWnUNbQYIoMxBYrYTPGwKlGRg
kod9DhWmP/8ULbmB7XjzJXItmZoSjrpl2NgU83jxvPikzB8dPD8VvoIB/Y0mtmw2
PevmpBR1xB/nhWiKmvbJUN2A9skOWQLORWCg4WCjhKZWytybCoQZH6k3PmlfMBy8
jxKzMzp3s9fJCIMlQXX45F5YOCkQ1a3/17o5OJf13/lYUpObbHoP1uaH3PDCkxLo
y/xVvNVQbezYB3ejTtBgYQGOLfeVshEqMLjG6XwtbO56I/Ex35Bu5JFSQlga99Bz
NeLdGjxIC96yNes6ylr70jXF8J7EpN8umhEZYahUoM6FYaJZD3D93apEtHJ9eIv1
6XMLP/2f17ex+Sg3yLmlFnsxMjFMMctBnH4zbdMZLpAiy6areK/K5HK0hqaB/ydk
IILzrAuuTdGwLgv8H858PLzn1ieyIEaEGv1lmOL6P/4xXylxqk/YOcVvx0g3XoHz
Pq/GjLLahJup8B+2rwPsjk0JYBpEiR1jeuguu8TN+Pnoi0bAd2wEHop3t9BX3YrD
7/ngaxP0dKUl4VbxnDhPRPcUezCq0r5eA+ow+9TUzQW/PKBgwDg7kaw9c4TCjFyZ
jUXaCod9wVbNK8dzKdkigHD2hUfRFBl1QgbSXmhNc8fWhjriXKYtza6pnm2N6vVb
VFj2/I9iv9NI/tUXVIDnSC0Q3pg2V6hLq6eem+T73rcWY3KmJhOcSnfI0zkNe1hM
exy8eojksciI3A9i/Tt7Xhpa3jeenGU+6JaO2AUoz7ZMTpSbv+8cZ8Su4TCbkMet
HXZMsvTvYDnxQGVFU3ZTpJojRUBJGaSH7VW4sG4l16z0Qv3KY9onXa1wLuiuGz41
96zDCt294eVZ7Vt2TeYun1VxA8Z/VZ7kL5/w8dvMxI9GkvLhbIgKV4t9eA90OvIX
yoDq6ZOtzJJk9C0s0uEQFtsFVR+ei2BPE6jyYikGgIt1tvI9lFZ8e+qJZMxsoYfJ
1AVIiWiNoi1l53U2CeaKa0jUJPVd+lEzhuCgGo0tpq5RhNPb+7GjYDZyDsvhlTLr
ucwmruB+SyNuo8Z58caIQBc24/J1RSKGFNSTROd7sBN7E09rq2gdKI0vARS9jqfW
gxqPyKpZIoFSv9vrwnSoR0zU4G8K1C25rcDv9d5HDfh8PGaIRbjPmLEkAhUokQ/x
wgkBZn9nENZvWZA9rWQFBKi9H2jda2PqYIgvEevj5t0xkEmWJlxLdUCnR/rNwylR
nNB0KMDHaZToPGbAVYW8j7w6BwnmAZZuRDRlCfdg43xadXjZqJb1yAnAPT5A+bnB
NVeZ6pSZK3kATXJelzDdNgcBChxKxnIjv+NEda8WCMGEdoTaRt4sQUl0moo9eQlx
ZjusIuXdEncJH00xkpluQVmx0AulKwxNP5KxZTFoVVjWQGuLx1G/3L0yfETADU8H
Y0YrUp0py36iF5st2iNHa7lbmBS74j8Y7E9tpWUc22K0woyNhi61Q6IhW0GoVomN
RByTf/E5EyQHkkOjsJSgn1cwmXCZIHj6Dz6YS8Uk2/yAeA6WBAzAlxIyPHhUXZ14
gk+b3l46zaBitMXYNsO3gAQ0E/8rEWHTikcxUNKt9ZYhiIOL7qbvHC5gBbYjEpyv
8G+zdPv4tta8ZMiuLrPfoPZ+5s6EcYXjTpyO5AOf8I7WBLXAOeob5mh5UqoEkhAI
5VwefcgevTkpennr4HGtPnd/3E7pZDlXcDkSsgyf1ZUaCH0OHiW/5OVqz+YIFdl8
mluXvUZPU1SUVWwi4aZY2PHo6xzoVaGzKyVzX6B82YSXFIqROimUdn0GV2TI5fsf
PwocYYig2i05fh28OTdmBk12qWfI/yEuJBpOEdiFlOUlEKWR0CJ43ETSIdG7FPt8
DHEXqyHOqu+bqxsmVvH4HIWw9uRUNSN4PYBBj4i+NsK6X8ujayKtz52Wey0bCWnR
GAaLzIVy9ame+X+2YjN1HeAfwRK8BQ2ukpXXowpk76pYhebZIpaQ9AraxhtcG6Lp
26gz6Zh+D6nLV9WkGEBKdLkGoyZ/9c74NJgjWmIuThPMLPYQtlWwUn+3KI4Sx4iJ
lVxzcFZuv/SFIyPa2zV//V5cn4nuLkambxzphkAXXyV760U4Fol41+hackk3f9cf
gpPiBP3/GgjV/23WANyUXJ7AOSNoquUyz8KuaHQKFIKB7IoDMCOgBbK2gunzyDMJ
K/iR6ZXsfDG/nBRnzIB5kMz86w9AiQi0ev8kOzk720oJlwtTj7+gH7arehWBkqS7
HpidV9UdEwK5seU9UgKIVQNdN3gWeYsJjRipsBIThnNbSwO/3QGrHC8Hxx2HRbcb
6dkkyB33t0QWu6wRjVfNo7DkP/iESvsIKePL0Krv392v79nGDm29mCxLfKsiFpdL
hyJOnrCpFYhuavyi4j0H4RqWBHmXPTWWUmQju7/THolT1fNHx2rEjdCT/uCLRY1N
6mU9lA7AqcAt3q3YsHF8snlveHXcRpRcmg46xPI0vfEb2vTTgTPdgM4dPsiveNbq
bshUtzpBtfsswHq70C4vqIe9ttZ5gpgEUTIDEMEKQMCe8qBG+Z4J+SDEfbNuIGWR
J6y5/WmefEcI2uJY79qujnUxQIRjLi73hepPwsT6Qhe5+oo15/Tsiq5JHSkR4KNp
ZWdreAZJVlvNjxHnoROtHSH+T5UKZ5qsDwNgdPj66EeYFCfuYmY7sm6irpj6p+d3
5VWasZgVG9oF9kDZsi/b7dOdzyCd1ec+cxwCl71iKT1xg3PaJrzvN57a/LvaffXi
y89DpIaA8YePrpwMzt4bz5n4CJjtdkDYOQidLyl8LIoUMpyESNX/rAIHfC05Lgdy
9ylI9UVqDQ4uAymDoJZbUzwDbO9yR/+FAB6YTe/C5J6PVnaUC+kSnZohhO/5t3Lz
oJ2+rff5mFDdv3sDLxftwYYXWsvDFjT6HPpR3MGlTtPWXz7emCcFKaS4UYNkY6Rq
i+lcxVa2I2hWPjERDGpYjPsHlvqFSb4MuFhZeOUfPxAnPZZ9GFcJwZqqW8IkQZXb
/trgz4X8orhnLMdmmdH7qFZ/GE8OatcgQ9cGOnW+QBHrmF3x/3qrnbdlQF8Oq95x
M13INaTkK5CjRHx6bGQpa66I3/vWSOgx0+wIFd0i+6gm/+p5tpyQJe14D2east3D
SwNBMa9tCtxDRPbifHXKZ1Exa8qxgf/PaTqMIP1ra+xuCjttQ6eNlodhqDAjLozH
Qy8Ruxjjf+wmjLm/A8/XtQaZMCibUmPSXCXanzI8f0gmYgJ3radtIUn8DZYsswsy
LY2CrtTO/YcOd+4K4s4YV+7xvIQLZtDK/QhRAvtz/+Q3sVV0AdRGFzdKuiMJ4dmP
j+OjffLba5rRcB3teHVA9DlspXmRzNMhIlRs+MsA6XIm7kz04EMAGfmzSV+8WJsF
xGKtDnMvQW5w3R/g6GyFwiRWa39AeBFYT7wzUsF7ZikjCnruPlcL7ibinONYRCvK
0nTENFpmpiTit9jVRwCpGlCoXo8c7UHgaxkRuFDYIWoZ8XxzaVd9PRwepwqa/pjZ
wQBWfTqKfcO3FTuSMzTTQofqu1JUEl3DMiO+glO0uzLSKVBPQGMShafkkQAchxJk
kb1l4ISZ86bZucHyYVrDMztYeimzgeULw9Z/dHUfK9E255pkqrhUm5L3X0c/EZ30
CN+oUN5QDRBDzqxfeTeR4DjwrUzSvpyE2/U/sXeZ/D57rIzKIiffNMEQz5FebXPK
6pHlpUER2TAOnHihHHEZtQeJqiszNDTKQIwCRfjU6S1hnGjMJUbLWINTGW0+3syt
y5AU9kL3+AlH73Yl2C/wygG2mBeXBoodx59XQNcGL2Zy34c97b4hn4TwiY9r1LRL
ti1E2h+Khvh1UZ7yo0nMvNA2z89vRCAS3tgcnKLMTLU+ntn3meP9fEXsGbj+G7ww
phbODdqBQ4JqfOEtx4dF5AKqPLqYqser5w6THVI9PGCsZeLN54kJVfs+nwWaGqoO
vjLs+Jn0ODSg6oB8qFgPpJTN7uPNazr56xAdhPldTbhGF0RulT7/14aRowrxBd1t
t86cYrwbZCzv+1XQhgFWsXlIoM9KHH5iEsdUYNPdgQjdrQ0WOjs4YViKznJeFSPC
EBgi5Sq50nV6ooGAyJ4rdemc89k9EUlq8jDX1R+y7bqeVNs4xtcNqqoi4KLuGfWN
nofsfeNqOeqBorAUxdg4meYtnDT0yGjETd8GBc+2wVZIT8g/qmTPYW4HvN7oWt/c
wccjSg7e9epUmBpJujleuD2KM4PmwW/ebLsFF/qUc5qhGlutuUF8L7f5JLrCNAOD
9Xzeo6wBRnnZRnJA9dARMM1yiNvEc02wsGm6upmUZbr2OVSx0kTpdbb/GCmoXFU8
io5LvtuEEo7ahw1kP9XPg2dSLFxHZGG+ZRynL9ITa64I4T9v0X+b55BWD2MigBdP
EfgmESDfu8HHgHNwxT1p7Vwa1PT7n9E56375JQ03DrzWlUGUn9QyTziYrBcH7irl
PllXGzs8UopSBurPsmLSflOPJVJ1wZoh/lw6wV29vnB5OjUz0mLXoyT8U5CMJ9OQ
xbFx/dGQcWtkMFFva3cnrt7+JvMSJdsGWNkQnCYtdmZyS9aUb0mFb4NInl7mxwFz
u1/HQdhdymGm0Px8rIkkT2Ti84wx3YQ+S7l4KHzv/LCPB4OeoVkAxIgyEJgX65u1
1VHgiQgRxu8cS4S4Skz81W8y2pHCvEy5Waj/cJZDpyLVbN1+Sx3qDNaNcirTF7/Z
krSl62fX1BVhZ0856wg5ihMEy/i9bQEHO9PqgSbRyCGx4nOI8melVwR3hxDwE6ZO
WE/9DlJxqaa6WZC3CqedOIPOgIyVWzC6ZvNOZ3PozHMRbggLR8RL3A1LQhYp57/8
6MgBK4843BS6mQGEl8QX/Z/8L9uv5lrlQ87tO6ZaxwxWRSRaTyQP3zAZnO67NaAz
UbpOO7k+QwiIl9yz+ColO0TqdZfR72K5X23qJr8pgDWmfKMOfYIm7rfjN87ciwc7
dGzGksTTkSWW3unGOTnnCTUewINT6ZQ3PcFmD3CjDGoIGPzmAALsDeLTtJdMcf7G
kr87BRSSKl+OeEIjHTn+T9xZzSNIE0OAQTQ7Ls7W9PAe17L0ZlBPrfVyIiugGMkH
Q/Y1pP290OALexDUZOewKPdnVeDEHLzhG8WyaXtR0BqHkyhwUx4HhRSxoaxJ0XUI
X/A3hgtnSFcFhU55N0lr8UDvYzUwlR/nvZerQm5W+LVzkKfuxXHXwWJGzrFomTZ3
UF5cXq2f/iFZod2RjDy0vdMDQ7zcw2aeD1CEws6tC3UGQyEwW+Jd9rdqNTygHN10
MACcCPuBgmz+oon0GWEP/UxzkronN8sW0qNXwjRXW6psepEqk2q4+fr/MwE++e2Z
0MfFkYy46QJsEG02vuv8ahgZkQlTuDF9kkYii1fNKmOzAndcyIoymuZkNmv9fcJB
psCkHLb6sf7GAeivNwymjDCMbxo3UdM00F6GPdXHYVTu2fh79iwL5KnH61K1fY9O
tr8fJ8Wt/nlABB84VWobfTJz03LVf57zBk/WYe65UWC3wlTkeV9aXs5pvleDUIQM
cw6OoQE4NYpXKRcEJIohkkEj3nGS5nWTloDcN0v1yLwVUYZo0kTvlOEuEQ3t6fow
anBPupH0AJs4Gp+tvTgpBfSNUBSF8DFnXTd+WZFu/++XI1O5PcIt0OKTMzgxA+ML
M3dcnm7pWatfT6R5SjHrRsBevWq1qG6CPQfW+2C5pRqnDj5hwry5EotCl5RwHvZy
0Q39Ik8Kk91ntUB9DGpNWy4p3jU/p51DVfYs6H/E4a6bjt0DpBvi2QLLR3Ql4T4s
0FgpvtIZ/d6Ln+5EPvvLiwUtAzsVHXKngj/L02tNK4iwLNjG5dRiVWpf8xeINHgq
uAeLjXYu6ke+xWkcfm0D59HfgeN9seq3HWhQLFmHf+HJDCTxygeud0kpFMVE1Trm
3afMrDMPj2kVW3K4S11iIcQF6qbbEbQTXgbw7o/FUcP4+MqUktN5ZOCRltjGWWj2
eGBHscNMyuE0kaPttaDhQU1PQ5/Y/+A9kYjIt4fAdpVYMSoKIJ4fVjxaxQSOKYJA
sJf+SsoX1NsXBkSOChmv8y9iOCYGDyRkWlOw1+Ong9q5eRljaA5WJJj57TTMLDia
aRBeEp0QmwjtBu1Wc+ZcgzkTHBcokSaczrWevIdQ8QN3frKquc2gc4a0NSI0naN+
31pRLxDWWK4yxZ4GWTZ3JJxWiJl9KuLhRY8f/A1nPo1mbUfsefRLtC983KM2aukT
b3HptjjOhovgLw3MljkEceVTHDtKRGStnUG1YpfyFhCRZqdjl5F7f6NMd5PPdsS1
ivxmuA3K3czSc6pqybH0B40PR3Pa1lB5nEDntya+4lqedCNNb9egkaX42YzLguI2
zBNUeCc1fmVJiuE2I9RuVSGzG3q4V4LKT+P0NFEy58YdHdytHkHgLKLB3JqJOaAJ
xh72XBE2b5PF+og5vM5yHKjSI7v/LuzVJXgGBjKYqkCaqp5Pnkxu0gm/QOjFehAe
a6OQYazisGQbEOHOw1V+a4DGBiwF4RVCQOPSkElrRPUrsIwLxPVv+f3F9kT5nEw1
hBuxJo0tlJOOmKkhp++8YLC5/Fwmncpc4dV0mO7DeUSmbPbZWXzZPPrjMpe0e4O+
JiV3hlSxHDEC/4MuyfzS3uhYXNTVEGCT8gFmHS6tQTVPGvGeOZGwm7aMDMkNAIoJ
ileqB1f/hNqXA1wVPZ6C/76+O6ExgWaPhR33cGaYy0GYHJcYilWx5KHXnbuNCBv5
QGEmd6KmkW3b54DBwPXuKSljin1Nl1Kwkefv9AAMCWOcGMNHsyMfI1O2os0iGvvG
zz6stLv5JeVsBA1CmWX6lHz3QjK3Fk4h14whZ5YkR17vpY4cltorOkdc0C8UY3tR
2bgHZoP7961OawzQUrHNW8900Fd3UQK6L8Fi1lr4W5DLI70zjHKKfWNSFPEutTuD
vmp7PfGMm2K+pF+jLl0N3eLw+Bww+p0TCITVK/EszvCTSj+/wjHCUS30ZJN0HguU
ON/khC8Pl0+dy6iZ2Ao+2O3hbnHBopxKMVr7X6OwmDX9UE21Q080iwSLcN6T9UEK
P7uqdyNYwYqVcviQoXEN4c0ZL1A/1xRgEAXnhKZK0IFKIecBvRC4+vaohrFUK7j2
5RmzNxZgblxY05TFk9FZRV4dWQ8Te4UPrCipvZ94k02HrDu3ZiF9+Nom12iXwuCb
z4ndx4XK5tLa/SyirQtlZQbEHA7N9tsOe+ya+5TT41KmceGRLoVvBodePQC9ADjv
znpid2UiOkGubZjhjd6iMp4U0XMYjMmTGe4xcZCtSFYzyCry1P18X6Z2TY/eU7lO
wGCoS8Q57nOJqnzxOVVuQL6ytIbLw1J64Zk81x5Esb4NrOkkadacAP29jiPKXKT2
HaqFM7K6aH2UzBaUqLvSnJKGPXoiGicpOclLUKpTO55DNpPzY9mE57Yg6KUe47fc
ugVTWqS/Md6mZGp4XlIk+RoAYUplXyrQJKXXcsdoCuAcEIRY9G/X9aexE3Nj/lSd
oBmv8O3PsQbT3nz+2zjpqq1u2ga8on0OfstGGk03M5/lI1uBMBwkFyDA0FPHV3yp
0JNtoHTjNIfUpBPr32r+FFkxLIvJrIyD/SD1ufdeCaI82ny51sb26D6A8Xx2YZqj
Im76gCKTyOTwkE1uph65LfOS4k7dXP/R6/dS9OGFS+Keza5ab4kF/dst+40g6Mjy
3vJoOopiBKlh62pBEFVw9O1sIKIEK4t2kpxZK5XsG7Sl6GJjX/aPcXgmE9gQRgoU
ckyr/AMZ9o8N4GDhDxlamgtpl6+Y1DwRKv4En+C59ytw7o6a5sR00Q98DGL/fi6D
fF5nTL2WaOMwtZDhj2iVGb0OD72WDvflP4jqTnelKAjk95Er+dQzyPVf8jUbH2XZ
c9MiGFfWjelfI6vOZ0nwrA2sLwJKVQNSEUIAliXH33a/asseH8EomOxoLPsoQiCn
mx+DT7WuoP0igVtbWmGR2KC3u7eRFkSLapWf9hWGnB2sQes4CknEvZ+toCLUWQOz
S95Dj/vC8MhFMhIWi7BqHvfFD4Z6t5S+kkFfBHOv+KVKfjGIr4nLQVtAaalxh5Vb
kSHsXsz7dxS15lUJ2T4F2PBlyfAb680PRzTuQ3kpH3Z6SefqEpRFlO0D5l0xy/3t
CGFhLJMPTdOvoGw7rC2QwCRtLf74+xZUefQ4HG4YCuttmUoNCambXYlGFybvM8AV
jQfERnQuS68cEYwQeu1JjachX2nr2dJxxODI+0SU6AdAM7UWk2vImJHesQXI0O6E
TK5I6VeQUuQpk+ZnHUle0murqlG1iLtD0mvXJ3S/9iQdxTj6LXAjmBXM72SNLHza
hsxPaLzVSfVw8I4Hiu5ut/PjkdIqbNXzLs4FfE0x296bD7ekpO4tzl5Kc/sg/E7n
JfBXPYN2IMU5y26gpdvt4PzRamnNiPGMhedOD1MgvW0yia29710inhafpzoa7eVr
IDsZ09Fudi8VBDF4Xz4meNo83EWzoq9kLtBRMWS0zKcJ0hJ+pbUIJ2etW8RBsNt2
XVFi7TpiE/vwclh0iNWdDuZ+3WKxLbBfm8BSXDy8NYiuSQu3T2qTP3GYZuSlo/lb
i/mlkekGrTtmXImOgJa0sG/O0CfSegCStoCahX1jA0cznyRm7MLpHVgDZXSaOVuL
W4F85yZV1bmh5Jcs7Lgy//EQTTHs6gKLOLvC1CXmNuXTDPhWgj1pPTuP3FjA7nwg
b5u5HoE6SlFxm+dMDRRKZCAfDHo926gmFjOpRFrG38Qp/s/3Fs3VCWSyPQJclTqD
DQiVSJNPPfJP6eNSJZZuYBPCQAOyYgpRwXa9z2s83VCbIXayY0hB14sk/OyIlGgr
OV0vokrSAZej+mmIzeGWBjsamxug6FnNFU5gOOgY4E+FW59syZeZ1TPLcbC7b9GV
aQfocU7pA++8zNB2jqKod0dl6MT4rk31IiUtWVQAHsK4AAOwPY7P7nzf+xf7bh3l
5YfxeM57jyt1VER66lDvVXRX2Y4LlzUf/HCO6ueG6rSoFuXQMHRUcqB+dUoBIBVI
osj63YSbvs1LNXt0KZVviW9BLZsjZh8j2jJ8TFCgEi2EL7IDGxJwjpjzFhdsk4Km
va+bP3AGWoLOtnSxdOVYk8wjUVu65Q6qe9cUPsHMq34/gH5citfozIGa5ryqA2S4
XwbhTUkuTer/iAS9IEdM5ONgLluIShLcSLfSVZCpxDqf2W1N+cBXFPTtNA2YEyN7
2xrTuC0ducri09OC9Nt1ruKDn9LrRGC6YMV2U8ztZmRi7lpJBZvdklDl/e579n3B
Nh8WtfVR+3Y2L/Km2fd2nWdmpIxHF7745PxZRfMGqJPtU/cgyEn7rTZEl4ecVHlY
hgVdQ8CLtpmQ1Y03AGQQgsenoAkh32i5j70CPBy6ipxNfrTt1Q60yU4fazr2q9Lg
6j6VKyzBE8eEu6+PCeEleC4sTvaqEKWPlGEawMtIP/15bJtvFB0XCX8zwJ5lquRk
3h/PAZizRhZ1crTcirDNXjT6AYUisyJr81h3FQ2DjpfVbmdoBHhzuqB24cNk7ZwR
3PPu5QJir7QLK7vDjgj2okgfn4a57X8VI3q7tS56NeaR8eWRJWi06HabR91O/s+C
IkkYyeMZEF2c2dGMTEWM5YGoITK0CpaApmsruR7tGu3KuM8k0EY+kXpNX8IcGzRI
2HXqKvVtcf1b4H/BOeaL6OSNV92qJ70jr1J0nDrwtlPX6IbjLN6UC3y5Uv5Gl4xI
drKjDzs5CoYNH2+DbYil1JEUJtTxF6kv9kHth6J0n1hENfjpOVNX1QDU5gLDQcqA
SQO6lMvuUHUMNIs6LbEOAMdxzs++wjYn2ciFQE6s1tuEiD7u9glbQnEAH7tf6jrs
Wt5SLZ+JALTOEVKCrgAGpIDKadU0IpY36SP9ycTalrSPkz1EBROxaEEmCQO3j5nK
ZtJCJBLZzcRvTmxcdHg0cbkbatS9846LtLJ3bgcX39kkANqFLai15x3F3HFhvJRw
4fx51exlQDVBnEOdXPdZRMo0oKyZgXinPheljybn7diHf/du0LPSMMwlrnhL3l8V
hJleYed1NHO3habExAwnjGlr8R5ygG3kljcVWg5kdl7inNOeL+uOR8S9xrzU6QT/
xGPwPPyHCVYeoG0qpswQP08T1d1dBJEp+Sbw2vQcfzbRUEgr9e2GMoKfAiR8ZvBS
+qGIsnaPg+NR6tzySaaUlvMNSi8UXwfz1Ms2gpMVXGzXt05vfb5SORF/ymZ3Zq1V
7AoIg2y4gFIe7bV3ZuiGZZXWkFZHw9WxNa2K1jeuGoVA+gdBfMJvllCcZBUNc+fm
0SEqtHx93KcFG7p9sIGhRn6IvUOM3S+YWG2ns26k2o7+ldiYdEnU2C+JEx69WtK/
l0jbIbZBtJJDQsN25fvgEPh1MQvu8jyheUxRU6GC+JbAGUsZ0oY0DfROuquJj9Le
NCYasdFr4dTMqJk/EuKbFyk8faE9WKBIxMHJckmmnjUbU+UDd3urKWYhn2hd/ijZ
q8YS8gh0jD36VqUShDgHVxLbMify6aobNsJ/7Fkm/lP3loDsIpS4vZ0czvHnkgMx
OIJx3VjKkUKNwOIfQBJXCuuk1YKmTkE9rW2IO0RBRMicmXgtZ7C65TH7TpPgDgfP
a4sC0IAFk5s2AK/ihGddZdtPXEM2N1yh5l2sk7Esb0azXnzPx6ouFdufkKrRlZHa
W27HhT6l5CG8iIjr6dw2wdIsb94n1eItTJbBeqITvuOffmT8c65n2yMMM4lWUcna
33osAaPBjZLGZDoHxtIzGcfko5eKooFlbYvCjuTY29HNZyIa3SIdS4D4wNE1niKD
YSyuFTpBtjde2VBMH9zD996wQajs/dfSHBol0+EryUc1/GZ5+FLl5kBq9AssP1Ys
nk4z+3UDrqPcaV7lvjBxNGd9Go0sEiG2xdqc+yBel+KGo5ENL9m/jf5jYMiHnsMn
RbjqtJ9be0Rp8S+mudyPQyGYv3gBuI3Z3Wu/bequ5A7eCzikVGc7he9Wy9biioG9
QGZDm2wOBaIg22lrKUI1uvV9fzI0uuKJyZNW6M233o6j+yn/+ov15VnroKN6uYm1
OpVNwV+FHM4YdzBdr0P4zPD2k7Gn7btxtt7UXR/R8HOepqusiilaZ6fC4fgZ9a56
8eci/q6WP/663gVWslkC7mIwRseLASJTp+390k5HM+VBMZMXqmYajYqxvbPcf9/D
DHybt7p2tfqzSa9A/sGRaY7eCm+xY5Eto8UaKhg0vhQXrHazs9r0UaEgxZOVSppD
3DRhtkUHUMeJLT7TKXOhvMpUN6Itfw2uIsnrIIBKbZ3mrlVuV1NLBExzobdvDD8z
q5EIGhacKOMDx66pUwlioucDNdKZlg6Qo7INqiupgpcSosfleLSZqbMdOEyx/dwa
kMxKoX5nzpHLJUPI8Wmm6c/tD1ACLqzeA+Wb+S72mZDVmLGh2KkhRDFmQVb9lzGo
t4vsrqTQrema5SR3LyJtOpU9vFgnL5pGAr+DYJO/D+/y2hUBkiaopMYbOE0tvjyH
RGI4RHKlrPRcVPn5dDqAhyG/zLGmg2McZzVkOuCULPsmgMdHSo93/MV7eJnYfCNe
u0PS/pOpvoXuto9WCAkhRyoWODB4U90wDj/Kgz9CdotLWdXVBBRxl9HnEycjFwNq
/3BRnRkygLrcPrvXIkfspbp+sZK3RhwpoWbweTlAnlpdW3VvsxdU2H+2W9TCHTd1
rXHVaqhFNSoAnQ/Aa9VrbW4SJHv8wP7DJXwgOq+Qf2I4rZXXZX/UP76tPYBGTOXI
lyYNP8/Se/7evFKj9xJjWFkKXtBbd0mTJMRBIjJXn//yt3eX0gokqITqYTL+GaG0
Hq94hIg2M5MOEqPKNUZ2t4XTkeNdqqZLxcNj+4Xj0ZV1+QpT6ic04ebNJWnyuUV1
rZ3fNT43NBEguMx335vCyEEJoCdjBTOeDp8xfBlXeK9u94uKwhbo29wXyWFGGM6r
LN7eyktuL1jKbOtwNK4PfIzfq9ud2DyiK8eXS6XNcVMs1TEolB8NWo1hYOfndevu
5ds2Nk6Cb5rGjvCw/UC4/ujAoC4Xa+Bl25F8ny8JwBJNWCIPkER7CXRE+WIZYuHW
Vz7Zl4AEHIxdIA6ELW0KE5ESSfWl+Nrw0WaGyJobweQ3gcSnE+4kWmygeUQGfhZ6
iKtqQAIdxPCQYyDWCuJoGebcyltU3On1TWAmBYkMFLRg1qF8beUyyB5f4x90PlOO
KnqEXoBnRfA9c5/FnX/8F3JkKNPaXFD5lcqOhyL7kQ1bKU84mlCM9Tm/WiKaUBpy
IAaWDPUAzl6vGm594Nx+wuCMCFwr8wqFeF2/70nYk0RX35NdQ0H0xQe5WKUz+R8g
4r4FgkFIFpD+1mCF3xNC1W8tGOZ6oozGeT7j4CpeexSMxboEShNFqJ1Pyn43z72o
`protect end_protected