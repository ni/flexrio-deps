`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2320 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
sJVlH+palpt42Vz8KbH9ld17GZ1B9nuNYVrSZ3Nf3XCx8sjSjO90bT1T39xTczad
VAG8kE1a3ev4dluBEP3GdzJ7/T04ATjjOrAEkAnPvW80n86hFPizAkqYbAoxzrqj
Y7h+UbR6EbSqY2X0geeTItpbIy9M/DcgFDccYB1weYIgeUe95J0ETGjRvxy9gD3o
A0k71AmlXxWDpSPiqPo3TA3TReEOJrTnuqNXdlDuM+Nnu5V7C3yWkSsxfHHYxA9H
oKdSFZpIbgNKga4jgZgA8LePvXnd/LsmG8SEGFlr/ZthYKRZQxWUoLMF7qhV3W3K
2jwjmrW9blkC7n0cB7m0Efr5bfOXTTyOXc/0lBo7ftXwiHdQtz+ZEVtZF/kYK6OC
E/LnNvq00yUDjtbIlYGy28RlbCfOvZMBa98jPo9n2GSMjs0KBR2NQyNSYRra7gqc
V0mGgFphmoKJ+n2Izq/y7QVrF947HP6M7JkWw2B1DSlRkH3thFWloAqAsusvpejB
YrfvXt/FJmJlD5hKf6vreIY9K6TnWDxuc3A6+tYW+NPJmKGpfWkvIWhWU4Wx3vLZ
NPZqArSgrzR4ZZM+I8WSCuQDcDcGb46BBXIL+XTQJ82/ZSq849okp1osnjwwu10a
4t++ZIGjfORPmi/HqLA0jckt3VlHbU9C+9PDB1o/eoeGiprqBbiZfyklLF+0NV0K
yrjA4EVwwGWKcJlt8Gi5Lgx+AElsXSZHpL1cwXoyP/Ra30AnKiaHvbGQI06MYXOk
6OtSbi+yXVRsD2aitx19XILjKkAZy+I5PnjuUu6y3nf9BVcTxbloGuT/f1PQoHZx
eD1LHjGXrGco5VIJ2vnG8eGIhAhsS0KeJpzLh/Y+RvT/Y7Cw8e6KUcQoZFB6t1IB
zQFEFY6s37fjnHAy8+5vxzYT1oQzSlbyN9+yb66xWUL5LIf00+5XOpViQJD0t1GY
LC1BnAj1/ScU4RloccyrRKMXBEeL1QBoZ5dBd7e4sF5/4EO/9RZoJMbYHAihdQ6o
03RgEfe/mwQJwqJUPiyauJJ9xM1GIN00prkyrJ5orTO14pIKRdOX/BI8zj7GQ9uv
kEqytRixK44xCUEoSgim1jmfs/RR8BbY9/5jB3uicffGpgJjpg2I5qjU2+NxNk2H
tNJzo5Dnpi7cIwGFCJp8kg4KXGsmZCAl9rm6AfP0h35A1z5EQb/sO5JxBiMl2UOJ
/KBRdYh3pyyESlSy80rjQYZefwX6bGcBlWvpmj0g7PVZf4d9U3l90Qm2SZVCHzzi
PaENuVrDNeTaChIYY/huu/E1cxPrFdkRzPBVO6Xbms5Kky1Foq6URPdZXlb2jnkj
mpbd6XIm26lRKpN4RGhQqVDA+czK6J5giun8c3Xw/vPdlO1sTCHy9gqKPcPOD0lR
8bZYON7z8Aab6A8JPdtkKMRuVUP5x7S0V1BKEBaRz+vahxkvxvSXjFPVEz7wRilO
rHv5ta6wRr6SXF6JA6AXWE4URwULlrPDagbn80h9LZ0ouzcZxl12UzSsjxPFraKq
xJV1TwSfG2898+x3z75wQsaJ+KVx2nEh77xziY4tni6xYWbKXOBsjQ8xAaA5Dqm7
lywGUNzRl1e129EFwqTJNTfDJg537Ab+2fsBWyfgTRPeEgR64folvsihjwnEgJ+9
g+ZEfffkGJhIsHin81Tc+Kqz08XGvXKPnYNQAWOoGLPD0C3sGWjYaQzTNESVbS6V
dRD57x3beq4+S9wrBesXGGgdXDeXTdu2PAk8uNBQ0QzVQb8Avj/5QXkWpvP3hvUx
td2oig5bTM3x/CV0GiS4qEYHARd0yOxFsgv6diqXM/m0pwN9HjTysr0Z3S12/LxM
Gcobo88Rz3HIDIWjCrwNo73UYOoOPvTGfILbDIKj2BtgshQ87bKuBK8OhpnzsXbs
PnzZ1Wktt+/VMqGDzVekDF/dLgsV4P+/VMThtRHEpxwk9V/5a9u0hwvV4osDXzY8
MgeldynVJiE5Y0uOJtrcbq0OIwJ8s2ew/28nnlglbtXf79BG/hpv3Zo4xbpEyd0M
aBlFaY3PlvLdDeJO/0afSX+dA2ghlm639FxsUeBxxgOYbBe9LNJOR4Z5yzA1jLrb
RYhj54be31dZREvSefth4CQ0yb/BXlqCWQZHRo4B+ITQRKisnAQMQ0/rkpAAXgN9
DQI58qYgr9XxoeB/ZEEEdw5H01K5rKi78ziJAJMwgaBPvC/mVw1LJxpb/61amMf7
s7ZeXumG2U39gvYvJ/iLDNRRFxLxBiI4zAAiob3sA7Ubc0FDaTdlGtrfRWnGMYM2
VP3etxiak2u99vseJWe/zcKWrW7x2D/vQS2R6KWnUBBNqH2I5M/LMFey9g+h68V+
bIAF+42FaFW+y3cz1yRdFM//haAgGjiqR66mJU4VpnBDkUIppIB/YlhJHoAc5o1p
OqYWRbfLN0YKPnVpW7Fz/BRR2naQGkEhEFeEhHHqX+4pI4QQSBwzjzm3J7VkPK59
AF8CtWC5SnV93mmy003iS07bU9Sufvzvf6w+LDImXdUN4/zw7DGnQPk3yy+LMkcV
B88qOY4W7YAEujzKMGTp5zGGb8MUU7NccnwYpzIm+hqe8NchoITmmBqHCU80rJy1
T0tpHck78zht2roQU5rA4049HIMDZSeo0UnimXXQMJ9mD9xUQ5dogTAa0nSGAPCu
H9mnOi0Kj682PN/pvRzcNLkAa2zBFRsLOTTQ4ty37eJxbx4yjbhGDBMLW5F2hDoH
LHVpIOLgitCs/n46Q6sXIf8VsFQycalbXpUlJ+nDe+QHHMUJsxNIHy3aDclwywW/
en5VlUNtKvZmulXQM4TT2zbtjGEGY6Ap8Dp30bG4NSlDPvMi6fuv5cxu6BpXTTqt
GTJ14REdd85fa8oNykODUlHbrm3Yfl/AuvIpKEaIrtn3q4zXRWmSY7VNjEIi+1UX
FWR5qFqgPG+9otwDam8wMw==
`protect end_protected