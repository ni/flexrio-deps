`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36368 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
m7OJaCYG4D2XeQKzWhbYg0V9U021acplTU9OksDDEFGyW+CsZvnZOCx+2SvRB3b/
/D3a/1OkGVzjPWV500TRuhNR263jTAkZ7YrA/TXoRVN5eoNexbGPf5YSizhqGIwL
ce1gARwuYyrkIqB/wk0TVgb2HYwOLlrXtMkFJx6nuQQ6uxwj78r9G/L8ejdLkqTR
UDmDO4TqJQjfAJJfsVmT0LtxQagObLKWY+RSwrrgOwarD+K7DtjnFKOddETkzOUp
2i0MEFPMCMCfPlk7U4HNyj2tZt+CpkfdP9pOtPp1l7BhRpWwZqy5y1KMe8IIijJL
dzoB5Kx8VbEnPWXRw3H8mwxPFfmeCC2nyRZZXbc4+GGVpKe7+BDJdZC3rgZEV4Or
UAVDmrvofyCtxjQYL+adJZuVuGH6GYBFRrQ8iRKUKa582+5xQteilku5+l1/LiQ7
kcJ7r32qDkis3UO7/8nZMuqlYxc+N89Z8V2qUsTz1//IqVHLK6SeKWscma+7VVob
doIVlI4NmTT1WUWU8Lx4hkpfqOlJfh11gZRNx5ujNTdmu2aOWNUcGdXWv0dk/vxr
Zw20S3Dm/i0sXO3TQ5iJpxLHDp3YBSKzCywqaK5KtmWC12T51XqPWmpx7TXp2cyw
Us8UJRnB2ZL3emTC94PnWVoe1B00LtPK68vf9RhWnRnjMW05ZV6cgKvckpzSw8sz
IzpQdd+4qSmqonCGTIZaCH4sAm0eVsMIkiS6pLaLfLHz1X7A3GWICXckLA97trZx
5i8fVNYNnYVYHod5FT25cie56/pdkmGkZy6I/RpkNtyBHgdnfigq5CwL6sotR2IP
iT8kdgfSgMH3/6kDouqQkW5jsYBuwYjQfjDhUZlq0EYskgPkXSyvrtFN7DAQ1euc
KI9fBD0AdGpVpArHFSmV1Hlh2dD9PxTS/v3Jb32fp/Zi4S0Jab4uC27QwbLP2Ig9
eeXBsexiJDyYp107yj6gKiJPwgBcGMQWFs/mCw9y+XGiJ1a9iYNyy74aBdUDwcxa
6JnKOh3Ej7q5qy7MfBSLSoRsRqUW+gqrjxhFJyDAslYgytZ3GWDbsytNQTw0H7sO
Lck7yOpcqCnUmeN2W4meCEfOaYhZZMWY17fgcRSyWi/Y2RQO+TvqfYw1xu+aGEVp
Safn+wa7XqrvbME6NKLafDlaHHcfc0z4UCjmRTrYGr6AW5wboqRaguXlSjBy1TPw
5ro9irVhTGQeRfIp91Pv2t4JfD+2Mbkebis/itroQPqO3es+tnp2LgYVtizE6zMx
ZpoUqLP8D/H7Gz7oPbjzglF0u2pb22fWAbsmrsF6lgiaMgrham/WO6iQPum6lZPZ
INuBo/yym37BrefDSfw3Z1dQ9USh+aqMqrsRUS+TVn4jVLlwEmGRbfZe/4W8HgnD
XsUR4pWKg2skPC4f1IdSPzvKMYHcSwrizIhMUpDIdDYdQknzNRsSGKNzKuUm9sUQ
iodedzojXQCVxau97MUZZxppi8DyAMW0uBkDMrgvNDz2D1hmcYycgTZxQpkUCe8j
jJB4tCLEWaSDE9xlqq/KH6halteyUYaZV3jjFrO9Y8kKiL08CwEpJ8ldkPxosbuv
aW0VAroqgKgF94z89OJ1o+gWwxN93Erlr4wZnJDpcqJzyiZXtL8onhN1LfY5y3lU
6a4rGAiUH3T7d+uUZ9GFcRPvzzF1VvsgK0xzw264Z55TGlw4fKTBV+JYGbYhfcJe
pDaUTgs6jKpfKkEIwBk042BE88evSRQFRCC27rVksqfRr4+zEuiY9rMzlipuW+sw
59zWMZW71P0UREg4CVkpMAnM1LW7H7Yzw/4rCrWXA7yCPhgfVOxie64YjeGxZtak
NHnRkqJOnQOHk3xejq/NjzaMR6/IMdb1NiQqp2iHIHHjfgD3w0CjMIqzdEDMlsuo
Oz3Wk3Xl5BeYFmKfquYVS9US+CPy323CLXzsCTenccXHYHxyaDET4YPqm5bEfVp2
tvHP3p+RJH3RyemoKIa/QXQWmVmP8cfvtxM4eCyphMS7tl1dq45JLO9Dz4iCfBhM
V8IDEHoblcfK1dVmXvOJksmSgoGGiH1IkpuQdVDK6kPY8PlzN1mUC9WVvjG5af1X
V9v2Th/mYW8MIeOjnA9Kp2+/JZ5oFn+hWtPEGnFvniWbvHQ9kR0NGCySvzEya5kY
h0+4f9WL8rCt7PS8P3fDIVvizLPv8chXr2ycGkWHSo2OY9ZIWCy3so2SmKgRreVd
k+NSfuPX+5z2dMqwFS9VSrAkQhUVe9IiB9XL9o1d81poHZ+kT3yFexnXxJZaLYly
q6NcZKePX2A4O1+QPo7JKsn8NKVPcR/LX6++TmLI6bjtJVmd3i4UbmVYPyQjxxkd
bhSSKGZloPugswGAuDT9QIQhy4uUZOTXsdmctGtPQb/oN5LXoVPjF64zTqBFwpzz
mPYc9ZnI/VwOYHg56ZLPxL/7ruOet12XBqRJ8KXPg/JVq7iNgfz4Ia2qPeSy+J/w
bovg5APqL7ojCpZkq/kHBUVjjI4EoVod0QHkTZD4GWEQDsZWeyUWfpxA9wPLI6e8
cUQAPiQXk6jrqOmBHIVD+JeHLDsbMa9gHVyfNpO2Y1LvIkmiDXu76OcOLVu3tMbH
gPYIm0CU48hpDWJvAqQgKABKqyPwhIhFkMxLAkNlnKKKJ8MuzM3CKB6Z1aVfLAkj
Azet8y2seeSY+XCrtgUB3mse0DeQ+hmOP4zcBLXDLA4d1ZCkOfIX9qXjwhRGXhz5
s8/GvjlUEbwCOkIxF2000TgP3oBSNF2SwowZhO0RLzE/HhmkuKcyYhBlSd43kEvA
D96Paw8vKZNJPB6M3vxNGSuxmYya4hOfdVu8vhPv3A4oIgbvxAXpNL0ME4HGPFf8
yuBY6eRsCAiqRS7td+n5bNWBIfUdRhrk+MqsN7jEzuRm6hvCzb/aCkhKF2CTdqc+
eapPnB7tLyGzJv4aZ0WmbIegiqC3h8TSb/M0I8ttwzmW2gevjGyKD2RJgNVKCPCw
XHnNmsHzmp2SZk8c5TkvKnXP46RjrLsVnOHDOQEdtdmgDvKtwdjH1aQA+nuUZACy
3Ke+5UnbvcX6PQH+OWFb4PsWi1Wvo6UTiCfb6HaihN1Ol5HuBrDJclMm9lbEDMYr
1HpMDgZr4BxubQUCGOp+kG48UJmTvC8t6D1FBkPAc28UKlPIbT3TLYfk0GjXrCXO
Z3zuKyA4Iw7nVU+a7sKH1FHXdjBNjdhvDFyMxmT/lZemiQlTReK1ZV0si+UPJ7QM
bbR7Ot28QxbLkvvU8nJdS2cMeJDlGqx0vZy+GuZbWvmLyYeO+yWlJThRQAh6je1l
eRbHKYlFFFXvKAPYRppDBVZVcbEeB9OHUCs3SxEbLT2Uk/72MkDZK5fsme1Zua+Z
sjNNxJ1JZJshAw0jZN+mqtqVTb/F+CKg3eh3i9IXLrV/4f/8E6PDGLS0CnTvx9L2
hGrBYm7FJK61T0LHKjiYy/ewNRJm6Em9YvBER1xjLf4liJIyqhjfiDobkezgMinv
B7DUrLnsLZ+t+tnWRxEh+RFg4zjSVosnCSXkb8mle6u2u5EawadNeJfBRiVhYVwO
pfWgh0jN7FOb3jKrlSotK4ptAcmgtC43Aj977aHJplGy3xCMd3tgs4FPICcKy/Nr
oMtLGokPT9H95ZHmfx9fLSBRpMTrT4xv9j8o/UsY3E0kzgpftpSeNFMKmXkKbRem
utLmInP48QSSHK4ZFnMxD/ZvGOtlvUCX8E1xk0XdDB5QR4Fb9vD+udHyaEe/1e0F
73rh8ZcwG5q1ac+3jHNALaUUdxR0hWI6tAMTwCCbtnOCj7cyEASHHDbbKatCilCY
zEOlEmbouKlA9ITOdUKe/mey7x68hRzqs7cQs/lRorzkcv/xx0KmWhjBgoeGdhyd
iZPtStRxaBczvFa/mO6aBmx68KitOD/mnNI4gcrsevMGJmcFn8GkTpxVYokAAk+Z
ZQxXF2ZUPZjpRkps0+zNacdtKbQVFqkuGV/I5f2IAhKBZtZ5MqEfMzaA13QqqObW
guIAGt53j08Q6vVIo8bsMBt6yRgoOZsZLpczznqgkYel22amR1xZpHd2Xn8QnFv5
fPSCwY3OxhPxCWjwB320ALxbof8/wB2xc2j7d/nSkkbGcT1wAHrt1w2SiL5uzEmu
8oHLO3x9NO9X+3Q73De6HyJ+ZHJ4nw2dvFnT4dA5/z0UfMZ9AHB3PgeNSzZG1YTf
2xZboncQFr1NZwkRoDHnlYCfuzB5CnsVdeoA0uVLxzMN2aoWO4X/b0VXIsocqoVI
i0iNOA9z58CNKmQT05BcC4ZhlAAmMqUxTTOiFytgQMAh7cYQUdsAiEL30O9vRXWT
jnNkZv9IaezUucMrwvaUNLHVkMEh8s0IVPzEwG/3t/8HT3O7eiHONdlgepmfVKRY
n99lQQ9c+D2eZYz07tKMnHbH5avjlxz/avQ1lvd47OfUoSA8Wi8tRedMgVB3bCev
FOz+bUExPGwe7YZC+kiOUY9nVLHy1NE5p3hsb9BM7GADO7qrTsSfONRfccIVWbR4
IO73o0IT+Ws3w0BPi+DtX/K1DrNIBCMdYPh3mxAXwgMKfLN8bqpp6eL72iVNwKrr
HOv9KS87Slkg2i/ZcA5/5MVwFyXY3FigiE6UWpXg3BbVgjyBDT07B7efbUVLppOP
kVd4sGtbJvN2huKzCLXTR+/Nz1ZgTxaWA4f4MnvoVUUmKVYTz2ePjMBN/N+Hi9sE
QcVjNNATbcvfiqrNoyiMghuYEVQNy8fWV7dED7PQs9qr7XZuWLVGPPnHINf54vSc
63dVVOet0A3focCRxEhLnweaKA0JD49oBFdrfpvF77IBFHMSQapWKDxnMCacjl+j
yfB48iGcGzdt9sasWhGCh8aoEWe8AxbBYsbChfh6fpnqaVJgWK5M2TUbMppSV6ST
7+0lKkeWi2+KYPaSpLgVEg04+Gv4CIKeiMd2zKgjZ2AEr15ogKALpZ0V7JPgavsN
q+5LVBnuZJj1c8YRgpcLsHCSM/ympmer+OM9NvEWpx0gCjCU/pHChIIq3xVhbZsO
/0nroeU/YsEtpkfh5oyEOoUBgZJWhYjPKZrUF8+KR4OCVy3NQsiwltfBsDjk58nh
DjmxP/Wn8sdGsnwcsYYqIZwaQFmh5pDxf1KOZlk1u4t4qCEJULfW9qdu58Tkzm/O
02wqKhHNVo9bjlM4ac2Db66F/yBVBzQJH5Wt6xmURWVnbtDDtcuPJK267CCOnvpt
Odoe/f9bUFtav71c7xYIiEAAVeHLGXP3je9CQVV1pPApktrCbrLOudaGLolega8I
azA9i95MkPOeDnozPcikot1HAMLkwhJYoLFlekYZo66/em8eN4opbU8P1k68gvwl
8t84n7fqsO7Y4JJe1/s69746bNn/nmj5okjA0lW8vz8gwxqgR4EdszvGxQuoVnBy
SKhrZ3Sl0DwZkeiRtmfOCjP7l/QSDnG3/rcwg1E7/stPTcaDJgzPcdYNsxP9tp38
Yr8YQLlSTtN/CriTz1z33Wgz+WZ+EuiZzHiMnYDpU96MC/1AQ6D2JbYQovC2NIXN
fiwvJlNuwh0/Lec/nQXieYzvH59nIRDY3UksWu+CUDvNifccEeRzh4nNAnABcWJc
YEVuJESHHWXz/5M24LpkKTA34vWJgamK1YAkn/2xhiAEH0fe4mChqk4+g8AhDIoY
1lmAFPa/dKwNukxUFgKgrWFRFs1JiAz2BDPqDNa0jZzFu0x607nEYEYH6G8ypAsh
+BTY5fGftH8z9g8Giy5GZosvaoc/SnUmCb9djJFNjdLzuP94Yn9ynhYtqgVLWE5O
VUs6zbBDhVBalHSOmSEgo/S/TLFjNsMcr+V6+JUIbf3SuJ21nyAw+Vcygr4EoZLc
+m88icZJwbPhJT+1INEUC+2mSlcDCtND/zZOwUfnw7lKPzx3pJf8jNoCF8Tu6tlF
SShZDL7CQTaCyBWum1jBB9FrnwTt/s32tD94KacFZ+9dddaspgSerl0uQOW92AI4
klMA3vkO2iBNXnSWGt6b1C9gTKyPVwpTs1y45vpy+HxwqZEheLFnwKNAa18gA1vp
+DW0fGJ/zepqOhaoA5eew0NJhp5Ik6tqt5Ng40cXzNTQ6pr5LgDVL8jEB3GAfKDZ
G8Bf92nmQL1yZflSeVnP+/Sflu6d9fJvEy9gBOkneF+DmyK59CGp8U9gU1ghJq3U
b31mwewjQkRyFDgMvqZhSY9EarHw+PNodE/mohqY6q5cj/wDwImMJKDrgz5gCn/G
zeUinmcBzjLXHHgiQ76l3QbZqvvxKdIU7G+M7EECmbWJhv974HczNZb5toSe4ToY
15arLLbEPmYfaPz3oMEqqL278n5m4y/fib5N/WJjcRvDF0SN1P2CmDJUv+dpZdMX
Zvbvj5myIQokylt95dhFegodD0lONN0yrMuLOCRivvsWxZQgYUr8NZBpO80MY5UZ
nmCBeIrxkbHfcfyL0lWVyOOm1snGlR/4Xg6O5p0bJB/Jn/08Mwc83YA0qLR7/QlN
1fVA+l8KH2bgPtZOWS9AOzoog/KxLDqeOU/NlYM4gInhY8alaM6kGsBrkdRtqDjr
bhQw8ZWH3VIoHAoh81Zh6PNZ75PwRwjRKe5AG/smm96igw7/4FTVmpA9q7vsYGAo
HVlnxOyT5fsSF7K6o1obE7NbxsNb1ucQyoKsma9eOTcUIc+IaJuL8X/b6l8EFghb
DzKGwiyOztm3bCxJnJRLQhsIB9J7wFXeqImLUD1k1CjIDlQkTXFm45u/KWOjwij6
OsNkpLrtSJT8IcgeY5MVCMWlZ67bEt6dOLnz+Ul7qO9IamCy0rnoDv9fFnG9jh5R
YlW6LfrOAteJ5kbfTTBT2THyt9RBKkbg51KxR18XmEtpWZzGJ8yl8tzckQ9JBSWS
/sfsbn3/6NOfXKxSXPrivriZwq14CjnyW37VSZl+8D8y1wbq9uPjsvvYp2oRhasi
0YPCH6ZaNZJQGQnx1VxkYOKoJ3JWfV5G7wg4BEikv554yx6z7OVXMTyEgBTOLqfR
UPDmtGd+D7AJXCoOQGK/TsZCwGQ6xsGU7AAMULhi8Bq+EfSps0aPlQLWOkGl6n88
FkZwPX6m5qact/wA8TXQvrV5Dg35C60ql8nwVxPGt5XDDHtpfWmrkUX2ARg93Kpz
uXdQem7SO/aCDjNfti3wqM9Bh5Xfp9emrWOie+CW8SGH4QjGuRoCEnCmaTReqsOn
siKs2KYZ9lCgnfdV/pr/91erFIyH+8HNsZ1T25Db3YcBKvwXYADOBqnX9QToCjLi
1KnuPN+uqofobaJQt7wEnQI3VoDhXLOrVOc9JaFG9JmahNtEf4tTYOV8ZPN+cT0Y
oCu15afIkAj+dBuVz61X/wFt7wShP5bxsbPg8lexGqVJFUSO9fvAGU9HfNBZdn+a
xTgzds3kcU9ymU5/ZaRfoVJj6vxxtufWn9D2ZMvspk6qknF9fSW+3WGsLerIAgo7
aqPHjAT17jUrghsH5tjmmImVxt/9AoqWFoOvzpkse11IZhlyyZe/iE07gTEcFjQF
j52WPg+5b+dYo/N+pkEnp1w8sGm0WNvXsHiDqBQguqZZo6R2IlLdXulOF0Qas1Tn
ZhQ2d32Wt+eKXhbLaAm6TCykJk7jPPT+4kl+SPaKmSHD4X/kX3d8dDHeIxvXvi1f
xF+Ogt+cPDFcwSthChjFRTPJdtGhGWejFM2VH51Uc8jtK9gcS69pUxxmqj8CazR7
/FjO+n2AH38nfXBk93EV++ZJjRIhntYd40y5u5eUa0Ann99/eWNahY+10dWEZEqJ
czYEZpmfyZn1Piiy+Fn0avUKWRDzl2ip1G9NPNIzqvNqKJireVoWA+G77SHGXcfr
Xr0wKL1bnhABD8Nx/sAJjEi3ERexdu72NwQlXALmf2o0OlA4RRq28/nh/Dih7puB
qIqu1IVSwLpm1IxgSk6Lg0cNtBCsQhLC4qxQO6KR+dRi+rqdPwXjPPOV20la2mnN
jDE26QIlrX1F4D1ehQSYlGDsKCV70/e00wdNfeDb4JmZTyAee2z423JmQzDS0aAT
JbkcN2wikb8xWPtSGMptOAOy+K3aWV0hn3BZBsbjS4zfvPT2O9C+RKgaK8+5E/Ti
uc0eKeE7IAjtHCmQRFTu+YcisJQkmi/Iz65RbieYoZfsRJAcE4Jjr6SmTEFwrQN7
FYVfwDZ8D3bHN1t2tVZoTPuPrXkfEhnlFD93fzk37v1cxBYCESRwvEbWuUCyRL/k
j/PKp6fkGO5jDjupJRLgDR7mtCymT/aSZhioar/54HbCURUwiVWQHuJodqBcTbtL
RBBy0hSHHU2q2vwLMVHIMr5y9YUGyiC4hBjtYGdE9N4EyfhQUvgP9Ebd9CB2+H6t
4iHInTQfX5RecGB8Cn2Ghx5NwZ3LLXTc8CcgDCSISBtKd1UzayoRrjNFf+CvPMc8
lpIHWm7KRD1rgFsLoq41lki5dDjWzWTXQ1qeTkDM0K5DbXzi8Q1lzzSqitcdvua8
j4zqYPvCv1AB62J2HZO6+l3KoDolvv9eUrJAoVc5nPW6jM9DCXoxfT5cEg6buLF4
6saOvSsrb14aQmStc9Nw0iaYab89FcFA1EtTtKsP30dgNV2IyWNIKYWpS//awYxr
SoqJ/hvbMY02ndUKM66/P3pLL+LHMbuu1x35zhE2fKKxfEGN6kiwgIUCz0/vyasf
FZiJ1jlQBg70l8srU16mQaPVhUuY5tgsHCe/FSiX9p1WLo1v3I43VIEoDweem7AO
D7M76GvGQg4akxht/gRMB37lIv2eRArguEJYWEYazfgqvG5s32eHNv8kGcvcRUmL
Rr5mmpTBkaX+1OkZBnT6DSl6StTIoeOZFpZJuTCKY1JybRxZrFW3fKIERKTJOza3
0zT4uPEPrnlHJ1t685d4XwcNtNamXNrevFwvBGEMbSw/4KudW4ZQcINc4LlDaKg8
iWkDCBCi3bGtoDb1y5HlB9qReLtmhGfr33tK8hQ8tPw3R+zfEyogj3mo8dpEG6cH
OUYYl7WLGD6xVFtD7KtNTaNa0YYtIYRPtTeoxDV6eNgRUELYeLOJrCm5wa0zBH7r
49T/8T3SWcX2dhkby+3XeY8dmQUA2X6CHc0WRSggVy/LZThTNCjogwjgXilzOgcL
iKE/RIjk4C2E4rXJEEZUn69eaYkMZMe589CwKK9IO5T9G5m9CvW2zHo3xW5i+PG7
iyVcw4rO6cSXCzS73VdBxXM1Zup1NR/iekKW9MBbw1ayBtQ+BmrFKV1mluqoVNKo
SBKuvDCvAROMQous5isL3wMa6Fliy7oqDIM2fgM8bvZVX0l9mCZy66FwXi6xTrTE
XLiyYmm+D6zk+kiU8rfcaGrljnU+h7IWSAhNSoBtUJYILLSLe+fJhtuPTaTFdafE
PGigC+iC1R5wp5LmgbxC+vIs6T/r1M6rmProSTyvvYg1EFi0RutdruMljkhbAcO6
RkRpQNAv1Mg9TYlbObzXi3WTAun7QKlnM7GikU7RFfx6o+nUtflJFRUKB2mrHEew
MduH8JCfDAByltfNDy9iyw4oD1STZWKLkeJElNNU7i8pF3cV7afwtF2xwKQTeNlv
3Wl73CPfBFwxNtHdH6Vn+SU7ZialFh4KmC3MijUk0cDn7TfIT5wxoqFggLgxOaJx
aEaIBuUpD2tVx5mtSF2A1D+FavPnOjN0B4IOCRsvkPHejgCji2WXLRt2FX4hVYEU
QgIxQ2gGpuNGVhyRY1g59II9Lgl1b7g1ylwY/Fy6gNyqNc/rkdTePW7VB20dgY1o
Tw7zZuKTmr6xu38NIPoAEKsPCDoirnDPw9X7OLE8kig8QZdd3viQHjZDsc/V3I3i
6pOy10UryXy6IqRy/qciKDU5bnEeU2cgh+k/346N119jSonv0xHROlvSbcSlXApf
9jP1W3CrwSa2TwFP+qlkYGQURywl+Re9Xe8H7I4OIUM99BuabD1cgcONiQ4zLES5
KNuI7J0+x8ZAd48gIokXVEuzjxap5R4q0JTudHqSCMB1qlF62S9IKb85KjEcfO9B
aC/uWc0lEY+J/2+OQmNCYcsjYagvCIm2ohzejihDm4aQ4QHPxsODEujW1e6r1Uyz
mgh+l8VPOUxHYIA2TsZR4UgsUfexOti8ycZOsZIrgK8ad+CcpI1KXTI/ciRSHlna
bOCPEb0E76jfNR+hnIhGnFztrm7exo/a0uhcSgiG9/i381lsTkwG6b3a6fWM8bAK
A3gZK+azlazavmGwu6YFDmwAsUhLUip215ExapZRgG6nTInw/VDH6QV4oRvuxavT
PESl7AQuyH4Hs4c+YnOKAeEZbxDNMAhIsTg/scvxxG6oYBCA6/uLxf8ax3Zm9SEH
tbjpwg2ETrvrg6o61/soDD1SbQRSZaSpmVA02GRJt6Iq0UV9Hv1uUSOWt4skOurq
P/MPIGJB/Wl/LHaZJtdLAv3AsD8pSdrE5CcDKK9Ex64TI8Q6dxke0NralaTMyi7P
Js+eJHQgXcLEJPcNTgn2nxnYP9sX2R5/5lP07AAGIoXpoqoX+SzTCC8+Iz3JW2G6
CTyZUiyHobGUw9r1NkqxuF+svQYCywlDFcpjInWtQsdinl5RirE+cMeS3ITqP729
BuF0Si28MjcvSYfa+VUr6yZeYEDw5aAJEzL/Zih8pSxbSzETGPM1uGDSc+nV6abp
oK+wXGyIC2XXGCZG8a5eQs0sIHQ4uW1L0OX2I6c3AQj0M4LXMfkyM3opFP4o/qx4
oLR1e8f4ftd2O0Rag5n34m8nwBWN9P4227IMHSXon1KBfWBy/U9eo4KaSse5uETj
iAHoOgjPS2OrmEzDh8ukEkO7IFKOMVdkBDfOrC2mwr3j+hTouF2Olqsn0/vnyqb8
ZfUSSqsrI6kauzMuO4AkzgS/dAWN7Yetd7uj3vzuGlRxXz82jsEsqyVSk7mNT1OH
jf4a/wwv044OyP664nT9SfUlEbFVtW52I+4RJQyQXTOk2M1oBR31Du8g0ELx9lYo
7z9Ad/826YgAsORyFYvBY7rmD8VBxleaxpjIlswjbeGMvV40lmvWKx8S91mFCyQh
1YI4AkPpxZJSrIi6uXj7t+TmUSiqILA6B7AHgQ8nBBsygCX5aPQIVL45wX32LuNL
YELvaKlhGpMk/ddLeKXLFnb0PnOZKB40eX+lCLrkkQNEQfAESApjHZer0d/htjNQ
8ZuXD2i9sn+gGzwroruCdOEdMclHMQrb+vMDxLW7OU+lQjjvJJpnN3bKkVK6pUSF
5Qv4y2jO2X1tLzqoiWvsLzpWlbsIqUcNlz+VgF9jf0SbhIo40YS8rfL+p175Jx/d
XCws1/FrQv9pdJ3P+878BC/cepePW2hmSqEPqcznPAq/kqPWHFsU/nrFmdARQB0V
Nw0KnDno1KdfTc8KUlZDJVsNnWFKFALn9ep7LLXLP0i52QmX7x2u1yWAI5KXPz0D
FCWjoxqhvgIFD7BuUrU0JTCRbDhJj++vuq2xAntKlw43b7ErrAjOOaX/gehZvW0f
Dcoyl8UYRzzssxQjr8iCH9BqdJRNESs/rk/k9kdqVeUrqIOtchJjIlu1yZWyDM/R
n0Lw/4sS/x9n24Mj3EIZPPTz8iqXO10vRAPmvsXmrAH7sJ2xiaBfCc0kgDmK3cK9
Fp/DOnoG42hOGRYMS7HKPvJr23vlnA+D/ZORQPgZ9zkirQHiUGWkzlopmsaFt9k1
ZOy06Cn2fiVCFmDk6dAs8HFQUVKReGTOqGRXqgoqjL/xYH03Mv2dPqRZ8CzF+G0E
168oNV/nPmcsBnQJkxmnsD06blWSV4BA7HbN2xhAlzyE57wYhbnRJpx7PmcAYqWs
XtZB9A/J2CsZrXOoO7v2JRqzDCpzqNdcI8lBnykM0ie4/pQ8RCjZO2/aXBE6cL1g
cJtnehVfiMZsjZDzj0wXua2OQxkZKNUI9jrrGPINLExNfCJZlE5LIeTuMod11iJ/
8aVm2xH5KFCKjjWZVpNF7pOJsh7lOIUK/yeJWLrI1lOvcEItdtu7lK7tF2t2ECDv
I/eJbdSusVwtewFh6jJlFwFWbjchWDtDjWWOxOU/l0vmzuPb5szTxcICpUKlUEe1
T2RIEpvew5LJ3UGb8gzlxqrqOJDJ9T8k6PhTZnPh+Dcz//FJMUxe5qGPDZbY4fBf
qGwiNp942DYpZfS8GZcNs9SLUKgssWYBBHFxZQQHSuXuWS/gvjY962olCKFQgCTN
X3D+mtYnBGxfRmS9S2qOthgeoibmW8Zo4VMsho5ZoIFsx1MgSO5A0nXzjSorvc1y
On9epkJPCyeNiU10X57jy1kQyKDBd2z/JyFDZTTunhzNf/7C3nfldXBncG3vQHbk
7xH/3P3zJF0fJPSxYlnNCpA/R/924nnN28BATkPncm0ZYuU/LQVr9v2wZLINoW9M
s16shODaDfJqMryWT32j5BeeAudo8LTJfLudWqItbKv/nvKsdzLBHsJk0X6HjAYS
prWkkCXk4oP2c1aMhyFhQDxhUdyfdgBeFQdky9aQoK/5MSUxQTEOH+PkChi+BHts
S3njWtciz6wAGCsOmjIXTMf+ODdD/63f3taRR3LfWTRbs9kehSCACjEsscQ7V/uw
Ll7Sp329lxtzWUkeSUZExFfIjfeVPj33QclxsnAkV8LrxzgHL/0/rY8RhfXVjdyF
Ed8AKUgKBNExc17c//4mY8STJZSk41BjBA4a0rCIH/v8EynnKYHiX8V5n4miittu
bgU1sTMVPku8BYlWmJvJlWGKV8E6PNvguFmhckGRpCF+/Qe7PUl0b12woaKsr8Nx
+KARpFed60NeDYq/Kz7Nts+83ycT1KRPBVrx5+UXFxzGFMe23Pq4/k1/MmeWkdAo
TDXtTAz0CVF6uoCr0rEtnKYYJogtU+96tlmdpbJRK3x0EQlwUHBKP8Y6vLW/elrz
QA8/AjTprK4FUoVpxV/BjT/PoSXEugMsS3rb8G/B73ZC8yq+i4UAaechpt1dM33z
u8gTuELmSV5MYRpOpb+9ksLyaWKVOyjXjIrjFtrYTGpYFtQvaFGFFTwzOtHVa1IZ
MXWUnKmxYXEl10BZd2m3Feba5BduIksFCS6mRPd6STaHWFsnUaRmaBebWSJVofHE
zG4a+XTNcih97Nxcvnpvektod37XtMr61U5AIKqLDJxJgy69O4na8JgQLP6wjzfZ
xoMC4UZEJIyHJg7/UYE7j2yQqFs2XDcvIqCaLpzRSiIMF1NvYbmAYUKwCyYx4QHC
tcleSen2zNq+1uIwBoB5crGvdIe0DcM/qODfbTkYyBXzu+hVamK3QH+hGKa3COSG
7JpV1IwNHK7qU/eoZqsW6nrab0cYDv42d2451IM45x0U8+2r673cv7tOi1YSpAM9
sbbV7l33QyTVG9L56LCn5n75yXbkaTltqSD1diRCqLLz5ieWzAJ6KrDA6jTDqBQQ
Hm+HXwhO5qQYzbRICBw+bEit5VMcnzHSRP2mrfblN7z9F+bMk94jQgXydRBp+CJq
+4BK5nqGHOEjOjQYEm3VK29lDKjWLEE4J4ulYZlxNAqzFeaTblrEbp0uDh1Xv2wt
k+LZwFmxN9mojTR5W2SIOxy3rAcsg7lrCNOPRfo/AXrz+Rf+sB+kYyFOQWKPaseC
J5LqoeFaRBw6y6678k99nch7RQyM3LhItBjjDKLMIoChaFed3aAnwcakByGsIMm3
Z0j82pVU3/xsOLgFwUXKJ77Nf7PGIIccNIn06EmbMGuDyOyxbYktlVdDnNy5hDRn
Q8AMZd/EdSYjMndDwrEe5rnPf4ElHcHFoSUfIWaaWSjygjidqtSg7/unOjSdiRg+
Ul7E0yjOJQ8nFByHqCAEkw3qSeHcYX5H/0+AwVpETMvtUGLUnCoS49Vs/CMX0kDP
theo/E+oRnUrYd0Xi4n3mI033mN3doWh9Cu8U2mMBMnlgH7/Lmau3cablSTjGxqq
jNZhbmRYAK/XbKQg6XVS113AduRLNZ9UTPAiFcBN/Cx3Ip5i48XHe6SUVsWO25Ts
0H5/f/eFzO3F0FqWdBgS+vCkJbql4tL8KH8KWCqC+VJwFugw4MKXTP6voDQg+hRg
JypCIBzybvUSlD88/jTs36FKVp+XfLbs9L+x++5XMLtVVSloCFHkYib9J3aGKOxB
9vJhcLAHQnd5xmc+sfzWtTAnwKQte5fwXvWV2XBVwV7l3sdiRgE8JC5/+qEvzhp9
t3srODksLBuQbGs/Q2r+uHylfTfmxxsrfan7v3Y6L3yXYLCJMxHPk1gs42LR+jhP
Hhtn8uDH/QGjWbcbHJD2g8C+xlYxBd1MyXUEiMmjSMzXrNw2dJMfurSLolgQVEbO
wQK/0wMFqFaVQP/gF0iWYO/6anEsgRlqvLNoOTp9dX2plPWc4hOG0c4ISpkpO/we
XV4ItXTaroIB2u8AvGJuLQgfKM18uuKIZYx86poRKk9pBoIVQ8I8QMCGm+Jy7uC4
NM4+an/Ac62CS1H5oUnjky3n8k0vtc32/VphTqTLbH9SMmewauQwkQNHqOcswgYU
CPbrsdF5ZqWBAfVPQI3dP325Jrx7j38/wxpPROlpxCVE4l9TSbQavZTOEhKIOPON
ki5nu0FXlcAWyBZ22o5nqfewY9qCaEFXxpVp6C2iMQUvEw4gvZS+ulDgNvnuXpQQ
rlGwxWV2ANs1F5bZW+FWiiEuOeoW266cTYUV+5VPgRkraZO0EtTvMu5m6TyAxnUa
B8kaZT5AmiROqaveUaI1vvkKJTWafzvlBMwvYljNBNTP41P47HI7T0ADfIMeTANF
QvyU8H8ENM+6QjZVsYDkUh24LzX0C63eFfFMrAPQ6zI/ZO9yD8mz/itfAdfsyCbD
qMgvlZfhZkdT0l0I+vkASmk0yhiwQ9pRtjuIULZ4O+tvqb8p8ocLgYk/VK0XKFVc
Ui56mKBea45Z6oLggzsaYO/tlwNnj/QdGXVu/w27vHd87S6/LjXx4G4SdefchQGw
VO0lhCuGxvejG51yqjl4amnzhPRa+YfqnFbc6fBay6ZwKYZPhx1kuN4coNltp4JT
8fR4DxVHp20G4vlMLa/si6ZbtrTWMrPVa4XjfIhjtmScs2colR/VY/zLQ8UEI8hu
b3LOHtm6o6ar1Wa3oLsuQPyD//atncqRNyyZ/WVe+S3pXgD7hpYdMo8l0C18TGhm
3MVJrjFlRe+TOTUHm29g38v6uZqVoTKNHmvPqlFJ3NfVDpCb4jjFDw0LDnBjYyRQ
0VmDWEvsa5tEHvjp5E0gKBpkWVEi4uRdlT17XYXTGNcFhJPsDCaUb20lnaMZUaVB
QBxZvkIDErfOqLI2IJpXyemvuGpDPFV1NndDOeBiITmvPh/2hs/tRZH0ABjeUpNR
w88UAxeCcOqUKJD1FhtXduvaSrwOQg8m7i1G8CJiB2F1LpWatCtjD4xoUry7esJ6
+AStMdx0sCXO0eUUs6zzuvcX6fVQZYUqoSDFg2k5Ih+FmSgZBcQQcGb1602Yu1qI
zpddYMoejaoK1O2B6p+rOzdTGezBTZ/26926DmVVTusduqUr2ukxT1ngIhCUwxdk
89amnmqKbZE9bApCPW1qwARYBjU6E3a6PhWcLb8PDitK/NqJnryfApotsZjcqgRG
ik9ZOHVLWj6J6Cy2oDQx4QCMFqTFw+hEjKZmbqgsoXMBiU03CNg1jT3cL9aus7jG
1taTpxAFSPOIzt4FfSgLoTGSSrJJ7b4KtJS2PxehfCmRKXMAMjhTBf9DtgwDExrL
8Y1GLjVYmpRj349JhnXhwZ/TkOh/nHJ8Pc3bUGrz6xPU2DdLgEtX1kuo+XG9mlPT
qOCeC+3cOG7DmTHifXBRm8UOkvo3opoPHQgLDu59rHbCZLr1L4crGZk5wO0pzv9J
DKEBqtIfk4EeFY8+09Ja217Tb3uVaz22+g5Z7+Ig90dtypHy6DpvCrLmLgJTiE5G
hn8SK57GSQuF2KW7wTrFI8KrPHpjoXOh/ARdIwgK5tpQdKfPUeXgExpax02u8Q9T
wEc7T2WHrz3Q9JrHOzOR94orBicRj5I/Flj8ysOvVAToB9D2UkgxeQ458HvG5WH5
+T5N2j/9bedWlFGo09G7xW8uFhcZN3WefE8mIO7szB4+74Wf7QE1QTEk/TyIC74C
KqCZuPfMZwoYPnwa0dhdr+UGAeTtCW8rwZdG+UQTrU7KB/vTg+570rPbBMkOffQB
kRxkx6pnrqSbTWlgZnuOhmgy0ft597v5VmeFqVcSwapaafaqv0rbS4bsffq+xoir
PXVn77ZmQyuyzGSohvu9eYTDKOnChfgZtMvfCkAGVtn031k6pEVANtjdz8LKBin1
uqZA5gp554CgjNHPLIHP6cUIpKbieCo8sVS4UZspjtUrQnwmow5iweA/sHGK/qet
cVSurOKz63GH2YS9AA0Dtd7FaHAlut8rhA9tySYchlr1E+sdS6mOBUv4jHWiPVp8
ZqREYLJ0CadsJfojNgJh8MKnKGmA+u0WyqAu4tkmoshXKbaQZx5jFMkKkeX665l1
+WjbHHXcca7QRtNgh7Aqa5R61mzHfFD31MvLXxmFnSOfwtMlrCEjO8HLsVHLXJmw
FgYgIsAlRlfjMpAZBY/4Pc1qdapRy7G0/G7rKVEV0wcUgdMVmW3NReOmGSA8Ia21
eOk5Uc64Rd+I/h1T12Ndo9CGRSFnJ1bv6z8epg/5i+ahk8enEqVfXr7IujTQQwIZ
8Cv7bXE0bRXdVjql6g2CIuHQEGrnyjEriW1lNg80IURL8PilZM7zbVa5zz19sYLi
QzlLr0iSv5kgF9lEQg7M3Y1WA41JTrt67GvVPGaETBW4ztOkfhFQTaiQcS+YK0Db
ZJ9NA0rzwPu+7tpvJaF4vmlRuev9UMgkb5PDKFeUCXYR9W2XFn0uxPtwAdQaKyjP
QJh3RcHKvmM8hiDv6kZke//JKecyV/Ea9GJfFu8ief9lWUzPep3s8R463ekXnZ91
p4VJ10qwTypFcEv3W3a6l7scIyFnrVUx+IgJ0x7RfMpJa2IKZzzmtpyFRGvSjjYI
AMbSpP0gtn8AYdub+pFR2NkvPSyKLBfV3jlxClGFCRcR7mjE3ZDL3+ssINKJ44Zb
pHcimx5iHXbFqZj5wMbdJTmz032+ztgEMmRYKn9wuL3r4ZakpOmPFsr+FCwBnSLP
wsChEpn+umadA1ydFdIhE1Xs4Db+jmywrnfCyh4k4Y4a4kveNXAWGkqZrJBdEyaj
69otrumP8wUIPuEk7fhaXIPv1ZOARXMKUc+9slAGQ6y/tTFF2KFqcOqOAlj/uxz4
angsIQffpFLbvglUxWJZ7a/uacNZ+zZmu5mOlkkCAMeuw+/BAs+3oqy1W9cYtByq
BvgOSHVEV113bNbQr5bQ+l4sJxul1Z0w4UtLLHDgwToQEMFeJrHUZzg3tGhtGsVF
+SiOQVmNvIGLdL81nLd89EmNe2x7Ic7X687z3dNWkP3zkfRAtFx7kyoZiase4gbG
M3EktW7tKF2v6C9Jfq5p8/2az4nAeY0z5hTBUkVk48puPXvk9Kb0baW25izGS65n
6O7sy5G0LtDGX8gXMH9ufVoj0rtgSR5SpAWlG3IeWVrVm24sej2FNxkAe8WQuF0j
DZl8TwRy/SgrkkcnBeDrsSmYIM4UjXekjUHA21bLIBdmnstxzUzeEgAgWPg//jQz
0qAggb2w3lGMpit6u36neyf1aBLxDmmDH10apDkaj2VfhZ8tURX0IA0vk16wIiMj
ci1mX4F/Q2fujHNYqgCZkhlEprrVywZjlTZO5SZmqAxmuXjbwa1q0toAGlQrZD3I
u9J/2RLygcFo7ESy71qnzhS9rS8YZfS/hKXgqgtVV85pf+eA/kociRYA1LlxN3HH
BIDc7+Z1rZsCjmWl9Ol2sWxwhGWiTMbF2weofOOePEA+0VVRTthTaUmQZOFvXkJ4
qtwkfG+PrNy0X5aHSrxEy1MunZxS8D4tkScAMlLY7KCkw1rxZphNQqH24wX7XXAf
Mku01n8EkpsstfwfUm8dhOoHV8w+C9TJVHhBXLSVgU58agz9ySEbX+04UaA6zWnb
wt+aKFcv4C4XizPbSDo0YlE8aPZx2ti31MQ063ZCJVbtON6AUxYTlDFgVIWu5A4z
Lblb9tCLzhkBMjrLZplFNZ8zIdMvXeHRADHamw1sQRw6doK5UHNAbJKZmLmr95GE
GRVyACC0JlMFAnWoaZ1Zz4/UJzwsHVQOBZaJAm47GzSsIeCM2JIl5/e1L/pJmU68
LnJUzl7neXE1UjuUXTaOQjX2XcekpsSr4s3Q0f2YjNaPIBGuRIXhrH0yrODFk01D
MbiK67299+9eUzolQlYtdIbaz481lP3m1ZFP+QsLC2U5JoU7Y0nDl/PaoX4tBLsR
LhlVgAc/OTQxxT/Ksqqtq4gDeC8TsKJ4T0T/ftRSzzq1yB7dQ0M/xa5W/b05ge09
XoLPyRjqqPs/UkGroQ/8QqJbRKwU8XMt27qfHO3S/lgPj1drerCTV04nK3akRxTU
cp6DmDbWie8v8B/mlBXVK5Mh4+lTUQglup19i4gPJWlmx/DuRIPqjU0xUoQrKNal
nHWMV0c6n617+oD1c77ywV4WCKOwNuW2NgO8W2+j+sTQkdXYkcD8mUiVqvHaVOO3
RVAlI914ZtF5Y2p6W1uYYTpRN+xXZ8tIVax+1BBdTV1vLlM93Id7CfaG08UQhgDN
k0IRe7jZIjR/IMYLZYfn5HlKnBUZJcvdq0ymZJVainw6ecJ6YfGi/HGBdTNQl8D5
AMAq97y3KcwUDoyuncvsJD7mwyNQO08/M1oRdZ12vPJRh+6bXectfZiPHfrz9JKM
ZgQXajK//vy6DnAkmUNrXKzmezJj7y370626HEhw+Rnupc2W5XkmrG+I6SRPLUdK
Ts2cPRm2eUbao/tm5TmH6Q1nP/O763fu7Hfs0884scjMLq5TUUhzOioPhqfuFuCg
QXdG1DW4qE3Fx5+Ue/HyXWp2E3cO9A66rftKYeW86UKZtuK/47shp5nE6yILOsVs
66SpfGQ/9XgPFo/ger82iUO6bmziFDfdYSkVPrg04bnwwDgdV3J4uXjfl7wQOTu1
b14/RpN70gq6Qh7zUdsyyDzvwX0OAPVr3xyNzSBKVMgOKQLrJBi0Fe1STk9jEMXf
ZyX0zlD6lUDryBVw9iR/h0kaPcnLtUHz8ns/y9Agid8PztbbHiPxdIprhGw4G9hR
85UiryFH4CEESwmbPHIVLW7YJ/1kw3Pk6dqmgvaCYetetUr2jcSMAVhmWZfGEugR
6mFBgBLxAeauKeS+ciInLtvSPQuk7iLOZFDo/i9U/Z70ffLWhcMWJZ0zOGkLHA2C
sIVb2L0WQ/T1HPY3Wd39j9MR90JX+vMNVo8TqBtKy8m5ikhPkRQ+NcUqEJ7hUJeL
K6H+uRgkmp0SpQn/edGUGLBaQm7xI345kP+Ksxpg7qQmzdjrwp0hPBzF9u9lxjhO
ZafpAkR2v2lA6DsWu4zHU6rg4sSl4RqhdFP1kurDpnRoGE4wCmXutWGXvF4vGu5a
05VmrVwWMJt/+AGtLbwBfqUb3FJaD9GLjjqBXI2fqb1NjcVkM3vUvTe3oPEKeiCx
ev2OChDOh1tOP4Pay2+/9kk3iresjoFb7d99D8kegtbs47flnnNsJyQDGlZAlipl
G2H/cZJvaJzxeb8Ev5yPulDS5j+PuBO254zmcQuevySicK434fvcwMA0qU28BuHq
YZFiIH2ACff1LwaUh7HcsOv/sGlgxFobclDhtsLhO1xF+bIARkvd9+1gUJpJqeWo
LMASei73QKX8elwJH2ku1MaVF2PmKAIbQL9jyp7+yoJuwSbR9wJ2N50HJsvEgLnQ
JDJEf4b/O/9HZh+kZb2MqNCvhLvLWszdoQE50bFMz2g+ob3NO68coqJtmIQcIHe5
QOfTdHdooyQXv0Ex6mvPvd/YtE8C2A46BscQ7UmezViWOY2LYFL1ej+z7Bo0P+er
xLtNA0pHLfn9OBd3Yrg5iC1S6BQQqViPSL02jVdsyWohY3S/aqrvpYT87ITI4NsX
xcqIjRUwYjn6kasydG/1562gJdxDXkJ0Ptm/8U7jBHHOkuZjeYlSseyVV712w90W
Dd90/mw5GNyEGLQNAXzYOBuHVs5flvxru9OpGxrAb7KCae4SIYPgMu3OrM7DDHeJ
FLF9/Fe3RT+5lYB/1+HtDvCJhE0y4m2iY9omO6mVL10GmYbSNh68MqXPtB4IuAkO
V9GcpmNO1ymlJt1Et2PmZWrtat5dSpiN3wKlHnnP5JzQR61z/z996YUWFFZZIDb9
KrgEt0KkjSB2kxfooYDX5ly3COyzJarKTfbQrpc5S3miruBQQfRWRkMd/5/0ZvvG
k9F2F1dKxc4zMlQiwUGLj6WL8V/HmphVs+OVp5f4bVvhpXPni625ZjCDLKfZl+XL
SyTIa9d6hJ/i6JFLB8BR4ySVAzLl2I6TP3uQqWvf2I1Q734T75RTCfMSG23vJPk0
7l7AtPHumdIqYoqJKfKA4tg/voDfj1bEwoU+de6HaT0XpPCyeajeFVY4iCepKkkB
qfp0p9pdis0FFIdm3UyzCX3/9oh/dRVNyjozirTIx4+TXObh3pOr8lSdiqVUU6+X
AIcd9XIp8XzxlU0gDNgHSPfaTsxUgYqfZxpzwFzuusSria6doWT9fV+a3t7xv/dv
QiohIPkdRbjANmITPuoehRRenU34dawlC5/OnygunaPtl/4eLmnxniq0s/fpmDuw
s/3DNDRuSCYdHwkIff5vJOaZLEhc9yyRJuUh5L3QPdLYp/XhlHhsmBdqB6uuh+v4
5CVWz6ip0pl7Mru+8t1m68YJycrcBRvxceHOAv0YeV8LEfPMiGdVlAsy2I9SOVuw
6kmfi8J1GrFizyujYBDE9ahSq8c7zPVpiqOQ8EtGnU4vt85TCHvU40XuQEsPG4Ap
mFZpR7GntpRjdGNXT99J9tdk+a7or6pDo44ByQKdjGBC3RR6m4Q0QkHLOSs4qdMH
MtlI4XrYiMvR4A2SMWNoscQnYXtAAsuoYV9iz7UngPkA6pOPTK47YblvkDitTdaJ
uAJ5oD2AerApXIpzVv9SshZE6rQZt2h3ygLJQJBqcRcZaWV5ESSouSzpXJkqm88u
tk1zGDnjfDjciykKSqZmDIrWAzGQUvp2jNb6lJYzzBpu1NB1Kxy1JhStbaj9MyzK
LNTn/Qb8hnmUn4/5+ABLVyfwnI2ApxEcT3yxqVksqK76ktU/tEaH8YzV1vQQwoBG
9Nsh2MXiKXu04kBV4xcnXPYnKAQqMdQngCNj46JOsDvld1ujqxu2/KvSzcgf2amF
lnRIZLytxdErvrx1Hvd46vjS8iNl6eEQfdez85+r3N7TuUp2TE2I5+N/D1IuYbfO
zYiLSnsmH589Bo6rNJTD2fxeKjwlO+3ndG7l6x3HS2SUQBIG/b1TYxQ2eK63Vxo2
oZaHj1GOnblqlA/+FIPzXv4ntu4kBZmVmCSskjdrDLQyPEIxeDFqNfVMS/Sx6+qJ
ZmwDBD1NyiWLHHy/EqGbYE/bow5W7i4KxlRNqKWA81ICZvtrpjfnSHriodoLVBux
WiDe/84x0ZJ3hSjGDEZ4Qx7XrpmbrRY6YMWxN3Fn7t/jfC3KJMJKXP0PCLXAm4NK
XvhWkLbpYeHDyrlSR3yH29UQTKdofyhrWOJ1yP+W0vG+wLaneAkRT3nTp9RqkrVf
go28pPOSeoe4+zGwZW8rEkfWTvzOyxaAyRgcJ2KY61MeqdsVhxhnjRVNBT5ILLCe
Y8Z2zEW68b1imLer3RRjp3rMmw1T8zcPLYR3HsHPydcmh0YB+fN9kz0tjCZa9Yur
6m6LAn2PcTq1Mk5muJ6JFWFmvEgsRpgkRievki+4A9kGRwYNtQTGZrbcd19+jMda
t7ORxkmXMrQA5KqsMr5ytxAzqLhzM/Nu5bgzhbK6Sw4fQfyjNHlQpH7kmXiEUGJB
/+vAMiH1ecy4nHTEJapn0IzSDhslO7cjCQpRg+2RYrBWRmaLMgSV5ryYK9X+IJ+4
4koWZ/clNrnV1Lqu+Hxz2LDz9iku3jHR4RkcB9Bh1WBguDqRXWD5XOtiItGXxmHJ
qgBwbCwVSYgpvq0yDNtgeld5diN5mRxjV7ga2QPRI2kBQ8nKPx7MFJQnRNubhOhs
G2nD/7E6jpd1gRyuzYSmFqMUwsk0iC0I348IhSpNGiA0dauq8elCLBRexZ+ej/Mx
+fkjA4LE+az8DrCGVjpZGyvhBrhAUPAq2RvtWe9qPBb8nQjnY1WHfhzVxqp8eCXE
jTCIi7G5DfzGQiZGCFwZkpNnQwxlIiyK0K+aHh/Alzo86kaNQxq8h2oLctmIRDj+
B0/cNIldgKo6sXg0ut44GoHpBOqbIXibT9qE0YviL9Tgm4DNU/8bJbuG1pGtO65n
UcON18RRtkE+LHs1Yy6B8Vrq4AGLwDuxQR0FQTO9hheKByviwRfIsHXms7RMqNid
NjyVdr+99hh6N2fOm5BzsFJAhvESPsGvGSI/BTAEkSAjcemnv+iMNn8O4I2lJ46Z
oIDs83pnZnreji++KdQ/NUinoxFHYpzebMoSRJjXRCXSKUCreil3M1JSeBtqeccO
2rA5ubzA80XWjU47I477Xw7P8KKfZf+lc9LsBycJLdid3ov9vRjxYvjxci+l+Fsb
FZ2VKdPXj6bdS7X/GP3wQvzhWoLzgTUE2jEGnpfCWAkRrYr14WGNvg7uuMrTBl2c
J6hoyWC38kgr2jG719DnmZ6ZzGEtBy+vpK1sTt9dPh+R5ytuFkwkbZq8cL4Z5gdN
+fLeMGNKQo/UMCiC9xJop/U2QqGB8cVzdtak3uOUDs2WfVAZZLGp8OmiF7EFcFFO
1ZburYkqzkKsKRMYQyxG8hN6kgYrcz/HQKl5eFIZ4WQc7y+urbmDX2jsI6Uv9cu4
0E+7Zv0HCRZcs7XJ6X7A7j1coVGsMJ9A3tOICssxoyIeFckXzAhzkB3H3VFLqx/L
r0w0pnSD+kMs7i0bIn+Z8C+oRB2k5m2vplnkjpBhSYtIV9n0B8lnyVl596620X4N
gxzXYK4RI30tBqqKpnJ4wG1wfRrW77v/k5XRtBs4+gCTgG6a9IXNL93PUzjwt6cN
uNyxyz5vJutg4HmwR7JoPRDXRzOPuQv4dde8RVwhUNKJk7gvB/iW1egMKCdzXkE2
cOch/GrHdMlLi5Ua7WuUT5LN/vREhq+k3wQOeenuQp7VHN8Wi/jREQo/1py7O+Mo
omojHtX1JV/RqJCp3jrRJoqzjJwna8IMOs6pIudDCYlilZ58ibtDyisKVo9UPr+z
b/s9FKwSC9LHVLyb4QA2TU0pmRVFg3wzfxs4mL5VAvetJ3N91iJR3z1FAmroE9Y5
iVGhRiqGR9I9Z+RQzLReoVG+EcWjlof/mi3Kge0Zg7i60MjVq9L4aiEGauziC5g9
/boTJ4fTzwuAFl9nZpJaSyOm0QF0UzAtd6hrSvAwgLUwSOwaZO9WntF44iOc9tu5
FgGMU7UjwZh8HcLGQfhFD+bF4iDNt9aIesSwhIzPoNDaZ/dirkBnWqmMXizk3veb
DBMz3XS4576xky9x0IRFokjNpaRVmOg0DIhWPn1fvZydeoGZFglwLxRygw/C9j9N
a3jViqR56aTnHdCrX4Y6NJ2dU0PNv1+gz+I3z5AROP3AOCG5rZH9z+FrO42UAEOm
Di1U8l5RhgWDxaIWFOW2LR+vdSfFlyW5PJlYWTpgW3DUDrJ4sNBg8WIbT7A99AZh
DviqJZ8sUHGRvkbUabzx5sPxYVE9FvAuLXvNrHkT93fSa2hzWm6uWKUw1Gr9ect7
8VmjcGnfYpMfrzMVyzE7Av4qwxRUyTDfqEsra/JEW7JkfYnamapF4M9TpEW1o//E
L0kkj35fAiO5rbDec1WS7B+qtPOUtFZeEhv3ydKhqz01LHaDoznVD3azkBtiq26W
RQkwAnJShjAK22qTjdEHST8Tks8i3pnROuO4Ybn7h7mtzGNMkkmpnAEiLLB77/F4
1CVTWjEV0OnDF7jlPh8P64pMjNL66rOpIBhLMpEhezrGnHh+kA2u7YmSb1mAHzhu
zeYb3Y+e+7n3AUGV30ZHAU6RQTLhtIXrSg62UTqSd25hV5Z5IePdQZjtrkhxy+j1
jReXtjQ4fBolXUHamqwsWIOEzaFzLn7Q/LQISBDlB+JWVnXB1iDFAvKW3h+9iA5D
e3RhRL3Tco2iktj8Ybs88xthEg57N5Y0SaRSKW49SPOOe4eVxaX0hNWUZBk5glbt
oKQ3ZyJ/447QrwNiZmBJmf78zfrivYTEUJJpi5pr6rrBoRBiv9rp1Rdraw8tgEDJ
Amh/BtUVZJJ7x7OWukK0rrVRbMqUnjIk96wI1pStyF6g2IawoAPjX29PFFk3UiJ1
TL2LjcoI+/b3HE4btyAfg2A9Wgm7vBofiStcPaoJl5IzLulQ2MCCFcdPVi2K/YNb
fVKHDUpiIiZMXdWdHTAobN04knX0kyRkTVfrl35KsYB4E7DOjcumzlvXeXYauk3E
3FmoqEBoAuLS1/O4zunvzyBDr2UR/gHVIRXAnc+iY6kouy3PuG3mx2N8OcocUvLp
/bpZZu3UhDlorLItgBzw3JhDeydqfBh+YKVxIMJcYDLJTBF+gPjB3kzCTSYXv8iV
KS+AxGdr67n3v945YwVoWhqZDEHdDOCkUuVebHfe0XWXOg7LXxTiD+exKoEmPD9F
5N2sLiuaifGW0kJxqz85YKrQFodFUlvxI+g0V+uxKr/Rr7NGaVeyECVXBZ1qBUFw
di2B12gtwkWaGJn557aaoQ6pDuB2wUMVgYyMjEVvfIWQe2Z6hcqZ3fqeu7iKcVUs
Lnwfmx3it/ywvAoRgmzDfTUno2QJGeCw5LxkvI7zY81oD8tg1nhn8tg07YScBjHR
tnWOTl0oX3BOcHooq3UmQz6G/2eJKAZwg4EBiykfv1ueFO4mGbFp6pe0cjTr4fzb
+G1reXFUM02J3qi+eBhbVn9Si7FR+shDRo+PJyg4HyDFkHmBBtDL7KOxhjaWdrKY
iYMH3xiJ2f5VmJkJfe35zbEUz6Z8s4mMmFbMUCfvR8vXj1IC+Pi5orsbgXHffVsX
CiQz8+thQrBu6bEWO3+khMKcXsOKBXHzk3aVLKYpVIpEVrmmUEdjXG/nQ/drAuoo
iswX9lF0aLmU/JvCRdAtDfr2VhSaHuCjoXeVxpsTxkmWVU4u+lU23gh5HAJ9HPpR
ixVmh3TU0DKh8jqESLVSU6IlKRlFAuutkVCsOP4+b5HeVI6b4RDmMrnHSDR0m6Lo
VlZWJLmnEliE6AOaAa7ad3GswQBj6HBp8br2u5mHDI6l3BxaBxg7zAEZu0Qnlnbl
2aGcrjbmQpsW4Poj9GzvXsBdkUIk+YE4fBzvfxglY3Ci6D1ZkdkAHn9wDQ9/62CG
YWT8aZmE+01RGNPL4Uj9hNQBLL5n9U6q6cfQ+c9X2EBexdYVSW81lXptuMXIjchg
GXsw5YVUz09GL0XaIkabbNA/2nTwEbNKxJ+uqhQm+ZRypNj95okfhFFG/lUs7fgN
6Ud93bqUrcyXlw7H91umh/hXFkV5xR4lU/mMFoHf7loiMOS8QvmIUR/UQDQV0Mck
OX1vAyBH2VRXjqYxYxrTS0LX5eFUGAd/RgUygTWwSJkgD8U7ppDi5d+ObLXSb4MR
PgY4hcMAHnA9cxaJ5xYdV/GCghtydoQDVmQQmqHYQrlfNLRVjhwVMXXhqJ7nxSqm
bQh5x/kibV+Xwap1HJCbKS3VdtRnmW+hNHvCGPCM9Ke2icsOUaN4yS1lx6NvyHXx
O4YM+NiUfLLE20p0h7cPi7V9FuXYD6oa3SYLQoDteyPiZpS7mk8lE5xLYEuvC3/r
9Wl0NJ4pEPsJdKbEABQQWF1YrHPQsHt3UJzvAb9YhT3NN/HXZVG0XfBAIMNnAbh8
vMAWsPemDGdd1jcoFime65pX65xm/pSmQBFy0wyJL/hIAQT40GchdugnzbR/Jib8
wmWzCNdOIr4wsh/kYuA+KVfeoTD9l9Wx0ftmLt31GnkniGElTR3tkpifOvX+rdMT
KSjTf7qI3TJniKD9DosWx+eK7dFQVtx/hk/IYtpeBGbwsgd0Emixmgrl/KtV8vaa
Tfby2XdDSUZX1+AVi5f+XaCUUZSTUhpc7ZZ+kfrT3hBEBPmX8fSCC83jUt7yo223
Mi3d4C9o5yiV5Ivc+bZmxbsiY0p3N+ObkvQQ7xwk1M6ncR/rIkVZ373t+jpqkrkg
kSJvCnImokHmALhETRGKGw1pUpCkpCl77H2p2TLHOGbrGOLxktSXqOqbxDXIjXMq
niUXQxCheqrfFB+ZY5YgP6lrWliu5JlG0KxwjmNPF3iyZbDn5ewXhwvsLxyq86wG
QPzmYK8HcTNKREAUFPvkx0d8WzAbGUnck2lW/wQexnUwhrAByZoazydIK9BkPDtR
En2StODflcGiKfseVPaLEwD15cr8aPmdVgLAdfKGy1sLSvp8YEN5OqLn0bGTqOMj
+79d8r0SxLAr3LBcfCq0mMg+2VpC/eTAWCL5gbNVWVS/DGg7JCtnr8vKWg6kis0D
OFlkChbaATSYuQLCP8SAFGXarxz8YQvYXcRy1Ofna5dS7xb6/y4UA9pd56mSWn+S
b5egbwd9Bq4P0xKb/dQTGI1v8M0PbjOu4f+Nv76MxoMZDHTu9IR23x11lAfnnz5x
FDACNUTxBkQqLQTDdz9LErtVOU65pUes6k0h9ozjvUrXgT0HzsIrseycAHqFiyUR
ryNq/Fi4JqIK+XYkm7OYneazuJ+SlttIp32d3UKvPy7msKv1o/Q/2FF23rfmRceL
wAmle6LmFqaU3qF8UahiO7S+icl9/wRYCOrmn/euvHm4WGxBaQPHxJvpyFE1+C3H
hg0ZkXan0DICfBwcax+D09M8coppAlt/kkkJEi7PHFJ1kXexGhnRJhsNanXr79q3
RnMaBxRfwjBg6adjwXeLl9yy58Ae5i+hB63SOv3i/XvHaZwm1+d3dDO8szGDI6ay
f02Yg82VYvOLIBPjpFZ5bwdbXm5nDkBbzEtWC2tfJtWkW/QjBYYS6I1X43/BQnf8
SW9vu8imjjRThJO/6hWdWWID+XdYBkGDGGcchdFa1toi5AlgVZRqE7b3xjAxaEOf
Px3D7J+z5clben7zcW9l82EHsD730HFuBLMCHOCbbNJQ/w7PmL3Bawq6MGb6U17c
0FJMcSHpOQmvBENDLgU5oqPgWF5Vjr0skycFLufKLJA5+gcA/8tDi/cI5/xSRA5K
rjk6p7RXSiGKAMm1OupgCvFcNtM6L7+o3kWZuxNNXUlPTNTkuz7tHUqPGdbgUIum
iiBGU3Hg0YdM2pE0Pi1HqvNe0NDCjlH1EFPQS/6xZgc3B5ovN0SF8usJ0b2J7xiM
vEV377+eiqtpLperqQOw5z4Mt7AFXVDIUZCgRzz6jeyuA4kexcnR5gVf2CmjAYAm
SIqurxRlrcEXF+7t/0p4Ys4cWY2MjSY7N9d81EvqAyEoxNRN9MJejMDjp6RR9h5H
9FWmj+Yzq0qfMSj5FGz2amBTc9snxzwX1T09Wrw3Q02xS1xBTI1mxZWjjiP8VATQ
3an+07/ahMQ/7YIJnHtAbeal9mpod6LPIJ/WCYeLYDTL1T8A5FiKAifx2QCVYAqv
WG0OACtql5Lb7y7cXiSRovEDvnw4XpR6lQMtNeNwn5w8M1sdDOCG9cDv92azdXdO
eenm+0oj78yyNaoDvJ0+xHdC5PpJ0Soih/0QsVG26BQrno5E4nevmEvcVfbEbVkc
s4l3YOlkOgutS3Upm/QKzNm3dVygnlGAAKdpQgWl7c3OF999b37uUJ59NaidQl67
vNN8Kr2GJC2UEdyV82VWBMzN31w/nheLNSdelW/NylJ0BSwTggXYLDUXzD5lw0nH
9aWb9G+gcIrpnwTZvNeecApiLy5F8br4JuclK4Xl4r6WiLuGAkpI31vQclMJkB80
uuEeyQj/8khBpcIEvAquF9eBsQXT93ZAVrQmF8citDctpAXFzlFfpRci3alst1gd
0GVnab8YSfBjyALo9xflyRlFfcMYAtv2/qGUdH2HZphxUR2PijPGYqvMqik3tqw1
mNmeQtfx9cdVrSj6luGKv4XQZoE/EqWDHOUPn5+xHJ5TfGlzm/fIczxfynD3j0B9
mDwq/CEOZfmH47Z0p84uQngXT4BUYRSPbU3ygrO+qKv5MzuZv4C1+itERoYzbYI1
4C2afCShKl7Lrt6lYtG3j9XNUoyBzPD8A0sm+G/lWvtYYieMb0A6y1UbHzMAkx/4
WoEVgIeLAvDctcPwtTYXQPPeLcCJGQoED1QkKqgvye5141Ze4UJb9TrB/SJ0ztPw
8oW0j5sDYh3xryt1sZngpcaPq/aSQKHM/ku0A66jWeOu6oRQ/SYv58DnQKzIQY98
DsbRfnwOmI9ZuPnhb/RImSTVha/rCvWVwIm98TCPsZc6TyS0dDpIqG9zDanIf8cQ
HPq8W0WthNSHkwYSQXiQavGnzJk3CVC0IieMjMR7JQaPKimkly0m10hF9uMiI8Zj
6fOcyEvdrsPf4P93Mk5VS1wmbFTcy+nBn4NWn5qxwOduzG7LV8+1E6rxZ2lxAU0e
UAmgzUPPSIJQToE5/3wchMU3Ig36N0UF0F0NJ2c5XT+WqYFoMY1bTPku36+4b26j
lS1QCAvJiuVoF6ix7ilA9TpCbKSq6JYXrGCX4tVuNwlxU1ZdeaWW5PAj456l8ZlT
MkLuEoP5T++J0ihO1txlR3pOxf8dxODpNlR9ftqFyPeWARUegV/6YtCx3psfuHU2
PUD6iZSUguGKskMbOttSppXNnHE8+UOgZm/ryV7+igTTie59hIzXzYW1LDH2LNiI
qGgNA5PntoI7TSXV6OolroOCpTL/3ec/T2kHYvSmEKLOUElB8dM9cFOP9ghQjFuc
mLUBEHk97yd5aQqv/k2iLz8tSdfbV5J0GhIb+HX5HVDh3HkHE4gh13U2dzau16K6
gd324s+55fteRyWgmrQFOSxkWJ1HNpEB4HJrdIDP/FmjlC58bcfwSzyzxUCQ09ir
MkVM8KRGTx4NH1Ei9a7yZKWEvOnhUqgvtvdfjzz0xOxTTSO/dQH4ZvWcf9fRy1BK
SawMif1u2SfysGqRR55KDWhWPleR3pULglLIvxx4rUZdDdtSw7mZGbZ309ZsOhX1
SON0MdxMHGp8XfpHiG/8iYWfKQtoUA8kWdBBX0YKWJ8daJQBbYC4GJK7DoUiKjYB
J5PtElTcd56MwqhzBzjbW7m0/sCmUi7FBtXvN62Nu4y5lGI1yGH/DQ+LiX5vqCwx
bhGxE0JXWfacNv8sh6+WPv8Fe8oKgbEC2zywgarO7xNw0wi9d3WDl9BuYVHsmjk3
4OWcZbGT/VtORSmhL0wtWYoDkTqeGvS8c0IbOSoSR+R/o+z1cpsXtUSokzbwwAyg
4qC88hY+nw6pDTGN273elsmhvKemgle0Kwu1xGLHaSaHaYSzisT2Ge5vFP9GJlnU
0faKwinsPkoOGYZ+XWifzzIkLc5EzwGNxOzDpYzv2sAHj4O6RI/64VRiwS9FyyZM
hqyPleVlHO0nLaL+SYBkuwk1DT6ndw51f1qFlDPF155CqLD9Lrc2jNYc/pg9b8yL
yn0WEdRE8B0UrUhl6Hjv+tVPfSrUCmnmLf8huhA3Z71pRBESvFsX6e2WlEUxLXPz
zG6mf5vWZuJyYoHVF+s0K2vXfVAHseluz4hlYu0x3y8VOWqzTr/oLmF8Omj4qxL8
6eGvNyO5HcFOpU6TCFKx/D+oxN18gK9ajgpIgJ/ChKL97bOdvAMEiEb/iNvAsWiQ
V8/pdcGuXepSFxNEA6kSKv2YbsAcjY4PpF+F3vK0nZ142vi/mN/TaMXLhcmbIAc9
gZTlwyJNBJNeHhfRPgBR+nWUd5OSzGLMkSlvJ1Q9K4d5lcfs27lZBSmguOZKwiq/
VzobOlLIngfJ/z7zuraULhuvm6pepUIIW3ViDJ5b2tCjI+ryPF495qyW2eogovj/
e0Z/4bW9wicS1pg9AZLbB0ggOLnQ99TlKsFbqla/15ejZ4biCr1j+AbI3Y8oQq98
2SdxUCY1BSaaDwBfyFZe0gVR8OYsoDeJtuM1hodTc03o1kcJj/TpyjRBKmtJPWHN
tsHFt3figFmUPO/ugh7Lt2drFxy5lN+0RgPWLCbS51l9lDeuzOjg4LrK5T95IJpw
8ZRflMR3ucIJdT9B2l4jh7sWMmN/Y/tAYORVqWp5Hzd3eDYkStBBt6NOs73HSwat
kEcWp6932p3713+znjDlFFo00CAmOhMyOo0+9FJKjZdM2k78K2FMas9bO+9hx8a2
77jLRF6105dnIj4GAOUaoDQQQaDkZDLkvf941d12f1pwZqP1mPISlSnTxkiWfbiU
OzJOb6B+FWvW6Ix5YsMZZREv8icaodAr5RHJCKFiJOK45ut1Y0ztXAvPwYHxn4Qy
igxdcEMAza6FDYkAFshH0K0YwM/2EM9SJNfBoJPQwC9X1EQX7jW4Pm/oDaOc8uHg
/23mMORueLbkADbXdS73GkJDw6E+awwzMrttkW0O4RP8DdWA3AmIYetGJDxRI//A
WoH5YgPsiRSLYPOfJT/h+ICQRFqRDUL1QBbEFpnQNa5R7t+biujP/bHY14ju45zS
Fg5FYOu4JU16rTWw429kGGnWwpvXgcVOll/UwrEt15LVo7jnkAiFgU9Hu5qnKnn6
DDFJVkxcjJMEXhMG2gTFSj5i04LFwSjGQ/zI4wowMIT09wCHMJz2vuD2WGNeUCfy
GT4RTFhpTne5Tx34K7n6pZ9+hhlwPhoT/5pPhJayTFM4dORvapqtet5MCAdEO/4/
mWTe5YDtGAMbHKXvZ+rqh17+qhHJC1jrkqnYDsfAI94mHBmtlF/QPsi0A52n9k0s
9bjLX+OAIPOUsZAi61tbcSfmI5M5uLnWXA4J2quOY5vI50k19ThprN47BoMJ059i
4Xh0gqp5JAC3IOdn8d07pJvr92d1YLrayW2OXj8fUAfKVsPn83G3sQXBefdfO9pR
xZ6YIrYLFdJ9AsnKeXZScylyftlOjQFt2wKPglafgZfX9/1utl4QX9k2x26gsDdf
MV/QrGV/sx2GWCBJr9547cuPsgihsljDBFzt/LcPC/l7FpvSoUOLIfJuq8LEd7NQ
DGfxQ01TJDEZ5c+cWD/KsPMKJ5ci2AitkSnxpbsh2ZtCu4vVBB4m/7KEhiN1PuDo
1Kli9CV/5CAZrc5nbXAsOg+0dMMMrmoYeXPuQIXJjgZ/p+7VbqkEZj4I4cB2zAUm
4rfFFJ7AaGCLDMR/2iZzIHN54vhf1lXEP/9lskxix4sf6/uv+zBKZLhAs6UlBcqq
q707n2JvtmraI3gnzrSWh/NceEoQtW0bi8BfPv/ojs96PfR2UWzICfzNmNBpA05u
OeSRasla5psBaFcx8dChjmJNu0kXzytPMZfwyE2zOdnQVnaaOvf6sXMlIEjdcAiT
CEjycFwt8VxdPXLItsC/YbBmzM7mw1U10RBNDaml/3FEHXI8XOrGYtKhamET8aY1
J2bVlUkAVrYQwSKa20VaUUpf4GFuEQi6lV6A7y3UkT8ChiRPLDwbBZdLiSFth+PU
byyG6KN6LI5hN63eYzH5B1EkjNFoC2gWIZvJG+igzF/R7jnUFM7eX4nG66Qjj0T6
AYEdX1PFHiXzAy2WAM4AQNpLyS550HIwfHtusVB6hTuu6mH22biLCJoe91ldNzJw
m9uJ+6uKdCQlWfidJHssMVEhqJDicdtQgqpI2PMlfXFXk9Yd78euKTYYa1CvsW5N
8yWuQ/9wvlguD7aLh8QPDJmbd/pgFkgY7B1fFK7YT+SGCKGajQIiDiyE6ZphqQPG
tfZIgDfpeVZABWpK+GfKFbv/+d8217iybhBPcfklddP8msxDKrS38GimzrXPEL1u
WlXXCHJb4oUG+YpxRar1wum7qr3di6bxG6ghpBsdBbxf5809XNCO5SO7NwiB9VOx
bKkfQpr9pIsi8FF+HlwvUq8XcuuPBvf33aKxcSFfNo6bFdd4qybLzXN1UGj3z8/W
zpwd7bUJw5cRT39txT9FmMGxQ2fs8QrmFBaiMxVeZutQkHDdGudFnTzNKy8YqYm+
tQTULfh9lXpS+fM7HR1leD+B0hC1fhTOYTwzJyGGNMDko7AskCh9I4RKMJbV4/gG
RgHFwY5FolBYdOcezCuhqhPx1mgWA8ckVERMjPFff3F9OYd4DtCFD0Ghy7Rl47FC
0DPqBmpkiP2ficDjQ3e+dohDsyqT91O0R2IXbvRi35yq4A5iGX/XIh9sxuKsCPls
eqZWn3/6JbuXDpm/KsZ+GhGYmcNWahaRFlNiLT1hI0miggtmPg0oZEHumKrQM4Er
5qLB4PDFXdJYRAO9U1A8hr1/MtKGi3L1vUngBQISV810P0Ea/378xelVoBtwWe0z
7p/rD0Kg6y7sidT/yiwmTUsJQjxn/TujLZVAJK1aMZhwCf0102TkF3n7kRlPAqcP
MkVJQ2JHOI9w2euhyWb5KJto74sAoQonsDBiHJgW4MioHJW1rGgTpSfIsA7eEOxr
bmdPEI8jkDfZtKFCxjWq0C/aAPjjechIIwckjwS9Tu3O0Wa/5DGDRqjd2BgHMxno
wcwUTbq2c7c4cZGH7km2v0ra2iuFu7hYUSpbBHM5IvW0wn1/lTBqpT0DrHwbO/4N
wGHho1UdaNj1IbaXzibOaYQPE7CuJt2742IEKId5GYDYemJdJ3eKhCS8NCasTPiY
0FnW2kHoDb3PXfCgnU4I7TRrvljeHEZ0+6EygbttTcQck+65bfHk/2mcwm6UehAp
APhzzOQkokES+5MoOTprsebt4PQuNVrHRvC5B7HDpofEX07NroeHi37DiwTUQRTf
DSGuLpIeTHg1dp2+n6eIkKW2WHR2zGbX/2z6SL18p+W21S8oX6l44sh4flRfZqw+
MfbkVRhvpjVPRRvxUxEqtjLU2olqd0YFnGHBNafPo5rT10r5z2GP0aJAqf6x48fm
8htlFGcH9PzP7poMjaefkvr6xwllo3rMbaS0siX/061kOdqomQCgM1lYsJ6O5Biz
VigseSYMDPZLS/wzZ8l4t87FNRWZbrCgyLyDiOOTkYTWNc0BRxYu4bkSWZUqHU9m
eEh88TwBQst6bsXb8itJWcRWaq0ucUME48O2x8o6oHYt0XrMtQJlz8TQh6YIbBYm
fsIzYC6afTdxossCHfX06wCnlwR459aLk/1rBF9O/mTSQPz5lYgiOCnWDO63OdHe
+Qy2ZcfsiCLRC5i5DPmcNxlsVOsleCRCblAEsaqMoPIgq08Aq1KmiV+U5DZLuUfm
W73lGso4ukOVRwiA4IUpEVIfnQA7/inTnVXJwF0KGqlY2HgO3xQcq/0Fc/MEhApE
yy0S7+DsRZBJLNEOvG4IKUkDNkCsLUezhuLWwg78xu2W1DfFS+5wSXzT32Xq9841
pZ27uq4SmCiIA1CLnwgTnthNsAo4/vhmlKJjWYPGO+jLOik9iftfJI0ezQImZa5R
zl7kAHP4R4v5xME7PAodBa2VTesWMMYgwooH5M2eqWlsH1DApY3ejyDeZ60NgFGP
QEQ2O8PlAeqS3U55eeiRDUlb0L4AJe1KrSwfFXFxoRNyzqQ6ehSectDwJqJ4Qx9O
Rjlq8fxj7zC8fg55onIqENMmG2NWihBq7mkAOdRBiNl/4NA/FnnY8gSaXf3agsr2
qbIo/3k+GfccyNKgkNUymnDXGCOPJhWkBjSOUxvjSDVR6KZ3sRIPcA4/mYqRXiWW
YLDfIdeHp2sv6gPHUVt4ctQ1kCLwfPBvcotrtCi3ceNRKyJbViy8e+qcRjnF3BLB
h0BSV0zmtpKeFKJbtGztnMUfWRIEqZAPiwA36IQmhG/2jAhIW1VXz2bj7OcoVF7P
/3VgMX9B4cPeDZyHBtWHpGm4sqQTRHzcku1x/l5DzWER9za57i8SGnwt3zw/TKfy
8Wki7N7uiDACzX5lfKw8S66Gb+aj1tmCENbnm3rvqHxLdu2YDwNAY3i+1yFtu12/
uASK1gjKuAyEVF/E4QjO+EV5vVYxcYZciO4ps5erQTcU2bje8sfe7Kecsj0PxqiJ
zizP1E+jQHQTDITkJ4vXYvPbyfzSzluxRKaip21qTkhk10eMPMNwHU24W2MaWn+L
nuUrG+rkMVhsiiHWL4L7X1juLFZnjtS+tl0nDxRod0dl2aT4QZPECVMMwN1b4wyR
FHkxK6OYfFLXPtp4F5/f6W8kJa/yrrgwn9rbZkvM4oxAGQ4f8rPsqgIkT3h6GrrS
l0um3/F5X9wQcLJdoaHSA3Fv3EkCHmAAjAzhD5+LeV1B77Nk1k6GSmxX9Mfvk20c
7CyOKkoSY6wyW6/bZk3UhrFR1sDKV04zxNZC2Zex80Hy2peqBjb+OIjcNSYNDFGg
PwKKPaEKI+K3rtGQ30y/HNrRy4cOhssMYv5I8AExw5hIUINJsx9DOTKxN/usnRce
x6EbsF40gXPVsUbjGbcO/EzC4t/HRoCMdnQNFLJ/NOpylvJsVmjWmR1uhtmjpSnh
vGQqBBnUofs93Q7dh+8xT5gKCKNb9wEfeN1Uhh2FLkwFIxOQzVwN8FsVKo13aMCN
ka87EPNWaDNvJEcu5Xhukk1Yxxuce1K1bNlGIfB/Bz78KkJUiLAMaema3LgcHNdj
EHPYWsgXAJmh9HYZ2P8Wf6DI/Sjvhmg+PtSqJssT3rU28deY1NP+uj6cN77Rr8TZ
qkTlF1s5/qtC11DHVv6eazPBgXxUuAFTCVngaBZLX5XbhJFIo2E5CqYsyOVlOu4v
p8EzID04YEImWQt1KO0EiBFkofFSAExbgC/3DuVKbKs1sfaekKosOS3D3iz/0sR6
rsl1309gjCETNzxVx2MCUaUpUZXt+zr6IWDEbU7H9hTleqiEtGkr7Yy9IiIug9zB
D+ckNbOcc4lwE6pPu1cMQ9JZcuJV/LKjbR+tWDWyffgHVIMXefk9HkMbkk8JgNJ2
hPUo9gQS9b/pxtXTWY/tOJOyoFEUVaTgr5PcDrZsx7UR5NPoH3BiN6m9LVHefNgl
3c/ZYAZC79o939rYgZWhUgwGKeV8Z4F9OUa5i+jVvX9DnVGPQu6u/bkt08cJX6Dt
QcYhIRTpXrg73m3j66v2ahWUQ1Qc1Rh9YnlgHinYamGRhXYxwi15rlLz9/NfPl5L
HjQESlfqF/uIMVsnSRd2D1sxZVsaPEpbObhc22DMYUaooOT3bnUEOmPdMLOYL3l7
E9qVLj8+KecaEgOtYmsAhUW9zevgM4bT5+9lWjGQeFJrofTo3Y2c44dX1Ctfo5RX
4Gx9BsxpC7Fp1vYGhfiARC+fdahQXmUlC9hEJRnKvU6lCCM1tDs1ci2N5vkf6ubH
L3qlhGOUUSHoVqtIWyTgY4eunBKTPMMydBI25EH5sz9xRPx9dOs0wysqa1ZyLvu2
nLiy9ct/vAoQCkVTJ2DaiTK6+e4xKIB7g0msKdD+//Z3qOeB+TsUFOi2dkjx67MV
5TuIvZ5QLQZlCVxQmZjolL99mDzqzEwGRawqCPfCFrGcsGmWPejh5qD/i4TpQyGs
SyaDOiKAtGVC0t/fQrr1lXon2Ql0XZUn8SLA15UGS2pS+5j6lrpBCzyEgHX1P6PH
MS/vuI2yrp40GsaJHKuXuT8Ef9bcfXfM+F3cd7MaKExKlm62M10OqIY/gdg34X1n
vfa6ytpz1hcUgaYL6C8G5/V1SmwkBb9nZ6N1kFMA90ffyRVBtPpmpmZ/3zkYlTAP
Nw/V6jhaIu+ZLv8bBOBN2Rw80XaP0WL7vS30i/o8PaDuDmV0yaJEpaRZm9GPRl/A
PHhbAz9BnRvN190F/TT8rmc/kJi/hchJ+m9IHe2WrJyFKqXBflQIFiLc5ON2H6Mk
tTvWdYUICdoQEBkJIzJ3yND9G2ph0mEbhtcNEhEW4Iez74B+/gKeyCJvE8sBi2+L
+/kwGfJTHDPc17AUiRtOZx7a2eEfijfQcwBkeTfvLJCU8NP9MElVFO3MMBTDyzwQ
kzrT1k62WvtTlc6Ftxjl1xdK7Q0EuG0CjmBkh+bjgXJg2ufpF+kfW/D3TMgv1sC1
bTMJMvPZEugmMexGiucnMryumCu0ZBPUr8eWqwrz2GPDwX49SiZNpx0RIKo8rf6h
LV+hjr1N6eZOdj8QRlgm5FLG1NBFLm669YORoHodbfJ4/mPhA1668KRGk2Rigdym
oo/6rmjO7FMV6TbyAJ3pdv7fWh1tngkoiQMReo44u50e2PMUgelmSFiVNFCKq5fk
jACn5MO/LO6FbIbF0SEmTA9Xe/jLVFs63xXWsnHs8CZ0rIaVfugHSCjoz6H8Eajz
CqMIDF8aqNWfnwBL8bncFXkOeLzsqmvZzuy8J6zQuLoGUwXdY7eVULC6iyd2Or+J
wWLW2kcFHyoFLGeuquZs/FurTVZXN8QDjWXV3bdHK5U55Cir+AeiWTErijFHnqFz
u7rUvjMQKAA+AnwyJroiUpcHqVWVjr2yuttm2P2qt/O2BZHwMyy0Z/XyWLlbqolp
Wd71ebl7Zwb3ECh9yyao7qJBO2D5zcf5vBjSk+5DCoBkg06SgAE/kuWHWCark3UH
CdJk92YveGacvD0oXGc3MHOi/dZQScHEzW76kmz4URBmochkb5C02gNEL8q3Woes
VDvcO72H9Eoq7DiXMgDZ+Jt1P0eR+EzPGy3/p9bonrjdPOoMhNYuhUdxmDpBzEXu
iG/fAyU8OEC8qqJMpEmo8tFeFIVKCDCWP3nZmEgP78x8WNrUSl9u6v63dSg7X8xG
BZe6GCBpfhLNax09l5Si1fggLbtM4IL0tqd1ilnBinb8Z91LST3//xfGC/3t0mcG
AwC0Rh3qJANrNmGyS5S2xyeRtOvTwnbBMAwn0PcWA4s/viXsnfR+9Ma3dIbqI6Ko
WXTr0haLTKP+FiIMOL/gPK1kq+tEz5HcYM8KgXeG1NebprMhqgHW+4I3d15SgIal
69bRq4Z1O2OyVPfKeSomQSZfU52VRWGovZIfI+9BEy/IcKyPP+x1lSVbFTSrNKuT
3u664TP8dOAlzszArPFUdialC7BeG/5Q8e9hYR1FjCKuBql4TjHFtTJek9g7LdAR
skUzR78iiwHK28wTYVtm5XgbaveF/lZxtPrf0D7/W2YPhKtF8PYhrj+vKn03hFvI
XT7LPCcp9HSvqKUfWR3ecDqMaAYKKn8/FZlaKTf4oNzxg7jbeJFPUEIVJE6W13VO
ve0rOIxzrPKqbvYHxQ1huk/c+IvqgL6TWx57gNoPc5jOiEeWVWWVM3leTHjqbLbK
f7quvE8sWo+ECFAeMCVL7WzdFUSE9DXB6HXGJYE/FvdOUWBQIhoB2ve0TF3AIXi/
qv+UT5K7v+phv1B0miejRD9Pd1mw6RrXl8+Zl32o/hGf0FaqIs6cMotnKUQlMpW/
Ty27RyEVaUh2FIml5aTjC5FmHTjwv4OiGNjd93bvXjMYKScnrxsGYN6Bht3JUam7
OpEchBnCwpUvyMFrcUUaiWjMQSQaFONTvbv5wqlr26Cebwds2j45fY8BbaVOgr4C
BVVCy4QHxb+nJZPBswr6DsU5BTkLy33Md2w1dKnBNimmjH5GLE1zhPHYKtjhcwGu
ng29KuqYpwBuOQmceSsTdlz12nl5TnSN6QW7XRWsrAa8mzP7OcBvC5eRUKBUkW+h
wqZPp+aPAwGxZ5EM27ATnwfa6G+QTUUsFnJPmuVvOKod7Ik5sYsICtRL58HPjsSi
pT4LVIhd0VoqCurCNL5yS6WCz6cmf5iY7v3aXGxeDXdfaJQDXFRNR/m5DhoPsHDm
U6n1QsVEyf/f5i8HCjRM+lE8WcEZ8G3rlguioAbaAJMvuLHnN0ugxn3Rq/hsTScY
cmJ7AEMAFyJdzu9EKzuZXnkTFKOC0t7A2cWnsYjjzM5ffTA5RxovzxxZnzqfnuqE
+k0XNLOEiawXVijqbt1V334Iu1C6oOSzTmkJWV7mbsft3uzawzZcyag7zc25opxB
oHqpkBjW5baQkjBEIlIPfrTNecuHrfQE7yHoPHhuyyV2hznt5U396ycqo8ktPZr+
oHMXqGGMase9WHvtXLnq1ZSQEGV/EbIADZBRXelqJ5c8+JBO0Xn0cMb7MeLxIMHb
ZDKzDnndpx/2fu8kLtJgnQYcWChD8Ru/qKFAlgpVPT6tb3KZu64/UrBNDcHluSL1
vEs47ue2E+jKb6qabKsclFWyOvkq2fHhBsAEue0r+p1n0/jxOb3QRRupDicZRkxy
u1F+eqJJKmpfIfhuaV/NbgpOcyx7Ns+oIjKhHOEz7FTLmC85agX2khMwXO3oosuV
KuYsK0W/zCkAmnzq4cAdhTUDLCIOd+Yr9924EsHUZuTr+VpTt/iMEb0ppWKKTOtx
rZMa2UESIHcmSew4HblYsHXsPsSR+39bfRhSouxmMq0Fi631JHCF50HmZ62oyJAg
cXIsiCjQK/ZW7RfzGC3+6jz80jey0i4fGwZpKDBlTyvDxR8jQFRBfDspfLoUyvyJ
4yf5jhd6hmqHoRItGuLvMb6VxnG3L4wl8PnMyhNJr/wNnr+CV6eF8MeH1yKSONvw
BFhr+r2GCOWBWI3e/ahdEn2PkOqx0sZ7sMcUHxm9U7aX3ZzjIYJfP+jBKFUpFQrb
DZVnWb/KpBrloifE8u/xkvyeEFxiaVYEWP1o8bC0C/qVbigLVKKF5GhI7wh6u8+6
se8JFI1WIHr2BrQ9IJhiYyAQnHOB3QvbVVJpNCNLjLPu7E9z3UWJMaPOY7eS2jzi
dmGxUfc2A0tDHBU5diW9utjcwSZnFL90I7GCbMECSpqT4eDK0QvQcKwIdBEAXxnN
HQQ+HUhbt0jAqeJ3+feNNmbi/931O9fsKSxx496TPauBpRlPhLWkK3kRU+fgVYsM
07W0BhyCWr/yr2T7Z5MKJxYdxfiIJRYxfhF7iWsjfA65udWHLL2vvieXGZ7EnvMg
sBrPRQuKp/mmDbTUyxYMc64BA8o0VIBlw4cg9/UGYsAMlopj9ewc/Hm2YYLH/k9w
9YxtuMLiuxjAY6z7gxuFIUu0YVyvobbCKRLQKF8Uj9A7NxAMedBgnCy0Siy0Jn44
TvBJw6oAVyZchfF1eXjzkbhOlSOuoZ0fRuUzQG65tf/jMu5YFoMuaJ9Z9UUzh20o
5z7p8Qi20jsCRFO1SeMacJjuETvPA5EBuFPEtK5CPJAxfAET18qNgAdpB/iMAoVo
GKk6C+PnhgbHHTrwvTZYZ+S3pgopBGEzAYXrezqoiRZQ9wZDNGXVAQUWukFDrTmB
U193nF5g//TJEmeFWKP0EZ45wUmK85G40c29t2MtE+ZEnPTvaGFp6etSUsFZogAz
kLM/SUssAxyYauufKgSzmBDoo6prGSIxD/c0O5tMTOzcM+TK+uLXVZVM28TFF922
RvPrioJmu19vkBBQxklpNum0vpykueUSf44SGe/KNN0s/d6BwU2ftKQComqcuKWI
3aBFkBy06Gu9CaP2Pzmd+7jkN2u64uYSjP/mOzG4hMbsFLkAexcv3qRbIx+aZ3ql
ZFWSM0RxJn6vh1iHGBsd69Z+lFMsMLyluy8xb2gcUsNPHFEOOuRAu0xXwD8/fVGk
4fwA8TBJVfvQ3fsnzOL0HesjcVDAMZEjFl6RC+LATOcRa+thyYznMIrOrS7YbDoY
9WhsvJFsgLU/73YF4dP3TJXgGIdgyEP8g3itWQ2GeJ97U8ea/0VU6xnq6ojcxshy
QeaYOMqlgd+AEh3ONWXzcS2JpY69Ag6phsBigS2QyQxtF13i0Gko32ThzGgGKN0V
v/eifE8tekh10osUA0pQp1E3ZavNzToIi+0eLxu8HpMGdp2giqU10gmndhYBF76+
VznXwjjZZQ0mj7eKTjRUZMvBXplHfwf31W9KOxu+g+7foptL+z2+wxTsLxq2+iCL
OyQrrUjyT9SABroK7VoxCYqgBq/CkSzna2KKSrskm8GRParYWdv0O+PTKwGnKA40
q6g8UzC1TYjF8rmKHgWmPBBzYkHxXYq292yQmVBOw8zbwlj/nZrw8LsDN75rJqY9
WF2yyg8+SMRhHkzreVHh5OC8BHf7bbgLR7Qmvil8iU9pp3s/Iook8kUWD21A2FMa
wpfZuCHyg7xG5Vx2Qp5eUFG8nCGRbE+d/wjY0RxrsLyc8nkR1rmH1io0iBgZ2kI2
z4vGFiNcf9XWqlCeTc3U/IK/RTTftwBX2bonWA1wRGa35yQ4jFCohS0PDlStBT+G
ndBdsJYQUr+ErdW4EO+Lbu28Ml5oacNkdDgtk4FL46wLoeujLgjfVzd05dmZy2Y4
C/cEUpEoNZogceDwdlB63dqGoMQ1KKVh7/49kAdNxgjlNDa6ZNKgmHNK6o1gUzO2
5CI9RGVslRdt6VXuQE6QT8sKFU61/npqq2zEyDcbcEBOIzaI9jG+lb46i1DDDdvn
5jitH29hrl1XqQdNJy1ORc9ZUzEskrm7xVy37uhWGaOLKfEu/3xJkCHfxUI+iAQU
fqjz+zLvQmYxuaINQWCXqIraGBX9+fIt8U9/msuk3rYCXVEg4Gc5bWx2xplOj095
Xu3t6mThM1UBNC+YqxGneAQLPPeqdiSE5lbu8zcVRtKpjY89LJUFRHNUcshtW/+F
Y9+22nmyGzXldZPs8GJ5d7Jd+9rxL+4/zbLWujxpU/vNk6b36rXb1kddNcOcGc0M
SV56rwQLXb035aoipgrd+VBwZCpzfluv1BB+INOpe/Fmf/pg4oHRgYAedARCNZG2
V2rgQUFy8By9P84FhbFtbkqbZLZsLWM3V6VUx+iT1hUln6AiehXiKxirf7JlyA/1
dYibTzf5S/791houCz1bbH5Mlg1Lj1SUHTXW4ik4KbncuhqC8GL51bG//CWGhChu
tGwlTIgQQ7DvbVQyHoaMLKYtHFy53JFbLANX5i/ptVDxgrwGDgEeB+5b6TGpcBt9
dciyb8kNLpv6gl3HcuNDxQRZSUVW3ZuyXIrKjZ4zc2lou9u5y+iKC5uZUrRee9/W
jsFK6fEGjj4QYL5HYvzsiudyVaxCzaR7IzfgsDfFhlkT89knerY6ZETKyR+EuvRb
86hpnxcc9Pd0eQD0z5egbY0sKklZH3Spm99WwMll4H6+UlLjirkVqSYih/xRMtFK
HYdZ//lTvkZXPwTY51CJs//QmYHy0Yrra19GBxVOtS4L1kuyC6hBodyAfbXh2Wt4
cc0rucPrNGv32zS6MA1mOO9z3by9oia25PYJw/7AsdB6IJPWQMart1fpCwKxW3RJ
hAWboS0gglD+g3767CmCVCL7tMADWlL/B2ZlzmKKXPYtg4l//J9Jn5Iu4cG/AnFL
hD0i2ek7ubd6BFF+7iSGZfgxdFtLppyiWd97mGuMqUMd91KnlRq9WeLk88z0z51G
UzX/jcnoobgibzZ6Dc5OZd72jKXkRsyOY1cpqTSNRkQu7D6CRyWoFyXludPH4gD8
xLc6A+Ef+Sg3KmQXxnVxJC2C9HIJRfcFG0rvx+mMsN/6EsE87/IJcTyn84HwL3XO
Dmb4lmwjXEyW/IClsqhM8kVriuDnkM0qU61skn9C/lGsIzsSeGhDa568ezP4K8BH
H/391Dj9izkUBemy3EfKKiQjPjt+HAIPROK6V7eLbCjZCZCvhGrTyBTPAjq61mV7
4yhOMgLCTRkfwZ9RYzQTk/ISW/F3bTyo8dWulueeZGodp+Em6xlb3Zp7bv5rckKg
+B+fkww+3ZLz9sYydUqghsbl17y23AZJ2Gsl6bOOpGNqbYMG0yh7pUjGvirvwRbr
I7SeIZB91LAK/Hazo3S4l/AePM8Z1zlC4YgSp43awyIOWqbkwTO4K0RgvkHu65H9
J4XVUgqDjsliZb1poBnTUSox6Q7e9e+pn2YI92FlMXJqkSMmHhhLNXaavZqvoqSM
GewbOV9DNVsowhjkgmihjArPh6b45oRUxYbITx9nYMWjf2qhNkkmhR7mFgeu33JI
mIGCncZNmYPzhTE7EnLgrhp4CveLmDUF6yOD6/1VrD3HlNXPtfZ/a0MvURD4TbhM
Mahd12RuWVRyR5RAXl4Rvr0zkOlaSSdEfDEPCVIF4hqP5Ni6s+FaGzN9h4wQ5sAS
pXRbmPJN7H/piQZvgQgZ98QFFs2/ebc1Dc45MopL10GW+Z+MDyYLP/6C+WtiUCdv
pyaVTg4N2PplODG2qrIosmwTROXhkw6AQDGdqJAXpdfQAAipdiRMJW3sETsJ8HBJ
w5EDEUH5yVoOx72A8U1nAYPYbwZotyZcJLD+Jp+mtH+AS94XG65JLI3XtdbJMwQp
otc8v5yL64OmPNA22a1tQ4SLC07zzoHvbMAw6gc9IgkaNQHlz1/zRFP4kDcMsE9F
xN4QpuDouMYbMo0y9YGbOlgJpUiI5pcd4FhtvBKnZTHbsdRYkrnwa01PYH9llK4Y
XAgX3HYlPYJYNORqAXwC9wcQgON4jwX0G2whJEb7PVKrvGdZHfsOLVTHUVuxKANx
3wc3/IkBwmJmzWg6swJwmpifpWCT67zpSi2ioBcSbponSdMP890qv4pJ0eSYOlMb
rdDbqv5R2yuDyx6N/41nEU7b+cBDwxSDe3c9zu2WWV6KiCmwajdwpsCLUGdv0iCv
+x5WG+PbHl3fWnqqYhjOFGu8LO0Em+Vn+3idpmWx7DJBJngor4UYdn5Hn07eXbS6
gwYLTBpzUMuvftTzcGSMQVvdsBEMfyEWKgDEVuVqueWYptAo0Wjj7ddO2xv8kZfp
l9ozkXYcKl49fVeEl2d0g4yZEm3rX2HSv8Pgo65pqUJKAi+MFlDg15uMYUiVDUTf
UY4M4t+IrXyp2tPxdq/5vqA89rIZGNKNoMvigqxI6SvQIGcs9QEF0GjhqoVtnPR9
+AP2Y0EPhCQFSvuKouZp1pmyGbR0qTMwb6ZX4dO7pItwshfcPQX6Z3V+jP4FWOJL
LXOzGWdBZt6w15bPatQ0lB5DGRCtZLDXScG+PK17FvBR5zcVrIp7UTWMBz1hLcHu
hFUGEdjRF6hcubMxBz/nElNDDEX0/BslKulMqeqsG9Gf/iNgnwNmCWsAbyN0E8b4
HkhksW2LMvWc8vh4kheEZ9rbmo1HnqRlH7nwdJuRLG8GrYwlMwN8Idr+tRU0v3ei
pTiKJ0e+X7pixVNVOlMblrSGiT8QHQeTu7TXwKznDj60H1Dh3+CCaqKvif+2YL8m
MdpCH4RCXpSsYCghq2ZX8DvQJ2XQBu9oQXR9Anu8Fl1FBE9hiDijmg/iAe7Lyv//
0ZM4gKdsen8BfGEyZ9eZiMxnJgdfTEojyCmraf/MZRZZRXzv4g/c7+BdrXl93jgQ
jdURMPO4qXQGnZlKnLNxIOGHGKd3HYyPWIV9nD7otVkCdRHpwixy+3vX8cQunmGX
6lLnsUZg/xo3zmAIlud/qjmCPc0zImHQSeyUrPpyDG+Z2p6YChxBf4MEnSdDIc6G
PE6MrwdrbWa2PijA9RyEANf45DgHx7G7Od2VuYWSJVsVuGQgSTpPpFuuDEc5OkFx
Koq0XOOg20TK9IqV+tgFXO8cydOrqpC5u2Tov3v5lrBaLdskalj6dFv1w3T9glU6
rSa/PIbaU6HXX/aSjymUwsgiRHKQRBLMDNBtxaoJHEfFeYw1z1oJsm6vA3YhQPQ3
+Ww239bOG2K9laBuJ+60KWFbGoWrL+zfqO+bsL6QmWzfdme1YWI/nP4tHasYlEFn
iMlZ4k63LiykaVse88tVbPWtrWeTu44ZITKn1cvCyqZKLZ+RUjRiGNPoGST8/n/W
cmHmKVgVjkV2m/SxHCb3DTBLzrrRw3ub2X+j+CvFqcC2gTB28JnleJzqVGvrykYd
ND/oJ6BxAtuKH52vsGWt+9Vj62Izc+racA2PupVPtuaJ0q9OsAw3td8URdEbPqd5
NzKDt6z99PN5cI3LV77pKUzpanTFzP/4Wq1tH+vS9Pj0uD3/AYXEJn5260NVfJCQ
RWmTWN1wHI2eTDhozKySOGW6VAu4wPuKVGhV2xg9Kcit5waqMjukxRczEUAOt3bi
CcGKldcmqxH9x6sVZ3SYqs4zUogyxgWsrqDBQoLKUI+Qt6g7QjZcCox758zrLbhK
5fGibx7f7PJcwaS+3Kv7Dc8KXmbw7UKCg9y9CPI/PyIVb9tHUXvlKrYTBcvv3zeH
XyeWf5poQKno2fKaFsFFvhAOJequJmWWzcAkXZLm6M5laTZhLbW7J3K+/Frsxz1j
zkxELjzrgE0MEW+l3wcJzRF1wogV8uB/B3JEoDZ8Je1JNQ3wmoe1zUy0WFGJ+2lI
1o3nXGlByY7vN+gRZd80UTPBFnAQW1BEy1xDtfcxfcHBBWkN/MfAwqm0gwfkw2Ij
tBH6f7cO5VvaPUA2vPWbL0IpbNQEIBg1OP1eUUo57ETYCAp6FBzgw8lVkyKlXyBq
LlRjoTSwKwiTvbYO9gw/a4m9pBeoBQDMkXWFqSEn+KWT1yOh7ePKA2oV/Yfn5ncP
PP0+2hWqBe1kGycWa0zOrlty2+gSW6PEATqj43d9lPVvIhuXcpx/U1BqOq/bL00V
tzSj/zRvHEPNJlDzMu83s+Vps/izGL6axsPizXrjmsnu2kMFWkFBfBJySTvoVmeU
Ns04+iT/ZuSwGDBp65DiEZLBpTnQ0DkeX1avJGvSWgFQ9kjiucI6CsFBgEefj5BO
swwRT8Yv7qSGcLSwIkVKeUhimqxkn8eUjSpVdh/e2oYnEeHV1n+kdxG03RGUjnd5
F984mSos+1ArhW5DDgKrTRo1/jiombZFKS4XsgECI4rKI7jIpidDkKhS4sxl2TC1
PalIhjomCf4WnSSkH05HeGw2mTy7R5pVF1pR4hePd+u2kx37UHW2mJtxLc4wFV7/
yu9NeWlmykpJaGcMEsH5vDCGPC77MLN8w00EvGO2c1lkUlgmdwLzWBqyW5TzRhp2
HMYtsfMjT1gUyafVSM1y+bD13+XnzuwSeUd7iLIyVMEslcL7WONWsljdViIN3Im1
OaF5I4lVkYXoCnT/bJCDfzGH19JN7GDHx99ua0LZ5pkbTUvjXO7WC9X2cRXGlreQ
m4TZ7MrmLCu4lzicaszsHbrtAiRc4B0B/iWew4K2FrmKl/V/klSuZ9beIziSJg0o
/OxEq5gtItsY4iYcQu/M+KkR63PNkySaSrfuusxfscAat42lVQHfrKkRfhYkS3w9
L0l/i73XSNcf8KvHMcRcjuMxWkj67PfpsFxqL2g4ze8ICT1iypf5LnhIsOZ3JRMA
6d8VCVoKTvf5b5xFiiAT6nT7ATeX6/UIeSQi+FRFtCF7IhrmXV/UWBHsbVyol6xq
Ax9ZbPrXjWk+3NPCnbZVdrpO5YyM15CA55G+M1tActy/Mpbu9RyerIPUzl4qYX9R
gcP8gpfCGFd+QucQeXz3vKnDsmyGNwDTwEw1hAfYGJn1wT1bI8aFKzo67tNIaz9a
WwWzdMtEtnG04IbHBa1jPeRs8zH1S4eTiHOg0zQl4VCztdyHNgqL6Np2I8BWqL4z
mDuizkeRFVdORIlQLqcF9jw6Nmd3Fa5eyKsiVHiumM6cbDhZ4rU87rHrbt0v4i8Q
AEX3TF4Y/ARP9t314dvNcupuFMFjy5+EYOBKYClfIJiK5SsU2P4WvFErIGvUe71m
CtSwcrXqMXZsXeIjNd9yGIUdGXHcN6MwDEmITERORRjrUlEEEpjUWDAR+wIVOxOR
ElI9rv3Oz7LAlXeRT+7KTuML7cbjU4dNKK7/ZUVUGOgQCJqIfb9k7raovfNP8mi3
RCikYRuC/JzdyIeTs3zGU9ImYQGGeUgH9frBMeD+JvoDLXaTb4FXBtvSUeGaKk57
AxmxIBwM0zUGhvJBPAbUnmVfQ01cUMN5ieuBDJ/wzGnNeGNqfOmKYBR1EU6NN/dF
L0gLtMlA89f0VWTf3/h7H1KPYvNNDBANgK8ayDK6HqU3h0/mrTOFn32WyrkRgEBm
FxeGr3+6vcm1biSzhuavet4g3dhgxLvwclhjUPRD9rhp7AJVUoKf57s6oxU9QmTR
x+kqdG02BjXSTi+y0C9E2bYwb61chSiq/y5ZcnFIXMxEphHC0p999aFtmPDJniqM
A1mNhc2bK2dDXtyu4Ui9skttlszUmkFPHmdH71xf+06ZyZEAQ9JmIKWyyzkLE1LU
OHXDB4sdHAF6jnwcW3uLJso7FU/USZ5RFJrwgUAcUI6jeholmxPIDBIVt5k/9P/l
FghsBnrN6CnBh54bYGRS/eD8e96EJqIBKUA2YwT8P8GtjKhQXJLD35B6u5Fql6Pp
enzuAaHNX2yYUluY9dbhJcN1Ic3R7ek1+5FK/PV8xk51rH/4ofpKCPay6eElQO31
3MDVjUdYkZo9wBLKREqWMO/1PjbYAStB6W6e1crzCSWcL6jHQJisVpD3j96yVThW
9G4bGFMumfiGLxrWzQLTSZX9ZYg6ZU/+ps7vGtxb+ljeT4RgCd5vcfO2jmWHM8Ps
/vFtIqQVoS6ubDFRuCjilt/27jmdAjWeTCZWlwmwZar95C8wpVL+IuIS6QyaVxEG
rvmYSAtEph5i7LuI45wTv9kzp499ouqzI35g7eJze5IvjQuypShhrP1LZp78pUOi
+MttTmdX4qNcmK4MgiSOVJpvnkzBkQ8I4H6ECTGF/zQr7/lrFoWzyqToZAL7Y5iP
h8Yr+bmBaRk4R+N3dttaJ1RMIQu0Hva/gV/6KYkmhH8DmMxEGyePqHYt6p3s5W/E
Wgm2V4MgQfYFuYaMagRJwpOCY4kyvCTWS8wKDoUMLb6P7AjVNi1BHpMzF8dFV8sW
9KHN4iR7vFNWPN3tj/yJ/hrGNHBLWqu4Y4YhInF4QIi/wk+2wPhJ8ouvXBI4BhN2
WuXelmUnUhcxhUK00muz1KQM1taQTG6cmbWuQnZ/TYNquxmcGxzExOI1prOOIlI+
mMHDy+jn/W5sacytTMlJ9lV8qJqXnu7zDsEuRSI7dSR1LOkqNQlMK0WruLhmuCML
4aInLcmhyNzg8GyNjrjl83Q+Lyxw0B7RARBNuChJEGT/+JUz5zN07C76ZR/UTC5V
HTmTRL5UelVp74lXwTNeJd22OGQ/TAhAVupkhkKPitBlzSyCUp1GWOeCSmyW2WQC
gy6f/+iwXCmiVh6gKYGDLePuIIunNskmr9HRZ7W/FtZ5FLmMQaujb8CQ52Mk4dNf
zVyJur2Hqw6lcmP1S8fFtjMVdcIwTQQe8Vi3W599csc55/lo+FHpru9kxQvP342m
sdYMQUwLdybJOVzu7eUItA0VZgeYv9duJlw8/cZwj73QXe3CN2xL0pfpEhexdf8A
LeJuag0zXa8VaLGp1NH5MTZYiY5JgLm9gT5p6t69Gc0vtj+MYmlMmBpODyKeKNxo
8l2m1yfg6zbErRN8e5bcrJ7QiM06o4TXOycWta9et1CQpx0X1IUb7MZZNxAmC4At
r1K35QjBV09GDORvQc2QKdo5yJPsYfTMb5PnR2NDb8kjsMd5C0JvcQGf2gSS2HUH
wBer/A9oTjXX9EH6sFzKey8cMgKFRLEpausH6jmS1zqT0VdrJlwDSM8FXT0d6KcZ
xB6AiJi2VKtyWABobhPbIb7lZ+f9WLydQKlNSWvSAQIcltKRrIuDfMZ6/U+RO5+M
P5ZBegFk/beP+Kg9SJ8tfINQtr1hCHtM5vTw6MNWzVXAESUX0HlJ8vdb8Mye04qZ
4EIUO0yGgAcnZZZO0kkAiTUaUcp3sdPckNzk3xdp4ObFrkTXu68GAKj+QjThWCkR
GK9yDWmLr2FY4pUOwYS/OsdznFDnw69iF5AnUr55z+Kn0fz3UtRKz+C6nZM/s5vN
9trf4eSMEFJ39YWqG5Uc/T9ZOXY47D7I8hjsjbw8PLoITbwi6z3KaDgoWB1r19vl
vIFTwus3xFyiQDZ9QOcF4R3vxhgcJ9YEXmk/1hHoqAB4i6xl/jW5Su8gwBJs56HA
W3atXj4ZPR5KAxTUM0Qn8IgJFGVROrVhI9YgeH3cdfF+Uyrkg0NtClIO19lbbVCn
MuurBmA4n1w0Tz+oJNAz7FtSQnHn+mQCDDg8kykCTh33us1QY5khE5+fEPZcTtC2
B4Vg/bbHppP50voFQOnbGsRFbnlyqjjZlOCDCG1K5mOWRde2YSOybgVKN4JDwCFe
DFJSUIZ0hCnynnArqMDXpmc1NUYcAKrxGwGE1w9jIXplvFN2VwrEKovVv8Cn3bGb
GtQbIF6fzZF2LbkgtEHh7keiiZxW8AGIepAPwpBuj7AdPcOPauAmchDt5ptVAgEX
wnEGXZwLzR4nhNAK2rWfNga95ew2DUQEEmqlsMwCXSydKDyYcfAByKFFjSeaqU24
n7CCJZyYn8luYqSKJ7fa5X3JxxKxmZn9i5mm5Cny15o=
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36368 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
9GNfeu2LhBO1rvG6TqMSwGFB7dhj3neA4P4KFvUBgsKAs4NWIdD+wRwX5rjT3Eyu
beyrO+B4kpsSz8kFkVVkiiaruAqjrZhTzjbaeQaeFLbRuNdzK1SDIxo0luKA0giP
Dz/KSt1epSR72zuYvYHXnOzgBMXSq9MAlHfSpI6bcGEPMkqqaUanPtwHS3rthJ3F
E44LTDxA0+2vZe6TVcIxYZNR6nRL7rj8XK7l1tI3NpW+Tkzq56EEb/hz72KXmvaT
29hRgglXxxu/JsEsGeURVftHvj/H230s5/m/6jfirRmakmQVVP3dAGJFaXTLUr+s
ZX0S8uD8iZlPXcxvgMT2eupozL+jXlXtijaMw3s6BYpH58HgNd780HfkvU6xM8/p
J7AAabCPeGckxLZVD6/wjn+wsKRRuQLUDFDLzkh8PVRA79h2ExVJB5P1Fs97aVT+
uwjF62XBE1fD7RuDJPL3nqP8ICYtejuuBnkCB693IPp8ahO6Ynt/Yj/3SBYfgrY/
zPb3GYiw519lWcB/IKmZTSkrPfFkyw/xx0rMBUVOcZ8Ic5SYA2Sg01jb2K5KTOCK
iwum4JCUV1hK7GvoSkyALrMih5ABo5XDF0oF8X8MBU15iI/pncbqp3SpdUGlLYjd
DgitKsXIWtU9yVe6kSaLU8bfk2ivxnYaBQNodGSwcKezOkIf80WtUAd8MZjujsvx
YisfmLQKkVLx79eqVUr3DJNVuT5c8K3RrPTl/srIx/tTGZ6az8y6IJiQo41FaPE3
MFo1k11tB7xfwKPsBKh7yvMXq2s7enftxymW01Huc17fC3fvDVTC4tDbO08UQPZu
rQg3M6Gj3kpsGqtKj515DpXrUi6O+QXs6auJNLqp1TZvOnCgUtQTvcPlp5fNBUzg
GYgH/tShpMdNJKYaMOIjUiS2F00fQonj8dH+6kTZ6OgGjvGizf/DMOEwvuBJibLv
lADtFWDLnS087UsaFq2DDEE80XaxU9aXO4BSk1fQjnYoGprDwqvdm3T/8mZtwmTY
1A0ykML4UZcIvntyekwDJJMZMrLZEvQyc3R1/+Gu5IOsMMKjdmxZvTJFkCqKI+cj
4wbdxmIibtgRWJe/vMHmUMpYv/3WQOOzMEiq/mwdMtBma5onhxfbt0Ey025o6OQz
dKVl02d0/EOpE6xU1JhVZ7uwXFLRUsQHtAWNPA7wuCm1xm6SeuPD4ZYMd12Onv3Y
pvT98GTulun22r9/QNR4gzX8knukNwPLw0axs7Sl+1vtqJVzLkA+qkSONl2XXO2w
lHA28+dt1sDOojQRx24SL1Z8Ayv4dj6b7jyTIVdiRi7cxPbGPiPI1yOgQJhXhaMK
a7RYSR9PHQXlc+InQ77/QqYWYfSLXrZO2pbA5EaitBIAyEHcRTFZA0Ts7TBuZ/o6
DmKsdrnvIYk5cFaAWPaEzFUAxC/zkKWcArlyX+6O6lLkj8/KQb49dR6qlxqsuM2K
AiyT1+xWzbj6qz3Gf3S4x1FtQnXHh+J4WdWTdWHu8Lx3p+Eg0jIolmfPEVbLjgO4
d7z5gYqyBwhc7oy9ICDRX96mWVm5qk1OU8z5CI92wecELxO3txu+9838Ri+6L9Vi
bfCsdmshYwfhSlOJyFrOpkOWsYRl9wBZXa8vdjUZchz+mVeLlUWlavN9TgtNi+7P
OCUZtxHQP9ycROzn66MspUg9CQbl2bnahoRCUuBLuuQY4bLBsd/FZeFnbA2MbN0C
1AISFDExsHFLwS9xjRQfXAF3BfV7a9KClmpPUX6qPEb4rhbzgTQzUJPz3gfsvlpC
WHboKqvo4bIV+Zz1WT9equb2bH/YbXDFHPdzJW+QyjxmMdbf7HdcD+Yq+4s67J3X
w7BGvAY+O7vBnChuXoEqv641g5+4I/LKKw4f6pyv/1/H48oL8kSW7prRjvpfGITW
S3fdZpncWulS1WiXIMBmSZ0AOadWkaYJHYXCd24vGRhPIwt+HX0oyLHXwoMZjWiH
AzI6gEJHOp9z6ej/iROb4+ZLpd3bOLjNgp/esp8x6wsaTsTFgh7F2s28YIW8SELy
92lkY0mpxiT5mn59VHNzSC92Vk+fRplnn1DJrVbixoV1Onn0JsEdr2UBRwsNE84z
bmWpSYU/HnAxkM0rV42Ii6XK3ywgklVLwOk0PESGhMrvtD9bmNwhMSo/V6KMgJlD
KgN4D2hjvexOr5oa6/yJaduigcaFitUlMZ1+Eia2Uph5d8x4bCNalq+t0U+siq7B
wIWgycJbOvdCfcioZDodwHN9HMpLl0zylficTdN2lDeBcio6Jp10foJ3WEoOcm72
VGG2rxj4caHnPvBW27ho8QfUmhttqvrXLgc5u0B6T+Yl+leAx3PDxjPhD1ixG941
pgueUuJjHxz5x1/XXx3IccBCvyOEoPWY15Mnt8Z5rKrqXfLsgpLimAWgTh/tSrNO
JR+GjF0xtkyLx+Ryn1CSEV5NjEHKQEj8SnZppj8GTHmwI+YnaL6fVt+xxfgS6daY
QJJOG9FbOInfC6FD2N+tz4rqKYe6g8QB2MgZUM3vnsTpDvdTb/yHWeB3c6WTVu0K
YUJmoFdb67FdkoCrLdbgUPwfFildxnk2DyzmZuOF2O0Yatn6vRre/Go75OaKoiFM
L7n8H7oklnNa281fvQaO1W4lJU8ulep3sdKTGaI7GFXEdfLzLRYtu+SWvMqFyalD
WCj88E/c4DMZyXbA9DDn/UHOt5VbIFbY9b8iZdTswir8CeColsUoE0ojk2YuWlF5
TmF4npzzEO7le25ejQNvnqLkvJLkgTQS/vRbQGxP6S7TpGhVIKcrw9U3yLTMfllW
VRcN9Iug09cPO9zAsL2vrngwpEqhRxI+pdKxuBzlOwsIXgLIQj0UU6ZFd6OysD+P
kmzlaeUNus4Aht3otJCFNdQKvfZSq600mx/99XUSfU3is48O9rkLvNufgsmpdKHL
d3X+WzzIFVbewiPqogs7wXBCCnG9Zr2Vi28733bMO1qNhjbWxNGOE835ojxufOSd
nxifCVufW1jDWurw1jf8SkAWGLtHGdJgdoZA96XlLThv+OqCWLH+xP+lc+Ybps/d
pf8uHwY/rUoddzkJA/1yddt3Eev9tcIB+ubwzDVpd63cjQD3932odP4x/uzfj0S6
2MgwD2QoZ/CYuKq/9n8aemiHiJ5wTllXE99gP09ynxhUrFjI1oyWi1wOaIkxrTbm
muxPSiMWWkJr/F2TFXF50elotJacoz2m1ffCxzXeh84+JGlCqcBIbiXgmVE1rOGW
sXhSu67ieymgsemvXSicQjLOlXHm/FwWrDeTv0wc5fq0T7aPi3eZKXbOHtS3Ay1v
CGv1p+RqiVR5JQ0lctNVpf+U+QgPvwduErRx9tfM/fdsnuCOhNN48+bhjlRyHGnj
ClFNKIrYi2FnUGNpikBczG4NKp4Jd2LdjOe3IzO0jBss/uA7uFWtSExIiMsyWCbz
+Z+kvnkBBEv2a0c/4434C+df2Jzd3UbMPlSqkw6KtXn8GiV4GrDGNmuWZL/CadZi
0EXc7B/IjsQTsInbBDsSqU0cFbpYabqYEHkljACrhhuCgBvWj9HZq4onGY6P0YWe
GeAt6B4SuuTw29CV1OQ69S2fdktzADOzOvVlPVUlOMqI2JBeg6+zqAbjv9/gXnYF
agZ7Q53G6utEXaSDhsfcHURpQ730jgnRwDEOzGONnPPQ/uSxJiTp3O2iWYG9e2pV
B9Hc3CgPEnPDF6RiqhNrvGeGE4rZJiwFwzFv7nui+ar1/OiW/ROVpL1Zey8Y18lz
Yfbir7ddLIzCrKhqUDKDFQfrbkL3w8L4OaSNBldg6HbgWC7EqD/B9fPSnJrdrnWo
ZYNvh3v8VxxAfsINkuh4pyYSATgGOK4mGO18IZYrpXUoIGvaZH3q8GdlrzVZw7o5
6yH8pN9t5XzZPPEvZkWy1j4nZx49yKbPeN523GDoMNiYRpf203bnPOBblEgw3OkG
m4tQPiSeXDzzUome4MQHDfg5wRA73STpbXM/SeZjS3jJTIhBCA5Y4nVBl0JSfaQj
Kk7TcHwG0NRtkkHT2HqdEXKvH0Xbqkmg8drCskUrUPPQ4dokRmB14sDqegi0Dd+b
QAkMSjGOMQhiQ49+qh/E7K4eBCUqACsJTb4ENmBHv/3dB0DxDB4/yQwsSen2lRg/
ZWae9wGtZsHhfp1liGUF3LKU5Pgy+pnaJDaAuiqpk54VhiKPKKoP4Ps/M0KMZpIL
jp+aZpYlljhJcV6PLWpxj/PB9dfayfTa0gmRkuUZ4Q9mwgwih8dyOKco6585T5X1
hG2/4wuQqyDPpGNtIjwW+EhwFvkrp5xEBp0h8ZSdqmBJrkm9u5EHBUOFqfNHOd5B
96lRfc+QeP8kppWHTYWDysD04tpmYCRReBlywZ38Jem2Lkp5cBqhVR0MvD8f/3Dd
3RVDxCxLzRaHvHzkNz1gMbRDVk+WwJfwkA2MIso5Agj3SWeMi65xRdfINDqC+g48
pzxaAXfw7XZ2t/r24bbnrcPR1rfHMFod9/JksgncnwIAIhb/XoRkOjvR4W1yYXeg
QF/fu6liVk93koeUcDK3zNWfHmTN6amA5o8uunJos473w0NOtL9yX7SN5eAjrfET
PpYEOxzoHa7pscBhsBPC8bGcAf5ylu7I6JQrW+7xo5ZY6fEnv/SIbQkFYDlINPpD
DWwtoVPMbCDJu9nR8qwdg4i1jqe3zEpfZqjwmyfd13CkiKzAElr3Qn8GeVVRPAZ7
BD8mOzG07R0XJxvTOd5Ko4b/1dePKNfIU6tm6fOWQHNzOGE1g1QYHW2dEDfMd7Aq
257qJUq3kNq1o4TubopDRjfRR6doXwgYWZiRzOYOMz2uGlSCPhprVdqswp2dBSi0
ILhOPDffvD2ElJdHg/0jLFcSV3zr9OVpnO+NZbW9aX2E8WwCG8jyNEggLPLYiSzt
YJUmvXdn1Gz+TOalrNxIYcqUj4et08RR3GdSpn1O7IVeIV0K0KcQsgXMOT4yd38O
n5Pf7IYr0uws2GGRjD3bUT2UqWy5MLVssnmx8m3rjBGhiP77mwOvCtsMjNa4CGNO
G3ZTTpccsMz19k8k2bcJSUkUaD1IVYkCFK1kK56aG1xo20Pf9qIRNeB5aO3dQ3dZ
dpXZdQIU63uxoLGV15K1POI5nOH9/KZOwSJ+GOXyDM6empgoUD0R6osH3c4ibApy
cQ7WJBX8VrbkqdRp1Fv5SYNrrSVUjzSuRNjFsT3f6zLJLw4VnajYKvla3M1Ty7Bq
C33mx+Ld6fv8nJlS4XJoomIRgYEaR5vRQ+4jjjAgr/QDknI0cloJTAPy1z6FejE7
b5skqXRE5MDc0XFVEGGiKndFH4VtsVmV3vYK4GAfgKWiEdHTBMVsYAVZZN4nuiOA
QW+csNrhChaTXV5n5WhNW458DfDvnCObUZ4+qMfmLodY40Fh/JNdx0t+qH3TW2qO
/Rw+x/YsBnuNLsZbwlqe05WEsx8eU55otlv1wdqWXVH49vZDfDjfdBWS57YIGezN
GBMzajgWJ0aInDQwh4JY6Gzj01N3GQKaDUeMXrEMVYjQp6TwvJpq0h0R09IPwzpA
naY1qw/N8eMUnhbDjRyPZtMROl1sL9imjRcwEIUUsAmoyz0x8RvH21g/h60lXlJo
VfUcPOe6zBx4MtLgLwsN4sUm4BfUZajOtgcUJQGe+UzLz4JrDMUkwoWktjFGwqC6
QkQprzUUc5TBTmFchMp6JiSzhxvk7UY+LA7GtHfKr2MgSk0BVMwoEqRkwpQ8CKDb
6ChamLQxjt8kVZLQ+AvzcWpuAXY/Ahv/ZlxV0FI+MUMsV0wZstD0J/a3cP8eqc0U
CEoOwldj4DoNdowmqheITi8lrvcx5btlPCMSO6dRzyDqfq76kVmdGZ9PhOn8nHEa
JVTtwe6ycxC1+QU2neiED0a9ETtRp1N8NGwRpki2shFGiNoOGP3Sk3PADMFS/RUz
sFKpOmVsA4ZC7e7t1yKgLBamgmD+URGXiAph+Wk0Y1gG9Rz/BkXnhEHPLKMj7moO
kULB7scWiUtwn9eJlt17yf776TUaGfzJ7YFAOg35bDaPurCeI/sJqSd9UFhodpFA
vpjv3diuhq2oUNikgRFhs65Si11M6YWl6gCmweb44OVkDJd8UN5Xat1EitftdMxt
Ax9FJ9T54QXDhGJuWL00QRhz08f/ZyUA1IrRECgnyfOEq+cDbkzCXh61P33dfqf/
oe8u3I9b624Gc0kSzOVZapRj1nbMv9GnMMv1hnXECgQFbHWnoVFB2jael7b4b7Q0
4oyfJ6Egae6R3JmTTxh7GcmUk59vDdX01YwxR2NuXINfXGJPvTO92gbdbBLAhwKj
+7U6x9YMX5BvPUySzC9QBtRIAtwHGEsmbNRYe6bm2QKQLJpqn8DlzPWnSANPsdod
3vJCA5F7yRbyto080FyDsnOOqZAr+cHj0wrsmcyYSjUbN7BvnLfh1CjeOYVBaGF3
lq+24ma+RK3H1JNzRGw6LmwBphPMMnpyyfURZVKrGbdvIKXFJJv2PcO/qwv4aiKG
wvdvbsLEMR5VlVPJsYoLRD5rcf0n0S0cDCrJJ4vqPj1FKa8Xn1ptnxcpWzVjZm4U
s24Iul2pB5fj8iX9WRaf3V62igszNt7I1A5epZufZezVzvU4dOXHJkINlXxg2kvY
ktmh1YXhz+aI/OrKv7wKRsWsQOUTYmP2WY6X+qybHtTlavG5+nEoQqAAhyWK9V6p
sklsh0kc8QPQ1sg7PKhdZFnulwWOV5lHD2EG3gDQRBJDokCWK5hM41Zx2j8HiI5c
uKueueAbibfaBLoA/56ytuBE6Oh2Rdvh7onetdF7BavufGiJFpD+DHTSqMFDnHZf
wycw+za1ylYXliP4N0iCR8BfRF91Lp0q0FU+vxBNY5BKX17gDr7iWPv3OHsF23pE
RBQhbbJVipalvVxaLHhHexYFtxtX9NRDpZPHoklBixHpqizzusiHypi9xWMpQEAs
+gg+2qGHZ4kciYgxVCl9wc7q4yL5K3eXel1eLpMOtib6U9CaUmP8g3E+tLMX2wYE
L8Dq/KCcn/aDCrUd4R0RNHEsA4ZgnJAomUiIBtHWNwEotYrBfWiCXk6M/r/jVjN1
fBQDe/P90KFHm5BGZ3wtKTrBI8QMxDuO4ncWPx0Yd3E2OZtRrVzGm0QPGgLpC6l7
nHgZ7Lq4y3b+qqF335MuEROBzsfyVywveT6mpSpCfAyHAgbiS2jg9nOhQP+LtBw8
eA00O9NC4nWxsmiECpGNSWgGgjgnAaFuGe2xK/jpgE4Gr5Kqj/AdZbRWjIurAIi5
UsocaalWAQyT+ht8OmRKjxgqgxgVj8Ywxv+Hcmz1JVW3hJgMgG3cZ7pUWqYW3Bs7
5d7Y1QfZZQUX0CkyUyoUhgIS+bjmF6DgrOHancR2nQ1MyNzeJ9IkJ7gXHOv/M53U
yRUAKJBsiHkq7gl85uE93/I2BZwfmW00GS6mGHNmvF3hK++wtXS6UtVop6DAGXa0
Njfbj+TXzIDZfihc7WlgOd1Iqv1yHeGPE5ES2btEIKPIwg6weG8UuaUaVZ9A2BlM
29eqhhLbNQcQhpjzVz/UEMhNsK5IDMVi+dY4MiRCnDoqfK/KjEAmZy92jxYVsUrs
TT5+QdA/Rck1SzWcaW81sD1iLF9hpfkatI1PE62TSVmOKlqx/YIGVcEZAkGssdI0
VW5Wwf6YZLk1a1Cp4zALEKzpuTzNQWi3qyy/dFIY3NHncb+cPlHA8IxBcNzwNWcr
4i1R3tcyv7cPl55li6XsSLgCpcNyHLHvnSe4zT6KYR8s6Rav2Xz5CTMt/Q5KP+Fw
twyfjrpnJEPnLjKUayHslVyCe/zeMtqLTSsKOlVn64+O4fxq8aCQK3CpH6XhCUiH
WivWv7VORt1RxYQYqd1dUUAZEOGHM316IsDtSwAXe9Sbd5jyIV+trYiCAwQkda8G
oelFwjONaveMP4StgjBmlNUY/8h5XQu8PKuB+iRsix81egLn1DjZW2T+bJtuSKUQ
8qa9jh1CtYRZtD7B4afqTuZ15XbYK97ChBUGyvESaBCquA/NA1+JoTTD9oEuMg6D
q1vZNSKGSKof1xWKX/GfcdputzqaLTtxGXIRMfmU5FqSzueYicMcQTZv524Sz81E
f2UD0DTrAnRN5hPYNFJt/Nd3eXfVB9H7jV1Vz+Rpy7C3WzVMpy2V4ZQEuA5DtCOf
3PL61ULaPAfO0TFVmXeURvlBj8Kt03RMF/qCRIoIjlSxIBC7QaTnfq5cO3GYt3E8
Xfv0JFaUZx2CF3XfirAOVKjPSn/iw1iwe0r+F6V+0mBVOHtYS3ifSM+WaHbDBC/N
MYE3lOZm8w7yd1UiUxf07cwuMSZcZDtUKIAhJ6GQMcPhEdApGjPJy4Bfm3znXJWs
ctFTpTfMAlMSDpovhnnMgD9NadEoeYg4aGNhpWcHLIA3YYL/PpxloTxyWgWqA+i6
z1qdhOlBslsIFed8/SLPsb6ZBfDHe0hl/gvBbE5zSq9FVtcHeDDhayt/fcweCr2Z
vz/WhK3bk3ZALz2ra+RC49A+j9QBrVfgFUbTl+aVtUyZ/JFETVemvN95fP3S+kya
dG6fHn05D7KSIZ/UL8T5PQnC6R9IjvBAFQTt3olHK0JE6awifxGejQ0GWRlsTuEs
ULUzG2tt85qYLmXU3jxPgo9N5k8ALfw/gbVkbNFONB/a28V5XhE5LwjG3PPQoag0
hKEWgxkv3B9JAo/f65Sp3dMioDEvwelbnVF7niGOEf9K/J/97C3a6jg9h53oFn6W
cN0XT8X/tAyi1/HqiXwbKfTH3SBWJ4EBBeEB0j24DpiaLUJHS9yoybdEoarad88u
WNPE++tO8KmDFBEJ4etmuYnIUf64qDuoRENV3otc/8ZtiCpUUn+NT0zplYRG5a04
Vy8xmyNIZuJ06PR3I8hkGSYJQsVwtVuAtWKuhaORcamAzSJnNApoAJiQG8TDI6PN
yKqA3mBIHCKMnkIaH7e9xdRpTs8cFH7BXFIyTFdIdt0N9/A79cgOI880yWWwfB9u
MEeEA+NGK+UkSiTsysIHfGdMQn3nUBGPNQ/JLjXzfO3cOK6qTdHpl66jISgu8mmK
x6KPAAmTrarOMwgGjhgHOmJUsA2NUMpV4FAv/XyNBYzaHUUDSIQ/8qHFNHCQHPGj
2hEklVAvN7IBVH7JptM/Q4qsn2k/PmI+jZgndQPpJrujICvYlIGiJD0jV9po9zwU
cVN58hg0lcFZzW21jSYA0XU61YoUKZGDD5SvRgMV2FElGfnBKhc2Lm0VX2+yJPNX
dOqITHl2Yil0yVw3AX32r14j5+Gs+E8xaoAz6LisRQwIjrUmLytTciJk7lklAtPo
rX3PEhxuY9tPiFXl0e/MIjaHV1wjYdTTpcnhfSG5r//3E6asWKf4IIdZYlDBr0ga
f48RENnzps84CKei7VTd0Dx1uhI0BMQXjuoG5amVmjPRyhLwukDbsYCvsk6Io9WH
y3EUvoqSnQMne/8r9nHpt+PSaAb9yE8HDH1GqBGc/Bv28hnd2DpBY/lsyW3PTetg
RULo/ZIrYEu0vfAtS2EBR4PraSrPHndict94MsUWX3uI3x33uR/QyL0FnUZIHoR2
21HbO8R/0ioAcbJUtZex0edVxbhUBk8yhoRbb75jVP3D2Y+7BafVFIbReAbnZOGb
6y1BQ1zFgzQICEGhkGjzvNzcwJMeC+owCdw3QuRRwMqOy+WYnylB34GxW7RRhf9i
vnafoaTY4kU4iRXCb4B7vLzxzQ2nw9qp1AQ4FhhwkzTiQHBowgpcH7HfvSXvzn0r
PVy3QMpjNNqBMqywdx/F0uNP9mcuoBr+3h7evKr9xsfxIJmDW6iHmZlFgnDqIAfd
td3Hz6jg9COkZvnWLDphjDZ4QBSqdnck3rT28+MrUMPIgyiA65TtljEpbNk3lfgl
KXaq2VhBZmAbpwcZhPPICcQ/DYHQUZjTRtmxnVsluamjrw9i1aggB6uJmO9aFVyO
zJHEyck4t0bfivPZRVBo8x+qdf7Q/cYJuKD0VrC+x9RZDR754aZV2w7ljDMrR19n
mu5RJb+sS3FNImEvX8ZXdeigOVCUxBRw89/murjsQbcjASGLmXm1iojY0kvS/M/q
KMZy/VutohEGN2lfQIQhWlGZyey/Cw1k5ME6+/WclN23xcN4/oOaPxSVSv1217BP
SFBMjECqM7O1MwH+hwotl5PATmhUFhS+PJqHnV6ZiwUx6HiiRcsEPnMwzClyYN25
lON3DQhuU+unDM8swufPbWXVXqXoK2Z9jBjnpcCUpd6hNg5uRJrKYG1F3RJYF2bM
YgR9AQAcmZYgzjsyWH5KNoTamcTZ/FFpXwbmj6OFQSvIryrEhaInplkixZzDlD3R
qK4Z11CnwiMJVUG5EyWAmRdorJiIvdw8qDCjjwN462wEdwSS/ANFQD0JRc5wXhmA
vaH81PMCeekxIzXeiwUd5c2VM5QVbTqEAZ5cHRzwveooNRzplS7UMM6J9/FE66KI
drSxCcpgj0UkdvKxGOmy7Pe3qznd6dsYm8SLUrZVy411siew1DtZWoTLedx4mHU/
VT8/ubIsxsix2BgxkSIpRPcGCe/H+oiF8ZuhmEpSAWbgJzaqf9+ZJTJ3ibX7vcSs
xmMHs0ll2kFwoX+lsmwmWzLf0FQdVhMNSec4RDemJ3xGqPEqYGpmWLRM1TmHiile
09XjW/r9Re/2lVEr30mNZxeVZZtejpWTvXfaC/mJ4lZmqpkLG7Le2BsBYa1i+2PJ
Snv5fTN4MPkz/xqRLQcc08ORPMrWntcwOrzzzdS7YJAqwIqiTVW0e/DKHTMjunC+
0m5ImU5rbLOmdIMDZ067Xz6ZGaZXyRcNc+sJXD5Bw0urxJxoPRE6uhIAbswq1lAF
ysQUgT3NPBvjnm8e+gRnFDnfyxWTF0KIQARGc+yhUVDYEROrnsLJq9DNq3nh5cqO
4D6XO9C3ZdwLqMgZ0kMWAK/W3duQRoYBtZ4t6Xuqxl8im2UfLrlJZ0zQXsd5WFLH
wqTJ6G1Mp7PcWYmhvQbyQbSiBr2B49fiaEU3QkfEPGKnHEPeng7pDahy4m75nnC9
7TaL9iSE8bvuYEiC9KUi+MFIUkmZh2NQ0My+NHxNIFJLJmuQd9vWOLzb/4qgfWmg
BpuiGyfKgS7C7gd0Laol0EE2z5zULOnsClfydZ2yPYirqb+ouptVW1eMh3tsM7Ep
9iotQfErMLWk+JzgO8DKnwaMVtH1rxKz41PMzJsdmoyFEIXKHfRt1dNfa8X5ZusY
Hzhap1FCe6E8ddinb+TSR+ld3wU4xAv0OLZaHcLN5VcRNhkY8hBvV71DT+t+o6Rp
Zvcy+tnwH809AHWXj1zaP/vHRn2DOJDr7VXmlVPOkFPhiGDo/JstdHIqzWPs1Yfk
QS9vTpkOVvm14s1UXGJcM/GRpPGRnIuiO0huapRFSkHI3lV+/UhsokRwBndQ6Sbq
k4Qz/6DsBQuq6++cV1o3gr/zdX7OWZbZSvpI3lTS1bX6+oAgwpw0qxuEIX96jHMy
gG2KAWikveE1ww9S0W3c9VNN6N6DbLidzAGFzzuRxgCZIIuNezLvDT50iyyxQU4r
d8XtcgmdcFC7iOjiNZ0GSlEngg/ZwgHIuXFBzEm+ZcUfStg2UadrlaDZKHI3DO4I
yYxPymFJVu5XNi/viqK5CSRLZfUzH0Z7AjxTVBj7RkDeNwGg5sTjejU5akPfo3Nb
/VtEN7vio0eO8BfImkskZMmHNf0x/aWOaPA+d/cDJuU1VAY+vhTGyDCXnVe3dv1F
4NtgaX+kqxb3Sr13aGOBts1jvq3zYbMdVd796YBsU3lyxlaBecpBZoFS0OqeViWl
V3FnyG2xoITUjXBZTNOLQcIjx1JGoDoRze2jztSrzR96EE7a9D3C1QZ420+L6o0p
hpdKdfoLKrzJVtn7IZYfQ6TIOkn3s7Ct+W865Qb39D4lPeslvh9k5feK2DzfOHI0
pl+KT2DiCltuckzLsjPIaE/HVPXlWjeCtnie1tNR1Y/sKzXENUWgzbjxQbBOxI2l
V+6Jq08a+VMXUUKICmNmchbUMymiZLNF3KRuk9+J+DpFDbGq5HLfzuYQcu6V7n3r
g35wqWUdReuanwX4XA/ctcuFtoQr8JiU/sGcyCMz3htnXRh2cxVIyYxceJY5rMB0
t4LTll2qkJwah2NVh/+eoCqbASlBAnW6e51bGrrhYO/9CgEoVpVi1w/mFijfEyEG
ohYN8miHAp7u3BDNu2BSk5aZEnUsRW1w3Ifc83ppYJKtdvX18gdr0wlJZ7aZ+2li
godFYK7otuzJC+OKr4R5H/CsVgonsmBHLkSbsOhJRNigUhJRryVO+NGYBL0PIrlR
uRA70DEzGxolt/FcT44+muxxrCJ3O1/qE9QhZzboXf5iJ+1Nf5SQRZL2S062/SO9
IoqL9cjQPid3HMgddAOA3hJrrcGLegdVI9Iyd9b/9tN3FybmyD1Pt6B3qWUMeMOJ
bOz35//8TCGkvUG09TGpP3+KlKaUTljLa0DHIpp3itmAy4D6w+I6hbnbqgGm5ye5
bKz8RKUF8bWdzCE2MNmY2ocaciIWt5dPtK5LYyGWel1KoHz9O3DgAjVddD7IZtGo
at84tRRt8e3lWGkR7byQpwlo2PmzJc/OzoCcw5IfupvegQ2ePsMLgd46v4nWMLi3
LMPDfdxFkvI/J2IWvwJchGRRyijHsYts3SQvfA7T76ghLtQyJjir9uMk7VvDc3/+
SU71nsHZuF6nE0x62P8e1WHir9dZfuBaKsz6he8NT1uu1HcG7s8ZuCbQVoXlcZ81
XPSyqnhrHn7wlWV7EWC812rNp90b5pMB5gqQaEOI/B++CeuvMIP53R4FBOnAqZr+
EEKWZgOne4TeEfFQgiYOeNRGTfFEgVGYkN29Ta608H5QuOYQJNt+sdH4cUeP4zi3
b34BAFQxeJogWq+hCldSZhwdbXNdjMVsfoELXAaR2vEndqNsJkM2BpIyoqrp122q
GudjsjLwb8We6OeFVJxMT5DVoqXQgPXrGEDlv/GQ8d97u+BM0tGwC1foM8+qdojX
bRHgK1zAIhv2MXh8RpRTD53BZp3p5IMPAGJuKefm9UBb1zreahC7Qw6xnD9lcpj8
Tml3ZJPM8/iEiKCRrbAXYFUrw+sX1E6vBqsEnROjLDtGC2+AmSy8feLGckBWltqW
hxUa0n+vsyWvShwL5bKAEeMM6qY8ZPfGvEmvBaxqRFAryIBYbzMEcCdSQKSL+wFe
xmDBujeNPMlQdtYLg4o51HDJV+nvmjcOTDaUk1DjCU//vVcPgM5FDD4D7XICiF3x
l06Mdgpc8NzzuQmttnRXvCECz3i1jZvPdWIp8I117ajvABGL+Baraeb2pa9aXjZr
u4SMZ3WjKRpP5xNA9WX2PW4HUEM9yLT94S/uZsvI5fBzQZp/bbhBPp712lNSeXb0
yjHfxSMHd3ERg87SeXLUac/IEV03BBRyH2/9I7Vr/kG0Mgt8vGLZvXxNRvC6BEWs
JAE91hTrpuwDTOPI3/reDykZowAK+/ld5sSDlxHFFBfNCXcDv/b75olP5K5sps6m
Ehm2nOJpCAlDQCxocOhCD6a6LCmf4Dcl0AOEe5Lj71rmPi82CL9a+lZvdY35hN4Q
7lmOErXaFR9gg0Ry8BYvo3P7NyOf8X3hEBUai/QZWkrMYE457YZ/i+QMwVi/2yrC
WrK1WTpSQm6l6R02w/zxYWCkX5SLIIc4o8QNZCPvi+t9LIOvdlltZCQ/0ucCUQC/
noEhx3cgbn+9OF/iMBzrg7xQuOrwkynxP2b8cANQ8PRHUiFiDVxKCEnFxvHX+ZTR
84xTCpWhSl1wL0hR2t3uTspkQBl30AU630qP0dPSlpjGgDzqSNcpP0Pqymiyxwxq
uOjFfvqwPReWqNscWRwuM6sQ7T654HnfelDrB2LWb/UY197I/LhncLjSYgxt+7NT
b+N7qrbx8QdgY7OOFU3megl2liWhCqSDvs74yn27/FxMABt0nGJPcZaWulUu6hsy
1+aQWZgdoPt3kPFU1PNJXyAKEqPX/rXcpu39yWPNbbYvIEfb4Z3gQTMrtufq7gjJ
8sHWKkeLyBH7zAgVbn8WUZI8pRi/18bD1GDqN3jeGgeXZH8+mhYR7NhV0fap2F1s
sWwemRpPx2zxD52rIvAok286mBUl0UPiwoq8UymWjxnTNtP+JbJGIWyeKTVH8sGD
r+S08Et8JL93i0Rus7r4yp5sCZS46ecgC+avLAxXshM70/ydMJi2insNzfUi1la2
wL3R1SxckJ0vqTOU6f9yf50AGKnIp/KSDgUbX3X0bZG4Zd50S+MulV2Y4gkk4Sc3
w3yyT8+7HekOaozNCU17n8zhTe8qLeE30ux659rFi9LATLAPVscjrzd5PeD2xxzP
eSvC/jy2S6z9U+gLxwI6fSzy2jQCUq7dmlpBhKJT+7JHmqv7r+HxyCDaRubu1rLW
6DvcGpUIFDFXsO5Vdzc495vaJqZ3kfUS9RZFM3c58Mds3mGe4FXuhpvFlxVwPvIr
WTBMnfRL+SP498XKOmn+3wzMzcnuVIP26NOReC4VFRcgpz6avp5/iSMOG0pDVqiA
dLbCQsyjhcckPfOVIxXBcCM/LdqGkrvml381y4RrgZ7C2rVHzv3s3lqU/1ZubUlx
6pJkIaI+/bmGesvD+6lnw7XP3RH3NWSO1d8Cy4tV9ONNL6jzcqTMSMXBYtf5LeZ1
Pz0yg/UM0/QxAoV51Zf7EqnZ4Nuuk/51Tx7jUyljM9UaJ7h2JR50tE1wOzAk2F4t
HWrj7Om6yQuEy9uZAjhyoQ/OP9vORnR1UD24sh5Yqfg907Ie/+bjLJrXdicf3H4K
aZZQsK1w3FfjELxHnfcE35cBHWdxO1eSQH7boLe4ndCywQKSfoloVKsAnG1/WQCu
1aFYFu/GldFxm59k8Bbt+sTe90zzNnhMcT2X9MXCWkngdOxzePujYG79MOQ0XDEv
aibg3xypOc/yHbN9qLG9+FX/+P6GeCtiwGEkxXYuzC+XugZ11Pfl3XsK06N+bI+Q
2u5hbae7F1lYvVK7T9tXj2e/Kzn6qSDRLA+IzJzF13GZwaniOcRDUQ7toMmA5iCM
FywOLAAMEwlJpKc8yTJclrcgxgXFiBL8SLXDCH+NDBp3yv1sGwLMQFGDPO0d2SQC
coppoxYrcIWdtyBT+fB0wxC50Ag4u4BLHadodp3aiZS1/eIBC3a/1xTmldbHKedq
fS6bHmGD15Hh68+mtI8YtUp9E71MTy5G4JtTV60r+R9P416I907AonmtpKGqrUhg
CCDi7cipB42LEDhF5fce1LLuPCFXXY9yFsRvYta0Y9f6shvO5n6CPDZ7/ZkEeQtS
J1zKtxhSU2yHJF2pj1cw5lrmBiDA4B7sfQZ7CorHuNI7JhYr+3b1RPZ86R0xbayb
ivBQR+ensgK1LidFRi7t9xtSfdjw8L9TRcthBBzb9+QbzH7xc+f2kGV2nxFpELfM
9SP5bg3ln226DZU0QAq2GIoS3TObnbw8XCqUxFP7L082vWtzGsWKq8a/mTb2yxAW
IGjAaddoDqOAnRjGG2EmnmNpFSJhuI93265KRBjiOwt0MsEkxSYswCM+ItSXZ4Bx
dUzZiY7u4E+tMxYWGXW9HdPjH3nwbuX1sHFK7biwGtRwoFaGCaXthSCwAR+I6S7s
h+ZMiJgU0EADZl0T6O669lK+l33tHH7cbXTrvjakprFywvQ/rkW6ydYnqv1hkTmM
xx+D0vf9+7flYPg2fDAbami4G4CRluZ2HpPOkUXGl7N8SXMbt1ln3khnNf5PUITt
mPdaykvLQAdXQoG2z1SXxH1ngsIF0vN5MSx5FCzkxiQErvRWmr4UI3BpPteYU/Il
NyXyq50Qy8j75Sh9uW0rAiBPNjfrYFUVnfT6bIH5ZJiDIKe8hnb89eJ+RCxS3Shy
PIHUnjjlEnyju9teflgvdoBS+GQyfswhjXvJGmxmDwSq4hbc9cLiqgVswb+M0aO4
CPzJn0ld+xzl9oj8q8TM7JRMgomprnmgRmaYotraG/tUu1blm43A/+aERR6bqYck
yOduMfi7fzoM5VOXN02KAu0BQnXPzfx4v0bFzYGjsmkEQVv8FMG/ZmqE75I03DwB
FyaYB4eo2tF10h2kdr0lsJeS3E5shKGLip5HKC4W6seAk7pXXECf+W13IJfggE2d
Dsv/VpL5X05uqcEpolD4QPC6Aig9wrtWQl7EP1+AOiCBjxOKMlBXA/7phe/PAkAW
Fg74/JZdlQQZvj7ERLBC/zgflLepcX1HRPPE/Id7AvJrsk7u4aAzkgcMHZAS4MUi
nIlZaPG3h/MUyrT1Qv/Aq0/6TjT/4f17hfp3ksyzkrKauasp10UNgs3BNiJZvYV7
GtP/lqI7SR6DrJY10UayPnlieiBEj9xOv0e+zdZ0TiHF27mDbZWMxrVrWAU8ZVff
Dj701lHtsiX2scAqfu85+ahZjHjAw+8opHJb4BGqcSd28UY/p14m6CwmSSeexvRS
8btLY4jRYGa6s7/nq072UvGX93vT2lJwWOCIvqvwe2Mt0dytFrgCWx3Adq5CUbk3
hLtQYLEUImvd/0PjpGTRhzs1Va9c0N8lB7I7fWPTcNJe29qEye+qh5fUzUK6J8t3
ncLhtU0BlcGN/d2Bi+fSJ12EhxC5CIWhdCEwqVNKiuiD5d2RcEnm9IBGTL98+fci
7U5OtUWLNG/NMj66MIsZ5xSPII8OrQDHkD4SDAdXEgafq7elPyxCf7ppl6GVMXSd
EaqWw+65cvkajWFOCmgSApNKPqn/hsZZU4TV/1saSpZTL7sq2THgdXsD2LcfZGA4
DwZn+YQYXZPAYti6xVpMdDtCfikkwcOkbEEORQk0Nn02HxMhAbLqwoOwVt7vh+v2
Hag6TxPvDvRkKQSNJylII2468xlh20PjTlPsZZE6zSElXImr1IUsQKct+I9FosBM
N7RJGB+a+xwdnGoR64ZeqQh/iWiTtF5A7TonpxHXbZLBYHvKTnoGla06IP5vWkQp
ntS6/PfZqbn0I+7vsxv8rRfIbrWOnbGZanOH/t0tNb5n5FtIn3+pbt3N/kk2doMD
Dh4SbuWbNPR5ENyJ4Bt++zMGhhWEtCj+AtA9+Rzz26yOUlWnRB65Uz7fcHfd4wke
/Wci7rCK+s/YqhtyZ2NJZStq+1Of6jrKhZdAQt0JnEpD3c0h5yE3I1lWcqwGeOb8
aMnvNC/JUNbgVz/l6w0Pxubzdx5PVPs5MaQcOo0pJZUgQrXVqPZ0eYwpgKjn4RgI
6cMT35RQuObMV1VVm5QdlGWUo6ABn69KqNJc1op+tQJecYvtFDWynscJbNGAXyiz
167p5nspUMO8LlJSwGp4KA2+FWBsrQc+D248pquIhDj2ZWISVec0hayxHSo4MQPq
Krs6ZXsKvhT6y7KOxhzHsPEpn2JFAzZsRFePv+iS8YWihU7C73fQ3DnLnS8vY61F
IfmWb+XshzD6ATaiDHovCu9ZPgM2trJr/1TA83i77VebMMdiT1P7GsEiIpVX464t
DmZfBZMH9M6jTdqxgn1LRR6KR4/2CtqwX+K3hm8FPWBSz3UbtM0sFlceAgZSVDOe
vCuv1ZztlwtK9fl1bYJgfxLMPCPRzA5qklCNP+eteyw/dBf4FyP5HaiVrWJjesHP
3Ct9HacmHci+0QQ8Wr7xIEtm2H6WREyulpC7fg5Jzr7MSGjT9HfYKDZoYJWJCnJ/
OinHc352px0VwHle2u5UVuRqh7spyWhI7e/DZ+8V1sLPa5gl4J7S5aBolmM8xk5r
NoG0iO34I5aDxIc3a8GTsokMJtddKtFCVHKPzKpX+wSvPNtM6vQ92HRGAsYT4WRa
z7gqFHZY0mvJ5rlYosmDB1HFFfruIg2k1Eaa+rovbKnj0juf+NGD3ze+bZ9ReYL6
QEG0Htc5iua0D37PauIHMDzU6bxlZZK9s/te0wlxXIVR3+5stW5LtQVhQsknpOF0
PPX+K3BXgS9pgmpgArRFFlZs0F7LV4D6X7QUBaMnOdgv0rAR3/uZbOXQXvwasxIA
TvMT0IQFL89/Ed5xbZtrxePRscDoMY1xq1eCs8Esh+cZR+KBa23NX3aGwJ0aVLx2
aBvvm4dLs8RFXdvnpL2AziCJi1r+dRRM7ncMtUjxSmb+1PJevw7wKp/ojfyLV02Q
AxOt0GgYyqnlRvl00gNKCDvfDRzl3+DzLRLzBUctwrFtvUZR+f8DIliPbw2nma1Z
jp0sedQq+AkjTm+//D8O4BmU2Zq7TyGIurTOCf6nI9Rh20tvecZxe3KWBh7QbH2M
B68DbcANLUT2we5/vpbJ9Nyc7ecIvMvc3btLVCI7ieZCq5naQlIadKT6BmpgAmC7
jexl3L8iW9WW2RAyGCzif4MVKeYNBJjx3HHlKvlHe+Oe1C3nbhogP2hCsV3AVbXd
+bRJO+mXdUyWUthpwVLWSIpHailedppj4s98HIuRQ0BcXAvsG9OheY54QfEphRIM
zdxmk/dR7OfwGnId1a6C0W3k39FLi4EMShBMOIIFr+jlfVL2ty8q+vX0DJSMAPk/
kHgSppChgc5SAIkbLaPTklpmQJ1Mkqi+NXxzh4EpO68NamDuv8t9mszI22ZCMm7T
tpXso5AC/3f7NyooEauWWB0DV1DlMfmzfrEHeCKEFXe4lk+PR7pFJnRvILxMyNhx
KX23R4UVoHcIw8ZSV5pNlnWpFqKWWiW31xUddYa+zMKYL9Yph38kUZAmcfI47zjj
pQSjJZmfia/ih/FagVX6H0Or7BlKothNhZjiTVT2qwYXCMJiMFfrkDAAdTs8Go8v
temOUsEP+Z9Vxfm9Iv0UwBaDCj/PyjMpDitwg5Zrxosf1YGYXorIJmbLPvhYdFJ1
EvfjsU9XNQwohAs8huDShtZFsXSYBUxN4BU6HvUQOrcy8HUFzjMiOejP0c4El8MH
Akg0Q6rlR8MjP69UR/JcwHi5Ysry2bUGnUQy6LEb3bV9XlftYIZT33XKnj4oNKRu
BAf7M2976fwZormIi4SQl4EZFsm142xocvj0jN5ZOLRhPDCHA5NjVWdHOMuUTPCu
OGNrTSnyCN1W9TeQD9G+FXmCcT9xcnFisotGnyjuLmbP2OL4M3OIPZle4KpiBhyh
sUy5p22xxeQ4ZG2QWCwYyEMAV1zTHmU8VBLGmyoyrbZ6/4ygsSnr5EPZUyURjVqU
sAZLeSF2QHAlWwgU6V8h22OUfKXcwfEOz/1z+VcaGCbdER4f6wOS/Txnyj/JNlP1
7MKrBk/bM98Vs2eaHtiFYTEQspO6gpG8hcQCJ3r2tsNGizqS8riXLtogLX7m3yQp
pZ776zoUfgCa3KZwGIzrjIZQVnDmSZC1SJxJWHm8U+a+tTOL/qJn4BGAqb/yl16f
RT3xdeOOuNlZLXarcah0GOmWvBIEXlrUH+hJL2yabI7M9E7ZVSJ4mTDHUCvl9kkS
ZjhxpbEKpOGNcDiz+QwCd0DfreehuoRiswvSsuheKAGcbEyxRBr3AOU//DVy3V1R
MS6I7ocR8qlVNmJy89mBRiSYC0+CxoNBTJnd2Vz8vMH35q0I81muN/J0QCTdHMoY
4eIrqXqI6g0vn/n4iP6dydqO3ZscFmOvaaiMrTtK6jqLm2NlYlTRNJKs3HMewOQa
CEXsQsUAppYhrJvOb1gQksqonF3om4ThfS/QeT/pr4Mxylaqe1i0O31S13hfD8OM
jg3+CZCxeR7zuJ63fio9MIZKGseJi2rerpkxcAcc3JDkT5BA4gjlx5GHbbnWm5ZJ
J+CoqBtgQFQ85EatiqnyOVbyH/L4+znIVfskpHP8ADoGOLj15f5rPt8i1K6gGYxt
FI7frmXnU1BKJB3vR+DePJZHsgzdDJziIPlunCbe+xHO36Fm3yOgrCGMGr5UxRkq
KePBjWzroYyO2gRO6njVOOUz6Nr3BUBfT7c3oKKjOouk3m6JkGp2/zP5gRE9n5hi
tuk1WoQ9+AMxGCzYoFIJ5kSOnrTpx0ZbwEL87qo8lkjiA5eDIZBQRZ5gDAYrv+/4
cy96tdYqaIUHv1WOc6GBPnN8bw+WTsY5iKi5OQWohZ5/KsEVDhF/U6PBsF23yxVK
Onh3ObgSgO32j3ZXVe1K3/QpnC27UrDBxnyudOl+/iO0W+SKYAVk5vfcBKf/s0IG
B/9eyAN4ukeQkGH4O/H/EmdIqgJfh6OWu2hsXdKRaAL39YzIvCXa49WsipdSUwya
tGUgkUlSAO3WgwlKMbthKYB36Cz5o0IBtT+lnbqX+XyiDLsrjXuh21LgIPjaWgsD
wnqflrH1ozUgfVNzwx3maJpXZWmFX1BucXBzYJjEwY6HQoD6HQVLqlZF2JEZZ2Y6
3rNi07u6QiKMfsEUpIO12orhJoIbwfQqicPwDN98qM+n3prtPdO3nVJdqn5gCsnU
3ESNwqAsGSSuQKt4TnJRZd2/GMwRxdIB/5aoPv9TAZISqQImI6Si8HHCJqEYwVh3
gMPbFTntazSNIB7FQpAoZZirNvjoznCfydXdelb+SgL8YtbKmhxvhom9LoH34wlk
K1UfUrCB2Vpa8+P2FnxtY2iNgAUFzu4RNqhq8kirJRhTw0jVX4ADUv96tnkZJfOh
Ixn59xKS+fQTQBQWUrC1xEi+CeYksl4+qz0CRxoazp273X9fLr+IlHXHC75NLndC
cUypWhiK+KprjppjqAblhrfH5zlkuo5+3CDPQVP2JtfNnw3UtNCDEznvkJ6jKCAI
TzfC0WmYYQHTH+W4b+sSXb8Mf2d5i9R1Tn6A5WLS/EpLHMKM/VT97aDsYzgUXN4O
bTQ1iqgaLnu/d7iO9q6YrKmHADL9+GeFjYgaw+BMEehippQvt2/blOK3v6C9Jd5M
ePm5V+aedJBQ+w9s39cGWq45d8lARbUBQ48weABIeoSO3toVgFAFljuVHd/RGNtW
Iadph/esd3GCo5+icHzlEmK3SPmn9TXN7kxt76qQ8c/6int+zU5uOzHYxPGqenC3
hcP/a9mdrb+lLWYSOirvFew14aWvNVq25a47YdXOG0jrDeg4tycgiroxJZsh8Mk7
3CTmQLcCLcQoeMuE69Rb7awqe36BI9bqDg0lddxL5Z2S2fzlAsIzY2jukFCGGXpP
DVOsVnYAt+wLbHScMDO9UeZxWW/qG9l87vdeDBeC4+27s7S4j6s9xEnpKImxcOgR
j1LuXqfPygNn7jJLkkYpZ/mIfPRPq8tlsWOCXGebcGdbYPJ/TT3/5Bj5OZAQcS/q
NZoAJVhbU7CNbZfvRT/uihmDq+PrhCBro0qQA1tVUIwi0sXyYXl7vnRTjqAKRZsM
IUokcQf9AokZLkaqlRiFBkaLswxmKv0+k6eE+CVeR6po0rLmxq9ZHhY+PDYV6qAe
aQrfivfoOBXZRv3o53OC9Qh3SCXQHSvFF6pLeaYZISnorqy/DUQY8MqXeAWTlczT
zv5bFmyGp4DuLG7roYKqa7/dWg5GZswja43Ce8tRZWDVkp10+sNswkz559fJwGRN
j2wbWdhZO6cmIQPWAohY0tWCzOnKQjWuJSeY4Q/33fGbsaVCazlRnN+suRKVRjPq
J01nvJJlKPGz1PLylb4vKEGcPEq8mdAmc1E4ZnmHun7h8M2Ee85N1k7Q25giuq1c
BEwZsIUHCvRjJGD9JkqzExx4asrH4UIeEIr76EBDjzjQ3/hD32T6CKJctC9c1Q8C
qUHxS7vrdIMiulrtH1N1kerjbgAVB9rm+ACSqoppw8MvQlM14naHPT7Y+9YzUwn7
O1NXPQYk/FWBiScwYkot3rMoVkai3oIbkP1fL+05hJ29FCOAJWBCmY+FqV1cD0cC
c1xVffQrc22K/ubyL+Hw9jIJq/MG1mW7MJiF7AKR7vF+vwTDViLfXl8GQfvxqyCw
gNnPJ+/NWFDyJAEipAGYSUm8yYkLOI+u0AjlGt2FsAvWVHJ4laYWMfna86ad4/DA
Xc18PaFcnJAYhdWKOhBa0Y3mUQJi1sCTHKQSYVoP4CRGsmCB3kK2mvdNuCK5THuw
1+JTZKlc+BOMJpGqDP4xNkDl+MgPmSopcqoAS/BzYUhI8WsiWBTQOFpvO0ETEHFt
A51U+TCh/U1ZDFG3ABrxsElTP7J7JkqFrFDPoiavNZsHbnhLWo4kDhuKeCPtpn9k
kmNdWwswY8Kql+yOSqn2PgE3AwjFXS/WdYfa8gvKN31JggjuIZq/BXPauYhTjjPJ
Qr8S9nOBc5e+UO8t3M6nmZpLFHCHWd5A78f+m5x13IrRnQoPk4i1vGVpk8lapm2m
5LfU2SxDovnHMhCKc7WzgGKzUxHpwejWiRusxVjxx1C6t54Ty0DcgYxBlX7rnkhL
o6jnvaFjFZgkdEW6SL4tFqFKOuuMFabAV/Lrb2C1ChLoKnRbl3YRv4p+C0+4Y1W2
EXiSBESb5icYqRgRrBqVZZ0QiI2Wno8cxCqw7qvig+alSnyyIYBHDOJ1rcLT/5tP
R4UJNncq0Awy28qUEG3Qy7y0Fi4jmQDajCVi72LD1unOVAFVff35C8ddo5eq3Lpi
K9EofqR5svorxQGuttDIeqAzSZycnN2BOyEoDUD0cEL86oU34OGatLxtFzgTLaHa
GFGRAc+MljipukYCOoA8COlguhn3BpO+wajuCFaQHkQNdvfRYh25oLw4x34INVWQ
g4Lhbmrx7zMvFddZFCRdCKocoL5IRjIEYloiTlUTO8y8ZMQe7SCOWEf+2yqtRKXY
I7iqQDq0H5iPocSsXBF545SM2McvLQveIVlHN2a1KJlYDn/Ipt8RhJ/A43J0I3Ph
FOHT4LvOd3XaVsjuodOOirOHzOga/qBEn2jqR24g0hMiRsndoZnxFAHo5IXtF3DP
Qc76H8wRUsAFzWTzhiALPG6ri8aa/0yWV+83Epkov4OoMYq8S5C154IC8Xa4VQba
kX6X8uc/FxL0yqC528570PLXVNPvXVDoV4xcTYPS3nU+XfsV54Sq7PgtCDgTRSCo
t46oAgSOGKQtwKZJUpL9HuY95txalNhsb9vew+8oX0RL2EoNL2BRngorZ1dnvRIo
leMaypBFmOPF6jG04fSdjqcdzecGh1NW4lCvMMf6djfVrfcc6YFQCTRIm6Nda7I/
lXzMEUF4uGBcGM1OPP2MktQ7CqAuWQ8o1g70VOPcA/3HwXXdb0Rf7J0axftCrDt8
VEpwSS9hUfvEpsKaJrn9QvLIsPW3nR1U7rdxhIQZo2Gxwpmgtbcorja1i/47GeSq
xXQdhvvNiX71v7WnXwKjkbsi4+hKZ7QWCjtb/0VPYKBcO4wk+fKyrEzWmRCuKbv3
XvNNrgHAXHR+iHrJCCDKffD7itGzgliabtAWCMlTisxxXdtkp1G+2mCOw34MMWYz
hUg9YjQs0LJyTAf4jYrfrjD5J2lr9GsnU8GI6zxHP/QwYrZDa5B+3LbuqoNvOaXG
qt4kPCNx+OFF2ZTgQg0v+NzlBYYkMy+0sewH2NvRc/oFSi6oNyODZVxTH3Alzywc
fTBa8nfpirWVH3RNUwVGsI2JKtnVbfvyowSxQ3H4uBcm9umTccB9dzn1r1txS9ry
n855IU2GSL+1ihe91XvQDfa49tMIEe2OfGvCPg2pBiYI/4GzGi4ikTh+9qrBPE2u
cWwSAvrFB6CD1N0C4Psy8259UPh3Gz1LTCwLbUHSXr1RgsgarXXfwi3hCXtvhwCd
CIXdyuEFk4WCsK4bmTXO/VGweXCw7B7rn1CxtBZx1ZyF70qkDaxNzY5NDvggUrZ0
LMjhQKIZYdIeAY05jQBtZTn0Fux745Qzfa6iBad2UtqlarK3k5WlA4b7RCBY6GHP
KhKVU1F+7rup/MVnUXAXxuK9q46yaDgn9XNBgjpuXh2jLrlWsGXA5iruXdjtgf/c
WwEfgHBGo5CxY1eiKSUR8xy6E/zhq+9kFSUHWXJsJQsiIZNzk3GEUrp7Y/PazK0h
TIPiPR1UvqDoYi1ZXEajvHarWfLb3E+Gqdoxqu4oUj/ZuYSGFaN37G3dcCg8bEYu
noneON+H7Io8R0MmSGOxFnlXuOQF7iXaaBYNRGlErpgA5ePiKN0XmAL5M4qfk12h
mhrhUnmxTDuFl9ccVvcQb0B0OGZvhWvy1NWERe+N7Wd5vmm155wEh70eZDhIl6u5
VcP8ZJE5gwGC7O+G3izKgZRDihBXeRxVa3lrbzwrLwdjVj2AZzCNn2DMmCROyG2e
2n0ckZLo/GMsmr0Ij5wTjBSwKzQ4ApHL3R7bsc973QLZtNiILdAyHXwEB5zkx1uu
ErC7bq8Sr0f1rul2+HsJwLL7Uw4AQAgT6W0jvm1w6WcUhfZyf3e/CALS4sTmoTTT
aE9wUVUjwKWLoxnq6FK0mZTf8stYBpX94wh1DFl+dmYEPupTSSjCjvldmeimtHrw
9K3AEx1o7R8OI8XPwKm+DwymxJz9s1hOi+gTR913KWylzs3RcFgPr62U4eEhNR9x
aHV9NCn9GkO13fW9gHs3kWudOMqhzTNi4rsUZRbrldviFXQWo46DFUQ58Upst7Sv
idkeuBzsh2QiXIKj4v2dnxcLflTgNLhrrW/2Ulq2A3RHC5VZHrcjLCZC0GuVozGc
6IjaQRdvHnrQ8Sa39ApVYeyA4xHbj4twVJ6TmmJ8rOMS434REXSZPNF0m06iwoq7
jjYIiaM4RbyrLUuzybb/pGd3ROvQWdTQvWRmfYd2WCON+khIhd3zxOKmdZ1ILiWd
OBbyVy+n8Dd8fMHt8NnXUChAOPOoaxED6pRJh4MPIQ2zNye0pIv9bvW0SF3p4ZM9
0ZOKT4B0PhYWV7rWLFQ3YGBFpA+IFtsyRl6XAnZ+db1QwAxqOy/JLq/Zhm2Hk1eB
voemOwV+nXjEn1I++b7UVlghrYZetPDl7zTssrzJJQKYfGgH28N8j9+xeJS8Yv4W
GR9k4zw/52iHdXy5bRIo9wMI/zuDrrEgBx8gsen+tGcbNqb53tezmkNh1D4vJNm6
O+wLK8QDphKelHF32QT+3CymDu0npnZug1Cb5WI+CZ7Im39fLZpjcYT3sSMPi0Fz
OZwNj44hKxX39RJ/AXNvvkcFJqFBxKkogGULWUCSBjQKab7lEjOrhNJgduRQyJPG
536HRJ13WZXiVxn0nSVNON2l7goiNUs9u+9hvHNBo+bTGbe06Zppwlh1LBMwXV7Z
Lu7D94AZ9EMy161HM+gd1b/B43gl0ZGtSUoqymWgxbowIZOthtw6uaomIFvMYis5
g8fk+JVa++c6rpj3JKD4Iz9OhfeqKq94nbJ3oqZ+gcbc3hJPPntD4AUp93v7wA/g
taJDVi99CDJA/zuwBf3FmsHPLFY1mU+KkVl4v5cU1r54/eILWl3cduh1RkS1FAGZ
3E0CzX0bCc/JE0v45pkOFSp4wrU4PvRa7zyleAnu5gKnGLMJtzqjkSru3c5/fJvK
/3rFvzFizd4sHKvjmw6db4pqylDHlzgSybg8T4ZwqTFT5wqwXe2klKzE7HQg3cdz
CTRJ7hn1kTFuiYe8u2xEAYpSy260ziOV7ABKMxRLu2+U0ga4jk9nnuXRDMvbADIL
EFaCssO7op9La+pk2fublN0+Abcj35E115UfofptVP4ocu4X1UEum7WRw7YRUV/m
ZsXKQm7f7Bc9iDp1yCcL2v4K6WVHLrl/2s2IY04A2cHWdyn+5eleppjKXQda3Qkg
TyS+vXS06oI7i4GGg1BKtTz7G7jBNtoSGR2C5igJaVpKvYof5rFx4JP0rrl5bmve
nDvjGZbzSumMmMH1as4O7avt/BK19lFlPvI93pdMtKT4I528+U+qzIf2W53E9KFC
wV7PRl7JFqDOB7kJU3qP3n8KCjM8M9P9pGeCyc0yTLrT3MvnUyiVq+wRll5nBD2F
VJD24yzBYqIbMr2PMKNI8QPlUDiY4sPWMY7mUC8GfWiziXffPNDu6CyUGmQqSZSS
F02cXXAUXknCzOGQKGeBJ1BeJeSboX5lYLE5WGXBLH0QQ7+OO1080iacW67YVTk5
tDQPtu4IhJoOK15jRcg2DyxT53sQQ2lE5Xh8jAKX6iOr5ddQ/Wc1YSs4B63ayYlx
XWquUoNP4h3qEa0q58v4P1vJwNNdeBpwQqj/eKxMUZ6cn03bOq3U9mF+ytz/zvEz
X84GUYAbpiXrBLXKnW/KMFvPKTl3aB/wdVSx/9nOs1M1uHHvLgIMQZEv7SwywXHd
rJZ102hFeJpxBqknVqMhfyY7t/WjnMJp0/sVglk5B06v4ViToYvFWb58SY5v0myr
Uvv9cy5VyklY2uLlIk2bzqGkrCChM2jV31zH17f7bEN4Y09FMXMEeZUWprXjDgqk
lB0sv4QlRDQbfy2RYbMNSsIfxwKvgnzEaJvVSD6qKjJ1KFYfLbY16svP41ZFGanJ
5ABGhnjJ680uf+DsgjbT2tojxyG5eXZcF0LvSgUncLUby7ZaKsAzEwm2lRVDODZy
vNBPh+rNVf+yEC+fLIsEo/RsdY/+DTA0aihujfVVYmG+U7DlqER9ImPnXUTQ1/BD
/FJN22AK0sUmNNYr8eqX0LNFuF1oao0YB+K433C/tnBRNob4U7X1TnLKfJQIbqOF
I20cOKBtpYSS7cUjMNCyNLkrQehNq2mfjmr4Z226nckgNQnRCMab3UCAr6lkveb5
f/Rx5BFXHr8PhJ1toSm/Qp/HsZ5eE+YNBMbifz2Y7Qm3uNyfSGTQB3QK4XnQY4CF
WYY8Zo4OyXQncSBa/vkpSbXJTi+DGHhFxMQTvXk+cGuI5j9NEeOARL/wXdkzl0p9
VENw0o93Y9eP06wek+R/CqYUIQePYKCmGS4ref01XlhBlg91cFbSb8EJyS5Eq64Y
389IHS0+byWyrSSOuZCX/1jvux730zeCgGJessmNyXod3urRbSHUwzOodwLW1COW
h4rwZtLLzcb6Ybz/2w0Ff83VTS436ZHeCjouI3JhiP5MGNGrTH9EpvHytZdfuO/S
Z9Hpa9dpcl3bvvhRB4UYb/jREVdZ6M7dAYFlsZ3UNZVXComzdMYGX7hA7Rxc1qmm
q84HReZQrOMMVe35yHEyIt43K23zYCJoU9gZVoj+ksyIosUR7id5TpdSHstSI77m
gv2+j26ipiZzCJa96elVXrvJf3Zhm3Y42lKpRa5zGhYAyNSK/brZLAxlGAVy1tfu
xJgeWt+5vri69UpiYb0UfU4+uV0O89MVDfxfRWqaY24mNqpuUdWRlx8eo/0gYdSw
sbM0vTBns12QFSmhAs9lph2sRv6dDQ9l2roj6aTS3FnYnLPXatmn9EaQ0Mcqye6d
sEg81U/543jVw0Cviny3pcsft4ARoa+tqVhASSxFmX6URL5Lu/pb0VtgFn/9eJuN
i73qNVe2aLllzBXdnDFRWTOEsOdk50DNwSUq5Bc54ba/vXOUKO9dmULYfU8KHj1i
VBwGCzKLT5AUsxWKXDfCY0343a/6fOR27MZK3zOGqSIECoJXJ2k0CSfFhEEwyKU/
v56dYrVo81e6PijYtmMUSsk0SbwU1tX6tZDVHvuITJoPRZEm04xUM9cTLkO/WVNg
IFEYQI1upmcREGj7F3PYM4KfbDnh4tiWCMEi0HXY3xZ3vp2H1VdI3yu2iY1aXEK7
xvRc6fkwDHSq8vp9Znwh/gslAaUv71bbrT39fl3cH8Zw8Fi5JGyPp9BZRbwlKjTi
dRXVe6E2xsBoJvyNQ9KXWlcfxKElpcAMkzbDGEKHN/OdsgiFskY8awuJWhw9ohmC
VDzcUiExe4X+LmY1y0bFTcbCDt0B1WSh3SEzRqlxUf/OWHX0fWjAruRYb/B5j4QS
depXt4vE0SYeWSb+GmNSUNaXovwjpqVIpxHh8SojvtgM6VmGTajZa1MDHeJJ688h
O6BwIUBUJqbDpQ7u9DYNaXq+EAiR2++cg9cCrbUje7MUwja4DXE4zOWmTTZo6G9Z
iq7L0DqoJ/gR9Ev4LsmtyPOW/oWpyK4AG50FqVmqzPWzvjmdVXzIxIRRLC4+86pT
x2X4+Mrfmp6LXIsWj+ebz9cKU+cYN03+LozqucOhDhnLTAU9qDXuNwbh4BrgdXaR
oCD1lSVC/0LEk3h0yumsJPkLX+wBMMH869Epj6dPxEAtyrYNduSyCGE86170s/pC
9qHUMqMwdndFvxhtxSEYBK5Rm1+XU8JH406P91d1orlNBcvQMqBoS6SQILRfLwGH
GuT74AY7uobcsE7j5Z2cMLGjTr7y7szAOn5e2l0wC/HWRmS4TfnQrccYocFpEkQp
KzVn4jzp1xXpyOBKER3xoBvU1KtLamRhD2ya2NjcPCFDuqul2e/UE4F1sciciUcX
B6ZkqO+Ul/fFjON+slxB8LoVmL+vN48VTRHGN/knxBEXHVBytYhxBNY85mPoC/jN
QvBGBSqhmaLxoHRbglCMPbE1JSBhswi+Fo9t3n8YF4I2O7rHraXyxDP6t72ttzke
lwvkFdTYLd2aJR3Deos6aoReRbAL+P1CC9FgqfCIMPL9hQARYNKwWQqXEqSgBOrx
iTVDSLRAO6AYIILXBxpdc5iylKxsasgQoqWOuDM2gJHFCn7WX3abtTI/52aXzk48
CCoZdgxs5/1eQaBh+ike4v9RTEIPWmM8xoW4U5UNd993MIWNFtVLAweMXcYsANkt
AOMcxzHzJGp/tDcV+9gKUZzpBE78hsjsRrcplQ4Mb0Qs6joMrPcRkIqGYh/wqTkn
82T8mTRJGQKUlSX9LiT17qbuEulLDz1d7ubvVP1GXQUL9vGZvqz+fZ0y4VFy5p9U
CgFlsJigpIRlSXP/ONsBxXfjgVqF/7+b3j/W63Ru2MxzmdxeoRgUMvwuD8s/e2dU
vx7NrNcyLib4xI9ZX8LNpz2BcoPIjBYVZGqADfNdknx+WDu0hI1VNDzSCz368YOf
nXG0g77wyUfRsb0wxCgPZk0pzPAexWYY1G1KGfI3s+AQsjIMJ/ys4SfLlj1HU+tQ
rq/2ZL3zYjM3EI6fPbVvIDtLjeLP+K5cU4XzVd52yytquK0FwCun3pPLWGxRVjD2
9TW93z5661/0eRf2FlLoqNrLd7CcXuNWct8ikmXcMAYFa7fkcTlKPry2DgKsG6UT
U125PiK3PPzRAtC9nT8VurJ5nXX/NOb4q5JXisaCQfAgW86PpWBSlYHhOw1qfHBs
QniCNdXP6z3gVUWZIG3aTCI+m/GQt5LoRlQDLw+nAoGLaXb4gTirga8TCGMw9Lrj
INJYlKq2l852P6zmK8hG6LZ3xo7d4Cu7d95aYB6J8ZkT382BK366t34PcYvVvo9R
jOsVAYjUVf6Mz3KjCCg6j9V2eZLgK3ZZ4nALy1wNmroBbCDL8/iOzAloPqTiYx/1
J8dDnIpO6e9iSWwDuWZ9lpao68/zsKlN9VpVPZpzDZdK8iRHYPdmOFFBVl1b8Rg8
xvjDFw4VVKhrBInj3BxbMYoJbpSofxuBmMH9AHXBKyd5G8ZWeTchBpM5Y3jmI9AT
sFVCUG4NHw7RqM77+azQDbrUH/Yot0SyBzxzmnkBxxXVcFcHJhZgOLX9BrKfTV84
rqA6QzT1ZV9H32GlvFZyQUmBjhaIaaUgfT1jTzkxCOs2hUYrAcuYuq7FNz5pn/Eh
Z670yyg8GWXnDJrPehGy6Q8Qp44h+d+hsMdfuydGuW+tq4DENLZ39vdmwYA8GeMy
Zfg7nRDO3Rb1IHJQOkdM0DU/t+3N+xrB5joUBB0pzSS4Dw4u16EGOkSrweaIwSWY
My1gCIbkcxK1zCNgOzygmnfCPTb6yqyl2Vb75MUh080U6roan0FVuu4YeOQns/LE
ez6hQwIEnJC85c+ceGs2ugfKixgqx4Ib9kgv/Sf7eWfU9vP93UeEM6ckiD675awL
zhzAZwpdJTI7c3FkGLTbLPYW034/Xzg5APUSi8i06Li4uiFply3WC8HZ5uqUMWc5
Z4mkIUA15lOP06H1AMePVUvk/2WQ8vGVi3CI2kprRG0SNbPlgiJ/fTifr5ulmSE4
mBXZSP8n5DjrSlIPOOxxcQMBrlWqzeOylOvkOsKSKi816bYdWhMCMKF+HvPKW6QM
u33jZKcMYHQgbQy8ZECBO5d7BEnWHYUfb417nZzBzfKEpGuLuz634RHkdD0FRKCx
y+Zk0sRTZzXoR0CwYmC+rgmXhZEiugluaehNYthLHvx6f16WifvNv59UBVyuFNkX
EvsSihGmiZ9DuzAY3DJeBFmlTH8RQYbgxe02IX35+TZaGNy4RXSxBRYI2tbtcX6w
BMkcFFoAlVU5/gxBznjXakOWBKB5iaZrRGw/5vvL6scYHg5UEJIEYAAs3zfQtQFt
W7JwW+9ABywoHYzdeWzMDZyrz8X9UK3qUVZ8CmfTAlgqKqICN06+2xBlmok7pwAp
BlMkKA3Y5tDbX3lXQOiCMckQcD0XsAGQd7R37JFJIgY3dWIQjLgts79JdolFs+wD
3G4w8IPLxvu1JdYDYmQA0Dk3a2tur0wLtino72jDUGP6gVY2S6A5r1UYuJ+OvU4+
wsG10PLsXqahWChMZ7dcG03ezVMrpgtz7zRDVUIpD45rquYjTxd0xrjymFIinovA
bmUmaxuAJ97DNWGyCy1mUzpnIys5Ny834nY8abXmF4AVAopIFXrgBUhwokjzzhr9
TtZ7QYxA3QAtmOFXn2SET5iMgeJiUwLj0JolnX1yLm5l2bR+6HSipz5r2MA+XVpA
keXzOi+s9hLsw0CDTDgvTJQtxXme6BAk+BoHD3ocPys3EkFlSoVDob2Q8T4vGEY6
wCf14S/yqj33lrJOcPOlLYZBF7hOGKvZxA7UgiSAUas2yT2098gwD++ocgSn/MyI
74peMDUovwABhcUX+3AZaQHoTH2pqe8Lxqc6p4rvrRZabpBTHk9jC0CybC9TN2uh
bFl0bacy2AHqWbd5F71anyCOCQTkNT9uSiZrXszHlriRV+nzwjR0vtKvkD3/R9EE
Z/d2MKkUuEed6i9Jzpk2Z7DwfoV/pXhmYyxVACvw4245THuqpjxkxHsDh2CqqP20
jen2nCNZoQLe2nh19rCy7+CZxu9Oybt/SLy6b1nMqjMiZYTPaY05RuQvFBDWIdtg
EwDHsldNNrwOUR6le7TvnWlSFVdw5LcRErTHhF1Uo19qYZZ+ese0fUfAaR3xzXbs
3Q4jckeecd1q1sZm7hAVf4rHQVkjDs427pjSzyzjCfvaaFVqjzq+VcRdONEV+Ho2
YQVvsgyNyXPz9LRJW03FK7Y0eKzXB5OtrxQVKdMDgCpiR0GCSJ9wXFrbsEhRf1o+
JKTH/qtSaeMQTNHaxbxzhNbYuJfRfLH/lt3GIUeyTVTTh5BOw/zwYzab2hpflbO1
00+g7oFnQDGPRgr0lFa1Y3QDAkHQrjjXWKSY89Bzr9hCv/C9Tphvo2HuvNVILMUB
rpLcplCkhhZTJkBsar/XHIF+XFYLOYIOAYnpi31xvsQ6kSMQ4Ncv3HcGCWQrIi1K
NY6xKk6wpP6ULpcpgxoIXcfKFVklITGTzfv9A7WR7YWR1SlmUM2ep4jMm9pttH4S
GMF5WLt43mQPDIE9vlWabTXTLFdYSGR8LZFUDO11sWiu+TduAuEXnhRFGetn1uu3
Wi7QHJWFwxB802RBB0BGJetEuPQ0y2o0QecE0Syviv/CnbBLHHIrzUC7gknimyVy
5UjjqOOSyEQRvV3Hr2rnzjQEVay1dUlHUg1SJUZSf540yP5guq7vfSEMyqIngbla
ZLdEYXJn9g7RWmfHijuDRFphB3tkKvWPixwMlIGsyOrLw2CaMCEds/Onqbl7TRwx
2BO5G4QP0SZt8NQxqLa/yQWwtOqQ2iFJljQqj4K4wnLUpk9hQuHblAmhMTVXbAXs
n6FuHiyvzKi/jov22ruq3mY3NwzZPu3CPgVXpZHYoZRuvlg0gUjW3BkmENM3d4y1
ah+Xn8FOo3c669th8Zc4Jj0lFeME4/3qNLfapKB80h/g1gEV2/wr0dpr0VatqPMa
O3Vv4J5jzAl0fbghjjJsNCVGJzxoveKK1zrJ58zh6QkAEXLvjFSGX2CNlbbWezGu
DkAlWBhhMQjOusuLX3IxxKHHnGK9GZbZmGhpn6Wdc/9H3xNSFZ6wcOaGjdF4FPd+
EixvxczvsV2VGMo0+4rAqLh/SfvkCKP7U0Fpg8zwUokcc1DiWGtJZD2vHXInA2AF
hzTUjNXcjuTO7NfgY9GT2ZjO85vB0TfgbE1hiURE5YEXigkfhhVHgEx6yD/6zqfg
0AUdayIM+UQq14wclZcLECFYwLyUMkNY7t1lHyK//EVDe78B3eiudygUOm6UGA21
QFVqwV6cX/90BdD9cQNfnT7zLjvx9BgtnQDxLtLw2tITQ4vtMFwzB/n6E6sRlouT
zGvdPGsDW79DwADRqJSH9qxPB/SFUJ6KHNKH0VjskDh9WftZwyoYO9q3ODKXRtoE
6jQVx1NNTaqYg9eKIe0dAWBlGux7uPIjT96NyZ5dDhUotsdoTExaCh8pkRF//ayi
JJ4zP9bEQHIg37ouEkt3TL2N4qo802d6aSuif9OH9Zse4XB4PJDCTZK/1ZiXuO+4
oXXFfr4dXDhg8lXLWdx3A2mjzqlQzyUMnOpK27CP4NEYD44a1PlpUWCj0cYfiSUn
qxmTQa33aWPDUObtof0sGBVGWZu66lo/a910/irrrfcjE06VEAFC5H7ZRIXmlOlO
jIUZ+VBQ9BPGQiAJZzjjDWmoNNuToZHq5pE3zrfJUz3m0hbThMlODCpWz6w50Sic
86wo3mDEOp9ezZlKW7nfjkf3gCFFSFfR9AMZteV6Ikf7YF3vk2qDdwgfT3m78orN
RSe6Z8GVYKsZuBX/QFTQE/JN9bXf01vvXk/jUMO1MxxyOYXbCj2V8tHTdLUDZ0Fk
YkXQb38fQdRW+VA4FXv9iQ6/bNr6VCjWYiiX5i+DeSafUCRZBV9I32XnQUjW7huo
ZZ51BBqrKqM5AA+MpbY86isdk3W9cPdFoiDB1x+dBB8ViwY2yRdd2tjaohijqM/s
jTAUoRiUcIJmA/YYj2X5si4fvOWMozK5CJ7hHVL4E0h0Ss5+nEG75zm/oKTQrBY1
o2jpOtn+BRaxiSe0Gb99OVXPrt9uCXp9f4RE60GNA+CQ9pb6Jiq+lYIaLAlWtCcO
0dftLZ341x7VWBYLD5m25dTw3pNvZpx0+qZmqCTPU36Y5lRB/ueQ4pwpPYxxg0TV
27cibhT7Qin6oNwo0jM9n7TxWYB81+4c7njtoBdpgC1pDU3Qh2DfDfX9p3W2TUp7
Qed9lbqKahBui1bxRqGuAA5ZMt9kh7k5ac9Ujvtsfv2pG3qO77mdl7oE5VsXYL0A
XssHC5/76RD/yuZWClhz5Ou+9JN2qLqOMs1LiUNM+sb+R4ttUcGRrJvqoonnSKr2
pSQpWrw/0SP16bSM/SEqs3MslWJxkeenFcZoH/xDMzAp2zbeCtktYitpvecRfW8l
Z/b82lD5FJV0rYqvHtm7+j4n7HORP9lUB7SBblTmndkHv42o05+ajrF11F0JGQbl
wLbcuMbKL0HOqKt7sfARhjiNxExE/I3YsAj9lPaKCK4aSm1SL+VbTsxBz48iABLh
9633w47vSDA8iUxT6nd66jVrQbgdOaZK/8GgxwxoGPlSZrCV697Iju8mEO14m5me
Wdrk59T+7OtJjNhTTb6vtoGinik0kOvtsQdNAnRgjdE3pBUaLc02xhbuehpuL61A
CKXw9jYGlIu/wicuwtTz1OwpnkLTR0jq2bH/IfTKP2jkUKDvjd7SibwwWRr5WbpK
g26UG2c66q4Fd+j9f3zGuaeiP04K5n80XRu7VcXWODsXd4h7OT1gsALqq0wFq7O6
PjJo7SZ/XWMoujsjpcTgK8eVK1SUmMU3RgdT8Gan+VBBtl3NZdENa/DvgRW0xaug
B5BRLxO/9vG1urs8TKc8S/SOy+tcNJWy8Nou3E0ssC9VepCLlZ1UCaCcOnUSaDv4
U02Q/E/JlZUVDknAVe91KsTzBlcyYtmPkPvRLdUi/qiTLX9IGtZcutRbhXuVQMfY
IgL8MRygGFuUdKbmVwYCovuYLIV+5zPDxGVgUs7uyfz3lmCCbgLFmEUZZa9Ry6ta
Weay9krANRQf5u06rQNq3ayZZ7mC2oB9VH5aLBJJHVvYkrfgb2JywRvwABjlqAdi
vmy14a8g5R0GYqStItguC7dHrO5lcSazKg3GnYKw4rEyw7sUa/GaHHufCmK1I3aV
djdqqBGpxbKIMR81wL62asVm6gUo1Q4jRGVR2p0eC03ebvlOPn99SSTXvVtXNhdN
QUwEMrTNFA8cOy1lqynlUXivpEkWO/2bwLajlWedN1JLXZ0TDVErSlDCkeDHqDWe
6VSBtFgJxhRi50ljBUHqDWbAX3vdO4pNCogZDXu04nVztQfipeKXUpx95P9OfUtF
9Gqdgw8vrv3F+Ze2OYMLrgpTnAyjGGOf4PIfD+rakszr3zqU4GmE+Fuf+uX/iKNP
7XYCoq9aXh0Xf4ElcLERAzI8QFsCsukXdaWZFaO8/Np1zadqUpTEkZof/I/ex9am
jzy3hAmC9nlZD38/CJKlLqUTi6lYLCE8mO8OG+tSK+h4oGdcKsjjF4E2DHlq9rhI
wzbmXO5KNZqT6UqtVc2kuGBP1XWGb6MiHXkAR2n31/C6oQnnJQ/eEA/CuN7D6PLG
aqhmcpeX81xi+lPwK7PtvCQUO2pXBj7/vDRco+qvGZGW+k1NWhOth8PhmPfpFLW0
Fqlt8C1AE+pf5/kOLUzge0IeeY4kRDYo05uVgQodtC8TkiBZJKfzunkfNcm62q/6
v/nTDtzcLODPSreXNLAsS7TBBlZYQMzO9bRPFs5ckyF7s/59/D8XdV5mkA434e3S
WBQVDFiMY2aMuHf8vhQjVT6tzczkXe7JD0zVTDzO/5NNcIrybZdSV0Q2xBOiuLUx
Cvk6RbyQEoiV45yxgqPx+kzruxo2FPfbnxtWubslFPLC93cla0Vce/lUpB2K77up
ctzXIcGDDUWPlV49NHRXSBrhL8nnwxLC4IK+H8EOHqDB4gkTgXzE1W+DwemO48i5
gnyLpIUD8WGBQdXVNhK+2DYcgwdZcbx8PElcija6a8UJVbhmSzepGesSzMuuXGff
FRizQAPxzWPyr8h03aR2E4m5HLRK4qCN1osW3wfnmbstHlf+zNMuB4eBuRTYIrm6
+L82jDmZOTAMIkEu4GYxnPZ6P4VWBG9Kc7T8WMOTFV5Q5+9B4RJiHmDkE7+9uLl6
CBs35tj7gbvSX6ZtXeYHslZaD2d3M/nV9x6/C4O166iksvvEPQcwNCiKHFvKm9Kn
99YYL4O/Y0ad3QSuMBPRaJ1f3nIq4Kj66FNUgJB2Ot9z0IEFhBeARy/rwYXtsVVJ
XHpiVU4wn6uRqReh2Z6cECYhp+F65H7eF01JkGFq7agcfbwJg7hqRBniHM0LJQTv
YLjZONRY9IY3eHzW2yZRtsChGWqYggKgGht83rnL7Wl7hN5CYAKBwvK0oItzTzdI
9yhZ6epQtEev8rPZ7WELCGk+yh3N7Aprzi2/97HYTBokfYqZQjyAij7nAWkioo4G
5VpKOWT3IS5PLSd0NmHqaVEo2fTMFSkeT3TFzRaISFt8WLC99PdgD7XQBGyXfvmJ
WmSGGZ1m6AUSEashzHq2Nlq9fH422Ncyq/RbOf2VgFC9Iz0ZEnz9sgqLlSZZjwTV
ef93Q0g/KuOTBLLyJFuFYKkBDZE9DDvQ9xWtnGbV+qup+aQGSvjfC8m3bGBVta1N
Hw0YfGYb/E/7ENEntkedE0tmkaFVqbPRcKcBMMGiQKvy4mylwKiqeXejX/CCpERQ
Ta/mVKsPPW5fDCjXHH7ZZLvNWWBm1sCnwhygllwJOuqgwT0B7bqvOpgtiBafVgWy
AIp6VyL+va1/EsEILA3eYdqZm/1u0CAxohLc6L2XdEHLxNUfnDh67lSAzI0Mq47g
3iHTasNJXHtIjxeah9soQD5+1SWWir3rus1hvqOsDlsauvFnMjCeVHUoJhBr/uO0
ZVZ+fyM+gajEE1ZU77LI4utqThl00TjVsGInHxRsWowCHtUURCMeyAMuBIMS2fa6
FWwN+ep23dXovmo2YHujHtbJJb4sWOetDJOQcfPltErmvjynwXS3N3i3RnimKl1G
LyiJta4Ptu6GoyhdvlgXsv7ATtmz6UcNpp4WX/NTk9WMFdYM8H4bMs067Tj0CClE
n3/ux5UOqyRn7Pg7qPySoTGNKxcAU7MXeORV1CR9WJd7WGYTm64pAyJqQR6vR3oR
yJpn+IIkT80Qi4Kg8k6qYAei8vBI3Xoy+RrT8AG0c3TndlBOFhNyH16g0Iizc8oo
201jJFHvQbTUyvVZQWe/xnOkOitenF7bz91htc78DXxngp3n2lkxVHKna5leRLtX
hXUmt6rDz0yy/Y6+bAbWfhMnJRg+5CEbwVEdXrd08mdYL18n0BHIgcmmfdAOo+97
frODqaTbkasLIc56DpTvqbsLlYlxTQvqb/49HS6PLZkrGVfGa9dTxKBOzlY0SmJ5
woHElx4tBMftRiZs/igOlSlqNbwayTmFKvBIuIRCsw1wXYjQLmQKMD+X2EWHcnXU
B6nvCRsZPInbt/F2ekkeSx4sjNQqdAGalxNdrl4n18rvZ3JrekirPGKIWr0ZZK+S
AjCdd1uZKbbq3ofQ3WCwDYEXj4UIcd9rpvjYQMIj9+0Uay6RInNaP11RAYJSqQ5q
e4sXiKY+Qp2n1/UhzWtwimHy/VjIH1RJ1yF37IJfuQ6INtCYcYvwyt2834WVmGlL
TydvKKey26wgerTrvrRbLUlSAQgNyLK0nTeamsw14jg1HBqrO+h7rwyIo/tUNYbk
PEyZ94FgvSjL/0xSmgwqG8HVrNuu3VxF64G7pwYsveKdkrfQUjDSe/fo5QCIziQG
HCaWmI83bNi5mQQucTPLOhAeK7f9w/3wcgxfBUFSOn8UXQKlEcB7W9oLJ0XROd4D
/GRTClyBF9NnGFXRys0/5xMOiM2Mw3jGcxuIxt8I24Xv9eHdohC9bTS7yh3QSo3v
2F1zvtOfzLq2rwSPavsVSqYextBE7QoVjdP7sXft0NOAGmXYN4TkG+vxmCTxfAXf
10Oor3Qk4Ew0dN9+mqCJw08ScLcKTsmM4Dw5dnHGJ8WggiiA+V1bPphC6OOsLQ1t
HiN2x2AlnbIHbPI0J7xNOiudg7Ja1W1ieA1fs1+HHzRkHGOV/TyPtKwsoz2Xp4eT
Yqy0LMNuLuIXoHMsXQ1TDHlNcG+DqMPizcnKZBZAKtQ6DjMIHxWrlsoh1lcC/6BC
mNwn7Q9w7Ik4Kk2v8iZjcuLM8d8E0/FomPWMnJiul9EwZbD8Yfo6HFdIa2ihwY1G
f9vMqz7Bs5ZmomhS/C7gsVle3o/1Vzq6H7WQHkd+9titkvgAlhO8KYIkOHDp0+Dr
J8mvpA1LMWQDQ6D32qlx2eTnwYPW4ueGCaEL5Hb19x0XRpGyrnMGM7IGyJCOYWPV
kGp/CrePTWu+7kGTMjLY1EN/whnSfVUSLXM+jv9mj+o86Qm/xakf41/Phk/FhXII
d75YiTss17A0nJsE/lV5R7eFu7W/9ARPaXlGoZQU9D0ZF+Z+HqUDIIAjdEp4U3w4
MlDNVYr2XuxCh6OUfcsX3s0rdhyoxpSZhQOWCa8XDt4YASXIQXlWyTYv3tQwtIA6
XtkzD9pCD3tMaApyhEDpypcJcAq+Y7QC6aGaPVq+hQ8PTlO878oDOKJrC3nqZ15j
jeaOYpgesK65lgUp+fkFhmRva7UEZgXnwU2F+OaLhBk2OnxaP4n/G4m8WYjl8U5W
98b/MaGg9UniCQHccvsep/KzKCneQBJqVJPcyJOqpAZkw2JhVInIsWpNGoEbYRS4
FZ00zd/BUeL3KGYPBxUUSJWuRieBu2UYjJaC7mBeun2LTPh0D7CrGncU0gRKgXiH
LPMyLFiOgTebU8OPIfKe3Xu2hQQZoDdJdA0M7yxlmCBRaTKaBt2wtVxOtUYY/kLh
vjeQNYQxuLv6kJpMlyLjXCTKyM7xMtjVlJeDjbqgiG0pL/lO7OLvsuyM4OUqBV00
6ln6Fhwlb33R85KUquktr4XeHsNAjBPS4Ar1ATgWNnZvRMaqTeIQUAhrb+nOJRkU
gCTj1feY2Vv4BAuhC8WlmCSaGGOzcLCBgDNOMiHD+K2wVO0vcmVAeM+J9VSlalf3
UFa1VItYX4jQfAndMBYyTbYIaUOYshyKKD6AizjufUDiw7d+ZhQrs7Uytzki41EU
JK6xtqmbLiA0NO3UtRuUvhFvvNZakVXqUr9aElURcP3PGRnTSjDYTwwXkzJOnaK5
Gk1ZxLRTDAu3DeN6F3CsK0L45mIDunj/rqgQJ2Sgs7uVJwh7CqEqejtsYUkDE5rP
6HsqTWxmzTIQ7IoR+6JRFkpx3ZlzoDsO264ZoD5/QfQjIbFvKyZnP9phk8ZfeqJZ
q7bEC48JWMrNCa5rBEdf3b0k+bCeBOINHY02n9lof5naAnE5908YY6VqJ3ZmleWV
C0KSnpruHZwXmC6I24SeoPBP9C2GLDaNkT98FGHHu/VPYmClnDcHbgD33HurX08H
OOGGZbP0CX/zJC1EjSxSODxN1rn02koO4KehB/SxnC8lkgwJM5opiN9zRHu0d6lz
GodjjkMv4pnboT7N6yYM7owviOY/CIgLdHuZY6wQYVOoxdxeHa/Ax3QE9uYTeBFR
T/UGAb92ryGvvYFqi+lmpulBnOiaIGpvz8f0VF6s6o1nf76U/5SBO3arbwb/Mpsl
I1vsteSeohGu7Fr3TMpW+zFEtaXX35BSUAVjIGAr++5oS6qo+Pvecn9bhTqhg7CH
TgdygZI5ErX/CVpQ4ZYTA0De21rQidMPMpED/ILAILt7SckNmoux3JKFqL5U9Gjp
dKPYYTngYg2qaJE6t6E4vRx1KBvcZqRmP1hvnk8ju6YxQR8KuPypxAiRGRAy9+vj
gvKOtMqw6W1//iBwFge80PvukXbXs0XjJ3rlowot6mFxcg7Bz7O409d4kb9VfACQ
c5dC92Y/xi8NuDoTfIScCMmTsVi8yNL1S6DDYXiYqD8tGvyjADMVMwabAK1wPtAP
x62E2O9ymXmTeEIIGuhRgqvHWOb4t7AI4Ymhk7oytaA7lJ+/SmuONT1hp/MBaTSr
Ujuxsw4Twh2AfOj57n5bFzIhaBeLtAQ0QfpuDsxyXNGXsYVrAu8MbJVrqC+/mAmK
zkkaIa4bnG7dlUm/728NdxX0BHMV4qkRk65repp2UwXB7+vyyiWnxPTrFnd7mxyM
eNV3GSsbA9lawnDKQ3URYJq9EbYz4sl/7KcXzDtUeGcCDnz1NeMcqmNLRgo0Gq5W
dMPFGE1aVh0ddr42Ph+qej1sjFf5om22N3uc8p4U3U4RqKOr8BIeMmB2uykVMYYV
7b3RrfANeP7sWbdRxmwJhlQruc8MOaS2LI8PuB0836GcSmdagaDbFF/k8Zyoc6lF
KZSmwZOJRcob5DGiidY+ybvKBhlNgvLqhva7rSD7Z02l6Mgst0P25iqKvHUqTkUD
OXZGP9aSSyUJJGNcgO6myzO8qjGUkpJGA53h9pfYJBCcS0qxkfsPDT9lW7ukIe+0
YAM1bWFGeCiUShhj8+iHfk3GZnbpUV9kUUcJDRVDjaaRevD3Pi903SFU/g37plfX
DE1PrE/pBCLHQwdH5ysFKKMtppZ1Qq3QG2VhyX/QDaZbCaAcJbYWJ6sGkbzU+umq
Jv1yCJTKufUIQk5CCE8b4l6/aiTVQ3DPlEEBGIC64D7QWsjRNzUOlJHvGdUF+Y+T
ynIM8jRgvkPAv5tInt+XfdnlbueV+OadsdYyrkK4koKAP3cWLq/7joWOIY2YhTU0
JGrSd7M5RP/cMHb5jMDFXBWMlLhiJ/wJxtUHy+ycepQ6cFRFxQzlyneyZKVViYaI
faoRZK071qgzMeRxa4xBvhP+J+xR2sik7W7OPwaXP5k9OOtWl4Bj1V2DcXvgT7o/
W9pzLOnY5K4Czcd6AGgVeUfe6TCBXnWUk2I+U7DWqHDCUtsdx62ldVVDQU/b2aCT
SQLWKM4RlT4xXoZrtdzdfLtLOUI8teCYU0b2UNNlJKKNXOgxpJOvX8c7CY9TZ3/b
PIPIOkM2aTDygWSmduiG0Hk5Sbt3m0AGG7VYUWE/qqjMd19SZSCpsHIvijld7Ma1
2Bo7O6YfdFJHN/hDtkHF58xG7viIgqDJTdOw6aMsqIgj+0KNBqW0aSTMs+RcgDit
5rHvY+y1J/6hCc1i0hLJYw4qHtia+OV8Z5AqFim8SPdwmHNxt/XC7vs5g6iovE2W
QfWHrLkqEc9jMKgxUx6gVjiLVhny2kOb4PpuVHtxxQDGjoQ9gDQ9pDbAOfAwkZz0
mlRMZC89dbj3LqqKDYBZS3Erjf+ZnjnGA5QIrLCDo9UTZLNv8GiwVj4fEnzzrDWW
oeds9KDq35uzSCiP7wKsqo5vjNxKodj9yAphWY0dG2V+2rrNxE8rDKJE1oANYlS/
ojmAP89b+EuEB4pguZYDNHSvwnLoL9q0Dec5C891xsue/xQtRYx6EICoK6+/a4At
W+7U/rKVZqliggYbKBhf4BsGqg6iDdAdMBOQ5vddIi+36QgN9Fme23nbq6rLdI3x
ARwEhJEXv36tFwtrdS9qWU6StUNiefUnK3hQgSNzXbGBxyLUNbSHFV8KnXeJF2Oz
6eFdxkH516AwYkK+4QX5h8tNRwneu8tPjOTIT+SnfQEca1FNl38rxTG0anBmV7qP
vDoYlHYBcBuzO5VFyFts1Owcc6pYFtbwAMA7S5BKn7UgWH8lGqopKwU2/Nt7o+h3
q67QmW9gthcpb1K7AzN7pDvUkTHW6yMgIgjr9dzwCj65GmKzpejugN1COjnDF5Zk
CeCIWUSyaWIufApW7JC8CABICt6ZVGHl4+TxUVHiDldVQ0Pr752fioxsEbPxmSGn
D+vtGrQY1BkDNQT2Q2C6j3TF5DwBNO0E34a2SxosAJO+HuQgjxwd5XI3LrKJMX38
kwse5SEcI0HSIHgCCQR2D7uorZrRqqC+HuYjQMdV9KuzsVDNecQM1+66uPIYRo+I
dGZKlo1tB6H0Xvj/kLSfk0jO96EsRLhRZHygidm4s/VCwmiyqutSDG8ZDwGQ4Uv8
kHULePJmCJ/sBZ6TKbNGDckARZnhHb66aZOmIOU3U14s1ZjFJMpxgO1A7FcZTq/Q
Y06Q2KBgonVcpoZyPs95pfZDwbP0f6mx0EQVMqdCmTI1UWrVq3fe77Lot3NodwFq
11B7ZniStdioc7UzVJQxCPu8krndpwINnEiwM47CaLeLGCGLYc0fmKD6oWDFKL39
y5d/d+C7cwpnlSlGyGJmhGqPlznT1VrDm1a7zQRoucUUfKhRV+vYEpuXo5dqJ8EM
NX+4uZ8QZUB4/a6+RDOGX6Krsyh3DE9c50KJCbHmx4SwHKe9SqurmzCqXJQigUHF
eQV39Uz8dWUG3Du+SKlvUS2qgHbpRoyvCbqAciNvGcfrJAM+6dl3Dp1DYjdSvRME
WXgfWQyjIEf+wIrCVJ4NOhD6UM68dUVChQnD6aMBFke95kKFhyoqV2YY7iTMFCnw
jNyTKZcMg5bv3TfSXumVirs2un1rbTZLk3+GHp/01LgIqjBv43MxD5mUgJIEvDdJ
31mHyULCcsHjm0FX3ZP4SdmUze5BVYW81jtT/x7QdQ9ufbxJ9+tYV/WeRmL9dzhI
25/08t8ovba1i1Dfvsxig41O2/P2T6s9iNLzlIfEYvOTQ/GOAh9QEV5xoKCoJGmx
n/LaH0q2qJ8MvFx0B605sypbX9xf1nf/tE0U5Ts6i43QOmx3jm6pCoUVVSmBIvB8
pGW4WN8AjDKY8YUhoJJh8rhHmLMP8WYWYY1zSH22LOXBnaAgq39jcgXGLvRK6Umb
nnDBbKVRENm3Zq57NEvw4x+F97HPu7bsNsY7sQ6cIwX+oG9c+4xSeKUiB9GQgbPH
FXmG3upwqu9fpe6/R8uYM3Zb3do7ke0L/hSXuVYbnqiil0g6r6CSKlyFTjXg1873
mb7uufiBuHbw/vDIFLQjCzbtojMollHMTCU1FlnERQo0fFeAVPZmtLDe7svtOHx4
wuXeb2P6qLHU/y9kZ6GseefJq9uhEiOpfv+BDj5DjrC8p10yD1gBCfT3iM32oLDh
Pgk9oUX/ozb7e+51Sj1EpUF4WWjlpc46HUznX95oPf8+vRBoeaWeRlXmD5k8uS9q
sVdf1/cuNXcJeAi6EI6en4JJvSV/OBW/Yc7OjWFQ3+5ay887ZtUa/VdqDnJumZYh
1Xkalis5rruE8yRUWOigwErC8Q67fvR+Q/XwagIlOUaKXc4RgVH8R5VuAjVf+RhP
2yONaXHKXpymdT5cILVsOGaac+U+8VuiLrTl9QqYwidkEUXF8T580fDaOxreBeEB
XUQEgPQGuljFp4sFSJF/cviSr7UanEuZAxY00Ary0nSd0EOicUOXUp1D1H2RyIxX
1LhH/i+MCuGifimvEWvIY5qYjg/jYywGh5Au+G+b0EaP5CuZ9AHfhj4lGf6eWwBe
U8xCbeDcDeV6jVFVM9LW65srDUUo2TnjLSw+gr5AfMCq9n3b6oTPAgRuQdTrxDgc
xC2AItXZMCgkA5PR8h6gwnvmM3fbUhw8/dhoakph32Ab5ieg4L3fbcCi2uQfP9tr
8JXV16JCZg8MIYsnRPpEh/ZNLQxfYqmlD6Ltn/OWKMU4VWE3p+30XwPd4tS/6YyZ
d04wuQ+COjw6P4XplXJw0rWR3eHFwWGuNL/TefIp8+vmssmSw3wo60Tx0roxL4nb
LvhmXfY7hj/HG64mkZ6CdXEr66+9IKVJjtuDOv9IjFlcfyHbNwjGt23pCalFP1NU
yhjpJ0ezdQr3riCO2tPgeYc0TWOF8eX/L+R2R/kXl9M1u0IeONMf3C+Plavm3V28
2/RkxJlFdPds9UsShygTr0qgdn+hu/Dul6bKtbNvIypKnAemuRtvlElua3orvB/T
xk3bMkvjpG54mwkl0mYbXtjDsGP0eDylXcS1xn1muvZEVyWzoYPK5E4uhWmaEcc+
QUFtBuQHrjudzhQG1wNfWEWHHiNBajSnzKEKpQ9Vz5gLQQQ3L0GBTtMzh19Q/e+Y
M1aqmYD4KOWbzVasxHzor3nXDRp3NAft7u4LPnKs+mLujOvtXR1BjP6/8Mftxou8
0tmEa1jtdhTDPRBKSAhhKAs4UWFJp/u/j4Z2y3kcYY47xcAMaq0PEBiWs9/jXOhU
h7VUe5f+861CPvmB9aDH4okFLVNinGobmoffcFaSiYVr5WMTVoWUuVrXf+x2rrgv
m3I73srCJzNaDhibDRPqQakgFfu1H/a8LX8G22xmTrC1FPJ6cWPvpNnsEbrzqdx1
JdPN6rSjsn6bWhnqGbb2CgdwR3tMiRttHp3L4t6rO+jxY286K2kT0KCy36kaGNFo
ef0OsQiycCGJnXG/SnacuwHbA43ouR+ASXwgYbTxHnoHRmJCwO0GuJmH3uhOP4EB
KOvKbbHFAN2Hysa2ZNE6v36wOpkZecy2OXL1b0IZJ6RHoQkuTDRb4WvNUP9+d4+w
k9vQ050tYWDOMp2lI7OGes2lN2oQ49mgjBy+XnBAQMX/Z3+XLZrD5xT9rkKHwm1L
zcUwJVXI22motr8Tdg+y4pQIrlU7fGAhY3j0F2U7P02iI9aqXtfsuMb2Us4lR4gf
9InajJQAvmaG0o2+/NUUT903OkavSYhvFyO/rQA3wZN7FtFI6AeNg1K8w/r3QWcf
WlMezm3N/RWPcgzwpuxY73MMdCBPO9lZVOcyn2CgPDrcsYvcvBVWQiqQtFUteHzn
Su8kltrsNF7/OVUj8nDw7yFaNiPNLLGGYL8Ns+pLkKrA7yiOpNkGm8fUveFa4iJI
XsSh8CvXYUpZfzPwYeyVOgMru7sdST4AzTicdLAzuOnS8VpK/ehH2bDu1r3tNLOr
luG9sNeNWEl0rvYl0d7vzA46NiAx16RuB5lgYLBypL8o4kvFb5K+6hyOo0OB4LdA
cz7JeI6OyfHI/lZx/59EdYiM2k//tnV0/5tSq3Itf9cA9yLYFN9wK57JteDBi5cT
9gHHsT5S8td+IDplDC9qbpWDx+T4LruqYwc5nv/gH/8jHZosibNdUKlYFMP2jjBI
Nj4VfKaMlfc/2yxvkM9W4fCBDSNWqDUYKs7nLKVe+TKH66m1RR1UTaZX0OfatzGy
fyCNTDPMcDjZvpVHiP6N/+sEz9qU2dBaKWJoihe7fDAIxpcCiaTkJ6Za7FotMkxs
C78tBsVkmP1xUM2aoIMi+mgUmEsmf76GyayV65IgS5J7Io1XUbrLELl1XjI+6dIn
WkfWDL8mPJBeoXlvByO3t4FWxVbmrWJ31ytHfGE5lf1LWnob6iO9RAARNSnA+xJN
DOJ6nigBDMCmCIG+HqiqFunAr51H4kdJ+nQbL1I++TLC5DQX4cEAo7pxQkVXXFAT
3W8rkiDLGxoru49WbMNTr29LMQ4GHiNruzXGsXoEogG6rnFITusn8LJEf5WLpwww
CxAUiWlXkW1ydTUdz4CkN3rmnhfMNw8nMKPHOI9YmFWcL1kq0VSUx7chFdyYwN9u
b+mL71m/ZYF++V/p69k6tH8J6HByMsY2YI5PwPluKm2D+mUWOv87PR/WHl+6gBOn
nqOCAZ4Duw15NnkH/6oznIs1ef0uzyHolYYt8xm/DjukChTLkZXjRFcq1Wv65+jU
wNxfYvixH+cjrEylvjn1ZUMY6UIWZ2Mpd3TO9Z6q4mL4M0IY14AsiVYSK6F4YpGD
h6QhE4Wf0iO+nyrI9K4MwXtup8hEj/P6CbKgV+GMxGmwjkiXa0jZ++2NVh+USilK
1SjEKYyX1ld5UBrciOGFuiT89gi0UKd9ahvpfqdGsz6c8a/v+Emd4go+aUW87VLA
+FDhuny9PtR8y/SCqrPbj2fKpjqpoUddFgSBNPbHfdofzJ8avw2q3rQKQIwIUtUc
6ZwQkORtU7GjIqFXI7qKNYrxwHLjMhXXDY0VXI9AJ+ycP5DXabQnzQykDe8qpjET
M+hAIjf5D69RTBmkdPCeJZmbG8f/cfJTAbEe4Nm66iTA4qxXcnOHEA0439tCYVZa
NcWpRj5jUGikWIqQsLF6syOYgwOtScxWsr7vu/kaus+M/eMB3GvsvZYSHaX8U4eG
prg26MOB71sCL009Ilu8/GhBHOfYNlIxdmr+G7tBxfzylfbgNaRC2zFxjed/r5/z
cTqHnRtfBZCePnBYgVWYDMuqEQieSfn89bblLBS2hWuW//1oV6XkvTSwc4FN2VHj
2yrw2Erg6jfWMOgloE5iRHZfgjOrmklBml28jHwh6Zm6hh8F7qm4sloEu7XCQRI3
XCfMCATakBvtohiFs9LF+Zt3XFYm2WEqwnIIrj+EwJhtl8CHEOYuyrpbbfRKRk7j
1+NOCU8lW939PiuFotGI50lziKdafnLClg3cgnzfi7ttC8Le4sDqo5KvPVuiXgWE
W6HEBYNXgmjQXGDNnbvE2DEApHoOl4Wo1sk9wemzvjqiYEQNzJqxisgfThcl8urk
DLZyenjAR5Wi3Fb7gGSEFvp9oHXGzkLGj0sRAqdX/92rxqtaSXZVSE8ZUiCZWdYv
tEGuVgykeA5T20QYjjE2WV8t2IJ4SMOBofac6D9EdAcbpG5dGbAO7ie1jTCjmSXn
ARJ1vR1TROqe2cGW2kUuxeUHkst1nuPiFa9jG6DxiQABBktcsoagtS+E7jW4+ymq
sxQZCXrEns0FCUpu2ROkYyBuQDrLQqIw5kAlM7YvN06Q35coi2UgIOiRR0A+fLEP
XYn7OFUlacmMkUzRdQjmZNVFhSenm3c3ds1CwCq8Ury2PdOH9fDpdVvYqXv1V+o3
nChbYyiiamradozvCzpfl1a9Ey2yz+fK7PRJcuRQg89Y8m0Ff5KsNAI8ND7PXkZf
GaCfXKmPVcd8wrjpJOmvmfHIFylNwrl3etd0f4eSIIDPcg3q0GPYLALsaKzbUn7f
ef2gdT6br2GlStWaABOavcIcWssDnbeS5u1nytlvpsc/Lai/5omOdOBrEjeALul5
C31UjyumZtnaiS3f0SgoxI+OQYJEziJ+Ap6ryNMFFSARi4I/cmSSexjnQUXF4M6u
pVd7XXhafqPdlquejH5jI9ZBMbJXv0kL+wvBjysff3UCGBm1fP+i6dk/rFTKidsA
jhHaRoLdia58mFojKuLDTBax9SOT5MB3fmBhTsaDvuB6peZZ/xA7RXBT6sSjykpU
DS6wvZqFKldyrV5K6y6gQ0+ivzxpscOp5Xou4QjbZW90U+vVbxSP7gTJr1OtiwJA
S6EuhDYIiqG9yxJaVrbm736OFSb9IHdpvtPo3vOra/F+/810alF3ql+dOuItCGXz
A0opueqHTXgBewI8Ai32S8UDQHH8l4GI9hmfvyA1zEcWEQxWlUavdpdp5jbaYCgn
EBfuIhfGy2q75dVXtpG7Dsjp6tdDYdG3ZQJ7OiMqvWfS0Kzw5sN1EV+SKW51M8ci
J249TR67SqEVX2SfiEk8DPuHyu0E3xVpqp0L8vSDUo1Bb/MH2cgUNFK3Duy9LWQq
J7Ow/gPnmPj+vRBydjzInTxXdMe+cu0HUoHGIJelKxl3KdLHdZ42e2GCvfAv1ioN
NVb2O0UEPG45wy6mOQg1chgw0UMPdLxBkCDc+MXNQMfZtxbpT1EbmwNR7HUtObAi
FPqy7DFArAqYmEA1Wvopa4QbkJLizUqpKUYEMpdZ9Ge5t+gYYBaOdsC3/2f4h9Yq
nf+NqLh2CnKQOe9HraqDT4De8b9+ra8cx6148zdWpw9YG8nBfCrWjheHAFWN/nyd
lq9O+C4dS4k5RBixvPnl1jbjdQr0gZdtEZXqhiQPszBEWA9xNUEHl/7OcDRNJ3vV
0FvU/ag8CZH3i3alYiug8Gflh1ku8gM624jNbmwfH3irpsGQG98j8hM7FHC+3QJr
S5VdJl49sGS7vlYa5cMZ24VrPFAST27alv0CmkTZTdUpWXzo2k/hyyLsdBzWT7+c
dhfL6P+XlTQWzk/O7uQvkj4VKOy4Rdl8ofU8DQ+Ha4Wfn7Am+1gv2VEkB4GjuzpS
MVoJ5MbGdUsEt4gyD9RKcheMR6/TGfhA29Sn2ADioKGbXgUha8KxVZAyZHs14zHy
OghHBJN7d6GHHPiDlaIqJhTcxZL8bV4fib3HuLYvp0DqsMXbOEaYzraF44HlEK7r
3SLRmjzZo88sTWC0jpuHCiFVSgt7gAMkiTz0hczkjojPMetdLgo1T1j+o9KR69hz
7D7opeoHBcucknUs4pFwxp6TGqtfSz1eXPCMjIz6B1hGxTWkG2dvAvZbD5cBT5jZ
UWOAsAD5MyqDOFlAt94HqSNDdLArmxJGG/WD0NQ7Uarbzb2pp4A4TWHu04ujyDW4
k7Q1PlmT593rhIIxX0Jx9v6hDxC8YgPGNQSJVM+ZkqMDFG8AebCIg3/vzlMcOb0m
/o15rVD8fBZZSR+dOXcAJgFu4N4vSIfYbzSwrYJrS9gLTJu6Z0GxtyHsvpnl9TLA
Ugb+3dtk1cTg/qvQaMVhFxRA4EPgngLnLJ5BUgL4oHVQhRehI/tvEEiFl0q07p7K
OTGmOxff/rYlMhrfC2oCayK7qYgCF6/ymYjOJYG9p7hIhI+hHMXsMJRmxR9XvfTz
bh93Hx1JA01TYCr87IHcaVRfMSBXsJLfu3JTCUwrJdgiHwActsLvkqmVezMln4yA
qHHADZf68arv8GfzKUPaac295IZDjryIxoM0v/KOuAHjrdeUqvEgV7kVG7tuBxcA
Vmv6xaE4cno4EZnOFoR8HXqzzSBZPs9zlcIc6XazZoy2UKAtKa54Y2ZkzF3XuODM
0H5sgf/0KujctQdSIf9kzeMMZrZiEz75wyQVBJJorC6r/s7HEFLB69so1bOaaro2
f/YFYLZyefUBGSvX403uQGEENijhYc0QHM2pDHkYRwaItuNZw6V4AjSDEFSfvO6K
ycq19YdLH3wPodLI5XajtEKjozjugbwURzDfeXOkf9DMlHZCKHduchiwwM5l9jvM
PCy8+3m1JhrMQRfRWC7/ej5v5sxYZrjwCIUraWPxto/2SspEWQxdPNuyJN3bbbDL
xrpCZi9+nwBj+VVMoHz1yBF43y/LqSki0kL9mOGxDIoKVfHJabOEb3HZCLzgy6bl
nyxeJHfU1cjw2VG49EumY6/SjWD+7v+3tyyfOncELIiwWXz+RFhiCS7d6EBBIdx3
2DpGfft+dBqSYN5e/Kmr6i+Aaysb98dVYI04e9BgwuQiHbcPMAauV9qP94TWCmY9
aNYboVF3FrgOBDxv+HHaiRmLJndj1FqfCqEK3+turNUabutTLCmK+dYoJ9FZCd0b
SFxKcLt+oVhagxysYIVitOAYvnirpsziJ6/jGpXs+Wc=
>>>>>>> main
`protect end_protected