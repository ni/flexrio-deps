`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 45040 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
4NAZGBPmQSC1EoH0Jm8NyFq7LL+I6XKWaSZYzH2Uo/uRl+mJwOGFU2bwyR/UQ7dZ
SPJ5XMUayyWPO3HKo1oVMtbquxI7WowsLxWi6wKnoVbPQOyYfg7SZ0IUiswTBg9s
KDBtRPwzE/UtBhTT7IyC7TZruXG81/AiFxvauxJCNE71WY7CC2SL/UekUcLLO6MX
rNZkX2gpNGmqxcsexeLur3asWZJDvuv+/1Vhiu73v87PpT7YU0RKsK1WkRdO5P38
HEdEOgf89lWtVOv4zzz8jdZ7A7dlhipS1HNQjKGICSc5ZfoLVZeK6sTchJJE1sBr
g6lZT4BtSogXSHQmJOUaj/V2BFOx25bi6mbG3McCk1oY0kMP7sBYd+/mCOpK24Fb
Jg9hEy/M4J2xfxCFpr5XWSRbM5cewuGE0Mxc/U30BpvwHAgv44Ot71ZbuJ6eJ1jh
QakRpGYCEnyEyFRI8GV7NjyDyUVRLlk1BjUJ+/MVD3ebl8ercj9JrNrDedP0H8MT
HFQWUKtBSgx9O5f19evTVgGYu9wkrkHoxvyrlXKxlut/D50Ame5oTPoD0GDvU11a
7hGxOuZ8hazQyGmM6jI4Ku/s8+ValGfF5aMdkuYJs21J4yimAMoRIFjiv75l8ode
kMTlVscUaye1vOKx7nwmwJ4WcAr/7XCquqXgfJ31YHP0u3hm5ae7QMtFLNs5H0bZ
rCmGDUOgzPPgIRH79GxZ0eeBoGvcpDRIB7tTrNRN8bJBMKbS8kNrEUVw6LSJXZnN
1PALQSzkKPxNZqHGyfHLeOxPHzYir4wE6WKG8hZkgkUopnRBmiblknk31vFL9mjj
qecdF0/hc9kWtGKAbjH71uefxOY/oL1qwMegeSGdjY9F9TTASZ0+C1Ct4WicNLJX
ZE5x/kDZhVFKG2KnD0XG2g3zVT77inZdhExK+A7WbPyDt0DhKrLZ5EcWv8sbDi4v
e0PIp1w8h4TwYtTAARtwJrW0nI960yuPvvd077rj56jeOerEUmQHwd448966kRqG
5fKKNg0qiNS7Lr8afb6dZ7THPTsq4utiaLA7tcA0uvHXpuw29m1rP4YAZHVs1Kz6
s0JasWvz3x4j7Lk6Xdni/sYr7eo/A//tGNTDOdXnHbI8ACQ/icgyVU7MZwNQ8bvS
9zZLLbDbaOHIA0h8u1Rfq3FYDrUSbGI4xXLBkeiQg2BYOXq60v3L6BViFWs1lpr+
QpZV4TnCjzvO2hd0VaX1Y1rlT7malEBwTA43RKUPq5wIDB9iIwCAtduvgx8rmnhL
iNmJFi5Gxgv/+PnTlQNfFznqvefx4XGJckyC/NxzXZlQa5DiZnc8dbz/NKa1Ud0n
66bVG7mgJQIcxCaZH8lb5DxIZtpWGNjXy0SEWktrKBiOXS7uVGGndMsHp3+HtgDT
RNo+aOZgELWse7EVf6mgF+2cKxdl3Ovq/Kgh373CkVPBtJyLl/s5xSxUzmVoCiEJ
vAUTbBg19bS6YuwTmQ8Wu7hqQOtrzK3i17bNJd+WfAgM71NEL1ZENJr+DvehFtlQ
inLMe4fwpEzjpVMXSm53tM0fdoYjhlOtkC7Hku8jUkbDPUvBT0bWLakXdfzgT/OO
fr18V/i0Wve4gOGSmYPxC9aeJ5+noDeYgIAMhwmdxSmdSs3mp08BNfkgqiiYNDqy
DP4k0jXiDI0iS+HcKXJYIuDbIldhE+vnpEyqVFigSU0ICloJsZyyAoEzgIi/bHw5
J4fD4aww68vJBBThZF5hkzg7kLoGHA9F0PMRJCGziqCYwfHIJxasAjM5N3kY50v/
KE6WTlfa0M2rYniRfkLR0Swk4yZU9FWWXhUM61l64XT5y/g3lxdNFvU7eb7lgGtv
M/33poP1uJQCJOl4JUP9dyhF36zhSa0twIF9qtIE+kQHf98kW/LHH2xVPCUgottV
dXImr1ZufSCrLEqtGYjqRJnOJJpzrRuJ8wlGNGuDdQtWB/bB7Eu2t+ST0+VJMOBs
n2p2xpnDCG4oujc8QbNaxbcIFeFGiiocgwOQNSGcIh3DuJSkRf7Ny6nBlQbCQnzL
paTD2PeiIOQllZ4NaFKKKpk0xt1FsP2m8zvbfcMG52xJQz81XgH7Dx0z0lOjHt9p
3r5Lio/f2Q2YRXQZWOxMvrdBfBSr8w1G6jRBacSTVq9lnP/WPf9uYDe5sRLUNESg
9yUiwtvGZ3NTcZjqfLy7mFgWQu/EgFJW+Yc4vtfG99j2iy0p+WJli5TNusWLn/4h
Ehcu66avH4ur8BqvNgYCuLhJxmKCtNEi2H5W873ArZmvOWebqIe9nK0exf+5s3RM
kYxBoDPyiwx5JCnNgxDU0A1ZPmPt6VyFcd+Ioh/cZO1HIBW5/JkCOFBGGTTG3w88
37frUGw4lfj3jKFKvbEOcDUIZVOZtIrTR1bMhWYuu4Xwpd17VghSLmvP/kHOq5Ac
yGUfBxTV0TUBf5/2xsneOVeP2ZVF5EXzNXxBlibWVmTdEHO6P4tknoY9KOF3LDfs
Z+dgTWlgK6HwiGiqVmCnLaTxsJpBg81MX/v3VdPB7QNGgVzwFnq5EjMMpBrrpVm1
oVhKDKlVxIQyKn9f9b+OEfTP2tVUJLPx8JB+EdQ4bMRyO2kVkjEoSw6rR/DULhti
Kt56Gt8QaNH1DAVe0p8uadWXiAMnIzekSWm/UsynfwZ6kXf/fTauwWKIK3GBpcbk
1xcyilKHCLhPv0Xy8bkAdwNEeFsRt6ihQy2M2ujVz5B0kAYnCmCaXhRpCfD/Gm/c
bbfH2R3oBnRYeXy3nGhSeJeoAeLGUgB+ekRXn6z44TsFcSHVFgqOO+wEseb02ZUe
ZJMI/WIwM5u986FdbVh5d1m/ei1qkSM6VZlrvY37A1zegBx5qhf4wZQaWqqLHfJw
gTAFvShQPWw6iqYSZL0fZJbx7BPdk4aIhPu+W7uZPp8Ne45jl5jdj3xXPuA5Pnq5
MyfUZfmzfWXj4MCPAA789lVDhO/G/zzunWPbHw5RnWNLdeT8Dh6bZXUtHbmkg0i9
ZGDjNUcEXye4pMOdSBorxIDsa/LNRV1YRAcY67wqkDjCf0ShRB9nFYoR+5iBT8os
4eDcfrSciNF0B7ByfTSUnmuOhoaHUvZJRY+47RAaxTgWfCulkaqiH7AkKkDb8uZD
gDsMJsAhrnlzostf8qSUkmDwQSeHYGIFXL2VzdH9B3QopGwsPZIPAGyrw+ceyC73
62jP123tMEb2qm3J6xUtoZR7vnO6GMXp2mFiCX9jR47vgwfz9LK0OIPls5eAnEvm
kCgWQilx6POWKawuow8QbNgLgWzPwkYHnkAchapvxou4SxjM212nyh4imHxEtA1J
YmLxXeX40jQV1AatW2AOu2Q+AhQT9Scwg7pkv0hxaoHqgNQ4+pGZ7mIEOO3NKUzc
2cwy1ztI5BR5CXwghPaVus5IZEWwfxjs/6c4mGHdPPtBTn1MHbgUMLsppqJvJjZD
rFaLaVB1OUwyHVACm0Ik8+GaRzr8HI6OkceOmvLt9CB8UAbf0KAwAOgqmXrrqkcP
Gjv7risbfsWFJGJFKH1yDcq3bPyaKz+PuI6PabPm23ezivA+prxPYU7E6aQ91u0g
VMv5GPjFrkuK4saGFODc1zpgAkvLtTuiMdc5YNUaHbufkWZTqAbRDKQq7pSamudz
+5nY0RRBpYBKklDD6mHFIHEFoBdntIxhydK4gTxRJAWB9E2pn0Ac0DQTFeZ30HQv
8DhKZjd7itujfs8ETtUlUPLPH3+jIy0xPktspiuAb5lJNkAtNam7TE2foXn9nS27
729BYoMfgRvuNuoa+zhegicFjxzqhhyzgktr6KwBKQlRnUQCks2Wtk3QP48piUFL
GT6jit5InCxxECTMtwpNEt1eW2DS0oVlIfrBD8Gn1BeTISV/8tlhjxfqsDgtyVRE
/Rx6ePYkv+885I15AbLTba6Sxj9z1ndMbApRUBnzse6JZuOUak1MFIEknAo6ZBPu
3zB+nGcjq3oRN9iLYj1hBTCnyEB4OlASzJFyCdtUXN0Dii5oI74hW6JVegW+DOx/
TVb6QW2IloyKQJT4RTdUCr2SFotxSdi94j4YXVi10VUvLdbp02QISsqS99qQjp1E
B6XKZje4S2Hk2bEHJDBGvuaRjzwucURmiDfNPlC0OWJ5++5U93HrI43rgkWg2Lmy
S4NHsAmnAM1Y+N7ail/8lZm46HGfv+02p8zMGX/YcoBoBixiSTUEeQocjWcPn7dn
Ccx1m+G2bfKWhvu6VbbKH4rVILLTG9l3kZ/sRvan/ZN8dpj+8oJqYHAgEOUSg8xJ
K03tW0z68xPDHZsMe/CLplN6+ahbtXDAtv0opZjfegqfqHkO41rtzLTHb2tEEXpj
iISw4vuKhIvHFT8AQ7qkoxDZxnKJidtOTXr8YIhseTI2VOq96YRF3UzZERAPsHlE
9/H7oSlW5dkoIYm/gAJ0+gHlCVl0vwQ3C4205/fuqi02T5OOzjQlwI2PxEOQPmMQ
ZbN4iKKx6uDw97dwUpWUVxBoJ2Oiv1jNqQzM34VgjdAYPv/ApFd6cxsIP8GNrPKN
K2UTJ+duKBI7sZymo1opMYYqiXBGLuOqkZuOLS648mG9xr9W7COdjJ49VvrQEFX7
g7JgqsfSJLUlgbPuKhP7ceVDsfuA5E5IRQpghIcb2VuMa3+o8Atu7vPEpWd5+hDg
LWDHf0wYnazjB52Ryst92WYmRIoVc7b6cbObXMwGsB+1Z8DizHAYd3NuvOiaY7kz
1doKm2I9Qb3Z5ntMw4hkoNKOqavd0zSgeiN3mq4Uxi9wPT9MZFT51kpkNQrHY0t7
GtjS54t2Ct/dPdhrPmqSvvruYPpruiNY5BlZhHYsiHkCG3+l0dJaetpWoWzzAnhk
emAZcmvmD+oXYBob0aPJg8wtMDA+BgYw8ceMDwog00rKMqsLFbHb90/V1ou1M378
+NJi6gYzrs6tP5uRgnNwlffpbBjOHc+bEKSKo8M783QZ+GHrXVwZxsftsQ7OxR+4
2rPZ2+w3mQzGCqmsNJLTe5ctc5lITUSHCCSxLqo3f/sQl4QCHnt3TGWHX+RJoS5s
ka/PgY8b505TY7dTYKUN9BKb41LCDZLPhaBArWa61lRrOpnVIfDioJ8k6vteno9x
5R42i39rWaAADtaVg/qyLaOUK2cZqb32cZRalIUnQrsOwU2xqvBIFOX0/Nh4UH/K
dlxwbqDIRbNjztOVu/KwgJOYwEpHaJ99Q8AFhpgpnGuoCNRNy+gxg4kHm4VJ5ZN+
8vQHiqQCcF65dxIbJsfPlBtHPtOmF+IRsiuaN4dAH0uUtRBX3iqUVvXdx3rpSszf
vOa5jJwTz9dfo3x1oy1KB1IqIU/cpMSqMNeavA7NVF2rjDsq9uHjUzShd79i5HGa
DbkWw+B9s4fSzCXnnRu6t2I2UULqFt6PxH3GVAYItbQkVT/Th06LCr6JYtJiuHzX
f+uCL66B64/EbLA0I72vuOFYlp97lra3pVgfWi2HxrNWT9XEARXYsCWm8XS6aUDc
KpI1JMIRYudq/LJuZU5QSvSv79nkZRlXFbEOih7OU1CeFLMnDdBP/7cl5SrttPR9
UtHJkA8gQcS6YLe3THJ/jn3QivnaApizyXLhUR1GaZCNurX16m8BIVe6Ity6P/nJ
H8mCTZ74ZjniQAuQdlAz3lDLpVajbRpMglX4e24m6LBBJZwdm3ulZbizhnfEklwF
ezPN6mM00xVjAcgX41xZvJggh38+q6qIVy2LG0JH3C6cJA4rdY3pfgxDQpvvkXX9
/yvWRfP2qzhGO/9yKSAoKJ2HUG5nj7X8SRQMKBFtNNFVhqxMUcPvHqcwAuizn8kM
iDV3XsuaX27pA++m7u6mY4WEsJAkEb28YS1ZIgeE8+UI/VpwuqBmhJjtgDIWD669
Hp1KEarc+PNygEp0hSvKetVaY7X626dMfgkHrikTLyHDChzI4WATqQKJdi7+trDY
O/P+Kr6Jso6yh/sNZhBYRLAGt7fhwIoOqtEfIzD/KIm1qc5ahGIGFM1deRIWxk3w
pNFjR5uhpW5DeTKyPLKTWSierTlfjbgBbqrhJaRYpeAOnNmuf3dZNDn/OvNpqqSe
aMxH7Zpn0EtiYfM/utxuVDJZlO8wd8a5LUGj0MMnzQLxT2e8/BscVSvlxdmd7WYd
LZHHGKrsiTyrrrlB/EK8hMIUM1rMwaE/NKFq2+AU/fDxCZY1JP0kcovoi9DJpjGf
yrhuzC/5COxAY5PAjA60hp/EqwQQxrV3+zegv+a3jlJRk3CIZUhbyabQfmelqmpz
KlASd9pzA4QFF/hT0WvpMbBgfxglWJMEs+2ZViRvfVMVVEjqBlIp/IX8iHBYc6C+
J/Dr2UzMq1GrkHlHhV/GVvGBYnZ4/EaH0ufIl09oeEuKviK8QWiF0kuaPBOcr4nK
EzQ4KIeO2oQ0D2uQ5vTQQ83EaTr8iZG7C/6PNKK5efc2UXDaZ5W5nrDaAlAePrwC
KDNc2W0iaCAdfbLON9Q2X7mPiggsj/Mv9P/ATuX+BszeQ4APVCgqm5Imc7IAuYPg
AnUD88qw/9Vrx698EPxz9WcHk1Tco53HfBJ7zHTPW0IpR5IX43jU1HDHRDTkTJRD
MLyD9r6ienvwKEV4ERiK+oLRPJ78fX1gvCg7f76FGYFuvBA7DRnuuwZ77B9agJy8
Ml6ucEd7LunQZe+SwJ1pIIJIGW8+y5GKQ0gOeSgfXqjlHI5QIdPy+wC/ph7PDTsV
hguxsC5m1ZQmjigTA+eb0Pu4jLxVYgqwI1sSzCcNFvpqRmUsrGw/Ya5Z9AQ1iUl+
J0b/RrOidPqenOW0paG7e4RA8dp4xGmIYcDmbApSt+u79k4OO3jaIuvhi6YnWc75
PJ4EHO2AmRUFl2ccvOtvxkjkij7smpLjJESPzNNfcMEPxT6H+8CORXDuW7+dwE3L
iyzQlpOMYaEYV0jXbsds6x6PnVKdhQe6/+nFdMiqFniJvoapLR9AlcHW5Tn0I0OU
5+sd+cFPtT+x9nqDw0kEbdDA/azOvDlK9YZCsbdWM3KV+mQP3TekTXOx48VVmT4S
TyiUBDkRBBLZpKPcjsANdaDirYIJhCh0RxZ8SNGZHzOShGoGn3H/I8TA2E8ZjV5f
c+ydo02SqoXek3kAsmfzcVBOvYWc0ILuHvzOtvaehOU2eq6wF4ecaj4B/UJdOHRZ
g3Nkj5mLC1bxwyAB84KT5pDdMI0MS1QhyU1EK8Ztol5n5DWyjq4/w39gxMd0fVIy
BVMEr50wmhCGA3511tJERXKedM6N6GLv/UXzdYleQev/mJiUj74BTd8mLg1olC1A
kDF1VLfRncCYnz+2futK19x1yxqelMofATLBiM7NSMUcL/NmSnRGX2YeZ5ihTQiC
F6BWb02VlDfT04v1SJIBHY7NyBX8LmC0uaTSrHWt9sTNEYtxkcROKeQcYk9AZxxh
r2PrOkc2CbTML7nFTUbRHk/Lx9t56cMFRHogpnUMjVudEFtEtaC2lgh1uRha/o3s
G3L9jLMa9+qMpGpwYBd+vVJv0hSJwTwfX0OfBlxpQknstRn2qFR5kbQSAKO8tDxd
II5w3hSkFTUE1ioAZzUptJxY9uGOr3EANUMZ5Of2Og/2pPENyIpy1SfJEVQJX3sm
4FJkPsSRoVgBUzwi9ND8PNNuUZhYsNjLnPCOITB9brfXbSATXOK4UExfXm6uX4pY
9rmBjUqtPM/fmPKLDz7WKU54EBSe4ce+UQmXJQqu+lxAbpYkucfr5SMOyjcOYkmN
aThrsGULKr7s34tqvWdnfDD/89zWseb+Jd4dZ4JOWJM0rMwJ/CGRyBfGHS0dSo6X
E+n4IN+HsnMVFNuClYfkFZTObMDKXo95tN1rwyowvnnnbuAVgX0vp/athyoltS/5
RGY3LPEk79UiYMZnyBjwmQiWgXPMxSytxSbnR6kGzj/p1Ywq53N4t1QxVRXrAHtQ
Rwp/VGTNKMJomvzNIo4E1C1t0Yagex97/yNO+r+FX4DlcZT0+5PmHumHjYjDK/Z9
+/lnf3h8sn0mvFSDxw/51H6bJKo/BXNLk8UTjYu2GDb0/w+vlYMm10JXC4ybwlWJ
yCDILzpMARUcLI6mnMk+MCnlI9DdaAksvw+dT+5pBIfS+QYSnqOr7GU1Kt/ALrBC
jHb282nrUdAa3Ep3AbFEEkZWTS2E1V++PieSTc1hjZoU9dNa+af5NgrS3TONOXNO
5hNNUpP+dbuNFGO+Ka4sDyyg9KKPp8obeQerpqRHQPRe2Dwr2eYHbVs/2uZ0j142
ij3AHcdXXXUqSO9B7hkPlhu94LmgvtQx4YTNqNjm/srtQ9/0Ltv70M/KgjKMRh4R
RqTTPIJ2+GfHmXTwkNKRA7ZoHoscw7liFcrDQCrJwOfvXYi8eT2Ldz+IIwyjmoUb
fkbX5liG66TpxTtUmHF7ajF6bwO9uLGcxYrw3iZEtzifnlPZuysHXslProiCJ8uk
ZW85Y5BVFwZ2gxSI0AsDw9pqpc1vu6ovcsesPfcmmaOe6S+EQs49XO0vHfCjHti/
DzNT9zsOk0HKWTWj6kRtDFHZ3FDGqkr6FuiADRC+fwoKWypvYax8Y69qI+k74l+p
A+rDZPaeIv/9aOrxmz1eP02W25OEbcagEw8Prrb2w7gZIIk8EpsShph6GT02jEM2
SZ4QuUZ2sZEdiGmTwJS6rCAiFrIrHFs0nCp1Dnta4Os/crnBiTgchp/f84USNmvF
qbGx4HKQA6vcUS3kxlZVeHzbVhjo8GeH4WONnLTS/eyzl/eJNTSsJ5DkZT+YMtxu
STClevxLRotKp4XBz8FUMmr0hMKZPn+PaYbd7WUppe5bf1okoBdSHVSXu6nriHFF
ARRkeZRyTBJ9c/xAsh6d1F15IYdZGvpA+r7MBAHSjRv/gcAf/fCABZdz5eoON2dS
x5RUoKNcq9QhtWDgI7MAN6rIp3N0+BwjjZ7NmaDw3OgP5ULJnXbHt/pkMXW3zxG+
4JDLTKFggVM/3hiiH9V56ewRmN6GprkzkpTRtF1mwqjKMFHlgWAM2hNth3jmFOHU
O9OYvOx9n+S2984/opEfC0B8VxhaUzlvFtAnYah3qs1dHi+hGS2sOKci2P0VH8Cg
wfEzpB+aPX8a6+3qNg6fFijEU7cwPesjQvZQqyw847opV53b0mgKwOND69318T+X
5O6tppviU4wNYT0UZcUxPiNrJjJkSQLdu8HyhNjTVOTmBucflOvhAgT13rErgG7r
xwBrQAc9GrK/7pFLyfOAn6Bk60NBD5KxKo85Xxsks8/BlgwhIR2BWaiHL7JsX3J+
C85byNU27SknPmleRZEGH2EF74fBlx+jxfOP0blw71n6axNJpPdRW79o9PbftxoF
uqANoofp5yAaQ16XGIxEMizBkh210zASLo0vcxN56LUqkAfqF8WqAIfnaF25rnf8
hOXq2ytr6x0qwHfXYp+tH2PUE+ayq31vhKjC5I3OeF1qabczsKX2Ch/OEWwok+H8
Lso5h0CUCeUHN0eoakFRAd49D2saaR3LDjUXO7gWW7itF3PbO5AwMFdjkMzM/eH0
TClVZ5lLqI/KWFl/0YAwJ15BLL++siMG6sQvBD/QmgYak+RWLLOvKghAGfmNApmG
HL2yTzWjzuZmFIa9bYeuASraoB9gnWGdlEs06kG67tCDFHzSJq4C0YSbyzVafSrV
VQt8XefLeAEamtUAL6DNCnklE9PzYjSQ6gs97Tto8Jvm01YPVOf/2982adHZwg5j
7BLHUdqiCQJYlhrgm2iiS0a2jcsAOiUXydy3UlZa+5fleSkf1h0IRH4+0THU5drC
qS1kL4X1ST2vDSQSIx0m5XY9GtV02avU+h8DTSw+n5mySydouLbgSQ1BhaGWLNCs
/bV8OBj4YQ0XCWu/TfP3mwtdzo3241iRZJ508L8VLWJ6Teix9KtJQIqPNr3TUsxX
wSv757YKQG0CzjByazjVD3Y5U5GZDqJ7Q4+aURsJ+82831VYpe9o3fy4HFPDRusS
K5epRJmowbPi1rsEAi7vfnuqya0g27g314DwnOb3GIZW8RtF4UslN561zncONxm/
0DdtRD/Y9Bkiu3E/kuWDuj1cqGl6/j+ZpZ7pJJKGIHV5g4dLe+H94BFz0w3XIxlM
Bh+PV0EkXQcmSyPGgRLsA7dMb9Hg8K0JLXjL78QVbLWsc7SI+Vu9SuaoyNKfiuh3
t8RLwbo8giBX+1duFFKG6QwVKGsr5V48j0eNx9RASWWKBFKkXWZIF94DfuLrlxBW
sCcsaNCwMG+kn1Q1U2zCIskH0rTAPU5s2dzohzUpvdLDvnPB+s+L9zSpvyrB3p3n
e/JMKwqQuC0JPog1Enm1TAYr3te/qqulXPT6HBoOtvBICgySt1jlktg/RWMoxQSt
3HRZO8Ukab9alsPe095hgSRpLXPPpr+0UGrcS/oRwvOgkq49bFA/HK9lHHtyOX0N
KLX/oSxDWJLkmrVdmdUPwwYgLXKnBwepGTqCPTy5P9D1vhMOJpAhslrvnCHVWG5U
jeBX+e2HHFmkoTMUbF1HBevbmOlca0Rgw3rhPqgccjBU3So8yAL1J471U0NEHJ7Y
zH8sPRd8gPmHyQh6KKdXKMkPscVSeOd3z702DPpdem+u9K2rli+1BoYLkGZMKdk7
VrcUphmLi0XgtpW6YGLTbiQTC+gZoCGG/67qNT55mD2+fBHmm7SCk0nHr2J1SDnD
X+WRMDV2GvJFdU4nqU2rit0hhbIa5VCgIjOjX58wWCvL1HvRBw2SzRPCrsLy9P++
tvVsJgq2+6cgOo+9T2kRgExWQT3V4u9BGQ7ps/jZE6sBcuTaNrRV4f/uxOeNSyJA
FIsHAGhRZ4VMyZ3zYk4fS5ZLeUphABO5BBfoN3WHjtaINHRE+iOQdHpLE9A0wE9h
BC5LRlvUaOtUA7TAfQcXemCKhrSoMHqm+PEL1ENH7N4ZL4x2CAjZaUil9qnOp814
sh17rNPC7FCcG433z1+0mWYyo1+7qZr0K4wr+vES1uGhaBeIHTXI5e6OkoOk3atY
oDuFnaPFZN+SFtS/Fgjmj2j+e3oOUBDtJu1L/ipa1xg76qpY3jVxzArX3ULwNPUf
zrc9tccmHJPEJ+4qxxH0i4Y9FyYt8Qf5Y+H4d4gV03Pc5ErJ//7Fx2pFxgGaJ1Ad
sp34j0UV2dww2HfYKopPRI0hAJDox9EzgpwXZWY4ouu5BGkiZPz/KLqcfDb8lVMk
O1GUToEURNDOqIZ4jouWIixtsbe7+FZlXnsrxKeZCxhKrukfiEjFvd0QoxzRsTlY
Ztwmasae6I4mmysDoBYS5UyjDeMD6ZZx+dO+sD7MSDm67yDylvq37VUqaUjN8DQr
MaWxR9HR0647Z6nupSUVpMXuxWS1Dgxm6sKwbdXallBndY0Fiei8xhlbHh0Yi79c
UC/GA1aPKeh4suBX0g+gy3Xj8G3qPNx1vUedH4UaJ2S1eB3lTNIlhMs2Tleqlob9
YttHb1PsiVmKWB6yjL+/wwI6IhPW6HBhydVQfOxLNkSSY6PO03QFBLkxDA50bPpj
Jb9BcIR0wlljPTrYYQonP9vRHQQkhDjwS2goV/LmPF4Btkj93QxFfp5CR68BB67r
gny178Msmmvcf70QAph1p5lAfcW5Mo8CrrGApZ8XV8r25GHEbDtLoZxP2rtafdOZ
pNkxmu7+W8kDFIQ59cMsYq4Z3yI+ZBMCx3wmfOdty9tngAGKldoMrA+OkP1CsWIJ
Y3V88PAToNFQSB0FJ4LUiChSoR+ljdgMIj+yi3ojNyR4TtQhwUShvR4s1+/qNkG4
RqeAgJEaATZGq8vndAQa69cqnOm1aewaqPP3Awtc9d5+jzKU6JTcGLWzXxCCqB/2
fZJlO6DZJbeLcWeMRnBg4oKqYrGojj0UUIVQxOrX9EqEqISKfrbo+F3t6adMTYMZ
GGGBw6n9lENGtZLstp0+9h87Y/7IGZzW92ZOHU6RticTyZIo3C5vNgqRRH+g9sp5
lcMS3sPRJc8xjAdWt3B/t2U6/ps8GjMLtKmWGEDXjGbX08uAZEOY3i4s9iR1N9/J
iV21aRx3fYSgkv53HmpJALicSvs9VPlKblTYmvSsTu1l0MCgCbGlrYwXrUGgEOwu
MmiBHy7eZkqlRpEr63lMsEkC+GaolonC9m5cNF8GFjQBG+YV9P/vLZaoqfi7ppPw
3ccgdNHFmrAZdXenkaYAmhWSwYT3q48L0W7yps0lWH+B32zmaErNLNRDZbI6ZFxw
caVbCgY71Ysq8k+f3jmmqW42G6JgVxAsTgPArmVc/h+DQ2MvBCO2D9T0H7p0GwcH
of1xwxnwfM87X9rLxKh13rISoWE5cpHt520Dnn2LJXj18Z6Xp9jRSqRCEtvfZyCI
elb0bsU0u++SILK5fskDoZg3r6ZtOyzuvE0Sq0Lbl2j6qGoi164RKPRlOcaozDcM
PaIXX+KEnOu+moZ1ZBs+FHW7Zypz/shCgFz0L+FRTntgVJPg2rQhcHO5RQadfXED
CACakQDpXN/Gu+folFRKZ2yqyUiohKlYnF18NN8Hix+dgYKmXrAQVB60C5YccZtm
3GsCu6CohVdIm+HRqxQtZ+Zdq9906nzFHGfnDOt7jnhknMx1tcvzBWNxeyEm8LLk
s8jsdRj6MT5n6Tt+5q4C69JlwS9nH+WI6hwqQRG+bxY7fXUcn+RWgXCKKM8G2GQr
T6x0I0od3d7Im8hXXDIXvIyX2P8x5HIFNpPLNrOmZUA4JbIYRB41KowlZatgHaUx
ssOgwwUFr5QFdUEjNmhuAtXeVWVb1jcD7jwGvR2piPAq3SnvpVMwO/MvSB37Q3uY
WsY3bnnSBUi0zhLyO46ZSr5pGKLuO8cjAyAZQl8VrAbUD1HXRKBxjRo3JoAplavq
dDSsaiu6/erJvVXP3HSaQKaj/MS3og4h1g5gYGOJ6G2BNK0xL1h/O7eyZldxNCnh
vA3QF62oCcOqulkcMaPjXI3XyUuPdXLWGi4rREMzr4csRIwiqVKDRI7sdAl/E206
+14Hl2XN9itx7YrI7VHbo4m4NNAfE77GxtGq16pKfGyFkEmiY+eup7hGYB+BLxlH
2Osq5AGA3r1fMk7sd/MMt4tJnfXwjfQU55f1BLYGjpHN8U5H+aCZ4s0mxyqaHjFM
e1IXyQ9SujANnFWgxeRjFEHfsuI8nNg4OXVjxvP9Y2GxRS5RBR6Ei+Ue0z+QcbzH
1qW5skz75EIJxFpqudWHnRKigSLTtjdBtmsAIwZsKlNrhcmk+Q1pIGdWo4M48YKv
jtBgzcqB5UjdrFAVKfbx/FN5QiI1JwPvBa1sD0Bf82dWmEd5UBEkrbFAEN9NeWYO
WIyzp54Okh1L351xiZrPQ62ybJSxrRpcyN5lyAYEDxD6mCRaekp4ODaEITGraPJm
+TomFSYe6OgGqVVwp7JKzwRm+Z51Y6ZHPgu2+nwto4X9XUoOLOFSo9cIc6LOjdOn
DOFF0cOxBHL6Zrb5FBn3H5zUTDowC1vX54JExH0WG48ovDTyMclPFjttyJFxeoeb
VSIIdnr1q9fjnEBTNQRuEkdcSOgaLrxWCgq44CPCO3TwmZ0ZwGIOak1O3d4yXx0p
PUeoyDcSfoQDkUNCdwD9EPKTAQk6QCvKEQ25Zdiy8x5LtuJzrWw/iYuU+MPRwGrw
g9KtGCKAnVwJIRzw2r6hJrza6lOtHrpbbU/+czflJqjZAaNAcnj5O2DKELN9m7tJ
8cVOfGGYNttL+dxKIkgWygPSQwaPq9IdMUV6S+e5GrwJahfTtBcxo1a0p8MxJaJB
wr9HYTEz+TKmXHqx7o3kmDBPmqlW5S9d8FCaMdNYh3UfPhOwzaMrPbyZZQkbr4T3
bAtiiqPHNxtik/fWDML5DizCrZ+oKKo/dnqez2ooSqeEbDhtXJuMThCODnlMXfoN
IvnwOnCUJzCUGudocRyOzK1pv6TAHRTw0W/89jXXQ7XnC2RZxPWgxtwQ08sAWtBO
5KGfEYV94g7SVEUO4vXZhZ/kocfHtNius3EitBJ/+ItsMhTUzygeAE+rE0FNHorE
C3HeBrbh7hLgY4cxmu0bU91Dr9u8Q2oVnsnGSV9Qo9a+wbR6MYWtSLkKN91V86t5
urOXEoYQO3fuTTHGi3UbBwdrDCkZcTfQUWUqpV42cmYSwXuhKx2pQXlwaJCXe4ee
C6b9yvHKYWWrYLKBJv+wZG5wm+5kRND287EDx6BFzXV9V2Hv+isP1vRBwhqZHMTc
MbYXIcXd4k+RNi5Vr3UQijhXrvOc4ENsU1L2stSop8LH4pKCkmbzFJQKZ3UlAZ9C
cHQ+sVf9cWf7jwPIcAAJtboUsYp6I7KaeRgxLHNXKrmfW8A9IvDXVHTMqADWYSYt
hkR7N6Za30tTFceQz6coHZAZ7it+ED0GYn/f8jKzmk2J0utkZaMxAozLdCbWZzJD
9qqZXE+CN40WWUb6CpfOfJm/ikfc3DMM7e1RRQo7ovU+Al6bTOAO0dOfHEjuini7
R8biYHYNPtnTsie+4arIIOTVnCpaJpVRjP6y9+/AjXtcTqjSARb+xEQTcVFja1AL
CPMePZb5mZB1jMDxh1acw2wfS3uLinH0b6wM2MWYNjDp5RQPjE2+nSD8qptJC1Qp
6OVyAzzt5eXKjOIgOH5P/4pjZ/oX2zzm2c9V5/CiFx+8wqGx1svSDhZTV5I5Hqof
RUPh9BiQ8KmaG3tOKaZqmk5uR2tPjN2/g3n/B7BzqDZhmrG//tbdbxsfDBs7Uagh
k9xZapvcN7d+/R598gZOkmxD2GUCcB6J/n6q06NUT/L4Mc96CpO7PDpwwWPn4xpV
xqhBucqSeL9CLDAT/HqpGOLxcElCdyTWUugSoQYReLtECxSdpjGkVbPFH0WyUnNi
3nbTSQ+lRfIjMoNHWQ7L/Xqqe4ONyJC9CfxdSA5g5+EeFVkQYB8/UY5UGDa/kGbP
y7jw1Y9ybWcMliKiG7O59BIO4d9juq25yD/Ge4fjb9hI8376t0/xxHBKR37r/tPq
9PqmEslNnz8Fjvruy2TH3yyOkAXc8E8SP2VABqMveWpPTFvKwLTcsGvXBrIpWXwt
PACb5YFF4UslUaE4Ta2W4oe2n4rpCPNEAQxTMiLh0J7qXuylGaI4wlicWDCrAFAI
AWe9dmkvXTSIxXs/z5G0TMmIvV42hX5NskrZPQsjvqo4nLnNPf1QQq/S4Jd3rB6x
gvQO+nM1STIffFcKaspA/oLUlsJTEcQCzAIFw6nsYTz7GGYXe9BJe+eCgy/iA+SY
cRo1dteq+AshXi8+4balP2pSycX0Qmt0+Ds1IZ7rxUelWKl3FHdpDwgPLKjlVq7c
T3cgGQ9wi8NJlxMbEX4Sg4UQO/i58e9ydtRvYI/CgODAPXKmEfv6RamLR8yncFst
o7KV0uW1wvSoDp9dGBGFlXcnHA+1z0OVg2INMfulLjbuo8xKNKfcdoh21m+JiVWI
jq1GGloxXiTsKKlMbHG+Ai54JrX4oJ1d7vE8LMwoXdS2ByyPw7HnNMSsitCdan+9
FB5U5nBnqBpajxk1rQ57iVwwK6oZBpB1s4vt6EjeDTExu37rDzHFvWdoOVDMn99S
R9vxzohQwYx21Mi/ovS99KBowOEI+jmoBY3dPGn/6VKu32v1OiYhFNncicQneazA
GedsCtp5tXfzSW6CrNsSb3pRVwITX9PtelOi8Zfix1UIWSTTRztmy6LKOoqz8jgn
nbr6ltqG8wBpCQH5ZMmc8M7PKvDHHdjS/01gZSAuXHAol6B1O1HeIjFBuF8/URBR
eAXzaqT3KnqyFNpFgdCkQpsUvRgdTShfZytA+xXz3PlQl51UKqooiv3phmS0VaOn
ZeS+bXbTtSDxoBYOf1H7sfs5ElkRSd5V58So2L2ct3K/GKkMzPG7ABynWfyyejvm
g0WdOz7uCbtEVh+KUUl9KYHvW7enIt92psyF1U+JfyUfTntdJz5ZuO2pnGtWPb9D
C5aTaNxSCrmXI4RPXJxe0sB33VGg75jM4ZD4jG1w5O82JP4KBtJiMvielo2TE9DM
OQixiKLipVL+pXgtXzwP43LI0qawjuGjRIQuS9kpD+Kui1q6Y6eJFyMA8qdS/uGm
B/8wA3RjY9dZ7T7fPBgedVlmMyXxwggxBV7cv2UmCjPYYErzx0FpVOCED+ilWxGz
n4Hi9sBARJdv5/IY/HNpkQAwHJADWu3r1Y7E2meDD1v+e8bG+w8ia6XLGHvtFz+U
nBLQ6MTu1sPx3mbLw28Ujgf6Fw4jmDT1sZ2JQqHY6g6vVlCjz1RxUBhYZO5BKmH1
BDMGbOP4at0JcLsYcA7wnNetcF3xW5yNG6jamjEDWvH5UiJQYlr2QeXTHWNRFm8I
/dkN23h7l4TSdBphpcqBcXpV9WdIl0YK6j8CYi3qmNxcauLps40lBwViKZWpwwX4
u+iVPXwUq+SYhmCXOcHNiC5o6HS4uYyFc5uuvBhnJTV9W/UmMf9TjJbW/081mgu3
6pBkkeXV2YTH9X7M7f2+bJ1pmacgrLVzkXYtK3sTkjV14kRRsrfBXF/oC4p6w6B7
mEF2Gw290BS+IsM+2WyOQP1ZhDX/jWbYQVCFG3WXS7YSUUhOBunFcNUBRYT8uR2g
PMnFS2ojGodTcoXe87559+Y9/itSs+3PdNx1kVTAx5PtljQGKNF7hy2pArE4FiQI
3v2TksB/vAiySqZ/i+khUXcLOusr9m4ugtKpv575UuPahdoI4F+wjbKsUM6pD0pG
hAwzpRZ6AZP2jEMN3OY8mwr9apSVnRtclJdoKcEVdFQJMWd0lv/S6S5CdJtzOSqJ
Fc5a8B8X4lLz2YU3jw9kvr9beU/2FKzJxJStqj+5RTpHvqJCPmU5C6iP/aGGtey+
6On9lhKsM5pl9vc9q347k0aTCPCeOO+yDPGD+D4OiKopttoWCBiYlxYU2zICKDeK
RElc9FHiyQjd5oPIfao3mN0bRBuO24r5ZLR8NW5R618zZ4DHNVyD6dDk3N7d/WWj
Flj3xHyFU1Gcl7z355n4wAUrBjSDtgEMSmK3LqldIhpVVZcjKySlZ1HMb39VlNTD
EjbIX/CV5GZYzUrbxZndXOLMPtYGrRlaFhHCDqO4IEChcolacK52OQ4mU7zu+OJt
FFEWK196bZZC6kXiQrBm5vHkF3TeNYMgjEFSdh9j8ZzFSdNA9S2nkud4tj00D2KM
fpES7A2ZmztEaJo79hgQrAR3n/Vy6HDmpfzS+M5pabYfJnVKilXWTZZN/K0+8AR1
w+KAsJYpz5s25RbfPAMO/InOqjklKIDbu5eHUcTrHhiOuPitTvkOHwdujijzDQDo
zJmxHNdRi8KuhpISzn2Sn5V0FL+v4Ndae4w2HksKTR/0bZWFEd47SvoglQ9nQy25
vkhB+Lob82hEFJW78/OAnKQnqLKGS0aQSeIMvLYXcA4Lfk16Q0Ziq1ro7TFSjo6B
Unpc5iYS4wrPBxm+mnpWcJUZ0i5VpobS76ujBQ7DfkZVerZAGuGU8JNQpozAySzg
9nsTxMcA3y78HKE9GnJ/YSLItpBc8psmm4HZPUkQ+FbD9KT7GvBR+JCZQX+l34oF
5Nn/ATQiDEuxiInJ4oyhFnF3q7k7s4ZubTc2zpW7vBN9HCSmbI42eThKYJ/Aui7U
nsm3zD2Ht+0dgfU7PZxJEXETa+0gMKAjABG2oibCrzp59dfWie8k7wcpgKwgu9A3
EE4d6yA00eY+qH+IYpuoXJvzFdYhVyfwQrIi2tOBaLKYfPmmglj+NzX4e9sxjfcU
N5vOqKz4OAMP5voo5SB+UWuG0zF3MWhLNgMBUjDc1R0wNYeegXXBZcydhZ1GGkl5
o3+ykCozDSjwUM2EA+/rg3Mb7+cni+IP4+xAE2raA/4+Z7OHledxUQpfxzLozCau
i3iG3YU5M7II2JR0UWl5ZlCq8Nh/QL7AbV+W5ELI51Nx1V7G87cRQoWEHGHZU9RR
8cC05qB8jsg/BlBgFo/vU1EuaRTh7jRIMyCl+1+0R64dckl0o/PFxqoHDBiB0RnC
kik7+gcBXVLP57HznXDRsaO9+uFiwRe5OETurFPWdnbsE5sALGybyx9zSQ3y6Kp1
eMY4hSNTK+PyMt1UPNLvTf//ri7kjzAjKlZ74hm3ezrsHrfOkOIEKkBCfF1zrU0C
cC0ob1IHKbNkSI+9kpiILGrkGg8sSBCzjF53Ydtrs7CDMDhGTCG8elmyZtrU4BPl
EJwCpVuppQ1/vJJryo3/5SQW0SZxITKJffO9rK6jvXYWQVLM3tqYnZiBywIhhsHK
tSRbP7aXd9Zv8QFKcLhtAlWhbb3jNTB69n3OOOzFWH+VwXSt/1OH7stUIfyxFKj3
vm9dXoC2N7S5eR3ZCcsKx7rWSI7a3ugbI9jeE4yH+2KxImdxfLjWdzqkKdc6jpRr
/i2JAc7gsJotgc9VfNiphJLEDJbiEJ6Un77fqgsGp981+LmFGZh6Y6x0S540vBn7
L6pFLHCVA+x5VM7GU00vfawgmgKSRyn/OTuUZHIunR8Z65CbOGD0fdfsY+gDAksA
iWkAJhA2SeIleShymnLt2jDHjvyHsjaw+g7cD0tIV0eNeCPXCwKD4MY5WQy8eXNk
Wyi4bne/3bZVNKStdnFVoYw376UQrwJwlafztmxIJoJCKIZ0JWUwDaypjoGraGL/
Uk8HdY/jGcxjzRUafB8SCgbkAMX7lNbA9pNldMzEsHfYVM0yoQQ+Yyt0Yx4kFw17
ih28HeSTV5/So462Psgm1TU3bQhBM7RYF8lc1rVj8Bf/ShhZpz0N0VFa5vOy8iMQ
/JsVky6lSvnZYwQxJaVUMoZDtfe/yYHYL8sJ1Pz+RF+UeNgyotOPNNuSPq6trZi/
tPvXCZE1WidlowfIPzLBB93iDQaI1yHJ9kLKfDpLdT+izQc4c7r+a98vdWG9rcgw
014qYNW45e28TOCAJ+xpKsC9TXwpkCKsreJbxLPf7bMWHwE9iiuo6J5gCASSul03
JfW6KwuMBF0qqc3FriCySJTJbVoZnPK4B0a9RqIbeqHS2oOMTXHpc2BfL4giLYFk
7X8pufcMdCCjkZumBA126hx04A8w6PP7sqktIqxsc5fhDRLeI7I3lVZkQ4uCXEL7
18rZl98Qgagq62G2kzClFNtDKBcs7Blf0l5lMnu4Ez6DCN7wRCe9v4NXTVcKtuoT
Lkm4pAqkvJnB0molOJbrkv9Ai3z+19j2qgDDUP85InwbsfvIDmRY2SUGbZF7fvjO
3wNycily0S8DMPsvocJBgN9G2SYSFhrSe/Low5uj5SKnDHVHonD+muPtHjfSuTVA
ttp2P0RC0mVxNEu1aLDmfb4wz3w5C0y/J3jTG58fX9qrty9OOqkMe6TJypHYs0PK
FPOLfSLh966rvE6VrUhVlVipalKvwuFbuRt6JE/K4gYqKaIoczw2DRQPzIOl2R2q
4NFgNCyNSxhcF5HehoO2zgVlz1GxGfcS5XPkqWln1UudMD+yaupE87b+IdIEPB2I
pLx/KFkzOwoN0oVv70zW6ytwjb6dkzpV2S3WNVr5m0c2yK4JYlRQ2onSOnKzshvk
q4CPCiRmGNsgpmt1q64AnjXgQfsQm/qB6no2vTD736ntCYJJmv8M+3FFeVMGd5Gb
Qm9GUNv4TH4caRSGSJBtIwPri/zcZWBAXXCL2fzcAEAvcjvIAxHIbiKJJgU4KHOr
I/SNj+oXbRF+wE7Mek+Jxv2npTzWvxNHvucbTmk1GUd3pxpeKgruPyxYGMCFJxqM
Q+8jbpKJyluSrMUkTpNg0Xw5GA57r3K0F9Q13TWUZsXIF9gYy71Ig8UVYLu6hym5
yigGyFO5Azpw/bqhrC5akIphjpcXc8k1JIS3zpS99yfLi1GwcPVI8hxJJr2svvmG
RheWPjqYyoE64sTf/L9whqIRQ2ErST1a7alrkMzaSYPGyNEvanrXRQNWvxN/Ej6J
c500NRCDfYxI2yC689Sm3GuCZHRruyxm6JEKeko4vuTMoCn++Ow2DYOEv4sBn5ah
jMk4PvP9pnJQAtidoKiN0/W34y9KEibYebcXDaXoMoQ/lTnDJ6XgglGk+VDwR+p/
1R8WGKcSoxOx+4fXZuNTiydAjqUy0/o1IgDsr+fWIQ0k3DVbxeTf8DJ0UTSXTL3O
nKrZFv8PzdQ6hNcdtM+OrV+JwGen8VBpt/HRH/EKP58McV/M1klRDE69GINRRKub
11z8YC/fzkLazQ/0WJGtAtU4L2zeauAS/8+/P1rDSBaFcVua01JY99C0MmfGI/Vs
RH+MNxo09LKPqgvCOwIY0vFSrM6zMw75YHCE0HiVXOR3OqI4y+JKE3gbKc4L6r0R
SIBksIQRLUl9YPRDkynHKRe2NwZS+8LQGgbRZFP9JlNROekrpYoQjOOceNvqPPSN
slFhQkYVCtVF0LMQb4bTYJohavnBp569UYlIIaV4UBMOMVAP6rHJSQ6tyRLbKmBY
iRGKsUc2nK42Bp3HXm/oc5Ax8kPgT16ty+Ov3bac61XhV2+Q1jJq6c8DHH/hPKEw
CfGP1GV+Q83VXCVaw0BOSibxyyQ5g9Sjmj3YVlfijFkIzMeVXSYgXcE7qZI+oiw6
SFmRvQ+JohL2yT+0CZ4oMjlAlmQw0S97kuRkbmdbt+c/A1T1gMZ+DdrrdoZgD3xw
gBbiFRDa4tSKcp+iGDZ3Ip54jZrsG71A0CJ5e3gXg83NR++qjfb9pGkLFHORolPq
rGy/LhyR3Dal9utASZ4N/Gv9H2be8CnELjrI13J7LysVxgIPIbeILzsgym6g7CZ3
uLiJUINGcYNkrS21mA/GjVdxRs5sLVwiAKd8LnDsnV9a06wzJvJAp+wLZ/qxLH8z
H62+612yWYa0qDplk3h2k1ZeyL8Ny7xByD4e+mNb5hDErNrbo7sfcTIB3RjK+a3a
pVazRjwAXZuNokZD8u4PiiN69aNnBknQktO9RIpV+Rd4cHcCoNG6g5yCC5CtjdM7
6mHtpSMQrpH0AjkOYukyBe5meT/F803fD3wQ1bMhfXPsBRWIw21bjHZ+wOBSxJZm
544wjmA/Zea0mGhwuxNF6RL0iaWmCu33n8d3NnrzPs+wlrN8nR0ClVW6QOQdPo67
FvNFAukzjjyva8LaHipBD0/HQjNjQoKSx8QggWvK/eyiTh0/ctkP3J27wH7Xw2rg
SpwYBq0UTElm3hQIQ2hIz6AvYCJoKghw4x1mGxx3UFjemP4RtYfeqNJDuCbj94mc
rEz/q4JjjTTjiwlh+JU9Ys5k68bSzTMfghYUSpI7VN/Y3JNPShZrVezKxChfWSmP
7soK0KZxPvxHpfyW+cef6g6R1xleZeNVFp6KIck7JeHNzMptYF4+3EiW2XJJq2Wq
vncJWRQrK6Y9EcmQZ+OSXmFgJF4tLqLPL0sN/5UTp715CU4pK8bvdLWYdGa4ZHVP
A6mLmlkEIzcAFZrSpgMNGCD/e9EaqkM1RsFj5T/h/F1XhpipbvQTV3xPVgxChpU4
zTwQqh1gAqljnmRc4/Klts+64LRCYDyp/+afedxloAOBvY2WLrZD1rqanYrTkqDz
BvYxq2zSbs1Mv1ncOF7x0hJ/4JhjZjCcjiIxhEFPh6QKGLwgJfCK/MRE60fzxXAY
E3COQSeza5A8s9zI/dvfRiLPCRlRqeBqCekNdFmOhxZbH6aYL04R7wz7MovafgKV
0d0M3vuYvq7a2W7pF/z5ayeerUflAC+xbCGBxWL1kckSgUIUxYm69nM4gE+u+2bM
a0tUYkZJqGIXcpJ5hGYDeyJF2ofzjPc/k9bGgwZPHVCxTUWomaPFAH3SAmZ7+eVg
cWJo10Tudk4wuyeMCJ6w+cDQgLgYg3iZKuCi1bYSmTc8liAjrgJ4Vv5JcBwNWkja
qMA+RBsuGs8974xFa21iQRbYR7XavGpYQAXsJIfJfIjMjyNueiHeIcdO4PMBFfhq
EMveSMkjLjHD2aQFnjsflFyyvDF6GFrkLwvclw25Nee2LIG8e4E+wustBwFlvGnp
IcvQ57NYqRJ33LU48932XhGI7wO9dl3uZUHwmOFcRrVjdx+hNxJkGHseL/sPHmIE
LFe0rAXDT5qbpAAeutIUoeS8GCuS8J8U+j7JKCjK16HAf27ciVb+8MHPggP0Kavr
bsxiLnmoWYyBIImpQvCLjNsUAs25DdtHms+TL0DWQ7f2CCVW5jy0u8t+YnXZMQtN
eR8eylK+pUcola2zAyJMj6A0TVj+z5ZTt0R54nFxbh2TBunB8moCSMzw3LEAb7dy
7Z+M0XYcFWSKOxEmtS8Zmjk9rqDLlAUWvXAseCDBv9zEmY+EG5Z+MdevlK+uq09k
ddrwyfmxC4ZkyRuibU4Kmj3CW4zseBeThxJ4N+DDq9GO+tzst0EK1HcMBw1dIA3e
QZbQ7VCijzGKIZkK+2TbfQY7GUs5vLUWjtfDHtlR9RnXmkUmntyWjfJmSE+UTUSm
mfh9TPk/3v8bT7qtVrt3UWfIf2Ct3mgWKiEQGo7daJHxmQDC6lSklHm/SAMYMYNk
rkFvDa6AtDq6nRlWOf9U4o1JNqPBAhalj1NMKrIlv1UBFnjYdY+UZO8J8rlldBwP
arXFY3Wq2JA+P/Hb0NzOxFW+lWb/NY8ZuFWLRCIuInXf+88ylIoefgmZI1gOhnDT
/hOXI4doumRrcCjjtqVuK82FYb6e5n/JpelubydYvtZnd0zbPOH+BtnAknOzpzKS
3mwjGpxqgcDRur5oeUgDrVo2sdkVqoIP06Vu5c7VB+KtlVgwojRlTn0+Mjq/4JAd
UsV/5L1waOovSCeIjoTwuaF/IylEw8oQbZfoVtpvVAFktNDY/9T4tn8L3KyCLiIH
+8ChLVBH2ZezYx3yL3dSNX9AY/biBBdc8aLEkDVnKjtb+dGgUcNoL1R/gRaxbxZk
FG2RUaHTCXEvbrQKfeDka4UJBVJjg6tEO/gQUUvtPzCJcSgy/tzNPTOl501GxN7j
uxw9ZaZrGcIIkjFT1ajCl1MrUDWjoTnrQGhImQIpvovEywroJeBnfelFXK9lJFDP
tUvk4qA1LmfXXnCCbqyhueLiDtYujNOjxo4Mpow5INGXNBIjRbToGS3a4G+M6mW+
5NP5ed7y0UPx9tm0iIOT6c6aDDTsPC1JoG2N9/g69FM5TnOmdjHXwrkk4aFPHcNb
bsQv/fcOplnv8FBEWOW/Agaz4xIars8GbgsjY4Ov00+u6il4ffMTNPXdJZfAVU/7
YpIko/monVAufV3iiGwc8x9QkxET9MTuf5ON7kn4Nq+NOWLAdzS2UhAOXBpdAHXu
iSzmbe6wDvAsHcPzJUICcObg93JqJ8DpZTcIRAwuAzZOkYnP3p3tL7dFCtxJg2xY
4mqKUj4/qcn66p/JhY1TX9EtdbMOmVxT/p0PdViBXDcCTlLj6xSujo/R9tq9L9eb
/oG+uxSF2g/wn4GdFnG0u1KonRYkyfFQPjNfvqt/0sLicfaJhhXKhZi0cI6+Lfgz
AFnicHVkrDN9Nk2f9+5JBwVExDIZ9rKw6/maNaIe9ihUXnEhQ7kOS0Eq+Qy/m1kL
ZCe70UtV4aDnOYVKLabMqYmoiSccIYXDFBEeuiswsu2AB5oE1TGgnKQEBXmbx9lu
98hgVn6dTN4IBoxDNvfSv/9o9bWeUSzR+hql1p/7juwc6C3N73sdZ9GESIBInpW3
uUzyllvcUYJpENX5VRtpx1dgK5tHGxEG+3hi8MBZ8QW/vyQJsIEyXdVWBFpf72OQ
vsaJlF4NVCteXTYVbTUe8FGMT/3eUH00ylNVsHrfbJtorZmpmpMd7gj54mP1Sv/V
7SUxBwp1KjHr201YFSaPRPWnszHhJkDY4TLcJYVQlv3yulgJAnF9mvWzrL8gRb+C
h8K7YD+hZwH4ron+XZhm6cL9K6j/9h3P1c0+lFtXFfdxYSfXJG2W04oOTt5fCLoK
ova1FUqDrPNg/9Nw3yRIo30Ehe/Ev0hxbZaO9LLXFvNdFNFomyCHmusUYO3nOPWX
w4O4kd584MHtWcMhPPe5ozoLUBrfY/Y35u0PL1r7idzkTx1tehnyEy2A2Q09p3/3
T/34Gpj8nkoLgwcG+uXIrTK5xECB1XU9TsvZLQe5a+5yHMvrhIBiKZpW6zehzkaC
g6hYbHr2ivtd0Q3tqdtip28WobZF/gZcRdzQ7E0pSlhMXbwybvZmkrhKr/p8j12Y
YtmPa9WZQPWHwuZsCjZebYTDQ7uV47bTxQOurTign/a4KukhpC6xhgJZkuT4ldDh
Twu8CV+HuWl8aj6rmljdUMiE2VIPuiuo+5FIOY88e6/ovN5hG2GxA4ElrRh61sQQ
GoIosveF82E94pi9J3uumtanHklwm/vjHkSdKz+DQgTkXwo2rsNyqAhc1XZcfiJI
1NnkeHEjQYZrKz1SANzYOwLp4NjtFMrmk08kMWGV7XHV/G6468omfSjJnF5ranpk
ssFIsCTDYVoMDTcj9s7AJYpyrWlHmZwGBL1rYex86Zc/YZoQa2XqmCIlDNn7OE5e
obEP80Z5kBQeKZ7b5rU8L3Uy0BQDHDyhjJyx2nKdyPR5fDnsEKX+3/sPJembPjMZ
K1PydijgXRqNJNKdaajK7mQAL/JO/niACWz9QaD8WQrzTCtohjqqqE2Izf+fr3Uy
oWMhFHMtpfV4bUzBjLiEO470KzVw9g6xs5+WH9A6VEsl0WM0k5xUKxoK8EB/5wzI
PCNw7TnH593+0K+1b3bUwggG+UnpYw+K+XV/J3k7sFAfR5VMuud+3PAnYBb4X3wz
LnXNZhZIUK0EFWQ6IooxEYPILmtdYgx8hWcUkdyCQvx9Da4UvJlJzMMxiV9Smyvl
w2T2apEYT64zB4klQHubvJRLt6+UHoUEu52/moDb1cuCxpWDLCgEuiR9F0l4muOr
f9GcWuQlLxfBGulvAyvARtocPmDA9H2wL1JEGeerd6obRTl8bi2S5rBRVPlp/Fkb
ebis+w4Ta/tJUB85VWlPrYHlHSK4JeLpKlPcZIqa8QATaHnnV5mViQuX8ttZEz/j
4j0q5nad6uNRlJBQfkCteqb6SMiKPMYcx9tPusPx7OWyZa8bCZTs3FB0wrl+6TfA
xVm4CWlS7hlqvTMH2KEepSVK68O7T30HmtaaCSWdDHJ8KaUGfZhXNreQZ+3R3CJP
Ju6w9LMQm6VgFWM2l5EddFW3kUc7pkQBK9Mq1YlwQlouoCIstEvMUE17pqwEnKJy
qFkF8/7gVkoXaMfjYw2MXs3HtOlum8Xa9cPPCtnqi/pWtCF0sQIhH9zlHGa4a5jS
pxsuVS6seRYgk3N+gdSf4E2gyJvKdGzhjdwAMFqqoa7q1OAp7jRY2YNxupPmFJL7
ISMQrvFf1fqyN0e7KE2kBvw2fTg0BNrfAnMgb47fu5YgoDQH1A7PqcSc3tPrkIay
abMzQhZc1TcxTcPk0wBSvp+fILCdvLUrevzVlRnxQEBYnR3v1FDwoM3aFrof9Ksy
laE7BGtkLjOLwwawj7OHebysLFpjRrAMjwHeKp26q74DE8nWZAvO4pX3d5Nzr1OI
p6SlwYLkt5XqXGk5dW3yBYlK55mW+PrOt0iKSEMykrlk2st1lcyQn1adLuMUm6sI
51nPRFPyds50l68u0bTh7+ZKe1SV4693kHPleCo07ow9hLJnX4rMRBafme47XRoq
KlbdiLEAXgA5ejWCabDcWyC3W0pCp5pcygoEFZfTXcPOmn+2PzbkGM+//ARGD/Hp
m5Z1l8ek81VdbLHf+iDdt0y0Mlv9IkdhLb011kYxz1051ZU8FSl5mJhXrCR22VJy
E7/mxdDazabuQc56UXjRA8hKK6F9trCeAlY93FE3q/0NxQ+3MkPHHyqAz4PsvZ96
GcXs4PJgxd0kSVZ0/Bb4BHXkCvqWr+qK2qg/MUkYemAy5hqIJKlUHGuIWmwaPcNj
oMCc7Qu0eYhaKCrL8x8r+MI+YBcS3/UHQGDVdE3Rd7/gev3o+ASNbx8wuztiN699
AHDCEzmzFMNNStUHyIstw4irgga46P2J/BiVB4rpA/R0oyHyXnVhHhmbTuLdSxa4
RJA9kzkgDKXPHMw59OJb9qkkatWv2mVf0hbZ4VUIphz2mGg8jQ8V7+oMDPM8S5yh
tnu2ZwsT2DLvdfr6VdWxzUxp77YpfHvVwX7XZqnlJMjgZbLbdu0aJOcNuhu22HZf
SctC/1US42v9OgVzA33aUAP/6oUtsDpjNGqy2xFqLSBbwX6MM8sO/5m2IY2a3kbQ
gRvYW70Jdf9AClNrmiaoZilvKYm20rJn/XB+PY5ZX4AmcfENrvfnbMnyHsz5wwY5
vP6H4V34sYFC/4IJSkPXTf0fx2a3toMltv3wD73R9JA/tOdCB0aMKYKMb/20nME1
q7SFwLZ6bRdmf68o01fsXaqtg0wN/ls+F1jQchmlr6KuNyX8jUWm9hRkfv4TDOZ1
9HcWJkscMI7u+JleIL+8xQVpkYVPcdPLYCA8RQx6Nuwy3Iy4SN1H/YCOILnrFTdp
b4Ak+Merw0Hr3Glwq64WhYQqnIQYEBPBezf/9aRZ2Hu8W8iGdvYx1ye9FfhyhhF9
GUP8wOGEQ9OGbPia5ulbWjyyLUh200qGJAZHhl0DEk6VTNoM7D5w5Ahg5JCblrj3
DZU5A3nsxC315O/A3sbfUPnbqNl/o8DIxMf3LfxyylYTrbMCVPNNjycoTQMGFopo
1V/Kn7LK6gPEdalq7HDQSGRVUROOLststJut9OnjqwK+Jifd9C8MRKa1JZCBjAR5
uNO7GPWmLyMdOrRfFc8yq0O7Sh2JgpoL7wEv+ITYLvL4X1yzevAknH1J1Kh8g5EE
UBIAgyxXylcY3RVIUUldZpdZnxPgttJR6NEMkcWVW6a5YalrNExKp8o+Ve6Ze5M4
MWOAgeygNzSmDdakLefa9BdNKeeBVLTRL+xyQzQBsZiJ9olyTNiTHzCeDY+sFmSt
7Waq8ltqfgBlfasvzUqCb7b4vS1G/+UaYs/kATaXwJZ4Ax2DfxUwBCiPlzIxjNzN
/Zcc8xzkGQpamNjjvC5s0ExCkJOjTJRKid3xcH5ebcXdxp4fzJrWoHFuKhMK1xAP
CUkY4OD7upwLyFsyULwjYLm5R6APoYlXGAjNceeJ0doraQXdL/EV4Rl+W8e4893L
Y2WI9/JDbvpYZe5mLRwhJ5r4p4rFMjVvIRNodptSAptVmH9K5LFMUerXzrgnVYJz
JbrHxFxLzzy3iCrPtTQ6UnirTwoFgPEfqLR9cK1mJldsXolv3WCEuxu35qjykiDq
3CEQV0zWxni/0grNW4X/65ANNOOjbQtjkuBJzjYf1SIa03loYk1jtl+ShShgTeUx
OrLLBb0uCrX23kBQ+TQbPUvYUsrMmE69SnuUQwrFsq04DW4OSiKPwUKDdvxlvAMb
eJtLqRz3ey85OhmNhvUmx1WRQMJ8MWySXE5qm8aGb4qHdn5XGKZXT99e/Ofyxtxb
g75UOSmxNMkglzdAzHzE9NeK67heYwU2pDlr2bgMHVo8M3ndvJO7WYHdPNRPh33C
6+0u0urD6A26ix2zCupWVTXo/paUUUhgsteMb45Y1ZJC0Pv/asHGDHCAe+TfP86u
wcUD2724MDYCNkCQIzF1kKhwH9ooUMnQGapLWkJ+5gHD367Jp/vItU373TVbyqbp
aqOIifuiqsJd45aqfsKaYLox3IV1liHecN/uwJxWlssA0olvZfO0SoAWcKB+KYVG
tjInOw+PPYB9vDGIm7tWntpD4WBRzLuOlkLPKxph4STKjN1+Hth7E2EsrfgqJbTT
TzzbrYJB3hcLCxYLsbCF7OyIeIQCuXlrEvglQHO/L+vDz3kcJeu7RWpBtgyViPAU
jqlS4YUFbQkVIRXPtKFdwwSQVIdJkg7Jb1l6TFcrisGI/lPp/pc3mAfo5CpiGrzt
MHrw+OdVV9YbM2uaeyy7zYs8CGjnsXLLZdahhbpn1oc2+CxPUGWlC2QRoxYHyc3E
TIV9cpjp3p3sWfw1ZfabnQJfTNxCy9vUlbotSasBhNw4zOcgmoiwrkdl0uA87PQd
d4py2VfvOaOHPHE7rCIX8UtEhqvjErFYDAWBtEH3ZxvCZRfv+nw0dckocr1cYff6
KG292uw7gqXrznyKTZAov8pn/5JfHmbtrR/t27XI57l0bcg2rKzxu1FlPNNjn0dr
nzyCD31cN6olC5fp4nrVFuVD2swVRBQISBpF8V+POkjTOqJSwkr5sYIb+wpCeJgA
BaoW49Cg61bVjG0hgugxmUGTM0LfJhBRrfOd33YODZhPjnneVTsFFhNJyYquJJaX
I8Iyk7PDkNdnasi3NEaOjBuUkwZpRXdJESM2+6TiGAggN86s/XC9uZ9R/Ha7onT+
UsuSF+U/X0eA5mymrsEKHPjoNJBMyQNiWtAxCTtVfj6meZiuM1+jdseeK8JQOCdr
AZ2R3f2fFA4epDgVvdibzhkGKobho4PJUM1y4iyHmcK1GctaubWhOUBR4zAm+fm8
Ngru1YPEoRM10bW85yHvomyT/3OEAqrRAjUQ174NdWMRWnVXEmvoQVv0X/byxA+N
Gi7+eCNYLO408v5A77vgKYGDzN0pTKbrqFXdxQaCQ4Fg9nNe718TmLzCvQQEcuNI
ChcsTSBZZ403IMyVAccWzx6BpKvu0GzBEhAbhe8hMEKtTc/Yd2aiTxGb2pxvAcI3
/nTHLGltucAzOa/OMmjq2Xe0JVvdMoThX745LRJxxVOP6eTczg3v2mzUE+ikBkX0
WidVzcHReEhec0JlKQdVoKUGUTbIoWWZQR64GQ3V4oFRTSTNnxYYxd1HDdaN3beT
xfXzDJWf6p5n5+FAfWlodjSE07gE8LZ9eBGtgj5Ncy7dM5N6dSz4HdGt2zFzny3k
hgdxTF/1MciyrLMYYlOC8O/1jTHqVNHk8PiuI0KQUwtfXGVnqSpMOC76mzKDMfKw
zEFIg4dffxC2+/JqoVVbZOXOYAot45QhZeEWUcnA2D3Pl7pvHikb/L11gBK4ZL5I
Ft2A3ZJWQqlyVE4ZUDP3vhvSj7WpnCDqKQBf099foODgqi8V6FE2YQGVeqSbWsG7
GgPpboH+2sIldjqL02LPYw2zDfJMd+jtuqBUXIrDkrnpVClztVJKKSb/7HQoPDNB
62EM9wflXmhh4I85aSN2zCEeWt3KCHY7qt+Ntfjgj3WC+ledO0ruqgVPteCP+BWz
HeRNAhphNf8QNEu+hI82IEy2RkgXGfZ//QuOvEJAl4XaqpUMBaXckObd67Zmn1Pw
z4xLSnt1qiT8RpwO9cTyRGE5FYJuSzUqvN0UKWrVeXm5ci/5O7cPNVgq04qrCniV
OeT98GTIIMZUo1daVA1kKgGVKzG0w/JAImHeoQmppI0XakS4YgOGkrDGc6y2D/2+
3v9ZMQw5/RbQ4RFsJ7L7tX1Z8H4A1BFVyf2xqg/cxle55+gdjummNRnUYfXhzzVV
amy9YWtvD0HjcYeqPFGZd+OYMxO+PNIFNklk68cehdlveHgokclCvgZSSqUZXND8
eVIVmbwYKGP0mybgVjVk18TuWHwNT/3iUc5rzb9UT/qha1B1tfuL7NZn6zM6+mgx
MtQoOkJC1CIehvVXptUCWbxGGBsQ7E9Os6HqIBk4TY6C3dq7Kre2CFLJcTDiVtpJ
UqOAL6/+gQWyrjwBM4xmWKIJ6jxVnZIBoReds3k4T6Z2QQ+zvsXxUZ2MfyPYEeKg
M5BtSV+yXui6TMZwYYLUEKGoiyMamrhBaZgnfYWvnJuWpws18YiM+5U6bAIBRVfI
3gAX7o3lQnVbpYlxKHdkQWe0tj4BzbuHT6jT2sATOoThIy81Y0ugLvK/BqlPDuJz
iNTwEDXTWeW0OTkIOwGFkaRT4ALFOf63nf/MOW6aX6uD+W6JVriXiqveqKgotJfH
bKWXPI+gKUCE/JToOfrHELUNsN5Z924Rf3Qzzul1LcJB/378/++rbAk0hePADhRx
ZHX7lOq8UPnxEmjtGCNhSxBjv7pXMAQX545DA/xWGnTQ6IS4Kzq1ZqoSLLvabmqt
wR7u8AmSEuId2oIKvng1Bs4PxdtvEO+4Vs6dq3/ay+mmkiBgNvBRI6I9iqpdBZt6
QtKLoEHr9CASVR2Jqse1ILWDv5FIBUIcbpjdJxSCPfWs/bmmTqw3/DccebJk/R7Z
5YhU8ksYDcv7gXvv+wRhL/INtCAj7A2VUVFToerhfhiO7G81dadlVUNw5QxqFSN2
nKXBuTmSEyx0PR1HilqRtF8I9z1uvieEL/UU6rPSkkW4q+LxsQljB2BAZc3GcfyA
hLuE4+NM7eJ3GRxfKEStPPs7li7WhYObGj1ctcjn5Yca07v1Y5Z1vA4cNyBnjGoL
WQaOkjd2F9XPAKopjzmMDq40CR5c6xgBW5QcE/2bYDVKu9IPQHesdejoRa+yAcht
9kSAWTFXc6hkBNUfLLEHmx3f4ldSrybeLlsBUgX2y/2Ea66wqxZpKBv1pSmSgp00
SUY+W0z1bFi9zrD7khtPzHHJIW63USJyyEhNgosPc3sr8rlU+0KJXqzOYHb1dxYH
tQg/3dP8+9j8NQUPS/yrU7TBzpuMmsG/jGYwhIADEKdzNyCmxzRlq3tB6rxpTX6O
WKgmx/xrcJJza0ltmzlpDO3kDrKGXxtv97bURacJSXW2r2Xa/biOAtTIUmH6nm+p
inv37DJr8HZoeMTwGSpL6LS9PtJqruNH1mZPffVWsnQN1r6hLzEj+PbXwWv1RPU2
uTfdWlnYYn5+V4OmzCgsEYPZuhAgd6CZ3DdG8gEWxImNu0LK6NMwZbSrJaEzY3hN
LrMSMur5Jo4LN1gWVRb5yH5lIbrRHlZaqa6JudTC6U9yz+cew3LCv5FxX+VlP4zx
kDyjaea+eZNMjrgWRT4UO4Qr3fCsIg04lHhWmA1kD81aDzJ31RxRGGxBp0FNoRTQ
BPtUojPhFc/J6VXjtCoarKMS3GF14P7MdzBJSJfK2M/+NL42yq2DOMahR/hgvMoo
0TA1T/B9ZBWsMC00qWccHoyCOMI81+Lj0suodS06uWTD5j3xqS4D2D5W7HC2x8wx
4+dU2FO5QWt101uoaRuqxomPAW98m1sroljYSaiEbuqmvQb4im4uJpRrxN8hYJk6
upwlQuVHNscM0m38u09uSnDpVT7PAVAysgUSCl4pzVAPyTZr4QjAgk0jbnCBhNHl
QZCAViRt1bWBoWb5GuNzFYXA7gx8nw//wLK3KcfGar6WPgIqJ+2EVQZYtgcXtW+C
RPROlwMdCOrqevTqZHq6G/OeBCqj6z3eZum3WcphXjlw84YeDHyAVyX7BwwprQuz
u62Jle0enYh4sPImRf8K76hSrYnyi0OernqQsOlax18DDyUm7YxEcGGefqvkQmpA
n9T81WEe2GhoPLTkqa5C4wdvKQU8nc0n90zwvudGaSHz4u4KGR9jeGCls4jc1aPR
gMm4il+rF86HtokolM0rt/n3DPvrFhe8ybyp9FsXpuTCmqops49Mn6Kwfu2ghWZU
xPZyVQKpsfyncZSz7m0yUIPJUMs08sEY1DfB5btvNv3EehMXjDhWKJHlSrMTpM3z
7vsw+Hr9PZlBILG2YTYrvwe82Do1fXaissXa3vRN+gDwCX15aIn/JFkUry4MDplv
LWbruBWesN6l4UiRtx8+Q+HTwWR7Ko1CpjI9xads/zeH+zkHtU3ICyB6rbR0ODHw
KVz5QinbR31J0i4BO8FtysB2zV8Uv8fzktj3fEXCEqIn2HG8WgPGgH9Lsxxd0TAh
eChhs7CfygwJ8zZQDAHrfqqeKO8Zt25cudAEqagZfSz0PYceCziSHS2el2ftGgFs
bdpX+zrytqFyR6aKO7M7BqtrtfjMZeuxHmeLDLPAefcbjjPRPKPuxa0nNFKUZbKl
tcZ71PwQVYb1bthTSpzVSYscxBw3jUE4iKS8OlQ03S0/0HIQdMX65H5H1Oz4FHuJ
StK207dJ/5FfMxLmhtdla1GL86zt8GcfzaFMrBkDUjCnjTnamwOBhI/tClPWBu63
br1SzI8cnPp4bJAcNh/qjeqUW3mRS8yIMTrn0UoRJ71mv/ATw64uxRIepE7AnM9j
RpqXGHDDRdapsn2lhm9MBhcT/QC91lJg+EXbhDspGiEn/iYgj5W+n5WSdICZ6MgS
y3D7skrkPv7j7AgoMNoWPzN970aOaj+RQimECKRClteLe3tMkpZudxsyvaJV7+Da
jRh2bkgtF3FcRUnBz5FraKZ7O9K8bHpkEo0K3BHjVuoPvlL5KblLbaimapbdHQRG
cS1Vc1lliusB+4u0c/X4/amG0VfdvwIxn1kAeFI8WPhebPOSQ3kCfLQoVg/jwppQ
CqTdRA76mNf085DT/yCzGGC+rgdJLMN+FhMfmZbvY7yYc6/h4XXhL8l5b4r93QXd
Fr2D3SNZ628CTEl7SuveXtrCwTbfdkyvRtCqNQ9/+zA2f3eXUQ6u4aFDSf79MuDj
2TCqLsqteIsiU6KheLkMO8DVjT//TK4yCNRXkUASrKS317d368z6nCFQ2vqPMB4I
gXDIVeXg2bY/Ob9uQSaMeUWM+3+Q+Z4/Y7nXhuzgmqXmiDWOb34OBigIQZ3kCZxI
GukYbsw8HQ8E0RPpAVj5B5GeHnLNbToSfotsX7GWWKrsyFIuRIkC09XC29fnEtyn
JHlNN0+STrsBzlIW65mLRg1zl9J1UxSNhtuSRh7Vcrb5lo2ir2ffHDNl1GnUHUjK
nbLaJcA2ZVOOH5m0pD86o3BhmCn317jEHizsBn6qGQfN3KCxX48o78+VbhDyQdoI
d1fxXcQFLvxrLz0gqfeL+h5zkwsppKtD5q+OBmvBI50cEsGA5t8Un+OMDeX6TvG1
8NuVphITzZ+o3hSEG+5hMNRAjR6H8OkyazbiBkUQM1gJuB/x2vLoCgG5DE/8ejvI
uMbM4vbZQ7IYE6AI1N6hh0kgIpbaduYarDhtMGnnuCAHtz1pJU5RWlPh8EbVvnU0
+XaVTPH4/tDJ7Gz6iIUKKLLb6aQI665Niq5Bp6ekmzxtVjKBaITAf4ZCtOup8p1X
uH/VnM2rkERdK6h6iiB731JuDCeJqQ+xVKRYD8FuEUEjjoowbXPvNR/cuqzMh7R5
DqmMy9aC/ZloL/x7+K87mZkVgNc4K52I+aFjRXWwoUF4ivSh/G0Xx9+zY8PMTQmC
jEbig5Lg3Dl+6tjzWTEO3UXyWdQYmSfPcbJlDGxChfpRf5D9LF+u4EJ6GVmSLZFF
3xtJgVOwf/ZFG7UEibtrSu9B9zKX5cw+SwBwD86DHIOT55SCnoo4Yw8mjtrRlB3+
O0XIGut0Bfj8f0mpxpRiy6UGLcryAUpGsV3yEOxMQbZteUpmXbTmIxrA2BElo4/R
0l8DiYFKyixq8eofPCMur2m+K9ItHfiMBYUyL2Isr5o2nl+wB3gjqkEfRqtCkC0S
2XreRCpNF/NPpiEI69xeQ+7SVNjS+oNuZD7eCW6UUSs2QpD2/YQmEvaHgyGWmcic
yDNIZ/PTBHiEQEEi7V9CmGWqByUUl0fEumB29dj5lSoefkVcChv643O9gYUgmuwz
AZSDfpfHgmeRma6kMaPLEWctw7plKiSGdm7LzDuhj4SELCoq2GouLUOWwYLtuDiM
PeF1LKXfL/SUUmXVFjcq/LhpomI3eu894Y6lBrPEJjHQdGZvr6Z10cP9yy/Nj36f
SNd5wvIH4ZB8v995zftx6nzgWOL9AWymgdrCaT03aD0MJHIV38Q7KEzND8XeLQBl
V+4NyD+Htm8q7pia8rTxgn+5RAIqSnFVIAPKl8WRuE6tJzd6Y+UT4n3kay1H8iCt
i8HPCluNv42xTszOkLX+t1pl5qjU0N0wSc8iY7xOLNg1wL23eFo3qE9biiJHr2AY
SI6rl0rkdIAXLItOBRC/1r4wHayTLaX9pM973Oi/UT6+qE29JTbeR+AuRJbptxy1
/DxJaapf4vPIO3vP3m2e0Bp38gi3gR2OGcJpP2NYB09iBpFoi+CO62xznap5FE5D
mielZuN/L4N5uTjw4ZL+FRCEhuWYFib/bP36M+EkJd9xLJ0N2Pk5JreJamVstP2U
Jlr3ykRjPcChn0r8GQCWQ10uz3Tz029PumU5+zwrup1sZt5dh8h13iTVryeY3Pz/
G1lT3tUIMR+DFfHaWYkRccVmslFMNT2WUM9V+nBHL+V7XVl9pM6e3NvpPgslmZvm
M7CFdi66ikRNkufIeoigajiBINma2saXomk2wicPtpUbxDZpd958ty3xFuve7dYT
7Cbdkk/pxpfJ+IlKY39607b5zO3Ni7ibS+gUR/hkSV3gZMaFNPSiTIRv1fQ1jQXF
T+OVp3GfNcnKJanklDYujPLwf2onwHfO6B/AF4L136n8jd38nUHNnd0zJKijFCZY
ciHYL0P4wcRy7H+4XmnGjTBv62Wf4qMbfTU1l7wF2Fci7QLxnJdejS93elRbouYi
u0yVVLQEOS7KE1cnx2E3EgF1Yi8+0twKhoD1k6cKG+BR1rlLDRtcjYtL3RARhIa0
2DGVHWKI01AWLMk4AVL6Z612boKmJD0r115xJHJycHCsKq9cHh3uQaghdC/V9aqO
mLN774vnYhrroGOZ0nOk/0y7TIPaSke4lVaMY5U67d+9qVyYD8twXDTrBAQUs80Z
oFY6gnFUcHFgThWHbtDKvMQ98RK4KejNfBRR3x5yhXAQlCwF8PaCeorlxtT3qlb7
mmlyERarCHIFy/qHOP68TuHIb0tFGyJok/qlv5hZXZc2eOJ5fh9lrxSN6ZnG94Ry
K2SKXngk6Hn1XR3kIyr4fyUt9p2wMaGI9uDjjbQaeGLFI1n5t0OM8Cebca6eMb3h
Q2p0h5elt7rWvXKsJp7nH6RHUkNdVuWggdgxYSYIUqyHrOVg/Re556HhOM1jgM2j
O6OlvxprVUEoaPzXzAhKv9tzG0GJN3nDCZQJTGZK0GBuJhVLzFK4evKYXSKOT37s
FqMEIWrb2knFewT1I/l5ostn1HM0t5ukmfPTWWG65M2RG6OSbjGZcmPRaaqkZUbv
X9l9S9rrYa7IwWGYrGAwRPsY5Pz/XZTmz6gMcEbo4F1x3Y4zlNusH/YuZh5VJGN3
B1iK/tz0REYWSQ0wtZxBgXFaLNlCHo5tlGBLO82T4so7jNTlzpuwyVX/vsDWr6eX
GdXozB4P2M94UX5D1S8B4dhonXOmiKT0eWmWMn8XhT6QRSVNFDL2C8ly9HX4BeWg
DuihR1aoxHvrhvC6lbJRe9fzjDuLlo+UpV1vfdfAlPt/bw3KC9W4xvSFbTRJdZEs
rxP8GHaimaEpbwJI0N+CL8YKA8a9Ytm6jY2MPo1HfxDaVD35hDF+dCZd88eX++sm
6q8TrFFIYMGipaVa7/XRj+vAzwVEZKQN7F4dIws0NiFA6+azbhtdo0qLfjiurjMO
QqhMKdZQmPIfzcqDuJhMHygFSjnhrqeJXsvWPv1b7R+cW+buYyzogmMV8fP9VyTP
yySS/qTYs2P/e/g0a2yrCfYt6rjZSVeKDN4ovHkLb93PpNAidxZB0aFL9fK8SPwj
nC6BV8s2Tp14hbBtU1TpLLn3t49laSFodTnrqGUp7ohwgV9u+ovDz0klopY/Nfm3
D/+mrC0G8PntpRMaPsmVripa2bizRlxq4Sf5W4PHckC7/jvMUoKiGCFQo8/4Stqj
MbhJ5HWAx0BKt/ADxCXIRzMJK40wJp2yt2+R4D03jzCmpka8cAbEieBgXHiJQrZC
X7KEFtJEtFbv+zkRRucA68vtGiDgouVQhDmcvU1ubKZLHMdTUYqjalVd72DnMUqe
Qp4TZRT2oYKilNhn+Mb7CpWq8MZt8rTkgQADu+RQe8nVqLGRbvccQhzgKIZaUXBU
DTEHAnmpbmtgjOZCeVJSJy4rRXeJb9lb2bOju+AwCsKX22BBhLkoe7zTR40f0Adm
BCttijPJhfsWNZ33y0i8g6Rq4M1WvRkkSawR8f+Cfg9liemFdg3jqa71od0ZErwt
6Gj1s9/VmrKWHQ4gyFbQ+F2+n/To/fNv/R4fmyk9LMRNs2hLe+m+xOTiG+kBan2D
Sk9v2+kZmI74Kw+XGDr9fDwDvx/nMezKqRjwdv5r/7pYiOFAiAH1/wHItUEiwtsQ
uXJmowIsVMaz5qWIG1KkNrK0C8cZYZB82vqz9+4J/hBWD08jrWUz7GqtZ5HHiCRV
vdjHDB7VHPcRxd9t4zpTadscRqHVtGjKRTG07rpuJp2BIc6bTbAq9d+LBj2h3rlc
cKgFzstQ7ingV110p0nKW4q/u89z9NajFlDZuhBSTx9zCI3nviJt0tnknHHmW27w
B1Z1+5QXQ77nNDLLqafOYjGIqe6gUeeMkajiZR5ghrdzyhAOLrYn9IOmLudLdcWd
EaJIPlYP/e+6Xp6ycj2O84qz0qAQhyUhGxiFkmukJiDTS3FbO5fWCyEeG9mThTrT
Pd0bkG2D5GhpoUBus/jz5nm5U8qUKVgmAgG+1QGtaD26WGh37hRyW/q+L8+2FRgB
31hhCb8W9T2GexLEN+anXpZYPtvl2emLE22R3pGdJPD0lI0LEAiA3HbhL4CQPJ1o
5bm4ijMeA1Dz1oHeClgW9Ztkcs0aPNUHwrvT3uhnAzUojzqaTYrlBtfg9T2Xp7II
2/ssQUaYvX6Hfvuv9heIC4ZaoZcKqlYvrBJYvhpNR00xHZ1O7yjcwibZD6LPQ/5B
hVnA2sFvAx+IjFaFHEixL6XohZY7J3WB0HmTaVzK5pnZtS+Uhf52xebNAL4QWb0e
NxS3CdH13FzWLc69u3pi9hLqGfjuAGAR+/ocHASfxY6SNAZ4CTT2IPxxiW9OQaPF
+gjk/DoaUKidvORiNpbvb5heUmVgA1k/gHrfjwVam0VxGpFXXRFdqIaTIkoHwM3L
ZETWliq7ZQxiPUt/VyTgPB7s8MZR5JL+fZ3GtZgBHKf8gIKi5e/DJkA1ApkRwRA/
wQgtVDqdoF7hjmfnff5afX8tlPpkeLg05Be/c7ySNvgIt77NoMoyNq/wpcNGd6Oi
OdK+Foa0NuEV/1sy3KrIOgLg28FCZxp3eCeHldwdXWvyKEDKpjgtJkS+0lJs/Zs+
WmhtQpYKc/Vqg4C6oUdF68uk8kjYEZDpvTXkGbZR4MKrp9GVOXvLS6E/G2PMQ4Cb
ZDvXjzArCPEM41EoqLBDWyJayOl88tGBHTtDxiaey8QXbA7xhS2MFdpWCCZMuyGy
ZOz+DwPB1F+iZz1Ifxt1OVN0onqc0XE2LRGHdHGoNGAMdKiHGLJYwnkGtwQN1yGN
VVb5GDCrQBwDlvbE2TBdvuwPX2LKHwUNj9cX87VQ6CQlG8dRnh3D0rHGgQunMt5e
u/B6BCrrIVq/K/MSeTCQlU1Vo++E9P2UrEBLvimR38AHWvxwdj27zYiifeK9kULC
Gc8C9kTZPidYRCvCWTmtTXMP+0YH0EsPC3LAZP2TdAmSVc4HVnlxrCZTjkGcOu7c
3tm6V+4tHvdpztODw7SilO4Y5Y0zAaH8bGSFeYGjQWhzGfv4bbrUIVYJSm/S4bt2
W/V01E5XczwWDLsnuV2GKn3DUpPDha3/LPkL0vNvoWwrTsUMsIXE7IbCndwEtESl
ZItqbsQitdyEoRs0YM1hLig0gU1CbX1y6pds+2dWKBMoQIGA++6BeXexPi/i4LjD
HQJnapDaR9irDZ+XpHSlkdum0tytkD8te3DLTP03vwRlh0fK9bh6QBihce04+/WN
6HjTRW98ehPCPl1l/RXDnfYsFwTK4EyT7s+hwGWquK5vkh/N3jJefQJ9UMh89rJP
7VS7uC4jBx2BErTW8KsOB1gL73qMvFk7YbQSgMNtolBw+y14q9iT2N5I8lnDJPuq
cUEuh7Lh87NcqAgDQB9Ai05VLVXLp/rZp0fIWbT9bkp1tSjIHlji14w4O/F4CASU
5ThSbHeXPll6eoctk/o2gy8VlddEmahAal2M0WRSBGgIU85OoaWrDcFUkLJUdLc6
S9y5fqpfruIBCrVIAzU294ARthrlO/mWEfVxlmQwzwU1Nrj9YyXrlZ8eTdFhKNFX
oRPHglLwAXqWClgUExF6nbn6YmcPg6scklF8NnI8MzVkw56otxYL3Mm7aPMDN3UC
KUTVfB+Sn0E1Jj93C1x85E4KMLUrAZgSNnh5vriRPAwCIbJtfAWRJhoBT6AfZksU
1cpR3ANK5vTf2KwgsgvWDz6WFuStNe4OcNlw4NTX9+eVMcXIWt0/sWifsYV1O80s
0/h8ZBigyIxG34hIeQt6PoT8PnFCYMz3LgQFzBBfJgmEQrnCITDEnnoNxdZKkBJA
rgsp9pJV3xa3lRe9upPoVlGAGmiiM6jcotr1naQZazNI6aPVxyiP6L/5DhguBuyJ
Ipk/YkUXMCcEZZP6s8URldPOKf+ZN3AWcNh+D/Zg1LdRWTJewP4VMA82nZq7vppr
N5eWaxQveOt4vQHHqGxsY/qZSHTOinq7TPsrdYhLvd6PXsV1fK3C79ZeO4HkxeyN
YaN41JC4snoAptkVuljVyWBuOlKHKz4hj2pq+xz5dwVW6A4X/eX4q4Cvi8JBNAQR
pMS0nRe/p27zge4L54EEXYWx9HLFr68PMR3Y0xMAOeYRy+PVBhrHah/ghR94fVX3
iZvXCuaQw9r6KtEyXKUAdCBy2UgKf9lE0Sdv/GIRRQ2O+ojCQctf4J8xkw2GbJbE
rPfMvuP8nyF/MDKB6dDOOv6KrVw1gnUPkpC1Dv0jWS5ANTaeXFmu9186adgnUS9m
x0YGiqBzt0ifZby9FsMMKI+6If1EvI4BTePOZfOT8GFPLFGBqydtrNntTO49kz7X
Azu5pBD+r0aJi31ondOOq6YXshrJWkZ0PSuSBLDPsHwV/EBg3/KgPo2OPNGHMb5U
bXh59eDRQpLTyxAIFvzIbZmNRHSLg1uHynVI7CRPPcLWAIF5ST7sTCceq6uhvuBK
16Rdtc1Bu7xfR11m+SD4qzVaQmDM9Xv13rZkNFXqsdMfNISf5FRYbFtA1TNIL0Yh
x57oyrua7mEfq/iSXIjd89ZRMMCMAqBN5rEX1S6K7kosanmy6gvyCacrXf6YqIPc
wtJrMkpnFJWNlML1Ew6xmsNSg1RMtT7qJ42bHReraDgeU+gZWGBmhoLLY+RA02Nt
hPzOgbko6kWcsEe9jbdXkeqsOnUk2/c5QYWDJO9ux9XUG2FGAYe7X8NY8lFlJGRH
kHONKJCksF6rGUYd1Mw2HBUDc0vHk9LOIksnPYnxggf3k3m+E30bb72iJ46SJnfP
F/1qspnMqCHpr+1aeW0N09UQakJBQEk58niE9MGexWVC9rDq4wV9N3Gf2Rp5z0ES
1t0SWQRf+OLP4/jjs7fObk7PSIy4ItZvV6KPuOTMlBkRV/ehKU1cnaJx++3/nZ78
SsRHywr2WzsvEXk1yHZ8VNdCjPDldzyCBQuyfEbA5mXiHw2n7DcGyxBY+FED6cD4
v6UjrTkmCB7h/0s/7isfmAuiWOaq9IjeFVwLnYAJp0KjwlFpCLfZUBqet20iMaMV
oxv6Xvrj4bPTmUE6Ch1FKaO2ZqnWE0Veomvak4M1u9zT1LcV5Buoz9tZ4jYci33k
d2QOEeqdKLBDZ7sKU04IrPP6EEwiX5iBTQpwWGbsDQIiBmXhlHHcoMLi9gwnN4hV
JB2nz0gWEYhnun1cNZVg0ir1FjTqDlHEXDXv5ik24p/AIIJ4m2Nj+ygraDkjAGK4
XfVmVdBwcHTUnerebWTPuwOlPjSu1fy4pXU2aQXGdaIRXrEoZaDdLg/cr62LaxN2
8RDF39C39ezY4G7ob7SQcUG8oWsXA/x5ZZg/tATclr1M+fCDELOf8RX93F9LIvBI
gOWGNHhfI2B0h13E1pUij3Ss4+wQ8LTklFjXh3UoTq8rCgNSAoqky0m687mrm5PH
JxV1WxxE1uXKw/00ymdk13iUW2RuDBgrClaXtd36wmlx0BVsENwB0UFVJFLCizGM
nIShpHEJrnVMahXC1/MuVSeXfwx2tnmR6Sxiw8xIildq9UJcXWmsv8ushzYYMWom
i9tqRL9pSsO6Y3wJFWttcmFmYPF671jrhdVEKqMDFgIKcaNnTIBlXs7hWDq5gtFH
4dI2/hM78gcaLYYvH84PPIG+q0qKvDIIpymrwcMaxuXquyfAX23wWWkUV5ssD0Xd
vofD8BDfFjIu3c0NNfgP80261Mvux0Eyif3YNCia0BQ7Qo1FaF9sVjlCzPA8MzUm
snVGVwMqGT7qQ0AdyFTpx8IRc7pHqYnnWFUMmmlBdhp7ffdBu2hD7qNNLRuomZ8c
97HOo064GdFkrok7jEXxqcqEDVwGinjjyEZaiLg2D66hMuKsmgh3RDfXhD8pgNhv
UT4pO0DWqRfSomn2lqO3mfzlDj8VnAMPr6eccsI+zAtdZj5nWLgGECBr5jBfV7tG
53cY5czNlPaGEjxim9jy9THEaF4yBem7lMtWA7rH6P1VAiagFqxKps5fMkAYMmKe
rbrqlLBlx6f99npvd0UDieZ55WxZaK1s13K+B93OwDHhgiJOhCs306nfRMLLjvnm
cXfxta3AWAU51cUCfvHfiseInCfdHipuKg9ofCkwTbp69my+kQpdEKOGG7fGODsI
Sd82fgiTU1JOxjMawIeKN0tYeNt8UZSI4JWiB3LZsVLv0VJ3hG6ZBaRkOAHtpVU4
7HCMleOphqLTyrWOf9tkSXs5IeApL770eMuWV5VF0c0hFuYkzpT6xMV9mIxRMAiS
2GvlEu7Achsh328WPUNRzanq+XvPrjt54oznLhqM61npZMkCdXW1xiVMC/1tuN3b
pIZbnI/pECrKUaGPM0JOQzR+cpS/ZGThF2N8BxWl4oqNjS1nyRpF6NkLNmU0gJm0
7jlHzWR66RH+FVNAf7BtdVNWfxEWickLH4Pl/CpYV9yR7Sx6hKdsFwOC11QbOnjh
vFktINwJLVQB/vcx6dBDNYuNUHuLWKSlyEOlcralNdnBcmaJ/zt2IgxHuDO07Qst
lcmSvrT5N+CoN5/88qeb0VVPH4N/Q2fOlu22zmwlRqXuRxvtRibZqwBSAfTMlQWA
mj0aKlr7U3PL+vsjMehtHdxv06sFJL/X5UYzDG1+Ta6IAESrdLNgIlqWbhUCMKjF
KG+XzQfAdCHV//5r1rfXaxlBo6cmRj3LHBCYSu8s0nccb0Kqui31u1oNtbI0cS4h
e5fb8EUljjAzWBWHTRj5yEOsNqYFUse8ISSPAZmYKG1ydRkGl3LfVuMAZPYJbwed
dy5rXfX9DZpRUTNcEwTVYYnAYrjf6qNIt0MQIFWsR1fB2heuF2A8gWkPg7zHR/zA
MkugV81zYT2EGOGjak2nzy1YjM/105CcVYE49upGr9BkyUIdeWWXciDuywa1T4hr
aopFvdiZORZe88aCwQLmLrS2s7/e3ysX8z78CYX4F1OmD3FCoIzWQD7svVa5oSP4
JVf/rxR/ZBVec44NbXKTsMDI3Np4LRiBtX45g9NAmzka01HxSZLStCdvSGxmKu95
d37Ky/nZQAAnroooi3CZcEjfiObJf0XENcmGALzg1E/eLCeyhTG66K2Se7gDc7Tl
6CDRrhTQajeNovdmskD3fkc+QTdWMQ0KoKjdbMLQKOjWC8wm7HGoHtE+aGgcdgCB
NDIjgUt4n3CiVEkix9qKZr+bCu1hD3ValAHDjnchIKGNy4S2Qz8mdMZcLki+kira
rMKHXvxqBbsYJTwdukHuxuD4rgwVer16UuPmwIv7WzZvSC7gRMTVvY8PQzPBZS6q
t0b4o2eq1xQAdsD1LwD77uBI6yPplfeVh8NmE3x0kNPI6HVt3tjP9swwxhqq4G89
5DmMKifNiAhFZKckep4bVg0HkKUPO3vM6y9dnZVAPbv/CpuHSi2EUxP97dqa0qkk
eIGobl+NNgY9GC3bejt9VkEb/wfdTwspGLOFcwHSlJSHlhySsvCOpsJ+POu9fIfM
h7WiXZ6k2W11tKmfnitK6496mmdbHegBYcumcrzzyi3QcU+9VF5GSu1zpP/zjBeW
3dvBtqTMLWzamjJ4csqASNQfNCnAFOsvWtGyCQtkRtUV0Sqr7AMKmMnBr8Y7NWic
6KmDeWsN+aQWGASgBbRO7gGYLAbTl0UgPq4TCD2EZT/eBZ15pNZQeYqoJ1AWLLrJ
lMIHdJwU1xHB51kO7h0YUTui8u+rE0FodR5sNlholv1oP1flBhKly8GqP4wVit/Z
Zz7guDHZ+vQ47qjHTVoJGuCcRmmkqDA6KVKMLh9K8/GUolfK2CWw7VOHDVuYTLHl
nh1fUYjEM7cexquZfwskE9ZTBMWa9AsvCMr3KrQ8OGAkcD/upQV4z4udYFuJVd1f
EgpdfY6PCV3+fJrf3qYl8dve3ddwmG+dfIl3tDI/f5n0Uy75goym45MYrSAXpCpS
em+3p3zoAxJltAVoqULU9vtZ8xjuEqiUZ719HGwRzxgQyPLHXau1zH45HQ3MFrC9
ulRstuiTnUOgLYyb6yeMMFyh79FRur4pPL6Os6CxpJUwnpjpphfZsOc5YrmWnUnU
I5f9RvX/VhWQu6/ETJCWJeCxTFrTLtRUJr72zsp2Nqa3hFjph9eeLjDybIzxP2PU
Z5JJ0isw+HMVC6ZSXUJBnn+2Agu5q0aeYi1wWW66tj2G0ipPDF6ni7L3TW5Y6xad
DfEzmf8Zi6WglYDt+B+/QMKf3ECRA8ttv0U42SvdumCacrO9o09wtWCZFVcy9Ju/
K1xAVUpCBT5busuQCEtt1vb5tlulfZikDGnaWTppgps8tL1B7KgseYd2VoQFyN1M
4w6D5shewfag2kqRCBifD6eRXsLMr/glh4Cb2WbqDptzTUwYJq/pGnVgaGWhTq1C
H8aBk/fSVlDIA0HD0LzjAvldKaXoM1MXzD1GwcqN5IysEeSaShDQXMUp0aPbaXYa
jiA70rjFzogIERQny8ry4OP8ffWWr4DXDXq+qyDfgSIT5sEU098NkvGt4xI+qo0K
wplow4bi9+Gzjce0x/RN9DZECe9UZt404muWtAeYRslSXCGxnKSB0txQEqKXUR9R
hfJeKTnSwg3H6SwM0ooN7wawJ29Ng1McPnf+ifXxEL74QVSL+S3GJbs6BQLCrQtm
1MDNWyg9XNy4O70g7iSZZEH5rpb6fE1XrTxUrdVenqumTfRCU1y6NbP9x/crcl9P
IOJ1A0tkuO0s7M8KdQk4skkR3kZlTlgKtgwooe4Xe7uyDY8ubdsegEh5pTnipvOT
5QFfHqj43E/wyFpovf1txrbNnXPERWIkNW8W/k2k+b7Yi7qqKMjwoj0OkvjWQJ3f
wNNkMG3X4CsGwYLA93Cmf/RNmIEfXs4kEvfxjJwNrEzjEa0DMPnymou36anygaYI
JVW1u2VnNh/n3WbJBWK695nQeaNihcLylEm7KgC6LFInXCspu5wznupWRUsTNG1w
fhSjLVVnC7dMXtNdfCHomDcwsPLhQiFRx1s5R42v2qkfudT+XJU29riWnshWzPNv
0xYGvhsYAjfr4kr+7f/ovxrNmGKdXGMiZIbzKPk50GCVLPXpjRwd/XrR8A06lY+Y
Xqxt8FmTnY5THXR9FyUoVyhhGnUb4ud+2tlp46Vhbq56jxnHkxBtaiZ1khFnjP+3
ZIc7lNJEtyPnW7PzzYbjxAgsuKKKRLQMBiVVKPiR6r+tU4axBeFGBiPDoXbolFuW
YztE375OuhHA+UQ7juBpOPv78cHGPLk4McoVGDf0KFkLE7KMUKCNTsPfO0nNHmMf
q+51UJn9Q5l2DKMH1PTkqk5nPUM935mANlE6cTQFv1Wj+sN7vWpEhp8sVpcgx9Li
/QTrJVmRsajHNk/IZvMD1WCbwziwqxBQst8sBa+xhvdYfabeJOwguOYNVdJh9vf6
O9eS+jLB91JVY10PgcCC9qTvlmND7+j2VM/wCoS7O3e7f7ykxq6J6Ub8cdq5v4ws
n9/gfY1S2wDy4q3l6cN8ALPtDivD5I/pXyVaeu1fSLNXWKCWJH3/nFlKsC4HEgP7
ylfJXeSXDciIS6e2B83tIBjFcn3/Bkr+cIgv5tu+fmEZvfYx2QXQemu/7VbhjGS3
FnXfQjgJfu01V66eQ/uiPaynkdrna6gutrHRKRQhiOK5lkbY2ctCghdblqP8vAoH
nGmamwzx4zxcqdg9nTDXrVhPbNQ9FlR2LsaFmpcDYKo79HMm8QDfIUn85Pdi+GEd
yWFaV0/HSdypYT6nIYvYESUouSxPNt68T9omgvbW4U5a/IGf5/2F7SdtTXObWoqn
keHMyraw9XLWBOqiH+JuQISo5vecA7J19BG85DWMsSlVUPGmtacgQAi/0dUvUyD+
ny8aHNq43S5ClU/F1oVAcA9e+pZtxSstFNJuEBP5OkfblyqiBx5bHX9h1xsMy9Pp
kMShq1sHm10cVAs6hARAQgKCkl0Bm8kwvRLLXjyC8GN/e9yui2fhixGOMognGGrH
a65hMxnAxTxME8Ih8UI1v46MSjGQbwXK9DeM28ND01qUuEmQ7vvC9A4quIe+PHTn
rcQZgMM2gdP+cFUZoXRNJE1+4f/vxD402DDnoSR+ogLnD5Bfl73i+1m2Mpj86ZTH
i67pHpl9M+E9hgSQkHeeQ32/ye2Q3ZJLUxEce+9yxUtzEkg0rI0Lkbt2ZUmOPLLF
VVRvTHCQaYc+QAUUAuAuo/JnDeYpep69N9Y8FiXq4Ds1dbzWBD1/vPgJ728d/54E
hvjWdaxphZotQVQnVaZEqF4C/6YmZ8bOnmRGM17PXKzd+N1WHbpICd30AS/B/ylk
FcXJC6s1V9peuJcdHxLo1zq6BdSFhk1c0kGCFt9A9UOV0CHn7xIARRq7mVgqYNsR
4GKV0a7GnPH2LmOO+MKP8ORlAH3qZ20P8AQXqUePL/9STO2PNAcYiMLC13qG893M
zeg9q+4xSD3+IOP6t00R6suinOWa23zDrBriHjZXVag99byTO7tXjXwrw/v5t3Ju
no+0SdXSX0l8SCzNzMLRPqMIm6uCbwNzt7kyRCn9o/KVZGbjs3Jy2A32+sQYLAn1
NZghEHCbWbd1+hAICLPi6BXPjhQ0c8ho1eP/2yRrhxke2PNfxsCHm/IY3hwifZCd
ZzzePN+PqnHCvZPQ7bvH22JhSz/+FAlk55cvfFyqGrC79w7+EmJWn+LYTm1jrs6D
QaBGjexJYbQZrPBtOseV3VeX5n4/ZkHIGP+3Hdjsfhi2xPYTnwJD8lPYmfpS9NM+
AoJueScZZn+ZYOKFe8Qsw/DImuLr8dqLd2EqKTFyBy0J5cW3/RGE8akx/TYex0TN
riOvr5fH2ih5ZkOEbIlURK3YrtPBv9J5j8ohouiiuUUbz3hKYcZa+r8LNDY+T20H
ZcHa38JJKQuthkaoMtJBH6rpibFxmSE5jvQnTm20LQf6f8w0aaWV4gKk4hTBiDhq
+mOeumQxoiH1/60Jjb1jWCJbRvpfnM9XTNOKS435WaVJFlm1mlqDrCCUHZNo+MqU
PEY74OStiIUjqoiWOPGsZUCwWetpKj8m0N1MbpnHaHD/N2IltObOF9kP54/sLdS9
BR3Kg6EEat86SwaAbwM/5UIEKiHPQdv0c1XYlUyfOM3m8XJXJgRnIJKyDJxFJD21
wEOBaDRuxJABm/n2NUCMj6cO/xrW8o/m0Ii+Qtakwy2lzQGm1FdDATHS20E9HVxo
h6WhBLG0SN2a2ws2kyf4CXQZkjaLamTJBxjNBv8ymxwiD12t1sjyKWOnEtHR9vmb
6uD2cz7n1gzHrf14LXGy5EUco9synKYQqJIq51FVrqg/NeaJhoL/dDMSpWkgYgMJ
HKzIR5ZtoHnIzTvqB0JrKUM3SLs7mWwI4XCf9y1nK5ma64+SbEEp4m6pLj1vsV4/
ASIaa6d3d+Rw8UgU/y8XhmAIRZULnOm6NcnIybWg2prJceO4zJ7+YLPfRpsWZhIW
vZE2a+tP0p+Hi0ColI6PKkRAquPYbJhEkXTUV1dFH5diaLoUj0sCYw421lbb15LZ
No2HQ+vJMAHRExE+LL+6lZ7FdVdy0GGF97b6d2THGd/G9vcE22Q2yQED4xKYyWBt
Hp/KV8ZH/mrIMwfxIRsgVUTb7T/q3t61rantsOb2R7cp4wMpmvUydPMqHs55vn34
Euy8rKfkLC6EN9G6EniTeBLGyq4UX5cxuesG9tBfbCeHga/jjGFpXM1mxwI1gG32
qvw+kOG2neBFkmGxhUkdkXPMQIh9mPGanHcx1Lg7JjVKnJisAXMjOF810J3ifUOv
3fScV2YMp7a4x84FI/M3GFWy0tPI1SeBF9avtWx6XlCKs/xrPe3MKuZ3Z4WtBgI1
0PRfwTbNdy8guLvPCAvaxS6vGWeEupE08pTbYxscZ2L6NcCFJYF+c5Kw50E+YUNN
Si5se+qCEeQMy9qRRqvAV4BPoBTytMx1319hHd4JGycwTgdGLeGQBN40hIykDQ4E
7G/F7YoxlDSeZlz+qKmxgLOIAnOFzf47RhRxLSEBIG53DuBv8kXCUy9OGU7Q8IY1
LddOVOb1ry27DD49Q4KR9/tmkOdMtpqyncTBthUzkxjbXx+7S6c6Dhk7icF1qu3g
ez7Jj2BQZ/cdDngeYNdher48cGguObp5AszlUzvZGDWgED4JVIyKdajUytJsszGj
HLXC32Lsjj0xYD2i8UYKLhHu5kW74f6lm7oM+xYtVvQpE3jxFE8HpezwuAwId6zA
3ReM3Wo0rsWTuJwawiqBLlAm3zurpx2XdC/vZywWy21va3+8Rnxuq75tGXHtbfb3
++Oh2pm9kp2nMBB91IiMNMkkL4/YnvZQFohnSmlplhzTzD80mjCeaLltYhSkqYpt
2FW6HHF+zX4sEDyWA0ILMte/RbZTByEt5EKPd02QC4hQBIRAjDGZ3JfslfndPbNr
QKV0e4Ruev/Dot/rT78ZWhaY1KxB4bHuW7dBqaHn0/Pf4AAAazrUuWJO1HlTAU/P
Bk7kazEvliGN3NAnp5yIkMsav3ezYcG1dNkxt4YYrKzVnnsF1O6yZs7zBB3rWIwG
4/kpOG7ciTkXiIZ5NV4HXQFPtY7xZrdZPssmqUYEJLC8B+23oMrKil722o8Miqw7
b13EQ3aP9lb7xQ53UvtC5ml2yOtkp/faDKoJfBTADT72cZsOBwMc8xwNw2QWKlrm
uIhLVVbBtN4gJqve1Q85I2We+DXMPdP8nlEW/aeQ1Z7jc1JeI2mFAvRI2YTnkF4+
AH2wP54m+A88WtFA+F40FSNtTOXNannX8Sr4NJVwtSP0FQ/g4aTLElogjRUXwe9b
IP9uhw9qK09jfYCZ4CzSi3B3yY+qMkJkPPpwzc10CYsmma9kt2VhSGGB50xw83+B
n4qFi5SQBJCM2RcW18szWebtaqOB2FJDkzJmDJi58zGLaVtHzmhT4dvF1pUdHNZ+
TDZjMbpEaXK4Q80bCkn81U2g2QI74UTippsI8EnhNgqFTYQVc79SwKIQTs++QHz2
b96GFTZWtCpv6bVQG9d5OmOaQtE9+k4VhBGcTRrsuDtesx51F4T4HhvyjbvWjyoE
lkfUdv61GvZgqEZNIDXLg1umbhsau9jwtNNg3kIfc9oaB4VM1+Gt+KdV0TgK4fPb
LLHJJrehNkvrykAZ24n+snvspwVDH+b+fTl8rkiiv18thRkOnLIf/adw5Tcer742
u9qQ8unFAqQiqOcvU880zV6PmFExNYRVQa0EI2SsfVvPBCSc4TgVEIuhooapIM9W
o1Efgrc5koCdofl0UxIqNBx9YGjHlB3TzqDGcyFQru8tmuYWzoZosb3I5g3MBvTq
jUOBnB/P7L8aKIoiiF8ilH31G30Ct50r/ORUi1r1pef2jk4sjEPb630Cfn5GhRqO
m2PTkE0o4NJQbKmtG5NF7Pr1vHetJMIH3usOIR45zdg/GqCZtwyg1Pp8YRgHNvEi
246/wlBM7s0McSj4hTUujqekyK60lf0Q4ssNnCA52NuVNmvu7wOxxtqNusujWebD
UMkKqrhG81tsQ/AgzBEe7x6mBuDR0EVUVmCIKO3KF1U3IreGbVsbj3SmuLuIKsGj
UU9h041z+LLkPCvNDnhQAlg9UrRq2WA3aeY1tRfb8K6TI+aHyROCLAiSShFQFyLP
cGMyXu+vfF5I82tfXNgJUOv41n/EpbIdNdKSiIORoOryNz0LjwPNo3H1nJ43Jacm
LfzctsUxTWNBTUfp9q435C8O1d5fMI4fiNLL1USM+rjXfhkUKZ9+71+stBfHOtIm
UB1SmV022tflqDmNk7URI4GPGVoSy8CI1s4mArxnwnpjT85HtcQb8RgfbGbK12jF
YwEaJgxzIfCCqbJVYilFBAjWEeFBwWfegLPE1RAjqjHAIVym7eLS8Z+fzB96caY4
3l2sHYVNM2P/b9wf3Id7U76U90gQkjO9ZwRiHot/Xl8RR2MqjlZFsi/I/89N+V1s
47R6sc4sl7IdBFwhk6LFB+LqSdjGGus8ivN3ydQbfYJs91+lyxFkDJIvlwXOKBMh
1YC5WVNAuBGNlgx/DvZ3Efv0KGw2P6hAg8SDytW9E1SX6sqzBRzPNbH7uqVwXRv5
TAVV90HHdqgpuNWaIPHgo/znbZD2xOjVJZ9SqAZb/3lne09WZiKXBMm30C7RHyih
sCMgEFarZTTvZ4WOnmip/b/csnJo7iWlR6YLAHuMDfWd4kFejQaGW+dhHkpeyqHB
cT/Y6zKmLKGo5vuWXOC/3/qFkecFvoOfQqcu/KF/abX4OMnURyVi8AAY99MDcWCQ
ak8fGzJtkXLf/bxUPkelMejMqgRT30VBoRDkG0OOqL4OTnbcqflI3Mees/73QCzx
ncrwx/pSavx5MqcZ4ClGmY4hz1cG7nPn8+XSvJzN/Kz0OrKvf/ETXTM3Fne+AnJG
k3YzNGhX5zQlkLpZvhr8OaNP/0A/r8gm2bFvEVwbW+kmGBoOYe3QJg275TY85Hns
CG15mwJ2cIoK5ji33AFtK1zTcaLmsLsFTh5rV1tUUmLREGSWkQJrU4+Bk6M7fRGi
wYru0IJie6pTJt1xo21un/RvsJfEC5p4APqKzGFel4bFOGMZ2S+XowgGgrzFCIcq
AoC13wITWB+pHhgUtYYWo9x6kPZWtWdf3BlmPrQrsxWxcpwwbg8VUUkwHp0sZ5FO
vJtRqspGFHqS46XpYPrXKL7LAza2m68O6I/J5Kr/g8VOgq5JLbGJpm6wwbMCcQa7
iGTTJQ6iEHia6zcnEz7gcqr4BCF5qvj39BDPOZKqhFTU1wpCqaXL+35RsUMnHCBl
T8UbJ5S9kpdMdf7OaFv8U3GEXHa498pnFvlTL9h6CiFCsufJsrDZDxqEs1r6HRM1
yjX0BPpsNvHe5g2LuPw34+hYGI+KkTWIC+DMt2opEGc16ZbkCulUdQ39O0BpL8+e
iKzwQ/CVFgmZ9JI7HVo1fKEveLU4y8CMtCPwUQllBG+yusWVXhTrky4QHlQl3Xk+
DVKUjenNPBtW19VEOKAWyTl1KFAOztNHEwOjU8VSmHcbqzyXv/HMlHQ5ZWwPAXcB
59D5b8nhUBHK2c3IgujHWIlKrmLKPj3NB7meNNIjgagVSXbJLkCO5aL9wspdVySI
etvETzdUnfZ+KUPznz2eIs3OrSKakFdXKgmrI0bp5ZxseGeMzNRYPdCoULDmTXBo
NcHNqkdZ2ykL7Bt8lxR5Z1ipyv7JhoTxJ09b3NFpg3tBrmbTPYHD20hWGyLW/Hsa
tstoj0G/sOHKXRrQsqmaf0cVlhAYh+rn2IPO6LgHKxcVTJnp6vKyy6WVGOXUBGd1
p6XFedi5XQrBZsU2WGE07pw2FpKa78c6v8kUB475wKeNz/odAZ9KusxEKgu/AZzt
iYMJlvgkKDPUufLaJgZ/8O8hdu7UwsIK0VVKzPIIUKlpHPD2C/vwWsmVLZgYEhzr
xU4H6WoLEmAyOvjFrlBT+yXXdXe5V7hnDl+nuV+ujZ++n4PiN7NN7uwACyEpRkA6
Wr90Qf/7C8qJ2tHZlOvaA4qLrZ9JVXokNL3+U7HqeFyNCgutPW1H45GYnzk6fxdF
nD8BRVSNZPwVzi+HPNjBHMH/wkDwGICXWI4XKfnuvd//tQQRxOESCHsaqSa5dau9
Tc8vSItXl0kdv3nIdAc3U/eAQcn5aztFAnMgNjD/YZJ0JB/XZuQWiiEuaYIk4rzQ
7xjnhteBIHrzD3RCtq9UkydhLFwIMsVFNnETFjB8wxyDbRyQJFsuCdf/XWaoMdUy
Q/go7Rkc346uZZUxX1SEJ2HWWFuUCUsAda9rlT3BUtdQRnc/a0k0Mt38rkrWVeeR
u0I4qG8XHl3zzvYNB1mBecsRqsajI7SJiu/dQgbM1STMaTnWAVHDUMpj7BUEoVIN
k6S9Iu+bdXa19SWbYO6vrKfbLIBOZCeFwvtvhz+yYaPW6FcpjMtu8TvOPbSV/YJ4
Y6SWZY4aP++GhOzE5ih8eyg1rdYGMh56NruSaN0K8pgOTJN31y+ovLkNl7apYnRa
+3HQpXKIWX3+0U7ii9VujHCsSjjhSYkba6SNriu6i6xm4fS/18Fk6qrz+0ikbjBt
qzTOQOF+iP1b0vBWdalqLMruiBekGwGCni6z4tJEZXkXjQ/SYeyu0tEBGy0E97br
14sALysR5xvExSAVAwE/XpYE0B1c2AZJa07cU7yEPLeXYa3WcvWyBtDipWKPEaXC
L4XJeW9weCqLt3JYygt9rW4C2gyM507Xu8OLxU1uXLeQV9jRwvShcOWwV1ZsG9YE
xPR2ecXrDk3CEp/dwsxCU9PrNq9/np4u3fz+haDIweKSt84Yo5qyEy8hsTi2sIRc
s2xEQZLTmCiI9dYi4z1knODhkjpFjIiicgRQ9OaNEX8jJ/Q6LSaBUBxzttBxmcOK
dQraL1te6j4zsCfXPL8FLD/Ap6YReYaR039GUvjxZ2m+0hIWokuqmUvJTPjgpIlA
Ah/5ccKWT1rnCbaDILd95ztqWapA0IdouDwBJtYZHTziwEyGSZ4JnFJB7f3slt+o
h63i8etuNb1HjbNA9X9O7Y0AYxvpYZ6yWGi7Vb4Yanw/a1QTQaFEyE3K40y+WyVE
kQf7nMdTWf/R9TBMmSLu6QUtIbKzkgfhWCxf4m6sR1ovgyB0xKNlT3jmSFQ/2xQP
g0oqaQWZ62J83UvB2QXFhI890FGrJ8X3NI8wUForLBQanTSQ8iRYnKoiVpEbwS79
jQWmN/NdGCPF6jkBXJtgVGS+vDtljCpFQkoHygAX66MdVFs2g6XvWFWqk9K+8EB/
ABKskbeXf8XxUeW9blLECGKe/ryaw1WnN1hUbh2SiL6l4Qy52b4J1AujmuzYydJn
IHogk6bqatpljA+3phV4mP+YGuJJmB8KXh0MLPwlDS/VplqxUAx9LJJ3KkQdD42G
aAJDNI554ABLm0bKZO+TM6kpc6s8S/3R9PXHcMbOFxaoyRgjfWoRpOPCa222md8W
kcPi4LpHyQnnmAXoJxtjm7eKDQo7CZ49q4F37zNk8EHS9Nund1+3PcvIQySRoSW3
rGV9VHbZew3AZRAxc/jD42RPV62gWFqYbWnBWVnDFZc2NT9sLsscHkpRb2kK94YZ
eEH/oL10wTjNHDEB+hUkEulMbdf8F5G/DxP2LbpBiBTVVcZYm2ZwtJgvVl1J+ZMY
i6d3v/6iVvV1DbZTilliqfCY9UHn8kCKMfrNZO5lbJ0CPQgtwfazDTeu6LQqdxSG
N6/BshgpV56j/BUcnZX9wUY51hwSkvprsjqiJ5EwKapQzRduakNYfth+7gBx1Fff
3h5G3RrUxsLrb/t+P2Znhp0tlMhflMdURsDNX2Dhsa4ClNEyqws0RM1IjLR3ljR7
iF97NQLWja+CuHxcfSy94EoFo30qrRLsQIMntxJ0TDVJZVBtTiK/z6TbzIP7hPt8
psdopkA/+2o+i2bV2NqY2JPNpHKa5GSexSftvUp2iomWwMr+rutL4KCL6c+wcHMG
GHla0RMNrpFV76Gj3smyHqbSG+X8QEjUB+gtnHRMQaMZ/gOEwkthXfUQDzo990nZ
jvTjUH6bMrNXypESxAPrrM5nwmOj5s32STySv7nBxbNyo6aN66RmxMhryudwnDuT
xSHOGD8YTkRx4xM0+3MPHMnuOhS9OmC/wru44By/CtER7aGHyXvVqe3KqFbBTC+k
/d4yoxJOQ2Jjegk4kJB9wXPIQk3SxghVscMFKY/Nxiyap3f+p4zCgxcFHt75JOeb
cBgfZtDWGru5SidL+CjvTwjS7L2ewwXPZttlRSiGpWCiSVc38+qfbrnmKesdKTyv
vwXrmzgWCxxjXdP00dw1rERRtj7IRcRsxdp2T1PDuVV7qnJP7nTWvitAyqoX6YOc
SytA1BAS7mUnk4tQboet3VrIJ9XRZooOHQNnJ7ldHCp5thu6PhLnEM14ifL6ABOw
eujIyt2CF5LjAzxH6kwn7rbBZ1iwvl3NZcLfDy+lNO5Tw8f1/KAADPx10To0itDs
C2RyWCaHejlPTC1LAch8JQeASocB5rYVsvw7YqwbQ1FaFs54rgNM0Ng3d2F1dfKS
eTJFO+pAHROeB40dnCKcR8pwufW32Jf7UAeh/yKXKeFi6fTKliyTBX8mVctRpyc+
gA6mzZnARkkKx5xvHF7PXDG7iDiFpazieS8pIbqTbzIctb1BHhnWAKUtcggEoEeM
XlUODpBlnj3tROVOaeUzPXgAQFiUG/WXccE5qqO6T2ZN3UjkszIWL6QC3akF7u5x
ejUdrwqLvsXFQewl5o+tzFKcmAzvCuhELih/QYWMbiemmOjfu2AFiMvyUhSHF3uU
IEM+PIgObpeV28f+KQhF8Eru0vq+X2pPuF7toxWEO5zyABCOcLoM2ggY2/797ToB
RP3T8eJjWvtlZOVV9VgqvjW1hytKlMVd/44Ezirp9YSlyblkbqIxa1pLLimZZtIq
O3rK0+zOQWVEFK/rsLAT8uNr5YbDaGN1U+BmuijQLHA1AZvPJe3kNozygU1V3zs6
i70CK95nmYiTkGC/1OWFg2N5uIwfysuG8frE8dN4IPdcjWP2sk1qrOEWa/UX8RUj
CXuxouZ/uuq78UwPxSpWP9nN25E4qvBLtrTi2WiLnJU55YXjui1Xs7HZvI+wcmQK
35tVMpdYpWnKDgqQFdHNUcMpdVqtMrPBL49nrr9uXAvt4auYphAvJwm9sThfEHV9
gfGCvucvRtDImq3ksAtEfNI4WJT+77YUiWtKI4G9TM7pw9yuNqC1+b/dqwU12Gdz
NWRKGpO7HYAYqrWJUCSuaKKMDmJnweGn+e9clAD3XUEH8NdLlS6v2AFlxMbc+vjU
f9RgFTWBXLUOfKxTDUjiMqXDU5WsEDYMJv+lKs1sQLbaz+9pOmD1NFPzWZyRBX/Q
GFo8P2h5LP9oh9Imb+drBOTfewIa1xO1ZEOdH0CLUsIw1v+ZFEV3/K9ACSzKe/lW
+l0dc3/46SoxoKQj6Bi6Sk+d60gIDiVR7g8WRlJWSeVWlJrNszJnoYkibPeaN5/A
J8v0fnTxlAcAzMRVwcWgzHUWaIK30vuN978WFljjelk7AzSvfsGYrHOpWpc47VDs
v+Yxjkf1ikyHEo4JIo4BNA6lwdz0GjLRX2VjbaCvhmZKRmtHeft1vAIrCeBRVDwQ
Mf1uCh1EmN1eabJjyA9aUX0BBHCQYZ0AtU/o0QxwlvP6bFvnvMPTrF/VjOTl9jZ7
J6rejbLXGbmLadL8BC5tWrGQtqyCJMzG4RE/xU8M8jrydmHMlLPL4i0pDrZtmREe
NvoiHle2MbC7AQEzIOFyHpBTYq0ZO3LxS06aIHdEU7UYEiZgILwgtIMLc/F1iEPW
pckX1tjmih5BHIhHLOFMe+vfu2tyZziyxxtpMq0x/JYhw0XIJCPvXwLu9lBWcvBG
mm/cTK6hzzkWjkRuDUqlViSgBXSVfn+wFl1ozyFsqoGbubNh7M1vCdLFrpgd7eSd
xf3fNTajtBbjb6CzgfCMzgz6d/OfuGkQQHQvjQ2eSh7Njjkc2+R5yTz4IRa+bn2I
uPcGsXYGdyGlEYUZ0R8Y+etry0bkpg6XKVfIMp3uS4d+WVf5BRZY136oyu1I1rXa
aQWv3FM+nC/Zl2wU0+5yUZma1rbP4hhQDVu/77HPaYGBtY8rvkjFI8icgXLPYDYc
5YpVQilCYpUS3AAUyxS9KY0zGtmgraY31sAJgXlC1VHLK7R/do2//as/u6pXp/x0
R5B5yrmc0msNeVrV5B2UpoVTp6z6iQ+pHn03yvwgYtVP3Z5vx/IZLePHOwXOjBsv
f4wmx8Rmnjvn/BqPTsmYiviX/8EVZC95ocO7P0Z6R1vwaA8EXYtFSq7JlhkLxa9/
v4h7o8iXsWdmt8vo8WbU/s28t+sv8j9GLdLNgIuQcZy2Ub35p/x99uuxWHq35nTd
KWsFWKsgukIjp279Cy+4ITs1H+bb+ORGEjkSWRyZfAu0cYV6mSEh1/b//rUThkpx
uBYCxUL+sMh64x0VdUG3WJ/dCFQUrL1EZRImW9WolX2lpyhN5v/Cl3vOwHbd4cQV
5wGAyE0J/yJsHZUoA/narcPeSaSLfWKUVoSy+uK/brKsL+o7aHNSDedgamGpxIN5
YeyJy8FXLq3O5uOs7OB0saE/luLdVSB3Cc/WvLzQDxu3WukwXxM6ejPJXBYuSlwh
0o5cZiDalTFiIBhY1PdCpoiwvP67/BUd6XN26fr7CXJUIVzq+3GDLoG6UCpWcpP7
mGOZkcs7zSp3yLU2PC+ShqJqGKPOD1aF9mGtLJ0vuRafshdswxi7torN1hNKBlHc
r3Rfvry2iKbLFlkAmvB+/bdbjCIXox4qyLa4nsMMLO/dcL6+ST9nrI700DRgHsbR
dcus27fCRQ3DRp7sO72Cs58r85MDFyEjkVdC17psz15qKuWtl2KysB9YRNjPePJZ
+/QbHsLYeCxx700M8jpyHvqLScpLzHr3jMPSSBZ5kLfYS3LDU3rb/+sUfUnio3Zl
0tlcLUcy9dgUdiOzBhR9nG631t3DKO4Ib17/eir9FzkCI+PpGuCW5c0Q3Ks5k+gT
OcQBwd1+xjP0T4gOPaZVJO0U8zk+ULrX7+WZPNFYoPZL8KZovLAEnUN3kEwIYfZM
JhA3gWF56QWSmQjQjYP2uky2n6vvMQlFT4feLkH9YbOtfOYaXeVmpwCMWZsp/nPi
wcmlfNi+2PFSvk5wF5WIxoGHv0SIqfgIgfyBr5/UDTxu36Edw5SIWTfvs+ykN43c
AWqPSyMVhP1RqCgLjUyqC3O4TwQ3qR39e9nBQGvduvwAbD7P8yrcctfXiUg/WxwC
mc7S5MAGCyGR54Iu5fcwJD+hoO1H0ShbAziQT805VwYkYYMRVfFh8U4ZxCnIQqvg
U1GL0Ywx/pl9jq7+tQp1BHxS8CSxAvVcYYpnGJASKD/qOjcZu0GCl2uhrSPWvyXF
0PBMnWOs4gvjjuFs3gNWoigN0xJy3boARLQloainPgZ3f52engkBc/5vU7TRNLGQ
pq5Dv2ZJKzB749CA/0ipcmekptMd42z9ySWmGL0L0Z7huJsJyPPLHPWGasKaNprK
Rmhx3vMT38xrrgTPmlVkXZU4O+Irq40ZFAZgIVT+iUkC+p7Hn9l4YA7m3ZT5ax6j
zNHzVBpR7WhdExBkJE0Vvt273IwRHe+SrQlc1Qz2TnAo2iylhHUz9A1cbf9lm5aV
wfQQZj0SZgw+7GipV62sxfdCHKyl2C3E4XfCENdfdhgI0jWX/UouVXiUZSl58da4
bmCxuQVVG8hLaDfjS0yCMCzKE8/9dXSfhi3Akdz4T195c9UcdZ1iCGFKp3NFPJC0
FBVcqykTlM9mCDAW405chDx8dD0f33xwe5UNV0aE0E+Pg9blVv19WEpZUX/BCFL5
JIZAZrtZcQsXCNKOCeriiOekbcqheOVvULeoc/J1dAV5p9fiiCSnL/nVQNldLmxW
4wVr7dOSaMhqpyKsW0wq+g12BfrPrk1hPxiIjaHkgZYcYO3BjFT+wb4T851WTF1o
cdwNeh8uQdNmqykTP7eKiZvylVHjYDy1zudS0OAqPPSvp6Y4K2lRRRZjo54Y3mNl
R93qT10Zszc1fk6W/3lKKQK296wdnDnOgfGUBxWhUQNcPNFOOJsp2U6IpGlwRD7C
8P7YJvlwPhSKfEqPY8g8yNnD9PYXq0zbtnjB/r9IdAi65Dqxx7NQwFuC0IMv8jOq
VTSvKODsdL8cbQ1GBzEwCFOhuoSkTA+knmIBNMUc2SuiGG8y/uSNpyDFlLa+XRYC
DTv3xVb5I+Z4pqHlcGwlUUOL+JQpEVOvay5hBkqbFOLtzosNfnSZk8ukk7q02SxO
ZK5eXJcTNNJu6019qOJwzMwJ76kco9KbA6pIwv+esOKo7GY3NL0gGYowZJ5MFJo9
P4AqmiFDIvJxWM4pKo1u0aVXpNEoQ6x64TbKpBp4g5DMom0MvdWVlVmR3/dLMpMy
PnYf9VAighR2Yhd5Fw3+ycG0WpRTAfKKk8hUatprSA458tznO2Y9P664pyaSIHs8
+fdg9Y0t+lfXOBZzW/qX1oiKnhLsTF9+i568s+ax2IMr6JVv8RDaHeX+0XAzS/xZ
/SgSY+HzFIBa048pvLCFBNdlrlO+OO5tbeXZ+RPf/kMOp0cIktVQQwjfpssMrAPG
LrxrZbSV/R9R/VuSAGRUWMIDwQr7p2XK+h2EqoQLtTQkB5mTvLOBl20r5LMcECnc
bgZe8EJS+U+ZXlMfhNzKQ1IKvYoG4n0iKWphyzM8Edz0EYIJWN3DJys+VKi6S+p7
r2uS+x3DBqBboueUp/D04LYgjmxXP7zPsdMwQ2JcyofPpvm1HxCZbxuZUFAZNKnp
oGMk9YmNTcg0lVl0AviuuIGJzCPmpKTBK5ZzWu/vSi1uOxgoTFFjlzZ9s13N9vqt
g3Rhix1q45avkEb5RU9i+eLEkc+6r7pEEqVczwdAYIjGCOPghUCNzt4iVm9rA5Yd
k9xDVFhV/89yByqdCNURHaSfZWnZT/MtSRnN7qofRd9F6uoOcyXjowYFqXBEzXsD
GUJ16bHiKOjdNA4tjxHsAJylsjIRu3opsOfFVVE1xK6U+iF5FJPGbGH/qAq0C0HA
alNedEJlpUUswcrJcuPsuqXu13lBsnbyTDof3DDvqPs1ZzCC4ImUpuvCqDT+sq4q
NHpZplM43HgVtbdLjirvi973IRV77qBIcqzRfmMNoAwVGYVWxkIamEb6bLMzRu8S
5PkzVxGGPMbd2jL/9APSHbGl0LuMqwHY1TkcxKkrBm/ucIcMWDAs0PxiNETnKkn6
Q/3Qa8WOYXrubKlV1rxSBuwV2+Qgvx3jYLn5cy8QOr+oj9pLqKBT6+XzEF2/86V8
uxAofWoqKYhdfFpX/4OZDvU7HlK5IB0D9jaTwrQoPp9HbpTAZa9OXJrJY7U0LyG4
LFfffVpnmmFNFpIfunaUtOpi+ntcabc/KE2A66OvOhcUrJEoWVgH+O8VZD+lkrI5
dElTQRjuzlVT8Js7+hrGhQR+i8+yxPvA7aUC9fG5D1a+dvIJ+pJFmsUAa5bb/TGa
zknjox2v2W9Ss5ndCM9QUYCVE6nRvFtglA8ul5B79OMA/dZrsAzPzMfJhzoukCuR
CXM0Z7Z9mYvxRFhanpiavnY8W8OqI+aDmCLR7VXdR21f/TkjXf+rxBOW5IL53Gvb
ujlmNTBck8Ipv2FPLEpr+D6GONQDyDOtWotE2TvYtUayIojjJGTEHfCb5FCFLJfx
QzyFhFZ2MU+dlwA28UfAe9xBVRVOZJErf7HC32HaWZuKl2FdjaYFA789HGJ28LM8
LD9ixf9UzJs8azTA0fE+IAmozFZSH6wlB/HPobOtlnM7Fw/OFJucdSVGyuwKJti3
8j9+Yt8KmoKMJstEM/SrzowcZA9xjXrdi9078hvk3dthEqa2I45vXTdDLEY27FlC
itGiEMBvwtlZJaveNzOWz98kRdfkK7jc9HNGZyIM01fvk5lHH9c3y4YBHzfxpyFY
ey3Z3gGEYZcf+U9XZvQjGfGPyemN9TKSRr3/pkVEtaGvjftrakYf8C4o7kTmCx8L
+yGjKVboJGRDlILRoUZlYZ5i+7U/Y1wCI86PI2xIyDSXy9VtLGfkDh32f3NSwCgj
9KFKdUp7O4/Xy66yKZaFHccAlNyBb8Y3hEXVfT6CxwRrpX29wvnRbghBPEpn6oLW
b1gHHtomCZGvz0C4fwrfh+H7Cb4Dvjc3eFxNJOX35+Kl8opVJOeifHJSGB59/0qG
KXQZuFBhzK9AOh8BUddZaM/vfK+V8bUXv7uehkARSVQyX6oKnzg6230HF1bNkQt2
nSjxAIif4UlGuGGMwJBzcxK7VstsVtATyw6Y3pZW33kxhs1JGuCvURJ/FuANTwzc
wTcBPTjIP7EKEGaihLxBYuV58WF1xRvIZ/6KVY3aapyJA40RX6pTq5UP7jfVzFAa
4pl4MrnN2X0OGTDie2NajzZxEcYjeGqDXHZVzpbfjcw+xGRpZEPJshJiMueV/dkx
+shHnPgi8qD7AuJXP8satmoH1DwDgctK5UCKzhGVz4HRRYcGtOgCnkeiUPZHpKAi
aGEW4W7Xz++8bkEKExMnU+/oNQyz8KU7quqIf7B/81Kv8XgtsVLsIzJfId8m0wtN
o+8FpGzXhROwXQmX0CVrozsNGoOc1sNleixyXv+OG5ZByRjZUv+ebzDkoNF+JtqI
0eUscOgQHQGpxNo8jzjRBf12x5aPIe6gGLGQ5G/OQa0a+lIzyAlVnOIdsGfgCsLK
BxG70mHUdrReyaKdRWcBhNDJ1DTba4wPNcFd1iPI6RewDIV+xKIqoC+suZSWN8f2
WiBTNd2wmywc1gOo3fciSNRkmTUs1oYnYurf/mTlHuJGTiyyRxps8esI+B82/av5
Uirb4e7aGYyzj1grt69tHkk7Xoh32SyupXneAiUsr1W8l0YnsKKzqQbE/8f4LkTK
2v3Zosw35QVv82TPwLw0KTlrUM6+6Wleyn0UDgY/61r5mXqaymsOT9SfdTf/D7Kd
1Wxa0DSfpl0z7av1SQZloOHJOhD4vn9oznd/v7fVSE0y+KsFsZf0VDfIeCDnglfL
y2BsetDBYBaBvGg16uEfw3o+M3NWgO5+ZFPXt7OBSgslNbQNXzShgp0uWdP4iZJL
gOApdDHsZL0dgtjvJ1ureZ8CQ2yB139Sm3Hmuk1lyH5ipqmnJEsnnj8Lr1GwfSaA
hvqlmLMcisFwxgFZfOSwkcxZdERF0vAX6iVkD2Dhn8HhFRLwXSBqyZcBrygtLkkn
EEbBZvS0UKhLpLqk7joLdxchuiBm+dizcyMmXrj0vEr1XxLg+EaGP3aJ+QsYfcSG
4DEKtK+Gpk5peS1zpIsAbn7ZQ/dqbWg9UMszd3VCkaqDROkLa5c1IImELSOwCveE
72Md+deGP8BkDNkG7IFAkdHvmVmYcXEJrIrXbZ2CLKVGSoEM3ktdbUdwdL0Vpd2P
nuVDts7+i/VnY0eN2Zycd0t40Xo6cW4+RanSR1NcDOBR43d9+MWzRcVyd099MBMS
I1GprxKzF5TaOT8mrxKlD3xItlbXHBH0jkqkj8O7Vt5yDB/L2j6KGKbxh5yBSKUH
zMLKGmB2UeqzePd+DZhEqqSY6gJZKVUznl7ktqmsx+2z6BWmFPtDoPST+wVXgP1B
B0bh04Op7v5s9YjO3i2nwyDPQmZztkv4ip2Tccd833/h/nsHbJWYkr2nWZ4A9+iW
y2S00SKD/Xjw6s9dXZsZUnJVa35cwagAexN0csdBRwLLYR/nqSXvGSV5CXVQVyB3
cpgeCVFE7S79kMwtrXW4suKqiamym5BUeBlop4jMeF8ZlgW9glnPBzzsUMiyuhMC
U7yUHcR5KYKZLOoMca3hVUXauleRWDz8C9dkOFArnk9kbJkGI4Q4I270J1QMcX0Y
JVqHc/wk3o/DgOlAhZbME257yz4NgbSH+pkJ5sFIjr+BpE4VKnR1OBpdM9ICFf8K
df53Nqh1iPxHAH5v2JG5secsKQbX28U2yb4BXBxjc8ZXBaCOqmfRiofXZ5Y265n9
vPmocfXbL/pnyaS3yjuVRA==
`protect end_protected