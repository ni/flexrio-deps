`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 45040 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
HDP29p0vLOrNPcWDOvry+TF6OCVUU03uvcyfNvkFCIv/qAnD8JWBJDl1WsVCHZrS
7b2LKCSg51osBTUF5thf3C9s6nt+3jXK3Ekw9kSX2ppvhevckLgbEs24nkO5txE+
9QeTaGVM469gSlc8TvEVxpqqORxwjKmtxKNvCose9d7HkioGVmB/n4fDvnok7ab/
NEI1/ZGCELu49oeWxj4TrIe3chOL1oYpsvSAl0zbh+aC6hojIp3zBmbRj7D8esFI
iRgIw3wizEInPhkvnvEVR1Qnz0hKG76PGWflQb2CPIKxKcD84MvykBXZCTKXZy64
bZNrVFDgOl6zS2BYSaZ4r1eTrRvemgMvyirHke8/afTW54vrl/CQtwtWKhzwbA68
WCF5QoK670z7ERHKcxt17zBO+wKM44KSWSTvnoy47xweMFp0fxqPHspiwFbS5ooN
DGypVRvcj9XdS4I56TxPNG2TvpM8sDHQzxpCe5lA4+OC816IXmu95iUgZW7AjXVe
QB/q2LJikw4wW3HmQdG8m7MFDO5YwIQZffxNXPQkcoZhgiSchvnSY+S06Av8sGoj
QgOx6r6wchl/fOzsagpEBmNLhuNwFErpZCJPnh5fvU9HEMPwF/fzWB/+HNSCg6Zv
3eQQCO3emq+VwIWF+HdT+oIa0N6Z91OcYOuwBsw3zeA64GZK1uorhb70QCZUG2Dj
y6GGFW92QRRA8m0x9suruud5m4wGHAZ1eO/ZDc1EyOOoA85BkaV/iQ9DpIJ8HbAq
qNwdrNJw3Uz9XuBNd8FCyt6wcO6lVldn3ATUeRTbcKFKDDJKWrQmEraZnz+twx0q
RuWprPkvMBQ+QpASD+IGN4RoI6iet4maWZhoCXIgn2Noem6s+Mtg/ZQtGJGhlE+q
wkIYLZVRLytsJzy1bZgW2wyxNgOED47ToXbxo9roNXhcjaYCV6StCJ7ip9PLq3D9
9hcwhb5DOYREfpbjKz++OTZV1HhUQIQCt0koNpbo0Ck8xBzFBLPQoi7MFqpQDwgQ
cjA8FTQtqxv2FqmIJ+6O9YPKNLVxqsy8b7IKINWQtlXfv/K9oOogiX81QNBf7sLq
SmAxIvyIT7irczrdW2i38gYyB17ODqvrOl13T3AnHZ+P+fwZFYHn+Xu4iRMrAooL
4jRwRvXXoQ+bhH52Ztq72jYq0NmSQ+y4WDtcIu3UG5kD0ggYC7JjD/0p0b1ZoyN1
+JwqX98/b0vlKcEZK5/mKB2bt/k8pfrdMv37J/vCONrw7TDuZACxg3yBoYRujOcr
RliWm7AkiqWeVdwMqbFXCFXe6g9CAuQongCaqgAkTXfo5AqGW0ZJ++gFrJBPC6d0
3NW5Du+H4qDDhw+1BCuLUgptWCvxhCgQpn12znRSa3LNbXvA4SrOWBw3NQh+BGyb
7U+/tnjwTpzK1iKK2R2gnPSu+G0QObLy03FHCUsDg5yN5QDm5tyaSKoUcYviCC3W
KIvn16A1UGoVRqVQJPikwP/wQ5VVb/DOu430LpNwKXGNBDVCKD75iu8caGZyH3TS
TFH3JnvKsYeGHwe6/GG/3dGRsgy4U+nOW27RDHXwepRzetXiEe0SN5AwOQUq10DW
3C03/fj/M1Scr1AzS4QUMNUXsVT/yVQnPX/yioPP7s5CeaXu9YeYcxeRTdpcM/kC
Q1gKsloF7ULh/JC2wrRQPgadSjrs0SNbXv+cC38UtzhwwJeXATsu8VgVKa6ECIoA
FrVCvgTBj8UjS0z4nqtRb9rvpeNPi9SzkUXN4J2aBa19D9jza4o9YsV0E+MbezKs
SAqiZW8LrRsUTJlFA3rg9oMpIJum/jBl/L+bscn5C9BzbNgwGQaXZrNJROyWlisI
+8xdHtDEA4YCgPiWCLuhE+eB9QZWd0m3eoGBi+YOFBEOXIoVhr3rghByhoIdyFNb
8hxtYAnYX+YZn4gX0yvWjkLaQaKUsySDhf8LJ/j2apEegzCFOua70eTAbJZygp6K
iHLKYiiNGdTJ2voqGz4G0zy5ui4ka9ZIdHRrbmF6JHCxa441su833Pf+7H8u4Vt2
wiIaJLVgV7MBE5XQtYBhuIKvfhgxkzU2XA0ZWiZKLyjDsWKOr2RdZGiOYi7BFtBn
aRW2kYYK19g9aM9tLHAFdFiH+WSO937mWHiQTtzeHZBi63S9zr4LxQ+vljvBZ1BZ
g1rB56qWzF+szjFt4EaHVZMm79No/pWVoOlh3mUJ3VAdn0Wnogac4AYWYYbKRAPB
g5hU8++nwWpiJ8VyyjckRhjZ5vNQdiE1PDAO2wGXD1pKV1lYIhBFGDxFsQsujTFz
ohU4QYJnVD91FA7EyMW8SUDwatNMbMm3bs53Ao1kTxYUmGwqA4CDX8UOKCUPZ/Qy
xD5B52/ODI25c+Oq0bhh9qT4yv27/Senk/PNcvPOTU9Ym4pLPA3xndoLacTAEhnq
KDnZaChEGVS2UiyONTMZjlDfrWzo1j+fqo+Qv737rZY+pAPX2QzkT5vGiJDCTGc+
74claFizWVGjmH38fUIflO0eH2v6V3/druYB+0ny8E/8SN6+2MVuvj+g4veoDGNG
Eqh2FMjUjWpD3yTV15aCqg7pYJNxJiL7wrYhg8gpqIR3w4u5DTIn5mff+wCmptdZ
PNu7BKupvUbNOJqwZxf1wS++QYNHye/Y9s0BGPt/chUp5qVZSSm0hF7Cqj6kEGun
tdvfDL35QXZadopg5zXy9MYyJP3pA5n2YEEI6y/ffuo74j9KvQAmva+suvl2LFCU
WeciUK6o/xZvC+TulTvZa4J7EWUbRlD3LcH6FeM6aA1jx0BXx5p/OPDkqF57EEDk
frIQCrq5lhuFd8tbRnn56/dDat8nLaSLnouXVdqyS7IMkX1pNHzheHXaDRqUOj72
qqeI+xwzIuKhemt7REgI1o3LNFSXtndaeVURO4cdEVUt1oOtLaQhV49H3hfDNy52
BuYcRin+sq8R+K5jWdgU7mAhfi/BY+5qmszIrUcC9zL0v9y/q02lWGRQofp+Hv/h
+XO/HIV92D/OtKmY4uB6Heg0UAX2QQT+WDekBnoOpVFqxa5uXvx01af15l6mlqXF
HJho7fJsY7HbeFN3C5vH2hQr7bbUZpPWOYtsMB1eK12j6KiL2tsPDWmOYO0sJs9F
ovzGM0u+izGfFU9RzmHnhslQ5CsK/4TNlVqpxGeVZQMjuq9PyCuPGd9Hjd0Z3E8o
zHN1GTNCzuCYQnseQ/umkWThE2ZtRFpiyatDMgKw5/2Kf4fJ6sRuVSW+N+5OO5od
yiELToVJSae7XsmJLH8++m2qoGssJnwYyyUAsMgG1kHicA0CUdBWP6fIIvisvRlf
cNAEnrjO7Fln9AyHNdBT47CX9Pe8/LzbIxfaSFvdvBSVA70JcvIK6oWERpWLxf3I
AsiLFDb9HaTYQjb1HtZgxz5KTdyl2ByvMiV8vDOZWbWlVJYga3dBBdqmbtSTlML4
YICSDTFMP7dcRqF7AbmqPjWWE89sMxcVuFy6MDtzTusZmoahXDrRzqbE8XCBXHeJ
GGtxOAc5tt2TZKEFNRn3KfoKdZLtOh/2whbmx7nbwuGpPdpYw3XwoHVw4TDRmjfp
426f1YrCADyLQ5EH5UaEsoEYh29jLcyjZf29GKjw1aG8K4UyLTsfeA/weR10P1at
INe5N16LMc446LrrlN5wIpF9HsGpl5CDZpfGwlnw4eWdP0xb3+pD2IH4nlk2Krk9
3kIlpNOW8zYOHWKwtGT0SGQAItHiFDuiBZ6V/vi+bwxxbi0t4DVhvD9TgvLJF5QJ
w6WU/SuWVe/MU21LUOFvdfzMUyPhEURaFIZdwjYjcNE8BkHuNhicF/MfKdhkCTWe
DIhbyIZxoqALtDycwoH+7U3hKCGPRz8g+htzM5eSh6/AndRK9o3a+WegS3ijD7do
Ylot5JzhsQzMreti4knROpmHBJTXH/nqJVjMbMbKeBh/r4531RGKrkHmFxbPOKKR
LOHC9wthA25vAxHe5G/411YJ0dItAs8ez2x2tSTbHzLMtcqGQFMq72NHyaX0WCbx
F1AgmwKkUc50/+SHrkQCfUU25daNMJEbD5VST1AhK3dalPSmXKhyo3DglqT8S7RA
xRzVLNAxnmBwgp+MaEgFgeNKtr6Rgnb9RVPbJiePdB6NMh4zDewf2ha7/euivxIt
6tRkdxRHyZEAiGOkmf66YWIzNeuy8X/3pzZgQk8j09tHQ4w1mzrejvm7jLqCrT2f
Azioja8Jga3nOJWMsn8taTEDAYEYprCQL5yKcUGnmwYE6Owqle572cFBp95686Sr
5+XHyzCS7duc6DnQSLlCicWbH6V1Xxek1tGBL4mCfublR1Uh3xvDOpI4hDg1eAhT
Ayi7dANbup0yS5zRNmSuXXgzPW0AMfsx2l/MoQZqc8VE0DwIqVDfFuiXqggmcU5z
tx7kgFxVCkLe8VPmMdMQQ6zYvvTh6QsQQMWb5wK1hKW+c/UCMcgYYo9duUnc6Gn0
1WuEmqVirzU5GjthI2TBZ1ZpokUqdFrDxlLO26hap/ArwC6yOQSa39VtKYbjUse5
UettSSOAnI5WaApPKlnXG/MKYVjUe7X3N5sutFDdLYFjbaFFkCN58+HoYmZ0VJVk
GXHI4L03ECdH3GGcldJ8HXgrjhxmwTSeee+WsyCZrTv78BmtEfv32HSlAMycmAJX
E6DX6saMdDIaYYreNvHkBKk72UOiQQ1Cw8jI7Zp2tnBRb9E9oO3rwDpVf6DecOKb
yx4oKpUS55yvcDletZoVm3qcP9E5XsQlD5wTeyjDc30mlRJiEKajzhiPg9xTuxBk
6zIJwXpVkhntMInKAzwjbGjeWpR/ankbR1gOVg/Yd7BpTWBtuPtSFy3AkcJ+AyFt
O1f+NA7QI738JKq+n/ZGn8SauIO7GJVywcYdm2VbSyyOIB4D4QZfnNJs9mvWrgGi
jiAR5jZls8WumT5YukeSjTvOndnt1NPR5OZAijcBy9YuPb49Hoz8fp+hFaACdKo1
aHSDqQQ39dIZp2ExsyNx5zt+kuX+P+BOji5NT74epuO4BfHfwQ84Zhczi4lsBcCm
B+Ozad25x3P203CoDt/KJ2SO0P1Nu2M7uYA3eQeLgcUNMAZlCsbJa8wlerdcdyW+
nXgV6rJDDpwaqZoiSgwfnflVIia0NTqx4a9+VIs0jeW5OLjjfr5f4yXzBghcXXJR
uepJeHBOGAxzKIfdkzxIFa/9+oZb5Rvh3905pPy2yXSKxV2J4soQKxCRSHOvvzJA
vLYqH/Em9ij1h6SmhZ/eLdjeOA5UiAnRbqohsoOFDO3QT8zSMrjTonOAwK6h4CTv
Yvtt2NNebbrGJYRTFeI4vP1y1uD6mkYbN+IIhoAy6BZNhiBbH573td6cT3q8rlIg
zy/5+YRmYBwmMIfYkechhEhbd+cCv/2p9i8GdYCxkMuStTLXWv9UWpZaW+1j0RIa
4g/hVZbQl9iwzE9KKnl3fiXkM2t8SY+uQY+lfat3FGK4G7Y0wR7mQVMnqSBCxBY4
YvyftH03GeOZZ118ykqaAaBzZdO6i5K1x6jBJe2/9JDXbkjkxFJROfiKS8x6ceOL
wS2SNkxQ49EtdLmic4t6nqsue5oYXTAWLnS7MmCrmg+s/5bfkg16lWpP4jYVn/um
5rFiD3lsLUa0kYoR1B4d44GGWfRgwLlcyCi2YwJrib5SAa+R3ixdeDFPJNu2O1NL
ffRaSG0GFL7eu5eIclZYHof4HIx2uIfI38TgY61mwh/3s0P1UApbKnSqFhojteGu
o7+1FhQCXNw6PR+2V6kvLazGLunQl/lpdmzIP5Ao6prPRaUmrKnXeseuqYIhEbqn
K2irCqSLhaxpsy02j5Re/s7/DHEWUcwEkJ/h8vK4LNXYQ7xbTAVw4gqCu+a2y7de
CswYWJzWlmpL8gLOr50Bh5KbDxlenO8PYshuSn/z362/tvpW2/e2jL5iyvyM8ppt
URyqSuZRFnqqVo9zWPrTbibbAI4pUSlW0WIVwahRHezxJRlQIzhZLyCJ+q+/MSxS
3w+WeHtj4gbCMwEJI+7Qg0npHHJvfptfPdo7O6oCJjF2iA1aT4MhLQcKwmwcwGd6
sLynUQBuX0x3skQDt6r5U3RNb02tNoDERhl/M4+XUfhHWKAtQakRhSZ6z3xQKn2X
cXwpfAfly2lumPoYWYZ/PRKXYCf/B0SnFtAcauOb6nlp+mLv7dd6bHlTlIeSyPfX
XeVwAdrqMTcGcxihzrAh8bQ3rQ1wj3eUwOKo8YpMgIgNsgeOgJgXkqtecQZHjhmu
8hvqv02OW9t20gYZdlsjj8GrLY4M3KFIyVFxhJVC+gY/j1Qpsg6naHkWZK/ftMWE
9F4hwUh/GIJC04zBFBGGnrwDybNIYiozCqqdIzd+KOJ/vu2ZzBILTd02mbh/kIWK
qvly8JMgUHBmtjVz/EP9mIX8mmkyKIbRWLHS0m4tAiARDxkQhH6an6mA1FhYfFEj
n8vAlb8BlSHvbHNPDVsG3NONevAFWXauHjNPwMkERMuF+HcsR5UCT4aoGcN0QGH4
2hfhnNhJufutl0KUMDqj7j4G5iBf0qNFdXb8gfpVAreUXTjoXsXL1b1cc1TIYCGt
/d7AwRx+Yjr1JS35jTcm6a+1i2glBdhza0vcnRxQBcPhQzrFoRnuoIAyijdEpYGb
gO12FdA/8hupRj2GldW1prRxAkaQPrmjRePBpy8iKw5ghfVIlXJdcGlkEnMb1aLM
bM8QrPTaWut0CpHmsqXzTzv2DU4laQPYC2qqN/o/mpk0lERyIuQSYoyZYDWxas9O
1Xix8rwzpiCBF61dD4wXY0zFuvYwJ1oWMW6ICDIeINgKSL21OnVWDU5NdXXbIn07
q52eI06t5bZIFlra54WmbjsE/XCVwq6XcIheCRgvIhkZJoU1Ui3JVKU0z+7mBZJX
IIoAOFWpOYKuyILGfbAGsSEqU/RjM+F8qoJ089Kvys4PCGdKzXe5v4ZDOqGyuX9Y
oPGbQaerQXUHxSW79jqbeOWtuNztjqn+KayRjlA+OwdjqKA9rWqJ8uIXsI/Y70HI
BL5bYcAxK8ldt6MyTNumhhhONq2d/cBh8Iax1+2qm3AKHH+fRTsyVXoqxHeZi+pi
2E8Gaah43S6pcsv3TCBrabzRc7M/4mfJZSCMVXWya7WpjEOKBp5gDiGMGfCjV2GF
pe+tOKAMxbHEkgdSNHPQGGZ7FGPCIUJ8GWmKvXVzbMQEMR33/wF4eMo9RRSsXpEp
vz5J7J+AT9ljn1eL4gYZ41flVRvQXh/Lj7BZ/xlD2V0ehmoFVucELs5Atbqo95Br
aIJ8H+XfjXfs+rnq3nkTvBJ7VQOVjlULeLAKR410UDQqcaRTjlFNS22FSXz8ZQsg
5zqrqtFoF7KmQYHyXVrupN4S3zaYS1ZG+VxBlDNkyAxHch9JssX2rbRvgqDp90+y
72VqiFpSuiVdmn6Y92ju10IXoHqTyY9GCqhi3oAmD3TuRfLngMvVqbX4nbkd00SR
BHCvWhXpCJuSiGCltnDASS7dIUaz+Z+A9WrUi1SPTp1G+aTgTFC/taTM623TQOvY
ckZ1ROcYvGdz82F6LzmkfIKAVlWTZJcYdmelSsvq+zb65Kf4essyFOvoNfkk8GsP
aBh16/LlXZFQ6thWS3imZeOAPvTLkTw2ZZPe4YO1FXWTY3x2lW50cOR2oc2V31eS
4aTywL462o9YQpkOV3cwmQAn9xUdzZBRRXSpY1Gn4ZPHfuAMt0u5cX4f6tDLZ7V2
mlcqJPjsHcNrV9Qu+3pFtOfIKTgHyqN4oI/aV0WEh3xRJR9E25xTwlGdrCigSyz2
/AthmYnkrA7lhuHqQ49xZGzzVNixlDss2MWwjfFP3mn5PMl0jTinLgC0Z3SfhqkH
4sC1UnvG10ilHLmhwKsVac65QN5JvqtOr3ph3eBeuIyrf8ZVKjdM0Ik6P32uSExq
Fdq7j1HUHHif+uBGX0KKHayD1Jay60H2ajt3DeBS2OSoGhIBczH116VvgxByy27y
r2ngNwi+N7Gemb5c1B4xMWjXEX7eb+AhrN/4bM6+TX+lv58t07KtdNFW1aVfgILA
BTpf7M6qfVhSluETbtjSRZHiBG4MkJYYZ+46/M/JUF6R0D4kRqc528IwzIuEQ+Sj
RYHYT99EiVZhUMq9FsCYSJCZqCfObeUV33uFZ2sPJko2V6psXeyOkf/lkqYV8sFE
y8Cjy+E8f09W6EBXsHZs4UJbmMSxFoTjeDtWHu9Dd568C+N4ZabmkOWbjzmsIp1s
40LpskTkMAttWIhnyJRmA/hyhdM9T4Nq8qdlqYk4j0hQNhXtqUgBZvw+ishiPDD4
sFfAyDHk7FcAb6JnqsFXQKCveohIH81j3AnefHjLrasfIo5ztI+jjnLC7mjrwd3A
JxTOnUJgTBHa7Bkrq8dpe0RrJKewJwr2Hx0OC+o0dhfQ8zj6xwSJPzc+l/0MOVvZ
vSr/eJymHPUjdebKbTMlOvh9aCqJTpxD6aSTtdukmUwmzf1NoUQ4Q8nuWB7BDchX
XOrtn5r1ZX8xOdmAPts0y+sfzRdtw/tduBgMi78GCJKtAMNbXgdqKxdJGBCP+He0
7XOsPNQ/8o1CIxY4CuQSoPhLckCNKOb24GN+C8v1cUQunnZqEXh0+teKo8RVDbG6
/+P0ffHTkaud1AwWit0btBhMQyAxJh9ehHABm5fUrIYls9al3NxGxSg+ZZ91YzJ5
YlgdMQDsFhf5s3BGKwo0HG85UG7u6xP+Q5WJqXRLhydockN78ifXDh2dnWcqwXIi
KSaiG6pagM3lMBiV2SEe20iqZoYQv0M0n1FBra7uWVEESFwE/RXPcf6MBTgn8Fb5
eJjNTUHxIFOw/P4zM8V+qSbBISvn7fPlMIQNKtMJ309T0soLFH0Kb8SFpPCsUu1U
TQCmDE4HyKT/cBlCxDOIE6feuWIWm6JdCu5JJKhkPMdeL2nLUmbpFCB6vOdCtQpX
ASZokcZHwI1AIOqSqFQcsAEjsjbUb0FZDSb67fqaVsz/JY2QEhC8YUMf7nGECz05
AVSA2oAu/8iAkO5AHrf5QG1+PYhZFFxoN/9FCdrgAbPjdGfrcRtW3H5WBmaXraQn
WbCulEltdjUdwx/2BPSLZXVIgO9CjSm1BUNnWqBtIycJ9MqwuUxa5rOS39LbOYiH
9VIUveYs5b7ijYq/uEZDrRxjAcRKCF4q0DbvZUVJzZHKGOqoenRaas8cThBAkb9A
fvAAGiDrNjT++tLSId5q7Ipjk7vu15ETb/GSG8xLpJzhlWXjhM0ipRMFigZ0dJIA
yB9ikhp+6yUJq3psdNYDhHAyLjRuCT/O0PROB6GADt2c2papySt2pcGWJS9sdwgg
l0u8rJYP+ayUKcCnqQ+sPcezKftPfU5ukiE6ADngzYdZn6An9tgEfw4ZSg1bxsgN
WD/ja/ZZ7HFx8cnwVzyp1AQVWk5YHTeOPhRnAz1X9sfJcr4mcvL1MivnNGWNA7at
Ayqinw+dZpL5UxpuBILJWsuAwO76sg/Q3K35aFTmAE+SDDomryactMxU4jOnClNW
y5q7/3/KPeuc2tcmXOx3QtauDQJytGh9W1FXq2DAmN8v9jgQ9hI/Fo0uxB1OzaCP
jjLB1A2mz9YtbgEqF0B8JTcMnG8+jhdQXCqVjXZeEHI7dTQXb4mRy4bYlGf2WVIR
dCXy3R6VFeCApasG6lPv52g196H7tnxHO5g8gIGQOdsQNsOd6APelVwYIGkMFSgL
MoG9swjtsMdIOQ/kI+gjocFqWLbuG5tHEK0sbuXxIez8BIlK7eMxbPFyRDO+vx2q
gPi8HTioCx/keGcTBq/QpIpG/qEskUXH4KW/nuacJglvl6HkI6SQEz/GUx+rRSh6
YE9n3hk1/yfBeZgc28q/w+QRhcJrGQ167IUlv7lU+ZTvxEwAVr9RtMrcmOc27ylg
Xzc+lfr730liXRrV3+R58FFXjdwN4lp5vcd8nuaQes1ZzYc3A4KEPR+LqL6zXqjz
F7BTCAYKJQf4BcPGoNsiUTKuhDbjIJQfFFQg1p8CYHg6qfQc+D5raRwFVF/2iPxP
EoYoqJpTWKLxGWhVZVuMATa/ze1fjhxJ64X2o4f4XxI5YnBlD6W+51TpTJEPcF0c
/AwyrIsEF0elXWgKJLk87fn2C1xL7mFVm7VXGEFSMP6QnufdUBv+kdpVoHYLR/NN
gSNJMYjhxmriOeswBvy0bOFeT9CQjN+k+saWqdxxBVSJ8T38QjwXaMSbDZ/ElCMa
NizcXAXQy71W8Lcw6ep+FbS9DeZoQtgnp74eE7BCsVIAjHpVUk99XrTGPgRL3lyG
9WpO3Y7lLYOhoOiLBaJgKmP1ZaA65zd0+H/lxsbiVHSsO8HVHZQChlz0MhIzDs0X
5+OkRqb2z/1fKKfY/uKmWpr9TMT9rYqly4gLj4X0x7vdKO+cHI4GMCQcaNrNFKwg
rzzhU9niHxGe0ujTcGAFACvUwyqy3HWqoEbuiqvRkH1VP6wdPPBI/dwEP5HXq8Oy
C5J3ttaclVn4yl4vZ4/CI0JtYuTqOqOEKPPVBS+7J7dflBAI2/J87xTRIGIM69+Y
5ioRPk8eGMa2+aBvkZJozbv7QFeW5NN6wK5wAnxknaXnP6V+I9eXA11Fr03Ka7VA
x41yiKKkesXoeMgmXnFy267/4X3c63j1ZlX5lYsCo4gBa8+RJE6dZm3m+VfrRgQS
wYWp+NIo/aAfj5ZWST/75+o+2jVS7Xx3gknZGuh4N3XEdtROQ2AIuxLMW3/I2U2n
FTD6icv1yQUBB9pBNieIELJ8DDMChplNuWoos7fetB3EP3zkBenbeOCVpCAMTtJ5
JIBsFASIz4d8yR2EQQind4pIqqLDJ90lsZee0JHRN69PLYm1EiQDdg3FW4RtjaWX
Gll+R03H7JmYkbE4YBJj2wggD1SsGv79zVqMj/O9SF595+FYGCfjrdbn36RRefIO
mEJhTaIVRsQTJ8fvpXopsOTae5G+whaEQJUr3fLdzHEFTshQxfZm5BHSgIXhscpz
auYSCrOSv5QjdC7FKywwo9NZ3bMfYoiRd7OcyA5yQ+2jYRZxz36YCAPAeUOtcHVb
YLPoNkC93H60SlmsswBe8DNxcb78HjeekAQqoqMwhpXHDItpE0m5M7YJ4cgoHUlf
KfwBcW5kUakewbiVOoHuM8OYi1pjKUp5adM0jbCiBgx/J0f5M3UimWyFfouWsiEx
bxHivBkX2o+wxa3DWySvRl/9itnDwqDX0C2EYVkjeZsf7RWaaifYripvibJGu+g7
qEQOuUMsMsVhMmY6j7GlvIGRH82lVQzTNmHfmTq7EAmtKd7OwXk2nVix9B2C4fMI
zfZc1FZYS49BQM8VBd3DgP9IKmPrmt9uApTxdpjnyDe6QSaDlx/fR/vjnVlPf+34
paGkdtST15BUxiuWyU662YY0geiw3M03OxJkR0nKYpj+kkqzxp1L/0KV7zkLWUOn
H5puchrVHjnxhVRtIZbzFc4MI/8Jz2oSn9mGghasa6FwjdBpLMeuDGhjWWTbZ7Nr
hlxSa4NurOEvEQbXaHv80Wa8d0nquELUp4fB5XR46/X7ZEbESGY1MloAXk6chKzQ
QYsFooujqGh78c0wIgWGCpEeBg3RQRHc/yVdNP5WpshwAO8fFL/gA9A0wLNOiO9l
PeJ7ciK6nbkmi5UR2rrHx/Dy2aiYixTdfXlHsRYiCMJNqK/IHIXN7NFxjry4+Xcn
5dRKDBqo0z6HTUbi/UYrbguARiH3i3M8d0BwfcNmzBGDjh84nVraLxE2sFhJy9aj
HLlEKlgr5e1s4BkUZW5wQ5wSWB/7I6BhF95Yj/jLrSU1R6VKWHw1ItuYhl53V28Y
Oxh3U1zMb5gtyZcmjI+MNdzB91u/j4ozHS12zsVSzN6NfVr0xAc9MmoOTENTX6Zp
NBhb+aC+4Hy3hqVmPZT9jap0Sj38lqCY9xNMnUsjZs4Lcis1W/lxoSiNsjK9TXjf
iDGnwcr19IORPHClG8ae08g3tZO22XF6vanV9f5OzpJVd6scZjprLBHfTBEeqfYg
XoH25RM8JrMRq1SNeXptzOV9GiKnCS/Qj9Kd15ZwA2RgOPb6tEj68lPal1S1vspK
h6VcRATddxoEzGrjkYLiPlvPMoWHchbdOPh/0QUdHQj0NW+NMnMOq3BTDZ0pYsJc
jj99AgaLrbRP7junuJfsXkEELO11eIm7bvq0a7h1LfbqeMdyHy8CynEdkQnmKTFs
QmuSKWUiowYXb4D85CVubA12jBOTgD/3sfdvwpZAkKTTHy4gdtQOwSKiT6mWm9Am
q6VVZimxhPWpCPqreyzMfSbxCWkh3WzSiN4ahRPAkZwbVHGBDKC9jtsEFkLhvd2i
0PwgneX2yPkOL8REdM+RYR5mSmgxHH1gfbd0jlMLpmV/U3Mk9cco47ghqJFaCytv
jgdjf4Ux2zkceCHmZmibBgiT8T+j3ljHE4EvBqcrf6ikN3d195okw3m3++Zt56ab
l0g/5joEo5+FOPa5Wc0NT9UUYOoZHB9xkQUhQZ3zJ0V1Lf1tnqTO+fCdasiyXLNk
yNzM8UtfNPgi/zZgVn5fgt+Vc3YBRiSsJblfIXZ5zpzSoOtIUzaLdpslubVU6izj
VL9YUGuUgxd1AQuhUuqlH2GKou/FP+jvW2InCJx+WtKTiU6fO5E8bp4qDLYWBkDN
rTLY7Ux0i7z6eZ+Qm8a1/qTcTZ8dzkAEUHw76XWVJkl6IfaBtAFFxLLfkVs08MGd
xIz2aSmMkETtiTdjesNlsk7agUap7+Gp5tknpz8+eVESEcd5f+BmNhVm5NH3nfY+
KJH+j96m5n4z21rUbooD0R3A41jXnWlRZJ9QPShzALZI9762hanbji5M3FA89cT/
mUp/BackKV7n2n4I9P8c5uUgkfC1vwoygfQkXgViV7/+qz1ug+cJGderF04r9yL3
bMluozrvcsjdMYn49O/HOg937VA/6twQlXvH/TqQpbVWh75U4R3pxYitLEkLT3GG
Al0fMMNCNlMyeyrDVWM9Htiy1LDuvYPtfDTMiaChMdltRpV8e5tH/ZIzg0jixjvX
v1I1AK2EKEcA/MFROCQdsplMS+6HCQip5LzM+zA0IvoBUvX/HJgiPIkrPpFHgd6+
2Khd8zJY6mZetXNrMCCJzHsVpfvyrPqnApHjzN3Ii+53r3iTofh9HvaT8dHztP1o
yP96lsopv52qlVv+BRGpaAgKwfpjGMOuIi2kI/8BlvkHkjsH2I5frKLMJbbidis/
HSY0pKrTWhqqQJRuxJyDy5V68HDUhebQ9zb7dnGUuLkJN++a3ZK82HixR9rnfvOK
DJYxLkCMVfIRohSW6xIdjUflqI8EIj6g9+C/7RrbXf8te1jPXJMS/pV0h4Q+3Lki
O7TPjJjeZQbTKQR9xIXyJqrPF4lv6x1jGc5twRW/c7CNoUpHXx74cG5szk1T3/x1
N28tgMAQWN6vZ7UYgf6yKe0VhGzr7K6aeUGe05wri7vxanbeTQsxXqw2NcvVHXA8
8SMAHZgQZgg3kBuv2ShayzkgBEMIsYM2wXia1drg5F5OhjiFomORrAFXEImDSITr
UnTxFV6BpceokX1oUtFG7uBwRyz698IkdqaNx2iIFto/bn4aVXMdfKkzFpb6Desr
01m8Z5xvW9P0ChU0PRCG2ON5Y35syhWrTWe14cWVbregSAHs1TO3T1FcPttLeuky
JBTniKer1WLYjB7j/1aenNhI7l2w9f6P/EfMtRVtStM4jQS/zzcFSzKv/8kk3F99
qLJcV0k0rvbM/+GWnQ7ssU9mWlZ0mNpN5jKq9+fniijq9Hi8/pSJnXyU2h9BEEcr
zsFrXkTliJYB2DHfVSVIkkvpEYLpluSBdKA9aVf8Oc1lTSDaFU11MztsrESSy9ON
FlJSsa1fCxs1X1Yoxb/J9M+cgZasVyJzAnn/qnKVK3cX9590np4HXeqmsKOf8pcY
fOuss1avBYZfJGG1b2m80A90S7eDdZQgFbaO8zQT3KOlWK8rAwzI2VREhcwsC7jZ
gSQsYUVq03BPkdRgrS6huICrizw998LC9xNb34X8VgZKEYGUCbzUlpQFM+9fQFgm
S31XANwJEQtPVwzOjscb6M/9aXMI+IReG0jwg81IRs/1KRY/oXx9FO05CgrMKJWP
Cw0LKzerzmdZ+t3rvd43PFKw2gx/QCR23oY7szXY9Zleb28Vlc+r7kzB9gfxp3tI
UHwWEEJaQNwtz0z0JmBq7JCeruIhUprN7lMzJLECLEhma5JTpfoJFdzdKwtuXout
KGExMyNsjUd4t/6d2vbuGeJeGLrd9uOS+LFZ31xJQQ3NqTUzUCgsEhOFDTkYpuCy
RMdyoa5WAuOMzJVSmeniARYihCFqzF7iVR9PFc4619hCJ6v4nW6kQJm4PrF9/ULA
vfH24LBBDXcxX9TaQXaNgmchUkTqJXq2rlAceZ+hf0IRhWpI291uPHbCRb66Ag+t
aLEklTFweQ9wWiLuytTSjRmaM13h9qup/irplz5AqN4Eh8XsBmJwNVMCjauq9ECo
iSUKQSPM5CSvA/RJ9JCJz0ZLVDHR68v0rq3E6QdYaX6RG0BgY5sYj/DWdBwtssIV
wVWdkM7nJbTevjE3+woHty5NlpmXM/wY7OHv03V/Q7IQyLaOLmoIJfVsKRE0KMH0
4MFKgyjE+nTqW/A49eKk0onKr9Dgp+KD3vb2Jf4E/34KPPSmQimu+Rn/w/Gd//W6
RJtAwzMiKjnu3DbvDmsbdj0Ljf3hIms0H01gsXkr95K9yuqm4hmDNgFSm2lQeWPW
1Fn1VWi7t/o2Fe9hrrDLk013QoCJBkuLAaDbMvPWKG4VvKrqcTvPP7S9SdSYfluT
aeTle5U7VMENsAtYObQBOnOkm9e1FydPSRmY/ATggKA/7N6FYq6TNMcrKysTtMiu
tcssE5nSVDoqviEFTh4ITIpb8TgYOA/QGNwyS4bA4tv65eGD8Xbnib3n0jscKjT5
+aUT/gI/rxP/RPYAcPe7rSplbMYWLqCJbg7iU3g+2X4CrQkfCwteytxxMmpgRJaF
xEzRHlz67Jvm8buxFY0pll8+P50UomtFLBBY7glsERKLoJzl6UpRi7aSOuVGwarC
1182Ohf4DO+QtzplQzFru/zMXEnoNUwQ2z3mJz+BsQbsIoOh0zoweuKHILk2qRU3
GKIwv8nemGUYGBmTKD8Ciw2LDQUOWCpjZQwF7eQLFQ/lPehc+DIGSLawA+3drJHM
QrAdLDx4E7YcTay+4lg6Lzlr+JKLOWqtu6l6IqksG0DvQRrtiu/+WrpdWL8HtzOb
AH2oAouSplElVffGlaUdmGGx8VWMKrRGfTImT+dDlH6xgcmXff/K+Qg/wZC90QNO
9cb26WlIZTnOhLmlj3ZP50zdhXdqAbOy+1M4W3Cl0BpdNm7DXgubKf7d58OfJkH1
58sreb+/76Dh/l030L2eNNmurFt4LQPspBaXJmDPgDrY8xTH6sgIJQG5SSj20341
i0wcHRXEN+f/J++2BrHcTDkjd3PTCd6nBM/dNgRFB4HnF1Z77VBMpjMYYX1SajjI
Ofpre1l51wZMCOgCxZxKkduWv/nW5InaHlFeZBhktskdMy8cdX8/TEQO6HodrtHn
KXcG3GvqV13rZPi646S6lGnsE6nP/E+hT4kC7jfrxfcEB6ASp9/rGa4n8mWb/KgQ
HN+AADphrN6mBojePOaKBF2LLMIrnlMkZBjU+DHGLus7SgR76j1dx80s3u3WeZIU
t1JXH8lz5kvQy/T3CDCYqcK9YmDQwBtNsbGs3/SdVO5+emiqBe+pGZE2biXrHIAS
jAqOctn1joV6BAI3j1j3ZLZnhIbI9DQ9397JQVprmoY1DV1to/7WXtTsCtmMAFqB
wI5R46SPXS4QWiBUEv8NZgybIGnmC4ZImrBMilAY5HQ/MVA28Jt8pskV53f85I9P
M+cqAT23kwoePlU9IT9diz3VQuJkVtkz8LA6mXs93xmwEydgxk/vJi2W6Q3F+s01
PwpctHRhivt8DVhU9Pm3ISSro163oZwSD3NZ90SpcrbxtPhApcaNwZ3NSImuZ47x
pyBNSdnTnFcJkcZyIBMhxa8XKRwOeZTN9tGWKKo35BivDWLqS2tGdiGbUZMRU0wh
/4Yipq1yWg8fnLFsP2MYaf0YfThvSGJiLNj3Ccgm1Xjm42PGPOkRnZPWMk/9SFzR
pRHcKJkbpVmBJ9gum/TeiYB7vXRLNQkXcNAygptG6A1cNu18Nh9+uGafm9wJTjBS
omm8mKGTOjGZx6eRXroaXQ0H1ohYtaKW2z6z3+yQagD6YVhi4S6Kbkave+LofhCw
hlOTH7Ht8iXFd92cBeVyD7MWSCQuMM0Xsi5yPgIFHizN+L3p3C7YdV1f1OtI43Ij
wjjHUcEhSFPj6NK57vDjLi5z1+0J/V/6UBZf91bhTfmVXUoBFZJthcOOGnDrvVHU
WIYfXp1hCd2Gq9OXL1QLPZi0/oBSyBh8gp3jVB4p7kKDp/7LZeCpFumIYwqdBQbH
qX6Qa6RiD+iOO7xoV+BIsmMgc8ilLiLQdAWWldzMG6fCuJcqf92ohWlJic9VOz9j
rBCBYdoyZEmzuDQ2Vobkpn6XfMBHsgERgiv34s79JXOA8ntnA9Ew+Az1r+aeSw3y
puoyFnrxY8GiTWr5qs3rCsvkbNoKiw8Ug9D5qeuVx0hk/a9VX/QjKoJ5RQG94hY5
PUTJCt0QgXuuPaEiT2LoKKATOIXy35iKAc47jkLdCxAmz1v+8yaAcjLjKMqu2ZaS
xhycpzc8U98EUJOmdQ2RuYMX75FeQjlTBSIIEsjadKz7pqqZ5FsdMMkK3yyi4bGG
SLVCR6Up8iHzEqyOGUEKeOJmonHoF76b8KXyGXEyJExfXKDnbdW0NNclaMdH0/lG
c/rQrsk5gLZ9Givmm7SclzcasU9AcjQ7ReuEknZhq2Qt6CxYaxY/uPpx790loRaw
gkeau26eY6r8gqz2FPuqCxrd75T4VUVTDtP64tgoNixpgKeyia7DuX85O64NTADw
ojOZSDuM+vUqtv0Sf5GJY4ClwZVYvoWOxrmnnD7a9pqylE5PaRFnrKuDwuZEgGRV
WW2GIeehlLuISnFbx/fuUzbxYt/SR/8whjjau89RYdzNuMEXR7Zm3LgRqSBa93DI
6vE5/KMVkJtopL9xyvc/bYOIhbTMd4EnQz/399rXK7b9FvMDNluMLRk6kzOL2hwS
LbkLH+GXYd8yEd5MRvNJ9fWHe5H60Kz/ptZ6uidka8zLWYJldMG47Knwnu3DVuJD
cMoMrgrTeBGd/8b15qOpMAH09uFJhnSy9JkeVIJxPc2hyEENQui4Zo6ATCNnD3tO
nZBEMIlqeWXYgZ9QewORn0qlOtpGKlisD49UH3NPB50rjSdCr1jPCrsugdSUlbu8
djj5VJpPqYrCsEZZ4xDt/NFqpf+2yVQl0A6vtQ7q1MO5ODFo10YLrROzClyxXSaD
+gJGJ65voBNij4GAcOYBE6+N2p1yTZUu8eNufJxl1TWxFCN8AMDUwzIxlMQVN7U8
qyxEzRk4KyS5eDvPqPyjT1leV8/IasMQ41PcR8f4jpOO/v1MUDHbUeXmD+5ZlGlT
bqTxoUzcMcor4uEoK+9Hzkz+tSNdTD+TX1NZ/wGpROSVy0AchTEse8rN4D1/Rg9Q
xQPv24iAKxOvaP1gXD1BaX3c6PP1qUacYFHoV/DeHQbQuTf4RSSjv2N7Yo6xO0RL
gmF6ABo/mSLga4wyx3mq2J178x1HwGvNw1hTNjrLFRKCD1mwViYoVKe4c/d3xsED
H7nUH4p8kPLHlTTOUHsED975koUTmmZZOIicT43ONyVA/6M9Zk5bupgIKx3nxPp2
st/OjoyMcNNBhIBt+FAtsReT5RXBTM+O2prbmOzr+hbpU1xrO3vO0YHSjaPSje0/
cqhO/L3BuPUjRNrjzZAGuL3kCzzrbUPH5B4pWwH+439bT+JyfvyVKGBLjHC3iDff
/bDMyl+YZS0eddhk87c4aEacUHc0aiZEM50bsV0jdXCyS2fahjii4zxt2TYCNTyN
HZO7n2IG7CugHjT0lejyvnP5TuVHi4/iFdIoStIgVHCpPAd8nSTByawiYP72z3fH
l3zgCgC+V9KwWq3oOx88/mn8An0qP7txB1yF880tfE0ede0Ij8HLD/lZPZ97AFUj
mTiZ/mN5Qyv9h8dgWXjy5Aet6eBEuyCcDzzTc9XTghIxyDGx9aS8kkfndw4d3Geb
xDuBRFlNvQKFhExqycHpnCoV+waSZvHJOxLVC78JHQT/MxWbs3vNlbvSHU0t3f0x
5nLtSdZrQ7QfpFs2ZhpUGKrjCcgjxWtRpV5bxFkxpcghdkF6QyH9ZveeGg/EgZac
teymy5z39OSWtxTLV5RUKZCtsWwg0EywW0l8YcpXVdzm8dzu2uk/d4lqWmN4DNuD
o9ZE2zxRj7lgP74Qlhd/NS2/5aOq2OBNsSaBf5kKpBxHnP9OgsSyeJu/KqVgbdOw
rPGCjyQhxC11PYS4bDHAoyuDid8MeLMfz/Nu2DBGpxxYxsNsWfnr5SJjhx2O/khu
lYxyQgqGtQ41LA5Mq+rVhXRIBw3fcLv32wJJV72DOQaSjp8vU5+jCPIqEy4UH4LS
p8gUc3pjZX8JMolJLwpxQHxzaXQn8aLvbFtITDB/1QlCf6LwytlKafdXoHKAPkOC
lGypZgDnlowi9pDCmNCUQy0SqUusDBS/sHhrQmeubCwPTaTmrn1iKVaZayx3ZHWM
Ay5a/J9eLnkRUPCp71Fk+F8TlbtCm714ir15MeyvMEITzNPPxEs+DuzHgwkfuZSV
VboEDfxOpbzd5PeELf9qYOtVrgDxMnr81tW5WUNBKV4ldUt1A06E3x6mFWxbwcrw
MafMscAxBacelcGwt9vCcyPBMWkMChgNjoS2GqpS4KeVyVmwaEBjB8PCOKRt7ALj
ayO4uKg1s8DVDfEIcT7N/iuMIjH5B7NuRFPNA18YqJyhM2LDRv/bi8xk2RSig4a2
+LBdQsI66XRgGsfYem+Cp6UEf5NBCA4W20Wmwc+x8CQGiHYpMpexChg06NfNlBEx
bZAwbcX1YYopHKuejOwd+NVImpuFtdQ/jWWxeykbMVYO3jjjAtMUb+BTM/521/Nr
8jNZuKOVR+EG6LWzv7iDxgmBCbMKQSs9yz2TZP1tApndftJj3f7HAIH3iBqOBe4M
ro6S4UT0oVOVqtSRRDAoPSClrvG27uXn/E09mi3r3ZEKbqlkZ9R9wR5rmQSt+bR7
AIGxoonsFxm94b+atBhK9UQtBRMMCmHVE3minpA8arYDxuWft1sVKoPFWbF2DkKk
V3uDTzFOdGnd6YkXgXRS1kE6zXpAx+0OH/m9LV5m9Qh5HJ5Z9LPCOg5wdcstJm42
NzWbTno3t5onaKVhbH6A9YZB+C+7alSKEWg7Nj6DeApbYwf7le77aeBf6ofOFJlW
pcLNFZgkR4WEZd76J6GuWdUSsnWMIvMQNzNF8bstbOF69DYg6KoH7Zr+JlA6bDnI
OC2rG5HZrQxTc9m1RPogbK3Rk+JnYx4Tudy4x5Rx2v5L2LA4mFLubfIS9PTTGs3P
kkj2/qJ2NYkw4p3iTKi2VcoC+HsxNdWxG1hKDh34HT8fV6xmUdDd9PD19xRt9Uq+
erj+jwsHPabEw93X3g3WrY6KNsmmZmbzTHUiD3tn/d9dsav3sEDBbFsGO7rBbcKp
7oTwOQrAApbHpPKcB0/PLcf/sK3RutFv5UL/0/3MqwiY1h2z5VIpfy+QE5UCE3o+
oLx250au+I8o8EGA7zzwtgViDoMoKH4z4cisDlmoryuqSilr41rgRrfDDta/Zp/Q
M2JyCdw95XAkrEU/8XQLfgUzA+RnYEuNsLFTbGz11Jq+dHr7kgXCQdc/oM5FdNmv
GBDaACslmSyPM8WDautYP2wCSugNGbF22y15/4D5/8zfIOo6d5+nYCMKoxrOsvG4
n+GTb3aZkKPwxcwucqHON+0s+CR9ThrnXjpnMHwI9fRAy5R87RdwmUTHvLFjyo+a
LgfN7N6VkcLyJtjXQEvo+WRhlZNRExvtboyWEdiyOjwH+gxwjNZPGhl0EjhQEaJs
65FhFZox03FqS0/GyoF9K2a1cb++M4+qeArrBFEKLzZBQzlHwDQMcbRPt/ZP+pHE
FEA7rGmOIMj3M4T0dAXNYaJzRn3WiahIvHrQ/F0zfgizaY2xOCI1BuojCINE3jDA
/JlLmFytAwD12FTPeL9A3aPsAKwnZw42iJqrrcPUZ0UoI5EVVlK5W31IOe3Nm0cG
T8RDH4Y7hzbNHR5Ac85OI7oT7kq1fBMXDFd2T0XZceRgBFqyRj9ks4MJHUSg04dI
3LmHj7FD7Ci4iG7IfS2SLR8tlS+kIGRbuEBCItddouE6JBk0MyQes935bHiAaqBj
gBzGqOvhBIoqe8dbQH4YSmkXialK/qdAUW5wBJs3Kaz0efJFSq4ggfq9UTO2CmnG
+F4vFu2xfgDSfxd67nkncsvIYP/4kSQFME5lBap+QZzzGt2DX40IUwGLLwAQ9mC3
xmLnkiYluZmXtkzg5b5bl6L8VxGLf5lL9UOJtwdc0bTHns+gRGOvRQ/0uXbGesLY
MTLMFgDNFhFfUB4mftwA5N7bGqeQosLw/2yQTP/Y8Mpn1ZXw8ti5A8+b/DNTZR2k
L2JFUhKPcEzj7tlK7HSF1A0bvz313zRGty8kWBwQ3KTPMFHGNxOoVPfEYjyueA+Y
ya3qaez3QtPyKf6cmc936kwEGI6llncUGEqh9bg96cmLll3Blv1qBruJySAV2YiF
GXg5nSdxn4Vu90vPGWgq6VwlJu7jo9Yvm8i/YNrk6zPa4aiKe9cV6NDfVPpeViRX
enLffJ2ewlFGXmvsJAlURvxEiqdx6Fjl6QA02QMwtnCtVX5qGQsNrfgb3JOLv+8v
RKVFNVqVSssyRQkgtSqiSrgQtevrvTgP1Qf4fO0M/Bcr5k0CiP+AC98vsY2sllHS
+JXzkjvMBREP/PSb3VRTmTWajktLRCjGF0S9/YhyIcLi0EaJEaogu52adTeN1OWY
CzbbABm0ffbBtz6jWoir5DZLVHcz7oBrSC3ensgTkBrPhuKSkg28LmUYCLlOALfi
+f5e1pNoOJ1gBnVfHddJ9389Mhvwt1oAX3seA/5HsXAUu33941zz+3j26XTQu6oC
BKDdoL0KFTU0O9zzpJyEiN2Gxbxeu18u/BzUuEfvFUmTmFRTfrfHogrqvPH5X/oo
65iXYAylpZEONnwgrpCbuvZhDSQdT7ZsGYTQEVbSkS8DTnjudAeNh0oM9TR2irhb
O9dDdzJvZC0/JyOtghKYyzHv6nLlA7GXCz9fuCaOnEDsHh2gAk6N/hgraC7jKnEU
EcVUhh4wVz3vG6pwUdWvYngPiyRQgrD838H3yhT0a5VcQWA9lPeEPFkkYgg4SnV3
umJcWyyCrNvISWc94HKTiecvsFRESC5GHyYpZvtDVn04Xrtxj6EFcF4qMSFVF/c0
2y1j3W3H7bhDqmci+FKmywe2gvouf3s8UYYmtHH2A7O0RHEyhmlD676adUx7+MGZ
Kgpb3m7ZyGp8Qd6DduHuXt3aWUUUiYYiXkJ7EkQ+L+76rG2iRSWPNHC0p9Oa1a2J
srdONu9ewd768qPY5zL0R9kBLL4dldFyWtMtw+V5Fyr9JE7HpDwilEa2xmXHPsI8
j5JgodzPVEoiIDjmU+j1yrCPx56zGs4EZGPxVpHgk9h6PZFvYDUWQxeZ44L53+ze
7g1B9UIWYqHBIq64194DreKFfqGvPcGuF0QweYU4WjLc/8S0P5PkaO7LdvE21wdj
MNLRFhr7UgCKU3gwPA4sIjPfCfPT63RyIPuAuqWqhapQx7sJprLbKEagfqyZdPBD
n52A7s6kMo9mYz8qHoHdNZMeXab3yTFGZQv/DnlEFK/eI6mAqvI2rzXHIrJ+9xoY
bubZTw2uxfrxAattvo+/Fan8Bzsl0ZyigCpI/J1Y2xVqv6IGi0zxeSbsItsRfa8D
2BVYJqUvOaE9XJ04Q7Res9+7nxip5Q0xnWJ94NghYmwwGMmaZXMonrCCCDz4kzgz
B960xTPj0uQtrgL717dY0UnG90+40MQ+GPg9ZgTLx1Ix54o6rQnJqgtaQaKzBg9w
zfBgIwhXCRwh2Sij+W8XM3ulCRIxYmfG89Jz63yWYHkI6OsLuSJdhyM7lv/25QEM
0z0Gp4jQgItcoPiDv5v0jRbidkF0SF3CvAeQjcY0Fz8V7TtYBKdnCqRyE7ZpSGxi
SC1q1LbnlS5hFO+WjooxZajza0qVm2Ja7yFRNejuIBgdnPyb/oridDbCgAKed/BQ
OivTVAy7a1PsCpQbZfI7BPHotW+wlF4U6IHUfTO8Gn9PJ0Pew9tHPmog2Zn6O8pR
TcT7ZQuQWhBwf3j9xUQaFRFYh7vbPjcsDDQHTcCXUFN6OdAjtgfDvxMz6fUmkIfT
P5mo2I1M+VhJCn7qGCqa6m2QysAcjxtF7CJqVoaqKHT9rrgrQcUsR4VyVQMJxauX
7sc+nbsvtvcRX5XuwvRRKLNjzlk3R70zbZNCwIaYeJLu4GwNEVieikTFlmV/5ZO9
nz3+OKngyasekPKZbAADsZGwC79pTlQXWLAphjqefRJExc1IJzKNtBNd3DKgBVcJ
udZ2kWom0fhWAlFgOriLvTEfjwB/uYcgGp8S9wLxD7aOlVH6Nk/HLh0eJ7jFGxhf
pJxzYKG4aPuLww5F+WrUCf9im2GBbxOxCQ/A4Ppy4fg+TG6yuN+xttHfpxlulJ/h
pnXRzwWlM5g8HFgkFxy35k8aVlka6HPqxIMkkpcuUXrRlDLkVKoMm/YCSjhPfiWN
sEV0RaR105gh130CMS9yvDGRFU1Kr6OGjh0pKPqA806YirIj2azUzY6BjT2LkIFu
M/0JBsYq7LuXSgYEH76m1VWJjtrj0v2+xWDXDULm7iWOWN0Q1MaMyAGfTvFl91YQ
R4b6z2suTqWFNThYKJISGuKvIEUwvuLcqfNBinar+5uWf7NsDfBxZneJG/1jdVEp
8uJlmdWZPXU81VLWGHtYyGEZWSTgUEB9pjuwycNXibHPmGU45dXNxXg7/R5JSIes
XShtxSIsHpOhnFAe+C1GZIaRe0S7JG5o723ds6wCD++KzGoWwR1AqtT8vHNyFs1W
PanmXPrB3chEOwft9nw5tstz+8G1ikBh2YGk/7GykKSgPIgIpFG60YQ2t1o6OjnO
iKuGBd39nF8fCBs0NwOSMdUCiARjRjPi9qw2lQsGI5/qDpnBFbeUx32oJNP6uQB6
WgpPrtoLi+5cAyMpD+knNjLA+w6byxFkkswx8Q2N6segMLRYZQoguJ2ZdIEipx0Y
qZjR+4jYzhEQ1MEVtDhkNlEpc/DFh2UL2dv1yOESHpoYQvNKQRU5xZqafY/m2r3I
O8bkFIFvXwpXEhcRTWEr5Ik/dMyw5Vzorx3oZBZ+Ka4GTJbSYReNha7qSt9VWR7T
/SXBZCYGIpO98I17YMGFrD52mgOumK0L2F6Fm82BovK2o1Qon5Gl/Eia76y42yl2
zf2Qmd2D8Sf9qR3vpcpQuhOyMgaUR2nZDYt4ZzjbRo+OsdfZPcblWv+sYd7mZ5mP
KW3OaiRaUFFonWtTDXKj2/lkXDbVipGhbxZH1TDCElPh0u2pRPC/NAIxc5GJ+PMo
YwH0yHA71iBShsOIzEbe2lbQTEh8QapLd5Bw6VUobYTB/AiuAcQYDEMH4tlD2WT3
nYHQKYO8XM8pAJ9xRmlG76WPXE1F73DEfBtyF30pZU7kFyAE2ccFRp1a2EdiIZ8K
LzEMlrBChTuUVo18lY6E2lXqm4ltJPNepMMXTvZvbRa6BsHk4IPtFrPWIYN9HUWR
OaqDMkrF/6x2sSiAzSQ8csSAtHJCFez6Ck3X10+ofFSb7f5ty+coydQyeglIcnKW
9OfT8CcsRB4yN1sFhhR/fKZlYfSyCwlZQcaLGrz09B2J+otCHcgz81EPxX+UtjfL
Qao8J07abOBpgyR3QoBBKPjburKlC2I9WyPmr48o23OT/BRiKPWIxaOr1vwYi3Bi
tzojdNA2uOTkZDE8CeerBy3QSCZsNQybz7VQH6KvgbBFrreXa5MZe32eP77E0gnZ
RyoOnJKTsLTrfNDX//7VKhyVrDV1RmriGq8HPMd39xGWaehER7hS8XEGeGjoLwpH
y0rSbhZNMIP9GBIyem4+GrE3jgUipeYxs1F5+jPdXOk2zADg8jIJRH+IlcVvFVtX
NIUb84oaLzyDOcS0hzjK+SVCX+aHJB3LuwrxJuVG/Yql+ZdBiPPgZNnnQdwji2yi
AzGk2DObZbOZ/2gZVyNFZt3hYxy4WE/u5SqT61NWNg53TZ1GjLspGTKlrAEuC2AE
1DN2A/rogDblubX+uRstirAkQqpFQygaU/XKySQwlljCUeO4vhS/4CoCElfaSzrw
xx53t2HID3daSQpZwt5T2JC3YNTUA4VvvaBtOH13EPGiRGLl4DjTa8cn/PTNeWVN
QZFV/hYZdu+V4Ic9GLljUTjfYvfFYkp8WFKEzwAZ8OeTVAt5Vhb8eSUYuCYr8cDR
B4rzwUn0LbyjpTfNlJn5d4ZTF2i6NsdS/Fz9Z5xjZBcJy3I0cyHRB4urZLu6kZ8j
QQ0I6xLDzJdMexzz7TwYQnu9DJZN4Vgjg6VewPbYPckDWWSbS0Yk9Fl8zVep9nC6
02AeVfCAwWBAnmf1ZQ00j3n4ejMFIgJ/WZf78k+Gwc9W/eWPuyXSLT4tf/YD+WxI
WDNV76r7TUZpoSs4lQMmJN89t23Vk2PDlfGK1kUvD1KDuXBNKqNZgd66ja5WVD95
zuWohqFuDCb3X1KSCiI0Pw5FXqDCLpY+bN3tO/3D0ijtHNEYhwsoyt6NwBoZ76HP
qV/FEgJ4pYkBnw77eHXaUyx/JBRa+eE239thJQaSbvsKZTgel6fM9cJU6miy0jw9
KFHAXS2FAVtJZHDxI9GPuNrLaaS7lg8kryQ8HRWSCDiboaXeOL64H72SAklJ+bSN
xlWz0y4LEW3n8HJ+Wy5hxAlrB3X1E0NjbbyiJD0tDCkDJ451F1ukkMQw8r57UjZ0
FC4K1HggJj0TGoNujvVwqZEOFSe5ow+6Fg6jEeZvKBRlTRXxa3guEXp07uoOhhX4
yKX8H5O1aBwKJSgYD04ATlPS7fA5YOQAu6aTUipLyxy/+vRx2uAmHwyLg+2shCEo
/CFVWsUX5Ym7sgSXt0oGnBhtCuyaAMwRZPFSl/B1k6ZVe2Ei6P1vGwZMWJwMyPP2
txF6NKSa7Tk/rnCBbwc/ib7xG1vvqwkFPw/jxlD4wjcBL8FrwYFtwYfoATUyiztF
B3AVntwkm1/QiZI2QX9YKwoh3TkkzBZmsaE18jXsMmtFH0p5sJicQtEEg10qhYiQ
9wEYpkbjVPKDJVt4sb94clBpUfUSRa7JMwdJgzbyCONmO3Weae88NWF5OmB1d9TE
vQUSXY2WypfD3lfUyVSStll/HzuiDm6Dc2JVJtcRFWpOZMJERE+JxkHzWXjxnDtY
H4FH2LHNTlQnOEPye9GA/KmcZpzq2PHaPwTbWxaq3RAHmxb5ZjV8FyXtD53H0vln
iW9ZdR1P+ZRO+QMdairvLdmjYxjO6gAnWKCpcyq/QUOGEz0eigeV7zUWdmSI/LwM
QbuHWudyd53Z+SLVuXM9XEqX+p6V30VrYcD3ACQLhey4VNJMc9RTr2Hu3/wxwPVi
6p0S4btKE1USgOwtQ86D06Ic04Fmd5EQ3CNTnk5lUBxxcXcjtoP8DqOkCrHWDWKC
eyAUFSwlWCMx41I/8UCr/ulkjVCNOa8jNgSt3xSU8PFbSKvXyCEUHcVONYTz+h35
tRUtQR0bWGJofX5gwmDm8GApI0gXfexqI0VS10KEeQyEO9x6I8DcmdwGsyKbJzRZ
AorHzrflPSC+3hR1axtMv9vd8iSBIPBOYdvktvsR4o19TK2Lcl3Zu6192i5M2QL+
ZT0zhoqLRP5WleorzDv829Z1jesh4WTJHzLaViOmweQFknWfk1E/TFywQO+suq5G
g2sA6ojxxMMPUVvBhsiFzEE9/m98l0Rcv8t3ioVcNSAgczJcNd6EOCea+ZZkj4ZG
HwqUH/jCVqyWjfpEa4NhptutEkXWSq+wCWmPmKhNg1Wr+FTjjGj55xOUGDRBMH1h
S/1CWlmjaBbR0QWbqidJMcoPK16Q6C57ivPj5Vb09oIFrZtCk6DKt5sIHY7X8yY5
VninRqGMoRnJQSOEpPga0T2Gz2lj3mq5GAzjBQEY2U84ZAtNn4jYU/rJv1UmTmy0
TyvxR9gB9DHe+9tMNRkKH1IO9SUgIIrMy1SebFOFiIFkT0PBRUMFtsIm3rFh0Abu
CZIyzeHycVCjODRXGuT6DT3BdHjCJAM89yEiq2tXpLeqVgyYethWywBI0gJpG0d8
F3w4xA4iDJlIxTrziUPNatHOjvtfwqikLIzwUNxY4usqKwNxPMyWJi1uEEuTcs2z
+arQ5kmpgOCeLf1gHmpRMD+pW4Tn+KcsfuxRcbzAQDcn0/KoBf/vdkb53TYARGzO
Gy8Qsw7w6CHRktAn0R2Tsnfbg3rxtb3sDiIUznLrBjjiPc5b9kHUFZv3d1AV4pzB
Xb3IYd4AiGq0eQIU6cmzuY/emwMzJSakplzNYcm73Mcmmg498GUKaBPfdoV6vWWz
ztoHswJuYjVv5yrJWEFwt6RsBUL43GETgpexDQ43tONlHMfsA5Xa4ZfB6q6ppgaS
0RbWC9kvebBYlD3dTzB8G2C9N35g6katAiksyRjbPL1Ck9ey6hhlZpqTQJ8BaiCY
0V7wkj5vnGaKZUpinBuakPzKK1cSkpCc9VbJjyNw/yWCN9aGJv39pcVdDz3xX0r2
Jbn0g57EtngascHnje/rVovrIKyM8G88mk3lb1TyTf/dfAK4EqyxXdm+m82wNezH
YUOp5JtbQ7GcPqTrrNv1vfOTymToAjz8znTduBH7Q1YItUzoGOFE1X18Bx1s84zT
4NlQ6s5aFephDHehNMLUb3zN85lu60tgmyu3UYH/vBcC2UPsAd5Rx6KWCWyLNjIk
EP1N9ubBp9G31Xb1mTWTUVgE5+vIyZ4nUggmlXiEuw81BJYRkJ/EnLcmP3w8kDXd
bq1+JwbvbFtnyaJ55YpA8qsXielxlhtq22y6IL7quI4AGvp6KSJo0A5xu5IJGKWd
k+hi9MwIaZ+0MIlLJwN34obkAOZ2wFXeoL8eP2Vn2GsVgTjsvtNvOmt5D+KgI7s4
QAGTnAOn6SPKjN8XHIPqVl80Ude99of1qYCFDlCPLhw9uASEVWVj5T+uWhjc24Rp
ATPXF3uik9UMXTjAp3WTOdRe3dKzKUdD9uqcKegbCJpdo/XYwrxIvNsa7qOgsLQN
YgBToJK52Z4+MmjWdDF8mXfIfk172mtJBfGzI+YeXzay5BqdPKGpI6310ML4PnqU
VqfAqmIhEM2pdmRb241BwqZusFW/nN38YT6Kxty9JxUtjxqVR0HR3EdjJDq7cmFo
GcSrUU3stkJodcgKbtszl3qATwQBB2jRiBr9qELnt9LVfndEI3QpavcxGX+VPSg4
jrGQnNNzwTniBJq5YItwIBf6RFF2JG4Bi0mNd3xrpkvdkduWtZJBkt0OtX3HJv6Y
JVy6WCDOKfFGhH/cDMxlWHfrV9b7MVyDBvqxsDbpwKesD07sIos27BrOs6nMwwKz
DL+oRh2Ka3DxWDeJGRNuasnRVDpwEZotn/NfIygAYpC1vQwWym7A4Nq3qUt/1v4/
JawbBg7jXVtudcqVqI/dHJOZbwo0OpvysYiwVeJpdtVaHmXF+IaFynxWqL6aDiiz
eq6865pJz+eg+i13Q+2Q4vsnVN2w+3YfHs+WoWezj/vzqV+qMp3yDdCC/rS+oYoQ
ioHuMg/aDYfQ/hN32ZxqYrAABJQAv6Qv9uHTNcpfbWsQfZWgpNyjQj46S7O1HCzF
cbnQws8PqgOLPGcilf8r+tKBQbZyVUvXAcf6T7Aj8I3yr9X2rY2At0K9gTn9AqKW
qYyValco86sg380RiKoClJVBnYZCver52elTxA5xWZhEvo6ZylkAomTkfD7eDB50
L9T5zlEedAXs1L9NsC+diXXQbR4fD7fFC3VXMoFuTtJdtASFDvEMXBnrFfiM+ONt
1pR+wj791Ad1/IU4qn6ObGtRiFFukbcoCEHB+Exy6LFo8s84MVRVCyzg7xPnK6nE
e51Iqa45UTGhCPbya6iqYDSqYKoK6+emkphZEYZlOkRMnKdBLaUyAT8fXBHLTJWr
UjQC898mIP3mGq+As9YLPSf/l7eXy6SozypPo2nwlIYJRHo/exgbIJwqW7f4H3fM
vBR3JvuoYASl9eJXbykX1XZiwsherWumFAaAZMC8kfVEMzneCLpC6V9yXZqxbo/s
Y3AOC3YZcz7RBR0tBBpeznHTIxhbfWT0wm5tyd+HilE+8FGogYtiUoiUlsUVOjQh
VUVxOojsR6T21T2SYSKSYNMeWtB8GNDZhPdjqM1XEHTg3zhERSQuq/+OX9azlQQK
pCH92wXzEkk1ZQC6FHiaIiopOYnLO1VRdNJPyEAeGW2L5b8tugYZVTwz9GO4d5iJ
jYv/TudVuG6DugkeItCjQQ+nwtONpEkVXWvfr5+rPLcuV+mCZOQOwBMf86diKgMv
w06SMRb86b+hhDwEJVs0uyQRNHugv5c3EN9wQMRGxk/VL3L4jTisWykGdHyPuZOI
HiBiRQ9qPIWQgZOD13skmbNesBgF+bNg44u310Nom/FWavgCrrqDdpY+GaByYSL1
scIOzSLKjuvrQLoJWclr6kkrwsmcdQGFJp5E14TrroMWymZkXQCXn8C4u0luyjTP
pK8DHoJIGp1scf5YqOsKUVb9DOq0Atd3om5AHef89JEfWYpnOMc3YeaHxnen/N9Z
d/zMw25OfozK/ZoZn64Kdhgi1xBM2L/gE3UJkfQy8zVk7EuUEG3m2d0S5VeWu/NH
yz4kIY9ob62ncHapb8UErqZ3LozTI7X16wb+AiAnDziJQ99dU4N9Pro0g94s5kMV
gSQ2bbmFUChPhedMwn51QysE0JX5ICTUQ2/6+18xWzIkBWQvDt/1pT880P1hchKO
bxLxdIKwMBUm28LcwCNpXS8+pbtJ3xGmlXLMEqU+OOLYtcmZ7GsrjKRrXDaotJap
Y1UlFcSQJppaea1E2SHnDqY50iFypOHSpvbeIu5dcCBDRdQIomkC8lCwKhzHzC/f
duS0HB2WiYvS4Toy6vW/7fZSn2U7tZoz9gHDAoZmr9gXSEqf835ccMRigkp+fFi+
rxXG+5Df7pUyaFg2kpUY9aXFiFpQrc0uAvVJDQcF6MVXpdN6T/DDmeKgToz9S/XR
FROBgoJbGCiKNtaEPo6E1EVxE23s9xHMtIKq92vT3tLR7EKH0wC+HfgwK92xdY4Q
XWPeay3Wk54FJ/j+Vk/h9Y21HCny1auOuaHnqz2Od2oXxI1C/ywoJBXzJgN7QIeD
UzQ2DfgA63qID2TEgeTDhhT9GhOd2oPEIKERXpRBDDxBDEo7JddWO9ED95xgkBH5
sMMGjV4khHkrTL3wcDzEs6TbCk3llflctiRALcnvuwThxPyZTC2+r3rIJyOyc/p8
4xUiR2FWSxmNvE3Lg5wXaP00L8AFLxnqFgClUqcQIEjP+hVUQIauD+KhcA++zpA2
FJlPXa7cwJyUM9MzbI09iPfUt6I3an9+tSFnh8+4vfeyVL0DnATwcpawkiKLpQBi
yxqSSbvNhi1x900ZbU+E+R4wgCwbiXkOFydDE3172wpukD7f3Ri5k8tGk/wSMMOs
yga/TmcMO0+NerslkT6JGfLJtWKrQfq49tGr/RA2v3PCg2FrNHM9aBjpsF1YZXTS
evpyWi1iZ5+9Ysk3HvhfpGpIEXy89A7TCbtYxZpeCNHCWRbKYHIAeBgYz9/XQfF6
8SCuR4VU8Li1e0M19jb1Ll9r9ls4wJF8ztM9FxgqLGQXTK4giuZsps5VG4dhwfoO
fJtH5vcYKRgYv++LagVtx02Gt6FB1VNGWfbLITT6BwqeFDP0SWm0pYf3VFP2zOx2
jZMsahqN3+WxIMWxyh9Rf0LeHJif4AYvYIs/wjTMTgEQRRNbDd7tzzw3q9Fzb/F5
+n+h5wbHKjNNoc8nHUSwYhFbKvLBy2DbQ7FU7bdOE3h9N8Te8FaD9sv9G1PC+h2j
SvBzbj2l3DLtrtcvU3DZxb3az1+s4G6JdnbilzEcrPZVtyo1SpBHWD93p9ergXhs
7+wtUA48LVeqhE7a4rg/oLIhlEeBuKRjLNfS+cDeBNJkF4+BxR7p122qU/hxNn9S
lU+lzqcm4YvpEG/DvZTHBkuWgPd1N5rREdXnU8F64BDzfeEZ8TSUFkNj6omUnqGI
+1FOyHrm5CcjrXj0YbcXFW7xupmoH2HMOj+njxjtr8Qfs3x5+fMptf/UcLCv9Y3A
cbk1W1QLjBcSDZCfezBVpUxEQJG/oUfq6+aM1H4SJuNjyQ3pSzwFuqdfBAuHwH9b
CXPNeEnOUAax06p16xCPSCy8XYO/JoXW/Q63JNLgwM9+flBL42SkGbvaJ/56zqXB
zaa/xjxgzNzXCbip9eFtrYkRoaJkCk4E3oGwK1ZAtT9oN2r9a5LAQyMB6s/ajQ8Y
SOjaMPlPzH4DZY9duFrENJ+W/tD7yaZDMndMMVG4g0/NGojGPaXoD9IG/569k8tI
MTss0xmPYvRnfszIDZtrKdfCmrd0/vu9DJ/TFcBKI04PeLtDEQGQvgFOcnZJIDM0
7I+vSFyuwgo0SwW4e2mVyVgSNw5dVTjUZbEHbvOnA6rjdi7qT5yoa4xynNbPMwEz
4lvnP9iFa8JENEQJYjPcWEJkM+rNe7zWd5PBC59/C8hMJxqDsORPhjoQJtomFc5r
ZF/J/DpI9rCQvrWAcu0p/AzhVUorP9ympNQTroASUiQZCeXKKXCWbBls78a5i885
1hJGhZoSjYolLMizs1DQhUUeOnuCW4MqrhclQjXcSzRkISPL2Ey3uogaLP0avhE/
AXYmX/HQ8YeDo2j0GJKQy28rdFrcrqadW8BgCSbGGvkfKrRfpk4VWHXaMIL6dZ9R
fnz7qw8ptmnp6DctOPjRGiH+dCrslqsR0SuD0PPN0Ae4cxdNhaaxq9ius9OMKSK5
8aXC+qljQVDUlSrmjmcMGE4+VcekLggtGlQ4VnnPv4svCzoFeuELDszqZuhjlWng
q0gRtUJvOhadPi2Ytwwq5aAZUcWUjVYmn+bG1H3UVM1FCm4BhmYR3U1jcGpdy7q/
Z75QseSvDm392RS3TPx6zePsD38T7kkjyK7HggGo+7lB7BcM9qrggRr+QGH+/919
6Cr+Do3iMi3junTXH/HQeJvdyPkr/WM6mhkgQSu2fVCtrPNiXqhVR/4UBvZdy+oZ
M2itTbUgM5ZJNozLpWPngwFudnJXatr15Fcoc/hbJorPD21X1HcAVlzUiSERGABt
mxHNJMndXnpMgejrHy5+siFeRXMFRwzxq+WNrBuK2wQzTWdK0HMkh2fxXsYSqNIG
I6t9Gg7pxvfgZ2BrBkG6o2MI6kgglbE8h6L2f6PYJnS64rJS8/oKmMO3bmAnTnEE
XokDOq1HeJmqMTRZpPTQGijRAyYqipl5n34SS5TaxOz+3DgAqZVI5bbuK5s3CT37
/3Nly2ckI9nCS0ReNPMMTWZEhOj4BCOzc/H5+LnHSF95AHAjxage76hgDxqyk00W
RuEn1mqclGbIn3hbiN/t99qKEppFk0WgetK/Et+X2gPbkgweL3yfiJQ4a9okLjA5
OTo7CAGVgct3cSbJwlHalLsQR5cpY1vEXfQdshsnG6/kdMKhXVbMmjcSVk5WaA1V
1sdxfc2xE8URAIi1D8pWlLETgCnWpgqplqlUCqoOyHmF6FBrcIQJlrVOaOl73Aoz
TEm4Xs6eBtAJ8bXif/jy5DcO2PecX9DopcBh2fTOKntcHbEPQj2eN3x+tjn/fzSG
/adeT7WggQYjFrqeyVOlZxTicvB/2hAZy+DXZOfo6pLDuWCOEGlLvv2wS0XxR6et
g6w3K04RJ7KJaigquo0ZGkcLrNd8m2OR+/ROtfEe1MpA0yQrEmjBgMY+r5swFIMN
5MLf5NCP8C7xh8gbCjJBkNPX8rcau9uhkdlQz8W5BclZoedG7hD1rGiwZusFnYXO
XocHg3+aIcpnsAZoeRkQNojxwHTtueXcg9u/QnGjVStgxMR0DgDZkwDU40eAzOey
V/nMqlh1z2FkZu1nERf5121vvbn28TfkrErHFRGbE9W288jQcsgELQs5VuJD0NTt
aZFt6l79KqEv3HfQn9ow4s7aeEDA4CFI9wfuxluoacuSb9WTIkubbfPpX99+Cwi9
c1ZtWaXlyLT4Er5LuTVCrc6a7YLEj5Dq74rC0FmlJr8AvPasiOepS7PNSzw3aKjw
NbyNbjx8pT62bdzkaItjZzqpau2d0xJq4Fp45N4cS+Ozx9WkNEJNI2Q31+xT2hHy
wYbb0j1Je0ma/LuFlXGYLG8jBY4tP4ui34hHeI7kmXwmXdX1QKjwi0vEI3F3c71/
k5+0N+JZzThKMhiXdiCBZEyDQHBWhSUmQtYj+EhjhMExedEu+HMNt9pz+dn6sLkC
WMxk6u9cO3RCJa0+2wH2CM9x5gSeEBa0xLa5Rma7EshgH/9iTfPaZJ+m/IBOAH1b
Zo26nqzW+M6t+uxbzPfUlJRRgymdtoXR/I2aC4EtfsULWWzdovo8exBZ5iVg7A6V
wOTq7z5OjfvVYDw3k+8MWwwu0XwwHlK8IvcJqLBqZeic9AyGt5DPsv3+6GbgbqE+
VhEJo8lQcVrAxU9P0GYgoS16TKnzvBmQUErDA1m9p6StyYsp/oqYhrM6gl5mwsT3
dQ4S7ya/EUQ+8+421Y31CFHvXQCsr73yVxdAbTKq7cpd/kRwkFelwiinui1cslY6
3RLbna05crM3xy7BPT5ccQ8c70GWnPwyPvNJW88M8gMaR5djiBBdwqf6kISddP2+
wIVTVSjFukxRcCpEG7EmnTmTPp8EGxM3MA+C+b3zo2jqwb0oRzN3ypbpqi/nXB/+
tahXfVm3KZI2vkC9tHfwwNcWdN9Z9tZAJHPTrNntFCvxJlhZTng+kHPYl5Ubxqo6
ljMhEYLSnJDWm8HfAVfXLkrdWRMiv3drJ2QD222POYgjja1b4FchDoV5QtWx6crK
+qTtTI1Yl4fv33Zm05FllASBpuf3Yl5FWbrkiCL/ISt5/1vHQDkHGIAVpB5Tmlrs
ZIAsGw4NVWLIbL1GaHcfVm5M4gJbUSI1iTMkfAU41B8/FUwlNECNXy1CBe7HAK+E
XzV7XnLzydhB3jLbit2jgK5e+OrU4MbI0kuZwpjzJusuPQVf5LXZUqxo1yaMCJWR
lOCwHUSHknEdJ8hD0Z4MyNoWuYLPT92Yc7F8gGqZkTo5ppqaQxX3cT6/xa/s8Zdh
yQ3aOOrUCJcvh6VKZlizUIArwbh72xzTaFfdRN8xOLHE/5YjRKkWIAwB8d18iH3G
QWBPwKKXyPn2+VAOE8BLErHLMqh485gH65HCQnMpMn1clxnZtobHb5+t9gIqF5C6
fBMVeNaDHhBE6VO81HCu2vgNmovb+STg/0zEcfHp2VgAY1aEs0TWQtOZor88fVPM
yu1X2+mBqjKmeN33paZakhlgW31mSxasqj3hMaFUBljgkNkueZKzc2h91jFAdTCI
b91Q8PXVe1+qjMEsqmF2jzxrJH2r1Pg08wqbJSVbc6uuuPN8PX1+t9o9/sNG6fbT
tZqSKzsOqOxY9KauWCsc8vmcqcVyogrI6oFv2lz7NBakX8n1UHd2+B0QobiqtyDl
b5Qh0wsbJeEW/KEY7V91SMpY5jA6PdBuVuBjWgPJR3Jm3HgLkHVp513hdKOhElqD
tzFIV5GXm2ekhENqy8kzy1/DNwrgOnU3luTCFrMv9WUZZGrR7TDcINwBprqIHTTn
MCKXDdRMIbg3WQhfpstoqb1nVedBgPOHzGENwsjNJ6j9HziAOO3GPmoY8OCdvdU3
ZpsuqdkXFNJBmw+8S1c7e6BT5HKtakfe4UuSCfWH6QlZI2SV4JpGNmeC5j3BAeNW
01Ifc5v9yXWgaaOLOXO0DM5CYtW1H0s43nVAkp4bjxTqHaZdjnOjfSBNLn5K3rXk
aEZDuLjP9zec6DYebxy0/KrmzKVDtnAjTpG2Xfl0LlpFNGyfNWp+arYOsTlqqK5j
blBL4J2inKNaFEX6k44AvSAyLwLINXGZy1Xw4itzKxJSe4PsENxjFaIccepXM/XD
Jnb4GtXByQafHjd/0OGHgYV2ct3CMZth08BwMrZuc1E16TC/6pw2ejo+xlf6cprq
8jHgdKdybQUsqJhHkrLl44LcuYyHGnDeo2SZV2jX0FFTf8UjY72L35i9hrJWMwyA
G44hIPJgQaW2qov/UqR2dL05KKSUg+0WY+lLvj5xJ1PCbQ8FIHtd7ICdHebKHr7l
NvRqmTiVFj58NjBDdahGF1udgIHirZkpk7oxZflbeFSE8ORSvmNfnxQvGXYIXvqU
doK4XTsK3Fk58oGd26eZ6FVavfGRUQZwjyffiJRkcXAhNEk0Cyy5uyNSCwvsQUu0
H6kUYH9BclBKjY/9GsdFkrNvS8WvYoyeWh3rXyYmbt1ewmKxhDfS+j8P1w+iYeOD
Joq2T9AUwAhaqmdOw+JRyXr4hJGXcK+x9I6cD6P4ndNd5OVI7kl0VjvxFwBSNqLg
8t83Lv398A/vH70nBo6aM/GfMXVAfnfBW/3VJoyYiFs+5zS9bOMKqO+Mrr8Q6grA
AaBtvBcwMk7UeCBCd0QnBRsfEy5zqsBNbKV8cZSR2vKWD1Knv18Xay9+KW2FLLxj
AsKuutqA2rn2QFr91n8Cd2dHwPdJhQanmjVZ3yf1zltzi6LPC78ZftSMcv3dIKt9
O/Y5GAMPPKGLV/5kECS/PRGyCDgIU9O19wEu5JZ2Qlz698q3JsXYdOg0J7f4NSiG
4GPThVuie9urthO0lkds3h9TI+P103leqWRfxaobP7MsZIRYNmXZh+m1iluTGAEc
ATzkFCoN4G24clB5grfUtOOwmliut1IPt59DRjM5VPYIkkGMoDDSrX/z0VxhRgPz
0m8F79jEtfv9TYigOakfALcArfeYzGMYPHuIjA/edO9k+V+wPn+qoNLars4PI9qX
C/cB1+q3Wtu2BkXxB1p2B8t+VJRB88GTCKPOHmBXYp+WxTLPDUCyxcVpjQPrkGhw
dMGL7Q3Uu8378Heyw90Rbk0unADsPMz93PJ3uaYswbAbsogW/sKa7a484Nnzoyfl
eWdmFprf5tG+qtuUDe8u9IUdzqJBvDjwIhA78ie0xO6VYTToW17+JV+xi3Tk00SS
0p8HYW36XQp2mKdL2RSqFpPrNU6FTn4W4JPUKGzz7saSt5GUJdl8MdI0r5P1kIcm
+wjugfjq6+KCaObac5OJZqusD/v6SG5VgMdpZ+C43P20t56f4SdZQtqkTb02s5Ne
1d6cdVz2kBOHmzXAr6CQgW/LKm1Zo1KKZ23KaGaEdK6L7n+SJFIkO11+nECazlW+
widxyke92Z/R+Pjis4DIZFepqo8SyM48EZrSLLTayXpvLTVZCVmtRpVttlBKCrnQ
4rxlYb+bu3Cnb71VUJgwAAy9F/MoUcQH+cgK09zreBIza5bHhT9QXNWJ3SS+lpbs
FgBUdPAzO0iu/YJm7wKzp1SjzecxClI24dxstI5DH8iPB6MM84r9oZxBqSApiJwy
8aE9FZf8IkdbiLr8cCRhQDHKFK3c5OsJ4T6/IMFKAUocQ8RgE/wquE5pOt4vAffn
AyXfPvS9E8z5ScRE4/9a2sSa3j/WtXqLUM4gaSkrm745pprKDn/pXT+Kt+y+aArn
bnxd1nmWaiYsWV/xH5LE7eOMj1Z971iwqb1OUpAu9HgHSXh00APKOqMOcks+KzcB
rnJS9WnBKatP59Ib4dIZVgD1ZjUtq9PyloGy6rni8P2AeMUZlcin+pyKzuBVJGdM
5sBdgRoI8lIZlj3p5+NNnH1a35cyzU6OO1hG2PdbffopqpE5FhDlC2DEL1JT2riK
3yxclwYUJ06jFzpK1lr1pJ+YRFiXnLcQbmwxVZm4ApOI8T8SvHN/L4ppUsk2Q9B4
E46n4dUmqG2HExsXdEspE52NBxNl4mScFw0R6WM9nl0TciI6ZZ92y/Y9eIpjuLLP
nTxir8YFISTiAnOFtGjCjYukV2JzookopgZEEwI35lyR6cIgBdaYT3ggoHEt0oOa
wetHf8Dnd5jPRE7D2GJ2+T0f1ekFXq1NCWAsosXum9B76kthUAn19MYPyUO+OHDJ
hE9sqVXsEq/6keHcJoXfp8Hw+I1xhSUzTSzhOAAHwn3YCgHDANwkHyN0lu7Or3rn
/LmQ4uD2VWaLHyviwKxAS/gCnknlXylrB+lSx3IUtxmG6BAsceiOPbKsZNOksVhU
kOkQELH5WTlgVRyeDfdIm0dZxA0S2SxMCF42jZhi9M5N56oc7V0ynjDRp543tsfr
HMZomyYd4nO0rTW6ic9p1Bmblbig0wCDIFKH0p7M23jRHlPOiwCutdFuEh1zOdiK
Wjq30LJLjztkg1PbbQ6QB6DqLiv/DPCcc5bDO9UQ69kRLgn5RTL3MVMTITbWDEjA
sCDINLejBJT6NTMUZKEM/qa1+rBtlP8ni3B1zu4uBTVGImlm4YVvLElUCXoFS4uR
0tz8FpAn2WSyE1ipynzQ2zHkwETo8oJtNb5gromFi47IbkFqmcE/oyUxNiO4QqS8
DzEzLuIvcKIKYnu/pyFcaFcUdpkjOcwj1VJdromyTfH4gwisjuCF8Qwdd40T1xsR
tRnxRWH62d3nJvI/0N+5lue846zTLPVRstlY57QNvrvo1D3xGI9ZmhzLHOnucjrh
KLmoEGKIPnT0+vkOH4D8bV5pZaXwRgQPcH6EtXhYwWYrNDEzPlMpGdPmwakwVYgQ
dDiOAnw3buFSmy5Y7Y+jnt27SaQifMG/zEHwWoW0Z2I3fYp0TvRqV6w+TYcLwhY2
pfLchUqFRV7uRgX9svOc+LdNDsJpI3RgjkkGfTzWbfiHgqor22BDryjRu7catXFC
cYhMrhF0jXzLSI6iAROGuE6RsLUtld2GO7j0kblMKZckceM98ACxXRylq0rIHdjM
muOIWybTJRhYpP3izUog9Y5yHEcSZbcqsu3BIFJhuGn9ROkIhiQ9MGY/g3TjHgpV
maY0eTHW7u89PH5opBmYY2P69eaP/Q1kMur/deJCmgS81M37UMpn6oUMEcsoIlu0
85wPupqdZbMP56knsPGLWEZdhCtLrOL3rvXs3SFzRB7sf8C1/mnqRLS3LgTz28E7
clgG0mEapYuF3EArT4dcSjzHVSFKkki00Kmp8KKMs+c5sWvQjilwRqYNYxg4O2Y6
YNVU4BPEkMU1bUAqI0+KYKWXG5IbhREHOlFieo2XpNFdAlzs/IliTTPiSPvif4vE
lT6ngbMnx+TclBSnin/pGFdFncPE97AWTCbDpkHXs1CEavY1bZe9cP3Ub92vY/Lo
m3Th7D/ZYyk/oPiKa8Tzp2ZB936ntfs63JDZKE23kgcX6jjXC5ZTSkUgHCRARl34
o2R+1GXUzsgLQrExC5/fW8Nxz5wPjnZ+VgKC4uYjRcaEXwm/0SEbEN/szWfIroGn
ZtYK3ZwjjN/PFr64ycxCt4q+72y2tTAEEg/Ss6aHyrY6Cw+W+/x9NkLjNSbCuJ4p
pxQySRADBhkkXpzIX8NQrkv3VzcjAzt3DQnh255JEESP6O7QdbPCjBLYgUnv/ols
GoTNalhF4CZUoBqEfgD3do6jDkDHFKxmq2RIR1Cn0nc4eh+O5Kl/ksb9P6t2f7+j
1duL7zOmrNoWFucN9g1gRJEpBeNCs4lsZzwjlwNua/pTS+RjxwYI/gt7I3fsI80a
QstzVXQKYzcKXlfWc4jt+YK73jp1/SAnac84/WM5iwSenwKEK0mPHZynxR0NGBKI
bH08aVwbkRD5HNcTSQ0jqRK/8+2t2B5HO50zEt49dgQc8PaeWaqeskVbogIxYpzN
WMF4O9OQZ7jgAbc58ERcEqEpUpglVyk6bYWPcWa/jatHjZv+yQPXF5QsKVnpWLcH
nw5u1j9FyJC4Ntm09k6B/lO0wGVBXus+8rqfTTMPLkbeURZ45fr7YALtwhXiUEGP
8804CVQw87HRkmEh4TsjINDSlxRoj1JqZr64AD5XDVXoUKmNBLa2s6+po6jEGotE
kblXzkiJrVi0D88ep4qi8txMYH4smBJK+eF1+sWsnl6xsPrNiY3XoUyIqRtWfC2U
zjg4iDpBrmwpWkNjwKu3dgMS4AEMwbD47F0QPu7zpLDKM1b1dTWvBGW5Vt3obA4J
VDrV+CEOK/b2ELpG6OOepaq9laBxsIcRws4phJZKwMqem0hQoMyt2Ez/Kz3uNcCM
vZD8r3LNZdZYA8pRxoAp5lmaNrggMdeUs0o29eC0ltf6lkdtM+OYp8neZiZukt7g
U0Ns6nX928dymDVfe8klRbfQIVOC4WrFv/UsVXL+ajy0D+tvVbjei2AsA6F7garj
Gry/qMf4F2IU/IOV/HNzAAuAo2271levxWeZ18X7oTrEX/xGgFb+qISi3VI46CGA
Q5x/Vl5o3HdBD8iRyFunQ2/hz6XPJKwcxKViXQZNYMYxODk3khc6obNaZlv5AuGt
+dNwG02ORjkRAW+bAnGOYWolPYuraaCruSKbDW5dozEHuBURTB5ZXLv8AWiKTO/P
hyvqiS9/E0BmBofOo8OiU0PBj1nvyDDBUJAAOSshofdExFquQY+P51VLXp+1SpaK
U07T2AzjpS/BVvpZfFFmGNtdfA10FRhD/eApgDvbDiq4CzPL0O/bYrEEw7bfd1B4
nu6OwO+JwP7yJXlAuXEJoCUzI6q6Ra9I7gHqAicvqY+h/TIm4xzBxzmteUiNb2+/
4G+yKGPnLAwxR8dXqV/Bnz5+sHPfIRcYKCTpTKhFv2MeDWu5UiSx7yNV0Dcrt2IH
JHmTuyYl390Fh66Ib9MYW7IlbyZTEkaxuuGLbMsJ73uL8J/70TvYcbVqHDkpp3TD
6hc40gP0tyz3E/xjFdu3yT4NqnqjRleNuHpaQ/uKCQmt1zHB3c/AgyOeKcFN9qU3
7+xcj+H5H9d1uYuPdgR7kKDRjOgK/psbPTSSGgigM/B0bQt7B4rnPoxFv6ok0AlE
9RO/djklEzsT0n0lUSpfkNDmlHlFk1CGoRkLVWbZhZg1zojA/UTJs0Kj727oCmK0
bp4qTRVvBDoxEZB/6SKgwM5/8SJq0nnnQV1CR4GqV8qtB2xN5SDAfqNT+w7R5mTd
PGCwzKRwcK9l+NT/MKfHcS5yhJgD3lhY30jzMXC2A+BwdoUaGXsbQqqWbeA2/jmE
bpNBB95JcqbVCYG2y2CejMnCyE6mS5jRZklGzKs84bfTYfwyQfpgMK5mtl+0t9C+
NEaGcf3eUnlk2bcOtQMll1+UQl/Bo00SAPPjS36arvkHW1FmaJEnRqcDL2TgScAR
uHQr6FYKCpPm/lOMtuI40YawinJwe7lkIfC3DQXOSDD/dYlhk7S0HSBzItGx6B6+
WpJJG3xQ2jCN9MOE7p86Dz+F/QFzqBfmVNkEH1B99n/wL2rCHtkec66ECJ6+O82V
1Wg8Symb3Notc9aimITGGIhYPFL09uqNNCS+ZHJSkkgMi3Hr5Uqn7yvsao+dEKDO
hKjj5IKNO/Q6Y3rbDE16rI7cTUI7AaZ/+9YudOB+dGCGg6R/rKTyVQLd4R+yur/q
R774CZotSBDeHWx27LQzRK9DZhnk3PVw+ylRVQtrmnh6TGBhTbSnjVco+gqzysGz
FoXfG/btnObRMY/03qaz3VPawmZ+TkArFCdwFZ3o5YeS0ttLLIfn/PlqfL7jS1cs
RdPnB2fR4aNhutHKIDWLsWl9uLIrbHR6F9HJgjpyUUYQ3Mp0sffiB+oXe/nZ0LOd
VpEZPXShYSYMtEOXYjohuF9eiWHdPZekgqo2c9eCNG+kMf4tXqlSMl3qlnsWwuvi
tzl4Ict6kqjmxSB8hcAOKcwHnzpZIiBWR+BTQLGodwhPr2szB60yPLR67RTvkEZW
q1KJmucMoaySHUkVcuBha262DavvLVtPUFJ5bhDPiZIyn2iMcFz2lXDFVb+G4ggN
gZNgaDl3kaymoqXBo6CIwBpBmaV0uo4YYGy5VxNFzihcPvo0Pgw3k9v2hV7X3IhU
RlAa0Z6tnYGKnGEA7azPgF9CqWaEfIZ+lbmYYz2TilEk3Z/bIJC3Ys7rh+CeXZpG
t6bYZs47MTcrzqvfnlbyyGoqaKjBX146T+/IZQWrAnyEI/BJeQHENjG10VlwG7WZ
vDCdR8kqOFz5jaJhgasee8+wyeL6NZwTgYGdDdUEyI4SkVQdyW8yx9AWpKmpCFM4
k9yN5weFsrFTulGX9w0jNjC9zfEP9iD0rQPfFRdc5j5GS9QOh3ojwIlVb7mQhmBD
8crE3v/ihckUXMHOTdZnuD5L0Vc8TLwce4AHejsJ4GkW8l3RO23nW8ealLeaEet+
Kao7PvHGTOhNm1n3A2MkLoFUohilY/72HCTasNMzW7UIi5belQTETdterf56+kzY
UPozNzkEambTisq4DMuJESdNt0qIR3oeJvFvbpiJP2NpqFOvW97t5ns7vYsgypOQ
urEOLcKiX5tLf0jekuGKfsCtOYqzaqQSk7FO+AGYsw8ON1B9sSk8vWb1etSvIljV
zm3ypZegz2J1KpLbRS7GYdeynn8I2Cm9dfXwd3XDR8/3YPNDkwruPh0wiwrqUQBz
n85+UIGurl3FeboSSgTS77ScGZ6Ggb5eFy53htegCuSmVe3CrVI/yPzNcEk+VtZq
QGl14v4E99yNzLOX18FgLCX8COVf4gIZHnuW1dFvC68y/NGFPVTsCOQ3ieq+DoVr
zIFExZd/2lshYYJ+fhGgcvJC24bCEN5xzeUiC5EiMkiL8Rfj45HQSK6mGFa7i5fD
RJZDMpynoTOUqezXeVcn9DrmRilycDJ73Qq4hW/As5B6pqIqN8bCszIEgIZBBCsO
7FDG0v020kIjGraDThUOZA1vHCaWLf9eSZpRZ3izFQY/I+iyDzuiixajLsXMtROt
xbuT4GqgWH8vF8U2qiBptZ4rNyusFDOLlWt2xiDq+xWkUMmtFD5hIF7qqiIFSQN0
vjqBCvom3z/OsOTOsyzVOzu0bFTV2sT5c91EpwKzzwB6RbyJngDJ0okxZg9aJG9x
4WSjLO2UzpTPIJKleK+5JD0HuB7FkvuqOdAT8MtZsbUpf5DVY80YE/X/u3i50VbP
YsElQG+3JRUf1pS9sn3un4cJWhcJZqAHMymeskhbmqXeBJdEewzinYrGl8AhqKRz
k8L82BsS51FcLQIGUNgHb2OPHNnZ/Sc/9TzIJ/fhgrAOnBzxDesW4FuPiWw3htTe
IvhngZz3yEOEpMxvrba7PGHeHk+guWDOXIif9EE1NL3k2KL5/eYlhhiy8wF+GIgs
LCBHgixBwt3Nze8wRdSd6emHQUT5nBnIO3yV69FlsdsiHlRrO4mN0FWfsXiFA2CV
uaoXFhOPzcDtaC8em2b9WnTS2d1nwztmVWLRxDxhwkwJ4PvklAaiuY7TbFG4M9EZ
rq8DvrEuVCILy7hU4WPXu15bURFvhXCKpBZE0M6Vhm5V2IVuUHrYe/jYp+uaTGql
lBB0rTSzIMW7pLx6T2a/eONRNsHl6z3e2ddO962KYO15M5gLEBu31x5m6BgnGPaw
kStOdNC5ahIJav3H//wZ6FbYA1mtw7bZDc9StnDiuRdcdrcxSbv6NfNe9NK2Sk1w
hAVwtmQINF0bscIHrnnYWbp9t+DIw7J//Oui6d2+1N3YDC0JMklRyS1lByo1/TWf
CIGgKCefzhBmvV4ci7DtpCQBjmQsK3V0D1M7GnmT2DZ6EQkAxlqROcM58N2jmc7q
11vHxwEOkDdmAGfEqmqz8fCQU9CqwF0LENLIgiu6O836L13NYzuZOy1vFC17MsJH
R9H0s8oEQDmu7XarB18LTHhh4bwzN//ZFOmrOLie1WqMfP9EkMbYUtZctZ8o1W7g
FZCH+Ngecen6EkCgbQ/5o7BSM4cdSeE0QG+P5BkkYJdCQvoQPAkRdQ0zE6A5jas2
o9fOvLftNoofjfoB/DUdxGddB0SKSm3CQxpYqQZH9ITi9JlMsIVdlWjlj7vzrspj
0rHykLREymnDz4trzaHBRWXwOYwynFzbPwxyOS6Wv6ZqB30/HnHp0DUlb+sJsb3v
KmKkYBuYSCwa9tEB1+p4jJGt2L1dAodty+bBkxuHd3ZHSip0q+BxEqyaJOgEbHPf
yRo1v4clcyCp+usrSm25jcB5wXPTzMSVOX8jNuwKND9lwemuGlCdoiAj3D5Bv50Q
6aP2ZoxtVpbkRvvz+W43Ad2JFVd2JmUctp1Af9PXrc23uLCSnpAjOWcUiyUZlbTs
UKpox6Bn25s8Vx0eaifpsOCFHFSGhciRznvCX6x+8ExxDIpriqXiTvttX3Q9gzcQ
+dT6Z3bbnWu/U9n/fScwJTXx0EG279R7PrQPxU1PIjrebxhl8DtnpqoGCFMM4OR5
0tAGuQSBKH4qU2rtj06w6rIewQYS6paXI4wB22uXEeIEU/ek/10Rg0YQN/Sd3Vii
2Oc4n23+pPpqWQ0paSGigc3skE2ktZbOhCR5xTnyQFtJU3nhoPkbWGvXYE6SGwyJ
n5t/cX9JtR5BWNCKGeRIG4Ta/MDlACRg9xaVt3RLdLhrjdZl2a7yrd9kfFKCkK6V
/otXn2zR5T70WlFZ9rd14uCI8LFgeMgbL/VwZrrGKSbuLzVt4j2HuhaiRFP+c/+5
Vqry519+zZcCYM+O0TcMXRdbgd6boer5uSZopf1W1IaK/zGnLswH8gSKM3pFfEHb
ymMM/+kSuL6RkjRMjO2f7XtjIKrPDjC5Fxv8Tm9kkaSmN3WNn/ryGIf7kLbin8Hn
5x1pFIuObAZQ9gvMTj6HSjmdb5bljSAUysXSmT01/tqzizjxRkxG5NfInQh8eL4+
lAUvqG01kkWmBd6afTaoExrC22O92uZnQGQru09hSgrElljyQ3CL4wfvnOL3IDNg
1FJUtyJfAwK707h7taEBiiYiBYMC2ihafPMtUmrd4BBcLlicQdNEzjHtAtZn7vz/
pptcPUbslOKgL9rSKG9Auj/NYqZuJLJsEVTpts17E5vjdMH94tzoGio83LwuQaKy
LYYtTwef8a3yXAO/54QSenjHTpyvH8tv9t69xLorq2iMBsOHFXRzKYN60DDjdBE2
T6cbZ9oXijyLXtSJ6sqw+iMUXrnzmDNWLquzZJ87e2pe6JqgfTVDNCE7ZOTBhlgV
TOHRAwu8CWjoWg6VqHg/HQAMm4lbp/BlK0ahadvVAf9VrOB/4hzuWQqwY8ggvTif
YbTLUx0ApG0cwrh7Y3B+LNOBEqUw83Wt3nNgc9FgL5/b7roPdlqPvBXN51G3pPy6
/3KofxBGSR9DAgEwJc7TguegagzXCZWPmpdFXWmaqZ50u+V5/hrCkkavSH192mOF
yYuuy3wXEDYddPCZIr+GpbYnrs9xcZcJwEZlWRd2lZV1e3NHfSN3yayyXK45CmPt
khG3du3z4GeX4oQuDRgzhnUtdzgJxLJync14Q0LFQkUUif7xXDza5Rxih9V3AAW8
Lj7PyQsgTZAqYgsRLU9C5h5Yz7zniP9+hmI5wExdQfY4Mj7lBtiVnfHGtnwMSuIz
yTRU6lKUJ56zgnjG127TtlYEBgYdwXReWNbepn5ZSJXaOhQbY+G9IV086xUSvWS/
5T6bLLLXgXyQqmfhCSngBGf+gZqV83YmyXUkbVRy630amVQ4X7M5/4H8GWPwmsVh
eObiqgGt6QJwBfQumYBygupcxYmu8YZC2fDNkzMFX/xaI26bueDnMZvCjLs8ehqF
+wptHJgwg79nfj7zKwEOlqq7h7yZJ8v746wc6EokdfAiTUESEi0DjCNaMq2Q6TL4
OY85QwUQ52jcn1qfXUDIBw3GlxGwcLDMZGznfx4shEPH8WPBQqUNwX8flndvTh/z
PLBcECdB2nmu8w6IuRW5FsCYP1FMnopa2ctyBiCbFhzCUF/zboviR4sh2mWrjIBG
vX5ddPCYpSm/BdfuwYORVWpuYDB/PsgQ25iMIj0Ojj4sW1poiQXPDUdXMRS6lV/t
+IP5FDcD17oYKE6fPd7EpN5EEhQvZyYWpwbARRnzhT2fz7mVbj0PzMXOcup6JPKA
zjC0ozKekEkYTUgWL5H9Dn5r2oe3X6Mb3b5dLopFdZHMw84pJ+PkkrWa4BXGZWGG
JKAHYlywtUHoa5NN2QG+4pAb4YWCPCqJF0DG1jXwvZllWoPeTttjpnOdQ2G3R8X5
5kajSeNCgF0PnTakgVytuqyzqcWUI0hi5rmOJFXlpuYGX6r3CKEJa+2kk6NUz+q8
NrsrvwoD55At9WCRrWDqAaGIs8HI301ceKU+8GQXpSKyzUarkxli2kj5+0qqxVD0
bIdZawMPG9Y8hxxgmAvDi4QDy9u/hDaCjvQcuuFrA5v+2UdUOOiwZZukfsAcmHSx
r9h1T4DJRbrJ2AIQ7ZcQvLHtnRlKr8Sguf+DawKNteUbe3tqKQ8oHRGVbOtU99M+
K7Vw0n2jsQmk+cuB4Wn19EzvhXH8Xmw8b1OF3xW+igq4ZMdjmGIteD08+v7D7ZdB
G5f8E27Tthu+/RHOPH62ywtumoDacJN45ZIo+pjARw8O7DGYVYpWWAKhK/+OKCNQ
L+LWARsh+XRmkaCS1+PlnVPOsmlLsgTuMeFIwM4sXo4IYhTWgbhxEHm9YkYc+JQK
+nSBXQ1NjeWKiEXs98Eo8UUbTajCLReJ6Z8p5En3/E2Twwou71AUpQ5Q8kz0HE97
2YixccbT9xMQ2v1TB66cNp0K0Po1G7JGAbjxbhdOiiEeCAfJXPtZKpvSSbHldpnY
W4JhWwFMMzaEd8PdnScFO09qiO/EtaHCe1HSD5OIEA1S0KK8zqn0alCLJ6SsRxgb
hN63zJzhak7dvuLYIhqmsK1uUhDVC1VmVBAugpIBguhqP8joD63fCn/dS73GpK9y
U1fwgazipFyWKrC2Bxgw8RaKaBLXOUfzK9t4yNuAD07K82duqUglkSa+OZ21wGWk
6MF0djxwL45tmtwZi+4GAWF4UtbFsU2DxOBCbm4/3N8GTLwBfFspseUoxhGbsbu+
7mENoc5uYa5q+dV30TFkiOA6tSdB31yjbzOz3+cvqZqCqq8tfwoQJrSby7WRCcyo
5NmfhoqJa2Ze7EUzCbmrTDGrKiLvdq8baM4eisxbj7saRvmiN8BLNHV7bzinoQEx
SYxMh2YqTwX33nu/MCRKB0JOUMXKF/5gsebVwNo86bQF2lS7pMCNICoJsroYUljx
eZYrhddagWy0zAwJZ35yOjbO7ZQCa6zF1KHVJU51c6rLtT7kqXUxbDq1zOa7xyOF
EQNlthy67SjIMPniRVdXV0sl7hyTedVBg2/6hAwio8jlybioNPs5K4jvZ+Ee2jfo
pIjMtHponGIr8vZDrHFUjb3dHNNE3CXXW9y8X62xLWo4bZAI6Y9lsVrBtbi5g+gg
8dxJqlFmOb97YWZx7GRIx+L4GfVOWB7yvNup1s4osppNKUslthoJljKOqwrTl/5+
+jZJU4cdmt2llWHlCwHMWa+gX2Fo6BR/+xkRc/6o27aWSL89qoUE8vzvDYZt25X/
FGVcG0/y8tBbAACeyTFRhubJEWV4iBrghrfxyWAB/DVDUdb4L29m/zewxAP+/nGa
4RBG9fpBrNUaLoybH73REL1uILidafScjGyN7jxEVOIx1pYAly4yVn0lOCBONN5V
2k+2MP7e0xrpi1/jhNFapmmDaYAna4mYa0BBuCEOl1nPbpmRyHZIVkjJkJTGXJHM
5SZ8fOULm+UbdlwW0fBodKWZiQoC4E2CwdAoqno9qPZFmHDlnHkRf7F8bz9lo+J6
Lj3V957NucfXukCKsWDgTxy/ECUSeyJo0BCrs4GjoLGy4kROhbZXaqhFyne+pv7v
/1ZJJTXo06aitkJ8VxERZf7pOMsAI3bvHPY1A1u8bDNXRW6jaEW1GqLZboBdJ+/H
rGPuEyQK7TrcGxRm6AjbL8q38CABLpwRZsFwmEku+YdqgMLjXQO6thfDRwy/lALm
TXcmW+DnE49umil7N8ne+AcpZI1eSmGRGQ0+eIfgIqwIZOj4gsONJoLMmQ41SxyU
POicACV8WNKzJmOrzPeH1pyrGDsdDD/tU0MX4RrTY+YkUwGyzG3o4CVj46dJWnJa
jkECk/xrvQQQmLwobjT108UN18tuuIlwPv5CGgOYBw7twzUNJoE48NML205msxa1
ElLtl/NF1hh5FP6P2c09aGKdDmfM5ecNy3Unsf1gzc4SSiOsf5OpIKggyqKH+7G0
TcNaO1bxh1lZAyojIco1FrSXueGWRJ2ZFAM6OjmazzWpkgtcx9BYGr17PneZWK/S
NOTBxTJb6XJraj7Bx/tpaihXvd5+U6TYxoZtFQJqgX2lOwgGQFYTAkY/F6ZJ784V
yUrAl9RpPisA2JO5bMmKmB4N0oIt8I2evtg0fZrDQ7NnhhzpbYv6fd+6Q9lY6fqs
pSLLSusyUqvW6kwSgXrxd1c4asrMfYAhA0my9DAwKjdqSdTlQ9EWKks0bh15dvmf
+Wt43o8APk8VbJlmzA/rRmIg2pyueK6DL77NDWWIAdbVL3UNE8h8nkXr6JhiKYzM
8vG17XatYvbX/U4GaDKfUVWv5QFWVWCvz2MlhHBtZN/oW0mdmrVCcE2P7w0BNINv
/yeGFJB5fVIBsWl/EDi7y1TVT077I3hAKuJP5yqeSqX5MHWjPhP1r54I/2cGMt3R
LpxegLtwEarWvY18mAjIhtrl9xj01sNGslOOL+cowpoCg5btv67IBzdxQMTqYyoG
kRKKO0H4RN+0ePlipfQHmeTxIRM2xNBPtIhBfnj9fDcGSgHAs5WINJ9XUXoaEtN6
VXu9avisS4sqD1pmdtcASm+H0DIyUko8cDqGNF/Zf7NaMajtH/e+0BWrduJW82kk
0m5xPbqs9C8Uiz1MVhcrMe0Ubk5dL5IewHe4WZZ6pDtmWtzb4EKnLUwZExWDwO4F
r2d1dLbS7qEam6enq8q6080E4eF9p6qB/P3wLN/qzH6F2rlYH+PgjKRLYoqCx8Ui
yV41H3lnHF+SepY8E28Pz8SDsW3J7yoiaHR/dWXB8DZGoLVWeRJ3n+/hK81W1saO
/fjKDoHHNuuFuefccqmhfU61Imh35mUj657bwyIo1hmVJz94cv1LXMKah/SgeVbk
kSJpowad4ZyPGMwT0Lh3Mh2N0tVtOqok7Fjiidv1iCqQM+Qc7NzG5VCgkey+k41N
gzH+ljCAcNPMzqSHEmY1ewg9mexkCc2fF5kqwFjPeqROe/9e+pLwzyao+t8100sq
y9daBAysiLjIQbHo925hIzXAW4w3iMaLRoPECq6bOVVXTZ0zFi+qRjnYKRYJAUBp
FfeWT30VwGwjEmZwS4lnECrgpvYb7HIOddIBUkGnw17wFCDNKk3vQbA30zDrSjf6
wEwZm+nowmdb7f63Imahm0VflfYrvS7jtst0Ai9IBGJ7N3R+yqJX5WbVKjsV8rXT
8AE/9WItRxPsgfmMcGMK9dS7O/VmHGfGDCgY6w9tuGJXPBz+Z50mAKs797qHiMyY
RfDBisVGXG1GBz8q7n8d1qHFea8rhKN6WPQR6RPWRs/8sRP+yxdKvNf8LmPXNZYg
XreCAP8QhIKQq7WO1tmHI1xd9j8pCVVVXlkjNiZNcY2aK0mELXT/1NxSNQOp95Ff
+JO8h6VW8FmBUju84S2hv5v1o0TtvroQNGWTi7eL0RM0wtqg6Kq9uXnXOK5Iz/T3
NeP+YElnuVWvr3FAy3r/rnWVba77jiSj+5SbVzswikrYDS9NacUs9APXLm5HPFXZ
JivtMPuxLL3YJZN+8EzByKSy4zyRRbQOZMG3S+aPm6XODHx560xw8sgqwMHbdztB
YeR51cFlLY+IW1tJGAgonsdAUPo9/u3JdJ8zR7o9/hnVj7Nw8R6Wp8geAb5e4NiE
wXaGSkIyNh0W5txX2w090+Ov++MwaJ1ZH/aQKkxFPWqEHcWRX7wolt9+L7hsdE1O
fYlIhNpic2ydE+BaVsbuoNWtUHM9QiAHsrTk7hN5hfB25IcYjv15ZgzG79oyoyFI
Ystdmksze2kxRfbz/HCTcDTUQs0nFjMS5xszxMOp0TTRpXjWwehb5M0psmRK5geQ
GXwsYHnm6NC/7SLgJZTviBEcwUBCFTYKRCmZnqPPzFVfEosuig7eldsvt4861P3q
PzWhVPU6ak4UyOvZgYBPVkQCFRCBo/QPaoAR7pd7sjgAZYnekeeuCIh1gJ7KJtH/
+SNPvU8khyJGLEa/RYx6B6fF1SZRFxP63TbyS1rZ4HXZwnNKKkRFFZqDVSGDtNq2
ApBXdOsdi3yYwjvLS9vZTmvH7scmMOE2FneZN5vN6RuS5vn+YPwDd0Jmd/jKPR8O
piDq1eVyYZ0V1gPA/rLto9EmqgB72GvJVjr+uNPjonxeYmR9Iq3H+XlXlUSD+Pop
obbBhe1FqRHphZjzRWhRZkAjxEASaeAKsndMIajVaMdZS4li9xFNQnTQe2/DchhN
MTJhDXpoPsUXiygbWBEzCkLkN+Kz3JoE2/tJsNbyZVlDHwk89SiV8ges0M5cvY+6
i+TsWBvkKy+ZAwYvG6BicTH3vu/eASpQePUPQLdGXWU1+j7ufNvf5NL5Hh0AP2Ki
CiKnUNQhP89oIQJArtyboV3WkXBQ5QZP9o239Tl6es9fbL4k3przX+y2xB3nXUNK
7FMqF6CPZsSzDJNJyIA1hkcXH3SGfA3KCO1jp6/Pw3oogw0QNAxtrycvjdmawb+g
L/jVH/7PekiYATM1lB4RP6igto41vW7hlvy9dRLdy8qZ9ZCK9/IQ4JhHjUQu3Axs
hLA/7OcjxSqkh2gyGIuoY/mqloQSycEx1hxpMQ7m4IduPhYyNncpxomSVlZZTtNR
nvBOoD3bXUolq5usqwagkxLUwG21BliA3loxlDs6yk+cG+/rbbBGLA1G2On27ua+
+8gupEVZxL1dN+ILJbskpDreTo1z0V/9N9T3thNyEl2qSRw3l2kCwPUxbBzJXjhM
JVOjiWRjnowFcC7Vn4fP8t8U4BssQrNFifylbclrqRema+5CXAXndnviiHBkP9jF
GFjPMMQJ786N3RM1SMh4JM7Jjf8jV5DMX7rXYV1gQGvC1TAu89HN2R37+lvCSZPW
EpiG3Fbc1uKY7rYcfnqn2msr+1SOkcjBD6mRgKgeOBI36DcaOYI2zBfKcYZBZxR7
AfyrAOrsVf7YPKHegumt3bXSBoB8zIEroQEjgT63D84X584eUtcOO8idjmuhtk+Y
ZOmhMwIIcLar3n75H/R2fALoc+ldpPtwdROdxkzdwslxtBnkKjg/vcV8m9KlaZk0
1kfqC9/XBhIRs7zMxyObI6t8HyAUqQdvXpy5BbTde+iWzJ5Qx24kZJMCipGAK3WA
4mCirX9NEhq/vX4sSggq3yzmZSLVUB5zXebPNVP4ENjzdnRxglBubJLCknqLYwGM
SLGLdzORoEz2C+5MhEz16RpcuHI7KJf9FjtHB6E6BK+q5PnLW0SuXSa9DfPVPomU
FnwXFt+eDZugMXwC/Zr7EnzIm88jM1/Hb6biGrHpr55wGPtGvBLruPVht2MC8VUZ
OPVWSboD5uAcqaUQLCcvXBckl7q3dm5yXxLHV4INW5AJNJz/qkyGZhLE02THWTV6
Oxs32u5TA+WPOXNxiSLfYDJmlW5zxKteOMZt3EBYRflCZd1d2bsaonj6bKQr3k1L
pHF/x5KvnvtANe2j5LRBxhnQihRQrHYOe9fs/+DOv4sVaSlqcuAIc1GOOUrUUni1
B7NifRkBn4JJBbGwEOGqMiR95m//zm2XH2NwC5SCKYJ3Uql1TkzHUog0mmwkQgh3
CIjgNCxEIKto1Rz4wIImR/Af2e/5B66EQekQa47m5cK6SKjv8SxPVcKyEFHAkcio
O/XcV59wSWEiBYY/1MG/Mo0s1IVx29Ap3L23BVxip6rcUPCdHkNXrOWgkVstWwGM
+qRUw6yLQZqOvOjxUJBq1ZXvreHJYMIBcCQ9iG/33e+vgIuiRZyLT2WjcVs8Ni5j
3NVj1B89g6hXQTjpgeH1szXEsf5K2quNYRECmPfkQp4X4EVQ8pmwD9W36PGbhDGs
TrTEzfmbmSn/DdGn7tiGSZsiJ+F1ujLHcAXrXX02WilX5KvJygIEY2dpyEZd/lhl
IHf65xxeFJmKo4X7/5VN/j4CJSjhBqOTqonPhkEl3I1Uq12aKi5qfjHtevi+f84W
O39tQy8Wppvp+zsUHF6QIgGcwjNiKLSU6N6/RaiXUlSeRji8znrwtQ1KIB320oN2
8Sr+vQ+WYkAMU5axIc8Jlc3bp+741Bk0y+4bpWVqjGxykNPS2U44d7HAm8fE2ZFa
nHtF2y8LlACnD96TyUCcL1cWAMp6l3EhZ5aYoFDUrJ/s4y3jGhBwJ87AJJHPx5ur
czsh0Nl4xtPIIlM0xtdECrbBKSCi6R1tyevAoAYQNj9bhbXBbGY68x/9j6NOTxU2
goxkElk1onUFBVaB12FgHcXwJFFvJZZTeEqAHGQuQD6VYV5n89S7BIdqCGWwrT8B
61YhCJXgexzNA5fBG90snxQe2lD6JLbJyuE0UqcpTzn7XbE+WZf18jxJkXb9WyLD
tT5WjfAPozO37N2dxYZogLp7UfqVhUlZwWesXfHfxKORefG6F+iBVSxMFp3osuJC
V0Qke132Y4IKjeJvuc/IH3EFD1sO3+oV08NfUcfNNCuVAC5CRNkVmIC4+RV8nj5y
L7f/wNbH2Ty6WUfjyS+Q9Ihq0sCw/RnH084RBPASmp7u4og2j8bB64gvXgRP4evh
1niuHB1ZYpuURaTLBWYpeC19nMVL6kZSsOAayoT9P/aSvuGfdlfw1tAPupGjwqYV
nxNdMXV+XtZwcDobvWWXfyvQGCRDOjudUJVhO7ROIvSwsnglOdDfOZMrsoo0/A/Q
NcNQhNlOKy15neVWygIUbkNY9mf92BGPm4G8FhVvfY9JJmWIEqCpUix96aA7KXjr
LOniic/DyaAAbj1Grn/dzxSLc+3RdB2Y2Qx2OwnATOLAX4umb6HGyZW4+ac75/WE
E7EHbQhyYu5Nl4p2d503POPtz/smv/MPdhIhk9cvz+UfMdz1XVaV+WOAI9fLajMl
tGPkUliBPl7UTO+nu3n4DR7vNm6rIVMQ3oarRhRD0m0Ga+ytTOYkruqjj6M50euf
vvUChO6g0P+LWrCfY58ozmFy/xrtObDa+Opgz/x9q3fmvhr/t9cIF8x2zEnUzYA3
GBnl7Xr8sEELGnDo66mFO6X7nXn8KeSW6NoK/qz7bOKIsmVJsU5dw/4xxyQGg1ds
0i0km/4ghPtX1gwdY+2DI8cmWUxQFk1VXA8yxPSf+yY2YI7e6H1bELqlQjW6SwLv
K/4/U6Ptvhc24XJNUbYgJkP6z+6uUVyie2YtvPS2GdDsiQk493fS3Y4RdquGki/h
+K3sZ+Ho3nh5ysxbUnnTJIQzZ+sTDOdR3mw34gRzFVbxABjjqM28F9VH/dCSOqpF
695V/rnm+/qsUl3I4FGTxDAKmZgBCCThbN2l02Ic4bKaV/ioU04cpdC1iP7u+elp
t6lo3bkFKcavINvyMS4QMCkZEaKmVQp3m2KSc/e5sYzQQuv8KcEQKtIuI/KZi32B
CAukoe8JN34ipBFWSxMsEmCuPh8JkvlcwBPTA1GYwtxtYAM8i6mRqK0F083M5IlA
xVFjL1eirEXOIcGC3JIrUFvAwzRg1j1cM5DwJJknPpHONdAh7erxewz6tOSm93tD
qNl1b0ZDqDPUaBdbD0JTwxUvA+zN13if8w0v5sEad77KiL8Fdj18+c/5ErInZCQw
3Ch6M3IgTxiJLsgnOkwFNJ1Y32ez0RzyU6VL6VrUSzq0V8SRb5YEuxMf5HS8Gear
4kacW0iLaxA3OZg5zFoBjCKMQOJ5xR48bdSu1fatKa3IFrjnw1RfxtIqBbhBndKn
POe6VMLeRJ7Ok50Bt5x0sZV3mDhSwhg8xrURZxU918dyyEdOaIWlaBRSSYOu4+Dd
1W7A2WW/Ozh4DrXE/lmIIjV5tWTMa+FfNpup1rf525Moi6FI0vbokxxzUeBWbLag
f9w5l3Y3T73TVyzyuPQe47+TvBr4kR94Q01fx5grRPk7tzgNTVdovU+MDz+MRFSn
hj0Bm302Z7SKtqc5SP4QSWuFW0bQs+tFSQ065f/DGerWNZcc2m4x32wKKibcWFfa
KvIno4a/FmllFbz4VSNeGoQNWvmvYzzM5a9Xsw5h8zzvVTdbP6ygJwUkOMTZUlmx
EvjVRaM/LJAGZHaW1rVXm9SPOJN8eXoWijIKxhFrIHRjeMaok0uI4u1ucLN15Usx
yXSTrJSwqBwxFiI+Yq/6XHpqeqEePWElW2Zos4FeqU++AfkArWJZQGbndNmHEYQW
vjh2aD2C5Ne0M631Fju33lmYYh8u52Y3HJKKydDtN3RxLjxvq5vcnewDbVZYMgQ9
qidWsqR+6VvvRL6XCIi7+idqfXVftpvwoNLbP2F6+qj6Mp7FmwI6410WDBmA5p+j
KObjlHbZnEsQWhwLcvLjjugvfNhi0h/VpWDiNq8trlm8mvwg6R9vGOZTftsV2n7S
/81Fazjn11UZtRtOZ2dXpdVSCV47DYYSqfdQUkgqOpd18BjYeWz9nqXoVkDOTFLS
uksHHXlTSNHUMjsiBCDs67dQLF8biCF6Yq1yy+1ahH14rvPi3lLeBUJ+A7Du83kG
np3gEQCv9Y9hTs5cq4WXC+zvvtG3W/DU+RDD1WvZlLuR2++hmOYteUiLov97Y6XO
hnyiI4ghlWcXL4TbyGaUe/wRDpoVGk+NTZKe3jHTwjIfFftbH4VMEvW8RhYX85vx
7aTo0pK5Ek872MkM5SQsDEB1JZl5qUP/Fc4RXrp55XxZxZrsMq5NQegXVcE9a+GF
lJD/ENmYzOIqMSpK+haniXaZJMckqie9TesWZmNxYrrl+DsKIwEIQdlOj2Cfzwga
3I+DMgQH/JZdO3Ql14iEKvoaQEHfFwxTGuUbN7xdeyFgayEnjvT/XETrUViXfWra
10DtTvfThHUN5OWs4XvkMf52gFWzDyIrHo+K9BkZZGZP3vLleVyuW9+m7RtuiW7s
A/f+eeikSPGgpCRjVBT+QmTOssm00ycveBVgTPACpca8WGri9e+OBLdf07QpTsDQ
1hPKFnHRd48q1Ac8T0qli8nJueXJI4533DEKIEpCkkfhSCQstiOX1adwSSaWpu2D
Uyz27OreCH4PTDXqaIwmNuNDErT7mW3YEaiOjUT+8cEf7D4zrtGbDq0AtPmtaeQ+
xIyXWEosWV8gWjgtzb3NdEoEHDbpxeQB5nvLkDk6+UYEziktE3CuQzigqwQhpzHN
ZOI5eGryk+vPTyrXcb+BG8wn26T/kaBW0zG+lR+G/n9qBcuZwEDnB93RmwztK++J
Tu4GlXWSkqvLzMtzhCn4bZHAVKUrDe7otYVKRzTfz6/Fn/jS0qwUwSiqz03ohFk4
kVfSKLDn9ydQmdeg7DgyZ5dwkA3Blx/lgCZm2BpYgYZgzlbzOxz5ptPkouat5ZYt
ZxHV/Ldrar2miYJ4o5hMUpaDOpQMx4kZgUK14pFmCkuQMOBMrx64bhTs86px1CRv
ehKAvnH0Uz4GvarKcIRrODMX8S1jdfB68kv5sgF8Gps+gboGaObZ8bSOTcO+Ktsx
qV3J0zYM697RoeFDeD5r5mwqFgFhqUJwfCTWb9Ix/tb8trCvK7OFtRy1StisxIoF
3d9+V5utrOiJVajSk4PVs0WCAGVaVuvAQZ6Bwz/EKNxqKD46P+k83HCbLDC0EMtU
n8Z59dVBVifipPLuGAv83pZUgeTRKNjMzjgtJT6f58F78h99kX6kaZUunzPjJm1G
pzZXzA/DgintVNrE746z5hFckkuv4usjPoQq5Tj+v0q274UeUfgy85MbWTBqtw/2
whw2RjjKDTzzesb5/qykWNnttdueWC/S/r26H9eDN3S/4g1rouDZPbFMYpCh2J1r
OLCcpBwadeGuSZbDxND66BchBtuILJ8dl3n8oDFpckS5KjsRZRSfnsFpLOnVGQLk
3vwj9m1Q3zv3GguY2N4/cjdbFH6w9orYbcxVXBLkwM/Ee8hffVgPa+camom5Ghgs
/CwpP81uQFs5MRBtHUyYgxDrY8hznWMOWoO0wB8SJWRJBblTwKXkDDD3n6f9OEfk
ZK5OHe/E4ZJ7TytlUY4c0AsdJR+lEOWEmEwpZSXyuUDCASn32mD31T23BS43QC5/
COWQF7upL63sQBGk2hCnQfpZ/Uj26IBrlk1QiAXTnhos1guJ1KBpk3m+99oGUHHp
QJfmQvY9ZJj6lRt6DA5xtsAF3JGjn6l7VJjECyWp50z81P+eQAfrNB6lsPoZyvb/
+qRB86x1mIPfCE0hpE7iMmuichxkbVwYd9jePd7IqFSTOK0sYh6qcGjQ/xDSRA7s
R7H14k2BDiV6RAa7aEhyYEr5X8Ba0RNLJM0BqWKuR5legbsdtQ5UAlmDSjfTMjwI
rznBlGxm1Tm+NvxZeayD7cyzN+fk73HV1Tg2TDsZ5VztP/4zIzKnKQa3BiGY8zNM
nEqletMPySeIfUmeitU1h7RLQAAkV7+FYBqVcsmiArAs/xuHwrisK/nsOESmguUU
U5TFa4A5vYNl0WK3gqy82TWIhD3bx9sac6CPeB7V+LWC/A7CxMFNv9q6QBxviBAq
IUa2n+ffpv052fTesVqhoYC2lGSLxIPdqQuGqG/tPsHYDb0Idc9GqGVz/G4ywf0K
0teX4DzkvfEvOLaJFQuIRWUOvd68C4XIh1YAT0uothBxRZBax1067Eecs1WtQW7m
k97IUN0Hn00stmcXal527j8T2HqxyuwtVmiZ3OEXzJHaTnj2zIIEeTQvC99VQKrO
5Wk5iOhfWSxa0JtMHrCH8UhGFUpENFhJJU/2SNt9EHaDln8d4cCHjCm11sjeRMEx
8532MNmR2CiAx5QGHTWlryw/v4MDBf05rm7lSsL+c4viJBAzMq59SqELnzZ7TJiP
PropIuYDmyc8AUva8Nc3TzDrKIZ53/6XGpStR5WGJjCoGS7VM9v9aW1vIMOp8ABO
5czo/SEKk9VG2d3W6aRh0Bze3uUCTe8vbYjocowSLveYwoZXaNiQ90sHwOlhi+9f
Hlc5uN70UUrbXjOTtjoukipdYBnndbd2JwQ0D4A2zkUcso3C2zyq0gwB4mSqCj3D
at+24kxvqxFKg+9UUGVDRzWHl9cVEUk2N8/G+3Q5FQVIQyxfGlJ60iwAFBYeM/a8
toQigt8xn/ygtp9M0EclpNVio2pOHgUKX4C5I0JilT9JbTlsqRQ2izc+XBAYo2Kr
Rw62PM66S4I+9Dyno4kf1+M4t1ugq0WLOOO+ZO9g91RBK0j85zdDNSCgqX+W9Bot
9FzoH0f8YVoN04y03bxrq6nqIMuHUBtX70dh1OBC1COP3H6ODt3os8PNn2ehIPM4
GSTI4uAHF+jYeAdZbdKX9YnQKEyoeiQO+YqhaBlA0gAqtb/TD0d0eabwpzIXzl5z
gL09os/oL4h8LwfSerjx2Z6rHiJMO6FZLN9WAuc0IsnnWlhCiY/2L5v14v/0pe/R
+GP/DfDUEDGAtaqJFwncWr0RQqcEuuJ6KBnhx0SKkRYZdqjrFpRKwi9PaqqaBy1W
KE5nk8L8Lov+x4uaB+PIKoN/SqkrNRDbNgxsipdGO9MrwjC677kJhPEYPBLtgt2L
JyrLtNc8//RgJlwRzjvruzramCMcTE2Di/W1L2ps3hujHBsb9S1iDt6N5U19sD6S
JnPywgjNNoOd6Yie7hYQq+LNPQgsxRhN2p/yTVLg6f+KqSN9EtmzP6lVzWk5srs1
4VuTBDj2N1DEP8Rvm4GdrE54MxabWc56ycfTJTQ3etZmnQg5Ge3p/+enu9uSCYT7
gYEVoMkGKZj+Ho2yC37rNE1KdxFs4pcfjYKKGROHQeyDZOy6kIqvE2tYfkBwqI5O
ApUT5Dy8Hnx1vkDWBDbREXWvii0L3teLKR1pvh3x04588qGQYoayU69e34kH/RXA
Q1I3h635aDJPsNEXgC9oUmHW++gibZo3tSDO2dYhkWJKiSYjX3C7643BD4kGvvgS
FgvPdIakg/CVKZkrwdc6fAkEjYMiu90/RIXMDp0826G/kaxqtlVynzt6EcGN3YLt
2b80o2SGlAG0f18o8ll2p9HM8cCSz8MW5qX/zIz5urmxnA4ZJ9Q7+2fQ0Q2S/qE8
OqyxgyLQlTDjOGMEMyaQJ71Ql8YlIDCZ+8yuZMkuR7gcr//86OmGrbE07w+LSYIL
de/89bv3J5AqgBIy0pW0jDQASusngjD0xx5tflKnpp/xpPJsIfY54wrtR/u7mhsz
KiOm5FBPUmUQ8LDN0EFA7f/ecqPlKR6fr+W2jNgj6jXSZ+Ag/4b6kdU05WJgOWCy
cGYlg9GOVhUq+StfTiX6lkKbO3S4XywfI4ool3KdUvrAjp+IMx5Ws4okzvig5tZ+
fF2co8IXnNHhnaxTRxQI4Z4tPX6XkOaKtuZ035WiUPbBuc3VkSnAcQyxb70BLVIH
/YirYvDFyFotX6qwdAIw342kn8rpkNPUyWztDhKOsw5Zpa1+dVQWqmWicvV6R/Qq
b0elOBhVZ7CBWtcdmLNOuGyR+J1ROOYR62OBv6WdTlMYeNx9UZl/J0BsAB1PXtZX
bbqvny9Tb93HCMjlYRSlkNlGgTUfmJSNZBjX9cUhAR6MEKILmPVBw3ghqSFqBvkj
pBGzgJe9lISxR6D++MFW5l507a2wY6x2vNdr7J5FeHPv7kaKufZTBk1tG5nsSOQc
/YesnbpcSoGYfrFMkAPgtd4qGxde7jT8ST48fBOy+en/CIzcj8eHbYF05ne192L/
wBKOCLVuccs0Lix7rgZT2GnYufMcHpTdPQGswcvIkMs3uIqNjKopAdSPuzgru8vl
xjUAtbQDOA1HQU36eAgZdAw4+bSZXjPoaD8DzUhVLne3aiieG801PXa28TKwnVOr
m8+w6zY/yodg9Wg0LkFUaegT3CJveVzot12/+aCK0Zt/eFsOlZhWfWhv6xnZpuTZ
SLqpR1YeZGvnXQHXeIDdMGJ0/4vP2AvdBfdi7QTKnzUhpIHgcDYj0ZXCtwM5rsd/
lX5uFTyuQgZqWyXXlUfRrTL2dUd+sg2Du7UOV1PcggZ9dnQTYGluoYHlFj0KHp0s
GWB/gJq29MYKqZ3whkjJGYr930/k2ngpO5k4WocE6YSJr0f6FJChYN1FOpFNFJuA
GdkMxmX4Tvpa+pNf3at8KfjucqSmBSrN6ofhh4JWzF7hqkbM2VrWyJjS4v68yLLp
0B3pEYjUv9CNq5KFrF/p2htCkY4TuuhcwenHadT/uSudvEotwyKv4wfNFNYzwwWV
u/AMvauDiGxeYkgvltsUrQc/FNScCqo6B4HqJNRyyrlGF0VRA7EVjv1viutin/OL
07EEkXUCm5LiJ0nCk1+QK9J5gWx55g8xe1YVc1mnONex238wQKWFDyxv/jbHHvfh
BZFo/DE4QwM4FJCtzG7gH7JQIwjjcogTr4a2w5sbkbWtJapeGmIAKsM9ah/gQi33
CGPYLPH8sA3pL6oJ6mMGun/Q8TTkN3K9CARJdr2p2lmlUZKX4VH8NabvnJiSxglQ
PS7QCOJauCNV25tj7RV4NG4QBV2BSWm5U8LwxHh+5lf1fvzMWM+1Y+DQJwOhMwex
wAdEhSxQfDCfmybkayvknullZhF+SSTJKWV8PYE8AkizjxVl3ZV0Osb6S0d4J2LK
cnczAydFM/r6HbgkGPyUS8Zr2+DQieApOuLlOMTRqL1KTng0BiOb8fehkqxtYXaG
nkw1OMJKKynAANVafu1PS0fGGHRGGhSKkMhCyttf993K20oPbtB+uHnS4AMM29iJ
tekHCSsTD0ciu0BmLVORUgqdnBukOd/6KRdW4Un6zAVpUZX5O/cc7gwJgg9zInQ+
RCEsLv/2M8C/1l3C0J076UEy66YTnMI429R54zGAOkMx6LFEwPss6MZH3BUzn0x2
YtSGbVqIua77eJpICB6e8eon+tVi9qY01F2A6Nnwi8HdXOZuaLY9FwbnLTOmfCEK
9wcKHxfFxk6/yv6IuBMhbFYBxmoYgCKznpWKJ5rgGvKlx0iI6Xx7/ICIKOYkaANH
CvWxmur94xmTlPwFFWKKY94KAAF0rUZq8BJNImPMe918vMLJyVLlnSklMMJ6Xo6P
myTecaC1X4NOk8Cy672DELl2U+RUgczKUz3JyjVqg7Y4INZ1a4ikBdVvcR93ZHFN
yzVgdfotMzzRsD3V6MAiQPApG1AgulgveSAIrBG2iBKabgpS87u1ECJPiFd6j4aJ
3Qo9TaxUQN3itZZLugoi8a6jEwE3LdY5gfGLFC2clmMwvMFnXJh7dTk91OjYJR65
13ZnRUPLVl8rdK4cMrS0LYM/q6umNmua3ErESqDeaQTFETzlDRj5gZLgVqZEYWnB
iDzf8FXHRjRURm5bu6IeW8mgwu8r3tH2iuUV5rxFwPFwXKJ/OrJI4qhBPIWG5yIf
SQPfmTehC7ajRsYjAgd5wlfWJRYYOJAchiLLTxLE7HsxA+Gmd6DUxqtQT8WmfROx
6h3hf369qV/+guzi3LgjMHTf/nXg8b4Hjyb34XT3J6DM94Gn4zGuo5nlQivFSZzo
kvowGaxUIynD5QjHDLVixV7ywm5Dqiu9DvtrVGvGAlfV2eA/WT2FbDJ5uKXpQLfh
UwenAIOZD2cXgvfvojGaDPuLj3kVBCQ9+eUxzCa38468tU/DA9AcioGSpbf30aKU
IK9b1VbPR8XnW8BPPGu3pVvDeopRxAIOTTY0QPWOboCaDAkVkfXkRI2ZN9Zo+rHc
fWIs00bYwkHRb/QkoO6XduOvxLmkJMoDWzDYuoEMH439RvFGK4VyoGvk5W/UewFF
Kk/QCtqdi1qz7nnAr0Uq9i4dR7dp9j/2z2i3o8J+vBsWAOfG02xYLavPkBDn7svu
lQxry0JBJAP6wr9aageVSy3Qy53fMOLdj/rO0l1l20KIykWc8EgXnlyN/Gb9zu1b
Pmul55VRrI/YCjgvqhc/5a4XMAkOBVEt2rZmC2zzmxJYb/t/ULKSaHCIOp1l9Wvx
UyRxHSQMmU/UfcsisUpcsaKHcXdYcvRexzxgEzQpnFXYr6oF9DyANMo8wQ0KMQb6
c0R6XdRHfVqWp2xLu584PyjNoyGYDRVQIojASBKwXqnkB0rbi2Sybj4LXdjkWHzK
k8ffBSiQCMdtopcNxFWJwy5QIwf8OFepz+O6mX4PpRSRwEh19EIXSyWyHpWYgoEm
ahGSAiJ+zIQzmr+c/YlnvT9+Vl5bCNXqRZU9q+BL+bCl+7h0MHT4x9Tn13Ck61A/
dgey8/fctH8vtvyaRSWXBx8FiL8HahuR9Ec3nKHlitMLsPMhVVkt0QLdyulR4Ygk
tDh2OfX/2ullkw8+jCEM0+7izCxrgNoOo6K+Ij/qfZwEh7P6aVTl2RoQytSXafqI
J7Q2eBfHI7Z6bjx7ub7QJYjeT6/urEacE6Ix5VLBsutU9tgSUM8220FI8CCVv6RP
vx28zOR3JnAC4135645p5i1anEbK7sZNhzW0G+mI05tDEbygfROk9tUR4C4BGHI7
STwY33JqgeWNIG//2nsv2HCo3uF0FZzEgmSsgENacTmAmA1j6uLF36b23C8mUL2r
0NHY9+XacLeSW2xDhuQ8lQ==
`protect end_protected