`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6272 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0gQgIG1mJzulW1XOK5NnZR8
C8XqDUtXW7uOWTnSVqbIbmtDsHrDP4hDy/xrzKHF192Ay+3WJJALD720MJgl/Fb3
WX526cB5UnUBzP08hqAcwcYyzPYE7rdK1TGn5qcZBi5AanQ+EAOiFDPzJu/OtV1c
NuJ3fdtyDZjNeBK54DhADn7AwXFIEybbibawP5yvBm+hyrmt4WqW1Q9qLfjX9kNx
crxRbBlwm2tn4/u5mks2BTzAbfcdF3skqu7G+++YH3L32WD/4B/IBSrekJfnhBmN
JhkIv+7FWgpi0BirzCzUnwBnjnSSLohbKtwtvyV/ASrSj6yFWDQ8Oie4f8xncZxQ
0JOIhXP87gKbECixUehhTaNe3qWRIlC6b825WiNFMeTv5rvc4t6E1VGx/SgLTMWy
N6oInQPafoaa0zZlnrhObos1mLkhniTN+VomVi0O41SkeNU6zvLJ/lDf+bzjdXOC
z+Y+mE0we83jmmIvS7MesvIpBZraBP+KTwIINp5tepkdwpl04ya1EbXBpNbwKZBe
yHV5G5VwvzhM6/NALGaVX4jrLOa2GxH64/dZnSsWjNJZE1OFNPTTsarzo7ClptVy
WCefArUvbV9En8VTA7n7OhYOg2dAWNjMlZFDYPRlfVdvZD3nGD9EHuJhJUhCfecR
X7UdIqOvsZ55nY59FqeWIH8LijRExTX5ffZu/EGIq1ZFctWpLEdnI0KrcL4W/u4W
/7sVwcRROSX1SY2fbBuk6AXir4jXU0mv3Eotlv4tbTcOKdUPDAAGsC2miWNMO2Df
b2BIjhacK30qOlacowH6pm2zuf5C9ruGMK0ecKz2ylPeXWYn6yLWg1o+wJawZ8NX
fwyiP8Iiln4GTlcO0ZHkserYkV/Ip/EM06D59oAhNp8oOlyZx7OrNaz5UkY85R+I
25VSYu0EFuBk+vAYF177d9LvjExc4GBzOxFaw84HFkjVwPblUfNHqkx6Bj2JdXCR
qf4+YHdzyYTURMpiRcVVz9stzfvvHZJS3m/s5W+j7Ewun6PKrCopAnyi/5+YOdQw
I+pCGJvgb2jJfdHdJNAf1tLXTwAyECz1QOrtwEhsAWz5FAegGFMolmOBQKMpndp5
kW/JvbQu1DbWzkOrufrLn/wCeOgxHWo+OW0wEvnoNBwTaUEQbHafeHzZV7u2W1ba
FN6u/8mIxrG9NOHbQ1seI46YaWce0OTLOxzp6PuYz+8dfvOjT6IRXNSYbycKQL7C
CjNNPFwYoMDFGlvbqRaYq3+rvYuA71sjnS/gl2Aq01M0DEqIQt3cieo4L+45zfum
M3ZfKc/T7n3bzC4krWr+gWX9DYkgPq5OtVd5YLlsWmLAbTRl/MVKBwtpMTnKFg6F
0IK/muvd4/OE0GSfOCzW0n/qgsZjIx8JB6/lD6u5Z5qddNW3eOBgLhF2h/Rv72Tp
KxyKbh1q4CtGzYVPyL8Efb52boIeeBNCKUfvJZ4rHdvCr0mXpL1F+Ddx4IKOIMMF
cF2LVKaSI3P6l7XF91ax7/jHUpYtkECubCspsvI0hEZFxXJPQ02ifrSaL6HUuKJ4
P0njBWOQBhOZx5AUFZzmw2PS4+dwddDSCkalcEozCFUBkfnUGurWcWmmgaZCN/X7
4yhYqnDI3iTA4HqEWYxxro88SZSo+SBJQ8cLnAfgmOSJ/bO1RVke5YBRCcwUYBLd
PzBalcN9ME31NYVKp5F7xQVLsb3IxAuIgof6TYYxpV+8Gf88L+0FSoIhIXrujab+
DaKJhclLHgjMinOTndFP8dUkj/0HmOa8AYkkk5mseTQg4SkvOERKUiaGgGEclVWj
+kpwnouVAyPZ5bynG68RaZbBKcVEB6YPt5fw0qUghvZThAp3yq4J/xGwdV41aG6I
6esKzs7UpNVCTeFRf0lM8kf86NQPSL71FKnHLUAEcsCeDKTeaivwSU1cgRyYcMBS
7I8qv6tVb+rZFLZWE5EEEJDVLLHdkF1ArJli//KCJsYuvWxsJ4o8OgI0TXVUzdnO
6+kIr/GF3OthVf/vtxkJRbRcJboVp4nt0Viw5ZFrf2xp36hKaHJwSke9MqmjugPu
VgClXuDh+C/8GmaIVaHYHmffP90tjQw+H7NErKBzaFcKv0CFxS+rmj9leJ8axXfu
Myq/3qAYSecg8JgEU5RSCZHpE59VURjs+/Y/Gvo24ZwKAx1XKK/h+YaS/IYjt476
U7OQ/I6Enb5Gjuau6MCyZPkyRSwANpwU8dgsOFXW5f9ODxOYLXwCY7l/oTeAHIY3
KMJFic0JDQnTOEbdWWRltOT/aGzuKBB89WS39Lc+ydZ9Xu5D7zxPx5kXOdra7Oo0
HO4xEVqSCz7LtCps1gZoim21uuqJgMgW1aTNigytXR35nNv0Ab5aVa9CFVgyN73G
iwe2ENvgmhYQcXyFCwc8xopBZNmHHsd+2vP/KaV4QhyjC+uPKgXfDWGaa7cIJA9j
XWnFNsMo4w+lLzbagYs9n5L4cpZhUu552zo5C5VYDJeyZaBIZjlYgVcAAvI1mXuF
mPQr7A2vn6WBc1RbaspTxZ47FuwVu7inuf7uP+XbsSPPn57yKvKLuEz6am8nfeqR
RMqnuigc7qWBG6aQPi76GbIX1yirTkdkEfQuC4r3CpVf6Ln2O/PePH2Hnm2H2pcj
QXtU+Fuhj/sPFJnHPuB6Yu5Rmcc8v7MMR1RibZ+2MlBVJOn0s1LjYBaBjOwQpDDm
nAYf740W2C7EpHoE8o5uHgU/RnsITwpNWJXPa1tqvEZq98WAM096VMGLGDgNSQsu
4dfrxszOYdDUzMaZSOvqWSPS/0OVe+nHBUqdLVvE51vpm03mHUltVWGyLT2/B/A/
HdVSIkg2w5eaG+MKwnGEkhHYxBbBAVqKQ4KsIhWwkWZkqJTkXjF/WlFlc8Ecu3eV
SqLLB8qlgncX+dYEUYsA1i8C4XIk+yME6u46VqVqOk4Kg9yAK1PeVU3iU/NPp5of
FF0VvKbKpo2XRf6OOTFaDZBQP3Fdlik2LaUdKPPsEdVVfXBGW7n2c3zW/rYqGJMY
+WorJ1XJ0/9erfRXVPztBtHrTsJ2x+rEml0L56+O07HrYyOMG2eWZNIisx+Edzr8
OYrGev90LEdSgABMjJpVe0vNuhTVO6ilda6OafpNbpbk8svL+8tTt7ej8eZHsUwo
6lVNfizmGoNxu3aHYdK17CRb8o2gS3ykzP7Sea8n2ZERvOX0gdXLpg9ObWo4/UV/
3h7vU0r0Cyo2YrTsxRH/W04IYetw7OEi262rEYWhtyARMUp1pn4TwqVr69pT1utV
nn3fEyOftM5Bg44KfN8JbRsG1Ti5cG0P6PBLebu+qsS4wbpTqA1R3s/1WmVa0fXt
G3d2X6k3U6so96v26wdvQJPEGMZ/d0dS6f1JA2RzxO2PJXjQiaaKPwrvojoRtMHP
97bhobOgvC4vlin/nOnB/1FJ5zCx0Fpf1Yq/8hAj92fVNnVDEMjHY0ULDroqaPEZ
dpM2Jpz6FTFVJDC4HHjn34jT6p9oPkJDsiMTdo8LyWSFn3Sx1Vrltb86arygK2m/
w/43LObgXcMJ6C5G55Anr3UUZ/+SOmfyZ/V+Gj49RPp9+b1K2QmziYp3HmiGAt1G
OpzYorZbR+lqIUbuNKX7JexXOUazlOIGd1SuPt2Gm/BSMpsFot33b7oVpdEe3osC
VlB1nYnlNsnBsb/BUlhHTSfjyq0F+wnQn1Kuxoq55TbpFDiTUJQcUPLa26bQqASU
Fym4UhofgIsFq5AeQNGWx51BujTFFvfufDAX3C98i6Q2d1HuJxdz4HGkubi4l+f0
LEzw7kwspVqOziTKNwljff6uV2kNT34Q8kYpvleihsHiWnJMNtMBuNO+lPZlMw/O
SxGKwpwpYOFasA4Hfpp1CqGCzfjP6pYsyGl8710c7lPtc63lVYlexlu5CHQD9Ccn
39Hdh2P2eHBUJHAJMdoLSGd2YiWnAp/LvDny5rzrq9ELbhXoyE+VKDmw8f1wiJOo
EjNF9akuRSmDOAku+kQgHbbLitqfQI81KRd5u/T2naY3BullyAWBncDq9yrLk4n5
Uy4AKfqSW+BvKFfsklwcUYHfZRbjrRISan6TOzy9NCRJCcQj9VqxmoUiEHpZqSph
YA7aN67Hrj8kq/S8EDkE6pgl9G2R4tdT2dMCZpFNlESfkc1qCB49Jf2K5PDnLRJz
0SR1CH/xvkDhL40WBobfOQRLG2LwmsGBp6dXTNX5VRn1BhywMJnXfx7zH+0daHhb
Wn+7zKi1JaoZSaPbjEUNpORXh5u1YollTaMqR6qFix556YzBNmZN9zvZpejojk4H
obKFxpXDKo5TfbQLVN3jQNwrBoUut8iknzONWzps1d6AvTBF/ut7yihLTBhH5C8+
y1R+7jCYVTVemCX9L0VXOLvGyPPqDI3bKD1JpR5HsCAmbPtYHV0A4cmsX8F9Zrcm
oat1ikrFivihju6G7sd/Y60n2gTsYvWAD/8lfUi22fvn1si917u6q5IWeMcEHn2f
+MGaTZHNsIfPnRIzRPUhlBEl4zucwNiAbQEnHCzUM1VVXHW0phgl4NQIrd9HaSLb
F0SETj1K9Mzr4YooJ73z0PBBjyOsgv+oQJMBMxftGDxt2wmLRlPrxQLI5xmzEkz8
o0mnM3LYuXOsenhWceGLJuqMZYLQM1YTAVWpKTCWeNE3XVvo84HCe1hMdhptJ9a4
voS4Yl66UEJdx9gy1WEUmoIeZUbkXuXEAKXmAAmIrb0RwPxcT1KHlyjRR8xyGAN3
V4YiyGQBG/mKUMDwOxISnqbZcWHZiSkb/ni5QygvSjOpF2BM0SoAd0faue0cGSAO
C5/3GWgiRH4RTbX1K0qmqs1bLUiWo6zG0c/PFELNdVwkcQm26mnQeFxwUYP8yfsC
razUU9EkQfQPA5aiaRuL1UPVmrN+PWSQ940OoKppQ69mbbp8B34tiFDPR6Df5+DU
s2HFAZN25RQGGGPJmDoKju0+BZTQ1sZHb2D3IjH+IoPEn5EmOkQ0SHg4xcU2fjs3
Fcf64YsOEvcewhJBxc4qstxkVRQeO5DIOCPZe7UekuSSMZgAZohcQi7r1S28sLnY
SLVXlkWkWEalwCvNBBbDjCm+ynLn2VvBn2BjzEeJORpUuuAsG5J6hW+0OqnLehbm
x0fLtsm4dkfRnE2ZdxwFmEcH8O2fb3U/ro2yPQrdPvqNAQVgObWCe52IBb1j4HU5
XURMl+asoWWbibIu4lgjNFCSAZBPqQRAzHTOeWnG8Lm8IqWMgo/p8Eoj8F30mDn9
jhceIvvtayxeX3FK1sAhvMXMG2KfDCDNJzUGS2yX+pN26/C1f4DQbzhD5l1AYxsg
SnqcWCIeEiLvAzIzDneOB88+HsQ0qljRAgyRjguiJfiPC562V+sRGqisMxxALpgV
OrKq/gGgCWvC5YUnha+49CdQ9WuLjO0xI/iTq9UpJzciCgK8JaPD5WejFbKSlncq
MJPE0dcWfhZwkzFLGIvet/SQUBBlQsOGbDapr/JenDmQ1rEkyrGwUszkg2RFBVEA
vYh2XYY4BiOeBMH4WyCWMJDHDezCDClIT8phfW0xgxq0CkMPoUjAyCjeG/69A5Z/
AiUoHo1LXB9/ZL5AZV7YfpzqBWCnRAFMxJ6TrkAV7jyMW+2G/HYoyE/B7vXTrzq4
f0nGdDaStH05mVYhxmubaf3rdm0e7ckC8z2adpE1552cRgZM1KYs/ygZnTzKThWq
a5Flv+04n3p3DNXVUkYUfJX46jfA3xO5Eibs1/LdVRJt6BpA67ijlbZQTrLo0pQ0
2ellmsq/gg0GFPLG+IvRKJWEvuM+nzc6wJ22Z9hBc0x3EE3H17n8/PSOblC03bKO
EwFdT++dEWSOv/o3Ywzt8sI/Aot7bgCK01hab08uUQofICgZyEQ5sbqZQmlExF3P
tYrKb/zNEvWMcv2Vzu2rIScwN1qIm1ce/MrJhFoZm8CrnXwUT1ofpfwxK6dI3MTP
V0tykVAXn+iq6Sgi4MPKEErO9RjHrUClpcDLV7N5G2Z8Vfd5ZJYqYOUEBtoxoIxc
JHos8pKUo5jQ71a7eW1h3TSp9IXv3T25YdGMEvIg/jSLEU/naM5+zZ06lHZRh1GM
5JEmoewX1G5RBsEngje4pqPId0ldWJIX5kk81Byy0VH61RWQe9E9we3pPGsa4BbQ
6rbZ+HPtU0ikoZ1nazQBYW37Z4oLDGfyoDwh4oVVm5r6tvF64dnNPxLjsnIlwdif
UFcaHe6WXQ7ep7sg8RVFWYB6D/d0h/jbGzYV+xbNlB6zq3qdt/n1pl5T2rmEtcaa
+wCQAcdkYvwNImPNUbEb+2HOZbnkJWjFGWaPdFCYwZxKZcqntHMmf6EhvnlGvf76
ORzKolT9MsDgmA76olnEx1ZmB3MAt5u0zEcCp9z9UHE+OXL1VOy9tmRnJpgk0aWU
ptN1dj2H7/g1gvF3c41YzoJThhRolnke846Tdy+Z7f6Gy4Xq7lKFbHNyhewqpl3M
S2clQkFjPPyA+7UA2gGGGJudDzOqgjIKMkCVNMsxlGtY1xtrun0pNBKHnfveLtCH
VI0ZuXohUqnDfQNy4D+kZ32nyTolpIvUCAoEBFpKLBADAhffkTXa/M7NMPTxeztG
ICib23hJCOKqlGVjs/VH/DA9UnhoVhZ/MxtDVbKgwWR7T9NvQH/LnLQq4qywh/W/
uCYOjzbEl5IeObPHWWA7FvsDtyyXQkZP0DAw+GTnUPeXziXVGET+TH2H8Dc5hUFf
onWMQ8l8SR3+1hXM3tnMzzCL+Bw8dYeLfYQ/LjXHuWU3t7KAuajpySEvUyuHPmKp
jdbn1xe83SkFRJYfNVOQ8QGG5tb16WQMyk5OrvN+2hlCFCiQzE2l7dD/EpwnVSFu
cRBomkJm8fHXPu3j9PhOBnb321syk39RfKMvcYy/Gw6GJTxRiGEqyra1ao31m3Nx
b3wZkudJUgHo1RWJMajSmPDao79OTeU1uitA0MqjsRsVtrj8Fwoy+82PTav9uquc
k6xnk6YE6NtFiEBQxqvWTO2EtQ3hfblTGjKoi2I2UkRmRpzIkCoMVdB4IlK0Z4JN
Jtr+VSRy07nuV6jbHKpGdDVNqu12hPi86W3565S19yRgCmjwy9H3hjy4eEjBbS6A
yrEOcvXmm6oP5GPUgBUOL00NswePZEs7EfvjyW1KJeuucrZhQpFB0ycYrm09CIv9
JkdaPV5bxTZjJ6vMui+bWJntgejDj73Odx9hiFst1VMwqBQ9dZ5UzGodIPNl9GgN
BFf1bG1/p3Aa491yYDfsKxNR1bglbCM5BAfRdAfBF695kEnlY0VivTCB02aC5g4j
qopV3gsvNPwZPDYxvNRU7Ppe9ZfMrfTVldNWP82GccrHZ68JwEjqXBm9az+AP0vZ
Dijd6nbs282ZPW5skcAB+uwD9ju2DEV2fXpnHdjOZ8Ign/umayvUwUzTU+14N+/l
KCd+GZNtWAPizSkpVU7o49p2Kmm3jqorcV868dqyPoYFp9iSt+PMalKjea2sPZOx
VbTAV1TDdIvXVaNZ5e/AZ4W1MlUz3nMM6jL3niToCAv8yEf652o8OEYCATubaBhk
dEHRdeNHNHJe6U9nyELrYRtm/GZmfsIT0Wb1cNJlfi4TgRNB5C8uqoIBSt6aIAoI
slV3OSPaaAOG3jlwwyeAFVe5doT4KSVExKRsPSWJKAWn2i2wSCZy39dxpcNyInrI
HdF8GAMHBv5tjX7C2S+WTRwrvjTZ7IHMwBg25CenyJWU85b26nzY34ALXLI06wR0
DUV/x46nsYYBITfYS1K+w8PU8JL7i7aR40/zyJAumtZ2SzmTavpUJcP0Qf4zuq8C
bOsgvUMTAPXhtkt/dU55cih4GTQIVm9E/i87C8cuBaGkjW03DAFKAYXXR7rjtZg1
VOA2lXDdEZIAQZturCNooKc75PeoanU6IhiQd+3Yqa0q1Vfv7mV70NWPP5j2g6NN
CfUcwnCyrtTw3P45Nt29+edLy6XFWwL3H9kVwYJU/i0Cz4AKhIwlmkOM6XVyR8Lp
Nr/zTUW4bTjsNnTHGjRk/HlRFqWtX0oR6k7kM2mTP9mT8zyJl1hMMf5DTGHmhGS5
Jky+bRMYOvSb1Z8YKTz7iWdLyIgtNaDhjJZ31hcyuUNZOdg2eYsv2a3PCznU7rDE
lxw9lCzp8TkBnR/UfTTzy6b01YR33E1uU13/KetL06U+06Bhq9A/AiWyojOY4kcD
C9z3wiEhvRNK/TZgsMJtvkUlrw33Ms1tc9ojSK+tnJY=
`protect end_protected