`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6048 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
wi+1jnavnbnCeZr/N19tUuyGkUR3oe6IyK/JehraDqRPz0l+fcD+tfxKkW5Zif7O
kr9Buplk+X/FklgY2b5yyLxM1HxcwtD5n1JCTeIS/QeY731V3PH3IVxW1QnV8O6u
NaUWK26feauHuok2q/MOYVmE3taw60r2Sz0rUFW3x9E4qLsoBH6Ia6chmMLrKTdR
3JXlfLpKypSG26VDlSVWBK4E5Znfkw8vEMgW+0IGJ0koxdRNKzdmyF1TcrbRqmQW
emPk4yZmaP4cXv3SFq1ISQSeiNk9Wzt/utcBJ4y7j+wCugj6sR0QG8ScEmAd0neM
NhRSCqg8d1ezsIEQ+vXeLL9c5dWxL05LhPwaqV21KcQUvzcHrcMPu5ta1kP/pboG
jhZX+Nb48/scZWjcqAXqLcIBUJYBxXh6ojLTLfoL9aeMSEpvLKaqtIp5k4XosVtU
m8Km0PVr6kvyMH20mwPRJQBFU95cDyPlTN8XwtL/NOAQwnyDwYm9TAEFRw5iSU8P
aijMsztlGTYvqXBBC3Wk0mdZhv2IDmQL8Ejw7gywX7zIJIEcqUP32kB4+sl1Tbz4
YgnLTkfBUCAql/dZpqtbpaC1hqH4zNgSfITvIXjQ+D6Zi9SUrbPiOTtC/xbyHLcI
FSE/rEtxgGj7zZ7lnPLGOEZJUlyCICirlNjj0Jn0wSsIArj9AZOWFJdzGnQdFhia
oTbK/4cxhPnVcv/gfxF1eKppb4ie8Et1xOYHajT6p0hZQaZKIulpRppN2GqL4Jzf
UTQHQkyIUpPQ5kHK3OT9xrFopl7pNS+40+FMW12EHq3llfZuwNb4tTXTXh3nU3bB
5cf3Iq+OS22Na3e6GePC+ZsufLHjZwlmlB1/hF88Fwz7h4xhDbR/HX2SmXHmVTNy
Zryl819ThGqyKcju3pAZF7uIllF/dXMXK5aU9E1BvveENhlt41d9z8D6/IwRONcG
5yR39GP+Rpm+VQ454laqlcE8m9Axa+IZvk73cVJejgxPn1U0huK7wy+Jciqpm62R
/vdA5rUN50I3fBRHXABRrTgpUZEjLOjafXSBovzSVd5bl571WXQicBHz1gInW3aN
Uo0go+5JsEdGuXgW5Dlm9ccVOruX5V7iqqdSvKfKyIOYUnl8ME1+Z420SrVHqtT5
Qb7aGvNjD4e7t0lL2mUUlmPUMsKX/HFcWY7vNYZtX3Sj3sqVpZLVLqAwc5eQX7K9
OnrmW2MOs/Cuv+A6S3jb/keCBOjlvBs7/A+mMV8AZ3iztmCKnIaJvmTJ5+IPPfgP
e2d3GtTCFYNlEsvQ5EUjrau6gtXcAkR5MwiV14RORfuw8PYrNLS2WFJECPR65+Yz
1oszerR97E7EdoUgbsw8DXG/9Lg2BxMPC4KI2zPJcqr+GlwoF+4xhoQaksOg3GQL
yYkkFkiN/VBadvqsogwhjLamaZIp6pBgrpafrAey0QUjrtW3TMqn9FRSk3VIFL/W
EjEzfSckhL0sH4NTJyhD/nstVBENos9/1lKX1h4d34S+9tMKBKTTurI0qloAspDa
nnf3cig9XqfVad+3wMAmCZA1I3gByIQ89/4fdVNp8u44jVjlD7naGFCJC/1o42Jt
h5L1ae6jhBOKi0jhsxy9u9gtFBTXZQ59uwMjt0j8IwkcGs3y8Ju4tjyNISdLxd+v
rIeyL0RmdGyyRExu0WMs00Enf5rWvcR2d8U1FEGJ/NXQh6ie02XOBn3/ii1yxbU/
atLfINF2E+1YzIPgoBHGnqR3WVh2xNRkRDwS8lpRKZsETTyWkF1y0XVU55nu8A7f
r2/ALV0qgakf+wtYyaKknRKB8uXZnauajzgdizXwixv4CTk4iVfDMoQlEPEb6Hv1
TyZCJBIH+wyjwlDvjk9mcut0MP3umTMAmaiVGYjelIjdaBOtC/y7ehAf/WGUjvjZ
XdsH0GdBvg+sG9pBrJvK/zrrEszKTpAI9qMtO+CRn5D2i15TuDWy/rzIMUCGpy7p
kJ67SFecvHOirhZ7YHq//BXR5nSDuNZhSKCgk76m0aeGQwA7UHDQ50Jcs8SgrXto
wJ4ceZJ3m4pvDEOxKeq5B8dKe9iJKaBBQak1/3SSpix1MSSw27Ma2lKiXrM7uGP9
8pBaF6cB5RzzF9FQJQagWOZpQgfaR5au3LzmUNHovLLh0Gw8hunnR6XX3DeyhZ9t
eVBG0txotTP0nMhI3seXSX/qn8nSSQ2DYREtB/tRHfLCZcNkhT6cuKMUTKKay7S3
P0FMJGcVdNj7tRh7Ep5FPSNxS9I6zehyLqEu11GXCp3d2aQyF8ukZMu2o+A2KN6p
zGbnBMKtIoiSxmFRN6MPrr5iQ3x5TEheMPa1NrfHgEjE4Tnvhdn4OzJgNhenPz+M
qZxViBHL0VstQ9KssxuQ6RSko1/vHl4JkoF9vbIFGN/p49WbpeQ1saP0inU1SAZ5
weAAUceUxwmCVJuPUz5i2ClmIHUCyv0VROna+O9KJPoGS/lnxBtG69eH6gE18kg9
jwEynbOjXSqiQcTUYxVym3gEOnFJ0l4/oGJqi7O7CKoKr2O0o4kZ41rsarLtafnD
PUvtLo8vUu2Mg9q8gfS4+AaX+CJZmwMhOMdCOLdYYH6H2D5dAkUr+/YgMl+py6D5
N6h9utnaldsXBC1bm5NL+0/bRMD9H32u97Rgax/vYXul5cBo/Si7Xp1cprS6h4fP
dxp6SWS12GhDqIGCGZwK4ZvgJvD7/f31fsgzGnNQIABABNvbIH5pS/YyQoszHI2N
sOpa6ue47fYipessaf4cUC5IQoImpLMtFz0Ks3ViAbGDUfpQsUPRvpn7jK6xxKsi
S18lO+47Deqz6Gj17eZtlSuP5C/mEWeEAvHYgNaTtQJkbkEbEqLcKl1KhqFJF86o
iycKpFg+1w/D5Cg4bE4+INmv+GMU0mWhdmPIlu83WlDVEipBOVi3sqE9WEQgEkML
ZhmhuNsYerIQ3RMRfQMGOUL8Y7WkZ7xKtYzvOinzlwhrK6AOdLG3lWARK1yE44/u
NojOBf+T8UJsw/Xyq3vLivsaoEa/CD2jyFPZsh4Cs7EXQ28yM031+8sqwPC5VMLL
2gHhYKpxqzpBCuTVJQIrRlB3PiiQjBSsv3NGbWLTwytxea8GMUo7yhm31nM0cN9l
piw4GyJrwYn4QDoD1inPqkmJCEyARbFulA9YfO5BZnbDaUIPCsPVQuqTIBALNQEu
y7bx1AhTvMkHatZkSKLRJt/LQUr0JZqR5I6akQ2RBiIxbSf27YaW/tQ13Uoh9lfS
2IAUGbO8XC0kIjunav4SK6Mb63Ql+/i22vglp4LJ/MHwOxXbjqaCC2mFJ3eHeBod
N9fSr/nVobR3s7XfTGdTrqEGhWj6+6vjeQIWzv6FCO95PvZAUDnSWeYZkomtHHCm
6UkoFKVKWFDik0du+jbudsfIYAZuaZG3H7Ntj4BPIDdGAtfJtgTa85eZ6Kfw/k8S
aaVK18KML+R4G8fRYDWlY5u9BaEmNx0F3wadiPrXbXmkrs/YjZnfA9iMmmw7mydN
EWlsV3rN9Qn9Il+Q8fcZGIFtkVJzYpQ3Ir3MeNSxm7E8ZhXD4VAKzD3wmTNZM/V+
yKazAcrfQW/V3HPgoDDhO3PPCMA65FZOs3QeIcnI/k57DPnxU2bPLTruuQiaRknk
HBAbW1tnT4im2Rae/RCT0kzx005LwqLL0yoKBo1dBjFpm1XqgJAOb6ZnEJgeCmAj
ZpJ4y1Jtf4h7ozI+zFJTdJjtjqVuGdcrv0VeTo4nTBZNSnGwPwYMB/iWg9uYPGbz
PqNMlg8yyq6d3AzqCf/R+u3PHtDiKGzyqYgmui+5UfvmQYecEfzKvXpHqZ+AVUa0
hx2rwRG+vOgHeLEYELEF8G79IRcffpN8zrGj5qPojWExOdQglKlPXUlePgvvLkGG
5eUNyilDgAM771cvagvicQyelR+CeH+vwI6EPUA3/Gtc4uXxa7dThgV7x/nUMthg
e39wBXZftx62wGFc0L5O4rki6msldLDAUsOivgk8azEvvqBYZsjc+DMapZWfTVUF
JPgsHT8i6HQ2I6K8AyUA7pyQ/Wvb2S/5Xhk1jS3S+EyFvsq/yhZc3wz/6fjE5ZwM
SkL8Tqh4eYRxDJeqBFCTxwCBy+1weNWZnKD/8qNBWU59ZCKXuut1veJd8wFkSiBF
orKO1G1BAZGOGJGYOPwpcDOcQBaRMUmPsASqaWonMPhLhQnEv/Kygu0K11/DxdjG
UdpQMgd//9EzEKLX7Yu+ElbN357PzDAgDid5b+svLbbDKSxQIEtWqFhfjcs1HKk7
IkljAVGdF6Jss0VFWKJ/3CvAiYPZ1YZ9Hetdwd7GL+BK46R7tbuqjeiediRr9BnN
KVwYoztu4Y7lCyehK9+RgZ5eixvyzqiClXbljxgLPHHqjbbrL1Y9jkhugfuALwAX
dIXnzr5GqgX43/fs8XorAoUVZsFelt9LpatW4OzN87NZtOViulBH8fZ/95IvM62a
Um4tg3/P51LR3GG5xpFMfJOLz2P4YDAgtDmWylT/0K0i0RgeXu7G1yCei8yXMTUw
PNUE4wPWDHG6L6np94UyQkY0/foUsDU7qqLXVr5bdJS2YG2vkuUXMsgenKdUpeby
RjQ5a43w7vso+bbe7bbkIA5Ti+di/FVOYY63du8W1/q1zK0EMctT6Ae1jngHMZjo
0zabAB1TctVbOhwBYGHhZFW7k9yTCzSggG161S0PD4pa/+W2tRaAeKom6UehTHy+
/aInJXTODgNs3q8WVs+ckoXBrng7Hxkvx7kCq57rTJ2V418j+GIEWyY3YwRpjYuW
zL1uP15MFO4tI8Ger7JTu4X7vLO1RCTdO0mUm6A7bK+XKwtqhezqwGoaAvLz4NU5
ZPgEJ3RefQ2e7rx72sN2zrZlXTLq4iVKeXNX6VB22T28ULq5m9tRWR1z/ptGGT47
Ty26CgerXTdnAmLPFEw1YCfms/VOuorlRKHYDe0nPjde4nOHq6++7HffFWLAAOUe
bUoTiKGWQNJQszoTHyp8NMyPc/ernRvBhdnE5lrJFveYuw95NDMDobx2ck8TpDZI
xmxWVwNb/VsdhmtRBeNpO2tbBQs6mogzCyro4p9mw+H74K4gTDlMGy5QU8R9sgd0
hxi4NOidxJ8eF8+z207MKCkT9gp627icITYJSIUY2EHTGOPqAAswe1f61W9odTbD
ebIxe0NBDm10ABEmSoJHnX+bJIRKf0hUzbzthxlPLKelpHOjrwOm1ppyT2XpwsHa
PH1mrLKjBGm6imf5cv0UzkSJe4+mtiy3jjONwJnREUjDQRZ2F9x2nlJCRchqT/GX
GnP6+34kO9kEXIWPwGfpa9Kq0AuyqUOKA+jVZMBbKHl1tou09ZiHu3ZwrbQ/PAEQ
3mmNKdS0qoINo8qRTUUdqRA9mLcD1ifuH7xMMxJKvct/gV5sK+tBA/HKiRv3lcxg
FR/g3zhwLxUpF6jLODizcq2yYE8rFtvhqHGk9N/Q7SN6JMg2T/pK6/YFWQ0rIr9A
oYoxdY+RweZqw4O0+EF1Teuo5pcZjm05hR01TIYRXK9kPvdDY5YjAmJNL5xYGLsz
sAWM8WAPSowOeHEpw38fDXaQ7UEFI1fTZKc4t/Ki83yMQXU0oqLSyy/3eUSMKOx4
dFnf7NdPN78E8gtUlFzTZIkN4wacs2Vd0KXVARYx+lkEK4QYva5QpdP4Wb484Bfw
bjfQLOitvvs3Fc1MEKlGL5onvo52ZtWoEI5Hc0BgWPr0hrOhZlLqGWkoqMvwAJtr
pcJyJZTnJ7fWSVwKekV7hPpE358+IQnefG1wZCWhMQQjPlyxkWt0Eg9AQqeDF/Zk
TGtSI50+DWfi42AFT0FAvh/ifW/8auT0s4DI4ItMh12O2Il6CxfmIptu7MhILQcS
VyROKPr3YSgG8VH45mHHLkgkTbHfEV1+kcO8rkbfSHh9hID2p/E9tlp0YfWCJyo/
rk7fFNobY9/M0VoiPbZDaWkZRtWbzxFw7R5o/HpfwU0lsLrIg/ZpgOdm+ln8VUPD
qwVIQOLUtOmJOEqeaaX8ap/NHxvsmeTOmwzSP/1sU7ezr/UYkb/Rp1Dbfkj2+j8F
0HgRX6M0vGPbQI3NDfpeqyu3Y3TepoPQUREXWdfBqVK28ttQQapUQfS9M3nY12UK
zsyhFzeb1irkNuhQh93VI9zafABjg84jOfCKNiaTgT1bqyK5zkz8851h9UxoLttk
ENQqU/NSvkfoCX2/eIPO4TcF95q/4rCrFRppmvS1XwbbLjr2aqzFZ4tw5aoAI+oP
+tuFbSKcr7NRSIvqVhFtjjUY83Hi5D2aWKpsxCJB8RipQ/9XtVAe41Glgsbv3ejy
JMV1mx39nJSBxP8Mppac9H/BHowvVeeVufLMxA0HOF1jkUdhbahD8eNBhGyxAaX8
KVxH52wYAvWdvBehiE5SsIxZ1Uv7L4hSkPFdVeSC2NbPkc6WSVNM9D1o+P7+20Tb
fPJ+igR2humsMSZyb+mU7qSeMY+AooIdcJRE4c4MlmjdUbONpt6J0jyKdtrgi68z
IGTSwczaBcs4xdAPHJyeiu6BgtCT0ahaG0MbWhqrxratoF5ZaHUC1/qhAp8gj9K9
CXiddVMYTVZM6RRNos8ZXZZoPgz6bgvF5OwwBOoUauoPJhoGKtOPDwb5eL9CvuqK
FdDI1DgFdlF+q2AkWjMmpcnLLLBMiykXVAREHE/cSDkva8BJNC0wzwWUFMvIhet1
I04NHZ+/x4MEz8fV1n1JcqIH2wNfErOThOox4pfJ/I+Ax1SYEmF0Vdcq3Yx9YYj8
6yRXAHIIvilxnQcczo0S+ji4+ZzW81mtYQUa4OUY6LAhIsm1Czt4FQ5HjOgYpV5n
D5+yiEBKpo/4hCGjuBGl3AYjlV/5M1wLTTP9i36eXFd+TktKgx2Q+lq5ihS6vgX7
PblRSESJdRz0AdCMeXMYrDuzWPE3HrA1mFAYAaDhX6XmDAIdc18VEiptPPqyjVj6
aqL5HG8qScw7i3DBkHMlNHF/u6zzMnGBghRH5vxbFSQoJNzkoC8dhBx1xGWQj2tJ
+PqFmg10cKa3KOl54K1e2PAWHMCseqeDj+lpa1mt4SE+m6KVzjoGyP1jAo9dUZO2
bVJD0kIYGbXSCzioCetgOlIfDU9bIvA+7/BC/AufJ16bTCbaUs0jbqxRAnvXNnoy
SJZHy1J32KH+O+kkIGTWhBYTgTP/6fmndhuGkfYQNDZvKxb4TwR2INFJjIIFyUqC
tn7M4Ws1g58Guqb/dmfbsjCpCnXmAY5vAer9U2GRcZVQHwdG7LuYTNvSIyVIcWpk
l+g149FtfhXGbrro/ot0nyUSG/R7Fc7iMR2dRH0/KOhNV6MF3EWY8a9+VzxGc7Yb
xp5agO3zop/H7OfnNQqoDD62/izvIqdMc7XFa7eTJvhDKrYUfc3drGJP9cxNFlLv
L+UQvM7FtoAsQZzr5/x2Mp3HAF6ujmXwGiv1RuE7lcZ1FCEnA7jOPb27FmV6RfiX
Mn+gRa8xD/qzh7QkX6KI4YNgRyRBZX1VbXgNqpsf7zXvg2NCFcxforJOFBEDjWHK
FJMRbjkmfYVDRUEYOEyqhXnaWWL8oj2gnNvqNte/D5/xeTkPD7hS3KpVq1s9JfKn
zBdaSKK7nhBcSu82+Rd17n3/tIwbxGl8x6jnluOz/t18Wa705YlCI6aLWAZ+OMRH
5xcSZXN63wtjN0iMFAnxAyEEDDZvDN+MKNMNzv2EP41xTK0yvKiYQG25xhZ33pP0
XjKDyslToFzTw1m5IT70XTcD15f4sxeGI5V2O+WFBudyH1/482fXtamcQ2haGK/8
iwWAsQw1ROicjT3ODIKVq+3IbXBEyyP7SAWvw+4EF/jD36Z2IDet+sIn2pJxNzOs
AEwrVXc0M7+wXoP68AzESTJVExsnve773DSS0RSY+KlvDkmagjG1V7qe2pv4ONP2
`protect end_protected