`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2048 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
XKfcKMLWLY4TfubABeEmfqhUJojlGPVKToLETH2dxHjJ7GM5uu09n24de++zV//r
uTRw/kchxZ4G2F8cE7pAOWaidx0I/xR68LlwGdf3SGYubWXtFblwx2K3K0Q+tSnf
qYcz2FF36fMptNuuAyN0YSeCdScVDHDzsBUazpZE815+1fmj95UvuTDXXT0pQYn6
HwVmx7P/ekiUm096OMrNK+durZ+/JVRAXCzhA9fxXyxX23LCs5kWfVOKAGpC2lXe
sMzgznqsbvtCtjlgztY9HKBtgFWE0dTKC1aR1MLL8kMhQGqCPmg0+EqMLXegHOD/
dQPTHRRvdncwG+ZU2eASoHumZDgWAlJF1TifL0I1xwxOXGwdcNIABvS+DBupXxVf
M0c+21EfdXnqxqy8iKEWasbiH+0uZMzymuamCwm65iGAoZDnmaJbETXeutX2R5S+
ES3Ky26X11YBvUpPZnB6SL1eHdn8teg3PAz1du+9Go/o7Q5DyhutsMyPafwd9L9z
zHDq1AKny/r44vj5B8uLNeTCMvl5C69wbaBy32Cq4su2TQgFXV6KbiMMsH4kPx2j
Xszfk1m/dEV4kyNhb7P0ZPe/sTszuU7ESl20N9DckXC34G5Pu8klxjvmjpIx0FF/
m+8YHlmG8WwKx9bJ4/o3E9RH1Kg/jysrdJIjwyISvTawGOYmOh3RPuEJRxiC0fIr
msPdsfW3flBOvS6pxWG4ObXHSNkwFNAUta8t6dCU6nuKk8sVtBD7dL8otD71M6ad
PAFTBsKJBgbfRU2Rk0Y9hDdOhcvwI/v1Biswq1B8chvHvB3KcXrYNNCDf6kjpPNb
ZL1amkSBa7x4Ji/pECZH5u4sWuk7qkJH4xDJfJCZPx0e5XJZcYORf3mdqfatPBCe
d+b4SuNpWC11Myq4vm7tO+r00sLL0uSplvoq4vs5z65/0vi1cAPDwQny2YA0Izvj
x+wNK0MS6YWsBCfm5Maxu3gZ7zVxP0y+HpmSzSGaSh91s+NlGVfvSYCKZvTzuHrt
HRdSn1InZbsdWC3AyFL/E9DEuGwLKwtEZcd/FZVNa8YJpO4l/yC1FCUZeLjRsAFO
4cxywuXOuwFxP0n2R6/SKrXLtL4jCno6pC50bILReqBRsx8P9zLmDKHdVNFM2g4Z
2L0s9rQYC6LjNYabnxoTYsp0EvMmpA7DRi1PVWSDfMypHn/oSgJHJy+on5FvTHkj
RcPogbJWo8dl9lc7BqJC1QefUIfPN6s0/KsrO69zEZb3nWz87Sjxz+ag6+5KfWjk
gqlerx6E7q9o28qMEyB2pAhYjgqaE18RtLLjSmTvcJEHxglYlQ+a/FzFghjfRGsZ
xItDOqBvZ7DPOf1UwkfD3Ifi64LESzBqyc1EdiWqlX0I2DI2tymwhlIyfDN1s7wW
QdremxjXuExHHg+Ha3f2k1gGXv8rg2Ft8X8ueLSQJdJnGG9qgQcB+Nf00SxR8KAx
DWBJrvlD34aj27P51C8SSVMfEwoaMyuBem3uqGfV3JYAZJIPYx2F0kW6wwUh1/fc
YEd+T1rQoclsYFE+gzGpE/DOT6jG5U3ZkNCV7G/+4oQWQYa7M4dRotW/Ss6DMHjw
/RyyuyZC/7LycQE35ftqAesulfIzxEtg7dYkmfu29lFSmk8FIJf3YMDLBetlzCZR
+4VIt9IUj/LMIIqSgurvdPQvOELNlfc2WsJwgo1xz9g8GAKgoVSyhXJzn3jXS4PR
1j5Ko1EmzJohngywqPQv6Hi/rhPmc4qXDinPYJ70krxXWpJAZEfGlb6YbWzVhN5u
F4jaChXg3fggK5fVBq48ivXgzp/MW8taBthRhBL6jwZcWMMjtgHb2Hg9iOYguupL
FPCxxwiqTvYKI5KFcsC5Ha/Yog3HUI14x+B3OZ9YHrItr1wPrUbUvUoN9prYQS9/
wJPvpOS3Tcgo4vJkEQLN7Pt5Fl5Eg16DGQLyPqpf42UJrMdgjmAR1AeVjZbRLjnw
SQynr30cSgJVDmD9bbNJHOVp8g3H8Eim659kNoSNCbp1sQj7QbYzBdQPhUv2569J
CXoXldL5UUDv2o/9l/qRxoW/b1vDXDDWgfjW2Go4uTMA/sx80MoWj1jRc0Bv7j10
gFkHzC/GiSU6BpQXk0BBsqi2/jKKpZ5PsFIQQLsuhUba0ADGXxnxPhSAj12N8ZSy
7gxU3uNGisUTUxWHwVzl2jsH2Dx7rtiBxUR7l37xwja5HVRfFx8nUpfFP29IxAJJ
fM8xQPq2IjRM6kNK070HrdA/CTb0uvGlrMryVILdrH20h5MyDCjmuy0Jb/hjJqTC
hCzERBu4AiWlUFfwiXk8wG9Aw4zAIjjcE7xaZ/2STC9cto24ebDh1dKH4DzdVwV9
n7+d2Oqw8nOez4Z5hgSYL/89pl3XOXlfgVgPHT0Kx0mrQ/Gfnkg6wxvlkrTo6s5x
JUiv66mvMTGfQw5uUMN07Dka29GgBZyhJbDK8ROZGf3ldqBJk2nzOzFO7ReAsTsM
W0FLg8wUGIrEO5aUDHscGsmj+WSIh35yGd7OVr5oWRegal/E5Os6C/4onFy1o0Gk
F62tGHccBBr5/vZZ2Ed3Subnq6GDR/dfKvu9EJhOBHg=
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2048 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
8aCqQ2oUxf3QHZjuYP1t5PlLWqhUGxzWKTeFtW/SNHy840Kyjqb+kPqidgHCoXX9
Bo9wl1YiL6lPumNznghJ9c62AZd2mTDWx1Pji4vrDM1iZJfBr/rvk82Vu67anXjD
356jS7yOE5F3xOOtg0FNDYiP98cOEzRt6Hx/BhQTfdG0xEotndvubRi/t/eRTOMp
QKR4yje356uyNPBjEGm45AMQHIWUv0TARY2u0qu1OHFla4RimJIxUtz91rU+2XR0
s8pAphoFw1isHFOohLWIiO3neH08ddsBKHiCQIEKzDALVJ8kyWZRMoWoFJVrGrmr
aEfekbdQvFYgrPgR2RrMmTvLC8YH6AuRQLhy9EIvl7Fxugo/oxza3VtEPD7PMY+2
qvoFN9a8425h+4WgbW0D1Zi62m6px24Axz7cRJmJXWdJmMJJNbnYB1DxdCTUNsjA
hKn4FS8PfQPFS9rTEQ2wtBltF5ygGyJdcZRTwv6TmVo0nZST1tmP8lcDvuS7S+gq
4jz0O33xc1RGpmkbBjVNgqlB1dENRKBI5rlhoWPpWkS5EbtxX8blyHqPIzywuIPU
6XZjVLqPZh4E6dKy1s1ydYnn+qqcMcFAzmOiK7wzJCD+/wQsevC5vTFcZ7Tnja2p
n038J11FDr5FUhAC4ptMXOxeknB6auvCcfACw+y5ZzDD16wHBHVMcqvdBpygvfyo
lTNtj4ofCVgFZSTSwf9j37ohdCKtChF7zVZuTBOFaUX6nj+3lC63opgSrht9NXwa
XHYKpM8B6X+cofM1U9IKZIU8HOG+B8IngQyJ81kbojQRdjEcu4SEG88LdA5fhoCP
KssE7pokX/nhVkyikBxoW/ouk0zsUXElmoxEgnBSsTBWWuAHkWBQ1y1haBI1rCY/
/vvtJAhzfyN80jWEeFFtzcvsVjJGld7/38kvIoQ5LMvkl38Rxue6dMe4aniiGkzm
WxsZ98SUMFHnyzTl7EzCVMXYPndQfZC6CApRaaBQOpFS1DJrdkCtZlgezvwzdktU
yX1a93thbgMwcP7JMDvQ7aS/RtkvVxl/NCKYWvTLO02VUZugP52sxOoqJpf5EXaB
YFEHd1mwZraydbyNKqdy0T3Fm0HvHTDetTdvIv+X1PS/5IX6Z1rMCg0TuG7ND63p
dWOQrs0ZYi/a6nmtwh/YUPc2th4+TCkyuAPsy7cdgLI5MAKtKTeVsAkjyAIJpSyY
UA71v3nYWLezTS/oMMG324ofdXoYCdaEl5ldNdInqPiEZKQBn6MzQmHfdcC/8a+H
gP9ad28rg8pG9Z5LS9pLP/qHiI8VLNU4vGzwisSppu1XP6bIQlyp0IEEvB1MSS3P
MZ4RoWXby46GYl3N8dWdtM2mjoT41ggrI7J8shSCGj9niAHpcFXlWkJ6g3gHLsbo
UJr4qR9YbOiE3WEjbM9wFjNv5yys2e6gfFIg43ZDdyb6JMX9BMkn42L8+YZ3tAKB
ITXxdTmEFM/PsSGCYSUDgA8fQQIdjtCYUUtcuvBzEcRm+CqqjeZH2iEq2noXPRSr
QirdGhFJCGEdxTpUfoPbXWfRdQpXDGsxJ1FBQIhWNebIn8426XBwHxdPoREdQEEw
yn0SlgCE+SkT00wjBNRjCP14FSM1u5rTFmyJ210EQQJYHD7SgFP6QNXPI0kCGO4L
w8YJ5R+Z8urqhfOQyKH1Iio2gx/AnYnDtWHcgBNa+hw2X3G4/iNdbHECXej2EjKX
D40KTD53p3Uw41WQ+bHx5njuiUXSJ83m4527HAK9ascPEvsRI9uGDbeuhlpyv86Q
+jNwEhdmDeI3WpoggAvxbRn5kMhNhnoABI78Ox/VSC9qH+VUyQ/v3EOOguGMauet
UxmL6qRDrV7nTxGFr3r/+YJ3HpJTwZCGOfZy8JM2sw6cUkoFouOOQZPMnKe8UmEm
9RG9JKsOayowqOdtNsEEY3PERdGfyDlGxhqzj4dyVKpOUZDjv1Wgc8X4wKZmDivj
ftjfEj/SV4ED0kWnOcIfFg64bXSe/Dytd9DrNp7+O2yTF/AOLGPfoCBzQSZjXfWP
sl0tC7nrB7fvHqEOzZ9yAnncm31KD4ivIUEl9/QByXqxHKdI/Dt3kmLtfyxsSDRR
Zw5mfNlKtNcuTBTGq9vncaqgymK63eIglX8k7eNIkuFsXUADjaUBADLGAR6gxOGM
GugunzYcV3gbLmtN4VMaQdSrnTgNHVpLGNwdw1/NGaIiZ8XKO9ajwR0T8l5fue4f
45gXJzZwmrigHUukgJjsUR8Nd7qdvRnlS0ERqO6QoqshQ0qgVdrLKrhljRP0IhNa
pAZgb/s1q3q8Oe3om3hlaSOmHmnhER3iL49N6w3RZF61ntjbosa0J6QRtE8yR+xi
EitgMPjJy86V7kTE0gSQuto6HxYn8YQC6eW3Jl+Cvmpi7tqBSzM4Zdxdwuu7JaUF
BGs2V0S3UKYk2hOrU8mXVxta5eklDM6HbX/DxKke1rir3apDs85zRARXSAh1elcP
y4+IWRA8OrHcnkQI4aSkGAOomJ35M2mwnGH9oDecKMzvs40WhAdOlVIm0uX/Ja9r
m4atlAqIaclTC2EVNawF5El5OelDWgkMrEtVV/7S/iY=
>>>>>>> main
`protect end_protected