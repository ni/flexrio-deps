`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 61520 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
VKWNRQF+vfUNEEp7apOJOQf/UlabpmNZTJNZwgpTcLKd2EvkABc0iQQuM6nlKONr
eSFEgEtZeD8uVo1tk20jifMMf1O9EV5ZfPWQKL+4mQA2VCOIRIVN1+wn5oBXXIWB
yqblKGqJDofwlVKD/jQ9mDIevaACnlAIgy4UcO6+rV2VCkrQp0hZs55HpJ9cXHBB
eB8j7ZZlcSo3WTikmpsCeCEr9pn6J3WpnFvletfhMMj48qcwVn3H8jereaFw0rpU
lwy91IZIxy5LycXNpn79tVVhjK27atLEkwvkWIujORguNtaFIYTR2QE8z35ZyKPp
3UC/P+UwjmJMFrJ03HRD9uKPmsAIDLKW5+s2KaBy7+hFzvWS9nEZCpZeqjfyt+/+
B9PBrDu4gAPBTaa/BU/CwaKyb5PJ7VmFKzYuo81lH+8ur/axdvxLj1Yx96GyHFdV
QgpQrgjuE6FHECAJgdN4NSGoMQRjI0/uKuyF9HkNBWFimjyoajVYG4fcUAfNT99H
emooVR4BZlDykUw7mEUpqVcj7MhK0Zyv8Bjfe4qXBWhQbnIs3C2enSOAzMYATqpd
hYkjUrvfT6fC/CKC74DNQhHTVHP0/Too1QYSkC5KtgvwyJ85C/NNjThponTYcXBC
629APtAHyzl8yX89ZNoIspamWXGeVzV0hdc7kDqFO5/pRF5o4N7yT9sUtKHgSIAY
S34zeKXm8mRfG+NEzarMKCjBWYoF45LbxNzKA3FkK9QdebTCBszVTNTOUQqDvWBt
VZEgt73UqaY2dyspQ/dIhpWCzxKvNfPNoMcpea+7VWhInqsFA5nnOfF/Wq/iPjZi
UVudgBgpmywdxH3bDxVBCQb3JuNO/V8VRy/7N11cDnRcZeGH2eq/dOF7oU3xqZlg
rb9gO3AcviyiZ2gRVu/x2xzwPBv2f4OE+iICQqRcEgDPOpi8ExDS67ZaetXauZ/m
XDEZ0X9YpdZ8RemmBBiUKj0ab02ADXWa47MYLzzbPxMTEoJ0eo186zAl7vgmW6zb
h6YYJuoHnHw1nUucl84Q+k+UyxEh8iXqOvtdquC7iszljNdcu0OWDauYDLzDQDjO
WmGtkUObaLbbQzonxK2TCoJlRmVg5Opm68/q4WepLiJ2WupX4UZztKtmCaFbetq8
EQJT9bXOH+zZ+dGFgWi21hsUevbZx5rSDvNcO/UELqireza36qG4+EFbgUEh7M/2
Huj7mAks8L3VPzG219vkU+EsQsRkajxRuHo8JQELl5N+dThTi1ymi0CS4MaMa0Ak
1yui4Mb5jTJRRLLBW8JglF4E/jNJsxyJ8NHhAbey6gmL6rENhTxIDwi89i0JJngp
1G/9N27Sf8ID9c+s/VM1hib7o6Z9vcOEJmNfUHYcC+tkhh4j6QYSXNS6zfpv9R3D
kGqIiOFMwnbo8gNFxxjSLstbXerZBh3a+dUEFKZi7sPrh0hHyYQHqlA9Byp3SF4s
0AS7iGVPzlAnYKZRqbRMg/DxH6h5RTK6udsS7d2PGnc1ESVhoSeozCxDIIxp8zik
Qszv7yBgCrCaZ9u+4v3yIT2jFnRFmTsw8hSp4ebljcTlVHU2UXFF09TtR0mNW2Qu
p3VgG83dsQ29HyXvylAJxFuA7vmYbc69ol9ztMtMAfXlloPfKwVFtXUzvqgmNvZ8
66ODt/I0q8CSwQyEyLl4KdN4t/Fa7mKOHwu7xlfhZmT3NWphMeaSuJKozUpRd4Yo
lEzJs7MWa6ZEPucolBCblZkT5fS1ZpgU68bKZ3+3P3fL/K5d14O50p6KhSPqL4KA
ycOXwn0a5QhwoET2B2ytaDc9CB+bhoajbLgXKsizlW9mViX76XFoixUE52GowRFh
eyRiN+17N5jzNXTvn0eJFlpRYgKhuBVFvKenblIZVmwXTUD9Osvw45nnr5qJTnaD
5mDDJpHlV4ZUXx4CDGIBsaNcjb9KE84fs6PylIQxZh6CMBdpmcCcPVvUAx6y6XyQ
B45YQXhBmXpaeDQMSk40TdzmqBFWQEjXTTtiZ/mx2B2evHMVSr1Tu8CvQKGpZ3rS
Y5SSIv73mMgLHo2Ysf5nih1BrjfLdTO7z9dnQifODygfiSuLteJtA+yFC1CBAFZN
4CC103pEd3QrMRFSJfqkCfhSt+DojXH0zzIzvlqEyA5dIgpJem0Qx9RfJXfwlZNx
nFyRLAiU64doWL66kpnWq5TqY6FDfdFhBACYJ7LeG5jtPAMQwAAynQiQmYlnW3Sq
/mrM7BGnnfONVeda6yyVc+I3zSUUQx35c+iUxuMfHxqlGJV/xPoPp0z1Ed3+aExd
4092vVyDa7brTjt4ly4ywBjF80jMQ+/ZtZr5a/d/Ku2DADozoO1VazDBg5uB5AMt
hDRI8S2MTIf/6CN585lgx/EuZdTIiYWKxAs1gS5JhhBr26ogqCSw6B2x3QPpe9hL
TCM7GQ7HFxG/Ck516idbXNEfOt6RUtoSUqyQQEd2OntEuu2CTr9iMEHhTj5SToRs
OF4e+jpRgPPd756gDeebVHWw3V6k4gzOr7NU6gzHKcNgRMrBfW3TQlLN6GAF+NtT
JUspTGxgLMFOLErz1P+atRBhtygoxmZCVOxgPs4NekN1raASs9JCPlqZS3s7ZWme
2g2TH6Y/B+TF6OBQlDIRMKY7Sv6jl/Znr55vY/TXOPjnFE601gpAb1CevnUxCuSu
oMLnD6bnA3DWoNTwnxKG2QVYDWtVzV1Beqi14CFNuZdoMA/1jMpdiY+GeTyhJuPV
o42gFgSfchtKfjTlaSr3hcpuVxNCOC1Hx3nQwE2RQr28YMTENlvlivVv0KQYO3E5
fl2o2eBZOD/f+z5UMMKlyjV8asOS5Fi6s7e9UOljcbCz/+ObRTt+ks6N0JuieLgz
l0tCYDnZb70rE5shJL32reglNJt3oFf5l7gj1R9s9m7mjCYImiyxiJ/MsXRfA9A3
AI4PomEWTPPRF5zMBFRoGtvIdmrWtBKF9U1ugKVcefM2Z3MRse5c7R1uU4p7b+da
TP+hGsp9sqjOw63UDDyex8+ATncZ9OnIdX6ZUy+Xq9o3pU6yDz7o4ceNSeweX79y
WKbmeTy0pu2CNeSrUnzRBWeuc9XKrA+bwqZ0glIK5/dk2WKN9pnosjow35xks+Jp
IhVO9G7h0ObT8X2CMn+fA5WNPqmCNlXKTafcqyxQp23RqUeXst4TjHuarzl4rFHL
ys8Ta2MEYVYuzO42oERSr/crst1wXsnMoB66wgBbJZRBPHtm2lon0MvgK/1aBRJ6
iHn0aN2V+rqa6FW5Rwz0KODzwhyzOtaOI+w5Nq+678B9ZjeWdktj6sPzwE1QryPv
HLcvxg23qf+mF984NqA0Z3lAQmOmUncdKITtugEEDlHXLmT394A8GFYBT0Oy6wKF
NqRLxwrJ1Yhwtp7Xflii6cZpophXEGDWgHJzeh5EiiuN1WA99i/Teyu3084sL/jx
BDMbB7kvp7aNXvVILiBmedgeNjNSVBUDuiwUsRQuvGuQi5Pr0801GDfhVpI3K4In
KcMUo3UL+efoXpl7xrRfgoeRjIsoxyKf25JpGFVIXpBAEwQIJGS5HNPv7the/RnS
sQRV3EBazCYqhedZu97zdnPXwauFIdXeFEmd2U8Ej0Ge5bdwM+nlP1vOuDGFYecb
61vhkkGP9i99DZYIwnSbVDXQpsEaJ0C8XKuaK0nLWYFUfWXJ1wfB+CFeVRdF/Mjb
06tfyJoghnDUfybVLboXVr/d4O6jDJUarU6nmXjZOgepgCBaGIv1E/uB2YhT8HZ3
7F2NVlcNNtKIuClfa9BpV++YAccO352hgSVA3VBBUiwjBw5uu04Xtml7txak121Y
3xWSqSaPQLVPCTYzLFbDEiSChaphIU1U5kE4dUUZRtObEJDxONUCnKebw6kcJhaO
h69I6iqm11hybqBuGsRU21QqzNS0OxGzIZBg+Bnk+VcGxEzTnKq+PkQGLkzr6T28
7LCPHbfM4Omp1vv7+tWULmehp4oyPlU1DtrZB1L5kt0unUGupEs7JupgeSS37Ww8
1bh79S9CTaCs0VM8Gh+aqF/tABdB/C7wTb9AdjrXW65C2zfvJgzmZyszyJ7nhk7D
6mgMBfm3J4x9H7rMB4pIsrF57OI1Q8IZX46ze2jy9V/bwclBh4Z/N38pxaT+u4hJ
gSnf/zdOGjheQET+99ip29ueyqRjKA0+MaXsDmYCZVwFkXhQkojyE4omyjVJNV0t
JfFa9QoLHVM4f/yMkZ5aVuIQ/ybKiTlOoN0F6sIhLnoQj4FI46sNiXhCiOeMNaRU
dP1FryfqLBZIZ3/AAU0LFyI/jN74+5tpvpBHHFoIZoUXcctOJY9DIcawbY+gf9DL
jezXA+d+RtukOQJ/H3Ax+bct+98JOtr4ch7Nc1tpKNK0EMQf/QVaebqvyhM+rraE
8AonBMG1UQOccCc6RbvTXwZOdnFxjy3gtIcqE6GIdUn2OHJRCKl3pfVims/T8rOT
AYTEPMkaynf1Lw37hU+AoqirXWr0b3USYFxC5s3IXUbxrs/FoK26j75095CpNQ6+
8gDsriYaslMPmosBldvNr822CTU1KUN/tteatpKqJAxThJlxV2LC5aK6E54Xe4qF
xDkLxgvl5ls7zoT6nBzr8Ll2ZwvhtwNy9/q4Jb19aVtsSNcmPlnfxF6N7b8pnkVX
v6SzXpjgd3a/MH9EZbaOPI77fngsO1Ockv600LkiiMyvhwuLOPNEkDd4vanUTixT
CL93Ky3+Bq6P0JoUNtCkRPThQsNnMytR8NhwYHN0knLZwQzRwNYQv+t2CFX4EDR9
oYJuKn6WU8ZBAmz8wVFuhE6E2MKZRFL2FZ5eIpMqIhL7a1DugRnkcQsOPunhxaH3
/wGUaoyDJLq8O85wfZTFcIGuN9inRga6w0vvOHKvj/xbCe7+kj2bz+LehPMyNsdJ
PbCzAiveU2GVn9QF0qA58dQ601CYomWbTvtlDZsiCVtWa0Ya5HytW6IXrrAhPI1G
gID9JIgAWA2wx7coh+LbEEPc0dyl8NOCDXUhG6sYoZv0wrXAU8a60wtHtx6mene/
XNlNEuoxLWLPuY3pkdytZ7XKnqyTNrn/YJGFc3HcJJ6vSacFUTr0wgxmWIZPHruk
YHl00W8IB1O3kaLmwmSnq9w/09SkJyzD5PDFxjHWZIVpM5OHajv5Q72CX4xSYVeJ
UUQA7ks5aqrZDode7B+TCFGSQodll/KwWWn77ySylKmV/1036xDI26knIwDcy9sb
9LpEsvH3WV53ylsOKw9W4OMrNTom7fRADMHyRDxythiQ6CLrGd+Y2vPFT74Z0IHh
QPcMfy//uqVjkflXIpuFW+RbxPe2Z4RMKEMsTejE6LCx41bg3OHw/pdHHp3IHmm1
15zJqGbayFRr7T9CMTH/MWOIOK3lKFPMUWId67kGRRSTqaEv8E2BkSx1EOkjA0fc
v+28QZQ1Gt0lQkF7q/TL5tBrpluGcEfdmAEb1/BCJhiJJN23p2zLiRjFiUlvbWwM
lC+TLE/A4wW1N3dZraZ+6aZHfY9mBr/gqcft9UveT6dNAbzrm65MHCiulJL069qd
fvp4qXNJ1GpMBwIlqDkDHxBmolTKdYIEg7BDFH4FPE7HPZqk5AVGKvFxZiS3Z7ZO
Y3By5zLMM0M81+JISFpbWsx/3OpL7+wYf4mFeIZiKOqYlHY6rDmU2bxS1lCSjkAW
ObE4PT9W8d9SMNzKBfpLZKpDXNLb0CPyRcHMOpGnotgC4qlVRTWJkGsRsy/MClaJ
3krPQZA/qQB7ntxdqI5rn3RX1ViTb2BWmQkkW5KQH0bKt2NP/bT8KB2GNZb0VcIl
H9XJPq8v2sQQ4Cyi5AJ+V6G2z/Gy6eXtjxXjf3eicaV+znjMzub+5RSdJyLLTsQm
fuytTuyMc2843kXHbjy8LjtwKe8eedhY37ckBwIhA2Ti+6P1xFiT3kCj0ppUrafR
tow9NNzZrXKFgJsvLmaLzvkh7xvqtKEHNsYB5JyTlpk2ent4sB2ztt4RR/vgavpn
tc2EFCzyE4sdDZXiKcBIz5499kjgU3g88om4XD5UplzflefaaSfvPCAo1xHne959
i13Lccx62Vxyatsy9XQzVudNBwdO1rXKsaaHyCh/yxTbHNl+V/q85st4sxaejQ6h
mjJXl/OAPmFKsjbpkUKIx6yH7LS7P4FqKr4OAW/CDR3R0sX2JgWa3A1xLV0lKYV3
GvmJu/o8qnGV+n/2w4CP35pUq1mF4hon7UaAFCWYdGschwqZmDY7MTn9WDigq056
fyJ7jZvUUNCAZYhV1PlmG7FRCW16EVjF7vqpXsK8tOoG5REezzyxsBVJeC5IEEa7
rwmt0V/DAZoxpbRpI0Z21c0MX03XDCjE0cGWXH5KOANnGkFBrGX4xIkiBcYRQNtK
b8rL0dVFT6G46AjjSJDtGaLQV8ysSBuWXQ3JxS3zX+UoL06Ucq1M5kr0rOQ8umXf
Mw9u7zPUbVnRw/xY7OMRYNuTIUKJa/X3JBRKVj6XvNtbm6TbHbJ20fVjmz3zBKD5
3e9DEUNlHj7fboVQ737vMz0aq/n461oTS9xLrHpaSjnSiME64PisZn4Fl+I46rsm
26pJUWrZN/obvQ/1vdWWEx6gtMRcS6bfPfL8OyuEd4XgkXJlid4LVZw13gdTifug
YILKvN2KNXiZ6S3VfXPoFZN4JR8orGNByvCTiDP9sUFMPEEFbwjb42TEFDgjeDJT
TM0I/6pe4+Ni4t35KQIlqlkME1uC0dwSO/gG+BJcTsr9+eAzBuPf2P/0Bcip9a2R
skiFoGvaifhaP3bsud3Sn8Ma1WnTr61hTNoO5od7VDetCPAT6mktedQgqDdyZczF
eD8L2NzjIPCk6iKUdrRFKvYxz6AuoRB6U+IpUDAzzRDbYZ4izTcJC8ihqriltDuh
ySkm1AHWosxKuIvwtjM/D9KHpbtCW0akRDBbYcN0jQmDo5bP5BJxG3o40hqXstxB
UAm8KK/oTaFRFdCXP/wYZXneMUWlZl39lkaRlmqKBX0FgNR30qftHpyxCCkXpSlZ
u/RbLoCxgkOCoCMW4fBUSFV+P6AHj4bTxfbkhaNwlNB/R+l/01fx0sM6zLlOxcTZ
Q34sJmPqOv0vUfptAGkTn0e5ldGQ/F9q6p2uXyEGN+hDSj0OrpmjTBqBPJpDm9fr
63SaZgRZ6dwnO85JEbeyGzbxThi30A/CUb0yRW5PbxalrTfZNydb0HcAOdBkfA1I
JdUc3mC3ZCJcvItHMA604vL79lHBqgIPVyqGFW9PkqvGCLs1GDEngd4+EF84oWRx
xa7/Q5QSo6kvlSjZ79KE4JzkLySPg0vzyvlz96UJ8ebeLe0+IcDgD0XtwwgUFhF8
nv0jYiDtAKm0w3sSW1SWvONFyDIdquRbyw50zG/mmKYENQKgW9uUOQLUAjxicVH4
CJX+bGnCqPR4HSgl4VqCUOWYZVnTnl8vBYZYKElNlzt4nyjDvIT99GrE4/1lrkfD
3FwsVWLZ40JzjmtKdb+2EeuIB78tashjCzO42c+/nMgYx4Ooba3dJRDM11119QR+
5313bW6Y37FfJbzvuinKTtA+0GYvwPzz1pdrraGKjKH8UfRKtn09C8F+oE0j1MLC
PGCWJv0pZtR0HbAnFi8jhTH4PJMftlv6fYRcvQkWcO0eZuCBWM2Phfgs2ge1icBh
4LOhC0rLfYLZbGZelNJfzoFZLLYHIYzTbEnF6jaT15ZdZmzShQpTsVRmHLM3jKCW
1EEnwNVrpiKgbQ0IqqAfkjSqHBRjY22LO6bpl+2mOch8ZokDhSRHoeHruaZFkj5V
GKXmCaefgnxUkxxvLj3dahJl/XhOZNseZDKcxmkZ63n2XVV9vASQ8cDPA0H+2Kvf
YR6fp/AJgNIinHXUh8GggMPwsQvp35jyyzyjs0LEgM5fx+qO3f+rP8dXAVGV7ZiD
iI7TYrIqfLTTN4RYDWwMnTbSSEseNMoaeY+SK/yrWSisRJLXiTWzhPPvOTzKM8E8
wO5u8nOM3tofihOkYM1LG6fumfqXKANSo8vBFH7rWNV/5ya5+C8GtT7flIA78/su
mbIJ3jq+RI7UxC+HUAxdsJ/Lk15iYLmlFQFzvGp1OjEDDR7ogGPT5Y4OBW9p2ihM
T1PeV9exrtzy6ygg4t5c2sRoKVyWpTacXJt5V+aXPSvqpoTf+PWWiZ4JyEtvW3M2
Q6VuWbFTXs0oEySkkZY/nms6mtL3R/4YPAooTJtg3o0ijL4ALRi91lpdtwUzQSx/
bSqsB4ZILBH0e8bSTxlTzRL4ApdP/xKPft6yPbOpc653WhHcXswmYX1uXIZBBjIU
4L7eqwR521UgJGKajt4MD5gSMbmqcNUnfRS3EiHmmQylbCgMYgGQH6Zo3qCF9+NY
oI+TBTErtwx1IZlymEJFDYgPxttR8dT1INvAtnU26EpbtddSBg4fndi0INR9cSBC
txuPRxuWF3uMCFjH4v8nxMXibvufkfYmD4v6B60pa/2HFlXYVFv2ecSrARnP/PCh
4IfWHUPmqGkL8ryANJwJ26lhHWkyyyaKehH82HhB6OrOjusoFKID/9hMk2hp06AU
80iL00F/xYy2ngeVmJrMz8wT1RZlMTzNoaqS0tJQBUkM2izzkyqzJiaK1/c4L0DS
2D3p2N9OfdJcOb1lyjiYZHIcNzU+jS1NLxLlXa/cGkmlWL1/YCEcBHPWAkFmjd32
lV0kn77HExt17FL+itwEziCIj3Gn7Ke3zoHAdfHc+aYM2Xj4rj63Buu1omyHVUDp
cDzK9BnToMscg8TwM/kUPG4KKodqnQD06r3kFz4m7yolrJee5SBF3qgmGtOXtyQ1
XuPg4YKze0BLzmKXFDeX9DLskkTui7ZWou7WzMFTMTKjrMyFA2S+rvv5d1SMBNZ1
0NUVDmz9YuDSQ0heFRCTP3nF8EDk+c5mGzl6d287FOyt3CIdbV+ccqo/9JCFhesx
maFU+hgoVTxUzslHu3XZEmBP/a3raY8RIDYhJFRHVzjn6z5AVZCe3T3CmJ3khh0+
+NEimrvZl9RQZPXB8jJRLKnUx+GiZt+2KstIEYWCt5s3UnGrx8dVwsH+ivAsoPMs
TswRn8MRlqBCzjT0cxCFoZQhO+dGNtXTX1OFnujKLP8bWev84i14k22j9nAslCGO
4dmWl9IpxgkcXs1xnc8KcgrvyEnjxvGroc0joeJmabtoTDinZ6g8O1YNE5B9ksqr
9ZWFvTj2jFas4yw3SVkPCr7O8QQ/XxGPjqYNC2cWu/229P6+qZShPW/qpRNv1X6E
M/YzSXl79rz3mArli8a7MT7Ad5B595DA3pfy9RlpevLvKtP2awg2PLUmfZtTz+I+
zlxxrj5TZ65+JmW2X4AhXyfw0brovKKWJnkR8dMTwkuoPzFG6VLBYY0m6zxoFkf0
rsj8WeLxCqpM37NDl20AlkmKdQahXlRVX6fXWM6wFchgWlWyc8qGtDHgjks1rxvF
dzYNF2WdQGkijTusGmn9s4iaxKj74eZATLKe1dZETNCV8ZZ02W2AukgW2th4gqVq
msxBALLOlmfcJj70hLrgeEBb+AD8Al3a7uQ/PWjo1JOmF+Zxs11OWKSzV6YTqtNy
vmbUOjHwgceByxUQQbiHomX4WywIXNI3ZE2ckUdLQhhTYuT3DnS0LFwXqv9HeljY
nzJe9rnefOt5kK59xnSlvEsSwFoJR7fU/JfsdrRo/fuV9RoUNHt/Ir3B4utaQPf9
cqW6mdhc+as9d4DaH0szwHpyu7REPX9WCZYVYVceeh3BF8ZugXK3NN7wZbm6p0Nn
ahlvU0GyGE06XCxjLxNl5Q5ntmCkYIMB3bO3lt6iNRh0RlbfP//g20UBiadNCnSt
OCzQTGEGgrQYi5Fzv+3uOwT1rOk1fxroFmjr9OjCYv2D8ZydTYvUDqQCUCvqKj56
E0RF75p2tMQgehRprRhzt4Qup0dGdApO46sPC6WOuVJ9rwIHOonT6DDFqGbvL0NS
5GmiTrooWeMyqZFqUJHw/bhmJ846cPKaaryGM+zwZSo5fMgVU4KfOpWdV0DCH8fU
HbnLYXAC5aefFY6A5xaRJjcq6i836dH6V7YfSKopEZ8vnc4kohEvtaKJT3TVheWX
fbnZVb2i7zF7aJRYCFYpt7Ffx6Upd2xdS9QNCYiu0yE0Kt8m6IP3ppY63osJ1Aj+
IA28Ym5OwlA6FGgOdHiEKW/08Jp5b8N5vEwuA+Wei2VC48S0koS7ng9bbrm0Qv23
f+R3CZnS53VxrVwayETrSrxGfL+O5DIDPLSloQnDzfn38rCjLBEoZEgXmOBv5oRu
Mg69NlRT7fju/IgppMw0hpydyOkJRhMtDbjJoKrYGu8ljbEWwKX/NZUVLGRE/siN
uoD03GcPeh0ouHDYmVPYpaC5w/FT5A7Ngim0oyDmXbUFv9PRH2Flx1VuejQgrcf4
rf4veMuQNt2sKcf7ocSg67KQouiSU6OPQpuvhz6HHIeSGumZz4xchhDVGnM1DqJJ
MiHhjPMETLcU8U+MOVguV+lAwZhwn5E7WKixVm17A4eIp4bSihXoUgqGpk3hk6fb
amP56UOGEXP7dZPSlPu3A1t+6DewLvWTIgnIkagwhHB4f+7YcUg7H/EH8/KXhd3W
h7RMqAPgVDDqP7SH+qyDCP8iFvXs3ZSIx3aksJQnjzxeMCCazE+1sODv/Y2w52+0
OEUaTWlj+KkqV88iVtEVEzAQSCSRfaRQ85P861ohr37c3ZQt58tM3D/LLwRzChzb
PLkskT7+EJxlrrpFsZKjKdBZkhzCfE02tPbaMvRda7LlMTgfxQjLW5nG16ro+FhU
Fe/CAGMoz6OHxXcqzdxaZ88Ghi9N3OZQqeNI2MNh+lEtu8pfjqAodJIA6ng5va2A
XyPdJyf1DfjSG4W0cHJ7NdgSWrpTMXVTnihw3Oemk9gjdTL5JY4KzFWIVdMD1Yzr
I+URorCvI1DpubKs3HoVoorE2dIxaaFZtSZUQbkS//MKVg2v2ZN0EdLD/V5irofv
pzFZ5MX+Fo3sgCT4ZN1RSEJrS5hJqFaZ9hDpwl2TnI2wIH09LackqHjQwy3itJxd
PU+l/mm9qI5JZZO//NjOIkG5w1H9e4Fxh2zuQOTcPhcxkkoH+H5sz6BuugI6CSGP
zR9uBVpx5rvvYMCsR82zZyfsSRlLNHJV4om0boLDcdfh8mUHZ5PmBFJh8lgvb0/0
do8Z5h0aSR6QK2P+ZCKhEjeOHbnNY1mmAqU1+38QBQ9IqLkKk/otfP+tCadLwAKK
QhTFzHB0CXps+T8xGsOj5azya0EDUuIgKYn7zb5xEcUbf59QGy7wFyPHYzLkknwh
17wxTey3bdVahK09SoicysY7tYRMI7pMuRvouc0zq9U/HUJL66lU9PvU4yaoh0LS
dO1hKcZIyZSvM1gDLjLWFsh3GMGCs+eTWDTvFbUNASJEYXuVXltLenmCI/Z7HZY6
r+U9D4h1q8NWofSACo1nmp9o4bhVgHantNRraR9+ut7NUmwZyewdsfJ8HltiXnIv
0Pn6IC4815WB3twWgSZKvxHC3hVPm8ePrfZovUzSbn2X8Eup8bSwpUqFMD6UcHoW
z5zARk9YjDLh/w9IrEqOPmkz+H+zFOKuGL31oIbURN0QHmK6tJd2CNrZ5JMmLdeH
+wkNZ7U1M2RSevKbrRaS9MPXdS28JcdLLlTVk6jj13W57PD2gmEluOATgCzqB83K
ECvAN1eXYWTBhVtWbqkOuU6v1ZwcmdAf01f/UJneGB0nq+pRWod3R1vYA7KVNR/y
1TmXgnUaX2SGgrr+IRrs1Y66Jz7UF/GMkuVZinJWbIN11EkDXG1wEXe5IQa8G7LD
rNIz2dDE+b0pHtv0qTQd6QY2RWHHwo9QZTlP3D+CWniod8MV6dpZSWVvcLr0ugxq
lRE5bJWAbrWaopNXjiazu9QHaLpbdl918WwI2Bhd7b3Yb5QRNue9sfCxR/73FOpM
pj3vs8SMMFmfJYQwdnvhdAybPdWOscopn50jOX2Idxg44FOX8MNjRQwQDGKIvdpy
pMvP7EN4nFWE6SKsyWOTWURIOp9zHt+STpx4Y6Uv/7BK4JGeOOnLrkJ867zEqmEc
VPDZe/Svd4UNAWZpdkBxxrmE1n4r8Uobdt/ce1E9rtRXkzQqr0q94+616HmaDDVI
LrG1wzj8sCMWLl6y2q9kNsMGvK081aF579eHb8QfY4kjozTAzoL+OVYaSnaUuUaM
tsuaUMCLMclVYHL/6zgzyOt/UhxcLwIJHQ2Q+HrDCpjN0V88YkSXeCw6Q/0fNYTF
9UWJiMzIosY5zOCIe1GtHPYW4G4bE0fJFsnh2IvDq1nGF+8YO7V9uLDhkmctG/ae
untwU2Zi9QXBLUmq/lsU5+fN/vPhexcZTnOy2n1JtdXErcVj8i/whFd5qGie14ci
w7EvurZaUwqTkD7y6dWvl0/cxbOkcaGuyXKkTlUyGJs0OkPIXPH4TgAL1xMu3g5g
zPamEmJiA04gGT3TelsW7B3yVzPNodvi7xA4VUtv3Yv2JNJEgo6AEO9/BHvzjxun
c3aYoYqMO45EgGWmW3/NUALLRyikTXTVAkj+tdKpeAfgXyLp8tkQsZQX+uXzz/nd
UgxpELmxw6uiHrsMs90m1Pl8fiHKifHQCLbRb1iRX7YryNpmBgARSgs4nDv95dYz
0yZc7LZhvyu/wM4fDi6UzMHuSaV8mJb1pubJoEVSvB+gRqEOQv2FuyZ4MDdoTnUx
+5bkHGeEXqnJDRuTfLiR29VlIO9XxFOqLrKSUgwGsfkt/1hyUW+svD6jRQhGraVC
0MkryNMbKQZOKXOgT5FmspMc6ApsLpVZ+tC75nWcE6glB+f49TRtfl0lwSw5rYmW
9bBhhnk8nem+moljC2yATAY9Mf+d5JMPujphRFu/uy+w/5uCarZGc5FTAVgedyC1
X16Vbw+Fzj+Wc68F8MAjsoGd01NKy78ovmdNHJbKxIwan0wTdTK7U54tbt0bUUe4
NlfRykN5F5WO68fAIGAgKZCh4cXxPGQ42VDDnTqkiTW2mHz2XYZpZvmrVFfwmtwu
cWvMh/UmygpqY2UijVDXvdnEboxf5Et/DcsiJHPA62cwV371lB74hZyDmh223o7O
fv2/gQfHVKLdcu8a2iRLgn+7T97+81FNEt3vMdfx1w1lLRdREETMjYl/GZ0otLV0
NKxo3UC/Gmc93NoNP4h5+UJvxbMyCGreMxaPsUkpzsEuoa35lqLu8QHgdjIWg9Ls
nG4kLwD/gE/ngq+09lq8jSMy4k9Cok+H//x96IKK9DdJN6Ea8BwasC8gU2GvlA9H
OayZvL7u/e2ckh8O/3AdFp91ytCU3pY1i83v70fPyPgisaEwlGuRBSWkG/MYoqOH
Vgwq9ioMMlEql2oI06kaApoJGFL6Nvw3CoeE9QgzMk7uG7cU+6p+H5GuEbE19es8
W/kPjF4+VlWmubT6Dfpah4KnTRmJ7LPWyWTPRVGo+9v9NCIP+y0YxkhS96tGGB4L
S+AmK44zS9IbGt2l7Q1T5XwjIbSzuYJd8FTHWAK7DZrqoD+Td00V7OkDa6lRzRS/
Uaim5me2TdUYRwr9X6xaHLe0vjyai2efxXYCoTMBUPaLJss6ZW/bOnXOa+UjunfY
V43/P5wJt0y4ieQC0/fqX4XjwsA1wzTXpPUpQIKudddOnooLV0TtoIi4BD8BbTK6
dlw81EO0N63FmYaunhk1/J/EF8oRLInHTVW8PVvRUqpG4ayyy2kWJ/15He5zVMEB
xqKyofmcxATz7HqxeqYW1DuDEjR/Im1YXod9ZS7OWkX3KExWokZytAhH0OFsZ3Y6
DHx4Mi7a+XdV6mnxxhUUjIxNr9Ihgpw3mF0C5Na3SRmmupme8UMEjUIwsXIj0eyf
B0n/p4YeQS7rjLLTY9nqNu10L63Y87j2ZYhPrwSJbcmrrT1at3JbVXkj920YAqVs
E1V1FdSKF7mypbb9vf3UPN9fRveawz0jkvgWUU4nmUfsbyL+tXOj3RW9ZqJrZLpw
LiPZ1CXcgo9nZrvLyzuHK7PbenBcIKs6/Tsry6vfxFQqqfNnjPnqc3D5CMVaDd0X
NicXNvxbOdI0R3tLwPJ6UDUMqv6uauWlJAyUEQVhUb0OdUv04YYNJshwsqvW5lhq
y+zwXFGg4FnLgPRdmOCpQRnoHHLdbI+ghsJYJkwwxIdutMrxmBfT+E6BGlFNbI7A
w6A40vK4XJxDsDhyCUBth5Zjp2qZ+VsrDECmtpQRHEz4Z1oK5ZM467idonBPJZa/
p1GM5QCFcOP+p2j53mdzAO5eS7DFA1hBfDFOojyZSI8GajXvbE/SV7cWC/WO/laC
r9AyT4JbnTFXSA1hjSsD8Vn/52Z35WeCkZrMDkAF3wFgXI1VKgIHANAndlDk0G5F
3NL6mpbTMrW8UZgc7CrROqHoYeycCBMvGdOrOdSRc++iMeym03ZhQ4sUIemsMakD
UbQBxoqivQ7XmWBUhLpfaDlEkR/mlkRK1+ugKuag0qiLcref7o1HNAD/eHu35AFt
YsZ1T0TwVSLur+c4Eo/NOLU+PVP5LFgjSKBvdsuyPlxinxwTjz5Ar9MITRedXV0+
chmsNuicD3eLNnO/cUKwemEQrEwVTRI0g6kRO2GS6a5mKShgG0psBWiw/lD0pS7z
BZ1e86vxlmhW1wF5tA0FfazJ5LKkLmjj/CSLHjImS6cnKzbA9wtWwf7eyPx3FJ7S
J1+i5HcIhgcgDlbQZtynUH1yXoVpwKAFXu5kYr+E86J3vLYYAdEQsztMYZfH+slI
B5vpwV6uGv0aWCXVz6fKYEaGKExVSezO5sFB3apLHFPNAxGYm2Zfr5AM+C6J2tx4
T0ooVV8t73UwHnCPElsPOIP9y19dDNFXBuRTiBYaEFxKind7Rwi9gC6rcoyV0HG9
qxf8zET/JnlTC4qH7oUelyOCehAi0M08owtQaT0OR9avPs1GPm77K4OgLVKMWLMr
c+fW2+X25cJJmuOBv2Ga6rKzeXi37oXP7qXM5VwfeWACtfh0J2WgbQq2AQFuJdcy
R+G8MAMKdiWZk6WGloRn4CbgsVZnpxVg10tNr8ikNFHGUbYz33m9WE9Vg/z3bzVJ
150pXsyipd80M85+kKLxIny9TkTSfwRw9EQGoA1EGdGYaMprLh2ydvn2S/64ZoaM
C+afXdu4SMJP0l/whsp1+Fwpem9nnaSGit+/vRBeFrZZb1uNrpO+VREos5l5VHBu
Cxlo0Ol8JLNA6ObnwWBYOMVcdvWOWzLyxVyIB3nXo56T1U19xgBEmZb3xdhBJO3B
vAJcbKyQs0CIYVq8I6yRI+9oiAICh3mGNUyDcR6X5eUjO624nvVHeCzDdGnoy9Hb
m3qbaK2QzyfD/LTKsXJmxeEvI2xzQsrY3bvAWEwfiZ+aNq8FJAaF9UbABrQeXaBG
66P/iUBHvat3pGkgsdztPBQSR3v630EFPxyiPKDmfEoWJRPoFFoqPLyI/r8xhbhL
aXwoQm9hGnje7Etc7ciHEo6qhrOoRtBpmxkz2CoFjuR4sFz0miYGKlp8rjTeSh0s
D4+3hjomTzstwmuWUEgTqOTQPUGf6ijkQQath7u4vpIDJS3BhHJRgETX0jjxVQxC
fGjOv5Ua/uQIj+KgwM596ns9pDBRux1qsdGPepTvAvHUxpZ2SoiWMkMqETkNrqjE
5IwvF+dlCsDCuXlxL8w+eQG8Gsd/37b0Y5AYzR+SJw5nh+6nsF3ClmUyleZL3EV6
Yida0BOSUzgrKhquBYOjA2w7NtrWHVlGxDvVEUImXQZCAYGq62rZe5kGQ4GqKAf6
tQqJ6+mFWjfKsAkE+aCufV6nHipF/Biv9LXq1tQMhX3CTGdzCsp6pBOscXrMNbaQ
8za110+0zkSX1Ex2MrtzIEgqqowpVzarFxb/S2LaySHXHeWtqygWeE+uc15R6tGY
cLHIXtvS9mBAdDFDt2RAEzGTqcgBE1MW+/HxtEWiwUyQtioLeh91VpTaKEeyZX3F
aintcKgMnoCCbKCl/KmbLp9BA/7SF4poWSl+/d0CxqW0C+c94KzFu+tNwupc1OP4
PpELbjSiYVNoC8sSkufBFHG4rAp6/Ab12focfZ5hIBd37O6bnv1DoKHLeC0pLPmK
IfK0nOoehcRvyCKgvKpJ1sejkyhQ2on2fBRbdH6cIQh6oiNLmmkWGgkC/P/f9Oh4
VqsoTRRMWmMxBi/BQkoVCD1jwrRHW9dlHrC8ZM9ix+2JLJ9IR8SCBr94TmDhv6CK
AxzNGCfMsss5xTwqYcbRXGY+bYOa5n9s8JPgvJ2RpSXcBD4gpgtuFzHMsDbkHnaz
4JslAfYgi1cnjxVePMl/7lWOZQI3Zgy/BKIVTy1+hltK+V3dusOGv6nTshGuU3KB
/CaZUtztiQ1VES9B3t45bp20kyZbIyjVOpXTcMD8rXNaAWhioJqpk0qrXm7vDUHS
9dqnI/ync9sSKfSPamz3Ti85614kbHsRG5W7kLnV5+/WBTgNPMiT5A6kRHt6+vid
EwsoAfadaoQ+YLqdEBqZhTCIwBEzyV+8IK5hK9XHRtD+xC5NEvqxPx2XpzgnpYw0
xZx0e+5Up0bFlWvSB0ziLqffETJfFgp4WPkqtbFO7dvmmTMfWovG55bcQDH7in5D
tVHPspUJPZ9mq4sj/JhopZyjsyl68Eq66pISWfsEQ+1erKrJVIJZO83RgnBcIccg
8lXRaiZnEN8Cqa9zX9UV29qljYfnZk2JyvJV482DeqNZCsxNjme7VEbzlTm8fgVc
Dv5gS+ReOdenolFnGrRlGN1nDW2ZGl5MpwjndiHdjPhPLYoV6hBLMM9vEMwu+97m
ywkijaTCMMxWv9NjBwmq5ZJcWS41YQ9FLmgasufT7GHuHhcnxBrrtntFfbQevEzP
mZA3RrTelaue/+6/SakSkjqcDp8+wtwI6nqPn0DzNty3XOSbduPHPDhwsGzWSo2u
FYyQBGB/7u+T1QAhCDP7Ld63xUIbZf8J4DNaFeLyjI+j2920Zuqdc7Z5PtKpILxy
FcImS0a/oYjz8zp7DSAROigsUfLBFdFkLJhmkrRtUGnXkYTe1uZkXCE7wUXg7yUn
rIVc5vrgdXh9pTTS4SvFs22AQV58mQLvA+WbyUenLiIG1mx9i02CESLQ4H3j62ka
x03mWyXkW4XbxXnChpqc2fwKWSeGKICexIaBGdyHZHI+feuTyEcz7+UTdI05+Pbd
/msC2aQMwtwUPnE2U6xSwHi0MQlkpL/voKveia4aPeeSC/ACMU/NgBw9PHjyyCMC
X+cTHWn7pDwtJ2SXbpL35iQmtEiTvJrSL56bV4z1y7d3YQZkLCqabZ2GwhQ+HNCz
wPr/0XQspbd6TrJ33axwGoGtZKmjzMSobaFT7p455yiO1lj15927UlXCazamuDjp
VfmwtsMF9Is/VRGzQJt+wyvk4RZmrfxvRe4AWSViMsDHcCDJZbonvaEMJZcNPRMK
w1VOG1wjilrMvm8a+0HhEGDBIfkXR0sR9S+9bk24/5sV/U+Jcu1q4nGrzKuzECov
0VxJcm1jaa+FCzm3BlHgDrLXjmLXh7QUQuuzp8d61lKgBbVsc444AiqyUPPX0fL0
HpoDVQAuyH1oWrRqICL07mvW5OffhSDc6algewbdw5lw27dtskJAV1NkOiIzvzGV
C1of0Z3ylUuQXQvMS/JWu7FGSlAMJiLzID9w3DP1Rmup4ki2HcdrlePwhBV678gc
eTndzO9+c8bPjEXu4ZTfxJq9hY/b/S3UkcXVMsU2gc7ak9jpcLqYFc2hl7rUO7h7
EaJ4MnpjwnanbVTpDxulT7Hex/l2FmCkzya3eeqirV4wIk/4phX/w0d2+6zl/ZPe
d8vKUX5pvuzFZ2cwbEutRjiKi24tcSiR5clh8KfrjWa2fBRcZ67YD2xm0trRs741
O9J1v+T2QdmZk2ZDauFaZL7qui7G62xEXQ0rGQe6nzge9hSYPMN3kul2MCQX5H4U
2jlXd9v2VLAs5BwUBeKbuI3/sAbXaBCZg3DO9Pj2skKdCo7gv8iP4GTR167K/xsu
03KYEg28oe6IK1CAVzylL8bRZzcG8YNd20qSwvoprxyXHOBlqf/VDdiga+wy7V+a
su+JUDZLP6r3h7aA0Cm7IH6AvUbO97/RO1XxW5cVwkZDwqp0Ia2SjMyjsfUJxjAi
tphfssJzE72kukWSuTBSOANxSuDjvjb/cGMctSzRdIESA2g6HEfGEFPoWefgLOYv
TKlxoUO9emTLJe/4t5r5bMNiPS2onFJVNjZ1wB5DfYMeQwSJyqVLiDJ1it6FMbrT
rZcpEeUUJ3IGuAXYNXIxOQcCmbdoS74Ewv4yQsV3mPGv2Yq3MPZOdpX9ntpDXAJB
tkrXKEX3+l6Aq9yAOGo+XsVROKKy942YucAOJsLWbcFjvDAslMI3vA6tcS+pso8w
liAnHxBH4MB/y7HnGsUXVti6OB5zDdszKqDnHc8KY3Hm9fWV06FDy6h0acWe3iRg
Yi4UDLsUlwTwuP5Z5XUxwS0Tlyb2h75OygWu4kL9o08pZI1iqxnBuKXSO/tfF8l4
jmrpITmhGvWY/tkLNkyqgKAGlMnkc4iz4DJ+H+jmNaEThcyy1vDU1yknUxatHIE0
+5rkL4BzkL2NgVSC1gXr2WI93CbkkrIUahF0kjLXszTovzSFH51KiqDGBtkF76hz
cVVZtF5vXVyuCJs4nX8gHRU7535gruasznpSWSxGC1905kdiCsMAeMatnXrvRQYE
Cmhb8OaFfVKkgNTQvcIx0s6i6+p4ZsCGtHTaPN+8kmAmKDUdh2V0TZCalYPoG4Ry
fov/Mpz/jWVDzrN7KURdPp0N/7ZnGNF2he3xMuvHazst1AYkJRG4NQGxC+JTNLJ6
RQUCTSvSi2dSE2B15zNWaencLq2giJL2hGrqq0L8W4ac/60hmTTQSKYbA4ylS2pD
s+q/TttmFzW3KErPAY2WI6VJ9ITinHdrnqbJajwLe12T9OIjZgaA9HsRoAYX0Xgf
QdjotKovPlTYNIxUxPf4oqCZOGyJGk59QNVtiFZ/2mkD981lcdDa5rh0MsOTITNI
cKJQ5/Plt71KlkwObUI/KJFuaIYv7RDDGXIclPBJo+icnKChJ8oaJOkJvPUl96bi
8rCt5GHyl/OYRPs09XPG1XiTt+l1xnGImhuCGsE7CzCoobri5EaLemsOvghkSqZm
aH8wt26S/GTq4Tmxv7pL0Dm4phoqGR/F9EZTqMM2/61dPocPjj7d2yilf1S4t8Tj
s+pgUytxXZqX4oSQ6D5ru/scCD+EI2T6Y+wPej6P82LDQ29ip1KQOv+aZKIy+4g2
v5uj7iS/QOWoNQDwqDTKCKhulChsZWMk0WY20e4D6Qmb6QT5iqty0u/ldoFxFwhd
j/bKcnVXowTyCbjRjKoAydsdyPdxlaN2YV8j5aLkTic9sbO9zR1nGOeqzy6Myn10
aHbVeE04z7f0EXERBqKoUVeNDEDFASBB/9LlYU/wjn3alQ78b++Ct8F0U89rTNFT
sBBXK50p1+OLW0EA1x4OI2eFjEsyMhqTFVkMSqIBV+8VF/mIM+57zmDL4EbV6dJV
QxMuP6EKA4YDT+mDvFZ1NwBX8ZXuR9GSjA4VjNZtSnr8zsSbWElSWx/rZQfGOnWe
Zvt2CSMnU3tG4h2mBBPvvmzCdYKBNNaBlzJSAFWWCHAfLOm2yCBcE2zl3vCWOH9N
t79LVNF6ozzJcshi9AgCxYlxTUuTzXzaxxln36eJQh6bBkrTvaSOgqiE2OoJnAE7
kZ5+VI9fmgpYRxK74qEDOtDpdRAxXUgNxgCWvqvMC2MQOJxP978esscOldwtnsrv
k7+p8S8N9lYETsQEIekPAsyxthqkYNwMsIaQ64iOUKBxA2XhO5KwyWApqRn4P2nF
IYZvACPKB2kUbnBQJ8SeGOQ4EM+s1zaIFcvXGzqt7BdHhttGkDi/lAdWOqBACdIa
lYjfIh9I4kYFCrzLbXkXRlH1RuTFho7GLmeXQNKpfb9jfAjv7N9mNRw+xetphV6s
oTg7sWzyNLvCEcmLJsarjWEVS+zjpcTGxwc3UGebCJsC1MAnbyMO5BgVNixDumSx
EpjHUzyMyP93x9bHwmv8ZgGrrqrax3itpCFyJAzibsJdShgvVd+f1QQR4KmhJFWM
3HaGjE+MGpLQzWxrzKGVp2hzxu79PrbQcRS7Qh2iMXDwd85YckzIZ7xBw2TJrqi5
zy/QwuzZW0humZxmYHtPPyoTOSX2PSbcI2EEzko7/Zq7K3L1bO+VTZ1tSWXGd6TR
L0dO6krnKHG6dgklzqf31YSDcNYkJ5xkF5aDGR9/QYlpkdTmOePPb1oHhL0zAXxT
rQ0Rmpc4e3cTLjNo5A+0FmaJGCPPOFrX1QW/uBPNCLy8tTCJCRscLBZ+F1oAEnG1
F6IoCzFJbm1tx45DfzPm0b00xu0/+/KcjEvPYGUi1pGfRnjb6zeq3RM4SgnUxcZQ
sttRpoAGldNXkaFHPbIlRKrRPltcwOYVeFcEcGw21aAk12zri70p/TYtFqapWaZz
ODSXIrjkegq6/LAi+NtAubDOlolxwUwNH6GqgJaGvyHgKyznkluGsUl44oYHVgnt
gkxd3eNVJh/WnlpoQ+IRjTAS50CSsMt6PQsAKA5v4J1Xfri5JGpBGz/CDBDdA/ss
v6gc/hMZewN+lpgk6qkM/N3YQcAI61zdAc0ajXI0ZclMB5KH2Ou8EOfsAQIXWXYu
DJrgCl9CiPCjs7rE6fxzMu5J6BbTlX2qhFMmbquWk5dX2vLtnICGXdlMWTSak/bw
EpjPyeFwYi7HbypO5ooWH+H8AV9q+bZB+wF+3JiotFg0bgj+eMB9QoS5un2T8OX8
CxN/NYrOJ2w4WQEc2OHMd6f5mXw0OfVyb0KfmFgXWpjS8szSTWHPRRCkdtk5r5Yo
1JZ6VhT5VRvQh2HVIzP3RukfmmDDkwyq7bY4NM0jiosuXk3NZYWlYxjB9wiiADyr
crcfdjd/azPRvaGtWo+Stpp+3/6VFDcUyItZAfOcN/z/Wdnr/peNGV2Oh/tuY/JJ
wL4yYjJm6ZkaHZvJdR6fbfGugrOUVw+mQ4WAh19Z3baDsTVfUHphLa18HOertu6E
V0FnNW+VChriSb4MyMbg6NmZlq856iZBHp57A5bEuvBGm2fdOG1hxBGM6DohwiqK
iCUSOlJsAWCUbVpd0NAg8OlU+iJp4SwkKkYh/BW1E3xiFPxiI/y3o0dWgKW9xgsj
vuZHMpNLrVsMGBbtf0GfVjKRqn+zyvBouqJ9IFbL0Z/mluyf0PhOvneTJ9jtcKuB
JozaMOhwF9ti1cOdvkbpW9PShGJ6dh5ZDSGtmFUAZOuH3JE3y+oWhXhzp/JnImQC
yR4j7PN8/FjSu1NNqhucEoioBASxYZd2+/6frLuhnkmKS4fzHCnZiTtcChukoFhl
AFrfqIHo5bMNP71hRCtuibhWlySPCWMMVC9FIE7GvMCcG98h5Dkd9wh7gs72w9Sq
jLG8Vbj/a4JTI5O5o0T9T6wO6eQaxWaFufQ0JBYwM7lOAcUszUsR32s7OnOtnsSH
2fo8ouWY4PsdgnDbfmmxhi9YM9UlihluKnGyj2U59JTNOjAVmMyKUi0FVyRsJ5It
EdZYHTNkNScYhPwnrZLdQlRNRq1cKV2n2ikwXA+j2po/eBlAncQKEW6j5fBVItoT
mLXzEPTg4jM8Zr4B9mdBH7sX7GUNoJbafOXirgDrmJ3NvCrkoixt1SGMJN0Qn791
7kTM9EGdzOVEAm5c+bsnMDO33DjR99u8TxauRNrQCFxsR1v4hmOtYtyVO1YwBhQb
zymoKiLyYXdGXBz8DjNG5FVW4XxhqSf1bjKw98gO5Rm5X+49giBfu/n6G7AzhXil
QhToOpzBcbR9wgzqzmGGHXYFBX/2hwOXjSopEZIvEea7WAN9JGlMqeKPXbpbmOaK
zLtHpYgJgWJIuD9tiuREz3rPWkixOYHdTBE5YGpjumco6hLSB8qREz5UN1rEar8U
0smsdLtXmTeme2uQrGwpFUeBK4d/pHqFhJGcZJltbXCqtYfVJROkr+SOcCIwrY9V
/0sVEniI83taMI2oq8tKe5dpTL4jTEgfih8JR8B2X3/ZfqmfdhyD/FUXr4wKXgu8
GJnSdlMwmNGqqgAfhPY9y3wUOBh157S80L0pwuwRmkOxQZxQEaCofUzz17+Pu7SU
MorKx++QudLI8SiEhPqAGK/iYWtyP5qMgAdPT3BDMjdx8pHr/rCQAPWhCdIB/Bc3
9LtLfGbN7CUia6GmeFYH8mHVFCTGO16dBpZMcqlKOgUw8A+z9jhXdJZAHBvsbi+q
QkA1VTRhcN2Q5XegAVjh8e6fm3lenNE1mcxJZ8dlvycJgzl6IwZ96AgSOFZ6kA7R
LRxDHbkIgpFetcdqp4W963Q7bUxpDG32wNw2TW6J/94HhPE+Fq6Wsq5LI58b6ZWV
9E5Zirn8LXot3uvm1bQTH/9BrHNOFkDDkC6AFFJ6JljngFnoYtb9/+a98/FVNj6u
bXLbYkXlk9DzJIruDOBKZDqJdlgHhoMcczUo1+/ladtVaSnVlKCPRMMGpulH1YaH
W5q/mMws61IQfSXG3y4Ir1RKTqSsW9SoCakvJk7D3LEqF8eetNIWvHX6TxtBQcmj
tDLqs6fRFcY/Zogz9IUEqoxVPp9S56PpMKMW6z04ddmAg5s1PLV3JehatQbLj8zh
TM6A2wizZhAwHQl3jr663i3dTthXNslOwfkSliMWGEsKmcKbkCWbAE4SXCwMt9hu
+IvfKC6S0AjihleFe8vin7mB8XDKki9xTXaxu3GtBuTgSD5alPtpcWiRO7d9xRG+
m72Kiz7wpsRKOmv0Huzaq8qhn1YH42hFitwuw+9mxCq+fZRyUueOb4ao1zn3aNV7
jTbBVdj38zyHpXNqKODeVXUgo3/ni6a7JHPxxHRXs2rAd11RwZRZMbj1jVv/dVJ2
iMGCr2aLHLMU7wa4W+s/eEyXM73ZivR1LJSHk7HyWrnal0qbFasil85KgEDu05zC
GsVim69aMuXfI219r5hmt3W8ssvrSPAjIEBHNqXZDyNp1BPX5yvbyzArngtG7e5b
Z5xPnV/b6q2tZCnkNegzh2LiY7CDNN6JYnjHyWTXL/OAf5jchMCOaXG53yeXC2pM
D7sjaHxPX8Z3ZqrNFf0XdY4kyvyJeo5vykiDQw2M4XYGk1TnI5sGq0fbnsK8ftG+
wGA+tvxFqQMMo86unVcuZq3kY9/kdOg5ZfHHSk7HIMKbBz5GgBpLt3R1GkASVY2l
acSk0V41cs7RbUmS2JK5b9+Fp6yghbJQoYVzK7L8k7GY9U9K4TY60h9CimmX3y63
RKXur1D1fAIoYk85RyZo/+WrQNzfmgjXxAufwssCsjW5eXhb8xroVHPEHOU7nwV3
To6cs0yYbg43s4mJSmlFOiJsg5nGRx6Daf1+E793c2fJfcM/WPdKheToYE1jBZiK
PIevDMEPx43WIhJ9Wk3t7JatpKBRL35L5Gc4JP3BC5P0xTZImDRECe5gmOwBdpWh
S0noqtcOxdjbtktreDNZjdNhGkNm7oH4TrP9qFWzfnNB6IvxDhMqEUtbSPNCquyQ
jSDTpzzQ0EELft12QKLRlbwixsHz/qY73qV1ejFqeen2ZvXAoM/tS1eFOYvAr3cR
psei2je5639lulUmUE0aJSclh0PA194s66mFLJ+S5ZCI37sr0qEjqzQ3089yGhL7
ZN1YxC23WYEQRLZgB0LcepmqmyWUCqIKNUkMtmGnP4miw2Z/zrJHDBKez8aq8low
AyHz4XLroNmvD/bAlbU0qm08XfG8lHrIMNSrGeorxUOCh+DqQWbfwibxXQCK9KRE
f78oTEs3RlXaxQ1b6QJY0Ln6sEhG7bcHtBwSgKlpsfBUkaEwTAk0eq5tzc+qXJvh
LcSuPvL8nWVwc1YkaBQuThAhZXJ+fn6uy2eanMP6dFqsO6uY3SYW/yjRZ1nBQnCh
ihFu+gyEOWZxO+80Qh3xD8El1QqBUy8SzANPBiXZqIz9HiCnbrmlrU93IGGIIIbA
x1tXEOw4pAG1ibdMcXm33H8sFcZnzrmefHoPN7kqo85IrsnHHeOcs3/qYt1FdjDO
yrPjA8RIIoEdFchxi1I62gGWF4upoYIRNWLsEsvVarQpiwfQrOtEHQq7kJaFyGyH
79Yw/X69/8qNweHiG00M8/YSTcLudaSIBIlf56XW1BHQjOwCNOwstI3qiHvXmwv1
HCntAwGXWjv4lWVJMsQBN5JUQ2t0x58CP2QYvN3PgS5b5FqqgMfdrKcydWOqMnef
P/QPIFDa7J7SPstDTF3APIUn3o4ntwuuZIn3QE0HZdpYqvw18Gpky7FIca/lyVbW
MnhZdYFFzDoSYtzLwfv8zvhZMn08bSIqUkAPhqGPq0XawxQ+nQGtfHIwPz/DAxiM
1XfAvQZUeyEkD1BDhREroj2YGFNPlQpGsMhFQOsrXITSQt7T7KDps5RtAzbZH5x2
w9XlJLx5aibvUBiJcMgT03Zw+ERyA/uSLq/1snNpXpjOjYnvClnGAK+IRl9G5Fg+
Bp8H9kVFTT3yw1uXNT6tetFWRqq+GhV8pzVY5Wx2I8MLdMxHwe3LFbeRnmtUlA0x
1ks369tF1r05E+N2Y8zVf+0MvdiI7dSX2KmJoLH3Aehh941b87txfH7s3t4qcY9P
qGciffMqCM67RlK073R6mCtEAfKVqIkG/tTbpxDhDKBAUNz7LlYtk+U7GKJerzbC
AWYgpmZllHAGyLDsz0QVp6rQutJf54FnGBchspMlflV94Ai4boGw1euK/d/vU4jD
dS/f8XFkee3FL0pabNYS3m7uLs2oXrlRjRvemayOgYyCnxvOfSPXUNxpM23E4Xmg
YtmTyYL2hfLz3wU/3Ce7Wk4FHF6OReDwprTpyGDnI2AvxOoovZuYFT6tNUI2rTPk
tnwMfxi4C4oWSn9X4QgyIGI0m+DJtJdnzbvrYm6VRXj4UBvC27pixgr8NYXZfn98
CIpPOV01QkSBDyVvOLXJqHJckNNWVxhVPxHS14JuD/wpiQLzuAAXZFHfi3um+lMG
TDyt20XZAxB4AjYWjT/NW6gwlbvyo5evTdgryxzJAK0zacCiAX3nkBYQssjVlegR
lj5SDV9YvT+SlYUdqT3jy0M5LX/t3PMQR5RpAYAIE2kr3OR2Y6OCAob7/6Y0Kb8B
r/iBhUj113qp3L7XGtFUTFMvnSAFfu5QmvRerpnLCj1wsSXma64v7AQ7NoItNgT1
Ao48Owc5J/KDrBZStNnc0DG6KLV9mdX9SrLpRKJGQhmD6G8ezr5RFNpP6jJInoma
rxUhe8Vjl7jGkcLHNOFZkRLmI3nxLbckdaoer4FV7uQ0KwXq4VYiBsDKBhaepvnZ
efek7wrxymw+zDF4y04ZpCHYV2yic9X6uLM7ZSg8JUsa0lOLtffLTRzlmEXbKP2Z
hUIDFiyBq4OACgujTjVh/6lCz1xb47kSYHOKrj7zMAsaofRon656IyIsuHbtfDli
LPG8FF81m2sw9rfKYAa8/qUrIDAXwC54aUlWiEOasG6HrZMjWkwUrhFZQtu5I9GG
+p/KVo2Ou+fk63N+VJep2JDFOc/EpBsRY+iD162Y1jFlkAkqdrDX7naRppi1LK5Z
66zJvtitXcpBxRRmRHPD78B+Py02yLtCVbs1a46bhs6zxKYa3UzEsdX1z0yxLeiT
gn9Ph+8y3eAIhCMqlleBfEqHDwyr9NSmvgSZ5mypaTTncu5uYPrjh8Wkhn5bmiUz
x2Y8b2OcuVz0uANgDgxQf2xTDoydQooFjhjQxtfK8xCEKjs7gsO3kArHItj6ITJ4
NcjfKuIxSqBbFHl9ud6OjfS1Rc7lCEGRRSTMK4fIkhAFv0uhsoOZR5qjkg2TYKgW
9/n6iw/57wICKrXrlPhsJTAbiJipwVOYFZ0hTp68W414yiB+1WXBRTjGV/ImFqDs
hCNF9+Mcxy3pSouFmbe5QkfxGxf7bD2rLqeMa7Ljzyau1bH3dCXmtRVLAwUkk/52
r84OafatqPEuVEuhqwm4lQixJNvkwmagNdbSiEhEgvK6kwSa/aoyI2vVOt/rfuzZ
ru0zAoJskhqDt9LXPMo82SiXwtVZRVbPCid0dBsgdhNcPhJGbhL6f2LMI56io0VT
IDSgMkkT5YNJt0aDMLie1zP7cRBzvBJvZi0CxASQBiIjeZrVR4s/YqlCTJRYYKAG
ENH+vA8MzuDxEWGBsN19KWRtasHpp9chK14sagrs3XCrxx/ORRubLNfR4hFJizFP
DXq6tGBi6dyZqoDaZdCZFN9r4m90isvz28tcLOnvgoboIv/OT+LCb06fkjC5Lf+r
TGKP76lIE5kcVpmJJHeumZ8PmU+DbTRBM48OdJqgyl495ebLi7yRD0YpJqouVPLJ
dpfH6qEsKAIcvIn9x5btMLfv1PS/LI1pF8miwFKs2GyvVNI490vgotUlunn4RfYN
u4to5CYxu0SkN2tHOsbdTepQuVtua4iz0bF4loywvGeusaDeA+f7ADs1lLkV/fLT
xVaT5UsKa80jbnG4jMa8LYPHZRVgTTwpD3mfG+SEMIFl5vJnknGKkJtzIrXjF3wA
L6SBxJ29lu4wG1Zdaaw7hf6J+8JisJHHPuIidsVSLiHaaid85uxwtXRpRx88lF2h
YPssHeZAW9U7eItAJ6JdHYCnC0X3gXsjRjkT9KrYhZ2jPGg7T9452mcKGJepxQ7b
4T9RXH5zg15sSnBB6Ak9UO0sIWXS1pVLD1nNNz/s/6jmmO5Jdt3VqD0lsg99AO3l
b7xczjTvwexputhw6TbMEMeqLGBAa5vwIQ31LFDPJvZr+6Y+ON0nPEtHThFmTGBj
nEALI5mUSE5OEM1ltjB3bezBJjjfv6SbV9GFtPPmdME42pZMQzL8gdlbrr4DW/ke
ZuKKhPnqSs6QNMp0D6ilUsKbzLkL6UK32qmgNEIGR2Ja7A6RjiVJFlEQDlIukdzv
Plnq5XvdJntAiC4lHPXFyI53c0Okm7uO445KIt7JdfI69lNaUfHau9YEYyRpg+pw
YC1w1BVX5E+mr6W4o9A8cdtTNPdHnhnF5+X04siOb4aFq25WQ9Wea/F61anW67QA
IDXqKExLsiz5Ii9yR9WGZ1uc/98swbVdKvw9WhnitRhUyl9fOeN+motUT6t1KGqJ
NCgs3SzAMAfiAXmnO54UPALOGLcLLi8jtBxwfcQCAadz7WZJtXrf+kUrr5P2sZgD
14PTlZF7rXHlxneI1nasLmHmZmRlvy3kTJ6nKzjPI7q+h0D/L1cp1GS/XvvSNBv7
ItKa7qlwGolrnNC3Z8eEfPqyP/mVuPWh0sL8r0ncUETT/a3N8X14xqPytuDXvtqx
UWE9gChVWrQECI3MvZe3ihW1PLAkM8BUG6X1EbktOjSAokplAXXJwOW+acS551EZ
pWxdHM2qovRxkmP2YPG2B94R4vBBiJcUpgm5azLSwUX+44CdBB6wvyjIu5yvJ1xw
oUEjb++snHFOpcca3WuGpr9PT6jlowYZnD7Vdsq6szr8kY2HitFRQ/JzYwxh+IQu
BIde4y4u8ahxxeigxPa4wIQWgqq3NEPefK0jzd6S60mUBMgXkZhbK5izwvWfbzx/
MBKBc7t9UwESNCz6dMvIkyKC3iFxHhVHsMep9oFH0CYlnrpx6eFRbmaV0SkbFQ/e
KeCdMbpEXoVe19iz2ZvDcEeK/ujIvalB0RPwp5EzQ126MrRJRwJXnHrAEflRAtMS
gV+EQqPwt+IvngMO/ybHOaCah7/wwGyGzM9Fguxj3yejKJUmlqyjf3tIsBCQWbGY
HwG1CHQAQHGiUsY3Z70kXs52FUAgHOW3MRxbKbwtNDOGudafQgEUrEn+iAPyZejg
5Gxj8dOrzXrufAgHK/+NIyMii0E3oHfQdZVCyZsk+mIzu/SMXeauY2m9Xb04T1gx
Rv+QOvTDakkLrDOrdpfwv9pn2qCwe/uhYmFKddD+WY9gUWQU3oAmx4S0ynPdxc7i
N0tKCptfNQBOKLSK8GpuVYgF9nPnUyZ+qo4HXplSrPqmKQgJyeEvZ9BqGlN/9R/T
jxUZYB2ZbDTU90572Uu9lwkXW9dio4Kf8VvuILES1Na9oTyUnLQvbPZ29UH6drKa
tcc+HPgRx8fhSev1rvG/1qBxNDa3rX8lmqKkjUVUER36Fz//2rzTVZD4pwSiut/4
9K8/8FthrHkpV+KYR0zEChnZ+eiphBfHnRmsdR2OPSZw+CJqFQGveV1DHinMB2ma
o89DutPwAP9yBSE3kOStR23jFtHMv8udRGqJPiVQZsxvd80oyX8ZTVnIg1RSh2c0
uuM6cQzgV/cVXNQegf49jfMM054O8eTaiJ4w0eO2LDF/J1carrqXtDTxkheENCLN
5mBUnBXZHmPGeR/TJTpAJsD4DEdHLy1nJfHbAFl5Kv4LNmte+LoJ15Fuy01JJ1bf
4TdgztDFy/swiy6hhtXQX0Rwp9TGeCbEsZWtfYD2Mktsh1OaBtBnu7bKKP6dZCNt
QWdA3Euy8eLzLqzF3YABCQ2LJSd1gFaAPkovpnSM3zef0OXSzJYPTRH7L5kXQbnR
J66P8bZary9/Vg9QqJLwk3kAWryVCv6oi9j2G7dG5V7iqI+oj1LNOPogO8inVWeQ
yvqi4QJ8k0NjcjcEYZuythvoCU2KmzN1Ut0okoTuv0N4Wv6BJxNFNeklXxM3J5/p
30Cuhhr8Nr0UNA5fhOoHGLniAmqbQjzt5O4O1VFPES63KCt3gY3aB6SZQBO9OsI6
1Vd3ssOpCROuUnLw5mR9qcNNcgXj/7FYaPc5QMUd2QvTHIbMcSwxCTgPyIOd7clh
LyES2J5a+VqmRcI+IU6MCsC0pIW0AfO7DIleCJBQ8YN+EFc+8qvzwXOa7H/ook90
MrXCJ5lCrpugSnNkxWb8epcwQyJrJtbuDjpnzLvjzTghvw392vQG0CP6+uDiGR42
4MjbN8sLSi17OwgNm5BVrGNxyzoSiRP/Fsx7aw3JbHO/E7WK+gQmYu4Z+7VhjGMB
J1bIZ6KQj+Vl2Fb3Oow5P3rytpagfMcZ3ko8E7xnYqJG8Msv5aUX/g5+1jJjiW85
yjNRGGCmolcDId9R0oqGc/rL5J7eqf10O5DMnIJvUEziZv8O0vNqGr9X/Th4QqrA
WUGd2IbeqfGJ+E55hvJdjN9J9ix8ZBpwOX5ZSsazQ/eLHf1lG0XFBD7rhwCf5xIX
VBgmoTk2eSVi44nMZ47I68v9qGtJD9P2MQoLnZ5kXhk3UrG75pJSkbBT9K0hD1YG
vtr4rJzkWToZSriBl5UIcDdwDdTySQ9dmHvQQn+JCoiCaTxLYxtvSWpXKLaJcJ7y
5BFs/y4hN2q+HX8cWdlq2iOdo/fVPd9UFyafVgTfDovzfO/bl7TsWikDk22GUVTm
yQetivwlVkbd+vn1gZjbjfbbqTISUdd0DkmJVGakL0jCnM4GHbLI7i3wHd8ZvJWl
HvdCihhrcH0uSI7gOdvHl90Bzv76SDF4HXr9edEiDj8wMYjcYeBLk2yalo6z5MIt
yGA6YT7jU3gBTrfZ6aM5qwdXzA5iXdN8pjU20iQOho12iktiAayP7kLbYknIXxSl
6Gn2k5JmBMf3zTKM1ZWL1/vqHt9H+8gizAA0kdUBnWoCAmQb4ppEiSOxtZWWcy1i
07fRVQb3BMbmTmeIB3wn5qKTFW4ncRD32VzhxIgl+nAkarouNHKfBfZQ11BM57E9
QC+VVh+oi4IhZeFvLU4g1COidg2d9zRo250K8sjr8coiRA8eWDq4yR9TT8yk6yzG
c8yXhkjJV4u946H5IFPKf3R6Pdkzp45+ZrH4RYd5sTmA0vlzsdro7ykb9WOaGQQe
/7Zuq+saFM70TENGi2nVrz9JWN6A8v/q+aaeyUU13ghNPAdlYdeAgfhNfAs+hLWT
c3rQyycILKCXd0GU6icKaKkE/27WxKNKhg2vKlg6J2XgFXepfWY5ibg2ithm0Bxa
699k2rf2IwPvZjLWRv8FBjhGyEZWoDZgawHN12s2ZGZa3e0dQAqw1SqAI2sDOfr6
uPxk/oJ0BNk0lYYHw9XOSf8oscf+wSPOU14Q7HhinJzr+oJD5/olaY1iJfI2xC9o
oTQqSk1OimR7R2yecerUsvKTH2tNicnmj10npDBcaMuLWfgTEN+bPCwm2z4QTOmp
5bBalFlZoD+LrBEcgjJAaMlAzll3ann2rlKhCCgpmAqnTTnqlbHrlb6wfcqyd6IZ
4Kd5o1ZbGQ6hzlKRXj2q7MvdUtyx0dfHJ/JNpeLtPktytfQpXFAHsUHblkrQ/6Yd
ZLw6DScJN53jNoSF2m0w1CYmAYJLOEaMOY+D94D7bQjCqUEsIuk/9t66kUTocX4n
iRj8pQiqS3n8ZvqsFUvwV/68rKwjnMKDIwgDjZRMDl4e8+9er+EL3QrzxhO+UYY4
IwQFwuxjuPnNqG2hhs8J3LifWewJpjASKVS0t2ogEoMG1SelzVuwMtABikdxGOZF
ZXKLYYZh1a/VvnW+9QJuOOh0HvcZhzcRKrCRaZ9v3hyYev1uz8/PWsQk5fJw0Eoy
Uy5JxfUFEjtTzDQGKT9UuZDmIOfSehI9M5QBQX5t+/GMPpqrU7xszPzs7zjSSiKJ
YEdFdm+SNCmwBBLuecnJbhar/BUuPpxA78zo86mKOExViNDSDkdA0ad27rOe9XQh
2rKmog/H9hfaN4LUmd4gOJn8FvQKOjHoGy0X6ln3BNZLpcUOpu9GGbXZQSQZB6D7
Tx9HQJwZ8sYdwy7Q/xA3B1r0THCoxFb0FqLpqzbc41NouxMtDSjOFD5az0PvJG5J
E/y7/pN1dY00XE4kKW9+QPZe77Sh9l7oKyDpBRGGxHP3nnI6yMhvEYghdiu1vjUA
aMW5PAnz3RLX1hPB3ELs1hZaKpotqPKH/i98YntwSzN+dMeapJ/4DHpjZrlVL6k3
N5BR7GdpDzLWMSsT99dq1YqmdpMoSGUKz27kiuNkjuZVoosrjpv7qQ1rvn249Kx5
amz9UbCBQXWFt5LhPkvXvwcXwIAuhUuP3MPpt36SBKBU6zQK49YruV4zK3Q+Cqmv
MejOv0p2vkSuPAa6yausjE2Pg/0Z4P6v63QJXPv7b2lQQZo+TQF6ZEKAXUrm5ksp
RKP3ZJeyvWjtm5qkwfII1ozaLP8rNGd6GOOEQxcHNY1/OH+g4LTHXgURqT8LLiNB
lNInlESNGzy5O56mXktPZLy3FI+ufbHN9UQSAbwpILuSgIPG+uVo4rKHH65pdXNv
fwyrUArwXljViOAo6KVwtEUFJK5bU4sWBXlu7nHsaMhvzLij791kb065B/63uEgu
KGfg6oESDPYdbDdIBf13mpwj1NLbSGb1HnBJ1K9++YT+vekXCZ8oL3tyex/wbrPd
RdbLAq5VPWd4HiFEOwPxoAeKvgtXIkm4ryodGXm/goevV8bsZ4XbvmwRPorvdWqy
ntnz8gpFyVzoFctXJHzZ1KmNC70rUxVVO/Mh0oSgmIUczCiUvEONgF1rBcGtAvdb
0GqpSXJUN6e12gJomF6ok5Oyw0UM8x1lYeapb+McbplyZ2YYbiuv/PETy62T3LCg
N2T4RTV2Sz3mRQU7FiE+WL1h3GTqhHWYo+4RRoHVUqgFOjIioDdY57hQQV7gc89s
yEyF9RSchEpdGg/5aorjfp2mMhUEylpCh8Im6/MzMjGAM84zio4kQfB26g5AEw5d
jkKccUBeBxDfv/sF0OO+fCof4gQ+k+doWT8QxQk5X5DelUXWormUZkreNVY0OW5R
lXaghzMy2LJLRezutUT2BPOHtv3iX0AEU/XdHY/rCuLEyn+dT0vLoFKKaPK09sZV
V90bnwkG1usnMBPUdve1viUW4r2Cbp6U09lUo5TaAnFhox9CgdM9JM8Ivcc0SnO4
u/SiUKTL7DMZlR8LnL4BPE6K5LSZ1Rp6KErZ00qOvslqNQ+elX7FRHXeUJ5BCzYN
eCkaXr2auRL4x8eGKzexTIVwuWRWGshV/D/Vk0MWnTcg22wyvacjLDOPZfzQlvHW
Y+9KxkNfgYli4eUrcR6gQC6zYeReX2Jye4ImPQlJ3euX6FrMjjkXYlCNJbX7b5pt
Sl7jyo5Y5S8HT1OkwdlWM4MSTW64gzvXvEk5ZtoIfC62sQZdob/68+UUa3B6rC7L
bVoRAhZ0JRCHqDLPzqGB+4MbkBjY2B0QJNUVAvw8vple3tM5nskmuCMP+0fU0RgZ
2QmZsAP7mYxf6+3+gnKve2POMZpdnonCksyMHsrgLtP5udAH1X/vvz+oWzyb7Wzh
2l9lQFUYXhRPalmK8v+lKnw40fixvN1HPY2ZJ/iHn/PsqXfdmWmqUSmd8DA5Fi65
NjC1Z4nepi4xhxsTF+DuTLBoMhxZSAMrgYz57RrqtHdJvA1nzDzD9yVdK0oXyPE9
f7RB+M48pqve5miAVQqQIXIXKhlrGEhJwGeNthHRBvt7LP6OICFl2dHxuSpsJlBT
tJDOimK98haARr5YjmrScyDyid0egwiaoVTteDplsiQ6bSI0aJBbbmIToqXD9rcv
J41Lr41QbGNhNbSM9f1/93z5p/Csa324THlNMOA1woIygq7d2+r16WrTEDIvp1fC
iTxnC7XhseddOZEBGSYkCVXwlhRayn+8nNxSPIgQWTMjyNwTj08aHTzM+cDP2B48
6ax44dLB6AXByk/npxrgfShj7WffDvxZPu7Ejm0R5ndg9iFnDviArMXT9xddTTH1
RlYV4OPHJmqvrv7dgcjjWvXc9qOEdqvXif5bNuvjNO0CrxFVoHjZ3o/m8GlFOhZs
CG4vQ79EEIAhzjj1CDwGeRrWElQlVARcuUZDKIT8FXGarGGMy17fr7Q+2Lmizr/Y
PZexjYJzVrE7kevAIYb4bRONH1kOouJnv+Q3haOx+O8YzVGOq/IDRFASmuzCz+UX
sLaqK2IvIlPnaNdvCIClKolD4KM1NP4fTKF151oXoSov/Ywp6/qlQOwTkeuvbOp7
xKKv8WUdyMbIlO/rrl4pXQNcTsmoSlh6PNJyqiHk4mooRR8kr1nLesTl/Z/UiVCS
Ac4JtNccyRU8jKE+xlhGEs378bzd140dsqXzQIxwwqT0UrAjRQ5IXL/T2Gxw83zB
TNQUbp4rNDG2dDW4aiHCicgVgiPrc8HY3VIWX3j/JPkmYJPQfixhHbzBYaNEBgQh
IiHgEqoGOwoelhAdyB8VrqQhJsDa6damooCaEcP+nMTOG7DaQp1ohTv4AAlKGGAw
kcWqgni83nSxXhVmyEa7z02DWyQQcyvDekxoN/cLNf5rCXdd41+Yvx3TI7C0zvH+
oI5CVRrATykTwCvFq60AMnJollxSWQjnAW/XFDeWyqpkXxeG2K2uHeaJdkLPG6IA
P2EFx7k/evB6ZmCtF1vXbNAAPMjfCiyl82afz7zhMxlU75f8o6ROuO5kMu6WZoSg
+ArZvrCH70hGRKwg+xoFIIj3JTMW5fz0I+QZWyTeSJKmGiVbDjz8c7TAcxDcvvMc
EdDB9DvdLYMMIX6Qi2+pg3K/DE2UT4gdrbvE6BdyoHN947bdb1mrX6KOmR9aXpcK
+q7N1SvmmtHB6bQUd7Vg6gJDGhHrKrwkzoLSMAWVqy1nmm1wUS7TwdbW7SBW0mCf
/umGUK/8KtZ0H9J3+F49BDa4IaIUZL1Xh9iWTlmV2LwlgAS+J6DOMs9gdyyaMTJS
bAMN6n7Y9/ebkhIJrxDkQZX9rutRg+driTDg14z0c7+5CD5qA2dqTYU8Vhd2AKrh
L9c12Jk5yWLLCfcB7b2tbjhCC1YfowQ9gE3qaQbonaxwhBdn0SLJ5KkBp7g448b2
LOPPSM+i2fLZ8d2GiHi4ElRlIgh70UTkJgPr2vbv5O6BXlAe1qMrOGurqKoHxbPG
YHMO7V8OE8QfR30fKoUXnsZoWIm8J3DlWlmob6Ge9zXWQ9r68GV4MZUsUg/U4LnA
m675HR9iyLqyMakh+Iaqg/PNmt+xXdynwyWKUh4ouq2AO9j0m5j8Be/V/VqTpYwb
4YVnpgsane0RUbEN2CHWh6zLdd8t6yO30vRyAONvoVxYXv12Ycmf5IJGTZtbBM6X
jQnOnxhVO+fsU0ZNHFlhJ1YTQTznCKwbPUGcGYYBfRIwQDufo37ynYtXAnz4wxMb
xIHLmUoa8Y2ojg5YuOTO9GzVGosg46FKx9ar4WkFDG8vAQpsHsPTwMRsWn1fRp/A
OqAB9ZqZ3C9gS1PIUSC24kOFatStP9TzV488pKVQirWUswMG6Q/JH+L3k4GgkaLh
b/3idD/9kKta3JFi5uiMVQmtKmJoBUx98+UkFcB7wUhQrolv9Okd43nIE3muMnm4
sf39MOwWpPZCs98CH9euWFYu7PpehLRN/j9FZ3g3sEsx1tnNgZwIgqkelDhpLVT2
T80P2/Q9r5OZHjhk6EVqRT+0ckfsujOif9bFM5DFJfOFOiBrWaPbXguIuqY9iFLS
TNlf3hzkmlZSuFnRBb6/p/STLwumx3zRUnlbrnWOQCc9Wai4Xax4Jz7XOfu2Ec5h
51Yse5Lpl467KhNfuZYpbaETx7KYCsYDRkzhCK91QCd9J2qyo1jvZ4dhIyI/BtR+
Z9/+yPuBZ/K3O96MVDuEwYxJkt1iuYEjjTP+IweLsCx6sD+79rFM76K1maKnSK3t
5H+DvX4yapwezytp0NApX4NXkXuKV5k+gXMFFHVYlT5Gju1OVbNgqTYmAFZAfZhD
mi+S0vMovYW9UQp/MhosztawYaFjTHDjR4BVkpZrtIdiHVb/RlA+62jyDCD9i9iS
xQfsUlcujf5/La7EfGLRvtlZe8VDhb28Dwhnr0fMYQ/5FL9wVds0MAs3OR/Q4F+N
EVNOlbUlDXhveOzzYE49PAsG6se8O0gu7y7vrY3kK+geukiU0IK54SiLMuSTuI3u
2/NG3pmdTZtLDkdpE3qJsQplJ5hIETtgexvnDJc7dtQJRtwtaM1fSKsJTAQb3oN3
h92w5pvqliLZS/zwWGLnnUnneHB6wTaKgjrvozV9YCLAedX8egvAjJ5XzkcA17U3
DEanZCi0JhdtysVtScZkYZ4ITg7OyEAiVGn+Vd8qJNcg2n59SOGqwIkjkXzFYZ/v
UnfRqLlONO6LgrjE8jzQ+Oth8D3wtrZshQXbkEuYhRAnsMwWx7tSrzt+9N4Ynims
NEe4sQYnyDq6aWf0HYvFwUlCgmdmwZKXTCnwMrpyr3prJerZxbgVEgfMvMH0DE2f
5+QCf3wgcdy7vaYORtb4IcBWQd+EQNeRD5Yj41Srn2eIaOqlYQvjYpjq11Ckv+8o
Zf/Z4CHeLJEP9iBo2X7EsqbJ7nOBo5O+z4VY6GghFGT5kr0hSIaWT4rTcWXSFu5v
loQutiRnMeQ6oR8qCE8bU+c2PpjnL3BJEzjl2CFc3Q+q1Ku4G4a7uYyTWaU5R7U6
NmTUvpuqTkh9mc8YjR/q80mGRy8/c5FxzYpXTAixn0cqCDhQ96pn3x7aelarBUbM
KQ6Tf1TGFu2GEzM8oZDROt8Ypg2+0DEO6uhxauQ+unBfakY8/XWJd7WIhfM/L6sg
cXoEbcdvg3p1AgCIWkH0l4ytHlvEcfKueXO6lj+Wthit+onms3zuSEU1e3QXAvg5
Ya2aXmmsEsaS+lWZEcNqieqzZccC0cm0pglyXpdBDjmUVquDYD2ISSHQM/M4Txvs
DfkcRjhklaRPeODbkEBmMzlOY7VOCf7mZdOv8oqvb37O8S3XuTWlGeLxgs228QpA
hmQVPMKB8Ezy8IGWR6QZPhLZdvYdaHbBwZ2ZokXgd9ogGImW8HgksZNOwWc0nd5A
h62Q5kCijAVBS0NtjgLD0dS7BK3stN9jJBkpTmHPy6pWhlhSsdnIzBqsvip8M/yc
5bXzdngs2pE2s8u+/Xbi0ayM/duBfOqAoWDK9NQY7uftVhRSD29giYpQDyeiKsB7
25BRJ+qJO2IwXnmwqtQBIJAmmcD/g0jpdLAwX3SCqX0aYfHlQI4GRvsBDzozP0gK
ucnjI4XykGNwCs3Y2moaRd2Z5ssKecdTuab1/zUpuYd+HomEeyzTh4cQqe/k+VKH
X0iJJYLf72vsaujMXnQV9OpiBQDHvhpZieRwtF0+ymVqavf2wZz4JGvPQNjLnRSd
5JcV8z/BDrpLLcGEsgw82Wi03ukxlblGSWuV02LlhgiNerhoG8BrzvzerBCxEsSZ
v8CkORVXwP5nwLkxtNQ/kX3edkiaqNCbSNUO12PLsJwgEajKOqdrdsQZE7cdVwhw
dxVsY9UsFWk7XBe2S7iiHBasyNtVWfBxQZIRS9KkX4xGomSpoKi6MoYu31udfyok
qReK8ErV+hDaT7OimUGmInY22RqXXs4FRccWDVLyLydtUhul2QP9NWp3okJRAuh0
E/Qr752LWss00cP/WeQ9NfjZHFPt/pmCxYy8ENzb5uwE87TAkJLDCd6opgaLa6nK
e64CVqGocMftI0baxArP6muzRh2frccpxVxRHYSgHP/WAvMrmqVm03qI65aJQtgU
yW3uheBVGRyhJoYUotyD05u6Y/3GA1+rVqx2muH4yvz7AVfxkMh0WsUCNqnWZUof
a+jcslsahrE+KAMYDsTGLeVHtLKMbpnceL5PQZjngCJTCd17Z469gqMzh9zku3nz
TP93gGy3kXGgV4a4FnkTmZQeviJYe09lmiWErVOreSBMP11vfIhQBkxNF86B6cvr
RvhxJgPjqsbjAVQ82mIeyw8v9sAXxVdAJD3Fbk3w19CmLJnWzCSwie3dwUYtr5Ln
s2WOCRthJDtBD3NGlWeoUtrw459vKmK2Kr5LYMaWnSuQxy/wCOStkiueAf06Mvt4
CWQD1kH4Y0lIovgWOHaUCrS2X7fONCrryzWfbii0au0dgOnbREJgVKry7aJbZu3s
zIEPiS9Kx/f+0rZ8LQOeV55y58za98RniOOhUaOWRrd+3Yq+7u3ueFPaPonFNcdm
IJNvVroanxu7ow8e0iyUHJ2ftNbO46MVWPtIZTPtIp5WZ/W1YDXHkK3wPDlVNOo1
mX+9sIZbCER6I3D/x4uGKEoi5FKc5xAzAjPGwb8GHqPEWfRWLgbb6UrGvGSubza7
QjNX8diQrQKiddi8LxvPUQ5tBM4V6yjbW8e9Jydg8DIOventft2370nyY5sCHkk6
Bs/JHcfjIUMZCS9RKQdyRZsns3Apbcp9+czCp9YEEEJst4/b1tHeruGAT52LoIG6
fAtoC8YMP7ZgBmBY8QgfE+Pa2lcY5/hfeA+muBZrCrKNwIy9jc2IT5VA/XtS3lTI
fTheFl7rjUlEGHbjxLx6eVIz5oZtoF6hu/m/kSi82hbHPCJ3tbO4fyNQGt/tnVEF
rAsIOUnzCZH/YrcnDE4t66tHZgCHUc87nj5mIwRftRLwZmzizLEvhpfZm3/V9uMn
VXO7rpYlv88piR0twP9lJ4okbVfB/4KG4wouSmUKkPns7CxDGA4v4NQvUoYFeSP6
6znzYesw8tWq9H3Crh2OQPpY5bLvQ1ux0vTeXeoqsQ0cImUWgxRswN1NM1SgxtUv
WBlD8x8VSgHS6XcgunF3yFaC2Mf+koC/8PrsL3acOojLRaQwKdm8gmyn7qdO03ZU
AOvUZNmvEGrm+tSuO/qHyYzsL7QVUp2Ob+xYR6X1GqnnlDK03r2ecCMduhulh/dr
N6q0yC7rRegA1bkoMu9fLCFZC4PmNjCywlwxIv5cNkiAR/yT5VugWBKk/TrbAzuF
8Vd1rgH22MNhn6d/GMx4LAJzO4FmHrFGBiJ11z3flstuKrAADzi/MY3i9gYqvQpc
Xcr3rFFDWPDV+010Uem9PZafNMZaT2Gjs39tzwseS97riyy15H01llaP6dwsQ0qB
mha/dDaMN9U3I6LaWyW4Eah9R9jpLs6meKBSKpzNU1aqkxwZlSVGXEgEpY+CN//q
u7F2ZFyTPcyfpFH1+2UBJdsv7jYR4C5f/VriOMmJ+9e6kCDHsb0jRc04XHHDH8JB
F82RozrT9Qkdks6bn2q3s8tLoHGV6TvBCflpWwXIhFAknnpb0xCjCwA1LQ1mOwMI
w8UwhdEoH/h8JbyUmVzPXwercz3PeD/W6sQGBIlraTUyqt0wKmRO4lcP+l9R5gEb
jqnVxNAYibQj30NHCAxD37VwEPYJAQAuuuMNGzTwsZXvyO12j3Bbs34eOLav7Glj
xH4PwWAX0aLh6jm1vueH8ecl3j+KMJuy9+dVe5KCwN06Z12a/7vf6t/qH0FJRv53
3AGCUGB+rD12DmGul7YkixNAl5QioizsYyvwApYtJ4WpQbw9sOGYGxYLOjnDCSZN
i0pq76LWHVUa36bpzhbjDUm7slSMcDuq+k98oQk2lYgZzzG/C552TK10ZwkfiJJ/
g7KVhvWNleFvj/8P2HBKiyOqoKFbr0QyIdNl0548VbuJj679Mpkc7exiZOO2abIb
FzfxLMqwH+4r+5xkAYhdt1bm1bVMFa6CeQdzhl0Spb8HOLQKduN8rSc8ceF098W+
7jaEQkT9t+YvgCZEbkdG0OGK5CLKETkLBq4RlURUFz4ryAmSR2eWsIcmnWuPTwq0
D9gV1MIMAVaXdIebUSWMpj3kM+Hy7t3+iVB83HR/P7oLVdV9B9Q1ut7URnnHSb5i
I4KY3QzE/8Y/vYUGC9i4m9p2EBEDf22FiLt53Gr80BjF8HArONVnuNvCjtzlTNCe
BFcVejiLf57+MPyPlQVrSIZUbdAzcxlZFrGHlvCFwsLxBOyVIYdn4uR+8G2yeKYX
plTxrDsZWQwhJhZQsCj9X2dH2p/wRB+4Fl+JGGXEEzhCQTgGvV8JgPvpuAJy3ggl
zM+HcrqiyahkOCELdjcIyp+LGRi4ZUdP+a4mY8f17YrvSK/xhm9jpSOGGavdtG7X
k2sgUvrz9yEIhhgK5IF8zCuR3GB8+5U/OsGU7Qtlbj3EKyWY1x1i2KiiGKWybwvZ
XhFu1Jdkt9rCnz1vg0hWclO/7CkFfSvuap/0qRCC9c07dhWCc4VwNrf3j5JJ9NrR
Z6D3auGK2WEfqE0X1A5szfpVJMt4aNeTh1u5wMY7s33TJ4RNiioZpDCbW5y9OsE7
8EliOOylWtomSNq2eUoT9ATvWVtkHYKk80HSR443N9QzRgsKx0HBhch/+WxuB2hz
ShzJrVUsbHdjNo+wA48Nqtj1VXFSfmpwzTcWVDikvOityzMtTmY3K8j01Qll3v45
DObtcdEDMKJsppR9q2ZenH9ly7wjeWoyRRfkTqeXWkdlthqYW064xWrgRbmausbl
NFTioOUqJKosYy/1CnAaWfXwuUd2QXZJFNZUGG/7iCUQDtaup1JKQZe9L3tE7fI4
2lu05Ph2IZp5FKI/2eMxseySJGGmn4YzG2IAsTg+Yj5kZWI6820v8qU8QmL2vdOM
Pc/L2DuQjikV6qcA7uVaLy4W44dZ9980YPTqlSSq9LlPlVWRUh6Bo6bpLIU248/a
lASIQ/sGUxGAxNUZTsQfMg9av0mE+4nhBYPp4jVjmBg4KBW8fyQvYlkMN2aDZuku
VuRO7rlKKsk2SfW4fPkDpRZIsxWAUa7Q/d/x0uFn+EOCrZ1cs8l5ngIKo/hKqreP
P6DPF9FsReBBVT45YiAIozadODuA+p8lP5oAwtJxj7iHw97J+Nds3lwgH3081v7+
jnAvdvvZHwFREu6nuxPe3cHSsB1ypROUGEe2CgpuD27sT9SShYG9UU9Z2Bvy7We/
j4Z5djXo9ARawgCgbeQ7eQiN2b5bks7ZphZ9TyglCPLH9KPazMnscjjHX6qWJnxj
FDdith3a6xzb+Bpc0gi//asKjKEqd6pnY2ShFqp3nCuxqdhyGinW1VMoOe0Xj0Vk
2qPboZYSFgpJ1GOnQwwvwDAXSjo9GDU+bbk7Am8zh9H67xDNhulyR21qg4BtKbde
uozMmzbkPJaQXymMcDK/usvxdsVEJ+TvemfiYlSKq1tuuG/AY6RdqktTD+bpGPOi
TwWhHMnOLW4i09Y2hADGNyJ3vqECoPJQC5/UXL7amtpZVbBhJMF2mIYNStcvEAjP
lPkEwCKW4kynHPsSSEJaFRQ57XTETIG8EfviCkRx+OZSvIdF2c/ZHvSTrC+kKQBY
3uzUeFu6ghi5K5dle/KeoY8fGvzIFzPsEjfpzKBRBkdZ8Zt+L4lVYLyIjRs5dsYk
bGynkFI5UjDhl/lcFcokUkW1tDwyetHA7ySCqLN28T61EgsH4HSwQ8AXW3Evf+ZV
nxHfIUPftHPhGTmBMQ0+DOll6a4Qab+OEorzKHDIQlemXxDsVvP0qTi7MBwMpcs8
WjGJJYqqSgPIbhGEHHP+/bTtsvjgk1qF378bwGPvtDLlIHCbxS3garNPwgNIxaid
P2iVi4sL/yNREQdKa7eMXnd7BrL3u+rC2Sj8/BUle6CwzAAo1zwDJGWw2DQHNtoE
sT+hvlh9BXabWaaG2BSYRT2PYTpe9t7SWGcIXKBWMiN8Ug1aIyBr9uQ9D0Z4XtId
7p5+BOi5y/u2im2hvMQq9zRW/HyUKwtCM1QURRobAflg8xIYEuSQ+QQWuKR41QtQ
BCi1L84GJmm0CGi9FsLptVka7lY7DSw2NmKsewoK9dFAZj0EXTXmBe7P1unxWoUC
Q1g0arge8CewHKa+vlBrbb8bjKkkrhMdj7BQI2hD4a3s7w3yknAePO1e1PLeeC2K
dgmkGeWBcezQp3V1hKlYD0bFiDuVs+nosm1ASqsRV/cLzHnBnKj1devCiNc+J8St
NHNHWyS9gRpJdsXopOCNYf68DLZ0zXStCBT1GLAPCPnDaJh40IaYbUXRGhXzOP2b
U0xF95+QOpHzltj/RnkTWQV3ymHVgJcraSSPRzgYpXZSIozY4mZLldN+IZHnXTCm
ZopOoUITjjJ2/INaVQakvk1DrRSRwmrqjVZOT/2Pp7AYiXycXqR4j5eaK7uMqmPn
D0Xtk3tCzdEVcCj1m9dChnJbXtOPpWrVF2AhxsXfONUpywBmpruySqoSv0iUlxHn
oJdnSqCJA7W1L/XcMpWClyCi7K4OS+F1hOFzbFIKI/zEXKTsxpZ5/ju9+gFtiplF
WSIij0nigUoKgR9rFocTiJigdGtcU3a5ORVRzK9LCrAr3nNT4x8u8s7YSbT0rehf
o36WXx9ZViZbWSiePuX3XOesP9o0LwA8GkRadspcGFzwKotjcI7RzfCFV6DxfppW
BIiLdxtQWywvhbDMGDHZX1lRbRb+oAAOMmzOFridokySbB35MLCrYCkBgmvI0cai
pWzy7uWLNOsDVMVeyEXo7I+oB/nqFYRye0rgwVJvT1uHXIoBfSGrhinKOhsKqhnz
C4iDZC4WfuZbxRB0CysPkDzAG8Edeh92pGjQOqT+nyejbN2IxV2RPBwv/WF3CJqk
dBv+XLhjqqoanidQ2/9CW2wf8sRd96RSEtd8QS+ublTtRgsJBMjHXrnFSsOIixYm
2Rx6LFeviJoEFxganEk4qPcfOBUf6eUXPGmRP2T0btoxgg7p5KmawTVMS6Auz5qY
wT51jy9mh7A8HLOupYX6tXVUmBzcstcUHUrS8SilBhSnd0nOLP2tF/yU3x/5B/o4
bPv2zQrcESD6PwJZEO/8pCG0AkGvEjdleDqi6CgSYo1nQzW0vOKa34mF/e7SuaZP
WJwRmTANjvgD6o0AWgdrzNMN7sDO+/e2zjtkfgYtAbB/9ZeRvMRbZMnohLTj1EMb
c1Mf+ZtDILBBPTvdyWlfioFPpNlY53X+OMmij9u2Z8EU5aMqTe1FrrmAhLcUzi+B
KRwDl3qMRkbsmOUBYDChr037KXoF8KaMfiUV7jWPlxzFBLNZN3HX3BAIFqAq2NvW
I3ABEvLMoDh5t4ra+OHQITTLiL2w8aB3hTE20lS7aXbgCFMetqALP1h/19ZAh8dj
1XZOl5wldVKqWm35tUPHxZqkPJe9V1i+zbB07I9PySXuc8118YZcK9zTumW6y4VJ
R7xWRD0/p8FaW0DvZiejStZ+P9FLJwFdchTlzn/OkH7udS4APP2QQjQ15c9fCLof
1CyOEFPUcNI69VDzbjAvons9VD/JkFGTUhEcuKvTD1kXu8ytwGmxCQ4RhWlKlaNh
Sq0j3GiBdxCKIPqiZJN6HQ3lZWlklraEDXeomHMwvYiIddh89Mi6hLrLGW3L5HqZ
+6Nhq4SX/w6gCoxLsXGAvTpVugjTCPleDuKwh08ODiA7/h1KL+HSK2MlWxT0tJWZ
Mc59cLdG1crrx1dsth3zDW9EN3v6VilQ/yPGq8c57X47FZ2Kc8bWFeBY++j9P30R
KwbrqWKoxLZNJxmFLX+ZoMbJPCvaVI6GJKQ3slk1n6p9+DorAms7iEFtuVGKm6iT
2LM4E3AjCBtlHWTCFiXzRCq91aKqqJjI9ec8AgXHR9lKZ/32ebkOEnLwXPEri0QT
XQwuP8NRYWUyBvVA4XUiww19z3xDpf3ipkA+46Y47pOXN07HH4pQdN18cOEkEQVa
wiAjxMrXevLu783b6mKUv5Se0hwY146WY6amDJ+fzivLFeszCnz9gynjs8ojI2ph
Q8ySsj0lVrQo0vwqiwMF8PRmI+1y+9/W5xat9wNgTJkXTOcZu9IPkdcy6TbYV9MO
6EJ5PpxpJMMbW0TPcv2UBMMRB5t2uYiA9Iy+Yljl/tWlz4M+wzJROr1ZZACtB2u2
Lzdsr1C86SjK8JG7Pg1Iq2VjP5Dcrc4j4OLPgasktVccqiChvWDE5WymNBmQKs5Q
Bp6C3nHhq044A+d3idZGIVCB9MShfe+7JDqK3BwC1RABTV8+IqMjRDq/2jtLBMzt
wWCYghigAmLttWV4kKuUpDLqSOotYsVgNrIYSQ121967MvBXplsPZ+rQVrCYOZ13
qRZDyNqU94cLMLKoE/djx1T/yLBLLkpsdQXLBgTwt8T5wHwwTbUoLntmbSm7AfI5
/znTaKl/iGYGpVEvwMgqXu6xn2s0Id22f6Pf5UeCqEgI81fo/Xfqjf1NUxGG/C5p
fkk7g7trRd8Pndgm0mZLWvpMEchGpksT0+R6ojmNfEJqR6QTRTpVcP1OVkauegZe
keeckEZtACHQt80nolGYQU+zye5WmZe1deM72/+7qBLBcNiZEESRVcqvYPejtoNS
PO79KA5aPVOz0+fOpB4KqmitDs11wDHU2eQ4APtdmLFAL7GfBOjvRq6mRoUp9qq2
sy8v2VfA+D1TVXguaMLFkKy9U4I/X3MYGGqFjty/rJI0haama8qRhjTrfAPpVhWw
hXv2k0/A482Pup7Hv+YqnK72RfrHlDGd5gf3lOe+imkLFSYDTjuym8y8YZ0t7DxW
O+KdNwJBOGY1q0nrzkGwu+H4E4lhlYMhGNklRjMmjdz8VcezxzidOYtm7fInIvbD
81P5CN/+sIU4SefPPGNJlLVzxGEXWWOC0X8QyGdKXmptKY3pJ5+2ThX3dORCHIRl
eoCY9Kga5/amr5acSK17B+wmDFv1OSRivHHTVAKwRHCpCZ6xfJ/W6smHYQaN6buO
LFXaqkDKPqbw5gmhjkCa/w2E4bnEyAlCWck+kPxc9W5ptPyswb8V9VbiBVsox8Cd
f+bDbksWJXMaTMJ7PtB5+gkkgdBE5QTJZppl0lyREWvkv4mG4rBihhEzgG5CEvY8
SQj+UEMcPRjiUZGmwy45QFoaCUCahBshtzf1tAnV57yZ30TcdELFpsF6w+eFrnUF
nLJAgDXwFZQyeFAx79AmzI2Fg04qQnwOMjxYz+qz79yxiUOlm5ewZEcg0FG+yOVa
PD6Sb8lmtZQ+7WVvg4vtqScT20MBrK0/qAWbHoNmidookCtHKY8vTspnlAKrrdiH
9XBuMWlbLQJ0Q0iSY3CF18w2gx/VMyP86Ake+IioRs65td5jE6qOMShGyPo/vBM0
qWz7VsgRWumTHtODzTAoESO9iJws8omLdNVVkoqCqQbP1mPVRJvGEpQsUfh6qgJ9
solTBHiNH1ogg1ixHXU415zV5ygwXcQOevQxQwnYZAJFoEqVZ/E8wM2d/s3pxLws
0vuyR1CpRm8kJYzRGZvvgqWS/8QQv9dl4Zdpqof/YStb01651b03uP9IQfFNZRIS
K/Ate+8BqXcnGLFJzNKnyfdQFZTyt4iADOzuwYMxJczqlDrEFEI9D3azX3A54wme
myQDnh3i6s01w2gdK90eG3oy/I5xnHIbxvwvjE412lIzwbywNfHcXnkNQQOk7eYZ
hCjC+Wdr1cTEld6XWixbP+L/p21jwyosvPg4z4dHJLEIoi6iTl3h6yyEBbOaiVD6
T56mid3IlKqONmiJZatrM0KO++95RjwSD1VcKuR2XdD79x+Lg46jLqp9FYhYPTeb
VckYR5E/9uL273HnPx8LAJMLUrV4/8JAem3WjEvC3EyRuGI2MNOBYerO2unAJLHX
LOoDgnMIw3evOA5uR8Cp+dmfhDsXYtFWD7KKGBo9Dl9xD9insNibziKu61kKGX1r
wkDrUITezxAfNASo9nK8eURpH+NhpYtsyKakMpqolVaGlMGHAK0ov3RgE6gZjLwg
WWNGsc4/CLrZREmTuP2uOA43yFvhUK4T34Rpe8YO1AT5mPwFHo/T42Ie53nGh9yX
d02adZL26ijwXEiuZ1NBXmIV6yFMQU35D/ihGeTq1K9TWziKwE7gDrS2yswMy3D2
9I+jG8ZBWJkm6tD6rODn58h9wGcKhl0XzR2g5XXB+zXDc8JZ++z9nJ4bwPb6XyT1
B4j2Pj7h32sPuv1mVnwdMaBazMva4pL2i1KyHu7IDiq5JtY0/qucAD5Ct4ay/h6W
JYXIgzoe9xKV3yXPh9dLPtSLOcIDVpdeA0ZJ0Sa/EtjZgYlnLN+c4jzIXuR6cPx5
siSI9KUk23cCMK8BGruMZr9mEablcVr9QZNbMWBL7tcqE4/kqRHlLaerEm5lzTou
2ddNIJz8y2bYZv4oBskYAFSGtNmcNKLiqFdA2QDs8UzKCwitnYReiHcdYgvN299y
VJJV4BJpw2/91bgSpfIekSG4D4KxZUJjvFgoPvsd6GIGgFZNuL4stGH8jLzPK/cb
WLdhADvwuNwzjqj8rpceao0AcD3KWCHh/xgAnanKA5qP7BjTFu7VJ2O+qBVSmfmW
MEhcvTckWXF58CJL181ac2MpXIe538Fa4o8zSHO9eRLkeQIusvQUjK7Wqmi7ngpf
VoOH9jzFD8MtYyKnqFml93fU1O9X6M8P1mBiJsh7C292yuo+/vIUYT590BbtqlJq
8lQEfU0ww9e+N855sj3q83xXQnw7E0HHjbzx6t6mpHzuaQZyrWQ+Up8OyV6uezWD
/5GscGDKqkC45JRtCNzv7bSZp/2pDWV4Y8rLcw2G39tx4HnBEAdAtRW4CcfZzIWQ
1esIqq5zbshIhO0gQwzFYaympA16RZWhSpySEEPENlByizseMkVxvnoH4PS2t9Jw
YW0PmbkUM9ev/XNtP6adxsvw6EyNqCtKJOiBnhQH/lXLd6AtJE0WBoezbh6srSx5
BzbiHJFxP2GFopBSpG1O9TTCtLk7XnnTwQ7Rc7hySXRKuznUMsipuSOvrDJIMRN5
v/xYeGMN+kJNTpkKdek9I4JujqjMW/Oy4pmdjBSpoef/IRpD4z62Ph2bZyP63S8q
GCTr+bHAFHDTg9FUdnQvVe/WPPrkl2lgLm4AynbkhjFRWi/j10hGmkGPwlko5Vuq
avfpjyR+P4sHIDphd+iMnq7Q0jCbP67KgqiK0A9X/uBaPY5E/BtTujkrXEKTqop+
7GcTp5GxklKZ/In5wYeBj9EjIEXd2IYXgokGuDTMRVBx/W9v7njCtCDMkvewtzYy
CMI8C/pphYEO5QPDuIMeiepERwtRHtPbbycLemYx6RbEKs6HcAz2BHDJInn3w8MM
tI+bWATTL89TpPS1rF/V5bfhy9wLzdOe0DlLDntmXfBS0967Ecg3DMdhilqyglRR
yC/YoUNKTWQQaCN3go9ZCKBOpsp92FGlzL5WnCoNC8kcXo6y2DG+6Sr6NxxOLOvJ
0hG24ZMNXPK3HKOSakfWtpHp6Dcb8RpM8GasF/8oRIocAuo7dbUQQ5fzoee+Rky/
9FPk7OrB23M+1DtyLrNRUzFgJmMqwyEuk1dUaIGMyZOUg6G0zroVzzd1rG3HOl5q
g7m/AFw+nm9XGLJ6+1azEn+7UKxsdSt8CCi2URka55EzsuG5jp1AKR4Bcc7LWG33
t0+d0baA+H3x5cMPSo8oeK2Ivh6oEyV7gmvcvhj2b/cdcQxv3RHDHnUUK7bgpm5/
ifYnohk/EGx8h4mNVMbDB7B1NQS9/wOCFxBHST8Dv7d5RY04yDi3l8p4+SEvrwJa
8tQXGA5C2Ikn5ckPAEJ7LzcepxrNCuGqz4AgFomyomIiUzuJT+gxIhfxUJIT+5+o
iewx6uJcKSy7PCxSkD1P3va++2NIrlqN7xhIXmSw0mlVhIRGJDFoHu4EHggB4+6I
9q3COU+8yNNY0M1cO9vNLvcoudOiX2t3lsudRTQorL+5uYZB6T6sfVvKgwo0gpX9
Doub4YSoLlZCXKs0JJQGuYn8yJy4N00SFUzwIRj3ryhmK/scefZiZgbQixzxDFGE
k8FstwnogjNCYWljiL5nuqei7o+1r7azpDMpZoBrNlvmRX/yP2eh3e/3Ukx71HkX
o0bxBRa41eI948ZH8npKE2/4DMp9w3s+T31Eokz8TRTW1KTNWQ3CfIU1DayaPKYF
QhhMzIvTIeJIdNPWQrWkRXYZAXCmjkMCd7BcztHo6pJRhqG4CcoYWXjjJZdgHvNB
JTqZgOFa+MfiXCWBeikzne4BMbJjazdX23unogJc5S4p1RMF5W6Mhs9r8tQTqUU7
8c4/0fxDtt6pSgyX8o1h673gkzdmh5v032kYG9vvJ3euxAxpZj3B/gM3DLYcSgo1
hEA6n7C/cw76nbRchut1bYwCkgWa/ksXcn3gvC5v325nxeSQV02kHuKredad3XVm
U3o+Fdj0Sd0b85TbVukuXORarKu++KuxixKgwjQSOeEfjewWH9ZOS4ZlwGuSy9B2
PuZnwhE+B8Wfcxwf3pTfkfDU9h1v53/WYb3ZtFOyi2s1kgDVt5fqth10By6RXmdn
9O8AU6+7xLW9GdV5n1g8D5sFZfgZKfibztCW1o2CriNxk8vkPY6FwGhzC/h7JKtZ
LDP1evu2U6jBV4O2elZ1931TjaCxBPaBXfu4Nn+4p/nxm45iAFPOu4W5VCxtqwRm
Z73l2ZadZfCGgF9tU5K8RDZE4JSmYrD+Zm74Gv85+5EZtqsJlNqYfHPNZcK8RAXx
mC05sP7+8gYjyqQW4oQwdG7TJlH62f//bf1WLkjBZateJTyhohNGM21LI15dFIuP
vF2uoFwBuCxipWgDzAUkDZdtwrLG+Rp3eMNTPpXtTMfq0W+kr0RZflSpAnDcL9qD
dwdaXQcKzwLrt4GarPr6X0d355uB5AYFpHmbp60Y7RT8W+FMdo9bI5UIJvZvQiEV
/Z019x8MvE2Bc9w9BBwkr0nsudxn0U1gMTURuZFv+lkyEOzXnROIYwoEBNWTGR9R
/9GyVkav/Tdz0w4D+gq71k1aSr7JGbmwditdVI/8NE9RV92aAf4IDe8mczjXYHf7
wLyj2KEG62684F9I/kt+oUxhiM04KKLWYjm7Yzof2JX+hqDjQgERR4ZtfNEGcu0q
sxaz3B0MkzEsYIcHrA+WVFl0zmpU7sF0qu+1f6BwY/z+fqqZWLryKIUOwEs9TRfH
qPu2dycBaBy+91rfo6zl4BvMaDog4KtTMsj+d/YS68GhG1sHDkbUkoIt0rJ23QB6
Ux768pr/lwXjLG+ifkXRV4IJ1hrNXZ7Pvn7mfjhfcfO8rihsVJp3fXKUbnTuvrGK
Mf1WPqJXQnPiNS8Wq//ilhHLbwkgoSmqiUqAjA23QOgcah9OZ2Pr3WllKcieLtAj
TqiC/Bh7RizlA9rYf2DuVBJ8OyPqhRm7L51defhhCV7yCPVL9iK4bMah4r4cpIyC
C+vxuZUSvXlol2/EEpC6/G8z12PO03fWZFJyLg0ZkMWmHfB/t4PS0GEWL/N6yHPG
DGE3vq8cNUfzsC69gNB6zgDmmzjd2dzgHJ/qlkL3/eCFmdICo+Bt7yPwBEPOjyPG
M8RD+sLIILXAIskSVHgI5fKn8wCW5G/qvb8w+i9QNnYDB8Kk3+Mu1T/SXgaoP87a
VcZv4IIFaSawM6ZD1n2HlBk7uCWBWVyrH9tLG14RkvZtEOmf4YBYwCuZ/6xL9XZE
rr4ItmnCTi8GTJv4g4Me3plmOREA5t8SxfZz2BCFmUFRFVtcE3G9n0tnJiDxIvzB
JBpnvDa8IuAPNjrOoUsVEZ5Ynmba0rsZJZ7ngopOt1ejnlCSTO9LqxZnAW+OTh7/
UNnv1Vb7RIKuMpdU2tKU6XoKu2yIBO4+Ps55q7ryc8jLPr5ukCWlYHhWY+WO6BtD
q69QPh7bwNE0r3aj59idYQH8h5N/IYnGMKX77DZe0AkhzhHz6YSfEDw1Kg3n7pGV
aXg9I1jXjhXFZNpd96s1XRczCqIOcGFdZ3EyWtgHpY1A8RVyFc7eSmMAZcAosevh
uY9C9rZkg2PnUpSB7TSESPMNHN7IzsCRCn6oHlT0CkPiBxSt+5bbk/ahG5cmSMQv
mjpVWGiOkVnY22VYEwqw51J+2PWKjicS0q33cRp4wzgmijoC8fJt0+qgHbvsRdE1
qMkIsUu92W0U9/y2nMYrFlGl3MIt3d6rgY7uYWDDO92kDgVgLILX7cgftGtzlrJO
o4mu7tDC4S6TRkCTBc+GP2v5+cNvuxXYE+HFvsQOlO/Gl13aPDwq3aoCMeCeVsxx
StZDAfsDIGoc1h3o5ZorWcBMCQ/7aLJrYxynq3LfVmUkUe631WU88IZCIMODv8uR
/BRdwI26w7RY/3rF8tF1eps2SfjDNRVvSVi9Hjq86nwqh7+LyF+cbXC1SN1bX70Y
2IqBL0LcGhJD4SGVzYYCb9CwLkEJ3oT1NjpL92jXRvO8XlqT/3rJ0wlUqro808R9
satdnXJSR0UyTiYss8vYBH3YM+l+8c9DVaO5Ps1IZ/I1sXl8rrFBeqRXFWBpH5tB
BKPUkbgPtfGC3sOuWE61EuAWNeypT8Pdl8hIfsU+uoCHFvgzeqXCzwkpT5aYEvfp
6Lblmwr85DhawevC2vu5/rVnc8UhibpN7nrrvGrJP6rKutUminHiNpS0bIo3wRlA
33LocM6SLJ0Xt5UZNJ433c+zJtrTYgUgfuPWVHeTDtKx47qKNeL2xUBpzanEwp3X
g+u+/mGQMLfD7+RqPskAGwtUNOnnmN0+cqKtahqr/zBSgAAnn0w6XW2G4srQsu5R
QY3RMXV90S6Y+VANdtgFe+7g8OGF3GK/aolomfwX0KkaEeu2mof7Ay08mB7MtRlJ
f+i2N7cMpVL7Ce5olObYgrePitBIhxm9KGOycIikGpRxR0TgpU6ZB/y89I/mkcNj
jSlNTwmf2N7dz//PyT8jZC2zN1dyGfRgusrtcTWtHdPiiJxr3CJomnazvIZEMEDJ
mxZ1L1cL/R19+HM/GLoF+GJ9cOg5TbIncit/LnY1xfPgrnl4DIIKKGiu1si5jwaQ
xcQcfUQRwnk3JQAg+kfZ6QQpYcOLZTaKp7DTefNRjO+Aa4kDcel3ODoGXr3HFLdd
j7kBWQXcKMuvXiM3EhRkqkI9M35uu78wdSda/ZYczX1A1l5x/TSZbMW+QsjctTQl
MB6e5urQ0O4Sp4scuKSW7BKG7P1As7ZjqvtCpQRv7Lpe3j/GrEHTq5RYcEykDhro
WPeuEjcyJSkIefG1C5NY3l8T15WBwrjjTgK4cq74vus9WS/aPJkJdhNLMIgc6Uwr
y6JNL+g5lwg/+UcPSEp+UuwDMHxE/r5J1Pjpqig1dLE8LkZgRJV7lqRGDDrZLXaM
Tl0wPcLPV3Lg5gdyEavbCPMOfaAAmSBTUiBxJvlbJQFDuWgybQxKc2aA6Wy/CirD
vR4VJCQ2s+zb3jE+QaAx/EDc4bG+J4PCv0PC5oWcn7FP8Llph9LQUWRGNgYt4MWy
vDe7jza1KdJjGVHeWkmzjrOqQiybsWJgu+JbZuQUwyr1zm4YtBarMAQYFeRCbNVw
30UMeYjkjrbCMDAoIGkfoXFIppkUw4qUG9tXmXH2I4nXcC1CQAcdwsddaXqofMDg
/DJhed67QwMmhgGaMzNpe3bzmrQ1IKR33g1vqQhDNhOew4sbAixBb0AU8SRGZXME
t25WU8o8KD+NTJ1r7QA/1e0btsHMDtd3EjR+OKfUZfVf5jzaFmdvyBWrOfPBCS46
btLOJywEBVy8gAxqkVM4Q8lq7qFNk4Tkebg0d6zcnPmSyU2wXkpX8tdhSdZ8UyfE
F/ZQIbzY/E97h5OO2F2XwrgvEho04zFCCSbEd44R36TFSurt5AI0W3aJ4+kPLF8J
ThecgdJhezqxD6uAysJdgQv40RJVXClSv7YxNvYurGkUbzkI2nCA+smcIE6DOi7Q
9u6OO5AMVtlr+j/hxlpwmyjOMYDNoFHj6v3mpP9qhNbycmLwlTuuO2EQWxTG09k3
H/AGOsjK62KhGtd8n9mfqpG9lCEt88zGYRTqNNhLUh6cafbqLLbZCNyVlIdwnL8x
8drO9Bnch5KRZodQwBxEbCfkhNE7EDlXc2ZWM81tjQa26Ig0oFqs3aDy/2f25nz8
qbpLs8iEO/5xOIHTjfpRwXCjsCmAbhDs0oEmHghaweYMjzr9JdqsxTr8Dox/twdf
iZjtGPA/HdU/F21mh/P0FCd/xDf3UappFxjveTQdo8boeAoG+4XAuy97brz3lbb1
kBFhOubcyrfNM50JHxFA4CceF5Yl0uPOGxP0/CzOh2VpHE7Xt+E0HnNG7DpwHnVr
BHhCUKL1btTh/1B0tOgN31d3vSzmgl32F/dKCqhWkkk92+hMIuGYGxtoXzWTaIjE
VhJTdZ3xMW4kHSYataUdKod5FJN9oKU/u0WbuYCWhaMtNnWv9xJFkHd75uSVoYtq
6YFcRTeEkGxQTYH2/iSiUJNc3aaeYt86H4nGFXYIczdqCBHxuYUK2ovYEKj0EWSX
X6RY87Re0kGwnbnkpHkPOVPYKsFfw8yCX2Lc2M2hfnfArtZg7aEgi2e9CHvqETIp
yaH9E7woVKHSea+JA36LAQOORaCOzExFi9vhnJGXAekTEQ/Qsvp2B8SNE5vUpvOh
VD4HC67XXDmbK6aAe1hvO0HHn6sRbYyoZ8gLoxw3gUFc9XCyPEha9oRs3x8ZB8fe
lNZxCOTTLf7DgQxY2QszVI1n3Ydh6B20pPJTI/o3+68zmiZ/OLBb7VVvYd0M3bMS
boWyg3Yiy3cLO0zoJeoZUHEtwf+oLx7nkVgSB5eg2ghBzVnAwEP8tOMeOkG5zwNS
oe9nqCE+a70jvod0fgRGvqxPPEoWsbh5n2bH0YNIvPqUZfWOrQXU3QSNDxAQJduT
kYtNHWTBKLYOEqUo435FHfUIZfuZdA9sd0FiGXbPhd+5dqWDS7VreWpeBHBV15fe
YpVnjNVGr4PJ8dO3fS1dvgO/tRiCwa0iIaEh9n3HY0Hq5+AEq4tNFcDO4lSvbHz3
AmezkmPM653t8ONd7fCMefOPPHo3exevlhs5+YNGYiDWbpXWq6XMI+ZnNirA0m9M
W/petS9abzITyyLt/cEWxioZ4przblo5EflQmetYdBOutIfyNKsheqnIXkULB0K9
EOggODwHNQ4yRcMadpbkqbYhKb1fTqETjGnq13e7xYZ8v36fh5BjsiiRyFU958i3
1b7kXgiZPcOtvDOTtsH+krnE3Oa41vJm+kQmixPjPZXdcZ8D4cG60oVNPLAjkBSu
jp1XRfQKYc9nSxQWfXYRtJFSGZXP1+sIN9N/3SshWUxZwhJ4EMkWhvidS2E3Xt+p
cnXBdWGPevuY5bJGdQP/3v8/RRPHRBoRQoiu6rOatcKnSSBx2oomksseEHGAf18c
tUtj+GuvNjHTsJyNBwJBEsKYYEPbH5aRqnWQnliiCj5ZHVIkYfrBQs3uBuqocNFh
w6awpxQww12uFPdyt0l15kEG5cYr6KH/c2rH1O6izNjL+rB6wCX9OOrLs9Ay7T5D
TwSK5ZpCY22borjW30ymWtEqiKzKMOTln7HPfzdUQGa4BatEhLOI+QevZnyvew3K
D0n63cCGgITInByYxLcqn5k4Pvh3EyqwbUX4qLz3bWGjO98YqIet4e0oLfK2ROKk
1yrnGJTLU0m/iGvo0geZRPD2iAwungZRaSxVHcIB1jsjYQaa0XI4didUa15FBoKU
aQ+KZUenFE39++X44rGwceHGVam91PTAjN8NLpLoVopxpFYGUAzJSYbd4+WC/Kih
ZxWzlpmp18zgDTK2FPx2TSKp8sa7qYmVP42FUvCjapHyCJRXfjwuv+niVR8R3cnv
6Anj4tp5JfJi7OB3inkK8jeMNQsClkQpwdNEKP8DO/0LmmkTdzPAzFijbBfNTMkJ
mCXrG/WFRYpdqtnYrFWiNbTrzGRkfmgo2NRdrLPnmFP+j1pAWxOjNr2YYpZLWi6f
QF9NNSOEhaaOFzLavl4PZJW1R7n9osVn3zyPKvSoyyUnts7/myNNSIdcU5KR+cWi
urasYorJSaQjIKBIUodbcRSVWXamAPjdbmkVA38EoGss83odCcNpOU3hn+zdf8M/
gSktn2CcIUUR9g/uUwfh+7W99a9waPNmZ8o1Uk9R+wRky2KU730hErLjki5xqyDO
gn+MPSruaD4YH7fGp6TGHwJ47RaFTRMaLfBSDwJ43aOuNU520sw4somCKcOZYGaM
1vtKAzyctrtLm1X4+bcxcFIURHXoavDEeamHmRTK3180MXAAU1EeW7/QRLzDn4xg
U6zta1FQLmlDTCaHg0i+9t/fjG+2MmuYE6H1DysvNdk24DhLHNU36B+1hXdKfq1x
V4a7da0Gz+cx0mHMMi1ZjmkBQ57D3OpdIhdcD6nUfdQL3oL4huqYwE1Gjtl+A+5q
cDTff+N6pT4sfvRQi2hvyWuTYlySnl5gXPfUbWvOuEwlBwZfrLUmmSKr2/yCaVnL
G2WsOOZ3f8yffv3NR+3O0qKWh6yglSrNNR4+FrgM04LdrpcFDrz9684bZ0Z7NKca
Ee5IcO0xfhOgPH2JJDyojWQuXmbgHJkLOYiIeJFVf60+/ajr23Rl/C8UbGPXMT84
3bVcC/DyPpJi6RsXwAVd5AVNAMyNIWNEDRtRlZTuMLUrLnUR+vVQirdjZlStHjLp
fQL9A4x4AESHhv5qQnGt7VE+f3c7eqS0h5COYIhu91+zlKflKRstSP/kKXxSdcoo
wupi3SsfXXxG3ovzUSwrSy23ZusFzcwXnqeh6XICOeG5lxcPdESGQNfNYbtsTtPv
0pkyeafBzy/cRUMVbWOZZt/GLwhYRiVo0UKtpa7PbXWv5y6rf12Eo+jiwylv1VMo
j4GTy1qXUi3WVsxzagN5yz/oX1/BvKMevRhX2OGoSeHgCCurdQm71qAieTTOGEXg
RKDaZ3yASXShoGdeBoLuxl9ik4WkbXEFT6W6egDMb+A0XSUOrLhx/ORbxoBaIjyW
ZIphXkYOzcbtSdHXZxRo8or9coSqdIkDA74gInxU8RlSJG3lxYj5/nyJlDg51vIm
WlO+wsbC+o8cFrpzPfkaobJGgb+kjA6rP40ocQ7lz3g+272Qvn+EYa3gCSC0/wbD
rCdnwTnr0sdZUCl3EgccQNEZe9bSlRRKoBt7ChZa6AiQNKDFPo6YCVjWGZ71lPMt
/3cV5DOgElcl+QIMK2KCp/vEHX0mpfA0SFx2OK/KRFcG4IaYvpEYXIDV46i9ntTf
GKOqt89QlW8g+V3EvP54eqDmTgw9D/ixOQYrhRKfJBR/hX7R2MhFq0Mh2udMj140
dawMf2QkD02fcgpWtsxtmYrFGvHLeG8RPsYXQSarodBPkQqEAqtpRmiVwUvP+thH
q7FU0d3OP7zf0SV2gpABWybpXIIDms+zjkhTIhUw1MQH1qTOZ9wlF8KYutwbsFdn
0gTWq/3KkXnA05o6Gozun5Z95rXsD7yvJ234Xu50fev+S0AXR0BKxqL2h/dRClDg
iu3adBxCbMQtmuHVN6hG8lvpA5VLsXc5XONlIJwgbKlFaRaS6r44ZULelYP2ofi7
pl2XFePuDAIXRR09mQiZ6SxqSMKSqXENKbOSqIIu7IfZGY4w+w9Zd9lPsAgfyWlS
BhDgEKGEdydsVHVEu3zb3T2N/TyaUHL3mJKe96ePe+vQa14BF3qtWpOvblouma6P
OwCGUhAcX6nYKR1ADAFC5oPAkll7+/V5WF33rXOxEdR2s/pFG86cTIkvrMzscZVW
FZPJmb/ez7ZrtHNHDNLtA74h44MRYw04jlpT0W35IWJ4N+JC3qGDUW0z7jvVWBoI
CCLvgl3vTQisdoFzeo+s1xZ0TOA9YGofEmRfmCAQGCWQT8TDQOsJyUTdqH/2F+KQ
8P0EQaG+1iPV/il6mt8aSU8BR+1XH2jEJzmHcGRvFtqXSBWhp7ucQrhf/g+UBtwv
CpXurAEBTZKdJiAUEdA4KRbfk3GWPDdwwftvdKSIxGehxkWUBuaHvKX6hrPvrXkL
tcPuuGAW5EP/YHr8KBtaiWapmFbT8aP4GyjTQQyV8lUIPQr6PvLaBqhPq4dKHdhh
6/naEAsmhghl2FUifjQdl79OyllVet/PvN7sJUgPfvrx9opcmf3ddma4OtYpHzeO
dSyRIlfOqkR02pSj6g35n/HPulo4MZY7oje13rnKLdNXyMDH79CdQJOMcRBlj0Nc
cRVOtwjCjxaN2fwZfm9/A6TsrzsoUiyDNnFXsHqyZCUoyodkmowEAhDrNqdKp7G8
O45aaxPTBMOOR+PKldfIcmTdj8BAnVNBLPUptSY0E74Llw1gdZvbeYKeJ4jJkSEG
33iVQtsWSGrZFXeJwZHVRiPLNFI2ZxnIMQsK/KZMObLJSWk8h9Udr09lkMP5evsC
L9Z+lsy04yCNpf8kZFjIo2IyiiKZuW5D0xX9KadEbp+ymGF3AeJ8viImghsFJkhd
E8uip3sKRiM+sIMIfZ28w35sUzJ6u+oq/JYY89+sJdftlqN0yk80uZJMGWKUnXO7
U0ru9gSrwpHaBC8uWBDCkJgXisdPgwkeZPA/KylYZY+Tzu7+UQvqxEuct/cs+10q
cOJ/vueTojpVaWOdjsCck+4upCr0I0bYyozWLUSwiRhh+7DeozBjtt7ixbHxj7nX
LYRf2WiO83hqpiNvEf/gWjLHrJfUmTITlEPInOErm8w0Yem8UhEIpUq/83DBkLTw
kM9CRU6KuDEm+MFpNK2rzzGJA29y/u/fnFPaz8H+0F5+7vgnWGzzn0aifx7ovWWb
Wh1mL+rsTU3hySVDa2lrZHs2YS+b4/ZR9K3x6YWWmlGINvvyEHB8Y0Gb/VZ05B/R
lFyiqSODgLWOoeatCSc98sOm5vDnzEsZCqzkW5oRPhyAnroXThawnSUJiFx0UrG1
85kGZINDYQs/h0nAoVR+VlNm83xkss5Kd4ZKoLwNqIZnHAQwEXzy8831D1CEV1Uv
O8ShlDp1eLYold4/1eaARhO9oEnkbWz0PBp5C5F5uB6Yj9YHt0VbsMKa54AaerZb
05XewsVtb2Bafj/feC78W/bYnghUYe9hjfTBMWGgmZsLJSme/OTHwIrzZQKUSISF
2LKvARJHOsFjY6OgLsFGYILws0kzEIelxLlTvnWMIUeA3PLYzYfifpwOrA6vuz/F
jndwkfuPgntS6Ypj7fnsTmtT/JqlqKTWgUlKblB9R0+6zBoYB9LPGF2T3cwZYFvq
csIdw1P2A/+Z7a0e7OA0uHfxyO2cKhBXGk7mVGRONwo3JlQSOXaf0aTdkQNFfM8d
Z7a266LRQ+nQvsmzFqriE7svbp0HDLdA0xTA9ZVojCDPLntoSzxYlslolfYdpMAK
B3wjbAMVb43pYOAtDUgbGROGKVtcelLKrWPdnn1X7fmGodTZAtTIJ08BDk/1Km7c
nk0I1kb4AcGcJrnARB3f7IZm1cbSLEzxQgmjTHtvKMlYnNV3bi25CUP/2CPxu9AX
iK52whVQiNZ2cft4mXBwqCzBCE6bcWr3jxmImnZteH0vi53D2xylVN0zb2yeodbY
Ilmv1wUWToa+4PYw5rIEFsq5ZfM1MsDuIUE2QyaVW89oZwKMHToMdOig6wAQ+Y8h
JiUXy2DjlZbMV9VEw3FShqz7rkskMTpnSL/oKte1KP/0bouOOLW1uePZ7jFPDXej
MoVBIGtqi23ahH0So0X8GXgHnKfZYnGqu2av5FvhT81OMYvNkhKrhix4Rt0WynXk
A89lhJDuWQz+XDX98MFMZJu6FhiiA7aU1dBZdwOGYv8AT088BCF3dtUBu+L2LR1b
BFN6lk7CldyQ/VtT7k7YfUliuH0qLiXG0yZV6Cj/ZX9cIJizO8p/MoDR7ua4EJB9
ztFNUEIWmmnIOr7FSqsqrU2wbbJ+7YP5vx6Z4nlKvb7kPH9v9v1PkWOqDSxj4gJh
nCZDCemeon2CmOCHi/8WVkFtYmE+WEUXbc8lCdM8o5244Z77vXQZ3vlOxEsXRA8C
GlP/nK4flzrXqhDGouqLU3VLYcm8cODAqN0MgXIFkgmaGKWl2LXkc4xEBgHIWEGW
jSZszDMUbVDtbBVX//mz0WSKhdGFa0C7+XZR/mhvxqfsj1X2pbQwSi0UyfZUX7EL
Z1nfwzhPq8tX+oR3TNcF3mrJDx7jyv5BXQfeaXCd+3VtTw1cNm/vbmOrexVwMZrz
lagMCYe4ndVRQzAj9JciCbN1tLQOggbH7A0RFkUMBuMUM8DDcvNtxillFwsKHykR
MGX4OO0qD8jIt1wLPA82ITRAp93muSVEf1wbtS1aFSostMFQWdMBYheaprWr0kYW
M0Yep8sMeLYIX5jw/NBkpfDU8mU8Ypt6nXAss//7rAF0GAHDeCYS7b9k36kHhziX
NN/pLGA9yv+WSyrKP/v+ruEZ7KQpSpeGG0EOl6Qyr/bQ/QmpNFDnmwWNE4yGia/o
LAtsxHK3pa62qRdwUD9RsYPfuV12KDvWLn4/PiCKbTbKZOK5OFhKiMB7naMGqD9H
qPEP0hY6VVwFjjr8oq8rw536VaWzoMAtnqe8JYVTgURFJ4xr9+/tcl8R+7doUZvc
T5dC6ejjHvxQ107thp/+L7lp8Gh3WiDkWwo4q3u4q+lO6uaIcSY57CXAGGz/IR6C
KQoCVBJDT5peekiS+/o3NwERzuXw8HKqUM911C5FLOXFQGffGWWXaZzpkFpj5Ata
smPa4pavEw4+pI+JaUKKEoSejNEP08BNciRTf+cmefBWQH47M/heBMGUjXg/8dSo
5yWrwuSyrwpftBUuOw5Oz2DTYdONGF84ZH1ipQmT/5R2FfnCfYwV2FFVrIBUEDv9
H5iFKHMKDgNkLVUZHB3mDcbxK5wUMarUy2mx0zTVCMER1ml4/3acuwCXJ9jl66L6
5/jwbrSQD6mDez/yezObP8zQ/+16dCNQRIluLbmtikztWCcnyv8ZCM+dn8ySQ3lM
Imf89Zqoj78X2mS0CDucl3AL8L2WOviZV2AJt//cuAVfKWkF6wZOwW45vSAm+ZV6
nOUtMIeSs3jh7Kr8aO1RAanSVll5L2zB6pjb5fKNAc86sMUPGEqmwZemRZ53fhDr
KQt2UOCunhOLkNMuQihi76sVuAC3BbAjrbInLBxuqECSqlkzLCRO6pxofTBFNn4a
3Cf+tffMZ70Z8ZgXu9XniRme8qk6SGS2sMHe0QuJE5PykQ6t+yBszBmWgFBy0Crx
hOFEukmJi4Hs/0+sk6baW+3Vz8GEdhb9NCrBZu5lru9/SZrn5jUXQZDsb6qn4nlm
vLMzt7n5PzPJ5pSgzwToxg/7VgwnVlCql5YBA8hm9jAUOTRC7Ob/SgLmraLOaiRd
LujBsYaJyo6yB+kr97efgrkOSRNuPUkjMftSAkH8w+8+4UKPkSP5qeAwBuoQrxb8
ag+IUmee5y8JxRz0WCNj1Q75d5MMUhhuZC2NnBVsj3qyctCuazkx0Nk6LeH8HaxW
pSeZn2BSdnXoy/9E5MQdNGCXCL3mLkxb1wC+jzZN4zZdwgbRY05vSbt2WhO/6oQF
EQEh4JYQNl9t/GQE1cCCIuG4q3O3d3u7GRHgJ8PEY8gh3qfNrYxWe4BIsZAd6owZ
6utHKAn1hyVKTwy7bdLA9ERrx1dIW2MKQQmMHvmgB1gm9viSHxeVxfkYPD7z223B
hGQXKaO3nWzO2ehZbAW2R2VjN4Ab4txqAofyVyWQ1NAqI9XuqQDwo48t8Kd4w2JM
kBE6DbD0fZ3qYT6UumsR4muK9+2/0QBu3no0CUOxi4QCw88AJ5VBb4svJx0+mb9I
sBXteYRkgR6T5rRUo1Q4F3YIJ8E6y70e31lTpy8ufrLRwPp7paYA3FN9+bhfX2RR
Ki8luUSRUh5y8PwM4jz+kLS4N/ds0eTg6fT7/cohAFE25LuMCEfOOJxoWs6hPtus
BcyTxlCY4LCAqd/GATsWL/qGnBamMjjiOnY8bTCiFMFelxnl2ZxF4k3cEEqWLdtN
KwOQ0NmQlOolzDe1UCNdCVuCpveYE7LtddJ1aMp0bkGGL7zHVhUQDKv0Ualf4XhM
n7/98uGn2rnHTSy9WfH1JYYP/xZa77x7sdQXAdL5bPhF6KK4dGcLUzkV06bv/bkq
YFOk2M6gMp6mKpNLiKqkLXq33+uFbGQ7lXMdUyOoHaG+mwQoawDCukRslFJXV8/B
oUkvFCHvVqEHY9KHLXcrQAh2WTcI8yiJ4xo+DE1J44xC2TK5OZ/Mo1hmRQRk101A
4hytqTfDLcXQ4nbrDcEGVG98oYGCKSxEmvyLHdd3EwAdjj1i0rusHA7GGO3PQ1tC
9vRA+GZaDLzpOI1QgkqlldpwQORDLvqu16gbsgFtnZaiXvVsDyALEm3YO3P+NRdU
1sTBuSb6Fl9iOFZ1HM0WhOAO5m7A13LhDmSgsRCisr+tjsqoB5rQoHbRQ5t4SQoa
v0cEaJTQ4U7mZIyH88n6pKAZKuOoRCKrcX9hYKyqVuEicMq2J48BdKAtsW4Dsl4T
h8DTDa7g7+/3nDYZqKopTadsql563W9O9+ggIWhspsyLIlHM2ABczYvGJc0X9Ghd
B/4OrpucyD4F3XqZ/2f074IRV+RzuYcCsJ3d1QD14lqotLqdtc97TL+EanSufTPD
mN6FIorCpXe/jDkWeUmfzUD2ovmqO8QaZJ+jn1inziC9ja/01JVL//n0ku2JTSPr
NpfrqgsOSp/QDhHm1Pbx50FjdaBq5V7374/xb0q4pjTk0S+U4Lbji5V5r24Tta13
Yxe0QnTQU+Xjoz0gpNcK/qb1J0uYOqxuB5owiXRghfBnTwAiX2Uuq4e0csNEuon1
k+KRha1k3+k+rsH5y11zSNOOWIigw0kqQ7pzNsUvRJg2H7UKbFBbgyFvUYRSLiIz
TcLSeiRZrWe2beq8VYBtzpbtpBcgeWtzPD8zA5/JSbwMVQIb/cew5QAD/eWI6gUq
1BIKlRK/EaS125K6yapdkFqW5ck21M9epnt3YnBD/IVDcJ4dvleRAYi73ZDaeo5x
vlvIp/OuCfVb7DviaYJ4R1MGoz91zM3DdAY7A9Z22vNptbTh3arU6U+4YjEhttzv
IImCbZ8qDnU6c5zuy+pDJ4IQ6EPdcpCytoGT+jW1UditKbl31DVcG0FZ/nMRCmIX
YEnZdGLCEn3C8dz7ynoCxxi1XZ0RMOO8Xan5Oc5Pzc3YhI6qZwt6T9LOrUbzwsX1
jPtdlAPC0zIUqg5PYOl8H4q7auWuZJ/uD9ye+udvlguFdC+54N4JuJU1CaWd/SlV
csfTyXiyJmZd/5z1mAmZHhxgTWr9A0V7zWHL70HcBF2XTz3RtWrjXPmNfOOl54Ks
vpsYTHs7AOLAIAYsiIkj2UzGgY6Nuf92mEMOKGa2XTlU4UA2stsl1Q+XYIXWdm/+
iLmwAug5RlkuHl+35+lP2A/phZ23C/hTsfTHCREc8/bD6bXUPLOulLyS9WoQbfSo
NarLHGalpyCdylTUo60jS2Qr0XTmLW4a+HFc0A3DLIntdIQcPCkk8p6glbvxNp3v
pj9zdwWFj//OY2qEvGWPx7oHp2xa9CILyblQVVtHOKNrrFb25lSKNFhlhMZq2wGC
E7QtPS1pXutRS343MCfsVrRejyVTs41MdMjirse1Ka8HnauDLEWjgeXRyiUGDcpM
1IKc6TOJ3G+mzkOc0lHbIPvxVN6p32UQNJ1fnIRuG+qu2yngR88wu8lhV+4YhNn6
8wbrofgG0JqBMMqeMWO7UVzN1Ot5IaNX0ASv1ukt5smGNQWMGf5MgWKQhFBH4NHX
rXt4l3PPThbYgffBxmZHXVGIkVM0OgKY7u7o5ov2ACoWiDdDXArvd3X454rmZybn
S9St6uxf9KCOtCSh/YX6Z4y4Uv8fXu5UIZ+ZPgERy79AtAyAcVJcbPNFCIpI555x
Mq+UmFQH66wSzxHeuuVmdkIcisajJvFhCI5xVeT5pbEk/SUw9uuA9L9NmWbQaxiR
INQrRFKsAD8ARzaejmGPQUQjSTTk4cChM27uq5zJFlMeDYWG4wKxfa5GNTCN09wA
GFTFc8NHekk+c+AXNVk3ETJ/m1UbgwhV1cFdHuw6B0dZDfXC6GxaIik2VQk9Y/Sm
G1t5CoD1wXtB6RaCygLL7LCfz+FMxGLXwUF4IXokHaFUpZki9fvPg5sGPqjR0BMV
m8kER6DqffrMMxg+f+4uexPvuJhgTgjnzh964X1gUVNT32S+Ci/f2LLWivD3Qt4j
u/jLnfEKFSCRvM/NrTfmgi4xiZWmyVYKsUArNQm6xu5ADpmIBHQUE6R/TEtA+A5v
mFcILlzi5K0+aW18ufcNsBQffK1KpFbakIVDRBgDTWwNvk22L3W5xkOpzQyaVvn/
hDckz8m0pVj0Mji3+3lwrV6DHkogjFkCd6ODhM58Y6g78yXeRB0IKqKJ4IXN0TPM
5xByaO8HsKzXmPcobjgwPR5c6Wdb/fd+mdOmz8YmQI9Nd0tL/RAK1SZsEV+U8yDo
8Y/EOKSJdpdhTXc7epuZZ3vUCNE8iIYk7ks5AZ+fo1d6UWNkma4m8Hnf4fw6b1wb
4aTkhkDPh2+qBZ8ePO71ibw3Z+nYVAdFu6OqFXwMrIIz7LXLc88xfgJ5U2AucY5K
cnIdS38wtjV9u4M2+RU8/8yYY25U43tN+8Asll7zfkFud+doLUWmu2Nfl4MuDRhY
w4fUpoLWdqK3OZAFSBFAbSqsy1TneZ00PV84N4AfWLWqQnNYKhaHZHLdaJ8nFki/
ht5Ma1SkN5CuZGHxoRdLBMV+FHO+/sPLTGv8YGkOylVHd4AAtcCXn2dO/+5ra6mj
ytn8TChyEYvB2+oYRJePrIi0I2J8mEyP/4b0UmObO8DkH6gWda48hkYYHFHsHnjU
yw3hLhYrM3MhhPiITsU3DYFEJgmPUAPIcE460VNb0OqysAac6CcMhoVT4sBDqnRK
OOswCD1wVqUJmfH4uOxHnA5TDtOL1bkubUaSPC7o7UIZaQD+M7LIKgiKuIM//vFa
3tY23i2lreiPdZQIBQq+QGQn8WMM9l9ZL0MSpnWflLJSqdbNUL4Lm8HwUpT1+8vY
KzsNHEEU3W+LT6poeKPQMBoZAk9gqTbQb06UAmUbWvG0OJN1xdQYqe5u2IOVnZbd
NVHF/IlB1l5bfSZ0meWVwvH8pIKHdO7JqO3Lsx4zO2bWFFHX+JHRSSdA8Se8k4LO
i/+G2vw+Obgj1PF60t0NNLTlxkyV7cs5/wqRhPHzxrHO7BTkdX7lIzXzJEOAsOAC
uSufA8dprv6j3RiAAsW+p+3Jb036J38yBkQnkxIGlQxG3brYxqA8Ly85RR406gTA
QAR4k2tpOxRG3vqHe+Mpud4svtzI0pS7+cX1DY3hlnvlvPmTgnv7A3jgpn4qr1Ce
n7PDeYO14M/7y0TKAKzQxzsc2VNb/IIABD0rj6dIjf3blXgnRChiHAmFcQJkCeYD
cOVc2zJSpEN26L6LjS/kkFYakQxWemI6D4P+KcZDmbnH54pmG0YkoNS5HLGo7izs
ucRO//rQqIHfAL90s5JWMNUUpJYnUnu5qcnOJ6k4tfiXmeyx8tbaI8XtrlTvtBfv
uVBZucm0ICX3KcsC3SobZX7dlrerO+hkLEZsKKp9tSroEIQzOXaJqbz+15cdzdFA
hza7Ix08mg+d4TaxpKRDZ2iZ0sGZ3v086OKH+4U9nr8pyu8U37MtpBpC1WJyujcW
qRPgZCJCFiRwBZw/8rOpRTTJrvyGUgVRr/YqEBWvqrbFA2hc75D0gyKAzgOPKNnL
u18USMYKdEzP+/wvlQukQB+CkmVM4cJ/eAsVU4Wfhr5YE+jVXfhN+rmR/4hg9UOz
+3iL13rKrF2VJmt15tZ4FrX4S94LqjCLnuvKWOgaR3YoXRqXLeKvObrn5BAmw8DE
Wla6f4343B2CkzjeSrD2PBJy+Y1b50PDLfEkx/VY+NHUqGXJ9zLqx8dqOBVHjWiq
IfjkX9p+NOjIwBijTyySu9eAHIuQ2btdR/Ph4eYwjIdoF2Ro0dVCC250agGaZ+8p
KHul7HNcakIgMFxxdpNVR9cN7NjcPm4vWebxwhUVFC+ZU6Gur7NjLVJogeS2+dUc
CkUsn3MwkO4Du7CTfVtf1bkpKuM1VHJIqmnTkhdK1j7/KRdKvLF9aP038Q+vFukk
m8uFxVfkQkE53PtWmSKnvRm7HOZ2IuV9o9LCMJ+aIPxAePVt8U7CiygL3v8asF/E
dLWK8B6YiF6KXxqNYfXzZVCj8FjKlJ6RcMi8cVAlRe1eZOd5CXcEDMyxybu/RIJh
3bMFfzN0n/swUKkXjEs1zF9h2kCK/Go/d3FcISyD74rN/qNAr1azgkgDSewXE0AT
DJ2bQBZg4Aw5lXiWWXhHXGx/QBtf2m0nUrx9SnzlaPIkcB8V/HAzk4iHDBdUwzXl
1tJ8Db/GTXXgEV2mBhcF/6rg01FMNcHEAuqfAJlv3XjybEsz4r4GCMj9TNmY/+6Y
/OndZezROdEGDIvonX65o05Pga2V9pBt9TAXn/SWqc60aQp1n0i0GZqDiIgqCF+E
urrGVXrPhO0Q6aQoGwClbm07PT6xRHlKiwXIur5MLo/elWxoAes+NosHRCjZDOvk
WXOFWnJuaWI2YJX5hZCYPiY1G7qn5sQLORoJDRkz+nMbIl509Q0cicP90KxLcJtC
dH5rZsnBJXPt76Qqq4m/ysP37p3bJImp6xyEuLYaCibIxtVf1i2hdx9dg8Zf20Qc
ReYSgSrz9yhRjqJVQC0H96gSGc5tqiQ62Qo4n2l3M3Eeb5EkP8w6Uza7Zti5EXrK
kDwdg5Kwm+wBK7kCD0uxbmJWI/l4u29OflJ+cqE4Oydy0ob8oW1/p3QuZct270rQ
1lJ1rS6RSOH/6lWUJRgAz9v0i1u7yN1wJtEF0pZuaet9fO8jJ6k33oHUtTamAJIv
EkGhPzxlLBZRcCy/PAU/bfuSOv7tMfW7PsajniMOXMrbKXdCHiyijSD6v7Fesvdc
F4NuKYl52bbMDeBOSknJlm+cfjGL+ETFFDt6ZHQwIapbOcPG33XzDIM6EAH5fnvp
900rpQ3/9SM89Ernz6LKCDRXcUT29YQJ0HjPIeqJGCzSYcql/rm+x5ysHOqDf+7m
v/ROurqpIkcYG4F+WdlFySFAIVm5jK2ZHB5Yj6RPnuj3KE9sIHUiRNYjBX+IXd3c
s/Xv5xd6cB4tSeq7ID5riTpMp+F3/304yfUHCLB00ZUqCKWEUuUMtf2XyC+PeR3M
0U5KfutMoKDVzrfi/ze56qnTSOV4+E5bhzPz3oTGPPbI6nPnLQRIrZG1Xb/ER9Xd
D8TxXObta2pTHszTp3aNPio2eSggd0bsIfYZlDksqWx7AwOMBcopID1Ouzc+BM/8
8FEHyHiTk4ncxApCMkcIoZ/pVUQiIPprJQ8HW/1nTbwVr5Ok/xttTpLDQtooqarX
jJBGb/602bJSZxTQSu8Nq+xmQZzmf7zEItcg0gAbfzVRvH3yh6BW0azsE63TzzQS
RRBDLuH3yGlG6Fle3Pggzhh32pZHVVF9TB/CSOvIJlngmrAAqR5OGpCp3s1nvY5L
NYvFRr970HBYtWYciARaTgOQQp2oWyX2nMo3dXs/2ZfApoBa5z0mhkzsPlpolb7q
LA2t4IE6saRQS9uvSBNwE73gQ2Y9F+UXlkVKtusIWywh1dhzaSvpS4m2IT5iQfZH
8TFH7Ivw1QC6BW1Vi01EcDi4Md6NeeNHjJ7xjxuahGFI+5qO6Ie+SIYcaIV7Bjow
s7i31ZfLQ/VqnJuBcE+H+xerllULOIKdlj45kJgbwDoDV0eb8ZpGqdHtEoC0o7DE
3vBI+SAnxxwp0s0sgr338t0thC/6Eo6KMZcvRWYcOm1KLwLWixZfWdATPHr3r2JJ
jcfvzFrk506Nu03wsVvnIc2MR76V1Moc1U4zHAeAGb6fhWeKr6Fv+CeoNSRgKeZ7
77lhbtukSA6UDBNDP1axWPqmSAtvaQIQ8J9YHEJi0Kd3WQGSHNgPyQ9FEDOFwJu5
IpjxLBHCkIlZbYto9z/2NmVie75gj5o1cbQBQvcNE4Lca9lgSXA7cCwkIiqc6NIZ
87EAyF5W/Td35rLU1MZVYB5F6Om4IPTgMOJ1SbanViaKNwaRWP9hgNDEOEmrnv8S
eflOq6igv9MtpStEP0OD7wQicL8CI8euML3kFG/aTtjC6zMcZOq7nxunYtATET8r
k6zqlEVK8RjBdr7JH+LS7W7NT/sYpIA6gwBIvIW+ajtgmp2MuHealB1Yt/QjhqWR
WEhrLXpzVehuLmQpObgMyJXohiC43i17bIs5jYDXqXv6xClPmTGcHiCeMvfWC/Gf
38l7/wP/BTwIKbr6dPjdWc7NkClM1CXwK5PWZap4rpzQfb8ht309TE1NFx0bSnsE
cxc6Ju0JVmYRVFHEb8fnWLbpK/6BIJOgYZiwCpEr/7x9Tu4gRTPVXD4TX71FaG+k
n1w66VDseEkTs4zDgRi8/alz473Xe8gjbWaF/KaiJbZe/+2NVDj7JowbFMrbtsy/
3Ai/PxulXGv6Fp5wYVDuymhAGA1BsHCVDdQKsjBzeH1ezo03uwSJHH9SWxL8JdSL
htb07+WAvLx9Yx2x15lGxKJJ7xZoC+4tKVRBeLsL+3kYbu8T6ojJGiij8AFgTXlB
+tQ8s/Gl2v9IHpTAC1HSRwfng67HgQgyHVKFrX03ohVXZ/P/T0SacSM/UOXdZPL5
bIIzvZQFdun0YPCEh3QVOH6cdLoO4Iwv5FLnO2CT0siE5XUUNNcmcM9Ffftn+CM2
XFpY7lm3MTYuZPMB1x93/VQ0vWcpyVP+qL/enfTpIC61XMnf5/8zjLxKkOINUggH
ZIZ47UhRcyz+JZ9EcrJibCuD05apvkxDd0E5tiwO0CFiBcGUOzla/b8CF8TPQ9+H
nDgj5qme0EVuhW2yOPNP+OMW3YRGTK+AHPVSNbRWEErevtjlojA4/tQA3wTKSlup
Bxb83lMadtR4X9ZKXybOi9uuxLpvSORrJa5K0yWrtf/hor+WAvdHPZZ0ecukxPUp
j+JEuGs2cHgQZvmLaYVDTF2mkj6vd95adgqTRIRW1I5A934NUwNv9CFuCwxUtCl3
2+wvlw/dNR/GJfkamhpiRVBFj1OoCKFJoCQDdIT9Cs0VSNlD8mKYSiGgqObNwlS3
9wiW49iGbrgs9h41ZIZTdgAsJ3y/q/3qu434I4t19+JR2AWQcyj9zTHozrL2bxHT
0hTiIpprXkQMjD3dVfE5uluNIlm1lBMrk6/8QgeO7ct0+uCRYkryTytHZTRnhn9b
Rf7MQLTmZ0RyS8mq5Wu8N10oUWP9SAxEqXR/lNm7uPrp/w0xfK5iN88ipvuus1p1
pwjr3K89yu0l1qZQyCcinkFbXZZro+/l3BU388NyrHiQUnsQT5kg1nO9Q+77S9fR
znrSxeGsQAoeqo7BbqYmYT+Zz5X1MGC1MUTtyWAK9rxpYXSLLzg1sInHo5soyyTa
Z/dIWTJ5nRXc7tQ40sQVJGLOFhET+NBjDTDteWFQm59gZXIlOjybKo6bzVheMNkP
Aq0Rxc5UkstkqssrvgSLcV87EIbH4R0PTv7wR9+OrdE87cFlIeaM7jIVGdMfq24x
tKiLJahrVYiYHvd/fsejgC7rBDDsh8+HYJFixliANvhYZfIxaBbTOvhMUyGVJ59H
SihRbxeyFhjMcelfGl30mLwSDhoqqn2rFOZTFmYbaJNVZvnxZiKzbxVdyL03VQoy
+NDO1Y79I8ZTZf5ljHFJ/hLtu2xvMjzlz2DkospM7mR1JCHCQ9ChGE3Dj8TaHBVM
gHhP1PzN9TvzYNU8/4jrN5CeiRUKpN5Ag3/PHCrU9S0DdSOxF/QbZfXeEA9h/Dw9
xBFzHG3lEZkZqaJepqvU5vAzhHalyxgmQTpkui9kzyF2VkxdN6HcMz0QMvoO/A1/
l4HqmTC7W+zM8djKB4XE/Ai8J+YRPHhaISbercYbN6Qwkr2cjKMyFFxd79WvZvL4
Jje6ku4Q6Fuhb+GarW6NSGZo0AGHJw6rgPg8QOOLXTJG8Fjjs19slhG2EHgjwl/U
42HMrT2Tmh8ZvmUlwS8/up+7VV9Aslk+9IU5BS9uuRlVtC7FMQ8LORbKa2AgK6HV
MH+ZEjfWOfIM/6Yaxi/Dji9GHj7JQ5ubukam88SC9bPwF2KJkHuJKOtIZFQb8FGj
PM3U2snO8xjZ61SeFOauGert1gpybZfcXuSD9bPmusY+D1fqQJr2KMgL7VbNOAkL
qFrdnD2u5WFwyLISPjIu7kScransYPq/dtmkMiCqHOTOVuJC8drW9zwh93/YA7vm
CrZRAATx42ynmkavmdK4nmszMdSfGuuzTCtLonRgWtj+uCkzL73q9FOiCpnNG/BA
h91aFauwMAOv4wVgW1OS0iJ9qStRI4EweKfFx8b9uK3VoxaCMlfvDS+tYrcaOfEC
L8yOQmPzBJj7kKzqVdgr051VRPmDcOdTnmRkyufSnqCEey4i7JWJkgD4gjVt/Vi/
Zwf+covkAGgQymevuMv/Dx+TFBTQiBUclbRvPZBfglCM55TQM/OCKViIA8+ssx5O
kMWM9q9TGMdiFrQyQMMuG90NhzFPMGaMy0T91HklNjAv3oieNtNZ+y5rLDCnWyJq
wHjt+tN8x19oCt3nj66smqjBH2xH2S5DZwSHUhN8KEvG5wxT9NzR2SzY2NXU1Xv1
hp9RGLFBNqHrDF31NxC1z3cwCknlerM9Bq09rQoTd12SxKin+OoXIos7NOrLZI7e
ZtUVYIGSK8t3FbTTNtrw8npQTlk7pjnjHRmQ0e+lyYkxJQrL51ZArqD0fKSe7ElV
0517LR5OgdJkK+JGSY/BMxA/jHHNwUFxQG2KqzjvS5EGQeHSylCnUe3DtQF73oB8
K8/sT9IN3Bb1WnBMcthgpIpfeqiKVNlHC61Fa9DmCXXjbbomAab+MA3WOy1R+fK9
ShiQiYvqhn7v1DKxEV7/O/8xGzQDmPfa2Yb2OT3GImeng2d4cf2etlul4G1AdYb6
bSD8AbW62bDF/leOSxMzYGLKyhfkmnqyiJ4yCATQVdlxCJLaQpnoElSivGlD2gha
KZcBwupqVOWu/nbtCAxlSN+X+QCf19wCzD8vW+7PRXrj0sB3a+EcmSKlEwMfQoAQ
kkpgdojl2hKtpjuDl6+kbVvmcjj/mzvb5FRCFSseavCNAQngDDqobGBMPJwy86sc
YIDQZ7efOLtfEbzh2C3PLml6SzY00x8mg7nzyeaNdw0uVTwOFa25ky1zNktzC4C6
tIm2r3tGprGMf++/u25GUNI3Zfm5Hpugy8WT5rpNEH3+9qGOGMR3f27GQiIPUEYd
YuWTFmnt9njuJrb5jo0W5jmOFVXbKu0sHT/MKqm+i/X1cfpSerLMFayB9SKFN0PJ
fCpawy8Y33DPxZi7KwHKEYhW1rLa4WUaHsoVGSD1E9YDgBn+cix/Fsw449KcbCiv
uYGSASdfwpNk1Tv5fPEDEr8hqocBmhsLAFz8kEsAA5o0QE8A509S1fJcNZmjwrAl
haTULir6WENum0Cg9woT8YkC8il9zdN/8vb6r7Tb2gK1VC8Ci5hVp/ogqfRB5xL5
R1S5S/gFb2HTYENgLfh65Nn+f203R6AWMXzUtGdzt48Iek06dVl/v7jUR2SI/U5X
SrxiRBb2EpBIgJCI3gsFWR/WqbXNp5z9lCgiPVCuDn0gqFyL7NuoJwLMDazI9Std
Mb+dpHSAW9QswPUZQhDDRENOO5jK066lyB0kfVCkej6X5dlQRNUH9odVXsXJzFxo
M0gpTycr4NmaNEHi7gGloESOK2ffHebiSSMFlqR7NankDv5OUsygeC7RoAmc4F1l
80b8D6FFfJCpTJw0fuJ3deQP+cU5Sm5Fw+QEWWB/HeeO1Mx63pSkiJMdCG9C2nNB
iQ77UEUhFPr555eqtsveI9ijQygw7GjS5vARcEnmOAizJ+ml4Jt3oEGMwwcDG+2r
OzCYnSMBN1vo1RufuzF5uhljzCb/qO54NNanLcvAPa2jul+AAdU9kNbS2qSiw1r6
EbILzBlu7VFDf8IF4okSz5+4fST8mJaYEOrbAgE2gAfynBKzfbfCfMiggN6WKCr7
rvG8Uuk7+q5JK0ZqXcNcQ4/8rTKK2AQU3wW2fTBLRbg1ddrDMCrdTlIX9/D3bDG0
DC6n2zA5GGJM4nt43Gn2mHeF+ETgA2HVmmj0RzMuP7dIUQYblUIVqd65EiA10/B8
dpMMyTQxEWmEKcBNjW6pKwy4K4s+UAevMxeLRsaNHQJlXSBxwJttQINBjgozAYRG
S+NJrzdKJ8DYzD1GNIbX+QpG9rg4FXPY+bgUBKlR5HH2ez42B0PYuHL+/ts1/grp
pr3Ni1eKrE7R0GMyinUh9tKXBgnK5oxEkSeD1c8Copr96EwIgterISWRmFhv/bZz
fl0D3j5Jcgfglgo7bQWzw0nzGm78m/c8EMIeNkU9a8uucABr8PrZv/uLfB5UczjA
PfUaPu9qwPcjlOlasjnyZjp/8tWVyWBX8ceK4SmPfxvaT+AYXW1MjH8GvF+2fnyB
/zTC+mXfTDNa22f85lQAacJV+6gGuAGI1c8SkKcizLPxjg5Hogj68h2laEOsJJAt
P6qsuhe6HklyGbUT2gizdOwPVk/0rXaIEfdnd8tUCbaLMOmfkdBQRLfzd4uZ52TG
k58rgfP20+4baxvf7LK7gBzro9o0Dvlb/VjrpbNNLdY1Iq8JFq8HjTrhp+9op71R
G8uWyJ1aAWw8LfWbXqTTTCpT6lZRw2H0Db0H4GLDrs8wxqD8IxC2wkMdZ/xkrB79
7RbeS9k9scMXCMJUho5CSvGDz+1flU0FOabAM9JcVHd/JNCZSAeHNFC0lu6FmAiG
aksFdJ8E/pDhrBJJVcXpeD5Zezf75kg55ryHqMDPtTE5tnAkPkbzTGsn3JPNrNSU
8bJGcL0p7fpB0zJnaEDrmi88i9gnLQQu72/9X3nVNWa4Wt+5j7cgFaiXFZmREOJP
3dEg+l8LbiG2H21b77qNN9pqjqYcwSxBbBggcrM1og0R9wJkl2yEmArmuIV5BN4R
azQJjCsgKhCoubwEt4KrT9LOtG1vwf82JiKInAMXc76qNOHrh5CwDcoPsEoNR4Rw
4KmKxYepmaRJvHiy6VL+zLIVJsY8g/5jgyVwFq01wRwO3zDnZ6fpPpOPjhmT40Jj
Sq9IvJZmNoZB9Ej6W6KocvuuTICQO/jT4FGrMVHKP0wOkmT0/cTBXocjgaGYuNv+
i6EvOOQTKyjr+eqPRAudRXEysIjtuFrl2CuZaEyb3SATg95ZK1Sn6Ek+NhDaR1UC
m2Sn8fi0yMgFbGYIjhXCeQJD2JwL3h2/O4mE7zkC/6T+bDxTmwkLQbYyoZgqgWvo
UN3rBw9L3/Vr4UIEPme5GUGcwP5WkqF9z6RQAgdd3jZdgUf7yFa1jZE/DGlZDRYb
JpE5pjDBUH/SNomVNuhHefFQQbndPPRVWxiYGYvcvl3pqm0LDoJVTvmvRnS2xbaf
8ZQqHVyfEyhuRRnSALZn//lKvBbJN9w/PD4dZeCewuARpAmWmfJAnJ6caBbRZaV3
DzddlL3kqvKH4iWyvluHeFNVP43qkIeuRrdWvhmOd6DtxfZ9ZYV+3g0brD7afvg9
o9X7RBaDtOuJFBG2+NlEunE8O+WxVoSjQqHZLinVebB4gd6L87XmNosvSqNwJKdI
2yYcjt806BhgQz2VxIT5ATiceJRT8b1P3pG0lRc66qtuke1YCYhKid6YfY92616C
w5z7UgTK6r3QtdxSAokOs4kUZbTST9/57A5BFANB8T6JTBaFpwpQqhGTecSMSIUH
OYY16oRCSnpXisDw1nO2PsJHjAoOrp7Sts7U8HA03vM5Dc2q0RSFump46DvqCiIj
kIdQWOm9TtzLgLDablxpBDzp0/4LIKYBMT2r0Hbg3zr1oMy/BuojmG7PrVKstoiM
2WjIDMJw5Chw4kWOybe2suLcEE+4de9ZJZYThVWMCcRHVuT7xX4wDOI3lQ33zwiW
JyTRj6tkTkuU+QXsyiZASfkTKbuHZ0320JBrWlo6Az9+1shecjY7iCoJdvMS8AH9
LZO6DqpO+8ZpKo2FviEBjuEACwO5FZ6ELFlWwLRjrHSWW7rJc/xMfIzXM53Vqy6K
1ZJn/tYv8T2UMMft7/A/sbdMHi1lv3C5D/J9lM41fZNmIzrfmRA2mkyuTLDG+qXN
oAecPxciSaH4y6kdxJZyiYtH504lQGgxvzvDSCqD0Ylf2ETUwByybTfUXMnUxxzT
mpB8eNAF8e5L7eebwAJoW5DKtrQxIGfvcA4JgcC8HPgfWVJ8yU/e8C3uLz6YdlbC
SadO+/2Uq4+rF52JQzVDhxtjb4aYJnMYjHkBZA8olgnlaia12i+TQnzf5DzRrDWi
MOdIAbhFyKrVX7XW0G0TfD1Bmik6ixAvxiC5XnIhqCbMbXtYTnAI51T1tvl32igc
fVgwadHArn6M/dtFNXjVunD/dPWBwFD0GhGYQq0bTTz5oND80mkQw2zw2Kwh3j0R
ZK9LdtlhcsIrl3yhqv7rBiYTZoot02xVM4A9K+Lj+EQ6OjqtymD6Pt+gxs4rDjv1
SX93q4Z0Gpda5R/OXJ7QVDy+5URBkcxBpdh8KEvEXMCKcArsNSpFPG2Z8IkOwBu6
uMSO3JvkZKJvvdkNVOAm8P3O5JAHAv44xOMbf8Ml2sok0lPveWf2jrftKXzjifEJ
5zM/ZrlYa8jBtUrKWdrNF4TFc4HypB4XB7ezpx9DyPTckQi0QYZEg2biWnXUgOd5
yKaSfjualdnWtils3LACmuTguJDXzjGKIq7M6tjQz4ld/gPsiHnmoRGRmtzmsSE2
DfXO6UMn0jOno7ZLqeYn+1lN9EaeQDDOJaQmf1jxLedQ3/0heHMXv3d5tOwTc3YP
AnShsm0iQCpYXzXtEXbFKuJ8OE1BNnGCxZJn58udcoVIdZZ4L5lHbJCHFmze3+Zd
KzNpkZ9UUVaSpvNugf1tVVxj7tHnE2n+ynjl7Jo4p9hYIg4FMu1aNuV/peIaZ8xl
2SgIlyMJQpzB+L2CHUWo1cGRoHcyb5YS39K5FXmtRfwhc4M2EcIEZ8cgHl43mo/y
GyuCXgsQISxEFqTQZwlVF+fCWYqor4HfbzmC9CLP1Ao94yG6cQQxx5x3X3wFyq59
tAmBqRsKmraqwYL8y3Z0x9d2juD95W6ERbt3L6tzPK/FZ9b2dwQLD5lOjpTBmaiH
kHuWwCleWKKjZrqyRO7eg3rrUHS3s5TTpxtuuuMF+D6Dvw1+LbE10xWlcsLEXlgs
8CTNN4GHFqtblfnpCBL0sbRN10Y6T8MGZlqjLjttO6DEr+20fs1CSeZgM1Lhpgb4
iGRCw4R2ACu42h+1KLLdLhPf1bOAn6e8IktkCPVVutaLtCnuXMp/0aLJxmB5n2X3
4JyNXhv7Z/P9V4EndERqBKCwFWXwC/dN4oMglKD4ECUEdXUvok1I2UTJkvI+t/UQ
qOxTb/S865Uzw/aiEr5KOVJMuZIbDFc4R1pmeVxr5OAP5RYljzrIZmEmniVE67ho
u+ZAaBWlmep0EiKbZY3+PlT0fMdeyiePGwQYqgp8dBqkJqC9zCys40jUN5pBGqyW
Rf5or+xuPIgy+QWPbObxOGTJBRCViuYWq5IwnZpbkzAZUTUfp4j9ig2ZucG5jElY
gspqKvfe/0rGMdE7EgCh3N+GYqxDlbnVuEjhJDfEYfOpJMuhotYGxc2duUP7/MQR
X842JVjnilNPz1n4NnO4HVkgft/3k/wYvS5QjUT6ba/8FBD0491xKPVNcyhHjNIO
eJWhG4Wm4xFs3Lvd3qzS4vIkH70QDgpdW/4C+aqqi8+RlZLlkxLWCmyRYmqAM5/s
bGPHnmdw0YHUwdM9tPWi9Xt39OfZIf42tvDqeZI6e3PLKKDB0Cx5e3Na/7+W568f
6zPW8VcHnwl6GPOWU+RTA+WNzvwa9k5S9Z1MQ+HgR4S2XGe1AJlso7DiAgVROKZC
YWia+ve08UAs4XhQ9KY5/IiimzGnnMaXbifMpQTIklk7DF2reZfmF7TUaSxhDpp2
3EakVdZp8OqQ4oVCfBQVRVcSC7Unq/6L+1k2dQyOaCZbAV0dt9OB2jUOXvhwd+fk
SZUSvOqnM+6/o5LSy0BMCWNO0tKLCHuGDdCCVNqQW03jPlKEhXbso8oCEVF/6EnK
rMyZ7JxYXLtwDdltfES+FH0lHJPn4SmRh1ZS9sYL29BoGGNeSh8agOjV/GPOwTtF
fOoDJ9MPJHgnFiMKaZOCr8/YWbaaBh38m4cRiZNu/9tZ1nOtatAsaFJUDRZLY7wt
1FoQWHJQ01ix8iIdaWimHDRqtUwvQxKlbSPLK6T2KVV9yezt+sYTMHVgSjrBtzM/
ko7w26raIRgqn/z1hWdGcYAZhi468rzaSJe/svoPMFsyaVh6ja1NV92sGkbtA6T0
aVgJJwPjiusxjt6ywAZerUy/dyHM9Xpje7KHlL01vi3bp9PFJk8vFRzPZLMGJIAa
h2j0QfDjPy4JPbZwyKVO4HeaIpJVvLUc6S1F9HhH/48bRS3EiEz7lruelDKv64eE
kRdrrL/EOOytmAUCeNhXsfUrGcNd2bH0UJu2UttrkeuZu1OpK4A1f64LAxun8jfg
WEMsZJpdBuk2TKTmihoDkSY8nBi1fIVfaRR/GNkhRzSponWCdrcmxdZQEdfcFePo
BDOGiZzaEZCQMmrpWh10BmS1p2T7S3T9sORtKF75JA9o0gdbhmPCCTMhoOS0j91L
82syE4iDHNHDIrZ4y9+FqPF08RPl6E0NKddJLSzBW7qqVyyMh/YrsMen1F9Ml6cv
R5k6wmd7B3hZ9obFTNCL/CQZiV9H94MFa3i+B9AvAqRYS8Wh5CFR0Yqvzaza68si
4zvScBcpUPIq3EtyM/Yep1yONOBvY3WzPt9KMg+Ie07MgslIILi7JIalcirWxAU3
4DlkWcLaVEntpra4fQtT2+tcYkCgWNpmgjGEDPD7VXgF0CZshZz94UJxhIfidkYz
7mFiYKh9LA4bhSZ7ubbpSGZforipuFNR+7uHjXnfwt6Gq7uqJzR06Pz6f9JDpc0A
0I6j2N7ppjAmO+N5AysK8NvqcYcsCdUjyQShf6bGq+zTVBhEpwYgLD++8aC0pj0t
lptpJK2jjn17tDSKSjoF6wakFizgRB/vJx59eFQ01TloGvZVUpFbytKSBj74k9Gh
lluGVVC4NhhmeD6b+Ndl0EZO9UObmdY9muxoRC3WfXr3efJ07uOb/RYbILMzAeCd
miLEmjTeV3Cqc7QzS6LS9gPEU10SInjcylPQzoiaPu4vU83cRt581hBYz/LF6E5h
fhaU2WbCOOZgiepJtIzWSZjhcwWvr6OFULlku8h9SoKCBpvsHy6wtucfd9MBdwWm
br70kTDkdOHxzhy3CiwuQaQvpsS0oa2FtzKhZ1vhwPjmKgzH2r/GiM4U8M9lwU96
lHUvmtV/dQUjg0/SsBchm9B/DoEhpwrcS37M0Ga+vdbNlwyj4yXLpKKIfarznu9I
339DkO3O/4YBsrwRc+lPnvscqGkaoJfxlR2mMWX2cCnxFip7TzMBxScGRu4aNg7L
bD3FrJ3d6/QhmIBT6aLDoDc+4CcfzBIQenu08Ber6RUxejnGA3bG1CyKMO7ZfdN0
56XXdXeTMibJZNQ22Yb5dqlOTupEN3xruYIyXbVdjgQ+GXNiO2W9fApifLY7Wfdd
Nz4yPKYNR9gYSwfNKrLBMQ4hXW77ZoFgVMHjE4wNYBqDaUrqhIPXc7ouZZiQH/Dd
GVNJ0C+5oJaAno8Q3punJ3C3dhWFd9m1Cpy5VNm3hKkAyB2HTQ7l8IONFle1J0V+
+O7yx/PPYqpDOZKaqPSHpxdJecOXS6ZoliohIzdD5CInxNEQLS+eBivaIjXdjtEC
kVLfLbQJxnakPD2v/qd2J13pGVY0ZzIRh/56u3cPoRHmlp6MG1rL8KNBkqU4wV07
LLp+67F+dSGmY+mgwUXV+p/btMToeufQ+uqDAyFlNNy9mrrUEKz/gsVQn3FJog6G
/hKoc7PzDHAJ5fdEf8Chi3Bl3C1q5cbNjAVf+8CAXNI84m3ZMl5gL7ecO20r0eqn
bWv565sEmyCLjDYGjw9Pj2+AlB+PfTihAI4M4NtBxp4hsrrgQqsjD7o0aVxtxLjU
gVGnm9aXGB8Q7MyXsfyXR7xWIgehqv3HQSbjQa32m5e4vScqATWxYiQHExIRAB4C
8T6P9QOvn47VhY6WlAX2EUaeNCJAYlR+Jm1Q4zrngKdg3pOh1TvEcK5zqFlH61pl
P/LaSUt5Y2hNkPoajOGJW67AuH1IOMuR8cPIr5T6guYnEb+Vl3KUaE8kGYjrqko6
PvOzwWZH7huKifI24akuqjxqRJ/TqY06PbwH2PlVK01QoWQNhcCjTOmxZD8CUfvQ
C9Jl05FRBX+3xK0yZ7DnxSPKfQ1aVP9YWIi9n2EUd2N7cLBtQmIbYv6sRS/yEC80
zFic+4vOtLtjgeI6cxF8797qU1RF1A+lfO4fLXErG2I9zV6YV3FXuLsu8SkpvbbS
a0evuEwU/KwSuu4ybV0dky8c9YpJGbBymOHhkZAGl2Q8X8iUFLuYs4X+Au1od9pI
JQ2zsz9FJUfpDm9Rd8vj1qaQzcW9fhLMdO1dA3OyvoxsDi4l5xUsW8HFpTJ98E9b
Jxw9O6aXr09hlWs1cZrxjb1FsGkXN/by/rHdeIRr6p2Glm6ruZ8qQuv96J1Atmw2
eUFk7zet6M5jhNz519PkK+JtfyRqcBNUADelOQlWpMA7VAhZUOISKUTkQb9K5PXp
7twRALqW0MLfNm8zAc+WdDmKRmk4FpS6wY/bvn8kZOsr1PoiXBybBFU1AY1T+mvf
PpdFO19AucqZ/uhpoXRZBeYN9X1pAqQeUQkbuagyvJRuZPtoka1Fm/KVJZhbCHBd
SwA42Ux6XVmT3/drUSAS5cZjKodn6qQKTakLgRngrl/2Xs4eVqa/Wk6OSGBZBb2B
j9uMFZZ4hoTN3hkhxp9Zo4rUojtRTNi80E0W82TPVtmWYVXCMwe9bcLxpWnDI+/b
WazValuDGJvPYl2tb86KQhOWbmNrrPjg1P7o6GNWT7i4S5Byj9MQHscdcJiz/663
Y8lRnoR0u6Ps2U+Da6ob1X2Sa6hX50wt3V/OyQwG3jHGFAWOCUySTgyLxiz9ukGv
lupDFDzKzZ81HRdB+w8uiOzsNfB8FD4HGRJ/iGhy9BNMlnx1cAfyuCDMlPkSeuL8
rE0TYxRhEwKPhrRgj8RZ2lWKnQFDLFGk4xQHPWuiGlPwtbNgru7vkieZV6A2AxGY
gy/zgDRgLaySlXx0muZ61TZC3vB8pYN3zyB3OTPt3afNpz+mC/SqppQsQeVBJ7b4
ORoZWqj55Njp9R6RY+xJCI6Z3gem0iQCiyuOt/+8WDJAP0sK5Ls9F8P3nnElm4k0
M6fzulQ3sY6cDp9lZVIj7FI0n2UE2Bw/1hOyNhfIhUptWO22XxnrNAXI2P0/RVSA
a9rDiIhWtxTjNTfwFKhcRrBuGkmxB4R5G4B7l88KNh0qyYyApuR5XsFZ8SLfnKCJ
3mTZMHzb4dakIhAPJk5NrqNpKTQZw1zQMsj1SNPQzIitqxJiA6RrJ7hl+g/oDech
sYWINY3QsWkI6JD9ceiRDlB3ypLq2wbn3kAxSsNUukRUEStr+JMTiwd0wiHnXy6d
5HPxZbnujtQ1HSSQUg+bIDQQ4rpYpYgf5nd83PjwmX5LdnK2IRtts8BuDGQba41O
3IIVrO0MVEEvQa2X/tgwgZsmqERMBhB2aKDygwi+/8i/vB8TbpP2/Wecyn2tl2MR
BgExsxFaQ82oxikenOK0nK38BRhhuRl99OtqLGzlgnjUPNG5ishaoR63gLc+oKc0
8VNvQ38O4UwnvC1Fy57CisJjunvzcY9e0jd2oFUOz+LzCX8b4dJt9hmuYR0czQDg
AWI26qgCcAXC2hTX1LKHFQzsFYFjg2FF3TYxPR52yyl0Ix/ElUDbwDUmyhXGzRCk
83y6F2XMCeUPSRC9s6CDesuPd5B4F7bGGaTHmq/6O6hywE/nKB3RMJLc+Rs9+QLW
hm3OMQwh3PUL6wZ8W+9nCsSJhcJn2aBsnL1ZvG+qtARavxH60vdfr13oRJNakxzd
VpjTrJhPWf7iamF45LvCd2xtM6SBgO27bP51cDUiDVp/t65zkJuRJ6D9WWRdmPKW
iQrVr6k9/YWZs4Lhkx4jHINeVpYqRzC0gLKK6edRBg/h7O1Cm2CkuMKDU+XDluMY
Uezmdv/66ha3OBKOoV6XAv5+utzQWtvubsxyPi3MjiFjaJ1EA9xKSkFJF1L/qTPt
nPvA399zGtaaxgwmkoowOZWU54ZdVkhoffRxA3L/cNQEY9wiXEXNOIg7gHj00L/I
EKIKbK8lAHyLrfjl++g4Gw/F6tz0uZXZDvE5ZG2oGMzBgz0iN4N876NkqralT0co
joDuytRu5uO2A9lqAmiI8w3Wg5P8/6QtGVkCIcf46/DSfZeAxXMp3uEzcx0Afr3y
vWGkLawq4D7pXLcuPf1LRiRTu/9zD+w+ZLHtXwyVa0Do4D/BnnumN7HXix4I8ywD
fAoADr5P+RbIRezqXd/biTzjAgJOpDqB1ezOKP7lJUtiF0JVnSip4D7KExX5kpHA
On6Q8lK0ClsyYkL7JbrhJjZzuceoSeTRQHu683l1tlWXVnpGgQEzq+ahl3h1eeGx
T092Dvt3brTdn8k/Qi7iF5flnr7WqozmcGJp+n2phZZSsy3Chro0LNwYyHUHVmiX
LMr8sit4i09asc99KZj1/AIjgfeEj7pRQQNzWNlWM2fWEpMI5gL0fD057i3yYM1V
HeV/UVw55vTGapP9j89pcTBU3xnh2pnPnHbKPedI4zFHYOveEQ0AJwYrRUHNmgUO
NeFjvIq5RmD46c6Cp91U9G8lBK856HbKST/EQGKUHa1/Yg/BZKH6Dnwew8HmabNu
nx0SiBe/Xb2/5UQOiWdLHZA0XRLhVAB5IjNdmNdgYwvPwtTdtbKiPE4Qz1EVK6wZ
bqi3SRDLlxglz8BpNAf/Ce9hmYr4IaVNmAvhPuWRtmXYq/Od2dinw2A8Y3q79S+E
UodGtm6YOFrm3AG4Na/e7U6meiHFB/wrOnvh0cNxIPaUiTRinUvizqYNHvG1qLsl
pen6FBvZ6entE5Il4CJy6x5JIPBrYVym/OZ9d+XQ7qgO0SDeUDQCyWi4xsYbslAY
2omfWCmlIWB5s+RgQ1anZ3vn5QBZq/NPfp5RLCcIjHnBYDx5eWduXUOodkfwX13p
mLG3TRMlAYR0LfZ011cbv4mZYYPkFAJ160eEuV57umw7fkeEu2QHXwNyONtlf0y4
YDjSFvaNGievHCZmPWeS3cYt/iSYA6ZE6DTW1d9KRc0NjIGiMNVzrPXVGQyN5nmW
ggVmTtJP8cJL0IuBzeoTobf5Wd09lYyIVFcGZf/6R0w4EfMJOpOf13hhDgOfNMbl
nO7r5f0n2sxoF1eDgkEOGrYNeHdD1q1qWynqV8uQGBAlMbu82pUo+Vcd4iFLFAEa
UgDlzei05fGf2b6ElnY4Yi4yJKNf3KXcqGSpLy8III2VmRdY+rMhVRQoMfWAuWT9
QtP7mjqpF49T+20FzIeWc41O6jgxXmyCssDfXJyj166RaxnqjiDUyQmjpa5XKwce
sHDMMjkL+TZU4RzWBM+Z3t+yVWcgZVvumAvOpnastVYOw+rCbA2F6oFUOAt4izeJ
mm2jsiY8w38qcE/j94VuzHNYY+3XSqKlxty0pSQREHWqgesrEQClGIx+zFZHBQvt
V27F4W63XIxhrflrE226/On86QahMBIfG3wPsmbpgn2aSKF2GvND2HpmlfSihVlZ
7No5TO+F2bQslF+vaNDD9y6WKHuSxO1X53lRyxRewLT6Z0trLI2i01UjntxMNn+d
/u5aFt9nFv0/H8GuoKlUgSaQTS0awg1VFlec6K34nnPU1GRxCOsvRxmaYAEN9xau
PxAEHyJLp2WG0xoxhZuJp3wdR+7M5iKpD8nw3wrUysTx7E3a4GXHZTYi8qQRE8bL
ZoIKbn87EJvVpPUdxUaWG4fdf+VRSv+k2Y5Yhm3OJfxKbbNVyM61rI8spo7gm+OB
IH0Oout3Af0ewszQM93P8PA3lSLx+igCGB4OXGAGD1lMD/Ivq9Z0ln70TeKOphT1
vZdNtNmqKWBhO/BhR88fmNVAD0udxtT0/vTc79YUlLGmTkX1BZpbJ96Ib7raXWBi
sw/RcLb5+Pqgclk1Ta5fqfkXc8DVQOI53UOtYhgG9UbrTzCciL8ZF6iVdP8Ws8cH
N3QttAvWNDX2NgO+ooDvyto5lDJfcwo/GymbOmqmTIhHyjv6VXfDn2MmF9DQwGvA
SR9NhihAObEu/R3AjONC/Iw8UPWinXdl5ik9sWZZUXf0PIx4y3PbhlO1haIpEQx0
d86qOFkrXPFoJ7+b8pJH+M+VSqxYE9pQztqWyT4dXehPUCrHpM1W5KHoSp2qmAyF
d0wQSzhiIWOkIX0buFFNI1QcD1Obj3mH7FPyEzafgBpWFWHWgn9CjZbhtoZS0nqi
IbBYePPxJZKYkF5VIkkCYX/ELMGcqo6v/TH9pkcisSRH9O+uWxPvjasnEdsmeW8r
jT5IxKWhxkGYZAWc7FEffsh8xcOeyuolngWovFhet+vSuWvrZaf+JjEhBHauZAhU
xzmdwayqkQqZdGdZ/1yKpqrWhsBQ5tL1HC/Q7/I9ErKJ65hqx8W2JwrQSZUeQ7qC
8Z4oQSkeujYZYu7dWQuYqM5N0h+oyQxr0OG1T8S5bG8zjUFIYqjvDYdhnQHUtErr
NYVHkRwuEU/sG/PVrWv8MHjal4mIZUvtd7wlS8I4REzjyL73IYflqHShwo7oi85z
KRA243XNF8RD54H0tIswse4FX8grx0RFmQ29dPBrQrFxMuQYiZTJ0XNmqlvwY+Kt
cO0WSqNHnhts7Gn6VNMD47T6t4O6ntb3n7zGXGOgj5IUgKaIKCQ22sMcbwCpxScT
ZKn/ocJryX5w/grcFNzzly9woRpAIs9upunxJ1ibY1HR5aB/+YkFenh40SrQayMh
eVB4dH/wgLc1QVW0Jf9Z60oIZ8cWkBH73Rda2OEAJCRWRn8ParOGwEdkttiOaGTK
0sTvetPWSR+QHBprrODptg2NjmYXcRoxJl9qqF4uOkHCp7qDc85QuiuJ38Uj9Q4K
3M8pXWPlSuG9VHO2tFr4S/iAk29/mtVTfUysA52Z2RMRgrbNxKaN0JPr8jljpoEn
0lL+cJoFYd7JsZnHNny9zo9fjhDAq7mIJ4PQmfgMrQ0TOlLxS/AKA79+7Ss0mjuz
pYQzS4FzhrQXo7e21vYIrYHGfuriCvmPYXh6RcmMRU/dmVTJA+8lHmsJPDQeT0Ki
9lRkrKoVFtOVNwPT8vqOVGk2nlaPXMh/YyNaDN2LVWcphpjPepvw/IDRplEaMpc/
lN03Bkjxpw+NyNntCHo74VR8nB7R/zN3tliLlVxwrAKeUkMAC0C0Mh53I9Nu9IWd
qStzloGDGfcVq1cTUPh4LRxr5oAeUApk9kj7NBjy8qaVxrIfw87KZ+vP2S8A/vop
XKUl0qLXfnqu/+NL7xSm/W4FqRBjLLvFIg5UDr8uws5SlisbgvBXkf3ybXFx3aHn
Pf3tGVLoljkVNqNIb/z0FRN6HBFEuJmnpwN83rE3MKeIDZxuoPPJZLLeK4MgX49l
AqercLNF7GS75ZAy6Cn83l3PxH4JqIHqqLb1y4HuV6S+kNG/JJxYxsMsGy0Kb04e
aNF4EcHaVUVO0t83U9SXEwT56CHqZVbbUBeAcvuYvJKe1Fo+7RvMbiBMUslwBOVb
N9LkSXuef/x/KvBS4YZUK6TLQz9AG/EEarou55mXTBp+y3xWfF+0cXZocm1CHM9V
QHnm+yLgdBn0Dj47Pyn8/vvPuuLjzXjkuxKkJljJXilR3dLa5IZl8v9hySoEy6tU
dXfd1EFzLUkkqMo0JDyja4eQxuYRY0hv3JDeku9tdF8YNnUDEzioBh1tGP2fRw1h
soHDyrWRSt3ab0bT9nyzzqd5flKwMaewaECqGmeY+wMBzPHNY5Fy/GennT/4lk2d
BRpWC95FKgrEuiub9vYzbtn+4GZoGYKvAa73t6ZYFf1v+Y7XXu5Drquj3dP8d8B6
wTM5/J0Kia/wQ3ozI1DudkVTUam5Mlls4KZPn9s0p6+vSSYeF6Q4zYy0mt0LLtna
1FxQ+qEPN1NergCv4kKdF9tSbUwQgEgBVmPPsIjonaIrma9GfnAAvElmuurXLgj7
1iWwTbi21+fQvfXCRKRQTx4B7wzFaGFP5zNhN/q2JneGWCYaSU71Oieu/aBWq0KI
WitO8sj6LxwV/cVhpu0hBWIDMANwIGo7spOBDsucSsiugwxCt0VYww06cUwF8/DS
jcl241wBM6y7Xfxd6mXif3ZUTMvqeG9/cCLfUHAVYIP+UVeetYVsQ4dnUqPPgDsX
U7KbJ/CNc0OGNbEUzWvFFCevqBwADTovQ6a41tnxk41h0stx4G0pyXXO0yDG0e+H
8vWiFzv0z/Z9r5XdsPs39WWlUuF97elyf/l3b2oXNWlLuqqDc4BKJMt+u++Ai9vN
S7JJPG1PP/ouKY2JQjRB+lDpow28TmhTXuAQLoORaYCGoW+kI5bb7KYxh90+yKmE
DMyjdttPO6iZfM7ih/OrRAEOSqPXQz0YZIG2J1dkgR7Onh2RYMzPac2Tm5PGg9oT
UqIvUZgq/QsspyFTZ0tkN4b56JuBbfUQ2+UdSPo2QvUCZYVEq+2HXNOJo8M4K7mV
pYNERSP65X5VvgMgn3JUS3s7x8cJ0jmPOajlVCAU2UsoShfye1LZtjJolF0phU2Y
cY0vd37oJn39IPN5Ocuend1g6JCuiLzzqsQiiwEcj3m7giqS0Udb4wLPAs1PPtzr
mL8pBU2m+nnzatraPuLaMFNUPOocMzB4WoNRtDUpjtfqg5a6zz4KbN3YkhTs6EUj
o6fteEpda0V2yRT04/kbMxb/W4kT8jgHDm59OxQ4KakBNo2cOGYbnVPTmC4i8ck3
1I4DwQvnHrUHwdjnuPWZd43mGKekvBmE0o5NaRr2DtkVfHGUoFpbTJn1H36eznW7
fdr8KuLqIfHItbEmZn1oG+CL85Lyvnt+U2sBKoJo7kMvP5dGOqighSD/z3CT1+49
0fymJl3Rawkn4o2RjtePsHINX6BXfHhbJEosH4XS4HjLloQWbHRM2J+hvqemURBM
rzp7o35xryT1PzJ74edM+3O9ftcEqgjXRfsnjlNjOCs=
`protect end_protected