`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23616 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
ztM98AhgdU1yftpoSvyhvE7pwbMki4Kc9TpPfPYqGtq662XXhj8Yn9jNCSK4Onal
btl6pgXFaAzn6xIqxWZIKO++JUv3x3/DO9ro/yyMaCxOY92ZgN+UuEIKRTBdkCtC
ek+KInvUTERhlEFzp7rUea7XwqqBN505zZLt06IH5iVWlj9jlteFHBgRqYuvyaXB
t5/p02rAiIK0BEjgdtRWUBP8i4+/6n0Yy1dLkqBqIu9pIIcPaoaM7PKXly9f8ReD
cGxaj1iN/l1wluBp5EJuEd52qDQKDkA3DEvExpqR3Iw2sMGsIbuVYsJJA2CGvhVw
ABpOIzeuNRmSHlx8kQcBiifdBEHkCQjDDtkFIj97Esnay5CGAOR42G6IpYSNJa0t
9kDHU02RwFGVaNNfqCNdf/jvKWDAcAzKUqIiwQWOtADlVTYoFjUGMvbXJgmQxKG5
SsJlxpeYRfV+PNYvkGDdlRRZCuvTFkydzEWGkGB67qjuni998gTswq7JyxKHrK63
ddx8gsKmVwCN0Tqvi08kZXKE5qv/CTxrMz4pDPAzxNnOUQfLDEKIjouhLus9nauF
hgZJkdwQtw1jWlIBnlF/G3RTGYEJ6E5hxQDsA2l70441Gh71jQv1PCDZ1c29dR6k
2ZohpD20NgeZZ4UzZRFNu/aZtwN92LLSKWMmhUXgECpbORc4wbg9a/7k2+0bYhWa
WDwT9bNHQXFvwUi9n/yOyVqjpjCwsDdj4HOaTI3W6TPuyIVEnmhxh7GipsE7PL5U
fl6yclsa30XQAaS7Oy/iaeI8p1AxANH+4b70Cp1k0mv5Pwyeh1rjKYO0YA0COn9o
lmEE3VbB5gbG6dlOUnXgN02XeiZ+u8kst0xr2D9o3apiKmqDYcob0gjzp4XYh3IA
2jQWBvDK3T7HtV/joQPoPihuH4/Ui175J9BeAjC0bAVFEls/2TKcb7jc45ssvq1k
3iqmZrOyH5MQz8o3+Xu4i5POWXMsEez5MfKD1eIfaOdtdo5qpzEsqiOoXjWnOECO
Am2cfa6YsVXl2GveL1+C7bH1Ps8Q+gnGR3cYBy2Os+We/Gfy+joeA1ZcwhVCQwkZ
wp+mRy42eqi3VXhNTu3BtBzIkszDoveQSk3Oku/qbeuHna+SN7IhzGmVQ21qmYYc
VRXBQgbW2wrLmrxaX8nDMXloIey9fQr5NxxVrgtphJ0TWIMBC67wgmb7x1oHbX3+
PESPHxjD4K1J5QjBmSMS7CnE6DW2os4UYMpX/ah0+Teb2XQRzDfWfImvbXu4I8dK
51Vcqu8WYYBtElynyetlfhVWZyQpqsCVMbrGBlHbrNH7nv5zPNDi2w1CjZV9LWAq
jEfN1/MYW+Ara/DcrwBrePqy6UK0wEjv8yL+V9vKCIBRHx4hFPHbokk6fVlyhNdi
LzsnDwxR79IDUL8C1hi21nO4SZQrdwjbjMGYfolbVliR33YAXJpL7ncmuY7+PbZ2
kFCWj8RZ6aG3aXdAURS4KYSsmn1IFskldYtsqXeR2604QLgZIvdFpMInHft2tStj
VX2clLI/AweU3C6suSEl8s8FRx9RvA7oA7ii21vLqdLSzvRQgq4dPFrKVpSJKCzF
+iOfbCXvClDREY2eo14FVPokCw8dVLkgszjIhB68ZvWJp7c1VXdeO8BVVI1kksHh
IISetiPBqV0HuWaHmJh2NeIP9DcPFkr0UNzNyOGLh8kBo0YF6yPsph5URy2BxZQh
B4BlGM3NNfK3Ia4ar57SBDJ+EjtgO5wbNI/f24npphK226HrXxRMgXe+NkknS7wK
ry7NfFc3jEidGs0XW/ooqE234z27sWbAi1Ug5emo51tWz/5qI9F4C+BOeN5TUUZ2
ehpmEAAuxgFpwNdo3CK+McXtI3AmEnIMtaI8cCcRIFuzdgZ2CNk+kprJK+kfqSpL
kqJI/oFD/+XglqPzYtOgS9eyIHa3AEeYN+yYFsINUIQsYty/QwyzPBx0SAsT7aht
+rKv0tZwQoWlhueUCzMsUHUp58Z0I6+GfTWcbBFH4vxMmvNiRex/ugRoHXL1q2Kh
Muzd/o1AqNah6EYdM+hzLa6Iqzg6ptEXULdR1urtFrPeSonulThL3Mn24ulh6La1
S1RSCtTtOchjbOvHo+JKqLWxajHvR707z3I3KNfE4n5mDz8yYUGA+b0tfrMAsSZ4
QBsdJ4apSKlBW1dZohTZh6iQU2fzfDNB6h7kscPkXRFmKWgm5wxPMd6dO3W1Vf7a
4nmZqlhQkidlFG5Vhku/aIZx3EOSfuxzt4iBcfb6y1JQM5FsJTeqRWLdBLRJ4x7b
3Cc8KtbivJrpc3uJJOX97PNhBn0JXIdJ2e5BkTJSPPyrToLPh3GERrQNTk/FdFF7
DPlczh24vrNCJ6JeHnZmPF9iMh0bxXXwVAgSL0PfI9oQiJhM6g8LQxyKP5A9yPUt
tDy8aQu2UGuWRgm1RGEfuLmYHNXxdnjvjedgSS0HM1+EqZqKe5bRNGV2LETRhB7n
e70/vrfFC6AwsXAfzkI2SOzJNVGZFbb0/kdaIiNhI5FkcGJIl3VTUTQ/aTLRYL8a
R+M8DBEBeiOUOMt6qvZ2MPr30/CR+/GS3658THLr/UOh8HJkBkPCH3LamSOF3B3N
I3Y97KXKtcAQ4YY0JLYy/V+8nEpaL11gNqQ6i666IWpfCPvGgcTc5EcU+J8VEizI
2fJN5SSBVV6cxPKfrkrFGDlOdT65gk8W0hJ28SwWap8tZeI9LrbnXea4ljeEvjsb
cX5FOWmld8ZWqZUW0m7qekyUobuHw4UQoZIkKg26Y9+of3z+s35QyOp/vNYUZtgA
O0ZpOIygF/OvQvvw9SD4xf50A0eoECCvNlnfy/dneFOAzTQDkrbdumsFJOC/FVWH
t/7TVtVIqGghQroN+5uuWqU6sLrlPOJApXT6AHjQriH9tOkwr0odVMUlMUhKLPwK
gmVv+gJWUtA1r731Zl4KUB4ETylk9IwAAoXnr3d0gNcwldXheb028AnNzIW5gPf6
ono6yji/mZbJsesycs0i9XPXOZKWIuMfZU8phi7jgQ1FE/9ImMyzlaum9700RV9K
2/dnpZMga4G9ENHeuRt5kaE3Q0aFCkSvNOi5dFqImO7yBostQKtdAdl+QcO/bUxt
SlEYSYY9oFi/5F0+nAp6tQ4g4FxnnsyKEvHiRPTwGOIrl/4WNtR8UFoTLQGOontM
+7lHRcLI0I4AQP+qDbRzrb9AIZQKHbHNgvDgoIHBEyJAi9QgNHDM/0Kil2vv5DtX
JMLpupoDACx1YbdWUmdjY6BwEfi5JzKLt6YTl9nsA5P5Hm0nvGzOHEJIkHqT4OTV
E/Z0CAR/6ozBqyeUUyxBa1CCMjTkVvqQe3yoEobnZw7ltFjutnN3rLFiy/pSt6Qj
SFaZeD6B8+uYdhzJdZ3hpJEbQvvL39WAuxlXvsLz7r5AetXxJiSUxHQu8SuZL66W
9ZIt+W5PWXFszz7grfwkidlYN6fJPE8iS7VViZxi5ZvsH2uZxTaak3lPA1GoVkgt
/uxPlvP/wPhBXsFmQydGzkKi7bkJ7hkkNV2I9uX93PlwH4ZQK2GCGqr+TtTtMqVn
87TCgHZVwBgPE+YSSAk0TEGGype4ePCddNvGV1zdsE9ILB7ObXdj+zsvoLjIocv6
aK6X5xQrzK+E3GNLdzPHty671FiP1ActDx+W4zdGthqEBywh+8ea+5NDG7Abf3yQ
KvL1WFaXWbgEU+glr8YiulFITjyqL7cRJxK1auG6qDt+/R+pvrdOW1YL3/ywYh+v
TJ6jLI4Ax+5ql/Gf8fvsXob/VpHLKd9xjNq7HbP6p1pjcff6ZIks37tusVkNEGn9
Bz0FXh1ul4860mt43dcJlEUeeGR/o+bY87Z1aahGHowyzeK/K35FE2vXorDeZCqd
nNjWcDTCmhWsO5FxQKMQY8Mr16fS+lHJGTwBpd0X/oERfsfHgSyMJlJA6uKGVQBn
xrKhMvXS1s2qqmpGfINe983US72AHzbYrXHPfivEa5LwB8FnQGyYVNvo/KiTeGit
jOxasiYAovRDrymzzg/SOpAkuU2KjKjyGXQSGWhyPNHmYsc70QZyOJa+Smx/Cz/H
BsqEgfc/VbSo3Ayzn4CaGIrU6JGvwIBH2C8u4EZdvpD+fzuUmN4Q+gnH23zj+cFd
ZZatHRTYiC8DQp4R8HiHVy8V2zQOZC0Q8bqXzdJUZEmeccuBL01SF8Ef9iIudCYU
Gcag1CwSmuLItUF5lIPAGOnckiG2B3rPGvhOX3w0Q0iPrP/BJICzd/w/6aMxLXga
Lm4VJiYbzLTChLPLrmdrxYFK8eH4bdCt1uxDSyvEeC8pNkFzWZ2sqwCyXQjL1OY2
FZS8lSDQUeYHz4odkAmvpMOd/CWdXb5b4BiJU6vOQMCS+z1YebCn5bECFSNi+JuB
HTzP5m5YXPd/miDYuUuSUnc7IZ2TYHwSQJ7Cw2TZCnDjpOmdDuP0exiwQ+7ChIS4
kvWEDoLqtSu5e5Cmw3l5euj6278eFR1lBxtk2BDJr893ji32qOw+yt2pAwNtZvDB
eH/xwitWSxkZavYL1ALgHEAjk/0qBq/slsL9uPuC7yaurKoh2eaZSDaNmWkNufnu
gxNjKyYK97udsUY4hMgUWR9GVD3M3PsSmd1KF/LMRG3aiPBQ/utjz4crxdCQXQcK
aLJjM8TXxbA5EJVYTLVtC/aIUZ/a88yv9BNwS+74rj71OzgnhSNgxFDIj3vTfJlx
id9ZNHlqcNLeZmfW5cPjQ84hy0xJYqqlU/EO1w8IyvdNEdUvIPuFIpDtWS1yQxrh
StqbqdfGWqgiuv7uUiD5P5o9gyojQIsNyRgvwlUZB9uGOD/ZNaQQMU4UzXctvC/q
d3/Hu8oz2herHR/Bb6yPcmwl6qsorMQWQ36aV9JmBlrO5+KN4GLwBhzmMPEBWPGe
m3md9UeNVwjOktQGQMdAGANHBoKjaXz3oxYaT5ZwgP/Gq3G9UzF9XwfNhGvuBfh/
t6TIWUPeM0Cn5W3NJPxJj3IAyhSW8tkGLcaNSjDRaFYmI4DIdOOqMaduEbZU+V+z
310JWrqqn2RgqkxGjxZI3jndKAEM9+DC59WvP45vHT5p3wPnPfpT3m4Gzv5LjRGu
sdOFhwEAzO067hb4a2pkGbMGjfJ+hxgT5lqwEW4kjcpwVHF4xQXPQmwRIF6YBu6g
C+3W6NMZyRjC1Onua+fvc3U1+FMkZgQXbJB0Un/fgT3IANjKfzdg65aiHUdS2Nar
844rRxbuLNgY3mY8Q1gMte+w+EdElSX46JXzP0rumgZj+p4vKrs0zfscW4eWu++h
EK0BvpWVhcCr3hqX9mF9Gh2yVfWatEbW8pPXPWiSbzQiQE6t7Fvwpa4W+vbnUoJm
/ZWDqw2iHVaDk+9GrII38PMswyRs2DzFMzhgkijv5jH1WMUjcDu/TLM/BgsPsXmU
la0QLgQztl+2ivhWZPSIcl7AzKbz5BvejOfsCqg5gIrEUbi0LzmGfWiXQyhb+rHY
JJJP4r/EJ3UPLoZ9pkOqHRMiUbQ3MwiMnXNpWUURe7INNPSmaIev9QjqPH3XmqSn
jTbKIZcwmQdpmzvFwJt6yVJ9rMXyygEYTNMZ7AFZFymEILeQSZCeUy8LylLrO2/Z
PtPx3MQoHKWDC5Z/vO8Zje1TKnFHgY/m0PBlhlu5O/l9vCzzCd2t6gH7ABuvR8u8
M1YHZHLZ9hyzVSTnuI2hPbCzI7mYzWmRoyWST7iu74od+cjb1RQwyyqQq2coScyo
a3GrMvs7bvFBRvQLCKI9nWst4lX8udDylQ0MUpW4bAkGrSsZPEUWUR88k/c38WyO
vNmARYcEhdHYz8zzcoipqpVKgHamUAQR1uM+4wxnVlzVQkztD3bHZxmQ+9coHOoh
4AKIFC61BFDzPxknDm9VYc5SKftomeX18npMdFxSI/X9EnzHlQLKWxVyHM23ZI1E
s9TOMOHBo/CkGpNyFQFzriNjDxBhJ0q9c7YpSEEUHOMzjRWwwXf733/zCpsYHsLj
52H0QadRZBi2s+SjURQx8eLQJwsR/VS7nSqrIsnT4nshtL6nE5UCBprYL/fUhdMX
Dx37iaMB6ZfSQ/kenHDjlsMds/xwwDDqTE2kx/pEDppemeDFO7OffgJO3uoEpNyc
NclLN5YZc7EwulrxRixQdULcZ2/6CVdN0u1eSt+0aEYVBwcRe0khb3yqGLqlTjrr
t2+jWtecdw99hbqkXxlDzl7Zj5yRQwR5eortMsHhwToeJ4KXksbECN+wiW0h38Bd
l85nXCrdfOVHlOBhdIr2L32EVbdK/UjurCIw6IE186UJLLD40WoOtTxeiv+N+egq
hYCwxn7kTtiTFT80RpjtfmA8O/g9bDXo602F48t1ggd/kTHD97gN63mxCxJ6i1Gq
XYHk5xY0rU5Be3lekSaVAMDENM/6JXetAvQydSvZK49XEenPPgSQlFbbeD84F58w
P4da0HP8ysvFbGO6QWjafPo1sdiXPhLcq7Qsc7ez9mwSCEon/+b+IMXQzk3gZ9+a
0lEU8Nwbr+/RRnJzaHAiG8+7O7zdWCsSsEGR5xv2HHfurcmBeh/YZB1UspqHutxz
X0jQbFkZ9UMxwcIBbTEWFIeRBBa2s9L8WKUZB6jWqB4fb7JmH1Wav16mwS3Q3ADa
OFvkbAZd7qHRKZ/BwTtbGs0y9EwOgm+taAIJgRcYyaYMRdLNYcP1aSxvQdlJtuyq
2d75YhjXFIC3rAca49VVJCI4UmfjtOItwl+VF5L5nbKDNTpMz1A7GJBKIve6Y4g+
xZlLnlqM1mzjKaTy0LAAg79zSkEZzdIpTBjhSdSRPN6vsTBae2qGoVIqlmVRvEsc
C779kfCT70NAiLlZjj7SK69ipNvGTyMmTNBH5JwtHtaAGfN1pwo6svKW6o5oIOeF
GgYjWwGgOSI9+KEmRwywAks6tQjCYEb8aXSCUDbccmGjnpNQuoR0YKD6sVMxjD0p
3ezPyP6h51OpWErhks1eaJ23Y7ODok5iO9wY3Mrxoni3yw19RjD/pXh6F1kkeuDp
CCulmikVVXFY7Se1HLA3YI67s/O0V9QE7QJXDRDNrrUQpLmu0m4PbzNsyZHU3T49
X3yiRvzh25ArtyOXocKqUF4BzuCRse7Z1OEw3xzsAgCcAUZHRggpFQ4zIoH6myjF
Iwt1WDtRotxKQSMTJ3PU6laz6Qkvz0tv0ydu9QXq0hXlxSQeeEHmyHii4fVZH8e9
RxogiOyn8lW7a/AZ802p/MXYWNgKdIpJ0/qb6kGvgfAOT8Rrbx4YSW1suqxBJXTM
f6mgbyImHpq3A9OiNPSP9GEj9pg8OZoQgPJ+PbO7YjF07xYM4b2W1unG2ch92zKu
OX7Wwa8v2SIzWYiodE+atfzB+h6asUo7dbP2IIX1GYfr56YChzG+tviIriEjI2IX
cPSXxmghFrjt96b+KkIFZhqOVRyxm8O2B4N8xo3PQ5hOq8CAH4Uwx3ReBkTyfIyA
mQsZEyrMWns/W8hXbbZVnJBo+DamwN6sOzUJRrikZrPITJd8+B8L8g8qhkAl0r/J
OMuXBK+HzmeTMfimfzFsjGAu0Syi9rM6eA04pk0ISL150NgOxgXZ9KYcEevnRj6S
neqFTvXSrMpB9vhfPR8jxd7yMekhErMeAcZWg+wgoq1XY87jrn9RMEdNZD136nEt
62SkgDrDetGX7xfWFaXS5UdVUngXzu3A27P4W9PlNCzmHiI/yYKK2z9tndJ2ScLd
Z2fsB7mf3w/zERIu4Hc2Xr3uv8CUhLBP/YTrwxVeJN8WlAWcSq/ZVEH3sVPP926a
VdRhmFEQnwfZuXzvUzm01zExMLdPc2R4d5zT5YaqUWtlfhgaspIdtevtkHuJFFs9
GmW42WozZ6NhhQwC6uo5oB0n6L5Kvg1B3yev0vKN/XgexQHsJEZzqtW+FILpHYbv
4lKunUzw/q6m5iq9BWdDEb48xwk3eDrkQGJTuNnAslAM5QmxcIvhLzCuCwe/CqyI
pk69CW6FJ1F73d6zA/pFUSwx+vqqF4KfhoQi0kUDImrTWr98O1M70PrZktlBCEGk
Z2JIfGX6rduJte1rIuSCCybKnqhiQsCZj2gVA2S8QLqHqk2dbHHNtwmZ6l9RPjAK
7HjdpOvgjo1N0jaUWVZ98llrBRzefyyWgUbfNPZSoM29jJeYBzzjBCEWcaV1jQBL
YLRwmbBcS+84Metc66kdYTu8C1Hr1Vqican4uwvDFZs73IRRmRaDjY+9oZzGpqYi
ywhOM9801V7VWDlnYNRNZljKBf20PedTGHeG3L4NvcQuX3z/UojYwlCaoNu6QVrg
WJ3Kel6YoEABVXH6LdEEHn60nKiOwtqwQGZOytSnKOOlOxn7vOSgYFMnesyVuvka
hCbiml3MSWCpcc04AWFMqsBemei2YMHFsGvS3W+gW5L3Zlz58xFbohWW7PBo+BAz
yCK8qgKJRCpRzO4HBOFR+A676dua8Wiggr+DQV78O8q+C9wMDuY/6K1Z0rVLojgf
/jPoFIAIUTth7gSvwZVIfL25DGtQqFfgoPl0Bv3fOk7mov99StJobmWEteqZsT7h
B5/VNniwcEVpEmixUYxjUh309y3BDZ6UItYwNOO6nr+1V7Ucff5HfSw7XXZXekhD
Eyo8FSq6GuOruHwKvRVuajIqSS6pWcwqIg9UB6IzFYIGFffjzXLwoSVDEWj+qUiQ
4+pCxeVsuRnRU7OHSv37aqW2r1O6Yn6CoDgOd/vnKYoa+5M0QekUDGHFyMAWAzju
qQNyKJ1qdw+R+Z36pfBel+L7HX1WsQwueu9UFppiqHBcRGy5ZUERcDEDeUWcNE4x
ncm489f/Oylx4ZKRiEQKH6qu7VT41VnTHQoZ7Mq4TyOduzpjSllWxYQNPXn9sSZ0
FNSmnE8wt8P7Wc9bYi6rgxF1xG8AS9iK+eZqfF27FezOqzTDJ/qZt1KoY7Yc0JPE
WS/RoGmASp5sVzlh4i8nWffjP1PEjqgeiT6DlFBeQIMe6JxzOudQ4iqKeZgKY4Iy
DtvrBNv9XlNTs8yIi/lCVbZm2I7Z+kxgbUQLKq3qonU2ivxC2wOn/Kxt/83ZwX01
I4/rsv1nXID/qfKS1ZrHSBZSG7BgXbUrElhZAAFNJ7eSwJWRyOckVBOhuVUocSbS
5TQU6SV6vMQiYvyOHuGo1qOr/Jb2U3OaNP1I7WiCoTRE0sg1Oqo05zXk7tg1ozK/
vgzBfyJOpiI2FIkPVF2wGZj1clUJR0hi9E0aaS04+U+2eK+HyFxIQXuatOa2x+I8
Ia87EEjxIPqs6+HMPrG6WQ979RNrx+w1EeY25IPW7awO09rPxQNFX+01HZR196no
hc/9TO8pzW+g1w2Fvo43tqQ9D3LKOvB8fZO4l+L8Ah+2Ji0K+bFaAvsGttBRh5Dh
VQoZyXzK1E4pCD+0LUxj9M8gVSVhNZbxwl3O29GJMKr6xX5Y8VSYPp9Od+7D4YZl
te49lfgVtoDHdtbYY7r1w5PL9n0shpE5bygO+f9dGGNy1jqRlThAUD7CJM9ycbPW
aA5UCm/ENRHvY30KfxQh3075PSrIHM//tU6J4W42P2cmptAwzHJWq+HWRqJvbeFA
Jvt2rI/8T9QqowkjZp+xRpvZQpq6M+6ve3Ujjfb4b2eBbEh2bBEVP05TrfFFJctV
TaavD3VIVWbnsPfbpH7i7aStMCfK+TdEWjytNIgrJHGebefnrcRJM8td8eOrUmfO
+Zy0mLetTe7EgVI+Wg6TmQJTjkIBIXmw4SYdXk9WC17zYzR75BMtnFA6ueKtFM99
YwGdnDBVDpjK2cCO15dZkODAIaMM691lRvzpsBl1wYew+SIkZnPBhaSCew0Nt/cd
Y1bfHPWATTwGgpwAaynsLGkbdebQXh+pYMgldfsunRwXsvRN7vKJsUwES4GLNWUf
oSKUVpjUus7aibxS9LvPVX2+xJMsohLEGeKXRmZRdXCohkEUcDjOON+57zeBlFv9
nvQqTEvFTxlebnvo8UbscxTYPkMvHB+gLmN0xl8VzpcHmYgoM/5Aiilon+ag6PrB
2O8V+ogaK7Xi34WN9hDCl1uKzpeik3FhAvWPxj/1TpINseb7a/i1W/4YV1zyIcXS
0peZCrGq3YnoOsosruddTHp3thPl3Ai1SuP/JScpJ2aeUwxE6AoBZU+JZbo9wWla
j2bjAauuCg0ySw2WIRSnMmQGHXt0ycGYhhtp9X9vE9Vo2CK0wXzpeuwuCBePnV7a
r5xjeEAUsgrx7eQbFNQFPDO4t04bEhbGRflSFsISS1UMjy9YBe05UgVu26Un/auT
AYMgpVZ9nUWNj3M/i7N5Fgvyh6evk+WJ7QGJMVa694btvoDa/gZm7tt0jv4HCYpc
N/YXqU3WS09x/kWy+MCaVGNdU0+DplwMENLK3F8WGZ0AbtFPfKhPL7J/BsYmXWxi
5cvJ7gz//+OYhkfUYq+q88vviE2DE060xV6w7AqDu/o8Drh7RUlxhZ4+rYxE3Uwz
YaRgwIrapVHWwxZ2J2q6y+gHce/2/j4RXzlY+99MfM+FEct7UJbHw7PE9814pONC
VbSmN3ddzvFN3ORyqH/7pUsU1T1Z4T8OmdtfvCeiu7CqLWIPIORrWtbGBqnOEbDe
8OxJCxtvND8G1uUjAHserDUpsbqBK5t3N2Gylroeu033/YlQUvWHDrQeqkwujsbp
henHnZyxk773g/Nlw3CcBJd2vr+bbpyqwwJWDve/0exvowS3PzhaSTbQWx2DJLs9
EE7GlQ3zHlUxs/uQm1R2Mvg4dWBUagAGgdOlaDGQrDhGmQX2Gsm5b9nIDCNxnI8d
1WNPnjrgNBtJvm3J5Hce91R2b9xI1GPBvP2Sv275+nNQvT43iXyaxY9bXLCGtJBK
OfPJ9Ri0mH7uA+O5o7cc5Qcji0RYzfC9ig2vgqZWZPpfvSL9MI8Ry0ccUk9IZsNx
515OMnDZizVR9MpQtNUpo6AaL7KhBJBnYk3hlLjAg93bKM64STtk9sn/t7OgnJJY
SLmFQbWvKbhCUhKVHxUvhkI+sjGHfDAklAKeHv2LzgTdXbWR21ScdXVCnF9mtn5P
CXBaGueVwHPyDPSGVUQX+D4BPqoa43qkCkGr/lbu1HQNaXodAk0StYPps9nuzBLn
m0fCWkKw3mfBK6Bb9sFBXGmeiG8dFQgUMesLqaGbPaPBmi6J910eg9iprL70zDt6
K3ofRduJxTmV2hNoxjZAEpMQmTTfUPKTW5T6JWsdUAuu4QKKh8z3qi6nNB6zljCx
AAXkOjxZeP4ziqmDkueAJFNxWUKue/u9VO7tzhNr2b6olbYcUrMdLakhnEzqd8fr
DnORy9KQbgFEou0yDzBztNopdycSF/sgy7ww7gRXIvQazNKy5boErShmSHEllKjb
1jWbn0WVMrBWCRHf6DoOTqG4pnb9eH/6vp4uUw109yvqvQ0jTJfBDFyhHBSiifAF
2I8MwnPCoJZ0tmjmH1jC84zMWK2+kd6hxyJNvzCaTlrfFP2q7uzXk3WtrAFrLbM/
jgnKY/4zkmV1PJ+B7K3k2O6r+drQyEYkeiV5fzUp2P7DdABRq7q7b/gja6YId8nc
H4yC4SI6iUGkfFcircL9HEgIbjR+BFzSWicAGwqL+MRRIfuCxigvef/V+0y1MS1m
piqbjMWM7RrRVKZxegbQIw5LkMDXVSz2SJd0vdJL+lyer55chW6E5Oz4ayWiczpT
SC4Sq9OINVVunv7aBSQKzZ23ZFCyNdgwVp0ZT09mPd2Hc5PqlqX61YHUN6MQ2DxS
Rz7CuiLsjtCnUjUTy/yOsJ3A7LSv3nXKBQ1tNv/5zBvD+qNOdEMK3z2flRockkKW
2+D0KT/xbwANLIx4gr+MCAve63qP5bfm2NQjLsPj13ytOwgbT/ma/aunuHksr9Ht
pB5ljoSX05UnwHdefQ9BPgbgQSTzPj2/F2LVre6YYVoAA50yFUSAMZZ/M5S9Bidc
qMbF7XysQIJoUnU/RumjFNNk7oOIuC/EGVy8xmMg1yNogIGjn52s/Dvl1vuPS1Y5
WbERBwq4Hm99yKEaCArOvOjqN6h+XnDEOZSlup9AjlhbJfPJAzzkvJl5gphGGXqN
SGajmmKrjQDVtjhQfkVSBXGBD+7+cvUyRQfImh0aZbuBK5F78xtvME/jGFDhyf/U
HVtaxs4Rh4OyoL6pGRA8cDSMuxJQsNBlKGnP+rt0/XzqtAxuUAEWT46myxq4xq+S
bOYYGUnIv7buhepC1ykizvi05aJEDmP2S1AwOX3o7vFyI6J9ff6xIpN+Tq7Zdd1Q
s22UuQqpci9LZIPVLCX+K8k425RajAustAMdkILo5iY6ffvtp2pgJuDMbW4zUj5b
4n7E0wqF53Sug5BwTagwQOiMfrQSCXY52hWxziUo9lzv5Y6PGgo3/iNmRoOIri1f
jfyxVJP0sUKMn5IJ7W0ovJwYnVR/nv/0gewyc4fvtbilkLT76vYYuQd5aRHNzTxU
4yBH55/Y4kkj3vzdpoKG7wY97eWtbQLYhh4RpkR7PcrsgIqsaZ5WIZED5HFhHgb/
69gv+Lx55FOUJvZusvtfH2mN1m4nyr/l8ATp9bOHn0hv/JdRpM9ZzOao2EQHxJ3d
dxIA0mDZqzd3Y97p/wwZP89o0DT3RpdyhwW9xXLfpoH6rNcNMDTc+ePbnJPvIpHW
DX+DdZPtlk83C4xIzmjlou6l25hhzs8h8njW6Eqdl4PWktXDUiG4xZM9zRnir9Bn
sJ3UCntNV8qyKK29mRt2dxz/uZMXFDYBbtS96jKwosPYE3QMNhjISBfsDZEWa/cx
sBFf1BBLdnxhvVa5x9kfFH3TBwPQ4RgksOTJL/dw/KX49eXpUKie9skc4Y87fQi1
LSRd74KZvJNh72+IkggNnZdHkyeVwHOD7VXfL/gl8nUA6lW0F68o1uQXA8JWbEXh
Rtp/g5G2NM8eY4raqlkJ/m0U5MeQP6NsNEW3wRhvsg4ioYTGOTZam+ATqZNNpgzI
upHukjT8MkERTFrDDYg2lpJjBCQj/ARlLJ1166SWbDdN3IyL/lD8jy1ohQA6OgWV
Z0wQo3KuAZ3+ILXj1LVRJAR9fE2O0tjEnxXIFT/Atu5NfdRHS/wxy0NeN+vsm6GP
SSXxEk3KhF9qAW/mbC9PuEnkc+fKf7/ECW8msKVN2rC7RAMuH6WEn5zc+5OIta0X
pHD0jfwLJ9ddhI3t359ly+x5C+WLs5y5j+Yfw6K++1hZ+Zn58/NNPFP5kqip2//7
oPsuDLhbIDFAqxKaulysFzcukFVNdr4HYSQeI38s6//7aqtx9sZ8cbBYJnORoISL
HCJhfp4xWZUTrK/1FNlyYRdaiKO3A2hxhBsXPa6ofcw3LGSjB0ywdeggZyNNOKmH
aNuuM3u0ouNOwkM9sLEUHvJEhthuJc4S0hK5I5DvCdVjsTvm9nvR08Gr+xolzZJ+
0C8jaab1Jw9zjHqbnwQX3mNH8HwVxwYwyUjOyIE65yV4HRVqVUSa+1Cw7kbaSRAq
zVikohr+fEC2dqngp+t2ZyhCpDRiCKTngJkWQY1JetFoI44NVWrknK+h48qDTC4X
vz8LdKKg3zTOrxgDeuf04fyeGIMQcULSMrSPE5TROyVV8fdgrQbhSUupGYvUnR7K
LXjQLdmDozyWShK2/cZkw4arrqDM0h3tvAp2pvjgRVtOPuBsoZ2IdKDpkiGJY3xo
khd586wEW4cYkcUgDrgOopV66QLJ1tIHLFWrTTJTnt6ejsv37OKKX6FS2qaODAWy
2zEIHrKBA8ass6Ru/wID67R0fAi0l/AXk6A494qsD44rLg/RedE0yn8eI17orR7b
J2gpdtA6EyCX2UvnGTCd1OdQUx2/xWKSKPECNwe3qzPKfAFJBHOb4Szk8hVKVQ47
hmLBK0ypbnHt67gSKuu0nnJLB1ChEXdu5IQcPmmZ/3GWlPxYe7xbJtuxTIeGmtPW
2qB58KEOdzyX4CvYdKcVkMPEqY4o7MOlAcqEDOVod9Z8urmy4Sc4MdewL0QJldp5
9e+zhKBz1FBJvDeW5MVZqQPMKrEbtYTtKWi4B0G2Zwe3WI866M7dTqlg2cr9Xyc8
N5AoRFxyb/IngOyC6zg6B0P+OxRZCbYoO+L2H1zzL0gyGOfptZYy7HgBtKjDwChy
iH8XTF+6de3xFUPV7xBq06IsZBDlY4OTUike7v7KjHecPx5gljq01XHRntHBiEMc
a/LEQVdedzshrtTqkGRBZZvw5ndICzQ061PdcpM/xFTp4nI95SCYbJucI05yKTMP
ABAMEH+oHbDx5dWbL4FBjB6ypcOZg745PvVZW/BNTOKcvWxLYgu9tciMFVkpHX5w
7h2olpo8VQU4WkVyD5t5ldH+UTh/CRsfjQRmXp2Cr6WX774HX+Adncj+BWAOYaj+
VrCemiYkwAyaqTVRE35mCLRSsLefApIwmbK3kFmli3j/PnmtFfrfQgdsiR6ffRAA
9yS0PPWp+675V+XlvElAtHi7pgdFvqKMS9sF1/Agv7rYDUzDYJwZu/k722RjHiQ9
wp5A5NHQDTDRAg27WCT0SKGqJYVS5FEjGNP/7pTypoiOq1ola+U2opfC3yiTN1mJ
BOUy4MSvoZEYhXdRt1N1jF28Kq8XojoRcN0BQaJ+3nthonIQQGl4iY0KSy5ZaMCI
lPws6dCpSHIrtBrEQ+Hh4zlzKnkB9xNqCRTko78ICvu+6m6pwvv4wMJySs+CtCzX
TGd6hVa0ebSYeDYOnQ6BFCpScoWy2jUkwSAV1EmHlCYjD9RtMi7zW7cspaWgCvjS
+g0jqUJ9LzO2qWgKGhPYXXbSbrSZe+vEDg4LYCR7THSVe+J0Ny2/gLzqiWFkzV4Q
2DWYWYI3R/R6as8TUhFqq55asKKHV4rjWEVXwoz9PnuIb19Nh36YVPxm8prLs+ZP
PSxCZKShWxLO7TO36StNgf9qXomddwlp665hvh+YKizx2tsl5tcuekCmzDQ7T5OF
aM14uR3R2xj04FRSn3jC0WX9EK+0JXrMD6+sfHhGeIdt2DtCptqZK1JT2Gdq3rxx
2RvQOXpCib8CFwFxbdFiwBsE++b+HH2/ViWH+2jBHw6641Y2uJsvoXHL1vqlQKkZ
qdClnMnaJary4A5LFX1xRxXdsCabaZ3NJrfGE3BWvcHJOuOKHD4aEAfZvZrKPsUG
+LX5WE0B73CmiiEa48qjmK9HFUXvmys+7lDBVp4n546hxNSLVuM1IHehEwYuGM/4
PNtljBtU3wOUE97I1Psh9dKUTYSDpiZ+guyZyOJoJCHuyAz5ng4USthKjHhG6ige
8rwQosK6Mxf5OlshKMFMQj/j474kqjdnb6JnqNe0DCpcr8YaM4T/5mDu/V8mlUJs
766HcTHqU4tVtYdhlQg6jBEuA70qcZdDEMqArnECQf/8cIKL6Wrx+VrCR12aNHsN
2eReJK68xvZcVTZ8hoqlF8oKB6ndFgtqtbZX2BSwjBczkKry8u1WxPoCjXNoypTo
0QIOjQatrRiH11Yb1yjiHU5r8vozET7nW3Oq+2pnRPA8gKKUizdToXM9aQHf9bGb
qu+6P8s+PHcvkzDjQ3sY0Ttc6r2uTEMZFQD9WdAyhrxVX2alwhM/eivmIZSEFESk
yDwuz8egJD30FJ+MpsNUCliINbEDFkbpCIL++mUFEdAzcqaazWx5z5ejHYvANUus
8C66SxSd3nk52Kq8ZbEX2PLcxbAN2sn8aMKjP2wTL2cjv/kxwFpcCC5545lsiMn2
XF1gxXj3T0DnOUsFdRlXN5tQYFzBUpeK2IR+y8TYdqtrVaJNDxMKvXXVfTHVIM2Y
GHvy+ufFOs8k2cwLGepBz0qIZT1qGh+EUBAlTHh5tThjBF2BsQ44g2SBuTydCzlZ
laXDk5MTmEInbZ8ASdnepqA0cmqMeecOkSAvW0TKhi0i/fX56Ih2YV1DDXFSUJCc
/amSttUiSOh9hPPddUdatRHJcc//UmpT016bAXNv6hsametyVg9ChUWWQ+ny5RzE
3qpyx4U8SiCdfS5dc+PHM/7a8vMUeIdPhWXneMko8vmgU8unmLwRM/8uV6CUJFuD
dP66hCYdqe/G/+iy1kXzEBliU9FKxe2Mm/ZlyzGJOokIuRewXGttuyGqfnxmB1zh
xIh+s8FDj1mP+IEVo3iCCwYDom70BTNBoGtL5cRW+ynIfZrPidKZ0agLVuFKLaMf
cm6pLBUdIF/X3UrEOEUN8DdI3Y34Pct+DiEgNkRZNfzNVFuW8hFM4MQNiEbQgr2y
KJfGW7X1U0/3sUhG9p7eQessassbRMKfxQ20z9ASvu2HcUA2CMmUH+amQ6NdL4e8
hYF+Bpnc0FqP4F3OAOc+JuERdSi9Gr2iDogPwAlDICanK++aL2Jj/i2Pg7DwrbBH
D5CRKcoXrw6Lf8rz7o2M85Z6VlL6r1a8gTyCLvcmEsTMC8EEhJU9KFlU7sKdwXR+
1BfKLs+oVho83Wli0Gtm7/j1ovbKA3Hk2iYOcwNg1XhfC4+bGeWjahZjlXEck3+d
3hYAg6poE4uf0vdlhA34CfPaJTPhnjcPoPBj1UAxciOhsRQvyMZ0v/LjCat/jexl
Ppc9Wp8vr0klrVnWizNlor9asMmCJH4AATp2to+sn4Z71HKFwwBdxQCYq4iAssqR
rCuzCy4N1WxpsH6SSXxGay2BKwzVv08tUzMrv5Zo2sCre7VaqZsniVnxgurszTGW
56neYFH0zS5kQCwQJsox3uTzATtJuOz7AHkyNwN/ikunEftyixe5rbwkF0ZuuIin
6QJqCWP3TcGjI0++ahNcAGV37x9iagHZPfaqy83XBawv5bUBGISigQCm+q8J4eTu
/BVABlg31oWV4VHf+XqEtRy7ktU/LWEzjjb2+GUL64bem7KvBeVzYLnb71X8+nof
2VkK4GDJuapSefZ3o1ZaXj55iDUTqSTANCSJC8Z96eZpi+6+mPpcOjzDWN1ypFiL
/qv7kl61O+zhnvWY0tYEEpPA9Do+WyQ7YRTsjhBcp5aL7HlJvFpkc3xazZ5OzzJ8
yzrfbY/FHexnKgAuMNiM8RoDh5KOv2RNll/hgAywonmh7nyOaGB7yVe6aqHrj8E9
iW5lEdsIjBGk7IUIzwLOnDEG1emqiYDM1xzweVLGfdYhe7rWHbNPcVEkkZY58MHD
mwc05gVZTXCkkwMw+sjTjlrklws2HhR8g+ytMonQnXEoEInYsNbbXJXYz2Xf4fjz
ziyTmQUKBn2eQAnaBiNOBN4aUCN5aoiwvjIx1nwEgxlI2eLdYUGZavwtsLD1uXlk
ymez+mlNuNAOvunmEsJcY+83MzMiKYGZ30I4tgRdB+qsPZmTbXdRkQV4gKgKyZCF
YgSPph0AuQKEls1XyxHMMKyCZSpS9I1HaT2p0dlaVyM/ygRDInQyKNY1XHo4wiBE
XkiaH5kEOYOnwuIOTIvr2vtpTG/HPrG1IU/fekOdzghZXxnDn29NC1L7+zYL4PYm
oGBHV7brDVqHSpymzNE5VCXSGa1+D5RagviCmt1jhlx+yw8sMTyevKOqTQDmQ8sM
XtMHPSwGdO8oFOGQFjNhUVsiWvSsD42ehroXtoUvTOcDvbh68C/EQz1Pl092ADxK
z7UWtrPTLNyXE69nWGE6du7HSoswEmj6vJ8kR3DUg1Jo4JfQQWnkOxNHKxVkt9QI
/l6hVhZXMjgNySwCmNpR2dBPN4rEqdsBFziV6ogvX1pF2pjYedWlPTR7qGxmxjIL
DIoUm/ME44S2P10IjpWzHRPOtQzFWgxTqKP3sw+9+Zuqeyoy1x2wFab0MIwdIciT
YpVYHIRPpMWgGEhEi9VEVPqMWg7+xnHUeXolNdEW/bM4P9hAOylY6AKUmtZk0KIG
UezWwP3M6uFfcQ0nPEUCaMeROYMK9b2g6tQG76SaS5NyUjANyfG3OtynGQaTeBUJ
uRH+007oY5b76UfdpCdfGgw9L7Xo7XjJY350x4bQ6Wa39f8kEE/XfFfbU/AwZ/ic
N/AGu9cv37mrfFbtxL3zB8Vbg+Ruqt90rWEbfDUw0wqRePYb8NyzQUYjJFy2kXqx
WSPM8NK9e6qrPhGNEUTGEiFe4IKKzr+LztlN1vq3XyLwgXMSNo50dV87bmBGqPTU
1WItX24tYkKhYw6FmF8zfnk6l9IEKshglWC8ZAaidrhvEQVivRzPh9m5TEjoUS3h
QfyM5nXXhAWhf9p76VRQ0lE2G4bItIxhLf6EG5696eFBwlMYipeC8B7WNQild+T1
l6+Jx4fvvAtb+ZK2WUm3OWhFcPfJToG1IfThplmE+wGfJHctb2eu6D/ubnfO9Opl
v+cley8efnPGeNpVC/01UYBHSH+TeuwWdwX9DvVW15NQVjABwphOdk8YUY3YF5t8
558+eS1ZcG/xcYr5rRmUvQxo5g3y5p9llVrNZmHUVjNz++45n/lIVKSbKDdf6qei
fGR5I80FogtZPG1kzNSbDAx9HgvfDbsDzuGbkn+BDXmzc1w3ifcXzE2GDc+QXlYT
/ueBbH9cWfFTcHsYqOY1pfbLaB9EWR8kNcQj9ZEXzJvOCumUyTZHG8GWJ9Zpj0Z4
nnmF7H8KTwkPlZOVY1btGOs/AzX9tkEzXDnROt4pygLWxiFpAtJjRM3eZt9EDVVB
mS2CQd3VO5wym2msxDC9nMoeIeLe76qU0U6JKlI96OgMHhAg1SICWQwTfu60vM3O
C3Y0ed9DC0vu8d/G5fpBxOW9thLnkcHQZmiCnk64iabSqPW/nGqhz0V4HwDrjb00
OEBhNeCYwxU60peNB5INWypWA/IODwJnFsSYW+k8QBCpumzZ7ggT99nqJAFjeSf7
PrNZeV81VVnxnfHuIjW1fVx32GJQr/FPexEX7RVUtYo3uomuOH0aHNKw7DQU05C7
KJXhCn1hScK+yCctJP14dyhyNZmYRIY2VzHp3+aZ/EJrEgPvCWrBlTnfGgZkfEvf
YYNmBnHOd62t2iOgAEgJ3Yx9ZPSnrJHEJOa//AZFdV6kymsHHIu0tYIZyGZOn5w1
mVwSGsjEYt1JxvOUcgxqRwOnf3IIbXLLEhSeMwPKUvRDklwBXM4I22MqiWWSNggf
em6h1CjOllxUij1Fy4SwaGnBOw+mQCr36Vsf3oN4tSogEaN4k6aIlRynDrS2wM9l
23U6zILizmtry2z1mmZM1bgC8DqMhjCSdaHulAglRNsDO19n4pC6X/TWBVuolzv4
S3pWir1nhl+jTvdnrJd4q1mEW9K/zn26K0AaiCiX1e81euPU9NrKabDzVJau/jEC
gdRiuFiKrHyUM4iGoK6VM/HDrb7UsXCfJI8Xnk8Rpnybml4WwNZiFd6JNKBOvo01
khF44uw9xLggpBdTnU0L7BvmJ15VtYFL9sTAe8vJyw2MlAX+ODYTAWj8AAlg4UtI
o5J562+peFZvRX3+FK4f98LmvYhmHKn52KqhxoJQjdhtxSwKFvhKXGwUzSCqZuux
z8zNy/QHr5Y4ANLaNgtOiV8HqdNuWabTUEyM+hNX2/gYsktZ8WIrqHMD7cMBsEtY
VGfMLwOHJyY102qjDaryUJjtivuJurSZ5iEVitm3IAbc4ifnlxIQH3Q8ZhB06WRc
yjKno/uyuGxR3IkuULc6+DJrnYEQS4FZMjMAvK1MtZlc6dumQ3yfk1qB+Nvyqj8+
nWwwk/gPQWUurm3eKSkIk0F88ekskLULtZz6Baxd31eV6y/rbmML99polN1VucLu
moHlLPweSbAmpe3sPRILKvDRExIA6WsqPZvNNoq8+fyu83Hn9BgZIaqTecmjdKXP
TXCpVLj2htaNW8OzraVqCv6Hh2lL4g6U6TVE0IGcAeWjm7Snliz6uv1wlagZ1lwv
nYFXpDwIXSial+EQXm/xVySyhq6NknYl7pBCSpvYF00POE+p8OhGN3A0jfUvR+RE
vnKExteR6yyoKNOZE6OvMVQLxF4CpWJ6C84LI8RDA6HqAUWMSzhkjtHMa34QMhbC
gdEql1hHs4w8sa7ysMZ9Ph1FahcVQgObi5QPjgJhj2zQ3cKoOKb8hRJRf4W76IVJ
gMMc0r/q8qmpwESkTrvX8vlH9JEokWJqK4JdWpDPHm46bqPLlVEKSjKKX66kU8PK
Eu7JtFdgL2t4PXk1roU5Sl6I5c4ifIhGFsFegSnQLsBW/egDPKErf7dygvgtZzmM
6YvtqGid+lIQOO3ggGzwoBY9zYz8kNvFmnxoq2OEv090be1SjKdoJMIBIbLEi9i8
4fWqJXtddaSbcVWdOeDTx7abMiJwNe7H1kxeowtx6VkAjFNbUo5O0Gy8yYIvnqKB
hXbua5ZGNySvUrTpT79602/RVO/advEcFkkylHb6FJWJkSbG+z/RjPrbJzlDuliq
sLAjTcd7u/4tfspw5HYoLOL1pNh5eUql1KcZajjY+SvTInfWf9nt7IHYZV/9A8Vg
2vS26I0KsbEFA7Jvo8Iy6OeTYOl3Gee0/0Mps0QqlRDU1Eh6WvFqzUP2Jxs5lUOO
iNNmC6MCby31A6HNHsM5e2IoDf105PNy+79TN2V0qfKEmaFkklH1eaapeW0sDf9f
xJNctGdTcLf7TNC/6CbXwXsXgnOCyR4HckuYF0GdJS0Cd+NfQCcmN1Y/yGHKeQD0
rdq8GmW8GL/ZL71aj/N38XZQ/+z3dGvXnADr6WRBzI6hZVRxMrV/ar9awHvSXsKv
ZAJEGolaS41FqfkbUABbX3xHkVgWyM5xQGbayLDLCmI3SP1yeef2WXfdNPk6Fu8D
YmpOMSFgT0bIWB9o2+B3dinpsE3IUdioHhe6/U1Ngxb8Rx6mZbwmdL09nT/fSpmr
vRo0jwuIdZBYQUCx6054+i4i5iGbv4LRFhXs9FWR2PsxqxJ0gpWEec6K1wAjrv8A
WpEvB4rX8GxJeKBYqW87ckdd2Dnz1jkZmJTEy6bux3B758n9qlu9fMj2ym8HlJY3
gqOSS0SGFTzACCTpCOHJ95YWBYQnhbklpyUQ2YeLU2d3TpN0OEwOpu4dRgugYeS2
YnHEYRg/nLuh7t8xS2RNR4tmRM+kWcqxRP0FZD+hHsEQ0wTDZTmRDFbWf879GdMn
AobGjTbiAb055rC07SLxc/PXzikhRxW8KdWQYXdVhDlgGGMlDrhixfxe8DU27gHB
rOyfQ+AEJdW3+NcLJZN7GOwRvrDrFo5aL/+KKe5+tlLDV3RQ+bP/jsDQl1a5o6Px
sifVPb3YAz6XuP6KxidWNCOcmTx50XdyU9h6JHO8OtZBbcMoKXkh71zun/uvISL7
f6cZt8GdPMLGGEtQ+NfFcyQgJ9saXRnJrux2TMsx/rLbrte2DyDuCN3oJbTEmo9E
SKl58OJsfoUFDowZrGSEyr3HcyqyBO6Q5qrL2+cbTNJHtZVd32xRI8ng/CtDx14A
VCHjTFW4Vf4bLrJQTtFU0Qi/SePNnHMR6Gz57STuy+2FP9ZCvVwpgC2+/mo3/qUC
xQB+/cjIo2bIM8O0FVvgVD94meTwhjAYO3W+3GlZUir/xhFAL8HoiyHCoKEdYHM9
iJ4QJTqhCbwUm+e6NcRU7l5+GqU/30tjTYmFD9hw4OKOHrUZH0YbmhV5sSCfLC4X
2jkMJL6b4PIjjUx2GP5wcqMZUdNmBu3WNAY8/eNPSzXPr0YneBfDkPsuCNBKoN18
SwuhJTE1vv+PGr6jKf4PJrllwObAhrpyGxSBG2qUW6GB5fgMTLqfGhuS8BIXSNcl
EH3p30AmWmBeKtnvdJVKqYPthKnvRUBOfijmi9y5wU26NcX6utAoXkZtsJeEqAjn
1JNR4n6na3txIwMm0th64EmjcTDUQgLnUJfQeRXkgZUnibT0Ria6fD2tH7LXg+ju
DBINcybldxsBt4I1ASW0viAX8kPG5xK7tdmi9BhsFXLk9e/45wGAmU9q8v0n8vdC
y/9ky9yzsDCWqSy11GnXSKi1COqk3s/xUpZokKcOJm341DgVKP1SIQfvdTjA+e7N
gUkYqeSncWv/m57/pn+H7N4702whhGP+4xTkutokhAOOYL+xHb7UjIyX4pDQEMFX
nfctMZOnkbk09DZaVFLxOo4GB4moKQViv571LFssu551ZZY/W4KFbmB+WSd0MzfP
cAhjIw0STdkoPL129ofQ+zsOjUKhnvd/wDgOtTKqAbJHCsqfodvLKeQg+e+ep7ei
vbqoxrN6B6Xr1qdocea9Wcq5IbqU3LFNj+sYgM8NQjnfpSEqtyrp2hQGlAjfw04s
pfPCUdd3hZEJ1gzc/2k8g4eTHBm0fQg5y4OyXj7i0BmTFvgHbvs8PaqLWiP7WAYp
dYUwPRAJCCvZCdJQsuX4etxP79QLu4FTeeqFrAIMX3OwHwNOasAHkkG7OQFXcRDU
kFZjGeVYXLEyxHodw2nJMz6DZNKTGn1+ocXPRcQ5LUMHNUa/T3YiTaPuub2cu6k5
3PGh8NledZaEH7lmq2lR8aZ/pu4Zqdu7LOdT+gNL8XW2OdHXmFhUJR+sA4FKY8fX
5LcTt1ibwQlGUDIJKm2EfDxqhzMJFrxJ2sX73qnEYw0lgXA+jhmq87C3NGANXr1S
cSzvf/HkIwV4EbRBJc6It8CdXUbJ3j1+J4RMI+QYh3PkZhBoRGb2m+nI4RGlbFwW
HPSKz1Iwo/Hpc2Lq0pyXcwlUC2gEJEa+tvCYrQ3KdS8GjqFbj55dsDTNRu+MGrWz
kE1d8aKPYUsb+9T5x+W2f1tUjumURpH84FGM4U7L550yblKcS8H9LzI99Ym5Eb3j
LjRmANRl/MzdVCc2YBpOf2xVtty2Oc1pdlRNTdPWAssEtsHVPENlW57s9Qs6F3Q6
IeMNRNLOT58yO3+Z7Tl8lG7XKW0ydrKulVo11etFvU+hUJcjV6FcF2keXhVrGIz4
9Z5p0hdEec33JATxAG7Og6lWIpx9Tfu6vpU/6CuILx+eowW+mYd9yxM3P7pXH8sq
r30VczImR3uFzTys1IfgCKNc4YZPQX4RE/KCLWrwhLP/UCFgsHExN0eZbYQ21abW
9DMkg+ZPA27n9RzBMbMx74ZfXDKZv1RQvk+1sRTI2/SgCylqthIV3vJdoyt9VMgI
CCLX3Vug2UcpcbuG4LViji0bAf6tI46l+f9vPMS2UXJqmZcz0NjSfVx991Ad//El
Sog7TtFJ8gLFOuBKyOkS4xYPKJUxQQ+UfD9AvfSIaHyjlKPw4q35ehyiXg5P8QgM
UJoA6OIOAdUwAm+91NxN9ClM1wDRCBGfyGhxmoQ81/fIso7zE5bpT91D0CXW4jsA
q4ngmwGfrh+M81rLWweLg8df3VsBAY63893W/yxj6HG5Gzn1+qfl4RCGfkc5xRc6
Y31T+es/tpNXSOULIcHfLY45U7YFlQj+XGrpgxfTQ8iZYbDSj1HZMFQb9aue4F8B
/j70Ml+oq9/0I9GHYDKS+KeBV6xLFdOoIRoeWmZ1Zgz7VEDG/Km/TBkY8oNrRUyJ
LdePLFUQt/zxRcLEpmga02R03q+lSEhgNmf5Llx9v+gToneQVwxxfFGGQv5LKk8Y
GPQjq9rW5qc/sx9zj0OoULh3d+5aEdNK6ZL3ooJyUuxFvUg0xArRUAly5VnY8cFM
i0qbDsjVsV63drW2WccbF7JGk/5YkcUNEKof9hiyg2qwG0AuCvhnqjnN6TAI58AO
ShwM8i5JgT2MoXjN5eNat0+KmDyVAZgcdaVS0HKcPmp0/gPyhOKXsVK5ovoclI0B
6MfWugxKEIc7/SNj+xFKZ71+PD2e1aedUbwt7SUwe/thDnYO9YZuy5u6RARqaJbY
80LnzD67uPqEeIgsPmasD0RjM/ZjzK/eOhbTd/QohF+PEsTPUATHZNfLmpa1qgTg
I0qK2piYYcOVQK2KtY4+ZQUNG1BzsgAtABigNa3OUfGfzmtVhzJshcWHfOXIo870
ZzJfQEtC8BYEbFvidhLBlgSQXW/Yny0wwcAj4MTxqm19cTprQRT6/w1Bies5kA+Q
N6JcEiCfh841E0oQJT5Z+gI/UmzK8WO8X2MDIlvzMqNX25MG66hsI5eR/Lmy+bmj
qDmO27m0xNw3V4nfEhSYMXdm8/C1gl4GAFXHwsjRyU/xRlyr/n856pn6OlPfDV9G
HAPUim/52rkk+/onrTrdDKWF8ED1zG8fHJ1V5zgQSdoM9iAm2sHqxkG+T7Vamn4o
hwCL7BlMaj6NQy2ZW0VB3rxFVUw6XpOszlCSMOMp3q0dbz7L7oPv/Bor55ycrwcg
CH0YfFyaKnxTYP01JetO6vOiDZGrrrT6htaKZx9BBYn0DSYv5puNEq7DUpS5aLbZ
nyrTlLaxWijolFJrOiEDmTRHjguPYuZTezfnPA4Ys/m+KwoDfVeUxMOidtld9aSX
bhlH0tVS2LebRlmi0j8B1fnZIk8q84WwFGn0i0kXPjq//xCN9+/+SuZN9LqGhq7t
Ijsxrl+d61xNv0KJgVPi4NIa4K/mMnl2DsrBLTFQOGl+NZl+YUm+o7V4FWRc+8C9
f9xY1PJQNB8PzMn97EuEx5V516T5kKf9TKzc2KlWh0x7aWQKpZ578DAffSPJ+uBH
FBOBDN8lvrDppEM9BVArix+mqY1DoZOVCQs0MgBjrqKJhGd0RAi4M9pBv1VnyTyC
Z/bnRe0WI8Ov0DtJDnF+lL8a3l4fddlU87aJjZQzLscXGXbxRDxfDVI0YFdOHY8y
BQ3r37bW9J5qkhsLP7zCUvGZCQ6Q2HobLmjrxNAEXpgl2QZCsomhDQ6aGG4BQJ5H
XfL7nhmCDriEMMRdC0nv3+/Mo0/61XK3e/mNuZm+o39TumERZf8l0LYuYPbin2S7
gWExRPbSDiStppHmMSw8Ah9sKbKKhYDiT9V3YFonwa9MEBUhdJmn7dA/JBF9mlla
Bf97Eo4i5rFnddobvfBYjSY8a7Wap+lZ+Itbk/D7CkiGaEBmyDwbd1LKOenNEwkh
jS4CY+OgHqM9IYIOHYgyDfpk8uU4MUrM59RI9UV+SaMFILy7tWz74uMNZCbfvVhn
CNvlQT62jrXlHRu1TZ8N6r2TAvAPYyW4gBMFbbLqdsjNTdQpOFI6uBRAR1EAaRpQ
6aHewJJZWGRHz6sRs+89IpV1XCyR40EX7JhlZVmKHXuZGClJMXUJ9HgVJkqL3m/8
8NbHklN0BRv0OnzP+ttO/4gwKsQtdDxLjd5DcdCqf42Ybr/+xOeJYsrgUkiD6wd9
vfBYxck2/r7bKMHFbE6zUe7bQQSdNjbFnUymSkatF84cJmb6SienhwbAaEOVla8I
Rt9Fdlo6yEhBO7+k1Q/i4zXbTv8n/WWCYwAQWnmkhnyvgL8ds5hL7eAv5jNMTAzD
PTTs2taaPzgWDMflwZ/4BN0MOkA8urm/b5Bzip8tpjakKBOJCZcPJd1WMDHVMS61
iRni2Edcoj3VrAbUi6nC4EPJ8jffi71k1KgwB+hMvSD50z01z+b/Q0QxRLdNPLTL
CvRkIqO//2QjfwLILEtOmZBiyqcui0U/df6VzL1Uxi/ZNPExZd4JXuax06k2Kyot
Ulu3aigEq6A08UkIIrcd0G8d32KKUu80JFlfWwE5aBb6+bipsJEW3eEO19KMUAln
AjFsEHHaPQsGtdlEid1g7Gdd7/ywmiMcNnkz6MthFWVP8/ZeVY0ebRsYm6RTSYBp
nGg+unsrPbtmy65Yr4LfOx7cOBO0kIXAZt79brJ/ZksoFjWjfTL3Tunmo1AsCekA
pMVUE4bMQga7oQ8q8N6VsLhqESeZvkgF9gaDKQsxtl8DGNajiaSEFCeRWutd+eER
NE77cw4Z1qC4/ZfjgWRZXXOWHjqMjoLP4dDJVzJmNoAJKXy7tGbsJ53BOanUkytV
iVxCLpQUQNPBuGvzf7IguKVN3rqeoZKsHmm9lKHhxDtX72dUW+T+cvqcXpHXTGkR
BKvB/nInTWPSFDElJ6DmY5G19KHC9Q//OBUnp06fhnm+he3ISbq1c5QJuPvaMvpm
xt9Y88JTIm8TJyqm0Z2jWTNrndYkdfJFUcvcOJIJIFXX+FnxoYCrdSbtAZMlEimp
XC4JzO+pMuhnbDGqM5zCpmu5tuqgPd7nZiNaii16JTJO29hzJEXzqMiR9wAU+IBY
ys7vLox2ghq3eeVnZZOUSVAZhdeHI1Y1KkDc5UTvcPWc75lX49+MZg9EEa/riIAn
OJ3rx06ueX5xGfrj7v/3Rh7U64Sahv4u04WQYdyEwFBtt7QEKEIdWGqRQ/5N3Yw0
bOXAsMU47HIxsNsonmgqNJ18NHiDe2h2bN/SotQjViEYG7ztZzXTRmwsj0VZ7bz/
OIvA1HAN68Fv7rBoOlWxQ6CFBXpGG3qYubqNN4l+OPlbf+glsvWV7FtQvoyZYVmG
4S1V4IZeqK6/kAhZYurGrkelljAmWmv8ZO7hIz0nCZwJJ/83It5ZTDaS7iaWz0O8
tNP3XnoSaQTDfsbeit4dpEYTLPEk4IfmArXUEAH/fPfB/Q7Kpe2CRNJ1ATR1sbUn
FqXnnymWZBY0y0X2vIk4UUOLyIabANl8Ec/ntX/uXZh/cLNCsnzOIUncFlmcOFJS
YapI2xEMZTGPQDmQsEuJrSXy2A1lIn0517zRM37JkQ+Uk/ivviNTiD1RRL5dOEiO
RrWcsB9jRFHfLoFdpvsTYbRbFQArOwmjPcg75wMUvabRo4Kg1W/4O7A7Ogw75N4a
rQlqesSV25VDrc5w4rSrYP1bzgeWNrZOoglFRysJY4Acfx+XDSj9KPkQo1PajNns
HL74btB5WqwNuerXuN6w5o5ZJDAysIhymTtr8PJ9/i+PpntI0gjkuyNIgt46dolu
GS4S64MkduMIX8hURhvcHP5EfvHVEdVqZSddGuWNG7ujrlUCfrzxFldv6DSu3lzS
7oFd7g0/6VybjY7iIJ1DWUUnDTslIcL7ICGEGkTMUvsPvJ64hr0QJPnPca1CRDeS
k1+LT1H3zLz2RKRX0n4DtkMQ442hy91NfyHLwmgRnsL06UC5vOYrhCYJpxacp6li
jdEL//SIQSVySsX8R0K1lXJ3tsn5YBgpk7o8ovVVyt20UAXhkExxpUwic/oRwBey
KiBit8GfeaUWID4622Y9SZJ4XBPz3jHk4i+eRMJL5Ssqh6wt1lLlIPWXKZlIuGVl
BUrrQCcoSvmy4IdRk9Hi6XfOBYt2hsGpIMwm899I6kbfILcVnyvi6kxQ6jGHHkS7
DdeME7Be9pbLCP1P8T/Bq/jb0glkALGubZmWEsqi8TkNzUd4y6VM6Uiq6TMPjTHb
qbAaO1egHLtQQjCW/tue2dj69T+LBcWeceRuJi1Da3Cbsywk7Pys3MkWfIQX8MRO
iVpuk6/vs3kEAXjb0QWO15XMyquvs4jdUpp9O/idBaXnIKj4iphmMo8Dc08IzoDE
XZ904RBDB167hglgcreiEAL6tQlKLFCRIeIrPqxAtJfqtqhSDTznn8t1u3MIBvmU
Wtl0nSN5WV2p6F1XwCrRU5bZSqP5QuTmxSVVFOWI3AECvWeHhNrCFXttCiFgv/bB
5gVG08qZHuQFsPNp28XpqNYK6JEuQSqW6Qj7yvM42tItFfXycp8KCnYpunkYUfdx
B67ANu6xEvdBpLBWdN+7CIg94MvPW2o2fQm0yf6DcgZW/kXTmVMcGL2ap463PIep
YfDH9Merk2JehDfhRL6tYYUxjFWJ6A2BwuxqkvvNkzCRyuqIGeaJDArQUz5utJlz
zY0gIqgkqR/FTSoWqO2orqmlUxby4o6ZqeNf6XXmh+zbuTb5t/bZnDuHTZ3klCOf
+Ebc555ldDWvH30/LAhJ0189LJ7RknRzstDnnahh02rLWRSi/jPGzav7HzirrWB9
E4Pe+aoYwAWyUV6FA4kbNju2s0c4hLqPIBMYKA3bKLalDibUHJwSOBa1H7g/NfIU
b1at+Ong4XcS3nD0rpAmMCXmkakp5kCxSnxlgmtSE0VlWCC2opAMHic7DtuXEByc
tFwwNLLrjg+21+pZTXMqkxVVWFQI8NrX4Ms2W1sS0XfnQNUAcw24LyU/baEf+wyd
hRmgDslCic9kz6gTEouhX+6Yr5/U+HdKvsfdKSpHF9Jsj/S60a9214rxbsxPt7hS
/eI7pZC+XxaNUwoLakP6wp4IHuC0mLgOK7vOGq14Gds8g3b+wNvvICLdSgMw69ol
R8BgkYGi+lCfMpRp8pO6q8by2dBUQtSB/56qPGUrQ05o8JbNLs9w3KpRcAZTg0Br
DfsoOVbqa3eqTjN/t08pb2lOdQfPcQqxInkX/bxlrRhSQYgYSAcHt3Vu9OQBkqx+
dpjtTHkJev3KNVewbMDiuin1v9jUeZTVjcoI/IkYFzCDGBD4GMmsf14kKNe5NZ9h
2V9gK2IB1r3ymfL3p0QiCPUiqKtDHpE1u3FCk1VmtVl8EdTjhfcE1bVTEFKIkkpc
J+OYNTIyKKBI/GrlbI7m/VX7oITRVjyxbCBhJkELAihkakmy3KFe6cO452I6BYbf
SNte4n7LgL4QoppcqTCoj/v34mlWZy3bfA9Ha7UHb4c046EFGcbuihCkAitWwMgZ
HRSbiqXH9e8zr0jlJEsnOc/GpKF5eGM0wj7VJLjLLLEXTG/0ELcg239p43INOtYn
GGOuKRu6HrsY+dRL009pG2YDEFoV+BsHHoM6y9U04KL3srOSapl4zYd+k6uaz+jA
fXI+BbSPaoguY+E70PXaLfjr/qLIeaWfcXNluBFG0BL5dYr8CxLwUByOTPAmuonj
0muWj+nFwNKhz3rSLRz+krXlXLJr3XneqYcKA6xYQis3GX9Zblsl6QSMJ2XTWnXY
oi90D5ybWAmuBV1l3Ub4pbx+rA4rxDeQyhM8/vq8GrX4/GNKI94sOoVDSDQ9IwQM
VxeLaG6Q0Iu9uYqoNdefKgTtgmENUWtoCk+3UfTkgyiaqyQpQx3QghW/w1Ypz9wr
q+ZAN9PKytFeYBMx2/uXRFN3M7nN9V4icAxQeQIM9Sd63MzD9pYbN5H6dGr33dGE
qSzRKpjpsoOg5NHZtbwEftrL2dI4I26x8dShySgQiUpjpUs8ytOxJydrfCAdLGHn
0+KR3yXuJO37Uk/llpY5DNtOGzJ3TXyH6bc6L/pCrmjCLXYPSgCW8JiXRi2ezV3m
YiNDX9US5K6RyaRVLIapwKHv9zWYyxvPf3rhsIaol0ZJIuwdslUI0+e0SJl34Ig7
MLNZgUYylAevHaPnJjbQwbQuWt9Ljl+mPle+Vi0wMuSaqCyNRiX4qoeOpQXw/VVV
5LYzUmSzoSzBpfsQO6CJEcSauvPWvyvewNOym/zX+0ZGi9Sd7coeZKdnIBmCeAjw
Kps672OY2aJmrh3NwZBqKfn29SHlQec+O7nR42c94WEPKurq/wlVLA3q6W+W8g2l
EZl2pfG4UJIxu/TqudUqIrzEDJXBCEtbDm9uGzPU5RAAYOrnlrKG2ar37Uim3BOZ
Frqp5uAT7gSH7UEA6g0Gtt/dTc3JGhT2niSCsZmYyzjtWjD5uM+BJ+kzykXxjXjS
kU3CSnNyaIuBHmMXq1C4gRIZzGQhZBHBHBvOMvatcdyMpgubPV5q0W6tONthBzdX
pyRiZUsoRnzBoUJU87QzauhFgeZA26jVY5EIlHUK8H7VFEpEEOa/zqYz8gqchz05
n3fWlJs+nWR7veXwxTuOHr3oBSOyAIJXG9daQVx+asVQcGP7FmZbA5xGMRvPo06r
OMFf6qAbfERUFy65DL3qlmR2Rrp0RF+qhJ5NXeR6hKshYQQJqFVJ6GIZkGpFPKl6
LJlvL3fSzXEjem4vZ3/A3yRQ5p4w52bOOOfR52bBm6bOAdLpbvYuCn/u9H7veaY7
TYwwySKY7xs4LQ70yGRIcpwe5eaurhMno82uDSI2259mh8T81Ajwbkc+QC1xAzbd
E4oXXXyHEMrMOqtkjDrSm0J0t4OqcFH3w0kBBpwJ1X8M/t3DebQKplDiz+x/luN/
wP3yrVDQMdQQ2+1nxz5mmPxYRUWDXryuZppBP4uR6VAmCEV+XCRvFLwNsY6X9+qm
MIUNSyPHELyQrAdtGMgVHC8Icc2gqzkZEBFp1vCC6olV5mbN3G39diIYr9Igi92P
+5nRXQlHqWhWdwOQHRxNW8NMUqLEP0bqgd4AA1cjxqg+D7b0IwkV0vnpKykLX9yU
1clsv9TQ5cFOvgfDwRg49Q2Ws7Nk62IXOiSIQj+ncO5lQOIaNMLGEzvI6zSuWf+k
vL+zUObetpv3LUQlWKZkKrv4HgwWA8b2J41E7XNLaLSYaYn9/pdqri23dXn4V67u
9hiAF5NODzb7GRYZEeWI5DCA6gCcoQmA5pVJR/EHBhQdUH5oj8SHN6O6qthvI3kt
Ir5TIJiVG/svs52iG6E832A5f5Z5ZASw8qVMCyWOlR+iUVNC6mFjJ89KGy5F59JC
1UwYo39E5XURufcy67ltMp6g7B98rH7QGL4wWIsr9eee9v7tdXu7klbUX6UMr91d
Rwlyt0vB73Lz/r4qYJDBMuC8l7s12yPplfFqGDqR0BkV4rpe9ONa921qi0nEBAVf
Y/mK1AXEVPGzkQTMxNGlf7H5nd0TlQ9KUOJpHTB9lvc5U89G0o9hg0e3PATGYNgZ
HBioYNJLQsUrHjpeGqv775a/rvlwBCVtzcVehQstJ5SHEss2kSKyvUx3NvhKXApp
C0uxFdU0oaI6k5aXk06LuZ+h7iChbhu/t0fyOJv2LZk+FqK9Z+PqfDJoDV4TjkS8
1TD8HtzvEx19xpkKMEpxiLWDAhCyR9h5wiNKNTNidUNu2b6l7639P/A1C2sizVZr
hhbtNKdeUNHtEpojIEJCO4KVyLL3e1zVAMlTorSLL2IacZ1CEj3sKrObCKYJD355
JI3HAiNErV0FZk8J1Wz4QjVV7OVvYxgEWSZclgWASt2CbCm1+7awisUee6qnqcV7
RT0Zql7v/c5BeRpKdiwHS2HyhJpsfoIrMYnAgbDrGsGVmP5S52FShOGZu6PfK6Ix
eSrctE3aRshndYt/5qz7vvNZpt2ebxnLfloYRtSKfzF1jfEwKyCKoBny562LGP7U
8czM5ubsjtaDMjHvC4zJ03mNMVkoulId/PdlgwkBUdhNNdojsGvYXptWKqz8AGVA
b6w2DtiVzC/D0FoBn7UQnpQRJiCH//Fjvp5q+PfUtMBoyWrU7YTC1VEjSuShHL8Q
JWyx/Qo/oiVg88MBo5rMzJFO2Oc83m/oJc1RkZZlj9NU6Og/YMxADDBcgZn+RZN1
y3XXNg6PcQ3gfL9+yivvHuht9AiSjsTwyvfJQFendiu+gbnkNAjgh5yoiFIR1nn7
4rUkQ5KaIO8aOYad4hW11H9zvQzxf5EatX7KBz+3atdsGb8Vdue2NRFoR39RfqLa
w/FfhKGHZQP6NaBc2g6uT7xZ45bfzG3ihXq5NgFa4f/TbDONf6fsTZ0hDYcqAA5V
`protect end_protected