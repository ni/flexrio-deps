`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24384 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
hRRAlfE1xLfeNfywbrz10BBIxw6Wt6YaBaqf+6cdLYcn1cCfONlyAbNp4WmRVGE3
rCT9p66b+y9rgc4clHHc8SZmA0VdgiM/CSZr+XpVtM8KWhDkPAhwg9iqgYoJ7lf+
S4aGwjYlvcrPbzLJi/82OO40VI+ZYfIZdE6tHMOX7PzsUVGgBAH6xqE0fuxACsb2
tyr4R2eMtiEFLz0d4qIf3kOghUSwMeGhIFJWFDt6uE1qSexzCKQ7vGUfJTgUCDtv
t3ZgaIUlJ1UhoE7r79Fa6yryr5ZrVauIqMW6eOU3VfvAf8zCEb3K8rM7K0DkehuK
u0lhB/XfwDnQ95bLRgXVDwxFFDOLTMGVp87ctUutFY9hemBs39j9MJcgpRgSTK7M
CsZ636th1d+jVMfy1z4nM8RZxhdbXjr8/fsdrNJxs4herwt054J1rD71zfPid04t
eJSg9WQu30m6xGSmOtCX6N/wSV2zdn2eIYe/waZ98Wxr6Kj+3lU2Exjdutz5Gk1U
Y/MF5a00NVHGavkdA2kjGvBiadQZ6HwvpDGJC9S2fTqqjqOwj5CZzQc2t+fm7r2L
Vyn+zaTQ2bpudqjzoEdzTzl5tiNvPZzt4rGUhwfQvnTIw6LBqWbikyM9/Ad8K4Hq
3PeYt4lNUwCvpq1Vbyds9zd/qjp2ZqInd15QmlDyU1a5HTTk6aNOay/TMkySh/R6
y45tpRSNrr2pZVm2Gx3u2wbfqQP/+h/aUzLaEwtpv0SZogOSCVH3bn70zD80wFI/
U3uLBDOBSAYfZkDWfWrsHk4g9MN3aqdVKCkEGzbS0qgPvUA0dqE8njifIZCQEIoK
JnRY24Bq1jKf9SMPn7yDsR2CpTVKcUJuZlhhebl70FOxZ4MVEcbmMZmMDFe7NQvz
sLeDcdiof4FKIuU8HrhkSzMSO/Kh2/xVaxUanx/grLcNpz93ZpmmFDC48ld6FF9v
eTolCdF+dSd4YiVvvI0o/XCG3LgyWufx4gmgRHYlFIHpsaytqasHBgrg578rRtxS
bn2gK0i/VseOHYuBW7ByNs9Q+VrRdoquhSSxu/RRrebZMFzpPm5kfZw2jkNTcYjq
k/ttMKluhq2qOSQnYsdxBxpACK8xgwxgnBKhVD+VPDqBO0zejwAixRZXwrCSjd2/
3k4Q9qbsbdk9Ypm3BUpP6F6iikrieUeTOHcH3qh0DPWn2RcYStEMO0CjnOVLxM4c
067QA1CJ1qBIfgYVkitQD2CqJ67aU9+THJBkcUyYqtgYXJExjpISUL8C/DQfpaD8
hdkOHRUWvdU9uPZzWG/ZJFxYPYiHKODf8ffFBI9G3s2ToGJu198pdT91L34Jrqyk
KuCFts/lg4smbVusngGLrHZ8XiXREJCh8fTkeQWxpbl+29mQsijD8UNfDXorY/sc
ni76RwZlhhyZ1+5hSOz2sr5n78bUflF87bUtXj/xxUBVs4OBt5WiKPZCAVj8Lltu
U5rGnhXdqPz6Q00AFyefS+ShDXoT2t+DtXthcmxasNgpVIeonNuTgJEgGnjOflxP
z5dnSGsSy/ZSEmgnkmbKA6Rhv1X3MjTl3GRCMhIoCvWgIjaRVTJExyoOjkALH2Hf
VDx17iLMEr+7bHRGRgjYIauVghhyJKl0D5BlYZNzdMXYlep4wZPtbGqBV8PTca/J
NpDqPj+0xa3lnLm7fqJVw42fWFzRVnvgPsu4E+erE6xWc+2Fx4oNlI1uWa6ZDemw
Z0Hxi9qFlaOVMsrlr43PoiYjPt7hnKOpT4Ec2Es5dqgKqkgYXDmlVEG74Q0xN82B
71xpwV4c1b3mVpC8gjF+Ni38blLkANZcdLrwW6Q+8cMNQ3U7F9SZfrCtMfqH3mPJ
g5QwRRjIbUZrYJHteel7ivfQWWXNGwdj8tx4wzsl4z9XC+ptaogVJQjrKuUTNnL+
Ce5LEKu5f41XJn3Ta1s59FUTYz324g5G0QIpCpCJT7yN1bZ3CeRRjacJdq813ZhP
tFqj9JBCkoFVJrjuF+UeEG7ODEDhSukS9LA2T2UcLB/aZ2Ui/dqlmLxlHZn4oxpr
Q73AhHwmtpumf60P7zCiceotYbd1XQA2YzGvD0SAvSHbj4oX0qfa5rbCkb6gPCgr
Eo8x3Vi+KcRvnBAhvbBIoXdwx8hcW+PdCAZQ2+Ms8FubvM14Coh9PSrJyPJASNdp
UlRh7bG7FtggHbwfX7mMb/9u5VKEDAhQ+6WOIJjH/kDHrln62/Y1LhpZJWhfayAL
zlQstx7Lt1r4fHEY6PJLSADtYiprVfP2+HYyEvR0/qF6bAWa21057vuMWuBTc4/l
Sfj1i15X0M+V0JvIZOCJwEsTedlCLlRbSvWO4sbyRX2za/jgZ0vLnn+SGH+ksqkg
WipoXtHWYasN0LuxGSHl3glAi9BTZBC6VgUWRrKB+ll0ugohD/5o2a9N6/5vP6eE
EUaw8Y/Lgfy6x7Vg8ib+qLgj0LgWA5zVtYXpqOA2/wlbm9vTaooTvS5XYwyJd8Fh
bI+H/cNbwX/3EIyLeHcvaEdobZDxMoV7CftBPiIbV9S8l885NeZytayUkX1zAwoX
3eqaToLxGU8pGqxQG3LD08QicPrCcnKhVTVRHtCKg55KYm9vLWa0d/YgOtWBJQJ3
RipqY9sNp5LoMByYISWl6zfF1fV/vUg4tl28P3EhhC9cka98V4Z1G4L4HRXOhjxZ
t5RMVmG4swxDok7vnUurNSeDajPZZoiDS0H9d1ZzrI+EyjWEfnACyQzBUcQobq0b
+sMbJiCz/Tlq658tHkJ/ace/uL7W91FKO2JgyAAWAio8RtFJIZ/AqGyiD0ewbwnh
eK1VVDV90C27fX0VXPPRFoEquL4vFtLRp3LobRVOkDXjNtgK46AN/tASktfG1ico
Mf6qduDYpK06KaX4mdfRQcoWcIHGd6IeNJkbC2VsIu+Kp2wtrmIvBdRaAeXNN0yS
gLaD9pSlVBfN0o6DBxzrRATRNwxceQRZBTp3eCENc3MnIstyLrVOsDE98XbbVmoz
b6B8y7piiQOPzbosaaOp6XhAUcbHk9pAm3KmLJTw0egrYwZ1yLHk3s8Kd6UiLwLJ
qFgNkKrsdv3kOADKEK+cBW7+bjQN4ZgXMTflDvQkE+UJMfa6cUKy8HzMF8qSR3ET
qEAqsKSpaB+kzjbyF+gnehaqmcQ29l82gXDzJIe58vR09qRXEHweqFGDjg2Ld42V
mK2hSTK5Axn8nRWZ3FSQBVrxLXSuAGtTsBMn7Nx55HZowRKzWZC+Z68/FVugh3Tm
pN99sU5q9QxSRi6W+9K1iDA604vZ/9PYr2YRTL3bD/EYmvTP+8x1j0B5/MmdRAq7
tB6Mf9awXUTVhS59gHf9glJwaoJijAzpMEV8ECKoMfXYdFKPG194ETQzpxS/OWdN
ffaTBOCPi+09u4jQYW2JjvdTqNXhNYcdeqnyTbRSUaonAOwfxskSpl3mfqd8Vc8D
jfN2TPm8SOhpLtiFBS6fadKEFiyhPZCryC5pZZrF3pgBX1ZNgrJ9gGFr8rp5V5WP
P7TjMN+86vreW+AyT2eySmpIa7yzbSudxCM+OIKofyqUdbpL8hDtOTQHmhzIZn+U
zA1CyLuBC1hXzNcMth9LcGZNka6tWJ6e9mNyZoEKjlRCv3mNNF8qNvIpFAVOMjc3
DByVQdz/e2sXfXZO4QkUED34gbpVVjhIwqpCfSOYH5uoJH9wjGBbI2khlyxXvBTp
ebx/iD2+PexXKjcaXEcPBeG9yiDriC1GQ2fCTRqBV0Oc7g9GNtcGNsG9du8px4sT
rYIFHw5TCAZsRxcHJnURhPA3g2QX/tc7RQw0O4SLUt+wDq0MCHB3QqrSbTWSlnAc
2T6tqtzBeQFqlk3p0KYrrdXfBJTcL1M8/HJK+UdMxJoi4iRMHpPz0bT09NZ/eESx
adXhtqUtn6Vt/6NYAVRBwIuQp8wrXqXpAFNLxkBwBPqRB2R6nIigmAn55bpsdh2s
EVBbUH2jWl52NsDHh9oMZK1ATdZF95LmEXilpoL84nujtagfyynhQ2m3bac7VUjZ
OXtgXancJSvEds4F+LEUKvG1Una7A3ZkB3bK+v4a4kHx85tZz+jk463XTt0kO87d
6x+jo+XV6RVbgRJmPVcz0JGTN0US4dFv8TDOQlxjr5LaDPzdQi1TULJ6gSYlGBGA
xmKAVbALzPcTQFkHnQxWUpSZGss2uj/mrX7fKkhOmcaE+rBdaCADXYrnUqqIiXlT
g1nlCWDH/L9q441St5Q82APHsoFznWnzI2mcDm8tU1wy7QdYUmT4fokJ75rZv/Ok
/EWF9kF3/JTAzDnZ1/2VEl87dy135F23h0Sd5hTRH6iYgAxG6kcq77amKIg9/pcD
xfc4AjOCWHlLMACr0yObPFHso/PIudhUSGvdoJ0n9VwLWQntvVLxklHGykhchkKT
li+5H9qULBoHqsjQq5d3yfeAc1BRVquuPH6C8Tx5f5l4kDsia9NPovNA/VB1djcr
CL88zrzzdW67OrrnuPUJ52B9y0+4Rgv+5BoeBmYeXsWY2GZ3bdXe+NJP8eZrpgyR
amS9cpaPKFICzgjse9LjnBVI4X5ivqHpMFj22L4GtrytZyId6GcXKQ63zii3Ipvn
SQq2fTr9s6FCeqLkyyv6CcJNvvj24KUgk+LFu9kM0o4qKMwpTuphwDNQWcD6pEsk
o/BFHQoHTqGuhAYP2YCX8z5MaF9MeTGw5Bbqs63QIgnO0w8QvPiduU9GcXw7lEqt
rDt/C2cIrXSFm0h5KyQ1Y8caIpYfB87T79MnOSsQiZ1J4U61qKvVeYkjuElANlso
rcJOuQwSUjmAfc/nNY3GdiprZlLdRBWAI66UoBRkSgsB0OADfSZe2YCqLf3VAzc+
aJIdYq6Kb7zBsMdlUrDChDCmI7Ftm1ll+SN/WQKnMDCc5nQq7XhkjBgNFSj1MdJw
U6YcEHEPHCsNl9FzB4XvuPGmqweDPoNCeBx07UQYx/+aMYtT27mJcn1EQKwiWKtJ
zZQvo/GApoxfnOuhPUQxkwmMe8co0oefTov8ksXskatQEdggw34wVbws2Odx3g9n
Ul+oKLHItqR+P6RH6CJuEM9fa52A/JJW2KYlBEVvxxQF2rrnoKk3jpJ2ALAH1aZg
2qTFB0TWS+bPSwnkCP29QvOU5cpvgYs4Th56X8eLmzG58+bSRQj4ANh1bV3cGmzq
9z3QCiLY43zpBhoVLXFFE/R1PPBcuRHlpNyTBdPXC5+nfU8KH4fEzxr12BHxyn8A
dbMogKh2jUWtzW9OlY4vxmWzwaTTfWCR2DThMGCgXrhs5zJZLVBwZdJCL6DklEco
+qcUEYtPlYEJ8ZvXTq9OqPocjWHna46sXgZXowLQpFWiH+WivI9KgjMBrcc8dvow
l/8oDwqN/+P9Ye3LzgboY1uzNAinuMCtRfK08tQkxVnnhuf4xWidmcuptoFqIo+F
voGrcmG9OCFf3OjIOd1SEakWdpieeQGagBwcnIwUkzVHDe0WX8Sc/XmaCee1VnGe
aNRj1uBrp2SPHpnvPrCJqCU3l3osk8iJ40Njqvcwlk+YD9lnOSbUQTcIYGAlYxQl
beQlMgfY5eQZ718lFF2ogliex8qcXkAdNt1Js438PQcWbMDpnfuBObjwhycNM+aH
pGHGeYuS2GoUPiTinrT9hU+wjvYGsN2L9CW8K2GJCQZbCBOq9sFtsLqrPoCJmCvS
EWRMM0Ry6gjleOoxp+ErK9Mh0J2atWga84Qu/MN5UDArAhov8/xXDDmpZl0ErzKu
iuRoKzPQDy+dRGuzR6IfV14GzRP060H6I7ql4y/YdJCv9xTyMUzt/N4ApzgyA5/w
hMXRtHaOUJoVOhIdTitznP7JkijAJfWdLaAvGuzRi8i171VxIKuzAvtn660ATgqH
n7Vm0bClNYg8OhiB9/Y5bt3HHLAdjPCfEiYhwyxolXezWeXvsy9J1IKHWWLql+Ip
5erDy+/JYSvcRaATvXCjOMhFuFNvYwVLVRt/tCRRbQbO/C29/fQU+ph27laMWG7n
2JW8s+FoZ/1FqOhb+YNZGQAmVXDShjJYyIK9X2Z01pVytqGYeuNcFyZlnWbe/gIw
SxeSOlyawY9vFhBNOXAZXBRc/GrzoquHFDSRnrG/H41Oq+djwTnge2xJrUgaSN1V
vm0E4xl6ZLiAOGfMKgTcBG455jePuRo5TDVD6uppiPRXa6uIqKP/3S0/Qk7FR0x9
7vchiXvIzswTR9T2cyFdS+xBTdNLVAucLHpf1V2uGTNlBze1g789fYrWnlQk2WDf
FrHkPJUy8LUppBCPWJGkecKFvk4du9UGYuUSqK1fOAwoEPA/oi92HobXTKa1l6m2
xafAoY6CKt4b0Gdh/I2ybV6zFF4vQtLU7fOEliSSQ3qB//wHrqsed6FEIYjCS62E
FzrcSOBYSw8LhNEGs+/MdB5kyPyuoC07eODYLQMqowZDerhm99rGm5R+k3vkZqMP
mMtsYS94fwv9J5Sv6oI3njKvl/19qE1idDcTJa0xkwfYznS94e4X6257XxWIpMPW
Z8QPeUuXtnqmkOnxfvgJk4MfE+bUWEXB9fXwd+Ge7P2coAfVL+qZHYo2KwwMATJL
R5P+g7sk05zgkT3GXPk926C9L152mOUzcT9/WqqJq12PBjmpDTrhYQ4NvdbEToI0
M6TsTuNaWdnc8Kq0St9nilNXy+tzqG63XPzEgDlGjl9lM81odOKr4OScgxkfmRMu
lg5TRjvPeUj3xOc4YFZpA94zPKgtXjfOGm5QMsDwztc1ooXBKYLRX+P8VM314g6e
H9P2tgioTlkukWosVUx+zE6yan46/8Xk0qka0oZcuJB/qh3Dz/7y1OnQNUqMW8qP
WKi5KV7eqDmkmrPyCGoUeSqHLsEGTAL91Vw1x53OlrtKkvhHRx3diSSXYORx2Tfv
eqJfXneO/9EjxD/GlHp5vJfOD0KsO+6iU8nEWzRZDb5TRLxw3CG3RPBdeFeleTAJ
M8a4Dl/UrgN3Ww3ZrX0NsW8Mo8iivT7K0WUoyuWXfMhGpAN7lwJnc6DYA1s1F/Gl
GoePrcb7wNN3njVclPZLWUjbpqkhVf/+K2xeVnUl/sUDAWmSKxk0rY/08ClDXbaI
hOD1mz20z5lbajk7jEmfRh1ltUt0fqamXVRcLYZ2DNBJE7cHabDs7RjdqIOHSlMp
ygoixsQZetxtcaGWWt7IAZOCZx98ta1Z7Y45PY/q4xg5092yCi+2reWgANvNB4Yj
GEV/BEr430LXO/9eDuCffME+mTGM7WBykLs5snJe2bueBb35Sd4FJiK+q4IZ0bYX
41xDENagiN3bIgXbb8IuRIQlLCEoRmdQ0p1uzgGXxx3oQ0Suf1VbaebgblvtHM+P
JzkkMaZa8dNZ5pDPaqsljNo44aEQT4zCpd9ihCj9LxsFI1FWwWWLC1QWgKWaR95S
arWcQKUS9JAPbyGDs0oOqknA2l54FctRubN1M8WCZFZ9jU+PU2dqlOj/YmCWhe3S
7JaNJcrGbFhR6Kx+7CzDPaNE08N2F1xdwQeGlxNxM+xrpolbpovInkiyzSCwVKIm
I8lvi181C4C+UnP8xLHz6H75PuWpB7WkdQAHJqWu/YArx+Iq9m6sdr6ltge+Jt32
pPoa2wVX0c/Qo+j1eX+ltZCTEek75YPkYnenQM0n9QMJ4uhgdJIvkFC4rc4sOg0B
0foM5om8sRSPbU6WkCDAXEWuwNX3+n4JBD6hnUvt8eahAjuRqw7PoyfP5Ch881c7
uQxgEYiKmmm/gmBPj6+Q1hivwF7WnDyvTcqUKSSVly/g8qNweHlUmznZzdFEo8Kc
cSSemKhTjtlzTEbHql2B0vTR+NLJJ4swJqKE88BKSaJRj8cU335jdM3g3WtX/ygr
aMgYvyJCJNGoVaaoLsUeoe6+/q35f/CBeqevcskiSlap/OuDBazZP7beeCbln6yS
bOJ3fhsL1JB6N1oQFwEJ9Y/EhFneHUaNyRJfiyu4jaTyWV5tNLctba0M/WGBwY20
vRqJAckKVurSwIStJOzbnZZO4hcAXnd0hPerHDKPJpSFMfWcYs6gXlkCsUQtq0PC
tCm2zfGMDiUFnpjpVylriC7gUf+MHptPS5Un4UEcsXMVg2ZXKii6yZCEMgUWzA5M
wz6GhNS/AwxwWcceRktiVvmxU1wIezFKBCeE3u683qTwWwg2hgdJYuW/m5A7zmfe
QZBqffAJH5avUji3Even7NuPrmqjXP+z8xZaxFd0K140Hybe6/66lkKwjLjGvD08
nCytAE/tRuKN37QTGR0KsECBO8O42ITb4V+2HF3UfxFnuerPy8oWvmHSdAJuLXte
twsHT45ZcycarnNjoaEZ7qlDWPvRLwREZVYyubnKOhng2hh/6WSOPFRWxBSHF2nh
fED0id6U9VlGtES8vrOlJjZyPc11ahOGjEUHTClemSqbLJwFf2/9SbQ3O13wWctp
NWX3uG6GU+CVFyFao/zpoh4lwOBXFR1dALINWXVKhffo2NGNLUH8z+d9T0ZwVu9W
/gvG4Ojib80VEnox8Kkept1ynUt1uu840UJwZB/hO+I6clK/6DWw4iF9ws7qRrh3
HBoqC8xrVboloznjNQqcOnJfavWA+wocZfa1KkGa96+HdFr+vCP+kH588xDGRVvR
a2IRaKrbal4C4pKSmYk2ycUkZQ9aeGbScZcjD0h2Op6QByLlG5/mxeTvpBn8VQlI
rikZAWtWQE876G7ueEvsX5fvYV7EOUVmPm0CPuqk/7ntgWSpK/F4tBaMq45PRXsz
LIXk5a+KtQvpeT7UQA5Ip/VpU0x0jGCv2eWMbQgICFqlPvyYU+t7mCm9TaPOKc2X
OTi/iTYFilzW7XuzS0sn1GjUjjW1KCmFXIWVB+uOyAV0V5pJuhN2SZ80q+GRoGy7
iX9F+nfUEYB9hybk00hOqvE8MTpPMitLPeLrs3lBKp4WJT4TRarte18dkzhICTmZ
F0GusNRGN6iMPHnSAPqCNzbpIyTdfXnvCws/ND1RMM6BDd8POYluki/UYBXthrV6
DY/1NSZ0Tl1W0jTlUhNSS8P4vEP6MxDLqqGnr3PXMaokT2Z3lnXBTfs2di3qbwFl
Zs2e+7uAFLMOb2wzvu3rPCoh+woALVhPYuXbv2sDDcSnQQ+L03OkKfTmN4gPy6gr
tL8SdIDsjQ2WSicLKS0HurjFvAIE4zEzFtX3jWQmUWBWU9SPyUQvZ12/BlYKroaE
Q5xM+A0nmc2yy0vyjFownRpJFm2LfxkVBWY6QP7XPVg56vSoI0RXCm/SNeeIOq+M
+nofv6nrZlmuwXhaVqJRCWYSldhZuq9DQ7BAN1gAgc55BYedwy3vqQdXxi7zgNkc
7rii4SzGAUBkd0zT/8azycjPiF0rzbZyvIybvFPkh5+agM8nT7lUOhy6aWpqFQmc
TUKKv5Wh5m3eG63w+cqIPqo5rU+QBu0MQWEYtZTSgQcieMFPZrJRZPqlw+6LStMh
A/XIVjnh0JFInLNXSBWXPzClh9gSeyA8TZ89+KtGbuMZo05xgTIbeocskxrkWOSt
65tMrppG0kSyNnZGppN6zqfq9rZPHhDCZN7wYIB7tizc8iMYpIWPgzrzndWgZJ1k
0eLDw+KlZuUFQAHZAzVBE/KM4AH4TnCI2TSet9eRb52ixnIUCWze4pqkkDrwv8Uk
+atMKc+XHusKO3ZSk7PNbo1pTjNfIO3CL3RgepkPPEGdzBs7fAI3o6Luj7a3kyy8
djd/6SZftmT6yGIL95PkLLB7Ik0mwpY3Y/vw83o314NOdaOsryBnv5C7VZUIFap/
IXHg2h5FyVPHOl8mnP/c7SqiOAeGtQfq9UfTs3R8JBcDCMpzCAdgOGnPscT9fSW+
6fcagj7OBd1GEBBUjaVyfOKSok/uP62gDfLI8VUMQrenZ9r1KkzjLmZa4GMy8/z9
F/CGKzAxKu+wHZJgIFPxwBEd/px6FDU5Wgr7eo0EcuYM2p09pscYuSPAQrPVOtY3
ULRpziMIN7Div8hQCZdelMH/DgPSXBHYlNMv4Xm4fq7c+8/Mk6qaHMb8IgsLx44J
zJDggcZUt6MMGVNuFDTRp3eldI9wTtHNh+ovT1ZpQzTZG61qSMSHWeCan1D8k9n5
CEipl2iglm0EaHkSaffuHAiTPV3ACGWUX1nw+MlX9ckvfGelQbYuiccsPGBGa3og
1usuk6CHl6eyVP2CXFqrH1gfHeBwsUBJKELQk6PysF3RNVc9KQLfmfVsPjNuGkZc
6kaKM/2qTOtw7qAza2koPDmW+FqzwgI23CFMXvH/oe/YdYiscSNbS+e89Z5ZHgQx
UaMCqXaAZZX9yxzKmSdSKAQ2Y08KooCwW/rSzVz9C6tMCQ9HafwZvWEvJTpuMUjQ
sczPvw2mqIwgTapHKYzxyRSJKE2pieMVwfuYRpw5cjrd7asA40QPbYLEeTs1FuiR
PWvPXa+RgI6fDtAFsJduzZM5SJkg77xu+DUjKTSkI8zPubH4Gr9MyxqxAFjsWwM6
6cVwNZ5eXwYknnDT0WqJNAhk5oRQtrtbwM01Ew9xBSEqokvsjOmTV7QC5uvhudW1
7EgwvqWpRypajq/PDE6tAMKjsvwq4aHWnenl9DH8yEGb6gO5GDzmLo/xWaS5QFpX
y2iT2p8YDLNfdi/L4zfPeC4A718MPOanhbHT9qmBBfKxKlTZlhH/neWwJfY6OOt0
6MMjt60OWbvylv5/AJD89GHEOdbdB8y0IRPYLxD0+tGT9WR/pj7RwDS+8N+xn5Dx
XRX3wdOsUsY0/fq1dDAO/OTsatme2l/9DHNPZhguMOhOPbWxcse3XlCtwPkmXy0z
GFbRdpvP+/858t6wa5n6GywgIinVIH2zNz546aPWCsi+52K6n4ifFw7r6GixY/Q/
9LElLHnpCCyXOBUCwgfpIEbdRVg+RzM5QeKTy/tYCP7uFUR6vC7/mL2Os6MRIBiy
qT6oO4HC5ftR8JMSwb8D8CUa/t5BggQBHshTD3B8TsFCT4fKDyludmHPuSwIpH8l
U86X+fqD8snhdr1G/32jxUamoqGE4ufYimOJV9+v6/0TxS7r9nNCNEwKQcndYOay
NoFWbwD3Dk7sc9Zr61+SyGGtDtJ6EFKlhtNcxndLkyO29hU0aOjKmNh83XBKBuMl
Kt+BCIL/BbAKDwd1PAzKxKCSA7juN7fWz+0urUiFTgrNxkvQm6mO8QnqoEUPfZwz
19IziNjt4ojFwfvgX6zYW5RDyImx5j6TgdPV40S5ADbyAnHBfp7eBFCMHgALvSKQ
wPCCb1UpSmZkQatqhspipKeTDxlpd3txP7tI2uEwyJH1WUZ+vgPj/G3J2OFsObvW
z/E1WGcpj3GlEbywB7RTBiNse1rw4dwrZrmCaJoE/hQB3L+mV0cPF1Fq1Om+TVbc
DIsM6E5yibLci3b1X1ngsE/LLed0cSJINnuHI0/kGl1VXf+8fZ/1v9Mq8nsHTytL
cT6OuU+JZQycj1J9utvflg5bNNaS3wiokFeQCwRDhi6TxcaaGK20PKpCjq6aOoqZ
FHmuXwZnCbsRMqnpFY0pjDFU8FGFD6vP4Nixy4vT/Hju8tqY3g+T+HXHjBTHozKl
W77sFOHQNAJ9aCBAQp/vuG2HV4A1ApfcbnM8IG/VlPuIEBrE+MFN+VRvZiset5nH
KklvEM4UiDfYgyDu638HUVi8P2DkXvcsYHwTPMv6VscAA5PoZYNy02EYVTLfw/pl
A0lBmnUKIAY5A9GgXzXNBCfZS60HkMQhMSkCc0arQK7U3aQHx7obLS/QR50ZDKel
t3GGARD96MKv6sUeDPvsxlOMRAc8OIYFFNDDEQ1SEdGn0Evc0b4caw1EetWn5WDf
FyxqTF3D97e70kZkYCE2zoig4v0CFiMRGplzi1ChvmEWbY5iRZY6M/RSUE+rrFrw
KZwUr2tge8kdVc7ugVLfCqSnYllPZ9hWBpjV9gtRe7A7vIXm3m1nVqxxhHSBNK+j
YxkI08kNqKp5Mro7u17hM+mJ3Ey1lhWG0ktSmjvOktNcbv76KVqj1AdQ2hUv2ZUe
2K2KPiorSIeLP1G/zZGiL++jnV0d+fDla4WKA+yVmtiXvkCII5pM0zzrSQA1UVBC
C8m9eDgQm0sD9oThZQrAugupbX8vqIpBrs97fC0FpLMJjcVr/uG41vyhshHGxZJ5
u7u46HvmWIT3FANrVkcx49dF1INyNq9oPHtlrBFKyo9gfjZL3XqR3mwHuOh4fHEa
NwwA7veDXi4KCpgz3COyV0cvtFdiUlfHxd9w3nUteNWM8LMjTgpCDRzVQ5Gxp0AY
QEuYi8HBsY8YL+taTSM9dNzj6ybsxC+k1mL3GpI0xZ6U8HDNwMvbcJQBZTPSflN6
COo1OUuWEXlAo0d4+p09HCE8swiFuxv0+53kPColZn8CBF0oad33aItslFFNcjto
TkHHMb004KeqEhz99+J5t05+Hxz91rhJlKFny5xBYdR98jXKvhhu9mq9tu6wFkRG
SEcBYHaQtqyjhGxqTBqHgn4xyvsl/p8CCOyu+HCdUZQDv47jxgH+iNnVcMXNdKZh
NcxoW1cYA4S42hN7NcBfkAqpLWZ2H+NC2IltZcfDGqS+tGccBuCt4USE+HwseEoJ
eXsQ6ADiz5ylGncCiAcVbXnRw1Ruyiiz0vUBgaAeBJSAivKZEuZGYaIz3LNNePOy
f58O0x8rsEkiFE1HvZqqOE/Y5oZEZ7S6bgoXKPQwZmrFUyc39r3VzfiYn49Dy84s
nNPKVM9sSLC9f6/1eRu8Fr+CWzDMaRBeV5duxSrMSF8Wvn+A9+U5+dgvKNYZM9s4
igbByceGu2YdesZeXiYCKnpp/mxpe0w0FiNDgytzAZIlJJ00FbVKGFR3yk7iIdBS
ipzyg/Usp//F4TBSxJGrQq0NdXele0WdjnKf+xZ+uDF/U41jqSpHkcIRRPVnkIEn
49HZGDpb2f/yCpnodcrfVqlaOi2RPfsUIXRQW01uuxk9Tnu2cXm/DVCsV140Bxp4
S8sHLZ9pgsp2kLGh181ya8ext5EwLHVNmmBShiFxaASTKaOpNl+wI9rGmY+jRMq4
LACIg77bXdIbVK0sHp7/4vtXH9BZ+c0Gx1Zkl+EiMASROsLVU7yQXA1xYRRETjPZ
Xt1x/MqIDnuKCFAwpvhGnEeu65z+hgmfNL4Hjt7uNoQ4hjXo4WWD5CTssylbG8FW
VdcQqNnQiIo0bJHQLWcoiqRETHIDG1yIvJ1Szlqo052f8PrlFPtqDftsA+GuR65/
Bf5Z0agkORBjfcY47MpXWfpbopEPq4Iu2fvjC+7QVFSvMUMM24dTc9QP+ufyFVic
L9WZ7y7GKYMwqGljAWr5tCkkCzih+zxUyMkMpw9Dc6w42Bk/XNFDEXeqhqVPxOp6
LPjBqGxzG3IL0PdiBq1K1luju4ff41/1RqJyAm2k0UFeWj8UvRcmNiOoOky7zwSe
/8Xj5e8aBNBe83ly+DrtF5UWxKm7Mw2ZKTqx465TllBa+JVgFHafmlSpvnwG0+mR
7k3q06x1wL66A9guXLt9QEuTETUzCfZgGzpdqux3mbmNN/qcdfect9TCr4T/Xnn3
zAT/npUUY59f5j50rkXyKqJOxRNb8Uc7w5leFOmkrhAZFKgaZifp3FXZkHMS3Hbd
H29zpvnsfCSZ+pdRW53eLPbUi8vbVlu072dJKTiaWlisup07AsUjzDIaZjg3AUyW
L1vee5W6mwBG/N2UiKWSCG+ALS4B5cfXwDE01EoniGKG69L3t5jJ2hJGfC/RRm3/
c7YY6h3zTWPZXRHfYwcHWE8rtXOegiiWV/Rqbt8Y+0+hByRtW91TLCMKAjVb18Zk
6D4maHUJC0reGa6DZfbPFxGdvMMp9ADD5INDqd/vG+fOn3jE1FbzYjGl/vmaFxM5
8EM2eKLl90hYKM6Jmj/0EYBiBcpcGW9+nzk7CzFYcEkb0gxUL3zvzCRmVjjZ23dC
cNY//8K0fjrZ3OTAb/DLY6YbHmkvG03wWYgXVKJMsWhqCfRMQTxkigf828yL1KYk
NBn7FVXwiMvOe1NoFVgbS6aadhCLN+SH12z6dUM8RVJ7qCa2Z+4vlXbIGo8Doxge
R3HivlCDTYXI1cdlC41aDfmVsX+M3w+Hi2QkqCklpeQU/nYZXPpvFR840cb3caLL
BMiV1BwvcrFqSLwuP2RhbGMjkrdqhBvybpM0/xpvps5CmqwYxGtq/VS3gce+ZxWg
15oakFlBEoyL/GTgLlDZ9rdg3tFd5NdQCByak66aYpTLG0JhvndhH+kOvN1ZaeZ5
TTqOTFp1I4PjrHfA1Dv9dkw2iDfPHnppM+cbKdoo0d7ul/Rn6KhOGu6yTUgHFGXp
Q+nNzEPsiIdT+6uuQSBBHz32t6QMBUSBF/krGQbMvmtaIdbzg+qXlp6xOCMhSbLY
qi1M3Jzaxo/Gri7hMf4W5M0hQ7nkvUqKuNCND528N1Q4viwiFt5z09pEcg1W9+XP
atb9LAWZe5unO9UQ+KMz9bxpO/0n3AzrwdC5Crgo/63YXzcKvJbM/udXois/ro1t
eUTyOmuIfNnhf8zgsyJ4eo5w2Rmk4kbcIoUogMRyM98EsvzKPc7OV/7IbR5QpfLk
eNBxBq6hTaGl5Gz7SuXSsUunGnWekRphByC/BfYsBpVbZ6t488yGZzd7yzSJgj4L
cAiUL++I0oOIhtYbbyPzlO5lT+PUjLUBd+Buyb4unT4hcdnYvVk6KsRGFSSyi6qK
Ktn4v8+Uwb/+rmdujNGmEGN8mNijRLbE6z2cIDcHWxXni4y6k/kZsWrcPahdBMeC
Ijfayhc9wCagr0hbfj5uRY/5Oee38NadF22vdonLx8nL7NOqEnYpQ3IPjXf2dbXJ
BNQcDb0iIUOjrhzhOH71MfippjHoJyz0CsZF29KVqkf9Fgym61lh/Ukw2kWfXvf9
Znp0jwLk/fkZJjWrlTAVCSmZjh9d9DD2bM97vwJBB/NnabWorcNduzRSBJ+9Cb0v
fh8k57OqwZVCC0XFGbb9MGe7pZDr0pUbJa7mjwYItPh9dX8CEJtCZZqDHy4H3iNx
B9QiQ/Vw7AQ+F+aTfi4ppngekjlvi5ybFXMDJYBfU4/S37A1dNjfQeVuwPpPuntX
6UAtQaGY+8PE+uBjg8dptT7uPDMNxcNtzRGtf9+mKiPHy8Rei2NUUMvopJO1lcN2
5BX3ML+RgiURatZGAh99IQLHkxSTDuLly8o2hIBWnNgPV6waIAfruwfLoHcvX3RC
v7lep/itigzY724Zt341F5wXzDsxFc7mgl/vSjSx3KvqSIjR6k/+boiHNjrnGd7N
qFFWlPL0vs9y8QElfTnoGXdhyE6yD61YnQ7MToEXIGnUENNDrwTE7qkhElGNmTfH
TK1wXEIDu+n7G1J94i35bBWsiRVkx3oRh6x6jrOmcsSPxvO0Ap4wBvizEIviLdYE
V6RKe7XpSjBXUvcz2tnIuiv2Z6DcRa/ZQcVY3rXFM1xyhtGMmx/AjYUOwTVw0ydd
j2doO6oSFUgJ17MO+8vmykGRGC1OwB9divsQgmMvt0HEOeKBO9+2zUJS2hEvCUWn
ep8Zb0963HPvlkBmP8lXmP1Mb1fYMRr9w6vlqvNlPh24mmJ5Tc2pw/olln/aRy+M
HmVwfelkD3ga9sQbdPQIsaDM70QEhvzU8kDw2lD98CdZuYKrURJWklw7erXZQvER
4yAWluJ0YHdA+KR3mqAxlS3/F5AOsSGCwB2WFxE3AyISXG92/rqrOWDYg45Ym+G5
zxjHlfZ/p2lnSqWs4uksQD1eUon0KOAnV8HHwdDZ2yqWG+rwQX1R11mJweF3dZ1o
z3ChZMs0ejL4NTosewpTAk0uVY8gR1MqfYGk8uStFEFjkOpnk2h+CFijUB23bWHu
jJtj0iwc3z2wKCeJWbh35pGWT1JiVgD290bnRjGVzOy1ERiSKErlIp35S4tagBn9
G9eFnntyFb2j2hCTaFeNtGaulS6DipNk/pfPvCvcBGO/frvLQYV26Fyn9unUtni5
0bbzs4HN9lwiL+lLo2DSjwRzK4OzF32n/7+ba5n19X4YHJtgHrkz6A20idXQVcr7
4kOFKkLmC3bUC2XD/gWS/H9/ZDT0t5eAxzyBzj7fVoIVGkTGz0nFFS78jTdJGVmw
7Kyx0iJS1hn1fBgOQ2ZBVO0kKCHn+/Gmz7mXdtMxfahOVeyofW0RJfUQagdP2YhZ
rsCrQEauHaqwjpu5bisKOdyvqWk9Cpg2xxgS/q/+vi61swa+hQ9HlmTlLEEdwTjX
pafclkSOuZ9heBnyyV8o2dlMXQfuoCwre5Fk07gXsl5b3YAbPG1cfWQs6iPhc6xq
PAsuMtQInvLZS47Q64zfWKmqAm4v2VB6ciVZQQL3guT4XQYQ6Xv0fG+DhrO4yq+P
xe6LJGy+7nlMhm9fdTpwXUhhI/WwCshi8JgCSOfoeSz1P2IswY6ex5zrgV587N4J
ONSJi00gOajiapgnQHuxlDnd69pCOV0aBBrxib74cD7Q2Dg60BgJt1I14jMQbXEI
KJlaajmQas/JqoDEJwPzuwlL3dZ/b051YvhGDEQSrsqC9pWogjJtbdadExc07e3k
yqPv3kjXAooVtEkc3G7wCnekgI0E0r/JJRkOM5JCrRXqJY1DLuXE1Bs8qV3j9ur3
H/UWgYDPTFzf7+XtPATZ7D09FPgjtGKhlkPdKJL/Xi7riqstRWFgXasJ591KBSP6
vtBDj7Nwxnll96bMH68+TQTXaghpvEKDXU+Kc1V5qFQZvtxodfY91X4H43K2LLhW
IAusrIpBUF+l8moYY3BKV59IPAjWwpPSK3g5M5TwKEfYXAjJg6+vgxxxNLjFVHos
xKuNFBYb+503XKYPUhH6SxM8uJL6RuLXfX5oBIjzTuNpxN9lboMM7+cwr0W06yKX
SJD0NkockCLZRASLNjOESJOouAJhoQxtpprL2hmaVmTBLWrmcarCApC4hHjwlEAI
S6Aik12wC4r7p0+HcPFpi5YALZbAZ2wqGIqCbeWEcfoM/QZc65tv/OQdsdWzWzS0
6XxUdh2fCjItqt0r7PayT9iXAQyJmZX6TWSk4noolUorvzpYaaur7we0sBunLMU2
cgfDLk/LSE2eHTVbGJlu9JIg9+Zb1X9MFWVlxltJaYRMTBynDJDCJiJoDcIj9L//
g9aWk9LwuMXD6MfzzJkZOS88svHqe/rkCmpTKZ6Fgom80+wHfwXhHYW1pRt3adAt
y1aqzzZNgwqxrZqHfhfCOyPeciK5lHblrj1rjL0oULpz/vrscV6WjQlhXzwHZe5I
K/T/OSPViMVf38cCqjTF+2czazyUqZo3wnNVIHmwFrzfmOiIA7Stf1CYIV8fx4Zz
e5ntwsVtWvOTNR6YaL1WEoYiCuqxSMQvcrLopNlVHpo+kyL/OW9apI90/pmUsqhg
cKcVb3N8uMjYbMPRXgDNMp1nWDgDJx15Z3fv2Y7fg1NVj/CfepXdR8/TDiISliek
ggfnMCHgElRhNRGWhlgAVI6xnzftUakHjhCjrAs730fO4bGpW/skvK44973VzmYe
PtyDs4DXLxsyjUpxjOWtshiSNtY1UkXtFirvt6sZQkGPUg3r7kR+EouxjMFlDNE2
4xQUCcIO82bGdlUzwDIG3W/8Bvqhb503tJ2H9W1rRd97gfLmk9YcepHRYDfniz9N
s/qsyuvI0EwC84Fy+ZQwx/+aCucyoKMtQ6AEdA0421SIfqrL/LngkfTkQyN5HsbX
fOs79gXT1nTifVi96yw87HMC8sTXaeHu8BHGCXamMoCvnCHiKhCB8GsLPujt0Yuk
f8O2XXqVKtNLnzy85ANtT4p2DiGmoVWoF2UhGreAvFuHZOBy6xK4sOI48IMkzEEe
FLdkprY+VoJy5R4En7ZhKEBiJ4AX6Z+4yo233pD5k/vVFX3+sQz85rJ+1hb/G8zn
0ydUX3xlVQBv4pIPkzp7u+pQwmA0TouBDd56PR2BHPbwPT3IS7168QXqx8xInueg
qWvv++wiHjqwfpYcqwaN6mzkw6eB4G2v9rURRcagG8oYK1vQHU3KholP+57q4qRO
fQ9eJmaDJeLOttlIGcbBhm7aWLGlSD7qdDV79Qg8mxy0xoxe62gWyQLy5tTAs/6D
tRjF8PmF5Qlw6hrNQsbAJS9mS9ixKpNr74q79GfkIVEqMaR0jcipomDA0jxLDjBO
RBxXlfNucfNfSmshj1EBeHuZLSCcgwGYoz6XepwWn55VmAc4BgvOd+0n5684dOJx
k940fh9hxvd9Ekrt+M+8h77ffwSUMop4uwJNaXXwwDLc1LWWiE3vQALTRzg8wwTV
rH4PswSX2P54YDB1rVnCVWsSyG1PB1VH01X87eDmMTyRqMJoqZOz12dDI3AfWjR3
UOJ67J0pDQMzpJ7uzl6rfkN0GmOKbl+mQW2PTaVM0hhsOXZ7f5wIR2wFQUQ1K+5W
DoZ5zeaVEVgK4x0FXp6SU1+260dr093fabutANb6HuRDEQNwCG7ggF9ygig26vuz
AkOclGKaV3en34lKkw9UnpjVRYGXvWLYo0XKW4HVTAc98Kbv3UKHF06u4jn/skvf
BlZmZNip6X04lX2PF23PYHEhc2icwlE+n6cbQXqnG8arlFF9NcuJPXAC5/u751oL
OBBw3ZmUSpArEOCNMNfke8aSKuRfz4q8Cj+9+O0fFJnPLQ+zpcr0KVwOVNvTacLX
OQN0QyoFkDiFmGrxN7HA+Q4VfeNvqzcv6SD6m2COhbWAHVC8A9HWBSe5NdCiYk5B
SG4QiDb0ElhY/ZQfZjrDzxYxBBrmfT04lkbs+pXQQJRs2vm0zHDi4KzxuzgeQOlH
hqDK+7mJx4UpcXhSiz3eSQv46zYOpB7t5tIZL2FhkCm6UiA7jwVtRaXaIlmmg5Yf
MWKsfux1X94M8ZNXOd5YTXOfEC3GSfjLxNdYRLGProWXlRLl7z3x5xPH6noMy416
LEsNGGoa1NbJ8BpFVXXTi37Lz1eu0awoAB1xEDuesLkGTc5iDuzFPQOGD1iXKA2b
aHk+NIuZdGglM2hnguymMpkDJHGW0I8NLzHVevTmCdLmJLGYwLWU7s7FGeF2kT2d
/DR1xtOGaK1seyjWimaJweT3q2Z7tbaWuKGTuSjqjpPDPlKWOo1TJtcggbgkrKDL
yxIrw1EhuagbXs3IJiu55BAMmtQgpesv3pdvGrL0hL+uoRo/WuUyqMCmoiQB55wr
QqQLpwwZ3bjNV7JjtOHuxDz6E/fwNfcW+UAP9+3rWxfx9lEyzPSPZKlbhx75kJex
6u6+m2nPMRKPX89WHI/lE37V+Bf6SngqRKe0wGubajLBxKiVA++XLT1brC9jPe4E
7nUPzAZ3oG0KirwJkHDSvQH3WyeLd6aK6HQz44U1GolE/U88SranLUStyTJlgGwG
6XCWR7BGy26uhSDgVaRxxHXDSYFveXN//6XCsdspHezAY3N3x0PRx2H7LWdHYLKP
aU5ar7timgy4uR7fpJnTVrWkSfEdUM4JDo1JzqP6c4xAJ4E4Z6jACRsvXVba4sGN
COcybjW4Ir+IsZ9yMf7wIJ+UQYFc+rCLzrqHoan/b3ARUonJrfY07xxP9qeLyLQS
vZqdyfQPTOax05QiNwXH2cljxsUg6anxxT02a6DZokwnQa8MSHugF+TT28iVY0cA
UnWOhzjUBMsCbwP/hEOT+X21aIQRI+7ZdFsAiGMvm/wW+JT3k7XkqIhJd9ED4KWR
Yff0OKJpCLlAxg7EfGNqm3D4aTleKWTr8cI4h2jG23EkfDRTl7HU1FHMuTzUwyrF
s9JqlcHUOmfojMJUsO5Ilz6MZkBnBmyrDEB6+VjvB7OaCAcNXbtnVKuB6xs78pJT
jo7P58x0QtAbsHOa06fF2qiUg9mIt3u0/a+PTNX2LzbjekKoWWhvPIs9HqKYKOCV
PozyJZcySZCN+KPtuRSpzUZFLR0lkFTGd3Q3FImzdRCHXOp3Q4+XsCaIY/CD1K22
Ah0u5ZAm4LWkxqZeHULhjBp8RgqzBrf0pWaMUIi/H76C4st8Q2GbK8QA0vDDsQHe
amMYZahFI6xnSKiOJXbKs5OcQjR/MXfwXrnvh28iCMDcqKDi8M5gV+sY4vC/9vXu
S75E7nuEJLsQwxAI1cGHhrhvKvg3uw6y5j9UEA4fOh7GaOzJXU0Hl6jfU1q/eyX0
41OmFHEVNlNpjsGCsoMOzYsSjQi4iBjle+YosgGcDvnq46ocGXMCACrwSvcb4QwN
DCGrPz+1JGYf12jbNXdpbPfZ5g9tP31Tpdn5PVs0EtM/62pWciomv8HE6uvrM1eO
I9eCCDf9aDQKgY0UKi90a8HpfRhFejgmymi3f2xCtJ24iqKPVyZOrdOnVvOEZFGZ
p8JH4hUHd3DFttWY1soo7Cy4Kv9M2HV646BsohSEqB/tKiPWRyvIH8EFOjYWGgXE
DkZh+gdRR0AQcXe2QoD5NT/6gyPSYpP9s3McKQL/BJNw9e0aHqr02J6ZCtBYsMxF
eScbKaGHqfbPxFo46FocRz9d4gTuz3LDcjMva2an8Fe+sObPUe/hmLhHNU+zkjYV
4nlHaG2TgDkn44xS7DW0+mgsLsts6i+Kl71wqH7eiM8+c/Io6mFidkkIMi901JxL
ElSlhM16DO7AFBZ1mfM6Pi4zOBtPdr6nr2yyLSxUX1tfm5CtjtER3TLz24Ni5xm3
+dVN3juudp8A4IiDkjuTozceQJUrrXyiAaLHK5+aq1dKO/RPrJ14jthE2pWuYcpR
5OM+eX8byE8jPBPLOO5mhzA2PfOlSq/8tB2aZQ997eOJkCXi7Vt/QtlMSb/MWnzA
2Dgf8HFQAeOqA/avzIz9koLP9eAlKrNLNz/6L2lfV4rJdYW90v2Z6LyUWKn0o0+t
vjnR86PjFjvsQRfWDLpEtxjETmYAYYe101wIWE26bycYsbsyvCNOT19xjCTBc2m2
Am5xIM4ROtnLCIsL4++q6aXnS65bZ1AzOcsQSOw8ZmN4zJO+HuUFthhZ3KG9xQX3
UfyoMLT7VTgct917lgfpWjpr3RdrNkNtPHAyiVnY6CmYjQBKPjt7T48CqJ8Qc/2c
+X+8Z+V8+xVpjqO8vTvJM1QqWwLMRv3XWKqMxqeelQB2ggemrUMR4qQOny8qfHuN
u278ZYsdIZs1TQ38591OGt/5CAEk6rvEEQhhCkQpPFDRxoJqUx1Wi+6ReG5bi47m
i+njAmUGCWlGyGYkJglS2ezCTFHO4Ui8wGJLj0l1s3s+IK2v0Djfu/qMuj6EsVtw
Nb+gEYWezCb57M/69yAMO2kd63h3nYnIt1Xi0tJulh4O+tI5t3vOFsa4nBO1hq+g
cEuJ+OTGQ894wY1OzqebgkWS5/iXehv3W868fcGgpc8HKPXgcCJDYkkdfWNfp/Op
6pyMsJ0LPhAstgJT7pyfqQKdo/2fCxk+HLMV52WGvkAqvhfpvqE3/Z3hcFQXw45r
NgPbaC6OvsBDh6b5twi7eANBSFzaJxWkXiaZBD3T9yAPD3kvPmMjbeo1I0GL9Rxk
ARmqJPjsj2phhYrhY28p3fFT9VndxED5K/YkM1m7Zyk8AsZtlj4uBWNbELOejaG8
KCiCaVlXkbN157CPMl8LvNslcVRh4Ius0B+ryH1QXcxMRQ9Cb7TWB/k+mBdK+UlP
If6haMyRLuw8UdeAORmey8PvJUqY3Xv2C/VkNHVQFp6lq4E6l36gf8utc3D5lEel
SVoQUguAIzUpXkx85XznMwSEtfB2Az5BAVYW6u/ajznvALJVDha6C6vA/RvzDH72
/aSqTm7eoVjnkD1tJjr+H5TWrvnMXbN4RosupU719OrQwfsQErKEL1UZQ/U8kEtf
yACiu1NEW0qmUEMWc4fqhEWbiWoXPsfHXm9aafFOWFSotNWIVpspM3fNjOT8DiV8
UsGhHdM/EU890scEgMd+Th/Fb679obi88FfRLkOzBCx+2ov6hGcPELv8bQW2asFy
QidbWORWTm40xa53umSLp2l8qh+GnXW/UoFLfHrLm7Ydj8svEtaJRp+cwRkpGY6i
p+GhpY8ZB6WnEZy/oOkthh9BZ3wXjzAMpOjgSMXtzSZINK7JzgVDXR2TgtRy2KAS
6SC2fdqim7D59QL8oWfrfdPEUgEOWmmFBvkd4HbfJ4eLbGhhL21E+MNWOOv50i/6
J5Vb/yY31SV/zCv451QAhQi+9M9eQK3T38PFliQj0FN+HqupQEnT4zgzJjs0Zph7
SAKJlUa7YEO8vVBfJ9vBiUcWtWteZzc1QxjMGT4/OuAfmQ0y8lWnQ6e6KMhoCIoF
vMk8IqV9qlD6S1L3yR3saJrgO83hZwxCju7KFl3EgjcwgGPRsHdD1KjZF3Cjz8h9
2IN5xS9aSxgmfY35jB66Uo3DI6o8c6HHZa3AMpuKL4FGA8IwaQcHp7sXNSP42VJq
tFbhskrhIMfB7B7ldQ/UqdOJVh/DNoE06INWXelVJYlyLbq4NCFKJCtnNHzGThlI
q+BOe7MjsGvRfzZts8uskLWrHo+DfaK88cWMeqs6TZ+03RiSRKARn1ufOtGZB39I
GWgHfFdNDwwJvujiWqi2r+mQoiHsQDrnhQZc/fMKuV8iRD2plojkl0KEhgrv4Hns
I5ZTXnWPfIfnY+TeAtvUVPCWvD2nxYitHUCuesp3zHG0lA9LtE/UDhbYD2wRosqK
kaRovUMb/L1Gm6at/2d5zLEyKc0LD9TvBZnGxElfTd5C2TrHcjelnKlUz0333AJ9
qOTHmxkZxQbBqDY072uIQ2k5K8wqzLMGpeQ5lf5tjRYCldWwYfDwy64z0kNENaXe
ludGHpEoleuyB3JgUBQMPqtUwLQHq68D4zX1EDsff3dPPF5XKPEkD856HmO22jnF
CBYVSjw3Uu6qhapCm0LqgRQ/qejZOpWmz6RYuQaBAwZ7pTkbi/LEup8NmEuymIRC
DorFdVHktLynx95OS63vgE13NNrZQJXaUVTZaPZnwOvyybg9TwJB2xgMf8TJVJu2
n1HhedgfHINt0HuSgkvh2DW0ekBHcgt0WrV530SVkRyD9C9UmHmoRnagPeopGwl2
ocT3SFT390xj1BNDGLTuROKOytqE2timn2wrG/aS+XcgG+ajpY45i+pHsXZLAMoa
tQqju2F7RJrmfSSXHiDvesbVbVrh+hlMnGcE0Nh5pX/ycXwKar2ufaCg+YiSrGvK
pfOS5LxxCqzq8GPc0tQ3wcNkwEEsKQtbRzULoeonxvzkq1h0DWhor/3Jipnw48Zy
sCz5k2n2X3kNEGmTLgbUfUFc1tQr8CQaEMosPN4ee5yTb7RNCPtuahOBCp/8QwIK
5D0csw2pJUNCgLeDEtLeoR5nPGZve0BNiAEkbtXuiTWmsV/ov6ORC8G0hWrX6GT6
aiXl9w5oPfRk5ucaS6aaxVgcEj2Ll6Evp9TyCbU8pAkISYqonuBCZ9e9XljfJ0Zu
LXawOPus/f46ukJlo/KWuSblMPOzFeTx8rcrmKrb0oKABFTVf50bZgp4sCM8Vu96
66czgl50rpbn3lJj5Vt2cwqbfrQoXr7sVInLee9+RubLPUCTyI+HIR2GMIFXfarz
mL0GA0F1gZS9IHhBWSfDaB9/xHTdmK4bqGVzf0YsZOfWpB9K4Ryd7eBXtzg8xdDV
7EBIYE1JKLammh8IxG+KznjIYp5K/pKrQ4+JXS6bYnWiARVV0Nksyv5sQ1x4DDt+
8EzE77oKhsAO+sHH41NWKIZVswqWdAJ7KXB6mUjAsExRv2FjbqXd5vHFNOG6XfaO
lnItDrMp2TwMP9RQWNM7hOtifYCAZFa4Of7OXBiAnVOmqJRNHZPUvedMQYQFDxKE
5t4/JVX9EBHJvaA/m//ilI43lLoillOGmtwQo5ozu9tWADdoMtWmuM7IHLPpnM9k
aL5VZAM3ygdxQhZa+MMKWOdeDFAP0Pm3OK2xfkdD9xbwwaiwnsi4T6YsfqOKITv/
m9nzz+NYec6G2gDC2dno9Q8rr+PTDjzD9QAAhmUp+krURxXRC9qzuRRnkzFC1FVP
3PFRS/RxP7+hG8o9Bz2xHC3p+vHxWlKiYbKghyqkK6dWTDT0njohJxnlEcD00xHv
oEaOZTtePuY6ZO41ZVEL4qaVnnWlmaMLBJoyjMGQpQ04+aP6uHV6E+MFz9/knqFd
8Z0HGivCSrWfjTOtKWt223g1RtAdNG4M85ySBH4o+QTpa6tlzFopvx9yxNx1/SUJ
HEvZdRXrHhP+YeNB3QJWrqUfMKO5ZBUDJLFN21qsLfH7ZV90C5H5y8RaTvh7wvwB
yA0O67xclYKwnpuwB252OanfhojoqT962OzI//E+3F/bDvp8qdr9hfuTt2ZWWFrf
J8C0g7qqZUt45p2C4ihgsNrno6mNO7Pu2quR0mxYyXZ2iKn77HldF+lXCI7iKn7Q
5s880Y1u4uTcWNSWmBsovvj1GryO+jvAb8vdTArlSIPz4i4ZhyZZemo+a8TVpmrc
h2CotcaSF71jX665tYOkuuyvIrXI1MKA9a056Vv94zPZj8/gFCfclcqgE12g//47
0F08I37xPZylC2JlUNtT836z6O6HVeP9ScUiZe/8rGcRhYB5gqOCRdcGEkNE9p86
oJ3hjWzRP4wIy8ZEwHo5IZav18WT/NFIVf2WynA/Q7YyHTicLWS2f18fqCuGWNhz
UjZOuap5viGXgdkfRsObt9H0VVM8Oph4qms7keQwG+1q4sz9WJA9YrTcGGHmyj4O
ijjjFTkR73FSwu/6hmrJ6G4mUgY8oru9y+Q91GxkqaBuhDHmSQrUQs0f7Q/5YsIK
saDJsC/qQPEIdI8AFLvCQdDCagiZjeMLFlxLRZxfJEynzTJt8lDkxsjsG6YaCk+N
bdUSRDULNOcn3Y6vUvrMiD58uQe0nQ91BsKco0pDEFyPS927bz+/nqKUiPE9yCdb
ajnF2wjZpQybqhZubs/ysm3KAwzJS28gAiYSyvh83qrX+17RgCZTeAcw0VtrrJWv
y6lMTWkw3qK5bHGcE6GR3Fk/Tdk8mnboxuVUxRbzyaU+FKritPdxAthovWhmiIwb
rzLn5ITcvC+fwsipk81p9UZUGukCSWzGtFtJCJ66UKb48zlWpKY+Ue8cM/jil49n
50IJHI0JoTcw6Qqemt4lNFd4TvKZ+u2YRIfU9kEULj0YIkDIohP+E3edDNcYkJ5I
UXDKOag1miTlo9ojH5hd2bUlKN2YLxqIhl30hz/vTQQLsSx5skdfkJASVTZpJZqa
GFD8Rh6KR+i5fOP9I1alX+XMPCc/6gQXMBBw5DZFGQsAygSkNPIE2XxH4jtc711l
5dCC21jhCoKD0pdOPgE6YvQjHqKibgAjvVv9CHzNJJTKm2EyzU5jy7iN3Nd+b+ry
tkNKeToVw6GydQ2jUhJ7uCUqToqZYwPcuqhqBWIuWVuwYIHJRmQubhWrNlhcOV3j
vnaqxeed9sR8VS7dmR0W0vyZQwJdN8UHFoBoqVujALzatCsCbZK1AnrIPRubOkck
umpjeRnqfvdx8gOibZ63dnL9x1Sid+R+fZu+YucrFvL+TscO3IyedecqRG88THZv
gud+KhT8KaiqorARQZwkwubC6FxAy3oYvpLNv4V+ocDArkCNgYX4Dqen4glwTAhJ
AI0LKxVRHYzGpDAjMg6SrK/CoEF4IxQ6Ft5RWaHpXdnJFc+BpeuqW0/2kKwg9DTS
0YfY+ruznDTK7Tu3Eg1hzlvePrjDSxLKYcAMju4O6qrTjxn1g95uNvsl+hJlxj7y
ETZS56wVyie/pFp+ScvUgmVMg1ITuovKuRSms4SXjOs6lO9D2+JfXz0RfVEf4QZt
mK7d1REYv44fObwRLqEJXkSYVc+QBY/OjjQ24ZzlMmyIhL1rUxNpjCrcbF9VDozp
sQymKRKSArIFl4IbGSEtjAW/2z9Lej2KKD10A6hMMKgNVRH5H6LX8/73uq32A7Q6
Axl/xDH/hKSCSK9ULhl4vDcWKzcC3tvSudX8wyCgcp1OH3AJzgUqCab9PYXBio0j
DfcXXdtClsc+n+hJFd3U+CgG0MjSM5LSOkD25iD3vOhcQabQBB3JonA+uJ2Ujpn6
3d/M3uCO6eQ5dhTW9/4n9a5XPE0O6rWViGym7Gl/NCmyp7HvociBLGMRGVEfCm7Z
h5DNDBGSu/+G53X4IfauAQ/9/QSdbrTYKdoRZjC0HZOmgUSNyfr1/DWbexyHc+E6
HnpV/y/Uz4IdEGqTbAWYVE3lJXlrha3Bu8n1oFTFGImYxR+HKJ/RSk2RKM9xjmnq
CdSTV4tnj64RrXbsv607G6Ei+Ytq29MIrYBoYEjsDnqXw5I+QTTgwD/Y5fP1sCgo
UcWkFGNyARuWsHsUR2USiE0TyoQJsTBwrUfWrOdFzKz7LhTOgsNHWhGi38BOEYfe
e4TiRWJ2sGS8z63MMOHdeU+uK5dNaKKd9NTwwCNu1DnvPFv9xpOGueB8QZBdJ+UA
gjdXqeqCcoNYuPH/VA7qJjzWxa8bvlIQPDI0XYpE1echph1nI83oGMlWCyR1+7ib
wPpLvcI7yaVCFsR/cbMle8AuILYEeR7n6G0m9pvBdlML8YSIxSD5luZOrTWyPVSo
T3vM6dRdiSKe6gopDPAGM7BNIOEVLY88nLHuy0DbMpwY6XHb6ADg8/lOWBsEXo1p
IwFjrR8tSaCMn3B3QIziO5Eph3AtJaySnt4ukpgDaxIqSZuvOqIL6nmMf6sC8d6l
BQWao2SW82GP6SNO0iSjipjdBldEKrDmipx6yGRVsSbIU/kBjNmR0rjmymBYMXJn
1UBzzrH1agg9ZacRDkJZYwEkpd+6ZvjOMegQVlasENzq/w7xxLAk7LM8MjhVsnfy
GSaBLK2FpKCjcgb9YffMBHCB3Wiz+B9RbOGVNN7mWbnx2BHYk/p2m2FAEGiaaqvN
GhpfMgyl/LCeTHQZvdXqCLNG1URIGghKxoQqfHZWD3Ad6aIIMZ5bRlxMB4pXcciv
kbYYf9jkLmPKHcu4VJgZdaAlAx/6Q9UQJlXagPAY+JWkMAx1Alax2PJeqJ4h5XQ0
18lKB+QEMvnjb8ffrfs6ex2gJlEEuZR33RhUI9+LOHoRzU6NGP32YvHau7FNK7kP
JL//6QD0Ztce86YdRFEUdX++gJci922UUx3hap0TXLFgeeIq913SBla0MNFvLGrg
bRwJSL2vtNzZ1M7ntBtFNZogzkkdne3+/1Dh3MPFYrtZ2Q9S/RuO5j5aKvc8HaDq
AoW7xy8WhfKVMORg3el8D0fGcJSNx68SbGwu7BwzurfmGfQV+8ZAdjMpjDRtRTjL
Co+Nlsfa8iUgdUkCHoYBCnw62D3GHTlqNtaFzvJI1k1kyZfqDnQmMsZdYwObMHbc
PZX68Nt5Gyb1Hz/QpsxgjDb0g18jJmPI5rhY9dJnsvWQFArzK7jvMQ55J8cQzx00
rfCnOUBQBtpcp04dvN009pjGtqBEB03YdqfUeSIb6wEOrEGvVZLl0xygznqpBrYm
Je7NXPbnvLJ1+AQFXrmx466DNb7uz27St5rBpaO3NlLLu9/PqSxYII/hMb7jsc4V
DnBoA87Dbxr4oce0cUZfa1L7gZ8Rqi+kJi59qg7jGySpt1Lp1JNhHefPeZRvAa9n
QckE7goRboWvMpH/YXgaxoSO4f8RJxeeBR2TMQCk6tYG6h2LqnpyvQyCfNQRuMdd
MS7i9UA/XAoVAGV3OuqnHyPK0Mg+qnDEbCLy10GKskdYgsNkaIOot8hSmUA0PlIr
T9B5GTs+KAnCYZcEmTNU6R4nV8TbN65Wy5VfRq59eX4TPblSjaL3RCx+gTWPKRH7
KqBzjAWsBej2Ry9ymPaXTGWvcoTxYL/0Ah5L6YZUECX6Ko8Xb8AVhfdtUByUj4CK
eQUM3bZj5qBdI7qhrn6tr7k+fYepUqfvEQfA2ZYFO0ep2BIJUL4VKohSLx7S2Jtt
1K4rUc7keFQjADJNwVQwynKVOoIvoH01D4ncSXq/nxxt0GP3NWwDpRC+AtucfaPp
pWJLSLOZPF7nlo714unC+BTuERunlsfVdFhU0u6nyzIj1P8hcTUYkACMQBjZXtXV
fdx5hshdvfXnMA/8UMkKpaQywJhHHHBCbSqgF6+ju/3j91WNMOPrIvd0IxHSTjKX
+HgqSmRNrNEZK8Nx4JY65s6M1Dx9CFKLmEhdM/FR6xH5a/1KCREZ3H9wjxE554zP
5UWiC9MpzcB1ZeO6Y4UqpFq5HHNb3vjkKIy/7MiEHzTC1Q9qQuji615LBk7UzEzR
TzTLW6M7hvfsov8aiHJcfabuBVEvhBozP6FI/Y6lAuNqnsvKlqa29jdl0QySd27Q
aVpug3oVO2pBwjdARagqOaHV96g48FBULDxf6FK4WcrsebmMac3vUKij6uDyPrfM
wsXi18GBYfR3Soz15PCy+00V8PJRPX7PlJFLSf7qn78o1kOoI2H0Nbx6s7lY0Xxm
nQUUqL3Wx0K94fktz5l0clBei6ZSSUMp27fhFPVQVHjqAVRXOygnFmLWGp352Xsh
KDNylwg8RAL+IWC0JRgDk/TrZISpSDzij9Fr5LP3xdYX1AGgKRb/lnaNrtBcEbgb
ItJO7HM8OCcCfHqlrWVaBIBQUGJxFkty0yBpTPJSV6mSTR1G4uk3y/EN434IPjLZ
PuFyYJGeAj8eEl4DcOPptYB+ukn7KSuLI4vc1BY5EV/8p+p7aiIL9U66XudWXLQz
6FMh8ASjs9I9GG/8D6jFr9egQYDd7LJkYTTKPMnOv8IQ8QDGEjwjgkSQMYdPJx9E
0pqMETmMRArOPbB59hcr/yqfz40njWywGVVwIU9d3yNVySaB+NUzP+N1394Q+4th
Y6HdD+ZsrKB2oza8YapBwtvL8aQbpYyDV0AB4Bswcz12Yh+faTHNml+yvlX5yS20
YaLtjsXdhcXZQfM+ahEn8MKjvHlWmW+yob6UTll2ImWyxR4YEu4WeBMM+sgQz6L3
ozOI+//KnChURIAW0/oqo0d9QyWcrf8tVd442D4Nz52r/dpHBqlE62MYw6hPgiwC
EusKjAHvhhQHkvL2KkQEiQhmvujkiTntW/EVT19bm/Se7/7VGVz6gqz+z6m5uglK
SADaLW867416aIv4WfUq/Ji0pZxod7XUYm02rhAdZfpf5ohvTP/Y54MjVYX+KNla
R2MP5qGCNsyMC10j1qhqTgmdWiM9g1+JBCltbyqLUkUDHK1wCji6XrzfKtHkl6FC
O1zGU+4WirBauo5S0Eps/1crkT34+yjU1lWl1LEy+V6i5hSwUq5EUtWbNZJZDC17
BvWsHqzZU8Xm3DfKPV7VYuDdta5yKgX3Nur+JKBjUNe+klcI2YhfwYnOs1udbv5O
gQkF995jmp0DTqc545O9VYqCzt2Wcgbu0pryDu9sOlgJL6ePlelQEUbbsTnTigNS
7gUlGnMO1W58DAuOUrD5EdxbpAJ4meAsWrEqgl6btiYpoFXNQhTOEDTl+nqty3dx
0h6CgZnNE2kn2iWe+gmqUkVJM5IH7O9+NColse/rTCJ7zNNkq8OMVxz2kjgK1gak
sXhfi5SBMy7Qf87y1vZUsShERSLBd8jJgkd64GKefF1UZ2ifZHWGjIHS4AL03UPB
0T5cvLNybb0ftTiBV3tEUnuHYEyHbT21QTkZuAi3PimDbPQL821j1YUOEi7/mNZK
1L2nqjAMRbPWuz22k5RF/IAMFbFmXJ48b2lYn4uIBOBTDs308y1TDRh173Tje7z8
7ivZoXwrPX/lD62JGC/txFCWjM69q9osthEhFib57qdRAwa1L2wJTVMGdMujfWAS
r+SKRr0a5RJAlDEjPz+RaqJkOKD+gEfbJh8lz1lJW0tVGMQsy1I1+0uBEfqSN6qc
mAoCDZ4AvlMArhgPZGYge2GX+lcg31Rn487imqy5ljAPhHt/yU3NWnHRQPSg2por
4W67Qfsq0ShOxoBf+5rerq6qkxuYc9ShzPUpkJ0TkWPBCkCx0Bh8o4M09HiXzoVn
ldRZVUKWiONFzYX4C805OQJbFNLGUwCsoNvEX+PAuX5dlT5r6QdGs7x3HkPjWVwW
cWbpowyTPT0ri/UOba+iXxc6XvmwH392kHxzX367P9ZpJetz+bztk/i0QoNQiRu2
4x4prMs2NtRgj5u+FhKispq2wfwYOr/WUc/1vwZ8Uh640SL7Ql4HrJSFqb3eM1u0
2XmANlRATsKrMvXTZeRZ25dD3oRyuTLnuNq+JEUXV+GwsO+owam8psPEfCQ1Uibs
OKYLYBMxkancQU8uZzO8CVlZNBwMWgxm+uMKNte8WP4fAC1GPuvTRB+Sjsvnemly
1oweq6wzu526SO7lVt8vUmFHXiXoza0P6dIkjlAjCFVuWguou3083G/Dzd/OgItd
cW6r0J2nwyQ5fBuk7v1HdsCeYKv7LWNPO9Y9UHg9f8AKJEzbop6LC/jP+nXoLFmy
ba9iK7T95HceL0zEL4SkOdeV/kAOi8oRHvmfH85MQVL4uZUISgfglOsQ7dcwJbcw
qhKtEPSAMuiwvTxu8DZH4MSelfJ7F1DIAkUlKUBs9p0igZ4oUly4qKzpAUQrSXj6
ATCi7YSH5iWZQws0skdd1uc6cj8DRx1n6d9RJLAMppFIWj4xVOfYaZAwq4kwe0/b
1zfgphiIn03Z7ibwSBuuHYT+NdOQzPQXuCHeB6zzlAHX2xKzCkOGvDdNPzI6w6Jh
5ln8gZVXfcRLCihRzxkng+eh+mSlZ2FLXCv5hXXhJs4GB8uZ1YErZv61ZKaO9g/G
umrfsfJ8NL7fSaY1VLq3Y7QCQMEZXoyGNaNnnxwPwzgEqWBM2MzsxskvvSCA4n4H
0E89mXN6Bdq1AGGgWVUiFWYtkd7iqr9/JZB7aDQFh59rGCogEJ1tR6Q3v+dRpozk
F+ixXkvfvyojuY8KmWBnEOBTsf8wbqBrMujP7rlVDYx61aE9Swjtli5G13oGEV1I
XRdJCZYumIT565OlXceBlq4ZboO/9zM4ctuWUAgOsIVAUo7I+5hwC9Td5fJmzBjp
nECKECFV0WbVCSQZsaJ5kzdHVPL570MSCBqArC/jQ+KBWBCpht2WQoxiNV3QcSLK
DjDqrcCrin1BuAWwGla76qP/C0r2Lk7jGkeNpn83ITHbvASzKEYsuA42byutoORi
GONHg8BdoFrygVge052s27hszfXvMf2uPsuwJxxnl3WDO0aDopdbCQw+ihVzpkd3
gvt7SWc4zrRvT3vst1EuikMtthwdDmXt5LIgfql+l2jGzRq6CPKzRpSoktvAKFDb
P9QHbGMnZjtHwZ/a2qil87JjV2uCg9AgzEkWmXyYyQ+wwE56GduZpfQBxT/xyjYU
vnM0yzAtlv5+4Ws1maBGjn88ZVvQOBAHHzEbBu75Cp9x6CRRdKdDFh+bRhepqhJl
jUH/0m/E+oF/qjhi61tWAw1Xt2MX9NwDKWnMYs/gh9auU8lmf6upf3Ybd9A/9OZz
CMsqML0kaG1YtKbVapME45cVqTTM+gSQF/8M1nxw0L95ekLy3GCLubwss7sJNBup
hob7KWOQ9FmZlFZw0JLutnMSi331udsq+H8RxZLnwvnstF01dqBRIU/Q6D+8MmSG
r/adTWTX8915JwfzNgEyOLsglil7DVvxzJ6Fu5vc6OIa82jEMTMHKahCadhr81FV
iMjXyV+d3owBW71oD+c4RpZ08oMTEyp+tYr1Z+xcHFsZv16k68KYoIP+5xdyOKa2
LAz4Mrh3Zye47CvWskufLRYvyaK15eWW4HoDatdPfrAgER//gzO+uI14/dfbPryN
xxkQrCrcO0yBtFoq63I0+9lX/uTfPXTFzdBs2Q+iu82wR/uib9dmveJsfifwxgNe
I/7HNw1Y/KkNIKajMJVL56up0oqnzeqZdfr0ql8aVOvSDLSgkMnPaP1Gom2Ok6go
FiXTYSp2lX21/5YGeUx2IPMFQvzw8jffuHFYVU0QET/LqKiBovk8tMvFx635A0fu
T1dIEmcnXL/Emta49I4z/Wmbns95gyCIh48vW/3rOpX0NNKhYZmndYKORwIYe9XW
p0A2v19fm89QiRT9RmxN0z3LxoVNeMSbFLkSlIZYCokPnP1Sx8+qv21vFA/CWop1
rIS4xWnyqH2Yx3O3T7R/tiLrXptDE3a8/VbnBW2OXms+o0ZQCb1uzyPxabgg+suK
fRPF55NHQCjEocPc6fyU9cntlAmfF0WJ0d22m/stirykMcLMa2JE4kpSlDKer62k
y8sF+QBPnEIR6uSAkjcRlvlVvHbTm/MjrR4YRFoPobzGlkDp3zIr/8LQde2p4sIt
ZGpOZM9Jrib0/B8xduWoKTLs02NxUjng9FejTQVY23PXWSo1tXI3nRB8z1APUU1S
1hja6B0DtY+N4DtRPurFI93VJLH0jNa+whmuwKIJwEAyKg2pmNSE+/PS7KRYakYX
`protect end_protected