`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 45040 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
N+AbGUvfDpEoMIf7wLov5TPATxW2RnKa9WNv1bhpcKqpVKNluQ2Ll83g53BUE8ek
VfH8SUiKewYI6R2zv51K3gGo5b60FtFxIBJf9u5OFTeNMU2is9mYbc5oqGzZcYM3
/yJ/KtHRTe+NT3eJZS9z02TC9ddFO1ikukW3fiNiXP0uQRb/rjYoAMuKj4lBM0Ec
to+bXCjRMQCA7isQJ3/Krkvhi71X6ajpnYnuKyyrmpNUKN5FVNhRdpJ1pI+7c0zt
qJ0r3w8yhSAeDRGVVNd9MmHyYD/nBzTBGYXCV6B6uFQL6+RH8H6C2KnI5cPTvCH6
HNsGdQAIQec9lM4BXVf9lpZP/cK4ApuhnTYpd/c0Q1SKn55D+/84Kga4FUW3xFui
a2tA+UX1WoBqqk4SEyjJ/2RNmj8MtBGEYJO5z1AFuJDPuDD0j2cWA5546wz5uFja
wFmYmw3M6cwwBw/6lbM2mQimzKV1g81DaqnmFnnJW4wTDzeH3Iv54g0RvbBIm1Oo
x7Vsa6BsnAqgNZV+XAgzN7dh+mtb2+JWgNfNpSNUgY9w7pGK73NOq9jqGAcUVykZ
8rJU6EetA+IJsF3AqSMcO7lFvPFp/jG+DK87858Lq+qIwU43ZQBYtw3vxhae8BnW
d1eHigvFcbHMTctQkHvLORSjfszJGWbdQlSa5R3vLSHW3u3xhjL6Y0FUclbKXbRw
Q3mrHYZ9wgKr1wWWxmQ1R/hDAvkG2YKkqNBI42yEmchz/SJGtERH/gh568SBvT0H
vLt25aPcyh9njrzIG78VBd0qAKHSJRMRumXnuKgLcyllmC9EgEcmj8q9Zfh5961D
eovkrtf+CXVlA593O/ARCbeEvWHda541rVdYrvTU/7ywskZtDsjOGJQop2JF/74M
EGDKfKQ0jMWD6CkMkyQmW4ZvvaDmMPadRdpVNX6Ey8s24syPa46QIJUCcnUYTRw7
MEew0iFbajDP6rw5WiLM1xA9J3wnhKKlV2shPdMYSptjjg2nuWu91BCKYkN18ykK
2Wr3TvOKbma74BT0gPt5yTaC9ZN0PMar5Lm7V0aO8+SSbL7iSOhCrVjp75HZpbtp
V5SNs79p3L946y1hTFONmdPp7vitnTn4FLEtYBHLGNS8YGqCMENQAdC9iREXgISd
dZI153WmNCxvxZw/O3f56qc0ECSjDgFrzR5hIqySbW0NHcaFxIN0xm4amBGPUKRx
lCU0niXdvx8VjJdg0veh4OV8jRTfKoROlYtlep61kdcxOqPNAsEt4ZpO8pXLRt6q
bsX3g42ONPklK/uxwFzJ0fNcPaOELWlYgBpw0zbEn5KZfmo7q1c/XjSGnpB90VoS
TY5yqGIUpp0B4m7n7gBWDpzcY/7TccjuCwVLGptr35n3NzCMdcA8Ok5q2zLj5xzn
8+54fU0zoUkKQWtsovHOvSVacUPjMTwN096HJK7P8ZN6qobNmPHwWaEo6IEHLHwh
wzjc+m0nmRLKKluS41A3E7u0kA+3b/1uyA7hUbH1pFVRZWh6Tij/tz4FqQKmh3u2
7y3s2yj2dWJUSGwTnqfMSnjd2Lir9KjIN1AzsYD7seuWxrL9q/PJpNPWu7lxJKW7
rCrcSKRb4XBVXsZ0SubVT22ZLea8RYBTA3/KZpUdyRWo7AXHpRSOHuGxL6nQKy6k
TUHbkQF0sLeTRKrEgY1IF+URbspkPGHAbJ0gyg3kPkW+ZDXq/R4T4ibJ/yWQwgqu
WskkmFRCA2l9rdJaam23VzN+hpYp6u1EuNVTgAWZBqoMj0StpIx2UEodko4J79te
4pVDsMjupIqgn+ksDtA4haAylTnQEfYwqlEMi7xMeMrnveJkc6w7Kp29vjPx6IVg
3QdTOsGElig8oUKyW6Ztj7y3PfZ97vK6cLS91Hgs+M4V3zOx0bIX3xTWHJxujtme
PgHuM8zbMgT2GVmchP8//R5S7R6Lq8Wu6lhWuOh8V7UT8bYEaB35t7b5dEAj8dAK
ZfyoyxCpH+eiP26JSw9zx04CMSrT70sCBEx2EjZXL9+EFUrfgBTt182CKSBFrjZC
PiXSCpz8+jaGba9Df1/yUokTU7uwLgQnupKfp/jeU0TA1DJj2tIzk3oShd+Z/PMy
4NjQIsbeAFEtW8pCg/z/nYtn9eOr/5rfy6WgE2k8ykVAqsho0tdSnn1Vul31E6/t
XBCWTVi+UV17brJXwdwfzWardolBo94egWaHDitUiPYduqWUoJAbIRPKkaKf2JVE
IEV8iqJc9vjIsoKvgRM2XcdBOYcZlKnQIzsk/J+20mrkY/a78VRloVwu/KrmSekh
Q/9e7vsd44omsqzF0FaoeEkvSsEqkh679mszZVNezJTW/dwaoM38Bs/SOtbPfY2s
Ad8luLl6TVZqp0e+C/kWHY91E6945fB5z8rgxDf5fHvL/1IFK9iE3h4Zi7xVswFy
jV14z7zH9QJJEp2A/st6TULVdUFx64+LLE9fi+b8vO37GWrQrEtGWw3mRUg2wtPa
F7JqLPL/dNRGS/lE7kqmuDEwet5LdT4wBDFOwTJuuTvNGSxMMgmzMw0lR2PF8TTd
funNKqdBwCrnIK5DxMCHSTMsdLkI7l75dBQbddndJvL23hDv1WFaYiKiT0OHlLxL
SE4j5uxOGTQ9SK3aewQZiL2ruRh/d58o07f3eOEntnA5t7iZ6I7aQPO5kTlfqz+L
3O0dNVR1wpex56+lBvETGgFBTj3zalG9RWnokTbQpCs8FstV1lMYXwtbIuwdNeag
3NMuqTrr2JkF7uyZRRfP7Z3VtQPfirZUuAj6S5J5Bb56xMdbDj1Tu9rhst8ul+97
Z0LFoHa3DG1uSSEoEYnsCMnmqtuTUwuWldTH5y3NJ4H3M+/696jNARlwo8L7c5x8
2D3B6t9R83VxFq2MsixDe2jZfwiSeBKKGr1Jm3dnmTg7HDPZjpFLFPDp3sI8hIXA
FDkInTmiLGGl8qZPANGHZ9msxoydXnO+0g9ZbsQQsHcUnBm3gWsGFvqR0auDWnRt
exWHMAeLU13hjxoPa6OBKLsADL4zXkx6xGLQBbM2U5o3hvUCQoNe6M882nkjjOoz
Tvv8iOddfAzpV7FWhcPiwYOwJXIzor75n2zR2tW+JyXQLu+HcYngmEaksl1/ejJc
GBFu7HBQ2BOSXmRz+xkh+IV3ycbgdNmZQyWT85pxV5Nbs+rlwuCFQHo0FX/cDY2u
xJdrkXjpdR1J3faayEhvfRRhJVQiEdzrBynY8YJ6QYa9Dz0adQ5syfAE0TM5m2Og
G0ODMzw4VsL5Op0kbtnSf/jDlftcimDXr4wsa8MZPKrmN/RVpOPvHpHywBDjabl7
90WZb/TrEjE7cgAj1abGKYqPEks3qRHjBT+g3cF5hkniuQvR2wiTLhav0VDvPTQK
nZkghA/EN8VFJJnbFvgZ4672jV/d8PkRs4JBl+z5M/H5RYi3+tfjZ/OVH1llP1Fp
XkTr2ID5P5+6Ya61ooMPsYPdDBESGvMVh8YXCSpBXgR8WbpuLYWX764QfA7yRWQU
PSm9liGXXjPMYrVY3H1hdcvMfwsuNGAtJtfJIqgZ0/ifTnMZxFtzKyeeDvSUKEyN
zdpMnJ3SnonkwCueoV6BwEKDD4lnf3nFbgnKdXVvNqN23NJ58nnEycnsLoRYikEa
vUK1e0N9QBALx3MlDw6pDi8AWP/Wqch0qtFQ5t/iNtSKVVodiuXsqS7G3rmRfoIC
14/lj9Nj8vZAX/dqXSzXsvxb/ndSnc8l737hpOZ3xlVRgO95kaON17o9baR32SKq
xEIpwk8RNfD4FUQdNNiOq8d9GxbmtckXrehJg0mj4/+nkJWxWu3lq5pBjn8MR5PM
CFrwuOGudFsVAFjoJqKRHGX/TITU/0sg41Futm/YrBjQU4Ps3aFwHFJJWm+Z2jVH
wdoCLlBK7LziFUQ7y/zv8GoUdBVjjZygikPCnI3Y9p5nypzuyzc7zjUGXBOf77dU
oD2l7XA3n0ocbmBwK/uukAlO408q0MxEom940ZhOaqYpxHcru6W67zI7yqrXFOWV
B/NP9x8rzgzfuUs7IQwloR+ipvxlQ2s9DcvZPmr+sbPzJZ85b2HxozAXqXf2uQLH
Odxqd7K3eWU1hKQKgFLGtlZ4qWz3XFYLpxfoiKDZM3T/OkG1EM9aAkeGyhMrjaX9
dwqgWEDQLo6p1N4Fk0vkUUyw/5i3t/6mwpeuzCYRt7LmxXHsW5ZvmAr1DL6YRzmy
jd7vjYS12FiyU4wh1o1s9IIexXeNT5JrQKmiuj8H41cNn444gHJV65k0ixCT2sZw
hCb/1105qpb3Iug5yjKVGpp6JkEmfMnKcqkOV7Lq5yOXT5GffuW3Y4pXOdWpW+G0
sgQO9hRWM21+BGQRQieb3YvdbvuwONbl0nfW3nMOWEoMVe8EieHC7bZM2HabG4Dp
9bHDJocO31FJtJW/1nF3d0ICwZlhzVHPW22iBrJ8RS1Z8QL8fCR1+r0IRv/qc2uO
asGmfLpptnruigwVf2/0i4cndgNYEB9tXP6j/zgt5B9aFyCayTDg3LGU/fD+DVJr
kUM5VDBQdQy7bOiV5Kbt3vw2HlrXDutxKgN9xLbeBsRsZXnZ+iAFT98RMCL0QCAY
zzglfg2LuCOC31+uzNUScc79GvyGtGlOX3FLSpgbfO76jm9z8POyWHKUc2ub9tEH
AG04ixYQqC7Crqr29hvWLc0q6ozLAB9/5jy0lJ+/p/EauwN/jZhrzCFSiRV/Lg3O
H3sEqcIo8idP0rd1yPd8CqTCBvuIkbtGdIUg14OytrWvIQvExm0YrVm5qgXeedne
/dxU0UgzHcyXcorOLMtKogZO42xxKvj4APL6xw7rZEja4+XUdghB7FHvXK/s3fe2
AuMpnISEvk+uXERQKE45PS/OIV8DDY8nOSlzoUDEY0705HKAzZypGyDykKw1eV+B
dOs3vQ4mZs+Dzf15mWoCI0B2zf8vC3nngeMtI5vfw+7awHj5rcwek1Lr1Ht+hOkY
JxwsMqxBGIC6HKjnMztAGcOyilZ2BZtW9fnDzOUcRgUPpzbX6e3pE18keW+/CroK
SIZxe+UdbXwlTtDY9Xkf+rhOXrFQXM1lt+09WTKN9mzIG/6LFsYacXwf7zjN144w
elXN8Qi7ZKnlqe1J8nsD2Y5wEC4WW/uGNFBwG9pBZleFAG5Ycn3nDe+H/Kvj0rgB
iA6ZSnJHhMrWLLAci29pXh6OjFGsSsJmOFAC3dyXD5Ebvfg9ZoqMjtsZgmtOD6Rz
T4TvXWa71L/fuj/EIJDFzwqKimeyVzLh2ah42d5V5pzphboYIE18zmbcFAVyju59
iLY7CGIG3yoHdaIXhkc+TfTwbSI24u27XVEAwjqnv3lIVWX1YswRlUOCC5VlcE8/
nGeaUNNHwE7R019t4VAPg8LuTmXcMCpA3lPjA3YkyGavVANIRa6XyJPl2mbz98df
nSRbtf5PxcObVZLuwCmwY+YjLVjpiZXXfrH1lQ47cj6PJBA4wnABYQbngIbnj0Zw
LIDvikVGDkUGD1u9JP+CavoyY6Sby1cEN+YEHDqNhz9K++5wQg2sipOFVyI+6VkX
5wOT6LNkBaCcs4WJxdQjA3Jlk2i4ret3tNmBfE+cmm9zUBXJjKzUj8vRxYcUO6gI
5gz6nUGo64x4ajyE74Gh6nnJVmj7BxZzrkmenRUs6z6rgpV4m8jtp0TASjeqyvvB
hKNH/9gQQ/rXRcTPuBaN/opG7Tc6OVzdL8DNt6/XjhNM5HcYmiIRU9kwoPbgzDS9
vOO1lhyIJIO6lHahlsQoTxfaq02Dq9w+PKXSEn5cEr3sbEMJfwxGnD9mykMkA0vh
2Mb+kIVrzjfy8dSzB1IawB3ME1Wu0iy8tYafsbkJ2KbEVvhmq1c+CZ5EwrkJ/q56
fzUzvuA42uzpIsy0JTO9uSJ3WMFrytJ5RnxyGcf8dM0XhiU96w7Dy0DrnNdJmBSU
Xyl8D9mSMasULXgfJRloqmSCYXkGI2vwnkUahECvKpDBysRN3BC0fCz/F/nv4fFs
YC6moBkHSFLx+LTXvlh9WA9MVuOM7BGdrCx1cDHqmZf/w/SepQQWGbopULvQebyM
aroQYgl3qVuUxVihDmYXe5if1ibxX0fop8tFmo9JvcckBVqDD1f3U2DSIMmIKN/K
qcUKoGAHTjsiHlmkjmsAyy9MbsrmCS/cYcf4nZfVz/TNiyGv2dD4/5kEMwvQNd16
+ORvb85bxTYQa4P+NjsMqGuU6FKEfMKG1D/EaZDgci4XBMBRYlyJZ9K/jXroBLjr
RCgpq5QB4t5VDBq4o1cLfAurS//Zi1sb0n/9Oz8gQIMwmasg54Ou3FskeGxzPSHZ
Gn+eOCa6uzkWWKcFtV85pAoZzLD0M+h3XKlpYxvJMP5prf3uAmYWZWuE4eYjVwS4
K6N+nf4hvyegKunU0Kk0jWVtK0qZPMSdP1DDVHTXblRhWm05pwjIXkU0mmu6ugGo
a8cWju5nolmA+sBV+VfXdX5NW8x/XT561SQtdw+2Ipt9Yow0/rVg1dEE490Kq6O+
EyS0Xmmsbfslqn4pEfMSUFTrMvA6NqMyrEQE+YeFs0qRsp7PNdABS8ShrdT7SJQo
l6f5+5U1NvS5PccDViJi7r2ddj4TIJLHvKAK3LlV9/X0DoodhSL+3KRvEmjEqGw9
Z2lHWub1a+9VelD6Fp52u0O3CA7wz0DgSvEuMOfmThQAEmKQP4evltHlO17C92TE
T9+34nL2sLcGn9TejK9+TmJoRdB5qoJkdNmIO48MdqIXUWgPLKE5DZ8sFkeR4FGD
zbN3EvfDCVKWX+s94yAQ/5ugndwY7aVx/r6tgJIm6TjWR0N2L8yQMzqvQ3DSLsgb
p180Rb3UUUWxns4KnA4vN020yXQIwK3pwL7CFee7UsDENGmZVUUP/G3XyvY/sFBz
njw/eBGd15r6G3Ypa5bCyPXJVeyl9xE3WQEeGXINUaMjqhhxM6U5PTP7sro6WtMM
ARS5RtEsZJQItzrFEwu93t9hNYFaZ0rDsfHS8JW24+BJAKnLSX1ryWuNJ0dcgDip
mOFEiGcLPfZIDLGzvVCKSd613PtO9iWXBbGHGZd4zOdlLEwgU/OtTpmH0mo75+mc
zlryuwKcAZbOa1vd0LzLe5j6GmclfTleMzZ92B5NJ6KuwBIoAYeI7faeyp7SzNEx
ER+V92EvDsMkdbIOAXLgfDjm5DrYL+aP0RgqXsbtwf/k4KTdf0wdW1XYsFWOvWt5
yUmj9JrbDMTDsQVFKfen1OONO63G9KgH6J3M4FQLXn3OFHE3/t1LxgvLP7CQnwh+
utNNNe2QybJzvZ2get5OyeKMJ1ORQsD7WH9QsYa2Wn3TB0hAqhxzhvWci+5w7m34
LdPQbXmjK/bHmdf6Ne3rJShoTp8COCOEzNGodfiOA0uu1lwz9CcdrxLN1di/Yhe5
LBg2ZpiUGwMP4jStTv0qq6APPvM7Q5LLIiGzXEnm1OrXb5baGirBzIZdAp2gBCNY
zk1GsRiirhqRArH7dZNskniuHVmjCebythSAO00UXxHEFoTnNt+Gb8o85ehjthqI
nls0l+tjqSSWlkb1TuoKWLz6XYd2JgW1TO589d1U0MztnzNg5fghTX5DZUBv6Mkw
UV7PsxcRzuxPiuMxV8M7pE2d9qzXIzLFVIgUx4rBnstWXZ1SF3QfLeh4FlMYOm1y
xFjsBoSW++X2EIXf93P1ahrabEK3Jnk1L7gRJiL34lkczU9eN/hZet7muVBSkp1H
dqS1/gyawbl+U9s8iHmpe71Gfb08pLwKQT566b9qsZqlbdUBXrnwqt2cJfbeh05x
zGxAFqfgqrM2EwT0vWHTfngPAG02Hy1mU+wOoRqAejE38wEpvdTWUhN9jR40b/Wr
dAK4Bs4AVLraLVTdVDtOYVP/MMEH1UJYkGFyBoYgyvppoXfMZxP07FvItWS7AebA
tAL0N8J4mCwjnUUs05uYwM7NsOZlBIEU/ftDKtqCpbiWFvG4ne/t+2agI6KHZrjV
7ymmAwMBiTBWWgZJou3eJAcaMN+G9q+O15GGBB776Xk76ToG94twiN0m9zdpAyvx
S9jHqC8csGN1slTQYAXq/y0EFuc0n+TZq9JnymQYXHkRi4bE4hBSfnH9iGTCfcSl
poyb09JY2mVkX7OKif1ivEboE5CTGtaK95uFU3TB+mi1wAMX2E3TnuVAYXSB7u4W
kuO8iQGG6gUqYozboi4hp+PD9TTexo+UgKg7RIIBrPn7N9oJDZe06LlN+Hx0dLHM
Q6trZJHpD4EoRjAVicYP8uyzXzbqQm9u7TA4uCp/zsp0529ivWcS9vI4aJAI6eyo
nfWJhH0WMh2m5RTIboRh6SZkUmRIZ9TW4X5SKRourDGCur3Po8MRHUxkYFifempp
/2xgIiG5DYO8IhM718mYe7+TOgFa6N8Yn/PfEazuQZqMlb/BEws0vklH4accW4kb
LvpJjH996rKLieGLpVZ/cZddBe9NHichr009EeYKmx1j3bfPROZDPs9UfzJvZvd3
eHNY9693SzRR7DG6lLfpdD2iYh0J54zngJAKTiSb6eT7pYwWk0UQ60KFqTmox2HJ
KrFsupAC4WgHwQ5zsYoASwZuLiSscrrNUgQ1qs8Q2KX75v3Ey7sUtvPYnJFG+FWq
NM70X+aeoLRY3uwod1y7BcejNTFIj/036xqgZP7PxO+TCOxx7tq6BXJBdTPlKUJ2
9LmwDUIwYT2wt6C4duZm9Sq1+VQ3Ph9IWZD08GJUpHSfTavMAQL2aXNKdSdzpEKf
wpFCVMCXFtEi06pHgMlLs49Y715vWfiDbBTCPJc6H8HzueCYY1Ds0Y7qGdTl+F0k
1HbfOzZE00PNlv2pwOf0fz0CpeQTCdHSDJzrgtxUO4ioqCz6+cAXDi9UpKiHz12D
8WVF9po6U0nvAnz4K0qs+VPshlXjER8z+B+39yG2mDgcPdV4zvvGlL+ONsETHLPC
N8hoJMaTC2gtrsOlNcBZLjU3seNXIPVhOj0yZc/u3WJqxH4koP4Tm0bKes/R7ov5
sgjJx2LMO9aJloqqYMQQFhS6MWi/8xeO7iZnfZsdhfbnml3OuJ0KclhDl0QwBDuH
svpcx+1yUwB28iFOkwM5Vd7LRJMigN9RQSavf183NKqSKXsyUNSPG9fHp9AOMWf2
OwcjkKf8HqnFGtlS+gmuAaL1UUKZ/Cv+QhU6sCw4krhX4ZMqCfG8eT7AyU2XK4QK
b+TfF3axhxrw1hzMlbRD2EbhDeTlG4RyHaNLH0bdOSpywGYzNOq3v+Ehj3maKEz+
I32zzjKJQxYzaR7Rfzb43W9k03IlEY0WtYWGVfmXE5FUSHw/tTdSD7CnEL3BpiwX
pb3bvNFjDrrLz3RtZ/NDfP2kQyrtQJSliIB+Ch68bpztI/k1MJHQ7LvVyk9ETpI+
LLnf6tI4JzcDlFApIPPfH1Jdvk70vjZ6XrCXhUyw08iFmnkP/pwqA7MWPzPd57n3
31/0Og/dEsoHoOHRULgV66Dv37p5WgSQJEZ/fkAcFArP+EZcWX80lIYKJ3VLDQsL
PjIwEgYWQ84KgdXznkf0PP/DFcfCd4IWEVAVUvy9frtlWt03ZJ9oUL5ylaK5NcaX
fXtqmT66EZvJpQUXkRToSDO52wpqoXQQOHmgd1Z0XzsJdvPW1eJEwTe9jrEdlfi4
grhbdivG8DlXoHPwBBKLgTBR99Y7Z7BLftp3uKZRBIpjDAMtRt0KdyJ94IUzQNXq
DbDxCwUbQssAch/k+RlOoZI4+vbE67+Kw9pOIe9UqFqBiG+CNUoSUY0e7xLTFg8F
0g33P+v9sD0/BT8ED9jl7s9C+nYd86T9ruYwR2C3BYB6+27/W+BeUQUT07WOGCms
1wrgouJArxZcl/wyyqVv9WVgMevrJLeZ2/QM/i5zI8T3ksICfiVhX+vBr8rNlFOA
7hCwoZgvmify+Pvw7pn/O6fckvnOJRRm5MbzZzkwe7+/gwK97aBE5cUqWlcWKc3/
VAWvzwT6czMSUnxWNG21K6BqcE6B4+5v0xkqw425dsrRb2G3vLbr5mrf78Aropcx
fVqfSEDGQWvMWEPplVz+d++ERNC6kTPGTcXbk+9aMpCKYbzWrtnGEI0JAmnD8PBl
2ZPHIzP+gDRdCokFkDk8g0z/pD1ATlUeSntX7VUD6ZtFlIxGBhamVN9BVNAxzkJT
R2mmvoz7CTZ3Wq7LzGvYA9RswORJ7bryNXo6LtT9U/XJDp3hb4d6HlSrfBlTRGZw
PexI/XCx5B5mYyo84DLUNZpLYNSUpf2+DaeNqJQgsWoEixKp+Q7eJzqwaELHZFk1
l3mrNQSrNTtYlTwMkYcRV/Z0asZQ3f1IU2NHwkquxkB14umh+2zvHn/zjxJ9hwSE
mMTN5kxtT9Y5U/R7mgUuuDc2C+GwRC6whVvHMoxtlDLQylDTa7aENFUqMdGDukBC
m2/93U2pVFmDsGonSmGdW8ULhLiJuMxA5LHpDQPLGAcHt2q6ymWts3Mjg2Rmtssi
bTWdgrQFF9+ChxqrjgObOMx4ffg55elukK6KAmJH8DPc5z4x8Ux4ame7Weuh9X2j
HTcWyGQJS40kfSycq2PhvrXqVfMUHZO8/eRoL7pNX2Xem7g0x5yQgeEmr714+Te+
1zJdmvEK+ZSUHt6zJq8nQqfZfwg+VkcA872YK+Ert/AD+UKwKdzTJawad3rncO6e
1B7YW/DogOp/ENrGt+38UBn+nDlaAdBFjI4qaVSwDLHSFlMX/oM6UJhmo5AvOP1d
loUQP14i82kA2gl+Ku0hTW6FMFemCUxQMeuZ0XTVW6gLUp+GkknRoweOAHXGHdut
OFqNhQ5wG7ZLDpzcToirhvZhaqf4XxK2R1w96qRIS9DYDInqjg7ldfqXEJTKcDdM
DgdTVX7FsRPtglOGBBEsRjmIKakAdV2+T27vKajKRB2CwltO57LJPceMUCPliJ/U
s2wrqxO5OIn/gqb1W5aFDhXoFREhXWC6ubOzURj4AN9juQesFGbKlA227aikSJ48
PvRmYbn6HuxROHFiboC63iQRpr7rTjL8PJ3PikVT0814ZLrZ4TK011uvTq+/1RdB
dTk778ScVF7L3dacSpkpwoL9DY9GxKe64frENRvoLDNGF8RTDS3zvXC/Ab/HhcTQ
r/a0Y1ZZ8GLBrt/8imfmhdzEKfOKYBWik5dyLBPXgIZxkC7KEsWNnBlSOvzcuYhR
YAiJxGnCAFwOF383jR2Jpbe7jeHrWFSqf9T584PPpo7/37IJeRug6zoZm7bS08k9
t0rTIeTq4ECdfQeisfyvUOXUk/OdrSz4Ywwd2Br/xw4+HDc9gRi7XgjP/ryfGzqd
mRg95LToh8hjzGQm0iTTjQVs1+yuvTAZ/C13fDTFk/q+zH3VUGNr1F9u3TNWKsjk
XbNPioLfLye7QZdINI2hx90nKvu+V+Fr07Fe3Zsn38QyjyX6clxAB9c7JcPTFOxl
WMyJAMq9sSu9eR63M+0k0o/fzYcANjGr5qWnlAzGJMWouf1/Sj6gZZWwg1YdzXjH
te4TZdUrmyDn7ErxmijGB2poFvA66ikK6N4iAxIWfbbJHXLjIJ81a4bWZ5NiP8b9
+Fk3yTtBCTdIH61Y0ZFF722EsF8/5xzFZVN7P+hKubXQ+05AMXQ2l3bU/8mB5P6q
YEItZ/FDBWw+1sVWsEyXcu8WUAbK1DuZEDRtR68liIGMmZn2xuYR0nYixLIVCUgb
lWtVhTdKEy0J8liLaDm3oOK8s1YRmcA8++zKakC2otxQDCfT+/unt/JE/kh8+ovw
Cs3htWHdlm9ElvnUtUJtlfDak/gl/bcpgKPN3AfSl0jZovRfwkRtwyd2lCnD7yTb
aKJh2l5j0mQmbWTPGEIOgsPCZV0FPLlWH8g+4wBsx0sI0n9oM+yxEtdKKfhpeoME
xLMsOSLkWpsHFRRtYDP9UB/SWXP088pDfqlL0WRMyNdq2mM7oSPCNYZmcmWUywlM
4oDU052mihZiqepozaoZctZjI6IVVto8m2+7wezz2POCNBRYpRSAop9caI4XCPmz
CSkzkAHzeJ/bY7DtS82Ai7OywbiqFwzNbbMD8uyfy1OgaX1HiuFOAl4fAKIqNWdF
pmBmtkUV9d8VtgcDfHbXMnkkjcIWsGLekTYRbozpc7ncraTbS2eAnpdyEwdjmPEl
Zb+B1FF3x2VixNwrU0IkAuRrK0u2lFNJJfFyJRdq0aYR8qMsAY/z/8VQ7oU9nPZm
gDYcQl9o/mgt9wntWFtarQdRhluVwhAEwKhu5ydQlvrjLUXKlzq/gOTSskh1wd1z
y8jyfI/QrhPN1q4+g0mh/lJfhPFz38DPjlowLlmd+aXoomJMplnq5q6MyqyRqUIC
nAP0HC0h27sQxQOjxrZv0dtR0REPY80wC8F1G9k8Th2zIFcy+mPcRprafurpbm1A
yolsqxHMMMqm6YoSltIZaaBW898XN0Oh7Gq1bcJKVHo4DDRX67YKmyqyDiGircwE
ZPw8pZ5oOM3BfTSHhnu0PDKZW3X7M9uvJH3iUVQwsbDRgvqq620+kzB1HSJt25jz
Lj8hPFRXMeZ+Gj0ZDgFKADcyyL1sl+nZNOW5sgKhqK5t9uNYBYetAfJCFvTGLLHW
4sBJzyGTiXarzof1GGAdKGxHnnl8LffuWp4dEeDp/yN7+2ktr0YVbDshDPYvA+Co
21boBVig2p2uMZbinGkNfUe1S1Jnzp+EFjyAdmcvOsgNJOkXIajfAMxhu1OIPE6d
GCZJMbVRmJDJ6/lZNIIc2NPq+ekJHROwmTadVlJddkILWKBsK8/Gx8zdakrY/IHS
oWw8eqTEkrHU2hio6SdsH/4cCBcqX30Js0kKNvQWAiDUstii3PxL/gdZauqvz+lq
nYhYd1pTS4gpUr3/xQJNwszSlqDxrIiI9Rn/kz2ovKOLCtzhrB7Q0Lphpg7Rn8ta
U3S4LiJxAHjC3S3jWicoliVS2wlIf5ryDR4AcM+cd+J7xqstHkg4ZqskrYlTBSMO
m1bgDLaJ8fyX5sPany+MOHTfynFvFePvdPCd/ZmNKJCigMEiMr49JyUQvth6x6zE
yb8UuuFXGbGlRXYZBpmV6W+/14IOsC8tLGWB0zrvdKeOQRw+76/FVFs8DCpHfvwy
NFfLqf2uwg8WTfwmVoRihJ3uhUWfOFrx7H+3jUaeF53M9lFYmv6fiYEZmFEeCuJB
Wyw/0zyJ5YfT0JTlxQZERizW0A7EJ2LYTfz7IaesW7xvMNBh/TxbzJptsYiPYaD6
M81Iuq5L/ci8Rp43lHN7LU0yP8jxa2i/oqdOqm3WviWRnytw5QwJRtcauQ1FghU4
zyp8lHSozNIy8b2QPGrA2SGx9qwmU6i0PfWdNPpNvV39b/+XdFncPzcnTXwZCCaL
Ou6lmMZM7xZehVJEdH1kEZxqdbzfy4ET+8w7ucJ5P4riYs7n5fVtuQrwZEj4apXH
wtVVAPMQdwbPK7dwQFuC6ykTkKxTw5dFXEgQN8dzu8rYM5gb3JKN1EonnUXmcJ06
Q3Yva934HjUIlrLeM2FxITqpXiVG7LGvEnl+QL/upWn6kCRaXJ71p07xHctNaFzN
WdVjbRjRJcew7UQA7adFsnLphjRftCM1wLe7nYTrlu+C9Kj4K54kYsSnAzgESf80
BqTsEu8stceBFzZiCJMS7CQ30xJUtbsviOTVyvw7LlaEXCxKYttMqerlJLSIq2z9
Q2rEryDyCuvvjVK0hSlmEViGi4Zy1yefYdZRiEfR1YHBuEW9wXkgfN8KGn4WVQyv
kqGT3b4Fd1SgZalMWEh4pmptiJW9PBrr3BZ+T+2wiQwuuuELb4yagGtowkGiPzRq
VOzBeHYoKjZIQ+jRZ4UgODIs1NFOeEWo+0ylRE/mDHNB2gBPQVwy+OA7ctRZTD9z
TBA+gztjTur527ZRBw+FyvhcteJVnfENAihb3LHKMAwsXsUDabzyM8JtQtUhX8VA
y7/DrkcEOhwq3+/VZk1/QfAWl1D/qtuBdUbXQoM8NaQFZGHndk6jH4CQ7rpdgpHt
HCXys93TEjEzDz4Mi6QYsizkZZMg7DD6O0u57PmczwErIcE31TFMGBqoPct7GkY4
blisCAQoYdG2zKyGyMnkKIo2sT2eM1eMguLdxq7TJ+4ThX7d4bCmpSeO7Ij3xq6n
JJfz7/yrmW6YRMuqYvUw43IP75FRkO80AKr6WLNdLp41Y8asP2DG7XC5O5eCretd
iajDrP6JjWGI3J0Og+QIt9+a9jGgTHdXYWoscIIAn+SiiEYEiS0oymsmoyJ9zLkZ
ySr8iPH3QGORxFAWIrcaI4RHDZpRss6JfFAiSsnTXRfGLJbT1dJGNPYzZwO0XEFu
vBkX0egD2+KH2IfLhp6M3MLM8pkJarPjZUmJ0Ee5zI0YRk7xihqHf4EV+9nslt4a
43oqyEGTp1K6nmoPfe2zkLvsE3RYSUe3w4v5SNYinfgEDZmAJAxdG5ITyrbHkBLn
8bxkBtPQIPT1H9YQHhAbtOTdEYquac0lYsRLMOzG+rTfhWHtEnhTEuznFquCcE8l
mf62TkL8+a0AO1BS7AK3H6Q7hsASOBEHXNO8PU/1oCDqQC0Ca4voUVXffxOJCwlp
H8j+qCpuvQF7MJkPhUF9doKnxQM7pjSJ+KCfYjTLC719wBttPe0fzy7qjs3DRxDM
jscLWRxS92ZgkoXK3MsyNRgfGbiPYvNtYd8zegQWvBFpfFMDrgLHcIlpMIBRk1mX
60h3EEl5PvxsYcRKB35OJSyqcInitz9rkkorT6Iz8sW2pBeixDVzTkHpVbCfBuTO
LHluWk7w6S7N7BEwu92IJp9jTFlfkgzbMq9CIuQcbWuOJ1BzMtxdZMUQBgAF2F6M
mI6W0jQWO0tR1YZQFrHJpKbBHCAzcgGnseNtUQIh1Ngn/yCYrOGDWl8s3D5dVnvJ
nckGH2g8DJfbGTsS+Ax6psviqFjORuXcAD00iy/PqhuZxmGRy8OPrv5neZS8OG7I
O7OtZpw/yxHDSQ2uG1BEZd6Mv4SRBICkMxVf1Wa+W+SsslL/2bR0+h4NKgUw9OUC
6DuGbWrP2171T+7CNQKKwwJrB3cORj86eDoEjhzY+QPuqzmqkvz49zWymvP6Sd4X
dktUCW3lLVoanIRoH4Zdp+fVZUtWn7Ihs5+ZQMXdDqzomjBBKJPT7vKmosLsw2Vk
/8Ihs/b3xWLBEzMxPXKNDNb4gwcEuDoC68ewDeifb2prbpJTfkg2k3dHxpwj4m+U
SzOCMYFs3cdMXkZ6nYVikW11xl6svGpiFff3yocb4OTn8RnTpe5k94Mru+EANjjS
iORGo1NwVKJvMpr9U9b/w0apICRpmEhX4vdKVeLF8vTl/hDm3/CAuzmSTl9arcmT
9QCSuduN9yXEYnIL2ZdDRoK33uq2Em8G98vhccd+jzjBUqXdArLDggZeiqEntrxz
r4F2Zd/7S6e6u7LSnjVXkuzpEOGSGYwIF2uTmcLL4ALXCXcbhWgsCJSlRe9SM2bE
44/2atoAP6+RwSKGxN6XGn+GmbZk0VizFJgndNpH2NaG8iLL5/tkBFZEZnm1AR7N
zMbv0K1HqSDYPLvYeHEBRF3m56V00LxqFb/Jn+4HkdP8TqJMe3p9RadnKhQNR42K
mmvwJ3SFyjJOu4ou7bacK255AZZptKVjp2AZbByEIudh4X0PIxSKiwyYesjaIG7R
dwoPzTlQHTHpqFMYaGv+Z/cEj0I/tnuwMeT4Y739F6K07XqOKerbWVgIwzs9JpeC
3JFtTtGU4EB+XQUQSeZKfWeS+DvVeVUI0MaIrWZjUhQwjdKA5bEwo3eam83fYRRu
sHt4BkKrztVDiDfsyzAitPXj83Opo5JeAnmu4dMaefq1FnQ2CKiAwDEbeByLSpva
nl0etY7OkqupbroJsnygTlD94P/IQv/DWHGHYJBPDsg/EqGd/o6+/Fcs3P86Vb2S
cpP5PFjw4FE4BK1p8lu3NyvKcfr9Uvq3Lqi3Bh+43S29AzMyPhcrWgZp6UyqRAU4
KpDEVBX4PvPl1S7tAf5us+i1NXfD9TvsKeahQdkHdU5n2g3tQv7WjNrBHCW/LIFx
tzzQBoBOYnKRR+v+hLZkjMsjNKXyJ8EP0bZ/yQHNISfDRceNRQ/t5Aataf5rnxkr
6xpLWHM2PiOnGc64y22FNNxNDcYJEmnGLMZzbkF66zz1+pnZc2VWftWwzuBk3rMA
RBGhbBoMeFf2n3BVFElRweabqUpylJiWhhnaPBBIK3YGJRhrr+Fj3xOwAVInA+mQ
MyslpiQV8IVFj+PvgPop0VwdYS9FXkfbGuU750ZgUz7cMhR7Qdj3Pum+te2qAUFq
tCiFFcf37DflcYdiwFz2o55VJGJMursho/oyXccSmgOdjPeBceYr0kQ5I9W4FRnW
aG9Ls3sEjXZb72kByUEiUyU3xSF2QuvOgYYCEhfYf/cVENH8klXa91gFnxn3u/Vd
REuK8Pjz0rL8QV2umoO1DqenKnDhQgctDVlf3XbqzMfdcgZA1oRzTBXyASSrTv5Q
AoeyGFBrQKZpMG6EUTri1FFuxoll2HjjsDMgLyGsueCgY4vWRa/1Lqvjl28FZF9t
lRtF7T/nfSwHw78xKI0pjrqdMfRg93ACEaOSvIkKZnRAVBZMcAHTDhNlsdemnBzO
BIbdnOh1NXGfSrPj6YXW9gL3FQYpPbdjDWSnYROu5tnNvSzDuKq6JOsR+EZBumAV
huvYfUgrd2oCkuFBSj99uqcL8pxty59oRT20fMUJjZ7QGspbe2MTgB8m7aPNshBs
CCSaE/kEcnO45UkexqZlvmv7GSgdnbNPnO7ax6MIYTG+daptkjzZB53OoHc5seYO
j++RrNoz3xQ12a4b763078Cz8iQxfzT5LSRAfispN9AckarK9teoWi3+bS0WH31F
eXliZp8KMy2fhn4yjSMepEji/LEmFKRsjRmsiXT85sduKCA+gOn/mlVvsPCsaVfp
WzjbwfaPm0aWr9FDAMlOL5UIEL3oJ8JR5JwqYtJueTB36FZqrJtlL9HudpbiZQjY
2IiKcUyBjeodhL7VKSNzmpVmqlrb4Qs7flw5ktdmwUHyUohjgZaxubo4bklEIHog
JiDHthwengNINKZw4FjMXQZ1dLdcFrfcDK9CdadPweOJeMPO9ZwlvY7K8zobFNqB
x+mQOyzSjERyPfkO4R7HRqr1SQ3wB/7tnrkM2ShVjY8EFkzsIQClW2PAHRZ1vQ5z
VKzq6VrL6lJS9buTaVzXOExiz6ufaoKgU5ygWmS6//G6oIMPi3Pe7PMeCfsmemac
BNDphvoR0jjSHQc05bV3ntTwzSABAXPsXvPUb7/5NX4jpgdRbvKrjakxZ40j/hSF
v/BGdj5yKYl1DP4eGJZgZ/Hcojtkd1uLALdIs7pcDwbKWcZkdgi8qhHDIK2O1OIm
jr9xyo25g6/CyyEaOXM39CfQyMWqHwvsKNju1lpbqFkUn0qypICWRaxTM9S+PRqI
uNmYYvQv131Ilxinyvs9akGscY9fUk2JOMO6kJRhxyp3uzW37C65Obi8lrIUJfrv
OUmtUgQ1pN4dN41kr+4XrwN5UxKocOpbkIBkL+iYHFjGtgPI8LRhf5Gq1zJan7jk
URSDAZL6pneBe4LmwH7/a2Y5N+gssSd4u8/4lzoPxMOAA2U1fVTy0NU2/svxkGFx
KWSlqrQzcxk2TMB8C+/KMDMBIbi3UYTpISkOvzRN3lgJ2oReg1DNrj7JxIdA9q62
4m/wfUk83XfJ6Kohdqe6tSqRH7AnmxpCbedi2jWLwUaCGyc8c28Xkuw4IHhpJrCu
D8G5HdSDKrfVs3z2NNdYNV7nC1it38eC5ubyLGwWmnWhKKVO0mLXF6eQuKlKtmGJ
PK1t3bHgGnwFBd3lG0gtcHEUij/di9/ra6YmESxaxR4i40d3S1wnArY+e3Zagi74
/Hh2lVNd4rmfReErkvbivPQOzbHsIQM2v27Tp9kr2mvYcpzNiLWqvmyOyANLAz5Q
qYSUjMf3wKK7KQgTUILxY97hVdRNrivmWr2N/5zNImMG0h9+aMTFtQ0SFM17Qr9Q
auxGwSuUGV2AJ5xzIuA0Y0XzVt29ZXye2kEncPe2ZIHWzOqXfY9tfLkCO8Re1Hlj
j9KzSP9F41JwMeKppWmE4mqSjh2++Lxi8EzimT2PFWlgK+Q3+mAvGJvhqrwrac6X
qO9us5e4HTcRcVniVOVnH1EBlrgUaGWOusLxxEZHTJA/M9OMNHtBm00HBRwAyibc
A4S1TZBnX4rIKWFK/lAOPrrq7xqOeGjn/tSl0lAEh4XrgzgVfHzHWd07G8qcspRL
EvitxIVJCvV7mS6FWWYr7WXAAc52KPhloEPwjSRC7/k4KdwQbzXO6LN9lG2JY5ig
S1GWDpZqrYqZWj3eHkx2zhaQ3atOdL288HY8E1PGRnMiu6A5XgzFRzlYcaDWd7tQ
iKVP/kL0x67iAFDD1DbuqCqbFt33TIcqMzwf4sHcsAHKlJCPExHFfj8oQVTTuMHG
Glm1EacW5DQFr39HJJcWi+5gxtI/RB4G/VfB3UeZ0DVIbwaYkRTjEgM9cmcuTG0+
QKv4O3Q/FhP1nXHluSsWSLwtcH1GuOKz/T3e6NVFfUC+wEW3iSNBhxmanEN1gxxC
8cbWj6dm3Bn9jvHyVvQhT1VVT0+O2lstVJ0LZPjvWQqM1NdL/9RsSF3CVp9Wlzz8
8Xnisq0d/Lyk7zunugQRS0nPO0ztK2UW3T47LrQlcrpwCV5B/bln+RyTQ3rXNWLT
NhZ/a2waZif25q8B3voUun7ji5qfzBq4sx29yo+zfjg9mjMewqLAIzbfaF6hUrKI
3/lHdVhtoEcm9jIPDws7pZ/Uj+M4eX7wfcrrAlXx+vubdaz68h3Wzwk3vlsJ78Jj
7eOB6vPUVeWIdrX594kyXDhvxRnE/9Z3H0yY46DvdpCg/J+XB0kjH1xbiR86qsK6
t4O221isCUD5PISc4gHMp2+LEPWZYStU40T3uDbpRh28QW4nx63QLpKjnKzOKK/c
BnkJMu1GN7lxKZZi+fC/J5GDAUEeI21If58pcsEzrG4cUK+YSuEjAKldJ8eSIN4F
PU9rZF/jLtuHgtkD90u296EETMR9QKCgJDGGsMkS9FQeDT/5Noe2Bt4Rq6OksMnq
kRBE9XZ5wTJryTFSdJOQtbFu58ZyfTlfY5py5nt4MiYMVTWPRkTO27MCkbGREw+A
8WNnIRugxMLhDoX2YATrApCRmTeSHS82sOkCn3DThPZ2KcloLwsI72VVbII1+V9U
C9OUqNhFr0eIeYbBqc4nbYd+jwyjjoY9oZC3tH/h6usUJaysoq6Lvn20oZ36uU6f
LoQBKz8eqoZu+qbV80hKuf07l/RT0QDmRjCUrPx2ApmYUtxvXENqB19VpnkjDU1i
/Co7qcfmoFe7D+OqyZ3VhrCseE+A5WxtAxhrLhIRxSEI9kWfMSLaNRnZgqa2Rp1Z
Q0YIbIPvjXK891zFkwUEzYnXvx7VltCeS7Dk2CSlJ1hwuR+QCXNnZlqWwOp8+B1x
ye1ZqHwiNrBqi35Lyn7c7lBZ2Nlc4VOlh/i1gdmXMAaXYjFgI82hZMKK17Y6FDuD
xlEHBkxZ9UnLDXO3EbTeZql/POa1sXNzTYgjdd5ED05LrbIXlRSkeK1K0gjLyqUk
hLdrYPlprLyLi4eN0hLQE8ZkfF1TqQ61x4FflY85E0dF67XcU6C3bm6iAcmgubBk
q2qf+imCuSKIh2fXauFG5T60RepZOdLSJxdPUhpuc1DQiPpA4dvf80i/yw+08efq
bYoItZPQxrv0nPWly5Cd8s+q1m0tPwc4wKw1uFvLwVNy9UGRN+jplVs5jSkiaIRF
QlI66em5Up9Fzwda0yXaIZU/+4f6Igk6c7D2IMkKkOeK4FZxrnOQeUmaCYc6VfdQ
0J9zyblYgTgeL95SlHuSNTwi6FyN3nDVf9bnwL2NdtF0Lke+kotKGQjYKnoDJ9GU
gTJ7zeFAaZ+DtYAvgGizD0Y3zqu3K3AzrUH6fNcvSV40B2SY9VCxmjvkKwho6tUO
aesI08CZUCk2MPrufi1Cn0agFc/k1kDk3VCy3AvOl6sJ2GUtXWYICH+9xQ6Y+zYZ
xsOQYHpCSwQddvW+HrmRxM3J2xgfbPc4Btewq1IBfEyi+30TcnrOgxLZMSFxfiJn
h7VJuI6xXJPpYwYSWsqT2FOioEDDEb1shV+yhjXIK/aav1gvFC1r7Smp2eux5U7E
2K3IUyv9iDBhOBdljK2HQJIez+E8bsqaMhLpDTI0WTkSYB/eeaLy2iC8ZAIVg/zi
WQYRp9akgnj1kWwQLqgZuKC2kQGusImONKGc4ZRhbbsnlD80yTKMk7SIltSbtU0N
fzk584e6nf8m0UEoFIrhZBckuB+FlF7jKfTMnUp6JYNhhYdZhvByaVzf7n9YWT60
Fg0Gk7U6+a/uTCJKMObIQtY4Blm46cxt/7LWzccMz1h7ROccyVqaaaZVLmlE1LKs
zVstJiv50hvJk2GwCkQtCz2hGyq7ka5u3zm6olc2OmmtVPb9yYksIPX5D3azRUxR
2+GgDRfe2pkcUMlfEBT5HuvrZ8tbHbHLdPs3BWhcEFZTUJRBd3YyRjMksW4hCYod
voE/8/aGxgMm3GguAceqDxab6n/Vn1c1UAcklMAHfgSman7wVoG09qOybOS7OVbC
dX6PxE37V/yESseRAcbcq9rnTCXkc1vVmUZ/QI7Yryo+ZHUlHMcoNVEKtBuiXlIR
cyMW9CvghVPH/chiPECD2tI70X2eRSh6A6Qn2Fj2lyuTLKq7zacsQkXmux1b1Vgw
C3m1TEMO9ohq0wHjC+Kzc8UBIv1unW+Yuix7p0oI1+KU27PYKa5a6yEA00Xkc7mw
Pg+XDAeYK8rvryz8ymz+MNqbLR4rxz9JsHK6qwieLjBKo8t5ojL2J89anlMjxuP6
I/1REMx7O/B1SSOOxHyQ9N5k7SKp5nzNAawIgc/LeRhDtI3QlRZcImA9Lc7fcw4E
92UVSyBTPifAjxo4l8HzTZ6+CaGTvd7vjyIsuauWFU1EHcNqxV+VgEHBEC/8zH0S
w/KvVRvl4EHy/WX7SBbpqi5yhy3tC5tcIT72gFlbF+KAaMm1R56P7vZHZXJeoGP7
tka/RnTnIrxeFdn66uNwTyta8GyFpF0IZYfgeCR2dgmZ3R7u68z7RPgYEfxKPlQ8
BqgfB/OXT3xvY+RUAFElqskq6kcAmQf0YJKmN75pblT/Re1slFrNnT7NRCUWtci+
gmBC92PuLlAVcXlTHs5oL7jP3L3CEgAfdxTN21K+M5dxHO7Sr4gkr43xHaX+WRAA
GQS12X0Ud/eIZRDQ5qk5BG/dpnQJLuCw8ErefNetnOwP0uFauXrp+k9SgeEtHvEw
BUR6Xe72TjBj4anVUlRlTHSFAIsUaHOmfOAORIwRBS7UgW5X2uXR+yLrJKL9wZgl
bhmu2O4Nu7IhUmHAH6WspjDvCSDrf15uNxDiJvh6TYVD72l9hBFgKCmblb068CdG
eKXuAb3HBmqlU0dnn5j6Etdf2zOrjtQnjnES26KXScBkKmDgKIZQXFr3pYcVQQfy
vh+7gWRwUGGf/Tn1rLbCH9TJkS51fcQPquoPSvJohqu6clSio15lB+BT8AMPY1ra
652OMr6bjwassJFU/j7wid1uPfQS4VWp4Kxz8OAsBk3Gtx7FFyAFXjzH8vTqv/K6
vyrmQiUrXtTOgdqcR3rzIzsilydFinGzKlo54pqMPpX+d7WZ8ISrbZwcNOhASRx0
pbCqCyhEpv0RB2ZjAb8rY9CvTwLxqVhSUnkPEILlJmuP1dW3PeiFzMrK+ZSpBAy2
vZrW4Rw1gEfDe3aypf9ddBtd/fMXHfDsSjRpUClIa6dTWhsa/lCYAlrOQC7NmdN7
BEYfxRTIDy8dNEBT6xrr15zRQ1V+OvQOSLHKr3VnDm3wOPiikciNbQ5nzG5+eTkq
eBv0gSNEFtoYwxHnaj6pHiXhLYNotC6VUAguCdt0lI7GpeOJyAsRcq9K6ouCDo9A
0ISbxfk8WF/Q7hi9o1gspSTHSMRAEVDdTSprPLIgRFWuLUErrp7w3K9b6WFQEe/3
MFZcKgfVipXq+H/jYP8FVPbWFxAW2Epg2mCO37ZbpYi3Wt5LiwhP4oXm0ZPjjxot
MX8IeZ0qcaunu8ZdV9/VQkkQzInXzHvgYzPKqHsl17MjQYocfcYqWiJtu3Exlijy
eKLdK8p/L7JWvzerj41w/XFir909LEPA1V88DFOZHJKQTJd3SvkTdr4tsxP3Wdeb
x1uqOm9oHiJfSM1gL4WjWpwI6Ij6zMoPCxY5kniJDDq64MDuXv28gWgMPwakhgD9
pDpKYR0l//y0V8rtAduDUtGzT/3sZJjHDp+9lmDBzvc33ybRP8mbO6giLoTaGybi
y/qlftUoPXdun3AaFva+ZG4izDD89S4vhwlSla8Q7T2PUaqtjaonfRf4GrmZnf08
6iMJo3J5s7qBGtcmI7WKt6jaU+QuCrq0bSaP3shX3iqvfdkN/lkwrBv3N7ciVrpV
ih4Vf8R18hSKv70NE8NlYuxKpcjHDWwPV3qpYmKMYFIFw1+z/JN9m9C5GpRwS0+A
erRObkqlvNbTspD6RPz8+xsTssTr5hHTD4BfdggrNT3bnFO7OutXkqY4k0mLmu5n
FK7mcPyzFpbEf2EquG9p1Yf48m5arQGNqr6EoKV8J132mYc/2kSv9JGzL9C41Tq6
CgyaVkT2wvm6gD69zqiVwWm7CYRsgAuWPetxYwKPCViUWxPGAHqjyND7U4jFOyGu
OZEhDUfFft889JA1blTZXvoWeHHkiYS2H6aFAG4tNWgfvRVVlVfuI1PrVrBfBXLB
LKR6SmfzDZGThzokxuPTRy/iX0tJgZR5uwsPG644uwoAJAr+AkK3gYj8lPdHI3HN
YSLTWq2R39nrFDR5a8q23Ag0Tb5C0juhTgdyvco5RLjIUU+b3wvjPQLj4WuQyAEv
ChA/M3HOsIFT187kzVS9Iwy6BI9WQzHiyG81mt6LZlo0dsYJAUBjUeidFWhJ42IZ
4Ui++f8e0dRTmeAqEpng+oU5jytwXX8/oqzKy8FhlLhrJ1nd7ieP8WyI88EnXH4r
BTRNrMiU6cU2Lc5rbU1+/BXRXfYKGtdsfopIeKrYPIoraNHxbjrv0sPFeDPdmdU6
YE+PzjcvTM5yN4Ivw9lXYSUMvZdkmvnkYm1KEI3/O3KCcXp2065+s2QAk+JgBadx
rzx2PfYmJdjJdCmIndK64sCmmsRgTU7qqIEIDh9q08V3e/df+vaxsj/9hzLkoL/p
azVlukMEZ84VVV1QbYz+FVqYSuFgKuajFq98hzXmc9t+QMBerRAlATM5khObvHTF
fE0om0ZPjDUmEt8Sf0nixOicJ95A1YXyNZNNZTX1/YYh1QofV1dOASppeNirl05T
PW3rz9sW1nLkLhmul1uAo0mxcN5r1k2plgH5F/tBXIPsGsHDuH5DHEoq2vBjFxUH
UrIjGkCMttsvjCxC2dNkJkRhvilo5PktaCnICE3A33OQKg8TcX/ggOpQsx7CjjUZ
JEjREdFKihC0xW8L7yHubKwKq5oE30L0ukg503UOVvJIn/uE/vBrQAVMi2YaMj1E
iQqdT6YrQdrVqRp0E7LQDV40+X8vgMb3I9qaHeSdIpMPHj8yMmTxZtdOxeE1Ni2f
vRFiysG0i8rDVgWE6QtcbIf2AwtmioyQSK4f/EjQHHhTQ6iUAJk2XQHaSsVFoEUG
UQ7Y5vyEF8IAWQ18U0q7oAnBFLI59XxAvn8rLhn1PgS+pv1L8ujo3ifGXl5B68Fe
Qo+crG2ozdp6QOD515ki5yjgzeJrlTZ29uzmpSPXLqACD9spxqf3yyNpW3yGUnNp
k2X7BNOPpPHM8xQpdrEesZ0R50SUvzCu6ZSmY1L1JNpPh3QaSyDPEYgLcFTHKstX
NaJzhR+OJtkZhYx0/63wZjleDJ+xFOtKbqoNto2v3euhyhgi8dAV8tL9pKLYaMEj
HULmEz6TkMdP6z014l3d3H9de+MiVGagRcQZtt9OMG/z8fbGWyOkJ6JWaEkOqNYG
MRN4+yzMLOmAdv+m4hRBWNWmvd5mfjCQ59S15XPO8X8P6uEu2odoSaxWzWTewLlv
wqH2qCrp+JYVUczdY4h7YStUZ+Vjl3bj8Eq73UwnNJPIZgs3xOEY45S2uqg9T87v
Kb5XtHS90ribP4UF3c7JjjvH6dTWBuUkmroh+mqx6lffnVDSzoEHeHMRXNMqMGM6
1ducTZCaWZNXsyV6TU/5G4k8BacnVa5AlJVW7uItDunWQ9ty/cVkIc3IRJ3/SNdc
MuI7SknjRcscmWa99diEpWZ8MeHm3AC+7gFvRoCADDp6QPF35linj+21vOebVLvV
gGQm0WoIVwjszp+G5PmlxhQjxaLDO5gtsnQO9pWFET6NfFA0HNmQDvOfsE64Y5PY
VOlcSqDpbNOt/mPk40/56bHtp4EoLhNL1kDP0iklGRYFTSgZ7SaW+9DrF6ilIsDS
pJU34TtECe9njj/ZJnMMyzv7Zl3p+9aIm0/Rsm/fH61hpVD0m3QLV7tELGZF+eu0
zRQXhvFHcoYPPB6lp+4F5+McoP4wgjEaI/5DkH9TIIZFn+ZaqBO1plMEUeWlahiZ
gA92lkuDvfMGxugPikCcw0gI4t0y5WkpbZYCXkm+GTyUpipehvKZtRq7r48ETyP7
OEm0o9uYN7+trY5wAhilinR0UwUWa+D5WCEXNyPq6cv8nAKYivEUb5MgS/u53zdM
s/FoSs57i9DlXr7XZ+WtwOkDsUGd2AKSGRdsD2MrdLLrxmWp+RinZtDlu7VCsABh
IwMCAh1VsYk3yxoACPHogP9vP2tsYxSrULGQ9mfzQGD+9j6zoSdDuKGFwBxpLiQF
KpfIEfCg52cr3E5DxAYiUol5S4+65cfHxWfM+WBgsVTCX3N9e2w1lAETO6evLjhA
VkNUUHBe8FrTBbppcuTbapJF1GYD3uQ4SGYO67EunsgvooBwNF3bib55qeLQRym6
lrySEX0P03GjNa0i7zxlD9PUtW/Rsz3qx2gGteLJCIvh/EtJIrL8PTZzvKJGYIKi
w/KBdE74EGAl5ZOEKW6YN81y9l8S6CypXPZtfBl2BLiE4JtpG8eAus36NU3Yg+wi
ePvvqGd/bUSDlMyH3vAbA7yrqm+pbEU1v1AfWkpCm+KOsQyPUhNarsOIYXDfE+6c
LHNx/jmCk4exFY0w4chpcWg6JwU2pUn8iEPOzvvpsIwMshS5ALZwPzdEKBsFQ6Om
Tj/bBhJVcJj6atGVnEUjnxLNr7DwzRkHeAQUgSZqYgXA89EHgQMM/dLixQ98wrtX
qFw2FqkzaSMiyYlWRF+QDQli4BXgh5xndJY29UlMY0DW6wgQaUWSzA5Rfvr3dmbS
CPkpS78vXVNk2UQdZ4g0HlfCJmgP996BSPgp8i6Z/g8OCjMDm1E5QlnRpj9LKvBg
Q3u7TCgwnVbJ+IHHOOQMt5Xx0B9KyDZpCMKOlR4YwVsjiGNB5LwUhObvaNzz91Yy
u9KfcmzLBQq+bpjloTpG7ERnMKBse0i4e9xrO5tn7PK8KvGgzspy7ZgN+fyNzr0o
6IAc8bxMXMpWQ1bEIDmrDvOe71J68Z9wq+3Jjv3PD2VsAryRkHIpis0k9KsOBHxl
v0puXo4S8mUjLZM2qN0u9kNMhJCu2/AA94Ctqr3KWYOSgMlfLpBEvz7uSF/+lMns
sJ/Clehjl+lei9/r3AFkLHG+r4GU3mR7Qwae/IbfNMM2stz0ylkYTK5D/A30TYiX
QYdPcMeSdYkJMMvPGpmXS3oDklqeJnucQA/W56KMZ2uwZ6JdBhl4lj21p+C7KqHL
BROzdv5KI8ebcGintRbkPHE1BDKpw+zMT1WkZGgIKqEA+d/sx7IjkrOsMtVpt/c/
+z0+XFxxoXwSAGRY2TcMLjg5VAW30jfYaFCd6L4hMWYLYirBvB4JqAQyURB7QdPT
apond+sq9QF2vx6NHkcxemHoXo/fAbj1Qxi7PTcs7MotUfAe37QFqMIgtd+ROTHD
Eryh5bft8blx7XM1qlJggFhdsYWC443tUGJT7j6WNutY8JXw0NOuG+6zGOR7cqXm
MNR9zapQbW20BV/WVaV9KShoxSwyTO0E/NwbgFBTEUSV01a7/0JkXcZALWxdGLh1
GzrZyrvwLl7dQvuc7pKWeiazdALcruaDiv0LooHfuHIObTte+H+b+raaLzJqPo3D
+C/rEC4zYUMSOPmEjpjtYM0Oo2oeX/NetMZvAHvYQNfb51XSOLFYZ3sYy/notxSG
2sMbmU28Q5DxD7fPdEwK7ha/xMEVNLnBA5kujym1UJUR1+r275rH1EBH5ZwpvT9x
xe/fmg2r6bAFoErOLk+CvcPdSeykxhUJxIHLm7dNCE98cuYbZOsM1kok8YCbg29c
aT1bJz+95+JgPNG3+BdbmHmrzOxnd3aUcBcDi4Oy2edlVQXQHRUEXKuRTnH37muU
U6ybefMEZpKmQuzv38k0EdXBdy9lJyW7NSpuhq460R70QvtyXHmT10A418etmE/K
ixpF+KSm10fG0i/arp9cALK1mlp4Y3cEFLFXTFOMTFSnKaTj0WusJBRnFA329h75
Qn5RBvd8jAfNWhIJ+cD85iRBwRmFiwr2Qv42p13m7IuTzKkcc3mIQjp8jHQY1HZ0
dWEKrAYU9hIQ4j+6LNNFa5U8iZpyMu3wo6hGj1gIvN/zTUcXKZ03ezKv5JVrs7WG
V67jYuSOvf1u8cZw5zMbDSexHPu1i7Y8iFulnFTvnF5LkBzxk4l74fWF1/EeCYm0
RRqAqim580q4QquD5n7VSUPbohucjABi0Nbu3b1iW7vgIfkJqk0M/r1148h/Iuwh
gsSFYud+TQf10I/ic1Q4ChNyhWTXzTqJeTtEqcSiKJhY0DFmEsdaUwy+UtFq78uz
9S+aeHm/YsADUAM7DBK6VvMoRsSbhnS0pRQaOI3BMADYtuCC7prYAYc/0vzTzVHf
hEVjvQQZxw0WrWBmTjIClFKBPdA3JiUEMjZBdWy95amj9cPN05DVc3RvA/QuCtxf
iZ8uE61gGCODTi5UzY+OhS32x0bzXT1zbkgoozJVDgbERS+Qe70lgWzD4089cRGj
O316gIzYqIThbLCTD7K+HTdPKP8p2qpt3b2WDdr+q2d9pF6vdvAyi920mygVnE7w
EJRJIrjNSqi5xqB5yTPz2pSp6DA12OPLMfJLq1KWHtcvrjrcofRN3/uoWa317SZX
Yxn+gw0xSTzMT2f1hOrKJ/2AvbyV5AgwmGpwXzuptvB0uEWzSzT88VDTGPxsPJGv
tpFa3Y9xLTotp30VO9NXohVfs80yJN4HoNjlRBLfuEGWLFUHbBsjeBFhgE5vChnD
R4IoNlF/quV+9KK7ESXcPbnSDh2GBKj+gdXfzEkRva++dkb+mNH7W79BbZ1FpFUK
cd1vpB6EJmGDhgdphPOXHMyg1DNvUJSru870LfUM4qeIZTgFl7vK6Ggihgsbvnu+
A2NMFO4fCfqAyp6CoJ3uBQMj/W2B2+J3BKDmQi0BY6bzvkYls3fYMbtIQqaYIhPo
34DLbVbNwFMXnW2/mWh1YvqlWev5nWDDoDdsfqJUDCAQNgIq64mgYXIgSmakj708
K+6QV/9p3GMc9q+fK10hbI+QMJcDDuqHd6qeRbMPuyUcNFVh0/VMhzE5xMYRitlB
Q6pAB9AXt1CPPDVQ0FqhGh8c7QPaO/ocVRNRo13Gbxg+VQmWDCFPM6doLflLEcgH
qx0gtlus3IPXploefKuo9AhzCxT4bUOV8y4FQY8L35t8AV2yKQsPAo7XT74Z2qyW
4Uw5HnReXRVXqip/EWU1qjx/LH6srVrvioekDnZrbNG/2nXpsGWm/NtxYu0U+cvX
PYdhMszNiEdNYncmVu3znrh+whHXBNWh1zYihlqZRVmmwc9EZ1RIgxfWcK9WxkuZ
AyGJvKJRvq6g/h/42vaMM7F5xKjsaj2n2Zm6nI0vuW5WptPZGyaOIu2uzu/rCmX9
uv4FBh0WdKSdo7qilU4w6oC7GB5B4yGf5vIMP4zl4jj3nyRfuiNW/BS1kJcy0D7L
aSCCV0m86pyjeVN1ldQGnfmjYkrGJeta3Y91HvMX7raKucLIA7ge5gYixA0Ms7sR
0PTT4NGpwuPWS6QkqT5FB85VwLC3pZZ0MpAEylGb3E818Lw9MFY6drQKlyb9foHv
AE7PMOMvwoefW9U9li9+s+Xu10dvmYHAQ4VOJ0Y9ICi7llY8+qyAxQO95BF8WDo8
n9Xx3/6wOwFahItEDqU5o3xd63yq5QzXlYsGGbU2yspC9GxtNcZR7GKhQkaf4Y0l
2x3rCsfIiwX5QUNqJCPPZxmM0kOg9LUYZa1lITfzdATj0ZCE+Vm5VZ4Xq/rJvhYa
+FZXjIGGSFlZ6gx2S6vkg3MtGbC4YIKcpygbf+BaFeiqrXyYDSFtb1nr+a2DPS3n
qENUkI7eqOu3NB9b2OfgbnnvSdcumyBxUuqfisxFMeBggqoJIfn0y/F+h7evVPCF
56oAnl4DJ39s7+IcRpWT3v+xnQAaBDJfW9h7ayUTfJIS6Q0h1FiIcsit/2LFeNVy
eAX6ecz8mYinUHB6KWgWJJ46ocONlwJgKdWYJ8XjC2JRoKuC0zwmuXrrbp2iDrk8
nE7dZkaT3ZNEx0RbnZWyF3V4WSXhaUYwbfMTwVRge4KyDADF1855BPUP1+c/W1g8
/54uG91TcCedVbujbHn4BeS3TNPbKcIbBy8som7IUCDfDgyswOxAHjyfoylHH8QR
Ran8x/+mDjuwxv4ewU6mWHHWkC7sMta+/DbNKfXv0LIidX+e1Oa4mKe1mVPKscJy
5OAsxILKPoD4ocAcHXbf9H4ZLeOojMAgXYCQnFf0l9h4Ib0JWi/oHOw2e2dIjUW7
Su2V0CYCma5u9Qc6rUO1kRDvjSLXuHnNpgZuWBrJL6zkfcM56zRSMibYePQNhSnp
fOhOGIcPjPKdOuDi1ulAv/u3kMevrFI46M50ktQt9r9LP8toip+vwrVGx4N8Ht2m
tObv3JDI6jU+KYVf+UqiSScqEvWjxsq1x1cW4wg/U8CimuspLum44pwlmJa6e154
+PN033BqRe8Rzu6pQv203o0nLTy3DR4To18JqGZ58SEdfIiBgWSrHgb9ulYZTlJA
uD/Aok4bzQxlwcrWn29lQ4/APpmPj5b79xW5SDC9j2HjDKaBXZ75qFZbF37SP1Ab
9fHu4FmmySewJoEGRqrMkA0xpahofjZw6hMheGr4U+JMKPHrWOvfdv1ailSqCXMc
I/Meji5613hiXcdxDrPxhKEQIsMDzGnb1l0cYk8iTnDi7M5f9yJdyfEZyaiMn+0C
z9vqg7GhkojpW181Cue8llkn6IQdJKS2DdM4NkWnUsLs4tK7ZA7GqQhKcSm9dUap
B152TJydQiy7//j9hlQjmCMOkA/XYFt5eIFq2+gn+d1W+9Aq2nnpL3uGwLUpZuc6
OP+YlDPBgyEr9JIaoF2OMHx6M3nLY3HMfCg2y5AFntIjEr9F75QvYWHjMWOFOa1D
tYGRhidZbxVhd52YM/lkEFoUK1fxm0xTYyzeyOPGAQasnRka6mEtaqS8e7aj+0t2
t2bn72M8W/Wgz0xeRxpxPEbmZ5uDmoZjsjLyloD3rB2cK62BGh9VwCcDEO0TImt7
DiYGknCQRwInkz2HhfhpdRMHP7E9F8aTNKZ7OlLX+5251sUxboslKiaPeRYT5W6M
dweqyoLYH8tadQhdg46Sbm0Uwn1lzTpnHRL2FZ/NsSPd82p4Xl+PHorkutz8qlXj
sHid3uB8E6Dh8zlIeLftDYLYOZrHZ8lWK7sFHB2WaywRXOcmCfzyh5mDRyzE/f9D
rxLs79rHZuWeW6t3wgbmJ6W6gBJc8zb59sPHX62cHI2qDp5s78dCX1rlzMq3BLF/
kcrMFH6GhmkCIZceNKUlVXegqMFRzYbARVrOT87okNBhmVqxWDilmKQ8YqcTRG0t
BzYAJVUjBXXvayTL0sfTflSVmECIUL/hv3xB2TnMPLU6NuF6grH96AmsgARV4pHf
HQIV2iNWBWCB6MicMBkx5HGrVw8U1y7TKjEfbw/r7pprPKKcfFo1SuoD1EoSDzmB
gAg+VU1JGOYrTteJnkR3e2Hc4EKH+qCi0vcPVyggwJI6yRLBlmBGRqhojqsNsfIT
Su3LL1xGmJPKjJZCWXGKiRS1NDfrJxbu8x6N50xGqBJW2yKgy1jIlwxg5VIYsedR
e4rpf70wy7DwEeVZxqcJw1dMBHP/E+7I14mbdcvOQByo3IVhaJr9u921toG2RqnG
fR0FkbjGu/Oa51frjjWUSihKhw0NRHHINVPlekAYiX8ZvAVVkTt//KKjLoJhAXLP
3aSn55KYDd2Uutpq/BzbE9QK1NiKG/KjhxwhHt4Hnau0Q+WtCJkcItm9aEOYFnHi
c4SczAxVlatrtAtRmGy3NssOFya8ey9p3+t8XQyWIx2nDN91lDtu4rUx+4R20f0t
TH+xauPg1IH9beyhszkTOhBL8UZCjOmjEdHB+QYJNI43Mx6ltkYHl4n57Vi5TXes
FYPnXyrTay3t9b3gDmhjw3HFjvQpGl8+FHK7mkCGGTBpr+ru4cySO1cKCAd4HJ1n
M7HykYURkBhK5XK74qtpFiH0XhEhc/WVKhNQL7C9HPGdRFGCL8HW4RsKxlrQ3T2i
fR3NPIyjGUCrkE0wPRG/TOpSEFycB/h5aLvari81QIeKgOC80Z0jUi/OVDh1YtB9
q3UbgAebC4Yxz/+cKW5K60cAlEVhqMHz0N0ZMc6b2a9yWPsY04lpxU4E4XxVwC07
TwkPq8KVHBTLOPYAKRbRe/Sf5a6gbbrdqkep2Eiri0cJTriTf3sQgntWHUie1LGB
sVsN8FnL7AAlQp5/uyxpcFmGDDgm9UPwWfK+OrO5r5S9bHaE6OGgOwNSVZ1rAeVo
L2XswFgrFzfE030OQpn1JHJddQaU3eyFzsDHgQifin365i3e487MRzhYzfEfm6uy
ukgLtZO77LRuEaCVdNc3l/ewJG4m1YlF0/bvlsKlPdbnp7TBGW1og7rXJEvckEo+
WIjw27lcaLl3EY0RqRoNCqH+MX4fesVtaTYjEQCyxX1s6e3cQFLomANgf5LTjCGf
E+cWjHKtRnltsrZ6icOicm1/IAxJgQm05WnEskmzGgwpzr/LUPM48fzwtu0IzWPF
FV2uUPcxz8mndzBHTT6bI5egQOSSw+bpq5uGbUxI8QIc5xbLl9cNrnnJtM54wFq4
6WEAZOQllBRJzbkKh0L+4GKCHYPxTw67Ghi12CSgRYxkvdetCoAUioo4mWKH5EhO
ERlecdTSz/aUwTTjsK7O9/iLV4rL8ny7li7iuv23sjn46YzIbRfr/M+m049E/4Pc
hwDcMEGQBnEV64ksP06Hz004EoOmnvxtw31K0AI2qQg87Jp/1Pegg0KQtDaELpcg
Zt4RbwnGUCHTo0+oTYx2Zi5Dha150LvoIXKYaMR4DuI/TtTdXWvlOXm9Krq4Fs6d
qmlS9P/jitFPK5oh8eHnGTFvYgUu7B+Th18U9OflIhM3wfW1uPcq05/jBvhqIdHC
Nj8ZEd+8j2zL/v1pmoaXlmzf1fnEpJeDgJI2dHpiDjLS2gzQjOkAy8MxjoFGG7Jx
NYD/s2u4jEezf/pj1foy49s3TFEPDjWOssxVdA/jZLjZIsJSHJJEKNW5sS5JJ/fn
8O67WHUld/YAkuXsOZfa+wHVOz2pZz5RKjY1wHepURwz+GddleG9W+oXVKjP64XR
E50JpeWapKAaclxWc6z6OQQNKDa3WIS47d+QfW5R0QWPz7iFHpMpMRji7hu5gh75
nEuI/GMQ304AQd9TeXwAHXesayXxtvSWqsyxI2Fl/GyqzZhdcnNqFMYzJC1X26n5
y+ZnH3Yel6I1OFw42VNjFSeRxbQj2/MIGnFzMZCeft4e1Dq3TDCZtWSpf/DC0erh
L3jpfR1lZpE0qQKLlLMn1stZF/gOeKmbapbkyNK7ppdcAhvJt3IfoF07YTWaPaHE
+bJ/R051PxHbqen/yvx2qAj0g7jTDSM4qnGDIRtErWMIrtKYxjTPOCvg30a/VMUx
L7dkZEufUHelmAkkz+ek0s3+kRVBfoJ5vfjfhsBb9rbS3EXB3c4jcHTEsAyK+0KY
x/IN03Ap5qGM2k8WNQLQQ5PK1Mn9lZGKyoeEiJFSnWGsWqetUIhrJPA3NTtT2GMo
4sQPq8jxGb4fIZj7WJuY7HD0CiW45fWFpKVVq65HMvH1pHz47bRV6z1HA23BKw9A
HnUY0czjOVDFy3gO7qzh+RqAGrqVwy7aE6IiWO6ZCuQCYWVFCpCqFGjvy5X78OaL
SXN+xpdid7bpxzL34oGEHBXdtwlGhSnqSKn/3y6eTadriHb53BkIeeIyBUg6e6Gw
n2ivtx2ug2xOAvojqvQ2BQFRyUc/h5JxR8vw9Bk0BalQZ6QpIQwcfTCtrQJYi3At
7drWe2EUT2MYQXosGy5i3GatloS7L0RHxcf4mHD8+RiLEyrGy+8J4V1Ijz6w4KKE
+QcSx43vRw9YiJDi40mjzFjVrOQwWqFuVzo54f9jUDl6fa9u/3c8QrMrG0ci2iZp
5eGotIOzRa0on/tJrzBf8lgaO1ZWp5/MmVvHiMLzGZWeu6jnrKp/H7hx9wgLQl99
LrRDUKv6GxniJK/n/yCUIrFRT3zvd/UCgUP3e35NDG0jPfYwGn75fSFhWreSWal1
dnZTAsmY0uEJjRPpGIKlwpM8LtxfZj9iyKTrk5FCWpZFib2FnSqv+z6u0aDIsl1D
L+74JeZiGLBnv8m0YgQlVahUZhGRo+gNXb508DJtHIaKDF92gFr6dYF3j++wDpdQ
uTsKqYwQc2k6OpNr31BXN20YS8F94iD5CoYOGFGzYH9yPBqGx40H8QNC/oGC4IRk
okvN5gTOQ4zF/E+C/FWMRXupe67BXjIg3PmzCaxqQOEdjVRRSHU1wcXcb0hhZV7l
TdZPkdK35iwHGqf9GcJjmE4n91egZ8pL6mdqPWNlHdu7mvEJX2JLEgPPmXw9nixl
/V9evpUbwenaQvyK9skBpoQuogZuUr8LtPJOM7Ww+bkN9zALeoQQzgrTo1YBHevF
kXzsAlQe+nbq0gbus1pMd1zAkFa0EN3h/F4ZGWiePUMzADYfZIWJ+DhP3JSIPuP/
j8Y7IXd7XdY7lf7goN9pB3BmKzlN8RBFKFdd8LOIEIjxEkxAxsRPuKlgnhXXtvAQ
HFQ8GyaLhlONXb3zJZxYckfgiDbpW8YIrzD52hr2+FtBhBrRN3SI6mjeisG3ilr6
U4rq9/ypl8systSnvallBPaH+hne/CfHmWq9w8oCZyxGm5oa7orn1TtGuEU8/dJ1
J3OHdT0LVMlmiwaHabjmo28gwwc4AqvmH8AUYHsb8Dut3+M9eYrI+VKL6/2+GbJ1
FS+6tycG8C5QeTjuONlphyZyJu48kuwmXOb0x4x2TjoQTgUTK8UKKAFLnB+9QRZL
1Xb4Or2bWwXKJdE+MMGtDaBjewMeisZaiGsWPGNjfC5ibHi+RX0j8zZTEp/KeJLC
kCsfFm2GPolMiyK6dJYlZLShthq9mmehzQsNHBjGnnkqQV/DvKJTIXyskt002NHn
/t5iOQmx5blUt4+euDD1pUb4u2m+9upUzFj61GouInUJQxU2ZPMv650Z15ezhk3V
rqwJhciFRMsrbo8Aam1vCw1zLh9+Ii9hgfFhzcxbJjsB9Gk6aob1hYfT+KeSlMxy
Z9ChMuC8+WC8REVOIf6YBgQBylEmLXeDoejrndPIJMredwjoKS6u1uulJ/Ig6MJ9
b88ytTR73pGEgVrLRKzLWe5klGYr3rQ8spMlo0yYvtx7LQ6qFBLICyWghMjKMKAC
0pqp5+EPDMfzT/O/9rHe/LhCqmlD9Z69YF2gUGV3ua8/2XPAA1m0qVqT/8dRdlzd
MOxUM/apFjbOCpt+v1CPBC0pL1LMQXaCoC2thObMiYvFhxITqHSzW++0v1/xTzVj
7V2Xt/26tW/mCr7GBE4Ui0BnXqiYyVAmf9UW8T4ACL22Qf8FN/aTjYEtpw0Ey+bO
DUUwPxYeI5xxKrgc+xDxbtXmJRe5Qbp96oKoimSd7/wCH6lL9MXu98Yu5bZMi9gR
qUpCc1kLls3Spo7CLa1x137pRiNrZtDWIQ98WQ2EteavnisC3D5suGS6+eUKB9Jl
vNmcpTsK0FxW3USque+SnPw5nJf6U7Un3MqO9PWD9xqSY4uYwjianS+HYcX2a1dV
R5pWaO46l+0P/Sap9/8NRiSgOpGd1Hg5I4GeYItt+RqLlCW+d/97xcZKhXV8lVqL
SQVCk2NnQmSG2UaG7KXViAX5kiO0LhbCWoslCxAoDilUqtT1d+Sbwu+QZXFVQDmL
kC+5FH4ek5NCksggpVwZbQHFUzrKCndPRQgXTIGa3JFRhcH8jafD8KLT7pOXWvvp
lmWhyxM2tk+Pl9TTwuVIM7av+fldVK4GlHiksnDqRHineLn1r8s1T/w9z8snvR57
E3FepG1dPdIZxfAEKshG98miJePn4BQx3CSEgdZqrJr8hEXVWvMbP0UjTCFvMqH6
vRovS2YSszGnTtMmbCWSqeVh8tIHTWkpIfZmTzxVlqTgbnHlBkdcovWBJHIJGtR9
f1m86aB6UMQ/P4JoLpYnJhDKz4sAyIxerGYomPIJ5RWTNCZTp83ioGvPV28IU1Ff
ar9u1kx6/4d0Jn0+JS5wSrGf0GTVu+M6uZPCZHyoDL+IirrQ5SZ1YXqOqZOFpSRo
0LRsJLKOvKACJIoBdlMTgJHj03Y5qzm6a2OEMVHVDbWBmahaQ6+ABMNlSr+DSIPp
sW50tI+OYtu9e6XWFQIwa51Oio563KypdT/ojd67j7MmBJk/thf86bi2E5lB0SbQ
dw8yeg99Dpd0JJM+J6xO2WnwldYzbRY7HjiU4DiqHkUbiDFYsUNd5Aiu03SGQaq8
RTLovVJ+eO4ZVQyDT+6XQRN6IK5yxj0QxAb9JXN21S9JCCsvm9ebXyr0sT6MtLHm
q1xbAv6irEXJ9bFxLgSNoEMMjqVEqmdgJaVwYEDG5jrlfH5O5p2Jznvl3VeM/EiT
0QbvMDs3IbcsUiW+Lq7oD+urKxwugOCinlhJz9ykO/6aimTorLGgRpy+TBSWRH8U
TKYXQyR31H+1XvJ/u06Qe5FY8ho+AP+/Tr+it9d8yI8YL9xQbLLu2+670wgl4TFT
0iBK2jubsy4zhm0LjuOeFYuzvp2VRgfDcPR7TTFlkgxXxiSylBNUTeBJHNBxTW0W
L+DxanN/rjA7MIs7nSjUV8A6XJ516tjyDpxBM7lqRV/wS+5BEr+HYDRBO5fOzxD6
HN8XLlMykU0Er5IjkLQlLXicvqP9T0fyjGDDTyFFIzLaitlbyBc9mnnSvJ0KgVYT
A+fcwZp7LmD66F/mUeoH7yeaXKIlx4CE0+afKF4bzB40atOwNoRoC/IpXKi6ugc0
by+be9pA2pKsnyzM1fD1VI5VrHuwnZHZWloOvSBRpaY9c8thNnLgyb2pcy7DoZsd
bpznowkbdN6rqj5cf/EMQzsatXhO9iqTG39rEEyHsKCUXZpJa6P0KAu0y94ig9Ty
JneM+RKTqblGvGN6ylaIySpP0brAvGxa8bWZ97kHpPh3W0pcCmRw6X52ukr1bkD0
qTH4gAXa6YS6EEeifxr95nUjlnTbZxA1G7jwmotWV7TjXjpHlgDqtCKO0+aORCez
6KC4YbZBZPSUvwxD3MIETFqO8iBywQVJkt/HRWo/42LUAEeEIoN39yGqprHM/T0O
q72pxfghbrSJsG3YB1OpAyJVNm7yS2i6OxR5Rk9eDG3rsoMuAzFUp1CTDP1KyDtB
ZIwFzKpVFtlUSN90+SFUEpa1PR490xpdCk3VAjRuu5YXvllz3agKP255UX/p1vrP
CGpHSoSiOuTrVJd7ppndLvlSr3OWw1eMvireLyMjGjqeC1TKTdTXfJx+zVGWeZdJ
W0i0NhTfWyixg0OEsZ7k0WuXRso19vW8yeB4m1KjUzmR56VUasL3Bfr6h7SSppzc
iYmtZ5iPos1oGE8V2yfMQb/o2QyJftZJiw3MR5hGIdwZd6SFzpSjhUiK0NMId4WW
LIfd4/jVxL1lx2OdZjrzLaZ7k4CqtAUTzk1ZGM3iCTwwrlPA2hBDotwky0/O7Gb0
fbITYGGboAaPAtnMUMD83WcyzXWjei2aNEa1bJ9752yJzui2u/V5mU+Aajsz09CX
vbt1OgUj7CvUbWpldU/mpbTO0Z0FOy/+5RdogMZ0bQ7uikkugGb0q4ZjacjHkO/N
qMvHwiqjJeTrLiVqcIPunfWFL3X2jIYChQYh2FkKKUfhwjkcWv0IfU4VZh9GA5wc
gBRc35HUVNuww/8Q2kB8qaVwubfIrsmsW7OkoD+V4yOfugsRSAKXxvoXFsoRkBwC
uj51jlURyIMUoGM7enKK3o/Q50mkH5LxFLTy8PoOkDF3pdgoiDjOjK8mGh+KGgR+
d0MW5FOIaVnl/az8UGMCUhNXuIV6F7Lk1wCsGNELK0p4RD0Vhgxp0TDegZEVWA3a
Th+axlNWMfQdNit4DBfG6FfULAdPoL7Dlt67yCtnWNiPqPWEEEn3vIuMAIrM6AFL
aQ2JLUviKY+2HXo5dPjGmyeG6Rnxzf2zTZEam5uBrTc4LCq2osCHx7J7tBlBlQSM
lUMOyP74PUgPbAZ0ErR6m0e42PECSfb7Is2EOnDd3f4xFVtersG6WSF3gYKHnmTk
sXYWD+MkQkwaKvqWH64lqCjFyQw/JRO5vHV1wLdjO9RYNo2hqIb2PNR0Mrn0cots
cE2I0K8ZVDRwMh2bnIWmB7ypjKcPxbmPWHleutUxMqZFiIlpd9lGFUOvrILOEZd3
JN9nzOtzlHq2iQqUBMupU6Zb5oVGcy/jVrdTL8nD59cdM1audZN+fL4lMVvfL8P3
HfgrdKSPLhwwPxHlcEX8gy8pMEMLVSLsihppF2kC9kAD6BQ0hs8qmSP7GBvw3bkF
6/jkBPC2u/fh67Oo7aMhTJelTjTlCC0HpIobm83CEsAYBLPvHeTdO88ahvSSEA9K
0/THxKbhadG9P/yC4YrEzGqh9uVuf3U9gjd23PkkSfpmiirtuTlUvThMSEPdsijl
XggjM5C3KsxfZaWKDYFz6ZeCiB+Vz4rwe9LWpeYN5uaKJM+H7GPRXTNPv8kQ1L9V
HnIqQ3KmuWECRu9HZ3TNOWBaFYbu+W97wYk/bZs54cEQkryGxFqqwAIA7F1tXENQ
2GWAB6oKJk8n29HjZe8JJeAvaq7r0PfZisvhmxVCni149OLOv0oI6TyVdBEdQnzp
lF3njLk2ccGHj5M/NXhqcl/30pHrR92DUSZwkcrrMjdMILswXn8n/Kmwqxmt6A7/
TnaAeWdbMPai6dVaSHglM5RdlsayjYvTfwEVowD58jr4GNQvQoHW8lPfVwhfeSaN
wI+08STs9nyXUzbk7Gng391u1Kamlcr5yBoixTqfa9MLVyp7Eel2XGkop32Zzei5
ptJqYeu4RwyXFh8NGzp43mPMTUQ+FZ5CHGHBLWx0Iab336LFIo7fIf0IMZHIukXP
svHr+MtX9FXj2CTqb6W7yB05xQwS0sJCwV0z5ogzphOVLCTVm2b4nHCIynxiHlyE
HsHzSaeSeSwmbG2metT++SA28Rz4//tZ/CiLDJlJwFKk7tEtMmSzmn70q/Tr2hRg
ifO8KjuNQsVBM+4WQ8rwJTFlaCJrB34ZNHG7W/WatLqBwgfL5vojakK4T6czsT3H
6ANO4FWx8cpHuETWxASpBDNwy0KC9xDtYBD0KTRsbziwK4yMrp4s3YS5uAAN3xgW
2e+gUe4dcoxwv9z/NqhmmLSRFUEXBjCl/ekZldc0wYGjKDQuIUCNA2p9Q+bQqHPH
0UQKxdLgQ8RU5ikZzr8yXO9qIz6WcIk1mnV0lpzcXEkZhYwb5mKPK8CWEcSI73uX
jrJRiwtZC07btodbes6GNNDOtlNV3+9Q/wmZ58qmIBH6r5PTEuaN08toxcq6gBMh
ymeRbKwULbO1w8hhe+Fgxkjte6OPM9Dhp1jvsbUGG3xKKDnkmTZf/aBQhgY1ZUDv
MqNHUpyoWmfKD7EFdoUXoTJ4Kkp0/JpEIQjTHiL/syd1BhgSfspCnPTR86cY4SaB
CWgLP7I9M612Gef+FcjlTi70DffAU/iAwMmg3N5tQ95PIglSKoiefq5B0MSAeUVF
eWpbseSV/FVf5bq2MX/OsVPur1updXKc9wYTL378hY6Ai8cgUkvUGYL8VITJXhZK
JHG0cBGGBlTiHrreDGJzel8ymJElE8m/NeunchQxbSY7daUuif9aL3jv1n7D2zxi
AI7INixLYsGJyM7yA4s/ali6nVpWqxoMWgD9TcDkyXgTDCeR7ekAF63k3RKXCW3R
Qgt+XYETMwFfa8TvsWa7VPNXwFS6XyAHkMfMW6KHFncOxfZwt+OKJcbXlQupkuiM
TPfCBQea0cXySm7VnhRlMVIYMuwbhTbA96ZVcjbosH0ZS8amFaeQ1k3YDWlynj6L
AERHvsbA1CquBiJCNZu2bnBx3qbEBcmzOlhIwI4M+k3t+E4q+VdNx69sSITyV50y
QlNdjQzSfIG6PH5RuKznB2nWlTOWEA8tXwrrgI6wKvry3UPDdcYTs68wZT2CBd2/
QaxbphC3p2cCfCKXklPF0MVF/NCoTtCxNM5W9r+MfeSeM/14dmK+hZ33oWLU2/Ju
vI02IGfD1QO3WZPEbfKjZ5hy0ryyUFFzCI44xdHBx4CwgZfnQIBhGoNQq/UUHZei
Ln8WS+QbK8KFnnXV+bjjfuLytT78E8bDXuzfF53+8k1FJLi1p5h3msSORYRZejEY
249I2UB3ZCFzgUNSNHVTe4XZEdFsiLRwkih3K9UIXM8tcD7NZOHE/HG+AwM+1wMC
DqHw6ojVG4y6IXB+ENHIf3y/jXlstzYRnzIVG6pB/uDdOWChzB52URP693TBsMjZ
kTWmUTyPkRnV4dF1+0Re0o1cp00B5gT629QJH6whDs17qy5kWG3qezJaN3FqlnPt
a/MGYjTaeyxDzlJb3K86Q9DrCg7y5UHm582t8PjNE35LGQ8VVFaIvKQxQ70s7cCO
oEhpV862Z2RP3VVIRAQdrg7TkidcrDEkCT224Ja2bQpmVdyeNqgvqQPFgsLesGGL
H6XvtE8QP+gtUbPivXeqkGlHbc+d6QbP6U9qHcIMd+PlZLgcWqddCJTkxG09Hdqj
Ej0cF02YZrS8q91e422pXszUscNOMJpMgobXy6YJ5l2vGH3X4BEz4lGZfxkWbp6i
xMMjM6Ke8nYijJ6D6meK/f77ySPlsisppKsSiF/DtesldyFRqgz+R3dh/SHMjn6Q
yzpmoTmvzlFLYAEL05AJC5D57aMgqR7ZYQO3AG/FqMCsMA9fSWY7ERYwYKn4MHfL
82SFAy+iTJCv8MFVqqd2326p4jaic3fX8UfJvap90SOVpi7B3CFtodLXj2//uC2D
R/1tjwtbPaxVz8Xxi96TKNRR/QPft4ItgUwQ8zZ5sEwn9ckWWSZIQmT669tGkGQs
etT6hICBykOKnYDdi/iIMA3+jGwIW7BxP/Ed1kpsINH/0Ls5zZoYwOEYiK5XuDaA
YnXlNCj/NSXgSfEcxveUWZssKoKXBHb/psTfk1ZXP9OGfLSJTmA0Jp3YXF1IpS1F
38j4TxHiSHusjJeCV6DDEMd2KVad8Pp8iU5LQB3nqxlA0YTYPyYWv41sB1rWYH69
smvfGrUbZ8LeooiUrDs5241WSFzqDTyXATusu+99YnRlwPoFydckuYLc5U0bXvov
iE2h4LE8j4nyKORT82qMT7M03rArfOtjwm97Xq9J80B10Tfb5lxYsFtAhIOkOW7v
wGEsHBlTCcD0x2IjD+NJrx3XVrR/4xhF6ng0BLWDVzJr3TsomQBs6Y/Mo53OYaR3
mHVoGIXrs33OZDLb1aB0vMLk+KjnF1d2RmxBBRj6aMsRLOpTiwKH0rDd+OiCYyZq
7JzKrQVAwtdJ591RhZaU526byPaEpS+4xHjhBut5AOA+Bp/INL85mdSacVaVttSL
hPF2imTS/ACq0PXHW6yB4CEp1063Pm5LYTHaJWiXKJrDNFtOIZ5zVgXu0r9Y66tI
Vp65jOTLejTeva6Dpc1eG3Bj17OLZFGtdOebwSRP/yk8eWsX89e4rh9RotSY4fnO
Ba7VLO37dAKzKLL9v+yi6UpqChpMeJHJq4lnlygDbp5BiXf4XLh4h1amnAfK8/jp
a+eA8ZGfAFT6ozx7TSPID4qMRmoQTEZFk6pCWuTIjEeDnTrlrND7JgCZQdpPhmMZ
3EdJlxBHwoV2Lc8dJ9Dghnl8OxaWYy+rQ/KIiT3wLnEDGcWUKIdamJGzRox5sAei
LkBuCGpFgQbyUGY1aEhvqBuQfQuFTrmjnCTFv49hkbdnrUefb7Ia0OlDeFBNWkh5
ynQbOVWXuSeKOJJHzo5g2BUXU3ft9LK9AsRiqVu8uO7eNXql5rKmdXJ8tew5HP9X
+bfCEiVNOPFzn7QU+q1IhKNwJzCVw1s9erVcZIV1ntmriuxIml9u/Rk1mDVrF/Lz
UJMl+VVfr2cHsuy3HRqSat2MedBmL0MuXvl5yqd7sBwCIPuCZDoVYnwl2b8GrMQH
BcfFgLn6VypMLeNarXWYKvaefvwn1uVcJDwy6SCZ87UP1hz7horfCCf/XIPhk1mP
fVyhy9XdLyX/BRYvVuf7+ruwndt65tKOYafAz0VZBI7GSplQSz5vBBNUhXU3rSSE
PJSiTSYdiWnqw/ZwlZA+/5EG+aWLcANojCJLXZdU9EqdZiBWw56C7gbYx4D0h2MN
WCSmiwL2BqviuBm8Edseijov7Nco27Ta8sObLHdgiguzB94MYi/g2nFKL1j7wYww
1VDkLLyoIFz7FU1DIFMrCnYRl/DnIYPGapSUONz3Ctt/EwDrahgUfAZtTNFY9645
5d7m/C3wiEl2zsGNGAfGXllKfV5wRNKf58O38sKXdwunAOneNiNRjF8VQTvY3BcH
Fz7K6LqDEumcfyiwkbhIZPPHnAbF/8j51JxqQnLR/jg9VRxMizcEzuDMZOLCevi5
00LRGKI4fZONWvslHQYSYDBxW11AzE2SehS3EjSFd1HIKjQ8Gmb+U3YLbd1Ur/Uk
G3Rf079Yttusa+JpV/FEyi7FT7WNaKSstlZqxRXe0jjvouKh2g4e0JoUCS1GA53u
2uoozdItENPfnBVeSCZgcggJ59l/i8HON2e9lVyL7H0/GivYHxlmhZEGxlZMGwuU
qGoLwwHCEnJrQFgtMWFmTtiZ1OwXigKSh1DUEvKUPTlvyU6ycTL3Hq840sK8mTy4
Et+mBnOKTQqUqzlbatFZAljNWJ+d4eq2F8sH2WPbH0UHcfiCNmJdHQN8tQg+W9Po
Of0iBYQ8c4c9/zZOhmiac9wbCa7Qdt1kxgtHifrvgxojYhVXfxVjLMonOE+bdaK7
AWuCEyrRbIRqcq7xLwvNihZ/ML7DeVzH0R5Fv7uohix72SeBAk/ncfu9289hQ6Jw
nw+M8x91/MeKJdiewBorWY/B0r4FThkIujjGa7kZvw2Pnubm7WCush2cBnYcrC0H
JJ5tkxo/8RsWekkxoEtJBGcyGh2LjLlCER6/U8H5sQwiWTafiFq2tAmu60Aw5gYk
4qaY7ffPFr+kszn+zqz8Bdd/cZD4GlJm4AGh3D60Puhl/IgE4B6SSDhLihykBJN/
lHLl44eU7TiTOJ8r8VjsZTCs6AOJGcyzIH2a5OQSYDLGDvJmS63jQ/cuP7n8lANe
C/eogn4wYutP/r/t55Xn9A6uO6vS2ty27TUpvwvxixv0DyoP9tRF04MeMDzwRPTq
VJx2vymUjqqZIaJliaSvP80syRR8fArSJd3M3vSqiactyTUD2hop+kNCi/5XHaLO
6iBptBX6litmuaLI7i0U+uPalYzKMZinku2to6Nh3Zb9SGAqU5yEahNfuLjGi80T
JIcLMsX12owK4WxEsmvl8JMTPTHplsIOdwM4N0JFCzFs7j9TaIgxDoy8PKZJdSPg
g0rqDfN1CymA0bR8w4aaqdnLN8aJ4IdY+QXjzlhrm+WpIrsnGEUkRNEPgGMwpQT9
sWhO/9c8tIJyWOB0KCIh4ZHAK7XTy5uTEwYqZfOKfiWZ3oLe7D5gYdmHSxr/5aTh
N/upE5PMXro7+LyLL5ds46gYhL5drbyV1LbKHomZhMPt9dOslKB3GDAT9FMbsnMa
j3+K75McRMRrPMZJP2VhFi7CiJLvLWuGw06YXMNIXePE8eU5Bjt7Zsau9n7QueWa
JH5H3bVXajnT+DELovmrbjdVjhgZAYyCmunKbp06l7GOgh85EJAN4CPR3xekM3C3
yagt4dpMVv2ttFiSxJmhkEImPVQLxREyxj0nYBaAW8/1BDl6lOSmziUnXqFPJRpf
kEy4YLZnC4X7ZC4uTPxnSJTjEyhkhph8ZNxpelstS5t5ckW8hLsiMDddw8JBsvdb
nh13A+78DshKF/EH7UBYEOXyJpLHW6C0ckQWddcpH6CidDueMP/0guW7cHnH6EAh
0q7YkylDvoH5bIvMqZE/PdZuQgCvTqFQyGlSqv35ayjyjbV6zdCSlilq5f8uTrhS
6Z/vPLUBxRoEge66EBoO0OxEvYN1U0fVKyQ4ItvugmYLMCwYTpJScOkROFDGIqQ7
zraJlqlHAASDT53+fuFbpdOyF3+EXmJr0r/1DDTIOKd/ZK3tx8UAd2JnD5Q/VdYB
iPRb5jvuss5ioYM3QZaFr38Podz1Wti6I2GA8O6z1vlGPmWD+wfqYqaYu0me6sbg
YhmSk1GnYCr01+SQiBuCPN6GUQs9eI9k2JIMjeVHsOnfL5yT3CoExgnhnrha9bNN
JRY9aNnm8J6TmOf2wuiQHhm64gTHs8NyaYK0rt6a9bNv0pB6/c2pvOGWPc3EOaGz
LfUzm+ALZ5wA7Jf5iJiagHRXIw2tGcYcVXWRA6udW2BvdSEGUnfGJvYa4iLw1ZJr
kg/fyb66t9RTEn1DSH1bI44qbAtQdWoYMcKNn65YK4ePe54IfdLLki99fWWJU2Xc
9oclm5+FuIIV5OpkvKYw0WyRa4PCOzsCarYtkdvEKgz57Mklwo8ttq6GeDsAPr6V
I/MZNKfd0hf6oGOm4KNSrF79Pf/7G52TkypqV9WYXBpE0gIQJqHzUiLGwi03Cpsv
HFz2kPhXF+qFlbhBWEDfts+WTZu644FUz/U8A4l5J7QC+PS/lY3OdgBjru3tDmcf
e2GsWnERJawpilX03MPSnqwgh4PJpziL+tYK4Oh87kxGTvyVrrMUmNHHbY+xTnFq
ObVP2e1mqp7uVIoRXNm4GDrIDIqYdNCGA1zsw4R2Ki46Xay21G61njv7zVjC7+CZ
LQM4TnCdMsLKwU6F9P7tD+H7rXsB4OMWVDfsINcqZoWkFPLmBXhTQAxvPNd791TS
Npj6Dy+TmordhOb/tthNJLIfhYljKQjHotXCMmJnrr4SKzgGHuuumUZ1Ht1HzWUX
j9H36pzBccLDVPgZbLQI6MKmnwu4UGL5e6FxTXZuSUYZe9VDr03ARX/yxqx/xFDc
wliql+Q2q80kO3lOy+Po9WVafue4fMqQHp946v+OGnfgVMVj6VnmqxpAOFxHzN6A
N8ihL7A1NmvZgwqyJ7gp/Fqn7z/7MwMxgwZI9BGoOwStP1FUWkrLKbiVF6DuWpdY
W1VqNDhIQRkNHgMVM+h58BO4NuRgX/uy7Xzb35bwImBkNiux+G1umW1s3uHTyquE
7pft4wa7FLYcrdom+HBvMcoOmE1X2AZ/YC28da0qtCuK1Z4fy23iSYxWkdgs44uP
RHHtoOnSJ/f/J2/Bgb9sWPBQD+xOIZ3axGrvYV1VeF4zrH+oZjNp5NiF6RYzrqWN
/KM24jE32JY0IQ3NJB08F+h+gph96qPvAjxu5dwGNArcwpaAcyf1+jrqW4xYB4Zd
ZnUBWcvS36As8d23Wc9jdzTHksl0+6lCjFjd5fl6oaw6UsQ/43bhiZuqGMCpxo9N
h3yyQ1SopDfYlsnrUPFIBj1mUoBnQ7Gz1RFQbNB1Z5iDqB3qxljEvTlmifkpICCV
kZyigJ4keyHUIoRTdC+0xmA5kJXId9B6pSAQ7DijTc1pmohymAwuwSsZ9LKebyAp
i0gHXVOkmIF/1Da878rmGZCeJoZSLSOYXCJrLyyYK5UEvl1fQiQY4X3V1Y3OEgU+
pbFMdsi6gdL0DFUJrSkNHHkrUUrSpjSug1zMGiu+9ZeDFMlD7IMEqtoS3I7hvuQN
d1asGw3xaPhA7Xef8ebqtW5u4uO95FqvbIwF3NBbc/jE0xs0d+QFCIXo0l5+wVTe
i0PhCCXvICY92i69u0JWduuK3D9Q/fiam8Q2wdLQtl92FlX9T832xGa69X/ebHds
sb4dZPPQG4gSXrAKPjA8XHrdNt3F3GWgjyRTJLzlXmk9rDdp4ANz6t0nwmXNM4pG
Ff7l2YZw+jpq/Tj7c+qmCVqDOaUjfCC73WzriPYwu010WpLO+E4NbXwrY4oJVdQH
lHuDf4LhbJMhxq4aUBFG0YchKVjSAGJ5a7NB6C7zUKoOk7Y2V/fY57vSo5+eg7FE
kkTfaQcdfklwELRMgArdNUzoEuHN6htdjaRL7emmXkuxvKIQQQiY59g3cDTzZvF1
wafPxPXodUAniGNlDbIycjwStbmcITtqpG/O0o6LGrPiJqeU1V76Xxpl4hOuvy00
QEaZJw6iEdA1szuJsxqoe0xlh879DjIoZrOo3JGZ4UY6HBBGFhU+0/K+1zbws7qT
p7NbkRtalABCNGIaFfDXpAUMaBU0+19afZiZB9Nqb4drTkrWx7EdWZl6tONvpA97
7QfbBqIaNpfbYKB4JPZW3zY8i8VqOYY/vKzBcA1oUavsFFTiQyx746pH4dYdiJkN
ApyccEYtFb0RYOKfEpDQBIk+XODk609849C1bu2EvMgslIpsyT/1MK8k1VTTlR4N
s8WLUb3TjkmTgSAWLPblwGo3GCV/7+zVw4bJ0uXASICZaDCcqLMz8pYw1hEQ19ds
uzKC0Fw91NSUTtF83mmEyjOGz+TfVriR0EXwjfz3HPVXu1Ip2W7GGwr3O/O+z1HD
oxHxzlf+y2ArVuVPwljfNJWjxPCeVlde31y76FL3uaPMuJVIi1rJNX2+2b9R5lxC
cM3YWvShlxlkB3sKS8B2XYxhY9QopLEDROYEbzwosmwBfUJF6rW6GGaMT3XBJlzz
Y7WEZENSCo2Sgrg6Y1Sumua+otS+/2Uhxato/964x5QGO/vNSwJkNp2MhFPVJkUT
s3DrBc2To71vvi7fbkKBPoIqxiIkVUthQP2FCAxcTfNRiVeSUZRODP0q/v3o/8Ld
NWTVkOLSRCvh78gKWHXQEFVGPT1t7EYDAz0Yz4xkdVONg1WUzI07mmsb2JIJm8gh
iJs8txhwefPcLea0UKr74kTRiIbu5B4vFpO1uWb3iUgnzEx5UlQh/YWT4yvaXAKr
5c/RxlwJW8hCc4kMMeqhIY7nlHRzY2/h4efsbZ/Od3zi1NIwibisFJDlHgUe8iop
7YYsLsnd3u4emYXDpIfw7eKba83yVtSMtgOfJW/lbWo7N+sgUbWKGW9rXN69pJcq
iU5Gd7m7nDioWs0Dj+UZMsLibpq/MMNxaIlPJ0oxoMkEg8m4LRBL+DCSQiDy93I4
nK2L7OZZEmtMd/yg0FLjTTdCE3CsbZyDlJ6CjuvK/LGpilfnWsJmsrwkgREDXwnJ
qEfOd5Q8mi8Nto+6djRhyqVXXlIcB7MdmwDA5HOvAUkIqzzELNW7+B3PQ/r4mvII
gNi/4h961SKbALbW95y3KHt9+r3C0yMptgzK812xMBP1dr3ShrkIkK0Qsvntwr2I
UnUOlSSRrGYDpIuuAzDgDfbOCMCiMmFywb2R8avq+z0Trmrk77E+QoOMAgdTdxFd
CEDfCwe5bQHakMN2kcm/+eOjGx4eUsuRkjitac54EZSsgGlkobDZ8WE599SumzIB
I6iAB5cO2h7ZOsomMf3S/QBhWkxAATSEE4J3Vh2YJ5clbKMfJDnm6BML+fGzP/76
UPTlJa5p8zLX3QvpBj5meNbwT+cYxk8x39KX7EPe26sQT3MU9LpXWKqT7+s/EQgw
jgFkg1UaX5V9VVPERh25g03HFWHbCgxZQraoyqy/qAzKWm4dCO8R1pwYZbXYYVvU
yVfPFFMqgUr+pOZu81iZ1DZZKnnYoKpiBIGDYLJWIITjBW/tgNPSZ3dkj7EdVNPU
3Kg5NQ74Fs+7/qCkq2omYZdUbLxLlk3wwMp557nvau075sZkwlTtt0ZGJX2hD2GK
i5JeUB6YstZ1HW2v9SVUqBXBaM/pceJLq0QiOxzo9vxtAEVwoCcA2GEmzd3SBVyJ
4XzbVtAI7D9XyekGvPXB99mSSxdgIepPxK1eYMFvAS+/2xZDHzTDeVs0k4qXTv0W
QZxQioHVWNiBXRL7I28qzU3e/YIZCjKZWqVh2Y7+kdtEPsJOQOoboWbEf4bvcc+A
qroDw78vmgt7s1vKRKUvFjq5Dq27Y/1juhi9TxKYh2uBp805LvG+Exdwr4JYX+WK
ArtuHE8FgYwn5KaiXFWfL8jnRfQBvVtPV1knqKjRuMyXXDkmJocYH+9Ng0j/mlfo
lmGuV1Fr9VN+A/WBWDmkn+sg7VvZPmiMMKQmC1bGAID2Fd5LGWqgbQeWqTICZPPB
6y0C5aajmToKx83RyW+nD8uJY+m82UqDG1PJIxGQnPLu0MZT3uSVvG8ZvkZZeImb
0Gr++lg8lYqj+NWMRIKjAF641mXO2aBuySgGukebGFQxnRwGUHKDWi7gKVTfiTRo
dA+9nFKwfjWZWgoLZdQ+2e2cb3GOlB3ou7XFljK+iLYnouNPa0Sc9g9xCqStqc4M
AMnymOeaCxkyiD1hEKjqe2AzbKf45Oy+uCIAiNbIVJn0XnQmk2jphVU2m25Ry1NI
DFhHSGIZGVI30/NSZVP9w4R+/QyzQgkglN3ZjLoENv/oNK8L9ooMDN+g6dirkdFH
yNRfxDeIId9ykdlaUxAEtgqtbn5YsotWPyMpSWq3ThFUynQEVDj8y7oPMQjDzWLF
M/8tZ2f/Mol4PCLUa6lyaywobt8Tbj9iMwMonQicU0fHEJDwha8+2NqSYmamp6lY
Pkv4Jic6Q9k/9REVvgYCSCRd2C3316FaxBqe3hHXhrROYI9+PUzyJdI+iL7qZClw
JTA6OxJoVCksT0ePgrCMwwmGEi6OODFigInybPFNqC5oOfdYTIbDlSqz2o7hpYxm
bS65jERINSWHCVRt22IXfnvPeFM22RrM/0B4unjv3a1qNL1rbn6+vk7gzsS6i6PF
b/EXaERcEoXDxxZj+nA4o7C0iPLPeO0zIOS+U4gH0Zqj1maovsupX2VlSr6LBy7g
qmL2UKHqRWbkMZHsIEYkUccOcVVXWLwwo62SaGv7ybJ+eyRWSdUCXFG9tMWGxVi+
e4pnQ+FVsXsZS86sUc12BBM9fT9fek6fiLr+gefYxYDrdA0NvfNCL6sNwK5MYz9I
lOwwQB5DYE2vD0Tg+jiTesnVDVsj9v6011pOD3TLVMOiQyEwFr5Pjsc1wlI06X1K
ypN0fbW7S9/sGeYZ2ZpqdWlMgehd9nMHRpIm3mEAARjOTy8CL2jnUP460GIuTUAq
JBDE6UnLrEdu2WycnewEd3VDGjoHL0nZe95h9nW56JtD8+ycuy0NpK+DCBCSYpxT
T+fEswLuTwUPDgJcJudhsD2IHbVacmX4dfeh798Z3iAh1Min4686Mp8tZRnt9UMa
4GyV909IUIdV8VfTJ4Z0lqf/7TFWi1E1Mb41NIaHG+oLNgVUo6nrqiMEA87JenEs
9mYn6n4ojIYnzJHPS8ifjj97mPE87K2xtz2F4jxLaT7gMjHPT1d+VQaqP1xwcpLg
y2zzVcKm6aYro/EYCIphVCCwZgZZQNwXU9omfOc9D1pWPQnAaVVViskdT3qJeck8
AYgnoYIIS/WSbvQYt63mXT7EGC7sS0gzla1WRAJY4sf2hMDajJjtHV3qCl0LF18w
HcEZX4Tl8ADuSM1AehNw3bCKM+m5GOCViMlBLhf7VeSKZBapSvBcTzppy4oNWToQ
76mRCePU37t5u5I81/LeaYy15AKTw8/2wlCWl7W5iSYCv0CjOCF08qkYlE4xmTvf
jyr68XvE8hxQyz/V8Qo+0Esi2gDQo/KKJ8+boWPoivr2u9yp4IfIVPUrrGOOPexW
PwCtiBLTawwWl57m63WE1yL1mO+OXrwD9gQbnJ/4pnld/pRICawHae1pbR/7tiGb
I2Unnv7OtVj26xceFcg2qE7f9n5mfTVmKG+XjmOAdxwoI1p1F31El+dMGNO7MMEy
V6cGvWOFljC7STqyWe/crnNcopplwSnyVxrkjvAjTD0yomQpFlCdbt1284uIbFE9
Qn+RJYOc65c2wiGqIgAhLcuZnzIzQTQW8PM+tyjTCWjhwTrGT+pAfXRg7OZQYfnf
L3oAEtmpoUAzec+jLauUW49N85wEnopnZzb84DVKO/dDDOyD73rRHRE5L3BPmjhX
wISiRLQrTZmSipAlyyelt6CLZ4lEKoD+gjrfeBtDIhPRpFC3RYMhyWQ54XEOQzW0
46o8z3UYG6dRhh8KPNYcuoqRaXs85BU9aaoGUzKAL9ZqSnqdhbM9cqSDntw7Ed0+
ALTYdH0UKPfmnpDpMZsjPlMcH9sOidTN1PBl2LxeBvpOpXB0G9K77rauPw1NdtSX
P4TjCtxp2Z29RUH1gGSfgoDgsJRIixbHFCPH2zgKaLamz4f1ZhhrufrR1kueaQC7
IGEi5SmJFnGFPgT5YPQrLxWZ3tCCE9teoVmai0BnsMlXEyaGxtwYQXb0IGIxLhc6
QszGG5OWkO6eenf+NGhCDs5DvSzNx+cla/qdfTuXR9VlwwBGBmvitNP9rBp6MnqX
WRWc+IXa/Cvx10Sep51QXi8r0BztGLngWXnUcUZ/Iw77fWib+uT02Rq7/7nZfkgP
GWGeZcEs0gVISRRp8CXfwaA2goyUVbMpoTl/7ml/s/oUlv6mQeL8U+zSz5kOenB7
BuvNBB+rUm1BiF5wvl9HdemjtsMJEtbonyr2xEVu/6q8WaGW12E4XK1/qivPrdPe
vtnAp8FP4cVyawwLOq4ZaMnHa0RmgMLH84OB+reXWRnVOgUvbXvR4C4Mq0iD3gGe
2RLq9lxfK6gHCyjuYCt2rii5sgdw/xV3UuKp1xf2Wjwiq88j2l/EpV88QlfmUnAi
OBSalvyiwz7/Dm41KCSaWA5vMwziFyQ7UdekiLWFRVGwFAM5VC4oHhw2uE0zQ0nd
UltOHBJ6H4+PejXx2KtwWxDeJli16QGY6A13d2ai24O3ZN6BsDnJRX2DCxx6R/8p
09X+GCYSbj8FAUOemgrQhocn4XXWgUd2USw+mzwOX9dSdJHS+PrT1dEzdhms8OFO
QAHxFMPfCzsVLuAit0S1kRC2a0Bu6QoCEWbhMUG5Q42YH8l+AIQ5wbHnDMQcwL47
mkzkVJFM7j/ufQmgxYvyEzHdpOyQZkZUn1slup42rGC+pUXlj3Y4T7FnWGbYD3Dn
FiasSV6ROmXCqS5RtlqK3H9rTNOEVIJlfH+zbXAgYQpVd7n5mvEO+93gW/ll7g3x
E2ggYjmqxB4I+pzTwRtOfBGNwqBqVt1dG+Ha2gcO2DZ6Z9ZJtz7x6VrYq6W8QBsI
e/dJBTeb1pKQEAzktXkOBSqGrgaxWGLGqcmh5h4NCNgW5d7mqAEtPpujk7+T6DCh
txzNErXIH8ue0mZbIuArIon4dALRg/lq8f7jq48co3aQHdC9U1HiAds/hZ9E9dFl
DChEWufKWuo44YlhH+9nzyNNCRRm+WSaXN8+EbOgzkXk4TnklH2g7RisWDjhRRLc
U7RRM5kMAxwsFV1rByqn3IRJ/sq80XQINzytoA4Nko/yaRUtsZA2dqB5kCbeooWs
alfoU6/etyi8fMYuvvmrAS0lgXc9v9QmWS0Sbd3C2br2HDpQrglQTGmd+bhE/PJn
PCmdnXlRqotwvZrZEf/fIpGSoaEsAt43TnzHsQ2e0tx1jGdesgzjEexOKaOuAyZ5
V2klRM0ZP6PiqWc7XGAuFUtexzWePA2eFhzydIv9WOq0UTOprj7lfpQeyyo6X18S
H8ZCiTJIPT80vi0Wlpx9yIt8I9inmB0Cf2lTnev9MGnCHH5HDkh6/Sr6WXyVnntc
qbMcM9Kx+gZ3r4403elpAt+/KkDOWlV9Db9dvOCBaxDCcyUCYot39LPpGoyPQt7K
6z2tAlAe2MzYnPZm+yJuuDWx3E8RQwz6ttZYG0rdtfC+Fjidccs58Qkemy3G7WnH
r7HGJjq3NVhLtuGuEylpVBoxj5MGw6hhsnZ337CByVGb093fQ/DYfeCsLbwSpNV2
xLj9yuLi++Bzz/0hJ48dhFiSrX0bMjFeTNOFJ7nj+4LHrkBt/8Sx7SSXF4F0RGio
NCiZhtkNwH7MT3baGeRJymy4Z+Rnn3Tymb2aBJ94BqMZkbVF84OLqqqS0IsUx6ij
Tx87HR7tFn2fZi6kTLcW94QBFwTCTiAqDx2IWZKJOK4Bv/aZhJoovd/EpW2T1SFr
rjKY0PPJZihJmR4tX9UsIcFQC7yrA98QaCAp5UFKOMD5PY1KRsGYUks1m06RE6WP
DcfvkXeBFWGMjFPGRIgYQKGHg6F+Ar8TTRMZOGUAtMLJCHkkhvj7CHMbySOLXrX+
MHFTgl8kRDmb6cEJzYTNPO3yJIYS//6ycSdE9npbVLrZj4Ak4A6mcdBopjWAmPfp
D6vdMfA9/iLYTGNh7m79dRD0cV+XOcsKrefvUOMp4qu5A+MyKGeIOAPUj/mifhdV
gt7VPQ5w/Pf/DdrdFV5Z53M/izeASxjLplNPKFwglZn0bQsxVj4KnNrjYFrt1F2p
9XONVKzhAW39bwH7Msg0yU7cl8I2MaX1qMf38VGMJi/9jDNTDnrfa/UvQjVe24vK
bt0HuvG1v1z3UdvGpbZPxDphHeP2V3ASG/vsK2fDzO629WIz+IMsSAsj/UYGTSN9
nXIS+EZRSIAq2bLvctCvL0HdLi+QAkTR+hLAQs5QxOsTP6yG0eFN/wtHL85cWwLj
NRAH2Vu3J8nKpINU2mcKgLN6Cd9Eh43L/Jc5O03d7OFXQ0QW0kUp8Lu+pr/WhfjI
I5FUw0OGijyR7XMwuqEjEl3SBeC7N6g8rYvd1yVGacSMhA86gwsMFtw6BXCMPDtb
KWKTD5+KKcVCmoweyS3vtrG/yUtentEoNisZ8klv2jRtjfb2YTTa92i4X5tpMRiD
BeySe7PVuqFe6uNZzdZhAjsdF4OdGZzkugk26Kk+CeiCPQnSH28tJ4dcxyB9hvLN
3xWDSOmLN3bvw0+LNV1LFWK/RgKOOI50O+O+LaVi85WNWCThMVRHsg1XSd03efH/
pGGt0uoEih13NC2DgpsmzSOnFEJ0tDCT7IPUa/4O92twp2dstoPNsFdS9wYMSfcr
DKC3yGcWP2QsH44mpaCVrbvCXHzs8zS18z1L3QI0ewb/knMUVOu/nMir8b/aeLGC
wOOXggOQ3KnW8MYd9igIliJ7r03zdU+kX1kDdyAJiCViXNkZ+7WdYJZZqC6AX2c4
n3IcDKxrhQH4Ez0wTa+XmfdYnQQScPlkkniIlTLLJZGXWLc9QlvixpsULhHSgbLi
/2neeiAru3C9SQLUFcn6a6f3652wdF1m0Zrk5PMRgK/o74AKH2qWeNvHN9U1tMQc
rAzTgQ8ejPvTbAeIJjcxTrULs5xkGZ7mkkwJVHVaBpG2U1MsxFA+vpTKz+glK/Z7
q+y16jjubHKyD9FEWpocleR3zFB4iyLsW+C8pgN6CRdwQ4ROUd8N42AnDdBzjkxq
IURgbz09Wbhkf/6t9tZMZoKiIOWFlAMi2gP8+TlwXifSDTS6JYo17gijppzCacj6
y6aeu3Dfru4+2Ehn/flRqTsUj7zFwsJU8fBGb+v9ZK+S18CFmPj7pk1ZBZDakfhg
8XssGS42beiSphz+JR0eY1o8AdTj+lOFXLKQ2FrIJwWReoCyybcqEjn1AKCiLS64
kxK0prW3wHW74K0m6LkxU7JutWy8MLxeGcYR6qz9lV4TtnOlXzZbG41pRGa/tXLy
UFZr/ypV1VC0HZ1dVH2Mio+m7OmVQsqCzmcRopaa12HA2rBZzAwJIp4zcx8PPRE+
cLinaDnZgmYMjg7T0MysICFcAOtWiFONfPy816uiDx7IzypF2uGipAIlyA9NZWeI
RYUwN7fJigeBMyLkp9My5XhcChFS2+/R8NJ9oHkxv0opuGccCh5uXKd/+X9byGOF
65Uw1tEeMYgN6JpT14aShG9T5HpCvT02/MN/snHCLszUHS2fL4zd8dM+HolZRKev
wlqyrFgiihKTq9Sz0RPNaV2RDNR40B+UPZ80efTlTFju9zBDLVxiv7ByyYZwXUYx
cGYuosdtqzhYBzXrXFDmAJna0DIaibrO7yW1D7U7eTjJgTrrtGTbGvTwt5xM3qef
2E0xi970ZpxJ1LgjYgsv01JbN4eOCdtBP52wmzPXgLULMq0GrAxFXcvpmsj+WJLi
MQq6qjGBahDDW+6PQYl+uWJbws+lE4t5YWUBz88bFap56RU3M8DsdS//1kXayP06
pgny6Tm/4DYyaWobqTu6J2aRIz18iWwxDk9vxinYH2pPliAio5ACJ+LLXqg5+M8G
Voc6cPJ5GhTW6rikfNATtSMNO7McGjpFBtg5uYls9dIszfJswoYpcdirMVz9y6MB
q8YltLebANq5ZtGJeAnK9PSg1QteUnFrbGpXA5oSceiujURHbhBr09srqSeVDMHw
CnR/HKPMAQ/tK/zA+azXGwTEUp4mSer/M3btrsNez2xlf54PVdh4QQ7lxceZDFPV
fV7WRI2/fbccrZK0Uyt8CKDAkR6YAnwDmvIZQMvb8KwR7sbKTcpaUzDKuEF8/zzL
xAugY/h5kbg1KVGo1V1hZHcBMBPKJD4dPOz3S1/0VWedqXLh60wb2CUQOAgZ0qlX
z8ejUAv3RGXmpK2ii8BuVrylQO5o0huwusfrD6FvTwPIvwiXvLcmqHelPKowINHk
SebrgBxquFcrhz4eKv9kOIy8kCluWefY73msksCj9KhugfQuh+H1+20rP958j36x
mbUetQiUSY5DV1wksX5gfum+LuLloR9MRfcmYy0fT4nRcbLWM9ZLYaMuNAqCo/4y
G0pUq/yPaX5wgi4/wPVtSaNmyvX+f+Fw/K9Iy0R9foOqr+btPY8ipURZylNdq1Ve
nte8o90LuKYjFQrxj9ICK+q9xdP+NmWCGQuTh0O1Fyg0HyubBYzkRIC75Xlihe6Q
jLce26AOqo8L58cAGxF2ZFjFD9a1rdpKOSydKA+gUpLYWVnONkVsu3qTqG0q+30B
OOW7ApiFIf9hDmyWb0WUJ7i9Gn2j/hRrPGEAsk07CocYNKe6f/7T3ymf/HAJFwPX
fFXpnFB/+BWjhLTvYsbVrpWNf4PdaHA7Z1UbwKWCqD1Wx51UE0JkyJKF3pKFiuSo
AIe3x1qy1f3nztWR1HZSIkGGZDscqkq9j7QiY1H9S9HjZGx8al1epBC53EpccXp6
v5FvA2B4E3vqNqFx55/VckEuz6kYvDO8/UkPG71hFwm+pCS1g2H2bTH6y0ZsdmYt
HEbOpc+HHxBN6mJFsvjbI7RqU2O1s9eBXLnjlbncnifO5KOHpZQsMxw7Ru5a9FQF
1Cjrb1EZUyc8xIVtbjFghobfkHMzk1ZJtS8ovjXF5jrrUNYQAC6VyEJ636gmap4o
bxfZMmiVmy5e53P5b5N1NKf4M/1VPVtLe46C4LNmCXPLEC52v9Cd8q/AAw1TyWSr
Wn7UUz+YhWGdzjhg0+xB5l3IH2Y3UGshdKiwwxGJJ9s6CDkkky0huQrvxU1Gxv2L
O2DrI9iKYw8Qo12qjtTsL+CgjPxUfTLcZp8mA18vIVPqNg3Z0ywTOztab4i7ZceH
LtIlWdu8GOIUAnVRjjqNCqlzwxpGPuEv4ohnzgn9YryPySL/cJ/7LJ2bxqqIY5Nm
pxrO2c5D7dyRoBPovVBBNcf+a5IHtelywgL0XFpUfB+iDwNdzeHeel7J2W/dT4z4
v+cmIIydUfuAe/4xWqhz7IQ8Raj0kRQOIc54bZA6mlClk+eCH5gIZRFJCl9RpfUw
j0zjgNNlC5K8rXh6/y8aoivuz4/8Raw8muJXOVU2gKw2j1oLpjZ+9I9E2KdS2U/o
CL1rNJuh/4JgDWBYRGiZguzVlU+TxntzOLzuQ2+7sPqKD4vHAo4WSI03ny8CCp2L
uNzPoeDMdCk7NS+LjVjYd8C5NRoKhVcugDJMY+qn6ellXaEkDTuOn9NmjxOBmXHC
SrRpxXS5SV48mzdzlQWPlNyd65wTxEwBUZq8oP74ujkOYq2xvRECIfyt5gTAA2K3
VY9N6jd+QetjRWpIlFLzZwMzdOeJ/vfdSpGVOj4SetkNVT7tfA7SV9oknTlrJWLS
/Hl1kDDe5CuAfbLv2ftLljsPLNtF+RvM8umuuZdZk9E1nvqZHS60hKvdkuhajPG6
nlQut07HIxKEPfK9EFLR7623Ez2D0Eks1emtmZ65P60Iu2ldeXM5JYePhttUVQlw
lzzARGS26z6oU8saAUBzoGQR4dlRKQBbgDyrmTJZBHg1XFEVUvlYmoQw4CxVg/1S
UWVTSdU5pZumDfpgixQXG+4dGtFL9VqQFCieJxvZXGH7wAMh9Cl+/Ns9t1A1vINK
a11WE1JdmUh2cuKfIq2TKUxUSZMXRfKJORqSFBBDcEtLC284LXd0eOpXcd0v9DQS
6tt90g8AVCz4051C2226pSVpsbkvCXXAdczfJNBEYPvBuy6kNxVFFL5N6I8Qei+5
Bv7G/cFKIWfysx52t8G6eLsQbAMHVjnRgOA38e/TC7oRP0Ki9xXA/7WXlaVSwNWs
5vyaSVY0uRNy5m6g60r69JCT9CvdI0xo7GLOkraAD1p+LMRIFYvPivoMiYoyWYuZ
bivUGpzl5GaIjQBI8ASj34oMm6YYtkRMUUdx6qK61jjkKeZDpC4BNhnSFwEuC5Y7
zJLBrNDMHbG255nuw8FM9mpENKqUujt2oHwWJoA1M05Nh9uVK69jmgkQciU4TMdf
YN2MHj7psZsyIgr49kEmQpiB/afG36/m2/jmJkSmlICayciBAjtjsAuQ2NlrV6W3
Pz0sJ71OG9b4qHU1vPPUBo2PC/+FPI1hI6jp+fjdDjbOvLJz5ospHq+UMpJVl33x
E6HkINtMD/Zyix+7adk03CeTSA2asl+yaZeS9YMH5/5bOPuUMoWUqtZqU48oSyCN
DNBgMF0+eWvLkQXAeN2G1Ct2Vly720BJF6z+lT0q8uDpw6wNk3uvzqhVgs5IsZYP
7xYhbcwWBmE0U+bfeFn3FbFEPjkfa7oXsYJeGU/W8vQ06VmPmmvPhxC5CORvmIpP
kVzqCM1O0wmISihuOdv94SK9dDkNcPZP/YFmOyz0N7NnJzQlRdKzkTXuH9waXs3X
6J49/4NLz5372CClCoP/RTNOUCN39l1BbRBL06c4jeJGlvbAdq73S7JpD2xmWreJ
Nhx4YDGUjQ2g4RrziSCJUF8NOezihls1oBh0A59+LKCr+YAWPiJp7tFdLlox1xWg
0MQuxsqIXbLKqPyZNQMmODLQKymbM72LG/iUoreEQ/hSkA/HtFhH39O7mBQyv0Qw
Q22aUWvc7O4QDEGIczDOsvxIC1ynPOdKfSrsOM8TbhsHgw5CcxPrcuC2Pc1W8bTu
78AOAurbD7b3FzEHzgdhVfD+DoXI5FDnSXLCDG4yY8G+n3sESLU+pZxxX8vSRGX1
Jbr7clRn7SpIbdDPF8O4+nxMkxBCjBfOhMeczpC/rDd4LMPWOxBOp9Zqx2ZWwiZ1
xxbO7nR3GXGr/HQqZ7vWZAN5bilyOZGPia+J07bonksKZ40pMj3E5VD/36ui+9KU
N7mbpcYdXJW0dQZ+X8gluClB1S/2ow2HhsFVnNUkZmW9O6JViQfu09HK5PVLADod
9K5HhXBtAViYz4deo8Y16Ar4NTbUyuEPe6hdo0dorgDcGrnXlc7puuMJmS31DLjY
dtE75itclD+VF3pkkv7ItKAXdmsebJpNvoeP5Gm+je+7/leFpLA15pZBuisixRg5
dllSC0EE9txhPyRhrh3rnFs6osgSMquJjCyZwTvIHQed1GUADUwTz7MNXMg1aE6B
IQkGcV/atCQ+1E2IVqFjChsH6actzQmyH6CEXk6X1kjTBqDM94pSRb2T+mjTqmjT
HyFR8jCyNwI7KbNl5rqYYAKDlAayEVvP1H9mLYCfye90wvXG4nLedFPweIwZCd70
NGd0M6b5RrjxsZ0TJ51FamAtvYuJN1nwWhq8jaRch07bk9Jo3mRxrk446bgfG2YG
eaqYVyqaJksQGDepmO+3Ncc9txOCpPMP4VPWL9CaCyTRuUl1CM/x3GSuQ99yzXoi
EpqnW/AlwtcLNd8aaAb2SkJItF75uR3xglhwydDBeTj8cdZlh4g2o1W5wZq+kc2+
neLfMFB81s4HwmUmmdOyPQjUqbrcoKSpEdR6qcrfaOxH3hTc++HBdv822esA+zhI
beBTNxqPp7DtOaOEVTmTxDZwRSU/6BQkUPlCuVfkqLbbqgOsapFb0EQD0JdS3gUL
0U2iN85nGUQNAlQO6xNmzdxLJMMloLCJk3fWOOGGZ31XXwSVg+4r8hzfmGq65mJw
+ZrwN16YA7j2qSw+qOuyR794aeXzDKvwq99n4Ul1sL3GF/DLUtIND4njWT400FG5
q4teUSFVHfywjZhX8xGP0NlV1NFslqcdrMxfcC1pmPC/jPZb/NeG2bY1NXPoOcqr
vosHj8vkxXS+bKZ12PRuqU+3NhuqDfYD1c/vlqgfxJbo0vuf5H9fnNF2cFVY4Nh9
5dUAepAChHW+DO75AM7P+WetHS3rrVjgxXlHw51wda3BFaw7K1qRsOlpW/8AcSHk
MmY/Z6t8EWCgixDJW2uLeXqTq47KKBLEm1psqpYISZVU3A3zPSAhTTsnH8Gh7O3f
PfCPxE9oipF4b14gDbEtXNrX8wfTjx966wFr1Qdl+3N1DdXaRHeMoyaH0RiIu6uH
eEbyAMIKEBFxef1+Q7VBZcONoUXGJuqBluNoBD/VPsDcEHKzdprcMHx1UOOYuLDu
ctrin/nYnBzY7eAMVJAHBz01363hjfMzjWJ6/PvKwNVaNE1cGsleBIcNLmud2aIq
8mMhCD9yMHERN5n6PD742aUCgJxL5ilT5gnVKd/CzlQ8eDFoBA8/cM7CLYeDIV0H
ggm5PUgS8D/xewRTVIxnsdePae1qJlxuKqmyHPyYH7yp3KsmKNSpqNHvI3aJTcti
kw0ixkfRPHkovdxvZfvxHI92O0mTLZftxF9Q7MDA32MJwuy9X6YGy6HG6a02kgVQ
gZlWtAtsC4CrJ6u8oanxJ/XKFKlfKVwtLLNf6EqQhOku+nqQjYPl63UtVoFW4rs/
25dJ7eauFg84by3ScUnmX+8FXRoOC05mcJg+0uGtAykdqBIvUQLHsdbDV24MOJAn
Ou7K31ee2J+RFQRHmygn5kP1W9f4uxIOqzSb8cq8vTT8PlrynJBP4Spvp6NGGThX
pKdEjGbTl3uSVkZyH+/NPQe0K4vZz3xO2y09t116GRhsCQJRKq6+5e9Bp6ApuRUz
32DbvMXIpphfTEVDQ8LS/nR4VdyE9HXgKjSA7/jZu5RmzHt/Op4bDd9MzHQjEdjt
nAP0thwN769Vy/6r+ad/dyRjxIx0EYJMrJjX3b/YayfdzaGvx+0tP6syCkHn6o4X
UrS4aOTHcszWgwXvc52WqvLPZrXb7FtkRgC3hzXKW76Dii6GdvYjhh8ytIhUCD3s
lxwRjs2pAVTAn68qYohnodNvTAWl1iqwHCNKnUx4ae7hw9A/QLA692nEXi3u7b8i
DUZl/YMZpk2Kpfh6e07iEcX4ThaCu7TIftyeUV2rC6UC5re+qHEsdnLTzZo0jhI4
Zjtu5SqNzV9raiS/AkZGZn5dCDbolTP5faMKuXX7D/Zd/k29ypRBH0fosRYLRYoI
HDLfWdEfXaZpcAAbEiHDR5Ryy/YjARHomQkdSoXPDhCx7DPrTLSfUJKHkf1z64PB
0ojihaMwkrUDO4R+V2ekGRg6XPG7xgQAxU2GmKAi3WEdNLzaoVQttZwy6JAjJGA8
KGwFnXGWXkIxIifcsOSzhHU7nxM23lAtTruZmeew3/6vdI8tttPfWGAPFQ3Clmo6
fmikk/gyA64D5Gwybf977FdYSM4N+JrnrRA7EGmg/6yfEMDcWBcT4r/t3vBY0ccv
zMYk0Bglau7Obo9e5QUygtHkaYx32DJut6VxiUZsjm8BtwP8SIvdKDYmyJyjM1I2
CljaXwY/Utwbze49pr2PzisMXWRlcuJOifsQLXp/1EzLsKoiFYZdYXnlRZ8KbCld
fUzzdqhD91Zu7NPMPD5U+NRsmDpSR2QM05LsN087ocUlGFbEOb4k8Fz1j+D3jqTi
XOq0FGMxFuwo2Yd+y81slaxqJbRY5WypcPdrfnl+5iNOtX/tDYC598yz1UDm2LRY
hzXxq+dedCn1eevnulaBBDf0rO3ORfWf675fgeObWxTff3gH8PYZIpIT81lTsyDy
RB8wT9R6/LdQdPAreBiNVzCILyN3Gn4UspVSK//CGh8U+t8AwzhXj+pXzOAC5hxM
RZG9AKlitM5kcWFVBRQFGl4PmXHC251ERrSGxUZ3jmS+9RlU4JRSV+0Fs5VGoMnq
m8cOlNOCv5vfKT6JN1R8i11dpLiCE9E60hoTeSB+YhV7VFA7emluJGpT10HEmwmV
TWybSCAfFy3HhZ0o1Q3raIEKwJ/dpO15J49RHwfwHv5+p3/17Clm1d8ob/pkYKJc
/qdgDHNV+FLCx6L9wrSOtw8SxavcpauUjOIr2Rng6VTxqLfDyTHSwyEKcVfIia0o
gpS6MysCFBXOvy86j3toj1wKF5FTDBvSO7/TbK7RHcZ1JzVDbUaaY2DQVGEPR2+B
1Q9pA836B0ie6+1kU1MiF/PhHQuJMSwG1/mlkJCR9x7TpZ8S/3JvdLvW6p30Vw4M
Ssj9woLo7uIguknkdpHhEp9IniTulzFUqxU3ZPixQWg+AohtS1Az/qwQ+5hll96q
9//TpkBxaRlYWfQuU/KpbgYqV+ZpXZ/e6v3RKBhZ79XQ4cQWp/FyZGZ6hm62LTUr
5bI8Ne6y7WdGIjVkAhAWrtmZuQqpnrpOAwvWyYxKVeRatQ6iV0tCOR2puC11/RUY
q7/o5fyvdVpznwmTbSotNDvdTIQy2Rqo3jk5jK1fXDTwKsBo5xG1q6xcaw8yKLEH
woep1WV8Zw7v/PdGWL4xQw0hsBCJY1yrUE6P2RHZwsM4FZpLfoU60DkeIoLq/bMR
7EkluCsdJQplIE8BvF+Ak2WO5kSMefgfQTQivp1QX0ia3ajQf7oYozWH8w59zUZ6
MaJ2aWM0II9iMK/KexRaVQ9gID5xj++rE3B6CuMCfCXtf8PBTm8UxDmwWzB5L6Ye
R+hP/Hzg6Pjcb7vPuRt6XTDEJ4P0fkJNIgVA4bQYqRRxR9lWq/5wLLU9GrBR4caI
q21WDx18y0A8VjYloTsrXRH9/PKqTB/o9XlpDtND/EyuPreZnDkIN1W6WLHJlLmp
ELBa4B5Zrfurw+o3pfRYheX8mFhfkgQRIPfRjbHGMjXoytIpUgL10TEHJ8xhkJAR
5vjnDts8qm9YN6zCaCW39CuhY8Of+Fezham+y3YjEuGqxHsFN9JpyWoz/PF0g13E
FVk9i/TGrHxAF+MJ3lvefg==
`protect end_protected