`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12160 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
ZIICkMu+S2rq/yOQyqhpupmJ1IlVmAI52F7eUhB0KOSGuGyqtv6SFvqGPpIVAJdG
gHnsYaX5z6l4/EXxEHyv53+e25rg2CmOMevXkeLbpciLaU9mGVSRZj9KyOIza6lq
Mh44FUy87XDUCl/ZIrJKNEdalEpdupPY6kQlEwprPP87ZjRjRiiZBpnG3ojhz/V7
97+aNqqo/Jlaan0IWCBh2gfHuzB2wCXttrwvKkDTohAA3laHpQU//blrPVJLCEb0
BbXcXBXBDq51PqeE2rmSECaKcFj0+cJpwWGOLODapMyGuc0tiWCojJnSJJSxIM85
/ss0ZTPwu4BsC86rlSy+UVTalJUnC9hU216sLAyroz4MoUGaS9KQRqrL1wsGDEz2
kEJ+uqa6mNLnst6VdhcRTYvnJAi+s+cbZ7ZA8YmMbc9ktaLwkJT/ySqbfWdEo6K6
x24t6CHex4wSerh81gZc+w+0T0LWZzzkx9UNSXiLwcp584R2UqB59kc7/gOh4tzn
kfdvMEJTt/RgoUibzSpMiK/eE4g8NyNhERKZszDheP5gDr5NO+40ZMkKq26j/vrC
zW9SiPajoVR8CUAnszkvsgBfxWRZw3NMvB42RvzpkVwbYKVAgQG5ppQXPaeRfnCc
y0tVkV9ACcL/mr5qU4JyEcPrV0/Ko3c8K27ZbIcPZqcRMyyfC1S8k1+FzL8wEsdg
l4S3IlZxQpYdga0asLgJq6oYSObbvOwVEsDWL3dYOmIUwnXU4lxhiAirrcleSBpF
qHdhZyr9Qr2hZGG8TZQLnmLFDyjQBUgoUU7khAFf4z68yH/2VFDknZo5y+gDqpP5
6vysiu8aCma4NKWf0rbBnn1XlnhXG2X48cFSOSVVQ5ZwdiPzoLoSNtjvgQe+M+cc
6YKTRLx+vEdjOADT+nXagX0TNrYPXyP9nhMHj7uAvfNPOAVBcF2VUwG6Uql8GutT
jJb6ySI41k3yjJ9+psyR9zhXSz9axJEa+InRD3q8mo4EgXfP9cMhib4bMMMv0g3M
bpsnTbMNK1L0J8X/vmUruHz0kjpdBwduajEIn3puAB9WAHE+PHBDqWIr3Kyjubrl
QBDtjq84vf2QHmJdgFkFV8tdJ8wE3WSmNtRisHrGXyDzropjx8JX8OzIvy+8XXpG
IDUNc0HxecOOb+ClZ0Hzpu35PxnQTslS69gxj5C/hNZvSZ+o9AxRTXIYmM+O7+Rw
64VjSa8b60+8Mhqtn927ftAe3X3tRJn2NIW+X/A5gQLzTwH++Zvxhm3ykiNA1nfZ
vQTDZhc0CEujFsIVzBm8ap9jHeOkS21MTBRu9FCtN5hVP6cGZcmBX27/yHiJokXH
6zCJwRcTbnG2HGMW36NMAbPjfQYdc5hrlpuIajozMZpO8ma5uX2OKql+QAK59GvN
jfFQytTN/bqyC9gWq1ewOe2aC/WfJ5hCDgrCItM1eGpXUWkK7x3zc5nuIBRtm7Jy
D8uIQ0vjTdxCOskhvbCfEhibH25ZbPuaNigyY1OrL4XtGkz6wFZ+uWSmHRNj9AtF
rRdz4B1gdVugW1zFiqBGgxmxVm6zBazQ508VfkSaCU53bzKMzfi1AtUcM+kFXS3R
IqwsGCJ8h+c5tmBARuTiEQeCnRXA0ky2TxiZfQiB63XlU2aTZzrKKdzXLaTlSgfn
S8VgFNvpvn1X4w62li/ojVU7ir4RSLSNDWrEzxTZtrpZTnzzqfYUfGtEENY1vPqn
lGyAdixTZVgGyhJmUg9CBcRX60jPp3J4B1IfQu5tIL0C7V+UiPlIpGvFPGl3Lhj7
BGeXrCApbvPEsxxe4jMLDY9z3tG33NCZ2ZCAxC5yGI7EKXd8CzH+Puk7qTfeX4RY
+cKelCYpUQKr0tCPCNE8mHKn69nkltl+9mqRfqNVcYQfRBBInWGh8Ezm0RlS7BN5
PS8T5IkVvMpyDpK460AwUofloyieTZQAOx9PEloN0zOQX4wqKPKMck6oOVzanJVb
7AA3gRBANHdZTsk9uMPl8fUYdPw4ko8ucbCB4GNxaMJPMzuZBdAwcI7phnxRXxKN
3kQKdBDO/RqLQNpoxh91T19ezw96be+TvHJrZkfvqnYtXrtPlvqM3KGTGT/Dv7jj
EySH8ky5SAUOZUZVJP1RWzvPedhXLd05lXhhXV67BasgXOcKx1y1YEpLtxrzyJKN
ae5orMlBshkKYwFGTbg21td6LVDezktGK3L/83DJZ/EgEm5FwxdaAOP/6PSk8Ti0
HoVkcqqY3kMOxM7J/pdJ+So91jhcA96yOFUdLfOWhyYdH68W8A+oPaHXPLw8lS5E
w/RRnTebCvqScalsKLRTrfWZA9qOeAQRczWVZwnAKVu3mA4j2BU3n+t5KGnrZ/b7
+hn1LLNZQyqVfdG57L9nABAyzGK9dF4W/NA2ZdTgDqyusIyyzznHWfGpX+IAynt0
MHUISuXlXgvXLHc0gg+3qrvIh00Yspgsr7QZPqa2im1Oi7DyDMoxHbQ/e6p/dDap
a2D1i7WjbHOPkBXuzVZHGcCOH3dI0jhreEw+LWP4JqSRxZLErDQJx30sbNGi9it8
BvvZVchRjssTQmrsT+yYi/m3lPZXhYEpymklTDNaNxBNk1/fBUtrpRMpoeXjFXW6
tr5bAvMleeB5DOozupUcDUjuI+zCoylk16y9//bj7smwNQrfCVBtWYJ6bFbYF5kl
eslfFvLW5/45QG24S/TfUB6Q3RTQy/JDBh6w8lYPoEr5WCO9UWpl7zNmjVupMiD5
CaEjXiUwiArODDsUt5zck436jACTHhZiGShYzQqBaNnp4IDi6lYGIsTJnywSRc68
01Z7iCLrSZHov7GsqRDWpMcPX6+Brn5yJjUqvoq12myqvuMKWcRNfNFkikG0/8t2
DZS00UeKGPn3xhJIAcr6OpE1Arsa64gpsQjf3MFwvNPsn6H/NXSDDvyxT+Yd8sj8
d5vJDNLRYMRFs/8o/99DAOscQ1u4gVrlGcQi9DziXfLagx4t5aNLHHR3XTnCVJ18
1M6ekUEOKwNbJbVlVi5xoMZArfHj8ubmpIHqRh0qaE2LBmkwtiSyYhX8w7t27kO5
zuAPFK4AB7D1UXpvm/bzjRftAQt2ve7GxOaxxsOeTYVlyMwhHClEqUXqVGai23wp
U6XEVAlO754xkZtbWbxBdsIDM1tpxXc0cfC2tZaNrZAaxu7KYz1PJDGKLx02etzn
PqpqyZWNp3q7CyvFYB//9P1BYwbpgUmfkWYjjtDLHSxyf7NCYV8P7kxlW3VdvemS
uWS3GHdSqHFvNy3IOjPR2CpnLRrTo6ZZp0v/7CpL55lhISAazEwnh/vfxfyYimak
dh8iUQbRyGalIjaMjrIvldNAE1KE6uz2Rm3Oc1zkQszoybEVks9TMphAOcWbIUiw
qOTVHjQPhEFVOc+OvQWeIjbQq4rPbLOzbooGOyQYeBkreD5rPfxix9PbNMVEbN7X
6jh/65NlMUs+IHTl8dQu/hiDP1PMgowr+4v68i17Vxak2ZKJBSLkBZhlEBGQicA+
tk1obctYCRAqs89t0kLFmMpdI6haCtQ4htQaSVkeS4JX1gpMPWB+qbn0TyF/S6Kz
4c+rcY7YHi+JburG5M0zzKWBiwffMGFH5kFr7gEu81geayAxK6366GDl/Ug4zuTW
8kcB0b1nkAGyH8guKtpFwWjBmvuXj9chp3WMI1dGfPF9QyhXKVfbD9LoAnUphKkc
NmTiLpCV6DhHTVC6i98wzNbr0BOJ2fKqAwjzVnkoSnPYeSJUUzaeHEu1CKi8111Q
hGIShtynwiYYHmWGQH7qPeedQc9cJ8BCphRTo8SEDpp7vMceYSwZZUu8akgBs33K
MgiTW3SgNdcmrfEUac+WE5yEvaPvcRqdQggzx+ZH7LTfKPVKelMgvf6sEBvH3VPP
+5jliin4Tg6FamO2Tlk5ieg8KxrAPaE9RHXgdkpxV/gxbnb86ZjP3Ek2OA0TIGIR
ud71qFjltEWvTQry7utsfyvmmdqvIrFRWuesGADTT+y1mHhFH+zMvNFrluHntLwp
nQR+EUS6IKjd5/+ruL4E0SohD1AfHhIDXyKsPrP51/HeblI5xWHswptFCoLaMRME
meRckiA7j/3Hraty5FAQZhJ0Vo4QFL60Gz5EA48qUknxqsSj3mtc0mLS39jbcMYH
UK+lFxJ5/c8adQwxUjRnpvRuBB/+dpvShrvH3vf/dmlOXeH5Nryvueltb94yEfke
qA7rLqc/cM9QSdu5dnl/ipsJsWWyfCk+TixNraC3mtTV2UWnC1aKfH4xV5eNIAF+
TGavNmKFRc4a2DylY2p7EJfgszJ+dA5XHLouMENnqrVoImcprTMfHCn4Yd/Ltd13
pCpAXMbTHCBpeCn568BHXVYi96ZGCPjUi3IFQNhSuxBKFfCHWOoMCqopLVIRC9Pf
Z7pAyJL+hSpqZOG/TuAmblGc7blOuISubEcmW8yJ4tbKRJmZutGgUBDwx1WZvejE
4As80JdW3bDv4dwGPcDLASaQpzBCz+d3svfNClLE0Gu0/5hdpNeq0pp1f7BKtUKo
zQJ3C1AaRCNZ9MnqWVfF3Q4tjCSG/NcoHBZf/mLZO/W0DhLlPhdd0KG64LgU0Ps9
PZTzRQhjK24+8chyrkFxS7kHFW4SEHr1vczAoMj9HDbjmvKFr8p0rSnnPwWT+/MO
9WowcnyRdA6zpE0+jqz+0zYVtkVGotkBDbyTNfVtUC6Z0eVZNIlOcm0A3feTucXz
fFS2NJRoBKdHSjWG/MxjXRkAX7epL2JHFQGikiiB5Xd3dVK5+A3a7D3twA1duE2X
ELLHxUX5UKLqyz46TxTtUwIMc6il9d1QfKusDoRg55yzhb0YbiKwoHWHyV2m0OYi
OFOuy2EhNDX34TyawYjn7eFFwdzgIK7DgZRwWdiyWQkjWXq1ZDOgWaQiY02KEjBX
j2LujTXRnzWYfqx5B/q6l9ysQu0kgkHZZ+GoJMaxZreE7vDhHh2WZQEceRNY/Mfy
kR9n1JJRWsvp9eACzQtVuiqClOZxnpDgt/+eWsIhDdk+HA94cXsd/KZ4aRcQAdZu
4co1lQ0ozPGVXdH2FEuHytdJb8Tb08nqQery5fQEp+2gbs1TZBG2htpxOWms9QPV
kg56IJ+TRRgSGbFkM6tLMzjoKYXlTkwJ4eQhGSmcwTx5Pw2XzsSq1uFj0DROEOgQ
ToSruC7ipMbYm1q74taGEM/nYk3xToDuG1fZ3PVt6+LcxBDQRuGrjrcV87HoqgJh
kg4Zo1r1H1kVUAEbWomxekTnsQz7bV0l0Swqqw422586SI0rY4QrVvgSVxaA2NSX
gxgAteP/81cV+pv1l8/j1v1/rQIusD8s5/zdSRD7hfRLfPrxhnOiMz59/8OoSCc4
4mGKHPb1e7Xi71z5jn82UObRw6K/xNQnD1Hl/gYpT//1XEgFBpIrRglMOl0OuXqw
xxq8uRzys0HmUDAxf4hoLVlhvciUnVF24ASFVFMMh4RyQB84baZob67v7jlL9Pu0
B3M0ga9ym8H4SHucFMjeve6jiialUaXcKz87O7Jaxd+5rG4FyhI1Ws46Tg3uU7Ff
0GT+rj5qxzH1tY5mQIZX4h6pGg+V+/BHnP2BcgTp9rQ+3bapTuzSNsB3pHmacSpF
h2JXYvtFdKuwdOh00fyzXQBLNmlLsZUspqzoYjPo/vyJ2uMIyCI0LFEKmcwV2aGV
0O+2NWiQ8fkp68BbmnoO0+edCGNCLuisp5J7z2CGC2dFDEGa4yItsLpD3NT4UyAI
veIZkHDvRNTeLECEx+C4Iog6AtCto4JQ+eIfjn/q3A+jliokk4dzpw08hAtM/OQ8
Ja/kjdCfgNVRAsw+DoOqIwtisrK9I024w7Yue65f7Qu/B6sdylGX0aSkIllEl3kl
CG72jSY8q7H3riSE5eW4zQUdRbnEfe5/dwep/BWIDuytda36zM5OYboUyv9+JM5E
VcIWfPuftShs1vknsLUhLmERM93tG5DWyk9PbJj9wxBfzf+U+afVsl6FiBiDAILl
qmJFbiGmFjrn/wA4TrV1Sh0k5VLZqSO03hH7CwxBolgh3UjuScjel0sxaZOqZMwD
qP7vMBIB1K+dcSxBGccBdGFhYUU65vgmv0oCcIBDPk2hNyjpiyCixrgZZ1c6tMuE
45lBMvgFTj+lLFY8BQbRrSrzODnMELxMuwVABNtgI2Mhd1pVm1kSq8+BO50pfD8J
aKgiN9x7niiJNonfSfy2iCcqy0ifJ2Bn5K1EAlQP4BimbIC7Yk0bGqkWKG+5Ndtb
hkhFp2p1Vk6j/ZsesU/RuxFrILzG9aPj4OrFH+hkj4QpZP7oQJla395EzjAxmmue
eXA7/uEQOoQJlhOLLy0HLmFuIATM9v31F+SJTvD0aBO+6fs8HcGC4rujFwGOuYkE
JSvTVcTywgjwpYTQPm8jbd+iN78O6Ity9u24XmF/GpKrl7AEIi9zl8L5ZpYbGFRG
hbnv+1SVH9JSM7Tm1bMkTxNBnmjTcealJn1WZmwT/k8rDwwfDYXQMBdghcegSN0N
3aJUO/3OrpzlKIC0T+8C/7WC4rhjMmT3G9RNarzhxNmf+fjY5G27jg288xcGUvqs
/P+Utl7inRpL3AZb59Pxf26Rde5mZUzQ5/6qrt9GUyUq2TSW1GzDlA+2WhnmlGkK
6TvhleqbizuiirH+Vk1nxQMuyZygemET89j5Ve8QbkfYg92+I4UptRkafMpnQYos
pfdlieLXfmvQV6aONCVlEEvqijeY+LeUubsAV82iG26BlK8JKkpL2jMwZUXCH26N
HfrZ0CvAPeXEMGEEzPV4uYuuJWKWg1sj7dBL6b0KEZ4/6tlK4aiKm2wqh72iaiR5
eYW80sI8F3Nyl7bnKFY8a9AaTzALUlhtDdx9+qEn+uiWb79DXs58TRizD0dt3arI
cJSyVlbc0jNho2TjtdO8qVhF6RVJtMaD4oOsp4yFlCpfwK2Cj5DSnMuVLSFx8dgv
0h6I9WeJjN2fNhDB1Fgy3VyzdSye96e/fZ1fu3w6iDebxeryuIbm551M9wWJdkVU
fqxeFF9FVYHBTAOaBZDXUCi7bgBKzeEFKUcy6yNrmdNji7zOgddrEHF13wIX9h7V
WL0rHc7K6sjg+j785RthmuvuJEuFQA5+3Rs986N2oXh5wl4uwXDGxr1DpknM4NLP
Uup9+jfnuyGf0ve5J9cFiQrPQvpE/egbISIxEQrHZhPATGuVNzpshVCkCLpULvPi
9c37YnMUFT0hLsDLc1GDC5LF2eESZaNxwLL/sZuu3GlS3nT+vbNv++meCfasyQy3
XDfy18sc6LxLys9j41+tLsM94Z6LkeNql1uOZnjBaJuq0zcXo+OXGwyVnRy0A6fM
1MNXM6i8Ryf2Sf1FD7kgn8oqE/nFNVPoXpBON1mw1iyxKkx2zuyIZblUCZtjPush
/UP7qA0bYHyjgrxMNbHf+i1RMB1em23UYN1YbBIOzm2JPsYXlDeTWrNw0s34LKm4
NLyq6Zl/sWqmBo0NWlnli5QBaVxJFxydvT7Rz9VR+0nO8+jPLlk5qujOujuCGXVx
hV/461roFG/rYxlnPGhHJkVjkHSZ9nfoAkFmQcb2kPeLIhoaqCoyz8MRwXZr2vbU
mefFLOwJgbIeppH7lQ0039LQOI/R3ZBeSx94JUumFGoke2j6HpShx97xWoJXsLhI
2Vk0D81/W4ju8tybd19jq9O0fmZI2zRfxJ/c22cMyxPis8eTimN5xSd/pyN6LpcJ
PFD//ssSqTB7pQYIWIrLM2rK8GnzHbgrpMK/bi9Mp3zfkwTcOqunk88ujeqoYTVF
csAfKgJ5R6I7K2Wz8KKfEOdQE1rPJUVo2vF7kq/ii7QgLMugKp1uR+yR7ugzTSle
RY2QuvqBLU3lNH9TMe24RSaJuI+Iqjh77QWu4nYrLXTnC0XQTTwK5wnQdGOevRmo
024pkCu5nXGl4b5iGqsZchDVoHugmpEGqR2ERe2OdhMRpGrq7xkgTZ3aitq+5jPV
iFpgtvg+GK/izQV+/DhMPhgBFbYl/ovzqA/SVqs9mJWnZ4Cd1Md0SCXm4mHVqvGj
BJjcGOSSV4lTlorHi2PDO2aBX4IOyDYRV45Ofpp8bhDQNud3YxIe//jHdWBzuz2c
r5+fQlUQ9jEQZcMRcZ3x7zcd7VSwYfb9yN3jq26gMGRfiXJ9Tzj3rfbr6Zt2DHxv
YX6mSzvq+zrQFxBlo4lOB7teHY/TBKOd8L4Y5udkIWNbHj/6HYwCmZu5s8PenSXn
gxHj5/6iGCr+OYqF1KFK1xqdy9IikkD9XMX4Yl2AlUGW4nC25U8MJExYipYoMdeQ
0CPHbtHaPcdPt81VBkndxc16WfC9YIb9QAg7xv8CMdqaSm8s5JavQvKrsgFXk5ud
KJ6OssP8yPajIGOLmFGDRb9/FpuKUVrtd8bR4UzsZT6S30cTVThInjvCjl6PausH
sCH+q+zhc/z/G8908PRhGRP4Qj3Vq6pGcDSfQbXE3KzJZzOH8P2kLFflYGM3EOTJ
HE0kYA85A0BGjPFpMr8EAAzIV3dxRuPVUVzGgwZ8gzQ7iTuZmsaH453zfxdyrOkx
Rl6w1bLnH09GtFmP/5bocbR5mcTd8Gqd/K0ajH6VtCko4rcEPOR5U77z6Z4AMoJd
gGqASDMQT2cIcYYX8poqYUlAjib0QHYOUjU/4ByjvQ54CYybgu4EHyYp3klcY3BY
ZxzHE8We/ErzXuF6bgHMcq4y6bH7kSwOasOH/eMXw6re/KhxFngDfjzit6fXbXzf
6zxiPGfvBrzowaP7yrVAqhd18l2fLITrin7tXCxWAxS51KVVkP7gr2XhIlUd+JYb
9eP8kyI/hc+FxRnoHK0AT7QbuYWoyJLNO6bJK3EbGPKNn9Uv3bvkuqUGBuWJ3LjA
lQIlFayJRR501jiBwTdbQbfbZsdTYow5nCcryQfA+Gl8uGaeaGedCAW390CMjZ2F
C4uMTn6GB5BCKttFUE20q/VNgqLl2jH33BrajJPjpNZ6JTYXTghIAjvzUxUpL2Rc
akIcu6w946rOx2t4r/1KFfFEl1FeJieIyiGl5pzGVc4ROQy6UcUDBqBbEzoiodky
3bs+aV8bsC5PVBbkdfmi67nsiRy6qT5s2f4/ZhFiIFfj8rFfvoxcr1LS+YunFeUA
0PLnlgKxXkGumITrQgsbu+fXDHVOGQS6qjah6l71vBrPUvI0Eb6oHyqChIAYe1AC
s4CqBFj5orGdzBJb0CjLHq1LU7FdeTioWhKOLgdQ5tfg1PQ5ZlOE7WI9cv5/D1KP
ESByT1yHhNd6gedNI8fM69lA3B1wlZWs+EtraryXAVNGnKfz+svvsGZcMDR65h7A
RzDlk9j74c4PmTPWbdB7ikJUZ9tU5m5i0sZMYC1cpTeCPEHIe8W3asp86uTKawZA
c+lrbJTXxvyvKdqwNMSR2HnNsiA098B205sTzRy1sTMeXwkok/szqdHq5AyQSA5n
W52OOJPSpUU1337Mmf79lD/1F3xEPY4yffMLkrTEcjDVX3O71jigPbxJ3crNB0JL
rEoSPrqJ6aJuyFFuSu356qNX30b+B0xuwc0eUYsuAith+flsYLJqW6mWE/ATzvwV
4O1rZpZ/LYpjoTL46FqH+tfKNFgp83rcvkd/+8fkqSqoUIBk+PsKvpDjzG5u27/c
LknsPBnfo1GfHOQpGl/bX163HMwxAdm9wjvJLNnTFyDt243oldsRo1E3S4seXzVh
krFA+RS98PRprsTdBuNW0IyOGCsjgWvgKSdlWmPqeOn+/N2QNTp2os4e3/dpxI+l
DyAUvzq66Gu2ITGwhakEm1/E86TmNN3M0dawUW3tHefKaHIx4WUFiTFkWVeFIzEt
hC+y0/3bzMzc2ZAywRu6MNKZc+OBr1ihlXNhYBYhwgdxN2aChMqPEDTsmSO3A0+a
2t8fyE5rGzcB2/SBhS0EbMVU768VzuJ/a7GDdB83vJN486TAWiVIc9NO2DW+cacv
K7DZuw85On2KLwelnCpjt7sQBXO6PLu5kG0+McNYF+2hrZC+QWR9yAL7Ru8GBsd/
FQkk/aUiKKsoNHkFnvTaAXtgornAxlUAomXEvCb/9yKjAsrhfdIZhC5/4O0FJhox
pdUGa8S6wa73jhXSgPlhlzo6zekENF/PMeOY5vdfWf9gsm9FIs1y+ibnONKbXuX+
juP2OCjcldqh4de2RJ0c0afWjHYXpwU3LpYWDyXzFgGZAzWwws2AE3exGrGeGOVj
QgHpusxik1y2+rjg5eBBC26t90qi+uSjQPl3awKjs00DC74u82mGC2g0rt5Nf07v
9e38j/hzT/HrF4XoTE/IlDawg6AZ7c1BVD+7BhjQFwaSu5fr6UMWms4AAGwXL3mg
xwk+ZJubIJ/b6mTwyREq5b/h47nHbmwt/3R+LOC7Rc5IZIp7iG2LbLKO+rS/7pVt
NKVl4k+Tre7yHBCAJ5PBltdHJEjxHI+pJn0Fs9EYCP88eNzcSxWLdIR9wcT2Lj5u
sZTljj6h+7DWfBTQhoPxxCtg51dJ4K3FbsxfO8Qc/Y38NhS0T/i6oRC9Mg+SI3wU
w/DnavuXy8z1s8pCmLMTXJYhXWlC0HW+dDi0vosMuwBNF2a1B7AsJHZrh8o0ozq/
q9NHK0Q1OjcmXDJ8PMGjXUiLkNl/P4LG7POGJ7ayx6FIB/mTmoAWJmSf9g3cpYrI
CzSXTHSlw/R7mbR//DM7E5WbtkvcOu1gp2/dKK+Z+ugMzlx3nbk0g8XgvmUfCb87
89XzYsYZfPgDr1JFknrAppslPi7nOzVZTgTqJChmHbIWA+bzew19YmPUF8ujAhOI
WUbcKqLwwUGYLgv4mQXEq73IISb8trsMRriXSuJYG89fKaJTX8onSwYqrnmS4Qqf
f3/H/CbBR69rHbAiGD/H4t8E0AMjuLVfKEUvgF5akXyTpi/dc78Cphelu7HRWI07
ZXubCD7KZ6LD8RZ0RPnKJX/3N1lLheU1EtHhgFz5+GjNK6B7qdEHH71EtuHzl80f
cdhQueH68L2J1nIa2APdSKM8jblLHWX0WnNUI/yXrKxCfpRpDxqvkinL+Go8bsAd
YLGPM2iXgkgNrhtoCTfRo7QBiFzEL9ZhfUkcMQDujdrtLdPuOmpW5pHfXkh5BJtW
ydgpoSnlFaL6ga14jjov8xEwTXJjWVzHrbhErAlrdvw2ZoeylFvCM88EE322G2T0
UeBxaf/ggEtsXCMhJBAx+gY7dGsctjFT8Q3PYAxgFrA0y4Jr87FhkoGxC/ej38ZQ
E4c1MOWj15KMqJGWHr2hhQviigz6xzcT8eYmFB4i2E500GT/pE+h2E3VO2smMa4p
1YnHxxOTH9+VxgpyXbk2uV7Fx/7OgrnvLgf4oXLhajt/DlalYlMvzBDe5ytyfX3A
dsEjXhIph1xWL6P8qWehdTcNBa/IDMxuorlFKn63/la5BQYKyj83lc/7Hj76fliF
35KAKpRYervfJvMOKvYFHhUG4SukcPDRTSYqMSSx+N9uM9KksFJyOJqOGryfV38f
wxTwL6bFeWdoJ6i1GjwfpAykxQkI77HTcjJrGt65s8h4LVaNseJU00TwegUQ86gs
lGOaWf8DeR25cKKNvRz/lqcPOVvOBE+GSuhn7zIep8cVXnOmHcXrXF79ISa/ialo
sP18WHWbBCVt17g2qB2ErCfcd69+j0Y2MBz86c0fljmIIq3Edps72KqD6A6OY2Y9
3ZB9cXqYnzFqwhtNgzQCTyWyhxEjLes8XetKkfVccp3uQ4ZaclOciC/Jdu/KoXJR
8cjRyb88Gz3SumRKLEtMAJXj5Gp+0ut7t8Rx0kpnGKsXAYokd5hWJL25SfPAy8ky
S8Lu/Ht+lqX+QTLDoof4KK05HuMunuHapIAaBK9KKpRodYcVasLSUDgbYEMjvPTC
4FRI3Em+UvV1Bjz5tPgtfROZWUy8nZs8xQTFqDX78DC/zR+r0s79hMia1aOpm/kE
oIAUkmiNdVfVd5DW5amjcI/QU8/JtGa08ZWIdsSBOg4HFKy4Jnvv2TvHmnePt45b
EAh0x60dAGmsivolgjKQGfUTnawNqIIcGMoa7lHyVWP1psiC0KOtO6Q0B9A+P8sl
v3LbI/3LJOG7B52y7IGqTDk08pQkp2ljVTq8ph41kXExumlxzDxaFREM63pxvY+C
HGfE/yWJRxXSKv7yJTqWEtMj6iqb45B4QsG7rKMzTxhfC2fnZgE7q4OkPniePayo
pH+/79TbBAS4NKoBCiWoVelN92FrxtuJxahY8T7EgH+ggkhvoYhC7TgGABdku1CV
12hfEk1qEOWrWK2As23IakGdOpDB0l1Gm00QkEVTEvEqXFebTlCu70+uWB8Q+1Rx
e9D8zyoMnOzqFbV8jZXG0ZugL/qTFU2noqGPoUarzh/PWEgIAWOIC1/WWK6rhBlA
Zcdiz6RLmZEc7bCQHRTThuQJVtKfCEUryTImg9L9gA05yCL5mqJxRFGp/BEUGApF
wIVPw6qOJU+/yW5Cxt+7cIZspUMncp6efC2XxTZKMw2BRJCf8AVRawVMTJNsOEt9
srB9ggdAGP3RGtlWtLFPf84M3aq9tTgQedO37bIg+hY5YLWe+0qO02sLfNoMvK7t
HmG1gqUXx6o2HE7r4HSYzn5y1Qj8oMya2M1MJ/HTazEWGhsRWLGy6TWWylvcw96U
v0/uyIHp/pNf2gvYv9PRXxvTaPLlaqG4oOgM3KI2NbK67Z6YtXbOb2wOWZ1eruc9
u21dSDB+rkQS+JBg2EShJBWXM2RkCUBHMKxD5ZVfmY+XItJIBMJmtt3knXrb7LUE
mtaze55C1ds/xYwAzg7NRuFKeB8VJFYnJ9ZQJ+cXFRmftya6hPWzlpEZZ4XYlVrs
z2k95DeE9DaXGLnlvq8VluAQtjx/yELXesYyBmQk3S0u35wCEf2vzYFFbWAJBAfu
UJGCMtYT6A9b2VyT6LJ2c0qeNRM+02wR8nV9niCqGOErSRXzSSibRcc+Ly6wmCnT
fQhRtpgPuNHDCoXxRM4R8BdKAtJwWFk8nO6+ZNmLgevIPcFBEFmEHzQEGPsiIGPk
n3PXqxqaGaWpM/ihf0F+MeXFj9oY9QQlusODgeefG9bGzojs6d++QmRpDiOBBT2T
SQuoz5pogulw4Ne5Rmns+Otdtu6V761clyIMH2Zkb+rPKm+wacMRhp3RML/tGoNb
dVvrWvyItcDXOpF33H1iUNk9YNJMHv2YqQwIeKlctEEU0HAx+7b7m9M9CseDKdN+
LVGHtfjr/X3e3P2sHYiXR0AngpktUNlb5Gzq9BiRce1r/DYNn38X+8ZzBDvLOSLA
Tqpj2Yo40MWtmcxE0VJcnCB6QWvYu/yyDpXsuAaMgmymPG8g8imAjcdkJohzxGFM
cuZBhwHFWEefi4X5ZqKjV0zcuggyNFEYyQErJUHhDHYPivBfgjV385vajkhYby2m
AI3rbEQGVjdfKVDbl3z/OGS3KiQ7Dq3WxiRlhVtBHHDIeLMBbYiJ6elGO+ZwI+8W
yyVhZQP43u+UYpt9VNrvzBNRd1UmsvuOC6zoypgXU+AlPacXJZQB4ceHR65rPr6W
7cGHnHBCIkfB2ltKiaJQozWmRGdwX1X32PMQqr/MvMF6ofJ0vkJI16pjIuIzcEpk
zdFDuUs7gYPPb0zdUuGaPLJJnTbmUK2URfmN185ANb9xucx72QmP381SAUcrwB3m
GhGPFzZ2wLJICJs7+wHZnXvzWnXupwRYf6rIkQBMXybibil61oW+mfeFPz0UcU+Y
yJwc717Ygf3arb9dbvk9a81OapqOxB0DfqoFlMQY1fmpNxVFhpfUwcifkgvdmg1M
autK358c7ynk9mXG6NoqK6p19aWnoAQj3JkCEy7S3OpSso/6r8SuwTKfCscMVViZ
LZ/qXHg+O+l0aeUBtAJs8zciEqVocVB9vxVU8uU2IZuogBM3Rl04x0s7WEg/Y+Z7
zOmGE13enm5GA5YkQpAfsyGDG12jRcOUPuJZb3l9Cgcgzz2f6DMQC3QZT/xrnwOq
A1P45fOYgCCkbb7kCKIHYk47jONQu+wxfvFGmhKH6liw7cu4GI/+j/gEsQLHxH5x
XaI8AG9l4VR786ZG68cIIpJNXSkyVjFUrtXvSboPYakEq0/rrrbul9im7IbWPGSJ
X/Ij5yRpv/WT9WStyU94hYsYkpQ4WIkxJMVREDPylv1owZLlTM04hvKg7e5COnwl
EU8e3uNLRBzGu1WWycCUw4TVjsn4LMTTztmWHZqYYooy/IjM16NHyx/9tjTWMOvD
3ZVeX+ZAvtWMQc6D84dfmaW+CKz4CJYE8qVQAzLnbugIAbOjqEnZCn9uXXdV+RfD
eXz6fjPfndM0ddtUUzgD2o+YiHRJ8SpUTcMqtjlLlhJrC7M1gADC+Jh3Qu0t24+f
XRaTlQKz9aF3YZjOhgx3Wp3oohLOeLEF6E+u96MF9+xnoGe8G2802qbMkAhyT3k+
6fzDlM1CgSMmFzJb+fowvQmprAaoeQfXgIpOvyJFg9ScoDrAgGE/g2Uah46zb0iY
iGYREDRwrggP8T43oRBd6c94lkGZT3Zo4QQYsHqfItfWpS6y2AIWkzCnsWykrQZm
zsN2LzvWR8Fth7beGEMuQLNM7Y0Zifb/dYAY3kmFyKDgO71WtexsXoY5uIrlX1Im
OdiXqe9GJ0ceN/n+NV4yGvvUzdMAWTh07cQFseEqfNHKlzJHYffDYspe8yRnHw9G
pP+x3LVe+18TQH7+ubWz7pzVODrQ5ilMtoUW7Z/5TBsWJ8OcF7fpAaTteQjVDqcp
7LQFSAd5csjoCRnEq4W6O1UEzgLA65+QuL7em/HtWWXz5S/zZAaH7ejcDUShLwFh
jrnK33rnBdt+jVx6LQIzZbL4r5TqWHIoFn1ci6CH7V2rm3PQEJPMHqO7kTleAUI+
ZM9MOnLcfpJrZhz1/OBtrBfNdZr4YzGUVjxeaOG9EC3YTuIa1JTsMBvKGGC9PlaJ
7kaXE24jEZbUdE+XOOen6cuRMAcl33XVl/3XLXAkgOPB8TQM+GdgCHm6Eqx29Ysp
Qlltpt+E0bdVNIl5k+NmB7lipLO7by7Tv+lHMOCi8xrBh5TQg/FlSwL2ZqOnwgGz
wCuw97x821Z33sEOh3cjw+TFiEsAfOgoE76XAtVcrARdj/16DA1NtI+4UHLZbz6m
YIfUsw88EEqt1ljiVy/mNsmJnrqcReSvR0NME0DLOaZepAUqGzsCsddbGQoY0VDm
xpZ3v2Q5dsbF2Ii0RyaDH6atS+MrXKv2HaSKsoRuSNfrE9qcbrn1sF9/tNoP9glS
nkCoasRW7jaleloAweH/mgohMaKYEMslETm1QSCqDouneUsMI4FvrnwFofgFuS+U
oYrbje4ZfHTgbF2sik7Nc2InLviKl+ShjSyBdRQDcgL0q397jjUuroWdvANABB9Y
uQpD3Wzjj5EfY7SJZzavoSwGAOCCpHHU1D3Jn6/m2s4hMC2TYXSC2JglpzJlaUqa
cxuKzMc2A/cuJjcU4P0XJLc8UfVjeHox31zqFBLtdIMGOmbeR/29DVvIB/e2x+9O
/8INJteU2rAevHyjx1NW3mPvCTDM/i8iaVobSnCEOzoFoLf6kUco28bnrK9/J7aa
B4mOjs9voNYP+JJdaiNcaPVCGGQAmIFu146WG6ajO1lwvyUc63Nm583I8SujVEIr
HW79ioI9+WCLQVgdQsOg5qIIkViyp73TiQEjWsD7gHWfM+hhYF5cbPYDbiBQqCep
E0dPKYUCL9cL+n4rwBMjKKx/nLyedogvKXI3t38/v5tpbrXJauXUFEhqDfC5dXs+
bV9YECNjs/lHlvzxU+vJwseYa4kSn9B/wR7VypVEowrsIoCeS+fsettlGiOQXYBy
+se0nB+ihbJEfjMMmasyTR8CkMnQbOhx6YERCjqE+XVhY6BqVRZwAEo+FPgIE8wl
t7QJJ6oys0F7YauRGpf96cCY7KvHkGXDB5D2iDcTTwvSJqAM9uyAaScmVzDPnFQB
Kgk/MCmvi3wHZarA+FUngsi7qdespP5KPCcGAlzT5QNmOjWdywccjIs3Xvd1d4aM
YVu2pQeL9vcSMMQwLpGzyg==
`protect end_protected