`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 50560 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
GgG2UXwpbWAyDgGIJC8iiEUFn71cG1bxQH2TmDv1l4sf7RKD67pmA9S7ibKAUnnn
A9PvL0+WAAIcPNcki0ZLjziZTc7Gi2noUKZcGPrU/j/k0VBbOConxruBuEbu093v
Xa34gSM8WsUmb/6vSF3CGqqMgn8/sd+ZhTZtSR96RvpnRob7c2S269o0BvX5L1Ji
1Q9R5DjT5H7fSRGaCrVsAmPM+1rPvxfEpiyTGrBlpRXj8iScifkpmmVrjLVMRmu9
sgT0LZmdZbKnyifooyMmZ6L6Ukt8ma0xVAZWBZbZ+wZ9SrGr70Ndu7pWPK4MF5zK
PQjF3+A/9KO5u6PcYct5w5qNLTtslvu0HrXg1mpJ4qJO4jfZ+CIbNDvNzky6Zjwz
z9mvoCD9VYw85ACJu+RFJRf+Vyc6EptPjl/8CASZsWiq7aTOYUU2kuo/hNHp7B3c
kNqW+yEWzE2DfUFOyz61upRrxqDlr3yPUPRyBgE0xMXncIfXOO1AAXT2ynybznwF
p+oPIncBVcQuWJjeFwGG75A8HjAF76mKpRtsyKFmKVvwt/09WvwRw0cS3gvI6VIH
s28kK7nkbh6RqrJQzItcizLcCswjy6AkgPh/FNJhCoi88pTkPXalSs4f/W2ZXA1L
Kvd56DceAcTFR9loOgWol4YuRUVvRfMW7sn29od8pLSCvG12NMcJpqyWMOdooQbB
48IUVt7Yx3fYBPhjLZJnV9ujfrkFyCWSK8c93pjvhUyYrsCUXyyVX9hPhZb1qTNA
WTtNjzx0CIM4EvAHCRmFTZTxEtX5qLJWauEkLEL6x5kKR/XOjexyY5XhLLRaD3ol
Yc/gQA/AdC1Dz86JSXD9G8C3do79kHr1LSihVrWrA3qbFP+iQfexrZzvxKfapnhA
PzAVWRGbMxVPKkTBlXemRLBsQBbmlrdcMtix0z8SAKRZ1fuKzoN+7rfnAmGIKu3I
CrAVv+O7GUafGsQNnOFXn7OunrFtaAQgEv+vH3t5jjVH75gIF6K5Li0mU3UNjoYh
77O+rBxK5RyeYASRlw7zQjpH5HaBQjZd9po9Mcy9MFdMDufU0e9lMGTZMTCoaH2O
niFA+5ydW8Eh9G11YN34fM8mXjRbEwDYe1a93ii2teJjUeeCkPf036QPPte0bdeI
cwzMVHLCRDugtsDrG+5UpiufRSztCxBJZ1oYo/iuBo2DhwhMK9HFrcpu+XNnw4mM
cD4w5GhHxOByNMO52QhOUniFWdFZTsnM1J/5xhOglm09U30yhSNIaWDBxqSeBMZ8
nTMQZIpLUOXiT0gLyvMUHGRuo4CO2dfOW7ZNKvFsDQ63/+KlB7uUGdWBkRYwS2q2
j+KgguJVeK8STBEGtwbMiZJoyazc+uSSqVnaVvDunHPffi+BSyDuySVJBr36D8b7
L65JMxm5NZy+bqTq59N4MzWzLfKvMiGCUGKsZ8QMWHQEiu15D4jvIDHVJGrRHt8m
DuBUD8EGSwmInjC2yl7eIEsD1p8geZvLCXyZ/jU8ItBLZEDCs2E+qWIxsbg63PZ7
2lLcQ2zoeJPQ6+s1np/kVtg8lb4bfXzeYzuYNzm0uQoF6ONBG3MEuQ2TN55jiMHP
zNc0CnZvSs2UobefKAF1rd6JD4RWve8qnLhIA8aIdBGbm5eJr965AMVpBkTtKY4v
k7bWkpBnHhL7aBLm61q7e0eRrqm5MOSaWL6tGwHaUV8f2JmFRWxuwOwbiYSMVPmf
Js28AC3b8IUefmekYg5TqJmOll9/yZWa5xl5FVf/r8wUwfN7074qq+alt66Qky2T
m9xaqWjbG+hE+hiAEgvp/pr/qj5DTIUo9136fM+RTvvWd/Dzuph3DLuJRl0c3y4H
vdktRFxjPJWKUAe1Zmwi3oxtAqbBQXA5UKKEO9Hm/PA1wLbbi+SDYNZhRiorAEV/
BnV9ROhtUsy8qeHH4hUtQ3SFbXRQda7KYpOCJBMczOzgt2KiECfTxxUDerMx4RhN
FLRigxKZ1NIRbF1qQjXJS3qYfuEUNC1hbLXsLAOqCgaKhjanzYETlIM7uf0cFqFO
ENMAsW8fCIe9VN2lRdJZzBWWkbwOhMJwNGQtanJD01o/Bi4l7g57UoK88F0nbalU
1793eaZNjK2WlysIl+vlt2szkaXAVMCZviHmoISaFNTTyx1xwXWPvcKZCvrdoVBT
hh2lnRhUf2gYw6aOEEttkOu7ZuKocCUgXlO3mYiwVEHHYLAi+QATHQ6eBC2Xz1Ty
pZQ7HlxnewVkUQGKKBSw6KP6a8vCAHqqMagDHGUUph6XrJj2MOKQGRMIyFgRvaXw
i8wmrKzj4WtAVf1S8t7Fb3SkNxxRMZ4awXGf2ddWqvF+thfFk639xAhhoX1mkF+q
C9iWX3aMjEn9zAWNwgJQmpY4+tkO0scq5auNXr39MGo678GE1zPvKtL+xRFRa7f/
NYJoFkDP7RDmVp3pyHanDpzI3t85eLob0YYKLANSwUaPJd3k3GJldhKvOH8CmDHc
6XdPo2jAbFD2ZOsQ2X3BU7kiSoRLJzyeJrvYANrVt0kXj5tFxTs/HT6R7qu70kG+
zNJaVWOP+yeRPR6CtJY+i4OI3WGWftJz/Hxh5RyFRCsvKU+jgFS77v7K2gtGh7Rd
59ovYe4Y5dUotHtu6+9cSJATMOwxujHSc5Jh0KRX5yK92fZY5IqyC7koaHIeI5PP
nfe5bBPRcXktXCYXFDFONahZcdPYTWJy4rYp34jz8H3nNR5HzP4mr04G9JLCka5Y
tb79Er3SHrnTRcnC4wLmyn6YqJ0i9+DTjdvAEBThzlHWLlikKH55NP66L3/wENO1
YltIN4kM2gQ//AnAuCVuWoy3/QKDkM8f6qiHFgGFhrJ/vqdhbAYOnRWEu+zD90s7
pjgfmNWYrXNkUc9OqFNlMmRm0oqrBm5u9JgJc0UwYVdCrpNxspza8+fCpek7xgfc
NfRdS0dOhEkRNnHYDnuPrOPDY7s2J0QbGlB1WC9+f7uTlnO99GwXvRfLajEu7TZe
vlelHF/rYOKbc0FGOBtbJQTcpgpp8ipEWyzbhMH5w6uA6TN/OBORgUAeslfTmAcO
3tzu+X4kxFXyUMzbpoeCKrAoIKA3Nn4tpKHbXPbQAw8QlPzGIwSRwBN4c1DRhMV1
j7GAkfc9L34KWeH3JaZ//8iQg16pl7clVHWvaQl5AtBl6ZlEtpqne/vqDFTs9HPb
YaGWEarvQTESLE7zQDFusiWVYlQVdhfzOF7oFVTSvuDKucyl5SUMyGiwiCJ9+E3L
PA4K3Pmqo3Mi1rkzpeYp5FJ3hb1GVyoV57opKolE7U6rSm+RE2ZlsOcUwLpvyRPC
6f92ZzFGZB7Cg5NRDHbjQO23ajttCMkPrMzlJM2v21vLmFUEJZ9mjO+AmQ6c6wi0
8tXNonw+XYtCL38WCGRjZUJzClAByzML5ZUHAZsMGB0w95ZSmrNOKbsH+I7N0lcm
5cNCTBx/lAliV9B9UHuN1un/nWrjVkLuyvwJrGwIDTpwoE38W2Q/cEihIM294gbH
5resOp6JNXJrT4DFPTrr/K1A4w0YRuy/nEG5I/e/KZ3q1SgzKLU2DE+JvpGGbdRo
q5vuEBOKtyh6ywjjI1lZxRJ4yPrIwooAjiC9LISHO0Y/jw1maNJAEKrtxsfq2dlW
1b/yPZ6WoXLxo389yiz8IzUex2AWuxl3XA57j0jBFzuLrMwe5DYrMrxrD86OCJRr
FkQHS+wzMQJ5nYXGpZaYaKe7C5WiIAKalJ2nfo2YF0S7MeuMsVMg1WrAWxCQCTqt
Nh9c9k2FHMKg7C+an2Lj6pRJd7TLk6q9CWsbfl0cvyc0scSxDB1bUwYDbIpmW0mi
i5hA+UfT4jRn20VFXMWRQ/zU30zHbHOwYy8Koe8+pXPU0F99JTYmS00rcrq3m8G5
4fPMKamw1wO2rPccIgZxKqcHVlj1q66vTc5ClNt0BY8+23xF2N+D8f2727iTdwIe
JIfSwaJwvXzczBjKwzoIgnvxYndDLdXntgMWINXKqoTuxW+cMtF7UF3UtNw6DOTi
e071unkr67RxzdsCmDvQ/TADhAwkyV392VOwstcH+eR/6997HIKp7fZ+rQzQjJdv
Fz3k1I76qc20R1fSbItRnfwLGDyQYgLKmPU1oHQT6IXt/AdbwQuZv0835Tqv7qdO
S/gg3VXZ/A2/B2Tq+TNV2Kj7zBX/i+b4vtoSWfI6MOlliDd5L97izUc7qo3zMULK
ma7L1bvcfSIvv20p72iXuW66IQEf/NRyjhZJbl1TXOzgv5+Z7+r1glWx5k/NdSRv
cNz3BQ26Y0jJw32YwsBup7IvWx40Ra/1Z+j5gXOWqyFD/ad+sTydSMLkZud524eU
g8KObvy3uSI/eXSawV69DAXoY9KzK8LUa+g12kSzXGIAKpTeXh6q8+iQOda+xgJR
6PNGn2SI1GuO+yGu0nmWa8Z1YTrwikdmL1DoYNM8767E6FPMRQ6YXX3EvMIcrO8E
CJBI68sQvOSzLthwlwHUx8lWFG/3885AO5v8gmNHa+7Yje89D7TvLO9yU60wV4gZ
dGu6lnczYYfGi86UNYepjObDXck4ZF4gXpcpnO8W/h78TgUOIvcfs6Xz4FI3txdK
aKkW3PCjEQMy52TYlKR+8wtf5EuhAIhhwn4uT8dmmH3JCi8r/cS6shFzFvMed2HK
faR293aMEhBh11UzPRx+b3ud2SA+tFyoY74XJL1q08Uj9Ch+aDqyvKs0venj2hC7
/hWrMIj1vMT7RsjeMslyDeKJgAGO7AUrKuU67oY0PDN8lgCvok0Af25RE1zBSFb3
UtPx3iM/e6M5IfZyezmi7T2uHduE249ZwgLVtkJg1sl+HjXkkTIBuNIC9klVQO0u
kgvHZKyj8+HKA08wuSzGTbRpaMv6CHfD1Ghg8Cx0MtA4ERDD97y9RSCMHr7XnvNs
fPZXX15trf3cykwx++iCv2zomm8uk2SuanCZG2/gSnA10D73e3gPTXCQhK3oc0WH
BN6fTVAIFOEAD1eOd38D8ZG+nfaNqN2UeTKTNDzJ4YVZMa/D+dnMUZf9Z1pSW6B3
MUewT5lyv/lp3AzL+VM2sZHdPFnSsGnY6lJkyUAhGPoALQvbO5ljy/SWD6NwmBwp
UrmDL31NA6xohClPhXdIBGiG4tHUOJSasTF97YifAowsqaIvRIVoX8pC/vPwhe2J
AGVGQxRZBZVlro0CAEWadpj9i2yrYxLJpyRBn6kSUngeoX6jl5YwiyPlaaYa+1eL
16oiR/T93CCyL/qxyOl6MpYpWHQkJCDW2pKMPd9qvVBHQFnqAdvPnbVVLQ12CT/w
bmKGWoLKBx/wwHViTKxVpZZnsz16ISFgPDoQeDEhjs6W4kMf5exW/Qv2nF6QCEzY
+FhO/H1NxHLG9rE5XHFXmRISYtkKAQyPfZOOU9bvpy92F3vh5XXweGOKoZQj0rYs
d2+Vi3usMiRdGfOwO80mkiXvAGDMyghZikMaUnIvPrdp0FrlSubZRWbwlYxN6Fse
iLBHVeMjnxWvzdSsfN0rHFMvpQNoy8i55Ymp66GlxDsQ8AQRkmFbUGVmM5vQwczK
7m0HvJeuzo38m0+XsC+rB7ujfNCxrnQh6pp28kNAjU4fdb1P+vKsFa3Ts1ste9om
BKg+fB33sYoNXM0lin6BHMtfCx4aG3T4qcGQcxndFTj7y/nbNTX3klu37LzOVv0t
0BWJLFgGqo29ADY0VOSwYi+CFUG66SPqBzrYi5kwncvO5dHVEQ4AYFWSn95+oET2
kL1HgitIqAcAYkUhlOTWO6vZPNV2kbaPuPP2osp9BWxbMHg1exn0U7DR4zdVU3vC
kRR/o5AWjBa/WzmNkdgXUROd3tpIAteG8U8QGVHFuOllBjJLRqvvMSMdwd9ZSnqH
z7Sr6tnOOHvtyY3Vqk5E/KiEtOAIkVkmEPoJWKoGEgbXs8HCD2F0eB+rSCHL2MXT
E7CaVL/sL94Q5nhvY8g7LxSYN3fJd3jYFCW84UtLWOSrF9wfO6bDXS7pgz4mhxI1
bg0ocXJ1d2bXbZSKxe2xPeEpGsjcJ+SSUrIkxdmVpfhjH0v52K9bCo1KoHRsb1N5
+I5vofc7D5jiVx84LV0K7Dy5mIghxZGTVv6mm+YNf6iDE/AIvNlz3+admCVrm9s+
bcGJQx6eOCilzkKCc3XSI/F9SvJAbxsgZGw+YSTtX0/TjiEuexp2B3cJkKxatH+9
AjT5Bxmg6NFtklIqBDWz9kbpuWCQAbHqngDjrUd13wBPuFKtvxgFH4Pfl7+wzqbO
hQa4MErWyRPIw4K+x1GOU6kvI3E07xRpRbl9jW0hiLJRUq/kgfnGgJGxEgs5o003
B/72Dd1Zoc0t+eT/I3FrZLZDQDzrGH9r5B0of9I7zd6IflSXUPS7qKCWEvsfrJ1M
a9SiKSwc2rohOuVMhSwDYHZb6mItgh5snfMgpo4cXrjBSTjz9fHtbu2MtwMRn/9+
6QzqaCMpqRM009CFA91RCWin2JDuHazfmpcr6j4yIMly7BKHF5fjvlh8nAOCgmtn
+7kEleIWqLsRfHxVF5P0SU+Ur9NLw+vXb7UtGdInHs7v/6yJKFAIMUbymYtkihNt
up5ydqDwsQCLtphsiJA7IVfCRikwbcjLuJkMurajXPHbn7XAo0/4SnjvFIkuqvFA
N41SvZ2UZt9io+a+D+sTFO5s37Xl1nfDWkRqYE1Ht4R3lkpKTOJ3u1085ns8Ot1Y
DHlgUTaimBAYg86Rlw1ivWe+8hZPd0b87/6qUoe9imPPKw/U5/Uzkgn9Zg+3AT4r
kaCy3OfjHDgY++mvFC8X2cpLC/bBfMKM8YhHgQo1P9nQNGzVZJwtS8rFWCEg1LuN
S5NwggHW1EvajA3WW2PcXgG7Gkq2vIrZzEI9GseqZOQpX0ecaTMrcrqZ20TnuFkz
qRM6wQZ0enDC3dFG+K3mGgVvQcnx0Snp+D+TTr4pjL64Ts0oL9cQqQ1WtqmFfELV
BCFEY2Dau9Gf/CwOM9VcTwOBQVZ7ZBInbBqHETNCMP1d26laQwT2VItVzQ9Nyui5
gth/HHyIx3Ru8vnq30b1Vu7Cgve79FwNb/pzeZtHe69Nzs/EeCrq5e/kgRaO5oAF
xN/UJsU6V+Fsh7T5Mm4k8mroPkfP1nePgLGh9BSZHmDE7oBZw4yBtHqcjYvHcvfM
9mHUI2BO07C7Ks4AbLizfZ2mstCh+nkyzkgm9nbqqWWuOj2JjDEKUWIxwXJKkXYR
hNR/3Z4owOcdDYKJEhFOk7VKRkI5HeQ2x+EB2JJHteidHtG5XN6BszIS5x342PnI
CaXFwj0tgbbdavd03Mx9w/yKkLNhw1t7F8yi24tiaWrUUmwUgCdBfWApbDsMeFWo
DJSYRrXO0W94wj8jj5kwgXtIq8mbWiXwULpPGtb+Di1OAOF27REnWt+KDUJ+t7A5
QnAXfzLaS5L+6c/uATln67qAmHgboVn3pRYaxoxv/Nzm25m1/O8rOZRnn+QXVHMf
bl8/xagfMRcHZ6nsIWGk4rRh5a2h2XIHnW2ZkzDltbAswGpwh72opZ3FZqpAA5qg
FiplrJUGfFtg91Th4r6qOel1WnIJWXp+IZbgz1a5zc7W1evO1WeTIyCRoLNlvADI
OK7/FLmz5Z88YIRkNofnoS2BmBn9tA/WSLYlpbEDckFlI+ir4GHzOYlVA1RbCsfp
nlHaH8vVOSNpA6QAmvZ9C4gX7oOBeIK/3nIh2xyX2mqHyBycOYW8Eqco9fFJJe6y
WrWZodFgnQ4FaqzMjJj9tBLEiOdb6Y05nd68hXSpA1ENV4ccKIeduoFM1BvX6aHd
9HAFrY1g0VVrT7jWlDQ0O/dLBFgio0TMeyWwZ/X+HwpLSr7x3Ma+qdPBL99zqkep
vrtltQbNYev1oMJGJUMUjYC8zQ2HVZjNr1tvOrPDweqFCqN6k1Ed3MHwPPNRs6cF
+DJK6cQSgsl4+1+ikgLTxKViBSFRAIStdt9ReNhTU9ghwYlow0sigIJjoYz0eRB2
fE6GVbhio2ctM5S10J9ifWZcuKtNF5KBaEugCcnQkbLgXz3ayBAnsn6j5prPY3Qs
P99t2rmQ3bIDzhjtGXq8VdylWyEJBIj4yUAmgzWRj1sQxjeuiQzddnstLSyoZ0e7
+PCZ1uviIHY9rTLwpaK1TVK3w+XwaKKEMwc/pB4HZORoS5KfjO0rWPQM9y3rO6pj
nCOpFFf5Aa4S5bDBpGM1EzsrhgK2MH12Dd/38RVMUrRWxVznq3m23i4TyVAO8C+c
FMj+kuzc0x5xtm3cYMCk22dnTORz7TzOiNdOepD1LTLN0Lh2hiuF94fKEZvg0kOn
Sr2A/uYrjLtXLP1sY0uBO1ry7pp0+dVi1OwiIWe88cdCSE3g3TF4KUp6Q973zaW4
2CC0khGsafBWR9H2xH252gVqm644Xg0Wdd8MSVXCZk1ZqD1cVRlCisw7wbNg9ZgO
0gGds9BhbewcCLYshbhZHE2xOg+MSDiLVpJEPT18BurtBrBbJxNXKXTJW5xoW665
0gb5c0fpGrFL4AuM11PKKUOcf7RLrpFu9rHqzRWMb2JwtnCyakIaDZMrBhOsS8Ib
EzzpN3nLaES7WvMR+eId2COgi5P6UPUp3VVPthhZtIRC7ar4CegcQeOOIQfCV9it
x0Kijm5yPiI7aNhZXyaN7nYEBVM8/lsdIDGj7rHznqNsi2T7mVO2hUZ3fhJA9g2E
KR9MyNhnBVqdlV1CQhILWqa/OUA8+MyEKkBzuHaBjHChRXP3hCHN06iacggCvsfK
6M3jx+lRvehekU4J7slJH/jJ4KF2qpw8rPrVTajIsaY1ixNTpbFzMZj3A2DPUfwv
UKjlvcywHGAcgllSJQpYrmrYE5fP2o2rCPfcUXSvMhpQ0S8A98H6JqeoXHix6X80
Wbk7HT23Wg0d0iLf7YjEpQDux8xnKFNe2+ATgSqGK8ogiO8KY+3yLcnN/FaIHr3f
1evOcROvgquvDwupkwt3dBtv9IpfRcLwAx5+l75kMpeMnGDl42mBs2S1RvBjmxYt
uuarupRhqCalpoCtN5ITVzUoEiSXng2NXqnTCIFvw2cq9nQXbc19E9Ihpj/claUP
sYsWNDdbEO8TfXOc23h6FEjLLtImeP2NDqDxMsF9qbMj+bYTVmpEsG6NftrTqUUj
iGuFvcEs/vJCaRyaDq7vO5vQwA1hZ9iRpce2YfKPjwRelbhCF70eVxKa1xloQlW9
Knp3d5BFfk+FN3jjv7UsxvXtNWEkvUkAJxrcy/nBQjkG+boOUl3XPNukYn5vI5mL
LrPjdeBpw24//JQp2Iu8tYPcF9cdUNWVnPpR/oMm/wU2sSkJoqQLODVtNugQzG7t
Im4qlHTjzak8cKIcKWKbuhocKGxWxCbNcHhAwC3ye71AisWOyrmFUf7CcbH6JuFS
0Mpjs+y0TFKHa9F4B9t7xdBMxejHvD3IOKH9a+wN/uHISR21b1InQ0g3BnVVHXrm
JzQ6ADVzjymqYeDu3nI0Qu2vNlG8GrfOPj9ZI0r5B7NeypfGMi/FGY2jc/fPZusI
c5gV8BhixyIQy+FDMSAzFuoChwYJUw/rSLz+DX0haTgVPJPdIuAYSGYGM0dcTvkA
OrEUVg2I1exMNMNiWnCYS6LKrHz/xN5vnCMlUMsUD4fzOKdY9IBarua8K1Vte4+7
AIAhm6aclr3nvqpqHTA9GRFiuqPK40fWkckAQnmcOJIY5FWEQPAu/BNH/89HcKcM
foIpd+BmLbWpdHOtUVdLSPQLEk0TVEZvEYLff6oTcwFelm1G5WMmSpuQeAwYBiaG
LfpiKZZBM/Cm4EQibyQT7Vk3TP+06z0s5rPkPaQMOpan2wHOCDm+vdTV82/W8C2M
8ElcNcDjNs9Y6NHcJnn+6zK3ah+DXePyhU0gmDB/58eLCHB7cw72wmU/STNO5whq
4slj4ZBaQVfGAMe4IvK6Q0bjmaM7mIvnOfMJNEKh6nVHET0tL0OWoep2x7V1o/UD
KYnKohFrxmx0eIFv1vqCjnUMK4mfaqobrn75J+HWKwqEoCsW7H/wqZX3RyQVupUg
h1flQ6ztekkCa5T3kqztMIONHLrnj2DclUJUCnHRdexN/FuRjnXDWMGj0mxdqkLF
OZ4CeJu4Y0wmf2p4p5VUJcoiGI8m/v3KIU9UBsFzKIq8exdf+qS6PJCQvdWYRzHj
F3ZA0D6nGjMYhRkjlP8AvoDXPusjwFkgCC8a57yIbsN3MM6cykg8xedYo1ytDWVj
jDwbMTFdfmw8z0RxtkrhGOenfp8XDKul9tvbtP5FwR2/0VSxd/2hxkBbBEvmYl6d
9wHtA3vJWaC+zPuGfLNnXJtqrq/JkxS6slYEHdqOwVtWJ6sKtzj+FLYQxSTnZl6b
xQtXbAcAVwWKuCaLboSKJk6vODoZqRzg5kzvQKyT8GM96JZhlmStSR9Cfd5QezgH
S2DdPgX0/A6MFcgrHoOrMNQtzPzFO2IYWNvMJa4uUUXrQmWml+I+Cc+WRAER0nU0
d7rQ3c8BSy+zvsftur2Yy1ozEVl1bD4m9aBHjBzhtq3DMHpCgze3FW6Dzd1cHW2s
hZOQxG8LvPxkM9ow5kDrjJWQhisHh8ewDev4DuITSdamFJC+0Bp+J1gvpVmAWHW3
jEwdT6bFCHyhpiKaUqru9rX0QiNCUFP87BdAoHvEsth/j6H9ZQn/QtyBU6Ckv4UW
4dopFZIDBJd5PVmrdosYQ6b2uNYdqRkTi5uCRsc92KykdAqWJWwZSndYtVTAq8xI
fK/ULzzmX3cqQ948KUQakj5y8bncoQB+g52/510uBTUGSsxgBu15FGFzNlEdiplI
sb/ddLntQLGn9GQ9obdLhPq5rlOAz+ckE5h3gIBAMqZzYca5YRN/Pvi/LQpupkj5
/+2Bwe3qiLde+wlihcBd4lwFk4Zm2ecYKhZ5lBDdufASt7pJ44vq0g8AFriOsgXt
83qhfJ1fFRDK5cDHWG19UUAdhtsxhruS/9KV3sOWZ7FBaxHHvbO2oxkvursP9/nr
y+nDXsSDuTaAWuAMGSsVLxiMmPXxVcp+hMScFetQh+rwiSfHQlvJ+D0FT7YueMec
WYRyA2rXdYCAx+hkx16KECy+oJh9PrVrfmjqGIp22vYKUPwC2FqwVGbx4ZgRF30G
gRW8s247LUJjCHXF60KCeDLDgDxK+GoLzhhp5evRg/8hMd0CzrqhJQJoAfB6+lEK
HZEOLUZXbUscv/RfQ1NvkRexuWAgMz4AoLk6owAm1ePt7XcoXqH5wiz8YWXa6g/4
BT2M1LOpKkl1dKSbgtJxXYERIV/g4b7BotE2Y5srExclWul/rdFFNmUi9cT7BVDY
2UKA9NerfbmwSkkMX2uyBvbfTRppwTzm1tWjRdiqP7I7aDn2UyD4Gu1dTLulhe0d
FIyflfF7i9mwVzWB5ocW3eCArbHh2aIq7wzqXfTYaFaKQiPB5LcU1AN+q4VDpK/X
aXqACwuy30sOmBOeIjEK0kGhoJt5usBqdTM+f9yOR5vxxUAobJ91/Co+w3q0N0M5
YcQddI3fGBQ4hbIOpt8S+YpoS3Tved7PnRsr3WvkpzsjUHzOSR9mZG0dlM9CRtF5
ENaYhdRGdbHzNRZr1adeGlQBcZ0qMkGMWi8/08qbP2oiXUs9+91I+vkJKFj4d+TB
8vVrI/IJVO+RNaqjac79X4EtyLpPImFurfn4ZY/OVVeKbOKPiq05E1GNoHy/NJmT
FTsHBPK3rWsXb8UEmdbsvnNHJ+UOlFUmOdkl2VZ+TBr8MHIOEW/lBu7+CK+30beK
8r7SpFLCVFZlio3bR1qWsCnLiRb6DvZU8OjdJk3sZAksMWUOirHDEIBMNOAX7Wzf
MgcrZTCxri2+mQbJDV0u58EmpTlYKmaSwzKy/0xVuunWQNtxJw7TAGpBGHcbmJmx
KS6qhgIPKqFf+WyPaj2yMjhln72oIbRV1q4rbDPqjbtN0YaGcSZeusBK/B+OvkVH
96obyL0in2zFrBj0N4k8w4TMeqEdrrhTk1hok0o6cemzOVTqhfJ1+q6P0V7KHYJP
bY3H4dMjzRFoobjuA1CeMNSKyND5mqQ5EDDIhPHiSqa+7CApVcV4LjhCKSLdbfVL
7qZirEhljdQuA3XNujQtqPeuRwcBgovppYBAWQRS8O06uvbfdEN8cUHNj0v5PAb3
ut47cRfFbjGoibQOJKhymmFnhL01CLTUi8Y5IjgkvjYHk/y5UvlzGWLj31QXmMiu
sZb/EzR0Y6S/ZVZ1VMYEdGzeyZMhuncWZQgEKN8iDmZg1N35mnLKWG4U+Go95HuN
kc/8vO73znzYNCDAjKPNqKguc8NH7kvwB3UEnGmsTzKABnRBQ5sV2ebLbGI7O4qQ
t7Oih86ypXb46dfyIQVLG+/w1gxfgaGbXEQMhV+jbopLUQlbMd1Fac+sFNOp5AVx
1DYOpQG3JqDqvzKuSMOPwjfb1do65KsWgOhTAOm07fjRygjXuiQzvUYfoB9/n5+6
O4+kADXQ/o+rLB7BdXRirr5l14xIyNPdqhLRCxXbw/lxXdl+YVzsIJIkR4V8RF4u
1tA1CfdfXQ0wiq0WkmEQZt0g4SgairE3Fsj7qTcLUWSoe41PxrsvYdFLpReJwtWx
Ib2P1qVXR6fwmEXOpMHXIo6JbM1Lumv7rfeb6NloaqOPwAuCig/m512tDkXfJ5lj
wna4sHYbApBdq/NvIniv2/37TkzeLP3uGvAnMYWY0BPnMCqkU/YqkRkSi7o/nTlv
fg3BIQyMlLEX15fz4E/U2slrpHotmWs957f5Y3B4EPvhHygbM5DU8BYOZaaTp3qy
PSy1LyrDVdfGXTohNDM2p4WtFscj18oqgxkeF0x9Nrb5eVASmQCbrc4XHIhfUtAx
ZfdaDNmIN/ayR9N81qTfUNNxE/6gHUkNGb7b1Oau6OYPpNjZnKb0EZcdU5AxWlvs
XtSyPO+ERvA+7AhekReJwXrU2ByfUmjyVlCurNheNo4WVlX9jeUBPC2moja33q9K
IFwnIYZuEMLfKZjyxeqJJKhvgVQ6U8r8HxrrV/YFuvji+IbpgTIBsj7cPF26chAK
vqC/zgReoK6hI94D6fYxV2OrunySidBZaRlMCoezA1rPZji56cq2vyCAa//3Ic9s
7nEounW041asexGuqTudWAnYA47KG32z3QBC0WK3/pUVT5elaljc/JTa6JcfQazw
gITY1/cW37JjcO37vYHVtc6jxXdfTHFYDBzg7nTNmF5jvLRTuchZfh9oK0pu8ke0
Vbp+mo2t0kdiD3OQcMzEp8hqBqUdpXAsbXZK5642j3dYvsRRuUq44RyAs2k1OWor
7/vbHUtiPwkhCEKEohJVZ4AjgGrKbw+5/Ph8ATi4EBqEnTdGQwE9jdRy9z1BIedV
JHCL/XJB9nWD2mIykNNEYtznKAQvL4ZEFWVVTiWkmeJEOowDL8O97rSlKieTnWmo
NA5UZdBc3UDLIL6No7M95oFY16xUpzOjexNSR7hrt75tJNvtDczYkjWVlxhOe/sD
VMbz64Iaz/aEjtHkHHzfQMM9kqFZERke5VwNx51ziTAAElSEN4SjJNKOSN/Igotl
KLdSnWXsPzQXPbt6zo0J37FMsfEgKQVyV6h7LoIBgxLx2pEdIpreEDE6f0AfM8s5
RUQb7Yrj8sh75g1a8TrywtR89bOXF+HEa68QRC9/If0UgGmVYGmNGgJtEIEfwUGQ
2L2+YXAFc64uDaxRrbxXVekuV0nb2RDmIEBavyi8VCpNu9RYXrjftoDpyFnt2VAw
1seA1nyTD7hcVDaHy/1n6kj9OZOFO0//fU47cSERVMLbAI7SojFPtNfVw6i89JM5
ildSe4y2sCWFV+DE2UuhanMYEf9w1NmCgI/1uHwxe1kNNR0VVepwuqJPENB7R0pL
HZ6LV7k6Fyl8JH+8uaBwiQys1v6CrITihBNsEA73Tham3HjSXUPDcsC9Dfmsox5y
m9ul/H+zmWJq/lX+Db0r3cs6md3vzX1+uoa+XtKYQtdsqLWfDVX6kaq8QgWcOmWX
7thzDDAoFG6PvA4Ld/nuJts0PS7n7uomtiHZS97rErMSI2JJZ3bjaLGZLxQGWYMc
z2eTfbLN2E++JRpGFIUpISxYw8BqscIIK6Joz8kd7A38eGgorGVIqoy2JLQvvd/K
BnJY9b5MiXHfmWX60W0HSESkKLBNNNkbqMZXIbv0HzBVXU0y/XanG93cj9gCw5WP
KV2/UUU0XwFbrocpJwjX97NBcI7dvHAyXqJUJZ0vtvaSh/mDSwoatX2UoCpMwa1b
ETe2bTog4Da1A1DlZ9fw8yq9s5o7LxAwyvy4OvhrA5TIIyV4G6Yw2Y3JKjbQTWUP
F6s9BNGd2SSUTalB8M5nrFzvv9MJh41EzvIvOMzv/rUnfvi7VcW3Co386BdneEh2
wX5dU3h5KUakhBua0ZV7jg/idnc0p1ye/fObv/9nHg+DcEBjUT+iAjciCNGJyuBW
W3Q7LK6egQSHT4NGrgv1+RK0cduc4vZvBcS6DrzPmLmM7FUwAO8euPZkOcL9QtxJ
gI4q4S6xhf0pAD2Tt/dHK7b5oOmnf47gDzRlG/sqqkL1kSZzyFRrMHJdqZEptzXO
7zYPT6nUeCQR1ZgYnbVfIPcuUgALGi6l8Xc1uMNymbANkoFLK10nUmPcZuWrbUNo
VpFWmY9wf4JnUhVu338fK/7MJ2wKqtUWvKK1UQw+hCW/LMTls65eCR64lDTGnOlr
erKIybVL27GJasa1FQ7NaMUmSWlEsFTL54fQsB1uAFuVaeYKkDANK4ZrOfrFOzE+
Fr2Cr/BN1YFGHvT0TQ5nT8PXfCefhS/IoLlDdjy1nB74emYXCpE3wgjZg6hUckvn
GR/Lu6vTWeO9iU9O28gioGOcT/9U+aZ3CbdK85JUWSISp6+yZ+TGsdKbofz/6qRU
t3RwCvJ3ej7lxT43IKSRBMwEC8FUzpeqXYjSFZKGwtZtqzsRklpUK0muxc2LATEy
2+evXzLdEcFCwz3B9HKnwuoLTcveY6XTaqugMgcCO7jiZKbijBuGGx7lWSU7I59q
flkxIwfOi1LRKdqAozBxsyM9QI94AlbDMmR35/4hyr1RlGQhviQ7nhVfWLCqfkfy
hZ61y00ItnY7O5mo6lxUbxx1/lEeZ2WQsrJ8VSWQeZQiZC2tulNplSEGatms/9pS
fRJ9tjEQU0FykUCfIeMf1Sk0D3A5SAgTe4S3DsCWmX3suTJKZ2PH2BJs5FzbohQT
C1WnzWcJCUP9n7d2q7ofnb1HlhSp+TcJOZFXoPUD3WE1X3wgE9QXsZgK+tQ5clVW
L4GdtaNGsqLulWz3s236rEPsArIntTLwZxnudypIgdpetHrETy4wIHt0uMM9c4Bm
aoU0YeV/PWXgi6pQDZjCvZlLEbltfreoMUmsEyyvAHJ62/E1MzMDDx1AVSOKdPTO
Vi0DYVWKLIP6rl2kf3sloIHBsoYMzEdNxQf9rkGJer+YI9hS278tkdH/qA3b1Tld
ZpAxF3nOh7k0C+wIbrTKkVqAe5NjVYyKfDJf3GZxf1xbxBSaC8rVM1bxyBTeNWQT
1a34aVpaoOwOXZcGzwKNKxVqAgBUp8qBenX20nEPgK8WBttAVF2MdnsKixtLP/5j
HGvQj6BLjRxOUczLWy/wyeZ/l0TZL8KyftQIG+xEEygj9trfSwJC0ew47fY2HAh+
phxwHE42TMOn2JWjQ4GnZUfDcD/txo984nP7WtxafsRq/4Pd2eNDkw7kKqrGX8fK
l1P3kjFTDZWS3hVIHuKxWDuRAAzzOoKz9/8yJsEEHAy7Lbdmtcg9DaX+rg+S8hNw
zINPGFQl6UWkY5aNPj3CNJ4hCLasklBOfoh8Ol1z5LvAR3KxWO27kHUaiHcxL6xP
hWTapL5pg1hA4ONOu+xuaxQyDgGlej+0oaMsTvsHn6/51x9nTLusuHCe/XdAJaEd
71HhvtRSsyze3cK/RMWaza7+XiAKtqKCCekFfhSzgJ2TmaVWZP7GMDUoTqxiEWWS
aVK3LknwZqMZ/VV+PD7zqjkyY1YBkbP0nqaT3KOcH6fiSP84nh5AK5V62rSGPzyo
q/ttEefJSHTS5jGuXUhSc0tQg1Rkh9bN+vPRClneL9rm15YIcQg3lC+v19EK3A7I
7LweorlB/J9FcFA7NdxuiXaxZDp6F7kw9R58Ybp2FkLC4VfkQVKZdQ8HS0KONkvn
QgM93PGNf1n/4jpknfX7PPIxZgQS0WFnVIfFcqKTEZ/wOAMtu0qLJO2R5f4TmX5A
28BWIjwi2/wfIiwifcVV174XbnE0WTXvAkcAv/4QDh0uWrZry7q/XT8zLlUdGzI4
Oax8iCWvPTvRpoeL2agP+QsomISx84x9NCSO06jqU5vgETWx4X/JaAfc8x2XUppi
IzV7IWDVatzL3E4jcaRFzoSALZblOeLjKqLTD/2JN0m/mAYTYwtFd75Oxg7V9kvN
mB9Hn6ncnZYS0mEE5wxEe5vzCtFYeZsoaNPr7GQFhbQ8qlr7/CT/IR/rw6ItDlgJ
jn2mRuiTBYVf3dxPFO08tw1dYq0qUuOtuj4bv+ZlSv0UpIBXRBZNbZwW2XBC45kl
TsroFJjp3MTwfvF9hjzqj6X5DJOr8O3h3fCiHCBX9kz8EYEwrKkqpbM9Nj5Rov6P
8dBz+pXhuvXnm8Ygs9M/38iu75vDmeDR0MqAt/PKvZytXsXatBrzA5t4ntZjUAK5
z2x/O8ZImKEmaGY2EMU/X+YsxCzLjw0ow9qZ0f3qJjHzeg7S8eDPY0R25i0Afwdy
Egw0SpTGLsrasd0xCXwu5FvhDwDy4Ok7NRTILCLucZFlKS20Bst96f2NuCv0JmsZ
16+X9zJosKqHU0Ncu4ZJEgP0YItsVu48cdY8VAjHVNqMWvIX1K3IPVrt3oO9J0tQ
WXQ8qndRo80AkeIyMG7kxArJREUQKVMjlSj4hu37sWcXPmEf1coCb9c3TtydNWyq
ItKmmwOltOONUPAWOyJUKlEr/sxiG8uA2r1asb8/81hanS+TvYnblsZj+xQHtPvE
pH23ZKMTsJHevUCm3lq/t5xsqXZd671jUeL0JrrrPqV4dR09LW+qo4lL1h+awtYd
uG6znrs7NgaDj7yIMY1sTBx/GW8cgyWVBedkveue/ZaFB+rxtn2l8b/yP7AUzVln
IkB7agSUcrA9hbQdWJL0DoxKAW5QUbqNClBezG4EkhRjCKHU5ogIwiuTIz2IFqDF
s3rUyktJKWqGXHHN8lpozmA4pkIfYaHHZR7ONko8CGyyqhpAMPIMVYoyeAl12vzl
jfMmiCWYRQplVDxQ4R1DQ0PFWcteANMLDumrQ3PhsMrmgY2AcJ1PzA6tgev1QDlt
1ZW/auu+6yQej+UY7uG39iVOe44hHc4nIP2atWzT00TEyo0I5pRZtzpUTLayPsdH
IBRo1niCfXbZR36m8mljp2BdCoI/FzAk/gmWw5WaDRElehjcMRysHWgdqN+v1GfH
0Qu91ovtYkYwinu6FRtbpQkBxhaBBPAM3jWafIRt/nb4pL7wP2PDwMLwdmfiT/aO
3NO0BevTJ1BRsyoBg9L0+K9me3iBVNtVIWIbDJ4DssO/rdWHmcHdQQlsSRwvpBRk
fqkYfY11vwVxq1DFXyBrIAQuCBooGtaWcaP/iDl8X8Fx4YvjE+QnP7qsaEUMfO1Q
JGc3vS5PtIu1nU1CryrVA7Em5RV0k1Ad+upJK/VzmISr09tnemxMvbt18hADE1B2
cc0dflcgon3bQn1O/zZChFcpwH6p+pP+KI2MYGsjnTI/YMCYV1dMSUuqUdN6aZWK
Ksy6hP0M1Uwog352szuULMjPB4Hpjmv3TSpkTULDTZn/gMXHPqhvtGuil5h3lfyV
S4n37IGXKTrD6oX6N5R6LlAGNe/0vP2Z0cCm16RdOlNTTMFRi44DmZOrKqlJwUvs
AwQ3/sk1ATZ4M1PjtntyRrvDlfwS75GqOR5ah0/RnHeJw+KC+tfH65wuPbHWn0PK
pxgG0Fz+MreyuHko93D4+p/X0DYyIBphKbPwyd+m10EKLNUxWR+G2JJWw8USSWEM
DhTR1AooPPjn7i4/UMPT6FfmtzbxrQwctY3targg8VwMEFVU7qWESnoFj7jtBIb0
WXeevgPTU1qMgAOeFw6LgF+O0C5VvHQJYWVCGCvMxStaljwol1uwC6gn6hrGGdUj
Hu2dmvek3agaMIj1cW2ZNpj+9nj7hMdTJHtrm3pSf6tWTKmSZuUpJM7HJYJxANpA
XHFFuqvIPS34cmmlky4r63UOKAbZCiBVFYNS2BBbSi/TLceui/BMLU6RBGuRA0Bn
5sJt78Awh7KlC8YFRyE+LBT5z6Uemo2S769rnRGMZ2tBU8j3upMuR5PrxwUGArVB
Fo+W+xqRXQn4YX5u4myGufCeDtu+dxA34ryQSdQXEukSvWX+DZnXqrd+/uCfORey
hL8t6DiDT8s8I4F+8rU3H6uFZ2Bh6kSVDOdBmMlnbx/DJGIewZEnmnbAFyUVF5r1
DNVfRaBaHpk6VciyBZStULWRaEKv/GcA9UDUk2xJVpMoQfvcNEXtyxTP8eV1WitZ
WI6s+fPvXWCtDCYyYORiiyWNwAxtSq/+A0zUo1O1sFErWVL4x/jMr9sV6cq/Jf/9
YWATdlRecxzoWJuyn4qQMZktk1u/QAxJARCfwri+U79TSuWurpkbOi4i9OErxHRq
3JVAiAyMQt0j3291HsB7BsYvJILXVagWI/0hZtF3jM/Ok0aEMJgeB12iS/UC0OH3
vkGUot6X5ayynJuutG8yha20X8RQmZtmkabIQzjnIPoXo8eXcuQbKH6ULQeU/Yx+
rto//OnFjOILziteM9y1jvNXpaeFHVaW6tw3gQHNAKyjEEbrmOSLUtqXybZ2CfQ/
YmAa15sluSBZpPpJNINbtKaVC7NP8iPpbbzHbUokM8+rWmQGwnZ6bXC0EUpbLgkJ
5HcVBilfY1koTs3k0WRWmWa/MF+Vhuua9Tx6AELWfgFqEP1Vea82Is3bnRIDoIIJ
I7vwYl5cBKNpWzZepVQ9rQQwKQWjhX92bLfDbZmdVjClC8pN0cFUCCNUbbFUylDx
XvwohmGqjEBfTMS2L+UAtUHzEnAcZ2Dd7IZMTGC5Gjs7YkACYz8FeO8DO0MxeahI
yHZeNePvrdkGGzIlvkGeDS6H+DPGjb/ipCATuGVLzHlSS3ArupkLONUsnInE/VvF
hfr6nTtwnkEJvYIhUmvZoC6xiT537sigk6NyAF6ZogBD+3bzNcT0hTROlQiiDnfr
yHSAY7L7YlX4pttl/hhd86SWBIBJjj42sstBC66syHBEK7N/WiGY6o25sScr/CdT
sq/Yl5JscnT7FdkyxqzAlDbqcveVobl3z6FY7WOIKtziD0N8nO8ZgS/YiwSZA+aG
jn35Opi24aOf3ukLwAohlV/N7swu2tpWX//kV3zcnRLSLz6vO5HMN9Wl43O/CREK
Fuamhnzhiu/MYADwk23NZwtqpJy6eA/zNr31g3XvSxAb9Nb0wP/mh+gdpPPZux6d
lYzS4MVkdQ8ECknki50G1VVqjEdkrLWo/uy+KdwHIPG0UIVwELcEayuwkqHrtyO1
9eAibwi5XJezSUrnu7sOXoOL5EJJ1Srazznv24iCTaZpm0IxTL5WzN4q+EoBUTWL
jyyXK7SQ5V8wDA0g+IifEuhE9Y/Gomw6Rs1AyjJcoG5EPRSL6CWUFC/bGPzKOB+N
qOz9Iz3z7ZjV54MghFS1YCGXgNXQ//ewh92hBQBYC/A7MPeuFv+zqzx34uKtvaQW
wbEWfMnxjamd4iLtWjz1Ol+deSdoeaNg+NEUuaB/aeO9bBbXnqAW1gmw2Uxmkh5q
wd6YKvnWOOctOYmpa4nzc+X7llLf1iJqI2ZAWYvO9jGqsIbgV6ITwG391cBwg2NW
6C8fhWcxCZNpDzwslsknEXnBoxOLMIK2YaevYIWy3v7+LbfQ9EH86aouRLFBXZlB
kqvZBD7VhmJWP1ipmg2GbXH1NvixKf72yupfxarRg3hXoXWZliqjXYUjT7fOykBy
uBoBYtNnj12AVNrAt6a57qDzRee2Yv5jMcX8QIpjp1Q+0BQi5xEFzsTczQxwGiiG
jFrNCFBk9bqUI+zShBBhAtm9flyEZ96PHcfOGC1lZdHy4V7Kuy28HdWNxfAXh2/W
phcfIK9oKGlNPlQHsjsUKF34HiecuqyrTU4Z5QjQ2p+na2QDczsfbw9hvPiByoEv
wn3wbRYARk3SsTk4W5kb67MtT+9GUU3vgLGWbkEdp1YOF9ZkH0eXx5cfhoOlVoRg
eJ2fHf+B44NWYNZRSF3ON4yMiWQ2poSh1m50+dHoP45HeW82WAxlFT/RRy4702T8
qBSTtZnY74q3MjfZxMEjOLgkInVSTrbC63ncUDfh0DlG7R7KY9Wq7I93b3VSIhPF
C2GPc1oHmp7N7D2YI+GTJ02NWFw8g8+G03sH24UfDFXOJCC5iG2gFG2sY+QvJvU2
pJtduHRWs8k3BL2REKVE9WV1xSv+ANyyALaUOTO35qx9YqpkOSI7IzrMGPS//ppX
xw4DFVa31NDwMAGrZPTy0nkWt2jp2kMILPlVQQqt5kpfmoDki2PSs2cMGXEdTQLY
vuOoFSBYeAKPwfEjDvuJcpRCh5PUhV2EpC1IrnNMJDl5UCvP/WvVm5ds7ZiMbJXY
PT4fFSyYfrM+t3jGjaAqQEnIzl5v0qGFD/z0dC/iwbZ0QL9eMFT9bWx9U4o6HJiJ
9zhboH6eog0+F1P0sXTSHP/3ALZW05VCg252o35Ue2HkYOsGuApVybNie7jlNA1A
o8exRHIZEDYk3cK5JUAbOatjyowU5ZIOtTlUmtxdZGziwc2t8BFCekW52TJ1tPPL
EfyJLEhLaJ69s7C96uAJ8T07VLc+hp+nfYcFeTOP/2JXjRZnaihsis0C076RhXql
hMy3rHDzk2bitbqp4tbTaDiUsCYSj9xTKqhtfwZ0c7FilA82xt/lhUAlEEmJZ1JM
CQVvzPl1lFGWn36IaZvJzJ+j9yCpb5ZGU5uzh9rsyE0yIKDhkZ3MObMlJXn+AkM7
F0CuU2QGl3p0GZUsXELPF1yaW+szWLQi253l9JXP2LUNdnMuPm6O7SBdH8+6Lw33
QIeHybXRW2of0Pz/TQCm1FGWHA8D+ElnlKq16x+Tx0flGyTII3NEZb71E8JtESUj
tUV2serPgvtaW1sKy60FTii+Yxsdb4e11IObOHxtOfBX1+qlIuU42wGbULdzwfsz
alfNxUppSMx8cMp1QrzG6wiKKku1hQ0EOlqZOG2GNyqayeSyy9rSzByhZGjXOrQy
1t2dYcRIqCRczgmYUehg+/ED1vMcHucuomop8fehrk4uShN1LyhaS+naqzDqz0PA
v/cpJMIraicR0nDBvEK0EOkO5UybLW5FocXeFCh2so1jsfRwk/pGpPqOGTfJnECv
qhbrqcCrMNonI/oUlauq50DAu9Lfz7LBPxzeHT/UMFBaBW/YzRKQ7jmIyZXj1+ao
wJcLzH1/ILcMfil8rTvezVbjaPoxVLgfqQx5+8Sja62WODyiG5R8feCr9EJtrfcw
Q9aFU8DXTHPQikHw1qQgWDmCjT1oP84h8p06ev8MatIhU5RBqKNQLjGenJ2mqC83
VyLGLd5jgYHW4O7f8qwCQueT00hmQpp05FdtQLovIwGKgcTmRW0IUarI7iOKk5GS
UQ64DQ400w5n5QFDyGPQzjFqR5cG9nxE/W/rkMlb3PZhUC9iOYi7q6bMPBA4AKLb
Zt43TD6zbN2Kh7raNEWE/UrdYRp/Lzp9wKGBXOw2FhBDCzUPfKvVteE2IdYO8tmy
CcVPS6sYdO/jvSqC6TsJe48AKwwjMn+aoac9c5DzzI1RKFENEpgiFj4AJ5rX4ZES
N+Na/v7q+qcSDaqeJqgXmfE32fwNPy+YcWATV5j8bgi0jwZdrerz+UaLDPxuklWF
7wM6VrNQwFc6P9Kz1IjdI7rLIxZdPSGECxb+YpvD0ChmW7JvEJX0ftGGNBM2172x
c/EPS9cM8ikoQymRO2nU1jYqV76acQyeLgGJBojjrNRITQQLiy/nStD/tcS229MT
pJse/oJ2Ub74VXH0cidOHgnxjkZmRfS1owqbaBHWwBvOC3Xjbgv0WirjzHeaAtp8
2qPLDkFXuBDT6lh9hcw2cHdHlSXaVt6naqMA7suvL2o+Jc8syqnYcivyrr38qCIo
UnXFXCQD+b8/ZmpJVhtIQDhXQJ27UOBjTG7DOZi27w66u3ExP7AyQF+jtam2P3d4
q/FXzAzG7X1v/BFTFQKKfoJzvbpdz3i8WCrKHI2JPD4L1XEoUo8yHaArngN60tk0
IJCU84oNPACW3u/LQQj+pt2anznZI3/j4aMAVT+EY4WJBMvkgly89Z4sLX9YrvgF
9qAcVZzcr7JL1gTkvN/OtspNKuGlONCa6rNEzFevQjWZVZwNH3mVxX8FWSDB+Uz0
m17/fuLgxGEW7RrFcFUFb0tTiKi0wOcVkFacrXTZqOI/2L1VA2ZTcpNymMJyo+S4
+elsOA8dl9lNhqGcrZ4dwJUOMtOsKxP4tzmFkUezFqxbZvoE1vt15Opw4YI6Sg5J
n49isbSBWb5FY8jtOKpqL5HzEy1w0RYaO5Q89oCoG6pmg9bgiBTDjwCwB2Yt8o79
SRO2Z9Unx6coNPCuB/JbTUCCuxJexpTb/evRNW53ytsPSnOmHoXwqSI4/FmxLBJM
Y2TtCQ+Pn+0HXSUM46q55rPQ+PCzPXrMUcuVvDAJY9T71/hydLXzxcsDWhDQsq21
EWjW3n9Ps/rmvjASVYgS1hd7qLFTW3ettN8irbqKLFEBDdAP684hpZtrIqhX3XH8
bNveaZ0bvk6wSDkY7PKGorG0eY9pOuNxvGmoHA2VVeCGifkpRetaq71h2pFl9nM+
QSxfS36dQlM65UOehozEncKUE45Xg8cKlSL0vmeqvRf/OwVOG1AhOCSco/wnKI5a
PQ2wqBjGk8nZ4HhXFo2c2coGXNBhAmzCYCuYLNn/bdf2HqCQi4cf5kCjYThK33qb
dZ2Vex0+wwDRE7e6FNbJH5fLargoEVg3P0OteEwdaQirtltFU9oyZAxgju3tHPrO
BaQdqn/qTnkg6m/wp9oc6VGcChfqzZAlYDtqodaa+bjIjhk9x4P1Mh+sFV5ZsBeZ
1h57Ax1XdXuneHEq5/R2GiS+h46Gp7TVM77B4g+sCQMD5wQ8sIDVdguZhceyJjc5
fUQJwZad/zgFUFN8/SxrbvSPikHNHYLo8/g56rVaAKc5QOb8f4Dsm+vI2OuMdYiY
Ozxmwd1DRC9BuJSAes9xewKkIXa2ocnRxTXVJPdB0ZcOGt5428Y2l9Q2+eUSDf1P
/MPCAr1MVs7l/uBzZWAJFZqxYPWdWr7X4NJlV2KUSZllyrrnuapQVQysPZbslk1D
4bSSgaW9lL7Mf14rCi+E9EW660ou5eM6eN+g7HIy1YxOFbZvXcidyMy6YMa1dNBK
CgXWZPV0+YbgBHjdKSBfQV4qdB7JW3YE+fjsjgL6P6etZKgM1l9uoIFnJBl0/qA/
v6NHDkw3gurpe0A1w/ktRYvw6nkzoioscGHvKIyup29KTjWk3VVCjYkOD24Jkbt7
/Y3tq3yO9oV8nmOwOGKsnAA+vIQB/M2WEGOetmJfs2F5bsB6WtFt/DzXihD4TxHr
ZhjuYv9sAenPHJSs1MWLE8i9bK9LfG+yTHiX/3geJf99M0Si81bMdRT7EcupCuA2
LNznVayS9SdhwB65t7JhfOTtes0ClJ1joJVQxQ8VbkU8JyIlifWqG/+yigMRMzmg
5zds/VtoYzA3hYNB2RQNgK0DJwUurGfBf/CabL6xLbwq4RTMGN8Q4fBafnjt8+Dv
2J6313BJw5hfwbcOnbaeeVCUechc/B95jUOO9T4g0s5N8wFwTh/gbLR4SV/5+P63
bogdp/iUhXQ0cBiVBuEBduXILGIt1Fdq+59Ibogp9e48F6hguGSheFxyQU+tW4PW
iXUPXkyICSzLe3fgewJOL7WjxC3IP8DDTEoCfpkQISqMsctWqZnSJW/V2IlJDPiT
1OELdVjtBa05doPuJbp1T/2YUxg3R7wTbw86KM4l0gw2FFghroqhHKBKwT9oWqPM
HcBWgoxmEIFhR84DPRIvBMXCNYkrkfo/5owTDMGaBi/dUqY2QD8RrFGhxGJfLF16
AqaxMPvFOAztlc9K0+XwAnT6Q5GhXVfmFxDMVgJBJyE+ITt7OviOwzbFWkukHTiC
/t/5YxbiltiscQSB8v8nYCeFjM/aSUv+uatfmsMxLqsVyVxNAJKxYC6tGHR5l86r
FhXtiaACx+/TN/2GaiVCEHEx5UBfOQYB/MlGteQdU3X2LhM2YSPyFx8ftvvuPNNz
aUqhT0UDf3i2IHoUKiDjmkE4TmaVLu1EHHMSzX/xKCqAqy+5qLTNwfiOn7t7+E9y
cDUWUhX0Vl5x2uW0JLFUWMMdR5tdKRxjWpiykZ3ZZcqC5hc4JNkFjrp6PavYdI9Y
KaqXHAHPYxbzCL8FAdklUEW6dDxyqwkEt9e4GqEAohWno1U2T/iIFFRo6jgjX51x
tqUagpQxmzlE0ax4u5YBpTsnBK21Jo/ImTXdsitE4y0K20rmRti3pIvHdo5FY0Vu
ydsxGMqnucUBunJE0+Tmq4NfSHDdem07QImYJ22Kn83MRKFDmQwPirR59OxPhbGl
+SpGenQa72FgFs08COhRqJr6gTuA1u6zfklHumJcIT2e0TcVm7iNnsplxGTFrO4p
EwekjO6tLjG8KJX4/wlzFHAqC9MkvmPkGEWQEIKCQMaufo28bAaDSowtSvp1osk+
TzDAW14fGlesip+0wA7h2Cu86+tish84TtHGYgGS5eCeWnfYsplG9G3Zg7qELZ4b
mlkH4aDK1siXHu0ERZvD/nqwX//XKLlLzQ9G7qB4b7vrDIvkl9XzY7meJP61jh39
SGmC5F1TccRlI1clMPp+ZBNqdCaSq3wuFEPR++7e01cD1ENbGsbBdWtl5uu8611F
NP2+l+X5HLeWGgYt39MjwrPd1Rq3gQAk8ZtMCwBBhndrlTmVpl9wO0N2TwuWvJJ7
60Kw8vmKjZT+Z8VMhIIMLhWcLDhMJPykzJWhvjOD7Cwkrw//RxKFTmA/27vsLjfF
rLKdbqVbLaBChfHdPgshTbIASn5MJZSABN+RGcyn0IKuT402Ozl0lpfd3NloZdl3
WEjCiFZOqjYp2ehkgpZOpcH6fUYNfVwSbA1E0qEO5qfHLvhFhVR46hjt2sIE12Gr
GsyHWdqShtwyO+OXjsiQr9h1T0ltSmwr5cBSVDRq7JmSwcstxAmoK2UJhbntW7Fn
zLVsAOgPklvVmCj7BQhuqzVRv162aXyJdbrHdc7o7q99QcJJb2q7Hx9gEJB2rG2z
3gqGtxbctApe8Rx+YZNQrYHeIwck2w9a3/bXXQI0FmFYk+fLbc4PCceYXO5/bgKy
uqihA7ucpGyiloG3W63jig0FnQZGF5Um9PWEE2KdqzaoG+5TvAKDq/pyPsfXNFyI
h8+QPqPfgTpX47KbTIjcsHJeNpyiB5ko+oorkCDbbeHRZaNrlT3y695T450tVsQ+
ViIcdbW9M8ZNoM4u7xYAY+jS0s6ieAcJ3eI4Ut8iSC9aVq+/H5/foo3rXkCngqHe
g7ozOuMRoFsBQwcoOkzRdS6mzw8qaxHLs4wyWsFg7RzcABOXHmuS748HMfoJazcS
3LI1zRzfeWm91MYMM7LD5T/T/7QxQASXbzfGvCreBaBTfqj/ti4I8aWz8TT8t/E6
mdF8JfCUxtcj+s2mCednxJdGOu4peQ6TcoTbbiQbz21OntTXAdvl3ObSVm3D++Na
TiT1ooqDKKgD4YIvj9vzhBJPbyLZkjqlneLTKAW8s9SYdfgc/Zr0KuA8XJv7yAeM
sBqwh2FcK0o4b6qzdFm9t8W0Wtpb0eu1o08qlu4R4Wx5aGpmFySXBu6NgVZmZQ03
T03geSjtzOeO2LwhSutW3BEu2pbALAhekhPCCC2UPgvh+ki+hM+pn2QdA4JwdX7l
wnh04PRMrwuGXE5IGaC9jMzsNVxHDkjIikYJ7+hRsFvTZhMVy1hh1CH+dsF4JiYB
Ka0AFwcYVqwpfhfDFey/0OB6xjcxCYIK+doG94RdUOsl1jkmF3J7HE/nYSGGKhcR
xCBfE4s0ozVRYJXm4x6wzlQeheoHBpOwp4Ugks+XJ/2IE+u/Ajn+th/2zFor+8Ll
Ey+Chq/5XkFq0tW4A2mZLrKofVSs2+NniaiwxIU/2p09YN1EAbQnB7/E3Ad4uh1W
ol12s3mLl4mu4FLc5eJ5PUs74kVz8uZi1H1AvcYXtuZnPKuyrGFruwLJNyp2vBH5
frtc+T/q38S7AmvS1M2rI38mn5Zc9lXPCl289/rM1dVW5rZ6dTGnxoOLTYCw4T2k
wi0T0JO3c2iUYY0DpV7UJC8nxK4XUkGiDRso72iZ8wZPmJM48f8v2LpgpG+NP0uN
zeNJHlFmExIm1ux78oJ7jo7J3EMZLm+bqU1/emR/yD4sFwCIp2c1ofOV4skcVn5j
HNaU9gSPhmn6ZlRL1y9tcjpfBBDAMsm9KpDDzRj+Gd9mzlAxY9gobWAxCpRPZdJs
gaOn5EjDvEns433DS5RTvEy9eBKuVuxo2IIC79a5c0lLUULCPBDZf6Qt73jyzRWn
sEm6wVvYutvuf/jBmhDGcpYb+wS3kq6OBaIgfCe/g2CsZkWbWrpHGYnlW/C+e2pU
eQtDfTzrZtMtTXKBe6Br9/ftxydb/9AiUMGn3s2lQL+84uA/B513UlyQQ1US24/P
72eLfw0RjMg8zcwJx6gyCy1MF3y11xRjxv8QhcDcIfdJPBbyZ01ykOzLxm31TN0k
nWxEKiOMpIExIyRUbif5fSZe18UAsUobxBAvn7l509MB8xjbJ+qh740Y11eTudjx
42euIHhXpQNSi+LN/u6oUAmXnLOdvJNpknq1IfbCS0wtGbQzeDA0WTPagpZ64tlw
Tm0yDem1z/v2fB+b7G8mm28Nr0IOazhqiGGPoLts5z87bcU/H5IxfghHmVnpr/5A
sRiR8hgUMVIk0HzarFMufVe2SunKlNv+QfCBS2004k4ajK+gmgxI6m7cnpgb9wuS
iu6OJ//i1IB3+nh3fSnz5L7DdZCj1/mugCVDHRCu8nXMLAfZomCd1BnmHH6rXVZK
ugSXG0C7GNY3z2tDAtKfPPqVED/mwDY8WTvUBcZMym8vZL616tWjwRErJoEDGljZ
F6wd7iwiOrU5iYWmzoJ7ibpx37ErnE8vYgjQBDiice26PP+S8UF/fQbTgjlhFX3T
C/7Z02dCRmw/7Fqh7TcgE4GtIt9jBJADEPQCvrr1Zyf9Y4+pYU7sAbJTHngKwOtn
5wLrui8Nb42s1rLbyoF2yBhiI0KsxrQfXCML0qjIlhb5fyscfl0N4TePbcO0puY2
c287xTIwswhe53BXiPifzZKIR5HPpkeSSeMIqPuJM+LvxuNHpjZzrRteGe773eWH
RlSHO+WumCJ3nLFn3MHOB+VboLTMqgqDXsLfGRxojrzfbbRyYCpsWU+ODjgLSrm9
7V/pidrjbUVMJQN5TSSme53VTNLhCc0IVBQK2qjQdDrApU6R1gj88N+9Gv0JIgPy
pgLIYkeiy72Qs7Eh8O7BvdZBrrbupiY/9YZKLjmN9UyhVG1TW9zUnQSDuSFRBgz6
uclS+p7bvN0mBKbTCWtAGpEs6r7DpyoX7bhM7ceurqyxB7N8Qm/OFEcxRWHrpaVI
S4Z1XSg+7Q0n57U2vD84D+/03JLQMfPSvFRlXPRMWmM4NFBWik31EqAd9iuH3RLK
gNrR9yooovGM2DZvSTAmm0s8YhpFT07iEw1Ji2BOY/GmDL6Z/8vNtxfrzBsE00vH
/fZY+Md1pJlAw89T6jDcyiWVrtDWRO89j+vT/25uOwbtkJU6srHHWntzmBzGeXIz
pExTGkBVgwOv32GssgxxeAVyc8rKMm5Z8QF/lxviZd2PfrKI9Yw0kZH6oAdK3SuP
Hp2h8ROUsaf4fUmQ7C5fOHBVOzTriKjuA2RiBUbohwb+PX5Sl//Ttqv4RA3IoJxA
vdT98kJn6gGiBbD0xVpy5dkGOBZ31lZnL8/EWXJ66KLY92scje6teaiYiiHKxAIn
K+WvqxEo3K4MzjNBT8yYGPIWgFVz/Gwe9VvRPXw8rnLf7bq9byUB+N76p+3OluEi
dmy0BZNWBv5nVxLeGZDqubFcVPzGeh1jkLSSu6OJ4nwD8cXzKgM7k2nWjf9gLBhM
/R1zPlecFAE0cI0VsZ5y6lSYz0z+OjN6AkPPtqkor/ijGdL4GL/DPxEdDETROUHt
AvrJz0HoupjtCtTTrA48cx04VwjWhwQVpVLkA0AqjRD6KHFEuZC6flYHgGzts9Vd
LXmE/kYgPyh8uN0y+hzr3UoFZp3vyIZd0JKZz1ITuCFjUlrfD4aCcbFeY9KgsfmO
oSlR8bSyIA73FyINtoJGJu8PpeehkbPLICjYjcQtBlCHhfY5lSgZcmkI5vUjbMq5
I0RbMmpbE6BkaA0ModDcQe/A4yc5vjaTlNmHjOmXN1WDBHVnK7B5x3hlWp7Q1nKX
WVXWZ3+54/FpO8oQQslKHRs3QmIv2krVbNgtyYT2ws+jVYabCAeSORiqPik8Itdk
3V1+IMNHRmyUDFMLGU4tTCUIswe9tYj5bbIjJZJAlBzlO5tLPSvHSTLQHT0hKe+p
sRrYOivFHEkTY3sF9SNcZld04wgHl1fMdyBkFIv3zXhaBiT3XO1+wNdaGDXywS0v
fWf+Em4PY1OUHoEt8leaBco7T4P35mxCiS4LmVU3BCGHxly8Ji942vq33+O1/Kpp
xNApOx1eXe8770NITbAcyq6hvwAsd52ktFR5UrqTdrJPknoej4ijkNNOFgxss9sN
n6uc9JWIDd1igaVbdOh/DuaYl6HZpcwyMY8HqsLCtNx9nIHv2HceKezcOEySuDgt
Ss9d8tHsOLO4KeIQKE5FK+bigM5LkXc3qdU/cvN2hPmEui6gO27tY1WfqRnBDIIx
V3Y/TlyNhn4IDH3gyrCggoIdg36mX6D09A3KbQGjCS+8h2k2/MQA/3gLGbm9oB+J
dNNCyL9iyZTGO3le4tGdVKFn5kZJKp2QG4u5rCG1DQMVd3AvnLXpnb0PfCyf5SuL
2NhdcrmGTdfI4IXn3dW2DlMGLImKxFlsTspFr38XwXgdYGAVX0RD67Ng3FhybDWi
BSTwx0YM7BYtHsNYIfF9l9wlIaMVW3lMZBnSWV6WPAYPU6C6OdzuuDV/izm6wzZc
QH/OjoZX2GaUOhHxk59ovcFvfO851O/ytWpGPdgEi2F9Kg7Ev4agAV+Qa0HqNznM
s4vyG1po+QcyzSJLWyRiBgl+K6iT9SXU1k20/i/0RyTslVObhBXJ5XahotyaEmhg
PN4fz0Wu9Khhd30j7hkRn2vNUbo5c0KW2GAoRCl5MIbhxZCFqiMRbxB9GUOdH15f
cdQfcxtX1OT5wWNlnSuDVe/BIf2IIcVD4jGgW+LUng5iXIMv6JDSQOlpdNnFSm6N
A4tzHu1OiRg3p4t5CbumR/xkqVhSglRdgzamGExVy9LUhIp6PAatH65MXdxlUnSb
weV8XmvvqV5oi5vuD57WlDNu111wabQFEB38+6mladntrQfbWLpmstc6EEL41KEy
RwutvMf8OezCy6fG8ZHQbjrM0cfZR2H5gBjeqSfji8zbQiIPEFTG7Xq+rTCSs21E
DXxCAJrbdyneeLj3iN4nnN+cE3goKrB9pGDR4utfJ8GlrimggpTFRb3ThmTCKkBD
WJMGXrC0hAaf8ScR0NTCy96R3G+s2TIBrPGv0dG1gmcyh6S/2M8QXZdwAovKjhdl
frVjDBHcBTvdOO8Q/+sInmH1vXxrqraltlRgwk+Hdt4j36lafuh3ohxkhTo/TXVH
atnt1XaYYmpm0fLyswiZkaLX4ibLwQtCmwvBzD7s9wCktWu8qKX8UvJMQwanIqA2
rmokBmtCAWZT8SsznCxmE95Q4tpt7LsGaJ4K/3WZjU5lHJU57jWpeFt4pojPmv3R
2Z8tCfoM55Zge6Q+WeftxnTF+EyA55TgyaMYYU698zm2O6JJe7s+j6Gerss6ba5w
lH8u8XV7dupwoGMpdQ/Q3OTQn1OiZXYqN0IIDAfRouU0u4joOWwMPJZUOHd5Fqee
yIcv8RtuEfX63SLAHPhV6fkJC9p11LtCy65D83t8EPNBwueym30BBd79YwVVDbtK
KaL8qMz9uyxt+WGHKrWS4QDayTEgyCgZKKRyrKAUSwj0GdRCvLsw70TfCsSCIiOn
xTpLyPjiOLr5svYP07qeBg5oRXAktjsHMxSdUnECiSL1Sfnt7mu7G1xspgJ0Jj28
uwH6WjpB8oPn63FQyhXsIZeSNGYsehv0trpKSszfH5ryxF1yW9vY7tbYnOQvUNks
j97A+pbSCWqULwlGnfL/Ax/KjoXbAhvc6dnevLBY1hno2SMqMUSVBxXFIdhHoTSR
oJZN54zeNjcpWpAOtdQu7BqTmvDYW7JPcdhx9ZutCzgAlEObbM2FteRji3a6vMVe
Wewmm6DFU6rDmCR5oh9cRJZ3R6EYzY0YY+W01Gg7UcyXCzDhbaaEdcKKZx6/XVDi
yaNqOp/tkFU8qREoeli0ho+KP0SzXrIw5+uo1D28lFhgwwLRznzJ7b+6MUvtqUmM
07u92lHg3qr/7lJOjjx14bq7QWhzgIh8Q3SZl4oFc7aDCSrwhNYGgiJ4cPjLl53l
xc/HOBGQBW98rkZSLsfezcNdEMbou5yZmkcpCB90HRIm+SbYGUWWuMw4KO0yP0Vs
Iom51fDZ1aKmrzzBUM25Vhnc26yM6QBySBBa8lLGUbMuQVreEUVUpMcD9NuNYc/H
AtoenaV8Vo/2IOSeU50IhNjbCZkkI3oYTRaJerT3yU2kGULA6/4V/xmdfm5FLs/Y
dMLcWiJIzjLtUAEGhG3hVNxUfGwzJA0OLXfmFOVc9u3PFlzcaKq2ORfBGAsxSQvK
HHmbvQjpQRXFlX/nbYsOV/c3Q+E/cnArZn5jjn/lPTat8eZLMU/BPgRlLgVkG2Td
qWRTpkiVJkhU+c10ss57buqJgtf1i/SysdWMTG/aewkjlVROvUEC/7iWXgTOBv+4
6oQAT4eLPBMWkBpz5P6w1trvj9vg6k3RmWUAgm+94YsyxlEqxFoZRqrHZnvR1uWw
RRNi38//tXKaZ6oKfGNy2h8iAgrrVxwbwaGq1XQtxUqIeZvRo7XD04KeHaF+vjG3
sfCjmJW9eFFzpzo5od5LhFD+qzBlq6rNcKOgH/hPsL5OivqDuZiPafZBQ6s3k1Q+
UgG++btxfGmYQFzlMx8qd2DKL9h+mY3U7zMpIiLNZByV3gkwwQ+gYt7vifwmKPUq
0e/eSRZdtGdCrhLOk5VwbQfnhlsotAUt1+E4u8X4k3ITVbxdI0/pwUelOWlm4ZWH
JIY+1Kag0/wDkqbv3D43h0xoI7hrmtlzWE043h7ECuSlhUV+WDIFyDoNebQH1Guo
/VcqXhPThS01/2LNaPcbc+VeJz8khLnuJRAlL3QG09fzO7XMge2Mz2uUmkeDZkHL
6CmvQ7V97uAf/LkFVXQm1vch3Y8se9/Z9JwiuybNyBFZMWSumYYDJFyJZaV2IS0P
by/lXkdk6T4HFqQJ4TWDm5x9T/L26L6Y4iYcCYKM0UrFnKQvLkT61PFSHRNdkc+C
t57oR9DxeiztonWjbGnkPIGubczIu19nXhW8a3CjqljC8N6uXJeGupg+cxkLTm8i
Sb6KWc1sZndYk8X2elDVygByPGrbY2aGCyujva/MI9WwiiOdNHlvFcbxRaqdcsRt
kbfQL2nxMEvek0T1dLeWL4niEqOVqdvmn+wRXCO7I8vRt1NdSQK0HarU/U0nK3TY
HNnW9l/IWcjuWFpa5fPtBuMSGtPZykBW50GOOHzM5xpeeVjV4Sck0Ud258PAhmmM
yS9beJXgTnRuF7gWD4wfFyA4AqlSLgocq+ZlxbklNyqhdLSa2uf3gaeL5qsymUoU
LY+p329ndadGm1pGmtnxaGNcJkiJ0pNs9wWFUM5vqlxils4oRb0I3eC9H46Kaxtt
wx5AMA4rOv0MmRevk3Pxn8yQbrZLj0bw9Z4A/beJeWMtuSaX5mWNrHEid7Ks0nmu
IloKwxi8Y5hPggl2R+4S8/lziC9cPYJdQtfR2Uy65N++7U7jHSba/LTz5w/J52Sa
YPGtnFVkKnwcfhw+GId5fkcn2kfRAsE0je1KpDO0ksBOKO9IWb72TBJdOiJAaaLf
DIwsc4/dqeYYa8P30X/U1eGUY1PvBAGCv0iRJS4iy5HAHtyfBokye7ww832eKE1L
82uejqnU4xU8juT4SfcvenXzk/YfWMUgEit/1mipF0ep4Sd6E6bAJP3cLZnaHcvQ
sozsr9SFFGWbcqfX6JzGmdTspmHcfWZNgJuGkEYMcerXdLS8PRux1uMTSRhnoTM1
mE9ePU84Gevmlp45sKKxfJQllVLMqfV6/ZXBF7fWeJwCBsMH9+bSHByYiunavOd9
Debweq5fNhPE67tseDFCD8cGaLUaeQbZqtxskBTSeC1irf9HnlDrJPoTVvXGMXgw
Vd423bubob/GnlG+W7d4cKYuTne3Z5LZATd0SVkosh+4kvlq+ZXqRCC4AehcOArO
Wtdw2a1YbGe//Z2nBnX8ndsSeraY/FntbNMAi2IKDelXaVVA1Ja5FNirOiJ4t4pN
gjhXgeru9kVzksb/U44jTlsJ2IfTIb+cGCLqyOzKjz6ispOw+g1PYDtJ5yQ4IYbH
pmPbmnxnfnbRErVM/CHjAwzBexrdSFSePWn2hehhQtTDX4ffIlTcpFnUbInEdwP1
hNBc9p184azQft4rvHqEgXx+vZBwcD9yZRhHvpNrTXaRxq4m2Q+tym1TTJ7fbpO9
Y8RbRQkvjBmf/lXbBHDFHtoRzZjUcv8rRMBXedzc0eQOYzFAOBavQb24mWxovj+B
YdNELA8C3v38wqUa1qs6rZUQdJLoS4FNrEoY+CyAksBOYgrZwc1InsnHOgr2Zwk6
0Ntpj/qBEIcXjww1PCkj/dOCOr78ZzcRNi11flca+yEBxRNNqXZvkE/G24NjDTSb
ut2njHETIODCxYIRUQAF2xcT0vfp6j0aQIt65zAHkM2LRCKSluQ/CIlTIUxGpmwi
z8rPxuefBeMNjQseYi8UboXojvbQavwBKIxXq3YZTffDxzxpL0Er/TL48/DPDIJT
T2oRhR/TAd5QOBrb2DlGNyjTnWPWLtjeevg5hcyV3gxc/KEBtY02mlnS2v91ODn+
vrZ3YAgvR240ou+b5SpnTborCW31NC6xs7LxVf+uhhHBq5yxy/A1YtF31nIu9P8m
0NiDpL3OTFbeS01Q7S4aSTr4i1JlgoqfAMjZvf7Xvd8NBUzDGTEkU6nRgYc+QvJ4
0I6QeHKCVixHaaBIRRAMww0rwHKQCV7H3lgN/PhzIIKxfP9QODSyPCwNCIsXlbMq
Z4+46V5e7lpdeY589mpoZNt4UalC9ZQILBgwCewPCVr9jcdjbSqG1WFiSM5van6h
hbcgq52fyQHj16TG4Yii6Hbye13x6CK52ZWK/XCu/jwXngG4/5LjSOdBShdaBvWU
FYZKKWEK9WtNQeuKG3ptI0AAT4n2nEoQCnW9GsgE0nXG8G6yED26kmT+3JvFm0jj
zxpyIM2R7o1f7FWzZEe9r7FSQtM4AaV99ZkLt7kLn6n1KJMzz5eVOpZI2YJzMHV2
NO1/j8xObgFehzAtj1J1m2qQlNdy4uytnwsLXxlYsfL6vsmfdH/WTC2ARQLDOwBd
T/BrLrLVMYw3c9utzAri4dJK2V/8iSUcjv4oGOBVGAC6D9qea6jr3yqTYpRqUlFL
uEdzwn9cNbZzx5ihuZUdxQTP2bdTUEBOqO7TwRpD9ydCbozqgqZXGj3s2eRIliSX
HXtYOxHsNVYTy1Kq7QRKLQoTy2H2L+Gb0prBvJ7aYKK9FNESEhQGNoJNSoI9xAq2
ETH1fvWK0PFP83IREzzzBFFqiL1n0c/hqTQba5845KsXOP5j2AMBhltKo8yRb58g
T01KqFRQWjDzXzvOka8erfllckyAmiO/5bDLVpaD/scNHCbpv2WGcgyRr4R3UFni
rG9E7AW/0Q4qWODRzP4JGuDwUpH2zsy6wCgWj5eDhewVFx2rJMKCbTmQMG31WYCk
HtVnhOVn0Z52iXjrjY1EHVoBhbPgnuHUBF4R7WhHGWmKAezZMXarXhJHxOS+YV/1
HyKhONjkXYgSWJbKSf/1+pNK8T9qRN0HSsuGIZofWnY6wd1Y0SLaApn6MWsW9i0h
m7K/eFbVISxHDvYx1dZIA0eWgX6uXqjaT/a/B+8uiC0waQXjdN5bGEKaDf1RCDXt
JvyoAJWErQ7KQmheiXRcxghdABohSuDPu/QzJ7riXv55QdZpiH68z3MQBWMJ6pkH
fGFh08muRiGzusIYlws/ioHUo9fzWXKzW1a+THrdLUSE1IC+nw6XGxRWSQRZEwbp
t/sm1yIvufhzjSJRaSCkZqzLOyfd14PekSjV5wnI3ME57BaFhrZSpTwjzwrWPKUB
KMWK9+5TOHZyluCmVF3o7RmvAiPfBFI9NduM+WTgdALUvv3GPGO+oBVO+JuDnPGI
h0UKDk6l+yJQ30hp5Wcc6JMtGeHdYrMt/C3mjxtt1Po2zTp41s8Dd9FhPpdJq0nt
6K0r5gl0uHKfLpqpYMvxHZuq8mKy7pPNyuaBVmv5DGHkuHD8hGOeS6eoPpTAQV9E
SVIUJ/SkFaJxQxtb+jp68yuSAQ6eepXJcTkkJf448/yergC8ZAcMh6i3G7kkYN0z
Y/KXlcpEMa/HE3uYdA+bqlm8iY06e0l66PUXmC0bL3xHKgb+q9sDxmlP3nXlwBQh
UMPFQJQe/SDf0zRC8MYOn+WelVxLytdHd1oOsJ2ksTwo2/XF4/kjDjdHqv/kb63J
48xoqnctfeOaapuRUzXH0Uvtx5bTqLA/lAxcOAtNxoP2ULbeKTMx6D3XJjXxujFf
Hb3bXMAnahM+9iLzRa2fUhCtetRhON4K3gS1HoIZvZSjx0ZcAvKwFlDapx5+fmWp
NJd6yF4Hee6KOfOZLEnnm2CtGt6btJDWH4lFM8z7eHo3vCSrShqn+kv5CuzlvyD5
rLFp0bs37oIcqMp2fsQgXhpcKROAJpdbJ4JNUPZtfEKmkU+QwdIqcYUU70bA0Z0G
KvV1HE7NetW5Nl0iiw56IJzKb+SI3AfaJy9fk3Fmh6ueCK+dp3f9uouVts8YFSO5
EApEjCs5EnRDZiXAuFzZpIvj95QefCioR4IjsrVtzrPNeJ8YfkKDrbHaF7kVKXSg
WLu511yEFHyVNCeB64HmkTS/5jC64Naymi3PWXtrVG2Xz9Ysm5V5BUh/D4VtQ2sO
I1SN1t6cIM7S5OszhqzZNS8yHGdShDdhKegGq0vIQVcxDXK8/dg2rS/Lep+nB3Ab
91gNIpP36FexhylzZfKGtpVMjg44Idqq+CpZGn8nKmeWxsTtZKrz7hO1GFzVRD9f
tI78tAV0NGuTA1l1uHbdUFPEEHAI+ExutvGkb3zXpORdXIG/tFCBmOxnmE0/8iqn
E12c5kzC2xj2lvQH2qUFaumRZbl93CxZxoiXK3PY33LGSZrP7K+9ubifT8X2BDTP
p9aF83HQuEUudW1cEmW9uaHstYNQWW7o6ssRj5oPd428jOLtacgMs/lKbDCKxvK3
MpYbL15ZEe9Ra4cbZ++QdM90oZNHQDki7taC462Ejkoo/V1aNMFQSgvCMiIaHji/
/gwbFKkVma/h1z9H30O2Zakc8iAlZ/1xYirbR35W2IbOnBMt/d3jUIojnTnJY7Sx
v4odRMix03co3CV9Q9ibd5A0hq1jC7zD481AH32hQXtK87+1bU3SNdj87P5BrpSp
0SvNRYRkynzRdtb78iLl7B4MvtEY+i5YQIopN7UILBiOWmhJ18BmHTlXy64RgYkY
NzKRWN09MLLvUvg+8ZXNgxu1sKFJcPOHU1F+iDXaiPDonZQAal174E/hPKO7/DU/
j0vuGWV0Z08LFGsDz+Y1jqep7sSwvb7fEjs8LDla/pgo5GvtvSWrdom+aaIEU0JU
7IyvtLHFo3ZzhimRqtfwyIqxPXJqn2UhDzfpWecBLY9DjMbSiFmUzlRFJfHxg6Ge
1lOmJ7ULmmoJ4lgLFTfJtEJTYvQdHQLUaNq0Yp4zFkLXLGTCWdbM7r3/q5aULL8W
/0Wedo/tUAmT1i7eVYt4xgzbKn4+LKGtdcnCfsbuc1lMEMCrPC5XLmp2Hzs7k3vR
x2JFYnT19jSqamnrfYl89zW2cHpcMwysYPLVluJ5P9eopw0PdfcO9HuyklEvEgfK
8ly7hFkwRuwj0ptceEIs97NdFBWoomMYHMgBnf/E0AXUZIVGbyc9gQmEFgtrSdeE
C7Q48fnxoZnJIoSEkWYSVWq9VRBWlX01mXq5m+YMuz6k2pneXAkCPVN51LCjkp8M
u8H32vmnawivt7hgwEsSv8EkB0kWKf8o5pABM+8Iw5ZiTDBzGmJHZCLGWy+XMF0X
/NxIJWxLXx+vIHkB1RoQuyoC+qi5GUMPDfI0Cvz1o80z6ue91vaniC8FGWwCulWj
6ltKPpgjnCQ0Vc6jcU20P9nRHWd30Yjpz8NP/qL5NazJr6SgjrcWl7jMpeQF+GDW
kDcrtkRllQAcnok1jG1mnCHDfl4f9DYxS5d0Io0XtQy024o0V5lRmccgfaPmHx0i
ksnxkNXIvQhPVbnV8n7kLJS5k8Bv6HnjgvZ2YK6ssEtzCpzkq3XV+ZO1XWuWfHl5
cxhZzpSM9J7RcwCZV+tq9ExYUH/d6vsyGD7svYbOwNY6tWM8dK4cNvZyfutPDljA
T7DzM1yHz+sW38fs7Vrrc3fUne+/rbzQJDFnuTF+UCtyReUPwzpfnF43SPQWjiuX
38VOlt/LDAX82JQP1ZtE9nFJmroryGe2b1NnYoCzyLTL5ufOWFbU0ph6rVxnCrOO
+DVknYwhSBCTbo/Woyy7udEPA3CMh12DiR7Qx57LyTe0SQLReOUZrV/YzRjogxtU
wPWXkH4eqZ/ABbJuYSWrQ9EhVp5DATEjOwt3JVqJmj63vtBT42UZs8o3fGrASAmT
H4g/1+fk3b89gENPsLXb21+QaA+U4oUwnZKofsdKxNYjtJqAEHYZaKG1PxxpjvSQ
DuAm7OhlMrrqVEMfw5UrtBjupevKg3HcDjmBBTcU9tudcZpvh+s57AsjTzGlJtbR
aErogjgwA1WxwARs05PhE+lMc8E5TkXQZ8lWjetAeL+DDVNfJizum/7cKcXGYqEO
ypXPp5UB44Cd2fecMAMRtTi0TWO3ls3abuDd0Z2YWgU+xAfnFutN4T7dHSqWemQA
QXPjKiHx67hkBhSEQr4qfhOxJRt+BTEelU11432ZUjQm6qxefKrTiZbcZXfD5jPH
KgI13gsLVmysqzaWF5ScSn1BXkYWMgcPYotBHsn05pH74m19zMn7TD63RYBByahd
rpTLoTcg4O/6O2moTnpAI7Enr1PPAf6oYYJtqkHOuzm2LA62VWRiPmv6GBRRPYqw
7ABa9/B10BMBkRDU5qEERymCKbcbpMr6WHMdLUqD74YhyU4JgCoWwgmmkInkAAku
7nP/n61LpDlLLRlWiDcxhxItdOU9pEbEisONVTCSbf8wQqd6FzNnGBM79Vh4H4ps
zGE8x6lvqxbaaBK+tjeQednJ+H1epkX3myLULRXw8wyEMWaaDSe4vU1uBZA6dMFW
68gjYOhGFyRSJ+KIy/OlS3AjPS1XFyp808yGTOEoGVZ0IBkbBFNDXBjTHhVBo/Dq
gD5w1PhduxDMmC51rJV9EBSc8bn21zD5lC7hxxUh3lJYO2GyZh/VH8MHi/iAEu0J
wQlIiZhi8zJ0FxMrVPSQJdwjPNfyrml+H1xdzc5IFoozIpGiQaAxkbLiBU2cEWAw
lk76n+bt1PgJlvbdmLcpEXCHZJSY4m6qXsYjxibd7UGFGXNBxw7DM5ClgR48+riG
2zBfeZ9g5UdFK/ktEjh1230vHaPliz0SDKhgFaPmtQa/6kth3Y3zoj5iDS/JL1No
Z6IOFQgxTNpsAKPhwjIf90EPJmMgoXBcWpkbOe0Tw+IQFmlHV+nRBcQZwt6KCRTE
WfsTwMDHXPl8pSelyJboKyWgKxMEnw1Gp3JwKGMAW4bAbQEhmlc+W1ZavV302yzf
gn3xHp8QKR+jcUQQGMWvE6hY6zDwca7A1S0v27Rwk9Yz40i9QWHrRHu473MNFzp5
NehY4UInlbkWcCh3HolkA/teyoYFg6jP67Mh4+aDbIzxQJuBTcS/GTQ7d0wCWKdq
VkA2vbdmBUnPWWdYBCqWdDISm+J+OuVZsaQk/NXwlmt2EeZOa0vMB7OVoC4CAD5V
4EzjFntFg+34F1+cMnLV7I1hsn0PcRUR5bszF/ys1wwdO48gb7+/+xONOh3bX0l6
tX2SdUsSCvi0qmAdMJ9HLyMRmIEgEBkhspxywNhlSV2r11u6N5hqC4oRr3u7GGdd
X+mdDWz+hjU4jNdHX6tD3uubnfAq4VPr84Bu9DFUxTN/+0hNWVswWAc1a8153YPp
oZob1M0yY3rmqSERu3miuQ9VehHOp1zAsF3MUYhlhJc1hufAStQ4sdHsTcozf0np
oAp8g+Xv+OYepeznYGwtEPAQflppj5WlmMwCiN1ppu4Hg/ugDkrFSgSD+jLef202
XshYmODcgsFP4PRC3GIzOm9IlJuuhNPR3EwRq7kgeDsTWwymxRIHMJCAnUGSSfCL
irbF4aIxgXEvp8KZH079SLeAjWJoD1OUwZTbBfzudgI0wILKgp5v/nkjGc/BydEf
sN0G/dE1zSU/1YwplsHpKrLzEPZaCaGoPEFPKFTEbIvwYdN2QN1MUeLr9nQJRqRC
l8eJYXzN91tG/24W118tldgUY0/0BFgSTMPIJsLakynMWkcDMvB3P4Oi3NeNRyJ1
kBvodnvtwbaZGLhfIyAHE3DihTp4WzwsWdGT1QQ4/5zW/crDUrBXTD0yHvLtzjyk
z1uKJhgtK+tEpNz0vctVVDSNAiYXZDjGrcA+iU08GRYMr805ejLW91D793H9upE7
utNf+sBd01tg+eLHW/bmAJlvjR4bPY72z0GYPj/yg1phwSdFa26zYh2NL8JNdxNu
7XmMar01yJ4hphmUs1kgYyMLwCMocNkN+pBSGpK8YxvH8q0YvO2GieUXm9aehA3a
IFP25Vbfp7cvhVPVbZllF0qgIDccoZD3+inOt4iKkJlmnUu7suuoMVyUfYtnGB9C
rjhBcjDebL8C/wFaTSmwzgE52MD1YGhXGgfzR91xnk5J1hZYKpp/sxBL4vxS5ioz
a9VLCClxFc/DCTy5GJHbSmxwb4lRtN1P/JKlWqkrOkprttrxmK8TMV4IFZFbk1jV
Rs3zz7GYqfz7rt6RfiI2ICK0BCmQX/Dg6KKXouJB1ycVkAJA25bf7IylZUWbuBEq
hEjjvIyJ7T6JVZT8+K/V35rJZ0mDEKsfDpyP0OImbWBaHnRIpOL9nqkhTH5hNrKs
Zlz6wsUds9pe2tia00bBWydhLfamCDOQAPwugZzTicwgaR/h3AJCLKL9mTH5KQFL
88VhuY1y52ACKmIUV43VfvoNHTkvax7HSxQp4ccslDe3Xr87rOLWpnLCACoG4tI4
woVu9sLV4dIu3UoqBnBp4fTyoAa3M0pUxwrJjWC2NMaVHqNnMtKuFRBrLzEjDXPU
WDcKZYzvTQKZPm9eIr0IY94k/h3il82uLGX3wymgF/QHvJaAafuI+zoA94A1PHLI
HhilWNbCdP3oJJrMIqRIGX7EG2z+lN4IHc34S7ZeXzECT3iINYMoZ41mH5sOMz9o
eJKDVCClRbIPjtXhljoghLbBDr6mHwAqlZgDYxCSw0vsJwpjFCvFO2zbhImn1S4E
Nw3JWBzAnMAma9EfCvMHyBU3V5o8EX9JKeZFAfQnfyH8cdfWvVkPpIW556PVgcqL
AiRRgl3cnuZWrq72jlf4xesH9DuLfV4FKvsYlThTmmvxst4t4VrduRlppUBvdYjI
PkUQvK1NwzhjSUCrZJZA14Nub39ijRe+vyBEBbqiMOHd4wDKjcyp3pkkdaSUr9O1
Qd0Ex47xwxpYbyNb8AXOvqkiVoH6zv5dg7YHbvV7zMG857wHEuqiRGM+hvpV3lUb
181efJVnqgPGCZr2MUmuslslVJ8DnaIWw0I4qusdLg47Mn4W/yvloHV3A2l22GQt
RP5VdtWhNZYi2zbIcunzYlOrYvtavj8Hk5s/bjLFibDe7v9PKln+9LS4lYtXABeD
WHxLP9V02kUyWhBSQBHbHnqyn0DW2UlXBxNc8SGUFIRTxKtAbh2ex3epZ3B3zxEy
aOm0P2xulJne1YEkYZYxk/RCOxjCQFA9yxsfkDe1DVAjBaGtV3LZ+ivgv8kUEdyR
Rnxk0M/J/yEa7qT/ztVCYs+zzVkboXt0mIMtS9BvfzAtYLx6X7lScsCiiWNVdx4I
QqvDuKkSTKKMmQcfi03qfAYOPT5qbQs1jTDBw7W2/Rbsn1m7QFrArRPiitGhqaiS
sS1ErcMxqyfQ4Bj2m035AHk55OnEb8yuVVfGPXlHsUo4Ffm0k9UJZsyAi5J1RkfR
GMMmEuQQ0mq5WVLuxBf//ipZuQ4X3Y5TATjGZ+SKKQhulzhBgIMb5hPLEAMwxb9O
azCQYkW2Yoxi7LlTfe6DNBnwsIDFXXTzxI65JJxP5On3yc+CS8fWQmaZYTUQLJFC
Mf9TNykK/cwsjz3YpRlByDP/OdTpjVyKBv8/Afbe3V0qCvFQMR2FBOsrGBQLcPpy
3BEZanpoD+lZ7ugxVn0qlixlk1x2mCdoppVfpp9t8P6djP/xAcNjeo9smRC5TRpZ
nYx1BqIjm2tEk4HPb134C2fOdmbmvSwWFM1n8KgQJuBqy4SlucFS46i6ptVxQnT3
Geu8sufCqQhaAZoUwqMPKDf4RZ4Gt9sirDmaFWkBk4GAGb3hJAKDxl0jPuqlIOBe
pN2QfBSRZyzicB+r1BN8TdUOvGPAkJSU5hVNEMf0w4VAtDBL/Fr2r1JZjbA3ouQV
ICTYCLJwwZW0NYZO4NLr9fZ6+ZiooOIk8Q+3+YpBqcgzfanVv2MECC8yvhAacR2E
UAwaSJNME+H+aCd9oAMuelHWcVLntxy+kj2N8o+16wASUJca2bt00OUbk4g+Ef4U
CuUXwHQtoK8tSiHsYgAF/k6hcjz4MmgO3hvP+5ZYVTK7WmizSsoX/Do/E87prlAl
hca2cBtYS+rqATL4gmc4DY+8pIvwfjHbRncqeamwahCuO5hPVQQgtkpA4ZuCIfq9
PmRrFsSWA8am3/WKei+P7DPceWsI5cokqN2fkjLQWU7LSwJkxbkAH+Yomd+VIvjb
G5l91oRFjgONqce7SBxq/phjs+0VDzn7k33pNxabrN4LB90kFu5N9X2DNJVRKkcS
vCItu+PVVYPrW8UvxgjeuvPUga11BYpF+q3qZwE9Bgus8JWGwM+fZbjSEqWUKwei
WSYigP8oCHlzbh2CFoGsuyO0b3Voas2ld+YreehhF7KbdvqcQ9W8P3wht/X6S6+S
f7C7Qy+L7eR9U5Rpo1urjkdfNgkEaHUJ//sKe0jqFD8CElf9o4DbIQ3P5y3wkiW6
+mv01Iczg1xfQW52HUYIqp0CZna2uDrVPf+xsYSksICFA5761/kKtBDVrk2IVv1B
1NOYfpE0hhavjCbhXEUfVl5DJdPC6Pq13KtF9RtsJ+eJd1lOF+Zitp99pRQX48t+
sO/JnzyPOj+NXmpog/B4mJRMvstHSIttwza0O61cy9MBYemcQL2YOSQtQk0AbS7r
7F1PO2OS9WGibit3vUGPWq2qfa7mhWyjFpH83kEwctDvLL47l4HSltAVTOsoSoCQ
4RFg8Nb2SNnwccrcyK4V9FXYdgPbahEDMSWBVB4AOGYCSutd77XjW7+z1HUtpNNo
5yO31Kh5Rk41oZGSs74om1kcOH+KX31cGKQSJVJ0CrUsmkXhvKO+PzJEkS/6Ol3s
MHYd9hrZdwZqtuUP+hwX7k94npyJDC+z/Xq8wzki3COEpwnhygi5DtbbB2Z0cl9U
oPVtUxrAX0bPI2xwgkv7Rx6SXdhv6IMwwAiznjM+LgaOBG1qbyrAiEFeiwKexWEp
C8xQgKwD43O1SC9+udTjxepom0yEG89ZDMnCU41uMnDk20dZWWahYf45BMrTyrlg
n9ckHgWOsS1ImfG5QNQPf2moK+lnpgvXtUQmYZggF2XLx5fD5rj+tNpuIKPKPVER
3ABMDMyg87soJ8WpMuSefS63dqtUUQ/iq30vYqA7S1puVWjuN7pLwlTqiD7b6ycz
ivbQ8R4xrL3QueADVh5DPaXO4hmWjWM/OQvPQvrd0X+J5lizBtcoOVQ98tMidGPL
thYtb2hBgoc++Ao7C2KbPRR87pLSqrG8xdAh/Gc7IWUXFBnUZNn3vPBYb3MPQJns
MgVnMkPNgdwXgNXGz81sZ+PchPuAHVwOg0ArDp4fkb1kVk6a50YQspfKij9OtAGv
M5pNCXeVWdIKNDWUh6DiusyBOmnnYf1I8jBNjnqugYordfYFH0SwHFZXt+EEefoT
i05hG0QJ8a3eaGUChIm3jS+PVkJmS7+9s34ftzGhjiO3+8LKA8BAn4e3Dk4n/yTu
MOIY3VAspPSCQqr7tWnYwD3pi3Zm2cFasQE/ZaiXC9YJfYkA6wAHm9mpp2OjFApI
SaFsVrlW/mlyrSQzAUDCU6VFj5PjzJyYguhD9IP6rHtJgnrmEw/xPsWa1oNXxg4V
5BEn/VHB8iEclzXa6cpuHZAYQ0HWkmlDaAaUepfbsRQT59MDHDR+CTEzeIH1S7e/
ykMiCS3FEZg/yBcMeKxT7juxpBKjAksszUXsgPNPCRmxaJRSL/SJwOnEI0YdlyKL
f/SoZJqGyfd9/g8nt+0W6G3lSS6Zzwch/Zjix+X+O9fAF8EO7+1+vlLVQIISjeId
S6Kn4ohxChFlatvOtSdtOQiiGcSlUwoQwD+maUVFHpGjMPqr+3UEwfvFA9ZqGvGd
D+iA9HZQkuL9AIV/lBqvl3NZNP/MLytg2iqPFBHJYX7KvLk/PW+1ON1afmdXdOpO
kFTkdM/RdID7BNmwTTt1Z8OwZq7eYSf7GFcmwUk3Mgjx5ci3FR+FhGFpRPX8TX8K
TEfSa0cu4JLz5WxlqKxbcz+o9uxBocch+hCTLxw1WtMnWM8QRg45y63Y/RaeEUNz
1yU2NS9iKTVW3t7n5nZ9pzpAKseFD4l7xBsT4XfzYWhQR5udpV6ps75V+XD/StSG
3OsUQPFkJebRBvEk2K+IalmS7ORrfdXeCsCOL35fFPFrZYURztCqb/zcPWZC7LrA
7SEc2GJ/XTwOZJBavSvc31AYR8Tt8JXkQzKnJpT3bFzBEQV6R6wLEa6rb5m9Eh83
Ny4oPIDwOJ6oIM9S160sJZInBwsD5Y9ld+zoq/UyGe7+MCluWSvi6QPWKVJg+JWU
FV/UWXE7Av4GcVgRCEB+ObkRtSuJSQW+SxUz+eC0LhQsy5lZqo5ZTMZOAnzpUw7o
IfWHMVqF9LZUzAdZjGCCqOuI2wwnd6xo5+M1QQc9q+ccIePrvv8S45lJcOMWzgub
AeOWBR36USmxoIhM87FGijTWtmQbrZyBhI8FIutaGJUpq8hfdq4YvMAjtMB3iCGL
DDIoX6qTRFGw7n2Hlh2qqpy8ungqv3YsnqJ/bHdz7isVBvFJq/CM+72Pm+t5btkF
HxquETwjTsBuWXwZ0ACNz+FaUr4iHpgO9AN5ar60S2/HHbZp+FW/SovKHZiWeMQo
ZUuajl1613BINQ4cKeAoNeusT/Wz4O2b/LsK6J8wY/nJYTyE2LCKrd4uNqiX5TV3
406IhJXyqAPUAzt63yoEnH9V8FrFydncGftcNRREJmulkTgNqL+aNGIEcWA4w8el
k1kgaGgXjXSQ0XqcyHfOvpL/zPiMqeucI2m7UCfXlUncgHCBKDcJN/yd8v+pobeK
0L59//yG9aoM2u7CuOlV2MGCzJfJBk+1bVk7n/uO6mr4K+26Ew4MgwZGsuURx1IV
r7xnmtFLMOgng0xIkbLzrGxHoa+q4egnQiEg8mjvaf4O6NYPDwxwVFLe+9o78ADY
AUr0+UG6J5OEkYpP3bwOAihVnRypLfLAjAHmtVYzNDxc1u3IVaKQ8IrcnQLfZcnV
9k4QDNL/hS/GyTKVokdnEM0JsHTEyogGRdkY6H1ZyNoZSFT9NQoe2gtYU2YfQDCH
8VLQ8MbpWC6OF0egG92D12ktmMK6Omlh1+1C8vgCKsxGAj9teL0RfRIs9BDcGrTx
/KN/ON8pGHmQg7a2n/pPyLq4LYdTyCtd+OHw30dLsIzH3tP9tbZmvP4fthaI1Jd7
/9glIbEcxlWmjTm6mOqsD0epk0Acbp37YhTttw0so8QLMnxZNHUYAQUBmi8AxvF5
U9ZTZLHPQBCOL1Ew5C4OFs0FoEVrZdow3AgmSgFvwaya8HCkert1kbhLt2fty+J3
okun9/PbttTpVjNi3Pl8Ic5SV1GD4Y+FDroS9RCnBFSYljOtKkX3OVai3gysZ8os
/REcWtht2EowTrVvF1/ou5PsBIAkHfZY4NvBgp3I4DrAg/guctUrgqRdm2bIjHs6
I5N3LOmet5W5fvwN6UVnhz7D/SKjA9a6FW7A12TmaGxyaJzV8PaponyIEv9nZ28I
RagtB/AnXDrEJJj2sucLqA0yHdXhhOMAc+r+0qF0HdsiedKAtxSg9kj3BSziW7GI
pylvwh87NJE5LtCMhmI21BuNQkXAW4FNcP2Bv2/e8htmDMWTphv2QjZIVQKJezNS
A7bpSwB4c6z0Ie/L/xR7JXYqGVxQgfmDJgoRTWmO2XpMgOFkScj4aUDX/ETlRNMu
8FZppKVJ6Undsqyqzk/sSnVwZZXtcye9EUl6UJ4Pnr7miNF8R82FmmaL3hdItoaO
b5UB0jAGNG7QS7TDcv7HmWoPP+lCvouNAWpI0yKfTTZjOhhLPSgHtBPKLumbBeg/
v9Y/QuCivHg+U06ThMGQInTO0sNtDV1O5MZ7aveNbPn7ev73CDIxKMG4ygmAxPe1
I1U480sSJT0gN9QyyuIfVXBDpdDFp5Oa+c81MR3gZPrge8OtunCiCSAhk0V+4yeh
Qk0vNWkMdK9eL9pFeUqCur6c3g29dzCY6di42hDoTLNKwGuFrAjS9FvRUzCLrtoP
3cYKGergwSYhMZ7cvdhnu2tj6XJ9HLi2ePs7XzH87b35+Iyp/TAJ/eABLOotp4RP
8Tcl8vY+bkXC32GD3d87Xs7i5p7wypEa523DgHSggABSttmxD7M2g/i+iv1zk3TS
UAs/SJBz0sj/YytatkmfYKphaGN9BH8I5S1l9K+O3NzPDqWb6ZTmmR2j7bLHKGAR
kX0FfmEV70i1YhAC/19SAT6bTrD6Dwua1ZCvneunghozLXLkY4fyfZrNrzxzQHvi
S05DjFf1fJI7qdN5uqN9U/bBwH9Y7/eqxPciCVhkQUl06s+mwMBN1EC3EOeZJ23P
64PKRb3pemz5faKSOlL2N4ijQmb1rvCpUfNF5bAtzZoLaiKz6W+LGN/8D+m+HKPa
FUIJz3UWnV9Yg+RD3QsMmXwV8wSVvNK8EPyQkzQNKAJQ2JeaHUZ4bpVhswsvPD3e
bR8xRB8SY1AHkKRehmdTrEVfIx2TJ9zm9umZMATicJhQqJMJhVswZS7M8uczm16J
2f/BYGZF6yAlo7KkENeCFUSP83nFfklcpEcXDGTy1ZjKKvUhUvC/e7mhYpUFObI4
/uR1SGPzWYfzIVZmhwWdowFJFTu7Dxo4+0JP+xifoI7EGvLg1RWUCFpHg5u1JlBO
dhLltxJyrRTI2dqFpZ8MTVYgoNm4EOhrENlybMgz09sxiKDxGAhCNPZFSVRmSQ0d
BVOL1CxMe18tv4k7irb2zdcGqMcGqWrvpvnIIhn2klc49ndfM21lpNUKAxI4YROT
LF+cMbTHvJsrwNTszIZTGE6D7TygT1kh/VHn67GL9nN01l72kq1+V5lDHAqxKYiT
//QZ58fiY4C94rigmK9NGD/YbPXZp0luqxHjiAgRu2sWYUi7MTQnwOffid2nprMc
4OusA9bgnrOo9JZ/qSio+Zlt9ODCdShLQDfHf2h9MXyUTNK32Zgp2foXF9aO6rwP
du47X8VvzLFwpG8ViYr6fQkEs0j5aMS661J/jpq8J5i5SebJYaAZtcuKJzEqZcHr
ooSnWXYE5Xd/OE9Fbd5Lf529K0dkgiz/v+KacZ3O/fmQDLgbreT7KoUhDgLIR8HO
Sdhshu9YkJCZMYeu1pAE+WP/fTaVKVCGi7K77cy0VwwH3TY1F41hILPtI7OmCkrQ
pVeWJrDNLt5G4emlGno2d57V4C+8aag1zbIBoHn4nvIJ6z3z5/MwuscZ/Yxa5FaF
FE8ngYa3ril7ws/bqnvxwoXYE1EFhdZbTKIowFouu3IzNAmkyCMwK57D3sPeILmo
pIMpTozNVqvE1QjWH8iZfasYCDI3Q+szAXz/pDY62CQM65OopLSaq1QnGfSkq8Yw
Rhs7E2pmINmjxRmfrS26vf38UOukQkqM0G06yrqYxGVNyOHrKYNfXsuX07ExGtp1
WzcKbwDOF68Ff3XdZZ4HMie1KtYrVh+LkeC8oEoh51LzOAIkfAZK+3svo7X1r6IU
x2jp4H34UCv5PDE/qxw75fbUFXIZlYvnRbOc29yR64nQsbY+FSaDSIBzS9jEA8HW
Wq6KbavOM6dlHYj3CvGZHZJWpJPCT1CM/zjcHc/qVmq8S8hdtFdY+05pI5P+PMF2
synUFwr5R+aNFwNIJKm8noSIhQgXtOxb8zMhh0e5WR5KWmkd511hBfhKYjJIM0L8
RZ8ZRHwsgZTJZpnAsQUxVmpKJbkRlfPOMLrb3SGM5lHIPiCAmbcBH+pJYE2FQn/M
M0sXwSLuCMD66QnhAlm1x/tjBlcwrpQdtzCHXNL+jnjRtWXnAiU3QollsYx0G7Ea
1qqzf/HF1pGQz5f7bxYRBpfN0h5zbVOF8PH1cMGSXn8a7h01ONw5dlPmxtKW26P4
PP5K9ok0aqLGAdmQezY176YmAC0rwfjwA0WPXq+P5edzKY9/85+DiMpY//h1W0z5
EUD53UjdN5Ocd10hG13qMH2gscYcQ6nfXncwKRlINV3gIMzTsuuh8wus0FxKX0iF
3bRZe54UYEshTiarQ4tpYO/+K3gAdDXrdXuGOuOynW3SNjPRb28JOg1NzZVk6CN+
7Qad0kMLk09VpEBtoyfWWYoEU1A8FGuBEd1GAtfpkcgkpOfBDiV+K+lDIBxqKPgS
Go6g1Y6vvU5rjmRa+9C4OWcd/Kd9GcKbez2dRR/UxBw/7zL+cXevhAsDJrFcwzVP
tzXfG5yyY7z7uzjPztUIQ17xqmEyCsFKhFasOqILD9mK4jHe9xBM0tM5U48qMTFy
euWZA7skC3firwlGC1ShsOJicg5Tvoxddsrf7F93lsnn+6PP/ecoZK/hXoT/k86r
95jZAYrzo20UeS8kBRY2ug+SdTiWmBNiW0uDatn4TtHixbJx3YrntFWdmJZtt2qF
u/HtQ5XlQJm7nqj9k7uj8ZqKd7VLjEXTkGhDZvmyhHezl6NmJHexTaOoTNBXu246
nRKR0SrsegGZ+QiyJZniIBAMGWYQHf7DChCzNDdRlFa4z5ML+UtgpUmbzdjxghOD
CbYK2UbRFP6x7jd8Mt3su5pXgBDXiBY85dlu0qlHh+EEi1UiXG/4pHOGolkJSYyn
lbJz2++SnyMEzO2slc8zq+76BXVu2KAN/iuEHMGBy5z39k2uI3i+kYRfZX/G1jYe
+OZ+yyRzo2LWAfcTaZipbNQajNpyoqRDIfySBt9qog2zpM24JOb3k6xqM/Aj3a1+
hwwDszH+29floIt+TPBtlCFylIjLiM6fRnrbV0x7QQclOfzAUjymjbCqJhkF0IAY
/9A82wHP8ZbQmSR/V9VUCZFrvEvLDNiHfyAozVTOQDSctbnhYDn+FYpPpYyrcbt0
oc4WM4B4poxj9f8CAIUfNvf0cw6KDd0vt7Rkzwg8c/l61eX9+RGffIQHRp7MMu0b
QGe/AFjUa3TGlg8nEdoA7j3tY81Grhv3UMiXVasHMpfZP23kHjXz04nVD/coOOg5
uFItSQVsMear4Rqcsfr0BJTe31H2ccQLSadJFuwunzU8kMU6LP97ZWZKMkhD//Bp
dbQQCzXWUqhu8idIQXOzRVkrMBIWWjJgYS7CqNca+y4tbRO0onv7XtFkiPZjrM8F
vxdIidjlfZ0XlxCVgM3VMBGTN+7dC7oYBDpHM38Wi9i5ZOezT0QPHa0ptbxxXfbx
xn+tbg9/QeqA+OVTj8CxTzS4E0N5OoAjpsR66CCOH9HGK31C8u5OLDrwbj9Jmutf
NuvAFJgfLVk+LFlpFWBZPthTcMOJUUmEvxRjSqskEd8NT81U9baGaKaOHRr1ynh5
dK1nPYIkXJzF5y2h/P7E+0ruGPP492w+F6c8Z7+59A/bkBjIfUno7ByObmiQXKSv
vcw4OKZPuQPJYi5x/uDb28GjVaqeSLPaX7gNazonIPi9cdBTYVyTM09uNsIbmQu4
fPbYMLfmU7ZBihi5rdQtdLBQFiiQx//JKtTiDiM7ZEv6JEaHGYJXkYO5es07srVD
szNOjT66WT6ERsPV32YyPpL1XO7piExi8e6+Txj+y/OMa9qKBVwtcqeGYu622epx
SnI6DvolwXT0l/bPnzjxqon/eXo1FWHx71eQqqZEEaRWWBPT/BXC3K/r9iK3vbWM
wpn/oGW557PVq5Dwk/ziaU3kBa3Sy4dRcU3TZt1CO6lc1kABu9bnyE8viRH3/sWu
kPX6i3UUFLpry4SurhyH0uA43ZCYvEV0iZJSWiquiBK+dx+XZUXTgQLd14jyKlTw
dNDEPErdIuZmfhZCkCAN4JnCX5sgjtnsRxpJL4W5ewNAu7tu8NAy3QWOCR7BfwrW
hefp0g2t2J95ZMMvpw2ei8+33vdCjnbQEXcF2jRwF5sADaos9cTQmqp4A21j7SAU
aRK163FMsbaHIdNVYwC1ViHZyqkdAzH3CUfTqt6or4q0TMv35n7a/Pj+TXHUsJXt
GvH1goZuQOSIPzQdpRiG7jMHTNawoOoXoL53eYi3qpfXlRcoVK21BpgRkcy6fLY7
KauFe7+6RPhpUT414oUrdaGGKuzNORzEYAz7makOYpScP43Iapan7O/VQf+Klt9b
qNmNNH281I5KLWmvj+LTSHYztvog32SJNjYXIi060oeK7wvnRmRQFah+fnGsrDWs
cuyTdRIYdQtP+WSYBldzztxomo/Yr/vTZHGy8v7so6Q1ed/PgUYUVBgoPi0umdP2
E9pNI2BZ3eQg5+AXhsJ1RPZBwLzxk3Tqsv7Js/BxOG3yWH1PeYBzqzxftyfbCHS9
D4tGKp+IKvb2hvMa7OXLAkODussNIRTYUm4398n45UrzCQva13M0oLXLUkKsU87X
rTKdD3y5g4/IHWBwETzhzjWcSgGBSIS+dCPa0kz3tocKZ0/hzOv/oYSzMBb7pAS6
Epwr7WfcKiKz9JTpqXDddx1iAiExOCYSVXTAWDlcdqn4IZmfHYZ2uCnfs6IjRpr3
q4HP1Ec9jjEtbCHtTd+myBgYoQNzEvzbmDmJ1r8Bb84EdLfeE0sBrMo7OECJXYK8
yvqdAaN3omeI1pPAR3NuZNtjtdxEjvG5X83CnOvGEYW++4q0mFVNtyzI9trHm1ng
v5NqKQZVEAKiTxFDWnCa2/3vbVvGoyY8godwKpZHzL/zSGK7dzwkZ0TlLCIdbxv/
5Xncg9seSdZ4OdooTM/ToXfUMFaVY3Z9kDE8ozu5oaCTSrTy4HEc2Hp6nT5NgzBS
QyVJSSopQfJbSB0Z8s2qiqWTfcHF8noZH08F6dQY+8hgAMCpgP0U+S+KXSlGqDkU
/sfVqTcgCmqauHJ+7kZho67QBFkSkkkCmCBKLuQxA7PW2SYKzhXgLj5HAWOuRZk1
ys6iMbmXaJAEzaTTW3WrW9yboRvPMZX094nphBLknKWqp77Qm6tsYeAOl1QPYmp8
URXrvg27JUXGC+WWQEeEFEo6NUPSGbOyyALeqi+4JKTvP0g0+2AW/nT4B8jGa9lL
SxMo5nuVzkzu8teXtm/p1I5m1qgYHPtWF1a9VbZFIz0eRcKxpnf6Rx9o/ufzAlxg
jqae0RgK+VrLPjaNYehHc/N8YmKQDUBq3IfvHmJhFXCn6YS0vRLzyfuNFFj4xu5W
U7jYiaTKOqGg3MBshwQ3YYQXitQ54rUaPp/iP3TtxC3XctJie/D6gg9RUki7WHsJ
R+S7q31aIu+pKsWf29HVtkzMy9RwY3eQ4HubSh+5o7LgJwvIrd6QViJRoqpXEu6j
v4Kc7s9tyrcqZLwG3Bs8oaUllp0mKJikJshZX/eMSrqWNaG+79rs8ETEnpEPaK+b
If/S0Vl9GAVeuzYJevvhIsKugUJOLmbM/M1Xr9grolMmxdccvxDzDayV/0QvdkC4
4cbqTDkp+OsnfpLheWhkZjVIHkOiz8c6eYA9Y52U2VUr4NI9yZi4cqiTnqNMUahf
XUjn7wegTRZ76zAEEVEkcpxqW057JKx1wS2bI3HOcbEcG64IDOjDwo3FQHlQ1oxv
bikHU89DcORaiGzA/yAecWNS0pjRZ0YQ/dBQd4gPiDS/KVroGDNOOVVpQ7HX+Qws
ec3iriwZglFQW9wjee/d7TaZmP7WK1+hJFC6t9OP0vHoYs9MbXisRbUcGX9p7okH
SisWj1CqzFp4aPXR5uF2Q2A5WeM0/89CUs0+nzJgcZdWTGYkx6XqJWTowEk4klm5
s+GWxZy8rBF6IMBm/w58lHu/0j7d0zlYDCpshAh9bKncy8Oa2NbRgBH58rCM1U1G
IHeBrsZVKpuS3+9TfTXsdZ6ffdgEza+k9rOcjKoCSCkRoJOV2HrUdI2lhra8lgmC
RJLfv+DSYKJ0q+80JXVxhMRFNfGRQ9AgX17EoTWfbWLTdBxJkM3Vh+Z6g3fjS33F
up0I6Ifm1NU1/uQywgfN7vnTGtB0TkZpavvpb4sQfNODu6RoZkvtgjporUVuQipm
uk5IaR/y9yGhwSl4Q27yuTeBgT2SOO7H9w0EwXXNe1LcS/MtxKAJh9uMXB8lSIta
QjBSiogiZUC5ajM62JNxzFXiSUT+jfFezSRPKHQhZOjf1bUWtBAWYuZK7mDL+F9R
HdQRoSKsjZY68ZxHImRkQAu+2S9yScuXYHOW1f+skMOgca2Tza2Cv6lWvXAkhxqJ
VvkAuHB9u3fBc8Cr+ZskgMxb6HCyd3LgUjPRH65iApGpfR0N+wx5O7Uf2f4qRZAH
qyevkCAkalT94avqfb3dgUnrz7IiTrdrUr9iGsTW6F/gmCrz3baEHFnjGmvwElAm
j2IMkQAO7h/AEucZQD3YGZMj4qjg2D2vdvavfKbNB0IiPcaRKnQZqK9tqwpchs5G
cHnk5UYwFYxo2bTFTHPlT88fPkDSZsZT/fp+4Ps6h3QX/sQ960k2MF1KV0sVvS7R
dOIABocR8iSwa9BHpq4u+3qjcW76V796Y3sVXOQSzrfP0WcxPST6KCB03xSS6jTI
zvzyMOIeUf2FNy+NbK4rhyUD3Y225zRA96w6peDvRYetoMOQgwzyCtSrbT6ywkE6
pO/OPKeiSs+h+12e+QV1ao+8fRqiRSQW7pnDmM78ABKkypDSNgHNVApK3RTovCV9
xCLpULsnOdFGhhyLUWSK9Hjz+pmkrmDw5Spc+xImztkRiKs+b2EHcVEbxxEqhaML
Jymn8eH8s88fkaBjIyxIlOw4hkhGABwcG2nWMNz9BGsYpLTyfJ/ATR+PBQclYamb
+lvODdbzTQ5CUaoOqUXAr7jDiCwwCK80VeOgS2JVhmiLWWNSvBfy1Q+qNMc7a3Rg
qixbAKTzsNGOFTlT/3fUOsICz8XicoFvTs8z8ZgJjFMpKPy0Q4voA2ys5P9ReQgT
cmp9u/+TdnSuX5VaL4CFoZnhk6YNuWv1DbT0Gi9rklMwLIM6nnasROvNuwDKGzvv
0POx+q8yw0N+UDAkM+WtSt3CK2MLgUgfFkMmcHtNl7UvQXg5nLsBs81wNv/ba1z8
BI0R6ygfvoB4yjcly0zuRWkFuSuDYKMza0qVqC1dT97FTCYXOU7DDZ+K97NNR1V6
IYuOMF8sOVendMFTbNs+dZoMvqRkD/89calvUYBLYygh97DDmi54K7Ong2tcrazo
rVuQvCmwFGt7Os9N6VOkUNbZR/qyKXbx0DHPIJCdaYmbPX13+iqDZO04p0lY8cJ8
hwMuQlLdeIGQO2Q7TyLQ1QbxbiLsWNLPLV5x+NMoapukkaS2eSAYmfuEYDVrWErM
Zn8wx9ql4Qpj9yacSbr8mhS7IGPAqoS+oglhZxTEcszpdIJAZVrB+BCzEYKqnL7R
VVy9eV/1/q6pYQJWR/CO9/0fna0EHinaFoqogO8m39F/fKz8kEYePv5ccZbJ1buc
7JfqbL294QOCHOumC7Kt5GkT345srgmRS2TAsW+pB5f3KJiQezZedeR6GGuYrVii
miXC0ndvvEUnzXcFakbyOZCQufuAJZQxgUR8oCJHTc3x4DD44xMGOjQoowJo3ihg
0hZ9iZm40W0aA2QiJmi+kXRWG4241Y4CSKoe/zLxs0tU+Yv2GBlcQv8IvWiNtMMI
rm82YRFrZrVsUG85VWrEXr7WG4YRSDvVeYZK5YDEm97Rp3MAC5OWTVvNZ74CWSrV
gGo9urPz/slGrilNh8IZeXwmsCNtkJXj4Ks+S6c8EtpTnFfJBR8PZuK35ESSvPSu
arfZnTUOGneeONQsj7jtpkTRDfnMNLmlJyql3n6hgg3fUJL9Q6Xxa6HagmUnIjH/
xtQnYApmmhoDPckR3qg1++NfrQEYAp/n28CIhHvitqNom/Kjtf0/RSzD1zcOj49U
VRyWj5mzGhPa810JUHJTbnMWx9z/NpGVqPsi+0jVUKiP4+bPHk6ldSNWhZFqRT9A
daumFQCbZfIC2TG4IfCYf/wGvshUqMF/jVLFZH/0Fd4wT/X00g+Zr6V8P94ScnB2
zRR339RolGYX/Rbl+U4jtzW06oF/lzGXdu3nIVcgWDMGdR/rX53q9Mimkgq9m2V2
1aytjKXPaaQK3vgab7ALJulXhC1SfkqjkSZNApaK5aDJyQdc7IVYOmTINfbueSY0
HxD5gpG6mAhNwNDFfX36w0I5+rzKkekRxNVW8Hs+BCmw2rEH6MPEk7x1ClFetDJJ
vjFb4eOi17Gsj4khGe2AYo1kAyNKcY1fJyl5Ot0cxfkNm/yj/60zb696p97sKgON
QJJeTruVGLaMHOdAZGRYkf7GSFjdUjWGdfvUtSePUAs/oOF2stjyK9sJttKWUJ1z
f2c0tG54RUobdFvHg3Z12XLJrnndLlnwTItzOpt0Rpn0SAMR3YR96SV6Sv6AsHMM
jJafk3SAoyeHF8fo9zHWYqhw+INrknZYXWUFyAFvfy4L6WhtD9Zzy3pROV5NOhYG
FtmkRrZuxF/3F6dv92SWbykuFbjPRnJn8Fe4UKkyfb3AeFZRtFdCGUh28seYQmS0
YpSaRVg0tope+iaxyNbJt7pGheLiGhXP5IOQs6cVx/sJvHSUqrrggPK3yLd9cR1v
P8wBMNTT8/YzuAn0tT1ZN25SS9xcDZxh/UoSYNSrwaAQ6LMcORVuG1Lp7sMY9QSR
Cf7d24bqs9R0gech7MTTcrHCTs3uy6P2UUkNF7q+M2NLqzLnc3X6EoA4I+WVczS8
xJ54G11W9T2xdVtPN+DRYy1Qa2wZZOgWOuCftX6IPq6aqBSWTGV/DrePRr+eHgli
qGiDJXvIlHWfw5EztHnRrhuSLJH5Cr7ylddobkTNxUICpGMibt1LwL3UGybsiDCF
e2y9/Yd1a1u2kFZBmSl4/C1hr9ff+1A3c7Vpo6PGLZCDctjwgkYNP4gHcaX7i3iw
V5Fyp5mFGSSBbOOJss21RyYKqU2ogokP5YNqveeATVlCMOEzcMi8h1L6OsZ3DUe5
Flr+Pcr73PyK9qqoa0VID/fbcXA0hlLUC7r2a19Ckrl+hDoeYlaUqR6oI6b459nw
xT/uI7+D1ozhs50Qc7khDlGL/rfq02GjntI3SuEaHXYRnjrgHuFrWW6SWe6Fq11h
h4OXoDSAKYhZroki7od3uYPivpIY0PqVLetpbNpixYBawVuiFCUJ8LqGb13ycieL
PSP24vQpkhTEe/ofcRsqexQ4yFtUaQQ3vH1A3zuIxleyEg+blA5ik6dedloNHhJ4
2U8rdJoPbeK9s5lrVxs+wVRh/KhFEvg8hhGwm9rgm+J4H32oQQgbWkDePQwbO7EG
ISmaZGKc7zdt7CmTEEc1pK0txxthyepOLVVhB/i+vpkG2qgS+d60wTGdljKq1iDb
B5TmNerB200SKHWjODFtW+zN/0ej5I5BSV89jcBBD8sMyKjXR4H4CZ031bTMHJW7
hCRc+rXeOSQXlGHnbyQq/uRNRID/pL5XQ/s8S+6pGgwrYstYt/fWFOFSSos0CHI+
IzAYHv4Ce4Plbp/ywXVXyNrTP/HJTackReS+f1zgc3PCADbfiVa2uKrvDZ48nKHg
fPmGDpvM+Uqzi6q8SNI52hBAWsa32nuEhJmX/kJGZSmy4JCiamh4uBCylp8pe1tb
xOO3byn9m6cbmRnD153iJEy0MWso34KgqZIebTVqxN8x5cMZRa+NVlnWy/yM74e8
9kL62oy09EXzXIp57xVhHYz46JYXeIPLZmwLyXVn28HSPLxzOlV44taVtwbmcNi9
TPxz0waiJMsW1uHdQ5shQnT+84I5Uc0D20bu5+utNcFz81Z5njCMfq5iJziXg8xo
62aIQ+jfj0grdGqFV/1/o4FDIVIMipJJZ+CrtoAzU542B02jHXU62ua4Hp9S1hHC
LlGO6xA3WMRwvsKj2wgq8N5X80tVQwj6bm3qGF4/OOFWVS2Uki17QoKKz89XisB3
kxytjHEPETYUzZZoaRoMaqDDqLvL+oSlO+HLKCrJrG1gx+8JfVCOZz9wAE678Q5p
6JegFM+FjmolMWd9GeXY4pT70sydT0gpMfUA9Q8pAYgaZ3y0QWD+JpxJd2jC66p/
iURtnngvXwKtJ4Soic4JePwwt/tPtDlv4Qf53KEV2wYC5ahCvpBgFdYOkuU+Qab7
T2yXTrkE2n9EGgAgkYmhStbqP8njltRXPUR/cKyLwhQ2tZxo2iaBcZ7wW7xA5NcU
zdkuev/QMbFvoaymYyixi3DnyXbyjRg2neIFVNX/yBPzEOgqk1s4kWpbdfuv2Qrx
yxfLlrlHVvFzj74akNHwemY1J8Igb/zN0yxPBTsqTY+xgDydfzoO87dqfUq6jHiE
EuvXedFCy6NxIinbwSI3yxNhJyYKSOi24bmVOcxVEVOGrAoqrZy9CieTphtQR9F+
5Kn6A7UVg1lk/nZWRAIrZYj5y7tSFdZ4mpyqkLKuLEPVc98H5c5KLXkyt1rPs6eB
uRb51byeKdHq4Q0HPINRgyHn/ri7MZomlCSXUrinxkmFSAtpIS/AqUC06z0wykzA
y288iSX7pSaEDUV8qv6LJWGlNrokV92EVEKsHqSoKhcw+c1wKSxTO4sQddWhgfJ3
3Qyl9RSVJfSQP/keExDPaStgz63kN240wWJ2e4EmeEwXzSaw+3+pPL8kd1rOVgTD
placny+2bTRgZQzXdQQIj9qLEBg9JJitbIYhgnbyXA1jL5MCGfi3mzz3wY5zPOSf
o/oO9K5VucLr3Dhk6tkWX3KQIm9HtwLwurJnVNFj4e1exHEWHM0xUO3y3L7+fLUU
aLc+J6su6OWBB55pPFDBG7f+OOp2pPq/aRennnRqOSLTTWivhxS/HTZ1E3JaWT6+
ztLxFh+67zBwHUU2aL4UQf6ef85mljZt9EyFzDR/4NgOEmO8L28zStWlf5utQSyG
8dDcnK2jkpF/6w11KJbHvap3BvQbGtwsLANl2ii2XrR0t5FeTdSh2zsAulPEFTMR
HWQoWUwdrrbr+bLZJwABipD+Tn3odHVhMmPXFyYVcKxUZcmT6W5rYjBymtSra3tA
d8BdSXGE/suemHIVss5+ZANeOLP+scGZmKZ/TCReWXbFW2d8QN/qYiG6TN6Y3jle
KKwZkdnOlVPzqIDFbzsQ2HLjOJGs0ZZjpPPeywqtKoC7TFd1gx9e0Be5yLBjjuyH
+07nYL6VIiqEHtSRc0wc0YWrFFGrhGKu5BEce5KOtGtNcbUPK7DjmXUQ/T/b4xsq
i4pGhndGdZspIpBQgirVRyASFbUBfBUHJg5pTXGRgitFoPEzVn6dr8gx8IAR1hNC
OudgUsmrtGBFs4LegAwYCbzgfKV2If+P1OOSgvB38q0K+O2nXUJAgPL/gEF2dWDu
iN7GHAAZ2Hgmp6RqgCXc3+mUfkmXgOcilVpWcV90BpQw1paPfFxAyzv6ojhOeEuW
qEID7zW77Hxo9X3sRBnywgQHk8tdyMB+zlBfGjmaIwXyBVFCrOWRSDc+JZmU5dLm
9TSBzwDlZ2ziRyGphYoOxc7K245qlO8fBRd30NAlFI2WbuuCEREs/QG+oymJAUBe
QB0UqQbDwJghqJZnoz6YKhjBHkHiHGFhHNFGDpYd7cx6jq2kk8Dfl2XoQ128tttn
st+I+VRoHqKpb6wrGcyVgxDRbikC+rfSxG4FinElEZPFXvpeDJbkvsrDpEA5ZYUI
PqnMR3hIHda2/ds/WpHFoIbEztnZcui3caXA1BpKrR9z8/8f1+f5/2I6oBUfpF1e
4n2JGZOMJdlq5FFISS4ykmrsFus2H9RfPsaosxGm7Ve98b5dz9XntRMxJFYQaBcV
azRaD61kBKY1jQDKdx2aTjfmsBwIy8QTTqNoSql8omPs0jEuX7D4EyqrtEoTyAmm
nkojDB8g+k9KiMD9V2pY5iLG4Az/o3jyH9XNgsF8oj3+IyQ8yNEHIfxe7T4OOoP1
NX27Yn+9D2OviF58mV691eU9bKILrvE8yj28ea9Vxb8GHFGIu9KnJQvqkCMTIC+T
78Uq4ya6zzyH3xaZGbV7iqhUL4IvqGKJD3tSRD8MDk1lo8QVZEQkoQivqXarFgj/
GlSO4izxJ/vAwolX/730sKuJfWQw9NNXwn1tr9Xlu7I2yQX7/RPIAlkIpCGMex28
GzmM0BUVdMfbP9hLbgkmRhQxTzByCs1yKun1mTzja/Q801DbIF+WGUP8TQjUesQV
4tjsroXX1ONrVTfiiFRe7PJOyLGT3XwaWz0OKYO+P1VXYeqBeAaSM3TDWi2qvBCo
5SXSxFSbwhbH+5UnpFCCweG0Af7vLYtmCQ085BzzyrAkIa1WFVUTmVva4bQw49cn
6XRE6xYKNhXjQE8sFk0z+NXGRM8B/i7eA421Xyz9BaV6vbYLURDx3WG1brctdeY/
DtBiDYh2ndjimlFG4uLRzE1C/NA6mNTXMkqfD3fmG75qH3kqXJKW8VvJpnDbCYxH
B9C2EVA9TqK+vVoFTCY3tRDIT3FMQiZAv1GITIdBAODFzGQubxBgYAUjOEojDJcu
jGyD9DZGAe+JIUxvBxNvMPExr1FAMDp6LcDtad0uNLl7TUxZ274fC54fxH4Ejady
OmWpZYq4UrafGHGJJAPM8QVfuo9pNdDr5JmLY8uqfcwnJSmbv+HtJxYdHHdBZu9h
RbUe7oMMP8mJrwbhy1GR98SoQ9P54FRfErNLlyGtsb6UKmLLmM2Sjp3sr6i5h+09
3eF6mTfKfmpuVSupErIkS7DdvJ3wt4rgiUBiv91Q5zu2A4hOHC3E5OTwyrPQrq4/
sKyhUf4Fx51TPzm8V40eMeY/ZiZm5hldT+T+ynoJMULJ8Ucs7RFpU6mtZpbERQnJ
ofY13dSXq0Jhf0+75u98eS6H6xubdtDybg10rbm2+tXlhFiAy2/DMAP/4BrgbARo
I6BSguG5DpbPUevQ6sdlQu7kHrLChU3vF0A71NQsv53NUJKlRzmTz3z6v5VHxZQ9
ws+LN7oD7jCo3T4dFU0/sSXgpHBq20B9SLhZFTGKYZtc1Abp6Od6iuix1KRcrBmx
tdUL2JVMzXuiyDNnpvUxwOs6rUC/IP/le/G9ape/tcFSSMmBTpQFJHzTiP7c3Etj
tgLuSK3uwdnLiSi3Oget8QVhP2ij59O79CZ/w7cQG6iylBHSb5XLI2T92q00DFW3
CO7qaHOrPYQNE/WsvKS47tsX+PuzlAEGKzg0kgti/sx9EeyiFSoyMMWnDWzLrvAs
NLYCYstGhjbmg3eescPgPdYMW0YX2o8y5ulEShauUW6CbY8zxXB4Dc++0e4Bvy5x
5ed9chD6cDJT//1qxiW75PG72HZojJkoWzon7RhI51vhwfpshI57zxB7XpQRsWEN
m0rqqRMQjSSwvwCVmXhWQXAUE2ygm++C5tk9+WXUHtCLl+3k0+dxLdCMgW2P+LUK
xytkDuzL9hJaBPHef9C5qLZsnkyzzFCQkBrq2GDYT2Z4hMSVp0QZZVLW93cxBU2C
Js0pm47QdPakxC+TVmS9xHpaf8kn65zQehJqejnqx9ozsu8VT4LxYZlBscS4fqk9
ClbC0J17NetpeJZ6o74vuw0660B13pz/4D7H74c3Aw53DU6KrNYaWoeHR6liTX9D
6EeGHyItYjNRUp1abFvAdTHLm/AJsETLxBWG8qhP9xaxnT5aMLavrrSmWGSpQZ7o
iW7iQpOGnkMZ2hy5sfjgItk8KqMFHj6mf/dnJEfnG7hSk7j9todl0yWiE+b7I3Vz
fvVz1J7X3tk1e7fEdp8oEwo1AaP8nUR0G7W2LOGXJLub8hGG9VgN6Ughn9bPG6mp
ghMc4NgHBLZzzfk/RPUXodSVYsLC/oi+DbrkDltFWeu8pZ41jD2kwpxhR5UXYj8q
J+sJsoW3ZJEgWKAAMgvhWxlmpurMF5m2aKdbflPnJE2Zr88VEefjvbgoAQEmeY5a
PnVsrCXeWLJQRaaJGe6yCwT4ud4MZBtLMtowXfEwPFW2v0OsgrLfrgrGoOGJJ/rK
AC32NjMF9NRc7xJUpCArWUmbRwBVrVJvfybEMjApbEwcmUc/dQ6MlVPcMdbkUpKF
b47r6k82kVroGEZBrQruZ8Z1Zo/osfFRuAF4iO6t4qEl8j3mg+FdqNhkQCW8XHqD
5Q/diBNDPy4qcB5y3nDwgTN71HLH3jqlxuuxdDvFCTWXEngGs35nxznIWQMM8+24
LxOiyRTARsuTDE0fIT+efjj2+MacIMJvE0YMPUO66srQ62zhXQfKBOy4ftZc1P4e
XuJjRhRH/2SeE3zKgfyIhuB5/QTMRZyLiiu/0U+g8opy3dfEr/LO1HrzaAbxJfBC
vzjByLr1rtRuJD5eP8wrdtXN3ap3MZgWuzS8+rXPH8iR9rXWPL7mC2JYzacwnUeY
onNscvxNskKxUlgLC/lkSwKnBJjslTcir2PznoDvcgO+hutzYFbX6V0jKsOy0tt5
yD6l1AeA2876wHncY2DgDcxDH/oXu16V9NDo/L6/nqGMgW/xaSaNyze9ecUoiwop
4D9ofLjpdxY23Wod+fpGX6pDUm7nO76ZNKR4D36sgWTBcRvFkPW12O32sv+LUVV3
Dtuf3zd9/hDVsaQvSxnN4CVEU45IXEdaRmqzkE+iOVN5JEpkgF4hX36b5dbq2Tgu
alx8u3MQ0uSzqvlntR+YHNbUSVeEF4/uda+6di5H6LPkWnwUKVIZAUik8QKFew6A
19b8W2jeekWRA0WB8l0ohjGdHK0QWikWSvgt2nvSDZydnKlWz+veQZ/sAzOHgrf4
yLRei4aM027t5yohLTTkuHIrJOSDm39pa3TtZEOjGPK1PzjNPINR8ynzLYVCM+PW
QpqUXiXon6FIVw6JTlHXqYPBFe76GI1MfxXMzFSPkFwFBmnnJKHTk+DOqepiH92G
qMLp+TrNhXEjfw2nTeVzZFuD7HmB4WjW5vJIBwiIHfwUJw47dEkId6sBuM5HNtNA
8av6TV9YXUJv9lomAWWI10jg8rhUajdoVmzVyLSlPIPmVv+nDBtUZMPxyNs8ln8M
rUP919Ncrv3TWajSGzfoDMBf5+mrMPSFRLGNxBXClcpmd2TTnfjtTD9FGHf1RbX0
f0hsFje+hfKgH0fdGKSc6xAq8W4VnQiIXTS0WYk7wq0SepqRIu7GmODP5OctU+FS
ydFxM1uiC9q+5kM/84E9BaLlzVJTaR3yV6nAAy6pjwCx7vMc0rgm06ZWhoYL4Has
4jer17cgmykm14iB7ZLonFl+vOJ8TJL+ztZ4oUiuAYrg1OkKHRqG4eWIvF6VUX/4
YfhkDJu8atiUPL/RPGnK8OmzgcAstdyPH5V697QmojmDtEBXvrgwApoCnum+POWk
IDVxsQAqf6O93S/YazmYiTUGr6Z/gM0AssgIX/UWPT7voJnYbJbKoEwOPT33KnKl
iXWNuTg0Y01m7bJWg/ObfmEHSE4BP83JDoOIgOiqtWdDyECQdrXNWHfr0FmEexGu
Z7IWt4Z436fuOYf1FH3VkIGEz+OA0TiJyRB1vkldwJaC9TnMNQbl88SXQSEBcNdb
sqSOpudK7iSU7tdRTOPJ8UTSnpn+Dj1Vn9CdXo9AA+xW6lwN9/+M7mJlQFyEhwAo
CVoO60b+OXF7WyaqSMDJQGJU0lT/AljOuDQDXv9rRtbFireVCnWo3J6tiXIiGqVB
STE0ZUACQUbbaXLQOg5pwaVgL4ztESJjh7nfShIUW+W7/u1vzLC+Yi64XKLlUxQl
gOAfNi7Wv3SDwOmWDA9hyTeMPZwASIz38as6p12MYdbmfT1vnyAYHkcq+h08wp/i
AM4gHSOXU6wFs562L7QPxIohwnvVU0ENgF9nyHzFTk49dwqW81+L0iBUeH5UShgq
e6BdGfCNWZM1grQ6ebLrAooy5NFybbdGc3w/pcWBj2+Rls1lbtWNLrh5w022+S/Z
yzc4rMZxsHuTbljZKQ32rJq0iAItOr3n9zcitvzmb9qE3X3MR5Bav4mCRFJnH99a
dz94e7bIu1KumdrC9+/loj4FGiEsGGi1AiXaE+JII93AdkGHNTRPiWcaL9TVMX1b
djBY2WLffWrwmQqKC1WsKXdoVrFl83NsB1B2cIGSxcHC36Ra/NDZp8th7T81LPaM
W+MLJT7/x5klsH8Jl2R1XDVSJMZSgQrdP6r8XR42u3ep8BLDU01JiqxH/tTK4wCL
q7JGs5TUMOfEqE/5IfDC0fq3HRaBaHoFva3cU6TeiimmQJm2aMgYUKeael68Z8cs
3sDGAuyo0zHE9j05gUpllp2TbxNvmqi1tz6Lueua8iYxuU6YT3CaM3ebNdi5jZA0
oEE1dNsDFkDksgf7Od2DoIiqsJh85LpudUP0QoPw9OKPlKfGD/iA/9yzFlUTth9Y
dO6sDQD8Sjbe6XFLD8nYVcJji77PW6js2JDcVjfL/WGWE/txJpJLzja7sp5hr1pI
uMZbgy4RwtU/U7JRbvqNyoTYzt+h/MeVeZ8B9dUMPgD7P8OS7C7ICV/wL9Ax3b0y
4QZgQkj5Km5nTFjHJOQcMG3v5ZHVdDJa5nPRq7cQPCE1ndWZ/OE0fLlLEx1gI1cX
pJ+VqyvlElgWatVQUYQdBv1E6QeDoOtgbviBfP/XiTQOe9FykX5ig67pZVHjR42/
XyuzUkMEWA0MxZDLmCADotgz4kYyDXkUqheXNCkxu2mtyCe2/EtDOo/C2QS+evxh
Rvhf3jSel56hHs/CJ3Gi1FEWCvFLQu1T1FDy5gUiiCDOClDdkME8zuKVqdC9hXJX
q+2iPVZgL0MbWN53sc+6ftlHz07rnSvR4RLEQkqXGwDRsiJ6Bc532OwpGpQozphy
y87Te4whDJAucmCME+EbfoMxHFKuFA8VamWoZTXrfdSm5+2Pp4yuczwDE9uTvlts
vRbbeS+6BTxk56TJE20aXC6TnrcN6hTMPU2OttrQIGMFJ3jDR/BBCOkXF+cluN3c
N7QLBTUKvyJnx7OmZKdPqQ2lhWdFnHeWQS3SlXJ2H88Kx6XjOKmpPULWQnD4l7Ck
P9V3JvOzd68tPROJJeT2w05+OEe6QbmZ1d6bdIER8SlOGIexE2d7pXqBExgure3v
yS2U+haLR5Lob1/Oaa7JkuFdpd+2Sz8S3UVVKNdUl0mmB7uIKEEz8tc3pOxCZZOr
Jm33ytWi6Af14QxaPmeqwRHkdhmksk+8/EmGEUI3PCEQKA5punHDtux+LhGPe4PG
bs8LgCgbWnDYNFGMfdNsl0XZjza81NgVvwmA69VHawK/OEm3k3fPpV9CaQiUuuME
/JpLq9zm0fW+HlyOE7jKEUzyebYCg07I1ch/MwVLF0kwv6wh8MpjBhjmNnrclhag
34sRc51BnO+FAx20OgY6OC3DrxgWL06UdzSC4qqII73WiBI2jJ8+30AM4AvV9sY/
dpU1LceQgpi7XnTkOhZPq90lRQ+t9gwOFAjn6gxbGyLrYZ3JMtzRVxI/VQD+nJBK
ur7/DlL3WE85AqIa6R48p5SLVugPy4OHAQD2qQLTImibxvFUdc3aDGF+TPg+5RXV
zPXldSKBOB76XHFpAhuYKYzaN4r4YwGEIwf9XgcRQbgTdbX45sYrQ619SmNtFcdQ
EUgUhcC99xwUEyO+2aQORO95+eXaAVub2KE+XeW3pcgXfMFioUX3UZlm9U8Ek1bg
V9x7keAXXP1tcH6PJJPn6RvbcJ7y36v2Dqx6cqVcFYd/98WNDbbSqW6J7wWpW1bS
s3VYdlJ4QuA0nc+T018i3UVyEmnh389M1T70NrCy6b6Siwi0LPaUHPNLQ2vgmV5R
oaRFgDZqi6nudwxroBEQKO38AKAMa0EAYtPs6lNP+lCWg0wQrbK++NMFZw2mqbjT
styyq5TAssE9CBJy8LmUshxaTiklNRjUPJTN8wxQ/mm0oOBpkneHjpARzaT6cY3a
RK+GCahpgDQzhaADaA0VgoPEd2qJJJJUQFtMiYwrlj2MmiR7N/urUeXjABALpHxL
P+8VXd8tVdPGDrhOBPYbF59Cfgsl5vk7ferdIYDuvbLSavxWjHf1jj+j1elQCqkn
rWQ2Yf1gzUrrrfVZuwK9OBRoRcycQ12AlvXISDcdSUbFbpkHZ7SZSi7LgO222to2
d63SgzB79ssVxqIW9qrpwKxjnNF8WSD2dG70UDiMZN4OS+NSKbdTNrcbRHX+lw+A
fSn2hQi3/u7gGtRvs5V605GnsirwQ5+9vE90TfXSH+BWpEHZtzkvyE6F8F2x7MDJ
01w0G/tlpYxg46TF8gdQIhvaXbHbrBhuG0SEuUsfQNFgle75fKZDU4u1I0nIZYeJ
Th/pE4kFRkDNjq+WuTwr6yAQ5drobVUFBiGOvLRUJCt/x88WMJqlbq6VwHsn4Zvs
bN9+vOuNHRGj2lKpouu5TAWngeoCA49la/xV15W7jjmQoRN6aM1A2T4psiip7dr0
0KhwjPjVR/PRmRvmgHNbC8gm7jWHgYg6jW/3l2NDq/fMMeIOfWr9rh6hppjOqtEY
ufZm5kt6BJDKjcYIAB9fT1O4CXdiXXcaDbuSlQh/sqcNJl2+r+r884nPIA4qr4Vd
44bd5Q4FsJBYlswhtxopw7FUvY3rAShunvm7fkOE1Bk697w03s+R2gSoJUIJv3I1
cpOLJqK/4LbLrO1NZE1sLSwjBc5ThbiWJ0Esx2O/S9mb1y1GpqpNZifOe4gzk6hY
WkX7SJt6YdG8h3LrtBsC1N7gYM10gDmTqs6Ky1kl0pbgUzWAcGpLvqcIIS4SUa4U
/heMxo9RrgFwmxjW1m5WYsg5VqvYlrn5X/zOZmVo7C/rrwTv6k05j3FVVOYJ9WZP
JqA2FnBSGR9kgUpO2FH4mVnj0dQtF3hXuWJNuHA9Lo9X48pg0niX1/P7PdjnhByx
r0wlx7cpAHAzYn6lHF45E0D1wE6bCmxa0nophYdgY7vprn3/O+tfHpx9qp6HqtWD
TFpjKTRBql4LJNf0GQqZCgfPsxbVtAKhHVWcs14caKq/DuaohiyomRPKegj5qv2h
gozD+LjrusiYZ4mRJpO/8rOCFbILqJ6lfCZkmveXXxt4ArqIq0Cklgq7bDw5I95y
Kik5wO1ZAca1238A7K/OFVrtc8k88gpCTOzkw523FwEksPCilb3LQAsD2bhvmgMO
P6I9KWpbek56w2a1yRLF3tI1cb2qyGguJUBseEIBxSLoRJkgaAb/kvGYCPB6n2nd
y8FFKMMb6kSSSrA9fBgEt4C5z++IXwrGd0YXxjjabDKpgmW5Bhvm7Ge3G7ldpDco
IQ+d9XH3nqtqxCkfmvWJdGnDQ+0ZZvmKX7GWLZvFtqVOo1kasME8MYLaNzkLxuFd
iSsVqLOsfewnsRvShx4oGAy8UnI2HgeCGFl1w0Fm4ppVT4o3517kR8SqSnw5Ckdu
wKZA0y0G95b6Jd5fd/T2Dr5P2hHHr7ebRf9PIdk9SQHy6XJcfPFNsy+gNMgtvzP+
xfe+006yxyQR+z1cdAnctT2jJ1M+ICUmcUt9ivu/tFeBcutmRT1gnBDec6FAXC43
hRO940B+tVeS4Bc5p9G8tK3wwJ5g2jYkXc8Xil27SUNCVgJ+rkAqoJMxpZeVZL73
a3Pz02pZ9I8fWCDDiO+798cUAcdS9jKSGEs+wl6qw8u/8vw7pjYwzLgZjCpO0Usq
H9hsCB9NWp8cKsMJCa8iDDPjNkRPqTRziAqMnZ0UHWfQ4noSE1Ky4tQd6RFWtNd7
O7YauII7rDdwS2QDqoNdlfe0TJN2PmZjPONR5zmgtLk3qbfg6kNIy8LeTB/nUiiE
4LcpLDP7rzCHrG0MZT2hMPRpMnsxBDrtAdW1HzMn1YfLddHI3TabefvUGe+vAbfM
dD3br7TLEf0KjJAJdqtlb3aiZfhkCBShwFUDoggVtmfWFPiXGu2MY5UIWeYMY+1s
AD0CsPGqwnOnb7XeL2zdlGFl9x8sEN2BZ4j6MpIHoN6UBBDwzn28p2K0BSx3zgC/
rpSn+uESP36TRSOGQO0+8/RocqWJKXQVfeoYVeKKazM7hunOsJeBxe79C2yL6B3X
zx5YbAvtrw38/VzOcba3R1spnO+cQ8ne/KHNnV0SLlGe1GCdm9U4HAZWnRPVAR2n
WPCoQF9MA52a9wPUH4FPeYO9HK2Fu23cHjNS7Ewpjtoy65Z6VXQG3DoMVuDnK8fU
mBDiPlQtEgpl4urmnlNrfzukZZt42YaFlqU/fPWafz/z4W6fDLl1GYfwbLv2+gK0
fQP5elPuKjvmDZIza7SQOrBuVC34a6RYqC5oTjGpYrZCIsDiqo7O/FOAlrhrTZ2/
k60S8UlXTsEqAiJ3/nYgpAXwqRWvzES60YPzjCUmYZ0TIxYQQCk9OgwEwWxV4qNC
O2N3XMqJByadRPf7M+9Q/VEd0Dt4aRsA1wWeyc7HKq3KlAnRZ/NHvV9xpGSFIosG
8hy6FoIZ01bMzF1BGcJ84Mh6oALeWRCBvywwcAJU5nLDERSPZCOlm2EHFWlqPQYU
nT1hDuec334JKCNa738Z/pgRFijUmmW2F4OYFp74Aw7BczPo+JoJiDGxwCXettbz
4OLxPfXT1Eboti6AGxORd/RRMQaZneGHqwpkzJEQvWDGG1F6+zGeVDmwbLjSafgo
KUaWKIugREh0yOXAd1p7NpFkagw0Kdhe2EGVgcRhDvhKGnFKi38yjUBkI22PDUUO
XihAGgaUUiFXihNY1o27VqZcVHJLXG3P05uzrX+mmEI022u/rsPCcmBSrfUredGD
+qDQXT6Z3gDsjdgNSRdCSSvtofAhOV0MOuucdyiHvEtTP6jyZnoTOSgHH/OFuR2l
WaGUlIarWOcJxUMAtKzN38E49zQW5ORo1zEm35K+y281kdwPlFoweiWLYUqGclHo
z4IoMxjsFA6Fc6sM7DBA1Rc1E6ylC49IOewCE8S8wE+M89C+OXOUVTForT+C7kBh
3Yg1tZe4yQDFMFYaEk7no9sHzom36+fCFoHpNI9uNw53Rx6oTmECKjJDSvwfk/1D
dSvd5eHB8erUu0tISX06Ka5GLhZI0YasamUXO653y7i8UZ/KjqsXOxSnRkYiFwxh
W4f3T5SxAg8AZtmRbXwwHeTWpB1Rm4dvGgimny5mMdWMj+hqV9CZ03s9Ky7K1DLg
XLI4VfbFCDZMxHUEYc6H9VugCqqoXUkJ3J/jORyjkLydZ9bjSrxb3fHISqYTXM95
AJlDNNkiZA1hHQIrwY7ggfiFK7VheAHDh4PkyvyYmt+JUtD9bi/BdmlEXcPHv4S7
Uek2I2bdBiEEiMG52eRh8AGBTMRGAcj+XH9dcjfSgXdxaRM0Dz/lN/l9RqmMs+/G
zBi7/Ab5fhvKNPiJ3dGvNf/U3jL0WlYFfLw7/ApTTwq/wOS+d9a5+NJLWPjbnEg/
lHFBabRNjHSo3QHpQ70bEX3vwKrVbu3zgJ+UaKRtNpC5oPIdShQU+d9APfhIx7Rm
OVXICVYPcfiD3jzVO24zqPRYotgrhiCK8MKpMLfwzh/R2O5j21QRs+9ryylHrCfU
Io1hROpUOxxaJPET7h3tGA5YU6+Mz97zhVUOqIZ1M6pLPeP2nNU2ZLDSi2E/XKCc
EOxqGFQMH1HUknwGewNqxi0f2+Wa8DT8Bg9W2dAz8B+YFDXkf9uDpNX0Bv4JZpFg
19ooXORC29cYrvrd5ivdjAkycOnRjnQLk7tZc9A/QSpxdZnxdx8qndt7YKwfu3ed
Ob6mphGeJEdDt8Xnq1JAfrqt4l/703Hh1w9Tf69bFVj58Z+oKhbyALQ3tHV9nkYL
TFhU2rhRkRJg05+/RXciEfxftW2VyvySU3JdAdAeJx5aLACvhFtXQE/h/iJOfd91
UffSsVAx8EGYjmoQ6mM+jtoZIjWfqp9yPidSasskv8ASKu0DAjhEfgQmSAP4/Whm
Gotj1aCZoZcNFhFW0c7eVRqQNeC8QRLenfC6NODKI0351Az+BrXTbM3ZKYVZKHa0
IBoaqsE92PgUJazKMB41q6QCA7vNgCUnQPAhNe4FXm1WsLK4LukYAuKqt+oUNgoa
1AUHOEcMVtZywFIYmz4VleB7+9UbQJaYTZD+KxtBABPfzbRU4CBELwpaU94g32E5
3PSlmIrMVtuVfRZQj7u8Y5MF2jJqDG5WL6VT4eB245sKSdIORdcvci24E3y3e4QV
XsoE5uo26tBnWCHMf7GLpw==
`protect end_protected