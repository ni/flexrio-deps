`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10368 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
HdytKcppDjja7VfYQkCqvOxoF0fjBeVs/iYvAit7WLR+DVCdIxiZlfjLG2HSEJsY
lUy24Nc4DROXoWutwfvdWNfmLQo0b0AGPygLbYQ3ydlZxMsze86uF/bt7EnHdKpI
cAYqMFAX4UUNHB3WwYVKBAKYMzjZdBdiPVZ7nHd9Jx0do1p7IkghKuWlE4KLiW5V
gw5EvtaVtrEX0S9QtM07Im1b9oQ27d9souQGPqf50bZ4xASnVl7Ex6RUOgr04d2d
2oZ0cF2WWROZyochHp6/oBgXdN57VbTAvIstEP1Azg274QLUqH3JlqXQedf8XfpB
MQ/4TChRnO/XsDhh2ZEDvoaeuGk8MuhBx+ledys3ABWA8R5137riyEQwO0u5jdlB
amAi/AqMQ42mQm4CteIcpps3HlDVqpX7RKs1Fm/CBNhkCb/heJm+EB+1UwYGkoBs
42n/u/TbgSwbvvZpuK56HLkv/p0gZj3HFIyZV6tw8OOh6S8SmEkElcPYtP23DVeV
BQvrpYGPDTWYtmcg04h9RbvT4+JBtJ7Oh+9ehVsn1V1JgGc4WYk2QZ7BEJzhu7Zy
c7wVc7T+uOTcGqIDpdX21E1d9rzP6jIfgJVfikN7OPGLma/H7eeTLo67QQrNP0Fj
RgK7c9DACfRwJ+AGUiYfiu8s0k7rZG9FZtjAkEY4X91rOgfxqjnFTZlkICOPOi0y
bxcsN17jXCSwfdvHxmg7ZfKSNAAXQ2cEFqQecAZaV/ChYcd/sFerhAFe8708sEGV
sG+AIXAKMXVjMlwePawkeQnqbXkkI/tDPGZrRTtw038Tmzy2LKyssa5xjt1UWeTy
pwkU4MzVLD0YUp23Muy8Gl3xDxghi0FhmDxOSog5o8K1OH9CcMVja9rpH/d+qgGs
8lKaZjntAxoNVkKQD94mW2+6SA90xHQ3mao2jSCW6uXN5geszZbnHJAL+aZbFJ2U
gXG9EVMeunGkIHaMEND5q0Z3O9EDRCkJL1qQnNJsTBGJhrmvUh8CoB2NT8hupvXB
i4mBqTQYGhpT8YIijhEpujIdkW/bD0JJCNDAG8Y4fNR+Dn3pggUuj1Ee7POtPnEe
xT8PBPF42rCDJYhrCpH5vFAycEgSdsvYcLHi0xikViVkNLs/nOGOcUuwsCnkvSr6
wa2URTYP42v0GBWdZmW9gFD4+QvpXLVZvqRl+KRJazFH/yRksMgDmitCZLUbv/xz
L5CoBpcxTFa/v9TxI8DnYTwA6cK1RxDcc9oMEG4LpoyllaLc2M4lKqbS4up+twnk
dNlypV080GLvAM2R1Q7/WUAgOJvmGhNrJttEI6WMbVR2ZoTA012asUYkF+ltwnV8
2R7g9Vn2Vs0HAH1y1UM+6HM84juk4oUjQ+P6UzT8YYDFmrjyEg7W4sux6asyH4xx
7m0XNY8/jYAK6KXURP8mX+sm/bxcWdLA5ywCoACUmqNfIhAtW/TMnUp96HESC0fL
Z8yDv63p5AVFHj/h0j2i98inBXnEJNQqZbhSDn87PZ6HgbBSeUk6gNK26LDo6QKj
tCCyYVbGGy7BtCwcaUP8/NkbOnb3BUoWoyHOMg2DLU0TzVhQaqu5jhqP8XzIM8bz
a0CwKOLjRM8c24iUmUaklvAz4rW/Ky+EnJ9r7XZtJMA+lL7ajiSFEFWJMzkvhU7C
AAolOBpEYTzpNTiTCySsqzEj1YsNizzjM8JXXMlvXQUOQBIUqJWgcJvN9Y/V6F+g
rRgCrwKNZW5mxywjtAkcdNHGBAGmmYTtbtkNB4HpdwAL81iaT+SMGMghooR4xHjn
fcQ5tWpPKt39W9fGJtq086tejQYaCssMENFrEsQQC4sXJuf9IkaeuhL2oEQNTcty
r144oDzcmTwUMZChL0lI6W11tPNpK6PjPqDPBJ/5t28FWgYorC3XGJk5CKd78kaV
y3veG5dRyrTwI/QK7Rt4TlQHOiGVX+OfP5rH9OFJRkEHcc5xc7vrhQk856Epxfft
DAUi8TtV7X/Y+TyfKBmyzbKw88/AOKcl7bHkAC+tK0auqx7uTjL+dhXLGYhZyZRq
cwVnCiHC/fzJF9dxnnHqkcg4zToqlZ6jLFy6x8hbV6rBxclcYXU+iO+QTn4SjcP2
0DeR2vXhiKttJeRLdtlVpxdzZFfbXGaoIgN0OB0DbLyH5IBGN+KrxkH51XdZvktS
IE+YZvaCcvgSiC++ZGmYbnNng5oAWL5CEtpoTl9L2n2PhAzjdUKfQnfx7x8Vk1IX
MEDd393AqSjHpF/d1tnxTwDHyP3hYMqjSM+Oh/3+d6y3Hj5gB95ZFReMr7RNrceX
2+ltN5VQVfmQMsgkifl14/pvvThjrHJJKPpmVqvWH2+ghW0PC1+z5csSUn2iMhUZ
ey6HFmF2I+clqOfHC/PY0YqK5l1kC36Z+2qSr1Ke4Zo9diPPi5F6JZqgtCDfJkv8
MTpf/AWxHdKz8Q8aNgc7f/FQko0wTV44ZSMy8gU7cx6f9IEEXwi1bU6KHodnW6KQ
6mBBR3RDzcYzvnDl8zY+zk5/MJ7Jh5hxIDDOsOXnwJ94IHIaMFq5Ub8eEYFoes2A
Fka62qv6z8V4RysujVKofsUkrqUmC7U9qGYFbbzY4dmspna0Rbe/81ZRhmqwpiJW
wTkZ9Qm9AYaqCDt3GJA7UesmnJ6wb7XoWc1oDNvdpbGUZxWG7oltq+2DpUbzXmA3
OXaFe1CPq82myJST7lb2Z7m6GS/ngZDiBjEwD1+xwySOOj9jLdYrGxb+AA1Jg8bz
VnsSI6bxX2I51Tnp8OaABk2lwIMpovCVSN2qrI3NBWuTJHVHw9qdl//ML558cGoc
xE8hgR1QopjxnBb1qdvBHkdksUzu/mUNE1lkW+JOOM0i1/UccmDSm35qU5+xG1S3
UHQXf17QoBuIwC5B4wz1yZXDVA8JujqrD0DfADHE12X0yNUgqFHJlo9RCtFkg2Ne
Mg1fsUYPRInG7JVPWRM1lxsYwCtLMGcQ66SToT2NvM0HM6xxLjKV6TkxQMOiRjb3
kCUMOBuL2D2eGdCJbnC9hf4Zbjn1AbljUA+webIkXc1xXngEQSExHHqSFKzbEjn4
S/d7aHNt3A5DmKcvO8Y5OhQ0/tqCVw5DTv1sJzEivrANSp4gACmERsr0+RBSD5hr
did55KNhH1IZj1pmYb0yS0WnN9Cw3Z84t4iFgnUHNgVlP7W37XdBK3TSPcuW+VvD
g9I/NCZKdhakWoUCOosCxqeAs8egQ840+A35MKpDfzsOA4tOZcXlAFHDg1IOQap6
g8UjNHEQn7BvfWA4iNx3DAeLOYtPIg1tccyamucnzTecVcjvRt3/9bKhK5K2XfcU
xG3NdOUpX3UlFV1WA2jTgirWNWiJ/X9hEFXWefJRXSouh5PsbG+n2y6sMJL+xhq4
m1HvuYpDhUxv6q688036GwnULQI+Z1A6ex+FDegyuOeEzfdCaNAyWsL73AygJWHs
bSMB9mhCb5wQ6RifgD+U7ysLPlq1BTIEVN51UdQdomBNK9SHIMe4+5tGLtPWoH7n
N5Ju65Oiyks/7sMNvshi3ot2Unhjd/vGgmd24jX86lZPPSZK3xNvsuFQbvHg99LD
LPaZMnR7MtSOmu/16WzN8Ewo8UIXBv/5DBvWUw0UOW9XFeEKTsmE/ryNL3cEGsGy
F+/bkkbsZ1FXmKqzq3oPsrbajKsU7av29FPj/m+ljPlFcZFS5q+4kV7j3cl9fHwP
3vouBJe6VNuDJ/1Se+JZyT35P3qNKO249VdiX+H+m48wGNxc2ogZHPoV16LLmpUz
IfbO1DchYcpRQ9ZkcH/a6ie98Yuk6yVmsOKDqZFxCRBiKyp8gETrm0aluIv7h7KQ
2L+GDsvlkxnsqM8BxA/nkoAgTG/TKZZVrlRScS2pmhMNwkXJ0bJRyInNAVc/CC75
5rnJqMSAoFWGmND0Wk/iGWsNhtZNvCUPv3PF4Rnj4FaiNy0CZsYsiCJUXZ4FMARB
YeOYORoah3zpj6acIwW4Dh23Gibhgqrr/GdDaOPmyVKseXQtxuOg9zj9JBLM1D1D
Mb/LGCDhXGwIoSJEm8J/RyovVimqaoBBHW4+8gKv539+9J0/4PoTVKzfamVkHBlL
NazXa5Te+6vBbzCSewDmgi0PPC0t83NUAUOUAneJn9kKqUKKpy9e39RudXv6BgWQ
e8l4xGsx4WzU/CSHuehKmTBXgOx8a0jOCi/cJ5jofLuj44EFuX19t0IF0f3f4T8w
B/drn9s6Umiau2vCwbWlTB9cfN4LfHaVLvKYc7X9Dkmow6Fkb4nqMgiFwnL6Aa2Y
djEUMAtYsHFxzLCBO2C7rUWXZ+dY8IyKD1G2x4LJ8lskCQQF2/+ActvqsuCG8ucC
uEtCT05B5IMtrLGxa6SUW+7MX4WuC541FmDqThuqgfBSwXAm5KtTymG7UyAT4iUX
4Fwsgrr0fTCz4U3L4hdPj/CTWDraZqD9yQqfUoTm5cEYEtB6h3WnbLeLJrAb0H9v
P05RDDV5BImdQdYn/P6V2fhmHi2uE29f3+a9CuLJcBF9zH0x3la5vbthB7QPRvki
A+XUuKEP6wu4zu6kNEj4VuBgMbPlXE3yqFleSDpO8+MDMxIGZes3F5iWDQss5oaP
rXYj+LtX9OFYMw/w8FqHrzyG6addT+i7QvNFzL/OTY+jsbPgOc50XUk3AAFS1K4Z
O5p5nhLOLhZ3OFRxt7vDAc8pQFECaBCREyM3e8TDyKAexaGvxaJJjO2oillebh80
Jy9kXAgu/E1U5rVFPtxS/Clsud5Qx2dux9X7yxMbdn59qJPz7YKxRpnp/kxHuo+g
szBM3ROxB8h97X9rgyS6XaCisb3H52bbFtQmi5JSjRYY9ROOEgDXIPoECB5jw7pW
1PjABZ7rtyy/KhM0t+SakVN8XM0k/ovuUUu+2WgUKYFBncLspIlareIAnv3O3uv1
vg6jiQqhkgBmDsd69Tbpi3R4j9blihxuvWSoGTuTkc0SO7+9xpeVFHM09eYV0qSz
5Ezz17Uy+XngpYeBBMqZYxzQFyRF8NexhABz82nyzPEDSXF3FaRRquBrhPuvwXHu
c+KKb34Uzm4C0ebvfGdR5qoz1YAkh1GB52we4/bF66v4yvZ7a1E2G30opQgTMa24
HA5FSnBJXYEv99Swjyn3UJ8ZZdapdNxohfex1HtYCyG4JMCs+LqTNSj8TNr554AP
mvujKS28Hu6MZxNsfgv4FNmI5AqYqydPVvBPn59AYPZBpPbO4xACkd+1NIETB1t7
tYHY2FznPZ129noZgy00ubBDMESy4S9mqmadOcFJxoiC4kyx0YRhwLQZ2J0qQ8LQ
hkYcZwRWV3e5xprGftlBPfB8I8eYJn03MVXVV0P8rJkhhyiwsXruHH6ejfrsq6TV
hS20SdSPIRiNLbPGpphE31om8E38Jl5RvczChOBH4aBMZCe7VOGLX4tfapsTGE5j
570ngHLmtpXWL3d6C8jeLJFpPC1jJzkjVSQydp5zU0oz56LNlIJ236uIm0ETRzcq
FaP+0M+rmTBV7ql2jrql/Nob4o4fG3VrgarwIBPTDXH2mZlkO4Ux0F8GXUDzPAmF
CNDXmjK09i/QMNZM1uKnG4PRju8jlgx1nLBthiaAZXjFyaOzMGGLbRl6wKzdqYSs
tlzlHKj21fhQlC3KNb/+jbFtMeKhV8FYdOeFpvSYEmO43tlCAaOvzQbgxUAOoe6s
LAsrr1iXZNlA7w9X9RkcEKD1GcM6jwKxl/DkO3ImV+C93xaCAQGF7bWxERMeRzUJ
cZLQOtG25QOelTAvX5JYHomdA96RkwZ2kZDmG6FjNS78D4+oeENo1rIs1w/f+5gU
2fsh6JuFt2iqtvHGZqUQIzBRyB809i0mimE5/3edDbqaRPhZuUGnhnyprCA8+BNi
a/38YRuedxsmdWJdWA+gRK3YiBYaGuZx8ZxLc3LrZ9wRMhREJQrUj/tbyuKYMgBY
yOif9wmFFEGEZKDU1GFO+K/hKAaqHCaQSzjXrnCxYrAHLMD4A68PRrh/IAnMnxsk
2QVpA5xsbsckLNoBP7PPzNFFZ4PB7RR26QNvmnuTwOX3nIWZ7Msp4mjsGlzH/IDB
5USU2ILjMzoLAa3KN+iy4GCnWLOm8eOIFaJgaByXC6WsSHdftmwY99kEOAjc62wM
7BPRQTUkjiOVRzs8ujpinSmf+S8WQI69aWZhLwSVFxD7CAcTl9hLIImz/rnjtQDH
68/NoLeevDce0QG53KZpBdZZSdyvFn/XCjVK5hKaIVPtpBaw/avfp5SUMSbO4/aT
dkDTpL0E/Jah2ke1fL/kRRGo1E9YBTPhzynnPgK5FYanzjLNwGzmdS87jSeuiSgw
wu1YAN3N4C7aTR8rB8FlK2TSIDTJHy39hsAAT/cp32xMgHzz4D49ncYdcw7GpiQY
mOEJ2+GZY7BgJ//zwjsl26IvVRwrnLtZicmcJhzesHe79kh9WibCn5bibHkaGvXj
O7DJXLOn5OFwHQpRC4394WMltlRuM0RBOIttUUgAuBeYACTJ4C3U40W0INr9nFCn
uYt2+heNiT5rjuFou4anXjx7uDEJPVtaoeeUV+wQl4zjjJX2WrEtEnEWzBoFhUaP
NU8bw1RI16W7FEEpOuxTsQUd7HrCjSF2khVjzyO4sJhwwc33qQW6JcxX5jEqG9Xv
PtLUh8gr9J81qVJTxmu5FvdLv7NAtYkKc3+yxUObMxJ4DBnyc0jQJSrGe/sIgA1g
NfP+GBCb8X4dHEPpQmTahSKG8RQCtCuhdTF7W1sm9JOxC1q6VO7Ov5RlxaqqFqJ8
vphj9jUiiL4kzZ7j1oTHPRhq2v4p6CeVS/TPhXkLC54KT2uc5SCzkcVpG7dyvTYB
MulLkSYQkr49aNd66dp+tps3WfElesJFx4nwcjJ7N3oHahF0G/6Gb9t5jSy5HZU4
ecuf5ilgQsNTGQDnaDmbBGUPNFA+DMdwrnDtZvIVb1IF2luiTM8Qx6suyM0c6/6f
ChM/ER59mgneAV7OJ3IGAg1jsWYS4/Ti9QPtAb1Ug+BP6LUXuXL4vJAAwcc/fewo
msE+SoUZ1bQ59S+uD0exa+bqWsbBiaemdKDSWtD4F3p9RiY6V83aWRthPDmnwMd/
su79iuv21k19Z3vGK5O9OyIo9XJgR5Tcq/jsFhLmoVF1BnaoffsM0itUXtiNmXN+
tfJIbmBl8sXRpnFyVNOOkkxOS4LB9Qyv7n+G0t+LjXs8hp2jjWNTw86L/8rxdy+e
YUGo/5BqiSe8FEfFomsJ3r1nHiqufC6p6PzrKiNfqeLqudiIsDOYEFfWbydPc8/D
T13cl9LbSxNi0GmCCzq+ypHtHt5FfU4gUfNirB7gmVN+0pjPS6dPXu0R6Yi4qUxC
JXX6vqKSeAAf3Z9w1euztqc2nurHEVwSn71mPyuXM8mr7lORevbtzcd66qhD4FqW
YQjFy2xiMGSd+cmn8z9lj76II5OR0yvI1CzRu4ip9vQTjxB7bQPoNEQ0KJnEaGhE
js4+b+FvcqkC75GIIDw8KYs28KcfeSpi8i6pko7y2BVQ64Tngn5OJzr03fG5RXZJ
+Dkw0RY+9iRmycbrNLr5s4zMwMtjCOXaWFVm8uhfKPuanmF2H/bRxL7mDibMSByd
5aCtL3L5GymDnG/p6gzG/j0rOB2IS9KiD+5EcSUqXTJ2vKTlv2DVZUVZxBFimw+w
bCSxlgh3kPyYB751Uh25oOWmlhsXDA9+rn0Lpxr2mbq8oClhjYcqUkfN0fyHCQMU
Pu9qhTNXazHWpT+Pe5J6zpg+eNvlyeO/jDBZhMpJFf8oP4ILLdUov3vcmmCNl5CV
YzB3F1vE8gpmG33NWySWrCXcMtLkPEhB7BLKrtN/0kINsdIY+3aT+w8/u6Wb7Qdd
LvbW9MDmQNOgyCYUz6HVyRfopHGkqHx7X53Q46vEYt5/rTSELIc+12PLrKxy5NmF
OkKLLVwD49Sv38CURHHRol/oqgGDY1trglqUijRHVD5r1xIR6jIMsf7TaXwEvq1w
NgtRMqN5cYYxmA2l2gGMAHPy1S4Wlvw1dK8/5ZGsTtqN0QPPP8s5Uog/K5F1JAwc
8UPXpNGbX1DLPSHEIfj7g+jw+lAss8Nn0pU9rB/oZihkeioCvkK1TfXxG+NGGkc+
QmIzBZqc2LHV/DVtJmn5MIUpmfzkYaIvAqvTLu2+dNRBVWjh5qy7gUQurUq+V/4b
75Yc7mNsgnxwx+64c/XwQWWQ5DT7Q0FMn6wNyIYAgDct1eYW/wWhIsGFgFJlGfn2
xZ3F6yFNKhWpoc9tpEoyNYLPlIlh8DNgHoOYwzJ9PRxFBwO/f211gYE1VRtWprZE
nBlga6n0pkt3BIhSuOJ/JPRE8JnGcpo7E8vy2Zi5lSnE1Cu4+OL9E8KxHJGCXsPT
f10xOSURWGX/qJFF/mFJj4CO3NTAhlWZQQ7yiCt2ytH+1EVkINnKPAldRRkNoveX
FVOa6v9i27RLsruBLv9TCLLTtNkzNt+Yf36Ve/abzVNOOt3qI9a3YXTGYf6VWDXi
msBMDZoVoz59V6tSOXdNuX2RdGMmVp6Ber7nBeq5yiavCs8WrL3KcfKDMYY5QZ8e
Mx26hMsoPeMua9lwcAa02EGDx+x5pOfYV0PiFIP7tPsWETfj+k0Wl3Em5dVzb754
HgL5v8DwFIxy8Nl6u1lezyqBv9Au/SnPu++9x6016t7L62Nl9y6L/r1Z2Y6nYRTm
czwJbxa9aNVaz7gKIxY0pYpEwygA6Kj1jFmlCB+FTP2g//ir4YvNkxBtC7NA5OMV
G74tTIHuRafeQrpdWCMks7C8rxJyWGJ2Z65FoQDwpN5NuUk1aSPpXXj4OlsdZdN5
WTYVQT13i2cyWzGhnBsvJHGRhGhCvsLnOK4MbqOu9RGShFXEy/An1/Gl2mgjJoDb
H2Yjxzczc7ME0i+dGsOsw31Whx84019z6Uid76G02zgWDoP0hRHVv/3d3ZN6q3Qd
+PV46XhMw9WGu8MTda6dSlbDpqS0e1nDvOwqhNTNy9qNgfNKt5BvHkubPMC1QECg
SoyMNJkp8babeIqvCkTq7rq0SqwLW7YdTrcbLeblLB3Tvio7YKbVt4pdPcJQsngO
gTN95mB5g69YEo4hFXkNe2sFz4OPCbdiCmawsXpnD1w50uK6x2kYCG4LwyJjWhds
iyx70mX8p6yAy/+Cb97QkKesIh6CFL+YX/RHNl+vbDuy51M+sh+34toEKAzXItcR
Ql5ebYTVA0n+tVJAhiNt09LURQgfuzEJ9GVpilIAzlYGJZUR782HgU55NC1KISvj
LBh5AQp3NGLXxdUOogaNEqYqxZo3ZdBXIX2wDl1k/ebvagCOOAodZANRD0/rYRdO
+avwOPpD+bYqAqQz0JByUDFwW5wCnFOAH4eVe4Z3MM/nZlQN2hQ+Kb81RK4nJ3vl
qAQNVaPpg/HMfwC/2YyBQt9uHxwxL/R4yWEf3OyXaxfNncLGRw186cbfr12yjPk5
owY235MW/EQ7LzYPueNx2H6Fu90OPo04Nv49po7dfOw4pbwrYPv0I6URGMY5tFrY
44VcyQlPNDKcKqtVBQDIQFo04YMcTnfouAV4EptXrC+ZjdVLhpIjJRBHRzN2T0Wv
pbUyNfARTyJZdBZyfT1UZF61AFEzH/qTlKxGJkRXaCSdTpJkvseTPMhsfB/UWJpY
MCiWPs9NV3fGpD6vWIZC2mJsOx3QJDWpeCNUl/SPdyUONK0hsKU84cSeq7zw81BR
t3ilZay1yhqvlazFmgJjq8HUVW1ZVnTDDQ/RELMDRYZdnqRleFFUaD5tILhQIRjF
7w/qAFAHzVssPvFkh83WMN9HlTmAiYLPYgqkol56R2w0dUvdGLOHFE8rNTmwXyjm
UK+CjRNzKQHRZn2tjD1gNEZFHZ0j4q5dLOMly/to22MpXYDi+4GZMM7b18UFK4YF
2PO7b1h6de491i6Kxek3o06VQlHCCbgX/TpACWOAW91k1kJ4ktW8bQIrc/TijFEZ
3PnVBZ9ktmGidjK4B0TaGWZqJSSWIeapMsYsCXLqK4JnDZe+6c6ooC0amZ6P12RG
qqgSFuw1gDCKwQTFaBLoz04+7snVqPyuwgv/4ZkEmIdQ7zkMjn7VYZEBfRFYQzR2
g/1rszzEP75tR7gXBDj9rlbHKcV+bsAz0j2F5G56CnO7DhbL9LPxpvPhmUu76pz1
stEfJki6wkVqnHMbzI2SRkR6jYVzedr1hzb6DfPePfaSShZ+X4lXY56PYxsICahc
vH4DlzgxHcpJt2N3tiBuLw0RjdfWsMEOvDWIM2Kfm7U7F440vgc3v8g1JigKBtQt
onP+jImeMNlU18BpOd9dJHWQr8e0xrm5kXR58IwJxWTpB6beU4iQnbZpJycdBJM8
Ri8t+haParNqx0rPC2SchFwzwy6zup8cCX6oNZ29ySZyB9f5GcOIOp4HEbLaq8y/
wWCPnWqSWoFT3kFR28ky3lXjt9+J7nSqcHAtsCw8p9rwEs8xitCdRn3xjqKOhw8d
GRqW5NcrUKoo4ThYsYQozzRxWahZGcGekV4CUqJB7iE4YR6g8bf6aYFbh6uFgDLO
D3BF9FEz+3HCTpiMp4APnRZ1bA49Ww1A338rXiHpPZ79T23mPKoj+CndIL3PKMGk
Q7GeopoVQFtfgh5xRVFiNIhkwmB+pZBSg+BazNehm7vv6hlAOqN5IqtniAceyExR
ZebearErCll2WeNZ1i8HcMLbIaEJyf9nYMZTgfEaPWe+djuNX69piG0KJonhszVv
d2Z5Ko5EjFtVU0ZIuKXEBaEP0CUvdIrNsdruYf0jTttSp2W4HdmRUHJDgOcs/FrF
69EMD+ymH+YTKq4ChlyEAok+Uy9NoFLXjdKoEbE3Bb1CFwkcL2uO9+BBxKlY9J/2
vpz//QyVUaouM+DwYkRBx6gBtp/FGmu2BN+zllIwVJ8ts+WnniE/08WSTZod5yLE
38kuWR1Z7D/X5hI1N0lt9jTPeIBGAcu+iRmhRIBVnX1D0Xdc+UjfjQnT66XdlpBu
C5YZrArU5z99k2vZkWVbpEoeShqrGAl+f2NGAuleFjd7+MmTLIYTfev3xa8k3fJN
/PmL7dJ3UHWLmXTwqx7dmcaEEVgj/ak/mqbPu++vQkEIuKtHzJ5rYIXVSaw5RzDy
BVXVsqEXpRjYVkScPt6ACcQPhddxKIsxYe1EX0kcfIGUxG2NwfbvmOv4XKQrwe+3
fNNcySmM1m3Z4aShljfeLbM87bNdYKxrNVh+g3SQpgo0gdv3se+IiVq+JixJ6ofe
FUoIwWrV6i3r43TK6GOeAFql+6OWqoTHQ4j83m0CWKuh20s9gj0VZyW+orsQSHCY
AD50OJ5wNOhHhuF+KXMTFjlygB9TI1+sksefuAi50iWZCDlwyf6MiBP5FBNxpI3V
aMJC1ZEqGfZyxGG+Xp/no1kov6IYwtH8GUmwcaCJWnK7KDU6ZRqSUceQjlGiXQ2h
I44V7py5CYDZolE6RMgt6loFOwduPlOfdMtcoVWKJII8V5EsESuWyqdYvyGmIqm8
lY5NXSG9QkwLksVJXpVTj7Dnadn+DLlvZ50tPuMGg1y7e69bU2UF3nKaJWyhzkWH
DyEmv1ndhaamkE7PvTZT+SIAs6Z/n8N58GZ9KPjrak5uO5WTaAuqC+jISLA9OzjI
XyE5Yy8GX1dL0PftjijKmrn9QdbpA0rk28TlnwqqbUF9rmiOApUtBYpx3bK1WGCI
WLEkooZFqaJyhioie4+FGMSxgkqq3AuKSkviWx9Q/4DRd+S6caYJWD3yLjT+CJrR
BFUnnQHcuSq8oDJVJbgbd99qqThAcDsfb1VMZICpqd9qDs8ek97X7znshawg22Td
AuH0aq+CGuNon0uwJyrtrh+kf1DoSBrs4gjiRm2EkeIckBN+x6eHARTfenrMEpBA
LD7ptYxrdkVa5u5lpbZ7bWFVpXuCbBkcSiOCn0Gtp/w+24XXKWo9BLnZ9c8Q/tVs
k/oBcMvBL4ToVgxhDXOXy2AF5MU/x/3mU5FEG/AyrW1cRdAuvoBvO/AyMZLpAGN2
KdRpRMnGlR5AkfYZMjCWsgr2VYPr8g6QbFtY7nP3VXg5wnNf8agIjc33hS428FTH
MKW8UOjYyH44JeFL+pm89kVq8NO4tgLItorYuAp6WtCBok38ml/TVdqUvodxsnD5
AR3/NyWWW0bVsTs5PRISp3/jOuRq1ZphYT76ADAsbaNZR+7fM7sQEHJ1d4DuTIGV
BxhGAOcZHAKzQxemwlTuK6B1CeCvRV3sFr3QdW8Fh6WpDWd/KV+ZsIlGwaB8JBAB
I34VIhBnJeTDijRoxeIx58PVMT9/ZDmJJLWfP1OeZal5/iJeuZWYyexXzam1qnFA
KXbxAF368nBAydlPoQcnhi7nn3gsD7j6QI9YbIwWTsrEUeU4DSEof0K1QeAIXgEo
1+sJfM7Zz6+NE+kBPydGTYwLCKkZMMFEeICEuzYvJ6YakquO/GlCJpx/dg5SCM/0
XaeODBc73FCHx7hPFtUDCi60xBGK8pRENulanNWjLHWthK85HofQyGoD+34HT+5D
XGMqs24KRRU1MGTE1iUm4CGEYfzgK1fKRXLy1Fj1THHv9RT8qgcNNhkPfD/Dd0oK
CsGg1pjupvTJGh0hlYtvoK2eThA1F+uQ5DJdhM25UJcmoTucKpsPF4dxERKuEhE7
yOGui8Wf1HlF2CgT1vW0FybtD3vpsapSPuf2taNvVgXjWAhSyB5Mt8CYaH85w/29
jBSMGlLFRbyTs0m+s+nZvYdteKI5DslwgQK4eKLLZkRON9BpuRv+TAvaqg2m9Wqz
XGEiciv3htHTkH+nko3SKNUWMG0F1eoASrmYPCCN0nADOr8/ch/6gvhKAa4r32s/
/uxV4qf0NJ01AA7YhRmjU5vNRXyKh0dhPNPkvOEXEmGJBYog5OGAhX+vL5vqy4C9
Pgg9kBGhMd6y43M7c0vA4hr0X63CisFMkmDVSI39hwKurxt2qGqSOz16j5i2okPN
CijkyKPIVyqXj0+5eMDkJ/rm7LUn3lJs7DSkjPMMTqmKRSUbD6qzbRGbyRc+TTry
XQT6FjpDArQGVUjuJWgt+0ImgtdKLoSlHVr00Nu2zVvJLki7upvtIhiIaU8qeD4n
xLjdBt9eG5t+lw+ppQ6PsdFLgPP4Mn4X0crOX4X+F7c3wmSK/NZkkAXKC/4B0x4t
ZIKDnWCwyH7j3jNQY67kEd2EI+BNLgIgBVBkhRzullsTdko3E88nalCOr8fmWtrv
uGYLKY71bYX8lI0OElvZFir8/4Kxx9g3ryfB/hz0bcHJBVGh3GNEqaNmPsP4zdFw
Ye+496m1Lig6T4UroTQyuFZFKqPHiGlo/cftyydZenBFiHpQzrieK9vtCsrgGCoT
yyovqMOtfd0yHe0+10ZalOXQa/2XAxHUp9ncxKNgoj16Pk0CvB4o7DQ9fYKnxwr9
3cCFladPCfuaDLUJDz+AfF71l5CQurVy/Wqnk2rqkKljsG5LdyRJder4GeVgMtpq
r1zOGE5pfw9+mLxSOU+JeBsh9Eiy6RI5MojNYl9I2PbwbURw4v9K/MdVyDuk0any
1ixGnxfydGaLu3EMOylcLLm2fKKbF4ivMnhot4M9qPh6NXMF3+vzlH6nkaJHzDrG
fPgkXPchLN/dMlPnggaTvHoMSrywERSZUoyKtkh7BsEQpRNx/HkJ/KRqrFka4KRj
`protect end_protected