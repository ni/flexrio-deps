`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15696 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
tJDuRBxzolupxTryvQf9781mFEFjazTxPfIJf5rF9/7ymDrBzwAfvwl2pfBKooVi
6JqtfwdyH/xPkD0XNyLUhP+ZxJQAvBE4ZYHEEdN2mcChMd+uj4LTcqrfEM8Lgd4K
49G3xZrgUk2jq9WIXU0X979ECNHhjUGhP3nB19QuiJjh0TAwwRKMFZMdlsGRk1JR
tMqDcJrSJWOYvB+7D4F4nT1oveEkePJ1nhxxg7jDytUtHwy0kgTFuTbke1HG4V48
DiMIweobkAeg+Gz0I0OxP24CJHMUUpCDNKFSjTkZy1mbyM8Jd4geRBwk5KeAbx7W
QCclG+IevJ6rdYweNpcTn6UU3BV5AlRPxP/0k4xAy+z0RU+7n5wiAfN2jQ926TjH
5KiPcRrYg+caDUwNzQLP7kjVpikofhpT/UEEH26lyTLRRjtVgBoDd1aS05vSCWqI
8lrBZ7eMlu8bAstVdgemvSOx0D/LJi5FgyFaZuek110kV+d+zqvXx8T3i+BDdb4R
5r1/cukUX57ks/2S8Kb/i8QG0+656ivNYUVhG2NM4aJtv59Rg0rLdeP7nmRY1p6K
rNLBU2HWiw+jQSeoSWeuUDtLdCeRr7FY89x+mqjmHlY5B2e89+U0UjCBm1j3n6mt
LyuQ4sNSIbqncBDzHd1wBo9VUwmrArXLuHvdfG8bmpkgl/wqC1baBAW0j2ew/sZ1
Vj9PygC183K1aIgDLmXeUDBP2unCWFi4hwssCufk7qRlazBULlvIGlqQKzdEliJs
Vi0Qx8Y3caG8h6WOwPSOKs/I9KXL0H7NlsFzcEMBMu3C54/XJ/FUO1l5kG8RtNIw
NN0NYWLYjDMRTqp/vxNfF5rzxAOvGaNShf4kad2qs4+Zk1EF0Et92n0mVqq6GRQq
CzPuddoO9qLq1PCjIEVvuzvKEI5hdbBUtzi0gS2QXCNErOr6N976OXSjbJ6guKGI
DPE++zhveV7DCEenBRSXfVTmSwnwBuReBnietF23ArhXSslhpgrUUEI3mqhNtxcp
stfFyGLGzqn5Hy57NiDVXCugbfVj0x+mDPI4IQdiqV/u29EgWWkb4CAUI7VzRKsN
YXe+cpcTlHX3Bgs1Dkshs7UsPtts1cVLX5ow46HyYqCRKsH5oWiAxgcP6KtTXvbN
6XHBfn/Ca3oGnI9x2kYSlTgM2MdRBIZAJuEPc4kRmAPYqVHvlrAgryWuAmU5edRp
GvE9cKul49xZzcoUwbyjCRJ+CjuQe6Zu8h3Z6xrv2OEUaSJm0KX1tCJ/Dah6GbPP
Is/b4Cx28fc8mqVTiNpWXsSMWg77SgHQlMM2q/v/2f8+s/CXhiOqEPhKQOEvRWe7
naakXhHDXgebcsJohVoJeAC46m/l1+DO48DHEV4SaYC8U8mBiCPVxvp7S5sstJkH
5s6zpPqAARirGfSALA98xmySCDjYrdw++n3hvS6Wr2GGkDcSMJ84DdF8TnrknfdY
RtoJo0OZHRKxx05jsQYlWky0j3AToKw0fR2Gh6WW4RltYsp+TgVAz+J1oayVCpvV
CpdURIF+Uk+SUPGiQtGj0pM0lsnUlTXIt9puFyh8vIrwGFaMif/sijiiN8uZrDZm
QQtd7Af88hJy/Kb076Nr/MPwdeeLygMgTlFQLYLKYV0LlmgTPdRqESXrXbM09oIv
yDEpeZ7w06ToMWmTkbc+oH9zdFEA2cE0BX4ZzSNtMLfO0ZbdwfOs37UteFUJHyiZ
eHw8nu6EhYIf0RVLZZDxZ2V64LyL7TfRnav5Oavm7UhjoKik/cCu7V5p12nGxKQU
jRKAPTGeBvZGiVW/GC7KbZ6WjFkde4RtJ1zXwbZgIfHP+5ffEC9akdDvVZJVn/WJ
66pLmMu6rvLczpsyGwcEBUGLqkyaX6nB4zLFnaWqrgqAiaVbdDz6AVrrACmPDMrx
lHfCMNJn8IUIbFtBMNGN6EXtp5nY8Q+RoXRmNKBlF9xMSE0sgeSs0bjhX2j0tjMT
5xQ5O2NuwgDglKrN0wIzndAlJhx28cjGgtG7h80N10C2G8/fFpGcOKJGvqtUTojW
wLlJvmSwLQH0d6crxgxOIqDw4gu1gsuqk2lQLvzzZwLLM859VhJN3Yyv1dAKgnEh
Pb+7cAJD1LFwoFbqSc17CG/PN6DWgwQ32NQhsq+/PJnsLv/pWK9Cdpnud+AS6cPT
fXnkM8lt5KW9kmEq4YrFvLPtycQxMJMQHOD7M72dl2v+TaxM0HugqGclqj4zJjlW
lqCKiJ+5+Fej/HFA+K8A/L9zJabzHUgnaScmgCNSfct8NFAZ6uNWiUExKlTZSL/t
5DJ6uP8vsR8VFodhyK/z9AREMZDaSL/QljAFIztSGxj/DSEz323dYTGWNfrW0zv/
Vh1DKK1dttV6iqZAUxoP7+o0IfKs90hdo8QxmE3qKb4eOXr+GGR/bPQ2kfffwHIu
489eY9hNw6VKp0eiivSfavgz1hRA50NcNkrq8Jhw6o18nTsupymc37NOSQx5iyYq
vrFDEjnyjdfhwIhqHRmrNtz+blXfJwz5bIBWo6yuN8JJoRt+O/sBgoaYHlqUPf20
5LaHKVv/LQ++Xcd5VTLHwee1Ty/+qjL5rMS0FrNCYpm1ZyrDewd2Ih01eGqVqDIN
NerEhXshM/iy4q88mm4maf/LnsUExxKjHX3W1xiK2tbUyAy6WCLtRBYP551AJsXk
gMmXmiaTkIXFhTsc6Oq9M+WO5jhPlXXNGo8PB9+KJdNemUFkZ0m6ZG++YAKPZuKx
xxMOnGAkJPVntN7jx1tYhOHo1ieUZtB99FKZ7U3myAx4R1+xqZcr7oYsmpv+9BbV
I7Me8G2ngAtvg9/HxTI3v0SpCA7n5MUHdEHCrDhAKcJ0mwQZvByidbDvGjcSA4sF
cH1xfSXiwgvu8NWW/0gfFPIztsj55sDzRe0mTzFmGzWgl9kOrGYd6fd6VCD/19p0
ka2e4UX1A0LpBaOIET+8Fnb+FNrO3vx8+Tq85tOu7128d8Bwb4KWxKMFrfXIREhg
Hz5Si8X4CHXfKQceqAafyrdsTJHnkTYdV8f8Jj1WA3vsMFSKFP7tJz3ZDEVrY3pT
HMIFBT0Lk2WB1qgD1qn6I0n8s9ODcRWkNUi5T5uQ3l2Hh71EbLN3lADEeDzwH2fB
qKP3yNuJnvpbO2EbEVG7hgBotxaUMoLOAtmGwrB4AbvUM1xLcHO/C+7g5MNKbjYa
I70piGy1W3+bXNj1wH09hbcazjsYQ9+5N58ZaUlUN79uSQMLU1C6HFzVd5qnaS8F
cGy0IDi31678BD7yaQSJk8piMQ/p+kihh4dKUl8MAH59FZ5M+5hkFQMwXWbYnpys
rtXoJGMGm0w3ZCCKlZrj4w08AcfqDTfKXxNPdeMaOyjw5Ij9hpoBDGw15l3zCaRb
Jj2LPg1V60O3YIQ+QEbIPWNCNDXcPsDAs3HHIr+Wjafx44O/xNtyCdbLUlE9JUrP
XbQwMtANkrbuU0VieC4X4I8uk7Ub6EWTpaHls41AziZkv/sV0OOso5hiWEuN1sVc
UQ/RCvDEA3JcVaUkIA5QL278/TwgeKSUReOZMJE1n2UZEk1fAHZ4lM9YZR4rditQ
AHm5b1ceGZRBk6p/XuBuQhTmDJgxGv/OaieB4H2Ukh0mtR91O+rXqDxMCjj9ndtw
pz6FKTsBJ2dmx6jb/LxL5jEiR3jI40QEcPpUSnryN6Ok9Vg5LNF5jKyY2lgLzb5o
BBmzzc3rO11mKavEWk04ugXnEQpa5Imc85BBvJrustIQwUVf+jjK8hQJrgVt3IZt
P5mKFK6kWSUJriAE40R1F5mBsKUgQs+7Scz8uke643DSmg0Qylp/aojXNbLdiCwV
XlzkV8VkI1JGYCdcS7K8hFZg1rfkkBj3+I3/o3sZ8Y2ERzcX3cOlKXitftvMD8K6
GQOePC4pokEyVpX9LwSOJ64XRQcZQmKVcSmoist28zsWvyuZfBMUGqrZxhFoTeq6
aMzMKcVEAZXni9Ds+jUuRbuCxB4jXV2cP3TB5pznmZl/lcyAJ1RyMnR92rtWR54U
6TY5VVJ8HaGjJ7pJA1s0RrYkn8ZfiNpzJpzojo+TiASDP8oK2ZkUp5wxRlLTHpDI
OIlNI2nTnem2AblvRyX5DiGIiHupT7OYZal3ncnNTHDK8o1pkeqCe5Tlbli/m3qZ
v9fR72KcYVj6CkS9QI4f2ftz1V81s5F3iw/ZlSUfGE5Qs6kxmTaRNEtLMwOEPtrx
Z+TDekIsMec1oGgUUx4HfJTyHMsc6h1ZBSKHN7xIJEO97AUskV4J0tu/bSsD5m2E
kcNkK1s8ghkDRqCfzpZIhl/QzLA9PVPQEA8ws8g9sWO6h9FPYTpOyLrlPcUXVA0B
+XknmIvgCo4VXLt8wwqrb2Rl2KCnls9XbMOTN/fsZmrHlyhSyzUGVYi264nsGwt8
8CKHKbwHEbZ0FJABC+MgB1Lf8O+ZeaiPW/IxVMyVaacv3/za+bLOjERadxnKONn8
BLJRe3uBbDB6HevciDKbnmFz8k6VMeSN9iYHdSPOdFEdFfZDOCNlWrsluZXUrXII
BMVm2TVMPhafAxSaY3wQZWWbAIPdOgH3Dmo8O8pWqx1Qvpgzla+Ybfe/JuQ8KOfJ
EHgVuVeIIM6uzXV8gcsPHQTEXblw2S6SQeGhBJ/DJgkWXaV1PUUSjtEal0N6DmDA
UgV02Rri5cR789XlElcLuPzDdXpqFt9oUhr9FX/0/VGpS6FAffTHdpkmAPEt6TOC
KCqWTp33lbKSu3d4Ktlv3O1q8NxDVaG8Vb/O06RZKOIigM5XJWyJaL8B4Q3jlSKm
icUgIOfcgN4tTiEehwsly9UGpR9vnm07c8n7+QfFzME2IrMd/QVqurEXHk76ubg4
nkt2XF4Jkb4H5kleqsunxhNZHUU2OzxM3ikxkS/AiRalQSb4Ar5yjSTf6yu9zrL4
kGj09Qg5WYO0ACkm0XZjYOfBWsM1N7odc9Vv+e/Zn52aZFFIjVefGVIcBQp92/Us
CnW29eCBvWgdWCD4oGYBfVZZSt2pZjCGb4QEDbttIqQcyXKotcv6uFUT6Hh6Jtb2
lXrGJNVruoR1Rg3uZq/NQfevFSyTGfzKbFU3hiVjb16TrkYdABWvxjFrmobOXw3W
CpR3+0eybqxkrTaxCLERXjqW2AgAjInG+BFuTBc2hYrUuthZw+BcGbQvVlbP/DM5
7rjcwriOfvPvEi8ntuoJK3cSkkrKaz5i6miTE4z8xGscchz94J9oe+NJy0K24mes
ujWDLBLQsnZtkHHO9DwSbE+5n6rkZUil4DRuJErTqikI+LgsqyOAmiv4fFobMdBj
9DuKWjhq6FS60FonBBqf9/ds/6nKhc3bxWjwKVvfXcCszww8U/6SQzUEQwRTnaaZ
Vegk9LSqpLSfwbsGnYB19GNHil77kG2kNvQBkzbtXqNukkqLjmIhH/rIadrnhgk+
q2Qzxt/nX+r6Zoj2StkImBoqp09a8X7pgw0jhXz6JDtiZq3nvpVA1Ni3q2KVBMsg
tD6WJTnWnTIWR010Qh9ZEVjVmDp81NpgJMEHX2dn/4Zq7MsewpOHNuS/dLSO4ukc
hH7CAcByFsn3BSZqXmnZCmA+L+/39qLxMmkWA1wl6HoJF2U/hK97Udyed6iE9m9B
rLxodkQhMWg2hz96zyys8fXzwdsMjplH3NJaZFOsjySu6e119ayEfb+wGlC7hFes
fKe/zejomnTTCD2jv2rddfxmmZK/znQtwiz+09PCUQYUDIw5yB/xgEIDEmgxSRNy
CleZ6k3gzkKgF11FLGja+MdkBEq7163YRU6YKaUiO3V/+d2mzYoIiPQ8eqVB7b0U
xg5DNvCEoi85/jjJLK/D5v8PaU0Vy6ufyDWQZ+YhCI/VauO84YWTDjHzULDGf6xm
Y9+Ngv2IGIA087AbqqahNUFZuLbWgvCV1i6JhCNniJfC4cG3tSRxc3VPHkShXK74
K8YC6t9KMucWWguejfbDqY1axtHrUpQ1gs80zLSPtVcS5jL0aiTF6mOZoL9F9/ez
hina1bXF/Y0rhOOG2Zvk9WqAq4C8Zlx8fM1ELYYaxOZJ/y7wl6tq1sEMuPmJFRVH
YzLXf8nk2nZaioamarIZ28I/8ogKlMwY/fVqwo2eN1LjpWV93JUpGmLD6cjU8TGn
1dUsDetBpqFTqioaSRpqKOJhMV4H6MZqhns/SCUEWZHBcBMHEywOjXPz7ATNNHDv
vb+VLohSzyc8YwNYBL/9tvLfoSOcmYVg69BXYmyPn8I+2vRmBCZi4OSTc3anVxJO
e04yzVeP7UsIsKGiGd+lW8LJ/8hluzCRfcE2btAh03o2zWva2Oa2RDx6WpPvqyiS
MQ+lzPyEjlH0Eop5XMfBO6sEW+XaM++yT8joWszLqC0SsHdAT4pm2zCwsz2fX5Jn
T+9BDJWsOKTsrEj6461MPWfI7Q4UyCf7Sdh2PyqcEHlJSneDQEtDLwe/X6ZADEBb
DcGi4rmE6MskcTPeNjyUZP2v0nYBvBm0Lz7JpwITHzuXHcsDkhvmeIpQ1slzVXkc
j0zLppeC6veYnnBOVPWS+Ybw8hrMZ+FlEAprOb/eSFkpPB8bB8gO2PruB2A29nMS
DmUimJ3OT6ioAH9VXW+yeW+XQ12LGMGk13GPkwx0C0InQ/LhvKeB/wP1rOpZfKos
bGg4H1TU9Ftjm1/j+2jWEyC4Lt4El9RamLzrenEcO/OVqBIV9uRenrZoJyHwCfWO
PIcwHHfnKzXBvJH9sqgcYuc/Mky/Va5BaMXl0snfXFjnKoMiyg1zTlAMHEDV2Yr/
xc4RRI7kay2DieKrPk+4D6A1p7eEVISiRJH2U5O3o7tpzjGuVtnvdBFtRqalODsB
RBvCE7Kqa9fVzJwnDFMWyQYO225PClSvi1kTkZCWljvV89GgPKvEHz1JaHFEskqD
8rR9y55S3FqtAAkCJNeKGhj2vPQkR9zufx+Z1xtSVO8LWV2BtOql0xdvsEhyn2QH
+iF98D5GiNzbHYOoATSBZQbkg8didGUC6l6wpqe6iusuSoYkT7KoHk7CJixwfnwG
4imBEXOFiyH3MOK2QqEZoGpwLzWAkXtT4YxzC8O9ZdYRcLSrgr/R00YIOTbEFHK2
lxl1ljLx3GlGmgY++naffdEGTfeu9O4BTa3Fy+0d+9e6ln3m7RHAoznqYhvn4WDt
LyTW2uP8D3X9MPWxGcOWc94T/lNBBov4se1MtKbH7LBG8TKOYTTXAdIK8cLSpw9L
WAoF1oSV9m9KdVe7b6Gt64FiSVjZEzjcCKgMfAXOrrDQrca2+T9pTBVj6qZQdNNU
MXJiE8F/9fNPlH74xL98RCcFUnyomGubaRaOIT+9WdA3bMYGRXgW2Hi9BHdDgVLF
kDhThyR66UPuwPhcOI0ANN0vYCiLB1SR0fck7JTP6PpUPHz1YlyAC5psoT0XUvOB
yuwMGVIdcRYdCSj+fjx6dmQ996CnedWuYnyKP2+1a7PjOjru9KijKg4+qgwDS3oa
V7Q5XwLqOh5Braya4+qM9wy1WuMSCHkRMpjSrB/hsFdyeR+a3TSiR4AwDPnGQtto
+NyZi04snLUPpTjUCD+xAZUoa8npgkjQOyjRAePATebxCjeZpbEzOCaR46AChbm6
TTdyg4RF+69kQU8W7ebwjqrHq3yk+cNdQbJQCt+XW49bUsdyK+IBtAPcWYsomX9X
/EhN3WGZ9/0Hs7+sU+BUjAQCGUkazrG82Lo3cUIikes00sclHfQXcddVVYTJjeTP
4GFC0enSPUr7dFABFYL1scWYL0mz3n9tB7ugx7wNoJDE8yreLJZctnvEkY8W5t5g
7+XoK7CXmRuiLt0rhn8ZFqzd62prarvmGwPaLRHHC6KHgA7jYJdNfSZboM/p5n37
k90BnP5IXfbnktDWvrIhfZzVjgPOyB8n6OABv3mwkkD2nEmgw3xvxVmW40rUOc2v
n3bSLF/Mvo1L1yLf1jTC1KOi4nD6SipP6kTFs5pGPTA5CYFXUp13zW7cQvlYyFfy
lltGPu0vWel+xkhkxWefX2dDi2gheXxzqDpwTuHMQ9vuKFwBwegBUq6NGJtid+g6
81lR2sSTuXM2jBf8+ZEI9sT+aK+tZWKyZIcdYzLaEhEFelNapexc4Cpp6UQdNHYk
IVw7xmHTKgC8+rTAISnFqQ1DN7PPVAAPz9P9gLfGOFZKks/xXZ5djI7N7TCq6orq
6E1ANe5v7nr2Ceo5zwh9rNCqUKKkOBZKTfb7CNLL2YR64OTzRI/n06OUGfPBse6j
NieAuZr6+9YDyGbDCEBMfse+YTDL1hbzo38raaXm6w3J0w4py7JHuWZDAYap9EI+
DCgWEuQ7LwkDKVjDYqPdgdlsRJNWNWM+cy1bPVbUcbWUjh33o8w61oABnwHmBI77
kezv+q0koNN1c6GU2FQnQZIBAGOoMuJsAu/4hNH+Qhb4Yv7I1N4A2tFn0y+pIdQ1
eYKIX4mMo4QR43wOSGUgt8CTlNVo1+fGF2H0Uk56GKZVGdDx6wNDOZST4BrM0zNK
/4fWg+DKpOmjD4SUTRUmf8Dm8sDLdlM2QeTUOSnWlOgiYNom+wtOrPW/2FHBeUoR
hOPn+6XnI7gsGhxxNuz2+6xEJwwsUNSj1zP8PgHvgtSTT3OeuozYs31zHpYjkvVm
Vy5iBndE3naGtt6QOB2SUEw6KUZdRVIEr3WzM+LNlquEhuTwhy0W6aR6XjkpNbeh
++1+LNr96HLKG81dgdkuwBInu2kAl2U+BSXF3guX6gHtPn/n7swl1eRRnhxEKGxR
hBUN0E4QzALoiMz+JXtNch5DaAFCYh1FxN4A/JK7JPiChJO35NuFyDhE96C9zpBM
rdbLjw3dSBP538L+2G9a4GsL6xKaq0WQFH9zh2c9mPhp58BlGJf3+VQ9QCXlkBfs
z5TLjYKehqF4A5S8ChkdIgvvd10gX6QDkiJv6TR6M7v1/Jmk8U6XnT3Rmg4Twb+Y
hALNMpw2SdUKlRS9ymaGur5PWDZ37MZqbQnmsFvJJcw0w8HBSpP8gpcRTJwoy8s0
X8cMMz8N9Zn84vdA4bV1GPaK90OkqDnIzpc/jJ0z4wzRZHEtYgr3zMufXJ7bh09l
W7UwOFKvFyg4ldOlxIp1eplrmy/9enx7fBBEhAX4M1NpjvnATnlHPYhxCuBoMWLP
VuH9Pl8NG/5MaXJY6cGUSR8ubFNxFYpYdfvq+enNeLW6C/bD4KC6NwKiiaal1sge
V0io+8pJhNxu6VthJiHwR1G44ToXzf1XWu5JHIT247PSy7zdSVdiLAy5Kh33Rmmt
XMJQ/LWfHXQPWwD/Cutjs5vio1MRgaNB+YGPCabsvF/Sup2ZStW5sYV9SHUZw4HC
Is02L9muxInAn65zUy3CVPQmMOD/1xFPDwiEyzgJKNmfTWgPSIhd+lsQQfcvz9f6
NkvodJPcTcWpe+B//qd+rYXwUAYdQO5R1f7YbvHjINekmDFmFS6UF/Jq0lKsH5SG
TGgInfKIKsR5oecjjTg8j6gLH2GRXkVrTQdZ3J+c6hWa15FvIPbT5PKVN2jbHxrF
rv5TLA2GUNDOgCABvZBxi0NjwTFLC/BR7IfcMlH1nCeNgZl5VLRDhhxNZszFj+AX
u37VVImJ5RVlPaP0lcj2vbYCV8aRxnN2T/fN9tQY8dNuHs7HYHlvW779OEz5+nvZ
/ZMAqsnsNzJmgkZi0XVFpdx5p5q5H3eDVu3TB7uA9KOlkHXr/x5PWrxfVcoXNuh5
Z3SySOKve89HLO3Yz2Moer11EhwO29alw9E3Q4javz5RRh8NUzShLbFfLDpN/QJc
JpgbNznQYm55JhPCiwU1sw2l2beG1k+vSzyc6wC7sxr5C1X2oLlGf8RlEKFeczx8
wfCW8d4gFvLEEmfXM96ht2yhEw5BOVwDsFcHWah9MhxmNgaVC7BQwsy9Aiz+154C
S5q+2QVo7R/kkqUyXnGy6blv3MD3ANrUHHz8YKHslJ1VZSfbC5Za9llnO4cAK4Oy
KcNpp6wYrRfMZ693DFa5bKYw9IDD0/TemRCUoERTThgt/s2m71rtf8SW2Enz4iw7
NgrHwdT4ohM0TU/5BgrxAhociFeqVRjT4WOmfItnqrGzST+3DQ8pgK792Dy/vnPD
jRlh5kcsjS8/REuzrMFDGOWzJDKHZLCpoPD974Wd8RWP6ZU7Mj2km1YD9tMG2TwS
Tc0fYY+gpXj5jpF3uuHed4krW1YQXra3diJO0fDkO274ZSXHu8dHLNrqKLwN8t4w
niPswEWjNWGnQ9OoeKyox866rbAx+W8jJWyrz5msbG3W5gTAh1WCvsNXp33jZbRc
eFu9YD9a8a+VsEkXvm6w4Ah/O/DdjzCV1wnGp6fjYVMJtnXt7LJNxXreiJYnmKWv
EcQRy35YpeTvqi4CBY+5zaI1lpdiD7nA6qTH8P8i8d3kYTTC6lkNx618w+rzwrlA
S3cJsoMoXUlvUQtepG9tfOuQbMjbyyKS/H2GhBupd3ehlKJOzn5/J61ZlVhxBkn4
s+ioDQFe40RxVqDJ88tX8Ge1jyDEySs5wUfv0N0rSRUDWnK1B1j5njQQGAkwHE/y
OVXJC1Aljh3qWZ0fSe3OG63TECrPzm9c5F7jebQ8K0imJY2HN/urJb9dkRcrEcyM
YYsj0kmH0HszhXMbYvkdHoHd1WpVGorSazmeLvnXLfSDZGjXTocNM3KH0Vu0J+ZB
vKqs7jLDkr0BMVcfMSHWjnzLZNakrLCdcGxXfjqKw4pJ8Hn5wZd7kIMtlU9Jy3Sa
PulsJ1MI7IPR37HAUgU2GyX+IaWP4n2qvSGdtKnRlR+suW88xR0jNneuZ5KnqhiK
EYoKsa5dxOuigenHcGFzsE4u64R78uQWOhVg+v1ed/vq0wcNDvHgKxTFfgRV3X2R
VpW21HaYpe5GfDFJyLOCtbL14j2ycZfAkOQYMOUo0cwwCcAqiktqEtXPFnOJiBK7
8EE28lo9DeEjRhaoTn19wJ8V3e6xlj9wJyrcrpnAdMhyRooESIkmQecgMh3ydH2/
sVpcEKBPtoOy4SDskpSo8MEFH1lBt7Yq41cP8eazeOdhmPKm11QyWUQcKUwtbh0n
s7pSVWO0Bcr3o7VzkGugSjROkwj6Nq3lIcETlZXwZ4A1GQZLLxZImchKD0iNgG9z
367epFrjg9S16/UkKoWh8CD5LHy5LsFpCHVjhRiZ03ZH3nrNs5TIte/KV0vVfOCb
aOfe3ujU6BU4bts+mXK73gu6/R5yIPlzy0IjCyE6LYhN6MPkob+61TEowtw5q3Cn
833jFiRfBBbEyHOwCBqA7YJjyRA7IsD1XEfSXyVJsIGdZBsHQjT3sRg7IGtdIOUM
kO5z7P2ffELoqxc8KAbcAZCQYQ2CmQoxUdmNOMNj6GI7IKE6p6Wkd/ySgdW8CXdS
laUnWEe09AGO5jmKMjwUamoqa6VkOmBAz9jy+0JWSeiVgJr5A806SN19DM/EW+qr
RLK+PZSfmmUUFYVK6CSpD6aSFOrUcfN/2Jje9k/odWT/elCxTskKrU0ZZjBkwH3Z
/EvhA82t7eZUj3FD9rrBdoN6zLeqR1Q0+Th3klUMK8XIJxb2/z4cOEs++UJAhQbN
fGn/Db1FbM/BBWsrD44lRFf2fvgx6j3SK72GMLDZfo08Lkl6UReOFiglMVofRAnb
upKSdiJ0Yawla4gtuJjs8xJTP2waF18jtDMtSivtPQ4qmeRd+HsOWIv4NbwXN0Ij
1VqIDmcj6TdJ/GKP0XW6hV72IBi+dV1UsPw3TNl0CPAJ9533yDqzeJ7OVsU0KdpY
GlCIfhRC70g5MWtaEpuUOYG+tada49WnHrTzQSpo3hVg+vyADfA8H52iDcf2cMQn
gDxmXwla2YKZ5D99cA1H0upueoGapeuM9PRHJvRu94q1+Bd4+PZb7sqHHnJZi7Nn
OQdUgYgnPSqOlGMpBc5mucReCNVAPvbo1agO5jamIaXxxXYDEC++eK9qDIp0tSKs
NtLeI4j4gakhqSsNogKUzQNXNxjCCmpuQGglqySNHzej2hb2d8nCey2vpkV9+XLq
MDZrI7ppmud3IP7VIHiiqYO8ytpQGOKEC/QM4zp8uhnU7a4qk9zBb8/ZQNTR7Z/M
Dn08Nze0IHv86m3fSNT4ftHAp4DsKPE9ZJJHzQrWfk+EUxvHK4/5g0a3F1P8bG8D
sRPz2+bDycV9HBZJYo33yJrcbidTr6lj4ebHknlVZcBfz7PNjap3DVqPV3WNF4fs
DFtTTHYA5a6bEtAz+2hVjpUql9e/ii8YkS39ibXIV3z25HnwNrXgh71kl4dkeCiG
ZWRKfcZ3pzUy83KiUfK8ImuRmoyCpjPbwjsr3hWuga03fpBB4TGgESLdCTEquHKH
VYc/5Isuri0sqVqLFs26V0s/2w4772++lcWxoWw+1mCho9Xbi+FEp8wxAJ+7H9y8
6WqmcEBi8jaJ2bgsZX7xCnpUFxFpSZvFRdFyf0QBVBG0VjeN6mhybS2uwXv7tm0I
bgwLcPNJT5C5i1wQ5Ms1BkYW8hQ/5XyEPGquIYLxiSrD8pNV4xGUQimCWcDfbmXf
HUbgDaboe8+cfKIViSefYcSpqaBSljtSW4v16llQDNkbhjSbB0BED4UfgFqmYvRr
bDDJZOB/qdS+/i7ovYTH28pxBXeJnH8+PIeeeFq/mii9rsBPQo4Pqs32/aoKt8fR
BEN5MyF8vYrDjEWjJSVFHW0IgiW1gDfRuCsFcr4PPKIyNV+FmPqNxwo+Dfuq88ja
6S9HfGEgO8PjPntm5sTBCIErhvj5pwVWeKEWqv5tRgfKAJ3fSHgDhdQzo+O2j1ms
Jg6nLveQsDw8z1sNaTOC3RWTim2LhxEfTCPwjLVogjCMNCWRqDDtLw33oesIeIkp
Q222tkf/BVTMox+KYJlV9IW/gZpkIij4imQkY8MWyYJgzkNshxmlTcU+tsouigTJ
fY2A3KDX7xpfK1BXrCdrT1dOjA04rUP/UbPoI3gBay2jz7L49ULBqiyer5X8YfyS
qAbdULUgRKniEhwFuHUnYmqsFUXBEiRYclFbBbvhCi7J7Am5UpyGHm6ZgPfRXXjr
KiW3zxfODFneaapoj0qHYNw3sjNYwZLTtgPXFnDgpxIHB7PVdxMn8j6Zrj2lJjWr
GaJRzd4YvPOip+dwKXD+bdk0yaXV5HYxXr92/+/sNjgoOm0RZxa/w8s7EcB5PEM7
Jxjgx/MPylz/++3AkCIlBZJVpcpORSprSD6GuP+sxXueUAiYwRZ8UwRN71kGUCee
IHgD+wiRkmDTuNShvwwlXdRz/GE/Q60NxNjCGu/Y5xUntAo4qI1WAXI4InBPiZGx
79eqRTevMIRo6TGHZnbSI+sujahudM6uD3wjUONUO1AVeswAWWDcADITVRUx0WNs
IV+kHZv1oY0kv0eNJk5CsFl2zWlvP70SZ2M+UxTA6jN1Branv79W/n6RGqwRVen0
7S4KxLuCaA2v7Le7pI6hdsXXgi3sypThMbOr7uGfFBsLQdnzJYYU0aT7U6DCIjgi
aScnLxa5J1dj+VfL0+jGxDVAzGP1bDQCqamBl8z1riLMHAzmIXvLl8M8UNGN8Fg1
lY6y6BMJyqho+bVkfNdGvVu7BZ4pz20cwQMUhzo6MqKZdtRMLX8kqQRuT9zLCiS8
+IwkLr491iSlfeOAEame9yAT982Uvn1+VboiZUPiyfEAZ5ZsLGiB5Y6QgkV/s1ft
QCb6U6JsuYCoo4muGfB5pCAXcTkpXw+/Xp8RuBqD1dL19ncS3HqJA4evVPxvS0lC
sJJgs2sPYdiD96fAbQ0z3yuxUW1Vnj1nbyQrU2qmdDHYHqc0zHp9zQNRMu8/7/Jo
FEvIJJA+l368S2zwa2IEENzF/430ml+24qWHecWHfhMxvhFSI77QnIx0Jf2YdPDC
f5+aQbFAKebz8L2tdQZ6Rx1UQlvfmNuEJ0ERNH4xJ+bU7Sinn4l/3p1HRXvVhHwN
7O2lEE66V0lO4nKB/1+ORnHQfD93TFJpHD/pJsS339MNRgPHP8QCk4w4EbqbptH8
rfPm5/L5pxgc9SHBjoGLMR5hhSAPjAkfrcrzTmI3CXQOX5md9JpHBqELUWgF8gHo
62wa0dE2QxeSj5oPC+zfB8XaAWJgvKr9oGEcJ5p7kZAnA3N4X+50NQSB2f9Q9kOG
2MyMZjEYLuDcFT3JOPPn5Upm+2SfU1ndtERW8uTiurEWYEC9vPL40Qj47ijo84+J
Pck4nX267d7Q2r56WX1UAO0qzvDNCgqlQwpNXUvongm04NuELlyaTDNtFgByM0Ma
7tnd0zn9mbe8Hy627x8GfSgGo2O9n6HzbMIsFX92OhrbqaFpPb2BZnU1QpHmX8AL
1XOFbQf6Y9K66+hqZpbn7uk2qBkUU+pUudRJsyQbxrS4FNcKQmMsuf/uRq5XS4Tp
G3FQIqQdPRYm8O4dHYCvHkD8yevY9z/N0i58pkB0YnHyozp3yKJbFFldgSLA+4ep
I2e0o6cKTT4HtX5f+kEtwGR2B7gLZo4Ye2FvrMCM8bPVGfvz/7XPgw06kTYjdwcD
yvtTTaWyXkO2oeP4TLNc4BrSy5FiJHKSgyF88kQqGMUsZKrmykFSXoZeMvodUb5z
84mPD58yHYlsE0MhgNLcCRTdzWq/62/A61mrwNxIOgfSTUw9WXw+5K6cYz5mrbGA
GRu16if5jUGTIwO7fFSvuJqjugIRGR36Sjk4xV1rCvifEq9VHP/BCiZXwyd6P61N
2jvEL6PblqyjPD/2u5LjMsJdAiQLE1QM2tG5HhpD/S7Uerx/99XqSvvpp8SmY7UW
pXEEr+KTHiS0sW2YT/5hzhkHY852dDKaqHcXE5JUUwlC2zlzAIcmCq6Z7ApTDqmi
QPUg66FO+S942PHr6PJEjtmGKcvHRlyEpAnMNCQ/rQykP8yB9st9LN37esEb3XW9
Mz6Ak79/S3m+8GlyExkzk9621i5tSwOBFsuTGkoKs2Mj1Z5RyPHRK2YxbBh4W1vl
uYoa5uHo+aKgBnorG6+L7zaw1USMHHfLjQ6MH5Cd6kLj3IVVNR3xEpQvQOA+eNEt
JR4ht83o+r4I+d2e1+Gwoj9CDUpJVIMpvkVx7h/WaKaNxZ54ahsGBIIhwm9nnlxY
8PwqdayKtZGieXUyATzqls6hB9EyH0Gqm20ujRMfRx/UHhaLkVFUjUJ3u2NtnMGc
m3VDYTgN/c9phJ053p7EPRR5bGh+vJ8U02oYPdKxOQgEVvHYjX4wQk09ngsdmxoG
u43Kvf4PsEStM1MUfiODKbbDCRjTAv9DqnqYu27MSr4d2XJumEsiAQACdL2DC6Zp
AVPfMHwrmDfQxIPIrB3dI1rn0KfcDA1w6wmZdchK+buaiwRT7Q9Vx+5QdAofnU+N
8C8naQ+kx1telLSVvhwN/LgHrlJhT6uNXlmnANFxFv6NqiQseBx29G6zryDjbrlF
EBIke7F4RoyjaHo2+B+ZRhseAXzl/iRFmLpDfsigz6oBUTyUAFMWSz0kJ9uiU5Bh
P1jR0YSjKd00z9dVCes1HmloZXYdhD/pYx4Xy+TaGw4++XiHTiAmSDvxPmimwFJz
tIo4Kz8icJJCb0omE5+rNir9aqTts80iLVYmnQ6OwiONM7GMF9uXnmYckDIqopVT
KgKs37vUIdAvVQSxiz3Mxe7ln4hArZs6+khfbfpEJfUy1C8PshCbIw2Sxa+uBNog
cEseqb2UFn1Z85Ag7TMRGyYQZ7XSmYqR4f/6HMGGSi/ml/6TsCHzYQ4Mjyc/Ye5/
pIMa4aZFSJalHtV8gUKbyvPqnbASD2vSA2SRs37K/uUYG1Wn44t/r/glqThzhPU0
0JoGZL4HfVZ2YDP6iyc75sVy4I79hB4epgV01W52Dw6X+nfbzCLZSEKbWsM+F9Vo
k8cWQC2k7CN5+NVBFEteAaVIoHFe7AAoNX3C8vizjEDjH6UN3ncz8ieltYZYPeRe
AF7WttLBBXiJ5QTxPS0GhcWn9GVhNj/kkfRqs2rhTiSIZdUNrRq3uqX18Hc2mlDS
1pQq/I7higImPwY5kAPCxEcJVQbRvDxtHRcexjKBEKgOpaIDKL+CIg0uTnDH53Xz
K+hLzK+9fwzCzS31/Sc6t51fYHljaMSw3dxzbH2GzWOYcJkT4bgpdcGLvRq41WVe
+tUzOvZykm79AoGXVikDgnkjBs9NpvlhnKBXmsd2P7aVYFbUKUW7gNg6jDcJgCLj
SeLT1se5nwYE+ODA9gtFtOv+2PldbO4ml20cW9qJTzO4NMW8siz/hJzsLASwdsl9
f4wlaachjJNsgDVwXqJqokR8x3b/kVdViPZPJSUAnfhtD3Hx4bEhd8C8ZPpIAJ71
mwIR2RT7RzGqCEoyFXT6ELRpx30bnXU+50Vt42yV94PBRu8o5dcEXFa/lh2gSfWo
3hQJsbMJvfy5o2RR3gO+tn6hFRVl3um0yt4JfDgoJdhpN+mMEM+t9XWTtk7nrrno
IwSmkSxYJ+IsaY4saCjjy194jEMvug/gUNiIQVy7Q5YUbYMfKxFm3w3NJqBm8wLq
ez+M7+gNlWm4bfai1RdDDRjbpqVard0gbunPTam6Zoe3p6XCo9f5bfLJbZuM2o5h
rlFdIRBg0fY/xdVyipphQSijR/H6uEKN2Ka+mmKl28XyGceTu29QnmiKq9uYPAQr
fRjYCaATeS7zuCm5yxJLj8AJfn84qqws8+I9gB393cd6E7oeL6xiQ7+t+ZNDeMnW
LNp91CglABC18QI+8+jKV4w/BaLphkwTRCNATz8823ujgNGhD0Y4Ma+dRKJoPck5
E4Ci+dMqczosjWGG1AAwvbZWbg6JmeOypR53HlVM8bQULOZlRyXw1l4fAHS0X1Rt
gzOFDhOoPIlddiUhDFUZ+gzQkMKjLydPSlvvO8rthHDjfiWEFEtlCBe6C3B5R/Ht
j4taCUGYPXtXcpo5B3Vhn20p32JqLTwikAJ+2g4NpkvuBTT16npBeulCafVCUG8H
+Efk2gRghAHYgAmY4zOpSpR+Qt+jXybXBElLyT2/O5WIwSqKBzWHYB0spp8VTlR3
Oa/z9WHWvq2mbdTy7ASf6mVBNhjLYXSoL62zZxRvLXf4ggYqjxgU0yC/LiO9rBOh
57kEcRcBCKxtGKeZfue1rnvcTR3Xb30NwHIPwMWa4ow3F55K5ObxnBNYUe97bDPY
g2VQ7lSy7sOlBTQ1IRjcMk18XJQlpZP0F1lO9pWUIwMPeJyyuwu+4N4O572OOIVz
wC3NLZYq8fdUvSf465BBvoTcmIRDY6MCNUGn4sp+8mmKDwVG5gdJT5cEfNQK22u+
A0zT16NZO0PGwtPAa3i0ojwnVf+R1zE26lCPsdrgC13kQoB2Vxfbm5xAHrYrmUjf
RPtbnTxoSqhXecfv6PETUPDMufCP2Xj1Epys68lQatitnxILnPh5TvZBPkmY3WD9
na9he8MTVGtQHsWYfIML1qtOyRf9kVhnXF2VFZ+B2W4ASOlSv0Y2RQLa6l1EUCLT
5UzSP7hD/RideZrcSaOkmhAkC1MX6WnZvJrOY0a9ohztGdzPrt9mrMUvzSwWLABv
VyDE+RvtQjM+OxoLofzlxxuVTx0lPaFjMruOQ1aDsEt0zC3trOQMQ1o28R2kco2R
KjMrMRyZ7ajzek2O/J4tvvHh6vTd4LW4otMGnKtcaLc/k+fERDOSLaQcu8vmfUqL
TNPSMB+M8WPZoip/0u0YbXMLl0UragegE0p4Ow2B8gdzGfE4ljqqmPpEL6vzGP45
225qDI8fbZn1htXYKG9kn/VsSlfGqVX7Jjiii6VditAsyzUbU+vybkPRSUPibGOm
bEREDcwRUay4iT8IcAVN3YKTIHpoQSMbMopYuhIGqBXJF56u/BKnv6M/C2ZX+eT6
1Qv5EL62TZcYrCZPN1F/kaFHZhODf7wCZypHpON75ufz89dZGCw/wX+vkOs4Gt/u
vFuWe5ur+MA4EaE7yfM9JQxDaFXH6jeKbx3Sljufhon0kSz+0dOfyXo6+O2DQt89
LfITx/H1taqxh25RBYSFAh+yaamQL5VLnJUwa+M58sAEjrwgmIBWp8zIL/OQFYPG
3XNrfJ1Gu5Q5Pd5cK6vBsMC09NqTKRXTUzAMfGWNlRkKUKeS0wpUkn5ddoRjU1tU
vVTeXyCCK/A4sa1NkZsLSvyhvnqJd6dNaOz4XcbaWGWcjhV//t8ib2CJfyxW7zI8
OshMqeIitAl3dh/GgUHGnme/DvntBa+tLYZEDonghyJT6YVNTkjn7uzFr1t2PMYY
i+/tW+gXkI5IanwekoJMlqgOiPuWPoh6mwmPH44NoT+oiE6w3a7v9w7TqrI9UNVD
hJijdVmTyoojz00BZ88206Y1J0JPjV+dgfJPaWeKb56Sv2AgBg2vlASGq2ZjS9Lf
PB3gCiN8FUYMYeO5J2gXZIJfVlZgYfG+RkeghkVh1pSGbvvenAkkbJitm12/ibw6
ogLnYHyM7tw8XoGxRxdQwqtzI+E4yYfSyDx+E0WSU2uz2jwK2sDT1pV4kcy/pNrm
W2oLPBsHK4fuem7mCPYNHr9SUgGIDQhqXg8IqQ7SlV1mbrofysxTHxYkxQBlJXrJ
vaMJPpZg/UWD9ZR5TumvKQenXSlt2+ECS1O2amy6+evkj7zclAStsjIr7+Plx7Om
fu2Qz+mfCWm/Z0GGySaA4PyPKg19mPt88Md/Twn8TAsA9PH1LXxXY/Z4Us5EKphI
eA3NCxI2cTlAA7bTxX3y9x6ciWL/f26UQuBA18OFwSSPehFysmjRvp1gH9DzKn+B
UaDeQjYqyBylaWbyZaFExUGe/ikwZSbZCcdL945IGtPYuvdqqq4Co+Hi4WylyqDl
RxB+aiWTsdih4FvRdTfT1BCm5hwOYuYLVpvA+zkTME+6q62g3cXyYKMCGXgsCCMB
+7ZtYZbZYPGAO2rCXAlrGHT9VBEcMQvujNIHiFFvDxL/chHXIHWNtGS3N16In/lO
bzhj7kIBKn8i8iy/F76kO3hgvOyhA9YLyxjmMFBOlv63QqLfV14F3M4BTYyZbXn5
suoJ96MUQSi0eIOTz0GVB4iVhMD73+0F8hnYXTspBRbMT5gscg3uP5ZRBXu8ag8P
M6lSxBaPBUb3vb0+np9CMzndjuBIwVZlpWGKJIUVYQsZReUAXjaS71t+GRIH/dFG
ltZBAiIMfIoaNIsVIUA+8skUX26Rg1tS7xqWK4xdlVTuo4HcGhfsgHq5fb0pb2UK
2ycnZMT3zrX2y20gaqFX5vqWRyUrEbOBzP9JRvg3HvVYEOLoYPx3TmCUOIcMaGNn
yqBGW8qtCiwdRoksoLrJ2WbvS4n9RoDMLtGFJIftp9rlKpFqBUjnkZvNfdWNybvk
xTt0J66rqs9U2xiurNDE0i+84THUWc41GFWKY52lRP6TadYarMo65g7E3YjCfdKv
4UeemOkk6VYSQeMti58GbBZB3/Zn0kJhP+m91Ujyk5b297ENh0hkGakzL8OWzdRh
cFdgf0rN518CZcfIzmp8ZlFCkIjq9hlHLCyT9f1SsH7+e6Kd0UUGoIGmpI3xoTsj
tKJVa+1LV5CWYazhpPSzxhH30wiGH4G6MHD+pRCU4NZhzqqXyP9xIw8bboTuj00Y
iZAkdsEEI7RpI0DLx2lCvRJ3/pLHGyoID//BGYM9H1dh6+nwFBWC99a0b26DIX+O
bLo5JvEjzmlk99xnE/utabURrdcgNFyJ3VpHpNj1Rwe+XjVjgIzS3QXW8d0McME7
LGGcQi+QAQg0aXlHLX0V5JZJ0RoJJakQ/vJodUmJnmNyPaNzhtGUxxTOSKgQ/kXu
nRvAVN1oG15onj1nFsxGm8zFkswas+I0vlPfm30xnME07X3NMaLEUpmqxa3qsMEv
neVG7xhiD5zC7vcqcxkEMY/0F3ssVx0DOhoFjIP+ogXFHG0tSLDZHO4f9AHczxji
N52kvV6lWEx7/i+qfhrvC9zzlWoMX/tqOVk2plntfhqeSMqCU64RkYQtYKPlTtv8
fKtSYtbAGqbAUSuG51jf5whkxmw2w+LK3lKTGLMilNALMTq2cBfhnvgq+53uzjME
hICZW1jEWKdH6c2IMPWRtXIL965ZaxeKZjFYMp514wHRNScYH9T5GbxwbD9kCwqZ
/O0cabBsLnEAielHKLdevLS+In1XQ9QbKhLC7MU8pL5R+8khy7aXc8hkxPrFyF4J
oKFvMZR0ZNoYp39zCrB88rpMh4hpr7MwsBw3O9kK7NAqZSqUhuNwFaoi/Vs/CkIS
SpIrqFISzCrVHeESJTzwMthQq8fCGCybqDSU8WZ+RnfzsxVQlzZjTu9c/OT49T9R
dlOnRdKp8GDUYVYCNMtME1dzT7C5RE4Jd3+Ao4g0rAx/s2+FUY592wRz7/QgxKX2
WYZnfnZmSwvakYunFGJz/fIoPE2LECz/ahnO6TamBc1m5mNiTk8agDPLiCVraSQk
LQ+S+Eqs3uGHuVUQ5YDBFgqVV/3pA7JuiHcqoIPBDF/WVyFusaG9MKKdt6dbZxdr
PNdWHKcpHSGGgy25eUDsrIEaK4wYl9CvMUChUkBQi8YZqql7+mQEaNQCGs7YZ2oO
oLGs0QEnzbn5QQS6QMMzmn/JLLhMWAXcb90g2IVBZeSa1f7iPPgrNtoQ/IxhlFuR
b4eGJWdHPcHDXQ+4JJ5+gXClgMXnPg+IYM6a5EaF4CfpgtG8JA/d6JfyThpnAxRh
gHY6+SOp/bXDKrlOPdiwC1L6RkjL1avqNKuA/E/oy8/c6c81sE6u/Mnh4vQVmOAX
RUNFaf6FXOSmG5f/VhzwqkeunlSV8e6rMWAzK4EKNX0yFJo+IAOIxpqQmh9mhKZs
`protect end_protected