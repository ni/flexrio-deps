`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6272 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhEl66vkmqNIpUVBO9a3D9et2jagLaXHgpCw8XU+WudeV
UMm2lBGTBxc515BEC0lQCVpnkonfNFmyiTO6WTIU+l3CRuYQYiWu5eHFc9yOAEyf
oAZVUToxuPleCTG0sdCo8c8WANyNS7rwlG6cRVexcxCw2li3yEXFnm6XM2DwLWig
CIvGKsHo5JA8vsWXJN80KaLs6JbddY0a4StevHHuP8m9dxSwPDrA95FAlAkrJ2nR
AWnoIDI+/jcLz1oJRFMFSoAZLEb5lpPC9zLBLZwP3xH/c18Zf2QzskhFm9dFEoSt
v7gKtKXaAKkp+N2qmviKo6Wuc7ezZjXCCS8hLzyP+rug3toLlh3naM3awLENhBf+
JwifmceHM4p4CMj8tPEB+/CXmFsKXfTsr0nQt4MsNcNQU3+1y9k7XlO8072z7qcA
xwgifmuscMhWg5XCJKQy2H64b+4Pbjbi9GzSCLCNtIYAZ43ikqmb0jC/bU6XpaYg
W/TyYQaNs1aPWI2uz8juuAZglUyyy+/A+o+zboLxnXcYdGdJeTUmSIbuwQq5AxSK
7Ww7DivAdHe7Q/bS5Rwe8NhMMw4/uHWEuJr6gx55fxEtXmduPkDoTLEry3RV3Qn4
E4OnJsb9TmYlbD1DPmv2AWOlReKKEWGvZYUNn6l4WK3ipTndLI/sWdoE+iAyuZbl
6lI61QW3glsOMyoYXfRvJ+n/nS/N4NblmmUHY3GmEoMK8pcUtIA8IDrUHVzzoNjB
7B2TSm1csG6qyv+rdth+qgV2QMbzWtL5dWfkdxPOmOrzFgLuAcWSYAQKmjUbL6dt
fq1gouR6QhUb9jm9NCyofJvLoW4/3Bo2T0GMmMRs5f0AAWmub8GBEtwWv5wYPjn3
/VkUEQ0UkoV2IzdGsZEYFOiHkHys2lFtRFGSZtC41j+JW6IlkfRXM5lh067opuqF
HUloeGYD9NdWNgXAfa3f8H1JU+KRZQoz9GSgmV9VWL7g1Kv4dBgDIq8PzdLeXkPi
OMF9ttiE0onWYhDQP9UQx4S2VcFmjB3Z0lbQ5dALQ2XRx/nQ+Jv1aFIwqhLEsunL
ZPcxO0/2xtqm0k6rs6VhgzFnmSHIPGZVANuNsgULN6AQLtB9Gwz3TiXgLc/GGtGf
GXb+FL4vjLB4ASWT8PxwF0u2p7ldSYDy5b2bUtDb/XDMsd2xfJV7yvKSkePeYu8D
y+CGBlcENmpIOxz3Whoy62Sm/D8j2FMd9PNyET/MsvKeceO8vXsTaSGPw5M5IvlB
gFSzS5yq45GLff2gljFGdm1XNIjk4xaKAdeClHsq7EJ42+rHK/qgAGqMCmbaP7MH
rWZf3Eq8i4kG5wGvr3m+XfEiX8MuQ+WNh0LnxzWBLo/Xg0HE6EJp1+vPGXLdrZ30
427UhirT7hfYnsKMBG3FTkQ9G1rzxxXSSWy3NHL/cqySiURxnPk6qKudjY8OYKie
NN9CApuOTxndYNHe8uDvoEGHo41t8VMmGLBYn8Hs2aAuxPWrBW6+K9gVwaoLF5kb
clUKBdvrN9ejkjdI1fLnOg8KYjNEAMPkUCiXSR9qCzmRRbvRVP5l1XZWhsjOcb6b
UQHQldA4r/HVEQf1gZfTlb4YytAyO4LBh7djVnpwTYy8hgwBYDiHkeOlWd2n7lhE
DIjM7s/5g2n9kyBejYuEMPi9uncm6vespej8sk55aPgcdsxS9ooej0/dPzymc+J7
IV/LO4vTXisCM4PsVrbWCyXgfyH0GbSNcWJNGwjUM8iGo2vS6aagqSApWruqAZna
FxEky9uZhLH05ToLQVqOl3GVkF+9/nD0vKMh2itVmVvUJBGp4mrfSbSh+xatKxgm
JPpE1Qek06+mNnHgAECoqfxdQbMVCXGGOEhpSo5hs5BfW2CvBEZQZHj/mjXhO1UU
CEj4wNNMtDC2dAj+GS6p+4QWa8o9lyN654DcSMlqCDkuDK8M5lcZbCKxjqnsyFdh
O/Gvj2XJrZIWU4stHPLXasgC8C4pHkeuPA4AnP9PpmXPBgsMPpIF8kGH4AA2ybyg
eNS+LHMTfr5ddZSWlkiFcpNoynDUFdw4tWMZflNLSgXouB3sf74aZQXDnrpjD8Yr
bpPDcYY9NS404rCPhBnpgWNvp8aObKVJ700GWkXfMaTdMybzIdNqeI5eALhe/+sE
7lP+Welfxw4tomwU4ymcPc6UKiq1jPBsh8/bePBfhoIZzunKGBoAOJf5ZmMXCi21
2SJQYNEag9o06LQhfKC8B/LfAYr5pY4g5u9KEJoR9jqRkQmPp8KeBi+uQjp6QxKy
3Iwhd7LcS3RLsH5xX+KsPpKLcgC6O9JWx4a1PP9oIe6yi5C5vYkgRnmDB0BZdlxn
BgWjRA76umhfeN6Gj0GGOfqH1LPHCdQ4oPOvmgku7A41IEmADezoGbPr2v+Bz93z
aPCX2xQZ/jrohccR9qkz006Ffl0XPv7BOv00MmqUC7NfOpR+5s7CoQM8w3bNKekt
qQ172ksfb+GcEpjW16wdRIpvsQ1DHbMCGNLIYwakwL97mceYoXNPTxODn93VBC+w
+UbNmi5+LX05q5HdUARRBWin+zc9HTUkCU/G+QaqO6hUQXm+9Yhh1LoPGez7RgHt
Z5VdG1nljT9+dbLiYy2UcixkkHBxQyHSySbDU78c85Nb+dDa4s1z4IthLKZLfEnz
qd4hZs3p/zKT0rL6BQpqOL4NCHUbQ+MZLabIghpU2gtLz6KOxqR1/4XhRtezBwL+
Cdldu2Ld8TxZX3JpW+Xu4v+nhyn6v8t1aoW3LET15XhrCJ0imRIiJFCcpOuw2RUG
IWybsK0umW9NgYScIS9RJeHlGxe9xcoJUsikmESz4gJIMW6Uca05wQS16IBEmGpH
benVAh6zALIXh2M9BtjYohdGipv76bdvFRKFS9LvoKjMCnURpK+cBzovRM+vNQWf
RGcLjj/yEUqQSZz1tbE8B0WXtxmM0XBcNWSGFtjszBVCstpRw5qTzBIsX25j6mqK
h+8ZavEyKfBupPImQgIPs1bp1n0UCkZk4nkDxkzEI+RHH5aLxmT3JJdS2vw14/CO
b8th11lzKhpRZ4h925CW06kgTtxsJ30hfXZPGgmlG3g7balWyJp++Ht98XBMpAdg
xcthrbkEnqZfXGGUHbkTsVUMVKy+v9qXtPTdfd9ow4HXsi14D5jNi3+2XgYIR4FH
znBQxpRC6bD5c/9q4UAmB+Bjcm/u43/djDK9S85yqfWIRKogwCJk25lhHSe0ra3l
MJwTl8L+WUfu1OnvXSX+qPtg1hYKoeWCaueAMWxNRo1s9Ny9jKxCQH0o06Ft9x7l
dJWV/U69pfKBAPGD80sIELzmcaEPQMn2KFq6SjUT3s/DvPp/0a8TAX6gLwMuaefn
f8lmT4aKIYGRSOIcoscqtgrV8vQyPPF3a+slIJXzaeUb4teQ+XevF8ZfvFptiloU
5F9YgIy1+Xg0fzQ3jFekgIv+FrLfwP8IAvrELMxTBaRt5XlJGiZpjiQR7CEcMkdR
MGd6HUGwPvturkrjGANXOUsbJ1e0x0jyAxfhN3i/NkjUIvSrBQnIcxbF7qd1j28G
RJ8xsbZpVVeBmFKv5TI5QwY706HhK+41suv7gIdIkCfedECuq0xMu+U440NEGX57
dXAbmslv2EBUpbV37WWq61S83JPp6wJPvcbXTKCaOAcyyZ9TFc3KqLGqyT9NueK2
OFdtJb9Uw48lreFP7J21XhR24vT7Rva9zXItDxr2sHKXUtpqOQtGTxNC6y8VaPUx
m8qQ/uFgGKZ2bZOH9BQEasIzG7HLpjh/MNUcug722QkjAKQL5EbRUi1z4JAJPHok
xFgG5bNyl1uiSEa1Up3xGOe9yG6Zg8ZymyfFYK6CcvB2wtUDhyf/0JcGZ8pamXxK
5ZqbcRVoKCnctCRyXCe3AY4rnZSs2SRPDSk0jnMU5ldt4DV05P3aUWAWvG2RWUAT
RwpAKqA6NLe4ATlaRDA3NO4bIhW/VIbe6EGURdL1mpaHn78FiUSy2bgLzj3qMil6
AhP1y8K9PU61vWqwRgpILto1rAUqMVFw7gDBY+TiS2u7WFBAVoBDP7ursdiSFyen
53YJQQjP/bSzihO7FVXcSAY1Tyu+s2q7yBhySsbQRVY/Su4ovf0Eod4Y7Cn5yynT
ARVFY3B6DViZ0TSHJ0i3kunycHpM9tt7uT7ButvZsP6HhtgNvGiAG7U5gO843rry
SJBaNx2wCBRugaI/DgAa5E0HtfKNDR3jLEehH1E4/3T7wKi2E7gTByH/wR2QbiwZ
RKOvmF/a09ezT0HOM7ia0UWLfv47OSN6EG/lQHl4Y+0y0VrH4CrPvBdAlHN8wuhC
P5TlqtMQe4wYy4a4hoECSjgpOSQaIP/vBCOCA0WLU2Jkh4M+UVcSqbqI5LuxTeCW
G5zhh9OoZa04SuhgF0RBPQQ10XdU5lk9QhuQHEpxkfi2pxYy7pcPR60nkZegfEZc
El+GQfkF6rq1AdTe882xfx0KFeszYoWIrJVCgc/hWz1IdoN2sFz4QS+TssffcLzE
OYzQv7DC3vxE5FWMK6qUjbvi17oM7KclG8aPd4gYbAAy5d1GuPYHgz6qEKnia7k+
I2UjOjZBPB68CstStAGDWX/uwbLUuXmhPMC9CuQfnm3ejW3NJ6omIVyTO8Hhl7IL
lFoKt0ja7HlwxeOC2RyAMatuu1hdl5xwNYoiX5unvW9ae8SlSpGstLShrOLz60jV
EEPu+nwB7JTaxaHIusYhDLl94tn3B1W4aNhCUf9LHb1HIPldlnGgXAtwJLHIxVIJ
4mV/AcYWkUY41jOjdBKfmXXcbPHNV43I/krkhiAkHkbwqAg257u/0B92QTO/qtZ/
Y4FD2fez6U7TdwPC5ThupywhLvnTSLZ5X0YnVdu/9akXepuNObAL31oyucFj3SlK
P20MfyP/GiMJdhZzpotG22D9Imsd5qzUNxnnX1jUIwHiIVWBRzomU1E69irJlWNM
rZyrRXzvGYQoc89hztdk45Sob4XezDkADoE1IKX30l0F3PiI06YDr1OpltenAdIH
JEaJVxidGdyyfKfujhH6zD7jS8jlr92mIDRLYhWRUApKW/OEpygsUalEQe2H3mEV
GCISZ8upsVhnuVO1oe/hKCS7ESPEwvK5Wo/jML1I5Yt8b/cvvrnAvz0cRY17tttG
Zm+sk7wlnkTViiRsA267OrW1oGHbXKnl4rFFxqqIK5450kOGP1jenHZLpQV+bwms
k4xjBfuovcIOrC9v+/1bnDEBKgz9HbbTmHKqZtOG/vr10q3tedmuPH7OqlOTgjKT
n1kzy6xJwtCU/0IuAZhg6FF5CS53t0J5cjxNGf/EULk6DqVCAhKNcbCFLPOUNVnE
d8SqZ4BFZsLHQYYmtgxqpZqYc/WlGPRtsljwEZmal0dvH/Mdbw0WEtnWIuKdbjmJ
9Wes9rGFh1A/hWGJxe1YUiZI+Vi9IUFqW7qRWcV6L6BjkGJaNWchmRtk7tOIJCei
O+SM3tNYH9MxGVYe07LRka5Fs2QBMC9jTmwuJ2NQdsI/hu8w4WF/1qQmeFhmlWtb
W/0CyDGSVPSbB2a5j57lV5eQ3OabO33Bhxu7++yBqqRgUeV9Lq7qO+NTCpaqJUQq
K55Pze4l9l6bELmBc3KFf4TMjUo0zY2bTDfAAHiO/6qFhkOCARP9Q4cmclVUR26f
FbG0WkBHx38yJP2bJ2TsG2NT52y9OWEwhJ8qufn3gFNr7mrdr165tRMgZdliQbT7
PRs6LLGRJxeveHqHIq8cimYWEMaDIrMCEvLaQwpLsUDOtmRWwfz4QCeANo7r0f3S
+522aPEWqDwPbGjAFBBS/kppjqBZ6uI89EcueLPF/VBJ5ttR+yCcj05cc1p/NBfS
B4P3z4GYsHQi0xKGmZ02Fzrp1g/VBArhKsc5Ax/WOWaBAG7h79hvuvddQxcGO24e
AeGShO4PbwvvQ2v1LCtkilYx7YgGhw9+f4jlEfaj7trHBM6hC8ZYGtTJw6k8OQWF
CjfAQyMldzEXutHDUPFpw9cVa9GgvZVXI2sR/ovoTcTVeJgozRXe7qWm+xizzrVO
LVk1nU9ysPjM85wWya2WnbUqf4AxSUF8myIFX1qZw+Df2XHr1ge9zL00UbA9SKkB
xsTz6rRSvN+fuVvcFjpTDfIJS06rc9H16bsfkRsdUfTryUyF7vcmn5IYJOoIVuCm
Fq67s+LKs0QO0L4BJiY8WbKa1QgeAzvyr4NWskufS+h33dt/23uGYjxA1mL6/Ze+
JsRYGtLLASMVJjXaaNqDLmML6+pwja/dxVKsS9/MiZ+l0Ja+y785i/9iD+ZqTYAm
y/bCPady7+Ysfp7tWgAzE3t5YfKMXR+91g8J4vPMdCMYKRUNItIHKpj+MeqSoiPG
yimG42nea9Uge7eyS8pyOM5QIfSdohwTwmjjIanwHQ4Up5TlYj3Ktcg7c6uMPeSe
xSpadcstCDAZQq08jWQJ1mjTIspLQ7ilZJWIijmkfLEex49OLmszUHtdnWcQSXxe
sS+j7bsuzrk6JI3KuvdkWcGJb2hcIOmV8+O1x35hM188tRIo63Pn5SFf4fG/rRq4
0+nEPvxt4W4CcvSMdC1SxF6XH+n6lZRL4AKOfgZgQwxMVWrInZ5W0yCJZXUgA3zR
vhS2nhWYmBzAZBiUIQmS+5aPinrwi9uyiOgWoQxIbuLYLxCSV7hvJYHMNHitkKe3
QFZ+EMTTBCkFfLuHRHfrMP/RloTaSBVLBmG1AirD10oZFANlVdvisgliCozLqp25
yRwqK7LvR/etX89nLxFxsdnpdnRBEP9ZG9dqSgvJr6gC/+lwnxJOLWqmZ4XngfUY
uqpbQ8etZP1LcncZFkwpPPQ7a3W/wbEGsPr+cVJ0jfxi8IWwQ1PXwRYMy3pUJshe
L7IoKJDSTdRYbJg4aqJ0/4vPULPFVV1ReJwncs15j1h5bKXNVg/XkCwzO8CyQCs4
/tqI2HbTnM5TUM3UgI6w93c848h9WdqPBZkZpLo9Csp4O/pHobGk31c4/NOitA+P
zkurnhE6nFPFlGf83JSQSILWZN4myEzRAzGJ79/lF+Bg3kw1zHpJ8GTJlOnRVPv0
+3wa2Ez1t5uRC6SFBsFsoPGxgnq6WoIIWlHimpWANLj8x1rEv/8HtmaflTLdYJpo
O1PS90JCpw5zFOtVOAICk7y4lkEWzkXKoWAkvAXVVfr0yDnaiiWlKCuN6wpHOpxl
DIDXYkIF8rca6jKETJjXyNAx2K3ZN6IAoa5iniodiPBszmp29hqL+Ri3DfL0Lco/
vZopW1aL4BAPLvP2+CbJtgNYqCN/j+l6g4SeYPUkIszwkvR1fYIIf56LNo7NDWmK
+qqDCZT/6IEFe3t/DzEC4Um4KK7/Lqs+f4Ro3jbY/+62DzB+1jp2wlHRuZsXaG8A
ZW9FRqJvfbOqFXUPhgQEocXTsrlDXoPX9ToM5rp1WxWnYOZOnffzUvUs8KMQcTAs
umqWp+MhGOKy3z4W62t73fv0xWC4+bsM0+PXGIXmovxW1NgOQWD3LMsH8d2BTZxu
IkmUcTdXiObA8uTmk+IGnPY6Em1BFbTRImBWvuei7BtD5UEAjk7w5gGzMB+rjzLb
lsZnl7J0A3SQn7C9kKmw7wtkeouJ/3nPKixLu0oPcs+T4eq5nPVT/dpi6lGg9bQJ
0Y6SxQK0MbQsHyvx7h0Effj1j2BJitTkO4KdZEU/9lTly1p3fSI+DxMbKHpV7uGQ
FWMXJvsnGuIZ8FfY5cwEjeZbLBZHoz4yTziBamN4YdRfPCb9RmGfFJrV2CU629hr
IOYl/f/qXAFfSrKgZpcABNTwTX7hik9hIx2Im0mpziRsdc1kQUOOU33yOWxlOmTW
g9H6+riMSoZr9JYz0U7UxubIHr/mOQ15WyR6z2jIBuwnPE6EJCP+BsNc9AKzuyxK
uIEVc3X8Kcn3ay2U5quQRi0Bk8gCp+asHM+ApmCM68LqDHf34UWPQsJTdOS0qA7v
74kkdr7WrP1Hl8eWsTv8gOYDu7l6f8uZoT/QD0ifmjp4fYrKL2AXHMs3gQyPh9yV
9s4vDa3G5mZ0l8b8bpU6EumR0nXEArIZJ73SSH7L3wO4ongJIGlxsDVjwFpw7lqS
+zzGN4EyBh0vXjb60NQ9x5F5Jd+yi8PKD0u1tWtimoILhhpUETbJRvE62PdU50JU
aVd0nk1j6blDkJgWQFfv6P+y7cxZaAYd3rGgq0DXgb0=
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6272 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/T97rZhQva68T7JOm4bkq25
b4BW57ADAHEm2yg/Vzsfl3PNZ0qsJqYKXh6pVrKzRkdzWqjRoM/bKgPR649DfQ2k
Kfv5LtqyjFISBSHkxN4Zz6eU2NUjQ0WIVTXcystkTjXUVIPcZS/7LO2PDt95iaoa
NiB6TCi6hUARZ/UZVegZ49GH9mm/EaqvFxa3+bGomgCAXhgpnbi/za3yd3DiAlz8
xSfvjT0kcblcmamHJYrPAn6MrTfcziZHqepmFqn/K2l0QgzGMqS2OpmLgZ+qOkOy
VOjUvNuSQk4teXVIeStWGfhd3bUzXK/zFHZ/fzZkBEVPq8qzHeiAdF54iv9CP1Zl
OlaL0sloZsrJiowBAcxxTLiR08yHDTOyOE0nQ2S0Bdji6APHTd1u8jEYhr8f5ze2
OdHwDKcGCjNlsUR6nyyDVFuUpGEHg0EnLrRETtssXEaDedLzEGoXST2Y/sN+ubex
NKlm+oAzmYncMs82HtvgQqfsSErMCsnwcNRxi8f8rMzeyn+CqtfOuxDsWVm3GBHD
AbndurTIS2hNX9mao5nL2NLMc1+8VzDScfcbPoDpEncsiGTKU3zVaXzVoxT9SIlA
DpXRrktOCqjttWLNzbk6AToFbG3iJCTNe6OzuATT56t3O8ifL5e5ixfGuGxxFY8+
T23l9Qgmw+WNUj6YnRn8wUfpFRWoNKqlMm4TE6jng4JcJuS/cllCDQ9MiI16mtwX
kGl2oI/XCapXxfpYA0TacnoZT9UtIBPFRtgzECugh/fJg4N7oIX9IstCKr6u+enY
DGMRgJDM85KAH27UqFL6BQ9PWrtH5sE+LKhWoKTl/tTLpOhFpq7yYI1umJ6Pmyz8
BkT/Cb9zIaJ9F5GJYkKqSIoIxgrosqtuhmubfRLH9LDqCDUqz3TkUAMcZpINGrKW
rTR1/ZsdeyQLc2QJZFhDf87AZ4HvWxVIbyAH6tgG1gruXQqg2FQEhgmAy4gfVS0b
R+xGjJNdM/qDL08W1vZllPGg3TGIVphogY8PHnuX006Q/kf8zd1JrMEVdrNbCHRg
/GTcVM6eX3fmuDRv3vaMGD9IPwd87lxx4ZBFDZRtFpzTvg55zC9TNiVP+BKiLgeb
sKJF/Sd8+4tc5b+i2wvHM/feB9biYI46lIOkF8aIkVanlvqUXZgOiCNidSPqFdkU
KmvCGOBKv9QHpbEkRJ86WBEDf4MQwypo7jT4wfTGMTFFq7sn7i9G9NouHKYJHG6o
77Bc74mHp/v/XpNvWvyPmDsyh1zyr/RVxrRKsQu/2m+x6gWB/l31OzRYuJ73x6qF
mDwuVyI0JJDI30YfOG+u6fAQ/y0GHLVsiGNRqzqNRZ0QnKYEIp+wKSDfw4UBHJHO
gctgpmLP4Jq+hAQNVa6g8iGtTQOjJ9/+hPDMKTUJx0D3NnZMMEFHZl3WZNJizvcY
2wCkXqZpSuO9dIaX1ZUjjNqdheIFKSlqxKngrcl0C61uoi+VKEzyj2pzGrxXYibY
W/5s6+T2QQX8ldmjHA3CN/Rbxl9UD8jAGE/nQAWfgb45nJ+sb/YTcV2/zOuGBb7T
OrXrG2nc2KhiIJlBAcABZ8b9cOa7FXSlBHDVxqDV0oOrVlazGIFmNzVA4oTiEhlW
OyNbhW3+3UaCB0sw5ehz4ulAH5c64d0mhcOUFvy25Bho4znB7/T1XkjUAB42CClW
fAYJ6nLaTWNZwTu8UARjCL3akJrOaymIPYSfNOAN/JigMTRrHDhVloj2oN1r3ycY
rWXp4yymio2SrildzZ/d3ZxCdqmcTOqO9fGUi9FxgkS5kneBnUrLbbnawNnIpA64
74AXFp7FqaVOQry26E6MhgXsZR+B8EzdOGWHuFa70Uq+XW1CjS2Bh9Ks3iZNJDY0
K6Yo3DRp2aMTk8TFav95Oe19MJ/UO1qTKdygQUMkvowU24ArP/n8xnCFuwcD8ylE
VJJolfF2VOKhdUaOZPmG4rHE2inwdHcN37g3hLDAVg+b7WWqVOXWflP3TmTtiAVo
CdolcOGG2G7+dCLyXE4JsIhGceHQ4MeuaV81esz/ifZ7q2gYAjwujpHgCWE44PWy
+lGMCFwoO4npuC7UDK6Ya6+EbBEALlu7dKtzy8mu4tOLayo02oEovPSps6A+DVzk
Vn7YvWpw30WfL2Bkl4UAWzaCNYoVWi9VD3OAb6HaDPkfTgNLxPhH+hC3+lfOchb+
XNuaaImL7Mn5sl/u/APMQmgLX9V70CXfV4+/sZ7qBUDPOmBbGMDKM4qpqiysRijT
rsto39MavpUdJcPSqUg8avCN4785IZXaKBesTuyYBNfml65TWhZdFjh5M0jz4nq+
48DgsHO+TmgS80Ox0cKU71k/vzgw3O6Zp3gzcYK0uZV8vyQw2MZUQD7dPmXFRjG/
qLie59JFF1Q4TcFgfu8nBgqY8r4UHMVK37+JjabzgyKKY6ypPIP0f0kASv2vFRdG
lEUetHOWNtY/byAFfVHgcu/8y3ppX3RP9+evo2OboMN8BPPNTThVfh2wsXvA57zH
J79NKiMsSiO9gKYuYmTMpd1lOm2Tfo1EplRi+YzyDofFP1fWLlmKxjP/vb/ehrcJ
hkSFzzPGla0b3ogOrTGv3UiYQfLpuZL2/eIYCc6FHwE0oPixQwawXhH3KDPDl+tu
TOpSd3jS0JwKrJa5lueaDmFpWWc+hOdAMWn4DNbJ14IiWfp3EBegdHWPaCtfuwmg
lMyvwAhV/LqubPneX7dSi7EBeLqWYtA4qdUdQJ0kwGMQPj5/W3P2E2y8Wo7BYV0t
6yMY7ecRLfir7egcnbzoCbXiCQWcvJIZSViN+J4j+jC0o1Vnd4WHyHhMQeXFXi7U
ILljj24rTKtsFRR5E1gVaZUGyYOv/+ab5BD6BAwdEXjnzQuEQGn4ZD6XZaRf0+Fu
gMHlguxscGkLv2IPYFaG/lxgA3dNG35aVHITDXiIFmsE30TfPbUijIjSvDXCn4OI
3GRvrNVIOellmP2A1+qj5Ti5sbp8k+nKz2dASBKYXRbb4y9FwMqBGJmVncBc83tX
7eIAZVZoM6LVzUpaSmEsoCNpXeEXSk11aBmbzaDYmSfbYPuBFdhA2U+EFQ0ibx8z
KsA7O/xt0MVLXK4srI+Bw+viED78DK/lK9GUg89uMYf2sitYx+ga+tDw3rgZXrGL
01TDnAX0Ssr21vdwxiaz/tQ3GliFtTmnV825Al+5fm5YVWzjGAiL4cf9tHnfXcgf
yTVZmLoPm37XFwkorV7L+3hFjhyKj17HO+NXTqnR396YZ5o7SMbx3qrfDTdBVo7j
Ix9w3p/btJxtZhEkJSZ3tJhq5202HUkoofzT2Rwj18A38DdrjcHxNtQPSCiklLVm
wi8svsJz5DNugVp/13HZSC9XuG3W2Z1EAhMcVd+3YJ2vEuO98ysoWdQOve3cXndo
w7Naq2mHkPVP0fH/tj9lmvxvxl8CiMGdnZP03ZnA2oZVaBPYTiiUXnHqCCJlmiXR
Xc6GtPj3kb03zrv9t9QA3e5/zpNofNhbT1mw3C6TMtlYHtdrbcH1WE86JhuSc75h
Bo6AnQTqF9nZLH1ijGTpa8MDXuJzsMiEWaxg70dxflcqatBKn4ZiZWjkAVsDdxjr
53vYXqO1vraa0BrYqQIttXtTi5iDlvkXcw7+SdGxFSDc2JBjHVAitVlYOggSdBMN
Wmek4JmT0ZN6A5xDlp1f7SgApr+TDsWxpDfs7UejRCB7nUP/ZHi7DGLoWFsURrnO
s9WRI+p9Lfr7UlGeQAzAPtjS1WTmZ/CRdMuLd1baMRm7SOsAM8zmvnL6/UkkIzmJ
Vp+gX69CPqjc1ED8lth4Fa0gV+iTW5pXRV8WmzsRZi7hEHhl4gs7ReicqoWLdIOl
J4pojprZxSgz8TNbuMcz6nOI/0ySH8esE12CV1RF8hp1eShCnakidzRjfEou9U17
1gDfTBTkXPuxNJ9lzvnOgDZfb6quipygj23W+ROm/QGSl9LpnhmY3VQGVv9Sxg3j
4Q7DrLZfQFIRRrKiZMoUwp95U/hnrsA3YKQ5utyE/F6CGv7cswFqBFRFiH9A4uy8
JN8SENpnz9rafMtXJ051FQXn/B5kp1A1HG92QPsd4dmG89IIKNLsdZ4n0pzbXHpL
q7ibtgk6IoUkIsZGhe3X8Cvc3oZPlcsgW8FWQvfe8pXXxZpKOU4NXNQR/GrnP33b
rOhvdljE1MY1SKA+S25W+MBDrCfgYggRUFmgJz/i7ghUs+MLZMVnCGVffW363n6/
FM3usBTdwiqIQhVYs8CVKJI09Nl8SObB5/AKetXSfylN3881KVi5HR8CIgmtD+BH
+XfzDV2W4EyReT4z+9DTOtBe7cX3C0TmQNxWc6MVCmQw6RZv+jlw//HpPNUAU8Q4
o7S505JvgQlnEakuAhPbJB8mHlqjDA+/bELERs3bCEjWC65UyccCPpEq/xlrTaJ6
qNS5/9gta/kkxOrUwkVBCJCDc6tq/oTVYsstrCl6wOrz6qUVGeuxLGxD0ZMHib18
ucuVgGW0m+bcPvFWc+hQRP584HHM4hz+Dfa5Cj+DXdIHUlO3FH4I7ULrZw/rBDBO
zlJQmvTaU05OTQJmvDkqbWKpHZu3bv48fLYVyRmPc4z4RIitoQgxov/RTK0dBx0w
yldB7XJcj1Qek12dT3m3/5KVBm7+UdYTPyVpAYHiza2s1g14z/Aac6tOoY1HAvvE
TcZzJ2P1pOj5C8ez9Ip2KwpaDerhs8iAQJkok+G8QY9pC/sGgnpTbJusjoZIldc/
Q1OwvdjssW1tXKlRq+qMMRQiIMEqH1YXBluJpZig6C5HMLptVqh8uranlaBlbOx5
MmJZJPJzgLu8XW/B7lMHoMg4wTdIdwb+6SzGKq+komN93iG9RBnc/TTW837BAmfk
Z1Cc8T62EECBcN9ToZubVJ3+sdyWT9jpRIYWtqJxmWvfxEjdk8uK/CkGZFKpSogp
gMWAJVdR+zekCAhTFYFWcEIgnZJF/WxuASwdECXXo5Vk146pHWRiRGszjdL9L87a
bLk5GE21sNKykSqHslz8GKE6Kr6bU+DBFXthC5iLGFbAstghd50hMpUGkXx0sc/Q
dd3GWOM28YK07zUp9XgRYwoTAdPVkcYxoCDqoNzy5qLjLmrCRYMP1m5CZlCbCSQm
nHptE1+ZIZSGffrm8ST+pCaWu6gu4nZuaCV3C4Mf2wo2DEpF6M05HWTFdiFZ7sbB
scbx51W2mk+Br33vVSQ+42au+ZaV3Cdy076cJDkhCpRn3rAMR48Brl7SX3ppIdcZ
KlaOKl5y5uZe/IjZbsurkGSSOpn3IGPfKQuYs6OeZDSLDzSLd8QS5TykcsEwzHLc
lYxGhhHC6ytB+oF5H4fY0AC0FPEc2Ux0w7S6PAMxwuG4jGwvGXnGAiiM6Clo0hVI
MLQxtfIoUwmAdTE0O6FGy5OTlt37WGy6Tpzen7KNDsmjjWw7Z5tJ/mOT4E2mCXDd
1TrGTmlGn4y+CKHIvmyQUshKz0Z6Um16fSc1HEeFuOKXZ/yI+S2nryyVd23F7AH5
RqfIs1bBN8YY8npR0dod50etRe5oESkRk6fUQMkJvKkCOR3B+fwuQgvi/OPpV5YS
xdSkxxx/YoSSaefZYEC/09UJWKVCPpeKEa4Ze9XmL2/NHYFETga0zBywVwCnvO3c
N73qW7AwGb6JmRwUDHPlpjSkwdG+Mr9K6qvDBHWWS7X95USUXQw15UBUwMU6XHaD
Qw2umt/C+YnhUml8ZOI/kVyUNqIdc0MpR2VAgFF6GNklFrPZPN2YTeHYiyuczJYf
j66AGHzHcEcq3pzR07s4yzj7iDMYISlWsWokFWdw433PeYoJW2WfbAh2XpQi3VLx
SdkKQf2Nm9qvlbH+c3auZG7tjG1Y1iNmwCdTBWd4JTPZVGGVbXF8KnZNTlF0X7I7
oCogTpGmOse71ma9Go41xOZf1xvtEs3k241mQXj+D18/USG+eOTFzblP3VFPPit7
c5ZKInjdJFn8et87vp5DbrV1h4LstBa1YgKtEyw1qvq4dcOQnJrYldqwchvLU8Bn
wqlqI1XjrArFHzHOzW2Z6+gWwBYQ4pN4T3S06BT8SiL6RpKqjzcUwYTyxyneffnX
QKgs5dEQ1aTnsVIIwXfEtWhAtOY8UdTXMwYSeEBiEIHP7FjEMvkkEXoqnaLIVHox
e9GnGHWdeWBRM3EBeABg8L2sat2CmkIzeBjslOJ+vPV7dK8Lx9eGp2r0ApvKWr7E
djhGqPMAysIAO64RAn08BrwqyosYphHH4TSQ6REzDP26kTt7bhZxdd81t2oZ3kEU
QlLuo1dDGc5mQYtucCdTF55NVD58ZqLpxIRoeEAF+Fc0v7/KzVY3bBvlxGl33Z/G
WiD1jYyIiCTWHzjUxKo2x555LsVCedqKes+bTX1JBjmZaE7oKnL1e7Kljdkb2sl7
wN01ihBT4iks3uQvgZQ1Y88NL9kruEuNosoSn+90bkWXNpw77nII2b5JRFt+IL1I
EF1WBgiXsy/cj5EmMvFQONh2CEm5NviBCc5/P51vKiMKiJYeQAxYWSw3tcilI63P
ueAFts2L/QJVVIdTsjV5GYk47ISM8KGUamOAOJOstaH1FezO4jzRyryhjgOnuzlK
yApGdtVXOhwY8Fi+k+NxwfkGTgJDhaNDydikx1PDaFz/DZKW18WqJ1tJqOL8pLJa
8OSoenUXgUnzqXMWUHMzauA6DzV31QQHhaPPE63WemRkSJMyq/JUb6sNQE7du7v8
ob56m2txYLhyug56JsSAX4iPvqzwhcbbbh2dOlRmqAY4EQhgvb5y4c6/7aF6j92J
lQ8kBwRTJAg2FjkS0hVvf1KBwhCbhE1j6FeWPuDOSw4luNvyb2C+X2/vWZvu9T0e
FusiiZ9tsdOfjBt2MAt1ks/gcyF7qnvQ2UuYeR66khmffdi5Gfhn8bqnPC97Yp/8
0xyEW/EqoIlJx8zi1ZQ3k/SjHNjoxncOFpvM91FbeMxelyeRK87O0mqMUJ3exi8L
iAMd649SgdWy/locx/KLMfUdf/VWSAQW8EID8IgqKuUISXsVxpzDGAXVT/n+7mtf
PNKhyQLzdl0vEvSDpKLZLxe6mZtf8si0bxtF+F1YmllKUpGPvE9KD4HZIChWhKo9
Ivy4okTRa+rlmy9GfUI9m6cZjnJCMJmg7SC2y0oJb/DHEUnKyu/XTCJMSP9pAufZ
IdFrNv2ScaXziFgLP8na9w3dihTh7DHURbopwUTrwwcvtFr6H18+FKH7ymNoesLn
dnFZxin0fdFJOIbYtqnMRTsszN/TFGgOmdwv88Ntni63ceh2I7xw2UXmzBCXXJR8
hO+eQhm+lkOiPt1E7jZlqk7JIQ/Hf/PzEqWcJNC156op/4e9PWzU1F0kVOeTv1LV
JUe1AdFjIcbuexnF+aMwyIMnuoAxtyZovi+rtnDiZWX8dn2LzYpAQcE+3Zt96e/a
7tUHarTZVJ/OpxbXunBgZtpITzocCq1Mnsw0ff/gONOBE3R3yBPlp7EzVdBL/JkS
H78e2UVSZRg3/Lath8AiZ/ZSYVUv7oXoZQ7Aqj7AYhHYJiHzSW46Mv3aUhw4wJ7z
6b83B6oOYL3Y/Xkrp3cpw6mW+g3i3xtK7VQcZu+YHUrz8uxATAqBMI+wj7RgntSF
WVE4B2zGcyLppV1TLL/5HVpn0s2d63h2OLGeboHNWoDW2uftiCMBbgRHOWg8+kbX
IJGzzm7xfUgDPH0nUCNWR4cy+lhde9zC8JQBzLnvWDQ/G6RuN+tui5z3Z5tkrMtD
aP1sQPCYSZOGRzq75sJZIUuGrxRX+SzxRj61Zjm7FDD1F1MIh+xApunWqGvNAEXs
HXreV++7QfEvp3T9/Zde3sG0wE3GzRu7DA4UL91bRPnANnarQPbcf6zUV+GQZK+y
vhxfwAHHXyH+/l3m9UKrFfgFyv0EFx3A6sRrMkX+J5RtVdB6fpNanlzPeyYJ9Cpw
IybGZVk+wwrep8DLChYMOczrjLnNsV2i3vwo0oQXNNe5kr1cTHSA/H7gRv801UIQ
N0DNgaMCMMUbFzbY2p+NNnT5TMG0/Ipg33SbK9TNarty4l/WAzgJkIM4D2Qvh90o
Hmev4HAQy93n07yyWA4B3vcWowXFdkcTS1jIAMhkL/CesI7PvykwBQ8cblgghRQN
12sl8I8c+jiB98skAKV392wSyznPQQie3HxQ1YV7lJbiwdNjWh1NCDxVb5dXJPOf
BNqdHFkH/c753+W225W4X0/TzncOOpHFd8c1fzAy+m8=
>>>>>>> main
`protect end_protected