`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1712 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
BD0Uso4m3HP4S9U6YYcCvQAFlC2m0s6em5QZNe/LWu5k2WqCepqX8FetIuIWKXEq
gk+mfHw1+8MjqVnPAHevTF4lHIjxkDwHBxXocDwPRrcpwNSvNaOEVa2Ptnnw2yi2
G5gczVxN9ZSGrlvn9HvySULxFmxU2k+p7wFAdIYnkhjXhJ2ZGMFn5sCrL2QSZQTG
nu2gLiQsUKR1vtryGRzQ4mLvaG+htO8n5R8ujNuw26NWHBoM60BugkPYSQEWk99/
mVzl3BRRYw2+649jkn4eZsYMAfexabClL17GxP2QeOE52RK4raESmGkzTqCbPf+t
ISg2yB+EIVeybH3eHzG0kUSQDMXzsHzO09uPKlTLWQrRuyHVqMuI8LAswKrF6IiO
q2/QQVv9kgAo62n7PvItfsEd9oFbVXSlVMlIUdUcLn14U2c24Bjs+BJvTaPW1B2S
GdHhtOWw1nFQBQXjuqZW5LOHKDvlHeqYc+VSicbAwCRfOMECyIraaEiBVbUOVIwZ
Isjd52JfTbJTzRRdwFaOf4Uu3LOj+whp6KDp7Vj/ojIHHq1gZL7ArT2QMuQZwn6s
F66NGzrsPb7qLHjm8/TXRkwhbSN2gCaIPs/sWoWtMQmuMHF28wjr6MPq7vjAnAcC
xTSdmrqS2J1FRhYRcUO2BITaTSxFW63pvjO0SgKCmkyAnl5IMtXRNqFN6lU89clb
WHvIECjN7zA2vLDC/YLFOYRrGSy7QE3wP9mJ9/ShDyC4AdK5OXWQhidkke3CMQAO
0Cjwhk4bP5YDjlw9r7et+1X1H9//bWPbekxqsIOHuAfZJTMIV0hf+Piv1EsoNARm
UiB/ZQ7xbLVrD00Au97YKu9bum0F7ZSUwOboIR7efDV8jbI6hND6iJDoM+MvQWxB
aSankzJEtYllcAz/au8h/r9tC96hVw/NjUmiNlocqyp1kY977wU+cxAOkwDMZfLb
8sGjr7W5H0N+rB2OyGVZif1ZWLlOSOs39TQUK42jaQIFbXykw4yZGHg+EurFmCcz
qYgIi1rnyUgwpzBOmnOVRws/xLoc1Q1ZHmLzzHz6OK2mXKTEcXa6+hgSenG13GLA
bjUVAPoNJFUejEjL5NnWtZ48gPgWlUghzWBU/StP6BWUssD4qjjWe8Jpbdyb3NPs
4bxbHFNU09i+7fO2ZOE3bpsNWx5QLqZjC6oxZSbldWoB3EIRhecVOqEGTkRopcqD
mvrkgFqSmVzsx6jT9shRX8vKzM/e/vsd7VRNEasnyuvFEGCQjnTVc/dDOEIzuuT5
AIuuuvJ8wDw1jkpz5iafqnAExrF6e473bS+p08n+J9qBhIC1o4MDMCKItSgC+Xrf
1chLdsFs/yUshdQLfIIJusqdjx6sqKJl1CBSMnjZhuewzkgMwBsRgReDcnmvSevq
8Lv+/rXK2fEvzdMztR4tbddlkdzOrP3oGR+AdoFxZS/lWJcIXXO89MuiEyF9Abgc
7Js0PxW7AlFpBQRixYm+rYM4M09hnjHwaPQpI7nb77AQvokaeoQ6jIAXtZx7z88N
PbVqSwD5iJWUl5XRP80pKxKdK1ocUselnkw8jJQAXurjv8GQE6qfjxsGtbBkqaq3
ffp6VB5Dv+AR1UaWTJIBEWJ5mythp7QFIaa9YyldGqO34IWMOX8HwW6HC/pxkniU
oEUErUv/P1Xv5ajrBLhbpeOtH7uDbFs8g47ZDmDLmbr0Txlcay/rN9tnuAAVuBYb
KaYTEOY/0rPMLV9MvQO3WZRzFzq9Zaw6A/EAXaNh3sD22Pop/SotXlA1Lcu+5n+5
4iodfpU+tIel5ZfRskskYll5a4Mo6XTse5CAp+iZkXKPtMLDV9AhdEuqk5r/lzzp
LbLmMQAhGVwvNrP3LNKf3Qt0BLMIrvsu6suP5+qji0D3PQ3Zlrp6QmtDqqUvfoLd
sVTodatDcpoBKqUUN7hxCfiIJoO//qMG8VepvRT4l/+ua2HMYEuqjeDE8+IV+1CY
T6UQSyeNcBWKzvK9mgvagFSk2VKxlUTub1l8urufuz/m0TbwggzKnBtTvBn/lIwB
/EBaNK4IsrtADFm3hOHUHftA+9hn3VM1e44vlv4mhVAGZYD1mXEZ7Od3myD64h+A
d1V8BI8MkTD+mWlz9SAonifoy2gPxA2WbcL0HwZxI5Y=
`protect end_protected