`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 61520 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
TDkIdcJUWDKCGvmrQYRemIBv1SUwjycDbhCTRe6w0cUgUCWJL7IL5v3t8SjuLI/I
gQhulak4Omt/X3imLuuitMkOKaGWla8zo0JjsJTQs9ZdttAToI9GohYvI4F3g1H3
Os8ckEXqZQ89ALnPY/fFXpNHNhnB0Qj19Gfeeq9Py2P3kw5CByVOkfK0Aphgt7MO
1RWexg0deElaCVUimD6LLOgXa9VRQwCmhxFZyqEmGMtBfvmiyRdGh/gW0Cxw+nyo
wGY0ChroldjL3jqliaihll0F/AoHbexglZYVl9vvqv0UlXoK4bTDuiYJ4HnoDe+c
icspZa6lcdjAoJ+pBY6hvxp/obBvVRtolOWm07MSCCzXFmDI/EMAW6AGYUFMFtrm
n+9FOJWBgz5cbhVlzy07eWrd/gE2YhSABSkIwtXL71IxvcKzkjLXzuUae4st570l
nV4KSccuiqgo/t2zqbUdSUrV97sJdfVCCjotPQauPGMk2Nhd8Xp6Wi6TCDYY1nM1
QMBApZHT7vYDS6Kz43Am07imr70Nm12bvpnx0erkrEdn3UYIc9egIxVH1SvlGBEZ
qc/oGi7CQdhYML5Q5yleqQSQLIa4AWsyXGTWNOVR8h/28HSsIeq6ZHRn6xgB6Dl0
IwqnoC2tzdLT8gbH53P0phRnn6Lt3r//sTEo8uhGZjulfS8/IFJJDMudy3oH1DCk
nQAAoftNVcjbto7Hjc4g+EdhfjyvfU9s+oRpbG4snquQMO3Xe8UB3le5A1NYEqVL
m4F4mhbcLT9Prc4BJU0rfsmrwMkgfLgGbSTtp+7XhsfUhEsDuMl23NwNODOGpUlW
02Cm36VYcOuYTo47W4aiDyZrALBafWr/UGx40u38GSMvd1qvLEI7y/gCwCrBgrRK
BZ5s3TtON+zX/Ke2XDqwr3RwAxFSH4uQACpiMobWKhDsk8jcNPtLUZ3j3zu+Vrer
1AokOpKzH1HWk0StR00j35qWoS677lTzA7EDjWks3jMh+4dW+bKgtFWzsoaTpWMZ
tZrxEp2f/i0mcHVovzAEPxfT74LxhfJEbg54Sfr5FaeMhBPYUYNRn+DcfxhASk59
8cOvRdHhKKvcWDLQ4bYa2iUjrI1tLJ3UgBYIyvexdRki4tpildYNizVcY/wbsIs8
/OTWEgPvjwr/zr4O59aveB2Tbwc07PjPkkN87q8Oamiy2k5eujTWEgpMaTVk3DNu
jr2PoUSgLscHOXw60VpAS3v5+/fjx/ToxfEKO7btUlXJZe1MRlF5sy6TS8QKMo7A
aXuW9V5w18aaJHQRzkfPH3e/rehw/SV6iWteCQ3Q53C//GDc4fQ48lAlGzliHnqN
mC4w2UsIFHku+w+tMWoU0IaVB5Bkf181G9sbtXtU/8nybT77zr4ip9EQXwPu6EaL
jbOwxKaTek0lA4Fx9oKeOYipWfGgu9V/gaaGUa5aaGA1gAoAx0txLSTury48kJuC
oDX3WOR8CEOUqgmsq9Z9WA6+bTA35TjAcPbDqVZ7DIonKLbMYT8SpgFksLCXiH1H
rv4Pdxhd7BQNKJOFg3kDV8cBrx7AGn1SepdgwHc5x5jm/l7IlcqGeZZOeW31ZD8S
6PRiRSw/S1SZrJvJrZA2KbUcunbx6HgatdYNKXnrQ0PwjO175cq5bv7U+pNJat+y
7mEiB1uEsI9adFMt2REKNr8T6NzBYg4cRZB2lJ2wc2F+IpSD5yRq4eEv5f1Vt4lQ
Ky23OXnSSSnOHgsgM+il4M8FrZE3cLcvIOSeuYaQ4+v2WD2SA7/5goaJdpRuCZWZ
7GhjUlb7SrjYINPD2LBvWSasa4eWQvL/q21AM5CQGkjuqjS0sp6ABXUuzqP6OoaH
R2ZOmNkMuvhtbe9IDUd+sqWi9njtV3GHDjG6m04jEt+nttWSFrB9JJU1qILHK4SC
XHPA+PJqo1NET0VseMwwEE8bYD2TxMeER5VsDfRIXihRqJqEwJZZbKo8k0r+bLeF
eMujqe3hGxlifgdbt+2lXGxwdEJGZux1km+aL41ypia3/5CvGQ2u25IK5YyDjsi/
ggPpIUHReYY6pO8LONvstSKNpBt+8BXnPRiMhRmgH3V9E4wfQXiK2dQbWghWLvzM
C/n+EtCzX+yc3nTXIElCncgj+vUGc85TqurGAzCP7dgoeKNfbm8r0+BPb4FwaoOH
27hzk3Hevu2y7t1Eb7OtANsM3UAcp1mqP+BQeyy8o1r58I/O6PReOqPMCtxGT57v
+rk4zu2tui4/TTVd+QbSQAZWfD2x3ucpUkr7Lk9qKLzLlEnXNwEGaJjYgvVIIrPs
IvBbdTXvbVMnkYh8aGac6a+rNnkZEGXHO9CCPuMYHMttM5qTMea0OBHxMv8rC+aA
byh9RSLg2rBASYjX1HC+oMWLOqP9NV/GYuljbeP1jtcfECzbc85zV8WPGDjaaXOR
INOV8ZLQfS9T+lY7eyRThzLLkrZyM4MdubAAzz257zMPBXd441LzIIGIKTfPoCsw
0pkh9/W9vqLwcuP9ZUCl9uSvHNIfpAYG9OBzQhTr9JdXp+a5dUfEtMH5ifZrm9/9
0hiPBYgDlLNOSVP97xqPYu6oXxVbRi4O0mxNvNUzpkezqTo61Df/WNhkQ3QHoMkQ
iHVf8EkX9hw++2zWNpmsQPOdJWvORZ4RNEn2x8LVmz5qhC467ib0HTuxnSbG6lHe
ziG1aOeSGgybZ3sJG43r6cqOju18V6HesY/MtOX/ng77MSUuR8cEKRCuX+LN8A0r
JZZVeQFrQqDE2rI2EcFSlqqEb8/1ap4ZlJh+sD9vVpn302ZNn6eMD4fKRj/qUeBh
SwYc1kNKBv10iJl8mHAbCuuxfKnYdr7Ex0ZB81c1nz6X0B8HrdAAQ2qef2U41v91
x5nEPfp09HLVdFMZo+K0PO6KaIF/i9ZcdSJs/G2ZDg9mZy2b3dxUK9EtfY4hfcgq
2oKJxz9fwFxvGe6UGK3Tmp8eb3LEN+ydGG7KbCuDFua89rCLHV02Sh+Bwj6XslGP
FmChjxec0kno963KzIHKBu/sPfvooi5OYq7c98H821UZy8JqBfXb1jOv/RDMunzS
XoyNejkcgX9rmhOYEh1/vk0CWkyZcpdPZ4pBsIbqUPxDkeoE3mokvhSTRnmklWDb
qx0V0XWPx/gtbIH60cwG4+FMm17gz2S/KRbrGlxTRoxQ9UlDbFTGrhgFZVG8SuLB
2uCe8YLo0Si/fu/XwSH/+T/HAo0cOUK5ci7Aqv+PB222LieVgosn+w5xfHKQnVDx
bj5o2v4DUVZXEpN81g4kzdFHBZLsI+IoYxzTu/xLpztURMDVSZ8bhC7vRs3W9ZeI
huGI4teJ9nNqVvSUbHPDNdW/oXwtXTKcpubjaIGLH4ld624FoQLJw7al9XVu4dl1
maZHBDLwhc4pUWmg05bw4bCZmKwBVTt1yV0XqOPFvrmaoFVK5jUI7pjlRn9vKag3
8qLrsS2uGelfP2JkecL9BoJMWufmIgToCEt/ag9VEypNvrZarnIRVO2eaWE0ohog
kSAsCDUCMOZBiF5KiC0cF4Re+bRHHs+H1HyIq29Zwh17Jl59DT7PTOOsxKZpZNX4
335Rh6vK/+BVMcfRizy2LjJ04xjoJrcLT03UahHF5JzwFUTENCwZyLAaeuSX9xq1
A+lZttM7lQdw9rmuwT1erVW0Hf0vgdvpzpA040plry80S5W7wd2JMhtzsnZtajrs
UDHq9eeyCsaFLNGcuq8pPJ5UsVJryI1oYbjywI1AN1mSL9Fyo/rzKXnLP09DgGYM
jQbmdqMhsassNhi/ka9JbMCSC9HprlQl7jwDdgwvUTSQYw9S+K5ULOtAFc1NN01u
ymEsIGqzVwNswbM97tOK8lybjOiDUOJJsytnJM2kR2e5ecNQPZlaasXYvfrTW7iJ
k2OcxtuVM8TMU7T5kJIZ6EMS37vUXrcchw0I0W1u1BLyxZhJCn8Aksy9Doo3mwfX
c6PK+c/11wRkTXbsPynqP1f991RpsnB2H5XcRCUoqlf3kyYgjnnpm1SK4sfPHbYI
yIupQb3ef2zgzM5AZmYtgfRSyKesNmx1YW058M+lWzI0gVHGKGKAbAwNPApwx0Vt
qe+Wjl22wHFpZBvKqlYsxclybPL8Lr8CQIZmzGzVVqTjp3ZI/YxI6PkvmqSCkwGZ
ihiqhf7Bl4UJDTlIhPzyz41mMUAaRIJys6z/2T+Idqz0LYEoMTA4oEknlvwD5oWm
rgqO4VvjL6VTrF0jTxhV+yKxtoo+/auBt004Vhg54tNLErIpDzHlDUtrFpBliroS
qJaEbxw1q4dF4ivH2FKxOK3eFgFrh8J73rAsyJPQ3PgK6X17ylaThiOBnANe/UaL
/1ZsXwgjNtbYJC5Ff3rOnCmAK/ZC42frb9r7FOZr8r5BzPP1YjIYOhygspgwKXS5
bo3xlh59P31XsYc2+ovlA+fJ3upMUmKCz6JYfGwC6NurtbUbuYBqM6CT+DgR21az
Z9ajAZ0rQ/eHDfz+fiBLDKOYlz2bU9j8nAOZM1BKXChwKbfeT4q0rdW2DWRfiuIa
riEWj6j5buqXPjOQ4md9iL0MuC4hebb2/V00lZaKu21LBACS2OectaAgh4r2YEav
4tXtR89+ZD5NCrxZgpk976qPOyCwzbROxDuHWpGKOxU3DncoOO4ngFTngAJRkf2h
wv8FgApqzzUuMmMc67RpM3IOdbAQGgfGuN9vRQ4PWyVCDgoTJaj17j+VaXJyYhjx
ZyWj43Mr6QVOzufrRlnMKpCuZLeeBF7V3VAs5LmTWACn4qJbrwD6lPpR8wmpXaq0
/Qp6dtxuRqPsRRFGF+mFEWccc7kDpokEs99Cs0Rbvo3sjRT3rKB2PymYotGkwcCF
1ldDOPP/7jLy0luH1oB00SSvGEkzBN58kmPaIW83vPBUzP/kubS6RGrt6nGcbOcx
98Mo+SPi+msWRBdR19NdrVzEhvySkZOoEa4SarF+LQd0MA8g15soRe5/e6MaOfI2
rZIlyQoBCUNREQSGkMWPhScW44uMqHmy9YT0iXytCyq8KR1ZYdQfQPKPuhTBJ0+u
rbQlfGpJ35uJBFQzUMYYwHb2Zg6/ag87ym/9C7Qa3rfb8/ti1SkrnvHPdcFTkA8S
CNGDBxUIt79CDMTjlnOIxPHiB8rb5/gb4IZjmivIPMaN68Zd4VXQgaUwBBnGz1XS
H1DJeVKKr0NnYjo+ASyPig/psh3TUiLjRJcos0MKyXJf8Z66VqPvlFNjlqGUDRC9
h8ZtMNKyJOEXPwG39uIhz5+b+amoH5sxopVb8ETOBCZgG4+YYlmzfNUB8kLsZuxZ
rT9e5UKkG4R01CStjxjzGuyMy6mMwNneyuarqTFDvzwt1FWuvjsEp52twcOJEvRB
744aqojLICcpUigF3jDoygjP6Sq756bYw/nYJ4E9RUq8zyhFi2yXQafpCGMgmahe
4GZaOE6Gpn3npyxSvDL2FYNHva+K2ImDSlgzccQSMHkas8AhliINaoXyRGN3Df7V
dBYgBP0lMxJHd44FKau+sn7kZjFLLKMoysuHaMeJ5pv+25PKPX03C5ADEjAoIeH8
Wfjx/N08vpNXpMCGb2Hj0rzzJrmT3yjAHokBr1E0dOt2d16W/JXCiEspav+bs1W1
2hyIQVmd0AKzgyMVnRgj4Sj9Hqfjxy7uEji+cnrWXYkGIS/gEIiepjp/CBQS23DL
HJEKetVVDUZrBjhEoGW21d0/65CbgyLzmb00/RbRE19VU7+zARlWNMMi7IZq+MWP
QbmhkNZjJQ1EhaS3JMfoubt9abKIo7Ven4UAj4V3O0jE3OXkYbag7NIQ605Qbu07
3Iim9GP0XST/5wuyHCqUtB1furSK6b87EZnBgPwb79xMoD1OZktvLvcnC4SNW2Ir
c0CR3jGWBvcLNLIKw4T1czDTriW6vU0bztc/hLeOFloti9bl9z1l0EWcXX+VxjVn
hRzMfxr8cYkZZ+3Ya/pvolW9otOFd3X2UvPbBWXn8cm5VYNVTmHTr0eP10flNRof
FgjxeGIKmFL3IGkZd0L5uJFo7CewfEJRF2IT3bI9kR+QbxyUtsn7gf6OBvuU7zsJ
hiWDAD4XgujtDFjpkPpc8K2L8zrbAgMusfOCXnV9tzn4TFGhVjJHdWPwL4YeFLc3
QqQ4PzOuxYmBP0VrLtWshxHInxtPBbEIkeufRQkV+owtHcb/LaxVSsFNhGm5JE0M
ZJXhV7STHqYQCbuq/SVKk1wqleHqtbeTtac0QLNm+Lnf8+Xox2Mriu0qwuXsaHzt
nWlZZy3u+Vq9INVK1umW9IMsmPJGroWchetYo7mSq14EQ1jPUGZcJ8SaeCbKMzcc
nndZgjjxLi/IMGzC0IDmtY4u5D9tZ3zoAkkPeYFVOBPBW69zlgreOxFQFlyIge1S
qdWjsE+PaAxuUhO2jLULjT+fNbT7b647abJWnkt2tOXNo5riVtuBQvKlWHwekeub
HhrA+KEbSd94f/m6Cm9CW5puc/JUFcz5tMjU0qd52bNcDX9m9WUeJygYRH7AlrXO
cA5czoxPIJDgY7iLLEK8VhqfR70Ysx2QUHgtYVeZOWrOAwqxEOEi89LyY6xAM9/1
lK3B//6Spv5ZAoEd4dqsvphAXEI/9wo+McDH1lCF0AQhbzynjc+QDSlc1/uOX7mx
ALTx5PJcansOG9twFrtfIIqRIfqMNXiE98ADO1Q+mcjCwwfPL4+rk7pY08vZeR0W
WehAryMTc/oraIu2XssA8MrJM4rtVhsBT97dmdkTUvQBkZHYyeSfyVJAE7yD2MpT
gfFBez0/zBLtIj1CbrcB6CvmdZ1FoHCnGNJo0jzeenRiffed/O4P3hB44i2l8GKi
2ijlafDFJvjMb49allPWvoQy+lpHmXHGuAFUMPzZfgdGmgyHUfqcAHY6rra0PFik
sbX55w9JRO+zai15qqqIFSM+kN5PXX1W/A+qTVYQhAfXL05euz6Nq0D+YEaUGnww
mjfWMuXBKFRhZWpow3UxVf24ppqjUfUsgFtrOaAxOJNAOxkhtIH2tWg8jEZ50pZU
3vHDYGMSFrvNr4iJn8qWia2oZvQI99fPbak8+qSZ81gdFxM8jhrxSmli7WuamJhA
ad4gcot5g39by6iZElygln26QIzLrZ+3UVbOX6gA5fBmyAcOf4TOvoI+YeStwiMw
BfsqSyXv2rCwbTV73GH92FgDKZqi3h8hvaUcW9753Yq4z1qe0pcmS6gcoIrF0A0x
Agq9RVBHwd7+WPEq2yys9R9tQTpakM9eBlu8CumN4oNcdhqEP4GxFqnzelMs4pSD
vcnR2OdghoUwd1UlhgGyc/Q9lTqxCDoiYQ/bqqweRQnWljo0RxOtGN+ocEzudy+K
qL9DLkg4aXc6nRSv0rbHhs5PaHTNTEmgkTz1C+JEFCxnDdyus+8G1UC5008dfrHt
AZ4GS2KIBo6GKwSazFdfHjdQZjy4+DsbQDkTAGocTO5nsotU+Aeg/JBFc0lonGYx
QXxuZTnQ5dSSST4H/6im+BJwhs8ZnUHCV+ZaPVkdLGE1jBf0zBzPY13pg4n42k5d
P5Hlm2/u9JONElJUS7UpYZ6fBpkDH3Sktv3Tz4HRkkqKM008OdivlWqpZ9CGEbMu
xATPqWHTIu10QacbOOUUy6PNrvaPsbuXsKG+vxcTQcULSEGEvvcpcpx7lyPMVfR3
bmvG4S7DbotHQz1UdeY6362201hjO5dIQy+Y+YRJuH2FJ3dSab+tZSq6v5vqydnm
7dpWXVOeAf8WrzYregEDC+1RMH2Ze/Kt4oRfbHyMIyFcU6D1hoYDbfHeLdb1GfpB
noLRk4igwcCOMou+85WUSG6O4ErVQnZfDBwqL8Zt5yTww/BGq9GU8i3k3kL5WLoB
gFRdHCjCNVEcyJCIL17fDSVazzVFB99cIWkpFiFInx43VRiw1AeNLJ1+PAzT1kHX
nDzeHOYmZ1M73cjw883gknB2kjkn87igd+m/sbC4YGBJ9IKhp80oMPsnF9yaJFEy
s4BKxvk/5l8SpbE0LiPpgaFCyB9caQ1lr+TJFdtZ1l748Qd5P3onuoJ6PVcVT29s
YxMzECpCtFu+5GEAx84ccVFONSFFxqT7z69kSnJwIJEMm/IgxXQpADkPsuLMZw/V
Q5cr9GHvPP4BcopADYA9vspI4FoHkrZBuxKEaHCkPudHPROTwCqAU+/hTsehgWSE
883e2eu4LTmNL6wq2Dwr/BNc/5ZrFcJOr+J1LQxxjq7CVossA1r6vuwO8K1RucTz
xml5nCFklv+XPY6d3Z31JrXq40/iuXisgG4lBqGJGrx5cYMdTGEsg7461CrP/8q0
LLheG/He2tKLKrjtznKK6X8SzlzckVIkcpH1Kl3rCFMfIMdAXiPwMY1WjAq1oB5B
d1I57XWc5kcMIwJrbDumKa0LzKWEXXXtKYwtwAKWhUmZJFLa/rXXr5TSr4u2Rhwx
3rrVy/iVmA9hNzCREF2ymYueh1gWpLHLSrE10iXow30QZyAEqQtzZ5+CmWPLIhEB
OwoUXve5tQgOlObRZshF+mP+DkBWSCKKyfbu7seoqJ97OBCTgfvojF+HkCkYATvu
A3xFS+lwtrMW85glGUdvHd4cKVXUNrI6AGief86F7woRXBzk4U7gqjWbVd+0sby0
Bd62iFqVN3ZOybTTk/457VBg7kglnh1EIhwR/rPunKpwT6y2Nthg+1FkB+ey9R7l
EuseL/i5KCD58KfSuPD9z5I+u/YFPjSaS4pTXA2G9DQ2lVlQMpaTinuaR2en6vCH
go6QzHC63y6rZ5Q1orWbRYt5PFB780PJ7ioOsU4J4PHxUPldQjzEhnwuq03IKa6K
RUEargmnRAP+qV0XYjHUcsQwU3OkLcJ6T0UK3gUC48TMeyYDRbXlF0YVx4pRPvgW
PQcumd/zJdcxzQp0Bx+ZCikcFn1/6bwvQ2kaSx7bIfYZYpf/FStRA0WOg6HdoGcW
banFe7R88n5lYeaTOBEZimrYRxG2GI5L5dmSfkATUyBgcVP9y18PTwPY+yssQ1V+
PJmWNiZAqrbW5dbtAFDhrx4wFbCyTQHNZ08h9T1ENDplNy86fKVsKuYrJ4SVPKEi
igAXvhm3HUaUuN9u7PHMKz7KuHINuWkdbhjl1muX8K2ZbzLXeP+wxEc33b1lrGWz
ofR3o+C0FdfZ5Nzr7+ixn6/kXaaPy/qgS0WwPlRNG72otX1OOSMOZvSnvSozb5a9
XTEmuC3iIlayrjx7pAA2gNlW9/nWwRSroJBRrtkMY3iBUERNc9/qf73sV48lDyHd
5wxX3upaAwR0j07wXGpgdgOTkqZ21kFw02k1sr9bSRxTYkkcRR6wk8IJIyn8CfpN
Sk8pA1emLvjPgHev986PYU8Toyz1TdMdpv94LUjV20Bqt4+Qv3j0xRRWmLSBe4NZ
qqcQYWW9V15/P3ZjuZSS3DOgwOj4IUKC49sr/9Vx/cXpL8ZoZHlte9SMFpnyE6+8
lKEOPtiSHpneZEyn1p4Lr3wuKdx3toLSR25Yz9cLu5CRDRs4M2ZYqHCnJfPJ14a/
H9DgwoPs+Jpdzc1tExsDDHhZBOfj9vfNvEgfyWBwPCnBDXwkZdDBHx6T2MJkcStl
zLLTfw76EDC9O2GqgisyZdNJ9AehbzSSz/pnPkBbGeaVCLbni0FK0Rc0u4JBMN45
kFepNvPNCRGRq0WbjKN5mpiFleZAsajx5TUjshR0eyFoEODDErH1ohkZcbyD8uVK
3G4zkx2otV/X6d/G8ewivP7C42B6H29j3Lv+kcz0lioDX4FHmlQVzgWZrwL+35Pn
+oOs2pB5msL2MY3pkwdfpU0uEmAXC776TEakgmRfyzVZqgdvUf/o6wfQtV4jgE6w
R4OJeV0WfQi6PBbAFtn3PBiAJpP/xQImQKnvy2IFukosQKuY3v5CUcKPBJFi1Z/9
6+GHRKkRt6Jc5EWCUxbDX0H4e2E/T/LnykchpODwynBQS2VzUmpd+1UA/anZs6ZL
1diNWO+/gKDrC7MmOrMKcqirdKtIQIDFfZqy7oUSx+wOpfJ4R9VjvjCVwLSiMdzd
6d996F53MVak4RigIJs2i3vwLBVO98RPeN1VsHyBGkDa5ltYyHp87/dcvsYl7g0h
/0Y75SMveFMh3CvmRuYoL0LMFNNDxZP03bPBQGLesx3FBwcbtYHnvfVaOS67kEJB
IvAmRHXYmolnG1mDkEWxd2lxx+JchH9D18CxO1iv0GJ9H89IbcQexnwJSxlZt325
gQxoh20O1VPZbfqJV/9T3G4B/qJC5Dytgj1+yXzuU98rO95ThuWd70ddMdve9g6B
/bHUFmiYgE+n290MWsiUyZ2obfGh36ym3zrkR8OVV5/S2/ki5o7jN57sGjNnWirY
EBabrL6YV/Fq8wVhUPMG75b+WA1qIIyQWP2+YzipJ1x22exC/PqyIOac/npQoBb9
gD/rTJGPYrp1Nmr+np/+L042detJhKCGDJpOhKSLDr+x5+WpQnrcGzVb21RibbNR
+kGHvp6+40QmvdpMK9ZkWVBzhHv8qxyIFPQ+kHOty6ctDuXC9yjclLgcUYAMQKdJ
nS82CIYVQGivsNVNYsA0pbAOkPTrrw3B9KDuNpXxvYgf/zWAiSLXv5/5P9l7kGjI
c9M0xRNnnIwXAPrMIwMH9jfOnCtsYc2BPI6k26IfYXYFom544dw+yYKoTu+xTT95
TyCbIkEu3mxAlhCCPh90yxJ57Nn9NfF/iWPSFupFYrGFF14zUdpEi7B48IYYThmP
KxZZlXSUNXIe+VE9tcN/pTBYIqqyWeOL+RlnJILMnvayRuBCocP4UyY2/Pspj0/2
yqnA3BBC3HZpULCE7YLN65TMD3f9PfnvEr2tRpFXdIrRhgmhmVVgiJhyOOm9mbBn
/gnfrZX9DyaEbo6LZ9/i7SYQkGTtfeHvOI19dVlvo7eYQM7UVE7F+a4TR8+8a36t
/yLW8EffPhpuog6Wub6ojAcXHJ7jYcCvDKiTu8b3ACcRhMreNfIYXm8c47lzbDGX
gBSDypzQDODnwW2HbtJhsQYdoazh6DfMXt4k6I6NVa3Ps2d7zk5s+PHnI0jCLstg
DIRtZ5/sW3hGx3jEzgTffbaVwMWNDzlelwmzLD6pSURdUZ3Ioxzeh7RaxfAHB3Ni
gQkVE2ZzRaoT+mT9iwEEpm/US5djhMl5AiYcwwP6mby24RQ+8Rw4l6x+tM02EKNN
ScyWxITB9GIV/dWnR5UPw64Wath7EMq3HJOe1/CcCtzQp2O6LogRsjwTl0VNYciM
iSvZhg4eta+FTNifeC4AhHwTbmIwyQIqBUW5Rs2AU9/4LntOH2HHY2G+mxHRaOwL
SlT0hYivucTDIj/QRRh/74E01DqPxRnNneLcvsEa+iuHc516FfTaAQSV2EX3FL76
MozFDvHBBkKVMUonKLrQylrzA4euPqBPKxzKduK+jGVMRK+SLPqkKXpQuSR6kYza
SvmjF/nATNokWGJ6ZONBbjQwtjslQqBElNk0TIFbMz284VJ7NWxlsdj3aWcG5yF5
+0lVqcoNMyiVngWANW06lnmY7X9OMdAptpt7G2KAyskPHBw5xLrjbM3AWL0U/47d
1v0QgKsTz8v776+9uAzrlq1a4aCHdeCODS5F6NbK2V/rp5Ogot0fTnCQzp3mIFvr
sPYFnnzUVNhyhOayXG189weWdfXiskjOYYzVadFlJhKSaSEgkNeThtgcZB5bbvnl
Jz0fyf3gBpQHVzNLnjcCKgNYsU2NyPW7mtrlMNAsKlcsHpRK9KjV7zFAfRSVVXVN
j6WeyFyRA7DiezXiju1SvPP2nArGBbNMesfzhLpFuEPsIe2i98zE1uXOt9eHQWij
Vyb/g6IBResZ6F56lNKv979dH+FegqF7MMqp3bXi/X6jJwJQ7Q6MaVAgZw5SgLgY
n1Em46K0KC05aV0PKSJTDy+dNVanr3dXlfhpCY/G/XSNPVBQZOnqn2XbOgnAK/eD
wzmNEbHw4GJgF5FpvLuknpePE91tentTOJ+e2fS+DcoYQNQ6Cn8iSiKQfdTLCWwh
HcwRDp4kS1vFtDhH6Uyl/zmL9JOF8N2U7IXUjLC5Dg7QBrN4jo6RyipRGCsM45Zx
JSqUSXHmH3eQouwXiyQF0AzfZG1TP2R6JBMCjc5cTloX+ClZaLKu0Ptxs6TzLyRd
m5lo/waYKxMAqO+BRJz9essVpdKFkQg2cmfIU1oMb56+Y4kdvnUteNyYh5xkTCRV
3lPqO0csLWTvpN2VDlUovrkCP0Y7debcMOE8WxL8kheUljwwiyD8ybjiCv2Y8rgA
OJGjpEQ92x/nMfpBQA8UAEJ6s07WBzFqctnpOhN3rKFO7n/U5dZyvNUqrejptXHT
9jkCWY2QfEpvJnoW3smIV+FW4oI4WTgXwcNkBmeQ5pdp0hYSLsRwC+UtW5/1pP9o
01ZVh+wAI3V64Qd8K5vhoXgdLo7IHs77k+znEj0L9DKg1HJhOmcAKpeEljfJ+Yut
9SN5Fff+tPzkWhYcF2hl/qFLIKP+3ya3Zx867XdwADRxA6XWrFcEmXSsA2cvMXAD
LVLAzMij/OKZfmS3/RinsKIr4SAsYfjpCQOZF7+1wSZf5QAuYJpvGvAIu5B1fGWN
EmJ2Qg9Gcz/Bzef/8BSSWwB1n1lSuuO+xJ9qKxSfp0QjbQ/Uw5glCu89c8gDwyU3
aB1SNv6GciGmU55AEEXUXvKkwUzS4ZvS1CQzHTjbVSVhtmzXXPl5BDcZSWVD/953
CHsDAMaIeKwBK+mkq3d6dviUCGn3uihUQzo6vn1A14TVaHf0avWPhTwj1fQKebZf
km//ikb6dMrOufNPHlBk01DLIM5+0T6oh8d8qzrBfwioTbbM7N6C/740wGh7UPHO
sCdwAWd2ecq2XCQyVmvgd1XH5jl76mAbC6gRbMCHm/+W6IflHSAhafKSehmrk7sH
gz5GKJaQaDr+wiHjxu3quBqaQC9TT65t0CCvHI8PLdbpkA2RjBj30xFdD0/F78zl
3gKAkDkvit9+Cn9mt5mTSfa7nYGrDpLB9TXiwzsnOF0da4OdRLKVPmE1Q9WxFhiA
XwGLtcrUXKjNrKxYEcV5qX5u69Etf4b679KnBsJtLPXbFVsmunSoJMQZt5OIGXK5
k5APGmH2dJ9V3GB9CKkL1ZBhxFMb+/DklPAaXyS0GbGXBARpl1rG+G/fqscSjSVr
6Timyaw1xUT3CIgjXYepzzYgGY5FissUyuIKoNSCJplfuf13k91SkxCxKNDbRSEl
K6i50XTEA60mhbXatKBlbmvavcUWsrsjMOx4kgJRa14EvTTOCgAzu0o+JOMXi1CH
LOoPhYKeOM1HTaf+25kXOdoaJawWGPcRhM3CwzH9aWkliItNpG7rJjeEfK4c/uIG
PeFft/Bjzo3gXZW4uPLHZJAswvxpINRq0Ag78xGp+ldAtysfBHc1IM1v1lbvWD0H
3CCtBF3Axb5/hiPzz0T8gqqAuqhmCJ7aF6RjiAERuBxE7pyho8wDyDEVMzGo04n9
dNWSzOgZA2OgoqvkoLOYcvzEhxXiPz5VZzcxntRdgnvxRm+WVuZOlqC2orktM9uR
1qjzDE7hvAHXHXvvfWR4m90VaGO87kk/PqmDrpfd/rbn8Wff7SMjR9PK62WtEWFm
Z2kK4PnPke9WApA4C2esvoSzDXgJnGNyC5Y8J21HvpbwXkhSPNHH+6KT5tgyXA65
wld8Ir3HbwIcz4xv+kpbPBi5EQjT+wCv1hff+qy80TY7jxKycuRSCPmitA0UCd1H
qwcJnIt+8yaljPJk6aHMJLtnGQsFVEIbs9XlZr8JnP4OdrYaum+6BgiF/bd9IYo/
8dgiffqJiimYNbZ07ErlmgEDuaSlK/zi2BoPXVjK3s3xQ9ybd3/B63hQIIozc5tU
BcvPpDeC4lgfNCBFDWsdjGURC53fFbxYecZb7Wmtz/PmN6WRH+exiYvhQZocuIV1
jvws+4Gctua0j5CwFfEmRAXU87u733IODfrr/RpUYAjE6ivupbMeCUIr5i8UUeVs
5dcnKUF2agj0UzTTjnnmN/d7MXb1oFdklW3XnTYcBYh5rNHY4V1SCyBg1IPlOx1y
+DKGamupgTKdUCp7eOqk6QAEQxRBxGt68TVULrdYwMopW5jeO0mMEVacaNdq6kwp
7dfMn08MTDaIls8utts8gQuEWHoz7bTwRQBkhuWZYWL1T5nNLil4Aeo1OV0POZ/i
zD/AbXfvrY8z4Y11WDcfNXpZZoAf/toA+MbLI+Ci22dBRwGSEo8X/hmeEYn81K85
RpCDWSA+p1MI7AVtxsetYSHwEBXiWjo5IX6lWR/wdtY5+2Hb1yevrIT58XM2jvqL
qhSCP0ZtOxEtj1XConoaRldU70R6rYqE1znq0lq6uJgVn0nIy8RZWk7+1MSqhYjY
f+X9zBgbd8XuwZPh1UITBU2+qt7kj84fxOWBf38SjceJVNlhCmTQGUO1IV6DRtNj
MrkMXhUayZ28ZYtqtre7Btn24PgKmuZWCyRqUroOJBHcLJvYjXJFss/FOsyI1rht
Pmu5Klq8Jz7qi4Wsf8eIsDNPh8N3dezvrzuh9J4lEcHYBDOT3t+52/VQeClu1yfA
+JNdJOh4/+7VpWyXURY9yH4vmFj/ZMHlPu5QCQtMCSP2ecHCngkmMff58lVJCygL
gyYz7Ioc+d2lbvanMtXpQfM0eTgceNwPyi5Ph2jlQXiMgboF/rZAoeXCHQfFMUa8
K1RTDNaYf5wcq37IalesY/dhl5sqfgZy7A//+PbHb7ZS8V6wXr08TZCZUgACqO1o
/QP1Hj3X+tzlQqXRnH2hxbXYMYUYsqAzNqiNBO+XuV8WHBmQd7K55tzSnOCwfpr3
I8M8DSuhKymt1G3sfb0HIHVAn88EgM0B+f3AKnbolKDBon7T2zcEQLZ7shj2IypC
BsOCDUac4RWDLzt/AFk3HKH96/JdmewlE4ZEx+vbrh6XbICkQ8l6AYY4VPDsCDmx
IolIC3y+ZxpxW2vrMl0fFHPs2V1Ut0QhNVqxLVrjTnwe/fwWt/UzOgI5H3bjU3ho
/IbbkBw//5nD7QoNpehkqu6JiGg49SY3WFb+9W0qPprbaD5g7m4+cBilT2DnfqCw
B7wRPmKQhonwaHRM9h1+p79z1LWr5f2etIMwlIYt0IQ4h6om0NzfRQgGrFPfooAH
Lj1w0j9ZAdaeVOorioZtrJ4FsvYke1yYnJMItF18ak/zo5AUQp8n/cF/2rR25D6E
wjj8Z1o2DeRDjzmzAEd3USGFrV+Dt602BRTrySZDyUZ1fHgw8iTDIkCQHk2FTbmZ
yDHwBANSVckpAnItcqsr3RmNlY0fcGfeO2FnHytQPBguu5vrxqQXjtkctS6BnIhd
C0uG2gDLVY8mOqEIjEpxfXQwu3g4tGcyPVa/h+ShvRyait2l8Za+SNTISlqUdpDh
bJICx2QeUCDb6BXlikwyOA2P7hG/AztWO66byPTMSE+cX2NNi4pe84/NS1kL/7i+
X3ChSxFyB+wouP8zlAD4HRKDifj2J+0j5IVA5IkTaqlh8cKO4uqWvEJGgwH+O8QI
n3dPvad4DaU0RfdDU3lP9eSNbvF+7WPm616uDpkVumNzCX5aH+NkOshodUpAaXHm
qvaJeQPYi6xQjasS5Vx3Cwbbxx9Om6uKBkDp8+Tz5DJkJNOgPiArgfS8dODDFkrg
AtXtV6RBb4tCB7mqYzAeFUGl/cwb/2IuP4CpcFkXVpsr5NrwPJ1EAGSQk7aHzUWa
toDiO1pCyY9MHxLYYL6P5fw4cuxenMSGtNPhVK13+kfIyHePOL1TqxiTa/jF03v+
QmcdRUilv5s9XTCzp0qI4y7Iz92ALwWSWhgiIwstQ5CF4Bzm8J7TJnQ7exaDMaqd
t4N9HvwM8Jglwk3vSosOUEz2UAWGmorca0Ag8m3oIl2m4vC3W+uKulwcWNAMexy3
qkzRwj6MSlw55pj0OHhsw7mImx4k3MEL1RVR6zcQpW/BTn2b1LsnAw2aOv6gt5WZ
qXNa+zYEvlanyaIP0dXem8eyV3ZVL8ozpmv1auRDFYOd7SUr/G6qgKPOIiIRCdO9
j5/uJ/CLXCb7kbok5gHoftV+iMZNN8fwsbca9kgpOrUQy7tx11F31F0y9XrEJt+w
CPrb0mDSE2Zr2uXm573htoc3FStiRiQ2kUkMOpCGqRvzGRLyvq0GXZEGswvjl9mL
kl7HMkwxsdNWLxFFuNZ8xK+XivoE5IU9+PLYK3jvES6iixM4GSC6wNuWLUC1wZ7v
pHK6l7Xa4BihZ+7cMhYx2ETiliq9h55v+BUhtPY1VjsJTeIJehxIdam5yqfxHKvz
4D+jkCiER+OiP2h+Gt2eJO2hE2oe7ryaqHm/oXhT8dIjKqeTZFk03fDtQuoUfLL9
TqkQn8P+WmYudMOC3cbTNGwACLzNhIen1ZkbIik3Xaag/eBfSbRa1mU0wXsqE7UL
2xZg0E6hZ6l82bDMqV+gAJm9LhjgSyj6kYQQHmdee2FPkggE4l5ZLqGCPWn+q6OD
yVEDjHKEMWwBCMXZ2gfgjWC42RSEjHrI/AHMktNTQer5uyi6cwZOpgyyexQv7Cgw
tekKTX0x4FHU8v4HfXGNU5wEz/V6jdbKrguDxw6WUBVPQRtuiYDSEnfCIBhxMhvF
o7HHv+D+aFAaWrykyrEFj+yKqNHP/6LGtAZYJUUPxrBztXkWQ9BFQ8ICIdqWAIn/
jKBYswUJ4dSrQ+fMaX7ZduxUqU8LjguRiZNwImhAwk1KizW50ZIzTXIJBu0CFebE
drU2F9O1UT2fSQLw10ADtD6PtyWAcN2Vs6KoQMYCV3l7cBZS7LQHpsTjB2Ie0PHS
fYfeaJk5AyO8GEdLAise8YUBuFLXPUHJyBH55SUbGPld6+aqvfNrlb80gzdRXwTx
mMh+Iw26NXI6Fu2gD4ghFWsz6fHNtqkulIPE3KmNyr0TcbVcpydsT6o1TWg4JU1E
ZYTSNBIM9QYRzez1xuYkuSCQPm4D7p9Mn9KXvpYYGSRFJeTIhiZjTZcwGSYVU9W5
CzSDTJPJA5qI4fuXSTuLzkKgkNmgaa5aF9Y+rjVSqdwzpqT9ou+sLnyrso7g3qji
p/IvgXMuRPXcKF0YQdtKxKr0OoAYAB58apP+ioINefcwiZBqFgx6uMEBq+o1JQvx
WlvPOfGRbJYJkCKcPxV1ojZivcX6DExquzemJ8X0ZNBrlCl0gd51OrPVQtw5NK6r
CjXSuZro44RmpP5KCbKC7mIx+in2ple2NpVnlS32wafgSlWFyE3jACWLksqn4mLX
T3G9AnWmvxWSR4Mgy/8pq+24VZL2mNReJSlyufBEhTrFD3eSqSu4bpvGLkHnmN5u
T0zya5DnWUGjSBNlINHWodY/mpciz1gTFCB6IeH0VOMGH1Ca1zVVCCigPxoKIQxs
SsmnSP71myRgRV7J1SZyKjTp7seOnS0oIXIltihBH4MjWecm2AkD0neYycMMrh4z
3NMvoZG6+SDjnnSfLMmV/1PP7oMWxj+zqNFqc9Kxr6pgijdxFMWuOooyQgVLuQFS
SBKq6B+lc2XoFwYo2bIvjbPBMF9zgVUfpSfwh41kEqB/mO0v9jXaSTOJyUmB1hm1
N6ZM3XaHKutbATjSKEWyYIBaatk8RYYgRv/55itABe6+1IMJ5sp1whbJM3l8oNti
1Zw38cezp6HF2yz6TeTFG8D0eLgdXP4mFk9gcjkqUNsfmtBjS0vEPAMc1YCBaipQ
wAiH8DXmXkQNrP0+y6cnQ2XLa9ANmiupqHVbsHG5+0akCf8uUU+E6aSMO7DVx1hE
kJeLHSHXRbdiiwMfb6PHzlbeGNlDFzZGrKXCaFm8wOSR2suoprccxjqn5YHLBVeQ
iKTF4bdplU6U5ZFLidCDn3hfos/cArHriemUCA9vCzlCcuZLy65sK+B7o0XsxJr6
xl+4Mlk3TlYLa+Tz6vj95vst5dJRMf0pszlcsgjdsoE4N4Pflji3qsrSbP+M2mBU
hdaNVJr6FT5/6z+FSwJvRZ5xIOoDNJG3lKOc+GbzTjWcnxdq6gp0tbJ0X457y3Pw
sehb9L7DQ4X28Tfwox2UYQGD+yfS0uLn/J6BivZPBeErVOdMVBAqY3qc2OfTa20w
HGBFQ6qVcsaFxBEVcDcW/9kURWGXRtmkwkjXfpSfkJPZgdwdl/xOcvFmYbwJLfzl
mfeQrz0wsSahi522x8lk2g7iZ915y/2LtOYH33L5bBxRoXj9Ry+ATQrl36oDTgn8
VxRNgb0dcy7DqJeQpGnFKk+dP2A2FODK1U1KOoWavNp2aBKjjbMO30ccbIPUkUrl
IUxhVM2NDdvPBZok6qMv1rfJnJL+fN7jLqqFytqj9mUW3E8nvfF7f+3/4zRlbVyv
L55dbDiF6jujIgs/h+lf1ObLMr3x7pvc20JfcHmQQxRCrRXgFTjnpk7GURKiG2VB
aYj9Gi08pPRwBIASkNi4rA9NfXCnl8MwJ83yN5C9bTHfYoVnwlL40cJV/lNS48Oa
mjSC2mkBAFIBbwhPDYcgO9P7uJzLwrx1UpkdGYQzoCEUTF8n+Ok2t24W0PM+TFJw
mT+a5At7PywsQop0u1lKwphspkW565LQl4Xv8SHWii7GxhewT4amOfG/m0OSEg86
AtNu/72xVAgnvHTJ4WD0LvS2pGELvZCvGbY73AaBSApio05zu9Kq9CDXzMZ951/0
KG2nRvBs2o1ao8bEyp1/JU86EfSiAawKl7MB++/2zxfcTiG0ppajxc/u0ivnhUTw
QlroFPzSRGCkLbrd7/U7hmV0/8qcituhcVmCXcEo0yn2pxVF03j5kjcwihv2hJGW
2k4XywX9BaA7JCItB+S3IS/49wnJt7Lnt7qJMOKZyLPQZfgcrKrTctWZc+Sf8rKW
78dAnXWHmx4H21+NVxAR2/b7N4c95t05PbUK2ZEQwgtn9rkADePKiNiwfWGQC8jR
JkU5f0hbI0rWtIDBSEn9b2YFv9JdT3zbvYkiWmP1Ig0dqOOewZAWr0OynuB+FAE/
0njTCwp2ALbgHBqwwWUkK2HNMTA4LwVWD2nZjND8XnWbjNn+S+FsdieihcFCijT2
P1Mdn64n1jw3KNYpi2MlC1Xu8JBaH+pJKfoLnsntfH2YGNuyw9mhOYs52gOyaAED
wL7up9sZrYDMHjimmQPdDbRAyaiVz+i8vfhdJPVdGP1kgpAp/MgVPUuIv4dKTTiK
rxkWmGYw3X6zzYr00M9eTYDLAKiPNa9IrzYSHz/CLgcrHG7XR3wjMMfAKXP/BAAg
efomGFKU7tqxbPcZHSgXTsMTWZhhm3DW7GrRh7y6vmVN/6JlwWHlwnMftKWLb9R0
Ii5eigQfJxwuP6I1+ZNyXGhjPTRXJwYzHl1RE1DI/fOu/wXunwiXNrkO28aTYsgn
iAR/EbRVoKvv/FycFzLAkzUyStWOzyZ6h9JAH2nsAtszAZGKYu29OyAjWQ+TyR0E
0gGbfEVHXXxQuuNOELTyHyL5WclKmx+STpxxQ/bX1eMYrw3f1DZFYYW4+T6iTRC2
R3cJtUndUlynHtEPipSXNDQaPqQwSHU+RSTKK50UNhQrVtTTr6WjCznu/jaKls3i
BnZuvAuelLy4ZRqO47Eve9lAgLJ4xVpuy0UrEcM95qWvuFfBM0nuyCE0RQVkDXa9
vYbScZASTlLnB0oD6IY67uQfiF+da4iOWQ+xP5V0xeWZm4jJlIG5RBq+9Q+rV3Dc
OldyuHcbrOpXl1PgwswKOOyOfq8ZbMv6T8fb9yLNGlXenjNqcVER7motKJyArdTt
MVRutEgRw+3COrVxxpn2xJ3Yw8y45+xbTvSuDDlzly9noBkETP2fOpKwazAEHDsB
m33QhrC8n48yF7c2R3IO9nqvjbx/NwtwrzpVnivwYdMW7ZP3Y4Tceh0gulp6oSBe
uR8P6a6mvh/SVDHI8LayRfr31pLMvORqW8pUqUtc+gDaXM18AuDLZzSriLTYqbVx
bIS6Ym9HWznea8os+wDan1sS5cm9YuJLZ11gljbkeMer/siYt4gZWx4r/7BQTTx3
xPTxq3zzcvIUh+LVbye6Mllxbq++75Icm7PmvsmAnqmdSFz24IIRuSpRkrPMEUdT
qp8HVOQPcRbrqvnpe0K9tj1imhcSlZp5LKhsJWpp0MQbuN0YxK5RQ6hetQSQum+P
w4XsAeNoJcBEGc40Mis5z3LhaTZ5FG0HfYYBCj05NB3j0VbUL/vgs9QODPZxQb91
EY/Ls9DFv+a3D9c82eQrQ8asKiZH5X1wl//VfQOpXmrt/mT9mtb6aKrOny74hgcK
e9ki4VT10WaCfSqTezWeLtTcAo5M5MNcqvaqO32DbUK2Wm8GjTQYXUK4U26WWA5t
pkPSU9s2lA7KqGgx1gpjY0UTTVhuXQ0h3zMHrj6mP+GU799/Zr3FCgHBVQXAjQ9Q
C6humOYUhkYdwXKSNgsTNmml3BJl79gTm7PHWeuXllSMHkDnXFUqNunde+5PrOny
WuJmi57XB0RmPR9hK6uk5EGg/68H2XFel3tGK1b4zOFuWAGJNN+AOLwMhOYVhAQa
oYL3wNYY+NsBaLqR42gJ2UXUdw3nnvm16qC9+8vClK5W26x/fiWoqE+eq8BLQX1r
SoO6U4BDRXOM5AzabOKrMgEUwiOwNerCItoeMRyjkxBju2dLdjSX/LwWkGwIoeMt
dHS45SSo2Wcb1dr6o5I/fQ4sKGbGY+INud9E6Y1/Hc5rp+bLZj12Z5yvNfklfXos
ZhMFxyhenscvMuZm84UQPv4O7cttgtu5ZSvLm2/sMU4Ycr0F6a5uzJNJP2IJpYON
4EFuijj2Y4JnvzWRIbnlgctHI35E7PjGugc/sTuViVrcrh9cVTpOtzQIWkqT3r94
Tc1ePMWhd3ZeYgTFecpmG0nd4sRBEjd3aAPNoigWkyCJSptR0E0fCO91qYXy/1PI
8MdWBm6O5zsPO7O0IBJayK0P/9wcjlHZ73IzyO9OU5g9iPFjnfa2Q/MOLaFNokoD
RqTu/yK2zKSbzcVZ8TxOAd7JfxtcwA5vvjiGp0NZR/eZ1ecZpRFbwU15Du8jBfkw
w9aBXnXjs+o/VLVlTOuCfAFBDgbMT6i4GdueBUzSrA4iJnZT9pLY2S7ELjmxGgDl
VRUx8xJ+US3w28EgPr5CFqXNCK6jeWQRz/GgzJS0ggTKgiG7P+oPrfQbe7pxUuNo
8cDUY7cuUFMVAD9ipWLFvmrFSfhFVDDPPw1zqxvXL6t2Vo8+Tyq/eAP2w+9+QFus
30bShFPK6F4omL7jv+0tq16n+4W1CUxisWpPEqE0NLeeftdymHTIoXnuLUGLZL4l
Q3nnLeUyGdKmcnsadARivhcipt7XK0RM51Ck24RMSRIT+XH7uWZfkOaBMng4GRir
WjmgFgIrJ7K09TsYUpLeqowrY36AaOOn+7eA8T+yOT3XiC53dWQVCXWKfJLcmpWp
TG4s7HnD7fcRxMCquAS6g8dIKC9igsQr7IaJcWWZuaUagOdJMLVKZlTfENJA2mXj
wtuXB3d2FhY3drv11+5++Yn9rPS9JVCBuWE5OTkigNMC044LAuAhXmkzLByFkCSk
vHulQbj2cCLIQx0ihquRgDSE1WMBYxeXLGWZpwad8GxBVLApEurL/gdP6RFRyohF
aT3C/l99d0GjAMN6FYipgXZv50lijp72J20n1dmRWsfu9gj0k/3i21ByA9RATYIY
/FBJQo3H0Qyo9ZGhaqCdENHMcPH473XmkdJ9filrTwdS+I8Z1FAtosSdw+ic69x+
Mj39RPyj79QGZhlAaqXPKZkB0jGZWZ63Bg/wMkIbD2+C1hq3/kZCY92QntNNLVt3
x/p5oADPN43BZfYLvb7fSyR0g+z9DnMp+zVz5ptMsZfcVN0Buq17dBWV9nSyXq17
Kga1269jm0lYVzkv0kmlHi8Hy7unFhP0eBEat+ZsHldDyvZiMqKb7Lnj+UU17RfO
x+TkHpXDfYqa8uqlkOo+UCnHc7dgoQufVahWrIXIvLSDYGguu7vBOTNt/QfFqlQy
ZEwfQD0x5dAJE4QjT+DqbnM+20n3yfpZ9e0V3fAaOjMdg7Am1rFQ/ihHZcyDFtQc
TgUNSuzbApyWxRYuxkkSpZsqMOtjRfUhdY+3K7stRQueZi/18NEE7GhWXyitufDn
Ux5jkixIPZhStU738IpNZX1D+W6RS5mUtAQxwtH0U7WN0+Cu9Vw+xrONVhsqRNZU
zx6CJyJbIFd/3tvsFZvzyoNArHOLHDr4t76P5KGXnbKDaSftK9dAtVOzctRq/cfv
GMZLKn/kqL666IKxo7jeDrTiYVXJ50NQHr0Je0t8NBCX6uBq3p6McJdBbRwOsSbg
lt0AwJ5krrzQX1U46R2ntrwkm2JvtP0ZPCrFqd8157dqkiJFafewGIBF5n10C3KH
5InfdXkwHGRJ8OcysoSh0OMVKVOTZavhOYjku8fX/YEnxf3wR39PMhSWb5k11rZT
BZdNlOa3wT8AHCrIQiEDJJn3DGeYoXtG6HIuPX68TPew7IO55+sPSxFHBAQXLAcv
gQUQoNyblXkgwkt1t8U8N1ueshXHJ1vnokB7QJzJ6SObG/qlI6TXlq5jfKlOsydV
SAbioV2rFh18rvlhAxvevO9+oZSXf3dsXDX9L4VCVK/LDaYQlNUXglLRILPUEW50
/pFbJVliMtdsZHOBWlx8K/xAihf6XjWkjeAB9mlxuiCmVHESZuSah8u+W3qLKky4
sFiqcuJ/Ta+hnthGTF1sJwWfp5AyefJ7dFYoq341kFeW4dZhbWgoQf96qZade9/W
ZklH5uoGqcs3TrMQ+dUP3MTyvdPq7UUoPeeuJAe4F8eVrryPMDwaHsN2aGsF8ER3
dBmqJrLqRx07wVhV312uM6SzqM86Q+Jfw1zqMIlJKe9h5fTYFUT7pZLY0DkXAdd9
riqtbzhiSJM6xB8GKaj6K/81hWUw3ONPqdhab4Y8b4JMzORvSAZ/+CdoOjXJ4mLM
RuCjPc7eO2cCjvDtJt9afecZ+1TUYpKNNMlVI9UdL/u0kY3PzNC0Wno8uziYG9R4
8lt1ZHYvxgofRwujLYbDUjW/+Nw/g7aLwzhKp7YILRM1ZDgvdGyp2bpMohTxjsq0
42SMImoQLdjoAYY2efrVa0NAXxFSDrQN4ehFZFlei2ITdG8v6CwxARCv5VkGDaI3
yiG1fHUVaxSCzlxrwwUR9Gg2a0hoC0VDW7orr/AHFxUm4iA5+yCjlysnDLr8YTJd
a+5kaEyjRILzCkKOQdcmoj6LOgvWbLjdTl+tVsAjIKA0dJQrtuvmLdhCcojSvIcT
FH8EjtwY1SZVNcQ69XbMtaAvGlrLp3k8EsOv0yrsW3MQUzJRROKRGCr/QSOa9YRY
HFnZ+AihS0OmekX4WQuy1zoxRWGL3JnPwtzYi/bZv9COVAp5XZtEOERCM9XwS3nt
hvISfGriMdm0Ep5kcZG2dntuO4SoVrYnsrPysia7I/jnKIL/JxPEIizhTgs7KkGZ
PHvrvUwQ9ubge8ncUWqPpcWp7XUNNpbwpkXFGFZetWLeUOgdvlFN5mvtPsaarVpd
jGGspq/w5EKNPf4hwz8JqCgnoNHhIOCP2nErq6EXLfXKwBwEo4Vt1ESPfWwE8IZz
o3+/vF8A/xaT/6V7OaW7CJz5bIUuFNLhVxE2ISqVJ4NUwCmbPSgNN1BaAyFau5Ho
oGx6EXh4cb13ohMHX6sKE9JuKiQrKqf+28EoeeyrSsDrYG1KC6RKzOKTGuixLlSR
pChoLT+joRjMDAZ1c0P2zagA4zcf5NgD+A2MhnfQX+Pko16veTiwgciNi9g0MgjJ
mjDDsFqQKVBi967J+rPrEoFCSDYUih9o2d4VtPDJbvMjFtm3jstQznLrj39wV7v7
C19Gv3WnOiwfqxMfXJUVJ7u7Soc7dxJuc1MBYId2JPmhvwCJYbqz5buC7blftSUB
1YhxUxf30Gk7YBas0WvfJwRtzv+EDJFjKOat2chq6ZxZtEcYGD6Hf9NW2TMlkBUH
Z+uffwdiwq41XeHL4ANsz8WyEnY9Ck7JsT0a70YoAQnKZfGsR7aeqvugze7u7FZ0
a9LMMEo8fw9R1FPSQB2C0bCzTtFztpo9+6udG71NkRG3eS/TfmEO8HTdaKpraNJ5
4n0eN/1bSlDMb6bjUbSxVetpgSdwN1bVNhN0pPDICHfZw/2P6o3y6WSfu1Ezt8i/
krN4fsXNwg4NN5H44Js2/2xiJv1J69kWxdLRiuWCYiJ2lUxrLyTmMiR0llVGqkUy
OajHOb7YRzOEroszqpxHGd8AoTOojS6aDzvebfFcw1UlTteQiJTfoOk9zAxQTglI
i77IxJQkNQoAS0GepRKYcMlG7px3qTD76QSIK6DKLj7Q0Oba6F/LWPrjc9UazVDE
gVSMYAa6bop1xmJmzX7SsnW3kIDfx6bboxhiPXw3UJsQt1X3lam7rZtucJ4fanH4
3hY069tat8Zfgavr9p+x6150DDBJSfd+RSBpP6rvStiqxYPElA/mkobLUvM5HLi7
nj+MufTV4vY5S4TDZXRgMaYcCOfM1uY/95ESMo9nTQ9ddJvwFWDQtkDI0tIWUETg
TdXNby1sCDM4fW/pGqeo37n8jK3cTXJ5x18yERLB4nj6c8fksuXY+cfFYrAg0WqM
3aRdNM51X8POeu4Fcwip3pskH4AI1ltjXUyRWHpN9GfUv9pHjsmc90k9VJra6pMW
R7B8fWgjf0DgXL4Yt2vxjmv9cPbP8GnOWRRPRw5jqio3XtJOyKMEyKLGDEm8Il/2
SW/DmrdVyo1USvKMKwqrOU6sUZGcxBPxcLG2vSzC2SpQFW5X+gx3uRdCtXlBcsAx
HAHoqVQH8LqPdqeVm+TuSccF4lcHvgm1WGxdlmVg9RN6Ts0AbUcFo0pvilmpemA2
ARFjnXjoaidrkUyBb81c/oP85UVd7JBkwsc8eGjaCFXW6XCFeZisc+8cB7a5Ygur
kdGbVwHVvVkRMuK0mB25Qxf5MhnY7nDxh2BTqnPOgBGCU+3OzUB15tOEGs8oaeWF
dhCoCllIslp0CN9oR0VTUgtyuCZZ45Olkri7RHE9k8gFplqEUpVhrXuMGTwAGqnB
JV/e9yPEaolaDqyLEBgk4PRGs1pqGC/cFZd8WG2COlT7LPnmvqvG2ZLR7T/0XLte
DZMoseUNHJnValP5+iWeUttLOS+tsP2L/QWUNSgMMFnWL3DHETUBfYb32y0CUl0F
CEaCfrTlfafgdYxjmfxgWZm3UkZlBTVTEQ0+RF1iEd0bOqK+GgXQbISDEKzB6z6g
lYFUtvgJ4p8NVEMuc3J6BnF9WhYu+i0U+fUgGDJsWw51ntrQZ2OS2vszBwlZOWgN
b5NmbNHVYYQoglYnoG8ivrmuAK8kJIlyhvxSPZE5wNplBMbPArVbihJHn6Ehkllk
rQgCu1wX+aV/1NfFLqsKqUR3ICFinBvVuyzdbcF2o0xgYtpXzGt4jGxWTAYKk4V5
TxYwtL+5hpG6jrqYrY3C6UZCnJlS+bzCyYdD13I8b5UK8GKygqtFul8fewwJBU5R
IjsRqUZJ+uKvjyySqUcKQgR1xIMsscgSgp/rl2VlwuubWpAiOUWEarBv1rn+GIUq
h59z7v70VH5iO9zHUzrEUoOdaICBGzc/V7t687Uhg0iqeLL4Gjvor9oX2nVp8l5B
885rTBMafKunW1SDioM5/7GymX/LC/AI7ZM28c6O/iJJv8ItGqRdf01MsURGzJFb
YqX+7tkG/nf2+6eDHmypDevptIDN9X2QB1Gtf/8Ix9SZ7dJk8qF0CRlDJQ85uzlI
F6wly8/4bRrWam2YWCPwEuEOc5Njk+yjyt26vAhKddQZZQis6GoucCrtfjfTLYJC
AoEX3zIFiC/CLjZXiJWZKAlwQ9vSUv2Ns7mnCt+z1UH6E93GJ68cMVwMzbvl837R
MUAwMzbBZJ3bwZVmn4TB5xYzfV2CzsgS7Gzbt99RaL5dVpWBAhkTn7uL+fEVKh4L
e/ggsBlEcEZlecwSrWlNg7iODuNifq0owLp9yHkhvOPgV3FcxQq1MmcxdHIZOJds
T4LN8p/FMTxMfo7qNw1osdmiskPSvM+spvw0/mlA/dR0FrhOan4x9v1CBKLLsC0r
sw+ee7C0mmVZASUpMLE26guvEqbqgltG2Jcv7kYEfh01+QlXEpsnMHcGKBRL3932
uJeKvaKm1iRkDtaHTrf4QEew4H1Dj+THxF8kq2JpZfWiKLFOoyxIZDxIlt1i4ci9
9Z9aWSWpSnc0QruY4UlsoezcBl6mIPm6HarlbnlFjAnXP3eH8tLPELCRmXCBccDG
0gKic9tFbtWKdxMl32sqV0jHJ51hYGvlJ3J3pY8WS04ibTd5F6Aw4WZZZZ7ahr0M
zSfXpgawGi93kjD+EV2PVJi4R2JZwTMMwocU+ntdZRNs456mVXPGdoC3LDeZNCZi
Wo32rP8+k8bGlewuCwJYWMii6RoGHwTN9fbxc9z9ZwvukSjtz/PCY0GqjhjzgOq+
c9S0ci079dV+qtLNyLpwtriN1Wc/L+xAFFLzOgbCMOTQhSsNVq5q06vur2m6WYur
ROFrvqfMLgyb8jGVjLD9WbY2c/NHTQI04vEuju6zXKrw85c8NH2SS0tqw+hYIBkn
9uuF3RYX+LELxzkO4tdVBTMXFLVYIf0XzYRMOzy9GUnyMh6czZHu4haYyqJbpzlX
H8MDga/Kwv5SioUe6OTTAwmzQbxnGaUCpqJzKzEKzpybuvd2LPjuwwS4ojshK0xd
llPYhWAJ9woznxH5OYENMRjdmJPhoO8QnTuptnx2xWlT48W4dgiSpLkX/K8OHh5a
O9poTw/Uw2p6Q+LjZNEmq8qgColg5CNjBlGr4/pjzUo2OynUzzB4KNpvZD6iTr70
wDgAGtWAuXPfiI8EXnY1puQk28Wne6cWZt9gcS5nVqtPfzcvOvUe0rGs0FXHbcff
CTBn/nOlf7ZfJUXMvQh8XQTSW6VnFrrS21tLcUyrqUTmuA5h4Hr160UfA4zjrSOS
uDqAtPtSJNPz71zNh3wjCWD56lpqEJ9TLBANswIn7mB0d9F1R9UNmFbZ+zD6LnI8
c5+KI4aEjA/DITjiB2bXZ5KEN82Ui2CbG5eyekY5Jkt+W4KvO5qynIw3jkBwhdnO
IY27iRh2sPsAeFQiTKV5YMjT2bZz3emvwlaPcZM2g6MmBCsBxL7exHA8ULoSkSPv
I/OkarH7lRXDKqn6ZKjN3VaXrmgbpLOzUXIfLaVVJ7aaorBx8Ebs18OJBXfYde3g
F/+RuKh2jPRT/zcumse4PqVeW8QLM6h3Fq+qoWdj7QWRr8s+7PSfK2XbiRcGREoI
pV1jF/NhyS7o2dzVqf/P0OrtAcx0Y7mTAuI1hgcjpofSE6woMfOl2QKSPmsIBjC2
npkXGvaxN5k8o//SJ0HqkjY4tyI/lWM6vVd0wuhMfjRnMx0Yg8fWElWOXtMaQQM7
Efjb34zhyXVP7Xsx1ccBOF3OPMgYaCvx9MTlgfowjWAtCrFCWL9qJdtL1DOo+pob
hjC++FOoEyq/vZJ2TCZH9UPJ9QNMYiV1uCc2cyrPL+F0DvVOjJ2Knp2bMwN9cMKq
2xvZ0oIwM0dqvQspTNqT4lacFTn7/lyAvCjaJzPesQpAPcUE5S7CN0DhM35zIRK9
mbkunPKbfVu3NPLsocgoT6bcugUW04jlF4GmVXqijKvYSC0YJkcHtynQ8ZNcBO9Y
Jh1wCIbpR91SNhyVNCiQ1f6x4X4LxGa6cJ1M7tp6Rh7zIg5G7dA+8K7GdBQ6zdrs
jp+iXrMR20DXgewSRF3WbHo4ylvVoGUgW+yL4fVl2rDSadPFCEtBpPcKcvZ2TymT
jEfczDVLRrgvO8Y+KUr4uE6NU/D7DteYypx7ONG0qw2IUs/QP3uoPoVzLsnKTjD/
mmuMr1S5hZGcsHX16ZzI6YEf/GgXKbEPNwruq8vi8CTa8T5x8FSgGsNUc26Oa1gR
3YIRWEuDFxqYEAwMSk1LviSOMT8DIBRg8uS7sE/SJ6/prlio8NiXOTpQlpSH8VKb
sbrC2jvzZidSIe6I61e7FkcNZ0ZQp6Zj6opS4G9gnHeJNgu0hoxm7hPb42aTQqpz
8uQ9tDWeJzNiyhr88Yz3Zl2m929Z+F+2bjfNT/RGuYOkaMQroRvPuH+h5OROVOWI
9ujOBkYsd1TNzr8ictiy8arANz2zITKHrDdpqT8FMoAaL1afaoD6f9p98oGnkoZx
hsgrfiGdyWUahkznj1BtaPrBXyt+CUh/mFz0IWmLq3vF1PBVZ7dIgIi3/Ywu8VKg
HCGhfdKfknU8AVopEARw5EReVGh5lsmN5VTsXi/taRcgnYNbjHRhpxvulV9mcLbh
/OsBKcpl1479Pce34k1F7CUuHGDEBKoXgi/3JOcNLDFf837sql4uiHNwPhN3iTKF
mGKSp/KyDeoqmdaFR90T11A1mZlCVA5KkGn7ozDOzHdDMHKlaUvMQzEZsBe6UHzL
8DhHjL3v895PnfPB1HjBk94L0BE4Kc/yd11y8Z71S61PEyMILXJ3nGVdFpCqaIlA
tJvxhKz6JGHZVL6z5TykTb56L7uTagY1Xx6UZpvny2VYZce0IoH1r3qnHEVM7VWM
NOJpQCiDyBI6wVdMy5rnAaYICBZaHyE7jtYw3NVLwnAxuYA00olradeDJPyI/zfK
RRsX8KUokEl7aKmIK7z4Js6g/PnWkIa9fFXAQFOZ5o+zHPBN/uuSdrThppzUSwDf
9F2nUg068PT8StLRFD3TikAhLwLWBdz0uAyPX+LmpBr4S7TZbewp6TGqSimtimcu
pDcxTihJYyx23dEHoCAOd/HCoDX8Hk1lu/SV4gRZ1wPeM0Kl2XCZjNLmwB65J1ql
oc34q0TB7UlxmFyQHtmuQ+z4EjElNb/9kMq9NwzBiIcDA70MxuENEJ3rymIXtfZG
vJz6kg4KIz1vHHkbbZKQ9NVR2bDzOCrLvh2U4PPN6lJtDBOlLxoWriBNRKyroWBE
+RCD9OE3J/mRkK0wNq5QfcpYT0YOo7y2L4HC0q0esddoXdcIafVN8Oh63VfhepZ0
6bjuxZDBZtY7zhqPBvOZTtdU/Bg1kaUWnnlqAvb255icGpaltZNxURPM1OH0IUSe
6jwyKZkoTQjQv8pAZ3cHjTsKziMCW7/KkAUDlT1p1sT0BNxaeRSf2KWfIx1fqUdp
CY/ii1XEWm8yhRa0tFV4bwfOtQtGXam04h3ckMOOplf8dI9CtSoa0x/Vv/THfXvd
SUI9DvsDvpAUXS8i79uGDHana+zJZVNxAKEyqLyzw9jftLIycM8mEamJTmMTTrY2
lh557YrXSlgPPMdR5qtN46iJY/jRujgdbzQzDFiGcG+/H+m2SzH2Oz5JmAdwPgIZ
Q17JcdMuswgGU9OziF0osXWIP1EWkwd2Y+BW7pO0waNWRQvI0oHr50w9KKzRPuce
0OHPlksxw2JdPdhTczlnR04Q7l9IBWSfkdZ3nciZn53yc874a3Sfm8ZBmeOcyM/b
d65CBgCQLsLXt8XiLpuR5uVNnN/Mg6xBXCODcT3J2h6I106h5vBSOlUHkJdPjfmC
bwTspwlAIU10f1Kw8PQ2p9YVu+b7ahoOvfxu/bk5Qi9whEQ8BFkYq/PrwN0mfWKz
Ola6+pfy1mYVZDEYDxhqvfHJYS7GdAfvv8hWNs71T6JZyzmDZ1Wn/MfGCrN3eobg
Xsl/1dvN5Zp0+YHFikUUoiM3S1SzmDX21bU9meyfORhihbqJ+eOYHEDazt91aM9H
HFMd82b7NbnMjQWb/f/JJ/Aczp7M8z2qIzP5rApiYjGSOHAFMr5lxfNi1qK7RgC2
NNl2oBS2WDi3XLs4zo4SJ3kpfHCAWFvZFFaYOjkDJQGtkHQdnTAq7ralizvFIRQl
smPN9U1fBFhzXY4Gxb0TRElMg93ulAs+6Ej76YXFB6FCfb+vrkwcygaasD5PAiEj
fWinlKh3VZvPARPYwHp8Vu2L2h6sIxM4eEdPyfLNPZS0BjbeqZUV/QcV1yJcwrDQ
JJhNxkotL917Rxq5cPbVgj5LPo1xWhtRyNP1kNOtW/QwuCWmYNqkSfC9yQ72VvVC
CGqFAllgq1mia7i9U0xN6L5np161A9wSlbHHmgIwYJsb1Pj8IDF5eHwzKse6wfn6
cWr0MyEqPJ2JV+aPwgZ+qEXTixZx6nTrGzKNdl0ORVnbP3eVUIyO1Isthu0xSFim
GWgzO6Jdj/rEBEZiHCzvtOQypD9Y02HzEg1nqCcKWvpiIzpAIcsFH6HxSPO6WMU0
oUn3d0kcBub33d59q1B2AFwaqaTkRE1ghkKi/smoJ4SiM+TXSrP7ramwme54mMQV
KKsSjKoouLLZ8FEe1TC4mpyI9w1mDjsGE/6bR4iZdsOPiDyj4Lq+JVjJyjmw1puZ
bOGqIBRhwboXrEb9zazq3MIHo3TBAdgDwKKykxLF+ij3Fl/TNeP2X64qhvkBhYyK
gq/iq7B72tdRvWqRrTn9jGjHOi6tBPqGSGTu9s38tJsiTKTcgQkquDgK3JxZq5dd
WdA3SzlJU/6poGRvZOH3owLafzDDD9nPWxPXYGRoMuxx39/5G6En2v+Is+hVsxWk
EoriA4hz3rMNTj0DbLj2j+obLW0v2WgvRaX+zLo4R1jptPgtvKDIeNbPab8/55Be
171yhmXZh8bZBCY2Z0x/0yYbVHfxzeuhPadHqITA72X0exRzLc2ZSLJu9Hr0Axfb
SFLliIsKaEot8BdTuFCFY8NZQKtuOrEgNR4A0ruSxUcrX9LVCFNZlWx1aY69zc+8
Qs90BlHB42BJxi8OUHcXshrBHmirhqsULEqJxqBc6zS9rKZupp5qRK8ok8H2ZXVz
8MLFpcVnrsC8qQPuI6hz+gUDmITTW3rTkbgw+8h6pXfHvZH0TXddPGgERqw3UACH
WlUBVIGNZo9BCJJkwf7pdKM0HDkNwH306GrNNjjjGYOM2qOCIx1t1IXsgiKicp1A
oCxrILvazgxZeQ8lLtlqn0kC56n6G7t6JX7gpgfsQcJRtQo4dGKa/sfhAIR0eU7y
SRNwKCjO7M2gJ6dNhzH7FOtClLH95/UiZLjDfZpZajm6jqwEa8b1SqkpYj1Smixx
PBPLESLfsh6HzFHrySF8cNF9OhtPioXpzxLQXQJ1ak8yx20RXAZawmmagEyeBUaW
jFCYgunCMKkb5J7VpXgylqkgKEeREV5bvCz3pnxA/WG8aAttLy8NKIJ48WzfLv/w
vltAgFvn4UwhPYT98f3GMgShY7YUUwUx/Hk3xwBUawSOT6nSX7ue+G97xex8f6lE
IDcZ6TcnnMxirnX9Ix1loc9ZC8BypjQ9fK+DIdyE1SsNJeVz3upEJHtPWQLmPF4U
hcX7MowIgeHH4uGzhZG+aWtSO73Zi8OhwRys4lW0itDr2X6uA86VFSZrQqDii5x/
1UJ+GSqfd+8oy7VAbyXfyfmcenDaSbKZqoXoPHnfiGlxTOjy979InL2+00JzAYTb
Sr4hI5xV5LTU2K3cgjPBy1P39B4ad+Yl1QMqGwrG87MpbV1lwLEnE0zPyTAcjdd5
msz21+eP7oulNIn+VVG6v56pxddWUb5Uzq+wLVT6r3si0gwPct/jAvqeIkC3zOSL
zcQKODHIvMHg2dygnMTKQQHNyR3y1Qx4C9Iv+oXZkvPeT25ANnoLTua4gif5zmib
Ws24FystED9zbxYrZ9XIn8spbmdXjZftImIsM+oERMx/HmHZbAPmlCJHohMWiUMf
w8Q1jiwroyf30/IscgnfR6PMgbj/A0kl/MxN0j3v504GuE5N8BTsyyO7UeyAIPcf
LfW54YXwVL4E4XR5FRxDYYeven+2nMYhM+f6m3bhq4XFiRL4GcJgt55LnjyoRiye
JJ74pT4SP7vM81k7AK6wrxRMF9GrhP4Bhrhhb3ZebiDlnF4vUlP9gsmDSuu7d06w
hVXPWBREDGjfYJDCZuhUN+62u4bSVwQHW/PWH8hLTM5X4pvWmAQznkglOhMn6qsH
ysNs83IqcpOQWBE4cgidujS/bsQvxWjPi4jJAbhbt0J9eH9wIj8ci2wL3zg9B2TA
B2DPiaHZZHwEmdwUD9ol9hpegJwe+tOZ0GswlvQRSv4cG4HmZ6ioEHOCtCIBH+Wm
ukM2C1LYr08k7Zt8Ii8hHsOmcohcfLrGyE7LaIbFSaj2hvBklFLxOYlSztEq5l8j
TtwaZky47XYmDH1b6qgsLKAur1zbk6o6l2s3Fbm6D0E6ev8KZu2Hape52rSNMM5V
xgTBoAHOeeHM+xlhvbyoYafqzu60UEpkhmgR1sZjPLw06FXydBbrBV40lK+pmYMb
2tYmRuJk2wOfp/B6EY07sses1ljJg94Od8GXpEwkk2jBeOb2XMavYdNJ47zSIapM
sM3xob5xNX1S62WPZZ86ZMxxCcsXEadtq0knem5NMB/ThBwm0XY0xaCTQ3eFlC5e
W05i3j11aNt3/rMhyfkwc5OwIsSnr1dKP1I4HgEVD1yZSFQQtsb/AWRvDMH2B6Qo
8JLwjlUB1ZCzrQ7nmzKdQplPgojIz7rN69NTM7kKc0KcbQ0Hpaqk4z3nicV0CT+/
CNOreAfcM02uCf8EsVPINk+yxzoTZCcawZuCqfB14GGsStWmIm2WOtyaVi4K9xqt
DwjyqeYpu7IHPq5oqbVQDBN4U3fkhSoqzDyeONwHWNk3t2KF4ehUNxkbC2BkN1Nm
Q9GspenBxTXgVmmkXmrqbjqJjMjwUuZcLUPsylF5N7RjrfxDl/4wI8WCqlK805O2
l4EAMznj8lh1c0PCoQoANUEZVzrh381TlLH/W+2p3YyMrv49jY0DrALfl46QddOH
EGX6dW1palfGbKRF2vmxh/AXojlUN92YtW66Yntvyt1D4g/k34WYSc6L86Y7HClL
qFTQuoDrblL0UP5i6BrBFAJL/74A8ze8Q2LgtO3jmVim+7/OS09RaQYszq6BM1BE
YHu/BIU+YBdxN1/S6Yr7KtSEDk+yWB4k3NTS1DRkbZJ/qu907BGS7jqRfvNhTXDp
kzBq5Ov7OVtZ0s60a2rdJd6BOXb/9B7CJqW3NY2dxzqXmdS45rvcuJl9wtOo/z43
0KA5eTwJe1490dFoLg3Vw6SerQjDfoyMVu9NpLBv6CVYt48f5kU7oj5SE3vpc+Gh
p7owQOGGT9DjNRq6oO/6izyDMTxC2Zt5WmpKPiUHdSaSLaP/I1tSfppC9FLbgWUg
6QnIk4ghCxVQCUZQTFgFGpTx/fRMIL9YrmZ+Qge5+2+VJHAPSGWQTNjlpgvbt9WD
elrmQ4GRWMUZiKIu20U8g/HEiV37CbuFrhJGqMYr2+QzqczazwZLjstLOXX3Z0cH
sNfrouQF7/1ZvgQfLkrCVb3EXRMdbt9dWL7XwcVkDcy2rPeqhSkoee6V4TFhe1Lk
fDd57FtiTe44LA9PfvEZucKw85vY3iJ7vuVuyNGh/2ve7DJ8J78amihDUB+7s9If
L8pEwQlA8M/kZeHPG2hgWqU02qdZMiHJjedJxpaAdpCkJfmUCXPDRLfE9DeX/24q
zrZCE0PbEepT9JoPiJloTTNVALBPOWJ+gt2ysuf9/L+5UofAc4v6MJk7ssg9jHCH
NPAoSb/PWeHeT+3A7HinAxPBeiUnwXXVXRhKCwrO+UiJrmDUhDW8DKEZhdb0vE2A
sUi5C/6iX5/YRce94kKbPNnRkqhUuHD1V+JEHIC0Lf8bnmQ5Rwj+KO/3FNKmO0fH
51n8qoFqqPC0MNSwfCpFbZXZ0yj/UyaAaaQR1YJykVnsM9oEWaraF74cTv/AJOzY
tSO4P0YYE1q0uOf//bPKjLCT+hLIhDPQ8EGpGwYQD2FGZBzurUKD8sMK9lvQRLU2
tCaiwsqvHaIPIZzpTu4xDJ/zWAkJozZ+NUFbB64wEsBe7O2x8d10YeDePX0KQEWv
UvQZnyB1YCJE18XsuEpf9XAPhbLjNGHwX4YUHHiQHXI0MwTW+cUXJBRXY458lkBQ
0FEqnGM8NsUz0/t2MWObdCs+YgiZaDbBB3J+JXMyrU8/UxZRD3YEo8sZzVNdArCc
0Exg9R3K3jEIixK/vXnFoQdBmtj56eX+oHTv78ze+xo87GcNb053Re9bGrzJyEZ+
GbrQuo5g1xYIqFmuhWGXN/WQBcsO7WWq7bZNuEmkI7OU573DMVJFxhcNIxE6S1+V
DiObNy+ZuxPuFJ8JjKIwgBqwOUlKPbk2Z9tbI38NJWlc71x94SI+zc3ZbgagWMoZ
078sj8EnXjj5lbTFgAmKz2E3qxZL8u91lDbWsW1825+Kx9tQh97glrkqUTvwkBRo
f08igvPe2dcpOvY2UKRgz15ysO4lJTaqMIGraiFBcBEbZ4b1XclKW3SCKNlqWm+h
T5KfnYxeSZg6czCshTScwUeRcm+1eNfJkYQgh3DChepFCrdCtKgzMDPEXqplBC1O
gp0Lyg7IVAdcFxA9GrBEUlswYjUkt0cwpOr+FMr8eB6xziSrLKJABq0t5ExfYzSB
r90PdLhccP96fFZPcWqmbf0HCSniKWy4oCZqs/tFeFYtOrBsDIEsX6ZsfcEk8Frp
RF3g0DPJLd3O/m9ZqfxINC8pOYk3lIJrtdxGGLgF+XgyeJpihLvIGqdwJ7NDsx5b
cTtCjNMjwfBDATandYEXF9gx/r9/skbf/ipikehuLJ5XXFM+AWUKM9XnbQem35Od
96yrYYWjZvMJnEOWCajb9kN45j9SCqNNzMtVDsJn2l6iUezZChu6JF+4NY4EQ39C
CrvrIHaBWflVcjwlbMcWCI8x4CLdy6zTCYj3Eu97gpg/0+Qv17okUyo+I/8mJyAO
8+7BT5BCGntNhY0Ha9Qru8kZQ4WccKA15qWZZjQSiF0AlV6fbgDpJgnuLnL/k0kw
zz2bR1HxaWi9aQLiAuAhWX5im43SRfnPkB9DI9OXyFGSaDiKJ2Chl5BW5oGjmQhy
hvMmR1voGvYWsFUxqibrXCbjzhFYqkku8Wr3xbF3BVbI0EkhUIKJwW2dLLjEwHi6
bkf7gSv0CBkoxr/jJFpWmQ43jos80ZdpfL2N9A/Y037hwlm63MR4zfxjFDTWUFZg
gwn4jTL5mA/SA8vq9nBakZi2rFTZcjCFV0KTkbz4pIN4g7fep+eLmdC1cEtb8BqG
0IlertmVfzjXb/C+wiaaG4XgSTBmo+2hglGjL36TrTYWq6QmEgdbmMfZRnkUh5QJ
dvs+d0CwQz3kkY+0AuLLKoRKSkXA8BdEs34xQ209xjie3N2qhSFb4MXNfKYOPYrq
tR2n1ZhvfwvlmG+nklCoPz/F0aSNzRK8d7Xy1lYxaP0HdsSVq3iw29xKRABzu25C
ysLkZjShCJT14+8d4mWa0GzPn6E03clNsAhH5QmdVy9P3MsjuWWbx7I7cklc7IJ2
B/JRbeOrhhAWCickoFngKiTGSPK3pOnljXTrbAmWKHou5af6PcP4zfnuaZeMXcX7
bHWi5nOAZMGv1drQYAKKbEn+NM5beUE9Rh7oPlhbOyIfsu8KttoG81BG8FuW2K0C
k7w0el0zVoHLNjYzglq9jdAvWxsFosarkm0kiqMQ3hi4oXOGrsyreKRxb/OEuEgo
bwLuON8dzn9ng3Jy/JaRYJBhaddbb8mJLFQHtcPaxQJPQWI8OClDGmKfAGxqSM0y
a1hUtbtmnyrYntwTdmwowOzWEzQ8CiBdE9rBapB7UPIkWO73keiNofNHmXWX5KW6
d5TGFOC6LEV5FKaTqPdt/sMOWTpYz+pY3AgNR3+QWiyTpZCiNrlIrVKvT+ZvJZGs
YeTh2x+i94qKrQpSNjRkjLF8yMSqi413ct/WYsBH1TgAG+Lvc67mt2v5m/JnSCcc
O0/GIZrYzwe9Qui7cLKmbc7cdpTljS4kvLRs3XHJsQhPaDeX5rjaIaedcTRXRDi1
ft9k8gj2+lx/kIRQ7+RxL5U8shvVIXjj85Eu+BSZ8ZFSglUW7ZNG5WBSB6ekhdpI
iVeet4sJfUeHgzf2N9ZLSwKf1wVmtluRfBPPBPiW1a+WHrQuJgNj38KFoBi6vFbF
cmOWa8DgCtF9T6mcNTiFKa5pGPfEyWUh7Esy3liHb/HiAaMTGCtZdfzHXH8Xnnaf
eHrENhUukDCzlii5gb/0AjGAC2rz0YzlttCQuK4nz6Ck96vN41nrHiLRp8zURoxx
Mrgfq3U3jpRLCwM3ouKZMsFS6o7T3TANz6o/6h+CAjUGFbgeALz77uwr3ftoaDuV
PjfcH+Z+m9fymfaicP8OjWh7mcxKijsMNXxX77qzeKCa+x05Dv55C5+0w8YKHXgY
r6xJcbRYzgc2RvtD5kEKvG4xC/NVzEDMiXvFIf8DusKuaZ/b2sfO5xcvH8z6pIzN
M5P6bpvbAwsrG/BEU29BzSW+f8SjM4Iig45SM3S6pjl9DwO4xk5kmG8gbzQ6q3Jm
ptHY3QngAsx0CkHia3yO7wNxr+4nmICWM1FmCDte85JHuedcNcNIgzZt6XMFj1/H
9bBlklhHa0fTAFZFU2GLjXL9jMGN282MVB48TylF2hXpmyXDFdGFQ9J26BHho01W
ivBnMr9yG1/j5abzmpGI+LuscDqhEWF2/1RohhcUZpyTs9+IP9IQFYhPne+8h9Bc
p+zAbNykjbrkVbJzmpgC45YQiQqm3YWAAdbsCneWeQNDRCkKQh6oYeH6sEyVXeJb
LV7rRE2YAfkaJIBSot7ugpjcEpynjf/xBs8YtcgHU6fNdZ1Qd72y2NQ6T0IzpOsm
DI8Jm0cH4Wg5TME8agBrL6WyYKoJWHjj/pA/TuEkoO+6epgk5FWUjm0VxrQg8AFD
yhq/z/E87211ZqDwtCppGpIENG573FgY8tpFINyrqUEAksmQsh+aEqmD40Yvj2Kj
UdP6afy2L3En7RjlfUNnXfy36s4JE+qZ/+tah8EYI4lDc7CfdHxxVFRwEZKFlLQm
rOwimIoyOI6kMWwHEBx9ir+i/umfydZ+oNx2V7wcaMPh7J79/wOjpw1pjlvRjJl4
/vjHkICotRfkFBtlDaoScFU5g0kll7qqOZg+xdIPFdHhHmAjX27YrQ1TMdEZgQvA
hM4QbqlynAFrWVhNKDlZ8d/oRYM7v4IwHRp2XJdB4UiCPc+mSTD97FmBFfvW3JM0
kjWI3FIKA7BUQS21H46a3oVicxVY1elgdbP+rFUkvY8Mv7N5oIoIlbx5ksGCEAK8
T5B1zq1PYYPqlcNJ6Jy05oWHFJkfFiuTijwN82dRnZEJzLRiXnepj14H3EuuigjK
bxYihzq6TJKc6ulom+6pS8t06Y6kz/4jupjmB7gQ9WczGvurzQEqd9NP6Pkp84fW
M+kjKIbJaK6isyZcpnA5t/D7PFNlTryilNKn1a6ZU4QIPQBjVyHNt96zS3Ln5lJo
YaUX9VaW2nkqyz8HUH3SlbfyocFELL6W2FK4zsPxJoHqXzxLiawd9NYwsppqzvYJ
vL5FNSCAS6jbc2F4YiXdYYKtPv4qZYLnls4ICciV9vQBq9lWt11CRnPZVQSsMYKV
ZZJXd/U7fM3DfZNZmdf0KjU8EmFADHsgIS3n/PxQ8JKPOC4vCe/Ug4bo+X1uibp1
U+RdLfGuw5vhTBmHOOTGSYASMt8HKvPH+eY3a34WJq3WPnifzx+JII4gydKQLAta
U4hcRqo1IBddST1h0HUevjecHhCi/tGVG5Lq4KX9ufwWjFdsvZ9qPNEh9UpXjQ4M
4OqQgBokPwW2o5NG0U3JTe0G8NMzjnxpWtTv/YmfwbUkGlPYvckfqinihsUo7M25
zUS3wfiKmeF/8ZvjFgLFZjEsYcEFlrVG1YpoeF3PCe8NppklIbUEltW1XwCdZuvH
CaRONoFAtQ5Jlg75arorBGmXXC2g3nuR0sFeiWG627VHuZpBFbTXtAJzHQ8gmc2v
8B2so6EvAmtKYEwaUcgReJOHzuJ5YZ9KRlFxCIPfpykwrDv8mMAYnegTzNYlS5aM
vnGSzBFqNGcTQw67dPpv6NjBl82ljQX9QDtBFitmgRddorDytimn4BQRP2iKeKER
YWwCN7RIAipMvFKHXehntw2tpQ0WRjF3+wWEg3YwBH8unV60kvM2j0BC14uU/Ymo
IhGqQ1JLFFaWoJKVaBM3aC8lfJChhQje0b3YTMiizqkhtejsE2QXvmg6HoXqqCqs
fwmMZj8+nXphUxa2XkfRN91SxH3tvwzc9uejjt9DWasBMxluTr5MaTGUPP5EG9s2
PnKsAHsW4Q9voo8umomWTHz79yiwNZgj7scgxC1F9EZ/3rSSfn6soTBnY8fRrN8h
p0UY8nOv5wNd9ws5weu+9Pb6JAbsZ/cFZKOKlT9+UKh8w74XoyQYsm8ilYDAYn6r
Jx/nThG63arx5krPumisYupxCOfvA1mgHmC/PiW4tJKWgkteGN+CVE5qWItsu3r9
L7Drrd2HBUS4Rqee/cc6TACjW/QgulmtKt43bALHWrzdupmlkIhFRI7LT2/IstQz
xptQmpf+7x2hhnOjlv4VS73+yoQiKiE+27swvY86mkNUUZP9ElC2fJ0S2o/BEGvt
A8doVtT+Rd3qOvVYXbUo1E47ZF/Svbv3D3nr1cP+5hZXzltmLJDg6RxSCJPDYW/p
gBe3JxVw5zshsuedi+o2hTXVLZIqUbUdj22AXjGEIqDbBHbg4wanPYsOj4Rsct8z
zC8ajQ1+hrhBsH+Lp9gt1rW6w1uFtd+aPeRw16zt+AnUuK6hDsg2Gg1hw5RA4sJB
lyz6UpMLOcRaZkRbceQlTYuYNfuzKtwbTpDVnLrCzWiq5ju8WAzZTHzRihOsY7jh
qJCGnRZdl705QjZFWlEsRu9yHYrWikcSB3oEo5C1Q9rIDWw2aWpwQlur/BTVdiqk
WrI8jBYbEzULv2gRBGcb5FEzjUAxvl0ALzQfrkoc6NGyixaTA8b4sNN/0FFInAeu
nQWWpHoSptrg7Z+71gmt3j+7WRs+ueB62Lt1HoUFniFfjA60ltlPbYoTyzFQ8I+K
VaPX8r6aW5BpE4KcourNBPL5vbcZkzQxJM634yeDM2zWS/U+q7rMrjdi7R/qCaBQ
4NcMpM5JjUi9eJx2HanaT1Nnh1MbJweBzHEFYLfeZJWAAvzuLLjhkmCpkiELvuaU
QizzFWG4a2hlp812lZgP8Ovaxt1EVpkfYe6pBLMNqSflAsYvAlBzyVP8xhOijuTJ
dBuQbO+WNZ1NiOuTNObtUJF496YqH1tXGZV9bBRee2zpBgBLv0hO88VmuIdLJG4q
4cgm+jDzh+KEC1cayV98Ga8nHeIw3WlR3fbYiQUMGqSa8dJtxv0rTVS9rKWw5YP3
ZpLJ6GtnWfDSzqtcEuwDKTWgmHXoqDSLQXddhcQNWgVCZ0OY9ZbZ4HdgVFnd3Ct0
s9c7UXM9mEeLah8Duxu8ne1olq49TAV77F568uIg0H/atsF4J8QvR1MqTe2P7Ovc
mDfpdmvap6d6f8E77jcZpdzpZp2M1ra8wDuxfzOGLG2xjtIw2hgdiHJaxLMGY1TA
Q/Qtwvx4AIlqmojBn67GgSFJu9PVY5QpJ9fExCcgIitIlyE1MJpH7nDSjBf0v58g
trNBjadsTDy43rwEN9AW91Ad6XjciMUR+5XSM4CA0/h9Uce1xD/o5PlndhfclRUT
viwCsQ/ZHi2ZagbLznLnk4qqwI1XNGp7ftp5xuXvqdc/E4Ni0pLZ5dGmtj1EH0WK
v6PnDKQzvcTBjHhbJk5+Vmq2HpgtUhNDU7A8zgCWIoOZkREA47I2NXwzpoqFbdtv
wibFGOnWB1A2GbQCQZOYC7osLUGbF++mvoDs8/MuZmydFt1wc/vHbC6Hvbu2dex3
3ZI5FvXxCf3fxeO4nRMaNlSYuaWA0eWSkhcTUwFQCGuqXKsVnjJBH4UP8rDBFUD2
GY5WTE1hOmyYflefEcCRuMy3Gm3WGLYHOpgby5B8KTTqNPMD4S4jtrJjfNnjVae/
G1cND+EEKsYxvKW1dYS6oeN4360I3VtGYP9T5ia1XDGDNpyj1dLjx5Rcl1vDLPtb
ze9PoQ7WFB5HERN6NQp8KGPZ7MCzsEJW4/yISkOzRXeNAoFf4jW08RO+wcThEn4Y
D7gmhjkZ2e9c8Jznny2ACgCZ47OJoQZ98J1w9I04Y0NrdlFBnU48aYu8Iq06AW0v
B5PW0IMSYmrQFTMjW01h+wBuQCvS78qD4CZKddsJT10Zp/6/xDMZ1gxrHMKvDJ9g
SRzXY5fkF5zMi0PspJz1dZq3XE330yZLCK8FI7wDXK2cjvzovWXkLbOOi65HKJg5
p8RrB9hSOw3bMPpx6oYLasrip/iJ4h70uXqQiE0SVUTkWxIfhJEICItLtl/ktKkW
IxI0KUlY2OYkeQNqfCZf9qxLG/69LwojzZreSBMLC2r1AEPMIo4LASbyIja1QtjJ
/ZVTAx+H8jABKXmz2eihu3SHwUT8BK/1JAYTOhFm1vJTO44XXsUTyvYE+Fig62eq
08D6UqLICUal/vIC3dk990fzRofvIJeHaLpbXeK7oQJwcwaJ8SpI06UXaLoHPnex
cOLyrVLWGSdpGcEZKWdio/XvNXjpLdTFJiIME7Gj7MiTJrfES/EK2+6Q0l7IiW0T
0tpV+GF0kW8AC8iz7twPCNQZoClpQMmq0TLR71P3tAAzIHSTjv7tPqtKqxg9fu4m
9ke+oviiJpMF6lm1a/14NTSQCql0a9P+pKtmRG8q7du+xeyV0LRZ1R+LWfZPCQOb
fkMUU94gIv/LqQ/IXSuq8XK9GdyknUVjfogCvooZr2tz0Y2iIT84AZTisCOrPEJ7
8cYj38H+BYgjfmgIH/nSul3RPqwWSD06zKUrNxCvezbLIdrR0Hdq5yNP+2H2XY+I
BMJOucOJwxRUey5v4oigrfkrgrApVJyYwTETIHdDjQzjURuyg3qyxD4XyhG2ve/A
xeyl1kllUyN4gkIWMRWOBlqHp1v3F4jjZ5XTsUHTlVy+WXYKAq1UlicDxvFaQvMq
F0MqJHMHpDbY7jko5zbmhd3QsEnPxRZT/6x/9P22DuTIsTtFJHtfR004G9BUDFTn
IERV4FS5gVg6XIFuDdzZ5SIpeSxNC18UNh+W/OU4zPPWBEfCu5e89y3nABoWwzwd
QqGzLexHQpBL3QfxU5hrurQYZ5xuYAsFLG6RBemrbCb1vt/a2yo9jEA+cXBy6JPo
NTYAsFnOkbqVx7DYjJQACEkQh3XCPk/JnWUec49mAiMCyJlGh8APPKPCLRPHel4e
LPpVmIY3xq7egD31pwlfeXYOnH0gxgHwt7fctmP3hNb6nty4vsvrTkeZu97IVTCd
zcwA9Lcuyr5T4yjBQCGf+14BmOEf0pTLXktcVBJQp7pHrZJp0bf4F0Z7sU05vcMF
CDqEx/NyzbM7+qoBFXFAa4ZHV72ZDMVtKc0Nk1+Foj8Xp6hinn4BOGQDsO33kB6O
q8HF0WbcgLAc8Rf9j3PKAgw6WaAif/xLbO4ge6iij4xMjzUE0rXPwjQwgRl6YDFW
qnyR7mTnv5sKuCCXY8TX55Z0/3lIRrLqqXsCGVn1O+6p3sTo549MdOAxyac3vm5u
UKrSqjjpr3b27CfKBi+9HpVsWia2f+W0JBQwweW1qNM4vN7DXi5CRjcgYlmd0sIC
gv/RsJwAdx3trViwCogb27MeY03XSSNJ6lWhw8UPb0zVs1s1ggzVHeHPozM/ysdZ
ZqGDU/lVf9LmxfNApIkse2VHLk8W4AkKeWGxFq0U94oiEd4E/i7wpxKU8KYEd5Zz
vrlPB0hMpzS6vAG/st0Q3lITBxRtHsPL7A7CxQuD/JnTG/u0IG5S8TKlvNd0H58k
nreqGJJftOFE64ZYGv0OFzL5KTn5NGHCGgL8rTJ3Lj7FZjeWifBvjZBVY45chMLW
uqXnItLySFtFC0sSXuxQtsgMT7DAnlTWVkBF13hG/TIpWuRT7pDqNGvyDVgQMp1u
oywTuCCMshjSzEXe6wgUeDzY8Y8wDjrb5BgEKv4JRsoIIaWSWltRrByeqMmG7jFP
16LjzNaf5ijo6nNL0ee31rJr5J+Q2NYcffEGNJpkMZCjTCgTCBVHryATjK+Rowgf
yFq3dT0+Sh7iKaFs2NFOk2RaAZr1tXdmCplm8srBfHfDYDVOk+EJB74mmiqNL9QP
pBDWdo4RSPgwEnfgRGr3IuE2gGBn3MXcFntY8FICXn8QoRQkvVc1hqvtVhWkvwGb
QYNmBwpyBm/61SOohrs1qmhxugAAEy20GVR3a98+2eHa9KIlkqPbP/CsiBPjl0E8
vpJ0ngSkonQVtXbGMKBsA/ALb20WL1rFpzXkLw7vYaTWXoNbq84Vatr/a8jTnZ15
1z1W15cD7b24D02y/k3OV4yHkNz3LTOlGdoYU12RxzyGxr/FmPeiF636Z1+Zlli9
nlVVRlD+XWGTRkIOFqSvy/emvVlNkS8zhnC2sBXadqufXh48tkt9qmsfZF5OijgV
V3kAKi1Nkcrv+xbDMIiUZgOElNl+huOuI6DiebtK9oqJMU5IzkFoeKKM4KjgdlAD
O4AZUiluQBthLkZwtIlCGnWlR2TfaZ9a0/YU8ix8T7nrXB4u171syQk+JIRa+go4
BRraTle7D+t2UhrV/XdBwwXlTUevMPblAGJmKQPb6ULw0NWPOITHmXy/zmHHBq72
ChZC0QzLTt780druKFE4pqfYBbPJQCpFVBPQQ2si0oRF61VCmQZ2Tm6zVA52Q9Mx
RjKPggenyfYxWAu5CAGqx3v9WQHTPuSo7FRXY8xryJnBF0n/ualnN3XeMdY3tCkP
vsnnMJzXpI3a/2qKm0FatH1JA+8jnNRa4P8wOxFRtzLQoIsqDLG/AS/1/P2kzzvQ
yan20d06CF/ZUxtKWy2orNUBLqy6Zfj1x1JcM9vV4Eh2QFSm+Ll3DX7LcGwC6DPh
E0bHMejWzKzFRxHFJqojncB5G2FVrdhce3Fyl75DN+UGzzEg0c3oDsNdMHKBsIw4
DsajBlMgclrw/OPDLSSiRy8A8X20HS0EYkcXtJJmxAtbbGOt0LejIsswAgB9DZT+
jB7sEWeudRpV4mZ7dICN7T9R9nu49EHAx0NU/wrD4JJlFdE2tlQ5Z+Q2/rrOIUtT
pH6N/QhuGqKV6rivUqN0sHa3wqfkt8JNlROuQfMC4N4Zt4SE2/pNiwCqHPmgyMZS
yOOm2f5V8JnZWddXLFFCxHHKyIVraEzOkxL8Jjxv4tlLJ78ujajCBHZ2TdwZ7HDv
I7PkFJFqK2qbFuFa2LGm+64Vj3aWxfEMtOYBXKB+aP9mnMQuMiNVEpp3KTTO8B5S
bdMM7GGqjCMSy+ESQbEPskisrtvGR3+RrwL+SAzvKpzxco2PhUqAMLQW5wT3C1GH
48/awIa8EiPopwgXpL4IWJP5RTx7IRUGOFeBYx1IDp8ged/TkDFmD1QRLDQwZQQ9
r4Vaw6/szwuIKdO0eUrSrWJQnltNfrmCy6E/HG4dWBhf2/h6Eqweo3hE1CaY1iW4
VudfEFZEIfPEovA4Hl6/Z4BQnXI+Uja2Y994PRwgOo7P23yXY1gU9wJagHOow4tv
9NMfYMNIzhw8TpQIsaw19VbcV8pinUzbkbEZflGKa/tl4N7TVXYbmw4SfiAFhDcH
liKEYt023Cl1uzetkF0aKXBy7A+ZRu1QTuh2cMgglYkVFhbWpkw41O+ld0wl3b6X
YpsQktYAJLq6Zk2omZDZ7k4/Ji9Z/F7jErZbr2I+cmHELvz9d2KKb5NG3DW4YlLl
gRxsBxXJV8qtnOF3Wd0FWXWYOqsId8Kk3/SFG9y/gw7qFJioD4AGTGCneof8NVMM
UWig+ntalxqNGgnziIj/qTQFgsY6gtsDVoeYH9XM+kC2hKpqhav6Mi1DKwdt2C/5
ZYGxVyEj80dbpZdPvBlVfqazMs/ERzCLd9ofBfAUJBpymdKqIEb1UCQFJLwFsdAj
lAUkNY6lSf4VbFbrnAcM7pheABpRxSdizbQ0UEAbQ1oEKj6W7MenmY1sUhhzvNTf
pSAt6OOh+N/fTVJmjh0bvrO/ocJDW8kiVUEV+ZTLH5fHNYwa6rBxbLMl/VTwEC2/
dDcFCFi0zietmneEF7isJ6WkR8XmwYM5KrPa1mrNjlsHd1M++TRwpO8QnP7kBTBL
NhymI0+nAqrYohhb2UWkgxUt30rKPQu1S+bkD/oVKnR3OdGoMxk8MeHHXXrH1kU9
udvWYpQ1CrGKjeCCi/XpoCdPzoqhcIHazPxXngMBC2PTec4lIBEFE9BM6RrJtDet
UYf1Kd/6m58sKSsJ3GWuyP5faa1LrQwGMufM9FHc2cl5vyKp+4wAe9zOl8sa+vrl
lRvy2ERpmJikJZLUgEOMQyG4jCdQN4CMUJs45YjiSMAD6/LaK1n3o9wfYnmCZEBf
yTeeGGb+jmS31OaNYJh2T5W6IeA60yjnsBJMUQU/4Dc/4QYDOF6faCEPrLVmo6Tt
XWdn6CvO/9eoIV2LFm17Ft8gapnDgmgB6bKkrWV1WnUkwUiWrM0M+h3Uc8mn+kbs
muUmsObP8GF1v2RKPmUF0aMSkLRFTTgOk5vM78VvnWZiXQoQzFttNLqnvZ4RWZ4w
toVvejSXc1KEzzDeWXrAzmSpAzZfQCDswvUx9FlwkTWZ0RkiMljmSGez1GIZFg8G
NoB6LypPMkvUSP4dYedbOc+VBkLMJKENgNC4zxn2KZ/0+Ibm4YInEmWOPsjbaUGm
TLx6RP26vqdasoQZ95f8qPTIBYbjrsm107twy9aE/3rdNZJf25p/knk1eJWiyBNX
AFK+wCS20t4nJIBmuVWW7m/lMFy96/QO0rTziKxs0Qu60DO22Dw5DUETvRcwOjbl
m6h+66j8GdwDFpHOPzgNtKEs1gKtld2LzBAXn9Bqo/9C4dJUUZ23P3zuYQWDrorh
8oyliQMOYs6wlJSlzHAA1GosbNpcAdxIPfhGJQBfuSJWx722KItJg0e86ya+XPmT
KqisUQPi+UfX1cNZVLbXaR6fSP9T1RGEW1UiHSFXF//YP43GhP1PIe/J3CufKbX5
xU0LwAWppysafE2ZPLD+GWjZKvTL9kNzPwx47buTvSEtP4/j/q+Aprm+gUhNRh3Y
lPGxWZsq29HzDJIajrFwP7SZQYimWd0ZYOB3jb5Uv7K0EoqzYtN6zPYEPT/Mm4q9
hV6AR1Nc95cNG3ZIAIKZFMjl7o8I0YeS72QEu0CnHvb+ykR8QITWkjshgcgLDvmh
a8kMl7bRuoasYls3LYyrr2G4ErCdhm85nYzmaM79AiTGQ8d0bWAKJfMvbqv/SShC
sWuqb4d6z8TijiyCBqNRE9+usvwB0ji6aGw+rpDJMDbbcPnsSgsUodQwyNI6M+KI
ta48v9xSc+9bxH/sVWHSfWx2Ktv49xDcQt24WCOXsPRA5cix+cN4Cae3x0pXoQ2I
J8wJPBoFzXukDaHZ+kBG2kD+niU7xX23bOxrJhktnL8FmWQ2n3x/IQa5XyYfzYnQ
vnA5C5QNFf93/b2Hh1kxr8VGhGHFZGAMz/Df4GNAQK7QNGV6+eOjL+Q1wcWWqf4C
fWPgiFPDkksQcyWkWgwFPvHOYnnqJ+9+CVufj0GFaLBW8RNw5wE5hqtAzPf5STbV
/JTkh5q36D2joXNNk+psqHnizzQ4tE16dx/APztB2zg0niU69k7BzMHA8okpQhVD
8sjgg2dUwYDbC5EoFuzAdkt0/N3ctmamofHONZShQlmuHrWLqckNugzAAvw4XKfO
DEw2gV25gqQ5ozzjg8ZX4/BYtpyaEoNr6sVe/MItdqQENvHodRSKFolmTqVKGj/W
vscwlYmqzx80IoBwZzgrLSFiw1ogfA4aCjPf8mJZEuErgXxhOPX9raHYiZxXWK/m
p4OIuzO4QZbiYD4U0AvsZ2c2LVKA5mxMJP0xvQnxJkBCHBuCDmE3B2iXIcbQ4cFe
zqxI0bveM/qtvwfwZ8boDTaoDup4SrVHDaixtmcKJJJOPkXHSeGV1LRBYT/PtnGA
taq70cxquU7Oi+1abRxZSD6OfaJvPpJ/Bvz3sR6uG/Gi9zE2sFNN5c4fkEnJlUZ3
qzjLuJGU7xRXZ/oYCfzT2skGOnmstzn41qQ562oNeDupreIhi0yhJL8+CsJZlIrx
P2aGFOulYVVVoAV8W+7QUC5K2VHPHfFwexA0xlhKMEWgXEljvO2kBWmPsi+Ej7NK
nxHPiULmsR5vw0WTMErGXzB4MlQvYvagN7sx3aAafdJdnBV/OdlHSzBDYyncqSSb
MA/X4INuOqpPzZC88zitnHECj6SKS334zW302i+PxICL2ALo49IA8YOVW3BG6/jf
4IBZzUPm6wDQ2NnnQ8enFE1OWMD7LxP0E872iwM6+JxiAEKVk/Xqy/9BcJOF4nkT
ecuYtZn/d2y6d41BWIPJ6pl29LZPkowb/VP/8yRTGNyKqvuTTK75YI4exj0Sf98f
5UrtC8ybwTK2b2x0PBEMPbXnywDVO3LPE7ejeBwRle4oeQ4P3YNwRLzVxrwwE5Us
jNS+WotoI8JvXYuBF5OY8r75oJfW1Rgy7cGmsrIOnj8qRV5GR9i67V2RKqSg+gYk
E6Dy9H/t/8o3J96huR9kymj57fMqoJAafHxj6gZsqncKA5th4lhJot7hYd18j1ey
BdnZIQ2JMX8g90axK/c3FUYdq9o/RWAFh4qeSJdFkmJpBhhmcupXJbWwCUgs6BxW
pATV6PssD8/blzNQAms21rFlUsH9/UlTo+HTZWlNofS6TwttVtcWNuL3tgUuxdeg
NgD4ayeLpKVf+4WlAIA1GQlPd2+DGQeU9aIcgbdQr3jktPwfNeA7Aok2RvYJslJq
nMZLSClY5RgUW9tlMDCqakH39+xcalVQTH/vu6CdpGZHszKPaOBetlt/t3SewFQn
siBBCYRQCdLQtSD4X/SJU+a5e09ndYEzv4TU63FcmZu34HKeDwHBCdaJv22XAe/i
obvabRDjCC1kuUH3vq/QuyXIKXdC26aEciFo9qON/cf0htrBNHnkdRhL6iVFPOlB
P/3Vvg7K6VWmN4K++PjQFZLAZnomMJ3MhKdsnwonleCnYGHH6+ridpAFYwHYlbeM
EBKCn6tSY8tKJ+isAt2STvBOhva93kyqlzTqJ4KDTKUZ04NTbfAkf3JSy/TLWkwp
BDJTcrzsHdxFjMABaV357kMNrdT73W+e32yDbElffWW5I7SIEwSnqDW6sSm0eTAK
WAUJLqlIZaX9qWbDsdyoupQrGx9flFSpJryj7SX8lbTUU17m2PeOiGZJ9FxkPW0Z
PKWM38m5HI/r0inceiFT5Lwv1t9aeMy3bfia/xYrCdhiG0GDeiuKwomkbjvnL9iP
pq1bkeSAZiuyOjzGpghtvSVhrncgbKeUr0USkZ/XYcuPETFeU0HRubxti5Xk8551
ky3g4SrTqDcoB2Sqilnsq/GKq7jE1+pQ2yp2OiY5RercQwC1eCTS4O+WDrUL/3hi
merouBxMoQwOyX2fsvoyfq3VxsRHt5F+FJCXiaIe8RQ59hikfsUhZ1tlRdoqNSEB
xWsMEhWtHl6tbRx9vk9hqZcnv0Do3YgKyNNLc7gQ071Im/H6MUBZiMZxX7bRjpzw
wRmhd9ll6tlAhklnlajvhkMcCOHC/O9A3NygCuGDKCCcXQLaFkf9b6XjldgDyTCG
fgydMbUyAGwAwDHX01n0vT1Zu4561icEM0hMtGuZlnC1D4Y549DGWdnPkrHH4Gtv
m+upt4uXabTtpJVztCrHdSwLGqlQOgiJwmNRmAoKoawkoZceynIF2z2h5uvZOndf
WoGEayj5lKzdeKhZBgQLUMSqYBnuf3g68oWv34QdfGeEMlRabIQ0J2GtOqD3njl3
wSF9sZISTQiXNXJSn5lgVaHZNhIO4N80kxZNDvPVozEk/i1kkzxfU9Eey4jMXhaj
1+B/SouPdlaPeke31LHCjKQlhrf7h84aKNYCLAyqvgFHmlFyad2aOxdA3VRn/meB
5lUi/dqenrewCYx60CB8aG5Xjko8B5ZEIuXUJL8js7ZaCFMJFNoXiq3LzwWs+xIC
nLxHMIDergfaOeKJ7XzAscCS6pcgI/Yzjt3EP+X3xAxR2FloTN/ycr1UleICPese
ixKWgmnixGRyCJduqgmU4N/MwfZe+PUAqNUzo4XryMmaNXAZA+VyXtPwpQWegeU9
EbEVFZ03JBKXjstAk+a+lNYIqDmkm4a18yJsuf3vGb64Zp1lcSRk80xNEjOFKOoG
IMSpiTZ6Jl5POpdNRj2L+CDKm/IJDZl6LCtyRNHCGltvGcfqk1W2DpeNnsRo4dLg
TzHdBDGdDicmCBHm2vbuHKMZyzz1TraCVAt4utjf1tBDBWCrDlNXwWMiEtxa3kiB
R1gMMXlyTh9RU4rRxWDRRY2t/4Or8gAhJS05eZlruFzhq0MStHRet0XTxgYaNYac
sBKJTbBFMIGxK5MVVgE6DlN7IBNzQlWOtLbj4bUxxT5WrklsyFgG5SahCLr3wuIU
2h9uNbGFELmM5khrF/8VLiEXeGmrsi/5gvlwxCCZcuNATLvZNKq9OzHzg/SDb2m6
T5MRVPAVYbS+87aqspSOAdRBheUDnCdK9rYzfhTxDLEcXbSwHxiIH7q+Q5bFiVSF
Fns7WygopFi2PoOSIo08+sM1I4WY0FvN8c6hZEoUx6/sNzwhRxLn5CTkxw/IrBMw
/GN+LBurr+dOA3gPIG6uVt/fc0R+QEz6dRrPDkBppAdtMTGlTkQnZUKMSJFn6wwt
shlGOSjVkh2gD8HtQZYZOhlgjjQgT9tFNL6afvFmpPXbq+d+Yjkpg2j14h3QlaM7
oR7ETFHdauoBOMBf4htoSmkXNk5lHRA0NT/crJ6/IgW5qB7Ax1WUPWumAAGWU+mS
n6YwpLjZJSHSN9Ulvvy4GGN6zVlMnBfLQIvji0lI/AVX59GLNn0BBEio4/1AuNNE
Yt5tThXckcvnA80vTdlKUsy8oFyaWxX6Dw7Hyzh+GO8dpqmC5H6GzBarTJO0JZBn
tcYMIOqPOpwYHYZB7Q5uuJvrACtMi7gD1m+2Pw6h5kOs4yucp/17gadHiC5duffU
K0hzETyXhMQ/GzZZ4d0LgWG43kNRlml6aubK0/c9PdG+hve1MrnR72eihDxaKJBc
Cnhyg7GMxeNbmmKPjOdNqbOe0qD0RGUX56S3vJNyz8XXO4zENhNRW/9085P92emn
VIEEXA+ikdCvhZ7YcXvFQVqtUbTiF9EdKFyt7GtlhcLpriyIZV/VSVk+8w280yEt
c3u9JIpaQx2XG/bVHTAxo4FNlsiwZXhdb+derk0WixZ+ORi4haUHwm9QywO0soqv
EPy/Wc84Z6+BtJJMUaAqxYRPaRLo1ItvmXYQN4e5rSbTVzZWVJHHMBrHDfpyS43O
9ozvFmEWq8nRKuvMhKncqN3tm/GNm+mV3PBmcjcLAgYJzNMYubuvxOBff/iy/c/m
I7VYjnd3TCVPqYItLQqSeM+xo4Pa9rDOJo8vOP/wLque9efOK2xpdFy612gPkGu+
ewU9LzI71wJySDxHhh7Za69rtrgfLMU2NPkzCbmoBX2zfkD9oULsWpNLzDCkZVGi
/mylHoiyTlCAERs/YiegMNKr2iTe1D9hZmSCihg9rjC7scBhVAcs3/OuAu4hkSYa
iN5geS/wIST//hfs9C0WzW089gmm0y7Us/WOSEHvdqU/568/TbBYpEIlQNBm7WcQ
RiaP2Iaj+/PzNQoFK4Oa+rB5KeA6wfz602nrqBwDNwJtkyGTfHYB9NEx3cEhFX+D
WxdDxuVsfxnA8IWgXv0zqRd5bQb7hQDA6i744HeHSNYvQQ39c2VfwRXm/8WYbdlZ
lens8wZMGXbiqcxGi89jkEpEp5jMhZ54YiSDfxABH1WYKATveecS9oowrgi6RqeQ
oRyhjuWtIlOSt7ndwj42yxYmkcUI8wDH09cl2viXMco8WImv97g8Wwkisv+N9jZX
kOAXyhKX6zmd7qeyirvPoohydcSNflXYCI/ZMLKjA3ieR6bqjN3NFvrkPaAggXkk
HutTT0uMt0QvxrVOm9Snmbg6hk45BvMFPjFVS4rAI+F9Vpd1fwO3gwWtpXKo89JX
E8QPP4GJPL+vf15m7qppyeMmo8WrJeVff0N4pLAaf2v6JNbrvFnh933LpHar/Ef6
8CqPJIr2B2TAOLpZJZsLGvToWqbTvPus1ioNLnQ5qn1G1UHZ3aqgvtz36xRTu0jc
o0vxjwiC0JZp2kcDAQ1B5hTn3CuT7RxrF4zJ01Ax23teEu6Hio+XJxmm0N0Br93d
j3eB05xoRCNPeEY+y+Gb4ph2tvr+4a/u1wH3VVTNQ4DQ5FyvUKnWETqCr5tUg3+D
O5FumchUPZZ6XTAyvnz8pGnC5hjSJWncmBmupgyS1iEB9/agKkHt+CeNsZOJksqU
cyYYPUC6aSvrvyLrm9rVuuhlW8m4Cf+DxOOHQUoMXM2dlNiEoSIHqTNAeTrb4ate
YpY8Jl8oOFBSdyKLLKhisdDZHhOydSzUUQugqGWvdvuPmKUWqLw3DptUBvNbnWlU
/Lr4Hl8I9DMATHnAIKq3OBwqd5l0yj2txcErxDXRFMWXQnwzWbFEZDKntBt5SZBa
kL5PPz0nSt0ucH6D4aiuWMkv2he7smA9sqT4MMOAkk4e6czHo+eEv0FWfS8bbj0r
QbkTV2yc6i64EiP+Yt7GuHDbL3toxlViphqgbU3dJqEkTqenQ7cFiW5yEqFV7MoJ
BYiERbjlrFPJIdS6p5SxumG7RdYGvKFbApxjPuD4khSCtheYEgKHheTUjJjOsepO
CPpoAAKt0Zo0p+m/bToTbDuqGmZlxhqNuUuJarseOtt52m4hw4gJZ+nQIS44K49b
F/X2HELDgNpyqSUDwBabCPHjS1FY5xqT/qjVeIP5xTsfbZxwwpp4QSO1ykh2Vcrl
Nh3xC1i6oExgV06OUdNrab1rhxnEwnTu01a/9u87j+JFc2IGH8qVOCI7CHT6tV7Z
tWCOxrAKZuDq1ESyx1jM+omhy4f2DWaDKi15dABRUgBLOlK5AOf/JBgFpxurpFgY
kydh1mPNIDfPECWh47MzRmxXGNB3Sl3VbNM6lu1YdluSyxoiKxgwL9awFNnKi6dP
S8no7WoEJojc2x6DNwZdkihg5JIEG0PLE1RVnd7GTxy+faejaZn9TPDqA58DQu/N
AcOHeKW2/wMo9hCDr0i8k8CNncW1tBt16JrrFvOJxteKk2KrsbCQA922GhpNGQB+
/8h21jAySUkUw53wWuHU/rinKqySSCdyOC2tnTmUStepvTD5E/GzYKJvJWCfizp7
TMjehv5RK1jxlGz2LSMxjtRud+oUl63hc0ri/+0z6vRK+7QsmZR+TzBKGPcA/LUH
OBKQyMfJ7jD1RJd7EeNJPyUZ0oxG+x13W3+eQN6uQs4TSahNPMTQx+0JFEaNI/mj
vcw5zrrLBdvdpvYOO77W7nhtukBjvIAm6Mwz4wMZQoYZQBAttOSvpL1EoMo9zLoQ
67mLn94z1764RJ/PgZVWU5PsHC/CmMUpWrGGFtaUr8AEvW7t9aXPOaBH+J7IhE81
kBREslrQKJkfdRg/X/CZ/ES/Rysn2iGYkgGvpY8t07bAQxRH/2I+lIk/9FJ/50V8
4HC2qHbfL3qz7LvQAY0xhvWRBlhqBstY/QaSND2hbXco51rMHcLo1+gMlTCoVJ9p
ZCJVoirOc5siVvtHCqm1YDkU5H9sJa9DYcGSlamafYA0JnzMXY0nFjv52wzZzwr9
+inaO7zC2yYiMhMUIo5rkFgmVkUrGMEZjE0mrDvJoxyUD3SWgeZkr2zaBFbcdNJG
6XZOLcfz8EZWqTG6tp5zLPE3nN2Igky8jpa94sLxBgSosraGyNRFVGUCZFXbNwYX
/DJvZDZUhNqsWlZL0UUn53+7hV2A15wD+c6t/kbxGxx/uVTfdRpAtN7YfyX243ds
GWFpVhodKYW9NvRPAjh4IAw0Op6ra92/uorl1dql67xOfgivoO0SXFNP2jRl5rtr
+UTNHN4hhi7CI6rfsgShCqtkcp/SDKVrnmepRkMmiBozhzYnnnFnZ5R76CRDXpxQ
LcqdtUmZdiL4u86njfPS6QDztOeiFGpJfGM/v6bYgmnHe7dmqIE/c17IQqT+lL8g
I71G9+v9S5hwzfk3Kuh4dLqy6vg8qmaifDN7KDiUyc9iSfvwuq1K5/4PZJ40VaPi
avPun9WWbwvf9y0BPN4BhliHvQW8HRPUFcIX5j+z6N/Aes0ueqxSMQhSCk2PiE03
cKFUuUkm/xG744iPdIIoPRgZWk4VFrR/IYAYZQ2nbkN6MjvqnkSBGBN2lLwMYfGX
nNzgxKiB0KUMFWVOys2fYwjkDLO6BBkk1G6BvbUIzJHpGAgdKujFrnWCm9n3Laqo
yBpe0TCGlJaHK8/V73h//5/9OvzrYAHp7vbplz+7gTn98nJvgta49rrILatfFaEW
Mn3SMT5j9z+1w6RuKpFPGU68rPN1aXD6Jh7/CXhU3wFjHoL/MSuTqvMI120V3/KL
2xgLH4hESl2vBaO8POtjAzC1y4w2pPXrJP3lBpFk0nsliD4wE1hPSeIhy9iQS0ES
Qb6Znl9S2j6mSS0x35bSk5eiGQDSSd/LkmjHXLIp40754VAHE5kZlPxCplaxvO0h
731bwh5T7BrroRu2EauwDY8kQN1sw7+PLWmhvQrmbrx8dVZ8oU2aWFPw+jv+0D+0
4VaSAoP+31k/i/nua9B4NYstJ1xHh0Jzts32lh5DoOk34CgmuOFnHNSKB02DBUcV
l53rIjj9dQLpJ4Nn+E+J6CmuPDj71xp68yqcj7iwA/o5p2oE9dY/OG8jr7DIbrhN
N6k84tjbbOuJgrJgmne3fQfLwibbR21xu71sSmvDdy7BkefqkWhfhWMJ6yZ861/7
KZnQQ7ray+SOoVlqj9IUiFOn6TnLhwP9lE9TtLSG/QtIQeUxcHLfGi9sOIvVQV6a
r17cLYl8EK9KsSfLwJpekw7a2jSSagUwr4EuRUO9afxZP5Z1eO2tiZG6EeQJXTgB
jluzpYy7Ln4tHtJAkePkEN9wCub7xt6zb+4lQzoot7kJWSCGzdhT9GwKFPZEjfXc
wTXHsdVE2q3m10HqpOdtAUfLpmbpDZNGPxqBtVSh9xgYyep8MKSxiaTzvt7/Bj20
zU+upV7snMFius0eA2r0ncNn9tyrkimc8d9obeBb1NdozEalcytahuWwNbFklmmg
NGOGjLMZBGRgkyyyt92BxpcQ1fhJncll2b9HEiqFqt2H692DbeKp+JJrBhrXmsnZ
uY6gQuI5+AwC90W7k1nesmgTr1PVfwZf9pDNrVlT1shj7EwwZ7Ha75hV9TmPYOWG
W6SJ692QZiekXkE9JoxYq5WyBHSNN1v4mlLBgXnhSVsaLT4EwMmFclcrcPihAXIK
uIqA4Nq0npQqGNHaRMjS2t0XUlt1hhvMvuHVa6EjQz95i8dsY9rIJsYnPS+ZNfh8
MeTLnvDwSM90iSByiBWHCCkg6Mb4oPusAw7wA1pEOXOwso+ipR6DE6IpWy6EYwaW
SZcbkuBC5flWir/xbUY+pdn4tM5HvfgezlQdn5A62FxPjFwnwp2HgDTia7bqMMzI
StK/yVWkcRQTNZgGeUm+qPCO3Kg24V7Qh2/LBbFcrSYHOifC9/XpPVxEPAH/knaq
IxUtG6GFu6Zsdhb9Bp9w4vOuRO8ydWbvSlMtnS71gavce7egl5KivIVgikKIPck2
0nMzNgeD4+o7p9Qjfetz6m4u2Cbk5LreDALy+8hpPeMfsjQqBjf6LnQr3uriMLE6
rkqc1zjs0SeeAMFlzZAzaE+VlixBIBHtijVWyHVu422bgFCL0/cInFmTTIVFjRTz
jxFoEbRXdqOnoyLCIKbD9EnCS9c+Ge/91z4PQdFm1m0IkUY0XVhI46HA0D2wUsq5
DgAXD7SEI2hK6x6K7eNecWJWuBo1bA8EhtZTFqEr/UpTxjP7bnEqB2Y1qPHPcEtM
TDsmTT6BukDkmLVf/y+dJJSo1CLNRXrGy/aC+naHCigBtgB/vkOXYzsaWLu4ncBt
TgeoFNLVlxmo+bGw9kWg34Af7G3bfvRgwwtx7QsxmuV/x8aK3AywQ3r3CBCUmK+c
nAyz9X4zoqYPtsn3+wK7UPeanEOYE+18+B2GVWdlguea/MNHFklns0PmUiz+4Vr3
mdY/F5QCRMevSZBctFOT43fOhogLzoSQAndDMxGauuF8eLziTj3NDb9IJSI1haH7
23e+s2du5DIKqRcajusA8mufAcMntNNZcGd8tRQcX0AlH5p4826xIs9oca7WMtuR
iVO9ljKBiHnxrKICAALsAbinfHJqlmtFBn3fIBdkHiA+suu+V1SYD+7w7Om/81ts
JzJ6lrJ6o7AxNX0AvL/7lIZR/79iuslU9XHQxVYmn/iin8bpCh0V3zXL32rPXb6M
bXWz3FX+OmbLPPbplX0ibSE2ad1ktJaRJXFfnvnsmJLtUVHDiPqwND4b1YxTYrbF
WfcIIL8zqlgYxr3kcESOHAtOFtUEPT/FAwauM7VU5SIMhrMthBwBJhvQYE9kuBon
blhxrKWrUAUQ5peCNW0ML7Ef1yZ8k8jiYPczDjVERtBnP6V2Pdvk6xfTKJC4zSwE
n4YAiERRkOXvucuLUlG+ajWRtssaZviNv48AW0Ov8+ttwuzMrqeLo9sgvuCJEjav
rt/9hN4FrOuMEByUjHfpj0lB64KjI6PX7jHRm0SygrFroaCgqcLUwIhBtsLSVYZO
szNww8o9W2GsanOxPY72Tqkpe/64n1OI9pimGfI1Zky6Ib/qaU/wzi2ECn5K2/nv
QcDOU51xEwDvYgydKXoiEPuJsZGc2AaNMit1z5pEqJEXpJBg0jrL9nSrRh+7JQrn
oJJbiawPTMKYJMQfS3Hj0hVDfgZxPFQf8hSvhA+GhO7eRJsBqCCKlXAlOkaR7wTZ
OI5E4kl52g/1Mk549kNZScqirt52rsvcg4I0Mg4fI8MQ/Dc/UPH8Tk3Dv1PEVohQ
gv6cCzbuAHpO+3nL3OBu5Uv6J0JF67LgVcXhnUtyktE4BgXedoz60nTjLI+q2L9b
0JSbMx3r9xEOw6FrmQ69SWuhId668zuTTs36fimNefChKo90SIIGoRsAZWhdx0rK
moRUv6InYApL1JcXGAr44kOLoQGzB6bQF8h6VCan/FtmJAo6grZST+NF825rwC9+
5hugo2jG5U7TWzxQegwWR8V1mNAf8i7f30lXNASsrz6aARHnupH58hEAn6Hdbm0P
7vgDHIFoO/eH0gtz+3imlHE16L3AQqk7ZsLvhr83o7OQo2fUum/uqHAgzMIy2pQ1
8OD6v1QF135VA/q4Rl07BApCD3mexufDnl3LW7z7VLVFYOy7IjrFnXuqMoZxRnkX
zcsmDMT1c0qJMiu6yewqG8jzKzScjOIAVUUo7kfu59QK7SJLXGyqVAQFfSmmCYKx
GK/Zo2nePMBoq1zDDbtjdRqlExp53JlKEOc+NFxucZ3i897XFW65jHQMGwbukJ6f
EJy0k4O0WddQfN/u2woRGkX60wYEgoKGdALqQ5VZxYolk315DI+nfgcZVD4WxF5G
8wmSLX3RA/1eH8XlBGAtHU2zxu6lIfjkvMtkUGvRfwQT4ikJMyZ6hKjkr8sMbuNM
+lMfdAw/84Q404WDdnYE4hTUJ7NvBQVqf+JcyMN3FmHSbeQcg3uwi4zrssjKhI2P
f68xtmP7VJYeVHNC/EYU7KcwOa9pUdw0stetY2AkvcB0Om3jzokZhrY58kFkC7Li
IYYBL2NKH/IaFd8kif5UDNllEs9A+Hzu6qc8sa0sbAWlloT7P7yRBbiOJPfrr9A3
Y17N6rqk5PKkDsQrgpf6qSBXOyUeTMK9lkWq30ExyXksXGN+KCYL0wys+8o0loBC
dHt3ZFGPGHmsSuix1hH8HDiulSs4qzKtEUaSWGOjdikUtzo4duu0/I9HdAkMihi0
GzaeOaARF3RrqOVTLO6jeMhnvYiI2FB7kXnqHP3i/z/xL+hpphbJWFoeGadDM0qj
aoqBhX0dx5Q7D5PPNHZzYfMrPABx/8skZun1eu5TnmuvNEeYYVRB+JSHXO06DAxT
TfbGJog1jO/7LVeyuW6w4QVATzmC6OzDhJ2eNDTS/2dPwDToxKlVQ24n35XfANxg
/H+nczCXnQu/x/YY5mII6UKYH6jsUaqp2JsPBhxYm9YOKalKo5RVgESWpiIGQUNI
HGi3Szze3gQWfXZJ3o6gQiiFmRtPMKdIC8vANXTOsPend6ne2AfxrgfwvQfqrqip
In6PpGxAV7IaL4NegGswtirvp5IxNbVmtQJcKXRu5VAM1YDo0M/D6eFACkw5vJ7B
bAOP7aQeMN6TgBhEXB/7vR1h1S7j6nAjGlpwk1O4oOdV5U5BWeEPpGL/0Hfb+e5A
BhLzhNfsHFNAmtWQIBXtE7NTmiGTfJFvURpPBxicaFdSACndXsN9TUnPJe8XS7Ew
OXtF8Wtc3cKKYPOFzY1LXNkVvSAk/PVlFef2ML/v7CSdT8RRm8E62OBVYPaDNk/S
Wywdn9bI2pue73QYFxiHKXqwnuWiPJDREAKDTmex4+M/p3FpkxvtChhr74M66Shk
NWOv/gIWPDIp68JUXcdE4j8DWEQthDGVIzdkxazNKJBjzyEmZu7f1HLjUN8JIqxj
q1QOtjzUbFOg55XTE4tTngvS1wiHVlMEoxRnYFlHrngQnYMUQ7qkCIIXX51ctWO+
/IISHHeivRcVnuQTczLLHRPd+ZkjAJiUxryO7KBOiJDZfitjUyD18aYDTP9hpcxy
XNBynlq820lDpMi4X6ERHh8CVL20hibGBhelBA6A1bHgZnuZ98q2+Kr1Q79LGpne
iOukyX1un45lmYXTaY2BVFfHgB71ZQ7+y+qK3ezrywLsDU2a0xiHopDZMWmR7ItS
PywzAgnj5Vk+0RWjPJIpy/Ry8l8VMT0n5/Mxx1U/5mkhUIVR0bjtVrl2xMoOCv/j
G5p9IsZ4rAdbTCDma7CAVnrHxpx27AYrCrTFJuUs7aNancpWK9zIA+u2R90JkJhx
48N2XRiS645J5Q1ayQ0CpMUEQ/vJHoj1P/xE+0BuIyEA/pk8/i6Vq8MeP1BQJYu7
PHJcQat2+KSttloHmnq7c6YtBCbouM8NXXywR7p7qWUDyJGmzNsYc9GaA3Pd9A+i
8Cshe3mqmc/deoqBsCCXahTMc8CGyM6jQwVFXfCoZWCnCUvzhbMx04HHixvgGlck
SryQ5eal2mZhk278VuXCXdKs7wmLWLEf1uq2odX3Hvwa+hAHLr6aT555PqKh1fmM
xBfhM1QY6hOATwH/qBqadCB/yX4n3uDjDBGFia31zIYvJUCA/NbAHwL8ymXhtV7+
x5Ury/cO+gqonH5RCPNcDlUNq2iqsBnbpW0gz2K9a/YVtHNahuy/7enTtYoWpekX
evzI/4payjfEofeQXxabXbUZXRUyypvSICogZaJ9OEUDJUGWcsp8cGkpm2H/Wgw8
tzkxXSptQTYcN7zkiOYLPYWanL/30p4Hta6i5pwlNarTSn+q1GXKoUkW5R5VTaQi
HcxAVmbMqoXXVMbx44MH2flxaQ7cyWn+9XCOGNG3BR4lCabiLDVX3LZpYl8ZUg9c
0kD7kZtgLLgbqXpTCOlnp6t7bQavufXSX5bWy1C615Mso7zzuR53GsLfLZGBiM2T
TDXD/LiXcFo1PX6kPVFYGHycYQqWSmULnDzz5iXhyo4HqhULfhpmGn8zD3U7gC6a
YJvRalqJpiCyalW6Zr8rt4loRk+P6psTXlU/ymhRPllCcC9bCfHQMjfnL9FoPWMg
tceiO+z4yy/SGVXCAf2JPgOtxtqVvbWG9LpqutSRFVMlA+eqMdgt/jPg+wpDai4I
gXXkI6SVdckHTBrXwZPCImLktMZsooDuUo8ynGWVb09gfPiSE7b3656fu7XbGRk5
sI4JRD/qRb9j6jlKDwff6lBR6qCWBwqx9zvbuo8gv6NflsxwiosTpnljPaYJniTd
nR/uc8b/S2xh11HP/EIUoxlGzBQkMqRcBPr1H31nuI8teHfeFeT5lYKV4bmAJu+z
5KY++8a8MmRDg2tz8GGiQzKmzsS/XGCOqUvAuBSTKdYJ+kl0RY6Rk6w0BnsfEGjB
fZFcn0h7bUJEejP5E9pQIYvkGQHSc9LCh4Q6ibzYubQUpQzmw5R6cPNSu3Fj+BRm
wM8JaoT9JuW2ceIYGveXr0/ETokf/To6hgSbJgRwL1tA8qr211gL/WDuYBSMR+83
wWz4lhU9a1q8L4hRIAsJiJvEEMAcxKIu0IdaoKo6aU0dN9+WhxJFR6d9PZzZ5Sk/
FaZcOewQl5uoGEYO9DUN4L1BJMkUdAjiYHLfRa/2MYHRFO+ZN2lVkR9uM9o+9H0m
szqITdF9rjSicOti5JrBG3ksJqdbLLev9iOpoZ9yqzOhYBzxzPeCElYa4iY+3U13
UihZYi3UQfV6ptGGbwW8/hbDo5oROH1fFymCZT2n4EWv/YMcIyR2GNXxfZ7h2aOw
Q7uDFX+ZrdQPDWmn45nvavRj/REuD7mwwfggOVa5N90ogJ2Do5DEJaE6NzbmXMZl
DmxWexhWRGQML4W5MyvUJNX2cG6rKinynmJBuQWL4z7jAllp03buJWbDgKtF6fXV
RU5TXPYqNH8Jv8j4lh6yb1QjMxSyFERcFf50jyujy5V0JuaL1XKm6c+xZV8RxQGk
vZtaWdHIK0Wwqd2XGjuDhLt67t1pTj9ZjHwm4njIUqxM4aGUcrWzLZbCByR9s467
tOkl+R68Smgtlin3Ke5s1OaS74cJMlKvGZSq7thzAhDlqdxBhyGThAnDwbeKcO/y
qhR1JmKowoJoK6YXSZZMgClHueDaNK+iPAF5o2E0dnQZIpCyp9Q10JldnzHpg7nM
bumgzmOJZiawY5vDVM1Qs/doIeA2AAn0b+13YFt55wliB9gzmigETFxnsS+Ya/UM
MqMx+12vgP6LUbYg0RyQKzw/KyZKQWSJwaUN11Spv9mgc/ulylrv4dRCX4feZe9Z
K0vYcgC+NsgeXTaB2Bz27r+4M4Q2Au7YhuZ5JtFMHqrCLfKNd6LIx/tFIA5q344c
Gq33Cv3xMtOsoBoJ5/NsRt8hmS8Zku2fTyIyvxMAOE9QcrRnjey6MnZviB9/coYi
kL+TnQSJbcvf0l6cO48na20i8HV/6ByGRQPCIkl4i+mY+wVoxIqnHhLN9m/pC4WK
0isTavgRBQGrj4oOAEWo1j3M0yl/sMZ27JMKbOSmT8XmjQz82u1lO3+ndkc2BDFv
AycsiM69EMh2qKPhRbCmoNrP09Bcbo/RdyxrWp9vntxn/oYus62rAlPwDN9C1v8V
RiRaF5AWlhLs6IUu1kzo7OXp7nyCpBxy7b+JFTvRUWwN9K60HOx9jjEbThhoc4c4
54MjW3b31x36K5bgWnvev6WL/ZxQmZwL/uPanUmZgwordklxGC0uPl5SVRtRf4jy
XekVQnyBpMWx7PVI4qpeiV+E6xIafkAhzaoCeUFSFqIeGAW7QX4XSfNvlypqxoFn
DW+3EVxsPeF5kVj3PbqN2EHHrF+129VT2rGN/27PY4FPR3dkQbUDYhNyumb5tOW/
LgXJ+2oOunvKjaA9R6rG5XpgpnVk8d74Z2afkh5P04WnTsWv9s5vCNG+mBF/zHKT
XeTc74IGV8VvTewcT6B97+71XYP+rwQsNJcEGaN9AUrqnc/nxlYLHTAz725etEgm
YGjMFga3AoMZbMvH+hap3YkYFEe/QBK9C08Y5AGXqLSL9WS94KI5rFn0SGguPIKi
jTPfMAu3yfH8LqqgCWg+9stbUJfTUbTbyz54aJEysK+Nl30xTPdqJtuAsXYi4eXX
LYxFYZuZQHr7ugLxD5AH6aPZmhahZKygEMFu6yK3XGelf0nK30K8iXszYwtgLkMj
VgwNmDQb9uQKEwVccB40S3h9HsXI4MfK9T+UfC0/qX3kRIw4faZvIJCLOXlDvQSG
ndnlnLoKphtZeeAaKe1S9EkhT+dYd1G79p0aYOLf2uajMoOwFizS20AZGTlzGlH0
yVaRJ1cCqO+9libb7PuRVLshzxyTnfPFCYL/CGw4HI3Cq8mWSOzpCLANIV3V3lxr
rO1t48Dadppi3iwnqt9vCWL47aQ5vhiWVyWaO0W4swDGssPVeQge5OZqhDjlMGcM
uzKdOYr8FRKcfyHvybiyeCby9SeUaJTgJ+W108yZpYhVzU5KYcLKqzGhaKlbPkw+
+0izOt28l/1wJhW9VVGs2M8mWbWb6AlEhAMsL1Wx2K0HLjn0Pm1ds3FiCI7rtmEs
3vNzWY+OmvKpNb82b69klFjA6pCSZj6noFKCcUbV1qhJbh8OEQn4+EFwTl2A9XDg
1iHH5g179XqwK2JKWAN8vaRxfBF93obPBBwbFPq6yDgPgiGefd04VTdG4p1ySKP+
W4F3OwRux4P9AammwzkSqEaAAWRq6zGMYfU6Tw5EvK9lmpabIH9X1VZrgLwnSPJx
ne3iWBwX1GlDOjHJGQMXN5ccqbkP5FAaJsfP9BfKFZZBCHHNRB8jcxrYRcoFWU4H
zsaKc8OAYob6I1jvpiF3Qzc9AVxqr61XBA2n/Ee2vHfngproUHTabwUtyXFmBTSK
GdObHrIf5Z1CsVMYeiAIksihaNOUXBHC9+x/iTXG04/L3WNeAoV012NHdlFDLoKB
PMYsF1zhm7ZX633+4UAyRx6Q1kcvRRqXab87dKSYih9i9LvolQ2via1Nhi4JRztB
Z/QgDpq1sw0vdaFipH91a+v/lv/8/LbryNlItJNyPMgjqlu1OVJxJlq0bmw5ntov
V9azNv3g3rADZ2Gw+2e6xzxpBFSDdv87mMxzUFEZLt81x1Mn1wnxULrWIY1quorK
VrRO/jQVeay+Cq3RmjM1ryvZHAeeUpzDT/6miTqU+7Mh1IxWG3W9Q9WbMi6+OZf9
vi4IwVNAaa6Wq2XO9UzuxUXP6zKO3K1Y87DnVgNmglamSH95EFmTSRyFwfsQhOOs
orUPM84cHYMLsd8v9IX5G4iLk26dWcH9MwUl6YMn8JvNj4jfbiH4JUvs7kTz/89k
bxJdMzIIKTQ5Sk1g46dKZMXEGkU2ojGwvj9+Ot+ZaMjO9lid1Jr4PKtyKpU7DNBG
RChY7IpcMiwbQAZaTLmAt//NyKo44ifu5Vl/RZOp+MaUdQoh4uwiUV8sqDyix90P
6n6A/hae1a5aJp8nz2jz5rexKUoT3e0I4Wm7y8wZ8sxESV8mxl+3IyRIrpt8e4XT
kDkiWBb+5yZRDvuLwv2ZX7P/108q3mcHha+W8J+7j/wS3ppLv3bWTmTrQBNlCMQv
giXeTkrWD4LWRzDolVEUVQhY0vy8iI/HoT79VvI9EoCS4y3Q26Ez2RQ/ETc6zzFY
khY0liDLVyZpPGosKX03jk+YEXzqyb00GooOvxM582UIixI5/kZFRaafjuozUeWx
Ggd12lvtH7D7jp4vimB/kqRmND6+DvJZw2YPEoK9YSnDAnnEWMzITFdLCIohhZg3
jMCKlNQ4ZJP/ENcJFnbSMmLOdD/O8WWSqz8NnhgY4/5UK+nps+syVS41n2LkAQ94
UGaTt3s4f88ZShlw4IwbkK5pF9ZkuWubfBEvJL/p0Ws44yZoqHEdihwIPAGlMdDY
OU8raPJagY8LXeJqKdyPJpOuamn8mpL9Lqt9bardKJgMGwpeBE1AG8QiRub+jkrJ
CZLrCkV7nrvzolaJFdHHpM4mwnIPpanciIVnQZSaA/bD1kULpyn6K8p+4rcKVddv
6F1furH7jnzz9qW6SXOEBRZapHPmAxmsTf0ezdFGbcpVPFDuBs2HmWqltuYIopyD
rpFCQpOP9sZdBuVtW5ECdoZRf9yhs984KVOkvjC1Wg6ewssLb2uy1+MVP7o/KJsL
b81Ty/DdkuEGDjjZwGhaOY8jpWTxEOHe46xGCtVqeAhoijGoo6BbzjLxdFb8+cMu
wSy0a19SWqMT/yymBHnNGMilTftex4g5y8eUE9NDRObYpVEiXCjZ3Du4W9d5DzCz
/a5mpjMGygGuKUqU9JpOgYSwsxbx2xk4VEiZKYd2OGjeZljcAF5KwnIQ37bxwKnM
gMrVcamsvIPxM3vKxXvOvhGl3eikv2ZbFCbBSvp9oavcBjCDl0EL+hktsZeLOE6C
3IFaCY9QuO8PQCm7gBoi1Mhp7Zp/DkZhSsybrTX/obuD287ciEywOMRPOu2n5UFi
ZTE4A66G6bzYFxMfj4005F6qrL78ZTrL5pfUyqV57tO7EER9RcVSjQE4knh7Z9rO
Nec9/i5HSCSL86NBBbXLpwWpB5O05295I4PqpcGbqiIyxAIKqKrj+gHsP11aWUmx
q+c2yN4/xEuG8d4AFY8FIJGYLgvbmFKPXmVzVJBPCI6VYCuAmBXHN26oqBvxmII1
ePpysEzQbzRDW6X4BoI1Bz8dApuR8x7ZQetDdf7N/E0mzfW9tM6gfcjy/ZtdtEMk
Y7YSRAoYO6dlq73GH9nCdmEIj23AnXW2ITxn6WtiYlw5EWB6G8A61ip2N4xbRaBr
+oRQy8znHAoLyHq9ZWLEPpOtGbO6TDU89+NUJz+GJZ1z/5umx+cTrqWgoAjzmw88
ybkjMFoaFeuR3IIZqY680DHt+Ba+9Wz8vdhOfqvztn6eHYfOBcjOdYpZCVWQ9iNP
tg6hIdrVP8+RXN4F0n6ShFm8EQ7sz0LaAwno2AJnORjJuly8WBp/YVZGoI4Ta+Uu
FL0t3xsjy+DrCLarnm58eXgLIDz1My7+1xscbeSfjln5xmYPllR7qRfYDBL5jtgs
66KUMhNbtk4b59E+70QvQ1af+OfJlmq9xYNzOE7yLSvlS9zRwZ6E/uEXmoaqVYDY
G8510fpFDgOm9UAyOPzUbgAMqF2L9BYoP5Fm3fWzcAMQJ65YyDT4W/gcvbAmhsoK
tYZjObN+kc0W5Z9dt4/gB0PGOACWik561XCJqD97AxKwY8rXDQalJyP6wkdojukh
XRdJb+qmU287VZRgvMTHryKBprQrXAAAI1OEDC5Q289j3EPNl2MBq71UGp/emP17
d02U9ktWNzAl52+3UxmqqP8YbUdPgvGeKJi9pysx/uZrU6+1rrq9MaHNFfh/Hq6T
g8HJW4eV7JbBrdudusto9bCZoC580+lOqL2QfHhSAx+ce1WsnQy+kYf+/77LYI1L
wA6a8BfY8LBhI3qgWyEs/RdZpH52MEUN0EIi8p9KHU4nEpzHpvFAgUxxTIxk23pu
zUw5A1+QAqqp7kgw0mhOP3ZTJwCXYKP7ckxQ+rcosNeU+Nt82VxUDS7dJXjyYCNv
+SlZxAmI7NnOG2+0MUwRygHFmrx7zmSjlHFj1KBSI2giZ3i/2xYsbIqikYI/f0SA
NZ6f5QOpQuI+CDiILCCuAtG5rg5K9OG1IeNxOwELJ5TMZ2V/imuKc6y5GON0Uxtj
78sWggCnRx5R2PrjvktdtI6HQQPO91VvEDqyNHYaFMoyzzhUl6aBhsdEQrZKpdz0
tsB6+0O0qX3mONV4Z2heyNfuWBGe2GBiN5EEMp0mSS09gT3VtzOmbNrHzH4rIEdi
ME7w06bQydAFheILrkrBIcuXO4/lBAQ8vy0xb/N34keufT0HyaZlXUdeGNWmIiNv
vcMoLVa3cJ+VHcjjCN7rL1RlRQoM/dXfVePwIJ7duzQTmxs52qFDonkYQA5vnNYI
2gzT8Q/UxJXDqdFbaNPfz3hBbu7XHrHPhkDvOg4PGDYuN88+cjZFvsAHUXLQXA4x
GSPqcbEElnCqvgtcjpLlNN/jzIMwAfdU/1ok79g5MehDQ510Dt7IPCZYpoISDiPE
BBKgLwSuxQ4oBrvpYfE88p4p/iF7Hj+TxxaewqCOT+QjvptM2FW4F68AkSTH4N43
0XHfE2MteqMqMtGrQmsN12rIri0Q1iGuhtoDHNZOYm+87FDx7KWwqs/Lt98C6/2t
VxvI+UnNxYYDCNHkSJr5PVv7tEwUpNDWI4MdRtSfX8TK7TQvJLrtBsr1wwoUCfSW
sGps0Ny2aTfstGdkREmiXtXAip+JBVhWTnIO1hc+oa3AHkzfp7HOBQUghI3v36rF
uLS3jajDapV/Pj+plZPYLW8xnlCwEhApGjZp1OSWODq4CfWwXQDrCyI3n69rUMYx
+iVHjjxhyJSxQeGJfeSX3ho0JB/SlOrascKUspRtdHx2if1IVm65lKba92V/UT28
vT9fqgBMoyInQmtZesuEnce6s2Ip5goim0mdd9RU+4KFn5kLBNJTyyAl9agGMMFr
Ecfd5VA18iFzR3IPzIgUWM5Wo6s9MeyESRtHe+FoC7Jjugh3EAopLeC4xSB5ZOxP
uCehBT3BdNmUTSDbZ/TM7KsGX56j0KJGADM/aXwqdDAbpeNCH4BxvSH2XfXKK5Yi
ZDATJAw1pTrMmkw0Ry4e8ZOGVz4k8BTg4Fslj7lasO58MN9qSOQY3xz7z5ZZ+LQX
jxndlKewVpJ1ourIbKyxVXz7gufOvOqG81MkDA0Ki8FVwq4fZdMkUMFAbsilQxFD
qLdR1c8t4vapCCN9+IBZyak7f/8FQiInVuSI9yuSUnJRu9CBwsv6jHwkQnYSGdKi
ELbcdaAMnEhWU4FEdV37vSfmaMclcB0a2tlJDdz8SVB81qSQXcdL4EQhGCMgAu6X
Xv6OkFOJc63ItN2mNCq7FuGib2XLgFeeWhPvgVNilPHjmP6/83TzCpCYgTGleBAH
mpwIYxJxNd/LSZ/+W31apJdlbWnqQMEokc6awP4DYzJnmMlSEeb2rmemM2hRGxCc
t1izWYbKvIghZpuLUno8/DFRcGHtxCiReHl3WS+/5j/qVqFO9IIyiU9zdOtWyTwe
hszNl/7anw+RRUKsKyP41tAqgYR+5IAzNSx8TgdDgiY/YWt93BylZCUlpzekkvzo
hnDJgb7OgCb3K/aIcCacCIG8oCqJ3kdNAzH4yqzoyUubCt1j1+cfCLHo9gxLepwA
5IjuYleGtfUParCXinpc0Bda7my65CxwKbzx9DD8DzOdQ46wUVXSDOZUxuHpRl3O
MeTdlSuALuRmEF7qzCiQ8kZuT4RKrhM7jeG+ZBzMsZve+KS6RzRlYZsRd5YLSI9Y
IfLHK97TJa3Eom/l8mpxnX+zaigSsb3VJxlJeyFSrbnvocoElBtwAdHWFXwtcEM0
7Nmj5wm2KbuoeDliePRZtCVI5CPmYU/jjsiuZp1AtIJ31ChsdqOfm7QLwP09GoRm
+fMrvaZoJFrEs7BHkVaRVIudTBxQ3VOQ8WH2BcNWy5ojOLZOWDCDMCMtkRwC9/9p
Ks3Wli2QJWE1l6guJtQPSDaUbysNNl+3Mr7LP6j6kulX9ikZufBv9tBFdsRF5vsw
hklTC6EeApK6S0nrtMH1cV/J6/KC7Js1WpLZRoPeqUHyhSA1Zm6J7k5sYeDA3RnR
wrGxNwiLfDWvkSWeF+cbDd3T+ESNPRfMICETNuYfEGDwKNTqutAziNpATssVneU9
/Ng6/Nm/bQPSO2Cl3SIHbaMuJ2hFceCd/EyTp04FDwciq8VS7aA5uh/kIEf8gvk+
V2+yCEKeGUV8lQ+h7bAssvB0HSINsWnsvrnUdp+QmMQfkAeYoll6byBLYYBQGdcC
SW1U2+I0hCFGtfTEJm4rPRcC5wSSOrk+enFVBpJUr7OVR1IqKlWhnu4LJ2IBKe8P
cl+aMwH4dDzCqnl/m8r8Wo3NWGsNC02DC0KvDgzUPjHBOZtQsonNEo9krH1qzGBq
7dwyvUG2wKyT2kOo0hz1ZMn1qvVvv03a7Gs6mQOgU7SdzTgFIyS9Wn2Czsvpu61m
pRdlWo9pioxkNq1LlwH85mn77m61h5gjpZeVAONQr3QBGWB0rlbI/RjtcDvqRTJO
cZQCmFeoj1wp/Ajf96hz9AqD9hRz9gpmJwXBINP2c1FBpTVzt3R3wVS++6JHpSZX
TFLGjrdi7C+EBZEHX0Xs43o8fBe7ztH/zlGEAuq+f/KjaW19ktxQ0c3z0FXJqbJP
i1JSzwmRTXTzEkC8+mjvL8Htslka99Y8e2uAnk78MIvB1Gv4B2a78cy3CKGVM/Up
Kdwt8X5xbMqJxxxZhzuBqzPQpgP6UrjT6dmxEdHb2G5gIXLtGEu45BP7gELz8Awf
Jpl0D6CeLvV/F98of72qHs+IIPAJEyoGtn0GZqeiMmxMBvnKc5Kl7PqRzH7Be0xY
9JXHEJ08PDZO4nQcG/afA4sHZ5h/6g+mWVQXIYDLhcSd+zf0Vwk3rCyN2z697Q6K
n/0EU+oSMHHPadDBWEi+Q5iaY7rgJVN5X9P1jgLGIs2QB4zMeNmeM8xzdSruXyaD
CX09cmtNwRK9SfU+neidywIgoNbfUq9ZEwXW5q+jSujTaJoxEHNmmOWQOZS3U1/D
cxUdy5oazCCU0BRyGMQFGP55H7OVCpcOC3Lgb+HjdvAbCKhus73/XRKhUsDMTqxk
9ABDMg2m+HyNm9GR5wOhBYcg69lUpTcu1owmyq+0uuDwvtqbSTj8LZD/OT19E0sZ
8iISDmQvp4j4tGl5frmb/pFuv6RAKb1wIJPgWhO69lKTUKW5x/cGWtvmws/Lx8Sd
bTbg1JuI77x8diIw85PQdsALMCERYLal5LRAmiIjsBNW5qfiOAoNV/zgPu9znaCP
p52t09RoIjuit0zi0MQi4Sl/pi1oLqJLxYVVLM8sfR6Jcgghm4mnQcgQawcJQChN
OEEN7uay5hrBW8E2dCNgvERHuz4Ur47g/3ptAlh0DqJSIbM55CGSHVmKu3/09y1w
pEq8JdaGvSN3lwlhAhtx2pYOcXgPjjMTmSu0iRLeVOdyxtwPIAwMdwL1LrYozKoo
E+bXut/Gf5eYgaM/JhbVxPf1Y1UjKmCu+YMuoY77Iyz/2XyNqvfHX9j/pTWP7H1a
NM2uIMJLXjQXzGmoLk+IHy95tsEjeHZ6d/3HBE8nhmXpvQdPAWXUhMwQbcLRdD8Q
BnSxH56rxy8lLVnU2OO8PTtglXkAHMORPorWM2Dq3QXOjxiFdXgx3ufcnNBYpW6b
d0Fr6zLq9/gIIN6Upl5pd5zEOlbMp9SPuh4+/K8zMqKUWhCiiYQhFQlv6JrzEe3b
o0d8EFc1C1xPf/+hWIOQrIJOkc+GSy9LrSV0c0I3U8XIJyj/2CTxY4TeQkEDhWMc
Eiwc4WIpdf5uRJNUjUpUaT/GTTjyhL7v9dulUbrwDeoC1DEqkp70wmdDnPlwt6jK
laD6vZ1+x/1wn8MPJxhEbRXcZ7NyTl/pgiGvMGoUMfZM7Uoy++mvexTXLi1FNos6
CcYfIT+nkWcEY3NhiZIj3BBxnNpRGMYDbZyZqfvUqxPYyeEW6b3UoWkHVBDbM2bH
Y1lRe+oAWspSjBOQF0bK2hocngKaHILmzWBr+0QtXr4vcXAOvfeRQh7DNA1670lk
8bdsyg/POODOVup+KVoxCKdWALci5NkOFfigv2utIVNJL5CbOZgm55ylUsocyO0E
WitwOW7kbK+SeDqgy78kQzBkIRo8YyredArQ3yHWYk3cEs+23b7BZgk5QVYhcsl4
pm4STE3KYWUAdB5VkvfUa52nwxGDf7gMWqXI2iVvl+ue2yx8fHSRWZwGTVVCosXN
mJEk4t8+1plzgyqavrwaZ8nuCJijup5e0iBpQphxjMHyBbdenlUF7qOG0coogIsY
FDwQo3945zQ70Y1gkFEkHMs/80EQbjYP3Qsxc9yILrJK0aATEx4kO1AJ/IaqUeEp
Mk/mgAYQLf7mIK2Vftm5zwTdQ8rdaE1gxD7lFrEOc5rimy/wwQihvvpmndeN77E8
dUuDPsG/EmvgEYVo+Bn4UFSZXWpNtK9fU4eFlS7kSkmzT9qXELSrtdSy15AgJrS9
7h3AGBoA/A2uGpnU/wQAXFoPHwoSFqJAV/6Hu16l3D1U0UAPm35pj86sVwG/Bz4w
4km60c62jIFECcEls1VQD0/h9WEUV7f6qOdeB+t1EM0T7CpVsv4HrkpBsUwHiwS3
YNYrUVpxQYio1WBcY0fVKLU1/kaeRgOALX0Vvug3L5xQXUbxJmyzmtW0TDN3Q89u
uc6TDd74DvOJaCFnExZ7It2zyKHSSVKQMS0Xa11ClC1ptvx63BejuvwJnhNp50Kp
nk23N6EgbCCD1cor9DLIOvimVRiIVGOyZWRedzZNiR+YJMfSehqzmELhdAOs8y6i
zNkwbQW/eIAf54n2BoXg4F1V0usRcfS/0spowOw9sAJc8jceKjiZx2Fh//skaAE6
hdjNfYfGRD1WWorKsz4KnXkucrq+4cIQJqTerYYHj5oWte9KB4yijG+MH0cq313M
leHb2U8dTo7SOT38/buNgxPZhfTdU0xYRtbV9KWdBby0XFVzjhSJ9roycxAohZYT
Ff27KLO8swh9nl+hm0ieJEPl191n15jauVEm6RVTRLHh6AGdNNkxDRIa8SWkmWH4
c38oFf3UEqKgeNEpVUjwhDEEsVgndS2mzRLOqmnv+gaCPcD12LpZxU1nC/gku8hA
ECMvLq1e11rMJyNyj1PzWnxy1KRm4chj1VrZgogdlysnCsKgaEl/lVE3qndk0qlE
X1CY/li27vcdA2DE8JxWFDNJPW/fq/t2v4GiiIr5vNbwVENrpJeOZ+15pj6qM6vk
XvfZkkVHvFGC5mWtKaWSslStQD35bsYre03nMscIYeURZ8CPIHLtamkefqeMCsHE
WsRaT/etlvV+wE/ONRFve4LlsrAQOZYOej9eaMMcN+LEISuOaW7cvygEt/TUSg1a
nefyyB2bhwNnBZMXCG7a0mhiwvGMgOQmRmCaptVkyfnBHXRYUSp9y/vJ1rCs7k64
+9OHgC+JaIjR8TI9ljAkgOvtkfuTpWcPRDwhs8tlXsVmhxGs/udfTDz1Bjl34G81
EfA1bsCWhsLRwSGP6wMSFIVNt4i0KJzLK0Y8jy7XV1wsGaKB1ZLmIDYbrtFhTfqx
hZJpO6zJrSnWUyQK83ATNw5pAs0C6IPLNmFHKauW8g4w8Sk5AlpO6/CiLPuaPTKt
uwQIQJVHxdx4p0Sw+ilL3bhLD1unUrdo+EV2MCwoiTGgsjVFHElJeu/jLeCybnrQ
/P0xFDOcmfY2zrOIlJKD5U52lYlvGxyeVai0+vWlcQQFiXS/IrEiMAh95a0ifeJ0
+xTi5kvWlykfNyVuOA4uFdPSnVzXU5cLvpBrxG2xbjA3hh5LTSo/y3nRjRX/B+oo
r5Xcb8uc9Q6gP9fh4zI1CVk0xsSSrsO4UPdo/sZkB3J1pnSfRPQRLMAngzhD2t4/
YSgQ+yoPu09krGFAiyMQDpiLMsgPFnezC+kdJ0qzE2GH5YY2YBN+doGmBSZXiDst
fM3nUkm6JoZ5Uu7nsjicfyaNyLTujkDd0ENwNLLW+xMALcQeOoWwGTpTA52zQgkj
Z5wbtghIjGX7nqSyhIiHkmRTvwSipW6Ut3iKcqZnDEHx3dFtVtY+CgsFZUJmN86Z
AR5H3+HOnraU7ygBbXgqFdlKzHlX9VLEuLvbx+kVGeTCCjaKxQkp1tw+LBZEPqHa
jrpVL9plQw2F9qNHOq3Qi+xzDUOuNoSNveoUl0IRxfn31hkglBrhQgeCO0/prT+S
peb8AGljMUmsIVDToP9SQZUycYO4ytr8bYaSQkKzQMeN5zyeZc+Mg2eJbyT94fnM
MKEqxKDhJ0Kn6gLgVH+y76pGnRovtjyDCzTX/6U2dNWLxN7x2pdsybGjkZc71HmV
SiW/l190ORC0MWkyMh9U6+jLWgWFVdjXoYKF+qcoQAxZSNhlYb98qL5RKhk2Xo8p
XSxqFU43VB1KNNqDD5WxCKN6ElDRGzGE2OPDXizIxcnYijdG/6x7wIzKkGi/T7jO
AA64VIAOLXGbXO3CKq+ClnGGx6I0G1Xi4gbK6YUqhyyM9H2uf9Rs4u16uim2/SCk
VScwFKho9vL/Qip7Oa19BJdDi/WAH6pk0sOjBfAYtob2mSo5itZILqP+12Ou06cd
G5MxquVjmWk7ErS20Qh1Emv5D6XPwWXWN3cIqBodmb41btYz6A6o3YzXCMIBFbe3
cillMFpxZ+fXxIAjS3WDej2yafO7XppbUgClG9Lz3XjVIa5sJ/Ls+iIyORUztKob
eV6RiLfzzp2KSKCGl48+CYB9YPapKV11epTr/HAb67Dw8BQUK/uzQoQmt2peWO/3
cCOlK2F1X7zeH7VYglTNeUZnPtYYkM0BHnlHUU6G5ru5AQXcYBKyHuXqmrzpYUn0
QjNd54x5yqa0RNu5r2yCPuUnOW6M+9OlI1sVMPjTsMBte3TRgypZAhTy4b2zJpbh
pQk5gDA3vHzdiF0yHXw2sv++5sx7sNG0VOxeAtpuIhLVQBUYsj/EB6pQMZndkWdC
Pt2ObmFIgTBdvzfmeIAFWSjZt8EkErT6BiguZnpAPTKRcZjLtgAVbo/5R0LAqhRC
LWX2Qx+ULIdGsR4WcuTKa7D/zfG4bJnMGDOvJMT9tdcUAMKBGi9wg65/L3KRNtkY
XITMqUcvmH1fmdSy0cMPFktS1jjoDTyjufwZOQBtLoaTEqGqi15fhY1bQR164bCn
g7WRkWDBVG4PrmNL740S2oqoPm8w7nANTnnlpfmbzpB215aQTF8dJQ+Fq3Gb8AV1
6AFDd/ff1MwVc77LcGOU56Lf6pJ0BfmPoKZohMVuuQLPkuTgwQKLeRodk02aPWPo
YTHhaWvhfdi+VNlxyvMn1eVU2VUd16jUbbmTdZExoOseqwWTJmmQoyI3u9qVhzvM
EvrJIbECF3lxJ7L+6ypIRLJUeDnVrt+P3iN9J3leFTC/LY6nG+HLjkOOQNNdmg3e
9oO/uKwmDndJAISN98pqT7SRzn0nZRKYUOeN6Kk2nF/0pUShV4fG4C/A+K2HDLfb
wOMoOhxPEguS6WgKHuVE9J2pwQqINQn652m/IGlDZugcvf/XX9rbY+1zMhtd1O4j
EKGPFy/YxP4fYa9hkDeJK/swQJsPqzna+tm967Ot2Mgl08PEAxmMvUGKD50a48fM
5pLJk6GkFuvHvJ9UxsVw1kdn7feL9E6d2D+wy6Xevkd/bws1fwkHWbsoV+f2/Pp7
Rok0RugXhEF45PLAVTDsguPW5ji2qF1duz4x2ekrpw8AgQSXJ6TX03RcGcWO011k
h0x4rfxKbfcIPiY3nzAkxnvz+/pNtFCV89E2as8kqjw24MiXcdBl2viw3x0LEkC+
LQ4ckudFQFx1rhNz0z1njwQqJhB/vR6NQACZ10uyh2nx9rUlzDSzMQxpUS++WToP
GQyocSBXWma1/5uyI5n8EiJ6Y2ttbVXF1xLy08c1k22kdUh6RpO5TYoRvVoTRWWD
HINmmFvrs9aZGfmyV796QPtfWiUBlkMG9SLvmbSH0puj2+TqhqnbpVodnn4joZkE
IxPCqQQ/yk7NKGkWH6tvsYEAZguBQzYZCYXVDzBzS4hIJDuhOdJhlknCzSmvErdQ
G114nyWeWMtsaQzCnwrwDV5quJxXoiugtTZaktyrvtIe9fWXwJiskQVBW5mEJw+V
weGvmUI7FsXBu3i8Cy0CW0GmA69rfScLc7onm16p187SE5oHeSWV1pTK/TYfYnjf
ZuX26tPxXouBSvQZ5UHSW6PbUm3Mrn5J/Wxj7hgWtcpUrNjdu5SKLq8v+Ba/nCFO
/q/R87CLYSrFG/Vp6lD6XUJlqXhwI8ebMVmkRteWZmTzsGyA7AvIAI6sri8pGmBE
Y516/jRa53S/sESwLrGkCznPcYt1pZkUGPma9kLrB/GEdHYwCVy6aS1Xbl0C0vbF
qveaEmrA/Ml6h437suBgBI1b/z0qhYxuf1Ffp9IMsEcBPsjro4hw6NLMFS565ZZJ
pVM7ScnV6SVfK/ywYZLAAZtv+G1d33aG5fkZ3fV4xgDKETfFuQMNTMmJK8KqWn/H
qykexJqTyI+t/bdajn022B8q5UV3dxFTCxGwCXCbQGpMOtimh+7HeRtORMIN52nd
qOYkuTg+cMdc+aO6hTuzTUxClxghJsAhm5XZk7hBEq5XHZMbVf0X8GonY5tDOTZK
BwVZakLA6vQB8WnAlqjtBPiyxmNtg1R7FvXYf4uordQLhJD8VDOkNfFRl1Xms0En
dgSy5+uNS2q5bl2arAtW6xGkhOQu+USC0ExVRo7BghJY6PJFPAI1Q7woiwF07rzY
7fsWugXpG/e3I9g+0bGrKqhMNFOan+6eDkPvIPmGglf/imGgnxKLA10lgcrSZL3h
W5gwjaV+o3/QAoVHpJn5A9VewgYnmHN7eFF2fIoXe/8/GvuFXN1j57A8PsWnBWHF
ZskagcE+4oN8cmRpXWJRNp7HFkP1BsH1gixOxMY+FQyGsyUrxSjFQkJ/QA+jddqh
+wg0aNUI2k4pgigoJ6Z1YPkpmrjpVOJDFC5s8Zif+SW629DDbw+/c9LsLhkHTPoq
kjDc2jqgh36i3ucYgPZnz888PyCW9OLZia+kfNkH3KyAVNaQPwk45oEuihM5oRfX
sM683Sy7Gg5Cmzyx3e16GcSoSZOd55xPpFoLOEMnPe9TkRiGXcq0iq+K7wLIxxZc
FVlUDhAdrY0zUXs0oG1Vmf7rQKPCXKG7ZWobhseGT+wVCu/URuHjrfi+evDL84fs
+U1dhQfXIdBhA4gnIlxb5HvzO8WIuAJBmk6r162Y2Qzyrz/71WtRDKjtovVS0Vg3
d/uY2ulwmgcMoV+pOyM+1dYmpsBl/lqi8SbZeAoUsyupFY8x7CtqqgCuiK9bTIZQ
yJTks/FAXC3zjPzFjBDGCRZH6+FMnzcapnAXsmjPjy3ji2yse9dmPopqd91/nKVo
dwKAloFmiBCcETt6l63XXCv91D/f5ny5WTdtaXcIVcFjBSs4ZrpuF/Huicv2Ibul
kV8fRBAlR+OMxCFnRr/aMLFw5PhAHPkARpMLlEiHsaL0ZrpRR8aKgsUTq0s9M3YN
HHN1varSAmCewCZyBV6bgGHGYk1ZGx+ZOac9fioDWuwkFW+EXWf84d89aZ/G/nwj
G9unHGZtnE/p24A9vXCwQeXFix6wvmj9N9w6GbdtRF0csqG9k+kzDbV6HaQV3iTW
CD2cHleP+IflKSEoq2agJESy0+0FinstVg6zlRaDLbj6+Nt/DttdpDdJzMjH3aNh
XBRQIXdEyrGN3pP4qEkkU05h7Sh2dqFjxqfpXmKP3txk4nEY7OD4pGi9EChuqU4A
nyHAyVn6RF/MkHgpiTDJF2wGVnFMGYrjupu27u9aVUJR33xOPnn1B9cXbc+A0Ule
Z55gIUCnhp9Oe1r/ilOtdSoZh3fWpSlu7rERPzywR6IKbmvJlhnqIMbYCeECV9en
5VUz2XdgHYwUuTHJ0nawLe29NFYRTz6OgNJjgTiTm8BnS24n0EUaHBHBVWm624a5
A6LW0DfP9WGmYYK+X41cWWfwt1v0TFlGq77HYkcsTYsMRtJVa1N7/vBMIWWbKI6O
25BUelZ92nDL5DcoXaKdksbbuSTs0PTtCKes3GeKf+Md/a2gCZudxoHaHt8sH+Jn
bsriC/iC56vEiNq+6cSMRvNGeIn2sdGdS+Sb/KdNLNmM1wkivbcbku8EQomLvMQ7
TzY90gg2RKbQZo6yDG5C6oek+xVNvXe3qssVafutGXCm/AKnTEXtkmUtlxABhaw1
Qm1Bj/oDU8SWiUScbtZnqnIq5hCZ0xmFaKqc6nGO/qSXXG58gAP0+YGMPX4ayDJF
99LpA4jng6oc4bPEVYXOUz6aS84QpHdeJQ36wowlWmt7/bQyPRdc0Sd5nqIbGjhG
AEXojqUi4+cMAQJn33pYas5C6Wt8MiM0TejNuPsHfrkx7VsZQ6cG4/XaCsJbIzz0
ufe/qIK61WxTXTbqUwtoqAJKYRgxYx1yYKHKQMLT4wGAVwWNqKTdViuGvxhUwZv1
awiGBVOcjCBQXeUZA8th4udl3Fp+5NxkOCdLu+DYJpkQdmYRpzOpTwXaKo73eCnZ
3l7XM95mebqJp6AM0htbYXQahCnMtYsN+/Bd3ODW/NiSoGkMGvwdfC9hlj07H7eh
tMTf7gxtEGV4oomkYZeseFJtHwrvS7nLVm0LJKCnASuWy6mKZ+d9zJYCK4UJvoz7
Kku4S7ZLh4eYCNwkQrMOgrFRzfg4kyPs34kIJH7OcEAePp/dJwPsyBMIOE58MVae
deqV73PeKXqx87WT+DJMn02T6rzzhsxsteIGofdoIUaKHegygtWzwkN7R6bPm9LV
uBkfyDV8GE2WD7tg/JHP0+OyRbKrHVkFzdphnUrwQqCCJw38Fms8q/WL/qkRay7c
OWcVn3jwDL0zcquEwNaxl+U4bQVEBn1D2ekGF0OTztTS1RU48g5b9Q85CXk2lGyB
1N8G49NC4f+PBPNXqWh9p+BTw6DeSNw2qJOJJcXpzhlTWndAK1vRVpzHhdOFAELw
pI55WoVmNfPr9dRJ28HmIRpEwmvTh7Ob96xrYkJLuM1QnAi55nmDA4ZIpB5ijUHE
RXg6PUlck0QT9UQE2YKRQY4Ewap3ARq73h9ccE/0JUx16diUqqoaT96GD4R79d8S
wouOlmVps08rSOqnWij1PGBuZtrBEkCho04ecyWD7e5Vl9ozmLStIQYAb5nnKz7Y
SxhxXEUY1ubK9r5P3hLl2uqmLZ2iZQUAifgs5YwM61AN0AWCudKh+4OMFziQaf7I
5Y2zv7QIuf8S0f7Ss2fPv7GUMmCWmzFjrXwEJUmI9iY2t8DK+Sx34nNvyY00dvZg
8g8HbxY9SxHMFn5P8AIUS/3yVAOSD2qf4b1FQ1DQvGfte81gSkthEV3VWK9pgOeX
1AT5oDNRT0R0gs/KBsnB/gWzWUmGuHRSymgxGmsneiZ5QbrHCEvtbTQsw+8JTjE0
7WEUI4i7wG+hDyDdLezFeCvJ254Ta68smTlDWYpzgEmM546eAvMwvnDZQkoQZT6g
n4w7NfT/gGRXlMbzcxj8sN6l552KCw71HVk+/w5sgCX/8Zo2XfHk4NL/iFbdsBG3
JlBYF+R/wUQwHPJn22xoaHaBJqd84oQ0vI30kqMGHXDtzvJ4xYGdJUyOaLVJD5IL
b8tkT+4lXrpn1DPlt4Stk/v46T3k+PS1JG4su9jerOVp8ljIc/T+HN5X8SXAAaoB
r0RH20C8f0ttLVJg+/OkeED9y/ywRNsI3+aSZSoeXHaNtH6E5L6KHA4fdyiqTpsV
8OVO5TcDILA33SbgT1PcJtogqMw9A7iu9QttJfrvYfQmRtiQVpnE1XR+GyUbCbjq
ur3Xtwv4fw+UcaZOTK5Wm4V6yWlvu7ZV+VRyb6KFrorKsm/CI97So6IKiy0sk7ej
Nh4qmboLDTJ9SQy0GYfkzTpahyDOqAivQh4DzZNrmXnbVqMzQWz/X/2dKkmsQFVD
Tmd6iIBvqR1RgHKtVtWFJeJACKWt/Bwyj19kOhaeUtTzXFCgFyEROPYb9B5oz2u8
I0XpBTIUDGx16Nh8/XinjrARSBC1v6vUJgPilb2GK70EjH4VKDTz9TWDkOXZb7Mp
YuYfLMPKtd9r5/SM4fXriF55d/a15rbiVdudR/arY50in2RjbajsDFEAMfFhTW72
oogCK1Ue5mGV5UkQM0KV5tRwKXFMFQ/k0AETfI9TKNGO1KUTLTzbq/gmfGmrtOhv
XRH8fXXTrdsTPjhR4NY7uszkbsa2sSuM3hsiz2PtmfDyLAsg/DHpQBvEj0L+CaWV
LF82p9/5kh4N9vIKvljdofFxpBIoirgiw5ALerhsNSGjg3j6FNqL36Nbf1hm8tp+
O/g6blvDBlSioEEX7fDtzID7fXbNFeQzrHob8zfa9vdljycWNMn2X6H2WhmhZycB
eo8vSwfVSCmG4AEQfSLLBhr7w1lAboXFwFgP0q9zh5b25s8fSbWbEBL+Gp02YG3w
GICQzgSc8dq/R2UehZJOmEpFyIw0t1bdtaAewAYNdA/krNT0Q7hK9tuRcpavrwXy
tj+P2lVhGNwqsQCSdIggm1IDlljyh399DcoQktOz4UoHu+KXNI+4vbPUIm2wItWK
sS2nND7RIvZQVum94ZIlPvovAts5CSbnpye1020mIJPHthGGEbv2RNvaZP5ZxWNR
oqWY9otzBIWjFXvUG2rILihRRaHb+yT+Pzoclhm/ZMYU+wIb59hvvBcyHoDB74tv
Bp40pPUYUw7ak0jI6LdVgLt/mmspvSeym4cqqKxK9Hj0tg5yWqh/rS0VnfWOuDKg
SnkPF7hgHbhpbgF6j56dMPorvGN5i+wi+cBWgAJ2RnmzOyp4k6eXKmAqQfj5Agym
Q2zeL4NC2Dx4uZ4y26bAo+h3pMgKSlavzbG2nZAlGWkhHzg4O9f9gn+9UXMxylWJ
2Q7oW66cG1vpyAJQSUz2xmsVJd8XguICrZJwVrbdwcKUiwECcJDpx2yjgytb3w2W
ol7WVa83T3YUt3e9EFeW+VjQR6QQgtTZoyJ5cXI27uj4phLm4lRkZbdqGsXDr+5a
L8M5Jh1pUareyabPgMKcuVITGCJFwFcVcHchznFgF81OvIn6xCfawuigMke/pV3q
oaNkQPSym7xDZcQ5ovgIUoHmat1gQGQdx8SeW+/9+x36vClmX65M6WIPQIHkzI+S
e0a8TALYyI1oxeLPtdfU0SDECJN24edm/n6QHNK2uSRc8rV1CWyu/gJkD0cs/dFB
7qayh0k0GdK3fl2prIwn4MwkkN6hgVntZg6bpk3exzHtL7ADxYup8XRNizjzfGSg
jK6CnQjavgUk+7roA8e3UJfpjpaw9oZsxBnIkWfV3nfPKd4ZIue2sb1e4oJc7iQP
noCFeKpR/P34TEOTUut6nqnt+UlInuxyNW5/hb2kpm5Zni/mRY9rCInIgUHb8AKa
AHCN2qrvOy4VdSB3qA9d0nVtUX/+vcAiUeMCjQlqtyiPvWbt9owPevEQYXpz9nF5
FWoRyFAJK0lEX7tlGQAJOMdhLYrJTJz+OoYP676G1N2PC2OIki9ripgAwahRP1ND
ARKm35C7FpUAhH1eSLJCUbrvAn4+lzL4UXHxiEO5bVVPRnkB144gdOjdv+nd3qmw
7r4rcTTMnOTJB4wsz+iQUg/ilnjAD3vUJJsSIkSd4usT34kjNoB7QJiwbOyhHtO5
SJDoAjFZsmBOdirge/F10vhczgfQT2Yyx9R34POEzgoMlwLX+PP/sRkVShNbn0Pp
t8I6uE41vQ39fHFqNa38glIux+90Ej6BC6FqNjwXN76FOHS9IJZwnoO1lHAmcLLY
ayiGKtxs1D68GcvJlorUIdpmAf8HskeAEi0uOQ1P2qeLC0NK2rwqJwq64nXXWqq0
kMx4DyDrq3MOCs8c4cQjqF96UYKGPEOI7HmDnMLRKMyHgc+D89O4L9QbUXKAqYPx
MsVv6PLvQOPT1990qxjpAISOs05on65y4tRBXeV1jS1XiKWnqvRXfAnINngsAZkF
kZGmjkJTUCxxphi+ToFP/QVRj3/uO/C7bceV5nsYP2FqaTSBpexqBcoe8QSukEWE
oW2a3qdIXrnGC7Hy88SldG/xDJlhevjfJN2XOljtxY4l/GJ////5vipjVEo9224y
LLBRsI8UPsvSll0ZXpwFe/lHITABwVYUlQJXd2psJ3Pw9e3HpnS0IK2ImbrSieNm
r8gxJUjD9+Le8gRHVBr1udSOAmcwFi6aL5SO+0V57ckWXYiWW+CmlN+wUjBX53se
oQBy+aK2bYlMK1G3Yn0Azy5TKous5iBG17p52x+SxN1/pMjArwrSe2iK5Sg/u2V1
z40Af8uSRspLcBWgIc+Z2QlA8t8AfaKL29DxO6ZHKrU7ho7U34FJR8lTeUOgNluZ
16gZR9LEOUhJmlM0KQuhAToonbvW3DAh0jJJsXEWMHnRPgFwlO7fk15pbEB4LaZu
ktEqssmjhhmVY1YNpu/2tf1MFbc5BTbBklNEXn1uVZXkd4MXVb5qSLC2hVoKKBAC
JnBgnrxSNimjNkWWTYrT3M02IYEjbDTA0MBmQh7PAKXvL0cFxvDTRYrBq5v41VDv
oSKoxLhSQyXu3aBwzTa0MyiICbW0ex6GHVhrwmHuBk9tZk9xtVSgfpIEYiUpL+F+
kpJPOGEc0lmgcXJc1rUwTjgK+2hsJBLmGik1PZOWxNBij417vjr8Az7+oWDVCc86
eCPY2wJYmNQefn1aiS80TLq6l4mnjutsOFmbAm+COm+HzSyP0y84qNUAWS2pRx/+
FvASBImYDIMPXQqZeEVxziouKwPcqOgn3gCnTKiHhGLM+N0DJPHEJbOxn/OOAAR6
pYmTTjfGRdy4iebJjILekY9rux+V9JNxTG1Vq4qA2cuYUPLvPa9pq1cPRyTvP+oA
piEifHmPjISwJq5USKqHaItKGPXk6DwlnYsYVF5EGBnKnoLXPL3vhyp1G7N2bUSM
ZSdGgwMoLT3+4LDb7MLM7dCzZ6wA8g4z6nOWRnMNftQAsgiETv7BKVx6A+HnlqNE
hVPTkD97TpAzKzcTk+AIEoDKc9q79OSiua4sr9v68I7EqIseOqCgwQ34qh2IdxpI
V76QA3lT1UBi0uOyTWFWrgRpe8uKPSB9PG8uuXGMnV3lCBDAG90t8huDZRdC9OdN
z4e5qlP0oc3Ntg/Cyx5PT8mtlm0o924NmcnDEAradLdRPyQ3H1MLM/k2xrIgpSl7
11IPgeZFVvI3SbueZXrWe5dqK7vkm6wcvZSuigdef8Zkp8hhMuEwI0aZWX+IICFQ
kCT84YRQu0tmRo1+N/41cU4u2TXIkQOjkAil2ogIgB8d/Gd70sE6TUkrSHJiYGd+
GCAb8WyY7bOc2UKTx2RPeAru/1Z3S5KZ4g5Rs+jN81cH/8dfcyeidDHZZwT8LEr/
kI8MTXnQaa3RAz6rF1KN7OQBUg2bVgXhLGNPPsYoEzu+GAE12wE3saef5wXZ2qqM
2uybk1Iwgh7o77hsxLvJntLTAU9xk1Ne42EzR57AcJTK0vOHDjnMItIM92csn2AY
5HGOMLjVX3FxuvjjSp1ZbdSIYTNorIJK1mTkAAVBKybrNRA2K9gS0CQ+cQHnhQCk
cCBtOqMasYioVIdFVoBg+BVG+a74Ob4X8+G6kFh9AJynTz0Qhz2+b3HuLRF3e4+q
KUAa8Eid5p1ADRd7HQ9XXJxQZKQVo4DtGvoGNmhINL+8GAFKN2lpKhIKQsztpOgH
HF/B9dpEzTYkuCQELfLcpNUsXnG/9GlrScaQc23SYnI6dGlT8VIuxaEUcjf3jLun
uciYhkm7eIMNhbEZ1o212t2KlGG8dhrMoGc7d6m8ehs3oeX5/ObCoCdi7b+Fb7T6
r3VMGkRWixLciuApMLL7Jg45H1zN0zbD1i5FnZBhlNoJ5Izi9Z7EMziDdqvd5kpu
Is7QVgxtTdyMS6LghG1Su5MEJI/XQJAoJwEbYIZFhqhiuvcXLGrj14TLwi8pCIar
HgFO4LoRdcwu8pGpvfaKMRR+pVxq10xgUrZEkDqvVJwiQTo1f6oOGBV23NSeKyGj
cTWV/vsCe1KbgivUvtWWpp2a0lFkfa3RTNeR553AgrLbbk7txrz2WxC6shNME7VP
23WsFT+QinniOrwBkBgllHue7sFpBjs+RsFxr0lR2OrMHbQJNMlrnkbzD4XG3Pfs
ruaBo5dX16KKS9vW7ndhoiibp45NvhJGD2WU4aYPRb4nCE3Ix/FzXYqOt/ITa+qr
yfpZD4ff+zdP/a4agCbo8xViE7d9UrEepCJbHjy6RIICr0mV4d7JeleFEnQnudWw
gA3GH+LGEVXQdJw3LPgy3xq2DxnmIdlzY/JeBw2ah/QbxzSJ5RM9zepue9quhB/n
FofTWw6wfOB0MrzGmm37QogEfCc8HPE+zuGK0TR2+HtCdScmv+wvbQe4canneeev
1gdxqeHi++MmEXZqGaTqjPb4A3OVKEhQUs4VE9EjHN70KGze9xNyFjn0akjbNrat
8FMyj/lO0FeQqcmYUqBQ47A179djoQU8kb6/86xPwakZVRERzVMJtbSeqA5IMf3P
0Lyp0rZhNOiXIIoiPUEKJ25rTUlsTiFEcRiyOz1VfU/xl3e3NqtYzh7A8uecI3lv
TaifTmIwf+USZWvlwDBb1N08zUczRdnno7eMyKm63XcQjshzGX6tOAGmzvfW61To
Sh6Ss23UUKAlQfo30XIJHzVragNMIN3lQvZygqVbyKeaJBhEI6KBc1WzYNGKt3VT
d/2e0e8OHOroP+Q/RMJxpITHEiBrHFbWuS1YgDFZT27GTeCPab7dqfPSpzpDAPeW
3c0O0RWjhUCeHsKrpHjHbf1Iz01dHhuvRAT8avVpbCre+YIVUzfoyS3S/e9/4k7B
ju/ER6naiMP33PtVkKpqmAL6Xlfh9y4gFbvAt9c4CIqsGbPve3i0/G2moFZLjo7V
wtTCMa5HH/pv4+1/C7Rlq1LrGbwx0E3eeupVkUwC8OTEv8dbz8A6hdg4rtYsE+mv
Q71U17m6ReZ+yiiEjF7sN1J3FqIgIcbnQWxtulhmPChFAlP9b6St3qSVeD8A/k/m
UMWKmlqmU68uK0EzraOxz33Xylp2vRSZk+ogsuhU9oCJgTJtkRX4fTHVJ56kdW7V
GI++H2f/48DA5HOTV6wLSJaQS8chefJKodZpkGF5SpWlfxqr6DRaVRe3zH/o99d/
6KyIp0Lfyi77xbIrlQZqRcV4XRBFIpkPnffrtPYqm1L2NrguSkMgAML8X5nb6Yzo
kHC+WVCEAxPHwh1rZRoWGmUDcoBtA3as+mLBL75S1vV4+CShums+F+n3yCpL4mYR
rPrOuB89PbsWh773QMRrA4B3LzNtbwBMDXAdb+Dkbw4yKqr4bN72L2tf6buyvbZ5
CXVt7jnRfxqIrU2c2y2ffl0k8GxTWP67/ef3mNVmT/5JC8ySZbMxpjjS9LhUDd0f
JlodJthEg+cLslGcVJ22X06HDICOaAaJ2N5g9sZx8TDf7/D9aL0ZqQQrAnWRTsqI
4YfX7N5QSPkrLTVGqqEkZacYDgv9L+qhoPpuVOXX0K3KGbN5IcVguf9Hmc2deo8T
fxAVp7qK3w4P0VALOEZLWkGMAb7NNkDH0WJbLIfrUqSMDmGu6nQfqEBWIwjz4TXP
i0mxDAL4iJ/wIyU43yO9SodnGwLk5+EfbocerQ3bsYwBptGPCICN2nNOseRB0Zp9
1Y4eyDAsqDF5AI0wYAbvDraFLBy2lvK8bO89LFRN88YKEfuA6PrqE3D+T/oo4nuz
0oCDeytMwITMDRJWuUvJzz52m9elb4b8mcCQJxxduZWY4Tkbn6SA+2sxb2bO7iMz
3x6lI/silbzqb9/A4u63oqhnC5MnRPO+zLgtyi/8lM800jwuyUKQckZb1KbGcXzk
9jG0wONUXw6mIEbKGlzHgMMND2CMo52JKAydzTjHViwOvEkDYPUrcMDpOHej4zPO
e/sWV4hVtd4tJYntf9l26lO5obSzty7PJa5zcwiVsDYPDJN9pVaAc3YO0vSTyP1s
2XxngDg2qWsKnGBdgbFQFD3yCabd9v9UdbvjtjLIEZIuS+lzNSuEyeVaqGMjD9ig
j4o4KWckNPioqnFf9a+aeUdhYjI4S3bVt6SltW/bXJ46WMv2/0KTPsFuLdzD2vZU
coozi7gXJQPuHyKKpZGbry67eQiqFlOxD6OGlxji37gBx5IRZ0h+0Z92AR7gVHGc
4WCcHL8yMBoFHVz9LNNg2VUBoi4JsKyp/MOPqRsQaXRtNr2sq0cOwmWr1SHM5zVJ
H/C+bVlceeonLyjZm4LWzGRyJ9lCfVi2R57CvmYgzN2n/d7ReLfHZuIn4OPA9QYF
Lq+I0jDJi1H7XSfUaqm6yzPEQz5QElLPT6vBrirGC6PYjlW2ohxES7B+wAIx7RVO
dK9qFUxM5EvFDkOZq1MBohGGaaCM/bVCBqJ1HgBboDasju4yf5JTEmVITxq9dOC0
EbH8MOSJWTcWPSgTnxXZ5ugD1y4omHl3W6rEoJkmfyQ=
`protect end_protected