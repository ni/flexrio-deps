`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5040 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
1z1b9VGiiW9Gp7THxpOgEcynjWGi3XZIF0PEbAAePrx+arPDK9UM9Jagzz3ASATi
vLzEprmKT/bzBLuD5tSXD2sRNHBu4QubcwQmu21fIOB/CkK/wM6iIGwIFqxR6xJ8
e8YriW3nZNi4FU/q5ffiVjX3AtyhEi5pMnykOFfDvm7TURvTLdOdv++d9qZQp3HP
cQSEORHE12AowAm8AOMEXGCDxfxtC+lNCgzSifO1GPoGCre0lJQx7Kx4LDt0Lk54
oeyuvrFRW2nmPQc4G6CWdqOskeY54CYIoHqE4bVRToUaFJsPmotjd4QHFHOrDZ0q
qjGQ7V06AM1xOE+UnVJqoqcvSLh5mJ9IHeRlWzdaouXc1rYPo+m4lUzV2ACkeyUr
dAf0Fn94gYVcjfMMy3mPUcRRFUwufUXyo3Qtr+CyN8b5fEioRW08z84uCcNgpnfo
EzqR3wzdG/iXMXU7azZWfh9KlcarJjtraRIbo4wLBgq0BTTcVCPTOnqnDFjKpIrj
ZiiGRZe/q/5bJOhDrYtXtvTEkYd3cZMaH2IHyuu9FV/2lb0cBV5kU54VCqqCx3Nz
tit5AkM2miW1yisKItakOTZjsneQs+GaO6DVplCsySGlthP0wvRJ5KafrA3AbT3o
DMGy/1FxCXkV6EJGTaVeVESGhyDyeAweA93WHHVmZE7SzRtsJMzc/u7WUHoF4Vus
cse45KQjaF4CpCh+Op2ewv/TLMsE+Is/YxmlINjEc2Y5qjtIAPG6T5kTKZtBMEQt
uCLIbZcOiGgoftOf0F4ZIaYLvlPS81c95uqmzyECPAWAz6Xe27C8S+Sbom75lBTg
zjZ7Ko7Pc6jeEwuta9IBSzwhHE4Acwt0fK6nrRAJ6msqm2BdV5M4RsqKqquNi7Da
vdiPtjo8tSMF4cMilDjpZDnDPjllisbq7fJe5OFTl1JZtR+EeSvF2KTZk0F36aLF
wlT8cBZskXn3sPivR9D7toJPebbo5WlY1F9naFJF8z3mPuryLAUzEz+oN3lSWst9
NJBiniHzB+QuiogVvtSNpBVzk5/yz7rO7BJckdTpUS3sh/5pNHizUjOKYuDBMYUq
C8D5vivd8w3a+zlpGezz7jhE/6abYbBRxDOqmWsveTjubM6TTgKVuFldzxDb/zrk
AsnXqqhq70XXPlDL2buJOX7ODElV/bDJSlQSwpTzsSu4EXHibWowtYHeGVATqQMJ
a9CSZslvosa5ZxMW4Qf2K6kAWZUXMOdzFX3cSjeh6m0KjMi2cjGczGXVN4xiFeGA
WhcfoHlUy/x+0u0+U4sNWrElkmgnnsQcWB7G/6j3sLYRLrvOtr5WTXdHSVcO9MzA
lJX1fuctxp9m1oGoWP9+54JJ2pg2D74Ck1+jU1ttw4F9qY8GC7O8mJltHNQ/CnP8
yIQxSfHA00VhHIGJMpljvhSgQ3AB3mAV/RT0Owcc7Jo1d2SoE1qMfw+N69J/ykow
58vbk+3Hzn2wr/JQePKckV114csluyRaeX2N4u4/LYOyj8t05T5zTxLZUFSAtlAc
Z1AuUJoilQAP9c+SD0UhMY3sSVmmSlRGkOm34S+XSqc/Mf1GF2JJpBufCp0X5kNn
wKX2pJHTk5zY5DdhSV467z8ffskg7OWDlvQjy1sX0knTXcyF0jAqzkrif2Ljmn/6
fLGgLPsq8NZXMQyHDmQBUa4aepA+Lz4aNH5asjUlxuSf6IUCV96egS02NSGg/jmf
A9qUeca6XPvf4TuKyEwbp++DyiHAhI8/PFNc6JGoCEVXFAC990t3rvrqxgyUYAn6
Y5pgXpFKF+XQZhIAhv3XlovoCgqPo3YJWq/Qiqq8pFE8UDN7PsBPqKa05mva48sz
M13owbVeY0UIlWk48WzlGXmPr2NqVNu3wt3BA1/xd0HORFOkkxg0E63yjHNqYdpZ
krtKs8GEH+5HX3BjdYtjmUu4Kp439gzfqdPrGdWkC/ruRfYKuq7rTvusd7R09V/4
sG/tol8UtNbwqWZdND80ZVkNTK9ad2NKcilUv7W6OfF/vhm0cOM1XKiMKh7BGIM9
x/In/fsi2jbYJshXF9zUUyb2U5a5kA+Ey70DdU4Baik1TtOPnxE+EfLIl4Ve3pX7
CCTnmTkihHOuxXbLzCD5txHWKMeAXYgF4fQNYHQpUBCNRxcAwA+nwwqVgdpyO+Ib
S1rdx0IfzAsz/MB0DVxfpwBeR+KQmEIqZvOOdCzdnfTkK4zw7N2YB4ticimXKMPu
4osxN/dN9vP+/uSX5AhF+QilF+52zvppGX2cygJfAzSBKUvWtrWfaA1pDWmbdJLo
dJ81ajljnVQ4BJX2LKyL6nVflddwbnw+VT44qqvDoF0x9zpRKQCDMl77obd2oaYb
/NuzN8AhwP30bHgmQ4Snxew7yonkrpnPw4YQXHGrfxkrskgKHX5YmpG3UygHaTEn
YGA452YQSfGbYUyPNr/mU11+6p+/+/vh2I8uZEEw9H1ZrU2hkBYmWb56v06rSsXd
QthaBhFdOzfukwm0f6Dp9ZtTUHce3kOiD4eCIxDSlbSxxQP7AyBIMBWEemaaTtvB
VVjgSzI+KHSk1eAuwZ2Qvqv9HBf7JhybFJLHGXXQ2Q80WRCOuKeulhJOXMNk0QND
7xqAZ+uFsxpq6TXZMx3+WAqa6FVaLYnQgRhMdgKgCBQfzRY3OTKXELyQNE/hECP7
+huZ/RBpP83J2iJP/gSNOEu1zX4xFGfutoASZV0z1jt6TqEFwApmvmzAv2qZsaFb
XnHWoItur2D0eLicTar/KFFq0TJQT4ZQWg5IQTFiMLVvWhGLdNJprjHR5yXonaP9
Q+QZ8Z3S8POGQ0+fQJ+khU9Rn3aFxmsUKkuOZNcFIynO0vh7nIHs2fp0aYnsLtQg
1A56kn/exn6ERloepRCIiSIWG9pEFO96RSwO5EY3xwiVkno0VHh9rJXwSpwX5ggs
Lm8B3UABavVaXPhpHRqYVFV3aPKgExB9X1Qf8RM6oiVuMkU5eZAMrWPNeyMXTsME
3VWqc9n999ZABXLHE3EvAObLwsdDWo62YcT81b91DEOvSIAGilvoBvS2hyGmV2rW
glG+7eufBjUS+J1d3P6+nDWSc59rTumZbKWFLKU4pxXr1EVI+3Ok+a+Y5t1m9InU
4mn2pT/hfgmWo88DuUBhxUiAUWXC5IUr5R0JVxKlB3Xjqsv/NciMABOb12a6yje5
D49CaVzOGblBvOnUp1Wqy55BGrmTOUfZm47cQ71IPHP83PLTSfzyvftOXzTzC1OC
9iigh5ASOhD3z8mHIM9lIwYJGAew2EFncjSeyBhTiikTnps5nl9AxWxSqRet23uj
81l96VYQ3gRx9c44Sdls5aRV8lGMsZ/3hqlgf4o+aSO4dgEzAztPeCQzzicvHZD7
4f4BLZIkwJ6fAsbwn2dx2TdRF8Vdp6WgWGKRIjWBU5ieYLql8lkd7d8c4NblzDq4
n1+HoRzR1HhtrUum4ULV0mHge7Hu4CwvTgjKv3znNEqE5rpBMANbgjwrB1ffgK9G
Grl6JZtmV6ZHe1/NVshWQSszykbsSFRYdbIk1jCCq8lnYG25vmMLF2Sr8FV1RfzM
mfFHmqg/T2VKdMErLXPeL71OV3IRmTqFp2nV1Yeq03qBJEaU5b2MrbpUgJK7R/+9
Wg1pTqDUWNsbHqOfHIh95MEuJdhRaJoKNOoNmeoFXE3IVSjiRfwzr5xP+Q/pfKtc
AbQCN9paPcRmBav4Hrlpb8oeydjrCIzBF1oc6/X2y/eaHil4r+j4Xqw9hPGY8zKJ
lYdf+ytp4QwtDbeMwXKkXdt8WxmpHLNMozMeyGofSN8kaWbL3RfFn0dpwYl6Okjp
SCJu0Q7ozKhJMh9o3Q07Umu+TSGvuzX8LPoWb8cl4LsjOSAPqZzTY5C8dfDxczZE
yinhV02rc3WQkO+M4i81c/MG3sKKRlL/Uj9udtVgileGUsZLBoiiz8tE75SSIrJH
4btAMxPrEYxq6ThcutkY4Ebt2omHodAOoDEXfrKcda6M7H0AI4ESS6yY8X+QCJQ9
vQ9ZK2ZioZ9SGhSMn9GMKcmSRbB85GuJ1h3q366o7ZdR+I6A6iz9h6ifCGH0jstY
VC2kN5pdjVoqe5sXGRLJ6/uChUQ99QghyTQWA6QZENAbTnoO/Iv/n4ItaMzH/Ky2
yKSm7uXeeyDbWpp+pz9/k7MLk4ncHsNbWCsjt3CIcXppQotHmND/AxAe+ZKBDMYN
ZnPCFUNUjajGGDYr+juP7wgr12MfBAfIAkpXb5r5DPvEQ9eROOUJovFfaLyQ/uxy
VyBLbQxbmZizmMr9p7xznhDAGWvDTTpzms161dQ2KWsQYetfdOwXIrJ0d8BZqyHa
Pqx9pNGGHEgS2TYBCeyo/ei89R3UV28Yk6pdl3FRvMW8oybG0hKMEZgW+Ghndp6A
8f2kP+oVe/uHWurStEsLdRG6lv8/xR39/Dt2nCDV69O47CvJUqAFcWz0W3RV4klS
nxELvi03BTNxbY8em+z7HcmYRXR0bYH30kgUWngM8hfsnf14qsfTuPMoOdDKwgaW
/sEghK1QjCkecJ8/lL+qx8IzLT2EDL9bUfgxs3QwhpXCenVYO0yvtcGneHQDghZY
7jBLDQCTupYyWzraZbxM10bDBqsfOj/jI0pYa9qz6jZewUghsKz1l1voSNXu/Fbb
EFN7tjNdt60ncqh/1r3otq3Tgadc1fD8mj529oDA9HoqN0pYVaauzWIVmAXNWcgP
NjA5Q938ST1VAlrSZYtUoC/aTDhVhPKYIIkKAwV8GiUBAnXyZhzFlqO/TNZPSPxr
Z5tsKlyygdaNThL6beTjonMetCrXZabO2oovBsQXzfGp2M7yIBMgUURws0N+n6KN
31bcBkjhswtXyi1fZhDzh8qwxYGHtT03zlQD1GvY5yVhUlUo6keTmnb8YlwE/6NK
G9ACAW5EEBR1lYelRepmw9+8S8icrU1uOnxxH+ekMWme28oim7Diu3CgSh9BN+qh
gMQ8u6CbL3pJV/bufgzlXvOD4nSnxueEZBdN3txDz5fkNFWv+GGfbWhsX+4HF4Jg
TUMUX/J2QvM2HwpGFtr/khUa2azrqhXwoupn+Hngy5X/3/AMEA6yeEwGuxuAjEaD
wpJhpiU2Cmw/IVEJIouOkhOwbJ0Ys7u6tAVGWq5Hb62brOho2xbhuJlvCd44dikE
vrlGg4wWZ+IFR29uurYTzJRBm3P6+OK9Keg3o1awZz/jv62RFvSBkhMV/mDQxDIv
zUHpIn2DCmzJYJhkyyyrFL1hG5GGx6BMcgStTPF4Zvz8r4dj8sa3OTkQhrPMtiNg
lMEjyAyhF0rpi4zfsfuRlNkeIGt7EnLgCIVeSuD/yM7wMlnnM3drxRBxUuCkExbi
U2Wj9Q8qt+0NKuGQSy/QzIKgbFHSrjtc41EVwGyZItxMTqy6vVj47r9PPtZDDWWR
Zagiee1SkQMooNrRr3azUGXA/xzmlW0kBa2wRX6SVKMoWlyKITCFIR9Qq+IwkSgL
28U9FZJvPV5WcAzsVL4nAFrgPar8o5EDNG4h6WYT9i11k22O8DQuurOFgmS+DXUm
CV/btuoIzGrIqpDqtUFdHy+F8Pj6WzRvY9VsgWIDYaz0A7TvnoXlq6YEl26DcG7I
4r7aH8HWZ2Lc8yLwD6j9WiRv2hr6PIwyEVI3qfs/fBc0qfKtUDnAV20g1zlP0F7g
BXIC2SrI7D4FDdTVwDzJGdV/lEi/FCoQ0xx5kpITQSBnCjRYul4TlEfjF42R9zBH
sIWj/S/hNs8ounZ6Lp0ImHC7YYClJ3ygaVoTKcJCJtwEzksBaXLNGijHp4GyUiKP
8Db2Nh8u9JOxbPV4T/7i14c012uXxHRE0EVRLtaY/Vgrqiy0BjfVqWvunPNUyJ4l
LNi5FODmfzl46urZGC6pnVOe4NbknX9F9Ro2W1x2kZu6cgVKKaVW3lodJZoOTZNQ
anfQv9LBWImO2WL2YmhLv8qRCUcPPtSMrh+gJmO9V/nlzs2ZCskFjHheAYrxL3ab
jK3ZqpK8GueEtLhSZNb40GFS98uNxxFE9hAM3OCHwVCK4cCm8j4GshjwMa6h+Qf2
cRcP2v0J7u/Jadzl6qkutjlGK7Nxbfv+Y9D4ui7S3MrFwDLjZAZfcBDhLoRa0jBX
k7GEX8Swz2lD9kB43ntfcCqJB55rbAK68YibMF8NQICaZv5yMEvk4ZN9IsDZ+fdf
T1sedOUqtTi8LC4tM/LaMAB4o6B61MekQEozB+B4pjng4sExJRIKH6DYKzQ9uthP
XTjtFtAYabOOfyR5ljqDKff+ArdCOEYYt66q1coHo12sJebZazAEiVfTcxJNxZHI
qE8OQgmjCZCfJ/Z/9R30GuJ2nwcdBXYRlu4tH9LVHgb0YO9QdImatj7RMIce4t3w
IWDkFWtS2N7cOzji2pPL4Sqwn9CCFsvFSxqDd7y/fYi8BjT3h0w7eWlSxwUeIJ72
Ip8+mXyKRsxeYDNSHbrKiAhESvrSDZLtFEAUT+jVVtbZB3kISDEEzpKpsOs86Sl0
2KOuMMshNmqZwTwrvqbNAL9aFWDcxdLIHLxs8QYtX3yKIOH2G2F5Ou6Jh1EhLUUG
`protect end_protected