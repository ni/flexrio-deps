`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 22016 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
akBpHK9XojjdOyFTP3pOwiHpqpxNBldMYd8cm1NSW7E7KX7wqi7k89k8sNITmarX
pxR8YZfXqNMzme9+v7CdY0CUpZNGoRbWXod8FzysOV+LB6945Fvbw/BJ0Djt5yHP
dQUJ5IuWHsgzfvkNt8WAvcNXegxcNnbj2PiNOLnBF7RrfYrXTeU2t5U/6FTo2GXy
a1opqsnrNLx+UXEH+u54pIwX0vCY2jYlsqXzi3Uy69TXmFP3cOZ7mxmLQd2+tQ1q
T2vzH426WraASLEUo48pEPotWRz9Jlb2uxQwMLUYwi2lKdDmBlgl3nsGCx9nczdO
bXHQ9hPNCZf5X0TOEZhlE4GBzWnuZXiKAe0PcCubbe9X2B/TRff4+O6bmeNROdZx
C6iZIv3BHvzE/E9ISMJ69B9YPz6AvT36bMB4VLf+6FYyoOntlJrTVrxpbFXqLg76
3aCxttOWoS4zIQ4xJcjEKd8D05xoFUDr0AqimLso6JVVz3S//SGS9U8KHk4rFSW6
WD5BJ2LigP3jwAWrQ0EoUbI0wyYxp/JeMvuVu1FS68Bt3AO36XT56Uh9sNaULVHN
NSVbsln5D7soe+bcaAJvQOMBPb+5oJbhM0OLbXxTRUM1EYxM/hF9BZHyGgl1mQ0g
dUr+7QVMA8xw/ni6QYbU2RdNlmyFVDX3EKsdohMynpqxyp9d1CAboTYqqIo21DeI
xU3cc0mjIe9gppPlTGAPW9RfQvu/Xn2GfR/bp3D3d7jMMjvHF5xANMwi4UOXBDOF
XgcDFwZOlZkNmPzz1uBIzXu1MlIKpvF6/DKDC7Suyvr7aOGEUuUT8FczyvL9w7XA
bGwCDKyC7IbYnU63fdIlvenmnKz1LALzSt+ZVmLOqiOHfFmkQi4P52aLt8GygNjP
shj1/pzPW0GdM8N+jdPb3WBnZH7rYE3BJB16xXPeNudGQ/PXrbkrQ7LGIBgwZuA5
DX+rnIsEDCrn+o7KxBY49wb+78HJvAmpxN5TxrDo1KtAIeNY0TcDQPs1BVvE6Aet
CMi7uEuzuDrIZDBIaWtNL5l5rwCk4yWeyGK1VrR8rdV3EA1mi+Nn1HggMez0/Af3
Aq6SqwMh2K1ijWUj5jePp1Wb87BbmnX+vQzx6x+kVMnR0K4kuvzEsAtY/JKv0QEP
CHDEtwR+12DYPmOwYA8FRhpVq5j//0PXfDA002XVkD/tGboX+6Xf8FDE0RyQHbGF
Ny1v3q0xK7RL/I/ZN5/s6y9qXKNqgVBQoYhWvpV1qnUUUFUGT0JH2R6K0NtK3yiK
xbdJQMSssHea9KrdpEniUuAcpX9ogQ4jOEKPHdOnHSIQh8wjA/NML1ll0t4Gl5ph
zjm0SwGxdAqSTM2fhakwIPAQxLE0MQHosg39j813+0/k8SafBBZkOxMPEOla6R0l
MvsqOafUU/oK32rndjRAE4MojXG9WgUctA9LpmQZ1+grOwTN5s8srrq7cqs1XeAl
TD6j85Iwh8ItYaN5XHAwBy3Rt8zU8wpNfP3jAW34+pWwt+iVrA78vcRfNq1ECOvQ
h/+c+5b4ZQxjXeRLFgBGpqFkuTVL85NEpOAioFdtXUsIst5syyq9RvzjLxuFar1r
0cPjL+BDe5pPXJEgWj5EhmMFaYqgPqafwArYekRMDuSmXdSfOAlw2HeDUZK+AI7c
V8i6R6I24gVY6qd1oHsizxwd6OKo4KltbR/Ru4z9vAPhPTMLgiy/eJ5q9YVp0JQC
ToRM1itD6ioCqrtLx6a6kVhYimLf0QehmfRjencLi6K9zVZ/xpdWfdCXzR0Qo9eg
qqmze8fBfoxaVG2SqSnZ883+XejuICxRuzubUIbeqNZYdmHyf1GMb8bf1iAy7rOd
hIsOB3UnR+B+BWx1lEIFHznduHdZgzMCqQGcU9I+56J2j5MAHEVjWdFurZHkIVM/
Ps5TLKJdeBxetSNWBn2O7OjAkNcHd0cKjQywWAl/MiQHixDmzcwBGSeKBs6mLQ9I
oqV/sojt4V1QMkxaTheTZgFyqsF/sB190tswizk3L8qyB7h+8jVoDpVsm4/e3i0X
Rxud8ZcPUvMc+8xXTGgILxK0fD2vKIc882HM98SmvzvysvVu7p0gLXcaTQ7sYGt2
Wrr37S0KJkXTR6kWsTwZ51Y79WrTxG0SLwHIN9P1pp2dzIQg6PqWxzNFDynuXFhS
r8fzBNrf3OAMGb8g7Zr/yCApILQysMo2DRKITcooY23TrpgRoBk83ch2RIv12tK/
pf8Z5VtmvkkeQ/Aq3kO/YXU1HJ9DnHmMyuiQ1F318oTPNe0plwy0VIpVxmQvaZpE
PURIa0AIsZpIxcHYpeuaWYBIy3E68hNYZXfSrRO/WOvFy7cbELN1HNjbqkqce6z5
FsMdRxuLJrH3wRCYlxaBrYIrPTRLObj6MgmHlv/MXla1mlhVmPJSQ9PeTxTrJvhY
/YCpV9ENZtuLCMkzZUSSm8qosPT8P7gBTFoOC48FZpSkeVX7wQonRsmlquOx4yXg
naMB00TSCUx8A1HbBx21gecxKEHFaAqKN0dlZ8AZyVf7L+NNtFNkRrSCkJPALfv2
YuVtJIs5+6phOmkwwKgkthpfAJm1lzRkmwOejGXz7eAKUw2xxah3yf+0rOjCrX0X
3BYBzYqWTG1kQXP8dBSDRbMUHWH7EGVByShtfOKaMZrPC5h77TsK0F+jCj2KI3uW
MOehXgllROszqhoOuNSPyF4BdJ73ZbyWWq/v3JJA9LjbQiH2Zc8O9DfuEAkZzSPq
PIgtzS2hsBqUYHShL4YEm+i0A1MahpOQhe7JvWH2m/aV+uBrjpW3qClxTDgiQGEA
XK6DAdwlql+dHjCPngAwZBDmnr13981Cgj2TNR9z7laoKsTv8VWO0ZiJrr9CLGj0
Pv1Lw0e10D618+3E3+icArygOyMEaFYLJGS1ZOFE8lwAWFg1XFfVaSDS7+FgFdIN
lo0T8tNyycsiB/3TCQaHpnrq99kUPcz+9v5yeg4pkqljA/ubtIQNvDFmXJ3Rd4wK
B1/1OSaedOGjmLRO6+PM8n9099ADEw99/rKzwFhLNj0EhIInrs6KwEQ9cTIWniFE
R3S/ATJWoeuYgwF3uMMzuZFOGNB2OtDNNHS5gfFJkvI7sQtp8WYKvApiUePBScCG
UoYBTxCUwcj4Ca2oKH2sDJ5P30U6ucqy+cJ5OgL1NjzF44SaOrAzrcE1m1fntdvo
wWWck/T48fFgPt2+bh4fpKMGaoJEIJ7/f2umPVyy58RkQJ9c4OycCSrFYHzgrNTT
8xqpc8FQ3xI6aY/XpjeznyUshmZcdaFRspkHyx9lm0InJI3X8KYMfWuctc9YlTN6
sQoE3S5uDSFdBXPQr2mSO7wGP960h+Ff4IVs4N8aPwxrxF+F5eqfdeMKv9tmkFyT
TBm8UNJwjfgQ1ump6Y0/y49I8h6adVHqWSRp7ibynws0r4bxTBZnAx1h9RhQ75B8
OhooK8kDD6QnG33vh21WOM++DTxYyS1yATc14Gba8IZI3tFN9PK+4QwgG2QvE6r8
FSIGPC+7J4X9kztimYqjyDqJjVoVmoc/c4newu34dwKZ4SaH6gSm4Vcs6HDsmck9
78hoNfAl8QEToYu85GDXDbtrp04im/7VUpC4S5zIf0JzgXlMKFZC4NAFvsgYUdon
gcBrp6olsJeryP+LKNA1wWhAwhgViOj/3T/PB1yCiwyyoJ1OnZsLbLfiy2nOcmVO
hI4FKZzr3zDTl1YfPYgr+K2SMHzt6qOZCHZtc2pfACEsNnSEGnte/pai530+fgIe
qaeeZRNwk3PiTLFeB9rsE3760dJUk+gtOhLiVZJVaDd2ICV3NsdcRrLs9cXyIxJZ
zmh6xOJf+MZEPgSyxlBgvKHDrxk2jvS8jwsaeLGbrJTXviuzmNRM1Idu/zv6YBCy
qQaFejwqN1wl3rMcl4kpjw4v1w4gcThf+jrVfKtkVSSpbd9NWffgSL92svFgkwas
MAch+zmlZ7SiX+59lOzhxfOSjqrd/1r4aDGOvwR9t+DHLm2nOjprrfa8kT3tYLAf
1WGi/iJMRLMw1H4k0XnhugiOseRXjoNSa4+3tgyE+m9rNT2zv+mkr00vRteQ6XfC
2ix8PbJtwUcbLVmIg53lEPpggjqw1E/ndqQUT7HwhXJ/V0pkWodEm4pAT7eEFHnU
tYhjg6DKFALe7BH4Edg4dZumADNYEA3V+pZIOMdONWL+np8v7wv046CEV5lKd0Ye
E9GpydzU5fYwdEcqmj4gERr1RRfnnU8H3014viOrbNRp/VyI5X1aGvIZmWR0JzMu
Np3WsHWfG2q0oa0ztC5ouXyOnLdaxQun6SMONJP6m4bNBi9cf79Xd++NdHs7OPps
Mk30ZTh/xDzNDMR4whvX7rHUmR8UU7WR7DPFZarP4y1Jmcn3Foeu8gGSTG+eYYpE
SG1KyVTZSXFx6RqZxcm6g1EVsZzx0xTJGT+ncW6LaAyCUMysmishnWI9t+VLKM09
2SfyRN1DztElUiHseBC4v4t+f7X/DehNVUs+6AJTyqsq7Lq3sti81k9QjamFuHmC
PoDD8gEW1xOrSxF/Z/wIWI2wzae6S/AT/D/dvtDoMU+xmWsS+fQRqbZeMNa77XUW
srM6o2EfU9elL0gHjm0RqAVoXdz3o6QsAHi/iKD29RBkHSd0ZvsWKVK05uIQIlrd
wEYpPviTTW9P9XvrSIkjYyVw8nSHVYv6LBVvfRYb6cE+uRquPX21IykSS8Rzt+d/
Q0KbQHpjecF4/ShSOXLzQTWjOKdWn5VT2m3w36P8/l+jotYw3z3Z61GOSKTH/Get
Q6cC+EPXVDKsMURrU5TZYl0r8F3qSGrZ/8YGJRNuJAfdGNBLr107G8ajdRJLTmOm
Kmnxib3z6/OqKtUzHdkhfype283iHJAvg5f6SnZGSsKHQRKDPDr5hteq0OGUZCbh
Bmjimx1WFzIH5R4SJJz9RVcvjT/Fxu+4PQr8qlcfB6TfuO5JYDK+Si5ZvLExnCCr
P6wvfS4ZNWxJ3jBzjM/mSMqZDbdh2XvDP9VrBJeAMvlMnGX6drLDZ9Q65P0b/FzN
9RVoWPy1YjK5lnkOQTJhcX3ltSh4yfTa04tFE1LGerjDjv3k/AmmIKomVzmA4uVN
L56v1oy1iQ5/oyXg8jgOsRJ0meputkpXy1Q8icipytK+7qWzCERa/Vy3lIpFmM+/
Iqx38/ytxlk9vtrKBKeeqd70k7NKwG8jlMchuNNQT9K94Y42JrA3dZB7xuzE3ndr
kj09v0e5MId2TCT4yGYeYeU0oo/UdiiDRYuMrwP6gf2qGPffjGywyAKZxx8Rl+g/
rOLHT3o44wA0g+J/3p0EXQWBAmf9bBoQ5XRn1bHmRA/yo74ByrEXaoDI27vh4ZPO
DkNFafF9p4RLpVwpO4m/4cNsaj7LWq9lYjs9maGS6qoNWdUk1pwz7OAbBSIQaXuE
JKZhDD0gWqlF/7+Hpt5xH7YOsJqwfnYVw7kmxRD8gyB/VxLtceWHM8b47jqkE7nj
L5DhNRD7P0kk8AhzXR4l4Yh+TraFn/PFgs8eypGeM7EZh9frUJ9JJ0MqT/2EDqYN
1FXX2TSPpjDmOYFL7ocW9paEmCCOS4Gf3OcmnJeIroD0SZrSSHfqQQas/kE0jXna
nX3YaamJzp+Dru4EeLdtL7h2kwty2iH4TVbvUKFH/aKak+Ef/sQIscmp1igGcB35
QhbUQjWtpTvu3+xX84aVSpnLDIMSS2rWjpuKSMwVURc0K5mXp5EQxHsCFNewrtHR
uC9tj9SgeBfItiIM78EtymXW2S9NWD1Uo6IQSb+cwYWC9kcYSR0pylEGKgqmaFGZ
MLK3G+OeA6sOiQ39wfeW42QkRoRhHnr/py0ZlU0rDQo1+XNTTzNrufugtoDpUZY/
6++XgNPFWVFw1qXMY9REYkaY/mIgdaqdhDt2kq7BqrGNQsjWbUd+aRvg/hrZkogs
Ys2JGuvCnRGg1tb4F18dW6qIk/xM9pGmBjy8HdsAGLT1GdESuOPb/1+P6glmF3Na
q8o7LE+/o7Z2EF290eAEe29zGFevAUrzWPGOcMLQvoTP0fUUDJjkzvZFNY5nFHfO
Ql7bZ3qeNznFvQJnGHdYF5B6LqVKfK3vBBTaaG2CciI/uJNUNhBVgerTsELdwDgA
ZAGL4NPARtSQRuENJjAY4In7ru0sasBdbsSX03MnM+wv+iZqdicAS4waPVOtPTR2
DaPK7H424ZTd7reDt4lbA6LjgGiRsjt9IJ2l4d7IExdoWM6QSBURNNO/nrWn//Om
DRb9BbPhZzrj3gyFBaVwUT3DZUsDExBhF7HKmYQcO8v3kYIKe8nzSDVsXIA61geF
Gq0VBnGcHGR4A8+pNebefFeP/OhT4HPW7gFVqK6iDvDoZW4PGRDZznndqCy3eL/5
pgdVf3qMYrNSbsXIzzDxPTTApQo10//9ty/yan1nhNe9ZJtAQH7E9Ys2sNYcKFnO
JMu9yA8EFyhiXCUeQ1zanq4yrx/G3JKYGJv5dqWdY48x5h7t5hYRIykL3easu7Sp
Ui+KYK71+dF62XAuP3vWi6aXEUXdoqC1wkiOc12tTcRpbGcZBYZXA26sjeLBWtnl
6qM3k3b26Nfv5Lj8V5asSQ+7Iq2vqj0ky+EigqNbZ+uQ4M7chZw+GOb1HV9kkwp8
STuX9/5Yc3dyuXwymqbbCWJxb4QbQ8eiG9tzqtDWvRVrJrmwznzsNh1jdzbEXNCK
epGSElv9aISPaQ/WqHCWEkJJq2DGS2RAAbpn0lqCDcpHUu8JuHJYCx6lTVi1M1yc
Si80yX6dmat6KIfuEoNWT1ZUoaAQctcE0d/T/f9NMrRK8jY0Z/vq9JEJePafcqaA
2OPresxZfBjumNp+Ea/5MZArpDuo/Ewuu0yYeexHgjywW09RE3MI3CasPzgfaDCh
84gE2gjceVqfOLtunr8QnvSq8hCzATqEK40Mibm6RxO+b4zi5t93yq2U7Xrh04PE
cU3ewGBgXR73w+Eg8X4dAvejIWsah1dlt9ICZYoxuZD822aiG4CaocK7etK5lGwj
+zPDRgnh6FQ9hycsyyr1cUrbQPXWvucG7RfSB32QlegOD4l3STMRc/Lq8RelQDQM
yKTiwAMn+OGELRVBiQqvEEVUrsTvg+5+27JPkB1OtB+FPoMPOG7cz7PycrzcyTp7
DcpQWZL95hFoZt2SIetXuattLN5T7GRJrhCh/VHe8ZSgHidKaDknpiFt1eIpQnii
U49noCnkplGTduoBn2AMr9HtM7VoHN/7pafgMd4c+BPIVGSwuBpqCBdianMh6WLo
34VXz/i2Ghte4wVVczjSHK/LAORrdYXcTEvMcDgWZKTKHi/rauhUwiJO8+xTxb2H
V+cZP2+QinMmnkGwUOA/omyv1DpGYHH/QG7KqakVET7AeHa/+9i3rmuVYkf9h3zV
l7C0OuSFSiJJJPqOr6KnB7MILMJ4XVv2x8/WNl4jzeZjz//UEgeAHKK0krssC60+
y2P5ulUhZNJ4o5jtkFr5lKDqPsPLa+866aqa0vUaxHDdkJr8e3VXHNmztHc4mr50
gVqNbO4pSw4Bbp0/ebJhXNxlA59oRvQgSn4JjbC4+4ukafDYH21HNWoxgxRqp5+i
5pa6pe2PqPS4hb8MIIqUC8rrU3RTLwH7YzPD/0z7HtZflSx5vqBMiSAiwjP6yIHi
Pm62px/5V20YK/4gAbvFNXg/obl1ButNhqLLoENohj485fCLs2cnd48h240jVLP3
Aw4OkFWxY2K4H6Cua0PvgDNd02lHTk6vlS9QSvtGLQcOYs6VWtuyg28eJrVcwPwQ
Xhby5t9Uig1kNH+8KLrk75aoExhfbnOEt9GdiaXKHbGzvfvTu9xo+IjHZ2fwBeSL
EYcllMNUkKa90pGP2hrQ3d4AuXHJcoCXRKxI1plCnvLcVDjNSeU4g4ZygUp1mPU2
DpTL7cpSMTm/RM5u8VfrA991gySCcXOWOLP1HRq06yOT8eyNOMgZZdGa0gZWQ+7f
0FrPCrEOIAgq2t/NkYMkgGin+7DgZTVxde/c8dFyZoiIHw9oojiRTzNz021pYLXT
NWh6yjPiuhlgrw1vS1X+DsuupZyE1CJXAPNgXIzV+Ew85nPk3t4EGGgwG7Q/AK9q
YU7+7ZhBYgLg0yCEvAj6J78bM83y8eBBic41FuqdL5TVBZMFd/5TLaMcvQiFB0zI
MmoiBNGQpsoCqJGWxN0pChjCA5hmIlkOYM78ptP0i+oTsoQYil+6zFK8D5LZNn/Q
H7QObx7VBOFKCQovGDNLcR94aiYICDFNeSJEtcUw+tx8wu20ASiSXHtQXLn1y0S/
Rw2x7QaHgopY4YITWKQlmsQ/YNDsmH7aW/+fCH2Fig3Ojx5jbXAfokmFLXi1qylv
YNJOpMMWvV8zaBfudtFN+K++NUZib3QFkLWb2QLmttilSpw0CqZB0ZAih/6lIZIx
MC2heG0yQDZ8Uvq5XXTCBO9T3EHwynrYA5i/ssyu2Ex/Ws0dA9Hsn3SbPLlJWv04
AldAj4Ej/STxC1GydFaPLYTfnn1/p/ehqAaR/GPEzciJYwjGNtQoSvDqAwsHNhl9
HgI+9TP49EUVfcsHOyTUfxe/4vFDe9dzSF5VaNAOLaocyxy5ZQPXKz2P0rHAukud
hlV9MDyyf0hjuQ01wVtQuvQwH4sZrcVgU4g95UJXpfsNn2eYoS2MbRl1a+gG5g2/
lJRBHqUpe+796uTiqA95dMCYwDyQw624O+LDgtFjNyx219FZPUWdN2beWY0HR57W
xRCk0UOM7Bsm1rGz+xkiMDvl28KPT1qSHrbH1LruhkcO+DQ5hdmEHYEuMfW5WXeb
/AFOE/5N3xDBkF0D6g23u193TH7ucf/6V82X94mUWXMx6DKYb/JbtNVpfVqfhS8E
F8YRIMxpFR/oLCSVMVEAd5koDGhuv5uJG3fQL44za0RkOURqOBGblYEuPmwkV0I1
nGzPL10sMeGW1WxT54GQEUXyOTyNLSrKxFR3GhmXKAEMJNO8LBppxKrgK7F+oA86
lpiAHxdEBI3Osve2dvx3La1lQvwtudAdV33pCUSU97aW31CSL5vm3DJWMK5OICXe
mkwaqvDRibmlzKgmG5JpftSfuKV5e8KsTs7+goiaHFHQ71WRl5ZtUvhOEQpV0oMs
1dwbnLYjC83yPyTjlXji6b/2+d0CtOh3FAiJgdJKfHoEnjoYHNSNysbPEc23aKWO
BewhfzWL/fdqArQQhtg8XFYuokqSUrTmuv6FE1ihARmAHpy/X1oqK6FJXsfAAG8b
Kn03NGpFk34wMyy0x20ODQ3d6DV0LnXi/4tt2P5IwOD0Nk7W/7K4Ialr6GEyfMpd
0zYXpf/lYCnEjaz1abLGWM4pMLugiX5izLUAqXE2ieEpcek3GxhKvV2zyOHXHS/0
LNsm5z5Zm30KdsCkUOccII0VMqqMX4oJ3D3PZs8vrqJyJbJax4j4nRMYcfPRuF6a
0FvhjtDbv846lgpMVllM0dUO52EL/hEwrcHrqAEzWkquDHoTXcbEpClk6d9zqgTv
Eoi+bVQKFYcxVOc2nVzzLxubaF8xy0iPkA56+1vAPiFJTlp4Vc7Iq9Oxgj7en0jh
KnyNdtM2K4YR2HEX4Ka1di62C5lBHm7uqKGcD4STP10PxZ6ghc0SaYmZyXPvSUsn
vriHD0jd8usZQeU9xCfgL8xcW2vsbbaZj2ZXWvhS4f+NJND/mMbTZsYivuOXPe/y
I6ArQWWqxOcagQdfRpUF0DTgimoNVdtwcRKPPIGC4mnss2kerv4HwYXFZT6LzbVT
RolzkQpXLcp6XEoein9vo4AP52zvFZ/TT9eWXC/n3b0tI9HRUTUhq4ZSrnV1cA8U
i4na9CzkhU3L75i97FfjkYNY/W8h8LGSYWq7whPysl6OH8aLm6ktrQqQCdDmd+IR
KiIHQ11ZdoSFk7ph8JGVX5TErlr1kUJ3a3D/Z64vWeif4p84ipdjzussE5c5/5x3
y+1zvBZg7th0vKLhwoiOHGj+n8qLTecyfy3nm1PFTGDljpxZWXgSW2FhCsSDMcCg
T1cv1uyr+T/ktFLrW6Fc7A9qLw9up3TyLuDpc8uteCg+cEg5njYjDpUiYRlWgoIY
CVde/iSub51BkKZG5ZWm8yJogxqA5dlnM0SbLjU8HNka2FL2+vIYXr34bE2ivJjI
woMeZMGG0hj15X4dc0FSccs9nm7wVMFGrqCdY+VeGj9gSL6SGhYmRCW0HxZIAK+I
/oO+TXPTS7v+rST5GaHDV7M2cZVe7F2fTi5KgmgfDK+lQQXEzS2LqVWWlE3YM8eV
s9zJ12l0PqKpd1VTkhh8EMV+ECSnZ4s+5NDFlFsoHxSD3ilac2IRcXtDil0Tjo++
7kT+c7uIj2zEPqdwOiq9lZDXtVbgXt0J8JZDxfJ4nJ550Ki8HieZ2BhRybuPTddi
aIIJM9KNLebso1Vp1TAeGTnPFKrHgNdbhvmtnrQvQbqUB6EJahq2hD9PNmnxuvG2
2+ttw8pa3HBhLiuT0viax2DWhOUhrIZM7+wU9gQGnJZqaY7/qMwFBdsBUx/SJVO7
qSzvGs5cgRyfTKg4WlmsI1SFOF8dPN+iCeiXljvSwGxfc13aSgPtABZcm6ZHYY5D
wpOSf9jlWxvVmq03kq1ny8cjU9ftamQRpYPTm0EPACtDcGhemFaUxTdhtCLU4iCJ
bJbronOvkY23TGk6+MOsv3ihX8Xz7YTm7EcO4z3Fzg3DtK0hVjn4VgQaMCvhhV+l
LuoeIl3QSM1a/0oXcXUcf/5md2t/HoVaN1leWs0V92TEWAzrxRPboW/BY36j8aQf
0aF2inE33yvWhohNNQCIv3RO4rl0EOaVF/qI/YWeFJlW6f9M4ZwHryNYL6pHyOxw
c84cY/vwJwv6XKp5lPFnBJVl2KR4iZelkQWb5Db/xjHVWH+ElJRF4uyQiVEAbpiU
bIpjxB7UWKdcMLVtR9tFcTc5X6jGX7ndes/0w/qrdXgK7h+6pec/1WQsZ1JoTi3N
gZnwQV1CPdAi/7fJZx2atHw3WbPq2NVfQ2roJ+2v6K+20BhNxTf5vs6RiTaW5G7g
Pi17njJ+QAlUT/9c990mNLCwyxzrJPTU1API1nZXBoUbUngUqOw5kvcFWyCgZF4G
6gT/sLRbxGsa5T0Drh8ptZcP59dzk0owhnqsLuXdM30e/Tb5vi3Cm2Xoa12x6EDP
GLvk7VjFw1IpC2D7a6Aw3Xixc7Ntc7rWD0Gi4QYWD2jMv+E77H0Bag/p4XCZo/7d
fORd6TW9ivlY+2vUIPH3dogLnLU3vfL+a+zAZHVHBkr6xfFmQYlrH5lh+Eue2wzs
erv/CpZDRksBRqDG9fSjiSiLbIKLCYz9C2OqeT/kG01gU8l5In/G8LBrGGEVqz72
BPSLnjAAqdnFIFKETIWBpXINVEGJlfgOQ3y0N6uLulr8L69lpA51W6QO7lliKLhR
ZsS9XHeOuF+qawgWcKtjV2ojuMcd2hFrlGcpricnttNedM5bxy3C9hZjaB3th5Q0
19TGm97J4OAsH3Wnoo+K/wRVncpYi+TSPKUC302+QxIMRJTxYtTbLRasqeJZyiV2
vcszav7ayUl9LUgoYy4B5b2IH+Wm4YLi91cp5YgnI4DacyXSVpQPlD1/ZuIvSb66
EU2NmXigwzr5Pw56XGYup/NXPyMZlLUEYF0/XFBuqkJOJAju68pI5RjpkYBlKYbA
dVns0N8uzLOmW6C5+Zzgan/e/DvHcnX/1VtvD90QepX4gKnTYIL5s73y51Y5nkus
V0MKLX1orQhcVUVkt60VRwLbHi3lDE/9KKhdbQsqmjJ+BOsVCZogPotKsR7p9rcL
oIJs9e7S5t6sUz8nyu/P3Cc8KUJDpFbwE1psKzqnD4ZMYhTvWWmwY+KDfw4+q7Pr
O6uMFSGECygHJyEIPoO6lyhHotOPvAb4NrrFLOjBTWC3n1VWcpMkzsq/c4hmLBsd
gtjAwoZ8Ledzqs1IPp2F3LfgS0R3JnJ0UJVwkKxeioxa3vl8/eOPMgLNt4QLbc4u
66mKQYpc8bo9Lbh5gxgjF0sK9I/URhZE8F9GYRzH7qAX2KHFfoH/TXyp46QPtUFY
oMr9y8GgYU5Ra8RM8z6nuquI6OsfFUzhB74MiwQI9zB6CiqrNawDZyOnWSthKp39
nZeThuC9OKAPrTGS8LVNpcUGGKIeoGLFKq5qlyx4xEPeSPhTSpHSzj8BD+ASXy3p
0rxd8ej7DlDOEi8jc+bGoOpdHoV31DeQ0E45ubVeHIHs08uhqX0Oz25VEBTKWONq
ivv/ok1EzwvbhsHmF7hsqvkdjbuJNi1Xs+HdT3tlF792ct5yTOpFsYaxFbSHZtu4
0t5nDQfNytSjWn3dimUZWD4vuG/7GNiafxZ10uckGyPx67EyCjM+T1pJcRRV2haG
so6tTOrD4ML5IGwHEkja0cID0WOxW+DjaIP3iGSN4sUrS12zz4dlbP+7MbPe38HA
K0rmoysnb2caPsjUBkk4tNxpqQNvDwKs6biwr8KiGjS/0XEvE4eQ5xj+pULGofsY
Qcr7C2JsvzBVCPz715a7DCBlPC0oIJb1ACBBlZCpractwy5nFmV/LxK6r7UmI72x
r2x8Wc9+SmGChnz9YYq9Fo7ijlQIeJ6sJEbnO4x5iSKcIONHn25UPFOn3bs0GeYM
ej9z75erDklS9x214Y7mbFiPXocbx0sWD7HiyIKl3VpGtPfLziXUzluzDLliKbaM
uyZYAbZVNRxIXhVassr52Qv9MwmYKl/EpjJcqgx2b+jYv2v29OcuzkP+2yXwxvXl
EY2cRPnWz15fB8xKGNX45J0Vz/KSPZ5a6QeD64nQhSIv9Be11iYoSmReU5qp5zlM
/4Q8XEukVKTXxv9A/8sVa6r3OB2amzWD20UZjteYsXFAH5fqiltTb7vPcpXS4X+u
TYLfO6qfE+e+VCixEgUU7H3R3EL2GxSuH+DByya+rUfCvk+uM1cn5RmpbYO7Mjzd
Ystw7BwHvLq/lCOXb+JxVbqLPX4atRmra4cfhue49pGRjhswqvw0mWBODLfZyvoZ
fbdZTa1xy1QjBO20uh3xrmXejJImJXr7IDzYOOVbnJPHM1S3F0MFxGsU1qtocn80
ZSvo8wlHGsS/sp2+DR0EUCPYM625Zyx5cejhh8azYw0A3RqWg6Qvgb+r71v1WlSd
GqTexAT3FdphM69xe0m+svisYd6chWDEONQengIQeaExngKqpyxUtWe6FfMq75Ys
ktmKw+iFppn9iFltcTZIbWq2wI7fKtiBigLahTlXpnGKb+QbS6QDiUQV3icf5OPO
Vx1l4bhEGq3jWXEHdWcVE2UoFQdrZLhCX6iuFRLapTuIyhXDlg5bU/EBX89QBCcQ
/fpQLSYLlPS7KtdNQvPjj7/X0GroYeNo99w01Y5HUs8JkeBcQmknn64DRWfx/p/7
IjIAhOZ5lXfWf0rwXmxf93O6ap4mFjSaVqYjDqJ6BhDj2/ODokFBV/3lVHklkI3b
QnIx2VkSmHl8++r0f5leKsdZ4up7AwokGkTscenG9TLqmGIIhsjg78Oj4159ow4l
mmEEP+YldG3OhmSy9HEw6XnUQjxyA4QUcp7scYxBoIaCUMXLxy5v8ypCeUt577Ji
64Z8ZURuBbbzvtVmg7DwAOVAdjyPUAoxuspeZ5E6siUdyRiMIdZ73Hp3HrR2vhlY
Q68WNuQDoRT6krbfaIzdyDEmRJDAWYiGygWtJI6ocDVaxBoSogVQIacSc2zzGBY7
Fk5nHjFCRfPtmzY/bw0fuM5xw7z2dR8Z51fADj3N65BW1a8kAsSbpolqkTDGNfih
QTmZ54kMv8p6X3yVhv4stROlQGhbOooH7FQnpkwgjClmXT5ZbHT89gD1t2xZYBQW
/Ccnm49ipksHez1h2Fq4jMmeZeRoX08GEvMeuxRKFZdSUeOe3AEZaaPTgqv2t/nW
wHE5B+38CvvYRozOXycQpYUN5tRfy/6vKsn3oc8k/q9CquRcnULCp4+1srrg0ZLl
fCM20iJs2JxX+zpfEcxZpLfTCXntTvBa7bvv9+jNmagwXpBEFz/Z8cT4eT6rj5En
dRdvocEjrXykL4cgWsTcQ+WnC1I4orsteLPB0zr3ushdaUAYhy+icH8zmrjUHi61
zsHusr0PPYs/7Bftz6kZcJMaSKrvGwSHB2nOv7H5ZvppMrl0kRAcD/ZHaztWKvfk
zzrvvoGZvX68SC5IjZpyAgBasgBZ1KM/XsZbfQxkIw/Uz2LDq43/EvzvIZQdexSl
GWShN5xVAMDVu6PTWE3Kkd1SroF8UQgH8w3SlWiLopZ1osQ7qe2i5IHtDdHY5OEX
se4ehBLYZQjijCp8EsW3YkSZq3GHUVByq1uXWlTVKzFitZ88al4VhvIWE3rLnWig
w3bN851WZ4nTwURAHAK+E/fSV8Vj0IPog5rSJDvgbl8XAxtt4voIt9JfFbvAtcDV
Uh07DpwYLH5r1xXu53U+bJYDfla80WH8vYNwhp99HwZnmvmPelPkJYLIe23+ozvL
7NtCBlDRtuJloLHh0M4KS08zleHZqeu+wKqbY//XVcMXZdQ3bxBkdprWTN8d3lfM
hEV05SAaQDR0D3R7JpuX6/alnl6Js6eXhjEIXwtLyf3ddkBN1G8ztmge6YMs4QL4
50Jy7IoQ+Alfwem61OMwUWe7aYRbg1qEafrNSTRVlrdUvopB4DrYg32a38CLjk1N
SJujUewf5JDCO7bqpJ+RmVVwHEAOygQMsK9yIvn03d+hFVO0SKAPv7vCEN07fVTS
Sc17X2+1y+G9R0TQjU3ULMHRgWGQ8dS3eG/H3c68FfYPFCUcJRDUoBzqzOrMv0ph
FAuUBDIeu3Ff8eC9xTL7Y7yWNaCX6GKz0aFJamIhNh/e4cJFp7AqVHzYL+E1RsjP
DJQncbd2MZDmb9hSKbTT0RQkNCkqf1XuZCAlIzarsFWi43oJ4k0huWucZm/HgvlV
XIj542sRj4C1HLGV1NPSbi8veReMgtHYE6rI9Wk4c1/jOtZaGNq+8zNfHwFEmz/B
JXkWtKjkgSaFHOAXC6X3nePMmG005HpzpuNpwo1Zo+Nj8YsB30aw2s1b6ETD57xM
e/kjrMU6JAVwLuwkktZfACMIBwx8aaQ4XFSl1vbB4B8HZv73+gFVDxBgPIqVKrEm
acoA2F4APEwTTtyXlJO05eOqzHsF8bCYeub/oF8vqvtif4NGPdSy2324aPaHD6Rm
B1ouPTPs38VIVGxTEkWKy+B+miWLWdpIh6B8lx4kzBm/GKIvY6YqLX3c/26E/MQy
MRONC44HUXnk+Xi8k/06scwzjW2E4RvqpzPMnp0JNl9V5Vy1RZbgoafXlSGsmGFN
LyO4hFZsIhakU3KBrIRFamgonLhIb2bsyyZ7+Q+Fm6LM8/wM3r1lUKe9F7zJE/FW
94XIL+85laI4eysIhBCTozPoX9BOtkykZd1hXs9G/0dS2NhO9nB9Czev00OOImcz
IFYbKJFFucgdQ39pJAv5Vk47oO1TRCNL8JA7bEI9wlk6zbkBMHlMjK4jdJp53gan
9R2NVQmi8WrP0319kSYowBIKxBwcHGYCLa0Wax3RkBDOzN6P+zWIU0zwx9oBVbhj
L88VUMcWpS2X1QrSCYXimkr7lZ5FrR+NANRtIW0q430XiNL0LRE/prkur2AL6LfB
4pmUyNh8evSTa0k2Bn/lqNih2F93enH6o0gYPlmhB1DDY1/74iWir9fr28dJG04r
HvhqVx8vVfe53XKJ/SbouCA8Gkj+Nc7YAwneqBhrEf1lDlrpDXHdiRDhdzVVIg3l
rzAk7hnujIUj+TnjpcM1tmkueMZIuS8RNHsEqZEgpbYcYtvofFFOzPx+hr69i/2k
TB1aVkFK1pV7okEJaNiFnmmI99dXQnuIjrrePNNAUM2tI93hmo96bseW8Ts+JZWE
r/zAo6wkM9LGdzInvIrQBe6/CRQILHvqSWLoXR1aniKQOUec5XvhNSE5/g3pDojJ
O8KnsQl5kKha+W5L5opS/QVmrx3JpkeX8/VJPCSdPodJNhc/DtBxltP8WFhGgsTy
r25bmA91zXmK6Rht+vTlgElYMZUuBKKLG+/CEdaR+MQoOsVj+7aW4jvUA495mCfL
P/rlphWgmp9xlLCzR+Qqutw/heVyFYALEeIKbpYnN/5uFVbxZMmcCCSIyzvY1LWs
7qdbwAuXty4VRfQRGDInlNfqFhCoJFjhGH7GnTXDHdA4Ab61BM97OKIG4K1kbC2C
bTflCy5AQn7MMqiZzGSzmDTu7gwkI3oSwvVoPlzw/8I2jcVpkuR7El07vbYo7nez
EBN7AYioG2gStvnW0MCJKxfHwpn3sdXhXjttML1AEp4qjCxfHK55ie7qClPOfFAK
BS37Fm2sBxNYs+86TYsVdFzMwavxWQ/PegobH6k84K474IIsjO4Ipd8gqUxooLmR
pyCAvkQjaj7zQcSS0LKr28VxAffvoApyVWGqSelp4ZN3hXJz7ECsuK9rtW6zCTlR
ITSNkFBHvWfP3VFRl3kVgM1f2PHqnZ04JtZkGsvfdzBRBDUtIzURp1inKJyXX3tv
MBY84d72oCcQCu1cMLdiw6ex3xa7ge7qTzp3ULLx8wvk2nQWyXF7tuWo8EfTJxP+
lX+8NWa6vD0nduS5dBI9N7Bhr3sE1qPzsfP6MnmxlwDpr2MLguRi4W7dJi+Sd369
4ardHMeouVBIWV0Qh4Qebz6eKye8oe5Wmo6xZ5rJOkx2lNqAuY2wdNHoo5TpY9Vi
dE+Vkr6UcQNlfN3y9j4EMJC54KF/WkxhMdfbowJbM/0sWS9L8r9sqiK7P6KXRNTt
7sgFu+2t8qA8krOq87SVcr242u3XKLvRfQ+MAhh7NlZh6F2E6UMYdTts/AhVgUZO
xgL2NlsSzgVBr95N9BCAUSGHY2ZvoACg7qWEBBYp9RfFyQCYwH/hYHA5YFuE3VJ5
5UyrwsuzlYeoW+OPYNYpdywIMport2nGFe6buXHippcNQ4XdMMgVArEIKvrWgRLE
VIFKugZ8d1bp1Cg9RKJugV6kI43gTIfFnGu1Wi2KK8tcptt57szggCvnkKZn8LUA
un+aGJhNAy/1wC2jMS+TYfZ2tOeBozj23GzoO9rVamCdSyslh00+goWL/OMpQkC6
KDw1+R9ZCL00h1phA9Br2eN/FDBTt6MidKTfeus0m7p08Wfk8pX8uLCaIH71Om79
CkyfAWRt8bB7N6wp+NUMibdP7N8FRRnRvCyc/98WbDS55HDeigZmnnRH5dkPgP7j
RjrR7YC5g5+P58m7Ns0fAoK9xudzMUhmyQQKOZf0fz5PDEJ5qVHPjgu8ny4idAgv
+c04Fgm7Y0e9tYImajso+y55Ya/6snbi0njYa3Ohrjj3KKvXFcs/AWxcSVb+9rdS
4e0Az2onw7WHy1m29pg1PZravhK8JtrUys0wxFtZ+B2ehabMAPmilpNSKG+hN2HL
xJi7jiZpYZSqT20SkOWey4/nuos6Q19sBRodDS6zR11JnT1op2P77MTu/ItwMiHH
2QrXnR8NBDSGxEMiIExam7gwVlRVRH1gr0cN78negU1K9lzZffa4dTyzuI1I7p0j
Sw4O/LyZ9xIuojIb4q9/JnBo2Jyjlg8gexdYgjPDMcZPpgDrYiuys3tLcQUiAGu8
bRzroAaUgwB4vytnnWmtWQcjphYVm02AHbrK1BDmTIXSOMv0TOKpTCfaXFa9EkMG
c5Zc49MwNd0ueyteF70J2AYf4BlT10GDrW8JdopdVvCkye5cuwlhhpGtstAjTJAe
vEooIaDGDhEi4PJC5BFwA/k8MgVKPrXJzyc0aAOJa0+1QRHDt7jnb4iXVAPEYfyF
HCrNRiXyuTTNZgW33LKcPxUizWRFgcIMNDvE2dGTX9WnTIYazlcBny7RnokDaT//
pSU3ayUouTJ9th77z2iX0eOmwdSjqc3XTxqzLvuLXBuyKcKSOX6IsGFdYK4BBUob
V0O7qBlMnb2w4x0uBdD168FRSDGTdidcNro8eCiqYnkuouQ+A46PeusFJVeWCeox
geAY+NQReV5jPlQLAjtQwR0lNyH/ivF5EgNzq32nZ6XH9Jcmn9nr9W/7GdhNDmLI
XWcz8XrJOndx8GESmj2ZVmnM6LeRXDHVO9hrqQiVe1KMsri7sqNrjRYGCXCnB4RC
WN59Suso8tP0F4QIIzc/M9LnA/EKpZ30ieCy4TGR87riMDkLhaiLkDIEhKGQjZBS
CAq+/MMmr0wnorBfBjsRPMl7FeFlhZX7VnebBHprkZ62Xy+EcSNlg0ezzTL4s01l
Jbz2m3W18zR6C2LpfNHHfq4giGe52I3u7NLKqs9TiMyS5ZCoZG9Zf1xaPG9jg4Ah
9QXZ5C5MDPRmZe08VtNa8A+PDPozOzMrI7XM9TJsmoBMvwJMWw0UBnLchiSvKwZw
JkwC5lpLOciHPgF6fA1t0YqwY1Ao3KxB505e0d9LYqUmjZYOzghThLQxhSfohmMz
2S0lj7KeS6WLsHix+9DvjFt1h41fzeR+Vii71U+0Z1g/REvQLNtgDHrNuLHzIGiT
dCAaBeDKfDbAnqw0mK9E7GxmCYFms97TwDRbTt7WLN+JWmw92drfVojtIALB1WfQ
R8vfYkqMn8pVPXf/hjJQpggZF+CAjBjDA+mPnnuKDpoubbToFsWkkcmZO/c/+/Rg
8NDpgMd8+j6MLP/bWwTl8kT2hKLlclSawDuOzIAksbxtHzrRy/RBAA+ZqfhQDAIK
5PTy2rb8A8LKFI3jqYP2VWIQ8GGur/1N4/lLUw5I82CWzOAESqSVuNQVuysKgCa0
Ce5bOPW4ZfSZZNENlsNrmn39BJPz7/bet2KmvigXNy8GZ/T8tF38nlB48IshnkFv
S84Plb5dbdXz+sEUG64MFNM+LJuMyWSz71DRObIi3Es+0TgdHprj+VllKErhtxwt
kbV3AYtSvdEfAORbz4qoAT8EdYD7abljanwuWVw2YTtDHqMtiSjplPSGm+4Pqeym
tZ8RiGzAelgPf+p7Pi5F3zCgkAvGvWTI1uLDJwlTNewbQO2gw9eb/eRA1WBFPFGB
xltrtiAGvg266rSvJLeaoXBhvhsqpB/52A05/mAFnsxGbtf/AsZzvuND+u/JFsfb
/mfiM9mdBkFTdP532fgmFSiG4Uxwrc2kEuFBmVrLrR9WH0MZPlSh08XldjFC5jb/
SqF4DRvUl6N/YiBaFCBtfluaLzqLYgbPH7Ve+OSei+6hDl2Xg9BiBQbkKT36idDA
xetmTOILtxWoCXXhCn15xf81ztHkhxxO/yZGch+vq1QPijERdLOT+lUCHVoWgnBr
Xs3+31J22Xjz27BtezOh6NH9qC7lofLe1IY6cdKlKOvRl7HvFvIF16X4VkJQwZoQ
w/tylyQdJpf0jXMGnsBUeZ1LbdYeK8ApBUOjgaaLe+eYzCpj7oJIkQcTxz8EDy5n
p+vdPC3C/ze9ASXkNymd/3gdUasumGvGmTQu8YWVMs/EepdBV4BpHzsXjKSityHW
qQ3XGbg+yyiIyBPus6TcAE570OnxiCGfe3HTMVsiUztWFlyDoXGolbka2QZhfSUy
dWUidFyXDKxlwovvs18MsK2z3tMkjSKIj1Pc7yrg8m61qFjbTT4DwKGBKm4F3q/g
GsT17W/gK/BctMcF29sREXs9jt4ndA3wjD6ga3r3OuYhvKoBdSREHWFHAaLTKxRg
mdcXgNoTG2okJ5mSOJyPUAyzhUpiCxU83maOoRIEZ/3IEe2jgrpL64pAPQLkZNyN
TNVJ0KciSdx2z45YWVa2TpW9ciXJeB+/J6oaQVGK54Zkt5g/TEZ9xxBx2/qkgAge
xBnOtzIqUEc0BxP+YX5XQSf9r9Y4azigW92QS8rTHI5ag/Y2CwikYr4iL/l9Gxdh
3y9Q2KDhvuVaFmj8ANNn1M8mTGUCcXZFVGL8Jj/lluuLK9wBPmCOeoHHyIZr0vpJ
fchcjO01S21XE7A5w4d+5fK6YtSHXHb6KdDm6rbod/9QGwXegCCLSZyAVMeILvQv
Gc5Fmq27uSe/Sr0BDul28szQYDjIKGl//7lrAGFe2Vw6LUofbUKXMpW7pNQgvrYS
qOXbq3ib6loXgBJKpZUmQT1ABwa9jwIqrM3qNILz7Kq0dBcMv3rpsH0m9y3MAZqv
9CRzS9rUkvehAGxldfOCg2mnXLUrX4cf8zibJHut2EoJZVLzXDeFB0jXHEPbRJQL
yTOMyaG1ROeMFDmvUXLs32ASiWMpLgNidor3z0I2rYfYxQX55kKeXvAApm+aSj21
Dx1yvn5CYQmLmtt/BfB6hffVM+ofzS4hXb6wBQonGJC7yD439lDG76QqKzGHSZ37
bV6V0GNz7WcNSQHETpTYzlS2F7Im1AiOpLKtW1UCAPeJE2zWufye2RS7HSlQIxG9
8MAp9VSyxY3fh4jkSsXien5Yobt02bzDV80N2+72nUMVvRZWNHNDJp9RT5sb1LGA
excF9SXlRvnFQchiH+IPhmTfbfwIbYBoXiueI2H2d1V+AMMLgR0U0BojlbvoYiOp
ZFVp20fgCgji1EZWz7Qo5pl/qeVS6ZGfOZqberPW+GOXdgvyU/S0YBAitQbrcVyV
rHw7kOXtdhuriSOqHTi67pkY+BeD3tBHNKD0BfPYWmpHnbkuZvXbi6zSxYx/7g6O
qnoF8h/WPwQ+ITrntsc7Ps7RCkoSWU+0JkkddHxr235YEctXrm7CU+70JgQsPQf5
ie3O6wuVIbOTNIW7M84gGWFm8gmHUxbiR7ONCn0zmb61/A0Gq9Dn5j7AqYS0/Pl7
A7XfRPSmbrXZe/n/ym0jvoIrJTHWrK/sgxEiHJYiNOi7ldylqGuYJPpfqSQGQbtr
TyHqot+m5V5xmMCAq3H8Ohl/5uooHwNz9XjZpy8SUPmOGGu4NPIvZ+v0o3oFZilM
oZ20tlJsq8fe5FlOtE25nvlPyqCW8RppLnuOwxq4mZCB6o2iZxzUmjdGB6Lzzu6o
2PcT9j7EQghyp+S8IStM0m58s7Lhg9F6F2frqdqLhmov7CnKMhmG4CWIrGoVHEWQ
C8MEXZlSubXZUtUhhJwGXiObAqcBMLdYwrl4/pKmKr0FuYTMIPlGSQk3gva6nL2x
o4HQNf4jznCnQFz+r2giPKDBCayCW9Q9+oXpWzlgWDAnOYQW5QXtdpzD0yx3uq3/
UYizzFR4TdG6X7/HlKzl2k3g/xpBsCmtIDd1wNO6BtOKgvfnlOjVi6+s897wSySm
LRUHG40tVlDZltYgSRicJMdaRk5GpwKOC6YXgE5B3jHBBb8FvYuxH3il/wIFPeo4
rfvfZagZJfG/y9KQeT8EVdlNIhI2GwIOsjFzBXjU1f8RNKUM+vgrB/TujYt4lD0N
voLZa+0eFqyVqIFuR3JGwoaQuleiVWfFWwuIazYAEB56O/nF9cenGFqGdL8y9/ui
1UpFyYyGRYvf9TC/jwVsIAA2xD2RpUvPQ60KONjxxIyZyCd4qVEZIGk+zy8fmHq+
/sUkcrH+Pj2bnrLpvKyNO2YvwTQu2W25t1wY1SVc8cUNrT8k+LvsS9L9U6J9YGGN
CzBkByW9QEb0PgMyxs25LqR5gwLlol2TtdFSAeGQfOpB7bK1ppMzoWeVuPfyEVx/
wyFByKa7VWPIVQZh8exrI11wxrkZeZSse531oI9ZVCgkEEUZn55rdD0Kros2BTCR
0NCtxY9Ft17UvP4AI8K6KNbKvdlwNm6ba9+fSTZY0XFHD6VxdNoPo+a7BN97QlYR
z2eXEMjDhDeELC/WqV+RGojRgyyK5i6OHR0Dkt7pyv4jb2UHiK+O2yUt9dVu/MnD
ITRjK4907IitUcq0HRfvt8v3hsmfkf6OjRai8G6mib9ukTQs/cgZV5Bu9h+9g+Ma
OJByxBmu3eQUqTUtdjsFUY3eOOML/Z8IscD/zoEBX5ikZ3uLPiCqK3upawS08nJq
pfhWQqrT6WAyfYIB101rZRRgd9/GFr+FsKkXbXi1St8QUgU39aElrQ9z53eJ+Id3
Sl38tq2eaxuaBl90H2Y3mbBcVBtcOjR0nmeKDQZIxvDJLxvY7V8bMBk170rcWRS/
b/huH7UScKt+IcLVwQNPs4/XNx29+gS2+K+YibWJBmfWn3zDcv384bDM2UGFS0Qi
vHosEJI3PCanrib8o9OevLDOFb0edy92J3c0xu6Smj93H1Pigi73n4cJbGNiyTFS
nZc6bKueHC04KmnHJiVlQv8GoC8WnJcHz2A+1o4qSO2+x1AtJ5g6b3xRzMtnmB8F
P8LfOc2B5Pn9n3Up+IcUqyIt0SezULYWI6RY15g4jcdsBQbNjprkvl/CtkhYynJl
bqC9MEO8sDuyfWd2JtQYR6Xke9+5kIb9mfodXpWMOpSRWfQa9NtEypAXh7a7aecF
GTJK2XI/3+aqMBpKx1GLKy8OMV5E611Z470q4caoIkhGZAr2vVyFOJcFwp0Y6FFP
ZXdxxkzZ3rSELg+BOQ0NnJDgE1PuZFmjnmgj7g95KaWs8vmVlcoOXRfrYfi0t6oK
fo6+5zYfKxyvuFnWzQg2aJTD0m5oct7ek3EiBtgakhErAl8LIRTI87pOYDj+qXwV
ELfLdjDH3hCgXZa6xFUO3UTxWMbVq+2c4EJ5cL6DO9Ag3tef9gu4RuGQStOhNwqW
59jgLtaUl2ormsKKw0toz+lebpUNkN46KKaQuiNxYSz5RKwXy+onI0p3+2RhQvMw
evjVtBUv1eQfR/NLYFqLI7N69g9czgH5dvghPs6RSzLWDbCnOAJ+Tjg7zB2ihpZf
xfqpQe/5mqZknBvHm8dnrrCD89KADWVXdEmnee1pmP+/IR1x0hQ/b2wfnlgDbD6g
Q3okU2l1uLuL3npE+y04ZloVlwQxu/6VL5nIaHioyem0O3GK03POkZPk5wMp2jpM
hUrhkq4/pf/4iwjl2TnJjhJGBrv8erX+69CQaNlzxexnvDXm3DSEy/6zdLSL6yIe
4APPCDZlJHQPH3Mg/tblBpBBznsd6DIyi5Qs4t+Px/0qJ2wUpJDwYFOInwW8NET6
g1ayj6VBvJYtgp3jn4NU0uj7lIH5qsGzP0EbKny9iOplMKsXrEVf4q4awv9BRr++
T4wvdPGiaJssZKQeR0dIvy92i2k/nQhBTQXgxyigpisCtd15gBnlJL4zaEC7OLAN
Hyn0VGq+ZJzSuFE0mHmHXhYRxErDhBJUlgwf8LmfRyw6+A6hJxN6j/P1vUTsc3kD
Dmn8HKJZeQcOuXdm+mOF4IgKhxQSUlibtQuy55v0snfG6hIzqg3y5i3lzJARXAL+
b+BPQsTX4ha5NKvKkq+TDinF4wQTJtzYAwMILIBgGzQOYU/FaiJWYkc4fSOq2+eS
8KSCopkBiYnb5oMCVHh8muT/A4iIpHSHRPjqj00miJB3rCEyhL5JCxOnsKHLnvPw
ivwAvMl3lKwjwLaN9QF1TySSUmhlFet6iTg7cWncc9VHsTopikER+4apmZRpMLlm
ko/Bu2YxP4fYUJkpj6ZphEjrgHjOkS4kRsduZqE1RRefz4vW/of30c99yJzRGxSY
b7U2r26EYcVaHLhoX8JOdBWrNpSeApRQ9StlR8yFbG3AkmoX735VxAmso14yBUWE
Q+tgeSjIEAQAclu3Gta7wm9PgpbGMUGl1XH8njxcH/660DVzn5kLqU1SwgPbhNki
J8zsqCNRC3d0buPX5YLZL4QpZOMR7BAie5yR3rZ/ZUh3x37D2DluxAiGiUMU8VgX
liOmbolDuvX2bpxec4vQX92n2txVn9QlAcQxVw1tL6qaGAdKXdNAi/mH7Tmt5QhN
VtlG5jJ57AX8LK/pFuVW3qvtvQ36z1Ekrpc7iJ/iZVaqA7yYVZNfWWSQJmVrRhWp
2BNJU3LxdW5t4ZYRR7cU1MOifpAt+1lDfMeUIetOgD2Y82Hze3C4vqKkBSNWWjyG
8NGsl4YR9cRiqThGCnGWYTQWfkvEF674HCYNI+RvLggpLmrKMisGTfjEW5G7q21v
83Tbc1FOybi36NHSmHuAWcvy6hSpTRId9w1k5CQi87Swc7+7htjAxO5aE6d22V8Q
kNoTJaTGfkMBDXY3BquTFjym101mtxCvTL9nVWSIViPt6Gh1EDFBYznFyD1Gj0qu
K9cLh8co8KLD7IewOsW5S/raeir4vwOcVDauBY0DLMVCRQRTRt3YS/zRRmBAJyB8
+eHU2gvK+1D1kbFjz53IYw0nsrh5RCeKx1QT7yOXSSr4NuP1gVGPTbwKastQ710/
4F4vA0Bdb1tEnLrUW5EQ4dYs8LiG0wbMkpPjfMOaw5XjHg8ZVdGcX8YFtjQBCInC
Jgl3Z1H6lfIM7WqIhPs+SWpej9ZvszwfyMLhC2D7Y0rLqZFwXMW67+ToO3GqWZCL
kYK7Z7SLLzaeMx72iEl8dawVeLukQfy4fek5USb6bcPPXGU7MdqbJ2R7vTgsXl4E
45zh7NDOtHq/L5Ad6RxWA23L7zIfg+ILTlpV0pXw//ixanuWemzX0uC9hS40qzDf
bR8/vigvwWNZNsfSMyznAA1wpIxZp++6ZlB48c9XiY3QhMKanDtJYmzV5FF89uiU
EdbM1MVJCeWDbct4vFmTFmu3g3ng7p0XxO38ARa47Fg0yZFCvgpAbj3SadJ2aCga
VR7Ks/eF3DcFS10hIQjy6kS7EgaWgGYIefkJvwJjykJwy9AwFjkaOxLyDFVZNios
3nvXPquURsU5Xucmd9qVAfuAQSv2ZtCsdKg2omkMlqvf7OS8SzaSoq1N+3AlWeHp
MmgMCXjTe+kYDi8xwy1xH+Q+ixBp7NeSD/OFr/XJwGviZeB7p5z+0VVXRHgKwxS3
YTqYXP9rq8xNl8OVp4x+IsKS9DJys2vdhgXw8r5DLD8aU6g6Kk4atx90Mph/dZQN
dWMWW0S4QJ4WokpgE7RafoNgV8GdeHW/t1Yy6PZZNg50xo60O3Tu2Sm9UMXr6UIK
a40AY+cvWZOTnFv7VrWflrKuR6P3ai29JdTQFUObXkuvtNmiNo/40A04nijIfMJY
CIHNDITlz1704nGlf+lFw9zSc/uqb5Vu2EXrEdYzmYbG6y9LU4LUk1J54TIR2WTM
lyZ6bIVeXxoGSaWil7pbW8bKcXtCdkRGExYU1SNEkUenxPADIRE/fheMny3LiPAj
MY42TUUi0XblpI+j31AItusZSQ0UtbfzVfPUUmpsMtpsmQYOPBU6GS7o2F8xynAD
GUfnk4DFmVhyx9YNc2Y2Q0ZSIZl53rcAT+9od9D9JA/xx4nlUWMxGyc3ivGL2rqL
oskgfrAo88mxMqy/PzYi98IzIF2aD5dtnZ37yId+6HdLpQp0fWXisKR905l6Tvdu
CTLEktJWG0J7sRhqeLJx3A8X3mmtd6dPtcAoky2XFzKG/kuPc8l5UvYCeYBDm7uE
cAhUDnfY2mLDyg8jLPg4+i/PK3ZTeN3pkmn5Z6XyhZjthyXRhNejB1f+VGkhdLn3
bK6xV0WsPaXaSko6LYwBb7u0XfJyRzZKfLPliX1+qWa6PvY9dgmgO/is2rLxTntf
Jv5epjU5LfGquybLPaG45JCNyP3IonYXupVWs06Nc7F2SuZ4FdKmRt5HQdGszD1x
83wF6MdEs6CQugsAF1KjpiSEhhKOyYd+Ois3AHVYOprDyTtqRIkzcvMcjU5N9VNF
HQRgTLi6sHX15qF/SAXN0dhNw+6lbcrGLqmrPnX8TRC5vDhnQznoKB33Mg1E1Z0r
sG816osMmLH0I0Ni9fKnO3lvLVyzNt1GyV6G4sVzvmLrbS+E0o/rR3d6gVEM3RbD
D4Ud05yJHNYAXNPNEcqD3cDuSiBTujuPncOBoHnCLelYFY3T1CW+zo9GySoNGMHU
jaswjjffZfgz557i40n6CAmlCiudVvfb6DLlQycQ/P5pQ3Xr67lf/00piVZsFNGY
vdbcMp6nMB//wi5tfLC3V1u88g8GAJWBky35ZMufSRFCAsVl7BbTsnheR0KsqPMC
0TwB3xxc59m4ha6FSRCWd39PtelFBYy2XNpzYMaCHW7KHklNSe+bl0AcZE9J3Bje
ru3R434EkYNXorkD23F1O+Q98S1mKCOGEbRAAfzE8B+8NjEwChFRyiuIDDjsChYG
Kd4Iyn+03mYlnOO0JC2Pk7RfHl6R5Ij4AplmJXo3gR1+woECejPksk4IANWNrGK1
MtGy9MRi5/vkvJXaaORjV0QK8v+B0+KuqxebkQPdvwHY0mkJ9db9aqbPldlru/an
Dl4EsE0nKE6w2Hgiyb+OxdE2F9IYXCnTR7fuS+8JaczQR0JKtX6WMIr87XhcYC/i
A2Slyi23RcEVbab5laMkVdcFKch7j+BgIB+ddQdzObocjf6lNAEbT/6OcUfhJBwR
SHde81mfv7nkMcwWDFanF8bc8sTnpX5JnNiwWDDw1r80/FI+fYZ5zb12EzcT8VBF
QGfbDJFV539kz1s+xmXxH6TlMKCMXjgOvJjF03VKwL7hWd4kUYk9H5vXT9aZ8lLF
P7AEdgNt3ASJM/gUF59r9aBr6omfONGz7J9N0H8RsSl3CGGkL+KajrV+uBa/cd5o
P4VY6yI4LFP+jRkazr9MaDLxG7kk224l/7He1rJ34gTY2f3wEcKhRiHd4iHCxZ/A
W8LjAgH7U8a3f46QHTRBi4LK9v4uOlciUW6YcNrnj31wGb3BiWFtts2otvrfkWgW
RxQA72eP/4QDNbnK3NFDzhmhFmhLIBjZGFP4gfPMgTZ4uUNhE97z3ESfhJgAu27S
0s+NvGnQcONOGxdQMljuLkaUiiacySfCsS7RdjEX9q3edbzw8fAxQGyryqsAEkc6
xD4AFAwfUUhcUA4TdUMMtO7NbsGiE3uzMmHBKGlrzJequnwmTttXtRRR0LwrJIyj
H2zAr5khiLfhlX+N0+6kMmeudaa9f1+xJ/NlCAP+4sorFZmE1rG7xZ58uTbR60Ke
WPons+G7KyGUOG+67dp4kleI/LWfaPxm0mhk8GC48Cs0i5lAviv8vMZOuruZHpxt
e/YZZEpk2VgC9QOKp/w+SUA08F5rQrbz5xwoWZvmjPwCpzP/LBe4Eozs0MJNpVn/
DvjC+HGSVgVSxhqJ5yX1kmU/e2CL2360hPiQlr9UPrmlEGoxwct3yEmZG9wQwHXD
bSsejb6DzpU7cbMmEI3d2R2Z7aJ7AQpyCGYFJGOI5bg4CQ5arrXtdiijjVHPigVE
i8++Gv5VyZnu4uMgena8t5KKVHDkZyG6AtQiA1qdLVmVfSmIURRsDq/npoymuoGe
a9HSLw3E2iCgfEatbmNiPQ0/uUfyfY9qmDNaMp0WTW7XnJDkmjwxil9MtZBwi/JG
+LuXbaVoEC5nA8Je6a2+r9vxJ0XGKY8Jqjd/wTxJHplEaOF0sduNrlGaxkEYoms8
GTmE0mxmxIiTCySqlIrPCfOjwbQ02/ynVqJiDEvJb22+0V2UT5T+1iyHJO2pFEBt
RYdlKPdNvPY0Ui7bw8LGa8CW+/+i5GbeXLehLjO2TUSJHzqHGCFnMPbByvgG/hKH
WLd12XWS6QQR0CvS7sIDMd7y+ZrhvqxpxbADriIWGLP84+ujZoKLdRcwgZwxbnUZ
sO92vv4xvV++X+YeScZdL6RHTSYkHp9Mp5sSPwIDFqHbdzuUdpwAf+66wjtSszZm
N5EVZBpyQkrsQA1L8prz6WF8WiHEXzSDZQ7vrvghuOEwFy5OyVH5BFJGp7SXjJeH
A4UQO5gx5P4/KWxFLKov9+gXlfd7EMhqh/BYmcM5lwKRfTm60oLUzn6GyzkDXPIC
AqT0jOGNgVpGgApJIzRzeifXYD5m1jd+yVirgQAU298j7ipiX61uUux2ocyXWZaj
k6OztWoU4toK93RCfqPtBsYNCGHaspqug/h7oUAtkXR9A0a/5Xgh07y5pP1eCsTk
dRhLZ6RwNb38h7lj0VSZfOK9qyg3FkNPLpEbDwBFOKiy2qYhZNOHpN+FdkJDZWRr
DxfKoZaheqN99xmAThuqqx5K9ff0Qyxeri/3TMIpfbqOJ8gbDldTLyJL8YB0KTLR
5baWi605971bd2Y0V7JW0G5vjvmc9QkHWddLCg6JxYbtLdopMDd/GX1A+xbBRYTr
R87WFpNuOYEfLEt1E/HahiR8JVaVg0jtCnmSbEY/llxOJwqCBFkhV6ofzioWth2I
UrFpxtZwge4693B19XGS2MKLRgDLzK7d7nfo0ml2U1fXOVcf0owvKAmixugzIEhF
ArugQ27xjLRmCfkKuSLaGhYzXGGz+U12akCZtMgD0uZmYkHHueTC9u+AC7YKv18h
SOrGhzOMtvwgvr+9HVwFu/ZS6yOriwuZSa6YzI+tVHYTXdPdtEcziLBr1EZT1Oig
oI5NxWoccz1Wbc2/jLr97lb2JpAk11uwu8dujMVn7IESM8GRdwzrsrRm81hfHLbj
ycvryrm1C3XQFnz2XwPtZncvwtnv174KJl84k5AUSSid1GunD3e161UCpLVq4+3a
GXJRQvRbK1+PqPOqwL/CCjn9CC09R7yTBphlPiBk7stzvZUg4PcAnK1aJuMgo8sX
TXx8F8Lxjcgy/S4f1SQCdPa4hz0VpKfMRPc3Seoki0d4hX3d+V1HI+Eoi03ARAtf
WQ7IDuUkOCMq+fbWOZtFTE8mpGRhsRuHCVdub72qHKVuorLBwZJc6bvBOp9bi55X
yGTt5UYI2rIfNtUsTKL1gXLX6aEINIhWrhB4iucX2eil9IjSnB0Qt0pCmmLwDO1M
heyoYPYXuSVzJNgRBaxWFC0ML5zabhUhbSnjz1ZJ9HBvpgn0oZ+UgpzwvAMiUo8m
QRSx3it8vx9auRiVpcYGk7OIGyguJ3k2tUnavV5P+KPD3GQBgkKwdoWiYBGdVq5/
WUmzefq0RgFw51LYSY/nhrX8nUyuMfqK1HsWjTZg1DpadoKSeiTY2ScsA1G040XE
opCUGmq/B3Io2AWIMNoC2k0P/fOCEN59Yj5PzJoG2PqTHEhKMA+fEFyeQySQt7Nw
yWwfKlaeHlgdHQvCe6nFM4/cO8DU2Izipm6kyVK5NnJpj0hVRT9w9zV1BMWkbA6/
jeqmTDRw/og7FB6ERNNCxviam4CIQiOGRvWuaPcwJcnsTsBM03Why38eC5kj5CDh
ayUgWE9C3zvpTmSftz70HXvlLyCeLzTy7BXOLCp104sYmxkkDr62/K3g/TMA24oY
xCb9vUILrp5xk4Avt2FpNKf+7S6LGT9Jh57vTZzatwI=
`protect end_protected