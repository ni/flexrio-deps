`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 13312 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
1z1b9VGiiW9Gp7THxpOgESt3+6sSIOLxsB+k7uXOpjZGLi6UvgQ+eWKGXdM0eoNV
TZYXrfHMjoX8bFluL1/55z1L0+6vAAJB9BwFavfo+4HLS2Sp99QupX12epbaHCBm
Jz99vTQA34xo3vm9PtSfHiINCrNhdbKCKFtYNGC6q/x0UTbua2hehrXO/IzY6fHK
YUnPWbXIrVJzp2NJFn/uGwHzLwAyHhj6eAj6WtBhkC27QVmcg37faSj4CvweQgCy
kloYnVDPlYfiSEg6wwG4rV/25awuyYnJjLiXLOOJRbhNdY+NmoCKJ8SgLj4I6Kvz
3NJzK6Ak21sbGh8s1XawHriDgSsJ0DGawSkvS/jvLJdFLBzlTeqM47Ktrh41rzHz
+QRRXWYyCP+Bwqg5JPtbZxDKhsHXNrEoDun29x1alAQoUKSwYirZ5QalUPE67Bje
/F1J3gkv1uO5916UXTWYYAL3s+cwWOsCpmni74kG6liaIgfDyXjFrImzwY27b5LH
Ya+Wl0aJHpm1BeSCpVYgJp7wvvDTc0QFCLNba/zJ+U3SfZbVhAWzxpZ67t7a8xHy
NPPdl0Y4uDAfmfENeIHBDObC6ii/1YCWP3rR5oaaBUHN35lkXaCkqo9bSYHmg1L8
iFI3O9xbXOQGqQWmjQ5Y563Uvx/nci1l/H6vxMHKGm9ayH8AEwQYUlTJmO0ZDEow
lcq+tj4ny/lfooyj+50xgHIxxxyMuZ0spv5QHyjXbHxp+0rvmnUs1j5ibfGNyV44
N1360BDMxplDX88h0jS6HNf6NhDeViGgKI66tEaxi1UpLnUE55A0yLp+Ta8CUKXb
dzV3zXvGEf4tM1kOf42xXTHHVqZekdOpGwyj0A6rYKOXlPOdpL8LBD7OImbNVyK4
K0p3Vgdpr0ArK/f3jo1suBa9g4aft8gT9IliZyPIpGIqrxZ5zoV5kSd0vyj6Hu/v
5fZi7mOaU1xcc07k3gXVEirzX2JeoFHRC4Oms2FD9mXLQrqZuexYjm88ooSjs8+d
9K7d/QUf2N8xLdIngoUy/JtzGIIgYM7s8u77sq5yQozqCXTze0x3FJ3fuBwMIjdY
vS2DjxT6TXllwuFHvWywktnOIpRHLVBPepwNXdNlkS5ni4AQF/EqCQ6BJGRVH9ow
LxqsEzZ36fUW4uzmhHCuH3Pr7UK3c49peOC1xBQMJKV/4siCJCa/qO841KdC2RPo
NLtOM8M0OMNvPFnwX1Czsh6tZRg4TRf/Tvwq6RB/pahK+qKAZyvoUUXZ/+uRzlys
GnnNucs8ewVkWpLmEwLvOG8ZX+cOfUxjL1kmTQqobDO+XbJ3aevRhC4g+0vRnGaE
aerurhXPJzTEk2QHDSjVhICorvK/1mpCQ1/iCvepgo1oGR1DU6oQdSdwXLNzlLxR
IAstqb6E5RSkUooyRvKcbjwDDOQgtBRR9JLEbWf0lZdwhiE6fq1LMjQFJ+roJj9R
E84D/GcrcYkuwbWkGRQ6UQQ/MHY9/IDFM3Zzi4AU6RZdHl9UwSBiVK1Ai8AX5ASz
oArFiratrEHxPxzhO5JwqH0yuVMv3NwmxqTO3EwxX3F4+0WKvQmmLtiv4gTiwZ12
EvcqRlm3/+oLslZo0O525E1oTMKZNzQWBmjlReOhUN8YtRz30TDa/fN2m5hZNcub
fivik2aPAz/8yHpLyLP8mFsVTGq7WLC4WH1wbQrhhoFFa0iU5zaMPCw9G6/ZzAVc
ckBbL++zCzDD1nFtHrVeq1kZ74HbaSE0JacVp/y1NvLYa6nkJRqCJRg2fA/EVZGW
IaEKPu/XCq7HQ5opBC2mnJjNczkNTuEDUW7tlsddJjpDmN4/Ib5IRUMe/0Is1oUU
6BPBQF8GgeKtZ3NLm+WIFpm+c+KU2ue0UIuHxkHMTC1rUWo+ozEvMcpfbQ9Nudot
Fr+BwOz/BoGfVo1lkJE4eY6aendKD75w+8AqwPQ04fkO9/h9kQmbihesJpHZYhje
J6zfgh/E7wBjCo0sUB/EsjypBVC6PTUqCIdughgy2NOItvjCa9e95R4m7Gxp/7T2
7fpwk71+tBaOhU8FlPeh5/ro62eXGajO1WECeos77hax7mWVOHnbF2TI+ji+ftwt
PXi4epJStN/kFCFwFbl2v9o7vqMD3lTNPNMpr5np3mlHpebCRJhpUU2DYcx1SJ9R
XFYfXJJKV9YdqpxTFWAauSF/fkS34xa6ASSgzkViV3pVQx4qv7HvZ55slO/zLz4X
12TpK0Wx7u7YCKRVqXe5ZXSC1LKqRX/yd/O8DhR/Re+3aKs2enIeeJPMoamrE/db
12z+Ss5zf23NjpA8o6a632o5CgeGetb59xAq0i86tmiY7MThSFHE41dqg7iEHl8o
+nt06e3izaMozxNwlo3/BgGiRSmfj0QMcObyv5jk3Aic/opRzLB3vjxP2h1Q0rlF
D//PYDDzlx38TPEFDskD1hYEK1TUjFiOCUDVaxFZJSCnaH7d5hvONh50xm3BdzkH
2k5tzuZs91JfZWYFeoVqPfEHe5xQKYwB2z2Lw49mus/ngewn/lGkRwdqYEwweUMH
5lkUg/vyvx995bALOgVILCPpBJ5qnN63wE7dHO85Lh7TIfAROZrBtFiwJPSOShRZ
qfOWiDBUkUrltkcQV17fPVIwh8nic7bzSZSv+1dvuEK9NZga9yeVcl5GWPlZTAHH
c1NZ/33EnhMMGHFoWsV7BZq/r7pyJAizGnIkkXmQLbKr3dsqFurbfOLVTADRoXDI
pfKG3OUIvXc47Uy8gnHPaQHUxCd+N7AneJ25FXuUQ+mMYcMVFRE7s4fLfwrh67UL
uLhK5VeROp7Ip9SWmcLJAQw/r0NMMDnV75UfcXxMDf/CsqjtxK3lU7S74DAEb6hc
fgQeudfvi3HF2X8u3/enJkYqTy7vWtU5Z9v/R5ODgY/zH0oYAcxRr1uKquOjgesX
ttI9M9WYEXGMwQxIJvf+QyGmg+/IcCAuuCYSGMYigXJM7svFmy3j1UXfrPXpwrnm
A6CPquQjNV6z7jhlEsS/e95EHjW0GAvihe4pFm4Gx6uu8//P7iGs/rhCA8OrU7av
lRSz94LbNeVYZw4CDfZMgmoSVyMycMFfaCcGRRuSms/umJXRGgbRA82XiceNwRa4
bhIr1Qs4aGy5c6ZhYd7km9vQu0K8Nik9JDjltAH5jpgHfuuGLIOX3pJJCyicG4vQ
bFx+ZGA+UCr0f1lrme3OddO/UWOMqTFB8dcuqG9e0NmJBYroT0oui4JTPjgvazq3
57yDZSYTfPpYbPwjxEQIIB18UNZVoBXgRPCK0F9mbjvtjcK31Xm/iDo2+gy18ktu
daXaaSkMB8ltlmOjh4bT7ES7xVHWNBm5TLOPMClN/i5dEUJf2H/VGSBbvnkTDYXM
zfOH3WvnGWhfyH70NJ8kpSqYhdcJyCRPndtCNkevRTqe+5t13t259mNaouQW5FET
ek80dsRS83QjPkCHl67GTehYlrz4fR3hIKVpL7Vgr1QN/mgGyubk8DJPRgoBb/L0
+51DEBJ2VJFTUmKT5dnrs6KZ6CTXgaz7b22A3UI3cjeAn3MZ9z+j/rkHwKWVX03K
qnsczaiLGX7bBwuXTvtbFcAWQEdUNQLKXcK/WpfTUwsWoODl9w70jpKwmjyIH5qH
QjSkDyrMYqL+GVhsWIUqLRcAZ0HI8Q5fPs7Ph3GBqK3Fn2UZMCIn6pAuIvPbOf/Z
90aioauGyynKUgyzn1rIP+BCxHGiIq1hH6Q0hv+/y8jWhWTaKbgZpgVM72PZku7M
W/jgez/bwSMd/Y9uQ1bNbXa0rGsEjumqNiLmK5sj1c6FGQdmyZ+vfGfPPSQ9mvhD
vm64qk4u8Ak6VoSQ57jIKFe7aqw/8jvtkxJxl9cozdwrb3dZEn/1d/sh619t+Iif
v8iiJPEQRTer4ZJBXqCE6Uq9gs9jPoxXe7/1FSmdWnHUQrOubI39HbthnJB+aVYO
bNCHJT+ENP4CyESzxpVsoDH9RiPpEHoaoqK4gbCHxDkfYvc+WM8oJQOYjpyco5oS
Nl6NFSI6dnjOSnFxFryD4RlEcAAGsljrEQ5AM7WxgB46stoj6E0Bje+HGRVLzrCu
cYv4VQa7R28Y/H1522WXCJvmBOqOVsfly9WuhSOBPP7eqYyG14zY8QlUgjyh3CJX
xd1y6NQCd+sSVgDTEGH4UiuNW82KhaSp2FJQqzDbCD6NTWq0vPUXmE4hyloBQlTm
qhlY3bXMb/blAE5+LaHtrBK634F3npiTyv5UfCQvaQgRBNNvvp1lxWf5YJRISQm/
fumwKNFRQqijBFQTbCExnA9tyR5BQN/wLnS7aTBl4J7RAx5d7T/eT/TPeaTGxzc5
v3iaKtxMjbp1QGUCCwhUvIdnWnPEAses6/yf+RPdJJcyR6ulfjNNSHh+URdqdgha
gT//iLTVz6uERuzVCm/VAGocMukKUtgc3uACWUKbWYSKthjTOycnDMFVSl7c+zbS
o27AO8GmepcwkaPvg0AUzdF6H2+NoSayf830WsCyY0IHSw4eo095aniJ1vptOJe5
Gjh9caKlBgjVKThBk2LZKLlEmpY1zqoLETwSqN8wuQautCNTjSGeNrLNJh3+TpGT
RgqN1P1dEwvPL41B4MGjE2+8JZOcnMiQqjc8Sl1HPfAqtExw4HZCFDzZSrWo9MD2
EZpfWn9YV8OcFQgh+nqVYNmiju/dBjm86Ne5oW6cGo+CISM8a1UEJimBi9eUVWH6
wPQaeiV0B/bxdKxlGg58lz9ytjO2cgw7W1PEUDKk2qO8eQ08TTLc3+j7eS8pn8GF
COpJlP1RaHjPXKh4iFXx3zDzjJyrQEO3uNns/Tfizy+jhgmHMlj5aGFgwZpzEL2W
8bww+87XeKltczC6RBnkDTUONSM/dn3RhuFqSQVdLHW2zcTWKzd8g3FUMP4TFHIX
PmORClkR/yt0oAHStdnIoRYsUu6SAEMcfYM/WixuRzEpQzkiuMvdbe+/OO9zjbcx
CadzCnE7JL+w29i7n/J1fQ6c4x9hJJnAt5rjWv6PERTr4I45ZyzmJWIAsf76BRlK
9jBU2NcN5y4T1QHc0ASfQ1mgYJ2Z/U5AvjA4lvEgX4SJcgO3WG1h0ZxE37YQH2E4
k6E+I9iKultlI3kBptstfSS/RkczKIKXbRrFLzuRUJrAZ6IV2mxYq7EuhzG5tbFf
sjapZvGmKPIlQbFYRiOlVO5uvSe6TaISuHrJE+8uuJ25CUrZVLyCqoOQaijaIgCr
sF9Jj1DQpKbP25z7zm9skUwWZSidZzd/ztpr97L3Zo/TSGZj1FEyaLIYSpcJrWRg
hZu2rEod7rSbTb+119PfOdl0bVPSQjCa5vTY9fOSnH3NGERVgsc+lhx220TMN7zx
9A3PTdnuuM2WF0uwliAyPQv0AR1HHJ9DwHEBAPEW/vnnZvbfPhzjEOI9331OF+9y
ncZ/XXRE9tJ9dPKwjX4kMpC//zsgy00NVXMajy3kvXKE0ew3Xmj6G0Awm+PMvPGG
QE6rSmTpYdhQEvYeRQzrbowyc7wDgTo4lA4ZRBCXv8rGicLxduNHe6np76FMV3Mn
3yJMvzHU/5zqO6U27nEmKfGZGsuDy4+xk19+rY6e6iGaOwg/l0oAEqDmlhKzuAPA
sLOWU/Xw387Eh8vqYxVhLDMACqbjm7J4XKI/mn72yN4K3gk6eEfswRwk336qFV+6
tCHCWcWLQzBuuon7GYbakv6xuKbULYgs4YbCLYL1BhciOpviDmd82Oqk3LRlFBWT
fcHVyRJoumLq7bP87wwkOUkM1Hjf1Qy76RNB4WfSxTvZnvWyHfOWYcfp11uzSa81
frWm+xvKBJQjzbYc9b3alFTaeE0pvFh0NExYZ4ytzJFw5vzX5updEjXLKrU61n8D
Ua65sOK8pyCFjqSrNvKo37lo9nPVI9nat1Mh2YxWilU0y/pq9+MSrp43GaV5cIai
j4VxVwldqDLoUuXCk5FSNYxFKLc6sIoJbfavPMV/vKKdGM81JFFYEHy856/EKi3x
rZ2tKg5nbJTFyur2uAasazlq+yBT1Na7f3AXphZASZFxzSs/+v7R9PHu0IaOARzb
4X4Ic2fHKN7qvzwO0ZoL6MNsqkrfSgj+Iz1lRw6qcLk42Lh1+Qp96D9rX9PpTL7D
fih+8VWYwjrNeQokLMlF652aJR2uCQLQ3mWYg870o3oSgF9uKimJgGsJvVuuVp8Z
mkEEyRQjOqgkZpndwoze798O9G+SoooKSQ9Or6BoU5DZZVJMwNHmxEjYdEsTBMtR
pyIxa7cuupQP1O15CM/NGmH2Q6BjZNVkBfoCa40HJjMhi2Mz3QtY+i5bP+zjOI2u
zEsVO+wCGLdvP89FusfOgxzO37tZGvfErC8zXApscWAIOFVR6MOoViEG8D25tKbC
bwKN/LO1RVwqKH7WR6CEmI/gUHnnwFuYR91e4WZqSHDun9LWCgQNv96SVP7g6oPV
8m9HdkBiTSZ0ahF9IC/dsVOa7/l63g8Tgno8qrvAt1xGGtkeOTSoKOaZ6mdo96ZB
j1x5kR5E42CzS+v0UwBUh7xcvQvzxofn3zAhJQ/Dp7e8b0EhdqL7llsWLOUMT3Fo
x/XGUm0YkpjvQveGBqNRTpVX2SPy8wQPqvXW7IgIghTtBBya4O4zas37ge+yklmH
da53619bjWyD/fzqEKnh2VX1Mw64QRjWK0pgkQjcRB1JnwlAj4cBaukNc0ul+YH6
5C+5cS7a8dSTG4cUUtcOkKcF15aosnmo0Phe6sLR4R3LsbcBDuw7ZJQL+ThKMHj9
6grc97K7z++vce3mjGhzzNx3Z/cfYd5XitaUlnzzfJVbvrRXYJGBlFXGJF9yCplN
ivkY+lqToyEz+RJXrJ5l45yaI59ExvGfPWTV8yeqi9RU3vjm8CSRk55SUKfPV1rO
0UDUFhcJZE2mEPsvREPa8E2rsa07MHfapTFgR69QNJtOBPcW62TrrZC6M9fDG/6j
2o4revgy52fEYLkz03rM5EA5sD/B4PzKLZyXKdyU4T2qenglzPZQmLI4OI694+ea
hbSobDwaOitRTRU9mvDzQoMPD9Ao0d9/TKaVQ12d52vmOHrdHjHUgJbUjqtOGXaC
AcSNuzqYq9pdykoIvKXQQshBfXVo+W6OSSq6IyOpZ4JuEosscNfLa567xPz5UyPM
RfeCRT0p7MGdQj8bSFuaCHiqEnjEU5BVWXiQPYjp90UTqgpQZg84McAQDa//WoWP
gUSxd43+tGbwU7rc17HCt9iwT+5Ypez3mCv4TS+vvOhm8AeuI9PBXSzjhdU894Z4
eyR+jbZMDXUgtskIW6leBJ6lWaDNVtQWY9Vu9kXcD6kQdO9pm8RB+mtBFfDCgFQ0
rVtRtfNf+wlPaMYTv9+v8jeyJKpVMjikex8nhGNhF66Ni7UM4p3CDYM7ftHB9JTx
gLiwQLyzJQ2dtf3DiHtWGuV3EoEj6AqZop39S8XA7T/kb03kW67iM2M6qAqo40b2
oHEkkkSWMOa3AUAmiPYB4nIVKvf5r6hlOoelYhp1UwtDSoIT3HT0A14j/2B7MQ0X
pyGJH5RXrKknWVYg3WzReocfwaK+qAGub8iEjIlmibMKO5Dn7DaHZsd0IerOuvLj
3geFZLdLrhdESsKGbCY8lMQLSwjzSw5xbL7ThD9CiXI2In0/3eE4wJXjISzsFvnb
VyJvv8Ndx9fgtTKXGlrMa/yqdn/yDp+fafKPUP9hjZzqKEHCEAdJaCslQrj2+AOf
4FLavF434Oi0yLldXURiqS1cDOYUmTq/sRGk8djMcxhr0jC8Ygc3xNuEfn08oj1D
oIne36sDS4+ENygc/bjoAQIP97yWPdmG1+CD8VyZUGX48YRuqbtbMK2kGDOgz8Ft
CDEVuxYdhT5amIYrpL+/SfI0O2t7GgRLPkir5mvLkRNyKKFeJ2pYy9NDaGcc9Lg3
JgyP0lLu0Dcigjo3f6DzGZu9xpMkr8rPmhrF7davVDT94pIU2CrCNKa4XZKJR/3I
oAJ6/LorwH0qzQ6QGpM8E1H/TjXXo0RJzeLwi0itrZux3Yl3tHE5oiVnpeJ9ygiI
nisziCDheV32ApCUrWYwAGzFTaSsManpSwdBKLsYUUvamey6Yx8XDd8cplSjIXnb
q5YLumj5rBRB1tQDcy7dtVajhUvj9CZ7AE0B4NULNR2OXg1vq7BSscY+dYhjMEWr
HcI82PRQ57o34XxHKDnYOgwx9gR0nLgNz0xZPOIyi/ywjTuvzZYRe0iI8Ad6IEdx
WR4/5Yp0SUfCe8J4z0Y6YalnsW43QojYal+odSAnflChGt+6rkhn3Lvnp7QKdVff
sEmMO1BMksJfYPxZn9yvwLWrLDRENYAsApMnb7YL3Ef9hfXZ+UyR1riXhn83MjIj
m/qjJw6G3ZumMx0dXyjm/7Zi+KD0F8sFvmXLItoaxOrawsxYY+Qm4WeZgMQa4HFh
RudbIhJhYhzBEp9c/4b7L/pzdcBVb2WUk67WSpSINhn1IGlQBji9cWFfG3pICJa4
onq1/b9kXScuvaLrMi3FKjhxQh6UWQH+VMF9KgUvk2meWeh8M4D5FpuOwKbAdPYY
0gFDoQzFm5F8sOhZQwtPuVynxDvm0UNYVR0YG3rwMatfkfYqmMKmRqDkNrEjcCvv
KYkOqpakpWXq4EfMGGHf7lqvHatljz1I9QLRiBzomtsfFkX+bqvQ9wo2twpQX/4w
1Ugytx1TgcUn0KPgLA55ZVl/1WjBqmMawy3s7sAIH8/orSiXhSq0v3b6YCrEF0Ph
7gD2yKs4mvTJrgCh6Z88i5LFsfOrumb0Uf2Nia0r7hGeyKJhHh8AdjkfAOrbpaIm
hHTNKsPoBDHKEHc+fTyxLdc7dGM5MkunhSjMYvr9wkPy819cht8QVE3BAi+ZKPoX
vRAASJbcX9x1EJ/wj+MRA84kS7I0nd8SjQyb274tZwsVSKlbDb3ucyWXGhF6Kjfp
nQcoYmzrsLPASlA6cvl1tXXU7S1eO+WTW+WacAiBPQGAcAZ1Srgm5cYNd3iXqMAS
+x6f83SZOxNh7OZCFd97kU4SWFx6KvQ7mDmYAT+BodMbQOYXK4wHp9fOlEVm3zf8
tAotZzBmJpm9tWu4+Uy27TKgknauYQNSIxjq3Jy69wkuziYhxCPhRrre0pZxHCFf
JrFcGdKq7XfowYNnIQrI6MmoTMdxFhC93QjPLII96yOmQswJnYWVmmpIM4i5Wqzi
eBxBWGm/avwc+f5Ah6KdHiuDGWhaaKcN3LqsxT3L0BRkB0aUo6q2B3WlsjLP56wz
bFG3mpFt4T1O4czv/7j6nCuNoEhLVVSkTtAZfOBy3z6Mc+eZKzgQSLudYTrMtHMx
U8cmOL9UgiqpLNxY1RVXeHkV65vQtvfSbCtZarDraS2CN1Zzz14uDeHvdK3vfAnK
n+6uMwhQVaAgdJcpCt9w6TRU0R15/NQCL5zwGeXx8tikerybLAG9UA0+CLSM3N11
+REEcC7gZeSAHRRfYyUkwDoZ5oVw7jTNBwi+vMbschtzskdKoQkHMZetF0WM52SL
pUiy3ZdQkQvFM6mKoNmdzZ5zzwLEGigQx+I2fdOceCj6I1g1FclS92/6HUyeVlfT
JTX/peSeaOcma1HGppU559FSiJCyWzvE7o4+79dIWmw5BltyOGQ/Go0A0pt3xDBN
wHBPZp4dSnjUWdo+tMTlhAH/WgYAEiVUI+gX5NFFhjO1Ee9k58X/hY4gfhj+ILjQ
3KZFtU6JE+VhHJSMD0nGe9byaX+xECHltY01fMYWArjG0z3tNMdu7p1z7VFJ87Wa
5/yx37U/hhxRbq/2GYOG4GkGmHsmB0O506ATHeNy8Sxm8RwzEbqIsn7W9tDF7Ah3
T0AziaE11ARAcPP1FqTJvMYfjl0Njwww3GVEPoyQuGxthGw4iucVF9H3fP1M9fMz
DeQgeUWkWOJ02lOuonAp2WNERr2HvLtFoPRB+m5DBiagUI5CWLITBksTi6hmsZmt
IWeVDWzCRpOzxglHk7NHVdRtEHS50Wx3fhIOhbtFDnltL9zOfIhHqF0RgmaRLmfz
nLMa+Ea8n3b1qb6EmKKTAwZ5o94sst4h2Wm3oVc/FaHgoAbFh0p7fcOlcJZkxYy8
9AnN/msPq2jAla2TgWA5c44wgU6Yo6oSSxQps6jifN4O+pUYZU4649Fp0NyCrzXe
cSEYPZHalreCqfnqiEA1sMzksqUJTLkNnEftq6wKMDkU6p1oeuQr58mk50npBc7E
WHDvvFIfEeTYfPGE6Fli634TMG1eIMk0WJeSkNKWumJTZtuvf0qAgFek9JnuuhUz
CkT7KN2d5sdvmkBHiKibxZLwh2gKLfpqzjG0yEWYL435R2HKQY7TmifpPCEbfftG
NIq972mFI+nmPAUbqMN2PlKYXJELKZMUrTwr+5TstX7hH0zUDXgT6pnE7uzWkUhu
mFNNOkZ/FQSCTvTgSt1Eu5wTA2XLQCxFduDg30T4S/z4vp2QeXbClLf1KGRaQox/
c7Ok/LSulaywQB21sEiYtOuuBBBbt0l7EZZCBE52xxEfU2q8gvfYdoD72rK1c9I1
lRlcKcUZTLmpDsMj4r0tklbNuMIkPLJ3VxWdiET0qTTdR7r3CKGvPD4qA9PBFk1p
lsWW34qJykcYhE6nFUapzjgK9QnWbh5hfPJMfUIjW/IfoEhlEBN7mpmalxsDe5+Q
EKRbNq8/ez9XA9A6H2H92RlyBBD/35ZxcH6fmS51zHjKQ1QjQBuUW2pB+yZWiDlk
mR2ko4sjzSZhrFlmOuFD/V85pVoCwTSP6CtxrzBmieFb+a5YTDaP5f4PURPV/QDA
KqkMaJ8Z6gbJPm6ZpPg0Bpfy1CpE08qhiP5rwxlznc1KWx5rOMmg/b8Qgo4bZaWn
0Cw03sRLtJDlK2/ZA0yvmXln8IqLF5i22bt7pmUwRWBhnm4OYmBVkz4yDft17Yae
5K3htqB9ENmNRyjUqW/6/qyfx4wLtOtkip+vmchXK6YapdlSce7574QGZ98IeDiT
+ZDeiU9B1YUBPBXIKz9RMWICAxYNcY3QVVBmQEwH2iFOugB4uyI8OUF3AzkiwvNs
pvwNBRfDExvoueZi9tnfnvQV173fBOOlcYJ6gJue265RNFZSeGaQnHoxYhhj3WDc
vibhggN7XDWvWm/95iZq7w+kA+0W685YwKWYFN1kz4obB3ngQVt8DPZa80lSjwCx
HzPQzHbCsTpGKjNiQg6Kgoh7wd7CojmxsFXzq91RPA8sqR7n5FodFdjBOVf59rs/
Ry+2+jLnNvb1/tkG7wBf+Iv1lPc6uLE04VPtF32wLUuhlNgnhsxV0yc2cuOo2/3P
j2p4omd2Vajb/pOMikjiAb3blRDpsh6FqNc6ggKnJvEzeI8zFyoxQX65umbP9Npc
rleAPrkuU97gMxq1Ws6XQ3G6OBfV9ouSC4YkIgd6CwCuoDl53Sfyn3x6V33rvGu9
VK+1fJBxdRAoSaz7rP7drz/j1zP2PjaTYUHkC9ycuQcfd/KVX8243YYdm9xwYWeK
ZYVxHXPI1W/1KHmhzRg9WgtT4XjFiO2We1cuSCJz6bAo+AE/HXqLP96c7Js610HK
zVn1BifPvZ3wF59B3TxVM4cNV46wK+2E0ljY1VjavSSUFf40DiCY8HlGouGUTtn8
3q2PddLIoTRPJochdDYqc3qW2sLpwAP3AzTNtC0eF9/HLMmlTNtXiNMjGMdhN9fW
1vHdhvOV63lHMB5tZAe+OY4Xp7Kwv8tJuV2hpTaJ0HyJyFCTXkbKVFfAeKq3cE+F
4rI41JgVPXi+27vcpGwoPE8gIdSXq0cCgdnhHw6d4J2rA2c79RabJlDXxgO1oZQw
TBSQ6wLokR8g4l6qScexS6C+rjyd7oL1I9YYko4uRuPURrqgrYumLRqQcwpjMHJg
zl46bB4DGXMOHAVnmjSlxWBwd5LTXEehSPcVxgjPSK1VUbgqWEa2AbbpYKLjqB+0
DhxIr0oKGte7bV5939m/mtYN5u7gAMDzhWvG28zXAFgcU1Ly/evftid3gvFVxWj4
ja1c0wrtbe2ULjcwcimq5Op3Bw9it3Y6MrQShPDy0X/DVIsyNBeHv0Vu7MZylwR/
yY4sVVqNbRCldpzgQZMZaqQ6Kv2gdprXnqdf9ekrLHw0B+W2ACpzW6bxyRBgh2uX
pCS8VEOLUxgx0EYatjDuTNJU+QCwQHyF01KKNMJCyEKt19twh5DQOcn/Qu1ohdnC
TAmOp3EoJEnS3hH0l97ey9AVDbTqX2SZKmSdAtJkeKTPdz2fHzKm0ST6RNbDxFYj
N5XZ//DJQDfEF9Lf8HBGN9pAxs7buuOaWVPxFZ0YIvfvGeouiXZsURKpg3h14Hvn
ER0vW1v8oU1gERn3JsxzfRcKlBTeRuWCoJjGWyWaOIuG4xVhct5vWUbuEtwjetIS
Uo5VfKmiO1x6i1OxTnz6faDRtZ2P0PzZSD08+nh5wRO8T7Gn/7VYO2zp/yGj4pwI
FZGpOS0+/XN2zgYr3oe0UHm5lUy4eTnOzJzxcdXKw9BxOm8SRccMUhcASn2NgFuP
Wz4F5gnbx0suYLMJe1ci1ZhKqaIAeM9aKYkPFipI8kcOL10BuXJXT1kwe9294TQX
QLiabaeAJZwj1p1RO6H1dCoCv/cqzu9UIB7y04m7uvGUVZF9V+3x2TzOIKcMT/bK
R8yJkSVu5Co7+lYICukm7hn2m1FCRNb3K/w37aoI6CVu1u/iHRkhP/yITgk/CoIV
GHpzG5Kv46786H8koyoULbiMPL+D31bohjZrLp8oUKlkQyWqgmc67s0V7SnRES7n
8LD3o77irkyr5pKZpGduAQHpVOOmsZC7wFkQPqyOUxSwHPE0oC9WAxzrbAOPfwy6
KTcLVkWEvRZ9mAoZfjtyQ15keVHSiBE9FplNKiJHh3HpoCg+k3eLJqK5/ZACr7wE
hlOwe2zU+LmdZt4atIlVOXSoEhXnzTrgD4DAmHc9mxHsQtoo+b4lzOSxCDVVBSPC
8sJtCNiEfkWB9POAneCJ7o1+zKctx47NL0D46VwDAhBIaltg9zYJ87l7FJCESiyZ
Hlcg+9zoh8AzpEVcsk9WtiDfhaD/0QeRYZCbRofNOAPCTwB96DgnA2cQO8LI0LH4
7qYLT5Ay7z0Df/+E8wxyQGmv/Ea/HS5Nhsdsvbkq/oDOMUfeNyOvs5f7n7TGmnWY
Ar/SCbWaxCKBV/d1ef1pfPvqrqqR781cBkO8eClFD8M3/YZSHtf605aIs9w/WUN9
sLXwfAK9kvGD3BinqJNn7xeZgmx8ujZwtBjgKyJcbhgvfci7k2SkRnv8nL8fgMo7
91opAPTZoTtoSUI6XY1JA1kK/tF+avQdfVaWJI7Na+57I2o9cx6395zZxb0Rb/L6
XnUOHYVHF67fvHKB7tKrau3D8xws9vlREnTyiKRPCvXe7Dq3wW1cb3K1lGpVRZjr
zGRxZZOyxJ5jG61wUzE/m60ut/65YkXh/PrjrLIOBbdJpUJtQQrNfIT/Nb+XXL22
GsfNqxukbisvjRHHp227ulSGbOJzJTh4VpYkXdD5SxneEpfY1msc5GRZNJW0+lrv
OePZXFMXWjVk+SmG49iQik85Ts4WA9CIE6n/U2tTgUK/jFhVL+CUzifBJX0wjtSu
q3tn2oNBTM99OZYoZWJtHJnsN6KYvuGOnK6VUvxTwYh5a82HtJcxk0Gmm/2aRYLU
bJR1hIl1NQJWLXTwysRHWkjl4kg3T3HrIoJe86rcQBmrAvYP2a0YltjwUBSpAdSx
Ne+eK89dxjG201KB7dDZezEzeQl8pUZ+Aq/2IL51Ih2uomfauCfVa1BSkb844SMs
NITaqasOB4oTBHPAU7GcDX/9u+OdaCoXDSdlzwt4q+JqupVtjWembtX/a3+rNpK1
ennoHlJBCDbzzGeA2v223PWCSAO6bEF3EMqhew104R3OZP9b25HewwdM8Wm0wDkF
F7Y0dBZsw2vu6LMR2NyIKksrVTv1aVAapenYj12CkwMOBltaZfZTd2L9BgjOQz3p
B44Ku4g7+iWdLUD4nToXCt7y/wSD5z2RzfqSxQETbWipN0C76JExMa3/cOai49yg
04FNiBZJA05JXl0yH4X7bT4OqC7RauDyXq0lIzf9MFPjchitGnQUxD0Ah5WdLOx3
obXRmR6fIchoJ8lx/7ISQTURXaqGUwVewPdqWJjyqxGArMNM/24Y85Xq3YpaSKNR
7wi8eHkOaSWdhTo9O+IkR66gcTd/dA4S9PYDqWCHd8QnQkmpSM0rJgkTqlpEQ7KA
Lk67OVRo9Q8Tr+o4/twntVx84ABveN2yDV2OamwFZnrTxBo9dMAmJQTe/8mEIvnl
zLUUEMIvrfwB93kg7oMHJ2g0JskndA5MHupyYGjpK+OM2l+R0051xXN3YDNRXIuY
l+5oxMe+dFxESwtFM9I6ulKjwHw8kACbJtumP76JNvOihXEZsqUIWWncgkfDkTmT
i/xYklmpvt1UDaIZFPnWsblJtTM+HqA0mbd/nBN5b2KWsOLWNI/AN3Umcu3HW8aO
pqnH7+PWGld1/U//ifKDjAtQOHZB4Rw1+S4vvQ803x9O2UuV0oWJvqYs59PBwlVZ
HyYRgq+g0NuiQ7BuoGWLYTG+QXjIBLxi4RlRHvZGwilJyyHrifYOuVjfQt7xMmrY
k8BrW4lVYmSU7D26Dl9TP0ow5h3A6nvOcaqFS+newjbYnWwbiXxodGMJf8vBxG2X
v1eSTs/U3wfZ6GLUVfiMAwVoXUS5VH3eKhBaW7+Njuca35/9Qsh1ZobFz2gCw0ub
VPKr1cLVLfkXcxs6JbVSSNUMcAAnQl0dwIPn1iSJYVpPtb6OLJBkSb6f1Q+/1xhS
ZY0ErbNnyOFNv4LjP2vFYPjFB8QjXKIVQaQdsiUFHpek/9K0CmCdo9QzaR1M7S/m
k1BHwK+m2Dd9GsLPrg01NQjpoDJXWfrqr+CL6t+6EEWBH87OjajfmhUMV6rymnOv
iuVOnuIjJAMCN3hPizEA4PPwYHChSsh69PoMtsL5Jeu6uIFA1+y92AXlYyJWg2La
uYBi2TVo0ML4W19e6uHSHTy34DVtz3KyZHmcFvlycGSxe47y1qo5jTQ7c2hhIE8D
61902mNrmX62/FDtx1klDzF5tc/qNBppsCX9MyyZd2OuDIPXwCoc6L28SPdeOkZM
9bLkQmHStfu5LWB1HmsUaNCFO2nohNieDqrIMy2P8KkOHps31vAoyvfa89kdSfu5
9kJFh9M9XFtMTSkSXPnKtjMtPvoTJmQLA2beDM/CXDShgbn6zst5h9kc9oXmyDFe
ElJL5jJyYvCVA3MYKuXUO40xg3hbUrnc64K7rEpm785BvjFuF+v6FOf3OWscfJxw
YXXc0lrZAQ5pqqXPD6m7Q0D2+rhmY5IQMqL0zuWT9VPG/JIVnzoc85g1DueUr6Ob
R/S01Xv7BvMmkr0bNoBWPlf2ws/4PzVlU89Hms0BXH3MV20slfOG3LOjVfG90LOa
0j37C7LQo4veWWajWqeSBfXjWvWLfz7VmEG/dWTeo7Fxojy14e7wOL9Io45Gj5LV
ooouqrRaKWgk5KUMNepE8yZRVOIk3Qwv+pVmdL78kCeDYEaeqJfwlEJu8XpQbKo3
SZq4Qj0J1j8Dy0pL0gYHYfeN1cFSr7dINFG1jSZrCUkKtkW1DnN6JW3RB4tyWwjp
tKJ/DoZySe+8bdu+DW7uAlrfJ+JP/GgNPzGoMf1VsIXwQWm+d7HPNuXTnSzm6rqS
dvVF0/II9txLDU435AbolwowIzW2rCb/Abofr6E3sQv2j66Hu6ZUddlLjEJzhyWS
xbx6V+mJYGI8KOQtrhm+xj4GSWrcP9oTCIIKgu4RjVXDjsriGNghgHp9NfkeFcjg
UxEOy1QiUJZ/RlFNbcAPvhkDLFFjpkDy7EWUSLKJZCLZPHtduMKbI71gZsotZHQ8
N8y4CUHKWuATicE/Ywc/SL23h1WU6LaP4HWOiP16A2IVusQOUu+0OlngOOzl/CYc
AkxAVaXqXdghTeqGD4eh77iBzj4rft1fHM9o/qx9bDCnlIfCn6Mg8gXSqUn08jzD
cFAIYvebSDg2vHisD4K9jkryFJVCfZtLEUCmv6YUdvPFWhd9sVVuEAvR6LPQ5pMy
uCN/iXdX2orc+I7r6UfSRhc/s7s4Cp+PTCm3pV6T7kVQSXiCsuXMbIKbgl9WdwQ+
vtb/afX9HPibp9YDJbAEPVgM3lmVQm63T87ncowptEAo2IY9odyshj8nKiopbAgj
FHdkARmsGaCiBwJlJ2V936Owkqtzd8P0/d5i1X1ZGLA35tQlMg9OS/+hOBqilUkT
j0FyDGnIMemKTNIbDsBVXGjtR4NEoAyOnfjWSlouBd6Jpl5kpGljcsY13uCOJ7xU
MptWYuOOPe0dwrsCJhD9SVuQmvcsXOzqiCAdkH2UHl2tYRd3ryRMowfBqif1KhRA
Z7q2M5GQA75hb8vgXkzketCoIjwyRBzQfFspZKNY0RzyDO9p/8ggySF30P5b7BX2
0JUMvBYlTR8JwRM/Bl8iMIQ9qjbKmW4YwwCvnQpTDSqjCF+PIWIirs5lGir0CDjI
+Cbwv47AbfzOifbNDGH+KeoiakmFWHnSQWiovQK4GWex+vYD4XWVaLRXO5l4xh24
Zvka6KWz0TFWrhnPdCnRKiQIMvg1xu7Eh4M3qglQWU3C3FCOj9wsXA9VCSXwHd8P
wugchLTlHLSUNtIf+yBQBJQcPDdoBYDA5quEmLha2J4AAxhWEi13ExSOnyblA8qZ
M9jNL2uHKOBcRtPVEjI+dfeGiCzjFuZWJWTosyKejEH/v4n8N06rCxWEiGt4U21j
6hL7vhlCDakZugTvtKtrhhENTZlFAJRjUrLi+yyMUsF+lNNSTWluggoFqoJz12UR
3tfA1UUY3SZ6uho0eQPoX4qsDZ+JjT3RsK5yVIIwoJhry/FZV2+7Y5PrW0yamHWh
z4OUr6hpgcHh3nGBxbz9LOWirIsNujDFG6pZe0xHcE5ZVnkA3pMy5kkRnOfwWA9D
+Hq66Ne02hhvrcxkbAFtFsPpbeZokcPYh34RC8JKafsxaqztkG24dCmeISu6WvnM
hgA9XMCx0uMB2TtlkgdANIlfeqzxTtEGuqXIS0jjb2jo3iWymv/tLtwHhzLKAQ+4
3P/efXjsrW4fNgSHdsf3kFSyyTQDKu78kwsGa54FmmMUitJiesIc6qfrwKsSfWnG
Fr9y4Dc+OzezL56TN3ErfxeJaZU0doG2MU3vho5GL7api9z1ZH0zhWMQIwF2v6Jh
/zTORW4qe5Bri/rqZVb8yRIZf7C6reBoG8JNwt7jhNNksU8HKch56/sokbfZ3UA7
N8rmDqkvMltkxVzjlYDb5xYZDK0MzjUaBbhjD5AOfyyQ/SwzC2hv+l8i/f9nWuUT
dssxpwioVzlHSfAJ+RqNcf2Xa5Lys/GmrLRNcIIEY6ot0jzW3nzTsXYtiuPsNQd6
+2vxDuBHkzvJFOipG80wF6qSqwcfPYb1QTOQYVEtq/UVp3yRahww2wxscNQpRe/Y
EA/j/q5jdE3nr0cTYSCwfRpVFyDmASVu1+W0TtfADM9G+jEvJON7J8B9QS+c4yCY
eW9AJFbHqHkn7h0OKnaUgQ==
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 13312 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
cjljSPzTIRTXBX/bLgom+eDt6uyGNecLxAWakXRtrG8C1K4PB702Gazgw/8AyooW
aaRJ6zM4bdQM+ThHKvuqqxmudQ71g0IufOwDyVSeV74/iD9SVraZAReb0bcelJPp
sfCMwtf53iNBMGgGabWW14nD63w64RzTokatp1zmLjZUXr89bu/wDjyAAmGmYJ0g
OeWKRI+Aq85pGsYkYQcPy5XtuPOwznSwm+8cRHRQsuEP9GNWx6SZu61meS2gF8t4
2KLG0S7ibCmW/8RqkC2aY7LQjR+W3pzA4rLYpX5XSb2S+niyCF4Gy3E5C+RygD7N
QW5Wk+8RxzrYmBUHdNtw+sQRLLr8+BFvDic/0mxO5iT5oenmBOknXSuB6qaGdysG
CWeMgJW5b9cvf0ddiyPv/43BnNcWIqO3Sv624Jue1Fe1M/WMTL1kxZcCwJjLkjrN
0W5YwD9SsaC9U9772v5MiYCOCSNxx/Oj2S7i5NWA0dDz1pTzbvzCgrSkciDG5+2T
y9m+mlUlzzA4RQVGOjJE7b9rd5ozHQi7UCLCULSmvDYAOrC9LdyKQLOdvsMJNNYO
0m3XT1tDLwtDjUachteGQaezJ3oxOE5N23y/3kZqZ+Jb3vXkxJYRMUiWabfDVLVr
D0jVV2D3t40gNkJXBwdbu46Dg1ppigRfLk35V/AK0HGyJC6plBWP0BJDHkiOiGno
/8DTq4x99bq1Hanc38XQCxiR7gfgHrOpahSMVYs7fJuhbA/esYz2J/KfYeHHShLt
hQPkUZkpbZOo9jqM3o7pEw1a4wWRXdUm7VQ62dFeLrWYa3XEWzb1I5JETJk/9Dfq
GGz+l2rZnNYTNtvbsop6UkhP9Ju9EdgF4XuuFE2lKGLJ+bX6wC77YTIVOFLH0Ev2
1y0Sa/+9xYFeBQOxKURfvGmSXgBQhoIvy2x5ge5tThS+dZKqAuGHKKYMN6tagDz7
p4TdoKUWTcF5wREXZ/Z4Hd8c9J+iU9rQYbObW248KIIVi0fVwaCfeWwynu/J3Kr0
Pv2+ujuABZLzTk9utl5WaN7cBg7phZlwWWSYmbPzSCs5AYug5AU/8EluYUskVxo8
fQ98dyCqFS75lllcxAdrnx8w1Fb7N5zm4EC/ykE+rWkZLkgowtadzl/3J/a5z5rT
wE1LKsaJiAx6KwZwvcwQt5YW5HbMvGXFyCKl2jciKMqDJJaT47JhK3Y65BV9NJ1+
TgagP6pMx6eg/c0BzN/zLv7DJaaZzFqcCZTiPr4UVlIyTnWzeVP/vTAAQe6txEFX
gAvwmA2ytQuR2hrMWVSHH/5h5rEx4pAJU/bQjE85JAHV7yEG5qek8ivmbIpGlb/O
Yf0rqchM9wmAmkuQTuo4xJ3B+FXANczP1arzA+rTD64TW6x/rqwGPO0nFLd5EDsq
gXOQ8qq2eK5kGhdAYHt0FbWV0Q/3p+bj9dVE+/we6Sb9rs5x1+vTSHyuRsKUzrQg
mFdKV9rW0bPDjL+GdcfI5uyhMz+lp5MXlpMnQwy2Vyaw9TJvvxp7tftFqzZNy+gF
rc2ownteLMQq+mq5N5tZbHABo9+aRUmhMjLo8KvUgdsPgxMMgAg6YORe1Qa1QrN5
aPrLi+7ncjar8QA0PsVVDOcUEoDM7+i7iSw82eAZzLaYVzIeo39LuvOjrxl3zpf6
MfTYqCWb30kWq38ZtbpWdbFX2RC9R+bI3P3aoML9c/ScyhqwYp94AAFe7seK/ICY
Odd3zQ5B/BcjkESGaATooAGk2gceu+UcbrSKvacH0lmSQbM2x/l6KNcu3UVfJxHy
YzZPk6b1D4NufmYwztCBrZ45ipDQJU4yRl36vzuDnc6LFerHjIVtRQV9VQOELq4I
PCxrTmV9Ca+fnVyBN1/zYnHn88q61i3/mio3E9Rm5VrffxDhaGKShnesFJLyCcGp
u1kqc04QjVUHuWIOajgdApbXLxYgzsafbqsLLK2DsmaEPFenaCmIHnqNRqtiUW6k
HYNz48Ryihy1Pvgar/xha/umZeKLiZ2pa5hxIbBVJMV/RMaMdiQ/3NfvkCtRDJfw
REwOccwqbqoyrRYRWlbAWeixz3rHfRziZWa/Be9G04ZHevgjiL2jtxqG5rrFeaUr
Kl1My+2ESmwXCQ5P+/e2E5xTjr7/ePERU0un6tnZyzJ8zFjEta67gZze8jcAts4r
L69XAK9UewgPGP4C38E6if30Z/evINxEQR6VrUAy8gdpDmdjiwMcZUGWL4jH88PM
N/yJUtuWqYH7fGuiruqrxhF+86BoGEap7YMwsmNz0ZGiE05gZllo8fysrj/5Uh9N
Fo5iYaYdLGxqDBhqLKROJjFjKhnpJYFesDkMlhyvDST6/LsUgRi6lqO28AEakrPY
gg0RXQeapUkigkSLlXQMKlMxFJaFMLjqTI1xq+c5ldO5N46qVffMw/1dhaLlPc6R
GSw8YnJt+flSnJLFANcgbVmdIr0lDUgxiYn60s7taGbvPRLIMtXJ0+VQb9wc0HMy
1ClI8S6u+7UPZrUKuyZyJl12qjxHj7pOs6B6xWQOkG/8mxcBzR4/m+Hpa5WkH1Dm
9a5CGCXJTp7AlgYskfvXZ/wjs0Gv9PuPhwuuIJsVBNNk5cmJoCXzSkeJjBgofZ39
KF62B4iPvOMdf33mt/H+Zi5dhkn+poumj4kEMvNCuxQ6U3y82L02mEks6fCnMynu
niCULxC77iRWLo17UPbNY5/mnVpXJnbu2xK25SqNYbPptc7vqbTN58RWppVT3Xw5
pr9LsdH4xJTQG9n09CgHiOHmYdtheC5SS46YB4kURWnyqyPW1CWsSUf4Oh+nzbm/
v25n7kp8J7nh3wgtMN8abnd8hFoqTgtUeFaKKUH3kJjvdu4xBW621QTdfrg+km+J
aAT+Mj/cRPinnOCcIb2Bn7+3JyE10qhLv4yQvzzT8GhEjsUc8UFup6AVh7PmIbrl
dogBAfKSASn5OEVT7P2XsYxBp766S8jfbIM3lKm34n3lx4vtod6zNQq80dp95fi0
4wGNApaJoYc6h/mVl+K1os2Qt6KBukd1MqKmoHHjSSb/FnucFbbaTmG8LvUnKWmV
sgYIJD8Gjvi5FDOZ4Wqk+kbe3vcMcg9+aywGu7eg952Vhpym8cPP40lrexxV1mAQ
sfJmmdS/3ODLvTUJFL3CN17dqQwevtFJWNmvRT555q6P5Wr2Eqqv6KkkeftWDLho
tOW/c5hpdg2iyKEzE4FWEsr8r/Io2tpzbc2SXxtXha4qYpqZKmzwU7eOIbXdxVlr
ST8tZJCnNz38+0h/gkhzdEuUBCrm1nmVgUkLc15sfVUyQJzZAMJLqGOf/iq04JgK
0UPiHJn/S1cQJS6gqVD44z7oJBb4VAomXKfwvNv/TlNoc+YFbemp8BKTCiqTR7eA
PfsV8XVPr3jr/IklaJAOBy/8YSiyNYhbQ8hp/pS5YF8QziEYHD45YsoScLEK1S6s
X9aq0yajKja9GJYnPscjYVAUfBjZJgD6d1g5WSVYemuTbeCPk/uW0m2Tklfc//Nw
lwzKF4JbP7XVQqwE08+iPhQJvz0vvkCOcJCouzivPefYmqNhda0ZyWdJTSZ6u0zS
zbRj+LikzJb0dH2CTgVShSD9LNuL7nVx4oBwLBOvNmt5DHHolEDzfT3bXzv62kH+
OLvKFaWZrvZ/C3VCdwa/PeO4g0/iGu+jfKngmiUCKWQ9I8Gd8Kh+CjNRtqMxzgOr
YGaJP1N8izQfoPuktKUjm/nMdFPNaIAIpsCR3HV8ydo4y9Esdavo9NW24y/Alnxr
p5NVbMz60epoLzHxyKLV13XKIkaTeIInnvUGIchGkgP5wc9h3j1pLZyv/mT9pK2x
1agrysuoOsn2CC/cVLhlm5AIAD1FBXPGFWNEXGNhwXv2OnmOGx4FeG+UP4mIJrw1
GiUyKpHdARbs6PfEWYGmKIY67PiWo1A2hRRSk7Jh4EuMl2OyFhlw6t6HvVEsvZ5G
XlWxwDKUZCjH3jq0Jc6aA3g8a3R1i2BcWQfE4h4JbZzmNJWU7obZeHmEIVRTT4gD
IseuFPijxn7mFJU/lsMjN3fxO/mm68+V/hfgu3gsNbZw5OqSMIycyrXhWSZtd06S
YzTJx2wRtSGyTQEEW2Y1q4Kop1zsg7T45+qifil03egghnp64kS7jvt+Z+1oTCDU
67mJBhN+2I0d428bgITXroxJ19uFeQOsqKiLhhWgw1VNlFxLPR+elCw/tKhCxNVu
MupJoU83dZS2wArOMjE/GUX+twsEdT2Y9Fiv67UBqy15cg9ebwFEL9JK7V5JFHi5
LlXdB0LrqP0Si+9hUX1MK0zStmTEb/h3Cuzw1VoPJyvkmvuGulk/wtGbhxTffeNT
3pSTuKf3oFqPZiSb2lNXmNTyUqFn8zMLmrEtxJ6NVDshLrgiG7ibNVu2/CVFsKET
sSrv6swmg3yGtgbgHjyEovUBeBxLRsBYPGeZ9XiE8gYIPpadIM0hOHks7kXvBFjp
8mnAEkqu0n9awE4L26gb+U8PmbzFJNeCRyyeHcB0HzRPsuMR8H/z1Rn19FiVi5q7
t9WCUYN7QnKDXjQhwr9FI8UxyrbXkeSQ6ai0sWKqkO+NXA8YRKVe15VHanz5vJaP
jWrWtjSwqgHl/WKaw1qz3afb82K8S4UA/4Zp2xoBg7HjW96/J28gR1mnAMt3J2C+
Yz3tliSo938rxgK2yoL7Vo8aH2YYH2aEnkqbiEzopHWMUG7mHPSJRIrVVZvO+PPo
c3fBhtlRHpYGIJF3Mn6dTkNgHTH6UwKaBWgjIydzaeSc4yeyX1St9efhzrfdjJVr
+Z6GRjnqfcbKzPnMqgrG+EXkDokU4JnBpwocQ1eGNUuwQ2ZfILIT4aPKcEixZWDG
+jX8Qwz7P5dOukrrmmBDIBZK8ATluC4jZna3sVJ6K5yBydMD52uOC5izQf3WAN0i
LiLiAcI4V48EyWYpLy4wi4R1JNjF7VJDVpORJpPeFX5Z7cb3C/yGR2jH2ln9Zbyk
x+YEM9Lp2PNeOWYqo7teoPxB2nRnr62gLhpOr7vxpMPbhgM96w3EunQz9MnK6s29
3eiX2DzQDZQ88QjhAxgzYehCrN8Lz8DUGq4RZ9dZbKMXSCzhPjSDz+wCfpzfOWQr
Of7VxQTiPLE58L0YHXJugWGZV2F2dbPVpqoLtzgOIixcCDCRszJJi/vGMbDjnTjM
aqRwpaz7wa6ZuuCOWLc1gqWv8D+zZwPn7UqjzIDNQYVEr3T60ll3BRrVXkZYGWTr
7hVqelM6QtP87GTsc5pI5tVZT9e0dJX1+hWEZtZn8P7q16sapeewiG4BYzHBmGIk
JAP3E3ZxrYvfygHZVamwgWSB2RYCcj6FeWZxPewkjxTsb/JhQMhQkXFOUkf9DoR8
tWpDpyj732Gc6sbcEr4jb1BedR0Dga5ywqR3rD2z9vwfHVWzKwxCPnaCh0G1JefC
r1kHjrSru2nVmXw2n5Q1K7uPufvn2Np9bplTIPBhIQnhE5lPr6S/te/nsz+YpgjS
mB8yJ65OAdzCE0EeZ21WlAUcItvIDWhKiDGd3+tBdx8DaY9A7Ocyb7J/TNrxE65o
XPlpIMPsDAjSATMvEIEJ/AFdRSSNXj/02ZLhWunVlBwDBrWxu/1/Bp4BQe4aD0SV
XpS1cFZoJ6Py5kCljLiGHLO27Wp1cWJV7k8Z0/ceCFnDc0ec1V8DkQgySBHIxz50
tFWuIpN+Zjh2ylhJOrY8GcOWF2C15E2o1QXNCx8hMIye9R1YVIhDAsiurrzYMqkj
3p3ChYPioZgnjNPwm4WGT1L8yypRM3wdoPUeZEjLlT4EzERVednR/i6UqDCHkd0/
2iVuMcGRi1J4nmMlPmF2RDuKS/GsjL8Vj6E6mb4iU/SzT1YkQvqP8awJI4GOfeBR
IxsE12yWDqqRggnuxYCKgzM/BHAPgzGcyxw1YKXYiWkx8fOpoG+8NhuMv/wWPzt5
DKFeb+g1xZyE02VtohgQRgMugdMLgaV41SqVS2//h2ye/LZkc3mjwVLWVlf3G63z
qPfSzdmKLPONhiZUUBSppz9Wcuapu4meg1nFvQ+bFn8H+dK6+kaNE+gfiDLAmjFz
ng09N5go8CEU72p6ohFtLVRVgS0l4OMVcVVcqch4k3jpGU8+qe1OSng0X0wJx7v6
/2DqhsGAY5c6/RKQGKZ7AiXqcIdXN8wgANqHY0UloGwrPiyjx6r99aaoqIZFAJEE
GUOW5H/kF73wdWsIkfV+MZM6eHU76MvWRSwCs3ArQCpsO4c61+33IWyxWXRzt6Ex
pGfNBKxtIlP4hoBQ7MliRCNf2fyPtlPqqojQRsZp5Mp1jcW1rzBfswwW4C3Nh9k5
bp4zXqNJi5Iw5s/lXPTU8xL5tbn98U2ZDQGLnis09gNz2/H1qf5tPbi4lRKmAZSt
V2lSOrhaJSuqZbDutc7khhDOOuotv0NpK4FGUfQHVSWLhboMrOyDje+c6YQK+6H7
05DnNboQHJq802J2XACZBrGNpIgU8rPKfekUd4K5y+VRB3u76jwqbNUq4GHo9Ywk
QThzUyvWpq1klnoeNSD9uQlFwvzrv7v+Rrl9LnZ8oYI5V+5vruwm8ksjznydblWL
B1wJ9gOwbsTjvcrhkMGLzXo3b8Jwbt6KMQ13Wcu4VEPY0aOtmAYqvPojpnTboE4c
rlQJR4Do5s2uGTKkJnfMurrWVpyURzwCnRr4TeNIMMQfJnID3nyO4N9PzFT7vVyT
mjmmBRFaq4qtODlFzVq/WbGiz3Lv6A+ACAsyjbdBL8/24LyyhIfd9jM9aQ+kil1k
qkgi6FNZuG41fSLlWSyoFU67rrGrZK2WrE91rXxRPZw/FxCWp0nwyEvqKNQkMDNk
23fv6n2MGxgiOd2Qglbs2phiF6V3vicSntDe1x7ih61XDMpPOz+yDrcOzfv2HyXg
QJWIaw3jDWtvhgvxbsRPyF8UzU2vZ9WKDVpWUrvnySmct5Xrt4xpwfok8wO2gghF
cQNjLH/M60Gt7B9FEXmjmvBN3LUiR8XaK0dJWQgblmOnbvvTCQPqehMn5dWqyjOz
dGPkVfVTYF9PGk0uOsQ+YEuaP/Mqs/Hqaznx3ZpNu/lQ4Wm+6SLDEl15F6wJZjGj
651dRXRaZ3SOC4DOl1l9djakjZmAtG+6eOzRQdelz/bjB6KPnnZ3Rzed5D/iEPw4
6QaBONMru9GTRQ6NEwyp+F9H1QJmPVjrpmyJ4RYdQEvnIGoaf2EgagbmpwfhP2EN
5KTcvxYq7q52jM0tR9sjHQoGsy4VIzv2TfExFvOJtGVORfWusqIxwwXCi1o9thhf
Xu76MVHGkKwop1+uBKPEtrs8QR9NjYEk1MC1D7NFIN9Wkid9wUW7zyZmsW2EhSgl
g7iUdr6Z8w+DpuOVIahDNBPwurwSKy+G0pZqF0eAhsIqdr0O+rTwUTn4cf3DE8py
97e568EjAOjHRqPfWgBoF9qp7LZhjLxnOqOgLt8ZaydHisxx7xDV7chCuHO/ZWQ2
UizvS+gUIkLLiumpy78ien8/Hv+8dacB/IfXZzSEmrif5qPBOLTB3/d9kdguyn5P
eVV0utPev0hrZafTk4u3ntSqKpf2vbNsi7hdOlVdluPRrXM6fjAwNYkcOP2w/kvm
qxfnZs4/ksQ52ujaHF2x5Xa3ZRZCmspKAbxU6ANhi62wCCu+XifVVzzZXVKKTQXb
IVsJfiiWPIf4a/hfAjRMsiDcb3uAlktdzFF3TLE0BGW60AtgGN1X0VmIw/c3sahU
eSU1/YrpUITb1ZRBM84WVcSUCG0GDvEwWJ36oEXRpgXKlA1Bt2m3hnpwyZN2+kbw
pfNnbCE5wpuK6+PAQ2S4qdTgyra1Vy4coW2lYIK0455C1kEjhnEamoC0nL6bZcSm
eWuHdtf2/9GTy3TW9Y+wGq3wA31Y8BZasxzl/Y8wTvRMxgs5B0BCRRQAoIVq4XBH
NZcxSpb65KdC1MsEOPUQYkwimjBGyttpNJphGxMgoNeBA+zx4liK+ihJ4u4kyaPh
8l9K+9y6gP8H2ZkbA6RPcbFZht+4yBJYOSx4cCmJCOXRYkHUEG4PSZ9Ttn8tvrLU
+vXLXrBrjVQrgrDSh3Jsk6HV1f34o69rmA8I4heU6c3JMiPRc+OfkOdKEcpNYNIA
9ydw2b+FAzqgsBAAR7uTe5pPPVZVNYcBKjcFo1eqRrY+6JwVjTJecQAOrb6KDqb0
55amSFdRxAQM3puaQuFFFJpN0wyT26EA/stD7lP5Sb2TQxAK9oFc10iB82rtYtja
ROjABNJhOM1jgzzQddsM2f5z9usaM7cPJeRbmWkOTxj0wpEOarFn2nZSeVDh11d6
eED2U+8o2fNp3qTOOEDEObkVcbu3N1AbL3Oy4cSkD6+C/Kzrr5ehuZ6aivGYGxuS
wYua/Yh9r6ap+os8uQlFIcv8YcT6ANP6PF4ube0s31G7bMsdi2kbyaGpBCsoZa0f
5eFpANQDSheLgrqA6g1d1mBHrH1qi/r5BHoYzeOfjx7Vy5eKt0RueOHNVeY/cGjJ
soydbWLFDMCf44ldUaJZWOm7ytXaJ6cif9z8AsEPMunkapmhY3lpWywrxU51FxDU
EBDfFVB4OUEiZnfukfjhyzVFzhJ1CHpCbzR3F/LZt97jOGdS2Xdq7DCBn6jE227W
xZ9Fs+oHM+8jXR7FwgMWCbmwQcvlJuuMhcImxs+lK6YcWAmV4P/vgbe5VEqwTJq1
Vq8GpuDCWqdEvngjtWs3GYHzitdptaAF5hGwhQ9GzPnOVP0f1pDDMo/TgFOKRmg2
98x+aTD+E1MowpDDGoLbelesxRObwb/XQjVFwvPFmBpxExaovIMhRWWZ/0Fweq99
8bXlfRjo7P7kSE87EfVBzfQsDgHR/ViVfdY1IZNnCRHQ478mEPUNinviUm3icN2e
ForJ8DyYYrbcqBtbmo65q8sg8dzddNUhmNxu1/1DIPYOAu5acrSS01RTRLSFL/zZ
kr/ZaAiZCJEBGYh0EBymcWZJJtsQPqCdvrw3muhr+fJq9uTbPNKIIc0oDqKro9FB
lHb4pJqxvgosWmzdxLxqKu3EPDkt5qY2XR5qAjU3Y2qQH7fpTcZwUbuWl2ylPBoP
SI0pDW/IoZPQcSwbFlAFK3NiQKTaSrKWDkMa9pOFbylrCLU4ZMh3LK+2hbsyz2SC
PjR7Sed2j0j7TZOEeu+hySj15gH0+IwSyu5CVU2sNzsgif2WGOk9CLkhVUTFLxlE
cDZkwRmeC6t4XhUKYehIu3x/IRyLD+5XOWyjuTii7OM6nFgkvltsPlZZj6aeySK4
sXHnamxGB2bn59dewrT+EPRQ1JxOzRis3SFtXmb56iFiwtqvpk1Z+W/w9VeMM7SO
qCwfxHWHaOV+Nl1IMsdT5n+WZ2dhJQIoCSLSBu+uCoph5V7YEG36LnVxj/3TRe5A
JgEtf/wpCWyL//iGouIjQz5txt1p/3MjYFia+0IWz2//rhppexEKGQzohs616+i2
pZywbSFWr2AzKgRW54tK9X6zIHqFJXGZ2HhfwvV28MQHqS4Y6oZQzUgxiwW++oUj
wRJT5krFi9BJvf6AUFOdjQMpmJjsz1hPpP8N5sVT5mkU+23U/ercu/OdNO/dzdhc
SLLolft6EQYxCrmI2UqjLiez0ugKNVc8iRbbhqQRmVNhp5w/jNpl4xBuXMviFy6q
bbIZJwblobHIht/yjzUSofqD+g35LSK9A7h8ahaok6Gz4xxa6cC+477m29BjgeqV
wwpDRGfsmS3+HsbaJsn834070rGUOEhb0bS45e3f+BbQwjhG6d9Mv3o4LOx960Lg
KPzoGmjJ7TNdkCkkV7jzSEscFyZpR8i2TmJS3fR3F4/d2AA9pSZECNWh69ISmFCO
4G2JTKtxU98ANg2BHCRpPDq+2/bpywOPdVNpAGn/qFKUTOMTuzlbdAFdeLvTTE1/
5FqiRiDslKZN4l0Bm/Jx5q08dKLG5ehbxxmLN718ezONCXEiHy3gUB7rWUX5b7EO
TdfmI4JpXHkGpPZxKURjR+lm1HiD3PiMBUqXBNxAZxZb5F2uW/PaalGFHdQifrHd
fevc9UgRREyrjIKkliLdADwwv8Dj9LpE6edLoynJQOW5qyeWIMnGUPm2hxUYGyY6
epG09dQ9Hij0IsIUu7d3nVB/7T1y34HPc0bqfsEGZk10CNXO9DzPYcZFMes49wDZ
DI+VLdS/MvRbJnzoyw1YIwqo2WQBmifH4HlGFaFj0PBG/4Bu0Hr+6e8og4prYDyj
z977dfpuncxRanH9Ki6CzR3sdN3Y32L6DJhS5ZwpH2A5SnzsmIokqdAT5ElOUExF
FxMmdcRnUQolv6d6Bdes62vWak1CEI1r/WCQv+fJzau/emXejz26NDhMxQrXuFU+
7PHTPXzIgqe1BEDO+nqMyTyXRde+76/uIvJs8KtZmqZcMw50YqgMJhVHzyOQqFVw
ejb9n2dyJHA9eV7kmR832GrJtczfq3gac9mxQjEsaW09sr8sHRJsSTD4vBKGUYwr
9D0sWi15liDbpF9uaLJAW6Km4YYB6Yg8wCSV3ldEWVvFFxFjemVN66jGMn5B+LFA
8JGXZ4MREC+sY4YWVVrHCMAC54xRWukz9w78cxchRXmYBEPguqOcgAR1ZE/CGv8l
6xoLMa3RDQaUmHRcZs/hg0kHtZHIz6xBhRqs8+cbj87I/PKjrqxexKq4FlwgUv0x
bd5jYUQ0i4Bvg2RcOPLDDZVCM2wrC5zfcipsK1jZ+O0mXnqNJSQvG+59oUbXX6M/
3mAQLsO0LO9tPOydv4F0d02d4Gm1RT3oEuOs5oI0Z68Y8yRJrRXIQV5FuLa7KNv6
XRTZAQOEMDpoyg1FgzoRS1zwS0afsNAdm7j329tzD7VhGeFDLCE3tfNVcRMJJCYL
wS5qTKVEKVnv6UI/BoZak1+/Nzcc0XPFyq6mVMPEgyvqsYWZ/sa6iHGhsFUy6r/8
2FDpVcndhqk5GTD4qpX8ziQkjOmsznFquUhCxMGI0t2yM/0FRS/LkXQZbidyzRJ1
wv1EJHiy3vnNU93J3tTHQOChpACmhJMQmfle4b1/KXFh/MYf5uyLhK5y7AIkvMmi
5Ol//kKGfcCi0hInQdLQ9O1KWDwtUS1zZTrpPlxOqX3Eq198b7MP3qDp8WWoFqqB
AM4w9R5PnX0Se5apyn4ONR2SdOWwdyY5j1qBCMVJwVK1sqTIJKBULV0stafy7X+R
YN32e3Lcl0n5UA1IoPDUgVxtZOYO3Imr3EOZYEGzs7q5RG01Ij5wT2SaueouitfR
USROt4GIEW+B9B9KwbSLgac3JlFBjlD5IMh18GnFMV1dlZ+jGPZ4/KrzkeNYf7w8
xOrRnHw2OK/T1TdTRaUw+oWf0m48cd8WjNyE9GqJq8KbeQIMvNLOHBIG3dbbYoRX
WmvJ5byLuvxyGrkeXNWOy/f7bTjX+wXJet8qpC/PF9jWMwB1JlYKArInVJKoNs+A
fTUuGxtD0cRFXm0q/xn4O/8BQV2/GvoTRmT2tWltzWO3MqucPtB+RWS97Ezh0nrd
rJbFk8I35P3FOweRgP6l+hRonrYuJqPOYPVjxj9Kd2XQyWaKDDbeNeB2gYEV7mkJ
l2uu5DJBHtiqggT2aHiL31qTU4l7UFAvuf62cy5r/WVOjqi/0hb1R1to9T0mxkG1
Tyl2Fhk40v/0FqxQxIhhQosc9ckDPIz0d2eYb17UK09c3SWXSexst1KUtO4WwC3g
2deCdoOwziCzkLZbrKpN4vLOCvTV9B3I7MRKK40spFuXJurLtVk6X/ltpmfkFGUk
76jwSgkn893JcOlo129PnHiO94Varu4K0ohPwMPBG0wHRfFOH++h6H73+rDItp1s
qmvHjZp6ZfPyiJ0ZdhqZ+QHddZjh/XLxAonKeL9q/LOHD8KFHfb6WG2ecatDAWW7
TtxRuPfyol/7uY4SNiQf+LgYBqpwRGFVNVeA22Rpx1jemjbrGg4kgFDaJSc9MkOG
1v3rwVHtYfsL9/34s/Prxq5ctn3CiLvniMRNubqGsWdXq1Cq4U+u9AU+zcHaja2V
odC/EnViW9i4PJ/zVLc+R7lY/jjVOFoI4UPiAQJ7urVRCVUaxqx8c6YODsasAKrD
Nz4jhrmI47GUxYK9FdqwL0p55K5lOi4zUTTeNvpm9158bGYFrPrXqqhnV4JJ46mz
ZjuW9qKIYfyBMfVgthTBjNUzm5Z/IMXykA+LQp+9qmgHdGLhSOZGkb6bmaQYiwik
3m3f37Ag/AaMBQgxk4ccStpLMYWi8NHCf1ZaG7s6d4c80eV50Gf52TwwMYmBuA5o
MQJc9IMkU4x+k4E+7L6DcfhaBkyzpXEmEDpTBei6/Me42iXlv7CGVIouvOcAw4+W
2mjRIGWVhWXhzXQvOsqC1nKDN6IyVT05KRucVFb/ez+ejPbFeIYM5eA1ccUUjtMg
aJTI8CCfJLOjga076in/CMKC+A7830PAmskoYNowDP6BkbhNXCVF6UvgE2uP+DiI
GYrFMw/CORZUQ4+IcbFOsDZLTrBkuqLj4Tn1TNzupZNp0yb2AAQ/MWJNh1ysrF6O
TF/AHQ8P1XNcRfzeJw7+7nFK4YVEqmuWBSYA6n16YIL1Zer5g9MJyU6g/uWcBSEY
zuC7Z1dH0GqJLnNFyW5k1bMYpjBhHB1EyE6mLIKnCNyj5+0cI/tYNNivSSXfgOnn
LdrxpkehWZE0gzbASEkWfOMFIEb0ibAqYcQuDOYH8L751XhajgBrrkmDPB2An22K
4L4h/H01LlEclmhXYEuoZgDkxrP62+rh+zinw8dQhUuaj4FJ5fWRWF2xyajIKsGJ
bXzgT+1prfl/W1Skd9Kadl0JvzFRv7EGResJJ6ziWon7qwUXmdElYsiU5w07Z0VN
OFYKIuDBm2vEl1MDilV4T+BVaCxUCjHhGknNf7V7CcMDwyshlZljVGqX2x5OwCON
T4tAi2YOa9GODCtzC0l9IhrVO/FcM6kUfDGUXIpglGlB9WZjuJP8Rd5A7KOg8F34
q/LIEvfn6UCXV3ohSIMnfx8K88hcA7GiAiWuaQsxdXo8JPnYwdQ/NjF8DWh3XImp
fwQYJ7It9bqPO9v8m6WcYh7ZaPl2JD6gylpvYTOS96h92cW8zZNtHVTt8us/6ljm
g2D3hZelDl+JK7HMOELCwp2lXZWlYDtKe7O+fqDL4undz/FL+HZSiNx1y7+8HSRP
TODQKUMg4GY8r7ur9jEel+70AzQ1jYHvSka7ZtKZ0QvtEfmirDn5Cl3MMRZJ1HuF
AGEaA9flB17liG8eBrSrttZuucSeUG0Run8F03WvcOIissCIWNwwC7X8gf4rYLny
ES+WRvyByfHHApHyI7JjyUJaKvAZNMHm2cHmd2pbdqmonsxEVlg1GwEDww4IjMkp
mulxddWdSNwRB4s04irSouWiHqhoRUSUorUp8fhifOXMR/sn81WoeyFGtBZYY92a
rgYDeZC2l2ETz2pXd2IgqEjRQl6Og0tW8puzu9686ZqSM1h2McgrQHgYd+7ZoGxE
07AOzY1vUcHXVVNf/Rvn661DUnNbs+RYyfzn/6a0A14ZVKjaYEOZtUedG7sfT27m
IQqDsgOuURLlmeVoTjssFrIrVjI4ZZ16u5noOwwOA4br0hsTKvKRGJMAY8JPTC8p
3gyOZYLNjkq23FnFl1EbKA3/OCpHW2D2Up/ilu2DcXi/8vgt504+bkzsZlFZaxRh
ca0dai+fPBKnGacdqO4MFpPOvjShwF2/r5P2UAeAj2pIckRbYGI2gqF6QEa4AUML
rFBViNi7jQxT8Y+XvOKGKlXAqDm3CnobYLZ8i1q7DzqYq2zokUmbSbsUyd6Uq434
m2MNYYL6SgE9rEnuUZeJ2e6nvJNKqp+Hh5l/J0f7NhfTC4QEoIG+eDBRhx7ln2va
T6kn9lmRKWGeI7m+V3iMAqNXEOHi/b8b+sd0DdUsdaS/Nkal3Efr1Qd+ZXXzJLqf
LpaGasr89PJoMbBQem4JC7sAYFLw4D7AV3tsgCzL/4x++WbeTZTrlUPZydsFmpK/
cCZ3d62nNXHjXraWWPJY7S4zXt3Ls2qpB1UhMG5PpFoz6/yNTftnFYFbRpyneitz
tTfKMnBnKpK9IJnoJJmafcIRa1iBW+L2kffCi2c67fvmLNTRSU6XVftw5PNkJ26t
iyhzOzeHaNL3g3f4CSwRXBzn36ZMj8lPNGxsH2uNTZ3XHCRYWHvPLd/E8yRHKAqh
DaKtaPgU0Tq7/TDM9vKZ7IHI27IC11EAWy8g3kiIbqNDM/IHobgMOO+R2lKVQU+d
AtphT+CyiL904dkYa4a1FQ6x8IcsqVdb7WkesSbglBOoeeHbSllUYFXehV80KkuN
YjPESdNn1PxRmGqWEArrIp2WxH9RRxOAAoJky+Is8QavF2YSF7stMTZ2JE5hEuoR
TELxdnKJz2EjzENeNRNy0U+NopjohIuP86KxRN/l7fXOGd7iwFumLejNkQmVrI/0
oA3shqAjD7Xwpe0OBJeovMRk6E9q7QGGM0fE5TAmqHz5cnzul5P1yf7h0IhlL1NF
nnk+MVBHAH8yQlQxF+aWyS5UiDS0wOJVtCrW2r4TFUDZXhLAhiTd7wwcpCO0K9IV
V8u07frrleY8oyuhvGddx6H2hdnZZA8wAPHxkuyUt7e1XhK5TvjmITHb3UIHi+Qy
LjhypuuUwPb1WZDzDEsi8eKjLXnvgw4+Taksjy8hj9zPlYR26ZLWBFJIzJ/HQJrp
JK6GDd1x10cyjgyil2fd+qYV8HXXz8ZhTVMEaOjoY6kbCxrOhAtAopTLRsIDp6xl
/OSQZ8dzvZFvwIGy6w3eRH1Iv+C99lBpCpPAf8Xz1+URZHZLsV4r80zXHdQzAxIp
TRkgVaUC7QzEj2ykI6RFoMSVc7Hrawrz2wjXrYxy9vM6SCFU9x+EXrHm7KkLs/Jp
vNOV/eD8mjdC/Cv9N2oh1JazLnjhyP3TSpgksVnq9et+hzbXkolmsk0BNf43aP0t
RmCUQyLU3MH/cw1Vffe3u3AnfRlzmqEwAD22SeecM1gYJkSIBa1Zp1suqJFSPI08
DWRt2ZlDt0z3zI26RgxlksPX+ZN35qT8pRpZ95xRoPxQ+PXPFtoR4GdK1KFjdA9D
Iw7UlItJsqT6sUZd00sMNvEk4W/2iQA9udK94XpBWmUJEtLC8Jn3iBf6gunPhDda
H21RRt84trd02z2iv2CzIE9YFgM5D70xnAYT8zhIV1xb/VJIpJuoAE/iIrg/6o4x
+HMvvdNjDTRjj8y8HLy4mKUItwK6L59juG2mFmw2GhYUd1zsCrtqPCPzLStIV5iV
PfZkGaqp5yduPoB2G5xuPDvQaM3DZs/Sy1HvVA4vPNxmQ+vaIK4E3IWb7zoJxr0H
sfcJtlk9V5vi/A0vLiRhm9PGbLu3krjPvAXLUmheptVLdH1YtQrKvaq4OF49lxBs
hGEQM+gVVeXTJxKPf6pW6bR9lGn9e/INtMDvWVzxEgQX2CuIFz1zuUQZpvY09Py6
8Us7Ran0Dw7bc6t0tPzrcYAlS5roUsGC3RGnzL0LW+5AEEsRQqSxOA3raPMPAjHe
rFcnQqqvHa0fvaBQRGqiaYL/SBvnEHzxCgtD/5EUAIB5jxvdeP+AlR5gzH2hgtWc
6hyVZQ9+DpKkx36CQsdIRS+k1IrbDCNi951lYkNG8aGz4ti23yT4dM3Edybxl4Nj
rcdLCJ2791RcRtQC6bZcITHvKkmJTKnr2A67NEEzApbxH+aeKBFYllidGRTCK9GQ
4wHOumPkIiDkzZUhtA5ULCUpYMkI/+ykX1iNprZorCZ6N3imCkajoLQt7KIrwFu9
qTiAfP/bI9iJihF2oPiKD+PQmbU5XKLwRcFKOUZdp8oYfJMAOb4wU7EIwx8Ttdb5
gIaqTuEwCfz6nTAb48+RVmnTKQZI/NrJeWfSWPBBdngyowdbLzwdAVnF6arUnxLK
tKmjkNj88OwOLN/hvCwLOKOrJNvKwW+q9EEEM8d6neVeNQARH0l7k5bdTt03RPqJ
h6/9dNwIbgiBR33bDMOciNruBdjMhAUhMI+GnGea10Tu2LXg+cYSKBuDcgEsZ+Hs
Bzg4fVFqn5XV0MXit5VVa2bONnL1WxHddhp2uo7+1ULEPWylO0QbP75sNVSd9n77
ONlf4Qsq4lKlxkb6+T/ZrSLOVLNIKw6ysvc74Qe5+lqRioKQrUrpiXYZlyAETayR
/TRmxKs4u2QhMth+Fi+bCYSHAVOWbxggUeIGmU1deEwAXcGhxVpByRYQLgZ4be/0
aAMEN1LcrXTxOmFOAUu4Ay1FDVHVTlr9/2BD7Jx4shN2C5a2Jm6OyXbq52xRfbCn
Df7i/VsdY7bABVViK6oP0h9Vlt1XfGJxVGnbT/12qzhg9krFdZy6hxealQFQhQAn
3grrWGcJ5/+ZFH2le6oIaL6a+8ktZf30U63pFQGb2LbbJhJ7UzRmlHEBhK6RQRNL
EbTViNDJmAVbyLRDvEbGp+/RZ3f4VbuB+AQP7jtGNbJmcYx92OX6/x/FJxNeDVpm
kieozyJ7YTh5QW1sAYmOk3MTa7Uftpp6onSGLzqP7yEHVLsKp3sL1gu/+g7SvIFG
ROdS4Q3GMlp7/6jO22LZKotbn2T2JMWf7GhUg8ia4Roc9jYEtMr7lEQW4C8G2T8g
XbZAL5lGfw5/2BBmdvWX5jE7sSHhlMHFvhgzeT1917+5xQn4z0BRYLIQzuh70IC6
LTMrHHrDAnjxg2woNA46+SL4GZzyuSR++8G7FLtNTiatyQxzcySB438vPiK0iWvI
P6f0HCMtn1R5oAReGVKs08A5MYb2JflcXh+mUmSEOBr0E5gbsqWBydDOqHW7JT2t
j4+P4q1fg8380W0FSh+b+9d3aOkqM6CPYnfkgFY4RQBR8wBfFcOlo3jNnX+AxgUU
4XDU+bBl/GDHWexUxzqsbkXhi9yTFOSI2oTTZRygKE+omqDwe80LEXnsP1+yQirC
lZS67qfnKI98nUgHxIpeU5tOnZjYXUE97gbrmQxSARwH5n1+9+3ZEfWBCfhWwpFu
U+crv1K95+k6UdBA6pyXbtrPgHCtkdcZh4W+KHxBDY7dUAScCaRxzPFqqvfl82nD
7IBt4GbPn1lAPrpJfwuoswsAz/HqpKrx7QNOAiK5uFFa40nu0m7BeliSLXPnDvED
tBnYKPBYMSjuGWyaIO0jUBfu0xonCrWIg1t5yNjIXiRgk+AwTT20AUMbHgXXtdge
KoWK1xtbofM6p4d/yJIYqrqDkjmMj9WdQX3T1ShGFEHOzKhwwPTO6x0UpYSG5C9N
TIMB9h2HVnPhto0N7TYbNj2ruWt/iINrn1NF501itf/MNjMPnSxHCzFYYtzcTBhL
qPG+yDtZZpNo0wqhWkjAqykQATrdC3QzeWfo/DmQ8LatlGghukq6gJ9Q84ZzcqQy
EoOO+FbX5wWRztesN1z9BCC+GYKBKGh/Z32Rcki/kiAlFx7A98x7a/pfwzvda1lp
3ONHbL81G0VBA1M5r0NZs4QDtVSZ9Aw+N8WjFKbCXmn2p5szIIfHfzb6qxn0LRxc
NYPnmkhRq6PF/BADQuc0siHu+w64JH/O1KrfIHnTGlU6vx9m7Ga2HX7X26P1XAIG
zVCmR2BoT2A7Y2V0wktI9Q==
>>>>>>> main
`protect end_protected