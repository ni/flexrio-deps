`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3824 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
LfLaKOw3utJqtz02pVdKf7i4qQeQssv/p57ETXHUVsmpIjY+QRFjkAIRYMxSOt3G
wUrPhvCBcvoEIJnA3W3r0pQ2N/s6BaO9AVudIdDM7ayXQQ7Mn6EqmKwVbfvTjYSm
XGJHOHmny5pC8drRLwPTsZx1xD50sYkbh8q1zx/r9v7kiOg07VjBi5WukiBYyVSo
S6lLIf2tIiTkDMXZtTIyhc2kkWUZ0HbGxlnctWg7P3vPR0g9H6zXWFJtxZ2ZJbkm
8w/OPq3CGqCEMy61jL/mklsUTZT0OaLsC7+5ZCUFKASEXL8pbUXy6HcrwGdbtS3W
X5ig9RTIJ58gVPDB6h8+BQiIz+dQ9acJ7SO+0YF2a6F6xUkaU74vPBy6ffoIvbZ0
BlFhGhZlfW0LQJg7RAo0ivb0xSCun15a770Xot3KEMmFu75Ae5xbCQGXAucX3zKu
CfOgLYARYvAmKrunIJebwdofI7W3pxjZ4QZUm9QaLlYukBzFniEE+DfsV6d5wt+T
EN2jgi7Hyx9cAZ+if1KPJAOmxH5ZlujyvvYoJ0QUBqGfYDEOaB2rmxyJRa8xQrhY
OsHRES8CtzwgOG7BHnyF33UUUe1ZcfzzJpxZlPNkEH4DjFzA1iy/M+SLcg/bIc2k
b06FwoLTTTlLoI+SnYR9uvaEPDLX5mlrZsfcajMSt4FcedIyqRe4YRa2gqTyolH4
+zuEDFrMdj+v5WE8odJNTbAJLDWLAeqV+RIJ062mwRDKUASRd9DSCkHB6LgA3Vei
y+wDW4hNnEYhM3c+IN6oirpeYcD1mkQtfRCTzp7BQdDE5Hj/2XnPD3fucEUg6XrF
azkAaiwuFYHNEZu9/dEliFwXthTsLLmKGq+HXFpwpoSZ9QGaWKZy8gFghzlmJgHy
+AqgohqbPBG1qYIu39AspFnszkSaMtDNEpPuB+gNGTfER99HWQdq23RKjTmS2N5b
6FRepUtCgGNV+xjg2zE1z5oaVvfpyHbaz0Ze1oSxaxBcUMPptkbQT6jS9VF8HaZ/
Spw4f6nR+VEJv9S6Uf3zZLPzClK5jZ3gO86Un0GV/3gV2XB5U9hipWh1hLOjBpzq
J/I4bojky5Z1JbxaXyTB6AQ+6QGZXsvUydxGNzw1mgVpcPQoolTF+WblIXDkYaS0
PX0rgNJXqlFsnRmrcxWr1haiff4meCAaQ8/9/MUYDNJUVyo49wiXHuMgAFl2DTAA
Y91jCWWoRa1gYwZrTdterOAcRf9fvSNo5Ltjo/x5KPRi36LWsNtyEgWV+eHLXC8B
Cznrzhl/fi12J4pQJGwwQZTYpjHuEfD1liPdBi+JM+3qT5vLrYMi02sS4Eh2TNTZ
bqDndhkQvgXQ97891o38WLpIlzxp6ZTAMju/gxALGZzc7Z7ymvlwGeCzBBx6sK+i
oaYfvdpZSMi5hKLUbHMy4br7iQ/VcPud/csVqCbBpsJRgXwH0fuMEcnNaFsWSv6r
dLafqeB3BaqG8+VbnY5seRavMZaoVk4idfJbTZCsGiSw7dtZbk5L3URbiPBHTDKl
6EPHA4zYPDEfTaBOF3QxDGg6YisWJafUR3gjz7s3K6ir8itEVBqIjscO2munphW+
qrdjw2YYuKNXQ+1ds3GovQkltuXhVjw7YCONKzgEC+ATpoo5SCS+S55v9LdzIkwD
5jTW3pVIA+/HJrNmHCO3r0Bp7xeGOjO18hgiWRTlBfL5A4Jmgn71ej17w1zW2n7B
0me3E7j4tnoTOzbHQinYuqQ3+lUde8NlzMWHQe/KW2KASKo+k1WfTwYRDOK0Uecu
oQFleG+842snhiO3PE6BMaTAIkUDhrpZaaoSF4sTKS/dGRpoVZwLQRg4Qqr9Ivyu
c6MbznCzoZPLgd+6ZUe4o9la0IgB8oqNa3K1pUCZYv/lE49q2mHz8kKfNyIkFWIQ
kQKoZbXN6yPPLZ35pTeCXK0nqLtPZtfeEcH4Ckho2lDohZFYdUjkHXVIgTkUYQJc
NswF8cTWaYMdEq+VPIuvHhBTH0rS5UB1gYxckHi/awCtanZ/b2A7uDoIZrZYhbBY
R55LZSHXmp6wQyaHul+iE6V5uB/9u+jD56XlSiuJSqxRlLTtnA46ql8+AZQvM7hd
Nw6pU2skRA7knwVfWp8u8Q1x0G2xKG+HnLpfbGV6E+wRIgObjOqQAwY2m2T8cLL/
Kh7gFBzLb8YGy+de6M7r84yCptiPes9OswtU508iYNhpr/GyLj6MbjEzlrxMab7h
bxoc8Wy125WdIF6ODUleKRiFE9brVXZJNSB9sFmhHyjXrTjTrFJOUvSioATkjE9H
kPCJXz4DUGwwciCcDBTp1B+vKFa4RIDVz0Y/dY3pepTtW07d5uoMEj6CLi2JLS29
8/x1iDv6Be+OibLDbF7plYZ+MPJB/5Ho78x3p4EN7kCm8UnjLqCinjDPduoWSJUx
n+oIGoe0uJ5i9eJURI1HFbZmjkQGW7NWsmS4OPVP0vDIQoikqpGvdcT8UIuUm6ZR
Gsv3KUNAgGO10LD/HBbrwCfhKw0ow+wlgxWk35QxkVbJUHMg/XaN9lBLL0n7hkei
Hbva8PSv74Mmyy/UaBBLhtvVSa103tzY8sY3c5GjreX0ZuL654ksmOuJCIPv1gGD
YD3uTk7sY4H9JG8VNC/2jzRF2epkq70y9oZpBFvo2MSCLbQpcYfi/50LTRJkCQVs
dIXvwmZtFfDj+xoqqUn5zG+OV/KWsrzbQbRsxfZ+Bx3h1KgUZo48v6BattriHimp
TPTbUmJ19n9GOVFtfNV7P863KQqW8ZzadxaI2bvC50FW8X1UaryAvhSzWX17M7FW
v7MQ57CoCFTcFQR4t4NYFmDYG7iEHxpEmyMNZAK7D18to/0z7TgAOtMDeS350KYk
47F/ZVNsDzHi7yQmti+10uLYMHrXo3qQ+o0RHkO5n+lj4egLHzoqm1wGUyXK8GOz
LyY8owsNhyWUUi33li4vFAOVkBsJHGMo9M7eCz2HMb7Vl8Y+3EZlCC1KmL4T/750
EG25u0ZBSp1DPhbTCgt8W39dy5BiLn958d2vhA4FSFmhBTCi+t4tL+ditixWb0Ww
XRiQNlJQgrHAw6pVzNwcBOynHhAyP83CfPjG11J2DGQf6rquKM1nzio+j2ZbS+yR
IY/vN9JPg/B7QvYwmRSJLReXgfv94V2180Y/V3emh3eLgWWA3y+AxhcjjudK3QU9
qiW2BMGxc7TuDsRUpHQYpxYxJ8no9wz3M6hoMpYDsopjjFHiPOeBt2HDXQNWfwME
v+Md8XKI4UKDZOvkpYV1gS7rZrE1w6EWi5YCCec6xZjUhqmpJi/5epxN4PSo8uf0
Se1yKTYe3SySOzWs7H/hCRbczuduJj/AdH5VindVtN3rBUUGJUeYyJZuuu8NI/s2
9Y9Yvm+wO5MxMtGprMysx3S9v3uGkdvRby7lRkmfl/ecMdPEOKISI80ulNrm5YVW
Xjb7a8sH1GwxVSZsu7FSuQlA9cZEgYZeIy0T2cmnhtrtPRhYsh0Em1vbSXzxLFUd
CRKrxdE0wasiOWatcxGcR1ERKUiZJZeL3YYeNra/Sv/63yPyNFRV5wtm2zFvn58i
fkCD1v4xCV4J4/dr2tdFnZGkD8pqFrovyN7Nt1bJHyQCgzQCfYI3zszcHGBeAytD
T3+WEbhSaIWYdlJBDXK1JXRQXEmdBfX4t8SUzkopXKc0vRhUY68o3NhIZqEeARcG
gvM/619XP0BfHtbju9H/wZ2EOfW6n+8kC/vJ2ke2RJsnprjYjcfYIiirPSRgC/YC
FEojitdcGTuYChW8u0SDxLGCEEfU4AeZIc4dsW4/EwTz8G81eb8DK8+TJRetIHvN
wPoP17f5lOnOM41XL9T+V8XOpeopmukpxa40GW8u04M7aYyppVK7OSGkQaiAIJ1i
jSJcXLBLjIHqZJvF5iTUTzT/mRASW75uC6kGy5ADIqfQgl6cpmoGlmKSC1vS1ftu
Dj7oO40EYyOUxMc/47kRQvukg3UbojVKG7GLiDYugJZfw9edqEBeTJwWDRf+ImHt
qVIK/wgmKmM+sW7WiFR7ixOU9xohqFK/2HVRRxoBgq1+DSmvkUEvFLY1G7j42FMZ
dlvn8UDrnDOyWT8BnlUIRz+mU00x/3UaqntSDOl6T+xkXFiCEUUiGl+BjdEq4EKG
CwCDlgybX97oPDy3Uiyn2l/dhBTbnktL1+HVR+MZq1vo6tH9nvYvkTeApluU2wjO
7O6Vixg2bPUj3JEcY7gox8fGNH9krA25hPKo43QReCtPi1GyBIg3oqPOO2T+LX4s
eJ3P9jQ9TUIrPu5K6slMFMmD3PEr6qpnflUv08N+EtSNdIpW+lel24ssvOdfJZOf
HF0VuMogp1UiFqG7f2s9JYR+HS969aU9D+3loDpmbz9/zxpfALFmJBSatzSB0Y+E
2qqpatxUfPjs5lLjeWEKY0XUBkw05xV1eF9NOb5wU2am2bHLJYsektabDPuGRSI3
2XiqYF759JikdI5ATvAI96bG2MvsDqq4arqJUTwJkWba2Z5nJ69F5zGYuQdszyH3
Pg+IF2nF2qzqFGlKobqRSWV4JU7+dhENygSAq812PElQBNLjNLB1GmJkSTaRUGPt
xGu9MtX1pyHbiNpD6syhlzvqo5QJoIk0ULHqJI4m0cHm9XkbsCYFPc9YaamyBchz
EN6+I0htgMQxXHOCMJq6uF2xT1JPP9vlo1EhMXWCajp/Cx3pOIoufFml7OPxCMQ2
iP654ze74tXVaaYSjm7oeDLKM3ybKvidbjn5obJ3ZxRvtSVKJZiC5bgojY2acwnG
+ZoYQgrpOeRrnNPjCXekIea19wRGxpTRlTNh9BgydXBpDbadGsBCcFHoClJWmKvD
lhYzuGiTDy0FIH2xwjfRKlEuZx9JRON/ElJ3U+IzOZAWVe88GJ6DOw2JqrwimUmY
mOskJqTSgHoZEFzcRPse4uKjLZY3+HOqtM28A/lvIwY=
`protect end_protected