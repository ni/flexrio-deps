`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7152 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhBNVMbsl6PTB5/ApNH6uD+DTAl4yTWHdDqal89lO0QMs
oiUFbXcPSlFGfo4o/eaCazoUlGAb56ydabKrt9PYHeZ0YG/vO+GPFN49lAODzTTP
Sm1ZI2N4qGSTeIq1lCpXFHSkxiQXTjhJIo5EzJfBMGIQyC09moANNYglVYv2yYZ1
2tySVBA2vZe/uGdgOnQgpcHSZkGsu80Ff1jw/+gvPE6fsbWj8k0spAOLseQtr4g5
ewbC+mLZRdD281xTHa5e41Zdpxu4jPcU2v2rzberKzsObuaXSVG4gleL3jTccR+f
QgUV9mQrGziL0XIYoK5sbsImggr6Qg3y2u6CKMnFaNHhjeU5U7SeggzfV4JE6ZnV
KHAbZ8xkDJrAyi+vNQ76hBMwLoNcg0tjC2fuTTRDal0eBph7SIHLl+2wgAlYQhGD
dHQwCtKfET+ZO5ZTftb3xZB8dkQkPMgegvRC+fWJ/V6+3oPA96G8VLOayRq3LeLY
pdAi2G8jLfb0rt2f8qi0LvUbyVyr4/UDCqC9ReMwSQMReBJ05kqrB18Bo6B5Q6Dp
GbjHfjbGhsrNsq2OIONTdevGelk+WWpQmMtWZJfDPZPDDyyx/c9h9TeSWylM9GZy
9T2znaZ3xzE7DQlmBgs7ALUiU3AzRqPj0Dsl/6P4DrC1ripaqRycMz9RSVIC1flw
jfWBWOUYOf5zvRdaVB+uFb4Xwt6IGy+8D3jQoKxt7H/bahC1g+sXHFyHKKO5zkEg
5a8TR32OdsikzJxev5vbyEq3WTaR8XZIcJFljGTU1DA/DLmww6tiwI/F8egkgRdl
zcQploN5XgDuinxNHDA5T6WdFi3xNmonuAYUotyT+bDb0eHiRaeO8cRhjJ24DTXM
EX/DHJ8snnSzuTLryxE7w71+5FgyXQrYCDmrhfIlXf9+X5x0xFzQqjmSAEUtU0ss
rb5cjlvMrLjuB7sTIrYYZH9MDoR2MW2sQvVhsRsZtbpixRGlNTXY/L/Na26gNWpm
2oQv2olfVs6r5pogzLSeGfm6VJsPkGnvQD4N5O4BfDZs/nzqVr0sVGj2H4irpF6X
sf2TSi2JDFAxM0Ya9wUS7kj1rW9NTXPOp0Wqjr6+Pz1F2XesfULP2CwfZIsWqXv5
vKYmj4eN66pvj6NqeaFVvBR/1z2d1KjiquUyq2hh5tatXv1tcO5RPPfV0xJW3tE7
820hsgrygy+jUFuToK0PLKm6+z8MOuytXlYW0vaxAQByNROLI9+PJkc0TabiVzzf
inM5mQC3VrFB93CzoOvOqK/qnkbsOugyfkLfkoTqCOh0aFE6Dm+4Y8YSPDDDezEH
96GQsZ9Yc9I+SMu+AUQ8mno6ZDy02TdWaaJgY+nADG+/9dhcqTLbeM8PG83q91qQ
zh1zll2osWOrN6kL6yRfjLueMKJI4HvmHH9TQbkh4pNDDEoTdAawb9mYG/8k1SQk
8nuQz+Vub/gVulogLbyH13/W0O8cRsN4OJKSy7w1NeJlWuMh3VPyZ1EfBWY9C4jm
NLpVsG0trvOwDl0kNIoIn3CZp5XOUiqnXwC/WKOX5S00e/600qfQKuOWPcUIdlGU
TK3FX/CGLmd40wDUvoUFnUIc3+iYjw3b1Ih/1QvMJya8g7c2/8ySYLPhBPevHeRd
2UediwbJafXUUmZ7AYYSPfc1e7BkfqHCtnmkDvFYNIPXV+YWIZfaVsjoIxxLLguU
MaNI65kcOv4kqmTy4expAdLNK+F81YFQx628hzs8R2qJqUoMffJOLfe6xUeCwkfx
2xhW7yxCWvFrU2WXtCatmSd94287iCOW6r4S/UAE+7UKv+Bc7NaPJPLnS4QigTel
zIpjPCVNmRlleSlwvkVV/MZmfQJdFHKpLcgyewEJJFwb2m0onURRWRzwXOLF4kVj
CpvGOujWxh3fWcsub1eSrMuL/0sLp6fh8NnM6e8HYJBy9v9FZnnqDQQ8jldiCSsU
LfGii3bHJQ/ttYVtalSEgZUIlDIqn5dlOQw4B4cZmrIRCabRXpFW73pWOLJN8YU1
BX41+AGlp2nI0AfetHjp9yhfu6yBHaGYFETHKNuwGC54auKEm7clldlnWmDCt+Aa
TIdSa9jrnccPzX38Cvb2TqMT53MWFejI9enbrPBIdjZsPr3IkHkH9YsrT+zYon3O
2ys1V2vCfnClnUD8Pui62MQlJIBiH0/8fhi2g4e+mt2a55gEBOzwGUi6XWIz0OGv
GGzB6UnTraLwLqJHWgVMbLbQYgba/7dEXTBwnp+3r1cyO9EShi6t/OOnlLkCJ+vD
Q3c0CI7LmcwXlV0TRg/vIGD8GC234CDmc0Ym6CHYDD26IOaG8am8lTEdi4Sxuh6y
3EE660DoCQvTAvgqxmYC8dZqflqKHoSvXDkgKF1fSy9t1AdvyqY4WlG8QOrHwD2n
M7Szt5IzEMz4onKNGutXmv28sw22p7uqo2abKSb41bsYwyTvs2+s2xNOZZrKVMdd
Ilx7XC8jNhWvJZUib47lq04OIbkSuHiji4euxdnUk4ZgtUwGXuntJv4SqaoGb+aS
ddkIPgoNFGlXpMRtotB7sIXDUGw5yp64+rAcnwWL14HeYhpBmsMvMt9Xo7imJXC3
mLO3GB+BsY0lZ6fmE13bx0f3HMUJZANzRdlRB/8oKAlWsfe1s69JosQqHzpwmgVl
C7HsjPrQLhOkN5QW8ONbKnSBtCzrUuoOho+j23nwDFWjZSvfWbXwGFOahupz1ugn
CFdQ3oRurY4WuAN51bYriSfC0ZzcMQOa6HeDCR5PIWvv9oVG+4nR8Ek+arlZzU2K
21P2oF6a6MTLnyEae6Bf/qo5+OIR0qkzRb9Mwy01fm5h5aF4wqEiPBUZyJ58cEaO
CtGQF9WEbP10i5l7h6aRfxM/Mc5VwBF3a2SPyPfk+wV3O94VX+FnXp+tpizsOijB
S78HJyQC0RopI8KTBrACkSsedkRpR7wt/lL8R5n2loplCf2sXXKksj+jGTYAIRVx
K+gywCPewBSBaMZhAtsA9ZHQ4CTHE8ujohmXU5imP5wwb0/uQiQmFlIp2EdeELhV
71BWFtbq7yTl+gQ64cu3fxquJosYEZZEgj3q9V9QwE5C3THuxB4pkRnICjTLJk5u
CD2w8OmFYt2fMCukr9ZVfst4Re+VPebd+mmodSizf80bcwZPz+xrZlvrUye9savF
VjKWQLAl2HohxXXbVLA6Qa5XnexF68NnP37Hc5iU+cGE9ijE6yowJhB+DAk3b46Y
7Kc0ERDEVz4dcZ683H9Nm9z6JAm2qsgysZm4hK+JHvLjtYWlOk8W1+4am8L3T0nv
kFch6XOCA8HNu8L5AkObQjqigToDrMuBrRJUKJWmCWJOguZ7iG8MQL0V2tD5mJ0H
dmOm2mCm/hMc6bYWX/aUPFt68uYPW1JVQfQmOWyozJJ2T330axMz4fYM2A9grPq4
1te+BgWfV/WChhf2ioa6PcV/vuGYKQHhEld2NvMB1P1xGlw4ut9g0rTxDyUNLU7V
0Pho0nUPfOAlLmn0CmC8hoAmU9fQ+yUsawdNDmYBUZJ+yaBOGaXKKvxmYumX+Gpa
DRX2p7mDKzvIqE7XEhIKzYeY6kwhZ6apfWZTuw7KfvUazaT4yI0JxkfALShmNFxH
i8CNwDsYRnKauxFq5IO4TS/+g10fwnNfDglepf2HzsTAiwSW/3RT/dU3b9v71VIq
aNH77cHSy2+zEf1CiiX06Pz5n8Qzh821pJSV3BSIWpkbEfnwwT65XyquagDdgpKe
+0KlNWsTSanPf04CR0pPRkcGyddvG9eWqkAXAAWbJ17BEEos+pwmWz2/s46O9JLT
V1bKNI55OzDttgEqvgHKi2KgSQODkVirusd3OSKDMkn/qMyVXhna2iqJ+UKiQgI3
AZtzHtoeGjytl/ZakvzMQm0hooGoY1wx9+JkNUM8QJv+svue1w5j3l/DHDx1oA12
bWbrFPOclO1N8eOo/JNF64riI0soLsaG+2GJxJr1ldg3j/Rc5C9PWft+U85TJl9r
j2QTGkaFMZsHtQZK+bGuGUJVJX5f0OBlyoXwdS12EjqBoxabzUgNdCRdSOp9VoZB
akpAh/vqhvYe7/OrqyOyOfoicn3D1Zt+ooc64JeHRZOMwH9ZWksdoIKZtAUj5Xwq
bLA2LP92xti56F0E6pREGl7lbro0sUo1iy98PSrtDY5QoUHAqRo2dDmrC/bKu4Q5
LvLfW1UxHc+VJXA9BTDnBhZtkiihluiGN3ueda44HCIHzhaX5Dv0xhhq04qGdLfc
AGP3Q5hV3QrztQQRVQlxKVI6STO22720u0HhAs3pv+FiUSW+FoSIPeB2lc7BytM5
yzIV1lOlDM9as8RfOkJugIHZQvm/O7NH5Wu6Q7Rrucm4AonT776/JScD7OItU/N1
6J/LCSxuhmy3WwaL/l4uP27jBe1iOKEQTIGMtUQljcO/9DtzzRFRXl07MtLejCxR
q05P1SZJR+a1cJfTqNKE5O/YQKc7rmb7bOSAeJOg0a05hZ634YUT6aq6y6UcY6zI
0ecYHTd2fBMZc6e31HYsuwL9usCteCH5eRffRxfvOr3yniFPqJEoR9piG7aB8HhN
xsY1sLd93ZhAlXu6Rm0l7XfX5OBGo/6sK+8ZGNG/Fs6voVUDKIS2bAGXnWDBVmG2
Pp4ph4MsrxZchGdC9PjNFUKJeiSpPR2SdWobodTavCl9DoqezE24jidqexT+q7Wz
UgzgX9I0SRQx5jO8A4oyTUcmHsGXMVa7kIiv+zvXw5fiIt0HaXL1c6VXC9W+0OSX
hgjjnHswh/wv/Fu0Y5SR5cOceR7OBLQkIajOWUhJhvGHsfd+h/KwIsmfgmSeUdrF
EoiapKWFn0nF1+zK+t42Q9zEBcOa5QUHPO4WNJT621ipIvGBynNdWU0j6JnOj9Fw
lysiZkd7614DB0Y1LwOHpfE6X7ud9tcp1QF0fTzutSa1pIOx1YrZ7fOPriqe1HXK
+T3tfcMdSwdkDnYmTFO4jp3iqQbmKGe/iK1Yfe7G/q4PbR7/hXvvLGLqZ4m/2a2k
CD9TPNNBQrxqVCvZ1TN+t8GIzAXYjALFe37zWtvy9mWJ47YtQXPsvLXE1aKyf+Sy
nUfUvn8ESZgzsBrStBI5FiiMzUSFrlYC0DxmdvSgWW2aw6zLdcmce2jydg+VtGLR
SgwoEGKrv9eH0Kk21oQqilSHSSAIAfY5YpJ2E9/qAG9lpUVYWjfYqiw171C10sBG
TX2WrE8sAD6NjvL1PWSiSqVMbfb/FlbZfgiVg2vSBPld7klciJ1QrmsZ8nHPMkM+
VE7o4bmTtKH6SlYBMhsiJ805D62F0USakEicw3/7C710/KspU5JjlDYQQKC65bUv
OQA1/WCpOSMax9XV0uOS9pqZbppdDvHi0zA1Pr5LaaoelnWP5moE79E0XlGD33Ep
92RXLrNDJBkCPAjpQHcxHmTnaM5vI2/7T7ihIi1Yc7pgoJQuRq0ZO4BoaygnsT7F
q3MlTFCXDfUa+u7LHENnXViFIVT2dc8KdMaCgWXN06JO2e2NoroXlOVHhXvYe2wk
DsmFgPvxgErzql/SR4cds1rcv/ljKedlxe9x25+ReqXRJWIqH4qOwfAt/FzXlSjp
gBbNYWyhKDiGJWQUblkttlqd6mGI2Argl2h93pbf0WcWGVeuZNsQ8wRw5s+lfILl
GWPf+kd6cIfSAQ4U/Und8mtowhw/XXyevnwkGBjFZ9lkLe4NqwiLKRpy7659w4n4
UsY+Flz5REEPtqY/ZZmTq79Mk+i47DHwXN/hPOGceSamJRF1WYEM1ctiHc3lHE4v
E8oEEUcQ6Qa7jfwssTjqjWGcNDgnx3b8WAhGosKu7eDL88Y/iOZejU+r6h0KJdkn
bnoQ+lboRUavbowU1iEKbmZu3Bt3eMZ5kQiP32iIs0HNfezwiGx1dhXjk7Ea7EQr
7j/yqKhJRP1DS430tAZbnJq5JmNiOhjvGgEIKQT5HfG7hW7nmgPeh39WcnD8WoGr
Xx2EN4VAFtMsmRBPqbUTEsjZ/AhvDIa4tT4ROzpsQlzZyLVmDMJArpLPPZwKnlCY
92kzRwc5n3Kun/a5ubDd+IThGuAldZqqded7i9Q0jVRiT+SyHxdo3f1pD8W5X1tF
8oVMdJYv9uapCjN5GhujZfw5z5stiOI6vxFGZVi4F3mj8JgAK5atc6QJXz6oTD5v
m7h1tOzxs4JE4dKZxiZFaNzpYoH5eUjoGMOE+mdlfc/iHCOWCRV36pz+KWDk+hwk
t3FWNs9PINKfXiFEuD3uIpAH5cI8dWPBwvAiRClBsZmWg5XgD4Nc8356yM6584JY
QPcKDTei6/kmKoLHH40+AODqMg20eT/lHCiKJBx5ItMVgK9wDSYm3EpY+oJyXyO6
4FyapFp8Sz5ZmdrGQSMtZKinL4jihIbjwQr7H3UiE8XzfcN/R5jcisOKtI8Mzmvi
6g06i9B2tfqoaa3mer6rgxsDADiNhN8mBNBj9iJSlLme/kckkc2v/43aBygVvMtU
kdWopZcnXS9mblhJEl6GvSAO2ovflP7tefeApyusJw+cuuGJ0mh9r9m0uaLTtzWd
/UBgdraFZnYW0Rj4GHxMOYeeh/vSRUQwTrGaBnd9fA20CLEgazowS6J6VHAC5Mok
JpM83OYymHdc+hhWnJVDJZ0tPMX7KIg/ogleoyj8plPgFfLZvcevNs/uKB29dWg9
4Y+0QL5BxagRd004LoNWTPE2v7X8G26P1bQDA6VlxPgrciwCjaUGwzD/mvkmfo28
vDDXpxqeT+oTVqpVOVbXzn/CbwXRK+1fdLT4yq6SGfkP31X3rbkltUoiku5QaIV/
oJXAwb/lGTIBtlxOLTh346h9XX3H+Pnon9glWtYSRqF+ApM0YmohtwjTlNfjITwY
G00udf5Z1IDvv3GEIiRUrilM7CCmmVx4B/qINzrNC5UnqC7GlA0nAQdTiojbEZfr
5cWhrX/C58+NHsvjwcyr/uea/vYFIEZV6TvwBhhxXCr/3V4F/+gkPe4UdFidajak
AEHBrQ9kOf8RjKaCcPdDfUg+9hyJbz+J8+VxR5Sd0v6MYnmNd3ppss5bYhKaiE9s
WYGPC9vbiHKJpi8Mcv+91zeLiBuNosz1zD6ynXMxVZ3IrWKS6VVoPffSBxgNFsrr
53oZeVVmgkqkHdMI6HImfELs8fW1A/lJaYJjeNGLn7qZYnwhS/ojMCNOZf8IVfmg
iTyqAuPaP4MBTLzqkjxe36d6Cuekkp3cWTVUbucHdDZNLTHxZR4rTuygDzE+ZN90
lPit9sHgNthwCohR7LgyQ+LVOimt8oAcruckrh0PiKFXkDzeNTKgYI63kCA7klbL
fmD0GXZ+qAOaNP+OokmwWf6MCLci38tuTyzx91H0mHyDbm9LNRnC2jzA2CkLnIfH
jYooo98yJS2Vx/k8UXEVemkYtsgE/ahW1oAh6VXxWv682EFGnvQLBeGKbm+UsUSE
ZI8ARA4I2wNm7e7ZL2H4FJ0F7Oef2jLVBfF2JuXjdIUj6gNO1PRsK995VHSCia0E
854T7BD3Js+Q6VrQKnKtH7URn3DDtDp+YtF2bCc/BSn96WzqwsDMbj9QcGUv1oqq
wtx+E6obwp/in5kPZLyFgbDF4Gef6ZjnCDvebr5aPDAxmyCmMWqqW0tVVlvfeMOX
a40le2McjIiBq5FMSrmoVAIbWR685v/1552q+Wd5bblUcDnCZzyJupRVCXXLB9g2
v8HbxxyRk737VjMsOgAMBxrn9ohVsn6OpfiGzU5whue+FX0BsoDEipGYDFJxRW6x
OiVIc6JeLQLUkMUgQypxPEFfBufaIjfS/FyLw4UB87E7JswxuYL/B/YycQKnPUPv
pR569n3XNngho7KDQQLfWTGXJQn97ze/ksADkNc3uXhMGh1RDVCZKWWHxmGtVrgS
Z6BG9RtldBdYYKjDZIgqgPXhXqHikL4m4TnmXMsz4oDOuK6WjM8fbg9kMG5JdVvP
E11iUkLP0ZrxkrTCSruE/74gGMNnaUMQ2uk16jL8mOCeGa943tPtQc8tJNxlG/vE
Lr52RX4e6vMezFQ5/BqWXbaNLwe1qPq916kiIu/ZP29cWp9BHkITCD2voViddKrB
dV3UjfaIPbdTjFr7N21zeVWwztzTy1fZHCBbrONsOUn91pxQ7OmdgMwVFCx46QKA
2yI3qRKf4I+EosHvhkCpE5lbaTT7yxY0yFu75+ptuSu/5LZ29+qDNi9N/FzqW77P
buLx4K8MglVLMXc7xDV/fbOJSiVVSruxrg90BXUtowIjdO7Ri20vR889/ISXeE0i
nE4tI06VsazHHkyIBQG3+BhZ+ZKUm4k3Q40ScvOmkj+VKQ8FtMIBZePVAJFJ7TqI
6atYM4/eLgL1BZVI+ZPtiszvf+S42UA9dC5mSElER/3aq+CDFsSzp1hZt3f0/GYR
qbBUKrB9ZRSvZsA+wV5s56bahvJkJKab12RXe4g7tjoynG5z20zUFw1GDrOgX4Aw
ZiJI77awiU/Qwij6y9sdbjWTShsdjXuNOH54WEnhZickUzrF8l9l2B+3BdC6tyAj
f6l+ALttdRle0zDqfv0iN79T9d80x0hZHcaxezMX96EIferB0HLJlHKdH5oDqVKX
NEDidSiYgLUFOS0S+qeo/LNagsMKt5tIdmYepg4kkyE2mN2i85MYsspPJKE1BrIJ
dR+hgDsOdXvmgEWGSftxRR37tmL60YbtMYfE65IFQtW834wxwNgNbSvfHaNfKWIo
xZyjrT2jHofQZc2kgobAx3T9kNvqEebFJ2gXa8lXB3zyj/J+O1Exsz+U8Oq2u5HW
jGrzsRog94W9Z5cGyCoDW/7fH1oPmCwjc2PMFqp89d2P8VGhlxgPXW8nXFtrEjPJ
njhuPe7JHMwIqhyaYAh3kq9O4SwEoC/PBCEdWkfMLyteWe01i1z0O7/GFTHdR2Bc
TmUCkEo1tyiKvUpb4PRyf785X8tao0lOYzZlKCW7S6OPpJUNROlQ//6rQIUfu3Ds
mK1Jjzy6QvNhVBweqKHaKzXdOyExJzejRkm83ItyQ1SHqlJ02o0PSOqYnTLxvKhs
vYguaB2iUTnq+UupiyjGt5Ow0eZI6kbvjRFDV+uJ/J7Je78mvdnWxcF0S/35KPSM
//ek+6LzxDpzt+eZyu6gOo8rN2Arbez0R4Hxu5tcDQYjYbQ51o4v5bsE1PX4JxWQ
JpfBAC+GhxgItwfAXevsuonnVnusCQ89PU/9aSjromAcpAaCMpLV2LYZ6uDvIZ0p
OpE7PSTsgrKdQjYsKGkyIfjs2bwKRvwVsJs1DNZ6XpxXZuQ58XgN3fMqenyYxemZ
NbmfNQ4xbL/hIDfAXpFiyG6w8M3aoVlhbFXn/7Q7+COxOe8P4tzVtM7as5Xk5UfP
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7152 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/T97rZhQva68T7JOm4bkq25
b4BW57ADAHEm2yg/Vzsfl7TOuMe4xzV7rdHsSWg325uL7cBP2fSPzF2gWAp4T7wq
bbPFVuz2tGJOVgHyu10KCAeTzHBIgZDVseiShxOC1NHe1G4CYRrwsHXJM7dvm/2x
i5lkkO130ePVBAFUBj75eBf/oK2I6yAUOylvmbxcQY6ux7JDhgQ6jQfQibkw5puf
BGRll4V8fiw4AWLLuGqIH6A13gu7+gAMK1EjUmYfCx0YX5K794rwKM3C8+q+a1/Q
dmC4JCNzugse1MVnEEmi5T/vLoF1MFMA2XMuTHYR0OhbW5xJEz2T32oHLR9VCrKL
UlZCXSDRKjVYniIlanoPX9UCHR+Esh8zAqKwyI168f3gwvj2C3+/ZCY3RYDgEycl
bg7sSCMZHvPydSENnaM9H2JKfEFtUXJEEFmkKOg1fF5RvHdauxce+lMwPYn1JkyN
jIrGLb+/4HbvgVOHLjJ/qxY86Xdgv7pRNt1EVO0pjdfyjEpvpqXchfS/zR+ksMLK
S4Wv1Bw+tvgEKmAIH6KWyIpr2MvvcE0nq7spnMBPP4BkC2NmTu6G4MBWhM+2mvgZ
udOkfnyV2akshU6DrY5OJNaH7nFhr+lnp5ZF6YjSfscFY5rm6Yvt9X7lPI1MtYKi
7pCURoyLQkxBKaqqYJO2uKl4U10iMotjsNOVs9I5qpTHCSaxJbTx/OPM1P7C4sG+
1qD11c4GFBjaAtrA8KBKm6AjPZywbG2sCh+kSpN/iugFcV/awsNh605lnk3emgBB
hYrZLBSzJjjV6HHaUL2p3TGQohRTorR4D9pTP7qgCk/ERjGWbFZ9vrfwtJP63p+s
3AOwbJllR394T54U7xDJGJo6DNuwwPTncMMZMLv30s0O5DT4yktnIvWSDz/HQrpJ
afxWG7c/L8C4QnHdKNq0EPlehLg47g/7I66S6ct1+wiQCsyNkAUEZ2EUf4xjR4Nz
u7cZsgAcQ/l/V22mNh7CBbIoXNa355wYTeXz7/ZX6Wo8J1s+3G9nDnlnnJ45bg5w
qDysE8sny32DXZIDbCFi1/mKT5zdJbvdoBo2qS00XjlXTWDOFsPa6zeP2/hqLg7e
T7PbNOsVsHMdmgO2nOnFX4jAytfgtxU6HdEcAebSF/bst9IjFRPCmDeyoOL4dkdC
MNscKEhH0FduepwtYC8l47Jc+R3ljm+/ZN/mblpmRM9t0jz2HYQGEdHpH8DjUHJp
/I8ZpNy1KGqgBrhZeCkuTEh8PjCtcNYPHggJu8jPOL2rmoAdhabZpc35URTyMkl2
fN8WNxOZY0fPiPREaRngudZZqYR1C0k/6V8WGD/6aDKLPM8a+MKpGSXq9iBLRBQr
auYX9hMcCifOlpQFhRPQMNxxG7DSnEIkXpiTqG67cAfm2PFf8nRaypQH7LN/VhKm
nuYacjbaEWnM/sQX//yu9IXsStU3ATvUL8s0h2Q+9/RLgFNwnhzsd5FmkeNaP3Gs
VADED03ytxCNlTMrFSGgsfZwHJ1SycU9HDCrMrdVh3fbF99TZEkJhEPuICbp17JZ
UXgJ7qpKuqGyx3451zA7SLwVKLFQN1Y2frrmLDO/fgL6hcMwrzsMrnkBKyrLLgoY
BIgi4rX+X4fHbHcDtr0F9gkfW7UYrrpGeXQI4ANxW0xqf6yxwBQ8OLpNQd/WMXCG
5HUUAN+QIbUPp2yCmWMjG6G3LDUsPgj4j0DtYas3jVsPBbrsuyMC64XEj6rFehy6
l9yqmxvU8DhFNhhmax1QjlUgtsg1EPW4EQMyzuYj+cLg+BnPdzOYqtD1r/1k9jpN
TMDP1/Io4mFCe+sBMh6P/1c20cVvJ/AQlgl2Ny+KvXr1vZGX8kHqfLvokcqfi3c9
+M9Rx25KEnpZit0elzOuSGghjVoZb7lUnuEnXfrarLEnqHYfPv558fBueZXpIjG9
O18sYrNUA+UzWxQxtA2S0t9ay75d+JL+6GjWWl4Cva+13jEZspabKeXl/E/i+BcX
IWWfec9jws02BlHEcfFzajNB/+Bbdy5ZElXa8bHpfRrUEFdERhoz8FEv5EIaLohb
CKQgFl6JWn6O+fRZJMk+16yG4mJsioNfZGrNEAR4OQadL+AbgGjOPZ4NoDmNb1pY
5iLw31JsE4FF2drD1WV1MO9CJeg+iBs2ni/RL6EkNYy2nJ3SiXY2uBKa1kiT0b8z
Km0LIKui1FA9unAkYx3cFj+0Bk3gRmCHbv7j7i7rBkzSbgd5Q8uYlR2KJL5NYjz7
5WVsPMhYQ9W639tbzL68RPb/OtIZNue/xbXsPucwqdhUvdg7GXatH4egB9gJnuJG
LudWm0RpfMQZpFFX71zsfmAxHL7HOxc3108W+9yIFNA0PLICcBS1VPfxiwMw12jn
Kje2RNnoPpR7dPPITtw3r14tO/7eggWPqMZEQUVoxII415RbZ70FXMV/KvPdCBoi
YnxmkQN8tDmThMk1B7q9Vr1/RFeRMnAid8kUWmaWnFcyaR2CE/yQyUhkLXP7wC8p
QkrCsqaQyFRVDiCMiAsHU9gi1Wg9coRbk0b2h4LfCTEr5yQEWJZYC1bwI263ZBe/
STMJt/T6lH0+5DUOwYsOtBwwVZqrERSThzhjnIuQ6QCf1VsBY8kFva1REwkphrmN
/9p0DxskS01piRxcW+1IGluVSxdcUKwfCMax7KocoE2JkUMQgdAU4+h8iZqyJwVo
6rEdijWp8nlLUjJogIcUrWIIBO7ioWJ0SDUwQ2gjf0OcJMsG8bAv1AwoeIb72IJ1
mydT+mGwV888LVZqnMTbsNBCj2Hh1Gb958Rb1Mcsk3kj6GlceLrWBsYGGL5rtBpU
8E0UWo/la4h2xBm8mkzhGduFHlCHOneGdwHDQmRI8zgKc2kzyKh8o4ikvihKiT/M
jRBCrLnmx6i6/S5MCqaU/aXMh+Om9+GOH72f/cQBIdhmuTWXYbqFJev1dtFXR9en
iemQ1zePoZgi2uFObtDUG28raNZ3mDiCsuhsnY1xfqN+1tEn6McPgzQxfZs938vv
IHCLAgw94hIL2tP5SdfhYeEKzutuSGDhjd8lNqr36aIsUGpIZziFSlZQ/0hy886Q
A58L/HJCgw4F0AFR0lgtEFYdj20XkkvOdgRlm8qhoSmlZE8b5R2aQWp19AEODlGB
nWFhNkrZzdBq3T++iE3SoVTOq6otFWZSfosRTHvpIfwz60Z2rD9WPy4MRWhOVvpm
h3dd/Vs2/92RPGDVn1xJ+5KDrR5oIBhWKTZZumOEuDIMxAhon8R1VzeRHu6/jPqj
7gPMTOf7wG9f2Uz39vuLl8N9MpPmHIRboRSovAgBj3fbzvsF/pnGAAG9uiztubsG
5+gaVSaahlQ5ByK/U5+d8rZWWjeUtV3iR673CXOSL8vCgEF0BzoHWQLnCWktCbh1
07nAZTm8PTLmNjhA8MiAx69bcQe+S4ro1mIruoLvBbsilBW2yRfqKxwCutA0ix8J
ASgGEGQBbi7dIeapUHpDavG2VoUSD7TZBjg67wMwIwquFBZwzwHQQA0VqzaPYnUd
yHv2li4j4NwrJEHkYPbRC2WPcnUx7XaXINgvWIKIkcldeDdKPRq7qz81PWncez6h
MbQ3aEZ7FuWWqs4+LK2yDESg6g5olOe+E/YHUMvj0yonQivis+53qk3e0Ed2x5cc
mLw4Mb2f+15NXXxa76th482+B/RFYdDIMotPezgP5Jv2VLC0uD5BJ/PQFPfMeAJM
IVnYPTLokTqmYU1z8xeEWiVSCgZrwfqVAn6rAbFHRvtuiB252mD9Zg7+FBEHMorq
JWVNDQ/av/S1MXP5Y4I/GgUFWhUSc2wI4l3pNNwZYwRLyiwRrZmZJkXhHv9NeiQq
gX4JpKNaAsP7qqK7CexEXz2CzybFv/t6NNFz712F2y8MemgaMASX5LOWQXlaF/ZP
KRc9A9eBExBQfu97Ik2ef/f50hlllNHLvu9UWusNK7uyFxj/2MKXctUfmhQ/Tdw9
wvNJfd2ZjNKsjGet8fApXd4JqG2ZxaQv/0j+E0azbxsjZWNeJwA5EqRYvidm49N5
fGQ0ZiHDaJUMLHPRPpj6tE4kuUswDOjebeCFFu/5IDZTCM60jiuLOJLXByUWGoZg
VuMqtfQxgHOLwv3r7L/LSwyenGpoP1naOfTuYpi5Xz3OnUaBjJU/VhkL51EbVPaP
xRtqu2cEEEX1+arrSh7f6t7x1W6dW7R8BnXFKFx/Kb+2uwHsCZk9g3ajksVtKTV1
/FUpdWNR2cPYFvjA/qp2BGaOH5vlelw9BzgGdgAhylRE9RXzci2HfPnPAZbWcpqu
RUUWfwQuHY07PPbHYx6Y5H9M56oU64TRw+OQ2FmwZ9hGqNX50TibjqGH2OCfUi1L
5rupToCjp5cUdTU/hmL6pYgNBACECy3Db/10J9d/H2VT2Mijl8LoChcwT4fJKjtr
/gy+x9AurAm3MINDRqFyRutnsLYr1e8sKdE6qDICc45wL/umB2ERthQ3XvSwhstf
50OKVPbVG9y9suOpFk7qGzxW1ItFQcDB+PxAncSfu5E5phcmJzG5Pn3BxaML/Bn1
KgSEAn0qSz4FDWahqEQkDlXMa/hQMYLI15898SuxkjnpMDvJ79ndsUesGscA4xG+
DixnM8c2B9JHGBODITQybMtBTMeUu0qq1ZzdL03N1qrC0in3yeHVvFdCjzXYR9Jc
SSPi67ICOirYBmg42B+4pjeDZ+CPbqpqgqKoH+Y4VLwswMJr+OIrOK6qxJzMwVtw
asCuj3dIspN1mqU+dbqLl3fCzEVKmXd34bWcULqSXp0VUUKKcgOPOOoKmZkMkdzQ
cSM3UGkR9nxqBC8o3V68BnyFF7OFoC8W6ftBYlmFThyq/41YnntxUQGNQScPAG8j
G8Q3LygzkpL7w2UT3E2Whahklk7K5phdeoF5k2RBF48ZQZWDqLKaam4x7VAVog85
RVs6ZD2HMhXQiaqqUP2Hb9L9BEth0XNENdCFzBOlnOAu9aD8NfMIERShcWbv73Pd
8DryeuhHPNaqyoquAYVae5mIzPXOGsY7G8vHbIoXfRyZd10r6pFJLEORm2G+EZjI
5YHFR/k2F3mYifs20cLOz0Aa3aZgLKOT2EweVn5JH9gqs8+T3v96v1OBOhrmCu9r
SkhtlPMByoekWbbZP11GL6b5U76C+Z4Vjv0BnItV9fDHb8sNGjhWWO5rQEJ1g7g+
fta78BNMa5RBFZJpBv3cwFFYVu6tJ4DfLeAzN78CYCelfgAzdU0u+EAFnvQIyIme
EbZPJ609zwPWybF/sdjtRBCtj3omPjjQBSHYDOPReTg38dtUCeVhj5O6B3wZ5PAz
xMS3rlxB0gAUbxDFe+GsPgxfn7jfzygZZf7otGQjluRfHBPZCzkehkSRbUxnVCXz
AihBYMMnW2oKtbc8X4IcVcBoNvFbqDUSLpIH/l0dpeviTo32K9AAG/9KSnY35BBI
qmJOY79wWSIRfb2luNjaVPtlW0WnR3B311dfS5zaqJaIIY5Cd0nMvR6Im6TkxK/d
D+hZpBtNatdRQyVF9pzNhM8CybYUGB996vCzZn5tOzK8OhyztqB1aTDzrwbI7oRG
HRlxgAvcWQzQUKek6d3gXMdEc2WmvNAxVKuT4xZq1cG2AHdW3zgcysh9ZhWH2IpC
+DRZZYwOYu0aF9yutYrWFXOcFbwfVXWIvMljlxtKAPJpow7B4xei//6SN2aR/uQJ
A7vcAaaVvn7mr3ZRPb5aeFIy0xqKWroPE4kFDN3fY0GAg3vRKPwvPZnCBdnTt5Kw
HrHXrvNRb+WHNCXqIEHun5ibbf+pSk1XewPPTQ3g/O0chdQMWeqSShAssi7CmspA
IOBGwc2fp06SRzK718t5mzchLoVmf1uL+umHhmebK4vVtxLFB+uRvo9Vih3fUeMd
m4IgJhq+g6/3TqNRFoHQbIBGvugjFdLHAaiRPLpcv/GdlyzW4mbKf9UXDpTr+5Tx
vSMihRx3L+SYSla31nBKJv2dd2PxV5QVGkGJb/wqiRbYbkCKIXWRCHABadzokeMD
ROgAUgLQMFrMHRwdVefkRlAgKLV435g5qqdY0hHlWs961rZA1JRzvOwt9XxwN4tj
YDXwh/kv+wl4L6S7s+LADv9yoPohK8KY5dJucG2r4EIxUZgxfs5oNM/qo2Eq7E9X
KJ9V+lgfNn2a/621QK1IVCov33VQsXD9PgZ33lZRszb+uU5vT/RetBNMqYz9fNT9
d0HKYOBNZl+KW//BNSgDDK/AzH5FqAOK57Z//2WjLk7KqPxbPROTF0Hki7CFtCre
4YiTbnoVVJxCph54bv5Am+zLZ0F2aoJ4e/rJvIboDZHg/OJ75AIgWXW5njfAHpRH
cAIBy8btQ4PcrfDNzgt/hKO9GbKFEDMhWN3Pq0+IGBOpN6jDiiOsmugaK/lXKoVe
GzlTbYps9vdyzckz7x5dCRYsUCgxUq2zw7XIq9DjTQmrpLuNel7N3V8o8R82eEi8
ODM0dN+hYagJd4XgH6IF6LgJur5k2ZNRa9E9/rxTvacs4EAwL0dHD1lJ2bqW1jTl
IjM9AfGdWPoG3IqYH2NiKOZZbMfHIFT6fkC62G7D8ydaFNqypRvC34cztKinlCsZ
Rg9ZqR7kLhPNxWU6ywHN3TW2QX8ACEY9r/fkpBPLsV+Lu3o2aSOVM6qyRmUjCjEg
pLRcSZJJe/zES5NE8DfVHu9oG9mwXlULZhqrie5mROHL7uON8TcoyMtynS9X+wlR
ZfBRLphvim9oIVUW7PqwucnV2863VK7UhPS08waT/XwHC8w9Lqhr/SJSpoD2ctxO
qFYiDqflcHd/vQmhxt/gez7CvhVEuI4bDYkfp64xq8gr2IBF5iRoVSnGAUKGDOB6
3eyO+5VAdM8PY1phM4HBn1KzCOlVd0ebk4RVwjtUK/gcCe0Znci1JE18lycxUgr7
RJ3Vo5BrUp07xYTqWggYbaFZC3oAdyLaoqvpaZ3XEi6A9oLrLdETb5ThIPG2gXad
CzaqQlJ3xydzN9B9/IroP2PGLFmdUxuXc4r6B/BwHKWJ97/oB/qWC25P5fxp7van
nKSRf5yW57gLXjfhlOBUnDckL9rMYvtvZFQIzqj5BoOk8JkT5F+h1nyl3HYHuFL8
Qgr7R6tPBQxfqCKm1q9R7PwTM4/1stvaXvj3mziawO98MlVnFDCHl74l0vXIiNQQ
//I2kwoyAtURqnp6E+VgObUhyEqrTE0ugxftJq+WMxFxVHAAEpDFWlZ9egEpUcFA
OLvtMInmRRw9k9YaWcerAJclzd9Ap4bX3EOdEGceAXw/hMTSQLW36z0q8zHGqYHV
Zo7uO2Z66RyFH9/BwmXFAaQtF7oKfZdwUv0s86+Nb0hJ6ximHi2l5MFR+G2sd0Nc
DCovAmSOeJxxDZtrCpv0cQ7YbhFTTOM/nbEee75dZ/MqVvwkoBRbi0j8scXK2ZVs
K6BX8oKpjijvEddbRms71wERnnUc4dBbZ4r/NWaDDwH1fNq2o744aOGeuaJxCy1L
3oNYSeMoTdN3VPQRqe/j84SubmyUOMxQKr97lcZuzLQe7PITdeaalpfAXnk67hT2
sAAkj1Qew6p3ERKDERJuUrG9NAb/ZmPrr3J2+LpOfEJgYRmHiU2MOqD65+cpRX2E
S3Z7YxHB1ZE1uaxZ3im3O0npYuT/J05HHOVCD1YfonSS7Dbr2/UlTDIMJY3zBb2e
JZSpjoQVMG4s/5BAOE7IOMSfAj7zVBuckyuzN1SpWvPwZlE9wa29uDz6LFC9odto
UGqR1PlexCPkJ66F06imdHFOnlHoqV7JJcfNqIKBvVIQeMIfkkc0pfIPGdZxENIe
tIyvTv2r4e4LQtWjLMc7LKuuTWLNIi3N7lVLWANVC1vxX+BNXZKVTj/wWa+y4OBL
W52VYU1Fnm+4EaTDuz4C34mbJhercKlLzgRXoMezOmfOpoh1rM5C9stjT2Y1Rkwj
Cvx/xVo/omfBmasUp6FAOop2dYntD6Jkrnmej5odT+HN4o0Eu9CLavrf2JuWvsLF
CcaKH2f2WuIwEAXvdB0A6R3tGwc4I311rqbYnbRc7VzFoyHMtMU0JKKyN14MqG/K
g7QS5kGZ/ukwa6WpGuZBv6COv5ot7tgvuoVRQvSnoHERms/QM2UFtJ40ntM53UOP
LyOo3bT/CSltFclV2gmOTiEjbjZNXhjp7mbe4KwAF44eVhNKF0cKwLgg+dJ24Qsu
3YCU2tLAMsOMJq1bAbjxmSRW0o5+xzEy7xlgsYhc2wMzzQFaCRnwvabigKLSEcPp
YI2oKttDX+3AWPm/BIol25o0siZJJPCkSfPk4UO7ho4bNrZxT0HAMdqzbx/pjBoW
x1mx4ojxspgYJccbzEkxvg8I/bV0ouvZhHmGxHPQbki2CXZWjVp1rcqn0+E7kOj1
QATEA6T7DeYYr6NHLF8q0uPv0g9KBl4L0+uc050bCYCJyX+uz0qfTxB09nf0sX8R
hIqpCht9l2IcZ4vpKqVBHXwBZXav+JlayPwvYHYCm3APsUtjSLlWqcxPN5Wl5lQJ
GFl49lY6ExP1jbcXMyWK+bTZb5HOXiwos9Wc45g70KLlq0+6bM6zL96tzHj2cwmZ
10DcAlrp63HRD8GCoaTSyj50nTNSKvTY4iJyUP3QOFrcykGlLe6jH3pI09kvfTDm
yx+QIvSLX27/r94+uoW427UcNwJF57oOV3gS7RKDsTrrpUTBCohXUSaCxk6Dg96v
FtgwT3XPwVoupyM+pt8lsF6mnh6RCIZaHaKJC/MF26xngw9WiI8Y6RGNp+1p8j72
Kj8qE+TM7EsUWUjxIt2m+zhnRieGf7LwAne+Gqy7W6GFo25OssKMfugA9yd905+E
I5uvh47SQb1w/BUh3OPn4GEZyyfjJCGV7hnRk1W48RZkYewBOmv7BR+AhWvXE6XG
YTLq1fiYgAXhhwWg8FRyVqPHJLIB1LuPzqWYZXh91vkGzmDWSa5MhfgDOKezTikD
ZOTmT+t/Ub/ph9k3PoNwyhxr8UtlQQIPk2aaLMQ/D/yyaWvuc/CO2VseBAyc6okY
aUpVoVd86Us9MPUXfosg26GHNAzx+RP+NXrdfSjoAMIlfndemEFo48JNYCZAVXn5
626gxP/ncOxzts7QTD3z/kGDOy6lNjNNyQN1hn7QS46o02/11C+DMLO3eg/6ksg3
hn9/r9hkfILUNGxBvyjf0paYVWqXdHPmOlGDR8aIgElUAQ59gx6ux7dbu9GlfZwR
EuysjjFJsWYOVd1H6GzekuVIdVix+BDBPDMOQ1VaQZZRULDiXvDIrWWCXxpgMcrn
mvy2R9VAXs7lAKM3sP5tOBjGod70WRQqNILAci0pNOiz3w4xx+ZxdHlv5y6pn9gv
zKXPah6Cp7RMsrNMjXBhWaPcH0cKQYIuEVD60DbCMdzRA+VBabeSnw/tZl7Py2//
>>>>>>> main
`protect end_protected