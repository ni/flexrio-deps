`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24224 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
FTGcP7VlpSOhasofAJvqcNBuJBWRM+O7ECOH01Xn0Tm+WrZGJkPWXsHBcpkyFYV7
gbD/F7tMdMevbNbdyoRencx0x7ZK/VLDBJLYH9E+VlQE3S4YzoOrwqGsO2KbbL9K
odPmJS9Ykf7HYVBSDbUsF2oBGgO/6/sm84w363fUf5OuOJ1FpQOd29tBJ6aGw6wl
Ep/ek5Ov8yUWXbQ1i7A05xa2ib2IUikRNoBdTmihtkikJGco+DQ/e8nSgrYxvO5x
SLoc8vD36mKk23aaYGgY+8odem0lUwXoTR/LB2Bc7lC3j8EBJIaVW8OnNtjd4J6t
E26DU5ipktPdvC/VdQZjunXcDUVfAPiXZ6lKe5XFHDL8cXkVvfirOPRQQqzZ1PcL
M5ER7drCEUlJJl+lR8JuoIgjSXVU6OI8IXTTTjEydtuEALPpSb76fkg+sZ77s9JT
DkpJWD5euzy49DP/Qiu1B46LFTsZSiMQk6nXpQD2uu0iTyW4b66wzhjvwjY2XpfN
q3YQpvXXAccbLSTNJZt9Nie5PUQX6KBTuKILksR5afa2NcObADSCzrzPUoWJGnc9
zpMgP4tqovVKFiI2WmQMXgmNVHUfpVrH9wGU69kBHwOQUyUMRJawtzwX1HRAx7Ox
Vt+SMXELRIhpGiOGLL0bEIztnESdfpBaa6USgrAHIzJTuizx8FTUg40pkgukHFO3
R7ezUBVck9pWSQToZ1zvqjIdu/XhzcKBch3COvI45lQpkYHC5dLcVcv33BWQAgcI
zBbrqgATQ5KDp18p01RB18xDunejoG3VAwJY0ZWLYGxZgdyHVxXF/qz07I648EqB
biuCpqUT2RBPpqqKnac+6jQVAJjeSPPkyvk3zw82jJlMVKZ9nYhScoJ+bfPtz5xJ
G+yJUIomrCE1IABq5IEdl6LpOGNddXanRPtgKHntrHy9yZwfnyvCK4vdl9Biyhi4
tKhtKvh0wFFe84QGFPsFBHk9VLa79KixPDOlp6C8Oc7X/A+PU3rWEPPDQhccJ+qk
vSuESz8yFJs6MQXn8qoysKdvclE4vpGrlgwSeSg/zTUHUBdSShlOmiKeiNyxe8Ba
dgyn2FLOjVNVJa/Wbwfuv3do5gaq8ifIX3mgIPCBRZVhftV0Tf/LXppBfn3cDad0
yRfEE5KGcjy3bArq30+bCiwKph6+bGntCR395LVthjX8C4DJ7n53TKIhLQiFJi7d
296uWrELXiJJjLLuXTi3OKf8y/ahyo4DueX1Q9hq2HGmu2ipH9Q8jvxASTbKknSv
wVQ9iNQ310ZcL4nJA3Mng3xP32IriYgAf2DPN9nR4U0tE0NOC7yPaJVFFRRgWFzM
vs2kR0C5Xfp0cnrx3iZ2o0p7pvk8tnI23t6hJ+irXvDvN4U8QQdWUrW9fIHgCUsn
9LgMG7jut8OiMOk/zKsCZRX9GVpxh3U3cGhYX99CucPUrYj8HReiZxUprjaWj5Gm
XgZW9RY1oEDUN5mUf1s1WWG9M4zgJptFXdEIbJ+5pZR/6EJPnoioCYBKTp5PIc6d
+ll2lu3P/cBBRXIjxmqDRGURhO6AgQ0bu12BE06JGz16UMtjVtEpWDUdlLOrAQLn
6wL1CIuW111naUVXF5SBNV4qL9IucixqhqTfjxzRRuntdgNPvDe0D4Loc0Oc34xl
ONWUNtGwKPKMGTAzQJBF7S2+NXPp/ABU5OvuXfwVR3xQ3FT7EpkxGN3g3RmUTb8S
KYgleFurQ5elwLWv7yBZufggg166iQ9U5oOMZ30dd2AzUu6kluZ7nAjQerrw9ppl
jbhPqiuUTuATqPKuBfsLgxf7sFJ7hFkcqHnJypp0cIIEXtL7BOTAmHyruAjMv7ww
2ReLk5VsiR2nzb7ODc8LaUNOnOiCHXJb7mEW0rMkgPA9nkOJ3YdP7qH3t2OLkrMi
AakIcrbPDSPg3Zm84oNF6CC8Vi1SjCjZPPu6SVX+QzRiY8XWozNWaaCetFUrR/sx
8p+iI0dRGECYEraemG5l2pTNGUSvI5uWCnmvANxB2IgL1ux73/al/Y5pNeN0HsS5
uT/E7VbAgAozIU1F5y/J2Po2RUOCzptou+EZgqKjcpBjxnIbB7zMFgpuWEok9TA/
duHRxGRhZDrOoqEcUzF2pdchJahoDeTT0EtNEtqdcLLHwE9xzGZCkpQM9BvZiDqU
VQbqMCS8EMbPj7T7FJOAEh/Rh9cemsZTemQQwiik7CPCv3PcU+xEX7z7+iQxlGml
OWXgI9gymaHQxyc3AjVIc6Nf7Jhx3TyxxyBh6tHccDB9bMo61KoZoff7U+8/O2l3
jHcJXrCJdLPAADNOme4sdmZ30IxyjEAIOeF7RSbKSDsU81XHPJ2yDGiK0mOX8Jdh
c0ESoY/kogx3FCmFXDvrmBnxZGOlqwXHI/lRpaiNTGZneNUtOXfwMIcmVlhWRlD2
KlYlI6Zfh6HIsIV8d52Oa6oqE+ig3R1KYCtuBB3PqqGVA3Ecj8imT1h5Rbtiw8gX
waF8QlTeCYkBY28xf7H4d99HoGOrEDEiOQ0LUaxdfiT6bn/s4l3sSrs5J3DMkcQJ
Xu8B2gwT7P8kUMPtcqZ2b2MeYWtA/JNj8x03740O7qbY1ypbQtsaoozRlRaNRqoE
0d/58NmFdqKQWKpByNrZ9/R0kUpPowf0GAAAIvkECb/pAWwZF2d6Kq/qNhwbZGPG
Fty82Lkp1UDMpOOHCCaOwNTk6qjCR/UCco3HT1W6ME7q4Q6+K7Hb8ADoPkSl/dTG
vSNv2dYo9zJjfW/pifj/hIT9WC32WkzPR1wyRB0yp+kRKYivSOilDFMyD1anf7+x
tSgVV0LfhWbkWL91IR1jjjyRzKDQ+2p0fzIS97zavwf66j+wPEDifEHXXHcqHoN1
MBSOeFjCcq8KNd1drZ4fokGxLHLxHrQW2xoH1MOeiPZRZX8zbxcue/ZFW3wOKYln
UZYkR1/Y9p93IJpgQvQmFskLwLlFws9z+mCq+3q8YHMAyfcX4SF0k4gWlvq9ZcsC
5hjpwmLiiumOC5WueTb7MFCAJ8R87B7VjpW0HkW1Fx1ap7omtlrkDG4QQbFjpwWW
Zgje+mMhXiGaEmmMlkij0wbozFyzjoLFFiMUpZhugpFEZhi0WESvEKXKQs6ioPHB
aDfUDBqv4lwWvHWwO6Zxgb2Ln0//ExAMTti2poC3nCHchxmSVrg3HFdQeXTVVhim
kSLrSxo+N0tv9YRdPMR3FFlq0nBLn2Y9r47cwKs+Yil6MCdMb/ktQX+g40dta2Sy
2alsHHcpDJLaiKMOo8z6GtBwSFR7qCkLIDFjO+ekU5gMs0MvKJuc8H2Q8MdmYaFe
0ZfYpDAIDGOZ+JFUm92W+TiojST1IlwsdZOjV8sgx6+8BUszkhdXxLJO8jvuLgOC
XnzisZCzyKRI6BXr3UZkLXtpGqhjai/dN1A4DxmoWASBzzB8hwjHdz3MqTSwVH9o
cwTU18fsEOfvRo9q3qOMOMl5bP+JgNzM/+hgYLIM2eCDGhM2CokBsbBCGUAtDqQ4
OSZiXVBbG0y58fvgT8iM/xHiZdrM71OoI/5JldpTLSGXsVUKoeKGYeKN/KVuaqGb
Sb8kwnQKIAbQZw3D1IBKsjEoaa1nP2SHSV5gkqoDePb9rECeH2IsEzAHu1Y2p+Zv
Ba3HxbNXNFpTZS3/AcAV5EiHFypPTk0LuzWrSiAF0eBslVB+eFLuFjrUmAgHfcsd
T/vGRR/HpGPzicNWRbGIMeXyNPPe06fZg9JvMVEi+Gu4+u3168T0OzQQ96tFycd1
7SC+7cDnhCV5a1CwkL8gL7NGbN8uaWFYQi++mK2TS9cUYXADPvgj38/FaVF13TXe
413ZnxQWaWQ3h0h15Cc5mYPAIJzQWXgRT98mqKws9JBpGriSJ3qvmWdQx5cZXtRS
+WwMsVSvImtvdX4zOgJBY4QrtsFKPO8OB/hj8IHGwxFcFR6KLkQQ80HziqkbjuGX
eiX1+DDQ9ZOA3Ew25mvLDHQLx6W8D23lDKmdYCxA1LHIuUIPqIE1YWCcBpKr0YmM
Gc/EmkaqplEEBAtq8pLKInFnBXDmMjfd0JX3+1x7J7cYlu/AiIELDSPb9Kf14r1A
+YKBx9ZBw2IFTMqIwTNOK5rDiWuxegb48elWCWZxOYU/TYRv1IAdJ/kD6LxODGTJ
Q7XbuYMyPfG/CA4ROrmjDDI5/gW0KptUlg5gFBEyfnse4N/ZFdTLud8UK3bNdJvH
3n6E4B9WrZrqEiCFmgpYtpiZd3JSlABCf5OAK053KJA4OqiOfJ8kAjsd0QuT8tjK
6eKlgBNI0JCtjWSIoecJGWY8qZ7TIS/UL3OUOgjocITiLTNFGOS77k7t8BId0hIL
FaRIVhXNkfXnzdr5PsKKkr/sh98PvfU+hDyK2Vs910EsNgBe2ZhPhm/rXFPqNc5F
O4um8GryJuJ6NmNzpSC2zG53U1taykmBpKUfImCGE4Pg6n3XtghudHHWSckBRHYK
jRoA34ZI7fa1Xl1gsiDkG8x3YfoYl41nY/kz6xQXlnFfx7DL0JBmL7o4lYVNDFXD
clAGUtNDzfsL/Qj6SYLqjSjKLIgyVJPSaZ1LeisEwlCUfiMyCPw26RngpijW7tMS
3nKtoBlbRhcnwlTa9zLLB8WVMt4/t68mWRvmuD5dtFycqlwhFtgkHuL0OoZnKlpj
M07yQGjCGp61c/PajFja5BpeqlhqOtzEtFeldLhjdEw66CeC8ZJcl45ppDm3eAjl
JG9iI1LWgSjWIA8Z77HRe7qG1AwMcKFEOSOzRmSpqmv3ZDaHorS8G/jwq+fm+WXs
pXptvrAaX43yBVHUDTNOr1R+2vN/gi6eiwRhkfiky0eYb/r+1uSVoaP73YZDhkBg
KeR709cx3/B0PcYka+5/r0/1gF1HkbsESwy/qzGg8fAIydolJLwP8MAKYTX0AtTM
ehs9eT7Ne4FbSwTiu7Tz0pCs99LkRRSZaT8DYzAeLF/5vDKqs49dmysw/5Oh8aMr
bxcu2dhKXzoAXan5pjGqt5ueTIwlrOArdL35oUcBDH8tUfFISBeWIdqIK+Uk3Qs9
NmzdAzFEyDltSfJAIZBFT35xp2A3HXKrP5bMgWGm7V7C4fOzwRhHmjolBaayIu+U
+zmzI2nMi/wyjI//EGyFG+t5kZVALbClLw5VW1f8r0sqknb7NGdehobhbLqJSHH2
n27AgSRZSAfWBYfj2eSk87mujQVXPqhGpOSyEcgiVS8zrcZe2VRFvq3vrpiTEbPy
Jmu+1aXiOPC0V5WJX8HEzgBZQHHQufqa9/J6PQ32TEdZx9vAx2B/mG/WmFmv+FOR
o9VTF9Whk+DSSqUjgaBS8nOZ/jU4oItazY0by7euI73LpvA38MNuEEmTcnrrAsnt
Lwes42bIwyU/enXT8pYS1FptpK17QjrhH4g+Wv3I4guPB/XuvzGb099BE3yvCuWS
BtIdohLZlg+ZfisbkLImWjNvJ7/q/48jxZu2W1d+RUX80JZKgJ9gXneEK5+K0hoy
7qYvVRLL36CzFV1WX/Ip6Ul9B6x11HbRCEsLaDa+7y+RsksgZ7W2QZyu34rszOZ9
ACPcnVPhBCo/uKEIBpa2PV8UbVVXEunL6+y47vaXSDh+eGJimMZNH4jxHpoFtTZg
NkURDE0DBNObdz9k8++39wS6Fauv51vbOqnw0o2FEOjNM77MA69ghW5j+799wWBe
0cW8iA2pxWXZMSP88NYdyslxi2jNqVGNT67Py0TFpZRkmIuNoqnGKAaUEF6XJf/d
FDLNCts91CQcyFFci5vgmL5EPi3q/5Uht9nivzgGtnRASh2TwRaZUn3+BsMjhOBW
2y77rggDZwpwxOWMNVqgJDkgy9Lb9ZNU6M4KYrbMv98RFPg8vY+fhZM5NUyNfhb8
BO2qfNqWKnLWOWkU5qUGQL50pCvTZO+KDfxf8MEOYZGaWiWIhx/QGD3sLZtSH7u8
Ddt9nLTTyATU5RvN4nLV1Wt76oVvjMjKkBVJ4E6proM4dI5X3PEj4zwyRmH9eI1N
zGf2tLbCdBcDLNPCZjCzSCRPQxisYWunbOwA1XG01fWU8bdBHYGe53ogDioQyDJ/
pshT3rzfhjJUjr4RBIr7VM8rKoJ2warSTz0d5mdURlB0IPugZANbQTjq7P0le9fp
2HlupMkQEUoUF0UL25l8s3AIiWm2f/UhtUKwsNSfetXMKOvjenntv4jgKiO3bFW1
DD0eTNKv3iUr3UvCh3WcszqE4E0CjFzBYOjmd71MDyYP95MrnC8dvUGl3tIyYeD5
umDeV4EuUpx7j7gP3EdvMhe2i/2BuBygINfMmT+5XoVVhEPS2Ncgrwo0YCyxeW+j
7dgxVnLjJcUlzRkaI6uk4guPA9HZBV/Ry9cMcqTqY2lcOaczUh7Z45ivEk9qRHLX
KbY753+o/IK/kG71Mzf40nE3EeDGJcma4zOdI1vZ4JY5azixkXDFScMpkq3KASMo
8+eOgaTHGlwmBljFiOrbHJbh02YjsRSpAb+9PKl16mzfjRbxe8vHK/WGhff2x56W
crkZ5HubKCYp+MCCOxgeTLrEGkbVwauaaSJapjvIFd6zg1gSyNYhmGDK8PUiV2W5
IuUxMimQf7PrMaGu6nj51FdGvExkvqTwEZpk/NCD05BfEBt0Rnz+U4nTdSx+FYhm
6kHk55hGhuAYwRK89F4l+QpfGSoPir1kkZB6QHpXPrBtK0W4haAk2SHB3upfOnWx
LVvptTsVA1fOacAqs7Veybv1zfjgTYWxZrZCzsGal99y9cK3oEiGyAIz9Vb0Xl+m
LrdFvldtNdztRYM1Ay6SDnJMS3beAei+hNPgdPWG6ElN5vOKY0vnXqxWCY2uHX6U
dkDkyKAx7DqrsnRCJeBM+bjgkeG7UdppvqCovf2eDLCGjh8eu2ELRm1J/4LUx1Uu
mYd/Q/wB26CBeH0wn4+acLaz/uJgyOwZFJqrODYa2uDaZ8Fybzcc5v+Tv6CfEBd4
vIaTUHd1nN2+8woxN+HmAHe6lRU01flwudn+YG+lDTKekL+KQs+Z/wmlgcPqxAai
wiDVsM3Q2K+G6PkiCn1Wa98KMuwIiyVsfdLDaCMcW9sxF4NBDi0Lf+1YQBvzV+tH
p4IAf7K5DVU3ZTKhTEbQYSk+u+NtMhYSA6Ui6wrtNOzxDkWSEWtN0PHCGm7B803S
1EY47HV0MiZ5efioBd5Os2pC+wTarzgKYykj6ERShrLt3ysoLqOu3tO58UQQcR4C
po6SHigW3nVUNtiXdpkxviFHPPYX4GyX8I7hqwNt6iRJpcV+k37nUgodrVe0MVaz
8/RLYIg2hVhUewE85y+qey/7nmX7rlmoabBG5rXjkwGVlDLJB9r8mmf9sg+gETlJ
yEm1HozbK7UpvulX/VyeGTzHEyit/qgkWf+/SwCUjWnMivGQ8Xhfjz2kFaIDOpQe
Ws9bcdgzHwR98km3oqFOsvkTfItsPwisvZpULa7sIc78kwH1FNw8inzuTIUu+9rZ
rdxsYWnPLPlhdk/JQtBFEh9Hl/8K8479vV0zcQ+Jhl9iHgnTCnfVgZfbDhE9KS2v
TwwvRu1lzbeX+77Ll6CoYljjqQl02+0NM65jOBliYE2ya/9WT4cD3p3h0PfkX95g
T7oxcV7C/DM0B9DpJIfMWCBSYoD8LPrxqXxugBf5PXnEHjatPTFWJ+NWsLAM1k2f
MtvHG9K9a9BsIaI3P5mOEeUzvfaUAZdEnQePl/6I4ZwhnSJ250xMDtlBBCH8Kz1E
IW4XXeHhHuWaqKR5jUoqxm7bfkeyQSGq0tbKhAK0fZjaqs5ynS9T7pEyLWxDAKrD
UVMnhBRFhC1Wn8fL7j9EDI33/JQI6O9qb9TtA990NbWVx/AQScXxtxxuOfbKCjah
r5l6DIJkIPi3LUJWufq21D/QZmc37pDA4vTC03EJOgIB/rnKWOtakSSIovLxFpxZ
s+TqejxFnPuGpSQlFZoB3GPNG3IJWEHBg5oFCxehn1rGiAD/UISvmn4j0LVbByOa
KaPiH8Qu4fO0aWAQKNzIlwBfO6UMtbZxLNRu/uDJHmZhcQeSEKwHLoenD1EyXC04
7JUIa4UvvXhajuIbk0U2udLC8BCCeMs/BV+mA18v+ZWTtKTZPE5D+eyMbGb5EPFR
xThHHY1bYcz2m9FDLhh6kJyMx2TJSmiYZNNwCVGr+C+LLvSlzyRyXdTiz+bP4R9J
l7JQdPrXcYuHE1Dat0zaU4TPeAqKDgHYSvyEW1SCqVuiYcA9i8r8iLqAQAbg8wf/
Qo0+zA7rsTy1kratUshzSRN8Wysld8tyYovbDBvWP1tIn1hlDT5xatgPfvgXjjpK
QelaGRb6qOukZBbmj23v5sLiBcgEwgd3A5Qs/FXKSZ6277lb0ymMimFIcnxWOCeo
KtxS8ktgqVDv9ZYnKA8ON7R2e4iTDukj/Fl+pVleMymIK7UNGftOEH43dgvgDTtb
Qtd/6oUzv155/R9z0KDba9kT7KcoaRwM/jK7JvJaDN65kqCErLZtryyW3NvZ+mwp
nyHYDiLfrkFVWsKhNvGZlxj79ctj0I5D6inDxS2cKADUJWgQqKDPCOy4UXse4g7c
ktsZyaAgHhs0M9ncO5Kp64bG/c4o13TpBnjjGrR9Amb/2lQm0plR76RT+IiFhfzK
gfX9IZQS1KNj0+BcW/BHtF2v6+JT7bzjHWR/dU9tgvnWEn6Kk/bHn9iMyINSuo1L
HfKb/z5l6rUfBidE+nyS2tWEvGmpPpBU6Gogo5MFmkajUjXTmFm8uEfjyMD10jcY
qKImwBfQNA2F8G0dccZMgCDJdY2HOoNB2+/O08xIBPtEv/v4gm0qS4D5sfDrIIPV
K2W1i42tai7nnSVystksThC0Gy7X4Cla0hIYe3MQsGxjonO5/zFzLHjcqAHD1mKF
8H79VGdZmUfv8QvJj1Wf8MmpspeAvlHN7gc/b1j+Y2ttT6kpRv3ZytTlPyjmVenp
g64uM5xxopVIjVPlpk3akFrHi/8flGn5Al17qSNy3expoAbdc6WPkFsA9mqVTTej
2bXJbE3mSE5sZ36u5aliLfB4PIp/HOAFyzs/wBC3wVzQsr3Nrm2C/T3NPfB+yEG4
XykDrEBJTv794PAeQCgoGCkbxpLo8q1tpgojFkLBHcXJ0/pzW5BnvW6zg4C1BshT
IxNaDvwarmsxs388BtkGjnNVV1Sm/Doaqdts91NqKtUlE3kBVMnh7QWf8IFxETVF
+QP7EqjtIqVaj2e/d+GydQagrVsfzIomq1n2Cfj0SmUlPFU7YGzT21Yhv/bqL3xc
/nthgf8+7BcM3BGKy3iyRGPMgW2ILzMRf6ntkW3eMwxr4290t2iSNfn+p5aWTMfO
4bjUcLgHvf9QEdpg3hDFoFmDrt5eyqPbLQj9luwIZnyzzD8u1n1CS1sY9QuMwp5I
rZ0n4aIJEGX/T29UhcXym9pq/VRYlugUdSO29JISrQBm+LwEn3rSIJOLsdmAz+VX
KCbWEKE6KcFNBC2OzM7DZXcaibNS6l9K4E8AzcR6MCMC/IvYAccRUifkjhrFSuVo
bJsTONZH8NsP1G9/EoL0sNvi/bSeFi7BXLnc0cK74Z2jRcrJXuL54TYgVH2PFo/C
jejhMs2vPa+/nD1JR6g8mnUBLIbts9sy2jSx+yEcKipMh7lngv7Vqt2mH0r6gAiL
s4g9ppm/OaEL5qwxiHiGdhU0XcRh6PUAhyS25kz0EjuQ+yoEYTNUTSU+bdlRfOe1
KihUv56CO8dpwVk61Aq2/naPpYGyT7kf4526owGf2sE3I1yuznKmfPbDpWudHEhA
IIZKeaZN0cwihkIVYbfk+1zMUoP/8r+Q366ddUKPdilxWaw+Q0IXG3tcZNG7I4EA
PXI7Dgc4AIwf47988qMEy+yWTsoPHLkvApFe6UDaf5zUcz5rNjDwkd1h6gsfOB8C
31YQVrL3J0ozvedIA/EJP7qpVmHDzkRmizVbjg3jOPKN0LNeKtL9ZL+2jItuHZ6/
f4Q8NQlyT/b8K46ABOu1A7SH/Sj0yAiprdPTvOxdUy+HwMX+b+kJJ/sT9iCclECx
66DlfnMloS6GzeGeTLQ29G5h0dTLC/7LlfECtsFiLa0Z9YUE3EsxdKPv8l/AXi8d
817mBGBRwAyG80zmZ+If925Y0lelsMUR6bnxgRONvYKF2HJqlb742UGgWI+CdO5z
LZYWyyan/hUqgowHxGa2ZUGwgirq2SwybkWuxEAQaOW6urZOrq+7NQLZAzo+YYFT
qBdV7U3ysTg4QD3fco9KYgB9lE9/oOyBbxJVvtAf1vVl93Jj9mX8kp2ng/1PbQDt
r8+EPd/494tQyURls0sdYRIxFJUPFOcsX524gTFSn4EwW8nHwdSjECGREG/dDWOJ
80uRzERXLmlGLHkv5tvTMr3gqSbUuzjatsKXxgT9YAkj3+wZcXhc28mv+kToIIdL
p6Ah6wIrd42B1J3Mj5x6KVXNL88y89KSeFum7lbbcC/Xm7A2jae06TDQRjgQEgps
2FFI9jp99itb9XvWwAT6NPCMim962Zu5KCa41poPBBXyU8Xq3FR3CpSjRbb5CziZ
ndL26o028pCDU0hS2MWeMT2xLzAVB3s++sNCUx47ZF5cX7CcErklmX3F6rXlR740
O3D687LHloR/TM8wMRJE8EpuI3Pgi8bo3yOmy/CylMjIqSUGuLuLyFOZKF2IhCwd
zpbP9w+DHMl4cFWv6EWZ/4DiE0Qqv9mNps5lceV0so4HEg5LIbzpbSOyuJTrbV6y
YOn7NCtvOXfsrsvGhLdM7caXWaJCZApckE5IdbbIvt9Zu7LvcqwHgHDA8rOMbx1v
CgPF3AbanI6E8k9qjz5TVQ5yU6H3fI4JzDWGwa8XeHke4L83IlnWjkZUlEcRRYG7
nalU1MgabKhlGa1DaM94mUybLvTLbyB+IOTGbH76SqszRrm8vui/kS6IxKPBGSA7
91Fo1JanDVLdv2Hpt27l/F0iekkUSE2gCfucr6djfegdz1pZSCW/MSggMtqTd+fF
M+pxLPKD3nIuEjs3n/NKl92JckmxKcIXzbNjNpgbDZiGuH7H3tfyrbuqn+cxIj7S
O779jqFNtmZZXdbUdfSpX7avJjGXi8EtHWG/c9CklZl2dqIF03z+NuVd3LVGYDkp
p5navBgAH6hzQAXuJRhMj3MxjLDF1OyybYhlrYkX981vpjIWoGXzldw5WVy0mC9w
3rhYAzAIWa8NZb4wze15GVo71MoUjNJUTB1/JJk4mRZHkz2W6qy//+hBnQEfC+f+
IO6LQoIj9GB83WA7n567tjrrcUV0VmZ90hITYddSpB8VLP+vsbb4AVac49HS1EWF
UaHxFzMJEfOa4vCTY4fZJxprMXGnds4TZr5XtoaxXTIsOmyu4RPUg8F9wiLYbgxs
kPlWAl1oouAVViOFcPPhxWDl3oCKEIXQ+P7/AbGKuuffBLXzS/LfZFnWXUlPcg0k
YJ+oNI2ecuP057M4PsaWSHwLrv5eMO4bXaF+jzhDML3lzOR97j4GpZZWIah8Bd2I
BigPbifCBZj0Yrg5W4/9I8coGeok1g1c645uTHPsz02Voq8/d6ZI5Wh4LE/YW0qD
tzADBmf+MCZzb+uu8Xd0mFAmOr2PI5zPqLn8TeL1VqckLJDqivP8YnJKRbKKY+4W
LTeKJk+3kBCdixcQiMfUJS5N7GjnSc3PgAi70ytU/s45ExgV4D5L8QsTDJmwa6Vn
PXz/gzTWFTVJss0Zm6COi4f3KRcef5h8hHt8/biuuNLAJ9CLUf5+U4/3qkUsk1xT
0AvWLzlXtGzlxPuDVk2rucsKcbbiKjUV3oyTSD+v5rELBmnutSweYoqyXllaL7xt
QR95t0A63ntpx1QKIzyZS7sf2x7iUKqCNTP0/nkz3KrCr8Y25CenXpMoUjZbp56x
0A2bn5G9u1oRmFMcGpeXgfljtdUPH87+fJWK4GgVJDbXUZi75O8U3A+qSptbo7tn
ECM7DzvWZRdIJZqy6kkGSgLXGQr4epcNOV3NVMwgqPONW+I+CutKnDVjQMIMkOk0
5uZ60x5sW+hqfH7iO2/E+uM5p8ecSChExPx+kfyqunaUeWnCCJTHTclI2FVCoNXe
Ha4mkUIqSLmWgeK/Y75sW+DcS6D4molLrL+7fyqKUPn2CIsZB7wicA6v0frgRr8R
RYdNChs+4hpW/OcS1zQOfrpXAUPgnEutzKudty7auWM7d/wbGr13X0sGadWurNeW
WVKzzAeLhSBPE5wmblgH8YOmMr4ua/HtZh8JSH/KOcqE0AYYNdPs1StkKS/oQjNi
k8QMR7I+iaTqYF2Ga6k9dOe1qyJxYCl4VntODULuzFstgT6nkC3djffqah5uBlav
l0FqKnZSVUIOf1KVPcPETji64CDwkGOFDf+Wjw3rclPvAKE4o79TkzsokgI9TESY
YLvPU6KOW5IVcVTGasoU8qJWhTXT2SKvr31Hm588zwb41pIISjxz5H264dPJSGxp
kjnFpM3+2n3NfJMeDJ7ic0BhkyxyribMfiwbitEJcvQqUccH0FGyzV9WkbWnM/Gh
D/0YRqgnuK3KnbiQ3gDiT4Z0TneQpkDDs66wKfpNWUIMC9cACYGIqeask14gZuUN
1zTNUYLxHqZXFGwYQOtGt9TT0BEpUEZ3puoveN0iBCjhh0k1bVCVMLC/dsIpghs/
sI8HnMNxFhKgb0mx2HPZy9gLRJiyN38rxEkD/6nUKMfxdsO/sN80dgZWAqNDzW4X
mvSsigc5tnGeJlsc2THFOzeCky71AwljEzBVuxzr0URbwsYRRt1BMWhJ0qa9Fg9b
TmRNLi6ypqRPpSeHwK8Hq3DictSQKNmhRvD79g+6FSS9CeptH8MMNWR4DP3dD9RI
sJFlhS2I35UkSO6oog7PgwDXJi0BKAD6dOP9C+tY1/7cB9O3ZNR9edq1/WPFNMPa
fjZJlSd8L0z/czjBWRn1P41yNc/ydiznOodE2R4aqDHEYWxb5deN43p4KAgPXLGX
lj6dWJdP3EnX2/fUBD6LUH3ueci39nkFFZfIQ+q1/f7lgY/yC105fuelDXEr3VPg
x9qH/0n6481ZQCYDFx2KpwzmuoADj0Xk+pSmLqtHGr+68EHbE6hDAJLjxsCVDoE6
TLXvgwCe45n+lyAAsBCXJ/KPRQYEmgOJiQWUoY5Q9JtAjtvpyatmzUsdIPEYyM5u
hK/YMNaFu9kz+/EaMt7Nuz0LiJ0phqMLJHXp8k4VGBxYM86l9g3IPg1RLai8U3Jk
Sj8fUU8ys06PnfP50sZNGDGKUjDJ1EpC4PVFF4Ryzy4kfOh24FPkQd2msifUAYCq
vV71yQdQ8D7sqL6jr4wKRd36duuQR2LnXSXerfco9GgeL95oQIiPDJOqczYZWznq
shmoHlSuznyqKjqwzHdN6hTF/l/XnF+MvS4SU7xCe9Yb8eEAv5MBD/KL2OIna905
NgaWvhoPwRlPqEPkr5YAreiWEiTSFPw4iq8jGO7iQqT0z0+DEIvh9YsmBk9pZfuo
g6YmVZdubbXLmR3TO1P7wjTReu/9WSb9kyIwgyO7tao9JqOskl6q4YBUPV1xvPdh
c1oWPv0CtUDCETZ/sMp/8381HNiwE/sagI/3PGMEoaAi1m6EDItyDtp8g7qwR90g
gUljq/jp4BNDfDRxSL9IoiideN06664ZwGzBSAqVk7/DtyF8OqtkGuhnWJoa9s5I
pOpwxLh+7bG2Ej/eIkggvfywGlH50+g+A7AmWqwb/84RH3ZxAFm9QoONlUgHqTc6
e9yqaNqXB9bDmFZgBpa+OGswLx5Y4v7s1eh+1YPE3r/7XCxF3C+IH+XbhiV2Diwz
zLOxJ5B1i1EmOq2kEYrJuxwIxku5FfL7xAPbPjmNgLFUWsTAvjZvjP//hVMRnkNU
qxk2ZcUbCLlT3A1CmMuzj3vp0fqR4V5Kr4qNMIrIVn2YcViEmAH3K7vkJVtIEqwJ
LUanmpVYog0zB/zn18GSNNUdDe+9A5BJguV96gYXx6t8u/n47O2vhEsg3WotR86N
DkcNXC65o2/2qIP6yEqlrNhw2lIuS5PYYBp9d979DT8t7G25/wwfdfOcvYpgNrxo
A/DySolLcoAUbNs4AbzzSIVbDquisSMIPaI9osdmthpmEUTJMbfCtLe21mmXiYtB
G749SvSyLN0S2MUETCFEAjVuCHI42/xcFGTLLfwtMk2FxYH0Ev/KxS70KlgGRE6o
coX5g9ET+eSuQLHC/+i6vEYGMVpvmn343sOtNJWrhDEe13tPf4s+ZD30/Kvxgxnr
+RXDbkHG5azw2hHEBMNj76emhjV08xdXkdLGuC3DPh/StKVJaEtX0k0oTUGHQRDR
11IOPnU/g8vIAQrKkFfNCOaREmcdQfMQ97RvE4QTNcb3YV1g1nq139NivFTNy43L
yNM2EKW667WNSSHoYSFrvtLSAo7elfTt2Ez0w9FKzfdzHL7W47xPJy5Bxd+k7+Tn
+wNHM7BGdeMJzVo5yF+unrdbQPP4uVerZan+4ekusaQ7Xtq0S87Yv/8x5jrcyisa
eH1t2FmrTMgbnwOlG3CqguoHWEU3UFXgm0C27isVU7fDuT8q3VbeiLUaSQai7gv0
Jgu5hpDKPdiVcstCTEprFBC62HcuylNxHCtFnqaGYkcTn4D7B4esVqLuEdbkdfpO
QSjjaU8d33gczMg3Fz/jezZTrinEThXK6Uw3vZuB74KcBboAnvyytXfQ4wNqQroj
UTUUE9VvxWYXFmijNcrzViF/hh5ALHeYnqx30xu8chzi0mdF1iB1EWR9vFh7DCcw
rws1qumQzpW22/h0IozaF5sBidepCQGHwxypjFZ/41a6wi/UYVEssgzggtmBpGx0
1f0IBni4rJktupikjJ0c/QV98O9Vz/KO0UiIy0WDpQm0qA1QHVYDr/NbgTqv39N2
vY9lZQBFQR4E8y8J0Sot7Y3ZYGHH+4l0UTpxSFUz0JMUFKN8MfNld/NnN3hgiXPA
YPm9E8PDgtnQ5YvPzdlJyFgcexM8LjU6XXTnoBfcoBGDRVIUdQUli7tBwwJQTwdf
igy8iS/uDucYnbprVIytdIVM3gLjD/mPyA5p0KQBgOscmrV1uRWpbZNHLs1ASDo0
y58Adl3y3ojkEjJSu253ODsUZ3wgAbt5Qo40MAme+90ZLvvHLW8bk85qnNQxkNBF
oH+N/GDrbunpBZSjnXE4yp1hUTdaUhQfJAqik1msUX69q+7vlZ+Xkdna7Iefj5h8
KEtE0dNRF1chTWlxCkb9IcZuuwLu3tsyKSCwiYVwmeoKHYPLIknw6HltTS1IACEB
PIAQPr0E5w+Fbu5HEtH0axUIKRUWtNh5j+yjRovB5lyiwBsJVllYGJFTB0dgEHsP
kCpsK9SCZLJni/8/326ZyXL4AF51hu0I0cZWvG3qv4kdPh97vmtOV6UhEQF2yXje
v5mF1+XavXBrg6y839qxLoYq0cbJSYWfBLIk2n/mpw4NVgC6QEWupj5bwQtmW9/0
Y57+WkGnvaSu3WpnqdusjpZbv6m9aMNM8kbgJwyOav0UZgARl2lXVaee8zT7NT5B
i4wFOC6ho/NaDCgwFBqGhDh+2UrTj/WGfhChjs6NSpnbJSL5OIJsQxG1YHERoy1L
hVRJ6CJsv/XvIA2Q7ad5+Q/zaR3Rnxk6+LB6E3fDzCVta5v9/hLS4NVxAMMxE6u5
CYPX6+VuKBJtnnD9uJypHo5lUTZVBaUlVbE6gmfEeYQb8O0J6ImEzLQ/VZL3ZUn+
zRNYnzVraEqa/Cg/OeJW97hA09eDL6PzJm0ZEJuqwv0UHRXoqkaRAAMj3HtCzLJQ
VxXYAHLyzgfcCaevDHvsiKES5qOlnNQuppDMPbbT+cATLzudt/Adp/KQvVFFC37E
O59mRff0016PMjvJ7qJ5BZbex8uJF8cKeVZtrRcQA5FT9xAYBkZ9qSnWPGe/Wgxs
NE7fFAGkUouxK0luecyfP/t67CzkDUKnBpoFASro4MnWI78Vj26tC/6gZWmOaUmg
aObB4BWT63slfG9eLYxysYJTnDs8+ogt6L+niUvNEOWZoM8lq8Vtf4/XAlGncNsW
hwBDh+1k7fcmbo00pcjYiQweQ6VQA9pI8b0eYxu+tDdAWjPowaUacfQUEoBzUTDi
H1Seh1NcRWC8No/Zi6sLE5xp4G0s0VMhX7KYq7bWjecpqwW1vickysglOF3DiTAg
leQ0xx3oEF5ZknfYtbJ+gyZQ9PtwUeywRoPAH/TtB9AyAZrPKbWWLF0zvKrobpPT
bsm4khgyQ5r5J+I5KPMw0JBizA+d5COk4rDrdA39MZHVT+r1r2fyBnii0sSYgadr
ztlTC4jmeuATVnkPWRavfUoXiTAU4Swtw4ZnQLTl8PlsBFEgErORyqAgnkXcOwvl
Iwa8KOCqgM02i2jPWxWtDhv1FPi2FiK/Crjk+Z6fltp1f/O9vezhw6BFxfZPChRW
Dcl3/nedANfT5pAkoBxzVc1JmtwfF6IR5Mg9NOpa9dzbqvTaL9pzp0FdPzcgyiHC
s/8uMwoLDWJsTenXzFiyUSTfw+7e3+XJT7jHPP5klzVjZdHIQxFVCJFFcCbno4/i
ZJ7TQy5FSd85KKGNhyLb+aC/c0jWKd7Z/+CvOcHrx2btoi+7cPIFKXzFNnllx5Ry
VXJQGZ+Ct74j3ouOhPN94U6CkTQkgnR/DpfF70mYZAuQUGdsXZTklVHAyZuqVjrX
TOR0p2okWKfaT2tpvTtUD5fom86/k9tCRMfseCYE5kgUHNxLi6yjdA5krtUCgHLX
dFnFqlQ/Vcb8xWYTRUd0WxNVOLSZA7PWKxQKHrqhdwHeLJxfPHELQDv/+jsDsnif
p3hBOt0SzE2uxAQxwAhGxNwyxWbcQyyognMEBrvlbYSjs+q2H/WVluYDQjs3q3Xt
pIEE3wXL9gfRKItX8tpVAkJOS7KsbF6ovjYvpMgj/NDkO8SZ0ktQ5Ou7cr0x5ZY4
f12jTTgWjnsPpvpC/aiDnNqF8Rc4tHASW3ZS6u1TZVd7J2D1pS9lgUYIKo0tT5GR
xDZRzbZFOZ0SvZovoEhivxe9r/5/fRTlCAHBBsUMJ75cERyFtgXeIQmczVLDmWZC
Ev6AE6IfnxWgTSPX6EW5Iv6HPILDLHM4cJ2HfYrH10V35vSZSCNbVi2GOnwz3OS5
uaVQenA6j35LjD6LVRU8mD+u3/RjGxm/TafuDGwzNsFKo/8Bq/i9cAC7M74owAe7
kYlJiI1tJGFMXoIAjlcIKLrJsrxzn7RdtRskcaF7LQYV8jsWq47heM7+0AJITAz8
gG1YfyLu12y/JMTpN9ga7DVpk+CrEcNZ0C0C0Q84xE+HiA8Jz0nTTuJuFEtRI7IR
HqLHuLRbAX+E6amb6idloe8HXAgnng5uo+XRSRneDZ4l5aCFz0hOjHmAcScGKvzP
n4ICXYeJLEXjkIqcBIzhEjpMQSX8uYTylBJT/Qn21hDrDFMT3kAvk3YN9Kc+XFD1
8HSk6R9QWRQQbHdeEbotymRhImbN6o+QqPakJ+jd05JzbssfPdWrOOeFsAqrPVwh
R0oyK+itMq9h1JDhNFYFADT8j9/OuOUXrlgbWRycCEm07KGpHFJ6mtuWOAgmf83B
Md2Tx5YWRVqBd15bgHLiN0afwWhGU5QxglqQrWc6ROkhfD9EYW5ipFXNchPXAj9M
1ZEFj5Uk2WNw/QXJlZHGpo9Tieg2f4LkUQ5JyGLF1JJueJZdq0dEPvekppM11XCH
X95RK8ViKT+tgZdwHuuW7+mu3B/lws74bKxJpaNdTqP5sEz18f7eyncUXZXVxGa5
1gD8PhsanwQUbhIlNCBsvgb0a83Qc9zZdp91iTzzcu2NToq8SLlUO9A+IhWoMxBo
3cYcfxhxDHbU25ANs9LMjV59oZxexOE40dwoWKZU8OhipC5/qw7Y2zEyady77Dek
hrMDzZj1BUvkYScQ9w/Pb4Pr6TGYDWrgrNafRQbYqJ2dc5/eEsYAOA659O0Nlgff
1OpL5/A/u57lFXdEIY2C4Zh+7cA7QH4FodWx8kjL/7OAE3+uMrbi+Xp8NPSsHIKL
FDhMgCfzuFaKbol3SyzlzMU7GxfmTxk0C4xu5wtJUP3hv6EQyW2FyxcAk6Asmrar
UMnR23FDhSBzDgCnW8uDcJLb3kC9rqEygS6wcMfLMwNKX5XBm3YihhZErMW6bUVl
DciUy2nrmPBVDb6868+1/YVLlMkcBb4tKKSic1p69me5zdT1r3usZyFQupyA9Aqg
2y7HjRQRlps8M/sl86cVDmBoPBSAvIbqTtUKdgaZ2IAmjvn321kUO4N8TAQ3rwgz
qnTyhSID+jxWQhkZGAvCGCpV6I2LGRuQUyU/p7Eu35dTm5LRVICcXpsttkkwRJQQ
3whJ5BBFK8gfhLAPy2VAnHiqA2lEFVZKMYzP/BCTynE/jlvuSSeRzRmUiDCE78ol
lJZesH1+nkHcEYl4sCWrpo++WxdQ7x/8duKcKZ4ShnCThEqIi3WwAMflE3OEYraL
pLyJC9Ql5lEmMI2K/C3sh40jLTNU4p+EBkPhAE+a+3JF85iakMN0tevh3ZF+FXqg
z69yawzGgVBekGblo+OkvZjwa+5RgsH8qJQgKsr4aTZI1lSfGsZd6kVj8p0NYFt9
Je1bpc9E6pL+T8TsJ23aDL65J4VxesnRhPKnhmRVbprj6MBJ7/Qt0eJ9Ltjtigrx
KguZvzhygQ0mWZoVi1d+p2PBc8L6Mq/uqUkhf/3P0hDai/gPT8zwoTBBpkz7z3bb
zwKzHvo+PtoNWACQUwXB4c7Yk4GYxQdPef1Fzjke/l8m+RCnYRTavD4hgajVSs16
HvIIzTIeBcgIA178FoZpXW7HvY2uXVJb8EI/ER7elIYShMHGqlcUejV/qLwFg8NB
hZDb23KO77ymLFXET50wybo+Bie6CxFfOQY9UxAOihpM/ss6qtzeG5FQSjMKakmt
qmYdxVzhckCQI1dyq5HU/vC4jIvg6BSdsc2V879gUMVuoxueoFXr1IyOLHwjrGZe
Z4pTCXYpQXSyr1yXfnzM7VS3cLZcIVOc0oICxZ81nZKMG8sjgV6y3AXP7YQL7nKz
xew6yh5HY4DZIc2Q8lZWlsRcptaywItmlHHElY1h6f+6gimw3p/YO6xbx7Ha9SKZ
8lfGyFXqFvtmLOkFkP0mLMxzws80KDsdvxozT6CzXGo0xu0VDB9mAcgRahxp6xtJ
nUg3fc6Y3NdrjeBhMNV9Hfj5VDLls4c2BVGr4hQs3VGvdWjO88bthGtzANqc4E+N
PoAPY6DIDJzqyEvkX0DQeipod4tlHl5aRvE8yD7DfmDSYTXjUNvnqldyWkJIgRfa
btA8KAiuWy/AEZuxR9GN1Pvm5tnzt6uaNF6rO0O9VmJ4c4IK7Bozvbf02ittYuu9
467lmoWBJc70c5mtZufST6uEwP/HWhVL1r7IEvjZ5+NqHgVZihmLGTEehgwHlBDF
/R2aCiRpl9KmP3DMMe/tFyfgVc3pnNNIMv7GyoZdg7MwIKYICXfDN1D9QjoQxZtG
/MSwbbESCEyvLChvhOJD5t+JxyKL/obR6wf2qS2+CTmwpkGUffqUQNSibAy4Aj1r
sH7RGVXTQFnpmXHAMhshh1eLjUG31aizlvKSYF+UYtsOVso2VY8UyeZJmr8rHGX6
GB71lyE1egQoZz77nXnwsMHI34nyQMxVLFuomJcRFDNY9fFhrtXLDP7BA+WQXBDt
awhoNxYlXgwMXQEVlJg+0zF5plIiaC6TfkNh77bALNufcRkDAKEKZk/YK1Q+ocG1
yiE9r3B0Lv/Ma7IgShDSHbmx7zqlrMOB/7E7Kw4M9tlhR3yXsbBeX295cOOwRWEk
twkgok9eJG5RepKJyICZsQQW22Bzy8qtTicxCtKNz71C4W7M47ovNU1KaEbgh1aX
wGQIJKjcRPiVDKn3j2bpPn+d2FxoHRHlbvLYCxnKWzWEvLNqgfzKp9n4JzS+pZaK
pI6pB6NSO7zBcKCYDrLoEQCqsiOvHrkVZmJR8f/LBY+OHUDmmhPGQvQIY2D25Tls
s3JpndtjI2hAqwJoQ2XgjjD0m3bNADanr30zTpZ87H+sg6tfQyUbakVxovA0LrmA
88lLn//MMPNab080wGjQ1C+ZhKDeXHc38Cwjxg7UC6et4TSEv8+vAq8zut2vLrhm
V4+dnYHL6n1tYTCHXMdXUhtxvM5Ns8HSODEbq2di2Qk0zgONF6A+mfNHrHChOeuO
9fZ4pp+Zhw/ZTOEO29X2uD7vTL2y7GToPsOep71HDBhC8TyhMkdz4in0q91xt9au
5u2ricDttfRlWTdlhrpcqCTVYEZHDOi7SlhozFMIMp2lDIFpk/kzeZhvyQNPn3om
LOi+R8e5Svfk2P3bGUkSN5FAJjzB9WZBxfMq5h35abhuseuNZ6WwbcOO9KaKHR6D
iUhW0Mssu71j95Dd1Z5NDexPY/q2QcMamUztCnnNwRsZek7vTjmEWVwlJJrHfO6R
1Eue/re8O/FJ16CauZZupA8XRWwG7Vp2bY8h6zGWOIiuWzitxmC2oD6F9NosBZXb
i0N5D7LNldRncGa+VQ+h3I8O/xF0+5sKOpeooXHPYq1nKlxcHG/ltvq8t5hi6l92
p6rhwzox3i8dKfsqrYOKg8YIA16W/Le3yyoTbb0ti3lW4SAp0jTcPXv2ct/IlV5S
WeZfi4lYNWfvTJNWClu47oqvc+FS2dJ6eOgvKWszfR6l6gFcd8iilobGrAMV4QCY
6Zjmo8WtCXHNYjmF8J3uFnwQoc+OB0QGwPFP1JJp3aLVbJQjvIJf5bEOl94S6B4c
j44V+ltEY1iH322zlBAiFMd6wUqB50Re2gP7TevR6t4SwA2DiVI2jxdicLv4I0Eg
7wRckwd7olrWV82uhMGpV/eafV9TnO+/3FpdvtBeI5yVvI5YCMQo5uy5b23udbZr
2fIl5zoURfTGihxtlSuR2L/d9ENF1s1Gcwk4/AubMmOA+BulicjexRrp5CHnCItR
VPu5YygK4BiqTukoJrcuzWrG9nAAAnPRnuA5a6opAk8hEGPug7zgMOm2cSwPMlBe
5na8ZjR8KFErciVSSLjQ824bgso08cTBd438cyyD6lMoLvuNzen35Je8uehZIMNe
UlAqhoKdLb69QGn997h1ATOING1KfkxXRsxLL5czO+n4pxwaUp92TE962Ut8Ow5d
Q9U94pSB8MZFB1bb1mH7RILboJBlVuzj4uiIIU0otL5M0RIIwZFYGLM8Gr/KCCbD
TnkZEk+7iVRIfLTfcaN3IjoJAmQ9xg8+4YQlKgsfCx0ZAE+6NxsppdJolJr2lvZ0
mGKVV8soHP99XKGWLqDWc37jzpljsxRPxw9KgFJR6qiQUDb8Mazn6Wyn43x0Vlw3
TE2zRbZdv6XJiHy5VW68kBHahXVRPuCpBxG1jD9+B4wOMEcC8d7rCTFAsDiQhKVP
RtMUg+dZFXgaDxEdz0cJNyKG64kfYjRoU//R+1F9g00yG3lOA+MKMfPjTU34cJTf
PhrxZ0ZYunu3tE9rGUZkGeRhZZTePJMGPlA3/4sxvUeb5Uqa4LDJS/NbOdP2rgAr
hO1Y+HUvlJD4gC8AC8Z6gI4O5cqAeVMgfXHM32zk41ousUvyuFOk0i6LyeZ4Fru9
JsQ7610VL+RaUPVLvAqRcf6lW2kggkWa1jWS0ES2q7Uw6txYjO+jsULaXQh4gKF0
ug3ac+zedxenUD6PNVm+3tuv80c4gIBSDS+wRpdROiYU6iT31BT3nd1uUZwIWQ1M
QVSTSAevIYiPfPrAIFGtLKcQyq4zmFpCwFHZ93atXHLNiz+m++IpB0TH9E3SX2Y/
59DrH34H64QRcID4DGDDr0AnB2yoAgVAp3o5lnnupiRwFkg6Svu+yZtdtChMEN5p
wcEsh1q4W0aIBWF0AT9m3huX6Ly//sJSZcSxyUdyEpCjVxmFNzOQAH4l/A5t+Lrf
EPSj6WxpqxEYfzKWOqemqxnuvc0gTntFdMAqyyW/srL4HIx8yXQqQS6KoC9vMAsE
Pb8GwzJc5uA9ajYGxgtR7oBUL2Vc56jwMdvgjTqsk4J3U/5himyQfs/cg+522Nfl
MzyIiXSqcxMmWdvj9WNstSZraFskf07ZNe0+3Nk/fHQm/F2KPFiIDa/LydF4EoXt
i0kAUq1y9W7ML2AxkbC2cBslURSYgrnxVeorLH4XP8Y5+qQvPZrHmT+N8Qot5CjI
+7kBc5Wza4s86fn4TUyqe9j4OulTmRDQvPkXnN4U4IP8SN0PJhT+YaBoyL++UfGt
Lv2tnJwvIuqBtqOGOsRiDXdS0jYdKZcUFOxCBkILPF5hZNSl30ICYFG5iZRf8S0k
CslG0MR1AKRtAtNHZY9bo9aZd9KeTeHebofJgfTX3+Tm1JX7hOJo5tO3Vse7hFB6
EeXc8CTgRgmLMw5mDttOZoN5N8U+GvT5OXallICJmoJrqHWgAaH3tOruQ357zw/Z
DNfhwwaVyebBBTTSMzmuDTM3FLvWGNNOn49vyc05nkN15rSFAyVkO2OXIJrnSwa8
1SvVDjw87BOPMilOqXKbHVMSLFMCnurgSDfmVpkbKeDmv9L2HSbGkwH71d4sqNxM
jx7QMP63qVOT2hM0W/QTXaOQg9a0ZRBmWecMW1mdFX4tBhJVJKyG15qDb8D9x7Hs
ySteNqBvfbKVPpJ5C/hnKydoGMcr6bLjQtWr0M2mdysdDE0c3z6GaLF6Hx/S9bRQ
AOMg9+t5p32x8NM0Uv8lyB4WCg5IQxiGmmDVcXgR1C+Q8pvWJ24MBySAwiL5EdAL
8JPNgbGiH8FhMBwfz/AdPbLfOpsVhB4D1bHyKVLRzi3M47/nAlUdFD0jldEJ8OqP
D1BJT0nay/+Eueui/snsER6ONbG5YII/+SKTwWGaxAf+BZ8302ok0qEf/2seiT2W
ELqBHmdsdtPmES9sNjsD0olQy0XNAzZ58dvbHz9GMVr+539l5Zl3+RHaPK5oEWEB
BvIhxXqMYmbNPXuFJT9aEZ7r6mvOReGRq1qIMHTM7tlcekm4+EuXxcpo+pYTRkcP
mTfsAR/FahW2EZpc8hYG/KGQZrwaIZrEB2u98Q/HRaG8KPFxl0ngl/Jo+BciLxlI
kIRnQsNecgz7suNwQU9+kJwn0gdFWS9N2NCKm/kN7D2880duzacX/26uoZ9kO2xm
eYi/gF4aPzMKkQSBM3IMh+kCZp6kmuUrZaYfaD8oTDQ9vCG7BGqwScYSNrGiEwfQ
FMSIzO1csvIpHjYDcCCY67HcK/pMh5hxQZPjt7xBO+6QgJRiH6rFDKkD99F6z6Z6
YvMr78/zVRVMFRZu5FJMalQ4xZoyLxdcGcQ5h5X9vBfAtE6P8QaSQc+RV12uBcQv
whq0vhxUKytubDw2c+yQxXBnrkEtDI0fhXZZ9cqkoiCglGmNTZNim/zLcNC6N0vY
Im5SmJhM3iYufNAh/VyRB2PSYg7R+x1vwuM0/qoks9rtBDJsrCP3E/ShjnoL4+a7
gp7EoifC2b3TZktffPUWUJdinu87JzjYHfMOgRjwGtfACFFd/pGfGWeQtdfBO6RK
drFaDNYQJPNqf1AiN3lVyBZU0vDpeOJQ4WbbqQ5q/WMXZmh+8CLpLnnGy2u65pr8
hwn7GZVWsf8uSeBQ4Yini0hhYClta1ieHzgkhDa67llTeh+ndoLBHULr/zOjy0ZR
fj89CHKfBs/1NbNkvW/hLHyqnnQQPsHnONIdMa03hIcYfUFUMFGHUiA9e2OyQCSQ
kPqdOmZyILXY+TEZo0j+sPLCRTz0ghkt/RoShfKh1TMvUg0Fk1AX3lj2XGdzBWNJ
Q8DeGu00mjcNF6OYWB9+Qlc8edbvPvN8XKk2sjGvn2N3a5EQyFaJGfFypPyLQ2UR
EyWQhOoSIRaTN8Q6YCbbEcMrjuS7m2u1gjWWlonVMrfcXke6/xqbUYLwDxxsntQi
hOdxMN9g3aSZO6lERUbWE7NOlgmsFcbiERBF3qcnZU6A30SCIYnBnZBrMXTzUsH1
lhf7hcIzGnVO8LKjFqv0g5hPgtpCCOLy1T3Y1r3400saXtkhYhsO/25JBGpmsanK
fHxSNdp9PJLBZXEZdTI3jbWFenFfCvcUYrG8txrq507NxQLKmDmXsUKfmBOuWtH7
7UE6Hsfs3zXWGAT+K8TZRSVF1jbRE7gAQ/GEXbawQiAnzcQ3pvIXNz3zK7jmJMy6
Sa7OfcQ8eW3qztNjuADrW5NR5V+R2TqFA6So+e1liLtin8/hlzYCmlK+lqrOEA+A
CUIxkB7C6w+7XFkXkKY6Qc2R3iqOrIxUbgiPQs9ElDV91IPdiUYldeV/bV5UecjB
++HHSVF2ryvz24FSUXHjtaiI/GfL9k90nepyScawELy2p3qat001sWJ/nNs+A4N3
Kt5IUE5qO7JsgKJFrQUyKmg3pEEblH1pTddApFirZoAPvc2vS08hHq+ss/bLdzz/
+9F4NQTQp40LuewElG24ge5oYW64pU5EEbpNdHQLe99wbBJCm3rbMM/QC/SLx/tb
7Ctg2xvhpj2YGJuELRP6TierJQjO7KrWSPKXxKzq2j8sf/ISvu5pyVU08v1htNzg
NXGyv0OlA5neKnorfe8HS0V4E+j5KVwRooSpEiRr9LQ7Gi5LcSNkqqZD1KWtCPKg
krzv4zP0n5rUu8DVrb9wdJmzd3mfEoLnusRhcADc+2iEsQ+NKs2zfhKKHFsVMXOx
i6AcA2alsRbErNECfQgP8SEajjof18VyUxScRShvw9UovJm/KHLhg6WkhEtad4lZ
OkXleLDoJuag9tz2VY6BleOEM7Y64PeUZWKVPS7kcyGUALHhJ1SkwCE4mV9eJlUc
u36nnG532v3uD0xaUUTWEcQ3oBDxXuwFC7RyPAcBfpCKrtjBsFNubX9eY8lRMc40
8EWC60SNFcrnXdFVv+QFXitOLlj1LrSGUw8vSjVX+eIeZxCG3nDME4sPP2o/FHJ0
u9xo//Lec8F03hOkUZVRT8p3e5tJ49Kbe4etOtEgjsyz/AJU1ZdeYHSyx87AMZKE
o2R1+70kd8xrQTBEyYNq+XYa5DDgxmiK2bL4Mlugp/JSfYSYl0Z+GDfv+K0OwThq
d8kWco/SYuRXvBQVV/FpDHN5zT7zx/3w6hVkexreypvdwbwTBJxSZFxYs11pqYrC
ePiDiXgc58KDKg+QEq1Sakq+ajTWvZ/pd9w3anFIXt370LUvwgDwND/YQQWXLkbs
qim2erIzPvKTA72J9DLZv3y8PDsp38jp0D2GSW4c3JqqB+i+8OUbzsj/s9Qbhbdc
41DIzgQg5LLRMTgKSOf+2EIYe+oJE3OQKG4JF/sc8vGv4HyomPKzmrISCZEhwSA6
pxhHpZdL7IoAp9Q+TcL9RtErkemqlWAhLtF2JVam5z4xZOfnRpsg8nvv9LhAu84u
Rovjvo0Eh/yOeb+uHV+FCVfLVlKtIUJaygzYIR9c9dbm1riXTisMToSJfyYx7wxA
F6g1e+p8sdf82HAVMES5NKmM+Axc/w4duzwXnqhG8/1lXOWlV75B3aBiKfQtPV8l
CmjjWTQVupzsxAD7zQdOynOi6EKv/RablUpBTjQRfqxyQdsFtvPAazuqkkJHgmV/
fmLSkw6n8OMQ1O/RD2KloY56puJy0nVmzJ6BXqjU++AUp+MLK47Vp6CyAIqFotwl
Mg7ynFXSWyKiBA1hjkSlzhcarI/7u/RWDRpu+MeqEmMUFcLnAMCgZYNJ46pwd6rL
R06blCmKSsCTMvh4/FEiO13Mvy4xVlQK3Tf5D2ddN3+9Di3xjuup7k1sVK35yJw1
KjU7nT0r2as4Wy36JOCUShxUA4wCNfc2onAuH2+Op409pf2heXJwgZ8Ei9PccyRr
MNs5ud+Q1WDbnhay09I/4fwMANoRS3tqxpWbXzGjG+J32R4z07I2TPdj9tJvVBBk
M3ICF2p2CVMIca61QoMfQN6rn+/o403dlVK2gYvz37ofu4tjLCwGoMMZEDsbeCF8
/RZ0qtiEi+5G+uTkZXrkhMNGBh5MBS+o/zac+r3+qbOCdJsQOkJ403rlLDAST3OD
iGhZa6u4oeuajD3YZB2i5fPMAywn1OoIjznQ99KFcx8/OmdJyAMK4/+lsxuECpyd
t6CpdusMew+fvMzB9hM3WMhNqCwSt3q4EyRqwYhJN6X+pbfFJ5YVSTS6mnzOizud
KkROWQk385BEKOaCddSQfo/Rjnjy5q4bsjH1qmyjKl4jQzjtkvPZilkntTwdS3xw
kP8M+vI/ZiK9tr7tmvRh+SU+Oq/8Bo0U1v6reaEepxZpqcKLjeYZpd6IUZ+rCzRX
xkXPAkWiR6U6Vj/8xlYjA4EM87W6qsaVwVQSlYYNeczf4QpM/28R7X5CyiVU/eNb
7pNSDkg0m6CAcUIxhx0M5itsRJzBArW5t7fUN07vGvO+lIUDlfwo4cuSMRXPxfTj
ypHbN2rnG6WYJT4yV7QVIBW1gtId625PCRYEQAoDeBF1q3+RGr5MHFNLmTSqZm/G
mKQlJDuEZx3jMSa+HWNvacjHmV5GH1bElO86cG94l8ckj4K/KKb2JqoMAYrx7b6B
QNQS0+Wdqm6DGrPz5Omir/CUNFFRkGpzTZjEPZG5BtzuPB2gZkITWkDsr/Dou2nx
Iad6b/HdA/C+ZN99o68kzNrI2dnmcy9o6KC2MbA9lFf1H9O7SC1i3+je8X1rnNm+
IH2Wm5vc2l4NukpZmrnmhPeO3JfyPqtCyb0qnVe8TaNSLgHDt3/p7TW9GIB8Tt0a
LB78D2IDfmZLleCtGRtyuDhIo8sPzy+3G/Lhx923W6CR1x7FrEPkcHgRqfazhxiZ
oWcbbPl2/H08ditGSwb6aOXH27xZVEohmor/27uUlmKwXToMGNrdX+dXj3IjeiMl
G9SOwxTyG8ZnkHep9cOu/sy41WiPDOq0qtO6zgWQF30nbIrtBdhyvuxn7V44Avjk
uqab3+0LNZwNelEpmEU8tudTlsRHWUvkGRqbpr5RYCU3IGhaQpwlyVhQr8AXxwQn
7Xf4jUhTru8fog50HMwJ1DhNGl5D89upBV4NScBknEpaaKvmWHMVQRAFjbEVGhgj
l+ij1Y1N8MC8VGTwNzcbjrSSS8ke6bTFUFWRl+Q79Vz2w6j5IOQcLuxNAFjc+SPA
SiNW4UVuLCshig77YbIpVgP15x4nv/NTWE5bfrOKmz9Z+lb+o8NJgYZK4UvoPjya
t7LEfLOVdL1l5VSlWbqRp0cd/i+kngpCo+++Fcf9yPkYA7YG7ohsx/9leB102qzk
WLDjfpVSACbB/qf1oE3mu9pZmgNjMWYW39NU2Y9MBokIxoRk2EVhypRl4kM0p9oJ
pDNka1a1IFacgUzLNd0f1J83GJe2e8WF6wP9nl3/YI1dCsK2yWw5AwBdhXMk+YjD
64uh8//Yij17JCcGySuyxMuGmW654hVUslA346YyBnOLJUXX7Myl4rtzn8scc4rF
Grna8bPoegsWc0l+CvT5p9uIbSzO0Le8SK5TV8Ry9A8f1sVVwtQcj+YmML0NlE3y
hJBlR3Bs68qAdebnvGHHXIt8CCpTQR22MmW36FxWXjjQpqm4cUyKWrmWbSatGzAc
eh88ymITTPsuctDn4te7hHeQYzIcyN6hilVSWkCXfEuCB901S71nZScPFEet1rXr
67uUKvF4blNeWbNxxJ+pL5IXjCAo3Oy7eqK/j50qh0BPvedRxYCWZXJ2lT45sntQ
73RrlqT7VZ6CAMAteR+wkx1NAyX7oeSwkDvt1hL0q5+VjCSdOrzlg6MEEHczCSh4
3/Fq2M0wMVk3CBqwXKRIOQ6tua4t9o/TtKPjcWeq0t345v7wT9CxAwLRLlBwE9EY
gw2B7uJJ2LihGUBXH8wzUbCcgyE6ZSWzxGsgaeQG9suztfEMPYouxa1fyX3xCBLP
iabuPJU3+ahTCa8zZAFgll22+i9NomUEZ6itnLdMA9BNdQvE/kNjS5hlbrsYgzJQ
JFFNpIS/JetjYM3Hst8LjTfVGNO/Ub2C0RJqiwaLpPjybrMyiINa264fSJ2U5aZa
hfzvPQwpDj2oIxX48q5dnsx4YKVAMSr/0D6XuyBTegvpdlWu6RzLM5P3fa8+Kpxz
AvJMg1HxCtan/CrFeVvPxxNvnsNdWj7iEKgeL9dbOpeww42WduKnCz4XIKKP1dDD
LTNYDciFNvti1xcCRNun0gCCqvawSyqtINMwuACP8ogmGyzlwC5TI85Wh5yv6ODP
DaWm5UWgqm2kuj7zoK+reAyalrzC3SjCkuP4pmHL2x4JhD2RJaTGqzBIFjLHKgsN
d00hkBnVGrDWh77SSv3xZdhz/U9/uGUD0Jrv2xZjXmQz2WLPBo2crd6iABxyH/wo
wzdsghud2BD7a12n8i/Mu1RAXI/DTbttM20Ryk3O0ZusvxqmfgrMCJbX5M5SzGEL
mengkGjQJBrRbEur9vWRdyR9o9W0K0Z2RcMkUdmL49BnGAbAQE25G+diNx9t8EsC
abnJ/qCFJnltN6gXltPy+3+7GZfonYkzjWyx01sRzPx4Zv5X0X6MYKXHM3JReZ79
jPniMXA+Ue65IgDRDWDkK/Sh6C1niesb80waDYFkTX72TNr8bOz8nAeJsQvhtjmT
d47QcuKEwhVYcG59CcUnkmky5g3ZVhlmy+E5V+jI9h5Fu6jLQJtFbuACyH/aGCKS
uav4U+6TipN0Qqm23RmYZMnLBf2H/7wHisdCXTmo3fYJM77DSkdw49AM83WwTYjo
FpbDEUIadaFOOA6jCoQ6/rsnaJT3djA4rumfDfpuJ0SEXHbUN827yAe23cqEbuyp
Px1L+AvRL2ewCZzEFTunH4dQzbgzvgthKJGhDAKPH+u3yOBoALst7SPvUopqo8mO
Y6mVEUyiLPvPOE7t9VzfwaIru7/y4cy+l69YnO4QPnPczNK7n05ye8wqYUECc6Bv
hwAWySBp9rUZy1UPaZpGU9uF+KevX8ZJgETMRVCHpZL8GuLgsrp70HJl5hUyHRyB
ZDo8moLkWuNm9vIZZRRXBA0i/p2dBwjbhiuUan0q27f29f/JYrlWRRj21nRbGMDr
BDBWS9SiG39YaFgR6GBogGf3sUeXg2slVa59yGEGRyX1f7A3P1hgjBw6SWB67dx6
Sdc1jqg9gRmeaK5Awou9cZ1DVypA0MhIzt7pNp4igdWQIecI7c/5Wq1RhHJSKYIr
x8SXGEJIbL7b2yUQwPKoAzT4zdmKNKILn4fvrBomBULv+aAnhxTpZYxY+SlblAYk
0Y44qZpnotdO1g82VhYvqBjkNv2U2xH28wjPZcedt18sSR+vnb1J/9nfbivan4X0
+9c1/vHExbcacpL9kxEudr/2JCtAjKh8Mcp/dze02zFgKMhKtUUMYHj7usQ2y/jK
gA48SqXlNdz0eh/iXuOJMsL524aYrMl+UHphq4VeCI9l33pK2fsVEH1cxldAC12m
mqPC3z+Ybk2ty81Ra5huMr332LAgDyDlzmcPXwYxkC5yC5O+gh4efZ2AggI20zbH
WDHmrReJNU54EY/bMAmnsq8vQpiD1JGIj7gQ2jmF7Sd4c9+zZa1yGeeAYNhKiN/m
doeC7XXSwfgDMzA+LpePU7HI5wZ6vgpMTg58/N8DZRCji2naqQB4w/c6sx0FUzVs
eg7LXlRvXBgzxsH+FkyYYHSE/l/V9L/LmUZ9iPzTXVmYicKPLx/AsFLoiw3lrVQ+
lMj7YHYD6EsZbkzU7MmKNh5jj9PQlQmLrHlABy3Rj2Hp9azjtP9eE3g1ZV1pLp3M
nTalyITkjDdUghGy1zNq5nrY56km0IwSxfnClLtz364rMRllLrFZjE0sYGwrSxxu
9GKM7fputH/C50ziAKAaVpw6qgOPKwcMTCWGBa3fXr2rcxIs02bAaWkqP7FsoHtL
1M7yUgE5s4abqvfxQ/nsOwEWL98rfTXW6mhxTJ/azek1U1isq+fEsAK1vHM7aeP6
CC07LaOU/P1CyoHEX+ICnw4BHXQTM8H9eBTHnq2pepWvVH9Jq6/QtkJWnGpdIoRY
EiKzRhR2CGbV8mPeSP6DLNdX/ERWxSoazN8wxh/LiLqvw3m3alEXDdkNxIzhHJrV
xV/DaMzySudy05+30S2s8uAXZkpZGCJn9oSqLrkOhzssPxnVYyD1p82QJXP9zelI
6L5ptWdRepy9LwSHByKiF/EHO/m9St8GLRK0rEPbXltshYQ9o7ZgpWxFC9jR0owb
Vwoyd0TadLEDQ1KkBrmt2taaqukuj/L5jcjH3L/jWSnsJHMu0Ca07LN7gKn3IyDk
Yvf8ujjNTuEEa1iiE5of26oM+jm9q2P9l1q6TBfiaUqTEnMWmjLp08S3EjtwEooj
I7QX0SNCci3jxUV0o2hNK26vgon/kDX7h18Ztx3qsUrAUWEGEMq3JXNAWm4jlq0X
os0pQZhBRXrUY1CqiUMkq2XyD0iXvl9LLsEwG+rNLWn9x0AnxX8jbKeomnVYqf2J
bKh3Soe7b8WbO+tBM3mygdjHquJm/PYNL2N1Mqr99L3ziPv+vMEaYDn3k8fa0NCE
OXD8Iy8W8DSQbGXV+upHk8wHUJNWaXfSGop0O2soK1wJ1uFteSNIjx/enpdqYdyX
R3RcvoTXVGJFxnWCkJPoSE69H/eT/mpu+GJOnqa2rNZX6mzgrSx2UcUfb4BiQ4rM
4vi2Pq6GaWuZsiVtLARY2NnJHiUAxPd7qclIvXTkXQ7s/req9StVc/B4vqKD4NlR
gVXzTTFbu4k10+FmiMa06319zT5BpAraAd7HOjgNe5sh0PZCVtokvj/8rPXiIAlg
lalpJ9CSY5ep0EpOnSKNSDW9q+U1UgpR7w8bnKjMEj5tuwTp5qihmP5Eowoyrcb1
DMvBx/6WfAI6v8vESQG6k6sxy3dXq7jZFtZkJmkpaBmMx+p8OUzMr7QxZChF+TRr
BblmhaBVcMlY/YEDn9/DEJouqFik+h+vppDhmZPdLjUEEd16id7QF9ECiYGT6sJT
JNRTJB8A8VmyaY+ODD0FqNAHC8XJT8E4a/onmhdOYCJrEVNf2O2aUm/8GP2WCS/Q
5oz5cf94pmMwJJbpNPn7p2lb+OY8Npxu6oeJHyIdVLU4iK4hONtx/i9S9ZXXe+lD
EU5Jy4j7AfHL7uldxTu1r95oFQ1CgqCUyC99lobFu8L8WeLO0MRJn9OT71cPgLrJ
EXiOc8JtD4UQGl9b43zH+TYdQW/s2TgTJL9gIdkyxdsZcqiMiZDGlujAfouBrLJe
hcKSOTYb/s5E+2NMpm3b11r6Zf5z4eNI3BYlaF99S/3/7DlLK08ULxTmlEWsv2ER
vlet9tJoPC4TFmIK7xsu09lbISvFSepUaWTKpGD0TKyFxr5wNNWGDkIAVg1TCbli
O8S+RFd1onG9wNC2aFCyvvIvjZc1du9VkPTZyHxY153ElYufQqKX74NfKPYQRO7b
7xAvh/P2BPp9znMfNyZKm2xHQ8aTQSr51PfsCULewmA59jVj37JqctLP/Wxvj3TT
nVcxAlY0XVlkeuvAgizW30G+++T+J+NnmiVl4B4rZ78FtS2erePq8ZSswS2Ttc5V
7X4gT5BHv3h99I7tCJRlWtqFSdPIR5sHn/talMuntSoAri49FqIpaYsMsEDtwzGu
MM1xy6Yh7Wqv/GPYwLnrGlOLPxovJqIwTb5YGiU7gqULKetG2y+tOjYBI1C8zwPe
CyDaLnl/ubjYNAeWBIU104xC/SO5DvhD6TtM3QQAOlVy4Aqaz/MaeTMxJFsfhGtj
ihiyDiUVu27gbj2szflQl5seT19ibN/tQRBTMzd1YrqWlekis0K6M+th7XwpeGhk
0RVHNmg5AQWITJzOPdksONjrk+OK+S5PhkT5+kmWfsFTH3F4PnCzu2FTKqu89Rz4
SBzXXl0HxKWjxUAY8omS/Lqxvn4DDn8cQv8PgPUWYBjMkaTin3nIKmf3ZP8J+4Y6
+DJeZeQ68gSIGzv2kadR8Aka5ZCOa0d0z6lEQ+OrtTy1NQT4HHfhr4tqqWMUPplv
137OQm5XEZQuT+VNaLvR7S6Aad0XBeSp6gZNkRldENA2+SgPG3SG3rSJcLm9B+2K
98Rjo7z1sOWm4aJeCxa2IVigTJrUeExeus8j51KICkfFgDJUiNUSjvYGhoMcYxVE
XJNp6zailm3Awtk3gjMZxr/KQBBf3u6Upq5aJqFY/g4=
`protect end_protected