`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2688 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
EumbC7jrt21FxnZykGOrrQa1pN6qC5rxxbL5T0qr4T3ms/XnRrNVIXM/TcBVqfcM
I/nXwpvppG5z4NsQvt5ONULvgBSw0qyshT19lElzorXwlbxKdqgLpXnKx/cVFzUe
X7YiOY+iiD6gImsi4T7SbgmlyChjf3Tori3hQi9I+XbHty5ttpdjf7r6UIWaf8+B
c7vmdGJd0wogVGNzECvKB78O/+pIYa/Y5AKy5fsxat72s3tcMXP7OZAjvhp3cDrL
Oz+O1ED5zDVvJNJe4N6eISF/tFvplrnW+7OEzMQOvh4vRF6lhxGnwAOcPOxjrkw5
5w4L2EWrRLlNxrqyWwI3AsTESO+EHdkntFaCMAfVOjTYOY6ySe91oABXH7h6llty
KlAga5tS5rKTtgDW1P6ADk22uCvyKRO/zD562ZRfvWP+Gd5NQfxyPPurjroMFP3J
ZOXsfJkjQEmuBDYYbsU9g1VPqWWXk46LtX5j1qT3LNBgfdjCaGiypbmdNByacL4k
D8FyVN8J4QaWTpd/TpHnH5dSUf8nMSPpA6jQGy4Wv/6PuoDB0vsDEP+e71ziKjpx
KMBiBRgy6TxU6h68Tjh/1r/bu/iy3S2vMsbqRJF5PuGhnYAGTN2baPMtewubl9tJ
/pP/41wiOM2hikgGk+/jC7hbWasOhc4VCtxaD3AzW6gymMLrmXVIQ2PHOiNvKckN
V/gM1GQZO5JOpjajFPxQ3ps01JfDalN2bOTbZ/bsUgOQqNMmO3ZefdUDCFim4f0C
j1TibZpDnqCrZ/DRDA/vLHBHqTI1RWcgElwpZgnVrV9Ie3vS+WCG8eoAeivve/Cm
EH+t5+/CrKlxuWzZVWFv5+d1NxL7HDy2R0qsDCLUZdXcu6bnwKi7BYCX6SBnTBCf
4cvuz70Iu1hpcTv1C2i7fpBoITRfvrknIVj/Q1+ueDSaTBOwgD1Z9ogw99+7Wc/b
9A3atfqTGQS86BjIKAiKhRMwmmOoXxyPDEi2bg4MCjdKZwU2agUprKly5qxJ9GGq
thUzu3tB/j+Q4FEknd+N5/1sbDmmv0GFghwzzQHlxLd85OO2HZKt48Urj5u4Z2LY
l8PCatZ+t+c55UYU1mz4ClFoU4VZFNa+3hFxHwJxuPlfBwmw70JtFbGxfGW7drYz
XdkQiHZkTwdqiR49azVcK5+/SjIyEEMXouk63p5rsgzakG9MhSsjz3xtpufFCVTX
i2OLLZTjnymUlcMwmMp6b/wU+6QvOH84p5W6RG6xgaiEmS0/AYpfM7k1LEx1dfmO
lC4huPdZ5XUTQe6ZvFMWMNHyO0SmjuY/05gG983uARV9s+QJ0S4GudedlAt1KVYO
weKrijDmguErGx8/t0gBtEHfK7jOuAIuxbDoWaa0JJevYO0qJUwVckkPsGbpXVbv
sE++vkVcL2X9eeUutUBGPFobMMG7+8dMfHOGOWyKnqzIW3EDijTR4vUX3pPNykLW
mMZh6THupkjkynq4mssYYCd/Xrb7fzviGPWNB2uTlpvWwxRQ4zed24t5LFsMgvb3
hI66y7XkQSGtTzuMHbD6UHMSTwtpM8Uf1T6mM17RrfMnmfD8SRG2G0iSw0iW9j7Y
oN8GN8TFOlS2mgU71MOoSvl+WDBTK91YMLrNoGjCAyyCr37SWbZVC1jxegaebg+4
BLTmaTnJgCN0EAbCjKmeEWDRZ0wpWgAit1Sa5eNKw/IFBfZ4W7CEgEkLwgg1z7FP
engsuKPuRxXoU81i/8ApkT1/WGq7/2JjbcHEV2xr33MErA4RGJYQmH+cqIcschcF
0fYggOToc28ElHQCD8Fd4A2qhFcjVCuZYu2fUv5a+FkiS9iOueajCOmGGUCnVhga
w0JxcLRkevhPceApJQ/mwuAg4fObLrtllBVntIFVgkCi+HKELFH/dJqmLu6PFAiU
uht5JDNOLGX35FxqotbbRhkj3HXJztxfBoUcGRCwPfXvQnxNfYlLqw3H2tva0mD8
1mV7/QtuKJsu3881GNd8rclg+xrcW0f4UmVOY1Fbb4gBcjt1xJbIKfHI/CdrOTvZ
DlYq5VVy7Bw9pYQHXSVanaBrgFfqmc7FPh2zLU0vX7SyU2+RZymZLxb+IOeDaSS+
o1p4x97Cdf7HYNnk7Fbb+/XG5ubWaHsmWXuIb2+FjbkSbn0fUDZtGl+e1NC/p4RX
lcdI6rvNSrPDM09PV4yLCfaXKB2fI05VWqTN5QjhSp2V13uT89O3wUB7qV6hJN1g
4ITP7eNNte01emYMUwVMn0o/Ql1DaQ2wFUBcOmX+T0756oBYscwxx2L3GOEtKaDf
c4mOUdpRPOfSfEgZZdq8DR9Xx+pZ4XQWox7u46GjwvBShF+ebvdS+M3yStioAIvc
9LtewAwJ5Ca6EQ6p9UfuiqON1s5EKKjh789VUBxDKx6NsIkoAZ+JOB5EBJ59zRzY
/rXQ4pCP/4wg+EVIwvf7d+lwONcTjSWFKNMH8OyNd8TQLsBtKj89IPW153CQX45D
z3tM4AEBwPmE5iK+mLP9T+VEnMlc45P74b0rYDRKVIstdwtLsJX+J+8n8kvn077L
CBtJVGigvoFmZEmytdwJL+kgyf14/Lppo8cOviSgwAa1FW45coLJixa+S77hm2FG
RYJWd2L2sYuUKLXKSnQlMGK/LRd9n2l7CCMHGmJftdv5neQCurHg6Y2wxB5JmiIQ
iX+s29sd4ASJcUvC+a1TMM39m16QOtfuGQxPmvx6XdY7MLeDSbLXvaVIRi24iCST
i1B5N1V/VUoxdK64CkhcSDiqHBhfUgR8wipFR/kWlnBdO38Qku0BknSbTno1cvWE
P1cshylWsoSIwEJW+IRRlNbyQ+rz4gR8Ge8J8lqvA9JMsguGxkCpzCF+EP9c50zR
f5XLjJslBt3BuOC1F4TsaLwWUzdcbMBRhM0EFZlLSjFr3kGArqS1xHDPUTl4KOuI
elhNU40/84tUjcaM1Xs/ibRisGIe2kzAk24dMyA7PeOOoK+Dt01CacjpNaxk2xig
euVM98vD49kCbBFsGxDB8/W9Xfe7+bUYEPJvrOeoYyE6CxsbWIbGHNCZnGWZjJ0+
/N1wyT819ocVKt7EPXGvpS5hVLKeWDtm0XvCqtiOrNoG1CR7oC8ooOpL1Oi+sIX2
piiqnA/UiXdliv6f+76jwIc7vyhaDjVVo3H0BVoV4pmY8TRhMEaZnVQZAXA4Vscn
CwqoWnm15+DU1H+Suu84H0vVSdSjtV6lHS8TN3cuFa61ysimLXPHnzjEEjAn8Ya5
N/MzJOLX/+yCaEcHnsQXqVBcNDoSf8pvsve8VLZUR5SW360IPZwgmDRq6fq3suUP
zyIZhT5iPbqEnGiujvAxWwW64eG6zQRyMNFI+hXhldc2gMyC4SyGHufUpUPXPWdA
K4nf/UKZ8hQmwcP5EAX3IYC8zXgn5opKr6dnh4LCOK2vdOFt4GDAkPfburXeHk5H
`protect end_protected