`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10368 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
/vEkqJfyK/81z5lf9X8oFYLgCdExARVM3sDjEKGfkr0Qb9z48nhK+5QD7ApZq5pC
Dc9Q6YRL2/hi+LwQVHXiYQrcDS6WMCoBH+2BOVI4Kw6iT4XKtsWu+QID/HJyJ13n
OXLm5vHhBpMOf832FupWLWdt0P9DL+9DV+FCTRmeg++lc+p7/0+j8A4kohpjN83V
QY9rvlJAaP4F0NoTN67/JYLCuB0AtOXLEYINrHsKd2oyriDp3jZCA9OasErbakeR
vKetHnSG+5CDWJxKfOH59LYU6ZQV+NVxcvtX7WviDCdAZlrMeYM/crLUof1jBQZd
0wlQlOuwhDsZ/IacdDkoPS61zexTAVsI7TmUuu1O6bqoJpP7wKd+7dmzfT3X1UpD
7GCk8QuYxI6qoxbMAJYLQTPFSpm0oZU+NErlxbv3124FQvXFf72QlecXVap56yka
qhGphT7NLBB30BWgeykQl9vS21A3rXyBpgWQRxCA8C7ABTpnzcLfIjGZgo5+HYwS
1nJD1VkF8DUvJo5qFLCPpzFm9oDIg6NYlTQY628pdSK2R3jtzq2P091uZgfdFC2a
lOXjmMD2JQaPbfuDneRxEFBoivHeLT/Co8N1salv1PVLY1So1EFm/vKhIeTfvFgH
vpavZn+UqKcj/v3CCjmHfqSeOz+DYQ9IItYEqNAvaQUoeTv/LGliaM1LkW0rsxBv
GTIgMs3R0smPJaQTt0v88r+OyVpiMFyFGSEOuHuvAvFLzbJsv9Zdd3XGbkAqaUp9
PK+SpWS1GXZS/GCvJaPb0cb4vP4IMPbnxeWbu+zMsDUEVsZWD7D+WTiUXRazp/gS
mgKxKfzsXylI8vdr4UzaTZWnDJYGmivWwQfyMV3RTCrC04+JQmEJzU0AoJuD1mDZ
7hIQ7im7isTaaXDsqLOgcBI6IpI5IvbrK8IZDa27fbE8pVebZH6cbLmvbd2G3D6A
mwSczyjPBAnwoOuNkiqD32aKgNrV5sUPquHC1nsILG24OZWtT7ZwJgZ5I7GWc2p2
Z/lVOPhZengY3AR+7xjxjT+BEIUg/wkp7MAwR59rJi6jp4hq4BtM1sQPFB9dzx7j
BEDeWQmP97Pu1qB6vIXuapYQBwcJjjPTq+E+tEBbnoIG3i/RK6V88w47uNtqhPkN
SSu1SNg204dpRt5+MXk6HUkg8JSLW/RmF1HxwozgIvEiIRmMsMkH1hQLH33NJHl9
BTd1f47WoNkdDjLYrTinSot194dJkZ5l4bkYzyBf4ieQYvZxU22OCtjkj/Le9bWN
xPFhWS1Hpa7JmeBtYn/hJ9QzTR+6UzKRp76/IfCY8oUP9XdqWIqPTL6re8++qyJI
PTCL3aEyAfpygYow9irwxO0PF+fsMN2lxsq/EACB+7DWhyFjZB7YYix8vKAmN6l+
4OX5n6Rv7EQNdukjpLFnbmy1OIuzklw4verQsNW31pZGUk5zDmDYkro0sjZSB9YF
QmVcmfj6aaf0BwiZbY+ih6kEApFYMJbpmCgsXik+0TJcqnzpNyLg1c4f9oCAY5Z0
YbaRlG183nQamgtrZiGt1MivklDQDF01+lG3GiYKi7PTIqacf0RJ635wQN1iXBkj
ga1xgHL1haALbAmcIV1DxTlBrdaOm1v6pem/2PjX3rGAgdu4V3n2YdWGOkTi/V/5
JvM3tWBa6oqU9kJB0OdyUd8VbumJ9QUC4Jw61p/vsek1HxH1hmH50ZEFZwkbhvoy
aqMI5CGaY4YR54fKB3l/8DW8G0r0Ukt9AcH/uOfkl044uc1PTZghZq766rsnfvBO
ZETSxJ7iuEhD2MXJfeoMz70tM5+bnxisyJ2g10TY2RNY1irikaWI+r7VATpXVhOp
2CMh6M1Uh9Qjn9DWCEksoUsz9DV7JJHQKQGzhb1PPSf1x+aMEDyWkvksumB2uzx0
bOTcnSg6hLHrziyXbcivsnoq+DHNYKG4d/PEbuuWCPxOf+jcE2EU+2t0rp8bukz2
kH8ItH6aMdRVrJNWZcjlp8UohA3aTPufwSRqSgL7DXXQpn+fhdlGOSUfoShCkFPK
MJnPzgIT60hc+i4T5baZjc+rnl34+ls1loPLPsVbInDlT90RooD5FzY3/rmQSQGO
30eRSdoR9Py/kmtuNh4gx4qv3/FF7iTa3gZokyfl3RBANV20qaX/GDEkhqt1B5XE
lnQMGfDlqVM6sQgEfSmdyk5gVqNfxi1vHJZ1VkfZ9h9j1rw1Vq275Nt/Viy+TAhy
cvWpcFtOhBy3wN0jXsB1wt58cKRHomqXiEXGKAG/y3z7rO0QY6UORJSYeS/3SBkf
FlhG51tVA95z7yoqRw0ns98BLd+PWtT7OHnI6M4v9GE0K3gWI4E/Qco6dPQfJRsh
aKIKJQtyiPtrS8PFRB9DEw2nY07HR99nudOAL8NYeLCe54G/NCCHwnyqMuUoNdcy
wZq3LDpOy0kIqHSH18tf8KJ0MiREDlLraHGcLkxKdDO6hxkaP4aWnmoPvi55PGYt
qfsfKkJqpbUEHabhimXofNGD03TcDJGPyUqbpIBy1IJFeOi4Xg+E3/8rn/etsBah
RDUPOzOZMRjlNalX6DjbFmhU2we1VyFnbu3BE7N/jCbPoIsLOlgROCggwAFR3Tfj
MUUdAEshHqXxNdBPJysV7aP7QTqwLgNEv/hw0JFiCSZcbOYufz0kkaFD70R/mM72
YTe6YYq7alWoFcovshFOFiCUMyRUnN6+l6n1mYYXQmKODnAmx1UzkesvotdMAH6T
lq9CcKioRDRv2RNl7QnLsmQpgDl5oRe0B1wYO5CegkuoO0EH36ekFFfP7t/WRfbj
BayvL3vGyb7CmTooIyMy2+NUdttye7JKpQZbk8/VtvkZWVSk7ktefZOWWaSWg9/7
8dv5wW4sa+8FOtIe4xOLa9rIIayBaE+w+jUIb6eOwWHiAyKj5bZ3IFNgVvKvxzIk
/tNThfB0aA5wE+bGjiLeeHuNvjjeD9wtiUo76FXOEvt3EyjVierDDFWvL4sCjWeB
efvy5xZBamaSC4zYTGNnbFo4Lj1V26t4g0+ceWtINvMctjR+sJ53+3ESUw2jlcRM
PIIU7sHfus43bQtWrJNW+JDOfAVBhMqCsTjM4PCz4Uo5Tkf8680UOEEQaPnWWE+O
z+uJxVc0bbTZ09e7xrcuslspQ4WkO7HSAuVqrf6GAHAqK3rog3DWasIzntoAFw+0
Wm9mlaWYCluxJEwX7Vj9x8Z2tuTCfAPDdl12mw9hDwgSyGqZvwQYxDyhGa6j6oNl
9B7X69a9riWdEGHjzyVj16Hw2bzA1nT4DndhZUaKAnko2ZWe7Rzez2NNVVEqPygO
cYsZE8Kjyq/5IgaVqVMDgU5/Z1jVLEWUsC10pvx8Nu+33GqfE6664MJiBqWVborX
lWuh5Gm4ENEzyaTPxsa7Kx8fkde+NKqyCZknKM/TwKT4CJM8K7pkbtQT75Jh7CJ0
oBkT0EbqleSCVRIvwndPHe6PPsDQR9Ws65xo68/eei4yZwAiwB4y5KU7IbtGOQhw
Jvap7k564nzQatmOyQ3vLSPB/llP3APmfQpLuEzJQLdCHe4xgNJXvi4HfwIPzJqd
QyerSieCljnNKd6+jcPFjar3QvLfBlOqBejQ5fiwW5sA/uXqsoRA0HeYKcYV134L
63j7e4/PZPfkJXp3ShkhdBtwKRYwKkzzYmtcWvUrM2EbVUw5LIUGv7v2NL4qqdgZ
b6p5tR88JkkYFJDyht8+VCnjakSYqnsMCbTf5zasyil6IxLyf0RGaLMV9eBjJp5Y
0iLrOExRVTyL+HZe1s33mrWCg/hA3tYDr2iwtxOwsyGt7utintLw9t7tCZK9cVL1
50i0+KwTdiDZdtYNoJ4NUA+N3PysGzW2Qb9+q6wi53eXj0M0J83klpAFDDOTE4nO
Gzgk8+20rSjxtUzfHAAgQWuUk8Mtma6E+wIXsXVtezqIla9YaazuZkc6oGwqcVyS
1LLBO+A7MLb49hqOJqsQIPWvI2CZ9aGOu3yV1ycjMQ+41Z6xEqSPuxtU4pEQCSPU
ZXsIBZZ9jxOVRQ8ND8ZNx2uqocDbbopPqoPQMjnKbBVKnDqbd+epWD00ODLK6V3J
OvD5yEOMyx27IBT02yVTcz5meA2p72oZjYk1o+IkmA8nS3uPGn12ZwcDIE7eVsi2
swXqo6Bd9hD+RCCDj2dpgh0FejYfWvWk7ScnC6zDFwhjsm9LPh5cbSz6HjR7HQUt
KojrvKBh4BStOMGHVf1DrM+iT/Cgya7zb0HGdR0sbO55IE9z4ZTyhuJebKlfimZy
jJUt0wPTOiZkra8FyzgakgraI4oMM/5tgbjDC5wfAfLcd9nFMBHF675Y959yLzww
VkK6zfp+RGeFhOL0PHs9UrqkjquBu1hD6Vpr8dUrGuv6bvxQiyWD+rQ57LWeMguv
4UjK+StU5x5eMwe5uzVksvFmNrnubnAaEt4pNRFHZBX9771gPWcgqWoTSsKZ1+jC
lFgPJd0ARwBM3Mwc6+UvTe52XlkO7wr3vG4ZOK7KJMpYC6n4cdUPUnpphCefsJaJ
n8xwVvRKHkxboKqajROKf0W7XAKaAW0AxW4/099mcDqrQa7geOwckDuJMp44Is7B
UvktUwZ3SkolnWN7ODB9VjIGEzff5+EXU8Z+seMg/JW5nIZwYVX+E74XnPzShKPm
rayu8b33uKvmPP+0qk40Svuxexc/4sE/YldiW1bFu/b0lmm3+MjPXAsU5cyK9p51
B20lBaTxg+yK3xLGga89yv4+2+pNjHLxUkCb+flZqkhCQExvaSvDpXeSMihhBHgU
EJPVnoI0Jjd0m1qt47UfNrUMuIBjG5k8a499hxXo/GDJbgVLc+Uu2iFGnWN/jspU
cJ653yKUPHkdmC5e7mM7+V3CDJ6tkDCzd9u8k00DJno9r2nVJl/QqShn/8avdjJR
ZlAtXVXvau6t0/CuzWkmNtB7qk17cGxnkX8KqZBRDY/8KqI/FRs56dh2dFTAEZSx
Du0PxbTjE5OhwvrWYurKa++Aaw7xTR13+T+RxzhkGPrp8zJFad4gUstEzEpdONtm
HoBago8GDJujQOclSVt3IqFVfs1kGs7OraL4nmVnAqqPFH4IeuklKmLvN0ekSfsf
q5esjT8DFAYsUZhYqrzwZlqp/8ECfHDqwa4pzmeNbmRGEvgfxhAnXpD7zR/X/jDe
YYq2Wn+9fiexDTUlDP0B3zXARDykftVQ8RtzUl4Bxv8h7xUyWYhNxinsy7R0eqnF
sYrIWmSpjmPKSpJqY697nC6POy7uCtxBL71tfvpaBnigwK7MYDIU96MyAbtT7+0d
3Pfz9bgf5WlXZxwfIZafnpyhIYJxxANLbpv3hf7jAQ3HBYAyiuBOZog8ve/FCfgE
DGSAnkHrmk3XeeP6ufXQtH+DdWwE5m8BqTbY811iu8PALUhPBM9rxjNESitAJslA
Y+W4A87VpgP0/7B/UcSc8rgtfZubycqT6jKmLk3108iBMsh33E5YOOb83RwPTloy
kOq3xSFI3Cm9+QSaZo63vA451ZYry307oNqEe4k7Q6mUv1IQADuLcuefgjIyQNw6
tH1TD4EtbTABjSRJ+qUvXJpSLgehtld+t6Dl22nmFVsmadhB5BkQGlUNfTX/uCcu
VSsHSCeLfE67qi68xObA6dpQ2b6nYm23kPAAFe7+VN5kh7Han1xNblwHZ48F4Kj2
T1xDOn/RFS7wsHTklfzn7ylVb902WA1pPfaRHUoVVLL0CWKFz2dG+77zlH6n1dHT
iV/e7mvcUhLCpag4w9JGhxH4QFBnkUWYsSwpRlaN0GI227KC5u/Qe6kwfIJL8aL6
sjfiO83GMKXBo68T98Us6yJEDm6WQW6nGdljfYtgur458TxfjjBqepNSRlPhEhuU
t1exiAVZv3Ia/aL7n2D5rdhQC/c0G+uwDpKDGcmKc+woeF03nIuwaViXimqDM3Nb
1YBrWgoavC1+tr0qJvlgKcgpjGAZ6WSUxMjmGg8iyck74lLJc8MUgqFNKr2ZY88u
Urhv1sAcvAFdHkX4Rw7GYFIigsxwbnHNWmrgc5jrlXwalKZiUReTbzDYJhg19OCT
cO/RE1hH3k38C7iCF19yVOHoGdcbb1JBx0xlDbdRofy/gKh9zHgyLm0Bd5rlEO3d
4VnS9LXuiVIYuMXuuEQP56Evkx8v7Qv+ElXJi7J9OFhW5jNWbfUxlwRt6yWoSxiK
2UdG11ZXkvZtnk7OadgQp76E4rzjKcKzmJkfDqFSS8P6FuNgDjXrugrlQ0wc5k9e
B2WR31IZdpiWZghTTnnVo3Te80TIJPjItyCr+RyuA0KkYI/LAKdZsUEySF+giKq4
X+/tkbtcT2C4GmjKPea7FlY3M3wRrPjDLB95/Kg/xXy6Yi+xqhocbLv2USeX2zoe
ruYasTNOO0+VaiBVK7abHVQTfN5GpgmPDlpR4JROTFdXSghub8EoCII2UzwSEfHV
iufZg7IPVgHH0bFAbkc4OydflXrR3Zu+80eFcnfQzOKxYKnW8S5ZMtCRsVgwm5Mt
mSMUjJax+Dp1FP+466dAN3dwREnfVTGflvUXLw0a4oMkPdQPYIFAwAtdF9fp2EqY
jgF6fODZstOsY5PGaxclIuF9MUAXk3+UjCgSys9uaUga2JVtmb1TMr5+gwxEITJP
OkQ3DR5O7u1G/0QSXINoUoiAonFvh1rureWa7Ivgg+HlFll4xjG1xNMAdTNhTmYk
c7UlObW7OdHEvq2IonvJVG4hW3FDtUBAQ0khdaA4uzpCy/q3bzGbIaBSBL2GzRjH
qBGBEn1BUXnX5xOZouFOM2jIVL2LFzZD51zyIvCBIXQdUF1k/rxdO1maCb8PbCIu
nGqh86sVnXIgm4WgoN3igDCqbDki/nZh6aJ/2/cERsqoUNKjJVQ7kZZs29YX+nuM
lFpodl7vB4lSqUD8y3pdfa2Qpoqhx2Up73NSuXIfFaABSdECILe095RWC7Pb1Is5
wZNIHPoQO1Vecs+lP0eGYatYoJbK50o5BscaEK6PHp3EB847gS4+s10MyahgS5HB
S+uc2DUbjLHOXGQu1a11Xw4up+ny4VATqcThbSio09wq8x8e26eNlpIrvIUHxFq4
iXnUymMBn/DDca0GRn2ee7VFg/NZazzl6dylemYfKG71Y6Z//YGV3BznHtn2R29a
f198mRkX2mgTApYuMOCTmAdJ5fV6IQuZFH1J6AAaAmJLAVRKZc2ahSVZFU35h7aL
ZHCj6sUFlgWYtfqY1Iocsbq+F+9XsBsEnDc+bYsr9uK4IqmifSdecKph+5XMhCqc
ZwJW9uw55XDoBllmR6f2i/h6bkN+oCWpk61hJu95APDpzfgjFSVnIeMgWdprfs6g
O4AQ8Lji2YMReH68z9mTvQD7ICFWxyMht8U6OYQL6cPpkmxlEFrPoCsRzsS6Upx3
Bfh4RdL+nyRcKvBjfev4Dx+HRCIc0GV5ogBj+QCBikE3gQmutbGkPRoVTJKdrveh
sQlcC6PlsXeI17MFiJGV8mykTKah4roAXlYQClGJZjWAfEOUxg64iWGAKhD8yCld
Zpx8XAL7PDMPqG7oCaer2Z59AQ/Tfrnp6kHmhr15snco3QQhyIF9J5/NqNLJAKiR
S2b0dwb0ZiXuO6cdlVaNk+hCTp2omtWqAgkhcjxWzOEu8tregJR242r/3DucNpKo
Lspd4+JRNOGrVhkJsYY2mWCm7A2vtW6jUyc2EBEmlTBxtmuajP3xIBmsivclDRlY
RBcLaO6CnrZTMJI20cgAO3H1I0tcUlEwwswn6E2ULQOOp0+eyeXKpXMu5ZDL/NcS
Wqe3c2jc1VXJIkdfGsN8AhqoIQYIbEdCrgBYOdbsoYk3qTLvJzNWf6Sy4ovELKRS
PFaQdhjRbjTbKZjEu8O7ioG7XEUEVKIA2jpavx9tIGrasds92X2kiyerJ4eolClN
shkvyU0sXPsMj0VK2+1+njqHJa2JOy8+J6Rg6vw21tVHKlhNLsA0yFUXSfuuSc3e
hK0peyxiK43ZX3u6KTT3MeYDkE0soTzQRw5Kd4qKYcxt5eFp7FRkxEpW2ivCQABJ
iL/XbuvMTvscNG8iCi2vEZ+5zSDBc4Z+3/LNscpJPK6rAZzYmCEEGi76OoKfFRPd
itByTS8o2keLcZPPlpmp+1jR+VwlkrI2tPhkiKhOO/3IqkZdJAMxe5tXcf+Iu93P
HWfP2m2zRKWKlF5zYkvT7TiE1aj9eyC89gdGnf6CrjUbge8mBnIIb0b7ttz/sJO4
d6JwGVzTnuH/vaK2uL42uJ9q5uxcuxzj094CfVWD8zpZFCRwmOjebeQbmMpiHG0f
EZhgxYqUrnIqWdQYfClK2KRSFXIMUQwLrSxLuC00ihRjEtelMHKIKXbM+5Vg+Iz4
hGvqmI2fSiYnmdHTTjCiAhwjrxItEFLoQ34Qe/DBs1p3GpqPr1rXFgiAfrs62fn3
d7kmuaCS2SuQ1ibVLcMxom6cDskopwY4k7yCmb8qdDkU1P+N4R3mnq2nwbpnVCIr
wBjQ5/fgrbvMvwXgX6TtEWltqYQkmb1dC/ekH7Pkj7cX3zMjShJzo3JJ3LZt6Z+Q
PZXEWvgaPL2ZpEvFET9W6FRwNoL1Ctynr+1aCif9VVFqRKqTcix5lA1qU9tFR6cJ
m+fykCtLhoMXw2vtIs2LUHtaL7dIXI1rbhjnQoiAHUp6MWKSg4dJWTP9trPQAtQI
dyF8dtrS5uyI4sGJUx/jc1XKBil6IgIRecxEumfrnZRaW+IS3eq7n2lZF2T127aD
WzMyDDTeVKNj7n2ccv54tJk9FybeqTqqlzu4YHONPjp5hDWi+EDNgOBlA0LH82pL
QxTgOxkIgSJ4t+/QuAeRCklpBl9luR3MGczC0IxvVMlPIF9DLwale62X6kelxTIH
5Od1gmldO9bf6/0X5EiHv0ChoAWf03YSJFZgXERrHFbIgSN7UoWLvm9xokoQ/AAg
Jx282fHloCGTzOtXGScxKvkzU8j7YCrPxIAqoxmOHvqDT+Jm9aotm06RKA4iZA8t
Hh4oz1XIMrWaHFy3fccEodNNStmKbQ/ycQL5AYkHUBq8x/Te1hy+GvJrlCHeoZc0
uXQIInsKKgSHFMzzbkAHnT1fkoo3oMFX2yWs7efoyRtistvjn7Pf/99t98Q7+vDH
6yTOvXBJd+YdIU5Cpq7srB9ym7CpvAvhXVjdVN347YW8g/flzQEg0hWkxiy/1J14
h0h68P9Ct0hHsacNOXoXFJ+VARXNZ9mOlzV5WgKEi8XSqva36iFB+wW9cthnglAA
P0jceU+LAUKDQgXMhMB+Xr8Mn5vzKyuQehlhxDIrUd4YqigQkxiX+a0d6iMEKO0t
2AiiRRBVYH0oUmBLJLdvyEVX7in0erQNrqhBHSSYyLZD4GPmlDk8fpWVZFXVIGVI
JA2yZRSju4XABdlSkQJFKM9fvZ/w3aZEEPnpaex9CKu08woB4YzRHaYHzgaAL2FF
r4fHb8QDYwPDSJPK8dcXaBY/YokJU4nq7v/NBue5WzFUt0tU4wstM2YwJ2R4kKPE
EtjN3aHg6MG6nqDcUhAkiJk1lN70DSoCl2DYPbJUCwu/lT85V+Y0sZxS7h6SHYee
h2GvaeF9b+NzaViTKZmV/Pt1bIfLE/SGYx7faLJjCNiotX2cy/a93sfMQcD4G40b
bDxqmbgqwVYX8f+ELf/SNMIqn2h3JMHtD7bFJoziSwASBHHbjb/lW8LFHh1lQRvI
fz4vTBUaNaLk0ntgtagaVI+0j/vu+eoCg30d0ED+/BhzY94gggp0bI07k7eQFGDG
DWr3Fx3GAog71ALZ2KiALJ0NDjQYzC92i+Nyn5lUwGKy0bL6bARB6qRXzemEGNt9
UIlAG+vE9QDCQGfFJH45Laaap5Wf/l6mgEnQ/GtRgn1zgY8PTVTG91Yi+2tuXQxH
KNNsodL7hT0DL1glIEffTGKAMwWXU8OVBhbL8egAp0yni5x2fJmoDJ4iFuRxeFKa
gzenNzpONDp6d4ow3osn+t6ZZz9s708znlf5owz+K23Rm/JyHv8fQ3JypcByqJUy
dPbztojRioebm0cIdnA/xk4wy0AO3YoAQYgYtXw0P0n82ssAcjqrEXq+6DaXZrxN
L9rsp3mC44I7VjK0vj+WhRyZF48NaAVp8S2Yf/71ciyUyxMHPWuqLCMouVEkV6g9
n/UBFutq/hfcqM9h2Y5qRl6QTasFSy8FZrDZnP4jM1hxT/JQdkgnSzpa6DPL5Ogq
i78wTVb3RtGhVNoddkVrWD3xhKTJdAnBAlobIlX1tUf2TmFe4qdUcMkH+MprEj4E
tRd9/CtkpLnqronggbBYIsP7tGqKi5DtalBj0K4MIMuL5SJW5NgpYFsjyTQpftHH
4446IQBbBqMRF6Zeld0FccAs/xUxTdwp7F+2/RAeOKldfCvqynWmfSLIxMqkSbeJ
ThfxZcVkKqwzi3RnujRVfZOOl+tqhRBe6OoLRlGONTKyb95EvBb1gRmo0nUG+MJY
BqRiSmxJVCK3QVy/qq1OfEaWT0Q49s9DYf2QmyA3mXhTtAV9TVFHYzPMke2Mfn9d
N7urIOePAVTi+K3Pqzg8cbhpA2ViKh4Sudj8GTKIT7kJ7bMR+UpoCH+X/zttGENF
Fgw8lxuMufNnTfRZa3hc7zU1lDJvkoTnAp3qRwhDnYhTmyd6pMOfqzVrIgqCHhKM
7HNUMH8G1SWxbGCJoTbSD74nW7VCSPL3LU5sDki3qe+IeyCIlHZ19FWOUuLQtTGX
OneULPkioTBIBbBassAeXIdAEouIVCCehe24ASAvGLH1qzxIPv4G76Ovug9SK/AI
X47+IStUN9oFmMEcBePI3N+t2MDWH0mVuDVwVqCMqRPJMPsKHW/HDdNWTqXD3wO+
xSksMUllEglAMVgWFMZX3eU3yER4Mt6BcDSy1DASf37gm8yzXKnq+QYr0tKPt1bz
p8XOFSJEz6yLcfHkmDlvahbh/S8fu27oSa5MgWOgaUPmpTgH0gtdOtOKDRWQqcBf
tlAEgh6ZwwO5KrmrfQARgMcxlSepWK61ztDWp+rDPWp6niCg65Ubj1CW9k9nlkAw
uNLdt/7g2dI2gCj8yfkyqaYi2dWaiU0xtsOn626RmbLVQOqNV7fpvpbISuoVsmH2
Rnk2YcITKzpn5YB0aFVQqb2AFqdpztuq6c/PIlzLeO/TkCoTxJC9Qoopccr2eCZH
Ut0SDlUshmCehi434IRyMVNbhSkwqdAgrIyWc9JJS5YAtYHoJdcJyT9DhqZTi18X
AzzJwZ38h+iRizyCVF1GZsBQ2mSq/YdCi/am8JWv+SohAl3UPJMOVlHFVOPjOWXO
3nyn8kNnLKazPUjMJHxu5zSWpgUGVggd/fMA2+cNAK7A20gkltWkqWksXOn5FARA
HfI/Svpf34YLLknhZz7KXF+ABAnnEBvSVt6Rr15Mx34jbD+iH2Yfn3wD/TvIutqN
VpD3kXfco8bHirPOg+N0ZRtNP5oZkvWCzD81tjudglIfFBeZw4mHkBJQf9rSOE/i
AF4Y30b9GlBIX2BLhPhwpfJr5D3Rot5x1yxZ50GQ8R13gg3VhEwDps8ysUpwQnrU
mOSYxS1q2luVMD9gVbWDyJt7vv8spk8X3dgkyHZicMqbYGWA6qH0hInGZEv71EWr
MW0bmB1m9JSH0VOJyxUbfQ/BgcFNFbilWkp1PxjxYJ5wy4nwAYLbYaNGHhPR9Yaz
CUULlkY2+k+HbE1U9L6Ab6nOx7XegXGjOtAuUfPhW07eJK6864zD19xrcqAJIXlU
1HW8XeuZp7XSWtpkgJ+Pp7I2KlLAYwTxstNFeIQIE8uid3KCFe7yLekMAoceo8uT
r0OvBAFqWERvP+7zITbPr+kJ8VhajJAE8fc8elGeVhf9ttKLU0vO5Jd1w3sJJ21A
+syXB03EfnjPv4Tg23UPuuchIwJ2Dh4pq4GK6s2x9oA+26fPXczJfu6przmt+H9m
DHIjcqsN+iZ1S5Ve+MYHGTCSIFhu7AyboD4mZ5Xz90DrGSnKh0cp4JtUF++SeKKG
iYt/VcurOS1qW5V473MKBm5pVMOv3RLpa/3vt3h89AlPBNjfi5dbtFgA6nxacu/h
QehNpFr5FLkZR6Zdj2UPGoUenCQlayP7PaDg4FosigJnmYK58r8rcgV7mWL1tXz/
sqQ1XIqucaLOCUFcriyAlOhjE3u8rVEYh/rMA7mWxMTw8Iwm2WdfvRKbUrOgLmCw
6alG/urhFeCoHyTybpt+Mtf93PWNLV9rMFFf6Qz6OUDNUwWIbPaTKvpPu9GlvC6p
UJKPE5qLt5sIQ3n/go8ufGESBARvDWGvsfnMSsLVlt4rvUzTeuDb1AR0R9dk3BPX
ZbqXeusvO7SlNJbT5HipxPcYi/UpKi0Ip/DN7J9mZrJvkNJKXF1yVmfr8f/BwcIk
EquKBepyNGd+BMTnQ7Ha8Zpz6Dmi3c3kn7JFxhIu20s2kgzZ7EPmzcpHvdyHdpHz
xzvRFq72pLAza3d5UQqrc8rYWOL7nqqGpQZ+7C+pB3JbhzWfv/xiIi3HTynC5pIC
+hcww5XDnXmppNjd2jx4tqjGkUWLas2/sXuFJJtdwtjl5jPOddeIkSdke5cd7hQt
eVzsiSuMHQLR9nYNBvhBTOxQwMqATF3Ok4XGqKgoeOap3WDYjhtgy5hhnlfJSCdr
7NtRJsxzE071VzE1PBWhkrGY/jmtp4GmLoXAO0eCJq69HZHAHVndFWcpaYaTvjrW
SDxsaSRUPXH6wh3NntygwRCOLFbiN+aLDJaX67xnOdFooBB5BkewV9jeHw19DMAk
kGirmnCdwMqoqFxYq0uLyPCQ+wWgsb4HdhfNk/JW/fxo3TDMGMMNdqFqrMaZCKL/
ij44v7nGCBb8tIiIsnUBcKlCzVu415gJ57g3h3rTtnnw+UPYF0tcpZr+83nw13Tf
BhUauXOTGkO9tO5wK8MgFMN8AYYKiJ2AsDbbVx4Pbjb/gCY0dZp6bXcGpGVlnozZ
FNZC/LT6ZozFFdTs+qYrqRr4HJx3G4Hwei4RlCXTw6CtXiiY7xWdgb33t5CXwNCC
ESWfkunBTe37rbZjTFykhdyxN250RtW6YtvUaANuw+26kF+MAWgxuZeySzuTGBRk
K4SOVKn5qw96k/uesnNCofXnC5t3670dzfLRBzCf57qUvbuH6ajpOm7qg9VCpTbZ
iEJbMWayeOCJ3NcGK3MZ64bqv11C1xzdMQRWp+/dC1J7ze88JuQPm+JB0OZE02Tx
qijXm3dT6Q2t6999MD2123x++ilGpVdemea9TV5JZ/RBFLtocsOIBM6BX1B8lCZE
v6SSoQnMVg/aYGTPlOwTyJdxy8pLefU8nPnYO3s1sa7iD70x+z+7AF7lvwK3vh12
4jPnEdx1519shIQyemhgfIZRjz8y3+u+NmI/Z2GPClx/pbx/bEuWCEzMkk/uy26+
bKZnO99cRt44UVs75lCeSo3sF2SniK064DUd24jISFAUNr49q1/JFZYzlhTgKdhp
92WCo6Ypwz5IDoerOVeKr5egiDhnUJN/WL8qSIre0WCycmq60gUe+ldmoX7m8mNT
Lsfl06NkWVeUlqByUn9TEbUCscOOyOB+ZYWA6OibII8JLK4G9MDFYKQAf8Qp74qo
sj4alYC1amAjCFlHuzoSk+nYLMwtceJIwdpeaiK0nybWLURgKkGCWt3ByGyeZwHk
`protect end_protected