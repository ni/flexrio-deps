`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4320 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
DBGZtUPdvgnvgIFp6VMrQUbT2iVccnzIQAUsmPwq1L14oYQRu7Dq2OpzAkVn70zx
JrW0jsyikefqZuD7EGGVOYFccwH0FTWIX4hF0/3GFfGZb1jkO/mnyIM45cRNYVKA
xo5My4fM0vOalzN7ltZzFOiQRLF8RlFVe2JxQvgd2umAgDsh+69UL0fcO6B/sfaD
Fx0OxPvgP6DmnIZAf8xuIt90nkCnT+dEtSu/tR1VLF5J7UoTAV70mu1IqoTD9K4l
/Me9Rni3x1sQ4AoCLQ6qWSz0pRhC1cod+bFlQ9158WhHFwIz/TnE5ZmWyfv6hzr8
zKKrmeys5vbbhQPMqobB9hyqcA9wf7Zn0ULKwQuQr4hTmg+ZxdRb39n/G7RBhNef
04ZQIFAYmFO10R5L1qDFbplZNN+hiiByU8V5m72dt7DWzKqtYMWjhdDQMwMrwFbm
pADB21rp76LMBSAGUQmAr+sV4iYFg5JPVPtJaB0923f6Mqhg+FZXniH98KaG45hK
ld4uHr8261bjHX1PybGHAzlIYotboY+3Za9sKulswTqUOxQIm5ssi5ZrUvJBSzf7
wWQNEpC5IYdfHzJAQ1TU/qqTW6nOmbnsdWvp3d333bMG7ATy0cgL6rm606MD2F82
qXPnRMNdRx3qli56lu06gKG0juUG9m4wxAye73cicahTJdQaMsamayk2JZdazvBI
Kh35P9VXkMYMMoxBAdiDwvNIdHern2zkYsHuOjETCvw9Zhr01b9jwDQYIQZr43Dk
WeYZQhofH2yGlORdtk9HQ0dnhc1pTGkGVOc3WqK61mjJNVq9UZyaXdc0/Pd6655z
CoF/KaqkqK2+b+a3nd2KXfNX3Go2L2+Bq1LKEU0SUcb0YSFmB8UbI0vxvys6L3PG
FwFNKpAmo5EuE3SsRAiPimd5qCDLl4hneeB4XSsgcvaXILT64gNJwtc1MuLmHdWz
fVXO520+0Vmi7jxguWp9XAUwL4fjhwUN2SXoHMbmHClvXHsIGCBUOhdO4bOcz3GE
WwIDAIOrHAepXRjWZW33xYpffBuX/6r0CUJCCyVsLp/oTJDixZ/0sxxVYH5xn/7B
kxedQYsTUC96Oq398te7brgZN9IgR8QHCjMHLvMJgSI3TFLRkL42w7ZaRnw8Rs6N
1ckasVNckq4ewcU5nIdDtnLBrPGqvTfn2zwwxaz/CY6g0tkcpuWgefSNETDziXTk
C0Ql6r5R3hps6ILjolQ9QtsIB2SSKl8zOdbNmBj6W2jGSOlKx2m4n3eHXN8cMEZZ
nD6M+yUFnncssL2oNEr/d0wXFkgDISnvseNls0vcI/T7Y8ixrDlXiYZSiJuJXty1
3ahR517gpT80kuQskKAKo9x+X98GlLXQAS677xoLTeSxsAsNfpjgB4WMntEfsWya
CcnU4DFTUE5JXI1xkRLgCnJfZKAeZ1jSTqQ8XAHk6Edply89raIkVRVRRbpB1xDF
nt2Yf46X+ETo19fSk04n4fYkLgrOfnT2W/B/A3Xg6zEh/MjmluWugjzlFWYQhA46
DNK5w9KTmq2AopYiz/uskEBd5d2R6BZ30G/oda8pQ20qwISE3sTTdVte1zDuTLOK
3VGSTtgFHRn7EKrhrrfaWby0Kfwz+vcCfP5W1DGPXyBBdcayeiLVdEnpE1WOuVnY
OYOLsHzhisrf6pzphQ67vV+IQ40n9EsQJAhW9TPPpVLKWxFCTxfN5FoObyk1egIt
OwpuiId5FWI1Xkr7FGpDt8OXrBP+DFwvmELYtEeUNg1eqKBOeBw7emkqhTbZxbIL
XKCXYUp+CGz81W0r6TWidECGR7Te1vs9+vv0UJPaUosw2yNo8sq6ueHcPDpBNQDJ
nwvpTfHuj/n2AISv5ki5K0NsRdac6ZSDN51gTNPzb295dhdii7C3IlkiKVShzzIQ
cMF2WqVwtdsP/ld11WXnXR5vMEERWvI2h7APckwokPjAigiK/dmUonhb62lpfsti
fxgbVlVg/rsM4x9RnJShzCSacCLSdTGr0vatYGZKC8VlhdvqF2/lZ1CG7vLaynrd
sdUYMzs4OxHmHW1uvo6vJgvwnfTWxDQ4aEMPcdA0Ja3SDlJiQTRzO5GFqIqYkgnG
9sYy40QQdWQNEJW73ESb6p4QQTsL7O4xXZaQhs6paQqcX5e+OKVTWC/6bT9+4XDr
E35Xpc66IJronHyzEKy+zH26pzDQNUt2xzO/su6hS8Jq3MpLduRhWU1wAoxRZNUd
nKn4Fx8MjwpgR7pFeCOfSwOEEd0rPfrtHwDhJPQlh9sqjHuFI2nhK0fzOsOEgxFx
Ps9mWC3KvRWHwNFvzN3Q62MY96YO6yrfbwcWCGGjIK4IVhy1no06GhGqt4Rs1Q20
C+4KAhBt1zTPxM0Vq/bWzr5iv6PPz20lD9O49ByUWUCh9DsTglLoNlIqREut7CD5
h8hRVQoVobyKhI+Iw18NlYnNkKiUPP38uTmUByQ1BLs3orWK7TKoIuocgIDiUc/4
gdKWjv0zcQsu+gV2tIls1B1MRTb6vYHVznPJmFJtArtixzE/WvE9ZacBRN1PQNHm
2OZwZphbFaraJxKiuhUYMLpldg/eVr8B/fCDCMeOiUlbk67bJzpo2t7YS37v3Zvp
UCeGMpjolhu1ic+rHS3ICiE+xtpMw8uSSjbFlgOha3VY1JB8Ts+PwPYkgqoKIP5X
wdTYAv5uH+0239h6xoeLZtcoGorDH8xfzIBN85KYgAHFe+TuZIJGPjXJAmx4PGVU
sKMhhaDWmt94gTvaWL4+HWHP8vvcT3ngJoftcPzqs2QwAnVsyQw3pNJL9+Ki9jJN
aeKdlLIBKyoPcnY4tnunikAl0rRBb/yQUavQuIRhfy6h6JgNtGeb2EvQFwNPSnNI
QLSNzE8vNhw92dj0XAjOnwR6SENzpnnd219NioBO3V0V5H5oG5mS3dFj84WiP1A8
79ziavHCr6cE+c8WT+s6Qw7sMRHP7uDwUx8AFwGUj4EbcjkV/Sh/t1FzeaXB8Dlo
5IeZ8LN4LuuZZh7Zr+nLVuLJc5N6yPvjwE29Z6pB8oZoktXkrm05wMQZmpgn+oSf
REYty8lcyndRbesapuCWZH3IZKr6fn5REFxuhxm/8h2UV1nJluUTnsNlslbYF3jV
0hcaOLbqpbuIIagQlZLLhs1Kj0sEWqUEJykZcRhn6qdBvNYarDV6ilMVol1gMiCE
ZYb2pRec7aEQTdAccCpqA0MPUV1zICxYet7mPU8VsjXofuegED1n6W613taXB0NB
WnRlxX1FI5FQKo0oRqpXq1VrDMGeU+hAHRqWlprLVaM3g/ypdL5zzzVa694drDyI
YeuAz3+PQdlsI/RyBKXsrvFd5lrykBMKIL72gSsorBsZMx54ruRhjPln1X5VEDl9
j6tBVUc9XLEiL+L5bct9X8BUdMvuChwUCeiW1hmIYI0ZVF6yLIyPxBNY83uyOORx
35YLJTfl18zw6mqVCbKA0CzEmyMO/EREPOGNej+L1klTmx4Vfy9V/PCSa0qiaZtH
wQ6vKH4ae20aOQxr3HeL5ulS84CJ4+hHIAqi6YHr61TeuzU51Iqcf0mNO98S9vdv
al3/Z3C07ARM1ehib6TDvdcVSZkxAyGQqpcGr9DnJxDE15VcUakGK1IzI8sxzETY
EzbvoEGQcWz1HsIAHuJQlrdOqupJC72dwU+Rm8ZgogNJHOrev1v61KjJWw8Npoak
/vbFwWA9LqlMH8tj74kIjtsFZJCcdVOZT1P4bVz3ce9ScwPvTdXHzBrazG/0287r
ghxWEQguy+8KaHRIwAB216i+xO5bquMayrA4cSll5AXTTA/j7IQSX1yefDPiWgFF
mn9/7RS9P+n2jV7ezELAGc4yTdAqHnv0d0AUfqnvavwhhLEJ+8cwBD/1VuTpqXsb
w0C2ae8O3lEBV2czdXHxstQX/JDxaMk8qryxMMMifxlTM4HzYLkOgN+FSIpc0Oyo
z7/YuN1A2gvuwlHweQDM93sD7jWUipQ6b+DuLL8dpqkfPZOOEZz00gAf2vF4//Cp
VPF2fEYNzkDMllt/ztY1Mwye3TlRwZ4n4UKBboU+KGbOonqaOGdGNTqYmIOu1Lrk
P3o73WjpXU/S80o41GDKr3UFQ6ZifQrhcgT+72pSJVv4v/jY/CZ1JXQJE1veFH2l
jeSHlM13xEOgA8ZZRDwu9RMg7bGhCHMnsHJDieQXGzqTL2Ff3RmcliEnrMPQpvEr
jHbvEHvT30GLNuggyUqOoJRiaoFBMbVTFyCn4AY9+OKJF1KPizK4kLZY86moqcVe
ev0QUFykv7S94uHhci8m6pAOexe1fvV/24dcmqsyfsnSaeFjociyf8/xh+6d74Tc
IG7WBmd5Xtp4seN+yRYJu8pNrwOEO53mAWH3MElfVRrOtOVAqYycM0W7LQtPuy5Q
HH4ooLNVcvGNnpsewsNTLW7wX+Xu8hc/uZkiHDmZeFytdc+kEAPHzXjTo/AS+lIY
dHX8cvyRL3CgwmH0pwAUdsOqSXe3xlZD9sDQb61qm+tdYp1dqLZKT/YjCMXMyNqn
pqo3slv4dcli3Rzw/Rdp16gkOD6otwvewTk0/OAv1mnL6srLXGjRlQhsf+uPQ/GH
QlTQtjMbCxyga4SQa+E8xc2XHeuCmVExxar+gu/ykb/o5Sc0rroGHcGB42cImE30
iFv/C2FRLIFCE/HTZLiqkFN14PJdBRaAFjepdudqQi0URN1CdtIrp5N8YxW5Y3ay
I2nDfAzFmTnCH0/nRr/L6RcY5lskdEC2D4E2Qhmf7Bnat3v0Ew6GWZZK/7xAE9Nq
HU6SAzlPcBivt2jWJSSjSUNhXUXRjXhewJqkfhUz+rVHWS9CGUlAkPUeK4iA4CKF
wTtjV42b5ThUIfL/Wwry2ctDFbgf3PXfQgYvk0/QRG6eJGzHheyvpceW/xJ6y1we
jZrbz8lZFXjrOAudzYUr94rul3Q34eJgchl1WmyHz79QkCKZessdKdcBex7aiS/T
huHHtURq4mQZHX8aRB5RKdMv8lTJkm56V99ULW3qroaAYOKoL7JtXU+GZ/bFf2pt
wdF4tV8FxrI5oZn2eJfI1Gqo/t3d+ekJD3RmqO31CtBWIBYvML8JGqXNgIr9SfxI
T5WtPCBoubBP5E9yhEAzLFc83RwplpJxSj8W4zTFIbjIAqdu3zOMcnsm3M6GB/Af
xUXvUg/7R5PVSx+Jh/dfBqfHer1+o93nXvq3DnhRjO5bwJpblE12JIAg6lpT3rAa
IeYGs5v0ramLfXpSEISpgmeXg0dj/giYaKgPucvKiILrQWnelcuuD0c5hgi9D70V
jbsu3doOpeoa47kw3sr44RtW2TyS91CYmUZHGrKexvx7b7JlRx+nNxZY1aXI/sTs
0UJ59U3gOsTQFlUuKZaK66Fq3PBm/EshLUlXwhdKObAqYrVG017lpin7jZZoQ1ks
OK9Trub9akZiGGCIYOR+ysPXRLwo0eM2soUqf4LwGjBcPVM+WpLwyWOXFTpzYgcS
sKNAFPHPBbhsaaBhj+RZuhfatqQggiFd0peUAY5Mp43Zer6Rvbm/ZBxUN03cwzZt
Kjm0wJffBo6F2iyg92yQ26WeBU7KgJuTVv6wD6HzUTwH8kxfisJw3a/2KQd19EJJ
`protect end_protected