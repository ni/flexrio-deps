`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8672 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
ZIICkMu+S2rq/yOQyqhpunPPNi/HmLul1fW54vDF71teqW7ZJs6XK4hCi+yFf0lk
aUhqruIeOrc+uDta78fa2OD4DOiuXW5mWrmGivILoowKigN6pkH9EcDYWYO25H7G
Eunp6lOaBSKFT7UYZYkAc9n7XY19CVTyHJbunKdYb0U/MIvJPkuX1YBLPxqMk0aN
8OpRfBaCGxMuXqh/piqZtK20FUPXaz5DNVe7NEzLdeJe12PlynbK6XWnE7XPDYJF
gnqrL0ua17IzYiR0oTr9MUnJd1YDXRoY2V7Ybz4o8Iz96p/4lq+/8WXYUFKtUZck
2GAOERcUYT5SVwy6qoA3BsFhSMNSwIAGZO6tbj+KmmGyJ5S+p+X/t5Hg0i5DUeQu
DZ3/jhmsrRwedEBwGkmga3nkw6JZg61KmQpuy1zRhDOwnt2WOXGUgnkP/uHX2bc4
IyK/VrYDsRXNXH6ItySyZwTbK9BAQrjLtZtb1FSPPre1KrTEd1MOeHZKKMOOv5Nj
f5mcjexa6kUMrbTdByo8HaHQCB5a38AWulRE9msJ1UZitHj/AvS13MMrxRehCZbP
9MVqUUfvGXgQavLvFzP78X+cNoEk4qWRaE+OwtBhpGgoVU2cOY9uMv9UQ0t3jr+5
lRX49xm3/QZPdAEqOaTb9vrUClSFxOQyZTsV3rxyQBNMo3jmYxNq0U+VdSSw9GWa
QTcnhequgYqT3+HP3zR/J6bHYO1+fj7TbpvSPkFuBu9shJt09SVjHoLCWkQB0M51
OTpBxKluDsen1JmhoOsnjZL6dYygTVVCr5bRa2ZGmGjc78GAV3w/+Lwx7oiJnjjp
zvCxU2LpycCOY7y41nyJYiK565g5VrM0ZBphGzavptqLRnTnyy2IuVog0vpzVJ9A
99k8BX/LJ6iN2pOpSJAozWpN+h7gETTS/BaFMOSPHH63U2x9RffJve50p+3Prq6f
EvgEjB3+qFY34MzOtvNLEx/u8s8B+sTV6MR1GBB+gKRsTshwf5PvXh15j7zcGCGV
1VcIiXiDQH/R9tHfClhSclGNFT84bTznrwcyx6pw/mDIHKGLYoez5ViyDvIpX1IK
Fah4w/5Usdx/7CcIBgCzaRzxBh1Uzyn6b9NZVCp4slwWpUa3tltqdzHv3HmWNFIp
Ls9g5ChKqsqo8KFjQSxWuI5lUFm/cWS4oFv+3is+84JRMm+ENnJebZkAYUvcZNo1
3K65kPxm2wtdde67Gz1SRvr8dmOQ59QeYgTTpwP5LlayYOVY2KbRC/kvCnLeo9rE
l5qqj0W89us0vxFdRLwjXHO+iKrQZz1v5+5KPkCVUR8kYM+IPnN7yDqO5mh3xB0n
+a482QxZbNx0ujcArrmWsNvcXwV5EsV6+IGJA7Boquo67l8uILCLbq+J2eVvafZG
mw9uc9Vlfi/wxkm4/NnaIYaNHSCWVJGhqoEorBOJWDg5oLJx8wsTr4RzUy/51eCj
tdka7/+11zn8edCFGCwnTnzmXF5CEUJzN5Yme7Kn86hekuxMZPlYIwqpkzr467JZ
hl4Lj3bCGEM8LDixn3rdzSnBR6DtTtYdknT1JwEbOO42H9flNMjWQ3M/hFCKi67C
KV0sZTEyb2h2OgfnTjivZskT4UXiu3dRtmFwxSpl14EvAr8FSSVzR1YEQ6ETD/kZ
WTfHKA+RNnVg70IpGRKJdOiCqv46OMJ/sPToyStOfzJx30BVs5iDwXpCeuJ7u3rj
SxflfDUCaxRegdwi0zr44L2hDKQBkk+GRBoqpVq9s80uInP7Gm8xWcMAH9nA8qk9
49bdkzqCQwudE2twl5qANJ5agPtoPyC4sIPR16mmRvuIEzoN0YuwzAE7p/IiDGP/
nnv3lwmQyWcAXUQ0T43r+nKlOLKRkU8kWBXwfyrUzz2UNFBhlz4QkK1fDBu/JMlz
JKsAN+gZSpDT0UJttyNwsvSD32sSvIDjA6wNncRu/XtcW6WECenHKP/7NqcbWIcO
7WSm8Xqe7ArHKH0RsNaxRF7Mm/tngRgNhw7zXLlVRaTCjT01gVuALEFv1xWtxXFd
dKgBaKcjnCqTmWdhR3MtEYqYmkGDfE6euz4t9/uo6xO0JpS8CFjiwU1vaTmezLwb
3z4ZdO9lwAxjgADfNq6gxi9ixBx9Jje6q4CF6SRaE4dqQQmPuKcVaSyFyY8E6yLR
q16yM3Vw8dMFiSMVeyRnqzPKbQELV+TjhOpSFCkED6joTcTORiP1uUGCRX+ibngq
i8/UwH1rebBU6ZEZxbYOGe63WAPUy+KMiAV9UaGBFXyhgaVfYIFTEHGcrrY/V+Cq
YUKXXg58heUYiObIQgfYmGZEetQgvB5PU7nhl2uDOXmgg/ZKwJjDPEtrjn6T1+4v
amBJcMqimsZMOB9WWSNvSdTGvZnY3bG/llbxd01bRlHjkvHglmraBBq+2fnWEcr6
3yudVAwwyMZnYMEiN/5Rywv5G+F507b/su/jTPO2u9Ap+R2wpSl6gK2jJ1plg8Hw
l9P2PQ+rDGp0kwxi79j8kKEAdX1wT/wvWDkhlLZMiqxuGnSF5fk+UzXHLnqXjdLP
aqHlmPW1FL+ir/IeT8pWkqleM53Hr5Ipv/kzI6q6Vzg9++iKRStRq0GuNxr0k81O
B5eJ783/AjevwcNoOw1KLFQJca/zWrkPOoKkG23p+2OQ2eyQj3k+LqVGQAcXOmBG
veXDqhtWDBk3R721D1bEaXZ4EXqnRd61vjFKj7kkkL+ceysVuGvkNZsMseIjo2st
ztQDjQ4cmb0bioDmTMUd3YOwhWX87SNSuyku4GUH8/5GfAOkULUgAKV2MVIpKytz
NaTCapFvb6pO2EkjYnWBm8adJPMv/UNshXZjfPTnAZ0HBsNdVPHn1e49w6OwHeEI
UChzNhAVhoVBMQnrV356Yi9BVbzcyF/7L4VJKoCdLd9StNzgeJNh5njOPBL4RBk5
H3JCkPkaNJsqAsWWdhtNL8HWg9HAKawTCb/uwy2or5gBcNn/DUTl7GT9VyTXYcAH
wY9Z2l9387ExOs2Cl/1e5ioPCssPLQH2dfyEMPdmvRWQhGiGSu+B3fzcjPMMb4SB
cSMHTeYcO92leOvlU1FvdwAnT4cz1/UgXYCp6hrB/kK3zAGHzN/4ewm2PlPCNo1v
2r330xw0qiG+5EFUZLDV59XGLqfTdFEaGihI7wadWzDxHo1YvmbckrAQcyVPUbET
0qrjyi1vbGOwUydM3ZcGaA++Bodx93nQS2/JLqjFjJmxt5MbqmW6MR+Tk52H5xCs
F/FGN7xOCNo4q6EdTajft2zy/E2Jhc5Y8yDL/RTUxldUc/41HODadYNCQhtr/1T0
vqiXmURX/Y2zyMvBStfKgjNPSBhU8cpb1H6eFtV7rLszzANdfy6AZgFdkO8DwwZu
qdB1c0amGF6wNq0QdV0KxLtRQcoKfGGIpoeqBXM85Kk+mk4bPo+zeMrUojhnEGk6
/0pTJY6WCy/YUp/2iHy2zgCXnU0CF7u7vcKkZBaMhCieUmDUyc2hxlpKd+g6VHOj
Oqp/JWc0tfnTlnj6zZrkEGEdEk3GdE+No9KuEV9Nmf+SgFHoRAqI3UQ+Pyad8A8G
+MaPCAxMcNarKFRgDyw0v7HqyC+NgRFKAAoEjfUHZi0bQznKVCpSJYO72VHXm4Yj
6uaicBtOsGwcHqh7q+knxVaAkPZsdMOTwyKcd9E/z7YNzaAKhwOiWfDrt2+kBSQE
z9kDr8Nh1uYinTjYh4GlzxborQmAN2Lk1exx/tvVzZPRiUy7kZYUOLtTFnyFhJQA
0C8/0avqVxUaEZ4nRw5Fe18XQL7UzG7kSvv0UPpTbZ2x575bG9M1CJjhMlORrj5Y
cXCCWJzVNnW8caxsvYb4hgnIRI6FzCB8hkHLG6b5IBFz49/dHQQzqri9HsebJNmH
9MVGVsUw5YPLE0OC2mJI2Xo5OVGl40N/7xej+MZPaUSmpZjBj5/6V1zb8CI0IrM8
0FcSVCu89/8tX2eLIwxSpxrpu/1cmZ/nwcQry9ZMYpEJBGWuqJF2oZh0h9hBf3JI
2thhGdDhoEPzC3QhxkWs0SHz64VAsNOp4EPIuKCrxf3koohkud4JnhnOOvvykkbO
+NYHxl9UXlEBapDN4WNLAoXn6jvIANRBfD7KHkP8zR3nGPUTinx+zN56qEHmVOAo
P5uPLIQFRa03gzRBP/DJJkLYWWoDGICdI4xuys7Sh31e/YbzkNRBjnFKYaKl1EgD
4V6NKQ4SP5mB0DN4LkxI7F/utMtB3DJ22VnEeRFRbx+bX4nZfv0H5HjwDzDQDCvg
TqTEBphZadvdayvGcYbqiP9K0pdqHpYEr9hMT1zYHXOlgFPsQcc0JbV9Qu1Nj6eN
HA8CMD7vnlKCIjUkNaRVxC3H2labTs2aaASpxwvGSTIl3JwNCRQsxD9lOTIgXBGn
B67ynvMaPItVmrFZKtAx2I+p/Jm5aaplybdce9d9WM2dVTKaaD6J4CKb1JaaKJSm
CRaagKLAxFUk8EPhTiWHKX5zGDMNAq6EWYo3OJcvOXaG5kRH3DLFhudjAyOG2CqL
noaXd7r03KdHv4jd9+dCc1SF3KY/JMcTMDDUmK31SSu5+lTN2cijX8zHpJuNdl3O
GB8Rw7rvNriQMFp1ANpfeeA+/O93dbY1fJJSK7pVMOIc2hHKtgJZocGIfS713QVf
gsM07T3uf1bzIxwcVuppGjHsluTjWTg0MFE+ceoPPJa0HlX3P57o/XLaMA+pmeJk
KO+grJcsIjohsSjIIjAcBF9Xp0bKxuIJb+0DiYm6mMWZXmegZ/slEq1q4zV2YszB
Lrjcv1W9lN4+lzwxBwYvGj3TQyvH/mq5oeEUXyJEyDq+sMLyMkKF6Yf7KR5o8b+3
RDEoQbr/9o9xyGi7qVKqi4PxBSWHfQT/87OmBFItRUkdxTVaXSfI/SeLPttgbWme
OMXdk/i2qfANqW3cd+N8G7XWmB5mYKrrQ1IqvjwEjR0QoW8a95J2X2X2MdD9Zwb8
1geil8hP3j2w9plzazyEUTYPJFsEGG9jKMYiOBrG2keQCoEohzAH+8h8xuqZJFt9
loQzyabpGotA3hY5KAPQ7GKfYqtT4taHElfuYwmnnnfXIQ3Q95vMLLonLZ/PVA2P
I10yywA0MHYgj+YFz5Q8w5nNDscMo6dR2DDPx9dCx2M4IxeGGQrpaJc/NvTy/qh0
QYfS0ZhmmpqTzTTOmx1wcHf/NumdrUJ1GGoyIgfQs6ZG+sjm5puqwxmhjvc4YuMu
JkQmeZLrRbDfLULiev4yZBqHpTKwCH2pvj7pGjEo8PmHxoVdCWDReiJ1wWxeNy3e
FV0lNA1+tYMK5T0hMTYNFXrnAsJbI0zkAzdVJ30lfk3OL9cPkgsyTOvxk4BJr9c8
OdMivxlpBuTzfIk6s9TIxuf1kedwfqVUo364S1Y+drhMI+WtXVwx/koBclJ0r4Fc
gBrfZqtr0w65V9MXGI0Ai+yYOrzjDCEpKy4MjOtrF4J7hRH0M69lKvgpkmlFQ2A1
6mA+4Ku8VZiKEjXKBr13qvOgsftj1XxdOve1I9bGTl5RkC4NK85UTkJ6qvwPoeqA
SVzUtWF8Z4bWVWUEeYfAOXh3UItd39qkyg/f8B9kkaBmUW7EojvpGHMKA2FYOBnI
5N+Goa7P3Q3fTeWs1f1OUoRFtaUZD11RH6Gozf0tVQimLnGFpCu+8IVJENTglHo4
Tc2kR1Y4jNuTV+zk1HqEW4D1CKKVlia+Hr+D0xxAEMcBFBKsdMjNaq3Ai9MG92Ud
Q/3DEtXWESFEsb9cj//EvS3xPARW7y+pxmN5GFvPSUm+mgpX43MgIaBQp+AUoO1t
/KXDPK7amHCG50MGPEGuyhfGzK0rqtJS7V63PM+7Y49TIgVPGrLmUF45qa6XGPm1
R5O/2bcguU2n+QF/PSXsikGSNq8uDY3EC6a8TDKvpOsVGXasUtlR0399cCTfacWM
excL8mqmhLzjEwtdjOLCOJZ2PzQriRrrrxspE4Mjb0ZgY4bEzjx0+CAgUIl9osOI
owVtSg+qFZe3ZxPPqUeskdZY5UkInTMYXjjggZVrpj6MV3bWfq/sXb8p9ah2DP+p
epxXM9BSw7QAFK6+3gVFFbXfFOXgB69bnjn9M6RqTPio02mwDbHWDICd31YcfPzc
ZVcdSHHFJnenWWkH6GSJmSDpXXWNFzIrSb9TH5owcr/AziHTs+I/jis4dBja2sjO
iYhd6uHJqniP1PQr4sH9ks0etPOgZBkzzwzcGg4+dh/+Vx65/1E7K5+3eb5BXflJ
ZPPbK+qpXSTY6eC1Rik3sic+vrZ0+Sur0yfMe3p8VfDflyuhMrmEH1ArQORifqUy
Zhz/3HzKxRjg4Cj5jwvqrGQpImDcZUbBNdVQIK1nPTa6PmGaJNEKfCidq0Wp/ia5
7S2ZOJf4RM0qTtlm9X5O94BslwmlMm8LprJC/gNRbQbOgjgrz7dX7PGTWMLVs0sg
k4fbw0OsGsDfNH9LrkTUiLeAJvPeoWlO3t502KSRHxNHF84LOwi4r1tsgU4gl+Lg
YKgE2OmrB9iWiHe9nJJdkPKvSvmCUAT6fs0UKd2cA63zgylvzLDcd67JT/2VvSfr
zmZY2qw0q4AmiGDOKZDJUd4ub4PJLqSjcNTPUnKqu6IraS3xZzkCGDLayArxJSOi
oKnF6PFGlplDydQVOg1EYmZVORhjw7noNjcB7NdyzOyunLrRjV+9uqtWKRJ4j9Bj
gNSP4OrN0FisaTAt2dLg7AHjCY67W5stEbWL1ecW8PhvfY+E+pwAULZGMMpdT4kM
caaXfA7mhhZBMSBaomwQDVeSB9cxhBcCinqFnDE/srjX1Bohxl7SJrJczCSnXgN8
+t5usJBJaeS5g2MvPts57Io25NEWuJxMFvRwi6xwqUKD4XQ5JSMTCv0tFCarr+Ik
/BGL99KHXmmqzyNYlIWSl36pRvHpIvQc1Gk6docf4FYXlA3ikvnugOXRVpwY61sC
WzdohJM/mezp2PeuwcVF2hclJKSm16KLGrXfJja9MwNgYUyMu+l/gDvSbh3WdnYW
GlemkZ4Bsa6evV79ahrA1RdamCtlPWIsLJIg/FsVaL4m/WMJxcZO717RH95vgTVX
bvQ24PGsWvKSBh1KIfpQAZ4eypukLgpZxu7MpVfUx7/VWJPzPXTGp5lbgnpjqckh
n4D+JH9ScKId8QSRKQyH0AKn/HNRrMTG7ewMgcxnJqCHlMF4MG0U01drUeCdPZqL
aOF3LD/YJnHqrdm8AJpA9b+A3OAEe3WK6j8tbDbFS8X3mCBpQ6XarrZin+ht0FEF
8ouG3Sr//OTaTme3zlURDWvOE9uPs518VPThvWVBm+N24YTXUG+EGngIqAHop9up
LuMtbWyllsa8IplkIZEuKi5440E9mco+Qlv9OvT2yWubZjQFPCOs1aqTETfBAaGg
H0TdBf6qZdZHBuZcZBDet49jQAhNdchEZ3Um1lCRRcDVtcrGhjGxeb46ByUTUQiy
exj1o+aZPgjuMI68ksB/4sjq39EYc7V4zugE1DtTu9ltQj7eOIA+yzAMqZQ/UVt/
xj958cxvC0u2iuXvOhWmnB6ZbWlviQHUSosyx0gBXNQ1kbhY6V6iRML37nzMVECj
y/5jV6rTzpbDtwfbBVWX3C5NrNQl/vvLtqIYAurIOVJ+Zvr2iu/hxdzcdR5syy3K
WeF/4Q4SvxWVDEmUBYDQsxf65QsRjrw1Dy5oEaQJnyEPY07Jl/mu9LPu7qhY60SQ
eNIOkFmyflaZq7bwa13v9/MkA55t5olZLkh/k6ziK8+ZOrGDL8pGud6WwTl3mU+b
uNO0yhcWREXyABK06hzIhekYCGOMAO8Gv4w3KNEcznOR8ERErSocoTCd3N36wGsT
6guGy4E3UakPWzOsrRcqmeQbVguwActzMnIcIt/hQHamy+Ftw8D7MWZmZVqMnqRA
jQtKvk7kRQyv9w+Odnrk6FQsHWaX/QpTsFVwjFpYZ+90MShXRsrfDNCLXVpXEBpM
d0AS0wn00+rUubukeK3/c1RUmUxY5gMAJDBzbyTD01d8BKJfLyaGdFdz59eWAlJN
4pEijIXwpLjeFsBJJcuJ/hPlXkx2Prw8JajQdxjBQ7GcUgeR2S8TsLGcI9UneAcs
+KzSrgqJIWuTUISY4BQMTslbiSg/lp2Sgql74IHaqzeXjH1BCtlpaLpeAlK4KLyh
N8CQn4XG2yU3FW5Jhoq7i46QKJpJmi1kPKkibQbZ/bOrr8s/RW4TD0zMRVmB00sz
GJn4r4XWFYk/sUKYC7qmeZ5kicbwlKwgOBmISzYT3aVYwVQqihXYzsOSS9lvyDny
kBhBTeav176Y4JdoKao7s+lssq9cYduje5NNH6cVcvdETDQWQnd/zBm6BIbj11/g
rbfvP7WV4xyGnwJYwBS6rowwejhO4BFJd13qwORBQLlgOPmW7+p+EhrzZjy7btAu
+Pp53Xrt5NBWuOiOqQspqBvfpCTTLf8g/poD5jOONboG1ysodo2+Q0RyQ2GsbA5Q
TjU79hGxbuQXXLHppDFYW8jehAs5lnw1ihsLwFAq37DRH6MEheqqIcxN5Na718WK
PoyBNx2qCI15XDGa9+SnnANyfaywOJeDctXz8DxZzas8OJYukN2CUqKJ3uxzrTUH
gtnM0lAeeK8HWs8q6Tj4TfZtwMl4qVlYM2DM4KCLTAEqCY88u8kRbSaTFhHIOlLJ
hqXni/FLwIgpUeDrnfUifE/vT26yDNB01RBy/id1rRU/DPyTrpyHiyaSw0cuqc4x
CuC+Hgou4vazH6Hl2dvViV7rBBHGMZ7zoLuxcCNVVvIB3+xClx5M9G/IevdsSk68
BeC/3GwIMX8rftqFio/xpvQ/34GMrzJ4D29nMnDSGtTf85m6FAZU77OTA7ROUYOP
jltMeUAm+ZDB1YxYrV4H1RemNFufc6/XfvsL7TcYQ4JOhuKUKiYyPvxL4cB4Flwt
a5ASJu8IqYP0K3zXhFScBF4une65zMvjE5TMBlPmFC0FRSxAuSIY1K9gZNtp1WgM
Ghs77+/mWEkpxOamyLZmk0jm/dWP7w6s7M7rtMkF29y7pYymRUZ4IS2GAzefiWdb
CJBKmlerqmGVKQpBdlqUKFQf7G1er9Zf7ESJ4smkX3oXZtQNPqej82Fiyh3q4VYB
eWAPCobuL3QWMMgCC+ZIev0K1z2jvavllchgbiUmYeww6Odx7STmhhULisvpOpLa
MAn03lGTqBmAhi/DY1ZhqWlNJcwDwxEFqVudgA7p3HR9PPiigMqfH/ZRliTP2o26
O09aquvwpoIRXIVUxrrMExr5YlCOTZ3l2xulvOiYdD3toUAyD6cFNh+QkbefN5Gy
FCZf1n7irWFO4JLuxJXRlDNEhmbvJ1jloX+0FaUyj6ikJWg0jdmQQtVsPJR/YBqm
vdm9G/o45aT7dLqJuHNBj906E+U0vT4rMFLbnB5Jp+8cNPgC5vPrXFpOGQhyqGg9
H5YaFqgUKg+lzwHgyV2mRA5YCa+gpfO9SRb1azXU9ibG0UjrfGK14ewRiu4eKT6C
2ZbuAbMMAtjQrDwIfj8wvY/nJ6KDh3U2F2pUVwha1SdDYpcujIqGIKZEUQeqq3Fc
TDOwDYXK9JRxxF8FHqgiwqa2hj+PImgpMlT2wzqccBxRN9kT7xWIc7BlZ7L5UHRW
sfMSpwDMVnfd8IDEkR0RMZTOh9uWEnOnsEn6RrYAc31a2R+PKmPIbCUcPPkk68XQ
ovb4/L5cbY8hpySUVx9MDlThTXrBc02wJDMZlgfW6pDLrVg5s1ZZUgffp5UzUSG5
jyaFNDAZpaPtchPgOcxliyntQFYhGN0Vdxub9FP0u7ksWdNgTEHGCTgjckPWYB/S
63zXgzIVDPBDirv7E/KzNdVo41pshdDzSqHW/lTD0xClcn9/rN8PP7D36TAyQMHp
Ar+IvDI6+YcPcQMa5lcll1di0X+DWNZwChF2O+zbP5a5wFOulRWYAykRWpyP/QfF
FW8XzfE4f/r/i2p0jqj3QZ4O/AJ6R42cEKQV64LG3qsuL9BJXskd9VSiUZOYFREt
Eu5M1L1MDgL2tEKrXz7lvhNQXotlZTLTYCZVN68df4glK/4iwvsegrObrcHXpE1d
UEl+gLiymW0BYb/BqMspU+ROqysebWdbAm9U9AACWC0drWLepnS68h2rCNzsd1CQ
cmNlLkQkb+h4GtHHzjyzTzIGtGrGbjz8GihbUNXoPnxdpc/nG7Fqm0ukHGyLwXMP
u/7W+d19DpKtCqPP0sa8ifAi7GNP9+LnYAPMvPNa2wVZHhjXb1K/7pzUyitxjtfB
9LyKoe9GViUthnSxgaKB9nC68gag2iLAKnO+F1T6g0UE5A5V1ydVxy4EJ5BmR35w
bIJKMRHy6YxHTuZfzh8fmr7h5fs59eSC4fQkyQKt4HumBAdL9tPhHFTpnCKkIqiT
JtSpaCdIxXDpsJpu48I7FYTJKOYUhucL7XBIg+ytYwhhEDd92GIk283Rb+6QEhQz
E2WYzJ4FjMsAtY4NwVEw/A2YMMRiC8RZgpvqKorYmd36LgWH3mVEl0m/8nabjw1Z
yrPCdmai7m73sDy9v7HYV6hwvzy44+hNZhv8PxROh2FjYDDFks6KVKhIenbM8tyc
pPMI17RQpKX3vqI7xyn2icsOmWqcpFEdvdv3LfpMLH/mTpV2z4fDVy0khIMLILA0
E1ddfs/rHjeIuR2yKLT7sKTQcoDtbpY5UoPqmxxkgYegmcoMB4+6aq8pI1AbvI7k
f5FJ8wGDFfcnMEpLF0FEfhH46zv7N4TROF/rHiL+ZuWPLYnJhdAsGTJJvk5oE6zw
YTWpntuFMgAt4h9KSHoDn0JJFgKgcRtYwDY+41NO0UkXYuHOstu8RBX968/AfNUC
CIBEoS+fUWXPlhk0sFU7xn+2WATnKXncRFsOFwt5koyHD2+Xds/d2Sr9g5FhAxvN
s97LdROK9pqptMWMKR0DFQ7/eGLcj61mpSImNhIDs8+L4zkyzX+Gzpgh2gk2yKIE
vqw5W88AeziACLPqj7lAdAg4g3paAcQq8pc5RE2/jcKsez3a44gx6U4GpGRb4x7o
VpCiQun+11vriztixqhyeFrLYV10+JsGDT2jkQgggybL5qa+nq4JbjPqZCrJfQOn
WFoW6ANquj04rm0dhNifAExlxqwuMaOObHZxQI2bLqyIxWzazF4gwkNg3xF2LPVt
wQcBa0cs0S4eqt6P+pagEOG24RcClnEufKQBc3GGFvHxfjqc4J7qpJW/WJMWc+T0
IkQFlj3dUfI9EvTOTK3Z9dVZDHvJj3sbKxrW7+joko80g6s9ZHYShvHvvKM+msgL
tV9QdDLYqYrYIsZ/EU0eUQAOPb/RfodYgpLGtSCdt6n2aGS+Qq0TGvHh4CL6dqtD
bOHQ0Z77/qTuNVIo3NBHuhddheqUiYo84ViRxtgrmMg=
`protect end_protected