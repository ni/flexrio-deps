`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 50560 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
LfLaKOw3utJqtz02pVdKfzJAd00IHyvKnC1DdN0hYf/8sM69doqyQIMtsRWVpRNz
wqVVXYFLneUQk0B1UV5H6de82WCqSouxJ3cJrfKD6olhbjzM5ErAs6QqJQGBBGyU
80UlhBASASEnwUn+ItMzRRfuRY1gVGNMLLY+xdYlT+5zSWKswSfKNZccQ/zzHFwY
/OWajG7bm7yaiV7Ldh28xCu/QAb4VYHPXcMao3api3HJeYvsQB5BJ5xG338GJypq
OkTUqskHs+KuNYIHDFyaIS7DRNctBTwZMJV4pWSF0y0gpBWdiK0TQOl6Zph+BRIk
0H1QIZayqk4/swH6FoptjyymDOmgZpd6WFGLprMJhEw2Ue9AXWoSIwZzfTdW6TFd
Xk9FMxFvdLyk7ljSEUtuGCU/J2tGIyZ9ywrmuTRCJZqLp3Hni/blwik2VH/MaWuT
emeUoo+EvwdDVynb/YaPSqooIkSeO1piN/vp/w+HzkhlCwWUyDD7gW3zSoIF/PqG
+RN6/xzMwnNabWDa6Ojsql8Jb2QZduBCNPSNnovd446MsiBFhxxlQ5A66iOmC/aG
va8s0jaIJejin8pYPiGupPu/fEjsOwvqK3Ljytuo+EnP2n2Pl84MSUzWgzVX+HxH
E3ToCIAWcrnrVcmzDi45aJwqPRoy7ekv2uQH902GTwojGyAIoPPu5xcbU5pb4WLi
DwozVICpZ6ef30Ns+ANjWdImYglo3AA0apmpHYUQjlwAIK+7o78FAnYX4f2Ibp4c
lPCj8vPWmm+ksO4AwkiYzvk7tgWpvkcbUeBXB0OrEKypykmx9UI/1H0zBF68cGAV
EtEFXzeFS7AQzLSCyzMOuxC5X3/08qi40flLOR8Ty/0JL7qPnQ0A4V/viQxfgWSB
bYcDgJd9URNM2yih6bfMtOFOHGOLvdr30CoAxNdwTzxh77sU8rs8TinbtDkpGknD
LQOyBIdDgeeuhCCPe4W44vMv8yxoUQBxqmv+AZoIY9yTupWKlTtOxPyTdj7n++8v
HQ56eM+xuWDx0LGwPccKKGIVCwzo1RgTe8zeHWRGHqy///yFBO0FBI5a449qtEYx
I1IZPzdg8xyVoaZJhvGxWxSIrd/CO4Cc4jp/50mmb5eyXmqaQgA4kXIC8RIiDmxQ
AdE7TBaDIP8ePuUr56rfxZQpvUoap8Fx2EvUsEHNRy31amlRAcUGGhNsy1M5gCwB
uz9T5aI3vWAF0fyfSJTl+KgPxkA33HuaObTAEyVJWejI2aNDxaCg3jK9CJwoQKxT
zY8+Ll8cOXYzisaNmL5AdgmXl7e0BkluGYSwn3C6NJkhc2m/ThJnw661hyrG/HH5
/kZ2qh40pFE/1dg8OieMjK6MrxerGIh/QPhSF1GTxx7G4e4ZUtK8CxxYIX5fgrNh
7dKVNxwo7+KI74ip49Jz+4u7aDdzB/k8hNMhwdnbC+XKN9sLzWCfrxUx1S8hHhvM
PTT7AgRfp+W2mo0eF6EsHS5Z8QKEDF/bXzKV75Qq5Ktdc+G/afzCBw5C9IPnmw1f
lv7LOzc9XSkEs6Qop6GMpO4wx2wks66Ds5vxhxa1ZVKrw7uJyxQfqEtJMiqxhGS6
ju1GjWuZhr6GlQ6JBsl4gPP8VBsfrxio66lxIInJEJoxxCt8wu91IZKTZeH8DnX/
3lZq8sROpW8NqWMyfKe32QfClwfennl6dnJhgrLzYcyvY5G4pFLRwpCIJ6uFpPuy
74n4eriMXx7Mk0PQUH+Lo5R8U/PMib7GBG2B5YD53jWRYw06DK5Il3sCIGY0sqCq
cjNlJnuREwe9QIbAgPvrn/TKcrBbAdihcRh+USWJCnsVWrD0GgX8mvZbJ96VhqdV
5emLISu6ZpTWlol+ram3+PXJSxAATb4KdNSZumxW9W1NpTyllATJwh5E+H6b5Rn+
0NGEkgQS4qCBQA6C4E2D7OZlGo7mibDnvPjm9IqSQShkziH5FTtVHbM4rXvlvb9E
QPyDaBB1nRiSsRC30PrXqLd6dJ5qx5++qx/wR7nHlD+kBPKD+Pzb7De8u0Xs4awI
Uj9Eg0poek3lbpRxqWe5DcCOGoDeJYi3zBZF4tBAqSLA3aO0ALGsFWZwln/Ch6xS
WTtID84EmM6N6qmTuIg7HDR9+svMpLVeCXgefUwq0m3VCM/IZibgCfAH4cXeuXnL
N8DEwTny4F5CoUO4ec53FkXUwfc0jQnzunfZq8P/vUcLXVpgxIxje+SwgcscskIU
5vclTM/RQPlEK4rm5PIKSuErGC+GWlh8L4sns7aGqhO29f1K9cjHptQm+YUQ+RRL
/C2DiTP04HClnLQLFlcDf0pjKXqRp1hewezoDoi6LfkWSDwE6v5+yHbHrHZklPdy
6/pW8XGMdVf9MizoMcZcUF738buflncQNjK3sNAIwm8a/4qZhUjJg1YhEb2HTlMu
XMIWrnZcMRe5U+yide0UzdYhKsedePSNc02PCRKq9GRT9+Hqhq9iQbw/PnaB0qIl
EIZME7ypaW5EriJ9Q8wc0f0NHa0A7AjKM1brF87N/xq59XRHRZZBJTTrSc9R+xDc
mR2+i01bTwn9guzMnYjiMD48b6vLMNpTmfr/iL2EWLj/CXQq+IWv+vdQWD7EsoT5
bkcm5WkEb5PM1hK/2ZjCQtZLYaTONbIDUtXMaAQngYwmiF9Y22KUoQT5wHnZAToP
qQY0+4rGyHtta+HKZSRhQxwl3GwH+9xzCELhO4rAlN5Dhpfpr3jCK+0yRINBvEFk
n+/oEMRTFVv8F2rd9wKFuRPGyftyORy8Tf1yVnJJ3uzJzGI5INOKkP7OuSzF+5uL
oTfKqS29lzjkXRS+cO7kLbYjtRnj75CF01jLSqnF5J9VYNP13wA71GQ0Xgfm8PHV
Ki+4R9mzYhG+PDmzb0rp+wF2het/IzT0ttyFU+0LkYW99d6z9hEVNqSqqyOBml4x
q1h+pL2hYE9lOdQtb7cLO5U0Jq8crWtHgN0tHnkNLTgXowb9qQHrIO8HjrzzxlTB
N4Wvybe7pLpBIadD9BnXLDPUu4hcFBbe5plBG8+q9I6PCzUKiIi2XTv8D/v+w+d5
qwwEdUEbcuz6385/OQd0p3BgSJZkzDKwV0zvK08YA8u8ZRTy41nbe0AZT6DHTg4F
bRFvstWTw0qw25CtY4cVya2gg0XR0Y1CtRXmRQl6AjOgNcLvp1JtnJZGSiwF3rv5
GoI9NZHOBJMD9o49dJBh7l0eKxO3JGC/tC0RsH2S20tpfTATtquJsr1SCXO6yhUC
d7d+wvwIFOrD+bOzK515QbiQfPCFakuNndufAl3tFJVJTmPTfjGYKYZ2OvNJrz0A
7picsr6wzRUQcLPmhKGgj3Q4vhTiJkUj2pRznth/qM+gB4kl3ma6UOKb6Os21j8v
9puiADUMLZakzusDr8lLTxYtcRHybPyTva++NYuXv0ULOoNxycK59FfhXs/G+MtU
NHDIPdGVxh4d0BWOq+/rMU7VaryeiT6A6WK1coZaYrvc0wfqXpTjt7LOUyr7jxqd
1SYxrkEzaSKO5TGh3TtF/lDdee3rDdW73UtRGbFGZ3atT/xhehftCpm4cdhr/QHG
bGlp+5Y7YMqo3nklX4b1yOWXe0MLUBo+Wn7K1dVXPyLtOj3GZURT9JLGr/m8VIgO
jL3jVCgp7OlA56eWqgN9S2Rbp1ulEcq+ROYmbZnkIM6UqfAW9uKZfAADXv4IYwuu
9T3zdQqfjRz/A3U/YAPOrTLdE6ZNJ+wTPRJ5zEIiz6HB3nNFluW3DnrUlR/InOUM
zXFCcg+2mVDRAqSVsz2FIA7sBTSbZJBcVTCnsFNfKiViRonvDr8wOTSFugaXeu6D
UfCo6TArrMoyHFrP5sPAJe68iIGjCK47cuOx7K9tulVz1gvdXGcvUeEWw+OUy4sC
CkzmM6VLCf3k38XX6/UKhwKgDCYaK+JZwxUTuUHWfCdjTMW/KALZnIqRbiSbLDOO
nyXXA8K58XLWBcG7pw63VpxMxpGBkWjMk6UWb0i8ZEfW1x8gab6C967l+tNsGaa3
DTZkIm6qg+PWGFEsycE9OMnHwxeKBfFnznlz66yOBwl6OXp3BlG1CRGO9EJ1Gt+o
G4/SFIGWr08vGGqM2+UWVxIp5Ee4S0lS0VjmpXOnridPKJFi7Nl4KDqw4zyD7d8O
1DQreTBdfaTJtENuxz7+MU6h7bKe7HGNoi2V2m35teSUZlIF7+082/zhznaYgwlo
4fDvg4GbFPCIvfcnluL0s0MIdbY6vbgzjm3B+FYIpiL58mVevQbGN6Uw0sQF17DG
mgMDcdWUydwEfDAgujL1F0bIlxSCpKbtBE3lNQk/AJdh0lBlkUePbmuxOymvt0r3
8fMiYIcfchGPnJ42a5dj9IpYlkWuW8C4nb7YYShUDo6KG5VXy17q6WkoE3vegQZA
rWwbM5bh6FLAVZFCCWKKdiNzoNr+m71ZPcIWSAC/gmlQMtp081ash0kBOUQKVzeD
JGarEZloFjSFK4xR+KHL+OrKMicERqFjPFYOgy+CbHakXcTqv3OYJP48+2Raqvpf
RV4rcvDOcpT0sz63NuExmZAedVpynWr/8p179Cz6H1AkwExZCq6MBAd/Hp5mHMUc
et/om6wCQg2WcLTQxV2fbJxLY8MuiUx6ZTp4nWqJkaLQzarYweNq88iUI6KCYxqF
kruTuk1YLm+MVbE1dJxUPaDjuStOHRiu7jj042d6jzyAQHdSpCtxItyws+cjxT7B
rVYBRIPWtVboNhRjw1NXbcllb9eO372SC2XRRGeUq3LQKIJrA3IU0DmaXeQ2TQZU
Q+ZfQhHW8c/Mg+k6dzd7rbnnzjoXrKGzHluWSKJlxpmZCJE1siZ6s+u9IVPG2zkp
5epXko9g45Gs5a669HwAMEa6h8/cNDqRN3k3Kq1Ad/GM4HmzqRe+yGOJvk8/BFzv
SrcLTwJy1r4SGqSQ7Rz0mqWYBQvtJJRM6mXLDGBXWSUjvHa8W0IPe+/nfb+jjW7d
Ps/kP2aM8lyu6vrCZZUJNhjMfSCSMWJGffbjPc/rvp1OMe7aVxrpFRTsHhMp2PGk
cJzrHuM3DV5VXFowGp93OfM3Z2MUghp/zGlfeOZIW6n3xcI4A/3mm2X5sAT4Oivc
H7QeqzG3IsRhKNOKBuTlmXZPo9NO3DdLKiKyiofV8nRchRJXiEcW6r79cgg8HewQ
2ocyJKQxVvVpFMdJ/0XJWPee7h5mcylOgd48ZA/ByuCzUTv2WqWmNrylYb5CJeS6
2eM+MjD6YoAUiYlMuscit31plkB6k0qhcka4+gfQAQ4MNyYiuor2sD56Z8/5LL5D
nYuFQ7q2KnvJa5R/lLTDRdo0wi7hOzzoDuW/66N4tVbJHS77pIxIEEBcNV6L2fh5
z9DTgM5gvI2Ji8BJ+shKK4fm6M88kJdzUMScl4Rl/rf9jKfRSFlIRR0CWtJuDZY9
eET4IV470Uu12xBX4rrUycNurmNP7xLaSInr978yWnfCTPHmdtYipwlr0VT35w89
vUKfsexezmxOcFHpWh+jgRvj0wquyQsY5iE2iOWBJdLATd+mwMNPD7OQipY05sQJ
GHPwhYWb4xo46bCMp61dGfc9R6iiZtIymaCNc1N2ACR3sr+/kHc3ZioLWlT28Xaz
1kAVRmLvFyRJ98wVyNjXLS5oXiRDUTqA3/K3jDn4keaRvNbBv8tc65tENpy5MQUX
EwonZ63nh6Utj7nBZgQfnCaVj0W5QXNcoOUyRU/YHuOQIBJQuzh2pxhuDK858+Qr
rRoTqwF07OJtEm9nsdyJ2mpvEeECkcr48YXuc+NOnh/jIvkYlxOBZMNUZysoJWCK
CW/41DGkxITxqI0VuvnY9LwzlBVBiE0bzTo7AZdUIDsfdBE8TpymNS6MwYrVjD3o
jLytzxyXUNGxnxaERBF1OQrWd7WXoN3h/zosYlWqHLtvLdRQNc4HkkJE/NjAsbSm
OdkbU0VF0U972VmDXQK4SHmMyCGUuV6h+JvDQ2zHRg9+WYwl+99VXb+rfgiyRuMc
b7s/hMMv0Zdl6O4OOBV3w22wBZQd6egSvqS6VtR3udC8j9MjfIvhUfBZDBqgts7F
KFiYOdniMzQok2YXgq/gN5bLyGf8J1B9EwWek8upaAAXNZfjkxrIfXaYCylGBdgJ
+bfmKmoWv//SRLUPAqcf70i+wNIywRFCZf7TM4pGoWi5kbavic7604HKxaC5rDk7
eZsXEoBRr5UfBFtezGetKh/7c4kEo+d3oAL0SCEDjKsHy/BWbnlL57Wr41wEYS0A
nPevL+Wz88XHuD8rWVgkqRjAun8YOaQVJZgB/6xxJ/qWb1QuieAA3b9qN+boaYgc
yRRlAHFnpOpkZ5yZtQEFjPZNNFDjF9PpqXzr3Ec1jAmyKoAeB3WIMSpkt2+lwX8/
kCfyF82UZUBOf911QlpdHdLJJUS/SvRC+zurng56Y3reInz95vYY5V5dMdaIik4n
9aaHGzu5sbnR+1hDKvJi+oi+APH0RTmR1YUoSePeD3w6xGL93BgbuPdF0A+KzeGy
Mfv9vMMpdsI1pqnr4tF39tQtYhJP9qhPeCs0nveKBoc7rP935zF38uGjtuDsgZmv
/XWenDYodr2MzxnXdiSi1+RFzOX0G+VITVCnmytI9Fbc1aJAI0y68f2rfpLAMDrf
WOR7GBXbD0NZmglyOdw5gOsUIYn6ujTCgr/pFFPxxXFGFwmP0WUu3yefXMxaviqj
YvGvLRwkGnWdgtwqVNcNF3yhIr8OdwsJmGqLIj34+VpiEOzo413u5mCYlsX1H1qW
JILQN19S9Wv8NEWSEELsmyFVu4eOiF0gZgx6Uh638VVPXBBcp53F9g18fSTHXtZ0
pGO0YJAVL3KNVZsbcopihhtstXxh6ltIgq5agVLBsMDbDSrU1LItVplqyoL7z77C
H1LwJO2Kov+evHGfga6p5KZLnJAO8XKeVs94bbRpiPfJHU69wbjSRZAVBgoWDdar
ElWVhed3/taDQ/NPe1+9SDOWOh6AItSUzl0qEoQnRxDh3qn2EdoxrlJgpYslSuqI
E3TfiT2keF83wmynTMSBnO5x3xvgEYPrIZXwMLSq4MCcuA8fYdMkyX9smdZ9MkXG
Z3pxV1g2GHufoUvQgNsrOSbQori8HdtD1xiG/yau6N8c2giCED7gnfQOzOIKy8UQ
psRU1Yt/ZKNEoYC4zOEZRb9LWk3x6aje5Eo9kxqlVSmgItqwKkt88QiZ9vrLuNbj
WXVDXTOP2oFL3Qdqp+4ojna5WM22OcVu8Q/alSWzOuwRJmKwku7GtyEMmuYFMExQ
4IGRCnFiZx78Oy+j4cV4Et8Y89wpepgL9HUsNiLvZKc8Rsy9oynfKYM43uF4Ida/
35w8n6HCo3j82dTj6yR80W64ru1cmFoc8haF22FRXaFt9Px+rzZNQdsybwkuoRgj
nJqamuZoBijnhG8EyQ/VSgc6Lyb+on9tXOoDzUMmIx81bpToJF+eJ/GTiHUMd649
/AtwVPv8iJBMCRNl2Rmkdk/YBV7RpBmBjBDanuQGpVoI3DJeF94ZbW4QhNFUqAwY
kluBPLjvbPjvpTHip4z2dWV5R3fL/KuqOgGiXErz/4Zx5ep/sr9jdPZp8Qwc/4DK
dvPGjzjr9ctEr5SJ6bBjGfoSQFWTfeAnAlv3H7Bb/RR/Po56/YrIbQVGtSM2SP2k
upzBT0OhQc7im1m6MDq9GC4RrLNLyGPC+T7mi1BNvAtOv5JC3bjbdiQYSTyFZ/rp
v4QrMEU9UVej9JLwQLYU1xvSYE4yGwfrbHsbsz4d1T5bT8yo9TrfyU3AJjaWmAbW
Rym7OuxY4gP4kEszbaIhT96bwryUDm/qv3jmq0bs8Kidjvd23cW/4eI7Vuht8f3h
czRHfG7Qqxzo2rPERPYmnax9ddhZ7Dj/1Plvv8fLtWb+IOc4b/E2lDdooFKfwdTr
EdVQQcIIOpYV9yZFC+E8Ld4HzSl7K1L+ITo0jxmUId19nYQpo+5DK/ay3VrFqDrM
J4xfGGe4k6HxFliu35QqVr/ZrtisiHvRQEn0UlEqml7EhCL0XBAC33IeppX5+C8s
4Ufp6BGY4KD9Q3EhnS8n696xDlGHVFYxzkwOaA/cZKmIg17jh8ZGwlTPUZ2EAO8V
KGVsJJylPYL3gCK4Tbokapz1uG7aapRKfDSZ1QUvO9rtdhbLbDcRD6RiZq1lN3yt
V+zqT0HWomSensVcpfNzeJTT0VPAPANkjImdVmZAcXxDq9rNRgKLlY4TX6Ef2ow6
k5sYe8PNBVaHo6mYV08FOCyNUdOyTijDffD/paIXirY1ql+r2C7O0X2MkVVadxWy
BI/2rIzR38ogEQcokhFs9Pf3gtICyXKARqdF0MBQao7cl9gYz0d6qf3s+IPmtnvZ
SeopotykhnDvuXRIckmqOfpBrKVusxWGvTqseAu1t0TCwJ1la/kWxgZm2iNiVcOP
X44F0UmL/x7N4Piq6hdXxeOA5DYMgwC+37wGox3SxMbZaGE02zNL2KwnXBFotSHn
DKJIO798pbOlmxOc3q0sZGgMddJHCaN+aN9JuhH5TAJigUeruKyHGTjv223tLupl
vjh+TmxjU7jZYzETXEfQQOuINiyXSRFFq5pdhC+dfTlr9sTTdNHx8MJIMtFHZV1M
KGzP5vWObKatX8gfqntR58JEKRfj0t4hKQF5Kq0vCFhVYd51iNmdXKMpON3D9a82
iba0oVevBLN/BbW/CNX4buzy3FUOP2sLCiZazcBV/YyTg+9cRFJth2JMx54Gs3wy
FTqvsYeIMT/STdpdVwkhW89JWT4vj/C8rW35fCmRit7Xr6pOpYDSpS4cbI0vWCK6
az1J1wvbk0Df8hGMQwhNFj1n357PKI69fB0e/KsN+ARhWjkDHASL9P5w7xZW/QmN
C4/6ljIKTkszB3WjNUDshY5/Ur78caLpgC78CEzagDAn72X3tK6EG2zmCtGZcq5Y
Qixy2ph4+Xcln6X6dNbZhsCPweBscDGYS9xqnF4jwfx8G4dWnZIYsr/VSplyQEEj
08kX73D+vA8Cpupb87ssb/H5M1WvyHgoby2l/hYs/XIPkbNkwf/n6Qx23RsqaWW4
d87mV0kTwRoUaDtxsGjvCCoJlC5EwN/odceflgEcv+QGTQmYzsOH4sqzmGAGu203
yrGJQCm+vI955gmIHIicT3V6ShA0SoLncQ5/yRYOiXfY28vtZEw9jbz3tEXtE2lf
PuIV/jA86a5tYV5N742RcDLSkIgW979gdm4hl9wVA+V75o7QSsON53RMiiHpiyCx
Sh+eTfCPKDLCUEe6NsEGWLzsh9HPdn7Tbpvbe5RAw7/0rtSbLv6CDMWuVW0mF56a
RboNhDD8IQbAfhhvHlKipsuZ5oxVeAEmk4oojmOJB6pbzxHMXmtpf65l3Rxh8vHq
m9uftpt1dMqoUu1G1utWdbmgw9cgQ2BD7kHPiEan7FYX/TrIqDntdtIYw/1Op5lL
d2dkiROapq5SyV1zFNAC0icA9ZABv6D9HsK4/AtHESo/VDuGhR6ndtrdGKS2yGt9
czjvESU7WTrf2/vs/7FfuhNmQKvGMuhnCKNFFo7TjpZZWfkTjhYmkOjHq822/fUn
D/sHrbufXBPYpiPj7LKm3bwC2G6VOCPwiM+XxbdjHwVSCF4aa6Bmalom8iZTo1kf
Ydmtd7p24J1OJVcg4OHrl6SB0Jt17Mh5QLEy6SjlWty/p9KDCLZSXK58eE4LT5EK
D2H3llGqHagXkR8qlfCAI1OE3eyqrLrGzsfZ0sZY0IFNikqRPCidz+f8/CgkImmz
1F9VyV3PaXVqeodMVM0Zx2M8NaIpxrvKCr5bf8bi3IpkQPpdZ4XFLacmBfU5H/D6
mWPOTMwb1yi5kRgtG4Jt5Kl5HjLB6uJtzZNZULoDHmk86xUZL/uQUzIhhWTn/TXK
m9BD5giL7xLe43utVrNqzM4N1HPTMjAo8GlVfcXuphoenl9SZlW+oezmyWsPZ2L4
pC78KdzwEIR4ehIqTq9V1KMhuWAaG+Yw1130qmksjdlMgRtewugo2AxoholjPxPl
20jiuAkvp+ADNKIdOcFweItntpqdeFOdJpVJJnWE2lVFqt1bLNtKRg+DN22bMv9c
pG2I77EifKU8uKqudR1GYwZRCBAy+oFCFRL7FlDWVCOO2thh2wobUjphos8pjLoM
KvRKD/u+MpbWdby0R6TMZeQay35kFz5rjM3ghCgZVC3CCK3s9Ed/6LqdTl9ib+Tb
hkwVW7OoazBaa6q/ScRja2rj0zHwiVNO56MkOBaPlOwidtlr2nmNCQUPeINVGwuP
L1jsX4VAadBLSwVO5H4b042gd8H5D87pEYPDOzYT2omTl7U9kHGJQATXhl+Ux7US
FNGjNeEyrY4OKdz05WLnjgzVx5tWTQT6UbIorMkHIEklPIStBK/dojWsTQxueqgv
GyL+X5Q55mlYGDX1eFNytBiUJGW+AGcnZRjWAArKA6gCdQzRGX47+R9Nz820tRRf
TyzzscyxS/z3DvwQMXJ90P26i42O1KOy6pax+baH1l9e84MJH6DOCZvUhcUbjgqR
zbfRino7TYVd7ftMeVMRSTf8opKVv6IXFOp79nkECtpOASb6o1F4xpFKgqK1uOLg
iiPfkhfz7I5x07W3zHjnbK9mehGy7pG9N5NZAlJCBXsVuwGJ6yf4KlpOF2lAezIK
Mj783v2qkVXhqoBWrr5EcxQ72Gh6ueyng2+WKBzdxvf5hxHnDAMt/j20cNuXZIER
gakP8OR6jTBnE+vebjm5mgQZkwfPHnmA4C7VmNORDpxMaFA7GOLKw2P8g7C7FOpZ
9p5CrLP+vYh60cCbT3DERFcr/ILPo9txlBQVgOkwZuGx4xjf+cEy2C28a7HCAMSx
vFBce4R3PrNUI3LqrRsDkMIWac0RqLH4Gm9y454IN/xFjhux7mRhxyubH99FTioR
yhVygF+yFE01kqhH6YzvCEJNepbp3rXVi4UOS6xPpP+0QSPhwKSHnfmOHjMagikp
ue0UODSW5oLzAO+mlCB0skHFo0VYAfXSP/aJmIU5JubkIEKqFwI/itSOMOd3uDPO
aZixxgLrU5NfNnSlIbHWGHy+qwGD/WUhih5jnMXWJOKOzjA5as/quD8FiFDWd3D9
2Ij5wgk4cvLZHc5blmm1RK14jRnb7ag87DvBacJMiCAEF7Uvfxqo0dPiSoJ3eMTP
l7+OLCCB6OQUy2eSPPGwzGJIfK09Pm+UG0NNaF2HxqPLxOMqWuAcPp8LTasG82sJ
zq93FTzmRZXNqrFoAJE0JfVDHbmbEV5zIF9tGcm8FFQP318iCrp6GIL7gETL4hFG
x5jiRTuJKDT1B4gJp7PLaAWPV6Rd/BT6+vmsBWb6kbNJDtmdhEXgL4mZN/hGe7gC
/PzTQpOyodnYeKu++VQfap5AbQTQeovjQvzh3cxOBVaHwsZY/LxDqowXIXfuWQk/
iu0JNldAtotPG6iUrYVmzr/vnL2KHGBGw+952k2rsjYev4+QSSOWXBu6DVAeCb27
IA/8K0qE5En8zGjE1OFyBZ2unPgF3q2aTXQBTvtvp0FRkMcbGg1LyE4ze6pi59wd
eUQAop8eCKS5wqiflNCgPLcudwEAkJ0xSddU3ltOjYo98HXOxTdECq22kC5Lthbp
/bo5NHRFjcEszRefbyXaCP56edoQvE3D7aC4TnhXz2WvsMSYPaSiIA6KSq48gdcL
ZqVQcilaaPeJBUZmeIaXXGjSrvZmcZLA2/GHebf7ZDwlO64LDZrHlxoi9rJGbh78
cz2e0BihXAFbH5dySFJ5pABWs+x/FK5GuW1mfSyasJsekF03tXea5D/Bmbddwg3G
t3xBaqjIwuYsULx3MsIY4bCn2gHhL5aw8FgBjVPL6QwDNV3PfHBqondb/A7/vXIF
OecECFHNuxrIUp7PZzqfLFh9apCQTI2cyZCKezXFobhDqPvz2iLcMDEfIfKqNSGd
+L6iW+9zmxr4NUqRaPpHyx18qZ4rOG2ze29vBVj/FCtDyoB083vquTiMa+Gmq0ZZ
h0EQQzT3nDsN9uUpOXHqlI5CbI609PYg8r13PY5mfSghy+ksZ7j4acQvciOpybMG
XpEtimxmvlwDU4mbkDFycHHxkmXbfHQilmtHUREbb6TNRr6Y93OFe67oNwDJ3dro
eEws6KxEYNlG/Shi/ZBVJVF83GhxAHrl7f1yuRehwehhBDwJZnS1EbhyEZNBxcQO
shwhO8W2pYCMjkwnWOCxdMNhziddyQ8Cuvlx0+Zbunkpok3XLjWcjPTG7cI0/3xv
I3bGLE/Q2GVoM1h4g1WdB/zyCZOz4/tOSTajXBQtLXlqroW5jLmflyleXi2D4teo
4IP30Q1INrI+2T5GJb+PrsSAcYPnLYEiZJk1Vd6jGnwKM89WXb+SOobzI3EEPI+t
0EhznCzn4Cfiig6UivBWzZXLzy3eJrbuXYlf55Z2lo2b/abSx8KlQ1AjQT3pHnvV
4W9eIkb2pbH7jLbM5fRtRUrLW3qJyAGQ9NipvFmXYlDKQCgyFlvqMy96HGxWJxP3
iCHrDm4PRLrr2+uJvFh5dCzWIXad5G6eJHq9EtglHe7QnQad3DINbdwV5MO3r2xd
Gies51qPlIg44o0rGzgrHwI5BOibOyjyzNlkpzuaGgDAZdVstKE9pvbz8prFGFYn
pz6YAMnMt/JEIWKwi6+OGY9mHOt4+m45yoPWYI8Ppk2U8mzciXfNNAKn8boIrwQ9
BUJoIS9bpyMnIOXsE6lzLvSjUv9Eanh+XVKMdJwlH33SPV31Hjo1DDXF6DSSs0Yp
bA0iw5k/UBWWUVedY8R4YMOngaNbOBu1D5QghG7480VQgfQ/INpdcibYyV99LmqH
emUwp09u9D4UqqareYFMk4i1EUB6Mr4sUqhzrTiVKHjvW67IEfPt1wrMrdAxITl8
rQrVTwDxtKSqJ/C5fW4jXBJWzjkZUJuGWCEzg/Z3VpT0k6cDRdARLRsrAhgQPulJ
05DJpWxlzUFsjj6b/2D/ZMRTEgXdnaLm0o11jZs7mN9W0YK/pfCnaI/VHDWv39oW
U2EpjR9lnJN2MrH2OHtcb+d70pv1V/f3bKXM0vcdvdBqyPG9im0IKi6ZMdfgDHrz
cW4PRXeP6fH3mXHFm+RvwJogvLW/2Jt/08672brX86pVQgIlNJ0L0hkhLhw57en6
40nHDtMpLy0a5hNvw+tBGlGz/VDZyIXytO/8JTQFiLiFmYcpw6Zh5bpbCtigadjx
yhIvOfBKH3RC76j4praK3PogQ77zOZv2nVwrtINVs0Q2RURxcwDGXVtBQ1Wi6Wd0
4W7EtViMSmY+JEqGMLKTb18ncNMvja2VAO/buEQuv7bbX789N15Z2lAD/JQ5PvXO
VgCbu6U3jK2cI4WA/uUw4F7xBRAQP9MdHSOnaj0JajkEIY59VLcFpK7QKAHh3C/N
6BMmeIuh+pBd632CW/zM0D+3FP2+CjSEkscU9d62S4I7ezmXMcHUD/P+ghQGZvIM
GzCWIoLwubiiQVVotPcHhk72ENEbAX89Y7FpT0ePORLxHiFV6iu+cui2E+X4NLlo
vghEnVwC0HPLMgpLc2LUw0WDEbq0R95+ZkBG9Xp8wl/o/gcvjDiz/6vayupxqbEZ
mcCvXaLGLyPkFOPeX+pfiZkv4TDlxL5fekBIHm9N8/zMtEw5bU2ioo4J1pSxugu1
Zaq6gKDst3avsGejuJpsG0Trjl6rX/ZqKUpD6lAuy9NKJnf9GeVNZ1/nHG+jL9dW
y9tBA9DUboPTZhr9nAwGZ49cbR+xTo65t7yPJ3vxn4deWdb7wGDOXFnNykdFZ/tZ
igmomFLyIuRpSju/znkMbScPsL0z8gnxIVH83FVZv4ZGJQ4ZRa+q4UVfuYGdhq+k
Bp4NXl7VFqY/lkNlKLZVu9ENAnIkM+eR4RTjSqRRe5ILtMAH42TrFSZzqDRMvhy7
q4eWJuFvZqRDHwdTiwhiq4jvw85kgqlyjy7yate6kgimNxwYCjIULIh688jWNpGm
dOcRu6a4vSH+rxOR/g5bxA09CluEBbOX4hLrOl/8pOQ0VdkDKttPhdMB7QFpX3M2
s2Y2Lkp+5SYPoDn7MXa5BryDnklv48MGTWilp3Jw+WtG1PlMzhyBSUGu+/BdcXRB
uft7Zv1u4M1Iaj8NKaUe8vyS5KuUMgEhdAgoaBqfdnYWMvMtM5Lh7E9vlkimbNmu
FJNYoXr0Bh6RMAwZc7TKCxhVdZKgIvoFqxblkq8s9SCLe/9x99kq8FHhgIgS4fzA
f+kxe8kxDhTu2rXBgCfvRyCvsx2cJ0XtwkJJb6UxiZf/Uhz8xVCWNRHIRhnt5fPj
KtuOJXb+Ye5tOFKFSAxJoRsknvFH46un3NddM7AB58zJWIYD0v1A7jv3i1GOp/BK
RtaNywzvzhP+GkDpdsYxKt2i0Z70ffKXyxvgaa1LbiiXIgIctmiTnzvjRL762HDM
iEp0e4Wh1Ibr+gVNDk42jrORgKnyTXaLYp3GCEkQNRWgtCMjxR/dImkhfo/v/BKK
ZQN/QVjrS6WHZQ4/VNsBM2rzlyhSx1UyYNJXRgCYHlw90zkMbRNKPINN3khyB70V
mCRr+SyArb2N77j9OSZJVxwXs3/jmIKtUcjW/pT2TKa5kzsPkGy+00VOq0WEjqon
jhf/k0foQdl3lH3iwEOP3MUdV7PR/1wlUzr10ItiX+PGFOVX3NRk3eHxqkSyic/l
NHPjBCXEAcdPu1Xxng2Q+Uyo5mDHeUXDu/OcGQ0a9nawnZ1/z4OfyfKPt+SG2RSg
1NFjJ80iQygBH/F7pQx40/XQdnW85qWjjZi5kI6FQN8A9v9fPBgngLlxnnhCDTzv
wa5Jq5G+EDKHAIKWuPK9w2MgnMGZpXtAa/eRvfb5i0tz040SUmeJuX1esrc29u0p
f9ZKkygcJYr51VsPLgIE4laFznCR2luumn1HjliJDNf8dShqY3JOsX8OTIX0fdcZ
dnPC5oUWTWbENnVp34RBryssqYvRl+TBzaIZZ4Yg1z36/aX2RxXB/jgqWg7YYjoN
b5yZqcZUzaFqw6i3+2C/sRL8s0CMz/vNer9e9Trs1u92ohyRTq9mktNMHrdOMmHF
x8uX2fjTWJwm9qJd9u99YQuCYLOqRJuXvPSyip+HxSuCh3pQdHOr3GRe55M/kBaB
YeCtHOiaPNWh8nVBgH3rW5MmRva6acw4/usg/OjsKYyeqYrLFC18GWBS4Vz+Bl1Q
EGtDPEvb1r/iA5fAX/ebEaR+a3aJWg9xM8ntbr803Iy7fn3jUmVph0HsSTL2lF5z
AOqTMb4iOhTuBR2rbj3yj4Z8qV+0ddDlzclbdtFCXtTRjq4HVwpf4FPqrCP7tcI8
n9nYXW2kNnw7vvORsZwRRinftT8QlirTPi35MufFuvKQ0Sg7NKtCW9s0+Mk/HA1K
+JYFOFJBJeP33NpD+eSn0I0RMBjj++ljwt4Nu/lIBhi5SmAhRT81iWVjvx0aULU5
BAJz/B+dPnQ4DiyqbM85hWUYgXcBSqmao6Gt+KlgwuXuROhb2XUFTeLxbuy7RfuL
2U2sv5eOwTy/3MrQ5ETmVNtOo6XU412yCet5engFROKcwMueGKd6jH4rc4yEjK43
bNaVneMYWCKp/LxDXgoZpYj1szFZ0UlbQ0i3+eKMEKXg4Xiya7GatSJMa9UHVWrk
Uw9NO5hwPrWjIsJUrIGrJisRlqxTuluH6avmnlmsGCGhoqd4PtLyUPdbw81WFy95
lSKMrl8bnVmqWAoftc5RTbsbjQ51VZ5V+mECRUdknMT+Jv8P4yyho6T5g1vYUHUS
U31jVDsjHkUv92ErzRzpAA+zi8QUBOKmy5LcKeQ1V8KF5aV/Lebmy0y+1Bm++7Uy
k8+cVrUe+EQbNrQ0nPiJ8/98XrTojzKsDc88SPAiot9OWsoYko2IEV1r3JHkSg7h
ej/VPPiyq8jfspgsNVm5bpbACvyzow4jH1NxJ4Gwm2+RfRBzdo2PisXrhQejGwjE
RnZig2y/ZmTL1TRmlEhuq87iXfy2MVQRBss1aXH/XvfSh3quXeLgFs7Ma5xrb7Iy
58I3hEUfXo6qRB5BGrGqcBcoLXHfrWp8d8TTye41a0LX+pKoSLw+KQLY81Huh8Q4
LJMUGX5pNA8TYlcDSHUO/IFP+ZEUIrrvP8Ti+s3ZanF4WC0psNzHf/UmTYiOnu/S
F01Xkf1ryRJulHE9nBPZUJGpvUmZD0FqJxOdiuFdAWF18xwMYd/uDrJxc0j0Y+az
L9hKKFRqSmUhea5Kn6HsxVwY0rMMHv5O01pRMX/XwT1KXWSyiAtz1CyBC7TwqU2t
vJd8Qz4FBT+2YfREEFgI0CQj3jl5YrA7yDDcFvHZi3iaEYDubAIpSJsTPjL+2O2d
S72gYi/K8jLCwJlF8xaen7xYpoDpP6+cpL2+LjbIT1SHk5QBgmoduEMKaBRW9zp3
RZ4JtS01k4q46BZhiGwgEkl6zbdCID8y5ohOzaH0IfIKNqW5m47o24ZIcQ1oCAOj
jfYPDSHE9T+0lFosWgn4ynrnEC3LuTYJsm1btQUl0tq2NPf91FjS1P6wSdUeSxKx
2VdXPhoYyWuFxZPN89JfANx1j4l/IimpLO+g3iRxerHFblqFclNulGoZGMkNbVeo
gTvPFzEbDRKTSvIGLe7ihS+KwAAAjtrbEckYEuWi9HLTTSk3vJGhlpftQSysoylL
Ijsti6WklQpnf37zLkvdJK32wVlpCKPgrh5R71v6XHTgsjrzEVaumJ+GyzAAW5jZ
57NGDB5WuCX4lr8prz5dNl2XXyAsxp2fyZEpBK4b/jhy0PUfbX8j/bZOEAl7vXOX
8wpcXBLQjvGTK5YXqiWPcFDITKkYkVrt0ZCXgqmZKAvWTwp5vKtXeXnaQGbB3bxq
a1pEVvrgyLtBWF/Veta4eXItNqz1fAMZlax0ynw48a/RZn30i+vaOcXsvYWkcN9R
ZsaUQiwb8D0iXCBAjJvTjQZfDi4q7KIgc2zytZqOeEzL425IzHTDtMoZaqrDgt0T
dfiOlbQd3L5d6CVLICn1wPAcX0V+yFNnp8/yVTtUWO8JWom7olbOPWYB93bRq/7B
YL5CvwXbJPObdLu6pDJrsTxg+KtDqehz2mOS4++c4dnx1LiyXHbzWW8+ZoCwNZfc
LNwWVZWzwQOXNXbyI+y+8ZnDxG5+VoeLkZQHhfe9FE4pbXIZJIczwn0cj7yRCH1U
wWd8oObe0Axeglf3Y5YqkaZZ7Iyhh4yEZW2sIX8awsnYs5rz9hqM4p1yQ6h7NDoq
sVMTQmDweD9+Vu+xWXS3Oz0sGu1YSbpsLwf59pu7H1NpQk/5Y11H2Gu8T+RQXHn7
lObQHwFHewhED2H2fm+yZJZtNbOgCU2cybboS1b9tKPyS5+CCLj9bHtCAdCApiaW
6VplueehnV6JQhU1Y+agaVUfJa5vxO1wRsklt8HBr5MtdxJlZrAWBXXakrZogNcJ
VhZLBq0RIuejJ6YXtMuruIoBXszHOK/pArxgK0HH8vLIf2Ilt/8HYkneYPfKQ5Jt
gPoR5p4vYiUVWIlpfJlwH2PTxld0UFKev7nOnOT76JoTWOtToIGDeOrSSpQLanlG
wB+CQJYVnkWvzabamagL82GHCDJTQcR+24rQQa3C+/kpdQySp9Rw/FrvPwm6mlww
5ImMV7Yh4p+76IrokvJayXhBHdcWkIKQ0MgrdU1/7L64HX4uv0IVA74ubxnE4H+a
TXkScVDhK02/Ad0Wvk+Vg+69S34vez7NPCeqnDJ+fIbCrhs+AoynAJ6e6RRpDzEU
/oQCJqXWKsCxt2F+Z5/5C4wzOKi23gIBm+694dHJPboQMO8Ads6qiRRUQxx74Qh5
4tbwjZ1VtBbmJeGrXtWNtnqMJ7BoCW/y4wkG7oV+UsVLrBHD0c/NhmT+wsZURuEz
tFfX/a+YBcdQyLLFhen6Jj1cbIVWzZZTnG3PIVXp6YrIJsLGMBth2/4sx38w0Mcw
HnwjxjO14Qr9gGilEYJWMpB/swGFQ+CPwUi20FUuze8sQOAKMuHQs2xnBI9obOOW
t+gOMttX5rQlIpUHuFLa35cXfsb5OHQnfV1ZrpLW/bpqUy59CeBi6VVj4kDEgQT8
Tk2waPlXMGhcubxE0fRHhFlcpAtxt4vl9q5QZqf4X2GgE+FmsOBEHBS8DfSen3HG
yEWwnJgB3lLL+xf65lECucAalVR0yvOWgkQSrOrYz0f8Ehrvno6xRdxyBpRECghW
hUIgSHYyYU5gNGSvWSbDrwSmPP9OCSYuYoyPNXIqwY/OZ5J8Msl+xJc8OL14pXHE
k+0V+lLpxOwA6HJxe6CjYFZDAcjbBdK3QQHZg+6HcxyYD2mauMRhRCxx81h4Nnjm
T5OSdVcnw75yXazsCj/XbIX0TQz+w/Z90bPEm+sLENuuN33k2Rm+nIHyRVMRDi7S
eQsEUIiQLfelAyKnIhCZRGBFgIuwS2I5WFzhF7+Rj0PpsT6paeXffJFHaBqsO16n
nsL+f1pIzLfUM+rOYg7Erav7tK4w4gyfmEqMh1L6nqp0pmCQwfqHdq9zB0JddZS1
z3PJ35dsTfdwbbuMdjog8brK/d7zAM7iv28b7K6ItsklqidQ0HnfNiQBjENzM9wV
Fcwt/qTc/V8bzhoAT/fYQfkXnoJ5h5y+7I4XKc0/a/sHH11SLNMUpsfCuAQahAxj
ZraUbvSpKP8GhlBQftrw5kJaPItuO+xK9lOSfgQueYq4ubIhVCQfVdmww8V9WWwv
oIxV5bQoFhGOGwWx2PVw0q8vh5mc1VVW05IEhQHPR7wcPO5PFl+a3vVFK9CEUM/p
GnRXbD7KJXJ7EfJP1VRG2a82Ny3zgFhzhV/mZ2+uF63vBQgMiLdTb1bBpMstb3Qq
iQRSvJJnVbTa9h1EPOPmXjgLla5xFBtFtIvRmW6lVOHU0DK1zfZK3N8ssmlKDBM2
+K3V6gqGGWJ7iIplW4uPtHcDEIxJ+rUG8Ic98s6349hOvDyh8x1Ww5+GFr88bgGP
Jw+rALIYP31+bl3EDCg9N+TKN8rP4hDdAdQRB4MovFN7IgtQUh1FuAD2JRWXAss/
OYUqSshWaJFmAPRjFuGb/TfcJkeEUz2Cun5bQyVMFKYrouUy3Wfb9QrAT6Emmb9h
6D033CiHVzEUhLPDSNh6402qDVpXYttTNYhr6/8uWvThYsRHLY+E6g3+gVxLYPY8
bKejCNMYAo8asTu9tZO4a+AZFzo/WSoFlAU5Ug1eCC8X17CwQaDW/XehabTKLXsn
n+jPjSCaMGMVOf2ubKzrhpfYvnbB59t+xc235buZA2DqFXmkiGI+BrAfWmSz7has
XhQ2jnwEzZj4Jyfji4bRV64ey2JeCygjQ1oQXVrlYZXHO7qFBEPOJ4njy2cvDeqi
GVjqEejtSKRiFJp9jNB6pasWu4epHehyhHsiIxOgznizt6JR9VvS6SGngVFykcz9
8QX+3L9WXSHu0k3FtWk0CZHJV49OUmCl764eWz6DJKfsi+ZtaxGU5d+/yj8nyEtZ
OIaIQb0l0kXktIE1FGCNmnZ1NDSfcoGD82U0GiO81Bz8HJVnbLkOunKfljKhYy9g
muM0t96IshvfgWqI06nnS1QViBbA+VN9aZY56zYApGVkMc33tPAyMpiIdIsNhJ5J
SxIj/Z5k4vJQuaXVfFy3X7RobXXNVvCSYPWhDmxEuIqfzIAaVQTGc4fynyidpy5E
7a5fnCVCBRokJajvm2FVafe+TpiP/FOz6EEjta2fL3krtXXatwTbGcNYNc3QREeR
clN7Zd82Os1/wiQPOMmO+IrrikRy90zuOfJWQ11Z5QdiPXzZPOZTODeWqfgc0bwb
J1N0XtHWngPZK/wQaxombie678LtxVoOYzP/t0iFQ7QgtwmRa11Z6yq8RiudeIZL
abyLWFGfWxeTDqLDXEdMBM0s8pPSzxqXk9a8s0H++3zMkG0YvipYpL2Em6kR9QDv
joJrtXOYZwDhBGSLw70XqSEGqhk4YhTiTsNThPBbaAe318BmTeCgdeTo9jCyMjVp
KMygd8AHxEeoQ/2vW1IFs1HxloiLp6l0nanGyJubmIX5u6oEtbGNM/xJz4GgQgxl
XWpj6wbkrJw8T0vl3cK5uxe5fkgHQTAhCYuUlP68zIRawhBb5PZLTP2GucJGt3Qd
GRMEFO45SOsJQC3677N6gY7AllyICSmE56f7Ak1P8sJTO/zv3Ra5nd5AF4X+REqL
AR4rldNKeNGM8G8kYqxwN6A8vADWT278Ird1FcqMQB9a6k34L55J30UxieUxppFe
4mSQSWsNdZvXDjWYeQsK2rxOj+RXrSns82LWavOkP7VSchaw+c9UlmbiJxT8fl7X
gymt7mUeWF3Mi3TdfFnbqf97ORarCyPVEM6J2cVE8J+9gR6YisFyWJUQQSW2E02Z
B8A8azVSLaI+QILMeola/uw/Mrjxoqm5Hgc9M11Rt2jqaoKtetth0JgGPRowIrLo
Kt0aFAzwiuFv959VAMPDTeLKlbu2VrsANV1hDN6BYuYv+Qp6y4CVeMs1fuuyxz/x
y7SDo/xfKGHsaBHAPUNQmGJ4G4Vp1s+MXOwKP/WK4d+Xm9VGoLvD7mjrkmIiEw/6
GDgqwBCfm5OIH4pWpD1wYzrwPOnoOaryB7bzeB6GKBzCNSFi7H0dVEQ8uwS20/Sh
HnTDgyHPAUhbkkPjR/xVCe4eiRRMI0Vm4+W0oj7W7XCkWU+ry3o9IUhuroQdjBZv
AP6AzFTy9Y7edI6gCrkfyRBjMKmHQ6q3F46ONgtilf8Zox4yjv/41TUadP+dyp8r
ZWhdS1KaiKQeUQTg6h8cvbpkSSaoyEN8SakUPvt7MgV2EDj0GL8Cujn8h5MkcEUG
nXNsWdzLVsBRcd8LJgu9+olGMQlk0kryBI5ZM7UCklIp5AKOiHzdb9iqpOgiNZ1P
7YIaD/Kb+AAOBbreHTaYr5iNXNYwfjtXDZNHpUgdTR/DZ4k8v3bO7sI4qW+HWBFQ
gdG/xlJeVFTniXdyjXzhSRoobL8/UqlBeOSrkQg1eEY+f69BxUQ6Hi8NsQVr8128
xRA+kfpYS6qaTAEmrufm4URyOyCPt4lAQpi/5fZOyAfdZ4LGvOj89xJhSmoV8Uiz
iVOnNf+M5fDXUOK71yLiaoOgmiqhpri/iyDqRc0r4UtQfJolO8EaPHsRnbwctTft
NHC/L8UplbwZ0AhLB3+WXertAducKFMl7oc3Q/TUMlqszxrOsagKoD70WXBuyIpE
p7rDgmdXO5D6rNrQwHsOtQ21BfSUI1OmY3Ta9gKkM8lzsEbEauM1qNCwUVFgkkPy
y0d/rQwRyjiUtZoG/rzRkTn20fdokycRnzOIkL4mjyZGXkpUp0bBQsdYikat60zP
Kr+FXrcCNEBlhn5Ao1zQ3mDkXADvMxWjK9PqpJ8RTs5NRUYIO4js/h7RdEVJ7RWi
pbDFeinPCwuMy6708pKzfGLymG5EBGvv0nzMhXfRm0H+FkuU3cx6tXDgZFq/gUt/
Ro7Xbs+PmkVeUcV0WrHLM9bOEjCffBYvw8ZipvDypIvXhkEl8XbxJeru+7MHGTpb
NgXSftpiuf1x245VA/9c5jf3e8zOJLs/7hmo9vOnuuhcozMj46caoZkND6S395Gc
7oYVluXFHTd9sjVozNIn9wdQJeGgXttRx8G9+qWmlQGg829+tRN6t9lHAHD3GK7S
S9/aYM1+VScl+Rwi+YMYvp4Y0Bi93vNvPfnOr8LYDnP1VG0EYTh02RdyEH2ojx5N
Do9RiyOtc0wubjOFLXRAvApdF9q1fZCpwXl8fQ37AGtl9/sE0kiWWrmIgeCpD5dr
LYfqzFz0scFrJWtTkl6NYxTxY58q5DELKuYO+hqa9LW1sheGVpfcq7f1WI74GPIl
KKLLvaArpH4i7VsV7XI7DgrCVnHLNf9K5xdU/UEWpam9U7LzNaq0rGjkXryAnl60
OhjAPprF/TRRiBe+T475QA6WVpA/iZxq3uYimEfb1uy0RCGpBMEshlMQgGyCEcKf
ymwWNtzohCVRX2Kt2Qn3pDvCI1xWsRC/XsYUAeOiXO4DloUecWaKhV3vfR2ECwZv
snlTBMCcIS/i0E947i9pwxcovTag4J4x6pSindK3qKtHe4fJvaMi0uNonyA49Byk
KdBSAhhoyQPWDKSmHt/6j0w0edLRxpAQgL8T7jLp52JTek6gaI5L9uNa4GyJS9JS
45R7g1wouOW6t2GG9KNI8N1ZdR3tEY7ZIpVGAxIPAlDRH3J2PrlRYOItQ2W9Y1+p
r+Y9+H4C1gvj0QkUQIGDGoqIpT8Ik+8ilqBVayaYGwDf/TEp6qPIrafxVl2mjior
coks8G7R1qd9KER1k+5dI5SF5NJBwO8ERP9V3LpUw1L55piYcgZ+EwrzwH7OlArK
AfqHFLrVP7JJP1vZcJnNLEzjBNUOKODcK+RtuB/6KTt9QH67mVR3T70qoa3XXRVf
zQULLeh01FzevHLmTkGXFSjVnXABg86s/REBtsJxwkBONzsZrxi2lq0c7kOF2I4L
NKBaJVamxq37MVuaqTBp0aThmpgkNQ8jG+fToQ/i2Lja92C4p6MNWJS08qFZ3pEL
zSjGrt5+s8m4mbHDdifXPoS5/eWxTBw0ezD/7GHN0Wi6UQvAG2Rfd75TnQFwGOkA
xDAvvJnZOLCZh58ynjKsEi1GrAm0yQXFxYPZldp0ATHC/impKXj88jqc89wbfE7E
BtAu5sdtiblB4kz9LrDc2EIV8RRWPphzVON3z0HPHMB43V0gF2ydnUb8rUirsota
f5ShiX6c7z0Qv8WYf4iLqPw2PAxwR6VzyCNyRPyltIPhuX2pQYLnMANbw+7ohvxb
z+gaC9b5Oqmo0H51OHacKpDsXd4XBibEHrpU4VzXujn4KJ/JyJyUIHYkwvoUYDOG
BzMBb7qDk9jK1khuzjrSShzesvE+I5v5PhnBHYsCBc9VlVzTo0CjXGrFhjDJJtHc
3DuD5StavNh6AhyRdKDJgXiV+Z8+hQdp29CXJ0mX1jE3DU8cGKWgiS9eF22CJX4B
aqQOiZlNum0lciLmmZoKXxv6TT49ShnmyjOohnGdNl9/7Tt8qb5e5MJMm3tlbjcS
dBCH5FDco+nzokRsrS4ocXLGnN/9uOcMxKmG7FAWntkPViCCETbOXj2XREXUPpW4
s/0fDq11cvmmw0Sc6/vEdUL/KbjdessvS8s+NJtSpsXqEtep2wrpJEeZatXDzDOw
rHHY2yV9jSyh0exydghOPvdop4ieYNomWgy7CEwzYiXsYvgna6jDWzweuHrSRTOq
FGfGmj1JNP8YvhvJLgmCYPTe+ELtZdxPqfww4mjZzqz5gbL8m1fYn4tk+71uh+FX
B80VHPud2+83VuNE6QM6b3cTaK5FffedLZxt57fDRbLRoLhAvy3Sp/ovryRNd23q
W12dsPNynSxqfQdET/EWkG3My1cFZ50wjkQBTGz2m+8aGYoMJqR0XfCetCJZ7bHw
KpIpwDFfoAvGxIYGIJ1rdlc03kUpMcEXK2CiGZOu/fXvZ6FOuLThiQK6LfaR00Sg
N4tkRaww9+GBdx7MDBJo7+mU9XUAkD7ijLMHXaNx6/3BtF4P/lJGqZ2wmGXWbvCN
53pd8HJpZa2bBpAfyKwutfZ1rTifk3Ixrw68q+kpB0QLHcRLD8ort0P5JOCXNsu1
KtfIwwFABlA66XaZ25YJBH2H7/kUrXtLYuvYJLXVI2z6dKfNUO/aa+vjVo38UPTF
qgLGhzeKMRHvw2lOWTWbqcmlo8sZqmfBh2qxBzAmOTgmLq0jykFAWsx4bKe6RC4h
HRIOjVokRt2PJlV/0bJfNGp9VxAPcOayQNa/HhYEzqfM/7gviwZnH7Hl4NrqVKcC
vULbmf4IkqSxSUIoemXAmDvM1j6NtLbJxHZKrOREM2gCxFoWqiIDwrUGCUMSzTYI
QdiWS34k2HyQGRZRVZ8cseDlnKJ695TUPFIWwVMfzxcn18GkrizHECKgppKifl/1
dQET+E2SuAUNNkfNSBFD3Qz79C/4BE/E8enlVcuWN9HzPYYnNWEdLA1H9uyOx61G
7OFHiAk8fFHwTJOkF6kyF7LaT+dPzLHykf36Z+tBbJlCC6pc20I2EiLmLWbKdgdW
tkNU3bW94gBtDxpNstGcXK3hQnKQiWoIBoPMA7x5O/ZpMxqYkdSvVAnhnGs+jGKZ
7skO+lNw1UJ1ASa9dqdn9T3eYm0zPzBMdiZEVgwAytCVsRNGpJuQ1CwuUiqhXZET
Dq2pjrQ0TzL0PoVfMIpo6NLfOlT9eR3zN+V6rrRM5RxNvi9JV8eVNJ+sM858OqKS
KWWbS7ZDnWesHfX68abedD2Vwlm0VuNLi/O9g1cfe9EqnK7CYjQTogHWqfow9KgS
G6sCUi+moqj+LE10tXCnGtMnZCUqs8RVYpqL7iUSbz0CKjoKrE6owqNG9admJNOZ
B4uza9hN65ZAgQGmGYxk7XDA+Gdii6rxpNyA3aA3dF/dAgKdKvriL+XeY/wjrOtg
NNrPTVf56OcSlYDzDTER/NRfiFJWMv3kuDSjBsj69WnT64dqyfsHwAZe6IhMs891
LtZ0zS0d1oSIi4hpJY14+TXeYcAF27F50MADGQ1zQMqKFuGsacro+oHoHzYdr6QF
TmFCZmO3JH+IzIHwIZSefp4/eHOTrLI0h5Y0QLbggCggg9L/ulgAWI/fClqqk/3M
6w7zDnj5Z4sfH+xKvOsAYMdDyOKHR3zyAPE7V9MvGYcJLwKEvwDNP/AA0J/xCsw8
9dTSIhqAnLyM29kn9FB8wopVNCYVblQx0S15WQ7PN4e0Eqj57lDBg30ocu3XiHVz
cgxCgWod0TjxZkg9GQ63kj9UXh54XEGo2F8z4FCamWUmkny8gqjISO2i13o5+/qE
g7LT7z74oEA0+2k4HpcJ1G4jPd0O143IWoVog0FvuqoTY8Wiw+f3IyhMrh1JIcsw
eANSx2+qmeh2txr59POLXfPCPGT/9VSQfRHNVkXQodQCJssAXWp8TDFEk7oY1ptt
GlC4m5BcSr15Qf9Fid2qotQHzJhZu/ldo7E0p3yXjN9pOzI7sm+dywq6bp2MZ4+l
HE4sxlKVGPbIx4djJP2jCyIn8j1yXUq+eCuQsXrRhlS59L87nthePS78ax6FpdoR
fuzUZCl4gx3fXXRHvPXQWj+nd1NT9SgxU8geiBS136wugucRdTG+6IBt44gzpzKb
mz9OP/5DG+xRL7GW94ju7gvMhpLz1dXdwkg67BvpyrNr/usE5QSI5Yz2jGW+Uxub
MEgvNzM65BLgAjGbGV9LLRnSMHir2q4+lyATwBCqubAyLgdcFrIjcDEb1+l4YEEc
DfKs+0V67G0Q7cmaUCQqf1zmXCy377PlHtQtPiqEsU9mIq/uP5vY/8WaQidEQNMU
T6Hhjb/dI1H+B4orJewqt9g1UchuQ8ICgVyK+1JVeWY3Aniot9cn7FZNllnxDq/Z
lChBa1aOHuhfuYzltPaWqhP8Wk/ctIQz31mZFbsJ21v1hqbExXr+Mfq4McXzjk2F
usEA1gWMXSEkRvrdVliYqObMGHmtpFSgf3FYmO0CRVcveI8AvXW+QPoDpiO4vWmM
b1w3K5SnSufseJ4W0DZd681JOu4oh1pUcjVrxOPt9a7DeoxpEg9+0fFCdAK9HZs6
nXnnYvkvRKOzWcOyLH+9YfRpOey+I7sxg0f5suW9NvoWcqtvl8lfUCGV9ht2YVV2
fU1sFeeFcn9MYsCx1AEfPn6jXLa/51ett0qdGJtFNIFlhw97/W36xBrA7p4vFuIw
71MRr0/byKsvCnbgq/MvMUlbJJAx0MNVAh/W1doHnSlOMqdQBz+/CwHNKJMZ2Nt5
aROpTbuSaO8eCWe8ncMifEdChbbJF/G8cqzQGpM0X6k+KZGykPH1EpuybrE71lNm
5gTVZorfmzBX81J8ng5UmbFR5FJfEODStXxeMHHiHKPCgV7th368xIIpRx+4OGYp
MY91A7ml6M+eua6WwHml8RF8dV9mWgDRvnf8xduaaH+OQBC6/5hOxeRHkzS0cHPo
9e2JPE7ih2Vrf2f97zcsxOYdRsjG9qHCTrCtlsBafgiqok2xQwzloeiiVYgUHi1F
vnk0H3dUpo7SDrX9EAk/PMOeNlbC4Hil1zBe577oBure9Pd13aZS2le+5vG66Quk
tOnXr/YXqk02k4xr+YtaoBh40Sul4iPg/Mt/ianf+NhUH3TKqXdL3Tjg50MyoeZM
Oz2e+I+Ew8GIEw0KFF1CFm51qd7Y7N1FdUoXjsik7BJ+7YC8YPUq5Rp7ZVy2x1kM
GsNDNlhf2xjeGvSD0ipvJQeHiQ60uhEM8X+34htJyMLLQufrqujLNmpMs/POI5md
X1vzoC6CiUUusPTLRGP5vtIdelynetZsQ3HWQ62oweKFuRsrA2C4qWzmdzZtndKr
CdupqOkD/N0aZ4MiKRLTIhg2aUDO2SYir2+N2RMLzHsz0VPHcyHWHUp7lqXyOgYS
LDlOYXLzHpH8rSEEX2vxCjzJZ/JxU2/msQhJuR2B7CcQDvywGqvMfsl3xjPC8Jgz
OodUUVbHvwRiHNE29BQsO/LuEUarhfMUp2lYZrcbTfVUfVEF3htcTVfss6TRBGDP
DX7Ok5a0HQ826lGWYkF5GSqBMJBdATi4+1jFkHwFij51i95HUD0iISCpoDw3ZYkA
Wubj/OBqVAlQZ7umfQgKpb0xArzaoOdRBh9MeB5j/0Up2KxHiRrKAm+p2tS5pG/O
hG7IoYolsiotXYdDn8MIzjed/JW6HaJ04h1zh4m0lxBztQygRvkj+86K/mA8FMmx
hKaEYdtM2sOZsaNIOSxZxkPbnTdN3lAc5atUBSBYtTXSxSaDSwGKM1UtIYUIkJTB
q5oRNptGCzw0f6YPuDL5HLGfvZZpjQh/ytxdHnximb/fXQgBKMFBM1VrxWqn4PYs
fkwFbgOfrDKccPqnm8hvj4YQ1AfdrzAeAylgzgLdJpUVbwLS2am63GajumyuwmJ4
dQeG1zBAv8dbXBcMrRUNyXomGo0Y4fe+EBKWfVTFuH8c6dYy7FCxVcsG5zIPQNTc
olAbt+3n85VooNhwiF6n5XqDox6obL5v2kMcCQmDDGrTIY0hyhs8Vn8ai3+1iXBP
Dhl4MH8dafKzF9J67maP5Q+sRkGIr9jWJOX+oo05b4K5vSAmKltAOOHrE7wUtjJJ
kD+vsrS/4+EOOnWIUOeFnW6XDnOh2pM4R+xpoVrYd/c0w46KLtKv3nL43w/ZYPDT
c7T3BAu81cUJwSwnvkHaXW2idiYlzqeFBI3FltzlgWk8NaPx4+4AXSudnK9Afwlh
tAw0Dy7GiPb0zwciaXb1lWl7mlui/w3rMKjqhKqQYnfk3pOLDaJwKh316DaXZ2/A
dMB3rWtbsSOhrGM90WjATfxab/LDsmX5/+54Fs6aB4dy9XVMVad55WtopryXeYUG
SiLLaz8wSGgPB0UlAPOOM3R3st9Bh7N67mTH66KAuk4QRLiFqjBbLTSuYac11JbG
fKMQV9Oy47oFxL2XfQyBB0prUkcHGaOI+Sa6vKQeQt0Szw6z07HK9lVfo+pInQ5q
7Vbe94Ah7MB/tUyCn/yHb9Yr7a/mh7ihCvDADLuHcILUOkAcofYXqWQVb21Neu1t
zfNZ1PFTC2qx5nhRZ+a1dSPflfJfL7RBVc94oKXdYsYLKj/ZqNCVeGPG5vz3ISn6
cNllysjoHOjGzfotMehiH232XKEYmNjyyLtkUYcMjcL6mDbRlJTcrpmwl6kXZdFh
GQY10jP7IceLECFZTX1fcdxl1AoeVGOlo4xozwhKpPI7Ln4pitmhNLRkvm/thPvr
GVkiSeAzKOLVixsk5Q6sTwRscYn4SjVRbS2yeApKs4U+S5OMiYX1+EJ4a97Ca6LQ
P2BQfuSDIQgooNN+pIYp0Paqz8Jix5ywc3NOTh26x17YXSfgbCgI4DOSaloEBqlU
nytiPHc/aJXvI4/9tqYGRXBq6YFVxkKsT9t1xozDkgvCrJzim+Vn5IfILGuP3CgJ
Y7JUGxi/97H1IQbdBn3PZrqxD7cgr55mmzo+V2H+2yqgC+LrhNRc4XrZNh46TtIs
uTYbRnnNUVaDs6NGZUSJJZCzKt+UK9dNR9d+ylWxijgYWHosBkCC7AFA7GFwGc6W
yU1LwY+3l1pnIY4TON8Z5wWAJXX/HUYMmJQo6f0isZMVIbZfZvxiyotRGQIoYJ4e
3GKsFDFLvVsx0bZrJcgiUg8CYFc60QLQTTBbBwO+1iYtcfHjRPezS9fdPN5Bqxv3
rzd4DOoXiQef/HWox6LW1ks1g++NYohiREUgE4RHS6lD9MDNuNVcaUur58pyAGCb
Nlqqj4+TbhSz272mTmMzN7vZ5X3gO6tIJF+7A6giK9WPEx/x2mVXIgHuUJrRHBZq
/pztL0W+PehlUfowvpPkbhQt5MfFon/d5ONwtAjb6xzihQpjEEZw1RvcmTxNQCHZ
k1T0T1JabGT+Wp4qJi9Pr4xGae8MbruBHqHINSa8bz/jDv+KR0RdbgVf95SC4mEw
RqjSj+hZ32ssAh8DCrH91Cf8p2B09itrBPrMMg3MwTntR4uKdwhtIFZgwAhRrlNb
1nFm0Vn8/qJ5B28Kd6VVHdKLaDjF0jGjB+sVnsqHxazZyqKNuTx2SONDebCVAEWx
deCf47oGXTiBnwyuDBDzlxwkI4Xp7XuMWVqGSK1NBlTAH071mZ2jb8Iv0ohYKXJq
OwVrMGzRuF2WUHPUrmnyJaAxPb8qbwVAq24XuQMW2tBEZKgQoHr2aE7TXU74v6bC
ebs/HChmFphxnCDxU44mx54TUXF7xOKbEaZK+NPbikX7hCEfSPxEOV5veR5Xf6Ag
uuqsTo0uf8+jwsbxhQjj+mGvGOO3R5rgauR1gVWA2PrPZrncjBAfjPTCNg8kBePz
nDWmWmD1/Jkgk9NKBIOQKXIbClJbhI8mIQECcTsHai7azwwzbynr8K9zQsxOpj/3
5wANUhW4TNyJH9FxEQDvWqjhhlEPC6lu6i8eUkSNnVdKuAzlq4hQu/Gm/ZsgvcNB
P3HNjJhqwkIxi6FNNpOZNNvXOQYvxZ/76u88/xdyQfTFcAvWGY+32CsyzV7J+mMX
8N9ii6uzFGdWTzJLUbTP4Z5KlC1YefT/xhNXWlyHHjKCS644Rzmi7BqbvOUjIN/f
8Ob1wsKUUUoDGX7+9SmSXX+sA6bQ9gDc9bQma9QORARSEc1ftsBJBk1jrrNpKXOF
WEdsUgi0oEWRaoK4VlX/Y7s/w2IIeGFlM9WaWoiWbRR7RhqB7bDnc7WUm7LEnTck
aMK+6jFOm3cTcER7iWGU7LUuxLeyFaEufLQ7cTeWTyUU621fqHkhtDErtMzMe7t0
6+msfp/58ejgqPxo35J9zQnVsr1ivFcNkG9rbv4XgGdtYcld4GfsRXY0yvKdROsO
I8AVKfa2eqxeYOwGhVqC29+m2jvXQZfFp5xmt+1Vh/VBuox4tF8KC+CBu25jaeeJ
xBx9U/e9LE+xhcWNTlr4gbfo4rGKLvZts35BvR7/+KH5vdgGSgeIJtipEditvJQC
Crt4NQ+KIfQWiGdStu5jeT5jMs5py3B7l4nL7q8VMmRPa47aTYIDSQhUItWBCKLE
mrZdyYCcSDqbFijf0hKFSRadMuHRcKyRuyH7ag6y5iOloRqjk0dVcehKj3lrbjM+
vkTn5oMozNHWkhsbYGNtLXeqTKwH8wTOVnedvs3198VVy+qaLCbCRagk1mYz6JDV
6W4MNFhWqKHqvy1g6+rkVyhhAeCfaLlSpbCEJxGVeEcn9DYXcVpislv4kXRsgT0E
tnL2+cQLb3NaiYKc9+0IMN/iMsSFUtNa2HbCSpp0Cg8800GUcarPjVJpFQepWswU
5+RKfyvdQrZeDtXr7JNxm0YCqdRTsHfkegE549rNAHjCAhEcTUfzuSZsQWp2FXqJ
5oA2ewH3Amn2rIpCHjNAbucMF8nnPoqapKKF8SCuDHqyMkzQrTajLGonzM67Vrio
JotfomdRrxaR418hsQE00PXW5V+ncHFh7Vvp8CY96QsJvQxuyXmuJUM8VcHfu8lX
BYSFlXtfT7SpQJ+36TV2MRzuMWFELE4AKb9jL6TV9gQ6RhmuNbh7oo96MQr0gv4k
D+pX1BA+UoIwlRk+MTFs5PgJ8KCIs9wV7URqhJ6w3KJtYAufF5DO+qHVBiko5Tx7
jrNY2LlkNsxTh4QGSfZ2YpLnk1iPCIIjd9xRz8guNXDjBMBb0BtcHu1NvNUZQ8FP
6Ogl+8c+pVK5mMpQSEVbnPifo7CJFhHrEAYrCIWsjRciM1Ukx8ME2qZqBwI5JOvs
9xUsio+5pPnsnXDuIyblTVakBTT5+FRtrfIyiNaU0ZU2OLcJPeMcr1u22JSdTYXb
/xKP7d8S5jTY3/nmUGh0kZEBgYqbsTe8PmZv2CGtgBb7LVkA2i/BtsQjfaOzekOL
+FU3Y0G+uKzFI+C4f35aX6GzI48mLvgFq9kw7pZuazoG86WMcLC0v9MpDLPmmg2Z
XpU+lOKDqF+jn/alX2oJnviLx59BgkhHx1YhYJ7UnBrkJzGaQUs9yDb8iFdePU2g
t8g7UKdg8hspqAJ0aDPN+PzgHQLxWnwVCNyckiq8Izu4yICQuti9JtAsTgd6WjYT
pbkdH/n3Mr3gjFvhydbDMxuRKPXwNLnuTL3w7gWfdBC3wcGDocNaKoZkReprwluW
0GApjVlDnIQrLF0PQCB0JSLg4fsOHai1abfoKEPD3m7ThTLbjgtYoN4/tuzmk5K7
qkXC5n7JXutavzJchBZg9DCn5zzI19z0UB5BuJW4FfkVJFBASV2m0+hwHkVXCo0F
F4CEoJ9Q0VN7CVnpaz/CFTNPbDzX8xzORQhIDcuZZ6OyNgER2AfVboSezgYokJir
v9SgSj6CFZ0jZMF86D9zyUc86i10KXbut2qPccUKU23meM401otY3H2fTdLBf/bP
KVUF7dLjWtQUopn5afEXr/xhdAW4YN/oWsOARi0HZ2THZjS+q9eZYSveXUNDAbBc
8xo5KujEHKDldw1XxQsn7PgrlBFbUiRdMp59KcBqnyFsDs7me68tPVFw5osvTZxx
YNmJl5Qh2Gc8UN+PmcRKFhVQhFicrQj8PrcvdX7emCXKGvxhAYgWJHdLENza3ha0
e9+hFG/2ApVdpAPzHh5UHEdEsSfdHG/udZGANh4c1m/BGG1ftTmF58W7M0sijCDM
dfInwZ4CawMgh9FIZF1NSfjLhDdKHwmN73hiBJ3tBinvzasoeLz6PjYcdwUt5ffH
O7Fumk+4wj/f3PQeopHiMWG4aQm0vls6xC95vfQSdSh1DU5JZP5CTs5p7wWWPJOt
odMgh1vqNguHWblAd7Zu7sCAVkp0pHJ11g9hE5ds/De3c3wgSctxL5k9QdMHAE+L
HQSv6ZB1PTAF8wv6vnaRhQe2FltwGaF7QWfnQR09zpY868dRswOeWpvDeioIkmaG
VcUxsRL+UUfVhGjtkNEepxLVWfzj+QZUIwmvvYW/iUAhLiGrkKDf2vr5Zt+6mhRF
y6kV0ljPHMGRsX0aWcmfnh30VH0JxR35A4CpLG3p0r/IfEJb0vFLxIP6jyQ2Gf2r
zGquc88bbxp0ebAukF+a9an3c+20AjOhwlAA/XudKUSAVqxf2+os/FOKP80uoQES
cl20qdadW6yOixQs1RfO7fSUvT2pbtj2tbexaCIybnZHK/huQfbO0hxpdcbexfrY
sWvTCU46GvX3oBTdrugzFfdbSjvWbTh67SDfGit5lGQJzjBdGNPHy+S7jJoZjvh6
KFG+jF1ANqfSjhPlH8cAE90g+uCeJ1/N16jar0fpXPWjd0ldmlSSodUXt09MU3U/
RZZMgEAoeDqm55fGVGuLAMpMNdVexr8ABY3NHth76cCdxoICzH1sEpCu8O0t+T42
1a8TbDhuMZkem2n6RuS8I0Xm9QOoc88tcNCbl9Dl/lF7pAY//GCl3m0T2TwDrrBu
DZNiDHkAL6xs+k/YvYq9fn3TbZgTJ0PB74JRFLHZSRkE/2i++QS0SazTAPgQ9E4R
JMCQ64Ma3KNfPkyKxUaV4LvXUtZKfDdmjsuOgCmgI2+oyzmP6Ms8tpkQKJkHv3r2
z9+FKTYcM6R5P4RZ1c7mZ/UK4qnghQJw258lY9XUUOMyC+rrSvQkafjX0nHyE+9b
rJzJc4B+/z5v+M51j4hsA25NLARrq9yRHVywgD6MsGrjN0CVjXYU21616WPxW9ZV
CUCQbjf5tuiqfq/ls3MmpiUb/h7uOfY1O/o4TrcvA3goDm3e0IXeaFKkBfmnw/6P
aWeRJE3sEYfyPdG5IbF9hgNYywI3XqXDwsSgQyyJwFGpYh1YelDu6Pip/DplmWva
c6FHKpvOjX70LQf3z/Undb7fYOBcWYAR1O5CFCYWzFPNKOjllkYI8uKQ7tKxx0GC
gsuM2sbbHDeJlpy2A7WGpy2tnJbeUPHyl+YG7rmSjZDFjNWH3uI5DAOUkBTd9bJb
Sf+hQ2yR5OrhckPRAiY8R8lyTFTFdc5zEqo+qnqysvdt5tN5mj9PI0YzYW+eXvQy
YZptT9+QT9PtibJbRxUfK8y2gYaG2X8QjXYyC9wUFW8EcILrSXdAgohiWOA3lt/K
nSAlh7KM/DvDsClnTJUhuISkE1hO8QcvytYOpABQcmK4N2vTRxLt9KJ8NxlP6oUg
LHbbxQvOACwbUGLX7twia1bPI2W+8jS+wbfSDiZp8O5Tq2aVnSN8PLseTWWp+ptF
k6QfV1sREbUfJX2p5TJkVS41DWQgF9oSQyFV10hDjqfODFajmwd25p54FSEL2zjR
+i8V3M1mvLcC7tQW+BrpR+eevyILve8oTaB5v9aL9rDadM277v7QTgMn7pjajRGQ
oO/9xQm1v3hAk6aXeV/Lx23GeDF7tYv3c4kWEjXoz59Z5wuGZQKJ25lV3H9L/pT6
aH6IYVBIzIUZzOnaucyvwH6k9VKMEE5IuKn3kgfWF0rRNsgDIWxNztUSZHVxkxyn
CbD8KMyG02csuDEesqNRkkn1fPI5NrWTd8zr5/RmE+RvG4sGRjVMUVCRxHyq7/W4
BwMBLujEyi+Is9AlCe1cCaB+IdmNUjJIX4+I8TP8guK59A5/7oyg7HC6O8ZoTGOr
ceDIqev14e3LE7KCkEfly8VMrH56QC7onybuYpw7x2btsVXx+tJAZ2yNYr3A1WZ+
hnKz6zWmXdJtUcKfeWjnWdS9+TiMSKbpK3SKtzRYrTbygnLynu+xtBa9PXzisMJU
aFS7q4OvmpK/z+pBrMiomhaQ0vZJoRqzRnjQQ9Ck4QVyxaJfRRQusVRTWnJAlcyj
DBD5eiKpqi4UKthSRmTqwEQTBBgDPexKfhXPv2MB8r/vd8BmXuswuXQQdqYT9kf5
zZApV9MaLzLFFjBDk6bf/YNKIzsm92DRTmSYgYH+UguXdo9ccudjcXgOd+P/tKHV
/r6tP/0oFQNeJpld5IuQxdj02EYIeoLnbbpXUPtBKiAtzPEKa56OaHsymvGAMADO
vZ8d8WtfPLDUosuSHebk7AVSiHdwsLmCGMTE+ShpjGtrA1tITKlbLeW8LmThxIjk
Ogv+Sa17kxH57lARy6uKISd+5BbrbSMEhzHDaLPePNSb0v1fxsOQ8wWLa3ydiZb2
+rkHTvMJj0qt+Oo7fMenBp1IezPVrpHt71CoOOGdP7P6/mN1wdCOpMAGZoR+pi0O
9Kv8HD35ZTA1GbdhnrTEAYfa5l2qL5IhJYcHEQOrGuSHM4MVWUpVlROF8dKTzBla
I876UPU13Lkq4qYABcIy5OgRyM8jic86gLs0WonWaO1z6CVpJLQt2HVHLe3bB86H
10Hd5Q/9WQWdPJA+GvNdoHelRY6g3RD2ehBCvdxCtcb6mT1sQx84CsFSpxdd9izT
0VsezBd/f+Sen6weoPFJVUmEzQAUmwZdPmhHCBwZeg2rzU8HVnc5OI4lBi69dJJ7
pZqhR+O2YQJcAxcyg6K9YOjMsoKyrIiMDCz4PJFsMpmVTUR7fx6DB2C30mn/wQA0
rYbczZ8YsggWQlSWJGSC68b9Or6iTPZXI3QmjwZddTGm3DqVYbSwb8Br1amRRGFw
3rGmErRHLH6ZrINbt6floqrs3pEd83ap0v7hka+GE0f8I1TP76JZOfHiUyvVTtnX
1aCE2Hem0hvLNEC+YQ4O1o6CrNbaVS5urrgrORCFg4Al/jV+1lWRCShwwB+YzG9Q
YpymI3G8zhSBZ5lX5gkPCEbSlCMpfNKn8+bsSkTV3Ls6lVpmq7Vm13YGbehcWnps
DXBbytcwBDdBSn8Y6aWM9MUDWA3/JKXq60egfXLAVf6SJs/uTEMIr/b3JZ742Ly2
dq/1m0N7HdPWQTMhgQZUxuNdCoIGwiXszi757bUnedIsAUvjqXlNHn6Frr6xIR3A
rUKbtQOMbHcFZfa8VtfaEwk5DUyY7BktrmC4EazNyUG/6Hfj0P9TkLPITQ7KFjig
Hdf0/ottiH4bknVkK5WGRN/Yb057UjMXgFAg72C6q+on4FjvaUjk587gRIeTZ2Vq
/UDnv02IwFSBAsqLv8XsiEwV5BXROs/w5+DlnJjpFrWZl5MWpBWO5k89ypd1sU7i
nucldpYSnKGZopC3JVNdwNFm4Fk4QA9gzChbhiCy72V7vQ2ubFSLLRhFYEXSrGkm
ysApglHjmPnpSPq/x3Dgei8OaT+CjY7WFbiPM3l6C0EMwCan1jJaQIyTeEZ5MuGQ
ck2mACzyXjMeWXapOlQbAeFAjgRSFILEFQDV54BuvMhAAhLbPByrztNV9IMqXpZx
/AwKFQfuyZHli1LDSmkXnV4kxm8AU2/OQv6akzPyUzzaWXeImgTKLBC4O+BIv+3y
ZRwWfSu3FgFQletn5qJze1adh29Lw2GY/H9Eh+jr7iWNmMXk0nAtGVP0kOUmBlP1
cb/36Rppz9y9g4hzfKpSS1aiad8bOeMZSFKWom45vFkpTpEqJQB0Lvqtp/pwUMxm
G/u3XSfXowIZ4WOC5pSxAMQGm6VqTH/ChUlWHUxCUUa15RBN9Ph7zrn0kQuDjBV7
mxzLSxWd7Iv3M7lB33mw00XUM8x+Tn8rzapcX0IPkybbLlv/omcZozaqb/fLu6zQ
zfEYq71y8Ff/grkArZUL6pamQF3XRH/tjkAg8AObVethWQdUrMpicLUvhMAwIM/K
akVz4NmCBs/bawCtRNWwLmZawm7WqZb1U7h0H5uiCf3O+9+F27Wc8jdFO0sYnDWA
bLC+/3GE3+U6vkJGCsCzgbGBPTQGKdqR9nnmCdF8c7923KNHR+I0cStURuYL+rDt
UpM3g5QIcCn2GajwsUfU/h2gDw13bkTDyAvWkJUMBt5y2S8n4EXkgabEf9ulfsjO
RB8TW7Lt5YtKJyjavjWlbytxLiazgoAWFtacsrBLf3eOZd063DjiDFF8/hR3aKNo
LIve/BKnJkl+Y6cE+rUNgx9hxUi2nHDFd/Vs88yZYVOIUez351XeyTtxxLUVVs9S
zif8pnetN2Y/x8mIn2qF0nlnvk4LUENjygKpug5NFsrsr8i2KcbKt3a67K7waN0Z
fDlwVFQ3S1qld7T8RsKkj4GyR+m5u/UwmTp9bDxEvgP3852SfGt1z3UceXwc6Kis
xKqc+evBADsW5pTYL/vn7hqttq23fEQf5GN7WcotPFjIGvqlM9mBjSKuIALvnJLE
1bR0toPPdHGDKz4QBCzWYuOjpNmqkLVjWfZJA6fG7Nc/r2/iYsdZuWx9tySgRsWw
yAlv/BrvsQUPqN7qxrCzBAW28Brq/T728DZqUCTlqrk4kNgV4a5RHdfsPpvWVBNB
J6dhKJo8Xk/wYFzgQNEL/RnIDIYF4eHE+I8xv78VcD9jwhSjYVgyW0uFXdKmd1XO
I+Oi1GIB7g1weOD6qZjPM3duWayiEAijFh2V04GOz472VkzzE1RdhPxpRhfXLFGg
swRoJykMt1t9Dg6ubUtFebmqkb3BmggN4Et03TYxUkfsXpB/PKE9bLzxNvoKPtOJ
VvE6ETEt/tBtRy06juekk+3PZGYXHC5q9umSzKsnJpLkUZe6LXwbLBiz4p8CxJLQ
mlg+PBw+TSugvCQFTRSW3pP3tA4XKFAy5aZbDheKN1HgT3rlb4g8kgP0U0T4jSIG
9o6eAyU+vvxXRR60DVxkxS+FvkXROXzCLnpB6ax+oQ2t3GXAPxapnlJoUXPql5Qm
Vas4qmiOYiUevbypsOuM7XndH/uyu9ddOi7kIdLgUsqKka8nlxuvUT7fX6VlyYlU
8eWGAzKkxrZrVhJO1J7OZfPFOKRNJGPJKuMLIJxhNKnJOI3Vgtjs23R5qkGV3d88
JzsD1Gb8IUeDI71TzloChVSnDdPjXiNTzO/RjTx2ckFK0GX8HLFUUSgKNA5taCC7
oye5IgW1uYtukh/ti48UsCkixMMBj3dASwVkLoDBaXdvCDyPrtoarJwL02s//NsC
AX/W+d7bmLzQlSJZxavbgkBWlXCj8pZAAypW0Y5OBx/KRH56JI3d82anaK5V4mvo
dTnZkrRgM3zikEgkhX3jG2eUWDZQN6GSWXKwceccUnRap1hCKKMU+/dxJf0nqgTD
iXx1tYfjlBWuCY4KFjYbQGxmbqge3/bJHiWBiHgZPSXZhKjmSCtEVf1XNLvVeEII
VMbidIppddw8az+EUm3n9P6KLZhLcZPl21QSN2YxgAYhlbbWC0GTMN2n/eK0xPnz
f6Vxy+swu7Jl9xUWiLPAnnghAJSMWTXVnwCdFpDKt59PGb9ikIeADsEkUW4UtIME
RR6rmdAk7SxefzbDKigLn3apr87D73/dEop+QuNILM7+iF18si15Udg6iQgW6X18
ifsxDesCfGPpiCoZzGvw+Phzp4/I3sYANpfHlp5bPeOSo9QNRiOv0ffYlkW3TRIl
OpovqYPiJwlwCiFyyzzWXzOsl9QgIkHE2USeRIQm15h0TmK0QzmLXVpjailN18uk
z33lDLlSfVLwSAhfcXSPKtgrAo9tZdqevTtyBUHeCcmCP5p/Mj3v3h+s8OrLf1BG
kT+Z9r/CKo6Q6YpLc1xSSxfuP9IPXgmjselkE0JQzjnQN6cjo6c+fUMmYicQdQ+D
ImIbpLfriKkoyuDqMj2lhFvnKFFbsPtY2QFh9DQCBiB6nZL/B5CBD3YAsUvBsQNw
hDIlcNff9GK2fw27BFJfjWHhoHpZMVj+Vu3EFQ8FG1ETY2zQaP5PBUX4yJ5+im2Y
7xV/7nb2LzMG32dj0Dowppwhm/HZpjj3dUYhpoMqA1brU0NFLq8NhKfmKca4zkJ9
VsmUs0dwFHDNwTsxJ0zeI/sB9HNxIuwfJ+XUuGZk7nqkIgxGsJP7++JN5wJ2OSzw
ajKa3Qhm6QkNDw2+ikR9hqi8utfDXwkERFS3YLNRL99G15Lmj1FKSow6ETOnr8EO
hRWUmUkZjZtS2APT2eOkhW74J+DBo44DaL2L3men23plM910gOisRHPhBtqRqWFQ
pcj3mYcVilK1z3JTgDtAcAxnpoJ2gbi96bMLafWG18CKROoX6zrcUqYdBYPSAt7y
hborVNB7Fhs3ukClfZk/oUo484QkqGKA9K9LdVJ8t4KF/wKua2ZevNzFRefyoLHO
yvERfFcMkS4/et9Al/LCJrdagsqtJDI1a6Vey4/3OY6xs5NxiWcQ/ibXGYjBrjzP
7r0pgqCoVdhvxQERUTlZ+FbzP6Vi7T71HYHm0FMOYdSi7Rn++pSSxgUpf0NmIWmW
HqxvH36qqY+J2CgCK6XUhM9BnFVB1iK+t6qaASIEI8/RvbZFK2txNwGjUv76ljfS
2XO9WvwcoAjY3z581UhK61HumsiFOCnoq0YuJT4uJG/NToieaLgirLF+5cGYv6JA
sjCIqBEYU07sO6mbtEN9Ztme9jLJZkrQGF4im4jywQJdt2Hu+bXyV8+wp2DLlCPg
wjAB8nu/wHVasVUxpi/IoDTgC55H8CNxnO2TdOuSFSaDNyeeWLsmobMCTbq+dgup
6WaKaKXbgSbH8FaVWCNFcK70RvQnXptxCkyf56h9oymIzqgt5o3ZVKiron0GQFTp
gf4+XjqFIPJbKFla+fECNRzgiKlOdAgj3vLSL3bwFbM97SzIpPmoh0jKXauCZF4F
PDE/wbZlDfeIOUe3uX8KwZNmiwhOWRDv8r75YUrJfgnsvJuT/pH6s3I0KxrXPK0B
SatcV7GpQsPbYNJyH6mq9z9u9T4ujZpK5aMjMRHxRmGwUySt4UDl4ACvdnaLYrgV
TBuEEVM5VW8xUlFKdBw71slAvZrrCVImlGAVYbd7VXuVj6cSlmHvAoAjOrxkWjWM
mPRyrL19lmDRQp3e2telvQy0wQOLgUhdnGePL68tgx2XK94B3R3IgbrMRU7P04ar
XBcGd1x49cdYZ5xFAtIKw0SSpIVripsVRpk69AEqMR+oh8kiH1vHLUZ1lPJI500d
5hBwlILPy5xdFUofBcv1aV/TgtxTZ32kURSDsMSqosBxXzWcKpfZqR5cfPFVTDNq
HRrHGxazpr3zqPf4yLFb9QDsjjkd/vxGbY6c8JNm/ZmnudzxdHOnY2qInk+E72x7
ok/9BhnR0gPhMsvLIRAL8NJqBtbAv+S6s0phw36YL4kktGxmXPepprCLztWdTL8U
cTm2Wm5yahBdrZZbU76Cgo9csDmX46yc/jHXr5Gf66bD0RHp4E/YRuwczcfeTpzS
V/vM6qTqZUZN2vqAQ/EB4qDSx9MPICyn9MbkkxBXR175vbYspVKOKPM2iVba/Ugo
/LX7lZDSANE1GDe6TxiqTkK/2XtRyZzg+O/uZ386rUvb1PngmKpbS09HXJqBb7Pl
fVAxHkf2dCVOGfktvDmZtmGOBF9chQ7bJiFSDSNBYnmeLVW2PpWmltq5kVXO3wvP
B5Enad89x7tbDGr6Vb9RDNe+ZFTRdxDifdsSyxIJcpFWun7GilNrQh+/zJv8ak2+
eritdvQU/l0bwz9QVP9CNxTMp/XItCuUpoG06ZNRzojC6ZMf6WjboADJM7raFtyx
oDleVxbysfFXnzXovguTYPZeWXeWIwvAWLvqS3bqOldvN7Vk/b2yNIWwKjhA0jxl
CttufmF+GBJo4F8AezCCZm3xrx+kf810SX8FhAaBP0T0LK0cV1kMf5WbrrEMu0MG
Ky/tXKuiqch7XuxAl/k66FY4dX549uKOt+zPfI80DcW3YMRu1I3qBGPK8VsTz3Pl
kcvJU/9s/Gn1cuDkBxij/05lDFvSB3qNxLXXgH8lK9SDDMWjejXCME8oWo8a2/8J
O7zpfx+ZZOC7g7DgREXOG/7WWHH4tgkv+5ZPiTV6oXr4i5IhsCMWypbCREPFglhN
8y0S+j2X6p88XNxKEtQYjDan4XVyz45X3N//N5XSJSKN0Pt8SqMpgX97SuMG8VwP
IsTGQgUEWvA86AKC6k8e4I5McR0pALK31fhbwWipR4cGENVQLXf5CCGtABr5B4Ty
E7eqZ0TCrUPINskwmb/+vXQqOiRTo1WwxyYVkQWvx+POioDHeH5V/4POxxW1m5p5
8MmY+TyU3E6zKeye1r6Scq5DRb6Bjn7BPcaYPk+wu0L+ve/128xQMYhO9RZKffyc
z3z7VRpltJZZLMABfZmcV4GdWixHIHoHFTbl+RvAt1xlwlRcaF61/guBJQzKFomq
8QRguP5Nij0zWpn/xc5x40kbBVNOYffjVZwzU1xdNfraGSENe/jHSvbbGOigpFgg
Oc3ovih73msIkZ0HMVTMxlMnqFMPKiZ5rXyECgcWXgWQFBbe0Ig2uotcKyOewIfb
RH6KCs59mhvktHehZsZm+/IVUkVbQxH3Typ00Y4HYGZOyiNeKFfBTo84z/CdQbtC
ohTmvp1eFWLWdNKiWhrYkd2h9hwQ8Ly1SJ0PZMFl8+6x20nutYJgIY5dFB85YY0x
oKQXLzRdLkhTgsNaWYGAMLu9ox103oVDCdQL/lShrw0tRg+WfIFJzA9KhyZduC5i
Vxpo4NEebD1P3kWowpLGrO2hkizXBQdAMg8hs7CxVLLCCAPXb0ZDbCdMwGTTVQPD
0/Oe9teqYlhblWPMkuNsvz2JNXx2PyTxoafq7qk9HRFvWY/UDXtnUUzn1TcXOfgj
xxZgSY+3LOYuhnRuDLNKz6NTMEGtusKBdQqLy1S82EoR7HDdf/LkmIUSKN5yWevS
Oh/nv8bh8ckBag57KTHO6gvBua5h+F82dkqBck4BDsL/W6CjSvMnjQlxXmCgCX7I
4+zZn2w9vM9SPZgivhANDncYv0/2I3RUc5ML3bzDrwLp2ml8fpZTqfUz2lYLMbYD
6sHDbAr/ZBpz1vCzOB4YlfTXK9cRtagHCrYOI4VRL9pzT6Y2OTlydFiYWnAoOfPl
2dDjzdhw03yQDQOilR9pbCLdi+cRlIXFRf+E+NH47mIXCZ0mPhjmaACIVeN+GP2D
iT3qbdb8F3JKe1WjMBTX6oX5vn7KBs23f8wbGw5+8dKe0XGZ7dspnyU1Gb6LMzSb
/Q4vupN0m/4hWhzNaXuPWzBLZzDVGko2DVZ9UHO+7f5gxB3K/0quvxHXduEhpq6g
d8Rs/mDYC97ZE4pr0Ll/b40tbzRv9V4hJ4xK5tpTOO9BOUnrtQDYxyU+0gWLf1ti
hoGcDzM+lCgKste+BxGINh5B0f8FrV6u5JcY/DYrsFejULC6nUtDPEVGExrsqW5n
7evmAeAbiZYRcyHBr1SHb+0Stvvs8nuiY+S+uQybBcxwDyu/seLIMRMJ6xGqhLI8
9jh3Gbxy+S12XDYAR8Jo2BunjtjOkXcT45LFfQgqGlO1OUqVx6IHMkeLr5yiH5ag
NO0x0yJdSzXLvCVB36v+jE0H+ltH0J7ZUlB+SlKw2dV+MIZyvWY7uvTH+HKKH8p0
F7FDiVz+yrzSVihslSUfLBpbZoIm7iwm1ICJQy9yVKUwiJsupfD7DqBYm6x3jblM
Ch9Gb+Jx3mv1ABBFVPdNQ4rw6FBJR3L6zf6ppjwBAbfDN8mS5aAFgwbFLcti2SoM
LudIA1srunYofjuaYyt366tG64zN9AUrI2YFRkdGDyjdHxp1n2mblUOeh0ZI/xqC
XuvkAKlpldgZAk28bp90iZnOskb50XM8dSDrAraPJKTiuJryDNhdihZX+gHAXIfX
dYcjAybfKPY1Wm6EBHfuGr7t+qxLn+bv0SwupEETwWmtGHzETVn50PylFIeRJ+XZ
t3OJoeD2oPHCWlUUjOQf5wgV04ImIygMbfro6J/ie57EZF7ex6k5hoA3Ja2HzRXY
l9SKZbY9panx0j0Q4YdJypVFUAu2LNBOkNEGJOWBh1JAxl4yY7oXBrspAX59sjb3
QGZIhOAV7HHqNYXc9yBfp8Elg/0PpbuW6FOG+mFWHnJgXgeD1vfpITSxdpDvJ3sl
W+3/YDO6Pj3sopGdvmjjGuhoDe9Bo1PJjmYfex1CdHC8jdyXc8i4M8EiMsexXfEn
412x2n9vTQQbNTDwG0KjxE6otM77SG/rTBnbcXNM/8T68RaPQtomkziHjmjAXxfO
TyiVh85BG4Jp1GzJBr9+3E1KlCSGHV9heKgkYbiFdrxYf+5hNcHKZgZ5tkdoyqR6
WAroGJrtnVgpn7s9oueqbnKiN9o/4O7oxmkFViJKFjwf3McQVNFAzA4NPJqvs0/7
SYklK8dpSZdigYLG+ReiB0zKeEMRQpbt7398dq8TOzyR8gZLS58k6k70wIiUzuh1
NTMVsk7prpZ/ZFZ3LFWLwEO8Zut+NITjqNrdI99bHGWB6Wk/Sxcy9C59XCpJXmnw
sUWvVW6wLBvEeJB7u0gESS27TnBj9rA6YyMzUb1E8GWhca0/OZZ0KxTyd2cVN4uw
mh0OSENsoNSuR1oLodLW68h2GAQZMg2hG7LZeaHdxDSdqz6cS9U40excpLn2REPL
JsjjWSiPKAbk8dMp8qZTaQuI2sfq/Jz/eMtJqwQY+P7fAUbPq6LCkeWntEPapT3M
wkIjBgRNxCBT2y/CYiOS1JhIWFnMcmhbVAjkl0jWdtUTaJqcI0GRQWPNbXA4Xk9l
xoWMSO338faFT+aBfxCFrsbebmFTcYlYwy/g8MVa4Aw8hSAFU8cWomkZqSuC74gV
dazS7E3/Ywtxqe4V82WTtX0HXSuXcICEJjlmQtwiNUktgETmQrGu/tuP8Q9kVDWI
NX06sKfc2nQvbgpp4smietkb0zwxWli8aNE/7w8RnsDrZdWS1KauWCUpKTJIojOA
fFfwFSn2RgSeQSVNeJ6qJBuMsBXm2YLXddT3FF3zllu41cH4WXX5tI1MIFCalyJX
kwrLCO5Y4soRy3efj3ZPx/CCJ7Vb8NP1fcBPUMkM3TrFo/BhD4SlA6yY3Tgf5GCZ
O11kcnECPa/U68IKWKrlPlR4j2iXx3igkI4hj+Z7TbuCm8sZkm3JdzaCuvUOf1RI
CaH7aCcZ2Go+qroXG4T6t0vQuYHtawM1RNK56KPtxw7DS4TtkXSb4V+YLsiArlFb
8YsCqzzx01/6domiPqB2VHFYWQz02GMxf5gLSX7+9Dqbyu1S0V/eU4klufuIQNI7
9XUomsmO/UjxDukun7wERWTQhEhlBjYBXx9OTvISgn8l/cwxw+uzzoqxv1/LZD4i
VyM3XSuQcXe0SQBqQxGvJymDWGninAxVzZaft4qVjl11EzY/te0DeF7VpvACksmW
grLlMa3P/kncFiu5L2jpjchtVhNWgYSIEExM+s67SpFFwWiRqDfudGA/xsT9+KaD
EiPRquG57V61RBKBXXowZ8MQPtBwdDhvIWxRrhZpg9CyRreMJlIMY48m0t+t9qxo
neU1Gx9XokpqjikMDs18TGdg6V0GErL4k1bpcXIEu25VE4fFm2xGi1xVSCSFFhTX
0ype8REBec68XfD8r/0oaKGXZ8B/cP+jzR3bXxxW1eqNnQfEOAkDoEJxx9FJIPyc
OoXTKjsHRTh/OXo+SCP5V3lIUsnFx44e9oy0KlSTMSLDSAQeJLc2AG0tIf7pVM64
IcXO336hIvhMkvMr49W9lroyNKPQCsf2eDubASHyjrVKxQLdBLrUrbCSvTup+NwA
LVdkxg+FWo7dDbHd9Lk+fwxL9YrOc+V/IwmowNU7uJbn1ZLBbj4a/vRmFaXuzLnV
HKFzYAELj0s/60WUa8CWL41kVtgvUaFLorJfNFzkMY/ofyq5yK3DxKtI6caUGKvB
9Pym3VR2EamU5tWgy8W2AVjNMSPCwY+xrve3IJFA9wEAikb0xh5cbmR+iR2eQ9qX
g6v8rH5HkcdSyOtMPIyzJn5NQw6GNSzjCfhqlozy6JZHB7eHq1Ug2A2rt3XyxQQV
4WnvbR+WE/AYaR49No0M3Czf4Sbe0sw08VCNChGH4U8NUERRR+02QtfK97/sSp00
X6EJQsQxR9KmIrtCWzx05zJHo4Pihvw0L9518RlGLbs3Bq7IO43PjuN6GKZbpnxv
+djLicP43tGdUkrfo10n3nCfzb3Ed09Q5+2t9sh18t+iLKsqJPMVc/pRSaRg9zL0
99A7fLga9w7L6CjYo35ZMQWa5xcle4mynYDLIcotQ6rww8Vfcr2EXaFg22DgFXOh
0z3hv+JQGBOSD3R8E333D8zj2pO9O9z1JIUUg4BCHYJlF9eRCUHNr/6lV7iIsw52
V9vVPgM1uxMA2CprSZsiC7b9lv3Szlup0cnpZY13J9qASHq7dWg/P+N2AVPzE1md
sT1F5tVlMAM+09vbQPcDSyq5/sNT2lbjSzz7MMAOvquTuMepTSHEuhW1Sf810ml1
AskNutp6hUMjuxpKq/1niNau+TRWNLvdQoiNjA4DQQYoT1nWsagIfLwQDUNJlaHL
gU6x+Ryw+XGv9atkij9Y2w4BPnBr+pNZdMnaj5BZcqtsCK5dI5ydmARxBPtfG1f5
E6eWcghhw5Co3U8zhDeUKC+IFZqbw0F0GK+yUQNbPGBtG74+KCLkPKPqHYplUr7v
ivdVLKA7lQu1yRJCorbFGzAimWUl6scSuDqBkgHZ3tw0QJgTO+dBpsA9fF/XI03+
6djeniTIYzTf2Z5+1Ncu0eL7sbxEGQtKhzR0x8Hp4U4Y/BAgNGyz8uDMHg8SZ9Se
ANHHYG/6txcLPTnpiui1BH/mww1W9qzhXf86kkt0QSoJ/M2As9/GMGRwc7by0H9o
kerku4JojqJvlBFkl2Djwxwki3ge1FKVX260+YaL1Rc50wOESkoyX8qxQMLq3N7X
hxh0J02pkI3FBa9LC5ztIe5rXssyHFyH4oOwlKqYSIqq2Tq1+Dr72hlVm+andqWk
YHy5DAFbq20WZ4HIhMXsqp3r6Dd6DQxB4/BgXo19lxZzzDAatHAI8VXdnSum+eK9
YMR3cfw/VFtzhYXyQkb7LnzcRjgqpODni5Zvmt2Ih8dsRe+dW6Q0R4u9om6oV3Rv
TBzZzI+oRvodhj5guiqpn+spVWb44gJp1IxfL3AvNpkfv2NsBmRu/fq+hbtMktox
og0Nho1NAD2WRN1v8yq3oPRYCLHsasQKuY6TqRCz/1y2g4ceIZC+s6+51oP4VODb
DcICkupRBWny0Ju7su1eozE4DMZY1V/SI83EbkaiLN5Ff5a+6qhd3VTPBwFj8uQJ
hCIrkWHYJfVasrTNhRq9nOj7OVzPfwRdB7grFX0vwjQkZGCOs5ALA4zz34w9Vnt+
3/BO47wekeMx7BCTdvV8cd10CT0G5ENe4v2evSofybUKADtPItnloBsMaJpivar2
nm6x9I5FNyJwd1unTO9oRtwrQqL9a3DVCd8WszPdxnpGp1nmZtpopWQefbv87rHW
52VTuD+IRql3DNaAd9hR82pDp+INqjrtfi19ySUq8K5lXTt9ZpJovQWY7h5En52y
J8qBYts7oHcrAod1TQAoFl8PBFDX2hSVOtS2REgcffl5uBqcO4ojAjY89Oqjgnvz
csXYE1JB78fLkUrxneEJino9x/j0lCuShZ4MzZHCs55iLdWIxDIaDwohU0DtAa7H
6uo1qckdrZiWugHAcpNmiF8Ddgl+v/Y35HV+A2kHNbS9M7vvyGe9tjC2lVfht27K
XpuceuN+tugQwnZeUJxud/BX/XaE7mz3yWR5nVsyjikjusH2FrnONtzq6lBSVOSk
4DqBYasDIQxpq/zDa7OCK7pTtrCupO7rwlwKQN8WU9G2/dncOs69xgnrPC7OPQbX
PpGhCRE/GWZIoG/Zz1tjZUizxE5hVoy+dmZOfLTRUdF0s9pg0qcIKTp548s6UaDL
M2GPHpACGFEvoC542Hs3Q/dBRKbcRsm4kgYI2R1Wjw+PT0+T9j7S/m3syYQ6yxiH
2Li9BV0Yjy90WOPHI1zWBH+HkQwTs6aEI0WIFg6/60eBNX/PUOE6F+czRb1bOZ08
jgHCi89WV7lF4swsY+788E5d8OpjUph2qdZcQvVZZw4cyQ5rayuAIeN8CFE+QcY1
WzfTwlH9W2nF0mv3EgNsdDhO8eQjlvkGkmDSi9grwdt7Mt6/IRmU4DE6zbvcrU2l
jv8wXEhRaZbCDoklUPFw1gi6EaD5QGXJMwdYPkq06tYPX4dnmCMlI1Rn/5L1ftyJ
ZtZzQytkmtOjolkuioV9N6HIT4LoPkciGraI+Xenx2tGvk0mHbdIL4qs5ahXXD2T
cpvvFTxmvKgNkZK5HuLdW5tb1IYOw0LO8SI88peS7uATafOAbrqZfIwMyGjFmkZ7
mCKVBaeXr/b3x2TmprXKeEoxnVfMzyHEXpMrxSt79aGc7zGeit7R2S0AE2FnZqgy
kr9RiuUQr9cvbQpsIdhfKzJv0h7qE3nuENJjroe537hSApfUkJi1SJq9vK7WiNvJ
WWET4++qhAJWVbMt9DBW9osvEO6E3DXKT+QS3r+SonwZMjEixQC/dC4/U/Cxe7Rc
bnXXMFZN7QrXoqC0JZPsOA3JMSx10A8jEJF4pq7lYWf973854W+kantf8WmUxaxf
6Wen2O7q6Wg118P2Fch1VQbNSosoUREl+CLJYzeuIXRoyGB6qcf7VEU2roxlCHZu
osdCTFfUgU1E1fce98kwhKn6af3gOJp+HG7OdbAhVk9x3gZ32e2uj/elHlDjoA5w
R3KlKJiwMML0Ni5MGc2UZkyxBIMugxOUW6/ec5b/1FneuQplXQzlTXBbWO6LzToO
cJYAp6UYx5pW4cPXpCptvn9rb82PIR4QcYbEk/rcmWxF1eBLgKr1WcwNrNihUR4b
ePaVyPVfxvAWJD/uQQZPW3Z2IqDc4CCvhragDAbtvVkFujX/S+168c14yKzg4rcF
bQpcBGVsxQEFdUARoV5JPnen9Bfn1bQDCoXMFNpX8R1fqJIhTsoA23GXG0Tn1wVR
dZ9dg64YUzlE6/MVRt8P/2Ge0g697Gp1eCk60m/SE233ptr8KMnqToK4MMpA8AZV
OthTcizDtTYH2KkMEhhSA23ItN7Fm2Tag+m+BvPDIMyl8IJypACvjoYHdc5neJFv
2LTiooLChY35faKXbV6qk5xBOEue6WhXsV4RB/+8onvy8Pl384sdG0g2G4ROOfCs
pDxYBgKFaJF19sAbHbNu7vxuAYfhfc8qknuHCBAwhL96sS7epFCSAnZm1DM6Uhya
2CtdpbEfc/9t8dtzSuca4diUxza/FWRIeUTJuoBjXcDIkrp0korOdg2qcFy2RoJM
GCkBHN5zaOOK647QL+olJK0MCFriOUMJ5SOdzqTihaZjtLO3XJqbgYE02jK5y9Dq
1j9xN2buVA6kTS+DzrGpACDPVN8fkLBNBSZoa6XJm0eTZUMxeWf0MBIqO6x45muc
sbXqZtZgCJ4m7tJdHTCEvWMQEbS5Ktvp+Hzo2MdKyPRz60SUVL5E2NFiLM2Mh3UH
JjL7apf4qI6F7r1sZdgxQIhLrHsS+3X386bjZP8xaFZ8PkAOFVIOv54hhrsjz5A6
6PyJoT4oX7dz5j22nrgBHpKqZAFoZ0LLq/3EWL6+SD0GQuZVAVtUP8wBs+0Bdnga
UmR/YhQ71qDJyHLq3H2RLcUpPrjYj0ilR/6uFDqDLtXs9j7xvdBHl27ExFBTwLdk
9c9ZPy/PJNb/J6qlUBj8SZFPv2/VIAB44l2U61Q0M8rQOp2Su41qjx4S8TzWVEru
F9itywtGjKIt8PtJ9m1dqvgrNrkoWCj4do+0JYsRwJQXEV8nrBcXFzPDNRI/4o2u
cuCVFc1Y/B59NKBFjaYwLIE4TBEJltG4G3FlwGUBm9x1zoGeJEdpCv2ngePp0fWX
yd7TJ8o7gDIGmd4scOk2PUIo1yXarKqGLIxjOkreB98d6SAsghWYN/+hPZshPdPW
LEiNH4nlYTSRz9XTco8cSIzbgiEmQtajXlf1xjrs3Q9uu3/q0XeyfBqpCLchDBDF
6vCLUbKrRCAKnPlrs06/m3OIFxNTM5okDbCAmWA5iZDI0yKDFd9WgX7OGPotbN0c
QztM2lALjLHHUAlqCU0GkZiVXM3f9BoUT+rTKEht28z+G8RCZZW+tfZQqIm5Pd0o
OWKdkBrCfgvEfb3ey6h0We78UExyY62/lH3INhkXlgeK+szYjciPCIPV3r00CtJ9
ass4pWYhF23VjeqAngxXxQbry9vxPIubD71ZXFVdcB+VGrG97XGArYQeTH1K6QQ6
JggdKIATOB0rUlruH2kPMASxgB7wqAixPUOk/kyq1frE1g5J9Du9hB3pVFxxujMg
nnmQrQhUCmseXGirju1m+3BzJC7a7eGh6cGBwnYF/FTZrSsL005W+2pMhp+u1aTt
JhkjRbV+iGLYMgGOo5ScRv6dMNG7M3dWSG1/h6YrN2idBN3bPBYiHaJ8EYdeNS67
TZp4C9a+sXtv44iK2F+5AKjzl0HXlrwBfbFWN7vA+XCPPkIeAkye5FnoRsVCHpYA
tbK6dMxi7XBi0ykdXNPPABMPXvD53y1ZhzFGl3AEyFGd6ApvxJcT8ikYEMq2jjxT
Ynef2pVT1UyvmKgV8JOzFZvOwUKkNxei/Xr2SERnY9wJ4nj5kzwSlQlKNOW/p0Uz
oW8MZqHV9rkFzLdPinnI23VXDxMGf6RMWhSS+IYiWumlFcIE7+giWiJO9i1gsO5z
sg3bU40dJXhlaYsKS+fn5Y1DQAoPTZVbtoto0GmKPoZEM7EH9ZsObzl/mbaQtmkc
2zLdt2MgFWeM2wRLeFG0x6aW9hjv59upj3wABVTeY/IuzUD8O/YljiNpZanTPJmB
kLdIb60JshsqEZOQLGAIGSy0yxpBu0q4gp2ZcNw1AjFB6pkSK5jWKcaiBUzVglAq
RwsQfITP6sxS1P2yIt4j98+bytN4MuftfA98vVFr3SJGVMFug6r+RAEFD7X/umoY
EUXc66YxXqK9+JxVn9VXVPRmnQt0tiqNxjv2v3NyegTVuRAgfqfsF2NrNwI0mYOv
iwd+aCYNuDHrRGQ9jd+Sff3wj1vX4X6M0I8O8I1xyG01ewJuV3Q0Go3n5t/MwLcs
+u4cHPi5DgCQbYxDgiZLboGDh8TvGMeGnB7oGRoU7SbL77DPZQRNIfAU4Qz/UxPi
1LlduHScAEiNDB5tXk6K8AR4i3jeHJfEbqjg0Yje3VykHz/ktkuawCOfNbyJQmgO
Q8vvLAWbdFMyn+ksU+SyBP0poR5hJb/QRiCc5EbFeCHo4Y9RWpnZGBbRkKGny/4U
618rcQ9cb2a1jo6c5belgIPFkTHzJDG41HVInR2TzxlGkaeSvLMZBA2qIL//L+XM
5mzA46tdO3sBMnv0vJrCbaWqaW5qb292wrzzr52zvSO0Bw7dniMsvH6rXvwhQHHu
IUdrdW+TBpj4gjYnODU6wHKM9OlF/IwAIgVGuokYm9Xv+eslt/L7CQ2ld6pcpRLg
i1gPdMbinWLq8m1SnsJhzzEDftzND/pCdf8Kkqa54J5KpQSsHDLTvAGzngIHBdZE
nLdWa/S8w23nELutLS0exCRGIEsU2SYdASWF6Q/e+tgc4a7w9F/DqZ1MBaapodlN
T8HydnVdKD1zRX3QDxhKIZTkT5iLlMts0MXKDPaKQHL/0GI8P4c2ujusMtdBSFlv
Sea+mrkXl4FhJ9Xoa87T2R2LJbP0spXVUXUn2b1yIyB0BZNun7k7DPBhP9RLa+yy
mg9cviwoBQIjjLvzfWOoqNYuWfAOJanMsY8kZ0lvh+7+awVux3lx7a0D8EZOfb4p
K7f+zGj4BsCcGjmJlylz5xkomIplOACEU5c8Z0xCKNNaOJse0BKAvnpZ/6WgiZ6S
mV/SAXA7uUsb8EQPkFS4cdVrZa079i96QMsYb8fbxJk48/kiIUdQE9bldvQxaUrm
hK37WlffBb9YDc62/ushtnZMFmHzGUM9cbwLO6cbgHjPxJ+DoDyRIdtuX8nFk3bD
5NX7jDOxfi5yTEuKy7E3e98Sc14zn0U4zJ6Drx/rl8UTR8wrZEK+LHV/I+LvSDZV
Z39T4N8nRILY9R3GpK+x98qOeurxHw8n2O72sLwzLrJRarL5Avg1mKKQjTaS9mok
Kv0Je5yFVwIl8ldgb7kqJ/09ySLCIVeSzAnj+KnNuPSzJcn6Da2HNRzlqxrM8Ex5
WpaLDx8wR2NSb+n9stFdNVoSlRWkmG69BSF+jw2pXwzbrTBYPIPWgvJ2RhViHfZH
Ym9mGiTIXdQeGMOf7au+JGmJVfvN8yQbEzQ+1kdQudJdZMp8f6efhv+d6/THGe5V
RPNovmg40BepoY6A1F73ymd8YOB3sRVhzqAC64RhrmEYlnqsdk1wxTtao/p6wUND
/fHrzqf7xOiqFcKqOD6eu8hQXiA8h9C7Clwbczvy8+oBJLqm8nrNsgH8xKSxYsKL
24Nu3NQsATFaQwFvqz8GA9lrAKB0uyv+R1ncLOSbfX3vGGjzRNYk3+1xVT2brRqY
P6QNRe26x/3BwrxCmFoEuXwsF5vMgKggzCjstIDcEJ/gvQX+ShUbxhQzEnLq7QcM
hc0UQnpL9fWGhuOoI6KnZllk4ysy/k7eYbRXokPoBeIqlC7nKSdt06Fs3YN77xSD
WknYAZQKxTFzpk61cv2OasO4tBtRZpMRkOLoPSYglqgreB8OVowIMAsLMfiYJ/5/
rMAfUXftTTanB5y5ud2qMq3VXSofGuiZm8uqaXkYr45ch5Oy3G+/BC986M2huhHI
aUey1GdgIjt3LlL0FUxuQfy0gjLeWZ5gSfHCB2XNZHw9cS20zPj5i7Il1x5uSNZd
A6AQYlf9TBvUFdhTf9j78S/29ocikxoCE/4uWIHOCA3duqGKKOSh6LiOBNu8xcBg
41gZyPprhPplUNSa/8lHTuqG15Y+LjYg8Z/7/Zkum1s8LGuOIzybe+zS9ycK7HC8
UWMC38QoUa2lfcjkWECvCgxbfvgfPYTdn6HFDS8Si1sqZWKd3K2QagOh3dVytNmm
L5ED5f3HQdCDtwgLIRBmojM0O4DyCK2qC21b0auwNn9RCTQeXCae2XHSaKWxsXao
1GVJ88ul5P3flTAzS3qYEicTwsrdlHHpmDsJHyDDM43Hqy+p8dIkfbgDf2pWCyCo
4ZAICSbsDSAsEawA1vVnLNJemsuKfYekiaGuxaLwppojoVH1OfkW5rMj7BnhgduA
Qb+Marde6riuawdAGbVH9zq0KiHuQPoB2RjB/23sSWugblK9R8K7xR3+lZNnFDjf
OxB9MZt/EBGO3NtnOs+WOfqo7K350BdUf299v5aicoFWRStmqdVZ4TPo7gp2m1SU
1cFA+WPEGt7q62cIwPvFiqb2kwIDSSbKZYc/+9kCwxSsdHUNVVM6zKurEV1IwQQG
zhTTAewb3s5OCP8epliFILFvkTK1UcWDsBJwh32HGcr1uEU8cXJTKTbCSVbYJ2c3
EV2L3PYe0EwiSnZF9F8OKaWNIWcgkey1vxeS8nkxkO6bQjdqBLMY8FZz3yNWgteV
KJm7du0yxma9S8xepeMudS9dFgUHQO70aHkMh4VbyDnuOVQLhl26OwHWqnmWF0On
oSTu9WjQC4YQWM6YkZxphUjJaYiE/0t1fQPMJ1j3BeKgpORHhOo+Cxt5ngAKUNMA
XqxgkDRL54+xcdNvsVgs2q6dKgLSk26qrtNM6Xs5JtVT5X1uUSxqmmS/EQe0EF3+
fREbry5/LhW6HSPm34b1WwPq7+v0Sh7mZc1tm79OytG6fHhoe1KlDSJXN+FuCAaE
pL2SpMqEiFmgUd/S2+A6aB6JzBUS8NI05HRrO8xyMuLbpKBBw+MY4m9WhPgHRNm2
ZxNNwyt8p6bMYpFAYjrKPpxrQhTS/ImG0sSDqPCTkTtd2QV3fF/49mzNMlY7ML5H
CfLaQIAExA7nH7hBJoQ8ODfVQgBiucJ7nlc+QglEWhPuCCBaZ8r3mm7yTQ0+uqEF
rbJcXhH3wl8ND4h68vnZXLhmR1KAAJE4jK/ZOlzQ4ErruKRy4iOKIAKZUyNwSFbt
NRAdr3zvR/yXPB30JI20w+IX4cR5GTgKtKZ/Vo20onc93IKVARB6nYBpX+HnXik2
By9vnj+jN9hUG+H+kyIwCksKiqvgu9wDRh62FmcNSMASiZNsUjt3fYXaVMqvXTGA
ckihcrsjLK4+w01PwS0v/B6tDrTnPQzRn5ctfO4pNHMuKm8y3AxECgjmDFniAz2O
QQTU5N4rDT5YLVW5/DI8w7CZYJNDLoNDnLt97Q4TysCiRg0bqlEcBkQCkomkdcQ5
4jDo/pDsIGS2mfU6GMn0pZ48/gRv7ZKq7km78uS0nQmg0qx2bD+27Bn4ZiIpfNLW
v4ImOBR2Ur2wTdg7rVTsloILIqen5BWJrrPqZMvmUY1xgTkEAOOctvCZ5FW81R1z
Ow72wZzQ8DqVb16x60I9HDTIgqwnaHeU4rFxJFIxv2+oN4NMTEcFd5TwFbbi7U9z
zTEANUcmDvNvkfuYCzAVR8/KHPtX/8pYZv9M1T1EmECtqvA8AVSkMhC355VF1tw/
0kVC6+sJHMNJ7DMkoOaf9D+/OdxJI739MaWhcH8UhEuzPl4lLXTIc+aFwfbVLked
3+5XV4kXPx7j2aLj23cilVaWVjar2W6N+6Z6fzAqhJYyqF0QDdAP1vnpK6Pr/fWv
L01ws1zTALxpAKO1GBM6RLVd5J/wsZOrWJ3Q+vc86HUfmmiDJGIxRq35DVf28ZqH
zAmc1kC4Pdc71DjiMTACSWi5dr71BrFdcZrZ6psSzDzWK5DhqLpPrsY/sLwOkYXG
cLIbI5iEHl8m6TAdn+HliWgqMTk5h1sDOlR3KmyeBzB3amtmp/z8mm22pfwVBIOY
SBO4CGSp2kKIKw06yT8ojS9aVcsfVnwKixNTZwbFtpRmez307NJb0MjPhrQUSTBU
xx5dkssKEVVgETWAzcopuJGlWq7Vl2unf/XvmvEw/ZNGjn6Hk61p3qsjbtSdyeZp
TI1z8/E+1BKizuzsCyieVI1/aoX0fxA0LdzSkdE6HuktHCO57T5y+qWJG2g6w1FT
qEePvtUopFWZ88eclYVwUGaSwpUm2abaMTzFoGcJXwUjKL2SI3dBV4e2IGFe2NuP
ZOWX0DiK4GiMDIn9shW4nnT46acJAcW5cQ6ix3+iGYCGteszkyC8JjeeNIziP7lX
8/2eRcwFz+wUmcg440br2z+gtGM/Hw2HemgfXGe4Q+PnaINNyRAt1Gm6nFjvyMNw
zkMZhGE3E3+MLMOxou0K0VKYuFjg8ScA8CRd8rYgFE2U9GFhPfaYjxbkSsr6Ut85
dcQzqIQm1SNXHA2DwPzXW+G8Caj3I9Hif1Enp2E2cXJvFJTq43WA62UTdNCY1Vpo
ZI7dINLr5QFGQ39m+pHamrJAA/I7OXkfmlB1VQEaxWViOJqGc8CyziCe/odaeI0Y
WH9jzaovAsgNDPoBNslUs+Dbj4f45O2qB8d8pisNxDLvf2L5Qc9Q9MvXV3+/pGJD
FC7mEq4yjebG/mG5y7NLjWpnKGUKdbIO+XzJxIl2vjww63MeMXKeKmHyF32wrDTa
mEZ03bt4Vk12r30MWlMvevM0U3DaI4xmfF/tfS081oOixX4nVGHsx/WmiLrH+5LH
jlI8EwhtorzR6i6kQwRV9xxmV9zuliv1C5cbCQ2Jv7x9ILVli1lSsTjrLPWgY3/I
oxFNRXeibeNuIQnRAeIqu6MY6yrNjDe5NUFEpmz0SotvHqSaa5OwAOqp9MrUBkRI
iwwuF3yUht1709e0QRIcpu1erh+6gbzigT5KsoWkFYdl3z4VjJo8B/8wKzuHJy7F
/4+80YWg4Qdghpt8wGJDnXAov5hajpInJ3G1wi4V3fIGN6IT+5XHAlIqfMMVmEqb
0i1qMrcYI6TfOrBWMDdxwH046ChXfmMf8h8H9vW9pVQ1LcaiVIXJu/quqgtUxosb
njg/mBXaHbA4SEZLDQpYNDm0ckPhe8DU2XA3q9suS2OGtAPN4FAIP8cg2dMdQyzH
5JiiT5tWn+zs0bA8RBUDsPP6wkl9PoS/e8Ucn6/amiqhsf68z5poy0mVEPqEnsb3
+3go6BP8oSwq8pJlPVj0QyCyb1IWstK/+pu1GIkR0cZB7BufvU6+yHic5EZ8M7iN
kfkx6vo3Pgfz0gk1+uEbUjewQPUb3HATVXi68SlsxLm88ffZXt9M8BfiTsbDX9w6
NB70YWrSDTLx9GKanhqWZpJdycNFbQ6SV96EMRvkm1gUSbfHtB9N3gXawC/Ywz9i
HJY8CLfsudSoFJvMkKk0losr+MAyZVs7q9Pwmbhnf6OkCGJsXeLGdxJIpZSAtbIE
qra2+3apkVcDuzGdd3o8Azv861iv1KbjWUACx03lAsPeWBDsybzgFxc7GU7P6sv3
XZYb9dYbtvtxDQxs1F+0xRY8bbybyBpk2lI9Ye4OlT5VHxjD4TaPwbj15kFmbKA4
TF5kFHh/HVPAIqQKiUImYsvKE+SNyxfoW1ruVSNDcUTI10yY4EaCtmejHZWc36lR
ZzsRSI8QbD+MLfnwvutDba51w05iEGjwWq9p7M7NgobTEWUl3PMuQOgrHmt2YOTz
M99RU+rdIUCYF9S7ee3K4WrFMweWFpx5hvFWmgz+s8Gk8P+449MKZC4DXB30krER
oK9/MwVBye2e27gNkkZUh+pPimTC6wYdwWdmJbQK87WHJg6uJCeLEsNvvy6GWAN3
Kr1/4qGeSd2J4r8IVUCAgabkaOzW02RymM/igfoS8QN/ryOc6HiIi/6vGmfSb12v
sbC13Ue0/Qt4WEmg5aO6ajwZuoMpVByl3rQfGxw3x/aj8Kw5JCDv17LzU4xnMXy2
k9nasLIE3butD9HWW9HPyfIa5N8DqshVSbGiym9yVffbsXXtsZlonfUnmoQ8cl98
L0dwBX40Ygcq6vWRSlJnGU5x+fzJgDLdvRC5hkt3691G4BidbDaEI+LEBORkAfFS
DE3lvSRe3TK5J4SpFZHbk8MOLiWj5Tc/bcZDyvxfIR6JD4vapstfkbbOHlEggiCB
IxH5uuy8TcPqhqjuwWLBWRtDnFs3YJSgcdI9VXvN2gs+dp/Yu9z7sscVa/IrjrTI
+Hesao4gRHJlPVrw+qZaZROIIwTPsPTr6cPRnUHhTb0J2eh/Z5OZVlerX1Goa0AA
VTbb3lIoE/gFr1wRVE/IlNcQHeBg2mZyfpMbkGSeMUbqDx9gnexXU/cwWBRsd7B8
RCF7znGJAWvEtL0lC0uEUxT+lqwmwJXL1ImHJWLN+Ssuw/Nlb+XVoJcZ73HVTYG7
ONVQwVYs/1mTbY1sMBXMZ9v/Aq3toxkjRdgDvA1o3p4KXKhjcYCFm87/IIcWkwu/
W/yOPea75pEqKkSCv7emDO65KDoleSNtcyC1bdIrv2Xl1P3hpzC9ifmON8n+T2/z
5GadTDAlpbLX89OnEPg6k37XVgsDjp5z802TfLi8GapMVs4O/xSDbV1I8kcT7kFv
FpCHchFv6X9I8K0xb3vJdtBnSpNIcyqDTYwsNAhbYj3ieQE2zm9ajmfX4Ms0t9lq
JnT2fC18FT4DxxT+jE6Zed7vBZWFZHtvNAtE9Z7ZLa7fwJB1Q8YcNyVfoyj1bWE7
sb6GPMGRcytPoVFiG+rfMKz5lKbc32d6xc3PbB4uAu6Hk5cxmiX5qwKvZBLf3M6J
xex7HcQH10tpxu8DzJhoF/kvv4t2bj+qk+wONs9u5aU6g7KRdJHsy0NGHmn2D0uk
hCgd5kNb4S62wRK/xB0E3Bvti7G0nlJHRZXmxOYzVfa1C/QF7/CZNUGidGvpLy6Q
KjKRJKz345zyIzAAArje6ZRsU3fePCoXviKdaR9L8nV8YEbCTtERiwoGURseyx9a
qrpobO3IWGxxXE4We4L9McQHVGSMzDMtssW178HRbAjZgVFI1yeIx2PhnJJX3bLV
fRl1GNrx3NRfjOJPkmKb+rECDjppzx+/CAFtQ58DLixfZziVyJOBoO3NOlB0twL2
pkR1XPgKDyIiP57RLGzhejQXq1lVzE9WsVi57U93Tl5ebQJ0iGsc3fport8rPS0/
KvUfKaIiwQYE/UceZvKidVKiAlM+Is0AwzIQ8d+qRJi0Ct5sYYl8wbQjC/tmXwMj
WUrs12ai0/YGJ3rrR8T4qQL0eCy+8PJ2fn0mL3xOCFOFJKBW8UJyoKGubmRYqJ+H
4VOosjJYZMjC4jOKkPL4U+8m/ukwxBI0m5XQFLd94vseoDDZmbiD/xWqBkDhVTCW
kynDrgVTI+cyl+7aiBOzqT4WLUbpmqvtCKzTUrbZh4/I972T0ItsLSbELnK2dKAe
jU0y8WdaAcq4mOXl4iad5mSq8NnJdGq7LQYjHzJDRIU+NscUGafge1vJqkYrYijv
Eo31K0HpUJcH2L7hiywJ3OPv1Vwr7oYNx0zT89P6um4++u3aMA9bXabWtArajc8Q
2QXW9OXucApe5X2vd7zmAO7vc4VblBlqxixeGs+cOsT0zWi1V32VtKoOv4E9UORp
13jlguTJkUh2WJTG2lUcRhyaoHzQTAFaXr3eAYUZLYoPDvB7+Pao2SnYGf2o9QzT
pHL/q3GjExBRhAvkz/WAHlOsYSMpyWCJW0oSkOfyo2OqH/GtvBt+OtWnVgkBoIhz
CT8mBiATYQoL2+uhx6HK/OmOMBbDgYfTixaS89FCnpK8DteJ61H3cqW1MXkSv2sN
q1rw79BwpThJwG/HxoQpIJNDYewmdjvIJ+3cLWE1H/hggJPyCsDNVxB4oqxMMTrg
IaVXPOoZ598w4QSW8rMiSt1om2DT18hgtCXwGq55y4vTGDsD5Avv6W3KlJfxhEzc
3K6ss3+lsgPLz8Qhmc3Imi8CCkoFCIQbf53EusHsz8WzGq4jQ3E7HYJipGbKgXuE
4hxlXvJTTgMb6u2+0N4rhz0Uw6w9CHdXLBiffcLJF9xDd3UhmdCQjYOqRP0kc7st
wK6kUJyq2ODIT6s7mQVMxQBfjUsVc3gVylMjfAWvSa0/toxJZJ4mnAvJLYU0y+Ar
aXtRiWcgU8xESufqZELEJsvf3YEaFe024cvAYdtqAuiBlmkvoBsGZwyH2x/DLd8+
MG5V2T6Ox4pA2iNgVA9hWcN+ultnGHXKlQV1ypm080BqzS9R2gdm2UbA7KUtMAL7
Dt41zqC/YdM/onQF2rYR0QsunM7o1NI/uvRqdFkbWN5sL6xj3dnZ+xDKfKvoqTyr
5K0eDpr6GT9Tipkgihn7W7J+2x3BNw1klCXUFGin2g/hOA3xh0gt2cU94gb+I3Ln
OrndlXLfDJNLUMmYCDNIHDobQuQ5BS9FpCfVlhaQeii+v3Ui4dVqndXvPw8Luvvh
0m4Tg/iztqfxut9C/0mGfMmjdbJKlgu4JNTl+OP0Ld1VuVjHSia9aaJZ3yM4HY+2
b0N79kR88mZH1zEx5f2GBElzxHqcHZIbueuEUDLsOplmwOY3/amU5FR1p7dksicO
8HUTg9/oJd9WMEidFhQdTBKpRPTI9Uin1EHgD6hN5+LafxalaMFyOVjQaGu3errZ
uy6YUffng4mMWs7gzTQ32I4KOL7scYE9NqH8h8qRs9UiKaPz82DcXd95tk0v7TKF
G+jD0RVAIYD/jCMBXM0trHVMu6Bbmnn1GTx1D5P93V/x5JVYa5iTAMxEyxObCZf9
W5G5507AiVD4YZ5nrfn5Q1/qO4kr9YkZJlGcGbwhAlMp0hcjTT4hDnljZDm5bo3w
0zY4Wdv+bAHagVP0WrNdH4cLdQ6JsljPHhNtz4C3GtOP18GM0fcTpUPdscJGLD91
80hCmrCJfFWh2qt1qFu6D5vZnOdtCd1QZQBymp2xtOxdDC/we0pYaVt6U0sjmJ2V
u0KzBQKgsYYtbNgILlJh4kQDWTA50DF5pT29NwXWKELAi3wCojKgtfkBljLXTpMg
lwAn3LaywoZz7haj8ZqScvKaco3kD28Foq/QcE20gnZBagyMM6P0J2uaTe1uYNp+
ecY4QZE7qJOrCjtwVUwQz5F/GtagJkbiON1VREzKNZl7ytIZnxEHd7VCNHpEhfqo
5vSGVCfzj53Bom2sP3t0MgF8uVkgKtbSfH0lTDAcabA+nf3SAF4JA0u6D5z021eA
52ZRtmmTkPAaMX3QUwLUxNaZ7tx6WEKVOpfr5h68Tgy/8uaVMTSsdZF5F64xm/Zd
QJQVbVszK8tFmzg4i81OgLj0cFh5S+cNCmHa5SH+az7N4tixFlM+anVxEnOmFJ1p
IxgWS0cxAGie3aNEi8EnzMD/ghQJmixmCiIxvTJRaZp6hs3tdqIxREm/p8vv5RiN
4gWUp2c76VqoCWWOLqNtqvPz6dpsuVXhJTLYZVgnV7F9wY3+ejzxrMr3Ohe0ERW3
VqOr1/lb72gODcs3JU7bEcf8wGwE+y27d+aoBg0PZRokb0br13C8gcX6vCwsCiw+
ciDkbleEFMioXezTF+4tL67+IXzBlKlhR+M6ehCPtGdWtUTPcRzC5vowIBiekP4N
jqEfky5r41uMhMowPIy0PcvYMRiLUQr0MqOtuIZN0S/dmT+5gPpI4BKjOAQu5Qe7
0pzngoke3CgMjbRoWZoA+fcUe109eI8ksqUlhdE9pK7epeieoQOqwJ3QxRdJd+uJ
nwQnaQIB3ym38rRARCggYq271cbVkF597YSHuyTcdYsdDvfndSotwKmO3ZX38toj
vfRgZU5v31nnocX/OMSh1DxhmLVEzSBzGDwS1mefxeT4r4wqZPkTq9hRE82S2mfJ
E7q4gblOVrU+TdftiSD/ZXeEh4biWhtyUdzY9GzyHQgZnI5h1fk260Y5jcZ+vQwS
VPLIB9xWqobT9VCRCxst3TONHxpqaSePxMhgxf7vFuP3rpvLjn9qC45nnNPeV6Am
1Sy91o8MXrjpEkGDIj9Khmw9gWYBlpBqy0sFm28EaqK5K4aKcXKjuKKcfWO+KUmi
xOQrHn/i3gNAAzYg8QGEc0eJkZcr2fpaP2PpRXdkymyy591+Voum+25mSe5+hBYo
/in/x7WdPWJ7jiZioGG1BYX6bsMI7CnbBkFYxdTvm7k8cFIDkE2efzBMOn3w3JfU
1pFJ29jlvhRWO/5AHV3SlFVNWwYLOXxE9v9HUjbgIZ76MxjJY5xyMvLuzc3a3sDf
7Y6bD/axdPoiSTPI6IWnwNV5l7lwgRFEP0o+hMuDRIVH7l24Bs+7niUfj+CUCWuF
iD1+9zlt2W7wZh4X3EPzyOaBKT/jdGqrc/jYpdTcrblB18u1xT0Bu4adHQcYXF/j
uPanrRsArt/YdkJlquk0kxTw7H6gaeWxMqbgMWP7UyQhwOoOQSImf6LmevgYfY17
lEX4QL7rMyVyczgWSDRyOfEIRCwRVnUUISWSsHO14Pmgbrz0YYbhuzTuJtxZNlnY
vbjFTdCTFhiH4GSRXnnD/6pm/rvStNJlgJSAUiMoNQt2EK1U5QJjLPBOuF0wmYem
8vDnjcVlRYMOD8Ei8Uc3iQxJllEWc6dZeqvgpItBJ+/iU2B+dHCtEoLnT+XtW1dl
eX071JrxqOELRWcpedYcqBh6dpFoPVKWqs/wgJqMI77XsdLs8wKeB9aD5Cq6OJt6
PWAzNEB5X5j1376i9u5vr6XO3FuUN3vP0jSB7QLh/PC4qDMsWMGr7hb+FsX7qvzK
yOnTyKqYBFqrcYrK2e+pO+RNcTomvoX7FY1o9XDHQEKPNpo1M4QYDgOT2+IHASb2
MbwXZb+26foBkylHDggR0/CQPW7be3u2KEw8uDncmwKLQUO83Nt8itqvYSp1n9AG
8DlIDGQAXWRYECHJyWqPsWrHXDIGpuQeh6Pyy1i53gmwpaju+KNavSeuUXgj8OBS
3kztmtOM0W42ebPQQSsQS1tO7b+CuHV5sf17yBbsOEt4A+ua+Ks1pcWAG0qKGAnp
CHabrDMHzbHSoifgBkt98H/FchFrSW8pP7lOEurdghF8S+WM/0b0cqj6DXfLfIlm
M4cmD9ghYOJwwuIg+potQXUO7CBUpo9iWygOVuOQliNwMaCYba+67TSU1BQyzyHJ
e0/nKxv9I/uBmIWMoTNUT9QTiwvGqolyKlmaPdfcRBSbcVQ3mfruEXZg3llnWFd7
WOkuL7vzX9PjeqoHX86wlgT1SRet2fPRok8PPDZAX7/Yi2Wv8avEEFGJI4TjwKX/
Yna0YXtnhEKNPfilXBC3ZmGgmpYvyo1LrRNgEfWFsJUpWQg2Ry7gVYRhj/OqQTfY
NFvZoDb70GhjMMMOLKsklKaNwvW7k7wUPWgrcBnShsAneDIPCjBr8ibPbiaMybvb
pVDHXsMWqlpGAs5vIwWpCLiQWDbIwYLOalemsi1qQPRyjDkkN5fQoR0RQYXvXtr8
T90JsVXVrqR5PGNu048PdgtisQJlSF3RkaoEkGO40EDzZY5ApN069pXdyVoTwUeb
36Hg5QtlozQg09ne4CuEIJ8x9lU0ltlQ++qryC4H1Z+EjqJIEtUKzyZaWTf9sRff
F95nc+TEvcF4NpDv56X8pxjooKJehVXvkSbAnMcoGROPVr+gFIoguZ08Ll675qjn
zyoVwmqAxINB56eJ2KQT6cphOqG1V/wK7K0mYIuaxLiULGuI617SqL81JI800RNZ
5yE162vSe6BHi4pDEl8E1fT9DvVXnNfCoK/bh39qtdksB1QDwKT6MTryjh4KP3XJ
g5qZeqdPlt2teaguB92j0ICeYNnedfK5r4PywX6Abo0+tYCGHYeqpvQeSTaKca76
TtBWzgx6pf6V2zCMzWToUTH1c7d9hLGFDJuejeuD6E43fHfB2eyhfKhdFekX94k1
s0ZPXDXU/uw/7+jDPEMRizXK1ZccAj/zT0vV+dk7FvMDXMLU98zVQedL91hmtbn4
SaGrv9LJAjRgGxWdPa8Kxx/exQksagn5UxVZyNXbS3r3RwFZyVHFlGyW1/sMMXeN
WvKSD8+AHgzXp2/5Ow7YRVH6vX1Ddsc9PhVKp2iCThWVoSf6rlQgrPH0bLnZpg8t
FhXIH5oLJZmp7NxWvNWossQYLn9rDPX9424Se4gbmuyKlk4D77BwkN8vJkUraUi3
L2h5apt+OS0W7QUhFy5ruuKCppqs8CIZnwxPA6DQuqVqXOXn8YWQ1ZIH/U1x0xya
Y/7xhTCupgxHOrXghSobaete5uG7Hy6dxLgGvyCwnUI0IaFCdTQJxCHI85YdKgHq
FKAHbGsYv1rqvpeddQ52gWT9rbBAXC8HH4BCCs6QZdg0u8jbwU5S8DIBpS+/4OgX
QgjP9v6SwGxHg3MNk4Ip/XVHMq3IOJvCL3VXPEXVC6dUuFsnO1E/yiM6tigykELl
fVqyKuZwgobHXIGJKEAaeOPIuYsoHRFZYtweoQ/LwR2FLGWLCNBfbJsIF9TED+kU
vdGvp6U88dZ+RdMGKTl2Ui83G62naPRYZwX3EFOzabviTBfyZ53bzFIt/2eNAw3q
pFYvEcJhGKWPEJwhELDw/y59k2h5lCl30BBVo2X94Lhc/JXVk7mpwX0JSVou1qwu
pHMwxWeOHwMYIKP+VXU1WG+ahVik5JO6h1CHFiwLxrPr8M5BT4jYJjBPr9tq7RVC
Kt5JI7nNmdb20obNxwDjwS0k63SIgsVUlshGQNRAerH72HMNZ/LfXzs4walTIcgd
uqDABu0+1CoF+Il/xCt/fOfqkMjQK3ZyeZvgXIL8SypTSAjfHHI2nQxXSmiMI9cu
cHv28FpdUvnsrU9PFAaeB7HzsU0neYbtpb5pobtyzNOXAo6ESdnr2NNgC/duqRyT
EzzWtK2I7bfOOHqBcLUBccZJZEi0nzuSa4qXub0YQIA6kTqKywi6nEeO3jlvy7BQ
vdHLCJkaIgshT2Ff6pGUfFrWyuveIc3m0bZzPpoR+f0dCGaNQyoHUoBVBGAUzioa
nQYIEJCPEgdwIaujgZjCaGFNb7btuqgAMqsgsR9oWRKbvkwNElruR0sizrFd6e8K
48EnAmNA7irf2WS4nhlsqQ767rVJvAxPq1wUItxfajrMcRDEomYMjtmiavdV23Ji
okK3kdCGpmx5ICS9JXLWDbuafvrZ8/81YPB6W0N83CjPOyKCErOCRPRlvTs0zorn
4MbTw0VhnkB1jOyW1UEOcjqxQaOEmUz9ErTZhM0aja7EMZ49yqw7btP3QzwqQwL2
2U+WLAPfvHtnJK5lISZZlDuMs6vKbKGAIbBUK1wH1Cd7yoKO0OYGiTSkXj8kwMrt
6mB7hG+KS3d7d5Aq3bx9iPhHll9VjXbVR+/vbqyKSHX5OgKaeSciWQOp9LloFIcZ
A9nbh8L6TRltNQZTsdYFK+r/EqmoJ1S/m05hzO+o1g9nMiFMq9+/a2e4BCE1Hsl5
sRU/qHa3A9gYAW8X82tObk/tmFByMLqaSWfCDRPivBoZLyU5sybTnKIt2bhR4d5p
1349pdamV6n41NhkVOkJBRVTse2O/opUM/suzWsER1ELQQBtx40ozdHMf6OGcJtX
tqLSgPXiG3ztPCCxZx0f10NuYdWDFJEIIIuvzGGcsrckSqHJEOYOHLZZ2K5c+KYi
YHxg5RknWLaQPJ1DVOZp2KqC9rOqRuoOyud/n23gmxfo+7gM7nHZCfXPaTyo2we3
xDq5ef9uPUfXZbTwLtBFHpio66KoPLU06Ur2AyPc2PvA0tnrK80qroIvUyKzG4dn
yd2tt/biY64WHX9qRD/1tLbqSEolBovXm7dBo3YX0oP00IWx/27cWYsHOx/SCGDh
6LtqRjoGX+H4dN6bxbep+LhMPhZFR+tML2fbn0xxeovU1DelxIJr9A8euDDHDlI2
TvXI1dhRAgDX0/Jmu61Oe2Va/DxUGN7yjVyWGrRBcpGUHcWy5Yeb3kkVi3UijFZc
BX19ZyEi7vpqmnctH0BarClmpArp1/iD0qHcFwi/603EmgU92b3PGIxVK4qdfBRd
ilXWQrT4Z00zxWsjA/qrZ2FYQGOuUE+y8Fb7xXgcPv4o6cea/sGzg2g7KvihEipK
koYtUL0sXmwiEIeR/BOe7qkfLuVPlk1NSZFLdUNgeqMx3wfP3B6ifnWgEouakL7X
d8hqORx91wMMALayP3BLsJj0wIZoEqZnNEahg/3HYK7dhSYV59ORhzxuQum1pNuL
ZCHfd6By6t7xBR+ObUZmexT2xOR1Q5rYRHrO+dSS05ylyLZgGIxH3KE7KEuyaNqp
sfqmUIF/ecPDa6/Ksbrg/xag8vf7EWHwUlRefp4g/BSe+SupObs26FIxxh5LGQTN
8yGezMX8ac43sK3YoNjlEig0jQ5agnnjWIOXo1CWcCH5mjfGLAQYymdia3sXJzrO
mC5JrJJaBWD2IHoPZMform83r1TsmcQnqrQhg5SbUJTGJX6ncjNbvo3b9KqX/ekZ
nhgK13QieHtkc1Dy/19/J6PWhCswRj5qmx1wNIlU7UsFtaozqG+LjVIu8j4ZatTz
JsgdIIJssfV9A1BFvJrNe3MkuNrhwaApHHlqa/Y/opKxw/zAq2WT2YzdExHRGFyx
1RrSp3DY4vDreTlKWKC4qmMlQwFuiYBzCjVH7bK6kgoDUhieAiAowNQYLkd0SjwD
xOEq7uGD8koaveSbyYq1y+leP1bm6qPaXpwp6Kr/8haX9sgQcDWveaMSa98uTxj6
Xt0s9oxC3YguCKMWSoRKo/qXOPkfN43tE34jmFS77Q9NGhEZtLRB0PaV+oZME5xl
ludfvhEkZdANZipPe2nhh7dmtCgdvSaGlHPPiF4e2eOOALaOMQ5bJmUEEuZ1eSxt
6uQDCbgi0fRn9UHJXL0aNGUfEy7JL4vgyr5jelldEXbSWSurRnVfT0hZic4pVtBU
w2N9MgogeGY5zU7LQlT4p9gctI2GR4YWOwRfyGlwH9BQOh9sEH9SAwUaB1elu2wO
RAuLDDMQdSiJ4HVFOu7TeoZ7FwekXtYnhXGpehrhWcTfx10q9JNbdX/sHU8I9D78
PjtbvMTqs1vCDtY3tpOfCFrqItIwLQBZqpxcQ3zoMIweoRveuY/I/3QP47+WA2dp
/9LCCQ395Yo7Q6jUYr53yTxRltwXSvTXp2eGhi3BCHQA6lfPkj/VTqfWFezmLOLb
7xonqUGcA0TVHe1IUKLFMnf2lIRj2mH2K9kcr+HTIq0wxMD59Q7UN2770H8aocAp
g2RRTk9+HJJt1whtrvh7UtxEBfbjYVDUNnCaARWzJn9QnQlAJrN/YkO6JYTYseX+
1wX6DmOPjO/TwOWOb/SzwMLbof28BT81A/Anb2nnO3vwrShNoHV9Y4QOPq5b3IuJ
K5SUPsTlAHlTdVAxzkgktOmq2rQQmYJFQTF6JCYGNkO5pziew+3dcmuI67BcXpyE
6vK9R2z3akQOSfhZ7R4GtgGVAFKJwXTote/NSZg8Vph2I9MmeYgI+od1iVm4m4aT
bn1kilgvNObbYiG50kkWTMndmmY/ohs94U5VfGN+A5vZuj2P6fZIBHqgF2+RY/Zm
MBsOCaQX4VZ6KbaGmFfuhGN407iTQEy9SxvtNWqhk1iwpbIFpO6gnpYHWBxOfz39
/Gwomf6mVofoF5GwiIpZJ2/Y7AovZhH2gZRCWl7/zGqgyp3IXANWamLqFUnA/5+d
mUwd2hqnNMpW6hAUsbd3lup5hmFbK+DxCLHmOVLa2EYluKCKBsu1oCC6znSyM6tv
P7/0QVig0F3DTgDVQC5V6LMK4Y1IUyZ5oC4Wx1Fkfj0+4Wz78KVKWmoWvdfEz25K
ezaDwLGksnZnLyWilvGCYuhNkjcdv3RWRxzcII1FkgKkv2SvqF2fyfhD6MFnnHK9
7LJrSeCFGFd1754GsdyDoJogKM9OL5IITjVwPCrY2BX2QuT4jToICt199ARodeWQ
M2xzgUOiYdEP/1XmlkhlB5pEP90dPItujzPkxjroXTP+kJuVhq/XiN6/Fay5iPEH
S4733/64JMrBsOtMJQyvr1nbEmc8AYfG5Oy/nlw1AP7ILgBLBDGKvvSsUk4pnenB
cCja7qKae6uemSXQCO12q/gLAKP7VryXeCyJsN6d3tgC7ImauyZ09oMkHpjF2J+H
6IY7uxW/xMmjl7ytU39/iAb+8RW8VKs/7YTxG4zWTewrhQLr31pReUhZW1/BVxrE
88hUQ2lofoAqcudmJo3B8I0Uim6iwXlwuBsNUh46ieRdFShI0GyXFaTpW5WsugqZ
X8qMhIMkfAmpIJ9CikMtA2kwRLAwttG7loQ1Lyxi7wjRgkx75oZR6osA/raBiFzu
we2FfhXJfJpYzNC4DdycrBs23xCy6wJQwkqCM/PwQWphtWX1fUfQAMOpgZoP3gsX
OMPGPUrjP73DbAlRAURDxX5wqRZvROyhH1RXajrio0hlkJ7vOGI9kMp3B5NvlrIc
K0EOUaC8fWWbds3wcI62JdwOnoRUV6bHoVai/JweDnnOSFfEFXAJXNKb42zmgHrp
fvd5Ysst/P9HuKfYWR1UkEO6+yi/2LbkQ7YYHHyVt31eV65L9YhGes1tVLBoxOZ+
ndpH+cKQjkBKAl+z/epDALAHiO7hnFY0dDracjkKUx4fzyAKf5NjqrcqP+qj6Qse
7WL7+UZJfGTxsNMricdISGqvQxs+a0T4UibDQJaSQh/hGPkPE+Ds/xRK6ac9uwVM
QK1c5RebZX1d5RYBCZ0Mjka5scKpPszIBykcNdSlfb78k88+aCbCN89xKuUY/OM/
M9h2UxiTsbNqElcxrT3PO8ro+bZg9mvCF4+Ivz7x+nBsbMOzrHe8EPAW+v1o0cpG
vMwAmBEzZsH2dvmXD336/09k9ZcrrWbdm+5zmb1KYZ8iwrdFNsYJyqHfi34lRrkI
MLqS9ijfp4t2AQcPsjwsp72zK0DO4uXCjhfKTn3Pqx9wHx4HmAzBq0bgQJIkBmo6
ZMgmnQ/N5VTCQZnR1BUWzWPzvuzU1vmu4vQB8XKimHI0UdxbL6wMnuNonmxB4DYh
Dkf1QwBQm6CHSsEhbtYZklzGDcEMNKSmMRu3456gvRBoxBV4X7npGJ0QK8OhYpoT
G0sUsf3FTF34clstvOXkgN+elwuSNRgwS/ohgUwdkNzJ9z3j0TOcMk7T5WSK3FOE
xcTKaAOcMx+F9cCHrr575oVwZ/CTKICMrsrSeVKAfQnOXJh01hZLqbgQGiiy7MXf
Dk5sh+oUiKvlZRRqDMLCaA2isjwgKcR6x77QPmol/I0XA8vn7Q9orEH6lFTphGM0
gS74m1xMXfTuBRf7GsPvjiuZQr2dyXxu46wZ/zY5Jfb6tLhp11t6Nsg03Eemlf+O
FCWZSQkMvjSLz2wufgC3mPcgHmBkq3QCS1zK8hhpH42pgS93Al9ntDc8o92wrwwr
RqNkvHLThCPbVKO+nQWxTETfHKEQashT+vQTdQJBDOqRvOmD5zR6FMgYttsa/1cp
wX2IZT+F9Pai63NrYpvpt0qgx57F5mQ8uj+TyEuc5XsYPlHQZ65tI1hj2c91eCnM
dn1EKXKIgEypU8zSGEwpoiyzs6cx1cPIjhrnNDDkPnLzm3vQytlveYaBC8yKNwH6
qK2iguLXHLvvfCv6Iq9tnS7btUSRFxuk8v3/+zgxbwHe8Khfdnwwpgsn0wsgQ2DL
CWkgVGgqHCOkrpS28SXfPAR+WeDUkhWzZD4MVJKzmE5ATsWaxhJj2XaRL230IVWH
lErtvvvbsixdR6WOleEtPQolR1YNpw2xhKr9Wc4ud2uwodgr3+2xhVCx0UuQCchc
/q/5jxhpIliESQUjOMU4EX4L4ozOES2nrDFpWxE7aGUS6sdI4OwQ/XbIJhEwfUZy
UYy/hwGYCDTJ2Gmgxr7dimvuvxeGuLR1UrDLHyE3llBnOKNOUHgthGCIP9hYLEsg
9leo61ym+VOnv7y72C36miFRNuzJBNx9TzEQypxhXXC02j/zgd2iL1uJmKPZPATC
LPQ4gCUJVVTdQVjm6/+5TLFNbyJpUWcaF6RZ3n6mlgFxm0FwTPMzIV43Y4dXFTfq
FVnlzxeqiAE7EGchK0ewjcAVAHzO3FdNOe9XWBcdeaBk3Oxx1kZTL5U/QjgVwfLc
lNsu7Qpsog9OCmQ6/DmTy2fm/6ImmJAy4+TlvrOVNZSENp5N9ZYZIfKyWIVgafN8
ZLogWlX0vN6KOXPcjY8YKQISGRTnml7IRnoixtg3nrVbNly0lipZyONxTXBDQVAu
pjLN+jklVNczFIpfTSdt56f9t1LcFVzUhV34K5YZD/1WysbPG1scJasc7PTeuOuU
QM4UHt+C9ADWCEXZBMpyQD3Sds70X9ASTapMiXSKnWPttKP4ICcZKU2RMldvCtSA
gmRseFtc6mYwlG+/jsVVNROzb57aIVjn4WF2bifNkoX4Pdvrp3QB6BWhZxXidNVs
5Q+KfC+FpeNahhijqZ7JX8mj1T4Gevsw2r1xZB8NBdnbXh3E3OSbfx5+0IINSX+V
1W2A3eLXmty+u249zAySSLJrAenbb2FH8U3jPUKMigH/X9j9KJlp2A68f5vEsgLN
EoWDYWG7coTq4AY5n2B4kv/8/B9p5KX1m85DfJRAPRobNuOzzlaOOnwH8axixYxR
VoIxkZNSHhlMXFAbudFOvlyDmwLXWkA52gPti8cQpzSAC2r6lgkalL5USQJd0rb1
RqAqkBPDT88HYsRfVmKzV03hf6fCb/00ObRvOsCnE/L5mE/3nL25EDFHQqVPlXsI
nuxNtxICJvSUjxBVkRE0+ti2wiU1FOy1qZOu0UIVlue0UbDcl1O/F9ZzchWjcCeN
L2/D0Atch3i56XjMgFmj/Ro0UxE4nRn1lGtCxPmxdT3wKs+AkXT0Uc+T/Uq31OAk
/OmZcbn5nDysz4QVIV0x8FS30zD7ppPEUAplwGygDi2pbW2AAe5S0lHGTcSIDoio
yLT3+ewmrB3FeCHDHJfyZPTbGE6qC1KCf0/cF4LnxinBN5KPBiCTNifhCpGyzDmY
AioAmI+DVW8kt0N+NPeBnQ==
`protect end_protected