`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36368 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
oDqealYugrOC+OIsTtIIFLhlPBm7isDA50XFCOyVcRqb9Pl3dkl/mnvnVnPBY9wm
ffsctela5c1x8h1ki+2yPRGSp5Tq8oasP9hf/89t+A74mWf6BVojgbJw0cLWM4qf
LeUxO/HZwmqnecmJmvDpSbP6HUmmfLiZUOYH9KkMyjAx8F2SyCCAkPaQ9AFaA0D3
ZZCaSA+1mU0rFHrcyxREy/HzW7YmTsTGUxn3FkR+sgc7kXA1iHxF7qMG2iW/Xn4D
dHWjNvgoQDb9uMVqUMRgyrSEW2N1Y3bnyPYBemUtsWQVK0D6LwrW+Smj6z0nPAr+
oHtszjLNYW+VOU3944Nyk4OCO+mXCPDG7hIa9D/5fKskfwj/QlyjKmn76skO4nhk
imJrz7TtedT1uwCP0OGeBGa/nJRIENQRwsLqvD+f0lLTQaES67iveIAuSGl0mKqw
UgVeh6HWg2YJV+vm5w/vnHVJx4Bjkp9d97aTYJsty3n+2sg9UNVfGBh2LRVJ0GHW
gaYMdUl9zOurrphxiKNvfStaXOIdLPRl7mWQba5KdH8piTFx9bx58bcivEe3zu9x
k47eBqn78ncvYOL51oa6ARvUUBxlVyEmPlTO/gPIeatWZuVzpW9fo2bqL45VZGEa
/au0zykxX3jgJMMhHu9smyNn5J/GKrQqi9j3O91UZMXfObMk49Nq6kFB/OtF/xjF
PVvAf06AIPXT6aZ5+KSEyFlC12/P8Pf4i0/Hob09lR2C1L2etGZrI3ettTOB7acA
dFneqfDi+E1V212jHbOCrHITx4r2pAmb7fsfz96JBv2cb5JvCzA+v0i1eNhdLVSM
JDcmyP+D0MV80MouXB3B4LJ9Sl14d4oNJtKlcWJQ6k+di2jPdVGrMKRrVjZupWrU
AsHP4cYQL9cSIykkKJQpKwyMlaj49k8Mhwj2NpxROP75cEWS2loR6xetbpBYByVM
DwFH+KFvUmxYsT1wCXTjV+XBwzm5gTHdUKRpK1MM6qg3+j4tG0YxEEif+4vh7mQG
kJNsXu1zUlXWPxhkFAxxBadsk/a7RFYnS+1hx7wgJ8qpJlrz0KxebUwzPZvgeoan
sbWn9wHvlgdWWpnJeREKTkGTeppd3Q8ztwmtpLdWO0Q9H/I0ljOeuN9bUIxD1CkF
8eigKMpAR3tGAVwhwT8IFWG6xD6F2flF/3oCGGvVNLwMockkgbB3c+Et3M3ndpbD
R8VIoOaBtHU+7bju06lDEqZvmZK5gJJjQMa6/4yTTUmh4f/uT8qwKT9naQCj+lrC
vRDHl23/H+Ni0aQpEgzyvUkyy8NGr5gnE523BXFH9xLU5hEhmx7VnLWYux5l11/m
j41UeK9q/nslJlyA8ZhffZ9jQb+fLwGG7VVNSuDxxrErqJ5B0Pjg6ka9y69F8ZAd
REj2meYxH6yGxczLpXiC+eyi4OBeCnIbM/rscQzpSaN2k0AwXGrHXZSM8EzqiEhG
WrjSzDo6RVYkJKVbJcZh2HaPACOWITE1Ap7iFmmjxJxvOoHnDEFfbPfU1TI/6x47
HVX1zQI79JmnwWOFufMUAXA6Jx/+GEZ34HMk08jqNW/zX7jOuC1+W1AF6L6EDyba
608TbcBBIDGliOBzbRUoDVQq2Gx52yyEKuxYX5UfH0i80xah2K6K/5shMAFt4V9p
CxS2VzwYF14+l5axO/DkvWDpGaEDy3Z0qe8EwJ09aEnuwIeaxI1frK+372lWxHjX
aK8yYmFwQmFisWR6gLbKptBwNgz0iTlsknLg1u5p4qhnh3jgsMhAkgvv0m4sNH3d
dGkVTlROkRTVwfaSWSRX2U0rNzZzE0soc9oi0A3bL1VeqNYBK7cOiHZYbsHnyrLo
CCHgiOVct5Cvu3G1DEUrCYVCzQ6jFvrH2bHgggPd4uWn9o5PqFRzTgGU7o8ncguB
LlfPJ7HiVDweuOpklxqtxl5wifkV/OAACvnEPPc3ZfhpFI05J1Y3IJSWqthQ/uEH
2Y9PbULjEsOSUSkIfEHvEcFnGx7HzS2V1nqhby1yzI7+Lu2zAOaXYOKhbc0SznXa
hNUJNTmTawgBZnBrryV8AoqpEMoYLP5PDYKKcUikNmGBiiPnafZgbTZTuqEG7QWe
TWQU29tKV12tSH36OqIQCzTW8XAc+UX5Pih1egiaDwbetxmYxngQA3iNJooBR3TN
KFW3KCz3qk+UMF8CVEQhPgBmQjf3+iPzt4syKwJkqx0pqgBcWAcBL0kx4hr7/Lo7
yEYxCagX93UfrmyDQh/NHtfD+IRKqP16gN+bPrHZdVlGCwuwJceVBiHDIi4TRRQQ
boaJwbTOPOlHPuUneAYV/DLXgU8IwwdBx72u29VOJ8kKnLNp16uraq13TzEe9jbO
nIkB6epeGBemZvjUJFxVL0qTn0KYGL1sU4ZX3s/f0ShL26gAyag/PrARlOK5BJEA
vJwIOw1lKkJG8aB+1l2U0H69KvBonvQoVAztlf2tKKQOYHWcxcZYp0ui6HdModH+
vo8MNNPGTB7qT6+0iFmX9I/qleC1JsBGF/AiBh/7pDLxt3S8kD+0bnJKQby5GsZv
C9B9E7Oeoug9Xu3X9ryOxslh1lG8Lx5AKIIJ6X3x77qsfyqPZG82yt9ajG7CnnKp
+iK+TKpPKZK/XvVPSs14femjWQ4d3Mw9ySJxT7lIZDzKr3AH2RkU9FVVdLbjEW9o
Ztu0yyPaDGgkKv9GoNYFh86eN4H5OCoizSO6F37RrnkT3w9gtNN5udrOxj9DK7FE
cCzzcFPzDRmQGvNaWIhjnJxDpporKfEBTUGSZRotE9cQhisB3wdQqnHWIJrJ2Len
ReanAhtRJpfIInyFIGYYBSND+8vkyAFv2dCVfEbcSrEXnqs0izgXaS2s6aTQaLwt
aFgi7DJqyVDfuuof8S+EbR9qm/+G2IVLtiLP4R/W94VBPXIYoIV/Z5oceGRLIZ9a
YkzSJmZMN5Y2HvH47u/pV0mrIIqELhAcZxKTSRbi8w+9hzQANjMg0Db8dTRYehXI
NUnA9Aufx9Fj+pAD5akT+TfyBsXRifmJL/YiZYcq/1AlRCgNarDnrKTm7h6ohBZY
tinyU0MaApvSs6QH/+7kcpwISLZSUopVkN2HY1AvVZyblYGVB54/iWkd61GCLbMM
aI6/WBAosr35FCxV7kHVAe6D7v8k/9C10ZAHRQ+S8b4cw8+jyNV/9BWPdmi7w8s2
qrLk8YQIsjLMq9lrFS5Bay+CX9CntdjGNwYuT/zsIyW/iaQo1YYU6dQiCrQGKXJ6
3KLVSawS+EoPettKG5R+MD623MFEsH3UyoFRgE9D4nDM0yGOfRhG742MKIiydoKR
TTmMIDmxknIgzet+4ezND8tlP9WVROS+h4LuIPD0JIUQcceR8NsKiDEv1KXPpPsI
eKo9EU+X8WJZdmfqZhI40GwqSEJExJo54PQX9cpYa38Fof5R7mmKZbtbxjyecfW9
Bx+7cb3s26omTQWDWP5Vv4faexuYcmHF5cPm5VYe3S9XGUVFZVfEf4MDZ0JFZJJt
ncey9rCihU2b6p6TitNHn1GiBM4GQ31CRskW86BnOard0sBkjPAb69NZHJe9O68p
kz7SSD5EVsHB5T6Yz0AbrSS9vlnkXK05fxDThb2Bsy6Heh7XfzCUipkYA7DIi+Fi
cqxhfWYYSFtTHY61A6jLAR26fWSbWF6ZhzgfG1PgEtvVZBRXnFyM+UscI/8vYWIS
N/A9U+GtUP3WJ6iec2p2liygo3q/wXArcsBK+NDU0SAxRho607A7uMMT2droxUyh
scx/VkG9MbE4rbvLUNzXcXIxJhOj4asjLImV11p54M99X/HUexQPmzabHyeaxiFZ
rGxk4IT19WNC5lO36whwD2JC6HS+OZDQRRCexwxZVeka9GCqmIvnG0mOEVtrVi5J
h3ya+JH5ougo9z6cXf24F47R6AdYKL/ngvKgM6IOpkTyfsxUvNlFf+TADA+tnBur
cqJzjRhkm1OOcNp1ix+Y5nBA+0ns96u0hIzfu4U8cyg0hOebUQ4vXiZMl7VSa/oD
eLH5+siXyb/a+4U5ApNUneZ8+EB0EAUjUcUpwSZFxTlU9TF+AZKDwWnOfWVNo0RL
tsELAg97tl4h2UR0luUqKI0LkTYQurhZHc7S0rljZXuINcio/Bt5Vngo+j87F+yA
OfSGf2sVCe6YXjkYFY+4ySfKhF3HXNPS7tY/V3ySAUe5an0Z671yWUif2Gb7ykg4
za3o6JME6k8bLGFOzyfSFu8dmuVT04D50uIpoZlGMOkJUluQ79fHA3FkJFEAlGxq
pgLCSFGkWU/RmHOh30aIFDsSUMulfy63Vf+gL3BDHTNdooqk5QWQTx8pGjAMk6Pk
P+Sg2hxDo3nO++LxWEbqWwzFHbgrG3DMUEoF41M5xdGYmiO6P895hVr9+PNlLRho
BVX9qt1nMWIrLak323Wha4rwbfTJQNNonOQhsoBPxNA5S+gLL7mVJJ428IPbf1fJ
hL38DfXbS3NYcZkkIslr6auHifBC+/dvCPIU8FRrspOLT/3Wy3TLJmHYs1iTof/Y
gyuEkdwV3f3S9NYTmxs0dzfHvOxVm+dE4mwP/9aZMSGx2XdzWjOb7e1LhE7BfoP8
9xAaXtVZtRQkozpS/KFqD2KGYI8InnxUdmD3rGuTaeygpjNkDuCoyVtMfNsG8xKQ
Yf3J3fCyJj8kUATdJn0n+YalEFPx/3eyJG6J2VFMAV/Z7E4ilwtWzmBno73WSfne
NEYTNbPGmmxBpyMHKkGA6HtoSpaMyj1Pfq1dIGVb31bNgoPpbkVzn5xtfoOVQGe5
mM966ru9HISENuRh+jFhHst+n2pxEemVVt9ffjRnFfchtw/ruWyHV1r/PJDu5J0L
eWVQkYoJhW6S9FrS6LuuPfuwcXiTpmSAIcu4X3/pgAKFKya674pklscaTi2rOb0+
HBxfSIFYNNA1FKcsvq3UzkCZmhB5ofUm5UkFEmJx4zfTIdP2mDONVu+9tTM7osSH
NTy7cH7XJWxTYQkH453nTdTkW5YmJVJeLAM4nr52NRD6kheeHRC5WVI1f7PGTPzb
BGokV3imLXALFdEsR1evvavcNEShM2J3PE8MNkd0UcsiXxwnAUIX53cGc0KAAA2z
rP1xNRrQg47NvAijjOKxRLmq+uadytfTNHJ7KuQ6Mdybs/M2ZET5qI9OrdT1ayVJ
2nX93tRxtn4oSeZ7MvTnxComHiUZIXbpor8Qo7NZnXZFQ2i+wO8L7zzOoPq+YOrP
gXnfNpta2ee3dJN8bliRjqv6pn6fupxj0vrmsPwVlV1QEhm0Vzw3oJ0TuznfTY82
V/egH9Gza4vnwc1VwwiIGmwGtjdMdY2bcltpeTUeebueDss26jcXF1gqSTCDqBzq
Qr8sf9WCapmnLCQiHxeI/8IjC11K3uD9G8/deMdcMvE07MURd8YikS+2zb/NxYCL
lIYlJBf++W9ZvO9NfA+PWBZZr+YkeBaWc4Yg5q2esnE1f6bRx88PQGD+1l6KLVEL
TPe3loyFhDN5DcpWw++nMINEtOCL/illlbsri128DBS+4xRwQKOZ4bw9ZwnzDK2p
K0JO26Y4f8mlqDZQh1zryMfhtTqhGQlvB6S0OE18i4p70k7a+w35CzPUc5Up7aMN
fIJm+PjzOzo4ir+g9a1D4Tn8RQn0Y3l7u1TCQqARfTTeT33SNxqknL3ImCPrniqi
5zLFOcV3YpAWDrQz8eSMHGt/rKwSX8N92ybd9rssQ2qbm2S40AYCks7HSinY4PSX
llnnOYY+A1I2uqEsMNRQOIz+y4pD2+Q2AumKGSn9hl4uM9++It6vHyJs6nYdw7TW
DgNPYmuH8OStYidrfpsvglBEm/OkEKPj8jnuIUVQai+kd+V3d+bVvhc3Z3xUig8F
pwOSiRh+wC/oqiGyxSb/iWbtzyQesIX+gGtO0lROyXBSwZjLn8h35mIrOr694TfJ
4dKKketL0drdLlG+zdX7kRugqrlvYN4UL4Ug7yz0bLg2eru01KwS+Zlodyp6OH+z
9qGH2WMkIBmthWbz+EVJJ3axT0zvBN0lNU+vefYMGTUpkgjOW0cjCWdSIXukjDD0
k5L34PMPEr1VTCBMNaaJgyoN8er5GnRIEgjz/R6x7XQcpoNWUpE91lyspUdWIG0M
Rb/Exq1QPnDWG3mYzi3addnct6H0Qy5sfgppvVz6pQ4bFfAB6Ua7mUx39UafD3sC
ZxxKTvN3jY7dJNH/sVelM7/FSUfjvsYAOlLCbBCA9sS+EIMbAjDFmbBBnZrNUE8O
epf3otl+0cNu8N30zVRP752nIt0rTjKKPRx9q7F0tWoDhRV0oKXnFErwU8jTvktp
aDuuv7/zWH/libRqRwHXZGeUFArGhKaWsTf3cJexw1OtC7sWvdV/926zP6l8km4y
B1g5ox3pXIw2rv57qDehHk1jv1aRZKorJeIjM5X7t5SIocaGFLiOijH3dyDfs8M5
rl+cDVpM72lmsh9aMyzic07hG6jNFsxtAtUmZd7zEcVtJ2bNAwx4EO/G5NY2p5m7
2TPRY4OEOrbkEZyeFqjhxdR0dwCuPq8+Thb7/7SvFd+nZl6NkTF20oECU+OmH3Tz
7VGMLMWzBuohejI/FYg8X8T4CsS5MpJUOjUxMzHd2ibTMmvfl+jPJotb4CDm9B/0
0q14CpwcaILuN5NG0NAxxgEOaljgcTs549QGBaOWkoLzbp1+lK+Zx3B35dNhKE40
jaXN6OcJN8R1JwsJTiENi9U9FILhlwfgJa6pd37HqqmLH6yvbtzO2OqASYPP5zVN
icajvqGy0PyS2TeL7Av7KbJghEacDE7JImNkFhfjeGEvoqnPXzczg8iZa3hIGSM8
8zzCiwANYhaoQLcU5WAZc0jR5jxnD3maca9OlPIgPfJ4rEemNpN38e1sWmMzHWF8
PDyBZz8K3PSpf21s3hB/4aVBXYgpCHbv5+RcrK4ELt4JCWNWvhsFTtHDhDB6J1Mc
yT0nu706vy1LmEdkw3w+HD//kmPq8/UNsDQYHFHnCRuMSdlu2C90SO+nvTjkDFGc
r1XPPijbf5xY5Ms82eOf2oq8c3mpFpsyRo4QckUsd9x2UCEBSa/v2z29I/lhQZZ3
BTASh+5J9877Vpjf5NVU/z+SLk6e8aqmgA3K+igNcDFI1pSwOvg6/kVqruRDkqwS
/uD/MB3tr3TgfRhkst9rFdKfKj2OGjik95f5RUViJeiIxjTN7L6gzTwiNEWGU/Cg
CXmc1d6yJTFkDoRmsncdQQ6KiiwGdBd9tvrTYCm5wWluDFiNq2B1cDVW89YXLWxo
pWMK7nv+8tPx2SUg7UDQHyvaroqqd444iNrMrGkPJuA6RdXMgCS9EeJ7Xe4nQ46a
1O4S5304pCCAYupxmDP8bAIz702LZs89V59/DRzdxeYSoXlajx1sc+tm7qnTkabH
gfUvv1+z3Hd1h7BPjxlckaWBE47CGcG9OgSbxlO2DlL4SuChdz1Lg4zUdkRniEFJ
a4ebELBNFZgg0RYw7aaW6EWSRUKi6sZsUV/PuOFfsP6JqFTf2tooPD3WCl+3T4LU
PMUtwlds5XZhvOvn9vTeqsm7MUwrkoAO7OacHZaOHUSdMrbie4v+NgYjcx6VItwJ
0UtfTIG7dELDC/UIsc0v7JKPefB9hz8zQsZScxEYMroXf/sIHtpL27GRuk2YsGFA
635y1kzkLd9li4/2/OItZo/ZNdS3BFXyxB8AabqMoBvbVOdeq+BMBp6zIMMB8TCb
bNBgpkTiii5FrISz2mrnD1LesJqMZpcrU8pfKqxZ8l+kt6AVNv/qcqGQqas75E80
JqQHhTSgpZgGGsUAIf89BDxo5LG+QDiLvcsgjgbcvG9kyCFmpx+6kodTmF4KScPo
jP+9LZnBaP4VE63sYIdBMcMfxlWm6r9118ziiujv+Y80SES42yJBpKgPesObXIFb
0HFzbPuwCjeWhs3Gpv+w1/EhqbEFIpoIjP0AeaS5hAgjGEKPJIzles6SlipmLX1b
3Cdo/NG/0TpUqBv3DpukEDhWi0OHZ/0pCyn6szg2X8HtOo2TsgkcFJCjI5qLgZTA
uaC/EGaLoSEIHFrEakZzriUruaGkVQbpqBuo84hV4r7KLK5iZPpGXSVWqYfzyUNc
JRxvm5KCUuu01ySKGkfzF1MzY3rwiSeuxENWlRi+6k37BO4OkjfTT/gSkBEksDf5
iMS+Ur2BZzV7O7/4YOjVSJNFIc2CzKHDeL2IdUOnXEyGNYSdyH4U+UbY7mbob2wt
MN1cu99ykwYN28vxd0SfmlZBIqAFyFMplo+Lv/ckBiQVlYyzvn8DGFrJrPcflfWY
ew/wc/L0BCjCtUqAfFfxkp2nr4YjenwdHWOGTRl782X5gh19Wsa0+n5qepxql07V
5LY/Zbq09J2fGmyrZ66ftnqvY5RZBCQF429AgKkjswwDgKKz2heWxoibwcfm1ORq
skk+T8CrTIOsVtIRdIHhx9dKFqQLOpy3PW8BdyBeJquTiHIHmIfxMrKh1bmLWOoR
wzaYNy+9yd89EDHZCrqp8t1ApuQhcA+ydTn44GN4qPtl5ZPnDFaa73TJdeb/BwaF
wUiDkKMBliW27Oft7mv2yJXqehoScx7W7WP9yT607wlgNevl7rheaZLTu3a9CTh9
6xysqS57ulcyK9bGBK5ATd/zQQdNq5KQELXfx6xzOBiaDJbYw+TktjYf8ZnnyplJ
ZRDYaw/X8/LiLsh73DXve+0uK/jO1DznbqV9+2krO2n5I6x/8q4m8y+uVey2K+U5
9SCu20XWRFC3XpHrwroddLpe6X3zwGdGHdHGAVbfCBvgXiekLHoDzfj8vLn9ml6R
9EPsJfop0rmm2/t1bmKcenbHdn6Kb9PFONgEKsHC4At099PE8DtFZgBwzkLfBcvI
xgCMVd2APuAv/X7MIcbwOKLYUmGzNLW4ClbP2P0nugUCUg/oAU65LUG2DaDFFpmR
g5ws7NR6oYaL/RY5KxetzDv0eMiAePPXnKLo6wATFlioMuWILhcCZzXgfU6+OeSA
ULJqlnmuYb/LJzrPdGsYFv/C1U6nYnWckRZu0e+08FdtQYqaAMydcxEhcDTnc3Hf
X/eRktlU/xWrWNAYh7ToI1AIRPXUi5csN5Qnh0KS5q6YVSNG4vEtkLO8CJ3btdVf
Rzls6w6NjbemEEjfaUYybi94foGTjHMro/PN70bydyuFRRLPBKqQ7RIFNLWPYiYS
e0a6sNhM2DUoDU9KcrCunmEh64vD9SBBQbqmE/jlMbvUVYD5Mvcm50rgcSpj7gBz
uuCKeaRjVb8oftrmNZUCILlsT90M/emHDpTyMy3/rOdhMd96aaeuLiIeWEShjlSf
vgnKLin/GMOWywYn00XlkeZtcy3UVf9lh/2YBP2hrRwu+ipsaAlkxoXOg4j/+Wob
zFekwjhj5yvpQrjrrtSYhXEK3+3fGFF2SYj0Q54XK/ghAUArDakJKce/ELnmC7iF
WXGGVVBky+84nc6aU/UVP/Ia1u3oPD1gVAtAvelSdpjXcqSW7k3rPM3+quUUr3SP
K8+2AXQ2sN+ulUI2JLskgvK7tgO2b88evDkEz+7Y3g1IK5A12sKiqvVL1fdTYm0w
gpg0jBcM8Nzo9LVAK3lubr+G++T5CshmXu/HznOwPUlQ+Q4JGo8uvDjBnfQbQPeA
FvUILVhXR6/nJC8yyMzRC8mytxGhY5Qos8jkTLq2MczunvtdOZsFH7r1Sc0xw0HZ
2uJsU4ZVWRZ1Bu39RJ9CAY15su00sq1I/NcP5nYLAcS2kLq/ShaU9/Uu21H2JTQv
kn3CN3JyWkZsO4b0VUH3rLHFHrCT+Gj4SOqxBwIpgtHy9OnwFzEKSWR1etxqS1xP
UxkDH1/s+UQVpcp6L9NmCkH4X5uqEkWZD+jl10oDt9UyX/ZQwB7TTqfzXmwH7bkF
3iH6asTHj0Gl9rSdmqwnJ8MqHRPI1gdPxS6UhUq0Dq1ru/9X5D/8KpS45/MkV7HY
WvlGbEdow1G0x0Q76R9LNU6catsjbtu2Sq41XHKk0UnzruOG+b5p8Jt4z2RsoakC
14+K+ahrXQaefhpxOVaO3tv9KqnJ3VkESAGFP9Zz4iVcsqwPdvn4g8zzH99DkCM7
aRxX3K7XIfyZE0XTv5KO/59oQPsu91m5Ek8aHqHTZYDrdbg/j+Ofj3SKqPozHs4r
wFL9BZfaH3fs5ZioMJXKbBF84jgh/kJEL6LRYyJ0efrmXjuBbUc6RChtuklhehPk
s7bBvXmUWPgVCv6uR/mpMwLI7IkbJ7pa6FKjoO+ek2KoUhYhkn+5VUPNCHbdAX7L
7oZ8H/nblEicZiaK3IzzgJshehSKcyqYqEPxIgaxEBg+eVa32ii8Eck3ZFDoZpB/
gTjmPuA8nQ6GWELu4OLo8RrPj+S9dPXS07DGMdlyLwEqNTALAyBFXPDhB1JJHOuH
zqxg7rMtD3Cg21img3/ElTyu6WBcMD8CGmcostlh51ohSVC5neu5xgRaJzrCoySN
yyVPIhOUE7Z3c2NhpyloY7dCK06C3PJgS27AbeaImYQi6k72lbufZ8/hL24s9vcT
KEqdnWG3qg/GP9B7NLcYkKfbPW2pXSmMWpmoSLldH96qARORJFNSC2OqF/hhD4K4
biS8tAU4UqFmm2cn4fCF/FGO9SO8cipiuyBDZjKLadJliRelM9JWTQ0Uoaas8mGE
Eu6/otsQzig4JIUWLSr0a+hdXHbFnebrL3flKq8y81ulgVgyMTuKqjC5RIy9soCR
glIbBiy4OfD6ZlFl6Gr0h9bz8NU7z3PgqAJvntSRYNXzUefmrjtayD6nwmB9SItG
TD+NJNEztsxDQLOnlr1C+CLUyhJtVC3wb2D9W6OBTmMvaIg2BINxF3trJuJ7sPYs
CCmHB4LlAIEVkKS1CrMSR3nucIZERfn5NL3JuV0AtyC1aPfguXle9lYvY7v0UkzV
fJzOETYx5AgVgRniqSBI9fkXckp8gYOaE18mM8+lA8s1b9Zb+PGwafBE/aH2yZIB
P4UUxR3cHN36zH3ATCM2RKI3TnONbeE0WTKskgqtvWE/NW78x3KUeCjFQvad8i+Q
WUMD9hU9TucDmX4TEKokPRqUhINKIYecf7IL+YHnB3UPLk7PdoJ9+nDMKtfcR4Ak
+FX4QNZtinNrY9Dpo0UansH02AxKl0Qbr0VkcWDePseZ9tRu3mSU+LxBgDunwVnN
Bte/y5wF7XmK0h2UWOpq6H+irVGBJgIhh44tv7uDomh51h4OOHCCmW0LSGXQGxMy
nA57EwS9z1tVcJLEljTbMbr7CotFklST+CQZ/isjWr5JR9kBeemz/3JPewEZe2Xc
xJAu7Vn+XxROrP9fzQDQe8JWVY7ctMT7fsS36F9kbODHmtKpmu+gfGEKX7fFyyiV
bW2ADE/hf8I7OnShs6B+DDIBIV3+iG8XnKzsZZw8RMlyN+7y8dvlm1sZKu1aaShM
Vsua3pssTRvt5qY1g+D+yGKwwkc25GTtYGjnRUWJsWBq4z5kGSrVOHMFzxIBSUHa
/Rq+JOBKC4XVelKNgwwzGZCUe2SbY6i1a36OTklV0DTenFpxcgTrvMgCizfGIwIQ
dzCliWhs04LaDWZWvD7oDVZuxBm4XJOsvfNzguknhQGdZ66B8AJzkz3t+ahAFL0G
nkhBG3hkZrBvPhLXn7wTqijPASIGGEOoOi3QjRYBVpPWamYoCg5fPwfLgx6pkjoL
3/zLNLHH4wflGHYzdQBHUxmavhjtFtJ19UTDsAsbRYfspI0CylMJtqQEpzK+F+Qv
9rwRvGYpV3M9eJc9mtfxmqg+D3ZF6N4bsbxYiLDIB5UejLsNexJi3yuyqU5c5Z75
j3ulDlj2RLremolWELzj6zym5KK5oS7a4QIgMVGNbyz+juzCKZn2fb6FpJEKnjx1
Do82jl22ZCdyW4qMFWRR54HNf+QpclqbsNjsL/32z6Yn5bbr8o9DJm3dqldAUQkK
p2yche3xJadXyzHDbjt9j1KinxoSOCUIIDKh3mkArwXRD9o2YpcCyJQPsLDPmw7I
tsXcsvGYcfpjiwIA8XBwAHuwEVuADZDspIzYcM4OaWrpzGjYyk5+eQq85TsyZ/1U
HYV1A0xvGOoF/UmH8Ur+ajnxECphkL0EAOSoxdvFpNZzbHuac2dzC92LSr9xlduF
VdbCJcrRY7LL+myq9YSb0IaxZ7Qg51RrSkLEQq0i01uIDZev6htl5koleMeHQ+to
twPYrt2/2a89SEE8aZZ/jnlShuy8Iq96GNlBW2ghoi3Ai/UH2RF6jhEFVdiUHJyD
WwFFErabdBYoDVOGuKpTox5p6luyBWNcPr5v63Ttbp16QpDD5m1kXZCG5zOwcHa0
+MkOshK/nvJ97W/eSvgbAw+iyRWyGwyDg/L6FNhyYd6QM2qfbhb0tGCPJv3JuWhO
Rd+iGwNS5lD9/uzXbb9IHWY2UiHLktG6v5zRpANWbNkKev/u9LprMjaH9w4TYB0n
zfeWx1jy4rkMoGpbtHo/I2ythEnZt/sGxGxB5nF4C1pjJxGWwGHcTtuhzXU1LZbl
RkUMU6Ivuvh9mab0X9BjQRXN868e1gmHn0IgtOciRz6jWDZWDAs0jUxg9fe04z4I
4Oye+N8wu1gXH41ZeCGlSyIs934WdxpXjczlq5MOFZxxG5kDHe0y87SwXyvJMMHE
Gd6eIRhp+g3uRDfPTHKfhF2OWo5fDz3QrZ+GkuQuB/yN7k05pKa66+XH/W+sKpQf
SbW6B1WF7LOcGszKmO2OsDvkNDKbNCaWkMOlOF8XoMDwImV6BjhnF8QtFiTEcFCp
GNJdwyMqAu7zP9lW6nI0WPKxYoYjIP3utuQoPMdsYZPIHZ7oJhDjtovXwYhdJ0+h
qk/mhNZj+vOPylrilzi+HioXMisNZMlMgn2yBnTWae6JfudBCg2iz4q2eyNVtsPq
1OR6mhm4lR/wBXUvp3TkM6AR1sttgkWjHMoIPVV+6sqhRfw2BiGMzDlEEd9k1yP5
DLDun9g35/dvOMQ4lFolNTVSQmhwv7CNItOpga7x8uTTSxTkq9cEmE2/P9vSCFGz
OLlfiJz/xknP15xOYKCbz12PkbZz2EvBoHxTxSbOY2/tMmtstzitZiasjEDTMZCf
6Z4z4ceuTqzG2nRfm4cN8A6DuWHxn02tQOzdSbvvZYnBLeKBsO7oCXK/bNUCYEnx
D+576hvsDPLncCbBzWP0XG1Ti9iQWg/bn4kam465TiLMtSTCWZ1CNNLVFxn+Rz6h
cSBKtXACtjDbkDu2XTwdpdSD3Qmo4SMRIpmYShOK7DDLhSdf9z63SXh24uHjXyTU
A24gYgapcsS+tHS9FzrJaktWeSqaNOmBM8J/haKj5S90vQgCH1/lus1rrYaDNi5n
Cr36k3CkMgSgmzP2lZf/4lteuSFX+InbeL0mkYoLMRXDQYYcEBpPBliOuUEXTQbI
gtrJjFs4m6KaZDRfrSZLQ6g9L3WkOY8mK/d8z6vdSSBHR9quRE9aZGuxsmgTulte
D8MICTx1SNnTc55bZ8ZajgjbSrMkdVm2qKTxNsOXIPvGw8NFWHXWmtcpOgV7H4Xa
Efqxv28MkwAq+66VhRxmbOAwJv9fCPQt3ngkXV1bAbvqpz/prxg85pj+T8LS1/k9
qBwq5bHWpcLuMS1qob9VUl9CyWb/mTndoPeSoKU5z6lSaktuCAL9RzqIl8PLkIRN
BEN9pqajqFPUEZePY3DcmWcv6g3o4q6oRr7WW26G/v+B9LuCF5wSXuImAJZ0oilz
9pnztB342OWJplZLq2YH5/piRiL/mB0Qam+X4SXveVoum8uKg6KqmbVNJFCbec00
AqK/3bpOhCsO74G9VrmpVwJLHih01UDlVARm2uYfrVjjzWsQT0ezYKkF6gHLMH4M
dBcIkjCklJ3NDPiLYE0dK1jEepqgJ4UcoDiedr3fPhsxb7+TZXcYJhNeDGRXIZb/
9XPefF7wJlwxOt45Aa5TwunFkbXccd+aazhgj3hf/EdyeXrjSKNCpX4zsipBGSAX
31pZ9OK53PRHGGbQP7g6z1deqg02t6GTwBOPJIzb1gPa0sERCMr8bs7xWnM9wUhT
maSMwj61vNmQniMxBbbkC2gOIcQrVrXivERVz72s2t+MKMMeRSSDggBtB0wt7akl
TzBMob4PIP2qXez8B9dn9WGH3a7mb5amRZ7nWiUO5FkGz2+Jlk3mYWe4ZC7D+4pM
/50YMtSkvaEpBjanHwalV8Zl57adxyc8p9ma0Oi2x/ot5cukKUyOWOJB0xRlE8O7
+3ajsCjJReO/Xcg2lHNHWPP7sqkIj2KgtS/7AHO092KFEgJS1czz0pc3O36RoP2K
kQ6CetfiZlJEJMEKveXizxNZA8bRMa9d94Tq4M++lhSrE749JR++fh4vX1PPX7ai
vMa+pi/fRq8vjEsbYjGva99JIbJ9yTzYbQ8lDpZheNIMJ1hBQQp+mGubfti0B1sC
nnjWjcJkhG7Kp3toqyRN/0Ilvt7YrUnbdjG5wvFt2K8cqIMlvUiugf3MqXYLtgMh
fPsmquBL1A6KEqcfwSWUoC3C7mcJN8S3h9P35YKfpeKUnkLO7yGws48KKmSJtknz
Z1Hq787tYOD1Y2/69cucUMNlmIzpZ8hxvO0tYdBQXkRbn/UhfACMiImQVzn+DuIK
XIhyd8MUicqAp2FUvvGkQasog4x1yJMRhNGHlHNOIu7bYTsW8sSQBwCqWTBgG7Dl
tdq7O1mbr/+bBzYl+k6SgScBn0YzzJDWcxS5AJ1TgIrse1HpEmzM0djzrOaP6Cv7
d9rVjxVqphpROiGSCxdAREC9aITKKYwMicz9P2kACkK4AboFNlLVEe0VNQiW1e9K
f8OIZEw5SVHyCko2F6TLrRdDkvAEOQj43Rrhm+2kSPfMeNzi6BWVHUUTmMD5wBjW
dT7iz1VxC3siWUPOXJsH6olerrVlqMIpO0hXPMjZX9K44NKZ9NU+MajNq9EY0AVf
CG5zVKM7w3y7HDTFun0UY7Qs29W+iBrQCQ6kYmLq1tuo+k463Rzv7fBQsD+0Ce0d
yxQAm0ld8kRa3yvFPK12JHJyOzVqACJFCOwO+eQMFwKN+lKmTsFopz1SkAqQBT0J
T5zzmYQpiWurd+nReqNwisIrolgVIN02DHQfYXHdvExhHuGUjQvlgRfYEh3n498X
paZ+CIVKu052aEZBRvULvVf67zUs4qfWRPvLeQRWP83x+QuhC5xFl+HCCQNmWXl0
9riiPViteEYJXpR9cY/Vyx/kWc7pubZukfdxQaOL6ka0o2mvd/mGwK6y0I5WokcY
L9LZL9+mXttFWe6NUIk4tJRj5moh+DRuOwL+HTVCUFJWa8Ai12dW+DmPzUL3NfHt
kTJF7GZ4pBlndeNDWjeAjR1O7vx8tyEY4WvoqVYzFrYitfXh6uH7JW/v/xbGbmxS
BxBTBLMIubzj7Tg7oT/wt1kqtawnXlKWTkMJDjJqO06JE+m2DywliCKMT1BWnD1V
4p4Fx7tLxgjqt8+3P7NHP6ys5kzzmtyVlAPSIn54fEnQeiGHOOfGqZNM+vezUHVL
5vpOCaj3FWIt+me1qrKN/gOWvgVYr+MsVjZUp4D7qPMi53PPnUsnPeFqgAYSWqfX
k7E6VkC3PXziAP4DHIIYrzG0VpHk4hJnKVGjlgLTC/pO3+IEDPLgi8O9L7nsuirO
2ytBcDb3luBm8eVTZ92pxYoTEEJWPsY119fMMQ/jb3X2eamqCqTJnEA1VySORWZ7
oUlHALfyor73HJbVRnYyoYi+g3OIKSWlcbaFDLgDrfF62U2rZrb/gSuY1V/6OY/U
mYLgL4aOScJJMcEcrTv2dOpM0kMyH6sszYhkFIhv5O9vLgATNkcZ0En7/4OC5i3K
MsBDMLNjOvQpiA0kfMljTZXkSY6pdWNeQno6Ov0WpUYG5WZzRGdLZZMbRrssjOQm
FoW1tDr74YNtTZFIJ/oADHMR0ItB9io1wk77sfkN0vRcmwJPuwZnWVPe+C3S/20L
+HZglFqnrZ1rAXBfDJ0j+NG5FLklMbpP4uY7kXJt9oEOKfuUXxtKZYAoxouZMDmd
KvkEQHLlhIt2pDeLUCNcCuD2hN8bpOXb9g9HffJIQcXWZ23+4Ev1m3tmZHw7+dQO
4S/4YY8BZEjLrcbmBI0l+wQwVc8wWbGtcnih+hJSIuaQDL07QEtXjxr2JcTO/gAi
0JVVoo2dKmJQDuhAAxZO+3hciXsR0R2wk7eY13LsHJj/ItlOPVNNifQzAwUDA0GM
XXhuvf5VtgoVWaEfWg2JKg6OzOrvA42UAfHkiohL3UvG+grDj7fdFqXf+Q16K/UB
BYh9Q/gVJmv/UL2zoZfYexZOWhJNPXAOH8FUyoK+I+NzyHiC2QAe8PNkpF9GPm8b
1EhovszYPBHpYEDza8NjnDBpzssoU187PlvTuQKo4805QWtAzBR/Hj9BO9QQ6sHN
p2gpDz+n4Ks3RBsTyq/cLrQ02Z73NvvuipogboEn2K09QgFjEqHojmTVXyvlXmeL
tTYaplNSnzHhW/liDl8fyJ1EgzT7zTiDKeUtZn8JLtub4s9qW68y8zF1YJpoIRmg
X+QOiU54p2BJ6j+nUR8V42/QSkEKFgw4lz9NoLgwCt4cS/emzV8N73kbxU7ePUzh
gpnNYJSJDDCqd5K2hChiMVvVcofN9IQaTUEMBOrkilvswdMXPTgmEoMNr5UgoQVh
gxkMKngKFyR+T/mLV+a6vp3wUKPvjGur18op6gq7gQzeIc8YAQ5EkXEormLDbE0P
42/hFEt2cG7EaqQ8Mto4Cu+SdHzE966YqbX5vuxBVY3wa9+Ykk7xdvU89+Do58dz
q1pxSzrNOlQazYG3Nan11Vjq1ZIGr1grBUGtUhjUKTs9mXsHIKVMU02FahZQ9En5
F/OibptsW1QDBRAv9dSQyYpzl40D1Cz34+nuJXtQ8wb6iC88KJ7FeTMesnKCPWOQ
Fu1CTGYlZvRBu4UmB9v+yNKCIlw3SXmBZuPPY+42vQdOo6dP9qr0Wqh3I95yzS5t
Ohu5GPyxb/3mZZf3ph4LD4Y3mB3O2zPSLpx1SLnmBtT4zkn0VJNZN09xzkiLliky
kD6CtvOYMZN2mQrt3gj20LdoOmNQ5ai8CnF0Bx5a+GCo/MUHvGfxj3ZREw+PqzZo
bEXIXqwtwt+wg8XNK8V7DZwwdzMg7I4+SiuE910U0Ndi1LtTbKTlB1nLzcdLVQ7U
xYdkFPjLbs8YCc/LFrT/NHwAndB/+kFBS6WPerE5MvGTWTGglZCTU2duQhTpIepp
du1R/tZf8yMVuZjUpof3Zs+9+xgMNwgotFMSdXw8qmuq+qVeIbj8g/nchO48iSh8
k+asJOi7jWhEgN204Nt/PmOroLUkS1uGCiMWiOEt7HDCTHNsRfiuZEqbQMlfk9sQ
MPQF3LWVa+eBR8BQcVzJrw/tXZ068ssjjrUY7i8QGX71R3EXQtEI0CEAB9iCZz52
qVtSapjBxSDaGCnZ+qp2cKtxrGFplWy+rxfR6aMLKHt9wFzWlpNuU08aUiIxXcO+
sJrjlFR9lh3tqdEg9+mOGkeBqcssq7xY2N2xSVAc3PF733opYYtibgNu+iXUip99
I0IX7S35jABI4mOe7k1ozJbzO2gW7H91eAO6Yk5HOQRZl0KMmPu+hyIa4VLKxu65
9nXLI8NXeHnpIk+MHS5QDyg/9jUVN+8Ov596V2qfbaZpEH9usy901AKNgSztahj2
7Zyt9sMkJQQH31DRwqK2QvfbI3mY6CAO/vmosUifxr0Vipt6AaFsw1JEh9K6GBLT
BHpD00wymNY3SlUkM5pYzheDD8gI0eg1gcH4XCRqmEisP1GAsKpQ6sbot8Y8Kg5N
g6YiFZbBrxgjAgy2RiTWNJoJEU8wXizoVqlqLYapLuB/FC4pjrK2StEM4zz3kJox
7FQTrn44NFGMcZ8+n80JSEPxrsZQ4DBuKzc1Sc8ufRRP5II+W8395Y1v3iV6leEe
nkTL0A3et/blGfoQBu0V37u83neejKN0TDaaDaKWCq/rsKLCndIpI9fE8dps6fl4
oLhWmHOFXGrFcZpeTjf6dccAxlvB0Gq8klx89YBGHcGQT4L54cuxO4qNSXNQSeBE
mkUp+jtjdHxGhoUtPwkNJX5f6X5I+ea1/RAgueWYXwNLlLE6T1gltaVzZfcOpgwE
8Gzb7QG0Q6K9XDrm3p6GADjWkaMb6gQPip/67X6vPGIAp0jeY8Izb5trtb6fTAGv
Xv/Wx0z2w2DoK/s4QQEFVAHVzb7hS/JekwjhxW2iPcNKyy6CyHDejsFy1FWEpPvu
G58Z48ATJfcX9tsaJNSCsrbc37IlXXwnDng/nZbYe7kLIcNh6SGrEXAc0NmcFSnP
BsaoETOM1PQAXC6nQBpmxd8oCMFuLFtM3Hs5PXaXSbm5RyOfKMxQB5cUAZxNXj0p
x+iiuSUjkcHT+5U5B0+Gt/VGeStknweXgSK/XJIrQ3bkn9dtLqenHU6ptdyF56n4
IQDMwxexmtphWQJ2a8pa/VKO4gx9p1cl4nPZdVVIurvrgdeqg0WGDVaVOI1HEmv8
VRW74TrQVh/LYp8zJrUkZ5Cbwuq59F+AbOw3MdwCjOD+WoYpK+Kj8B+FcOYBoBnU
odB532hWu+e0KZ+T9ubdi0QDHsDvaNKrG/2w1r77H2JeHPIarJR2iXjCAQNn8Lxb
10Qfou4eX65OSXCtlhKtMh3LBZUNL2L+WFtP8D5plbmafrfpHgIS31vVVSIUfmAT
zhd7nnkQ/XlfaDGzyG6ci4Q3ltooBGG0zuPBFEiC8DDv9DtnsTS8NO/TdB3An+0M
fMCUXpuOMYBiE6eCaDHx+3STQxmtwkoUgaCPmXQJNkdTU20rJbdYVNYnd/YX5RoL
ZihoTRX8i0cLKb0q++ZX6vaKh9oiivXTX54BuG4EajQYneb+95UGF6vaJ2izuPa8
7eBjARI5SzsyeX0X49mD1lIeNqgDWdwGZ03j1zcL18PgByOLNRMv3ymW2StYZeeo
obYgJRfkFLQEnHhizOSDyZBz3eBOKRxfpDR2PsUo/KqVQ1WM2mlMmg/PoGWbODFO
7KsySc1Re672NM97i0YmlyqNBtS7XO+Upr0tpS6Tzi9LYzCLJJcrxKs8k7T5AyBZ
FMy+ttGOzEupJdavjv5V0t84o9vp+kc/EZD2DAdxsZU3b43Os/XonlTor8SI8LYN
MiMmi8+Jj4PV6cXYuaCsujTqu9NT3IDswMzvtPHZxF/M1QX2f5uYi+83J1SDrcoo
QwSFt8FnEGle/eMC1LNk4YmTSJOWmxJ2XK+N0DmrDKdboqCesYjHve8EQNsUFtl4
QBzENQYLQboSMS5Kn1S43trTxKzIeSWJoGf6I9qJUdB9LajJcogZMmVWmfPLe1WR
fpmK7a3g7+dFITh0VcA+69ps8xn1r0m4iDoN/qJuaduFyNc6b0kQxfpbmUqg/T93
pl9/i277a4cvj1KBYbOv88eRZvtPGZi/xG4qUlT0cM5C+OVI0NhNAGi5jGCNB9nk
ff4iizrP8nrW4Qd2DtCWUfwC1l74R4GdDIufv2MDE8ipBWK4xO0Viqjxj3Nlg4HO
LQULxsR1YnvD2UTF4Rssfg4XK69E9IenGM4ZR3mwjg5prXmwIppAahLosu5QcTgt
gU+soyRkuuSVqJsFJcr085JBlkot9uExl0jHJfMc9Pzz5jVHjmF+Bstcu7unn0hZ
y121IPx0tRNuXZLUTauVjzBH+ImvBDLybotWPuu8t1UG8lefBSdk3a2if4YsRGvH
h9PysqUrv/mvmhQ0SzSfGP4cieoaCfknPkA0QaPq97qP9r0m82M7arvcpBTazuWI
YKeUi4/5AqvN3qJiaQIPBMF4WzM38X//+9nIsgBZR1rVyxCTbqywwF5TF2iEWwWY
CEUOVKvBaCv8+tigjZ+EFKv/1cqgAmHS+QalCflaI+cMS0IPaIWjWX+l3s0xtd6M
ynt0u91Zcm69P4jU/jqweKcwsiuOxcQ4oPNHzWzP4XYcfgn+M4tYsdrNiyHflclf
Mhq1nZcdkn9+v3hct7WtAWnFe91jmCpZNKmTr4+9phkWwnK57cfQTqMVXkeenQeg
JuliKbNTzYG77hOhLMLViLBX640du9TihVVqgQnbSCYbAkiAX8LNOapzpmd0mYqK
6PZYCc1yE91xLZkt116MWJwqAn9Z81u5rnOoGiI2c+5mbBbGicSHQSgqtrNq1avZ
PC5UDS2XX0RAS3NBSxf8hDOrX7rPwPHkkB4gOhn4ROBA9gilsuMs3S4D5BkeExOG
u4VJgv2DWvl+qW0cT13Q+0kifixSsFbEy5id2e0B9GsTcA5uqQABGjM/edp2f/bB
ZQpYsr1lWvtU8HyEigE2gyXHabr2iaxdWWxpZcuMyGrc4G1wRTKwBxZbK6PNeFWa
L92X/m4ZatvyfEEbL0MjvhpCoUHwnpY6XHmClYYLjFchyzATR4RWT9LFyxP+Hrvc
hh+aquV2H/awb2jny+PXci/eTIy9b/9CNqG5YeEYjQdoSg22i8ge2G9SSstpaqFs
Ov1aXZQG5nCEqku7yRy78zakhyjNBEEiObA4iapxJ6O2FX7ZZ2UGoUCiO6ARJRdg
DD8Fg86m4l9CBTsiQoroOLU/DnMMxFkw7hzfYidqJmBP5zvU0AQ9dHCeYq5paBd7
OWv8jwOvnH4kend5kDnZqOR8ORel8jcskyDmfzoGIJvGg42Tu3wn6AxehfDBkpCM
BRMiNeoEEryTNrw1O3IPDDLv9nqfyquKVYoTsfkI0f+LzuZmilLvHFqs7V3i54b4
zS9erTJ7X3HlPiNk/GEtW16AYcjeV1XlbvJ5jvEBk41GGBA3SLsS5tjqR8UzvlFv
Le0SNt6K8Tcjz2r3tJFyADs/D/aXTQ+W+hYYRpA5yUHwROyBVwOo73MaXB1vxj2+
S16RiAZC7bEHjaWBhg9E1uTdNmlRkoXV6aVOhATEBautBZVHi4l6avA7IyDmsGsu
lhCUdUXDmTksJWWltrPov0aUBZEG+EpTsKEPSfh6vZy81cWVGVynf6ddLGWAvE03
uRfJeJiIofRaCXTb45wG5/TTxDkLAFYmkwL3cTXB5u1MYQcuwTIgiaIBHTeZfheV
Ux8k4IF/HkCAaoV4Jk669/0pyOpttnLLWqtLjeI5ZdbgNzm/LGnjSzWE2n8cK225
q7G1kHQjfydAVQILIqt3Uc5ouWtR1skKraQNVOvtHt0eDX7HJ0bzvVQ8rcBIYtfB
0pcNghp0en3I6Dif5fJuCGEQ2w8Ptwlxaffmx7nJKrwZcg8etwmT+Bs/wG3QJw8a
H9tQZY86y0NqpOBhxuvKqfQePj2FfuwdOY/P+HrLI/CXi+Gc1s28aAa6njT/A6sY
0+T6ZWCj9I7rbl3NeoIys/slqZn/+kx1sR0+eB/iLnb9Fkl6KOH46j+/XL9NY9ox
5TsmUgnb82EywniMtH4UCqWbOu31LA58UX5snx/ztZOSYsapZQp2hQyhWUqz3DzF
FpD8QZl9RzL4XfABBdGWUZYDkm4blKZk60R4JzMlSigXNZ87qamkuc77uMZktN+m
cNYCmi5PCu5/E+jqnYGA18VvUBrdf4subJrx/Wn+VJs9uLwNtdxJUMq18dYTgCOp
fCuHOz6bbJ0D7iyTa4CIyCcd/yqjKYHmwS752i9izWwU1jR44mQfVU/WRZ/SWi6x
OEdkviKJCisS73B4VCzB3TGRBZ9vHJDGUtP9+3zx2HY9WnE8Sjk7wdvvT1MLoGIk
bXsCAk+YpzGDqjb9WuxLgJLe5cBDbevm3EyGayZz+SunzH9cI0PC5GsZshgKrIeY
A6LWXQ+d0txB0rQhvA8o4bEksNQcwRkY7hNPl8QQMu2ninpDIqEqHOxd3sdMc2SM
/QGJJXWcqquK84dpjDZ7DtDVl6PUfANkwtkF8usZb2MTAH6Cjtid3AsgLKLNkovy
c7zcS2m5cwot5IB6I6K8aPGJBqYMGXly9/vdshaeoxJMZ7AGujWGvq5znbN513bJ
9zG7eLOOOEXXXEqPiqLXqmrGim/kIqg5NhTKCcUtl0ShPCTbc1NxfwKgulcebQzU
7ZzlmnOgfG3cS27QwYkavPp230hbV1hlgZtNZCSOQbA59vZCnr1HZy/yRfxHrZ8w
c6UOU23CUGssJOxdyOLAg+k/99EHrU0QRtI6HB4MVwY7CMZydLeYazfg9zk0o/Q7
Bj5C1qO9UaZEdiDoypulky9QW1C5etegb8vcE43gbr9ac6pAAlIxyqdnv7YNXse3
FUyi16VdFFQ13mkiY38N0e/04NQ369P17UpwUUqO8CHQvaSfF9EailqKSTxIsVcV
dng88jP4wCYzPUQu2LaRo5LeJ+oxbvWc31vpkh7PB4HvOIy2i1ncu9ZwVPyutrbX
vPLPGWPNnCiJogdiVHaA5QBBDyr3QnTZJBYMmwuFtUes96c0bKLmV11KYhr67LpF
dD2g0j3S4rZuN0x+LvFpYYjWKDoh0CppoCwAY6955oB4CWhycV63RxcEbRcgdby9
pTbnsUI69VrFbVBCye9E5+RyP64K9VxlR+48m7G1LjnEyk77HBOCM8NSbc/3Ka34
g7YVXjIlMvWrKpM9B3DiMWOttXNTEWYy7M5IWcvYNKEc9Dcm2e7TwElUFFUWrmYY
kkERZgnD8iGqc+RxTjc2j4ss1ltq17jc7BHLTJqLRTiHPd6Fy9fueKPV2E3u4muy
OX3ImqwTODyVPvjL0RSVoLoPBlS5mzTtL2+C8QZcQUgmUHT4SvWvffpaUGVE+Z9K
oVmCzwyxf+sUEvQUAwvqjCj+KcgFYNW/HaSkVd5agTevXMoskPI0SjhLoBlojbtZ
XR7qPkuEYE6UZkBMXtTar94JvTgeclDvVS2ygsLqimjNoMq5aEEWlijv12SpMVER
0qgXctvMLwgf6JYP0kZzXyp6dxHTk+PygC0H4HKS4ogJPvojwYGbGOn+cg1CquUr
idtH0WYKbYhPXTgCU5QNsGVKNv5bjYtJ0K0Gmxcw9FDqDlegYlsv4UWaZR7ys1B3
L1sbKO4vuB5vMrwA/StaA2JCyENfUt5jauFixa+bFujnwUz7Z4DyWKxuPHjOQ8ov
LNbSdaEy+E3a7JbxFH/vN9STvdlQPLTUUU76vk7opIOY+VRdckfABzZATqDzhHrt
ZoA0P+rG3MoAKUMt+MxTqHARVDUCOCEU2gCYNh363NKhFVqLNGyqYyRgCjFqTgIB
oB5KlDTgDXTLpejva8pHzFTCmjoh1Yg3+oOr0YCE1A9PxWj1bVIoeUYIRE9XLHLr
MeCOaOuG4Y9hihBHY7PTIQGaDiIbEIJZ48o587JEffhuRJvv0uC2n8+sMeEEPfiI
crG81GLeyFe0k3QBjWTdGAJ3KXt9doOIhy67uvmnfQ+RSr+9YJaPXdcW9KKnoKEN
FLC6qxsqSyYt794R6IUZUXBJUqoy/vRipR1T5z/biYiR+2KI/x2gZjYdlzgYwOhV
rujMvM1z7+TC/g6fzj1hCP9PU9QlS2aaN3EsO0PYSfhQlqcne8kHcJoYFfplk0AK
MXXQ0TSOz7fdCUHlpSoAKF7W6ANDP82Bi6Nfjqida5pVunVp6f+jwq+3URmjWG3r
9pSpeYJE5qmUBB25k+6VwkM/TsHRVT1hj2SPWFjQS5YrRNAtMpIfWr1EkwIiiv2o
V1fsLmqe6liaauSYR3TEdJxDkJUPkbWhZwVWy0U+nvsR4A+5JOh3pnF8eo6EtqOj
hFcdG9VSzEz0WYohLqNjK8uXPcdthg4AppJuoLo0AKkwk02XVgwaIQKy4g99YdBD
5LHE78dANxTozhG/VuxN3u8XTQ7m8T9l7duItB0jBX2IfScdROS1DbogapyK0wNS
/UmLIrRk9rJy2dQIgMhS4ai369kKwVkljnaHQw7WMEej2Y5LMaQt53S6gzKbI0I3
hytWBrQSJ1EdhmV+KIEsWh+vHUc6fDmqqydyyn0z9vXt2ioxJ4HdSKkoYBJ007og
5e8RTXRN3fVgP624a2KdB9rp6a3xi8TOVzU+ex58zIhDWK/vPotBJ6QNgt0TtAbq
aFEwZaxNqxwGtc7w61eHgJqYQCUAkeOQxkFYQHMkSIyHxu+FJS+ePSRQKM+ruQ2o
d8rIKU2L6IV5vPn3HwklbvsuncORcy+vzueiCQKR7g4MsSMX7CMG3KJxdy1qJSju
rIWY4b+fC5yLjbOZNhhAJ8aT1JSqwLrxVVbj0VwW+tcSHRfadmp/WRy3NbI7y5Je
hOYz2bHJ5eVUWJyLaJXRMCNfZJ2nlGKmIvc2sSrQq7gOrRT2GwUkTAqkz2SEBu5R
lPpfHNALO/5FEMx+rkeI8UHbo7HQGEOYNXsGc8KDcnfnYKQanWAc921u6GUruMmM
6W/05XsyE5/Huo0sJn6cTPn65VIizhqmSQ4UvTE24tiFh6pEdvrZLl/X+ztpusFE
AQ//B1gjDWnN7XvHvuJaBj5X3GK36WSZdvUSFErlGxgpwCYSHPhLPLaTZcupuVOh
cVozvrDXiTs7FDZjhWPoFj1fAM/gQeqNGrgrswkzo1kvshwNfMv36mr/pQiIgyCH
ahV5scs2y4F9IW8L3r8ODjx5XhRAt6RdIw8RvVda+fp5dRSsOSEQKnWmqps2rVQ/
DbQAv6th0IzHoF9YBiCr5kzgKHdYIyDzbiEDvrT0h64uOIYrRn+KBSJsbqE88RPa
QUkLTWHthHUl3UvtwGTng9YsSRcsgW51yIIFpeDtq7Z4ogPskG+MMfzoHPl1cGBC
H/vu/hFBf/FikuGmtQ596ieGxOl6LjVMheI1DZXHhcbch+4knH2+pZdnfoX5ts/o
z/q+XgAyZffg2HairflZ8HHWHNFhYbrfR1Zu0qX0Bx/Y24CkjvutwbU1NbOSz/Xa
p8tq9IuZQhmAtu/q4aePpPXwnGeZ4zAvMaEGmSymMKYpg1OHpa61UNrTjNIBUZ5y
SCecyixoohrOk9Trsl/owxAkb8e7Ht3pGcfiClDF8lAltXobS8W9T0+7GSk1lgIk
/mvNn3VT/828Znwbl1QAJpyqtrZpnoozv5a/xRMWjkheemDXOXrFFeFqjxOIGK/q
rMld9nd1vLVBjnhoyltjp7Hh6Fzw4C7SY8uh541Nu2PQ3Tzh9GhCgmrCe09F+gPf
9QuVR6VMq/q4XfEl/G++UgXcHC5NVhxCGwAPeSbUMl0cRI2dvxJRavi+pICQwq0Q
YUNOFNNr6SHuOeSNBwk0NSQtCaESj31VqdCccNKI1ZtN9jmAP5T0IFYm+Pcggamk
k8fDj3YGu2e1LJx6Op/SPzUCRHHAx9isnBiG42CVC9OMhe8Ldj6sWUlC84fh4iQD
/5LFvNeqmQjkiK4mVI5T3m26IoNWBCBmWWIaY2xmJGU3+Hkx6p6LdyMl9VuALrFM
B1v4Oo38RH0IK2Y+SgC+umaZ7mstBp8VD8idsz1Bsdui2JkIRkI3KWEceVfBYAvj
LhZSyfewetMLEy2K+7FLv3AHBok7l4g87blyEM2cTMBEjMq9uDjiTgBXAEHJitHc
enMCFNywzfIz1y+2KjAqZ/sc8UM5Z2q1xlFX7BWlAafeetlZKgxVavgemmXNdC09
2vyIqqhpHL3aaT6U1olZBfrIQCqVtVLHx5G6AO3n462zfdvISoQFKELzrWK3+JEZ
1esCUMYTbUEW+TOWn8XURWI0DlHZX7fgHQH8zMQ9QHVIWReHnj1Ddm1RqBkc2KRf
rWnhXnP2pxS+XOlf2z/qAW8RIVZJBPK1C7GodP3pYsOQWiL5JkE/nMp2X/p077gV
rhzkDFXLyZPQqMgRq5roMjG8kSiCThl1IIttoKEfWSJw9aqyFj0t9Ff2yjzskkSi
ZIli42oD+Y2mvxzLf97nMgUwrW2u43QltRzIQXHJq2rikNqNBAgDL+Tk690BZvpJ
piaWYoHaUGmA4gbmbGjP0l7OiDuHvIKl7/gnH3hUX0x0EAuichNJdem94P+HlFxD
hu/O2xkiYelD2NDNT5sMN69NDPZsk2uc5gBLrKVL9UjbL6sp4CvSHBQikbCYE8gG
dIDq8BH67JlhtrY3u/FERdxYgPSrSzeNKU/I/tOWMHFbI9oak9fkJC5q0jZDmdtW
B5tOkJ/OcWyP15n1xMsqp5Qe9GSBXUHexyXx8txtX2oR0el57qFRbKR2RLwnhvHB
k8BDSOrocwNjnuLsX/kQanPtN8H1s2RNZkSLBTsDte2T3JJattK+GlT4iC6XxxIB
1VzTrt7DStDEKct3aP2MOIoQkf31yjcyOEWe9BVV7asecLgWVY4hnuC+bVdvwf5V
+4BwX6x2z3bVFVAMp2SIGzqGVYTh7gG3vJE73poKAuzMGVRQWR+8pfzr3jirrj73
tdO3NrrmDTc+HofwpAzPE0/zM9qSKwizaonSDegOykUcxwvXRS9+PZwKo/ndEL3Z
uLnkIY/7VxYc1u8v0jGm6ObCQ7+KuPW+55k2PgrQ2uOIyKjZspPsdTi9/NyAWtsj
J64lnymHaGU3cEO9uEajDQMM8szwHBwHRp81NJrom2KutGbuaGelnthA0NxjyDue
56ily8877kha28sbQVZl07QNkBU9MeNWesr3KU3tG4abuyoecjYVtnPJ12qxoPZz
SuyW9ueSBkSg1DlmtGcVY52YC1lpMAVgClD+E+0rpI4H/Yq4jp/eclTnGVSVsrOn
wxyof8sCnd7UvknovWbkXGhfTIJ+gcGan4vFh8jDYIi/zsucJ7NgnM3h20K0/vv+
zNZbmik91zprHHljHjy5kq/8pq5iBDWgss/TpVarmbvG0xud+NiruyrBw2O4F40W
sK/JNX8unrJC47EXI5Suqe3wDrwghzKA9Ual/Cv9+5Ty0wS4oWn98FmYSbobXODS
NJSpSoz9B88mVAUkg2pJqkeAPtxTGEk3t+Q9+0unNn/5op+aK/80PzQyUaTQYW4v
g5G/qwhnT3IE+ZWfYt08IRT2J+H6oIpmHsKoSFBXhlUqQb7XWH+AhTNh/jk0E3Mt
dT/T9v+nP3WKurB73hTuf2d7FhldjBo+YtIMhUENLS7ZqLhe5Vl4oqO/Uv/zcpLg
E8SQbP2smfoJBpo1gcqjDhymzrjyJ0VaxyMNekb6rWO5XayFh/2JYwQVqZ07f/Hf
hJ7gKiazjHf0qAfHGNUQ3zFhhIu3QXuc+/b8FPd8aVoxExZmSrQ0DRHM48X5cFsT
O0FnXjXYehogcA7RzpuNUulByC08OckplQJFQT98fpS/I8zn4DH4vzLqfzviNkla
8i1DN1f6O3ikRwYcygn6u+qhLqoXUR0PIZ4TYbK3S8vJc3hzMRAQ9KiXA5TtpbmA
xIuzoIq2wjgyejJSaLJtq+uTUQo3XrMzmgd3a877NKsNXjQsy7Xewif4vL+Fgx9N
HB+c5uRtq1TOFwid/J3wvE/sfesba0sOS+/GG2psWKNXJ747KoNFzy6zua3PE0gE
/aJtWlVBUQnZ/a36Bhyh+S16b/8faWoIsa4u9s8pnT2P2VMEipNfY4sejzXzSRD0
IW41YGU6oQs/pVjXvTLGddV+2WIY8aEQ9pfCLfscad20VCEIH6tywJ0K44tfLjSr
nc4SkxDB1lBx0r4GNOvmRjuRHFgwvuOv4AbJPkggYsXmfo3HM2wK6DeyINo4P8JY
uWWFa6puVt/puerjYpilleCm78kpq1osfLT3jf6+AwUxjDvoEzN8Oyt8Pz3+zTKc
lNhwnYKdUBb5tD9jLO4iPtXdImMExMatEyexbzvtWn9MMvBWmHuR5YIMGde8heYX
L8ZAlEVvSKD1opVeGl7+5fXRylII0l5JpggomKY+56S9TYbvxb06FciOIx54Wz0j
2YqJ1zb39BBmxFtEDgkZqQ53YKvazNzUwSm71SR1VVe0Sbt5/qbVa3YOYrYLoL9V
erR/mjXlamHqiN/ZHMYSpiwFIISRZi4Xg5bZPLteEYOIW2IJ5cxXc1GT3E0CyhA/
33LddczMrjkxduysGjmLy90TzUQHz+24e5lsdcR1kSz83jyeasAvAWsZ0F6uNCKr
tvdYDrzRsrV84v6s1g4xobquLQtL64njUjXK0SejEtJB8Zsna6FfZ5lXD6se897w
ZxpKw4k7N/Tolgf1rizySqNtKIrKlrQ0+yrNL805ihGha7gDeNINfvExxH3NELaR
6KZOcoqpV907DEoUjbwlBJSiAV5sQ2EGFrSuG2JuzqVUxIg2yxjpaQlfVkhW0l7l
8NK3r2yjf6WsSs+Ql7UkuKQu35fXnUM3eRogNQJbrWyVQ5PAAq4rRjmz3CXVqap2
xhL5TVremh1Qs8lI8YGmtUX37FFNP/99U+KSLB5WkiXfO+nDv2WDVUu13LEXf5sx
Bthi4bvAUEfgHBTarvn+/j1+Iw1Y1ZM54eNBp7PRj+Xltp4uzxynWh0s4xr2b1iF
bv27z9XWV5W4C4FWB976z2IxttRtrdLExQiugYuzJxXl5s+4QgAasdsk+zFBlbzt
cgUTUPbRUmVUIml3GAe+nF7dA4PHPJAFmph0a2NN+rv/aRU8AsDE/TvXpuIu/gZP
+sxkP84IAVM+BVy+I9FAeNFpyzM8+C9j68a7sAxROQ5DLI/dM7eWxWzXZ2CVfVcF
zVO2fLSgXjIc2vUMEofcuNGUu7iDTCLUrjk9gYc1G7eh5m7vcld8OORspue/tLxn
NLvyVhA0UQgwi2tJEUYGuOc0R+R7CDwHRYRsBp1h6AJ/tKjcXn+rBFwMFHEcSMpq
lHfFxd7IbdRznKNxvcCFN5X0Dme1iF1az3Mp1moE07gJA0Yc9E1QIpXYwInMBT0I
gvZhPizreOQ9s3UhocA5UCV7TD0AzA5cK8nI2RvqnZVedHLvwG/MQ1SrEmRpHx7x
LbqBrGOvPi4aEUav5RAXijNusd7Eye4dQLKkeNoLyoS8d2oDoZZ6pa0FZtMapmFx
kwZiR7Drz8r58wfFRUgNngz/0mAdzB2Npg3mK3N29njVOTaA5AnGgepmM0LU1f+L
UgnsQdE4Kw9yU/b4GIgvyqewUzQBmp/lnreZ9C9v60FURbe96ODMCqL40aYrB+vh
d43mfPQHplPj4wRPblmQ/i++0l6luPhMrDWs60QfYSBTycHL/3wgxVxsq9ohp/ej
Rtze7MFs8M/2/JT96qlxqaW8tUTZVluI9fqlL40szYaY6HjbSlO2PO72OajfJ3sS
30AbvXcAJSp0USPIr0hEUiikoNK/NNitM3eHCcSJ5YhjAypvfPh6aa+faUlthWnF
HGz6FeLCi5baeX0RYQ9WdFFZowc/gMMZ7aMokMr7TtJy6BbgKsCV6IU0qrFH5oMI
u+Rn/DQiqd4NPzmG1QIERnjso5Kac9J2tf/i84pXRU09cS+wm+CjfH6XiGOR1e7m
azzSl4EJ5PQ6pk4cYoQ8XugeyR4EJORqnEOdli26ygnRhVUYlM3FdrsSJbWbpBpO
2pOLlQNNHfeBUnMLIcdx4RkEhIL7DLhxLLLExLaNbfXKNPaNefiKBIwU6TW1hZoh
KheOKxofw6ASJegYUOK4PJLfKsmM8JK2GzXJpuSAMU3/bfRID/5Ow8pKITdEhmCt
Peivdaw9Vm41+N2KSlLH942yxYYkGxqhbssuMdBcicnbVKgbMM6rCxOSHsYH6Ved
bgDMspXHhC6yWlr7P7sy0Tyzl9CTttHKfkR7nU8UhOGQFEbuVoZSpFstr7Gf/DK4
/qpH0l1hZHZRaVqNSuF91A59188tUIxNzk6ieDIrJ9BAl9B42ddYTFKstREjwa6U
5eH3CIxHzF2U2on8w63bIgyxPq+t76kYCfEzCbE0/TP7yW3+w4oF4ivYkljdVa1v
q4Joq8OKIVT+SKQzcUTvFBg4LBNkoixdUm3miHCnAe1LdlboH0BgNuLZo4L1WiNA
CpOMuv1felg2zMoc+AiMrYM9QwQTQ3OdmWXiH5eVPNx1KmdzhYoXnHpflcddN7Lo
1I8ApccpUJ7geIsritmHPQ7cvGZKKpOUNTGxcScr9hoTVgPvHuHnYwwViTfeWWno
hJa4hv5TIHgYDzZctVIbp8W1+33scC5GwvY+cGoswgWab0No6Jg+y7XQ5j1Wh2YA
sL5AAludIu4aaFWFWu6XfPgwS5J2c6lNPS7HHEp8x2eTb47rapkj62HSQVlDnjg+
O8ZxC0Zcre94qdTtQXdwZB2CsatccGHiOHtZh8EcjhB356FMQQDhDfZhOq15AbCk
UtbFyd9b3DOVUPcsZ7sCa2h98YZmS7LE37nV0/tAgNPLwoWNNNHc/eqv97raFJRq
7apvFVxx0DhS2QIqFqNuzAJPtfH4o/3wHjUjHIofdz2E5FkP9DC95MYeY6HrxQDb
olsOxoQyD7EdFaHymxQv092VUL2J87vjQ0IgfngAF1c25uVWIGykpjmo54rBmBqC
Fsz+EXu2Eib/O92kGFsBmsdKoCXNDCJuZNgBdakzUFBD9w5RNc9Dq6AqFhBG6uTg
+M6GcdMeIiAz0V+0hesneLDrsO6ENfyPgoCDm2P7Xolrt7R4Ubytkqu6LdxADcMW
3JB34r6eaOEBJd0sJtWOCucjloB3eD8nMXJKOe60wDTIME+Al7kdtz0aHsjoEVlo
daILJ3CLEjizOP8S3l8V1ebq3LpsKNP/ITaMHx67R7EdrmTX8ZFi0zm4n880W8ug
XAlTTr9YLooS7JMJevXLE0rfp70DI1laH/ltRR2wshhuHDgewlThxNMLTC81veNC
rn+ojzZKDNmImWFV5Sm87coJCGjpx/2JVMaT9mEhflIFi7tvv7ZpJsTti3lZclze
hAilvpECzjCWz+Ekhr36/uKERzbWeA7JXs2wa/2UJe1+3G1nQbV7LnMNSjXKSXk7
VTgUWh1TPE0IoURJhAwf2Yp7yegjvznor0BQpQmaz/6gpbNNpHLBxUbMHUiSros2
feQDonhbb5CRAoaeSrN0p1lvJUXdBBOn/9KGBE1YXDOWfcGwbtZLKFtLLXzuqteA
JA3r5ZehRL2gbnPWPM5Pauv+6nb/OAk6yIa1gPGcFt7FB77ExfC9Uv2Tf6EaJGh4
9Q2RxXowjjwoH8UuBPwzhHt/dSBegrm+8ZRmogpjJTkt2DT0Cs66KBs0EpGuR1SQ
LAQAELGGVlqT10+s+f9UNs7p4H1yqEDToCBYnXlUDSF+uHiE6HXcTjM+tfi/b/Qq
sw1z2WkVGmD1jju3vJTEzKRsQV3JbLD/gW90Qc3YHnEicowu5WXP2RZuTuRQ7NHU
9cDb449gWklwZZ7c/CMXLkCVtkmWZtvP5j/TR2HezpHQ7mYj8Dg/Yyxlqe086rMQ
iQCgeXJdlHLuAxw7SVymWcDmwYtbhH/6jSsK15EduDS3F4LxxuWfwbZnux4w899d
yHTLYaxOVXo7LxHR4nGYTgqHrLc69SxMgEjT5SkBJNi3mEa5y7BOzD8fG7NpT3mw
ixGXzN4zDes4zCyGGfF2jlK16p/A9HTAGBh4d7kKQOvXWd5PygzC3H5RzSEzon78
tGarSKVdjB6LbVYreu0UPs9xrZgPHfsaTG+VZ8El3zNnUA59alxwnUhL+QpleVZC
khR8YFXhI6lSYccTRAdPLFXet9qFDzN571BWkL3E+He8UpWcVxEZ3JWYVWjkp3hK
I+gL2oicAeTsAWWzEUNwNYuV+KNqj6Nyxm7TL9IcdTFf5c8CssjAJ2N+bYFT/qaT
krRFgiWsmCMkivOjduv76gtnj7/AZmwHfyp87sT0WHZ6csZQVeGvGHH+PLTZ9i2c
B3q7eL8TDabkt+fGbTlHl2dbDagHwxlbNUaurFj81WLNJ6TB5zLwRjHBg0Us1kJf
mLuGRvgdp7Z6ujXQEL2vnJMGBf/swgw1fw/KZRrC3pAfqYUzw/aoIJriHOutNwIy
AOXHEBSNaSJQvLdCGMAaPSUmpP7fS6DzqoSr8J74f2j5VXU7zdJj+NDLP1lwEVWJ
Xw3KFIX7j8B2Rlm56NzPxqdJJaJKKao0WlEpVbpWRlOgdGP8FLfGOfhVNh2zc5uL
zI3DTMkYrO+rD2eUAkHmUw9Do5e5M/sr7xf6Y3Ofx/Ay1ppDbPJf+hvXcsF2T5IC
Q+NsbE6mC4uJrHI/MWYtSSwjv/tNttzA9I/mLsFn+mLyWm/IXnnBJJiqrHbJWtNX
d3yxKTP/SHQPsShXmDaYeMlYJM6FBTrQAFwDeTsGPIYVBwf+oxc8VehxRUmg/dQn
jEvDG1qXUQwVqIgRC9jD68WLWC6j31iBaFmwqDddoD6vg7WF9US6lekhGu6krFno
2x5n1MbeRLQvX8/prsDVOOP98psl4hbPhBSxQBgC0GgqSnOYFz128tayUlNbFB4/
liI1ListVzo2N+WHr//gWfTILUP7NeiMLWHODqSQtAFdfDO3QLuvL15wGKZTzS6h
pA9DK8ccGp0Dn0lTkvxo4OLAFw9kSyP7xflBKafMwLAECvi3LCFGa+uUcmuqUBAy
EUAOtz46HcstTSg6k34KYgASB9x1vt4PEuyap1d1IIgWyhOck0wYzgxIJ7lMAjYM
ywiu4pHrckouACF46VRgqpO3kYAmY1gPYUEUtEWXrpuo9nsvxpv9bbeywBgY2f56
imytkwBLl4MVRgrgYOuA0Zpzxpi+SNvdVq+PxGBrIoT0Jdyn64bYWKA1LETZPWkG
W9pJ+vH1cJpeKDkZjRNHy8RGT52g16VVrD+yOZEDUcLvCYPatD4SfduRnmNDg7Kf
lfdBaOVPloRt1C5Jor9zqGzylIB47gD48v6eqK/FN2eL8sIMFZC8YsLaTk78G4pQ
gASKFD+bahHBy0OHi3fqV7DbwIrG2qiRDJX+Rmd1FoRolyb3CUzfm6yR0Stwc1/F
XVE74frdmCyuuDqpIKjmvciOUG2bzGorOpUQUZv3EOeaN4vlTDA0oLZZptvqaKSZ
OGlFUr4cocokbki/ONVne2pQrQQx0pxKzCwpNug2yOeAx511etfdQ3Hg8+j/UyEp
67uUMZhfdGZQtKb5Z/60NFFLoWE9+jL0O1ar3S61gqE3IdryMwXyifrQQX5h53H6
05E98I2ew6j4LLAgCdXiNvW08z3JOCIEnryM5cXYtAKTifGkYUm6pNFGMrx7xo+R
ie9RBHo1lsPrvOEGHpky1bDaCwfyxBt9KbojLHGfZjJbvBwiINz1h+6r1DZBzFSp
ejCN3Rjcrw86Hk5owOm3cXz+jdQU2MTrFZOjyqT3SR0zOCGBsGw6xGEOqxR63lte
+udk9PLE9hftkss4UnuH6VFRaCtt3+FXeQ7LXXYTiHy6f31c9chX6m0i8J0tOrW+
maB6VsRsZhvbILdM4n2mw8X1IufAkdOPmO/qLHEr9JEZN9ov4my8CeB337pMVk8E
+R7lllQnxru3UGwtG5PXMwL/jiFlzP438ohGbWRy6cXNMxeroiNSkVWSdKgwFApj
/cTY4cBI1luIFsFOpeBEJ2K+NPgkIdN1LbSkF0IsBvcli3LkCrHDzci6HNfyJBb2
ejlihEQoToaaInEMUABXqxqpCQFxilWqMo65bvRdoIjDP2KiCjZ1AWpthRGpiC9d
VJ5xEHUpAVU+SD60QWaB1JLprGMEctdgLxLsIPViF1DJ4NxEPJQuCj1HJIjhhalO
gZs8VjKZMz0/UB0605ThvLOanvIqEhHOID1267mNNP7dLQP3JMJRW2On7W5T7AHs
q8VvLBnO2wi9M0qFE26TcMS8rKCXYP/EJPHKaztBOFSuDafyya4boRKVm+oC4AIv
ecShjQ7yMuvHg3O/7YCH5gK2mLfXa7UH4msu9BKE3w6dn48/OHzcY0K70GV3OFok
WR8ufIouN59Wbo6T7tSIIyrNyn0f+7AFnbFZiuSg3QhYVK+co9KhknSbvWs8rW4X
pjZtIuucSTJ78lFNN+eHwx4RV+5ENfy7Q1zS7OD+IOsyiCw0zHPBdgq0qbfRqaJG
sqOgslKOFW05cjAvSXyT4K6R7J0Z2Vj9OZq+PUIYyzOOBkKayLMq2Su3flQTK1pO
i9oIqswjzavsNlUNWIVuAg8qo3FpONwxvlN8quec0bDRS7rNnsBEmMm+cBdHJWSd
8TKTw9eVoB+PHWqNGVQ+SWBaopsMjxUgHaWX3Z/CmDFTGnQfOcdLGBPg6C8j2rMc
j3WMmOlN9WNL7b816kOE44o8e5/QziWrs8YZ5DPcc2etUrwpEw4ckPuMfClIj+8R
r+ipntm7bcMuK5h+cUBHx8SOcQtRmFD4ehIVRsDlMr0UtdE8U2K/K+Do2XMn+UzE
8d2tcIKHDkkUGpI5olRcwof6/QR9qk3nduC8UfI/9X9Mweyc24B0ZpDKSXBfCxN1
ro/huTheSG2b7QfAqGgOx2wwlfX/K1mJ8zBavL1Qys6Sn3cCgfWEbd80x9QUidgJ
l1sm0xyWKiEPOP5uLwk9DoOLIXtwM90Bb/CkyCZTqcYmvc+Fco5Y5EdRNXD2CoXa
0y/tBYpJu02HOMENBJ4TP5K8xvQR6Xt+EJJXR7dKd5orXVX3gxTgqGd0J5OgHgGP
p+JM666PN9WjtpqvyOv9MYCrbPOxW0QGraxnm80uVdblx73xp91XPp3ftR4zNWkn
WLqwJ+5+heTEW+HCg8tCi1pStS4rjMZHGMSexDwHmTmXchQMz5GhW8s9tfij9tCH
0Spw5n8sy/uXGBEVvMXq72uwC8SgKjgIlVPSfY0rra6XL9X6pvPyrI579AVDBbVa
HH0Vc62MyFntPm0BY559aX3Oocjwgxflbi1mY+zQrop5oA65zJ0tipRrQArmFIPQ
Fv17SE4MTACrVXtW6ybHUaGryqZ99xypSp7wZKRhD97LNmjhnNGZnSwfBYIAPF5A
3c/V4S5jUxaGakqHpH6LsDl5kQf7GkQEyO3XWm8mjg2f+2aHPYLXm6946sQaDs7J
aQuLgKbPAmey/JLMKV22ZyxaWMeQgkWsrb9Naw9mrUgUrL/TE2sgBEjnv1V7UkQr
IxdB184rfPW8tYA244R9lM2btheHlvkOqtfsrownAvoOvsRV4ArAlFHg2Qk74ZoM
W4y+NYC97CSYjLNH42ye83mCU9sIgVb0yyEOY6ak1A3xT9XFRcI8Ed7zJ4/3jrvz
IrHMdGoPeI3HW1e5FWWnFuihkkdeAsHucxsiD0xArJ/WDhDgxhVzcsq13X9mIEh/
l+HUWdnV16H6Lj9aldLnngve4etiODC9IzUVpYUgBZYDdL8bgioVjBLF05FBoG7y
AbIRnL2m85HsGh+K/2JSoH+TJEukNS+tUi9uEfooFBLDfKU9G5sa9l1C8aMWb31T
ViHSkYk5VQr1gt3t/Z7bAGRXhgDUxanO4lZ3AHn1f9NaqkRbPE4inE5wvqvLyOeW
Z1b6TfDAHp2dzQBqj64t1sUrMmhwMJjrdhAv6sPHN/cMHwezlPdD8nkGmVAdSLuj
BLh1uPDRPHmQpDwylEzt3YnrVmosF3Z9pHQYimq288/lIzAd94w4N90E8Q78W+AH
JLmcdkXfHjOPkUrRQG4B7rczl8IPXRyKcufe0SnphVZfDEe96uBvxJdm3GYClIsd
c2Bdx5KeUOT4QdeSL2asBc/GSluKhmAeeBX5XnEYwrGQUDF4EceGcVcDAaONLJyc
OOL0DEzd7lh35KQl+XTty1CKdMrGStYnTFKn3DG88beJCL6UXgfk4BcsvPCRj86C
MWgjTUJAC38WTtndJGN09TUBw38WTNtapeWwQ0gT8WjpJ5WVWDs4C2C/42DNPW8/
I9n8SYfFtfKHE18pfWTGaWLBtij6Stwm5cj1HOYHa5LWL4JPFkHunCVzocTbukCj
tR7XK78Zkj5Axjh9rTnW3EGT/uTrl5aMK/QUUf8YyEOfPyymTWtKK0THyXlS4y7I
oP1TyEbYqkHRcNxuP43SNgyHPV5Y9dDOltAKu/LU7fVKedA31FTWBz5TvvvFMgrJ
WI8xiKZf4+8qKfnn3ZhFtdPqjxFmd5E/Yr3qR7XWSKsjGPnaBR3bNEX2A437c3XJ
zZ8bFZKgb4wQBJw86lFIzNrM9UT6YcxT1zMRWhhYTQUFtGRPDFejTo8+n1YMMW05
UCfRsU8wU8EIJP7xuowCD4YSnnfhwZNCw+l/QXdJVPQm54my9YFTcgaba509aSdd
0THvWsCfiE+0kWX6nPDITt87ILOzplJ45A3PTzjfNMz3gHJkuGuNYJzPIo7nkS+6
NptTkOMCNJF6g5lAN/lPp326DD6OmNtPqf9TyUOmbTUVQOFBLufA0IiNP0DjHa86
tBXZd3Hf91ROngShweEIuLsGd2HOsqMeYDL4V+OtiWjR4UeY/vpA8ycUKzrMbH09
xzadqqQB5ldasZ/LuiE3j5p6vQLJdYCAMP4QJIXgRefOlupXgR0fo2CplXrip9oa
onGBa7Qlydg8vsMTbh1EWbysBXhysaJkzcPadxmZ9wqlgaSkxn1Ws+2kpY8fpCze
juMNtch7xoWcLLZb0CppE/x71aKvDNYvW4uUnMKjkaUA/Uu2v6qP7pP4Wr5O23tE
Y4sM/Ai7rFdwWkW7pZVaIKbd8ZWFE5t/HFcrkUyUZHzTqm5H+Tovd3ypa1ThrLtm
nj0Q5/WRIw2Ha/VqvN6O2oVkUKXPlOtiVCBGyVSTmVf9FRTFcMLiMfusBCmr5GTG
iOUcR2FQ6nwJ4gYy0OtZ6T3mHoqWQ11xscRf872KGw3G3+H5awvkCTuhs/bNutdS
9AtATmRMr0OUXM9oMg9K+DN6RkVYfsPfmpX1zU/zcVWBCFXp2vuTwbgplRVo1p+/
pKSsvf5R6F8XH4pFsUmXGQpxf2OVwxOTeIOZm0H9zTKOjSHFxxPyM/u8AVGNefwL
shWeIR+q7ytpHTD6MxvedmF4OSPaB3jnLq1h8SaI3I9ZPMF3m+TPtqJehBv+G5eS
Nbc6N0Tec1QNX4jLWZE3csNPkGaUjP2xMTA7oUh5AE4gIcNYPhBT3GYlVjQt7WFZ
1RkswW0AV9x0Itum+G+bhlCGnx2fk2YrDRaH7MeOttSwoDiWACR9hWl1RJ2mrm9q
Ivn+N6zus3Ikq1Euq63PLQOESyxP/KeUDi/ap++3i8tICzns0ZegXfVjhZwdE8vx
lSHAA58ocXKBFlljmCbTtkE5MK3tAHoby709LIRNVV6D6+/fVEEShd0St6v6+o+0
5QEw80GmbuW0E4z7Xu6Qp4DrodfzGJZ8tjvp0G+FeBDY1Z94LtAVMAtHgqiZODpF
1Pl/t7y9CJqJE9qVnFAdZMC23JFmc+UoMPCh5AL5r4G4367QSEFx9eho/zarVVQv
ZM+1PRYC41FyoeqcJ6QARgcKT6sFMZMJ1VN1ooWrzw0u5s+L8CXXevHcU02h7AA6
z/HlQjfjNwZsrO/yIoSckgaC/Nn3PfwgyfOnsFHBCK3F1RnERQFN/mOJuuZk8DR/
yxLephS7+sspBIJkHAngTiuAjPhn0eUXRuebNjxcgmS7cq0VNyS0CSWlF7ae1bc7
lo7GdxwUDL24F8Fz95Sho7exFlP1bb9+SfrVgn5YBxyAr77ddeUX4zy2h27LpZKV
MurOJx5BV9ENKIXdyDnxDrqrUE07lSjeEouC836MqmSIBebCzNLNV1EPNjvqH+B3
EZ9Ek6PQR1jSvBSgyp7iAZyDVveZyFv+3cumebsEVKc9VZoWgAB7tY7ihaTiV28N
KGDR5Orrq83h5Dh6De0pNiWcCkWZz4h4Jxltv5JnPqvtSEHB+AO4tMk3J6EKY7xy
q1m4PgZrpyNJG1wciT5RaO4GzULZt63eeJGbgYAdbcnr+Nwjhj0dbHS4EDLak1a9
6XNbVXw1y7q9Ok/BEJJUuTzu4XRdPlgczjJlspFVC90ehhj/xdEjsRPXYAPdmqrG
QTEE21eWbaXdTChblzE5z98Os1UEMXwN+AnQngWQr6P9VtolGIsUEjIZtnbVWy/0
uMov8oz2+fSpkizjN38nIGT+koH0vltgJdfjHwxd1eXvBWvxNF/H/PP442M/WNlQ
0wTpCd7RF4nI+7nJ8w/gt9jDEwT6biYc0oS1hM6Cdz+gXepLC3WszRiHlr6ph8Yv
sNFRJYBLeKIIQk8DkP7xP5cyiyoPf7DkVJP94uLIVzDItkGhWWaD4kaLS9qRMXYH
wjSOJvoz3sxzOV1WL6BAmu+P13Qsv7m0O7CnCK53E9dUtQH0zD1DNiQx8g4ei2JA
HafYNvAYIeo6oQPyMUEd9WN+5hGpCpfNRSYKXjWYOf4FwX2EKP6IInwoyFTVVvWP
GgrRSaPfxb3ZSyOnp0/Ohi05OsAPZx3GUDV1edOhWHVK8rdYfrRIyEIYTrfbrdcc
QmtIN5Ax8e9ZiOvjV889iy03/aKfIB6dlISqPzu3SyQ2FAvKo9Nf+oDnf1quCZfF
rzqhbtuKlJ6nvju4tnBYxiYwsV8Vzq9Ew7gU4XHfszScbwaPpWosgl4EciXrQNN3
RWJNl1MxN5q3c8OjY/4YF8gZqa0cIOMn9euWQVSOgOXJcftreCUD6vD7WzXs8FcL
P2jrGLAwuyflqfg0fUIPEux+uyGAe0Hka1tyRjPsnSFoNUEXndnK6tKtySMGjy9g
B/ps1NCvn52faPUaodtI+JQqGz7M1VsJUnElQzmDHtYlIRyXX2RgzZ6oEdIoPZlg
n9XofVv/WAd0MpyCy7VclDxRZYYyuUkDOLAT7zqzibvVjqooubYtLBiUMm36St5e
RyMw17vH4UcOZ4lp+i3Eu6jYPw4pOEYPym9fLWovZqcHEX0Vpcapzs9xevEGezWK
iQmSTkWbsLuUIy3a/3zsQuyeM9ccjXO3WKAW92/ZbDoYgqezzuS8Ax4DeyRNJfHI
8LA7vypbhAx6sN2wCePpMtOV8QcDgmtGrS28+ZbZr7vGyomBFYXx8FSyxyZKn9rC
xyaAtLTVCuO4f348dfBpXC9iO50BMOZItYMq6n56aVfHpMlnnaIPRmkaQD5o1SMv
Z5C1aXICZuYHxj2pT1uM5b9pkr+byWcV+6PKS2omc/uIbcceR84UMW1kGhTap/dk
KIVicAm3ePli80KZ5vJPfjIx4maPqYfaRvpH5I+Wic92lbRHWAtiCalfGcyKf+c1
072hl/VjFdF6snEgr+Xe/AQqtL8bjLdZ6DjaA4vCOBxLb5peV+w/Gfw/wptZxmKL
0pZHMuKhw0tJ7QyBKN3dQUrFm40dKOZEAYBHk6zA+KEZUJVsao7mHWcgZSoQqxU1
fwWGrdhksXGfZnsJ19vDcl4pfWtZfGIAiNOVAHMeEVLqLlRW+x+8RkHfVQUGb9IM
OUom6gLmE5DIFN3yLM2NEgdCN5iJ081hfiqTwItywGJ3qXf2ChNb6eYl2i3R8AtC
RhQvcXMI7gdaJziOCf6GiVXdj4ahBMJjfB7FXKAXJb1w3vEshM9Rjcu1dgfOSPPU
Xt5Vxvh6tSU2YaI/2mz+vP8EvVwlZrEUd7MfyPrzQbBBMGqO4Q2zK0N0QCgCgzFq
tMjSNPmTkQYC4wyyE1EXlpNyTJjl7pT3IY39piufgdLjyciYV8sl+BySOCkxCJ3O
2VL8SsL1vQGwPGwP6HPFNtlA1Gu8lWawK0aMnbTjdHOnak1rhdVKzg0C5E1OJHwv
Iz8sGRFaFVdp35I5/QXAk8Ps+QlMARz3XseCZS2w7WSo4c6xhQVLWn16qn9zeFf2
vDrmMmVpzGz6SRiZu2vb+V267l/ik1FRH5H+RsLcFBau4oJuTbMYT0ytx2VABsur
KPY51L9zKVH0jp8Vyfbdd4XpLJSKUOHKFLpWJ4icBUT13XOVoghE86sPhwouISev
BQQG9iojNcSajLmyw3/KeT9P3VThveS6NTsapTvfuVF8Pti6F1iOd8KvjeYvlps0
2zVzXha2uDJmg8bXE98tqgn8SjlOKhi7e5HkLXOGel4W48CoBx1hNSlehxUxdqnG
GBfLa9AHlaCrs65i8Z2bN05q2Y7LjDYE3Wq9artZM6OWcbE515FpCRYSyRB5+1UN
abQP+yRXAxP/Ivv1gs48eclfQIRlChM6Xzb482prOVPmKG2chZiurW7TN7yhbPf2
dFkNg1aXRUPIM0B2mj4Dv3fIt5KMYhxukyIuLQdnE8rv4+jup1DM72iB7LHCl+vT
0P9qsmL6T8P1MUZUwr5DxLKueip07cJmumfaLkYbLJMnOKTotFewYLWUzRCYr0Gz
H5V58H54+dWN/heR0zc175IFch0U4gc9mkQC4m4hOaDaBBvQGk6c6ljvtbS4FCut
2b4wtEmbYvHr6cxexi4JLz0M3MhFG/0gQlhVdMQz7LVRt2fQShrnUH+FgAS4Kdmw
ecJAjyjRmV4JK0Js8RssUnQT18ci5iTD0rS2xTKvrLsZDGEoZvnTBRYC28LE3gbi
B/MPDe3lUIuDG5bE2C9vJr/uMVs15JIDVRz9dVIUGqUEKWMe9DKETC9gx5/0KWbb
oQokA8LR/sgMmwaOQ+3UTmO4O2Wblq9RNZKczb8+bT/lJkgF6Cyr/cLFHAI5SZP1
elyhmQmL2JzW5Ksob4SMNP/TCa9JL4UbXBUaDpmuSn3EVXCF3jhDoFluxsSHip+7
t0KZjt9lb4MFDo7s9aAxNlH5FGTGDEWECYgd2U73u4ZZVis7tCNV/1DiYjxurbCA
RCDFYt4lvQUHCXycFLl9NmVsiK67jVFP/G8Gsf/ZzfJzFzEec91wGEx6owQd4lMO
wbVYSG3wy6fGoseQQixWwJ3CDVu7sUf2XlfS4cudYUGxy8lHDgmmHFK/txFiayr9
uhauviv9mYLm84O4o8+tb0c6OJq6mTRG9IOpzKUVdR1lHCYjOSKO5Lg0QNljvg2n
gINh6HI1XqDW7mWoyNuDn0vVKF4+gWSlaDEGT9jRUdJnNJUZ4cVmZdWDXSixpB2M
CkurSA0V4lrqZrdlFQn98u5RuD+gqVxVhRCLtzBeQLd3VgxSfzf+ZtSZd3/Sbq3n
vdHFUBihouaux/yJldgKRMlKqE0zIkjH2qsDvfDBvFWcMfQbQQ1dSMNoPfIXzWby
2BX/QordEgR3qgpmKTQs1BWGueJ39RlHhx2YPLSf0olc+7Im3FI0fTGYEk2ImFsS
9cwRXTpk4rjiLwFTvMSM+lXy3/ISEljCLrYbfxe01PfWRbawgBS2uUSyj0tOvTFU
lBXK0Gdq8FjnTSI+E0tjVE4NQA7moXy95PqLVHJbxZJFdEGY2n2gr9+/ZAgBs7pO
OVT0rtPFle0FZVw6MBnHHOnbKxvi8ocy1BkkNEbtNqxYVlpZ/bUiyg9VbCtphHL3
VvDvWBtS1bPbVD4K9ZDbo5uLTSaAI5d//h48lkD9NHp3R0Esexwlba1fGVxNxpNl
VvhUhyTrglGYskOTdTdGeW877XNW+XmAqlJFlPmErR70ApR7Jxm8O4NYsbPpJW2U
KcwwHUTN36agQ4Ub2+gPeOOZV0VhXzroJnMLVk/8qokTTeGM7SAxuKx2deB0Qg35
8iqpKUDQ80zBGkmBzUh31vv++sVQ/uOP1cmoxjUtfJoK3XQqUGaCRHRrL7ETUohg
Ghi/PZKtSRbiBjkLJnSwAr70pYX5xPhGPFyAosenKrJrlDFWTZvU3fyfGYR58VeE
1zMvobQRsVLMynZDH0fefm0dTU9WuB0FxQ1UNmZB4z0shqpKnbPqW1cyvyAotTFp
ZLuBSKRFutFH/aGLwfu483E5wJxHvnKXb7+YGMozZTtRkNh/PImCg51AMhk5pAB6
3YHZBHiH2IwG0C0J44vRpSV+eayfiWghdA28uRErChvDr9HWNeING8OMKrXwxYr4
EhbsunZpeyr2vDaR2axXe/HK9TYFKRqBxDiTZevWZJnNyTB1reJUohm5aKOxH5Sg
7df8JgIn1Pi+akHtzl5O07M+Tp8DjDgNarMehItNPOIP1MaJCyZmadDUQw3Hu3kQ
UA5iUW/ORw4Mn/7/V/BeZmRJgYaCiBbnVbwh3Go2+D4+ZDpeN5UDHB3BN+jV5H9h
aoDqyjmXi8mrsNagrMF8rzcMdtev/Vu72qf63YZRMrqte/uAmAKyqeeyL1gqPNRu
pte7XpmktLm1Y/vH3vHcjN3C3BAAGj6jYHw+0i3Rc72OIP9M1TignKOn3Xvh8Ohn
8dvESTbIiatfb1iHVMjnbT+TnrmO+24kkieAG07IFZiG8QbmNfVQqsoCjGsQGMHO
Uhkuyd40DB2uCSvOq8zUHNwThers3YUZRC5FgRfCndGpWPoS9lqt7iGYFnXIs4ZK
SL3Na7+w614FnLAxO37Ej9MHIe6IHgwwpuJUIHn2VeTAfMesE3MXwgHtVzNZFyJw
zW5tkg15+jnGHMzud3Ho5zy0A2TK/fDtsfUp+2orGKCjNu6ptmm8CMVu5bYX1MXi
RonQu8b736X2nAV6Tj8eKf4WaULmhhMPdJ3hAFwGD7SzUmIXoQadwO+jtHJBYI1b
/fMT05kw/MJyPrxh5mJiQEMqnq0ogHL1yfBhC0/Ma0cVkHjAy1jNwks6xp7DM1Q/
BdBhkqpLhLlGOvBKL0mX/dqcYqdpK0gdcRN/lSHO/pjvX+eLn3SmFxTQz98rK2D9
5lriu4Lfq+0C7NRDMMoGcrn1op9UlCKf76P1pP/pc/ylx6Du5MKXISuwqF27auZH
FE96GkZWNfjS5aMoW8M9viVhnfeMeVNSgn+Xf9HHvhU3ynQPLXADYjgG7RoS1ULm
1AfwEYNRpjM0Qud+AlTlZvAVhxsilYDTy7SW/F38P3IpF9BM2vg6bEXDN/idv0Fg
m/BsLtgcZekkrIGZJTWLSe/ahxYc28ykPtI/egdo46m21MeE1z3jEVoZkK5jFsJo
wyPCkb0cABdkc/l6sN1BbDNpvMJS/LVYU5mG9D0DC3wmyqAhmOFgr0+Hg85XVM6m
5OunxZboqZMwpBSQt7xsWRdVT2H6Opo331pnbAWA3hFp2O/mHd7jSpAKpgWn/rrr
5tyFDT6sGlwjeQYih/9TagzN4Vy/DTt8aEUBKRn3jEVIbtwpqiY1xZdHjWT0RsdX
Cj1E95AUxqJx30b6OhGg877SHPo/Ouqf9RIdR64XGAEo1ehBRJxLeUuQrB+BcLqY
8v6PKsJhUlL5/5k5sLBc29J8X7gcaXJfCiCQEWH+VzG3+rEKMrHW42Y6MP5uqFeM
i0+VsUe3ZUD8jQ0IabGWCcPJEh1TzAbniefaJP0hYLfkmAlQ70w7vp3BrSrEcVqj
vtQSzsT1xDIybVFRlpfGMaV1g0TblLMtBnq+dil2FHLEhNfQ2zEKbyUDgYEtYYFe
EYYZbVm75nT4kO3j6BeKhFhwEjanZO56rW1dC+Wf4qwZvHZhUD2uUigswPNb8FnM
rCYnG8tWlKA4c990KVOCpJiCy4erxk4PDo+gjA8od8T2j8yWC24nnI4oDA9371mG
OLy8gY73cmNQJe6E0927S5dC2tQ28rX9afn5hu4dZ5TgeSXNFKLJuUgNWCbajX+A
akKpc5UiPjt9ALGuS0qZAhRYHNpx4NJ28Xx5tS9r9AvmoaecqNjx/aabCu3+ZE6+
sEZ9nZ1DQyUCGZ81AKrW4z/esiSHckA8yTUL0XFxG+GDNnekatrwN+ODoxtDFdBl
/SebY9Rr09YTBCHja3iedZ0GtnBzNFKO4FTaUBOMGTP63vHq6QoVpZcZjCPO2veV
NS1NSgCFKEcQQXHYy+mVLzJIXFfOi1gzzuIid2FPSHAT3Roe8Hs2ZEArw7XUBiXb
b7xPLIqy4HDJ/FjH//eCPA7NttTnjj5snlR+SfYX0j9j8zpNEuAqLyN/EW3avdxe
WgspWbdXwDpUg+bht5NJQP48cAnIPCp/CBNbFp/SklIKxfAqTQyXGj5d5DVI0ebB
sPzR1oP55XNR5o6dotDbX0ES8lDqvzAOner0rGhcZ5iosT4Y9kxKBZNgbfLKeBP1
xVJb9RrggLR0qqqg9U8nGFivZ+1YWKqeK1VqM6EFTyIa+bFwpSe/0StUkuk2B1oC
mHSBEZAFtuQIEL6SLLNNEHaw8Rl/zv5tjKJ1uB6AniS2c7k4rIGvEnpZ2XEyhc5q
/4f9AAMcvkWmAn9+5GkwLisqGvMKZsWGrFij8EHi9MDogcuOaAQbov/T5bag2+RB
2WBBTe1ILRXrVc8cg6WV/Q/VC/CUtJ218YphXNZrE6VPz+kcKeUlzUC0aD8LZ0Cg
YlhLGFzYSnrECrAPUqcum97x6+6L8XDt48EMPRXCJ02QMVL6ls/JdvvaVO8G4afv
IU58ngC7Q8pyUHVHbf898vFGRL2D33G6Ov3SR1ef3ZSd5Nh9iDBePJ1Bk7sP+3cc
mSR/NFe2bf67L3hMgNVVY2QTOeyBVeWEAlxLrIKmK1IGTim6Ng6gheVcWkIhPKjK
Ovba8574FBZcZX1Rfto4lDLjsUHCB724AnNlHzC+aMppw1YMZUxKQJr2Dj2qAPZk
HqN9+EvJ2DLfomOKs5uuYxTZ4j0vE9jDK3O8VLkkewB+AslpLWQSy/u5Q+eP+oEz
uG+Ah+9f6Mj3ZWjTRzQ0SnjqMIBu04mVFAFK1YC0/fMPiXql50vuaZuBZ2RLR/mB
Hj4GLh3GTBqweGJM2DNYh/Yej5UIg4Ucn1RMdIwAx8yQzex28rpRxaeMtIR3RBRL
SfEPSZAGgX7LeR59O39lBUuyS0D8GkvEC8dn/YxnJyMyLWuZI2nh6erqhr2OiASi
xAU1slCEI/8uqLL7TkYOJkazBmOM7UczmMhCtFY/5GZnp6S4sUfWj4nI0bOtFJFa
u/rtvDJbLI84FDxWoIXv8gbvByHHpzk96K+p2Eq1N1RgwXTDzzpAS18KO0Q1ZgzF
KoNkQuJ9nEzut6JrGfYCqUuR1XHMxcgEfVRyeqD8wTxtt0EPIug3NeJ5sp2xYKvY
O52N39WHhc5t2aGed6QoCheBlPIWnamVi67+D/Thy6fqY2ZyqI68lbmR/VRliuIK
LrLR7DYCLjiZ9Bmibt/v3LX4z2Rud/7lOW6QnjSxO27y/7JwTXPsF73BEcahbhoK
ZzXmqphvOVxDehzPvIqhVsRV4ImGkDBJwUTmxVcvd2LmFfFRWzVmSgIcsWWCSIrf
gwiPckLKfeXvwBH6epBmbLh2+TCgTS9ddn7YHkV/wNMVxnJRL2ycyMAyk3iOH/5P
000LfYY+Bzl6Q+0yWz1loZnP8dI9+Y8JoFoHncA7Qj759fJOBmRtPkIzmGEOpn8d
b4AKQo6KEiGtrAyqO887y9BJOL9qR58srrKdX4+3wTediyJa2RtNK8eeRBPOnZYU
C0KUJLqaYSg25qCv6rg/N5FoizaTguEf8XRiZ1MuMD5LeQSnI67I07Xy1zX+yjPT
5MTxhuo/A6bVmT9jfFZO6sAxovrsoLhZVfMJyESR48lkRRDzpvUANbsT/mOJ2UfM
H9ENuXgbsxdhA50JiCdnG7ucIf1D5Wxm4ULH2QhMx7hiw9y4bdBEY71hYkzpeovo
a3S4RZrXstk26ZJ27lUs7Up34QiFoML4I6fh7jY3WCLLgf/cKP3nNnw95LwRPMmA
lclp5rW+aFgH8o+rVOWLQqVGwYa9aLH6BCQosMWZ4PlobVxtqF/ueSse6k4/+9Dh
nPv3627qy0hJ9ef702ZrcVF2kqEvr/tz7Nn5OTWl4ogI4MXMKScOqhrxfUr7cesG
XMaFTOsHWvo0bpciXiOgY3A1wK4tmrs5ekTIv5ajtwsp3Z0522GTSaMX5di0NbJC
gdIPjT03b2m2fdpnK651Ecj8421+EgQiyxxbl37TOGJwBOoK1FezRyVYJyJcZ1DR
qPJjBPnNXw6QtMrrsUjranrX+z1a0sVsVTfFkWTvpHmndL7yDzXhkYj2XlmwOlgd
5d03E5Y94kkkd2xBfQwm8rnNzkOmSi4H79Jq4zCLzXRdVSndW10vSVd9zzGPaoL+
K4EPu8smSllV3fkp9pWr3FzQj1svX5qor/x99yslCjjCRevo+5Xk+3Okc4+kAQQT
R0OfpiZkeiIHm1Z8B7P3pldZKnqOxrON7+IQo32kpPDOJoT8JuURvVZdmZCvAKwF
bKwQksII3R5/RssnSol51xwIA5hUYPgSN81M1U9Li9eN43u8ODmYTYcImREwOmYl
2+06MbMsPYJ0Ua9LAaAGcYvJmnC8g+CpWV0ItGzCu6wJEbuGhnKVuxznGxRVX43n
tL1FX25upSto/bWjeewDCsivlrBMLo1J8irmK1KCQGhp6eoxfswFE6TEmIJaVKe7
gEWJ58FamDqAv52dCnwdQ69nrgpLzfyOJz5med7eew7ikXZKj3u1nyKMnpdJgNV9
ugfn2wyWO9m93fqKsuLvpJURGEGWiLGK2Opz//e5+loJFh/ODCdthjVn59RM+3ev
Z6TN+B0ZDxh8pcdiKq7Ki8olWYupANbI3IYUHMlZpqQA/7WuIbg0ZE2AW8P0GNbX
U7ky894csoXJ/OPFkybylCOEfd9cTA0uwZc9Anx4CmJnoIuv28j1bKEj87ReCrK7
bEbLZeEQD8fmf0ikrbZ2rnX28AyqesHjQ9ajxYe2hJjggTcJPYzgrcgIYcL+vnlt
cS5Gp/q9uC2MO5ma4vw1GWyUUO+/voLdeJbPm8WC2bBpfufH5Y0ptFQ8SxsPNQrF
PplX5/riGbLntSQq/XWW7U6sH//C/6iYZzmrhdG7WmbxEuTFLQgMk/6wv/VjrUNE
liGPnCmq0P/7HgQkLX5ttsISJ6poGZ18kbfk7RwGP8Vm9AkKlx36AGrzD0nDwnQO
56+zlYUa1AaYoa91hB9ZuvumumFAxg/TeeVE23fsuoejWpPvJH/bvuhhLu73d4oI
IhcsAVnHjOzUw62uFgLPT6bSZgdqVpuKh7KAfuv7nVDB5TuI7RdJzAxJ/eprf0gi
G1tD4kjcclsCO4WR0OWBue3epTNloCDtGPFVxoLjuS6VFzZuOc3k99KEOIwOtJ/F
2ru6z3lMbYT1HmXnM4uiRz6g66tSxAVUF6MNsUHQCwu8p21iQ+7kJ6ZbWDg8jpTi
DnRbEOWmJOn66116OyzE7ksg7MqY1GrUxfLBiMA8JhnW9XB2CVigfIJJbVti/MaI
QyrreHMMxwvmQh/Vfx1IlIGSDoXFS/enMoWSas7iPQg6Y+DsED/Xug/R3UbxKlut
FMGAcy9nMYXPituoMHHz/4NuNYVLwoZwHedz87su+HgfE9V9TjIpcfSgjYmD8GDH
rLtGMTgC8mkAsw8vlyQpJwLvm3XS86qJ+/HOSc1A+eHI3l3ujELeiHSB1AonolnZ
PjJukS4BXDu5krNvy0na7kd4X85u9lg0cFcAzGIQpFPsHt/LmmiwU8+GM5nCRyWo
2BzzZByEAJ1ugRdc5gRsl9ZPtioFkj2JWvGrsXVFzYnnJnH4+4QhBmaUNWwgfxxx
9mpZY5sJzOk8RqAxhj4VHs5L9RVwy10mMXcOOrjWO1eTWqecTa3O3iFMTBvQgrfS
7q6pGiXX6MQ7LrB74EaAgsx6dIyMv+zFKpDFt64Y0Cgda/oYOVOS1WmzDZis0JDZ
pu1C98XPIbRXezuaclHpB48mz4r3vz9pjzYSBKYzM8O6xWFL1NDOpWkaCwRQuNFy
1zvzczqI9pFgugdB5mSb8wFt3RplvW1fpzOkE0j0NA0ZPUWeisYKXggEGhJGNAY8
bk53Nq1VdQYtjzoyZaLXBjH/qJJh8WyHHTDGRjuluL/jfF5DyaG4qAcCR4Hypi99
Yfq6jGuTpzNhvM+N2QAFkC2ZUEw7ZfyMI8E7PvP8wg9TbpqSRBnEXquA0MF7DF3G
k2QpUWIdMXBmlwH/6hVNYp4ZoBQv/u+1MKtsNvw0dKf3YPzeS+lxH6wDc+SYNCRu
wbFJOFoGdPK0f+dG9X0pXaQXmYGUGqujh0Yju9MbEgNqeq75MOL3GI1MKaY9QJ31
2/IsktGImgiUy9UNvn/NrrDoZCv0Qu5hYGYIfyMrsOjBJLwAeQsQ0k92XB/76yZL
YXGIVWJatRa6ehi/NOur0TcVaf179ebczGhe/rXiB477hx4DlzYu1tgSlsm3+JZu
79BN/PFhpJwnONjNIfs26bu9udhQyCiZfUHKaIrZuIB9UNmiYLmBMX+X0d3nAhpI
LWM2dI8CPp3/p1fmqfG8L4w0EDvs8aP3lxHliL9Eo49thyhWd0yFXhqPWNAxxEnx
kKCUoOslPZDWI/rKfzmr6HjA6tNzzFqFvsTu6c8MaRJIs3fVcl6B06oUrtHzMRWt
s1NSp6wBhyuFo6PX4PzJZcPAuV6CCQEPy95GCjuH516MW7+CUt+GQ6jDMlmlLwdm
Grx3ZY5XhP3s8ny9p21pMrMj+1L45s8F4KpYOCngDH5Q/klKTxE5CX01ZG9tHV5M
IlclgCGwmjYxEUu27GO8STpeF4B3IXRHzKVxzJfSl6zVvnK0BWmIyza6fI703kaP
yn8Hm5Im25fg4gXIhfiiH2yJAHJlYTTcx1ImAE22FTw=
`protect end_protected