`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 41760 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRmObns8czsvRiDtLMy5tgPqPJJUfbqxHLHroaSda7mK9
qS2YERM0dNRPt5o7iFWWN9VTn2MFCBH6BQgZJQ7GCNvM8AOb+gUiDbr1uk+GeFH7
qTERxzRPOgTZRc63tu5+m0+jqjZUmrybHTTaK2p8MCXGFj5rHjuJKSoPWDGhEIA2
sOBYFqufK74HmtkNYOTve0dWypexw7fm96KfzX748W5P73Y/GHRSncU7NAYkRchL
Kh3HdZu3bgwCUH8PbE6ljN8V2BlkgDKWNc2HWqEls/CbEl/J2LxrfVMDmOQNyaEp
+RlEt46qU4Xj7+kozGfXK6J8b4gKitKkgumh7XSxrx1n9+JHSESL0y5Wfic+9cYR
UzvSIUo1/zgp4C0swCVg57DtEVzcKMQQKcyPAJ5jue/8O0M/zjTbcA9VFi4cfAoP
fJsKqewchl6zAuB2HlAszEXDYxLtXOrrCapo0f7y8Uad321dE38TklTqJQjZzH28
4WOOkRMBtQgBHpOXilsjqFKb9NnQwYNuBm7WipiwiMBQh4w6ZZpZbnZgBRQuO8Ed
UXsbA5dvafX4AwPqyN4E1Cu8QjFrygHsoOireVRDx+2+IULXNnYOZ0hM8ZBJW4vI
I83t0RDJOgNMaaJqupEqApfhAE7uVMggbe3/hYC7ZV9i6uf6Wl3H+EJumvtLF4Lv
jA60qP71Mo69CR7PUFp7xJCmRkSR/WhRYK6VpwEBkTgbtdOu4N2sXpkemjB3gTdl
3JpIn6ZuU7sJXYRM/Mbt+HxgVusy8+5jegoxXT4Twb8ySBGBjEJUDLcY13/tr4ka
xQvVuId9YBURDqfA+u0E5toMucvaFAmv3aD0W7PMnwM8U3im+KSw5novGWWxH8aR
MphecSgYSQZHCBkW6mIDmCvR0tZ35UMy1R2yQbO+CCZEr9Kf+qolQhSSOYrZ6URw
oDo4nW3Xnc8nl7gtw7MwoYOicN+bte30uDiBvCxq+S09OenQLJ627JRiEnzz8A5i
JjeQfZVVrZQa6MJYOHa4Sx9hpdPRZ17/u+SF0ZSLyZsKwh07H9MMpPEyj9sbX/on
Ybb01uVn3UbVwbP3wIax8pYCjxLOps0XVlTgBr63loLiBwYk3vQ7taYcaux9Mwmp
Hv3V2MYiExsB1Qh4luYvFFBIW9Ks8Zcq/6fnld9lkKYeGkYmOedY/L1l1ZUO+TEo
I53dE7eGQn/JpskIUgtyW7ugjd3yO8EAd/9F9RYXaKsnNOphCNQjz0hEfm+HDaux
bcEjyvrcSVE16a3RHnL6D2LDECK9JV4fnPXgl3T+XOuNNwSCcUA9Ja1Zff08QhbW
sx0kIwINaKdlJyVe+P80PSxX3Q7D4x64pb9ngBR4wWIrW1uWbrk6+PpGkujQ0E7r
n3BAYomEonTy/2MQjSqyFpzLS838/Zm/Of1XZEd+5gXj1QrqKDfgBpaQbUbC1GDu
alXVGEGPNhqsuBHyED6425ZDRrdI3yQXt6B8GPCdCvFW//GEERRSNGyDR8YQUpeK
ZCEwcsqa0SLXytU2BWbFUHBSzyNEQQChyRyuSngKZePvxLjvOT6xka1heEKcGM4Z
pXk6tJ2czBINJSDO5Qg+20r52FnMHSHrBVbq89raXvNHcrHoD46NEUvBl0OMgEzQ
olu6jpiZX/JqX9FzLOPhdVGJ2aHH0hSLEUZ7vYBDTEA18w2DOAoCbK+1OZCJ0Nj/
M9ktIjgaVaAvSjbySexuOSv1jnDljJzjOkm0vdSWDL+96NwMIelZH3j+wA2vktxD
wzDJfK/xKzJR5oHLauwCJ2jrnZrN5Sd0XmAYplJLjCk2QvmK4Y9h+IIHMhaxg0n6
w96oMpmvuGsJm3/k+lEuLY5+m1j8cElyaJokL16PldLjatGUc3auvmMIgB9CCrat
y6Xpudp2nHnJANWLxapZsA8+/h/jQbM2KjaSPBwN4dwcCruToKSag4MblTKLaSVZ
PRhERoN2+MLWEPrAf32qm4eZi70PWhJfC+jJp4oTsVaoaXlaaTbq/eEpzqPd6YzU
FmNO6VW6WnlBlbWBEbHdN20r0CdaNHiOIxNr/mDPmT5QYq3Vz4apHh1ffIYBOkkl
2hCxTPqcogMi2gY/1Rgg7ymwU276FveigyH1oCzcuz4U5Gjvn3qTPogelhiQWQxD
Acj4KeUZaI5aOADVZzQoSyAEW98iniH29EPikwLUDFPIeOpFOayjltFGhCW2M1nH
Jg/UnnIXPjs6ELI++C2FevJx8EJRkdNaFl73nIyFVKbXlSAWRWzdlKXS+0tUO8wl
pCGpnWa8crSrIEM1RjZVqBP+WSqoI4gHimt1PTLJPV1MuwZUyX68CmtLB5rttvzZ
cT4uyTThJtWu1SuEdi0bbFUzzvrUInSnd+8OUZ6xYl2cBHb1Z6o8K7v22Zp9srZq
FvFTIyu6s5hftoCUxDINFFtP+whD63ru98eqS8QnaXB5BJ1t0u9nTgw/JIQDeXLE
LDTvjLna+A2RsVntxptvGhUvKan9MVZlK3KfxOLsdDWyGpgIAiZgMal5qC29Ms5K
q4R2X5Q9WlvU3fua+LT4jyLDNyu5xCZ6EqkmCXXHTn3gq1iH9fc8lX5e0nZuho1h
yLMxxEGoX6Q0Capzo2VE9FPWZEH9zurnTSG0Y6wGEJpF7CHkbrdpqXKGEnOMzW7+
VPID/8cnFGOGffEqtbU8YY5d3SH18YCxOIv5QK2cstwHQKXbG2VovJNbPfPyol2G
3l5cvI/ZBU8Mf9SPMb6K7LwFjp60MpChAERYHu2dxrCVgDb46fUsastoaxe+ZhkU
XC6txDZ31G3/9t5+h3UV4tSdXEtsIybSImS7zTw6b7FZxWdq7FUZj6S2cJMZJzlH
n4URp0jd2OXrYlr0RQujwLKSw16RN7C3vR2sRYsTcdw8WsV7LfRiWdP6QjGSbUJj
AJu2KEZVHUL81bIFftzSWq0Sey+v1DoEvv3sJ8O3IwPkZjW1I7VSB06KaJW5s7EB
aYkMnooEuujYw3uGqNwnH1Xpsq7O6N8czPherNgWZCr0oo7J9h28yY+pQVBImDPf
fRvRfPktzgmypRQ65HLN1XVrgIxrsFbfLLuPqfmqboyUJ5Etq/c5CPhAeqDssKth
eW3sdhvZJmkSXqQ3yZAgz+gfEKbRPTWSanYckmXb8X44nDmBxT8zxhlWndpF8RzD
MHsGO8tTTklsAvHkqAJ6LQcvBV349xuuvDoH24/cnqnbdsgM7GM8nYuDoJrZ2/TZ
4MrzQORV9FbLcc+YBSCMW9m917bCWrCVqAbXANgv+/aoP6JU/nahgdo7HnidFFi9
yO0+PFNJEOXlmOXMpt10oxl8FbzjuBM7oq6L4y3wFzrCrPou15vP3vW0G0BYmtir
b+2LhQ+y2GkWmzGjlZi3J992tvlS8bSszkFZaG2jRl7qQtTvqlZ3EL5jx92O/1xK
87Jrqb/AB0bG04eWiHWTjUUKXTb3+4TJxactOtuidPfzZKC1sljShqTL6X2F7+/e
RkNkTs3BLf9RnsqHI84V7UbttO3lq4uarPAAqQqKb6gs6PGpr3/Usj5O2TWxOMEE
mDNd+2M/oFf49y8jwHHvrYQKucyiaVgudqrqa6tS4Hihk+2oFQE5hp6XNKRcwOt3
GlSIsiJ0yCbo+trbBLXh7k9nwy3nKJX1It/9GagNqbnFifq2bpjxct5xEcWiEBiR
xn3AMae6fwWRrh3PmnlCGOdQWWQFh3vpAphUddq4jy9Yy5kSxslSZsyL4arq2VAV
cCiSzOW9hJtLFWZjtOk3YCaLr5rWlBsuD+6ImmIQKjN1IKyBQLH3Uj7VPoaYO9qo
Uv3nENvk2B1aqT/xYmCQJ5j9eJfXm3q3jgWMFpn4tGVIxA1bwGCdZZ2yQHWO8Qb7
uuHUrajGU/O6aiF2VmOOAp0zwtRagPzq/JyQAFAsROteC0cVAaf069l+sT093EHF
pqN4/JyS7xrQQ7HAb1htpc5raqR/Z0WPuuqxJOQeV/ZqhULAYE4fKTFaFmCk97CJ
w2CeFp1bWMWcMmPp8G2tpTrf1tzk4baIkWCZlFk4U0iHllqCZhcA2CoMl1YQmx45
WEVVWQ6aCmPDke2545EsPWZLW8l82fsphG51IRSYjQFfmmIHRQyImVI0UaUCBb3x
i3chA/l0rVqfdUKJAcAVaG1bI6jPKIU54w8Hi21DfuViDIwJyupsq0LlyG/K6+AQ
dz7j4UtzG8CjcuexsghyuezAKXeBNDMVmDFTDqTIlY0XixG0YucBNjMki3MJni0Z
cJn9rtdlDqOY4heHGfMYnnNBeqS6wR6dC8Gd7y8hgyaKW7EO7/853nI7DRV44FlC
oXSQCYAfsMV4PryECmR7Xh/Ae4jOOCy5b7UnOrnv7WeYfkXKNbgfIlIhegKfDa9R
hRHTnE7XznRgnHT3i8iVpic7xrM67sfxIGoCkFu0fTA2+PaTl3WLQBH1t60ah5bJ
sb2JiLFUpWwoebWQRB3VkXr861hOeZy77moD6VH4hBA7ly5AcRmTtLHeb52WmA0d
7f8ZV2uNeYlmSe6dmGmPi6z8aag6bEwbOZ8gGgOtv2GlohUzUfXM8QZgGZ4OYTKE
K5zAdEKjaIlBUol8DGc6n7+84thGwCJ1z4cAhdYOvpI6BKRbTB1ZIlB0bVzy3Iq2
t+JWDvI3kfCwXR7PatD6f7MQoyJOfftVD6k2g0Oj3cxeu9wQ9bPzZFh7CrnSXMNI
5tk2C9/WPoYMotamVtEL4oosqt3ntaxw8BJGiPMUOxPLTs6fEeS1p85aCsabm2vn
T4s/HDRmTsNnwOO3O4eYE9zRNfodGTm/wsPtG54f02Mvmx72Rn90uZjNA4p0lwKj
MZrtnBLAXLb8LYCKzD2qnS4uDHnkvKKYb7X0K8XdLD7OMBJ1HhGbm7aWEwAarFzQ
7tIbz150SoMwfR6hPLGW074JmYTkKdTJle+xbJrAQs2wpHzbTCMjU9N3HJPHA33y
TACxWFGqwH3D0fvuJErCe7bGNafqu5V9NWdwY+YcDGViMhgMMyP6rvGclYtmJCjs
Gee0PztgkolBk0Xt/WXoFSN2v5e2h3O7+GurgZJw0Eqe3P6TSilkoB13NUvrPVbo
uzrQGTQMXb7LYoCuGiRRRRR8YNSKK7oUCI4RfUSJQsqwkI3/fm1mLmBxAzq6H+mI
y9WU2K14SBenn/3/Z+hEhDhGxxY37/Xa2b/1uhnFuUPFwfqCRxjOloaFsf70QmUl
pIhpUFPx+yxLi1KQjA7yA2W60RPJ7Pmy4swmOhEeUMd7n3HFNsN9ZgHALvjS5fo8
WKeXF4PXiM0iccOPJabpdZJau3lTcn9pziiv70zL3uX5iPbrAI6BuFASZfzsSqXg
6bQ1XDlZqCszVz85kLoq16PGfftyXkscZf6/C6xaGLVGMTLt4r0Nph8o76RJ6r4J
xpxoSl+/uMAOMIXy7+DwiOLStWGPz2JdsYcULND+uz8kOmHM74RormCZUXRkQ0ML
KG8WsQVpjH2Z8tyxeszECeDKMJyGV1Q7Nc/DyATHu7oWwZ2NCl7DZvRZnPUdXtar
O3tk5WdUuBMs5KUtaEmU5mKn312NJDj3ZsAmTzvKc8J8VRxpm7MNAiUV7yGQf3zW
w67k8Vt5LISed9Ydvx8LFzvClFtGC6d+qaQ52hCfd2OAxAwmfUe6qCnXbgV7blyn
83bU3sycWfdkK2XiWc9lc8hCsjTmipuMurNfCwClYyFxfl27xh3N8T+9dcUDcmP/
xjWNXraVFKEbQr6xEqfcbYMwHq3LeR7uZwcYhJbjX+KOU//Lx9MhZsmA++Y6ZC4u
mLBTopyQYFBsAQntJ40Vg1llsfEeZB3kIZravms7KHPjLK2nxA/TFzQ8cZmW1/4s
w6hYvWdfBHjLVGnEg/RVJTqBxx8Wuu5BNo+o37qMUNW7ndmeN6n4iFL9AtNcVHZ2
vEIYOGpULCjfqK6+OWXP3pyaG4hmi1eJqHeSwnKs6AaMQO2TcipyJPNGJH994BAu
fQK0tbystIRzMkN2+3sO38wJkYDo2/oxoy6Dy3Jwa/8Inmyd72ymxdv50/cHPP2F
Dle7Qxo9p7pnSzjSA4R1IRMlsREZ5HlGSjOCjOTFX/linqd75IaMy5Dk8f7i+asG
iZo8StydlhWB0nCtoqvkGYzaNblYW8khlzs0wZTHHhnaoNcS3tVvmEH+8dGMy3NN
6Xh7qJ/U7moSdWD6WTov280wQC5bTtpbnBA+OTb6O8xh81bg574yxqYwCd+BCwo7
abI3tqS9I6waETJMBp5w4yqSPKATQNKouVr85ujCRhtvWGN4pBZYPNd7JPrtRgzc
9Idb0j22Wrvmid7Q8m16KDF4N8cEnxorhCrceq0FHsBS+o2HRzj8lYo4mSQdYp70
y3B1llB9TtU0WZp3K7gnyIoahwCGAPJozcuW5WDN6WdNpDXXcr9Q1PsFM00pDECZ
ojY8XtDIgPjyqMeYz3brghJb9cy2fl1PWzbS0Q9V2Hn9Jvyktz6WmBkO9LBQWueu
uwcQlXDmaqKXEtGwYH7Q9Cb3Dl0rWppdQgXRtQZBe96qeenFs7xeF3wupKZa9XFT
NBAJxg2O1BAvkR9q1pjX6VHs+Dq1sp5uW2FRfgHkJkxI6BO0XA6PIvMVLLVVi/lS
w00ULcg/Y8KTzxVi5MniRPGpzWR6jlGYMcIkuEP1aPWgxDkNxFTozPg+E7k/Fw10
gxR9EeaWJm8mz6lkCFkIMx/n+MhVmMhr9iMUHrlscX0uFpTwakuoEOWzQ3o4dY9t
jDnM0WZ+6O8ICXrbzMlpARXu0L5gSrcsDTbghPw8kCDeQgPh3wtX8t7wvPAby+8F
Tt1AJjvEmArVCc1m7MK9bX7+U7sOzYezIOYXAsWjl4WQCMcFqbJH4qyrmSUN+8Dw
ClaSgcoFItTf2KLm1MPysZRBdFbZ7IbVIRdZ9iZ7+PyKqQe/J+1eH2bcJjGWCZ/O
OSd2gHKTaaNJm4TbGhoucwsyYCfYmBiq4rHOEFxlkx6FyELiqPu0JcgQlbVWjUOj
oy55VJxsq+RvWHhLfnuHBIWqOyEXp37tSJsgq/8NEoPmQCZhm8Vm3tBbQi1eBf0u
Zc7Odim4KKf2TGBWbwynvRHbk7WDVQMxEJljHP5jDhI6wwtDUK/8bGo3K34E+FAT
lqLM8H1kJ/frkyCBdKXpXFrbS7xpl17QkKBufoAM5mtYhAemJbb1h9kfCUtfBGwO
hMdFiwpLcO+GONiXMR/F2Ac4SCHpPE6pDpYrDAIa+8so3iLLTgLlEpzWjf21NDlq
EMaRySiCztVEGwcyklVSimTSRqPDx/ZwNkhJ034EjE/+nwE0GBKNcCLa/ZY8BhJj
P4v3mnsMO0fEjXhZLe1+ByJLRJBbIdHS4eoSEWMQ9v55HV/H/DhscCClrWuiEBko
KEp22meVqKLqU75EclNIPwtQ0RVe3RThYyzzcv7cz2tyQzY4OFJwwCQYBLD6eoRr
m2UIXoFamWWUIDoojPQ/vodoBVS/wNeukyP9SsNNaa/CJxl9rvO1qFrUrFSAkQGE
b2O1P2BoKRZlvPVohe9XxqEr3fzJOMx5oowJg1QKlIxa35Ymv1sT8WLTDhJmm6s6
qszRiNR17e3gIOOpKaPIGGUwKeu2zKhoT+tiTDMK2HXET4tAkucQGS4z6304P5Qm
sMsfiwjucjao3+3PDo6YfwCN2K6a7ugNv70SALBSyr9wv2PSqk//gsUewnr4hUbW
99VaajHBwxhzWurnY9bxLT1tUuQr7Rfk8e0QkgNYw1/uEziJsyR77NOYi+G2BHth
2fxuUlJSl7S1K+NDcZWRbmvm+wXcLT+UOf/TO3OmMBoq5MzNYHM3J1T0c/xB32Un
MRhPWA+5cIiqf4UHw8bjLe1UUVNGAvy3uYqr7MA7dH7+6pmBuBs+RpL6dlAgkUdd
kH8kNYd2n5A51XeDNa7SRkjZbOj4Gt2xE15Fpnf9A+e80x3Fdnwo4bNPDUHSzKxJ
4e9NxSIvKX5DJsnjU8ug1ZGfUvCIrRYu4WPFYJx+Rgpyf5GGeUJ0344EmSzDjVsi
lBgRD1OkgfTzSQ4MZRnsysRBlwnLVLsUGLHP2IB0uOzx3dvBECjpHGg5SEU6tuTX
Ugxa0y9ZN/40lThipn/aWfCQyyIRMpDhHu6aDHjGDK9gY5O/QcxX3ZeL9MDYp1ug
XDfQdaXVFGAEOHMxsG1CDBvUi/MM421HFYVD9RgduvUeH3lb99vdq/QghZkfo+Ut
I9WBF6Rd7Sa+jyn870S/1FHz7PRTynnTLrVwkFJrYL5w9Ca/+9ZV5YSnrkJ2UNA4
bCIt9tWSXFL92kbRXCweT5C6n+YBq+3x+Pe/0PZTZjctJb8NZDANGF7UsM3MJWvu
ito/FZ6yXkSXdwMr+QPvXLo68M2T9OPveZ3Ybbad+dp+c7x5XfoG2xnclFHCxsm4
OeSOQAu4hj8zu9n2JakltrCAkqbMrpOs8QL5naWxqIjrT8w8BItEr7eldbgfxWtP
6+oZ0UfscxfbeIs1tTXSpXmgIypWwfqGHpJXOWseYDRfZV+xxXJ0Pw2PnNGJ2f+6
FHSW8DpClja/qUM9N6rQChQZoR1EMi2oz570Wf2gk6dqwm8Q2OuKBAF+tW7MyfJM
JEayrXRbkcAlIslo3LoMu3okJQKP6bcB9Mg30NtKN04TYiVQe9nvGN48aYlOOlyQ
+sVN3Uu6edHIgKnP46mFlGmYBzX1UZR5K2UWyFulGH0O12RvWLbGrKnZR5oeUAlw
1oC7CUTBmvMK4UkC/nYfEZzB/Xx/M28ibinsDQXfTaoyrzXAYOtIrOp9lzFoRxty
oKGfwBvTmTaHhTgI4w3G/Mq32+/6T0FHkX6N046cTSmVKhWVMumLrilT9tiIQRk3
kGQVFp7p6qvfFm+Wn6B2fLywghTJ2YPqTdZjFn1q1W0QxKOFtZHmQXrmEgSdcWA0
NFgfixA9crhCmZg09VjZzoXgVjCRcq3OXr6Gv2x5cPBiRcEPpGiO4RUHASXOYGi2
T7VaRMjMffbsE1QhtNxLn2Fgv83UnoTCEJNrtSrjuUcQtvVhySnped8YDe0x3rSa
Pd1zBChGnb8Z9LeVngtjWrqWK5dAMdtITqHvWbfVkr7+ez6PU6qfKDpSW+uNOKPn
UQbDbdzmjEK9C9dbTWmMRF5aKE0Y/DzNYQBOb/SzdHlaO7m2m5AgJzMmpFOIiJev
Eq4/YTvfmzJCfDpvI9B1gQtjTmylodRh7PVjaRnTY4c9D+vyKKOSlXWtA8hJvByt
PnbPXZ5MtlJKVz87furRtruFD0zpbLR1Ft258v0hj2uCVmup21LgdRdMuyA+DVkX
BRHAjm5BX4YN3gy22xCm1NCoepOU31WMUh7U61kP/kvIij40zo4Zx2X96bcE/uK3
MIdQrZtMQX5RHgVEXaHQmTas30Pkg3dd2utIAotd7IkSOLUcLDUnx/Sq5nkbYD0M
ytqE/gpsgfXFVzF4DbdlaagUsrOrCrbyMgTDAKQqO46ipK6kGbksbL2GHOozNTqK
gYBHGfowqO34V5UUtrcMT60614zoqxxrEobzykllRw8/GV2f8hOxQWLy2y5sdP49
1WFpItvA0QEIIk7dr1NdPutg0wjY++5+2RS4OG2S/pbzZzBkI9hEUZtu8XVmLH83
M1ah9hWVHuCbYoinfVbt5O9JowcXz2y0JAvDeWtZSWZlNTPeki6yssPdpJs2NkuP
9Bz+Sarw/EmIb/7tBJjUA9jBeZrBLdGUaR1BRzcZBR1AAdSBdTsX7w5f71kgBJoK
HNlVfPMT7fG+IFTdZe79KkGwpQmitpnttxrfYI/HLBK4/y5tittrVR1kwn4H/Vey
VNBKF6sPYDeSteH/gXaEx5ryip7gTtFwwB+F1jQkQm8NZKAIZKXuH84Pn972MlUw
LkJAhK20Qj4uJ+3J46Uz0KUtvHiLVbPL+0kktEvFzo+7oCOVUMt5UvPjt6+r+Yde
hGWbKUpBRQPqQ4rx9C4b8sSFTuMEpa1XkK8GpW5FDE00gsizbGRtJYMcsbWoCLmB
5V17y390B1H/IO4XydFa8MS7nhkPMd410Cq0v5Y0Sek073dlWnpiAPyxe2tfwP81
ttqehRiihD+xzUACq+Ki8DET1Wk7CwrWibT8zkR9Pe9/xeAt935l38xRtwiR6k2K
tv1C4ywxKO6gUpJYH0FSt6ECC8qNYNVGSSdAJAvB7mnrKl85Khib9ZEWYuJyMTe/
1yCUmsAoIBF0fEPHLEcjWgsp7ZFO5wc4bnodXf1/nRkYne/FiiuBRde0GBzm26pe
vboR9h9iPR6iKSRB/kKQP8TT3uOX/wJ2XATfEQCkqTNgovqKpZGZbgJay0Guq5oX
S/5XS2Xfgxi3Gp2ko2MadADC8w/e7fZC8WLs6GbbldZaYvGM9LFQKr2VurEhO4LO
eQ/mTWu0QGwO8MFTW26Xcorj5e5LeRL2krHnZwpEnD0R0dCv7SxR5nVbxIJUeasT
wmjYYhU+3TSNWczWmJ+ZXELCxeMHFrylzXuMT/N65sinpDX/SU0NIRcCtnU5e5xC
1ZEFfBeRToSlVGl3uH4zXf5jmhTd9PpYh0GLpwVoWYHCefzZmp9boavczZ8MpTSE
oKR20V4i2AlDFC58/PV8KRNxhSa55/nVN5KIZMjNNA3bGRdL0P5IyMLA0KnAkxcH
uu8KjBfc6KhqqzR5adUcdFFLpEmJ6EhOMWSXzGfF/+1FZPs8liKLVyaXx7pzH2Xs
m7xlTxTU9Khn+xL21VGTD45RO6E16JCgaJVpIOjHLAZp4ElOg7c3LdRekX8aIo1e
V1ABN3hbxvpxWReY8rH4IjfEf68uSKIdhH03gA0EH4TfQQBf/vtnIbFgS2w40xZQ
+PTcPlx72qyRm5IfuVdNqBjQe9uhXRSymNwxl0mgdMs9kSHmCbMWzxEFhaPAMh+s
RmhURLJWCPh7UQWt6lIhJWGfoc+llHVE3i9Z0WGQzA15x0urguLlE1u8tsr0xdJd
+3573aOohI5w9P1PomLiYh010AONJ/pmkSeauW23ApyGWZ3ATBIL8uwb3jzasrux
DiwqMcQfewH3wkoo5QG2cUwVZivOXeUwPCy2kXzaFDagrZW1beXWBzH9lmM54n3t
XLxTkNxz8aiWbXw4SqG5OZ54ukaEQ+r0vn5CzcAV18GthkqsH99rstp0cVnVpIAx
SWSvs/I92GCzRnA+l5ct72pC2+xzpgdQvuJQo7kJnFidueX3n5xx0lPn8h2OhHya
5iAPr+EcaCzAK3WkQO4Z7vtPjQz+38iFWNTHQiz75pciXgCAmSuCyxkh9vRSmHIt
Np9neTm77S8QhKcBiZdBLqBytpTZbfSMDeJFSV7eqz8hjtPKBi0nk/bAjb0tKFcs
1hKEzzIGuKkdGpGcDxL41tCglE+82MKmLVkCzgocFo/QVH1Zo73pQFQGVlBX+XMA
4YM3UCKDPZDrCA8GQ8Razis+LcVzH+mKI2Vz4Rc39gViADzD2W5OhY8b3nhCnlIi
PTSOBcmFsRF1LtYVm/ETCBssH5Xck3BQhNgFtZYX77fm6HXhRorsdM00wj5mutRQ
5+lDQw6bxAED7MuDLZ+4fDQlRkRYjDLYR94aYBJ+x4jeOlAxfQPnS4+0Ap7C0SVX
ivmMP9XiwssKMceLshyRJgegg8Wwdtk/Dw6X/oZEdqSH7VZCUisdng3QRxFornB5
3YmJ5egNQeT5hwbbNAFoB0fHYLPpfH7M6yFZxG0TgTUfIfmzzQTJBzw7zuyNrwEX
dzbjTSYm9+AZpdtU/o0ifoB4WDJi9SQWZ7DvUCcMT3OIl5218RKgH5uoIRoxy0pa
h8kUTyuo5pl/4oq59jD8AIzYc6Qc4fUWKQRnj2EpwkdV8hNHRwhdal4veSsncRxX
VaIQJ5CODE8HRVs6OLMRkjEjV9QWYc89IFx9WBxpgnrGRaZeN7O8GI3hAvookc4b
vpp5X6eT3G/zPt8IEAh8V4WaK4UBQ2sUPWunNOQp916TPOlTI0UjOuOiEzPwwwY7
hsvRvVPV92vUuVIi2yEs+OEBKhN6uWMEtLvRS/anfGsMkQB6m6mA7yCAI38zEcip
ek25iH5jq7zH7sVRExbTaogWxmeWP8scAiAomNNs2XKE/7tVDpEmTPcGuealMi92
/ppfmd/coU0XjKZ58eHRWqq8+w3Ua+FLQB4zSEWNmV+G6GGz07tZHH+cOZMWfASP
tSoDqEGHL2W05oxadZSNSzlQjD5oZA1iJaxbxthWaZJk8/vcW2Rl2g6J8pkdxOJz
PxXOO6ZHwu74Nhbb4ncPJQ9BjiBRKMB7Xd/ppKowHUSAB9grg4U/BvEpjItEx1Rm
tD/jJiO+/GsAmWqYfjRstqS+27JsZdyeZ5FZDCV+6QOoU5OG+mcI3OP2y1Jh1b3H
ghGYdYhZqpW0tqyPZt6WlhtJLm82Q0XyQ0008rBjC1+snk/cDXeh26mZFG9svDXA
eM6Qz+8Q/MEJSG+EGAJT5VgsLCEmwWOFB4gCTeWV19lsRIkzTqPjUgFgdHmw1WTs
nTTUiIbmjUrwKl50pdvVprk17a6pSu4TK9A8p6jnv9TyrKg8b2+WIL4uGg27lsCa
nrv28K4MsRSrxwzRpmKPmun9GAdKYokJqCpGDzFJ0H0zvc9YHzvURCwMSeOki1ji
/8mOjKmkkW5CL7+iKOwbIW26BhwBOagIYSnybU+G92R0QCRwz9IYPbbT0CgPzB7D
rrFWtPH2A2NcLeoSbS6Hagrgen5VJznUCtQ7LjvFlXKMjGY6kLBtABJQJqh58Hev
WEbXODOADKuMnE70NhduA0ZyWXGhV/eVLrO/58yJ9LDykqunf4b47uBRAyC/S1B5
Zar0myiny0Z+ucChNEPE1TMShGvu7bSf4Mo/Zi2kt/6FHtxHh45Zk9rFvhGfTGuR
6Vv5+xvetRCd3dlUmbuh1Cjd9bBVS9yoilohEHOcfSXN3j6DScFZ5NNSFRq06w4K
cvQA/9o2YLQQ5dbUfdwkoUbhK3AusJur2m21JkpFNXEpJDr0gH7H79NkEHOgGq9N
isLKnPX3V+4FWkrqbRPkZCqE8rl7mbnD0G0eGx/0ekKHcxwyFThmADCSieVO05GI
UNaZBq7hc75hQH5n1wwikxbMe50dkidHQqNf7tzjBeez4p1rlrC5paeAt1VNWGNH
wKV0fbZ1JqOo39tfHnyW1WX9RerV9oVgPukVZqjF3rmDp9DgkeqjKWVH7zm20sq3
W0uG3veaXmpxMwKUHSfnT2ZgNsYWqd1W0L5Ogzbfel//Q3eNR8Kt8GnI5WUADwhB
JNWn8qI739mVGGFApp3Iiw+nUv5MT9c4JYVfHjrfAXGBDi9BGLeP1u5ctJgAl3XU
zWdiq4WXOuuqIcGnd2ebrYQovhY4QoaA5y21W7cWe+FcCNL8lVzY6unmSRMC8qQP
OEdG+/kcIimDVVhjhqX6owqht3EpalsQtX4AwnSL74NKFuAxrjN/pctaARY8hxco
2i69A38suP534nTsNSaJVwIDTo3bi7yPcKmyo0m8mycoDtxeGsFtfspaXfUpHw5n
cIv8BH/xVwrZOdSOSFc8C6sVNv1DJvwJvPaLHCtG2vyssDBLnapESybf0QOG6Lio
FkDXvl2+c9X6K+tQPA5Km4lRONzXpSVCHhwRLmi6hNywQPl+FjJclvdOXnSyCVzc
4eA2u6VcmpDHrAbUrK9pnJDNWrmhguEsXsKSutqhrvI1JnsnACK+JXJtKJCfEAiY
x0Am1eNPC9R3TrINHvPkkR1yEVQxsCDcqqzsd1ibcrgNqkY6zGGi5NDGZQzHgHZ8
LfIxvhELS175g+LGTQZAQ5Q1sfnuzGAjLEDQlBXGBr3NW6sCR35+3CkDWSUIUUFa
da2qZuIUvj1Nj+LXsQhR/XNQEWGekAsrts1jMEnb/0ezmWU89B0p68/oBdQnJIwK
gBHN9HbPCNdbenadl6tIMbS6a2cYW2cKd+nSmGs1T+3KZHvi+2CyDbjBHhv8/Jt1
9Ks6/T6qHvIjKAEMiYqDK9Vy8U1jWIFgKN7iJ44OuwB0/xj6ktH3ODpKoqLJUb85
qyiwVl1i31H7DAwXQdeJSx9Wx8a3fptWE+GWBvzGshbXbm7hHXqrp7PWpSm6SK8U
9eOCDXaFROIIUwMPL+fDEMrnF5nzEw1LO9sfALd3fLqFhMGNXW5fiv8iQHzNRenE
fsLg+wQyAR68MtCZqCD6C+xUwEgYIRYkiN4sHChJuwzg82qCQtBJJ5Y27jng5BlG
lhg8b52s6Nc+/7pGY3eNnS6cD0/Or9dCfhzayyQ+TPlTHouJWNJbc1eQJejBpwxX
lpDNpQJaNRc44hgctM1Ro4yfPCJV3y0/sK2ahkbmk/tx+Xsrxy+1OuXyUjtZCe3o
8XVZNLAvK/92CjScWhUixuDE9XZuEbR/zPG4RmLPx11d7ODBOEvKYFLIhiRhyDeB
lsVpbih7vIUwIgR02t6UPL46rmXjfoQ1S6FJQrNQBCzJLcZpNuBEtlPxViOX7VXj
IaP+vOn+SqxCbvbgeSnsocvn9sO9GcblEqmaVSfASiawmFswLF255mBHJqZ2YM3T
wE3Ty+ZZW+udblTphSJagwMoLt0ORuCmTyKsTiHHKuwTS+/Zxxgonqvz4GxLIDn2
q6qn5IF31TrhIUhNM7JMOBHTcFuXW9UxfGuWmCFykt7zp6BlkJvnpAhRW+rhPj/Y
DlnoiApA+QuVWE8HXXC8TWi3SpgRK76rKe/gJPYbnCVkjs7Z3E7EB+eH66yyMpKC
mefoDWFRQh9s9jCIuvr9MOHADcNKUv2rANpaBk9K/lAdJX7/58YKLxvxXAD9+zPl
Ikpt1431IdwMoAJMKfIseBg5ZuWIWc16O1T3d+hgOPVzST27P1AUHUvsMK4t0k5/
BnW3IzPxPjhLxkNTObZ1B9E4mNMvzsMa+gb3uLjy62LFRtuQWPPOoppl8zaebOGj
Ir1Q+Tlyau+XAL4O1Ae6LrhFynLfl90//yUXIRNf4CyXTbKO1U/sBY6DKAxrUolk
IgYAKZVshUJkVwcH1ZyEi+crVP/nPMqtIb2f+41vjxbWxE+Mp2r0Eb0MTs5nh/5O
tX+NCP2OlFbGJrBEG5E7BFjo9UvPH4OlW9Qv0JcoD6GcQlWiFQwsed3YpSHr8NGT
EVeY16V2gsc1D5WW9it2VE7Ng9r450VpLGD+/d8JSN2GMp6j0A0dHGKISyVLvKAN
c8iG0Ujb8WmdFa4HFoOt8s4XdXuatdEIQiiobX1/6PosEAy3Hxkmp91/VSpcq/vv
xSw9IDlH78uhTHZTGwFHZVeMdrDn2ZFBARl/gxylSFOBgdu8E4Eh/inSGqsyXW80
RlPzbKjl5YrjXPttiaTWKAYq0cP9oIj3pvN6WuLN3c2zbbgSXy7ObTw2fRcuKPR6
SdbhNXAIrB2bKI6wqAhBNbQD4FLW17pp9I4kBg8lAYFjfHfj5bvitILbtoBPRvw4
gOPuoxpBkY6hnBSSrliF9lzEgTMW+X0gte1d/51eswfGO4/PnvwGoRV2PVKrerdd
in2UmMUbO0BhtA3V6WeeDRMwGsoqYHT7eYKpU8x5CtOTXw1rwbN8zx4Icfe5XZwE
f2RwYzQUu1zz86K2ZIbTErX6azhEMc4rAo6FEc70bo/dhCV/utXhuCNG85+FYeVS
UDNBZNREMvDii684BGS5XYRjCxusiqX4mv+3X7nvd5bqXsi18dpPH1XavBw7UTch
jNVRkmZX9hGjXNwoLtFIePKbAihzsZFCmcKYU02BXWYce3kZgYba6pMWudnzOrNs
Sad370uf+gwVymD6zKdTE2nYMPfJBqNrnUwr1z7Af/CsM4IeiNukT3ZcnLpR66RQ
3FiQ8h1pWv48JOKy+QrylzjRUAcW69jtzwREOLCVIRUOXM4XMAk3J5bRmrSIC2yp
f/9k1oOQIPaAIqH/8Ib4iP0yW1GGyoPBNReOoylaPKBhfD0Dk3AFaO56OT9cJpwQ
4nJdWcLZnbF+1998ZG7Eh2S9mQmrYmypg3UbPr+ePtpfZSytvqRHNWZ7vmmsocko
AV2tXGBMmAqI4sbKcNhLUOQlZWoxqarkehoN4EBCMhFAU2zEhOBXZjHNYPwu04OT
Pd1fqbvShHp3Ce8AlkntaNMAs8Ok1vBbnSbBAUOuz+LcIiZrUzeIPaG/n572bGrz
DcW6gGK1wvlqFvWmKJyqR/0Q4PDnNGjjb5kOi9ukBgkuNSgQT9uX0CCk3LMMzHU3
SPN8doWjXp+8gY8IZooirkY4/MiDK6HkRJGYMQQwkWw9Iby0NI++CsCwTjg4lrz7
srtf9Blh4lNNRg0pHNrE692raFoX9QP9af6FOhocMn56VTBhfX5ykMkWwSmqNIUZ
Hmauqp0h544bZuDo/oWJGsM2W4tEU/Y7r7Pb/KHdfTr9q9zxFo+p8oKCW5mP0bZi
el2SwU/SVnWxImogJHLmAJGSzRYgOoLQv2IQPoxEFwgD1zx7VLpt4ylRtLLeuqJx
ru9DajewQw9av1r9utAG3i5IZVITpBFBl7wEMzXjfPz7MWqZPYlGz7Glnc5/D9pp
w/wPJZKsNOKJwnJtJXvkSYnQx6yjc0x5i0UP0fu/j39Y20CbNabe6mfVU49CvwhG
HcB6S8PoMoE7rOR8WxYFiiiRh1miLBAPhVtNkw6dQOqxIIHfPUXVGGhuigeJ78wv
MbClytx0OzrgSiJWeIxDtjtIPLQTLeFNFZDFmKtWowyzXwPiY7OmixX/f5Fxct/H
QZv0znSKlmPbaxa9fh/opWaRMrWdbRVAq+s2ChU101NrfnhIeeGnwWIdFWkup148
Imn8vYTp4N1FVL/xaIlQMqrjG2BVwvBfR7qmsieDI5r10Sf00+uMkyEdGyHETe7w
bGqLodRUJiK3zMU66kF0rkdxWY2HEB9NJRXWBmNo4VSgV6SPGrYlRIY3ZcxdcWhY
7/lM+8rzTYhFIw/kHJt5F4h+lihkTzrC98Mxrfm0nu8phfq5PijgdS72BW12+l1z
rcqVcXrW8vFlBnQkniIs9nhpzjvq6UUJBOO7VkKonT9khvEwg1OLXqct9+m/i64y
OrZ14A7JqZvhJ2m6MlRPVLx8XkgaaVzv5+BRPqEJMLNxDO+4Da9TchHJqNjSqaUg
KsiKt3Dnpd6nm5vA28Vq4zY6V//uJQGbJbZ1c2LHAtCqhwS6rpzlajWSStZZ6h2I
ifRdmTmNfg7BYb2R1Tr/9tw1xUj69yvoEj/K/fwxVh5Z6W3a7Yl2pSOV6uDMfO53
aYHMVM7+hL3qcFYNpZxrLNF/QK7OtGbOSbjuT0Wb5XoX/eJsYX9xRj3gI84mZGXd
Aev8BSLCqCDsBCTi74f37rZcCxrMFK5mhHNwWEeHV7pJ8iMt61Tx6fOK2lImkGB3
EIqvQ5M1jffn2R6st+2rLjIjrL3Tv7D3MO2PPn5s94DLknG2CCw0hlnUfeUnHn+o
a22JuAZIghE1v6ofmFHg2gvzLbMvrxI3SWoLoyincQnle/SwmPdOWo6ejTiJKyLa
fNwHMsdZ6G9MD6WrbhVMrcQXokPLdNTwescJ21SwNbNPOuZu886bkHWNiQskHJiV
kanRNZ1E6kJBvD+viBp6cQgK9fV5BJ7e4D/mDIiPEk/hnRifTaPf4wXtV+JTXb0P
oCT8N7NofWvzbmOJxo3jXASmd4RdnHv8ORbYL5kDuP0p6m23si1hEEziLxi6TItG
kWQTAafdQa+spBjlB2BJePvFTR1jPban9OnRbEGWDDkSl733uOOzJisADouEfDWF
5F8Vc4WQ7Dqr5/HWZe8EKrleod+2hWcwEViS2VUb/u/7mQHSgUpQbfyUNGEGj7a0
lqpsPBcJpqAc9Tu2aHHXL12QVQmwgPLO2kF3uPOeWZuBGL/Op6lbMY1DWK4BIRK2
9ujVpIxc2ZWsuHJUmzbdKNTrIh9jxtY5GW7M2T6BDcwoOF0sGnb+/WOIs2uMUdWD
2OFH10t5Qvfa2mL7sKkqIPPcGZoQMWYiyp6npv6EzPEvJr36IJiUFwDjPziYmags
DEoDa2QGUUT1ZTMXCK5MaGB8VEQ+9VyL4rtoKlDcs4fFus/p0BQqin72V2sk4KQ+
yAbkZu37uGxrmDuQQc/ClgTK3i4tPEvWzLJxu0gEnpSNp8vKo7PQV0Uhh/QJQ83/
l3kJVnqzzJAZHw4SmvPGkxl4putRrQ3HSK1p+uD6emsDGqvPql7VPclWI695RNBD
PdsteO/5mC59NJm1L6AUIpWfUuFMxiOS9w9aIXb7cpb4MfLLaacjjTtMNV6dwm70
oXU84OG7XbQA5PS9762a0zZiI3f9MvjAb4ZBNOSDFr9kYUc7gvRTI9zH6wO8kmSo
LmQIYygeVO2Hf9mEozI25cbgmdPNsam3SqN/zwryot5MvJBsqzq0EKf4tMSpRVd8
TXxx0vjCWsR0gbb4iBbzRELMIxulXnBDeN0OsAWGyMlgGcOC7VigiJfszMesIae4
FGSgaXSU85arVX866G3R0AxMd9XGqWBt282qtQXLAVIXvXTF6n/W5L7JZs8Xec3l
X6tjR5qdvkCAoxp/LSDcpgan0SDDjv1eYCk+K/uxhiU6Cfxx8hw8ouYZV3oxsAAU
bl/zkynDOOD+2Sb6sjdrPGOjqFU6qyUO75/0El5PbvybgaI5JDB8DrUoO/4WHOaP
N+ibGzUAn2OjcvG64Gf9GBSJ3qCjgFN/X3Yh4fG+l1pjZDAvf4q5oPb7AsDzX69e
eR8tA6Gj1l82FuJntYZCizNtZ2dq3H5/h1bYXooJBbpeijfpCX4JromTSdr664FF
L1PRe7w41uj6AH3kYCRy6rvM1p9lw7LBNOC0rCQiBh/wL0RgwWNPmf37dGsokQJm
aUGreu6GlBgZS8XXmW5CyXKfQMZWjvm3ntW/26F65dqftI3CQFxiiENphadodb9b
OFS+ATRxLPTZn3VcavrJAUMvqGqtyBPYPhDVQhMYenlLdVlenyS1krbMkDDKpcu2
QWzcOIGGJgi/+0JpwoRANoAi5FRIuj/36bKoRJSyB6rCvjSxMtOd4h7vtyxSQOgA
wrhapcbhahEBfO0BNgsGx/k+XNPIzcx36xU+SaIN/Cybttie+sZqKPh1jXGjCT4o
31Aova8n9X4VPq1AVZL1GjSyZ18D78UHhDT9gJ2CS1kPHH8jYvpsiA1/moyruRDI
qQPSMN/FbqZTMCkZoYza56pKpqQSGXlp0EvTfE6pzPHfUqOLknNRFBW4oQa2zdP/
RdgdeMZKjfs2LkkZWp4xTEhzZg4eXTaIdQjb3XOvMTEg8JVU0zaAcCqpIioemskd
NwJ/u1Sgl+tIavxT9rOOToQkKBnyGMn6Cl2N6/uq2V1L879IKb5piMqcKJegteQn
LkvWcQLBvQtnS6j+9dFl0c+P1d9AwU3crtNEQZQOBJudcdIB0VZEmHwaAwxd+qe0
4XBoph7GxWhc/ZrSuPvIuJHxPwkJBPrZinqmfiHhPOVeVTcynaDmzqxoldfnBSte
LuhNFaPSe0kJO7+/vVMsFjukZkeTLfzOWVHok08uFv2Tj8nh31NdrzLhwDKumDwq
dO3GaWUwJhj/mDsBRdeV70mukVt8Eal6s7Vin05X/eWFxaR1l8vASqD6FXKyHBoX
Zxkxdxh1wMDPPqtZYxQ19woRvS2D3lKKlsTuhsznXQbFRi7uB13WfQX8+v/VaQ0K
61tg1XDj3BW/VgDN+nldZiB7TlirHJ7jjgymM54uSVapen7yZaoh8GT73TCbLe4Z
6s8RPW6LpPkQWVkLqZj17UpT3mpY1fShsBGNElBfBKsd/1cfzFdK2xpxu47Snc/z
jATs0JcmK7oFbd3dkcvnXukx0FSlD+bIsKpew1f5L6BtWyxtyk1fWYyaeu/owIAZ
IYtM9V2MjM240ufY8tLfd96rqFtwvnQCb3lFD1MkyiEd3y3Xx/reQLtM9J5fMwxN
AgyQDDdy2jzPt7ZScdBPQ5s+qtsLzH/MLPzav/LCIpItsPjeiD6wMbmKfuMQdXaJ
z+Q1xU+rH85ue9ryQoJrc9tLYfy31CfrLFTBe5l8tdvNbNg/eCd+Y+0/HCmHfaxP
04Riyihmy6aweLvQ8DcSHbIvrBJFBGfckifHxh7QeywQy8ZfN5Q0shGgJijDsYzl
oqecWpPTl9A0CZE01E+3l6c8RvOV9KV+j7pAt73R9hkNX5qbJ3xbLpeZ4UsETdq+
Oy90kEyQy2aifr2mjBHZoXm1I12J5HBzV8D+3Buj3/FLqUO86Jlkj5iACM5AHMKA
swwzTyyFBgSaniFQDQYmq6a03s/t+wmS8Z6gaAwbA9oEe/roKfmj3tujWNxgGhSZ
gGTGzlNmHcSFsfEghivqyGTqS0eM7zKU9VpM71cIBdn0kTPMYo96TzG/TlRwqf4c
SMYgSQ2+CWnX/SvMaDxyrkzgWMyP3NGXAzbrVQ6eWt8ks/Makjf8V/7Kls0wN8Lb
nBRiX7TFFelqFgSELZzFq7DLKhWd4z+Wg5wwrd+F0aSdzonIS+DF528JGW8qpyA/
ceALFil2AG4Y9M79wc/5f3o0w/DOo4c/tSAIPhZgXT0fYDf5FxEhJLCZgl0yiqyQ
hu1ZVys8qNZQU+7GFzYCkrsNqJ6C0KLjXfDIdhWqOoomzdnVjjGLcf9HUUKdwgm8
glUsA6dpJ8GcgvUN1nWRlCpll9Axbbh3Y05qTMCiRLxNOCVLRnb61YSxKS19IPl3
2MDRHXadLY4w3mIOPI9zB7CKR3haY05SvMOtRULXj0tD5U/m9TDbmHHjBgas1Ltl
SygrHBYeCnsjkdVr2VnLbS3w5tn5Izw9BwtwLdzg5jOWA+/Z7eAvJgsNs8JORbPy
WRKpNeuSvaZPCPfX76CjjNZaorCXvP7Q7whYdoSFQN1UCpLbZgcuJ3rcx6AdExc7
dMjquU7Q9+1Hi8RedfOXtl51gnrqKeB2Feum5AFb85NOstsk962TW0Yu8++LgSd9
kfuMWOftijV89CvMcCEGMiSm04CznsbqGt1y3ZeqYiDgDfoG2N5ruvycsRQcv/bf
SG5IW9AZE8i45/TAAiGN+OyFMGRlFzG2SPLtMBwYzUWS4QBx6OJpNC1CynG4wIUh
w9tipLASB2myx1FUNE0z5Tn0OYJvdDvyrXROQJwQvrwUoOdv04giHf/XFKDmdmpA
fsuq3cVhuuQCXn6rE/8uJfIMuK/tQTw6ETTNkBGzrQie31rkChCNZmNITAD5M8z4
A4TCZfy/LIjYJ4UwhLnImEY3cpC4x1/PJIvSZS8QH0NWuA9TPB/+A9mRWEcA0zJ8
QoRvlHlb+Ma/gMuF89UDnI/amVpPKIKvW0BeTVsVjJ4m8Gms3oKevngTUaUpf6qD
yFnwxB+BiUq0Yi63/bNYhn7Nt63REgV1ATvUhxOHMDWCG7GdVnB6lrsqkjEF/SJW
TqgzA4yYfoOGI8UXV5rPcmd6g9bXgNc1+zOBD43Um+FRvVblWaaz2gZAEudhktPE
T32UyLMAIGk0PihWP8ByVTpiUuvIcqyXGJB0G9bNXYyzlMWv02iNXsVXSAtCMdIF
huhjqgrnmrGGZnqyReR538T3wzsGRYSFjUTH/7j5hG0RYN2lBJp3ghJT9QPw2yjK
16CDRVhLgSXQ888W+uwygAUcIUmADoor02Qt63XdEUGZl+OcW40zuY+vJYKNm5Up
QAG9Id3/LYra2R5u5wMom6rlwfC6K0wk+L2KbhAlV3crZC3S8ORPkYSFMnf9yRN8
IWBu2qxFK1p6VLP+F9jgUcSl4lyylJycyWsLEE6cxdFZTeYv1E8U/w8HliXVQuZe
DlvHssrqofXT3jCmPHwBr1upUIjxVytE5kAVE8oAH/xY1pN2PjU0gNIHQgjDefhs
lty1JLhUBbSiNiuA+AQ1tkZ+dFR0xNJbOdMF3rZkgyAwhnaxZ2W4yj+5zKTF8JGt
R7swens2v8wmcLa8meE9K/COWStq6PMi8En66QXmsX2YBH2kL+JiPdzlF14jn8MB
V+v7h8TsXIio6+DiLVvLs2rsJ0kCxtk9YV6IYZH6l1oJ3lOjkWoxxWKkvNSEj/W+
Q35XS+5uNMbeDJ/fOBQJblFDW1V/C/J6f26+4KGGzujOE14wLgAMWNvaZnhmw1Nn
sfaDnNZmWtOPGXeuIUnphLjxIYXkXivvoEw1lI1CV3fDxaIA5UnmQedf8KsqA4Lb
7LQsoqwwOgv0Fml/XblYGR9ZPvs+VZOiO7WYZOzN/I/d8tsDXgZ6P89DLf9EYq5p
YFJcInQnPeM7Z/+l8208PtnDN7BwXQ/EMJ2duNaiZN/l3OT9IMZqf4QMJFxJcOWV
Geo7Rnwi4mgMIQ1lmAt7ldeqPAFkcEeAbYzwA9LUY0nAxC719bh8/pibTMUoFdH3
S6F4nySczBn2FG8/I1KPPvrkeZvXkWEmFZrcTgDwDU6jNBIqcrONhi1KhBdmlNHp
66YUvPXPkNPnQsZ9QtOGWH4GWr1ITIIN897seeenkxoOIRYP0IMg0NnUf6Drg5yQ
F5hwVrzE8ZVs602XE+k+hPmbz6GCm00YP+msD+y6cBvQdRbYfBd7WSMt5oo0sJaa
F7FMrOT4UGMKp+ug/VxVWlov8PXVrA2MVGBkGoJ0sA5/8DCcE0skqqQtNBGSOogh
uYG3LxZJU9yw53IIc/m4Tjwol26fTrBvte0gOal2Qb6l/bTyD00/VLa1edJtrZ1E
fNsXbmSrer88G0Av/UzDgjIweurhmWR3vyoPKqw0KZhWJW9ZSirafQNhq2Cy5xja
94cN4HjJL49NEPF5XDZtJRa9Lp52cwBQ59fZ3GMmFP48uC1NTJ0yzJkhXi0tyfGU
TPHz6OafwT2aC7YKYVe1HDBsbPCY5R+2U8RiXDh0/mNRo8KZD/MT24XF4Oz0rjo4
RXjtMJcMduaA83qKhqgW84+NuMEsnXmIsEClgtkxr1T/9YdOrNL3EzQFPHDq0Tyw
Nkg09rZtZnCw5zsMiKFFggMT3h8l1IZpPeXM5O0YpvssjOJEokTdNj70gCyO6IVh
SibGuvkvC6kvC0LlCTeaEPXOPrPELdMIBgHDm7L496dkWNZbgd7A60Zm3Ds3LcZ2
Psgbs0dX1eqAKtlEvrUOD9KMCL7CTQIiAZ54yg2Ft9VwoZE1h2r1EqOGNrvKAlhT
4+Ypo9WsXQi6oGSP7x9ITQV/BMr/3fCwpJle7e7wiv3c8Hz5p9AX1jmAjx3rfn0h
DvM/rTdaXsPcwXye7jGlgxydHuLLSii2MDDBt2MQyt2hqrdeZWAfUoO6KymRZ7js
fXE/WWWnLMvSiQNXFbTktx2NWTG3NJgXiv0A8Yb5Q4vulUxIgrWK1paxsVGrzXbN
Bu9nioT5W+tUqNlOHGA0+AAQ0ZGmJPslht3P10Zyr86u8oyZJubyCNmKV9+7EbFJ
CxivmIBFdI6P88VfMidvfyN5AOZMCm2egul6AJX9/oaItL6DRZDInpLHKG12PKMA
LiaJReMJA+eWTMajw1EUzJJYH2ciy6lj9VzdeA0Ch6ELqOEcTmm4SA23gQhLD+C2
MHAcqgNscYtr1cfc0A9PoMZtex+SG70w52A1maXwD/uoIFZR+91gMkm/qdRv6jI4
JKXlmOGBu4sTAf2qKZ09h7EGKlnoZ3FAhnUBOSdagHYr6cl3FJfCVSt+LxvGnLvN
XK4o+dKF+7dTRQbC3Nr9tON217hPIcFbDH16UGxXNGP0Yzr79kHc5YNNxeRy7TbE
cV4jyvSvkVr1a51vQI/GVjHaU8oY62vi4j6uLrSrg9wcxozxbxeWtGK5cSFeTQMU
l76rPO/TLf0/AywvfOPFxHy88vcxjVPunz2GJvbdGyrzxAsPSv0pj5JV/96GeuTh
lmDfurU1szgaTy9nilrZOpwiLhLWBK96U9bSAQoB+3YwqjUus6YyW++WW2wpb+93
pRfnwKrFys1Lwac+Xgls1ukcFPhQU6Kd3+68YwsP/A8nHv0g3mWFW84w7GfQHp+A
M956JPxciwUQL8Kyh10QZa8XY5dn8lkyNGsaVMeLSeRbjib8dBCcI05Y73aQ3+uU
a51CbKqr+Z6XyhroeG6POUIZYFfyWLhJchKGYgxFazICPBZr9n6cAbJtNpXCFKmJ
kuh6uQGe7PzI3OJnqm9i4Uhy1sZDi6YYBzxjgYbLKYp2z1SO60M+CuoXy38bSvl5
NeK8lEFSZIKrmpgCfbiK7qawH7apBestQMcYIrC1ReT6Xpkc4Fg7nUjxExMS30hP
gwRRvak6d5MGa3d4vidHpy2cgKJImkLSEHc6vw5f87shRvU/LW155CNz/vfHuytq
I/KlTbBUiYumYk25j9by2Bww87nXDSqu79NkK6eEidZggEcrBM74jUEdx6Zno+YB
UmkXBF/QYKeYlrlbDyX8CH7Om4xSD8CMCjMF9G79edIeNVGWPRdaBxMO5Vfv+VBV
+Kwdp9eu9am7P4nfbgbyfqRvQ34X2FiluDRUaLjEPMmfqrs96rv3HsJZvolzk7dH
EzpoJr41xgfBkCS8cE4Mksj/CDwXgc8lBSkUZZjvuMLwskuFPlbPVsJjP3kdf1R2
+kJGXCMLozw2FT2oxq4YhxOPNEFJ2B5RISPBXk+BCnw/KDR+BYMVCM/tRPbIMs1G
D5dkUbKG6jWuvG6YDjm8KE2LbhWzQyF07drCOhv53hnku5X3SNaZlzzTku1yVWVX
RZDCiWCCTvi39ajk72FxyAQHQnGYQH/CVnV8IowSL9ERt80NcjtzL+KmM0ul6Ett
4Ni2jVPLuBbsulv7b3QD2s0Ik41U0S8PNUKcuphcDOOCM6SJ8xc8rV8Nnt+2l+xE
GtTIRfC9tIkL6qos1uvkSi9rhzgL03ebq61tPhqYrExz2/QQq9PHvAXI7WiTSZo4
EXf5G441hQXjGqLhlmKsdMbPVQGE4V3ZP4OltBzO9Vxgr4ZE/yqHCvVp/4SMicmo
2RiTwQHTJfn2tA9qeuUKaeJCucEi7GwERYp8mfPvruAV7AQP5A+Vyfsws2yahWJI
g4E89hUMhvfe5GTtymDtvusAFxGMv+6tAnMMCCgLGKADRJzTecMFPKqP3ch/Nhot
XNRvswZy0EmCEK+wrcp1KO6ol1Hy1Zp3/mkDOAE1liJ41Jq+lhX3RE3tzDrIAHf0
sWBn9WsJLXQT2On0QLKB9rBr0YrWg9xtb30sHMdetQiXk7eTtr+zUH4h3jYa0fB9
+vvKRC2x0pv8NsIR6DJRNCZ22nL9b+iOyx9ZtOzw7HmRydvy2mcBhac3yUTNmLj0
XjR3iSSEKxgMY0xDPHq/5aTKU1pGF09lCPso3Y6meZ3vjNtgv1Om+uF3WMeXZewk
PQ79JyTsBQDrlgQo1NJBJpX+1d3W5GWCVUJdcc5U6MCkGd6ZitF9x7TXrvDxa96m
J0P/5rkAyu4Vt65F6woyNMH1NkuxRIc7nvkQo7EMqgOvd7wOyifoCbqtrjImtiKv
5smovs3GyyvjAzT/C31cZb2VNusYLqKdKx1I3hcFRSyMr80hChZU5UNlLyQVS/ig
xgAw0h+KOTLqIkUNhtrQheIo7zGsvFtW4g4uZw9gwPWfzw1JrAImBFTN31gP2fm+
ZduueQuLa/xr6L4oDiUC+UUKo732HLJdsfTzMPK9q40TZjoRC5Fle5z5w6SxbU7/
555L4gnG/qJaBl5G5NnXs7QK1TNYrbqZl+fNF6hW36kjgAeQ7JnhzeXGV8jOL7cl
K9tqChLtkTIytOwlwu2VZsjGAuke5/SL8sZw+pBrE1wNdW2VPqnQ3FbfGlsHXmln
lBqfeajmbhiDz9Y0u3InPwKFoFPGv35ANX4W09iExKYaQLSZdg8X2lg1gc+cXxwL
0vxeB9CBx3m0Iyu/VbiAxIM/oD3lF+tWjXWFFnqgTk6gEuUREyEscdVsPjFOfolQ
ogAQQHh7NC80bzyb+Np6IJZ4bYzTdBUe69xXti6iD/wWfe/DIRFBy79poeDzcAoy
cGYIzTKjKLWuu94ujsnuE8tfx9nmZnem1IqAnEqvcVaCLIkNSfBHt7TxdBzgKfDC
Po9K52zqMvTNw9lDKdbffUO53gEu1mDthDHydeyfsviMyoTbD23znoS2dUgjfkZH
fS5y0v1E4lLRdTofgaGZswmptVQn8DAZv7/uC9iGzu1rhywgtzMLRjFV6E0TWHWw
xIhya1cfM0GZLgKDfNVcjkuepdNzF1Y/iESZlYXok2g7euvMOqbAvMgg2R54/ZLx
wB7JecsnEs+teSfa1ls/m8N4z6NuSPF9SZnw7lItKWYNRFlf9yYDHTvilwvPvRim
P8qqN09GxZe0Gwoji+wZpmP8utUVfULgIkA5LMTodzafp3xBCMWzJnqevYQ2unTm
g493NWzTOB66ch+NGN25opUFPn6F1obrRwAHgoHqQ/9q6czjfSrSZvtZ59AUHeiw
qOO+A8nlAFKqVKAyJAmxz1y0IRb4hqVOOUztlW0sZlCI3y0+yXzOnyS7V5+ijrXI
Bs4uS254MGroB7Ft3nJ0WClpY0va/Tn2VB3vHQmx3wb5TbkaIZ9O7KYxd3olgsQ/
L8izTzjiGdXDs/AAYBlW3YfdKKETgqDhFHN4+1IS7oC70uFBIWYuGEEDzsreNDgY
18CDs1WLzVOIWVqTBbO8ZdMpq2hj3KFRhK5x/iyhOoVtZND1wtpXjescTBBWhiZB
oef8zuKraCmZJLatu+JnpczpOS3JhDgDVC50qTSaPSuv8UJL9rtGi/Zd++gq3EzL
CKIUW2NuGz58uvIcU5SbJjlj8JIC3X+dfCJY1kmFrGq75M1lCqynrcocnn480Ov0
dVkJvEifhUP5brvsOpnKEPYImUemWPgmM8Ank2V1KbDnhNF/VsasNptBXqej07L9
RWzP1V3vs5Txyo0nv/PBEM6flqIkX+C3vd2gm3B/FduQwa1hc6KejPlBEq5/dNIc
dpfUpjR8X+dYs7CU46/P3mIUzFKBCl/yC46afRuoFASquuC4uEvGPHnpGRE21VNo
cMtBQ9Y6AO6HTT+44A6qnr1uzouIF6IR0FtT6jufsO0RyUUqVRFbDWFdoVXNqyD3
V9sb2WdEW19HUUci1wLCrT4/tVLQysusTY+JgrinuQ3lO06b5QTeCPyzNKBgf2ry
H+aJuTkuEISc+PqpsFPKWNTaID/M+N9GcPQchl4RlkWwYxs9pBL4N/jU4B44uqlq
mQpJB8HSaYw2MXJnZJF9SSimPplpBfAZr/G3JrCN9ipdB8TmLpbWdrQcmAW8PGCz
4GtZbYcswnePzaANkCJbxTmwyJN/q97BmtVH/8SvuARZNJb6jz8bSz7TJKQgst+y
RTG20w+X6FbpRB4LH6tXTQkjOH93iXW5YXajmvGR9KOeY1/DVUuWDNr62Ay1GfAj
jk8dxDdab6q4NHcGE/TLFmu4yVTirPFuIHCLQXTjgiw20aygK8Dn3RVcbcfyM4Wg
5bfUbMvbRDbYJRqXqf2T41nn7axEUmhAcGGX3sIleMP9tJ3LWhXnXz9PV+Hyz6jp
+eQm3OIz+PKgt0NUtkaZXcXx86kszW/QNdyd7vwy+t0p9CztwfeehElVxPtT5QWs
9ClCwigPcS8WpdgMdsL4GtQCB/7P6oFWM5WMI9jeoZd1J6KaMcUtYS7Uzyz4CGCx
o/X12tw1jSbYiPtUFrLVwG9kK/Du22HjBHa2l+2XJRZDhAg2o9sFpflXvGwTmf5M
hFP6Y6Ujq0Pq44f8YSs7lgrAnZQLrzVZqZnoagQ+9Ba9t8yk+chONOUXd8WLKo/8
z1S6jiT7btPe0vIy5OjWIb7XHv80iUN5nP8FTbWI0VapzumZ0X8plKGj+HoMUn8U
e38eqCiQcybkcYAB+gwpUI4QJhoumYJjABxM5WqHArE9adKP2oKL2Dyu1LXF3BU/
+GKf9tNL2EWlu9LNYZW0A3orsBKZ0ltkgFFeGNuOC969MEXV2tsptwkPH6TLnZ3s
oaM4bIX+SmsSV/pI4fo7Cc8iloXKf94uGDHn8dLzuo1/mrdecskGdD850LqRvT/B
GSoyKe3uFdITVhEQMwEy9erN9tGx92w94Gxbb75NYHeSlv7C6tgBHvdq4gLMykhT
hIBzdJChEV6inP0AXsgSSu6JlWaLxb3AGiuiKauUOLIkSDzbdYnaWk1475j9vtkM
dxhJISioj4L/hlM+zfFW+QmME6Ld6RMRH+Vh8jdGmaW+tzt637V37cFoTmrfoLVY
44qrNoLPMA59rhbsdd8GEyFW6LCNUd8sbt/uj79cyjN8oH7fDMOfkv5ruefs+FpO
N6sQPOmzvMRF06IvxJRt/aAXosNCrtEyBKMTkY3ohQSQnyzs4Bd6d4TRgfQdTJC1
z28IrCopVzK1g2vFoT5DauD5OqMGdj/qouZ6V2buWCrZaw5df8inrQWEUFXGRjcs
ejlXkmpif/53srYqLm3hOA2OR3eCahPkVFdrgVdwphsuK/5orDyEkH7MMuwiDN5m
e9f2aV1qfww39OldH31WOVxblYmzKedPAD0syWopJhA+rJNw53Tb66Y47Wa+oxYh
AFghPE5m6sf0smMd/t0fKzDj8SxNOt26MYLVhxxZhMtR9AV/Q35SdTWydOKUjWQx
o9E878t5MZVSGo8bFYgu46OHsZSzgLT3qDQvqQC0mcZcnf70pheT1YO1Kw7eLlvN
4ptH5+yC+gVVDumVr/SUl/tpCtC2Sulbj4R3qO+OFSYYrt8Bbi9vyFfJjiIgYG+U
LlYyol7253VwT/3iaaH4+oWtI18BWXSqLu7BVTbU9HankpdrOeRWadg6jxp2c+r0
O5abs5l1SpT1CDa1B+JBMUo2maOahTkVnlepckPqg5kOYhO9wSbS/tnGCZPyAbsS
gw6H3+fJzfJ1HUfei0NRf1lYj3XvVnDVCAGfc/3CmxKbimTPlznRzKbOO1yS10uq
c1nAv7qX0FYjj1WDGL3mIlNrKhWqGdEtfluJ1A5FuyLY0VrkoXJF/hz8g6DFldrt
mFXDlKEnifZj/fFTjQ8lr+c2+9uEbMl1oLbiJ9FbqJwpdqv/2QPyWmljuc2KDX5m
SvXombR3IjF4V329GoKfEfdH+sshqj4+ZBN5/ZhKv1YFVP9BnRe6ngcdq5vDqnIK
gtr9oUDJUXVa8KYJE9wHn2JGRdo3wc9lK4CVQIf5iuRmUZJ3kYzNCjxymWwc0mE/
c78uP4PBli97Jq/GiylOYFv6m1pGQdwCv94wAs8idyRmEHxZObtetIGH/2WBbxy6
atE3DmQ9mFpY6pa26ZGJItxrUvU0JmJeq8Z/Y7voHS4rmv2aXjl1tWgRP3pyip2P
rPhTx+dYqZXVQl+11anFcnOsbhv3YKX5HhUqX+OKZ75dw7p0WauF/TxL6E4iuTjG
7eXcuR9c4k0LU2+JEgYCeLA7Bc7RIBAMnMnwa3zf8KtFzBotCzhObtoYrO2qp3iB
QkBixf9Osm6BgOZTAh9Mh6anRD1/ggYL2NmsXIPn0TGKExW1NzpE14b124fCM21w
rX5vz3l3peRyZGx4weBQ6UjHuWyqZRUaUuNSWUUvrnqwu85eaPia054dRTMjEae7
7fnPycLprPoYqgdqs4fobhF9T/Ft6a4HSNsiMi4ODmmBQXYSc/kuoYiGlZyaVnEA
hZUGNp2mEe7rF2SoBxpdnQIWtAIC6DS+l1c+B4f5xpXooOevcpJ8w9xOYSslncMk
YMSlEdoWBpfbO7d5/qt/veWrPBsTsQ0LHSu81GuXJhc5jgeW0Pw6Idy7U4qbMhnf
dEW0/1/yZIqGZodgJAJYAR2pB1ymjNtPXIZ5JLBKmD+2hvlg24CMdJvU6V9pjFVu
LkRxu3hsNOoMic0XEbi1wniU9Acs+nvL/DnOilirG2FChoDAv0ICRikV+A0CbvKk
2FDz9oGYbsp9BAp6wRa5bd9LaFfqJHYtoI11cmZvQYUSKul7tn667UPUVgNV9+nu
lw3bYyAXj3PznmifKuFPF66blBA5FpCda+7VdhmWvrAfk39KTyCvftSkndsYrhVG
yJLPeaSMLB3fmfCznCjSWi9PeaetFP4uMVl1X7hBpy1i2ZDD9WbIbfo83O4lzbpI
M84v4jGOdK6NJ0kEm/3KimAKJFQdLIBPgX8enBlJXXxlg/5mev3cYR2upU8tonJv
A+fTWT6Ty+jLgi0Rqbt2u1GyAJrf5fAd28tjN2b4sMwxQMysMOQEnevIwzvq0X/A
ISIQC1d5Fk8KFpLJJsItuBpGiCCJT2MBB8a5oSCuIyuJhP+iMYed7njlaE2dAo4X
2Ub0jk4Zw8EvHm84Z4EWxnAOGOtUdolMIFrGGyiXG8CvLO1NMFbUFqwTZlm7Bz1D
u9kGXh6mHCA2IRm38WpqI/RVxJnF6uuG0FthzADqgOxT6rFyKh3Yo+fl4+MU87s8
nDcbOiFaFNlOT3lf1eRswT0SSpKVWxgG/OHMVgcdblHngYkbA11Wsfe9gxBRHShx
6Y+yPgcSy+AuZXlA0pcyKOg21npa1U6PEhhRG4XPOUgVWgjORQHNjvT8S1JFvsFN
H+C5/sGJaL29UKyK5TUy/hXQcoh6xkDirTbOD1bVDQlM3rbilLQhyhDaqlNY+LuO
EnfFrqn1fGKHTmvDEn2yQ7iV962C6Skw+oZC9ST2zzGHI2v1suRjOb34YRTggzUc
/s8DYrVqKEaqgT/wXuorR+CO71Anm//aWLNuYRPcdMHVmbr8Hwq0K57Gaet3+1xg
+i7/QIBWLR0w50fvDedMtwu53/sE7cKjg+gpkSBBvy6Hzjr5L1mvYEBRnddkYAvg
KGLnG7tLRZLG8Ef8UezfoXGVslHwEC5wrTaakjmkBVhZ41n/ybPuBOgz8NvRBv/2
0wFxGob198feObtO0KhADjseLlRZFULZvtK/FImjpEsa0+9RHe/9M2lzXUhkoPEC
02KE/Mf8a/iaKPSdJdplORs1V4Sv4DxgJj9bRX1fsoldT184Q8XnOL3VN8+GadWU
NJTiFTMeClB8YZZoXwNsoM2Lhi7c3JT479aeGjUT8EVFwti+30pcIugWWhNrqDxO
6RzUA4hUNC5VFq0XSD3sSkKiBpHroPLTMQ20USXHQFcmhNN0jFDOoP6akCYq2rrV
UQADhA4adqHhG48Ozv3bNXYmlhawHVTUN95oNdsAVvK5kB+jZFcv+WF6JTNgtpPb
fE5S0clxggyU86zBmS4qfda4K6W2QPWV2wF43YITafkJOQEqSMx7TOQpDfj5BGXO
vh5/ai9Xdgx5S3FdjCs01dIdnq480snvTfgqxpQ1IR9uzrl0ocr8LD942LX0sNgo
bef2x1qNpsXlfmQpDr/uQht+wXRvymdmLOWYBnVPBWaCjMsHYP8Demi+xZPfA0RL
/yZWtK4tfrFaQe3x0AajJeVqH1yut2YLd7viVCa2ov/n9wXOjCmUHB8xprzqYxST
kXFtBuvtqIZjF18Rnp8qkpyopmuQuxLbrIIzcJpSHAtQHbAeW3aRNVY4IEd1z6QD
lhv9M9gJ5x4hXZdqyWV/ZvKckJ5SvAwxX1RL5eeZKXq0jnvFFgU0Ym82yhLaQVXc
9HYeA+7QCEyM2FVwHQwoViZBxjByooDTqH5P7SDXLBoSGhvFB7NRNdnzVHMliMgy
HG98fWfx3s1LUdpgjyoKXcgfR9QRveJ86ziJl0hAIibaJl7EH/QEBrC4IWKsOpvi
h3JJpK+pKBNxBWDMPuA9cW+L2RLCBdF8XDcPGSJxXytK196i2uk7k3YJXEqz3/QI
Ae8kuBC/4MeNJj1arvWJe/lHbW0sFPIxPUn4CuBJqKbCISIyssXA6tVKu3ye9wL6
9MEZtGAJ7BM1uq0MAHsfZ3E/9/HZpnkTWsKUoYyubUHdh490YTxy+dzNIeT2BTTp
CvemB3yJuDmCTr84gBhLDqco3upduiofAeQyXnPdvOXmUb8s6sHZ2PdBlRw7rbfX
ET8DotNlMUi3nhl50uwromWygvkYiJqJWBAVeUeWaNb1OSQJrubgtH0WCNVPk7MG
8MEHOdZ8mDmqB/+wATEs0YWmH9+6Ayyqh7mUzp2OZCAb0e3FZ1oKE64OytZPxi5y
ozxKhJIlwIe2hcvAohoE3d/UA7L6jbkY6W6Z1CKF3gX1C6XKlP+DDSttHdcZveb6
z/O483tNCBS+o8daBeBdHSek2Agk1JqZO0pIK4/t1xeOb5UQPKQuiOkBTHVzTDhJ
xiN0sHdIEgycPgn/N8xpn0B7DhT9bvem3xtvb6035eMmOUACJT5vQhdmYbD8aJsF
QkGP5fBY3zerNdWq3lpwKuJ88NXTTONLiPu9+oNK1xS8p9/T13ZGnPwzt7beicwD
YBlAI7oHBzBB55ISYup65WSVDtwPZWF3B63RqiR3JSAluCHKlNws61I6u4JXFPmQ
8J+ik9LAlVgnscIaGfhnCMxRheOq2KyE/tPQC3Xu57o/8wRZw5dQm1i4Rxd5XT/o
VllxPPCDsIxcbr4cEYm5c5g7QoL1U8mKu8nWEg136Q1g93OgqJnFAm4HqGmtiPdW
+7uxUYnCmrs1uDT3dIOqXGfLy+0UpO3R/BdzsUTKhgyzL/DpUs7G6ALprrBJ9/fP
MSLxfP/NLq3hdMrLLvuQFO9OqvwZBYx8pg9BvCAOZUk+1dEk1uT2PLxnqtrOP1bc
GPObX/sR6Q6GArTmn/cactuv6Nl2uaPcEklngc/Rigsv9+aza10HZtR2TVws2TRD
VtcK8VLm8ZidZgNwON1BX4ZIOe4H2kAYistBR9s/ErIIu6NjzqE15KB03Xvuu2eL
Lrhb82iS3TDcQHczLPVSM26iQTKLKfol7n1jORjjZRVujgJ5iKb0HOMpJze9I/xT
UYykjpWs+T9Eu3OFBdYwBcKGZrV5ksvzjBislyh8tFkkS3B/66ISYZKxoW/gQsEs
1dtfotKmUyT7uQYRZF6uw6BNnqcFO7IxoZxwvxjQ+t5hPq1dttWkcmmiXK9WtVbg
4gDItBxMJKqvhcVQAzpnbsaFPPSdlnDLt7FyxiSNuT/t7FomJwRwWUxBB8vbLcZw
XMXm9yOqR/eLDac9j/CDKFiVwbi46OGSlezvbgvOS9bBbimNAr/giOA9amBFt6Mz
sSBbwlF8SW/74WvkcURfFlzkmVBMeZK5JJQECHOIL1EhS+UZxlSmArBevh1xxsBr
UCH/CVVNbh75KjUkfQobBD0zOCym5hzHhFTG89cooN+OCMAPoY44c3+O3Cn9h4rC
JYM+bmO6xJJ1Y9mixv9SdovMJdjv7a41ZC8EcbuMsDGUpIh8RgmBoGPjtHWgp12R
TYo1rvBsf9a2/grCiZzcsv9Vb+qdsFoY6CWoEdPyA1X14Ohf2hrLNKS6BRCIi6oY
oTTB+/meNJPcYnp3wpLktwzc0qL5T3rBFJMrgADLsHchs/6O28T2tS7T9Z7h6pNj
WVt2Jq2HlI6DtxsIMkmM8oFPoHGKQ6SZcsdZ+Nhz4Q/UZn4gP+rQvj1K5+z++b7l
jSzcUibRgEDYTAD1A3iqu0/ofU72JlcOcSc9G1vmBOtSghJ5Fmn0Q4TLXjnf1fdM
dsI06e7kT6QnCmrDWhZss5lPHakviz2zarnKIKerUtC63VchD+QlEy7Q/8pggtI6
H5H9lkHVjV6n+k42/5AdZoZW3NlvzqSv3JlrofGOZhQCCknNgaY9auYhCpnUwvy3
ltOLcEi20I7DljUjbIBm6zYdpigkjQu1HHRQDeOOuxIAYNZREg3UPArfsrt0mNVy
jNmDO4xysj+pGv2aYqaJlrep7sehv3TlUjoC6aoKJqDBkBKttuBAmfpImhO4S6ub
ybdNN5VCOQ4d3liFw4CB6J/g6m8xCeR7idJ2kLgTJLkv/G4y8FmXQGGGjARrZxzb
RnpWRjx0pbXYrtqU8vOdQm5Aa4leRLJXeNGFnNbwrl2by1CtCejThJQdWNaEAl76
mkD3S+JyYQztjxgeT/yh8hEkl+Jmk54+GSaEvTYJ3SR+KVuVp+3HWtnoHVulqqeJ
7OCxVC0uN/p9mqA5tIJdlZbhqnA4gSC1nd2kFa3E78eLQJNTNdOyxyODIFX2uRKM
wjMsvRuQZFxLz5Pwo3ImFRHYe+fG/BjAz0JO91/j2Kh8y6J/aHUrTNtk8F9wY9F0
1iTOik5+Oq7IUobfOYAqar6f+2rZxIc2OkqOhWY8KofgWnZJlnioEVc/7wbwfwWh
wpL8SgpK8Yn7fuKGXzrm28VZZ2m36ELg58zPFO/I2O0dkOHhywhXhowuKQT6QhLr
jAX5LzR9LqqNggwoESb3lJI8LaKBqZB4udT8km4M0el6NhtDDoxk8OdphK1h5z6N
3ldKGx2T5YtWj0JFJN9ll1Wy2ar7EGTDO7/YL4uCVICX7iLFMssebe40lngWa/KA
2xg83OQie8ehfL+WZIP4CoSnps5bbh3cokxZeVMW4/G13mcI+xc2R6iQk/9tFV6D
favNZ76KONCB0GHu0iYS0TbyjOhGBd3L/Jy4gypLQMCg8WpA34HIIAZ+BZyOYrO5
xr9kWtSHoML/FQNm3U5KLgcs4reUNaCSTqGMahRnqoGNBb7CnOPao69xZ6GDBL4/
aW0abTtd7DNECZb0WY7/87zX403rZtrrhN3BfE5UcSKcJhSos7xH1LNOtd3sVgQz
HMdtxCSKmR3mE3fv3s/A7fQHGAloSq4BfUSNaOgFqy605u4hwbKFLhXEBJz17Fvp
LNMk3VPR0rZehpauX0M5DAxIYnNRXBlfQVyuKF6Tugpm5bg4tCDa3w7vBc8sO9uR
gaYx3WSn8fuLDTNtUlOAWOsEcviMPrdNgIavJGtQqehzJwOacg+3PvcHUkbbwrIx
ynoDjpwfWElIStxlt2tFW+6CtffdfejCw6v+MY4Sc82/M97NsUdgqgA/K0q3heV1
l1baDI/RUe5BSqBh2pVfRfQo0joLPxjpNheD8902euCkJbE1vccp6gJOX+GqKqGz
Ihw1xx5fbsVjC2B9Jcmnki5VRU50abpVhln5LQS/aiGcJchlCJyOdZ9yFEpipC7B
WCEViEH5iMTuvZJUtrBXbd2t/2O8lPYz1PLZi60cHmqnESW/P/JAGYM2v37UQ2eX
DBcAh8i3cZICzCuNTLWImwouC819/tkB+VsqF+tF/fg6FEcY7WKN6ZIj5iEioa/v
YbOdmPTj6Gv21ryiK/1HyrnIi4DIM9OpqVPsqxpHHmKe1klP52mLpIHib/PijERX
ecIWKRB+afqwQlxjxWC1sbTbngugT6lspFhI/hREMmAQp2fx7/6ZWauzOGusYD1z
NyWuoxpj6hadRaDfl08/6UyMlVYyi5X4GIJOLDCzQt0OHOnEtOfBYWxPPKLXxbJm
dF7wek2ui0KqgjRwPC36uDw+iTvMlagTjdAiqN5i6vZPsrlh27lvzCdlehAGMlzS
yzmnsy3huB2nqf4UETOIQEjp/29z2OFGBkb6mw8Bdd2vSRrvKmWAk7gpMyhplSTT
UscibbgmzuLYWAdnemX4kxfG8yKPa96jWnKHKWBt4tMP0fDcpIAdAuKx7YkxzmS1
YKqrsDfv/KQVdTks8SJP6mhwU6sMf852npK5cZwIfq9k05zMjDiu787yOY4G+oEB
MThEuWlbwjGuZdWJZRKIdqAGoWz5gdO0JaERgyhs5Xm5B6WY7+oqaRSjXFPR5W2y
JDyNbQfKkZPpx++fGyekRx9AExrtcYVxUNl+tCtaCxjFmaYg7Ob9sEn3/zpaFZ/m
Q+cA67++Woe8kQcmu1TOovm1cCLliyKUdqs709zq6cdiRy5vT95W0dHXGZ8hHPTW
Ld+hrb1pq+0560RR5Uqb/G6racVC/Z/U0oGvDl9ClNJJs44wnwWHgh9ZY0onEPe1
jVvUOi9d/VFAR2vYjLpkdKbdyqO/ZPFd3xdISQR++a0e4OtMzBMQdEKCOybXYe/L
Tibzb/Ysqjs2S9ZlVMKVlUNCF620gToGrUijBZ9mWu4ez0R7BffxpFjg2/fjew9+
mSLBqsW5cmzcwbf4wysQ11YETPiSQeAFikQdB7ZruwVPx8FcNVRdPr0BwKGQogQw
u7WBPXEh8Gb3BZxCdWTpiCVIZmZvmqOLkCMP9enioUjhwUyjC39k5WnRLauV2bTb
lTAllRP87l46TKEOkkcLV2Cj9upJIZF66Dh1i8zqiONYOvfU1ntGRrgzyQ6BzQVR
y95b8aDzrwTy1ENcIPUF+Kaq+RyT64eW0w4nFkUXkoXMUkxJaTXflW4sa0/n8M7t
hrJ+dUSJjrI8mEpqHJYNKwMMtaEvv8tX6uV7Wr8CgAOkS/p+5soFfEagbrPMq+Ci
iL06qCD/a5jP+FuzKD0UV+Nc65L5Rn2Z71AiyMczJfUFhMUxOsl4Zk1/a6K33A91
oSMKIcdcWcwE9NRWcZdFI3c8kc7xzcahiQkm1HzbEgFf9USspiafKfwsKC5nbPH0
8A131D5IvzJ4EALZRuZKOCEezIcDZ85uwzUOL/LbvT7WR+vrsWxU0nRDezcbKnBa
zRdbZsjN8Av+cUmeBTktBfkttl0vRm/NFqj3lqBLlUffS+Wy6GFCKEtZDlWwdt9q
WxZatj0QWWfbdt+pbGO2z4K2CF+vndfWYUcYOVxLz1owHiQGbTLG25qZagCfCwCf
qBeHwQa4Rr9+1ZJS1/2rtz0rc2GYWIyI31y8Zn1qwrWo+Qxhkm+9ItjXNwnrluxX
0ky68gtV4ez6y/nFXf2A7LHBHvBIXAw05Pnad7E2YxJawgmh8LJMQF4GlJhiP0uX
bArgzOm3AoMIndwx9qr6o9CmuImj6mk63ODC39jy2oc3WUS5fL+Y+xUPk16RJhMd
EOGwCjz/HmOs3ig/VnE8oCLxCi5GcY0yYn5QGDLXyqQJh+E/smoptkCpfGDcrTj7
T3OG3D/6ob6gBCkYc0ZNnajG3dMpXy05tosJ+Y2W6ayYmgAV1iav/xJLOZS89wAL
5ifAe4Ovd9nnivAcx/fWi+44ErT+n2sY2CxcOOqIeQXbsExWm4qIV/9TaeLofXNe
NVnZxqP22Z6Tj+MeCctMjFIB4MK8AscuvWbgYa2xCFP0volGM8CKMtrhZMx2uZOm
DZHhZatvp16HtqIev6ofZjoEfT8rXeGMXFlpnZKqptStXwRK4ZGMMgVWhHYTLAap
nTSZ0cgq8mIDSD8mJrJAgb0UiynoN/4bA5JoMvFGKq+uDn4ANo5+Z4VxvqWfRZIs
3skgEZeXbTGHDk9oPP0t1nIwZDAMmhg/q3EuVh8qSe9pLO3nKl7YV38E3h5rzNaz
9F7b4+FnGlhArAkVJrCV/8DDGPRvAP4EA1CZHvn5ViGdAZJ5y5KjUcHJTPhbwKAp
rzT+scMAYYQPDXyqLQm2bZNo9GGomhspIy91Pw3VV/r60a5v6zRPxHeckz4Ux7dC
kDG8cTxHy7H5JAGIu5TR/l0XJMze5DH7I1bve17ulEwK6OGzTNCDGMP6W8kOy2BI
N4CYbTt7f+0RhPcD1T7xFz/C2o0FI8mI+lRlb8eRahREaUjJ9IGofL9Un2Jo2CQT
3TPuhIC9BOZmpS6uOLWXjmnPLslHuGqLil+arBlC7P3F82vAbELJ/ubp9MJaltLK
WHZ4u4nQIg4H2hSZDK4vbT7Hbn72ABC5sfoGiGZ8lVUm5gfzyKujkVmFhO8ZcPHG
j4JhNRIXhurm4g4ZqBYHRFdxQXlPN2L2fW/q4SkX2qKd3m+h+sl/DKf019s71rY7
UscMrAI05Gj/RW9mneQQxahwgpRWCMwu48BiykURRSo2ARgeI0x21bBdqgMHKE8x
0uaHKmbR+JLCwH4ORnI7mRSyLSpKGXNwGqtrrvX7UKB5hWIPUYG1/HxJqQd96+Yp
+gs58uszTywDik2i/SU0c1+WJjVVIAn+IK9a/IpnRs6+jmpjjd9SA4AGSUqvHd/+
BJek5osEmjPmQeioF10rnIqCd+A7z+V6fDGf+oEUrtXohmQ3Ekcmczjy+fRZt7rf
F/c5ZtpQD3G9HUlj1bpRomU0brga8AIjDJ4HlBy20SRQnCqx8hN7B931CuxdLSGA
3ZTLNeBlN1M9OiTLX64SZia7AC24NGuUxWCCKXp7HGHM/YX0CgwLJEHGlCdfSszF
V6dZxtpk7FEDvbvsQDxtkeNUG8SBD0WNS+ut4ATIP+C0SG55awItrrRZ2624QILj
mKU1UvUXBOdsV7IiwyRU9aBW+NiGJoah+z1eqi3MgibBFIOElFg9lgKRwS6kLORw
LvO5WRqL979ovIID1rRMlakBtaQmGM0czieDeLKY9RrrlabWCQc/U5MTNpRG/hF4
VqbRdwEhVe8XhiUSqL75j9gKf6oZFFNJqtqARMHAgiN5+hnphYwlSU6sH6nlomBG
VbEnQBHlXOB2VoO3mYrbHknwxQqsKjBD8Oa886+kxCFX0yYQbpd1zTfbJA9+cjkx
aP9rxDgd/fGcNKA8Nb9BlhzlitYbVoqQ5cxKNq1UxQfrB/ESllj6OSt4AAMPoXN5
srEMOOGUELliflyIXwqoiSCqMqId5t0Zhu+ayqkx9ziOlxw2b+epRJzsWNgbZ4L+
s8FiJtqCrIeUjNAVHw2IR6PiynRQu9zKft3ZvacIEgI1oZmzeqmcbUuHkLkYO5jk
OieHNekuEzemImFkYZPkUq+x1nsUhH8LGAB8Y7wbhFYEfLG38PX29YoEDsdbWBDC
jpruJ4XjIwVHIjLNAglapiP5/dDD1GVZozBJBSf5VuBEDlbXJb8eiXjM+Adju54l
rRRlLRGnKvkrSFJi96UO7+NII+/+Ni3fpl+v6htgtiMKpFdbHskV1Tv0FPsBUZfW
7o+dADUZ9PIpAacTK3dcguCRAqCbfQg8aaTTZHkuD3hp1jcWOK1b6aKrpK+ordbV
2zrZ2un8AJ99YpCZGfGC4f5E10hezlxEOt0Gm4NMKrCOIqJvnKUHy3yyhUEq6FGj
f/CrQCsl1Fznu+M6gTBuyHhqs8Y4DeTfhp0QYTRV3ni27Yoyuf5Ewe6ofOPESFYC
t+kRxMb1VY24m9DKHAttgT0tuqvjNnPBsEbeYPAAmkf6XSAZAInGusbWKFdULd/P
m6hIO5AZZ/zx3eEi3CmLDyWq1IwMmpsbGmVhi1EjdZKXobiHCEGMCymoOlLt7dFo
kEoT7Jz37Uqom6RSd0mDFLYivyPtu31+5v6oVVqR6eZsCuDGEVsaMyiFW9ViLkXw
bbHVXohPs/+9cuXEBheSOnYOVR+WN0jn5aPvx8F/Cs+E4GRKSdeBNwl1ZtShhwID
SCXtapugmjYEcY6Br8EAUTl+9CdMu9gF4uRnSwTXVZzlTcSSSpmiDm/t2dzk9B//
gV5B3f18V2cuMsiQU2236G38YjkNq7O3I5EVhkLgPRNE4slnurkYrZcCZp+FxawP
8yFiwlh5VoKiiDTs8vOMhuUYbYaBVqeOHlh9Rowpuon3zDYdSWY9dhgfJJL8POFA
pLoqJXjPiIhpLYqO6A/cBmlSAF4j3cWKrhxSeXWpYZthgvlrsrczWowBRoZaTEzo
Px20rfgBtCzKUSe+cigd8PwOzy72M5BcjzDSB3C1tESq9XpHe6md0Z1ELRaVDv+H
fAnUkco+HQBiB0UT3US1AIDB3Fe6aaH79wClCxVeUJqKHgNM/AMIKUBv9ir2Lnyb
tcceAl9vWj5FPi3XTQEwJxxF37attdajTKPqr/BRIyy87z/N/rdVAz0KZ8n0P/EB
Cvaun7Qx4gsazp29NiRyefM+wT8OhUu1quNSE5ct9cAuWayvDts4p/xkNhFh9r0Z
/W61njX3N8l7B5WnUL1EtETsWDp1NS1VINVzM9wlEDbGACMCWhi4wN8F+Q5kMqDy
sRh1ZdfLcTblRYkUB1nNAWZryO8+p0e/QKg84LBma7lp447RzdSIAjvIIasGYckf
J3QSFrZMGZc3T3pajKIvy+IE/z1uYTud4uytRsLGt//QzebN/M7lvCQKfQmkcYLw
tkDhWxYZ/F33ndTSFHEK6Ggeua/qVE5W/SGmn0eT73GvadMmp10re2Oe1zIq/juh
T93BxBQuopNbSvFeK7OxxbqHHZARtg0ttYn10l/CaA6aMh4Ss0ss9XexVWuWxDOc
R7xfj0HFQLWkmauRPNnI6AdVIUBmtujjZBVraaLAqdokmZSODKGfvubCXwbz7Nds
kyxPJGx1qC0++vwVKpsOSsj50130tb+Kt2I6aIhKUFBRr0Q6mfxfosRdmFWeliPd
LYf1NWlQZfLNs06/h1pwd11yx9J6j578ZsyzfDqaPOK6cNUaE16sLtu75KvS8G5W
YBSjgK/QFbhCh4WK3l2UFujLeq7/SdO/xUkcRIbYkX4MumHuGGqeFXSjWvtWRGwr
lHKYJcmJAKPNAHW6tUM1nhbcwl9SMWiWRAbBSEt3Z1KGj/7bnewqQssDxh49YnO1
cu/WoYY7e9wDtaUWe0D4Pds7H7sgksu59nshxi9RnWa4HIxVzOtdR6dOXZmaC/J7
F9v37/AGXj1WuqKBnBoqJuyFE4fa9qlgsdwjgOGmPna53VOwZtANRdCKOX2tTFYL
bibNoPiEfCV8Bt7S5eWN/kGJTUYl51ig04QSDHvs+u8BlreSgixlc9EgQe41gMmy
PvDq9YRVzI/qetSDlbTyOgYIRr/TD2hanyPYEjwwiSYRAkkMntguInaW6AcJGqJ4
M5s0WfYxWas/ISZUgEyQIGgzAQbwqAN38+2YhUI1fdMzzPQafOwcrHuzqjW5+aof
l7C55HRPlY2QueMdMn0m1sw9W+U9LA7Skhai3MWuaB+QxT3UkCnbLJrmsCjAgyYk
OT4jaE/rK46/sfs+vwoOesysn5nTpnyGd3oR0lPh2ddnAqr4ZVOu8hrMtHIelHuF
CGjcvvIbg9fy4YhEpwn5w05mc/Lm7ptE778NguchnhrBoKRzDvyT4OnDWR4zCrAG
9u2TSO50zx50UY+f/Tbq+thxyqi1CVYkvYarryFIk6DfP6KIC7uICOb4vSgEs5Lv
5A7psC8HkciBKHvp2psTcZD6XMvvjPRuEWVA2b2fTzi2HGzstC/uAbdpl2Fw4en1
daw45XbbgY/Fd/tnFBRY4D8KHI2CoB3mJWrUueVwucnQJuhl5jL/8IvGNmUzFtli
om6tNieEVLbnI4+/LWCLrlXNHIZqvn/lppZ+kqkVjJKx0miaveCiVvtScwizfyot
GJoq8YFSrLzY+r7NTGN61ALDrhOzCugr8nZ2KomvKcmHWDayD6MGnK7ZV4G46t0a
DXG9JP3h0QwCS6p28wblDm6ePR1b7VK6yfd7cI7PSYgRy2HHv6EzVWPTwfnbVAnG
QTGd5Xl4ZrLLuDJ/dZNXbqiBmPQpNx1udjIJMux4T1aAL2fynF9ukO3vCkT+7vcs
k2+3h+6pe85CncryEXFGTBSNeKeWvmZVyCiE9uupJiCR86+m1/wDLSb3Ji5ATE3x
i3YjJC7SSZrGF1haNScU0VdzzU1gi6tjBd857e2flRBlHF/77OjR9aPFa2Yorqsi
uBHXt7YFITtOKRg73DeG51cf8cz4Kob2LtoND6NdBEyvLm1eP9BcCv9TW2JKWB3D
uJOOjfM1f6YBQHnB+oW5FZxTXucDIyUNMCJj30K3nnx9sg5voL5J6ckE+uWThitt
m3rQfin/OLPBiC2jB11hgT73VDQqU3oIEef/s0Bvk/2AH3xY1oMzJ33R2yRrlD1I
R3FfP8uzgkfIYEVcQ4Rp0a3HRhkAHD+vmZBpR/OyM55eFyCW7MuCGAF/fqapRMn0
em8dLsWPt6LafKwFADeVFogDBoHdmrbj7xGv+8ZGvTqtyNPjT/0DRD3hEwcdufby
6PZKvN7CxOqbuwVVT4ljmplY9UsnlnL5pZEB12zHmBDrZDd6M4VDdb4ixXdhwu/I
QESoO9A++xW62oL+vkQCCoo9m7W2G+5bmpbpqjBNutCBa91mlvS4OeTrORXfVP83
xbXgQuMxhCUl0g9ZLAd1H2xVOXr5eFRw997ysL4CyAavcVm28GogyNZEQmmF8oVQ
gawToeopQSVHheArfHLlfF+yOEBrBJoIBVqftztK4/1bBLLpY085cpz0YnAnfkIq
gQEDcKDPssUSvg1lawFZzgj7HgEL34QTqnQIg2znoPt06yrddn2MXitJ0J5fc8oq
496fQGnOHeQ9w8Ms7OHV3av4onkRcfpqmZiP5IbfYkj68OhswG1B2w6oD6w5oQkN
nV7H01lKT1cTvnJZUIzz7946LRU3qzqCEW+7afvt1hGn1AyEQzGSuqUAbMGan3VM
OWCouGVtvmLbp39znqvSxweXhxhAIbfbpx8UrPWFR0UTYQkTPZDzLavs+RqGwnZU
BWpjneFGoVzNSECC6cgw/EjbZNp4BGqBZQZkQ3HjntrRldKJSeN3DOnxA+uWXVLe
j/2fza0uWsq5DG7Kh/anKKMofnlomWQZSHatHJNfSj5P+1qxOjgM3/rcePvYPcKe
oPPtZP4gU/PONXgZPtKVNBQErQ6YD4Q78aFo0PSh8u1DYpHFC+oq9IsrdMt/Gdzt
6lqW3JvZbx++ZGTwXrizLKIlkLiESIHy05jW5f8dY/SKsxtK5jw37ZsKwjJwTeN+
TKHRIEWVyw+o7h+Y2RPBhIR0nwRP/5A0nrMcWkhnaT0m+n5FLNtor3dFPib3+a3N
W7oK1kOGLhPXs5Z28xSvBaDTv6cr7kbQmf7kCGyotbgItsat7ehBJdzgl65hiX3U
lVumgo4+jSEEtpypJFl1mYb5P/4kR7shXXOO8+u93Un+6XsEYPrJy1YnD2fxDwK4
cI99KgcOkVAcAVuVF+Ej/METcG7pRDp658PqKV+6BGG7dGoodUZLDXBYenL4pANz
rVru2rpXlSv++wNwV34/x0MCjkLbFMiv/Kuhd7eCBf6GvEZ4gXKBXkqqF+aLr/Pf
DvE91k/mte+QTG8YDJVMTX8CqjJAle7l2wR8PZMpOTsFQZPPiWUauSTDbQqXeo3P
4rV5rOdpsPHwZtnm0GU8WusRRH6OIPOOCC5twDUOjxEEm1K06tx+94DDOehN/Ywk
+aoiVIaJ3XtMF8kxoJ1WXTU/vN7SY3d7ic/qbUvn0a875I4K4ezMX288diIuukty
+epe+VWoL0eZkJdBhQTYdpOhRK1DN4NO8e47lqNzlKWLXptqpGasJfuGljCl6pu1
BgPxViJR5oBsJqlBktzYxZuLhYYmmBHj+N5391LZZdiuJOrfwBWQpvwowDeRdY9k
9us5i5X0kbMNZy4EfWDZGy0T8GekJ3A/etX5sT5g/j4XQ7z4bx3eRlplSjnnlkuZ
141dWdgSfvUEKq+U701eMUv9dxx7IQbomiDZ8SbQhBLWWImMbU99+Et4pVMuz7Vg
wwowaiG/72a0gBBffCHcUPb1JciQMXfOdEAOSnbsM1Q/lp8KHgO7WIettOx+u0E4
AXzKe4sAgYKDkQz4b9myqHCO7QN7EiLbLxlv/1TdJeg/AHyxzFfFbhmSNjLsx1Cz
OPv5Vze7lCG19vWbVSe+YAVT4SEiu3M++R3SCZgLaTToK1cS5yO8peLWThVsxHIS
jPG2+mQV+9DAOkjSek5OLeId+vDqoeu3imSR8Lor5nF/V5ArjWJb58VCc/4Va5Iy
BXOFBPJ0RyG8wyqdjWf7dnQkgr6S9z/Zix1qyrVD25+C7hTH0ZHovdshzUgMlT4W
4cmbx5+q0WzVVJC3hGPPhwIawN3Jq0k244xBgbXAa+80yB6/U5sSX8VY3nhGMDfw
7cx+tBwMrpRKShfcjM7T040GiGfSYfn/pJa48/bXZYJVvNfF4qigigc2Y/yAX+eZ
WJGf3ZM2gL7heypceu3Za5XQTklaKHK586K/IdtYGCEE52TwsY173LVn19Pnfrrt
wXhJRBT0QZRXSzrFqYzh2Y/R5LA6RNxZfz09FJVknyN5fDYV/Rlh2CUsLI9kexIq
tmkhR92CRK8rmwvZXnpeJszkWhtDfpeGkoTHEmCYng/mlZTrag4+nUlQ93+zbXUb
JafFOvTLSCmbj/7+dYPMMz8ekqNyGRyQVDw3sYOAfQtctxTI89yVr7j4aImOV5YC
YzquvzjZ7fNr9k7GGJmTbpHOJYr196QOqbWT+xrvCgy3aKjAlk8ApfjP1MEnTXjB
Jkw4iJFGxDGuvhuD7mIR3vsVhnjUuB/6crtMk/Z68Cw6OBI+tGHzYikaWknlx7p9
ljCClfSLtXPftDcIcwYRU5xKynVD9dQgBy9FH0tee1A0Y7FJJ/RHvswELyIGBwCl
wOa34zfR3nzWXhoFvKaixTzDXXJIUI2NiE/WZkB6ehc27KvgcNLusnUMr8ei9RBn
JvMkyX25SP4Gd+IHQNupv1I+OWcrSyuYO4NnJx3HYsYwSS8wmWkO2eJRmk329GC0
GWhDBnvVpZf9+vLGOvWdJlcU2nE92zPYYr0W3hU28QNJWy8TlsTA4Qote+GK+xZo
na+vUocfJEMSZIGYd9vaI+pJwYNB4DAGFjZnqR7n+T/Ss3mec0r1Xs982QcnM+4O
wp+9HJtbrSL8Z84FPj5m9Y6XUoZ17JDKby+Sc7c9mNRanUkPtRjY/pZl8+HDQ4/+
Uv2JXkig6ILlTRXua7Hi+nrrNDwET3GI7uALSmhUExSf5+OiO2JqzUa76CXtx9et
w7J1+bElQbbGZZND3FykUVgSdr2qfUQ/fb8ni/aEF9+SkOpHoW1n2L2AJEcVTz2q
oBrKK9FeCQb2zd5RlrUVfmRYJzWOs0dOTEMm1VcxdhLjHDK0QsbWvrryknjvUE1c
xmE7x1eDcKzdPGXk3XtqfsL2acFCt8dRksqttZ+4gW7X+GnGc//gNtaY0O1hlp5E
E/06yYZM0fihYTHdOuzzFwBDZZziHzq6NqLLBY+enoAbgCzXtdJC8Va+uel5RJnR
xub6x+er9F7XKNUDKK86TfYRPeYyrRTnb2WrXijr8EFmNLDSROpG937pPFUtN5Yi
qEtGQriKLxLgwwwQK/fb+9EZaIk8u+TlT0/cf9KL+r5VwVpNVOIhCoQ20t1SYlDC
jV5+93SiKrSbSRW5SKxb0/I8YTHhS6oMPuyIJCmDK4esv9cDOG50DIKMQwdqtlpt
XFS0A9ev/c1e1hKwmcWrg6xY2elAlKsEYusu0KuoCMIp3p8WfTEGW0AJvArCtC2H
9BtgdtYHb5nz1UzA3Iw8Y8hShcjV6ooDiPIUNtzZk1RK5x9WtSPBJ75JbzHz8skR
QBaFRtn9gyDeXhkG4Qja6J7/2hvFVods/LGHB7y3TTm2EMMpkqvpgOkd2YiYhlaC
oh8IpyXa7aE+a+UToXydxvejFNr7o8aL0C8bTG4D9jM8AqFtIYU4xg/P32CxtH82
GLH/L2LTrP+nh3d8su9YTcIGdrK26EPYKQDeFZY5EQG4aoM1o9uLnqJQZzpWfOSa
+52lwmRCsyqAl+g0kEseGtYVMr/y7J+wSvagSMC/IkvkBWATWCd6lK7TKYay+mgW
7nl2SiiUV9sBmASyCpxzKqlj1VqPO8WdYxi9xoNc2dt3mPT2D71kOnBeOpHuF2ak
WZHPrWJZxIZ/Xbz34VSO8aJjB56DBy+RPNzjgc2sbP8V9lZ2pYniSqIzFBxBgGUw
rgDductEe3T8IogsJwaxw4apF35v5925nAB12MEKXSR2ax59RP1sj+yfZtpugTd3
zg+kBLXZ9q48BdPy33nEtbIHK50V43cZQ6k80Z4BUED4oLpX5c/Uf9ttZ6NgT5Hu
KKEj0XN8Vs/EZu164FdawVAvHbh289BksOiOTFKRmNSHBNce1jtaTJm1nnJAnw+R
Fxe4Rvk2Z2YxTYJv+TQM6R+TVPgvS5jD7z9xBKs0RQwmd3bDLcaw3jcRbDB08dMJ
WVlbnuSUcqEEbyfn+70FhwxGwTMJrSq2KIlZTLpHkHiMF1dcKpySJJOS83tCtr2m
voB8L7JiYQuQ5FExWOg2zOvZFnKzDVsACCWd8VqLnM2x9mLhnSLqOoNO9RfSxZvi
ZDZtd/DgrvLZqVqsIDA9ZpnUeG94qWjgHkN5uxOA/kBt0CZcllc3R3XGzSLhZ2HG
qx+9JBIISHnlIojLFO66UW5skIqKQ/Ue6BszA0OeOa3AZ9lBbbfdknSFEHUCHIqv
I3Yj6btqlbdzBEJjlEgaBlVCGusUnJfTnsouc+ojxU5QBQ9f1cQAMv7M0VB9pslB
lIhAul95P0Loyo19vM4iYrhtFt1CRKgD4mULJRWzW/okYs2tB8SD9HJ6GNP9NTH7
0fiRKi/0EZIuCzmBZLHwqI7Qi2HBwo0Cwndou7NbDzNAMSl6IwIkHdIGc8UDUVU3
EI51tFjL1TtHsvTTNQU6vK3DezJkg19qO+MeRSUwDtHJZ+NPJNzoS+bwawupG/k/
Iq6U8LkYID7ngi6H7Yuoilorhse3Gjh0A6uaZ8DS7NTaqsR8kWrp/5JzaoZgNBVR
DmytenrYVdxd2pdh3MRyCJ9VYbz7HoMmzYagY+CywF7pJoDzkhBChEIIk7CezXIz
+0NvTD1L2MjU91HR8tROEpfKNX/wKuDRfjD0IdWuiPxMe3sjK8F/xfNe7uwjUU8D
V6qF91FG1/k88Szh0p3ka09u/FwbrDBbsTYEn1/Wn/z1TOoHAJRQsglTk4/j4T/D
avYUe0MqD49geLA9fz1Y53Bv4pYCI/UEN8PyxISsTardhIByIP4XH46X9J1bvzet
A4mJzJe7gcMeF6FzJGPU0joVzaMR+irKd4dj3p/eXn2MqScQ4c7RREmsMt3Qv3H1
ax+P5z/UrvnEoEtdkfbxTQFvjA83nOM8i4SqcIH04EWNXduoz6KQ+lKQ/5tuzfV9
kTOd4rgyMmCNwGlcHq2cG0wbfbS/4JIdL1YQZIqbKLAngjUay3j7uOsaWiVdY5sy
B8Pj1of4PCS/emcLhuAC9ytjIj2a9uc/UxHgz/jo+jxM0ou8Qgd6pfz1udCF4UiI
5Q3SpDxwBFTrSW9jJd7llOOGmb4RoWKXGoL1ir/F0slAE4O8k8bQsVyf0YrmPffL
Av3UehofZbJ4MnCIhiQ8TX67CNb2gCVdAablnMAdU1REPFFeTwddJ9wdFaumUAyK
WFofusQ9hodh2dJm8xJGa9lrWBhne+wZ+PCUbHfh3+d5V/vTk2qnGjWMLH4tPIiS
RKr+Mc88OzX4Jn5FDpCWbfottpWgqBcSDSO06ZuOoZLOD5eCthqRLa1AdzPDudkw
l1Fn3yHWIrAt/bQmMV+kUnQ5TxIUaFSX6DqufGz1rDynMh+OA/RraJ7iYXqhKto8
GFPocS2Hf/5xo8dVxT/Qe++xAGh5loMPFVDr/CqGVTz3JESjp98CW9jr1b4HASRx
3NFRfNWLn+ftaCaw436UEDG32bjRJamaTt3ItRbzRQbve5IZSv6GhjHYiY8qRlpq
vAhDqI05Eags8aGhrfWaXP7fiiud23zA/yoPkl6uBqWiBs3uqaNTGD8WEG2c3p6h
yY4GWJOEibnLinA2QS3+Wet/DhUNYCbZLOqW4ndLLypnxMv4RBTVkIat11k07GRa
sSN4C4a38k4oVgtYEvwrqgzO2HF7SWMOsPAEeYdcFYptB517yGhtzpnR4obcJNRc
T/taqi8aNOJLCkAEzEuZ8ANnG4YHR8Z8fXczTAMGErfH6HY886ysQ3cg0A2NtCVP
Ye3+cK932RXN4Sk9l9LJB4qt5Vq86Vd3Ei706YvAdi+vQFdIw5HD6ehd/VuCh7Bu
HB/x7Q7szdp1mGHOtrTxVaxR77+caS/RuXz7/7uv+LwaEw90a0R3+2th5bEnvxLc
OfCKtoPjzWHdKBuv4Lb7r7CikAzGLQe0PghVLYiM2HcBmIlbbV/RdRAjo7X7umga
+olTDjWmQXs78xFH37xy9OOANn8qrC7A1M9ZbvuFnfW18BKYUUST1IS5VFCujFqf
nfRVXiFMbM4DL+qbU2FKS5O6LyO63cUyGmG2E2+zEqI2kOH+nj5lUKs7/pDXSWHl
osQm3MYEMdU0Xtq6ZkJHC7vNdLdDOD1LjBwcPTFAdY2jWCkrrEecnpN3wnI91NE9
HY2gFVhH9XgdsKx97p0AIZ33lChTcULTLFnHVMgSzakwGmEkJEyRw6oO425j4cHH
YL0K861YgM/VzrwGhOdi/gGzu6L8YeQY4m12nEcCtY5maWnYOudjFUB3rv3HOTbo
sYVMRw3h4gGt/Q4tQOn1dw3IRu42oo9Q44loHsYglQGTEGiq/UXcoEzRFAneCGxA
cTnkGWOZ0hSiGWIFS92t+nRh7O692C/beLpYibRAPhXRfWKha7v3ICAP4PxVjPn/
0BJamkFTy6xvBzF86Rpy9TYWqfacU4vula9RC1Tmx8gmKEB9nRaMWRenHuryjah0
qBlLVFpuLHUPHipGAVj+LJ9h8wsR6A1lj7z2Jrsq+yvM0qmeTul/NQXRtXOB2FRe
cSoEjnKRudMvxjMR3IEFn8jgyJM46ZsuONLO86yY9EpTVPnMqWpuBjTVhOGC4pks
DUEPOp0pYjLV65HdbIAGsM4L6J8ygFomcPSPhJ3Mm9TLC4Izs/v4I9XIYwj0xJ4V
ThXjXG+9l/zXpgPJC5v4Unccj5IRexfwDd7lEDh9O1YpBRGomRyC32Qll2jT5WPG
jcnu6InzubR4flioMallx9dZ59F52u2RgvRak/nLavOnO6ekG6FQPy1zVkXgJzKy
9Cfu/306oAj2KBGcnMl2Eq34rsceYmclZFucM57IYSfuysROfGWyhb91nn5p/Va8
vvIP1JVDXxImyk12nGp+DnG0cveZHB9+b+QVQm66Oif8J0Tfwt+rUjn8zNBwCJch
RBzDuu0LAVsnqCoDdgeAzOXa/h0zn4HW7lKrwfjD+J1dTc5pI02PZApQ31TSJYzr
B6R8BRhvXFDjJLGMx1lQ12GmN2mC9LfepZUMzYFkFvkM6ikNmgOnNxmdTAiJmN/+
OMxIjjcAXY3t8mhxc8/fbV8s0qHOvNq+kmVIB/Nft2IFeCA9qbW9kb2SkMeytUcX
9eB3aFLV77CyrwEkFfMsMnjzk7qftBjGGkT4InFHsA9yA96/CvzdWtLfyuF+KhjD
y3Ci9Dmk1lewa+VQi3sNzCVhygVhkBZZuz67Bgr5pElVpIBVQbj0BlmYxztQuOu9
b8YZ9YjXVMIsKiOneQLe91X+5aSPkcFX/oukLYqJK/77b+N7q74j7FZpMGTWTb7g
Y4uo2Ir3rnUi8jtrFEDd3mfKvaC8ArewMFu7w7g1flyyCBRSx4cgVDbmnQTbv09R
l5ARzQDFArHctgCtYJFzga4vcWVrkmuhzHP3uX6KNLpJFHXrozuwk6/4zvfHGB65
sU6m1qMf7k8RxDLtdZA+lt7Ea72dtzRv3bPLfYlVn8vNyldMLZ07z3G90JWxMZXP
6P7c1tEg3Rzr8WVUfLpt74udQ1vxE9BGboyjDSy6xuUTgh2if+UZ5jvldXAc6wpT
36g2O7pJrWONDHgkvZZVsj/gkJ2Htsk2d/o2DhSQbvVBlNzsCqFyb35pc6aOBB3E
5f+wzv3VAQsHETnFAwTvpk2mRMOzPCJgZHcLYGfY2M/FyeEmUHyCS/MgmsU7oi5+
Ot0n5C2Lg/Sqqs82cLNmrBm3mJXYaLWBxsBDmDNY/r5Tt/yZtuNz4ORN3lhBUSic
CaORdFQRYIHkopUQS1cV8SfaXsHEIxLWgtsxCgCmGjQubvoPnlBIeNuBxg4+j9tn
SkyZeYdi6HTDmYi08nCLtXLnBw9Lp6EtqePrt3jHeiXpKiUsWYblm3TFmmAszV+c
+HTkZLJVyGHRbWQCqRk+6Grf6pkA6/ygc0oTsXSp3oZUDXwsMAjUCQX9tNeVjmFG
o6VP71Osj9yyTSHu46Rbuk3v6OeT8/Cf+jB0SAw0kDyBNw5CN9/VWknY5AZTHLSd
NDfyFyKlDhnYmQYqh0ZbTWk3XaeK7lQQzLqhImgwN4uwy/zWpis2WY8IGganifd2
CXxZk6WfAcRQDPGLUSIRo02UxIm3AX+lZ9yGQ9d7Y2afXGkav8CcnlRTkZdqYHxs
EUsz/4et6a+Pkq2Xfk61Jl102fVRYKtzIvA+wBU3F+0V/pSq6RfQ+7TmWRh+rULW
ZN5avs/v27AWv4dALFwwudIhNsu+Snkdxd4Tj7izOq7sKvfrQhOnmxuwZ7KnfPKQ
aZ5VMMqjlZm3rje1inXBglOmufOyDXovPW+l0a949ReeLDz3jDpm0R+yYTD3jnTl
RdF2WUXeKB1g0sjgB2IksFiS4OGeEo1M0ATgoYxrtGzlemgqbDOACoa9fr5whhLr
QdTntcB0Brc15w1s9lBFiSuAcZMgbKs7eQ/C0KBQZXcUdjJMYVkf19wBFVB3czmQ
04HBjagXe2Atftr925BQENRuPOHx51mL9z33Vfm2bxS5NwknVvxXFR5k9Fg9ZJC2
TDAt9ym78DeH+L9m0h9fcsGBnu513+4IenFtc4HmuYRp4b19PgGHG8U74pq36Y1H
7J4Y8WqfStqlDjeRpkpN+CnPXo4oy21A2rvDcwbZ8OyKj+W8jguzMrtD68XD9CJp
2HJJxHLRoz9f4de+F1tQ6g8DmWNRCbB18gFQD/ffhrHfeU5P3YgwtvFyKFtCE5wx
/TnghblMhNGMEEjdMBIg/xGdNnawIa40cLDbyuTYXeUwkOvHrZBF0m7D4POynuFv
8zAxO4q1BDz9yl7PDm/yQ5LIl/sRvZUIJGs2aOrW/vum4GuAlUr1vtHe76eiKKsE
IBf+VcVpXx+NT5XpM4ugZqiBkTNTZDAnSYvoBcAOXcArWtxjz6oCopMadLGZA02j
JC4ZIcgGrApwMrErovQfr4TG301Zg4YfVtLrihMn0zkEPUDc3TSk5K6VXxivP+6U
9zqhTcfOM+sTdpIRLM56E4VRpKY0a1kglTmvARBCJ9AFzTgtmLBxr85Y+cEUd5B4
yrVebEJOdgc8PE4VTsQdWRsrY8cyPs3+tAFyo6CLRSJOLoTO6PscAOmuwf/QlGmE
PrZv3IVwzBMxlq81uZVuQP3B5YljIxBROikdeTt4C4nPcqMReKQ8BgEwScvnOFE+
kkTAQVGInLBJ+7o8BND9mnX6tA5q1dFHsbopwpMD3PaJEQWCuSckOo0QEXjs2xxD
/ZKPP8yNO3c980PqhSDphfG0FLm//q1pThFR0xslOhitBAu1NkoVJvA77dZgKFtD
EoA90nX36Xtia827L1TAL5U+6qUnjV9Vx4me2CFxWxyQVxixiPTA+VGh7s+j88Mb
Kf/tuvmLzcXdFoCg/djaVD48pjTRBRz/a8NZ8G9Pr+iY/PkMoHGr8+Y4qjoTf0aE
jkLEkU9YxINE9e7V+fHRazMPJnxDqViXg7tnk67r3rCUnHe1IKolUU0qyU77XPmn
YAZqB39JgpxFoh9PdnweeoMjBYKjwBvO6oxnm8yqNs/qwRo7ujhTSQKQESxKyMX1
plA6dyte1qLUQ9iju7mxtjVIujhKYzX43kMbRDCyIl8Zv3AinUnBXuFJL5Sy2Enm
apTZokJpZ+b9/S49ZgpAcrENgVBu+AHklbK3Z0bRzqn0eSANe/6Ll6Wmi3lr79yN
SAs0SiXBj0AsSdrLjCIOIGg6Scpx61wRZLofiLXZI5CG9tNxoczkFdV1gN4rG5IJ
2V3F98qT4idc4sK/tRf0ddZxK3ALosBBtubkV5y45XlSUanUBS2D7YKsDofGNwrt
qXoX4wj1lhPJo+9gslnNsTTQBVDjqF0+/0bJS09MaId1vwpPJ1rk2KfwRcGxAKlh
byWpDusuKPsZBbP6yYtUkHjvd9YQ2+SbPujFBbaUSFXf1SdbIyyKoTkE/+i7K0K0
hKUthOHSABlgAtzGOsj6YTxaSyaNMvVekTZ8w/tGE1HvKyDY46Rcbu6kHv/QNgHW
sFXrVP0M9vEZGnx1A48WXN1GrSaJ5r6cMV8KAHAv5mt2fIflE6GrmxhP1Zpg7xo6
YGo53hPKCFeqSJGp8TPj6mABVGV8p437XplV81jQX/0fGjCXgBWC+fTTLrNoj2gK
CCgzISHydYjPF8KRP8/Nfud4yRcmS+QkkgkymUdBDty8BhvNy3fm5EE4KmbmaIyL
qEQRfBd+Kc8R/F6fnGGexG8RX323R4rEzStUncwHTxNQ9q/d1POzskfzYmvbK8T9
wiWsAF3tc/k9GxZJIrReZvIA1jVSAvDSmKFK4qPTQKLo7bVpyG9sCRJVGFecr1u6
T3ClpK52zf2f864FWY8PJtBw48wCIUw7r8f6C0UEhrldGjr9Joib+W2nJ7vaP3+Y
lY2RViOpkxJOixw003GhMbukctXNi0Her7CmkWZlIxAMBiFG96DDfGLYSPgJGm1k
b32yHOnEgLgoTdgTScV/hTJY2O3e/pZH00ylpqQ90uNxo6CSOgVJI4RbSilN9OZg
PtWE9R/q2cEy5X0vOm619cOxtfrxYlV13ek/cZa6zZ6o9uoBKC0aBfFe8OOG/RNw
cv9C867CRfL/X1uZiKzxn37e8Gjya/VKgQue8Nuv7X6xUeY8H7cOZj4HbLRi1Bk+
bBsO3yE+JssJuR6euQwt9zIZOmFK3PH905uoy+rupKwXkZM3xO7IDgicUjoaSnD6
BOCnXRvez7pB5yYglCSM71RwAgS1MjStQxPER2wTAGx8zxZ9ofp+stxdJTazRiBc
+LfqxItE0kMO1kbuk2dTwiks3qolSKjEsCmZqQc9XNcpiRKdInyDu722wgWUHzYq
jzII7NgHrn9qY3CQ+mBvkoFqiMDY3iBFNonDa1LRmC+b01syyOEy2/mFKgMxVHh/
LE5DY+dk6l1VHRBOw8N9TG4BKfFAdG955P8Cte4GZ1N8HtPgp4ZXiwqVkolBOUNH
kmnq9HAcn5/2Cv1EhXfefByBBpzMVf9t54H/RjGzRPmvnAg0hqIURY9Ih10/z7yb
KYHTlPBJzgiX1+NOPaEbwi2GbTdeKjqezKD0TWEkxwCy9Q0NwrCEmsRn8asHtaTO
HMeVCzDRsMPwM8b/Xa5qVtvHfUINbF6958alDz8fff5KdjERw7hxipjfm63JF0+G
7XyB3sbJWk9zXBxy7GxQqLqF+zZu7Ye1vHn6TSgN+orooRJ9YbHb8Z8/q0Z7vASE
m8gp83SnI9wsgf4WyW2pRwVBEKRaELIQPzNerlpYQI9qo5SmGVkbcQl1gUYIakgH
/XO7MAwbA77u0sSUsTzlgnHrgIZdmbpzkymnaaV03N00uKEQezDHwOCWVq40KYGO
sa+bf6NE0PXzyFKg2b0iHzX2JUPp25xvTmUlBXWAsI7UV1ak02JXeH2gezFYlSW2
mqw8kcMhzSqhPwS4ylV/50wIdr+7oG30hk9u8vAYM+0OE1/oYrikKJL4GET/GdiZ
C6J6/Lzi5i9J4nIAStR38IrP1LPol1bviwGgofOFB9fwcec4QRy/5tqJ4HFI/x22
Zjt/3mhByF8e16S/clU2oDWmxM4Kb6bQeuAq5138ka70xTS6M366Qr/v1J/UdwOQ
eIwZHBNDpZT+HVuI7v60vw9dWpSs6L6FqdMK9guTNliDSfo7FBRGHCiMNSVH2Iup
5nhVxkaCH26VGvAYYMsMa+SPDmaNWDDQoPXLbYXOAewK14M+EZpRZ5L1b1OUYBav
lxzSX/3Mec743dXDWhORRp+mrCVNaf8b3YbnWX/LJruz1zDlMt50q/jnlxRiGHCq
FNxOWrav0K3bj+tn9sJWSymbk/6Sz1hm4183HiUuZhJlMSiF2WGpb0bPt81u+Dca
Bb6bUJmtVVnWHq1t5gZa9RgAIoAhDIEj3Ss41vI8S/PsTJEzk2XRHWmsaMuhKnPb
w58r52F6C6XkvqQpG3VvZ5KhpGFnxLatoa4lqzXztyFBENr5RVJThNLqjReSamUU
Odbp1FZpV+AXspdl1tFFT35zgzHkov9umFWp4eSPwnbENRJMo4BDnu9jVkzYTwox
fuJGc90I9bg9CafY0dK8sOjv3mXk6nKw5iecDfbEpMtzjT2go9heCZRpZPkXfvlJ
JKuw1hKdOzOPg+YUyo4VD2uYHA4z1E0uCFdTFHLCaHd61ITLxQSIvqMDFL38a1Ti
rOp38ZSdOcm3tOWajB3Zxax1Ut86UgewI5zF1dN1pwpM3ltg0iy4xdM7lMvLwUGY
LFAj6PkfRm8XqNhOu7SxJaQr3UxQk+GipV3yRRXLFCaTzvZgt/N4Z3lyDKw5Il3A
esiFEnwI5DjUgR9bALy82V4lrJx7lwfhzemZAIaKwV22mgzkkhCHliOWCvEc62d0
IWbF1rllstxHirIiX9UggGbJb8xGkodcxN+h9IpnE51YqCXk9CkJgogMq0CGYqly
YC/Y4IPZr4ScW7jxPHlNA2LfIMcQ7/azYeaL/UwGyRUIQ+Qph4lkf/XDFi8pnTDi
kt4LRIa22lhnvAT1CXCQ5PE3KkQLTaLq4Dix6WBnvA/B8nrcFbuXsb9BjWW73P7g
7am+jpT68HmEcO9LsD9kDMz1p9YU8GMotBiU/ORUrUjpZgJOB/G2Fid8kJoEICYs
YaQuIP9O/iaaWxvA837B7erPADnTW9fsW4qT5IXbUDu5zb9TEnyGTEsfUIr8gB2o
PIKTg2v9TaCHbJRvVCcLy14wMvwTcye4dmjqyyF7eJFwdl4FMW7x2QTOneb7pMwQ
LveZzKI+juh0KCUjoc2xEs3pK87POmAXc8ZRk/r/9sg4dRz4VI09bCiiKGSICiz4
TtzX9Y8IxHrFymj5vDLFGGq8VNe6U/AyyLNPH211TH4yc/fQR4n0F+B3J6+qeBiB
GlzcglZf2pxKCXnETf2utsMVUlzxiFBEpJSBIEtz944iwjYFvz1DLPF55QyPV63+
N73qqEFU/KfbwDzt84tdAvA2LE6svN3nALQxdDea5T1k3vV8xQCH3eR2m9KaCMwa
ewOlfWLafmQoyR2MRIXjZBMzTYLzHouHj9+bpcRlau6Fn/AoWa7Eh5UecvG2z+Dy
ajEbtM4W4fPHz9TmGfzAMo+5T7JQX5SxrLMyK+/fSCDwzH0gLF4WcgJt9pd0Lklt
M/1otJzvl3Bg6igsCEK9URtoxnOpRF80B07wC/P72Nu4fGhFRHw1vi9jBJriauY1
y2Ok60Kh/gCDT5/AeZgVT7j3jIrG46ahMPld783eIrgC+DNsA8JabgHgCfkbk2uQ
13T+72FumaxXm57hmbwjuwyO35ySUJHuGCYPddOXAtkw3RtwHP57VEzdU3ew3frN
tEal02tKPeO0Hp6B/Io49PybC45zEIJFJgjz46B+nOh0FTb06YuR4FjdCEwG+RG8
iM8HLMkHYbz0JYY0FLAkbhlukkkEoM7pPNY3t3h16eQJjylDcStihWp8vxVbPqvh
YSLi9DA4rd3oO70SRcM/Pg9Ls0uVBbQaXDWbQeldjjbmwb2iNG1rq5p4Nt7CtIwQ
+epqUtcDAngU6oPayC6sU0lewnGHKUp7yThXGufWBFtz2zQl/bER9eOGgZUOy8pT
6f1bxdOWE/ezH1i1OH5ZX3KkIYAMwWYGCb/+EHyudUvMXplFEsvS2pvWV8wD6uHp
ZxRsNCpb9gn7q3w7S3AMWwyg0y13G/GPM0UCAdwq/+rBwYeZP8TNagJpIycq7WaB
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 41760 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
/GMbQK29Y+AAYqzOrLs1aUNorLKGzTZ27kyxtY/WKeVjx0eGuUvSSqqZKaYfxgZM
nbjRpjlgCxYgqhQw/Q/zfrpIsqd5qqGiMdxAQPutCIOUn0UB+fkjaTmKMLCIcTKj
1naUQou33gXhXQmizbNBxSigY3ctPuyH5yvopzz/hmev6WdQCtfzMtalgEPNZOJA
K8vvTh3CndRNK8XpNqYbAlCoBDIF357iMbp/MRim/MwWX1LHg4fZ38o/nd93VH6e
6WhUuaT2SX6LLBo542LT3U0GvMB5+TntV37zsuOko1QG88CNynxnCy1iRzGFRDSj
zMlfvcBxwtzzHwU9+iekCwH9tvuI45rIKXi5Wq7mpGq1kGVmxCfeYu/9aXaMI3ot
js2aJzb49gXtR09IAMo6NlK/GsaaK4xcwDTgmdguFSByh6c5RJGsR0gIZbWKK+Ak
SCH7LmZ8ONuWt8HUqogpGGduPMV7tb8YsQRth1+4d/WEFhHnris9wrqJyC52rCjf
11PhEuIHOgWJxGL4cSqy0RIyqN0ACnujvN4+CgqjduVQQQ9K/sXfQubokAIe8/uS
Htf/hrafMk0hYpPgGWsGtarpUHZztKljxqbJh36MecUbFhaY9UBgNKjy+dfRF0n9
qP/+SJyxBIt40T4tNNK0q0XCQoq9Iw3RKqlFgcT/Pz5je8RyyAkaPhJY9gks878Z
LJqpy0LL75xkoQCSlh0Pt8evkEDNsJTxtnDAtOMyLRN2pZQbswANUr+QOVZxzIok
ipPfv7+EdfhwdFJUJQpYRTgMspyWjJxLgJYWAoiv68oQ70rCC46gBQjqaLGSrDMJ
4l/DdMS3iPZseXIb6zyTo10hdvsEfMioQZ3P3zKEzMcup+Tla34iEPtjUaKG0Gpx
iBCcautbnU7qlP3kTpEqYabkM2qwR8uuJoE7sUOx4LJQVEXorpX3afS91M+Dmyvb
zo4lNG4m6eWAb6bY9UczBL0vYcUsH9ukQSHZvWGJiIMHtmHz1zcYR2ihi4YI/oRb
0POj/O96B5dDjGPXy6s45gNDJi+oLpOth6FNAOVsHhJwZV34VNii4Z32pQ7xb7+A
O6lWm6eBb1/5c+85z251pneiX4dO6Oa4EhNMZ/k4GoVgN2h2ogUvCHbNX7LNgT+p
eMvx3fVwHaJbg3Wb9IlRW6fGk0ZLVDI2RvLzCQ4L4nIhmMxqLn4uiXqIInmXWdrY
i/5pynGXHiUAJsx5Ox6wXHCpZOAz7NtFvYI3jcUzG/Kf41VEpBJw1MMz/jfJ2fVV
4pb6LOrnP+nPDY8FQZcc1A7z3fplaD3XXwr4c9Ot43a7BAHhPyDAW9yJt51QFlHN
VxbtYz18PD5TA7TJMQrWLsImyAECs3EzpathiH9D113gyD2CsoarwyE5vSVe6boH
7GRmvUydjovEWDzHnrinLSmodTjjPsW8lyWmtKQcXUNNfsjqmUi7U6Ex8zMM5Gip
mxAqWx1n+vFYRWporbhGlNByZ+4TB3cCByP+IgIGun0uG0ReUkBBIFSENkY5+2ta
RXJSPPhY79YgbRc8zSCIX2bLr4n5mIE9F9CSbbf1pWhru9QCd/7zUIPxIQ3n5bjD
Exyo0Q/GLVRKrTiJHHzxePO3yrs7r11WYOWqJHdSYFhr1LQWkkk6XBsazY0ZDO6/
vDgxwUAmKfn+AYQEyEYCW0wJuyiU4Vfs8pfllbfsvIB6e0NSEJ3HTLZaM6ylD0gr
7TNG2z9mfSu7nYq6UlpzldwqiuDTLiyOfwFu1RDtm6pXh9n2Y+9lwEedR82/00rO
QyC6d0Hd2tYZzLseipdyiDJNLx6CidIHqSbdVIizN9n5yDu2lbJcepdkQM91JMDk
npXMVuqSRgY61/M+G4Vo4PqycGP3cBJoAJvWYiBMpkC1CFfaH+PfWKhWvHi09Z8u
tjrLaudxXPigBANb2EKQhBsW70/jlS7w/2Q9UDkxhMNV307rYv+9g8ilumKFQQmJ
vFHfmlZkmo7q+PKXy6cx1aMWgMnsJGwF0UJXUbGLVjroD72wAQolziZH6HGsY9zK
Isa0JxMrlb74MLJh+nYv9DO/tUkb0yAcB5HShKrmwaR2q/6JP8OehyUoOj6PdAZ+
7RJwF2laWOU9rvME+GFppZc0G80k0FzPffvgHFcF1f2iCx801p/61O+Fm8CGGL/A
qvA9ZvAtkSQ3vJPU5Jzh5c4GCSsqRmfS+lJi8i7MdTNn7jyjJfwHm1vsOPwVKTF/
sj/+n77URYImGUl6UiuH+xEF0vT4tvcytFvF4i5mdLHVWQ8qNVt41zAZP7Ly8KJj
/rATIlRutTPPlgMqhhyeoXoP/bo5uDkdTFmNgza7tC718yexHTVIxNv4Mhuwf09M
uRyLVcvunnxlRW4zNXRq8f9v8Zwi3yIcg5iM0pbZlRmc50U2llT6gWuLH3owGN7T
Pm4jWTrIMuD0QAt8j2YfBvuG90YcBppRX4Fq4EaEuaQPzThVvWcOqE7ecp/Fsbgq
4Ar+7DtNYlW8zakpnFIuNp9SRNzwlujG28v9p8oVW1gpjIOVwmdxwJspmjD003iJ
QWNclDIiphYpuHQYBPUmn515jje/O9mm66/c429HltDenLc/tsECv3FvoMhe1TG1
JrecmTpJF55r9HSI6C+TROgVsfRlRs/y09/l9GVoNbG5cK/hjD8Am6DP4YXB6PKb
FtWs9u7wDbJpWSIVgk3x+9HGsY6rzW5JODC8WBVl/3keGjoVnJxCHnvOimELfrGV
knV0gkKQgBfdDYDeutjpBPZCAUAi4c8djqKLdFP7adEM7dUoGchEjUQ/5rnEt/va
/PGALP4w6HdYQzo8aATQhdjTbu2r+4x2afsXCpt1SpmLEIG5mMHs8ZZ4Pcvb3d4x
291ge0cRu5foCOFvnlz0rUBNKbFvGXW2zeL7MbDFKJvvG0buIktMufhP8Ri+ZrOs
QHCPldY0J73/1PYT2DdkoZUzVa3NLjtBhnrdfMvswo0dxKA3hlTeA+h/w3nlQo5a
a6xcRXtkAqhuEVf76VHaYx6olAqkC7GnzNURnWMgKrdAKbTfBTj7v6nRf0CsOP3O
xVB2cNUoetbZEYkjpQrjtWTY4bIFXM9MhkwNf3JWsLLuH+syyrDGhqBwVi0i9zp9
wbOYBtZ40TVUUtTjV7Fyk8Ccd6OUNiXbDvDEXLEELwR/88pxpOEimEtxmXQyTaT0
dGmA1b6+K4R+lP5aiy0XAzQiFORkJTyMtMCSNy7ZRB/3nPT0WrDadDSPFePP7CbJ
V9CgphS+jzdWRKLLGJ/UzgJ5j9qTho65UdA4B0ml3r7XBXcMBTD9cR0IbB8zpia5
Bd1uzeucLnwyhxjAgjRSeKDZm8G4wMEVSEGMTYsMVSCA/XGsrGl3bQ64Aypm5k8L
ZmEKOb7UK5QjmMhAmnDC82AlNAzfY2N1PQwR7RteG2XvDNNENLxzXC/wfDF6TA7i
YqJvZUWrxm/UGV5RbIT/Dj4kzzr2fYCmexPOmuvY427IOdaJVvIxYEikstNhiWSE
Rr6oKgOnYF38qo4lyGIRkiELSuyQL2lBgSxW8YwM3DYr+PMmmo4wvSDUVydC0SNU
7hZAVrdPb2M+fMXALc1TAKHP7nB2S52zcdbOaoLxVo/6wZ0tpkQoactlltmZb0pp
jCFbDZsDaC5VW/8yvSWrkaKhyemEaby9TZ+jFwUjBYhwNFVySN3yDf4c1afvzWW3
fcSnn2KdCYAKRMrf7BeM/7NsNeASQa1JHHyyYtwlv0Enzrl653SPgXO52xEL3edd
woaRgquVC/A3KrOn08iNuP0MCCI8cAh5k7LxpLp4vrt+H424rPX4zJGi05i4SR4c
4GPaewFOigD+79EUmtV5KK1uFtOMoNwh10bSQOWg5TRYKcP4CQkjEjPDbOOvNnFE
/l5/0Y+qkPuqZBz7rmUs7zp45HBQCKbmpmc+UWm/XW1IjGeXVHMBgRm17PGZdb/n
WuCXQd8BfocsQZeefCccjtrELdPX9jLR9e4Nbt4H4JOf+7fHYwsLJcH4f1tTkGsc
XDNMWLZZfaM0FcbpKp4JHHaW2zyMdFzjH7xzaXHIrmpvrdFDBU4SuDnGGJ+JFP2c
6t9TX5gPd5KSky54nxkOeu2dQjLu/qzIFPFdoRWqBG41vYLh6xxiW7W4l5Zz50LU
xQxrojcXWJ9bf0d1ja7pkNwcsp9uaSV9FmCigNErRtT6W/zi1Ch44O1HXAqoR6Od
7Db2CRbCjFf+APhRnmZlO1lvwOv5RWhqqju20Q1Ii64SIYWWHN9HJP0EsG6OOXqG
3hDgyLcvKiUYysjswbhrgrKa0TrlGEr6YIpsLCJaVPofI47WvIc1uhTXmgdy7G6w
zQ4L1IIWhqcskPEz27bs86xf9iWzF14jrjqx4IN/UVaOW9MaLkUkK3Gm9GR+LQN7
3rttECgWOmbP0T6efOi001b2vPcrcSjpGSxmD6M5PO03W3hP0tq+KGcPun5hICK1
CoWeG7vpcFAI8eDZ+w1QXXnSdKoxINGJcoMQwgi/KShttEuNbdHuywG3p/R+Ubt5
ZOzTZf01TOAVr9UO7CJ4OHvFC3q8f02dMrfEC5UI7jS+JaQNRm7BFpopRMDeDCW0
e0CzLDzzi093hBA1/t/G8NvzDcZ+kUwXeVTK9Uz41s3XvbSVVB7lbQPcoahvrC8+
nmMtN0tATXB1IuBbSK9pi3uO8C8H5N9p0FjZfWvnsS1J5HGJVOiMwgFKQtTvKgaN
tz6hGvrypKhfjuepjPMyL2JDHLODSvWRa6rFLRdJJuD1rYmZUAt5kqzh5dX48BHX
OPmNW48ihbcBL4acNHRvYjKhaIXn++OCjxiZkP7W24J6qqx9UIybvexz+eqnzOYH
41KQEuVMFFmX0ArhWvnw4Bn5q7kjHUZIi/cllAOi9du8ow3lKLXt+rOqyAPzvNqU
7pNeawfJBazYep40both6agfF+Au1c3GZpOc74IfHBScGPRX7SPTy+cllKmcLE1A
vTxi/NaB8UI2G/ktswz3QNTNwv61tzNt7gM/NTpZvJJNBMSNQRJuOUzJwxnkR6t/
iy2mgRuvjHpyoQPfIrQPypn9PbvUC+4K0KuHnJQPaDipy/gH2yL7Li2rcN2mTtcJ
QRC7+RYYb45oSGRppeVooM9z76w7wRa0+R6aBTVr6F5TQ6FwIgJXoShQIZcl1IXY
H6ofXsioIyDnWgwjRxlFm1AwCdEZqAcdncY1wPUAcXilnhLT1CwQIkxHh/9zDoq8
8jLxuaRL4i6/7BtdCatdBZQ/rYkJBKr0JfvVchBPgQclj2dJ16KSyFS4FnkCKUoS
RxPpbIXYwBLDoea/lNiCA9ahMBs3/J4rfKyC9FpMaXyFbrS3kLv/pwQq5V+sZ7OR
XELHu6pHBEWg588DXXZ2X4z5QAFtMHAaI7nSX7CGD2pxMd1px3Pslewurp1pYP6m
sVEe/hKblQdobelMmk+qQ+RZT+0HRYUnPmU+paTXC9heifOa25j17AEure8MOi2K
TANd/YA1n4Okd5m7KOkvuPIylZb3fECncVlwo/AT1Ur0JSzx644cWqo5EYbw5Ilh
VP48mw+6xC6bKfxRZZ+sLpSdkFu+6C58UGv1k23cqJE1jZstnEYfFQEXjkHn7NOh
85jwKm7o6zADTg/ps5xcaoXmMNXJ+3Pg13rLFeWS7uUf17nqxv+cOssuB8h9RUMM
9D4t/T91zmJ5z2Vt65ZLRi20aToPpxyh2UzMXEj8kJMOW/+BhQosdydyRdW3Tm4L
F0QKNpHxofaXthBk3DZWIL+PIxWgLPQJhEy7zWkp3XGDgMv/Od72VgbdJr6QPB9w
tCaNLpmGP4iI7P9XPtvzxCS3pIBGJPUqUFwH/+oz0We6YJiXrJzTi1F4f8MnqVfP
hM8HCdXNRYVPH9MZ7rZ5djFL/DdhiJp3V/vCGE8lFb21KUBKSP/dikNTHCynr5Pf
lNPkjd2Wp97HWE5E1BYU//D1CdDSmheO8NsFVMpJaC0GHz1FOxvK7gHa/j1lOFET
PP1X4aq7+FU7myF5CEU+crKA93lEtpfKGBTpQfTGIXCqpK/EkCoUtNDnELn3DN9h
2bz/m9kqLskQIBq61SSSEB9hDmXnkvlyB4VwPDjRL4cufZCWbYgGLs3atbIWw9iV
Jd2Ewkj8W52UVOEF3n+kUsXYzAekIfJ6FUMgScFPnMfZQ/BVx5jTa/B+nJ7Bh6h4
9UBWRtgSlIt5jOvy105uI8lngpl36QbbHiA4QAIuAcRA6zBcjF6NIolVpHaTFxJA
4IDIFNEykPAakgam8DoO+AWCpr/zoF+g1sNiXnkmHXOco77PtU3KBHI0ZcwrY+9X
U+ZlZvhIDXB3DssUbAo2OyUxarDrpiTvLRoM4XbzB7HiiG5vXRQqjEqaBWYImdRa
+qlR2ZOU6HEFSvrDYhGDHQWr+vqEim3dPLmmrR+4a/iFxub0NJlCDCQNsMdAN+Y7
fwmu07fqF6ZinG4Q0aMmsTTc0Y73ftzNUr1BFc/2t/Pl7b2OX9Gv/YDhvvAeYGLG
5TWJaae3ZDHaow0e6PsGN/cxTGZUG8QRbtShB7CZ3qBhXzi2ONCnS3rJUAtFPbrb
FIZ4/MV70UhNCqFLYpjBn1U8bdCzoauxT+XOKkAK47brWUr3oMPkGwrtbfQ7Yx8w
0hlnvBUYYYIRbgz1zyx188iaXabaFKqfVbSDymfwL3jkKDVtYH4Tv7pikfmDFuUy
S9HTgmA1IUWWaVr6toebI9j0cbCwYLkiTzbYueKuoSvgS5gYhotK1PmRjaUzTXFi
68/nYtj8DMMgo5OABZr+dqcibdKOF4a03DMV9Bpe+hBErceEeWsW8VkAzIxfpsg2
50P+FixSHYArdNNIxU2I44ogW14LRZqkvKJzVTWUqlYshZaSP2mvUV402RXeYeiP
2He5Yeg0B2wI5tGK/uzvkQ3DAM2+RcGRWTXq+FDFJ08/E2oDq3Xpr/S+AROFjMqQ
0VTNRpMWybJCtWnoaJZ6++90UIHKrejuzGJ4KzgdpHjJtu8mMR6CTPr3Q8claEfC
R+Fqa80Cbgc61hxe2T9GmQtDzuL5gptaXgXSIs9UjlLekVRZ226eMsWwAuE2Vqxs
jAmBwiV+mJHeYNBE5Zqm6eF9IfAgh7nCFMpT+g/tjG4Pobo645aYTTDYoMgCd8R7
caf+fdaJH1shzA1YRZrPz+GjwidtL+K6MZBHGQIuaPObReHj4qVTRHivNi6PTydx
YG5XElVWxCKrekZw7qJByrgzPX9IgXrSIn335ygImZBKHE+kBlRrA7TJPHJH0m2S
pc96RqUz3bs19k5Xtm9WFVuM1C0IujJloIgeBe7JEbCPzCb2XFsKKfGhkzc3tzMQ
F7mFfFusZEo6264RK0k3W3xP10qJMu+oUGcPcxmSqPtmMrzPaswtw+cp2LoPOgWG
39hN+Hf8eicGo4MQii5bBbE6RG4p0nGVkdj11JeqRZDLPdddjhxtQeDvK0A+NDyk
RIsthv+xrrJyVXuLl/3XsvEOPDFMMRqeKyf/nS2lTYTf+TB6/3aEnFI5juWmTfmG
rv/lU/TtMXY3yI7LjCfJFEtTJi+Q9cOIIgjyUn+EFk4R1q67J7SM2apLVljGT5N1
a8DfLt9XGTqcsU0r4VjnZ777FcK7DNce5tuiyLBLDkeI9O2v/qWUeMs0wzjS0JzX
eoFdpSU25rIMt9YKWLrh6PxqBX/JAWr7HhVQKIn4YhtE79cFbvGtosigZCP2MeKp
mmrh/rVYQCtC2dR7jXaZEWvAFZP0sqrx5ZL/dOudas/Jz6ErP5+0vIHmhzswBJ8O
0StX4Tnl+PXb33oYPTpb7Gn+eGFmDCmUWYN25ZhYStoS6ZwX4JWWHqE7deolYufn
O5XWKSzn+aRuL3+heM61UV7RZQQCbEHJW2UWuQroGkHwU9+EI36WA0zdkhJNtKcs
65i6rmltU7ROiENT+MHRsrynH6d+SMoMYDb47x1s1Pzcnfn+Ie26SjhNRfXJF+fL
tbe8+xZMtBVakadqpGHIH9WBWb8t8HipqTj5nRKem1SmlDDQCzoj99YDGzEH0Yna
ByFaVYTfGGnqmXnhfutHSh0824Kt5cTylw3U4yS2ag5SnPRMKhI61Bok+RN6qGpU
ic9ZZA1oetg/Bh5DyfsqU+BxyY+upm6bTTK35uYj9kk9Zb4R05g71MZ4i5+N4p1B
vEHnWp4fXPKg/5uZV7MOcG9HozbIunKgaOFexYAKq5CvelbMqkG9AGqQOqGa3UoZ
FTx9mBB9AYDzgG9mmwH3qRXKshPge3zpMlhlHBzD4bKt7Zk5XrHZ7BVAsKJWxAxo
WkwkyvZ5TZ5vG367U56/V271tRZhElSUTneoYdDsf34OCJ0NM0nlR41HHCGP0h8t
McbaEFaHqSj7snEfPxXZfHc5MhZE2VIor2tKhl7T6a6JeJJoyQ7LTNah0PYcBiLY
mF2Xsb+VfLUvIIVHnCkF7VbOShTLfvAFl7X6gADLpCgE3Dh16CSSToP41g4ct+b0
RLwcO1/Hnvban3JXyVARIz1NGhnnxpsx/6h5xwIfq2PFVzfa4/v1i8VfZrLvIdR7
8B+4fHABxKSlNvkistWOuItIXQDgAG82DQhLCcy84yG9fVH82Kaeu7D/GmVpJ0ZO
5zIaFZvOFpASVbX+FKi1eqiTcxiJDZfDDLymvQAhihks/VHbQD8yIS++4bNaSRmL
LHrl1uNh9NSkI4vG21YPG5icWempyZ+9N0yTwRNzDOtBvYfmRw4VBpaLNFvGyuvJ
++DEwqEmg18JmInRzJNjgb7CI2Cc2ZdU7QmwR5hNz7kmDH5+69kERqDCfRWdEc3G
VNQCakHs3cQbgjnQXLpn9Kn0OtCJcBP8iRPPjf+uhZysUvVIPPZBDWRH0Mb1W8NW
/fZ585J5bncumySRimOCR142Yd52TjsUTDvcJXURei/OEKOjn+AASkZTDTNVoJa2
bEbC/I9FUc8qC5+c0KrYKQltGrV6K6SjrpEcQVGOvo0hZYTlWB1mO2Ar7J6aX4K2
V73tAAptWLN7jL5NBIFHpxl5NI6rChGOs1/P/FF6uuhSqknLGN7kU0BpFHp8e4gz
T7KRwbbwMteWoxyjdNgeZ5/wU5R23ef093ksH1VL7ZdHl/udMCqgXkJiAM6yTVuI
JINmxS2p+AkxFMaGakWnXbrKpQlVnGmMDAGP45WcMLH8Eglu5X9Qbv9UN6CvCTmp
hJqSpIb9iRKoGl26P7LjWmbaZ0V3Zno8RUCofwO4RrDvtiLyAM49CX159CNnWTbU
+I1S6+cfIeM3h7j1JQ7Xi4sOKdUCHATsPSPkJ+7HcIKrwaWCB5sX8lkQVPHkIXRd
ikdoeTdrhH1ZNByMf+pC4uJJ0uleW9WW8uaDtNhuEHUH0vhb+3sysB1jG//Ri3G5
S3ylkPs6eZfyG+yOFWHWUUUF0Xg1H98DTClas746DQZijkVRYLQrBaygt6wBn2Hg
AzlYvvv5IvP5HEUWhhQaklkDAJKiZyutswxpkJhG82g7lDVNkVp7JA0AlViAJAQc
zj4Yuy9UwSYYfYkyRV6BWvquV/U6xna76CAGOSr5eTSV2LBiqSG9SljMZY33Fc/F
kbfFwweLWmRdfgrCvTgOXlREkYswmWT6r7jgSHgtLnnsiV+yvttD72dWMhA7gkrW
GTrl9n7/uIrNZiZVsq+/ncDKoGu5RRgyxcCwRsuUmqT+JofR2mjiMwVJYkZ9P8r7
ihTK4X8tYeM0+fh6Mdq1h9KIW0nq5yHqRZqa9gY0zfT9xV9/93+JbK6irCQ8WYVn
CvCmOloZzaXWI9djk3UgGJv/F1TnZuXgTER/GxjUtaT7v1bEmEBB6zpfDBorpsB2
rU1OEw2vFSo9CvEtu67A07N185UfYDExvwS6B4yfXe5ZUKugX5tZ+tt+IOS1GJ1H
sHCaZTX6QZiG8M8qWHFAOXMlFt9h0sgT4q+OqpACysjxZlULmxlwInS4U+o/XDQo
bDV+O/LPqHVM6x+uopZYcvO7jQ1WGFcViTYmDflUQSbZ1voD/mqNcGnOG/ZW1kR7
ajOQuTMn7J8AIPouO6kmYl3bg1oXW7N0o+e/M547YCJCvo8n/DWTdpMnjBUtVMsy
cmCpYO9kp0zzzqjMz2NGzIXEqNbNM4rqicHB2LC+zKV0Js+78Lp51EwJug9PMjR7
uYPX/2GAR6KXrNRcXdS+rbOEgEXldhh8L5C3x0cTaSkIU4Kx+NMTq4zLPM2FVesg
T/ak/VnQXCi34kLVILR8m1lz/ayQ97kuCg3tFgWKsjSNseG1gEFNPY0rBzxXHi9u
9unPVZWY20vnwCZw1bMJa/CkpumSWNYTvXG5R4g3rWlPkS5jaqSkCljixu4clslV
gfDmGXQ4neLPxVRsMws9hzzScBuxgytj8mhi9BeSsjEGUslww9cqjeY5pc14c9jh
LD4wTPqOqqkrM8SYSFnBl33ucBAqiWYPe8ZNm+pdmxBlD9G+K/mJ4rgCPC5ndiBC
XWycXc0Ubr9FbnZu0iop9TyZRfI+HloFlKn920CIJPICZCFA2yBYtPcUUw//jn0z
KkKS0neBSXJ4djIiF7QIOFAsCfni0I+aXN6+y2WVvhNGyXzmL/WLmdsTQ16Zy4rX
W4W58BCV9udyeupKkLVpSXE6R+14ZsyAjNvxWxGmzkGCLFVy7/s1Nr+lGEbBSTzF
Nr7S/0G8G/h0MBDPf72pku9OKm+B8lEnbvXSifZcb4D1KOCws63XSCYiMI3jGqqV
rVWAnkKJvqd+qqY8/HRL5m6zbvq5IkyZaxqNchO3uhQLxYpj8YBFLSf5W6+7jcKV
wDlOj3bUM0zh3JLstZDgx9fH6qFTpgcJIw3a3/t8g+1cKlI72Bd0KeQ+ds6NkdhC
jBT9CepnUYfmA3aNWEg6hJUdOExPtY+rGC6XbRZ01jb4ko2ZHFDtFDA8rf0pVjej
fq84iIr/sApO/8QctI3O4WQTEqw177JiWdT1r6Yq1OlFLSuMkJj1GPvGmWOFVk+n
z2YKCLsmAfvpLqheOMizm9P7UMlOXl7nZcCXU2W5uSQdRE7Obd4kBKsa8fAVTKh9
z7UOMGWszpCsl7iUkSiNgFcBx7Opjpian8Ii3SjbiFiS+X0ZRO++zIRxTHEpENXp
n3cKxwXeEv/UIQKHs/lUfbufMwV1bJpvLuStPOsAj6zBXH1PElfKd0n7cP448sC9
yYCdDYFn1oVioRyKHq0ZyZd2Tzyc1plXRHo5EfljVXU0/mi+8RTXIgYkB0luspmC
Mcxu8kionHfI8AUfH1T90YgQ7lIfsMJWBGjnQqTJo36p2MR1lRhjCMR9xG6EPzUJ
qCyVWBphLVlvyINWwt72QvvyLVRmgRFVrm+z8uqomTO9rgmEvDHYVQ+qpS5AnNnW
gp8xQO7kN61txmGqDfeN+O54EYgwUolTUtx4iyU4boqa8JrWb7XgyEbCOz+4R+Dg
hCL0pp3dHm7t4fmoWFk/XAFSmHENMG5HOBol56tKkg8EosQTsxTp5eh2RhX0qy/k
buE5NWpq659JAe80L6Fw++ZvbffrLkDqeEDQE3yO75WssZuCCgn/oVALNszZ30D7
iKkTKNAk6qPeOYSceQHQTsh85EkPZM8NJ45SWJrG95U0waPX2waGNGLgrKu/gY4T
+C3SDGlepCoEJFT+T7ckutd343IAJwZHUDyArP1bHyJWViU2kGPsonhYWd4lqwOL
Asea8sUrQ16tOsjRMvW33pqb+R5ZzEdw8czf2bq56U5RNoT7/O/yLk6x8h1PGP7V
xeRnmm7GaGSLB+IFEC4AyphHpXabm5rDXkWfngkgHeYt1l9hO0txxMcoeUF67ATe
llqbvCRQ/tnx7DehFq9sKtStCt3Yfz3Gh7RkHbWm2Qyyk0lSWBgZu0LiQF12D24w
6CAgkrW3BSQWkk43JS9ynwRDkR5PaPtxc99WqSKCyrXlNAApK5txOWbb3biHM1qU
Dv36aEHVPqXhmdwr/kowMXA74xRDpcJ8xZbgC1vE2kM5H6EQv33tPrjcco59zHMW
NWB55eBQmzz3tYJQX2RFUzAnJVLp1gZcf3iKVr8wVnvpsbhnrG3FD8hkBUGGBq1j
0t077xSBW57u8Uw30wgPFPWIn28wGB7mc1AydxIDtyzc/UsaB+kVdCg0OBa49YCY
0ZBmvPQ0mk53jVpDurHpu4vjln8hoN/54F8y0VaCJurVtmp8Vl3jp9kSitMpc5KQ
02qAxDa2fXui6wlerz+Kcbm5T0vnUZw1b75TuOyd/BFHfnJL6HvWoj6XzqKUG2s9
uLL0/Xl4H4EZA39oam0y3dTc3yqwaSpmOK20hRlEnInWm51HyOKppQUe4HzcBqqF
ZI3RYDSw72wPbQncg5B8IRztYHseGH7Qpm9RpxFBMPJSN2Edg7XjnylgtHxOzQAY
hzBmylsUrbSfbwoxPkDNJvwDfM6T+JJUfT+04KQ43WCOzn1E7GE50iN5b7oJejvh
N3/9R6EHtXe2xqITCTVPr7jDK0CCvWvBhtovXxHDvd3wF7wkGTVYO8BsHL8hedop
Nmsxm2kH8CvPhxc9/Ldg9tXxuTfrWje56TEyy598DLIh5YAXnGvc4vO+nH2Kg/Fp
dGVlV+Ntocfx0uOftqst0Pwj8gyB1tgLB/jFYDIYBJ8zs73guvQQINyw3JD4tGuO
XihTdKfuzW2KcQ9bf8TYSt7fHT6VOE2TOmS6r6m99zpmEgV9Egufjzn6w8S65Izr
A9imjGAf1yFFgmpcWJGO8vL4ezU/UTxL4QCzhfTAJ0+TWHLanNcYYu0d5QfyMJyJ
IZh5GdUelhvv7yjPZLsk73UP0gx1YhTxowtbHgfgxWWnLDYV8ODKKIZnxLwrVWPE
JlHuUfTlbnLRAznNYwYA230MfYKP3lH6BM/wJ3kKNCg3ETVNX5bveJX7XUZPJjfk
C/qmGH4BInpROAkmhD55T1feHSTlVBQROiZt6VLV3ZtEy5uT01orVtj/DULv7S+W
YpR8DhAo+nk/tCtGnVFI8hJfo8ARkfR0e7Hh3FlsZFeFGUkA+eaq8nWtxufw/iyG
q4k51wfcAtgBInJCWH/afOSfghF1baaGLpP/yrYrYNp70iZtXbyY4SVknBqQYzlG
BiqJWuZPUk31e2dfvMQlSrg3tKsoVCGJuB1cafrTdrWv4NHklObPbLkCQpC2joCA
t5hwLR5HgHT27zJlHssBAeie3NDTTz37EX2S70IZGvF9j+Qo97Nk1/b52a20zIUz
nXR421iBfa1KGOE42w3UjznX+96INpFYoyTXafT07qU03vj/wn/M3EL+ypscYZI2
NOkOgYVCVuPtVHbGzqNM/hl1i6aO7mpDYFVESpU1jz9fLOsELunTG/xf1qgc5Um0
A8MFuL8CG8JGV2TwnBgmeQRKZ+0DWdzPda5O2YZdnhmRgkAdCXmmqdvZYLRoEHj8
sx7wrGwm+Z+oCDcoxdqNISK8kvfYpr/DbBGZJgWEQikH4sLRlvfmvko9FGd3SJbZ
zaYPr9obQfYsTsTfTvIBUzWsPgypFoBcSNefUe5c7e2ZXQyhJuwjIQIlq3SsmnND
ggrMzhloqAEaJGEWA2UFKB2c7ZD3EKHeHzWyU2Dn/8cYNlLxGZ9uNtV6MecolbM+
MCjGugghsJ6kPR9JVna/t7FlHdeegCbtFTtBPsXJuB32AzzI43aYntwPwBa9sFza
Rv2NdT9p2GTTou+F3dpR+lr6C4qXgWBuJcC8e4cztEu5qKr4XU/rJdbpjtyu9w1T
H0WJoMWU+ZR+lUSZbkt2hM7x6kfBrRsFhT8Ma7DF6Mo1IXjCIvcQQdBuXTURc4Mo
BXegAX2xym+4hIL7tyG4LudzoYlnL0t6A/lO1g1WkHxPUzFokvZWy9S6FDg+KQrl
ZkJ+BWZ8b79ndPW3ituG8IyCle6kugxj9ERk5EgjIf+GUvOE1roUb/TJC/Zgyhno
xSkeR5zQwWvtooAY8hMX47PBA5/IAzA8Q/gT4pbaDqfl4QOtzVBAxfXg1gzUJ9vH
Q9PuRoGHsA0OuRuscQoK+OqVQC1kxLqwKeichTeuQGzxHWWI8KMXAkSv9MCguPip
cqv0fgrGwwfSDrIpqpsovtuSObGUTHeJLA3x/kOjyCus1mQSnpT6xF66gfEahn00
792bHcV0cssR7LfVUJ7P3ErMqtHP2/4ck5DegE7iX4OiuPuMcmfdWLK1J3ovTnYw
JQaMSp02WflKSb6W2pRO/cP9fYbYaGMLMoUbgtN4S1pxtFTxJxjgMsQjcCzHTIG7
UW952dOS8wvjELK5N5Rj9Ls0+mjuCSMZY//EDvlreY1CfwWLByVutwYYwk8hQdgF
2X7NONn/pqG0KFfhZoWfVfw3tOMpvRVc1sPUMcgwHFly1cUrUbgaYCcCGknWKa0x
ugv+y6TiYmFpmQhbp1zJsGGat0F6PP+ZN7v8WWP8eOhKM3P45y6wMIs1bJDn7bzB
m4DP6zNvdNQt5MoQ2WeGAZTJhfPx1AEa4hcWm9cyT5z2IFGzOo6SHFuMWdTG9mMb
TajbXwKoajCerlxACpHH07dKvMVZSULCY8WX8ZjA46QpfaDNsX5ury8ouNjx29qf
X57tBJYZQ0w3xyjOrrrQ+xWWc14PjbIUw4oT1pzLh8wmUvLNQnN+4yFZFmN9ceBT
RCVQSqH6ycDBaBvcQHd9j9iRVcvnCwxaGWwFXHp0RN1L1QA/06B2sgk+yVrxQiIC
Am+8WJ0V+IT4x/zr/7n601PXJHpu+DYb7aivNLCsmv1a8yrEwJ+puFS5sJNQ3PpH
VmvXuC9kQqMJg1uURhN1szCcRKJ+5IrnLt7jO/EfQM9QdCBNMUe6VuWQr6rFUDED
fvpUUpow19JpsMv4PzWX+binE4j2gCV2aDCjMHrSiibr4gjwp/SNtuKqnRY4/Rpc
XR69NcFKJJOehJzGSfxpxXlQLYpFElgOsJku/HZPNkmEe159NgS4A9XVLlgOlF/d
OQnnkWFlK0PysQPAevw39/1AqZwzBnSIDAPDtXPVKCt0jTkuYanZrv7T8KWUt5oN
B9WKTKGgOKfbPMKTlm1wIWhtHlObjBh1IjG/yWJ8nbjCUXwBncfip08Ooh3PgKSK
Cfr9VdjGyARP6RMromsfwLaoQu+hbkqLCqGXRv2y4q6y3jxxv1EG1RvC8PSw7yge
P7R/lGggiRUlG7sgli29xJOdnX1AuLNiMfgUXDGkce+2IR08co+l1lmkJAbwOOGO
fcNk5G9coxcnEZ6u99O8F6orWMdJFIUDHFl1BgRrflnpBdKk+EQ5OBlKqXLTn6id
YMzmCpZ6skIAqbBQihie26ZqfKBuXoTyJEQMQw3EDLJCdVLomLCOPv0cnqaDzG18
iVF8QD/KGDnpayD42loZpdDUsnllERL7xXwAm2trq55rb0w/XY3v34nyQg1JUE6u
cFHdKxkfPW0Wv3waxsGxYkM2Y2LnNX6ExWIYmB+5swF4PH29lXQw/3UtvhT4qHdo
xROsJdoJWuoPTh0E0DE1DBzPFc8L86eorsOGN2ftHOF1fPkKkl73co/sZdr2Jjqz
4ZjotOIgftgpSHwWvoo477UcippE37aSD3ppbf9qyGi1gylzmcrXOOhPHwwVe3s9
VavP8VAPj+cdZss6gUr44UGNiGbV/6ihnZAvLh0OJs60nOlM6pYKej3wNIAe9+1b
hPKMhN1Hnlhie+dtBnejB1+3zjVtOxKns0ZxtuMPoVNqt/BqP+kFJE8fnf5fJhNW
oq+xOdtf4LmndMe7X8GWDzhQPMT539CC6NKujHotp3aGnNd3nFI3r7xlNGejYvzo
XWGf94eB6m97az4byF3jOT0scZpJGvf9JT0MY5CaV9cvDjfhrLxeqKhsGd9HaXoY
OOYuA6Dw7DsqzRIirPbKkQMs4b/FqSpxd/ppcAoKkrtxe85ZNqw0evg3uc56+QUH
lABkFquInDX0uV5lb37shsOf2D+p0Q9v3Jm6hm6tw4Xh6Sq7MrgR6yceoa2EOb1B
wDUJt1C1Q2w2OqgpbqTAp15MNLPFpepulMJlMd7N9QascQx4gGJVGNbi5LN2w/7J
hKkdTv2oB6K8X5CWB7IvE+8XBHDCJZ7/MkjFf2dNgV6ncOucqLq+NyyB5nJ1+ovx
/GhmKXy8wbNXtEPczf4LZEtR2LuzYpbSpqicJj+s4yqtfEAfOZTpsqpDWFIIz1qu
PLG+nutEGhDuX41CZaDPx/U+/ZJcPMbaYJyi3bepLCoHWBlArpFsYSx7yK3s9vL2
vIaBiGTTgU8wwycVV1ANqBcbXzcbe2ZX0RuPsOX0hwWW7loN+IJ+QBjrWmRY4qoD
PGsi1V89X5MvKao1cXUQ3+qKq1ISqS95qq6S3p0ZpezDBuSzqjmVz4j628AS9Fsw
q7c+lfrbdcTI127bJlJ6oI1D4xNiI6uUChHpQeKvlBZA5Wb6EcQsrdE6xWnQdHpS
aF+S4hFWGTvKg6dlNfVoMPs+PkcffEWKmyqn+aLEPiscrVRod9V2mhIQr4JynaB3
gUrtR1+Vn0Zr238il9eNE95J9ci+QbCZRWWznMiLJGNZFvJwA5/+8PwfHRcLH9ae
ZKqa7rf4gjqYYBNy7TxOUSUvJsFIOrA+WupC/PP4kB0imYowTn4/dTxX9PaYcqqV
+e3uG/Kj3JIaqkzOEk8EdIjQBde2Dc145zzixJex1mq/OQEsvTdY2sy7ft+H6W/J
hME7pqVKPStjBtOFIipwCusX2rbZLGrmj5xGc+gV1h0gEmkzzpnHX0ael+nZKCNw
Pv9FglC12Zlsvc7+gCTPiwj8hu7h6e8WqxaimPSzmq69N812ICr8TEh2+KAnVOSM
qI0xR6YfX74CCjdi1FEA7doXW7ZZKlkRNqO7Bz33YZaLLcydfdFVQp6EK/sMed4y
8rJtUa8DcmF6uC0dCbo/Ifd5rc0x2APcI/kmLG/ASzJP0z0njaBGsz5wE/Lugu33
iy3rm8+XKlg3e178kJ7DMZX4Dt2RaXoFJa6P++m4Sr6CwRrzS9S6JhrYVb/OHD6u
4F19va4pGam/H+GtfoSABkeZLwvwdpyaxCVBkl2AUZCtU3++oNjxYiIIpxWJ05Vw
JExZDHhMUKkRT8z6v6yOvEh5AZbU+l08Dx0fHF9E/LW/QQj8YNoQKNWH7LqWnn37
gNy2n5xl/njm/58a+AXMwLYCNsREV+CmvfYBImd4vluxVfbOi89Gd8JyK+xPTwaA
TeNNzrouY02Izh14/Ibo3tVXwVcRygCADOOxkaxqZF1iqMk5nq447OyPGwbSy9u8
QmIEjNJ++oXQ9OHK0EsQIGUkFHpx7oQpUfy/DhAqpi3D7vTX/eF/iHdtCkPtfKnV
6zd5xIhdR/Fx06AXOHLWRloHMirt1WlIubMATQbJcC+ilmnBFOrvG/4w63yPEt0g
Zle0qtrYUADWD+zAjbJn4sqImJ1ERShQqyKkYNQ+jhW3YB++tP5NO0C43TlZYdKh
sfmnr2Nn/AihV/KuvfR9fmuuu0BoFfQxEhOUa4PoqN9jD3NYvGEDeZFI7ahYtM9x
/DGcaRJY3+U8WrTJ5ZIz2cu/HOq9S44Zpi9xJNlIiF5Pg9KTwqDCiHpA506XsZKf
LuXzgYw0OKtJXNToDulM3mphurLPVRT9mx2HWS7YReAxB1mcDqUrxIa95wjHJg2x
Q8RDxx6OofkLfl2CEU96ZgMvpo4Vm5PQ7zmYHTtUOI+gFqDr4NRfYy9a5u2QwPFC
eYfiEKRvdi72dFO97pa+CCmMST5mdLzbpGZKU/Hjylo6I7owAwiOOKp4HhAPnAZL
9XkL4PfWjCBVHWmaZueJ9faoDN2qR8i+hYsdGf9H5qPireH5UaB4CmBl/ItTaQB2
zYtGsgr7LJvtu1sCfgUjniyWuZZOKX9sbY7fjy7zBOg3zXLSe6XN8lM4Lp0P45I0
f28F0v9+84sNZFGF11s3Dvxc7T+JVeHIq1+e/iRVWUy4QX6wKY+ERFg29I5Dzhz4
aPs2D9BYCGDbm6gpUpvqAmRLiqQpY0/yIBTqPsGJz/nY8ppZ+qVSaMLYtN3VuNN2
ETt9MhSmvcChle7BjD4gYrZ3WjytDEFVECqlFdUT/VJr9C7Hm0TwD1kdxzvZikx9
3murUJIw6gDlSN6fZZRO6kl7ZvZdYLX+Pj9qOBvVpvTQr+AOsT1BoCRF6ek2686H
ujYxFlJndokDUgjFAhsyeML+XF1NuPkO0pBeW8q3ffUtEUfdQV3sXpgU6qsq99eA
URxeeWfoor8u707mMyLervhQmYQKYRFWjpD1oRUdWW9tmmzU8v0XbbNIJsZ4cSI0
/iTX+e8eDJ5xr+CyLuWQ3Ml4Y5DD4jN8ifKPQEPgeabEAy0VBIqsH7mAspDsenK4
kN17fBkFCp8tjZ5T4Di+lrmyfK0qGDtNB3w5HtsbnlZwxjKzS3/tzNRtcFkZgE40
oug5DJVur4g81B6oJMJ6qc2YoSB2PYs3m8VZfO1MO0YcGaPpjXPQ0eHylruT0zdL
mg6kCrshIy8r0XdGYGbDznEw6aeemxBXktged5NUiLZToby9zAawXXJukV3XMqcl
Ig2alnWcWK/N8KRtTyhY9jfBJ7o3yWgKrWqOHnnsueBrd/9NypOa0mdk3gXhzjOn
ZHeA5/cgo9RuqWeI0CpF7UBeDTeABX43PVCOXimyBoELYpAa9N5gMdockAfQB4uj
+wiTUl3gOkT/IhepXIZ7Eki7tIcq82SXp892MKd7YeX0zYNBV3ZHJL8SdBDW8AEa
bS0iP/jCiJXEJOWhm0SypACzz5y+eEHMtsqUhmA4bcbk+3VBCSmskHQECxbeaXwf
4olEi094c8jC/q+N3BxJWvCHQDNK68X80YFRQCgRg/NOJuIEE+rD4NO0EdfXyeJt
Rg3fumZXY81/vZ42GavEJeELhwoqnTzfPz8buv0/y9QYEGVkmgbhNayAaEawwyrR
1p456K+it/FKBIntlxKrY9RWJKVpNExFzagV9EuaJNCos/P2D0970pULM0gsM5MC
jYFqb2aUqp70L4L7RiWFXWOoAb7lKAU0IbnyDjFY2FDulRrPomkpgV2RG6iT+mcc
gzH0SzZr/P0s0BCO0Relw1p8J1Vs3Wa/KFDuZfPcJmg8L8IIWGW9Cnc0vVgqnsCq
nyY8HUe1j4XAJr4zrcdcLa6AjjbUEe9GJIU/VQHTPRIqWJ0qKR+K3cxGnxRJyP6X
K5g3hCIXqN/rMlgoDuD5CoVXA+mtGuVBj+qcPZaz28RYYxHMjgCu57hUTkqiCsn1
R4v/xGNxvXbZqRqa4SPVlzOcIDwvFU2zFn5uUBoO1uYGO0lhWxpM/Ub5NMWvPHW2
frNObCm9+MQiDgKHEZCn7FtbSsj6mFlF9XYIexS+7plncb8bnyZeQk13e961zwD/
s5RIdpkUXTa7zRfqfKTeY6JlWS+N1drhSa6FeqjQEVz3q0fBs6wctfZ7yOFgihoE
1x+n4nVO98Bl6xisL4G74nhGOtjG2M3lyWM7IHZZU228MKnQPyacVcIrJ+/42ALi
RywLhiJ2B0mtRQoHQs4rv0xHstDKNlEbIpegx5HKrmypYoImVmpaQJaEL8X7jwRc
JTPoZn4QZZwJSqw/rBwVy+VQKNTz79ywgrauBwg4AtzymXrcvFBSrbAtP6I9aBV8
9Nn+uTNvxguLgpKpOkSBST0xKDeWN+JVh8kWdAasTxiYC5070LTJLFOBQ6QiQIz0
E2lDMIrcnYKjbK3TS9SzCEIG9ychRJb5fQWQrVMgQvlFJHoDL/0QSxPTxhHn6vwG
aMMCZ1lf3HlZpFNbu/E2cGtDnJm3habd5SrdHQ/13HZLNLJBc0xjoLjf4W52MJKm
+5LO2HW7rwmw2hXl3M5l9fyYlgfTmzEwyAvsWSgy0SEI/bDlduCglODgEEXfrrIv
0uJNstDxoKJq/ysaSRQolXbcOGsZitE+ESRd+B5dvxeBm4parOBHfIySPyeznf0t
Bw4OGG6uwGn1Ks/SgQpyI2t6uqPzEUKLEvO2745Zlx12oWO6xtNhXkFuJZfls6nP
btfSM38ycqwX1BarIdWYbNEfckQU6RabeuZRY5Lbnc64r+wrzyDnobpowbxEzJaA
EeAnMWLOs7zzNB5CK9ER6EqVqgyiKDjGXKAtojzg1EYBHqpZWtrlxBPE0NphPHWM
+lIEkpQxeMTwr7LIr29PNbHK+/iXElGyvrC3bYctXNHX+bGlO12nS1RR9GpeobZL
lPb8EGSqgJWSyVuenCVYbOm/paTxk/2pTYN/wVvreQjo5/I/+584IjaCt5yjF/DO
jRDb20jT/J58fFm3sJ38VhTE+IsCqWSAFqIhquT9A2LzntiZMOXh29hKxvQIbg6X
WO4mgBD4KgQG+ZfXYM2fi66ro6L9DwZDzijE8uCTbjbwuzKbgNokTWojuCcv5AI7
cuHC+Hsb7wmi5o9KAVUXze4Aq7ZHtopwxOhgudrCegyvTtpK1Rllx0Biy7xMPnje
GwerM8TSZodz4Fluc+wKYsaSj59/AlWRxgkcnTE6h82tJbOzuIz8Nbc73UmfEX22
c028a8hbvtKGI8bhIyivGmEB52v0ECEDipijvMdR57Xl9p3GCt0FTvfmT50Gk9Hi
+WaMnykMt/GPGTQ9/HjvuWudvjYfTnmKdtgJVBbfAsQj7QM/EtQvdymUK3BTBT+Q
/CDTmvtPr/XHVW0Qhjahbi1NzilS2ZlQxk+6kkSGhAqz1QTvVd3Hx3Cf8T21VscC
XfouXNNhkavbTB9NJQ23rnS904ixapwIodHS2Q0AH2kTUwxv1V2Pd1aQEQz+8xg1
cuEs9ccCMGQNDKxkDdQQlo6LbRL2ZFbD5jpCuHSQEOHhgqlivij6edHJtN6HvXKq
c96UirfCbGikjgLx/Gd72GBSId6TYojQt3ncgguFAkMcalPVGZVqBbKN/RcT53Gv
Jt/yICD2oDmRlwmJFzOnCXRnYF6LMS1sa1eD8O4YspmDFictdZ6srMKHxBc9MlTq
EfyuHTNEjLUgHBZQ5uIbVIhzPWInez3/TIXV13Gp3Blq+sByjjOkWrY/nZ4aNGYO
rloxkG71XwVPG3ATIPdVu4KfeTSEELfXBhkF7bNSJaQq1tPbR2BVoqAYRcmU8Ai2
6JCT8JYLkxy6JGyGm9bvp5UNS5tp+nxBsRYyFEannY235Fr0ZisM6iAvjl6k5vC0
nMom5IZj1qJlrqcP7ZFUvd756xZA2cdq9s0A1WiGIQXR8L4mPgrhW9zKG17r68GO
l9dy42flltDRg89DDSpiZWGlRIYS96TKiC8bnFWsuOwVMgq2lA+bKKRwZ+TPyA6l
l523d9FhRZEaDSALgdxsIhCPOcUQ1/1NO5ARg+RSsezQy4gfpl4TJLmqvO+OQDg+
rTVirrELqDBGloN+CfsyO3kFVSbS0JkZWaDSGjgZ5TVGZSQ7t1nRj/FJDGUFd6+7
pKdymUnjrXsuc5lrb4QX65cQaFXECGJWBepKL5MYJfPYs252clJuqfCow/xkobUi
Ia1J1s+cDIU6zgGTfmoQf2Yv/iG0LBmQW+pxPQy1hwriO0OsLLRFGV5Lwrbx9SOC
1ViYdlaKiZykUpVBI5xdRzmlY2NQqD34RhE0ZKQai5TZqz6myEvbCoc2sV8MlgFc
tEpJY0OY/A3br7024jsE66mg6d7nspTgZ1ldNS6uROSzX/CTIJ1L2h7K3N6AChlk
e+nu2RGI4ZahCwroLe8Do8Txr0X7HtGKSsUEXrqMTQqKe4N0DB9EYK4DtLWXbC2U
W15kYcDA2pIMDC/SkE3qcgLxWzHey0F8HpJUsfhAKDjm73jgjB5zWUktLUkYr/3J
65Sbowcp2u7Jb9zpeFEBd/W1e4fRzHFzK5qxgi0TJu2hPZ9etLwGc3N9b6Dn1spG
Zb5pNMHQ40IRsszhIs5dkpMPwcnBpCUAXVXim9lmFg9JYiP/T3ImB+c4SGan5QxC
7vOFUGOLdzp0cNtYrq3Rp2qsyJIqMHvs1+dhKowj8Nu5g1jo5/+1bFUlNiSnGy87
Rq4GHYT4HUz5SqQgqqRl0+Sx3uVt33y0OtkC2rEgQG0mZVqmGGisKr3omwJo3gpt
Do6JezIGFTfmzBcnKgvtJsZV5VAaXNzRd+zufNtWwWWCV5kmS1TXqvzZNP+U8g+/
tvKGiqLpOwajbeseXJtLerTrOfQhOjc1YcBWaeuHkHWDdRSeJYaPy5GCC+iboCEx
GEFCh3+5ANqjvjkQC6P46TmhSqKy45WCw73xo89V0O7L5EhWKIBl3qc4RkLpz3o/
U0THXvSJyoDVT5Kf347lXjdkfARbow6bdLATknqS2+LTL5HIz2/R8St/9s7tKjY+
CLjGPZtw/OqIbp6cMBJBnPS33JuNKfSEE5EpYOJg/8TxO8W1Gv/J27gx8vI2JBSJ
xstTY4SjZyhH1QA+G+LncoqkJQrGpFrblfXgoJdYPKOlAB4J7fkJ/UE9e4frvANc
TUCloCnM5vt7G5rDOwRcoZLTOBvaN5K9VApl30kd0lIHodtOwx13ipJXmCz3eJ1B
7lQVvfEuEIyYMWcO7Pp+a8zTGldFhcWAVzBJvD0bvM5i00WR8aq8GlZwQC94+fP2
z3eOodmgCOFR+e2dIdp3MLvVNhQsDtEjGZVX7oBVz+RLhOC0cBHbQvzg+wrU3GPL
gpVvbBIo4rGVCxuCIZIYOMuCJ3Ns9d/3604v1qXsdPEFLezCLOuUpJwJuL4vxl7t
COuzGDT4XDgugLD0kkSyMQ85ezCLWHOV75Z2KSp1YhmKc6n6PFMe93GFg6oFiWfm
cCCNiZ8tklGesB9jGC48dJnzaNtufv+4qbC7pxIxz3uHyKakZ8QncRIemnXCoCbA
ufe0+fKcMrldyWP/cXtlgqlV1ErfEVJXaImKXKjfq7hSoZeDggb8ikEiIye/d0CN
QKxixzCbmIN49lmFhCsSW8oYLWUTuboYtJPzEeSWjQ2o35s/gn7SrEgp7HpYIjgC
TtT2Ot/IotsNjg5/jLVJkTwReEEzCic6VVGeJQicloLzgzHujXE8nxB6Yz+hgkiT
ChVN3HUsO0qAryjtNweffJDsjg9Thp+6H75fprRPwyYHNDKTQYDTFrLjKMREAKyo
25UlBViYbJqAKLBihY+y5OQWvn1mGVgre2mU7Zj6knfMJpqD1RxeSSI9Inrps8Id
mPV86PGml8wv/PlO6HEOKc9scFNtlwu2pV5TmQprpyR+N0roz9yhi5wt+q+cbDcK
9EscsDeOIiDVuqkuGd5cU5L+2hnPzrXErC9DAbRi+2RU2zbiOECCIHvHn4ebugBP
/F0CfjJijaJCmlpz6K8lHkLAHUpk1j07Z1wpHdqEDLA4vRhX6M3pY8tsHIF0w11P
wKBvI28WaCuoWZsaiKUKxdQG/D2FwwguLW1DpQCkptr+dnSj5cx0GkfKLgLP78rR
RtWi+4oVNJTXtpe0kgniUCvHgpEELnTimhRZVVncDkS3s3+YaD4PN/j3KiF+J+KU
gUZY8EWixnp+7YBa4nuD946fASWT0M0/5jTrGe3n5zU7qIIBTS7inzKg2LPNenrd
R5GXeN1T8toPARPGSBaq/dmKkjNeZ44Y7APvnRqlXA8r0wKuNcKQoBxmRzZdnBap
DEf3DNZ7A5GlAyG0SHUVOLd98n17PB9wBh4WGEHRXIjDDnHTrmENhLZsVvxqV6YA
IU/fqnw7yctbg6NgrIlFqn2JIeok0Zud0BwvUnCn/jfKkLgOVklrn9+42Pp30fan
KzVW9zpwAfRHA7eFwWZrIfpNAkyGjoyVXBx+Av9OXHdRZomOOnorJ6aHZmJTPcjY
yG5vT7kgCrFlly9VKhApDIauqbrExIbwDldV0Jmhw8DV8/fwdry364gEBIosUiJU
1X1Sa753wfW6x45o4u9cjDn6Cjh0qVCsaKo0SgXj2AGnjIDitdzkiEIpBVj7eVm9
GwL9KX21cuDBcjGdPkWjbHzOmuWR63AocC63K2WhJ3ym7bMIPkqnzaGguKgJVuoS
5hE7g0qKRBwrm9hPJ54HlXfsRtfc93pChA9LLu+cTY+InZ+42wCJ08E9RdHCktS+
OUVdProG2OK0I6N6zh74sX4gQTT6E/51RM8C/TvHdMu6T4d9NNNxYu3L+ZdYZAsy
5PTzbFpz/7ZH88p4QanxhrRxyqeUYbOrhVl3MD6VsHRaqIWafcMqjKw4jG8/IsX9
C91HwHZ35iXX5o4qixv5gC3nLd2JF/l1apszph/OYA6n9MwUzZrND04PyK1tGVNB
1QrzHUUm6/07hJ4oYV3lLp9XGldgxtY3z9c0MapHnDYNrSzsHfjBA1sY9c/eBsAA
+oj02MGd1xyzY13coecIfaRZEZw2HcwK5iXtdGxVl07GY2Jmk7MrLJsL4h87AIyI
/vDPeidyr14azJftNek1SYPEbR22Qutgsj6MVlSdhAuq5aVie9UPBwSiapCEuGoV
n2JVY7/T51kzHUFR4OSLDh88n+mhmy/NCrnAyAhy327hZoOAzHWzKEjKHkv2+bVu
BjHHgzTugD9OcNr0Rp5LA10DlV2ynen9W181rkibP7gf/csP9M8sm3z4AMdTsSog
Mjej3H3N4h/PCnAbF/Zy5c+2reVaI5HwLKwUWVjFkot9BjVQuoaw3ztybA5yPjwc
HfBJIAevgV5soG8WlUlJC13+mqEJhErG13b9IzrbLbNLrC1NJBLSAS6jjPLeaJ6S
YRXaXQhipEiWnwyE2zP6TgC5pv4K2HwqghBt3PnjlSkHnv114oAdgSaejt+zgGpr
o2Wp5fNLsiHeaVpKfH/UXYa6+KzL9xu0VJjj5X7VNkiKcBSHlrAIUlXyrSScOVrB
UI4S9x0Qe/xUGx7oImWAlqRq9nr1Q/hKZ9ZaEBXKonIXWVWUz9P9V62oYrrKSpgp
87v1ucdbbFZoczMWUYdfheX+R+5BN/myuXA4wWBte3lEBqL2oYfS6pgCU2ICcO5t
Emsd2muhZO06qeeky5ivq0/AD9sS0POvYBziMR0ELBOuO8kyzljIl4h71zywOiaZ
hTejZGUiPawfA9Gal2Uu01/gY80VUgjHfp8xz1IUXiebu4ZDQJX2C4upEgzjYxbI
vP9ad7CcDSzsOFB0lI5fhjmEuKpC+id7jTXe5tZOsI33tJZea09zUyxkkMsCzuX5
bpM7K0MLHKKFpDyGiE5piFtdQ8JsrMiqYEzuVJzkxvhlUp84rmnQXWmGVqAh0sTs
iY+FO5AZkjoZOUE0pTMSi7hvu/9JAMiOm35939sSLbhRrJN8i/HLwOz1Ga6o0lEo
GtUT0Sr0VWXxo4O/D80nH1HUVeetJLd3h8WG+lFhH7F2wtSbaUa9P36LIXtRYibk
uiPPDwyzPqnHoA2rHCKwTtrc7phcwxs5sUYw0Aqa9DqP7TkLhs3T5XViDzR4ubeT
406GkVXHvocnC3LBJncAgzCUjAhkr6EENM4tdUMzJpgzf+EfoFRgwqyF3uT3uwJq
END9p5tdXLHOiGjnIgUZZwR7ZiKrK9ed285EftroeUw5GmMYslC2IkoZX2245x4G
Ou4WT/i+nzn+sL1kqsFm47kOXhbPZnK9XPGHOJts9OK6CkhWS22e4D7kVLslZsjk
gDvDhUAtV4CY5NW3tOUYuhcKzorIlIAO2MDUuDUOyE1NhGH3GCJ9w0CMtF1p08tg
jWNZpU9DPdQUA9CVq/WLs4zgiRodAyQDcOsfj5YoxW0Jqcmo9D8MmYcOlozMRGBH
ZIcgTc/+GxyhwEda5MhqKYMoq01X3ojxNPXrIjToIfEckrm0KcF2mxV6SALjc5I8
DXxxqI/FUTzS8VQML/g1Xr0cp1cQ6ueJ4+9jYDG4oXnCthttuaan9orho8IP2Wgj
gJTwcFQqSa3NX0zKr4nButJaP1BO23C1AFMTBvbTpoo5TcXob9/z26IVq4npYV+T
+1M5iY/23K2fSG+73eB5b2J3NswOxh3S3fIuSUEFhRWzA11hYEqRHWHDxgr8HO7G
B2TznPk5yY7Ryxc9CgEopOpvqYyPiJ6FvVIvYa0/R6BsgwoK9lXl0ASDoAKi+OMT
EUSqlit9J0XHeDmF7n4y6l/tYWIQchKrJqNxLoc8eJwoPlz86FnkU4/8PV2lX9x4
K2T49wCW/zSWAhgSSiXkXppvvvTPQBIwF25I7ripWLxkjZ7ULEsfIpgrJh156SKb
I1lrkXVhjRuXpCZoic+yWzTaCfy/GtmGNn17bUi6pxW783hYiAfRkGzw9M+AttIK
UaV2lFOd6AtrYIssyJYXNIXKOlmAb1xsveeYg0ya7AhI7X6BKgouL/k+fquijRPI
2AvJTPiibmgPMzTKalwIiylgwiV81OWt5s85Ibv49wHBnnrjvkhHNmR0pMrZvtKs
SLWT6JrDIevwUZyjhSQPvVYiNbl7f8gaVs0s2R23Awa7Isk0+dDV+ge6amOEhxBX
EVSQzFZc1PuungSLe+LVvWETUl3azW5AZ5tzV6si2N1gpqKfepopM4y2d+NzQ+4u
Z7NcnzPfMDb33lhyL4ZuYYtF01Hl5nRRxNA4lodz2YN4Pn5SNsbXOuXrV3u/ouoo
xnHvBIwLzdM0ErDFR79sBAsdPgmFw8IT6Lf9ogsF/QEpS8ItrcLpLYcfizR2xad2
uEh8mmf7duCoI5c+TGk/scycugKHmdAi5xdSWpWyHJx4b8RAk0M45vYgR250zybV
5e65a+7rauqSPFRrvOP0ECpiLHWd91lxt/gDuu7GbxsR/N/lWmPnmCHAQGVBp9yB
1QJm7IM84z0QQ0cBQSxVOkDCE3uShisVgnSTujlI0FQ7NE9d2nOav36CpTCnhhg+
6j/Ap0o16vIAaKGtwZfLGKzfStZs0GN0dhaRN4IAbWWE9npiTYyo6cc4HM7fxAY4
zZHb2aLGOihEl4vrFjZk2oGA8vbxYgtc5pIW36/vMuL0zZCZohXLK6IYqPncuHgL
hZFP3u5vYkup3hFKlLSOAvzWhsfl75iU0jzmsbJDWFVHP94CVq54Ac0xFJHr75Zs
L1TU44tU17XKnAysiD6oRpu3HXI5Hr96H+VSAt5TBm9sE7O8RZsNG4A6wFszWr7i
/pYdoWw0BKt4DDkOv1VvKeiQG376it8K+miDW7cK/tIhdOxH2Gdydrye04Lx7Nqw
VCgwuQKg6MTXxT9Nk0y3S5fEWjm8i671vAFopPI07AByVbzUy2kGl9G30r7TbUGA
c2QQMduad5HYG+MxdP0yJ+Ip1bzgIXii0fBRlkXDCFGaUMs/sNYQ2RruXh4hOke2
V85LHqSKi0hbFW0ip3d36rI1nNVwG9Cwj1ASRz3Q1F1Rw9gw2Toy1LCgwP09Rph5
lhupNmfWEDwPpYM0G3tQjDX6f1PCmA3yoE1hhp1eAsoQJK3Uz+ndI0m7tiwqU0Ud
e/YlPgWtB7XWOxEBAEKk8ezImtjZ0hLgHpKTSrX1OD/wUh3ArEa1Qi8I1De17+GD
H7Jvjp+fNTkPmAz9OP2lrXe6OUf9NsNc/qx06j+j2rThFzkLSQQvf2yNzFZepKrd
xZWwEiMIy787S+fOM/8D/f/RTKfhcx0PIaVRdq48GcNDVBonz+j0oVyrkG/+o2zM
ApaxcY3y5cqiQEEjqm3NIVTLtVeXRgH4STddcEtAYtcR8/SLQBy18vyA/Ae8P6Qd
XUE0qGv7na3T12t3xik/HiMoThttiVjBmuxu/DeVOwOYQyQH0boTIMDkDgjxCllJ
0YvFeHmKA+WddGHFOJT2zLZKge+CRCAL+X3JVqsYBOicO4eupznbV5O11N5bi9gu
Nyfzc7MM8cmYI2FnVzOVbroPC5J90WWap500aN+UZ4RaPUzkdZ+wTeWgTrd9sMRK
oUrY5/GcUpB23HvMy4NwzU4+s5OXktSLexBq/3O3zIVYsJddj/+YHY0mFMULAppi
yuHwB8mUx1tnrZSsRPzLKbtYfEz7bDCszigSN+/Te9yLJvsZy3w3z+mgY5tjGA1b
7rqI0E+XEYCLjFkkev3RNAdIxvXZYeAzkW53rI/y44xWDJ1o7hPsdMW/qM/kkf7J
swet/hurIqgQEDO6m+tJvBvpt13SiNOaJbp+FStlHsY6einFzsg4kX7hGecBD46w
KmDp4YTw620ykG73RL0NdHP4pI8PlNzSCH25+J6+M0XhtxSIeg5pOVVbN/elL20M
qSbRp28AgBjCmN22j86W8qExrBBypjiLh5pRvQj8vAIfcV6gPPYQ2A8zj6RKf3Di
qZtheCvjziSJboWpJG4GVKQaOsM/VpjstJwgVPmFcdRaoJnyG+E6YPivKBqJAln9
0UT7R/C6GoiUr1D3WsnR31Jjs8kIDO/SveO50NAFSx/w86KQFeru84qZrvmIuUcW
e+obYvyJWbEwlvszdT7EZibVytZ2FFUr9jbOlEP9H8CPpXF5n5Mp/tbz8luOhykZ
+LdAXNc0Zn9RlqECjQ4SGrhj7iQz9DuBLwQBLP7ncPkQEiRk/brOXKxOrt4s60Dp
jArRsElHL6Ak9JABX7+3NjM2q2b2oXwm1vtPmdYlrLjq1ix+GclSKXSgWpbiL5Vq
Stu2ZRsyLTnOgjsO6QYNBKLoZj9olq46Bsw6AdCgMQ/6CMHbdw1EvBXoEXd2ogop
8+1UlcVIgvKNEhu+KuBGXK1MEf1FL1SCKXFbBmV133iaxo2INZihAqbYFR4547UK
MZprt6yZjTKwmaC4TwVmLIRvvCPCLadhbUGEVQpkvko7ScUll3M2EKwZB1D92mUG
4KzHM1TPDucDST6BKdrTeszU0+QLFfnWTCTNezk0zhLU5OA9hz8Ph0ym+jNE6l/p
NfRu+fwQkOZHndB5YFd4LvQt3ZBHx/RIAyzoMln5P7jw3VEc39YsjgUnyVevh3ro
8HismgvoxAWVP+sXlVa1j+jysxEYtQ9piEep1ICp6IS4mZohvtI6q2iE967xgMDM
gj+sQrvbLfT2u13gWhGrkiwfCvwQ2uo2cjP8h9r1ygFy9i8QZJ9LHxb4JRW5Fhtf
a6LdUVQczOJbriyW/Uh7kPZbcKxedsNfnxyNjV9iC1E30kf9ZyLkZ632WyIc7p8s
N/pdiGCQV8eyvMYX7CT5OecjaqWaX07NEIYGE2qbelmdKOb+i0bWB0y5dwfbb5lb
zY6GJBC+iphjMwkWu1WUXua0wlTnOVgJgu3ots4FC8ztE/DNLUO+9NkvJLVwNa6F
RalHRKKJbtgaKCi/5b7K2bHL4aIMXCfj61sqpf3mCLLdqZeb5a1xOk1ENiVpIS1N
fh1yFBeXfBKT7mNxy2yZRrUEK5Cqtz8T1yiHj00uR1N4+fVQyiZLjtgATHTrqgi9
5ZDJoSEC1FZxqbVikDtWPhnEpB39+bARUqFWtojf4WiuU3SZS+JX+wVB0tP1ABH8
QdNfVPK/dGGwDPycEmCdHlx2KBB2XPZj56YEINHHmGwck+6C8oX7JviW4/H70d+F
dHrwMkChpXPEbJkX/ht/i5f/7ScEDgflZh6E0iJVBOXJGYz+rXGYdoUYNWbXFGmP
kVfwmULCD2NqEbeTgPZbubiJi0zDEgJpj+QvgxN7r2B2v1OGbAwmy9ZWqDC9HCnj
2Q8zwuqIFAgJtMmxgDEIElVvzMnl7jj+GPABc1uc7DOcVcTsyTjb0jpleLzIjc8R
oMXJmGg+WgEe7IOT7gPmA/qVN2QU0hsBfvhlt/zZPjWzwmaxEd5xPFjYW+vjv1lE
GKKkkEt85MoU3uyXYa2KZMEyZzV2riS324NmPKCiXA/iBuWkmaJ8itK+3IhF/kv6
IONsoZP3IIDZY+sV5/juE94s00XWIM/d5wEG3yRDncPa/36n/1UXO0DwUooEefJK
vWsMMVFW5EwiAvmFG5Llx1Th4ZpPUj9rZSIjNKfz5cdlRJ/qXyYFKnc+TvfxjVH9
69oEJSo9a9khyid7XH3k4BpZyprkzaVYRy8LMIAf2thwJuwfJOuqJmSG7udwRRZu
bOQTdQjJelkxL6qKhEMHKWEXPocVBFR63nhqUUscfGR4Vc44UunKZGOtMp/yYyzk
4izIrvNzT1VVM0tc0gU1tEFF0sv5qEq7RiKUXU0a8FOtCMCNciNp/CsKp2V7+F6h
WCqwIJw6f9xu/yzHsVmDezNCZmLOu/rMmIvf+0f7GpCXUvsaFgUOW6stNEQAkj75
FAcoCEhPgTwgBy8tYGwKLNg6kF+IUuGEhv+CJLUnpEtkLWQ0zFIieOYrhm2L4xXc
5HPLa1433NxcFBgSfUQvJBW92VUW7rPbY1cCJfeKlJC0HxQI2mQFt/BFdQK8ykz8
IFQYFCDmwqtPWWJCZ6lr0HTOOHLRSvIVpPOiu2eGESX8EPBBmAE9I91fz0Y2LyKa
oNZiyhp9x6jyc66FfP0rkJNhrCVwyBOCgkpopsKlzzTMhOdIl5UdXFiLpBD2DxFp
3Nb/B+AgBtOd75t+il3GYHfvdkLuqBvTK90E11WxZU1BY4e4La+0DbuPbhlZbcMT
1E/yveeo+LrJA/l/Bs9b1LRamQGnI+b1KXjRm5eTHfCayDeOMUo1oniualANJExG
67TmB9rtXin6Uaw3WbilmGZ3/s0qXM5Nzuf5KsxbEyu1a4DzyJg0oSeRsOeb2FPb
ud2dJ/jRVdXERZ2KMu5cUEHLdi2s1x94W5Z6cwSDur1FG2CcpImBOvSmm5vT8U2B
D4zF8dbE9rH2YYXVJm23r++P4aFT/z1Ury6xDlmuMnoSFbdWcootwiY24CymjUS3
gN5RpGX9mJ0GyCkO6GbA0aVzAodrSJjxniF+87LmArvEVkfWgeSAtW8VzBU1Dwzz
jNC8jEpu9Xt4Mg0TKYZBnWxqvPreHgFeShLLoB3HMqfmHhFlMTfCB2cQ2CEf8aY0
tPbPxZIbu574fzC+SRyHvP1NxkwjyebKdMVSYvhDvTOcODjoQsEpm3mJ87ZrBShC
lUgnpJT7NrjkcDojorkx5F9YAGW6KsA6Fu9waWDHiSnlGcWgS7vD/XJ/Pj4lHmIr
Icm+atM7j6/nldqOx2AikR+HZAMRkTFrq4ciPrMINoVTf1jQBDcjZ7/AYDtXgS+Q
Y+PSB4ZlEZNPQLnQbMAbHjleSsdKGItw5odDv6VCtqLf/oqN7FhcyYYSJn+mLsbt
N+CB/ZV/xzw4Sgj891T6httgPjiQhmbY/gJgHX7hEwtRG9gm1JEkK/y434E69vL8
e28mPK0D8l/AhfkubjWuqv0iz3P/UBeV8MMBE8mrXgPjQa2PcE+gxKVuwNdCseYl
UdVKeTWxzXKklxa+IMDMdkFIuqy3r+wuIP83OYBwwUMQP6BzcRcaCR/omFAcK56u
B5qF8BodaDi9uszGl5Pu3NVhxy+iqdYXMT+8vtra90M5M5yhqTvSuIdwnAqk+LZw
GMGDtcL/Akv7RCtCttcWsXoribU4i7mRpNxppkN6Rt0qIZNTLl+o2V6+BmiEzxxr
eOAkiZnwRM7ilS8qIOPMExFBiGy+oOxWZnxe+bC9s8VaZfBYpF1rzYB0x5IQWHF7
h8AqTW3Wisw+OUHkwFLrHagQeGS+fttDy0nG62ARRvHt04AnzA5RxbxDrfb++Wny
T1t81tnzuDHAva9ZTMCdsRr1dv7oEe4RVETj6jGHrvwJp3parn05mLLBgccVJTmE
giRhbMahdVuXvnpIkhnUM9nqzHzsDRk0G0gKGz7Hmyq1CnFeZHIDXRVIcoRtlcV3
8FdBoBEeKbloODNtRdEGi0M0stC2yGuWIrVjuPJ5f6l4XuChzvKvpeBsDtpY60Kx
kCe0ueXC5AESHoxwdP+itSpw3s1jf6TWd8qlIG0w4IavodjUtoTSHGf0279Xjk9d
1E4WuB5lNEH8FcKBpa7vQ8U1OK6b9yS/3oSP0VFWRcTmTviUwMVJet5eyi7XPiNQ
AvH8nln9jOKI49iU/16vw7JZgvZt31javGhqKwikCpBlSvH02UGjby4isSKTELha
7T33p9bbUCSUn7tPluVTH+9/0/DqwmxikZrKdAG/uRAxo+BzexBab+EWivHxe7Ai
qO5Xp5a8MinDelkvqQ1w5yIyNf3E8z/+pL//x4mvhy54lB4b+T5nMKhwAUGOJ/xI
XvYN7j2s+Y9AxJMIVEvANOYr3EdDq3gdydhsgM/E5GRs/x68InNV/G33fATEtkn0
EDSxGsdu1gsFg07M0W2pXkjJKbZ8FNjMFRauD6iqSmXVNyoKXXsjLx48vsNDGQrx
dpE5/pHX4vcQHWEfSPPlVRSR6mtgyfTvpprbXAZP4y+kR/m8mkeAD3ssm8Jx5D+/
Wn2nHBcBlbhPrD7BDAby8f+glE7iqUnCrv65U5rUnhZBjNfnP1re8s9DIVN/Bah1
bQC1AGR8sKxxGA+93xJ3Kcg6u/qicbM34VnrSx3iVuM0aeeztsc7oy0kNCcsnwsX
VzpGFNUdwSE4/wtjS8jisV9X6P+yMvJasLhFk4BpKrRWU0AbgJ/SAP3KXrILQmDW
jYOG/ahhCtYKl2xgeK0JWEMwtyltb0QPVI24+HCF2iXwnH7ybmc5AayISx2I1I2X
cg/hO3oOle2CJ1qQtQMbnQHV+tXuq0gouA0072qPNQntQStfvO2Le2TUkOFpHvZM
gtcxUe3q51thd6gG4LhiMcrBAHK4bDjCCWSzNT2BbTib5DToWlBAiBSLTixK70vl
9rgY/iMNU1MDmChfPcGG+Cu9VMaMMI1TXS2alHJ2chL+ZDrK6FfHC/1epPr7P6+v
7XELd6uzFoz7S1LUe6CxH8jD795sE0GLjnFJ8imodDTLA8eiiRr4e3Dw+KzJzA2J
xNXotc5NBYqwc1n//2zodZ1llNTha6N0cyleZRNkULgyhRMl/MA33WZ7krKkJp2D
WBLy2NvoqCs27oldSK+RngVHaQQrM6FiOWRtnPMB9PZp7zcC8+jYpGrqDn040JKW
XB4jMQS/8vA8axpoBfzPHqdjOqS4gqxHRABSeV2o85YfnJVlPyYrTlpXbX6P7Pfa
WF8PCdb+e/aVgk37hmpKCCVL89laFWTtpriLaujmm96MH756BlIpPN7DMZ6gHdsa
w14OywsfSA7+CLc6Ebzzkz5KGITfjrv8Np/IMQxon68/tu76JiYvw8MI3rsdmTLo
n1vAIgRfm3SO4lTkIoejwC1Y0uhaSHyuU3E+07BtVSwmpnbF6IXwYkfjLKd/YBTA
AbTh+Tms+2FmYC0UdE85lEd20nNZwPWmTBAEIs8OZMbxAmo4FxgjgMr2gYOpa8WO
6S+drl2+koY6m37f9EVKy6sMVnJXSWqhCQ2+oqI7G1EFa8TwWc1huxQLPBZhgoRT
FXUezQEtWxHivXfXcAgMLdN16y4M7UwXlXOLsFt+Xgq05GeSL2GoR7cjZS3kYL7h
XAloMXkyfQzJWu0qhuUIvuS7UC4BFHwnwnMjWHnkhlM6oYMO+G5nhTRCdLQpXlHx
g6P4x1bPQnb8gSXPFku00muDshXWZSAT0vQplQTkM+9pyCT6ZCrTjrUar3X6Jm7r
RsOvaz1nKAHio2ibWNb1VLRbovRuOUmyOkVY7kExNjizzVoQHL3/nXIRt+IkrjWM
DPlXMg8GD3qd7ZgBXzAKaIXzixalmQTipI6F22aih52dZ7mtsZ+v9h4Fl/XU3loF
4agLodImyC+6n3uBU46+LSpFn1cqou5UATQadKoY1O5SIpHbeKwqW1bMK+2H2kMM
v7aVuXxICRCM+XBmJaAJeb0rb1de316+oz4YnC9Z/7y9aA1/KerA3BJYrTDGU5Mh
Npi3vlhNXeJXegXmYiHZf6xtwo4EdvPtr31odkWa5LIEs65nvJga4FKhpsJHJjZ5
SINIE0EZbnGwCuj33hr23u/OOHY8gBGNtfVlPv3qYjM3uqySu0Tu9hsTMpcB7CPB
if2aNDm/olz6kRKNgtSW7WvEOlyHvQKMVgW2XVadwmjuFjnn6gQHbAXNMqkMmV/a
r7vRmD+6KtHbQU3SgBnwOSPpnj5TAVZUQZBL7o99apDPc+EmEflc887jEihlWnNp
G4j1MgC6u2LoTKaFwpNT/ZAbRA5+CEGiOKvRAYbFnZKGDUm4LN55AmB+h/u4Aoky
+Z8XRHY+EiAtUCXEWISwSvbI3Lz6iVvEbndvxGkW0LCVESbYxK+7YOxq+6qCf6Sd
3xQaPDVSbdyXUe5kiPX7DBC07rwAeyX8rft7OG9q3Hw9aGgfzzAidCMoOCDezyfv
dRXcNEYaCQ5POJndTqo3SgqvU6U4SUGkCyKC2Fqn0y2jlGEB72CTKUjuAtaJ0x1m
ou63ndSJnIUpLpINY6GCCahq7oHFN9rFtn+7Zca+9RHpmwQTqq4sP/OJNkAywTAC
ugjL60ETsVWM+U5l+1OqZHtUt44MpLrwu+/udQkXtCs5YS2TzB01L4yLkrQE4ucB
Qcew7iFrib4rrGBvBJgHvFBSAGkV36tb9UVgR6EAdB6xJTtbOdVdD2WsMEhn0sQ9
ZKRKjE8Bs7DbI9BqLDb5rSAzglJeUH667ma7WJAudbaPmNQojaesoDftSGdbkLkl
Qw9SVozo0bftdhEpZklwRNbVI0VMWr1nOl3zEJcoNGQBIqge5d8IMevu2BhQnkoZ
eyGWwZP10wzoajsIMuzLEdo0hx08IQiLuj9EvWoDYG6WTRpMCvCs4lhpQdgB+eUP
nBCoo8JSw7SWm+rsI63tTSxTrA49Jw2d0lg4rwSJMi9pfgIdrVos21Nu7HkeQfCH
7rhZj7Z6YMmLHxZnmvfMVDWvWvuWZYREn/1zY2yNTmNP+peTcIgH4B6DXPg3zImz
YFw1a1ITK82ZkU8UBx6SVrepd2+l3oxf3WL1zs4GwWuU/RfHSgbxYcmSceOrqLN2
2O3Qd/SaG3lzgRQw8E13l1Z3F/ohp7cfmKqYkQ/LzTEdDS69lnjP6IBUcTcNFDNS
+2ZKlViwaz2r+vjMtA8WsOh2OMtfpWrDkbyr6i++dDdme0MATgpdo5+eeOpEhT07
asR7a3Ti7/t5+hy7Y+ThlBtm2K+Hjzhu4lhSx32Zu62HXZCT0ZVbtACZJMoV/yLq
6WvoUoh0JgxEFtP1oT1LFYCbZJ4/5f3IuVaImKfeedcG+H0Q+fFXoT3/GRSiM9xF
btwuVXpzmMN2zJiLDAKuPN6nhEs6AzDVTTCIc/ZSpeH7AYwtHFG9PDp63EHrYzeH
1JbqENa5olBwizv1OonkpLtke+WLB6EEe7OIdJRVqWdLrA8ckW6h0BzL7WAAwl+e
JRLxcmzNclzr3vgGO1mBMjOyg9I24IjCBGkstzKz/+xZWO7Rj+Myc0EDv4sTvZsP
ZZrSZecsD4vZx16OXoa2p9SePx0Ufz3cuvZ9JhusuYsZX7ct80FguzPpTHZCTXMj
/ARXnsqqr/15l0POnV+6f6HjNJS3+xEJbM42p9Ul6MBHdIRxXKV2P6vmTKByUJQH
TEcE3oguCSWTcGoHSWzmhRVlSfVBoyNLaC3BFqhIsJqQmS5OqH/AyfzN5agSboOu
uCRx311VTABkLQDt7a8vq8rABnm91ff+sLlRvGNMxpU3Ri8LbVMPWVxLWKUUwKEE
RJb1j1WyGZz/voN74EYpMcvtRKSlrMGd/qFc5nPQVgHRMEtlYtlQnSGwxmZbJiN6
hPbdKVluWCtLaZSfK2CYXtul6tfA4HYT09vod3f5ByChCS/C3BZtgQjK4EMRopax
Lpr9jIweb/4QcegIjwBdJZ0h2uVAs2s2yANTSTPh1g5XUvJ1Zb7lA6ZCZyIQ/Cms
+fwVPd6N5P+ItVlILlBF16yCTNzNnTN5qgtt9n5CVZQTROm6Obl7Vh37ksgOY9tw
N55xm7lWc66fHElTcxVoxpbjpZTRwK5AErg6jyAADBauTQO7WHg0Tb+9aEPXoFay
vzeuf6xoAkdmgvxX1oK4e7RCFHaQu9WqCZQ7MPPya42xRJZtd/FkXzS7Mab+6AQv
ScYlra0q5dVUpBzi91kw2pIhquw0USfRdb87PkBI/ubRp0lxTez69EsjgRzmtmRi
7Ud2HFq/Hu4nI5gKSRgJW/YHfgRJcUGB1WC7cqdMWOdXDpMPQN0C2UFBCVL+d9kK
HYWyWbyrlXFKF3T1/CA2/qZx7h4gkJSewjHKuCp0oikjnGKTtviOx+aVjVZi1wrp
tyDZVGFey+2PwtW2L/jYrBJduJfZj9wTYQ8c+f5VGcIa/8vuqLDbboaj/r4dmNBs
jL/LJQwi+Hp8eaXU1VfLitwuxr4f8s0dIPhdc3oosVfcfDo4W+a97PukzxAF7QMl
rxraCYF434uDTARugPaiXu03UUd1kBB+kXxvd/npg1bjjbpTB97i14giUj03uY1y
pgFrLE7X21jvq4cXcQ2/MtElQQ2irYuMMYPHsnud7SvmHGTp5m97FudU0Rj1LwYJ
1oi7qsiGpsop/6BxSg6+ZvyOp/oY0+fHv5djS1Y7mN7MC+HmWMcLMKEStPae18Jm
be8lYpctdAr0cxttaLjefoZceEXSwRxr/vlBXP9P/0D9hGWKW790y2F6Kx37wT/j
6Z5AzXlYweOdUNjowdqhEXPl6ykuxHumGfcxX2MHAaT5lt0uGgcVSI/mXRpIDsCZ
rkh6J/8hS3Yj8r+hX+GyXxZ7gBek/0KGzcVDhkR5a3bHsm0TkcCLgZCKVgE5zGxO
47IRhw4qk/rBdPBYCI+oFxwG7Nt0o5wBrKIV4pF1EsZQyK+4orUXy1TTymWv5gVs
IATYcTjWJJ+zlY4yuBqepgPL3Vabrn7LOg4Zy4oGsvGdpy39BIrX4w6FNjfxdVOJ
Nyq9IavcJxR1PsxNwGFkRwSEKQ/hYqib5p1i7KlDwDynbrKgt6gcx/CtMuvoqFrj
axZWUqajn+m9cwiuWY6F5q30JHLnIAqOH8TQhMHoDbCcC0XcDCVdVz7ZkSNnMDAS
vT+0Ay+DOHAyLGJbjNJB9qhIFQnMJD60QXo5IFuyjLvOw6PvmA+95UQf1SmpNpPp
1F+qPtuVuQK6GTkOhaQj/NdVQ7DViYIdczOGqMxmTanejrLQmytYbwZUr93tg/6S
SVY3Ze9InKytUuIK2YvH73DYt/cfT40bDssYyH7k67397bxOC5dNRs0uJnuN6WO7
oa6il3aVTygR8Sj4o/+KTYc6g4G0tP883eL0dAFjBB9HkBk70EIhORFl6PWBaY02
WvcK/ObwZMt0f4a5Ez3ddvyV0GFc4gPK+/ge6h0RiRtQZE+hzK4UVJ+VccfY+BQ5
Jh7iTXAw9oXPgS1DeR3G0RN3E8poJO85aJI9bmlphueep4VJkCSPKI3dVsrHQKCR
xvXeBC792knFQAUZmpFOMnvZ31tcmgPvmiqxRoXN9PS9/T3arVrbDoxq0zQHTc4Y
fEO0C2BY2sjHQfHoJl5zfLZunkqYuSix/5q/grzlB1rddC9NBjQZt7DnZFib/RV6
fM6EK0mpeVZv/hAx7OKSJcmwdnw3kSXH57ClRlyK3jx8GTZzv9dDTnMVvh4G1FmU
sTzqonp/YhtWzGGc1ICZ2lek1QGbFSuQoEjA7RRRZT8GJoK11n4q6+1nOxZAhX7G
MKRFpVDxt8zvHW+tGBdoLwEXwAwH/2BAY1XzMxJTdq83t5QnE2qTiFdhx2y/8fIr
IA1jjwAMX96ZtxgorbuOouEWJQzu/k52ntlnEG5yuGASzc9FERmhQUkFCTfWkeXB
eSsokd9yE4n46hqda/fdmX7hyyWScqn83XLsA/Jsp7e1uwWOxPeo5FtsRN36R7Tg
Fc+Gkubiumud7bZYXnHZb/ReAc3y9ltO0yzcXYSNqHsQ9iTFN28rfem/HoJ0/40l
7LUKwz1cUT3ejwH1VyHY/QoYY7Biue3LjXls4iBkh0NhGdTP0gYfG3n7haJmiw4S
T2BLiF7tWcoZzwiToo/UjVunlNbRPTX/EWqApzgZ7ZGagYmQJ5XYfAZ6qoc4PWfs
vZDWZcqRoym7fbdZ0V9Lndok7SAa3q2zGhIWic2EpaY/eUFIIKEp7OeUioJXooU6
Fo8efUVplOwqfv9DwltqJMhpYryJJEMcQhWPF7AeEddRznA3/dPaH4j8F8Ub76Wm
nAia2yeW7g2ltNl4ItkNJfNT1RGDjsj+Xsrhim2A28+TzL/++grg5Je+1XopdIO1
kFbnyq306TX0mcbFvHFSZqLZwkYXCCE3Z34kTk+bLNpwuLRKijXrqvX7Fl1T8xc4
/kIyHO0d/TzkjplBzmFUAdccsUWwmRtkLU5VndWhrLhRYC6Ui+GEgRUNv75bd2nN
fgao53ErgfUekwaXHhx+07wRFbTS0+yb+12erH9bQd7LEqMEgt/iWGZJSROVlAvP
m2lVEirG7QldbgZvGX0FnQ43O/fy1uSd8XbZ2mpJegxDC5Nr5BKLSCNVBP2jRUx1
wUMGhKILWDxEVxWCSbuEhc4hVMH01L2wVyjurwGq4xqDdYVZkfq9BK/hVvPpscDo
4iyiqqQPlzTBfEBiorUcolimIi9q2Ga0E854bv9qGaCxwogSN2h6rK9XQbDxEA8R
Ozt9P2m2oxmhPAYea7NuAPlyj2nZHvXQU2eVwLJKIDSZR39k+C6G4TBnTWCxSJJs
GhCxSon9PNFGdpokBBo+6aF8Qz2uyi4qB9ezqyXte3TnFwxgEIsr5HgTa1feiTHw
4wb3KyhSvx+kVMugI0WTbmjhEFmExjZKqsuwwhUefY2d5m3oslDOEKnKSB+kwSpx
ax0cM5ctVYb8FYJcHXccaUeYz+7/QqRvpbFpuhqtZIUOGiWf6gcOmZv98kDUOx8/
ynjpQJkNY2ZnYJbWFzOaTXiIN0pWqGVQ6zASCD846aukmnWnpkSqWpXJiqbkR2yt
sGwxfjJnrCdkJADgiJflhhXydWalDT1x6emoZ6je/amI2L24aSA9NLSmcs937uqm
TKzCrX8HNXpqO6wyJ+JQc8sEfJdR4jZ/dqXq2tlXTP0EGXjnO/upb1K6W8haMgjW
gs3qg5+tGOBfSe+5SuUihAw0QglF6D6eu0u+2T/rBN8vJhSp/FOXRg1mzBcWsDjQ
yXIEXZNjY9klqsDB1cVv1sXdQ7n6KNVqTMp8CJs7O1CpdeiBH583KY1DgoLjAHB7
Ks/qUFaYyJdwcMG2PZUjIfg17+O6iO0MDqyJ+Xao0VUwb7DbIOkk4/DBwYQMyeNZ
bdAhgTuorbisa03bQN34l6orTwc6+mI31cgHHZDrgmBpOFbI3xojTqT/9JjFlh1x
jAGmxhqnQTn9lNECgtAWkvVf2mTniJoweVLnjzvdEYPr5rF50oEWoZdfYAYa+7Yf
WjEfKSyhtD6DSfvkuWz4Myr7pdbwyXhn3TQMC/K4zIYKulTModaudjDP2aqI8mQU
Gily6VqiZ8IMol7AXl2eiF6Xod/bE4oeglvDFDIiH1Nh7bg7nty3F7nkLtmUeMRN
35/IsFJIvYj5FiMB6BgJt4PuVNc1i/9NTAi4aJGpZnoFfzMP7Rqwt95frpRmfGCS
VRQMdqa2EFRKAzohnVNrd/KqaX/0vLzxVRsJMaQlGb+FRA1E+jYeLHFla8BUIbBu
l9sGJSyJhD7Jk00Ybi6YyyCJ6TyMohYwO/1qRkvj+ueusVPB/3lxGaXoB/aw0JAP
bqQ+Q/I8dYicNhyXWhpkxCP0ZB/7Pq5hXv8tP6JfOdmQ9I7AT73Dmtc9RHG+sCCu
XHbr6HvThJg6vmfGtl/t5GejCRCEe9KUYSWVmOADVE65VbP2HcXICsG+Aw90eYQk
dTfB24Kg9YU/+4d9QevG3VoMqdCDytY4ZIZPIsN0EcfZjym5NjUnxuulZgGjwjgc
ukuGzMcx6XwxOzJFAUdoP63bTZdcdKPuZgOUupqFRf4WBeIMHmkmCqRH9KkDa85e
Jcof9QLhs0kjC1nCr+9GIvGQaGzmou9HWbhZNlb0bTEGKB78fF5b8AU+MzSsI/Mz
mvm1ZHyq0PDEoDjn5obE2azAMUpaWn3jkgiYKCS+Xgy5Q3bcX4HkHxjVZr7O4Pn4
FiG2gXpeSjZ45jMZNrWVwrODEyEd6/ud2hB5+K0itC/8xpZ1/2kKjc7g0eW854gJ
nlL21o0QRbpCZJiifXRra/SemSX+M3VT3O0SGYpqsOiWxVoP3lM+Z7TmSsoQ5E0c
FZ13TSpszpDCEZebddYcsm5FXdi+D0M3n4rU0QYRJj6Td9Fu2VGwPyMG/VFbi7yE
ssV1WVzsvJ8LbRXirzmMF1yzEmSru9zUzhj4Pb7gue1wX1alkkLvCVW/vRsjqBSq
PjsB8w2MrObeN0yZsy447p6dO5TqQGiHLN8gJ9/f6NzmqOs8tIRwdyzcZDF5uFhJ
ObuZ3sahWPiR0nzN6Y9GasS9CDlzxcXUcts5+8q6D563BCK2ZtowDfa2CkYRFMEq
Nj4A78WXnr5/3Evwfqyr9g7mZRaU9BqEclOMBAgp43eySic2PHoRK11E9iCuHE2x
viRkiwu5pe4LXuQV4jlsIeosvR8LmdJUQI8+krSgNxroJmOVCSQNYeiueRPF6GAO
fq0UHO5bC2c0u4dPCKzR2E3/Lo7EWrthRQ1EomzdrLZBjBvnik0ZUrn8dpex7lem
5tG8/4avAOf8qiZC2okczlZwX7c9ms+sNqCMfxhrZyenf8KVw+65oS7mhlUnE+2d
IwaDGqO5e6NnLLnCpKcMbxTrYe9irfFEzpI9llJ1ZXCNz6FfjziIer9SmblZfq1w
zfgzewdut75KCTwr8alViNNfZo4zVwOHSuHYo/rOFuUoyy9ackE3/JmXPEZB2SSV
/LtqRa2B/ZXBOVJ4K0Ew+9y27vaNW/qhgLiFlVwSVfv8P8EbN2/ss4IhJcXUvkXR
59j2YeraBYWuy9iOEiROY2GKISCvNgwhTCwO8UZQX+YZLcJI0PUm/r6ZBF64BwhV
WOaV3q2zEmqzQuyJbsIoZdcqzJ0Hvgl4IxSPFkJG01NAfBuTMji0qHzL/BozlolX
342iunV2sKHgue/ZhmznAEuNyd7TCJFTs3CFg22f59qqWfaEuCFtQrhaeO5DbPnt
V4l/w4k0H507qt4pR+bDXPPn4ycTVEiDGjbS0UAI4BoF5CwHLLXeak1aA9ViDxq3
daqaRI+a6JOCD4D3K4wE5AdHGY8V1q87kwZfCBO31jhAyb3mD/Utuc52vdD8AigB
hECnvGTtITpniE8xeH+yEHNWej1Wk66RTCsHKB/90GaSNIzXNfhA+xDlqJuxIfmW
l7Dr7bhp1m/bbL39ZyhSGb0GI7rF7iCfTT/nYNE97Ia8GFNjBcbYn2dEn6Toxgbc
4Hz2tvEjbMrhSP6uaBzWxL7jLq4+NVJgGboXhoLpAZgnBYnmQc0Q52YbI9+zBczp
3GEyVvjy3IbOPLWxa+vAw6tsTnk5p0Ov+KQ4AzfSsVF4s5GeNk5mfoHsn4S9DfDZ
6MoNBVVRy1l2M/gIfQxU+IEq0Yy+uYnvmQhx8KL2l9eUnPS6K/vIehYOuOQh+ftv
6DEB8kqgV+E/hGRaCb6UnPlpLwuw2SZS+5pwkfmg9N/MWLMs6hnMV7wKBWHD9Wqb
OHH9s6G/CYNx8NwOEbCpjiSVYh+zLAsaCqconFiX6QMeIa1SB/3bwlDEq9wq8DgI
TWPq3QUtpiCnwYPYtnAT291IidDqahUfvVtXTMNTeEXD5ziwi60gWylgsn5Frtwm
G8mecy6ZJh8kCRar75+YUIwbuAW+Lsul1kC3vbMsK0GyGLnrOPEjW+i0LZuyjfaC
12Vekg0SI4HcBfKwaCEfZQ0NDK/FHzAoIPaiVSs7NwNvLIwE5SnePET+ppWae/8Q
ftKEzBoMxp8fl4w8PXmRR9egZeL51EhNEYARgaAvE6Uqmo+5jMOjPk3wCb9nawtq
uAU2tnLx/VaRZtVLb7Ed08CPbZc3L9KYvqEoesavOhQ9shqE/qri4XX00C6ftRzH
NwIz285VDHYRx6MFwhKWfbWjeIH4zBMBFvleSNwhf5uIBmCaYgjYyweKfRji+jNs
X7OGqFPN3aFIWC98coeErniQG2eNmPdo0Kz21BKxPkepdoQH6wV3voDnhRCDK+U6
B4abCR+i51gjIqTwemCs/7YR79izYn+j3LBZvG4KbNu4G6Mj90qqqcD2Hc/wmQ1p
cubFo97A/Dr/E4Rq5hCAZ+117B8oYlWK3Qck4bDx30BuBIHX0+nCQwxpcCqT9YJh
YXfVe8ZFy3Nd1P47IF7iEcN8XzD8drlG6GzFDpA8vwDJOOwzg0b4vtkO058v5DxB
bflz71dFcu8BwaJvw+h3ITtVNce2NLFU00cGuX4AmKe9YO8GrdVpyC55VlaobDSX
DERMXYrbvL9vDdBcwoH/PnFq0akylEyfm9s9mVDpLX+ELNJImKjLRqO4eBm+NNNw
OtjXKgucDTyRxDQg/YfxK2yA7zK32P6Iz4lcRNrtDbRN6DwjcPYwdQThFvE08Ew4
608GKx8PqE9KWT0oWglyZu1VnPLzORdG54bpJO9jFymSrmcYd7sLBAwd2vGy7IME
fcCGmeFE3Qm+SvPQV2w2FXdd4ji9sYYvcuTOlE4RrrXw+oN8cLyfY4p4HmzAT/Y3
fPl1Spe0MCp/LwV8BDuRLTJA++B7o8lDvtk5ote2Zm6zwsCGDKUYhXfPJBcxW6Nr
5R0IdkpkuEbht0ehN522aiZljquThCHs93+pVIyf18aqwUenmsaPmvDhdTPULJUR
9c5cB6BP2xx3F701jeRySDoztP6NkyqR07d963ZrTJ42Le+dZj6VAEG4e++Fdg1r
NRqAchFwzAqs7IVW8FmjxaOqE9g1OY7meLNkATgFDLXeJM/xc30besBrI80GH9Vp
sF4eV3oSNlfyfC6Az0NnslQc7Ms9Gw12IQKFhTUve4jAF90MPbktsh4mVFtYqfv7
8Guu2yCOrzUfvsXQWXKa1s8rwVjmrC60x2yi1xWZ3Bi8PRcZtBKh4PoVGWTmZ0/S
lx5q6ep5ML3y38GbfRpzcy4xYa435nuLbWWM+AZESxR2Hkf576CRhYG4YxNpouhF
2RS0DL2qoJ8FHZEU37ykkz3pMriGqwQwHPi2JlOpIqhJORUNrZw/nXSni91OomcU
6zhTrLVhqE4Ew33GbN+0Ksme+VeL/6Fxvcg4LUNN9HgM3KlWfwDN05DegKkyNPzJ
j55VS1ULycKj5dDl2BxleQqF9xFf1ZsxPnSYSm7TUJipYakmpuaa64BLyMw2lFyO
W139876p+C6oyWSO+MiNGrrrYnlkc3zibfdqHq6R0CUK+i21KlcETv6T8m1urrvt
VjYsZQ3YH/blmmOYDMActgNDtEA5qENxMCB3QAzuDPYXKSqfE2pX1RK9fPvlMlHf
U520Sl057BAaeIGvAN2dp6O0g8y/OUFkix0NHb7zntj2YbMbq0Jape+eLq5IE9Xv
PVsF0jtWl49xrwdhmFKXFXc+gPDZ0X67Lx14cw7qtFQmZLXV/Vq/6GdWCNbZyuxT
6uha6ENVtDCOdiDwX1Ezd06Q5v5LoTVsBCgBvrhH+2lkF9N4ZnAZJGB7IGZgUk3n
CgGxyLNRxJJV6z/L0rL12CLkAHMGnOjBb95njc1k1hRqCh5xZY4YJK5zu3Llb/U2
eEB8TeRFx3OVsryvvxiXMMGgKAchRCb9HMkxlraEAjLA24wLUBBFP0F8e+gQb/52
6w10Ljqk0iOn5r7Kw+6ZPI/NC/zoyogGklF+b5YbPqPVi0DILYEbgBAX/9OwCwPa
+3PnhAlkY+leddP+Sappym4cIPhP7LzsEQZe3tbki4M3a06Blkid7zSNL2ha9Ugx
8RfCQYQztgN4KPLnq3cvhzbA0fsrJisV5r3S+d6dt2s1w/0blXA6UrK+7oueeZGF
sSmUbKXLsATNCA/Ev5EM/tQ2PNb99CdkkcPTlCcg+ANd9b+u4KyQjs28+Nrkju6A
a1b/92qHPVwGZU8WzqD2Qqd1NcpfcW2OvaSIwW1YpnnOoUBUXJwVyJVVFemmJD1W
vcbCZdFP6FGfpsYqBIf9m7eeZXPgnPmV7e6Oc8GNfTTX6a7wkfjjHRjl4vBiOFyK
w/VfA3SVW2FZHRfj76jCj7kpavJP8Z6Ct7Q5lubPsOI/7K4L4I/GXW8I3QDxepPZ
cHFS914QFEj3+oliFm6y1DJW3QwgpvaCKcZP1rVKFqOVeIZR6aafWDmG00q0Ahkg
dl8ZJ7+tgau/gVAfDK31pKCGTFuuHZpsx0ZGX/txVIqy8Ws3d9CCWBxZvaTO9sPF
ztOf7K7DSotHQ/w6N+KkIPDKNAw+nYSkEFppRu5NFZF7P1Y00/Hl6Gk5gWqiSOHs
1/jxm2BywoNTWqf/TdmsUD95s3/geORmXzsv3gsiY7dv240ZYyB/F3ZYS81sn5Yo
092NrcPtsDXbpiq5XKBrmdqHu29ClY7NuvXHjAL+ku+5K/UrkV+0JqvjyIsqnrjE
xg2PLkm+vqxiOVWqxgf2YQpJXO0lnbdx/OkcBydDCbQpg1y1jJTVNMEwpN8ssm05
QsRgI7evF5AvlrVT4Dvgf88c4DGbMU40QtoM6IKwcZ+xV/rUwqOwCuktmLP0XL9o
nyxS8HIa8cLKm5W2omD1jdTm4Wozgh4wSzOUpdNeN+Vx8l5F/+/cts+qf2QS3eRL
49qVt9IJJzwoIVdWGJnSo/rrWMFttx757YhxUVX+MF+7wsh7n3IZ2A0z53PzvPtK
EfDMnpXTOkzR+4tKxVJhCD6A78tVW0XOQJT6Uw3rRGVpdus/0F3BeB79b1O0FHSx
pvjS6jePTHzjP+JfSEO6oek5u9nwyyWY13kouIcw5zRbgY1J9Go4SoVJJnyqeKWh
52z4TdlCe1bRto4hXWTF99NWOIBjuJn4uDCHw4Ix+rBn0Sfc/qE+Y5jXE+dnHnDc
7OcdkZcvzZSK/ZWhTYTSqa6fe97c/Q027vE0pEFY7HYEg67NnEuxhZ6Gv13eSZbo
XBQXek+g8SBH9Lzqc+i1Pwz4rpaaxk7hiXwGDe1V9sWVBu/NThLlmgIv3p6DH4Ut
6mHwGIa2Z7gmUeOXzkUPxq33QrcZFYvlHmeHkspHHIlg0oZ3LXlcAufWveqnbGLV
0ViJ0MIZpI4baXfI8X7i6NF+F5KMzUoacF1voVdNXNO/HbD8+811gzQqbGCZ4Hx0
ANVy4gYBQZHlffI0jqyFz08LB0wVTDxa/77LkY1fMZE8cHE7gbFSDcEfZ1nsMzME
PCTYSfBD997cnLzpg3LFamNglwGIRqv3RoxwxYUAn7HVa8L2mCjKJ09kCKDnZadY
vEcn69W3Y3DWO9yGDaOHdz4kpFMlhhKS0EokTLcDKWC+BuZifNnkvZ9Rov8Nfelo
SvcRFcvDcPkvvcDzrZwQLyR89sG8v9v1USvZddIFGvF/8RCNMHnq7w8FZxe8oBRs
mwXjaV2nTM1isdUS0ARzhSiqMY8Yvoc09p6msHDhocGQ0ryjljZzaaDQ++HLo6kc
+tJVzY1NLxTsLmdZJzbn9wbGUeMObqcRMLHESt+ruAGPPb6E6ucWau/OVXzQvSU7
mhCeoFtKt5uttE3LiataDfRLXvonb9qSdr+r5IoZllU20IBqyCko8i5vXhHi4pOP
LydCbdrTQv5DwUIfi+EjfNWRg4kZXMD2z4soKNpFeONHvNXtu0Rzpk3WSrE6QIM5
jCm7KhpfEoofJ5ryFsmkKzbwuBXI2cOGa2CzYuluHkDgrmNsE5tLpbgYe7ALJ7NU
36LtqHaKHjdj6taTtakcEOQRzGlykkPkmnQSSLUTBTIeux3OF2XnXOHcAgTMd9g8
3zMTifaBKn7PCC0e5jsj4CMTzQtSirNooMTzweophFQ642m8aE885oi6QnO/BrKD
7yULy8l3L5nuwfVkicuDwWu1ZrYOGSNVJiphCg8+B6bVmV0ElbeQhYCLnHvvfV01
2Q6yptUZvBSnlzwetsoMYNByCdQC9jgTRIYoFLwXSIA/1OGMnjhztjtf6FPUmpqT
gxQzdaSOrCrb4g7GXfqebYBkrjr1QoQPcNmdLMrY2EYuEZxMTy1QT8B7PQZ85TMD
xBBY6kZ+UvF0hXdnFkIUthk/KcqUM57Tbi2G0YenPNboKBYaxQGl9dxZkfqI1g9y
mGMyD5e4+xbF4f7oF3jGNi/NVKPCN1eA7m33A8FvPbDlutpgfAS67/sbLFvGu1IE
kaBa2AhxI5aFhkrqyhcBuHjVpPFOc0ZZLX41YOKYlSMAteAPGJehzb+gxccinRXe
QHVluBOpv2AySquB9adMKhWcq5XHlVaHFQ+bt38H/2vyHNDyuVj0pxUITrESbq53
R0trSualsPitSsR2cY2wb12uVUq7BrmcNiTVLN/aEo0lQWgUW66hr7ErDhWji+5r
5+gvowr8KUR3fk7VzY15HL6kR+caKVHLJWR228xQ15UYbCrMQQK92p5Qz2rTm975
g9/BOwVXfsd5wK1g6mQw3dRlXOp+EwuZQe8xdGi+/d83hOHvhtW312yh0+zhqgwH
0X91uu0yiKbQdcxsCIMlXJ+B1oAvc+2mrH3FI+B5gXfcKvR2CDzOBYjHByA+YS/d
CzTx6h87+JGvkmxN79aeUBLjJC6ladqR51rGt5/cQqZ19J/iM+YT2XKXEPKxbxoC
EQBqrlsmJImhzK5TeIanC5fd7PQbQpHVPe0a84/oa0Xxhnf3qyBGWsYmTIEG/5DV
8zKJ7dxo9pRFEHZ6w9TYi4ypqgc1iPiXblZoQWAm8s9Oe0e7p2ojkBAVFqIUBLJd
w1b99GrFzhXmcpPSlZS/omWn4NS1T8ZG7LgV4Gmsu2QMHzQB+G1IxFZLKZF6kKrJ
17Pg4V6fn3U5TN1lUryBl5hKWKHCYVVgPv0bLnuDgJw87y6CdtzjgL4DOjwzyqXp
rMkYPjv27Y/CN6j+C08pw2MmJW7GLrXai1g5PlHrjuE2/zkTYwA0WHVyQD55d9uo
8vsmWVV1Ze3dLoJhJWLDSK8pNXP9CQ3D4Ol9L8hH9iBUBo92Ke3ZJhU6dhF//vVY
GAwKS4XgFktmVBXZrUCVE3bdYqbqNmmdVNvzxSZFD2T8fI+fauI/As+C2pdlx7Hb
UR8y0yQttuq7B5fgxgXOFJz7VU2HgJ8iqpLoimv3AHgVbh4YuNJPGmFHRoV5rXUI
lbDx3QvjLaBSZrj2vIedPqBWZs3crYoQaL8YYnZKOU2im7UivxSRf2q0Igo1/cpZ
DH/xNCOfOIQ1PDGDuRC0fpr5X2OsT8Mw/a3xcCds7/wO2LByHjF1sody/3Rg5vnI
EfvBhowc1Om4EkZGv7XYyK+nTJlI587szWFx6+jRkgrGyRal6Ql80fj9AaESEwx0
8XgVqej3P5ahfz57pWEOLsI7R6uQh7dIA8XBHqnUfxnC/ImZ0fg6PFOB55lLeZwV
cacjqnaj3xiS5lk5jF9TbcLdnlgbgEiUbYgU3WHf2wOexXuT7UPx3adOzSotwXda
hTazshvoV0YJepDU6oBoG+ZaM7S8UfJCICldfVd5OFKGg5MqMiFmiaglw7tWzTmY
3KAelKgTKmc77c936fuzdIiq/gd6n5luC74Q7v0K/mF0s88C8kZQCXBQfHAqwjdI
c1wMHV++ix+7LbuNT2A+3ye+xdPAt1ueGQvmZSybya4D5JCfa8XEgxscSAmOyY2P
dbDhVf9otoyQxfwvdXptX2iT6MTcBxnn6COwKYdpuOsNCDXKJ35x7OZcR0oWy/Ic
Nco05okVAp4bo/WfMdCLzzd1PL3rCRPiSCyd/ffrYIZGz9R/5RALWBwg3gmQWhIk
fhfUsJF2fTIoiXcq73amwiXGAL3erLsyzTHeCJlGfsQHFRIW9GbvJnQj069huMJm
9WlgaBjsEFkEm8HJJBLPfNbTsH2bR2RbR2QFf7RDJOsuSoxSxa8JbnrimYIoYqlc
EqloCB8K9S+ohlhBdjOVPK4ilMD5FFeQyWRqTdpwSrsD9ASrZozReBz2FAuW6l6Y
0T88+0xRcBpsySHJhraQVjygt8ASUIE3jiXym31pbvnf7e2lbVO3w+gAgavU1W4k
XyG2UWFiJ63j6cmGwZPi1ZA7vORWYQlZo5poeghKNykX7P7HGV++0QhGFqbNFp0B
voNjnhY6gbI/IOLqV16O4jQu/cmiMG8kVuvTSjRuhyP4WnzotqL1zZZeRGGnXyqj
9E9gFGepMCm367W/X3ERKxwkV/g4/EJ/76lSCQ35UJhh2eQpxMQbR723WPoD7Hd0
8XitTC50TakXKmet9UcF0LQq6WVM40yQyXjrvVmM5tQVVwKb7PV7OSg/5OUxNd8V
AMlgeMrunwpV+G5H47CjYVABwKGUYRdC1uJX5ntHw0OF8n+SAiyRgXKhoIUgfWVG
Khr54Tfnk4tFg2nBDipoEJrpxySml/oPHEo3UTyzDzpWsWvlMzfbAeqKRKRlDkbD
K/K4KrK3xY8ijVAJZycTYZ0Pnl0Vph4cM+kOToAUIcrY2sYShEESbsUY9lAg/Sl8
78NiYto6RcvVyXs8lwB+uEhnncpJYg36ibQK/9TIwskNyndDZvsYCl/Llx1n2cJo
6eCpUl0F149dxiDtcfGdef0De7ef8QBE/b4k852xuAdVInMVsp8IsAxcJM/HCDJ0
K1kKgBIxCZrv3wcVO+4qMqUUFeeTh9is37fgGQVqHo6wtlEzLz3RGyNS/hg42ckW
MJkjnFyisLXhTu0XjdEf8RcKyMfWGecn4+08pZSua1Q2mBjfCoDY+0MGeUJjrVIS
niuaPAjJL+RLtnpWW7x9sO5A56aTrMrpxGpOlFz9F8QIdTdI11C0Ywz5FMiR7Plm
kFzGkm5gsS6MYGwMmc0Pw4Xo14rYMuGf+O2ZkrLfxohyY3wpgMsDFnfPyNZnTMCI
N9550TFdSb7u66qIiJ3Pmq/lWhyZ7sWS6tCmvErJfhvm/hmUki8IB9kZzwvfFdT8
1GEJd7hDAglY3qCcDfCdCQZaKsUVFmtJbWRrBDRSQaa9NZIsRb2oZsS8P4t2K5wm
bI3ioWhuvmp25UUQefsO09f8U4d5w1l9rwiov1GqJKYScBIUb4QLUWdSTOkyRfzT
ESpi8juh78Uc4Zssbb0T48botE3fQw+6JbNrt2wMjjcKj/1YaHIQwylClajMJ+WO
tT3NlNsgdPaggGUpdKGTOqpBY86vAHgHLIKQ9TCNC1jvS2la029hzGZvs5t7Nkgd
fhllaPsj8BxrSVp5AJRK9+25gg2zRO3SXl8MJpdii237vpHSJGN/uCxvrTrZdNZ6
FOcrY1KEMOx5D5G9AUGlUXWR4iQEURuWNanROaudI/K7VSTIq6F9nP2Y7GvY0e+M
XETQuGyYLoIZbmgKaVx0j/7ad9dSatX7SfwOCApEd/RhdZPGuKppFyKrPbI9dshE
9VmgE1tEhtiMrOp5lWNea7+tI0TX3Hxjz3KEj5On/lDMkCSAkSn1j3vmgI36t7nW
BkAGkv4kF7p+xGd8S1NiwQCd2eouS9mWQGidNc5qATgKqeXzzkTsRF/RZhZ6eo+V
QgAmmOBOL8XcMfBI3B2bATuYEnoN262VsTXyZDANzeV0d7xOXL/uC3zdOW8WwCVP
b7QyfftJeMFQT/phJ6C7xiVvgU4KYGhRSRLkMHfJ0dRTGMwR24N4xowGMNSKUQL4
X9VaecRGcl+0vqp7iPWCA59n7deXH2BH5NXJw0zUtxr6zVNdme6VhanmvzOhMzeV
tDdLz3VvT9P/eNwk5NYFL7tzn90xBIqlb6BBIR32AqaW2fBI2+AN1iF2hg4yWQrO
k9TqWXZxzyjZpykFII4ErRO7EWqFc1/LcF/1L6P7SxksKMk8y4+8lHsBeUOy9lIJ
gKo31WGT5ieh52H0ga4lYE7ZAWZdtGqLNPOaDBqsfrarqbdyCu69BE+o+Fdi8He3
IdJlYuWGvbaaGL882Y0lZ2SPk9Rd8g88sFXzDGZq69uNWl17n8y1G9t3w/9Il/0x
W+k+OtjConzR47XxnXQhJFUHx79MLeeHJ+N9t56TkswFUC0Zej0ejCWZ5AsJEqkE
XiChtoMBz3L26wyuz6JuQYHCSOChPNUkbjbyNN0TfXPzC3JzvUFy45NG0MfkHJ2P
diQZ00zGWxUtPgMq3tUo++3VCCebPEB3b10eGhyGtjlBPYezp9J3shuLwy0/zE+4
3LYCST+2ANyCjmcdCVvuYIxBXj/sPj0DUXzPU6uV0EGLL5aPr4m90cNctfi6ZBVK
0N/mjn90ZSLRub42mImzZ7Ci3FiuFPkmXG28719B8fEYH8QC/SLp9RRSgF5tey+t
9+8afzG2qD5EqX0Br2prT1uw3Oh3ReepSx8af/wPV5BXIVe8IvhTOwZ+bpvdAIyh
rwUZT4M7qj1VFDzki7I9spdhTPwrqMYNu3wTkt5q5/EqCJU4kd9lnY9aHfPFpJAk
9voFwWJR/y3xFjXRX/gHmJiB6D4cJQ5r0Jkb/kPYjtx/2th2ACbqD7dYHV3HHm2d
9K8J9MsGLp0b4brhjdr3QoTOTKMvwu4BsY17adknytfag+yIt1DD88vq9eDhIl7A
8DOU48V4PdPZ0otSdXueoqhVqiBfpoZAo3ZrQU/jgaVdrIwtfNb6tdACWD5gMS/F
rOGxInLEPO0S9WYb19G58c20ARr/16j2Kf6+DGkkjLOdvW4z7WM7605j+0+ITYay
zRutvF+R3MVGkLdqpgb5BNaLIGLVFzVE8spXQbAG5+jQYn4W7qCWRq5FU6M1HUtN
H5cCxLmwAbZV7ZT+FAp//vaYscr714Z9J2dLqfQM+ufcD4aXq3W1C3uv9uQkgtDf
wLjSRWWvCQEpGseb9uVNWFDtE8TwMzRRrD/j+Q2HJQNo8pE9DtvwvYE/0f7mCxai
af8ibyGsAfZuwTtFsBa84kZQu3rsuCQdK1xQy2c6VFVTNPwfpzrorEACJmySzRQT
+kS53g/Eod6Wd2vv973rdtFEaBdMCG2JRKvVSSVA66YZt5KBgEDXkbU0USo+solX
aVF8tUaF3CSqo4628uvnQhihPOyyRp9Z0XphWwBwUISMwI8AcHtYnljo3V4h4Tpe
fmMz0bWBF2dUWdDM3JdknCrrZscbm9dQEXvVi8Y+6YHfLUd8V/OpIWLKM4lKIo64
1SMuOGjmyWwgTnUbgQL2bY6yQpUj5jIMvZRuCb73RPQSOCe0w6Re2EQp9D5O4cAH
rQpykt7zLNi6utMvAVO0i/amg7BEQeTvmSv4Qp2RB8OnYcgAoC38XhdVSicUwwEr
nRe6/md3ezx3uL6tmp3s2nzJIyF49fFFJo1PpgQK0PqsDCPtpazGBvAML9ClXLWU
9lVMM9XYbootE+U5sj5A78dP4KT9yqsDhIm+i4w6c4a4nJYteefSlAeLuWpc0t8y
DChRmXCPxbJLA2c4IBInXGVlbNqqZoW2e++qX9SdZKJ2F2G3bIrYHPcNphA/yna9
ecxejWRBybihJZ12ZE3535yEVq9oghlJU8hfEIhyuOnqzhumSe/oL5HyUULoLn2l
2tya2VwTgbQYdIi1DUDGgF5yyf0ZIxmuc2rhaGzPdUIt/rL5vD7METICMifa+l/k
3dW6xMZptHNW13uGcmJhdrDlJa21sqKNmwfactH/lTrNLqoRvcj70Z7pzuY4r4AW
jNa/QVdUf70cn/49giHUMMI05KMOYx+LKe89New+jTCb+HuVvQch6bfQAa81pUZ9
DUOT5SzWQjvx290GH0waGyCQBZ9svqH0lcAbsdhw+4XyZL3uqxMm7mOQn27DWsXW
YYb3l08u3fTbDm17/H+8LtbO+DO9J8ccYYRFbvWq44t/yaoUmiBRPuBrN6V9S2pP
X63iuUwTby+l72IQLaUYmYZLzfuUK1UgwfpsOdJmrFH3OITUJpxtoxMXxTU+OpJM
CaDLfNnFO424CRhoFihVlwV3BpM/ORq8/y9XAqbcBECO/id0GaQz9tg/VfEwcNzc
csq0v8DMBvkYU+INoDJ5KWtNEqM8yOvdZTYzcYMURiS515JBl3Al/8dz2+Afjo/s
nV+uMTmTnQz7IL7De1NCIQW0fAFFMoT9+/olVDvv5MQOifsPa2rywh9HPA2l7fCG
EGUd3WlwJNXxl6QSncymeW4EGGwH6UFVd8o5b1frV+va2eSvBvn9lsp3EGzyTQC9
X/McxXD43DWQIc+aSKtMT/XpvWT+QSmVBU2ypcd9t4PhVXoLxF3VM4CDgwRGPyB5
S39ZRsM1jMwnbkqndigio+NmH0nlZCEvffNbGfk7oi3wU0YCynirgJnKvkVkioqa
laZJniiE4rhKbKCaMit4Vg0GqnC7FoNWrk6fPo1P4FdmMxncnjnH1yJW2sNCFhz6
Rz7mA9Mv5juPBdtmLUeaYOHp40qnsiH3B+sGTNBBW7ftpUD5ZfrRYRnH3vMroiQR
yxB+Vg1r+A/GXAu3rD7+LM23g4frHNltfWyIfIh22HPPy1aeCxdNfAMaCEzCeP5h
9k9+51dCrITw0Hi6DDVrxWoMYcVeS/x6CfFHqtC+5I7T8vvYP6FEWhH5VCioMdF4
KFOcSLja3RrNAaO70KMdzCrxmkSExGSt1GEiMJ+xloXP2WVCQIE76nAT4/GhLe3E
sk5YH8iD63JvaVn4384Vo2NttUu8ttobAvHcJOMo6t58GypWADDTGbBb0gzRJRB/
D1pydELJ9ykJpiDVsEj/4+JlQzaCtiylEPZF3n+pTJDRCB+X10RWfHSPwaRzZR+V
YM5xOPaJ+Ggg5Jpg3VOqRZpozCb5I0mKX9nEwj26BleSBx+AQz3tWlHVudwpoIB8
aXTMwzgvWf7Q3BQknog4j6VM0C4J/5Ino9N4DbHaQsILerUhVgMVJZksUotMdAB8
SaZH4G3QAcHSGmJyIrlx4QI9kSdYQ9Jid9h+A3EUj/1QQcBLT3oE9jNpRiokK68s
Fd9CGT1w6CXHdplEFDaOsOOuSbXMxqbFLuwQAyQCTIH8iyOgh5tIAUnCGoh4/KRR
3YmUBRze2A0fnoFCJghfrD51QUbJYcY3vVBqSJEE+rri5zfaFw2Kqq1cMfHdtNp8
H4FQ1w9U5l3dlq48UQw63fMH9/TOc4m8Vv/MJ0ZgSa4Ax5uCSb7kX60NqG1hr65+
hZts5ncR+3XBxY7adnttc6mMDv0V8agGJCZ4Iik9niTlBntXaO5dQBSsuYEuT5nU
UG9CasqwYB9Cxq40TW+GbC9xmVqlmYbKQZfsCUbBBoEJ9CnMzwlb9hSnauGoKwLT
gTJH5pmElYYRuqDWuD2SMrRU0fGwc2z3/XzfADO5AKdR1FJNGF39Sm995qh1CQpx
0sII3zE15QVFhQ+4MCYNN/2GrGDjQY8ptH4zfTknsFRWtxMf71XEFJJkgo7WHkYP
JBy8ESl2nnmLM85828YtG5YHHVg3mZCQPMnSK+/S8suWMAlb09d4ItvoJJ4bY3zX
vHfDnQBznq4OhfDWc+PNhQUf4WC2Wk1Qp5uJFY2UqystM8NKDfCNymXX+XmFAz/+
194O9UT9YZwHwcnuWgy2j04wBRRwMQ0dwegeHIFoqDtBT5Cv7n3X2IftpFR+KBV2
xosKIV3f0AloHc3MUoulBeDGkpLd64aUA3Z5Kux+xzxQtoW7iVViGlv+BSctKg6G
qy9OCQXp66NqlN2Vb37KKbxvFzzGwGABpQQc+GwiPwrzZhLxprXzBa6r1WZ/5v5T
eJtNWrh7cyszz6am7la52dd6O5cuASew7zHuewwrj+d5fv1c9r66Luy/YLKwcPyQ
CIKVvTYrb6R/7wXJYae6S+TuPiVTCAdx3BDN1JGXOtAcmtoJT7JeJNEGwNueherg
GXarnLLPI9iVC6WNVjOEF6LxTT3XaAlkqshhSoA9nw1BC79U35vN67me6VedyRWw
/r+vpl932KsqbDp1KsVBVDV8C7QeBUalfRsgwj2OLiftFNWCj0Qvpj1XNZp/Mjvf
ik+8OGeBnEEpQGE9EMG7B4d9E1C8apWlYvAXEeiuyj1YOPoK1pn+hkyWUDuo8kPk
/+iaJ27OUl5oBScnip5lsfnzFg+dorzatVeAWHQlOgFpWNLZIeucPg4jLt69RTST
DnRtiwmePWqV8PSJ0bN7kggqAmoR8Uiu1IyJHap6KebRyqzs0sm67Law7Hhst+Jm
ZTowhJnl6oklH6aHPeL46F8c3VCnEcAaHqPkh8Bd/XDkFlw8//GOR6OcysmrR7pD
JZdYzxdWygWpIws9Fc1lRzlKgklN0P6a+OZduFA0/yIphVlZr/GHIwZZets752Z+
MrFyd9xZovLOHi2E9FLIhV4ZuBkJyAaz3S57k1qsEMcDseQBJeQDxHQq1GfnU9GB
OYuQIJHNWFgljJ1nZSRb5NETz36iZ4RbEsR/Dz/xSAQWVMMCcpMzdsHUOeKhXsTb
B+QVuoeI/RjfR2h8/A5m5/n/agUgBwB0fvaIwkd6HYytGSOiKdaDD1nk1z31Atr6
neFkyOfxv5oey+187ot9/RnvWLjz+rpaC3YPbHTR8YG/SInR0+3sdefXPYQFVxJv
GpvbSHqUuzXXlG+Q1uVudCC8Jvyyu/grOrht+XG3/21K7IvfvjRhe1uBdGc7PVeh
X5mLVHXgZHMKgaxZl98RQrXPHrlGTJYsy9BOS4sgp5LyxDWtFoWdLjMFobFJ0kEd
EfSvOl0gT3nMw2m6jKQHhAl8fy0fYUUjMssJVjR4zJAI9H75VKee38BAKycDtVt0
dd3hcnk0x0lR3pw665t3i+a9cBI+x7Xujqw3j8U/yXVZqGe8gxxByMVlrxU2eQNJ
MPzceM21gtEI7ZqFmDZlUyco6M9yChvgYExONKZEmpjR+qPByeoRSAKVeSdV0Gt+
cQLPxYN/kTQ/ldVHNGVEqBQsFWJGNngoUVldLD5wknvLUMpZf23eBsQjN573Jzip
tsU7rpub0Z2A/X+kbzuBzx66cVFNQtJ6eyno1vQ9WqO0Gwqjypo5o1r0z1ZAxVrc
yx4raIDvYWgh4ffJGsTwGVwyIyDk1+7GLMScQkzDc++9SxpEtyjf+i30K5lJj5r0
gXA14UA8sF+/BVZEVVOFBt/1OIEW2cKTtBvTAuXmU51I/GIc/gL9v2yS7aVnpjZz
Iy9owtgo7/LPCazeNULOSiIyJW1XGhf2jJqb9OE7kVG2T6i5Nn2L/GrAIhGb2qiX
QGw8GXEbWkHn3iXmNQtN5nvrVha81GelqC3DJeJSHLm2A+v0rOI39yfwF5gFssNV
+iERk7pLusBTisYE27ycrIeF8Px9mvJh+e/tw3ZsHec9H/VPiNoeCbPe1Gkiu3m3
pUfMy1+GRGEE+ooHrQ9SulV4TrrYCVWTVyCb10AtZTmWAE8D3YM/FsN6KP9mYiNq
UhBJriVyUDV1ph4Bc7cq7rSHeo+yolmGD08Ng7kBv1X2gE5dqodnpAiTr6BPvbjx
RPsiL5btb8NUsROqdJ/SgEEfikbu1P1VfCTAaQz7/XjPOv3EJ3DGMWM0RLVwe/Rd
4B0/REp7GY9fVDrB4qGuwDfh6f28sKiR7aAqatKijq1eSlObGvYuhmeXdS2M9DlW
8FrRSEVp0S3fbweu4R2zfKwlEVDZaNWWOtuTTcxX5pH7ThaIfG54ymPsyDkrZKfu
uZVIsH9oPdTgPkNbBOvNLuaw8DQVAW8qmceX+b6lswzetwfuCa2PgHcRYi9HfOcW
>>>>>>> main
`protect end_protected