`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12160 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
VKWNRQF+vfUNEEp7apOJOYZ+3DIAZ8xzuX6OZ0zKxuRMf3CFmE0qMva557bscLmf
6jlfngou7a5toasLObDvc+z01QhyxyqKkCE8F0Qc32gLq2+yyJBWHy2i28WKbU/e
3xXzHzYfoMDoUBAHsGORbfD0nSRkQIZOysMT0wyBUhJLmXidZRreKVdl0hrrX5W2
ohAvB2U/3+csEcEjL1QcBsdzn4WjzwpRHLTMl9GaDu/1WKSOAdU4pHsxsLlyD27g
tqPLKgoDiktBKlS7S0LdYPEWxjFpVQvAC2gzV0QIyuMtUXsXiOOMOoMy82A192F9
4/24Bn3NUAoRd+Q7vopuMpLHrRFXT0wsJYuSscA+7oGMFxeoNP/Yls5IfQlq9t7Z
3YBWXKVaMX21tqki/hlKn5uGrz6I1dK2DMoOlh8QPLXWunhqfmzu3WVyXECRvg0F
wQdpokKsPTwapsvLQyVjgVuy1HlAR2D75XzyX/cxJUDp0OSlRNDS/Kq8C3m1o/p9
Ub2usL+gdEH5quStgg6JPncf9EzHBulSPp80d1kAYYZXx0gc3nIszuJBRJaIxadT
OovIIg709rezHysXYRlGYPJuQVSzAB9SMbchU9S+kCJziUpTIBwRLAe72thuWG2+
QP/njlF7RSzfcq6h691B27bodqFT+BskXJmiPf83g0p9pZAFpt1uRUQEL7b3QuP7
ecBWSVvMbfCLbZTkpgOCOoxE6gs3FFp2BULxOt93obkCRuHOrAkjEHoIPqxIIQzy
t+fAUXLSKGdkhc4I6NHEtHE2FGeVSgXIkHY4hKl3Qofbizmd64rc1SyJy/thViFY
8mYkQ2BU5IYM2eTrxPeo9UVuJSxdZnZcleqj9mbH43g54E5TPkaAyxMPd7H/0KUk
/sVm3rLCuB6cSChNSS0rps9oSVRIf6U9Mpa3dHC9GkPQz1VF2VLU6ZdkDa3X2A/w
0Qm7HLS1UfKKzfykvYEx8tdbrA0yDS5R9pAkakh8/68tNKmnShueyppLECpShf0v
+s6sLIQZh3louB3NdKNcj7b8WnzSIaJ3vVamGEEO3KXY/zfXU3qhtLYdE6bHNaf0
mNUAm+ciFEwx73seOA4pc6Boxu0a/RXguGgG7zpvXrBIaVuyyrm9XR6TUU68VgE3
h5C+9gfIqFCz+TgZlEq58JkD3wbfUqLLBXFirwdwklS8TCDQqnd2jQqUuuBjQAAh
MlSsU/gXibk7oZ+fpkbT1EgKsYOht025uiCZOf5eJvYghhFX19PnkWY5oHaRsnQw
dX5T6L5l+I6XbIRIylcFBFcTgW5NnrYC/Faq5ao3JqTtzmmM1pxuTKYKR6ax3dBB
WaLu6kCSEspxFGQ09xdOrfHkSw5kfKVzdx18CoGVjQ8c5mup2UvrgqdoO3bbSJ5s
fHqZp5pVykgjAfCTuxiESnbfnuFCaFh2w6uzZ7C4+F9711X/eMOT9HELzPGngIgQ
lr4RC18uu/KHqX765IofrmCQd5OGnOuS7TEcpu9j+GdMxWEIcxSdvUEIlSz9TmmI
Fm9xs7bTkocVpQHcVIAKKEXqh9CIXITmPtyEwCta77QieIa+JdpMVZjcpe70iJQa
+1+HwqwGe0Q2a1o4iI6nlVK42CgZhsl1qGxxw7peCJoFNL7vM7sgsbJqRXvz2msi
wrtF5xOhFFQ2wIo3FXtvpoMI7wmdoopMTHOd3qC+0pIfzHBbKzmakRgPR25Z2WCa
pfxWhKpTm+TV51xy/vgwu6s7F2h2feJTW6rfrc9PpCqodMnonMp432sDtYRviMzT
BNrZ3pZu7y2zoPqVa9/ibdISZqjlVhTzPFupGy95zGhUpVTiuilh/0DYId+q0htq
LjD3ErVr9x7UUY+ucuKHq463AKv54OkYlyns8bzReEt57k3t6dTI6MW6K1XvFWQ8
4zLoUBocfo/Um/Mds5AO+H5wr6WBgGpH4xDOm5uCT08JjrSaco8NHz2TdjYX3wkw
zh6S0UrCWa/UKCAYx4RUE+nUKNp6gnLTtbiaYl5YGfL8DMdVp3MlVOnY4HZ5GeJL
+rNzsQRNWBjODHP/CxxUj3t6jGqlma+fVavse3XKg6cGa7JNPA+m0SHjiYJ7L1ri
W6G5I5SGZyAWHpbu7TClrXXcoeS9ieDbZPCmGxY2oVe9bqeDRu1dTTqBc9Jk3swM
+6BGn38v1KIzjYScOde52sIPbpE3ihq8w5FnO3vSeJ14SDrFmzqUDIHKmX88JhBQ
/Nim8NxGIgZKMdt6XRZqpwLaWHQ38g3rlZHXv6IlMjly+yWNMWX7o8O21G8w2jNU
TbEQMPucbPtKXjR/7w/5GLSfPxJWqBQBunRiGcImlix8bayW9c9rDMQk7PeZ5143
2wQiraAbwgjxDtzWub01vgIU6jW4vGTrzAAb0hlMCp8U8JgCNe4DiBnY7WVQ7J0G
xedpitjeHxSSlWEz08SGgZwi4VKjJ5b0FATBysmXOPwSz1lUE9xPOmExgoReLWCH
0l45HBvtVpifBHFlLHWbqwkuq74q+tWRfgva7o1rMVU1j9OhgU7jP/lZScCFtXT5
uQ4e7RVwuWQBNHEY/SOiFal+mawmjqWB73P+s23Or/PkyzSLkMLqW3UkVRffW7pv
hGzyT3g7YYucE63f/Uc0PGVvzw0die+T0s00PfBoev9Zun54vT6arMULvIaZRN3e
0w4+yqZtuSEBa4eeMFSr6rZf3zcCFk0anuV5og4FI2e39rSkhpluD73Tlg+h2w6k
Xiv26z3KR41s22WF6dHYXYPjZw1mqmxGIpaX3FgTOLOGHrcU8YHTg1Q+RiR452t8
bxL1otqscWiHFl5hKVVR3krf7nkZ3JdDpk1PLxnQbZGqmmRSvZq+k9/FAB/E5Vyl
O1vf4yMA/TZqqfD6qpjgJl+vixX81SskcxwfGbVKksOrS0B3LJRM2EH/oWDDezFU
spfCEt/ReUNr/QI2bPfOZtasPzXDiHTxLd1QMBxsqgzd9D0BbdknptD12ytZZKNw
3Iii4M7qNTd0OvqpjtklmsOH+fJ1+8hOboZIlQxEH1uHj4iixf0CQUFrRJkNxjot
GMnUJErPHrO6sT3PdyPxF3DAFcbwa7VGJfzwZwmAANELfDEpGFQYVkTjomvF8Xvd
CPLOaAo5oVrGPmnXAuRS2xqOim2JDb3Tqsql2T6nzADkZIlloTGZ92y1aJGUfrfM
aXdVLYHqIo4uOMTL1T/qL55DR2Vw7GTxZT/Sc6sMjAo7CK2AuFSJ1YCQk09QgFKz
M7rOSjM0N0AzAZohTAoC++hjmhoejzkAkVkWT2EledCRUE+f9XBROhYjmGSsvgpP
bP2ssEMxrQdaD0mORRL4MMIlg/m0cRZmh9rQWAbNxOSp/8gY8Gs1feD152s/U+14
tjz6XQ6y9EKx2UeQIz5JsMiJSl5ldPAfFuugG1cpsmT7huvuDmYL1zc3Rv1sIGVA
qYHNZPIqS+EfpCUcTWjr3yxqiNb8nQnmNjUDqAKQv+yyFAtd5ykeJlzvjiKo3UxK
c08Jzsxb0VzuJKRnOvDO6+2dqCUEW2B0XHsR4Nk88+rINsr2IpuseLzxzPh0l5fU
RGxbG9hw1qzU5o/05b9JaG4wr2Wpuv2X/oBwPrv+j0jShfBl+dEFXwrw4hhBlUde
8p98iX4iOwq0mKpm/GT28Hb/MBPwaf3HwFHB9pPr9vgVKs9VquR6Sl9c9qWD7A4m
QpvBLFPSgkRq2YyeBOhj6yHPp5XHq4/fbopurRs/U4W/v2U8qq8jvFvI8KoPy7ZC
jJcCZFAfJT7J1YmBQ0+QXktZ1KUNaHi470ELC3ukcPgl3tfO9qBXv7UfqSuMZfMH
H3TbYsC9kRpoNxR6Jrlh391epUf/t9vX1+kEViCnASQQ9eGoa8JHpkLcTt0Pk+ub
qyvpuvsQHhnumKiMcc0mGN+zoFXR+e7kuvk+K6Qw4HKISKYaV+9MybuQn5ZV6QNs
9XEtQYMOvvzum7rcwdtkiMeA9CnaHDbPSZTIXGEP7BMkBIrqFAE/+psflnRZM2T4
oRF/bDKWJZrG5LAlkVDc0EKTEznskUY1pAZMwDAW/AHmoPjyrg5KzB2XnbG05yV1
QhIXN8kuzW8SfYhQWg5/D6lJXU8JtIa19bKFjx2gCoD09WTE0Lde3NayrzNtRkHZ
jQHOOls/rvTJ9zV5alam9ya53w/799c0LCtOYyk2pazexZu7jbxzdUzTgw9jPjiO
HAfkIAUlIhU7fN5R1BM/zsZ3DZXQ2gfwvDXqrVf4pe17IT0mC5DFLLB9hr2EcF5Y
CtrHp32zpSWpfLfC5RltO0nF1wlTUwBIipsG45EIZA2INFYNVTpzKfPka3qnPjGd
DThSb3gNaxyGsjeY3qq+khtl7HMb8uipQaqwGCCJ5O9Ps3MGBgBBO53ewwRIcnMa
y8BZifseeIL+ruUWbpgyZco1bip45p7cua9SFVnaXgbcjPCumyx1VSPMAWBTAj2Z
kHyn8Edt0zbJh8ccVpW6hyIFog4oZvYg62QnKWhpoul00Z7m7HdDIcm3WVfqAfrx
l81wrP3Vd/9yi/c1kxuyx5fPlGvE/1kC6f2CABOdTfF26nc1Qk6YDJ489IAMZCqC
4BrE5Bw/ANS31FtTKMYVSOSFgrjKXF07NqKgcTvyalbM0FcTVNKyqK2e8ACzUXpd
09RN3zhhv2DjX3v2Nbois3+40LlGBGan2LZhFPG1jiy7Bka1RWgyMKKVbwfS0646
xZ9ZGVCTjHf2m+Hh09NSJjRELQ846RtybIlKpQq+wfG9peaHSIa8a4km7A8kOtuP
x166B1BNsDd2GIFc3iVIlPP0ZIAhCT1caFGm6IaRJTTmOVZjvDpr8V6oHArkzi0A
hgK8SnPjoggS4O64SWPcOizHXUXd7vgk8AY+PkfDiDAuOuvuACRJwVcl4IG9YBGi
vsPA3JBbAe5Ay/nmKWVyRGKZQXqYi1q9EwNNYupWDGUoXcAor1faMChY2zmzRM8q
NJ+rQkfIMOMV5p8LLBg3LBszntz6nYGsO/ADZejTlHZTiHXfLKyVvqXeALeisfJh
2v5oLkzV67j/iIj6QcezL+83dh8+DmqVOwTpFWJjlS5eWRO9xeWt6YxMtzuPE8MJ
aVZA7PDQ3EEzqJo1Fmo54QjwqSVpMFs/fWh5lXePjgWEyb7BJEC6Bl/1A1v6HqKB
drqMIENeyRpZ5EhdkU01P8I/x+HSICmit/W9sB2BzpALp469o874ad08gG0OXz1v
/CmRuiFXqW6+syEDdImKly/B8BoFkVtl0Ml6JP2aMuvuGfrf72Nfk4FJqkaotR4I
HvdjkATUpG09R9yJ2/DRVChUmDkwfFL97VqX2Y511icQAqhhajVKvtV5J+2lRk3U
+2JkesmsrsClmSqavLSEGo6oCOrw33b3A0Sd+6o1I2k37MryEkvk+ZCdZ/H5XtK6
vI8LeWD7DZeXog46dssZH4ypDeIbrvALsK2oqk3tIlnv/Jw/KAth5OlzzXsyyXgt
yIFNPcjV9BumbdEZNwfBKPqjPCRPg33V0W0IU1MGIaKyAnR7stbERkNkatJlMI6z
Piu2M7/WQ+XtmuER5QkV9/hQneGQOAOZ8B2GNoI4YIO6yXZjpac65QnSjlTKppGe
sbbyHqKE8Y24W51RqgRjwd0rMi8poLGryrnLq03hf9htd+FHFkCSyBN9tcq87ljJ
2UYWWOyFfqRdeGXKUaVVh87ALFmIgWnT33a8Ly4IkYKzWr1ZfrTW/V+pPHKSKhcB
jdSYY4JIGFmEVoiDp4pXxjHFcGuLzRSO3gGJ/1qMowAyirO6GkjspXhYB2GvJhV2
cHqVQQNqvDzvcq+lV9jDd9VgyV4NftGLbPdlJSNZNmc3lMnv+f9DJXeFpwxKUQR/
oT2+9eEMaYDd0zz1jLmr4GcTiCTjHR9JIHE00RcsUfmT+reW6QBeltxTjoDf9hFS
ylj06o+9LlcbhzORQmwX5YMY3U8LDCdF1DN5GLAByFBxG3dk+Ck3evawqmeGACbi
llgobKL9dNA3QcEG+ll/VMsdIYDrLlMH/Rchi3k5v2lh9hqfhEfcRy1BlY7FPha5
YMIzQXzoGAdfCTbeBlpe7I27CdEMjoI3QfR+nmYpLcOkDF7ntOk6Pa33opfO/qRu
DYlzbf5kWJqV0/4L3TRe4MQftwF5wbHvFPtMbCUwqgRUxlf9lKRcZnZOV/XtjjaV
kpcpBeQIlW3YcLUOVb9XTFp9/6fpokNRzluIm/W8yydyKGZyNc04imbZPFheQ8lp
scVeeZ5LNuFiA5PVTgA9Zm/zKOdGUw+r0sU9gsQObsYJlijBgT/KOVHUwsVx/apc
c6UNBbn/a/j/5CLMOGxL8qQDk+NxnghgfXqHUe9YRc37ZCABcM1RYz1PbBV/C8rY
bJ8q7mFQNH7z+L33A44LvvgTnZKfDK5rjZpQPnOoY3jzP01QIfdldZ5GouAEDvIy
nie9RQgkmiokOlN9L/ipELu/ya/zVm3RkpcFado9SCWzG1/Rc9HlesXydYJe0EOY
9avMKOKzpDArvbWxPMRoNkoSNlc597j5Qve6MnUgyuDUHhhjZQ+VQrUdMAP8FRsz
/LennJwXP1uEUaT4HX2q4jb9FWMiAdctQFj14m9v7PAdqwEoqAmY6poDqR5kztf8
QbFxbSK4axXSWK4HQDNLu+YT/rfNc688cDX6x9y7Ss6mN4UTlRZxcDkt2vi0IdyG
nb4IHsnQr7uVp686r1GL01intPRdfqY5gR55t8Vw3kg9LOgc9bjicVU4v1+3pzUH
Vhy+VFroyLEcxkIkt/VtW41aSrG+MPhEoCBu6UfjJbITr91u/9P5Gb27Kit4KPUR
ScQhg+8VeVXb92w1jwDsbbigm0lFyK0jsoA/NH+R53NzsBooFtOQQkTv9DU/yEBj
N4oFoj5o0AY7IKt3dBb/HVM4hhwL1N67RS3wDZIjPCpvBm4+dagwKH2pLSfQDu7n
d7u8JRdyW5Ri1cg112aAE9gPUnR0AjvZro0r4NOX1tBVNeye03EFKYaTRuu/0I2d
Bs5as75i17G6NkjUPaz0h+Y0tUjT98wMebcHntSwiWso8cn6x+iJKbAXUpTO/Xkq
kke8p9izzcmxJzNMc2vJE8Ku9GK5lUXT7eBI8Frb790CCB3SusgGq+Pwj4I4cfW1
e+PfDcHAYTLEQiiBYL1NTk2yEcchpFmfIb9V/MrD+EJUYcdoeNYBoQtt/TwMEeMD
+5C1WETZm4kX4+/pBMY57lbj21ipO/1IN6/QiJyXW/yb3hhDgpwxsTP8NnA2ljNq
v8RennTrkQlAGxof2snLQNjUF5SMICZxlYQXjSoGeHiwxlq1++JNStbrojSmHj9q
A5ieMxk67dQ5YbulSI2eykmgfWINmhvgjNfv1EfBsuhmKLiRclLUiBgx3y1XufwU
e1aB1wzPHhnCUrXlQXFB3N/Xs0VyMHhxzJhYTrAW7Uf0yX4vCVWFcf0gx12O4QhU
Wv1U1jkKU4dYhQPI3Yj2aLUrGusv9/6nEO4ZFnOwRXtnMDEVCs80MW/35Ep/N1UH
+CW0xELaSP2/hyz/bXXLCxtyP/F0axTG7W2OzAZO2MXCwKpcwom5NamfgqGxDV9D
L+85qXR41VUysR3IoIOa0B2zZSgF5gieX0YyTygYMPuiyNH45ajacYA0EQHKNpBM
SY6CGhvJgoVDBEKKaV5syW9QLBMDrQwcLAeWbAOdPlqr7rm+WoMxZqXdYWL1cSMb
WcF8xROAJxg5PucWkvf9MxOIBp5iRh5/kddMPPapKhPvElQfQLNf82x6j72ez4ab
OGmxXCHvifKle4Raz0Inn/rXvS9hZZHbc+HnthpDiHDmenmIN88tWVO3sTPeij+u
2yoH/GvIPzt4adOyw3kKC0e8mR6R4IOOZY/yZqlys+OomLqOof3siIXePZNfVp62
zyZm7UOoTe/quj9E+aBvsyRt3Q0gEDLop0Ah8E+DLIz/cbbDFF8bD3hLC94Erc2n
T+/FKnw+Kh7mPoA4sP1jSxOzUV2K6Bn/HOT42/aubDhlq0gX5LS2nEUkN4Yt1eCo
tdp6AVSdu9Mdlpes/xpUQh1G3HEEXlwBhokR2A0JkVze4qGhVz0Ok2HUbGnE8Zj+
3ne1ISrZ0o/mVshcnqG9GlGxIZaRdKM/zcoBLzXI3+bv56nHrJIr9g/5avUqCptY
A4tTrZKtezkHqAmjMOpC5F5iLfoNiBkTuBUM+gXv/v3JDXMaP0qYusJaXP2DEgVh
4TLznmWc2bny+NoYVAA0yMTF52mgYhHgSi2MIkSFOdEA2CDWwRS/II+x4SjHKM3w
O9Czq4HA3kH0Y4PXKjC90NcUYdsnWQI0ScbB191QG810j3+tk4pwEh756PMpWg95
eMECwRxuJc3xYAdMFz66/0meB5AQzguyivDtLcyMlQFG8ypaGQHf2+axOZcmiBg4
V/1npNmSPeF+QBr40DLmgRbGU3ZwmBu0Q4PKF0FZjRJwPdbSi7Q+hs4FEoqZcoam
xmc8gz6gUUofs3u/opZLzqk0P5+zIV8vFFL4y4eWs9KVYIrgIJkjYvmC8qenNGwo
6SozU1Djvl1LObnEWS89f7eP0Wag/J/N3qerk/o1CzDc+VBusykA+fH7NExaLM90
Sid18iW9tmngXNlSnHNZfjfrjS2x71XJ8EQLwm1HOHXfT1W+0IAX6iHzk60LkWtJ
3R4l+/GZAy99n/ODZQ8ok/81IfHDfOGdynpOn/rfpH4tptCUFAsxsnMEkpINq8V9
bGjko7QMSHXZXQFwEkTSpU4idKsWgNtXvkaJYjTpRknvhsZvsFpJn9dWxnMRNEqP
99GbyRN0Ta5e1+ComK5uVN8pRc3PtHSo8Va6Ws2Ubmj425chqTEoWI02vBxLY4Wu
N0WymqD73iZHMoU3SUq+r+vURGh+ynKRmqxC87B1RYcFUQaWYOwaYpK6zIYcqSXQ
SwWUajoLtxMBuYjZD0WI5Yast1ft0E/K8DErI/qeVc8OqSWj3y17lu3+/pG+66PY
4QAgWZrEzaVbfMpB5cdi2LzHsyjWML9YcNhTMOuXy8WaXrv8X1jyacokhp8Iwmx6
+/PUWAyrElKOxmdpyhhc89M00/sleK5yxZwd6UjU2HpH8Ku6b9X7a6+KyU828WP7
1+1zUkViCMD4WYPJPxdHDhiGidFJWtmFJw17Kd++IjyEmgwPQtlypNviMhgc17BM
F6khXb8bxxZh4jdc6tYoIfnFN6e79ZsIpIOcYmiAXc/FR0akWYG4oWzqub/OWBWD
dvwPI+pmQZZd/nZyiK/zcR5WPPbYIRXD0p2oIXREBw4Av1zh4H9GRcLoDpPPWCw8
95/Uw2CeHEUCQ7gugsvd+DlwBZT/JD/g1dyjuYFMIZ8x2Wb+bUdndHSDSUgILOrR
Rdy/vnernL6yiOgMFM8K47h8QDfEquk4b8wQ+AU4ZIcpCxHJcyRpiH8K/vD0iB4Z
V/PHNrbhpSwr6n+X6wNIwsp70r0Dx4wl+FJAZ6siPvpI8OUzXGhjx+UJQsEwThDY
5Q/BUzI9+vhtaOD9GidFVKBq709ldpDbeKoKXG4CpDWUglJvBRlWhbfJv0GM/blq
C75v/WhnC1ac2f+pRuZK9H6MIGQcq7jTf0goBFK6Uj66kVT2/VCpM5X4Jk77e4zb
YkvqwEYOr+IovuOm0aP3jF8HK59MnpkmO+I+hUy6VudpyTklRjzOF1c9ffHcZ7Gr
QUN/DrdWPyJEE0q8AwlbSjCRgxMQJJAqo6p6tpp6RK0duAS07gdXBWlzKBbLeG9M
2zrSxRIuiUS/FrRIMQXJmmTdwppJ7Xp8zU7vC3bYTnR9ecodge73eZhS5S2zmSts
xOZW9NCkk7GU0LTCCrMKiwM1gE6rL3dNCY1Awty3zKNgkenoYbHLOHDuCBBXzFsX
BLhI6UVG4rELKScz18w6hM5ohDUU2OYXJEUYqMmDsKNBg82rleVedgWFGy8RyJN1
2dlkl49UolK0pJqqSWGEhcY+1276fZrMPAzL+aAyFOi5pcR42kgkvXJWZ/VkljiB
ljx44Z5hsgsYMbKOTezBW2v15fL3F4MT/pP/hqclzDGCmYJ7SAnK9/LVJunTwKyf
p/1tzyow41BPGv/MI6tyHVOsmRH8ZuFWwC/XQ40VTA+mE5egpLlI749/WkSOqfxz
jueQlZFZV42bJtSUomi3pWLpoEnFYINZFv/P0alBGzkMobEl7/t4FjEKNi4LI5fC
sxnEOsWi7xeZyZD42tliEClSL+Yg537rn/ckxSUV7eeT8iKVbqBzyvAqLvB/jpmb
awlvOZePCam+7x6U5+TJzrJ4u+kC1MIOtpTsGqGA0x7oZMoQR1O/fql6ndxaNdbb
3cIFd8+5axC7aOWuCpAJDn5FjRFg1UA06LVcz+KyjbLVZRHoeQSaeTRJptDjurX3
qFpubcI+e2JjkKvNgLlpW8dstRxXj5pcJogFLkdLdHB0Ty1whuLyXioPSNqbtpHp
ewVaPVx1vMOXnBh3ECXaPBVxmVOX4vTy2ZeT5e7kGaB5TUXI59yOOcN6kbWiARtf
dpLp5JSu3SIHRoDVgPY9Df0/PVN/2MOfz9qr1w6BpAgRrIyACIJFuYUT6oaSwtSk
8c/IML3vdt6AZLjyxuYs4Dd1n+Moadcfr0DdPzm4tahkCMKyusl3K6pPxvfLhaHH
T6CIC8mslT7UyYqyzwGQwCaM7q0rfTQUgYL3CAkF+8Prxp9mZ2i8todnwjxGlNS2
iBlIOx+LJBqF0ZJGbrnwSjI79PSXWim/bAsvHftzEZmuy7pJrOUCo5U1YQ1SlAAA
qpjegjrwrAR6xFBw9EiNupI7NjeY1jwNQ2DmyacmkO97D514JO9RPjZSguqb05FU
XBV54NN31Z+xQ9jhW6cq6p2PwLP/P2ssxsZ0txuSeP6hQ8wRXlmLLFPiHdeJ/uRv
kk2c6jyMKycF8XIhRBNSRV/ioH7doZUej1RIN3VodKdsLRlSnOLYsoYkLQzgLp8k
xZxzqlL3HCM8lQieej9nCC9j8vnrKRWdSOJq0hRGuUl7bBXAy8nWSjGxCRpsmv+g
YfLCmBzZDa2PjzOupMrWfgUKA7N8ru8RjVKPp91Oz7fF3LTt2RtSzVhT1I3xHNz4
tYjbfcez8Oez5G/9APYlCpVI47bodYtPauX4ZGTnhj8zgd5ysrdvKK8jEUfvsWpx
ZuudlpTpmPMJskGRVKd6e2s31m/adaFsAJrlVgSZDtlPLOhWTg0xiytCocsRQ/fT
uoupHVSXCXBMYikza3sF0cvQ0EfqJVNhWlUt6lI34FA91wIQpAN3fqeDHmF1ZKA5
Y9bp93ETE1dk6xV4g2Z6vwHqPerJBd8N7HSIHrXJf4sTX6A82WFc9i44nCEujhk8
Ys3cDLpSYbcnese1XdYeQWl58s0RZqN0+YmRdJ9ICxAgUVg08aVRhL7ZLmsJ9FCX
RqhDTymh8YpT54yw0MbDuilNhUreCUmN66BqX6dFAhgCgtOkeJjR0mjFNEs8E4VQ
T6hdPIDJ+e1vKDhuyDo1uv3begGjDe+h0Ga6JwDKEJsnIMSZm6YXUug6mtqkhyAn
hcbSDeNkbLib2iLdUTTe6h8ZdZQDc0qtkomnv0ksbkfWXksEdt3wmZAEyo75M09S
eBktunffOWqJRItc2upOUAtrJ4NzJdMoVHu31xj6NEKaiWhJy/XR08QXxfmlw8kR
qRTyur6+jvE9vfOoXqPLd5XvnrHXp/hLCIIHfXwpAm5j8dOP9Ffbfjr4zt1Rw4s+
ETm03tFpLrsmMsk9iVKBeXClXQPo16SfG2H2nw64r057I0QVEH4pAAfxzIL6IJQt
lID7SKW7/D3ItOba+VW6/kz5bdR58RXT18RDq1nm3439oJRxHTSWB/Z0w/Pvwafo
hvKN+WGxX8Pxrii+aSMx0m63H/9jiyMcqkdcm+QqX/6mUNnqIPayghQnvZi/mXoE
bhCjGss2dE175u0iO04FIaoh0uzUnDZuM4YlXhf5BQem+YTnSekUUe7kdG7oDZrB
wClnfws3efp6QJMNmeeUtKl1tW2V8i6SrkHzdzOh132wMamB7ktg8bakZivjxpqO
nZHK9Y+o/hv5SR8lGsapdHFQQ5EjpoFL+1n41K7xBsvGP+1yxlYjIa8c3dSkIMVs
+7+57BvN7aZhEZQ45hdw2UcpuJ6dvzbAZHJpdaj/oIseQsb5ovWMIfZcP1UwspCJ
4lrP22M3vuCc6V7Ojrd7R3diOj/fKn8XfT8yYRibUG5u0nd9xvSKDvL1Pif+OZSz
j93pnv0LT71qdRp86gtT944GMpeMiq6/OXLF2Y3zHukjFb6VTG45j+UvjxKXNUDR
bV89lmwucD+0k3ISD8+0NHj0eo31dhATJ0IKCeH9xHjKwsELdYLtHtcQhAiFCGmS
zk/jGQ9w77LtmKuxXzg06suDIeTO4PWjPDU6pXuZVN+mwWvl80UANz0tNUqXSskG
fN/FoOGe29D6TebcLaxAYCLjxBtqWSjZtQmid0MCoetiQb7hfRFXRDwXu9TMB3yx
jgu0R23T1wb/LKd5YCrJsrJU3hT4s1JQ9WwrgWrudg+hcqxenxk3dbu9v2UdfPrs
zPoGHdW+mH0nr+YsdYnda/shaiGPHoYC/jZPOj/9JPuWMc7Z8SUG0k4UY1p+g/uA
FKLs9OtTRcWxfEGHcTB+y3cCr4EiZFaNQ8hCLYZDkcEdiSEP3ODozl5NpstZcQZT
MCiegahnEPDtLBYKUc/ytfbHO14UvE6pfVTdGfjhyROSlPkLP+FkcQnuInAw+UZs
jAQHFOBKN6NaEdnUnw+ocBeYSne6NVNIC6eSN1NupEy44+3xhrZFqckLTIo10A37
GEFGXc4KTcBN5Vb0CLMNo4xp7/GS9suhbo7EpaUQHBwRmtz72EPWPaWQz421LKP8
o4J4hqyZZVnzcZ7Qs1tCOMdHYdlzv4jCvItHoeJAIKSc95ZKqYyKTHdnBh7eo0P1
ExHUjZiNIybTakobBxxhPg3ttJm8xpkWzXFUyCAeNF5n5yCZw/vEpgJ+bZNKMuOs
dXrBCDQqxN/f7LZ7u7U1R29nYz2/5jdUhiQsyF4ynqY20usVr4K15TOC6DYXcp+o
mBC3vQy83KPNs7ipENYvTJ5Oe1r1AlHh1ieU/+JTlSw59e2THbmJgXktSGR7ERsE
NnMaisp3B3HGdXZxKVxxe8tiPrct4Ff9gNkenrZYSLGvVfsJuTy7xx5zkGKdsPyH
KWOjUnCQFilQOChKY9upXIwd75Z/HQ+PukWhb0zZc4mmIydWmow8aaSfw6gQXu7j
y2Ok+kSN8EMekHQf6vQEYJ502ikdYx9S5/Xt2joRYRRNWs8E2CfLKomNe88GqhvI
CZGuSd1axSRBUjdch3cEViQKfR58qRGoYzVrL7OEhwl3QTAObCmH+sa+P5zkb3xC
mOxsTESkjNlVTd/x55JNft2+lLtjmwMn6V5ASMDWiihW1fabvKvikbp39AQmsV7N
y8Z+cKu2x5yhR9vZO6S5jcDWOCtDNc813weOp5nduYP/XS63PrHY0RClbOz6Ylqt
mQkHyNVWdXQnoBZe9S9Ymi1d2HOkTeRwiZNYBIIFlVUPkLBnoGKFoM1ARLgdQ5c9
eGRymUpnFvoAi9Sy+MhHVz7beMVcQ6xlgkb5dm+/RcZhzUx/7vZa255QDNtHNKvZ
P8kvWyZZcoXQBFvVQW1Dof6t2vJQ75L7As0PzpbuElBaC40Dn3SBdjl81JpIAgij
JOiDrMtRc9rqPBxClY2VKJ0g4DTQMgiRsV5F5ogSzafmFylz6WM+iEl/eHYsTS3x
RSTOZAjNzVAql3agDEEfJe0+tDxIvriiPukCaNEujK6jKlbvrPCcEI6aXnJTFBlc
dvl9XUhQTjX0Rn0Om/0iSiUFegUDTD30bOTP7YQLdxQQzpxY2BBnVpDLq8e4Ddxa
c+R8cfgFdkwCI8OqRwT0Cxm2D+EKxTxI1Nls7H6G2x8ogNFln9sxfRaB9LaeFRvw
QCknSYmDd3Bcfxf1hMo61vQtDgTL8zX0o9kpELJEmE9/zH+P8CXaBzUexAlC89Qf
2vajcw6fi/u/22nnHAFeiIKMgxsv0goT/4sL+Z42QcBA2wSKzhjNHgy1Hz5uZaKV
SIlGXlQTzeUBkmnuS7ejRnJ8nJAOSkFcSngtZv5VIJoOrn6gLInErqfEWUnbqOqL
kM7w1ivfnu7i/AAcvpN4xkDRyn/wN83KxPCmux65rC5daR0uIeab835GKqfZhUuL
ssT2KmYfEt1KNnJxvXWHn2baHT2ADEVkDufaYFMe8FjpmdXa+bVyCi5M+1D7GWBQ
yoCSuVZmqOiISwxmM0KfcnPR3V7TABssPPzjPRqs4i4qarzIuKp12T47wAbUFA+e
6A4fHe1OAQNCoDbsnSzJF10EFAIxrPem9zKN4UviSTC/SWipJSahwP1PWtUX8ski
Js6F6Ql8Upqp2T9xbvI+ej4zSFwQ2xjZ+26sJ7neHZBVVTbU05xFeO+7ynPZoOgs
5+Vqg3m1OtqaOZAXz89YSgIYBBmWikx1dhvg85NRtURH6MLNMAWE+prtI1cunc7R
+zqFqiZNWBBnll9eTeevGuyAk4hZacuYocqCI5zQH+DmFwT5O2DXaC6TLb68jdgC
+Ess2lcAldXQqhmHMmEy/jHebB6UzhmBpHGSx3e9P0uJWMDpgHxG6+WJNJnbSnFm
2fjFGTvdyKRRXjU1qODBijg1R09rnXeukaf627h6IWcCIfRqo0nVLVdqQUXwooGx
NCFe69wLuvCemxZHmJq8prf1FLMxG+TTGDkalWWOjfjOaqB8mkRdc48sJwHi78ZQ
TAOff58sc/gSNxd/rOO9JfL4AmuJZU3mrMcb002Jm8mYMH6/Ry3CSVka7e7vwr4N
GkUt6usqbihz+4PigQfo7Xnh8dk+UoTcbAd7TsW3/1pw+q16DgRxK8R2L7WPlY7A
smzlfgQn1d/VJmm7GJgWHOvT555jVuO5FdATN7ixX0jD3OqzIFDdO74jCqyEy4cq
344CgCcFt2L3fYoebB4ODVGjAvVd7eXZaShr944VmtFvOBXGIUWJwUKXeoKYQIwE
HIYpGN/dhvR2O2hBKK4kLE5P68t5kR76bFKt5dFW5vLbXG7HaBU584FrTm+8W1ej
6G4MkIqc5okAsxB0Qav/YASyOc2LVLID5Eg8bHMcRv18FBGU5Ltejr8y0Nc1cjD/
gJ+0sVNoa41B4wONIkdIfphP84Tum3h3QKCkRnbih8OkfVlgZLh9oQy3Vp73wIZ4
Dizdw+kfPNClRK0gB3ZEO7UbliKLsintzcpLVdGHEDAM/45Zx7kvir9LXdFR72hs
3e0huyfnsfB5hdKS7adrT3XMb7rc9G/pgNh8V/mW1cILOgQe059w2JFdwwV2s6J4
86syQgp9x0O0/uqxW189gXrEFYLe7nd5/kB9hgaAazqTAKRvk4fhGrTYRrkTC6DP
WzcaTUnfo+GiMYpPCeHn2sWaRBg2+bQ1siSCS05ceri+XJfjiCswGV2pm3tv2yFq
y9NzsTYzcmhRrTCRi9cm+esDjmVfbCRhLUiStUq91v5+yQOcpaV/02SlmHmia2k0
if+YtKPpdL1TagxwY0qfKEIlTxuN1unQnXXhH4r7nKv7LKphz2vGqEkAtgyRGzIm
gsLveVmZ6qWkOJ++akMBWUp0Ll93PPCMU9HOFcF+/2QpcEHQDs48z6k3Gl8P/ype
G3N0pDAUV7Z0PhGs44DJeU0T77UNHaffF9FQvFg9FE5wZ7Ato1grHo31jlZKsH6a
C2iW5FcIbhmH+bKXx8MDnIQGhLnj9TiBL9MTN23l8ydf9CsPPoEYP1OC77xmRcTO
kyG0oBihi/+f2YSQQ9V/13LsFue+R3sw+++SteWJFf6FkUdnzta2WxHsbxX4s6Tc
JK271ctFsa67T5vJiwEIcvm9JDiUV77jJZyZMO72fqrIdrGcb0C43PEz2Idfv35G
5AfFTTjUtStpD6OV+g04mIEvxQa7yHIV+2CihtqG6rUwEyDXNekHeRONTOODYDEJ
+FS6p68++Fq8HYQ0nFeZ/g==
`protect end_protected