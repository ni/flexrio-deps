`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12064 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
L2bRNdr1lLBT0eERw3vGlCn38bEoEj3VjGQfkRM+fLz+lCMaN3JBY7KLmlPKxoxK
e6tEFLEMZnT3BWK1GWQnJkhe5mkNCbqtLmDk8PPli7A9UFZjdWvnXqSvFHa2sRst
ayzvc2pIaFAgoGanUl0wXjzNIazSq6kvlmAMPT+H9bANXNpNjaWNnq4zOeNWWpT6
CgfKB7/17zXYh9/q9o7MfF+dsqwpeBqpDjwmRMf93gG/kQqTx/Oe/FX628abZazr
OfSicHW/VSfMZbqeOqpzt7heW+/kwQoCz9EJgVzvpoCAwpcyXShzl/ntQ1Bbyc/A
uJ3C5NwCSMMrgOTnBZgG5elQygtALLZWqEykVRvzxMP0uDne2yXJoCLdytjA6pp9
ETEw7zUELLBNrvIbJKsswZWGTeuw2Ul7Ic+bCSJX2lbqmNQWQJtw+SIqgOrfSXDw
WCbs13+BiESMy865sYohoKOjLAhpNENsibeS/5FKkV97Ctcg24cikahwPgufYK9S
kl9k4wpbKAXHKed/Z8F0BwuYylI0yxKPxEX3k75fwCjpd+XFL0qpETsNQVBtEdTG
Ga/q2/JLl8BUtOjdw7iAvv5o513NviiqEePcuuoNsJ3r/hk//HVLonVtk2J48FF3
iwoGQfxR6cAQXJmVERxYnglYvOtwhBLmqMpn1hqsdHlMvkQoqb1Qx7OKaY9iZRjm
n883ykFEvEFGSefHfgOEn51phSzl6tnZWewsXGJzfUilxoTS8IIo9Mfxhsacmcfe
gyFYypdmf7T0PJ1NIIZxOMi0UGKsix7Abs2KWpcSKu+nbuZsplecLAqtKph2UI1V
YE48kgCVER5s3ZyvEYufTCc4+16CfjpbJaesx9PcEzERDOihDu8t+tG7/+BZzbeQ
9W6OAzvu8oGqDxZ7HIUfRzDuf3FYJv8eS4ba0tkhmMVhAzhjuOqL6u5aR/pCS99Y
avln6ai2lCjISdrIshzH5mw7Dd6LLtcTDhplx9g8JEEP5wW2rFstUF69etOat2bF
Pfc7/H2C2V0TE9pxboD1s33elDxA3jH7VWjbXt9YPMnGe4ZQzwEoyLg6UB5sNnnw
zz+v9rK4h1N/MQGzzYkN+Bgrq6B28qD24uT+a9+wts9QVVoDImBlznSEVAFfnDt2
9N+1Bz1ZL3UaJ86hPeBs9DMlkEpvifxxwNXG5e498nMX/ZN9h657KKwbQBrocEwf
0EWpy0xGBMFW2dnJFIXWe/7Mj8hGpQ2RhLtGbSB6cusdUJO3d/zQrB5wHC7YhJRi
33HoES/h8A2X2j+TtAn2ykIJgCMB6U62sYOc3WDV7Ypm1sVHkN0Wv5Fw3lu7b/A+
IRwhBlrp99c77Od3xz6VRoRLDesv1PuDeUhj01QOXE8Ae7U53hXf39BxzxVaacf+
7othhGtlUrBIt32Ibla28P8+1II1OypwH19OxXdZMuBKy74xp5evAUhGyygqC6gI
CIBfjbSkGeaGcJP5jQynZJcJKqephJSCZAtCViL92JFOXm29AldsiqzP6fJsKmhj
gqL41LeIqUkp3csmu2t3jj464IpbFVl9dFBRk7+2/uuB5GuwIBDPyaqmpNH9NAv+
bzNRficIImYa2W3WPOyyrJeknGQuoG1enRW5+GWf4hHAzGu2krLK5VCdBAJUcg6s
xgKhx+JrWSqGgvc1fSvn4KE3NgarbkHMQOMr/G3ykW3yJdOVMzXA+hI3cdTRPFIv
OIiD3QwRQV+1LUqMiri8uUhB7lVxBwmmP3/HWLm/uIBqrHsGw4OqE3iBJfcFp9v/
7wqT9a7Z6sUkKKsAOo40IfTBdmhxbh7ZlKqyJNb146AmwjzmQISfR5tBt3EujIkx
48uexM+GycnJwUyfdEnH54rYtPz9CmZXPuDDWrnlCsfzT2nhFCnyiqlZLwxSmE0q
vCvI2urmupO3s23Q5iD+zf1mP82EwJ/0jokS6bV7pi22AwP/livVKZsOEqT7Mt3H
7ViFJHmWz77kVlx9O5QpzPAjIeXo39Bp/4iq8JOQn6ym3ur+FTXIxKvFLWmv4yMs
UnoG7omKhPh9uXFsE/9pLZHNTWhwXAuPmD4s9P6tjQDSTYm26qI/LZ/HdXqP0Xha
9de1kFw3k1PKWP6zjeh2vGtCySXN538xQlz9vooobJR8OfL3KKsp2l9TrkW8P0Aa
vP3wGIoeLMwxGDdKCp+GTxbI9VRpMHHXacSVuHYe7kXOSX/s5zpYOpXmH00XpI6W
5z2unERWOndMoY+jL62Pts3fqz+UkTtRAFOIHzTDvaLKnOOyceDN7hcJRgdHLp5g
MYx/jxGS6cKAnPEwoJQyHUKm9HOrwL1/8LyTrIsJR4lsg363a5xPhrZkA570JgFu
ErmOTO17PNGvsD858irDTJ4Cobkm0GgP6FBjkl2HaRUCHoKJ+Ogpco7unatsWqz2
WvVMmDgkSunqoLnElFYlqCx/b5KcyfqST5/ovLSuIjPBKJ6bXgS3LvYgB06BpCCb
kWPeQCgQOygQKxldHZEcV5VZSOfFnBPrnsP8pW9ghYmz+lCONZza6nMZHabY5DK/
Tr/H2Bz1X8bcrXcN7YyGHJ4SHJ6g/V8nQKpW85Nwyl05LRDx+1/6TgYdRsh/2pkw
QuKCj40WX8h4S0tsFgBrGE41Sf2V9ZLLwWMsmqOwL/kDxhcE63baAWrA+0JVMvI6
IzlyTIeugyjoNVRk+TXJCBoqz/D0cGVvyu1vLKYiCPmOtvBqL+r4tc9Hy6lF/T7l
2tqOTbUdTXGbJlptpzkV6g/hjuSg3g6kDx5bsTS6b5Z4WeKrNUxJh/RH+ir5BY/B
Lfro3nDRAarBba5lchdjs4GjXcLmcO3O411XMVzLfJFYsH3P71O9xCXST8lxT9rj
oTU/82imPryvEPTxQu1+w09HSMnk3IB9DcQ9JVykaNmgAEISqZNaHz6re7YvfTfM
yIErApsO2ZCVdNu2qObqfLXgr6Vf96PeH3VdZNZjH3bSpk2nkJWntqCJcmUfk6Q/
kqbBx6uC84d25OV2Kx5Dn2OgFaXwSL0q4lvuG7BkRmZTUWINWwehQDY666X5B4Cy
btmcUYWmKJJS6SwwexVt5BGGsziN22P0g6g9h9w7eWPZFN3KNOeD/AcUb5M6z7Sk
gHGfy25kn7Y+zLidme6Nol5R+0QrFgFViNaYlYz/9E/zTe/IbsmzkYk84+ry2SWH
0hk0KClK0HIcJZLsJz/F8CPRx+oZPLy6q2u8LazR++zzji7BnDBKxTZPpytDQXhK
nRtW4zmz0IMhJWjQqsabWq9RMlEazS/az9DTNEAWvCsaZqdGwD4ED9XVYXtetP6L
mAp71v1QLozs4nynBFKUeJujpcpsTknapea/2ykEEVLXfbymYH6WMBXPQeawzI4x
VcsWlxF7n/0LFFuf/0ErEU4zKlXj2ayt4zSfmU5iDkqPEN/a+H9q7UAiGiiN2BIS
XkHbt/SZ2N/SHT+ur90gXjbIE7Gnd6SigMjt3f3+qNCIXM3Y8W4widVD21fyI0no
kCgOec8pydBGvSEOUuDQJyaWfwInIvYroi4KOdmJB/rPH7LlWo+kFGeGQLY/RskN
x497yGtzMCfaOMjYt50Q6nCuwmtnIw0O+X3RAFRrhefrIAUt5OJrbLVqKmoKkfzo
UiWqrp6sHPUAZJGkkYBNSFYi8JX8j9AmPNIt1mvrrmUXin8jZUY9xbtv0xq3qXtJ
09PL2+tuKbCvBOx6VYhYySjFQlBmUlnDYIypVQRig22H/bX8YypgwuIrtPY7qBgF
ozTLqFV82gyfXrkKGcOZa/Ymu8mvZat8AK5ZzGBoL5po3DATuTBjTLlvvekxnt3R
IStnvEw8VZzd0OvD13AvYaM8Mmx4WrdcYeX4tIIwBgPjrcPUcO7fDpBqrd4BN+si
OExzMv4nEOnHFbor7wjO/XnVdqDeL421C0a5g+ew0lwwS5NrWK6k3zk/mMmVPFAC
KJ0pZQ4zXtL+0NZzongzKZsHnoyX7K00Fk7lx1j2ebONB0hsESxU7j0in2DBTzo+
UUWGkV3UFCyGKa0bG9C1jTa/lcXlzietRkpvP0LPkWbZs9WdLiKvwvpeyQFBHOYh
hy2Zug3Kfgm2ZvL284yBFfua+aMvQydH/hoy6uOxUH0Qs7ieJWSu7oLtfr27r/bb
7N6S9Zrp29gKFIlWGutXQ5OcbFK1CKnS/C6aZgb6p8bLnTB0/hXyOxMTZjK7FzGh
4Qb2lFBmTnwe96V04dhOu7IjLMBxWKJrlbz14n8XlzNX3mlJCmpntkW3INl7Tq4m
uZyyRS4D3YN6yuClf+CBaJ1TIZN6yzOypxD6rKALeftZsSU5if4hlCbWPIsnOlv5
iKI5n3+cNUQsz1D+N9LWMbKlgrvNXPMOmcd9ayuoaScDPDiuw6vp0zzGWP48BDXw
Xoxttib/0KMtp/D5AtvSj7vULMquzR7PhaH0Lve3zUlXsXRZoJCE0cvSTf9tDgkF
92sNMVGk0ApLfWSBVjhkOeyMJB8QgJ/TdmQaFWQN3X+ktZqsTywvV6XdM0LDppVo
BMXx6ErFGwh9XQZ2u+xsLzBFp+Takm8633BaFGbpFBR/RmW/FfjB+WmWpLdUR7hg
KTiDbCFNdwKyw7/eqhgr+si4n3sPALHTxDEvcjcmTnHb/wc4PwCtU2y7rglkb6/j
OChNru5nQBEZPJxJv7JGz6TgnMwQLElFvQ2PDYz21G601dL8ygzzGhZ8NuCALeHk
B9+QgQ9JcqPN1SkOmJaHClMG07xfVuommxqqGl0EQSg30Ga2fXIqV1BGHc//ABfC
p8O+OyqbuyRWhDOAS7Bt4sTgXC7kfi+KVjc5fxRTRwk0tnd3JMURp9WBj5vDE5uW
+vAH++6GjXBMPgiMqMMiP8120pLDSaVuD005pgD3P4MQBI8sEbEg6WFWZwDwcCix
tiEtutXfCQCkpyzpBo2SCRNSbi7LMM62iCfy73twGIN/hbZABNHagmtc8dd5N+sx
iGiiLGubJ4/duxTMKgVH1+3fW/lX6MuGjgcIERITpD9uz8jaxZ3HqMyertGZqswT
SJEOZ5otTlyQPQqM4QD+p1UTQSLZVNOrUtoFwX5mmmrc+N/hFaPNdUsVIymUyOXK
FUOirtmp21KaOCXlnDTfigYg3jxNyqKD7+GdyWqKBhZAGPyvHyi1cF5r+D2GCmo3
0HhR7cuCyW0DDZ+QQZ3CC4lVqJfUUwsb83LIaqYjICNcRE7fpsc+tFaGY5lsoXas
7BjEhE3ZlfqbUARKiHMViaIotV2GEhDe7UL1dXkGbCkBfzwu2vGRleVKDRumQfMl
0zrq+xU0ApsB4aeoOaHWQ8Gu4iAOQXnd75rQqXtiVHqhXZEesRP/I5J3pHxXGEFR
4vFXjaAcPK2wHhblJAs3qDgc5LiGWeu5au0DkIYi/iB3eBqIdad+OWMZXHtayi0e
t8HCWF1nihJ9W6i6ZpG937hqF2v8gaabxIujRKupFZyjJHVSqXOEmaPu76a2lcgS
f5gqxEjLjFPKUMr5/mqJti1AiRwQmW9emCwG3AxXHSoHkZjoEZhR4vMJgpxa99ny
rdXZQOayz+728tGcWiPKwb30d047tYueeE2r0/xHYcxVLjCPBGkCB+4i/K+KoHc7
f8loNod4TuvfiJKMuVDC1u/VrHUX1+1ZrvYQ/1t9fCmD77ZOwlYoReCPfomEfYvC
ioMz/kUFxBOF0gsxjhKThg+ny8mvl+Ux+y0d/6l+z377lD0RRyNJCx3v9smtEF2Q
I/8l1aFv5SrUapfWxe+UAL1Ji5qjd2QpdFI+NSsS+ZQmgUgPrf4wjyqXRuXjUzOX
n551Gk2iqMxG5H8R8yl94UlpMFwWBAlKHLnmoXfP//N1WgCfn1/eJl0l71koulOb
9LL1m7vCzo2YcWJQ41Bemu5fL6HHxuIiTc33AJIKYgjjH8HKOyZ/mkMyGlxSKWBf
VuhLPkBnsHRQsQ95mNgSu71kdmjPlAiiLhcam7ksYKnrvue33FrY4gQcOreYyJnX
g7DFHdxo6nQ0omkBLqdiNoD0j0a0CYsgCF/CRSbRKl/IyEgFSza3mYfvNRxGI5+G
iXNLzUo+yBjefwoKiW0LeHBdjp7eE3ueJkh9JS9OHtxmbOAbvZEZSyAlZgLNmRhw
+BGBVhGqz3RT8uiBnWC4kHyNmmKBNh2O7mGDTDuEpUFBmKZHMo3V8DaNSd0uQfxC
QAcTgzK8R3GYqarGKiHidVVm/oKzEgoA00Vc8A92+w5yEmw2IVLfX379dbg4BLiw
A4D8C20mxK3pRh5MO9z8rZAR0Q2BPPHqLhdjcXZ6tRn/CxJCFui2c5Oxbyo+hDMk
Db0hZWR7NpxPuKKzx4ibl0I/6mCTzXbgDi9kg7jTUY7WerqsracgeXAq54Oc2ubr
9N/oqKptvLj2283mUaw0lihi161iANksNBWcX0x5Qq15IJlJJDSr/YpEmst9UZ46
sQeI+ZDDEwFCUgHznfiKswnXdfAYPqkiOUeKoF3Pu3DtRsuVLoES382JRnEHej4S
0lHieGFO3tRfC2MqCXYI3Ao1jaEKYIlrSn0SJa+Al8gr0MEP1sWC0vo2lJrP6k7M
uhVqPta01C/pSsJ2MVtCsspiKaVfXbzDgXASQaopr3TOjCA7m0tmSXcdYU9jzvKT
fGGqXzrq0vOq+Z8/VPQY1M4xjM63SoGYwkYR4FIQH2Fd7jZKtiepNJrbtnchEKxm
V+bJA0JaKaAb54X8hO+HrU6BrWxbVqVgeJRxiW8BanyoC424H/DNi7uRBxB6s4Zu
2KX9i1MkMHcHymNZ8tF9DUtMcT+62OXf0+H1ELbcNdvCfkXB+gmRSgWDcCmUgtgW
12K5ZzaQVEQAac4lGADi9utTm4ap5yhIlVE8DXhWC3kzX7Lvyug6WSJNMnHH2P1U
b1v+ambJbFXUJWGNCHL4dWecBWjSDfxnO0BExOJc72xCFgOwyXkWK9TNsJv5toxf
v8gnVS1vab2MHkSsQQYzDMHNKggrSp9zY24FrGeTeGQqsG0w9oPtAlVywA6YAoNo
iklWBG270CBIWdTigX25Swi6s6d4HwecZ0QSCifrGwsxlwrvdg03oqXii7EA8Jwe
79cUv+Yn6zQnD9SOTqb7Kq1ErOlp/DWYIYZGxTeVGB7LcPrryv8YbY7I7AfDL2PK
ojNgUK8CcMgV1gT97Gny3XUv1EKdqYHgvj5/c+Cu9+Z2n6ApCPp/BOwwXICCbL5D
kQwoBqyz3IMBysFk5dGHP27JdA98auzKuN1Ez2MELP6lNknJ2XkdcJR1XjKYlnM4
+p2IO1fcYl3DllUIPYk0S3Y2VswOgkwYdZnuW1XlgCFoltkASHd4I2W7c0VHgm5I
AV7uE/PbpxciMiYQMwlY1YGXFD+eq2hWcbuMWPxoOf5Uua8C3JVkPifWyCKhCh2G
NyLW7wxZuQoo29cdU4qYpSA6Hak8U58Zy/9lIkvtw6jXRSoIe83qyEiP2UVfBoLE
Zay2UpbXUV2FvHgOVYngsNRhsppV/CWh5xUO8rR3hPtg/nCoGFIoxhgucw94dIrU
SZtOl7gLVq4vEO/qNajr5Dvvq85blVY/mCEPSBgN0HqWm2CE0ptOatlhY4l4R9Ot
sLS986RE5T46K463nYHPwvnOKatZ8baEQte1OhV22bYoe2RBo8qPAxLmRKnfz9Uj
3UJ6kSTEquiSpsmU16cCqUbe6xBqLVaOVgC0CPQ9Dh+rKwoP2LlDlUWh507qP4dc
NxfJVOzKBOn7NFlKhtj42gSreu1rSz6EPY3JwcvoR/cctljVY2ZpCGtzzvDNJgaa
UHT6HzA9o5nXp7rz0lQvUUPmP/7i0/JVuHtrf4h04VC/bBDNQUXRGCMFKXZw+j2j
HGfKu3nNirJBmDDqfg1/wyRSyo4JaxYwuuRHTsoCAJY9Hui0KrkrrWqqDzJhE7CA
ZpSKDEPwTVUzd7K6Ci8CPTc44fqhP0tdQayEgjGhydU4RO83VmjX0Z1bHFMHo4a8
P9g9kAQeKgTE8Bg6NFOp7FiJbaqo4qbpHXr13W/drWvxSxcQ2q3f8iLHNnPOZh0o
SS61dWqHF0Ep0Sb40bnRDRLvz60koFBbT3eRCTf78INcftAzm4ZM1DP+MBQzKMe2
1LD2SReEMDwWtK3bcbwzTYE8axl9EweEtWL0ZAtKTZRuwqeFTcYkOfyYGJyA6q8l
pXzcNOuDiHazBC85nXGfMaKdf1MSSYlv1lFwXen9RFgh/Xgy4UBMObcLNEbcGYON
TzwvBSBkvVKGU4RHYAk0hcyyz5TAWDdeB4yADoZNPQCBfjLo7d2LHG2RA9842lD0
cYBXbr9cgnNNIeg6cY0H/WDEGviBsgluWB/r9Maqsn2MPFHBrIjpnAfBKgh5M5y7
QhlA8Tegj0nUx3rQSp2mtpiE/dJKVWiO9A8BMHbKhecRIarz/nRvRsIinN8NY4lb
HEoN78EdE1b4MI/i69Xj3GigJhIko3Vj9wZz9oQXOqt+6n9BvOTtNRRFrzOZD9zh
7bA0RQKS73LqLauWbLwnJPgVC2Db3DV3URbmuYlqZP7jfSyk+uuLHh4ctcX3+AgI
yqRu2ynbW3uHCUe4PoZ/hfqtN6yhNkCNm77+xULBI3bgEQs65mYaWuoqWmxhXIoL
SLfqxQtnTOarZ39SkA+MjxAjQwKJZr1gosSIBaHZ/nVO7Ufi5YurZSKNCST0qqF+
oSb+wgK0oIRA3P6kML1dBF7K7RWuzNJHUpykTfarMtL6NYaLbB9/J0PjR4SDS/a3
JL4weuIRdIzXT4OxGEuGWnS+I24ojRetZquemQHq89OmIG6KoUcrpooeUH8kTcoX
6+MP38QA5olx8eVVONaFBIGogo7405JoBbZ1jausJv36FB7llHSHJV6q63qttzmJ
d4wJWFRgL7AXPEBHQD0RqohHMZdg/GgK5Yp2aCD9NcyyubWDdlNFZI18GQ6+CQW7
5OCEQz11Puv8VB5Rnzv/648Rro02ov432mZXXx2gSbBufxs/rzDgH9swKs8fY34i
RJPnaDhCtGr/YY4VVkOSHriXXY236poqQGNKZ61TqNwm4Gc5p42Mi0s2URC//1FN
LloNBHOl0m914d7ZUKEMUCVQk0QNNQi4EMRJ8uCDEioN7qNy+Ok6SmqxYjNU+F3t
AT2uACSduux32boa+uDgdTmDk/Iihd7FTS9PgeKYVwY1rwW7n8KFq4YZAbu97gYw
rBenbcRUT2/Z7pwfmAEQbU6Mq8MNX88ZSfzMxfgEXs4CQp/aAunoADQA9llelqsM
iCGhmbJahPh7Tq0UBTYV5ZmhiLP4s7eAtIAQRRVs+BHiDKmYxg+Yiehj8INs5XAm
7g5Pa5rkLN/JNUDiNyWvuCI/mnFyuqIma/65FtKmXPMY1G3CY/Bs9UEGgErC56Qb
/IqGiXRJRUIZ5IzkClCkeb3w2TNa5mCirGjszvcrQG9l9Gt59+ckaQqWU6hgfsKo
HuSxJz1gOKzyW2DudghwbAumcW9tSk7ZoJM1ldUrDhYAXDwlQzSFKHOVDKqHa5Ca
lObRQBZzVvlJWORdxdnP8Tv0ScpuTCRGk6FiQOmMh90i9YlwZ4Tar6+NcO5H/wDA
5jpNwa0Lpap547X61/T6DesG/99yUVPh3E6dJH4gsz8fYO7nI8jWv68VitCgX30E
H3NAHKq4dym8/h7eUOw61zDa7zmMNnJvmjhUw3QsJSOPgviElvmbWnX5ZQf4z1ZM
TaBkOyVXE5VknsB7AQHY7EWfVvFOc097rLH4PlV662rJsbkViD+DGkSTp1MYM4cx
/U2tU/PLAGd3YT/2eLJkrfqWrBv7pljUs6/TGw3p+rfQGc0rLbGjVJ5xZgV1HZRe
MxwN3My9x1vsBjc8+PGrWi6ncceanQjuENUB0c+id/YDLsAblFATifDSOaNx9SJJ
IWcplTsLt0CQkodipObWiTfFCNHNqPZzlzfJWs4jhB89iXpTddTc47U1Bfh/U/lz
yP7Ie0Szr75eEVAkrswOPyD37emJddLoHmJmyowHbqlxRTtAAbTc7gSIbg97FNSr
NYsh1WNEfsyzxj2alZTXZuxzlprpf32R9aU9BFI/xhgfsy8ov2J9WEYf6cWpti2b
2+e3w8B0GkiewyjY8MHEuOJFffr4UeHvmB/uBT0EA/CNYNE6DvZk+E4w+KMwpqW3
PL4bST038b1JTQLqQeatTu1eSnZ8gPltlOA2FKyMvuUi2bb41MMhMvIBMgjJFCzg
9B4mUnIZO2Lh8ywFQ5rTCyTaBbBeYOMo4ISjIYU06Rf6ypfkPbOrv2dgdRFPh05e
cOzdWcZAKhbXxIf/eskFDE+TGr8B7WSCZVIzMq2EIjQc9uSOvLA1Umdk16eLU38q
7/W8P3x/6Pq9yB9XwZRBD5OYZ9yM+SCdn/Idl3CXpmjSXXeb14ODeNoOt9sMTp41
yVfOnRTV39kwp7k8NQhDqtfhi7QJWzTyRSFCrrMDofFEtnuOJ3viNveNKkUy+JeC
jqMdJDtR7Z6qMX26aoCb8Cg64w7KDwTYkTqwcJK+txEWJWrl6JRMV41gp0uY5l1G
MHuENEqQ8TN2XgSM3ggLhx6CUWyGldUdDoCiropqhzZR6zdusZhq/J+aJqhAE/K0
tPzFL8tyci09YsR0k47BUrVs9z+4dvDKvmKd/3uuJ8fa91TJl5j6mxytwt6WlPsT
KCxxEIQ1g1tLWGuY9C1k2DPjaSblBkqrcQpmuxFWlFirAUbQTdYBGh1UpP1wqXRt
f70cwFkSCP1jqFdm4bTolSEc6i/HgKws3pgS3ui6dSuPkKkU+0jzVs95g87g7r0D
03n/if3o1fhCIRgToN/AnQr+TxYGi0WE0QY86RTWB3IUQio8NhpMEjaZoeyugGPu
LygjOWVKGIvdxi6Bsixr26n7VrJjWwqC3G0i6nfGmGf4hHJaeQesUXYXWEap3xGU
IjDgreCoR7Qr03o7iLqj/AbtFF3BHon6O1CG2IiTYhZHBW5hXVZs5Fa1SqPGXnHw
GgggPxxxZLacjO9UYAnr+eGOaPVKrCDChhzqzUTxTlGzp2FX2MButFDUMua2LrtW
VXp8mU0u0J+DDsFHvImifQcJzpJIFTOXw9lm4LY2SY/A8NYyGtu0cGXMscoGrhe7
feZVI3xOGGIPDAQKg5agBB8E75ascQKgtVaLmsSrNJw0bxzTJ+tmQUo6oWo5TGQM
k2KhHfCBex0iXX8ugO/onCc/NABaXaTkc8dwWFhM1qETMSOmdfYi0pJPAiOXwRfB
2D3QaYvp1IIweQWBp3KbtWcmB4SdqsTyljTCrSRekZsPsBi5nCm5qVd2f25DQpY6
sQWwJ7mMjW2hQczH4BHibFesrSPL5o+hQtOG04AfT4xGrz0wRoCErBO0raucg+Sm
7+UWiZVlc4/wfHLd5TLRv5049hay5V/MoopBIGCbRdq8BPuY+r9aJtnQ9GhCe+Rn
N13pScWvg291TJ0m22K1qxOkwe6+iMhI3oPnlRxOEePVCb/Lyn942jpy+6xOA0D7
ErODnRqjUugsox1EMuCf4G/kuKT5NDQqx/vvA/XYGIhzmqJWRLrS7tXgPKS1KEYP
o9NqLy1FYBJWf62bFMDHtlfr5/u3kzvAzfzsDQXk/qLj2h0eLdtRrrqSz5l5EmS7
O9Wu50ClxsUvUBSRibZznytzIU3Vcneuoun1N2odW83hoU/Dj1PCV4CLqCb43mh1
gspk/nANiBej0q2j9An/G73NVtFziIVZMTdnyzx5SbeVOwzyBhJo6zFqgP6TjcZz
AmHfmZvilnDmrcATQ19T9ScdBPRwzYULim2RUQFdE8oIEcypg1BoIXQ0CsYz0wCX
skY8Ky/KlxK59dhXoUTWyWSqQUAVlSp1NXgUChPNr8/l8tOrf1SmAu4onbu3eufc
ivL0EozxUF5Hk7hXL7o8ZH6G4eF3Nf4IBBwZjJDq6s4LKgpZYvZ4rk673O/bwHZO
9U41fGFTu8EqjpkwMUseP8NObeNw/zTYJtLh4DdC12yWl1v8G4z8zAUh5HbFqtCD
H+6iK+OwPGANHKDnWR2uHsKz7YwuhLBjr0A/hpge/JwqU+g6a+PAqt5MWsV6aVNJ
vF8QFOCDzdPcUYVK1AUBrjSJTAAIF8TyV4jTntavBLzyIHisuQYWJIcB2UyEyGAp
OBTHm4mcIGXLQmBNoLWO2dXcbBKVem6oukstUywDwYY2d2MLq4TzlOBOYrmFuZvN
EM3p3Fcq7ymW3GxToxVuYuBi1qkB+ZZ9O/zocEM2jUmR0WE1evzfVZHv23HjD1UD
s+eXARh1WJOSVBVJhKa4jbu1MB4F//M41ze5kemVbQuBAOlWzXXDU6LTHoY7SSdj
YPYgND/+PFSHK6UzYVjUQkYLu9T1k5dp/holSUzl6C9iWSrZUhCrZqje7agm8Lfw
kWS0bYnBoHUtdA0qZFbgYNlqJTjio6+KjGwxFfO7o3ydmc49bS/jliC2XtC1+pxB
dO6rXwJrsvwiyLgqaStb2Gof0Oj9QCJXkDNBcm97nA3/napCoJuk++pi1/q9WpYK
aVd5SFLirC9HxPrCTsxQj+5Skj4M0TLr3gMtDNOz+hY2ismgqauoF/YE3oevs73h
RLDmlrNy2GFRIYW2/Jx9ccvF9d2lWNS215i8s0pqfCA5mwP3frmdzsECD/INxHLO
ldMa03F8R/42KZ4H6zH91lwc6qT+AtURqWWZyRs12eLCEPDbpYcRKixSxWnf9Pb0
6B7Vuc8NTVgAgrE8lTL4sV/oY9XfkPHDrzD9Y+tlrYS8Gv35rQivDqkzFzfcgOw5
Zn7Jfm2uNQZHWQREpe9NBKZQIwHZvY++4wgij2/896AXubUzxeW/MUNuwN/J2y6u
5UCz4Fo5KrGFbLJ72R72x8VULgUy80s34xyzTgPMi34aHlwHuBYebP+vG8lZqq0p
Mc/GmSD4zfgkGJJTPJCVW+Kke/sreGE8fHGJ48AJlGhear8NgGydCU1tMhiJVaNd
FdHONW3U9/ZChmub5TorDYIJIA397cVWaRgSDUk6LxD0K6W4R3v6fXVHyugPhYTU
dwMFqD24qa7crZRO2b8K8ep9IaTvxHYDWRpy8/u9p1GepHPouE3P64OetNxVu5m5
JAXjL3dchDoMhOqWam9hFj4EEJ/tQJ2qNSsaTaWgYP7Mq+vGAL3iDcwa9ZKxDNjM
Th6zvHzJQcHyXFQY5VRo0A7olAGJGZqEXTojJqAWfTjBWSJo8maDkaaYt0OnVkMs
f/IBJlYkgYgBZ+3vG65LWDxqLA1M+CgQz9rmRScmUJ7Da0D39tOOnm6s0ugLzWvs
M95C4PHzczFJyjssEaH3EiALfbhcnrml7k1s9jyc49n4+JxO5wicVu6VKhGEwCj6
/X6g5ySJ4fq4QB/tS7/fIVqU2tB42Tvq+VlXeyy+3TqWWgyd6Vcx6DhpDfuGL+KI
7GvaUwWk6/e3Wg8zsiN7wyyk80EPK/YYse26eAB7NZb1sCPOZWYUuKLPt3OcOQum
2JZ9WDl+RtBxr4zAHubQGLt3NNwtEWsUlfupFtt0E1BVuDpBlc5irMJt6PkEhF6W
OEfWoLGSds5/lqWHqq4nA05fAZ/VjwbzSktyXb2N3gerXdF2JMji43PqqHo9czHD
thX9SSUXPktnechkkiQ/42gbv67XVcwE83gHSSMJJkdHsnKGnb+S9M2C8aTPAy11
XwYYYbfNQugHjy0rzyIbelNlql5RRu4IbKSCX9MTh3WOdNo2JjsN9fBWwpChyPo3
w3NuzyqYd+uyNgmcUfbFEhol+Ez/HqhwdglnCPYLSHxko83UXO/T2FqnXc/iKhdR
/WEci7xapWpua0ewHmS2OTmVctYqKXQd7568ntWB+GjVMGow2QM+RUi7+eA0aeke
ZcsB5Fmxasw4rypdesEEmoPH05CIU7EIE4EMvBnTVKpPVBtb+490x4JjVUrcJLGp
0j7DzB7JEDF4tQLacuyylJpcZrEEfvEaCGISiLOFw3lSKkESkgAxkEeyyZ4NT2kU
7pkE1/z7pnqyBRfvKztZ3P70RCdYJ7GZe/Xu/pZXwuVJQJuwrgeXik+eQLlA+L8/
OaW4lq2nsrKJGsQUvuSKKvni7112uX6VvfHSaMDizkiTTWCISf+QCHvi2c69/L1I
78C8yJ1TWyu4mQNCm58nhjuZPQh/mJMRIQFNuM2kEe/R/r2Zf0gJBmOhhvqGTL8n
IgmfJN00IZQ5w/TUYsM7I2eoJCWPUU65ankU9/nOBsx2rzmAcIuoAI/kvhziTEav
IpPn3J+roskgqm9T2dOAj/uUgueQpFhkor6Q8KWtMxo+LuTIW6vE6DSGe4eDZR9b
j0/0GjzUmjb9YrScOBEgvvpR6/lU/Smu6efHaCwh2Q4NuzDpcrdzEWTgZggzCnXr
MxctapECJs+vX8b/p2YPrjmvwJl1B8ToOlh7CYUx6nZKmSs1+PrDX68IcnM95ZVY
8+OqMeA7l0DOc1qA1rs0VtCgpmN4cqahUea+5CpI+dU4aZ3rPj1PYd9gfX39+bgK
qxvt3ENt3gQQsZn5g2iw7QGRgp6UjedRA2qPz9AxKwicCUqhmZ17g0WW6fZakUnC
m3if5VTqL663FkYG/WZFWUWbpKAxG9pihseb1wNH/aLI6cZcWzFJeRl7rbp3qGKQ
+VM87peExbuDR4UBkzv0/5HcF+dJB3ZhlnHRYm06vxHtvHj07mmmGWoRQYBQd/BG
YXVSPg73ZekyFhkcpsXINq+bEovwYTe5ThzDvUece9ysmCFLefdMlX8gSLWy4l+9
JAWvaVKgvU/hOCWJESj4tuIMeYTpbtLISKbJm7wV9Qs7o0O8kbH+Oi+okese6Sbt
TqEDbt3CTzmTV1dDXu7wI9rbDpJEzRe0+uw6h/zZdSD0Iul0Ruf91M7AoZsmhHyI
sza4HayD3CUWw4SzUUMuk7W15oF1oMnLuHcN7kRU7w8AOsXD+Y+Lbn6tj+J/tSGO
6LYCmSZrRYvJuB3loKmw67i3/cjBBj3jtv7Jwkqrukl0ZhXLFm6x/UKl8vsHqqmI
tPim/VxWHT6F0+/AtsgU5nH/MzOka2t9U2ImnPOs/qvERgaSyXjogZ81Xxk41NE8
no6xEjchIpUE3yUaHpvNWUCiNpUo3ANt6hTZgI6vzEF/K06GghZ7n0yVtUs6HYlN
n0GXdApsViaUjhtYTiE3oHIn+PQvVLYqQoe7Yyi7aW+bAsF7ImbL/CdTeIxQ3pED
kYBV99rt7apTzJQYZeAxs4JIlLPgIuELXYTjoLttDdHE1nQsXHSE+R/nRQZNyq07
aQkg89WyUBbyweo2HX9U1xxNhTt7TDH2Tht3BNl/hSfaxDujorpiHlHiVXc7EuFy
FAjkSJzuY6wV95B2HvUMOEITrx53OiDxK65I6mqENk+Jm6X4k1UMpBuUEk5+QW0Z
3ZSaVr5h+fmvem0nb56rDp3Lfq3a5/DtQdA38fdS76hFE7qmzSuSEmFfEd/RPGR1
hb9GIT0771+t/R1LtkRifoAvJvZ1Dczcfpwa0BlY4i5rgZbr8lRed9Oqd3AtTdRW
xZj/t+Qu8cqhy23zb2EoKZm5EvNKKI4H6QDdE36T7tCZUQcw8beKs0kAebmXFRrA
vb0SX1rmKHRJ9NzlW/TBFW/MDZc7AnwExbKvuHFIN0KAzqgysN7aLEfp9g/mVvIX
wSEVYAsNMUNdnKkEc0L6T3QdZNMt3ZvdasmkfFsGs6D8XvoWOOir85Y3qMMacZ1D
5XHVIY9atqJtl9GweZEara1gWQFPGktTrjAjMeUjZUVadcnpZwW5R1Fdp4M+Z0vE
Dd7RowOAvrAg/kaqRbDzSVr26XOjhloVoMRnXM4AG4nxSanNVD4TGXlSCXcmFr++
riOBFr18ltRPC80fJozYbERKeTUncxjyJh+8fcgay2VK5b0Snxs8O+5x3Bt662eu
pODez9vEbxhHKgUsM3SWHw==
`protect end_protected