`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1744 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
sD5jeIt/NS2+ECTgxO9JluLOTU6i8aWefJdIhSEr4GLadlfhZm9B9mRu7PNqi5FZ
R69rvBeteYbwvcLAQZkM97A56MLVyBQ9/IhrYMM0p6KOziKmhpvmjvaBE/Z3poBF
5naPTeAfOy8UFoMxLDWS27J7UhQfDvnu4BZfwHjYqsOGqJoUC2DR/fFMfwHYeUT7
KRDMkr2cefEwTUNaMXnhl0ooRXZA2hi4XMI/9L17apIWrPR+i7HLzUVo7XvSYqZD
uNXzj9JnA6eEJfzivRuT+zXIKYaXHtj7fN6jO+nmidV7F1dIX59O7S31uFgVGQZs
lq8sfNdkm5dbSUPWAsEA/RUCermrJUYRsehSheWDh/yy15V953atXkttV87KbKcq
qPd60h17uP0mTzsfh1rNA7m7O+1iksyBcZIuhU3rCDjGH3As7WU98OlMzDh6inS6
gSqTSx7jgwb39OcoHzmvi22lQ0HE7IhG0x0g5pa6YotXPXpkUzPaP/4whWpKjjQU
a1u+3j3CEb6ucNWdZB2Vk9tdJQ7HuMKeW+vyt7o8Xbo8rb0qcg+2ERCI1uLVmubl
TIKbi23TNiwuAPXFq9B87VbV4dYSyCAsYSFkc4SSLdVwX6p9goiN3D6/l83BwKu+
V2lx1660L5SVDwteeVaI+NHIuwecxZexqjiafoxDk37PdyyvJ342hK++c2rK+FDC
x/oMuTN17NvQNu1sHrjhBHojn9P5RinQtEn/R8/Iu9qI1sCv5EzacY/OtxzTmNmn
6thTolpahMfdZaUukBge+cPl/P3M/+rCyD9Dx6MwG8Q3wamQYd3m17iwyqdkhm2n
jh2Jq4vSMtzD74P/Izipq/5NNzsiSVHdNZC7lAA77pg0ridU2OEdokGPCYd1FkEY
C2VcWkncIJWRH1RlMHlCqia8wOj5AVqb7W/9ZhYuQ/29PC1Qc9kYNhKNKt1v65N6
k9nizScaf7TjUSYotP+dWASMKftcNV4vRrzoreFgszV3WX7VlY5U3C4jWr4EOPu3
BJX7Mh9O20fbNZLIajBRsxHK0FfBCGINaiETv1+fhC6/FgkU/iIuaVMWSnIcDCU0
4RXSUMS1/ZGthTLV6ro95t7CRt+fsFSvvr8c+HLRCOkOjAncXGnSP+xLnQteR1AC
WcZIssJymQ+wZ1C/nITe+AKaPc1KxO8+UmUifWvhu/ymxafeZdGfmJOV9wZsY1wZ
FR73rq8Iw0NIzLbFjAjtHKWMFqEUQ5l0an3Adv2byLYTSJpRUgqK5uoXnLeiyRYj
IO9oA2PQWE8S9TRyOlim0HHsjdu1kIpXAyf2vknu434zjh6Km40PVWWx39jslfw0
KDgRWuepKsht/gHi4MWQyUyL4ZQVJH1gPz10QhIqZ2DQfyPmkCgRmFJQrgksJvre
L+/ETI+uti7z3D3wlQsaPLUmMr6w+wGDBEPUZgV4ClSRb8CffeJgkdzaD2K7JTUD
rws8ZuFyfQtTq6+ndSIW9GkQjn0ixxI/70/xezpcMUDpl5c3S+OS55W/rHffDYKW
Us9xSaRotLLeo3Dzu5elwayY+T0KLYT+CWWw5lD0In5ronV63dwIjDoQVReWdP72
uNnUO3lu4BNw/GXqPcUlvcz/II1fvCQKnVMVUVWD77t9/f+zR76iSJ96guexzb8i
/7S6+cwLMkNMvNnuVg1+OdxBtCzHEXWvMT4U9enfLAn6wI7/sD8Q7xyTXFCQsXbh
RDQUj94cfrfOTA+5ufuanYGtApiIJIeLfkHTu5J56axxRK5c7rAQy/D/v3GoC2GF
SN9ZY0f3lXcOKIO01w90KcEJnfzJLauI5Z8iP9hVT4XHx+RkU09N+gNiNeDSBmjk
4wv+QnJ/IBaZEG/4V7gQ48nwgBaR8fya4QF93xOgyFtexDclfhdVoSL7SFfCqwjb
dtf6p1xNNVRrzw9yyQj+x/+eTaaNZr4xzn4Ei71wGM/1elhEMn1eoZe3rvzuqJ5C
dh/ukJ4yNrPOAw1FlG5kbBqOq+aeg54u9lOn7jZ+bOtzIOTKbmsix8h8pgo4hBEY
NTH3knxKMhjLehABwRwjsXGSxFTpfZvfhELRkSa5MPY3nbMe+wW5R13wnp3+jcvT
0do+YzChAg11ijClA4vC0P2qINJDJlfJ+Vx5ac3+KOxzab26wd4APYg/tF5HNegH
M8VTmqt7tO88gd4DZQ/34A==
`protect end_protected