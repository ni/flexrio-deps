`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 19632 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
VKWNRQF+vfUNEEp7apOJOSVr78APbBZ9xN90qYKa1P4FxL7elcYiA+D6ZOBLd+xB
iEpbR2rlR5gpssiHv4YbpMWs2BHke/pZTo7nP6llGI2MAM0mJLlQiWOWWgO+0vVY
N0CiEtGv1f/WPksWiD/+PzpaXCPD1hW0GWPAWItpHVflsKN0XcBxTkVkD5pIJk55
+W5mUkG9ILJX8znp9YGKlv05dFgV+zfbHQefuNfqql31O/I7emdKTIbvg7nygSoR
iYnfMsU75BxYHR0gKwCT+5Fx/Vj6igw3ppt0GHBQ0uOjS2GoLkl4XYH+Daaq6n2A
v+iTTUAHdxKIHqRST9G/lejk+QNgV9m6RmCslrK9mIfkUKoCzEnXsE1oqV+H1AMq
RJcCJDd9YbVYanJazWj9SOhErFzWgrUzrPHff6/WB7Fb9dysxzmoGj+GYVbJ0RPd
g0NCBXQsaGL32xTbsjUaroA4sLU6QsDXeJQWsh2I1+Af8pZPziSp7bwlt0kmYWPf
7TIdJLzccr1nYcMYAVxLNnTI+giMjgTOKcpy7rUTooX6yZEOE0Ecmq7N5v/ERlZl
OgX1rdsAADjzia7h1J2gB7KHQxI4C3HYjW7EqdnzmZFcn0H+uKvUKbpAn9mf/DiE
fk/Fi1UJveITxRbksni57CFvdJHJltVxfAj0/huoNRpUjRlnyHs3lGOzEQlkbr+o
1nJMrWHRgSVKQ2ZpCUN3tPoIichVNidSqeNftgu4LSpraQyxO3HdH5pmsJue/g0y
2tgzUQeZGgSJ2Bs6QMHnfBVEDuGMB3/Rfbm8uUop5tvHdGHUMrjZkFSQG33Zj9X3
2kSodp+susmRGiLHErq3wMfmTSyCbLOJMFSqISIEdhH4iXIYkx1ViDX5NJgvZZHc
UPCJKdLOyQz/QGhIT4rA8h6G2hd4TcL5aGp3yqMxmdirc2hCiWk1B1jv2udBqO4m
Trx/qJ3k9hJNxrW7xEFuYkUn3tfiomAeY3vUWHNV/k+czdxAoKcBGV42jBBllrfu
Mc9fvbuJfd1fOrwq03GVZ+JBgho04MvuWGVyZvmb/TEnOv8chWU7PhCP4Xp+jYTu
OR2548qNSzZmF/3secVOXjiMOYZj+bTNNv/P9bAXG3Di4RZFc3b/NWfg35c4ncTf
Y/AYJSKS56hTHmrK0fEHJvAIAKBARAezHPLRskes843BfKejoLZ6MIjrJQc7DQIn
yif668f5CmOCoBZ3vuGNkP7TgDWz05x3UxiJqUc7VCFs1jPE1dK+EDm2Hztk9WOx
5Jp6uO0tYhKzLOl7ZzKCZZo0StI9FtTTvfwWJqBQyx2MFycBnXRJWmGyj0TKJbdt
JbdY3tpH/EYOTwwJulvOVHO58DMBE7KShBzhsSBdIfljJ8faWAVEn4c8QU7XAqXK
yuUzs+1ZuXF5AqLnhJKzCzq4BPS4fQAy/HY2ay4Oox110erNGBUbp6pRhWGhMRzW
/doNOQNCOmLqBmyrkF+WYH2YFajCbQKLhRjtLwkBci6UTCqQNroggYYurkPBPysB
/rJBHLIt4yTD1BBRxmQuYVNlm/Oppr6NvJhhJoufUuKcTpsxI1xA6vLEPsM1DSam
dJVlKxZb8cForiM4xfm9XsrX8JdE0joYNAhJoU3baP6b697G2sKatm3B7WIWlDQP
Qwxu+xyL7rju80lx389jjEmydXW4OlseddAlU7UVTZAh0OTx+4Yafqcv6LgzANWX
m8sXWeDNfnCZdWVsFAvHlIn3NYisKa/aMaYYDdRaQamIqL3PLDrEBbR2jXpiRpvb
eim+Ch0ip6/7bjoM1+EhyH4GKzWvA1jnclELpsWrKsHeV7dl8+zBMBvapWF3kCWe
8wFtD80YVzmokJmhj1yxmzLL2rZmiWhTcV9JI6fBC7eP5+n+RaXr589rGlqS2oI9
sdj/CIfol16OmfLoYUQQ7mB9rsVyER9RWsMsfPKMKbqwwPS4A7gi08NeL69/f7G/
OCC45m/PqYtmI0r1eHKEP2PMtAJu6axC1mGi+FDnDwz8+VPYYzYOe8Z+hJHQ68NC
X9QQZOGrUy9JoFetfx++quyzod4mx5bbBCg1kmmZPyOKkoWUZ2/Ghaf59T9p3h3b
ZWJS15NK9VtHam5T7gF/tXdHNyqpe9Yz/jt7WNw23NcqC9at4g3vAS6CnRF+ee+4
cJnkQkARgYPVtlZNjrKk3PhyRHKvU0LS7IY24HgIuUr6prcbGj5LKMdqBbh1rTaK
NwZPNDH3OVqUifku9SMjw74JJ9+EXUV14QP4tv8KW16vCVCTVUQBgbyNIXrk1Jfn
Kk2Ta5xHaY3gCywACYzbE/rlXPRcnaiv5twdayI/3HropSNdDhjO0BQqYBMyFeGc
LSfy6/BghYtbhCA/3eg4+NGQ7y+VA08iuQWao05PavTPsIbqJZu6BR2sBt7d603B
Z81J79Tr++cf5W4wWkf1sJexUyt+NxorHU/rYaQGyTr+BdkkC1NRwEDPYJq/PDhU
mmx3Jdv5vZCMaAUXHnTYc4xXlDYQJ51S479ptSkKTn587ZXMQKcIptlHBvrdER1Y
TigahDzGcrivWqScvB167C9AkYSD5rR+v/YdvNlrOHVBPACJiz+mbkemIz5zxslD
W2LdPeiKjrcbyEyBrET4ik/A/AzdpzawIuBxwGN8vYkjWGTwEk1kw19IWhc9gRDD
R79oTmjFQqHsOqAXm0nmLiN3iJJ7iWcHqKQG68jpO8ButanCrbI6cFrQUNednZR4
YZapWtlzW6OnHZUCYSgLM50I4O1muy8AT4qwCPKEu1OpHPXupicgA490venx2/3k
FApzGiC11S5hy4zr71ZMYF3JmWbprp8VcK3LQG9xuqcMdgkxCI3BQPeyF8qRV9EW
UdW/FOpJjuXksBMyX085cbX0lEoFordOdwKA6LLLZWOL9aKvPivfpsAtXIiLis7U
7Cvkwt/iatEnMW/qpGhwuXQK4iG4CGMR9Nqz7sqtuwa1x+zCpBm201CoqoMwL1+u
z8tc7+0UB0MujQQGZJVqz8b0n9mUAX8cKpXbpsXKNRam/FeN50WAbCdKpfDcNnhB
uqGqTM7+HVB6XfKDd6NzmXa8WtGbbGNW/tX23Ce9PeE8KYM+DS/czptjQXuskrmj
97obqxAxkvdt7xSPH3jfJhxu66y5W1U8AYhaNcN3yDR9VRGWyR7/NswSD6yBTeeK
qOEjZcmijF82uod5QLJM48L7d7DQ5GGI7XLeRQPjiddRGdlSQ7/d7AX91Bo89taH
p3IaXEgRGR9m8Mt3JDCO3+2hREmDT6PanqsQLyjCvZ6K417WE3MBRA0quOcKbsx7
bDiAWkxbUuJL9MuXlS0/qfdp+9rU3AYia7Qyku2WIrB+2MI6PaHWTXPUJe4xNl5Q
5XX/sN3JI6wJeXIH4mTqh06KoLOLu5jo173ZCX+naRMZIv2yoxZ0KgI829P7H5xW
Ji/gbakDRHkWhVn4NUVx96srplAt/czZ59pT8kwHKKtTBFjzKE2PVUfckFdMfFgo
7yTDgdK1+mbFrxv2HHURE3BGVI6cbpTi0HV6qhaYACoKNAUfxA0by3b0zASWOhtc
TDKYh6MPxPvluElnnVd66Lp17vdzj2SiOmo8/a0ykaqIry82NC/esIOL6aIcGBV9
LGj+G7DFowr+BlOH5cUSWDqTUgKHsqZUvCqV8fk3W7SbyPT5fy8MfloqSpqA/61r
Dk1dwFZX9nge7Zu6plW26aKDYHeb4YR3NFjjGUY3uz2+SGAuiQ/PfKwvEDaX6XsB
JMgIuSW9zzaFrB8YMym39mspoCCvvJmpwUMhsU4p2rT+dF7W1axbFbEOCblk2sDf
2S4U8WQO/11EVJpc3vMqSZPsV3a4J54m4LUc8q5XJwAkwV6o1wMeIRrZJYGlOFtN
vK5skkSAbalZc9UIgW9psPp6NUL6iDXB9KChn/oEDqvUVVQ9gAT863fL99J7WFjf
74XkbLp3pBJzpZJwmAx1aAFlxDgpwnKPSQmgb6lqoVgIkryUqPWZ2FKPUrx/2X7+
NWHfoRhr/aKaKuZWGST5x+Y1+Ot47jiae9OhXN643NhNzHAWPmLdkudUs6e8Ym+6
FDq68xFfQYEMe62mVNisB0JlcySJC8Idbn2okgbLbbVTdjy4y7RkelQev3nN5m++
dmhgSZnthbkFfrRDwd+G1WQqzFLQO9d75717zp29KtVO+IN27aQrBdHqKhav1MqQ
zezlt2WxXCo6SJp4/6/yN2U2sBQt9ds3qhrKuIfOFDzQdaJbP1TmGYAtq3mtkv7E
ysGuSPHPFI+lv5GmoVD0BxISvAENd95GUpXAbk5HF5sm+KUpGHe2ClHWkzOJg8ZM
SUMUgxyAlbCyGT6fCg5dAqh7EEaD8/a5IhlmTOrzgIT8O0IELRWnRrZ5vjT7X8gG
Kmowq6RwsPUvFPQorbKawK2nO5qxtlVIPLuj4xMbR0F516tAsbeZi0qZgr+y6zrV
DKaMbmQ+UYP4JIP5mVM6kgdI9XOxx7G5XbUEMrpXqcBeIYqhNyLAfb5G5Dg/XTCe
/kwp8v5XGIJKALRjnKeHhGEKMjua1b6eCBhqMkkbm+bD8/+m+MM8S67MGP5wD8rV
HD5vDwQhz7J9zXkIxOo4lRZE7kNByBgw9mXihLGJMxGrXVqB4DlNRPX/UcARvd4u
+blcFESzlytP3JLrsraA5EjJnc8AmCI23910bpQjdQ9HrO6KDvO9gIs/8u5hZIpA
BQPawQ0cI5nJcimd0Y96dONAFFEXBYw52TXJDEP8WDlBlqq2YtYXcEHFBTI4tiGM
AGV/hjpfTKKvT1Mb+CJKOPDCGuufTFU9Tk1xKZa9pT0PprqrQ5Nz4Cv0eUSOOyfh
fDhAfhZuGuFylx8RBmWgOeQbxqpj8UrN0lTE0mrN+iVtxEg/O8ez4THX2OlXSLFE
J4UR3Oef26OQ8lunJnrW3GAUK7i2m5BLdWIVtMGGRO0+1TTYFQg0HN7rjHZBedlo
13WLKGDXgeUgMGkVW4Tu8rDdqzyxUAfkS+Siq+GAd2fosKaGWxcDeB6GjPlzRC/l
QNkHexF7ijOJ/IIMrurDOP/IfdMJTwlyu5jQVEESVKWtvAZQIF1C99/zTHfCfKP5
t4wyTJkYTjlB984t9vZ7qjT3QiOEJkVVtWWLQ2jpXChV9GTIU5wmYp0wxvOIRGSR
g3yTnQMtCExkQfOEzfLvY3l+kCztFczVwqIG8WI6G+DBrDkFiWFxT9+2SENuANrx
7IZ5wcUI2FFkKaRIiC8lQr33pTBi24iOXcjTr8VYfCsVaTHByOwKmkqHrN312wbj
lp14R3eQNplWJwfES9JAhfTxKElzDKZXxk3G+AVtx0wyce20TNxcThmXI1t5LNca
Mxky4CyDYlBiR7JMFWmG2mmf7t3CYmOLCWfPDZKEUC1JIfY+Hzx+2TQhU9K/KluM
Zr9QwyZsMJ5MNyxK9VmUq16wm/JmcWV+zfhCqrnBAUJqd2qajTtc5XYLLmYwL9wi
gM2h1SGmYqn2wsrZWQ48P6R1e5xiFRidpzpXUO6LCB4toiTFwRiSzzphGrQiq/nK
CxGkYYuA5pbmhl+WpsJ0mte07lPYcq4Z+AVcmbRfUoAr+7ckX0g2aZ/9FWplXqYz
jzuC3sHbbiNB2V+UbO1Iclt4Y0+yspI+jPOYiP+uO/I0Dkkmv/wYrtv+CPOh4KT0
9zmiynSpF+7/yZUV3GLQBDUzR4vZpXXZOoTSxopdNq6yxu5VGXkBnH1pQ+bJiWRW
EUM6wOGAblnXtb9HFRpQWjqvyo/iyLe4/JQxn40pCga58mj5WtfVb0JYH2xcL83u
jgav62wkDUCKj2FT7gYKTbJbwhkV5yEKyWcCzWLSETWOakJ1E/Ew1IclBeCFur3z
BKTeX1c+ItIP1G2lVe6fLCuhLmwvbdsxw6hfUycri/7DyW0TOBEHzAMmJffUQtPl
7gwK4XOOfuvTGaIvEwrfKuwClzPug9V1VGqeeiaof2w0KNjDinqXDanPGQCNLkKy
Fhv4EUlOcts8JKxIoh2e9vvyBTMdKcLhM005VjFOE9jsl9pL7MNiza9kpuwQf0Qg
NZyxNd/C8VJfkg6xcYiuEVOIYu9Ocjqz9eksHG168ddiQzvcjn8w2v//lIGVaa4t
kTBZpnDNTloZzij8Dv15vMr0Rs/pOQEaxxXZYH3fYJrevoKOgJIwzdyMpNs1Rhj3
BMmEH2mBfIvpKUBsG3DgB3xPdk9uPOeHYhNbLqKy2zzc3CcnnRbnWNKZm8ZgWxk1
Adh/ydlhsguxPfTk6KoZuFZ5WJYUgOa8mHvGc478mlOxJJmFvSDrbjJ0fdAbcdrh
6rT1r25sic2KFzn0K6JSVHihaZbC58HTB6f++TQ+j5z97C6sj2c2D0O2Pa+nE6rA
SiG1/xFrXNqN/YZheb2grv3dSUN73KA2MkTAhG17CBkO99r5DXzcBq5LoH/pjRIO
QQgPi1QX2vNvDdE2iumjD5yMmE9mA1bheWRyW+DJ6VBotOsYW5InYBYMLvMdKLfE
yrV5DommD97dP5v6ZrQEv+WB+YzGD8VGKG/g71qiU75IgUq1Lio94H8iMIlvOTZ2
DvOqGl7RNuX4ejLZpSNJMxgRBLIfDMVeqD6FYnHM3NOPu8U9vp3Y6v98GC14LExw
J/THshtyyfhxQApe9xahKgW2sw57Lhmwtx+82PsWlGLFMWBDwHOgNzkfoTeuJ4wy
3XGyucZ/XSdWShWlp48rwK6XXalKmx0swGCiZ36DOAd90rrE5mKktJtQtaNe6Nsx
1Cl/VtZ0k0ib45Y0UwlbvjnoWhOdNzomJZl+hGXeai3gtfnKxbkKGPbVNcVxb/OY
NguBfa6ZW2S6q5O8ahfCWYZKXMBUhAJsR1V2KKanM6APpiTPLU1hBVKuadQkzs4n
KCnEAtQLPBQgpXKddJgkJJf+B/SQR4p+cwfJv8Ci730lRLbZr8yN+a/ZTzPUay8e
f2PAdnW1bSBFdjVTaZEZVviCTWgFwHXG6NDxNE/orAG5MJ6DqLJzNvLLLRtjToN8
QhWcAdl9DWhx2hRnXX1+nZTeET59rKlwzMKww+K80qISjWuUgvCFhWhpF6TP5ZHJ
PDLWfZ57UBHuLGxK0LqEZWUzncHY9vjD87ll/RpkhV2+I+3lEITIWRl81e1zV2TI
6PIsjk5hn9nnFuec61gTpSnx/xcSmVSd1AuRewSBzrS3aRKeQRWwMiZqeTLniX+Y
Mcr7r2wchi12fy/cj9WrdO3tkEBamgEMIrj0cIG4QOOcZzBBsUH8Tp4a5C7Q2ROR
0jipCMaPGGlzLXdKGFN9LtbsdKqQLc5bmLkr/upVfbfx2x2WtZkoEu7e9e/L3W+J
mU9ajjT+sC0McakdbaHtZCx9vQNz2wh7sqna6wotMr3AfWLwgU204b1FNO2SptX0
xbxOC6ZjGz+3TB8+qYXorQXAs4I+BjlcqAeNIpl9fi6Lyw8ALT8RViP/cwQ4iEwN
R/LSKu+0wtG7AHu/QRqOisQBuXbqxOrdYlc3XF64zvCya/AfrqG1Z2kdJhDYe+mC
Ac7qNcP1R+3c2lvvrnD38VvkxptsifPGnEzw33AmgpLToHQAVxh6s5DFl5D2rfCw
kd2+jSMnf2sASW15CxoF52hI7Px+a+CsdQK7Urv1WkwowJGaYCGRNsPwtW9tFa12
OqnQo1AyFhZo44fM7CMubA984X29g75DxY7iAJaxvaUa5mLNAA3zgdcuyqJ9vKsw
JgFpTuJm8FE7KRnKyCNRk0qD4da374j/CM0m7wrgFe9F+2TUMbfuNG+7dPx1IGU+
Fn9x2BgB8gENHjVJFtb0rhrFyfuX4v45csoTsGEaQaNNXNvQlkAIlvvWAJeQ6UZF
l2H3ZqdZJ3A3wjaG6q4CDPZm7xyGBdvnLqPXzB4VzTtVRlzPvenQ9NCfEEZpUKN2
GqM7E+ShhBJ6ZwSBnxJ4/QTOfjUR5DiZK0V6daz0u78nuYvWY6hiV/bFW3hkzi1V
J/DYrA3jYdOWSRU1Teo00dHkVljFQRt+SUwXE4S7xAS7xwqpwV8nUme60NpHFo7N
tTw1f8gJLQwVzktojtJUq2lJts8xx8sTJmxbqnZN/j92+Dxih/lHWr4lYrjpt4r4
VezqsQMiID2wMXtGNKWt4LChFAiaD2l0JZ2pFUYrqM6fcyYAjFsISIG2osETXMQU
59llXoEnGJAYNSyzC8PLgVIftGMvDD+jsYPedmvaJw98WQEdjvvCasCqBKa7HO1C
F4NFAPem89en8excre4cuBacI3NY5R1fJHrSB7wL4IFlzXDRezQwf6CCUWu/Z+xE
kinN+i13EOMWXTGjlyznCr5dz6zWMXwE+sr4QS+LdiqCelXk5Hv+0mJv4/J+ii+/
8972B9DIdZ1ZPqWzX5FB8frKVt0AMfotbPZEo2eJwnYIwPOGiVRgWmjjXTeujROI
86Q7Wj6TxpgNdO4Hb8prS5a+mKP5n8QUsgQ5AiaBG4dA6odn3PLI2JoE8AcnWTLU
9sPGzfqv+f2Aigjj3HZkmDUrZJfYP4injHmziZB9bqjKep/cAzPhlKgmB4XlbkQ/
zsByw0HsdDdYrezJQaTSZSJfW980/zUdLpQd1881zpSJQvuClRC/jGeSHvaFTi9w
x7y7+yRGiWjs6eYUGP9PoqJnj357vAfW769ZJrXIvH5j0sw8iQaducQ1NFM1XL/z
NHCV2d6+hxvx4e2kSW2RBOxs+4SDvk3P6FHwR7UGWhuQ+5LaXDMXHhhsfM8BLyI9
trb1z7fErg5P/Dm37BAUq6YXrIJyEBLGFpN3zBNdNexeiP6CMYfv3oHho+IyFtib
+4BdaY7TBJHhmSo5OYqmnyyoO0OP+JzRWGZDktlScR4SUVlsjGGzPCRQPSTK7k4F
wZWElMYq8fBD8BSsC60vOqLphIx+2OUGc6lKoHXfwM0QFSZdrwY/OX9xcN/ZYCRz
8G155P8y+7Y4BlBT4OXiIVenDwjHVEekOoNl8zW0TUQUNWa4ba5vqYY91d17R74V
rX2i99xAOaj5iHtJFr/bTNZ1A/8QtW0DTCyOZA8uoaeHmyY+ytKzcd6sMf3dlHPP
CMjO7BYVWCkP5yuU87wBS4SFWz3DMDyxlV4G2BcEuPiSE2JwVNbLiyU33azfEhll
sLzuqUyaEvUfofbp+/0R3SsTAMMDA5GV3/lPQInHlrRu9KC9s4PFiy2kvOVaXGl9
L6GeKOoBQGh6EUrCoi01hJENeGLuATLTfC8H2sDAytWVJ/QHQVBF6F0DjI3P9V06
OBdMBtcDONSsy2dUAvIu5MWZJpkluiHx3PUkxixf7UHl8/NpUSOTXa6GpSwhRKgC
x7N3+qTv1pIPJeMWQp/3/zVPtekC9sIp+EcyYP4mdllpIfpOMHMT8oBz0J0yNfin
CjkH8yfw2MxO2hLc6ATlKTGo2mOd/6mhjzQtyrXirFGy3iUnq2A8JbHIZf0FSevm
ieLKxkUdWYd4jQGW1tkJbXCUOMkUzDaxH91mISHyNaQr1/u5P35KJMETHn1VE0/p
q2zx2X0Mc41IfVKXFpdqb41ZSoO0wB3sWlPOD9f+vbb8Uz/zXcmHvSf6dpC8+8Y1
aJq5lNvb5/KdtSMCsxgMADsnooIE+N1QPHSVd5VAETzvFcr3ynPGEjI9DUC8J9ej
2hNnyzCR7fgnuZ0QHjQ1/s0/+NgN4NQkH4i2ejVn87GPIbeS8j+zesuEp0fijbM8
eH7YHGaiU4Meh5241ZsNs9PbhqYGYtQ89+L1eH16aK6vGHgzplHGNpDd3LkS1KdF
GmeWvzdwIGnDXcyY4zsE2uzSVDRdrWvhOjCf/4PiqIOmvmQ2rSa7QBK7xh11+AcC
6lTdrk9egDc+D27Tf0Fb+etxtfnmgk/p275UzlVIdWrdP/OEr5ynfiT5w8UVf+re
L66Mj/BBC2iYmquB3bfoM4Yw+CltMybAVdmKVcIU7Dl9qZ2aam+rASoWJM5yoKx9
8UZd6US9cFyjI2IBjBI5J9TvAcmR/Sld9/Fh8YUe/3GPbi4wl8P45d4FUlCvO8+W
FOBIeDv+oi2UeVRjSwoUF3DkgyqPCg6VXOe+vNTv1uTXuzElz/M3gzq2K+l+8ofF
iE2EuIqQmlErn+xkekdaPgj30G302MMZcT5TbziHBCa+KbMQX4j2kGntrXHdjhuu
HaEyKgIV8aOEzqt24pnWI+Df5y+GGOySkj//JBlK3JNNPJkMuhNH+sLAyCVRwG+N
i5NsdRwdyfz59pMG7TsxpUjz7KKMk6Fl9f2FoH/h5Im/sRlSkgyUO67poXyxCp7j
BCHlK6aTaGaquY04IlqOT1gViBA8AhHehIk8D9EVDfdBCb/te5+YC+hS9H+HEEMd
ShZyYRyTbo2eFseAWBaE09dLzmblx7+DkZxt/G3lUxXsvRn47SXMqEoNNbfpTqYp
NmFRFr16twqZZP1S+KZAa95wbUNoabfGPQsmDc5Qz/mp2q19W/n7tvQ7j7n4ZucX
lh7rUexSnO2+RWI6BKGhNP6ca13qEtFoXEQvkIp1DozcidDo85pg1icalbBNCfVS
+YCxjwlZcPVOcu5H2NNr4EZbPqCseZntFSA+o4h3ZYOsDm0pflVXhO5DkOuzxc+y
WU40Mz7tBYP4fuog/cWop+qxhlyvIwB+mc9oTh4SQzyo9PJJvdmVWZkVxbp9NVJI
xv41sW6MVqE1hjKC20gGxIAyYFpS71NfRiU3RQODSKo8JbrmCgUZ971JcB+Wtu+6
PsHD4UbIx8FSfeg7c96EHESDBfW2ZiRWkl92/xHDZd1KQ25Jp0QShtLN5sKrDTvd
WtDByaiMrNHiSCPH7Kz+Zcl4o7zAy5EC4St8/Pk1VtSE+bpw0G6G2PPDSHjEEGZl
sJafsF0z2UuMexiXvwUpIWrALIGUgSV59s4cmg3K26rntEYqK8l/Q4krJlQFay+5
vKxra0JEVInXx9PVDEKR902UWKraxPGdlI4ctHf+1D/CicKEJDdnUwArxRJMEmdS
4/3D7+BV5Iq2m92c4bWFDIrdNYJ4zNsny67itJ5kIi3wS2ZxVKLwbwAuktLwX+lT
JTfaAx88ka200b6SElQaGgfy3U6SJlShzUqn+fuNco/LHkljgDIkWS6SpNYacdfl
XrxBQYWh3TXAaleaz68So6iEhR+uVijDWInXb/gCjvepbRyIxn1/odeUZdZJh4df
V9LMB83H2hMihOMGl39yf4BVXWOvd7diQ1Xyo6uwS8szyHCnXxUmEQIKbuFp4lC2
vIxvPHmXtOR77kdpwNDs2v39RsIdeNpVDy2mNSMQ7spqP90uhs3qtRr6lLNaFdGz
1wX8BfQUM8s2XatQB6CHQUNpko617nJFZL0XFEmw+m21dJ5jjixpyiix6xZduq8O
StCIjuNkguKUEYkK/4esvh8qoRhmNyP9JgjHCVjdBVYB2hzbDmn6Upg3YmCWSgi2
bx07Tdk4YNXgFiQNaeWKDDW8SVoNJ7gtiEOK7Ig4g0rk3uykHVxxs30wqs0qeI6p
kUFe0KWU5FZdC4WZMwk0Ns75/Tn9c1wKI3K26ufGaCILaK/sJ+Y51v9d0vUgTAVd
Qcwm/xnS2hq3qw9YmBp1TEELZrCOzWZ6OB0Isbe61g/jJ+C7AkiabuS2KnBZs2Z5
CWCK7JZ+ZxzTM3MuYtLgbB7D0wA/4vz+DFyM7c6w6+BuUGHehoUbjNV/EKeEaY7+
LYtbjpCY0bZcUfLyRCvn4x3ZFJ+KR2wEPxcYnuFlgK+ZZQwYbLEKLKs49EFBLiLM
Rrh1PSF82Jgcdw54jRQB2prjdLT6wmD/4xV8502Gj/lMG0/oj9gk9Zn5UzskBMKU
n1y+jundjNsryd9j9dWM3VsKgeFg2ifPB4RoilEd69piFEGfQXxZM3cvejsDXhkl
WT56lOiHN+ZZzYBJV364dJq85sysrfAYuEdHh+TXJrBJBH19MyKdRHqoICISsBIx
bSyTxn5I4guR4rB6slrqJBCQ2yWTZpIFHJDt35q0SuXRZdrYLqvf4NAxto7ho9li
OHa8Gp2PSxlK085XMmBz4jGaDUZmppFKtClTKWjBPMqtuT1pIttJIj/fZNbJif5E
JhqApsw+e9yTe1NpM38wAgNb5A3ZjN7AQSSBr0osORdGrIb1cvWaFURRAFdjijLk
I94XQOSRjCPTQqY7Sj3cvm6Rj4Ku7JOPWQz4zwscP7TX1BaWHscX9Nv72nrecBPu
7xPAjAbSDTeVpUmCWYGV/Q4RAuzWWllqw3bkDAY5SAdj5g5tHupzJY5uigTKWOxY
aPPNMJDUKhQPXXtrEO9BqwVZRX4Mq1tGKVV+t59EDavvmdK3tpCREBm7UTWJAVEd
0yeZXrtgVJyjGg3fgkGwWB54eP1pZzcwmXgnYehE2Zb+sPlk/h7wPKvcHQOrrj6d
zCLg9s242dkxeIuPb+XxFDjeGlBncp81v9PdXMAgu6y3igkWU1zsSbEzf1cYOkmz
W7DxyU4DLMMvNA/vdOOvQBKbNCd4v7Bz31003VC5H5NxCUVe26425yX241tjce4A
Q+dXs6+gZGRGh7aECHimiqGAUtD92UB2Q8j5gSpLV8QntTIjhuTsU/MzUWlNB8dt
MNLReEd4MVYPdWxJ5EDX9eiXdNohytegIl22uDlLCHFHXgWV72RCyHm1SAcewx95
FqXG61KNEPQXOyPDnwEvKOxdaeM/bSD8CAsqE3jAB7ZywoGY5265qNwhdAwk2+bO
XCoPoVG4r2IYDluhP73uhUyN29gD2PXSjVHEjy2bwjPFiOBH/KwD93Wx6iSEVJan
2MFm1v3yW8DKn9SJGSsL9rb6TxVncon/tseCblq+BTmTAjHaV7ZdespCn7jwUdse
ZY3nf6U9B4r2AVdMtf6fjz9tWDRMmMcAo6W/9p8+6Lipl6xwZOpl3+Vwy65ybnCX
o1rnF8+nv50AShLPEPsC+N0lis2LVPkYyxifpyz6w8Z/ZeVzaWdTf5vqg1tnSi1y
oPHMWnfKBK1hiQ7Bgj0HeSmcKKCxE3prDgMGICiur9zXl8u4y4SSiaeQll13lNxK
SAwSpWSZpN/d7d4P7/vfC72ph/Y4OGRzu8DQo2jNKfTakhhky3S4cb5ERy7KmLB2
MLoj9ksf7yqbCPahwf4MFkLDdDSH1qUNHXc2RxJl0zJMSoPLv8IkYeXlDR8nYLDF
P83u82LVLCMMRfWqO17aHNYWx1GA+1JjK66BsOMmhGhQcFonrw3fSFCFjwx9rlER
IpkxaJwTpoRKMlzUKrwWPHN45LhiCIDACWeUYgZJacEHps5M2gfBsYEqQQ4JVlG7
iprTzrLaIRdYVhR8Zqy2PZDVXrfrwFO8Sf94BZUTruZjsqB7yApurNWG69smPqBZ
1IJAew75YNbikiUKjvp9xoaeusCtcQ4Ut/QFY91PrUiTHsG0Fq+otghFn+pQ3Uyd
2XygCoxapa9CdlhkH2uo4+3A4kfD8JRiFKKiaYywLnC3pMJrf5exuNPKpf7nTnOE
I8oNWkRxr+b5AnrTeU+Bbj6qN1bIeI6j+n5Pg1xON+GYHykd92KWFH3h406jUGkV
17AC3GQVj+rRMX+yrDJC9W1PtGrfsD27aNZhEppUx/+F25dxnMsJgGTDIelpN4wc
RvT2AgXA86rEIgnm25s3+sE5uM3mKeepSOff/1QlgYl1N/OihhIdNUr8Wgy7PJ7d
yX1cE7HCZxFETkGKtkQDzc3+cQvwzTWQVopkhpDb4L5OaQvmMOzfs4KavpZ8P/Ai
2nHsoyK97owLqqyMn7WEOzqlhV55MkqNWQM5wFq4yL4XQ7UiTuuJFsMCA8V0HciI
XBzxKXMPSdska3UIEJe6E9v27Z5N35e2SPFMHW64IG17qIRF+/Abtu4KXAxcvHCX
FkM2hwujzWP79P+g8tngyZvIjgh1hy1mTlJ5xBPn5y44Ln5daXLCgjMc8SQT9cd8
Djk5MpZjchGlhiCp7jrVeJBpE/lBLKkwb21U9jcIbTWz1xm9hYxME5mfjSDU0c+Y
DwZ37iXpUhASp439waIl0/31h3Feggfphs7RvMvtgcWaO0YSuV4KT6ILGzzttypS
kd3mOT+NcXwsNQ9Qmjxz+0Jh8AhzJAPoBCNxDbKSUpIRinnYhpDqE2P8zNqtEuzO
EnjUJullB6qGEsHpdU0p4guXERUbZzPUgeffAGmXb8oYemInF5WJrN9AA2VSmIi4
MfdCbqAnemttR8K8tRFlneq4U419ZOnUzaAdGLYV5DD6Bi4xtLHG7f80H3i+fu7n
S2IWL3pmA0w8oM2/ooqbLrNDfolus7AEeL+pirGHZfL+vUlI5EG86O2ZBVp8v+xI
olvS//XXqMARpg24w5qRAT3JfuwXwlo1S2bPvQgiizyQBt8oMxMFUjR0n2NnenSG
NqYFSJt/4MsbcQDO8if/ilN+Sn9ZAzS1hR7odONWnMuug/di9Udo9yyaFW52kff2
rEDDvyWytnnJmNZlXW1mTRvsRC/mMyikIH8d1R8KXQcH3fdado1eyW6yRrahiDEM
+xPt9BHz3TCPoRwS9mL13UtUJcsqxFQq1epcQnBuPPYupzADa1Wr8VpA1joxyCjG
mJawlc38uJi1WdIeeM6TTO8OeqMKBdxWNdRAgCgbSsnpX8R7xwo2nF6nUxSs0e9A
wW+8v3AyIxFOSK/7nVbm7A3lu6406XIPfjinGxOEhlfom4R1Pj0NCzsHHdHkYEk8
MkjWfHAVCkQpofb055JntwMAWsv0Kda2Elsn1fNB3jDreB/KpQf6hOszxEWwyOYC
8m9bqhF6VaCd2bSFUMREG2Ww5ejZpu4feSU0N6mPclCYL0h8ZMr4fZy+y17Bhtgl
Se4atQ/8cSFl7KyKtaHH7NA59Uh7X8BvAV0gbNgAqtIqrxVFhaiXLnBLcEXwQ39/
ZnlbCDDXOOlDL3Ziz1y+J2MLJoDhR9m+mlC0BzGEMyJsJm4YYJBaoUdwWSU8WrF2
ZXvAxfFLWKZ9A79xZIFa8c2CUo03q/yz6yDh+uNvYEGoolCMwkG0XUw70dyKPSP5
qizvu3hFShWpD/WaPVaKO1l+SU0Qq5DgJJc7LurtChkoXHz4GLIkjE4UcRNSEh+X
Z0GrMaW6Jh9RPhajGQmz8nteiPVsOgzPAA0TkHJZgEpgprbW2vQ8NWvDtM1Pcb3Z
20b2jxn9XV6AhUtC1phjfAoA33E5cV2H7QuqVrjMgw7ZCjSv7B5HGZizkfTauFda
GngGomEsua6/rIhxwRop3UGI5N7Ft0KPw3TlrBJgoslGR1oaXZO0x0Ve4pXP8nI+
Pgkv2VIDyzUaRm3Of8OlNyQZafgIYEiXmezmchaLxI967g0THxb57z5TcrrHuByK
rqLzg34u8ydcJKBjkmOKIBNJ9pH0a4ORf/aaqfAYpZmLbatBfjem3Qx6e/CpoWFY
GI1IeA7MzL6tmKIWWP3xaacYUaJeX4oyiZH5+wZ0SCALJ9qbi0wjiPZzInEe2rqt
HfMb61eQmnYVjRImi2s5yTOTWwUbJK/YmpxfxWm3f3IIN28cRA3/ja5sr8dfADzK
ZPgJG4t/t/vUMuqJViKVuPhHEzGgMzF1o4L+97bHQC2ZbddYbGpPKRVOl/hcTSmB
RlUOwXwxl9JFdRFPnHV3yKsR/Qwp8EUVQYWVwKhiTGWBLEDiC4A7VurEBHmF2bic
TWc3DASPLhMjU7km26DMe6Flpb+3eiJ8l7NShcRQl7hN6mNve4ovZcfp4xrT4vyq
4hO6FaAxQHouG5+lwZ2AQSeGBj3BWanXCVvqXB+U9yS6K3NCZYLtEk3U9SVO7P9v
vo8p70mbXUKDU8qHHHvkYoiTa/wtMlGCiigC2vl4TPFi5cz7lENbyUM1w/vIrCjV
Ar5KJq/l0sToBv5kPcrpGZ1+gppPoUqzblYPTqg07Dvy1+lTlBQjfGaMKblOVitW
p0aNgM8CR+5+rSpfa7nQ06PzF0ajL4aHlyOnbSaeuCPEEWc/sTx38OkFhITlDCnS
HrMjEGnx7azuXizUSlLUZ6WV/lXN9pHmDB0SUPLMg9Q6iBa7yCm7cniGwBURMlpn
w78QKudlEbaJyj2+DegARoICXYwl1XmP1Q0O5POFtNr+LMmZDuCGX3hTx/0OEIZ/
WAhJBwlTFGPfnQKer3d4MUyK6uP/SY3+VoM6LXwYSh/Oj8ubTkuNqDs89Ix5aDK+
/wV/D3zcsoLPzDx3gbRCtSoXt7I6f32tEd6E2w3bh4D/lWOrJuETVq1hd/485g+v
VCQrpxRiT0OEgwtK9DKU0gq07zGoymvamGeY0VtAnq9saZt1BD/JIQqXC42haAMW
KI0gv/WucKPRd/dA3F7TNo4ljx5qsNoLCXjLGNKZ1fJqQWsYs4x7CFk6EpgTRhud
N9vRmk1p03Ht7p2XUakGST4s1DvsYVODOngCgeBUtZgd3dzq7FeDxmlQFqZTyCps
a+xm3pFWcXlpsTYlV7Yw8dwZ5cFcVBktFP2sJxkcbdWyRWLTKpbIJNtzSp737NLS
mFzFHHxZWHQlDwxgNUhdGMpVsk9fpqyZ0vw1+p0MH+QHwbi4xcoCMnzsAf45ZoM4
cJZjrCaPRHMfbkjU1Evr3fMzH+5KR0SBBHkNM8pe5ruBgiQDoRKhUDygV2lBXOQ4
GUuCFQLe8UMqbosIcPffElYLps55y/qohMWybekmIbwC/abxgPsYZj20z0prBp5g
bwlH0FVD/qHV2HOUQA0pvyvE4cpGs9+LMwAA0Mjc6S/rZv1f6Z/7AdbYLkYsrZKy
11ZGIbQhUCEfmHYkjiwcZjfNYDjMZJHVgQYIqhpPlxdRYTADTvZh61XzW87kw4Up
QfAcEmOJv5TBoNKQ6Zp5chdudMovhl/zegwIWoQaaVQftdQLNgmcIEV8M62O1S2D
Nk3Gb6RqafIeEitKXes5kA9rJoqfFLe0zUlByaO8qJc6U/5UtqBtgVC14X6vv+sV
qg4jhgcGHIZy6JTwpjtodDE70SO6XGbME7Taa/leWA/+bZWPvkshDNoGxwSh1uyG
T5e53yKewdyVkGhFYRAWvl841UeW/AykkzhGT4oVXGlxjjaXtNAwzx5rs593mEEk
qVb29xeIe4gdVCH/ozWotYeBjPp2t3IiXv+nyLI7NIWeyRWexVYcKDVd236AKR3p
yhBO02bR6kMdmaX+C413YIvRdVr0km6kh3PiGwSEsRNXVeamzoAk1xHefeVcp7GP
fZngwRaJrLtKibcIaPWHPa+4gsg0UHBLLykP6SSl0nMQfJ6RBRg0BM7PB94aYg9Q
4cp4sZyisGE9i44I4PdqH6ACJsFUqia92flsnezNYcH0Z3RIAyGbse6xpu/3dFLv
xWnJotXk+5SjxLAq39Oxb2OYuuN9feNw+gjsCWPYSuHnQUJcynkNRcd13UmPAbTk
9QWpV0rr1HbtXsAnDsW3jGkxeBtokBV2JCCZ53IVJvT1tsSpC5562JvpUp3+B3Ot
gBOq59SFxmOGO9diIkABHLHH55PbVA/Ahph9rijZpJ2MUDbFB25dtJ/zym6M7IUg
58/DzZSXDPMiJcEmPXgRwoPEoWsOP1Yi2MmDJIFGrzfpdI6aO2TILPha/Z6nZ1c6
4raQZTDuPJBPzgYitg5tsCAimbV8iww9ofFh+mIlWqUNxy/coML+MxAiq9VdoITt
PhJrquNQp/bpl2UecFn9ocq4dz0+Sh9O+qga15K5GcpYaUWYxQY0xQgJB2k+x1Ti
C2GlIeb9VQWJGQ8/trAgHolHy9ujTatU6T9XoEDXzAFpdjS3KZf1YAvp375Nd4ni
dSY4ayxKVIWC5C1TKxug5Wl4rDv+oSwGEimDICCBysnOfXCNqnx7nj/1mJRraWc7
4i28KK21uB5CY39UyQEaPcgymAkYxlqv8EhNEnO2Pgt+T37eKeYi2BZmoWiwMqyk
aTSz40H52YyLVAkg2tjxSa2Ih3nhG1W297k3nxV1UYPcOLWmj6JqkvR2o/mvRsan
LrkhIP2l4h021tMNilvQATCOys9L9Dgp8fcY1opiF3+vBRv4CN96d1iFmLzj9up6
QQc7pApICP368CDWwGSQJgS7A38CYQ9iLyDUsLClZCnTzvNRHDpEVd2IL5y+7v/W
/JonvO3SH8G1NEkCr8XoKmcX7OlUVww8zva9n0uQNaMcPxdnAD2LZMwadlwBS6sZ
X4rJbecwiUUEZQ17JJHyVTXasAs822ZrCXelh2mmGQkr64OZrTnJ7GV8CTdaQBcp
PiPAhmN5LaRAOBoakwNzOqcOLCVcRqz2AY7afYf1SsIAQ+SXskjK9X88l+GQFClR
fCiRf60N7v71DFyuvk6JjdJnwfsJMd+gLo5rFs1BMGjVfCTrch17B3NMyZZ/mh/p
AXL89ZdAo1USFfridAdPji7TxtPxwY6fZeGjy+i4TNuWDHM4ziZ2xN1xYykVHOl+
/TKpjnIBiVnFJeJPQlt49TjnmS4/E96a3Dfbd8V7bik7EtBApyK9wKImW3f2rXL9
Mh8orbrvlMdWctb02Qnv3fLaZzHmpCr4zh/yHBEPIvXdyKAVq98cS5w2izVpeiej
K3AJNVCapqAeOkiaYd9FlNVKZJC68XZMm8FqN51/2QG/BcGNgnt3IaTdnvjIe4Z2
UB+awenvGkcDm4lc6ceCYqqEWDY0OUF16sSL56oIx1XbpZL7dkCJpF51oSKcPMkY
xzwjf9Gs7pZjEWtJOp+mgwSBq+a/G244RoGu60h87+jHdHCSINlkjI6+y5JiEkae
wQNJOrg4KiUNx0m6sXwrBcS1HHFXm33I+/O9x+87Ly+VRheL9xiDbhw0K9ztVcou
EJQuhJ+c3rpD45GZhAFYExSSQvcBVQuRPy9R38DhqMptUjWqFuYIqEubWgs7FTM1
A/QGBFiBbIq1vdQuWdXW8rH6fyWgq6IjxDVdg8B7mu1oD5NIXoa/sKt/0hOsklrp
2Yk2Y5YwaS3K17yvbETbOSSpIvKW0/fntU9HvGVFFQ3saZs1ZXsunUH0GVM001vx
twN6qyZw0m4k1UsZOxPLcLZfBr4k1m7TGPc3fiWdwaFXxM8vqQjMhHzm2ZVTwefS
dE++uICJJp+CZU3Z6FpjUPFtSE74vDyqh36siVLsojBvJlYak5ZcAbxpw/46V0AW
wov43T/Yr7afU4/naLUDsfV5Mf4WX5EOe1fKnY3lyk8sZPI0+QO3xTF1fq9GdYjM
u2Ujsk2BE8oWPeRHovb0f4G55YabBjTq9UbTkf9jGVeNNiG5+SllJXKxFvOWf22c
hwYV6IkD/ZYKysT6MJidiAXqj/iJ5R9tJjZuUR20p/oT9q5LtcjMpbL158qV2KzI
BptAKY1g5SUGh3F6pHh3LY0BOb81v8zXqWs8pDLFfzqvdFWiMbEC/y90yur8Nj32
D9omjpXWhrjVfKFJOeDpGI9xOZxIrbR1zaKMSOzRkTwolOYINZUqEIwCEQFc1VmZ
A637BO8vdhl/E8NzX6sEXasUwdVPbnFvWLEdFgzK7SEcGzKXndb23GeMss84jv22
kcE8oD+zk9HrnKN0JoTfz9ePls7Ki71Cax/u/xDYWhZPxBjXBrj24QiIBqIPclKT
7q/+l4g+bl2mNBv+0L0wnhRscU+/xHXyP9MQz7LOFvwK5QuDK5i9baavujavSFma
LyFhIouig7i4dQh6Xx9dI24ky26zkMfXTj9uoDdn/c3NHrZb3ykkOtMada81F4uc
e9cAK8F2m5W1LSmU0XzYxmzkQQLfgWlW7LdLsGH8SpbWUXf5fxsYVVivCFp00XCd
U72q+0c6IgNr70Z2R4LjN+ZxY7Lao5WkPdMzMXKOW4NfyIzEmnjq4sNGrUFsbioV
CcnjISpNTgjvo8TgoYGTG8cuMCwOZItLy7d986I6t1wWVklIeU++OGMpMhk4zGEs
q+AjiTpKiC4ezq39eCDnxRtbMNsPdsIt0UfQVYse4nUKGvz5KogKZKQvHWBITcBH
5pD8xf+Y+SpfdHDEOV+rhdc7HkwxQJXCGgTyyQi40x3r4t3G00SvBdjKQTse6hsy
KO3y4HZAColex+pJIk+t5kZge1xrEK8PbLj9YApFm2owrx9mNPEaxQJ6QPmJpgEQ
7Fwh+dZCoIhnr/m0jOa4PjEn1Y9pj1aaGOCR8CehoYSwffEv7NyhVX3JfoSd9xIp
wmxSY/HcSX2gAYfM8FDrvHmqvylw0Biyb9pumhHwf4irknzlt5w5U4D+Q31qm5Xv
wx62o/a7yUeSjT+plh0qC3TkurNKvoBpHitlKcjsuj6Zx6bd98m62CmpXlWPQULr
K7GPYIVFQVuPCLYDdjV7E4ydu95ZxD4uVqmjwSVXJxWfxGwd1wp3qtxBDcCCbl1P
VeVqlZ6cTfelJPHqCIm/S1WVuJJ584QCgGtdBmOm78PVAJQNvx7V9HvhudQo8DLL
lskuvpRSJ+dxmfMqI1sAlgEGS4V6lUO+YX2/sBwjXsDeJxxb6HudDBJQ9R03V0DM
hcg4sJru7TY4+WsDXdvnAuvamMcwUSVtDMEf96hOLzvsxcvbdG3esfn4chCqP6e5
bDykD1fWbptMH+gMd3G9s2ph/4ftxdyKQlc36JnzbE5uoErmb/h0DT6HP7IQMLnH
F4RRUVp1rMqK+d8F8jU5HmiNHanARQW8MKn8hzFRqWcAh1akFPbSxW0LoDpXxHn9
NY+mc9V9qqxQryQPCzlFpkBrukuSLPtbMBG27GmWEkcn3X4KTbo01X7vBYijthCY
tUQeIOyCR5p+/ty13hUXqy2YttXrUT1nMbTouvvGyq3kj4MWorNAt2n3XYODeFCF
BosTewV9ULIETAvFyrDSm499eopaNRHRr2s3YuHQJfdWH1NXWWEnA2dQ/OY+nkhp
+9m9TJmDzbgHQTSV4Dj62nV5yMn6TTjlVe/owvdwt+6vhM3R5mkYCBx4CfuBy7sy
xbz3r1jublQ+sq47AWnjbODA+Qo/SwlE1gBUcjPoKa2y0bLO+osdJkBoyNtd//ez
EVropyZGgj3XWQL4FdaA9bz3D4dSbikSD0jmzstXHn2n3I+d38Uatp3hcxstmhhO
uPURqzR6q+t8CVu1xJDtWOmpgaJS5C7h5ms3E4dexl2z+TDLTcCpVIMiC2ueJ/t0
Ky5Se5fc4GAfGcXfsfRJSn5gwrNaD5nxxcrIk82+2COD7AO4cD4OGNIQ9Ir5kXzY
PZqALtyOZtUjG8iyJJs4IpC6UZGSrfohQ1vzQnA7lSfAUkcE/WtrI8RBiVbq2kej
ZdgSWRLpAk4CjZB6rxqIS0v2W6biRRnNE5eEP72KCbJ0CcCQIkKWLeD5vHg4wNez
amv/jbMnctIBSck29nNBwzfsZJqFq3TOHBxQee3pyIYvqcHee9mVL8DwzH5AWklT
bi+97tWskEXzMwQJEJjm/eIRnLsvlDt9TLJI+xs6CyrlZlHGBhjAak4Sty9UnHu9
1bxg+a4peUuWyzOtWdFQGur3+v6MXQOdtYUQ6XdG8JULoE29IgVX8eOhosAwYnSL
93qFRNEEF+eiwHQc71HtvAqpC2Q87mNJZD24DKW2/9GY4OjMVmMIGPi2hEc1+EAe
ECNuqbW1Tie34oUg3N0deJdjl9NlcPIUN46gkweplsR/JvuVw+sVDL0vVruiHOXX
af1D1J3SCKDqCl0I9On1tAlPy8TzlSJXB2AW16852ziK6ijYPWedwqqDGG1GiegB
ymE7LJrrOYQl8V/nyDDJh61xkDqLHhVn+92TgX1t5G6oGqDlurZpUvyM/rD7D8qN
QdG8Hbt52ZQb4LJXkQjIW39KwlcqBcnfkGHXuJqvRiQpckViBM9fv16/OZJOHwTh
q0Q3vd0aO3uK6H9T/irWv3CP/Ctjd3+kTdajkInMlUR44Ptm/DiQ0sfU8DAQJrz6
+BC+Cz+4IvA7AH2VsP4B1Ine5iu3Yb+bQcbNPBvOgXuXxx9fgvxuYN0ie9zTmUOq
AGywgv/eRaxvyYQRxsdojrrjkj7STjqEEO98cLUVxpONtHWG4nNQc4R7ABd1bbVr
07jyL9B0emwAejO6Wvb04BZQ2jVl+BaYyo7A67uh1lKjdqO/NzO0N9+OI56/v7Dq
pW4GcC4yVv1EfBfsSbgGkeenv5JiZXZPtiq3UAknW0sJ0Bzn8Wz+g5kKt91N8emB
IIw0m4Zft/b/jFs2810nN51QZFXR0LEKDfsTvzABl9NnTbM4jJq4EATz6QBzYM8m
AmYt6Ba4ZmAeMkQOkP+cEfPhz7RVzAoxqKpGw8aziw1Z6Ym0TRZh0yZyiV2O+xGi
agYB8cXGUIYK9gohBFJOBKQwvsvjhJHup1mLwwhOkP+1WkAoqDZQGzj5n+5UW5l/
qvlUelDXQB+MfdTyVocwKrLmpno8v3BcNcaS47ARV8UZ8wEJdzAK+INmI9j9mqCO
+ROeRCtgyNOdGcru7gfRCa3Mg5mRPKAfdQED2kVosER+XeBK0xJ1TlUqM32UtLSJ
PGKXIraexgIJCnbpDT54dKhwOGpVFqQGym6GXy9w26cHyJtgiXxRdwisJIU+rEka
ILDfmsafG4AUK8ZDtQDe2Xgg8u5kbcsNB+G3ofL8och8dhHRc4GMU3ISTZ0Cg/Es
RomqDjOEKHMFzCyXhckxzKysI6wyI3NVOdOr12+328t626HAHUqSPEnHnjqtidkc
hjr8HT9OvWtkwCSZ6GbE73wU8xt74cidcD5Uy4WIaFL4p2AcE5cf5ggwrD5AFRNo
Z/Fu3pqrbv5SA0T3d49sRjQgwDWa61J77SruMQLgvYqSIPu86csUmFJsI3lfy5Kl
lmSSXGAcZosyNc84n8UyhmMSOKK3vddwEI2vEHu3JdgIkQ2ptp7+5Rjb2KITjmXE
N+EFYK0t1TIgm3Lqf0rzuQp0L6UPpfGOia5NqHnzhMId21L0PBYw0eoUCmS7tLU6
wGYRZTg5A4HQUVdXsHh28mzoSdOHUb4YTe0UTua+KbRjMvm22WeaVjaHHU4HV5Gn
F2a73TVQuHm5uzMaLtzHFQvfKumBxNM9sZy0tovvMISgT02+67YS3Y/LjqKaDDzt
st2xW4e+zwm5uVXDdBZXTCMmcDC7wadCW27VEVPpX0t3AEzJyjFL0o4V3kricLIE
F2NIHPgZTFIX8As6pZNMv3FSFqFD+Fdyez/kEYjUzHGNXUUwkrTnY5htDnZM0ZZd
IcPsjDP/Llw527U9boJAvO4HE8+fl2YkX+nt8risuj2pj3fRqA4oM51a4cqywJN9
1U3bZ3Pdl0saGHWiU9qM7dTXCS9W1RK4mPpjnOr3NBXiCrV2pl9RwMqY0WuOt1aZ
PdA6qLxnXf16IDePao+RsY/i8SwOFQYAj0h0Vvfsu5C++btXEfvSXwPRmZzb/RbG
RtSrNO7xwvdmFnvPKTMkSxCqvu0Wm26xX8yS2KjqB4A6ZM/wigtwz6k1gCj8g/0p
xS/jvk8XgSz3wafvIpvigHWhL/cgzOtgoqEQVrjNujB2pQ14QoJwc0dDzE1bzcdr
auYbaF412UUhOgMG279Lqmz6Ex/TXTM1h33PNehZGNMErm0Ov4ixMNHszffJCcJH
6KJKQ5OS3+s7EV7M4k0te6x21D8fnMI8NbBhZiDUUxfgS6fFkGgK+RM81UfDfmrV
fX5nnvKiSel9fIOBtEu+zlFZVLHyGif7g05K+qapZpcectEOiWwBO98PgtncAhYd
n4hohisRycAW5YLBwlYnsCYL53I9yxDEm3S3ApOk/jNeAnQPxcwMVr598tGGtZFw
Ix55Cv2mo+P/Rcm7qt0bMw3Y9ci+qqo0T7DiHIqXyJHkvRCi9us3tKerS44qHt+C
64EFTp9ei0VFYBuh0jFd6h53gq44QhLn710jxsAcar+0uo1Z8WcNsKB00MvwauZU
zXgGmJ05+e/3vm6QmmzCsOsGEFF6ALpbjaymqNjKSI9CDsx2Q0dQMNYHdmCU9Jof
xYJQA/Iso/V3s+Qks1x44fYxegWHpio5ZyzjHPFPRqKfTP4lplxT12GbfVJEaMRQ
85ErALvStUekQ8OUw46VqrSHPsaUUqXsI7V2vxn2kv9Lhoy0Sk8z03LPm7XuORwM
PgeuZLjItW713C5wpeMfzVtwt1sTnUvBh3Ntu2PG+KZkmLkvGT8u3IMNaY92ZbdY
YN67CtFDm/RvdXhBPpe9T9y2umSu7VKxo7OrUo2k4lBF9Ny2aSqzlOZVPboaz1wS
iWo1lewN2O/vsy+17tT3F+YL29w3YpNr0JzhRMP1YbCoIucX36luq/OrvZNPf7TZ
JuYHI788HFRpsniFxHLj1D5I8551lrWztamUga/MiPxQ/GKDIhs7HHZljhfWCMi5
hYvEhwFNP7pgwZGEPhpMOoc5Rr3L5gw0KaTiJPt8ZSyedWlQx0KVYZm7I0ZjZoT9
EGLICZV5Itam2fnfB3etdmFQRyIpJ5Vw7zZFkvpqom8GWiKYs2a/RlUqjcLOJdNn
QXV2sT1b3/0PMiiHQkr/Bm89ET9d6hVUYNTft0WEZEs2a8jb/aOCoOxPb2iG/fnY
iZjrV0p26WaiFwNlGXpd0LjGm2+EEf3oFRcSPRspJ/SXnUmEWO6o4RKZZnbwNSgy
8qxucVvspyUlHWEU5haOkAbE66jmfzGGccK47tvvbOw2mltWKex/jT/qqE6xPCAZ
l8YKtTXTWCRvFGO2i49+OJEpEYPEKXyu9rPZNddlFSKGMGbV0RmdJwjO5E62K1Yp
fi96i8c3kqvicriyZt37YSKlsenUKX0Vp6VqX43vl/SZ3fJL0rgV/qzyoY6yVjcw
ii4LKbZfENXBR9pICkYYbQ0uRfXPQl8JORH/MidqeZtphxjbxOSgiGCLfzY3bKCC
c+FUaQSwa537R/MIqxU/mFMt2Gr1rsPh92+pTPNqOx7tPiLOsvbwEkn9tA1ePNaO
IOf2nW6k0Y07PxXuzBeN24+ngcgG9mvyWlsuBL02Fn81is5Lx5noRNL26lKvf2hO
zYHH9iujQAfRx3MTHoHcrZxeKvP1mdfpEuENOHVvH+65UK4HTnmWfMCEeQFaRwkS
kze+vzcZbYV5PL7rkEkZjumtKjW5uVtrgaxjUfGSBqAGqPL9tteTi1szV2GbKRud
2KdsngPtGbFxJqrKOZhkjdgspk2VFXTkpIT0Hs+7U7NWsI4BrzxNdv+6UxvQWuMM
Fz1T2RMgfEcfCjTu4SgLJzMoiserENO2IDvsxIa/AJPjPtrSuYgc/MX54qm/HRqP
hv0VcpPK/umnrS6YqAHVe/OuvK7ypLbQOEazCmtWzp91/Lad3qHBk6WznntL2E/m
8Jy7aLHcE/g/rg9ybmTXn28kT9FnbYJKIIl2lIwW05VnKKeYt9Z5+OK0b+q7Cnvx
J3cVFasY46Oc3BrxCDd0dlDNFkD56QOtsp4yT2hAdfqDKDGjkT77MyQsRe+nvC3D
ATOrd8xrTen+Ivu8hP8ouNhMbMtS8M9wusv6du91ih5HD3stB5T57dLWZ4Hc8m8r
vZhdIjXdeQH4heWl2flPByRIXC0CjDeiWVpE2ubeSBCTAxO+1zykQyi4QU+om5Ie
Dk2Dej31WIzdnJFRC6Hz+zypqveXWaNZ5EsmdmS9L3yZWRyfhCIdovWv0PTmSD2x
TNZI7EOaeQbjbN1FQKvZe9VPwIzzZL+wmguMoaugczhWBB1dx02BgQnDxSYDp1YO
2cwTNrkfFp31836MhflCe8DaFi8eHfhufcLYV+LYS29QhjyisSzWzTmKAsfceDKy
qJCHcL0Mr8ZDchugxeSB1+wzpTc++35dxYr6NU+e/KPRwU1ZDMn3R6Opc9QmAf0g
I0dSegrB7ACtoCCUVpr500LvrCKVbJEoLbFRhwtzYHPYB4bxyM+NL72A4MmN40Ny
QwtDfmrD+t19CfPwqoSLCFKAYW3aGhzho467jJd/EH/7SkWVvOKNGtEoz0h6Q8Ec
IaLd6VSpOBEnlE7fM2Mn2OAVLS7GeMEOPvSPzbGgw7NjqhMMVZIaWazf6N6DilDg
quCz0lYAMdnahxO6waAZKkfXA5ymLKlrTouj6/ng2N3dyx09BA2f/2MIixUbiSO3
`protect end_protected