`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7184 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMWORzZC7bo0toZS2Zods6Xs
yljw+BvqICQb54hGe2JGpCy7VfzPucQWBxxbAs+GRahx4zSgSeugyTMUqyOg/zI/
n+aj8gBeA+kwbOZMEZUXB9Bbb2CBzrv/L66g4kq+VXJMVrfSIB+F5/Q7wgl4+a+S
Sns7SmGzTrM2yelmt27qUNqYMPRZcJGejNL0lhxYI4AOI5sWpFqJKr7JL4OwIg22
kzC/Pzg6KT0i10NXHZVBHeIzgB5PLelpZLuSLiz5lhlAO84Dn+an8RuUd4lFoKc2
uFehlGLdoji4Jrrr+B7UP0mBMzU5fnLWQSM/osEwounvnlxXgqBIqMhFRMOeSv51
pno0igDmElJgidcxbejuoLSgxEij7LfI6FgF1tcan2wQDKdj+B7KyyZj+Lqvl1TN
CGeEqQAKFXCHTn29LKY6nKUeXTDqrpN0JHXwfUWFy+dK+ZzsxvsLdAourURFnEJN
ZsZx+E83g6JkPyyDyZENcYyTjGPZWwyA9VZ0nsGxgdzbFMaWimtRLY12L904vyq9
V3D0D1oYS0CFcAUcpSkLEHOZLnoj8FihJx2+HJFRrxVhKe/bbhvezY3vAZNpe1qK
LnsIY4pgw1GZSR65fRke22HqjnE2FCAKMGcVYMIq7n7PtO7wR3iYRaQtpSBpW/Qy
A5n28dzM47/M3jM8DUIDil0BOcZfFD5N/szym76eyZBQUcV1riinxa3L6NdpQ/qV
LrmgG4eXDqbjN2CPv4o5Qvx1lqQTBBJ8c6+C8VeHTKuwUOcls2pd0HbmY+HF2byC
bvG+DGgfWMVlowT4u7B8dkzRoZnk1Zz4noaIlhDd3ZmIbfegozDE+AM7yZyRrCDB
rfOBa+LTZdcKuLeRJRtMoJw+js5yD35LVEzlJww1d+fidjy0c9lam7SL4Bxc/gCz
AdtPUcY7YbrbDCWXXWKLHtI2BWkjL3zW2XupqAdA4EZRhtLAMzv+Oqmvl9dO10Pr
Kqacn1fn9i7s8ZX/rrRG2U+JwVWjIv2clqz+bsU4Bt20/4ugH36QTpUQJkU0tEHr
2UVfEhhsKUDDqYFnBhRBt0GOMO93zqCeFTjcmDbsLHbt3DvL6TWu15NIdbr0/SBF
HCvswgxOzBvHJQG6BWnATgqBN9O3/uj7MU7FGrVTvndr9GUIBNkHoGNwf0oKGBN/
VOk570vywXx/460LhFxyka6mtmm8F0UX9wz4Sc9L0ZQa4srdxVoDsUq2NQof1IYg
tEaeBG+GBTxWRvvqlFVBI8xa+Y83TtkuTvRZYXsJJJu0B679HvLWl87Bv88A0tUX
ke5eNL7lV/R5AbqZ1W/fOkkOAqPH89vQAfGFY4tD3km7aaWzNaQG7w8xJosODj/C
ymxr+cPt7lWbpcKmAcBtehv4g0UtDsZlJfp9kfZhe27FOVs9VcCLQvP4KOtffu4j
x/80YjSaRADXtXd3SQsrYSaJ74tLVkkZNxm7IlF8j28EkajEJpAoQIcT8HTf8WsU
oyh8nNRIy76S76JGqPOMZnU8paBUYU19D13V5wM9HL8F0BR+5byHKJzLmsMvh5AC
0lSmY9esS4vg1Zj+Ln2y89m8QEnX1HNk3RK1SqDUu+MpjzS82jc3ZpPbmVi2Cap4
tQ5qCcwK03pPSV7/vrnS2WPujNvt22uhU28Awm/51bnC/YjEmDyM8X5E6eiRI/Ni
G5UPqGWHG0UDCUm9BWrkNTRWc2fFFFnUONRgnCprXrACW66tb+9VSP3OuqGiV/IS
eqhg2e6SAcUqSKtcP78aa4X63m23alkHD3lsw5fx0NW8IYwh4phuG+4XnLPPz1PV
3pPWpJubujavcxFa3glCyCCI5WMcahUZjdyw0TNFp0Qek4P8tdAf6wCdw6BPf05K
MebIfzjcrsM3nU/c78TIwEcNS93NvfSUzg15QL6cQuuKZVhJswoG4OyoAxf/MyJZ
sR/Q2X2kBYEpE2i463dxkcHSUWmI+aqIyVRY0ZYagBviwlUxfwwpyv3MFEZyCrv+
JdjLn97Y3n0esaE4RUiD2hDhj8uvUtEG6hD8N7OxcnHwsnZ+NALcFIKFYzJi3HUN
satZX40rdMKvC7L0l29+V47BHvmPIhlH5Z0oBxucxRgvFWyWgPWy0tCkVXOw11+g
JlEQS5v5Q5bThFedwhrw2h55M6U/2thK8tc3JvWGW8wghbehdbKYkvTYu5D3SxL3
IBFqD2rqcM9VsnlUgtmh14+5uU5EiIKNYghh5Vd2AbgvUarhXvAy0nEvbzcDuDRV
QfJyIygdQyBJVyTUpefSaWuouizeIQy9kmXLxkJ40uh87j6MHkWjZ8jw00kZk1t8
pJNHd4JoNlDjOlBVFyQ7N4iOuNRlEnwemFlpSTZtWhimvM87llj02Ya1Hd43Gnem
vPuEzcSVfiPkUOBD/QhcWj4mgsMPaMYIcO/4hSIs7bLpEPkFFRlC5v7ibLrU37mE
IMK2ZpPxkuAecwTPgD/UOvr18Te5VTqVV6mS4c+d5o0645uELH8C4kaV5LYWGJVr
xqfJMZK11N2qXOt+k+o+k62KxhS71EKY1dJts2LJbJHmXGMNxlMZjbG78yohujL3
Ku11Xzci4lDMkr1BvgIv3CyEQZnzYz60a9S0Zjl5vgyaWmZeciLTu0X1gvHWok2L
U2jS6pLuYxHoBQDDa8epffcCD8xf4iZIWpffYkRod79gMR+8ZJyVbkoZsNp2WVnG
bCsPk0Bg5yZFosWuZQgnKKsL6n4GlchNawboDh9nCTaabBa2Hb74rls8r42Xbhm+
aH/qftbcXmzGupxHoL+PTxKLanENgQOgtFbR2VNuB3dhEcoGdXMAILYNLxznjtUM
gpUZjLWy6zgcorctweYi8F/LKc1xSbJ4lD3/zrkbx+Vv2mlTf5lMkyVqYsSoXnJn
i/QpOdg+czjZsnZWazpMFoWDDh2OTQLl3EGAX9unD+AfYVwsY/cqXvEGNWKDmDbk
CgjHq1wjMqE5C0TENYUuXH6KPnBRDN6XuhgHdpczbb7tUzZsRMbJ3Ad8BoftPq/B
Hgt6Bdizp8wikVkA9JQgGk742DvLWc/1jWZaFyMK3RmipHpH78lW8S/4R89dC35A
ozxg7jwLgdMIfDocIU/LHX+UEd5mgjYC02VSp4NnxLnw/+mDI5UUldmUmocDOWrt
aTEWc9mi9/hzE1u9kXhVtvImVwYvJEjEAutcPNvesqwkwShtz0A09waJjqnxSqur
tt8S7tAMo7FGxdply4jk1HTgnnzk37rE9k0VuyyWMqSC157LbA8EJ1RFJ1IAtvjR
/mR5rx7EI25AavhmgDcTAmlKr4MI4LaniKKmAE8418AO2Qsgn1sTuHSkTjJL0p7d
TemysUrmmMbl6uPHooCdSL+TableleYGgGB5CKvYl452x5DQcO/e0mN4xNSuNQLU
cE3qf4P/pKrM68zv5qhwXTcm5gEBl58UqOXy0KtaDc5E00HFbwyovQ646DYKkAln
FK98r+MyAFJY1ZreMkl8xyBbtUSHPBu42jfn0gkeSbkUU2xz/oK0iP/5nptKjp4M
98b6qfHKW8YGgxI8hlpXVrqocFo1FUjwLx1R090M5n0Kv0+6KRaPnNcR0AIjoAVw
IY+iGnIs8/K7lMGky21XfneOUUCBI9IITu6DGCENha69n0Z6jY1k6B/N/wMvQeFR
c8BMXju/FLbndd5bLJHsDXeqimA0kRvQ4CZF6POTY4ank4IFubLB7f95jVJ1cogQ
i/cTks5LmKQVqJhRWkVaHhx0s55XjDPOyzaJJ9U9hvUzMCHL4af3/l0dNuMfnSdx
E0GO1qnTPXfQIfSipXryQ3pOfWzC3aB4We7wwegRyFhC5q17QH7eSSzs7bqv3PjG
KLTM40kXT9IWJTnSvZZM1QSYVuLKfJodS3zxevEOrRa3tKdw8l31aTCyKNGhTavm
6/bNDvYyE2mBaU7l9v9dDV5nuoDPNnAPCOcfK6WIJEYACL0TUAegX8y6jj2HmFlq
gwGnoIWLBh8KWtfaiIJzHYvzPOVozcSuwvE73vZ8pNyHTk37F6y0Q97s7cm6yJj7
p8y0AZdJjRA36j+1RuU8faChE9jiu6eou5voxLXFo4cmDzjyL7VCxSXpHyTvv7Pj
H+1lP93rmHQRSdTPFikDgugvzrhXxsrgHjfFHMRpHfPwfc1ZZTNm0DB/iALW8wpG
rUDSBZYtxdSxwHHuQoXBTCyfcLjmY66nwj/w4OCZfCSwy29ja3fYuLkQQ0iXnjHM
jqQ808Dlz6yQ/W/Prj/+zs5qNsoXw9I39wJ12zdnAk0jK7lEAv48av09LXKJuuH6
PjDf4VSjRLZga4olj2J6hx/f5Bo/geb1/4KHuzXwVznGx1qTSvBi98YJGYR2kC4p
DTWiExyn0Nplzf66DKrbjGvtcqZVCEqBDZ4PfSDfn3Zikvuz4sO51hbDxccFhqEH
QRe0Cud7qzTfHuYPG69py1JfguDhg7+s3v1yuKwC1imr1HIPhamFU+nw1J1cXYDX
7dRDTHwxo8ZzJqsVkybAq5oKRGKB2ky9qoLhWEwfPOK+utc4/tVRWcKs2+6mNf16
roG9uykA1QMzfMxFmQepE96US19CoiVBgh68H5dc7wQIlynyG1+o1HG78i041t4j
PafXVtrqnz7Nk9/5dXNWFKCP8zk7T0DMriRkx5bW5xJ19rS2eSZ9u7L+vBlS8/mI
B7Csy68D6DNdVG1Uw4GCypTYl53n1LZn3f34dgGqGW8PcQamBSuYoPEpEuhS6ob/
BGHdJ38rSCP1p5hd12rXiPfCxh2iNPzFKjWoI/xSTOMX7QnINuzUpF0QXcW52LEW
bZ87mQhm+Y/VhIfUlytVke1VFCOiEwscvrZ0QXBQ4q2vfp1U5SE7vpVdBPgqtVTy
hurQFIZVkKU/CmM0yj5md8dagfay972xOaRbIgE/HoQkGZe0stdfG2hyOrUyykdT
qr+rMuVVtZbIkxsKMfL33VjgzgdSt8Xaz5wRQQLRFpNF+8JAUSLTMDvnF2yl/rmt
u1tML59fjm2wCs8d8b/3G383l5yJt2POXd7YazgYDGdtb1Ndsr85YMewnyWI9FM2
DTQwP1OTsZ1oIZ0FzfoAe3/S9U9wTirS9tkJ1yY0AHl5TA8MUAvHHLsSCwuPvswJ
734vUAt3dy5qit/JDMMVR7MOkiBv9eTa6ABr2h7Wd3jMZTwx4eN2M1IbujswuMgV
Q50U430DBz29OtBkq2u5ZuwGGQ8rRQvW8ciSIwnZVPStWtvW53uVDu9sJvQZPT/B
wIi2qGPZPG6nFHTOSsZOLYytd/bsaGifhgwEdOlEqfXxEaWtc5ZEBaIqwcEqZIFS
J+ZIya9d1CcmyyDUVkptq+xBd/kB3bxugSYJfHGm0OoZJIvy1naJgI30mLnzf5r9
c+bSvYZtbbc9fpfx/peGdHt1Gam531rGYZT6ExNEzEBl9cy1O/NPs1Ld4EdbUfnW
TSDKrQuMsDu6fx6g+760uJaCEi6UhJHhQOIZh+GdikoYpcV7ygqzZWcOpIx1pT2r
cQP0DizUIZRa2HiU3W8vzbuHjLJ89lY2TtvE/zcef69mkEtamco7BbCL9KSuuIQX
uP6x7ddO4biLXRRYjofokPxYbqmkK0vVGtNuQNiBD1THJvsr2xFwsTeU4g6/5YB2
prAuhrcLEUVQ8ZOyusAZdL835kVcmuqE5T9Cxdd6Vk+Eu9EIHYWfbDiSnnrqenO6
ptjxOPItji9f/R2pFeyjjuejT7wli6U73EI7H1LgCwNT3iAf73OO94eOFPuM1WK+
Aj+k3F8B6tv104qGZw/Yx9jTPUSw25beov56Nu/qbWzbLrNrqwW2536nVzS9Ri1B
vqyBjgseHTVuE6s1oMkU/cOSF+RhnYShxSiycnyjTJuksPbjSmxT92rstphAN6Uw
az5+zgQejC/2GjUFvmxeAHkIS+p0jILzViMwXq26GlV9ekDIJ63yIsajnzsmuA9M
8xxYyvVq3OpxWcUVTgqRX/Q+K5JzUmEH+Jp+EZBHQYeWNdN9D52FeiPCRCvz0fyb
roZwJD+PNzTwrtJz2rAsmbLwDO9WLdRT3+I79AywrjzMktDJcUT+zZlsUS67EF28
R96Erfu0zYs+psdplwAc58tpE0RlUXIhTU3wuQekvDI6V6N1UEVnNx0y8qZSBX3W
Uokz7tS4yJYPzN3vrizdLy8F57L12Phhg6F6k0TYRArvAudz3l4cKgjSyrW3tUgA
qLSiiYtgloHOKao885wG9l9FEr4OMqYAIA5BzxkVlc1Lm796/0hMEuZ77z6W5Imv
zeYW7u2lDSwrmdPjrCk+dy56UJE2NmkxRjHq+F5PL4Q51DE22Wlg7nfck5Ezx4zL
RSh3A63Yepaz9PG4wzKVvgGGeZ63kg9W5rNhOUVZJ7tEV6v7rvGhvCSukyt9uPLt
6vWx9KIMQYuM0A3xfnmj/OSh2kcSUhLRuY54z+n3SKEu+jhqFRp1/m+9MPHu2Hxh
uHB9R7lYQ+soUrw9rTyG2euuxlagKIFndK/6L4PIAUyQBWMsjWlQOAXoPqZX98qD
02cO0AH+bGylvlH6HNvDfTov0AasPVHO7jcIvhEx5WGx60q+3GxrW0nPqGTeTosp
gtfn59kMb3zDnWRzPx0c6tZaM2bts4LR71Nck1wssDUJQEPjJKDEZQkinApsmwo5
nprtZlLC+EPMfJ0Pr2XwcZNSCsN4zea8Bnyrky6kkpgeJRD8nDALvZBr59ZEuTCB
C7wgVA+gkcNxeNL0AI799NAxtYDhGj1L++rm5l+oz/9E53H6avG3KPHxNW/4y2ij
qMtEC7j4bSJxSoNZlUhcVhNFcBfJPoZpkPpynx8VMTHxvWf7N2bzxq5w19JniJti
Fp3SckSjSO0qk5xWLCTryE5oEykkgzKJv0+cUv80C/62gpulMDC1HzP1sTTc2GON
/0VrjkO/USJXL7+cy/VN+OiFOUppnLv16MKy/1cBxnZQ3oeU+e2XAptwo3l1RkZM
82XB+6C8zPqaNXMsiyu9GdnJcgv87Gj/TDU4pVPcSvIdOhRIQqZbDAc3pWceiVK2
6CL2YMjUmUH9zY+nLmVV77P4Y6rdX70zwj9nMSdFNel0ffYDwr4RePdRJPsrKw4h
K4fOYR/Hc4VwU6ISWzYUYx5X63axZRXDP3iAFw6pbxEgUMWTJFbpH2OFEr+lu+IM
EKU+u1Fi7ZsNIBLE6seGCKv/9488b3wKZVwYny4fgm01qcm0lvpEbt1cyJrYzARN
sqDNHQNI61eGlBM66OJ+KdQRkFZWKsmGq38mptu48NheAhhSCsiCfuQXlLXhpqcv
qqIrWRGlmY8jAHWUh4HXlChba5NcK6R4lW5lTrXI+tCwvoScz/1saRt5BHm4diOy
72QNqvVJuP7KZDgZgX48yRzf9HG2S9Vr27Fgyf7gY9Nw0uwd/nv1z+OnbMkV/184
z0u7hIMumnbKypWcbJiKaUNI44irTWLFXT9qn9Xn3U7COU8bZGk7WbNiR9lBLfL7
lU4iLkNYtCqu8m0Er+VlyJMy8n0vDcvn9S78h1YqgfCw3naPsaD3iwc0PABuYZOU
EOoZ1Gbdbzj+SXBJEsZghlpoGoGUoF4GlsmKPeuBnqveCGqU9aE0kptHoqv7mqhU
d9NUem/wrD/JT4avBEJ03dLRAOZQ3y1s0TJXFDwrH1wkBgXFa6rOUhiDQx37fRhq
jWI7UiPS1XRRrA18nUhKr22Upezrzf33dEvzDj+cmNw9mr62ZKPwT0KhylITfmrp
XoL5mqRDnLdQupXibYHCXbLWlpW6Fd4BBUpJtSQ50+ja0WqtzRv/95hamPHupMdy
mFVk1uZFBeeRI62t7BhvuD6R5WnCqWVmD62ggyLWidVpnkkvhnX97oUjMjtQ23UI
eOvfrDve9qM3zQvSqa1Q+nXTR8fmyibcPkmMollPqE6WUTFaz6IUvq/eOjxi9srM
G4bd8YnrCv8Uxt6cCw73IkXnmHXDaFzWR3fzG/TsIptZcY+/TyrxiXcsgVIJpGiL
aY2y4t0rB/BxYEmiHJ6KvaMT8EiAvDqwn4/G8C5IZ26xCLcJzi/txQmj0o0TJlTA
/Pa9393AQyodpScyd19a7XBdi+aVogjBaOUCzz4N1i+UokdZbbg9Zc22412iZLMh
9dU6mf1O833YIbzsWmkUoSjwvi9pfd4l5sNKkIh0S2HoqvX+g0YasfsEitA36aTX
QC+gqQ+v+72Tv3m37p2WAgxCqZ3E86K4oUuU8avWZDfRC+Vi69LKMvbvrD6Vini0
qWD8sKTvx+pxDQYyT+y4ceORfk9CCUsYfM6CRWe123B1eTdrjOeYxJY9qSWySezy
WBh+qhOC7Wefcq6oYoYu9NcdBPjWVmvegeGk5g/JxkuJzMXXiaXsQ4COsEjF4pP9
K/HIC7+DQ5hLAsq8OXOByv3+32MeSzQ/9Y66gg2enTwyx/qcEypOMdcOwrhJMoxo
MfbJH0rGD+3SOFqUknD1s2Eh+/nsq8FClFxzHROjbDE5FQNmp+NdT6EkzCecyD9z
ER86RikzIYhOzQHdJb2dtQWN4GLeYF51ksoFRDHLeUHzKVLmDPU1PTVElP+Sjjzv
Y5ET8xK+DxrRcG5FlexgJox2HORSYs88rD0k+92V3pcF+y8RWac41DWsKC/6pgN6
HR8GfY0hF1qXNWsdE6R+/hWUjnxGL794HJYENmzMSeUcEZkcul+8Ja8asNqC+GCc
Lq60VXzePUXG0/4NAW7qtOSq7Py4fbNRDseXTwU5D3N5+zT9ZoGgF431xlsOH6zG
m3IAgGg8Gk9qJfAf8h899hW9NHWrvP9p891xLtEzQZ34+ag22wjDOABRZrj6CIp9
KStgqehJSN3/RTjn2leOeum5DSt2M+DC8YbOfKMy/lYWZ230ZRIR49ufKU2nE+Qk
hEoezfD6JlSuq9h/ijMX30VX4U0ya7zPWY9H79KojAQnXyZu6R0AeVW2ZrgfNY2h
ArrLN05m/0o9z0f/flwzdGYV75mNYFzNmW7kKkO5YCCqJltRnknHalIfb/QM2YPa
Wuj1BH0k2zxRmLlSVPFJd4ktdPdjFpUiuOkm2bFbZPr8IFdwChU4qUMAA9Bzx1Tl
LlicGinvRPqVC6SLN5p+P57n0UcRM8RnHjM027SkMlvzKW3q/gekaa6ny6mIcFtA
IMvTg8TeuUStzpXyVImL3bP0cdQCh9Xh0bGIHyh48Wz+rRdaw/HF2ZOMknz2lWeO
J121hVlmXe76Yq7M68RxKJWPhg97NO3UKXiiMcg+Er1PYj1FiYOMqhH12znmOSjm
qlrRJGQBc+I2fjFvv0hcSIHswYHpSsTdwS7cINf1jyHxM1c/QLEywuEd+J6oEFGE
yWZTnTxZ+UrOsdoR+FjXN+e8mum4h0jdDs+pl2Tv64Dz06sU/BpaU8boSXaYvVg5
khZhuXGJyHaW3r/I1GbMr+w21Wi5VpqdhrcY3CSyxL4=
`protect end_protected