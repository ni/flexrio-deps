<<<<<<< HEAD:flexrio_deps/PkgNiUtilities.vhd
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 33072 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
gjQxfoUVC1+c91Q8h6upBuGUFNpvL+iM5pjqpOyQMZZWh+iBLZOSfm4PnfKtfZE7
5pJXsiqbRVMmH5EOA7nhC45gJZw8ve2NiQBDQTdPY8ThPpuK7iRfMYJfXOxk2JNI
Hz4IwZ6ez/ae8k16+3mojvwYwehmrijAv2PPl26hGWRZ+gmKYIwbp9ISC80S7GB6
m8vp52FsfYHVkjn9U1CfhdHT4JEf9E9jhifjflj9FzVHyjfb+fZVpI6BPDOzSy4W
zUAwXt/I+n+0JMepKH7ZrwvIZdqVVt2XvEiSGmB3/7PO7N5ZjaBpLwH8MN5aKbW2
k6iCM6MkgDVBCZIB+SMmRzpN+Jml4VfqJK6MM/gKVpm7QKb+C8wMRIsUYHIe0xrn
IeRIPXximeuFuvCauNWB/xkEyXNia4TRi7FkyzKvLsP+AxOPgmziXsq+jFe4M7Oh
VkfvP/iqI6SR67dKDafdcRWvnk3NUjJ7vVzehBV1HgKIVrpU9/MCzbdryH50XMl9
k6xWedYXj+Voxs2h/0VSpZcCkWjaNbITSd12NEMZ8+jFQTnt0MH1/XOoGNkpbUcY
0Cfjj+T58eUI3MoT3kXTIBVml6Eg/vYSWQkFmELgAyyLLIJJoOLgM4PJGTYNYQHO
xeVr1CpvtdU98woNUIhJoruEsaboXN588QNwg0DFmIhCzmLJC0PE6Rov1C4YjLUh
RT1fkrV750JeeJZjVlWRyqTm2l80gEd1qh4TLF2pqJmJ/ad726hr7UMcyXnXLADg
V/wkmhDeNS8pfnb7/zsRzVjzMnTuwNcDruo60eF1FjqVfXalBOw1LBJxqxoFgSxr
8Jx/LZbb5X602yRsiHDPEziSgP90JPs2qEo28iL1bEdEnoOOOZZkWbcOxYhD651r
1am0et3lugpcx11ZNG2wTFZ3Q/Z1NLT7jlv+h8u6IoNwaK5+ByfY46p6rW0x07us
bpf+SJcuj8qe1PZJu8ydL969SYMhzPAin6cIT2lG3XwZgirkVKcTirE6+YqFsl2c
XFZEMVjZ+klJfzImrT48BjhMkobguUdJyunJQz8E4dTzKnujfoycOv9MenhE7XJF
SskNTudv/eOR50xb6QpOHuNJTzW3hTgpstkMxJrdMw9gBG0mrnOsmszAtFuLd6Qh
xxWzeLwzwxcG/aIoFbakm6K2Ugbuxrnd2hceCWG2uWva1hBj/jfzDunmaWkrqFT1
HhRaUQi7pRBXefug7OON6vHtublFllb7YEOeWId/rpc2JdHV/A6VY9wbl5t1hojO
yX934255BscXuLEQoUfOpyutrFr75MW+9ueZwYHIdTPPa3GqJVJ7xYq9dEnNPvdi
vsf7Ll2cH6HYVqFft4lDeG6Jrnh9PhY8psG+mY+nzqJK2V13l8jUo2ZbIeaqXh2x
G0NoeAFCBHSKAWTl4mk1tZHtk0uwyiN5hwEXNNAhDVT/R0y6efqHjRup1k32iG5w
uNB5OHI/EpQ6UJFXvCh3Gf2r/3QDB9c4v7ZL5//RrtOKDRK/ZaxM1xfcw3paWcK/
87SjHTeiUcEQ9Zh6L+YHuKGRTUk74++GhSqYG2NNfkS+z8jTwnV9Gnbq7v80vtXe
yXkCApWOutdfKAJkK0g0rRGgNDBhZksoCSSVVhe4+0bD2eC7D2soYhOTkgw1Gm2s
GrNUYy4/sobeSveQu/QSKHiWaiRlRbfbZDBiXiTgJhD/jP1IAnLVA+zE7RWP1dZE
l3lTYSJGc9ayMw5uOz/ppzSAAnfugUxh4hJWD0AgOsSd4XPGfq7yT8lsFM8icCXw
jJM75HXBER0PgqWzB+50tx7Z5nt1P+pOXMpLBahRitfhJZjrGtbs8AP205yM4HBk
X4JKUUWUArhiV/GpDqvz4SkfJRwltN/W2y+C2j3jdqrdGgzzFh2J1nqJkjSRv3Sx
/lx6eQOEyvRfgKruhEHt9j9Uy2qbMVhosMpoEC0Eyh9/bSPXgykWpnnjNeIxw+XK
Xm4wVhjzrRH12IpOpyj93sb/7zIoVB2ur5OZKaUMEDww3GVxe1x9WLxj8nQmkn3m
YNc85uEzlkKH3uc8n1OVNYcs3OLbbuDSMGlu4p3S6EgDoF1A7d4OqE3CwUA6p2aM
IRxRfzLmtzHpN99JV8A1gVpmUf/Nl2zVUvW4YQQ64snEmYiqkv0P128+OB/rCIzG
ugwHUs4aqfXKcia6yY8h9lMNRHY6B8h0CZ53Bp9DQMjoqu0SXnwpQduYUwm8o3RU
fi11dZEZMi9byLJCbmRnhBUtAjOeBqdK8wmEx5T8ue0QP5jvCGWufw0qOfNOd7yl
XvWM0n1n2HVb4rSFluLzF696QQ7yjgpOI/zmqBNKg2UQjncq8jcluW3EM+N006t0
zn+6qCckIOXAZUHS98eq5mVJAno0/CiYN42Zi1t/dT8LaMhQioUJoFLbKxvBaL4C
jCmwv8WbKK3AjfLtYuuhL2Gz2Uvydu9fbIZ4p3ceeaT5KLXrTKxEut1Wdxoxv/Ea
oj2D9MiiLOZ4tsi4hzwZuU00uNMrjQuCSP9a+he/8OleeCGcmvE8r+fNYgkR6ROB
SqR990zr2ooa5+vN8+ALMIKgIb7D9MF5uWiVOUKbySrqA7jKdzPZyiXbtqJWzhV1
gkZfy4yShaJFyBrrh80sag90QS6pDcn3l7MN9M1OAfwQI7Ku5znjJFtUxPZHmBJX
hjQR5pm3GDUkBniUfINPNU0oRXdDew9/N6M1+vN4xTFuiRtxHeNN5Zo/o9fJsf1n
jKcA0jQMVJ7kVNlrCCQQoqzxjRBnCRmc5wNbOsMgpcd4lGk8odOj+Ig9UlWEhsG4
48Y8zLr7HosqAsSDgePC6WGJhEnOaHFXx2ePtV5OzqWnmFjqovesKtZhZ7u+wMZ6
X1KZgDutkwZxgcQ43aUSN0+8SNtRW/EzRhVr4G6EI7XNdHcxmJ5M78moFVu4am9e
te+Z+33uSNpxcRhpx6RZHO5DOvhed2BnaZZbnan8l2LLNs46P8uLmKXp1ciyEiAH
irgHasuQpWWGWhjm4hStCCeunpkkeUzWWRjuV/iD/FTdMc2pbz5E+29dykl3yqvK
SzFwTTwqTiR04/PFOyv2v+nSUYYKH6vIiHYOFUGWD9iMHEahd5QSQetXwNOIqpw3
EmzlZ32vtHzvpBsQHMuxwPCB/bvUjt+e+DNGOdL3ETdrUAOTbLTVQuTjPFSDYRTd
+4X+UaKpA0NpDH5CzSIVBwmqP7Y9RPp17KOYCn9S5JqlIt6IYfTJ8+No/4O9uJbj
qiBD+ZM/z9Oeyr2401xhvNA55S+ld60/jsvCcc+Ah6zGIrtUDEL378I4LdvjzPp7
froCxNJSgF1P0b2EbFgH4IvJPUxOVOnusisoaTfQ60NtNPlXQeabxf4cXXByxIOt
dxpY+8CyBYs0EtSfgmUb/tcw4k+98FefKmuopmNZQvibtU0GusebbTxrO0PUtodH
XC4PF2at84N89mnKQRRbnjSanIh54Z6869m4cE+L9uVJR8zqwAmiPrPxFhu8pVRp
Gb08Rvi5Z3YeW2SHluwxs/YiLWQmLtS4woQ26jZfgmSl4xkRBec3Mfjl8gBvTt/D
fO69dUa3xY0PBf6pqRaL88onmDhegbkGdkYy/GkUEq8tIcgJLLQb0ev8FZwplASw
sPBV2pqit9lT+fzCq6LwkQY97yQk/ehqK9lTDB7Uefz1P2bqpwA+u9b62JeBD5pP
Ue7DpMBMLuyPpCqfxNzC5KSD0k8EusmXtZz9kqmmoY68PZMTZWk7Lq4R3Cd0wzep
22tkRaVf62EJneq1jL77y3ETmMBgzoZ1pP0YMqB4GGHA5QbsKUvEK3nx8VtYD4FO
JL7rsOBxBGLs55yrMi6f1n6A3Jb7Aw8Obtm7eHbAhFIo2pg5GgTGcYqAsrbBZnbz
5NLFO82/1bZn/MZ3Zdj/hOf6p0FQhvczQxicNzxmWua8rmaRlsrn5IOpvFs0GViE
Ka1iQZTRORtmoIfaHFsWEkSo/zCQG7p6PElEct7zE4KPwUT/jHUraRLS+DDbuvQN
oFr4BnmN3FUkW733QnQH3EsJVyo6/MJAlWH2La7Zd342Aawgs2xwei+ywKQR+euF
W+1yqMHLqppxvgfIloNmGiTYWAUrWRflYhhE8hzSXIl+S7kL2ckWEsmwhlwws8t/
mwM6CE32eauQaECCvkeVn6MmT2HVOTtzJrUzRwKdsOIbpK06n2M1o52HjqG6Jdwm
mPuzSdcNk+gUBgx3urLYKEU9NkHM9RtSKbX/c12kJQXFHb6uI4LjTpJDlFB09hjh
iCr14AFwliTcft8br+j+8TDyD++GQJAX38G9QO4QJOgC1hSpa/gXwE5iMkE2psB8
FMKvqAZ7OCP797yTevyC10W9cOYBVz44CKS/xurycUWtlsA3ndayKxVmMOOIS0lv
ijzHczDk9UM1zjQ+xwzhAPPtwgmQtEGSpvPa5l19LJ2yQghMfegvMMrLzVZUXG1f
338FjY1FYG9Z4v1QOZmVpxgaEyqoAapeA+pWq17kKh/aoUl0Vr3p2w3UjnfP2y9A
efPP1Xaa3iIJAU+up1ukTiuoeKOVSRKjBNXx3cHnANWq3hBlALWEApq0k1+1JfeP
3bAAg4uytkxwu3tHEBK88CFTp0bL3LdZ7P6nggnGzTLIo9urneR0Utmm7cvxaN6M
Qa8M49bSYu35U8CPw6ZX0bTou2W60xhafKDjgz24zR3mDvoJRGwnM8ApD9QX8bqd
MpjspouIchHsPbHFFWyFUsbIwUrwHvlj+9WEEpIRPTC25sPF4mDSXLsCzK0oM864
YfFUerrDy6jfEj+vlzp/gZz/GyYdQntTZEnyQFkeTszrMVoxGpC7UlTlNOvI+OCK
0Q6z25C7hPNraXRNvnCLVkXm5ZTFBB1OEkE6LTYhqA1evDYrEjjqa3YM/RIg8igp
48EP6zAKvfscuuI7gj/JpZdSMezrRXUWHNzXWsqNBcKn5QS2rTicwcQy6fOo/No/
gkqZBT5aqWoq6M6l/AdytSYoID3HA435MffyBzBTwxzWArdgMFFYKBn3ocNRqw8p
H++ZYs/fud193ic3kALJ7rsfxqgaqkSNE+iquc0obZ15LTtGuFi70but/GOFfTUn
/XmVCek2JcfMMG5R4HN9ZqEM9qrRqr3srAFHgqxFuNOqgmgIZfsTRngNcjCQIsW3
PDbn7rT2aochdDXg1EfdEMFCTElxSR+IayEPtP771SvpH26XxpR7TwIXrif51SLa
TZQm036nuz5KURMXMX8zqexPTgAJOXaSYjx2ZXN+REz6H5KBhb45jcWaGfTlT8Wo
YXQlnlw18pF9HTRGTJFV3T0dPxZqwy0pTjLm5oEahU3Mc8hMgH9JvrROwvk+BBoL
32hyOtPfOCB4siWZ7MwwUn2kgaG0WJb2E232uPdPHYzl74AF3b3hyeHuJjLa5k9i
vvPJKHbhlxvB1pWCl8lVIyuDmg9WgJ5E1ZNVVZY7k5QszCNNZ761VNW7/Xxd7EH5
qjWUrDV6DzMxjRuMlKp2d+M3oZI5Fyt2D5/LGYbdA9x92LLjfLNNWwA82dXT8sJZ
WRCDaSNjUrCHI9fS4jquPCsH3EzbTM8/uiMfCzKPpHkXeRtwNvUb1cLOSp1oaLrk
plyxW/eFK6T7yZ4j0V5ociEmPOSYoilkcpeZfslVhX/IaaZCS75Fjiw671HqmFBH
lqw6zq15M4MX/FfgyFm4sJMoSjGbQxS9OU9uaV/X9qeKfVchnr944jnqmnovcv/v
934IeMm91yGvpa4j3aQyMrqEAcYHgzXHfPuV+1N2SoKuanwjpxmvaydiqKEmD8MJ
1U/FrT6c03L8BwA3pfQDsUPqzU8I5VpFQmY4uilUcvS7gn1ty7IQGVzwgiMJJjQQ
0WY+deDUJ11GYXY1VBC5B4TzEhoKJKP56/JZNQZgqGA8R9WY7BXSyvkYM5KyKlE8
Ryis2LT7nzqCzZfxUfH0UFZmKn6tcjFXAE44CohkFpj/IYZGlSt3Y6wScWwDAhiq
91/nvCCPhrHMpGGqbwVVtuMm/iN2nqzfpyeHkyajiAgNsvjj/hq/1wiJ/3Eu0qeo
ASdpHffPzVNSx9ChcQU8Px07zc4jyalojaO4iJRoAPhd22NovCA+V+xTc7n7dll1
tZo9OvP0PmB2C31E/9IXIV44x2cttZBJGX9MYeGOwbNUA8I/vWetaas43ESBf7MN
vwnpmU43AKvFQ6dh5Q7CGqqU123afIka2jEdZ5v0pC0r50/P/g/2GNLPKRWywVDA
HBfaiuU/1zL543uenrpXCcb9FIMNCEDLwlB4LRISLIj/Xe0574RlWKPrMLllxuQT
dUiDOOGygGx6O/VY12/J8y6RY6mSCoiSaUED2mqOVQZzxu04pmuNLMk7OFjveihk
LIRgRGSQx8EhR3j8s65jO4Obqflwrn6wFnrsbNVXNUmjLwv2Ip7TxJEYZEDgGktE
iNeNbUDj7mS6MqQxxueTy3oqdh3Ge3unDHjPGM+FIIQByCN8Mg7AIG+wVrafwSH3
iNWhvWM5HDd4e3VIxzzwj56wvo9+rZQ4MHk1gq/5llWZZiLWbIEDkZYJUJeSeM1q
ar9qKMFXyLVbRk52CZz2tdJWkeR4eDhbZRgYJU7fTl+FklB6GI0gegYkGULVMpiS
fB8xQe8ijUn+5VEae4BuyfdGeZJIecvz+bTBkA0dMQGYIlIZCk+RbhIz9UyoVrT+
Vf26QdfAzbb31Iilw9FhNDYWJ7hBTIh7rsjeoVL2kMofqz0f64/kCKw0tTawTQ8a
+08j/1EcShzz8gPKbFWrLOP4N0k0xWSltW/pwkiqb4+8kdZyQqq0+YLZwS52/Xso
PKLkYE4YEml6IsnaGyf8SFOX5Yps9/U3TX+QG2T7OtEUMPpHJP1mzxBYTREFKJ3i
NeJERX6zNSJCMbjYXneGRDy/hQh8Zyw0VlYg0awZMvKH6TVapjyOvudy4JI0Y3ji
sgVEu8NBBVr0KeXleOOZRwQskT5sX0JKG3azkQax0MfZ3o+FvIFc4hA++DXNf2ZP
AKn3znjWgpjhD3AZuNAcQCO4hzQeUDkGlOJ0zo79mXkVjQhI2F8hbfVDZ5/RGIia
yl623InuUWzNFiNoIHemOb9E6CjhHQJcwPdDUOvXucNSJMNhBEa6umz1F2EaAklD
UvtDoERb6+SKDeeAFg2TaV8ZLG3huYWIZogyFJc58EMW1a/xFJcY5Pra37pJCbuB
YG+TnPUUCVG9DVRbH29ysfie+B+NUt+wE4J0TmU0+h3GG2OjgyIdOrGh6dqbSdU/
l3PYyhqiSNN489ZBUo6J8EFWzBq8MG8akCSlrozjqpyc/aFPGdqmxkp6AfiISfjs
Md3WRSbbLILBU3se+AxjtcunQVUOw7i7u/28V1LB2x56Pd0G3d8XZlUO3GZvrBie
iwtqVjKUVX0btOPHTQ7oJfDNALMfkvLhl2LHmZhF4FrinefwFuVfzbWCHLXOw+uu
GXGji8ut8Gk+z2RjB0lxtQx3HY7fwSIHE6h0Y1S8ZEWhbdcwY7T0xyUT+ONBT3Do
2LgU9QBt/1f9Di9nhABTRgLP1ssO0kcoaq58h3lLrfGl1/klYKXtEx0GjjHUA7up
zoB8rBzNoajxSyFa5fNom+Xp/7ylIOWIrfhRUgJJrTAJXDbfI0/DYt8WtKvSne47
QIQqRwnxP2q7q+/oPpQiuQwP4Cnn474rjTCi404h+vAVxNbg5aE+PtLT6XAvvGwH
adfTN6pV4hEi07bWeyVU0i4Tk2ev8FWZLYrEELbvBB3YmnY5+SHgpSOm/SmjuRHX
M+09o5viIzhR+swk5HcVKQruWKsM5OzNlyrzCYDWCjfwotTVsGWe7/SO9VumOT/h
hcqJwgDdchUWn1Dy0wm9valepHK0YIGX3+OOTusup7MKQCBxoPc7ni/E2JsuD3eB
43+zVxmdg4M2TE6G8INNaAuov6MSD6ChAxEOSqiiAr+CkffCV3Iz+TYfccSmuXZr
jwozsTfRcM4SKGqO0Hr1phXBXue5z3+Hlz68/E/jiv94ZH0h1bSsC55WXqd0YRGA
b3s/SBO4HiHnXAI01/8YMSXouwRWydWXfrsxwDAhFrXwzZ1X/9Q9t9v6Hg500PoI
D/SP0V8+QjBWNUqio7Bgh6MtSADuDz1dDwuvR95C5rpxBPEwLHCHM39ocNXuvuWO
gllrYI0oxs541UtzJic4B/nEUi9PCL8kAa0lnEs8+HY+MsZjrDR3/fB0lin0rQfT
MVkIf6GgT62yHQROVaJNbYqhvi3W0pDQ0lWdLmTmm6a8WPHLgNm8+DlZPoXVeocS
ffvjC97/amyRahn5i/1ULBOu2WGp0WjSp/sUIERxe3a2UMCcG1pdqbOgOhmQ6613
XKWLlceSiTTqO1Q4vu68k9jNGtijPszaEXOGpZhe663mB9nZJ95LLZP6pkABty9A
mp7PuV3jZogeunTjIiivwkNyl6h8R6BujhddYO9W7BPyz9KoAwI2YIfR9g0N+gxs
YrQYWDqP4VO74Hr1VhmkbEttqZyiA2AISTbLrSfGEyWIwu+roAeqHYk7lE3HHzIS
U6gnNuIkQk0LQrE3klgL/v2G8XuQx4jRcIr12M7wxrOJTGVqP3ImKb3FadtVrM1a
aFP4G7ft0g1FQ8to5GrxXrINGKGGrkKQ0Dv0w7wzligTKlAuTs0UMPD42CVnANev
BDIiEJkqv+PB4HbiwX2pXeOIulZtA8VZveAXbKA7SDsrVijzpUuajIbhl00OMQ0S
4w/+Bjyzwl5bMjcnYDjjPTKdFW+2l7xjFi0LWmeyIRpSS/1GZ6tsSD7bb0nXWkTH
EbaPU2tRNXdfecjsiGzOHjnzOgmul8alDiltsEjZuExtedarLU3nJrFtOMMEIH3X
MI/MoCHzmZNEZ3vfYArO061nAGp/nywkQlksTFQ2fdILt8tDCuhM3GQAocwSaNja
xSmOxguUg6PT19UjCWKQ5QPlIHCododAB85RUYKqoLs4tsrpaTMDWs4H0Q99wxoE
k08mm0X7Et9nRfwR0g+DjHbnBafyi3UqrbusHzasrl5EuG/2ETz+2F14Ca54WwqU
YqTZL0HZ9xRV26oJf+ZGvHmLDJc4LNCf/pUoqZhGF1OwdQ72Z2LvQDnPrF/XmA1R
gdkFsUChrUqVx1nzgjchsKIsqR/DE0WMZVk8rkebbyL+VMQjxLPm/8MiJTVtNUjd
/DROP763fMKvC9mzTeOI64abw/zq3sZia15Pn4jBXEcOZbFQgIIx+jPH35Ak7clR
0aeNkgx0HArrLLh2b1bpJPHcwGt3rEvrec6hQ82MYx1kdEedzFFvYwP9y4hLiI2+
tN9viDWhTdTK1AxvAxnG2xs7nMUMQeUnQkNbLxlPAdmqmydhRPx9jGWI2VGU3qT1
vUIaFceRXH3grHJcDcl9Z5cVptSaSWCGIzQHSz6N9447aM6yVeogTyAyjmStK0qf
GA6rP3QjdK0IGAZQL4sqSjnbSHl9+hQ5JcGg549fdbOdz1AnbAKJUs4DElNLBVw+
9WRaT6NE9z1b7tKVAAs1GomT+2QaU28sIDaIB/AJ62Y3tM6hseMhVThj2JSU4eZj
2xaFouUsicItV4e8vxQcYoNO5V/R4jw0in6aYkRro2MgVF6nzmfKhbd55abhKrxS
hpG8COSekYLWsWOBiShQaA9XuZ8QxVlyMUSbt/zZ//mE1cwBtWjr0pdVYwtid+5N
wt+ZUmht1nyydrjycKO/Z4g4BsgQP4DS7rHN53ht0Acr1kkdAw0cREYA+GIH8MCF
/8IWIxM6nnHLFk5Wz3xoPOBXt8t1ibXYfS+yBO9tkQynLHhpNmMhhy8Nz6jH1FdL
Ez0e1/qwB4Sz1WtsTH4U8KtoyEw4CxEHEO5zsfwb6B01yqeeEy7hqiDnTM8zUwuu
WDq0gnILGAFUhFRmRp7SwhnWYk1mPhYmhp1xtkvj1COq6aDZRYZSSMhaIVcV1Bb5
rCukXfJRlHVGsuGW4rJEmi0YnkZS23JcPvMA6reJvYYaXeuhSHzY+GjgHgtyC0Vb
eTmmWhOFKJfZwcGeYTONGUEbEeWByArq6ht8Jp8CNq03jEtUBfuquvy3xnEHJbPn
0t0mXYFPmvO8hOkjRvfBpyCiOtjmAmeYUirabpB4zwB9essbgPsoW+Tiq/DZpNgr
eAKBN1kUdxBd/9BuiKmkg5KtDXPwmD6hfXIv/r/FxW1WB8zmz3H5yeNnMe3R9NiJ
BvmX+LJvk7zYBne27EuSoWv+tutHQNp9NNMkqkBFE57+vRpixeJuSO7uuo/tS4tf
Oezmmd4GE/dMButxv3NF6rp34gXBQdqD8H8PfRGMwKB5IYqX81QZV2aF9204xx68
makXMeDtSyT32g8S6roKVrsx5oSjN/l6fNXc0lY/cUM+gcsKGJ1lbthnaCBvcg3m
lJBSh2AYd8t5awGiczF3AMxGwNkFGjrerP67OKsnbr8PvRvEGoWzlhGhXNyk834l
mq+0jpTEJVF9fEJG6wO2HWvREK1RgJ3F7I/97LNHsSxztyzNgj7FYNhmGxYpSrea
T6r1KP0OkyFUyjuJQAklgWva817/k3lw8gx7wtJC+r16ZBG1smJYKTe4Kr2nMIhf
LM6yTipHWtu0bSjaygNdeZvA/R1a2OMFcfVJ1QXWbWH83PATzFm7INiUbzneJ/zD
N9nUudUOSIAwTlrvNSfLt6V5gjHbVIAAZTwLKYDfp7PC8nvuRW382DcthdDH0ICp
v+SDWRltZ/qhF76P6BdXw+5CMmbFV08JrdC8Dbbmq6fIGxLEliYBWM/6zyfyU1Pv
31rAq4VSbWotn8PS06BSN2uyggRtgnASETO2t+IE86SpgD1UvM3/KD8TU5XJomYF
ilpO4JnFS7xjlSKQeNhVDVVk0aIoZcOpuYwVBGBW+oF1HNd8Zap2q/snjNv9Y0pa
fea9R2Bg6wVWq9385rLPaH35O0UZR4VmYdaCuhhytlWUP60mPMTitd8iC9Dj//Iv
e4jrQlSQfQK1ZixheOz5MviGw+aOZ45JKxW6M1AO4jJlaOeDPCXGHXez9NNwz937
o4aGd58coFAdwg1YWSGVprFEt/ozYhMvO2CnJql938H7VJnJceCg6sQDNI5eESbp
ds0x+aVwF2Cy84LBKfv26pt0fdoeVaNRIkdBfXKRwEp31ybakQPJllEXxRfll609
2v3lHnUaeMfqW/eIlbwTAQo248XtLENw4s9I/ltmXyp77MAwHxWY4UDdaXb/++VA
kmQJ/uc9hgLd4PcaNOJEUWmG9CPdc+NJvZTitYmUL/MU2Y8VOhKfjYhiWVbq6Eh1
IdZCU1GnP4vM7nA9ivz7rw3dFhxwvtYg+ZubmPVdn3QwjX/dz85JtxlWlGd2wRlF
mNCntvD/LbQ55545kHdX21vrbZeDwYO4wZjNoNf98YuNSbogel3+2ytBeQa+MQlB
aKxaRLeBkOdCFwR8gYRWN/jFtWjdjjJuxrc2NaZYwiHYtssxny/PGVkLQLYvIB6+
UCoqEk2SIbNMH/Uw7ZHTKy5PYrm9T1PhfOtEIov8oZAyRXqQcKZrnuBjx2PwmA/P
CnkRVsJFIxugune612W5hiu3TSmwa3Salko5AiCA/WmsxMFnxIoqk9czQrea83Vx
Wb1lTt7wv8bCvIwYdsgTH9sScXTaw7IMFnThZ+eUPsAA7UW447ZHKK0nvgKhl2Dk
B7Z1w06C41DyNuKHESk5oaDNAygKye3w7AUCO9ymKVqEwf8hqq18HQsp84P0A0Te
9YTVMkoyHiOoxv3ufVukk0nI0G/ROsFESd95KihnygkofN6DaK4RxO8jSdimlSPA
zCSj8LnWrymopzw3gBCZF5EeJusNx4zJXX0B8EeX/ZWhi/C9FysuyrKHmkjh/KUL
ne7WL620xIiS+6jgqKYI6Bzqauh4Wok3Akz2AUbRRfySnh5rdNUdEB/NLCWHglSP
MbZ5tHlUdfm/99qGpXQWEcha8YaYj6CZYRDFqrtyK9Yg9s0dkOw18CA34ccEwKYF
1NJdVGQPIqD7/eLn51Ematt/gcMOxgL9pgVDbMnVTkxrR1h6dVZH6rtqfBlLLtPN
DZg4dUZQdxfCrgFxrUPmkN/tFgljl0KSsK5CZMnRu2aZwVCT5eeufXK1ZL/Bybir
UVp8U5E/0CKCpa4hMDac9FSA24ybqd521ubwGtHgmW5igA8pqEuadooU2rmUumRx
xqpXnEyzxYa21b6ku7I3lIVom2rSwvz14fUHniK6LB09f3uuor3JCVsWsF1iMhpm
cOsiigQkLe+n4g6aLP/j9Kl9sYZM3dHG5MLVlQkwxY88wiufQsNaHerTuuFtfhib
6+iGo6Lug0veOoG7KXOs0EfCje1sISpjWj36qFwWcfaSt78tfDgHh3OUZq9cpON5
TPNd7fORx5x0n+hKiKZVigAGULRJo6ZSwxgOxoSe7pyHSzDEO8EjvzDbEXPL1Foa
GfYxQh9l5nVSwiy+LmtzmJ+unoAZPKSGrtRiaAqqmhhnVCC8DQtSTfNM65ygxsNY
2Gs3sv7Ul4GEwVepCZMCXMj3siSDD4GgqlKrSkXcEhmmcY8QpxQx6F/rcPEzvtKB
QagVm1j1D+A4783rH9joktOzGrvke+7uMg5pVcY5HXxf9GpXFO2eC/v+X+Jiq/yA
t7gsZ0er+yTMm47AznQp90ozZZmtU81x+Tx4GYUEr4kp5dX+L11QakVl5jhsfj/H
EfPMknhxOdPiXYxHYYYIicW8FXYxUjk9ibRx6cFqP2r6FgwA2MXpSTd2DhCb/zJT
r26kYaiX/cyAV4ZmyVeR2e9SOj59nRn5fudlmLv1Z4NV9Ey5Fpq3CRl66WNihvn4
ik4MQ5w5CZ+Rn2ngDrF6yChkAsnu8LntG3TmB72ZlFzxYvNMvO27U5GfnDNMzFDE
Tzm8gO4oRKDKaukVqtZZR2qyQfgWdF6YjGK/LYXzWxhUr55qXc2rORlDSPZj9jrJ
ELZHkh/Q5VZdFsl9BLRyeVhlpn3Fo85KN6tW/FkEydxvz+Zq595bdU3qE+1QrN2l
dg/tvyBmUhD0qoDCa4oNN/xX3hGBI0YYZ9Nf6+dIqJYlI4+TABBIvjGROBS7IIyD
x0XptLy4Ea40lqlRqmtYuF0k0b7bKxX7mTjskl8ngjZJsC1XG+kVpKYT42RYOSse
6slSjNm5eY887WLcN5uflce6LhZ4oD/cVycwz+whlSEKhd7YVdnSll95ZAXF3ZMQ
DnpDehCwScPVG0jrrK34f1EBZmWZWQ866iH2p4O0oimYfPsl7+nLdH6uPOUeGlg9
5V7CrXmvNCTMqWVDNLRa+5jFRjbJvbTRZT59xBYN9CzcR/Y4e0gDOuHPEVWv1Y0H
NsCOaBkiFGgAEMT3zN9Bw75gA7fLRdvAp5tWdNVtHnbC5iHkKHoo/sJirYatTVVX
czsZ+Q07AVLT6Pj03krZsJmNCUahUnxQkngZ9NlK8GwykMz+Yrre1PrtT2kQwitw
GGPJbaI70HVXLZsYWJjadqEt8mS+pFJG05kekNMREh9zhRSY7m5FqMDJxZ8H81ZR
rDzES32MVwzDjQXhwjL13EldAFU5D0FKNKIsGFMB07iKEBarTDu54smMY0nxtVIY
rQy54ApJPxfJ5eM7rryT9d0ExJ9ydP1IXO5bUoOGtmceIO8yq4FC3H9tcufOXjMw
bYN50wF4+SRhD46OHS5E70Ee++Fe5MhV41tFRWvd1vI9DqX4b6WOJpCA7M7+g+Yb
DeGSrWRbfb83hTJuLdswc2it7XcYy0DWohpv7rEUvomHZzqUv5EH0lTF6sVcMHwp
DaLWNxRiU7oRW7Gkm8hOBH+RdvmjoxOBwAKqbP/FLR1OgiGqdmH2Uox6yvKJ3SG3
WdAa7JmHh3hvtpKmWjZS5t3DEtI7kX03ATqrZHXL6FoQL2176CR/ifm2JK26hE9J
9omiWsQb2TALv4oahYFwOphX9ZbKyFBgKZ8xHiJzm0mj/7VSkndIZUduCP3FYgDw
7q+mREdZMsBnDdW674NXoYAf5c7ERY8oI4bnPlHARyXwPR1cvn45R1hOrWEj58gB
TpRUwaE+C3RhaHumHHl5BEs4o5Bwf4muqwaNz3doL5v5RTyOQL/FkUE+jujIeOLE
zKK8730p5cHrF+OBrYbppakMbvu2IbKmPOqzZT9PXGTvjz2dxWeqr+D7r8ZLaNED
VCj0hJx7rzCtCwgGszKk0TMFb0+J+VuLesTVjf9kjNPzXKcT4gh0bGIY3AB4XR6m
K2X6Hns4FkF+StwluFVIIuio85RyDE75e2hc2aZLfEbUdmWnH4yj+u+ldh+HyOSY
RRUShyYOGat2ijghjRBQvYUQBzBNkwJAX2zr1BBJoULzSjYau5QknlinKMYY/nsI
lmKDHfxgHKYIGVv9fjCieaSSWa7cYEt4X4Q1fbrAMq0KjXrxzo6QiCnurheqKx0z
J/XnZixfKZnj3gGgBAQRFB9/a9REcsIxAoT1GJ1jhCjAd+EgHd5Zj7au9MjreWeb
0vrzwNRv0IONLC+ZSBpNSKh7GlN8tez0F/jza8aiYDerEDdcmnMfDeDtlCA6NOsR
wo7Cjqx5J8CbBPkSKFEhvdmpKyR7ui26qo1ZgBoQxywG0JBPTflTnkFVBCL89qHd
fJTyOu91CcBrQut/pi6pEFOWoB461s0g/7AAOVSoZLpennnyS6OzOhECFScBDdMq
oiWBsHGBRzBK5wmd67iM6sZ4rtXunNqTHbGtgKyIT7Y0F/zNJyUuztgNrBMGCL0u
pSOEHF4m47+hZdJ+efO53PxwvarMRsdyCnm6IlUJPQwQ5qS91lqFqd8p8phfNWm0
ZeirMKaCP1Ns7NkLzyQL1o+tQbRvyaZACAcHkG+JLL3MbXGN6TZIvp04kzyaJS/s
N4HF0+o5ra6L+BeZtrOLig+/a/yNjbJjGwBv6pMjIZMe/AoX5M/fwldWBRAR0ToF
CIOnZVOMPsdHtnV0Mpz8klibojZc1CEI3/wGIfvAlKjltYww3+plNOK99qd/UcoY
SMfYptPe0+DkGGIPHiWsN7GKjKsVuK88wof4EXx3Bcyb5xkH/+1mxLIByHcwd9g7
W4fM1/QhUTkn99Vct1B207A30T4W0vHu7eTVDsA1bvlX9qdmkKnA7XQ8/5lWGRMI
pZ+ljqCeCdL1aeLOlYGsJGfzBprCwhsIc9cnAGavDvo8xoo1XeaLhBxA07cjCOLC
Om6o7aGAFmBA91Na3rZm4hvdWEkyEG8j+WiJ0pd5AmV/OqE1utgSN9k6khbhbJTW
giUhGzcLPgpE6wmBjazMzE/nl7hfkAn4+KbztSxkoxcIXqX0GIfET+uH39PccTYH
jJgy2AeRsYPuQxOkSF/tKDKVEKuc5syQ4xUf5TSqhAH0HLgxXzTH/dGgxFVbQhOz
EdBf0jevmPIHAmzZ7zC6mAzmwbXUaZszXn8z0M9gjO6AykN5pSabRotH2Is4w+pi
iS5gHZOJNzS7AMfvTTnXyQCCtmAolkSi+tzaIbNGFWjN326bPMWVaNk1r/UWKHRk
7r3Bf7pzcN9Y7Neaw2KjJOoNQMvHxZgHnrVFR251lYRlZ4+B6TFBdOVRRUWm+GRb
u97lg9eGfuk2QcLk64XDf/tzz9jGkHhDdpfNKxP6q2RTp52TIWdCaVox2arKBeYt
6A6OcQ848QsrFNDfb69JwnFZetxlraIp4LUTlQrDPCwvod7PAM0P6wl/k+n2ktSf
tK0eLQCcsao+YyMywdl/LDQtDBnfgVp3PQo0hGwI6mO5eT/XdyiiwG7lsCeinPBa
3ucSPV8Sb9rV5G4ydSl9SfBBf+TsLh6zysvJ70RHR4Bj1N2f75/rqG3OzaWHAoH9
iKyoLBhcUw5PMtpPvPUT93myPGUAfXA2woDYTyHGtcWVaxg1pi/Ok0uAMlI36YP0
KRo06Qze0fhpEeJboSWussmz9lyZNea7zGe2YaQG0HCoqkNgCmimbVFYoV8qZqtq
422o3wtl2i+CFVLnD0/M0SaixhICyFWh3aXjb+r6fwb+nz6UXptjv8HBel7qt4PH
4bQ8rP8aTqhqbMz8Z3rcHQ8p1g16dlpsAJM4efOzxXMED+Ke9bqTHOT93Z98vTkd
cYeW9YQVsY+Xt9n6NZ2RwlH2JjsQIhyuZGqszyzBH7MKTifqDPWtin1sRpBq5P3D
ZYW02F/ha7NZ64r1Y+mKdBgAHooclN+/KKyzBS2E32oEvW81HQOM2a7H/OA//Ne6
6u7TdIW2bMQNuR6FFRCCXgAIxvsUAwQPxbDj2J/vcalKI1ZniYAflU45jc/446+C
YP3gUhlza5OBI/DiiZK6jXWw7yBv1c+CqNiiHy3PlDLMCIF8tlIRpiYDh9AISk9R
YhD185qCMHc93efbui/7mt8Nv8znJo5latLbsxlyBJ0NzUrw2hHL7XH/McMZn7U3
RQ2J0YWQoYacp7DjLhgeakf7pNw1YA/+BfT3ZP6a8rgzKZcpS3LbGdyzyqLBDopi
B/rWqTM7+V8DP53dT9gQDO5B/AZQyLYl4D7pKubQkJv7BX+0uUiIngOi+ybPOKJy
vst69lGVA6AaK8Faewt/Gi/AOcuZuwnb7hi6kDvRvhqkB7U/OuG7caNWGg2yMhem
FIVyYFDeWLPvFqvC5XA/xLYLIf/OKCipUBLWSrn6O4viPzWMagyhwjoIxoiLtrpq
lZ9ZN96PPdwRSfbEGqvKmqgzVLewNfjtMDLnPZnTzoSYPK1jBSNQhAN44VGW2MvL
MB6XlpecgZko2STDvHH7zaWksfLX2YeNiStFhx+rJ3921XX/P7H+AGZKmoV7Lobj
3zkj844ovjd4N9xSF5pstygG5ett7G36J92DCZrfA9Fzg8543yY4ZH0QjluV1Crh
u8elUSIRE1fj3hEljdgnGEiAapQo+ByncgvNhM+tvlFzL1r3kQT4RC2qB0BsvyQ5
wplwAi772ZDO4a48v7dXTvtJR1J/F2SMgrxW8BPCFuTBagnVJ8VlYXAvzdqMBkAT
cEoMqvHH2imbKBIc+t/3/Fs3ImnUOwPho4NUbMG9j32/qALaqbsv7YzhZZLUKemX
nmsYLCxIUzna3LdA7arX7oGYd4fjXdH5Sai8a6JU3oxJkY5s4HZZAY/dMbWvk49n
aJb1g1qbX66sdcccKyAxUxsZJU5qfzf5i2Si5m71qWWkyAex3eSodjkHt+37XyOl
u+n6PGUBqKuhoTN/cPwF/LEccce4I01sKw4YK6IJGrgVR79/37AdVLB8J3pwL3qu
8SYGMXU0NiEjZqBbCiaGeZl050erMo+nOwB/dgBzpYqYSl0dGNsdqFZDNxgYSB0A
gcRSZhb+GsMLqQanBzhJboAx0Ef0NciXW8uxnLuLNZd8s5Tg7ko+Tn81rWh0i8qO
o3Jlei1EmR/bT5df+drOS7Bf06/323AnSxZIpxOfAIkAGvVqAZ6tY/mAbFW0TSp1
WIb5tdYll0r8UOKmfQQ4j6eBkCWuMTVoGqn8cca6c5f7AarHCLlbdSWiU/JV9ET/
9IWyBQZqRhEmN5cR3FnoxK3vUciPQbUZYFoUWEVLuM8Z6MhI5TM27sV8fqRDcc52
RdONL5xlEciG6viDlS1ylJyZ21KVDqkau94B1cmbYMXIOQMmnJGFQhlFpuQzjKfQ
xCw7kLjhkpEDSf+tXwts53oQcGgAdkAoewenvjdA2A/qiFJPWvXkaG7q7pnPXxe7
sUptR4PaMasMCUUjHEQGnt1iWrUomAY/9tHc2O/xcXaSnhe8gdhGJFQiHAZ6HUf6
I6J4Qqu6mfQ6XYERCmVI0AjJ75f40jM/xUXSX0C5/kzpApL27U7TyFtC5oOO38JT
g744yi81bvItQEM+/Rd1SNx+W93imhDUZ13rNM4cpkIir55o+kzFCAQ99r0fH5GH
Hd0gCu7Jd8HLj1RClzrE1BxU4DyYPTudBpcPftpuD6BAbEjjvuBDNpVTZfE9W1kv
myJOoUpVGqGZhmu24YqpnNxSCU/jgHz+rzLvhoUuhvvrJM6SBX2gN73CmhAz2P1I
ssPq9erfpSDzSZ3bgbMwCEa15Jd2Z5c4hSeJHLHJLsLQrMptnUBDdrPlkCeka+mW
N/s9IbHsYWSQXBpP5CSvJChRhPsDUKEOYoHmplHIQkmPKhvs/hTID665qt9fD/hd
qaXU+pnGUdg9rPocdlIG8Wjo4uJ5RIKaVR49zu2cpt4k2JPE9Flu60kFNtrhYWuH
10QhCAxUoowp7caZYE0Y2FFifhh0VCCYR0hqEXUk9WcYN6szFoKJKF26vpxAj8Ma
0V6pSEOhEz52PYCULa7ijyeaAaPHuM6qgEFvD9JafbkEnKVKBdeSfvbTUZy42Ewc
OMv/pHkaEMEcsh57Zp3nVUi4+5fAKQGl1MLcFOlJ1rPqolytRPMD5cc34RULofcn
+mwUDncC+EqYPrdo9ZDXnyBg7H92QXgSKSw/QxcV5kqSaGi4P9fZiHqIkZShPpAc
HNMDWVGnnBQ3y1ZcgDTHn2rJZD/DN0rQLxI8u9X7yLvVFFjxY28WYWCAqjkZ8ifc
MCF7ykNKEqJeecRc/CxodcJ8PtMQQAsggwupMx9VXc6SYGFM7j5iyKohhCtewu6/
jGpWuGsTepfJBpYx16GcMqEnmTKYC0sY9eMF91bvij6Ux9ICxTdLT1YQZcM3auEE
vG/4bVc0tK9PNz9OD63aO6q3AQ+WiaqJu1tAc/pWFQHOBGJowpIGrI8b80GGXBRn
beLKFWENoOaUm5cMd9kVXStlZLSuyRYOoJ2QBuDtFYrMxNHWBSZV6GxNeO2gldmL
YX80lzBOWFJpjvoLZO0lxUYIOvg8c99b3LhxLwrWa286Hh2zCr7OnJlN1L0VcVRI
PHx3BL8X1AX/UcGT09RmULEzLbwlsTszGg8COIdf5Z8Am9GGawYfAIxdKnHvupp4
e/ksQZfbxg9VXXkDaY/aoG1ncBcOCi14safZJD1Sogc3i+0hkuN3R359wWawxqLK
z+L+Irdqb21jpPiNeZHgRqy5Ei0MUVml1HK6azFfkllmrxPYOZPm47x19mDcPJhc
7ngjBTvZQkJlwPidnM1a4FfFkKCnumGSYJ9vAepuMgmTXrScf3AwgKIo10CoQe2C
g6mWWkeAF/PnwFD24Ilrthrrlg4Jrg3rmhjHm14hQfzZGEDs242dTc0GirZj9iuZ
FaKMH5PR6XiYu8QMtCILZQ/2kUKs0QVfzITvosQycYVEPm+HzAuFQJpSpLmWp7ez
XEEAN3cgnuO6Sqn9/S5vtJ9SbhC3cHUJogR08shu8H/be97MiidtSOyyetgbdRMt
LAfu4S1jtzaBMC4q/jyYQgAIQEieYqIcnOXW1nxLoU/3QE/fjb7JFglzvSz3xFcf
s0BsrndBHvuz6f9Q34LJJbMv/XLKMgj0Kcv+UyttKs5nmMJs2i4njiC+K7YlgOMX
PO8igTh6g9kXwnI1gcMItFCF/uNTQrMGOUL6RKKYwEkRuG1EnI8iRv1OowGLvVkd
s5k2YjAcXzPSSEMgKpsBaNqWASKulLe1FeQZMXLwlBQMsssluwf2hR0O70B/br6z
EJDeT6c6qV/cTXPBipkQigehC9PyTIfdmZcp2MbW6WXYjMe1BF7I+JBrx36I4jXz
rmkL8NzMjSZHBz9654eEdXzBYIX66CI93xR/55xU0cT0+2rYwkGfdVHUgp+vJNdj
z/qGyu0RdIabbgI/7CW1gsQnBtb/hBQV3IZQtdQrlHbCBD/U38ctvyBbLhsrLdoy
ukQrORU9Yhj21hSn4KKWR0tCzb6hPXKpr2vSu5Kknk64r/P4eh3W2o7Rq++TD2HF
bIPjIlrpKPJPRiba8NxSgiYsHAAzR3HKveNSBl6ya8Jh6vHis+1maj86+Hu8r0SZ
qv5DO+TgzEoL44j0Pstq29VUUmMgFcXMg35mZAxoKN99Gt8fkbc4rdY6OZNa5+lx
+joTyfpfCmjQvlFtGDp8ECmBU3O0Pd66ppbKnq2Y/zWEc+lYK/qQos6rBMBDJMoI
BA28N5hmwfzS7X1vxZPQt3Grm6jPy7aNd9RPO0TzUqin446w3lpOnWGJTOH4gHpN
rnNQaiXsIlBaXvvGk5AARuYCqTqW16fnUI5XAr5cuidQy1pShuGyGmYDZ6qMp5PS
IQvFnUdiaTe/2dZaIS4+tOyWy9mi0PfWf++C2AseUhER1vOqkdp5SX3h5UYoMgty
pWwqJQvrrTIjCVocXFmeJ4hdnTm1a4VeGve1B99WkLF3Xpo4Aeb/pPNx8yDqct0K
gPmLSbW/ePhuk9UiyOgHUTJ6+FulNetigDwrjkZ5R9l2L5Q2M5E6hDErxwOzxCmD
2DkESxlB8YVlJAB0P1HVQ2hJeQH4iWqykDP+VqQ3tdlAxCbWGM75i1lpE5GgpwnW
tR20YI/jZ21CVz9mdevych9Uv6p8VRI7HkZK5yfue2dEefv3nYxv2k6EP9p9FF3X
vk6VFY0PkoarlaJIwjPFu4Rhey0oT27pCJ1pppv577EsMX59Fwlrh+DWQdMJgKk/
6KQVA5K5S1mWqyXMRHoHy0ekoOr/maCqkN3nU5RIf4ivmeSKX6rsbHmZS1LO+L4P
HE4uwDjr9ymqvLLrnHutychrcLPUCugvzpqBb9jSTRFHYmBnZiLMTDIUdd/l6Q4E
HXeE3s8CyLQKQ4fatoJ7U/YrrN+Id9CKyKDxfGRIwuODz2dnrufnVUIIfOm4Bk+0
BJNcLMMqi5rYMMsep5th1Z0/fqs7zSjGLQPn3YYYLE5cwFVbe0wgj2kLCMsT29l6
YDPtG5Nxvb5hbEphb/hZ4Meu4//wgeJrSR6ec+5vt5/yIIids7dDGp6nB9K0M/TD
7TYsJdqY4xa3JQx85HiY0lO/IOPzPl1Ubj78KX1X5a2SoPCap9Z1A3DRaQq/FXRX
5JUQuMqls2Idx642kmIkJR5kyCEfvu43cXKalK2tnZc1OyLHwqbCZEjdUMR0BopX
dySojOtPlnfcScmw+jZDHptD4ZFw8kqRHNrlYsCk9D6Ts1XIInP9RC13R3JPdwBO
PcjMmmSIdE3z9xp5TYK7b0lXSQ3JAegPqkaY0TWR6IkYsSEOMcw/f8Ew4beGjy3S
P17duRuwijA1jsqHebsuiDp7mr52kpTk1oF1Kdr/gNay25tGa1w9uBuhx7dIzoJB
TlwaD2MvAmBoORas4P0DEC2PiZl54kYJauyV5q4DCdthMU1w4ROyXhHFok2p4nFf
SrHbNRUhQ2jyTYjVpZuHW2D1w7rpdgXn9cEkWtuJDnfUhZQK2jbAYMSQe/8i7xsX
LtdF6Ec5qQBs/Fzbgy5biUAez8CpNpnA3FYNZpBHHTcNSr5t70cnPL7qL2o/EdoQ
AyuzDrQgGl1DgKaW29AEvOOs0PPWCF8aaTEyGlzCe02lofLWF6o3mlZ4ManG6cg+
Hek2NW4p5s52JaSI7D0xcUWdKiWVbhzJfpSjK/GPT1vbXltzk8MdoaD/MEFhMBSo
t19Kg/uaqBGWtlsywxfX3D+k40dBA9Z0gBZH+tuiUGq6WBcP08/ufNPGd7+OGXon
O4RBrcBfdg0gJjdaZKuuF3WiPR12Ofs7f5me3uI6XA81xMib/rIzvv7e4SWuzvcO
jjRDsffZd8oD/MuN73Ot/zR5WzEubg4T+pm9w7kD07W7oagOYcUJxoThJ7dh6JrC
S70o7hgWDX+rDiZg6jCgeunlNY2fdVQwAbgzwH50TOzPZrYo+3sonX/CC+5vw9FV
JPmVflTiTNBq9guELlgs+XEaB6zi3oohTQ57KmZP3aBtBPPvQQz7+be0l/JNn615
jzji+iOWrEh7C+bFAqiScSX2NpcN/Gtd7bm7PHWo3SvqQ6EAuAipIaPcavRhnNMC
1ey7AJWBxeRxktz5s7h4zwXRWJDJt5kmhqMjYrPdtM61iWGFLQwABtcUZn6uk+l7
T5mK2/85ERSjmIMIC3olNpmxUFxJ7ZnLtPmBGTSs6o6AEcHoz/3piJLxy6rsokbJ
UJihadM8x1leypm5fU0RLKzOuLaE/RmuI2GTh7P9uZyfhqvjf6a5cJd4yoXK1Pwx
KDU4YLP7Lp2w+UvYydCiWru3S8/WbIIiLDwfp1SN0jK2BpkbpnkTE/Wwym3FxnYj
BO4qRsW0ZkD46p28qwJpbPC3Si0ikQOpBSSoDFNxjHJwzR9eM22xD8pKKHJabrUV
D0FTgydf1A1d97E2rLk+1ppXCfaS6XzPFP67OSVecHuppXX12m9xdDJAAzLMFNDM
4NBHovXvqTJYr2Cj/8ef6RSc4wqBTcfemd7DvrhrYWMlisrpCnAJIcU5yuMP9VvW
aUxmd5WefKieGfndbMF04NQ+Ak6TPen45fBXwmlCF9BcRRN5OYUCcCXcYq1567eU
ME8MJCFbgr7AI668ZLh/Q+/j88S6IqO9j1dbIfqtGePFdvwi0cpnyLY4XU2WGaMj
ybbHk9DcKs9BxK3vCmbmvvTO73regoqYZORFj7UNUvwXmTpZoYzIE83gJoRxdtbS
lcMU48aQDX1gP+Qr1twaLMBZ9IZ0tXV0n4E66V/3B4sH3ivfFrCg5iUyajsWHzwm
Jkrfwz/m6JzSH+/3u6sTNJtWTAB90Vyk8ygoRTVOaeAKxoEb7bpqa8tJfBOJo0zl
01GgA8ZpUxp4sqLwLvF0c2zBlZBikWotBCeTvP0SYpmrrnoQRaHR+3T04KwOyxJb
LPsdzhU3LoIrd15yb/NzvMavbD8JTYJ6O4Zp4Zjto27iqbcwBzLgnepXWaIlesRY
3jMI24lJskQC6F28stEFGjAeWd5oKmTqC0iyAhRWLCUpgzcCaJJSWdtpAqxgfiOB
zBqna+sTKSkTf44JOhfq3ieV5K+sW8Q0B6Hsm/amG0lNJOf/NZIJ0zCYh33ZwDLw
ATBT25N7iI++0XKVVRs2tXM/sEf8vT3Z3Sel4e3IiWCpnXactOCKD13/IKYKfXgO
wnWfrmAnC0uwYXHkYkYE0V1c0yXTLnqiSqXR+QUU8e3jc9NtwlWxrf8FoNOyEK3W
rUUH3+EUkwLCVILyy8MNcVXiyXoqX+0/2xsWZ7BnCreSuaNXeOR2EcEJTu3Os+sP
Y7TovlVXFMg4+GJI46pOOZn4UuR/kMc1yIBSPsbKE51Oron9EPSTjDnKyDwfbpJY
l2pkOzmv0qFUge5ipnOG7he9MGFpOv3kVL9W7hYbw/OuFLSsik8YgNYRnBmN8tWe
gRCKEoIr9uXSJLbqXNV54MsSYfEEfbyGlTJ4vB7+q6rViBEMzAHiihKtIa9xztfO
H2bJq20wAx+Q39GucOuDyPt4t2Qxiyr8HzCfDR2MUj+Vw9lvxSijC53WblrylNpB
NHQwAP44cXXtmx6IcbQY8QSNIDB0VnxVDYCSkBsSa05eA8y/cbhH/DaXpBshCFBJ
s0GvWVnib+mEY9Jt0lJvlokXtN3arhdqbi8vDPoc4pUkNV94jq4ALJpdgsKJD4zK
kScqYCh4U4j2K4V5M4MD0WFyMsyqY7NQQKDrAxd1fvUg1tVHlksPKJWMAkr+zDy6
/sLISmp0CQFUhwHy9kOAFBcChcaUp7ra2sv/F7rrJrRvscy/VQg7OX2vixdXiYnx
jM6a41biQdvFdryYMI0JmS9YwlRKZI9N+28sPG8K4D8ilf/K8zaWktT+XfUf6bfl
RC0Tbj/z/fhf/sjzoDezMrRBkMxBIMWvTMH9uGYX+ldBKBzz7lTSowcnE0C6L7no
EQc68EEz2cov+4HysO4PgIVjc8HOkqZrjUyjnehxT9MWbnNCZEQ3wTQo+3bQzoiA
9Q8uGz8k3VxCGh+FkI9/+uysVTDQAzCGyACQjLzAFaX4zABruKjRAL8GDe6Cn4Pp
jb+xi+RYXOWA3idXo9gegJ54UG61f/s2vZ726DZ61Vgkz3IhIxg9TjS8c9yDE6ah
TNIY8Fw5IEchy/ri7HGcyGdY/tPVrQ2I6wPiRDQRsKN+TS9udyIKmsyoSMOpdelq
yMJzARsByQvNn28dxbdEa0qcnEn+gVCzhl8LVG6RaidKkePEbEQUG6bV8fxQIODa
hAp/aWt2pd+CN5SPBL9Y58lUE9HA0OLsAeIIwxUqLjuUFkWURUylBcsj+7nzGmQf
KhYCj0Wsu1fGny4fwgAIs/h+Ymo1sN0+kDadIOZ8XPLmuBI6XNfz1Wv0BqgLzZ2a
B9tC4js8SroLgxrAa76JrOAyf04dObV6U3Ppi2Y4RZzR9+jR9foWhxSEI8L1pwy1
GEm3LsZmoHo8kHmoWGBa/qbc5C4xcJ5SRBf65jw7OgDh98l1n/HOd6p1Af4xF8aC
qukDmQiaWKq0E4d7u32qc756HrNk2hnBzQJB34WBqVXjfzbv9FREnbSEY/oFe0bE
YoVvHc+kfrExPXShk+TMgVy/bDhe6N7+jmYafw88v05E1IEf/13pzQ3EzZO5lksf
M4MZOHZa9hm0/ZfhmHkMWQfwIMp0odYfDF0HeTgl89rVtAQKr3n5Bdz9CpsM+ULQ
N+42WdfOfdS/P4x//n/Irf+atbTNCbtGGYXR0BzhO13es0ccIkocQ3klGhn85iV7
tzNZjlpz5AgHnmtVPlZNUppUU7Gvzb42dbiFl/j1UPDgs61j8MBbwRq4wrHesBNo
IVSRqUdvPszgpDz1Y9WOCVaC1lGC4g0k/RlW9UmYWRUbmCGCixvYD+0O+rwM/YJe
olXZFm3ZipC0c2yuAwEoDKQ3LXUkp6sXPg/p7FGBuIUANQXSUNGq0OrNqmkYn6Hh
Uh1vHUS6Kg+h0zrOUF6j17ioJ1wY6XirJHmyzFIbcgbwWpV9SU5EyUYghKLkFpDl
a1zrWcr5TzlEsVPUylJohcBH9nZcZtO2nD+rbuFSpntLqaPFI5ogW204a08rPsvk
YP9VAZoGCAY1VzH5wzh95KfV/87/tmth/akXG5KEmn8u/vp1r78PhrlaRAHhT9aA
NuZFgtpyNGvL51gAW1MdEBlPA64AlQni24SwkX6BgvG4RwtXiAETFvvcXfktH+Cv
EP4GXV4YmhNGa5DnuZGehQI/T34G6E/bo1uuJvZb/R+K/nFM0B12OWJIL1kjlvya
kIxELZmEVmk4obvCS69EToNQsEZ6i2D2ALf5Qr9eGkL4PMvH5/8D8ugZ47/G1hnP
CH1dBoQfh+0wF9w2ltCZulQ873CaS+1zyFI9cAtxxyaqyyIya5mmFzotrC5AWr9l
Ahd+XpvZ8lTurACtfsJ0M9KJ4oEwD4zmGFOzoPt0X6BF8/RENFX8Y1GprRG8/naJ
Ttcr29lpVmZ1Qct+h0btj6VzvhQk/vPFoj0OQco+4das3eGP9rj1fZIOrwjgjdCr
jiqWNzefyllF3mNlWApGmvk8gSV47/NfsKbHSrr3IdzlZIqqhcxenuGg7SHgMLnu
jCKvNc4blzF89dEJzsZXm6ECykHcfaoIb5FyFcBDvRF2/7BD1e94JXr1cWL/A0/Q
4DIzjmyGPn4UsXgIoqy4vHv17srAybgklb8N/+ew04zXjpXsHzGtx5f55tfwzNbK
WxqpHmpuG/+bx3/4Uiwdno5Hd9bqy91jpl6UHnLA/OAV7L9+BOiCk7hvNvGHRVBp
z4NW8/uakKrjvIrfNNj6yrVzuY4mytBsRPK/EmaXD3jgP36aCD9bzlIsApp0seDJ
a/j6gUiO/z18G6moumDtw227WfrUC027M01m1be5LdKTFO2N4EqrDXYhcGM8Ekmg
efl8WfvT/0IttExP6QblhXb52WbALdh/ypkLtrUOHWwkZ5zl92M753KK82UsdAQr
OdxNL0c1zWmxntaa44nreIq2jlC9T4KXuoUQlsSmDXDV3Nq8OnMlV+AznzhMyg6S
qJJGIh11A7x6K2I9DNOwlXTjVJo4ScM+8OSAeLIRYTHoSoGzbV4FnbovwELYwS2G
BVnqEPq+fcd+59hFLuT/h0PxcvGDhN9ayT141Gb1cekFxVC0ggkKgwdotz4+GCwV
kWYNemTU1vSArvu18cczPoybAdnplERxwM2Vpp9knuXU3D0V3pBoBd4GnkzjVuW5
1AFBKHV93iwzQEuLvNqm88F0h0Lt+3XsCtb9Xt9I4F6l6a5GOEeKodH0DHSpczrG
pTZ33IZVv3DwPwgflmGq01h/oE92cWxUrDKZaVc3C7y1qC8QV9RjL+r/O6e/Uveq
UXzKdboZUqTpaG+SIAYRIhAJuc/WIHu3vvzfds9q+BByRXBNX0TFXg3mEkN17bhh
Dhj75/v+MW3s0SziRGS/dtLe1dRSwwuFjpXKWZI0McnwbDrnWBoU2dEHt60AE7bp
urwc9GLiFi22euZzZ/jxNOcdhn8Df0mIqyqwHazqpmYiqWMKzQqhOOn5aaZsApZP
D/hE6Rxcnl0Kg1O8v6uhEgjbTG6MOX+AnrwFgl63YYhcYUgueH+rcyosZoNtBfdN
6Kcj3Nb32lqcXDftg1KGGpPAjXK14Y617nG/SXRRdTuSiNNoF129Tld9WpIfiCXN
OMFTpA16zy5ZT2gL4B8GA2dlUwLbEUwfgdYqu+NBzhu17T9EjXG+q42/u96MntjC
N0ZKZ6L2q5qw2x3RByjDpfgcmPGFk9jkyuPOf8R1PlyPPbnX6jJ5orV2mH2HiTIG
QbYfi4UHtHtkCU3N7lJ8mo9VvU2oaMVzPM06hN5Gnpisn/ykwZzw0ntImB/3/K+0
QHcRyFaqDWIf82M6qDdUlKgtRBAI3UYTabhswS/TcQ7aUb4Wd0cX/Ey5Th3PaCte
G1ZW0nMIVyxu/+8omBPtumZT7m0GTHim91hG788vAoSZoM3APqr5pe0RdK2+7LLv
aG79LbqitpNRezr1MLOyIlERPdfj5YvFupLtanFyB89sQZ8SCRYxEdGveHA96OPj
1n62RJvckLSYalzG0p4PKcqshr/ntUhvWRcS2w5TiKTOC2c60FzhoJikyu2xdfAg
yWikZHsCcJ873kwhtQM0BsvtDI0BcMOkY2pJSGDl2D11jnKl6+ojVXm/Ww8qOlPA
TvU4TouICyoo8ddcFSH9BFVpKvTd7hzzNStEhiAFNZgy5cFc5dp+41M+vGpgh25z
DmGre6vy7Z5J9ZZ4s+GHaOtyiSZJSSmpQHLXO+L5djz+NmIdmBTB72SbNdj8X2bc
7zNj2Y84WLS6S8iYCHK6p28q4AGAfqb7KkYxyd7kK0yg264TMQxNTHYDgQc5AgwN
sBnaK7XnLQVtDZ23bsTgQPHa0pvn6bYst2LMy9yReg3Eea173Nna2yMtkJQX3sQY
9IOJeqezqhCoRPsN67LapmUEzLWo8UihWfbS+224vogw8KsnDx4w9iok4hAR1nMG
Z/RPc05vLGKmwRVSCRKjv5ZyixSxfXefwYHJa8iVgOG9+6fzHnOSq+kd4U7odJlx
Evf1UVKHHu+dWpNupTNVkE6NFY9/ee/zl79G75uIAqzjV5T1RpfxN1KWiq1Jn67J
OsHMuroJvsN5/8u/V/Ax6aseYeOGDLAxP7TTwJHci8MqMgYN64AuNnCZgPTT+Ryw
i6eekymVUlCp1gCGHcpSgQmhPpjxOyexV9yG+JGBIM5yMOs8SkXocS/eE5v8IQWR
OOUZ+GfCixsXNC8h1MlT+wvLN0/9H29OL973fxn9XJxfsGGrUbWlyY1yRrdGHzUs
+SuI9qTpnKNBgS2UIuTUjZBQn9EytU22wHcy0cj6BgseZxJbfZauNj1tQog6r7sB
Sed/sJ+HDlS93qHWcUDHuUSA/l8DMQ3pviQCKJaaVCUBtw9JVmqUCzf96TGOG0DH
GRNDWGy4jmZ8sqlioJeMtHmMd5Vg07G3zs1puARjr2HbpvksvkGomlD2tgDGc+Yq
Vw0rK8Cq8oZGL25ax8xrE9rM0xawIh05cz2enW4rI2YfvMN5/qqDYOM82YHxOHE6
L2BzE3b4263b94jiIsVY1qLuzlXNAHcDCDvS4JbBV99ouo8i6wI1MUp4VaqUaJPA
jJd2nJ+ts3h5qzsrv0vGGNIDt5AbpADGObfolQdxY26n1C9yhOufwQjo94Zv+Wn8
vxfmqXGinKI4Ebsq3xHFJt7BGN9PeK3vzd5RcN8LPwlBfzwUpMzVBSmoDSOS4HHf
TpcQamsvH/WSr3RlHC62oOx8vZcpx+PyMw9pseD1qpKdoCOq5TiaJNCN4yInYFbg
s0Hf0Qvvf+fwre5N8tr3Y8RlnvKpwBrdAwZNyuADhrjdi8jnY2KDZtoHU/05eeqI
DLvBQvarBewrCOu57rKcfVSEiCF5mZRNJa5fN/4G6BQXwxwpnNBTLcI0Azcpiccb
jbnQg0XUT18+27nWk+DxcNlTYeZjFdz0v69JlM9esY4SwUwAFyrpKYIz2Wqm0j3L
VwMPddvnfTIa4vxc2nBAs0bIUVjGoH0Yw4F5/ziQS5HowYsongUz/Tmkdypy0DoO
z5m7KpJfeTLm1s8ux7tTogEcRpH7fva0hNiRIxiftjuMzTDcZIhulpYHRSo4GV35
dG2veIUxN3ysGxbUC99vz/boL5xXk2A2hULuclUkyJ2ODnxB5KLzAOS5Y8iYR4ze
qPfsOCAerHPo5LvlGOdQbs32drTxM7lnwG9D7zG8Z3YOdnKAoaWApp2OEMqimoTF
FIdRk5MvZJadmt6W6x9gnedYGQ/e2tY9Ccv9/F0K06P3hNb5AwQ9rieVcajhivaE
vLaj9nKIJ7eogTMTKzlH/TaSHkU1AyR+I+CbC0qWyj5p1Dkap8FLEyHzRBlELj77
TZgvucEkp4/zj44xbz0LToqDUiUWWtGWIS/M1N8WiTSJJ2mdRnKRY34kjpwJ0EG6
VrXXb2JPHtatvpi1qtcMQJNRUJ/owqXrjOIemEpvQhSAzJtY2zyltdb0jSBx3Njz
SlYQDGXSexX6QXARkFI9BmqN5En6NSDZiIASVI3V/18wYC5r+ibKuxm/LTN+Pecz
scvwXft6Wty+9WXNRSnf5JIvc6pPUiFkj/Li8RiGmn3jZI8H9qrSwn0kPTYClqW+
64ntRgLnZLugTPj2GJvFvsz3ifoSJdTi5wLjsysiIJ2wp1g1keeK6hY2Gf9ljJrV
aSnVz83ionLU/yJsuB2T5GTirEnNpWEoCrAkFUl1avWcfASBa3+iNrRXO/+3PJ5J
tZeJCnANtnf7m9qBSthUPEhA4+ni40i1Waxta0riZIqBnt374WRg6EYCcnAVXH9a
TTrzK0oLKY59ubPe3vJhe1AmvvBFO1ICHw6nb7+BaLX1UWcqxfXTttPr2zkT8A7c
WSML7AYpK1ovf7lSG/NCy4Eq+ltkFwUzX7/9STSsQ4SwWYqSbyPpTJbihkjHIKlA
SQZr5EdDFfMFqLp9CgKkmHIPjEZyFEchvIx7UM6GJR+ALgHDPLJn90R3EklFgpz7
PxOelhQOS2RgxlsD/FvRiy438+bRsOP5FxKgv3xTTswkP+Jjg3lLJybaai9Uuk93
sYK2uIpZ2XDeSwmSmreCCiX7lDXe7OeUz1jw+A+GtMww3dFAQZ+iDzdxyVJw0hxY
k4fFiIw6jn//V2cuSqZ04mPAiKW3wMhx6nZG4aZfGJmoCB6zKCDDpO0uD4jHa4xg
gbpl6/CFZG3+LY11OGZ1Zly/bI/26hPsUGr0DciGIyZTy/4JZQTyZnpdSYJicolB
maCi9A9o7VwHUP5h3oRtORbXq0zLZNY0+T5DtGi/woLyWgKA4jDcyRaeltZj6eym
TpccyKooItxfIdaoUm89eZvgRaV3o+HwXsXsOkdLeBM1rzYlZU5bZy3wX+AS5i9o
4Q60clOfeDshYd1GAIJy6n5a+NnK/euFWUs/SGYKtPA9aS63UM9QtgxxFKNcn90E
tDpco52g2mtWz6s/B8NvU9vA+RPY8XIE73Odp+yRUSoDjtb+kJ9ONAUUQXFSxKLZ
VC2VBuI9vRlA0YMBCGgL61Z4OWpd8JmQbQlOz1htw7LSeZqoxC0nyH1duezaGBW2
I9A0eGfnmlsZUBFyfbhOuClgPGH8XCvvrX+WhHl+ptp1dalAd/UVIjhzPf5o74YU
BnJPEvGYG0MJ6T/0VMIo2jH0gWKAq27lMqD9y3gcLaM61aB5jB9Wl4bF1JTf5/TG
9NyoIykGpVAn03mNqFXFYpv/G0mPSqAos9oizxlCAQlFadbzI4PpIjd24dOkzPBg
Q3jC/zr/sVUiF6G+ZkJNSfvROWAacrPogyfSnWqenTW5Gqh0NLScteVF3HDw2d6b
c7qmp8SDQxkv54PhT1tipr6ef6PmIS5rxDnV4CFU3AmlehUKQQpdGQY+r4Yi5udA
D6NH/rV++7o+Kp5GK0iQEovSwS5ghg7TMP708cFiSrumIUVBZn7FD1hwoHKg0V9Y
uej8vPCAptytI9r7cyFB9V+QD/2kl2fYQTvYPtG/NcK4uIq+5vw+SCki2jYvswbP
Yli+STj72DXDLgHigvw+17R8e/hOKFEkwm2v7k2O4/43pvG1bhxsn8zapWkRcHZt
Co9qgLa/+xGYWji4E1N9aF10YcycPcr3Th1cWHCLOhD1TCwGR4WXKHlLPKHiSyAF
dSO8fYTPzNmM1hmY/0yc45zLnUnxpbTgpWgxO0uIeUFYEAeZJgsjaqU+QZWfJ2Kg
vScgHuMuXrcRErB40TCkpaGoFrlZJ0Rh0Jz0yZpilCt58N8IPa561Avy0Y3m0+tM
km0/EG6tAVnMhddbtmZCOTzG1zy51NvdcHVXz8R9HcfMrqyvZZS7FXciobFNpp5D
xp9ES5Q1Sk5IVyOTFIuKte+cslMc3S+y1DKzEJ3b/b4gdHmC0YPaiapwDUkJrBxc
j+Mr4uYDHsNuR9lZBCSje/gtq1BtsQo5SuayMKRfLfVlFO8USHG3bVvYjbySFRgp
JC0mcwpZmlAwhKHA/dssjfeo+N5s3O684yQTO60+WxA5T+qOYdyLTOnTG0cO3o2p
9SPBPXtb7k2GCNfVHWitlKZ8gb6fEJ1TIO5EUpX8oxIv5V9rXURiVvNKKiwB4tLa
+K39rSXZQn+69OyJl8k+yvuPx7JxxyYbFEA6RZGTqHDrv+cYBjYulkUsRSCKlIZy
SDmHTA175EFO76fvjYLjPfLQerDZ6oaWKlnBzZ+1LLHugYl5JjitQZXcFtW0sHP/
1z6tQeRo6elSIjJ0q+fPiCI/AYBXINSYPfvuq41t51MvxPmVBLRflRBK6CIxrsdY
4Xyc4GcpfqfzJhinFA27Xr1G6jaqHakmxZULP5i6Adm6hP1YsT44X2EXDL5izGDI
zuw0WMIczDbr0tEbw3YFwTpLPuGsZtadHxbti4Cn9TIMgqk0CytdTAiuZPPdTR0U
2xApxe9P0dWypZgoPMEkh3NuDcqPeZis6wRWIjZA8etFqRXNhtlnMMzlbDJ6mQl7
QtXaInd6kKB2w0JYv7g8ajr8Xjh8CunoiyWX01juyw0A977O52VmEvPmIakEwUrS
kEwKg7oK/8mdV8BPghEZa9SZTBr+NB2v0an+8pcl333M9HqI9xSGXWhufOJKdrYA
SiA8ktnQvWIFY315zdgaVsY/cl6jNLaoO2aqOTIF5FdrvPaQtq2lfPeXq4lOo+Xn
JtWW4p+EI0gZ+m6Y3M4/XonuV3jvLNxL3W5R5xQbYSqWl/rTBFAsyJBMTPpeX1kP
dBUrUlBBP+MQQT5UVUfT4U1/iS2X48TBL1v1y/BAvv61sQLNC96p8/IapQRhLrxW
j3r4WEU/Za2RQeWbW4LIK5s9B46GuO36JHsXXuXy7jwZHhKZI0MPRHs/Y9AOWZ5z
yHwkRwH0g13QPfXcp8lKBLFCn/s3Ed+/ibu9hdxfGTC9A37ZK9Oo+8M+fdMydLhT
i3mN7ci65uzG2jKiciY1juY8tx+y8pRIcmppS4zF3mAFELRKWUQzKTJ5PH9WsZFG
R0Atx07Fle0ptJQeP5O4KaguqE14xRxo8oAB3mopiuGPCvgVYCCcRxzyuk+HZr3r
g9mYztNMgeKu/zWsU7GNjGFqbKvfn3uU20hnmDIzdTfsAIn1hXQQUxpgoaAdb+3z
fQh7nNaHuRnN1cb8d/+isMbTil5srHXKwLyxx8VPP5Yqk735njxpwvtc86RK0xLW
MMKa1uaX9NfnK2X7Q9vKtXp9IPRi31QuG+eSncEq7lh/gwe4kJ/yzGBbg4YlKPeN
hLKoNF92ggfKA8OnQKEGOSFQbvOcUT5Mz7QcIzQ5FEydUNkHCDssv6H8+NLHGdTh
FflrqZSCNj6HBoaDTLhOoqxgg49G2NJ05CN7VG0zaKj5nS8b1JPbChzvHOsUzYa2
sxiRt2kBgajx7KFtnKsn+GHnpbfZ9zVakzTJ5GnkYdeUs/aw2u7PHxEojRZcwtJI
+SHBFpdRSx8nxjqU10mM5Ei1qgAJWoypKQaQbfycMD3ruTBu9kwXpuqoNizsPuAL
aB7IdfAK0n5hnB9l6u/Ms1HvE0+wU+W4Zxi/J/qrvjM+8nCWnWtar497i6q7w0A7
76va8/5AkOIHOiNX/I5kHpqKXZiwHNAn0artFzDlO0yd9LcYWhc7O4HDaA+Vlj0z
uST2GPRJCvjlvLVlw8UL8vGnhSkSEedydjNZB+5+p4eWwrUCybFYrn1dKnuhtcTL
+15EZqF30SH4F0T4/LCAdP6HowkuZmiOoSngqo3nCYWG4neMOjFaM0JOQBg12ycR
LWew6HzGMizmGlS57NC1/hUVh2l0GLKrmtiqSJxJi1XGoXiBmOSXwfqoPaGKOzPJ
4VANVFZprBNTUKJ51lwYgoJU1kMoyOD/C3FCW71iPwllxFccTcxpnTXl29HSi5e2
hOQVltdDQah0ebtt5DPcRlfqyyL34ed/pi56PuC71uun3PrubnK0MrqKscyK8uE3
xLc4k2kLKv1wdfS6FsMZsID+CtkWuVnhNN03O9vSYJIqamxyCd/qisr/yppvjFFf
AK76hPuBXYKHAj3uxsbZ0Jwqj+Hc1WFsvuGnqulkLB4agNM5KJlM9EA1S/nxi/Dr
JDOIKWewslxox94uXj21+MiTdoPR0VX95gn5UEpoyfSZAo2XgOMll7eg3hyjVCJ3
9bFUGX5la8+N5mipYP4USOzDTv6Sk6pexFMuylUiSll+SjIzFoDPLTNndYVZA0+d
ACwTCqTKJnkSpvVCWkBOEbLDCiOxqQ0h6Imo53U5zlG9U4a3xVSDYG2Lviq07JKa
b/Bh4/YldBeZKelKuRtSWiSFYJ1DptBPhSZfZLBpaVGYhwn3A8pJIg2+pFQE88gK
kv1soKNIIN/ZtrCfr0wGsOMkWqImNNv8x84B6lSdjabn/f2GZ2XSNiNgGkBxbzNN
0+2HqDSOhhMTnhx/76fCQmd5TfTGNARFoy/YEmOmkC6ZhIaNu4qZqzObkXGIG+ZK
3Oz0JyGXJFuOj9MHtCP8iqC89Abwi3OGmNp9CF2SAUpZNlJEqJNO8+Khx7LS/hlt
oSFrF3JiSgVHsJzGseNLl6g2jG9a8m4Jx4rfTo5uhgMQGDAzupmODV18ejN7UqPF
ZAUB4t44EA/a7r6iDHu9o5RKec3syMSa/4AtjwHfssP9LXlZxdDFz2FB7lLTai6R
AUYkRrEVMHkG55VI2A+o/mhDZSouZNguSBy73Bl8lo12jQzxA+O/NcSywY99tM3x
vl9G22PkCjy62oQOBH0e/C5Es317iO5K3gGtJjR5Xd714endHVWmvQHesVuDC0vL
yIPJm8CBeAY1OHf81WeQruH3v60xgUNKVwnn6w3jWkzLsTenU7Dd+4WUzI3ek1oV
URLIPBfYdQ0dBc4ZjD3yLKzbB1K9RLmhGz3S4hxeJkaDcWE0QKa5dySPEO0cYEwl
uVpiLvwOZgFfjom9eK+R0e7rbcTLAevDj8qRUaODPOPcIdU+iZG0KYcpPNoQ+ZIz
VLUnQpBDKsAExZUYtq7j2jEtBqbB+U5M9p1B/iuuj9wP5kR9otXbK5R7k0UE+kSd
6IoWQl6Gy2OKZb8gW/IGKYc8WJDs39UQlxomcR5l9ThNS03cS6y1t9+ZObyu0rVg
VDLjlkj3W8/OcroYRNHvOmwxHHDaiEa1EuzT7V8JSVvVOOR9frKDJN0FjTXFAZVy
JP/KZGLGNA8w/mpg7KPpc9Gb2k2lcyp5nAfJZHuZU34pJCNE0j8Qw8XUtiFWJYt5
8hZyI1M4PzKMD72NRYWVe3XL++OjE0V6L84a+2I8816c5G0G5/A0/TEqGIxJnXCN
sZmwNjGbM3O1nJk9lL3RLGA7U8J4lJZL+4WycoepCjOd4crCFwvOprBk7fgVu6xs
mrvZSuEuidKXtJtDg4DDJ0anFBBh93Jw62sFGbe8BOWwpg/mASaCVTmdG9vOXpdV
ZVvNTgDjsXFB7YOJgdjsMFhFQBt9n/VC6nr9ArOk2Mlsot0cfXyW/UDs48b8GvsL
YeDwv+ZicLzbwS/48yjPCSWbnMxPIaxVIUYt3Gth8EjTJJh8d7ozCJX5D56BJ6+7
E73kQra+iG/vV6MF+Q+Rz8eL+btYlHyDhUD9TjcLPrPuwWWxCk4ySXFDYcEP+bn+
RWTXAZumXuaK5Q2d/eOSCUew4wczUPIAdTcvBG/vICchrcUrCNH23z3CuTR5cwJK
dtBpy2RHIA5kS0LjtgwSIx9bz5vyR4GE6LXxDHQzLyaAX9RZysqDh3+cIsTv4vC2
B+NN7gkM9xR6FHEUKkHoNMzS3of7IKF+Xs0VZUxttKYAYwQXy8qcyj2sCs98+DEQ
Rv+yYtCw4Pjdp10qy9nzCjO8KwfFfvquAsKh5xtc7se1u77abNpdOrVPobe589Rs
2MsvW19fKAp11Qz+bVG1noT7IQ+PVUaxWtcerOyxA4KqmjqJm7gYXspOLiVjYx9m
MjyqXCULGl0hxEUNPIrhrrOGfrzEb0nQNER4xPKTAOFKa4P05k9C7UKPD3jOzehX
OojAowHWyZgGbQFOrHos9G+LnoKtXad9/4Gje2klWWTUolSIuljatGRG+SXhkh02
sgFBTV5vuYqiTAhJskQ99ylUNJWlFwB1+QETrWz7XDOyYwesPa6Ie7GbUwbJYckX
HjCp9w53+n+WjFBNaHpNaurnwKJ6whcAUAryLuMZPRKI5GyccgJ+kXyDjjwHQ1Vg
FYP9nNkU+dmphNU6hopRfmWi+4fBhjZnMMdEJwDhzJKypMspCa7VqxgPBP3IL3QZ
TKcjL3+n7BqM3CAyp35wctiKOMkH15+7fYiPfQ38mbzxTtVu4/JGA2X+YysNt9rJ
H92A4dsDN7cTC6ygKi8/fy+NU9vJrXe8+fwrdszzozJXH1zNe8hrQuO4x7OAmE+8
ih9gzhwR7jEu2CJDeqNNZckOArjR88zKdVmhKwXTQaAvrjtbc2smlA5m1+C1S+7R
ahZrRtLWv9hvpJtS2IZDNSAC4IodeZgP47dGdQ2EkpPjYbV5hZFzEuxeRkbafvPu
7coJBkorYFETw6Hohcn+T8MAps39iUOI0qFHKCIeGcqN7ZtK4BrmWWCFurpJW7R+
BSadihT0IRn/7KZYORfx9Ad5+nqF6CSiwCzSm8yd2vlL38KQjHW8curJsPWM7n5+
apXLNFsIbcX8CG6YafuXmVhs0j6gEwZK7mNg+vp93uKTdOPmd1JKwwwGPyqhTacx
tlSJ//K72+T9AaaQ/HYvosAsGHxJylaVtFskPEaUqwBoBumyJlS+GKSzxCli/YTr
tQIz8EumKd8HZOUnVI/MntBfDQHD9DTtXNixolTCaQYbo4+rZwq9NTmKJKFhn1NW
eFrRxkIDZmESCHfcjjwdQMvrFjUoFpmRrvpj/gj4xA30zUEfMmHdGn6md3E1hYrU
9V63HsDEVDt0t+FhAqQF2qfjBNbetV9XxFvjlOfE6Qy+AktUILuBJFWi4wEv70/V
VZ928D3qZmaljG7hrAo3IbDaRsolnsx3bWjdWavzUJIeHQeSczJjcsfJqxR/unIG
20zh9cq/+YlbVDHtbAhbW14Lul2knuCSh76IAskZ/Cb+HPd7TRhWGlhYU2EaAx2l
+BvUqcEC2giiYV7OgJ4eaI6rppY+S9Dr98Hr7zi0v8ojWgtvWUhRbuvqSigpuu88
Piqxn5hOo1QYqm+wMAq1Q5mgAXPHBVwVgwIe6P+co/XkDL/znPBAh34jpYof60OK
Lr3rKG/ETCxQtKZhVLfrpgRVqYvEV80iEuQ636bf01X7QviivyilcE9sLdYVp3u9
5wMf/my/kRwqaQ0sT3QkOr5uGODo1y6tLwpytekQrx8V6CWrNaIYujWhZ31dwk5c
ybGj9is+a9z+YGcC1EQ3EDrF/FbxFQXIyl8seBdP9I5HUPisqBC2yTTBiaZ7C5ol
IbfWWHe1k+HA7nqO+7fXRLr9Cxrxj9X6+rB3tLhwE9bxfsq2q2ET+BkO6u9W+TZE
MrhSKMPdIbGE41t91rskPYAmD0HZhkz8+S+eYB5cYVTm5QocgWSGvoqWk4JP6XD7
L7jKyfdXjI8qds1pMDjHWX9HcYWyFJGDavgD8DdWK0G9HO9vjzMYTz0JVuBW059T
v81fKqzpU6Os73F2xcXaZThPeSdnlSpxYzkTCB3SbEMD9zOlBz7Sm97ky6oLuEbA
tIobnbe5z/O2sxPPwccoW+cMYsRsrzXGuFry56r3mcaZAeuKDzHGUvLWkBMWmtD8
nkXGEeoxp85qDAuLYtZqlLctc2//vfeKY3pOPavrGObiPiSc2j7T3kVP1V70lsnh
pUwpcTj/L+Pfaw7f5W1t0N987k0AWACrsR1qCNpWBUJIrf22c7wwNwszYxOwRtqQ
XsrVKFLWUGbV1P7ytwkr/47i+tUGtJjYAbtGiccDSAlQW2Pja7saJhRBdGa3SdfO
cZ9tJ0lla05ejoRovDZGIv96Yjq4PnnIwe1Ob1g2GI/bnUVSadTP6gdXoXh+mmBS
g0pnX/iCrlIO9vnILKl4F9Mk3WeGAufbnxV0aIF5RjTCidX6Of8zxOzpm0Fe+IWg
Irm3fGqKx4zz/+Bi/r33DPzp+S2Eq1o+CzCNUwUIINCvIZzUy28/XM8cnuHMln/Y
VrqOscgzEo5s5IH9TPln3QHDIWptkWduDhCN2AfGupxYxw3QkH8NxFbVlTkFuzoj
AmmjLqco31vFb7kEHBzWKNHbMN5r60oQncNmP7NqYPrHUd2ZPDWysr7Jkp7T8qv4
oUSKcQXKcQL7rTGmipj8QBmyQ6aLq4LfN8Nxvpc3Pu/7sBTTrXW8wt9mv16+OGt5
Qobt2Lo17tZF5EUuyWGPODrDuwRzTQO53osFsLKvZBQRJ2QZkFIlufyyrHc/XbLS
GSsZ6ksQqNe4FDwFhBnDWf1U2HzzW5/IWcRbZ8p3ZVBUa5RYOHi1ElgDHrGdKhGu
53nsgI4C0cnJLNkG78fjXS8MHuSCGsvFCcNXIF4WvvLHfjWSHWrXxylNiV4NqbRd
PXmHpAol04iZ75YjmF+0uxZgGXTr7uL8S0Lh0jgt43tBs5FXD6Lk/dV+ZA5E8abv
2y0PM0+n6wOFA8Wb6g45gWuwD++wje8I3wAxo7jPf2wdi+Vl0QAFPDiWQakiF0tM
vG97bKHhAHmUXHcZy3oCh1VZqU3dDIkzGwZFI41as3FYzqPiZ/Zo8VOxFRjtET7M
WSg5ECQ8JgAC6DkQprt40Z70IvZ00Ya07mqmaiXAjVEGZpf8K9oOphPeWS2U/BV9
6uoLGqSHRI26vuUntbuYIV9axgS0+t013IT3uTMFNhXsAdHX+XT36gllb1XTGibC
BrMTeJzgzWPN6JFaW9S9zDk1AvD4hfkmz0OIpr3IytCBelJz81bhUx2GcmVlH93n
k+t2gr79nqkaW46jIazRmtOcQxorK/OWBX78r79MWLer5rsI5ybP6A9F5DonxnTF
/e8IjYbQU18G+VDxF1LGLDh/PkYVoe27aEXtB5s5zQ3miRL2GN2LLF/rBfFi8caQ
oUMTyj7fsU7LCyjfC3BfdxqDLem6J+wuNFUChtwRRNLbP2pLlmjzUFt91lTdcNnq
LXKFczEA5GtdQADrjHqx/aGlWJLjWLydyMyoedbBSY13Q2pzLh01gpdXIlnO8fpp
XbBdrM0/TvwKiC/UspkgRIo/mzi2QelcZ1dDe3lh9DdHOAsQSHqiixRQcAiw5uok
X0/JtVa6Z8zAojFafAx/zQQ5WxccFjh0Lc8+pshrng4Gn0rMNQxzJora5/XAfmR9
MRyKW7nZ4jPsEnDpAa6hnUHrlgtuA6WwtapfWUTDuWRk39KAm7k2EGoIOIiDcpsF
cCSxHZMCL0kPTogtV/YiZa+CzuP2WjfgWtD5bidKe4wouYyQINa4oYYq1/bu0JTg
imHNYrW5DWBs3bx1IDySekjeXGKCcTeyQ2PBQdz8yRCeghngouZxSx3P1T0SeyMi
ys6bOGiNKrxOVzVdJAIRiTb4wpYytUN/iIhIR9jSvgH0NARV6Ajll1itz8KxiMBx
NgsCbaP45VJmQBaT217nNC4UGuzIYGicqliiOazRB8cjzAPonnA9KIiHstTrNob0
GGikG678HbuEqeY0hJF3x3NScIbSk0Q/wzzO1+zNk/SFLsVxAL3h8J+z0EJ/EL7E
6QT7vQATJm/Y0UlczP4X49OZo2wsOvFQxG3dGt0C47EbT8XDDMv1VyEQZqzdAvE3
A7hSi0HmcNQD4LpGJfxsHQHHoYhJ/NicLoDJxvdcDTjEA5dm89yYPjh7wwTQg943
F3CkGUssMNzEAWQUA7SQKVbTI+3XqINhTiWmMc9dEsRdBL8CRTqnKFdPBPUJNNn/
TOw/4dVgUjq9Cy//954+FYwjUBfv8C3sDtZFPjNINlXEQLW2PoI9F4ZRxeu200e3
HOioQ/SlR80dV/hY2qpvJgaaz7Io6BRH8ePv8NLQU+iwpz63tTc5gkORpyG6Uma8
6Jdy8fOuQA5QxFobjIeApjMFEq7uWb71fnqkNy5ftiB34abhfyou1b/k5w8MzcqQ
kZZ/6xh/HKGvHNJM3AV2y8/zNEtAEQx8lr9Ie2mbHavj8zvEbPpjLrNz2Pn6tums
LwZACjPt7KtVdF/LJPQ14ukxdue0LGa0x7KKe44YtzRq862RAQjahjPoVoEwdL4F
FY+8H72DPlVxLFWmdLuLA/QROJtp3nQC11+PqvfP6lYvRmEhhnsih3E/w5h79mYL
qVklWA2eUQ05SMJ+ViDTNkA3X2gXWfRkWOeurFYMbINL2DPe5yZ1+lY83fwGasHx
Dig2oLXl2vFURghm3HPk3ULS5JzsDcTkwwYpb7uwEkYps93qhoRerXsxDB3dEZm5
oG22Ct2cQYrAasWymKvqNu52391mo7eK65vdC9FM/tW9bY2pvObDWJPiPqvos7+V
5VjgAlnV8rrqsXj+ZUhBKH+TIW442VmvWyYZ7TbRA6HHGK0xnCdk4KNUSkgp6nQT
wH3C1AR4H5YHAcDq2l8Zi0izHAzQbLxS0HMf6V3TU4A/MTObk5HVeEqzpZNk8cnc
5hNvR7uYmoZOIy8utVcq200bbfakDDES8DoVOawtLeFY3cEXjptmCqibNe0q0CFW
tUJn49BWev1beoy7ccCkqlybgxzsuzCx55T3EOvT+cbdI+dDixZxNohj3iIe/hCB
p8SY70Wye0JXgnqJFEPQ+StTbA5UbIVx+wxmkuJOP5o7WalkGcu0o3+UtKeE4tro
BQT5wzbZUERCYRL9CVruJEWIne+HQhh2M7YZAkDcB6nS6kUUP9bKlePdB87MmoMV
watD9abp2mpiunayMDS2VhIk5kC1AYEo++H+16JkmkKBSRgJaajuiN+4+2mUriIr
JCvbCV+Q02IPeBPy/2vG82huSNhQ94ZRdQIjI7cH9y009Oba4vxf7Wai0cYhClYQ
pHvLDCcIpJhdtFzOL89MCxXtCOKuXIaZQ+HHg0b1OtEog9Lc6NVBrID4QKGQjcBT
WKLpVQgAPLaIP1tSaN4pXkhBixazt4LAixSycG2dAkkJ9d9pKpBjElYa5R3DgPsL
hzstiosGAULWAaWokxUnmaMNTDI6+fohVTrYhAn9Y/duiGXiQ6INd7ON19fELp7Y
9mz1AFBI9UxA+A3Q3ERzOtfj6SNhMdBARkf3bbHp0Cg1gkqCXYQO//RwwcY0icQ1
CLVC2rsuPmHEkRuvYyydGgWeI/mVkZlBN9dHkkrKQqnD/YFDwjhGBdQznxpTk8m1
g/70vTEnRz0VMA4TQZ2tWjxfDCYv7UFFfW9ptMwgQKuf6sEMe+COsk1otW48rZhr
J069T46D5fKDkSAP8I4S/pT1Vm7/iFoIys23UmMTo35mRXXy2iJ9w2voXkYaVf/Y
HDtbO3dUwONKzRS4muy7HjN3LTH5j6Iqm/aSlXnUOMF5UesDCAsrb3bcr7noNAHv
kVhJdr+zJto44o7Tj5s7ZzO0bOScQVcMKV64C7d+dklFK/IY65T/Qf0VRxHZtVn0
sH1lbZy2UGnhzjkWX2y68Jwe6hbO26GnbwUjKhZ3cFt98FkKHw14j6mIGtbMDOH5
lKVtT3hgsiXumDJW+D5uG5OpH8+E/wHZNcbB3aCnRDfXmB3fL1KbEeZ9fExnWrtR
+coArBV1ngL2LFg2KZPviUXr+rjZ7/ox4u3b0qiMyBzwKhHx4VvZtAJZqq1V/2pN
ZdfpDmPAdekICJgOd70DLVkzSMXXrdlkupduSzmufIgq+WYwp4rlpFpR5+q9qUb2
IEATf2/VSj4UiHP01dkoZ+iQh4qdH1W/QmZBSdi4pxhXZR1EvXPvaqFH6FpaiIqt
h5wbC0w4H+K8Qsyft1tH3WCXodBRmQCYMVrI7Ho8pLKHZ4FcXRvAMoX2NdYYj80y
BI5QROWVW3754yeFW47vP6Qbo+3DuKuIaZFE5Nn/7PPR24/eW6VoRq6umiKgy1UP
tuW3eqFPvcctN/2ZTTLcmbBG7pB+fesZKmhlGZwP9x91n49He+paMvZc/fmwMC1S
nnPsMQOGsa72gb0aSShlK68aR4rkQRnRRlNV51I3qmCI7yERacHVVQf54/QvvMsk
O43HNB5s8/Ye86J3ZMMdLSRVMidbi0FDcOBNp2IZTuRw1t4U9HvGHNRxSC51vunW
lh+EeJMZkXoyPd5VDQx76AZxUI+dllUBz0pvAOtTQ+s7x0N2PSirpfHKPRkDA/Ft
XPx8KgN4PH2nQaQCc6DqpcLfYctpkv3BZrGLu81TMlTSiLmmFMM1C3geUDfn4Jdy
hOTqygJDmJc3ZG6+wyy6toD7RDTT+7qLDcHuo7PFCRd6MCR8kXLjfuQWTyGG83+0
uehVsLAmKho5S7fctT9IhFw7Kb5V0dM12XVaRlHySenfsbQoBllKn9KF7GgAoL14
Wkibgb6l0LgpkUn+idSdfU/EoBF4r1e651X9OnhZyUBJnLqwB0Uob4H0/qLVCRgn
qa6EzkBtV24MyeE+cpKIACWJKqX106b0nEjBdykS3Qz+y9snc9eEvNaEqZHKxtqL
wNckSVv8F/aa9/ioZWg3Ri0EXu7uInYgXNIVOVSOBTAAb9U/XeiUmzfAJyiZBLqH
ZhFNz/keBKYGHemxgbvWVt2Yc0s4T884lYUnAhMaMB3cMIIJFAStueaDyp/8v7C9
1zk3qPcO5hTbYYx6ahIxYrLDWb6qrlQ7g1UuYARq/hVX/ercUi8oFWDzIZk73HWT
k0xdp+gxtu5qaxMOfKcA4zB6J/y2PkdzGAZq9/PDaFyReQOIJ9JNePF/NpZFkThB
79HdP+cMQ8xwFNmuGGzFLbWREPjFdEU4Q/iFqKiFxOvJY9KR4Z78io1TgtPxXQKz
79K7T53X+wZUiF7wtASzTh2PmQUQalvIxllhhkbSjHvvsV7ELUA3QG67PUeRxaSE
WUcQd22e/w0Pj4b5++7gKloejDEVMf57Nhe24dQcfVTySggAFfAUsAphF3tPkeop
CNJfuMUSpcyWhZMTsYlQJyzPs3xLE5ePJn3ptcH/gFdmtq7EOZTo+0MvRmeLJzpN
uTEykBikj0m4i/QtJXXmSNjtOU3ck1nwUWq30ISRvWXx2m1QhdGrK0rruu77y1wu
MaJvrnsfghvqAYmF0FUSzoKp9UdqUQSOjQe0KuYfKFJ/2hXm5gVpgUSJVrbVPj4H
NUDPfVe8qGIExvNRKeTp9KI//kmFQBdTOdKoB3YMGsyHO2fS6XSfI6AkJBY80ef8
e+xkhDDvHY8GJrpxG+b9MxIUmW0frn6WlOdbCr/mjp9lYINUmI4AbuV1cIwekFb2
j3jL0UYvek71IYTSjHmxcc63I/WRU801Jvx+pYU/s5T5c9MeEemue8skCpdQKvYR
so5klSLF11QF4npxFtKn+EKsrlourLk//VndQoPE8L/gq1mKn7Wipj/GKAr9p+7g
RezZcvS6RpBcMoKL+pOmL6EWzTAry832LRPPo2QiHElq3ge1GdaY8EIYsh5GjkHf
iKClJBs1cuy8k/Fc6LK8A/5NfFPoRh77uXPwmXQdAY0+mzgqUrX3ym2ghs5bNNUv
yagoOD8ezLpjCh+7iNfBk/HFuol66zwXH5tl+JG4Q/Ky9qRbrLC5sTYUqG4oXZXe
SmXaaafqSBNwTraRV9W+2U0ROIvRmFirHFOgEKQzCeNU3v9rY1akfGG2D/Np5SjV
+ZxGTQoTd3NhuOfeztDV8FNUGfBrDg2IMltjNGI0nF7JZoGRVxvcWgVj2Q/Qq9Ki
S/MrSBUAEnLm+UAXAvsy8dyTreUebJglPjaGoMQBEWKy7FgLtcw1QmoGQoDoSuVp
dD2w6lnqO3tyPTdLuNFACZU0lBqks55PakbR1ig1xYilqBe0Ffv7pPfYSpLt0AV9
cgMh3tc7urP0rOvkJoJcgJc3U+J3Sk3uTtyTvQbsTwN7wzMqEXu2gRo2Q5FLkb+m
G5pFEAHLHduHz9UKDE9Mq5Oym8nKT4PiSTCuj1+ipkqmj+KcJdiV0d3tUFbOcMbC
/48FTb96s30xDJ0Z7OftqzdY7mJWhqDQDwCtnxuXsf2IjgFrXj1lbLvA7LVAxh1Y
uxs4PvhtinMdEgBhH+Xzzahz7il8phX9tZGpy0cEafXc12v7P6zsuT6l/UFqPy1U
MtSZ9sFx/0TnBn5BtP8crqoqn67cYuiF5GeOt315GXCMv4ib3xPDylFJPO2bQ2tw
0bxDdOTsXKZz6BKNYArO8ltTT4mJRbuiZiAKJOCb9EiidI40Rjh2ASEI5xCyc1Cr
iR1ooz7JEXW9N2ndIQ6xVz7B/hnOUjae1sbsjKE2Qgw/tbsqRY7+WSEOtOZg2Ohu
nGuIIfSvkWldsQtL7NC1To/BhaU2Lh7iYORqizuoEtOMzJ3+aOmKrmrVfgjgmicc
lxHyMJzogLb50bqEUMi122EgoI+6Q59HYnQx9g+yqOIVn5PfWODZS+iiU3GW14y1
e7qTSFIoMjdg8QlMO0REhwQSdNGeozGIF4DLOi8v3YutmyV3bLTiQ9sdMvYQ6zaq
kXusfpgXR2zfY7xdRytyi+n9eh4rEy7MWYKvD7FGLR8OIxe+Jzjnl2Ik4Xz8/+Is
ZXgRXLIdynVAaaXl4SFjZ5BPE6OCTdZsSOS2LtGSLzU0GUFRRLpfk5VZv9hsjKHC
/sbjHwGimS34kGDAwRy/XwIe0dvTUr3H6om9lGRO1FQNCJ2pk8g0NeMbJK0Jy3Ww
/+D9gzbqCS8tsqeLxXN4NszsPTyp8GL1pkJlDrKspZTWYQJ6fQBrGCD6nh8BvtGH
PZEDw89g/Y8wwCa9Y4/FZQko3hgu5YdJCB39I2Rr7sIwIBUZTLKF3SnA8CkPLd4k
jSzYP2s2hwvhYLL+W2cNP1H8t6CyyUazrpscBt97c2bDoTF/kKuitrRlgWRUiyja
yXYY/cRan54L7yzwhtzMyeDeYJRyeq8KgJCXmrK+zO6DBpcZDDb0B0+tNDEQVQ3z
dJelc9jXmjQHVsdelOejQLeOHLMylDnWDmmJ0Rp6VKACOl4R3yW6WC3ljTCZR+O/
hejea0bjvqwkfo9j7dQKQL0JPE7ZeBZQ1BzJVFrAAbMR2pGbDZv9OLe5RWbFxCrd
=======
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 33072 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
DyUmSSJKy9uR92lovAin2gFi/HKXuTYZ1sFuAJP8gdCyE64GNQTbvmHLwAtLvRGt
noHiL8G7jyrFwSQ4XkOyRoNTlyuMiwWdkBJJkSCnqzbV40WIvI1BeveeJzaCnDaH
66jlzBVnKqyKf/7T0N+EGEzo5m8cBbH+v/Q7TvN8HD3hioLi2MZokg9a2PWfA02S
gq+S1fHWRi2Py6F0or3DPDuhXVMCdy5+UI8n/bvOBVBWfTgbIGerx9H3MFlqcxdS
9ncxUj1ovvbWYcnduGmVF59ZJnScBoOUV1DvkDHLyzoUTkj/xwnZrv+pEUMeWR6C
8l73LrTisxYHG+2JugGzGjD2rOOU7uT7dOKAOULY9w4onBj50bfr/P0y0r+O89kV
lWkA6fGcKTI7dqdJs6UM8q7yW13GWt6lwVCvN63wU0vZ7ON5x4lPwx4dWkImfnL7
elGtAaAZcksVm9lR2hLonrfaDrCg3eJXtEkRqTnKc768DYteSwF/fTJnm7xto97c
o30BEtxw6nR5j6IecBBf6LcLAH84VBk2KPbQwRCDVnsEvYBDUEnjgm9QfWwVa3ek
R+1kQFqzLAbcn5Nplpwayh1OlQCXE1lZo76EuzuZpviA6iSxq5NrVtAc7rG2you8
Uy8m2old4GgGXsW4KbWvX08/Qt7js87DTVxJPVlQCdKm1vk6IgRk2X/O8Oc1PC2N
/YQ0K32F7TJ1QSfRH1cO1pUlLTYTE0Y3TNy/K7pyK5nLCrhBDkp2kTYITpkX3siW
M+fLHyVfLNHuqET1PPHwr5QYfYz4ZQc7kdT0KcgXbh1tvqf6zJr4iDFsELZUfAw7
ZimOhzyVt3nqja0XdEZ1ynNl1+GaP1Iswhi6Miu44QuPvlU6/Xswk9WOeeir3zrW
CX92scdTtzDx4waUpSGWT22B4+5e6QGcuo9RbKPrqTbnQtp8ZT2vZfhFCqCdt0zH
uD4TV8Hv75q2G7cVFqkfeCao7MI2Ys68TgjtLG1kKyg4bwz+hTb+KJCl8IM1xy7Y
7HqIx9/Gv/9v4xJVb2ZrfSDxAbUPDiD9ZCqEDTSFfLmWPodownGOKzWNmQUz0MXA
k28EQgh2z+YcojhGP/tuAXMQfgKLAMemtEdGGobQWagOhIl5QG0oLY/stmUjL+M1
WwQhb+bbp+4nVbMrPB+rfchT2d/6Pyi6nDBeaJ8lXg0AefD58I0vScZ//uvvzYPp
e+r7RGbjPysdLFsde3EVQGqIPrMsTYPKikPqGtu+t9hCSIG8k5kNvaYg48YfbkIq
PPr+d8XCQuI0aE3HtxXddUxC20OKyDiV/gSrvqHrYRQz0CFfP6UEPaVnN1koX450
yy0KgU9RUsAYd5CDgOewWeFECr+aXAs245umkYN5JqitQj4maLMsdddrdpfBG17L
EAn5ErT3/Bcq2QhAlcrxMwN2zRcGXXVQEcgz4DC7gqvUwrA2lmUoLrNnWuwnSuVx
04ug0TrpTTqfkWLHnIaPbpuK63av2adDnq97uitYq4L1+Hv8Ey7TETemk0dtWNDJ
dPyglcT+0xIxaI1HA5O7bgb9n4odlMXBlNyYA3B7KBJ/cMYf2/ja4TIfTb2gNEHZ
4kRA4jwW6XxxuHcO0X9g4J/59PMetI6xBpoEqz5F2WU38NVoJyeOwwrP7sgl0/Kl
ml3T+32WPQIVGgDbtbfYdGPXTVskfYCakIjD7EETyMcfg2zlFWHbjujzbBFOxjvh
DI2+US0yCkiMIJph/0bgAyudWTOAL17zNhux+XBc9RBplDGFMuzHrWOd7MaWi0jG
O8SS/uOn45QYiDqZthj0sP59ikxF4Xeu9dabwEoGB81EVZvZo+tnGqIP2cRLz4TD
KYlJZRT7aTzJz9xvWUICFSeyupMdJzwC4HMMBgZ78C2QJAqcPaiPZ7XetdZA2aQO
nmyttyLLrDSr0SPoTH/zpq8absQZAJqs0dXXwiVj7E6ej9uCXBLNT5A3QKZiT/KV
O5LqnpHDa2ThQZfSd+EsbOlCrftTI+Tp/21Z3nCZSYWt5g/1nxH1JG6c824joj62
/PQBjPjRXHfQZ/JJFowjfXvgofv3DsSM/fRQGZwWiAlD/KuB5jqBmOFYxGFaKGOM
5IkAui4xpMAStgklQxSuhItPNFGZVsgWm5JG+mp7k84oyTELTR/wselnqL8VwTpL
LmudjwS14GEfadWUkERiGY0nIbJAYH6nNtvdoEekYno/PaeC6mZoTX++7UKQA2MG
jO4c2TffSr+cYdq+IM7zk1guz8eqAJayWiumqcdU2IosEqaUfmG7oivPpJpd9QTa
4+hi0Sx7tauUL6AZHlPkZlR2RF76G6hCJOT1WgTaJf3CjYBS6hYu8WHrhUp5rkx5
zhUCBIt2/bIqrr8ERjvJfZuCOaX60K9jWpMe4wh4sO1lCbHirtMUUllAzkB64ji9
PCU9ZCs0QC2mgx6be/g/WCnqZ4ya2XTZZmVk/VtZXTVwJ3kE89Mb+cIjWMdh+/kq
TrYlYJ8HJW0YLCsaRwiInfZjfCG+guRg1wRo31ZdXkA1MtS4vKvyi1R3W1lKJrWZ
KUmsSQycOwuI1pL+VPRsOflXNL6+gnAZSwz2xxULKhoJSng5t0ElXTizAWulUQ6b
+2afxhWPez0Pq4kYwL6gV+81IeD8aZPq1LlqUhsVSyQZuSoNAoDQJPLLNwzU0MqU
C2V1evvxqdnBh/4BDwhQrlPBnzaw8jBU7fqSqaAsG6gnHJlkEQHx1/8+k7PrqKbJ
DKWIHg3/GSKid3KnjwbC0znEV/rxDUul7ThvwrZ+2RER3hqG14+htRnY3HbZCA0m
yFVqtMwe0I90cDTf7a9AjMK/LtVac9luKqXsBsK2z8JYo5NSslpWWxqeLYuUNcdK
ysA82255CsylZTUd8c4GMC0PiAc4jh67LVMED+jv8EVlNXDarUdeqTEomEXBgr0w
3EVPuBWpK8A9Vex8mdap4OkoyEIr227+iogosQN1HFV08u6LG89qd8BnBD2v7yc1
z+iEwmG25pMxLEFMk8zXqSOK3vqsd/tx5rRZKWI1RkJIhXVbF/Yq/mx0LKWI/n+D
//mtEPfuX1YzO08C+k1I9MqYEEylnEvHv/cWq9ZVD7Sz+BBYjM9nM2RzOGyLAY3c
fRA2SkqLnerWuELUJGzPoA4x1qnuWY44ZcBKTvUNxMtdsaka01TFvMH62j2G2G4q
iNmu2VPFLYnFkXsSULt3M6+b1kR1OXkb2u7XfZgb92QhTrlnjIiyhrBx2+qEof+7
y2+GJSjX3f6nETj4Lny8i2HrcaKeiwDtu3QLV4CfExP5/sJFlzeanw3MWUyh9DZP
ZDm4gdY+OdieyNcMZxABgVSgsJPbB9PQnMm9L2l+hElZEFPiF2+vPiuLXPv8Y63K
tU3vuolAVoBIpPCWw8qUeca+1zRvWJT37ev1V0iabJlFq6LfP2flj6mKX91CDO/4
Qh11cDP34B6AiLDnd0mhK11aw7EkGFnXsGS2vuQx74ECFHoOD+8rHFecT4LiZqA5
qlOLlG/vmoDdLqtIcGlOlu6GTgNX3PDyxke0OzGX0CwecjYBpQsSjd7cLTMd9ZpH
K+YVUhocHYHRblBd0Mb4s0uxac12mCks9rAaEt1S0UtRG1w0WYPe3+6dGBATDTkJ
ffrPSSAqiHAAoZL6MWq8/PT+48jzuKDa+xAbdmwMjAFBEeDTIxfhGeViaT2WEfoQ
TTc8LpK40rDL5Vq3OJZjKLDZeFQGaVS7DWq+OCvJbd3eREVVm2VpSVeALYVU6jy6
Q+iAL2iyekRg2TPq8Ty0BLUchL4hZ2RVgZ2VDW/JfvI9lKantNE8Luwu/pxUp0sl
zh4hqO15VEBd0rMQCbvSjyB3HAHtW11wvlow/C3MUaDUHwoA4mNqCCRd/LKFWT9n
oXwAqXaxS9aXbyz00EfEFZDZJjUnh7JBBPjRdNjvsNVaKPM3AnwqJ9nuYJz4rZd/
peOIJ1zXzfBqIyo0Wn7FDbVREJQb1m+vAXr7Cx/daYd/GzbAqsdHT7FvvHmZff90
Ai/HEDZbToTS9FjvlMjlygJMeWWvjJYnLiUp7J/g5vCLvAxAnxvs3lhAx8U1QF5n
18XfchOOY2cVDYUYk0B7d1o31wo3Vh/9L9dToifP+zo/89AbESv82Qk9BSQPuz/3
cPajmbCibXZARefdhabbQldrmvG+9cdJ+lj7NeOU0GYaqdBTLafM1P/GTeHmmSg/
gPIcoAAC/a86aySoaQJbc/gXjL+TBjV94JN4xTp9jc1ATnoy7a7yXTuG5z9sggqy
V7mrT1Ii6FIggX7Wd+QO98LQKDUQbC5UeqW+1gMIxSY3wN069DJE8poHVrlKj4Ls
CzEZ82vKbf/w//FG5MMr69l/kG1Bi2iwGjlScACDhXRgGRXD67OnkTUAOAi2slS2
etfZLSrGUKKaeA2rrL7QcXHe//eCDjaKPyxHL3moOnsVnL9oDzvF04UEsEpQ68xQ
amkY1pSbCwEUkHFvzyPX+qS2/YmcS2x0PTPbkGB0vWTOL0lyk1yjNqK76qDe3kJZ
j7BL6+y/twisq3Vqr+ohme6V7MIJ07oRWgBBztNPd6JyGxmJ58Xmb5TRnSmFXms4
Z9mEnauGyqdDi2U51wZuHiG8aU6S7jYCY7iBIS9BabXhlsBVcYzYCKf4cL+H9BDI
vDgvzoSWSL5UjmIHm5U5o6ykN+fi9+oQ0EyyI4K36Cg07tuQIguc2YLYUq6cAF7D
4QF49aI7aZ9Ha0vVpaBBAeGnDJprwrg23shQHmhRUf7OZFkyHTDMmUEmi/kmUCUp
Ks+V9rP/oGCOyeLnruNXUJ5mL81l2j/icq0BwfZtF8L29RFaVAiYLB85xVWfhJG/
nnmW1v1R7OJwuJpsl+6xH5qj3GpYqdg4vR5sftUcGuwMrlqRN5CeZ42X7MDUdTIy
l+3vJILmY0+rgP5UQLnMuuDL32xixivJm1lwcnjUwacKmTxyVUWl1Dopk4O7wUyh
wQ9geMi2vzrs01eFXdwC5Ke3sM0+1uEfSdxl3VbvDvdBf52dW229wM3nOY3icU6u
wPuXDlTwFwNRc7wydz1SIyTSkdCjoQ4CWndqtrpbGAsprXp5hNBfTtGX51n/T1I4
iwydb0TPwih8WQ2xzATmcBRdzO0WB3sHkZwCqK6RfaA/WYICIMFTUhZpxk3ofE/c
q5o8heCmspGDGehgKB6jXt9V6h/6iukHM0La7qIX2hT2c2NczokJDFzhn4M1t0+f
nH+Uz6qcELKbyNP1aI9iEMI1opD0HRcWs7CkW2xdwTUnVRWiNS3wtlzIkueT7WGT
gSfgwzZ+0kS8Q1nHZoybV5HiBNvjIvSYxSXcukxzVTeL2Smf77W16eh+tG3veWY+
W4u7Rl9ELQdK9FN4IpnhuezWahfn7+tXQbqzDpgeewH/V/q/RS3xjZ6HsuFB9MOH
N3gsQCM5OOim7wfDPTMMjY/4HeTN1Shv3gFVT8rm4SWODLx/6dhStUcXmM6+Qv7S
zMMJ3T+D6B+wHIEU3L4yhRWmfxpTLR9cGVH0bUtnAh8t/rUD+aXWtzPD5dpCESAk
A5IVkrDolUl0P58RMwMLmjomWr0IRSzV5tgHAG29a/bf+IxDUEE5qDkBhwrC1CgI
KiKN6W3siW+thahR3mixhjX9YRQNVWvW7RSRIhZaiggVxvLGDGdoO3Z4Y6yLr4n2
g4VQXGNF96Sj8OPboGiYIDST7ZL3APNccsa7NwEHqwraPBJ4+jn0VqncqPaXQZgo
Hh+FvmazLjptHILg5c7KNqN1P3svdixDCy9lViHYs774d64tyuwlb1YimYKueCzR
m3aa0XOkUj3cYYZ9OEeVo4SWg5qH5BnKa+6ZH/vK85lfywxMMOoB/8m7Db5GzNiU
HzgxI5k44h7rtkesIaDEaFpiY8rIHQaFxNZ5KTxduTqDhhpibrAHcjGh5zlrgfES
4rMrP/+S8XilRH1Ka82yS+y+N73ZSplwNe6avpt0LMSs1/tE3FDLCII+u6Bui9jP
lTlbwQCHtAsi8xoz0ryxY0fSZQRd8NBhtI/zbKlFvg1f9IR/63eRS6T/32iffAHq
WMYb/mBcFaZ/zhyUOqMn8GpIQ9YFOzttWqyn28KrXKzSwnBJndUfgO67hMMVDv3b
Cf2TunOztRzq8U13szhTcEePava1frhpFoXxarmxALTmHVOFGWcc5XN1akkMg6Rw
SRgeReCRILQXWvbYVXaF1fw7BgChnQDWN31xJYMRHMMSADOmbVoloI/2xlmn+yBD
xJ++HqVdEnjZg0hkpdX2y4oPdN6ZfnB6bAxDrnrMSITZeIng+VF9PxXrZ8Q1xchz
coru7zC/Oi9qHKa+oLjyQzkcLEyxyVmk2kzS1V/jtXuhwslW1c2mCBqwuPKmoag+
SJpe59Jd3ywsSnC3rUWXz2brHWWOsDlHvzUm244yIR/9PVHixqUTSkN0NpkGj0go
yOc3ZVEE+s+FKk3CsAjxVf5K1PYrZlNT/S6XAaXrtOO5sRM8Jd/4ocEu90EQXy6e
v98ESN/QN7MGRs00QQYa/LJLOI+lynGnoart0q+vlj6ysz/wbyefNrllMZwjvSFW
RtxRBh3pQNMTQu2ulgrT42T4aa3y+XPj1yJdUkdK4NzXOvOxjnJlkONoy2t+01th
eQjMIPkmSUxB+g4Ci26RCmyRhNQ4COpHpL0OJfUgtiwj+iaT3r91w8omk2qahmq6
qySg7wxw8uwxvgkOtl9ruH5G+3LwpohMzYAwNMROli1NZBUlHnaBGgumexYq4Y6D
/atQwHuL8xMigk3S0mnnH/UA3CxCfQeh92MxG0bTlAm4VI1OD0kVuEoHZs/HQc14
wD6lDJbcu5PaH9n6mqyJ5gAaTTAfR1ytcLA8JIroV052/72hYIAZRwO+4erEOlTa
B0dyTqAJQarltjeavm+agSFC87PGPqaVJTuZltYusjXU3Gh8sYtVXEXaZ0EDbTV3
B7QEpQgFUZosZQGfiScq2dK0+bZXg5MEvwd3uiAyjfBfG3JCZretJnPl7k88zMQc
AwN5nOMIcUj6IRryC9eOz5TCaWWBNbnAHhFf6YHGSXoAoD3S+4gTe6bPyhB3Ib5E
vNlJu4dS0c9xfLhBJUtk3ZLMEwNfSFh9F0oQbgFhuJxMzP+IpMUHJIY2WZ4Aib3h
z+e+TaxT6t/VSZq3119BtKWCFS6aDXfpnFtn17k/cUcg5tM27mwpDR8PuptaIVch
1JwYuT6DyuYMzTqLB29oJ82KLUBFB9+zRhPG53iyCSeoHX1FhGftnoO2F3PshYMv
QXXcZbfM3Dpylj7K5hFf4RpHI4nDzOnJwszcuEnfT3SA7+4nCJ7K/Hde7qluO37C
ZH01vdkNMabnGchyvycwqjV+D+XA1tknyWsasfXE8rAltSbb9B72SwaPX+MTSz0f
VNZTWFi0k61yV13XOqiC60VueTa/MOwIpw26n+9XiGTMGeZxGw1ZUeNT3YctfgCr
NlLjZ2eFYN5MasK3Bw2PRFRe08CcynOSfmcCnn/HqhTGyAFS8wFNfCNX7D4L/C7P
qutF6HOrHu1L/cOAxBGt+3olcNhkd3UPpNZPxF2Ysz7oVgaM1cf7IR/5deAdSyGM
FBhqFZgavSpvoYrbZw2hEjZ4RznamlrIuwL6SdpEYtl0VTWGxIhHaIPwwECiwoKj
UOHSnKxtijkYvSWPzVYhyC5CfOB2PohoyvALdDhMKTAoCr5PwqMdkvQafX7xzHfn
lkur/bG9RqU89iZV22h16THtg3hunnJn8cRUezDU2TuSOgkgkqlBHwc+44xfTza+
n6gxuphw+6lprE48EGVjxV8Tf17qEDXYDaYzFI2xLbInyOc6q1maPEeZDtFUGtKR
QTVMADKKo4k0slOoo5mU6ZqYDyrJfYUem9k/05Na+7c/mA1hGRFnm5kLuT5Q8txQ
X/qiJTOXbiD3xbCMs4QbTZ4IIAwEDtIIUZm/gVHACADMDeyGQx+Jm4h4PTPJK0v3
UbzTNl76sri3j52bhw/IT8pVGCF7IOfjbwFdjEyFEznE6gvBmkhJK6VTZJtOzimM
hUsIIFrBejGDnLXGnBcmlL2F5l9wcjS9DWNgC1cophlHpT6eQcFUInkN4UqyacWI
E8z3UQ86MraVlOPVNNxdSXXpclEfk9KdlrKtAYCXRjxhRA/wftVaCxOaAUJsr2oe
CHQDKb5iNWX47LyFkE+CeQshPnvwA4irapKNdvaL/eU8XX6/hlOgRZWa+PfYBiM0
o3euLYHvJEDRgomumxmqeVRTwI6K/k39EsjejrFEF0yi87EaJs7gweEnhjRLolc+
wQ1bpj/dWOvHIZQUdwU0yO8jU9c/InjYdYOYl/fO6a+LYPrKVKVFF2XcJT6zzuqD
2+7nlcHs3faK3YJ1+N/E6sZcE/MyCiM6J69Qqw1+x8LSbh4QdMuvJx6d8wDmjc42
P+F11ii4mH6vYJWA8ntkHlGZEHkIrQq7lmsrGlfikqcwBnG2Qp+BJLJYds1TUByN
AXw+6CdE3Y8lQVB2Ss39zIfC4iFV5fcPcSgzsLLq1qagtLnOp6VMkyDebAxV5puh
NpglEQ81tWGYxBkwV6xhKED07BpHQfsrcz45v2HXL3XAfiF+qQJp6ZiGLF5k4g2f
VChhpfSg9OOiJNqFuhqBQ78rx3Y2h1WueOg1ggrg5FgNSrptMIQnSP6M8Bq2j2um
R6ClbT0or2Ci/p5pM/B7Kiy9kHgbp0H0UZ+SuNV3xXFDF4ZD8AEWG/gSCfStuiO+
RZKIb24/kvLB1GpCQYfs6S/idxT9gB+B1h2jji1M8fVsiGHjbLXkX1lb2tuk8W4o
dyEIHazENCUYl3thwmOvNVvM3aEx4oofXxtUsfQORB51qnRPiqa+wpY2g3PEN6BO
6MZm7FbYYWXYvktqIl46nPZJ/RdkLkB3zH0SgvL++KSb71uOhBJc9t51ZQ9zRSr8
j9FP/PH87rYp4sJ7S/RguCAW9XWbtXUTuP+018G8moaFXwNlxb95jzfCDh4Rz/Am
PEtllOB2tpHtRllH3OjGP5bRkci98ihbsPW44w8YGcVy2gyLb+h4HUpGeU7mkolO
bNX0CEiQD22sHdm+mp6B2uz0KGIVTeNNusH7oow5n77zC8hZpoeGEd7PDN2Lcngh
12Tnf+6Jg0OA4YxTFWSaATIWaSywdBfCfN8hU6G6wo/v6IXitIAIML4wQfzK5E2N
CPOYBSzG7Y5PXNuRH/IpmR43jVitSxoA4aX20WIw35itFZkInoi4EKnTtiJWQXHq
xr5NkZq7goLwaw5BtkhtByxLclxaffWb3F0L8PZpnCSr+VmbdWxIHn0/z4c++qKv
0svXPY4RIPYn/J21qZNy07cSyr91iGmdfWOR/GKkMgfKN/qRMJJbLHgwHb8rm1hg
PviPTCimx7ASdOvmwDUZL2DEQkzwuFjUz3GbcZ1ZwMPmHvGqUogef7Zrw8OKp1Z6
Gsk9FiK57zmaRlgoACsIZ2qseSB3CCdanHrI1m4IRMYsz59/HfCvUCyKJWq2RSRh
4bwnn4tJtb09IyApEmX1bMVy7COTkjm2vLoF2uRfh7Cqxg8ezfy7chlXBbCU+XZg
s5NFB0m8knMOSLCgaYnt2lxJjg9TatBy7yyzRwMkIYdT8hjl8Dh71BCtTksyhH4U
qA7sQMCXbVu0jsQ2yMPtgk51/v9SEeXMhuzX+Tr2v4dI9awocUN1gKgqmjjezMhB
I9NNzQp9in8Oee62cg3+H0GW4arRFnFtnppXMiDZVyHGVOnEP+kPagENSaxacn8M
ekNjk1tpaXqCxxj2OpHZpifcYYGj3MRwNQx2Dk1Lr+R+J1/8w7+ldj+31LZkVQ6C
fklHeyoy/mdxNoAaCE8EMaPChS+T7lvq69VYjXsemRrRaGzh6hiYnXFYybjnjDqu
yboXa7Dnmk7kk/Hf+5r36WmJPAPAUB7jBnvDHLfcyowYyVCM17Jtr0Mo7ySrj5+n
9DKu11mmD4FcNsx3gz8suoVSXec2O9lFyMagFoq4dWCYn1FG2Epw49TfBQKVtdUs
bxJw/2Y/FcFWdK6fmaxAnO3Y0YNcstEjjyBEQMPOrTrr0WpAl2pUevSdFXcUFVvG
e8DvdfqIYop9otnswhVTJljvU8xzNLB1/5gtdZKqtzIc4nDiy95hB7ZdJlzxFwKO
1FxJiJ2roAXw0p2sINMb7xWa466QkOB65mjlXFtcL72gOJA+uqV81v4A1bWk2vgt
IUlFG/n5OTcCNaJrNiQ54IyeT1FBVEV/6933E7sBB4DTKxSfDgzNz1mAas/202W2
BlAdOUn2wFRQ8ZaDDvpo9GdubpTr34uGAsJY1NUBRZitxqJneLr5kuVmTtzkG1CR
My24I91HNjkENna75iVEvhyTt6NXLz0BTWtXM//v3E8eem5LbM91jaJyruCdh5gX
jz8AL1wAojY26VVuQUGdvDHIcSW+5ty/NRuz+sFua6hXWJkGg2iewRSn/e883Iny
FxF6ko0JYzBsscPRjQ7AVfTmriCtzkNQkKHW5p46qZM/S7wcH0Gi4GlHHjbGM86Q
177t/zngIHM0L0wNnyAQl5/iDsaasOi8tKL0XtRg2U1qOt80zgUwung4E9nA6Iwz
eg3ZhYRpkxvlsmFNfjjpSPWK+Um5WSv5Tbp1LvmB5VjpGHYa2DWAY6mYq2N3n1yd
TwWOd/HQzAKFekP+rqfo9O9kXahNgBSf4ASdDqPSXCmn6UIRFwjDvF9VDLZJLwOz
T6n6ebIvzykn8btwRo5vdG52vYi/MbulCjjRn0EGfPWZ6LCDfeBacKFK1vn5qNTh
30cyrTHI0vho5+OIcWU+XC8vVvNaohpm3HVGwrWcY/6w0mnzij6BeeNgE16P13J9
RHD446M9us+AqDAU2tmxQVhAF+bcthxV28wwtjSu7ayIg2dwo3Z46azSIrZO2xyc
9myh983vS2NbzRMrnyCLAdz1m3oQKSEqASEbFuRtsfdB6RgjdEWLvkbbY7S82Pfu
PRNePdQpzjjZvlHzhLlwbsGPkPCv6KojfQdsstK3kxUgnfiu1qege41bO7awqiyW
kM67mpVkkeX8zmgftNUxgs92WTAVJwyyqxT9V/GzTDU1uZEAwszJA1xJepg8/+H3
HIvCo7gWkzKPo+ckwfeOKXdIsopfROyHujJG47KK768jRupKPAm9C83g2Z/v7whB
Vmz1MufubqOJzSu5r/cQS71P1sAL+jcCXqEdWm4hrcw84RPgpLkZoZ7J5gse/zws
05R56Lr5E3uj91IibXBASGSLph8Irl6+Np09GiJAFd4c23HZqXHjLlevPz95bB7R
xZuHZg6sWDwEr5QvroFmdvE69dbkQZ/WR8cdgBsWKytWJMkMI69M1oqof59kl2ZL
g3IqkGtYuSmMZeWnM+WA+MN60cXPW5nogh1JKktriFhAZvSmASW8sGe8SOZO+Bm2
gh/9CGWBDVdpi788lzfsA99KrmkhsRRIp0MTfpH/CJld3vBqUivCnaHv5JH+6M89
zJbffYa4FoHkQtJRDOGit4t8LV6uuIeGCjAIUEnvGPtBMxUD54B8VyhymC+MDtj1
ycMcMUgd+oRv4Nlkm9MD9QxSPsu4aHui549sHBjUG5bcBwvSvy5pJmWO4x2ha8Nq
Y1pyx7NsOGzBGXbYvCJOGn1hEFE+oPz5MOxdwayVARm+uxBaOfcYKx0btrSFKhWH
9YAFqx13WK2epTZPyqV5Ift542SfWH4f8zz8DsR8E75bUkAK4UzIIfZaNpOmBAZE
6D0sIH3KDRPG7yJoLLFTVOOb0FE9zJQPqAriAzRf9DRzpy0YVi01IJMz3EE6dobl
mu+yt7yY+O0LP9jxSe/YJxkWl/lmt3SAxL4w28P9sO4Y9kjwZMPnzrS5R5X7XnaX
FVnlrbtF+53fkWi3V7f0EobnxGKXw5+kK0MQwrotvforgAuSGDZr9QDc3kqZb+ag
iQqHXXuuX68QttvKiyOCUphcss1nGYgnNw6xJu1+P7+qPWpSWBkbRg9eWXj8uL+e
lL/jESa0oYJ07S1ZA6f7qvf+8evBTVbWZK1qp9iwIPPa+N+1zCQhcuo1Bxy7E2yB
3WrnK4gm5yHoSf300fFwEgEWn3Ly0Wgwgy7X3NI6wNh720nECdyJ13jvVVfdPI1X
HMnEYlnthUJVJ94niugbGUt07wg3zdKbdZWm4Xb9ajZGpqt/pZzqQ5RlHhCq7FQV
TABWGGkCI6ZxDTb5IsBBCCyjZEUl+A2+Jdp+/Hnggnzsz+p7lVwqLZ6ktof+7vCH
NXHci3aLbq31A79PEmYfwF2SIx4eyGeznLlDJLVML5vQ1zUaIIgoQBKwXuE7gYYF
CC8ZMjZFc8xD12IuQUVJwSESUttRrf1jT2M28FrH/Z7wDxLuSQ2WtG8lZWRdta54
J+3i1O3VtoUEa50Rhj6/GZWMT4dvX0S8PIF9pyqs+kKc0cji+rwJIbck7IsMog5i
F8EXHEM1W+qe3Qy2miBYI0Hb+w6XbASCko7Yq6TmDLgd+XOKOi+mlVD191nuyPWn
pwSIlyIhx4e3xREGa+zpM1Q2nnzSjq/K3S6aCF1Ic7CPODZgr1dsb406/WeNJ6lR
s86mGK/IE5wb5ccbvIGe9+CiiaNhyo6JbrxvfM510lUxiiVOpbkH6jVXWo8U1Xvj
CqnDErrqoycJQZ33WVMx4LJ3SNlw+0nkcCom621zIJQNl7kroCF6zr0g5hJ8l4Ab
5GUSiDDDbN+YgBRBABcIIiAmJBB3KhawGRqiGWWCrUOimGlVd+dQUG8DyBBJiBop
hUMWurcNM2flg80Z1E4WxpsRB98mJFjED58Qe0tCpaw4qIz8AqsPNuURXsqbGvme
HE+Zf5+MjbB/QBr+LY6x0Tj01Tgg5uakitnuZiCT7Ja2YxEu4TKOWMsAkM/aXBHJ
O+8KR4A0hHDeIAdjRSsNPOQ1Nm3YPI4ceIgPtJYf/k+aQXIBzVMP2pz0Q7utiC7V
vvyo7rVAc+dTv+KOFtbgG+quxuRck+pJbWJVYheK3bZFc9Q1gymg5MFlsI873EJt
n3pnZqcUNOReZ04XqPZfwMVfgQa0z32iEoJnD2BlcmnrBIQD3upU3bo5w3YMRu+9
Hzbqu2EQjxnnZDgOBJmdHou2XjHDvoy1G/GAzTOy6UYVrKNIjeGLv9MRhIzYDnlz
Phl3tbA20GJsFsUZkvw2JMavilIZXWtGLEJ4nLN+Zu154J2gR4s8jtD8Y1iZiHNZ
/TJ01t6swT6q6knwaPDtC7LuaPUnz1U2zpIUKdAuR9nFPJ84On/5kGwVkneJir5k
YJ4grMPwOe62j66MR14J1pVFTzpUWrlNik4rqwjsZFdSpfIiGSxN7p+S2XPxb2iz
yLkbdUE7w7LBt22gc3Qzq87TvimeqpWySU+XEcADAhmZgGXwqXHr3cJY2L9ENJxt
aV1x3TQkN0fo82tTvz5gKqoayz5IM2ZzOKzGZefVhn11f7VeeGA5OqST9UIlRx8G
cPQkx2QW3hk3l7nn3GznfUXgFbkKGBps3OfNayTTNQt8MkcFbMmD8pGAtDrebif1
rwy+2lEoaUceFIzMI+Yet/IiTYqzhdh4vS80qqkSWLQ2Jwt11n7+cpJXmvm1JW8I
yU0H0BGBEzRI9wu4SLSsw+socd2Ell+MmZcoU1PQkfLdgBomWfGrrwq1VG6rMbbd
6LGzpnFJqfUFF7qAWaMURDcOolnPk8cwTkYN6YDzXtHGSDPJimWdz9d5nfhD+ewr
18mVXRs0dmEhAZXIGeuWksicmetW6+b31KQOwOBZbGL3m1YCQBy1zK5TyL1IfrUJ
yzL90GODikpdWWr99NS6TzlAdRsA9IwQWRF54foXF4Eare7PI/OjzrO0nBSeaRGe
eP6uv/ygMeMceneweBqbmnj3tvv556wYvorSrv+zyRMbHZEDHB7DRxuprPGCzE3f
AKDgd1xHZ5oPp2u1mmCWxK4/5hSszGoiGjGIcFvKpwwL7gKNE+e73opYar7jxrba
nyfZbANNSLcYrOf6O4QYyyVIUdQD6zwVKf6SrgB02z8mZtarMGfcheb8etXDolxV
tMXGoRuCQuKri4VDl9uSOiw5KLUOE//tPMaa3vsFUXhFTIfliGa+Dpg+G+opkRlb
cDBVpuvzDon366bduweAmW3cmqiBmNl5NDlatKxCUOpOgBdzfUQ1lmIrg+543rMu
UWth4/1gi1Uvdr7DDT6GLIEADgfHBgntY7bG4uZcKg3HhHGEyzxfw/zSUq1HtuQo
qeK3lnu7dHT5vRsXgEmQ9uZUQrOASqTKuqAIkXjYE111ZobGBNT8Un9YUhrcYvTc
CllkSoQaFI6d9AOdldm61Aj835d14qJWreY1ld/DrU9erpiV/aQq30j7KgHXFkJK
Gfpl8B+hoKZPVSwc75HbuwAFs0opBMGcloc+J9ncWfx3IXID686z7uhbWUz73n5/
jRmu3WXQJsTk9hplm0Gnn4hKO+8WP37zFswMLhexUXym93+cRdkwmwHXcg4I70Fl
jLCgS6xC36SYts0PB6Tx/soOQyLm3FhFLBwzXVT2XuSUhikBr3jMsDo6ZdjnbkqC
IjDJRVj4B9wIY2pAtrReqEiikVP3RxuYzyjqJMLZxb6R3u5rEBBow85Zoqlu4teh
MhAaQYjH/nJFlz8T1ilC3nMOK34zOsNMhydkGikfuHw/k2Sjh3CfwXOlXdoggoOM
iIfzr8ch/clQqxkD661yR+X9SS75VR+OsCYNaH9MA1vSWjeY73wGVChPEzFD3jND
siK8xRkrRzQECyr6nNCrV0a0nOI7VZ2Q2eKQDrIui7wCM1S9plBZn6//m2t2qqHN
Yl6aw8FkymOiFhQboJnaDWEQcxWUSIDXLZRed8sgBFHblu6IsuIlkZmv6JQ7Vr2Q
1l15O8i5K4ayUd8OnMwfYY8mnwj/j3hRfoARg2rGkJh8gIpyAkUvqlWc2TzbkYh3
4GJ47IOuS3QnqcPHrRDPaEnn7kg5Om3AfNFNDidO1gda6WUuvSFJSdkeeR+dcIH0
cwlfwDJGo25Lb5K0/YzwwXXI2mln2XuL6Tt4deODhuQADer4sW05tVwrNHGZqSxN
8/g7I5hsoXBJ/qp5fR9vmfqMvsfGcfdisujijueKNiEC3qLdD3EenDwOT8kpTJPv
BWJeE0Ermy3e5wRtDPKqFCPGtV6HIBAEKit0rBaVMY7LGQuuQ0tQxz+uuv8FlOZR
pVmSSHTp2p4E5erBn74S+2ArQesVidt+Ki8hkynrab8s0ElBr7DVFX40VzpKi+Zq
cqkCo4E02zumEReMyzo11Wo55FozLqZGgneFuzzkhdpV39/QRCoHpAmItCz+RyB6
N8U8Oc3IWjnzK3LHbsNWD22S5U6CXfthPr2KBK6dLzUSwgl7hDqq7aAgEguiThv2
EMcf4hP4y8o9oCpfI0rhUzd0/54ui+qaV1bFO9nmhNPNMjfvyyMCvgq5JgEJn3+b
L0CtXURDAb+CWVR1OnTxqUbPFJPHfV+pNb3UNYOFuFI2b1v5v28mDExjWYfazxYb
m3R00IvraaNb5YYhwOaGHclAzx3BEvWMqih0Zc2pq83X+hIF8E/SqeJ+AOTvwdCH
+CBhjgzu7b9SMkz/gPtmpwF7RYeK9IYlQksCaGbRfQAy56m7BkLkFvDDh16G1MoR
p6guIwyz9UV71rBnyg0BCHlEPkvAXUxvrfEdRFEEHOQsPFBenJK5AGkRzkFA+p4Q
Izkso2HKqZKOn9VtOoveUYJhBXJlJjDf3q4NzqWbl2nSC1dB2RlrOiWrV8DtKZu1
U+O4sY+hbAK2Pp5o2XDKEq/UxU0luErJON/WBYyXh4Fq1shfo1EDSSnIwHhB9vRO
LtJDD/QRUdFwPOjfvNK1iMttJW9qZPhF0dAxyfuf8B3iPhKxGUivLgTFjZk1o0CR
IpKk0gTEg+OKK/TOj93OMZiJ9rOdhPyn0+p4eFaBE4WxRPuRvn3PZrhi84ZTvd1A
wTaCixXVdatNfQMjAXBKte0aW2jmsX93cAco/OfD8PZOj9E4EPABTpFldEFlO2gz
1DvurI1d2g+TB3oN9zdn357p3QFg+UyP8XU0uMIGKu6D6R8P/0jpRlJYyTUn0Zg5
BQl6Bw07jldGrfHzGJOU8eEQVY4VRYFVgytuWBSgA/sZ7HF8P2XA58dA9YUrvlFC
ACJJMMImlLB0wapPHMpU9BKTE50ijgzbOQpjLnYZ+LzUwbXY/TPIf3Dw2GCuoGLK
OB3cavQo0uG2vLzqD7niYWUkRRcaPI3spewkqTnTt8LZdN0J34xKzdpaIPoD489v
c54nnnAkP2RiuPLfDlJ599kq/zp1T1h8GxLH0vIMgIqR5u4q0vkaSfXO/4vxUqmY
xQCL++Ke22yzcHabN86YCA1kIbTHHPVI4uK9W8ZZSIRMG0oHMvswDjNqU0KIubBV
XJg6Zaw1A9e9Xx+X2qhwXDuFn0xlrnqkUDM06vneV4uXh3OVpFc11LIVHvanPWu2
Z9SCnYZytX7IKcIR2LwLrHeyqcgBKITl4KGEAS1ZFsRC+tKoFDTPTa4dxcM8BXwX
F3T9t2ZJp/3OIuExw+wneRdb76fv5CFAb7PKdUrGABtnvRLJxLcXAIU3D1TjwYbO
GUyGbV7DR0xQe48eP3nZA0Mqvyfljm+rv/H3sFbdFZ+7C+YrpcwifdQ+z7eFe8dk
GqZMiYTjYFd5iMLiW69YdN1oC818drw4JXzrJb/Fp8BvBzbmFwLnb7orlRGhZ+D1
CKToXLNzegyk+y9xKtC96/EPEHfmBPrPyxGnfvnEoK5aznFXkdOWtcugyXl0zF49
sR7J+WWoMClxfTbcnc9WGdKsFElJEDxb6ofHDTgTFKPrgxxlgx/Uy45eHNK6zQHu
EBz4cQkL8gMj/pRKoH7k8tlvHtR0L6qAE+JCyukjUxT+EKDLcbvuP6nwZLa5MdRT
ETAr9/+wJy7GTpXgsUnCUmbVmukEAT8VueujON1IIWnE1zZ2aErNzlJjMaJ4JU8H
wPtcqNZ85SsW45hppixAR6VF2oRY0ugTcEsqQtHMT3zyK4qfBKhAOB0rbT8MszPj
pTybrPSryHpUPimC2Xx+L/2ElA98VMfaxIUfBJmW67tJDn6nlXbgjEwms2Fvz5Rt
oL/R1AuZyT9MgULky29pLB4VQGhJLtjKwY/S3+rldgUlYRr/r45SAoWBnK5Xhyrg
j7C++nKzzeO5xpt0OtXtSuAAdQC9hFfporHxRS4mzCnM/fFQXlWYjmT+bY0p9uMD
oZ4zRE9vU19AAG6OJKdgMmqBlTRf5dtf/4/H4aZpN5DBF+Pwz9o1l/BOhYMPngUA
QAVDgxiwuiPn4Gxve7t5JQfI/4QIZMCXY+Dz94ifMiTtL9kwL1WOqB6dwthf2GKg
KQQLqWXSNFvHF6aNvS52EBpeairvPuwcJO4Etcp6IGE+RegWyMII6zN4wLvhvVzK
aJoub0e4noyEMW1s47cGXYESiz3u2yaDBn4aWXO2PStRo2YJDZzJQBAt65dROAIe
GAf0geGLAUzl9noZLkSVw6W3OKh1FVas2WwGthoGP4Rur9QULlMhfWGsJL4BPodY
5ePYi0JIQ8VwFmf+Sdb9KaWrCJOvlbj6mBT7e+fJPLcC8pZn3Q//LDemFXg1nYQQ
f9NuopRvMSEPsYgoIO0eM6NZJpEKMgqd3YSL1bnbog8czG4AxR5WLr7ZhYi7FR9P
XEwFDwAM0oftFt/CjqDqtcJelGQSAoFgAe9RWZ4KVZ7YRTN1RSUob++dIqrs7Vth
AK7RqAxx71i5NUa8bpsuTDsC8zvoWlCI+If6S4PuEbKEBcAmzK0XhXVgCouOzLBk
4M8+ovF8POxJK+ykJEl0Mzw6hZpI8I2yg0aLTmLxHhIQzHVZkmtghGQQGQesL1aX
/MMuG/Nh1qcFeOpmzn7xdpGnYRI7rbOY9TxijllH7tWSWSe+2H6ZmXTeIA9QNyhS
SgZFIQGCsUY8jsT1qbiWeoB21D31pY9IElF0AIlwysMgocW0dOyqZ8IT3cHzoehL
sKxQl4CXqD+HzW4/CubT0lxirfk3YihlLG/xhjRA0PbTWY37G7ZS6PWEe93tJVm2
CczW2x8R3LryqZtqC24IJjt/SrbntFfrdkDNvzw4dVezeFI2wwLvuHocA2B9gYXH
ZY5rzqz3D+t6ehSVZpDKmZHPxQ6SDxLmly0iN0qp0BaJDILOco3NEuumyTpUWAkL
5wxyHVueO7QIijxYQusiq0VYMvaeg+mNDVS/P1prfCZpZvhG+PW3CH5UIlgAUkNT
4Hayo1LphPOr0+toYJXIKGeXjyEL7Yz53yBtnLiy7G2ogqHwIlQjRzRYKhximLSe
I/u6uYBDtuLZr8c8jEZFqtAFBSV5pIomVPBYETmNQtIu9E8xQ1kSP/Ef0de4qf4P
IWhqTV7FTxWSQVf8O4RjftkTNlATvj3e7pQd7wGRIQ/JZ+OycM1YSHYfqbYe80RS
8vUgoux/x0OJ7vAyK33R8LXBPT5dx1asUwJVrURyku+nR/b/Req/vp6OzCMpYnOo
7YJroliwJqw8rFGTkNUw1tSpp02skhduyJNQVIe4P+U968E6UiWtGn80HhBeNrWR
qUjn9A0Hs+BzIE0yoqAua/ieFlBWdyr4t/iA0UTEVTisXpH93bGeOEla5KFGTUvk
Xoyqq2JcziCAdPN+dGAeYjOxSC1JB0SgZQE44EQkb7v5YfBWeD9dLxp/PGULbWRs
R/i/0VNB5T+n/R2LKICRkteDif0PTrJ6KoBknfzGYVjFOjxt7gFFnu1ECwapH5ws
QuaRL7eq7GEg+VKmf1vvK6Wzhvh0M8JUYi6Z7F06eh3A9P4atqrtIe3/J/lZdSht
uZOy1W1NtbfWaSgE7HmpUOl8/bigj4smc1qUuH9+Mrvg9b82cUWTWnCkNULf4FXL
nEmfD65FOIXTmQVYgCezrsGp4Bsxvp1oTq7607WE/OPwd3crWktmHy5rVBVLr2Vu
Mm0s9x5PQ9Mdz3YpVKD6xoMdu1pwC0doSf8EdpFcrv2u0TLYHRWEATte5D2SkA20
jZO5rPULJPkIRqgd4AoPf7PC9yzjhH9yah8LCZqUDoUqGYEB7f5P3Tp/tYp6nuIQ
m9EaoHB+7/lDswlNZ9SZaA0bJ3D9xeFUoRPeFjGeZ9ymCUordoJDGjpCuOYm/ngI
mLvnIhmeHjsCiLGbmsmkRjCF1xrhLpCouzKAq8KXNstZgoiTncHe/cL5VSHG46Qd
W1aFRII2qHWHnUElKrk16/assTG6CBBXu3oXnDthb6pwDn46g6z4ZEsrIiZM7zbf
elvI1zmZVQK4uuxhj3bMXBlCpRSyn/Mt4Sv5Z5BvYz49iy2QzJIKi0no6E85KSri
1F+rZB9RMYgTMRu7xm8IPgy2Pxd91Lq49SBOPBqFoxosZy9G1sMseYmP/nccqP3M
RNpRFh3NTvpOcc4zwSh7w8VQweByV+BhjtDSWG4nYjxxyFqy5vV6gXf8HSJNnKb5
3HF+6xp7NoZG8DjevV1hpDxEMJtnhqlbYKOdaUZwq/BixUvZ8M96bDhYuEQXr8y1
J6PT6pDopY3N3oZWNS1X+Xa5K46f+maQfrt+evbb8wq1dxGvdzRKiI8L93xyvKZx
k4/hKli+/3GKMrHuMcr7Q+votvePAAV/O/SksRvnrKJrQRLdLgon3nvnLAIv/unv
cj1QlqPCRIttDTvGRBX/0EA9MvnnoKtcys8Gx7LArnFsZyH66hSVNei+NphkwH0Z
lte1dplmv9f+8YSVq8hCsfbeCY+/eRSOIrcoFWb9YSD5jwh/FIKu5ZCAkxxMCGbB
7/TgIkt47b7oIVsym7ah2p+FdEuhH1ZzS4h/fazkfhoLsA/4VqgpfhnCm9tW1zRa
2giUFx6Ib0jy6S0Gu3Lnv6kPo0jrOKSc1/kbNb/Y+D8Z2o0NoQMV0d+J+on/XPbi
gLT+tlueE48hOZTppQA8cT8WhNF1dNp1CcA+Yjf333Z3WWk6jL5qV/+mCtTPKkPP
9ElPQ5mQct1Awc6a2cKNLfJhVlDBCzfMmbdM44gohAwf0jsT6G8y1WLKz8uzJkr/
4K310gl5uxHvIxS41Q9CFyslpMMNaSiuv3AvrZ0XXO6tKICVzs90qPWGnD2ZeW5B
zcE7S5Z8rq+vbKYSmTQ5xhFKgjdflucRLPaxTcQpCoEyYlbP44M/iDuH7/DsUMOn
2jfQvsYz5p3+nU3NPDCQLLtZ7Mn6uZUICYmZhnp3htrBx6dV63iptRXNaUIuyDD6
4vnxvtjRtx/eguoeP72pYGwvzh4bFoKeRF06FbdYQPu5XRBaOfpXJVzcTMGgH5Ks
UbuQr4Eq/7DM/Qletw61SbblSqV3vCT9Dcimk8CxDHXSFXMYwWnEDSka1PKT10CK
dmxqs6cG2KPYAAH0+FxxZN7Nw/xt5zAPwBKss6qTNfU683vKcaP73E/vbffgRGxv
+UqTSV1YJ/yy+AFW0Ii2sTMfnpruJtM6OZeyvVAV/PotQDk59jntLRvnqj0Zywcl
OwVlk6No1WrmtPQMxE4drsS1YV2JGu5IF49spa2wxC3i2sWN1R1Z70z/uO3CgYGE
BRhyVc3Foe+FTJopZrtnjsuZUEeFGaC9W+6TI7lvaAybSu0Uq7rAGg8h8/eUCfrr
ZiK+Y21phLM6vMwtObPld1+VtRnjZdSjjRsjeTqDQYaAMhPxpNaf0YIwLK7577V9
BtsNPUO2RsIJuX/u/Ugqm4RcFxoGiuC5WNsPQoyNsJ7/E8V4AUgLv+qh8pddtBYl
XtgBFNnEhPIv+Ss2lb44D8nRWguUob6h9rvep9/j4+SUZ3HjRyWG9cu+rGgBnilo
y/Ix/OMze94Yt4L37/Zusc5vSq8shEMvEdugjZoGlkfY5wNjeSC7hj0fDY5CiKf7
9I6rZ3IOGYmSsWQ+mm4/EagPR4YV4D1Arfs93Ph2KdDhcJmq649ALbDREAvEYzJR
w0vBOuul9vbLbookiAHmHKGRYatuafoR+DpoX55Mh9V3/Pt07r2TWGyCG5khGTU5
o5bBwNtx1Z3lEML1QrNdL/V+LDssnGZxLpQ+fbk63CcSKx1QPji4+FciY7VHxGND
ew2pIeptjmiNyquI42xyayrl48xUhUm0yLBxADSHHHZpEO6Op4MyAzLjk0z69+w2
tikJQg4L8+tgZI+T2HwY2ofC7fk+acLacU4vfPLnFrFWM0cMPPdeXGpMcCwkcGjZ
X/0zY+bJhavClKwFy0Qbljc8C03eG+T4SR8YxARUzrEz1iUw7qT+cSymZACnrzJy
uD/HuHNsqB6ueiMeORBf4b2/8FcW3xbZdRgCgAHX2rbnKqNa3dZIjC1rnib5LDtu
O9SDY595czO4QdVIQUISf6GqwMKxpszJVLkj8nQYjIJqOfTFo+G8+NMS/3OK/fD/
4rNZF2sydb3+7ScUQ5J3axF4I+ZqxD1ZBlKqRFDexRRf//6ssBLkarfysuSFNv+d
VVl2ktpIrsIGwHU9DEXw1ZWK81VLg0tDI1ixy61Ngf0fZRRtF+e+jqAHDHM/chYB
eyUAepE05qubS5eB/ycgpW9AHd07xR+bpdaR7b+DSxBAX7U5bqYwxyyNIlx2zPFc
S4RhaFJlrkNSF5xaNbhGgHNO0gZpxJeusQKCfUpj/vv66giSg2H7RttwhNMQDfT/
Q1MmOYvwY8ion7E43RyEB39lGdIVEOJ9eKT9HWoVLe4h4kRzxmX5i8dcYixcmLQv
ICJNuM7h4s77tXDi65PEuS5IlZUkJ1XmzFjY/JvqJ8Gz2lFFbxH3Z5+8xSNIct+/
O0o5DEVagpXzEAMp0yEsukj8kXlOMrDojnUgk0/IiY8xvU+arM2JCecObMddbEk0
SOawyt6UB0/4vwO6ZnBRf1Jrff7hII+UIFMTW1tIBpyeITfeIlAgaAlizW7o2omd
1IKIF0Ar3kLWFT4Kgyhlg6kOOtSZLIyvIWGIz1Q8uoExHmhuqe1nNYeoV5dZkSFl
fRkKaIEXpTwBlT+dSDkB2/7WSwTzy1pxChd+vSdazmt2QsMrclxofgX7HPMdTAxx
XzIgl3Y7NhE5FAd6S6KqpHlmQ61oZYfcyMPnQvF+EVZ/+KYZQZHY+dU+vmBuqvBe
0jdJxywqtkXd1nh90g8PO4iBZdA7GK7h4leA7Znw07Cp7iedW3BbkK3iuUdJBHho
rn70K8B19ecG8UgBFOYvt39m1L1oUTvn3P/CwEIBTOVtpaTamGVgnDhQsDHAD8Yi
9dD/3zE+DulySQ4I746E5/UlD69Jvrj189NGB+/WAaz7ebJf5EqP8l15QIfxQRGY
lVylL1dLu2/K+yWvx1/oG+yYAXjLOX4+GxvUgyx+tRNa/VQTlrv/grWN1V3JKs3d
q3tIj5+QMrbNNBP+XWjc8Vm4bNG/2EJTt+c0yQMAev64qzZPJK55/yx7qbpjUulp
l5SDX6mMSV9b100/Hf5FPLteJ0dTRRdeo3BPUSz6t07zqDQe2ThwO0y7bEvhR8AN
SJqijXsFTlsKqFKS1g1azKoyZ1eAiSTIuydcGwyCm3hpeee3+jxMAx9ZL3utWkX/
kj1Hkh0zAjUYAwepHria7ogEdLyTeDajF/4+TsFCyQ8zDLsCfZIkbHhNliWwURHR
u9L77M0WyKBJ/hdKLhP6ai48dHiqYEnVHCGT9QfNJUUDOqfhX6HNcEvBiABJcX4g
OVvTkJ8NSNzEfaGNItidXoq6gAwtDE3P0U2HsuTEOAjfITVPzBtIrG55KEhjPMbH
ytvpfqa0gvoGdB/zdF8rnfkiUIvgyhZeVoAbcwX7XVKsmyktKxolCoMS0iYxoreL
ouw7VmMCF2SjeNS0ewX02XnjuWAsyZzkIZCX/eF1D6+BmlSH/4UqTkooG3EuIkaj
vubLN280+K2Ua9E3WNbwuIajupAOnpDa4a2oTjCYTVZyUMT09GEN51RLTaGehOrx
SVTd4dVliNf6GaKDy07c5POu3INsgI0pPCLKkbjMFyAV4bSiml0D5eM6wbNHR471
p2Fvzb6NPoFEQewezO+qOstnXrXCRyoLlQd23WYmip1YP/lNklxXJDkIJA/nXvJF
ZjF5UsFfLh7IBI6EcX89RLmI6Cr4hebUzm0zFOU14a8gZVSxg7oU+tb4jekVCCDt
sUcHhIhEiCvnyh0yJfbAoN9gCEcvA0xzpPVV16txNYPsHXJJxfK6+ihuyTWLeY7j
0YF2Akbym6RD9XiT34O35GkPq285Vool170IqhfwyydIYS22qsX5aP2WI0OoeIvD
SoXV+20WEYY6JG9YsMB7vbvZDcc45vThZe/31mLfsloqirvj41TvevFtaZs2QV1d
HqIp25ymfGqJRkx6i4bxlkl//lgbfVqsjF4QkUF/FZIeO60l2ywf58zZFiHDrNhj
yNJqlldz/sbGpXK6do/zGt2RwKIbqJDX6FDLf1vqzM9c3YFCkARwSMwjGZfIAjL7
7HJyBkgPOC0QjBaKQE5OjRYXli8sUY2Jq9BYxSmzHnYSm/vv15d9A80eBMf/cMJt
8ORatFlBO6qVKD8krckx7Lnnmqlg7Rgw9OHxYsw1asq05+XV6MbL6gErdWdFKOGo
tTCYVuSEbqmiuUe+j96PSa77u/DcbAJzrhjVLS7u74l5itIdBnY/WaGBBmUmxhlH
G+lwvOKqmhWs0YO1ufffpmPQPMie5s8FU4WzC9U+RorlzrAurHpw9LwbBCJxMyM9
7LHlfAWxiPmaLelgr+SKzcuQWsrEKCpPap8q/OItyJ4gp8cu3V8zXXmH3Bpx/e8D
CiBxKBDVK/G7FzJDF6OqoA6vInnfYKM232cpFVehx98aWnhns99Qk1nmhUzfos/w
zdasCOvG6YpnXLwCBxuS2awafm4+a4bolyqiB3m4w2dCY8X+jWA4qV0R5sNxZ6aa
lXR33HpqvieAc8i+e+GcCKwoUowz1mF5HV5vwQTSIk3I1nCQ/CSHdbsZ5axFNs6O
hnwQq/7ljIgkwT/MTkruuksrDRc6MqMBvO+ZrMvUTYre2qBINJ4JxhP3CAKuP+Aq
PeUNBEdRBs/mPZ2uqHLl0S1kVdrTuzNLVxF3GSLTNbpFVPGwBVE748QltPYmIpfG
bYyg/+lpjJR0bnM3e9j7BGvqdf+J8fsBmwiaWc5fLFx+ASDtyI0X8uruSwKpd4BY
S74zaQ59plHgA8Y7J+pIznjd91PWV/IgiYCiA4kuydgw3rKvES2Jhyz1n1buSkzF
QPCWlrASn6yMsIEZga/P49jCO65LyrTqf4ANxVuWBe2DIJW4/EbpJ7HD7oIlc/Sw
R3Gpt3VPTYdFJhMt4JOuEZ1LmmqmXwy/4TVujbdHoRdKDY1FGmYWb+wQTcyfyJy9
2KR4m6eaZjPdNfvblwQDh2+BEbu8kvKMEMekFgjSiKmYS6ZfNl5UlPhrzK02ec41
yWKWfEBXhpfQ38dXc+tKMyviF9eqQtU8Xioq3a9AHsLOHteOkIzbVxFSmdDecp2Y
/rQ6OE5ln6SXNe/rgHAlGHfZtdg1bDkvaw82gH9X3ec1RX2zcyYQIQ4nrUfKMFZu
YivYwfiPE0ZaCMrbudAGBbdBi/gAMIaJLYcSn01FLnWlDZHc4uGyITlMPIKGQ5zp
/D9l4UVQhe5ouuC/mN9dpfyuLyFbUeNDqZeMmx1ubEcLaTvEb/CLN/PO5dBa2gB+
bVfB0Drt28lHVqu2xK3qJTNgmGbqStvcN2YQZ9kWLSwLKe6wFQ2te5ReaCvAcdWU
wfHMhCKjg0o6F/l3sE9e9ocTLrEBc4AlVK/8FCmwToykJA0ruHNcwzxTKDVfbCip
vO3Odd/4ALYrH8kn7oHicyttj1MS9I+6JM5TlVgxI0oIn1KJ7T3t+PmFKGr2ArLy
B7Al5+HoFkEsAy2I5e+pC/NEWsWEQUlDdqAGT8yfmAHTbndxLSB1qGC943ZZ0plu
znP7OKxxbGhG1clP3Yw1dQKjD+FHDQL271YB31nxzalEYLmOIsj1iooY7yG/ovr3
PxAY4ySZ0ygXanUrPyyBVeuUSevV5iXsK2E6xpHj21kYRt4MFT18QHdAc2V5ifXv
fE+VIUNU1JXFY0y4uel/vgLuTwavWpCRfHMEb1UVjji1VlXnkWpxQDNrJeNDTrjx
jJGTONPrsjTjxl3PK0ALInPZSHKCaL+cs+UpRDMkZojtgw/mvgmflW0TWVr2S/bU
amF+FXrsCRq3ri85cLuey+hrRuzIKq7k1wWuIZbUSbGHLW6d4a1bp47WlRRh+Ke4
vMCyWEw3yIJTVHE1eF+TKf6ZEs8z6t/FQK/dulEcgxjv/7MIdeqqZS0PLdPfuBad
PPrXPs+WNAINnT7wSOxzgWUITDPBGjY+tg1T/MnrXaOqwmtXNlDiG6qG+XhWyB8i
EQROiWIslLquMZwke8HcGoKnVZgKsZWtfcJLBJEdjh6lu57Rx0TGqSPXx70zXnyU
H65lqDTnMcjW3if39B7X15Nna69Ti+bBMUnhzqWTRXmJnXIRV0PxdcNca9yqdodY
nOciB8VGiHkGQn8uEcyKP9sdHruanfn+zDpV87/6eVjC8R3tUsV3Fyj7rM7o04+H
HdOhakQEP+1/utYRqg8DWyE61/C3UZFQGIGrr7F2YgIUBOkByRIN1WnpoKe9PHJL
D3q3O3wxrPqBkNdwln6obYdzVJgS0Xf0o4dMwXYs7k3UZZPdA2QJHSp/uEVJxDGZ
MTkCNq7xjpU3bbarRrEohHByGjI6u99BkYxHfH8WRxC4hSocV2KsR0GYc+O1Yt8B
FXEb4dAMhBHWr6iMSJ8HPgvVdP4eK3ARdxFijdftujgV0bC4xQCIclOVcyHoXMBw
gZi9KlLhW7B13KKY61D3abfslETXMR+P56H+6MJvke0MksQO0io88u8wKO+p7R1z
q3ccbtXw9CAT0LRPPWyGVEbOPJrT60pIfXgae7B7r3Xn7nPW57G6LM4BW+sx7/d4
HsliLmeWMBftybrbjY1PlPYIwM7Naxe5VHM663opnhdnVoNCzBUBffb2wRQoqsvW
B6chKY6hnqbjD1CxGuL0xn7Hn+fW901sW1CLpb5LSrNQTOXQp5UK/zsrE6s63U4i
99r9vxQniZBDMwi36RVgIA5edbUmWVnutOi6rzJ3y42LY1tpusPVGjE9aSMKbwPq
r22hwSOYeV2MmPHNzGQA/OFK9NvvO9R56mpIjSxX6OJJIh/mMlwjiPAJdrTz61g9
qcTgKqpg7+feqeAcfIi2v4SqNQ3OZ+TLuruEW70N586W30p+Ij3RaRt8rdpAyh6Y
bOy688LjeVdb+9F5C0DeTKlvtcoNWZxqvztMxgc4VxMmAAGjQrN7IvCzVK01dLZJ
pa1HPhXp5LSL7yOm9B2ragb9Rtnh3zTNKjaO6qCh5m/3aEjU5wPu5I5w6Hzryuas
vo/e66g+EBdb5wBj0AXkapCW3f4rfqNs4fNnFtG0z6IFrEl+f4bidEqBzNb7UGWn
RWbisH5nfSBe2mpySEIyWKbg5/PbVfYj5JgwYD/Cqdf7Zzzosoc1KNN5gVfcZsE0
zsgXN9h3dQpddLdDC7yhkwUfYmH3RhWtWshrIZH74cWPS2sZxfE9U4AF/4QjMDk+
30Tbpew40CquuYfJV3y3EoX4b/OHXuABUHDHfhJcY0/wOPJsENXXbrQ57g7p5QkY
FIxvehGP3AF8ZP/cNV1uFcsfChPygfUgphmhvO2emgcveSxNQVM3OgDz5K+o7iiO
68qso0l1Jrt2dOUb3PQzHnQmJ0D9mtinTJf8AW1OitsgS6rQjJP1CEueFMsTh1yk
Xb+/k9Y5ZnKEPiDbslLHq8pnU2ye0sjh9BPpO6fXnE1SWLcdJT6QTpY0cB1TS4AK
h/ipjYnW8Cxpcc1jXEZBg39TkSoeEaiy2pXbRjrAT/nWf1aPZdstA37p6nO4QpF0
qaOTTvjp59C6Si0AxxBNC1/X9PR9q90lHrHqtZE2M+QBiN12ct5aPkOIzZRXzoih
s8DRvvtQteAwdjLfNwFPN0tLKHbyXhbPrXAFKiHYZmAHkdRhfN3LSfrWaeVo77dB
5hBsAkTj78eJVvrZoEXgq5/2gdDZUgMZcGoGh4i6KjBz+YErV980tBmahfTX6G8u
9+eZZYhknUlYPO9D+4IZKRde54DIKwMIQfxz+M71e4eCrwkL0sbduqk68G94Q5s2
7hohDKV1LzGbF+c7JDGVdCyn85k783M/46CTl10G/ilgDhzMaI3Oe+Ck4VMOuAiK
YHiGM3KtXbexvi6zcJEANP4mHARb1CVaiXsRPJ+VM0bKSgwgkwMwueLgUUX50JX/
YT79P04/8bC0vX2X9pzadvt/KbamyUZz14kFceO56BcIlcVzHgO75m061DibcyvM
kLVBZ/XG14Qh3kTXW/07oi4assqQb60IjWpYSy3nDIIOVClWu7x0bPh5JNx5gMCs
dXio7OQMd5RtGmSioyqiHvbSEwgdzqHyZyYWG1s/f+UdtwQuDgfh+jBGCexFe68O
aXv0ESQGg/0i//dlIsHPXtK81oR5908AZwjut2XK78/r0X7R+0ggrvcK6Km8rIbj
qstTx4QlArlQAZSt78gb9X4DyB+QPY8yhHZejmFGlN9hY2DNhrAQc8D1A4TQWPQn
eoUNfyLsv1Iu4NM4ypIP1P3qEJeH2AnOnfCbLK+aDszlqomFLb6P7b72/6f8mYNv
2pkbkaGSLDGVXx+OMHGZKQ4S3+JQrzb5kFSllLLquQ4t4O58I2Hqv+eKi86sRLTx
ZxuPH1vczGaqQcaitPH8sCAI9enb1umlgWtw1xsxDklfdHl8VGyqchCQqZKumg17
bhxjXqhyiDmZIFw4ZOvkE3E/yO+ZRvZI+7ACjwpoB5fvgBXxvYhLN+GeWh4nSACl
cLMXsghoMZBr1UWwsreFakbgAcCt2YmeLsDBggVkasY5zYzf1D5EvyhnABwVsI6B
CBUHK4CAgUhHEgdmYoigTRj3mYeD1ha7+JQ/KCMiDW8EONgUyDUrYpXXCqPwC7B4
X6C1mM0etN7/+Ag0c3oXG8ph/gZv4gEHX5lQ9dATNtRhhrvWTO9xPWjFnPzZb8bp
2IMXZ3U3T5L9OO9Tb3C3aKfTgpxpSkBGcf4gxXCtenYBajdv82KeSt85Rm+eAbKc
JFWFJV08vxdZjkDWxp0pwj82e/a9sjoxBlke0Ui+u1Hva2/lKHcn29lK7Yh2z/M4
w+pbdgyFrgs02s5radtWjJVlWnBlOwVwqiY0z74sQqvSgWuOvH6n/Br9xiHjpt+0
o9Bwk/d7UEKWUPj8ayMCEBewkCH/1cbIo0+YFIE6h2eygYn+uDlO02dIR7PBGN4c
8EdOgT0yanPhTOKMGlLwZe6ajrBcizdmIoFoj7Ij2y5RoQDyG9hLpoD3meVkFISr
VZuzKT2z1ZXrVqfWezPe7hNmqIrS5xqefMnODs4UrCHFV7lXvFU/MXDHpI2eyMsK
eKxnZU01PkrRtoBbME29lsp3BIUttNmH0KvlGu5ulGkFvq8uzr2Plwa23M6lfYtO
5w6wK4xuj+u+2OkgtCij2O82ED0kWUecqqePMGYj6FO3kz4b8NXlgPV7iVMjCW5Z
1anrDMIVE/AvOXNXQhBc/GS04JkuOStjgG8t4E3JjVMMGFgl2lHGByPsZVsp/+oD
6bc9bqO1/SMi3t1ZvRU2mqTkErCpjijGw4RTDm29nVLgQvoK+csaeDEAg5WKwgHg
+TF0i7pLNTdztIU6JaeB9dXevdChjG81Ym/Jm35mXuUBIeC8mS/afnYq3QCd08OG
lM06MOFw9CJv0+WmLHhACbxTO4A9GY3+dXsvaWTF/p8waRZeWp+l/BENM+jbmvcp
OorjGAMrlxAg1m1XVAiYoP9/cJoltJ8BGup/uVGEmljwlx2SaqUOaLGoTa/m4UGA
Nvk8P0ZDL3EqbbhQAMnyG/0WlZVoR3HYETyB71JQpzLcN2V4s7yHzrmWUS5hk1J+
KFxtYi7NqT/t0L3o7RpXCnpdqocyri8NeZl7w3aN4LEoqzU2dbVLyj3kUxFKYN0M
mbL/As7ssgt6RYyWFO0JlHHmHtuSMi/MPhe/8AReLWxfAcV0Z9Php1gl1HKtc+P3
5ioi7T6GbCfKzGtrrTrvO6gd/qQ30wkgpZCsKW+uV26QT6yk5HmExK9zTFOBJwTC
+3v5zh/ArZCmprN5fuRZ1RrzQqv3ygicNenUdIdWL3bvTjsThnAd35lFBs1z9tKi
38B9EzwpyauHDuf/ZSHKTd5nXiCrBIhy0cIdylaRH9CPpinQ6z8wxmBj2PK5EQg1
AEVIaNXm9i2rbhqXJdwjQz9yVpaa+WrpTnOASRUac4fK12iRU8C+ySLrVlW9DNiH
iJq5+PU+anlys+0zytibhtBaUC5+H7rFk5yTWGUc9uOalZ9bxt1xVwdFHMV66GVA
d7zcroVB6E/6TTR7DGwL+YfC7ctygQiwKjDAzbiial2zcOAYIqUXLn7YuEqolsy2
64S6tVDxDB788kz2ElIoBhbDkLP7AEFf46kz3sk6pS09Bz+ktqFjlnxOQVwPXh6V
Qk3Mz23RODWtMv8NAlDrgqUjnKI/8wwfamyBdZot+bSTK7tijH3VBjfXwxPRQK93
FmbZeMFxi9gRh03sTmL31XuqXh2Dbo7P3W6hXhQ3Gw07helJDIFrOMwEMm/pcLIL
9SnKYmGb1mfsmgp8+MVkCGFcrixSmSCqCWTKge3JHOWuqDSS6ZrONhP++Tw0kpXm
A3SjGuhjAt/aqXgqjWsjyt6zqTVFS0DxRoM+/SDXRO9dZS0xPSD5zZphb2m3gdhv
K0FsBr6VvA890H28us4uc4tAslT73kgnSAgZAe/kFcdB2UGBKy6HpLsb8qVg9aGz
myfTYG6bdnxBoBK4iSRU3sBunTS32GE2sFKWPs+mmGxi8vj1Nzxn21I+7ji1F8wn
YmqWePp9F9bWN4uyx39cJEDCLpJ8BGT6VQoszcpTkDg4OKw2KWFFmSWAYW/kJqzG
zsLer6ZkOEghG4VzGWl7fj31jxnaNoCvNrl6X0FxA4b5N4Mx4pR6XccritXYQQl6
t0gyQP4N/7tp27N+jRx2VyavwKlNYT6qFrfr7dz+yKtDRV55prMveeq9CjwqBuIO
02NcwcgeHq3PrOOzSg8MMmnQZhZzBniq3QtnfSG0Gth5G6UaJM1P5OwJWAlF1rXk
JMltUldtvrFWllh2oE10bERgMP34uXKpdhS9Vp8wKBr/UepgTZFORDuff1HYXkGX
ujkluNukVhtj/H+Y7SFz2xJ35S9Z5ue0rLltsxy0HVVu5l7UDrVG0sVlIf7O5DTs
cEFNZUUaRUJzHtWoyF/U4Ao1ZCgAZ0YSW3WGDhOId7lrvpj2bOdQpClpZqG+iagU
xl+j5vsI/JoOafTsVZ7zqRudnFPOie7OhTCYMWvVq0anGz4nIvmworHrApmOJ7/B
/k8WlnsSsX0/FeT3BJBdJjGfbBMuM8ZegFaoQo0UUsQeYviHeHOyCVsPp9MSiNbM
ulk9d8+BqU5k2VNTaf2YOXndlux/rMN39kR4zi5kE5u9FQUcBC4Y+9tQtLIkC8LE
9lexjyfn8wofBE4eDBQH46j0o7b3hJu2qXw1M3ObudEEjP/NkLPOcS3B7qMEijc8
TLSuZ6Kn6OiHXOPfdOlDAHz9K1pCpSuMoEWTQTogRvXDo2aucjyjNrLkNht7MwAM
RpNHccK9X7jqOXMnPLeXFTqsT3gM+xphH0dnkaaGPPWh0T8uAfdK9x3PSVgjkkH4
KW+hfVs2zVs965WDtxiJrL5+DlccLApEdTXMMXTjtwswKdGy+3vOTgF/uGt6nhgg
K7k8TzJytMii6KpGoaEfHA7cZLGlsM1Fp1X+siozy7oqS487j+PLr5MDsiVQvxKo
oBKQQJOgwc5VNBtV006TJJLIBjigQYOqNPj7dVoYrbChTUdqHOCXe9DG91qIvDUe
RSJ/AceDLERAeI9irwX94XlUNVU4NyfGh4f3OhBgfDDmhkwJBRhjc26s5EAXE2X1
yiycEwA0y1fT7tfoY1tsWYIav3H7dCnbWfFyqpTH4dPF8pGGGppFtg1EZGxBM2LZ
O0pM5u0EH92IVX08m1yna3iFck66KAi3ZUptVSHetGmYiSpm44OSXYgOR6Xlurw1
Xkka5uHGQz4+DcWfAv8zF59viN/xSFeRLwFjwfdFN4LgU3Z8WB8XuIy0OdX6mAyS
0w03D97UR/cG4R6xGJxNySNEa2ydgJ0Q286KCXQ1oP+lAF2u/5ZYdar7LRPryYJu
h/PfxoG5MayfpqyqXDiiE7zmanInxDOPIaYVTVeNOFwA6CoS1orQbtlnFTxP5iVz
KtwV8lz3wyzOks/B/v8F831paCrvzLsw5W4/bAGS+Fsb0BCHPqHEm1VzeK/xnlkb
1KqBG6undWcQAjBVKv2qpTeX862n+vEGqzXNnEMj73bmE3dnooo0cq+ICZekqxIP
BimpOrktx/wtqV1+KB5edZ98EUVkLQ1Iu46W91Qll87oh1RljtB7B3gyhRSRkv9J
xpEl0zWbRLd/8wdtFBqY9qLlWrS4EazCDX7WTe1HF5JdmQC6ghvdA3I71FCqEUig
ncq5KL/+fwwEJ9TtgGUNeTLWFqcFUDI7Y8B/Z8Lx++piickufQ/amM3HZDdFCK9/
juneM0aqKACxIzSvTaRGEAOuS9FXIe16uFdtIGYuVippiHef6eO2KB0HaM/A4Qfs
nYdHsa8dc8ozkCk6YpePc3kAM8t9lrQc/cfdt9lD7B20YJLKEpB3zZkjcEGTKio1
yK79NcAl1gIDiGPm/GHhhh7xZniuBkXHiETJdi/f7prb0kk5dREaGo02erYt8BP0
Z1JNzmb59Qm5WE+dOP4hoA86Ukg/EhTPZ8/9zcUMUgYZ71a8MgRfpT6stAfa93Ko
clQAkL8dOz36/BivzEdTVnLvAcr/zZXfp4j1lZEaUwQ9mSJNhPybsnaxhzsqH8a/
9UTITsYM8Bnf1/z90M/5mhuyNExVdf4DjtGvV26K79sb1X6xUK2E58cEu+pjsFMm
lBcBTRju/4QjYUdcu9vHGHGu1pelmPhB/1lH0PRPPX9ovZBQDoHjB611d0xoy8Vf
uedSo/JQqei8HZW8HgnbUEMez1I9FGdijoU4i78vbclLjmEMtcKn7tghG1bXoAwp
4dRfGMYDouD1VpIXxpIR2iKR5QWKjNEZ5b/h8ubBgpiSLl6avltsWV9Kv+/LCGFu
UGy3uoz6w8c2qOoL0mxFPvsAHTaQtaduc+7pLDFgU7amTfSPiTJKWWkgt/0K3fa7
2pXXM7B+jUjqQZ/EfQSHBaKNJnMCjExzlGSbiIRH4bECjJSK+Tj/7UAzopzQU40o
F42cykm2HE8kjT+2e6BlXMmZqAcBQH4TLNKpaLkWd9FJ9AJDDQhcbjeOws54OYiE
dtV9K5v4hg1RQAys/dhO/w/zbRVGlGGupOrqAIBLIXnSzLA+q7+tjX9g9ULB9DXk
GZT7jPXm08HJPaKipM+Pk9l5Owi4A7uG/cXttg0OSR3HTg/sEXqiKJkQTHw1Y6SN
rqMd/Cxpy/Y7YaxVFxwwOJDFA4sHbWKaNyLKcs5W58Kb0IG0PA459MfsSc8Et92P
3FRtJjkAIsXlQXPsWycevCiicuqt8D4j74iQdwQZxpKGeFIc+PrHWzAtmRdKltB7
/Ot7QN6Zm4nNlTDSg81cubZ3I1IWf0UXPJXmDFVt0pBD5yV8l+vjU2rUXC4wlZg4
MRYM52ymqpyHYdcjp98WkOZTuw6DAi01SpyxiVguSpXv3+7PEwCfQDxIgKLHzvrP
/XJAOJZXbPPwylNr+8MX/TsweBOEjPDFrkqr/w08locuzOH864m3bxw4uY14nGtg
qVAuUz+hIXpwuObjRQ85jsC/1e8jPdPEZJVb5uaQsnu57NC6LFdG6Yxk0nW0j2rd
aNXbjjNnlP8TvUIOvxcHYE+4SrgKG/QQGIrm/Z/ivcHiixhs1XEUfgA1pd8jnorg
H22H+RhgmrZursUgJGjkrQgxvx8Poeiw6YAkE6o06QJj+SXtsMwhOqIzvjwd1LO/
sJ1XzEAbfahd1qgNVxS2CNyWyIloScFcjCDlPfr4ey4wUR8uPRE8UU65ieREYEQr
/eL2vQUcGtVVApqyfavggaooEu6G8uzQh46hOaa1sL07swycUsz4+mlMmEHTBtjt
+cQ8WiazsLFu/xu68O6G7iEslzPdhWHQ9glC1cIekMWvjDa7FbtK30+z1MHb3OTc
My0S8ez9Txq50UvldZozXWOIAuPJ0QKPCi1e7aOBxDrUyNmsTCshjHrQS7hpi5+o
A/E9zWvE87an876rlW8cumA2pQYKLi5uR2ZV8YWaN/qxtxtg6o6P/jlQJqqdLtxC
Fdvm2Fp+iVe9B7/DMngDcxe+CCAaHPNIfX7M7zAW7/EEVUzUdqNjpZwmAcUDR0rM
DZVImjgLGIfBiTLK+/bjU4LCqXxxxS5d9X1nsGcjFypEd3YgSrnivbZoKcQFRpJm
qNshvlLy1/NP6GAkTfcFAyRQwnASsSETjCs6PPm9S+0HaoClrkadYJOGrzft+Ft1
UEN3FidruSYDYy+Xr616BaOL6NHsJRJmvDdjlFaOwU3gz3xDVGBRoWChYrVAVGWd
EeOoJKDnkUI7NAtDqeYZrZG1hKkqk3fwSBij9Yi4jhRHCcNfBlW1105aRD7eHZLs
LwSij+8TRQL/uLvmAZAOSaPi4G3ABhZt8o5G712bTmkCjOuCJz1k/S1WAPaDrBD6
QoftUdWHM2IHnWly7jwrZymDGozsnMwfizDHu/tON5asGMAwtt7h70vk4p7us0gH
8SfuGAHZcVn2dYjUptNQGT1BWuePps1TY4uJExDcAYtIuWDVtI0VJSniwzQIBUe2
gD2APQAE6khcSr2F9+m9ReeZ/zGmcYPlHUUnqafollwAaaCBtLmVL2O0WKnjl9Qr
SsmO1oEBwf0VMqhKR+60Xq49LzBAPHs4HVHcFt6H9E2yR+iFDdpBKLqktLrGa4aP
mKDA0zmqnibe5f6eF25NViuiKVf+Ct8ky25fCt9g+mYqEhLSxFXi5HOtUQcIvizl
bSxBreR0T5Ke8heNeFzvHo/BQ6Svo1kePnwLI3YcWMayPUjfW7KPFf1U2EOYrK3F
LslF3iO652oiopdQhtlUocmzKJgyyxqlok2Gwyyajm/Eq/wMIRRQd/n9YU2mQnr+
f/M80fze2JZNHnMNZlM8DYgLGDC9Z+SSHR3rWdtFNrImx8JW40wZwaL8xEMo4WAO
delzskco2A4RQCn9SLb1iz/n1fLS8A83p/nI7gX+TAse3CyAMpuzzCZ9p5OuVKyc
+9Pyj9ghQmXp7j2mGOZslTv8Iyk3vSjWzQqZysWY/ZKQXjS0Q0iSG32V4ctUqsNs
bjqFKvCTznzBysnRwW/8WqQIDPpahGtkeezxpc0X48meqrJ7fqvFoFRK9RkMZbGX
/FdldwFAxfT5kuZObAbeHmO9uiHrQSQiJGodkHh+240f+sy590CncTY4hLqdf/9X
Qfzre83X4m914NtObN66gvYTpUwyUhW6tqK5RvfzxHvY937nM/DWjbzuUsBNECGx
Io0lyQN6QZmRRt1X1l5zjjrh4Kvvs/PaSt8L5l+CJ9jTHizDoVO1juxeama0om+u
j3M2pHWYEbIfGRhV//IeeqlU9P92FRf4Jm0JkMEoGIemwkoAOEPdB8E5Ioc7UrMn
fTAEM1O8Bpt4jE+rPK2P17wenFTbyMn9ea3a3EpQZZ8asQc1QK/zChyHoN7joLNW
qdEk4hcfvqrk0sJgh5d90oLy6biHP2JvLczbKf6MKezFS+1Mq3NhtTayUcj+/EFQ
r35UFzres//0gBaARdob3U8/FvFtL3Lz5ppTMTIgdhccPxYmgMWr3XfSxDs+BZVW
eyYXceP1iA77Sz6TTMxNUPI2zfe7HLm8utTvJC2DMiUDzfIJwuAUp3xGhRlI1qeU
sy15kKCzjVVp96ZuDG+m/MsLYtrt7+raOKaaMlHQwgY+9VqML1VJ9ycbcqvOCo9V
pA7ch3WbiaXdj1wLDMtXGA6ASsS/6ZQDRYiEGcxoy1opgOoQILVtRwAEPpruDICS
RFKKDXTItxl8k4jCFom4xoIPqN20rKN7Dg3Q0UY9sL6Q7mCn5mMoqrgTiPdCdxk6
5UY1RSwuvxq83oDKsWNjGiaD+0w9XOTw+K/FwinkDbfj4ctebaHFlnuCJQKAlwfc
sspksrCBNl0C4omkF50DvbIMECSyAFpf7J4n/fmxnCWUkNYMzsL5njEq+NO2FXCC
JAK/lmZLBjgr1NL+0YnTn1mTBrsR0GmvxtFA1x7twXYYUBb3hBbXuzKuYMOfzS12
4GhnQ3loRDdlWZ4EHusklkalNa2xaMgylXvzhTgPzR5fk8t7HhFl8PQbP1F4VulY
Er8Ta/nwigtkoHrl2NB5MhfyJShYlGJeOUSDzOA7fI7x3Sk5aoGseaWCGxQnUXQv
zVjRTHy4Td1X0eH85CiidUhvpz6Xgkeh7eRsoxbNNsBUt8fRpyQHpJfMqgQLkgkc
AlLnmZ98FDlTx5TcPlYZzEUCr0IZ7CL9tnD+d3VLfGagkrsggAXgd+MdD8IJbowc
YnAN90XvM2ATaYjBa81IZoe7WbPjvevgEYcrOyIs110zjWIj5WIoRrcazPDHL/9s
AB2yBh2RA2BzEE51+oQZNj+aOcfhKDCN+Fw0y3EoVRTzJMTPjghd/lnJUAQMyDpx
FYcF8iUgGtw/hSdUGQ2dZdnee4o0nQMn7XZNaTjB2TLpuhtRxaNPXdkn2O9r3AYp
R83xta78p3Do2s+akd0XC5IoytBJonEahKzvPMfQxpM33TmkBsQWk7S4C20360Ci
XTXBHXiX+7Xe/LvctyAPX05KoBSsLjWuSxXM2e7XeXQqKj5YOFutZZdy3QndMohz
1/jzEi1Eom68RDYb5kiahPE/UJbSCs1JgpYXqjempck68ChqL22E8yzDHs4AJHoh
aEM6/x9xWneldB8Ojo/YPkmC3DE8laTXqZM+L5GV6Tf+5iXUcDn0QaBAmrPr7QPA
OMDsi37/5wU2CPdLtlWDEXelc6WxQqoCbkOeAr228dsQNkQsdTfLTB1JfO+2MDkt
0evNCghOWtDkqqJd620etuddd+hSULg7c+9HuwWXg8PFjHJvyXhQeoLWWkHKXaFI
a+o4hDTLiEQRgnZX5Yrlx0En8aR1WaFdUALCkQh6YInFG/AssEJSxU8kKx+/AooO
fu4Z54gOcbO+dcrtEJUIIDn61mNaEbH5OLU5LHqKwiv//7e7ZkpnTO6C9v055Iuj
PE/DawWuZWhF6tJiiUdRqzO2kcf1bxgFrPhv06rk0Lh759OMtYuCvc8Qeh9l/gdA
imIU2EjPYad263L+CDJo6H3FU0rMdSHuy4Ot9cv6+qILhoODsnZjVtNNvTUte2sM
2A2JRKAimrlAm6PJjmecaX433sRv3k4i922fDnsDQ77dgUOh4LkKO7fthWKqQw5X
PrQsgBsaQwFvrdiL/A5xhLmhQwz2kQoQlhSobpvPDYuIYIIoXSWlZkJonzjLweXM
icjoiyc3aTMaZyknWKLR87LnRoWcr8qxrWeHiBv5Mcx2jRdUbhiyj93QgjJSkXAo
gmE39CqY3ywrZXkTm718eA61rCPFuGFKHO7UnbMK4ufUuXUolzlC1ejhJSBNJtR6
EMWcSPnh7GI7bUf5xQ+kvHo2Qto9eLwOD+AI80dBB+K/4f4kdMHr241o2mupvQl6
ugFdCRtV3uQdbm5BiI2X0ohxltNb7V0EmCfRjI1Vu0mfbWY/79D37eFRBhKCKKPy
Sc8XAEGE0SDK4RywH7mqFR/aQSvsT+3RharNmbZvwDVYYAf21nQ5SaUk9nZp6xcn
z8Fa6Er/8+HPW9s2xiCtzRp3N1kUbbmMxcPZDRdqWbgcFtN5LgPWgwf5gpaaF2eE
Qs+9eyxmClOq0ZfHhHohH0g33g2mLe0tdhDSIYvCLUfe3c82ddIekmh57vV9QPXm
8E8BhDFU/Ctb9A98oDcG4s2qmLhnmCxZ4Agkke4QorBTizgOcML3Df2Sw5ZUEt0m
CifXZShrWgmJxJLZtUYGAHezW0iE3JrtXTQJrRvGcaqUEiEJmQg4h8dDU0v60qQa
0IdrQRkPe27LUgi4oQqD6BYRTHTzHi1gCCj/11jv1G3/WjBij2/ezCk0LnkQrEr8
4wQJNnaKdcSBb7zYDcFrLRIbFhGqW044OJNAJL7ozBdgIsMBNkQR9BEbDxX6LSPz
dQ0cgibg4Mhy75jBHuCo5vdro4zmOcq3INEim11iaGkv6e+WVkafKKGAZZeKcqqy
Qv5ezd7Hlkh0cqv2YBSCS6Ntgrm6oIYKMurAmnJq53nFVQ+IrlWv6ZW02DiHLk+j
z8nry0R3AhGuxTl8hn1Hp9bguTeFmvNeTwmWa0HkDLa22DhHeDA7N17M0KPHvtPf
ra25FJebePSKRspVg/iMrN6SA1EoB2MYYKzZ1EI3ISVxoaQEihRTAjKkrXym2Dse
RIOwTehRbKRkIAciI1EFyRO9vI4bNUpJyHRXr8rWHdcSX1Pi8r7gq7pjgEJwHvbu
gK6jkObINsWgOBdhvvN6z8slFXss6ErxOqj7+4bq8OdlWVwDgw7LOxmcvS06/jA3
kj/P5fVxRcbmdQsb2JZOUQgr2TUrz9BjTdXV8J1g1sKl2f1JEWUpgh5qZAZmF9Ct
cWfH8ZmfaHEzSBZ2AWTaOCZAbHAZy2dLlQNykG+Nl4qk45cTWfq7ZHqfkjoGhY8Q
PJqHVoZ6PyqBf01wHT/4ZDs/LPBgN3GnfkLqUpdhHnDqUeiTQOYvBqAXYStSiZVI
XGzX1Ot6DvGNJ8kgZ8bMwi9WyE3iZmW9VYxqAKtv+C/wRT7lpXZU8YLOw98gTMIs
7gnRqBzuRzpCQzLiKF6/xeButnbp81LoPnJ1RT9/HzjPcb0CG8TgsChAv39n5Xdd
y3InuuK1fUgT6Wk/Q1nIBtyPiCZDB1H9E88Yo/4S54h/jyu3F/WTCD83q1AOAQmp
f5tTW95NC2GpLSi50FbqdcFZK89rHTTZfOFETNQWmMlg8ojJnZ/Q3WP/ElxgsLhE
3U/FasKuS55Yu53pv2VDTZvc4d0ZIx70gKVX7iKlZJNdt8mLu7BdGB5Ctguy1DNi
hmZ1jah0UZ+lfRDt2XKvgaWrbP312rRMGIIJ+0XcyuDqu2gDDpoAYfyQuuc40UOH
Ru75oBnQaF1Yni0B2AmscMbS81Jbu7TviXL1SyV4mKU0ulX/jGpk5vL+vBL/5Fhe
0krrEkUw8kGZoTXggHS3id867ci+6X18o5bpkD73Xs2/jXbAyhTB+9UFT/OMVZnl
M8UeqG0hvy9DezTAMZJY9TjR6/ohn1mTA0x85MmOehFXumKclHVVQqUifmgAROgi
2FalQugAjn2TR0V0rn34R5xEPvTolqrx96i/2vAIWY040AUjyymtn06KPsBQDXK7
6nFcmwbDlmKxFfxb2yP97mGyoBEC7yA6KHbrkFjXllMVfUXYVszI0IpqXG/Ae6EI
L4/vAyjXSI1TXdsTxMYs6wy/WLQZaShkMdhnQU6Lq2jwgucWGnNVNg0K4BQpkz4k
nNSGQwECnvdNqUsBXwstUoUEcZ3ZJYJKBz23TF3NnKhU8eVXGuKmKd4cpLzEwhoi
eepyXwdlz242A1NcyWnn5CvGmGwwN5NwqG4zG2b7zna8x4GDluY6Ku44iXgaeWYp
TXXqJqhkQ49Xz0AxvNHAWjRMhfoySAs/KEz+mjQ6su1Xyjl9sQVB6JjDtKoyYdqW
NchWMbgc3olI/RbOcnkfP/ZTaj1AsXso4RYPY9j0w80Pf77Vf27N92Puv1dBOTsW
hMk8G/n4b/ges5wB5CBI70rEST/l7m7fTwIYsxsc/lollIZbAzyNCUpqzvUzAFrM
/lt/SmAD+I8y4ouwrC+tDnDeNTwy3w4quomETpeM3h6R3/WrUKBVp0DbJ9s/G6N8
cJ75ikLeP6feDCAepBsbMCh5i9ybtqCyh/Wwv8xyNL6mzr7pRDCz8tnR0dFCScdO
we2P49zkLrUJB6lKk7Jcl0C59ek5l5Y1vquNln+c6zYjkmcXezVLzYARodm1qPCD
qp4FaT0Jyk4RPz9MJyOVhTEyNhuhOPKJ0LP8FwLKQEwrI1/OJeC3od5JautfKwZe
EvS2qq1WrXdC7Vg+LfpWFSc466eO48eBRxXm2NUiUqU9YB64vFxEbPXvbyjZVsvL
WftHyrDhhPVM4UuIkNRzUmNZd4PH1z3KZKwVehvpkMSDnkMMqyoYlwWUm7ra8Txl
fbAmpviGyf6kdq1odMqQO3UiW2T1xzXtLPzj6BCpyp/ZU2YLNOau3VQ5hZkAJGnA
XZJ5iLpZY7SujuVKqjW1km7qrn4pP+x6asZjxHkS+B45gSyeCWlJzdAaCZLyHYzo
KYEcQEvoUDlIrg7wii5hF8YsP4EWQIBT4U5uZ6FIpW94j3LinMGvrvEFSbgoRnCZ
BvHK+qsmTxnpvSaW0ejtQybLZN/K6l0COqU34FazP+nAP91w3h/FXbBz77Gdm25h
KW/CJhsUpr2cziGIq1znb/hQEiEh52Lpdnw1diYul6VTCxJKj16FeV30Is3ywOCc
ZDE6OmfExaNjhtRQph83Ywnk1FxBTNMH1emQ0INEj5oQ995KfOepu1cvYKUwsw3K
9N5Yn5LMFvATyMbKS/jVAnG/kBWZ3As94FjClAFAp64Qu5M8ZYSF62d9tc26Js/C
8SbJcma8mhe5ZyBPVByo3IwwpyB5IPazSgcw3nwk1eps5X6OCsXfjkMpov5mxSd+
aBH9w4GK0VCqQ4vkhRjt7mMhJ4rOiZYwBP5gS7RJriYagtX6ZkcyU0UoeOh0xz5Z
+/+WgOrefzl6A2ii9ywsX11gesw0hjMxS522RrKW6zY1IdSBblMAb9RSH2tpFUt2
7JMXYBan9+7PumvTOLd/AYDESR2wNwL/LG0umPT2o4JvObwAJ767yg3o/J8gMbM5
s7YjZZipnfZu5pyeEbiiphwqsRU2xPPNjchwuo4L3jXCVYBDipIofhBvo/TQk1Bi
GnvDP4SdUFtHumMKOgoSibrackeZQI108rH0TyoL8t6cB6n3uIDYUpfU4tMk5561
LbFvBhFHSP1cCVcc4VFASI2LO9CM5hkfcIzJ54XPBgYIIZuTRe5feCDQ7FzZQKcn
D2K6F/nA0iQhLEa/zbsAU/jPizo28Zu6qkjA6gP3kHNmYrpsciVTs0vvSHtc83L7
SNicOHIk4/6brfK7xmgvIuIxM9WP71RUDnqJHNX+tWTf8hHro2sKi6oEKIuYulbi
pJnz82xr1gDldX669CFU8WpqnHk2+6k3RXkZdsEUDNumnaPSXXAVkqvYAeT+vGrr
biEfY3sgAOwljVC5siUlLqUvfrOCdIyvdVrFJDjtFS1QZ6QaZ6jE8jg4hs19QKMk
gL0i1/PncXYjGmuVQIdvcwZ0NE4gMTXolAbz7iYBXcRppG/wtW7ZS91jsQPqVYmD
R2mQyT0mr5cPmNzA+Ehs3+lY+eg1u6B2GbywIVVHBSLb2xeHsF+V4B4kgMCEigGI
af/V4xDlKzS8090sRfadlcsT6awpF3UWClOLFGNPzGWbKvktHJea90NNioVL9eV8
Xn1V4QmqtSRJ0Sm9pkT5NaAeyd04JoJAI0DgSIsk+wiagaaYKrKICTQ1B81MOnZz
3xVgE+fs3nBPIje/qpaEm6WUBdhzwqrX1dkfSmE1eP6HhcQHI2GefAGylpxJrPa+
3KjWcijB93o13FrzqOhXMGx+hVMm0iUTtB+9iwhg8VCStsqj9B9py3sfc91pbq/t
oExqSSghV85pl8Krp404DcFXFrwkbLhiuJZNm8W4813ACRBNkQcYuXBqlebuPJcj
H17Fn1NzF3SuHFuiPiTgS1GCzVqQQHbvjpD07xdklRiR3T6EJZqr31m0rmMZDwAf
d+m+8CBHLUBOzrb62DwLOn6P+1noQeo7cTOtyymtD2Knf95EaZWFCKPOcKsa8Qj5
T8cNJk6RcWISsT1wEgRDsL5Nu27Fmi2zx7YQ6HepSu8FFp7QBYsrF6DulP+42YG3
PfsvLVBKPGQ3Nz+HpNmtxVfSy0XRMzAP10uBuDm+24E2DYPxGoW/m+iBGg6cYiqA
CTLJ6j+to66GwMg0iXpbSuh0vU93q73QSkepFk9X94aIl9A3Q3/O80i8oJWutXpB
JUz05PvSWkyxVIZ8fEOE5EYAtYpreD9m9RYcVEnsM9cRSInPD6ZzKek3XmBpbHW2
PfZiOV/NZtAfjh+E5/G7KZyMbC6CDlOdwMdac1n6XPrW+jiWN7hDfx/g0KjcA72P
a1BwOFE4Pst/yjm6KrLY3CsCnKmhi6YUF6Tkua/GtPGNXmZ+oZdPjMAbDp34/ohy
0MrVhSeBYn15MBUjIDsDnCCar+Ma4Xmt/Y5QI1iExq5mCkowGjQgzdQmzgWaNnQQ
H/KjGpukz19t5lpPhdKfjfcCjonqwl5Yu/Zcg8ks36kqKgRpZovV5L5eYrlOtsti
3UIiRd0erxXE9X6zJKET/2uerBwI7l+pa+L3zvQHWp36h4atuLZvAfOtNiAYyNB0
4oCdEo2GF7/vW3F4JkCV0HbBoAejTntyBrtNaI2BssccjElxSFCWCey5X3YqrWKk
OKklHnWHxTbfcFSlRfA2jDxaLhKrA2bayt0gDq8BvduR3chn8vzg5DHkGQdUl6uN
CeGDj9HkRc+qKapEqF+0XEgqcMB13C/jcS4jjDpIHdUK8jTNvTbtmGPd3fhMMaML
d4OmNvmYQ+2PzJ2v3qftH2f5IYcN2thBFVfZ0BwrhDhA7S0P5oRthbUtA5d1IBYS
KGGxUonpYlKdfxLb4X4vU++JkhHt9HW/P/Apk52nGt548r7UnoQcl7Zwx4+SGhwp
t/kkBkgcou9tanyY8cioRdGVtrf/qOoKqN29b//vlnzl9RNt0h53mtZ/mxYdDZxi
UwPytC1j1KE9eiCu0cEsGGf4WjqzVzcW74Gv0xBLqqOg7kqPcsoPw3cZmb3aJNM0
H2kPaAcdxVVWz5IRysF283tCfYRKVcbAwGOHRm8Dcp8JDhm9KlNrV1XKfSzflZhD
NWs68gKJ8yxdCRVvRVbaqA9BEKztdq2ZtLUYWxgLQ6M8eoN3V9mHdXG72aPFRBAv
1eadU7HrfMskHHB9cbENRPYP7Ixk7/QplKU+eIzP6G+nXMDFlUHk90aJuxjDgErq
edwEc2T0tGc9oEtKT5y1kF9woIZ2XAwavC4vV3+CMXQjjQPmQpDCZsr6yqbMfSJn
SfH1R9EPhmrzIBeLIycxTqskcW1+8b+x3ueCrPo3EzVF9CBw6xV1M8X+EbO+iybo
pIo7fBiNxf7W6SLPHAoOrZkimkiWnXgMQAHtiP8U6Knl6bYsHSU9VLFwLbgXqQUm
wqGtwsThftqhE4qZ7kAS30vTXFoHhPRhssBAeTzLOFWXYyipGFYWZhufmJo6xuen
7IMsXkkU4dWkXKsO5Cmij9nFgwa7z/W8lgFDIbbim88Z2hsyK9oqDRY/zeb8IRB0
JQruQuNr9mWiLwutXpRZS2bZ5YOBHDIfKl7a1K87+MLL/Dx5x9v7S8C3ZFB93ff/
pa0r6rNfYf1SxcW8vkmIiBPoo9S9u2FNLywR4Mc7x7Cp1Ga5z69goAdtO8etXXg7
YK1/p9UQP5iJDN458Kpk4OdfU3hQ5Z92eZkKWUTOqErrtiTKyt9oDhofs+Zm2/yL
3T371acecCVY11CBB9ASXOpN8QXH7keHXuMHQXHE00BmbkgSKryy1X/QzTjTnsP4
281XlZkm/H8GMrSd500p+mMQBIMFLOln+ip814ZZgVrdQkJKHZxczjDS6S85byXc
a68yhvBJ7SMUhC5L31YVQeSOvzy+BgObFEchK106vMjGRwaXAGOBtqSgm6wvjfK2
WcgZ7tarJ7y3MbbEVAqIZBnhLNqoZxjX7KGjOqHuAWozA3NUrZCpl7ZunxjzCBDh
D3Ct4n/0znYpIYcdBrnzITFWaUuuCrBuVjYOOo0N+jTqid9IEpFo5DQCwJOE1nM2
8EA3y1RlLc7oMdv2aq3y2HcU7IABy4mxlSxVCu44PsyNVzmr/Qquga+9SNfwQcts
aXJq8MOVhxJU4yYSsX6arSIh2KYri9g98alZhELlUQ342YN5HmqpdipPWyTzep3c
/Jrrs5HzaM08VfHJuKCs367lQ/8HIZlve0ENmosmbZfqnROm+Dx7v5jkNV/D7rJC
Vcpcvv3DO70dRQ1HKO/vR+FSvmyeQ6okOjAzrEI+hzqOOf+CNiwuWcV743id1TzL
HUMAPT/gWwXrLM4utbGccd/AT5hloJ67ASMmNUIM7qtBm85RtKebVLojNM1JtX61
v8msQrmrDjyxx4Wulfl1QX4G0Un3U2y5qT30wdoMJi7Oi4FmiCVoQO/SrAxXcNl9
kEOKJ3fYQU2sGtAaZ657/6OU8mpTDD9b8jxtbL2+PrTot9LPfuFBMQCtj/uK3xvk
goAWgLqVWnD/chqirKOYIOFgDLXNwt7XAuXujKIBja7C9jCEzbnFd9xvQIRVTfjI
MSNTaGiB2+pBm7nAw8xI3vFKwxQLq249kPplfzdQMlsTSeH5pY6SWQ66/QpT1CWR
JwLnNOVhq02KcIQWvIzJ9sco121L00q54AwNu0QuM17MgLhb5QYg+cZqWaTA0M+l
5khh50TsOaH5gOvBHZagcCEYF7hjhAoB9ycDzutCeu/U9ZnC/LTy8rdqwvZZx6BA
lDjPqxes0Pq+teTX4wQgtK5kclSi0TFU1HYBo/Nl5hgw1HpatpuWeZYQAl2tJYl/
YgNb6w0EY0tfRbYHyrYfk7KFKxEqOW0OKbDbMK8YgxY4jAWGGnKbTIqUvFjebYmN
>>>>>>> 426889eb8ce467b9c9a9f74dd4af433c5046285c:deps/flexrio_deps/PkgNiUtilities.vhd
`protect end_protected