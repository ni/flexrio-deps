`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4064 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0gQgIG1mJzulW1XOK5NnZR8
C8XqDUtXW7uOWTnSVqbIbs6RIRkrbLkDIIzCVebsasDaW9BYDzIQzFvhL0e37lGj
hm6feTOkMDtJiCUUkWDYASe+vMOtN4OXj46rJUgvVEj0HA3hF3Q2awktwCLAcaQB
pdobFesoXX8mz4Cwwj09WXPh6KeNRJ+DROmIwGaMKwlrK2lwzEbyen1PaUPqciBr
Wc67z/lHHj4zq/tsnPiw7zNy1EONSNnrK5ZlLeUeJwGrQmeaBKY3t81yai4GwL6Q
sgQ4ATlblPpBQadFpaT3TXoaLfcoNj5btEgaM8k/ge1V2LtN0vSO+d4ZXVO6zhlT
6wJfVGej7MVuGHcUVWLBPH1iu+6Geog9FkyIuRxKA4B5XbOAfZkQoJTh9iOjoYYJ
nWUQKmFK08B5kI5PR1pH2iSII7s9ExI5GcyZtkem3xWr55wM7JlO3eyvc7oAru+6
uoZAUxyIm83D4cC6T2bdI1Y01OcE3Kv05raRuaMv5vVbo8TphLamiql8VQSTbyA2
pU4ihxvn5foA5KioBI7Drz31Z2pNLvV+8vHWcL+hEDdn5EfuK1IAjbT4gS99kF4g
BKtxy/BP/17b71FQF1/ZbEM8d9mKF9IwplKVuFY+62WHsiffwvpz8grUgtrAjLZl
c+lj+/W4b6cUaisDXnXwYzxxqyy88fitZsl9MIgYuN6ADBUI/JzDtkJ+zPTm8X5X
kHENt/YeZX//L/KJHJkKu1IdP106/S8pQByrVJdd5du9XgSxsi2g0HZZHAOTytE+
dZWS/oowxpEDXXj+2hpfb5zPdS6zOoXsvxo63DKVXjg7NMffhKmdsyuU3c0ZU3/H
B/hJ4y/2y2oVcmBPHRL6qoGX+mLrPr3Law68fywzir2NXPnGV3K9VW5OkII0yL80
HX2CJI9/V47vjv01xCkjKrohcskqpyt+V1Z0zbk/9t0HKW20dk414ukFISBKAGOp
uEEZ2oLZ02j5ZazipEBjkMiAWvHMF5zZ3VTFo6lKN6Uhqs7SKPfzXTls2nibnPFV
059TaTrPu8BGT9zSWiwmOUIjIZRu3Ct+MenY5Q1HfVSlJNFH9wySZ+AlGOxa6jMx
K84lK325+mGPQ8JtcrH7tWW4rFRAa9sh3A9lZuwVgvsj84e30wplATt3PmTf3enq
a1zwQ6QJxSlK2+40Cj1mm9/89lwMM0JzYXPPfcvUL92zH2OzItXVGlAanyEmlzFs
CddSSN+AN4NouK6xRpydcI4T8kJW4J5ZiOiWP1A71vNMMwRfDedK2BeAcSwphDEa
tt6VwiN8LPXj2dL+k5NFrjLSfXKRKkOeqQg7bIEG/S+v3EGaSm9ROkF2KDewZwTy
mrrdo9KNYAwnrbLj76CQ/FmZ0jA8EWHk68atItzjQ99yI1txTA3FjOIavS5wk4De
06OT8DSURMfqV0bpelL/QrhKU5VatBOD9D95c9AhnyLvycM4QZ/g4lvHvL3majhv
hOtpTdrxe0BdC+MSJ91PkCHA5TdBLaqxohUXQd4YA8t1udILE/tox5sHGZOYQI4V
D/jkTqrNP2dOrwcbk98MtafHnNFV7c46im2s5Goe5/U5BHZFveshaMAmA3xZ3amA
aQh+Gy/6wvG7X267qw0CyCUdxZU2IIFnelAlxoh1qHzDEk9yCnVSq6wuphYxC8IQ
pWV6Y4yVGr6faCfKASmgrqAJx4dwCaFKN7x++qJkB3dF2nWRVMwSgccIXNSNbGXY
sMl8MVivj/dPoE3xFO/FUQkEPKNe1+dpidb2CfeUDx3wQaBjEwbJz63fLBaqXL9k
VdGZ656X1siifEgYQzCHhmd/1WwjiBpgS9v28oGDFJo6caLJ3pNfN89lK7jdsom7
ZH7wyFId+AF/ts4Le5e6D7ajCiKIDYsgezKd6rLm6754RDxq0peEvR5YI7MFdxdT
Q3ts0IMTBdqTEBsmHaCY0sQypj/sj9/k/m95M4A02pFyqV7YOKPnXrFNcBESe+Ub
qD0dQsf0hVRYQ4zYy668tR0LoxOhNjeQjiAInlT0QRkB2bwQBtoHxapvQn6urzKI
4wpZ3GufzFYquWium6Ya3PF98LNXvK2WgsRAnyZHB1nJzZIdTX1T7EP7sstnwsZu
uarbI8+vpCb77NqX3CRsNGKXcXIjdhaDpAfhVOT+gsr3+Zf/onzIwHgN8LaHLVKH
oVu/oeD3eAQO+IYgc0EPYPIKEnCDn758IGTikEPln+7Driu+8kYxEsLeYdNA/Opq
gw1t9euC6ZHrs3ZfhdaJWO2QTh7UjCEeWylGRQwGplENXWGUBFPxkySVsO1S1JzQ
XV4Zy5T1Ww8rY2T0Du6M4lk9KxGPkfPcvOyXBhtqqZGWmo1Xd22cRTZIllAE8wub
abn0yVmaXQPhnznOdULlaakmGcwrQRTl0e3Rm4Z7UUd6nvWpz8qnkyg9gywsVao0
qeniwqniFWqMWMJEqNAQrx3ocJd1X19QCtJdJ2VrDWAHUxIZdSzwJkvejfwK5FBD
kZgce+HWuhm6FhApvzfdLTdYzNyEuzvQeQJdjE+ExAouY2G15iblYl+rE7yqYhn9
X97fUwHrqbZShZS8kps7rGceQ4UIwnZK28w0nT4Sx6y+4/EQSbWMXxLCsWWmxXEJ
sQhpRvHla+Cie9AyPQAYduPHm0Yja+TjOZ/6vSd/t2rwdazi6+bAA0NialMufIIv
9Mfc8oTad0M7DkCwXXIn7ouJ+lCB6qry5UFpo7VfXtsodUWfJI4Rw64oh+TM5VBH
mNeV0hJl7uUrCLepD08w0YCj82MY6yYUPof0N/rrXs7TZYW+Aa0njIQM5yMviakr
6gYCikLiQxIJ+U3Yc/ZQUzvsB46UGmso9GCSpYcVjc4lYs9kwrcwsS7jd3s0objA
lTBiE6sFqvZvYbr8LY+npxPw6gjJuleqmNWIumYzLK9yCdVgQpHCJn48vFjLEuVY
zZVp5hFvcb+LVSxh62HMi2s8rHDjuuGriAzfyExhNGaxHVFAc9Kbn2+eMpD29mQ9
YdKIvz83yqDVOXGOLQ/RHxu4MrjD0iw32buhOI/OVc9YiVz6SyZ8PMMILUfQuAJW
lViGZ60e4yaHjlJo4CZHYNdJTT0aAsYV8p9Aigan0636bWszQys7c2XkrPHbDDfA
r84DgYQCJdF/b/6pCB616vPCl+MR+y54ystIeQDEkMxNqZ4d7367QBONV/h99LHC
sw+9TJpn5s7B7TAf6hF+d+7PUhouQB5zn0SNM+rh+FOn9PBXuUX0HEv8kqCzurK5
UV+oq+Cg6uIfw52ghRHv+ORUJ8LcLCeYncYcSGIWm71sEYToGfLUggDX+vZxpEei
EHnkHWk62/ihDws98qAT1VtKM2N1UEh6VsuddhwuQGT57fGAwJaMWENK/ROLrLJu
J+SrGoPxxupHHZTdyx1fqNj39qYuQY+mrtCjRtEgMAxGGq/x4g2yjRcYpqzrxSP5
mHXnWbK5ofT2B1PAd3WgUB0eYgm1fKr9RshRfBJ6+XYSh3RU3mLTcbJjk3Mw+0bs
G7lqCFIaf29RP33sfYfOL1gQ9BO6LpkS69HHWHebGtCgLKsoYBZS0D7JTjs1dB19
DFd+ZAfxPWnjLqnfPLE4jx1IbB6cP2adhkQRPNXGrP1arcW7wZu3CPmfAxxQXiwM
NF0Dgtt76wuvlLC6TOF5B6+Z8WW7GQf5x82CQWjYao3dOA8v75go4dP3od3DEpiD
fdLj3FBBSl2X7PEJDJSGkQ5mcwdezoX5TsW0TGHw/wrygodSYw8Xl/YPuhMiMWIR
igr/zBH1hApwnQIsNtPJ05glyq2ACazfgKi2PbE8dlVDCjStIcIXi9hK67oQ+5JQ
ITIuaDvFv+70YrhstRZr2p0cxBqzGVeHdWyVbPV1hb4zhxLjGep91fp2201fASqt
nfDJ1TGPnh1aHLcO71B0VuA2jUG7Ioqo3q+rcyBFnOsQ/t8yZ5X4NBw0NCFctDc4
7/ZGRQrbNiizroKep0ItkCPGVrKwNN09Ore8eXCSDskBQF1Yc6wlUdzZNGQnHOsb
FSx5DJT63H+WX5utK5jKlFQpS0HVd04oV/n+l/eFYagJWvTP3BmavZOn8yesEFZW
06LCCcEK9VqbgcPFUwg/WTVgFQvArn0bwb5Ww8vYPjC1dssCnu6TF3Fldaqhv5so
edmzb8z4dQy7N066+Yv//dHldvwclBKKHeEEk4noj89fyr2kjNWgn93pHZOn1ian
OD7P5s88mOc1mtj+HrZOrSfzeXuAVTX0J4gF+TyrZ59aBiOVMoKW6iDRU42Noodo
7UDbizzzT2WwINwo3OAJCnTqOC6UcRRWeWyirT3ddaU/VVI51YN3x7A5RdZ8zCho
NbKvxlVCvzIV6ktPojXvvUanG5E2MAtkDdqMmhNYOanAg9sxD6z1GpQSQj5sgDcB
nh+NgpuJj4q0qG9n1iurTKPwpQNNXKB8/bLoGwWQlgNyfd7gtmEdS3J9XbLGnxVx
jZcx6SgjA24xzQSW5cXm9eozcecmZlVMbWLbywrJlFTmVy2r64V0QJQqCRpZxYa5
L4TB7hrhk+X9hGES852+XularAKFl4aAlZV85lhekVA5ciD6OTFB+Rv4Y8fIpkHo
tThA2lAMbmxYWj5/BYW+YSCvZx6brQVfL9gmXnxvftks0yPvv8R3SfEXit2RTzpg
c9/2wZGK3+EgoQDEZ4bn0JxJZGk0lzz9ZQ4S810eCKhwH0Se5KLLsL1VzWnIE0+L
Kkk1WOgROlvhI1yfk7wqOTU+Kttqs38h+mr7R7qJ+quvYr4AzRGASuTEVEePWShC
MS+akfFlzqJhtFX+77W+mxNj0PcOVKAyAmQ+JFHRDXy9CqZ3Th/m8nxxPSB0yIXJ
44Pz3QKzz4ViQzFP8TbyihN56YCQ+UAsDrIB6PKKt1/OPSt50Tbt/SKS42QnE1ne
TY/bU5vNZtMj4sSRs95iPGSzy0Hi5HhYo2RTXoNfyYQnot5NKCwVnxKRHALD5yU1
n6POugFMBgH/aca6WLD91e4PseOn0Za1jPU3nHBhnBnLpzx5kHP42A54XoiJ1hZk
HCgbf/YVHlG78DB4W/g1UloqeMBHcG6nxTpwcPkUiFdlLum2fd/b18JvQs/t97M7
JjaIVAH2zmdK66PcaI5GQttjTjwZ9wQSRWz7eSLKBTPMJA5iRu42yRuJ1FziUkrt
kO9lt3aV/6lHxHeowUPTmcpMFh9h0Kn9jeJOPV8fNAZlIOLQ/Sp9c8lEqpCnGRDr
e0dRjzVZ9z7yrtu66o9BsZvq8VYXl0pj2A5xtghrSag=
`protect end_protected