`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 61520 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
ZIICkMu+S2rq/yOQyqhpuuK69G8muJtMqZIdfbojJ8gGVC8zbDzUVXWR8VF0YYN3
muh7Hx1bxRaJjfX1ukLzqAytG6B4hBi4qZhgdSVnBVcpTpxr/pSmD9k4W+vpvpVg
+H6Qco5JNo6u2PJssDAEtYydxG+H2d4fLeJFc1/1/qP1hydUj81VJ2WuA/N3FITr
WT4viYW1CJLI7pzGTP7Ylv9QEXQzFDro0fC7AhgAfWFskABblE0A7RZczOBpBNgT
er3uv/+QFWG+q04Maus0HbaTeZK9JsddWJkFRDft8wmJclOLsU5j5nz78Ze0jgC/
yuhHRvLNAcSY7sTmbm3JjFB8cmQi0NmJHB/MSxGnuhtLL4Z0Mt4/4OTSgSOvD5BQ
HcdSpoWPdFGiV7HoIyRUMWcl22xctOvEfCFZ/ewGCb7zfQ6l1UTzj9RT8I0RZ1tF
7Sk70MjZfZdcTZtp09NMEn18Y3Zxx8CUN/yWhpkZBZtXT9f1TjwHwdlW3qkbov0D
A6smaluHRkk/hJ6+ywBH3ijnRGN5rsuX6a1BNQS7Kb/keT8ak26M+YUHWeRXF/ex
ZxUP2aRzdo6QewGVTF38JzHimt1YvGB4Wk4v+B+x8z0L29IUuBtBWbr3hG2JQE78
RFWMocnLRBvux4Lvm5OP0CFahpBlEfR6vdZ3zIs8o7lIFfYLMRsxQxwFOMncHbbD
abI76CgpjuliUFImWYV4Qp5j1S3+7SO87bjmg+XJqYKJA7UNh15TARNnkz8mImhp
G/E9TdwDYLXEy8eq+u69Qayo72MIR5y1570TfqAV27CRhRglT0hR+xSmCcvvndBS
cxfA8N8/wndMtRGqzXWoyAEEeFU3FfYO7RRlXcEm7rU/x7PkSZmBaZZYb0RlV2s8
utw3JVtj6bR7qnhqaziZ1PprnxhhPxvzkqMwPgnZz/T+EvOSSFTM64BbhSvcmjCB
3a6OhIyhhML/N1tW2qIEo97V9xuYshksXAKT5RDNkri5NcS6Lji95yVSnV5Yu922
gVFAZEMfVYqjLM25KU9RulCjfLg1pMW5c6z2pbgMy8aLgGSM7gDtSw+vKohEpOys
Hm8oeYCROKn+57Z0reRrc1cZNYFYqeaROVoXp5Cz7wbmS4qzRkWZ7wHsSJwnrblw
P1Xff29tRAWdI0tyZRQ1fqpv8tsuJqW01y4OL3+nDVydUayMvP/1ZU02KMsrOEyZ
70gy4F07WNNJdvDLMepxSzDNG9jt+2DagmwvJz2vEoDOrLzaGhwXd/w5cA3KaDdT
lf+Fshd3BH3iVxSEmYw3a1uc356IBdCFg8szgBRkXpjNYwDRvGwTYBAdBxp9qnpZ
0iAL/tc8XFtR7zXmObS5CFz/WHRM0fPEPNJyYH6tp0AbtUSy0wvc9oC1Knwo58K9
WLaRkyMRaX8Lu5ehhxUaGjbFrgSWLd3xbvzPITdLYX6nddrc130/RmMfGYBbQo6c
9YiXEdGqScQleYqzjyIzn621mVyySPBqRIXvWSWV/v2s0I19ou0qCyd4nlB8vzkM
tD8mQrIOaSkfkdZii37a2oYvUzHzuyYElrQ92zESJ5tXbdwk+32GJRbfW5TRJy50
a2jK6kP4JEamXAbN2X/c6e9ANxV+rTZE5N/6FGY0+DUg4/5d4ZbcEuKjCsdiGxjW
Qr7wsxolPiZwHC1ulpVt7YhOsOgMdp9wkJPGDOyQloz5qQzGbTEWRX6o3beO2+T9
AoMt/CK0DPd5gwYnFI6sIs6y/UFDR7zBSK3EAL9IA6RCgmIUson0UecLCRI+LQ6z
6LuGbH47PijhQe1wQyMGilPxUpgFXSs64Gu0qUtBPw5OtzLrywOCKEOtN8J+aOeV
rRxcFj4nnZAI3LwzBLX/Ol16kHKi18XoM/SMOhe3X6fFF9wCWASP20BZ1ouctdLZ
Kqjn5MRTlSnlRi91JteDmNsfZTAV/7ThwZfxkp502a15fm5n51ALrLvQ6A3QonYn
kiKRwGEGeeDWLVFphTq3NlSSY3W7ghtta1S/zn+wg3vX0W1dvjJPMYEglbUrITMQ
l24EcNSX0TkPL//D2+c/dFlOuUUsbIhIURcj2KUwW3XxiQ2/KE1eqPwbHheUztuj
gYuYpHrxsaAzQ3swG9IprKVa9ZaWQOm8NKMLuIgyYMdfbyjVrJOyHwgmgj2sidCh
m+PkVZ1Omqn7Z3xhwF16nXQaww3g9UM7/v5tRUhCZx6KRYQHLW+fFGSFLxjfHcbN
ZKLe5NOUGE03j5LIJytF0Jgs14Riod/rEfa96YTqe+GrhYVoc7jEWpVr0vhRV8+E
VeWtFegEKBzlYMy2z0cnW6j9aM400nBMLXBP1gmdwHNq8UvVFgsD1wbtynwCvQ3F
mlIgt3riolq+Ar65KpU/sb/mffhRPh4f20qb3UamiJuVfm3mC/ILjaMKfESm7YS0
YN9Xe1/VBVswPpQq2bGGDtGubS3BaKMEieMwFs4I4REo9QmdK4poQkXRV7Sdo2Va
3p49duRVvvTNFmLEjlJqqzQwAjv4sI3RLHRLlL/PPybuQ9TZzrVwUq7tmdxeKsS+
+ZTNJ9WYQPS86R2wOsKePkXTBMo2Mf4SV67GGjmQDJlXiLrmbJQu8IjH34oEnhBV
urqGoLP9nNIsy7dBmL7vPyqUMRcw4BWsJb0amGGgMlsfWIBxA2VS0aCi0oD0QvKT
cCqbWWkFdyK3tvjq0kH684sE9MOuXqdhU7IWGw3NXLBwnxmJbkmDCs6FcRJC11Kn
ab76189aleZBxOIc2xMkrhXtOKT4VqthL8wYdJ6EAFuOnflQQohrPw9XRCniI6cz
r4MeWlxSmGvhmAQAgtITDVTgtycJG/S8LpRpMp1f+LKMGtycDyZeznA+0Gi4x9nR
7Aq9SLrKMw4vduMiuYzUW9CcP3mLyjkdglR4rDdWhfhaF6V9x5UuYKrpa0YPKrJ8
EDCAIEOsTL29n1odJvZ0xpEer+q2fmpuDVDl/AVFVdXozgUQgH5eeAMOn/Hw4gRd
iiLt0nW5saQDTFs0IDIuPe5LNarb/1hRx5kT48hZDqQNe72NH1mw+gvKC2/RTWkN
56ph4YxFHSal2oVWSk35N0Nx+bgayXbeYJVohz/nhEtiGfXSNvNmSatxKxWm+O2o
APPlOKdte33/U4wGG05Z9hLb0jujWlWfRcg5jPQwyyYENYBXV2gT+PuJN6vt4BSf
qEhy73V5REKr+P2tOEy5ac22BD599uXHyvkxVBBWINTKUykQwINnq7qy7wnAV03B
pUKd4qX/T+NbeRzwTFpX67nFVmRmwnJ8i8GzNKM4r+yO5ujphxPcRFSHv/XAiAP5
4REvLcDk1zUV+yXZYEHuC4yuhl7JE3ZgXHEANRXfRpwyjqvk6OG623xTMh4PcNHy
KZfH9W+bk61vdKBwFWrszMwsrTRtTZm/iU+RwjWhV8ghFpC6rPxdrUY8JBaWCXF8
JzjnU0gJb+DEsPIapyj9M8wv8XLpgZXrxvUqJCAniqzOzxEG0jm6SaxkBb31WLVV
Iab2bRc0qi4co+dmx495z/7IUXRvy2VTEn3Ewb97SLSnTqiul+YKKPc/Q956Jc3x
qrymIz6XCTIEnqYl+ILSfFWI2bR1aP7IPO3FUvJvV7JgSoKuEue6jHhAfPB+EfQl
vauywSv6z6tLbOXiyalRawGg+ZcV3w8JrflnGS5khXHvxRplv63zy+q1KxavN9qU
WYIUdzOtN21PyQAoqRGvr7El62Pb5qoO7FS05jqajgrZb33JnFRohu/rO8sjkq3m
eNRYC6oGkqFaWs2l3bwNcSU1ek57qOXpV425PhyA0xB4a38hVxscbjYBRSIzCLdi
ib6hE7U1wxrg1MS8MUeRPow/1Oj92jtCQQBj/a++sM9Wsk9veTLV5s/sqzZDMBKH
sO4aYsvODGfLnbwMjdbA7H0rgFes2Om0FSHDBYQNu1XZ9TZ3EOUyp0rIAcUZPKd6
3nIA4g4gmNWGTKh1nI8jg8CPdeDaHrGFirH+HtJy+8ukyLZHz6kIJPi1x33X/pcS
Hmj7dK/ZEK5xQj6K4QO0793RDsRqyvaOmpm9z0qRKb7xdssYYoJVCW+ldPMSdK0N
G6Ydl0H0ECd3Mb1y9IsCRqrU1O/VsEhLX5V46L0swIRXlbNwcGfM+YCFAOM57pW0
C6MqloZOZwFfOyAC0kISfzH9R5SFm0Fj83xqSj5MnbvwPzo1ZwmEnepTnAq2BV7+
SUetDFYKas1WrUgu63PlY7VUrrCFR/u5XmH2//PTSYO89OkcURvatGT3P0RrnWex
hBUiTVVsWPn2m+KFqgiywqVMaOSGxdyDBXPSktcl6FmNlYU4TJlW9K/BJz1Rshwa
vFGeXnuHIb/0LFRKYwwDXsUhRMFndcRUOyGIKQh+kPpOA6g+XpHHGe4NMBELQU9V
vwJULaJwVfp+MWWuxzV+j6QLbd3Re3KHdU480Koq6hyaBeWX83Nn6TBkoqZQlR7C
wsADjKZJDnWHF2J/bzEE/gTfwjPr2w4DYW161LLjJbr3AG6z1OVUs72xHDKv+mYx
UP0JiB/Cm8w3agmHK7kFPINqDMPiR70xHQ8f93cLJ/AhIyHzmKll5FjBECnZWNqo
UHI9tN+UMQRkM3DPXVN73wfNNrBP3r2/kFdSJ1S6fbo7I8XDqiBjUiFJJZ7X1z1S
2J4wPcF6p418rVU8rfhbSVfG/9HKWa5bszDxhfYVfolyCB5qmScUCaoiLGLs/E+e
td5acBc005HP+3ok9voI/aaCdO2bM05I8oo+0T8RjO6m0XPolIlZBSsZgVbJeRt8
CexQuk1ZA6fIIgvKuEWFM7Zyx2MrEY3vP4m3Kf++QMlwuJYiq+vuajFJ3Ku6C3J+
4wPCgkjYKAbp5Bd2ZG2MLT4yCrOXlGwDOMZOumQk7Z3Zec8M2eksKDDxgkogLmqM
/4hXuSbeAKdt9faxbXvOxMZhJyCqAs+WHFDSWD7H5lzKNYb13TNDiZqsRwyVEhND
ArlBLlERX3fzKQe2W0z3uhkiRZvDLLnO+L2Tgr6j52ydjR7Zrc6U0fntQpdnOY9j
OghtVFHhK4J7tYjbGznS79bd68nQ3/eOijFo2/u0QUOrB9+IpYMPIRy8dMhpGajD
zkFp0oQ5+yT2Xbhenl1wUuPNlBKtSf8CDSFWoICgnx826YFl9jBx3wKfCuor+VVE
sU9DSlEcImuWsbm9ygzSwOUFmj1g5rCqGawWQaC19R/AzpVxJMfHoy/cW4/T83ZO
hBm+ks31PY81w1LO0rAP6bigQy9vdmXHigjfPyee1oIUDK5c5jMFA3JegkeG8TEM
gr0h27rLMlXYG6hGJce8tqsHreRyRqS1VDXM+SmzTJ1/sRy6l8d77xFyg5lyde5d
ZzSUsvVFIhlzRXERJSFJ3RjKqBdBl8hCb/CO7OCxnHjbUZvxvpEWfPW2RzeBlQeM
jAickN/qO9zGDQPisUlb0HjYuNgfJptRwiigCGJvOGKd/YClIHEXABp9PAigttJy
CNPv9y2k9QpZLboNS/P/5bocuAHg/t9wIGWe0NJeEYfOcFPC/JgVddFs7x5y/cY4
9pvPeEO0L7iS6fQfVz9hpr/VM/p2Q811fRpqaXh8CnfU3VtIGWvXwmz8wgRDh9j7
aksjqyPq6xogHzwWBghwul4wrbab14jySOx6j0eQOHtK4pgJrlNPNT6GPWFq2rXp
QexOrylw5WxdOkn8h52eVQyI0b9yZa1RtUxGReDSwOf/LdqksmU6aeWznv9xtpAz
Efv0XHdXrh7PD337Cd/1Xl0GOCAZk5aNlAD1ml+t/exhitgNSO13D8CBV2PABb1h
18f8CUCZMJLaX+1/HHog7ZDiqhgPMuj1Bm1ApwNtKxfLjExVX57OYROLxZZyy3a1
+mK+h07GwkkeHIaBZPSc4EipSidvd+Uf4eoiFv0bMVe1oMi3b7+rwqda2Puc0/Hv
G9loiFY058HHswackerSgXqF1hqpwiPmFVTz3O9qBY/dkVpWoMsk/SuqexwLol7I
6GeAPGAhzI+JaQMzsQtWooAPEqOK0iVhA8Up1V5ngCKPr89JVcSlz6l/mWlIR+On
QL9FcYBE4rjNKf8TQU2mn/exKsdHEBzFECdM/x2tPfvBawYaUvD3eLf1KS+kWMcG
gBrE+6efa/x0pbcqF3E7kePmZG4rG4JNxvvCVReiOJRCAK7d67mY67kJxGVrGca7
hQq26UMrusM2oKGTRHggTChCUVW6Gfzpv95mWFhlCcRRW9AO4YJ6jAdtd9Oo1Y/+
PNw8l1WhMZnIjde94unP6bB0y0RmbbejxABS1PDfLqFHA5yUf6vgl9LwgA8xepNu
fDCvQASzfelos8HQf3YEKG6lsKmryinx0C3ViIAtSl5XkwRAJEQvES5B1JooKYN3
/eaxe7IDIbtYfvgChDk454Z2manoZi3YGq4FIpyLb98PHt1Ti4rLJBd0ohLCKkNv
fQ45FOCyvegaMgTRWHnRVuOWIxCVwVVM7+rlHzBXzxAMQZ2KSvcp8Gu2pJ0E6AoV
/+8luk0HeFtKMAVhsAHPieRSyhhSHZYhGJqlGaHDcdB/QmRLQ/CEEPXW4ccpX/i5
VdjDQLuJTk7ynhOTo3EJ8qREgg5gMgSEse+0DDTmPFMb0kZza5VhkIk05EZ9u6FT
H8LllzdSqXRNh7uT+RlxjCwo989Ozbw9wkxEpaWWdL5m3X9N16KsFIV4CBG8Vchj
IygX4rcNrsggkXN5toiTcOtTM4W22PzKWnGSdQle4vURWbmRVd4rc6bqPcscX83Q
d+moaxldJj1vgkuIXO26g40ASJZhiWKW4TfK4nxys269YhnRH/2orlNIm2xGN4lr
/a0g2FqURMwZ6M9EzUh3U8O1KQPlIPuIuKvykve1G/xBRN5TPtvxyvKq0nBoQHSM
ChCGwGx+NO9rlfHJOouNCgmCQzeUwxgvrAx+MGCQgimrfmnAO2th1aMutScJmK2A
6Q6wCtPA5xELjYjmdeEvO/+8ljrAr2ZV1rxCmzxFJhUb7KVQWAANhuErolNllob0
sjtRRO+ZR0jLXs57jo31+EgPRXmnsCnzlvxHzqMjRhBI6zcI4QaCGGgKUR6polVp
zjDwUe8bjhoU+LvrAcgi/qM4bVQRsVSxOyxBDFqQj7MsTbSkluURwr3GSQYhjlWo
vkG5rulUEsaOKa85pHcyN7wu8yROkOdzb8SAI3JKPo8xCaQLpbhbukvOsdTDfQbk
cZkzXbdUDIhjZkw8bpycJdj6vaobajno8flzFwhFCqnM+U6RIINVc0OuQgDop9zE
swcENksiGvpWDwNcilHUaLSPi3ObIJLq3GBh8KrZXT20JUS9Oftl1zPt++0RwPf+
vRRd6BAC1IGDVu9AS088FBsT8NZ6TjHpitRSwqP0CDhl0latWPzj7rhy9vymdiDv
sWLoaPOVtkj35f2m/gB3+Cx8hebSCpr4l2DKTW4ojUfHcdNjqsnQ66TG7QhfMHsD
7vngi4n4YPNI5rFT3LClt/Api2RcrZG47Gg4fB1PPRUnWJQrVE3Lds5cdiSRXsst
Jk+DUU144SrH+gln9WjsG6hYkpHgfJ29Pr2Txb0oyzW56Oeh/v7fu7Ewr+lntgsd
FwDdu1NILQjsc33wK3Wpaez+JDOCaSBPLt2jbRM4lw1NNff6sJTCRRWq7ybLsrZi
/y7D0RJG89rLymZBqm26OQFMZ6Bta1YpvMmtHaJKqq7AceTwllY+2IhQeQDIiNvX
tM+wqrORV6PNsS/nccBxZs/qC+phNjJTjteMFA60sqGayR3rTYKOE/p+vxSBTn5k
oaBeDhF6BQ9gCqVcs2whOxOiD+WYHAS72bq6KQd/Weoc+YMW6ALoOli+kvZDhs8w
wBVRhnnR7ZUMSLPy/CKh1/zbP4/5Ymg+RHBfV7gIY9g09CVDs2OJsswIkVs4La1U
h67n4Jsv9eDyUxMwVC0LY7y8Ltf049T7aUECsUZnWzEO7Haoys40FTf0K5IyQNcV
FmzweO0+gHRLhqsbf1BRxaYOMc1X+0gPpDY2ddxZ1pYF/3PjT99egkzVMo6eaOQQ
eEl4UK/I5u7Zbfw+uGlULYR7FmObYIzH9Ebui4kV7yXxoeWmIKHDlIK9tououj5m
OFn6zbeRCysFX486y2gQ+YCG5pvKXeH+fZxwTikdk6Cblul/H1ZRAPMGBkdPdH2W
anXVl2Pg3TcXgqrc0sOpDyp2AzPhkA7osTE5EJt4dkKnyUBt1k9rpikRMNqKH+Hf
P1Ys/oJcGJW1ZhMQkGsoAzNHsshb/7YJTLnx2bzjRPUxfsYGcvcdEtTvXm5G03n5
8gD6TTtD2nWKO4uPPkXyu29ak0l53hf77lRau7+TPJyBvbX4ngQRjLtBN8MwHB19
tyAg43A5S5RdnGoeCft2X4w0EA8G/EjfBCxP3wA3frh8IgKwOjwZuUAXPgVLon+A
pViTzUszlNLhKzQ72gsloBScrqRrO/o4Z6i9qB38fEbkDz3/3LOKTpynMWSp9cC+
jW9JnBQSUTIvIUr3ncvYvcdT0N6Vtn81SnLcc4O6iN4XgZK9Y4zVBKD2u+JoNom6
13zZtt1o9Xq9qrN+7kd1PH0FSmxAvcOpHNkq0aCf85uQF3a6ZxSBX2RrJTy/MYHe
QeRMGN/jOV8xpi5JsSS9A8s9fRvkYKBl/JX9PW1jH2NtSsXsC6/MCi0iPgs/6upl
aTLlmmzBRikbkr643gYQ1N7/GjRWzSgaio5aOpxx8Xxe/hvc3KkPVdR7QK4HNTt9
rmqthGoQtD4F/n8FYEgDcl+80NV/q87wuZm5topElHjncbovzCcxtLUyRXqCfBCq
AfH4+Q/vTIKzZVTfS1gzMtUkia6ZL95D0nZ06au4kO7pHJu6gCkCkOvhaktwD91H
ojeJeyKbh8ptwGmbDy6tZXNjaco2OhIem0mfrnaNG6pfP+sxUtPAg/AToLaLjYu0
L0p6ooy3i7oc4dP6xSIUaBXYcMav3m0iZ4jcYgK9ZoCkaSY3vx+hGg0ZEetDSfS1
qczbDdgUpA31aPnl3kmd0qgVbz39rqmM4LXy9SQHxamqjY3CJGU1kSnR3RzIqlM0
9FuSgQ7Pc5wv/YF4T0OPbdhEds3ykOA8DkR6mCo+wGA623PFftDHxr18vBARjCmY
9+vsprIfSACwKc1vkJ859UrGg+OuPRS+o69U4SENhu8utlXbdplxneTSYJt60xLf
9rwrSYu2GWw9PwBs8Zd9SyO1wvR/ovINOZ5uSvy34SWxCAbANBr0gidt6mqdoZgP
vD6l2OipxDtMplDxPFOY/6PoSAR38Vr3pjaAgH+x4DDmCW0fvAJqsgiMy4WwemZ3
CDhCt56PGHjAmLxKvLB+IdyNJW3bPSFYOXRA1XLYQ5U+/Vag5Mdppx9m1WUKbakm
EUHoMHKfF2Y+0Ja6zbwFZb+h0qk4ZfqScANMTVygxy+nEs4RF87YCB59dejXx6Gj
d911+9WGDYkYoHWpSjDwuAKu0PN6vtXRCvWQIJIwymoLRw9cEa/hjatzzgtK9s4n
EigWswLCkvwWSUt/SMX4RrTnELnPuCij5leIDs/5wkW3xZOyVGfwvZGP42DhVphp
U19y7YNprRfqm4igavA7vZOWLC4DyXv8MdkDFcxTm2GdJDkDmv2ArsEdEKLACDkf
LucHeXyMNpcssQuwo2SUjwBz3/oDK/2SlAOYiQlmrL1uiBo3bKPPYGBsJO2NOzOl
jypHNhlK1rIeLEqUtitmRSyDs3tyz4rpdTpiAC6Vj0ALm/y8fHQAM+z5b3qJ0gPD
KYAg90tedZD01Eh9nAPXIXHqWJrV63LVtfmliNZuS7G9NZDRqChmFx1aS4BbA/Ah
KdZH133BetQrAUTH3IdN/JiRcD9Ur9wM3ZOk482GjYva69Y9NBTpH7Z8QpZbxLw3
V4Zh4dy49BlINeYsNOdLU9A9RK8ermja1zNEHg+5BLTxF80ujZi3+cq1q+5rYOpa
V44U1MnKVCCKOd/nU2foki01MP7E1VNom6Pi7ZhIgeErQKhaHnCIYUrS/37abxp9
/0VT4C62DrIIFKg9bIP1NM55s0y4kv4E5z5wfCaJ2VFBVsenfGTk4nv563admzbO
9PyT9OshzGPOWncvRZJilL4A/qG8g/+nYLTm6LvJvTgC2z5H3K16MpgaOUx3fSK1
uXgmMfLwtn/SHWrPtGj4uHmg/XWsWKi0sgqTeCImxX7MdGvOmTz80mKooizx8HzI
n5nY2c82xnFQ0DiBtG0PIvYholW2A3ip9bc4Q7/6PqU9XcU7k3q+FUJ8NXAxXOhC
FG772QD2BYCAVonRgqIFn9918gVjX5cuimAlyYwAw46sSDcR94S2BOFAv6OT5Veu
lV1XXtSHjOHCgIuZRfjNs0q77tpbtdboScA0eD1TOZzhhAiMH+nNSBK3pJrTqRp1
dXDOsTOAfFg9AlKjGLMb7it0cKsUiSy8ovk0+qdhe4dLJw9Ko5sbPoOMlARQwaZR
rt1IVxVK4ap5EpnVaU9mdeTODNXUxNdPpE/DVJZqnxgYSRUJUCVnb/lKVLZk3OIj
NW37Norshki5VD9GEI2gY/NJIVcr3oFmrvQnpPzc4j8BlVUytZsR+prbivY7JHrq
bcr3ZHlggQDvV61fV6Y9SYsq+jqb8/JUgAge05RCiwyqaX2DwBI8GsqelGS3wEnW
8oje+wmDUE+FClxlHRhcuFKIhUQ0UsjpYuhJaP30DahSDNZbCZBqSI8IdNbtNc9W
Kw2O4IoGdL3sPBHEvUBxl7nH1n88N0lZWsLmhuhM+7AvYfWjFeswnrxnS4UC8Jw1
tLHt+7es+5ziaaENE1ZQIxcH5RwaXrm+oc6ykQ78Xn46g++7/ZNY6Iq5BaR4MQDY
yVpJsbTm8lOT+/avhE88CmLS6QF58SMh4WmmV/tBClolsGjyPbzlgwWjsFuW6clT
msirv3JTyBZ+cz1Q9jhWw/89qo12cnyMUdioiOl1M+u4KMMv/xFMq5dP6wwVj0hD
9MuuqZ6KrdcF9TkSl5nGCvK7/28d8qNRU8LZtKZOiPqRN58Nf422H2cxnRrBm884
R+HnX1UoPADgJqxBLCDv9J0SAYzuqkjWljw+ym3cto4+e6k4aXjVxaqupd4w1yoE
FcuLw1idtglrOCVZ1dVo6wpwY7vGQCyLPo59hyASd8TChpd8W9WmeUJtPzxt21iA
JkgRrsl0nqB9ez8AXd3gZKRPAjKjbYYZiURKUvr8JOPeHMqptbXZY6CSkkER0E08
mJhFEiP7HrQguhlLglchBVNsl2LqtbZxWfzRhDE0vZ8CPeJ2rpiVrGjzPaJ//6JW
iIEUdJxM+0qYelMskouWTjrMhKuhmYzT7YsGJ1ctxIQX8pJf+Ha0HiGJ7i9TzaSx
FDE7+mwprY3yT9jdWTdMPiQfrbl9KhoK5GqTfCyDPmAMpknUJzWie+btXUq9HpGF
HxD1PzVunuH9Z2nuPhXxgyQeGC2g7rXVd5W6r5PHwkuc0oL2CylJY0gHi4CyczUu
Q6RSSQOw43ZbpKVOua5IdD6S9NovG9LwGhr/NFbhDLkdAKdXYZwdgbdOa3UoMEyo
IxlxUbXOz7Ag+j3+d/sGzy8tI4esjrTBVjjPodNPB0bGBFTDJTfPQ1o0/ui9WHJB
95lxEv5UxQLTb4fzD3m4D7Z4Bnr5Gw5S/pwcHHB1KeiHTZTA6GJY5GIQQzd20wNa
7VUYtifk6NuUsYL2bFZn0pS9ip6Ye+4lavGXIA7lHj3nPl1a3lTR27v2a+VIbzUB
YV4qIW0hZ2vCX9Coh3wTrE3DsT/cafxP6/XF4VkZXOTWmyZd/V0LA9auOkqYH1JH
Gn1aSuw67be81BkRXv+H+/7rtqX46YyEaFhRgSoueT0VqDdmPk+oK9j9mF+5BG7j
xLANrlj/bCJwVssbYCQmBXmSyvDzkGU8dw9Stt9LQBNWNLJLCAtDiZqCG81aX+CE
GnN8LUpiNzrjtoNDKcYa+uPGjkjp2G+MBE9N7tlVp5xCg5qjZ4X+cVWl9NakIDw4
Qcyh7m7hfTT/vPv2VKeLPZ/DVwbQeumn1N/q3poJF56UxNJZMSusCkIYw/kUyHIe
2JptbKTFlAkD+1jN0n8Kw4PrMUfst7w1lcsK+SCkOWXD2FZuO4BXF1SYmsK2hc1U
6fSa7U+/39gq7HfMGWgL43Zj1kto4NpN5zOmK3ThGGhu/K7R1BNiABbW80jFNWb1
hM1c01mPZ6f5e6iMSQ9bMa76yODow5kPn+XHU2+4S4pIc78nyLRydH/nkqB1BH/1
/xNp1CO8+cEFkKXugtvUuSF4kGOP1+76S4qShv01PB9njom4QWZJpXQSyfYW7quE
DnEFo+6TAn3mZ6Krzh0mWW1zO7Eelj3OW8zrpLTHMxOmpwqcoscHz0Nl52bcz3d6
BVoEByoctRR+NBGq8WcCVCOUK5lXiICrmgtbPH/lnU4VRnlNO6980sKeIRbqjiQe
KqpU8MfIz87G8FtuQXVOpr41CqBEkZ/IcgQLF5K15EuF8yT0+rnND8GwJyrWZxoP
E3hztO5uU6PrlT7jmVF4y4a5y+S2PusxA5SEyycyijCrj7cZwGgdsUfj86xPsnUX
bVn8wp6/G40WbcwXF2fWTSxngouUfakSuirHdrJDytv7yzo0dYzn9C4b9zsI5FX4
pDCTuxYipODtfdKV1VishfYtTLP0WVllqNqV0/xBrBWOFGpXVBAPQ9gwpL1IMLra
jrA0c/+N/JhR8BcWrQ7iFNlWhRb6NaHvmIKGHWXX1pcMHjrC3JCykK90yGLXWn/5
hAeryzIo2Oe3Gla/ZB1YrUhUsuFhPDRAMP/mH1JqVUTh3e4ZDsW56Vsh7c6vZboq
LG/AwIT4z61uFvfWhaJSjpxOfpScHAarb7OyxkSh4uXzPuGqin/2+oluQ7fcSfPb
zvQanNLkP+DYtNzZF45MZy6Lkmt7n5ixvMyTCVpiFsL5YzlxPh0wSab1XmlPvkPd
38IChvtuZlF4GbcCyJm0FevLfMj93lhiGeF91IxB0nqTNEQjDaJ+bUTGElaBmwgV
XdSFH5TxFK7/wQRHOLV8MMgT6aW5K+jftlJYDTT8gUAijhWVqb1UzSoLkB+AYoD0
rDjxFG7I/w+XoP8MpDhdeI0h97ng0WGTJ1ukF8rHeq44OPMiC49vtsszLqWQfJM1
+ka8yNH7OBzHMC01cOO7iEVUH7oNfs5xvLL/s/IdTZHxPUCZcKiB9HZ9i+a4RddT
LWuL8ze/kv7YsH937EO3Uxdh93dVsNpAGUuB1LSl/43at7yRfIb2eBL6vAM1FfB/
vEszIaOVHkogrqnT961a5gdaCGBgur07Dm/ZVS6iC2cK2tCeqnA3yU22hu7MhYb5
TxywP2Nh9KpozVxj0JEj89VzV478wV7nJsyNdqGl3ynjpr6Gn18sa0vIVAqJQSzo
YyIZtrYxNwPq6Q7kjMhpQ8vYqBDwrmF1S+tA8wxm0f10bEkgg76T4Unnju5jr7Cv
pRlrHzFckHLaI4LQUkqn5hzrqkswmdJBilxGlmcdQqa2HmbYNs04suNFXYb+55uB
r1DX2hsckCCpy3nUsmN1c72sdbH2SD3xC6PNzU7XHuYNl+qHgpMrQvE1hhbtQMuF
XfkmerYZkxwRqQhe3XmqsXU+Fmj8hExpVMtyeB+S84SU4u6NVNpwfgC0dx/BHREA
ite3fVAoA52N0ZT0vbKSI5fUQqlwS4RXDF44YHfFhM26C4VfCivl4u14Q15OBDrt
lo+OJuVBP6suGU0J1syLJ9xYd19fDl0oOev8qG/q4PzQz2xpOoKRUebxlOxVACvD
RXfFo8DXSOy4mJ0Jt9jx7foN4GDR12BDScDns49s76Jrlxnjpba7qjvsRCQZlHd5
wsrwuoxHiUYeDmgSzzHXcq/hwtcDVfbphIfUANU0Zq7E8lcHAYexpKLrmkyFBwqB
tpJ1/uRvkPZH8EOSA0NXdIdlXQoOBeMQAvqGFiS/qSjish/Y1Dd3noS+Eek4NmBI
92EgdxZAhnInMRDmR9HvBaXTqa8tGWPjGfSSn1wX5inOm8oU1ii6o9qMrBWqJ2cR
NcXPi3YbGL83NXBmjGEyQN/b/gfjTtqf8VjnLDBrq5pTXSxQXT2cYkTQYbmebA6h
0ABRjrXJK9XLstt6vKgDpfgp7AoEBsaiw8mVFtFvG8G+epWO3KH0n0pjetsgZny+
WOSqUKYjrCPAprGlKrVywvYTyw82RTFezWCnp7CD5cYLXpYoymGdVsCM+n+5zOpX
gJqiHXTjn+3bTBrFD4mGI78mFGmFYmYDHhIWOjAaZmctr7oKbItmQcplV1wALZB5
3+5xb3B/y1W3HSFjmlgF7Bwi+Ao4WjMCEdQO761CcBS+EFnV3pC/D/muxhgtAiTp
VynQZH7lyxixq4vFbh9Ba2PFN0/j4gbCFzhjBm6kPnH/8dQOXqxSzcGL8dWw1bw/
1iEcismNqMOOHhpa99MmfdVFCalpTh8m2Cc8ZEPCNLP8uWAyS+RdIzFLMeVbEnqG
v2eMNukWrEpdHcRrvlodhUR7KG7LwTnBi/Vb+5DipI+2xIJFG8Ig6eZHR9iTprhQ
Xm8NWubJXDSZGI3KMKTX/ZukIA60RxnN0dibT9tMKY99fZ9qelh3zOGlcYLUxJOq
2LAYQrJvWPQ10D00GkMsNiittUdSrwjJqO0iqKwdhUP9v4fQy1IgpcZel3nZc1uP
tA9hHfEVP7gOw78s39dULiRje/cDVYPDCfVPgtG9hDZQqW0G08GDpuJKeRTsa/id
fjaGoQDqk6MacZqB8YvWj/DEciGhJI0oRvEq0uzwxFvJ5ehaKCLcRrJ79SmKnEXW
43H6MqlKB5yIunOtCsGYuZwvFpuwXUd5gixWTmWutLN7fLi+G07feQuaX0bERqMz
hZXnI+vioueZhWnRVNHAiDtwOh9Kv/IUpGPQo8hqB2hh2x5Ph/KBfluoiGuao+7x
jcKwJOpnqPX+Jz837Z8rI4uAshOQ/hSYTF4YMBsBvtwLsqQ2X2Ggm2dCztyFUhuQ
1LhM3E5TOsXrpub7xUv1GzgGuFeov6TiabLP01RmVVDh7JdLClpLL0h1Sbn9FpUH
QPymLWg7nIR3PyampL5Q6bbyPJMZI+XqsAwaJNs09hm+6T27kRkgCzCqjA3RZRZB
q43MdpsCo6CDwfR/1ww0TF8E2kSejTaoDv5MV0AJjPNr4y2bq4NcOq3xU/cJTwwc
ISuVK9B2QjYW9DrrB9eU5r5ABm0IY4jKLEa2+T5EPqJHGrqtOimnE2ijNJL26K8s
yAQab0O9snsNtvRUVHPtnIuCs03QRyE+xDDewCA2bvkcyQ22lt0N7s2KY1D2B0yg
HOPOSNNSNEcfJ80QQF5Yu7YRItB63NBiiCWWNLBlLrbMsHkFWi5LkaPwXeT6n9Iu
eIiZiCC6Z9LHZfgy4oIfC1txUSzUbVvFPKFEbH4M2X/9HcBf84HcCCB0X7Hs2SPb
S+9ZPSre9louVf3jp/TzMDoByvEZUSt9BeFYcjF+WBYlRNQ594xGrmNjL2EqA+OL
kgmC8/XNnCkIobg4DXO9g0i9kX/wFR62eOJMPN/ZY3r8ma8eGd3smKxVjA5k5WG1
zIyBvXL6BnheGMaEvL7rOkK/Xg8ZdZgOBl0kK9G1FJ/6az6l9kIlg/SA7pUwyWJD
dlGJh3kJkS3zNyaQ3yvGYkh3QY7N+PKm0Xq9ss27GTaOc3DICT6BjFXRbDs01prv
8rieGJRGzdcRgQc8r00mYpVXzy13imNGBe7oyhvzhfrRrbTUzQiULwQec8mPrG5s
s/lyrdPF7MMnQJVgzySdlUXMsIPwsfUI7qBYQ6efd3ylLtUYKHV5jZnA0UvBzYZs
+0rc//X7zFgNIIuByxVcInMH+YkbFHClVYH3pyacC7whNLTFftu8QS9Bhnf4PjE4
obhgsot28CQav8cr/Ozmd2fhklpGOHEcYIpIU8TDwkVcqHLU7aMYqMKkoSODc4WM
Q3E7t15FePzTOsUwXS2vVHhBZS5REG+JOPnZsDFNocEHc0oRj5MAvhCkBz7VYHp0
xkpmj3zPH8f/jQDWGyIjohriegmQBGji6nBNX8mCq9sfUq4yDPy9lpjVu4WTOwnA
0qBFYphleySNGdYWXwIMX6fY2D4KrqwHTk3Nh1vXgoc5+H1vkogFkrnUipYoK8Xc
00YZZDuHkLcg7rpXs3ooenkdq1EqvJRSCLnQ9Z3jtw+oMnUj/H55Rj0g1g6TLmez
O7xwWVJsLHJiLZzIPogKpys8MFwYxi78OcfZT4hlJWWr1grB0HgGfX9lqeXYGP2y
KLJ+nmCNDSUzz4ETcB/AhJDujgKmpMIBoT0eTMNWZ3jylTr+iVY7u5GHXQ731AJu
Vb1FbRstvHVTgyye7LuS0xPG5PCl1fCfynngLybk7G0/bkBuSbwAxQVCKOK7EJKN
zul9KQJuIKL4VisQ7Yk71e4iPBz7bo7NJ7crwwxdPRrx/lrGi06MIKyXCnkTLTdA
gVm3yWIIrt9vOPbXu4T2Ru+RgoFuLX1U6F5/MpBYQzVnMMlk6cysFoyk78FGYZHu
594PIG2CGHVuecCznKVaplAQ9I5bFQAaWFOpm0YA0h3sun7TOV7dcUsgud3MSMNV
MbrGWvlT+sUIpolwHc0xlP3vvOyCPT/Hr7f4AhvrYNI2AdJ4m7KtzEs5K41dPj2W
aBpsOTe9cE4BF0Fyd8LRaRjS4q55xft04ZsEgr70hCfprkceQ6PY8Z3yEKT5gV5z
9btA8HuzOP9Lw3H/hkeGkMAIBJYA98+5wjdT+D8Wc2/nhZyW3qxbsteBdIWYxfA6
KUOAfo+ExKf2YUSWI52/jlJfRZTDACQZVNFYa0DsPcl801bxRKr+Ldi9oXmg1nyQ
MosdPT9/H7ff6BfrIdA8tjBro1gkAFofVysIPKacj+Zj7rHo7qYzof2ulBJDQ30K
o39uYY69LiFnCPRa/gTFloT4wAlA9sONiOU6AdpBTR+SHxxzh5Y3EGhZdBGMEBGG
UkoHhaJ7+HfjRGqHTraYzJRRT3FmqMURSh1H8H9kPsycbGnUSsWio2gHj4aJpeHH
6RgKIq9VXVi/ozZO1x7RW1UTm+mtXAr7ENx5xoKTJgKcAZDZjVhmc4HuFXEnOxgP
QLZohY1FePUpGArHtkXVwTsFx0RLX1UWTxBEF2lSEctjHULAwpHrk74+y2NN8BW3
w76gOmC4CwAtiUrYDTZq+OTfSQZ+3iw90gtB83qKwto3wK50Qr9mIIAopDEb0VH0
M9NQghJbR8e2Q+fegAJ5CLyJNuAO1/8Luut3LQvNlfX5/7AOE5SkD76beZTc1FIm
waXJfOaZeF+dAg3q/FQpY4DDzgkeqJAriJvKKFLcRrf4BimbYMWM0SR1G5Q82rAW
kaWUGe+ruR/QhDTa8fHMvssvrO6hCmrlYTMUdOauhTyr65zWr3JZkCkGC/bLSfyx
M6WQAN4P1rfAL+Z0p6JWxO1oHlUDz8BgsC7GmDddhTMpx0ND5rXtH0cJeev6Lnmt
Nrntz7cTZmitho2pypOIffQJp0vezS2RNWfCzzXvB2fQMVTRkOnTXKgCbNdfnAJK
4Q4eh7y+25hmyIOrbWg2bxlE6bMKrMZes1kJfMHrKOJCBfqAQsnscCsfU1vO2Afi
NE52/MA6kAs6lg6TRK8XnCWkZVItgtTlm0ru7fOYTwXZc9BK6skYgxw9++t8kIeV
4MlQclZdW9tK5deSgWRWa30qAaa3RRcLLMGAKzvtlIHGC/PPtDRyGJ4N30p1oOax
n3RPxWVX6aDQPuiB5ZpU9Gz3rNSCrDzNyzFqhiT7paOyACbRYq7Gu9y8XVAUdnmg
sZ51BPgr5VAwbnIcpXDQJ0nqmAnceiXNwG61LlpLJvOvXqXMn+o45cvt3/mJyw6w
2HDx18pav1u6e9vw7hoP/GIHsxY3NCJbsUZH+04ROqej3h512FDc36G944RgCuGe
DobefwXsGwEr0iUZiTu5sLTb27tgQ6QQ1mXlPgebY9pLpJjjYNK/GKRvM6mccmdG
nhlnVk8YYHyYZBNBcO/QEeSwJ73X2KHTfjrUv1SNaJIgNFqgwWVkkiuOtoaLxMFK
u/RMfIxbGTrb5/fiIXQNGZl1VXC7YgRPJL1S0gs3KT2KjRdO5q7gOkSBxHuUJ117
hgyXiz0oCaxJ8wgLqMga8BRgDTcuSd1Q7ARehNo0Omfr1AI/RPgJ1NtCB70ELh2f
8EHCv2K9c4wZCo85LYsAgHEhZ0nAbkxm97doCJzHiRyvCJCqs+rRxzOqX7d1mhrW
EWTKyMmKVwUKTNUXicDVA86uGoJVNR+7yYVQqn+Zu3GCQ3N5/PvMusB2vEW29Rnx
bYdu/In8Wp0+q7UWX2M1XWS04jA0jNuCnusvBA+d07HsxoKkjBkTyskKlru5eEVP
G5YMme67H+yjFCdbWIPmMoLvXmDRuxcDVqYcltPkq0DydVVSCGMQeE9tBCq87vWU
geBBpy/rC5m9tVgEXBTYaupFWi2shZnqJ+7Ep7aFGc6V0e7bjY5FZUb3nSRMPsPB
Hhg1I98hF8185dqS5OiDlHgSS4vdljGXTu6Duh/4E6r4vUdxz7xg6lhTnuaEsBGx
JdXQKOIDO+1aNcn/8h2zJhyZyfO97L6mKh/tvfvQsuw7SeCjS082WqPGvIz3Hp93
4KYXjR3LoqI3WzV6/6AFSBnOmRmJIVogTPNKWbanKDu+LtwS3GPN8Rh0BChSNYI6
2BDlZdqaSp6biTJMfvwmrbzPYmLO6ERpyKN51r54Dt3R51koPQzNQc94T9vUag8v
w8d5pdD9wijq3vIRP363iht0igKKBmw2XbJ7cu/o/3i/NpyvR2hgDY3kFQbvTi3B
ITMGKOkQKPukaPIOmxNTXDKAhLFuVJYKVDx1Ybk2uqOnItdXunGgbYZ0DU48wx6s
XobJwdzL/DfK/VJ4ytRXJzjvL+vmAvtD5O3+dvEgi6h7NdDp64EXkx1sqgj330sR
XP9L2wCwAEkK4o4jVtPNLcg3BaF28SDi0SifiwKCN4A432OZe4ZB7OTPB6CnNM6Y
4fT+k/x5f42CrFvW4Ai/SxkBTHRuBiMrgVoFuu2SXwto4WYfTrB1GQ4CdpUgIFaC
cqtUAQNM8BZHYSte0McFI2wU4hYGXbs1l0SnFXHSRtz4tJv/FfBcIp5mKhPNphWY
Y5TN5xhnGx4Zn3B4gtEHbK2yTukFhZmvt5Ek9V/kxK89cFca8lkEJwpitLYTRojn
YnoWdt5BNz07rHjgNsB3nZVff4KW4MSPO4Quq/QvotVHqkzxflIrYj/PwjqLSRCE
FK9Ttbru2Eo4Ey1NrXToCPDAG866nBnj9/D+A7/Rp1ki/jfv1zNwiirOJBZ+vJj0
ZjKm8HW05sN6hv0B0xVVUhPyr2lZOq0BqhOvb+gse+ptBqySx9nlT5Wwvf4dcEnS
mZP+WGSidQoKSFuuQr9AkQAvAqilNibAWfonNBL44aw8dYItjJ2AbFZOXzSJYVS0
7J6T+j2yJ55mBUPTrsE/DjiPEQ/u80e4KvthlewBacXzNwmtrbzypKEtgcYVlfNM
faUQkqB5YRnWo4zcco2eQdezOBMOt71RfuqgHV1kd1SNC6hU42eFCGClk3pP8G9V
HJLaHh5kVRyogplskQYMrGEOm7NySNMxAJcbdmEDudp56LAD80Kc7Lkx0TvdFm6l
iQ+uTL+0jFaplo+Jx5cioRpFZh2IKlRLE0m+c4zfOG084NN9fzzXFDPvQFennwaY
ddst9r9a9C8cGiWQiJNAumDI8J15MrEqG+n6l6xzHEnNLILa/3vKHXc6eMktM6GJ
9iurj8syhc/ghVfY+hZyWcyihvLCTNa6S2FxCYznLR2iu1wUvyUvLpBZ58pg+k5o
b1uhYd9GwYn9e6zbBBvKGbSFQh/mtByqM5NgOiGJ2su0KwmnOhrxB5tS5j5zCazD
qH+XIuq9cSC/Qy8yEVX/DlsgEOGcPBEgAQunvhX1H0cjYS5JU5IP1CJ6ZTvEh/mu
fKRNWLf2C9Q8Ub1TW1Cma9Go2QpAyVFUN/emE3cBbkao4ieBDYrUVXZWYqktjUGZ
Suc0er1oO0zkbR2bxxDc8U+DuIkJ9vf8NZ8GdmDcQ/hCQRPB5VPmOMtKQgjV4RZL
fcBWtVtoNxOknfe9mRhq8Q2SACRs9jFvqRh8R3SCP8/lkNnZ8FascAF0KqPJ/KH5
W/mnMzMruz9ZLifQX55d4rjqobTjvxxgiNq/LEsJhfN95P5Ph+aX+TqMNpLF/l2u
SmkK97nxWKSYBYS26wDWcjAvtvKpZO+ba4Ubf/g1mjlEuPwMRMZefayFnUXyHrl9
bm6uyDs7NtplzR1E8kTioJu4gN7Ty+GmTgIII5e/nc5UiI9+d4bOxxkuchKe64m5
ysZfGtrWT0ftRn0+uykILgwJpthjOvpnageTZmKpQAw9uUEHhM74wgvGxzg41+4s
qJwJ4+aVpI649FRPHpWElKNYP/06aaD0vYJlWRHKtmTBCd4tjnPuDmDM3Bqzd4Y4
wL7tYTY1Sm70NzemEiDRYdq/qNRVYXEtpsxmq1Pu1d11U2lk/LwFZUtqvcN9Uv0u
D8wlW6ItHKXUDEKrh2ujD4hmNAPGYz49brTDxDzNm6tpNFs2ItCfhr83JNmgycbj
eQHZHBrpBgFKehaeRpc1VcUBBobSgZ1nZHETZWKyK3bXYOcI4iDzkrv1IAUmhJXl
NqLDHgSmP/2ALBcYijMq1d8hb7CjyzSGV3B969qfGAhCjMoS+trTOcXM+6ohqZVz
leVOIBT01zQlBvO+5oVxx3eOaPyO8Irrad0UXGJICcXFFcNau9R2bPXB1DDaZ9gL
WH0KrJT/w6Uf/+pob0qNtWT3ERYB7UGrxyFyYgoc2zoFKv+FTgM0wIo86sG+F+FW
UMaRH5lPPx1MmrHikPFdU3R1XTepTvmW14y52yWq69L5n71HX2/3mA03DBdPeADO
ndrJ/i5hnmwVVMsj3f8dV2iYpZ0MFD1VWMpH5nvDbhFewli9j7X1ajeseMsTewfo
npHqhP1DrDulEEwwqv/s/8HXFXioMcvoCURkgqy7rEzIs4jdbxh+s3uhuD1fGlLi
JVDasJ10g4zSDuv1PXFCCRKrjsCukJPy0XxlLCPz7Hm3OKc/LGoGZu++sTD3A6T9
oW4xKQhD1jEFLTk56p5aEd2AkNVHp0bAGxcknGv/KgVjYCIk3YXFukm8+HWlUoJu
NA/6wimUjQxZRZDG212ibkYoI+4atESE+aQJNelKuv7BucxE6Ccg2yGQ8bkGyFXH
uXklAS0iGfOzClupPMHoefdZP77NqOoVf073sIrQupUOiebCSyhhyDUfl+p5Kgso
xvfs42nWe7DfS8h+csQYrfjiHJgpDcfcvEVHJpRodJ7B9lGYDWIEAz8NQZIDpB5B
crS38d9z8Mcu48ZsoKCQ3hugz/Et4qXtKhG5YdE8BEFvr8G9hCg93/9Ngn+F+1E6
1kSAGdfIZ9ZfkNmMdClcT0XhGNAJrCNT2VIiImHsuSZrVm3oSchnOkLbl1Deqn75
oEkiXhlLiyEk98PfnZNT3I6ard+6lCg4dLDL/iDC9U2FHqc5uJy8q+Hgm0MuZ3WQ
4Bz2smxtq3x/gPfmkUra1sx1HleJ6yDRdr90C9UpIcZeVucCvO6nHOOy98Wo0b01
ijluOeqHc+o+dokWukV+HUerHYN7ZWGQwU32DHl8ydJ75P8Q31wsO/okVGJ4Yhei
3lBAdwqxd593A+JZJlcqC6LmFu7SUJa8XA2Oz0Z/fJsixCy7ZBTAnv9ISzaf+lxG
sgnEubsmFp7blCd4FPJ9i+r4Cw4kxOChp5BAcqUs1W8nEpdXw3A3oXGW3FUcPtSH
lLSxvTBaDG8DFElrorJOAJBSUVahzFAd42fvILiO2DQB2Le6hek2ReDklFZasruM
i6g6AANM10PbZ93pAIuAqdLTicUWCcl8PApCs3Wzp9Yi5W9Rr4kpkPMM49ThzmFS
KRrlyyt3IG3q8vwgyfow83m0LWBBKKjHHaxbVH41ikEP3TrmSp3RAefrzSvMPrdI
tXKAhpI5T6N37PGAcmjKtTPFng7q6hkR6DS77noppBmpyBmr00k8Wt2nGEZZ6I5E
bvy9LaQZJnUipaMY2DGixjjICwaG2nnZ9tW/BdoS0BJbdlYA0m5VRKwDKtSUjba0
S98j8H1BNuoTn1XlSENDvo8FIi1JN1OVwH81wPnqUVhUczFWAp53rRNtGc6YeDPL
qN04L7NbbsmlvaRZEpSKG5ofsMcCMIMP2edxwKq5gYGzvwDl/jBUmClL2D9BituJ
iDmSPDH3KVwIHkPraFYGMrQtZFLgF2IBDXtsmkFRIl8K+qgAfrvK7NDPZbhKGPpV
kHH60JO9Ss+Fc9HPtad5s1Yebfj4QCWtplC0pFZ01D+2++HieObiIyBaph+WvoCA
AFEIhpRTg/iEncRi7w7q/roE7l4sKY7B0RHo1AMTUNNCwgajbuBy11OSr1v0T2XS
nCfaVkh/+q7yE0ip1BDaIWe2FLeZfIUISK34TG+/TNrzUeI0wnX4kOfeg9zMSj5Y
1hToqCjTKWLf4x87/tjBpJ562IVEh79QQOfevruU6wtUngoaydjxGjXUbYkuorYR
1tobv7+gnOjx9pofXWLBG3KfQMP9S1oDpASuRSZGqxxvowPuvscwmusZCYUkjwg+
+3vcVC39Ic+iBBkMUxMQmmwQdCK04YtT6xZWsHTqr7OVSjlBoEkRSP/HgQN8RRBE
h7h/sRvgsiYjoxm2WiXFYeq8Z2cHvgQfjxOtqr8KpqlHcHadMtXoDzauUKw2ldpo
kcfz3aX+jW9dSyqKhIFzfS3bM5ZcTg/WHaWnmXwp29O1+yu0enundnlTrLS0BC7m
/FR0XBAMFyA5ICRSiFSZ65TtqVzjMvWtb9Xiwj/H8O1zzBCr3q+dSnhj1xLvQ/Sh
CbFgPk/RlAeasn/UNv2fhyeOxZqtkLZ9O4TIy+m1IP6jgQoLVQU6m1/MhK13Dp4Z
O2H8/CPOMqClLcng3v7QTtb3C77cvyZ7jz21oZvQ/2csAxybtRERKFS/LOM2K8DZ
E5EPaY651e6+i1TDNCBjeVTEAzChmStlvPuD1HIlXqIepXekV0ckMbmpPiM6AbpH
EQTlTh/OwixiCbMEhf1+lcckYCFqvhPM9x4sCKMinzKFvBySzYvEVVRuNNTHyzG+
kYw4oKqX6mzSTBZFWjDfeQq6Lc54PPl9ehEs7DnDtLOV6ZVATXY4qt3WAWbNHisl
Jr5qNaKX61Vb7Yg8yq8QvM+JKlW4GW4gUv45631x9Tfk8NO3j7VeGvLNopWHPebV
v5Zl3mTv6Z0EaJRV9GohkreGnm4XVvBFC6VD9co8hWfVq8w6Brp8n0zxJYxkzYrY
IyjcNKIaN0srLW9LNEU+vgOq1pIezStyzggOwbenDemmiUoWPws8dGque4Vvo1oq
gdhEEO6Zvqq5wdI0UEwL2g7wAX6pOOKR90vxSLCreOz+apeuwvCABC+DKZ90agm+
yU+otjKFXg+4DF7oKUxpZKxv9lu+V1UI0AO05fg3VT33G/nT36xtmfaQM+Pq/Sd6
59whyoQaJKXkaOAqf4cpTXueXnnhb3XUnuEiGgzYdn/LtUk0auXaEwBZhL5twx8/
FiG9/p6etguaMbHiptDc1DADwBh3+cFKk9UQDTiNdet8S21wwu96+GCjs5j/Zdaf
WYnjaEvOldYOE0aMF2mj2bAi169Q/5CIPkZsRnMtrJErbIvJ4UviSpRaeP1DQRQ/
/U1U2R5RZpcPbVwAh5DZ3gtVeRy8awf+zdQ+jMVwtM3Hh480KtpvoVOFp0XCIc8p
yxnZa/kCrT7RmFbQ1w3im4S16NjE0swrojbCs1pIwcx520+5TzLET1azN4Ofy7lZ
9ebIMxkE2k90qqRlA6bwb0rdJMvuQPkwiPCTr/swirX7l4172bBxWzby6PoNsRxZ
jK8tOutSfCS9hJZskI+hPxg2DqDRKsFlhgdn7bgI2sNNfX343e9B72R7P5/BdtZY
zSHTH+qoj0IZwqcWLWhFBpqTquWuz+cFYvT5igVxuXW4N0Uujp8KkUgATFPOBTke
+HZeClPdxHTSIzcFH0xpXQcSgvHAohPq1w+X41yc68lT1sAXIEBOZCz6pDOPSvhh
kpdKJ1wN8IWDvvkklwtb51YPLFGvT84JYz1lleIaPH/YKerDcGrwHczgOBd2RuKI
eqFqTQNOvuul14V8sJbimC84K9ON+cLP3OyEg2DfEBYYeZzm9e/nUhiHf1vw1/9J
axKvtvBkkZpmrounO19ja+7tg161+YPlvPywxUHQpv3eA1vQW/Rnrovdds+cEI3L
hKJ8SndANSBJzsBsWV0eUAa+SPe6Fv8kRzfo65Wl/sVcFpYg/291NWd7341wSF4q
mq/0QPkpf63N4pVBzurTdeZNoRpnMbonNqGucqTfb2Y2605rMIX0Zya8Po1C4nAH
/S7u9mBuQt55Y+JAeV7V6MJaAjri+IZO2YmyNVaZeyfotSr3+Z3XkcxVnaULjEQM
EvbE/urtyzv2c2yEcKrI/TLrIP2TWyJrMcyeJLu4Bt0pnOvLueEn0iliAnx7Zclu
IxcjqA+M+6r1fWl5kRr8fiDN/Pb2RFeRU96hP1X4qUa0jEwKAdgqtELRoHyB+mvZ
Vn09/nN5s3q0gGQiQoRE8AvTNRfObf/bF1Qn7rep+zUfPTpeFvhRsK80+ipxNmIE
lbwWFwtExqFY1C2IZsHc0Qxre6UiOrjvTxl4G8VTyynHx0uSLawqOWGh/xVkh3cK
YXRy5xJEWsI2D0hQFpcHIb4+v6BrhsS+8Qj4DLYrUWBkgZSX3jMOioCNUsNsyCLJ
bjYt/BRy+5dnb8ibyTXGRmw2qXfCO49GCKT0IjZrmYJqTW5kX3xxTgNda6xWDq1F
ra+1IIpARm99c3v7Efv+se/zWlPHX5Ju/KaBjzBaLx328AAbRFRgXKUwN366zuOi
cluhQcILeC1UCIG882KbgJ7sCp+IUm2EX/IR8HFtCIh19rPGJi+tH+vIygw4j+cA
NlQCPNExs5uyfORGvhpr0ixnEtGMy8uW8I0hewFu/BoqJta199xdp0C5aD0JKHs0
1CtdhLy2ztSb92ydrZ4PhfolaNBIjryZH6WzGH1oCgzue1f9pbVNnfpoqA7lFVUX
QgtID8E9E7U5cBQYximGgrsP1Zyk/VzI0p62Q2ofOMzDjK8xNnQ5ob9c20OORrNS
7I8atArAsx62YVZcbFSLPrgYMz2XQ2xKcRUjPBrks7OKlkGdvqfAO2p7IOgUS6Oa
K7nr0pL+Vmvw+JWGuiDjMZBt3lEkKq8c16ZBO2LhD+pba9LLjg+HtiM7R7iP0yW5
jV5FDSyNTt3/1LYOMCmkaJp9mtpI8RegMI57WYjJo5oMBKZD8NHoNpBwkYFQfkEs
m0YhLYfB1KYypq/tnj5x/3HMo5pVakKwHcYR39lv+LocFUIXoI8JmWT31Xtj9Z/6
OdCNHPI0FRUx2VsVwN+YXpkeL4SAcdCpgHTWpL22babCXyQCodSc5/dLw4aA6VGr
K9ZsYrLo6fhc1CirHpsVxqv3jxTGWFfUyLFKhfmW2y0dVNsvf4aQghaLnTPtZ87m
wA2Tu7hvB4kDP9l2X/gqNRkNBIUsskZB/BNY8X16Ykq9i4jSjWAzMRQ/R1ln7KVt
WEB44Bbr+DrNtNUmsZWVNlAplFx5CKXXLxdmL5TxHwwromulSo4FwGLQsM7r9Swo
hosPRKJAed8xpJgww8Z+HiruI2tbHc+Mp7U5iaux0WNY/Ig04iR8B/3TW1m4D/8J
+Lvh/WyB8btGTgGSlniUBBjNBpJsEYVPj9xM7qWLfWnx9JtRuuDb25RY3W5h5+0M
nglk4/p2yO5V8QqYGuPH7gMypczcgNV7epMjVmrzJlKTuNm2AVtQf1Ec2wmY7tXD
2jptmaFzRfXpUnGGiA30f/T9xHrZrCkUUrj+ov5GW0tdvO+Iu4jS7J1ToQrrmjBC
mGv6JJMq103BsUzx0Uv3YgBTUNgCN/wG+w7jvE4cN4giSbGnEYX+LVCpkgxPV2IQ
MILWUkrcEGNyEoy8p+Ue/TElGpVw4EJBThfhufbGOwqzzeALjD6O8ie8uTHAvYCV
VMWfJSISmYw5aRNs0wlXJSyiJj2VghKoVhHJNFATZlmVak9oB8nFI10OwisiBMXO
DKSX8DQ0mAWngdYzdxAN5CJsM9Qy3JXFFbAydBv9Hk13VZRDW8MCYkSkQ4XWur0N
Wu8+C/T3qBLHc29SQCuInwSA9kPhLMqrjBAVFsw+aj0At2Xn+eLl9qogTHi6HV9h
lXFPWmeCy5szvMZN8q4wqkdg8aIl8tLPAl9J1kRM+ajt0nmwCCXfNWHl9Br1B9Lf
0CuRKQess4UrcXYcdFK7O6+9AvHOAQO6x3AKSM5OaKNkJlIMlEgeBf0jsjM2PIlL
AKf1YhafldSCp4ooRbTJtIQTZRxsQyjq4LBPYR42vQ+26R1OkZtlFI2nT+y8U9i3
Jz1/nUFPAwof1bHlmryeLAESZgewfHOGUdzk81fFZueay0nR3UgduM26RATuvo50
+c9GPF2FDpYcsieqWvZUQmsbggzSEEnGADoktbVTpVqXAdqCkfUZwiRBm4maXfKS
gh99x++C/2hPcWl2xj0NhCIv5i5pEx8VH09hVo0Awo5Ab45RmeHzFbecLkYtc5LI
PhCiM+LdlFYSeOj6pUD5OmDn+DYwn6zdhZqzU5f/N5V7ekaDt7Dmwlmr1MPIHJgy
OAB8pCnRt5OyuBKY1XVI2eOHfEQm4xqhWnb3Mo37IntJIlQzlXtchsfpuveggfiC
b6XNTyFFWnI0ztE7QihV0wi5sQvi+Fq1kNFK6FVeZJ1ydAQpohXfwm5WFDX99sfy
MP+u/cPRV75m4J6UhyiT1hwqSAWN+EtQFB/cbhbV01ZhmSU260jB0uhQUkPRjZ+m
BPn4Pby24g1g+EDr80YO6Ft4/C0spUpb3kO7qifqdADJyocTat6r/0XuixlJ05gI
EBD7ixSEUg5I8iu4r4gVBubcDvMKw5tDJ9j3kGcpoUaYnkJxWTytw0uVESQWdHo8
dshgCZrUM4vz4ssJqEihccSTJhb1CKOl71yxJNF91sXrS49xXyaGH6cncKVj4MdS
vnA63pzdqlxw/ZdpvROj7M/W4MV2ojFY2z8ZQ3lzBp2zPaeoDYfaYaGsr8plydVq
IDr2HUzFsQECJfJ6mN1YwpF7wf8DZeAv3GvQtQg5cWYzCM+7W64RuC30/F2YTOjQ
+AwyyyY+An6okfLrqfGyVk++kGUBmgXAPmrBVGVObDofsRr/fIFxi8HnKyIvmDWy
l3b+hwUKYihSfCoKcNX78MuzyEkDdidXhmzsEnSVTqfgwjtr/zQNdmbW+v7EE9eS
1XiV3W+Vi1X4EB2qYo7brndpBSSkMnbs5+x7igtFA4iCtWIkbZ/r/xaLYWbCUavp
6T2HLJLMhlpEhde9cJOlexGBkxfLHo4ZI9BKttj8RjvPlG7zTmgOIrYzGCPJiiSD
Atdv/kLkNhAC2B6L8WWRMGB9GcOyLGYobeDac6GMLhz43ysDyEzZa+0qnhyk70Nv
wWVUaH7BJeM0qb9a+t/jmaaJOMCKf36kpvAA22Wpm92f+Oz5cSuGC/LMBRd4CJEl
m+A5jsBpcqulSoMUwMNWZhatCET0PSvrpVyCsif/Ykl27cq0vdmCy/MATL+yLaO/
uYbLUyoyfFYP1JMorPODqCYQ4nXnybgz8ccPjxQl+3vm8iNP3MX7pMuL5cr9eaD4
gAQ6IfHBwJYxb/GmtvmWR2B9+mhUwJ1O3f3vkkzBM5TDIylWWNG2Kt9JzNgh6Nf9
E/ovYeT+BFPqKcLMkkHwZV49xrFTlYKQPsHcq8+0h3Hp9tvlRvCv/0Z7NIIUrkng
4QTH2efG8n+CsUby7JsgPMI69IUmm3h0qFtHWCljmw73rvAbAkqEiccU91gIQtkU
7LuXcXCOFTAPyUzsAzqJazXiEJKVFu1Ez0NzGLHC4RZnvVooHabiy2hcCfjEOtTN
0k1LHqiL75m6rQbipulML/sAN4PTZT9WKjmEPYfPvMgSNxrhwLBsMM0MRO2jEN2K
XCb0cvnrip9oQlM+yKD9N1lsHNUsk23CNPpzRbYC0bWzAyR2E2pGTMsPivrnocCf
Rfz0OOYGMy1OalAN9y3BWIwbF9iK+JOqaFOkkCRlNSY4XH/JZSSoo6HkT+Fq4OoY
lD9xJmlW89nr1QhxsNjqItQfOWf5YXs8VHKvrq8N7/BM0Md/ptk12qezD1tNd5tJ
WjrR5dap5Qw4g8XMNWC12gjSPDvjSRYZaFDAg2ARHFJma6OTB0PGZNC4JN4VV03H
X/sKtKBkpqD2Hrh0axgH4Qn71GMMEtDn7cAemxpz90wb9LfM2duHailHQWWauspb
IAwnMyvjXymyZmCXznNkiPW0ezieasDsaErVclXThmSbpBCwU5xI2mjEl9Uhn7Aa
FIO6XwlaCUaFrl19Gf30xQ/dCl20A4VnYV+GBwChxHWStVjwVP9P1Th32FztoRq2
YmkBsvmYxW1gOCoRUXKwBVYoWeHlOHjeZuJjIps4j3+WeUVWIdCW0n0DBCI+5BMB
i20F/M+54Gg/nY+kTcW7bQcK8Hy6BiMvmBurL3u8ut348oUve/lKQeAW/K/v0lnn
pB2v1WUo0kTk6R09rvcggkBpIEHxgA6YClHQKtTLWjcVnpZ8FHfWfmo0lVNuRwl7
Bbhu908S5ptSPuWJ0iUF57/fOBJLknso8cL62Xkd4RTHrTcIakO+qRkLDwW8Eu03
MQB7jbXRXoKPnIuxZ/41AJD4/Z412b/X9JE4o5sE0lOBBugI6MJE3pmbRgCIS9Av
NQmm6drMNZSI66jnV/skOehnuzZkM0ltHD1MpYdEAM93GxmfSQdITzztN6sH8Y9h
R48/b+BiFh62jtcayhwJneRcF3jHbV3e+9QFf4oPCdB64+RY20ye/sEm710VzM7Y
C4y0fJNctC009M5vyCjznsP2HtImgv4KFpr0fwv52sp9JU8wP1kAReepZMhvDY4j
K/W6XtRXvmZ2NSaor0oBnO9b6+5j8P36Y/iSpvFg83eISknigMMRBBdOYCPyJZrZ
fudgFZVBOpnNXwUZyhl8maYWANSO/SGWeciQkFo3T9dtp4phnnwtqQBdIoZ7WZDD
XIPh/ZOWj8+veGFT+SEIVLf1fIzFNAF9aGvWyS0UHIpog2/R3VrKKAas2+upr+v6
m6FGQm6D+FwJ34n6A3T+7dcymiY72dEsoikQpjPz4ZO+md+knOVEBhyWZ/JojI3N
1/KnMdswU/QGDJ+9Bbq3hQsB2ObCC4n3BeZ4crc3Gsp4qHx+FMZU/REz7k8Ol1++
a0mTab65SkgVepUlg7p/keFJxvKQIqCD9CnKkmL1jo0vNisH3UfIRSfP2kEv0nIJ
gWNYIZmS/8MatBiM/gt0XeSIeX/9UmAkYJEjmDlyk0Jr/zsSv3OB3bHydjD3GgX/
WOVTk+uB49SUSDhYX5ZpivLRLTeD2BwjcgnueU/HTM+Q6TswPtmT5kcMKw/daSFf
sgiDf0gs48Eyy5l6slx+O3JHLSkTsD6aanHMYbyIn3JnPXZUzXdm0hVsi0a9ChHh
fZ2qz7xOwNYmQwxhk8intezwyxLWYZ36lpXIykCbCP19embNLiRzeBMrV/Lcs/PP
WOmTHoTdB0ol+KaheChfGDsmA5aqvXjaOFVewU1661HvB6S3i/cBPHFMfxWApk/c
6x3j3qqJU61xrmI2Vz38iye6gaPEs4JtaP7Lso8vwvGixXCg1uhFT0Gcx5zhTlbb
S7Z2322Qsv30yE05kwd4CSA2fiWXHWW2+Uno5yowzW1YChyqHE3tB7G8C6JSuKVy
7kPvQQ6+IxqRBJAJYp5+QRgopslrzoUGFSHX9owoW8KxQ41acSci2TpimfbDClXE
ZaQ+KL5LfIhCAvSzZC5ta+/yPoJ2r/GkIXJsJBuCgaaz2B/mYdfUSFqsjDhzUM2h
rpHhhCZioAbBTGCED9ri6k5th3xgsWtxe2ZrB/WjCnjCH0SLW/YnCxoD0XJkkR1I
Ee3DBL6PaZBaSuNk3DT6eQHX14eexECsdY6WCn/PI/nz7x5wLpnzFWMEbrmkES7g
duxV6sl1JJ5qzKkCgpJGM8Q6bqoVcifq3NQOgA901dKies0nG48Ld4pc8M+OlbJe
dnAYv8ov4S57E2pqpY3E3hEA0qXs+S28V8Itv0Y2jcyZ3kei2soF6P/LmXmnprXK
scC1ERKB9mF0U8RJK2mteUkzRiXu3BlQHl7nWzGWEypmQQmpvcLV0cVgOg7JuWkA
pWWtxyrmddiXTo44KG+HKavzQ/NdvmWYPMRa45HzHZOAhHim0Wicdqa1bEDRjD+7
Mqm8yguvl437ZfkkkOa0QJNEWSQjqluqXIWfVTZwAzA5o15/fWEAzEhIAwtJTX+w
WnizoQi6Bxq1HSEJfuDoRDNck6LWerWCB4LM1PPMyvjrnjdiHm0SXJ9unP7+l1Ph
KgYfEtOcVhe5T5y67+e6hl/ly56EIgwxRfpSvDQtEOkzQzPwQxqWz8TzsYAeVkyS
2/C2rSkCOQmqOLkZx/BXk4FdTXDFNwBs+JgKFkF0O94DiL/ximt/iee06AXEJXz5
X+YeyHNHruMmg0QJ07YwjczpChZUdIVKBK8LC03pw1fhRKSPyrEqB2h7q7M/11qZ
eohBgFrlJHr8Qd7RcJZHo+VIwDWAFYo+HnouR7VQ9EXed3vN10ABcJxmxMe62b3L
AhfyVOPrIrcQ1pn47cmKgOTcYhbWHJhXlfzSymUV9Qoor3gw9Drtv/gW7ukqWSAf
8pB3B0+wFI7wQsexhGPr6mHufKUfd+MjwDAMs5d/4+Svql21GpdiRPIRCUGymfu5
oxyyGkvdAZl2kjk0/OkKa+V4ftjVCvl+XAMzzTn3rG1/DIgRyu1iNGTY65APtL+9
rQPE0nXnXfJ3HAlZNiPBVw/k4/iRXZCRII0i1RAYROh8hkvhfTgRSOpRIvRJfJUb
EKQ7aO9wCl1g8SnQxFtjkBaiPcrvYqnB0ItZ89+XslId/iZrvLa0hbC0waL6dsvj
05pocalUck6BdJhIkQSdbV7HfH76iTqq1LAXz4VpFhW5HOhk0B+RtM9gOjuGOE+g
O3fF3vouumn6kCXINLb4VAf+djZ9crjSkL199B0AkN/96pTHHgfPmi+ybxCvH+Ih
QyZyoB1CZjn/HY69QiPxuGrjOnqTpOeipGRdsCA6Msp7QmUjnCeS7QrWcris7d4r
uJDbfM7sLOArxvT2eyqvGgsNH/7NVVV9c3H5bGCeHZ0NPrADeqGyPLGS6T87PXYo
mQlCzh5vFE7eCILQ7e+5is1n+EncnAWWDim0RTZV+33bIOogblD2xLrZqhiImdqq
2UEZ/KgDijKwkcNn35dakwMFBcZloeNFR2tzGzXszO1qhmSTFwYCoUkh1MdkwqV7
mH6sPjsDxe7PaMfpdCNascXAR/YGAJhpaSJF984UhrO8Ukc6smAtg1EWU1oyRnG7
UHW47+mR+gfzes3gtQRM+kwgwJHPRmBRB50siOMMqd2IvGo0cp+O8Rwv98tjOFa7
zU9ps0gu6D39PUAGkF8qundrUTV642g4OeDbm/qC3135K8lA/GGFQxbup0GSa/Cd
53XJv7HiugOeHhbzW9bfGlDlO3pUyKNI3hzj9gnsfoj56yGysIix1ObhnXLg0itk
P7S6D7RQu+npTj6dH1rIrvsYBoF69Pv3itt759re/foE9uqlUvR7Ht9O3WPfy1ER
u1JPyxKCdx2qhbCFk70Iy/A6RoD6zuNKHoNu+FOQLLvkpIDwcAi7OgEc/hg0rRXN
rF+6rYpNOYaUwnwYf+AP8Cabj+lH4uchFRnGBZ1Kic3GWz3sGvN6QzRKQMt3IlqK
Cc7zj7ifb74tj+lufHVGr03PQgTe/+wfnHo0+62mJh0NmiYk0J0Nyb1+mR95lS9i
U8wNq95uIw/Wk16AV6NdjC/L7rjsOVHJNj1rnCi1mkWBo1QNU8uyXG/Px9V3mALV
xv0SX2zL5/OWsTVYvL6DFfawrAIqqUVLxAqSv9nDx/7ycB3gtIl3n4OjTA6XbjpQ
pgI1TafEsI2VsdmuPJwvmeD87kVqVedFadEH/0TRBHqURtJ09xU4uAg5z/ZDoSyv
DgGyfASShIJQQRIm25qd3e57+YXD+rv7BYTkiLWY8IHKqxocLrCTXa3qKZtRnKc4
i/tbWrMReJR/BvJ/VtLQP+34oTHrxqTVBi/YgnYkKqEyIRmrnMyARTPsYsyLmhvJ
mC7FEBAdbUWNdbcpa8q0d4knsWHK6oO2ka0lWuuU1o4AFuaWoi4Nmi25R4fJT3cg
bGKHwIeN5X4gYVXNOzrBpIstuQFbPId7CftOl7LAs1onJr74C1rPRVfgHPxe6MrG
twd6UlNL9ZfNBovNtA1OBKpV41XzFWpD7XrvfHgkOqpduG9xtSiwzigrQZwGdp6k
d2fCuMGX1n3028Qz6KVvt996uWjQGAcPN0fuJEr4UWFbQCiUgJPhcHCq6pPdm8nO
PDLiuUuVvj85BSiyaOd8iWse4eUhy0U0dSMRuH5eqkJ/zoD58h1q9oviGjgxR8Rf
NFW0L1r0a3CuWAWmho6KHjMgwRee5Ujh9sO5aoGuanP/CVi1TtakaLWPnYhwApXk
TCPZLp3+scG2+qPX/PBzg+zl7Qcd1VoJYm8ERQjpPXzeACYZ2yvnsjEoioz6eqvq
OoRYwb4Q4trwbJASfJvLIzGU3xEPXXqHv49y963CmqU9Bxh4TL5u8MRg3tW98k98
58EOkY8v6Qsvisc0OvwHq9X+UzYhS6ou5/anQtossCV5GtjoL7VPFfumbwZYP1hL
88EwQUSOSPoSgmPtGMMZLsgVfbtsAO0hnvvA/aNH6Z7/kccyiyQKvQkVfB6sLGEm
QADX5rrWklm8DoNu+9KnuyuROBR5TVJdiCgQC8NMNpN3VjDMuyLEHsPlon/u0OCH
QkgpnmsVmWQB7Q1X62grxAWVzS153WLOax69iGywYaMwY0O45a20cKIoOSX+UW/F
vmi8AovsfnZxI9l13ZfD8tpWxYohC5oVncS7GzhURIVgxpA7GaIae9cOpCYV1Tmz
PG+AXkED0PUGXWWYT2myr64FtBcvRUlYQ2dgCFaKcT0WixJ1xVMqrKiWTYim2+Qt
K5xVFn2TpfXZJ5Bb2DflWyH0W58I6glM9qFpMg61trubYbGT4Ci/OpyYNYAdEuCt
xfFyE5Uq/Uav7dBwEYq6SuWBJ1Q7YGbWBkB9bCloDHzXFw0HUsDhu8eXHDgC2w8Q
K2z2aX2K8S7VyZcsaCCnZZNCewvIdloFsthWVlZMxyUA44+2uDKwWGKq22jswQ+S
F1hg/3FLh/BTeI5M/Kho3nq3TUFuqO9ARNg1VO2MS7EFWsX8oO9fejmb6j3h1Hl0
YulwxTT0IbzOfBYC46ziru61LnDLYMBtqYEB5w2p9O8ijWlpMnwP/IPxrNzph8jw
wVmd9WhNBmjxCD85XAokLscEJqVCkK/cqlcZNtlC6eppiENm5zu0oSojXjWCoHUc
XuKW/NUKZ28nhl2ftuY7ilx3MspovgfZqfv8om5valmQ8hiaO8PZSIn1JOYm928C
QZOfpuCDSfoTwZzRFHfXAIplBCrqAinLZXW/AvwUcV8Xvb7zWVDH3kyxa92k5uiy
XT9Fl6OmxaCH4cNnj4xwcR0suwEU9Sp4209s13i8/sSYl2Av+j/L4ylzl7qG+YQB
L1LjzlxmZ6lS6WoAOaEwZfrLUVBgmwkRIuJaBZj9cNzUEYZCfRlxp2ZGHnFB8mwg
V6g+EKDaZpdYR6OyVkGHJFwHFlW/1Fcyb/6TbFyQv1BRE/4wa7Xm6gak8rcWcqL4
eWMZZnmYDZtsSEIFcpfX5sPIikNM+h05M54xGagi9mqabtpG8iU6xQ6TqdnNPKti
rtJyjiwC9QbxNXHGqhPUEO/PcqvBVpHlNp8uFpHnIHev9Rktvfx8JZen66zvOJTx
VpGlNeHKfqBXCVnxIcLy5ncROLEpg3l8/nfZsPKluDyUcI8w2ZB2LmBVYZZziKrj
m5fvJkNL16fvnGkaGwr06OdyMXGElt/hggvzmgX79qvwPmEcge3QYCSQR6U5dwo0
IncNxY6TiaGNu3tERfmoiapBBg6pl8N3Hh8gpoc/VdFDN0ncTEqMa/ifv4pouJRj
9rI+FifUf0LGvXyMsPNEUwV0sPnot0I108TgLC1ICYpQtcYiDzPzL7F7KUt0Qzjh
lxtP3pb9qorzNu5aWeKphmL78bFtd7AOhBQc40HLiBqwQFL+OnJHrL6k18eKmUlC
sWaZvuJ+52NFC1ldlVEWaX5jdwHjwrTLx6Pu/agie0JuEtd8D5xZ6xMrggdO0XOT
NAdwlDYPBOjWF53A2hsSv3rjEqyRKZmHKoDaVxtO2CULULS6qbnvddPk7pWfX82v
30PQq/YuDM5KR1Nyr3xAIW0l+EfQfiawylME4zAa5pbJD8T3sheGtFRukVaa+WX8
+eNgNxEbc1f+iAoiNo4iuEnlirXU3pSvTahH/3q5T0GyQP5qAB7QjAKZDmn1cdzJ
3aIk1Tlxf1oBk4Ft3O+Wk35rFniNCxWQkJd25RloPEtpVj2cEj4ybFl8X/msVBeJ
h4xa68TOZhXgJZuEG1wEzb9ko2cy/1uljYEE1sshqL7Yn1E6OcABbz76Iqp4eKTv
Nm+SK7aq6NOF4d168sB+N1n06MHa0TK5B0nqvQQHCxXkhk9YHRLPCWf1cbf4xxj8
pTU5tiixIybakVe4dvujXE5IyEQO6Dm7+jm427Xa3hFZuho99WOHGAB6z9BWjS2S
uXqbYZg6J5EebLhw5reuZCRVwU4uMhduUyKm5bkWuX6w3DKG5TNOs3nToj7nry2n
U64ggw5Ya5cpMBk8Vo3NHLksZ5SzjMut3Wo1ouMIuylhRDgkh7b12EPUeCa0N+RJ
LivQvg6cF+HKXaK+/cPPysmYioINI0O2jCY1ikuPGpROLbfN9talZFRexNSatd94
1lKyVggzG3yRpr39jYwBdpLitq+3CMzdyfni2m2kUa2obSodR+nGSB9tcLrNwIOP
Yj+m5VkrrEryozHINDpBSSe2AD0mOO2kxeEesFh0X5NfEVp5yZMw4CPlWIDeHux9
wfKhpq8GaK6oo7r/uBG1KCgKQPWfD2dQAFLkMgMnoFeuwpbqhcB+Iz9F2ObsAkkl
BT/AnjjoxEZLpyNyOzo1D2NVYUXkBspW2e/pTKKHDWYf1hOv1/IxQpMtZ3zLLW+K
GJ/FwKkci2QpIMVYGajSN1mYoxe0pghdrBS6ZbPwQ9laD6u1MG+H3dM0JlriYNYp
/gF2qakAGppnKQtib6LVxZa+1vvJLuc4kJQet7qVrO3go6XtLV2ns9xbh5n6fm8F
JcdOn71CeHgTbras6p396tI8Ax2X4JMgAWWHK6eC0RlChxkMf+BNPDhqm8hKggoQ
PQfmUokV5qiji2vG3YDKSRKNABbpNBGsq1+WZ+FJaNIZbyPB9WvTXSd7jxjKVUt3
4fY63uV3x0JCHXozfHDZh2iuw9/wZIc6sO8aCdYxghaurlryBJT1PFro1HpuLbOj
VuEpASkitVsPJZGaWKrfgHtLI9PHo0+6G6ttbURdGVTxfplnXfm9IpFjBxnKJMxN
q6EylwuWVNCfxeyx+71kY3OowvA5YAb3AmQ5s0afvT3qkPWMzez5iqnH8jDQmmGm
AOPPF4E4QtC39lrsMrkSVsiV/vgCkZ0vZ6mYr0cg1so0MbPNyk7I5nJ6wqVoRTxk
fm2FhaTGwNoveDMJzrTw/9zq8E8j9Eo1pR6BOx86sDJTzPHNOBh4fger4i1YZq+C
hF5C43QF83AlZbD4EOcrZrRTbXRFzCjEyYg9wUtJ+pwVVZCgbdtXwouu5YyNt8kc
j9CSUtzwLnPem2taYy4o3QIziS5foA+H0KQoLEus/SPX+QTnyeEsF1VKjG6IK1sC
Qr0jRZvQZ1dPW99Y1jnDW3OOZwW3LcEneT94WaM5N1i1YrsT9d15uZBtK8yGVCPB
t9znluR1G3+7yn0ffyk+oAjVXQRukoQq+LL3FvkQ20nbqyBzxvRG6KBJwQ2byIjX
ERI9Tzl10+2xwAy67nG4KW9RWgB+NZUi64aq5cjyY+zjP3gmvGXSE6C7q/CtfRBI
L1pu+gX41t1nUWJ6Q9HC7MQ2MSc14iUvpgAAXE9pZlt3x9kRjTLS4yybUojMf/Sk
kxn4yT4EqCUJppO+iPEHfixB1lZhdYx5+r+Fwz/QpYedgIq5BzXhUEZI9rmLigF1
8eYucYY00Kh8sx935a8MDyKouKw52gOpJmFLtblovB0krZ7msQrB6bRdj3PJAaHK
Zi7JokcGhrAVEWBf9CDgfQ/NJjIiDUFj1aImCFcyAsdh4a/DrYB/GKEUObB9YVvf
UC4VbYUCF8zsWHngxP29mGvJfa8YTk66CuHzeLxd8k8wvqQYM+plLiEESOgqgz+y
GQ+ZOdl0ZfGsUIfTPkd4vnsIPXI5BfdC07OhW4ErJHgUakwgKxXeIw58FeTndfNu
Q0K8UcapebMnMPo6bfbXq8A5YgETQ02tMREXCVKyW9pf9fXsxnNZgLvCXDbLjuv6
5yQD0xCH0NtwBTyq+VNh2TZNOuW3qoy5Y4i+69tkTkdRS9srdQvphXMTPbVR1/RV
lccRW5bGENEIhuL9qo+bOxZZoWqrXYU5yfmED7dGzJb3dXwJCF5Fhbyi7qLx8VtS
mM4CT1RbBuXwb7aPYOvZZOAyX+A29fnjkKAcdP11frLDG1WsfJfr8ZUYWCTytBfY
QclYDaLOTWmU0mAWxy03/9M5s3tLP9prQ00L/AQSPFiD3eTE77aacvp54uU6RqaE
8Ya8dqSNAWWtw0xtD45AZ3eovrb3rqKp7rGR5bD/rQMehaUfa7DXT0b/oWYLIlw6
msQV96py7UcqIGl/SJjW/chXyz6OuIBDEpRGtSL01OwhnkLAHNuyH4ykwbXGC3Y2
Hdk4JBfWlmVuSARgDNekZ4InjjFW/yrqX3xrpQkRI8Bo5ZmSlETIk6s5CczPzZgp
hcrOHrk70tjfHPomo+ZAeP16cDk6Qo86MDyVwJ0FA6bWj2Cxclb6pX0OsXfvd/5e
zcaoeDt65NXted+JULwrGvrByPF9NEWSK75yQUzd5PI2Mod74I9jPf6vsVJ6lMhE
phN2QEf3ZGTON79MLsb+aZIWjmq5yBA0L0w+dm1d6Zh2RvaWHgLVcEHvGMIU0FPg
yGdRzpsVrxF2GmTMrz1c5ErdlqEfS4G1YwGdqKr0UJsjK/zeCLhoA5eeddH7RXo7
Yq04JOLcMvn7uzKGxUIWjminYtYzsgo6CEYyxk/2UYQMYgAyquYw9P51i0qi2Mey
+K7pHA/9dX83ggTKZp11WHjKtV2j8+nxnfXbtVewzqz+z9kXArIKwmyNbwqdmuu/
hvtTnhn4pGenUnKMBFq6FSd+LKz1K7HIKAzQKtSrmQhxQ+APsT98qa+BA7UMqMbr
UWg9+m1aBIHJPEtg9PPS/aPTVeFVPu2lpJgRr757U1NBFyEQcXp2Zm2qLeiGmES2
5DIZB2qxzmQY3Ttsrl0OLkgkIvRuzk4HkRP8Ox9KJIJ4DIcZpgvteNaeMzA2NsnZ
04Tcsg3xB2AvlxQwfU67cSUGRIRRXXyt8/mFXpLZ38YwI5zGV4xycFqvMwCSO69b
hqUaKrTQiSd7sAeZNLCYvO6UKRePx4HDKyH+n3eJq1S5gvceNbSsArdGH593zg1f
8VgvN7NU6HVfh6Ae9Gw30S/2M8f+G+4tNNW01yU5qXIOIjnw5lSPpxkrij3KblVJ
Aeuq9YH1WgVIfo73OLkEc0v/E2JLnSVWm1//72OkqPhvDcyPlqaZXqfLSHL3DX5m
b4FKqlToQ8UNs75siTypEJaAny/j4684kiDUUNDDYBy1oCHV2FNKc2avVZwxgqta
TkOW10l3siSj1aovt+oQIk/x2yv+zCPhJDcIuj8UERXzxgrGdPQAz2FVFGK0SEw7
ZFFX5T5qEynVeFac9wKQQS98/Qg9mH9sLFoq5szENezU6AjZCTXi1z5ao5sL6DKU
oWUmiHiDCaTfPtU4H9rtihD30SuxtoKHjYnpGPp7XAofnVTKVhVkQcwK945+jP0v
yVoimbeekD6i20n3MsmNz0LFT9Nml2tUbloJPcXG2PK4sGpuEopBYHRlI+TxVTQM
B5HUOVsjIKE9FLG7x4IC4MUWMUz+chE9fWicvIMqDOp+fFsnzJFpRF4oig9aU7T+
QlD64oCU2EoOrxEPpNnCffknxEEHjm1afdvWLIInc11wPtRxON6NiK9th7ErfPD7
x+vynh2MMluqmdMj9U/fWWG0LcdMaV29v3xm+Nmd6PHjY2nwpNPJ5Lr61+XJkD8b
A3ljPN4XSRTexl1VxmWbI3NX9hm2DyF7YJucP6O/opJzUIlS7u+tvPgTynccx4yp
f+xKnjGITElvxPhT0Uos+dx/Z1Zc1Ju4t71UO7ig/cLOmQjhii7YBvJQwAGmszZ/
kPzlwv6IO3rIjp1QGl/0G6PpUJMN9HMxOSjGaorga1hKGY/PBbO/ZgJqVvunWXv+
RAtsu6cOg4mnQkGoYShs/g4ei/4mQk05RMh790wE0/4UOwJo9Av+pUxN6e5PJAWb
7Xl3SkTXiE20bt538l2ulSFcelaqES47aY8ZuTLalhRzpDejdwHAaP3gwKkd2N1B
4MyAipu5X+9bnPi5rSssCsDdwy69vLBWPdB0x7T4g0tAVxJ19j4nZi55793wkoRM
jw9+8vaREEvpkWyYdh70R/3sH5fL6VCKz6KnACoQzWb12opoNKCTa31/BUQGtCif
6iUF4jlTTQ7qq+vDaaPAFa7bMPHYhkJhFlowic6Ttj0NsN+SvajNI28AGGbE51/E
v98xsWw9xUx45kv8/xwW0EPAQo+EmzzSGdu7ekLKXAIAc56WICxGe47+vb1FiH1j
Bca86BWM88LRrenDriD6ciCTk5gzlYWtJJBsJjkMqHqr0S0LUlvlzIR4MxzcVClm
C9777e/BKAHHDyAsxaVq53Nu4eVIt0dnx0ZiNZE6pkbfNHpP6U9DuH9DNq5WC7O3
MxWttVvGAS6tqLw+FAbas6aB/8fpZ8kGSYwrV6CZpxBFCgOSICpfP5Zl77YmikNa
p+7puDg5Gj0l8bOuYQd0oMkJWrOulxHqBXulm+MZIrc6I62JNY+oZxteX3kFoDit
+3gcAqHioCLT0H68AnL8QC/CdcwK1h+nlu4QQz/cimzn3yYyMFdqX2cLbPAYv1li
G+inTeJLBU3h4vII0qWTdSQrPXpoVRdxfv6PpRvU7lY56/wYrfRxIwDKRAW6GFIL
sYTvXVdXZaWldiIbEOKlVSu5Y0ohdNs5qVXwteZDODxXTFvY73LSpA4+TMgIEntr
ry+rtEqtrdSaC3wg2P5Tz/FEH3/FE4d3ZpWz8hH5g44ePyfjSgt1+AokrUMVz8CP
xnXYh8YH+RG+0BTRhEhy9KzqB2O2rX0Kyn4HE4TmMEuv0y80FK/BumGaCmFW8m4A
ju1aNjTWCh6RZCd9XZsx2at4ldj8C5TTMUD8khx3NyRi2BM88RqIqBKug43RK21u
vcFFJ8a9B5ScMnxry3uiE0qpXUk3W2b5r7rAVn5dtB4MD2H9Ff957K7C+ACjiQNn
uu0V1/7dMErFqE9DzTHj0BkBUjJd0/PZaiHdCiRJ2AMo6m3JOCJbTd2/GaqyoZn5
5gM/pEpE/gCNg3ao2aIc6BnHGpB1rC1Pmamx0xcZpP3IVaNvJcnUKfiRB7nIp2cg
lBjQUvx0M4Ibtet4+Ic/NMULf8WWBjKYTNqaF+RvBsRAZpgHyIViOVdACn8kgzHK
QjSq1n/02N5luJZeDvQeklwVdhRWOLNstbnueN9ENTyckIuQhfk5O8J8HfAVVumr
sy48vxaQB0lXrEM+NMUbJ7NLv5vnjREk9QCdGfwWcufVzgvBKTn3CL4E2Ldb2xat
JcnvQ3tQm5c5mhKh9YsKWou2f5qZSkvEg2AQFp1OPGGr9KiJcABT65+jhYn34AiH
/X5D2lmJHt8TeiWOu386ivLVKgGowAtHuJ4BtRpE4L1aNoEl4XlrEbrHX9cHAEt7
v7R+EX3mNcsHrBFkeRuZlqJfn1GJLlJsHdkHVf59yMP16TrM7dscsbqRtQewBo3X
LN4/zjzNN6MXWmVGMf5m/Db1wIGILe0uXgZ/evgcPFkmpsM7ym1dFpkBY6XrZ+cX
zj/r0vKuo78J7TkVBRdTGpYu84oFHFQXl/5Q/1D6rQBC07CyAg7mUUbPNXvAI4fT
8yxm9XTpvZMy+UEv75BuEdG+6JwZNfDu8e2sgZu3HQmNa/DWuvxv59GnnDlxNsEi
Nqb7KlbmRy/sDS6CZKPXFulvtElBIgsEo7HIO/krKO7MJuPgFvNA/PrmNtaKh45G
vzq1qVgqAWys7oi569XN0kA/fXJLri5bAvmo8RrZ9Q8jBx9locmQoA8bRQUyE/R7
25OmzSb2Cv0/HlkigzKEqFLNeI3yk1LFjfX7MVpPE4sPaC0/pe+LzCXxKTjL+1Da
o2JmO9GybGDyNi0DgD+3S9hm7373aoBPbNpEWB0j8TNr3GAhb3OdXNflpYf2tDd+
UTTZR2h7bMMCvMsPoGIHi1GYgdfHFB9USFU0fTSzfc7wdkVz6h6TFRiQ8SGkCksS
Uvt+0fzidHGxWpeB8fE/0IynarDmbPXqe10tiov5ftzp5hQpsz2xY3mfMQCgpKXe
47nLwW1i1QsyF9PPfjIkmVzWBAtCOjUOWKw8wIB6ebqvN5KUaAQxy2bOzN5gaVT8
pfRahXeL7zimmFqY7GC16kzp6C4GSe0JWAkPFIHuDxRvG+rovmgTEjsW2nvabgHR
kVLW1+R5N3obFQXGrRQH/S508AZ83tw9cjqz/gFcaNLh7SMFmoeS9nIH66RhwCvV
QkNVPetbAjY9fKf4CTPun1eq7JvJBKW7Io3jOHtSQqoaFW+rU2JjMvzAElZXjHhH
NOvT2JYAkQBehf1vF2/L6qkkeZulhBkrmbki7ssDSNf5dnAoejqv7nbBW1EmYKK+
FOy4m92Oj9KJx3b7NSd8RihxYExKNTVSW1pQhYXoioV6JsKMN/ndPFTRMyKpb/CP
jNLiiX+fU6qOGlciY+d4XESB/iDasdqr2wPfpQ8WioLM95boqBiCo+EjR4XWLW3t
QJwtf6K/3WMxqOtrhFYkFaWX0oYM3eyp1359XCn3jqRweaXJK1t3LA16+FX3Vc/v
owXNww2TwIGok0vM/zzDCmvbJnTGY+AeZCF9uq4SK7CpfnTUFGH5Qq07h+XelJwL
qT3LGCaKUlQB+zP/7IvDWhobM4jGPYjOlfLV69p0wSSE8/llJtqWU/xd3IZDce+O
KTPFuvbveDrzrU6GtT7HtkuqGHzjO0FLVPnJU/06pfgk/5qbPw9vyCqt8E8T+dLt
flgR5itUQt706PaXcf3MENVxRcn60wKdp8nNUmJewlpjjoTmIhhGHIJGDS1auI/Z
Cl9OFYUMYMoQxqC//X7z3y7QMYcgedjdq5lKH/tgWZ/jJx99ZhX09ScW+lopdaJE
t9vaR/RNWfV+k4WNuJcuViiHeP6TtPlWoffP2QbMJssK/VoWYDpr9tPrxf3eqGog
FEDBo/mI4p3vrgL9a6uenF/qZ7keVbIl+eeemL0KlURHlaFWst7g8+2y7lzBZtu2
6+QjtMx7D2z+OnsroFyxuNBDGX+C8sDP3+s3jFdeifTRFiD+f0QtaV2gZ5NRKqNz
psmFOL4uywN5YTs4Eh/YZ0xbT9PJLBEgv/EHky9JcKgyWARdWTpHsC6kBOiNKtwK
s3d4Y1IxoEI5KhdDJP9nzOqs/NZ3MQMj52IynTTNHD41+U2t1pp+h51f7LdUB20U
fUux2KZMLHJ0aZgCw/XwEbtTtWBOAJRPo70VxkOzMOSwbV4ziFKtKqS4Vx0cQPF7
S/WKgfrXYX9jrTSWD1Mlh95PAJalxvQ7lPY6Ob43h+f85Y7Bl2SjBQTSVprtd+6F
GFFs2o+wWoBPVA4DVDdP0NH3EF8LxZImx0wNWk0RF/OXRTdfc4LpS/H6iq7qoEbC
cwhCZdEm47gfQXaJ/3+WejjVId/fKJHWNHZN16XP8W1nyeJ4RDJ36aEtpcWFEonr
ygSiwFzdvUBZrwWlT8KlhHc//6xD4l3vDhNXs4esEiBTXtEyTRDnDprkgXEH/gSE
HBgxYu6PGWaBIBCsvKWOv5zmAZOkVf9OogBfv4r1zQaRFyl7Y7RFPCiVnKUdMO5D
nwsxNv4sImY7i9Nh4mQRpg2BsLo2pF9z7sQ3eszvQVGGTQxs0Q/xiT1e5N6+ut1u
2jNrdb30+nB3867Fqe7bixQHG+IJBfhCVcj73q5O0tdseqKbK80reTc+vvQ+p+XS
9m05wiJMC8ccwnAriQzyLUA8DDadyDw6vl31sTGT1rj7R0iDqhGUc5vmCWksMCzv
h7QsrPbF9+MhX69Qpsa08dEFMTkNZT6R/HcoUT0IHFcvc7XXmLpeIG1MYNgXw8gO
WCzbBgVrwMdiYJ97QZvEEXdGk4ICAHt4i0lsZqei7YWgGae5yXB37+RPZ4h1YUs+
fRhB0geSLOgpfdWBr4rLNx9g3UEaDDIYG6Ehb2Sy21WAFn69psBn8mObO6P5pepb
rprqMuOjmAd4oxsP1Hh4MksfxMYKm8fi4kpGcw308zRmIlYUPh/rvhSTB0xoFMWe
oOSIybxdy3FkbbQuoeT6U6DZNXuELb5tor02sWnxSlwaEy6SnV8iDiJjoCQsSZKP
yHGo1rgbPWpfcZNFKN1kZn3gcaLiOaF/ua91r3yHxVbNEvUnig0GvYCLPyBTfsCU
Xqa0QpjqTB+8dYVLYSpXt0dtPqfNLXbbWpMbbr/ip/DyGi2qelJ513+oI8cUBbHc
Ky0t/3QbkgHpKEzj7j4C8/gCJFKxSXZCBqGYTnvNDUe/6i6II5w99dFWl6WsE6yj
pboT3E2qoyDV0pYPgrfHb/lOFFbctSapbwwemOe7tHUt1YIbQCTIsH1auZtwphaD
rlXVZOuo0sE040yLdIfiltVNGhOFL1bktwf7X1k8WBuJNyR/pNIq/9AsnJ3cAQXw
l6vb5rQLjpdFOmTBBGZbt+c5HoH8FtfsQTlVoNk9Jl5s8aLb7HO1PfOZHjlNdtCH
uF7PL/21m15QMC0dBNzczcn/LRl1+cERaDDQHjlFNN94n23YaIV7IG3QJdPt5dq5
ZBHfaXbFOmIKj5vvh5A/tm56iPn/3zB8SfxqEm6bHXiaJvmTv2KGxBmG6+nalZ2i
pfh99L72YV6tSu4gocilCzfV+SrhBw2uQk1pIf5YD/Vks5f9a+v3vUbu7ntoA9f8
BFN57mG/hoGlzSAl8X721nJpw/ZyvyE+Qt/EAyFe6waTOw/pqgfTwaXhPzYL4QNr
+39NwZJdpAFvhqWQQ0H4dImTPK8H93tFm6OnrikklyKw0KN+5LmeckUX8EfT/N77
yDcVlzj2KTacIpj0wYn6t8YnvHx0D11/CU/EY8RUFizNxMv6CUUdSAY+mhUPAzWE
h1CTz8I0bPXmywVH8fIRYru25aqSlQ5oBl9w3zqmonMli/NI2fAF0mfLwDsHrrBX
BGisPKjphEfiCc0X8VxkGGPLMsuhlnQJ5YtKRIKyhqIS+JtSTSezUibSMZeEhIx7
omqJj6sNFedOkb93a8C0mfVJ1/tx0aAumGqNwxrXpDjmc083JaQBgWJIoF5Qi3+/
7/J1gble00HEliuJVR5FFWnJ3mU2rZjLeJuqEscCLw1k2etuDeQrBrS0wfPIr+t+
LqrIG1Eu292Te3tnQ2uyIYbJYT/NH05dgM/7zGQqm3SOsV4LAsFEAotB0hTpifnp
w74UcbIJWyIQDRlOG8YH0/5rMP/MFOaEVc/aV/9TavJq8pQ0lksVK0vX74JgZbME
VD4/HBft+iGWbFV6Yjus9/H0r6Jnr4YAOlni7ACKLu824nE8hFhJXqeqE/quDwUM
frV1Z29/VaVGrhrL0Zx7ih86sH7F/v/GFX7wABSOW3GQNGfIpOeP6nRzqSIeZJMs
5jKWkG/SEuSWNZFKEzMDM8bLLrCK34ZB4y2S2dkNetYTaFHmHODaFrtHZxoHWRfU
GIcs/baAhcs+8QZRLrINjdP33FjfrFX5zLowlq31AVjh8j73gXpcXq/2QMtPpil3
c5jx9mtsEBFC+LDdSHL/nWQ8DywyPDmtZBd+jCDjG4FKiQURFloq8DsfHhxfFnDZ
3LS1vLbZDq9sCegLkqzK6ZLUfelkplxEiiIS7G+c2AHn6cqIPcywyxdF5wCydXQv
XMH5a+qUtDL9M0d8SSqw0rokl5rVgK56bWu/NSq4WPM2tBUUp8TtvTN/XjTR1uAK
4QLY1iCYVxHADNDZuxFBOnvzb2inBT5EzDduE4UXwr2oTNP322Chqwa5G0gP5mli
n7qQzAY7gYX/6+J1P0EQ7s+ScqWdUh8iNISChO5URlyfTm4G7/4TeBapm/dNZkLv
TDv+fGUGjMY1vqo3o9icSOnLfs4bn8JpanXBX8BGLFBZX2Dwd6vANDHrNblo2MfD
u6/7hq27BtWXw6gWp1gMgiQIGVCj19tCKjPm+mw72pH+uAqGKHYWg3BZNWmRo8X0
CcWQO7slxsSK3ckE+sS6l9MKZWFmYsUJgvwdlcawEbgVcNi5CY1gTADGbxXn5Kok
HAwC6GM4xOI59npXYG4hVBA3TThAdvGDCa8giSPySt/efQlxT420soO1sLlh+xWV
ZaYLVBvz6nwzdUkgqDRSic1jJobKQO39ZFw6IOT/Od63b9fCVKbMVfjWTcMSqdlW
aWiA0NV+juAVmtdPUl/xqjTMO64N50GqGW9ur73ZAQ1YJB+INkOlbpfXFm9Ky2bV
7pcBql5hMebw8k/Vpp7MmA3DbeVRIsa7VqOW9PCipWErv3jCJHZg7dJQR+ygO1zP
6MxiFoarViYjH5H9h42xOEvIkgXl3HTXLWE9Z+sO2ikyAig+BquU+qf6hg6sY9OI
UxtE+gulSCxmZqVsaQlpsM9MG9AfG773OmRXg5tWOhVTlIjiTQ74mC7S0KKFu6/I
35aPTiCnaQB0eJWBAmRL2Q3nN2YyRRs396gPS+A6mgSoYfXVp5ZX7zr2kGfTRNHC
+Klmp6Lx2uhT1/u6tHrbgKqIO9wNushVQTbocNq9ACRsxQSEzhsq6sOq5+hAdjXP
OybE1ep6Khj1qGkv7pyEGoZ+IUqI9MwJMyBpvgrMqx9m2Zh0U6vMWqq9DX8XaqTg
ZD/ZP+IuzQEdmkKpcyEVAZKpPkPDylBiT3sI4eFW8ES3bdUgEVP3bydjiSz93bIr
4VLS2uN3Ga1s/+LgUe3qvCTCWiewvOYikGPTxEs8xl4DdbbkCag0a/D/JBruGYl2
GyzRZqxracBQbq0j+2jAl9E7x8F5F5V9GkuwSKtEwe/mZUPhANFnhIx/RZIuGWSa
rIpAru7M0LAU+tq8gAwTDAKb6sKrZAg3PVl56TKxDeT77tvWhZ6oi3D0EoH6gpoT
pFJrhi/B7SG4hpejDy/M5gXp+LVWEBvvJ8xcQkHbaN104T8+XQbwiQnSHo+9a2+N
Nk0tkbjzBmWMthS9cYlHxSkPT0u7EVfjwYr2diZZNqBgMvgTadG+r3aWc/Dv/V/O
0dduzQBTrI33x2Bq4zuw8TQij8LtBJHsTLlVuTqjHzupCAxSrHZvzxFciMeNdn/Q
UQZM0wYThpWjKyugMgM2VW7euZrjE+xXMJoQV8zdqUzX1f1hGCwDbbLKjSY+IaMs
1CpJyhvrB4TNsM7PNLyilWm5cUNIR5HwMGQjMqlBjvpWZv+zq8C/UKe3laQTmrv0
d/B+rG/ihX5k0er1I36JnNEdLz8uM1ZSxYFSzzX5QsJaV1TWJm88Ml5mPeYcgIM3
Cvj116qYVobOPfOfHFJ8TUggqnmKdM9dps+CngEjtwUtg4dUyqk4elxBnyiO+yN1
F8BmT5YHOeNt129uZp+xydUTyCW2QB0nvonPs6j25prmIAD8W2/TZtqoI+Cw+EcL
cHlKqIEbQLb1JnEMgqffv7tK2dS+3ha3QqUAGBx2XBxDVLDMb+HHk9lkR0rwLCoi
/NFQZvQoIXqoboIFnQ77GQ8txyZ6rMmPBh17gCeojpHS3tuyZeBuOdl13qV8lTxp
UCBI58lcxzXWoIe9E7BvJjojHNdfJ3G6maC6dNNK2Fula1ki+l8TjyNNiXo9PI9T
/I0ph4rRC9kHZlm0tb9jCRiLaMUqpq6gGg0BQcwMBP/TfjPBUDfa3Oqg0vsNg5qK
RMUp4KVLT/1vjlbA+6ctDhZHrgBea+NMjtBUeXV3nOotEzm4nLbQHzpjAKFjeDXA
oROe+dcSFP++h1dACH8yK7bvbREOfICrzXt1w5mEqjKvk9NnLIE8s8Yt3ZwEiYR/
DG1QW2RICdelXnV7txpCGDm7wNOfJuLM6YafOA40G73F7H6WDOUrU43vmOYYiB/H
6PZ7TeuAmJit4Fqmm+VbHPc2aBrZlzNEh3G4YrBgF446VHXIdwhaXdjzL0PjoZkM
eFLa14vHgbD7EVZTKP7+ewxaBY4NAzKlOacuD05XS8W24evAqQeMHBU6Gsqx58MF
NtTrVmbZAhhpRYnTf8gIlwJJJupdwSaZ+/1qFgd9mm4wTA3/thLhCkxaSXnpZBwb
yhGWmJO+YYYrM3/LUIj2o9eb+MQ+t26vDcvi8uCFGMNxg6P53hp2GBq0ft/j0aJM
nzsaEV94mGEvoB0iRyFmsedi+GOdPzmElNqQS7TJLEAULAWcUDVPnZoNDesPG4HQ
M3UepyghIFRqrhdWCoqISVyMWwzoC24GXq9n04G4sZoWykqkFOxqhMowplDrPHPF
lrH3PqQ5cFh/JV0Bp6fetWO/kZM92Vre+3VnG1OrGS2x0r5r5w5xnTWBltRQSnX6
JSszzOIv3ZOSu1JERofK/M84PJb7usMknBIFD53+CcjqgVBPZpktLMfFY/P1Hxwt
nMz0/GSf42nNjjGujXeXuCjf8Uvp5dWrwT6KL1IBehDpd/p7U/Tw4jTg9WKJdo50
6D3R3Z9vo4OsdlLwmVpLJNW9KpQNjcer1TduGSGTpn0nSSWP4SU+knVX8hxhg915
09lot1/OA3hG8tQA/tfmBWz14YaCnHRWOXm5JR/CYYJVG8WXHt8E7OmNaH/q3Ymq
EHWsrBt2AAl2JhVK6fPYdLOivsKQCkUbSSipI59TgBdrrMXSUGXNMrM/FK30ddPb
1mFjowzzXYb5tEQb4cQuPmcrglYOpm55QqsZ5qK/1GsDUwPF6fryXRFVFoTX9ZM7
g8pG110G1sQyrgAQhAaRlygdUyXPYwpOybUgpproRsIOe+aZVGchIYlrNfrN18G2
002h3OpeqxddGl4qd4SWxWEl+Q0vBl82SoyF/XeoK4isUhcSMZ8jsnP96MW+zSxx
tbPpS4XVrfhR/uW4myrjCYlIunl6FDRIJGKwEGDg1UK3JBuBAhgFPO4EWHrG+Yi9
A/iVZqEfpUAe4dGOWobiZbv63/amhoKq1CjLuwm695bJBaWlgKQ3h2tJTc0nth9R
glOsZnU7IWBBaCyl+i+6HqPTEThE4wZ5DYTw+HdyBCTEGGMlxU2wzB9lDSUdRFqC
/cGNHtjdFU7qmFQzKcB4qdynX3t/EwblBRLnqJH494smE4+6mSTtyxB4GKzLcMEh
B/f75K+il47M/AysSVqtFAvNSKTiSA7SHodyzZrsZKLvm/1qQKt8VaFtgl2PEwky
49NbMzdjW3DzzCn1pPc4WoeOdZUb0HKWlv1fsojB5AXMQ4PadqzdXJfVUDqbb2xA
p5ghbbeRvqJp6mpEGjgH3pOvvPU921bFcts89RwT0fcP+V7GNyVou+TMTMLAa4+B
JZPjvcTOYQKRfsTkXmbP7cMX2S295IJoMoLXWkDkwgd7JKv+pZ914NbC2gfIi3NF
SyuGC3X+JEZvH8K1ZXpEUvag9k3bB7Dl0rg1nx4ZiZDHX6t6BdOTr6NhzQyrkrRJ
aJt7hsAFNC5MLiWF7BkwxxWNhSNERgqknKl3gGU6p0SX2eLdG/IVehz4RmM6j5Uy
iezcLrAFy+3LmU16IvQtzYmRQmFODrspB6skORQNpDGhOUR8peF15dAQJQZnLPWg
Kd76rKYYYPPg5p6Txl7xP4mry0VGfjh/yMmTJ9A7RLeDi4350aNaRHvnNA0yj6q/
Glvk7o8Txi2IysPNwMrJIyJK+1Ou7cwp7gbUEqlD4tXMlYaFX2ed+/jfjLQpXWRS
wpR4HTlOLhwzKTho5u6OVFj2TNXo3z2pcPH/axq9AqhKZ8I62zzzs0XdN4aCjPLS
miVzEuSerYCvNVdWl8M+bLQNOfCXzmPPQEJzoOOUZlufAamZf6u6//5KN8ia2EbZ
GrphQTvBx90JEDIwkhJaG/gvGZmrUwQ2UvNTEtS4G1578B8ZaBOg9B+SdqUpCxS8
8a7SWxwKQGAE1WabC8vfgwOiINJdhFmBRn8I147MVascJcyXAi6z000sDaYbwmWN
DHf/HUykCkxF1xnsi82S6kVxFGG5SNT5KXzbL4m1Sr6YIqd/dvDqoxkxK6UvSw28
tazlIZnd5dpkg6tc2EPEzZg7PFwurGUEg1j4lt5/uj6/PPuxaWmfE8i7vLUnvS/C
Kf+awh3OB0uAkUwVLbedEuhC0PfKOhlJJlXu/S6TSuz7T+3citK3iKr+YOIAQN/+
uWFjlFPf9GX/q6sGf3IOF58spZz4gGE+ZXkmEYS4wWsHl0P/K51Vj4Sa6F6k6IOi
Y6SEZ31jAH49TPTh9wq9Cbvu3gL8xvLtulVvIt7CRlPBc9TtSjlsuWHIb14wPlbx
yBQaTiB0oF1lBbfqLeElQFcMCZYikVexAT8RAhhGVd1Fls5s5h008V6qVhv9Dnm+
JRZJ1s/SMJAbdICmW4AtOJia8GVKap392b4d1nXTomrrHUD0E6OKyNYdV0lo4nO1
zckfvrWwG1qb3UedxUiYnfP5k5xn93A5F3fiDreu/ZXa32EWBxpKhfOLpImRFdfO
nIA0iLR1RAZd9nbwYBkgPRUvlCDN061/YYbFwWeMRlVustJBc5J2ANTqKSs9iZen
6TntCDiF9Qe50D+NE+e6YHZpqoq2msvCq1oEhtr/j6ZYJbsptfH2D57F3SpqP6+U
4fe1s+RdYYdioOutImwvrWDHkQ2Aw2s0GVAug4hzVWHjI2dj0acKZ1oc4D5m8cm4
JSZtEL0xdtR76QNoZy/T1mPXNiEiqTvoVaerCnaTYcJsTBJ5xP7F9AHrtYKQSFH1
oRc6+LNuPLSScOzkcRFn00gzT6FjaRaEUkFhTyL2RBDpKF4q7BCSUYKVp9FwR6ri
4ChNbNAIM4fbhO798Lwp+AQF//npwH/efn3soPr//qPvcbqcVrCYCTIoZH791lFb
HybHz6gC7hBd+o1AK2XPoVQsDag9P3IqJ9VJXw1+UZ1A1rtZ/Z41V1h4Bz1nl0hB
Gkog0lym5b8a/sDE1X6rQNwZust3bSegTnOjEkxqt8eG+p2adURH2J0Hdgk1c9NR
YMs2jYmnhqkqlscnhE3uR9NxVp0kCz0HXE3p2mm1+FpdKGmOKBbffJ03qOK+cB9M
uIF7ilprppfiGmsjZcCsWAFnhCpwsJuX7YORb9RmPSE9R1/23DGgw5UBmfBYL0L8
Vh/ElZ3dewaGWSHScUO6MQWB+Q/1UbWct4hczJehm0PcbPpVevwxAbg54r0Q2Qah
UE/ZZ+w/U7hsTXUXgcF6EhcwzFj79e/zn6Bl1Ehe96WdOMac6ZQrE1aTHhan8RxX
rogxpbkySly4OkfHjwEYbqtRDtDs7HXeTKC+ZtEVMGWyJCAoSSthkeBkGogJMAfE
cQ7NMDbFbCq+GxpFgR68j0xQeVE8RpCjQ0GACwSq034MTVAasLIDCET61/P1hquf
1Ul2WCA0JFkGaOd8sxLqUIhR2mHqA4LVhp7evVhZOLaVnm+npWUvBLXAtt/wSOzF
8D9XcBeFw6ZIeQqhtxcmxpKqmJIWJkP9+NwHs7dCIn0aINf1jA8lKfu+M2Rjkt3t
RZ06P7VgQrVOn9AQFruae4yOv5Cv8GufqjvXqpdeD29KEf+A/F3tMYaNzsgYlist
4pZXU2k14aicAOzflwwDXIVOZwf2HnHApb7zgIJl0g9Ojqtd5Hv16tX+Fm9cH1SC
qA6C0lMAX2wJT8vrv9Gd2NqpW7qNbafC6R82lIC739o0VhlkpHBj5Xjyw0qObBwp
Uz9Y5usQUHc4jRBmxEEoJnKcIoLDI3Np3wUAeTOHq5Ei3cyUHC0cDQ1OFe6YCK6g
P9aRJaxndMuCA7z7oo88Yais/lSJMeiwoWg/ipwHdIR4Ad5/LkTmZD+kutZGBMNN
i3pQSWA1VBsUL7ItCxxt+sy2UntyonMnbAlmdN77GEz4Brk2mYZHwVdNJfrXsRWf
+0nXXFX6325dRGT7QqodpT8io07PxeLUL9RiICxjpKa7vI4U1ngepA0oBhWYNxca
B17iV6/+hAtsCTUONjdKCvV5wM5pqc3FB/GFwxxIXPBAGph3J2dxsIyB1JBVknpF
Xevqhfs1eir7fPkU3u/SjSzRg8EVKvgTqT7gGPQPWHeou+0QRXSixUCQ2GmkoWmD
r7LYj9821bzIn2xrNoCea5L1LPK2mc4rk3ihutpYTK0/FdSlsBod7MjcwAJdFEzO
SKvSzWQMOI66XM8S0YuSuvQZYpQByGQm+6hudo2y8asfT/HcOcFfomSTk+5CXDkA
G32wKAKxJCNZMkXf3ZFuE14VDGQQVFeVmC+i7Fz9d5UJ1AeqzeXDr8wKnNQwBQ08
+WvJipTJ15cFQI0LpO8994U5bneMQ4svtfu6BRQX6Bn2Br2DY/JDWFyL2XELZ2ze
CReykSp93mvbYYl65F0hVWQNqkv0TXUPZDuyb21gaiWboA+vsfcbfcS9UnvX2jWc
hd9NNlNJg0SwtDojubq824aGGeHqOqV1MUF0y3zOUdvgRB6URUdIhsboLk9x87Lu
cvW3ge4IqnDVN4iRrFsdpyTCm7KkVkpHJ/CRqB5JTQh/eEoSNZhN+9PqL9ogBsjf
T2lLFumcUT6ciOGtMnry+aI+btxHS9pxhOmiBcLo+jdzyfkmdRT0em1i8wNuDX2e
TQWx5UFj2Te4hd9ygv//AjQVLVOwlkJt7Snv/Mx6S4icLZrZXBKiWG318Vw/sIoY
y/lwS3bwohA/yAXq4EsN1DH4njgRlDztCzrqD9QSDA4nTTaFPPgLraeqn3SLCzzB
tOpmZNHQbm5UbfxMRAuh8/60GOFFJq6EHgNxdqiS3fNRBQr/WN4yPL3NfDqeSWG/
cskYnyspcrOUJHjVbJsBJ3t2lYeVsdBjI6aECMYxDnZofLZeFmqUy/2EY1pAaVn8
oyIhMjQCw7jKKXNCQEtDX29zOEOKmM8IdftoSow/YJG1Ra0GtrCFCjNjPK2r6XeJ
S2pNkZVbpN6eZxrfKxCieLo6iUj2UrT/lJpDS2r5deaWRQGoHinhLF35TofV8jQC
dUw07etmhw+cheLHxsq6wnTEr6sUnnFN4QdXKhFIh+PN5sR+KzKoxSMPBCafnng3
ppmkt1kMIfGisGkbFxYNF5tZDzTO5BFT9I1eBiPiTZco8gksVEo9Fd4udSqIndVL
6xoLsER6XauBRYmyXm9lNeRucmqMTXtb0gDVDtIf2oq1EyUDnpYM+FEWty65qusK
UiWn+wuWx806ChCkrYV0VxbwmNmICaNsRGy3naerYpu1AD4198nnRl/y5IiNC85o
Ge0r4eeCSZo3VMT30fnpYKEfX1kKNt21kJPEymR7okPcO062V1WLK0pi706Gjc22
pMqT9HRyREd5fNoXzq7HVa1hD+U6ap9gbqmMppEL/Rb3XsNMiSGoUVHBo5uqeL8B
N5vZolqhV5+LrsZCYuNZlgQBhL12elI/qoGO8brk23EQrHqLrZN+hmm3g9LQ7FPA
doatjwAw+AhisV3DOKTNYvo32SGqG2lO35KqY58qQg0AOxdaaIf7GbtbmuSIkmYF
gU5DoLOdon1P5G8pTNx/g2FHy626xSJUSJ9p/7hnfK3KJCuwtgc3UQgqO3n0V7EE
5XeHbgIlL8d7PZyNhXWdHC/CI2uLRmnI/Zbl7J6yiVPCQt79GSbYqEOSpoIYcTs2
sHgigv/hqeaYbDIO6dwoO2/oOK1DpWeg0F6uCxY22M2o/HajViMfsX01/Wmc817Z
qsOUUOqUNdx07SG5s6sQvTMwvDl7kcTy0WlAXqZ5+wAj1cf2KoPYPZ2d3nSMcoJP
0b0sTlp+Q4qVy+RKYeeIPGf24E1uy9QIf6TyHOFRE5kkFdVKAUFipV3ons79MIIB
NYBk2o+fdJvoBaYQS2i+YMJrH8CQbJ/D2vuNBUmW4RxqPnkV5Ec7sIiFQHHAgpYe
Kyfi6SthTbx+u5u6ieJCnGaFxdIVBymOzIpxr0OfRuCG9/3K/yPllyFmvVrz18Gz
0ea55zejPlFhu3HhXikT/WFwkPwx0SUao228Je6h/CiwXGIYJ1luRYjPqBf8UEbR
SBU/6wNjCiJ+gLOqsRNeI2ekn4OjeA9aHzR5xfk+Z1c2AUvWyTCu7sFevC2uhqPt
kC4HznxzEwIpPPgIiFRCBgRAcYsGbvBww41wBb3Rqs/RHo88OBiUMzmw4CEgAsUP
/rMe7VQgevZOtHUlCgnaqSd174YWJFp1w8F24c+rKg8GxHMT7RxpG5/F2cc6UV7B
i8dJi4IQuASSyRfbXm+GcF69jrEFtmRP8iIntdEptTS+QZQhJhgaRuQXpyYGGAsP
F+PRHN+zRfhgjw+EuwIbAfURkeTSYKD0wkxymsMP9PsY0O9NTUW8GTX1I+9eO3x0
4qzk9+MTuuPAT4O20Mpl9ABPmJsvnSrv6OXgeQmranZ0kH3KJ2uRE9aFHiWXTX0c
O3TTRa6fe8knOq5DePC+ErBezTWroICKNNvNXXEshMnxFLTua5eLGy+sBEFd7ca2
Sv3gUPFLt/hwoHIdsiH7pbt85mzcJIf9I4TLcNXEm0QRyodt4+HoFWzVFfSpbrm0
qSIzTRrBTMyhZGa9NmQ2YLUv5f/QoqTLn/hljyWWyZVRV6rcx1l+cEcuwelpDSht
XdPXcKs4bCDlkY2t5+R9vUwb4XLf36aFQoLs88aGFDiH0hPaOi9xH7WvTbIWrAiV
4wMG04R41lIKsDUBo3APeU6+jllCJMVyvsJ5cQzX8q28kt+8Ua0aYTGXG4G5PJ9g
ybhmbc6ydy8dB5n6WKmcR7NHzJE/T6WHE2mTaV66Lh20ulW2k5JKBshF6jTe6bmg
04qqXUclUhR5J8lhzK8XyeOTBE2UIWVit9YxNpp4ydaJyji2SaKueF5NSrDl91R6
vR1PNR3cobT0X/1kKDcTJFngrgmnqjauLBSl/oeMrd1yUSC6T2E7f6BYFWNGahtQ
OmvKZJs813QP1OH6ooJ+Iw6Qdo4/Kji2Cqe+GNm4kcOeLZ3Y/omIKjnKWI6efFQP
u6HxfnxMng78jBWx48QoUxr3gblsS90aE2tKA2InSv/2l1kOmWr5dxFrldXzGLla
ESTHrvq3SwlcCviAt6yLkLvohsao+gqx6MsiNGtxeUVjdSEv6K5kny+2w/kpkyn9
x5+xVt4Nrx1DQAMHMHDc9pVtzlbxueOyTjYC3XW9KnnqHHI9G9tjQSH+k9/k5b1m
keCLytfDU6Bvzz4Vl4wuEeDWHuNynXcI7hhL7omuclMNDkY/Sc/IbRmthfKMIjml
S24tpowlUUAxAycR5eTTJ+Jx9AXLALckkVMVmTWTMHf9q+Qc2q19rsIKblPkYOcG
2ElgWGV2NcOycAQ3ldTZR1NgToQTEIw82aKbQyyBT3p5KiKpgB0TRcnNpapPUQSs
yFGOSR9krv+N5l3Jlt49Xf3RpNYjolAXZ2bTwaPWZBlO5pw6LU5KhQXGPraIMHBb
8pnFE4vQLNUGKq9GF0zFXNNh/pbA9eR5nJI9YEQ3PeUyzqVjYlOzmvnqM7mq5dvV
55rJc8Dn5q//nH4kZ8jczSsDWXqp+dn10X0pRtCz4Aha0odS8rBo4EOPBEMXfkGs
S9Z5LwyN9rEso33yc0tMsO5ZY+7O0e+bByoXlk12oQNZCf3sAb50Pk4wh+He5nmY
t7su5mJz9Z7jBWfLwnUq2GDepOI4V/BBk6RdeAVJjsgLdsSRdpCvSaHG+EktW7Bp
3UeJyNQUnrGuxMcKdBTZkxZN/zIeWrQ+//CXlVA0rtTbihY3dpXVQiPZXUX8+Hut
pCzn82szR4/avihXEITtNGppiEnlGh3keVtJ9F2YYEaVuPfTpaopclQ3D/vO6ktV
Ua3NqbW6dOnI+tOZsdm5JrM+tHwDMh+plQvX/H1KOyeyQII6OoABpChN3kQpfqP8
IElA5eim3lNcLiky4BCuPvQGysHDZk5BTcEYUqClj3Ywom77HMEFOLuhil/yK1xf
qenUyeKqOfXcbcvS/IbBYM83dgfcNqA8re1A3t4nxF/zDzDb7lzjfaOzevCguGrl
CW6SgFZ74FhUm2iu5mxEhOcuo+Nh8SwZEPoLsLkzIUJa3WCrdG910XCghwlOHETE
urC+GnlVYwinCPtsvmlM+CbRae+Kka2KCjaGeVdCiO+9rA5u90Hj1PsWEBoJFcbK
1S93wELp4947wcAwesxrrwFj9/vCR0EeQR5n64A3mVlnTXJ+ICryyN7QSF4McOLA
FAy3CmGNKY8QvlKtRjrE1zshXmPGBnyj8mkaCBp090lyHgVdMAxzV7cikY8v4u/B
Deu7c2G/UoV4C0o5UJpg5yr8xJnG6WLWi2R5XQ7qAVeY+oY+T/Ht7o40vT3O1DtW
yoOToqLUREi6Ey3ZrjQbYBYvayyrJTcPJvyS3IgziXAztz9QV3M3uy0SWXtm8uLk
/0zb4tK5/5/tpp7W2TFZvhO7fS1Zo7wkWka6izHSBixEfTFcXxZ5JUb7PG0Qq7o/
iZuhgfzM+MZlPzEVmHeXFHh1UMo80H3yR6eEqofBKG5ZMN5bEie+bvb4mpAJ0e3w
CrdyJblcXJbMj7kt+xmwvLAani47g4W8smYYxr86Fml37VmDVqDpt4rQXgXaEVH9
5QjyFp5UaMrexAQk6VoGeQezYkHJJjewffAyggIlQwy3xVFacPfl8ZoBjGVdIxTR
XUEmPgzKuvaQRsGrIIXU9wnXXyQMurcFQJp7i4whHZooNQhTeoz00fKwDgf/9iZe
uwB2VGo8KEJ3cTrRRGin+ih2japOtuk5MEmpaWPzyQc6LcHQ43smJLEcT872Gyi/
BbImXOdIqZDstbjOtthhrSkuhmIE5e0o0kGtsz9z+KdfBNGp32Fy3YVSCCMb4OJP
9G9c1cm/lY7g6cnMMJzBdj9YdT/JZdLNk1gs/Y6Iaw2uVZpXtHw6jY3aX6zcDk53
CypHSknGbZugckefXiZgWuKydg802rDeaZ5xHmQ9Ipa08Ri8Fas8DY8Pa+Rmv/b1
kxuzMMQPKMtIPv1HXclRDNpTOBi9H79RE/kb3PqYFCCysf8yR5A9Gcs136YWzp/z
RsXx5/Ssyyv2NU7iYw1wes3bdydEDwdyhmcEYsuRei5OO+IMTkVqH0r/Qr/QmspV
wu12jbD3Tm3zxNLX+gwW+bKRe1nX1pwM0cm8vjM+vbUz1bY2PnlxaHi2bKuiyPis
FS0ZDHd8mDS5o411yxGs2VdbdlqC/h1K5E04H4vDmWgfWSCOa9nvWChAb1Dqbehn
erNk9jWEZLN9y0bjh8LFJPAKvC0fnKKNNBycW+6tg3t2tiAoV3CC06x/DC0C6+l8
e0cTSb9VN1ZzkExm4fkDF703k4pYokJLgHYVlBSqfCRUVknrEp5naUEyvpS+a1Rz
ZVk9rGr4SETzYLrtdRyeeWr0Db+cX7Tt/E1wRY0TwKnJqN7ro7XjWfFbA+FRgHwO
EvA5V1y/0QUO0fVka1EYr7DoupTsoSyfhKBYaLv0p6UzZZ26O9/tgt7+mLG6Jrh/
ajGXKng5rH9fLITBEks+hnM8d0r8iAKiKoekJz1QMguoaRlcTscWEaSKLuHD0WC5
XcfZQKa+suQP2+Ega4t7AMsb1355SvvA7qX9+2ZqVldDDdFOnmvjteR+RpnqUjDQ
7HYLpeXoIj59WKwr6WbQfOexHuS1mqruA/72CwixSuFnrjlomVkxE9ElCFnGbxpP
Ephg6bky0jzX9ZfmQmW+wuwGKHyXNy0MactyzvImQohSiK9lQcdLB6VTUuu3Qr4s
XG0c9kBcSdk2cnPG1Tb3BLl77v1l13bSRC17UzZjHgV7RVf8OMz37S0pVxFiYiSV
1s9fRt2pTmHe4KY5//f7ko85DfUuVNw1RfNkFSit2r+FeghlhDswxbJuWMYb1HDZ
HayKExAlM16oHb9eqyRJDZBayTOruKex1LKj6dotdmM4qEJfSVbSmHmDQabYm6C3
+zoJIfiU4gWg/5n+TPb8nujC38wowipz5dL7LVxJOUS95CSoO/+zTwznRfMd3Imj
1V6hMtcA4LCzrWl87jFqDOeJi5DRFyMAHJiMTOI3/5r29Hn+qoIKw13xSkgNLUUi
vQB2urpETQYXUlgvNguSZ9aOW7e9MImrZ5IAXcBCzPagKjPXZQ1zn3mSsJqLQMIy
rrMFYEMUVIV5I5WdBs+x+Iv/7whK5oMyS2Khzje8gkXiW2wn4sr14Xn1lI8CfkPj
3DYsx/5HbCuk7oSMRNCvKrIOZrJlNDQxiDnd6qntshMfNUrHIUTjY36vn4Pa9POd
CY8vOgroUMaopvMOqmwl+87KpHTwANvZvOy5zOLWDj/+OmuHCvWWojjmbffxgqQ+
G8aUkOfmNHqZnkpJxlxksBM0SZM9TmwBky88B3EAeILoUadvDeSzbDi4SSeLZIhA
cFX84IEyzqQ/8OB31JCIJII40eWxaIodfd76vomrC2b+cSK7CXS1JMs4gf8WUpw1
U/JZQYvsXoZZjn9AfXlI+cw2XLEabqUV2xuDmKp/4dR1xejriUHhVFkys8HIHu26
NlmOwC3tWxO4b2hX1h09/An2G0M80w1EzydpdL+8LSCuhkEsYiQ4X2OMtft2A2HC
eB0VJdTO9pUL5piC+wPBULFUJ3ylrH3fxqwSw3CI6R8znpxYphgMkKypYwiDGvej
l9gCt2S2EohGslpDZBYdg6E07GnjwtWsBG37xU02p9uQiv8rgE3mWS34Fg2zLj3W
pL/okciPMAKLJVbX2oIhw0NppiB+j6X0DtL9OiHJCFEYStMQ3zGQdiOrDalHGE4j
C6Xp0u7vciotFmD/JfM/uhnQhZmlood20XnoX8KBUZb3iLpGmfc+Srq5F+4h7wY1
PVhWaN0lmj+lBV5w6bMeI/r0o7/2OMb7PXu71PU3+d1xlEwmNROlVaI4JUJGNItB
qRouLAOsHTj3ru2ctrTKNcRT2rx43tFKGUdC/krbsiQgneem+qcu69UkvN8HY48r
W1fwx+yRAl821m0cRqOjA3nNBlY1XihoJYDH8e6pd8BaeqZP2pTNuDid8Bkthlgz
nG7e0W+hVlkIiHbfGFE5o5PevdQCfd3BOplAUYEj0wYfxa5FjFWfDbJxB0KmuBkL
p4TUA1Rs0kzMv7fWYae/xlGeLI95NbX9B3rVyNIXzsDTmMSxKuj6gsZatAypaq9F
wIFOROaCPliTFzl4O7oHLiqYpKgAnuqRJUIy0ClNkPLKpO4K6oqJEJNDXSOL5w+v
CEHAREw4dvVEIGjofPsdu0l9AHLWggRPGYBwqmIaw0KLc8N7xqeboGwUzWKcKPX+
3KqjJB7JP7VpS2tAJ4tGugIH1h1Ne7NdzG0pucMYimBcza4QX1fHG/vg7qgY9P6m
tcUKF0M5YCTufjI//icZK1gBIslZ0yBSKnbASp5PmvHWJcxf5hfe8PgbBlNGxqkd
OZQnb0VSFt5IABUJFcAo0wBs00LCPQFRb33Sgj2SPwnRgcSJ08JAS0kFgKSArnck
ccGtLHRuKuSWszD5IL/YhPbMzM3jLgV4vR02JSPjLOPtbZPj2+z4fEBgyboKSjNe
Aq2ItnTqtcJG+8C2YUn3QcjI6I9QuND4UQ11/L1Vkl9nrTqCkrBBE5Zxu+Kqdz7x
be30vb5hagPa55nV1GwqCrhKmJQe6den8q1UFo+2xs9g2dvOug5MLzUGOJXdH7pQ
f89yBitzjzZBI4LL9GnI5KsJ9RFAL3vS3Y3Po67XmSsjsMlaJ3/ujPZY8jxMM8+W
2cAFtpC75j4okESfOTYTrsgoXTSBVj0M0n5afEwEYTJCV0Rieu0eZhAMXv+abaiK
h2uHsmcng3icYVKQeNZOtLkpfuSLrix5HpcKDfl8y10+P6dHiGyVnx/6cOXJsT9y
xum9xTjD3GUFr0a+6u1SeDVSLqVLQStF8JnYmZtvmQ8NWXW5sMT5GhHUatLL9N0l
+lTJN04nz/aDY+NX0OYUpktkIRcYWcjxAwEP4kxY2c/nGrRd3PvedoLF1p+OwDXk
+rmfVloFLmxtGgYF/S938NKsMGD2KY1N4V1lalYlRn4TXMvnHh+pT9LB5+73/XUV
vz1NG/6xNEql9vU/LeMa+DxFrLNpGFHNlSFyb04weNvFIeu3Qz1hXDIXWuJeWyuU
i18RyOwrVrdLvDZ0hSlhDOgHwubxtjUgD4vioUupWv87tU5SB5KCqIcfX3nBmIzs
Fqx5wTmCnGD82t0mgkS1baLQpQ5TEQSE+pdpcF/cYqIoVpR+5o3QK26ONdHaZRE8
8zO0Gp8bmV7SrnM6DgGq4ZGeoPWOGT0c9iZR9+RSV8Iu7kr075WXExEkWpLwC/N7
GUY56Acn1m8IFKb37bH3puLTYXUhmKt1e4cRgOyt+ZmiwLSv/GhIbfqNBlU/4vDx
nmq+DiH20WzARAvVOWs+kSdV6oC3IuCkfID+toAb+prWMLuovldd421A0A1AbsQ2
sCMfeyKhO4mv2BN8hiY8GmY4NANAqMfTwJh2c4yTgoZUSPbsHl6zswW+io3h9gHH
BZcBqHmMBolHdAng+Ju1m9edCYrduS1KYwlicsjV9XWL3K1rr4RAio2gLYQN1p6A
1Bo26FDFXcsU5kxECf7Sy59YLe7Ok4YEndOhy3VBLWZAMlVchQ1kA+y1X9jdWtvO
yex0fIAXu2fIKkB1TWTXq6q1bw+7zqzdDQWOwnHDqylY1PuC2kFxTOB3TuDNx6dm
iqW+mwRCCRylZVnZOI0FnOIu0mRqybhBUmK5tCjyQ+fe7JbESUUGQ4qtxYntJk/X
LOsCkdpEok/gpJg2uHUY1jXwDv4YsYOVshqbT0hOuklXtPaN8Rhmj/z3C9clgnL1
ozxtMJ6ZZWaqOwr/Ah0FMEkEOGYIPU7xMSOeWDe1fuxS0+er2V/WaeRfnE7nEmvC
IW1u9GagypKhBgS+Qre+ogc0OOmKiNmisRED+JR/mJgpOWlpdHPgqLnRn7WAhhoI
iCQEERA2J84iMfmUszzdsmZnkVO1YKcMgOqDoLJGrK46hEMF3JrFZ+aZCTacFRkP
12adxAdpbSfjW1BxePmNYLyQXYOg3OLaqngeD/j98gs8cLiPcnIiZH4LNcGIx+J1
4KYMMJmRkW1cdi1NZ1YgYXhGuWhh/bZCaPgmJrRvdenGdxDcIe9x9zYdrO49N6ij
0w+zZrrhQeNoIon33jFqlnhdEMWdJ1lZN+w1ECNU4pc2pHdYs4jKzQzy71cdX7T1
ze/X/0nvSxfBZqzIWQQWtRzW1a0wjS/uKEQj/m5eINjsq9p34Frw/adZ5X9PlZ3K
aUIMhSEAceXnEjWhAh9jyMgizkrQS1dmVVSf3X6KDg2AQSQu2n7n02HMsqzxEwNZ
9XfYd53jh6yKbUVYEr6vpMpCqSO65tJGNLXMx+he1qlZ458rlJNOycmvn8oHdkz1
cH3eu29K9pl30z3H751BfRNUzcKdc73F7KK6dLn7Cgin4QaBS9qkRkQ3XJDf776t
DFC6E2yub91jtiA2CdHIcZmL97sF+oyTR4c1YScl0T6Qyxl0pfOKXBWY0tZv7kWe
NoeYjE9I3p3DRYt7BRTzuzFjVu5qVEj1DCr3jUnzTATz6qsxk8yYZK5FfLAMxKc2
o1axPrXUGtoy+WZ05TzU0AlMvF9p/L3LUGxDXeYAeHYvsQ4Fz6cno1JeOfhaqkZH
9g2GQ3NIdcAFkUoVr6S7ks5I7pVqJV35fLjaS7JGdnSMPgN2gSVFO878TZI3qdyJ
r/TP6khdacRy2jGm5lMPsc1x7Zbl0PpqwKO0xV8DswRvHfRgafjZR2j7uV5gcWwl
uYmR1nq1Hxxny1hW60fwMIvIGnf0xITbSyjZiFhBfQchDfpLtMtUH1G3p3pqWFOx
nqr54fGfkcfn89x3Xc5LpqeG9UjaABzsUB8KYAEovxPekbBlUivUpei9+qCfDBhc
yjL0c3MLAjr/sYEE5RkMzGRXa4BUyLcF2BXnCnQNHgoBlruXfbaPZFma5uXvyKNR
7J9d8XatfT0jyJMJEdQPIWwrnydy3B0LrZQtvyGIq2TuF3pI6BdtT/6hTX/PaoLr
kFIe8yWbgZAQ1LTvbaSc34Dt6lwWCyeKjUVcQBbu1m6BFpPXG7clRDyE6MDBmdSm
sKWNTtzAknmjQuutdtcwyEmxrWT+UgHGO4OHXSBc+p24Or3UcIYA8dFdd8aFyyGk
DN93V3saq5MedyFNVf69Rkw9HLFL/WmDelVOsKMihA93UshTmXwMh219BzyaN/0c
N4ZHucXf0iuT3qNl8IyK0uZMZt8zx5g8agT5vDNs1eHo6XYgdkAdEUTM7csG/gAS
AO7Brx33JMRVZeXG0+VNH82C1mcdslo9BACEpezy4j011JCDvi3gHOpzMph7aQlB
w75QVD/oxFqMJykrDHwtcXbnvhKoL4EK76rDMov2+jf3Q6qnm+QePcbgZzuVEwuc
F+BCm957Ve0cSn1PU6eBObb+dClX8C8fpch8xI5J9pz1NPi2lkj/Oxrir1YSN2Bm
HIdjk1xcyabkkiunYPcWVu2AiwxWYCS38qLWd+kABhGWvLa0otWU0MI37kugAQa3
Di/n4rlQEz9JuMNMSPRYAUThCduT1k7FtDXJt7NLeNBL6QetoYmHiA3Nlfp5VKzC
cGeEW4J5mXH0XMdhLcwEene/lleMeks7LvCETEmG6tZXbIVE0rcRE2FqYM9B+gXC
Ru03N0E8a2GqwguAPJPVLogGDXvF+zHvaazAQsAVFVGvcrY/Pzka/N96l4KrHhwe
UOV6HWG3pv8r41wuD9rzM6Uu0OtIs8H0tqMJKS4VY6l0U4jGGQ5wJa1dlQ9zI+U4
iJ3G/VXvr745yOmtHKXFwzuq3jpn7NMdPo06R9ctRp0iTBANAMM1jC1hLlcfninQ
gXcB0jwqwS04zQtrbsrb3SvTWIZESRjkPkfJDP2zjgAWVWNzypeOUKdwqHIPO3Qe
XJ/nmFhwJCaKlsOJyXToX/FGKBVJFBvjHy/1n+U7dZjo67p+00rp1uZzILTSUi1w
v+Z9kxhni6Q+GacX4SdclDDrkGQdhNVHqzk+T6Iy90VXwjx9Dj0Z/j2Udy+DgnbD
oXvEXznjQ4Vorfd99SQi+Pi+QmoQiYk/dJMv0Egk5ocBE6bFgXTeYGE9awQ+Gs8+
CFVU/2nQMvrYSwhqsrsJ9KS6xJ/5PbNguRc2S0prsaxXBcF6XOV55s4xeCxF6F8c
slfPMxCsfNR4zcDVaoC7rVyrQdSfdPTXHi/nnrKDkdXYfPNxi2/c5kK4t7dhc9Im
hBr3Q1AwXmLBlhwaRRS4A3hQ9CqUB9eV/lRjHVOC4tgL9he7YrGwyTEsIq/YjS1m
aSznSN7g5uCILZNuSII2Z4qBRop818nndc6Tc8nu53HSHKjXbXIS7XmpwWbVO8HN
aCxKmfwH2lsddLqD+dvx1l19uX9c5/0TIWUd+roe4biP2ybMEOQL2EC0WAqgX+Q0
cUleSxzjAx2bvEL6AMGECXrmpnDP77I2v3dFwL/rgSTMthmcUBo1a5OmXP0JuMJg
BQgCmYkRJABzkPkycfvcTkM8P9de6zxyfBwqhfv2//EXiJTX64HH3fVDfIkDu9UR
oedNy3gqJZj6cURptXTLWMxMIH+7NYrQXStqFn3HqnMaLL5C9Isy/DrWuxw7Os6N
LyTDmM6OxKC2m0kcjPttDHXbYXEYAkZa/RutXuDoarQJ/36O4V3yunLSjmOmViQw
gW3eEn/bu78IxF/TnCb9vj1wd32v/Rq5Qxo+vyY5QcyGg2n4E0d/tyUJB3OhM6v9
+FtpopAZZJZBjGekRxW6uqDQCLAs9g/Td0c0cOvINSqYpMQNnApF8ie/gOB/S31I
sjomd4i2IrOUjJEebPGVP7jyastrEcWK0XqCRkDc+v0gXdrlCpuvnzUSDtJJhwvI
NVc6pl7mMrXDrQymwXv0CQutOlHZz2kWCxPYC3gWURPQD4BmgGwNI7iiQ8znJHfy
PVNjaLDfEdjtGW/cKdFuDtZz1tQhHS/kyDhmik8XYxN0yaX7vvd4ITCm02uX2c1K
DObVMuSZuWV34ZJmcFh8k8hqAE5jHhSR8nTqxR3STuz2w5dikVlgYgd0d4YvYLST
OIxNx4PIAbLU0qtpRX9eN6Z2b9GXjCGD+kWAV9jcyB6WzKcWJKlVqHnP21ATV4aa
3WVLb3kCGXaK1vKglViOkc7nRCnt/5Sd/BtbrpKLQXHD6yWUY8vU5db3ihHhU3aG
zZ0ZwpEL5sDgEtEDXy6O35HMoLx0XQeN3hMqdJ9UbjsO8Z3xTierNe4lFMCa/w/+
lLIl86mMCPYT6dXPeVm/E/F+PFdQJSPWoQPj5ZY08mgZKoC/wh4FLbfibCl4QYp/
Fuc7SKowVMWxm7Imuatu1gpl73gMJ7VAkJYNYtk9ovqUp9LZ/WWaPkfFYLI3QGff
nMwskPJdQHWZp2g/ZaxIXlrE8Yjk+XbNB3JdqSlelIdW87VN3yfrjT6fBFkJuORg
pQ0vHwY6CU/mag8eugwTlIp4WGcwI09hb8xgyWgTZQ/BwNLu7oo3RkRbxEO20Yrg
05qWVE/DLkx9torneh18t/AwmMDABifc/SY8UME37QkEpiP/Q2eeFsmrvKkTmy0k
Q8mNgIeF8NxuR2VGTdNY5alHKnt7gA6wnkexNtmPt0oeygSvMdJygXFrFFFxP6HK
72BV2UVVrAPVUDFOosug04vIPW7wV/h8er/t8YowvPRqRTx6eUylRWTsLxF02IRr
H4JmO5FneXhyOM9VK2tD0BZbiKaM7FxgkTGHEhJTDwgUgtKhpRQ/Zpj6hlMb/0ld
krBECi2tZzlVKUWwfEBRxMz5OvCij7juifUDjPJ7HQJupw0Yj0f+wyR0gFntj+L3
36gM9F2Ljq7glSUo3RMB6ygUJ/4YLhbElng+I2WAENb262h0+X10nfK0H7vGrU6x
HMEZTXJS5iGQ41VYK/dKCbxf3Bkjt8iPnEHrzeZe368Ps6lTyCSrUz+3j1VS6vSy
gEU8oHV78zUdYTAfDIAdprV84bf0S5Olln5+9nz3nIAHeWO6sQViH1pqZvsStc1L
Y3wJykJZRd+fsjIkUFQ0CYSVC+NHuaQE8iN0FDzjQm01IvJQXoUTaMyTvnTxQVOw
BGug1EOtOBupg/0ew3qq4/6j6nyqJS98AR8r7WJ0mrq7n/uueP59/Rns7mMIRbZ9
I7HrwXXKNQGyhrS0Xc7FLrUer2vQ63q8xMlSUa6uQGNXvCiOfdJI7n2xU1PKfOhX
kvAy4u/VAu5NI5BEo+BSM/N7Ulvn0LTB/yQP8Ts/nTGWBbCzzjOgdOUn8ol09UvH
qT1Xt9d5gKtNXK56y+lY5hTu9R4oGXrmeXd5MF9NSKnnVWf4ceicQx3/q6OOrmgg
b0paz0liTFZ9Fay5LSinACYEjFmzrga35uCL1ip+uN6dcdVQyhjmXY1hHcxTtPL2
CsUpL385gXop/v039sj4gYG8V1ejThY01PpPznvNecmOE8HxYRyhxl2sDlm4vEt0
eSM1bdJb5rX9ESL5PdDkLRMKMK1aJuC62u43TPiqRkZ6yIBvoLHNEyot/BEYU8vG
JuiDjyf/ex9uIGROjYpDV+BFw6Nq8iP2CWqvEPnGc0kE790DGsAva0pQX8g/zyS6
WGEwUmDBFw5v7e+qIklH4hZPkQGYXa6jchE4sq33VTBxUeMWMm+nAqdFbGO4otAn
rZRrs+BHcAxLDqbMUfitIVShwXcZ+1lJTKxn96/JRpNHxTkgWXUW7wJjRjvtmaMz
jU9/nSWLCx6PJ7LBGJMSkPZrqvNimnTxIAsYNpPaq8EkJfqWjJGC5beQudeSK3Wf
DCK0kspcAgVZ9dk7JyBaEcA1MU6ViOJ+7YMNfknTgPg8D65R1XjVpgB98gHLCnCR
zQTT25zSx0uefVCD2Njroxx+Qmwjb/A/GzNYqTqTLymfd31UxMXAZIuVPhHbmluK
RT3ECkeumixZy4Y0lsqpKqYwzn9IqY0jTz2q63bH2Oos0/JqTWTMydUU53CCZCvB
a0wl31eDuREOdO1vySBLBAISjkcxoKpbK1JYNXz140JjQEAuuaXzb8JfctN/Ptlp
dXUmQbe5e5eSSzfacTR5bF5XP3iKP32bm8nKB1Y3M5Ir7Wae17eHjmEx9cDT09Ko
9z+lNAVoAL2LtSODniXjSMYyTl1r+t5hghkcm9wLOCybP8/+KumATTKdcZ79n5mD
2aM5X5UeFFKqcQxcsc7IhhRtvM7smB+KD5UrDUPNv7gvjeVyq98kOQ312moj68bq
OHCkMihXTrEQ4LaERpCfyPF5dcWPPkCrc2pgK+6OnqC0i16eMD5Q83FqFUZOIsyx
JD61rX4J0D9WiLnEoVF9p9AqBe/gzrPGiELtVGMHRK7Cm8u1qtW0gM80RspT4/XG
lrdJsxmybVw+0lamsf+R2qLjc7fieeZPUAXMUo+1KfLTsGsDE39CcXeHCy+RqGlV
aswp/QWdSiW9/NPPSB/b3qt7QAHa4e7Ifvps/Qyyv1KEg/ziyMlfY3zRjFM5l+n7
U9+Z00jBIYSCxXlxDwL7byUzVhbBD6VpbgiJY0+4wP4ohi0RL3eXj7XmhEDOLRXS
F7GaBzrBCHVKvxiaaVgSLy5+Ue9S8L1igDB7vv4OT4xIdpvp7ID7XotWgDyGMbw5
FLAF86UFsXQQgt1EolyEBbORpCHxJhaDkwIsfZwX2T8y8IvE6Eyl2UORAWv22h3F
jJfDEr4iULN2dXJ36JF333Jh5mUrJ0zacm/Sc4+BtFfaLfWhuFsb4ZnGWpNnbcL2
oYTwDmgjoauszVsDmIemRqXGxDfuNIEgs3BSYuf0YxZU1NDtxtv2AzgH736NV3kI
9VJoc953k6/OhL1ddggshVgAdXKQUw19F0ihs0VDJlXTtpDMozYP9w30VdKQeGax
VXE2kn7Z+5YuNYC/KtfR3DxOkbAWW6fqqQtEVizXMLPjYrP0tE51KhTPAby3RpIw
Y7pekQzXLGwQPCDn7npDo0bN6QDB0dja0qKVmMWBFoPUD0h3UM7CfA4crsqGH8jY
mTxvC8lwTmDZ6ImCHoxl87Dm649In/LaBRNWP5A042WQ4gbyQrpS/R7Oa8SK/bfp
rOMFukZLE8nFyns+dxfF3KFW1ccH6oqwSqabJ6EDZayqm9E3DtmjPGceIi30EmXU
4g7ZW/B5zZM82gtxqAyNURc6IP1an0IeIKJCrHjYyStEku73BT1LJLZfVQjfAKzN
x8qxH048Dt/nYYvAu+0Pd7qxYffqGfgj/io3HJ6QiqJfgxzlZqNvUNttKPC6PzyY
2KiIxSzQCfUD8Svux/f1EfitWkdv1tsKHxUPtzkKLUXjLwIwwGLny5Y1OeHyY7ys
lKaxILHPFN/I2/54SUZFHoJ0h0pmD7ScNYrm7BvtAe5RJJ0EApKsXVP1ejMKvVkg
CL961UCDptx+CxJeJuaaRZGwf4Pps1uG7VcvIFfSYWfsj/PBWW8b8iWV+YiSa7Ol
Ehdo8N26/II5U9MqmxTJM54hvkmgft/BKb/RDLiAlx/zkjYz1LzrkDTNcUIW1+A9
VTuFdKJRdPQ3B4eCIJ5TNc9qypOaqeo3odGHG5H2M6FH/Zd1Xa409EWkwdJAS1Pc
ub8XtMZddLuXYBJ0yIUVxF5liNn9pp+bMV0AVVysUmUBjxo47A2rx20rDR9aSMPH
ybPyIGPZ4KDlfzmmHxsJA/LmOYUhAkeUXgQ13oOzoZnZ94YdJSg+pxwKpSeTe2gD
a/hOfo1hEAAl+DAd6ZRnCvsmTj5g+PSwiEOWHZft1AFkk/+0f6rV8L3WNK8j5Am+
XZhSP9O7xIl5orNyCuIGN4+fipbp/uf8OpxdsS8sVpEf35EQz8MvaS7GA//rOGVl
YcFH9cZul+ttQpwc2OPH+m0hNirFO9QGaSrQHh/it+H/oTbnzGOI9ZIGnuLXox2U
Y7Cx8Om4emNNjZvZiYu4qJF7l60KIRBehDbEh+c0T2pwBwdET//B7jtBZ2T2ARGR
U4qWX25KI0FuEnr+BK/a0E7t8IKktM44SBJX+zsiPrlBmPXqLEtTBMxj/ePWo/Un
P386PlvCl4HmSPk/X8PYs1X7AzC53Cv9aAN1AsV7fnxRw4BwCiPda0cII4ZCFPZT
dEG1t2MAa2APP5zta/GdrsE4gx3haFbybhoWQZAV7a5c2kR36yfmqtpPY6Wzb6w0
PpotOiQYuOafYvBq476Mkl8dOwmIEV7MiCIY/xMYxGhrWKqAzhxB3Yhg1f0+2A1e
WbEOjzNeYgl4zQHRNsoOm6ni/sBcTIZVboxfGFDQtRMofVGQDXg76yi20KtFSjiO
6Ti+ptqV7LFMsNMIBjJrzkju+n+oL7NSfGWF5h7Q4olXnGBZLq14Nwza/OW0gGZ8
Vbx6WaIWnV7v8PP62NKDBuZQe930SU0y2URUx0lLGFE9yYx+SfNl9neZjT/aX0Px
y4d/kS9zDGAN9KkVI6zZTWMnDVilJl6HsXYbrGiIYxDDf/DegWCiNhE9QhVakcvD
AIcrSwQolKdfCgeYoUEgUwzfSKku1TyS3neHYueIaf453/ABk+2FImEgugGjv4Qx
2auLAz/aX4c1ezdAEjgHLI9WvYyp18BMBIB3rrZ9kcRaplJckkuHJDYQECZ/G72m
JwaOw/XXVSKY7OC5ahPEmdnEyeohHE87VYLKLOCSlkw+Xegkfcw/5MFo4PrHsQsZ
ynNd4aiLeRcX5MhdHEpJXxAY3TC8DRFzC1NmGIpPd/lCOED1yPi9u8ievwN9zo3P
7cl6yD7BrhrUBgKNhmLiw6qrgq3SL5+6oCKmKhYeSCvVxGCql4f4/ah54nsZN1Uv
FT4s7Pz3kwfExuaA2KXtbpXvZVjd+XZKgoGyqyKPiP5ypWRfshHVfdj1Zag8mJF+
G0d7hI/RhuEyoiapyO0sJchRPMiWDGeB+fTI3LZFWspIUjC7MmhvoJ9tw1YiUphe
tbP+z2ZCpgdNUed4zXtZBUdWVv3jBxKPKJW8iyGNrcqvWrjHE6in2DBMBKqxW3Wn
MkBRYkMMEFMmsX9EI3yQhz0+08EvNb8Tg1+omyyirVJJLr4F0SDaCbhc4eMnpDHO
L67etVq6wqcgp0HE81GDLzR3FPzucfzqE1LQMpSKH4sEzGfy7PAzF2P7HWi9nsEu
dyP8HIrVxRGZDvEzGvCP0e/sy6TQRgBzyq3X41NOT7/z7mY1KR8Hrv+qcadgQF/+
pGmk1tsNTJheHWDRiXGwq4x1rPPAbsBCxTr1ob3LbHOjINgdAYES1hVo2FXFpNm/
cvn8tt/rlVRbzRFh7LtDFfRgOyw3GByCnZlQ1zaxeFN/n4LriEJWD+fUvvACKD9U
GvxHcF39loXCwgmwrHPhQ0JxxbTC3IOvhx5hUmFC7Pdaktt1zOXkcBBwclWiPANi
+ZsSTQ3/GH4GOX+rl9DVYCkcmVv+o6FUmSjzEpAsCw6Us9uJENQVHPoQG5sBUNes
hAWqivnJme32s4i4l2ZAe6Z/NqDr3OBdhzZ1KbyXyDCk6qX28mQhhfS0EX4siVPF
kx2sGzsz604h3vvCHEu9e8rrtpBb+RnULEyD/EbQXy9BtP/TYhdEWPpRuCeuQ+5Q
phFKWcAxc7Nuikp45l8oY5ijDlFRCXNhbc3zrajsHBlVUCZpU2MvP3RpI4MXjPlG
vNUWENytVK557R6BNfZ6yXN29Pvxqy43hXvR/STW+PD3Np/HmyMj1HQX2TNqe99F
u85phyaWikZj7Qyy/aQUJi3Mot3pNBEPCQFpKFF9O3gNFudDfgSdoMB7/cAtTaXt
DlwjV/ht0nBx0e7Da2mje9aZxO91uHniWfed8LnLne4KMg1Z0dy7WMm50Hn8vyde
HXl7ekDuSNg0NU4aVgBRWwbZSKRM+HVZt/l9GqiuZsgcoUuQWf8CSwQraFfBNWmk
Tt8jTrOU2MOG3U2px9TAVV+h17ZcfZfma7+aRV6/CdeMujP1wnBEe32hxyo8lX4g
0hIEXSvQ6usvgF/1yzj8zIhyKeBCrUJouJ9+Pd/8ku+oWZy2Se3RnQ4Eos22IUcV
f+nSAfdyjiXmnCIeELXhJgFr7Q7hoIH0zsVGoH4mEIbxR2/+vO6+eCe671Hj0XRm
ePqFVaitnguGt3OVznQ70i7qt9jpl/jipzfUE6iMBEBduQ1Ws5WT17oP9L7uYZwK
G6DLksp976E0T+i0Mm44SRsTLXNiFijzfagOwxKvXJbT5dfnkEKvREwH1nuuSAdR
lQVkaorQicfTFUtXcjiw9NO0ohND4CNLSVKRksenNW1JFx7iDgSPLd15U/DZ81VH
n+Oy8Sx5h2wFkbcM5Gqym8PwZXi2VQDsAaIr6mdlYSuvdH7xyoas5yDUt8m1esWB
fIPW2ry2h5yqZFIUIFuDTHE+xsH9w6YFkx198pjxYNcmz8EVD7b3Zfi6XVZ8tWla
Zc0KnbsqZJe0e40OeW+s2Dut3OlVZyglaTBppzz3F1+BnefCL+hKD5wXrcpmh9dt
HLbHYd5iHuhA2hcMlrVzPyzJkVlQ1vyRvluYS+iUbr2sgzu0gFCU/7QvyEHmiY+Y
OoIrOIsglJOxjEQcVOgENdOPfWeRaPLkFeVU3FzkabQebp59UZSHe5qVk3UGGAbR
CnmXMuZZy2gKBZSHj6erI0Hkg3rUYrHzg7CY1OFpkW35JB1RGGflf077PYBdDseh
EITySRs7A5u5Kdcn73kjrMP0PVYiFxH+E/Jn91q27ulsGSASp0xydxt7wpvH46SA
eZVs8NjyBRGLum1Q0vvcCVgGvfIuxQfX4tz0c+xODNagS4ZzvjMoGwbkMkOJKR8x
Jmlg9lskAll/7/mVeRIQEsqIsnYuTAp8i1BWuBaKafiIHbQJC0PIKrQfkVL1M9oW
DtgK7IbphXlxizNJb4cQeWlX2lKvufEto6OqGPlqFdH2nWByCzyoH9t4THRrXxEz
VVk6iYgZ/2GGK+hzFpFE4WTfeuy17UMtOCHzkAeO7/qhJtKhH/lNi81uSLLh+O7A
/+yNBw4alJN+Cm7j620akLfhFmlMtyqCiI32n993ooEUTyker16x13yHQJyi4z9U
VprG2xXTPpOdDFSuCqV1l3h0J15rgglZAvobwwLpZ4XMupcbGxbWEGe9RlPCVDbc
RvbMuQfKfWkSxv6tUrKEG46gMOJ81sIEPffVdNmHeI7WXAuEe7TDgCWf6JbAJvw2
6qJ3XkP7GDAbvcagf3daAlOg1/Q/9PQaHcCRkkKnZWwHfLznT9NeHm8rl0FL7NIe
2hC8i/RnO4hrhYPm+l0xWOluTB5s3elcpl27Q1EQUtHUoiZjbs++XR0IvS929G9v
qasQzk1Gh7AxoMo5DAYSumuHdyU4S/lfF5U5yaqh9ZsokP/iYmdQX8U7nemROXUW
neWEJFST6AGdFWA7I5G3iHen9I10Zx4jaO6zcG9GATYxRPGEYtp5P74wU+MQEqCU
VTZlDxj0V5Wkcwuyc6PYYVHI/yNGVkZDls0NW7xA3PVRTTT1gLgtGc0chJemNRKu
6JHlQyUYAJnA4lpOpKoPOxiGVPhYtIwfiCj6KMDwixTgH+2mIPtMRBATHtErLoII
a2YLhbtSAfMEVjH550huwxts/SbES//W48dESU9mTwWpZHluvPWdDvf4B7Rf59Ww
9+jAtxU0oXdOvFFIP74t8bKPKf+5rLpASOrNcFhjxk8eyeaBEjc184XUvrZJqoZD
BrpXVQtXfGCLjQWXmR4IHaYR7Nw1I5cXZzBwXuMKnb7boHNbNlOvZdx5yzz9ZN+p
lWdQe6OiFVMJllPYrO3P3HPbBvyOb4ylato2KLrzkJ8+ciGWaVtnso8PUdgjJdSm
SbgU5eK0xBg0wvJg/ueq91+tYTB8a3REJ8wIWieJisQAZrgNC2TiA7AWDkthlFhb
EhuDLskLuxwY4GBq88mEFaSuGS+XwQWfZ0qZvWclWwc8lYNvtjQ901Y9nxAjwwW3
/PBbaaKpsQWFdSRbHSTN9fgzu3AtZ7f4gLmTN9RbxBZyt5v4vV+d4/89MTwf9VPt
8gaTEge5FmafOVJ9D5ovm80CWyb+yN2ar98JzP535oElY/PyhdAb36i8t4fASUWH
Xr7eYck5Q7tq9osRjSbDKnd/kWYIhxFNNKDIYPpc8d1XRb14cQ4EjEn7QuMxj/Mz
GK0OlRD3o2D98b/QT6H4qe+nTfoRb5+6NvUc6yiiwNo8gXnK0ZnEXRUrCddDlvZk
XcPiUETDsBqwxAiTL1+gkr5KYnK6xaMDAf72M7ZS1zW+PMavmtQQLgX5A9U+NDEP
G7vJ8qp2JuIDvSlHgggsphu6qGgt6Tpr7+RcfwyhGr+cPS8G5xKxvfZQJqmdHaXh
fxziBOp7UW3t7BbgmAd/fmxK8MViG8fodL9mbX1ddBH21jyoE0En5dwB6NKaW8i4
5JnLOqddLwTpfUy9hgvGMIQKy+jXh0rAoT6vKHrwC2a+qLOEsfBa5atdY2F2Qysr
25U3AXI/gUnC3yRyrNNo0HCwPsyv2ZEJSNHTwgBiTSQNyQsDOmDH6OnJ0tsvt/M9
lSLk948g0rGp3tXquw45rd9qoq9KSMFKUdveAuVrGBYDctF8yOS5fsWsFBE4PL2y
a6q9kYCijo2geVQft09DNF1AXwWrAC6PkfDl+N6ZnHZ/LZHFfkjbjZ2CuJ6B921B
wqZwloaAaGO8dF7w5vNGDNziVuWuTZ7uVWXj50SlxrnIW015tWLOyECYO358k/Cr
jhpY81afoEzJgFOOdZY2+5qpmdbOCfyGNYB6TOrgnUmSC58eQoxkeq6H0V4suKlR
Cds4ZExpzDeZtnOYWwKGNv3ROB/DfUQX+IDeZn1QFT86BptjN/0JSo0qiZoP8gJU
W9OvLyRTGta09j0Z4B/CDOjOv0klaMMIEDnI7dVx2/ZXqBX8l95iof9BTYLI0c9z
xIXZRcYaZPK1JrQy98Y2Z1bmENkKCa7Qdb8g6bBeXEKxKdJ+90NM7drkYjzWjvDe
bCWlv/soBHhQYe7Slkkw4xmaiHp4TkRJTE1Q9cMybCSh96xwyEn7/teyMEtjN7vL
+6iecbHo1EJFZg3oMKa4Oa2YOLjArZqaPi8tb444G+ROzzYnqL6u8/c+EkaMJYNu
8WlPLo4CJT9JSR74gznjg2NeOT7cbllotiTt0VclZ9G2s0DifZSANZTODG0FT6Ir
F+nhjmmu8lNWjObWlwsUzkYOICBpmV9C827gCEk+O9ZDAJZEgRmu7iwpgsJaDxxe
hhKM9xdkRGDptXavKz7sY/5AUV6r/liFzMKZiRSHpFob65dOCJZprkfE7HO+RFeW
Kzx211ErceHt1RSXF6P4zqsC8n5WyWt1DGrnTKgyewMDqWv1CZJEVNMurmMAoNzw
rTrF0iBiiTCgoWnmUzgvhWCiNYa8/dpP0Pe3Leaz5CmxV3jCjrlFEynNrgm1c1MK
2ZeJk+JYgf6pDpZ9Q7LS6BvjImGXgUnHqwBeOZHeeuBiXCf+ic4N5qR3ZJEtg/eg
TSn0eIpvcsEKciJgoAFpo4uoBaqei08k3r4t0/3FCo0FpJXomdznb0wH8LxiT3Sx
zMkEndc5stDBGowNqJfzjizK0gj1plSeIvbH2Ac1A27VQNgLv40A6F2a7aFCD8rf
ibpKQaZpYGc/WvjW45wzSUhwd8x4c8X/OJUtJD0CKlK4anjYBHeHw0X8L1ULSXuk
M0XgNe0yqylk9jhjbHKTc5wGPSUju6km1zSIWuPKk0wTbGFv+tVHV+HE1AmpcJ/S
MILnwRSC/XshhObATO+neVXYxoDQeGQ3VjW2VHCRdFYSmMq4+mYVXo934kGAu6Ya
q5j+3BLpgRcJrDdM6j3tJuN3BaiRNAGvBE9gNCp816CudpI/t1nlFC9bWC78UmHN
1jkdT/HTZvS9+8ypSEtG+cwiXntCxyHho7tDmyzgAijmX4PZyp90n+V35wOZIosC
pt82UZ6oMYOYyxOIqo40JGJf+UMPWLRlWJbMcW3N5TKJ2v6xZ2O44njaHdPBjaaJ
LGdxEer6K80OlxTn/t685K/swQI7wq5Zd1Rnmn9RDtudM35BLLGCmpVp7n5+9M+x
riSZ4k8/t3VMCL6fda6jSNVfSjT5rhaGC27LZBdWL/hz66bJZsVqm0a1LnoFivZc
QoGH33D/m+oKPQ1mrAi4oPU87UphjFuBFYMtC5oDAEuG6aNHWltx/pQ44cpbanMD
C03e18xTpgN0avnwC23LbWmwVLnixSdYCLiG0wX0ZwU2Su0yFGuBnUhVi80Rjz0w
53IMsYU/V2Y7+eo7n+UZik4dSXRAkTJiog5J2BLuHDuGSK+xWTLmaZPpQ2VOxgby
WBJzt4BgB9amrTyCN0r7vzgjTtgXuxisDctKOm9EZ/u0hqGuLYuhAgds/0QlnVZC
/qEMFeIuep5SqsvAsADJri/oyXJGwil1/Jrc1tCLzOD2qWnwe4aGwhtEgdXv/+SL
4uZHkTl/LjPIfGj04Ont76TFmgsmRfjdH2ftNoCFGZeua5HkXJzJxciR6+9y9brV
kdWG0RozHQ5XBujezGIHQk+PRe80NzedSlHx+7vLf0ZoylonG0nuztloOfY//tpC
SptxvKPHIkX1R98ZUbAuZFIaxXjWAYDVgCJlI/ULiixekoo4Mu3/7/+0EeVSvd33
D0Kmb5xVSlqc8u8Lm9cFL4bim80oLZH9/BBEpoMLFi8zqjGG2mvwC9DDY45p4DDG
ze2fJv7bEMA5LtVhNc1l1aAJyzohMrs8hAoTvFxJtvsLXRo0KSSUFC8+frA7lrN+
PyMZ+/T7P3yBMID1/Ro9Qs6SMoO88IYB7QluQ+3yjo8BYfd81VoCFl86YgmhImzn
tcyBfCxEKSwedTGYukaQBuD9fa9aitGrdKRnHdBsrwl+Tadz9UIO79qWMO+3jGZb
jq0C/klnxXdo5ltL7cMiWgz5YZQt2bJvnJX6ZtEAJR+S6zsA6Ld31XeyQPm2KA3p
26jRSO0kYqCgTGdNO0dc1s2gGCCg+X7ZavVNzyZytePLcoJQdMq8HU9A15454l4b
SPKMpXdnPrLWEwJd/5acDrEodYYrDB+yQcI5dqpnPNm9f//ykbcAHTDdNhXImvmE
RO6d5QpxqQT5SptoHXc/PV3M/Gz+PQmZOr2Xd/+pwaLTwixnm/J67Mh1MtsSQxyG
1oP0/PxHKVKCQ88HzVW60vhYszCnpYMCpmhtby6FDGxSWB7wS5QuDQR1xRDvJxjr
3OyPf/AaevIRnCVWO+YUQbsSaQtgzwhNGCipvI6xGk97cdXuArMT/09gQHg+dx+5
cBsG8Rrydm16WgPZ3QbcZTqyr7n/t/JVG/IkZ2WKKv08WuWVWQVA69DZssDBOgI+
VTS5Tn60i49Wl1iuSIKzbA30we4cDQp5FEWgQ4H9n9qybCKx3LcZQSx3t29DLjdD
nclYQRDjwF2cQfWdryZXCP0tIhrK5pZLm6UwPajIYkE/Co6Vn6g9vgXXE/SKnT7D
kaoRGpAlFJYosEosaYtnhu2GVvEtzouyzf64vLytJVeTdUOHDwTxc45DnqE4dj6s
rRHF393fak/D3UCmCJNoTXwjxYGCjdlLXSrr8HhSeHiHpN84C2T1ZE6vkrVUpo5r
cfl113ft6nfUzg63TUAds0Xd9WbtTp5MVP/V35WWRipgFJyc5dFpYovyTLMqfK5b
LiuCk3uv53vhZakPb61C16WOPctmO1OlBdn+F+I7Ewc2jznDBC8JXBzIksqRyUw8
UfUM/j+WzhXp3lkYD9lpHzo5tnHWnRhV5Er6NhLEtBo2GPBDFzf7wq6g2ZFPM8jl
r9WkK1I5+BLhiltrsCpxFjzcvE5TbUByvVcR+bzZjq5rq7j7Yhk3UDfuiB7LgO0A
N19EHj3t1rpEQ7ctS9SxCVK+EnVushp63fGN29NQe3V9iVt7+R9RwMzy8OZJo4/Y
YQG+tIQelUA1zUO3/JYc9ghJIxTLYTuxR3dn/E8T27FigYjmcmSc6J6GAGfjyv9g
SYzVfIK4DNC10FU3n3Sw9JZYmvMZkWSOrEoMnhs8ODBlVviL2LxuL7DVZLJ06urg
olfdlsze2ytNqqADE1iVrHrS/gLGiS2TpY6XGLRi6YSqUL8NTd+uZ5+aUXz7DAJX
43MNas5J2wpzXn/m6ey5xcf+aAQtBSJhCk76cgUl9ZkXL2aaoQsh+Qxaggiq2FKK
lEr/J3JWJdyBp4xb30sStTPeAxhKUU2eht9GWzAto/WbqZxkWADapOqNyRPGfV1W
+IeeJw/E63w+dj57uORSAx4v1o1qnHP7JbMEHI859e3wIf5NxQ60beO2PIbQ0JNr
pTQvIvQvs+NLQGm/UDxVWvWtLr9ZKEdgyHbqsT/GY5ukHpQbdOh1lDBLqDMgvkVE
28+G4ScyqkK7EhUJAEZjQUMdBcH/JbkLOOg3m1fj+FhnxE4dQbRxMvXtuGQ5xiSR
KbZG1niuXmuetyFfG/w9Xk5012EupWQoxEOiKLWhLB6zMRALkHkAieWCgjf/Ndwx
nTF9syBEPzwUZG18cR/mf9oBz8MxDhWzQYd6iGlPDFtTHBuemkvGpqnJXnzIji1N
6/ACXpnS08L+f2gcqrQ+MTFhALeG0mRYNjdQY2gy9ssyq1XT8j9tKZpNadeR6MBh
i4qrCp3ghNTMkUZFrhcN2NBXROteeylfVC55yPek0+onGlejxNhxfAW9Nj9ihMKz
Hc5ZLjRacKNkYKIwZXDY9Wk8gYoXjEtEk6pHsBzgGIa1sAwjWZqW8S8SPFJ1w6Lb
fqzr3GYiu1fBdrUsuArMvMiOuPh3l9OSRsqWZqp+/gCmNlWHm2qYWP9XtKKaukAx
d9Jdtz4tDOLDaALVl5lbjMEIx+AtcgwtMZVzpQ46O8d7CrVJUQEVmW1ODS+YxTCz
vRFEAf3VErB0MOVHI2vx2vNYM9WDPp80Qm7KZAjH/EsZ+WNo+/jPEH3m7KcRODF3
zzgyXOsB0814B6kvdVYl6QvJNRtlSNO+3gCeHrpMlAZAN4Fztpkk7J0mV9iri3Un
n5b5EloFMPbWhA0BiyD/kG8HnmBQib+gFhuXH9o5IcdlVnnc1nOww5575J9KOAU4
5hFJ1pxQ1ajzraZPikRxrKc+vZDcr5MgEDyxQf7aoqqrdoaxlLC68kdzT24kff6S
X4KGBduxSM0LfvtUp7vnK8m57hjoKDNGuoRbu45ZMN2PbNvahOLp7bj+Gn8CNjt9
wA2nI/EFALoSc5IoJn8uL2DACY9Y2klm0g7p1/DJSOMLU+hlz4kT3xM8cgmY64LM
EOILB5WQmdCHlIZb4pEdchnUuozzDP5Gc4UouI4ADO0jWfljeHE0AOAvpFOG/OHR
5m2CnBDa7NGITFd42O3T9I8204VZFPfScRWIIBuUO5Q1Jq+bx014b8M5Jrx2luBv
ypImcxKHV2qHZ+F1VDWBLntH/ULSWI6XcYf2nPmf/qHTYcCTwAO3dBTBaio8Otbr
k0IsTi2do1mG+aezTAYL6KIutMljRj3fwg6wdk5vYkjzIYxFXz6yBVwG7Y6hYD4x
iO2BqrZzpbJ3GcfAIdaA52r/FKy1mv62UBxjSCndHr0vzQn3vwephJ2qAS8DZFi0
XJa5uK+J5l4vzgJ/8pGHqX6Jz3pfdIR02JfGALy4FlMnbeHle7QdqTDuaekkwH1x
G+LNCUu0b1yccQDT73fQfFOrKMbS1dPpf3CGCvsz7iac4KgIsnboyCg7WoW5Fu9z
oYbsBTBwCfT1im6WOyQ0d+eTYvc62uG2LApJEILs7x0pBHi69yjQVQ1GdK/vkpwT
T2q+Vx6gOgJyGrKNBI1t3UM/qJBrHcSJGwO8j0882ZPc+XBYwpAmElYxD7DJMDIE
djY5xU9Lbn3skDvrOhhbKswu+v5NpmvkVlTNUr6dXAGb++a9aByBOq6QizQm/veC
5Iep5LHh6DG5IsIKah/HFRkOAHHAb6Q14SsKPskjZ4fjbHfhh55nF75dwFdwOZFr
ABOqnEm6S8hiFZeJItCwYlleqVEhpMxpjkEmpD8LoJFAYbFvRMhTUTHSbhk4dMXs
TA0nX2LdfCGxrmDnxrbH54PjsGNv2Tal+jM7qKAThwXEboNVs6Fref3krBxTvxj1
FIFVLkCW1iFYmVlVxvxGUMni6Q2NPqIKbDldD/KKkpzlB8UcnhpRr3U7ubxKIIzg
qNKb30yuRuBu9LX6n0DK7hgY98yKBjzqs5QMVzqM65Z50pR5svmqvJUTB7lXFOdz
t1xh8R8aduKKcP2rNHsh3eqHnMgZ7yPKG9sZHh8r1r0WODSFcC5JzJqfxfyrfmXm
x/Cw1l83k8uSRAz5Jwa+OCZmx0URabQEVSDSOD62hie72zic6IlRNe0ysmNlxGyF
8DL5YvOLs+KEdq5ALiZSfDD3BXkLq6wu7oAg82x4vX0diltM6gdAG3io2i+Hwye6
uGAbJ/Ydb1aMogZywtA1CsutXJYEsPxh6qnWX8Cvdn4FineRJy4doGs42R+ogm0S
qDO5zterH8ZYdiqI9n20lDrVlRHQO2o8s+JOKlM76n+JmfRld2K3WoWknYZex+hH
j5reIbNlJRlvJHw/Yf+pJR0sL0Vogz5r/c0PANl8nNrQenupggwb1uGZUHCbT/AH
pcAr2vazSB180SFqsOf/JkPdl8N5Cjq8xQjJGkMHyGmlbfPJGcqUmIPboSGV57TO
hrpgWBMwYlQHEc5XoouvKaJp/nyr4UcAN52Vw7TONDgKlpAs2tSRNqaQJzWoDiAK
dT5K+du0FPguZthW05/dCIlqzXGtjSIs0fp39ptyN+mW8w6715LoJ2Wxqq6LMix9
o5mTyNaPHYnZOajmFTsph9km/gtcOd8wMTie51LVXtLfbP5kmmGJl3hojR03p+SU
Qzj2m0JGy3l4xyV2kH/vDyRjEoXS+Gx3kHh6PBqKpthVnMmODnruIoOryNySleMA
QWWzY3ml0sJUCQATE2Oa4sSQsG4avjaY2dnc5b29+4H1X+jbmM6TGe8/DMUs89vb
NAhavzf3uChIwNwubnCOStPsPcb2yOb7a5+f61AAZhTJ0tebh4bz02OBApPqN16z
1cyWycT4eBbLTZ32TqQE6THTGKgYgr1uPctE7fsqYZP+W76/l2i39GiepqyBK+Ol
jKbxwr5/jxtpPvxy5txDA9WWrthYAZtzD8Nmx73md974X4xnQWBUh6S3wB0tQpTb
5HVCNP6Fzmq37bVMp2TQS4SlGyyxThoWcoJ9JuNlTUKKvDCXmMK4pFBHFdxS0lY5
yb9aw9r8z3O3fTr4FOGzlzFc3zbmfZlx/w1eZ6gC7jSb1rYX06GtV+P8nGjqWj1O
FTruIPtkbyd+1CQCTbfwX/hBadYM+nQtzz8gnxKlU4qfDxKxyld0gRp5CpuzyMF0
6mfsjgsuxUbd2m0rS6+iv6aeWgtufhG9N25A3+tWpQCaeqVI80JcqqIPfRi11nb/
7hSd+45qgwOBB/w4H9Zfw0Y6L4HkT+w1ChALtzluMCyoGPjyXg0kNWJiTwlPu6ro
YsyVjseLd6D9q8nF73XyEMawst14l4p9i20/R6WvUsYHdi1PXb1LN0CZUTzbLu35
Dw2dzGJ/sXwgHXE4+/L669G1412BvPxAA24mU8lVJdIdMGQfg1+Hj1K+QE/oMUpm
8Q+Dc7K4Aj11/FkZuEFCobOw7tU02KKQkf3ETQfT3r5/qTt5JT2Ynceyq0hO/Z3G
7iwHMeAVOsWbvUp5GVS1le/iP/Jp7m+lnbo76wGMycwJXdcB7F7y1El9lOYVHZGo
lNlf6aTDtc728Lr5YdWYQpQY5Zqzy6TS7VCgvfoAVmsM1KmA9OtZaG4YDJdiB3Ih
Z8uYxk7QM7lSTFbcLd6hyjA+orGyPRCSa8g6g6VUs4XkyHAE3Z3gwAk2SWM2yZJz
J36ym2g/uwgGbvq+AnL8V4G3iPsnfXIaG38SYNeB9VK3S0RZy1FfxJ++yfyOR7Jg
Yygv7CprWVK4BWsDM44fNh834YoDyNLzZFdUHR5U2A+d5dopX52JEMHOgNaMu/fg
/M2L4yg3zCCHXzBBt8WSIFtl7o27wOSEB7JzQ0YNNUvPlk3tTEGrRnpLJam3TXn6
kYjYpALfe9GOoAMAZeKwjpu2HiPk4xx9CTCDWHLPYgRm8WdkWSSqoqPYtOCPLL6i
uOYExTCal8NYX0wSI49Usm3cx6fu990E88AC8QvwAlQ36essC3BpwzLvEQ1Av8w/
+wnSfC2kPIEnZm3xkKT9DJvhNprswH1MW4wHrye15r5PR5v9m0CdR0rIxPMlUZZU
UVQhTCYwa5eSUvDMfDgGi3oAIagf/30YAk0yuAnkYruQzxrknNWoPig9zlaT/ukN
jRt0rDWZI7qUGfvZ412d5/GF+iXBsHKL4vPVUDGZYoeQ6gk7P3RVKM0BSN73Vq/u
qUP5D8kacr3UpCtz81k7mo1ZriBCbFjYjfzGjScSK0D6Hq+SeWOm0LczjQs1s5u/
73WRtALsVDhYwCrnEBAYZS3kuWlQZL4lmcYLyVHcWxFIobD4ZiXJjQ7JybAmJzKp
HA6gdOFM8hikYYShM+NT75vKZNjX7NcjkAh7NY9YHTXfaJZcQ2CfC1gqEVt/Oer3
ijg6+4iIV47GClpjLZoLzosSHIve7mROBku7SfWeyHl2XMH/NUOpAW5abP6GnXEx
W8SIXSNraxDlmjQOM97dc3IuDf4euMPS1qjcSYGhNnYe/+bqFVLUbNaxU4QsogYz
WJQhQ4Y5ErtEMmEBYrpS9TYLuaKtWtIFSZrHW+pHUJi8TlVEmqvQigc7qim86JOr
4uomW1KalHV4ubSW2XdbrgDSKW55htT0z4P4LqdEdz4R8J+LKKkbBNXWJhhzV4Op
/ud3raAiDWOiV9NxwqAcKpDSJ0QyqRJtQ7X2/zuVCZ9vT8ApQGyYUPfv4wYvK73b
knlwqgI+f6QRH9eQ699+sqcFVmzSm5R/13Ud9IrsdrOdyzGYyCI1mdeZv6YhWDu8
cKhatHvwK0voKDHNIpQyJmH4Q7mHmXkDdzCWBPmsCb0bwx75xZR3XVeCjG1Ds6/J
7EIjPvXW2t8EmPtl7iX+og+URd7YLhj5HjZVj7qW/BZcVcjHC39254+tXCYooa+0
bLmFhE778/zqsOqQ6jQdyMnVy/F/9IDkuPnvpf6+V4PGQ2WZTdkVZ4rNqyb9vyoR
MGb7sVwOrFCdGwfbIS0sc9fQth22YYgpVM2XvOHcHGd7bTtQoe4/kwdqv7j3rduW
tSqlfox0pGgIc0rj1V4M0kktN+yA5dy3nGXIF2zBUxEIwindCxSkRx4VzxxXL6oy
UxFvnbHRdJr77JCByuwiqAprWoX2IzEb+j6m/LLBHm9JhWvi+XE+d4ZDavshRb/b
nq5ppJodB/h8jpaIC/dVPRSbgN/g78VwTh4Yqfkv77WDbSJtF1HrlDDKH24gK4P7
o34E4ngok7bwpMxrueEav4CzbdL72cFFV/jbSIoHuNk9rV2/R9PPJv+MRowYByHg
KenVzfPfQe8+Oyfroz3YlYrT+33rnDAI/WHNIBi0qGjFBOU2Yd7Q5aOjm6XX1e0h
gYKmQXWU37P3rM2FY8cPxxFzK8B0iAnKLiMTWPynA6VIF8n87QB1XRowvLv/1g0j
zswusy0TtQ4oODeT64Q2hsmlMvHWzwAbMvCKsVouhxagsF23OQrwnp0CKT+Oj24A
xltyAjqMIBC9ovepH6iL5xzocak9yPEXE25Dxsxyk73R13cD6+ieg7eUU4z+JDZE
z3ay+c5Wgzs1IKwMu/BFnajhmIpx85C18G1ysoVWEwAKSj+4mT6MK5Re2VeEUPDe
5wplBxPZCdJyjZO4f0qm6/zI3buS33OU0CBby8uM705mQXfp/q2vLofyIVx+FRR+
i82v1QuUfIVE9Tc3ciwZAL5l47OfrvndcvbYqO9cLj8AXI9Dzu/KR6Sza3P9l519
GzmTcB9HGnU6dDcp8Yo1rWXrO/xrO28yHyWb4XMV2WrOv/JqnEbPLkEL/lIwwsiq
CqWQb1AKsSUrI9REa0yIUs1w8PG3u5zuMFkETfVxZ3rQ5CzyPZ+PHyh/K2OH2G3l
9BCeGas0Z1XqT0xd+o5lWaWqE8dWqv8yvmxQoriMGZAgxtTH9lXIqqCml+Pu4LK2
VEWDw8ka0/BL0ViQiYXHm6aPCRV9V8jCQ2qBRIxLBE/yVGUtAvqujKlckyjvNDJJ
YEjJIEdGmTQNhAMwaTvXU6f2nRQp9BgVk/BdXwfZLxqyugwleVzaDnGKAtEucfO1
qqjlG+aZNDws7wMHL7ob09ZzDRxsyT5ru6eaO1a5CRL+PAHWXIp1ZWIIYuJCWZLg
WtfsVqkM4Xo1yHml8Yk2g9/pX0VdshBxrvwBKK+BHaJuVnMGVWmYKIertAoxF8LQ
/sUi+tW9XSK8DUx9kwzRFDJLf5rcyRPRhq6p3RFpvpJENH4vFEysTS3CVMnCCugq
OylFgllTjAAViP24aUjyTBkNKd+VP9nRn2oEgGipD6pJI/l9t9wU3S/RHnSKW1L5
N4q/4cohBONzIPvDavgLuNr1bpE11Rs8WzKzhqAj5W4EdRQ9mefgwjNnADAd7tRQ
BlQGBnSDXKxdLcyjysj7SQTMl+jL5XGJIqgvpWs++L5Z5225AI0f4T76xzLRB7x+
E5IaXURc5eYVYCu5I+oJdxTblewQRXvnMJcoTLpJ13MgQVrLYV7kUXRuFM2DCzPi
/m6kqkbN1VA8y1oZR8kF0SinE74wTdLznd/qorbxUQlqih/PQKee1Y+hetwbS3pv
Cq7wGxPCqDbClTYowNyoHPNrnNhePx8/52lXGpXmmCBZYGRNTGggAEFsh83wUc52
fbYjrUpVTDC6rnL7305dxijIjnYjx8okWPPv+5uPvu/JMlwT+qLFhFJMksZbSiSR
tvF9YeaU3MQQBwvqhtIkaBZ2kre8lkGzEb57iZRNUnrQDmJqfZHtUtdvm4HJM+Jw
zTQvVOAEv0B1+qXxXeir4pidbdwQw6TH1I4G6POLyrWMltcB7k7/UMLnv1NKZJVD
OliLliT+rwwMYmG6jvoMTWOFiDi7DeGumZnJ3RPmlrVALO72qWv0a8CPOKj3kkWD
8c2Mivd+1ktdweILeaWi5kjU/KLNHkcPnzd/FX4efX6yaUViNemoVvTCe8ya4kC4
GKcavBH81tSb/56BPjlc1sDbyAs+Y+oMTPf8WqACWd8=
`protect end_protected