<<<<<<< HEAD:flexrio_deps/PkgInchwormWrapper.vhd
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2688 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
eqFSpb+CvMuY5DmKJBrN+h/GgGEjTlt8UIqe+HyUAP4Q/D/UpHx0jBpEd6VKbPLZ
cqQh9ZSJzdjyXOTSWLBPWv2nkTnWus9+mlt4qgy1p8fg9rKYKIOLVveCIsVsKTA6
f7RWyaTGa4G35WbQmfkDzgeiUw60aoR8sj67VwEeGQ4ODbsRHusE9NZO1cPjulQv
1NnWKIr6asbUk3nWHI1Zw8XlLFJMy4RC7YdoK3nmdcFZZvgA++ZGtwD9mz2pmPZC
O3PAvBBJaJ0jzNe9YVEHfm8JnbKLYzdiX3eGKEjmNSwOFgRibrK4HznrMXR+TBsv
skB8YAr/LOCnXauu+wUtytsOj5M/kowsvW3qGCmY3NvNgQ7oAo6rMEE/HTenz3k2
9Z5AYzMA58/NphcDYsIZRff/YkZNCkriim7Z3q9M+h3Y/rIqeBaUwnYhVVvZvX8p
DpOhej50dxo/mtGjHE+467GiA4b45jtCxjGI2xDXRSUxVronBrvFfBQRxmmh1vEx
2HXkQvJEWdVrZdo3AsK3qW4qQqYUphisdhquf7oVNy9dKa1RArqp/ighJFsmS95O
KSazhMXbSGL56fA/4Fb/fHtektOmkximH39SPmgooxQqpZs5iTpIIxhnzOmSEY5f
mQdW5I5Dx4xKr43sdFU1NDOzZ6tfz8b4v2qTNuc1us9Zt6UnCBez6Z9MBQlTzozq
k4bzwW13zpgXl1E7YO+n3ppWtBHyvIz70k32K8uflcl48MbDOBKXSeckEe8T5zws
jvrxWM29eIbWm4bGDb4Vxa44AaV0bUKO3USnjeulhk5jl7uCe5kwQLAI5CQoxVny
vzK3e2RIk0iY1I6sdkms+cDrdY45zPlUIU30f90JQsmnSbon3SitqxCrgLADQok4
PvBuyN2IXld+BMlBoims23gC165KnkFkbhcWt2VxTlfSKOpMB0lO1adQwj/fbRgI
eibWhrjL4L9bYWbQWrXnHm/l0kl/+K54egLanruvAqfDOpxvLcnVr8nrYL+rwWMr
ELZ4cQJUqEhMFwH5/ytWBl/4haPIF+TxWDm7S3hhzdgwlWy4/TuFUp0C9tR5mJ6C
zF92+aYp0LwkQZsEnUPJJf5ibH8Qug0bwFQ6uTJyFDSYrSijvfTkEb2NRkmsrluT
rIWxE9dhmh+2xJw27K6QY0menwkhsMbRJ7EUwdcO6OB5qRGrVmf2/D5NdPKoBcbS
UpLYGr6nVmR2Av7ct8K9cs4QREdnFahLDf4t2b4esAZVZFfa66OBbIRuzQeqkyAy
yWcS9XX0wWMm5X3ZLuIqseiY8Voot70s+eK9Lxf65N24B1O0rvVqGJJmk0+MPJMy
jkMqE2s6MS90ZSM1cWq8O21Sb+PoOFi4/+oFFKG6GEFMrQkYKSEpQqR2oHKG6+Em
NKridFcXJXDaUTEy8oLzCqxvr4FFuuCE3hXNZ3S61uE6c6CrajEyl7U1kF8BFfVZ
47EqDnCQweWYe4aHWKNPYzJPCUquBx684G8XyccsA/1ZhlMF1+lQsMwAm2tOjELM
f38tme891qFEPR3wh0117KNCH4dASvp8he/J5bq1JBS2/b/ndBL1itmA2IGZDB8J
U7keEQ3imyYyhD8KKbEVXtgj2Lr6N5seDMyE5pLo/5DZd4MEXEbdnVNQ2us38LeC
lDdSLXC/fawKGZORNtqxDfDt68K98iwpeOi4o7/1T+ZrCl2frAtFnSacMBLcg4J/
7F93kUy22yww8UK2w2ejF4GK51LlnhD1qKtSHI381E3wYMvG99MkTRky2eRxWRGU
3mbruDuF5iRUeyp/Usbm74Cm7t3vZp8KBZUwtPDy243q/DsfGnUZK0NXuddPaSTG
5OwnG8NLV9TZt9laH6gYfp2iWnr9HpZDubxFIQT4RL738PUQGqxwP5mxwjz5aw/h
Qo0+gh9A4Aan9FlEVFsBcEqTW3jFZDvElxgNS6uqgciz0hzVUGfpr44udQDZ3pA4
agrNilxEaet+l2z0X54/2ZuuYxp9m217MTLns4J7Ju3hUiD0WUWA6HONFJyAJiWq
utWQc4lEmYmUsTrkEeFmos0N4pyVpcjH8nXmO6qXrn1szQnOfi8MhL/3R/QnSPOk
ZQrpejqoMWChnDh0b6KbW/C79wB8ST1cm/cZdB9Q3zmtgcDH5wwFiLSDU++k3KmI
uAHFhAaxYZgA9dk558VrnA802fWY1BTJkWfP6WVAJwXxR6mLRllTw4np7TOEWKkV
/cwPvelYwD5W9uILsmRPO03Jm5kydTUNWUMelWNgN+BUtQ8fgMGW36VC5j5V4e4F
0ekxHdXAjtLKEkD7F8nE5i+gRaUwwxb4CXi7QXlfDFQWW9DLvURgYsgEQ6b4hw8u
+Tlo3rsS0N763Xdpy805+jiOY5OeG2G+hNYhcqxLZR/Qk6hcCRyvBfNArN8tSDf3
B5riQSuSNmrlCp4zIDHdfbOKC7570NsOLKdwG+2REQavH7POpde9bLf/gNAoTT9H
eHOK1U0ToSvv6uOxRkVKTFhLo+u9nhGS5a8QbcA8rO3whOfkBkmo8jj3eFU90sKF
Y4iS1srWg1WEfvpTbV3ws2d6KuZfLTh/WPM49EDuTW4eJmQ9MqqsjW2VgfC+Euz4
r3luBh3i6LojvZyzqUgu64PIyMT4NPsSTbTN6g6zpPJmU1KPmI3PqHX4sSFUnNTZ
yrGoGeTVx5OJDjoSQ2+8TKLQ4SIXgBrSmc0MoesYymE/gIFiOmd5qfjoHYK9MJn2
uZm5HF41BCRFa2dW3m4T0etmfRvSgQIDqkQ8WMq+paXD7JutDVocDQ66u2bQ6NfR
ClU2ZAFqYa25HBF7av7ZxV6YO/8TabC8tbvg/ftiyr1Z6MdKGKjte3TmIoYsrQmg
ylQK3/ZtCsb5mZwaUN2BOuho6zVOTbcUhj6vcnORomIaV84mXxoI3c2wW0MTXr4S
nqgJvezrMuR7X70V6f189bZmIzl7ZhNjTvYwvMYpafxhGVSyqL6BtV8Sh39paHkC
B4emAuzY5NSvHA+brr497CZ0m1bVN/rPJo8RBNyDMX4wu4UzfNLwIrLeQZKX5ajq
2DR62dpo746EKQ2H1OW5pczhSWCAskn06c7OG8CKoG63tDzKvrfajIDofL4wtcSk
zZN3BHwMkDG5b2fQbblEVX3Qtr2KGb6ecMtHNgtllE5dKB4GoHawK3S43diXZC9a
dX0PL/pTXuaFNQRchztzC4Db1rjeegtdG7GVGM+jjcFC0T3JC/Nmc1rEGOoz26tz
qLuTh5cRZxm83uYp1vNlsHy5GWDkZ8zWw8UV+8zyMl0LJ1JQe53cRu/SmsHAXumW
tqzCy58uWvY8TyoBQ19DQEsaVeQWVabFrNdqjGD8NBT1+q8/EGy/vjJNop3VDZbG
O+rwWze0uT6YTvUDpfGhrkOUiST77RgfePAcM/vIBGcUa19Mq47ERBNAGuxYKr0V
=======
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2688 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
9oM3kKfrWu/c6xK6HsCF4eyCFdVr5Uy5aj7+c6r+CWmPcNT8O5TIDpxiODNEez5c
kzLLqCqBROpfptjXFvo5hEcitAYfbLFgBNpCZTF0QF3Y8id/IW7uGOi1x0k2cORZ
/zKy2/rZszESbG2RodCYfM+ZksFBlHBSW5OEq0MipIFZOa00R36v8CRoUOoMOT5A
U9Zfth3cXgsqp0ecJk74GEJxq3XdOQCvqHc3rMYIrMxDoTaL9C5P3QHnc/t2RMAd
yx+y4rZazeA0HHzR1NLULzV4ieZZstbTvDetSvAwdXh78bGuiJcWc3ym9BPiC+vM
d7lg26pEI+spB3SPyGruJcFcWHTY9HhrlrmtSOWSqLnYv4FMSL+SYXUKHIi8hvQy
+CuE/ezZqH95aTt9XXG7L0ZFy3JMGVfZ0fgVc8eSIQTcuXhEIkUtRDizuV97VPFd
IJM/HPubO2yMpJNfix9nTbdyJW5MH/HMvwrUv8Ry+9eq1IoGSFUVHHVMmfmYKrIH
rlnzW5Ksb8YqJ7JxnZSICqhj8fAUzCrijhAP4IOpeRbpDVvMc/slAsX4sveHKkdc
gH0kHT05ftVyzKCgYvjuUIm0n0c0M1TpBSpI0OX+vGHsiC9JB47NIntpRIdK+kx1
PdlhGJ+2ovWVZQ2QrLlNd+falXg+FyGvQJdQra9dx7UvqMzpW/HjzsFLc9S1SLQ8
42j3WZlrvdcUy25yghXTRSUmqhWknnVU5gfE0zQXxjXIklyPe4lP/wJBTzi9HC6N
CnTBO1G+nvLLfXs2JEeVfTsoydlgYWCF5A1vu80sCQ0kzduT+pPtDDOX79K3aIHZ
0R5LA1gP7OaYS1oIWVUFtZA9Su4K+0eE7ncwcocKOBhMmGxEAhDR27ZCFDPn6K80
yg53bJjD1tRR5JUrkmzkJ+HlKFj9cgWCOj8QFAqUwYPgg2XRQtn1dH+yN1FNyKe3
Gi+jDIwmEPcjk8JO8XBs6WbOxsMOXkDy95qp8oY7BJm/HUdYTFcT7UOhvGQGAaZb
mwDBivNQ8L+Q8I9GvI4XT7vZ2iEc1ftzhPsZnvDJGN9hjgDqn917pGfSz9+ggjsC
wuq8msi+zio2GSkz7D82hgw5+8DQpcwEKtiOtHlEs2bcELy41ULbrGMP4tE9WnWk
SkWYHWPcnG3e19GM7nJokIRtdeWUAJy8M/oOkGhWEgP1jMGb1qudFmVIJXKr46kO
hDnUX15fPB/TLnHH+FbQ8pe6TZzhDcf6lysLEq478bcAuErXBqKEPRwy+HJbgOLP
D9yzh1zWPZMXAgMa9w8XF71p3PhEGErll095YQ3KdnAVHJdv4I7Ed4HUh3bGpMjg
7OoIgH6RRSJevwzSz1SB4mca0VxnVEq54N9744oLdTs3h5lhWmpJl78zbqw5fLHg
npo2RvCTitcH9lyYZs/Lt5ygLCbIKWKnqqkpkNSsbqL8iB9Iv+te8ZZuWlAPJ7q+
pf1YYFIURI66pQ881IDNUf3C3RFDWennm+JOzol47Gb+2O6J7pJ8j2MqPL27iZMB
6dXRgxT1Mfi/UAtv5XCJOtyS6x+98MCJ99E09XM/4jMduRnyyhK15Kpu9a8tmAzn
Gc73IGqgKBuW9Voau87/Vo5FIbELaAIQnCQxjW6QGuCYKaV58wiQrTrvA9E+5S2t
vsb/0NXmN3ee0w/8AsgbTJkAeXDZYOzzjorQEFSeMLv51tGWpCK0BZDs1IljQ3It
NSUNCCnLZHYEssvrg0o1Y2W66uTiQy3Y50YbkpHtBFEPPwZJEisr27mudgC6UMHe
OfOqciG6viOV6lsNakBjENFahptLq10O+p/5z/5m2SeK7CWQNvviYmajNcKeSNZn
7nnvD0uk4o9c5vCFI4Sr3gHCpdm0n+hLeZmgK42RslTGy/UUS7p5jh6b34saa78n
KaAmydnZh+UsLHPnNmKWj6gFWUTIuBXoeaDPfqAXFM8tFeeq/E8BNbeVagcRrcQp
yBGqAfmXXh7HAQDvkbZI5PDZjBjD+mV8KIWowTKBkPFQuSuUkTo5zkKLIfMEldV5
P1zQiKzb/E30Ur0ufLwpr7uvV42ktEsgmNpVjauJZ0wSIjmd114CsdqcP+t5UTyx
7gFB1z4kfr/4RFg5y548dl5awzSMUfuqcc9gKDX9rsXqI8ZHNhHlR9QMDZSGiC8k
5495j8FTVk+Mdkm6KOcW98hfvmPSqslkk4vPKmTTG+/V5WCnScxoV+pf8EHC0Azf
75u3cy2uR+M51N5pH1IG0RUOrisf8kzTKExSIhgp8K65jmcthl9Iro8JScIvW/oF
lAh7zn5mccIvJvxZnhYnnXkUnf/PCc7wUpnN45tucEC5SVwSGQ5RMpjijUjqlctU
naPzz8vW9ullupLHIUJIAu/U4T8UR2YdobdMt7ZnwYUdyCGt0K2iXtUFx9rExs8u
ZJMEMWJHM25EfCGpAXexScMy+zhsGXPommi7os7iVFiV16cpwpfiQZZ0um7aLAgd
RRdOVXPF3qTI8DmTgCYIZHHW/oL+UWkwK/cyLUuj+zRQ9AJ6zDye4gWUqYZ9JAK0
vWNNubVSweDLTjp8HTK47b022e1heU/Rg8APrx9SztxSTM1EBiz6gni1SJfEwFeJ
Q3L5Eq0+WsOZW7LAPnrmMzk4qUWVfiM8QnrubG2nY8tYqeQ4vBvrlJ6H/9aJ4KTK
nRwONfbHou8EQ1DCjR1XHj5+u6uXHHGD3d5OFGRud7eqtUm7nyIqObtMwBWGYZJQ
En09QUtEhGvSTNHGMfkvPc+ZFJvwVjle5nAIQNgMYIluuQ0kTpIh/Rc/HiYFLufv
k4ZS+o9/To/L4PV86L7WBKIjZ+RHd8c9z5xOPGl9kxzLeQbDm02HR+yknxq7pO35
O39TYZSYq9S9j4xpwGK+6um6wi/pAMzlpB9zEIlcvDL58Y7/YvRwBkBFo8S28Pip
gW65Q0ryFPHPrnP5VPvvs3OeM31xwDeW6pmQpc5VOt4po4+wvTSuJb70nXzZdT//
1GCQGdWyc9j53AJPsfXTtfxFURPE4xuEyDOQyp6ygG7wtvf3zeG9lnQUCjpY/DmB
daG8QNI5sUqu4+YCTkjsreSXKE1UZjo0XaShsVxpetsRi9cy7aeh21REPbx6hDfz
g0bB+g5wsEEQVITr1wfQxR7/wfERQywma28sp3NjXZbXb8xJJvAqWQMKgvbTVw/4
IsKaBKQfEIEb2L2FL5597vUi9Yo7UxnJGO2mVeMQL3C92XwKK+QlZwJno/Vo0Oqp
sX3mhaLbAQvDzmgcpwvmRcTRP7wAAKc/mrZ/f8BakxsuA+S3D5n0Xm0IsF/AyHRi
67y9WLmFvciyGYEH+shHxV7NzoqvcJWV7VWzfnSPgnPtkACqAjg96TVXZC+L9yT1
IuRXOOMBFP8BYnyOefLqWCpwZhML6Kx5ZSU3NR93y8fgBYMLFs2qAtjGOpc3rwUo
>>>>>>> 426889eb8ce467b9c9a9f74dd4af433c5046285c:deps/flexrio_deps/PkgInchwormWrapper.vhd
`protect end_protected