`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10128 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
FPPR7ws3fN+RQyk1V5tkgDRlfXOeaLZ4kJY2DiCnJMipPRt1uzPT699R+P2KsTBk
eQzhVIdevoAV9JdTopIMhE393Uw/ZDtqH8wWKZ+e2QUyN5N0RnHno6oaByV5uNCS
5EcEuviIvTj3wEr0/bA5Q8AcdWzjUUigno2wKCFze5rfc+lzkiGznGCynY92KgvK
9aB3I0ElkqounKP1JqvOQ8NQWwkSyyU7dQdYb2MSATWarMGhLFH2GZvzOQORIwwH
7hq/BLO0WPIZLxd/VxPxegow/LJlDKImOi2Ik0vij8xxaWvYZ6cWPjsyys4j+odO
zKoS1ec2EFw01Ivr2j6hhvBuyNurNvZdC4uzimD/1b6jbk7N5Ey+RghvvNFOk3/R
S3GiqHzf8dve6dIZNb7k9AbzVjRPeHj7r+4iJ5dFOnCCvFByJToXYLVQI1ZfQWmx
aokIdOQj3dr2XA+nKWfHoDqnWnmT4xlTsQAkpntOMC9pjt4977tYGPhy1T+VmG/c
OykxqQ7pOzuqGDDBShupIgMbDxQotfhh+wwkLolYoWNHr4lx01gDKjro8VPhdI5s
YVjJci20UmPJYTWml9sxIJbFv1aYr03Xj56CjKWxAYZhoeYRKg2oZEur+XVqKwMN
IhsH94PS9DQQnCZ20FvRgUFR24OcHy0UUie+HQgB6GI8n7z3ES3LJs4NzQqoH+J0
/WCR+0+xx5DvyNAJ41HQtbm3uWzc8NVEJk4RMJkL9mJl2fjplSMclwhC4gnFi3cE
Qgo8CjCySjF7q0jl/ukR7pEY91Iy9OVxomeNeDO6l5pkgZhJ5fGbwYd1QjfrWg79
NrgrWjeJSg6+wk5z+TmXPasMb8lXxCe2rMmETRLVqvwFSqWAuTT0xhvEnv+yREdg
lwhA4Uc8WyJzf1/FJkVTbn9/X12lz28QoFOpSXOwce8f/HiUBdA7JP2zcgjii6XH
QX3j+QDo4ayurT/fq0n3MBj701vqX1l2Z+XDhRJIvWHYzTW7Op2ASSxh1G6oIemt
n60a0Njol/gw3YsHIDhgj0wV3LqChY4ZI3gIM7NJuK911EFXPrLVDKoF334q+vex
yX6O/6FzpaECRJVLJaFafd9W9bBYJ4UW5d5tETRW0OaXhC3YUMW1C/XAMDod4XEp
XCX8gh28KpayircVVfls4nTBGa+cpgbLnmPEVTrN7XKnlTOLLosGOuYwnjIaiHcW
JTJ9kSJqNt+KVn5qVECM9XPNrnQr/MKUpcWKDFP+ZlbL/P+rOgnV8SbYqxq+z0o4
2M1TWyB+dZ6U29W7xWaCzDDdacnhcu+GIGgijb9KtBrlZajNjNxiHqZvF1g+E7uc
vrW2NaNi2JMZFmfgBaKsGE+ktfUIUQx0lCP6odCoIw8mnW7Nm5MNG2dBJu8I3mAQ
ItMFYnUbtrPjRPvB6smQ9CKYT1gqvtzCX89latCD4JAUzK03nYC//GQHIz4jTqOd
KViZJ5yr65pV6NTBI768NCqYAle1Nh8egLUZjVO0R+mznzd10Hh3AUWj3uHPQkwT
b7a7a8LqhwT7UxILQ/rC/4cbeZz46qvqszngyU01KmP3yO/kbcVTYdYvHVkEIXTC
VPYn6vbOatM4UbE+dCg4HaiTFCfFDPnVQYn2dwllxuoVddPH1XzgHCN6Y0ReKFM0
XDgOrCFkn7Y5mKstX19c5T0rGsepIOEK4fIvGKtKgWGWMkLrrGM1b2YOj/kXmdjW
1Yaz+8GZ8a5NVAdB7CN7/ECxc1FFtDZp7l3oAFqhpky6M9L5uvcD+KTPG4qRdAvt
2ouDni4H0OvkU4v3g4PCZWxqrTu2XQqo+MCZvycOe5lGoRrLHk/uff1yoc9DBT6D
chrp1GowkdNgKQUI+Uyk+rjR+4Y/Fcj4xtG0nldumCfcc6kdDam8gGhURWyNK872
u8pkGx471ahcM+Nt4n7Fxna8SOV1J3T3HIIJLiMBjKvRESdOG3UOvbvsvYI1KAI1
ZEM9fkhERH8oiA5ruq12iisSggcur4B4EBPKtK+KAyCkQ0tkDi4pHgje247ef0WL
einJz6vfReiGEM+jrINmZ6bWKocrz8jtP6jnkPmwcvw+X0GAZ599JuVnEYT43KpJ
stn+pHnaXGmE1/0lbe4WOt0CmG4HSCqAtgD1mRyUAg/Kt5ZBNMWI8actowrTIuLr
9Cp5/tshxx17OqXH2V9GZjsTGe1VOArUn4BhxyGuy3c3HwoWYMxCsMF5ocOG2RbB
7gYjfwcLWfaumr+mwrAxEsO8IoTl44Ghe6O8hbEbUhv2JTlW3iiJ0TomV4OvbEPn
v2gHARoHgNXvjiiViqulxEZS3RUoggICpK84Bu+6wbfqBLd7oKOfXrXV4P5JMgEs
pMk7WZH5xbC7drMS+GX2C7peUllDZIz8oCEjGfyZ8mhAubok8Z1C5wqrcr2mim2A
QuWyATSQSPDE1Aw5zEiHbAZBNIoYFWKJ2JNGTRLKNpanVPUqxwJzprPvROk/McyG
VHNBmFfieyfeB1Z1LLSHtkZEmAHZuL140RhIHknwaRkCc867LucEwnLqigxNXK/E
VEQM8/cfdiVwmdE9brglYrHa45nuvG1+IhOuInHGewn+qOLEsIZ47/7o/Hgf+DNS
V/6lcAhFxB9uMLqh4iWVSZtRH+tCukq2A23BiYTc2Va3SMqWrBcTEIZ6BOsOaxCJ
bUNdJqbhUoVn49+l+aJzLXkF6bzJI6FuWpgorKEZaVc2vlzJZMOilga3inOmCwO2
S//a/qSnMI5gsFAPisabMxmLC4BmOzEcNQQ1YrwWkLJKy63xwN+ZLkz4mnWP6p1e
JtLxIfRv1i4zbDd0Or+Z2sVxCnRa4UZE+TZq7ZmwTmSAMCJBu7seP2kQB9+t3m2q
c36ZFGjr0rs33aH4pwMla46Q+kjHbFuMvAfOECeZNUyxG6Xoa3R+iri0nRioRzkv
QE8J8AV82u/z3inuJN4NIB1xhei0385LYomg7B7NNe77H3kMz0+oEsUynyJF3puR
HwcDuzxaAtR0W2l9/jsDmhqliOaUOVUo9QvuvQijbiNvO7JlanfdygGM7VuvRTM0
KVOCSe+qY+mxjXNztqajPAE2hdkNKdwNCs/77lfTSLfhoKAD5xZqiQFvhlv7bD7i
ht8e1YfJg3vC/+gxMzwrhIoOf0me0epXIsc4bOfQXfNr0/HpTT1PILxaregGhhlY
rcrxTpMtTHK9VBmVIMLKQgm/eI1ZxW/Zuyf1XReSgFROYIl0ts6qX+wfnt6e7msG
6KxfGgzYCHgB5KhRqHErPPrC0KMdj9nk7edTGCoVxIxOKdtD9jXjWAPmw10OjShD
06jo24Jbs4nhEppE44F4yfFw2yoshuKzgT4OnviIiyDZ/kSXXHHFq6ymkHsBA7/9
NDocoVjLBS6GAxL8FBXYvP7bQa3yO2SI048yZ1p0wpUM/UDnKbrvAIgqBIOOKwPu
xzda0i4Y6ezDbD/oDt0cQEsRC4flYsRYCGUq8mFlh4UmHhFnAFexQYwYGpOS8Vml
E3b9gChhueulmLjQ/09p+T4tK+u7k8KGeFD/Z//XVAMaT6lIp/XuGY4Q9LrmCYa3
utSrG2fcYnNL+r0uRK7/yyZPxk/UWbln1Xwj7BBQ3milrzn633wZQ74ab4gWoKnD
JjaSTEDzioufs7hRRHIn6qtQ6p7JQHkCdqDdeXo9KCQpTplw8mxC54fFXzC4eBVG
zAPTb+sSWulISW8SCaAI0C70KpjavGiX9cz4CjuE4v7OJ2Bl5i/AJ5BVmUForl+M
n5XDgUoMxc7gCU6/9QY55VJP8tRsxg0ZyLGVsL/kF2mf7vsxQpCi2XHAvy0ar1eA
qxBzgiKtYZFwrpIfkwWvnFhu7vmftrpV2VoKX2pPC1Pj2LueBHjpGDI7GCJRoFoC
WAcoWJ/BPExmS+36H5ldhjXpSVEiI/M5ZbINa0Z9ZndhGYieoTlZwGcbWAIlglri
XGQY2lxnsCG7AIiRXAVh5H1fdG0+5H2cENBxtmLzon5qNkSElX2zsLfnVpS/kgax
LlaGQPIes46JFPHBA9TLAEo+zt1csvrwKZVWJi04pRqdT66UBirOVYXoCA8mTotl
QXcByCNvUpeB1EaojaVlC0hSQdlWBeRYe3iEctpTtmYbCkMNcNf81mSQ4NozROfg
PcN4qtPb0I+fhvajh3cvZC5ZEhgdosXKgZS6d14hgvlWyMMKuNbV2OZg6DwWRfJK
dsK2hlmxXTEp5tDHAuLRpA0l2PHvNw01mlb4b+pY8MrQaKthd3qQ9bt/x7MlhPP2
iGajj6u3O25qdY1KD3f/oHmvJlETO3TZI+JWUpO9zTY+QJ1AM5tKi7otSdnF/FO9
ywzv+0O3z/cxdp8Z8P2peaacQgxM9YQtmnCYkeWkAetDgcQrVRNw51QiqfpFcIkc
j1O/aDciC5ub4U3Fs6AT2hHSPJpNojctMWAAxtk2Zcfoh/tv3uud+F/RNlg6YPBU
ePSBHcqroGTi0LuO8y9TTE5aaHAv/PqxjuK+Z1p3KkLUxBp+Y54OF6w83c3Qv0CQ
/8AYQfvmT2NBC+F4Z2XidaZzY7rtCkOdPmKZZrTNgB5E82e/CCfnj95JQv3LEgQF
15vKTfxWUhPoQv+sJHJ4BRafbrJ+hjk1b5hTxkMN493fSYRgl1eYvQ76xV3sqF3X
xTCwQcCRELZpRwoE9+6UaZF2eKJEJwCHFAliDrKuqUiWREL0p/MGRdrXJbvakLng
WGA2q1nbYi3qQRg4C0QhlfHOcKmOgbiYX4qqP1EVDazP3XgwJquw9MnT/NDQYdeG
T2c7m8w9sUf0cDWMrZ2PZOITRiRSOL6BAXVH3F+Df8H/YliMSfiIktpdAACN/CJm
J8EsdcZkDqCz71smQXBqVzEbGWsr9IxsWLgL9EhwBqRzgQPgEE6IOsvCOq8RLdCG
Rozpe3DoHffGiBVJ4ZaMOqROEZX2JeyePP3SYrUpAwDEi4weqf5DIzeiDSKzqHcR
JxreZB3BQnRrNLnAcLThXyXY5rvXl85qZER3qC9MQiFMHsLY7OtE2VZLYXaa+o4N
pPP5M04HEtskJmKEx+Titc1q5Zqd7YshNT+fiTAX42+/n+Rsvom1Th3r28vD8ONJ
hr8rjxZHQwILvuGZhPX4G33uFlDpPLIm/d82zQBRdTZpysf9vXoTan/rutXACKXL
hUYgKJyW3hSFviTLEwEwbi2oeANojxBfKa2Y61DOTpulYJ+1joMBSH1+W0EnxwYY
yHjjkt5ChyFBnf8BNVRIoFJCRFbZtkt1R59VC5LHMf6DmRMn/CQSLBRM8PDi0mGB
hkUQdA0M2zq1JxH87u7jcq32pz7+oNzxvtvc6d1PKXpPLQnG/klAbOH4T7fHvUPa
GszLAaL9ooQKowVd9aECN5oQMXfzYR4vtrlIdXlMT6UtqSOgu1/Vzz+madPhO5Y1
aQqEB8Jb+qwfXn+r6c2MttHwfzNvxIW6lgnbLYSUnftNrqr58nKWaLNUHQzA67xS
kWtJlrOr6VekhwCqrFixPHY/V/7Nnrh+7ZQ0ltXpzBrYF8VLjqgCvlVduLFjwgPz
t+4O7WTFhWLNt0ebG82Sgt69yU7+NseH8VcespN8heUQzsHFdkgD5+VZv1W8qbU6
0iljbB1osCLNNxZgR32Gm/xXSJyTcMbPg951SSadtuDKQcmm9iLldBlzl10EVLqE
/ptys/Ao3GCWw3PmOuK5n3chnjQpsR0UIaJCEOwM6OYaSSnq4UuCm7wFQpF2bMAa
O93DuAyvZPeACD56MVBgISsh5/1l6m09MZOm27+OuxWtb0Q1tTWbZBIXLsLAH/2/
CrhUgg4t2R+6WM6jpqvw5gRw3Q1ScRq4Vqt8XFQXImJJWTgidQCwtgv6KmOFPVTH
+ETIyIOooMfqjXpx8rCZMEBDHLb28VaxdXQbEjPdaijV/HLClznZ7B5EyU8UTt+7
XzycYcrToVIZi8man5+AI/yxkogD4AJXa9ZPzoe8G5eh3+g/58EXo2pxkpVQYPiH
pyUl9ZFwOiqlcb/Dov/+V5Xw9HJaDBvYufCHFe6jzxtGPvw/CARN3hZ8yc6bQW06
xztulIBzJSO1U4n6hJKcYXwrXOD6+JZoMYKT+eZDx9Y9vZyk7VMSnKamZ+sGerjS
Wo3s0OGY3tfPfg+uv+ErQp2jpTE2h0tcorq+G7VIe1LhrwsieS/Ftx5WxiY29A14
HIpkET6pOdFEiycLXrwilW10Itsr8zCud/RDJKlYLzWfVNLf5N12eph8T4zh3pOU
AMKMbbt7hSK7gctTKdSLdklErV+mJJ2OOSVQRLYgTxJgUcgHSurIct1CpQIwMUVv
TVGY6w+457zXj0nxw8XgcZ5gqeZ8EBsTM9WI0/z9Izt0C1ouJqXei2oOfah7vXgP
rK1vvZ7ghqNP103vfNHCNXDbLmUNNVQ9nXmD/1NiVZFkmISBepH/AB7XPJyXnMqA
rU1wtLNzUi3ARYR0RC6pGkNP6bQj2DdPBwClxsxGbKfccQ1jZK3nQLz+E71mlZ5u
F5NCQJ8+s+D1ZH63DVvnTa3DSVrnn7pOodX+B1we6Ru7coXHu5CPo87IRIkPceBH
Q4kvFjmWYfGP6GPWPCu6zDoLxGUfrgCpPQ+SEushpuARIMDLK9IwQxfgfPF87Ybd
gchza7wVJJEnH89UGqtyxfd3JErZNVTt8wEaGXapHyenjzl2heXJVwM6uEq3L7th
hwqkCeZQjx+25v7HbJKQXw8P1e2moRkzxsS/ixeChAi7I93Bd+kxbRx5/K6aUI41
lxOUl8AwPdMF+jTop+6CjZTVamzyFIl97vAM0go4RqSBn5vFrjvnL4AB59fqmj2Z
Y60exBDubT26NVWMMy4Zz+au68yWUauH9Av3UCrUkeSw5beupzNCjsBiqcxqa8Zg
ZmozG/XejAGTFiW61U+IM2ulLSOO4fStka9lkvnQ3SK3jgnN6sptaWi7nZp7vsnd
cXdWRCHIkB3dEhNhmQ+qW6+/zyicbfyDAeb4zMvdm0l8sdFpe+pofqgvDGWygYyW
xA3iwvFtOs64sQbaeYQT6s5nrWX1twmIZPsrBvPAvA3QkePa0r/JEt5RoZO8dmt6
7t5xZVGErVSRKQc+zci5bv3aTldvbhGJUTT6c+zh73Kk/l2+nZEfayWAOhcVfhdf
aTmHb+jwEfN5eNaXcYPo13Onb4Vz2ofOiz9DqYCCPkBEcLLeu1geNWfF0W83E5aK
c4T7EDCkIJN7WoqJz/UOT+Kd6EPeRdNX6PffQt3xyJAj0R2J/xt4h8WIocfbEzq8
XmablCPo1XCbWl2NTbBcuM+1yL4KXgBxmvhufcEq8x2h3Y5as6++n06rEl1vDBia
D0EDEY8pD6y6/h5hZiPrh8lI10doE74P1QC2glWAFdwPIFFT61T2aUHZOmx8QxJR
sqQWNGqTGL+FcArLnjoPxIJxxb0+OC0nWlf+j9ceJEdL6hdkNEnnXDNzboT67lii
d6kBJEV6o3ZfYGg2eXKr4U6q1vBhkFeIJznybEOThXpCjhVd/Z4UDm9yLa35lsqM
9hl0i6BFZ8Rw4w5kE48hK4I9qqcWhfUI0KauP1kcZu/D5uaZm3skqfugGweTu2Cw
C5bpOEH+Odlg2k89uMwBkpyleecxAAOsyQ8r1RBuAmMvOoXd5buK9JEbaNmxHtDe
tIv5tydLdX+O7q9kewH8CCXyfIn1KDONshi5LVRRMdXLlzojiR7AkN8CppfU4ucD
VL9rU9LaPlTQYZwDD0qFUWktkhnDIccz1h1SvDobrKDJxOxquwP37Ax9v5Q1DDPq
olCde9YFsh+g0GfvIDQD/DVD1KLmjzWZo2MfN8NH5m1zjbIXWCdwrA9CZllbM8Gn
hwfSccpODEz2sRgdCGAxEJixPjwhQXzrCVYyFxWoQ+khLPXYoIWjwlbdIfNydj4p
EzZ86bFhwqY6poZt7/dAT27Xu8I6/Qp0aiK41B5YPxraCt/4faak9I3BRQJElREp
guQNyV5f4c50QoEiKf9gbvsUKQ9E+w3itW5wl0KEutidczNSBu3qv7Iea90BkypQ
eVR+uksvNpjIdXMt+YbvkVdbXxwYb9hEibNDvMhXZknHtHMBJtv7N3bLRBSjC5nD
WdDQq4ziEUJrSZhTIOZU4EFHFgxxnNTWDISMb6gRsjE79lRN73yfmd/ILUpoSAmW
1Vz7rPVYZoWjTAhBnTvD3aqGJSV80owfgZDMrGSKW5WtVckVPWwFQHve69TazdFJ
dbxLJwkJDIwPZe7pyjM+Z29s89uveNMKo5pcDFx9mBN/kacQ77WgKOCd8eCaQocm
kR9xnNbEhd8OEpBDLVRsf0NYZNc9Sg4FIPZCkYb8ST+HIG18aDy12yw2tOpTisFG
XBZ9dZHE8KlLg6FXpmJ3K2IvrBeNPNqOZT+VKIi+UxiGghyFyxD2MSP226inyKI5
83Iv+LB++BWlfGp93bQxkSTgYSuDaFDThfGWz3On4CXXLteJI6ylEHqV77NxuVIz
umkhQ525zX2B5QsilLogVheBdQ6GM1Ci3il+bnpMRGQDvGKlCcExo0xAYSWKS10T
NNygcLAiJMGw9MKRt+HCCBmeZ1zKMBOOlBqIUizFnksJVTHHh7iLBkyZAu075yvd
gqBXOYFX7l974veCIhDXN6S77ROB6t7dNUawNbwSP012a2ByAlh7ox5T77Hz6le5
uhtFVLBBu3bpYB5/6uUixu6wR4R9CxFxmJbsbuae7307uuOzt1bd3vKWcWYelYYS
RicbIHOLCrVnlw+eYzR+igQrRWvJGk/A8tdjuinSgx09261nyTmt1ddGu9bia2Dy
QjByOnhFYE9FJhtuyAfT9rehnNeUhR7SZvGwRxYlNWtDVfor7w5ccNa36GjgrBGC
t/WDnukXb05Ccpwtc8SZ6dsk/hKaxZomw6U/CwyQfcAlWoBQis6UtmmnspgWzWhs
cAZUio/TM6uAGEU3e24U3A51WqLV6m0KfTPVXUTsnf9TUR713MhKqTVcExhjft/1
A0j9r8W33p/kFqb0Ql6jdayD0wWshH6rd6WOZJC4CsR0A+ajYY/YzI02SC0QQfdH
/klXwZG9IsYvYq+NULPW2Ph7aJ+Dc4UOpynsa2QovaJwnIsBrKBOH+K4WxH0mwpF
Aj7RcIsSNYr+iqMhy+TZfx0F0+Y0Glw+apqHglR+B+s1Fv1CwIEwbjkJVEL2m7AY
34P1ELYmp80LkTNCvTV7QXdigREL9G3KgbJtVOpfaFetQQrLTUuss5ireT1DoXkY
qZQ5abGslButLDYRFr8vsjwk3c4Vp5OXiigDc7Mmkkxeg0FkfXcSWzJqDBLrxkb9
RNYFM7EYtlMJpGsHKa4fGVzv8AtpNrAZfFrhYloQtHBCmeSXwuqOZBvGrvc0RjDb
l+OQnn4Jw14gpRn0psgpcrxLcRLLkOuonpGAEpE68nBN5JY+gkfVK3xfpj3A75VY
8BA3DoGOuJv3xlvGREF9tfhvifa6B6+0sETZO3ktipAMCWTc7HUIfOTQNn4hwJMn
COTGOKKp7iya/rZaS7bI5YwJUQpLPkNkwwxUMgVeLRfeee6pur4g2q16hO5TWEhH
87ZXzCuxJE2J1L36A+zdctaZxtYjf82uioHekYm+3OUlxwHr7LnZUWX+2YgsokcH
/kNIGM+qdOMeFwyAy/uNSSl2i2n+QDf+WYAZTD10C0YegcuPqzUjh6jqjRFtj7HF
jk7pIsUgZ2jREmD0QNeQVFhKEHcUPwoLrtVK6kyTyAbE/xeh2R+4SS7JlNx7SdiZ
LEaOltM3ByiXBItQ04CuktTjrOoAWsX0Qg177gvxEXoFjqnBusWOQimlJaJwE1vn
YsM9d2AOk22Sn5pyNHASqgRzrHqAOo1b5kJvTS5j8yYdwFa9+cd7QhaUQhkF19zY
a66yMGqpJHoqWqEORoRQP+NiqQXxzH+XIY3UpGChR1feaMxlVfBIMjP+D/kDYrbj
8Fj7Ajxn31P56zq1nrHxK9pRCmW5tEvmgLqibP7JxSiH+VDqJFeKgMDYGhnIr+03
IP5sZjBLOKerMFJNEMl861bQW9BK4EaFx3rXL78UOWY9S8KjAKOdLriq60izlIqs
Y6ZyiIB6nYebXi8/eZ42qLtdnQLSdIGmZvq7y6h7vqYn/RREM7u1j/e/QalNU5Kz
gw/dLBfMCEajlQPjxu4/kyvmITeSzrr1te7b+KF0bzoj0uG3QJdISLeKSYpStg59
QndHyYiNwQjmI9neG7eAQDxBGTiPPyyIDj1u/edkvzEktvq5NomJOWFZIZhXGJfB
sLWoKQUwzaTop+9tespiKfWGkWMnmoBrQCnKXPGY6EomywgMnqILEnRkP5hhIl5+
VNyLLItZqX0hDKWXumuJICZQkrLtO95rl1GTgjvDK+c1NS1ieNVMb8JfEWtyFzoa
Q5kmZ2VtO19AvGfY1OX7Bx8OWKedHYDR/mXWZGdCtvV7Imu8WZqRCpcnBLzSbMt4
Z5+mRtt6EhaH3j2MnPZ9Lh63LXSDyaQBzmp8mZ2BN4nx9Fd7ENAJJcHVJJv8nfSE
QFj9/W4waGC4zK016G/thKlJFkblReYpHs+QVwV9C3x7wvdTH+Zw1eAzatjFztWx
R7JHGSCFYaOe94GfRGOV8p6XXMDo2ROOYlmokQjbcagVREVRQUA7qDIlVHYibBkG
AErAouXnk3flwmckLO75EveOn3/6lLELR8FILBVXAa0XZvIspfwULC2i7In5+476
jJCsH12/aedUkcuPzcQpyYNzf4y0jZfCg87UpEMizqGT4TVgqSSiOjGSa3HmczgN
1ZDVn5YsMgiq6Ifm8Gl+6nn7XxDinA4uq28kHzz1aZPXP9ca6ak2XF74Pqap2hvy
NQy4p8dtEYSnnQJBmNmakymyak2TYXyWzE31F5LTAkRJePL+C70fNjZ/J85oYe6d
zHOXwXMsx3GQYsck0tgOAoI/ni/KglZrSj/ykuYbacQKbN3ZXwCDezom+6ZecOO+
nVO3fQc4xshZgw75axmqaCHlOAF16w4XPeA9xpxNRR+02bLehkp0qqnTAtBfhMmG
kBIY2n8SHl4pZSYM70omnBdzSC1VjaFfJk4h93rqQhdWTjwiDVctGw5MfFhBgU4r
BOWC0YPwXhCaaYmbeRgv3VNyPYvDEC4lCyEkoL94qWDTVBKKi2w3CBeyHIxJJEDN
kgca9DLuDs9JlD4lcPVSfpDaJdEwa5RJmjDBGO0k59cvHcPNqAWGsuCJB6wImFGR
zpaSNgVGgoSL64pSBeWPJ6TfASVKNZX+I1E36yWnAhWz7df3Q3Dbu4aoj7b75mtE
5Fq1N3B42pnyoMKYXHAZACuAZJLsJg1o++FGyuOa0M4L3+BBlrEpTvEqKLTA2qmu
o6Q9IOQjXE6UAxjImwSw9cQxVcR8uDQzqwHwqUKXr3UsUtajqVuay+FwpaTOe/bl
3ByB6RvcU74m1IFj7VYpEN9RoiwuDwobsXu1dNKHsUOgjN40g7es5vWphkiH7V8g
Mt0qn4shXniH6E9912c3gZMdnZQmcrG9EfYPdrmpw3lV+W3SmgHqzLnGPtvPL+Q6
ILyz4YeoEvuE1W/TF7J2/MEQeP7Jvc7zs3rSB5rI5+QPc3NqA3A1PnozUGvz8b/v
UNWTqZ4iaqVPz/abJbdyMifPd9P4x7UYF+Wbkz3UMAc+yGdgtbU+hlXiYbduOK+6
V0t7rQsZWJU950REnMrdgZg5FkbJiyQxrT5Zk5nJn6TeFqgb7iSzr95/DYma466O
2on6h0mE5KKkR2rx2pYx1PXyKXO3PKmk/lOM5dlDYwaq/0YHbO7vjKXNs6+QZekE
am5hUeFpyIz+iKzrvUbLzcXRiTz0DEqccsFkze5ehf7+2292P9VpzyiZW6fKvs8X
32yJjU1kfmw6nDbmdPsfV/TZcQo5gItn2LNmtXLeXds+a46AheUsEVU4d80n61bh
OXt3QHWnj0OxH99tv2I4L+CkLy4QCR0lhnQ04pP5CLEhaxDG1KFyj6luHxhiEUNP
brI/YeKpYImHUV6/6lBSZaRQyViXkNCOSJLBRbUN2WAXzlMGheOU0o5Uf6m0Q+Hx
xc4sGQypEhPVxso0SMA4d0NJyqj6lDtzykeQ3fbaML+H15QXWycZew0KdhzkJ2Tj
w6YuEVQf/ebZJyWkb/OpEhu4D3HIehZP4RDEWZYp0IMVvVJLS/MU7//rlzyHGm/6
k7FO67Tlu5N7GC6MJWArF8phtWs7H45RJPwqXSQiaINXQQ1baQDdUV2uyhvdel/y
mtAYLQjXiSSbKdC4NO3kiWXodc43uex6W1aPkv9PGKXlVohDAo3IPjL2keePt1cK
Rp6mQZLKro0H+qgtVs+VFKr217o+ow27L95mBaCTaQoP4W86q6dx4HerflljNuIu
8uJs+J7cKFz+bhHDeVLPgWIQZzicsseNSWxa/NxmXTKt54PQONuwvn4Nf6ZeNfYJ
jFbnzBRx+xQWCnkaBPVfmGnh72fwzRTHQN62bI+akddrcJ4xE4VINFDELYip/abw
X0bSJOhcX21dTLVPNKy/GZeHvV4LDiv5s7xNiJe2o13GcE5uAuJ7KasHJekEjtbd
XxL5CsOz9kQ0Xa+ouVqSkhFgje3bP08UzTxnqlY1wwU5R8M41m056SoN1TaVR4xl
8raDRE5/b68eXLbRQZzUvPkixyWTz9dSghjIcNtI+qf4BBt2JbfiBGyHoPU49j6W
6ZDAkEO4arzS1LYYPPFYfwfQcU69zdLIHt9C1+r+MiBxp5rFTFS2BaCvQZt7PdOs
OeZlw3AEqold00Mlh0ZjSRzAuQzYgUNA9SFed8adALjmIpRU0X8Bwg5SSCAZ8QDb
wLVP4bA82NEuxpq75t7eBXoXUie21asskGCo9KvO8JWB6rpNERnxr6NvqTGoyY8z
RhUHI5BlIb2DvMQQvGEtE03eCT2AJcqQaftB1xQPuX2a18htED6v1Q7TM+09Ctss
/Jah99bmdjp6YwkvkvrHwpcVa5I7XwUIstOBcypl1e6Nj79CRPjSegwoAvBVCU5S
yrH0jnWGKDqHP1O9zBCuiWNOu/Hi53JxZquAxmYH1796AQi16z3u2y4rdYCvWXRT
iD1m9Vu/vp/FJptg2f5VwIbV+VxkQKyQwbZFEvjbLqcoe5R2ZH+onqj0sf64dpYL
nU4owWjCVNyxK4859GiDUsuoLmkH5SOq5VjuwH56N6MO2V4DKqMhx/ojTu+xa95Z
pxopu3zMkII9cQo/vYwARhlbnBqLqNTUfK1u6/1Dc5wsM9XoNZZvd+P3w8ZhlSbm
/dyavC+GgK5UxZHpvXQvIKhTbn++uuN6pnTfDPMZbcJcD2laZchO8rDz7aUhAITq
`protect end_protected