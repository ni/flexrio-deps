`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aMReDmrPskJscpWYThVKVItA5gecPPZO1R595p0GoIq1TSTG+UxXhmmUXc+VYHJ3
u/C3EW5qePLufxmXxmhmDnr9U8/cYC1zLfk44v/2OPb1TBrTsludEDQZdGNWeV9l
cPUMSIfZ0dHXN7L1M1E2XtgoTWQxf3VDHs7B7lU2y9Rdm/ibz0fWMow7op2nWdD8
gJ4QlNl3f9Oiotp1p8vz9RFzzZOF5gBBslZxcTF5+z4qO2W7+xLByngthWm+exIr
3Pzy8qyUo/m2DDwOz3VJSvSNm7RUq+0/yJNOOz3jr3j7ZyCj5OqT/jDAWjJSMH+i
2402Un+wDMOQxi21JLo3cA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="5R6K2aWI3OdbT2A+sz4o9+2XAInTqB1/cSw5W16RnA4="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
Gm/2BIZF5/H5qen8uQizPH9RftTuEE9mgEOF0SqeOKegtP64CfvEUnIxj/ahmIpA
6xUR2v2l7E5duaLZh39Mc1GYsfqE91NCPU5whLaBPg0UuX4cgTkO4cYbW/7yvcrd
4wavUfwXEp2VSiN7EVxL8RcZTSMSI0Jr/aojiilFqVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="TEmQtJ1Dsm7TOzpJk/CeTSSFx/zKExk04H6I8sT4Meg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 57664 )
`protect data_block
nvPqn26PC4XWLLQG0Fq8XsMTlhB4evbpiwGjZroFFLgtNlE6bBjdtwWsB89WW4j7
jNfYbKN4sBv0hDeMH0AAR+8g+TCqoX7yLdIUd7aGwBUZJr6FdDs2wTUxRkXFYNTL
I9bh2qnrcVOdGgdmoQXI8IgRvh/ctc5C0Soo0M+FyUShhuF9y3TJibM0KlQ1IBpk
kG+8hgEfFy5l05aSwjh6jz+0CuKA5+muurxxVXayc1o1ICmcBbg3E1W6z0FBEKru
ZjvbILbT1pEV16fLcmJM/ujIoncU8y1KvBO/THtDGSXGcKcG9Phu9/IBnL3Az31u
oPKJ8/T+MFZo+usDCrRkOHszqIpSbU4owk4JSyx6+uN9KmSW6ODC/dBV98uSt7Zb
EYp1fVBm3CzvUWqkLQuvXv4cgkYZf18XutiEzZVTsRw2cVSF4d+1CuFoVjw+zDi8
wIVN6yBbAzhyALzlzkbJRJSdtrNpQRUR+cx3BMPUT4eJkq08UmOyzDPhULm0LsVN
iSgf1LvZ1NsVt0RjhZCeIF9eIkWMNLApfwbGm23baatptuA3iWTTyMJ5DZY59d0i
Kg8BkV4WRxGsYrvr0IuDmw48F/NyNxyJKZC4sm4O7r5/Cmmoi360x+yt8ojbqvQl
2hYL29eqZzRKaqRDyj1qJhgHnbEG8PKS4oT9BlcfqY6ZPf+dyPGzKBJEgUx5FiVG
S1gkfF8+UlKhk7sjMbtuVCKEJiWVC6xGIwgym+tyt55geCIt+Fijf5FWsWuN/6FT
5o9rRsIs6v4zVKak1qTicqvZ3KRtC4A3WC5MPoamvSCoRxtDrhaAq1VCdYuuBjrI
tvFteXZbD1DRLs7SR7xESoTjoneqhGUMwVWy+HlNp040+9eFoLot9LCpvTg+026T
z8ccjOkKR4bzoT6b/bqyBVTqLnld9w7L8ko1OXBr5oKRShk5TU4mXgzJq5++ry3q
KPCze0UpS9c2+D9LG+TNZhOBuNI4J+LOmM4Xd1sluTP8HQ9aGriIG5ra30JFn9X9
tD+A07roUoj/1xIHJLnC82TbQIGStqDdEi+Tm1q60E+YuKmEU/5BA7bGgMvJqF4Y
9PujFdx0J+L2vxt1q73+jhXnHqxhoas3Pc+0nyhE/8caNDanIaAl5kVjTj6rzQPD
iFC9np7DPTxHIZe34mmdTKSCHxTnflDEJEavVauK3bPUJkKEgF0EtTsiupkZZj9p
oHZjES84sofk2OcYF12uhCWCR9CFTiZlFDZpHHUxPK7yqNo9RnjkvQoXr53HTMUB
3Z7IwfuZbcJQGiDRIEiqcM6UdEUz1FpEPJYnsykZOGYFrzKSlyPkMoBkBkAMWd4k
SFgyXrqc3wnJEJDMNEk+FxcsJBL/7Gj8uWz6f8/jx/foaVN09heDX66GkRswq+pE
t/REyE/jo/zQEcX2a/PsT50zLV9CIG/344HhmysC8ZCnThhddZAge/+kTJWPwygY
+S+vIMkyRifTQzDgDPwYiJ6gc4LxMnRfJrjL7KqHMoK22Oa9xkJA856bGQRq9Ht8
a6NTV8l/Lnw9RRjA+wN70R2ycx/NuEOpUPCDnHkoDxn/k4X2/CjQ0tAhdnuQk3BP
6m9bQZMAjWLoGMIVUJNW2HXDBwZMmFjHjkuABSWKmKAZg5zQygh47iNCiowqTdd0
ypJjlR36O+p5aAQQK+mz/vMW2w55vInbE3elajyufZvRlhNjCMQFKEl6kvGREZAL
hSrc7mZ9nIeTtRaOt7dOt62m7b6zgrMjcfciqoljY4dJlfFlMoXF5N081VGy0eKV
yGs28y6g26GAAo7XF5zZYsbrycD7VZPklQFW16NUnGjrOe1Gohfh90iht693RBEp
UY20Jto/nU7tpmdTqgD/di5jXHeu7atmXGxO8+OHZaby85JfUmCw6+3KLeRc7fce
4GDhw4tBalUV0wn/n2GoRl6hmdTZXr9OISoPai+wHs9NH1BAGsoEnpdLRD/NkGvs
wWot3VXr2XIZJ6g9a83jGgiPRxQBwKMn4Scb1qzk+ku2odh76OOSBrjVjiVP60N+
kdZYWwrlTtZLb+e+dRZ0Qd5Dhtj8doMj5Kwc2Az0INAKmO/+vmVAE+mP4i38ks0S
SpqWNdoD03Bxieoh/ZpVq7Ttasm0l1I24d1dzf4rRFuteG8vDP2rWobaDWJVJhhl
s9g/Wf1BIazAX33fmJc+joK9PxCVY9lnvWpzkmnX6yK5IGHDu+LCsmhxf+FQuniV
tQXBsv/qqaS7VFCb10W4cdNRCbGvRbQUByC/XLRH+t0hlFQ83frnc0H5EI7NTrww
x12Pz8W31FZrAWWW0Oq07/gC+l6Rcic6Q/BqaMhvWxqTPtgMpROqHtMgyCe/o5KZ
A/f35wNuUdMVZM8YXPcQMeAmYJVoTmYyfDAD6DNbya8Fn8vmbf/wkRtlF7/K08XT
2OLitqRIebTw2zmwd6PXjwo/iwjQuEape/pUKBq51tMQp9t+VwEFhy3xh27oYlGz
SQ7tGGzkIe0rEQjWFIzZ3Hepkt2So5N9e+0LMLFfNANmqNkwMext7E6JmoD/Tg5d
V87pEEWcTEOa39y6GiDh+2FUQ0ABxEABxcrxsYa6xncLaupP7KbPq0945tdQts30
XmKRhazZ4bfSAuB3KsnQNR97E02rd449BxOuU/uPwPBPQoFpNCUTnINR/hXAxtVC
yuAMj/0W4iR4jMJnf5YKdWSMtNVIgdYkoUCalbkAnCPO3Ae1eyTOmpbEjYvL/iyE
a9exkjHYbi83MSLyJGLN6iL8XCjpdbhp5wYblsaYhnN2+ZVoFNZljaCBf0pY+/gD
6y3BE7FhFmlo3wvxG159IkenOdtl22423DqZ+skpXev0kiezDN6sEl/J9HY9vXIF
Yb/l075T0URPR2p4xa3mE7RAP765Eq7c/Zz2iWAE8ORLe7aBZAJOQgJNQMTTprsD
TIeyKVDSko81k7mpo8iOVggriVSw7qHS9rfy9IXutD+pCLxPgx3Sd2QC1gckcZPo
CdDXMzZw6oF9Tz2DIQ40bpnU9Gg1S4k/4GDKGYhPbgbSS3Ex06HEZatzkWUuizYh
XcnuOuA/FAYUoPevcypUV4JLdG8S4kajBSOnIMMwDKPwLKJNguczHNucXFTy0D5J
RX+omgl+Joe+fdaz+TBs6eMnx5ew+rpkrJSC0Karq/4SRCjXEa2vmukoTebFINO/
WYIgQArFXuYzLwILNkbkXkOGaRALPQkSZugo7rSwB3gP0XVfisrdu5b0tkmg13Uy
7suYLwqjVTBmIqCytUp9SjlrjQTM6g0wajyNb63+XQBlRsA9VruPUanooNjffspU
0LPhsgQ0h3Moa1RykPvPtDWrf70lHJQM2jpvr6vBmsQpkrubVbeIHkLKFe6JRbHa
2QFwmA1tsfJUf8SabEK6GmQq/LrZcgKoK5AmAG47HjpYASn/zcwnmxkDnnkA9DjN
AcMrhoo7DhZdPJPw1vftFBRV2mdLSWr8MRk7lGOWTlxrRb+yK0OCeM1Ou9bnuSF7
Gzx5jmqlEgmQVV9AYPhcvjRJPfkPankArCCAcZv+r1aUs4Y4Gnpvb+JoIKUTAtAA
Ic4jZunEx+gO9ANI/JkfZeNM/7mHVnq7yVAFrGRUrd+Nq9wlk3JYLGDtDHMtZj4g
KUc+vbRPS8ynsUDhPcbBcp4SUG3Ku4mHbUXcNw1kh+y6vpLm3dFnZEEkNFA5zqBu
2zPPP+OjQLMnNVHzxhSI/xPVJWOyuq2WNJPcLBHqb8RS+puNw64adcqLL1GYhAXM
5XjJwCjnk7UrS9IMJ6T+gtpMAYLxicMbNFlqnsTb7pykLlzfjrn5vZCJk5b+yrIj
R+3D0mrmmXptnkBsJrQeGv3ukhUpGTdLiOYOZgEjlcFPmQk9rpL58PA45W/17g5Y
ZgtzetXNfEH0lec8kAwzaCcMh3rZSoUxgBTF66Dq315BG3HWig4FBlqqpao3DWFz
A9f2U/g6eDquw8NhdIHBqloH98eYaTuGJKJG2UqNK5uhQgUX6Yq8+x31hUNN+dZF
5A96gJcqK1exBWLTKa03yeHSXHMqLu5ZodLsZvOuYbFLaNe3Uk0rjxwr7oiMJKlP
uLf/mUDknluAKMw9zoildlRDEjCsGWDBd+qseYJ0X+2BJSQGIh63ws/4M6mMoV0Z
UxOK/DwPfs6vo1wxKNXROBbbv5KSSne2ofk1cE3WGRBUR44WoTUa3K5LtSXP0IJt
hMdcaJrPiL0iVg4yQoefUl+ab5xfvHCJ7foMoSXYtQqwJ6ijTn7VLWnFB/iF5pQu
7teMoG/vfks6RdB2ewzeR6S9qB2FMdRI5+g9AutfqJbB+aYlna8wY0CUHoI+jF9Q
UeFIAyxdEEiQgudSpAII+kbJbnxtlDlDkqNpwLt80TTgNybw0ipEKAWohat1YKNf
iXFq+n4CvDsKsTtyM6w38LRFWh7NItwuQwbaDt6CS6+lP6EJhisrFp5YKsC3Otho
+txumwveNIVI/t7IJlVVbR1mWRNmVxE1EiwgwWpKJINQXlmUpjMKIhHLRQXMvEcO
TKNOkfavdBGPSvB71RhMFd0LQukZ7FfGBPi7leBUDny7spdXI40imAPs5ATCmdoI
ZN4tNIsKdgxVkh5N6/VMdwPAd0dwAbd+r/6+cd3I+YqaNv5++IGVjR6HTCGY4wdY
MQHltIE+nKVCJz1Ht0ZTviRGErkIrgQBV1Jt7fsOfrQRQBWCac4VS9qqtRyZigOq
9WcAtnR5dOcwGE7iCpoW8MIK50YK9ydy1kxgh79JPdcb/DJd4K9OTZ7X97VcL9jF
vvrTnGXY4nlnSBnR8p5MJBP1p8jGaWAq2Sz806s8gnARIIGeYF8GtlFhagcl90L3
enWYMZch10faZEp5NkvNQ8xi+Azslil71h9eStC4StkH7qDhxyIlvyASHj+8LBZ/
BXy5/WM7bMkvNQg7sznyNbYbjVK09ke9/bxn00cuqCsmA01OKpOLUdyOTGdaa3C1
12UkuzZvo16+SuLar3ltkStPTOjaB59cUZYbgm4Aflx93baKIQtPJBvyuJwU2Ytg
vbwwtW3vRaOnroOYLLj39SGsbeEOVb/QPSCLxNfJ0fIq+0beK8AIXgh9Z+O4g2Ir
hDQUfgJwbPwu+9PrUR6NyoDR8X13eCdbaMe+oJvndb+O/86kFN3rtZyFJkt4GbGr
gJ9Pi3/SUr+WfJTd+nTOJOlUZaYmRQHdvGWDA8CTfxi1Md/X9w7cRW8xnoYiyMXf
opeGtQc2NQvB+LxQ6+xlTB4r6WAscCJG4G9G9GeRJEGsRG8Zh+b3/AG6ujvOhP/J
nhvZ3hjWAI2+S7TbNPovNu70kte9+fD3f4G90pFBsGjjxyVhzvd0YlYzWMgKvYiL
bhlVApwy/JJnfG0QzGR13WmnU93ESUkjB8uDet/nbh1SExAeRtXZY+Gd7rvD+eIy
lCwmubKGdpkxfHGqXWZc2g5Hnh/NtdJ8Pmsbfsll6lqw88fF1+RxPwe3OmAxO0lo
oMF4zcCSg4Ba9b77glDkHC21VCOJOemRMsNJW5HConnVvB6txrMupQP2fma6xovz
7iwIu2ZDaYeu3nc54557lFMcLr/fhCIpZ86O4DnEXls28BmHZuf1QfKZ1eoAcCtq
H86PcjYRINbk6BRWKikGXNZEybMxu5/FSVbrcPw7+L0xQwTgl4VLR9+g/KLZQdXW
JYWnwREAEHB8xHn/delaW/0BjvY/EcScrxqgyvosANj50WTPdFqtHhhPpVIGwjES
gsrbd8gmh4X1z5odMHE6quce945RMlOl0IYXL5BgrmKHSwpPaT/ee3KcOo0as8ng
TaVSHlkwFL+G1XH0Zmq3rB8DCqrus55wgLQi7OU2BfzmsZ+oc2FDmL73Zw50kE5A
k5ZJzBB4MvEUXDvBmkOF8VXxT3j6IuFswBLBAXZ2qV+/yq6MlxLVp3Xs+SXi/B8y
hfHG/8jr+y21HS8eW34qbnG4kwtwbLFLa2Tuu6psshcO9FNxnpiYrlEmEJkBANKS
9WkjeQAUZIv7dtChHUjCLhON58sn7F6sToR/9K0hKH1fd3sfr3ksPRSmuMYt2hGD
rI52P/PZu6KAoJ1QyKBkQ3x13vXODxVizeBXH/5/prI2CD1/I7ZyHQUlFOV47cNL
+c4GBLVApm9Xa9uf/uLu59qQs3XBa622BQXp9TxKt33juny9nShFVq/weW6H79LL
sLwdTl4lvVU/W4f0xvOaPy+QIAxPv4QbV4sCSgChom2cTbig2se7r9S6xTHhoGTj
CKD5IB0hPqdEe3r5bsIgMpC+RpgXkQS1/irRZgmhqeMvbS8uK6VGrAv+CiNtdyTN
hpLMqqD/k8tmRe5cCaRszVO5lr2jyfw0/YLAnVeqsWLw3iwmesGx4QLisNLgn/re
scT6Ds5KYqydkAzBIRUXu7GupgU4VdlRfyABabaEwCXD50PofuK5JpOFgcMoDfMR
Nvmx0Y10uBcoiGsVID7xDcbbCEOGq70TX1f7nRqIwumdL5V2eIMqWE2EpDEsztFM
/fPDs3l2DJUh8QM5Cbhz1wOz+fnGUQEZwC6uK7cGaDEhERValGxYVWdIq2ay+rg0
8MsYRc58X0Bbd5FvR0HTwYsMc4Y4ZlRD0bUVfMXmAl6FgkkTj5yOelpqbXqkxVi7
EdjQhIZ9UQZVTKF/l7zP35N0lLd0ZlbnabMWdW0rgSuJ6zfzV6sSeRBw1o8ynFm2
9u2g1Jqgaykfn3nVKH/xDCkbwLj36diAGT/pEwogBF9ZxVj9IoEKenVBG1mx2YDB
d3/0a8BzJixtpdRgGcq7i1KmiEIPtEnhOtPV4LOvJQwjPPYOzur4OJJ8sqmszh8x
fJhYXkeEnIdzH5sfZKXRsMgv/jOCOBoR1j6ObI6FfTdETAmYphsXvRVbAFuo8+5b
LRC8sBTonicEISsgU+Hvm27L9VZqNSo+JTwezAefyE4ZYv4rMbGIzbJijwvTqOA8
s/wdSjU50lNLe3Ctd5j/9O1i5J5FThNI4FnyEXRAK6jhwQ6hDc2GZjVP7y0EMYgc
BOtMDeCXA/92HP+MbTcvHyoX8ZJc1a8FUFQ7g31jQfsO+jCkQ7J3q4W5nAkk04wG
4d5tFbZdZB6BzA8fSqt6RruSAXU6sv/NHkGNrjhFup55alJd1G0moJ2xtnAM7F/k
v1+2POia/kJI1nQUxn3XYs1KrwDoDrnsh7exNimKw/v9amcjd0JP4nz4e6g2DMmA
C1zCS04XBpyr2Ado67iguB59bD27PoxhoRlp95L0pv2U/1I/jHn+wSuRCztMkAai
9rQNBpAB+TX0458FAK3U0BoQ9ZDfsxuxDmHJkUngXedRwGHtOd4i9NVgZjNYq2je
jpqR9+G714K6flGWCyBWUyYutvl28thlBkGo38GahOJgBp23Kz++1XlizboLKPjO
NvXytYHaC/jW+ldqY4lixGigA4FgV1Ovrv1GxvH0Oek4iphPh75O7c914jXWbKj6
WDgqzVP0/fQkL31vYzUgLcJ/N594pCYlqtvyDCcPYgMEZCyQylDoLV4YI+28KVBG
Gpwcig6bTEXoKaKEPan9H6HULAQgpAncfm4Gmp6gmxRlrAD0QY9WClch5QF2ddQK
6MMrXCOwlrdk45RZOrQaZYhwEUiHx975juSvda3LVI1viUqy6D36klTzpXsxkW0j
FoDeWjkGwYt24E46SPytK+J1wKn2xIg/m4osI1i1WkLZSkJgfkEmS7fLmDOTNzk/
glXjx/FRta3SgiR8zjtpL03iU16eArLsX/pxDSRItU+94x8H3DYVsnRelEC0MFQY
iOOH0PAI76Z7fSWXAjvSGtQ+Eh5EbDuH1gQjkKSldsYYpVuQyI0ti3UJXyDfxKKv
vjl41UoH6NZ4fugHXw6zsInnDoEuUJUN2nNXaXWWX07pRxKOtYAw/0rMyxgynD+i
lVCkecijZU8JWe4v/UFUsD9JE4VYr8MINkYgSKj2BTAHoK3CJ6MyMUtEYhy1eiAW
SNfFza26iwBbWoMzAcTOSwTYvn2fPuAVuUJtPutdSPuy0/epcrSrYNavY8VH5HgW
9dt0nynwiC0WGzgdVgtvLSVQPWmCi8J4URHDe0pLtgtb2KKQubp99hmscM2Hy5MX
Wyh3ldJr0echyz6FmGLQkFNzUV2J+rqeALGSuARrjBX0DkbT0kto8YwmN7qOtTPN
6wOUkksWZ6Tgd6NIYxNcnbv0QJ2OozsmldNQmthZLSwJv6YIlr7OV8Pl1rPNkgDZ
0t8WCtUhWQGSXTJmiwR+uHpfnKMSy3VTcW+m4bIMSVNixpys5c6O+XaJVulZjElN
tBgsb9VCjiYUpPk3o52VLQ9p76kprCcfU4KqoXxQUiC1Yfoy1EzDFAZqctcbI3nb
fCWp7yC8vh2hgVi+27ErGVI1U3c1HRLHbiwP71qFhk7Kd+3QQjg8KsA5Sc+iKIax
ApcXTBgX32rpUaAcg/+oUmuzT8fvjh/IxBKbEc0wOU+LvZCxfQdCOnwK5U7z190A
OgXx5+oZox+rcapQ63PPjW4gTo8j3Sl+5LviX9mNP9vqdz/zJn3IbF/m5hiZS/Oa
lFOMtcgNW/rByVXpQJVFv5NDYNpA8Qqe5TyqUw9vK/s8cTAN9OcveARWaObjOi8c
Fp7zvDgo83YI4RcwV1xH0xN4rqyGseoawFReClt+7Xg/3DZNqeodQTSDBtRlsdD1
4QqZfmFOUkXjauCKJMuPcsJl/D/cQ+IBTSAcgMZhRbAptPxYSObUCt0bkvn2KHRn
2YN0P2cQseQwvXjVSZk2FEPMfsvR2ifcYDeqa5IJ/uWNYneo4Fwshvg8YElog8hf
w1UPRPfAyuHyxyc2ETOdW6nhu9N4D3Zjh3fGVo7P66a7Zc/K5j2SeP1iYYSeABUy
Y+Ye0koX/A+q5MIESm0ZzqEWc1N/wEazD36aTNIf2TXAbrJeO1h/vBD5zEr7E6rv
HORwLVYk8ROFjxuJ+eGAVq2yD3gSDKpgZWQE6m24ImVZhEJ522vFWhx10PmGi+qk
TZ7ivKuofNRLTa8gVjGLkvMDyLFyzoKThbYaOm7WkpHb0k9DElE0uanVvrjG6mT6
8FxI8M3HLDWTwS95jvvH85qXzDZJ14zjhZMPMIcT6Vo6RpZilHgtOOxm6C2Jhvl6
1SMFoFXfiRyM+/s/tZEzW1dggW6v6gd2HWFzdau0r2IQ4UClvqdlwp8q6rujKDzj
kEogGM1JkDne8Pq/RLbc36pTAN4dc595dRo6IM56ylEjpqFyILHd5/RnGtmrnL32
iqGAr17Ya3CLZCdVfogz3sW55Ech1m+quy7KRQU8rz6JKTAFXp7zflpsjWk7Epi8
F+O2Yn48aBGvNq85H2T/xzGvR+AYkvgnZTOhDGZJjtbd+oMN8wje6E5dBc7IaXzq
udCAzTHJfFSceJA5QKPeCdbZqS5gyXPDXFBGvPHQRCx2G9GxmG17LGi3qj7RpeT7
AV6jm1pUwk1RcyLcdK46fhK8fdMTT/I5RfUpeCa5vkDTy3hNOJws86LanXHxT2MB
12zYpg/Gr2GDvh6D64fg7ubMUkZ3MmNj8KERkc20kjXrpE5dimhz/GysQsasjHr1
lvmTm+QkyCDYhULCI0ZY1lDVVq60CsBM8Y9y2BVJ5tEamkqpebWVLPhX04X1Q1LA
kwU5kq4EBzejWMksS8kwA4sxp5tDnL1bhvD9Za6VIJEDdwO5kGnLZ3g43npHbDgZ
o9pw7udKwiFAi1JYpqWyZTeR9xJuavBnJR5JFBQYfxkwCqUZ93OaWPjpoorMG0uc
11yO02bOntst805shIgYXie979CkV2BtSFV4iplIunDi2pomSQbXSsUGNfyFEEON
skpIdIH9GjOv61K1BBvtwyhJ1/oil232VmksrJ2c21P4LH70/9TW26YKw4a+VCPB
3EjO1Vq7eI1YCc6EpQ3RjMFOqzucGDqS3tXz9GwDx/aSLuid8nCYr5wkpgbb9ZC0
ifnFEIyNMOBYTpxzkjC6gMLaRVwTvnBGxRlz7OZrxVl7w5KEV97GjyxZKmadg/M+
kZ3DSTv6pz/dNwKGX2EUdVkGjQ9r7sUAbvYp3BMj0Pq3WL294CcJyQS4Re6ostKf
RfJUiuiUkza6l7ep4KmvmkUev0iLwois2ZNcBFcXVStg1KRphlTkDLlym6z8QxUL
R69bq+9lQBzFH5oRO+QEBnmjQe/WM5IeTbxXfQuiqixYm21t0TYMgQeGcVoUqQLD
QhhZswW+E1bn60dfQV3Z8lIA/pmEcNsnmlf6fHP4J2O/C2R5NipTli3G/N/nK/jT
zCmaTh4U0YVODKBWS3W9gEvg0vFU4ZH9ROY4GLAtlJlUny/oj20Uldet8/lgh/62
yrPhl5oBmid8vVan6lLg48ruGkpkoSEonb5aj/tnqt78xq1hkepy7PZtwblqqmj9
k5cwPW3k6UShAo6ojv1ijpBE1exFu143NBP1f4HLBSw91wrLjylLH8Huxyol3WAW
hR4HgmF2EhoBEqwxmGBXZX0aDkT1dYEHVxRbcBkxIvnaixqbFuPpGGssfocXQUo3
VbU9m6/3GfJSaYqinU9qYlK1qSJUcoKczoBCyxn3zJk5kukzMGWaYCDtNZonHiJv
zbivIYrCl65zdSs5rsW3t1SNr1mudYwypiTHEC9lNaLje+HBZkmy4AuGl01cr62J
rMy2V1qxpaeta4BBfjRUAfFfPkmikHReO7m6tzm0eSbE8yp7JgerwsFVpe1jTA7o
mz+SKlUKCS/nc4LXXjFcGurwZ9IY3oK7U3lpRpUtUoQIA0Q0OSdEsntOZ2lRg/qZ
wv2f7kTAUeamzXzHl8iUJD1JKFEQC3wVqS6VEuvt5t2pMQGI7NWKZxG5IsNVInlk
6lnWVqsuVl++g6+M+p3IFMZatWf4+OkERnjk0owzCzB8izFL1ssPM3l8Ylcahi/8
HDb13361zVTgda0waqG6eyMpZtYpPxURE9rkzV4XzWEF2E4iTrmy3pWGquzLqFym
1AG+jNKKiA8ZY4vRfuJb0ZyLQdVG9XTEmCmqEsl8JoYVDJKgwOy0kGXc7VHOPvTz
Jadk9cqbJBqBEh8ks3YgzOoFkIvowS/vEGXOL0F9Y2dv4Qe7hRA8pNApBA8GSQiY
O562lTQTRCUdESfBFJQV+PkJrWRNCL0c4i1L0CaZRO2yXfAI/b4KLQmaz9/33fIV
6HaNaZ5F5dFo5retzw//sTBVmeN53oMcufTZ9TzJBadPZO90aRPiAOA1g+OqdF8g
/fZo4nBl+E20LBjY/wd/9l5Ml5agvZDD4UPK+g87AcOk+XmrvA2cg9IFB7ZCpr+R
o64w2cHXfPm61oUIpw7EuZd2hIF7Mn8WpOfaZuBvSu5MBr0bZuWyDbB65cory8A9
QVafXgGoLWixUYnajKQUIDwq5lsusajsda4/0x1aeVzYHqNCYQvQ9SQ9YmkL7fi/
DMd84+MWI8yGp40Uyczcp2rMAzuDRsOOD/BtEQVXeCLgp0Yrw+Mwj0qOi8SMpC1K
4aUq05NV8H5w5r4ISs76/NTMuM7Qpjc2fZHywBlN5IXvyIFPUK0eK+TjKUn9BlHa
X36wfERb/JUdjWAQEMZOmAHJSySzoALh49w6GOcDfz5wJqxpvj/LTac5jiDJOEFl
WfyZCHUYzVpdHBzG5fUhwk+bCSuEzEZ/8ry55lA0UNRCmqTPylh448o8tnvzTK5G
MM0FC1XxJ06s+QXyGhG7jLc8szZKDZKlYZCFPQOzhXg85/QO8vwMmNepRGg2IlVf
xtaRYFhz+eUmAem0TOYpjJ4NsbiTjCzspu38RFyHBE3ekXFmdM89hpDzZnYytl4e
YJVGUekKNc+zZey4RnTNRdi6Tmh6VZgXkm9fveEWBmmJr8vXOatzDIQc8w5In/SP
46kE+YozKWOogtsc7kwwpfIAuPt3D+kw+KfuOOOOJR8ELwumRbp06RFciuPC8e3V
yc7Ik7VP4xxjgQnB2z+WM7Q/WrDEBJNjIpk5Ls0uzKzqVeMiu09Mvuh/lpu8zFlx
VdsA9OOHC7crcM9TJ4x5rPi/tcqeCn2dtoNxGCqHOZGQBgvqHKX8WhOSEBFulOsR
qejh9RIz+TVf/AR32vCVWnig394anu9zKFZNOFDiPX4m25XrFfxOud5RdbiotH8F
unuYw5NSiBTER5mJW0RvZNb5fdrnML92c3AA8qrBL/zli3jwQ9PqlITTjqslR35o
0odenkrvYkBbzjlwp1avt2g2cfbvPTWgGki0u+bzfp5BmB6toBhBNdSqFBc409pN
8vXlEmaQUthSJ4ISeqj9rbkW6gvUCXufh5iQfXdmBsVnGF5rvzr2B2K1TeNFpab8
pZqqusuIGb90clYkA9SetPNkXIHSr7GBu0PrYCa2gzM/klrJgMdpVsgeptd3J1YR
ODJRQxtJDYkJoRJkEf4U29ejZvHWszXPDFcMqC4AD54CHr8RgaVOL0EMAeLN1y0b
wBanvsUzDZYAzwvWqJGL969shUHubYEJFyHu+5kotaXo03ZD6BXLXTXhWCNbXohp
qQ8xp1Hepx4rb/LFM02G1yc7Rx3xDdv3PANgQiNlQTaLY4Eggq+ixnYvMmI+4Hpi
Bcs28rUJ0oTXL0NvPlIpgGvz1iS7JBVlt6FVP/+eEf/rtgQiwXTrXBFVXBri5Mv3
p6A/oiS1wOoCbApJM2FgeYQXpTJzvmqKjYy3e9SrZKCQPFQBQ/ZYKODyh1hQzKoa
cZOi1kWwupnUsuMT+prpF2OYkrXryliZsWD5aLbvT8CF9QCXS53cuOkAFpdttnRA
SpwoYOhSmVqWvcuebk+j7vT/HS1Cc/Cf0Cw4Og/a/l00/acmmpL1jNoLGYiRv2p4
YXmJqDknlIX7n9nj9VesoLD7gMjW7KsIN6mphucgfD2iESs7Tit0uX2wJ5+l4OSb
2m9WmYyOV/td4QOJ9lzz3esOHP2Out7jFl+3mJ64lLhHKWauBYsB9zuiDWGazw0d
2cusmPbyow2Iix4vdkhLcxMSLGTTuv7pAmEM14scdix2h3Iml74HWpw1I0R5NWSK
AaFiVojoVMbkayeD1DVcqMcr4Mudd50+g9LVleg/zEEkJptJriKKv/x9DlNqe+3i
Ju3UylzCrJJdMhIYf+Ns9sB1mlDdam/7Pp5YWYv2kCSaHwmIqp2hStCsbHGlmUdF
K0Bajz+NILlX0xBlvyGqmdmb7rVzZhNzFwT4B0mdcFLd8dmit72mIua+tIVnxBfh
vUGXEyxYwEnFSvLAkzbYaX6oZVgbKKiDaNy1CdOtOvjRl5TZOnp9XwDOiIzJ2E6E
NTHu6bvpzixdjSllMy62VPCEpje14XX7vecIAGviOWohehcjyScV8ZL/nGcULjvT
p3I9R181M3jbzBjn1GGWDWUFboXoqP6N1vkK54DOrVH/gBdLVkwElEBf3zyLhxAW
jwd8QWAQrBKBPTOhcP0LnKNmQwnoYu5uXBFluHI2Ng9mjZG+4OkRtXsH05XxGPKa
r1yJIFvPA9MuZrSy9zDZMKACAYuOXDT7+0HjddcLsl+IfsDHdZDkBNlHASTBAkmt
C6HmiwjEtzEXqOqbQNjkTSJNpJdk7wGYERJTIy8wpyVgbUr8IsH4AXEap2UKXS8S
lPFudZXYeq6/zObM77VEs0ktYG7XX0coxGjiOIj4UmV9RsKQ2YB5AwvXperIqfQJ
tifNhnckcaPhivnRUKNkxptf0LWsPsLhqb/Fj9tA1V1liMRCnHPonomjjlo08OeG
V+tkMmbgVx73z+ChTrlhwtD1Ia26BcwMGtq1KG9WQhCrIi/x4SPYoYPGFqO4NtRz
Zs2D5X/OmeB3Vvbk+wCkUbXuVbLMq9YLYvSAsV4mZBODC50MaSrVIaQVkBODdxHB
Vnt6OAHtD/gnmVVzvyBh1GMDoUJoJBxIJ1eJG0Yl3K0SgynRg6LU3Y9wmeO1kgAw
z22WFIQYsvESXtzucoOXlhUJMOoWqF63dMGE4JT2wSxwShRSZypUGgUjr5uGkGJ6
LGaTn7fME+KqRRRm1JI2n5JwDF5/LGP8wQTRCpQGpb/ccXyUpNsHv84ksJgM+RPF
Bu2efMxt7MI0L1hYG5FvfYjmPhIGmqbv8Kw3HXD+adzmNKM8S/LHReznoNIsF9Pj
ZPcXOTiApNGuwh7OdJtFmS+fGMYeMCK94hzG9pfirLGB7cUEog1b9meUiZPtB5NA
7h36jEPt+HFlFnssZjIxvgO6KGRSq6c7fpA8jhBlNJ8ZU83UZkoNHcuVBjYXNAd1
mdljJaJySSSRC4ZllqmHf/HDVJHVm3YEj5nYD133HK10WqP/QmcaibXK8Icf7Npi
sc2JKDo0lGIayZsqyZqjZJBqs+DC+3A73ZYCNz/d7JKobJQA4awYDTQ84NbquLTU
6U54dTqrT4BLR6n2Vt6DfpGg/9AcF5yd9cZ+wNrm9s+jTck/AKpfdE4iKqINn9Wq
yisqseZEPzfXctiJ0u/v6IN40Tcr2nFblR2UMYn+y0B3vRSchvKm4lKH++Acj2Ej
+Ei88NyknKtn1zYXiJwnV2PQqLSJf02TRg/kQ7ZmhfJG6oSkDUbF9F9UMdg6d70j
+eCiSm9g88OIZprkJ/pSkvIdutxXp7WtOn0s2Q7fspIdaxUUwATUxTqMCTL+opqy
QDynk4AEIpXjXoYzjyEyDSEvWMohXAPATr8wjL0G9CKfKLVjoL/sq5pOocjERLze
J9DG6ZHIOhMONKG7A+1edd1GHF63WjjKJnAVWBZM+3tefL+2GdAphxRZVLh2jvGC
n+8d+nHALZpOSeNC4HmlS/X1QmGxZ1+ZZs7QLAFEMC9eoDE96X+IUY6mLIEzbFpH
+aSl7cRlhLLwhXZ2hUXU/uDp6hO7NZ8Yql23yYF7bxwJqDl88flSHFy3FDaqHs1Z
sQEEkxWfS03TnkhiPEpZaOBDFfE29ptrtJG1PgWuZJ2OhJZnyPVUHk+zvfV2pyTl
ucLYi2yFt9g0u2gcYwJDIUZugQphGnN8a+ediZhsRj/RqIjkFXcRGMBBNRlPyKOn
KdwMkGYg/a6srAjap7XJnV+cs18HQV/FYwbWsfputfLGEFfoLOyp1qouaINL8BOE
iw9T2tTamJSypa4vmQaSq5oGPn4N7aOnhdlcDLzeA+bKnMQGNJXZ1K3ZXYlN5MYF
HifIfuQQTbbUm1xeE7Ed6WFgDNR+nx1zUEJsDVnne+K+ASF2iIY8F0hGB+zjonyG
QoawwxaJMpxVpqEIiFj4IMsQyIZdzUkH5ABwOa4DLim86cTLWd32qgM5O8OdVxXk
tHkEJ9gK5qIv8bMoKVbhjJhmCrRHsPoLqTGp0zqXk5dUQPHOtxJiSn/1E893SCbP
bX50zVFytsg4Hv3wucPNluWJ0MxkPlCmLbr1/nlkxTFJctwU4j2ExuW2mh27F0q5
1FXfoB0sCUx5SfqQkF6ElvPajZjgKs8dvtsMYFKeH63e/9feQQg7k8umMd12j7WI
jftQ7aSyIvrKRnfhajpaMm6yIL87uMXDLsvjDCvjyvh1oXNC+V9VfNN7xX2t9Eiy
MvnPjH/gJuFo0uGuMPLwfv2pJrfsWRME2G0LWyE4iiHgqmycHCsY/2PdybDi/sYp
bw1WH/FyX2ww5WQfu0QiYulwmkAlTxySB/MjJoFlrT9PKqUkTWgQSIVI7OHXIhhp
2PSiepESRasLhcjKZQ5vy484jLkmNwGKRemnPtuu+ZTDzqhfgfL+HTTYUrT7eU0y
tmf005SXDfLB4Fe1jwPTn/NNk/+hQ3kqCFg9XO3OG2TK0OtKby6kT8QXmQIcjf81
UAUSCb+Qi/Hps1KXwyi74qh5u7HvfYsoqdXyIsWRSvuRskKr+Q9OFIpCi46iDq1G
YsbWMhe8up2MyK/nVh0saiJlo0z1tovaZbgt3W4hFOWXTbxRhfeoxpsuRnAkYHjo
WR6sOQzIAgVCW6XwiWW742YXXI+oE8UlUovnjGDx27FXW4ratAX5hl02fyyElFon
AD4czu1qlno8Yo7oRXoPCgpMcyAUnAP5L1IdDMPlqffGzPiA6/9ysvJOfsRtKoW/
kbU4+kDrmILNiKXcpM6nfX8OPF/fAQT9QKC/Yd807vkWeI3WiDiPq8SC2cV9J9fI
19au+jJcs3dTtTBr4ffTIKqmFpC8D5atqHy8ZTHoK0imiDfYjpFGsRYC0XXa0Og2
sd7fX8qmlWcAv5hshGBRh26DiVwHe9DMaBq4tp3/1+Qi1sJBxdwzPve7DQzPAz+E
Ekr//ir4xfgkf/q/mmLAmEbPwKLHbaJImDEMfMoi3Ol4F5C/TctoldWSCagDtqP9
ODWSq20BAz2IEYMOnJSK9U2+nGTL127jVagxP5VJL1sgsNAQEtRCYfJZd1cE4jds
oZx7isffjHQyHLHdH8rH1L6s4QQKAPb6v2dsROGVH23notr3fbYEl8py2fQZyJGH
q+yOANKe5C+LldL1oCaqx41nmI8cZiZcjS1JwTrcalvQxMqmocjgbLpI+bKlczTB
RISrJUdKL8rBibHOmi0Iv1J7iZel9PjsK2MevYfCh97LW3AkedTjjvPPKaUYkjyM
quwxoGUxwH/ZtRd2UV6UGCVhOru3d/vooTdcdX1CLyULcNvKKn7BPTtPnxCqj6Xh
fP/q6pTY2KOaZa8x4+kcHZo1QtCmTT1byT12wDdm2NMlqEwHo9MwO0kCQ/YJfzWY
iaKFb2KWDUjuFRJqXj73UjfdvmJH/1SnRriJa/CSSI5F01T7GZEZRsQgl/D7h4nA
4R4YxlA6kPO3Seg5ojHNKPIEm49rN0WwN3XJg+B0CtSCKtUDibuLt7wJP4NOBtI3
MrNgzAklZ65aCCqpikRh3t7XLJ/diso80fz7uo+U2V1aJLnxBXz1013epeAunOgo
eSYWkNEUza5pddqqb6347M/qLTChgBFIMqKcJC3wJRLqrttC9cw3QxsSoq0ttg4M
UadNTI4qXbRCvgNDVEkjORpZc5w8kmgYig+QsZOzXtrX9ctmCnypIROjQVxSEBW8
KZDKcmbOLBmVubDAhoyKyBbQXaxS0TNWSdYeL9mKijlfejFLU9hN8BalOoIpgeeL
wJbbtWYunuGB3BQnrcB/QLkNn2agJ97SZ6oH1T0t0w0TibJrfG0GQn5KkEFplu41
j2ePWMpQnBhuMhHnI7OJio7HK+9YfvRxllbcnonDeTZsEZjeB+8S+kiBcOrCLPqh
kUDkV41NnFs12Tth41Efsb8LnSuZeLp2TS/rXcLWNxLB12ZYiDTd7GWhVA3pc0It
YQudno0eDtycUGNQbGMXCQLJaYL6eY0KqOUlPHIpxWMkUlT0dp4XN0io3eeIyCZ3
rA4FCsOxK0m9EYEQ5/z0E43dm07SU958cBW+s5rnlrRo0o0fvPEzGYvVWgDLIg7F
vqK9vrZrdyt/FNbMdJKhB6q/2sHX71VOtPbfpYnGTemUVlMtbC4PbqZG9Cj7dOlK
Z9hiaeaOMsmO2mkMIxGB+VTylcIGvpdWr3D6h4K2U/GaprsBxEpa+5bWFGLM/bzI
lHyp0yWU1mMJiIwOzy1/31zWvo5wNs0I19SxMD7oZfvEDfMl1YL2R1cyCVNz9vjN
IC/yjAAHTsiYp3HLqhoHn9UZ1pEHNlRmIzYgA4ZB5t1ZR/8hMiFvanBmZ3BALR46
JtXviU3DYcpkwF6BITImjcNRJIYQUJxDTEF4lfPa6phEbthokLLlbIFB8JmcpvvI
fIwTmbLb1we5t6IqdIFbZ1bWe7TtUiNDktLltHvyIU0q9erNwEdibxASVdZJ39T3
GD9SfDyd3prf2TxRBjKdF7/TyvL4mAUb1mtjBGWnVICTBySSqIzVWdk2n3Ury5Wb
ixxi86tPALBK1YOxOrRloUthjy0XrpzEckMC2034mnW6d823iJFwq+R06mmB658M
86ecYwyxx8wuJioBqEtsaW8loSwf2vAlvFMAHeFdg3gzHPdJXsWc2CR2uDjgtL+T
Sj3wWmKMqh4ujsJWd6ee1IZW+PjoLR6fL5304yYuKhRzoW+uGcCARZ29yP8xV/zm
ge7K1aiX5FXM7lNkb9oFfaQpmG4Rc892AQtFBrWJ0Na79x57DrcJnp4YR/67MbYO
9UVej5tASi7Msbzoma5Nzfbgf+nZawLIvds/gfcA5eUZeInAKtYV7O12NCrbL6zU
SR7GEPw4mBrwKvmuQ13hYaK78ms1OkJ0MKaSyyngH4pSoYSIG8m2/S0SFbg8F7Tc
MCk6zebQFOPkAYCWE+/Y5kLxRQ2wkmVuzv01OtGq8DXeDAAcRoRlPP+YwORF2A4t
WuWUNMqKO1hR2lN0x58NCNE/eGWciWbHtzHaskpM2ox6LE/tqHMlj74MQq4DdxkY
biOUHqZN4pOwyoMa4GlranZ+OUKKqGiDkeRnxl/uad5QybIOscpmu4n+NAxBA1i/
eoogjnt+0S+htNQaXkznt/KozuS61KVkhwpeV+/3ttweOVKtI9L+jnT4AtVH1HOx
9iMl1AINky10G1sPGAoiL9NZrsHvYDH7He1FF3hopfkh8IhtF78ct3S1H2MAR5LP
g9629XxboelfeZoVxefcYdwGU3zsiaiUz62v/sZYJjvO+7SqLZEMq2aTDHeCGGhw
kDT8fyWLjG99ejb0rVcTpCrHdzlEoTJsbg2n8pJLn9EvDxDZ9m+VksTHdnboBYRA
c1/G7si0tixUe3xmHRURwBjVmSUF84SH05qFz2xb8wDYo2NjszsDH0OuV2d6cDaH
XeBUJprt5qtm8BSq38TV5Nqrn78VlhR0b7p+N39jMrpFHZXGMgiVHnr1QJPjHBJ9
9x3LmYbQsN9vuqQW12AAsDgPVu6pMli9ja5LmBcCq5UyummmAT5x2xYr/hYnTmGN
86aaPp2Gs4i0YdwnxN59RDojg/FF0qo1/u3q4cR/6xrtO0SIGFp8QlgoJzV4N8Vo
DJzC1ytTUvRdW6Ex8XTQJPEO4RbDQdkEuV7nHeoC4x2+3bYlEK5gvFVYoln/TN/l
XFsMfcrEqHmbEv8US9X8Zx/0Bq10azBI4e4mVWvjxBlffo1LTn5y1bGuZhe2mdiw
NR7iNTDJLMVXCyovVIJLSiYyH2FhagHkTKel5fVeNt7wiiiKnUOz9MJk3oIyztaR
vnux0ad20Z5/isAjkhSxf8H20JT9HfiLcOdjAeYfimhUKKSKOZQqY9assPxu7I0B
iESJKzgAwE0rDW16H0pROqoVu59Jy9W/b3GMy+BCQsXA9Rk+3SgHGRG4REwpFiTB
SfWGESgHdTeZQ/MPwGt4roJJoUisHsqWlI29LLAyJleyy/bEfrhSVSM9jHz6RKUV
Q3Q8rlrJjKSHmidjPK/yLnk15FX+WGPApfOczTsDZ7vE7kiVx6jf6rmBQBXSVutA
MCjr1WK+TreDUg/iDNDe5t+bB8VdWA6/eJeH87PsTA66ElyUjCL+SsnrrWJWlYUD
1yWRy5ho/ps7sV2LQDEch8Gl7DNAZZkbqs4D3punuHUGkQwTxjhZC2c8ypc09US7
/L1NQndT5DiQ9sgzOeZSq0KZbkdF+rIDFc/1bA60OKgrVe9/GKmBSSq1vvT1LOOY
TUM89WOtNITEIMqrkN2NvH4Sr8i4okZb9bmratTmDcFthUkMhCi+K54+dYFWZzZZ
3y9dl1jI3XkL5B2zI6B4coxgtLvhg3/SWS4Y0bM5AA0keo6u1/wd9IYCC1aymdZk
Wei4uwQrFMQcL7YarhpA0ljDOGnzD3Vhiqmbynjfpt8+6S2Gwm3loXU5eKO5UmN+
iP65MIEgnIKHmZLBpcBEDqLWQkS9tl///kS8tAkueE2iC4VyMABYb7BVv/4YYEqi
fO4z999iOY6OlRiecrQsk5cOsyYP35iVvwIwEFhvy7ZSWlioAyf9WztOOtRX+liL
4GML1AmAwuY4ZwM2PIpCCbs0WvCAcdsjeV84wE826rMPLoe/CnhKWN5sDpvLkvBg
FQeFatfH1V1QcNXWUk6KwPcA1wxJ3sSZg3rRRItulxYdUoalfG/0CBPPVpefmC6M
8p4/IHiaroavjfTYVc4zsYX5+Og0zZ4G3m7bV6H4yuGB7qatiKSEWtwASAErSS8N
6f+jo9l20G0JJUhzno4LveTP1tSztLw8lxTTm0lHPGuHGRCL7kXDi5wQFIohqH28
RtHqgN228edLqgEHPEhFeoZ1EIqAOqOjtEWbgxH7YJA6dwRJBKIrqeNAKR7Iil3Y
hPy3pa9052Np0wkkUruVUJBH8Lh/r9/Uy9a1RHTy0fBM6EVjp7SDcmdTr4X76seO
xPC1rmfGxp1nPHBGVqzEUN4lQGT4wTy3j89CUblWwODMBqO6mopZ+tsqMIW5/h94
r1EnAnyUdrIX0P2XqOximgMivBkJMMMf5Q892Bo7T4tWaEHUNx+A91Iudg9q4Xf/
oUqi8uIONjZgtITvnFArYHuN/TREEpT4bhCNgBTafgl2TIQ+w2lj6tc1GWZtT1iY
4YHWQRfD6C05Qr153jFKU5Gq+vRiR9wNtgxbTqQFtWkaOaXHU8dv5vkivcpKWkCt
fPGbC/gnM4HewroX8a9H+7dTvLgSNTI9OuyA31dcUq0lVi7PSnyCdjTq0d7LpWhG
m6fl8LyrIQPvcY50fx8VGViqppNX+pCUQtQJEny6EDB+6CvMYcnQ4M+RvpyJ8not
3uWloweDwm5nDmzmwQ35wZmqluKwTXu5tl3aowXhTLQ+DjZcJ7TnT68lBzDQH86F
UrCd01A+jQhHYBewBWCe0UsTjTZJYhbo0myNtNDwgnbPivLd4UFF0sW2fJhRz5t5
2dTKulcFlDY7HTJ/zpXl7D7mVPEtFFjDWSuMy28hfYOGns8qkMf9rdawp3UPp6I7
uVxE5zpO/nmlnZaPUh6JyhSxO79wkRfbEUX4EjMbAXR9Oqkz6Y6+LyAWxz67DvdR
b9ju25edbZ4v/naymb6rmksv4sqHVAACCit+yU7DnzS/0rJEIEulwRwiqycBw7g2
C4fVnWNuyscuGm1WWd0ceAxQVS+TOFSU2Xr0IvOWLStHOisFi9vpvyf3YWC8CJyd
1XHUuevZdXyOKEeFurJw6M4S3FJ2txd0yfaQ3OaYXHfNYWlhJh1AXf4WqklaJ8ZT
rPpW6+sU3iIIkVtqjzl5kqEAXrASAqxOc+1iXbSWrmVAS+5meLAdWnEDPvjyaXl5
2CLaW4kdz9phz6rtdwArEtw8JIF7xz9EkTSavA/nbCq5LhyoFKLEetJnnr+YCpnJ
TeZYp53RBsBolQaxmRZ6ZpyInn2lVmR2TNZcy6OUQGDVswpe8LDGXgoAuLETJZUs
0G5tkJT4dDnP1jLP0p8DSXpgbPNexzCDqLy+QLON9g/EdO+DInSSaji10KUjPDhh
Z9M25JuPGo4/6yJJaMxjc2maPtrhfobzG7Ncrlua/zrJy1GZ5vZ6T6FY9K7Sw2/P
aTLuDuyyb0RSvrxEp8J8zYiwRIvkt418FRSFrdfi15Un511YCPtcu2gH9kHNbpgb
jos3ecvJS4PEuKJrQeOY8T4m4AazR3tGCqzn6GLkULgf2ua4hl6XHPt/fyRAF8rp
/GK+hTZkvs6nCITbiXuk3PoLLGkk5Og8BRbm9vg2f8X0IScSRMHknQyaNVImLC3t
eaUoyUCRoucrEnfg7AqITjioL+H3D+YeQAJCTOjsEQbS9xR6esQdS/5qXr+B6IpQ
T77OUCeNkxOyBNvkKXrXz1zEDs71rwmcy/OX+9sHR94jJhsSzCc6NOa/9s/o9/ta
wedqkJ3EdiZVRzF4Hg7z/Sb58QQ87M+qjYUziDbf213VRo34Mt6/Y4TnfHUCHV2G
vI62aMX2x0UmAs+0xTXrpuvIY130EU/ML/lUk+5xJ31VbI9rVLo7XetrSz4HTkSJ
1klzLuWBF1VYqJBbqymT4ZgraQbIbPAejQUZfl77gk9LUJLCEDJHUqgfN2eODWHI
r6LsXPl08STfziBKLxhB25oX7nIkEOM5fen3oR5kKuqSzap1w59zxK2OAYVRgowD
hOxLpjx+3kPZGoAE6oFBqNu0iYPsroUWYw8nQf5dxyn2Dw7Ieu9lU7klwL9PxYsA
HahqaR/bQNXFBYgoJiv3V11jcgX2prTiSAMKTV05OuavQLiVzO6LCe49gD6lx6Vq
m9LXaD5PmHgXl8inQADgppM9sgk2BUw0rswib/M/gSsYpx5bob6f3mIAsfM1n/tf
K7UATIB8aqgk4H2HomddjTyNtdE2HDucVu7JJj9ptygzAWG128kDU83C566AnUvl
Zks5LNac6a1aeEDzN6150GCVLiZ4mj/iYUJ4Q4/5wuSDmBFznUapoK2O2Utv8S/v
f841y8XROoevgincHd2HNzQHVf8TXKTf5RzcHScPJrfeKwKgOAIaASsxe+asFPtl
bsqbMikpaG3o10YNA9EBOBhBqKLzwWhrTbjz7LqCEaIO8X7zU1kFdzIGrkFspQMF
Y9U2BrzzVG6tEZu38fMgyLwrUCNBujVPtowWQ3vCe4ti+1JALVIL+y/U6sqT6gj9
sQiBW8bLzrrj0Fk0sdbcDG47HL2RC6xFGIVsxrnO5kf+zUSOSWxhraxDU0AKGXda
gk/EI8UTsPrrwxNvfbjH4DT6AWUFo/gt0aBmBYZo4eLyhrCtHWM/7F6mPzeLwrVT
ENxM2hNWt67XFNtdlzIYZ77FsMkpZyzebhn9wdroK3OYW9hn3ncXGTH0GKgp5cIn
juzQZ2W9wMh9vGq2KVXNAeMmLbU6C95Ptxn9YsXPh5JyQRb0bHiytUG8vwHXM1f2
cR/exGPTXVfyohRSi92uioY6p9C63mUjeGyK77Q7J+i3EqNHY4OaTmoSKcPKhdVN
/Mh6rsgcnTBv+lQcQmVKsOAJvdftOmgkiMFwkf3xMyEymND+dBzzrde4GXlMKTWn
p94SLBWHtwKtL7AYaFj51Cas3PtNc4W5ahW64P3UEs9MHyUG1yNre3QCuy4aXn+2
5HsTcyNDeNX436CMGB15rTFJ0L/PJHwxt5WJrosj7I2cfstig21C05FYTsQIwHKQ
6KExbDwoOvq/unCKPAEQyNLcPKMt78tHHGSZgB+R/1JaYhWxmUEy3Xi9iox+VXvW
6TsLbeBv3i9/dtysLqb2VSSfBg5oTvXv5i3dhCye+BRDQGVF8DOLQpDzSMFvVh4R
JvhnDN6pTMB9TNR1xOhBBe/OTcEDJYL/WyTjQ6sjLEwVkiGnH2b53TX5S0caFL3y
1W/Pr/IiW3qztAiVoGG/THGMW0VIbVPXZ5LOv4iZCutELzGI1WwyIgSlBGKIJ+YQ
kKprn0d2IL9nbu8StBNkm/bZHHtLSoRhrvIeoYwud2ZpKC+ETAUka6CaUY7YkG3w
NyROEXeakFIuuzCd83dPPYyCRt0Llr8Qy8U67nklqur74F0XzX8tWI8phYpLKsly
1qVt1n3BL8ovipVqrWZxe0c37QPcg03Ehlcb6RNxrMFCA5sLLBw0Wv2WVqxQn6Qf
31lz6yRKbqX8/LJx9WNx0lA3tfzcDX+iXNrliwakgisgKFYa6J0FnD6snQ9oL41c
7bbvTxiqxv0SNS8TUdetbOhq67zbBBF4fMHPvY1krGznmTDh3XGkvdjEydH1TmNy
2hohzq/tum2sLcCR+TWSM2LjREeSvriv7F2wUJno5uHv3tDeH3LF94apQ7KdvwaL
teUIjNH1IsVMGRQ4kwPrmnFkH9Az7DGtvpg5fOd50DxnBcpoUKWeK32hJBEt4kt/
5uia80/7+NW6CUggeCvPFbcoSf06ukBb5kbDx2pZx/SA2Ibj1YtOOJQm+H5b8JPF
3AGXP9sME6SMu2ZxlY2EQcw18SpiOzo7XBJgVXPw0j7aMyTM6ztIEY5cGRxA/yxO
EiZcbOxtYv3i5gIgDUNcETnvaknLBbcjHEMgIiEpPHm4x1egvfS0L0ZU5d9dhFug
ALiNl4sX/gXUJAAuClBafYeSeyOxaFq+2ZIi0HZI5MKEoJy49myjaDAe4xRHnfXW
RF5z57bts8vwPGuaw+O9OY9eca1DfH5aOR7KoZkDvCqRgmsEIBoZZ5dg9P9gqL65
GJSvvQyXLTB5hCu5RFk+8juUg8i1pfdiy3egWWE2GWVkH7SlUMu88CyCX66WrbX9
U1JuVvFgHxUrcwErxLx0XQ04/vIm5yyGNrw8L7uyNIlqDOkPJLTHc/lIj4VgYCCT
OB6d+l+eKyAoBA3cpoJgX9BzUKRP0rSDLBikL2E2UG1SjQnmlCceZQAhe7UdUiAX
eerAT97fL4KJhoXaGXrXPdOPhAv1AY/IK2hXpjFpo4L4Wader7Fyrakgg2O2inwt
/At6QO4376zJgs+1p15TCqNs06KXGgi1PucJrlwOLTGP7g1vSa1bBJ42d1zhFpxi
JRRa6HTmCZ1GSkFtEBFHQuOWB3ZnmQNOF/1eUMmAJGu0f3BVq3eznHFejEqADgVJ
8+i70+P87EvOXpWWE7d2zH1q/98V24buk9K7A1ZmP0EKYZAd5XwdFFHWCx2sVisn
xcEy7TSI68cwTmy3flHweBPYZGGOSs+zSD5N8KzitbVAX1Dqgt/q+EkJ03CXLvgc
SIlxky6IOanZK/GHtEE3C45xpIEQXf075fgxD8NVLhP1lx+eMjNVOlabncSGPFL7
l85M4UQS0yBrlrxNxDv80+VEBteh/jxSeDG9BX3yqEiSNTQvrUb+UT/k4SI7ijYN
yiyxWEm4efB3nMgBF2qxuwGQYWXd4viR6CQV/g+9yeo8iSlguNFVyIWnAJftKKqA
yyi4294mJkE+dH2SZ4jNTFkjFX7ZEPlw6eW1UGgPGSOPQE9n9zj39oyevNYbmBBI
+iauCq3+m3R0kxqPRy+G6qHJGgNpQdLHLOAG7mKNyK3jMi4Th/d2GKo0uhmGopn5
HG6VwAlpJBxRSzI2nFNXMOKhw2Zvl2V9uwvUh+qWaAmwJ9T1Oofv8qw+G3b4UxlI
xWYV8xd/ZGURAVNU3YqxYGOSHp+cpXs6jiEX7RD4mWhOxDFm9MHuTgkqOZklBL3e
FBayxIZq3lMNpq1NpWitJeSD1AFIzFlYoiuZhWari5FrZTbX52j3frzs3K6b8TAE
1IB97WvQ2Rmd5S4pxWElgJRMErs8YtsTbmkp2mBTlbwKlGVIHd22K/aYb6w7Ua97
VgI9L6yr5em9XKyuG5A8gEw7UyX53oJaHQFRXcV2ldApRLCEZYzwBhtEEmASbGnh
/MHPR9pn4Tkmr6Xfy0n1RHOqkANaDY5lS/5iHyMUsAUxjLGVk3mvHqvRCSfLC4dY
FitPiuwlxVuVw8c0ekYMjr9aWrP9D1n/jqUwbXowaOqvxt6d1k/Z9IthlFfsnc9g
O/ZfIlOA8BuOF6Qgyu5om4GL6AlkhfpxGmTy7dOIrdSq3cC6vNwxj6JMojKi/Rkp
pwOoAuOrq9hCjbH1rb1YeRd+djmnGUqeN/sfigo8wGVxr/jwOlZJgweTCAUTQhcH
7wOHhsaYUeL8TFNUAnMsfEUpHai4QFjN2ewAJ4oVPkn7Y2Czox+1teDMZg/L3GmZ
EHottm4D5C9xnh+/0lLgYLgNUZD+mTds5Cmny6cV8r7xrecCIQRzU0D6z04oEpxN
fpSC8A5pxst+0Cv0OlfxcOG6blUV6B4A6LrE9We6qV1uC4RlCGky+rPBd/moXh73
9pH1RL5INJwjfbMwhXUaxmPCVQBqPQX30DfdSPupRAGdWeDqC4lO0SICfh4k2RjD
gWNf5kidt8SDgvumyFYopCrsGyxXr7YP5rY+jwQHULUjHcvcY14lyNO8tKHXtRCF
YbNg6BsrnKwoAgXCNmZQOMtr7TApaeoRh2xb1X+AfMj2Tqa2GxeOZ3D/P1MbHJE6
QMwU/K9UhNs5JP2v1QwWpSdJoFkP49vphIb9Zfz4CT38tlvWYuQEvfKZnaDDH/kJ
l+vtxJjlhd7kEmnYaNItfk8+09vMy9TS9oUotkf78gqXLGUSB8CH6Irrz44Offud
Oj5diOnDKQ565c46OLX6DJIqajBlUt+ZCisvZFUf/p0rjm9vv8+U9t8G6OBs8ApU
9HOvH+oSqUAy3DfGrmrO6WiIJolFcPL7oHjx/UFGmc9DPejcTZYgX1NNBMGJrf8n
9XzF76Vd8RWLTa6NCSTyb9ORI96VO3az9aahxpaYRNwyHRYWppfM/bK6xWQHw1G2
tn3PpNXkqnA8xUdscTJNZmh6XBxB4Rd4Tw4vH0w3UmkbJQWeMMInyjBr8Qes0hlE
/JzMYCg4up0IZfmpUUxy5CvQLRw5H2ZrLaIj8t6vTLHemHenJAGfQAiM5IczEqeF
l1Ao4O+gnMX6q78AFlgTwO2seje17dZMcDFdv1NnNoc2RQEAvdhSAZ6EPcZNLvs/
Mzmyeq6IuZMx4ssKIHHEV+PDZswTsKeGk9ithIKOlg1TpGAxY6Hewm5OZ4BgKP/j
U+PzjDQnzcE3ZGoDQfLiLY5LJqQ0Uxc7/Wn3XLitC9CCGEyjvrdRkEUBccn5EOg6
TE7ThDz6I9/NI6gbvKbXH+2wo1XpUVlk3mI8JHjrPHks4R69Li8Pd1cRcrukW16Y
1609DCIMgFyEU1xjRp1fQyVNb+H95w8ZXp18MBlEXck9TBw2lqFq4RSTNT9LkvWK
nxbjXsn6/SSztpsrIaM7PaIMiJEYJDK8vvBCGjrItU4FqJyXh5M8YhwMD/clmgYn
Va3Tk8GUo7FSvtv1UkrUlX3cxPPgr1NvQ/vjTIt3Hh0wa1InI2NOD0F1rP4th6QC
6z9ezRCBNrwJjykLPEpZBZk8WCVNdm1/qkFs6S+w757WpCb2mDGG6JtslVZNamrE
CG6JjBXbV61t7bdsI7CJDARaghoJ5YBbCLtUTk/hhCGcQki30haKiIUA3EoXnLAW
BwAPxh+QaIubyQfXwbmh5quTnzdTdGPTAoiHE9NwowpqrUvwQHJZwUN21gxoa9Yz
HBr98aPjNyyiLUttxvn9sW+g2uDykW/l1c5x9IPhQjqANwGcjdAxuI4NRxJKaLej
0lknXj8daeYswZt4TBzr177XAOKmTu+z45IFC9tZFqKJifBj6b45FosLwgs/jUyz
BlPPVqsGp8AtHcCksCmUefDGQSQcihR79gTcNXl3FIRsXja8bpaqLKCX//ubZvV5
oOGIWCzF8fI/U3IJkTI3t4q/a4XF3d6yKAnV/rNrzi+8uf1gbJvzA5If6fK6waxA
VRhcvlzFsBNKQF/HT2/TiWqYe+rparNjS7P8/jOmUNDrRZ1XOrRD1SMdQJBTlVC3
9wOthrP9tOzrLmrsl5QwxmYQXA9ZHTK7s4/JRkOvMhV6s1UQWg22fyXK3GYU3NW6
L6RHikiOvLbcpEAeQEIVwnIueR4X2gQcZff2Noz4xObASCPbMRNH6IK9Y+488s0H
TWuE7wXPcqe4+0XCZJDWYtpqL3dV/GMRBg0oK7UvFGZr95GM/wVLfk1DaNt9i6m0
XkyqKdmw//gheH26its1pU2fHCsllVpwavJdNrh1Rt6FtvxqqUoITHcs5jWElfj9
1AxGY3jU6Azf1kD1uoBQIVmbj2y4SSGOssBbq6EnqnfhmemkcizrBXTc4l3NNCpN
u2+X2UA6gtc8lDrl0WA1o47/6RbgxUTtgWZrrxOQtg4wNMuzZ27/WjTOYPHdQEGJ
o8oJ7/6DRyM/AEpieIIO8q1kWr45BQlv25DTwJIoRyeUK0MypknZ+3cgsiosgNv9
+5cnC4QTwfeQp5ea2P0yZL7iM9Rffk0WV42ZJ5SYkGsmnz0j3KFupe6LswdGvPhJ
l+ezZOWyxHyCGQbUiH/dUm3cJ8OWcf9T5meTfptuZe20p8HZKnsMjF4QuLN6k7k6
3egUuWqAnMhwoyAtxvMCVK6T8S3rh7jlwZJoFEzXN/zBracge3VgIHBlu9Hd/Nyv
HKanxngwlaiu3uo8GmheOovAC9wL9qqmorGhX3j7R7VsrKbQSRyPf2GdqAZGWvDL
b14rMLYeeaVwKpXhk2xchyvAKfvKAnffK1hlYAsyEogOPCKF9xRdFU7GCPUWeNwP
EN939C5R0/20D5CMmQ062XxfOxC+NHs5q/BN/HfsJUlJH/SsBoDR9Rl3b5JR+AX2
tR8naHvn561mYgnAygHYxaV/m0Le+i9tdbcpei37mM0aDTZa1q1NMeD7H51vXUCR
pJ99eWGItTNctdeRKEXOB2ysfiyoYjeO/6gvGis59MQ15AQHYNNQaRh3e7PwSyHL
Lwrjxm1v0HQ9Vfqu3merX1MAYwxUmCfpk6jprjpxDUu1yedEkOXazwSCot1lGGVD
eEV1qXyNqJy++syQ8A3GQSSm8DJ0YZFAseIjwFUi2pOsVtk2JNWT2wt7kBouoN9t
HlF5SuRKA3p/0C5m/1rv5+56+Iu7mJVPwfclVn8qpUy7olz+tz0W6qNZdp/Be10/
E9JxQPhfFNfyW2XE27C3rqolz6Bhln7tXrAPovLHOxbus6cjToJZzD1214jipI46
/nWnBu5WweDtr4ZYc6/Lx5imZP//kPUpMVZnIq+mkawtshhhnL9cdogUX4bj6SLG
fA94MIvcEw+IkA7JdvmI74AtmXfBaXlBXA/uc8Aun/MZ29O5VkB84zljOUuKS2CV
6qQkFBfXwucrKpedGgOEfgJXid+2bJorGJxMCWROBINUVwTDXf1qBrL/yi0pB9YF
dkm6DYOsOcUJK67nDnWOtZKj4jOEXrQS65sCHHIhKqOY07ii1V3tcJJbgsd7I7R+
e2OqY/XxZlNBskPnSKUSysYMU8aydpOXN5QD9FGxbGyiwoAq/IzWTYqy+98QTHgN
oUgcAiR3QEqhsagNabCsjOgHdUVL/PR7aUPsBd8ihLK/0pLP/ujbETA07tMiBN60
mmIvvrXH0Zfsg2sGF8S/fH2VT64j5yAI/4FUKp53/KENDwvVMPyzMa1eQYI2Utf3
+e+fgELwsYsGwEULBaLsIvitxYrqHS9p2SQPc4uHqFGgFme/akxHKPpCfwZt84bd
HzDF0zqvWbZUmH9mNEZdVwT22am+XmXXJzLLzyCSFexIjMOOKUH5Kxx5qXTdkMLU
bqIKd6RFMdhdwOgQGQv/F3xPpPEDr26KOci9AADOx5qNIvwbgMkSqbd9KSEBTpHy
TCaGDMAK8YlxplUbHAygTg0Jgq8df2YMLxuSSRcHJmwHg5cKYBtnuKyuSyxbSw4T
g4xWOgFws4LZUiOrnggO1YnvmYYpyIF6lifA6yetHcOFiQkfnJnAzA1bRUUOTvLP
O7Dk1dDqUD75psPrNPbSOho0SDLxhFyud6AGPPOLszOWO1ggoJHRm8NAin6SDdrP
ittoUBJojIwa+MWV8NpkpB8/PJtbA/CoBf2MsIPerzPnHAnWWTBe5rMLXXN7mHbP
CCp4y5vO6HgxgdyVJEE3l4yykFIR4+Ivn7FIVHIUsoK5ESw+0swj6rYI8HcOxDVX
Ff9LrvdaUh2dGrZ5wJlg/VW9BJf0zR4VdNiv3ZMaIAWybAe4+PVSM0lDiEFcKwFE
7LMyDerkRXZaSUuXWM1EfQKygIzdzGpD6kH06xjxedOil2yYRAneJD2X/SxgYsbO
qzPQOKLtgk//vyZX92SWgqwUwPfDCZFpUEcmz77BBpS3+Enb17yB9zNYBII5PAZG
ye6VGBGzGUUzYSdADkBbT7pW6NtgIvNbhSLGsRHGUqopufl9fAhNMErrzbXXJDXn
tt5AMzZTvIFBN847lp7GF8DgoD0+BYuUDgu6btgoS0RrGhpibJGLRrKEQu2gnR3w
qlv4hTdToSxgxGUWN3LInwOosx6cgtOurseytu3opI3LZy0xtcR/RgwYneC3Gy0z
Qv/VoTC2xzW6d7FDTequo20AVe9LX6wMvtSlWJ2pzXzhKwJuAuxUZeSXk4uZLynR
WWtZ9WVFkR52DH+U195a3hpU3f2hTpf/S+AXBw7hz/logepvy01sJhiYnDgdwb+h
QoeVfvf6MV9qGmK0LalHxL5xFtc6C0WZ5U2Zem2E3s14bAvlA/XdBJWOuVAr8zwb
NgLzLGNrTpu61lLzGD79AK5OnbZG5dhVJjuMpt0w87z3lLqQ64FDWYb801Qh2/wL
7g8SH9mh9cTC1rRxB0MvTqgjTVysr9pRGtVHkMq8aOkd60h/9ITKoycbW+CniuYX
WfRRdThC+JP0WyKKHy6ANWSEkmGyRNAgJFsVZmTu63ANEvZEqrYHYjPbHktlO/xO
k/O2+R3PoPWGtCZcfj0G4S0JV/yVhrOkCyu/BJUZoZ90DED/VohVOy88hVNy3lzI
ATOM4x/z9mgR3t9lwQMVnFuCsxzxGKyvEiOU2qhxm20mwhTGACkeQwG7AQdTUrtZ
YyMZauQtsryT1RS8uGGl0iEKDoCaml6wbdLhh5i7Lsab782w0XmPbGsHbyEIsTD8
EY8gs/RtmaiF5YAsdSM6iNyfV//n4KA98pvZ/5QWSbmO/l4BiZCwGXvh9/OPBy2h
HHtgwA8kTyAcPxaMlhkBGdZl4zjaU3MvSR4F/Vez5JuZOMjli4eGecJ57ryNu8SW
MyFasnox09yV3sfnmhObvkCroWDAUbZ93KzOG8P4qByYsqZp0i6eaRIixERABen/
21BuxV/X1wwPmrgPVdDmlWKDDSVW52Si2xj2yGQP2czzN3LgyMDqbTL47Zb7wQZh
/6T5Elf6bL+BUdUtW39eFWcIc3RlC1OiBgpjO+lH45MeIlwaRViYy/X6z0CFBExY
HUcc2UTkxRJkCz77tPA48/ful/kbNdTvdH/qfKtW6IyFTYGzjSVB/P3zzOKQuDcR
voh07n5Z19bqVqdfyx1swKmo9R9y8vGDAq/2UPdyv/GIjF3/Pbg+dQ6j0n/gbDrj
rAynRU7IY3uggUJl9x5jCXhVRl+HDgPRvdHlFCJmNYaexp+NhE1b23fTykfonuyQ
7MYNWZbCrkKpkmIHuqZ6VqpKCEGLusJsTBkjZUqqRZ064EjEDIZtEPjFACZ+dIys
6IkTzXzLHsn4cLEhaa0QbP9w6jsA0PQb7RTjHkj4UsWe+8MikQN4ak3AiR4Oaho7
KdB4/g9RH1SCBbuT26dM+uURUUABHj4XYo0aShwXEb49pL63za/b4FqwIYznE4kt
XDX0f/RAzm0JKHNpYYvCbc7mN25GpzHnG0VVxdEyhs+VG0FYROArwNuUm/idrth2
fAZtR1LNz7ET9fsSsz6evWSVLEV2mM2jpzbQt2fTrjFvr9xpM/dC/F0La/xjRjEp
Df6H5L63SY28qLsjlqFbUYByUMcJty0eQ6H2lVfCdo0+B9zHPhYKYhi28qzIQdHY
IDhommTYmOe6jIgxv8BdBAOg0LFoKPVMDeQ1/+jdAC3HqIJyZVJUvr1IGLeuyxkL
keFNBRwqv/2leYsZ859LRhcGBnuPX5VRGk7E8yJNVkhSeboLTmcj1EquvGRKKlGk
lTX60dqCVw6z/hpgUrYlgFE0IwbO87ZBEEebYmUEUC9mSK5mwfWdBi5OyzWZzFx3
z1rza4PmS6QlGA/la18Yk7y8fObekoJHB5TLq8fTeuMp96mSVIfeRvjjBBU5KdJp
f+VmQ4zrhDysPR60KPrFzKzNqKnm+RaCt6tI373Hs8h3OZxHfy4T8FmSxlEcx0cN
fQSULvcRB7HPl0tRvA+OVKSKr7qPjilHPuSkeqflBzh4SwXM+es5cxgPYnqy7CBh
Sqr5Fue45eUM3xzstxz5fobLPzYFgIgOlCgHgig40hRYYriDNqT1I8BXYX8nobX2
2r2fMyvbx62cgdV9UGfqgJtMVRbynMIlG1CAURn1m13tqiUs12ymed/H7H1u6ltU
J3+in9BjqMzIjVWj/GZ2qJZHs286IABohJhIQS9QaP9k0VRLggiLHH7TCStFrgRt
faiO+7i0p9B5p5VfZVw+79oVXAT386B/Po5jDlwkGnBYcIfGSXAYR/MzYTyqt81S
mr7d2VwcLohW62aL5JYyN/Yzo3t0uYpMoyyL1LI57NrB+wC/f91FyyB/9XbdgQcU
s9v3ED8yaS+B2QBw8SdUjZsVzyJeUDDSMWQYavxC6Gf1Y0rRxQtBUFCb7gCw0+Yw
raz7wCZIzjML2m9UFzADYM58iN8mRcmmU8ZpxTkpy/OC6DRFutsHOxTNVIgOsxg7
PIn95S8hCz4vPRICcrJZoxOZN+y8wTd57mxnJgNUR0GMjfsUyRr3ux1A1PTwbvgS
MMIV810N9C7GaF2togiDbPOnWidCh4HlIrryaohctRSKif9ovuyPxeaJ8Eq67oEr
pbHCPrkAu+Uz2XEfquDCCptyaIow9C6QvHTyI9MB4/kXIX8DQuMquW85NzIVFfKt
PL5eo6ITfaLHKEJ4UdxYM+Ona0dXJeWdJdmGNM6puD60LPRW+BeDP4UCANHJGU9+
NhzhoqwCX8bhnNp9rp5JSyQVv3SmeNRCGMekjgaD31s1xiSd0OrDdk6ZLlcQV+00
LaSh81QzSFJI4M5QLhmfsrOrNs94AP9J3OZkNIEQg3LcY/aorMFw6Z2OiBH0AtlL
q17NyJacdmj5spe3Ok+y5uSddeE4hlK5FgHMEMjfM8B5Mb85EUJh6+4IhkBSouH/
clKpN6Y6k7T0OjNjAgYGG/ewHbhvG9+PjssVF9R+uj0nUspA1OonN/mm2d/MyGgN
UEOFT8C1wKwg4JvGEuUHEQVsGZtWD69t1Bq4AanKtZjSpD00QH4d8BQxxkfhrHHd
jTPd5d26/91tBWmDsoHWdUCHsDi4M0+JOotNocrOuqvhOEyFLaIZhtt2/TgaMCtu
/ebJnS+36ap7sXlneooNiqP9sya4KEjiWivHeR6BKomdOGeOUApcF7QjQeAy2/iS
+bjR/Md6ipvkGhtDdzsvm9PL+QDiBJsH2SN7bfLCM9cC8rt7HQnofsfe+Aa5j6AF
CyA2PIFJj/43sKQQD2G/fJEdxWf9fO/P87JY99HeOpMC77072oZHYh+rkJX7Kvr4
Unywim2ftMia86dtFkbJvJrkTu8TJuG0MU46cNJdie+ltn+oJXKR5M38zmeSNOrv
MBq5GQUFIygJi/wq0nk7l025ERFjS/ifLTrDsVDBAYrHFUrVIe0obWZXPMTkikOq
kLo/T2Zffr2O3FPmsiYP9TFgcxxcfQiR7r7M1tZrmlKuBhPN3+pjRPbRobgEVjnS
7PX8z73BUyC1A9kMfV5PevSo3f0uhp7jfGkOoNGOPbFuypeaD9MIzmMmRwTOcQvP
CJIbKbJ8zbKi80bBHzCp+Kx58N6VCDuqVmX5xJhmegMY9s1Wqo273tkmOV0M++O8
KXpPe8LsbZg4ifTg1fYoO+RZ/qhYwWBJKJuUvSUYLkeWBEmY+VjZnIYpTml+FZoT
/ByEtXzn2xy3qi5gwjHlDV/AfxBgiGZMKKLqtgU4g4Q2e3/QSpgTtGe2AkWPg1+4
P9JIMOL5NLrZE//0xlQfdi6Vc5yIDrDNyvPADUAhdYoOf29Z1qy4kPAuMGwF6MCA
ob25+Zq96X8jACr+6o029cd9nAamozz0Vb63oJnQiOyAgVA0fKufU/tx8y5OBquE
GQpe4sU9XO8BnAQ6iuNS98eh7PrgaEIjsVb/WjYNwgf2uJSQw9NruredHWlZx88h
hjOlMthORM8U1SFg9SflxO6WK8GKNyp1/tdw6bJLPlqOUE8pDoNF/uOdIdNY9wPw
+TKl3IazZz1KxgLUQyJLl5jH9uc18Zs4IxEx5/Q0bTaj/+QnAcIMuKuHx8gcJPba
0oa/mqi0u/ooxSGpF0m3UmiIUf+aA67rkVZxYsyj8hMl4ONgnKJfhDaddA+e7+sW
HYen5ophus64TFUrDo7a5zqws1WnudqG6BI5dnRK3ryWHYoOhHXfunLhQ4/diX09
JxvJXVnOHtKq64GtdmfozOOFSbPAVLZ7viln4o6kfrffbkV3Qql2gLJBDDBghaT4
qSMIBpe2FuJGqa7V3thOHkUH3FtIKRzuz4hEOCPJuuw1rQnwdmU8sQDvI//xpC1y
MWTMyxr22K667YcXDYeGR0pvb3vxLIK811tHUbJcxc6Y3XXlvOAV1FPnFQ8BpLr7
e436zQ/opaRdZq0q67u2rCHqFQ5f2syXZBKQ4vip3NB8L3+ElFdliFOJPXDHU6QC
GGy9MM2jCb0c0SjYYtuZhcW9L0NufYZEx0eRfsEvtLTdasfOQN9artv3sjHigreh
WEJimBKkUh8adYrS5D7VVM0GCi/a+bVukumuZ1SK/JS1YsAAObQrN7SzZYnII8mm
IGAQ6xvzMPKLmcWZnVhnc7RqjddMhE5jC7vvebe3o2SMXm0U/vfVBQY51BTyPwFp
a2q67aMejxyNOLbw9Er4tqp0lSt4T/+ocv1ClLo96HUv0Q/yNxHd7fl2BRspeMC9
c85mHq/xIpGLrusZKVbuCiKj8B4m+o3VdB9jR1AatR4HmFMY/0/JIflLRF7rlf3/
Cdj1YwzZAR+kCEaij9N2qBYRtYFmuWS733ghyVzl8/RctgzwsBmETcKPYIaEMK7V
GRye8Ht/tSLVqf25uIXRcfNtAZZDgLcaEJGBhtyTApywgafocIyQkzYwtPNMdSLz
YHDz07J3BSTvcGKHy6xREkq9h7KAj1mpSz8kBIDokMbdhvc3uIcZj1gKv3L5hI8v
OMGnZLSnPT3Xc0Gi5S7PHazHjh5C3MmKCBtvQlrHlzD0HkTO6icTPvI3xzb3zU5w
w/bDMWqDHvQ8X12deZSis90S9uB9jseB0wCiP6KuSFJR87vrn0R4x7foABc/Ial/
2Lk6M+bITvHvb1wURVd1+Z1eSfm2DXTzQEA5dVkDE/qmoyJAnFtY7yeEBd19JQAC
NCy/5WiU0dGzAcjnmPQLf298EbXUZ/Ses91rcCqj3nu6D3s4qxw0ikuN90IgwU/N
O7UCP4XUXQw13YIpoUW60RrBO07QQ7x7iDjD+VE9PVdNIY/goaR4PMCompdGUCAo
wGdtWYTdZ6DhCpqA8HWZXGAv2JYhgHNDtuL8rooAz+nSaTv9PbHjYO0MfpEQB8wR
+rpsdwcF3PXWGezgD0CxSocrs2El4aJUUL9/CCDW0XRXXzgJamVV9sZSHJSxHDhX
SB1JOn5MQ7DwYxp8Otq8bidpKfuH0fYeHPzg1ET2VXYOGzN50gftZrdi0HdhouGr
m3zVnS5ZnBUHwgU6cumoLbGlnl5dZ0QuRVFDwjfhSAMqP0fMyHWoRwku5mv9ruto
ZMiUp1GhRVCUkhpYWNBM3YqKqCvaoVYXVnLWzPqlYmTXHDCDNRO5I9xE8tnZV9WX
6WpCwuz9x9IwCyev2WwdB5HLZB//bclrDDW9jZsnVY/qbJ+AAWpuObjL8qQ5D2o2
3X8t+UaNtGOKag1VpWXf+1vKP4dRwXbrTYwA3dLm7fgh10cSIiAwtj4j0cd7rPET
NU2IBKR5RNr7AKZ/g4tBzHLcS+/0yk+AZCeBPLgkmLDo2plo1CgUaSz5iTHk+RT5
u1Kgm05PGIpy6sreXZ2iZzlKeJRBLb2hPY6ERzLYUl1BJNvVKLX5zQhd7s03JMuY
HU8Dbrn1U+56havKlvGG69X0xPP6igp1Hks7ShhTMH4Z1tXd3dznLTGACDEvMMBq
npUWQ0n2k1FlsZ/OgrIRTL1mQbkyPqq6F20BHBlf6q3rZ8idCKdFs5OcYf3Rpy+K
mKNjAEGPMf4ioRilvdWyppV6u0RBR2hn+lLdxFTPukvzOfV1sUpRuhj1nlwS0k1y
kNdw+U3U6v0bxnOrsT4B2kQW0nGoCTlFjNRxX/bOuRTfJ6+Dwkn/kpLt6DFXE8Go
D6PkLUudsVYTiV/gJuYAgpxWXqO7DlFwssI9tYIdweNAn5Ji7PfU7ot1Ixfgb+ss
HOMsH+TqG7uFvs8nmBER07013J3UFut0X8xu2xnUrD/JOmOGR6S1ot0dauOyI/Xh
ycpkk1IviY/x0oU63gKcLLQHJzA7OmqpIb5c8Q0fxd0DvGjyMSrth3Kil/doFQve
mFd6Iivyyy1v9+xpqZoR/X5pUGq1EK0wlFf/1D8KLHk0TlyGbPebbgFuEtzBmeBs
idoCgDUAE43skJWgcXkbgyooax4yE15zreUFRMnvTFb3DInuSNFS698CZqOp747c
EovbO0K843Fv+StkLsX/K98DA41eLpg+GeydTuNZSPGMfMm1D4c1AvQV5LdZvhw1
IwLFIrrKQtqGOYwo9CpF65qeJrPtsoymD3gW42+zoDz25q2OCgYkeDoq26+NconX
CMbq6p77p8rOaVHGMdCvDm2c3Iq5+rjMm6RCb0Kgqc+AGMO4mszA7kx2mYF5lw/1
ORBifCrvM6bvb0tJknEcHoCiIe/+aOS3dP5fpv9O1ZiGm1yOESRZN9C7HxD/Z/Pu
R6h6Nv90+0yrKnA+8N4jSfnMUVvYEBjpyXfTsRie7YDZceGPReqkkL1VcVbr+a3B
nMq0Q0TxrpXb8erU3gUTF0iMWr9Dj5LL5KI9KVFe7MHCHEdsOoBwiphvlRTNjtH9
uowDGkWxOR0uPEdp+2EjRvoiiyEwGnAdY45KUL8T1UVRI/2o5xhpqDOuEqiii3iR
dcbZjeMzWJ5oDDTswWJFRuKK7kxhJkcac06b0TIoOr31LRimCcau085pIAyblYQ0
b2kskL058AA+HJi3LA8W116QHTmUB1YBNAO1kh7VXEfBTtvmb2KSFqU3KlEcm2kO
6XsoOqabToqoDMCx8D9yvxHdWIyEdbdt9ewN9BiHuF6khb+oRHUbc/xB7tSxENoa
8DOpmhbW/4p7g1BKwblI3sBk6pfF7HFHIKEVRMkgWvKuYI7N9ubDap1VCin9W0z1
mtyYula/byGaMs53ibQ7gqvGKP6g/KBf04H/1kbxoJakBXWL6NDvGfujnDTCcGSQ
hhfLJ62Wtx5VeLEBrQvaD8W/hBirK99JffkNNMKc/6oYzusp6DTtKCtLVBPJJvs7
XDDLseu+UApWdrUXcpR3TauXiujHUXlhzHwqsrnlJD/kO+uoMTAADfXWrlYuxrsG
YxZZzHkbmE4d/g0iLdQkmVgaSsCDn6pv40AeRTzU8B0+Rl6LcuHZnxLPnji0EqPD
ilm2or7/nvdhySs80xk213BbKHjopQk5STjAUjJfoXajQrWFqh1AMCtyRNbwxsEx
GxzMuWPE5Kwv9MWGwafvjdvau+Mcl3GRV5BflAeilxqueQbVQ5J5RaCQ4KzqV08a
+GX8HRA9QWIcDaKhX8klRfNSQDdoR+95LLAh9yApzo8g3xHhyNDpbxiVxg9cU5kl
93a8eAjplnJpOH5NPsQ646D5ppT/qaBtWhQp9jk+7m0/2VcX1YaESQEZlBtI7+Ua
s3kkAMH3AsAfRTLU4yA1egLMcJKf8er+nNvS6t8l0T4R5ZMU0S623Hp9Y2F+kciz
pWSeQT2WsEJbdTqWiv5zeKmI0vgtrAsxtHUTtytokk87mjAbXQxWNXiPeVf1g0si
j1ybK/eRGzlk+xvUNoZ7LrX6R9ghZzWwwM/+A73g1LS4qAnDd7OqlEfRv6Fxlxu4
J6YHLafNRm/eA3jzr8VWsh8d3KK08oP9kjS3jMG8CgW/LgwZ0w6FwJ0iCT6VT3tS
lbROUsYyZcdhwGMdNYxG9W4+1wBfvMIlMAgkqiGImp6wFXuRFdR0uGL410HG19Mr
Cu1AXNEfgPspaQp25HHaOZvXghy851vtkCwb3QyAIuL7KTSbOZcyQfgPW6AuIfAX
3c6RQZCnV2L5iQUAZgGt5rKWyDRoUDwDpYDpCfzAqzpfCWXRTX+5WqrDqb4ynnVT
G3RI4OFBulg/Scr8Lr/ebkAT4WFxDTSw0FMz4Cz/jASB5vzNaImqVCvyvC/8O30d
75U+mF1yWaFXZO7pTbZMHcpyVPIjIfQopaCgz8v0ngL83uh2q3FomffPM0PtF9qx
2ZM0F1C2qZkpNRaxLpTI2qBu3vygHn+Lsr8X/U4nv6ts1CZplLwMXDkRSuxOZyDD
0TiraDnfslNfIWxqFGRvAvEf1O2ezHsNaXQKNs4meX4+5FWiQ1su5azuiQFIR6OO
Edf1xZ7oyVsvS9VvHeiskRbL2O2bBAPoLWyS0LB1Cf9FbNAXdc3vcJlHknNbijFM
8qubUyDQcWVtTWOWNszU5fI0iUkBi/FaTYucPgXLspcbLGCGivkG6o8KZRIs/TVz
LJ/bLkvKtc8CLghww0pKOa+Hckvs6tfPQC5xqFP7G1uonp6LJMInU8Tdd028Pfd6
D33DEAh1Q5iRPBDJNRbSuo1NbS2znhRoTvtynjnzQsOBcw9OfVro1dGt8+Ozxym+
HjyixoO/mn+yhZonhZT+4ifn1QjScY7La7y6CGbi1j2eci1Gb9K9gbogz+eZltMN
GhOZo/DxSVQMK1MedqX8uJpm2wdxJTTmRxmvwpskW96GLJtAkTYY/P90VrsKEZbs
Duobh2rQmROVFx+K362d7D1Fv+ermn07GFFFkxKjn6ZVnkqG4UIqMUmvMF4MCv5m
9ki/R5/SVJYHrSk2UygyH2anUFqneF9ix93k0yElR6t5VWFn7PR29PlmRFIjOyMz
YbMwAT1mckynAIDfEq2n4s4vazFE1Uw4CA1fPr2kuMKcT7LfFwItRtqCZE5N0SGv
fPlikJRsg/wXq7PTbzvNFkWWlM0a79kyN2PiCXSKVChpKmM5YMIZchVeXwkNUyOS
jh1cc8I1eTAaGRB8v+b7pucvlxongrZoMAF+RBavSPzf4k2PIJFRlG6lfRyh4wBE
akl42tnCluoGhurscv/m1OJrB4ZXSoAOS6aJHWuco+y4WrISGQG8he+UibBxgMVe
jT8KGTwTtceWQgGQO9BU7r4lxrP9p9+/oJ0wJanfuoq17xG3/3R4QXF6RYDMICxO
LjDOcPlqHu9yeI6TheTPIkIxYMuSLJGX2qt1CVdckdQnhAYu0ZL5KGt85V2XqF6S
IU6ew6S7AjR1iLiWMjjwwcckFbzEIMS7vo6nsZzYZe5XXBDMCMH4PduRzytmZxOW
Z205X9PEuOYffTA2hAnpIm45CdeMBnVCeGEsKXj+aCVimUDe8Rm73WtHMr6AKj3n
SSQmiL9Mwq2Zs2b7EuX9vW8hRtEi9pRhgn+i+gShS7gHFAg2vtF3flHqNdHq/N1k
LM2yWrhWf/toXoyOh3+26o6GY2dugq28eH2qzz3mRxqqMDKatCW14R/GSA5xo/eu
eeL40xf7xn7EK+tK2FmMwYEy5UvlmdbvBqwLzFFOd8+/Lg1H669XUdaQ/M8ejTM7
yJ06bZOB3mL1IHw4zOcv99qielVwxUnSEQTwD5I7Pv3tr+zb+5b8SO3CRGvjy/15
8+Zsi82osODvkbvSJbpnv600L+NIj9Xip4wk5UKg8W1CEE7loN0x15dJH/A0lARP
3a/JPj1idp15ajo7j134mOab8G6prnYM27V/k7igfsNGM1B39Cehw1gViN3vp+dQ
Wn5vdLHfyx1WMQBWCTbKoHgEFrE4dzOh6VD3adKNWAB4SCRq5FyHSncWGxcVPoAs
Dj8NJWqB5oCsqxIYk2gKabO3xOs54+dyzAXGLuouC0kVenFPuCcspLlzmytQAwJ0
D2v/GLPlqcWoEUBuv/lgCR/OISGls+ByNRdif3gTj1zTxh2A3OuTF4ReuGrDdut9
zwqgyP+NIc/6mM6WLcjPgvSbzAajeaog8xuaiBUEyCpGdynih40t3elukdnS2CXd
letBQJvH5COQVU3ADTNw5tR8cNlqMD29OZZgsl/f3D0gcHB2DYwo0IZJUERD4q3A
Nog+gRMOgY7x84RQibTsxIxWoyZTIlUVIVuNSXHbkTn19EfySH0wNYi6rNh2aAJI
pBhsIZoaqFdIarixOt4l7cq5ZXzubNjBXwquV0WRxIrBLh32yTQUspiq6LMM2e46
u+Jo91D6sGRLjH/8B34+8tKfsNKwrEKI16C0wIWzrxxSBK2OcfnIEH956IH+LMb7
wr9rSGrf4c2vo8MfFV7jI3rv/obFQxu8pzkyuBbtx4H2WBQr1yQXSJ4rsk04dnmV
ZQ+z3L5uW00xQuZS/YhQTwqxuDwBVpkQarCKxR+JQtTcraBhZ/WXCBEvYcTap/kX
KHTXfuRdxmkPsRbwSKow2FO60AWacpukQDrgkeO0OWcbMW0AaCjr8CfCbU/UHHPx
FApMuxqcoZwGPW5gt+nQKtNBdheTajSKBBSl9RGCnoJpXRf7em7qXJtOcinecunb
HsIFLnC47AkQ7neOeRdizLs6NiP05Di2J3opXkJsuDZtM9K14BOxKmSVc48sP+fd
DvGrgnCzl4J/It8gj+PqPZUknVnL3H7ZNtJGXXnpUdkbmzFcsD0VxP6+e+gPsGYE
BZTRuwUeoeEyXBz7v46IxBuDHnm2gYVxzY4wFfq92PYnCxqa7U0zbXAFX6HDBU33
sQFX1EilUNUZqzFVKY57RIj6m1L5XZUN7POTaK3kG53NeFL5eOdt64EP2ac5jDEe
tAqxw5rlxOwO24xdhEZnO3Sr3igjU2LKYGdjoHzgrTHzpwL4jkhkNezksq3wxraG
eED8Y2AN9TRfazFzZ3IX7RwWjbpLNaaDd64cAcXibeTefD/0urijxMhuPrFPphfh
+ZGDM3YfRWLXfPl4QC4fwbp+VRWj4/J4oTzmejOThfH4j0LZaahuKa7mKNNHA0kw
qCwm97Jy0uHZZxOQTIwt3XJiRbMixMCgLZd5BOJaLU3Hd+ex/3PAqys4cAsVZsQP
B0RjTPY5BjOFIi2URjuR2+Rc2L1uaVvpH4PmQhLPfQdYHVwDVbcskRTm7kwgTQNa
OJ/0Xy0OxNAhfJ18CKnOOMilkrNHV4dRiFLze2SYoKfnxSAgr9SdC8l6xrBkIVLM
lzK0rCivO7qHMhYu9qboGE+LyB+C6U5hj/gkYBt2Nu1wLcB9OOvLE0/MsfLP8M2l
osGcVjFFMaYGmbd7wVB2nrmpKZp/zTagmHRBDgi7TPSdk0V2emqY5/+anx6vmlP1
ToGfnwMrL1EHvEEdqtgFKgRY5TV18kxdAGKwi4LH/CoezwoCyIbP8x2iMgGWYNAz
Ff6+idMJnuZapUFkZu7lz/MXIi4DbS5Ip8nE4Ve0HSEEuVjkwRbBHdhpZGM/+A7G
T7DKr9nY0zKPJLfKiRhGIc4ychxyp24vZnOtvzTKV+ow3F9dmzb26Tfyj7DY3PfG
bRcG1r0MCoLsizh9g+HnjGeSn/QL8POuhYZUHSiil6gIVcJTw3eWNJpyeNQvqebH
nq9KsPcecgLhiC3U4ScezL2b8zGxdMH6Ry25i+BFCHQ4L8aUsO30nT9UtAZCt3wZ
g7LSAkNXQy8GW9xQwF7EJkjNTTf7/ZVstD8sWUU9tQuYilJHwDtrfUy7v023JUNQ
iqKHjVJrSWK1dDZViJGa07ndx7mQ9clQbam1o4YREtwdoF4UQmrYqHB4IZXOIJbV
mX05vkkvu1r31zwH8ezqbQzkcRNcztXKnofd5IU5GbVuD9++pxxlU/k/xAYUCExg
nN0lxVoAW4hAWSIx87/4GPzMN1+z0RTxmhx3uiD4Mtd1Arh2CFgjZ3o1+pmyllO8
1SxEArNgU36G+EbrZoenkCQoeKIuAcY58XvsZLnJKMIDAXRW24N5VKyrmFn2B/zp
U5hA8bgWP1ckTphdcwYvbtI8ioxdjyDaf3yBjFXP2VMGm+/Tc1XI6eYGT1p8KhRm
1bBRXaAqIjN3o+cwX1NcTXWldF9YPhD8vSeUJXmDVU03v9R+VfemySYBWRVtErkH
aOj6t6E8MmWizpTjI258TRGqBw717IEaZKP4T28X/+PIJAfZN5xqIydA3HrnV0Ir
cQDoK/8oZUg25wTX1fyGnylEOKjScWZSdVkWwjiVLRObxOAPeML6MFeKVZgQuYv8
Qi5qiZJVUj41PLDoaAuBgi1VPJK8uw8zK1czQ/9j8iQNuBjgu5bPUbScq9VsZns4
sZADGRynvKqXo100rJC8F2NtkRlAU+kV5iyc3ygsjVCmtB57iA+nW0ut8VYbg0Di
Pcw9ztH/usL2bqBHnpVkxTKyVCulK3nppUT97qQYsdG+WkIQTYY4X3wiOBRe9Qmw
DNgdX9eiSQFxxKjMYhx15LSOtpanVlrqq/1Fu+E/oDSJqW/23J4CoQIscMBdXGIl
3TO2AntbNgsAw9cgviMHGfEZNrVXDG6l+pymP0CUzlEUxk3IwSiS6PmDnOMACUmC
yRBFNLj873mZzlwuuphKRKv+iVcxeK9t1YCw+oaKBnAMC5aWwSHwFO4D53c4/ptt
P74KXNXVagIVe9bHv6mujS1qgb9h4RiaBkRI2NIqWQmE5QYQSAgsi5zbU4xy/H/l
fDqM7JKsSrxRcASezTvtQ/7vwuMoqs0wNCPwu7srlhkEXzaALN3M8h6kddQaNTmx
nTbIQTxuuMAEu+TYNlhYO8rHjm/rYAzYFtxYQ17d+Uyysn6jNpftEmllHpqHXaCl
5S3Yvgy0sBxZ2kszOr7RfjIDt9rxgh7Pe4ShYPDg4gPKPbbT3szdg5SdydV+u3X8
Erx9RV3onY9P2p90cU4f599qNbA7TWzu6kBsRRPTCdWWKeUOOIdC7oWEd4R+IpoF
Vng+HILcinl4voQk7Yi2upxyTns++BbxRDmK3R9ZjrOQeDcQZKedojFeuiiYlX3l
gvC4lrbiN/nZMqzmAvSJhd5HUUsc52M/Dtn4nlEOy+y3sr5tQ+w2+dzx2QD9L7bR
8ZlbL+tDNU+FwkehlBQhW9ajqCi7EAqB3cCZ7hZjiCh9N1ow5N+lhQw0dUA96AhU
AaUnHgqbVkmV/hZHUbMWdS19KKs/iXXHqsRoiBuW4SGlGj5M2A5Eao4RQ8e6b9Ty
aWokP+YN3vtHNStG63L3QCYAh1YiQq9vFFRm4TFd6E2XfOp2IEA5Od88/Z6OXN3F
0q8WpfWr0EdDrfkG7fvUml3TyGtzPNaJEO11zOlgwY+2CbB3mNqX+oUDWa8j5TCW
4rfl6yrj604otoQtb2OlaAXgPrD40dEfpBQDXIKDLHOjH5ZlluWXZY0LuPyhfEK/
4XlqzRXhQ3EJ6ro0kGikZScjQtMuR1adNL22vz9w/7e35hWwjMUebbEjXpqXW3Rb
4qMg6cU8dQSNIed9ACt4+Q7Q1eImdC19Gzm4BfGCVGDfZMzT/a2QX8ZNLxZtLwXb
Cc2Abt4lDTbd1abLV1Q51gjDr1qWtrDx+1ZdSG8BNmX/n0r/by/mtn84mSvYug09
s6VOexfZe5fyk1ea86vgHX96Lt5tgCTXaLS+xJO55VT80BXRYr6aiEnWMA/mUwd3
ATkjxe1NlP759GXelIOSpEsvQ2q9R7frWpzgCLp8kUcWMcsCE73zN3USxnY9QbP2
bJRHEttG5xZQ2g8lUbSYly5Zfh+85N+ggRVVB2nngrM5ESRC6AqiUxqk/7QSf1dO
dMi7H77fFjRl9+dgMNruPFHAeSx/iEaihdxqRSffNOnT8RIu7JUW9XsZKIjb7oWr
xYcrqbjTfYm2+HH9zJnl/35DQEOHYPJv8UBmRedoTaL19ZvDjVWQF7dehgdMflDD
KryDbAeDT4WU3pnwlHDamaE64y6NPKDRIC3B3M3jnf33/KPvpcEwVXazNi89Vm+o
TUC8pLRQ3nYk0voWRupSZl9eEWvXi0ceawjEhonzxknFw5FAPLxb6E3Hf5WEzPI5
IxGmonQLfs1B1gpoAh7C7AJy4t4qTv3+uvLM6VZutWvJL9yMnGINbnVV1mAdpBHc
7PFEE2pr77LITYYhKxRkT5EN93qdpV3rbVwjO7xaR816wI7r5xev9LQSRL36eDLq
2dVTZE+AD2nf4PyzYI6TAU7s9I99OiFowhbwDDNEnT5OCUmYBlG11Y2yZgC+SRn+
k4aygNBBaQJ6XhGzgGYoVD9/DIEFooPBkKTHhZFoZ8qQ/2HKhTkDgw4BR2kuG//K
4pXEUWFeaUU9BtxkXXC0iDU/W/m0gWRq8jUdcKqLnMA1Zj3VpyH4SLj9TEN5c+uF
wD9yn4yW7eYKTgggwXRu4GVFT9oC242vpQqjZZOBJZjKCmkQCZl7tAgN7gVmuOHN
dlf4N4LRDXEjosvGvayKB1HOo11rJmpSqeyozdCfxS6T4Mxj7WpmgkZEzqXbv7DC
wQd+3WKrUsdHz0il00RpTsQ0japDnqCPNZpIcOOXZjTS08gMFJgmITjJNgNneUhb
Fmwnh0/GzW+nD6cOXRlI3M87SsDOTVaPvebNn9EnQXHoQcr/DVkqrQhQJ6Mkuuoh
wVwjKqa9MV93A/iP94XZUXGqbsQ4aJFFajdv1p0y0tFd8VRn0D7ND1zPncrMt9AE
lgDIdWfZfYK/vYzylNXg2XDP2qIAb8JBMJN95tgGGor3xCd6YZPXbnGUmMMjbM6t
g44S/yz/VHwCW62lv91IJzbkpPmK5k1LdzdigwoVU8A9sTUY/seaUxR0+H68kfL2
Pfdks5L+//i3UlfkWt5xP9ZP1JgIEaJvpAoLg1jK6taCMSpXeHfg7gMY64GJ+HGZ
MpvBVEaEaeVW71vPcFx9SOVYzrfVKEi/SaIBWw8qtqxRObMbu2GeLp7/yDXGRkuW
HFl6QgulWQAE+kRspeNm/0NOKr788a8ENoCQ2w7bTeMsVCouTwIebPd8rjws17lB
O3cJpP6PhZXpKqOxBeMlI2Mrn4glY/pP+OiM3iVd6A628IKzUnLPRfh5K8IBQ5qb
ACFjb4d5SJJVsuzbdRajVRvoQGCB64iPPNAl44SwmxiNZ05yWWepaNgJGrhhfGmZ
sfnuLz9Qgt3kjpNa6HbHgWxQPqOZfDldYL+4ZgojJn3zavV1S/RnIvZCPxs3WPlH
exDQih7CghBa/u3b2he2v6v8OljCLx56CgC4HgJHCrG7FawWJAgsCaJ0kJvuV9DI
ntVQEW6AxwShU75hmn6ejnyqn9wcFoB1TfwQwgwy6j049Qpi8J6zVsDCCgYJpSKC
59fzd8IqpJfAvmHz9sEiVmp4cWuUbCQTyaID0/mHkD2M7dZBR7GvTiike9x2n2UN
01NERanlv6O7YAZMK87GF9n9PcJg2FR4RXmOftaMPd4y+lpXL005fxWzFPSGLx4E
BPg3MkGpp1tT2pYyS5gR4I/z6Ik2cGi8IPpUl9ZUUwGNgSMa84rnBK+EXEpcjl9u
+36gvk9X7yhDRigZ0HRR3DLNLn1R2bSLZub4sdw4na8O+k1G6rWQw/BL9QmRPFQB
awDPdLnEpS7WfQlNoL9mAA88rK9DrQYGMf2E5sVfvEbrFAx+9Onhh/Luyl6vbOQ5
TDoD5Tnbjw7nXhmI5KT0q9+jWTBRtEE41mxp5+FK0QCGNVPD2W/WhmwNKxfAjP3C
SESgekXsjbpXSVsAvYmPYG3ShuEnETm+rQ3j1TFrKaYO4mmwhEuDWgWAlSpbIS8C
w9sW5too0bOrpudwVfezwnLK19I1H4xInd9iWaWlaFTg4clZ25MOs+hy+AxWCxs2
3OQYC1gYZO8wtC7CapsS0BTqG/u/0zR1rjJaAR4Phey7NdSzSMP4k6uMF+AOM5XN
jOyLKcA1mvXY+JIw2mw3vn87QZlEaxjTRRwGj3/wlpJ4ZgQK/M7xxqfOr3fhJcG8
qOgSPJOp9fLCjWvCxVcc68xkOcLJL0TxFsdJe/14+hCPY1kLy8EHBW/BJyoZANko
xei2tM4PsHMwWM6NgQjwCKnpy9vcS14toq2iZ+QRG2Hs4QEKceizsmlNz3IuMvXX
c7FcUSk2O4WcIZUp6uOe98PIpAlz6eZWmmQRVTvPEm5c2DDXpUQ89WsTmNZAn2aZ
AgazYX0SSRyo4XMuI9p6xBWr4cO1nvEpXXkf/edPdoTJhfKS9m4bvTgp/+qXLS+Q
sQOAqbdpvD2yVB5Bker7OmSqriS4pDQ16aVZsvZEdm2Btoe0A2rUNFLO2/biPWZR
PGlThPFMB1yUVn5soab5i8crVKV9+UQ1GkmiPYY5jhZsTm0FgA5y2i0soiqVzdUj
/7V5iYvAf3bsnUavIeOynszRdnyJLahYAJln62XNIeP5uoktxAPwWH2/sxuOdCZa
UJWd5KVPglAh9Ai3XxkvxJaON/QoE/GkCIgpQpQz5Abje4cQpSv3kYYEe9I3T34Y
mzEnLhyT/Dub+sUvuTrMVpsmiQszIxgJyicMA2h1vdbKEAQqizpTVDvUAF+1Ufkp
2uAy4fHqEkxVm/RZ325lIlk3ML4D9uEynWyy7bTiER/lIC2VmuZTScwAfRZeNZSl
JpbYC+qHnuuvmUzRI2qPMxX/Y2zbi5M4arOZ3c9YqqlXjVzooShVkk7ksC9jsXoD
uYC3IODth2RnudbItUS3A44CoVyBFVXzByJC/+Vx7ye/l1n25lccGNrKaHeZtISx
VXIEh1TJUz3756zT1g4cHLGSo2C6Vf7sRowoyOJSwKCRNKnJnYEA7N4+hOCpRCDg
uDIcJXD6ealQu5QJw2qe+uhEg7ivBjG+DoE+BX/Q4F4w7CfyoeM+P1RfxV+resCQ
1XLl26rmLsCrOSkhSYesbL17CW6l5PD2cHMbVNxqxYhDCGi5otOW2bybkX3I45k5
xb55wbCQLlTIqZ8ao65kKznSGtf0ilnsXsyqxilUaTfI3qrGJNa/ZP2WG3BR60oR
KNXn6BOpFfCPratutXQvNHBLPtdHvxELPNOkm2kQN39wM0tJLKui7smU72ij1GQ1
oFiWis80ItXnCIPkro/krAm3uRpVyMwqmIPI/houpYRkKnIMWEf1IR6OcKGe1Upm
okfemPK+tCVgFGbfCUhFiLyl0bS4sRk6jO7fHV02X3Q3Q6fLCUMt5WKya64FpRZS
EkgIvE059XKDyBmLncPHmoRoi+CE5Ru79BnAmLaQC7gAFF3oI60rlSfjgzWtW5AG
0hf4zpatziYW+S0VpSYFCZiWwjH5BleF71WN2BV6CHnP6InCiY2DYOoEhqlEKLBD
YYd1pLlmifKo0XavD0DftCR11Qzb+uc3ZCF9lRhKtnXUfRPceQcmRGSMaenNotUI
704zrWFC9EzBKMKy6CYJHFe6tLN+XMeC4zg5dodUS+aKjaWE6BCY/jXv6dtJZ5sk
bhmevZ/p0YRqnth3nb68vj46lgyShhM1yWOz2SJrpF+mAysLDvzZ5LSdTcKa56N1
sfsNV1vPDnPIOZYGzHQEtceG+G3WT8taTBx42YsvmnLdyPHsi8BDRVwaYjUyIIB9
ggSF0dfHaBQFlhgH1l4hNfSGq4XlO8puKm8jud/JghzqKpqO560Q50LHIVU5IIS1
odhsdix9JBjjtMVl0g7aH4iORszgVd7OuCewEIekUPWRhPOnIkwsCuOhxQbG6LD0
OPmvpyrGHVLWQ1LqLhJF2mrW9sdRWlYZcCCorX9zjM57SIT8D93PUmUvw7WrUpvn
PQcUeG0RGZBEnqaMFltfOP9a6SN6JgsraEmMGa3bUpa7q/xzjqttgFmQJXhiqZKc
LvQGap8m0bMeV01YvkyAZUd9W7GNxWIvo5P3WKWmT8qiM5qZd9oI/tDw1btlci+0
tEjwNapk6FkSLKKQolTNpYVo+ZmkxRvpZqy2Ci9B9BrlbEqCl+W1k/9XIaGBMMe9
8gT0tarsPNUsujl5Tu13HYHelSlAkoURFGQXxH+NIrgEks2pLeupsk/bjKLPafoI
eVe1fUQ5AjSQ7Qfg7otChqB2gO7/8oSzBFWn324sSNQAykymTPerhrbN0/Q6pCnI
8+LJO0rUQqYmCSEkzGuYAE9GTnNe+JphOtWQgPKZXytsSeVfa9FF3jIcyYEhOWSL
zb0BCvvM8w9IIGpAFgxVrCzi6zQKYQpLkUzGnWxBdUXpFbzOPnj5cFUsvtzRjnKI
LrFil3S3ktptqr7U0XGMls0+Z/0ykLT7XwAlsKJlvuRlEwXia51eVfdoe7Q/9X2j
NxCVjgyJgItcLFcXvSkdL/OR4O40hKXpZs405PuPcHli83KTUqiRTZVkTn33Le+/
qsBl/atzpztUD296mNYcnqgTpjYnKNl3imA15JgbWR9BBShXZUwlB8qveS3Uy8bl
CN+vTZZT4dtiM0Fiogzg5Kw1ftj4X6N4zg+qB4ExQlpLQF0LGqKfp2vu7R4uXrjI
SSJBhaCdcdX9QKaS7wJSs4fW5g3mB4B/A8RYoRnT4l0TmiN9trs5LCClVWxbP68p
cS5/oZC74UWiMDBtpCqEcW0rdv6K7yDyVsHHYXlv29L8eZJApYroVlrMye8GIqZ8
rnsp1ICf1nHevnznHEpQ2sew3DyfOXtGhwHdm+c2XBzUcAysAFUAJEHq9ixtCVR1
WjmGETva8NeeJhXrQHHY2g9LGboflsRdzXFE9n15JLYpVPi9biE4KS25t5sopXQE
OTCC9EcvOdr6RZMDuvKQGZLbSSfuQGS2JIHhya2ZI3ToUZFX7yiojfYHQmgGFPbJ
P9epGUtlzBzJYkAaAAeqo8p/bIUP2tdAKu2bPEOB89BxCLVA+ZzvLFD/glffKKhY
OnWKnKLyKK94EA6+z8vfM6KHuk4VCHjHMk+HfiEWUlEN7ZrVdNJX4KA+Yjxe5/Bb
E8e9X2Xx4/8uS1CCkjt02906dby2t73+b738uJAEpKMhzqf9N4Qxvttn/uYHwLFR
IefCI1EvWd3JJaPRwDLB8PQmRdYF49YM732FzLTCwn7jLj9Z1phBX0ukCcTtg1mh
DbyP8olDjkOVit7tsHPRVzspz3hOzTJw+1P98JgzdUSRgExZ+hvpo+vklilNSuSe
8lPmaeWIuzvnepv20IyHCqfLAEv39gBeCDLFM3mDT3vEgkbq69ogyKFTd1FeHjTr
kbg/6R/cgITx5ZFD4piOD+SYNLVgNx2g410AFet/lU8lSsRbxHOLR6UN5Go7jSZp
2vikCg0SfyrkaGQ6aVg8b+pxCDfYuE8CTge6duBtelMcYBtQ6pShSuAhJ18G17fa
OIw/1b9MbxArPyxXweEFFGsMsCJCRXGnSiJ2a6qVbURCu82XLkcuag8krUBNruyo
YqaVD80T2/QDYJeUb+9RJC/ZgWb6Hnvr97Cg/Ux/GsikjGIxMY18GrDfQ//R9KJb
8Mq63qQMpBKIcL6KwIK0VAjWdCAXX7kZUsmcRt1ta79Iiw87QEdexvxDhxszZuk6
fdD6XvUOPbLaIJqmhvLB1kFV+GcHSEnbdxtCS2SnJneNXFQJRT890bDk9y+4IQy7
o+5LHR8v3pgPDdnVLtVVHpdvGbNO7mUOVFnu5q9UTWQbqrzuNiHobAiip/KOoh76
Y2HJXdzF+z3CyYjSVe9ecp52zfTwZV+/ET/icBXgEenKn2/HKUalGrIgUXyXYNn0
IWTfN9xBO5Mvc42XA2XXJu33ZCQb50nf5otrZQgzlOGtKEvh2v9fW1kVPKJiLT6P
NU4F/xBGOo1lPgwGXCpcwHywI1y++UryRRcZAaHDHG72p3DDdZR0ksvOp8ZDeKR4
FKuaa+98e/wKg6/O67uAEismxlpCkxhBxmmR7JiA7YMeSZgkOEeSZU22KP63IwRa
2JaVuEufc+/+vJbOjtV3Cdgc5XtNAQZKWzueHZbat+6cOZgrIG5IElIQ4V5ydGtN
HvqIklfPnTZ/gZ+b+2ftYzfTYqAMYUdf2IgJsSbKR7bj9EGqPM7LEfadG4xrbo6f
CxUibnIUAH41jYp/aORJWn7hwW0TuJv+9YcaKA8Ub6j/JhJ/1s3+kwSbyOM1lfSo
Q2TSRkiNvYKZAjffvQruGWvZUZj1ERC0PqYJBSJ3qa6IM50vSpPZr7Vi2CcPusuz
fiTKjH1aP0DQP/fT/3Ic0glfECerALg4BZtuFVViZ0GsOjv2eITe1uX4C9qZs3xA
6vlVktdCzrtyrfvT1TCoKtMZsv041LtyfkC9PReoB7CPdbDb83GZG27lhOdIiF9S
RtxX2UEscfHkY7boBvVB9GZUpfrTjfTXDWQiUpJf8uWA0E1K34TCDC5sfrwVsMUj
S5sVCkqKwA+NLfQAd5XadlnwPE+ZqJct2L1PXgFXbF86/qapiyDCyF0qJwg4Ejwy
6A3nci7kvNCHh8m4kfP1YwWxsjtdDWBQGLIe4zfQd6WoookCxCb7RTCprr6KcnQU
aKu0VHdDWJGN/PNA9Lw36tJ1qSTzVK2/dV8IGzfkM0ONv1ZMGZgOclnKOKKkV4AO
CYA7vwLYNe7A4OdwovOfat5GoaBxUilRcZSoyW96DF76XzGPxqzZZk9G+PoI6USO
p/kIteljObTLhbmJTI5I4cGltIckh7uCd9k5NA7Hhw4C5xxz5xWejPp5TI8zpOM9
wHv1un3CrQYw6yTQ1Cq9MxDtQ9e0RjYAzDOsxAAqg7NR8JvDLWamWbwPBcqMMgwF
gHnj3MvquF7xvO7dJ3DtnC6RrJWVPHmD2O6xbPfvDkK5hQC6uIqDSDUUJTCcnVzQ
loRf/trc4vvz7sUTFP62Rak4dLf3FUC0E8R2e43U1uRKd9dWLOFpxHq3QCx2lb3J
vEc96N1x1yDvlz1tmBOo080RrQSvk2rk9Y9AF0exXS/gpMMoYF0+HgDOuBKDrIrL
prHsqLtqnJIGhoJNv0h4o4ZhGYo4GMc1rYRFt56ZjOK7dD2SGTKJHOSh2nQRIxFM
TXeU8jvIDWkV0C3vjLGxPwKnGjEcqFD9QYapNm+REare6MAXgXb9hdvTGaRLcoF1
noPP+zXhVUHsV29rzPEWrEJ1qw35WR4iyIwx76ZVlm+r/ebZD1WkGXpEWioV6rfb
DSTrUBN6FsFxQx3qAmwwxaNU1EnnJlo/SZb4pFo0u0fnWN65LX6DqKBtaOKQUI57
1pXE68pQmFVlKMZzss2ik505myc7m80W492pnonAlAgrVdMNNze7dzR8KjJhtDRx
cA/KqP7S+ACWjHsHNnBOoPaw1R9WG0Tr1zk+scPgbz4qeYvV9ehPXkzd8BUOQx+3
WOwnvRq3RRQrUI/8Ihnfsxswzo3Oz4XLHMNu6k51J7iiZ2gNK3aKCJrEHBGToDsE
S1H+B3tpmFdjQDbC2Sf2+CUZ67Suf0luWGfh6sGXut7bNghJWBaKCrDh3hsmWjkS
Gkr6MsD58CcJ7juCWAI3sFZG2tZy3XVMBfPr+MlOacfWrpkB/3TxQeZDTACBj/YJ
13U7MPZicLXe/yAkSIaTX56LkiEYQAfBzIjQQ7q+jTZt9ilkwkAMZVhlNyz9J2yX
/i488iPHjMSN57OGhN/tyqN6jgZwZJgwi3DY+3Hh93cH41Cyedq2l8RRIGiIEJ3O
hDCBc7aQ15uLHUhJ/V0Jldh87tWi8zs2XyQS8WOpjtHIdCHCUcWWxRCQ3s8t9cGE
m2RuZzcty6vEzCSPzdlTYazfNkWwfb2xxqdHy/9R+O1uYnbBV4cvDVpe4TA7zMWf
iJ6tXrLMWDalUm0ue0MyKI3a41OJl3w9esXIJcLuBGdWaC1b0DHAnkhd0+47JdK+
28YUZpGiFoD4MKQ4z4zAyfBaFGWv1oyt/KzJPNu8nClfs8tWXjeitgBa7bv7Cqbo
8JkY4bRxRunkDS+f0JxutVhuh/ECo/QouKLvmZ8S+eUY+AmGQ/JU1aVhxkZMtqXq
hp74F4eFuKQzQ36u4HoS4QCy82XtQLwC01C0vL9uiE/iBtygJiQJLqkKbpfZeNqr
ty+Y3REmGHe21PDuL56vZGDcgJZKredxY+9cBQNQ1ME9EnmcRfR8Jzc+b1ApkMMO
iu0Yn68LfUeApRaXB58ZUP9YXpwfYlDHSzNAiJdsnUBeMW7KP6sR+/4+CPbuiI6y
R5YVhpUXUP8eNBgMnI7yy6Jhg76IA+jxJipReAXuKfxsUitKq95CEsCc4UJnZ5V8
a3+CzyfxzFVNZZsZPuJk4TW/NHy6wRjPID/S2QtCWPpbX/un/Urv1i/YcDdNdeVL
zDZIG8vLvPnvU/2cfB0zj0FUtRMOIhHpsSyDKQa3BhSjeQOUgazI3nCy8JE/Z7VZ
APco7QYmatdNB+GFokAXj/DkJdDXamTBWDOzi6ytD/x3gboUMoPlfiLJ4MJ/yhVO
NIvZf8VHFc+x0GhlsqtZuRKoWAhn+M7ZbrbdkaVs4KYC2oo1oJyS4pNyEEmzGPtw
xEP/a/iacST5TVC/KrhaDOLOPaligfZd4Pkm2OJi5E+dGr4V7IjonLw45PncgzJz
FmWQpOfS54FgnuTMd/xIi7wuPancdPN+cgn0ELEGP7jK4BzFZjxPas1Hj2z36GTt
BgM20DAIJxQGyS/iu5ZEs0ml+0oru2GULI1v+XYG7YPFrJj3TB/poPVfdojIHTqc
5BUnmjX1993UU9cf3wUna5XRcpyYRSbgdZmRBboDWZiPjzHqZXxpgqCjkl3kUDsG
IVolrHTOMREID1Me+qv15kzoVHxb5RDcFxO8/MsL9mf6RlisXZWhnw/8gi0Pyqc/
GLdM9KKlJBRyZAHB3cUuDs48s2L0u8eaXOEvmlkF+lqRjOt3fvSAd3ydsfHvocEA
vx2p4ojjfIojfCpYgh7uaBYr0yfDOhixOGLRI0AbKp94XKfPQYmsWdHBOmUxIV9c
5dBGJn92zoDTxWGhk7aL9oebf3vvTtHE2DoV6OTe/3SCbHb8jbC0BZf2RrcDaHtf
I/yonisOq6bhQByydbcTocVhNIoy3j3HR7qPzF8z0RMeaVJKDrFyKdG0UPJnhW/F
Nup5FdDdH5BEHA+1o2KIiexWe09QRVB/xxBGMGNpKPpM5aRmjFmweJ0jQS7m009I
O64vrW8U7j1biKsNKcWP1YkTF81JT7gP6kTM+4lKbxALbR61uXquhYgBbRPtvXy9
Hk7FNwryukUE9qtyp0lPtBIt3bWrtPU0uD0R4HStCCC+sVcV+txzG3GISW2rpzJY
apM3iVHUjV7cEHl3Al1sb7E6GaUR6TOepY2EvmQTOuNBihpgou//pwxJijEblw0f
8iNCI1xwiaOs90BubyubjQiBynyQ0rdKU3U4KtqnNzg3GDoMyudW1YiMs0aZczqS
ch0Ma9IU47dDggkcl18l4xSDDBhija6neL9OrfXh8lVG/ARAgc7fGbRkn1bLPCQM
QFGN0B6SzggW6bOC+E35TUi+iZZ8QsSGpvZC8pgzupTCi4NkrrqugG0gsgrD3eJ7
aR8e6tMMtHWtOLnb/80qBlU6BCK/UEbvjIOLad6hIEdFpepuXxbxljnrKi99l/v9
SgoPjMri4WydhO2lKXaFbD2f8OSH7nwwXZztYMpCfySbpQt4VgYCapwiWhBMQ1GC
NukZpB1HB6RZXPQKPHfwTbHwtKvjLM1+EbuKb0RgYYi+v4ie7o3sLtVzPsVWeYvR
Jloc1iXoeBJC2giNlZtJlUA6ljJO72xzyrLzatylBDh4L16Rzw0AX9SBondE/4D1
IAsZjelVqLLW/7Ce6OCH0IX81GtykC2L6tH92x4ZLC89kON8ecJKTXPa8D9ntjwQ
4wE+bwlOarunTruT86c7vdLJdVOSGIXn5amgO9X5AKe0F34C63A7W9XP1hReGhQ1
GgsrrRGpMDPH+pj78NM1fxuR89pQlSCpOkwvGAmFa/SMMKxPytQVGWxMUEQmVkE5
v/PBcopyQtmOsWIrPAaMXC32a8vPCHjwZ3WboFgJBgLgNp6HXpdcdeHb3VKHga9y
wdKGh8PNeskqJtEYb9xAGCH4g4gC3311xC1y4ukiq+DYOgryz2iftXI/MtBs1M/s
4JmNn8IV9E7giFYN36CLqDFcwdeRrAoXIgpS0dX+NfT+Fa2LFFK1ff2RG9ud8Ywu
a5Y+IY5caJp5j4I02VmW4kewGsLc0MAPxkOzkzhRhIaeUy8BF9znWJMnG0jRNP8e
zDOqJiUDgcDHD0jIPhxw/NUeHfJqevAlojEIXMF13Owc0Efc/g5iWEWYLVjgUbVp
VYsy46r4efZpALla084kfJBY+tFZs8n9AWgLUgfA64/X0s/Z8uAsWe5KVRgG58Ce
RfzSeSbCiNYVG4FbYJIRt4By9Kmddi8ZwK9SABtKLcT+cI5DM1DrlAYL4ByIUPLc
UT/s9FZ5kTwjrbNoFchvi2I1/CDQghXA6vB214Dg8hl28fnjaJaDc8fvrhRMYZIq
xDAwXMsOcb2otImDNl2g4+j3MEweQh/N/X3KFt43KmG3IK1UTlxqPrin4TxQTeHF
YnCK3gb/pLGbZjyYpSAnOD5rib7X0u1KpW9U3NbdXP8hoz8nuZpUtg0eGsILPiu/
VGogiJtXAxp1NJmYDOR3+74vusFqYZAw6QubsYcC0BSd/hOb7Y/RGP8wiACxPNAX
UJTGFSdI6JNg+065VLZtCvtV2ACOIFAaCClXTKfeb/qmps26cmASce30rdSgKCNg
mTyuW2eO4kRA0SKTHec6juXY1lc1gJaMTwMcj4cLBw0fnpJSAxLNfp/Zm4lPNfXd
WR6/XmWrX5Bo87Fx1w6eEFHAfiO1nnQxmnOc3asSKWI+ppZOlZno7iDVRTC65JJv
oiqvPi/fVEbhA70lZTOjdqyFniLdPpJUYyUJJR0Q77sVRLXmJng0o4CkwArybgio
nIfji3AsjacNCBZ1boZ3uw/PWbEH+iO8CMSzxQ8LD7ZST9A3nnytK2vJ8akdT8y9
Z3doCEwUa57vsaOBLapeaH0caV4nD7VUOo3HeOIQGwXKQo1ZT4VspO22deEVFP6m
XAtSbUiGDIXJrKrI13ptmt0qQFQE/sluLQPPfgkzyyqw1z6geRZOXA5yiEvcBZ6m
UilTTgLrptBric4TARGF9EmKusrsHIGP5iV4jYMtVxqQa6mlzRsIDhLi9jJevisp
hThKFGTpPP3SXFyFQqEmfPVE0oeh7SSJ0w2exbd1MNFtKoIcRMKLOUm1o0d+iDKY
GJ6hAWGneZU1sSPUUPf6g03vboR1yXuJ8UBVwaKgJKLAECgeDoLiPAnk7oIw/w7O
NhNJ6kpxyx7h9iL5xCF9qgV1tIM5DlIAFXQsiBJ7lpZ/BlfR87ySpmhHaUrP4e9B
mJnGD9GxweKP/nKYEJVv+Hn9g/PtuF62zROXUG/LUArt7kM9dTE0yrV7ZEAUic49
Wr+rAlZxDAsLRTEemXCfvlEAltcNLicokz3B8cFZRyoNdWCH7Zikc/MEKJwv9EHh
GPAXPxSDOSbOGvpZZ7uZEXNm1DChZtVhHAcMhf3DW3IYLSmGzs7ddv1cDs+mTxy/
aeqQH0iab7sjmjf2rneoy6Nl6jVSfQxTn3Met1k1YDTsX8KdIkcjRQHk2j46ve+W
JCnLLTXQHLBKAc/fSlrpXIOTwwm9n+milrzXdVbAIRpKmgYmUHwVBu92yhzXNWPx
6T5AEx5MnDheO4fueKqqDJLN76xGx7p+kmu08ejoCCJTlhj02tFoXB8ZHgkrvwwN
BH2io1FxzGjKj11txoYtiw0iLVdx97NEAjHCFK5/HiDB3VXbCi/lFPmZ+dwdKtxl
p/rW1yY/87QsmhTu0vg8/+HcgmT7bKBHpnxIAGuu77waQO1KRrTj2XVQVTr+GLFe
xSiaLT3Ifw9/a+Te1ITV/sMVH8i5iaBfl0Y2VE2/rWsTC/PahCoHjUCp3V0xqmTr
lAxe7t1l50dAx2OpEtnZO4OsJAgaWOheAr1N9KE7h1O5tdhU3q5Loi8bA2B4Ohe2
QrBW0iw7AzeW4S1sBkzicCnpIuVIkJt7wvG20aCNFSq8a7vd9oP76vtCKyHVWRQ9
okK+/jGl0gAcL0PP6tXY66j7taIZg2kgtnICbdXF+zbU+Qu5o3gyQVD7iezBSuUv
xLFr6a4hH+tFNM+MSz65gtnfq6Iwe2S75dfoNXk47bJeSlaAqa/m0kZ57UGrVYD4
aZ0u0xHGth0Skqyw/58Igw6F66WlwP1ZPt0OezMlhHeVRAES8dq4K68x7kiMPxrv
JyQGKMP7Km/D1+T/uWe+//meRkLLBRddL3EBH2+Fh+e9FZoUfx4pDMIGY7G+RwA2
2b1YkxmA6jtYXbWRVqExhZUFoWXIOKCowRZ5gXowF2wHWVWL4ZaqY84MEzvoXW0e
teFMtBWykGxH4PzB34CLUpYgQk6LTDbJW75L0YWwcXSlBQUZ/xqsaMgzrWU+i4Y3
axYEHqsFke6ke31ZR1r1TSVdiC9ghVNOuvQ87cHemUEoJ814h3cxcelSComNVc7A
v5m5N+WDAZ08ajWGSt39jmafAs388ePcPuB7RpAGW8f7Pmv9gsr62f6aM/+zwO0A
bpfXengyYunwexrI9LNAUaf2axbiToIpETGZpB5/PokqTmqLQOfGAuRi+IHVBm/N
DxiYiIoMj1Zg5HITy2rYYUxVWdcViB+vdmd8Q/yvlVHecu/3ncSU3OgyqoLRnRSR
AQ2lxefJqRcy2MSUk7Y7JSzg1GClbGjYRjOYU6DRCgRiIjuCP5tEHY0j0rKkuWTC
Y2uR7d/JAFG+i63PxTcunFjtmOunX1FzpfPXyF/XZ7RPdyb7SyhTu3mn/yn+houl
g4e20ABrENs90s3X8d4yWQIQ3wdPKiAG5c9srLxZLAEuV2YRcwShP+cr1WW11lNS
Vby6tNXZXDyoPqwxJNi2B0mhWqZusBj7PrgqB0EkGCkR+ICeIgJH7Tq5y8Lvrfee
+RaDg4eJ2WxBENo/I4Vi47HW3kXD4hv+k6ZKjGG00Fb3aiK5+nTM0eMgwRZKd51K
YUtbrVYGZCuIozcwlonujtof15U5kgpgTyS6WMg+btN4CRTMXaxZqi2h6iLk8Irq
oAd1YmxSM/tUXQuAXm3xFUnLOsusySaoCegEMV7MiwqmtUCbyZ9+m5kEFjPX0aA4
zJPV93ws99UPBpi0ybfQQUTYa/XGl/9P+tDd8xviOy1NZUn+wy0o8xuxn1boE5Dg
U+gDIsXUymTAiuUfxK/o3ch2+nNrmQvMMlUuQC3c01eNUcazlb17X5SAXM5wHaO6
Jn6Y3/bjVgkbCAq4Ct4XkEszXpZSfOhiQmQWNvASl2WvnneaC3oNpb9QybtaE/tz
4P2chgqggnHp75h5kZQuk5GC0V80BGwvv5l/lZrIXO0VDDQ54QqZ2zlhsShsyazR
bc6QoHlDQzJUMDli2QkrYWRBFOpzy/gom7QWgY7cMOfKnX5ahBtmYMY6M7/wSqp0
KNlmdhD3Bek67vkqXKj62ys1sthMkGA3WMllO3TeJAm0SFTLGytQP6SfTVQQ+1e0
exzjZIItsUTJq+igJQI3ARmcM3S8ald+ABKvroTUlsLHuWU4FFiqSSS7/wYeIexM
042GZ7QtkP/IhUogJO7Mc2N4HJUjtNM1nQ3sUK6I6zbFUs9+BTH1VpSyHIpyATPX
MDylP0CQAWzGVigrTj3IeGL1nByxdR8T6vpFF5rbFKeZmhktFOtGU9mqDuU8D7xa
IQwmEXAzBV0nXEiglObaGJ4gNY7cvP29DxLWWk3g8NkIM9sPvzlrEsfiHK5tS6EI
DvJ/cVrYYgSY5Tf6iyLdJhbSNXffrZDZ9pcnrL++hYIdHPZpfWzr3nXqTIDx7YY1
RoJslvvK0CpaHh6/ISjaR70xCGW94PCViDayfrg1kv5xOTy/aO0jIh5lJ5oBQPrZ
lsu7Yeb/obPspH4TgyHugRyJ93wy39cvm0wXV4T2yrAWFAl3wZxRYwyTeayMoWUv
MJXwtGCKsRg/Dzi0pkt22y7mDUKHoyJb2tEMvWKVLFwboaiF6VjvcMfd7hy48bJa
SkTa94AJ3ingNfocnRb752jeDQG67kw86sRAGFExlAotg08bERO3sydbtwhCbFQg
GjADqjLgivTSznHpqPD2n49mdp3lJHHMpPqnw7Mm8MYTtE+gcROs0awJ7nm3g/pe
OFfZmqJytn+Rs7kjZn/FIOxgGa4Z8dAkk4SQij77MwQg7EytQya1A4079E0QD5BP
0isa5PLOJ1gwDG9pNjugxxEr/E7OCnvEJfdB2vlb0lT7zYd+wNp31Y3JhN6VuvNC
DELZSnhlf50wBWzjlGInrDguv03S1jFRyOnzRlgoakKfDO9yt45gnWU8PlmWYJb+
anQ9Sdn1HuYvBneOKHUIeXT9Wd+hxKXGNvXpE+iT6K6bIlPddx5cB1x9DgNjyNmb
AP+mCmxQOIqHDOzftZixIosBdT/p4I7Vr6xKAikqx97t/qDZCD7hu/U+Rc9To0FI
kCHPBMysv041auatFBM7bUsReDWQ0tRIoQIWaHDq7CfnMEPXyXeDGWPERULoys6V
148stjQkFx9jLVPmp0pk0TkXkYVsvS/tcM4tlVkhHqRaDBvO4scCZ+vV+ftsmTnB
UI+aC8UaI6gkHAAflItBrbH7l65XOBu0C3NO5fZq8Iw4D9cSG9QXKdIBIOIk6NC9
gsBugdVM6uJJ4CVXOZWgDn3LI3aZyScCSifLMVC0ozHtdrJprD4c35N62CnPCt8B
K6N8Fqi5aqmXPzOqLWsdog3g0Setw3cIQUVgfMCLZFL1egqk35AnegOqUcLBPAbZ
7EgHkA4MZT7Nl9WlftDl5jfGkFpkyjU/73/gM0mm3hFI3pKl1GxavhpzaFcC/zf9
Yll1iwYjR/2e0XuB3XP9y6pGKGQec0lIC1ugSF/L74UYywWgtAKUmCVP5Nm3RT7O
j4WtH+1usILePGQX/IXf8UIkyR/nc5OTOmTlUwN5gDi+dillEGSt7/NspRa2tKpf
7p/mqQoGPp0noCwKh9ucug/LHDeZoI90Xd1DRNKJVUdMEO1EFJ5ULXkgFhbE3BGi
ns+AdwyvrIRReR/UCLxDjjYc88wG5DBqHSMIYfSCdKKeWmQxVQ/P+l0Ew4VzjSWg
9Sw7VAlLyB/xlA58xnX4X4LW8zuiTiJrgjj7z03nMQo9nKVfeDLgsn0ojz5MmIuG
DVzXXIPSF0dO/xcfOEQOMb6546fOA8c/9AA94D9pwdy6XMl8MT6luWcVC/hb9Gc5
eIHqC1rOuXaEdoo9fPEjzZ3tEMgPVY/SCnPDhaf3jbLC9l3cGrbncyItWBFfD6YZ
+/k79spVqlP6nYDozwfwXOFroQajCoLDIz9INhnJ7sig4Da9A9d12G/iYxMhrAK2
7Q53UIyaCyNDGEUbU9oeVc8gzSiUixnQTppe7wM73yijJ6zdkxyV0V9001/tkfRb
SouVk6h95gXACukVFCtyVAyz/NfJ7jC3J/beGnhFm5d2IhLtHmD5EH5ZgVWFAxs2
0ogVas2NtY2Mf0NzRjJ/fN7YAL+A9DnFjI9K/lew/mDQa+9q/nf4j4p9n6r6ie+h
1E+zbiRYV01XMVs0m+YLb+Atx9s9qXXDSZcCSWrjpA3vJYCimiq3PUxcsq3Oi9p5
+jbcSSwcQ6Wv7joOIJvYLIw1hSBFnsLSw0845kJP4M8ewJL/XMlkdWqljfn7TDzz
KrhI81LjQVmWmThud0rUgena9xIJp0LFnKxQ7t1r+ejW/XZrcCmhhkrMMhZsDAyb
FxJyCBd/X8ndbrE7o1O2hr8W5xEg09R33Ki656j4C9zsNVYm2hHP8ihsK8+YBWkj
3SLtnL+C9bNvKtJfHSiPd0t7WPzSF+Nptgu9cR5jZvx0UnHPZgLBYmw1p4j0YyAy
4uVsAMk5JKbbKbzzr7YjBnLYK3ns1QgOrfufR+YFS2fkh87R6Xv2Gf7+hVloFTqF
BIWKMTplkPyq6rVrhKu8BTRhLCQ6jG0IYWOpoQlltPVUZc7dHJddlOLhvflIo9zQ
Oqte8mRAJSTxFsi4fIINbPKpbzo3/w+07hkZWnJAMHQE3nVPiKx/uGPEK0OzM1Aq
oz47UqyNXzGEiZLM8hpQyWAU7OQL91X8D1c7cEY/EUnJ+Uc6VxZUThC7Eb952kms
vUuz2kk60zy8cR3Lzc3h+QxXWmWmxGQmejBmNe+AZv6oBbSQOVJdiw7lmrJGgrfA
Vj7WQe9gPCaE7AeRZ7yrjVJQRWuggmJa5jSlj100aS7aj1G6lVpXUXdYcjTNRgtY
tTiVhXAEHnzEWwsirvzi/ltNOy5elL2U4IJEknOuT0jjCFaTKiN/qVEsvFmbHxo2
5WFRD90VtS8H1yTUhuD/WZMZ9K7gl2+31eTkrCkpOKiAihNUEhb9A5cjwUx9Mgwr
YIZVJD/Mgwx4CPugfs1m2dVoAOhD7JK+kjIX68ozRonHqAzmq334dUDTbH1YAG+l
D6IOXVz+KbqbIP2EdaXY1/N07lbMgnuybSlhPosKNg2lsE9CHUre7Oi0j4RRT3yG
9omMpBHCbdPbwOZyOMEPTt8Lo3pnvDFIi2V3+HXO/Bt9IVJoZuccqeeoIqbQyeaY
29S/4AgcepX8+yanPgc4wYD+Ch8VzFRz6IX+M+YzLXSYO2x43SpCEOpiciUScm7S
DyKoaSzAaMybVTT9lWGvP3g9f+9mwZCnnidJN3oZY0XZOyGPGPLj1hyva/dLGKVh
sAYYIGGwD+D71W0bXbnFw4OJjRW/IlkEJlysVPWmHeFca3LEfWqItScDjyukbar3
/+QtFeKjlPw8jZFWyE1zI4djJF+tCeOm+2xPEZPUMLh9EFlRIiY7X7pwsyxCpm9C
hxbLQcYOZiNhutcrgu8Qn4WAmeb2rRrgPMFRyURPqKTTj+aptzMX1ivof8MO5zUb
PJvnk4YGLyEvbeHpusH2VbvpnrNNBsNFLHbsyL+Zbn+vZ5I2LQkLB1/QeM+4fCt4
9tyF177UGiPuzJ7QDaY2ix/Sq2Sn/2ZGEYdbZWPndHYWaParRZCaadLSaTzVrfOb
7URD51OG4hxps97wDeMn3+15tupNBNqgoiv1BD8G2biLUT+fF0KrOgxA+02AqwSV
Po+XWJbbFaEbEZsMGsYk+1WTedttLw8xOAh8KrWsbxLSrEC1N5rRoaJoSKyYhOz9
XcQQ6F5LiyK8jwEjcGhD4eEyoLgXbWvVnbF3yqXUtjdQi9nja8nDjInH8Ao8nQx/
npQoIXBBeR+g1nzbg3CvyO63Ae3F1Q4dLEmd2V0UgRQWTGOczOu01r6YGxs0tPG6
o0KAmIHS59hDfX/pLvQd8CGhCSDBsGBrRQTeccwbQxySIqQ9NJzAgF+Ri9qCkSYi
QC6EkMdCpi1yO1A8ev3pKZcOmAcyvXoK+6vK+Qn5ldNEnxpeZuw8CD5/YTmCbewA
SPQ6UaGTppHws3ze84Uc58nB9EjgWDR8eA2t553GZkoSbor13AVkzXRZ9yJ6qnvm
sam3BVZRHyV09buu+PnMWW+OyCQJEcQTfGKnhaic4XI9Oale3lM6Cbahci2fyUHn
tGfHH6ZMWZ7aymyr1sZ/GfSj23vHCvUcRwWXqfxQaRrv8EkToiBVWCGkqAIlt5Uo
gy56525uuLeOo1yJvPWTwkCFdsudrQ9/0g7p2SffSHM420gy85Be2+pF6o7F42B6
1xnkrk4jyP85EsCk95+g3nBukqybY6hs0oM7IEx2ZBpB60Y0nnjhWEJKQl4bZRIK
YXW14kzhjYnVEbqq6z3MjoR7OotImRELcLdXBBo5OEg4oxZfA1tQxLOi87NapDdK
aypilsOk6vmEsyfXKI6EMQlA576jzStkgs5KakhJbvJd8/mT0X1WKSmoYE90oxyu
ILkXgO8Sg1l8jCoHqzyYJz2HtQjUgog6AN2zwSLHrcpLMIM58cQyvDkklhBteT/D
NMdoVHXT8ScEZiQgfF+xyFJGAZvxCUgkkKkxeNr8qJYpMCI6S5S4WxJQyLYnI4y0
e9h+6U10Nqx5u9w94spJvjcWNQfISa+jMaD22GBlVmkK1RCKDEql/V1Kbu8pDQwP
9LJhc32nzvf7l2MNgKvL7LMlmXtgd+G44Pn6P7vJTQrX4qwwzEpGBHEGq+sPZlzG
PnS1i5Pevv4likOrAJYhl/zHpT7A/aONqfQqpAARf2GQCX35qXWKGFvXW5Ply8QI
pjhhBf8QUF3mSUCpwLzZz0bShEoG5k3B+jnjQ0q56R3pk1biFou2Z2MUpJto1mB9
x5yLglUAoguCnKribLZRLmQLcaxrTeuN760HT7YyIaCFqx3JmvBY/K5myacr3xIJ
VrsHXJiGCqmxt5YDrkKNEZMvhrLLZ0OTDQhpqePBicWZQIEiDBXdkVYMBodATVFD
hDDlbCDnFkDWLSLcGgc6ym6Dg1leYex3EHx4xVypsKUmlMzhEd85xxQ9cQ3HEdUF
fNn7DcUwyvslM0EvR67jpZyPPbE4EYKzH58t6kTjHnr0QSzAEC0Lc9DS46GbDiH7
04OUTtBw14sHCm6JG1jB5Oqc/opgUYCv3PQnHtSIHJojm5adjjhVDBZ4xWGs+tUn
WvF8QmSGIweyNT9esUjFaBTlOmxvIWYiFJlQoRaqeMcBjHR7/BOInYzGzys9D9EU
OgN3iCgMU9JAWTR5IUR2Bi6ioFr6B13zD2d2eyV9ghwvctqHv2Rh4LEaPFF3Jy/C
IIW9OEPsNkqrkGqVrsmgKpRTnD+Qkbp/rsjy94q14zboHrw1JjJgFb94h9z+myGe
Q3d+NiivlA6xjMX4R8/2OGw0fwCmfwqeyFG88H53s6BxerhVFJNEwGxEzvOpcA1G
DGTTNly6IuI+b2UoBdPzvZXnFt3U0NKzIRRCwkXrit7NhT/tu5bKYZmc9Da6Ut+W
40iXpbpQk3OMcbzhkVBmV6aZc7tp1ah0FDFykC0tPqaQuF1lWSoc6AYITyaDILKi
pm1wrRVwUwcxRKqXdXApYU/ADmk1Dg2odZU/99dsTUqN5Pmeyi2Oj5ucNLBBGCv/
W+6Hm3IhFkVAiB+jbDMxYh8Mo0bPUWXUxoet3cuGX3bWwMB3k1zcHKw2raE8m/IT
lygMRdXQdleLHw+JXNLXJ6qskvZSIEG26mW6O56D1N9UIrzSyWBAq1WQN+kqXTp4
gPP1XHw3ZLVToEw1LYcNuyW/0mC+N+exvIpfD0iM0msoZW8xJZjkhJf+lwd6FGXE
L+GsVo/5iaP2HEsgMs4K2OfadX5s7LDKv7xs36cpEszvbEdzNlYLSkDaE1GUalgw
i10jhNZWUXVHdOErgD/6WeyQ4gM6J/MS6aA3h3vmwyw8GMUxJk580A5ngbC+ffYD
xUlapm7GiS4yzVbAesR8TtWqeXkQDxv9uCM8Wwz4P+qSr/RdPXWDkdQSZ+pzMJ+K
3SfZi1oWStmnGbz+ITms5g5rj79N3vScY9Zbg47KR+MtE5BZQC3kLC8Ganigkknl
aUtSZDJ7pUI2nRy+vWsqYxyZcJ8xbwR7sDSrn8aMxqdpaxdt4Ynui7G77c4Qesbu
MYMmgPwIkbmn9e4ID+Bz8y479u2/mVqv4wcylt51O7enDliP6wolKWmMIDGnZXZ7
v6o0W8GyZBj10WicVXuHB70u6KF8BkB7VmUS7wlXCZbdLfx9tstDicfGVYdwSPRk
LKIcru3zaz5/rgHvJ27hQxnxj6UGwMfdqp48e5VKkXHuiP4zzMiaQ1MXSYJcis5M
ctQL+QwdnXEw8GeeIeyN77XefKWZeBKpFu+L4HXwHN4hWP3EjXFCSCjzYU/RnPfZ
AFFX5E8gGDQYY/7sBedkYCs2bmjUrmjBcDBVQQigvLBZ5M1qmhaBwoSSUpwFM5WQ
UJWbf1Ntqv2RxlYVCl8wV47/Kcx4nqpRljXBQQWvJ9+QDYAUNZf1v4xrHVSSs/zE
BQDqi1CsR3IrNXhrhBIBgUjRMhguKvDAdRVndcA1paZQyZDq1iSliph3r1JR6nbw
QZKct5cMhm4g/GBhXqH3tSbQxtAS5/2mUqS9OvGhbEmdXijQKIRJ6KDzGSepc1xB
GOmJYWEF+Wkj1AzmL2zqPz0b6LcFQD5gJjfQzGikL9xZTGej09hyHklSMTN5PA9r
zSE3yhN9B0kZ93IPyZqi7F+i/B+dq1zTWm++6c9uHzvZXNtI5XTHNo1w8SWGYFYr
3353N5nd2zOnD2vIW6Dvy6rDS4opEMTL0YCnOo1vsNeYpjV5UKr6BZdVKkpSk5eA
tCZlIkCxZ2gQHAc8TVBt+RNvSPH+o6uBArMaqv4WcLyMPU7D7brkBgTfplHWyMFn
zkqQp3EwBWfVezHorxxogJa9hf1AF6UVpITDp3WlajSIXWHaEp9phCStNT+QVget
2sf4o5VmHuDrJLd4Yy/xcI+XxTHmTcYTobXVBt5esn3t2Ccg183QqOvCH3sqlOO2
5zfyNMKO/rUbMuaVJvs81g153f784bzKaBsWMFve/OUJwWNE4mxSbvn6D0s8dqVT
NTIxyiUdDzRWRORCKtLBf9/C5FKXm+YwuD9oVK3RA2Gfoynyolo7roQxAerYEnF6
AF16r+//ZDLUmXV8X/x4fWdcfh7LsnQK7x8i1V/rcdtgNrwYH5LJU3Uv0oZh7yFo
uQr8vDzvCTN/rLHhLLEfZ8b1vYCIIZM4ZKerzH8OwQkJnSzLpYEAiceYEfg0eIDB
MhGrkeTFRTsju52e+CY5GIchEHcpLOTiu+itOUfwBxCe4m1wIWx9A9+gyEe/qP2j
yrLSTExVsEMRfu2w2z1OPTENDVRkvUF0AKksf1IzHBvQ+ciI7a58VRcsm/zbybvj
3NNVaNk6778+623WBunBZKvomBAR9dZasjyM4UxYg0GBbU6QBbrgq+OIDK9zh5mR
01qPHEpcWrMAZhIpgJYDa1uNdD3IUpHC6UyPQ8mVjRJmk6P4/KszeaQVqmaMSXIT
RMQtSCXLwUeQY4ChOJGexVYJtYS4uEL4miI8VzIG6aX3acgyBeoRVWWBk/KiUPg8
ydrWSH/tgxqsKsx6HKKuT/VLXeaeWr1xbmLqBEYpdgN7qVTsu4ZfHZewCnLWZQ71
SGi1Vrfb3fMK1qYejXEwVHdHbmgPMZ4Yk0BT0KpURQmBM73Rw+fG5x1aYtT+pmUn
FVm6ZoNSB1iWfSybziWoTZzrnwGkrBtOw3how2SfkNGw3nm4jeq9L9I8DFXB4TIx
c52Q4rQrNiOchodw0dLE0rJ+MdTI/3gJiDQCF59wvolqMz8/iEecdFaF1WhFVB93
3YnQZ/SFVH2gfCsK7XMnTR8D7KWS8VQv4tyewCKuCszhtDqUsHoWwvBV9XNdfQ7u
E59teKOZ5mqak9qyWp8bUqb11zahVxrnfDmmpbHEV8CYSxFuZoNUT6GIgUK3YEPe
rK/d300UHvQZW/GBjyklUBnCRq9+W8QjAuttzlnXSPasavAUHCI68loacy1g9ce6
emvGAyq/rNprodFw6E+P4pEnkauh2YuDhyFzKNC5b/klJ3rGshh2c4W4TDmZJhAS
e+mNPZjZaUmUnv6uNJPyvtIFatTK4FmPXfBVb5ow3zIIv01BO9Aat1FR95mZOFiP
h4Vi0ohzk04IB/XNKSOcZJuuAAwKeyeRUMeO3CcrjqmFt7yqxJnh5BGg9NDnBFQa
d64NzHdxyrej4JoS5/PRa8rf8sUCIfYUGk5pUZfQHWeLL5k0jCa8hBieWy4g6T8S
h5T3UQEOKvmxJ4QlwBHqb0wEqOhjw4buUsv8gKfpa9kpI6Xm6NDMKCeBTpVW8Fwc
K1U1KSrpCeDwkfNEP4zpAiHP1nZFcOA+a9yeRpnGI2C/i+/TpMxUd7UzYcwc3yqC
xpZ7LRzcN99M75SMviuGncAVRYUIqkemuzCGR3XphioY1eXwYzFjk5z3Frm/DBJa
ojZ1w9jAaT5U8dGlUVwG/zKIF6baKmnskGb2l975LIKGXVHSnOheKkZE+Gfsjgz8
50H6buVbUJhvrdyuymItnzbF75c0uO8REVkiSbJXCs5zDx1aQloMxsLtLrro/ejE
Q/o6zm1+7lUv3SU43wmxfMHp++32Fj+o2jS+eL0tQduDRbmL4UBKsV+wWOKp7n7F
k7bxOudO6/XnajNkDGcX+HrNSmFvQt0u7HS9ScFL7W0ZuyeVG2pAKTfK80M6XHcg
OPCUXZ4SHIurgOdVQ/DK7BKQd38q5Fkl4Ximd2nZmIGgY5Zp++IwqYL8cC/epcZ6
mQcW51NUlQJR6r5GazlaFIp9+5JhcXLbBEAFZWuR9i3LTZmzjz+5pbBIYaHLq737
QVGkzw7i7IlkloW7CRAYiqu69UKY0ecnzQ7sUyLIwYVkDsC/x2/ez7iMZ8A14u7k
WT6tQSOljgt6H/QqQ3pQ3ka3d4RNkxS4PZxNqUjIyeWHR+4I+FZ8P5CG6CwKWNDx
g8a5egQpB0AFYJkBFOci9nxOP8g4Kkv6bfmMkHRQdBIexPa8K9acc7g/YlLKaBUY
xUqnt4Qi60od40u8sPvcW+daSwj/mVDDM+t/qqDZfChzRK1vXA+Amh2tZzQTq9nD
8JKQZthDDIFdN7bBhN4Iy+C/V+nzRyJVsCDWLX/zerI6yOLcmizEUYJlSEtJU4ER
MDXWUBhikR9ePvfRNLoEBVtyK+qLtxWz3hK0xz4qBhdFx4OXQDqxceAMkG56qsQU
iiXTZ1Jc/AxEsT56JVqCCRoimO9eoUbXfgCPNnpI9sIif00LU91Bi/U1n5cELmcp
N29XZ4l5Dqk7zoCtP1nKTwntXvJkCOe4Lut3CSX5LSaYzIdkwOpPM57BO1TPdpCu
GpfRKI4N5gwtn6YG2tLXv+nFTq45oSLiQmMzdo/Zsu00SSW0hex4IBT9FOfLRdw/
cwq4mTngWwetpGGgSVsHF/XD9N4kXp+l7IlV0Imx4ufT3V3bsl9wZi2REUO8sAl5
qMppIsmzeUQBsvHNkrRCSS6BWa71bC0gcAyOpjY3yWv0hcUUeDjM+Tm985ZQCVu+
3dl3cY4Lr4W16kPSDUDb7X0siVLTd6z/PSx3heC3bY0WtWU2Cv30L6BP1hBXhDkh
fqSoBBiqzJcsjJQ5Wr5+MyvdEVzKDooV4/ly3snQAyK4yDrOrR5/NLaO6I2ikz+N
3l+35GcMSVcXaQzQaKb5mLqDcQLVwjHGGuB3iH8ZLXaPOE/z4NNyzeVWf4kRBPus
qFq1GlnaF1jlgY0Y1OtvnE1LDQeCObsjaArfdKGFfr1iLkQ+rq87rvn/5tL/2cx1
pgyXzzjQHFjaR9OtFPs3i8H6kvglJ4GihXBM+URWD07a1f+aWI2CigkOVtiUzksj
Jvfy/vmHgF22cpAaIPlokDD8Zxc4jH3ejMm1hInRbVtVZOSyLatiP5H2TNSHgF9x
bp/q+WcmfVajW86wkxhdOim+ia2c1f4zjYZltqjwoDWBp2b5lr3pnnaUMYQVXRnj
WZ9SHEk8iv9GbkZJoqXj+IRQl+9e6lo9EotIEb7hxxzm17Snv5ywoKELz8HhAKCS
zbRhaQ5wYHOXtCyWiVOmfmTC7lQxCLLSE6gyb742oefULy6qX/avtJT27WJJku6V
oLZM9J2XGoSL6wTXgFz/gKOxnUgcP/AjYRNMJfwZKCRS/RiKq05HrMiKfNnGLpX9
Y6FwyfjdFEMU0ApgIgoOIbFw332PO3x8fC2K0vg4+kghvD4/591er55hM21aNxB2
BSHx18nRc8DquyLBk5syWAqR05JlxrZTggCdj2BRcXS3lStfyuo/S2vke/iV1rVV
aZH/1g4sZlDwkT3mIoI00QoMyngzDFD+r4veh7CKa9JXhAggSlYa7comw3HQU+E4
xU2/xtPSFpiQNTBG/f1/Zck7eAYByRafaFz8pHIttWSE/hH79N5MKCOqLaPj2ruq
Idt6nQMDWcnsvvY+Ko2j3kZoR9doK88bQopwMrV6hOqU7DH2tazLUFDcy5Zk8tcv
Vz5VDKy8o4InHs1Dni0+66CDw7SPU6onNKo0uEh7XbdHfrPhE19o5ZZhKNkWlrVQ
wyNbLG6kAQ/M93nd+W+jdg8gWttYhNPJ167id98Yxzb+XDFZ6BAYOdnU4hIfGRDR
7Yc7qrXKbmObFmD5vGGxlob193WOAQwvifJXiD73ZfYnafx1A9YKaH9vpniOzXGQ
yEi2x7OqkKyKREj/CgDVYGlnqEesbsdqZUNyXb13Zgxwa1S8wAz1FEXgPDXN+Erl
bVOAtsE59F4/iH8VjoYP3iGSFjcOV+zZvEW0hRdMD7jlGpKRcMUXD9ZFaSrrVBrZ
W1WNVYe6sX+Fdmw6+DJtnafghnIkj9NLkeEEwBV7HDSo8FfNLJBo2pbfm3zagui1
0Tt/oNBglGpiqeK5OOFQJlIYwReiDisuj0K4NYYqaTfvxZbAedvVsZYAyr9aXoGh
Fss0d1Xr9Iqu3kPWREcKW8PUH+Be8YT/jzeIFkAUxPVRfPKmuguudlXm5YusKray
BakW7Okb/MDq3sQYjVoZahetG/IvZoUinqV3Hoa24LnIM5aw5VRUrUO7xreyvpWn
FAXM4bmDHd2lh8QhZv1xs/n2HqVQHwoyFlqsACuDoNgwhWQQlexPdKrsLNfOd+0J
Ly/FkJJ/C2BBn6oj0eE/sSYQXJJxuBzuYdqLZdYJfJvjCQL02xSl1x0+qzqHYM/+
WIcZxBzruLN7zjH9OjoVK7+UJZVzS0xt0EX9xmcelhCVzn8TNofd50ucdM+eLQiI
jvbzBqU/nlNhYVHI1FGpkSMEvlpF3UjgDGgxbDk6HuphVmwpvFMF4rLet3h06J/f
G+TrSUcXN6yN4RIFvRZ9bbljiiBBSXArZb1lGxdnbbeXQx3F3QUYky0xdhlvROwi
Qwyc7pSjxTUfrcR+DcDk2o4SzWFTEQ72dwQb0urd7kR0Ni+X/RYjgXcUDOJ9YwK7
ufjaaWZuD5Vb8pVg/isdShmo4+0VB7SsAXQyV8vp75VED0n0IymRP9iYa4BWnBc/
b2OM4Mv9UdquFF0kdflbPMl4yxEB+/kYtQsziX2FZ/DIuA2zmovdkC7CCxHqGodB
7iixqJu9lPRZ7TKupy/gjZSwHjV2qYTnKT9g+MDMCwf5f6AuUgurHrrKpXm/FDle
LRHfnyX+oCMg2Ra1ljfRND3yNAFJ3Gi3mq7wpyt7yy5lzc7YfX9czj8yJ3+fZUsQ
kcaVsGoISH9/KaHk6G/3ll5a7MAUtwGHnNnTB1H4xPP7MVCfIEwaxGr2t7JPhd29
QSjTdlVnJIuzkClUnWX0qLm1nWUzOKA50DlwUf8KW3iUdJSa7wFYg4uAVOFNCi+r
9KeJJBv6VQ87ml3O3oNe2Xe93YLVvy/HJpxi1ccyy15C2PV7vslkJhIg6tlqoEa3
HIuEdb9ZN9an/AiNrsYzp108s0oGXzTXfy7WokrA4qzOIjUQUOBjs6NlTYRfIiD7
6SqWjWPZgvEqXrfRIW0ctsPrkd7MsRga7PqgMyczJ9oqRR7SbxW+kthZCjhIPkSK
6c9uiQ1Ln+zA9bsU8d/CgJYEjO0qIbI27FQejjkS6B9w4qChcrQstNvdxTxYiFBL
kGLdGjSAg2gIlgqfgHuQAtHyOtpZKIljYUm43TQcbTQ39ZnmM6kzq3OU7G7fYaG0
BZQlvM2vGiTDAbAfOzPSuUNUedP/e9F5aHgc/+D/zF1plD/c08HTN/ZcMqclvio1
3HSNOqMw9f0WP/aXy0vAyQcHWY0JcLzLtC3TpcBV7NLE69tIgPHkH0s9s4DmQLCM
pXKQyMGPTi+rvvTw1uusrLIwed8678pQlNfpHEv+YOS8nu8tkYTr52+XeoTERXcz
5cer94dkSRJb7HPCx/pzYA0XGzucGGoLF/I8GUkmJ8jmhivoul9KCuV2bGR3C0pC
vlHdDF8doO2ZK8i9nAlFkDH9PpxLH8gH45Qlyaem4nLP4Yj2huRpa0z8LSt5Oi+1
uEQsxiOhyNL8SqDvD2voOw/lLixst3hrkSuJGVpWWDRZenEQ6LG9D/XgbJabNg2t
fO9VVZthkR1ZZzYwf6FiSIFeGydpavEk08mEguW6NQWOGn7EONJFeRP3JsmDqH3f
ZKnOgFX+6zINkps9VTMpx2LcOdrBSM98CPXXoOYTddvh9rfaVWUrH78ET7Oz4/SD
pblVY+FQbRdFefGBuFP+2VJqOm8qEvzuAMc1xm8fAR2NUPMEscLWn01mTnmRt6HP
pwjH+RdWSL/wZUA99WEQU+gUsoIiiSrpPM88FzG0y1TI6UdrW0eDNlxwYMyGJk2f
kbgVVmRgYw6BXR03aEWG54KzQ87REK4oHRv8SwAify31xYF209R0+lp+cA3Yc2QL
BeCN5Q7QiDLRJYxUgl85/ApvUvJH4VXAn6pVpO4LVL8iNHY5d4T/QMU+2MqclYI4
ozw3h1DxSfpmEEYC1xlbW6gm+2MiAwiflc066rfvtrH9wDJMNU7hkmIHY1JoTZWs
APJEoDx5zuy1YgpoNyiqaSBirjSWpVXU4NiLYHQEaxOZjCIJDStgHS+FlhmlmUj8
w0JDKJWsTfLoBXJEWSblLNVdQQvW/18XPocRcbv3NMG3k5mBNohbXRFnyYkbG0v1
BR8jp3TB7j5RjBimjRKFqn3uDQbtNvgrXZMsub+UUwAzQsXyWGcHXcy1X2xs8r9E
mSHN0MLYQchsaGHDRHzkjhWBg6pc7/ca6GKcGFmYHFVETGaLFmu8AZ3XaAp8VcqU
2BNx8Dk8HfnDZRORt5PsUW0IlMCbp7ZFRh4sDk/JyRYybVs/p9C3HacCq3OejLO1
ustNdVk3iSGlZdtdxnDCjc/zWnwrtDJBoYrKNgYSJ9VG7+AWmaUOlEVBkwXbQbng
k71MnhgiaOwENxGu/NiDhLBsXJU5hqcvLTbrFpvzxSHEbqgkd7eG8nXC9+wVGDuB
L+iCgjHKG0eH22QGb4jryKPFCIopmW3sqZ1CF/Ftozj0knbC8aIxLCWZx1/xN37X
8YgqKZmA4OhFft/CXJvuBblLHbZQBYAkd882Z+TStwhbRjQUthHRbnobXlcRlLR0
a/JASk0yM//nd2XGIZrYuW5GebmfBP4T1GrME1mzROpBrCbrPgdF7dloCrJcg58Y
7sz+eLYiZYrwg/A7+jUGBAiAtywPOxV2fIAyERwN4SukpOVXWO/N6DPwvdpL1trm
gZoG1w/GvlXY9ZGOgu4P81Di5XF/wZGg0QsrRibl3LheiOf+we6o8foQ7XeoSzQe
AkDSki1V1Xln50hDM1wul8riAdJCnuG7I48mPAHqWMvo+KZONvJmTraScsRIAmtU
mIRv64x2MwvaAikrwSeDcoFGn5K7f/4+jP3QO1bE2/dFg2P4KA4koLC0+0JMAH3+
5bcJFNnz2ps3MFOIo18ojRPE0VI6vujen3AGs2Ek0eh4zKxBt6F7mYZMibDbi/sS
IMBL+Gc/q9HMBDGkbQisR8PwwCujnKdRhf2II8woUeuwMhTq/fkmDk+qDiyP+G1j
+y8XpVM0GTJ9W3Jh512XW8vTx/3phF0GdKT6txP04eVyccbCMLU3EExLRpb2luhS
lqmF6fprp0ZngCBvm78hmmRXaHmu6DcD2N1GRssooUZb/JAYzre1nP3HnPk5yVTH
zwsiZWTyvGBNeurEDzoshqQAvJYJecNUbqLWJO//fCRMtRWg0b1Qk5y1QBH829Mo
SqFzZTF+We8NdaoSDIBslHq9kBMz9jix5xqKTM0SDXjXv1YL0hRIU3oJ1IsiyO4E
6gYsVo8vRnZmArwFmbJqog/SpsXFWEjl7A5Zk19UlY9eh1pN6EUr9AfBBYwqDRUB
eHKpcYtvyM1lVTKwdYmAQiGkqjTz2WlX1Mi+KmxQ/qRHlikcr6ryHiALhqyO23BE
IQWGCZMATQ+kN5XQ69oAzkOETO7JKO2Y1nXJR6MVbbGK6pgdWRSKD63itfCnIhZ5
kwbZMlS2Y4otaxSSfIJ6/TaQfPhFFI96tcXdOzE5U2npaXYsI825Mp6Oat+PC1Vc
wv5z5djXBdIlJkBQxyVAMl+gdratzKnVkgbpxrIWyFLGgFOwvv6uikr7mXscmfue
mm9e5kRv8RKpxzo4361wRmfjU/6RT+C5Xn25c3WDQsO391ZBvxxV/cezWA/l5dXh
9GGOy3fHhbi7ANWyUQDhnw70qbSwjz0ujUf7E96Y3r7TJOcRH243PJ/wFREAThz4
/2bPzuod4e3T7oZ9vZOX7YOdLvjDXzQuaeacowR36bF2UtjVF6s9qKQUJdSK4xza
aYBwkO3e3YdQC1uFQ+z4WwsEg12kWzw/r0sVB0kyBh/AxHgvV4ThMLj+e+QP3/TQ
WeQEbhPYkLuAhUWIakhGzvBsn5cut37hS9T3r2q1tyTiHgoS1aWiUrTKavteMK3+
GArfd05BQDFI0oayB0TvE96O+Hro7BmSXgcVtn7W7LCQNH5dD59UCSLg3uZ655JL
t+XhTwMwLs4gpvcTRYGH7MqlGCz78fbkMssf/pzsaYvc1Gd4nzeY6YE6uG/GG+KR
X73OwZbmOApuKThur9U52hvqGVeLwIMpsk9K1GBjyZvlfEjishtJMxQa98LQEDNR
FRnSM0bqlzn0br5j4+FGUM4cOQ9hOndVdaoFU31ob5LlBV4TlXYj7xqQdxidm7Oq
YDdpXayXCcbW5AO2AHIROiFlQ1d4jYHOG9I3Ej7acCqJ1HdIrQgXPRna6LKh25mT
aM/JftoMN27SxRhUGt1x63ehyy6rlbf7MaoY112EyA+Ned/4ibKJloW0TzGu+Z20
1v6C5haf5aTGBxYFGCAKgUnVJjJEFqYFZtIzIiLEVuxyjr9OXZzd4SJo+6JsdjBZ
dsbxnQEtCLgsNVaD0yXtp6z0UCjt1j0Z66lqatnBtckXaqnMCwMMX8hu2jddUL9e
KXQNaFdHxdMgEravM/R5SLsCZhx1gaUIWrHxgL9xyS1k3Tho3gzDrCCpeCqezuMF
1ospeUobhLdkaREcE2SeG1wk6VP908YvPuTzFjKp3a9wdWA2OaCLw9cw1BIXjpZJ
RF8QLJ2nOWHfPKqZTyFj0hPAVmelDWTEBriFGLcqTXUflOAhqApdS7dShJxYtTo5
CNqtOVaj4rd+aq8NJjAcip4cwCb3IYzEyO6FZ8DRCRrJuWNuATCnWkfpkboNqQwf
bNd7Sox1jnMqcAdxaBksvKdF1tka37q2DBtnIEsw+C1IOpFJmWawfOuHucoEYd3n
DhLF7xrJk2OzE01SDlq3fN8asVcyqYkhjqWokdhuXMQdTQmPMqD45wiTaZxj4CQl
f+opifTqZR37NTLhl0uMSt4jRFrkI9Qjo9owA9eU5wNrur8HOrZkZqnyKPlDD4TV
hWbmol/7gvhLiIEvLdeepTc5uBChtAHZn6tBXH5dwlHVybT5xn8b/ym4f0G88OVo
TeYIWPng3wheCVwkySLAkCTR9WxH2IEAnVbfpfZv5dJVs+4bv8pP+mvibvzNDaK2
9BS+/lwbOY5FZIwHJNb37sxtUtXC8lMsH3464rV/Zr7KxQbxvmqMISPI9REHvlBd
CxTj9fjpW+gHIvGxbWIItZsXW7vQmL8WKLZQajDsgJrV5M6EzUsjAlRSRAznPdd/
ZihzViUxCHekkdNE1WRgBfzjtrKPyy31MjpMiTms1FvhWXIqxsix7s7KAPWw4ZLJ
6MP5utCufXOrC0FOl21Bh2a+Mzul5g4Swf/CFRGZVaQEQ3Apbs4SL9Ck/sujlpHg
8D0XBDEJiCu3aqp0GQfFqNjdlr473FvU0EFHjEuYe7hzSJf6UP+x+9Cq03WRjbtv
a1yGDftursICZFDn3qcF7qneqBD5qfg/m1u/h7q8gQ4M56366udTybNTtbkiL4Fn
9h8DWg8UtKyQqmLmkrM0om10KMRppV2DEqU0X5L12onYZStRRpgHg3HLQpan5eFm
mhpr72vsTMy1lwqYgqFSWUAC7phe5dMAlexYmKJuOyYjcIgK9551qCFPL0KwofEI
1LDK9a7aY5ggAzj9CVzj9xIVMlurnF+48uQaixcURLPyygkX92pGeO4b5ea3aB+F
ZonQ24wrcX3rMxihxGcwI/86f2vn7aVBg/FcY+T3NslfeeLwS2rSsmWThIy7Stap
/+S3yYwbpVXOFmhdQqPEHDsAI8gHaOshgHeEi0LQpyjcZZuCRa9D3Yd+20Ogg/Wb
ETVBfIPvnBJTdYAsprbLanbY5A6sPzePn9GZgSQ+ZUBJsMlnZDZtI9BU9aazdbcL
RkreLZYiEHtQVy3yNBi+ULTOey/vgzKgc9ywTjd6rICHC3n5fV619guQJuhXsfe3
QRGZ4876HKwkPnuyZjMLRJHd+PlIaf1y1gzcjHzpMuSwxm2OdxWsxA2uAVxmctmo
0Nmxtr4/fKcGzSWBa3/Ei0k32xal0ZmbhDARNxIX8IbEogduYn7Jr9l4NrDqMIpK
em2NUg17arPPlqhkdhsJslTHycTjtgIrrRip92LzXeAayVOKLNRgEj+b26tslS0X
U7djlhUZlBXiCxVJ9n6gxtnZ6odjXdzh5nQmjUAU+f1Y3ZkdkD6NLhngqaHiJEOH
wx+36Z5Zih31aNali0gu95bKGNRe/lJJICLFUd/qvOH0BTXd4QxUqLTj0Q54SUtN
evVLVSTYy1wsbqhODY05bh3lmmtCu1o3wet4A06Wc9YNhavVu/Zj022JLDWu5bWc
KbJy1g4jQgx49xoctkVif9ezDU3N7Own4FIK4KnquPxFy7Jd1JoeV8VOc8h32lb5
fadef3MrZeZaSXLX0VMkof8JAToxap5SEW9toJIXqdDTkkghQDosiMdqo2d8BA2s
3DjNFPIL8MXqGGRAkA9OKBHM19w2KsWigFhKTnyHDYYN5BAH18dr/12dfSKG20KS
i+JGGHO4iOjQEsyBjfcfYDgXtdF9fnGhHohhmmfPrN8HOF3QGbd+qHHkymoSmN9a
9uWKN+H0/y1SXr/KB4aGkuXDNz7eL0xqDzyQ/sr+QI1zISRyCTt2tLT63L0ZquUS
ZmYC6Neohb4jrnKgBtm3Y/VPmhHvdmeXDZr3pNlNd4muJcyEbjKCZznAztGycFyV
AxUkjHv2aaeKpndF9fiGFNXgfy8E8VrY8nGYkZ4nv9llqEOwDJzn9LC0V+crtMNR
g/WB2kKNY0X4W1fRRlT5oRUi79kQyni5ec+mANNfVhr7PFC1QT9uZwmDWb4B+XpU
U4stA7kUbAKGrzuQAmPrauwwyzl2zX0KPzWhc9MaWzWItT+JFqp1xOGq6hhUMvYb
89rQIXRbiBhG8oKi//OqgWApJP8e2YfOfXnc0WOU0xIaaGnEoC6LGztn8obqEGSx
GXIobfOh1vUQqhw02XfEtJVizPVnVqksw1wiYtwZAPJ6be5unC1QzUk3YoXPlgA4
FyokddPxGMBoOJ+MPSBiNyoAC3akuNem3xCt6rEUE2kP1F4M+VIRQ7yEqm72iudc
jXPrkrCNZAdtuRjRdbyKyocDOTBFV2RlhXaK8y1MyHBgHA5LQhQzxhkKds8yT5Bq
Pc4uMbkKNIfQ+z7DPZ94PrtNYDEkQ1ZYAuC7N6EsldA81kChZiPhr2Sc/ihO/jJ2
4z182GqrdyDCd0daTD8SvKND60szrrZ3PwaSp46mbBu5azSd7RhnT5Lj+28JILZv
Z0o/5GWw+ij1HQMKaCUMWfTCZ366rcSpaIAqmWRDOGN12gasEGTX/jDCvoxzgMP4
JjmQoJmsEl+mCIh6jhThe+6zdChFnSwb2jixuwPwFM/sxuQX26bKJrzXz9hc2FfW
H1OmRXENtP4fHS8ApMMCvPOxCmfdyGgkq5BerzlliokLzurOkBxjMlq9+FNIEilN
3+a1veCLoCVtiQH3gLVkT3C7BS9mrXLz2qFUit3anB+PVOT5z0UhiiDxXr6sMpC7
avbvrdvVAyJnpLSgllNgaVCy/fKmdTExo82xZNRMsgFA6qOvDlztL7pjssl4Jwx0
m653di7VQuFl8bG9LUShSZkhINLnWcGAvnMjmxmbTM/oZKWMJEpl19wKtuvMZTzd
EopX0GtpYiAKWrLLktlN9LMDzWgw99+yf6ChiJDWYn74i64CPdtUgN6MRD+quRrp
+5A9BJnjYRgn6/DbM0QafnrZ0gaz9c94m8dBvcA4umennBmPlzqS4yquIaPRIHbw
zyGjEnXwXBA1+xIAqPTKXIOQ6/xeAUkzc/GGEX5lkGAzC0M8HNNDrko5TmAQNB4D
a6M2oDTAi/9Wtg4Rc16Vhcgw9W1dGBtlGmdv3NlfjuDVxFntV/UmM4vGOAx729+Z
0vg9/uEYLHAkAhag61gOixr8IbyS/p/8QvuEX6tUKXO+/7HmQ1riJJV8fSDcuCnm
NcjinjOCg2doLwigDXbLHtUB3ovNQHpBX5EORsOd2+5K5U7RuLs0V/HOOGeEAKCu
y4LbyyOza+SesMYd+ceImXQhKgbc7e2BSUcOnpTSf6u0KRAMOOhXy3Oy44GTajqn
90S9iZJhlDNtbtFdIMJ8CLijqfr4flW2sl11PvoqAez69LqdQRAtYzeG7LCzZU5c
AyL52umH+CrLQk6nCAMvcaTpAg7Rn7ieARwI+4XuMy90avWJatQ2rXmJuHSacbYh
PNUyXHc1gTXGcPxnA/bMwoVWfllsf0NLp4XxN4MUdQU2XNBl0/wa5ys+hNFGK4D6
9x6cnvIy1+CxsjplzCvlO+Y/uh7DxWqfa4u+9r7Ql1H8E1UtOoUUdKZa5Ufq8fg5
DHmoZvSBKPLJwDufc6XQoiJFz721HvhDJ5aOrd6hIosLVuI916ndSsEymU1BFEh4
7KcGfjVAuhm+tkDRNseXGaipOr+Jmgu84yWHBmN5Yi9DnRQ+pR/LcVB/71l3IjAX
x2et+URBvj2Jb/i1EmDulBSNlOJEkrb6BVNueAD0JQFf4++5kXQaGlP1dTHDgdD4
+kJoNPCtC3BgV+1y4JbonzRCL1Q+tfEqa+/U7UEH7sqTflcwPN/6NoddRw7PE/Ax
PgS9QBHSYm4bjUWEKu7U7hkPnvDZxItSunqvDhjmhv4R5t1zSooBgnOUSUGHSo+C
HQdh00g89YSL/TV/fTlx+wjixTOCCa8jCWmI58xARSq0XdELjCmAflbdGaTtbSUI
aWpfoY8RhHj1C4XNQJKUANda1vwMH0jWEgyfm3uLJOXc67U7Ep/VGur5BAwVHHs9
lCQjIsL40DfLshUyM2jLsiD8V7oimPbPW7U4qukKF3+yq1UFPG1ZXeg247hzi+d9
VGB4tcKVdzJjJojwX5sj0l0SHS6ANiqkUGB0I9SV3Jh7//fsQZbknQOzN88V4wTC
EaNn88ZcF6vVyaZKV6tjXw==
`protect end_protected