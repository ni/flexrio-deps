`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Jm2uGAVYfY7w9Y5qKstopObZuZAEY3b/Io3MSEcWLhjjnKulVhCBBYAEQrAzzGsT
vMbffkdZgjdXQUg8jOLJXSHZ0Dgbnob2vlppjZs3bgyHCF7MoJ35E+LOsaLimUA7
hlqStcK49hR1hdeBPr/OwfT3UeVrRtQyq0eJXQ1UksinX1G9Pz3/CmcGfTZ/C72x
p9icpt0bkY4/1I4GBvNCsA6FFKH947JqH27OPACiQQRW/K7JToQn+1uhWr3LA1od
lbVrWu8PdZi7zW9gK3jiW5GaPjwbYQGqeGFs3bTKBILjb7sYHxfxw7eDLVMAIu5D
W+OTIN4JiHiE1gCnNEvkSQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="pm+c2fYA/4JT1uhlJGVUubML8hZi8lME4xPobg/m8uM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
nBaXksR//iZ9fraC7WMJWWSrjqRXHxmM1Y0+KKN3b10NElDzVNMlR76DLrcnamFd
2n7uzsxWqhhJR5LBl98SXO3Y90J6BMbw+OBG/MFM/zUulxh2Si5YK5G9GCrG9gvZ
5JomxuZFDu9CzlWGTuRUt6FsE4Lr6sOL1P+hraQDpMk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="M8TXDiNa0BVMX1P60yIvW2WA9jKGGy8GtbuPknDnC9I="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36704 )
`protect data_block
/5TNZvs8Nu0G+mfp7M8H+iVAGG3Mh5DYZ0Gn3rRNhV8b5CcJKgjQajrRoGl/gSxp
rBAhtT8Vd5eelHgtvBjpvFBA/EBUrRH6CG6pqRt9r2qUDt4UernbZbxC3BC14KYF
M1mXvS+9WI6Jij7CRa3IldWzDu0tLRweNOXa0jRfkD1+FLMPdwxFR7+XRTGjnIVG
O+fUZ1nF0rpJhRaJG64LWMoyY6WFGmc8Q1QdZA5jHAXBBw1WQApvYNkv7se6MmSv
kvis3kTrbU4kGwxcRxLAoacyb+Xbtc7rQUx5IMfVz1Pc9Fq9Bb3Ktv1zJhJFYgIS
i/VviKZBMG7XJ+WA//TGuK5Kv2ZYzj+LdlL7s7CTa/h3m5bPcwssv2aVck1k8oIJ
KpvX+bpJW2v92MNmNb5fMHM/TO1F5sScNNqIuApfzrLLFhllntEdcX/DyKObUqhz
ituvYU6kEhYfSwIyD4cSpn8bE50ijXBSB5LJ/5WK6YllsdJ1O756XYEkw5hDSx91
xu+f/du+tf+s4wGuS7zP1mIlcB7JYCTk2G0YjgeEx7TL1iVfJCYqbKCOVk8fOz/j
wVcQTEGf4Y5XgqkpQXBk9k+ZfyO8B8K118bdT5JFPYiMM4yqKSdkvaj5TRrSTU6o
KdQkdUwRoVL8PPba/xxfEWYiCA61irlgC//Ywn9AfbmUSw0XTLhO0yd+sr//dKEg
dgbRykL8m7c2Q7lgW7/iKcQqMve90uS9AhhWQubG3wdT7rF/50IjoRDducvp8sra
016zqhcWSCA1xdKVa/c9sHW71RLjBgDdBUrhibpnTFI6rFxtSXsJypvp7AOc0hfM
J4E8RwhLuiSoZYATZ8AC7WWzpawmxgWb4wp1DaBvTPVbQrRvG8jxRKzbM4II2dgb
Iz3gnnP5NlXarJMgGB0nrMC5Jey5xqHXPiMMC5S32xdyg6KEaq/jwKL4mliwTg7y
HX/Tcs7DM3tv7mjOJOwAuXy/yqlF/3k1gNjR01OX2fZND7EXKb8T264mB217wJjj
erzdO/EDCRSrPzA/wDgzNS/7E571bh2ou5oSjEZF0RwrszGBUQgg+u8thCuTY6x8
5GD1hVOmb1p5uK0SV0e1CyNzkITXuogk6RHIiDc7p8mtL5YJXjfk3m1Hnun6CkxD
/H47TmpsyLF/PioUqf4mAtEucw8mtqoiP3XHKQtJtwtmV4htmCqW+6aXryB3Mjq4
KKExDPY4NImf/iCIc81LXtvBYCPMBkB2gapH8MQ3rTs/E9QOXQoHnezJw4GV6oyp
W+mQiztMh6CgatnksE29aSCumEuw9p6UrqughL8aKyFYhV0wmByxgWZisRF5n825
SYb9SM6JwE37M0vld9gGIE8lkXqTVrNZ0/eHRHooqxNfby9QkyPiPPf2tRN+7aVb
xzPGKWcsbAensnDOzX/YiLDE16SUIQ+AgpcoHh5+N4qsJ04j5wBVVqKZMOMiaO+Q
8CDGmogURUf0smGVFwJd2XBUsEvFkcofpBdAq8bg9jGH4NwvWp1BMizdwRL+uKr1
YCU9CHcDYoD9/WLs8KuVHTVaMxP4J3nx0JY5R0UiZaEJpS3S6XJDwON3oI0/t6UZ
NQv/NdaUGTOkHyHq0hEGBFktFuDaIexkTTw5fxcYPbDnMUpw42o+KQzzpmMlOtuy
sWypnyGGUlsUKbtMemzy8nJvOx16hZaE2dPXT/S/AtNiWFtx1JBfXOVYGbaM8cnR
HB8FsZ7OGtD9aD81YI8epoCIuXZGr8lP7kxdCkjqQkZyON+gZGPwJjp398oFqRmu
4lawViVpVZM1P1izk/KXa30RLeHVoocapkxzGgcUClfKJvKmgKpypBUfo/oW24D2
K1MkCYmJ0GeB2tSIFuCuJ63VJ5iZ2JS//uUhaKKNmHDth74khCkim72OLBNto9C8
WpzbXdAPzQK3H2SraNe0ygTalUTakmznuVpyerEKAbwI4iIsQ83yS39Vcb8Q+KYp
ohvYCK24eE5gJTV2zTV581t0FxZBqoqgsS0quRqunkK1HTrkUjTFDb3HqoOgcEGm
NKIOxUZSQaPilL5OgC0b4yUJzJ0Mu+E5iXYgTE6xrJsPOZKOfDHkqmppb0bluzHX
H/dUx6Tywf5Q+V8q0cbv7aSgI7EJzqxPkmYR75AIlW9fl/hCS6YI7ilEfwsG+8XS
FOhfCvRGT0uPK9pUwQXbTKIMVBD13xqykfjX1D6Ifp4D5iO8g36qHsni25un5+oQ
gWCwHSNdpcNEqFEP7xuKMMsft6MTnmsiJbHu6VCZfxWAbyX4d7Kf38DskN4yWky4
PRKW0tCyIQ1crYHd5sjnJ82rNY5cRi+xzvYmnL021+7yu7pKATG8s1zmb6KIAdNK
Eab/nBAkPfbmghvMf3dGtvqKc6msgDZNPOJd+KPp3qhFrBMLhArQIZ60UDpLBREK
AuRo/z3QsL0Gy2BgKLd6lLIgv1SS3Fyjhb2JWGNEjLzCtMv6Hyc/ny5MZx6+ImDW
vibqe+3lPS7+HS43sEEUs9SjQNeQLepGDMWO2kHKcOMhmpEL5//0hZ5w0Vppesfk
gz7PshNGae/iVchdEFGPpEPyeJ38bmbotROeICybSzPcEq6PWJH23zNbi6gLwjBk
ihQ4UcLUnigv2nYWqRMxsDSM0DFRRMVO3uAWhyYiLZ0Mne0dXD1P0z9ZhLo3KbeY
aJTEZBC3QocImRtysbN8WGHG3/hkc3JCNo+5hNOAAU9+6kgAMA9sWqr7vXvSk2/D
5MEuoZex7soVB9unSzMMtL2NHP7lP0cz45a8xDWr1MvSlRNIFZHRTEGFSGjZ1zC9
cz7jwN7qjxFE5qV4r4a8cwUEyTfVfLFXOC1pFuZJFNior3gdTo9V172nngxxBZl2
SpgG7w5wqP18tEhDDSHQhPnQWnClSiRczOJbFxZxSqrQSN9DsyD4ebuuGz2uYaJk
1uM4/tl6LI8ktiYjU4Imd1xp6IEkiPOzyZm00UL/p+r1m3BVHekW67/fftsfu2G5
i/Y4jXj0c978JwUHpsbASQz8530pvZwv/HzGQ4sdPVhdoamXEPpNB6z5bSvHdGyb
rHudZqR4/KQ+9Z9B4NMzPUE2X1466gx5L4Hefp+r3o3JKFJOvm1eKqyKagu+i1Oj
t8bPE4Hcd/EJaAv4TxhG5WgL+WhjmmER8HQ0hxOTu645kchjTp+Q/6Gr4F2Krban
Sle9B78D4kPjf/BkjsrGQLAlGqyxkRT2sPnFnnakgQaFJ1R+H6b2XjUsX+fuFNEi
fyBQSo4sav8KqhlcCDacB0V3/t+9PtytC85AQERIH7iI6ocDKH8mzFobIJYw1e2v
C/rJ1cYyoL1LAVDtgtb9MAHnG6QAnKKI0N+gvTl06SGLbv7HY7p5xBDqV6VzxMzA
9Mmncrty+hO5kkQIzCYkgeKMXTFhMr6SbMJr6xBPWsW/1XL9YEFCExdMzic1QRIW
rxv5aG9wXKgNrb77W5hbxzCvaxyBRqhsWiEOExvXmPJ1y912Gu//VL9hyFDtQo+B
zLcyYxBKrMavRBjDP0Pk12uqxtPyYODLPZwc6zfzC1Q+dabazn6/CP4BwMZI4B8B
NMQrMFvTGpq8Y/tG83aS3xxfyvmcbTG2YvDhqQxIUEeswv3LYcwzNS6s6PvsV0rr
LPR8IHFFYdM3jeqEz72DURl4QgqvIv3tEEkAbY7qPN3SunoX0iDesLdsrqdQpoP7
QAR2AR5TQxaBf9Emx5ITzfpTPVvxs+6Eq4Lk+42lPtIib1LgSJWiA/GenvAHqBo5
eaH5M5Drb1WKbB2+wXrhjp6BgHJ7e40eAkjOFQMdJysZynLI/k4lCWDscxd7lMtN
4CYGqhfMM6RuPGIoPOF64q3NMlsKtZKjudOKHhS64zEMKL1EU24t9xDCXasTTMHn
NTi0HKlDmRYdi87Ujqu8VARq1/dj3UBKa+2hbRQeMyWyo2KTCcMYxbcB0BmFX+QD
0esBmySDVKGJJ+nHqfwYQNzSJg/3oYJjTreixXJ6QiHLctESX6Xa+Hp/x1x+fTZc
t9PySpaHnVE/ApVfX9O9vP7G5MsCoQ2758GDzVTOdGsrSF7xVBHKEePHnnIXvcxd
Op1W8MQFdP5R4iDs/o4GuyEdEhASr+w1TfSYGSj+nP36lCVQmb0TsAk8bcLTimx6
UPWy7m1ZF5iyGUhm8fTISJaXHb8y38EP/S+SSevIDPc5Pl47zSszW3lLFZUJpKvu
5ug16ntWrCPMRNA6zcjI0WUrdmNfnCFsWEKa3Yck6rvOJQZBWo8p1HpWo6nhIBNZ
32f0kkftrGh0R/1HDq/6UTwLLQ/hPslSQEv3Fu6Zq5PgszBAZ+rpisDNkZ/rKNuM
ryJMV7+Ywln+9mApvTRj8vW1CwNDa3qKxRQ2SBEFUGAfOc/515pO504vKTX9sy7V
z8bESu+qru8f1eD3CMttx/k8K5sHjyqIAcf7jc0Mbt3pO758TD9ylQskh5AhQ40A
KQeTxQoT7AgyAeuDIuyXlSiAcNUt8Uoj8GXIrqTpCDySree+TTgHglo5Pzhuze5i
rx7lz8R3HWHqd8+KHCFxS61uavPPYrNnR77yfkDCkOnUJCDCGaxE26nLzDFtzn7t
WE1WtcU05D+/3CcNHEJ80B0lgbCStZ0mmX34niAwnFNnRVCZQWzYyqQxh5tBL1a6
K065o1MjYrCk8ZHkqLmlBXWOtrTzyBPMSjaLqAIycjLyXISUEJcMtw2JYB94xO+7
g2Yd7KFttBJA29g3UI786GkV4M2CSezVzrCLOJy48NO8VDA3DFZS91KYwCBSCrjx
BBL7uAOeKEvwBBgzz//Wots4hByZcnXJR7HfnA2SUM+Urg0Qh1Kw3UNnkkvlCG5F
TiGMErT+jAxPqE706UmNQVj6L7CV8fGvukajpgSoObmOBVj3SUxT034SsYBvXEhW
CkHMmbAEmnSLs74N1wcc0Ye8TvxYydf+l+fKVj5wXVXiAwskIqr9Y7D0Yed4XppX
D29FXK8PdhOhF2heLnA6+jPowj9ZPaUJBRAJhLCLZaopX/MQXzez84jMvmrSwxh/
tXG3dYL1xmSPlEGi14ftfufjenJ6mrZKu9/4R3eStzUnUUrqz83DWqeL8glcnXMm
87WG3niKYIcshcNiME5brbgRPrToAlM2QWaor0OqjM9TCjlbzUDPgwMneKcfl2R6
fqM9VzWTUFHsswTDtuBpH2fnjaq4BIPUeulvxCqMQL6dEWz4JRAnBqGUIFoms1Cx
/NB/JwnR8eXzUHPZDAiOOfvk/eh2HWghx7HqUuJI1Fh29N2Nr4u/gKtHvsx8+bnL
WRq5tIPNcA/6/lhcTD/8mxlxBXJPRcFAEBgUwO3bNCkjc6B/E+kpuYmVUux+f1YS
7fHuXV+mGXwAr5L2G2O7+sxnkHn6xPxzu3cED6gRh1kjdPlyfO3usO7VTNqfyZqd
YxKGEqpaSCxPF5s/YrZpkH8Fax0UXIyRkrL57k2b7LwOJjg90l0wM5ET2+kJ9O4Z
iffrMDsfkFMXMnS9oXmvJGL6YM318rVxgiWX5ETIaabl9kRWvE467bR3xO/qtB2n
27wt19aHQzCTY8LLVfxCUvw1OX0UO5LyfUdHQ8eWK+iky6CHEau8VYyR7dEpcA2i
55Q38wkUrvigU+i0zibTH9jaXl51G6yH/ugNbf5rJGsuqPj/aoS8SxhmyquKwTyY
maI07KzgU/IdIYOzDEKY/xO2auWr4Gsmy3o/cgLsp4MOCaFHVclVpnBZn8f54vAx
w87bwEjC3XwoPdoSMTZEnFSP75w9J8elLGMlU4ES3x7dIHtIR/g1gjOrCCWr01w3
YQggj0LPV3tiXqCKOHueI55YP7gy1rdcfYSLsSncJOj+6+4XDVAe9c14vpETAI8s
EBcypQn4rFQDGoRKE+aQfsS1OzlP/QcmYThYStu5q9tSg53Fda6YepRKzMqSoq9k
eNKmIcSOGMCspzFXcwrwe+7KISVLcdo4o8Ftf3Jh8km3Y8xK8ktuY6j5X4Y5xJZS
lmLw0GGrYgNqVWTEMTcbRVVvQunn4GNTGCbLYKStdf2rZCZnKKYD/g+FQQOr5InU
cR+fd0hN6PaliTq6z7oiABfh7w7Q9VX6Gl8Gg8PCWEeULJAsWuPt6cU02tvC5rbN
LSugqKTXkRweU5JF1Rv0jChiaL8NEsemkck+7epOXkIGsdcaSzYb/PbXKIPjq4us
XNKWeklKq9GzlVMNqAI3l6GespUDMa8w7XwUrBMjUUKeL66HiERL2cacSHbZhAlq
FFGmgT1Ab6ngeQTsxNhrhoDm+9Ra0QakHMT6miGo9xPp+c0zj74ByCKN3JkXkQgZ
g5cfXyfdWv/QeXk1e7zA+zUnvT1VpvXvwgo6TjbSArxrfa9eB5MNl9jJaQ0mG70n
RU2icndLIyOP9ealzqkVME+026gq9pcrTGSGdRmC83VunJ8qdAOhP87D/EKMAOmJ
T4w9ccyvbslIu2ZPUnTQG8nF7W/O2XbC8yTUWYBJaBkQvaS2gjx//1av14VClh8X
p/UWW+oqcrESJlG8z7pNV/3gv1BRLmcbYTTJDcuTVtKsydopYDqwhckcfF+RgdRd
GsevvMw2ZPZIuhTGw7nKjj6z3ZVdpr61JsuTIJLR4jcl1DnItoEqFKlnsVaeW3Uq
my4L9eE02jgMteTOnzsYFxjSP0PyTCD9l1T6tdXLe6ySUKWEaMoVyr4jZIZGk9Kn
YcnDwU6aFPei3lsGXDssRrXTpq0yCV8TWh0VsXxGTe8cAWatjHV5faikYqpyhICO
8FDY8GT2bJaCWkGYq1ROwR9c3koKlyvfuJs9yPs9IXdBXt60e5nRyOHI7mtEAZWW
qLBVewExx4P1Hngcy/1c3q8+m1/38r0sUr1laJ5q6T5hz9cuKmXtPeUhua2iAlL2
8pDIDkJXvWi2SeNJB16iQVIJTFYJHiiWbhGITqM0jd3Fb3nIfrsFjqKymFyIUKcI
DDyZQMeg2j64Ml4EV89mNGL87D2HzHo7hQD1eqEe3r3eqJtvX47q3uTMtPSnFzUr
HgkcN1THtSfcRuC0t+XZgzaeSvfF547Z3hI6fH5E6sJVYj4y6oQ8RbXv3yJgddob
V4qxozdcnpf9NT4Jp0To6DdiVgfHPakSHXGMhdT/7N+ON7QeA4IXUvJnRrk9kKSu
HeBuTSAFEHBfzVGOi2WM3jb5K44B68I8stA4RB0gvMlHWwy3/HvAJIPC49VI6wLt
zAmNsMAuudV4HNuSoCri5NRJyyqg632rgDubm0FlgpjO+W7GoQOkV8kWzuKEcSUo
Ppr+VP5EBPCcBFlDld0Bun9KqvIzgsDC3JB5G/Io+U5hPloSk2HSMBHcRlqls9OF
cR+n9/nn8ayIC85FuxFbdiubadO7GZbYoIVvoU11NKgrCUG3t9/3BBr0T0t80MYT
Ss/9fNnVe3M2b2gJe0DaXDi6pGf50pm3s56U/FdwnFa9Cchlc6oKabWYhxnDOh2O
6GGCFmI+2rSzFTTb/wuT/QO9iM0n3gHegxecLSChdIiYP4ipGvzpgBb0A64GtKNL
4VBQQCSFhSeaTwYeiKNRm9/jfEFOXAaEMMd7SuC1ZBJ7AB5Af/FlRJOU71v5cTXY
bJ7/dd67ujq30LJIy6x+H/8bK/1PLfewLnGlWk+q3vg3W24SfmRfGlz0HIIyNVtt
tUmCSEQwtvuKE9k0WSQxd8uG/qg6Dyu9m+NDVKrk1IrB11uTxF71N27frr1QTPyA
3WfoFWHj6aF/UdcTPhEtNZNy9j0czmBtvWqEwLzHWpfQVs4NFYT6uinmeEN5asFZ
sy2yeR7al66usfUMCKixJdJuh+l6pQZXRb6nDSJ6mNQuoMXOioQ4ZTJNzqxdvKkA
CAavLHaoaYodDeRwxdOcr7rN5BDpradyPy5Ttl4aMUuZeys9hzHSVKWKY7GPexzl
T1w9e+hT0CSPptviyNuWWwhEBd47ouren2hYduIEpXLUfCVFXN4M1t+oCD0UefV2
EJ5N52Dzi3a9s/s7fJcdQw4eY1Aw/3U1OnlvSQV47tKmNf0MaosGOsdbGeE+mw8S
L/idvc28y052O0Aznq96xRjAkVXh6AXNYDzqJlrs9UGTJSzJBYOb8iFr90lCannN
GIFvBAoB7I7J5pyfJNDXuCBjzKYtDtEQ3Fb6uuWFVXi5VTfmanolEmd4nWV1VhHZ
TcJ0vZySDtpftQbRjCTVB6JxIAMp7gEqAuJfOBXKMXeOh3ua0hSeAA/nG50QKCFj
W/GK6VuwG8i3YsWzYIaM5gKKfDBfbIqkQihk/BLFNdKax/MeZvHqW601FrQ/jht1
qyYAdEQ5lCNEmU/NAVSAZniD3liQ7pMi4svYv3ttuGKDzNh3GKQggJ1eLP4/j3q+
6J1hqL0hJS/FuDYvmZH+fZVSG6/vCRBee81/GqbMWBcNK7mPk6No4/t9itFFNQC/
9VG1K7OrnfYfT7SYy0SlF7dXQkYnq/UIAspl9ZjhYdbhj4qczif8KVePXWg8HPd2
yFhjgPaDTmYGw4uEU3Nre8fS0D6BZDNrAiOCAsCjB8llSxiBZqz4w77e14NbZ5fX
ZsHWz22vaRX6YwJfdN2md8kTarWZTeHHjrNrwQ6C8hWGIg61pEkCE0fxPkxWtiam
vLNZapUPW5nh2jn4PrRWLNJO7xcyPeJPYgkmnhe/7v+RtIJqxzZQ77NXE0bOqwB7
paIKr7IDw/2qGv1OrevuG79xYmXOVtgiBI8Vm+qTykKHd7F30WKgIYIWV7tz8Pkj
JzFA8Zee5wI7oNXsodYNlyQY36QqEV9miEWJKBdUSe7zdIV3HxVE9nYeCNytbSgp
m7ZhWfKmmrKu+UI+xxbmeW7/PJ5oYay5gbSKG3RXA5SlE+YZQHI9Zs6nP+T/XiPp
yLsxsZd9S3J5vtQkWhP2ne24VqAfd8WzLESJYfEWDcegdj/F6ePP5sOnT04mhG0d
3IRoLsi9dCpUvrp2/EPh4iDGTwJUu7tj19r4Tjn4p6osYauFItuELcmVCvH0SEkt
fGmQOW8KgXWN+yLSoDYsEaA0+guzcX/T+HHSq7gYzLo1n4Y76E5RNlv4GKTuWwm5
iLlMlLwikeCl1CUPWNd+76UPhLRJ2li29PnZkE1rZ3CYN+fza9k1wPUeXoqpGqjT
jQ2ILr6XmMDakCsjCn3/QL4r8dsetj+qD/abHr5QT9MuvZiZ3DK/2GuJmnal84fC
EopRSO18LoayrAMGEqdxxY4TXPQhTGT7kqICvR17ZTo/R+tc+mc+TOWsxPbm3WoX
5Ec6alEzVnZxPhrmCtUDTPzg3ZtMQYFVJIwkin8O+kITpK0xbP706VJkv1XltDXp
kFV7ex7q4xEgU/ZpzLXk41lhIIRMqENxFKrE+Aj9fQFXuzYDuUPmNJj1I5HnpvrD
LBHlOOJnAzm9J0GfnjfH/ITtOD38pSei+T0uxwmbb5KNUavz1rTtIARFpQbXS72P
ca7aA3Dv4azj7XnzmKTLT0qUyeK65tLDXQI/lt5ScZFoJCHvObwxFUm3aiZMNk14
1cuTNVzzAorOrTsHRYP0XRX4UliXZlMoP2zKKhjv1neDAf50hZcDNXLYJSYKrEsQ
z9Moy+vVp4GG+EtIxyggHcxqs06lfvlpoYIDIEdfa84r/wdPsY6dqucoCeuczyAM
EXfqjWCkRntB/h7fmIkB1LDmHtt2T1mOu/fVDa+f02qanCTh7OeBBs0om3n/Qr5G
fIbVAiPJxgj/+Q5jYcQc5W0qRBEwLe93zOu0XNRarzyXuzbg2SJTP0WyZYs+OdJG
eXN5yAu9lOqBzEXwDDjkgN6/tLBDiYcwfS+by8dtLY+RAaVyz45/ilDtnHbINy5j
qWQk+YGAMVQzA1E3IQ3jO+r3zxzQyLEu/b0yWiWDg5ktXB17TZPnwD64W3BV+KFx
fMTVfgy2H+kilq1VQAgwcxr1Lg9ke/GZWoogw1RODtTVpWOkCuN2e5f6fXDQutDN
piaZ0LvezzqVcyqDkdWAs9sPcwTTS/3aDoMDiwIC33weWKT/0W2wuNNakCvy2fNO
Np1Qwqv3p1KG6+wQKpzvTqDj9WQiUte9NsRNSG6pYKgWTNDZBIhq2vygkCPD4P7D
bsyS4l0/oDoOggLNR8UN5tlNr9Qv6jgvHBVtcNAQTa7dXgCa00YzaY1FpBKtrdoS
dllvzC9CB3cNDAl8m3fwRGYJQ0azmhqe6FLN13k9oqDSNuj0ZPjo/fPKO9uPDc2t
IbFNgcPQYyXC85bZAVkTpExQCSG4/pl6haRgwkltniqIdT7+1Pv+pVk4FJG5wHJD
OSGHUNQLSW2fTs/P7/Ihdkm93zm95wckN7DjNWBbHnUfWOBVUl4oQ8h73bFYKBIX
SHgl8IOtDmPnUJPVSJiAtJMjsRph57OdfH1iIIENo5IYOdfsMwY++vAp4Ap+aNiw
vCDKau31l8+XQlai/nZ5HD/SjTWj8tDVH4kAQKml38Dej5x7rs6op9Y1YoSH1bI2
xJeeU22KFxUqV/KPd+PwVFswx6iWpJFRRX9KKrea/wc7GSx5dV/8ZrhMGvx5iS1j
9CIfwuc+nOpV6zyO5bbt+ZeX9Gq2hXlAd26+/qGTcOyRzhykfAxed3hRzXrtbQhc
AVw+tbKPS3sPZfbgBjvewMttR3mzrQsd5YdmV5VP2pPPB65nUaUQdqfDNQjJ9cPU
7Lhb7s+XyetYwlZpwzCFgHLP2eTz6Uo5w8HaMacjdg2ezF14BU8ebyK6mUTUoOgb
Drhhq+PRAbbEm9qXzfpdZO1hN6/+IYBTZK13HWtI+NBUTAxgv4EAQyCkSFknfKRQ
QJNIpFsaYQUm6jRfsRCoCCe80UFzpqdd3olvtRyQBO6nNx9+wNLpsFeOFwUIdR0/
qMrsDoSw3dK8POPr4b4p4JeonzIwph8Apc3+eESOTS83060Ovbuk6hZ8x/k18XJJ
uCdtUxEhkngWT/jBue+VKV2iTiTKFmbvNrUd+jvZtpsZwB7kT46RC3dc53QAIaEW
WeBt1XiwBggDgC5V0gy9zpDrHypRvS+KIxCW5BOi4N2+w8dSIDR4eYWQAjrZI1te
yE1M+UiLUY9G3MOWmerro89t0WrAIKgGlTqCsl4rvEY3yw4wZVdRqpNlN0+diqyD
fzauRJO6vBucCoHZ8l/tSXq5OoEahOKm4DiCMXEPkYeC/9BhWHoamQVhTV0iiHh4
kWzicFzZ6Z1PkKUAXsvMAAEfU8+3JM9t789HGEJ7/7No4tZQ+58AjnG6mhHWmmeP
H/MXlP88kNvEda/+22PmLfNH6HNbCsfw+2NHUXijXYmbftl8UvYp4oYT7MfWLeyw
N6yw8dFk6M02RUx7gIxqd69T+HxfuOK+E0e8K9v19LIls/RmAE1eEfnS2dqB/2uS
lzFjWYo5UfqQqlO9cn5o1wWI2AjsnockSvs3ezdrYAVB0T1slPH8QEqf1dMwUHkB
NQEkV9bF2NMbgXJ9SKeu3pnIREUqaPfehyBxxwq3ScIZJOR8pOQH/S1cZdeD0FKS
LyrED/VL2n9w8LC2Di8jzycOWPG9Dhtj5q8Mu/KDvrpP9rON3ibV1ntt5UbUwo9u
J8DP/qbfjvWtD45dErBb4Oo+9GZYJtNP1luBvvolTs9YvvYq+QlfrP0EuzwlnGt0
U/guLcRFVfcBxOrhE2/MF4TE+QgTcYYsKzcAhytYLVXe32+xV3DAFt0VrJpEld83
h8Sdfvz95n8GEOQOMvsbA4yxMse7Ys8ppFVh9cFJGwZrZ24S24AooF+1/jnssx+r
N+H8fOBhl5yEGK8chv/KRCaSn4aTxnuGCvp/lcuhyAi9AgVVz5f3Ok7+tkHyB1g4
cBOms3p6hkZ+EVIvlaHg8MPMJvVAJNcaUeLuQNlZEsPxam5zHygahbqZyvRBY13/
DONABnpHrnW9xsFl6j7geOMsrSmQfkC2IwUDGTGGZZFovglTEVRhya8AokRemjVv
hOWhgOrnOnkW7fmWmNikPgzdS3fb8HuK4jV7D1gDyftEWVln12naZ4zmIiZwwvgw
fcrbJaEZmf+5QcXuBFzl7jUwCzANfM4XMsQTvJJibuiyEpQCAMA7eT/iidXmsyMU
HHdO/RyqzlCBEs1UsEewCtB4mMQW92CHW2uyyxSOJP0opGn+vGRFjiPuGPSSESKO
OGPoTvO0S6zn0OKYjMKH+kOZvcGsFjXqfJKVElz59cCf9pUjbvn6Pq0stUwIZAvF
bRFj//Pj6wgMOm+b44FKH2Q21I5KYNa5EzktZMXE1Par5e0WacEcUEN7e9yqygpQ
ZLARkCr0taeEJMv6R3dRbZhfax2/F0OnRCKxJ1TPspLSjaxsQbgVxKfzYGxHWgcJ
N2H1c63jZrUGz117UYukhcEz0aHVpzPF06EKmQD8xx8pKiVI/RjE1EPhwVMOcdUN
8RtEHRuHyXjorCRtw8dBMIbzwF7rfLT0fw+7l4Jnmqd2scqXbwz/4VZVIPfCNq9d
iZiG+ajdzo+mdWteEZzTU7w44Kh7BSYFu8SgBAaMITDXsm27AdbnEKTrxe8qDQ/X
a6QOXW01OTU4OQ7EDhpJeBILJImy9SnvXMJdMR7DmEzmOIlY8UXq29ziB8uIw8cm
9nnfgvzfRbwHJth5wok5nAKlYTS7tBh+ij/v5ttjOsulXzA0xi1OHBNa2xs1Vxyd
qqbnKF/Di6bZpr1qY/dJ+FrqzShA0L2GzuaQv7dHUYzZA4W+1sY5FP4htYO6luZJ
ww2uYSSYwfue6f6ilnf8WQjeam7/h1nWi49r2IRQMq5J1yJAlUiJjIRqlwcDnp1E
ZgzkQmQ1GZSCyn+xHbH57LwQsK6oY2hzTses+fegAJF6eStzM36BvQyFGBMhcr08
dpE2h//aDybwWxYUfn4Pcb9zZAJP44gVjMZgmVwUKhxsDsfvnmTBdceOHaJsft1l
X2eVB9qSHZLB2CnF0ZkKGYN3Amkn1lUOdzrJRez69TNfcPa0KQgZVq5033FsjT/k
VO6h4X6VysCS4wWJX5zy37bz8ThmtI3BpRJDVsL+PXGUtkEosQ9Nf8k7Hy3p03jk
aRc3+Kq7Fi2M40DdhlkuUbNiZGaBvuKWZMfbA0xB9FtexHMMH4/oCdv+2NehQoBZ
qOr9f42R8Z18JRmQqqaW9JKPCbKXkdPu7QX/gaXr5DQH9xkAze6XVLleYj9vg1hC
YODZfVMgur7f0MjaN677Q6Bp2sjXokbmWPaFT7wlijDQT/zQqlzVrzv6TPS7skIG
/Qb28MSy/1dNCUSTU7lkNfNjz6buIMw5RDpouxE2NkX3g3Y9ASOMSl5PSBrvgwWp
QiafrnBB7Y4720haPXrhVdtSx9V4KG756UAYspqCzGQn4f7vivhkadhEDzc8MOWI
b/uhjtlt4TGZzq2vTV+qXkdsw03QdsxClVvgVnOkwuUpoDOED5HsnoauGkbkmBgz
bT9mF3INT9MW8aA+5XEzgU+rj3uVdJNO5QXRhTrzaarttUD5uWw0QsQBcjdFkanw
RL1WsuIovn+Gpme+6YJN/RJvBkL2P7sYKEINIUKDtwY59n+pXwGJeremqRDHSu0E
omRBvD1IUYDB1g9hgz1AZ5PS7BYCa5oHJOZ8Q14sjmEG1lzNxzz3T8KpLTKtuaBV
w6WvusfZwwPPzqtFhBj4pIvonbA+Exr8K+Yk0U9zNOn/KY20OfHtMCfHCvt7sg3Z
I0GMcalcOME6Z65IjdCrp6PuJL0QWXLrhRf1xpCvtfQGSbdf/nD7eLcU8bMHEhYl
HORS+ivNbYD5SmGHsrmG74xNMmFgc7RBjpl1dvkJFDuvEXJckGB6eT7rQAFgIItT
AB9Og4+MJSTZHeQs4GucdbqJ2ICwNeLwAyqkk5c0FkoVfJ5OnvrBIXQAFOt28cfu
zYuPJhOi8rElL6PjsSYjOOFwHhjk38ulmtO3zsRVIG4/ufqXAvERskdC/JxF0S+V
WGHBd2eISEhfTGKIsg2xCu+wkEggnmUVVdQOy1SxitD35GbGZ5Klagj9zzEEUBhS
fXEawOv9MdZzJ2aEMRWD00/XYi0Qw3rP2Nzb8EYs4jor+GjiymNqizC2xlZ1B+On
Sfzrf2CGO2i6ZG6qfbZvAPtVzCges3KjOTNeUS2Yc5pZh/EekPlndOhZx+tCiaM2
i45NjwXkiys2FotVMuN0WiSEy0mXXeZZxN/A2Sz7RDDCe41662BQ+/7HfNkROaib
irIZiZAe/Tkiwy1UcUYkougzQrPdXG10yvvo7ARZAkNOKKB7UVfAlS39b+ZqBvtB
2dfZI3fmx4/GJI4GHEcp9lgMaDpr02TRys4sYnGFJAKi+xVpwDV0JdDgiNZFXX7q
7VOaocYohfZX/+96rI3nV0xIBs+ZXxqcLVJHPXQhXxinBhTflioAPmK1DLykUwvn
VdJURFKQOgX7BIaT0zBA/VGW76UxRXlfYX87fxO+VhEXBmxjfD+eDlX6icW8V0yL
cDdn9Kk1MdHdMt9KfsyN/ys8gcU+sJoX/FOlc7m9BGV5WtJvBTa04/KXXd+ppiGH
0VjTfMhj4adCHQ2NYUshd/xv9a9Q9FTp2Zzgr7FWrlS24JM/CZOFFNJ/tLuxqC/H
otlLrhUb3Lhxlb5I4wNiAqL3j4cPhNFcmv5BIpKWt0h8W5NeXuN8RDh0QfM/90cz
NizJeHb/cqHUW62UtbFUlgq+3lIHQKaUb1RqVWwZXqciEvL/gzUa+8/G0uqcqXg9
Pqxdx05z3f1LTUFZUhAxJsFL+d8j9R7S1HIa8ZSngNOpDWYQ+puHRBoU4uAeHKja
L16p42NOHUcP7FHXZrxWMdps6Yrra2Nv7yEomYjKhbRzkMzLi1JiJTglH0MnHiZN
ktb6FBTdVDyCXkJy2EmogD13XO83cpKwpcjfjYfQ9eZsgeyLXT4D3cv4fQnd0ZNg
mKvRb/hxzSjFTohKgBiSZYJyJ+1CImXW7ldHJDiEeznyRuPuW5SKkjbBhxfm/6yM
/bWNdt4QBiHAKLjVs4TReVHpHEcnXAsoI/tyqpktR6Ryml1sTAzJDoD/TJHnHMKv
dPYcuedqq9Rse+1VwQydkEMhl3hdo/e9ZC6ZWXvqYQcky4aVpamkBs44DA+zxet4
ueZ62PP6tvYoqM/PZpNSYj3q2fqn++fqPnHS17Zb+Rj4/914ZPO1qGMbZBfbNVmR
7oH6WGf5lXcinUFOYgZtf7/oUMlUV+jQJncJ5fEV71tG4455XrrFMuuI5X/P06Nu
CEmmnzztx95A+JBFDFSjGWHZ0uTu+MNaL2JDsFd/D68bvvBVbLmnL3S0uJz0yLuK
GLquX1z8/UaW3WOtidFWE1zgmsAV05hMPNdDbUQmHArHpTEpj6Gba2UybCD4xBA7
cnYhiWQ+LFSi4Idd7z1kTEZdmoJRYyUcq8kE44Cvc6KEBOn2ZWJ/z7L5Dsz2naj1
SQct8KEfNhhHtgxl9lI8lCraT/zc+DuINz+roosa3YMOKQn4oashNXU/O7RF9i4a
PpIxUn5OrWfYA59yZiN0C0eavfK7+t/lO3d6aPckMtL1yWKaE7JFcc0BJ5BEHI2k
5pVlq5vYCiUayh1Cx5Cg98jb4wfp5rIRQJMRsfVY9UYXDL5fUecwcAYqFUrd2HHs
YZBGqfwIm89DuhfG37NDh6GTI5/ikfHYKGx2rKv51si6JH2Sybpq8pwNGy6lFUTT
IXv81H89JtE1EjfAcHKmQRVjc0bcwrXn69CTo9/kUQzNc9tuWDX/KhHZarQKP75s
m7cKDs9b9besC6qkNM4qgWjfLkO3ORlLw4gaabvXR9P8t0YviIY2ehksYKLPzd7j
wb4pZNL9f/vfyI0q2MSXph/gUvLLq/0NS4cfbj1o0OpDeDsejsco9aLtHmFkkoNG
o11AR62XDF36VzYENLp1PMe5rXMDDDfkCaaVv5+RyIz4hgxfs/4mz7A3lF2hwTYv
CrMf+8MKfBid74nZyvLxznDkuMpXfwIChVNv2vb/XNqMfKrVfwQHliKDvS+tINq6
i94azhQCo3sRK8BRh3sNCUSAPTtpc/eV9QFM9Oxm01JkjrINgaTGY9X2NDG+2Eo1
mN3Z4AMkpXVM6XHbURmdEXpnqPycV+HlVJ6eFe6h+KCODpnFavIaBpuBj5PsURxz
12/TSNDh4MvLEMNNk5MRvBXlJIQr4VIjZysfxfxeXDIcURFq3rjKtz9mDgUwrRtn
jS5P7cA3UXuxjHUwiuDaaACmTqQRisPMwXoODPHupgBZC0EALk7U6e8S7liUQ5ao
T84L++6eV4BUInbddoEDT5KolDxrn/pQDbhJ/tU/AAAslBCOxVtxIiL+cgbqMCI3
ybp9ZHn6RMCJBVP5T92HMb9zXHIW9BEmMPe/4jV+Koh2cuKP17E4cc7opObIsUTL
rxoOZJyhQUTw3Dk0MUvs0zdBm244VDiZkIY1KgZA+Ohc02bf/8NkfMA7AIvACiPq
fqXPGMlckq4bsJtO+21M5j88TzdAi5UmY11xPtcJf6nkgOccbPmR/c2/PyPNlLQ+
ywjJAqmbqt4iIX6/B2iTBrjPxxloFSe1l7wIs/Gnu0KYpUQ9Pf5enCyCqOPMNhpq
rKyOfDFSBfC0bxe6mSn23uW+q0UbitZUeV2ejWNtnq6nQgmszW3IoMnAyZhVCfxM
aXPmJp2aC+PNpBUNMSCmB4poDnT+rGU/31nQoCnLdgwKYNm70m0DauXlYDxvJRQq
UUgbyQIa1Q+yMe/tEyTNpiIiF8tcd/RVCYmnLHQryGfbyfnR2uEC0EqSEmeJOGrR
rNiFsBAXl8v2yCATwFjxtKVT5jXjQ3iP/9CVmSXTxbRm7VRXo+gnv0EWZF5H3w7a
KJhDDmNlmlFDN/iEODqD8K00O4o2iqS5h+D4t1NxIMPeFfU9Pf9RxLHo/bN9958i
JK+BnuhEO/yKsMGOud3iEWKOYt3aTVrAyqaDxRWq/bAxe2vZVMUeND49Ao8sS6hu
Rl+ftwZXstmkvbcUKno5UVJ/LciTS6jjDsFMqZtwF43rwn5+KMA87JnvZlcK3YOP
GArfptWAH+zpvvSa3M0eJCWgQyk6vOU0TzoCr2wwIYTidQn9Ecz0Gcz1ROpCmtcK
z1tKVKQ94FX8F0kwOBCPZ2NTBHLxIZYUbscjnLorJFlaVWSpoqo3T0MmqXhWEObq
u1oo3nMjM34mKfuimU5c0cI/d8/t50VpOwftXhjD4C38TjYMtDBh1av73YeAc7cS
vIIyGQPEyANj8kr7adrmnuovcCPrB9YjqSSRS1vHaK/qC2s4Dzz+C1QlTa2uaDjD
x76fcZdE8crza2jcWBFQ/vuRt1DwX6mcibnnYyU7y4EYxvZkV84jtwh9l9B/ABlW
gKavYb+KS3PnAdw7s13iR6lxp6baOzEDZLkURiQjRH2lTzyHudTqtBrCZqJN3zrL
J5dJYVqRDvN2RR/hWpmgU1Q0iHI64chZaPhbrcLxhzx/wOvZc/7uYec54/BG1lNs
jN2wSWXfaERoS/PMabxyTHDNv57kRFvJGXWaUeeGRNlIcNZwE14F1fQCoaiB6Dj7
6ToXnk4zJjQiSxcx+2P3IUjmbbEuM9cyYZdhI5Dn+12W+GI76KcvDzUnDRqNQgiU
hdtRlr+2ca1s11v6rTn6V3SRgRi035fyF9hkp9EH+17G0XNj+XVT6R8cmqp1tBTX
TH+rZrRk/RW/TjsPqBvMsMlE7J0zzuN2k4Z+jHfwteNUThvaOTxRgMZMbM7F7g4e
MrC3iyQp0evQTMFU3Jc99tmPLQho1GilmebnoxjUp71EOysmdmcr/iVXH/wacA9n
xce8QOSYPlqqm6vGslnOPFr2rES/1Jl0aY4h86yb6z7I/0F0uPGoZNyeoYseTiPq
PuhBSt5D0N5cWJVrFjuehNMM3uvrUkQaTBloxuk5lJ4c0/8HSIhJ66NbM3oCAhix
AXD9GwJTHynehh1Io1vcCg+wdJOEgfYOxDLIow83gBJfjy3UlE6feai3i5HlHpfr
OtdVffhwLC9OefKgTdscF8k5GeS+B37Ul1FHlreNkBv01ut7KrO7hp580RSUXDu8
3hXEMtWoSEFvpoBj6vKTgi5p96WV++Zk56RIWMYe4EBEfnaLTdLu/uAhqHvKtr9X
DRfzx53uF34+SWndjuGYCk38aUeQpwKNzjHwbBJNxXKUz66TkCbCrxjk/48hQipj
kckRSjunHxNqUj1q+BXw6C6bYldf+rgoxhYLVsyxzBqNQK7l3G4rD1EFnUkmi3DS
SEg8XqgQp0Dy32FMZCabgu720qF6SZbKhux2PnWXS+n8fohJoE2ObzCQh5fNy59n
5jGKTja/JZKqwMvawmG9sCWdCiBVPfxeUUuptFgWFo4/Z4abRue9nUiF8GZDnXyz
x8y7U/2bLs0vHCMZ9EIuSAVwPJxNIATXnpNC29cIgpnPj92mn/tmPLscw6v3d4X2
VM0GQTwrWxHROSjVS9EqArSvFR2BS49nmy3pOLLvLosyaEoc0PG0NDgsLbyzq7Y5
rpcCkF9nBSaMM+Hy61zBdD0TgzdDS89WpUekn/Csdf7YUI4Yhzt2ibQLmk6Txi5l
0DVT6sf35WviFcpsCsq+quqtpegHcfzAyqz6jO4M3k/5saLq4vO/W5MgFK+nWtUc
Cu/GdvM+9G7977WtQc+oV6L4KZSbpGnKp+6Xo/71uGkW7uJCaXIKbmDrNZmDITJ2
OUzyQbYRanoD3pXxlByyWlUUDxZdigbjQWrcw3kqwSjVP65Ik5uag/a3dJvgedsK
ghi/sCBK2JDN0u0FPx8DlB7A+2iQvd71XjsUyMEw35SNqG1M3oI0RLZ6zCKFt2Eu
vcnva74Gg3PWFdh6YxtMCMe7hm2R51wYpfhjTexUoTyhwxRyYRUJxsoDGbrggmVs
xPVK30A2l2l4bYGfveOGnhqYg9PKAKnIuiquJWXmfbbkxKaA0R+rmosj2qj5vrih
bMPKu2VSn5liEuWwUnCWicn72Y/qqZOQy/sGRJdUqvoqtW44SwadfWmHQL4l7uHh
d4wNSDfDLyWcK8ATSR4fmR0t6V5hSY3+Z0xV9mN/0ahFINW1IM3iVAJ/lo7rNpQm
TOq1Gt1Uskk0icFY44f8A11vG8r3WIueb9Qf0whvngccTSW1TqQU7hOzbtMl3UJv
H/BVAufjnSUWqs0z9ZI3r73f745Sstk9EcTHneJnWQs1WrNIyIIu9FM06pwvJwwx
xSjaInYlz1zKcxg9KfR9ZIi0kfSrZl5JFD66dlMruERGrXh/o/3xP1WAMOqPEWwC
W20kcrVBYAS2UlTGn6oXdpZMaowDj9WB4KOD6sOU5dgYXZ41vqawhUOfVY9AT681
XOgUch32oy9cENEKqY21qdUXFxO4ymP7/xd7XIjhI64ZAgVqHrZHxTlEi/lg5lbU
nENosrblQez/M+30F6jocexvLjZ9pxtZSbouXxUpBFGKDbnWZWDiXy3F3ddNpzFY
UFfghjnr8qiyLs+sCSD4tBkvzBG5spW77df7mya63dRKs1tFmGU2A6DUgoWbesVI
4Eov8H3tHd82QIIM3YpQ4tILtaix9kZTXkLOOmIbj+YEYznZhFxUdDBfkWrgjG4a
GPYOv3au4GUmS5Rp0K65ZqFvb9k/Z3Gb5afEsrIQalX1AzyM748GL0tLvZESGnuq
P5MAWctf6xPmiP0CKZRs98l4adHRyzf7R8ClI+L40UHssqGzfjA4R2YgQeIv7woU
qRGhe4cujkCgNTDN+Arz77oRxTBDS+0sef75XluSnuhTSBz8UCTlacOeWJMHZ1D3
v10TqCAgj7Sd4ebEnwZqiFTtCcxAautvQdQZiEJYUVAm+mr83ZamitLmpfyQuz+X
LlBHvzkDNLNALyNjVtAoAOxoHjBiTh66ayVgklMpb9jml1A+zT0HhrIEVbdnBW1z
lrFZYlwI+cMwE11wGOEZPz9cTSIohUQNV534fJWb3wkGpdAqGKn2fr3yb3sf6vzr
u7X70AgTon+4FRUsCqnKjalS6C6G9BdRXYD0Am87P+W/2GRP1TdZRIUVol44z6g/
/42a5AIAf91bUp+vhp349OCiw7kNqa7Bty6onPW9LyhG6/g7LVErB6vV+zr7RVnc
nD3GheMFatNaOJdJznjwscRCNfn1vPffu5IU2u8sJtNzuJecsMD0byT9/3E2dukz
gXBWNTwfrAb4LPlRK0XYJCTiYapewmVqCWqEnqBd2Fb2135zbXv0Dc/BL9uyS5kK
F+lW4LYnCHDGLiHGUhv2yTJK3e4dflx1bR7dKevdZnLlnbppfwZwpYVdaSLMBpxZ
xQgTUbYumle5dMISUrQDrSEkp1aTXzoT/e443e/l1F5ojwUS1Jr+LX50wztGkwxU
hdi3MECWsesMmB4kixaUXz12YCPqJtmZvg7ESmPsf3pUu2ZvjuEY3MC7dGKWlf+N
BpQLf6WzoDe86ujgcvbfmw9BrNZtgEg2oUTL+fcmVJYy5W5MxPebEx8yyLpSFRoy
4iXhAlOtf4cTRhIJoSxEgmOESKBvRrMNOC1albEgVUdVRQ0QN1gs5LBRkPfx8fjY
l+3KCJbLlDfLXLqaxOkXZcoVTNtqLcOFiDbvdi6lou13Puv8AFCnbBdVSLl0pnUX
M+cSguPkttgJ7/NoJ7y8T+DtLAZ05Qvb8TB5lcg3lV1xqWfk4McPCU3NuBEhs7/U
Ym1imLkqAVRGHrjm3pyJlu6WV4awo9g9MViHLQP7mBBYP7gBUZqR82m9216F8aVd
j4+hfGWywNDmDCElI2hu6G8fDffgDCS5p0vjXQSaCK/HSIrZOcPBUTm9Wn8ONCBq
Ffz4B5wX1Mai1g5nFjxGf/ZPYXdLjUEdyFOH0waVRK/NPFmzZh5T8n6eDNKWeVK7
t9r89BWOmGxYPzbtZda9zkO0aMyDRBGCI2ZeQdzCGR0vEU9K/sPxZX3ASXodmpoo
BfddGnuk3cdVmk4cfuBHKF/bcvrxwfDRfG4vc6Ea0cKcf0kgAA4SF3SJRk6XaJf9
rBl7NXJZPsEigeWxMt/1wMztFub8CGH5KTt4tE2UOMnVrF98xSUUT0DCzlmYlq/J
9DeB4IF/vTnbIsNa4mVeUBFt6U4ykA+sEkAwXfj3WgE3f4QnN5RCmPbm2EpEoTpo
allD1Duwoha0dhkHyPRhTi2FsYhXT+mUkqx/ckwQ/loJwtmbvgKDiVi0pkppAtWI
wMHy5CBz4/hKBNwkT3T2ZG1K1OT5j2Rpk6zv6eLww556rnkyrac4hnoE0neGT2Kz
T1IAALNJ6ijTOcVXoTw2QJIYUwqQbOT8wKHRQgSgK77iAEyycs4/0cj2wATxqi7r
T9ubtfABiblbOKkwUFu6g3a+YuV0A4J/egDHe9XmOlIajqLIhYPQ3iSkFUfJTKO2
oL9oKMix7uybEfINukfjFomsVcy06vFLHZ/z3QXB+DvPmrinZ26Ouk+D2l1HlYyn
DTuqQFhQS4B0y6/bRERIWjtGCCGwKLq8gRI400XVUiImTxNBoxDwc25uW4nzHqzq
rKoIhohNYxqxmsZJBMoLNAFaMIyg1GZr4RJpVNC7V++QWXxYskmPq0SPgTkk4Fce
sd50Gd8AFnyCCDkdn7ifL05z8UUXNTeD+R6yLk5QUAnTss4QC3M05EW6lVw+isNr
0LSmbLdqEJaPVTdLg/hLEhPvvdKFSz8/9kPtiu0UVwXs5LTF6B3vZy1f6NI8PBHV
OlxdWJcIDQ8Ox1771XmFQj8qjMdodj2i66nTaiiOagDDbXVsqLt17BQmZFNk9DVo
S+dP8VkzDQ2zxnY1yUXZV++UcgtuqffLvRIA1ClDA4LNzvg9Nd/ACg3S12a8eMjR
ZgkzcQwdPF6jOSGoOUh5rN2qPdPv8/KW5GcYQhdrDSxSNuyHk0HgJMkX05mgcVas
WcfFAK0mRCk60DbSRMu3THWyx08Ppg3e/T0Q6hmBJhm12RSNEOehoFqWVRQVToZE
+tzMQ2r7ZTd0iF4WDgB/cVd4f6PNFAC8xnT8/t7gsLhbR8zvA6bgpwpdKNnQeKpK
I3gwX23zXGA/LTLkZDE2J25xQO9PDJSxjseCgM9U8TgHIeiH3oVWYSESJqFSzxw0
Mo42vjXcJBIYoKVoBuPNm3JWKkmNl3xwJuoS89ufUL3RY9A04k/+UqXpfOJoCaTL
+g2Yfq18OHxd4Gf7JeowPje2AKcAb0jL45vRCdtKeiWXD2u4iTnB5DpWt2DkQ4a1
3+cnyP3NejUspLOuOBbBvV4EuK28/W4cF/xrLlROv5K+yLL+h2xRVxxXgTbI0GyI
jWWun0Gc++KoZTfp+Dx07wbQH7KwTuU9CDqM+E22ovQ4EncxpN0w3/5tilTAp/fX
regqyvnb/eOFRP24Tvss+1cbX1FPEMZ0wDxdhGjOQauJq4V9QzP9pFkSt6tgSWIu
9Joz2mP2CeDA+RMeQF8VIl9FzOGQZI54wAlIMbKwk9W6k8DGJVw79YqmMskgc1rv
7Je+66/KE7PFyBMFJIQTM1TIpOer06nVpGdkNBH8JZ5fZC2GyaLuwZ/KluJ9C3YT
cP2hrrzhRbfmlqbSY9xceR9BeXTe/zUPV9PlSVNS/b/kNPpUwQJ7DRtbnGjl4Duc
yT3/UURJVqudaxoPPDk0x4M5T1c0spoL7sdt1ezCq9UfGetmw8Wf96kNlE3sys0j
O46mbs0MZrFW8c30WBZ6sDPEGfttMTcdglv+mMib9qi8Zwm1Juc0+2jibK34Ts1h
vmKHGC5gTbP/3csBUKTSmCsxcYTM+Y325p5bOiyFKzBnHcCFLEKbgAHIabUMp1SL
s/KlHR4GSB3MRb0cH6frBPl/KtoxZBnRLh9oucg1u5bZnOW20CyJlhPPvb8rXpxt
u1YHSQwNqAUFDjbI3VdihWJmcLmo9buVo1wQXur7ixvPdyrQ6R4wMbHyPctHFJJW
bUbBhjxwQgwJBi1gdDLgNJaDBWpNntlRH+/PzbQoWdQ9re10gbPu+HxXPJiFuT8O
6wMkdQsZWtAIx7CbAiE0KhIgo9CbnvKEGJhjhEsbOLNE3NnHBoAsUAk4OiS29YaR
ERSCUJhfGrzlIRjenBiIb1y11Px0YF78nU7ALuGLq2G3qIk205dIZCRi2ZrHfc5s
2k8+cJppuzG3yjMlI9RoBSM4CmpPHqZ1BD3ML80xrQzj+MjuFznchp//MtgUH4Ce
LBvcdFVjy2mn4gA0l1jCMdExJ7S+lsUl3RMaSzG4sJMMonX3cUC+bI5F38CeZZSg
ElSrkpooUcK+jB3yHexNRnEJo8/a9o6/gEaV+stpjgGWV6wfMkAvg+C4t2SPd+so
MiGl7nCTvMW/xai9ncTMBco5lgI9/ZPLCqftaxRvD6IfA2+R9ad8fdEIVP1FmPdF
m3EuKQWF6Wa2L/IloO5Z13/fyCm+KlF+hNg3SEynOqUonZeq2uV12A5XZjidrq50
emd6SvoejQaP8myiWePKUz2n++eJGVQQhZH8z0dQir7JDKXxZNchlcFKAkngwv40
BMMszXzJ3MtWdG087kRIU7eP63f+rnjxLbCxTYV0BRQpxxIGQjbRI2asa7LNSfEx
UF5STYMxZMxef3HwJ04RWCGDuJ3NxZj91CdGwmzpqSRD227FkqHuIeOhrARWG03S
H6souMNW3neAQDiPTrp/sK6TGZRhrumky3LPYAojQT90+u92HvLSA1Aug8MuH2GP
iGmbzyto42qBiEC7tP5Au8KaXlTUfHvgw9OYI9H1juh6uuNufl0i374Pwhiqt0Ni
boKe9TNZLKKDV9G1Lgyv7THlRLueds1UQxMaCwNrvG3OyXtCGpti4lfMx6P2uje5
PLb1NPiNmjbgL8qeBC+/mQpwyaH3K3VDX0iX+GHzWDkKQ6Hnsa1JAKru1YIhg/ue
BXVJvMUfDDOaeKUuKsNmA5QrXsTgfPqC0zYFq26YtfuQ/hy8I6KznttGhpakEyxu
KeeeX8EwQs9BUKoMDCaQXOrNmPIcRivKSgMb8IueFORSWQUzTHCfya+7amUM+mf8
TIH1SzLFV6VqXGMKT8zgOnuXuorIVD3UgTUxXjcOPW5U21JPYi9WgaJFZOi5T2et
lgxfK7QCYB6z+dCqZc/9AVvD/Whve37Y2BS4P2VTNbU2vOjhNzT6T9WjquTMv3jN
qjVvZAb9tZbcIw5aODf1K98lHoxINiM/EuZq9FJuaPSmYqLL0XfbEAEyRf0C5knA
i1Fm7ma1hX2ogtDm4Nel+CIcJPyOi7nqVrJJ0jVTYy0Fl/IYJBqW/aYF6yVwN9K7
VrMe+inI6ZDgxq7OKLlT7DsEKneCH2sH/G1dNp0OAcDeH0ceLbxrGPTpZjAgEl8h
CZHSRMs8+untjMSEW+1intruFRCld8hq/E98bV97X7juP0+LYSNguZqUxDBZEmrs
UCphL/NFdoOx9x1bW7mbYESbOItAcgx6PGhdjmkzuMIzI3ibNApuvMGuRmyYu38/
GFm/q0esusucT8RfIe4X/vQ1AZQthN/oU9l3J8uPNmaG9QbVl2DyMcdK3WbDdnxR
jNztRgYqCIldsW5pgcQEA9YXtch+YNwe+zufX7DiZsMoTp4j4p48s2BVNh4IIdwQ
cHUKrrjSqwU3ffY43YgepLwjtOcw0ZNFseLL9BKe34FVCu6xDNn4xhGxNh6stMXe
OIeKf/rEaC99WFSoNC8VDfJvosMvl7T5q6HD61kC3QV24XcQR+KiJhZvINXLsZNJ
+4jTgmtNEKJQGyZnX/Y+Mi2IHSe6tP/56AiVyb4Wa57vL3fyHk5dECJUbUWbJ74E
cAQ9+gMSguxWX2IOEJnY8IETZq8/GMVgCpbgjt+L2uAjl2VnMZzs15df5q28RK3O
RXPey2STcu1zm+j3qjdv1yDlJoonpsg+9tSS3sJTpeXR7JXJBDCmGdx9V/dbG4+7
GOB4a1hQJ+/ryf8rHCIg/+voH3SDM2gJxpnmdW9YMkPSDcLXICV5m1DNnR7JHw9m
wrnzSrTHKrSj+M+OkBPyREgGmYdKPjk26vsOQXGEDUZFqG5QT/535M2rKTGx2Xqk
riZ9dOi1ppZbL2skEWQpygjWMedk086Radn0Izoa9TfmIk9qOiij98ibcRL0LQh3
ojAJXmHmOp3WionY/CgsxpW5ztBOOSCQWU5a3YFXykB1hzERs6BmBb9He9EqObun
+zzBe78pEYWbqrk4P0J1Zdskn2Z/KqxRx0z3CZ+YM7m94TeucMPrbid5RyxXJgG1
An0g+1iBbfTbOP3UK8/iOpmAp4Uj2jKpzLcgOmXT5hO4C0ordt/TZCq/jM6v2WV3
JVMz4ZSbKkSGgazjhsbocGI08wTG3XoAl3xcTBEpk+n8lkMi5so7T75cely7l/IJ
43xFuuWmoR4hAGi3PwCvcLyM+mBzJcz9wF1h/0R4P2vLZ0IdhWjwWIMJWxzN/Ic6
BAq8dnOA/PTyegKWv52lh9Nhr11Ga5f73TVchyPQDrPmB+iriXx9MztNRxGVyaqU
Irml5j545WlqSmZuKAcwxgKCSn5fSVwuKNkg89j6wNT+CJXw3XGjU2Jmq7QjFfMg
Y1zmJgF4PVlkNt4i3vHBfERGm0XC/mRMN785u5v2jq2U10q5KEglROSAuDwcKfUd
t1OKED64wUbduZTBCwK6FQTTs26xtxF4N1QM+xen9Ae0E399MrJ9UsSaZkqjldZ6
neT/1dCUllo5XBQhw7f1nYL/hnLKeQIR235mNkCZk6B4lo1DKyq9DNHcSNf6NgR8
w3/qrD/+qm0qsltJzmMK4+Ih/pQLcjZPVJffTkSgmkoaqi1y64ePBuw9W35eewoe
BGBAowflGF755T4IdgNeRlliZ/LdZUBtBOQtMpaK81lE0dXAaoPnQCQ5uvngSz93
M0BUHmIj4H3IRQS+Iza2WNdoxTODEoqGvA2hksl9dTKwPAN8CWeo2lNqQ8zGQcuV
uaSLbm26BYMHh7nxD/IdlrFl1606tQTATsrDD79+YI/5JepmOLn4InxoKFksIIIM
+fEz8yZqqLo+zRVtvWA8yFA5oeYemLJCbyruIj2JxJOFmZmQI1NyQ/BeJeCwfz5G
TgtROK4rp2bOcOyqrdPm3PB0vj3nI+/SeUf0uzM2FoluAZqorCAOk6NyBeSv0EJR
Bs3p52Yf4lPNjypFUCn37cnIaBsXpULih1eisHqGvjiomui8cIAVQyXc370Qr5D3
HaIFT7+75hqdx1QzK/988pq3DHuhcsHk5GxqR/PJGpcUmSyBVrv2y0bEWdMIpTlE
vX/bUcO0Wm8qO6T7lZDyeRMsLe7bR9VbM74CfHKyrxZZ9Z+tB7eHEkgD86Xr8fLG
+vhl35qa9QMPlZpKJWSo9p47WuDTzfeIXb3aOOALPdwBrTta3QR29uZr4JoLt6oL
YTw1aEh0a05Bi9+p/H0H2QGUKVDGB2JD+dqRgYkT1dhI85VHJDo0UAe7iIGaANl5
SyZVP7+zRVFqVFKebCFBO7sHggPJzFnOJ+szffUvrvYyJQw1RXuVB9syqbGHRQFU
NSjypxTc83WEXECxmc7gl0OL3AzPEiQWlLx8bBIU61uK9zGumgdQGIje1vk6B9+9
PV+fUdso8LvSXEqo+dZGAbDHQyt0G2HavTVg7mtiujLlr+ud8UqkQofwwQTJdXRx
mH1zCHl4c2swoyoTkmsGRW1QOaI1ImZOjvbERG53t8HyUGiL6OZm8C5FZ3iNfi4n
7o+96Qlw6TxOGFJp4rIsLGeMcIQZ4WoQbKWd6g66shiNzGkWtl3R7NYeGwkm019k
DZVtbR/cWo7s1ogI5aZb0rJhE0RhYZEur5NUHg3eCyxVyvikP+3Qu9wfINCug5U0
Xmps2C2WTmy9D9BIkKfQRWtz0CpSSBNnajNv6bgt7BFAv6Jj2TvU7ugGH/2wCFOG
gUdZIJEU/dnrNEVZJXu4bAyKGMv49s56SLRbhoAAgGaPOhuSJnB5dyVczsZWNdbJ
tTFQXDU/AKkTZjMz75ka4r4cJO6GWF3xN3UHHjJdsTg0uHpi8Z8mtBIzD9G7/sUG
W6xHiIwJ2jZnRu0VUPRxE8uH7C4Q3uc2dwd0poZydMG/1BghgeRrdmGwS+nCgdw/
/6AQcHc3W1qGAbXL79LlXkO81uyP5kqWSJHrEwgNXoUyl4Jw4Fz2D6qZlwGPuDWJ
BNEJRtTSSg/+ctvD73WA5mzAfL2EjhnfrZ7DQP8F5A7a5IhitCxzLed5cKkQzoJt
2GaiLLg1qTmUtR9e3esovBTqSdWXwvHYgbhN1sJ9+DJs5fomm84eFDTarWvH7ELO
jd5PoSeYsYAojg0kf7JsKnHn7twRlrnVyKwtc3i3Jhk0U+zl1Ys8w6GPMF4WddIK
ER38aK266YYEn1hwfSratqcJMEJ4ZT+P+OIRgX7cFMmM239YHtVGHcVOri1xk9PH
iNcOFiR8IO6LBj+8fIbZfDo+DB1w5P7ZaFVF8Q+o6t7G2/wKQnfTuvLc3xRQzbua
I83vSFlV4FriQWturNgL9kdcxaT35/FPnG+Tx6CXQpCj0aGKrk+szk+T2fdrlOkS
2SdnSbPX0ohBP/PR/ejYJm7BiV2vTVH6pD738dgbuAgElbloTydXMO8s717GUVmj
Ie/CDNKKIcWSlOoiigksb7Uf4fs+GNzZV+Q3KihUFouqBY/hXSfGYxSSAkdu1lLU
vJRNIhepkaeBalTMjEik19myakB+JVWlRHFQDcuGUPwteJAfXNaRVdfhZBiN6rC+
els4BxE4LNDKmPcYDHuqGwYPyLyK5SC76TAWxtwnchmxYw1ZNUR9pf4EQYhDkhg9
gdSNHxpOtRzL5jQQFTFs1zIpkofqhgBoP4hKwHZptQO8CwmcHlmLQ7SQyi9ssWNs
N53mvcxUOZ7Lkxi+4PJ3syq6VGmcqe5d0Fc+1HPzrfosKXjQURqD6mzmf5Pwh57h
EzlEDY/Kp5bKfKxm4j8db7eP1CtBoCN6AlTL3kWyiVsAJL+X/Rzembe8DHjWaSvI
bdZNi032dzA8zf+kLOimFo4ROCFgBoUmIdaY1q/kJIF0yymFNO2/h+31HeDFxb6p
zW/z+O5vvMJ8z3Ko3derefOUJ82K0HyY+7C/vvsiCj/DqBxbX5nmGGGlu6UPtYLZ
Kv5oAY24CcJhrgDxc9eEc+AtWT7hhYxYNTJNymx6hV+U/RDNsNFv3sqIjBKsEWeM
tbMDRbVP9fv+5pb1zNS9Gx7AMzgVo+kGpF90QHu+Gpn2c6BRDvTEe95q7+JAK9bS
m8Y7dsNanGgqvDIEehj5KO1PDtoyuxU9OPfYLrjoQiuht6Pd8yPiHWJuJtU8D21p
DfYMoNp91FODIvqkyJcTUyqoJWvCzpL6AuxOozDKDSRwK8T5NOGwN3bpVAtk6xaN
vAnIIZglvv1ZjaL2yigoN9xCmvL574kZRa8Gm/EVsY0MYE3NKeaMECcFza5Ntt7c
qyRTDNQqtYJ5/S588U0YhkwHbHiMpkgnmwunPaWWKBZfyBS09sBy4oBNphcyjnVM
X47RLBdTwKCSG8GUmAeXaQaAsmR3i8FTXTsoAKeG6UPnxn+BbnnmlO8hkWXxZLBU
YJth5fj3dLq2njPcpS8NSQPu6NL2efr1JJ6NGySv0jOVhmEo5zN34GD7tllDVbAh
mvN6Cw9ujyL4rTNyu7h262oRTkDAhlwbn7d71idFiNGldwJWdzNhymzLguw3npT3
fUQ6qofkUBP0N1Xfn2hQ4IE/fSH40kmI11ijDXc3xWknwsAv5+MSsg/jubevp+y2
aaO2mXiqXlsj6teASsSuMWAcPeT65pGc6PGBVr5mgjSsRswghzV1rL5Yr8Xstjmb
Gu7AwmVkD/5OzEyQniEEPogfEHFqFU1Tj4RoPldYIIb/qQqMVy5Lx83SDJS0nAh1
h3nG8tc4H79Nf54fmlWRTBXKMn1BkwFbMKb8WwIJGzI6cxSQd3Nlf8t10BYO5rB0
ZlUal5jo0/ehiLpEqIRTYpkyD80rdJABa9mR5mhsTN9/k2cT5WQxi9Y61wAN2MBt
qrKs09U6CQkLyc5RcXhKLgR87kKGVoM25uTVlUM1SBvx/a2MSlAy/vw+e+fdihHo
tBlzyYtAvzSdljFdTXXen6DK34GseOdy2UlIsvk7JQzsOx9BAs5o2gxjxC3a+wLx
enFjdGVjWb6QgLB7KMXXvnu1+Rsx+y59jzGUcGpmFLtkNqYc98lmehKsBBDLQ3ac
tPoPC6205IJu3CBWcHNQZCDh0Y2YLczK2rkGIjfR2ZB4GI7c6gDM+4jxZR58Dgtl
TaIOM4Dz1bm4Gl5PtpcIPG29p0Y5ZooXSOS8qkRfqgit3Z793yD4RCSfMgV7kBVN
18ikZNt7nYm/Dt9LkOjmg2dpKpQ7SMxwlXd2l8DBysf74nAtlu1d+ZaoV+PncqyP
zZeVinyZMg5SRIFPx9xhAD9KhgaHNYfp69udug6kTM6bjAHX3qrfSqout9fJ6pQM
nv8ZaDqitqzO5Jpo0lLet32oaQzBj6sKg+87OPCX/3GA6+h705QC7AD8LcrGj1Rn
DyzNVrTgv02hE81kHwXZR5c/duLpfHzN3bCc9P0TXlCNJFNDjhhJIA78QnZFVt+E
jZejYhkJpunpMKxphPxP3xmIJOYdMT79VTnLlcGWBg8VgghjQ+pWqrFAq0PJjG3M
Lqt0msuhCTLTL6xsz7w+Gc/PqO5Xmmfx+6pROz7qy15FnRqqEXLoVpBnX72l+Cqy
FEY8A9eZvEpHBns+9nbXcNehC9bQDV7476+Jv1qhmzdSV8qC3aXQQPU3T4Lamhb+
1aU7tnbfnuGn1ekk/nesnPvXb/cpvCma2DnwicZHD1mxtx01qytHWStPIglPKvBs
Fv2BOe+np9bCrYKvUE6OajyNgeaSupkTyK6aNUwvEp3K3TIvAUdi46NqdoFuMklD
A2hQk9Z/CYocQJepVnwBPid277fGjtwzrHy7ctflwEYh5Szybox9z2brIvfidNDc
7wBjXQ1HVTYcEKwaBb25V6eW5NRI39jmNUhFa8oXR+R+/XQVP/VUUdPMl9qOVTzo
bXCJ4pbSzAHs/UQ3DA0FJpKjXo3VD32u9HykqLdDscZlXJsixMwZpulMyfq7blNn
+3gur4KuktvZSgVwuX5aIHyHKpFVMiEbST5dQzYqYzR0l0mj3/nzQrDikZUT8cYK
5Hm8bovYoeqzLBOgrx+SEYP8Dx459zvBzkwJ5EDAS4vrbklGK+f+4x9VwEViFfo0
a6Vhx/ZNUww0axoj1lFScxXhcmeho0BmDCdpItYc3IBk+rIHdLF9I6rIif+7GK6A
fIn/By3l88psSCXlSncLHf07lInu9sgFU338NHfQRQ/uYxQ5D/qH8UrMef05y5hL
wrMywjuufX+JtlXzL0k92GHPozNNMrNz/52w5CByhrAp0j43F4YFFwIp80PsXtOg
flgcAhNaGhp8yyv8M+mItf6OODA7jQD1Xjbmb2mnJtOJVrRN8qMph/+mVs7gZrst
gMT5sF6iJ2Edr9Yx00kRVoLRSsLopoQBigBdE9uTmtO6HpGFSRtbIfwHqTpMXOON
6t/AwPYBwxpzFrSAiin34ttZ9HxM59jCuWy3XccGp3ljm+C7ndSu1rOQ6Y3qGjwd
LRiUv/rVU8tyDDfa9dwDIK6Mb20UScvPxEuKNofrKToI+qaNuwFmru0LZnkjIC0Q
qIr8PrYBxD2t3OfdFIbGRUZNHBEP2fpzdNVOYV+lVfKKz4daxZwN3ox7eiZad14m
zQwqjLoCTb1cQFXvmIRlk9wPcDkDIPRHvOOK6mDq07KlHoIwC8GdQDWrHFaOijDn
A4D7AALbeFKBpMV7FVwqP/HZLHN/qxPYsC80cCvXAvMsovH3+ivfQPP2GHu2HWZc
ZNvH5DsW19Y2tpjIhQTsnSOiDtRiP/5Dsw6mz08VD1yJwI2KjREROdi7sr3kBGeU
ICTommF/1IYEzzOwLR9jgeSO7kWOrYcBHAWeB2s3jFzpjU45O1ckns/UMcT4Ymeg
MKXc1M5nHVOr0SuPwCuo1rMh3804gqWgFRQVatBUA/yVSfC+LoGzsiFMbmpuB83d
J0Qfvksd5+agJXSe7D2lOr7MD/13Mx0CGzDnmHOicFLa1/A4NcT3CsCPzjAJfEko
M8JlnfXcqzSym2EMtAvODyMeadbEGNdegXxXaviDt/R8sf1Sjk7dh6k/NZHoZhft
/ZWhZqbuEoeTsPZTtkGVCCoPE/mGp42nh8ogd4Um/f/YrMytI0v6wz8UxXrWljvw
X56gmZ4G1krywomZqlx54r2qGpnDMv16h8q9wpHHu5E4nIuYQ7EXCoC86jCbOaRh
OzF0x7W0BMf/L4lvsTX+CIkSY7IVkAy5798CgfL41jUygkqt6b+mgcl5lAIt+CmS
z5Lkuq5cANQmstyalnYhHjwHa9Som7GMfu5VMf3Qn+V5qLfNqlzFGg0NVA6AvUed
1DL3ZyCUuVO1n9K+sfwEslO+fWZqyjxz7o3iOi9xJy0a31f4uUQ3xcdAhgehbdCN
lZXBh+M5NZ0bq9B/bEM5ZGnOBWloQv5927ntaz6ozDAWl2U2hgBixSoOx/7EjoDb
QlTnmwK2t9Rv8XrYyG9t0h8QC7RkWHtaGggKIYDxe4bEm/5JbJ/JfbZRpcbkxxkP
GsFfWfIgwmJx3L1xEvRyHrmXNN0NgV0EvU0mXVqY4tmvGBcbkJmpLbhGt33yXo43
ZZN9R7PKcsrIsdR3GEnTp/k0BUl5nqUQD+i6CoJRDC1AgP4jdvOU9pXSOzewtssC
OpGikBB37h49ANdjXK84ua8H/sucDzCBUVSfvxdcQ+2vesW63A7x9RfMdBk65du6
eosSmdC9Qp7koXgQ0mNOJHIkXx+7I8tH1YyLyW6G7mF3wJt+nXbdMEsy9jDs9+VX
XRtiwLjV4jZRD/13sK04Q6rafvQlFSXIPR0wStbl/wXpxrRVbs4RnkBRYr65oZCG
wYs4wf2Zxp7lZHX7ueh2zVKxMikeqwifDrALpoAzO0JU2cUBfh6HlCZmopuvWTna
0a6XpNuv727RE6YUEg2ma0sTNQcIqVnn8ukZ9M6Km+n9f2FEUHaIoMrw/eAWXiYl
Lhc9yy/4dhVwjXTE4Wa/fbPxbqzPYh5TCRig+vk2QAq+R94V4bDNkzC2P0SWsbyU
lv01L34ubWyw9pTITO+kNakGduIjXUhqfrTWsWKXNi1JvOEdgPtMlHxQ7CAnrCbt
94UMFwX6Cp3vtUnxVIkMWDiVh1/KnF8/RR40kKmvYojqlgOWlsM44uS7PDN8wS43
SH/F9RilIcpoLchJe3qz8huuvCyeHEgfWJBcoNcImDlpbx7omsceiAhiNes2w04j
Rqm7UR5TzpSpPbh0img3XfNhUmlxzhm/P/v4QyCNRrAXNaJ7mhLmhv1qTbJ+EAgR
UY6WjPCCbbj4rkI33SmnZyUDoJihq8UIgWHe5/XEcOZd1ZBlgmNblIsKvv2Au3En
GJ4ZsyXNz3klw/ys/jUdZGmwPle0zvVlITf7fxQgx2xXvvoArcmOf+wfhK7mCg1a
DaZNwTXEUDaAy3mrLKN6doZA1nFKQiJ6sBiYc0sQVaRKb7BjO8WsmZau7ItQiJno
518TeA0qUWKr469xEfDKC9XKziK4iHp9SQHVvPAM3uOTlaXGOr78Yep0gFmVeTIT
/+M4j7DpWiR+m+nUSKidfWGo3qCoscgVeJA3N+Olbzh11k4LunPqeJrm1gY5gjs2
oUU/zSSI8EEh6PQVawryk3Rs0o9XadvexxeVRvLjsGucxE69bggo1fwFkh8MOhzT
f0xICe2RlAr1blfcqtjWpEzccWqArUl1oWqLB6u/S6f0N0gNfPAGcRBsHnAWaTUx
zUnR6eCju/gK5jyVYLdAqWsoG+AdSJJ7fwupTSiF8uVnx3b2DazvbtQyNpZ1+CAf
4g+Tnotu4LJZB8VPhRmvH1Wjrv+uJy6C4B3fo83D4As454QOAfNM3vpWFSl7ssus
fSJionFjZPeesy3GXufVImTYAEe9TU6ADLKPdamfCUAR3MaGoy1seMTvcDDcS3uj
GEfMyJFfpwCoNzaDUqAXUslYZFjiNuaJzakz8KWq2vpSpEC/Th0Tgqe4TfpO/whK
9I5lcLKTTjF0K1lp1Uc5dVzzBgYt9mcyx1StzEqUur8aIY+l1VSyT5sSD+w4CNS6
p/X6TcO2EKeepGIO/hhmYkhNGrrID24Wwn7h5qlMn0X60NUAT6EBYpw8n2+cZxzr
w+aE3+2xe9Ry0oIsZrKQh2HH45JvASc8qP1/Fff6DYc/Fa5XEumg3pVkkB9DXGuE
cZ+Xx7sgD1GHEkh8wpORb1Y+acUAJjRc43qg+5E5bYLMBbnIF2GpxfS6tjuBg1sS
MlcBuW9ayKBNsTO+R6mzA9PRju9q92Y+vUQM/Iv4Yt5JW3/oBQkpTc1Bzwe9zdri
IiDFa9aJQGKKgW6rhgAnKAZk574r9dA+6fI8qtA4LXST1+UQnJXbldcgJGYfA1kZ
+eE7upYZ3X6NaamQirsPyAf/ehP3rdWgLDbqdSFZZehnmoV9cL9mOEvmKBDQG9b2
UpmBvUzdk2d45ASu1YhbWKj02Cg9Z4Lenv/4paMvhoqX4z23ZZGjNaorToCZuLmR
6XBcQeuKhfUtVl1AFB/yJyrM4Ip7PF0HG6M9mZS6wm5KJTSjhg5jUQ4NMuwyueMT
dVL+U8Jo4o4RoVPbHMjPGYwMuXsF9ZayLhpKMnbGlXH756LCVXqQYOEh/LeeqSMv
AX//u/yrRuJRz79EKLOzDOqyqhSPDPekGFYeDXsZaxIGr4eYELD0gU7UVh1tTXJu
9KRX08lxcpXAASKH/O/DMdhVQtqcktWwckuosRSuwe+O/O21TADFPtidWqS5WcZV
qz90YkJ0RxHX/PW2ucznCYT6L8IFuQgU4GXSlJHYivWrbDcb+vrSfXinw74wyTBg
0sPUcWqMkWGdr6Lguz6Rhe/KnJvYJzEnHEWepD6rqg41aFiZEK1Mmdk6k1tKrh5g
aJvOQhqrvdj1jvZjJ6chthgXjNQfDBdDJk8wdLpG/CO2aIER1k4dKHkwHYkY2HFL
iIluVM2GSanIGTb2M0uNOi0K5I/DIcNbevMdLhZh3aRVP6l1kWIAGw0xno48aT/q
DoXBCAI+6Xi54G8gOb8sNXh2xLedF5/ua1yay0CvqtUfaVabkfzQSV6gI3ZGGIaC
0TGu/xZSsK85j300zcX85CkQl9gZ0yi6kIi2Ptu3vi77HpAfuUkKAoVxn2sRp5y4
jve8S7jJ08scFNr/mWlrnO/qnq0TtdDnhVAIacGsC1PozMxzeYbGimy1nsA1nc8G
M5noG1fhwHGEUl2QZZSMMtaCNuFmcfg0RwdfMbQjdf7Yel/+xJSaF3gkau3lo9yq
aXItlDVU+tepELKHSB4JnxSnBsPWuJhaOJHgV9Bnn9AxPkGi1IRxPQfKqoBdllIY
WhJVcWQkwv86Y/8DI7DyLmbP9rUNeI7pG9WFyKQc7fI0IkHrcyI12No3x9bsEe3Q
GOcjZ8LQvIiS8F5KcAfK0p/jHRrXl3UwuI7NIDAaMfj2m03vXiUwnPvHGfbqP5yJ
rfjzXET8owbdl8mkjFOkrEYzVWSfrn9FXxKDI/q1JTLu5748dtIkPeShMpJ7Nr03
YCvkDkJ9l5dcKjlsz/CfxS+oyRPeSDikCLr76KRVRRU7y5ccDADO8qqc71E6Xaen
dlVG0XJ5LfrUXHmefrjVrtMHpHXjVmN52AXyoT+MzTZ1Q/Xq1xYnlyI3CLKmp1Jh
Fld/Y7uUgbKAZMoWBh3hbDU/3vqu3Zo1SSi+mvx8RHwoh1xgQj3JDVYmZqomqjMW
9RzeHCvMh+QYDMlMvPISOtANOHRlufQkUXgSP8jih8LiEDBIrz8ErnxduemKLKp4
1yd2rhmPBP2cg2iZN1oziVUIoOPF5KiyMpWLamVG+XqzsLnrU3/VQLLaNQvLov0C
NfeJJ+Zj7aEJM6zTCAf4eqU6Mqrgs5J8F62HI7hqQ1sdmMVNZzmAsxCe7CBDxDT2
DmI/qPRLZrMKVWd7JKmaKPNFqnTSchOs+d5cfd1pB8adbKdljaOBht0v0vzCP9Sg
3FXrmcy3/TzxOggL5zqcNVh3eYCeyA9aPKraSn5aB1TPd39b+j1Yzt8FHWAxmNrH
rWsov/lvv3IDF1R2HuZSUCSPy5q+wilf0kNhGwukOpvqSn7MCbx/QqbHCyPc2qkF
JIipp/ztjQeLxPHiU05PV/dkXn6limiE1iAfR4ag0/Aq+TYUWY7pVrYExe8VMo+H
FVJrL/poCfUDFk3YCQiO21NEGx2Wv2hBQEzXRX9h/2a5wAch2mwJCfB+YmFd4Ysz
kncyPbsyFMJWjMbplCFMbxFLzBmVKrxtYjb/2npCSRy3DHwn00eaLCibQu11yhrz
qQG5xVGxJ3phTP/oJ/RasG6mrtGteCpJMQBIgiYVbDY90OwZfPOvAHV+2GEl7Uh5
TojcDj8v5WMXALLmLP9ZCw7eBSBtv677dprbY1iCbI5gdpSj8PoWXBXAHkiD0qt/
l1kd+M++BuTDCMhVSdSXfc6agPmajJcMiLEupGAGk7l7jA+RI27hRCTXgkinG0XB
D8s6bitysLlG61G++Uvt5Cujv6cmnCf89BDk8TvUWwPP0oBItpNYvJ5230DmpF3A
JbmQJKAteNNkfb3y7oj2PiOziwAJ1PBTmwNojAN/oxuxpFQB9VWl0Dn618d+/oOl
ivWXdhmVOKFlTDR9xweaod6O6xH634nXz7ETNT4PDNlFawr2vsQhtq+tu9wUaEpa
UbpcvcDWbaLKC+7a7VKZApglIf8op6WuMTuCSB98cWGxCL6hg7cdQcW7GEhbbsvC
lWVBIIzaYQPp1xfdCDRRKzB8qydghhJpfOKBr+Pohr+V1e0KC04yPaf9ZQmlxamQ
SvyeqEaEgi9wPOZgfqzjEPWhJPr359Bb7KisXnah+2getf78uoi5zBHkXQ05JXdc
ZyS8tgtQFbgGDV1UrOJcCwO5oOZ06CTLH8UUH4FcEvuPLVZhy69jvGKENcxZSp4r
dJ/TSIQdZJj5mw2GJsww1BIu5g+pcqZ5grroKNRNCMsxjSBPdYB45NE7RhRWajIL
C4esP0oSIW4bEyMJwvDqe0HtzFjtDN9XRsA6lslKPdfi2EB39DifGdcEnrr5kEvO
9cdyunYDCYeWAG9GGWza4fSttfG88yYHpwJlsAzKL8bnDZAG2driAqKYRL1+PdJJ
iOANs6ZT5FdMJ3s0QddAQncLD20s7129XyQi0jhtYbWwLwMtNCyag0g94gT0ApBa
khMWcsgaJUZ5mPlhjOiaQMjlBf2SHfUu7mu2ykc6ztSsGszkk9EoPVBrO3T0WHw0
4P1th/nyUPQ4eMZ9AeOBJLzj5FQmk1+8NxU4VYk0jZ62aeN/1fMBPVFlVa86sWXP
mD7DS+myNUjT+W/TZcbFMkplijnhogCZtIktN6aOUYGPHbPz9DfEUvee3wCibd9+
G7IswN23q06q3PYwaIwSqzpy1gSfsO8V1O2AXocYpH5qynHxX4dSsu31ahLk5dVD
bDKp5N4cymZ125RKxD7voyWl19fKKPIiXKEaza5YT6nv6BBm4ztJgDJZEX2DlIFU
BtdZYccTVrzpPgzGXBdLqXjno3fyexcy+tEa/IKfL27jKNs+bv7Jgu00d0PSwFUh
xer+sjbJbSZ371pSHbTtWCYS/oKXnqbYXhPlpqE44GSf8LvRDwtsdbw2adHaYHBW
OmPwgPA+ZZvzNPRIHqNw+6AW5noRRlt3euSEDw4Dj9ABI5hmDNOHeXAtIXKyNpmm
ZTd/D6a1ZREDScsg2w+rQCyrfIQywgzpyPLXk3+KW1JLfEcOsS002xPvngdt4zqF
WXneJqw1PAHrwZpWG6KBXDPfVuJnj+o042EfV3bgjeH/JDGrj6+2Iq5kkSOTgxoW
UZPZx/SIgJ0fMpFfzIveQFP+62NyvPiLO0Q1NysI9kQk+0Ga8wWE33PPQ7HyGw5S
TqTdCDj3KojlkYw9IrHz2nSFt/oXdAN4kdkGJHdFwDKUgXLm2GpRZ4z99XkiY9dY
QqLKDvQlxUDJ0oSMsr3QhNEF7fef5L+8RCZ8mrn2nVFhbR8bSUdfL+jbTz4crVa/
xVSoO1BEUewmZAbARdlXyJl0j3ypf8+ozecRBFeBVT89J8/amEWtgqc7PA1Z10L0
/SrCEg5IDXT7Kz3G6PBOjqXrj3W+SvOiwAgMzyyxHRYtttnGG39PxuJQtjVxfRNs
xlkHDpdzT2IL+iA3F2DZ7KoHl2WkRFT2AdYiPkL31Y0HQOnrWRokoICvpj4r9YQp
PFenG9kChJ8Z8hCAFJ5oEC6EH88Ki6YpiNhr3C9aX8Q9GQV+wPuLDXJgZFU5jDSh
y3Zs1KPyF8dRP/ysbR9FYIobdbPvDwvVnqiqNpkJ+OYitZ9SvTJFHkKfkh5Nr/yj
nsvCCjhcOoS50W83AVknoEc/DO8ClJU3YQIsFcGm+at/mos8AlonLAmFsZDY73jN
RdPyYmL+HtC1yZRNRZBZa5jGH0L/9BP/zRrIrkdCp8pruSg/WvXA3YSaS0H+G4oB
yX2yF1kslP4261/iCNVqodnKNVtLnJeTX2uVwBg8mIBTS0Gt9ALtS4HqLaIT0MFg
N+cw7X5cpJlSa/xqrsFJWOrkPZYjc1pMsnwtITB0opimV4K1G3ZQGkCf54xjwYpo
JZf0Jz/HFIZPvHwWu4TzfvlvIOroluM8+avgidVABfZwn6UXgw5CI2NGMo4etzsz
EKVMQwCPG3i5oclcttnF3lohTng/CN5g26hCpWfK4lrEnc2U+7pgl5KWT/XviUoX
KRTt6AFR1fq8CbCF7p5pyeME1r8RWzKy+rv74PfU+5Qk+SOj583LLThwEfFAUW+A
asiri6b1BweT9p3vcrBCYdsuzyONs9QuQWU5bvpDj/2XxeM/fkhvzeZTXlGz0qkO
OA4Ww3iENkXKqJ9SGFoIms+ieGFTz7yoj31oReZtuKn6epmGeHcb0PPl43JWHEGX
3y+gjt2iLDuZowwRSvvTMrLdOzovCtRG/2K+aOwwQabjPHCsmFO1PFIDlxXIYqbc
8o1IMkrgnBktuqSBQy7iDPio+be5/Sr3atJhkaoKMNytV98ebNYRdnp6Z7rfyA3p
iXze6acGOOF0gxhsLig9BX0gi9PLdO0gvAPXN8Pq9kwye+2lywo2/NhWz19USpY6
/aKZErwYhFnZunY1JiiJwXVSaLxEez+pYi4G5zLEL8PZgyExKC110gs7LwYgvSGo
F6G4c+dQbVstQk4ZTJ8HGZZ7bJL15QhS/U8v3uUZwAYJJXtPexaIQt4O/mJKK608
ZTvm6dEOQPPWV1S+ICGECX428CQT9zvYdMysJGp/Dy0oHaAUKm9dubzXE+f5tlK8
p3TkiHx7INy4QrAu0a6NRN4uLvtchmGC6khCc/HErXBTNl9OMXlHmdBRcGDwZSZ0
DhD744yvvB5ZW/J68Il13O4+9i948z2QfSYmqMvFjxX7jcaV7lrwdkVG9Aq2+zyy
W85YeonUjcRrqt0pUadkjUrL5CiWo/8XKb+YCjy4JoPo3lgTgss0ZvzxAJXSN/CV
UqC+CtkbQphTwIdze7ykLTkB76lUda7Bdp7V2PdSx0qnOmStPtZfn5jYnpzRv/yP
0+7V8mL91WS0cEKTnsSjXzcyBxYhOiCS7YdnfrVUj/EGCfiEWVGp5AOkR/M9fA+V
ueP8/VgsUkiCaw5Kxs05YBK3lFH6c7d5PhQc+IRAqdg9h/oy1P17B9f6QC/D2ZFK
bzVwwedqXhLZW/CMP53F7atweyU4uqDc3Jp/U7NW3qtMEt8sxqwuS+NcQGrq/dB4
3g2McUB9oa0QzHXnOITvwlYriqUTnFkpxXW3xf47OICBvpLjIw8PiC2C0hwnG5nB
AnKD6Az5df8cxgy69qW3xgoeaH6/6eEmn6ellEt5RMZpy6YfQ4bOfvT5HBaZ9QZa
gwRu8NbsGeLf+rmlodFuM5uOlqCOF+UGY7iDITiJvfZdlBEFUOC+lovAlm3025yy
f8J+EkJjroJDFtqjjLTUXmWDTPboq/AtaNZAIBwt7f6vmHgD1pjqnQYBlfyoaDkX
vD1t8TpkqU/P4ckw4jO4tfeLw0zg5WX99M60MrZg1rKF7RgbeSX/OXvuH1fYO54W
y4KrmvwIZcfcs9l6RPGbgXaMW4QA3qumi3AZmz/W2yoJ+o6pEUsJRiRNtwsGaec4
oBlObrHwzaX1PTu9eAKmEzctjTvtmOj19RXRwBHTpC9VcQ8/q2MnBgG1Zm1YmIZh
w1EJoDSwJMFKKu9a1aCfR1OQ1/R5O3NL9TauSyvCutm+5Ip1hq0vHyFq7HWGnxqq
NzEdNY9lX6/MKeaoTlQGIhn7RXDLzLeoVm9QlGn8TzjCN77evPAo6bCjDBdryk1K
INRZGxMwyzudlRzolW+NLUD45RsFZPoc0Svyd/OHvaV5zoU5PxH/Yb7p9LCXKFWN
1n1G4XQWOGfAmGw7hURJ/T7Mm549a68lHabtQnVMG6yhMn6NM6JjX62uzD9w6Fzv
5IeR6sSRAObfa/omy01k6P5oZhf5CZGHaVzNmlG4M3Ybe1pwZWPhKuqayLto1SGA
lj0TykFYNitVjS4V8Uf6/kWbI6oI4wY6YQFsgudeOwld8bMdK88U1A6owYjS0hEu
YUGE9QHf9PB+MEVd37qnbusm+PAMAFEmVgMID0jwbXUXI02OeoPCqiRi5lfzzaLV
39b+04SeOBcaI2x2E2eTSsFAMTxSk0/6lgzTxDwlBgXrP7AJi096vJdQIZAMqum5
cxv9j3a400tj78VT50GHKUmXRaF+0gQ+heqCjT97RLBeB3JwwsrZCQ1KuwhrwdJd
8Qps0pGwiNJypiNJ5Jm/fC+kw3w4IO4j3QaNlKE5DrAXylLuAqVwUdP9RO5oVciz
XzcRn7Bo3qXAkkggYYToDTF51ZfkDkcz09oQvuU7yHZOF7VJBAWPF7bA6gnBnBxv
4r22c0VPthehAOyU56YXRClXD4D7ZeHmjEOx+KNPfqm5d/SrkSDD1fYY5+UKKhVy
qTA0VClFT7BDyNbnQnK3CQxu0Aaf5DYbqnnzj05Q8ZRlwKg/waIgZL7YNr1tMQrR
yzbIwc+Z+nO9kcCBXMxmpyaXfYlVi1WXUZ1mWGQgn3Wmcfj2YLnwRzJYuX6Enm3M
vWSe+0MD0DmYQZcceUvDaRCZWOPfMYcD43j+eVnZzunLSYuxbcR5Yvq3ERFu9Q7K
dAI2vaxWuni6nR5TZqybe9Nk58i2eUOOxctXBSk7mAvUpHIvusfGGQnoBUKydQl8
rcP/eKvN+KSaWKbNiucGkcviDCPEsQSQ4PUtDXXEqqYCB89g2zHaofFBFCkG8alQ
kLi3AI9QIqiD59UwZZ+vblUpHT/2/h7tgNluNTV13tlBUuwt9PLl/lZ/HFBfC7y+
QXHu7kPgHFrJbCQZYD3z/jDjE+NCTWZP3VBSBoY4f940rQnUCdUtx69fQu8Mmq69
qvKX2qCc5hhkOaFzgGQVaMjeQnUB4alxHbY0kjEnTOY1av0nM5cKoMJrLfDRxdcR
aHQNAKzbkD4f7MYzEv9rJhdVYgWQPKFruZe/0+CjTopqNn+lyAvE5ru65SvVNgko
3NcBDJ+sV/B9pkZW/bUQPyHBazfQOSkgTgAuFG6VilXB5S13J5+AgGEJrQNUo9+L
UeHjS6H/s30mY7RByW84ENTM11OZtyiFzqiboExB1rADEz8Z4YUar9J6gmJQnoQP
8DT+9B8pCzOfNqxrZu73ytV7yhuxfKmv2go+k0xz0TSLRjS1UL1uRoFMbUC5AgPF
IN9OnxtA/jvNfn8POd+hFqrM7nk8NxlCHBCL3aqcvJxDOltgp7YTOCaFkQI/pZbI
NFGMLb6I4GKT6IFG5O25VPafyIrMPDOEQ28bIAI0a85CplYiYKCxtU5DhRMypm9X
29CtGbB0ceAbdXqakLksANQ+aiLXjKTxEcQOPODtJrwH/Zcf8jX07PBgyIoaDIyv
qPrYl0Se/cq7bAaLqqO7hBY32H8fxzFzAknsuy6GtFpgu52dHLYFDLm1A/WG3qMU
xuGLIvpav5k1e8E+5cw7mhvJwBQU+l3FmS/dO8/8+VnvTfSCxHTOYUw6K9Cgaahu
G73LUCRTupEMDXA8FozV81ssJTf/2lRNFKv7/hk7Xrzb5hhbGZowRZ0qQ6m7eqMX
/6vJVm+LhFvhaQ9OpySUCTYCbC6fEm/KBBdP/GjLx7/KyPi3v+3FfdTBwGhmHozQ
O+zQjboPPdqva/tJgQrULZREEolqeBauz/A58Sx7pnC7WdorZJITgZZR7TR0Jc64
koZgvm1vU2SkdMkWiixqh+gTH3z8qSFmUQm7MCl68ARvg3px1PaFM/PnPX88EgXq
ExwghOIweg9OQMI0yP2Iz7OxQ2j/jz5CFSV/UTCEsIH/YBx54MAZoFtKZm/FQoup
61LitsIVYJYFyQUb1LLndxc668EzgqvXxwsRjOsKqvFekoiRXR4V8KRCnXfJloBu
IBpB5Xuv9NuJkF61Xal8s9uv1c+MXsZ5DqMYCv5RGq0blICgpAyEomYpSFgMj9EC
KkSyqDm39XnBs/HrcsBb+OyxdioNKnVKFzL1ANbr0d9Pivk/EGvtAu6FsIHPXtcd
rtQ+XxpMrhVV4Zp3nHezIDAKAVpTFWF/Z1N+IFAZP/Vt0xRUNv31GghCmx/TnV/a
dScayJG7c9YEyeehM4UE1pdZKQYjxlwxL3YQK3i05ub9J06Mje6bhma36hAvzScL
YnDHUUnBfxIACakSWCMmGFhhnB52z1h4AaK214J99N7kN9yscJe1UyPIIpIYhKm1
1i8aQ0n2wfjq/5OI/YMDudEoozae2rx3wa2dmJ4nnU4y8doSYVK2qGzVzVbRzAaN
jxaQoLWWHVXLRQWCp8w2rw8A8XfcKWuSoVUiO+SRpLynsugXpUb+i3Rl8lCijwPk
ZlIJPNFK+0g4WhLL1TZ67ettj0h2cOhuCVHzmnxgKUeYR9yLtSENdaWIbJVY8y6H
yqPAciongkU5ju8ecqKN6RZC+brHYof/fuLXV/7iJYlZ0RBI/H+oWT6SDJyEeSOu
1HiDnHp61m3Ap2mXZyVA7hPWG0bl2WBIi8gqorCNRNN4xOdxOIgFKeVPvY8vwrKl
3GFHZs8SNbGjBoZWpfTW6/PG/lrr/bn7n5X8Z3gZD5Tufi76oyKXB+bmRnb+57vX
APzvrpqivsWcVJybu5RyrNPOhTFbTngANLAwHgLjMLkXvA689DPlnUYkk5J2H1zq
OkaHyv9uOBdiEj0z8aX+1HPvNofVtPyNFF2xkdWHJWzTgYpDavmkymUZcbk6EQaU
Z/zldleCfjppqojAzeg44Ns+RVCLnwT5i4oY1VUORcO/H8bzW1as8jc6bVrP4qpm
zzHlf1DY1nNZGGOCJaT3jrJVTCVRVys8mNMOT7bUR9mL3ypxqzdn/titCsjeR5QF
Zw5fng/MMqBqMfYVQ7LcLcknf+K/seej0tlr6mNWQBpaHtdIVCVRG01G/z1CmzZP
qaAguJx6Z4i8A8/KpbpzCh1NVoFNr4Ztq8pyp5yDPdZdHs2G9cxc/H5I7UIjHWwg
Y0GCAhetQYWCtki4RjFF2ruflDtR0PaM+vgr8x20c56eq7CGPJlNwvnaXjShBCFX
j7VPHyj5c5nFg1leRZAjMxf8gQk2qjWbDI6yNABVBK849bbVq102SEmWRcWb3e4q
uq//BYaBRBsOuFdqbiahijBhB2OdQqWpg2ZCYiP3VOLrkatXPSyA881KIw6+XOU2
UanwqclViTh/gWyQjIRkv2vU9Kk+FyrSv8HGtq71lVt7tjq48wQwlsl31uehxX5w
WLkbDMhnEnT6XNtVHqriCFjnzZ6RNihv6eOYcSD/vZJF3s6zT5kbVaTG0Cwb7zbM
/Z0vmjSzDuNnNwzfAPRFOESS05rPaKd4r7PEETum2bSTyFUpGtwzgRQQXjT+9ulp
x0B8VT28IyskZHcw1+EKfZsuHiDCDH7ahU4CSUBRI3f1U3ZghoEZ7xmSq71+y+bN
7v0LOnPl1SV82LIp4cJ9IHr2GjdhAof9DFePY0lAYd9/qOsnW9EdV/M7kSx5J4te
eYsrlTrJoMrbf70njUGTYYv+3Zob+gO1S1bvuItNmwS+HAvlJd82wuEQ2yULffQ5
jcCiDZeGXry6N2VhRXnLTLakwYlott1m8P3nvWJFGhf+YCUEPx7ymGPuiC7Qyr/f
M35MZWUe2bdXg4Wanz504AXHvyAFuKNIFAbczpgTYlsWVVuMyzc50unJbtQbgHCS
r/UVkCJ9gwWkIao2d12MUNyjUukf68y15CxBXwo+DXIfBw0gF5w1w+N9JGlplhie
lspCyvnZFsas/9TLqMvjnvHFAhYzQ5OMnm/vbovFbn2CzdG2YHPDhlxpY3qH0vOY
j7cXjzl8hjewXftxpuFodMig/wYhYJ481nr68BMYp76GcR0LKgW9OK4xxrNrlwLz
kM3uM5ePoKRSrJi5CuLTi2UKZ+Ed2NM6XMaD0dbh0F7z9GT6zMINwVp69cie1gAq
/tsTsRFIJ90mVwvwuO+auGRiHbt+x+gtK1shptpFnOPAc/uoLm4gB3p6G0tJlrEc
xr4dtrkVJp3A2G9B0NsxBW5qrTHfNzKEYB/aLpu57xyjsj0/PgaoCBEtEm9mEc62
McJMBxotBwOYBUU0Y5HmP1TdbBdtuKxHZWOrfFJypa2twsXltHpBml8sj5wUVv3o
JgwmonyIPKjo+hWkQdPZT8bwYpWf0D2LJJeTnT7RGLjnWRpgUNX2uH8Pfwnanuq/
r/k2+Pz87UYs7SGrf7sd0dJkuKABMrm+scEqIroW6eQCI+wkMtkH+AN9JxqrwFbo
Y0Gnn6H7Yo2ffTIO6eD8EH5z6aPFoyOQl/v+2pvoFyGm3dsjBik+Oq15sVV9GNui
f9jkpaQMJlYjpEacCxnBZSqpZMQGtBmwnXxBAtPMlclZ6qTPtSGFWDFXJluqDIIR
FAwICMdVe5WRRGiee7waVOaX2FPYf35iBBVGwpcl+bFnSgSizJMxQVVPEBzroVaG
4trf9aH4cd1hctp+4dN1w+6mVM7qvOfFlgrT0lKYrdIYVhlD/5W83v3BGYeM3eeW
8zb3nACsQ2OQusVDrzbQBfizeWg4iqUZUslmP5mZ0K8DfOBfhr3XOEkmeX5dvtmK
4Engva5UZ5WA950p4iTm4YJO0LNkREoGaYR3jPRou3l92/0M4+Q1Ngwg+K8cC1v1
CvwSHaneSQUulSRB45GAbhaHXC4oMYtctDGq9rf5xpbETKkyOOwNwS5BHo79qO1H
FlrJ7loYVQZ0/KitR4S8gnQJ83yn/seKztdVrNapscYrbW9fCUudr/6xEkoFyuU0
pPmXh/zdRm4Fpq+z/U9RbjVFFDt5oT/6ZHQw0o64vHKcolos8BFrm19bH8HjoU0b
s9S6bGxNF8AzhWi1a8snjYjEWci3E7BbnPzoA71IR588Br9qw0RbPhJLgGhX4btd
wQXpfn3QRdREJUnhp646PaAiPjmtzoLvlSAydCIxGk+AakeO6hNwdi7Gat/+SL5h
14aFHDMVH3jBGhDXZjm/yszXNAmCiwXWacRH2zVP45kxNfdrjTyyDrGTx4y43t9R
Ad9NLXKGtzzGegY5QoYKFPdyVHURc/HQN+EzVN1eEvBMUdmN/I5+30NNqIiM/ivA
zX4pTFz9INeSIuBYYteDTw0YKAUSVVMRQAtiQY7jjbucoP/s6KClwyciBgRdUt5m
w2jCNfk5I9yybn5cLQzLSTuukD8112LYGzH9rw6o77Z1g36eEabPCem5/x3dQta0
BzJwvUP6qfVYOYW5mzLG9LcQvmLLjL/w7wuds3xKAg8JCKSlO8SYHPKfbnya5vJo
0C7hlzIKCF3VYaH3NJ9PXQU0qN6pK6gURmtGASZXlow/bmdVFvgdYWsiawdNzOXZ
651GSLF0oPN9rqk9BTS3HJxcxifq0fbwCVoqGHU459qbN77hq/gbo9pFg/urYdKP
DCWBhkRaQS9IExdltbcjzSrnAQubVVwZ6oqu8x3klovYuR/lfpcKx4jRc+PGjT6x
RgZ5LWmGJ+GNN4Qyfv797sUwjRQvGIyUhmu3hbY6esh4EDnvKQXob7RfHGyF93el
rn4e9mmzLawH2hrLRvBQlm275VBKW32phM+cRIbrYU7zUPNrfsuhGZpIODTOefkq
HygaAx+vEzMjd+t+1Bj35tDryFrlsFAsUywPPM8Q7HUH1w7uI0rxOKo1XydlzGi7
Uzpj4krcJn2xkzLThCdYSyFVGOGAoSvfWwTazTWzl4wmwsRwcUsog4liYRxVtm9H
kCkN1SS5YRsMWcJp2/9exMsfoDaL6D0ZwR3O7oiYK95E7c5DqXBA3HV0qo04WLzL
851DiunOegXapk/AneUv9MBOwLdCxFwCSgdj5c6eQeAxG7vS25gLR4lQPMD0JiEY
kuYnCaeoPMlftPwPd8C2VIeHuR0mfMnCqPyLnBJwNDsXTSD7WujRPRIkIQE8Ycha
TWPMKzuxLfAJww10xP3otmD7Y3F33iEvvGO7bv84/lwUdesmr0D5aCnPnkQmV+ni
sg4BjC3qLiyYMGcNSSd9oyldfyKA331Ysmyr2776iCAVny8coXVTfpDAwu5VtajF
zV7HOArTdymXdau3YZCtDL22ai/sn53l4WzgBa5p/74+ONTdWjJjJPkAuLITP/Wb
w+rcNurMpuPFhIas4v81CxukVmgbsS5Ozoujcxa8fkXdKfuYdV81M3PB9nLrVOlc
NSIXav3n9oHuw2rLKRjg+DLeVgjd5ZahxDYRFiAfol4lpOVE0o0bse7pMntaQRjB
DIJf7qVPzdxO+d3dHv4wIb6Jl8tM3lwqQSPXdd96KZyivDeGnFDzSOe3xKU2r7Ic
jMf1w70Ia6IfaTVYvBV2lN+P2kBQYA+ejVSXwHAq3Qj0SIzQkOE1EBTTIjWO86/m
eO64lIiTWb4JdzsNFzUaEW52Ti+dTHjQwYR4yk47TUxBa0qWlG1FuWzDViElfrSU
RKpQw4QvstS6iZrocyszvOxl7BzihDTnXHjhNgoKdzTWOzejh6S32+DfeRWM+TaW
uR2nUp0yw9byD+6WBBx/9gZfh75Up0j79Bke2CkqCO9ViP2sm4rb8EBvZ3LDqTHE
VeXhLPoOWuLZJyWZlPUOPSPtaFd6U7VfqW8frjo17Ks+zjM19b8DdVdRWtPS8ezR
NpOqg7u+fa+5EwuGNEHeMjxIVYt1fsjVmcETrmJQmgfG0JoROUznPq6MPLfodaEC
W59PmGv6aqAUQlBzNoAaJKdn8jurcKmcsRHpvZ/c4JPTLBIooumGBVu/GAmIghi7
ro3Bw5utDJu6t+0g4nPanIbV30B9ZVzubN7mb9bd4WjH4XAiEi0jXRjYebL9wCZf
J3kf+9X/wL7gAj3iRDuNtekZpUuxpwIED0eAS3AaWidEeXl9qp0s8X5VARqLIzuS
SK+HfQs1NvxB8Smn6pBOmynwSSNGZRdRsTppATqvgM3rfCma1JR0eG+nVmSrEs9b
yxp3UemhYnh5WUV89qg67gpwcOExbM5rxRQI+UZ00ioWobBbSSAP4c/5/nV/12iL
o+tuHr4x6cJPUnbF4lCq4ZMe88G+NTZ1aZSXaRcZ6l6yzDjokqIsUgvv05K9bK+4
2p4dHndYCgTyF++guxnOFPPB6UCPfh+zavlp7PkuNlkWVbUdXbq3QNgGLTDYi7gu
CzxqG7xSfagv8ku1LsEpBtEkw5ddb3USdp7vBFlEOe72Ve5ZUA2wYzftgPUOjgQZ
WJdXsYKhuGbqYfsl4B98Px1/OY3lZsn7SLdd1hXCoPTbS2kIb8Wrt0dHFJOWTWsX
q82eh2/J/SO7AyPF7GlZMDxDqbBKdeycLDEk38NoYyNdZkwnclmQkWlnxUVX0bCM
Binh3Y7xtQPYr2UcAy8Jy8Jn2JCCQAWvrMvxtzfUwnXCY1uR3yvtMdyyNj4exGJ8
6PmxwmX5QnujjCWG92ZZi69Z/0LclOuT6qhf0v98yQhrsJY2GuQG79PQYxaWGdpi
nD6nQBAwmmR1tz3vJ5BKYlA0CTocze9O1QwOGH9kDNLsqc7ohYthbU81ewcz78dB
Z/LsQYfzVXXK1hoBc2mtyRFBoQEeXaSzBSVu5CMXvUBkqrFW7E5aUT+asFU5Si6t
W5wMv04hkjVJsNAIskq+E9UxWAm+cOGkVTvU605i9R8vDxmY6vepWb+KI+28uHc9
5to0rjrOIjz0B9rAbuE+zo9QLNo7JKz/TFklt1hFegjHqD1DFucww71D8jnaRbXQ
ChlxcQ83sVxBMGv5Cc7VgmhHA/thY332A+WawfpadHKfgEXX0X1gUhOh9/tZcniP
D+ZNokhLCE/cxzDoixvrnmY6uwOO5tyA4zUJG/W00gf7OV/2A7UxzR3Z5eqPY3o/
g8qL2nKYVTvHA4suNL5OamSw488hAnB7nFnCZ527m0fIrKEVp+7wERNrWultYxJA
1hLKX3Us+OYsj+345gY8F9z6kYxdI1GhZOgg/GVZoUlOPXrGRqgsrx2GBcub3LC0
hok4Rcex7hEzvIEzHxLZb3IISgYY0M/PL6YFuWM3WrWCq3QwCR5LJuPldo4GHQ77
QeRcWtTTznk6VIZsJVt0wT3xtCMGDxaxjct/BSLV4fGCSdJXguweLyqToUkKQZY4
5gZC+7lROty9bvbQN5IZhmvlObozmR/c0KNmKgvBiPsXHm0coDAT/GIerVr3RcRR
WlNHMusY840yaJSQM4FOAWjwMf00OWX88udxFWLHaOVJEVWiF/OwxPcXV0cSQFVM
F0FOdS8gNmvFLOHXrRfndh9GC7M1icbPPlQbHzZM7xTXUMx84Hjxlee2DQYcfeR4
B16UD9NM12ulsMAtWaMcr0Rv+u/vhYebM8SsPi34QAYZe5+iiKmK7lGcTUEIQ03r
91/Rvu01hOuU89qZpPIXvlodMhZXjGKw/cLBuKUhdvaCJMS8xXRrCsDb1IZWwXAM
nF2Ps29/+o9RfKqpqma2euKe2ba+u7WwOiuXWRJJZQL4YocSK/5rUu+dIgptm9pz
CAwGJ3LHtn0KJQQnXvNgInrQ/Cn8AP+WDXzsxc36z3lXyR0rw0F+eqC6sJCX99Fy
vdcoL8fjgzx8aIWCaEjPZINZRkU9gDxyLlK8FzhWDCoY6ZcqUu50mr4izUhut757
jS5L5Z91SXGLwFhCTUCtWlSzelhDzSoa2Ny2NG85V7v2cpYpsnNQHmgByYBF0k5d
hoTfL1KVkW2UPYgjaCLSS4xPxYpAIRWVjVO5+rfpKBjq/AKlZTqODMGt7PWlqESb
b5RYJ/IJA1agjK25IKPPYF/3lkItiLTWvqWp4wFd35dkM6bURZ1O7Q06zL1wULp3
vZ/tTAmpkl8zFai7TZsJmvYT7jIheq77x4PKq1khh+oXn/xc6sMfwgthhNLVh6Eo
E8Icyt5u9xi2gj/9JRlr60oW2nAtp3bbbE7ztrbPq4D9s3e8zv1of+NLVWfMurSG
8Oso86Mu52GiTREwURAls/GLD4sdvPQ7usgLMhlVHxiVk0VnPIj1MEyHg3gRA97l
kPTLfkJLs2Z+L4e3oOpZDbYiD+fxKdk58D0Xm+v2dQVYhnO5SogCu8QkIK2Ysp95
exRPCLSMNe6hUqg3YBSd6iBVo4BDncLdTPh++7RUsXC0sJrVOpIC72E8Yxw2ApZd
jSWLS1IDGEPuWfIt3EAULm7kRQ3fbbOvnGaYVNn9nMObDRjQB82pHqX1PKKQly6/
Yh3yNoz3vL7UzduZPVBwbVn2WFCiwgpEYAZcnNKsn2w2h8vreyqibLS6lfXxMUbm
BVg9MJnxAEhyv0I2b7i/omEiFKO2+uBjf9gyzXW7q/4=
`protect end_protected