`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9056 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
yB5UT5oQgw999PzwDg9vEvcB0rfW+Guk7FnxwXE3uEyzsCQ2W3y8MomEF4yRASUZ
opgnzIWT1Mvvt3BitPnsXWyTZVRFPEJTOlCgNs3/cutzAFyHFX+MVcvFF5P4cDIE
lWkKQxz5PDsBxKcv5SQ0keLfBnVxOH280P4W/Ujs96qdACtqwfrQGksLDcgyvFN3
VoeaDK6TOas1Yw5QXecXaGxFVhKZj2XyxtS8aHPwJ0a2DFplxrHuDu5AVHCDl4Yi
6rJTIjmLYdUTm/C77nqNlSC2upat+5QcF7Si3YDbXO2H1zjRvBav5MJ3JMnXHi8y
1nhyqNqPiwAJmHhFTrJJzayKlunyFovWfMKtN95LfzOPYKUJM3KMx7SGMkfvJNGs
tA8Sq+HmeUrK08HKE9FDvyn5M45jlr/kdvZgcsR0Le916k7Q8OyvH3hZqIp9BSR7
WWBcxXFJ3bE2B8brqoqLHsazC01HNXP4pVSAqX1KqZsLdXO+H0Myvl+V7r7BgTKJ
tUm668mNtuU053drZTlPhnQQMluam1SEUnbKU3uVjJOgk1UPr9Xdvf4jJ282jUTQ
4Y/st7/vscMf0Wp4OnOZGPxOTklkBsznSowTzRohyxoQ72g3bmkc8GyTh4h30IO5
/P1i6XlvU5bAuZOqIMuF/oUhJhieAfLinCu5pjekHqTmKY9UkvSe920Cv+LqepZh
IIP61UCLyVN8pERKBlJSY3817WEz3lK3Z3QAnyWHWEzEM534oqxC6K0H/4+LEyot
KsdUOjxvVAepBcQrKJYa49lSia2IehxDXQhiP4dGeRn1jp2Tae+elqqF+g0neirq
BiTlivEC5hsY4eCGyci5CNP88P2eoKtAfu9HaKiOOKRAkPQhEvXzDj4JGTJkjbxs
aZiwCu3/WtD0VYSr9yx93ubc5+1gFJO+7WsUu/1q6zXyvZnWf4UeqHi94/pCXFOh
nr5j9693PXDmJNujG1SqB0s8jrrsO8HIXC8eZzKZw0IuvkCohfiEelmuKFKYo1KZ
6/Hu9XzSt9M3ztLEuuJhcG1SlXMoz/TkRBxCr2llr/tYfyMw95VsW5P8EHDfTlmX
k11LKyNmxiBzYpoqTdf1twMCR9SXsy4bFaXNMmpuph5xX9Ezb+T5cVxNczhx+KBq
L0A8nzs/1f6/07/r9u0AZZ/agStXHW5kZCrbVO7pSjsJpvvUBgaP2XY8KpKokSRq
O51b4UbPtjm7V43yUVcl4WG5ERBj8Ss0h9Wa7u/u8jk4MsXurxyHoX58DnoTesKN
G7zStyFk3+SPy0wi2zYK4tTdMjzjy9nCT7tF8/DynY1+WVsghgWIoxTLMg5UvzxW
GCq1qxNYyWz3UMXD3Nj5x8BOyIMyiESlWQm75F28FJ+otsRH0vgSHV9WjVO4zfl2
vlo+/MC5JKVWHEJiOK27vTmxucZ4skvVPiK+ZwG8+OFH1WyPCQruSrasBgLVkggc
Ja/U2f0OzkHQWNH40TrAosWnHE1jIuDCV0W8MQPdAa/23/cNtTXBl+t3ZbQsDStJ
0cjKswjMh3E6URArdWG6jqQoUJlYXSoLh9D/c/7jQefo+MsXNMHoT+XZiqvvP8TA
P11CKUMpbR1F2h381MuC+vgIEQ/GY0hAJ7RD+5Hqkgf5njhZ3CP496UAeUOIb+g4
snzf1GBs1eq8aU6OUJjg1lEoJ/v7kq1wWQkFQUNDtexJAOHzl7yeVSPiCTchIc/w
ITA7DAJR+1DtfljnJwedL1QW/DT13bMo45N9ZSYfMvp5T4+6dAU8skcJWZY3K2tR
LCKFj7q9MZkaxVDoFmmHj7D1YJPzgG1OWQea/wHhl/gD8pq3/c8WkX18YRR8MP+v
fHyOK3Wd/qyQaOSq+ADcRLm2NtrvUPeYqbBd6CKoAsyRUXwywB9WaYN5gSbfJUff
8K1+l1SgPYlg3I8Es1+yVUkCTTEKxeNFgkheq/9weFTC5x8pUC05dV3QaqNq0J/B
aKukSrGOLVxLtdtc5g2IZpG/JbyErRz+6kVty1Do0Gb+objrP1hku31L3ODNnRUp
2L9RolpSCOVXtTaz0TDYPSj/P7W4sVAP3ZRAs1EGtuOeAKfMMjD3SnqhutQtd8x3
A0sEjqRHokC00Y6EjGKyn6cWLICubmdSGyVcObTW7qfTk3ZjQ11CtdzoPAu6b1BF
b0OKohuRppOsxPrfTugwZnUdjmcQWcl6oF4aUmylxECAQhCfjSNUKMmSwUEkPBMd
oj6n2XX87vLCgQ3aIvXaAGsvEWRfr/oE9FsVmPMufEZX8sD8TWTLRIRI27mX/wa2
UIW4r7bPH72rhP40ARboRNiYD3eBJVEci7Ic8Qw711egBqe36dVAyhwKRYvrpctz
R1aVgQNDIdZLHdCbFUiFmd1KqK7EBnBKYPg3VnMC56YL0jCoXFqlKerG/hSNUTSF
9ZN7WI7fVe0TjG59zMQJ815XmUd1wLWJlcorTY/uNj4DhqWIfUXIYI2fL3wUDax0
Bd4kVfdbz2/IRhLG/TJXMJ9IkE2KEj7Xm6TISiILeEg4rcpr+XMKl5q8c16Qc97M
iYG2tZSQxWaiZDx5B/4FsFtwJYbZjQcZpQDTpQ3GLOmd72HROClp4q21D9txB7Vr
sOUJXTgXsXucXqAYy1UgUilpPbeqd36e6mXqH4vp5x17pHk4u1Olt5kXt0JgiGdM
y+Ezqd7KhW9pcwdXhyWgC5Jzs8kIaQVLHfMh97s4x3uaQdmtvRZJaK7yEVjr1IH6
kVWBEGr9UvuXGbKtT175Os1YMmHYF1HRmd8b4GoFKlMUzHSxBU7G2dCzCbiRsHPD
IzIcB390tLdsNofkZmihA4Gi7zbXHdRADAh1v6alEMZ0h8E8UhXkjZ6dMiermpUI
VhMmb9l79W+Ztz7q54jiN6CA0CzWTaTUvjkTBVgsds87YFojx+xFRl8ERW5UF1/0
OoG3Wtzd7wsolU+izpCbRO8lb/TPHzdGjL9M8oKgPREdWya6GtnIc6zBp0wPUJgr
nWo+MDOXyXFei8PxvKeK8/S8FXpkghPvwo0KDy0Yo4dhDCRHp2SOntl+18vEtvHW
2ol4CLBxOuXSY8DjSFJ5w4/cDsYmYHdEeFAidZee8BUk2D2djmSel55k7shiRqya
Vz8N+1hBserzJbAqB33ioQynVsEwVjDF9JwUEbUiL07GcBriMfB64Mwb/Ap2TnkP
1iDT9g2hbOv9f1hLGbfxiz+/aegwjft/TQhsG45cxKHH2rBTkNQqBXXrbKAp1Ka5
y0xoPqqAq9YjVyGDDlC/RHPPJhmI7eP0D/ht+1NsNSHN+q08WjlzN6O7tFAUe+JR
HkyDZBEZTitUmJ3u9ly5ms7U5jehmmiBGbPBKb2SW6qhi2nAUoEwLxWivEmIUGWy
Ghb+y3UR38NXJqqmRMuheUCHc+DYZYevon1B28azTvYWHPmgaNc6+EnQbmdZEqa9
wkFeIYh9apL5Qfr3HKtj8eFLIdvbm0FyUttvhB63/1reIJQxUaRFdazFT5Xc6IAS
4R1oNMDdz3sC0359Cv54exltNUpYOT9EN9X1DMy1gPFEZPdfZJ9VHdlIe0HKp59A
O6tKkXky/u3L7yUEQJ1ugGhE1dBVGuA2b1wlVe/vGoRfTczOLjT0ZGfKsAtFqV1O
ABAebo0pAjefLDyJ7/mKI6Ux9bDZ1i23JhvjCip99aQTofQ+kehEfkrsWIvx0mzB
dkI+JaVcuoe4AUkKaFx7J4oeJQJ7rz64DB9pCFpM8wwaqx6VoMxfS1mFpwEQY0lp
Npsb7OkA2E8X8oco7itxFVYuR/wv/zxCekRT+Pztpg2cKvRc/yxvSQMFR+JXrFia
FouFG/0jQVJAingzbwpwVsyfUNhoB+fSZAaMVlxv0ZElBlPDfTZjj6yR9/h8qOhp
LoroUTq4aMAZQkfB4H2rkV37j3OxgGoe0wtUB3QxlbuvJe6ctRakpHCikycKYuNd
LkUQPvbEzAV/s5gZN10qT1039ZQIObvPBDtRZKfgIFJLzbyerwLy3kxzH1v6EGk5
mQoAjGcPQl2JLcU6TfT5m1mQ/E4+OmdNU1AY6kdAEYvNbP8uJokhonpr5lfevncY
fhsFFzOb0W5vstbMBOMgNFHfDDres8GQJv6IJ4Vz2U+HU85gOwdPJGejqpk6wGNw
S+bxXshjfN0/nDh96CYUY4RWeCkK+j1qYf/OrAD1/K7qBDLLJcp8AnAVlhdgxFk6
8fDzMXRMZUdRDK062BfLqzXrqKT++KyxBRQaADvHP4yPh86eVTD3kWtNtSOMyLLE
cwMk1luSOutAxNfp720JD+2hffYZUThDauurwGsD009aoOvyM482Sx3uXRM5XVhl
Nq35IMfioqsc3eAbByfmcW5osjSpQe1VLeqAwIoro7gjiqaD3IWYeTvHqBy3g6Ct
nPyPyVPs/WDvQZsE0V09GgpfbNzpvOHE2oaUsMWofruPyzY5OA1yvFRWEGZ1JCDV
FYq//GK1YtAuWEQh9Tg0GZVbfnE44n08XTTmuPinTv6lJrncioPS4fDk33+UCcbT
k1m68VARY8m5h4wdDnIVrmaED2vaS9QDjb2lUMG47MxcivjIpA0QYegYlXUdOj8x
x98+5JhlH/M9x6JhIvGnqhNt0yXCvo6DE5v52TG2ErU9a8GdF53wgBLGQ3rG03dV
pSBIUGI/2tOcgj4tClnR9X5Lq2qQUXvhduPqpXZ63SzRl/kJnkUmdH+xYrNg3uVK
Bnd2Ef268hyT4kgsL6JputD25M9s0ZxNNIFcVFIlkz4IGnsZKwAbazyinbabDa/U
Nl0MJudPSBHiextXsXf9qbmU+BeJ4w8r1rWqo+B3LcAmeoUe5drFceunYN0eOaJB
lSDgRXxmzyeYffYPsuYLTKJlfMt0ACnN4qoLFeiUTyLBA5wkMYpmFBSMhc4RTEV1
18qkYgEqd5MDkmYN4nYk8/29o0pJpSi7bV66M5ONO5+MmyjdozY1XhXUQinjHtzL
FTMwhLPPzZCHEPMeY7jzhdWgl5S6LDDtaosIAXlCCP/N+mNhu43xMv31p9j16phG
hWjhNlLf7rAcL/fkMvgv6zBBN/E5GjcKYXwtK2M42X9nTfYrBVDN+W9j53lSKIsh
xnsxs8yezAWFNentUVYBgV5EgkY0WtiDAT+y1FNldPLS+ZFatcytGctUVWD7yqoM
8Hcx33hYVoss5m7BTnt8QaNbyiIx7Pq+T36hvnuCokyixUYl1/znpgrO3nQrQFBg
S3aRD5WGUqxZdhPJq6eqVXHwMiojj8UxZMUm1nQlylOFqPBRALlmW+2fgcJjb5O4
dxuWtFbtf/Jt59tqiWnQA6RomLPgw3c6yQxqgtVyt5avgt5QDDMzvFqpcupR2Bs4
oeXtLbeQDPmpkQ5pB76m7N7ITfJLXpvpYxbNBUPY/4HH+EdXA5n0iAMm8RJ+hJ1U
5oIaRKYJa1zI+l+lWtwZgpx9XsbCn7KuHu1upQDOlL69vwubzqOKcKLwFLN2Y9v8
zcu/9lcsBtp5Pc5Gil7hBDxX2ykuea/5NyTalBxrn5JumVluYqT3EkDE0pm3OU/F
Deb/A983yiXNADj10N0oMTQyiE+dHvuOSQzeJyxWlU8bk0+HRs1mGcfew13cC4oV
egqxKTcpdWy+A7D0tdzwXwvIqy7QzN4WknjyY1accNt013F7eff47PtnmerESVkB
lSJaScUazCWkHTQ0XBAp605dTxZxVxSyBWD8uNLB62JqwXBTFtlcb/xGy1boY3lY
kTmIb5mi059ko664iNlkIK4MPOwYekx7olAiN3iLAQj2O8Fn5InT3J7TbqKF0gRs
RSaJ3LwafZzkdp+C9gNdy+USDfXrlxmhVLtNDZO6+BX4FH87i1zsOCEcEVjvAqsv
X2LaAQNbV9CA9mj+A/x97eP8z8YO2WbaE7vaqhjeAWtQWBR94EVHQiLcz+sGvTzQ
cl43J9jGKLIhs63sE+lWGmMgziksEfQRQmLFnzjWcRx8MloBIBmKUUpHj5QcXsRv
a02gQ74Qyp4sYBAY7r2HPrjnP/6blVETfyfjDd1iYME/qrQvYlg4H5EyCyQzUTpX
Ym9JSCpG9QDzYU5d6gti0FEjZ+XDFzGk9J0yFpH7lM8sc76Tvvg4mFhlXrQ9+n1v
Y5TIHXlZLmxCEKWCKU+esFl4Bp4kk6Mg5rconpqAeWEe1VVZNioxWQWarPoCP9re
XN5xl6JTKcO75w4K99AS/F8tM16IYk3fVM/oS4a20+YJ5XtPPTbtVHfPBf2YbRHP
10EbTpuqWgDkqVDQjB11swQ44PoBSMbS+JVvZdgCev7h1jUY21NS4yU8FrJviquu
7Bn+vID+0LYjsRLRlxzRj6O5jpEfrDXOwTyIkPg/4Om3fks08aOLNEBR1tylXWqD
335sDuWGNX+uRHI3Xpr9DQxHUwhNOaHwuthSUHiMvbmd4+zxXmBSIj3MApFaalpD
w45tC9hMQ8L7+agEc+FnNoPJUfaxMlNWZlQRDnNQRmt10MdBxnr9FcAIV7P2gHej
EMJt1XpxxtPFqEf2mVPU1Ep+l5FPMQkJSTXnXfbs9E6RVdYUHmkNX1Qe6L7hckqh
zYUN89gY2wfl09Aw2r1sTP2nhcsAZ8+wM6yRNT7QzViK4PGY6tCfBi1TKqxZaVsC
KA1LkMZwUNExdZHoadMURHa2yLujXtgze6pzY558SAd+ycb3d3/jMr81RJlCb3sO
mcWKT0Mj7jXi86sjVmRriWADucAYFrSxMAOQH+SZPv1Dz4sgMvpjQOlnnqUnhCF8
k3DJ9JFU1kCs8iqOtHToNtLUioDUiVekqadI1KeWoTOhVnRAZWk9xPR6cf78pZ1S
TZayZV95/7Ikca+/z+FnxPIZcrY7JMxCVTuo1094OyX++EltgdvcnGzzzwdSrDKR
0hca+oj+uy93Can04GyfB/iiqcGaVwoz8feG0EToOqoFa7PF4yC1s4/QnEw/rk/N
sCaJV8PWFzyeXZWEKZ2Tsb+TAMnNYWuqVefQ9f96J50tm6BoHFdeYsADrlw0QsVD
8PpBXbcHUoFK8BGy/IWYXRPx0lOIochO2yuW+0ed5y7H4hQ4f3GhRE/j4fWxj+Y3
0GzIPTHw2jioqpSUe0WoCs1a3fnDay+uW9mIK8+NmEX1gL1nd4nsw2Ol72UFJXc2
gXHcpHP2EygSIfmjcYmcSE0spCCSlEBlM/nH5rixgYDO+/FGJnaqbIOWDWRWNipr
kTtC7gxqtLS7W41t6V0wzNtT19uVm391kBqeeye45hEMvlI9VU/frUXAb4VY9IQ9
5O09gcd2RazVmr1y9Zsfb/SwmeVenI3zHhKonSHeRon0X4ClmjMS6wmxsDzq204i
U521dV6qK46F6yDoFifZxIWJjHEp8fTljZjGw2dJv4z/znNXcElPSqCGPb9Zj/Db
TyGx+WXYae4Hchx1JRAZ2V0ZXQPZeUkw+DmrZ8vz9NcEG76Gk7JOoOfGmKtV1l7E
X6Wrpf31aeLuiGXv5Bjpf6/RY3bA5NCx3Mnr0uE49x7TeEfIv+I/AN6ZdkP2YAc0
IBoEAV/F+MkbBRKikxVtc5jaK8vpuGPAufa6AbmJdl5WF1JI129XbCYLD9jNYnYU
Ar76CYaKJ03+s9qUOo0dKSGtEA3DiRoIYLyJNBNM/is6z46psnDivAcPpyWZgFlG
aKmDWBNg3iHN53ss6tv2kPzVGyZ5sfH5YJvIyB9KEw/e6MU61chGUCIem7IZVUJz
WC7pUxlT7J6P0SN27aW5YoyUltqUaPuvarT3UbjaJhihII8oo9JM5lPkH594hIxt
z/kSbJ6Cp7+GOKYFhF6pZ4hPvyux3n1GbAllVyU5qlP8x5Kd/XKgoFQfMyvzu6YZ
QIdyBshRGzC+9XK4tqGIg4a/Nn4X02vuQbHuOnT0Kx8bjH7b3idz3uLSiA5XL7+l
fUtNaMx4KTUoTl3nbXxA8UutFlJ7leAqe9DvCSSgqSzlb0d/CxT/lIA0ohmyVfCm
fsVARv3ezaPU1qvZBh0rJlIRKH2Fcx4W8g9fX97iAQA4c4GRoMjr+SLHEy5cqgV7
vRVvab93ZRfmFCllHg8LTVjn4GWf+K/dm7UZKE+anYw0C4MoLS1YuXLqTTQWXa56
4iITHWQqsbyzX+uAGiLeJaPsvUQq/hNovYm9FxB15ibMMG+9Ne50FsYdp4PgipwO
O11kNLTh+W28IVQohAYYHf/J/h5a01H4hUY5Mfp4SQtUsQuDFmD7YjDntq+D0FuI
8bCV+4xboKxPOkAMR32K+l8VD16w0x4BRXyRIOia8KoHOkMBltYEOv1AqrZxD9F4
B7RkAcnXLk5hxA7zJzbJA5oQzD+8tUoX7oqung9L7YKAihQxxPdipSIMLZIjb8vW
ocQyyVYIiZo5jXEpxCYc6eI5I2VjgGeABgZwFbXOXnhfDoBgM0+SsvQKi6GT4Uc1
NkFsVetEE4q+xKq5626mmIsiU0pvXiWalUR1Xm2zGlzn/3B0UMfkYNJ6KV+6SJVN
CSbo1AJNqAn5dMhcBrXgveNyc71myalZjinODf1jNvUcQ5HVyT1/FNewlj3XtyPB
+OEpHrxVPut75nHxLcBl0bE1OdqQ6UI0zUTjFTpmsR0fBVwL/uuA5m8IuPR73OtT
Fqq5mhkzO54DCoqCYG4/TmAV4t/3O1ckfGt9gdlUlneldsj41IEY9VxH7h9rqEss
AFvXF/DEACSQROPlTBk2aDlMgxjOo3H9cpaf3JzoemW7mU7r+pUkiCxiMavqWQbm
2VqhJvMIwaYpRWDqFKR0hr/l8yMzeVGbBXAY02dCoPyok89BEUdmVFh1ksJDH2Pn
GxO/2cXbpgEVIcs1ea+YgF7RFIiMFLY/+GM3HpZr5SvxSSi1MsHnfN1lkVttMLnS
NdmRZ6WkEqTClXnyJ2CqcUiEkcsISoiUw5oLxn6BubDbuC1Ea+CudR0eihVAWAcX
1BSKDOWfgGn98uxTJLYPpee90j7YFNOV5tyVTupO5wibapsRf8LBOcknPA0vEZRl
K75qgGccNHxNQkZgtx8tVDDv6tVFWOie+OWB2vz9HBud2Yzwo+ZFFpxXNpc6KcQs
7mvLKKzhJkO/+k5NL4+GUcs9Gy8OEoW4ZQpxfBUB7Hqe8TA3w2y1ml3jUcJhvF1d
6y0hTkPvW5Ej151QH8WTanbrisPAjrdA5VNw1aBQ1fS6FtqURemdzX4ZK3v8w0/L
0R441LSkHGVqn0OPnxhkYQLhe5GLomjTWW6ED7Xhjuwrz/lV/z/GTSWrRilv+sH9
IcnQfPUWinNW1JpVeeGIel2BzMxW2ypOqdM9NJx7gOSfmPgKHNNa7PrrazcWihgz
Hj0tmdDoYverJ7lHLLrIOD8k4XgFSAI4pYcdcl7Pz4gMAZS6UWxwuQL9d9C2+iEY
AbHWQSpH8hK5BGrrJIOdJuyOjB16I3NyfIRNW1XBAnhQgQ/O5qcSAUefxKlun79F
kPvg43KfdLXbYpfv3/XrDb1SDyHBcPghabhRoemLnn6MyY604Nc/Nwc8/aZWGOuy
qSaDMiKqetyHhr3Mt23d2OVJzrh/8pqdZ8G04VKFCH1+cXiSYvfirvvP6Z4/Jhmh
3BtBW+yxQJT4aYiWrX4fyh/X4RjmlKKGp45kqNc13hNoDC8o7GNLYy68n3MuN5U6
s3Nr6+kPUVJBE4YjHZ5omhTtcyhrsPoEdcKwIOgfrSxIfgJ1/2GmJyxGVtCH2f/C
Gqy5hG6YfhQNW4Xsh1nycm7BEcwWgJoLw6y1GUtO/AZjLNJSDL+B3boP0gjy+Q89
g8HkoG9Eaj4OnmPWXBWtas6oQhJSBH86jiXEkOcuckLTHojPMhLl8xexlVw7D1rT
I2MRIdPJ3oLVHH5sdeJsV/PPMo+rGipqWwg78WPx0OM2TWjfiPGN60we6Yaj8nou
3Y43nNhElFufbIhUxpaW1j2/9CdiQERpO+WWZu34sE8rtUmcr+8EnFczHJoKeWZ9
FZFw2NV9/qIiTrBdeYkcONOiWQdMxZ3MGkvfaIx8YDe4p6a3XY3SpLukCUUVHBaT
wfFHv7HZPpdA0JQ6woNBH+zXqDSbAEMBvQXkqxk/+RLszlT3U77K5hvG+dADVcQV
VWAFUnD3KBoOD3ehceV/lK6GXSNhqoSWU/XZqBE9+Z4g76XELzARIgkA74MODruD
vd34PF4fm6ugWsvIhV/UxomiVL458CHaRBpg/6sW5/iNPdCX4Z85N8Xqv91/T8A1
399SOWzimX9ETI9maOw0j4YfW0d2Rn1uQqJblrPNWkIFOKApuz1Cg42FbeNgbXxT
hCIEhGJW4166CmEJlFuSa3MQjCO1YRDcc/1DHCEHDd+4t2HI/mcMHGHVDV35ECVn
xU18mfPjGHPxhtJaGV7VMCkpkL4wghwv/lR9b33ECPYaIETQRHf5uW0NEMoaLANZ
vmp/JVPraDA/QcTPn0IVDkzJvWSeRYlAXntbvBuv5Y6uecuEaEuxCmfdmjeBIvR+
cng8l+aV6I3wlmmdLTB4HD6GRhiS8exT93Aj8GTTTXShU0ucxfBZGVEDN6cs9Gru
vm1Uw1qVprtWjYuTtXXzhHB1zTlrAqgZnFnUxsuKxgpzIc97OsT87ATeZ2lcseY+
vuehKvG5ip9jAK0jQClrUnRzfwoRYEMjafoxmV/l5gnY3X5srLd/9qJoKW16A5G8
BTwR8yhfVA7BrVg2gC6hOi8BwLnZ+p17W1rgopPO1ZerFsLcVUP9dZPdCDCqAggK
5N9lgY8chWLlmO+6YUEccXp6H2JmSSLZ8XivOCm7XpcMBQ54IQxlv2lrUs1gWZSh
r677z0YxwRX9F9lF+Ao93C4ey/ur1unWs0k+J7W2lqLLXdx8HuuhnkXg6SAfML4N
usI+PVvdMVtmywPWsvCtQQ5sTwjq2DmERQm6FVGEeVZxlEwq9JH8TT322m9YC9qJ
xlwA10Ha7YPsB5GHiV1zvuW+rTFTBO5sVUsuM11WJR9bFDDmWPd8cmnLIWlMbyTN
QrdHLhrYMfyEHR5jBT5uLRGhkNmyGTMFq6S6aPyOURBmUgYd9qBj6T/JFjTXLime
P7OWfXueUqCyPBrkXJHJroBAEoVo6lEMcVhTUEtaP/O32xm0AnpkPyx/uS2Rbayw
ZQd93NOSQxT6HOGtAMMDc2cAnN255Bqn0gVDnQMghxPoZxhzfQ6ixQSk8/7B8bM8
gtgk7B3J0UBZvbt0vgNeIShqMpqczkhzWsq+D9Ty9YCWVbgNjbaUMbF6BZLXgxfe
PZ90jdgH39YFS8W7LyLcNe8KKQazwiw7K2ReQxG+091UWTMFcx4auW+DsGab1jQN
bM3dXZEtYiBiNobek9LHegD5SB2/T6+bfBLxBGJMhdy8ddEzGnHeG4BdTmROXq/e
mEdHHIgGiwEwly/7TIl8YlJWWtTERQWHF0/p5oIlPzbclhqfti7k9v7DJir3KtvQ
AN1EGRpequzH6pVojQDwgbeHR8JvnaKWM2wt5dLNm/EUEGGyBBVl7CAT0AAwtDdO
l/EZFU5AJLLqjGB120737e6p1Mjz3Cl055Ll8Is4aQil8FafI0Y64CzHq5p0XeND
E7qIVInuPpElklUuABnL0Xp/ryWJv9SbM6komPH8tWN/zDPBaXEScA5Wl8zbXpBS
NNRbVq2unOT0XXxGTdC4LwI/cJRCkdZz859+O84IebYDdcPUxn52gPg66cxu+BOn
rtSAs+9CqIy00CHJaU1VBSxg6cpljE1od0OLFnzEZ1Srx77Zi/QGb4il9dIhpUTc
Y78YNYQmPvKLdGMhYcrLxFJjf5Qe9C8jFCuuMLMj05coJpqvp6S2ULZD0vcBKTiX
dEuqFBWFnvKcfxkfyUbxhQo7pLm3YZqVguX5fnzktsYlhi4beCWGXRQg8NnJGLDy
Rb+7eqsfEUe1zeYwtJgM8lFFjWQjGpd1xcMF09aKkMA=
`protect end_protected