`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10080 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x76DGZo6eK2Dnr4hTEHAsoG
XBC+M+zTmMWEHYnyqWAYQQFwGQ21V8Ric30KMH/cMBvrvVwmNn6MChbyp7UzzT5z
bZuTFTkMwxdpYf1DT9Uz6IXFv44PTgK4I76+Qq78iXffS1BOI8hajb3aStH9LVJI
sioPL1Lh9/mt8kZfEbopCQLsr3Qk9TfOsu5AtI+0ki1X9NAbPqwEXdE1u5U1JXE6
XDUhTP3/xcUXC0/QexMXRHMwldP8UxhL6LFZxlXfMso6coWdxe3K9QrE43LMsXD8
zfqyCNkznL1uYGOke1ZAdO17pDA9tMNV1rPJiK4hwGQlhBPZEZlLTWRVJMFh+PDK
a1KYSDJk58x2TRC7OGpxP9dAMBXdknsmMVXoBocI2ZbQJOQ+DphSruCBs9Z5WnfC
x3gb61jQ7Wp4ynknblPbgdktaTwRAuHi19LyDr56HNBnQxJZl51uvKzJp67G1KDM
AYAuplUBlwRQAsFMzWLEVfDLscO6q6tW2kUZWCONOTUd121WYwnjxmbcWPz/6GvT
o0LB/qP05A5kCgzPWbbk01TpeQF2vY3DVAgPhrIr6iGi9cczrfXSu5V/4p1FI/40
D5/uzZDkUMcAY+QsDhJxiXxJ41CS8PI7reMCDYg0dZL9t/35VSN1pBmD+DZuOlc1
0WwqN6sFYwD7Eeo0wOoFyzcgi0gbhLa5nMkfI4NwHyhKp6+jhZUaz6wYTeLgeoJ6
McRYJoKZ+J04/AtAP68L1/eCzBQf0FlF9OuA3srcFaFHJrNGWAdWpY7xS+RKuifV
1e0ka0cFUglWh1vQkMFeI11H8Q+rPR4vn/BRL7BoXoCWtSZEy3EVvhUW4nkZFd5H
SVsozFIOVwuGTmOAst6eP01W6W+DMWxRLRETi8zfn6vRxAH/eNDXsMMMOszCa+vd
sZEWopZNV1cLSeg/732lhGf0+bhTe9AeiG/MXCWo8Wtb0KhHkgVR51ZGNgmkr4L/
EaLAhao05H/vf7sM0opYxoI9DXs0mEmhd4J6wwtgFdjxbgiyfRmhtAYdRiq8NnwB
510FdtLRL3I06WCkKMQ3QgDcOMiVhNuIYlMV4Jb5ggLh83lYoCeWm8ZScaZS/I8M
HOg2wa8WUz8sxn+79SGEJc6LDcMV6mPdclUZG/a+8sr79nWOvzhjn2/HHhb1Pn0b
++xLJrQgzEiZ3oxEkFc/g/L6kYLIfZQ0lHqe8E+jy+vknmfVmbxaEFJlKNfeuj0y
W75uhiY3FXUxc3KUVD/oBQDZA9tKMTg7DB7wnNAKcIlaxBPV1Fx4v1oF+6YYXN0X
VkMJh1EyCO+y1FDKbCJqV37nMAUwcELniLWF7yvS5IZDR72qihP9PHVCz8NAx7Ig
SDUPFwP6ab/627Y+OiZHdww8CdbTE6mrAlUD4l38PLVEpNIoqcQQPiZu1Z+yRDDd
qtORUfqkOn2KeawhjwYXlnQ7iau7llUUTJmFyncPE1vHfW1lOi3xkJH3WRBdkoiS
GDwNvFgFT6WDn+T6DIj+Yg8CpVHOyCeIfrWeBDSQ3nXAvb3/9/Ihqy51J7fhX+pP
w0U9HhaMunDXRWl9P4/TPUe62hUMDzwxOjkDQf/tYr1uwBzwhc3TD/7V3msyI04A
E1wnaYyn4xSI0/fG3E42Exczh2qU3r6/pn8PTO25dsryXBzZGrGju7NYgYKwgOEK
zak/MHPxlUZ4QacoDefE0xIZhGD8htF1pbVrZmNR3w0VJt1dhLpZEhLjeR+p7Clu
ga5lHi6wXHf+hBlcDEmOfVwwe8/CK1NIp8O8vCZLy38E4Urdm43bguTkZN2fC6iR
bsl+F4cuQJJbKLcC44I8lL2118g6Ivgn4Y4gtd/qXmqTizPL60zgXXY5wP2WVJyd
pSk1+ynF1O8Kf+mYptB9vUu4qSShg2Kw71ilXR0POoYgJ5QOCkb9e9wMY/2WtP0n
CQE4U8MaP56ltEQ+na+UJfNRaSPvLoV3nMHblvF72BlMwBF06qeJH6oJa4LhXmop
P80ojz8UDV0sXO0RjuCZxESK3ftuYnkGMJePFmNxqsLC3+0kkUSxyvBASNY8DW+v
OV4TtBinjkQ5vfIGv9AFWmre2QnOq62eBt1LR53xgwJnmaUEr26zRolr86lM8VDa
p7LmihifD8WKo2O9l1fdshZkMA7lgAEIrSl8ql8Hbn+/BI8E3HgeJ5l6mP4rqwV3
JkU74YC9aBU2eR2xrwRl9DuozZLcVcPdkq2+i6Y2p2GoAKPA08fwfm2uK7WAc6Hc
LTj/jFF9J+m/W9qrJmUuKaW7JNkTy08JUGDvR9lmB0EgAFlmOO/V9hwx9vRhMstG
knhpIEyAHI0hhHk+wcoF5hWoDsSuPh7O2B/4tj2tbceWJ2ES/imgD0NDznIQnUKU
kNmeqam34+z1jHiQIAzhEorA67fONItuGeqqiTO0j3aXYHQXn6IzhkP/Fn3w5ODP
5BfVYASSlpyROH4BaYPknZIXiCIUIonfd0lM6YXrsErmfseRtqnLyKm98zyD9gs+
+rMXeAnM7WwwDwvah79bPNYR5AmWSTq6f8d1teRQpUFCJpRuziFP20SBiCyJrjcN
jEzXRBldNDUQuWwb1EAvhkYpZTXuSEd9vBSUiaP0HKyjl6uXl1aBurp8RFyIJyIV
wX0NZLCG5kwngRH0PRbhBPw+xdqaQDKMITc/+2HyjLi8nMLC0yC3N1ZmScIgBCEM
RpDcTXeWnccuCa17o3XO9IKbEI8t5Wz4UpxPngxhWLs+v1+cAjWB3GNB7FEwB7kA
bGuneV27d9cKKFkOXjByCjpxKMyWCB4HimivsnYDzi0K+IB0sC4ilusjr4af2ooi
34IU90ttkhIPAe6h8Pj4Iy0DVcAWr3Wy/ioCxLu+P1K/02/hQHpvLlaeF4o8gMi4
FXRs3NhOltKxrfhUon9WgG39IDMjPMTNTTi/jQl4VC9y+u/Txn+13HgvMCvnPwc+
mcPUZn8tq+XmDVjMzFCQA74t8i6Vt6FyHsQL3BeKaBOcnyYsKIKhiTIGNu8n5x4c
EFALbjaiwMYfFwpPPGfi98ou9w0rrH0i3e1N8rFlb93NHOEmFuu9N5PE1ajoV8SR
yOs8wVqZyEGOICGSUEfvHFSK+buqUgCxJvLvNwPvRrMSGCfg0Jr0rUeaSnUuZxXy
Kn5/3QQB+wYMJrtk9/lQIr5M6rIpmSXXmHLxvqNgY8pst95WVcU5bWjlrgcejoPa
XBqlgMpV+H5SWbtHi0hu5Un9W95Z+gUyAyPtS9sXQ1PP3U46KxGQrlKjXPdetpTW
oQVX09jw81mhN4TFRyV6LnLD9afZtzZAwvIbRMY5RN8yhxqwbhdDncCjXAzwyjwB
QKp478y6cFXkyvoOGdf2O+9uD+jebPX4LHCguxkgQDBhpCOFCbPEAvpFBl7xCIKp
8Vi2dXn+77vr5uKtWemkqCX1C3/AghYQw5SKeT0fFVpzcJ928W+xr/BBOTPix9Tq
Qrn/yM6FWGMBa6eaNZW8zCfvFum+k7JcS/YFo4Ouldkfp+VVELrY0nF3dZc09epe
EM8VYTfehm/1dR3KC4vNjX6amJRIhZ/g96ON90o2GqQVeawum+W+49x1OAl+0AMy
P8MW+XVIoPULQuTqgtoOpwjBVPldyVYUmw3fZlJaG5x+L3OE+S0wvpm210WAD9gZ
IRUbJhCTCcj9zkG6P/oUJqznQXN5943ee/CtszoRQfzTnEl/rHTuDNOeJ+ZeHUfS
l8wcpTpTa0+cSDhflHDnKs6laq0LiyG2mybfko6YL2WDco12ztcKFtGgcD53B/61
ZKcxgMT/rt6T9BJjnit+9e86ortsgcue3H3VBfONO+mGCoPBA8TN87Yyu3KTyAhD
7pokoD5K7YhhgV13VjI/8NWfdr8g3G//oirvTnpD6eN4+7IGuet4LHyNr7ImSDa4
nhcGEwwLByLO6s+g9giLzDyPg19Ax6K8fsPPWFxHxFk4f86KU9Jtu/8MTIPZjnm3
ffaDW4GBgQDu1jqm+E1L0ccOCBig04HWy2tHfLTmkM8rU4brSliylMQ6fBp6qKGn
ve8ULDjjdjJ6CoAhd87Ht84Hpz/SrnCFpyt0TyGToYoADpxJfFXfyhGIpwSunrik
4+rt1u/QP3J5sqjgtw9L14KU2qbeRwb12J2F2uvuljElzyonnvM+G6kJ84GPI2DP
JepiKNJBeWpu4Glb0SRyffMuZKn1iervJ/8s4NQPzQnzDC4n8bBfKMNBnZAmJlaf
mAtgs6p4ckkMqzHvh15heWgQyc7qC3qp/gJxGv6LdZSlA1H5/LSjKxIThOpuPBg2
DXf48IVSx8l2m5cTH9TdpaAe1Qks7OIVLjYbb6Z9dStZcYywTh8Q+yo4S6LjgQ0x
44BPZhj1fhbU+5D1IrPAih1+tBbHS4qQ36VadVOR4SXj4Px7pu1PkeamBR7R2d0/
XP8ZrNWEpdvNyrva7P29sg6bGNj2clTFgX7yuR7kxboC7wHoHctumYiSJT/58kl6
jCF+oIGUQodnnA1Dq/UwpLt09yvgNZwqXzlhn+3vBAc7l746EiaWYjB0U8PR2h4q
GsvV7eu459FWRs/QQP6BhkkUXLJ8acn9ORABGbQjc1ER4GZhr3ViquIveSINtx6W
VqpJS72+Oy1DPHbCHcDhOhaDEJ35oT0d17f6CbvYOWxalO5KudzBYSwxOOh+DdHe
r01/CcQe0KROvzAMlZV3y9adOclror1+/bP3766xHYiLCwRPHRLxJQKMxwQM77K9
Yz/QStHqL5mMh7tuTl9659CKCO7BViRoRVPapyhkLoNi94ITx39p7zzMD92GN8Gr
ZRtGkSzsmTxBJMCXwIjA6neNQwJj0M0Shq/7L8N8xcJgHEfynCbr/A57UZ0jEets
8txj6VEXnYmCjol6VjqNw7SWKEnHr8pyQ4Vc1J21HawhsDBPqgIBkh1k8q8uOhDv
YcXQwmRxOO8q4fCGV+QumgtVpCoDNhZ6gOv+5VHIrCyGCp7aGyld0fty9x0z8e+2
sLSgOoUfnpFBlsrsY6AGl9gjJPvvlEyIkvElrqFq74dp9gmUHjwEFyThQMGTZeAa
Y1PUH334yaEkdY4+rjwG/tbHg2vdGJ+Ng6xI6cv85s1Y30kvbr26MwgznDvQUj6x
PA2u1gf5Apvz1mAH+DhInPgNgnHn9F7xPJPE0k+OqB/O0l6rVfnQfGzAhCL6vFDP
gB1FSnVe2637dWxzHggzhXL6jGpDG4HZF+77fFPQNSuakQW0oXyNKWXvryfbrM08
7LY3AWhJwqlEk8VB6d4bdsNHYr9/7dx5SrZbMUXb6hjzbnA/MZUaTsyuH3RMLLSh
MsQ134EA0yEnCK07Ei8xAitOSg50AC8VFXJlu2WEj/gyYBXypuDkqln8NdlB6Dey
8M1PPhDXRojZGvwa2Jg9uwbLV++wGiT2WrKfY1AkIg7Ft1qfIezg6ZSW3hj4dPtG
if9Xl8mWSKu42trOxDYrG4JOIz80/JdSxOdfSr0tFq0lMJe7MGl7yzJ1HgfkNuXN
CaPbpq5pcmGeUp73SGrtk8QFK53A3T+fr1oEg8cdrm/UGtpdSosCZVjqW/7Vj3Oz
rdTC8lUReUfuDlGnfYVWvItg15EMsMgh6UqCkIwXzBfRk8HOH0Bz7rhxIYBf19TM
Qts6UKfHWQ3ZPUFe4U90OFtqC9j2wX3h8G+gYOP7XkGS8myTShjRKuLG7H2kEQjY
djFCBRHX9L95XU0/OCX0IWRw3QBIAQPFY1mgT2ovHC6Aj7zCTCSDUgvmJ0cb3hBI
+hVw2C7QUXxEcWeTAEca0VCVbHKw4hncWnGuNt4kotbB3+L4vedI1pqGKdi5OEhY
9F3xCkRLkhzn8wnWw6EqIWqTosUMQgqojbRTFv6y0MUJKwaM8HD927zzl3Fh1gUR
hFP8F3kVNrANRfRkg0kQrnujEuGSeqSPufRAr90ogrcHWU4QzvMQJhWXzfUWtTpu
t7STufE/s+7m8Hq14Q3LR8JTEYkGsOPTskwAZsg+N3+bW2U43tSHd8hFMFtk5o6p
Y6Degl/Wf3aBqoLhK9aMnLB4KyqSsRz8J2tce8/M416As6AYdGYGcBxpaROj5UKz
mqA1tN5Bi86jn4It+Ve4lQEiJbrOOAqiXOrE7BsdIUXCeM1prT811cqN8WzMaJSa
IOCoddrTEc+czVEvYTh6EcitTnUbGO0cfn+JleAPpkEa980DqGChOOV9IT54XL95
AUxYv9NMGOBRLStauqtNjuoNQdmygfOJT83SZFGBPW7v2oKnFFXSnqFX3Rl0wf/L
YK2tvgh8W2yIfOK5nSEp1fkBy6BFs1Yv3bj3phonOiZtNn8Q+OYAxpE84k2aBSvw
ZT0IbqV60dYjyGR+PGSmim3OQjMT/u39BCqHM+UCbqFumZoTN7j+U54PEu4pf/2P
EkwvE9AFp5aMvGHPwgzztZHim6E6/ajkKxZcebbRASB+IPM4bc/r7/xOf2jQzjyP
hm88++SF72R6tMTHIZdhJ2KLSQ276COcnCBIqnNOCUNHa9GtBVN8c4ASn9bXAhNG
Ixy4A7VJ4EYXztHrR/GdJLcitXpPCnXobctuPK0cj+J3mFTjGRM7xx2NNma7Wwvi
bKASTGb1HB2ziPFki8PWZMn0JnD3G+ifWYemMahA3Ifb7uC2qBK5TQ2WiUYLOuXd
Pc5p+jca95sBcZPBM31IPeGGKeYLls8uJoa/VHfcUsOR778ak1CvQ68AAYiBMYbD
KgjrXg9FYGPY86PzyJBNwKJR00veYujvAhl9x52tzEN15fDVjHtfki2t3/M5Igid
69A9JeDdJEvdmdc62I09IKTSm2FrBEIaIIdsfS7/7QNRzQ3UlxFFXJNTL862g029
IIrm/H1BAJjW6/NC28HmbHOozWyJf2vOljXGUuZcC5hjcULyqxcdkFSIpubWKQYF
5mr8e8L2L/5Q+dOXOHEHtOpJIucdgR8iJ2EiY8jSfFxbMwaW4Zrn/JrTFpgffMqO
vfTPGcxYcy6VXZXPfKVTVFBEMebrJ1IapBHHzKd2j0wGPZJjA0QdcaDl/z+bxzKr
SQzpYPf8lfqw4PuuziJ00oRho22MAr5NzM8+BpTt+fFIorwHp53n8/fhl+Yyq5Kw
tP1ic3x830m3oW/Hsmr2t5kEAvnecZ9jw7nqquj/LbbBrgqf7Y7wQptvRu1lmDpp
aVQ/qZwo3iq8wXZId/4bSnsYofmlrjtoIcbZs7IrLZtjxnXDtv3JPSh5+B/yCY2f
58ZYLwimZTHvNE/dXxAYFhZ5dSRuVkToW1s/8VqajEWmuyXZWL2kfriKi18gak7a
dvbqy5R4bbJa4alEvpOTllhVRAsuZ+RddiMAY8Ns9T3E36gW5LiQbAMwYuCIkYPR
KX78fz0+1MHIWOC0bzcWweN9k61l+hlva31H6b6iI6A/XokAy9IaZeflqJQwyyvk
elsIqwOdiQh3bV/Ih1bPCKDZ2KOUz+5asSqzzSc9IwY/vjB+WUCaAh+/UmZeo1rO
XIi/1SHprmdZ2eY6g+IgCkh0cLvA88Ri7/iGO197Fmnu+tnaASXH7I4JvoZTc/e8
VES943aFF9JNkUGHmwRtCb6iNiwOEudJctUONC7J24ZNtrza5j774mXG8lxoXA05
Qduq6AD9OAcMUWTL4Wu9bagmDkeeqDC76+mwWBYDStq35Li785osO2Luyj6dEGUI
XkaWT53KT76/FwA7Pd2FBTs8rflm2Al+J7xbLVPRssKpxED5qlKFuaheVknvOqXd
78N0e+am0AFmj58mycIhtAYaDmaAc0LQ4srPrhtOBrxoiOeGDBBQOv9/UvYT8Ilh
ZEZUiOOJzQYiSxzIwv/bXJGwSOzfKieoi6UKecrjn9bH5LNRLtTdgHxahZcEk2Iz
agqUdKyOgyDZteQ7Y0zeegADakYuSNqLTT1mMuUuryK+Wmi86IUBkfjDHAPfsQBq
oGw+Hn8iGu3C1AInBXkFYcF+rAVpoHTckIAtQdiU26H/m/TYmq9/9Id/JrKTCANq
DSZLpS1245mVRG1Esujinf/gD0R5XzP2gWRb8dQwSau1dxu9n7ZemMtgLaT4O8fs
RxNCkHtFEx0TFHZRfBj8O4GYTbQugnF5UiW9iFDmtcPdQ0pGv8SnXE2WEiOOUj4G
4SP4Jx+DJAPyCiGKpvgh4QwIPFI2JF9o/u6cDompBIb0qGJMhsVew6zFnWj6lIBL
xT/ApSmBJYllLoN7lG7eXxXq9pjJ8lpDmqsWqGvPpXtKG9IjI//OD/IjdtjukjXY
UqtoxfyV6AdO05kd+jAObBhny5nmEz6oMboXLKQIYUj5z9b3dSUmWKvcedDBHrJz
181j8+QN0320b0lu13G5kwx1Sn4VWlZnfim/u0sUfwObSJT37DI9gSUucYhL/64a
9IZN2dVpt+SBcaGNlrUHw2oio5atlE3aaWZMuFE+m/mVrL1ryEnVjgnjywuYSHVr
r+erFYmGUbm5PQ3ylilTZgnlidJuEz1bhWUYjNp5Bnz/4mc2vT17gpYNzlGyrEce
vJjncdW5d8LrgwTwk4cfiHfPeKFhcVlVnTQogA1Z5YUkZKFd2vLJfxLSdU/7F5t1
Y4fJNv5nAN3ChavRf+2f1T+mNWZMUI6eVe7D1HIwJSy7GvAK/iqYMV+RxAxaHew1
Nc+AaeTglLBz21q4AO7uNTuErdhh7iBRwEn/te0Rplt+ffNKKuEXt5kCCjygJ9dj
IKL+gkwwnU1tYt5vYAdFs+0v2Zyem4XU0Yfe7HZC/GBYBgRXBzZvLWh1BbAxAhbT
0SHaD83Lj/KUbSHUOEGG7Ib+C9IoIT45Q37fpi89CLwL9TpnfK2bjQvpw/Z8ZfLA
YmWwBkvPGWU6klcKZ/s7m+UiHin15pdCyAdzZfGZP6TdyTFEvB+YZbiBWp88nmNT
33KNkF7HRQu/H6804+Uqn8VVCT5ntLqJ899hQEiey9mksP9hTZp8vUXiux22g/tA
xfdSKtkQZ80oYjsmpJQw03SIBAD1O5VXEFs0SLDmyAKhdOGdlsONdCYYOKDYQFvC
Ujt9XfX44EXu5W1Gf9+5yD5W2NRCUyeDGbyayYfRIvAQ/bodFbNxc9MUCYIcg1qg
tM71lnbnZvJOvnglJsjMTyu+MjO1+qnPpsErehPoG3F2uZGTfmOLCL+TcJNWGsuA
JXzJooygLfuLvIW+MYfw7unEl99gKotArr8K8ql2szg6ZEeWFR9mtXNmn/wAoI5Q
Yi+M4qYMXht1xnAT+KBEZngHRnIJdqZ6QSDjjiSFNnZwxb4n108fDSJFa8U30Pzz
bdulz2WZSajuwwSLjsvbNYOE47any0fbQMlH5+xOp790rttY5tKpFtHacabiudFM
+XgRFY45aHmuAhGcSAoT4R09xnCaAy5zsW9n5W6M+OrpyFvhZGQdMMIkIY1xmsbQ
F2vQPwriIADsiNmV8u3Q8MgDZP7vgXI9uRgiEpjXtuQwTxZD8TNIvPBZsUkg5UR2
0udo2IApXAr/SaUqIAt/BEb261aN9ZkQddQVGVxwEMadZhyYS5vVWHy4Ox4WmakA
eh8Nhxy+9toN3NVXWEqTA52E14UTlyk+hTRxS+a9YwJENsueRbm1hrL+nv0HA2sT
zmAPX+IZeU9u2qrdq7CrHmVyS0F8J7946AvlmmBJREgKTp78kho+5CKpT7ym5pKS
C7CpiLYOVfaLBUnIWaG+nYEZTSdwP5nHa+GobOYt9vrkvDiQbGnYqyxLiNAmRr9u
iewddfYlelKAxzLK9r0liIP2YOncN0BrYRu4WscdAbwX9VtSwMMfCXIpzkw1ZE0O
trU63SxadJCK2mptazlFXDM6g2ODP3u+ZW9gBeFRsguD0orIQdWKKjrkXtAgVv9+
baRqFiyd4qJFjTjWyF+WIUqbThD5dWtLWb4vavYL/FxVuqYuTNzJZoJzssFoITJQ
lWhOJxsyD2kNBUB0IVFCKRds5KgqC1uSoFbiqXoP+kazqU6Nsk43+F2WzUkc1boe
2gTFgAkP6nUzlCUrKFWu1Fej1W2CJ64xV8TDNh2qr6CM3UkqUAjd/w+B4FHP+Wec
KWw+uSioKBtPJJ0248xov+PdDw+VwTbk0raaae4jfO5BTio/IyOFHzwg88YByEO5
IeyZas4mq27eyqt0TYSakSJD9Oe/Ny6j675tK2DcpoJOZJq1Dpclwh/4TPvcgpW4
E0Lc6Izf6Pi2zZLBudMWPL5LRQEjatxB22DHnzwnNibuAvnHBPZvemdtmYCilkiA
zwOaQxu7P9L7GNvQC5/2Ksii3SVmrHuaqMSulHfS/+OUL0RYhA0ZAM7hooSlf6q8
M4BoHe8II0u37moNJRIzWQV+qpRNntkPEYrN01N9gAuFUxD88Mw1z9+RDN9tb30z
IbkxDGkzAz3OMcC+ItSV4nShvZ9Jwp6MRsONdHBdqRH3UsyxYeV1czuDf5z3sKvk
qJGeuJGUrVW+hjR3dxxv+ZiXqkIAqQ2an49+PLeMEz8nSBCdLvk6cU9GC7vsdIQj
hyV5FNwaG512ZXQZ0vv4Ku3mOdJwRipVhtDQJw+k2ucFbQbBdmpdJW/837q1h6ej
Di6sMqoJ33GCbrFHqLeCDsaNrpWf5Ua0lKA6UeM5thSMBTpykTSXgXVUf+M6eK87
KuEK3SKblP1Le6D60rViw9YO0VAd/nsBH4VtRxstODZP8dCBYiLY0GBIcpuMf6v4
CPwFXFqHboErHfFRlX/zzNwPPbJFFR2df+su11AqF83cX70K6ww6QceQAe4DTOJN
aJuBt9400at4YmWf+2fEesNJBxF0GzHL0kvi0+NP1bqP7PTXH/Zieq8b20ZHKbmL
xyL8l0hgjGlF7/L9cPEavUtx8glVqQ/wLzspz0SJsb2crOSo/Uk0zA4gODintB8w
MopZtMIUu29Ys1Ndz3j53z+DVCe7ftMMrjVUC/5W8nFamXtJnhD9fXmSld0eQgx5
PKEU9xbUKd/AvAb1+JfkOs+R59CArv3m/xLddpyC4e0V38aDjBQr7VL+S+JM9M01
nCGp/eK3G7tk8rND/XpmrfI4r8evHmPDCPd6kI2G2cj/awkIN/W7qs8O68krpAPs
/jXLLQLEI6F34Yhy/JwlFI43dsxQLlDYQe5zKtV22ltf716VDQhAlrw8r8Q9Bgan
ohLnysRKnIXLEZ9h8REBfDtQOLsTiBbdLxGA/ETS3ALveAyxdxc+TC1F4d+oILQn
XajsKLVTt0DRbHpROw2ZHECKGAdLGf93Lqt3Bc2gy9d14yrl1tIsi4GZgyqV4CKP
+eT31f5zxdT0Q8xxSLWKL6+DTgN1MjBI1kSX4FR/e7oZxxCKY2YonVJ8Pjm/WP8y
UumgKUrGqoAppEM94KpZvCQla3+GmoM1/cGwBIsdIsg1Ho5DN/tFdzpQo5jO0FMQ
KDc5TXXxmquaCbWwKM5iWV5sZtoTDtyzehCdNNTSaxGULyF5tFF7FNfMG3DdYENL
kvgT/lmSUM500y54If0PU1Tf3YuCNjpkJQCM8kYzR8oJ+FF698GGuhmFQ2rzQYrl
reSQicBE7z0kY7e8cgoXm4nF9DA1f3sTk8SPElzLVHDj+Zm3mxe/oIUx6kcy25Bq
BYS2898biP95rXOhW/5vJmYc4A909TikFdQfzVIZiHzS4EE3oHEOu8xi/bkh7959
oAC2FUhJloIlW2OGPFSu1oWjLSPwfpm0HBFWMt9JqNIHJ+9ObXcmRwYrvJXVbf60
2kmpYt32oXJ6SNDKUrQVcspXHilMdqxKdzzaBYjJybNyDI2gk1xkPA5B5ycbqZCq
tXYEc/1uRxbqzQWzueGL8k2pAONxPt39MB8GexalRubw94e7F4xqFbQtIUlHcfh+
F3AodiUSPKrQcAaVUsUiH9crQWHdT4D1hFKgYIHv0hv62kocweepkc2PehEEIOs8
JviSJRahhBKiDfB7QJY1rK1czHsmDdxXixHlcX/E4xOrOqRck6FaqdidaJ1p54Wt
Wa8xTFh08o+Q5CfEMnl2bKwsrqGz9dn78vUEftQ6QFuADTiOYZvh01HJ9gcgfNxE
K4NqSIlxo7JMN1VMxmJEQnH72Q5/zt1JvjhXTz+2rVEcwJkyGB0JUD09oQrWgtL4
pantHJDNRS3jpDCD9TmDs++yJ04lveuSmwHFAsgfSevnIkSmL7tmMCCPafrYyyJ7
TzFESbeMD5wIhLo97GLl25rtEQpf4UOTIffwmTF5Lsv+LfDSNXB0IuRWrve77Vvj
Y32H633Xi2LZW4tidBzORysfFAHf/jIkQRLGdtylxowVJ9uGv40W4KEcfgpTQ//g
Ie4BnzZeP1iXVGtfielb2TlQ/MhM3PJg+p9mUD6kaeaScnGaPCMhEpJtmDLIypWR
l580AnJoplcVNsyFbJ3F5+F0cUTkj6swCfvL8KL1hj8amRwDrp1HEKuGISHQ/OMv
p6g0fkSb/Ehf9ObDC4J99FeOvIpHihshL+U+sBHMi7FQO9PVKcUkcKxojBPFCusN
0EPU56fq48ao07bwVxUEHRNbguJCpnTdujx5JsaA3XCZnHrNvkBATbk53qPfAO5j
FadrEZ3VemXlBFzMux/I3ZXb3GL5PIgusqn0Vyz5+ZHdek37zrcHCqcCTF+/ZnGx
6ww4ZR090Pu2SCtgcslYJLFDN9sqaTZMp11zOi3v3MKmyBj3sbGAQqCOW5OYkc33
HJcfqyw0qVqEa92CXKhFmydAUbkseFka+b6LyL2j9ECPKR71w9+kDQjJcIlHdczf
hAzGhNyc1VP7mensw+lE2sto+827KPQk+kCpwzs0ofPBmTnZTpw0qluyNFKJ6RYH
O8fvgcbwIelJjql4CfoZnPVbAQzWdbtvSXa2VYKtZTJPXt0ciWZe+W7THXuqTJ66
UkdcreeOu58u+oHbp+Mx1UtAyBG5ggwvsAf9JypvSM6cbhm1VArAvy6xR7h24+xx
aXXfybqITBfYJuHyBwOqDqVVimsrqQS/z/G1LMA/5NltGQ8ga27lNYXJ827kCDTz
mho9bEhpzjPRlTsTp0sycHLTiWhR84weBHO6ZUKIjGUAHUEC/jYMBZ8E0aq/rE3o
cBdbQk4nPWL4ROEPHapei59mPXMkp5mx4eb+JRlO1SaSNZ/TPaUi+ydzepWOlW6S
AtTGcajbK7PJuDVlHJLMgoJ1qRkJ2ou1gX928EbuWI6TXjwyVdX6ELssNkbvZL8O
S4QjS1kBlMangW0G6cJNDy77YjycttOefz0pDLmeRCsnVZo2q0a7CUPU1OkJTcjF
DcV/jE2JDi5kjoYAZUinzo0Iu6j+wihP5L3PAZ45ThfwQTUBZ1NhLy7kqygRjub7
`protect end_protected