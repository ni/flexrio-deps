`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 55056 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
akBpHK9XojjdOyFTP3pOwuy+R7KjGyaBVxNfGBhVL1Q+H46rKLI5QUVlPHjWoD3p
c2K9dXMzmTsv+1Xg9HOJ1Tyun0udFlIRB29GQSO+2wJQaBDdPEW9dqI6crIGsmvL
O+YOHSRkpJCzgTVDdRaUtHeqYofhODXqBTLeeZCbJ1KB6FWIS5cEjjc4Rk/5JREW
5himFDCkKo9bxE/A05VnKeSsOP0ZbcrSVC6MsQZVBL3PpyCsVIfYaDjFIq3T8sE2
BwJtRUWOGwJRJOEVeI6kkOAlXqyi8yRXLS5D6ylAmgHhyEGPSBFCBzHVTq2DK1bA
DpkCz8Xupyu5R4EYQ1LhleQn3Ohqw7OjAQ97cOzJ9GAXAGd0erVBePCiAutRJx2M
t78OJWj/NynltwdKqhMxTZAj762tBQNPqzFHgFf1e9JwcTnmg7j9otP8ViWGjdWB
T9IJySWeeclmA1kldhi1P2qU8oRJDwLPxDnMbqg9CzJMy8L9QUCfcqWyFOllpMsR
uM/XgSc8DF4UKLtcE9zvrBrLO28aDB8PuESk4w/70IAn6lohmFzN5Grvs9e2laKF
cPSOt7e6jlJjqZQSSYkCZEHzUAh6JjgJhIlMhEskroRasxqBcFmPYNXtSjBg/18H
XSAdQTB+vrJmrRU1r6VZaVCu5+DnG4I/x9NLNnLYZBaiKb7EiOLGypRIIV1z6+ml
57YpMykc4HJMkHploq44PsuhJjSBJfmszn93GPhuu5nLzBC/yATrvrL3A9WKfVM+
ZFuoKVZTqfH1J8+UPaQ9cNq6A4xwFid/3IghjC9WmunSW3f3Z4555HJv7cAv88ce
FHZvwF3Z1aqgpLL5IX5UjOzlhHzpLGOqoGjWe0w3sUd1zW5xudmwEbrWGWkHdXkA
uImoAZ/A89WYnwCa+fIBvDZC4mmykqtAQ1fG38qqCkQYRUU9kUkad9DX7mnYko1J
JUhhWB1lLpzwpBhTLKpi/Sv+m8nRyX7mzBjHHMpP4XYe/OTstBmJDQFeFWsKOTTm
VAQlRkd+u1zqZGVcsBkv52QXS+lPW+NpiL6dsahgvQTqZWgtc5/SJLaR24sqImKb
68WYjxyuaHvbUY1Qj8oi7rmTqY3osAq8L+g8/Z22FFp/xqeZ8a2KsaWbv2rn/rH2
+9FgYKY1rH7xuLdbfViL813mkh10PfdHrH0WeVtgtFXQjj5q2dF2ZOb/ahm+6FB3
6ElfvXy4BRbNM3cmtY+ohzjnNej8hGXFuhCpEjsnT2Czd177y3FRGqoJkJgVhm81
ovbSFWb5X7OjmzQ3zibMrHFylfvPjMx41VfQ3UN8cT5l892ePAH6isHyESKs399r
9/HCrgTUfJQ+sNE8rmhNc8G1PTIeKyIv8TIzLpUxVDzBgCAgFCuCY+UkIznEvHFl
K2PFcL6VbCbXcu7VkKYByW1X3suv3L37PVcg3BHLFaofFNiJKFTOiiuz1AgnAZ4P
kHijDW1qKt2R3VBw5cQMiToxFTDDxAauC1OWP6Bc3mZm7ng09TOukJXyYQnrunCP
VTlnJpR5SH5bYA4wRY/XftCixM385tr+JAFWaFUl8ZtR2ZYaPjsVldNP6L0QVnFV
SCMh2D7RfeQ8aUn1fBNAErYPA/u//tqM67PUD4xbaB3fOcIaAsUclvbPD52IKlK9
mwtSlLCu4b2PjCZIaqlleDk5X5mvNzL/qKmOVLeqt7f19xrh8xuCijhsqOYhy75R
/P6Ran33ybnHLbLVPt24k3l8Jyr7GdRYCmvRr9xGWG0ygPKmlLeyvfZ4kzlmEgTs
aSY7fYdJj7F/8gedfnVbpLQAfBBAgX51sx0OiSsZoDw8qz8HcVF2IWK6Tng5yAhy
3iK7JZOVzr4EXE+SXfLp8wh6hWw5qUsIGGFHgLkJhLbFzM7w9STdOBlOcL0r2Idi
ENP4iHSuSnUpzz9SGLhKSBpha3z9K6ClufiFPoLxQaBxUOgA6qPvrgl6vnWKNCS8
7CrInniZ+ogDvATGNCc3nUxCWGBWVAvW+J3H1O9M5Fp7D9DKrTi6azC/j1X04KZi
U0RfPxUyfarpn9Wg7St3NOinUJmGn5FhxmrYblpfG0r4AWDQrw+71CRKtefm+pHk
c/wt7O13EXw3BvXqoep+rlzK5xhReccWSvBIBcHViULZNszOW2Z4/Mw7dxdKbCsv
1V/3FpSPpAxEpg1RUuAo9alO6lKGs5kuxOBNZ1WOvm/m9wNVmXYWcgWhrOCw3NrC
stRxAW79UHwKSnMw56ujz1bBr1hECO6TJ+P9U5vGvJAtVIQyJdvW6+B79ep0N4oP
aUvE/tdNxcbJ1UYc+YFI1OkfEM+xPiuCLGy87JzbjuPiY1wqlRJzZ/CpXfe8CZYM
Tf2fcMC3hUAnNKGy5trY7YbBcbYrNN6qj7mUvdd17B9Wl1meyN8RwAtoADv8nRiV
1QoORpw2s9/xY5d9JK4wcBTsBgDv8fjmQ13biTium9NchJMxrzsN/LxfySlnarKA
+cc5SxE8ZA+y6XvRhT+EHF28Fz8Ab5FlL4WgNG8mkxHnwwi2p9Oyyk4Jd2h58ljc
/QCE4qsTgvSDjExuFy2KJ6rziezRdJuKfUnPPzFz7pTv29fYkMu4EcOpPVHJj8Jk
J8UpKnQjjP/5C2R3RyTtPe4WFiLNmsA3oS6iYQgbo9a+qYhafUnPJQ/B/dWHvOsQ
OQtM9STXN/d4JTE+ShdKpVp7jc5DIttvZ3LPVo/mCG4asq/GxWmzJW0TZTEMrHrR
o/dLFYTz+Cd97nJhAdT3W3L16rZRdfjrdvWvaLTk7iwuuNtUuAecsNefaL7w+pQN
sP4wikVyWBopJzRcmBhcjLQm1ukL8Flx7PtrOsdDZS529EhHlats8sj3q0sVBF7w
gSdnqnqOlu45TQkBkF6vC72NXwTKahcHLRSp8n6mdN8XPC/XESULNrI4re/6ai4W
OIeVwm/RPf032VsX/+9cnr4SXaxk2GHNj7MaJe+W4ueo6ray/XQYDvk+CepBDsnd
Gr7a4mZJSqNykkaNRiOKBteMsUDu4HqXF2S1ZJHv2GwTl7BnvZAlbtQ4DfhBfpTd
Rr/cSV3bgzti99an1/hVSHjERH6BFpN+UNl6tRcGxE/QGAfZgLITl7tfzNOzW182
A/Ea02D0cCI0h69zxKI1leYqOA4m/y+L/bzVh4sylnnx36DGsm4NL+X8puGblFP4
2BrWT92VpLEBb4fGKvuz8T2ruWXZfpLCBkcAp/F1iLDxPVzMSkJYoH4Lm4ziBPuy
fvkdRKpbrXXnHXjdbCkMTyJ2k/O7PiHDfDO9OIP0nnOFUcolB66VnNu6WxRojz1+
7arV46t6zErADLi23pofqAEkiQBO3Jmq+RtnCklpV7J++O7jvzrImg8bPNQcan60
zBKbSzp+lhRCueeGFrDJ8YC+1Dv02rRN0sjj9r+rsXvBUvPi64aJrxwhh5tm1mIe
ntV3vDQ5+Vv/u+73JItW/bOHg+uL6FVIQz8otxjpn7r/7ikwX727E5LuAOEMm1OY
brIMK86KPlNV4oO8RrR7dU1sO4sSqTeTDsHcQl9TboxBHBsmA9YbvpZT/JQedIge
Qh7rkf98q4shfRYbHPuBXpypyHqP2NNhoozqlPTL2RmlxJEhjUgL8MEjr8w+wI9S
PxZl9nx4jamvj4FWndnjEXGXa9AuJoScYrwbM7mPWG+gCVWqxRgPUZ98PlsMcZbJ
FoPK7bqay44UT4hwFTjUPas8+X5esZ2PDgTfL8+5S25nXrnmvxUS4oPeNNkRHoMN
gID03zFFJ61noTbSh74gICuqTgzlFDwv0jrKc3pMHBivFkv6NDRcbItlFNsdpt+/
S4QWFiRrOcqPcprq6Vgn/trRjBkpAUJDkouxpYNvSEBfNpPH3gkHiL8gfOcR7xjh
XnO7FzkWWbH2E/JFJn11LCrcErkkn5qdzynSGeWXPXU8qmGx7dCGHlLaULH2iZ0V
Vb4nxd3A0xkBNk3D1/4hjQXp5303lOI5lp5rVT2El6lzyCxRCyC/cre67QzYXbtJ
iZA66hygyqrD414acHiCNevG+Iq2Sj4riQQ4ArM4XGzO26p5TiL+19RIhqivZalr
Cr7rolB7tvTUdTAjaTpIluAIN5lymcfxaC8x1olZ/yKHzMdTTp/h7eec8dmQPuZy
0OuLaQlEMlIdcR8cuODiKT776dq4JJiP2aqA+QrJtgwB55f2B1FxaltF6fiRbsAa
gmsnmYER3LzNP31RMaDwDtgNj+PaLNFFMYqJocnZ8HX3nQvvWE4k1cWPCEgHaA2O
4yUO0lyYBVZMnGvO7R+TvOL/4HIXAz2l4tKkXyDkJK3kYLTz0dW7HR6K0p2W/+Hl
kJ4in7xxWbwfG9Yag19wda2xV+Vee5wV0VvUob6GAVZqvrq9iFNMRDxTSw/Ip0dM
A8MGj7ZOycdg+5MHqakGLPFpCxRsOH1g8CCRKDn8jwAAqLKQ/TCEd3ri857Q/PMV
k4RJt7yVvc7eqzQow+KgjlW7/oPq7XR5p6XuVrfgPuIWwsfnb5S0Fm7ToRsNcws6
8hOLOi7BDRes/lJCqvsI5PJf10zzMn4v+/Yg1oJ1MospNgdIUsw9NEEVHQEQsSqz
u37iMjvEMSc+9tcnbcvSBM5qGfMqcqIA+ikgT7Yx+FKCH0pt9+PbCU88PxnHfatd
d7HDQw3NyFKXZAjluPFaihzl2XtFPGA3/hE1ymOTSLh6iPJOc8qt8dQ7jIOzuwze
ehcQHfKi5ZPLHOTrAGyI669xnECY9cmvzcjtCuZVrhowGu9eHiExz+278tdEZyNl
u0InpSdPdHz7HIGFGiY0wevK+zVfcR/Y0uxPwLj5FAaBbYdsIgXHjMj29JCuFTXz
gRPok0+Tgfx/2ZUos/VGtS01om2vTlLWCWGs/9Gmjo19BBSZiOgVk6Nx/MRnZILN
xR05PRtfvhr28NYKlB/9t1RnWCmSHQXSCanaEaEZQn2wb8rKPH+qdWNjDZ/TnKP3
NKUwNGBUjlMm+hZ1nwLehYyfQeSjPJ/3Zkhr8+WcVgcmXlETYLH83oGVgb930aUI
9Sai0jZZQvFsZjtAo2SzQoeotx7faZbwNFs1Ccruz41nQwZIPl4RD3cHJo1hqaRH
AgjjwC0FF+STtFwbzd78RazhcmTfHySmh8SaTMSghKv9hsCfxWHDGmxTp3Zv10cg
e4LllgLLsjGwpYRcGsRwQaOkvBVSFYpcpT+ETpm0FXGLV8xuKlBFpF+zsaq5M6Te
99U+BHyJJmrBqeh3DadNhtq6oJSu2vv8X0RCuSnw+AuOEZvGx9DXNNkw+bMm96Qw
1tUHHoYntP4ULImmIgDbSS2m0Gd2Mr/vgCpuVC5uH6tmb1dVT2t4LPl0BTQVRJ92
RFxpiweQMi/TkZ9hJyywRbkBKPvSRoVZLUt/8NCtNeuRm1IBwsLuW0MKFuQxileW
WSTrKwupykWDlfdpWzTeOPYOQyK/RxYoLKb6U8pZNMj+NAk3BUKJGDjxyJxu1RNf
5AByUhdcozNE9UDQn8cWJCuu5qi7D95WeIfqX6ne2v6L9FyLA+bQ960T+GVDmxmW
ecI7jon90dD7KEw9kXSZCATGnmiTTaubtJqZ94rVdszOkVV0XY6pDpD9bvF4bvt8
M/x/9QQcpFhRwXybhhpPALonaXSM04z31efDa0K6HXlNWwH862OHYqlkxMtER1Th
APkShNO+vz8Di8kCC68D0NdrAEX09KrFSu+O824DJNQKO27dS8uO4QKKy+WZAFXM
R7rvU1TUeidtxp5q8ggdsGTWUGWUndXKGA2qBq5cLoPFd9DmyRj1GqSvhY04XeGv
/7as6u6aoxeezS3NSvtKRQinIVKFiqoKwHJWoYv+SsA4Ufoc+FsLk6cWHmuE6WIn
VIYA47fjJNUziXAO9Uy00LobhVmnYmNNVvR9Yz31FOj0RG9gr9PfPeXiJ4xRQz6T
5gSzBIcpD4QmHIFSWFgvhQB1yZ48ON20b8JYEwRXUEIocfrzfi3o6S7ZyLpv062j
eTCCsOthbF2p74Z8kqHCPhgmiOJjQ1BlW+Og61b4y55U6ZQLy1lwox4kRgPRydge
mcD6x+JDeP3fhktcal3xl0bgPiYSKKmgUGwIV1VhPdrz4labUYlOXD7VlZC4gWb9
Yz9MJUElPpSKYL2vOgu0xmgQXb56wIQUt3+ModiYnMvXfMrHd/p3OtMo1DSK2S+A
6eTV+LB16XY7tso9lgYnUBfzNNKisTLSD9iohHXf/RRK19LPWNAyg6Ix2qM11ORd
nSNdZj+05T7pbOXTaiFVBUJm9VkTVnhqNfANaz6Obb0+thQ6qHgHrtQ3+XNjky6/
KsqoCT3Zw54WgGwW59rrk33qv8b4/5wZFpQPlUOHTRCyiRbPfLrvloqNRSUo7Hy1
zpamnX4I2EibQk9bBvUgulscPrZdB0FHV9s2hbgwcZoubTZ0HL8cVK4oBkliOewb
ueR7ouPpcx0pwb2+NUBeHNEBNr2dosXShVtJjMgr3mgFcN5Dv3o7lG/SermqCDDl
E7YDSXLPbsNrmbny4vsdiddPvD1vL7PJSAsLCGFxhJzvOgSoK33lFsqWsFKFFGIv
h3xmI1eYFGSU6RzPUutyEyhbSPNyjnisyxSLL7Q8aQjZ5XcIasR6t6rY4X17hCxr
E0hf0DEpjpUmiqr9hSVMKukAZHEsqi2WxkHCxm27R2GVU+TPD83il162MpCMgzcm
BxvrJJrWoEiQcrtxGRqdSVXQ9VHsXXycUz0OkOZHwb6gutn8mYjbbs9FjzuGoZ3L
BrDdBhgST975Y2UVH4Y2XP898WcTQLZQ7E113cMWWeiXoSuQIVajdnI/lPhp9l3v
8aWmJWOcrHuST9ALlwOMiAavuCQHGCPicCwq59bSCUkFjUkfsCKEHlZ8WQ8kXTI4
wTOU+3gcfHDLsTXvQOniwq4pJsUYGfdqHWYWmm+PJRTqJYN0vtzHPNE045c770wT
268VyyO43jDVBurtV7BhqoV8QNZ/JTstwUf2D+68kRYK3ckW82n9Q4NAw7vuqYS4
UvqF3DHG+KTOuKW5UKDkOeZwzIiHnqwEbE+cv57Zz9k7nlZFA0ETeB0r4PDT0U+C
8kBFVmA/cC7/DDpjdRMS/slPe36xeUum7fbPIDgwzqUAenDu99oMce1UiA6yTOOA
ZbZlreCX+5h6wpjDrI7C41WJmaVzETyqyxRLpXHf7it2a+EeMUp9Pp0f/Rso1Qau
4PkSpBEYcl3gmZIL1lnP1KYTpiGi8UkgD4kwRr5jC1WdXczM8jY3+YwMVREtUf1f
z4nroDkkAEhNLlQqmNcX7aai89kFu5e/FcLOKpHvhb+x6evvjYyISIkqetAmt+l8
ON5QEdPQFPtugrrRd8NnoEM6cjs8ouEAFAjRdd0hDUuCOtM/f2uvGqXRcj4UNn0p
3JfJfJHufc1b38ZyLCHmqJ6iUPucpCtwJJhHGYqvkTBHQDO19omH3UlZ0/X0c7Ws
g8NJeLwHLaI/X0WVSvKkddKB15KxsbYmSBPgRObxDMt3I107JEvEIl9SV1NK+D0G
pQ8i4gHJtuKAAAwIownSvwIjjxlMTcFGEZOFY3UmKFV6so998wR8IKaHWyySH/iY
o2r39sfX7UBz3oIoMWqYqI0HmugFCmTVLH8sZSec5qyk3w8KxtF1wD15AUxUq9ul
agNFvZiSL2Fxd+K79L4GZPP52rnjH0YfRE6TE3fzJ6ZymiyJ/KjpGc9+HPjWHE1f
k6CszZXmEzXzFYMndfiBTnx9Ks95FzXpXtYN6FDiKxyF+Rz66iLPNrkKnuL+JAvz
RJaouBRyVx4/YHYUsU4M4UwusRIAPnJLGMiTaLRuLXnaGkXrnam2vekPV/55lbHO
YMlUIi2TX6dvV3MSzAHIYvjOZE8/si4IYvKBE9ORRVqsPtMmKDE78yCQvg5pQWjV
yJOvbkO9SEfHl+lvpAxYvhVEaCILbjd3GrT4Ggl+6OtZ98joGF5YFVSOt05UCtkX
ws4hAYiE2maxknPMcxf2LK4NkkEm4elSYgdAYeYjweBeoYKDSsDCYgqFwf+/4qu1
LcAk3adq5LfPAW8I/QoLBbKg9S/+Mbd6LgleD0P8pmFfVyS9KASySluyF8KIJZgt
Bwo2nQ3nmf62d6VDb5JriZP+z8X/qIgfZQiBkOhVZUEp9BgODJVDOzn8BHFIKUNp
i2V9oG1zUGiW4EfJ3QibwOoP4jqqnYSbEjQlUSvLMeE1X1W44zGUOrA2B9IYmlPR
3zP4PjV2aq9wUEgjje0MJT+HyDuPjhKqtrzrrQDhkSBfwcklYrnCg0OBZugH3BQR
l3vVP97G9ZTa8SqOkM5L+E+5eWOjocKCT6uHR4gjxdkl2Hd4Gfjegwhnw3I0EQST
7lZxKjZPU/DPAsa+y8wKrf8+F3WKIgmDDxf09BKCxhIS5sJgmoIF4NUdcrC4VRyE
miuAAce8NBAC/ITnoZAg7Hg98PTxi96BoUP+7HHJ1jl0PFpxuMnJXMckuVFYmJ2s
5F4DjDEStgZMYUe2ACNXQicQ2r1iW/OEPuySFMw6dBoASe5wFiat5mRyKokqU3uY
Svw4gZorc8j4mHFFHvT6kGxR54I1IZjLQRQ/WQH0pDk6v4VuhhvTDc9tiZl642bY
FCQ2fLtLXBfyftbNGon2Th8GcHsd3RlUoa4cN/kTiC5llX8Hs5JVCnI3t1IALnSQ
qxRjCvLMjUa+smL3JH0mIfKglkkUIigE+ia7yPrqXcMVMIeWlPWiDF4Q73LwjQdy
SyxhD0GVI+YzVvY0LtZJoP0vRi7lDZrVlLw7LDWRVwJBLj2Osy8vOx/6zl30t4bG
v8RXaT3IEaEpD0Jna2nL6EiGmDHjf+hgQWR9/7bBKnDknGC5z/DiVpyqvcaIn4lj
pvTwps9/oaU+m2BA7Z+evyQ2ctkdPbJeopt0UIb9i5yPFCRH+MhguvVrV1bV1TC5
UQjBNaOKq3ncGhR6VCX0wtpyrkcZaJIbWLGcF7Tq3lQdMoBV5akmrMNt5gwIVNKP
N8W++s6358Q7E15kXRAXOEL1J1I6jnG4NZjUj+HeSHhRsHEbjBz9XSHq+8iLiqwj
1bArEaxQcvUbc0cX6/x/2prTLLIeNrGCEQmq4caDz+6DL8Bd1b2CAM/OkuWUt+it
eHsyIx8zGY/IjE7d19gUqnI97qJjhQz4R1O3iG04Pg10IBV3tM/tR7nIo3CytLvz
BJiEc3yl4nzgmVOs16UX2NKvX5uKcjqkG05XfQrepNQMrto+b+elBkyGz/NQ/XQE
szsPYcb6H9HY6eAq208w0od9JBEYO0QjXi48xamZrmkWy5mRd+jui+paQrmOr/sE
6oOuy/90AD7n0eeJ1L12eOuXjEOQe5oB5bxKUddMvmhY5a9nrb//JEk0z7Vy8JGC
3ytHTSsXkmtxPqxk616mjOFGSqSTn+uOrnUqnPH5DACNaN+gtMkviE0zoW0zIonO
f3zUUt8GHQ9m/vDCmS+uqLJojYtUKoqABrWNCCrrFP3kBacqeaBBWvQ9k0YpIX8k
xOiv9YcdCTXI5tjrIQvaAuH6qKdbdhVk3P0lZrfc4aMjJgHEO3BZMmbuE66VxLcn
jFZvXNjseHnssPi16XfSDALGuybzcRiBHhmVfyCBD50ERYpqVGr/0msSP+SW0XiA
qjA53+2ZGpXCyvdpqIEfbcELonjhRZmwwLvb0qqWgdjGGGFj4M2/dn1L5wHSp54R
Cpi41p7G7kUiwvJhO9aFcV8i59V5FA8jZilHcl2ZYOjLWmEN2PR85/Q1Zy9K2ff8
jwGpZEHaqtFe6AI6yE1HMY0YcRCnmqqQ8uFqwgnM12QwylNKoO6y3651lJaWXIRg
srfu+WAwZJ8sAyuI0rrDRg6G8W8ZYXaKLZ/eWy636rkuPZWLIcVjLqELjtHb/YHC
Umd19tV4/zWlkf70RXwhVFJN5JAo+sQYL9DZFsgj/BEqBKEXwT2pZGexhCoqZWuZ
9YfL5waVWC4yDnsxpFsfzM2IpcWSkc7ZxRcQmu++1wiy84NdGHdwz+rrEkUS93Rl
IptERT/9BVkbBVvzM76H2uPcpxDNau6VcW6OCFsIDQRGeINQ3OS4uJJAyWVW6CSu
smt6zu5p1TPrhVuPBsxDk4gXLdmCv8iNdeDkCPjZ5/7mkHD+X1gxexUn2kt+QyNc
Eo5nevIGh+2+DdvFOW6bx+xWBsFxus74BR21uex2nrzVGrMvxsGP5cU9p0pjElDQ
R0FkhpvHWGMtyJYf9yTGw5VlTl9O3TVV7eInJH5Pvjx5nDiYf+0oyq02b8POdMK9
jBR12MOGCv/jJ25FdV2bp0wcugwQLzdSS/TZYeDbwmeMA2mNlkAV+nZbr06c9jL+
Eo+U/KVcOsk1PvqwNO4OugQhfog2xMiGCJUpld4/KB6NWSLdNix5W10eYKrPnWxE
jMSe4OGHquuK/LU0y1I3x0rcxY2BHEznVimJphDRorbX8jZqzbLll+MmhrRfVLTM
X7eilPDMNoNBOP+lhdZbRDzF+cOD0t6/3Z2Wz+YqaTh8GrWfDiDhz/wq24wEIUDq
MInTyS+jAB1QcmwBbnLupes29eJr0dj+zBTurhF1cXrrwNSM0ydQR5T+ee+T/PsB
KzkAy/2klUgpIUvOJKmO6yyFvahzEDNKQsfM/fBokwm4q2h68Rx0W6Tba9ny47f+
YcZn2ibaLkpbcVKDxKwqY/jOTgS0ifa6PR+KlOgRjgNIVawTESrkgU4s+Ug7Lyg0
fvj8mg+DH+MyuOFLBcsSvn/MI1KcDzNT6a1i+2iiUFXBrVvwpFzs1K+h5/iVtEtM
/wUr1zA33cOizJlD6hHW/3WYZU2rn8JR8xi9gFTVYPcF1kljREIQRfVlPB2feVif
FSg1lALeiqZFU3xbU0qJcOuUqTOLKAYeDlud8DO0XuPCvzHrd5Egz0sC0DxpBfvi
KRONWFE+h/mRkbMH/f4ht0HliVnfbSvHMIXPQ+7AoHEdY6NXcsO54rjxTWUh10D0
hiabJOCz+J0Wa1K9UlEK3c6Y/q3+k0RyL3tn/LMdM1ih/ZSKEL46JBPq+iB3C7/E
svsKJjwtOy3DjRyruowWm0w+Mg2gv03PBQWzY8sfK/FQhcF9m3gpnac+pjKHP1wQ
fr7O7LrpfFIc7Rgp6MiJF2coWX8gjl8MVHThkpQQt1MlSVMALUzY9ZdxD0b7lMeI
cMlRAv7jSC48gSKwnHPqtq6AKcQ/5Xlf0bZ/nLIiMGTqXJWyXoK3XuVkXrj5iIoC
36wOCorhgYKv1gZ4G09G/9Ip9QKiFxprboegokTvtx1JWJklAqx+x8D/zlIye6OV
7/CJ2suJK7C9xCMhoXBC3TB6bK/PghDlsf+3GXruW6BC04pV+1uhplqXU2m85WEU
/dQCnOCOnavew8QXqHEApJZxrUZ4Xmq4KqYgaibsjNJaTRHwHNkdSlaC6pisLOzp
KjhgPJwyVjSg+576zO1tSuuC0DP33X0zd2s7xXjJ8FqXnedy47Z+6/sC1BoVweje
PzEQGHCOOIUW2aTTAVjkMRozcfT01D/hAjlFheNhdcXBaptO9Jel9dpr+SNNG+py
Shu2rUQB+a3kCKfPBeABNUc/7pi6osUedo6Rsf/2BDFzOpvZbPjPyvsTQMHpIiNo
MBp4/mloT3d3h5iS5DVZg1USfYkVvi5qlfR1GGL8PntT4WEpLDGtFifUTwIDTBCv
6l9FFxZB2ZgjoPtJMtVx70mJJ9F1boumtfPHAZ6qElfmjtpwdBa3F4OSi5sgdn4o
crrJGPz8xZEijHaNw+ZtgXaF85lqk7yiMAYGWQnvF72P3YFuW3Iqrh3AP0/nN3Fb
4NOi4O4heHz6sS/p4ulLxPSHuOftZCAP836Yn3ax+FJcHUGYBlyx7Ox33h8p/3sA
HmJmDN6Bt9DwMcj4pNz0D4HLjC2yAKkR45Km/OVd66EQ6twz6KY9GccLGMTa3EKW
H2l/yhD2zfQX3AgpKhh5dfRQLTyJg6T25k0JSJ+ZdrTsv9OF92K7hQqkHnv4B9fu
9ZXNOqCuPAbcV/De1zQclZZzTyU+y8ABUWqPAFbMUeCPmSiytLnxHfKxWxTS/US8
zXcWkiGkMjZt/arUzOAvhYpTzNqD1MWmuK6Qy6Y9Jbo6V1TVdSA84rCTPzzpyMWK
Ad/x+EMXT3dY1tI6X4m4/728XF7nVjvQMmFTqQABSq2yABAWiDAHmnhOpVwFHVEq
kE3EnXDUePmYGHJFAc9TIwjbJH/rE7UTlYsZaEtT0fQeps5OsQIvh/Xy5/n8N3+d
qgTni8yCFkUprcUYNaXORABMZmDBkLL0TRIVPJhLGbgRnCMrGmW1hj7XlNmuRvzs
ijXi3eXq+rXfOrzLYDRZcnciZpZcOmJp0BtGhh1BN0vJZuLfGS2JPq1I7Zw3Ayd1
gY+LVeUBPcNDc3EjTWsRUyYTvukAoteP0O4F8cue4gO4dXgLJn8O/U6xpxpqnjeT
lL4m98NbFZMmQ1RXMOUuKDFcVYKWef/InZ5HdvePgt3o+NL8s9e2na1YU8gBtiyk
UEF2aEeHieju1+VRcIkfevpO+yqyBA7U2gO6WkvzTSnUlsREj6IDme6LUdtOymKO
5i2JMSwxA5OsrPaWVxhZOTuzfxVcx5a5n2Yz9u7yWUyaYKL548Ez+bVrc5swAHu9
tV3mQQ8cSTlNf7e4ybZtOgtMa6pXxHunsBhpzO6W4stCQC1Xczze7sc9uuEDARiG
UB6b64Men9XKmw9biBQ3rCQiPylCQiJysJihqNORE33+f/tA8J2FKnBeBlHmYRDz
1hrs8eKrLtROAh8Og3uBAqSjfLmkmT0Yddcjb3CXb4cEzeVXOXYXJVRs/XiVYSnP
+NKR7QNfwrvl6IZKnrDb9QZlhujgNm7cC0q99wbs7RShAnQ9C1mTlSaZ9koBs5+J
GM97ornJFvHOjcIqMPvW7YyJQVaZm5u83VoSZIkjHWjGkW7okJB97erA3tZ2k4KQ
wqZsrEG69+jB5aSKR/SqyBzw26bIkr2f+BBx+x4020Gq+wgoffSSCSNkqaapAtn3
zIOVu5ZDgO28t1EqlvPzPY058jnxhLNDU+nIhOd3pol9ZuubYMDI/tAi531WfjLU
lwAJRGAZx2pC5s++gOPrQZ0zFcU+Babx/8QhnHfVtO41HJw6wC82T4uRoho9Fesv
Ly2Nzfd1OTWnWzSsMSem3cwtSJ5P2fwYGAcfFVdVirPZRxdbpkngb22ApFGZDl0R
7JfQBBWZ+rDA8Jo5yzyPV0frk527o0l8Xmtk6g60phxEH4bELdlaqUYgVA8VXm8J
aVvn6hQdDDxx01aJa3a8TYACo6FRu6+AX75/gkiz3avpZ3DU34ICl6xDUkR3vRDa
E0O/SpGyT8ZD4/nrbnBCCw9nG8ywC0XV6UUjDDffqouSgeQSdUpEp6JoBh/7iPml
fwKwsAyEVnfItR2o65JI5oGS4hy0ok8bIzpxI6yx7ZFJS9stTCL2bEagVAG7j88t
p8hpihdvi3rGBe2Rk4sObcs73ku4Nwt2M7NcRpdTR+T7u72MwuQbgkuv2PhnZA2I
Qn23F3ZXBMRuLScAWU/pCsDOjB0BX+1B82T8w6J62Bhkj8Kaa00lVh57m6Fyzeol
9J54mAgO9BwWqPBge+CeOOtGz4nlqXyH22frmFtHNjf00GxOmAd+Mvh+qd7+fMyM
Kb/2nEQvI4odPG4KsDbBl45NctLDBCwEOspZfBwQ/FEBhfSck5g0F03soohN9Kku
ofgqw2BuBIC1W2Pn+vMscshj8OeGpdrrJG1a0Xxe3Fu0kcGJsA39dSwqJjqW3QH7
Rp0hxW6nXmD+QXgbD2mZpscShTEaRRGcWGT+Ld0gzZ7tsqB5A5DjPCBkhYwnkteA
qnb3LKCh6KOglUBjJE6UyRK1Osrs2rOmmdHnyBRK2xiByFjh2HSd56xPDcHEznnA
IVFpf6iNjuR2h823DQwiBzkallfiOWjr2q05doQzfS1XZQvDHOz879v8CPjU3ZdW
AdwDjzo9G4D4Gj/i9PM08KCoty4JQZuHR/gquAmvAIwycNyVWnPFB+lgxKkw0tNH
HMeb/gllet5CQ4IJ1pDXf3t0OpMGtjjOdc6STPxmPzpGUB8lqLdYgPwQiUcBXX/y
je53lJ4Lf183YzM2AdVjnY/bv15+mTStU30EehTocNl386gNZL+E3YAnSw0Sw+Gw
1A4/Ck16QHc1DQhilnNDUDKTINaBiQqReIJ65vBOCaTlo54exx3D9EvpUQWk0u6g
gGjmJMVoBH/aPbfn2T602hIUj1vsP0xknGGsLNYLKouzi5ct+JjPFRn65JkJcbYM
ijud58Wd0vlqMfY2ykBfCYvuPZkRpiMAObbRwH/DzkykLmhyDtuQZuxmAOhTLIMM
Td4qPKDCODSr4PMTjlA4KjxeayORe+3en4A/bojM9DxDm18DyympEGL2S6vtHtvF
wQGza/hGp6mNA1dwS/tON7VdYJZAdF4XBTtAaNEN27r6PTwIiVw1Qh9Po0Ee6baH
IsB9KHb4jrilKu7AHJBZq0e7FPPY6QE2Jj76KuzzB7Ttn3BrW4Lnk1shBPsNQTLJ
4QracoWfB6xN3jkMR66Vg9PVpmODshWKY+waeNBJtLCywgXLVzm7diVDHpQps9qP
hgrRyih1X/yRXSVEQ8AN2eP4ysl+2MUPbvYDNIL3lzjz/PnJ5QZVZC9q4StZ7UGb
LCZF7lpn0ZbaBGU8YGiu/f2s5yT0bOSurcTF6F6VvSGTBEDuBvF5rfR/hZCuUyqn
2xidDrcixi+e3IF+ne7msmbSO+aASFhXZj4ZiV+alEuYFvbLIiR39iInh/DD1SaQ
y4vgKsEIROGYQNhuhlgGB6P+utAWtT9VJNVugAfeN0Qfa+aqVgev8QNZbX8C7UD/
6JcOMBjbHnyope0nb+PPHUwiZswuSqzabfotFMd8U5W6e8NBNu6v/VyMlJ6upHIN
b3SfNCTgslMVPHApFLeZN3y7t5IV4CUaQNWOMGFQZioPe0w3f0S6wK+nbJ2C1JaL
O2obHVR4pQf4E7eXmxmEWQtpNR/SulcX1AWPhi7zSYNXvX5qffJqj0zrQonHFdmq
W6d8rdb6izKaRh3lUDz2J4vI1cE+yPPeEgPWzwXIfVbKMb2Qy4iIHsqqjW4cYG4G
XQXmSIy572cEFchjFeT5HMfQe9NhUopr4gIoqWRtVXYZYMMaLOCrD4cTbTzB80Wd
9s9c+qtpoFdiYElup4rheJkbpbzAgvigwjfNvjQLELVi+Yp687WZrqg4NVyyDceH
130IlqxphcIpM0LJ030emqX+k17X8fgC/Ncf2wGE4XUNlxLziBVu8pMPcPfNlDPT
XJiyIxCycyAGf21dHoD8LfzjLy6/HBBTkZq4N9dt6R2IDgTCIph/DFrGBN9003Db
UYC5dFIE187I9GdG3spJnD5I9yeopFcIXliQemvKseZzjAKyQr+hIY6HtWfCdejq
ztCAARVLnxwcU6Z3pPFXnyCYVgIHUJeMOrMwRvXXVXO7f1Gf8aGjFqw3tnA5BcfR
J863Zc0eWY1cWVIqNRRhOe4LFvMYUKVTqTd/h9jDtr27si6iMiXCzE9vQA/PHVQI
DuCOzzV7oW/RSaywwRMA1YERy++dr39sUzhCA1SLdCPQhU+i2yfaB6rfF7ZAlcJr
1XjMQOkmK7T8VSxOsjGcN8UvehOknM7lvYaUBBrmpz1J9Y/Xc9W+bQ9aO+8kMShF
nlzlSrIThFcAiJwdH/9wuVJ+BYMfTrbMkRUkFfHLkJy94O0ipP/I/vK5o9RXHlA+
SoWPtP1gizCc98vIph+Y9y+RaCNv7Nq5TvZaCzhBBZknodfShMLUXS1o5QLSM+3P
OcSD0QL7prLbgeStu0kwgYDJr7OVbDxDBXeyl2FeYqmiid3zSz7O5FbjpIdzlQvz
zHYLdwuKbpc40ew91Ypv5iGGimRRcs1i+BGn5UzolZ09dMMPKUCbxxFt6Mgo+hY/
RLmVlna6MrizRokOpLr7iVKykTBlG2618/mr2a9ddF5ihuZP0OU8GEFCmfpvNClU
XEYqywe456mqs46rn0UOoNbbmI8wT4uwA1p/Q7ixS6I3pbs8bq8YqQplllGn9Jio
72htFgynORPVXTAVf1g5m+QTjsSEoGotEUo8B1RgsSk4u2+R/Xm0QToRQK1ET0Qy
w4MORT0ZQ3mtIpfcqOQ+eNJjNPKf9f+koGTSINRvC1grVxxlQoGeKG/et56atwI0
fmikoSfvnLT8ftd//GFZWJGXplhCNuZNcTOmtBnnwirHQrUMDhSeQRuQVuw7B2+Q
PAo/RtGRfpwZ82RO8lruqCmOGsSh0kai+x4kK0szuh1p6/q5jpVefHAP9OC3AClz
CUTeT29s677mNpCV7tIy6r8STlolFSAC4Ewo2HjSRALppovViPPczlEvlpiYTBw9
ILvIAYupukwIdziSVlkyOszZra4bvP5w16piiAGx0D8t4dNCY/VWhHEqO9Rp3AZZ
HlaG+pHC12mkFfFzaDAK+w/GkgNwB8AFidjZSGBXM3G+PWBpdQrLfxQdHDyqcula
l+fSa2JPF4RY28JBhFy2UVfyUcTdZq9VXIOolayWU6lvbpnua2eBltfR5HQpT3m6
muclCRMV0bhER98okKLOALwo9PQ+IKjG6oh0sW+ysZpVwYn+u4s9AdTSW5skXQK6
MWFSpCZT4dX3pOPhERQqoqZioXAmYLooKXIutI4fO2qwkOOSg6wlAk1oJroYpQxq
GAo9clFnBl9TnC6N52YX9mIWY2/M2awxKV6ga4OiveJE/ewOX/INglSUTWtcpREW
0lZt9F1Wl4mdkGFREHfOXx6ByfZCZlsbSjfcbPSyedjOvI44L5V1birNsYHsL32o
frPOgig82DXZ4Ev5cJ73L9XUBSr7hpgjse0+898a0JHxqV/DRLdX4PM7hG37eKSz
C721h/0lJtvmiFwNGJ+E3allXmOpnpghmJFVRYIdLOyWYRWvFXd7sSyIyY9/wrvJ
DkElvFb3vJgx1VM23+cpYU5wHswdFlp76sfICSPgM0M2Y+UUF3xBXcQZov4oF+dd
wMZYxoDJv3NE3yWurP/asHSFNXJzz+K6JRG7De45nC2hM47rv5CcPg/ykYLpFGN9
IKhxF9oLPYqvi/HONDssKfdrGPEAjSCW7K5b9kDIZuPJfg24C3U/X67gfEJzik76
YGI5qgDjbs17CbPJR1aJ3XxtJKuLfMTSOp1scztr2+z5X0fQ5d383WZZs+LluMC0
kGyIwNYj+DXdjMjUobVC2GjIMsmNguQQT9/VvsmWhviRY43Q20+Ibblu5j/7+SLi
z+j/GtJiJy5jYQu/0aTN2MiLAxfDrp6jJRhuswXNz7IFs/SkfJn723ANAcJp//Hb
FYJWNXMLzKHFt3AeOZELrdulEzAX3zmvfUEZqwzI/mLfymAPfn5EVeFJJBPwzv1d
sBA3yS/wS5YdC7mv705hhf5A2mzoDgKB6KxuQRx9r5sQj9pgdthtASa0TyfZrQ6+
a1cQ6ih7q4yZRSH2uygFmNqkd52dp1vXMeyh1R1KB0BMCJ708aSmBfE1N4sADw6M
CwbVw1S6tW+heIGwnuuppz2TWgvqbUBP81J2rC5imnRcaeL2Ncflc/tEtm3RXHhW
QrkQIrXTfnw0eAsQZy67nS4n1Gmpha854uMkyXtKxYLbAWh6uRDjBLLGIv+qoKFw
kM7Pq3iluhHtmUfxl1v0KgpuNbBdTjLLyAUcM13gklWWzQGclMxiwCvJPQzzl4ja
nQZaRmGVmvs23VRpWComBnXXpUnYdRdzBtPOmoe/cYcZvdUSQmHQuBn6/rMhtE2x
FWtC4vkS5mTbFn0f2Fo/GUvPbkBhzzgwnYeKclOV1KNPOCAdeEAwDciGP1XWxbaR
pCjSJEv8k+jS96DhAFQ3KSCoP+6RgEM+BlNMnx+jZU1NDWVvJjbJuz+fc6Hf3tEw
DkWhMXBznUF8XTZ05smGAM484z29uWKKn42g/n6lR3lCgd/EFI1j/WnSht70s2wf
hi8OOSaZeVQuIAOLLQbh8eI4y39Oij0mMSNnXG9THhURmhOoAk5LaZt/bRHx17KQ
MnIp5t6SJGGrwsoTinw+GtHO2wtXI4qYh+/ViOe1wDe1d3acVyBGjEfLwY+hYVS1
fiEhLK+Rhe24LSfqjVu9p/whCwLUVbAF6VMJg0pJEdeSn7x96pGhYZhazxQlqNCA
ngkLdRW97L6Evk8uY6vJSrGZ1c9Mr9c/VyoKqSGJkj2/pcJExgqtWjzz9/a6Ognn
HulFVx5yyil1j9en+WBqYSAIIpOFF7xFiykTrw9vzgQaNXIJ+bdLm8CR1tm6D9v0
0ZKFRpDV2lbW7CiaGg20h0FgWMDPLipGdI+90QPbAabuEWUBCfS5K28tG4pNQaZs
CDZVT3bRzSMbmhNM0uALvswIcK8WHgpEOkwKZrcVser7bMt+2VtgKOgE9yRLGUXh
8sivxkmYhnO8v15dhVznmFla9jYGmYtvvijkuV0AR/re1xuMv4be6tT3H+Kz0Ugo
74YKOZCx6/ixQDPLzaZOg/lkNpJlvM4gtw5UITrCsenk1y8sXZRqDh9PdkBaugEW
gtHHZjemYNZbzOcq470ErxvcIx/rJ3b0ZIJLNMkuLnWjM2oCNAjl+XvMJi8wZ67i
8fTXnwZeO/nbqLu+0jIax3zs08bjbYKBQttezrNA1rewXabO6lTp7c/5xOyiLCIP
ZxvXDp33DwuryB2T2Tc0HT6j/hK5RuPl7cW7I3SjWj7TvJDVrmr+ko5geso9oI23
LVkTbLfjxEphL5DNGVm2aDDShF9jJ7hO1Pvf2mbxD6dGRgdGYcHp/LkYWBr1gC1A
spyTP0BZB+TZLbh3HFTU7Bc8mdtrNlWHdP9k8N+O1/74EFWXe2io6L4gEGP8L7qU
OGw/KXitvivk7qS1c6HzTgZHrZBVxWGTEkwRPP/ipTJeNRRlCA3uJvPdun60moHy
ZPc2tDszl4+sVEz889o6vzBwQ23iy7qOqKd15n5KAdg88nyIY3UWsuBPwP5/TkQN
AzcNDRElwHyIQISkUQq/PiB6bpC5i2IBda4kLuKJNr5+PZsZNPm1Cj0hDvKPds75
MWzGcY//Q2LVc60O/7fJ0Ik58nZn5KsoFmEfhPxE2Vc2Ddz4w8CD+TZ1PBz/sozD
DeOBQ9/eYKehBeaYjBOTlNQux0+JOnq3lnnoBTjtI2Iy7ybyrA2ULJ/R8yp8bjiN
gHaEryQhFawE3STbBUOXp0DbGX1B24LZHZ5vry2Lvy9rJKCeQOJnEVBtuE4BiObB
sQ53mRv5BPnLDUlY2l8ERoiWJCDHJqmqHhAiwxa8CX0GdhANrtrJJI6l/OIOaU1N
UJyP4PumSTLmEJu6Q6xkBndpWSdo60CwfL+bNjuIBP2K7yPh8PjpUP/kP41k5Zxn
dVz1CoR5HJvFNrXC9KwdQwNGHOfV7L0osYr8No4aYxLaAkLiOpgJQ854xR0ig/Su
DQC9qhxlSEOFelxj+PTW3YHno+7gfTLDxOJ8c9I4O0t9rSizqi9d77XC2aqWzM2U
n5dMYdjYfgWOwtyxOkK5eLSH6Qf+EOxcuBKTuivKKJW+Iygyvs4qcjbGRPV3pQf8
loP59QyR4Przqe/vwad1ipE8mpNxFLeogc88V0hAXM75v87DJ3h8JOnR5FxSZO6z
eeTZj3bnZpcsBTbLISQztAvjd01L/ADlDCSPkwRpx/am9RZ47xqOpmKnebKeo/yI
RVzSe+4xDjE//48HxEpiBIzdyLvDFzkihRXkSC6cbiOhqMtcbz1HnmF8rXmkNSis
LgXyJxT83jvNA6co+iCPLrHIOCJMnfbm5MKFQk0Zp8Xljr77hj/yIgHHpQVFX7mr
G3SwKpSUg5A3gFq9PO022FNbEoqsLvI6YNLJ6tFwBKNoTW7hxVylsSvZNed0AmKm
uNOphyt/G3blA3aj10Hk5KmGLo6LOpbEQh5Zgxa6/wROiyZ7KDhYVoMXuOpaddes
if6WD7oNkYaITu4QGLRF0vKCFTUep6bI76Ul0Hu3ldqecn4sCHtZNjm8iaF3F5yc
ZN3vucYhGitCnd8n4x17Loy+HuLdClXCGIAcnN8fe3lFkom+OCjH7hmemMZ1j25U
CPrMs73e229Y32vmm4OkbJWImjneKySnKke8jifdMEL6RhtrG64r2YjjQd99rYme
OysCgT+9HlkLr4ucZg1HYFK4HwX9zkPqhAU56PjYrhanzvWPjyIvXAgEyQh7qsZH
5z70j7HsIfCbXDgcmwDgFVYRYMiiv4V/8ey+wsMy+OvfqfRmu4kqc4EFIhqO+bxb
7jISSsW/cPoeCKh8XGP7fq3I/ylq8blQc0Rez6NZ4s+ka2fIzMOyZg2oWDhkbKxq
zhVwFcnTeFKuaA3s400g2FB5Jj2YWwBfVvTqBb78MFtRE5cH71rnCvKSzScOYjqq
nMuA+Ak0EDqpvHYY7VK70N5KNo9sViwib37PpbvzjlPC+1KEzzYvcTlBgHBm8nzB
kRs14B6txE+Jj0SRYaCj8n2si8JATSz9IzLObo61FIe3a4rCdk/47Eb9MZO+lHzw
lYTM0U0+D9Zvh5+cW1pHMK78D6BwK9Rbj1QO0AxETjkpQHcD/qxcvoBTBG3HwNq4
xI5gVAsGhGOF8V9ArB7+7p6MmJmvpBgM5q9Wold604LYUq753Y3XK1niXrnmgZkW
wbLbqjKs46AftZkSFT9oN8566H53G4SjzgLo7M3xO7EjqUuCAXpQZiVLSnmhKf7I
AtpTsrusTq8ZW1QBzv3SaRhvvOf5Us7oYje+rJD0Nn1FGvliveV8T7WjWfsI5tAS
JGCAmSk6owjIuZgNZ5wUVZE1mZkIXQZNoo5n2AkFfwIcFEGhg0b17eqgLQEXAWXB
SUsOLeavFHwjvxL/ZNeWZ8KB24z9fJSIkeoc/CiGbTb1qE9o2HcwB+L5gGWRUKz7
IPMnE/xQTTKkq+1aXomaGosZnUez6X5jB72Ar0yAu61HGkJ1ZoIFCl9nDXpjN7sP
yYOlS5BoY3f+DcK7IQVM9h+bv/SUFxRjF0CjtedzuInufcqWjdh/46SSbygo+mJR
be9492PLMApJwP/JgDBKf8Wnwwx+06u4Xn2aLS3/t9sHBu+Zlkjy4qqruIr/90FG
SP89vjCONUjJtFQUVh5d4AuT/x0+LQTGJ1JhP3ilzlLOkr4cOzgliB4mjs0Hdip8
EGovXwDRPOx0f6to7DRmkgi4VZPkO9Bait2wEIrxdCY6/yGlpDq5WcwT0mVSuQez
M++6jTv3hEYBISJhezsIQ8dGNs+zlREvfhzfIXwQapSZDNBqrtOS1bv6wOYZevMQ
RQrLhTdJHD68GuCiMXh302muf0FAWZjXEaYxWRbzW34trVc0rxZqQft+y6cJIK3O
crB46RLiHpm2/aWW/TAFZFQAkQQAHwjhRLHZWHdRxTxq3nO6nxWdEWjxvGOkIxHd
Mn32+In5xvfBnIf3FPHKKRmSLHce568TDglFp60dG8o6W1V/PJQEEs/C+noz1zDk
0nlfxwz3uLW4dlnevuD2kH7CRnmiY8Ui5zGrgiYM5D+QplS7bUWpgXRDXUcdDaku
VL5/veDQBLXyGRFUN/eKLn/fYpK8MJkJvnjx2UY+cHs+C1WisZL9hN2uEi/gc6c5
xC4TOxrdI42dJ/E38Xj0mg5/w+kaHRFwP/Zu46iHmWariBqqkmQxL+Cp7WyRg4Cn
fN9q71lVYKDodoKITwjYgjZN0d7Jt6ghYcMu2KjhlGRROBkExQ93j+k0ZnW/C9X/
oJB4swOD5/nf2y590fEHnR77dwEC3UxXx37kqo28qFIhBGKvhAZfdqK+TlV4FEhY
ZAC5Uwe8eWfdM4ydpgwQe1sK/EDeUpXeeBin9/Z+hMKVPCijUXbI8eyOblD8dw5s
R6g3leBFmWKykIYs3kvIRCpmv2uF2Ezd5/dLODRfGGKUIpd6/L6cifH13HCF10MB
6XWbTxlZrdIDpqnMrR1TFtjZBLYcdrRbM4aKn6n00Q5NFyqmFMCsV1m1metH9a07
BI95j69qGjlqGh3m1XdEMb8CEpHa7dKKwjPH6qIMxYGNOBzY2dAmPP58SUaZL8m7
xkDRHNljv96CF8r64z6BOmT22KtcW4o0ocK3Swwkrq8ObRLgTg6hCrzu4b4Lzxlr
vdj1CD9oy1tJHjfQTbhDS5YT1sisL23HKs5zpNUASQ+SkRvn4Zg8k1zJaYyuge8D
2eoGWhqudUX+rLdJR7CuktR/cHLXkm1EtFyvAcBDzImB3HASIYuM/n9ANFndzFPv
k7odfYNeLXNREOEKmTCblL2s4YthFYYBxR2np1IUs9M79i9opTvWwX7hPjaTLyKe
gmolOI2AOPPHKPcnkdPZWIcX7V26/7s0PWdxEqWUJv0AH1M96E564acn5oUEu6t3
HBNlpoax8VTNi2+dmUjizy+566lrrMxPWXIK85fIk9SvFs2zWmXj0lknVs6TmcON
2IgijBrLtV/MQyWn9l2qor/pftnLdD13PxHNr0VdFV4Dhr48pYApRYibNXT/+Yig
raJfSvSH8D5+EoOqmCJEKdE09jdrDUMb+Vhi7tnT4QVJZs8p+vXEn4VoMlH1VGFB
zQnTWFXu2lK586HzEv/DDILDYPRY3ENkPiV9jblvzWxmvTKmd7YlVwnCFhlFMLG/
sS9ktPhZ5Uqb1KZnpAYvjqk62ZfOO1g72YdRxkXLyKsAnNw3tCOaxA+Q+gpRHR4d
Yr8kSBci7YIFGlf385kUA1MM3+/x0EhNT/0LuRgoIz8hLMpIhbAjtuAIGnfyY/6u
RYdo+WKFsRkGiFnYhxhy9gW+q1eDk1Yv9dD8Iwf9nsRBNKP13+6ajYFYDd+4BqXy
nyqU5JrYfJjWmYO4ZdOEUjAAIWBggwAmycWInvyqxuCnTSKpUwtWZCBAu9wmM3UJ
gTxir5RPyAsr3MmOJf+F/FG8mZP/LICggpg2vkEQXdpEnZQicTXWvm3gE+R3VtFr
W/F1z91V0eELlMP40MfEQJ8pREFAo0OkWVuFPgfgyfmI+25/+sc4xT2/fTKG4DJT
szVhJ+CPYnjsE0XBSHlNe1vWzcpJkphaXG3KwWELHCtiFT3FCRC7cxu5RHynolFl
/zJ/5IwjA78yTEUmuRtr0E80Gsdjlx7vhkbCoUDP5hFvOBBsjaUIRcP2/60KMIdC
RaNJI5g9WpZ0TjI+d8AhdbGrkvEcIqGTi7H78/TBg5TQRTnENENdxGZNvgcYEVjD
VBDBJAQS4IcKHvDD+z+IZ1Zz0t5AxPcZNwLkD1Dy3HGxuZzbTZWUKxaorEC8MNso
5zrzE+rrGKlKFeDeTAw5q8gY0TwvGVjYVtEtdgom6in5oPOsJ4G5q3FoOnjq1G8D
394sjl5+vrDrtGVQIPhXWQmGMC0e/OsaU7hLzjg06gZ38MkJp7ed+0xTtcjdvbW3
nD8deKGRRlc61EpUSu3vwA+HoXNdZ4RZ0mJWyDUVBgahQZTWjvSS3M6szkc7OHjo
w4CYW1lRjO7QGhuoTYwtWmrWj7hLhiqr1lIexqgl8Z5B4lq6LGLdQOO66fwnvsbZ
vNLt9TJ2+fxmOpmm4A36TWFVFjRPQquxaTy9bqfPsqhyrcEeY/CBVF5o+NAQlSKa
mYYlDtBSlJy0imYro8ETYPkLf6gO7KwFwwlrAjjUtdksG+mvu9dVNWoRzxP5HqvY
HjCt03jrwlGtCwGsM/3brWMF0JlydCwsmlKJZnwCyjNj5FXwTC7mcCCYwRu1kLt/
3L0LiLci6h8pOLYpgl16cBT71rIdKfPCc+n4O2biArtXsj5uGHjHQZEQzRUVe9mq
/h9NpjKZ4PwgRSYV/+sK0+axSHgDe8a/Srpz9zTZqactMIJXTeC+SUpMMYhIsSRy
1xnv58vl0LBrgHeUCRaerdNVRFbmosPrH2bGmpf1Mgedmtfc/u/nRaYW/NgDGXyv
/CY7ghm3DIfacV7IE1BrQtszlSUrm3mCRaanDX+/ITCY6IomDa/QH+cZkBaYZiLo
dhb7zAhrSBpetylXwI44DmKH6Y8zRnCL1YHo/C8wTRuUN3c8cm3/Beem75Zi11x/
e1tNdjhAwB0TJvk2gF47XPZJOkHKykfI+6GTwqcm0eikq4ERHWXMT9J8sQ8yBkhx
kqQW+e1bFvME40edi+qvvTI/YHNGSyuG+ICVOnIaKjRqpIaAaOCIJrkSJCeufpM/
byJ5cAFx3Nv0LZl1wGbhnbzMinCdS8jIJxSqvytTF/mHabEvcuAXnX89tErYe48Y
OOditwkjluRht2pnuGKKUS5TdwbUq1uNxMYToffv/Qkk4Yf46zuyNSXE31z86s4x
L5jpXRoaDOUw3G1Igz12Dl7Nius2ubgpn+CJxDP0rFV0f+plzNPn3UxdewSkF3f8
fbMdmgAGmp5YMtt7DFHcejpQe6IvVQNE+hh3jzl/61gkuFAa9LIyAhN0mMY9By26
oxTtM0X2/ijFZLfU7yVgj5zTvETwyJkipr8pcAHFe6mrYR/AF3FXVpC9duyPWoPe
eedOE0Vjp12m4ORzqwQE1LbyaIlcRlXwwkmGfrKp99EbBjDya1lZ63sBv8wZt8D9
PtGX+K6HnxO16jbi6x1BBIEqPbZGr3x6J63wNUlkl3LKK3s9oItzXh4KbaJexyBN
9xSNSK4wMRIlPD7LjoUhr9DbuFISB/idYkAeOjDgPg/fqPetYYuIYtMma26v4Gv/
bPl6ANI15CpBAeidKfMP7dVVwCJnvKfbLPdrLQ34caNAkg+cCsu4Jpu+Ej8dfvb9
Ynr4f++j8GsGVrogg7OruUc9n/0iMoIt1AMVxgSjltu3EWRjBwSIMW60QEKoW4zD
MfYJs92aEMB/vsV6p9n4/uAqQM9tjvdiHDF4l2/BGCE+/JrT0ANuTR7Hq9Aq5MP/
AFETuk9CW3A7SZWwm1BTq/77TX8ve1sP2gmovWLCQgL0/3GWcX5B5TKgdGC3ql/R
vbbhb9EgWKNg8rYW5rjx0qK1ATrIz0ImxDLrJQ68NGnH4akYD1q7/i5wLXLp6+dp
jjelV3m1dQk8oQP5LmRiFflIs71yiRfqt7eT8MrjJgJoSliVrd2R0Ixn+qaftvyT
CDL3qloQr7ODteEwIBVTZb35Y2Sg1VeEyJpKaTPdLCckTYk/TALwTi/Aa6wjpItw
UZmyj4Gp/iACj/s88JkSKzvHfc8l4+Ul3BEH2aq9Au4pBCOOOQgAcm70PiSAMM/X
elP3yv3U8oyYGDEHxVvVdAlH5I431DHgeAt/NabXwwEpTyYwaSSFywdJM4Uds6fe
s+WJYsa7XraYyqfiYqzO6ftH2aFnW0tsaXGtRQu/OMC+oqtaiuTYkPNz5FpSBanA
gCKjLfXSihKhismyAqaN/5ChqxuN5OAvOzFoE73PVQNa3+yngfZPZaz5IurRB7xe
lHEzs2xd9GgK5XL53U4NUkIVzB3K+jrcXo3jYrLCG2cl+KMrwF6xtrTzqIc82Do4
xiAXpTIvTsRVpvAkLcPNXSY4JYnpc3OLR+ufpGeC501Pl7s83Bp9qqf4w7NFVLvd
EH/cb7cDXQWAtYFyHNr3jrphY5VHhRKpLjwkqf+LmP/Dsgwl/L81SmK+sZQwi++a
2767px7gxLGIeNO9YqSrRYAND+ogK6hkz8RbsNwNJD7C9CCc7BTxqHEyZq6Ha/aB
hnVG5auLQGz6lqMoh9bceQwSMR7TvYfAhq3FoqGxRx2tkq37JTDUH9esJhi1zObr
4SOrKdMVKpEWMyhSYxO5iAYAcqNmlk2foenUDLI0qcRbiBk0q9sP6pH0l6kgprMw
Evi4KGnCOsS6ituMqPXuyh9h1nrGpV/6R/d330Otr1KNgRljXFQQv5nkhgu4PXqt
SudG+p0EE93YaKKKSgsI6ONUQxUu9EGsZuCMU/C/LgsWmfj5wWgQmiRzNDAuFzlJ
zgteJCBGRXf5/QoU35Tc1F/TREg/DG+gIMyNw4Vmec7aCLCB2g5nbYrNMztlFfl8
fOXYn/GsUYZzoiPUfO8+lfmKrOJrLcehbfsGa+y2q+At6NaLG+cBe0Sf/4le77L9
7xSTxYrOAJuSL+5sZT/wn4hORQUs7hbI6+j1M9dGU0u1BgM6iQRK3wJs7StSlFkA
QZ1Z436z6SbFHZ6LRgcWPgcfh7ViHqVkVNekH1Dz/bUKqtVl6vumKDA9tvEF36C2
+p6Vp7ZUwEQk6aUPBwIarLzL+u31d6aRr8izB/0HOycISwSRTa9RwErRyp/MSBa+
+WELSswqIl07I3cob2wO5GDFCYQysmO3UR5o8QbJl41L6V5ln5muOCH9wsD86ZNd
On76zDZTwhEHnJ9UhTXfnHIKRdQ0rTh6DZxj1Ji+SWEOSCe9gAj2B+jOALcQLC3J
lgasLcJApkLv+qEj9SghkmqXTOWEuvmzd4HKEVQ4yk9qvka8H5OYUrwhoxjrmuqX
ksaMCxT499jivabKKzuKYz67vdEaDUAiTKaO+JjWFIdED97doidTVj/rJbir6ptv
G6FWMZyBqUOmCa+xV21trwLo2GjPliwymlWQjXu66w1FfwLVuNHXKlWypF2ct2XH
JVG257FL9d51NCDYnT6TktCxbtNCkU10CU4EY7TcfqCAFQEYBASlwGN9lDrXdIZ4
swUjw792jkPB+XSmoYzLokHvHHXDOJSOrEkbn7r++HGIFOylKE25IUMMfbmjac2Q
qv64+VWHtaIEI+GI0kcpYw+Xf23Ce/K5zpCLG7tvoE0ZHn00f6wsmzUbKzyR8U7V
hgGNEL+zXT2bx7+YHs51YoOxoSr5ZY6t4Ww0kickrM7g/2Wm2hqBHDe1IHEItynG
7V6vd35NJ9J1aiuMcXIpP8rQs2UrsIvd/fTnHeSaVYtqWHI3oiVmmh9Tdg0NPGFi
V/CUSEDINxd91jRhGmNzfkcBL2/ZPhHwmRtjoSi1lv1kK4X6TkHXqN6Bsw+b6PDb
lyh8OFQw7KNHLGv8nG9S4+SkjT4M5j4aqAkznJ4I4titgtKUJoSMogquzsqPqGpf
7PBK/TbxxOSuAGwobZDm6aJgxLcSdNQ5vbE4VYi5cMlf05gj6Ua7ChDCi5ClXTNW
Pn4LD5jU9Ni49bbnJA5q71bi9SYFYjN4PlUvKPEDhA6mZPOiPu+7+wG2ywAF+tjv
TTzM/y8IVGxO8qyyIv9CTDgfO8MNOcYP4BUNCv6OS5xgXIAlnntX1Sa6qn+lg/Ta
tS9yB85aqDTVE/0dylz/CslZXY2uHe1JMjCeMyRb3poComC1dkTQS6QXNDBuApDG
PUhhvFtTq3jrEDO8hE+eIp6yEziZ2KRP6AEUcGXfW20Xy+SKwxn8QdBafTmSzzQ9
Gkxk1v1gC5CCkNHAH/f5vwwAIafMlxM6EW64bW4q/ll51w+Tyk90wwcBZE+0YM4Q
HUYp/psLHJD+FMIgCHtUKrwuqmmxcrzvCvh1zAoLErOzeeTiD3Vo8vd2r3zkISVv
P5rw7FInvsnRTDMibA4jy+bsFoLz+1OsQa/2LmbrysnQ9tjTKSGf6Q41Fbn+lmRD
8/AIBOPIcoXziDvhW+HeawkgWgAcYSK6suOY1WxPlgb6mlpTRAxdx6OTX5GRs0Ew
AjU5EwjKbaxgF90Mql0k9O5De9+/gTqVErTtmxg07Cc906xQBNXTqeBn31nQwlrC
PMnr/FsYwgzUwTJQew16qYqiGvOi1UUVYJ2AE9CG1Da8DR5UM27q3j/YSY0icbyG
jsxTfBtWF1+GD8oa0GzyvtDjec8drej6A3e9Bw326FMz2mIjpQ7Wr/lLDmmJfn3i
gwy0gHFJDSJw2Y+ueiG4hm9hcmgRoTZwlKOmM+jxJZ2NqPnqj9t7Xq2IavNBEZCx
TtgdBf7vUcchOeCJfSplcDEoGiCZFajQ0PslxM/JZWbef0HLpZ83orwcnFl1w2qT
+dVKeM9E+fnRNwDEFL4ZTYIpuGIOJpZa0SOwZkxZwGsobxGocNlcdWkMS86NPpl1
06paDXE+IZ+MVSK71pYFeVVOf/sFy1OMrDQP/YAKz0UycfCwrFBYg5813C/48utm
7WdmbPmhlMpjipgSG9h8woB7FMWr7y8EP+g7iRqlUZyAJuGKOI7Bv8grXw7sJUwp
ji4DrPOVa2RzQPAtJP3zwc6Ulk+0O8wLOdKOooS7WxDzuoUuHWodmUz76wtfaoS+
szxqaM1hinbyaJwxwpvtqzWwiUoBNG5aoOeOGKTP+ujrqxQ+XUqaPDHKH4F5uP5L
ETBuaiD6QAqjcSmd0vJ8YH5Q3ytS1QxMzfpt48qo2O3O1CGJZt1ObiAQUD8clhTl
tvk5dwkGMGx6hBFKjuUrxGEk07nAeClATqVwBp6xMc2uyKLRB+3UNVzXYhUrRdJJ
kqM5fzhs85xOFmGrUANOUWBWbg/djsPB2oIZEjbDxfHWqvDoVPo+L71FIuhxiUbu
bMx+h/nchufSyp+NwnqL8Kf9aulfwivqJdFF7DCCaAABjbenQTf5kcJxzSLzOFof
9ZM9jSikZ3JKNzrTZf9nX1l34D7ZJ+tRlWl9rm45iUELUiHVNeopdsWDij24rfG8
2P2bfJYayj7M1zS0HPmUkK3w7OSfcvZBVfCpV6YQ/duFqKZ2GD7/s0nVNovMgBAU
cfJq3g0PB7vYM44GnDAvjvaPdwynkK+BfAcigYfZbaaOj4gibKDHoZTxVd1MDUtU
ZlBwUemrZqyA8kKBk/Laop7Mbs3jpfjcW3YFhh7LBE17zyE38dPd4FrTiGwwVNVY
bOH+h05Kt+4Y98C3+M0XAB8aIZHkwz5qOPdt9rn7qchEGYZSJTQhRsDYfb6QmEH2
nTNnZo3EvPYPUUNfuQgYzY+BKj2q85S1vnG1354Ng12spj4TeUwfBZvaWT5jR2Gs
yekTV5mod4cADm48FVU5zOtfWYECHZ5EpT27W9mnmnZAq3IbT8DX5Iapl4aJ13EM
7Puv/Y9UEcwOhQmZAgMqkOPHxRLx4SeJRMmYOsULRc1aQvIDjMpTMFpbOquRvJGf
dS/U8KtcqBYVjYz+aGVWKYGT2dh+BLVZ6dMupXM6qksFHxcrLMuJCMvSwFyVPakF
eOSkILZV+dpxbvRbU6fjvirzYS1NxYWuLER4zYrLPqzT2yGTUGjiL+9QFsZZ3gMd
zSvir3oqN8idoAmpGzvYOZ2FY4FRV0/YCYNPmrjGkdrPfdVcFVMYWvy8V8nAR8a0
AXuRTf0N8a7wcyeZKe+XdFBRgExNDHySOKwYnqn6JFNfvd8xNBZ8fBpgJ5RWUnJb
veq7CCuY2ajZd9XkMwOEi9x6CnnLc23o6k/YQheMLy0uP5vmNlHh+PydcMvggF0l
026c3RsO4phopF/QFI1bnhfVmIIrkcny7jY4smSzu3yk146D3//8Jwa69HZhaZcp
SE0Ky1e81bzSDp2ms+Dh7O/EF8qU5EizGO0oq+vGrL+xUkmBBEEb/Z90hbifLINM
YoM68QicUOn+fJcJuhNkRdSS6kgHZqmL3ZaGC+cnsWRxPbSC6v55midqBoVgAM01
NWug8dSaZ8MjBjqnVaTAJSte9qLJXpIMsEnLM6sEbrr58H4FX5hIumpCWOAQ/qbN
Z63Zu0GdKrXXY4sE0Xg23ShmMVfi931qajajYpuDBdVSokjuCVeKxiAZeq8Kjf1a
SSbiG3bgEKVFtNuPR1mDK0qEwqMzA30VZP+caEe6RM9wgUHg//lfgs+sgkGmqcEy
yPKUr+x/W1qo49j9KvawYtU25dJHj3joW+DOqDryOX/vnLSQZuvrlQDqDC4Lln/L
+Uf11Y3BI7IMddQ4Hj3SOKNI7CVCp4KgXqjI6O/SmM1alu5pWNP/9Bisc6ShUMOd
s3kOkVT808q9HaY8AIkI9Zb1gyyq7n3CiD//vk8iX9S9Gzxn4XITPE+bF0G+Ynv4
mKrwxtN6+ME0EQ7ulEkEXb0J0LCa2pa4CCsYw692fZ2FjupAkfaeVE1dEmax6/Vl
8gDE/zwzGY0eBgHZAaqx5DQDldI/ulALJI5FAXomTYE+KBoC9W3rF+cFK/UWNTnq
KDRpOwQ7+qriROQP3KurryWTUuYG+rFk6ExrHS8PydTpKNWAC/dabyslx3WC/Hi0
ToXmlf46oolWdiesi3/W66iT2eS4dHNZSySoD8OWPB4ialtkqA+cu9B0VQcgzegg
VVFz0xwEnaqLd/omR9VwA09UA0e1au+ocRWGTe7X9QYz+Qfgdz52IBZgWkSJgQwx
KG165bs4mZDgzgo5Ekqj+bW1faMtt4/e0mwROlvQA6NU4owCuqrKSVH2/CVtnDn/
ZmSgd0ARrIBoG4px5BcE6wRScAyzuUW0CFumLdHDU/3zOUwz9AP5yYQZcqUTUzTC
/X0COKcCB3+eZIKClpnYJmyUdtolK+WOwjbIA3+nZJYb6KECa8OHOBC2FnSsa5an
JecZNGW0oRGQIwF34wZ7i6cFf375Orjh7G00eyie3Fo8NzvdP3YQ3rpqulhNS0wn
Q5F84m/WRsQvf7GW/LVBvxTFwzzozgXnq5vo3XJAIxqQW315/A6ujIM9IEzuieW+
wrbmn2D6Nr8TEhRhnbYsf2CwW3Gvfn7x/qfKYN8BxYK7aUzeENC5kQblb1NmNL4A
k7mACMftXBgud0zAN/DetflRf61XRCcC9B7oEMKxF2KqvoX8bt02+Gr/Qj/m5r7D
JYBBOkHDYdixLz1huONBfZsW/9E7Q4z38pNVmXQdlodw1Ajy2/86IEp8Cs0yXuCO
/eVXQI20XCWLpXrEghtkums7Nm0rYkoSUkqu4RpjRB/4O4Kah6RRnLvX60I1pHUO
uRgABULVOfCK147sghslHHKVd4MzAwByGgQTsPf4E1CAx7pcLvD5YxkHw6T2fJpN
hVECjm1I4iI5tJMuJ7fO7AlbA1Y+IGnAgTKa52fHVxTCf6jvuVltc85yFGDqSFUy
V71rOn1myfjt9mSlnOk/CSC3xvTTsWobnaH+n9zBNFaCQ16xYtkQCI1aV+1nvexE
vDWf5cyLu3efXBYTL6xd8KPFd3OaCJXqEM3im+iLB83AObQuGQn+ErTXO7SJANgg
pWOIbxaU8P8UMY3HHp/yjRiuQGis5hK1UqpJVWrf+oiraVe24iiQxAxsv5aP+MpH
mqubZpGy9P8IwitMZD+DGer0X/F0jJuZfwfQanVYh0P75bV020bZ9ejKFoP4abvd
X0bu4nEYykAuONj1TCZSCkIT4TwZJX73RjGK77aomN3k4W0qf6yjv8sKRkYR2Zj8
1NNUqGaELcK9ql0Iur8YjrDq02063XeocmEpnYpvlsQ72eGetub+Lv/LxUhSiCtC
YfE6z32n2sUiwRy1T/7yGFbMdIRKaQ9kSAtUqWNPewZK/foxgXiv+RATDgzlMSvv
0XZ47S1HHPbl0qgjR2AuS/4r7mt2GoIT/Ugi0LxbQOJv6EeOtgf3H7n6i8dmThkn
WGu/ORbMSUfpU6h5behAgsBTU+thibBoXjUxfuYe60TomaOmON8qgLjAdDGy5dPl
fG5a9qYJ603DBpZX3lorwRngCdQKPa6S/mT+L58/kJ5ZwDh2yVs8jFtpgueeHen1
eEGsJrxXcDY0V9BQmU/a18SUyGxTeDLsE6+fhOpA3GMQtl/Pe1LwiUSozyYp6wP/
E1rX7DNvTiSboX/cqCWfztk3dW9QXESz7S0FsU5127O3jecx/1qk92la/Zp/n9AW
ZCaFcrHPGPCnUd5FRliBeFEh/bMrJrVhZQbTKL8Jby87sS0RxbK8C6KrkTw4/RS1
m/7vUfAtCfKyNNpPW4sinQo8R6dokGxbJ1fJtR/evaGxlZVJ/Tw4tqaNhzLASHVY
VsIWaitg6Rf15ucCehBFp3ehC178gej8I29KI5W7mW5SX67lcBe0ipvlrbHGOfWp
96BKATOHVNfymkCQLY5Tl+gtWQxxyxnPO0YIngRky8YoGNGD9i6690xQUVqOrx5F
MDCCyt6HydJ3wcB+6BG+2vuojCfkW+GWxMea91UMGuzz78cpuxXlT/IkDZuxxVFE
X0hNgmxq1YNhIyBfqUSVJAiQqLQjayvVHbfJMerhs1SXLgB/omEdbyr8DrNMxB9V
41T61NQLPowTbWR4ICyTU8+n3bXmKn6baMz6mvfeQlYJeGu4hckNEGC9iS8Ly+hx
QKNmnjRpQ1zFxUaUrEleHnD3OdWtUcWcz+mFO1BQu3xL7G9kIzOXpC55mWdD76hE
DLW4wbrcCf1YXn1Sn3rLJtfQL37CWsFTtBWosiL/DfkdlnpsBlkUoJe6r9i9m3LL
1kiLwUtvjkRD7XwLFH8DvmCLQOALDcPslqwq5+jiTg9/5cRi+bSGEKsrTTl6kNBP
h58KBPzEanwg/th8OXEfFiwZyvo+X174FP6TAzIfUAr4XB5uDYwZ4MGTGnshNTzH
vT68OmWBaFGc82oPKv46w8wiARpeeGlhUHfiIcWSooXXCCms31X41dM+68VF4EYp
cp6fLFiVmAnY8CDUVC9xreIS/oC5980iRnOV2tQciEeyMNiRaJYvyG75wlUq/TPx
fI92cWY79TZPgTd1l+kx4dugHkBe9Xo5kILJpmE/LKbKwOxAJKwd0P6/GTnsT8Hh
oeS2Dcu0c+YEgoktsd4VhZoKJzLAYuvIuSf2xf1KhHT9zSinSK/5RgANbvJ26dq+
mZGBmO6m+uga5zZzwNrxf4J5i1neuj4/rADq6W1FfLlkfKxiXVmp1sGAUdNU4mIX
2kMxwTOA868r4wf5cFyNtmk/dIwJqd8gVQST+i+QnE7pixeUFgkrn1bDUoE+1zBx
GoOpPgpV+s/mMiKjwV5m2x6Cry2bjoBq7CCz8MzLmbOLXAWNzf5BXufjzvDxcnAi
GcEKUVIg9SUIViPQ7YEV7gHbSsZaOtUeoNo1BGgPUd3er+89O0/uIRq67eB0ejZr
goi1cHk4hWsjERXQ8JobaVPUcSeDIDD73KqYWfrJXNU4die6wn0NygmwWpB/UeRp
YbIey6gk/IOQ7E5/IlQsh14F9LB46srSDTsVbW1X+mDw6qxMu1yMhae5YVWC+ARO
njQZl84c0IpmopeyVn5O+UV4NLIoQ9da4pz+8SNw5CBj2dn46gRro93ejGcJtjGp
NsnS1nz0UZG04+LsM/jciTi+WLeLyocBX8mBMyL1b4oJjeFXbusrHe3FHUkpq6Ut
j6+Q1WJK1U+IU00pWpMUDp1Q1E3W22kNasNUAL1/FZPWqWTsi9pmc4+ETa+rOoYa
I+xpZwHHIlS9OiW7e7l2JZnCcpVlJU/1JekqxqDKy4PyvrkBAoNGJJ0VsWuosqNh
r5O0JlMmXtZ25P73df3OegDy/Zqt53qkqhCWDrn3yFxaBQnSygIRiWmvOJFkj3oS
9QSzXP3+F6WDd8Gh+ot3AgrSJxYnw4VXk3CRSdmriBIKgDoSUYSnwVLQMKZ+DI/Q
5lzP30Y+/KbbF4Tu36qxsvuOYgBO/tOif9+Y+4U+jGEzVjnzmt7z4QdXD4fIF29I
7wAWt/rPbqNvlzi9PiheSXRRM+nfZrkBxkY5pTyjfqmzL+8XlJAsCTKG5KaDA08G
xbXlSz6cvysHxKnY30idaatQFm+5X9XIAJmJI3uxRWxmmGy0dNt8Ue/dSgrhUUEt
3HkQwz3P3uXspE4qnPlL6deKrK0q5G+kVLgInxQpZRY77Ti5IoRVW7zeyf4i4tMt
ycNGMn+UwadKIQPdt70J6RssoQRC12uSSOF8WqIW8iXJYTx3bWPg7BRfOgDqhHjy
oL8msjG4+KDBsZROiNiNGK+yeiylrYpRqGgUuA1d95ar5afw4d+RwQzT9nx8Y+q7
24ngNYHpfRrvygHMgI58nSFMMori/2JNVZqI1Do2/ULlTgISubjGF8O9AcjxOXKP
TLIe1XiLq4SOLMYTiJSBM2ofh3h/0WNtpDQqjapBBiuiEeoWrlCk2t3EMmR2/Zzq
Rzz+UZuzMjS66L1b4w84NN/lKdt5edhpHBlV5E1gUZ7fH5WA9x89669x1ayE6W+K
61Aw66E4zvwq51JZbfzhO9zmQZxCTZYX5OFuNLi70KVD82KB/rJtpYMTdG5hqzzM
0xIphWQXpf/JlU1cn8GbowYZwOSTmc0zXqfgmcbdeVtwFiVZZ/F8rWNtsHkFR5uT
m3v1E5bOTntR+YIOgJFGlC0KyeEo2jV5rBjOSG/dt2x7omM39vVA3ux8iP0wB/U6
DPQPsAi1PRwUTAocB5ZpkHv//QdIePr352bjZRJ8QTuyf/zPugZnlfqS1B0FmMsI
jDB2ykr3J+u97VtGqsOxZvIoZPNTupdmh0Awek6NPYzWo/vy6kKDKG7TBASeX0jX
szVIXqE9YZm3lWIGqzRPOVxBuU6F5fiYU1u3hhb2nCOwR7nM5njrfH9MpTcvy60G
A9UBFuRWyKyUbPtqos6Evk+OGVSWTFM93dWFWjR7iJjT24Vr9HjRoyFdAlX6SECB
bTPd66qYZJ+wlO/qMz0Z31fXlpiL8tCg3hXvqa6MEWliGWw1B1b9/Ht/midpmtTR
geobeDrz+9Nkqrqb/PX23rH6aoAYzSaqOzsO0t4U5ynGuiQv1SymGCFe3CpRHair
wxmHmCkTttSzpPkaZeak2roIiKi38EZTY8znFXzEXgIDH39omlMDRgWzTOAyTuZF
in5d6z/4WXi1vr+2UcQLim6OdvrhNIbstrSDRaIPQMGT0Cb0tDjyTXUas3GiGJBj
8FM3rO/TrKIR2Ue/Rc2lUBSzSb3gN7AOcme9R7WUL3GNavMvm/RRRmxhl2OwreiF
G9T8yjm+J6rvt/mUD72lImxCh9LwQKEDwHFNj8CAWzWbefleqkqaFoO4LBzeFzed
vSzsygvlw0sAuYbba55T+YMFKp0OzfoHgb6CTeHF+bYWRbN9KZTw0k9vw85YguI7
tGRSMhSDTzizJbq9oy31/tVeRpnHZHz21xV0ROWQSE2yxB1fDaPtpRY0Pp3IBSEc
a6HG4aiXNewQRd5QTYc1GqEU/F/nE+frRqRe4FG3YhxABoGVwmmRK/GR9plVynJW
8+p3Mq69qMFuk0hN9gXYn5Lud0/r9PnunDg63UHyLm9+hcCIwYjaJMjmfZyywR1W
Tuhe2oqBnoO6WM39g3tz+RJtZIjP5JneLaADuPXa3QKe/gMTK2uxGV8STOxaFiay
u/CQTf9c+cKZKlLmYNcdrG00u38hHQpNU+q0H9ydtG47Cy9We9AGtKWn8tSnsSAJ
4M3qoKHhSYezuC/h8NWd/YofOCrvSOZ7G7vRFp7RTGplpuH7mMnBoaWmxGfIxunX
i/vSq+gLmErQbD7kgXiyXq/PnxA3KZgo/pa2mwPYzRB6NxeFj67tRbqS6Fj7vZ92
DfrgF8YpPemvote/O3JLWnYXwqm8y20P6BqsMS0vJwqJCUx9/hklZsVpUHwCiM8z
QGoTpmMHc6I7dUxjOkoFWCLB48O4OOy5kMuAdVZhytkDsyPcvmWt0lVx0IwjQrpP
Xl8b+0ifsl/YJKPMWZ8R84IleKNuVxcLLKk0SYSIJgGqVYe4TVrMt8oxxdA+62Mp
2abzBY7ljDPAaydgVYMcXHpwb1Lug9stDGn5OpdRXEZhdT+iA7XdARNB/YjTAsY4
8l+QTKgPrxp52sjVwskiJtuoQ0D86FliU5FMOYpy3eZrlMVAbseXzl51Ci6j9/wU
5Gf1ntsdtJpcRX9Mnh7kyDwDI8VIyK8CqklK1M+I2oC/AMY8H4gtkh6eIkdTO1uC
J6Gcw15/4XWcYKxcht75ivareaZeRVhGtl8DSQbPvjlZ+O4dpXEJtKbQe4bb+cha
loHPy8iJom94D3lcrukP65p5krx3zLBv9LRaTbYvQWu+GAejs2BC1Zzq/No26wgT
+GQDPXB3eE1o6e0M2432rZg8zw5fkDi1wfziMODZDxCz0/X9OMQqUx7c02TP1pIv
Ixjt3j9wCMTOQ2aNnM8WnSdUjkeS5tDNVp4xsQoIqcVn2JJUmU1Ccbz3L1/SacHP
X4KRKltdz7FNtsahpGDvNjLmPp7GRqqYhnuU1cyb5dNqTl4amjNNx/D5NBEioOQM
OFAObMGN2GjijET0mOkvhi9M+sVh8lCp8aJHgLTcytCSP3dME6ud+0gD+a/lI101
GB/wZLUdsaPYuGFr+7pm4O+/WxJ8kUebeQ9cF3eDCAovEmlfiEJettYQuDFH+r3d
eFCoNyR9LwpUHyx5Ia/5xWFVZMSHQN+EAKJlgRusta478kpMCaD6bl/lKnI/67B6
yblpaABoFsLuY3VyrIo1ptYehHNZklt6ENZIRIjt6odh0u2XMQzRZM7pdP2jUKVz
2nz9MouLOhXXLWgSEoydLYOmiEAsWIG04i04vTtamDDaEg/ZOMH6mYaJZM8CYDpp
Ib2rxyXWLF3TeSe0KmFT0DBapTDAWTbtHGDeySHayxDR/EWD1pRf/Uks6Ftx2qXW
CkUGncyvBWKql8Fc0ZHZKzrYDjEixRKJPyZ6KvwvfiDOb5YmeT02GG2IFxPMHiUJ
QK9k1TIPiDE55hHZfyWh7pe5ucXkRO7odCVzSxnL1YY/jfTHlhXVsLaWFlvvHizs
rZqt5VxQJO6VueCBTLLwHxSHIz1p/R5trwpjah/QHasrZoYBW48qSo9VC7UrAS7i
BcpAkscRad9yMB9jDlmFi3IRrZ0XFzk+cLeOr/cRWVj1MiT9OrxlpPpLVLWXoxD9
uRG3uLBtLlhRtAlXYHe8yb3R+M1IrqzebQwuMH2bqUYa/7is4F4GrOKenCG/zKS6
Qrke1QEv4WpBz/PQNX46p5wC4QsTQXkiWUL26LCyrFV1HRv/8tFPn+whY4QILigi
Rfuhq5yjflq2gtahRsZNNI2qSEmCH+RIVhtvCVMEawKqM8wfVFH7K7SksESd/4+I
rDTRLsQ6IT4+R7eWhipF0JzZUA6Srecnrw3KVtNoPAVEhnYsY06qxNywauyk1m/t
bc1vtmfSzLwc+yLpBCcznjW/UWEsquyTB47vljbUApniarakOYvW/8tN6uYN6fCq
cu22gV/OgnyKfwbhmOdv7hvQ75bVbEF8C/1fid2snUWwhsj7t8q029RVwnoraFP0
3Az4Wkz/Xq+gepR9XhMKnry/q71fyzze66zbBaqnFW34dGJ4ZmikUAPpkCaOW7UQ
HhLzl+8nud2U7nYDe24TEGU0cpGPUhguEC1ayuEq4e3TDVPyUzVnxlLGhDiYABBV
Z5ilfEj5azmA4jFfsm8L6KAQAZoVbFe1CbSb11LGhqSTFgHWsKYFwOW9iYPXZqcg
O+VJg6xe8ix6nQI44izLci069i3bNaZs8Q0Pa0jCNjZeFZE0Ngxwtj/6WGLz5u2n
94OVMc7Hp0ipNX+iqjOIhvy3B9x49H5NIDLx6e4Rlwk0p8YfRiWoJmKW2v0trZ1U
O8dfVR3ic5/DEa+p63G13iR3BhSLrQ6RHaN9T1GruNLuGfp/1fCH0n6PDFM1gDbn
rB6Zv9B1kI61zDME3Z2Fhz9B6cXtbKTQJSLTC1wfDeVP/p4QR3u2a6ima8LblGrh
wf6lPylU9VAEaqkNiZV4h0UfmTY6bJSILxDKGYrFapZ6DO3Lhqsgk1qgSZohhkE7
gSufQHAREoEG21DVo5f2/5RDNc0GzzQmqCSUsB6xjhrSPNlwOBdbZhjx3et8AX2s
XFxdgwtfau8rWn0uo3rpdPi+PopyefQTSXbXY05Efp/zCVgqQrx/w+YFXIzVRTgO
VRiFNFpq2QS9/IwgKhrhf0XLAma5sEUwskWlKokwGYC+NbbC2xCKzK8mouHYPKIC
CtbWLz5CNji4Kas1mNmzRVC/d25lxXEAPB7BAyzpy3LvBKK3L7FzHDkldXxLmw+I
9icvkeqbr1wx/tFSpLlWV6E2EBgGaytyvsbu2Kr62OIfxIR6ybcaHnpCQqTyi2pN
d45bIY0HsFqxKItz2SuRkKa8nLdJhxW54cz/hsbzIWJLEwSU5CdNe52JJkcLLk46
+KS9Zh2SrA+RIFb+sBDB5hpVIau0ffgKM2gU/2B1MfjvmgOxS8fLB3vrdBmBtQ72
KUEpgJ4PR6UdszmkyqMsLubpNjbSOgaoqSjFU6g1U7tXT8wnxdfcEIW4szw/kgDQ
glVl6FBOy27lXQHt1wc1FNF/AsAAiEMradgsIST4ggv9mIxVgZPZUGArPJV/IhaZ
n3pJyuQvJJVUEIR1Yw2Gq9/JpEEGMQn1CBeNeKK5cPkcHFLHqdRxKHXfNhmFtI/5
6dLSEz5P1KY5IeyvpPDFWWCCV4IdwU9Z6wNfzIKM5h1UMHNx/40P1klrR7ZLDD8K
ZE2NKpgVhs5lm40MYjfJtIN8gWX7mh8EysjF3xRB2cdyAyIMPTespybrRkR2xe8H
7PccCJEYViRw6nkJVIZRyjJIW9frGOty20b1wqzgcIIfgpAnXsuMWVe3YRGG0jrc
g+4QOgfWvDtSSIILSdQslzEuPUvfkneVvv/usefdie4s4SQ6J6tABcuwyRlTaAlX
TKKQbwcpat76kyxhbBUisTjueYXORpEju/KJvmjeh+kHSzfrAfCquPe9MLZdwM6E
/HqGK3mrg6AkswXwgpXtkYVhL4h6TbRB6tC3/KTwojrk2S1FhFqIcnLZN9t5hefD
Y0j7Sy1Y5mjW4C4i9qcQlkLUAYsxRsJE9fQVZQVtYvG6Ss3qdiiIj9kNa+FrzwUg
Sl79BDMp8yRabhODnMYX/Dns/ZS82xUvCRy8X6WNF54/0oTt64YLmHT+Z2NbQiEP
KojdLrNyrRL0Iz3xU/7AC8VQ32XeOg/+5TIh73ymbp8BksUBO14oGhPsSfaPxLqw
ej+NesDaxLaAZnUpXagcJqgFd//jWrayhROBHtbeFiswAvb3gMX+qFkS1DLa0tTw
+7X7HkWoq8w3bKjakOSiySktadRuBSvXMkOSTcqCcy1/okm/4AounqXkpLhsOwUs
vijmDfTR66YjH8oEwIXDv7zL3rSSWbr9sP3mqeTuGUfm4fivep8CiS7wvhwTQU8c
yakHKaQcUJrIgNSd/mDx7i+HSW+m5OdUtYAep07T5ot7Gv134FsPEbSBdt6yvyf1
kiitXA6b9bWb/jehyHBWwZvKfC+hugDqCwZj7z2hGAgqiMNYuUbYQTqGbBaxIDWZ
f61GCY8ub5MnHTMaLYB/290FtMDpknEV0NTiDasqcLR6vOKOPd90pAFZayT/509h
ySFiSFvCh/Luh4/6y4cMdraCDmn4Hclznz32K/6jjFRC9kg+2T5tQ/nR0JGTuCIB
iWAOhuZh9f2VeHo/X8/e4UGxmgJnnjnYuuxhkTFokK6xdKpDIyGYhaugi7RwHi//
SZhmKr3iDapySMllS1EAKALpM5MUM/DxAj69yZvoJfo27k3fKu1xI5AEqzAfifmD
Vaglq4HGJuog+wtfcOKHQuKofSfqZv0VYEzoA7eEqOxo72T1pGSKjLbb/i2hBXGI
nYyYkiMVZFJmggs6a/GvMYm1agHjV0RDpVeJ2LZp5AHJVeEC8VllPHrvrNF3iKvz
NSPsTMbKWm17hFAaQWG44mpm2XZJEafV+Hj8qU2mLhC+5vOrIkmxiqTJX0HfQSti
1NDmZXKekVR4nlyEnUV2WaXHMFdbvG138OPqgUMzUwYlG1l4jJDj2nstA1smOSwA
zIqnBNsn6Y9h+R/tIuzjxHGWj0/WK88nJEPbnZ3Ju1tqvB/yHPtrFTkoIVkJyEH/
H3ei78E0YyR3tihSE71G8LdCnOGFZMPlgZNn+v4IkeiidFJDG8rSllDJK6YAChFE
hlCMmqTXc0I4nO1ugdgrxlGhB/leXEDygKA82VHCdMpBKlTEwYpEKh9596Bpfzmw
avb7hqRBjwI2R4EYO/Ep+e5Qghx+i87OZiB17trBxYTgUYzhjo71z20Obvfnvr07
RVT8LfJ9kpYonU+OTW4sBSv/eNXe0ixkvg9m5secop0ngmNeqNIfQjpefm+Btf2M
rdyxaLUTAzb4sFGZ+3gP8pytdb/zULWMwGPGNWLcYNPhRwIFAl8UrH/gOrsDGRi/
FiwuRLN5z90zThqmQ5BT3YHyn/fifoSzc0DYcEoSiIzF0mk6a4qzZNVqt4L9UaHN
Ip1hN318YVPp8Bz+gdHJeyn+Iv50+avqB7XEqHQ8rZ50m9He9SYYz5B5LcztakCy
a+fvDd2LE8n2L9EsSaCDRsZdTemfmvkk8T7PCW809ilgXYyws7xNOj6/pbqd3EYI
t7jWIp5ee/rG9lBgnXKxflA9/ju16aB4HRprmouuhyF9Rez5Xshl7+dLscNl2gKZ
rsxhI3f6EdyOSklDHCqTvzW9aAblVQfXXIXi7k9r8EIippQKkkIOdiM0uwWUlke6
UW/l5x0D3eiq1vrOLCHNy8QuHUQU27kL2o3NS1ug2/HfJxUH4CEYA+b9LNy0kqeB
hAsJG/w7UOH2NJxCbJR05KzqcRPptnZGLw7XgSmA7FB7VeHtW9WCkEWhIa2dIa6y
XvOHCPN/gJGsrma3HjENG85yQvttFuSimH25EFEZn5zXS4KGkVf7E4mIO0eHX+Xg
vzxFPvrnBR6Z0+Gq8xBdvQpbe0stVqC5WM/DQvHisLk53AqDdloOcZO6rh7JmYgc
KmdF2SXZQ0LW/pJ+dvSnhEvz84JExTBKNKDbt37nhHKk94oI0nqZf4bEgfx22ovB
j1tKYomULxxrOM3ePEfF7ph800TLaRFWYQjdhffZrh2qoSskDlNVjuaYpYFXqclj
B2tQj7arjW5qeh3KEaF9ON3p4Gd3OAxH0ueAwrvR88CWR5ZM0MsveUrepkY29eRa
/aUY4cceFPTQeFFU8wIs2FdD/z7yR6bUkeGS6qruoDp+XSp0Utssc3mbjBoFWScO
hkEoT+O5/kyq81d/n2zrurd7NqpN2zizrgcBHyQLdCRLGTcFNsNvX+MNBFJtcp9n
rf3WdCMPc14RbJDoJZzQ8Ut12WdxfqeHE8o9KOCiHoHjXqCy4DBzC7JfxjENnTZk
Rvg0WQJrmEp2HxN7+uwZusduZaE5lRb3u7etDhDUpLBxO6HICaNkDUTLbsFG6jL5
w3PK+X8v4Yow4miVOYwZlvUdBZWQA5JwFyWHYe0sVt/IY+LhHSSXy0R8D49qm/+e
bOKE5a0LNVRs2+qC2NW9dMfpeN3dKHo3JMfzQEJM7aClUsLPJgr1JcrhoCa/B5VE
kCIH4HJVfKmXYJzQHJ2Hn3M8V6Jj0XZa1nULkAsNmYlUhl3H0MwThW+c9kFBNWmA
XyxwOb4DvT7i7DUDn2HyFO1/rPUM/7VmhIHLLaZcHGLVkZnk5eryB2J1wmMQYfM+
Rr8DUDtjaNR9zvrKgISBLodJ2b7L9px5xpTfqtU+c1MPmJe4svS1+KVTvat89KeH
Ozj1t2VI0kS49iYLiz/nMejt2QJfGK5OoeOLOJKyS3F//99K1Y3HW/WdMYez9kXN
ABFhvyRhvgGbH3MpHtXkJKxVSOFw6MrualxoOqq2ruYYND98Nvsxy5KFUgN/tbIy
ja/DNh7HgUCB18atqQDq3QBqc3+aWWVWRVUyTQ/XKUyzCJELBGf1e9RyLJV5dKdn
eK41bM/nT2W3u5oZ7XZKzW5meOC9f2bBcFE23qVXjUFfkPZYRCvG7IUfxS2rhCu8
jB/RcnbAZz43rOAG53WorSD1dk8/0llHwDW1f/jirUejEwSig8DqOwp7POxPELv9
oPTtetbbfHA46d6FFnNsZkAQYDntT+ZzUVvu17XdawyqIW0bpbmdbztuNKGwzbHl
JablBT4d8rT8YsCkGnRzvYTWXsAGatyc9Ch37bjUyAJ4ZDSshY4pam1X42ENQoB0
PepQC5PdJdbFRxe1XK9mSBPAkwGYU9jgD5yYIfqFTTddJohGx7n/KusdNqjpxc0J
LurzwSnqT1m9BIG5LfbFFvmTvjznnZ5D8RJBTdPZKCep9hg7HtEazdlrJcc7vQ9u
E9cDa9q96sWPOIJuSUQepV/0civusEXgnK3voXYkBsnn/xwlU39jX9TZXlO5+fwZ
7O299NCyazr+qNhwA56It64zQ2A+uVzFvYd08BB0xcV4p35LIGdVOO7akmWgcHvh
f25wNWEf9+pHTg/Ke03d2Cdmen4KNFvGaP5BkHLq9uy7ySwIFmSHORrhSlOagwEN
NP210P+yTUiUpfzk3uDAS2VbDxqpDOGEE5R0VjEqnltpRX8xKHehul3sGpqtU3Ee
szZpNdBhT/OGX5nVLcf8RboLOn7O0uHhgCh1OGnLyzHNlOeY83UTMgedONeAvMtS
Cx4lrSaOeAEUKWo4gKhcTunL0tJWh28APCiLvp+hXMBQnh/kC16fLBc0NJPrpJTg
Qc7TdbzkqRXhClhUm96It7RA8ecM1XZ/PPn/pLrb/ae1ncaB9Ii7kpZ8BDqr7+8E
21bQhtDSZu45qLzo6qHNPvY3kZTQfyi3uJVcabCHa/O8OnCy5OmUV5xBwTHFJUVS
a+JfGLCt119HQuH5yzMceJcP2zV1ZRnXgCBQIAhZd0GwJ/uZRpSf38wabwaQiwm/
zyxJ8uVN4bAkASOyB/avpza5Zpxz4wJUY2K8WGvfCct4mRkbxfazyk4m0UIS2FET
GtnbQlhBFPmYSN9W3AKEr/Kpmyu6J0Fw6/DVHtv/md4FVdi5NyzPScDl27vegfLq
cIdRBS49JpGsRGkdBpiUmnGxIINSKHp+jiPf7weQ9XIbChsphvKXVAZQfy/f4/C+
4/2BOPPEGC4/H3QucSAMtuZH/43hnD4mnVqWwAh6xXgnfMEaASUh718DqVX+Fvlf
FnXL+blRrHE8ei8CC4W6PZbXcDlvmVAcvuwWgqfR6VxPeqixZUmUtsM6uXBlw4Kp
IksmOvldNIDiEWgZO4fYaK3ie7T4Ga1htFPSIKiJaox6R6H6+XUyTqsHeTSGft9I
cr7a2YBuNHIeU3dpedkQHUjrWSvTI39haKUyTXYlf83zSPr9u3sc9SJN9XITKLjo
JKHrROWJ4CpCNTfuzYOay8ywr35aOIBT8RCxYzRJRL+ADPTQMnyXOdfAdZj7cZS4
2P18EXspP+EFZzKo/gT+W9h+7Vujz9PJIgvxF6sATLUi9kZcBeqTQeVhjhONoqXL
p2GABCCDL/BVa4A3EO6S3hy31AeMZJaZbBjZzcNzPPS6+uC1VOB1VcRzjhODRzlu
RHsWKu5jPEbdgehY8zpeFF5CzLmv4mdl5lMKhixjcRbNLkfFo7PVhfJmsTDO5V0p
VTYDkf8cEJbxSkJvvcGhSibsWRULePcDUXTQ/d0DzKi9xPuR29lK/zDMHWcbkVyL
uwhVtAMjCmPKP6AgucRHIf9ZfJzq4Y9jykXvA4IhE3E3ifM0hy1yXoelM6+p1qf8
Y3h/Ei3xpc8B7yQ8Z3e5xtXPZRbkxyocL6ec+rzklL/1gHDdTUnNb32kX7mnBbl2
IzE8xLYcBCV7nzAFS0JqdDNJ3E77SU8CoVriWm3UbXQ32UOOg8ShO9iV79kPV8Lo
5cV4PhobDHd0iX61rINLawjlCgAWQrM0D711aMEfIUH4lwK16gr93qcyakFqRT3t
1VG54mFtRAD8cmcFFraej6db2AKsafk70yBkBwl3B9GNP1nfcD4POpcgAkMkikN6
Yqb49wi2vGpcdccTjbb8Pe5sXOjEuh/YNox58OEX6cZIhOlCFnbr84CgAGyJpX31
amS0wRNpNvHzRC29oFEo1FLGqUwxRJG8WtBanHKuNo/JBAodqdFcCLN2Yb5pH/d1
f81Bvk1jFnZrkOmJjyEKxdrKQMA6AcgiMJROCphjU2unCOoGSBmLbr666K5Q/cVD
IOZJmsE6MrRj/0mlQyfsrm2xfYVDubkxHOneAvqSonFz3jJd0441bbqI/ZXL6c68
tjDc5P+LUIsc2+qPQ2xjP+tC6j/gskLuCiDrNKSsYDNRq2lVIqPxaEnq6rclDqN1
WKT+iHWhMN2Uxto7f8PC9VYE+9mvh8Sxtc7VKOMF3fHzHVOWQVK3A3UjTSM6dE8n
Ron15nTIMdN5aBFeKnWwTepOaKTV/UDM/mDkdFPNJLDzYHmO10zii49i5wkJy0fu
CSsGmYbOnKjZ2pVoZAtDqQEm4XTLXh976g7RokwJTYkLQHnz9deX9xCWxXD8JH92
uGpTCrtSOHj+eVpXQmUhNbtbWJMRGeBEdD/gxS3fRpuzGzRUn/xjmOC2JV8wvqhN
bHGXkCx7q/9PrnxQ7r/wTWz/thB7+17uYkLQUiUvqfJS8ixqXgQPOU1aO+JBc4z4
LEgr4jvJAW1EJQaDP38ACXlYpQ3/pkZkYKO7HxsqTLatv/5nntYO4oHlMCwI4ESj
XtILD36Tw4pU1c1QWBPJsZwnzemFjVHRE79KHrbu7n3ZoNAej3l87gtgdaDGu+s/
hanfSvkW/6rPOIu/AFwwPTRcG6Mb3TLnPp2yJhT9rOLz5v9LEFUzb07PUhoUY+Hf
OWAN9505T844bNcvmSeQrJNPykVxV10tEW2cBS2fwu9xjOh5hbvX72OZ+N8RLY7j
qY7oUUG8gDFUEIi8bEpbyskZB8kzSb2mfroVJ/LJjTpINpHq0He15hjRbGPpHIs1
93YbOVtg6sFpYFV4/A+KDCc1jhPi3/1a3DE2nd15vZ20ftppDe0YeaGMtOSIEZ5l
9xAVzSBb3Lv03OxGcI4kg9Uv8o3VSIw6iF7AArXCEqx7drGI94U1u1+u9acHXh8C
B2wDYFsrGcK8U0H/SPVaHUD7Kf2uMjW/0Olsi1cn2vLAuFtL5ze79ZStV8aw4MQL
HhekSs5njmBT7HwbZiLrS9KL2KH/21fVDQr+n7sgmLWUOtA9W+irSFN81uIydhQr
CVrNiPKTAQKMrb1IND9wc9RjJu4oSW9O0YGQf7Jk7GDIS20NiorwkQHYXrs/j9hQ
sfNmsrGyR3DrGh7YwzFw4BSUhz9Ub2EDFrRLr9LmVCHU1QYzey6IYpseh8gfcgkE
Jv1aGfEiw3NZJ/FrAEWnTwwCVAShWSI8Y+sMWyWO3ziOOo21nAJ5OJiLqbxg7OG9
5539hG0LAcmj+626ryYVEGhKCVjzh8SkARd62Pi9ogVKl73uM3OvFZnrssmDiZmY
C4yFhW2fNqx2XkNmLNz6yVtAWtLtzq+Bja2Y+LNrozIt1cOc86rAiS/tpvTmNjPm
5V4eZryX4jEHBYPH2oXlKphUrcCZRszg+1BXBvBskAXQzT8IL7uaKm0POOYwv1S/
grY9V+gWNwflAqDHzO+dw3hHHFGu3Sn6vfDcLK4zVO2PDOZknfEzLYXxy3DaxSx5
1ldvIMcbrs98WsDgA5w2AW21JRmPYk017QnsnZriu9EqW72qt3I6vqf+cXGdue1w
Fsz/irviTaL8vCd1J0syXYjyrObw6SnT5vP+XvecrpSg1hZqJ4v3UDMqJ8YXMGZ3
+p21y+CjuUZclAE7xeZwwCaMjg9rXLh9sIwRqwDwbDcspDHKvy+vbU0BmY62yt82
wQxUxt3GooeXaPMGUS8ErmBa6ooAdOH7FUYolbQsTjpGskpzOb6R2wROorB2bVoF
wUxveLs3eOsltNk8VqOun5YOvo/r0thR1XSZtvNkLfcCd1SwcP/fhQGl/bInRMlT
Z2GICxZnODXY1nvhN81199O3VAHD1SDhaGYQZ5XlCyTR6fjf5+PzNEpI8RTIPRa9
teXWWWB0NqffmdpJbVP8UH8gNxzwuNpp7MnOmzlrWjlDc+aTf3ae4/lfeofr/2FN
RK55Se0iKULgs9Eo+TGdyz8CQkg90eJyQWPE/85V3OMvGjO7t59m0Te6cHweg4wM
/rEK8XdeJUNTYwhDiraHcAWFI01a1PN4nYcN33AFjvCm1bBOuH/u+ox1uYkKryFa
mr/lOPxA2/F+DcWtAlnw8FzaPtweFCvQw49RELxiBHCkfNcNcZpjcza6a1zQUIqh
VhVFby45mdFjrRKQstQ0iedTmXQ78dtWEn/VwM2K1svwIJrmeBh4UJjxw4qL3Ix9
808ddah95wQGbPa6qZC/N2Z5CCJfw8QgtdSspSugkAT2CkZbMQyWbPX8vvsy6h3I
hf9lAPH0/Vk9bjjFCnEJhbqnE61JHXXPzfFyv9Hn/J6OUGBzrJ+i3d4SjecSDeN1
SeDSpmn94mPAsh1btWqIXaK/uZ7FLFzylbrgrCboCweHhiD8f0qQI/LFKNYEM6sW
3EZno0rorB6TM0gct0DabCVRu2XyJM5yB+Y9KQzJHEfXSgkiiYARhUodO/WbOKHs
Lv8pPHaJmI+xm6Zi6kE6/iS5ASwaid2ZHSdM+EsPAdTuXEzQFqUQC4AWPDf9tZc+
Bn/OB8YZSbrGMQ/SdXbbZ44ciArpsTIL26aK7qq4ga8z7QDo1ktMd8fNQ4gnR4LH
ChefnWmfNDhuowAgRc20NFL7pQxPEIcRyzSQL1dtIZnr2FpQyAKaJxKFn5Y6MYsI
+SVUP6/WIQjIBGqup7ZpHK0EE30NeWsfekpqkXluLapmobDu0qIPuBkcdUxzp+KM
mnlIb0+PwLEUIKLJUIa1TZCn32EBIe8K6Cm9ZsqkQwjeud+72e7S/63d+z5cfX6o
ldTkbrD0ohD2nHs993p4XZ8OQlfCHCzS9918RhUKVCRKtA9fyL7FS6oOlk6BaMq1
uR6RHSwXEcGU89iY+hqVFmi3t8Aoz3McIeYx4bRddSDtoYIRtggy0Y5n0h0fgKOS
a97SQMbrYgjw5jvhs3MF/tD0IuI+qSqXWg0cVYAkAFMrcBXNxYFl85+qBO7wpB6/
Nxf7F7dYfknJS+DRoZs09mr7+cuHlYYuNXhEoVkn4jjt7N1P+TjhEnLPjF66BM4I
4mS0Tvuj0AcMiCwtFmI84g//YSWCco41F38kBiZfwsSovGiYP/KE/lYeS7F6W2nt
wTwIAnWempWelilQ7A/DG4qm88z53GM9+JaWdl40PeQ0SHnb1afBVOJEZcIZjF6t
/2lHjsYTZIaAIB3gvlRcNhmbd6pCiNYv6GTcsvwNfcKXL+3Q3eIP+g9Lp9G6QSrU
mvNAE+rxXa2rV4X1p3xrCjr0oqzekKX5Gr2aB9qBVk+eo0vp+IMrovSuCinhVz6O
+Flvs4aJ3c30DgrfdOQKE7R2nnGKBHrN80OmULrXjk4BVMia+tZldWmelulZEI/Q
iSFNGVJ/vMUoyC5j1m6e0C8SXZD5D1T7tABJLc3EMxHM1A1vUYrseBvnngnn6RXb
hdT3L+cc83nlfBoaTlHDqBm/KRJ20o1wXEq1ztl6emabqYa/nG6cdSAqOaRuz5Z7
rTGWTqHnE+nh1f4AF4DqMhv3wBxHO0WaXwwmYWKMnFcDmO+xrSnl4EChN94rQiNE
c5V5LTpp4mYKu0FUas67YjYgAg+57l4ti6l1rx/dD9TwIMRrt+su3E8PdjfnlZ+u
2aDp+icSaoZBiADXvtgJLwPfHUCffuVN775NxGCRgQwPIm/YP4ZH50GFt6UcPcJD
HfDg0jNVdi33XAKzv1zs7PtdTuJp1y+spE+guLv9gXOK+DTUY1Vi7G9PQ/vxWmsO
wY6dBDaDMChLJeVHcLWo/Bm8hAte9Yk4Vzsf64F8QMGB1bi7jNuN5gXSPHr21ps8
qZLpihHnIVEMON7ZwiVQ8oB1hOvm+E+9HFFfasbhS/RKF4QYOChMR4FqJ2jlx5SQ
OaNON4AJfKZmnSkovDNrO3af1s2lah+5Szik15wDIvRwkdh7tStOlW4Vnv1/oEfy
iT/qfOYBZH+7rRwU2HGeVyboqZhuyDWz8OlR/LcIHzTMW3pXMhDc6rsMZPdkuvk5
b9oBh3tFcco6rmNQ9/5xGiha8g0pHTNTx0Ji6yrPgJ/S3tA3fAoVxusoo6tUwZ3A
+Wsvke+xwnXHaEc3P+kxRzRSt8SWlX6Q4Qa7cjoEdY2OZ/IMcwIxAtM9VcTC1qXj
a0eonNwI/utkxF6LFvDq949FdSsF8I6ZXXgYkxO5zBoTq+8Z3ozFT7Mxd3pLYKBu
L0fJ3B++cTAd9ER9gksvY9uXjFQ6M83jtNQALBfgr1bqJ7+0+fyH8OTWS7C/Dnmm
5DjnsRFOUdBCzFR3LZPDpmk39MjYlwuZUontDsv+LmhHQJGP5GtsgRZK8hfCtnL9
Mc11FyGHTx097F7SD/yD49LxTaDH8zJzskWxRBboPNhbDj9k+z+doDFK9NMjuHQ9
aW4orTlRffbIBe7KyFjOIFndHWIY4qwbboH2L5gJfyLxRO3PvRnacsJd6M/qPmlM
cZAaqMCiyB2RgiTZHAnkMb14+JVYdoHWwjIBtdgUCSwgxYZQ3tHBZ5y3qlFVeiTE
fOPknvOwapyDf5wWP8/CsCWiPlnhAG1kSP6VPPnKlvvVp5VlbhE9M6fAuXtKnTDV
rNkoSU4MQr7SKDLe5vbNGVJZTHW2Ow4gVtxR6Jw4yFWfYwy3rma7rfVeBPiVsXoM
QvN1oWkK1uIZ+a7C1i53dBWOJi2n2cjtHta7/zRFmjTi3SZmex3Xz0llovOfUdlg
f/dRpdBPSsygzH9s7vPfX3B7W49sXffF2N2fH+Yrb0oVSD7+OCJyF10VURYjv/Xs
fhcZFp7rMt52LFSD3gpn7/N5dBUTZ6UA1BlIzTKQ49cmC5W59L0YkdemtsjNPz3A
lnu6xmCLsl6tK3tJNAiTM4sE2uOnNgcuAvpzRmmrzEU3TMsIVKg0Hv9451QEJHkY
e1jEAB023Zddn2izMDTD1DAK+SLLZopLNVji9KNU5mjd8j2yKAFC6/+tL75JuHHe
R47zCCX52flY0ysHlcl79fFX3pHgRDn9X9skXXr7AND1QNCVc+rnLwFHe9tx16Q4
/ff1JPdFX+WmyTi0cTx+amZcj8ZEYFIb9vpaHwJ+o6bQYWYRu/M6SDhS0/h/xuuj
jNahq+FM3kClEkJXU/FQZujVz8rIvXnJf8WeJ7KYbUFhIuITQDvq0gbtrfFCHkFg
5rUKHdr8H26Qmdb0IKnuNilFI3lI45FKqU2DcFl6Byp4TUN4p9M7LCyT77hoMHQ8
OWKxu6hDse8EEb4CuT/eL4fX1gHF/rV4waDcOl4gJUqIgMmPbblJRC9zegZkussM
JMrrhVmLyWImf5zMk0TV7ze8umUG+v1X3H7kLUerFlJ9tegA0qusI7vJ3jy+45vm
S6fnIMJTSyl33yauEC0Zhfz7iMxdyTrGJIbKo9+M+WQpI28cudQ1eyy6u91h6wqc
P5SY+rMqQ+No8DQT6Qvw7MgVyh984R1FrpmE4U/as/dKeKpiRB6bRiSQSIW6dwMz
40Lrr3loqiMq4/MefA3+lbM3TB9uCYEi7ciniWXE9O4ssM8mImdW2g8x29IS9M0I
FrZPUyknGHZ8pmAnts902FIkwAVnx/22konlbmuFw+KeA0IAZjWPZ3a2L7ZOak2a
FYTdkLK7V09exozbrhohDgZOt/2SOYwDA10IfjMxloNVAkZCCAar22LfeeSW1B7j
Xx7kbpHHG2qo/E+tfGMY+htHc3EMSb6ph+9r2fJgZem2XWvimGpDCcZ0r7nl6Z7x
Do3DFbwi3BA/zWH9YOQV8iyysK2OyNEO+MijbCXDb2i9p4xPgKSNAvAhFjr/wkWF
8taSwt9p22ZBKpPkGeBA5g7SKk8vBn8tOC0ykYHIHy4rVzwtn63vP5SRDS9hq7nt
xj0pb/kL74Xals/a+9QOcsvcmgK8hOrpTQKzAeUcl/23e4xaMPWzeUEJ1WwDfGhV
Miy07ObRj+2QhGsWWePwuus5y1Gu4CvHjYFS6XFNVAX34ciX+TzlMVMarKcTVZtm
nfcGrWzJWIZXNQF8HAsOl7SRonEU7y9vT2rFkc+cgpleTtA7fm9ECoDv9tM+awMG
ajHxiVzNNZVefOzyJD3YkmwDAX/GSP6gBSFyI58kpa50PgyTcCX5B9b1CCOG7lyj
KlAdTAwIjWAI6I+VzsNUhE0ZG8vCZgi+dTvdrC9LLmWrwI8UYPcwn6HFqfj9iAPD
Xk7tBSeTvihN8i7hc2E0C0UUrpZBLt/LARxe4RkGixtbBDsSU/ptNLjM3C4VmUeW
hMLbnDXIAHNB0iMPQVCYF5LCX1KiZ1OX4+jn+7tvRXnl4lK9f9p8Zu+V8ULBHfya
yHnw7p8nG2q/U9e7gDCF8Mggw2QgK43UgQggmyDVj0Jwe5Vz2jvBx+ymYOOi6Na0
6Vy6APLT15w2D/Y0ayCkkFCENZdRgWza5yzuwsCgKvhUjGJgZSBr7talUjJoGJJQ
6qve+bjecZYl0mt6dQQVjfEu/wPtkOF0g2Vn9WR/pd+Cq9NIQXsSkwCJ+YvCPrOO
Vvx7T4fVIVeB06KPjVGra6Z7HyFY728g1XLwiqOhQCM/1Xa2pH1SotSco8gu2kF2
wXe9SJhit6lqEGUTBxOwXrV98gT3BIEeunlkjAONR1zgjfGvFgVvRcelTocSAk9Q
EcjwR468xx2u4lamLdEouw5Iqi7lkxKx9/F2RdgfW0cUl8ZT1bh6/w4tgitv/duU
uvt61i0832m450TcDlV7eT+g3fenYOiH+Y8hTYcmPzloR0D4E5kAxlPvpH4XPQov
djQuGerWGv8893r5VozRL3zxsjezsoUtbVj37t5yt4wUm/YsWRFrccsbKBr86Vba
GVGWXrkNaOJ1GheABNRV86bBnnXlO7TMewuIgr8UJ2+3C8io7tZfN86zuNUBeKCx
kQgt2SvUfkbESOiK7OHEmNi3cdZGSzauSCKXIfCCdhl2HeHiROMwbv1Ip2YOOeyN
vkMDXt9JNyizFhiPWtBGwF2kMUuyYKu3hqKuZLlqFTvI9Xi0DAEUrtdzjomw9JUw
dZS57Cm9i7j4dQzfuBVbSv5bGOcNy3gAkEZ/xK0PCKmtiEy3psc4+QuItxvSwf/P
IsFP3cDyzWEd8bC0UJdySjh/JYPSN6WmwgQCi6welF9KDj7UFwJeRNdS0Uc14PV0
wR7ZyXoh2tNBwe6z2Y/TI37tXK/V0Igc3g/ShpwVMv9F6RoCyvT4ewjp4wpHuMCv
H0l/4BqhmS3ou9AgXdBp1brFFbYN/O299GZaVe2Uz2KuGNiCJtmSGrs6nXxY+9SK
1QeeLm24eyPmSPJEr+GTP6LbxeLGM3UlA06CpspVUb/Qq1z5NsQWlCuOZbqtbKI/
AIwj+BRmU+tNztEkd1mqhLL2VM2LTB7Eu0Jjme38oJisMeXq7lhEf6xedrQmWEU9
AXgo6dRtK2GQWMEEyfD4JUbk31jJBoYYJAUL+0TDKbETbYhXoIuC6SXRHc6hMmyR
J0Lrr/gpreTxMzSF5GZAVUxk47xLp6LUNFyNKI3JRtCwapQLDk+MECCW34BWwEne
krIriSHFph09FYdjIyJXS0VexmWJOPmjJFYt9ToZ5lN3FAO+m2B/5HTtAfb6If9T
+45YtIbIc7IB1EWyYDXE0AyRBTrN3mGiIPa8KOz2ySLDLlPHhn7dhIiRrcDj9YBE
Rel8n5Y93W+bbFK8Q+hUAqBG8Vby8fg3nHiyHYL5sa3khghynm8h8IjoQd1qAl+k
Fr+NEP4OLTmTIZsQRhF3hdo+xSWlA+H8fS6b1RZ3QVuaYLQ/zMBmxm3GsKEYH8Rv
3revLsOdkBMTcVM39H56gzfWPCjJH+pUOrTBXHVMfOshDBMf7Bl4/poflvUYH+Lj
IP5Uh/mEEx1yt2Jl2Yzce+wGmxT91+ypegFm8FLqPtlUOfTPOxnOVbm7mMzgHelm
lkOBoDP3DR16U6oJ4Z3nJzU9EPolXGW8g8/7CQnXkGSidGdYYNEYtTUNBU9ZSR9e
HyKd1B4oOsVeZkiSYq3puQ/CKgMn5gRTk1so4sfjmU0SbnChwqBY3WJfuz2XGoSp
4y/qJyUR4/TJcp49xsc7w/ce+xAfkrTWveyl3ZsUFWUrsqcAU18mmCEGKBNa/Cig
u7/IlfA7ZAmfNtGOLg/i6f2MS7D+4ZzujH4sEia8/b6X2+mHaYaNAHM088PvHV2a
Xo64Nbj6QoJ0KuiFVr4eZqvswUULVhBtGUGkspsyUeXJngLlWvysXOiHlDVMH9mJ
KkDBMFu6c6Tix9oXRbAElZQBVz7lUbtJcD+fOCVZzZVfY67II/hQqIY2jNDxYmYx
po2ZF2FPdShdvNqvKaIWG18oGWFijcz+bq6PeEyCT81+IF/eDYtaya5F2LxmCbH8
7Haji0Uj/4ULBCYkRwGjOsl1NRQd+MW6fBu43MuvSrUDce1lnmkBpvnQFKngQPOX
3DCvc4vqfiOqY9j052rWJBP+2g4pordo5jQ7MSkLyXayTcWpqF8xydpQpULiQrkh
HWnNcW4ALLfaBejRLMMOhLJd4nLmKDfAvbPsR4NB2zD8ydzfRhLAh8OD0ljzMm6+
pKGjr3Qkjh7nsj+I81dUnJ2+T7DJnwfu4K75R8RIkIij8CjrIOaiZCpbZ9cbuslP
jSicuBoY11wIS7A+0AZD4NoDz4jU1OmnnRLTOWolk0akmbqTg1OjLPrYWcMRJ/lr
ipH0hwOmle/0rdHPxKuW7q5o6aDpwCoBw8ByV39odiofUbSAaLRWaMWpdyaAcPEp
T+XAW9/r11TrlrsAyrxHU2Oh/c+Ls1BusF7jxFUSuUVBJnhlc70FoXV1IlvBKG/K
7sgbEIqlagHY5fEdmvMtpDaSXAq1bO0rtTrZWvEe/ySN2ZOg95kPGiRYNL/smfi8
6wk3J6OBs21WmJQR4sv8GulfoZBhfqzD+iZu9ut0Ebo0g+tcBI8QfD/Laln7C8S/
crc7hDfggDTRpTwklNF2UrqLzGQUueSw80cFXuG0G6bjzcxoINJGl5Hupdx/ScWy
5usFb5A6fgCdpTbw++49doZpA1dzcM3G7rhPAII5PxpURPuZad2KDpPNpDrhUftV
Q37sEx2SnpsSGZFSZp+pclelCXNgE2f6GL1+2PXdstUNfdJFeR37doeCOXTf98vx
OctPbNUqOCdcz+IVeCuMUhkeJyeNLjs2vEUC6dOoacnZJs64Hllz+gQzWVWyYf+6
+HqbUyKoiBM59up5BvSBZ4dvnoa/cHmEgpOuLrwv2b8/JxLBQL6BAe7tkNWGMtfK
Jry0koLbkz5iC9Mfqrt2Tbjufxxu7Yh5fv/dBxrYqIGKYlWHy79p/nD1OV0adV2q
X5FFIoEIXScciZht5XsA2W0du8jMITvblzj67oiYhvws7lL8oAQ9mMQQVZ4OMPiz
+31kCOEgO+flMCfL9uQoP93gOJL/em82l6qzgYbQibIoos7ANdfXNrD6Os4r2t3t
9hrAwACmrhvOdfo9Lm7+pluTNFvoGruGIrT/VEdRF2OA9uW+AQmu9N1F6HReWW9c
B3vtxuXR3118lf/0OA34K8/RBkQB/wCfXXTORtEatkpcWxhlNUq87eT3K54uLbm5
JL4A2aBs0nCINr32lSzd3dj36e75CM08pRSr12N8hUzksEaEPXBjivx3LZICN+DW
/5DBIAQwBObUCiivFYlUGvgeisS8SPUQcii89W7VnTBjobcO/HDFVzk/Z+FD6eq0
U4Hq2IxfsR8thW/KsP+v7qLWYF2D2XOlv3u+CFFoKX5lIxu4DVvWQ8aVMt6pf6hH
wERea9Cc3fwAr1nQMMX2sstvg43EgFSEdnPPDc+SdQdxlxvSDm5Eg3YRipQXluWV
wPx0V79dz3pbWdNV1HMtKx2iLBblNZ4ozrCd5YGsqjqQnFnN6rMvD4zE6NaQ51nX
oUAxs3uxYDtHFCDX1jcAdtd8yxpyJxnTOGgdf4P7ryAmmERseGVgohMlS8QTM6ju
Og/laEM+D2+QvNbo14oBmztwuTMdGFKVFzPJyOcuLNw6VvEIA2Zt/xV6UdNvTt/5
Ahd4+8kbmLDlhKf3TdZblMv2l/Zgml03OUValcpzdDU0WIq24Zth6MH43H+NwxQ/
S7zU5/vMnuAPA9Md8Acky6kjLsBrBsDCKbeULyW7+HJoIRi2D/Awo6cvym3XZtQH
ukZ0ZTmm6u0Pdh9G+RK17ki7bpiBV/KaBmUeeYkG6nMwBdLwgBWIXeRTlWl00PRU
IPM3xZU5FLJ3I99js3fKCygrQ88+XTSjRgBOhHyNHa97fKyNQbHCYy/jUdzJsLDo
IOTZPm/zCE60/Kq87uzBVk2VSAiOZQtaroOH1Bdh45Q2FseCkoo6zOFOFEqr7lQH
Oopf7ojMt/1j2QLXcNlSuIGpYgBMPQVaLSz/0MuKTW8KIhsBVt0CjpvE33Y1aSkw
EFWVXjZb7RZG20kAYcUqyqBDz52ItOx0VFgeFda5c45pCJAhxkFNgYz4kb4RZxl/
QNnit9evJxvf+pARgdgn1i8Gr5H995a/O73iUNZ79K9uqRKNfwNMSkzQyot1Vyop
TPapxC//T0jHAQZ6bFraKH4fvarU7LDHCUMdXMmwAVkV9z2JScStSTganUenjRjC
B8mL/b0dK3atNJSdMPgDwSVu6VcolyZuJ5Z8+B/DAU4o5sMf57E6cP51Yy17QlyJ
aUKFn3qA/RlAm4cby/0QM1sfVQvqpwlq6FzSM2CTGPSsNGyu5vMvxR+PCQzinkhW
SKFx2oybEyRGFCBKQyOF4W8E/u5mHDZpVjgc6ICuNy0aTXiuj34NGIZPpXX5y4ov
AkWNoNeQIhcTWg/63JYq+4M1GU1BOZR1KE4pB+zaPF9NKUbk0xOlE6+d2f7br/v1
PhVHO0HvmQ0BZL32nTRabUMqeMZP8apuSvw+pCVi679GqqmW0L70lAy16RLF3YN/
avcafeSgL5svW0yMzHPD0RJxYB8z8mL7eTkWuGlZwE2xIOpYzl2LR5aOpMH7WNC2
nh56MuRdF124/iPriDNHy6gtsP2UTmZyCsvQrkgDjuIEi3SJyRMhQuIjdj+Y7UO8
PizoO6OPLzzf76GL/zkwfj+YVFnpWypZ/Lp0ebhTTgG/p9FKKMwJCytDU4kjYcqE
UbmZFhmZo6X2yuwEkO4iuYtr1NrCwQkzdJFOL8mlrJujwlwJZyFlAe9ewaMt3cj1
LIr2X40cwdLHcmNpMR0ed9UpUwE4KePdqgVif2mXAcuZY2B9YbbhZ0iaOyM67Or9
QoeQ+V0ucg3AK0+Hn3CNd+b3n0FmGnsZOg9bsnJ50ozO6MKhfk6CcL5a88ASLJHN
2pMl24Q8d36vX8sQdFvPYxvzSuEbwfFfycLZMUQf6iA+SY3gLQ0hACpp4cfRjHu0
RGRyjI2xEmJb3kNMsqBh3Zcok0ODv43Aa5BTZKKglgrvoPXsUsz3kVJP9opDnOsn
ItFuRRaCCrdxZjJ0kaeP9MHNcpAthkXFPQEolTtgQONOw2KsUe7KcyLT6cUFmrLa
Gn40Mvc/2DUvf/bh34B9cB+F1GZNmTCoFSGQ6ucSKlDeWangr7ziCoduOoGUDvy/
JU/NwH7Ews18H1FIITAbdome8+rUWfJAMDhQUdQtT9pRz5mSJ/kVC79EHM1QTYUY
pCixCxmAtyNp5810N43pmD+dymZIGFgZq/ZMigiI0WsyTrXWmSNPm3XD7yk/vEeg
k+o/v/bI2ItiJbHkQwogSlODFc38AoKWaBkzSPnU97uZDV00yp33GT4wolb7YnD6
tPzo1KGEX8mYEELviCBCrUgk24DSi+/msOFdT6RXJAnvN66YsNOEB9STAZ3xZArV
lCvddK/IpaBRDt6I7Be5pA07dsXpx47bT/c7D1HH+TsPMa6swkw+RcYOOc+4mf4Y
sQzaADIELPA9Jb1+8F7mF/pPcOwLO/TDs3njKgJqQ76DYCbFDOW/d5uhtUBIiOCH
aTzp1Hm1mHEVQ6/huIdjQbeWwIsbD+ZGp6nVXq/nA05e2GNJnQ0dBCW4G5VnCeZy
ph85FqlP5NLF03Q+RzUVtHedgwgasNeG9CH8KQhxw9rz+PZx5P24OcM2aDZbe5gg
4ahkL6QWf4kFNKn52xjzKc0J067LLogo+JkGxY48UHNLPKsTxefNWvCe1UvGN4w3
yYDaCWrumNGk4mMsC2pNSnXO4eEiTJaRq9oBEt8njOguHyXWh5SvSkGYfopgIREp
i0/bZK2owzR3oBwI7vmaG9OwwZ2sdGMJeuZxAua2gIlywu/wPGr1rvsaNJZ1Uc0Y
0cHHm37cg4/TcjZw/v0KVcbwUqi/Iytep2crn7wQCytpFHKr4uuwiIOg+s2PuiBz
AJjZxwNP0NoTubIBNHGahjNlkm9BVdw0GQvj4m1xykV6iG+c4uJ2dRrvGlPnWdA+
+0ETnb/DWHqCgP/w/oLLvNCGmLQNijnygDvDcdBtJnf7MB5WqcWoQZbVaawd/jON
Mk5zKlG07nfRJpJX6c5birKwfdmjyMfNxIHZ80EeDlXiL4Q3IzEcT/jzWtXTrhZR
fu7jQz3w+Kk2fZlMmt40QJDsIuu2nOU8UhMqMbeoJx/aveo5ngZ4jv81dGQKzcez
qq9d+XuxBMUqQvKIgg6QHOQnLU45K2M8oMI1Wn0C/hvsuLd7SlQ80TjCsT97J86B
+3rQHaz+sPVotSgF1ZQxI+hOW+EB/TuLUklMqIt2LR4e2LCJYolBCrzwXrNx9Fk8
+fKjxC+ZYUdWHt3ppLlR+iTthe9pcPrDDKLcO73hc7/dVW5oxenuyxqgjWXXAv4N
LUq4OpxDPfA/Qlu0G2J2QrbWNeGeSL7+xqHaXtHr7/VPtSBu73KWcxNWiCagiM3v
1OP8OQ59x/y4CDRWQbyyOjbFodUMu90YijAeEabkFWJscZQ2ttlVsZsl7sSJoyQ7
RgsQuFvd2eygxr0AyAeuOOxaqppQYReIAN+3Zx0u9C5Ya+Nb9gZ19YJ+PH+wccTx
6/3Q/y9uj1duJD3NvRajI/frrDiw/uuBtkaa0aVmhL+Gdqql+Y2Y99w2QfqUF1xk
lwshsykR9QD9wqZJgi/X6scAjqj8oc81vU/1oew33Db5ld0yq5gl3E947UB6SedA
O4xNtmACKm/6HkdP9yfPybazB6krKB7P1QvrqDeN+KtMrL3TqmBAWM2NZOCiTBsv
pHsgRnFgWFlPEOestbMWNtB4xkXAhZl+uGCmJffHRSnOeMJ84KkXVRNmkC+A2K5r
yw64k6ObENgpbzqWTd4dWIqtHKFKtRtZbaApGW3dOrVubhtEytuxEYqWN7Xhy160
nhHekk2SH7YP2l0p+ySvuuXsVGyQs/O0YYZY72HP6HwB5PMmVhVnI7JPTtzQTVns
WAO4xqSr418qkwkazSII31VfHnSNAO+46CtSo/PTBtmDGHiIUfOI3poBeQpblDsb
L0vmppHU9QohVzDrVYWMXgWjUmQfSQN89dMxqZTnEf9+Ep0xW0W0TZkOmyztPHeu
Ao6rz9D/8MFSt385vtjro4bVdNS38aDKulXKyHMprzdEzI7ZbzLySeDSMogvBrNG
BjAkBH2AE4Xj60T6wd1had9pFSO4GezKvKPNEKFu2hnB4ovJJkw4XrPI9Za6YH7c
GntuVV9BgP0xbTZG7phdOjAdcn51Rjy3i5oncXHoaSI5B23t4YDW+WM63L/5iOWi
i+Wync7x1I5rpVkKD3O/DktB46tUCqOfnJATKK24y4YU7Q38Nml2kkATWZuwQvcA
yThA93j36Ah0hy4gqY1UI/6+wZfh3mj729MWv3nDEkXp52n2wYAPHFGi3fMg4vot
wKWeqJXuR8DxGijiM5Vb7NzP+pQkI1aZy4r6KlF/WAntXFb6JyJllIJ6H/JGamh3
OomzA3aTaoCgYF+Vt6mk5GmQB65lZVxauWUmy3tLCcGc1UuTZBjWFwEW2u4FHYaB
M+DbpxHKyPvssXzV6T6ns10SmS7g5/HcHApYunogUuIJOn7Epl4XTVTx+BtHjMlv
f/vIeNRSNzcHiDjFHqy9R2Nlhj4IKUqMAX+o26b5jfwPJyWwMutawsXtigYQlMLx
tVeDJb1zErMg67epN2JXGpvBoWQW4A/YHXUXwwS/T7xEImXW9AzvPo7SVp/JEGIx
cDQ9g0vCseEaKGjt2WGSoijfbAANcrrFnChNqfArLto9LbqnVMR8kjxo2y2fpx3b
PyP8kF7G8/ERikq7DhqUj6qEHTzBNTarpovA5wZlLLqcsrXOn8x2OpJpQN1ePujj
i8CIMU6X0V+XWcjC+NLyESAtE2VauZUucPpiPJ+zZV/zYbm79WdFmEb8txn4FKE8
3z7cq6TVYjHUyFmIyZwR8Og9DHAPSCzzzbRUqFDts3VRrU7/wdwwAkHB8E3gC920
rzLtM0n2Q6cSQqxsrA5Sqnqc5fANqymHBr41xx6cI7kcsOs16Nc5Z7+YJmyhvcWp
Smz0/y2oH/byX7+GK/k00olQmHAD3ZQQftMTX2Lfa1DdVGqa/SKZwTm5c14ITT9G
ojNuw1uAgK1p3ujLSc/JsUMgQBY9azP6qJzolLXahiP1iERYsDT9yy/P88ZE0T6c
yovzEz4igTBc/JSuwtvuXPvkmZCqiQWn79GeKi1uYMy/YaHMC3QsjLxWGSCZbC+S
InJ8iujUFFZWzST24CIHwOB8X5IWrshHUaPuOMYflc0i23HkAkmgGLDEKj9tX5GP
8aCiibQNHBsqA5rzDm8gn3FikPDtsLDQL0Khrzakk3y2IoidQkqgjIUrvx11K1nm
vSq4jUJYLHcrNwFpKsIsUC+01Qa+UfesEqbSPPlEsFA1UNsZ1SM0wbyKcz6QD8AZ
dyPHlWO2J7Vipy4HCTHqsIYDB5f9cgdtAQ0oHDg0EuB/7IOrJsbdDkCoytzb0UtO
BHGV7K6Rkl5W5W9AYbBAcRlxFou7HP4MHXYetPeBp8ahstcEqxTVjiqhnEfUh5Gt
NGiCqQSZaL109tIPN2sOsJWgSKNR4hV5cNJ0QMNWWCXt1ilIUKUcvkEgdkX8g4Q2
jhF06pKACrwUXJI7nVnxmRhkEobyiLNRujTZDWf9ngKlW7KV1oi9GDSo4zgjAXrd
/xSBNvINYqVpkji2zVMMyv9mFh5vZ+z5Kc4SAdRaG5O6fIhh/PfViWAHbEvSVZDp
D39/pqJ+ZDDx7PFTHhZTy/erfBUlUQ2eRREIwDfzBM6aGUEkFtI1iLoGORYmYIr9
54jY5tcqW2+EDqzQVYh4zAkVNizEglABk1iy1M2MkGM2qZblbfYvRndx9eRzNZJW
76ATKQtpLZbzxMhnZ3fSSpp4+/iu1t+Ik6LuYa5pP367ooE3Kw54ijPHJDijuJbc
AiUR60AqoqQIESde1IratKC0fr2iYo2w+uskNdl6LaZIet3mTAtu+qlTC44Fgx/P
nsqZSfY6ellLaDlkx7KmP5/2F6nMCdyfZ0Hg5HQ76UjAjhS5LZz+ZBHSfUFnRXCE
jmxpHLQK6V6A1IFZ4wUweVD7denQAft6esdcvJ5fWwZrANsz1UmU/E4DND9O4H5W
KDmeuZOi1E7r9S4M0dRY0IaMhXADFDePF5NILMiVFA7DZNbipEfWXQJDq37RrjTz
nd2JqYdBqPoS0dGdIorsGfEd87d9XYXGOyDE8CxQdNCfob38aVEYZSJ0Ik/il0UX
vHIOs/M1Thz303A1YKyM4K8bXC8nwFwaf8gP0c9zMRzNuxiPVAAb34EmdGOi98pG
ivGy+HKJPQlMQrZq0/jMp1Kb1YGnh2/gZraOtXjVX/0H50iK3Sx8IjpoaPA3ZMLz
RpEeu/4MA0w2b0UPw52qnuiBWQhs1MiMfgMajq6owjjequ0tlwtiiR8oDLHoop24
n3kIFNq037DeCBPlhzi0P4RnOUIbawkUzCVfTcK1bjwk2MjdiqpebP/v49AU96E3
l3vkTRQhM/owMcs6qCk79IDhQXnk6ZEQEi9tkhFqZ53LdLBIQlwLrFhotJHPlnYj
KG/OesNAeshOQSaVVOE0Zp3qaM32zGdaeEtxQGhHsPq/8SBA7qQEK6y6yAzsTH3/
qSm45OTOHzcpZ2FiWvHuxYQCSdTCPwbUlSD0zA95w57MfUwYZ1zsqrDuMpLUjMhT
RS1KaiCKJdVmX7H+4ICf67BBcJorjitEmCKnMoNCayoahHl5DZQiL3fTb7t6qK04
JKXZQmd4AD/V7Sptk9VFgmJqOKIqeY4fdkQRiyGgTYgceplHU54OKN4e92zvQAGI
OfGYP4QzZ1WMOnNsr5Prjm0WqZizirkF5cMd6j6YZF/a4ftNuGRILr2fDA2eCRKU
J4nYJO7fKdn+yW5rdZh9CklBZLbVUJYhkDW/jS/MiKYdcvZ4miyAc+ceykOc6wsd
uiViR0RbJLAIsCk2HrcMvfbHgVPbUCpvjEvINaks0/C8bvigrqlAKXDbOXT18LfO
u9I6H3B2dlz5Bv8tJnt+6psIb64lqWaQ2HqvZKNrIcj3M+k3mBSqz7Yvw4COifSL
tl9ssnGk0y7RGfnUPq643I0ZzcfJqfc3Xkizy08x8SCBnrlgMwfHVbA7TZZK71ic
KGiNM54m+oVgL0i8pju2kvNPW5Q9++NFtqlGRlNicz5ZciGd2udjSrQulsd1KZR4
XQXX/BOAKxDxloiPO3lROu+5Yru8/Axlygge5J2n0DFcO7Gz6TuiOJQHNEiRQEnJ
r7EPwXl54UppTjGfBZ4BRh6E3/bYYDqyCJiWmT2XJAfbBkr8MQkmx7U36Qfy2gPi
SC1/JGYa3HN2m7UXrZUhY/6N5Jgvi1rNahMVy5Pq03v7pHIonxNTFg5XKabVvqI1
uM/BqGto3fQJ6kYP44ABmOlnWQIxDhhEOcMeUwdr9qfOUGAjfKZTQ5q31vSz9MgC
GeBCngH3vvRpfUnbDI2y2P5tQ5/gR/LkZfcl4yFJ/SEnIyxBRb6AphfAVgwy48Lm
R0KG8V6kdge5YoYtMQOxBmggkzvahh2GX8/do+tjEO1Yya6zlrgHS1GaFnkYAW+H
1sSZxuRkGpy3b+CsKbRIyqGaXwq7jmaiaifVxlBBKVnLo79TeOBa4fH3kFs2oUAG
ZA0C5zBtDUhRJwcSTsZLt3DMf09djm0phjdEdHsIclQE+aEMlyKaI3PNjAYg6H/d
v6E5BYZPYk8XkFDuz6AEFW5Dz8VcMD/ZMwjAZaLjiWVZ/IzwZULA1cozSTUMK24w
pvtYVlVfrkd9AUzmJ9Y9UGDiEo1EQQI+abc2qn1QmcGxonu7b+mcRWzcioiWp5cN
rXdnMBDS+EP+P40+oASHKpbxUYNOPVjv7Wada9+MwsiJdNIapNqXx43nNklUGmL/
Jlwem7MGVVEaGNsJK93Ur6tKaGxqeB2STtlw5HvXw7NLaaKkBl6/HD3KbCtLH7yM
EXWwWbDs3pYHgNcZvcw3oCqub0tveU2lybK15wVyDB5k2vPf5/Xysi9z6hZHgfHu
Mft/tt6Q1740VggS2lgtsKyvwt7YqU99RawWkF4+ahS7tODPK1R00p9sTBeRs4g3
ybXOjVm8//49ALeabwFaStTZ6YSS7oxRCtITO5xGyY//A+qao65ehbshVTUVoftd
B2VpFkM44eM6RiRlQKxZe+6gumn2yDBHb5xHkYeMgB0cUh5YAFgb0YtV2gNNShaA
FM1N/p2C6yMvWSOy6ZXYGTFA4D6vIuct0/sMs1YyVoLfCVlrbPx1VzVjC6tVpJv2
FXg2MqzPhC/xxuL7NQuF/H9kaaD0+Nu1gRiydSnhndl0Bw3at4xoEbab+HH8JyuP
pkdmgBhShNRInEVekeGDSUMYm4vw/FrMLX26iZjlmckzFwUam3O9Janwdcf7WZQd
OTo8dOG17yHXpztPrbEzDc+ubRsNbs7nRCxFCrBqxnfgf1oJpr9YBHln9t5Z5mL8
9VSfiwuUyj9t2domzdG3KMVr70X9EcD3eg8B16YUzuhBQYyMhDJf4A/iFk15PtL2
fd+krQQjtdsmL81hlrRnaas5zJEJNB4EQeeOKAmGPx+pOChYSPdpejnN/9Re26na
kMBP+ufZ/5uEDTmXXRwVO4zDNeO8V+Z1R7SmjL6IKpcA/eKMD1wTRkl3M/J//b5j
JWZvkRbvzGE353Slw2+ktG4Lwe90LibaDXHw3gJl/IsfKy56maLJ4e6zpztTrrg6
8Ho2c1qjpZgcwwoQYQoytQbS6p0lXJwrDz/QLJS/qzYEjcu5PrlzxbFjSBa9bBWC
oIPXSKy1nxrdvaSTQ1mPRYmx6jzMJnIyfFD74EL+ULtXpclrNY9ebmk/ZEAfnp4I
dGu6mc7k2Gl1q61rsh6N3GTI/VIfejhmVGErABlpd1cJr/QN47b4HMek+ac0kVeY
1fkeIvFcBiCPiL89ugVo2b/Up1p8AHaXOfYBsi/RKWdQgWAHT3IlVYnT1PZ4Q52m
rD9vSAscG1ZYTKcz3f1neL7h01m9xFuLHrVuHBzvfpEBYVh4GWFtQ1FPzxvs4qU5
CP2v/9tr/FZN/y6p/MiziJ0EoZu3QP+0GVklPseavmH2UpU9rbFr4wAc0QqVvawu
WqhIUt+yYI/kEO6+UkUVjBkf6zOQnXiD8FT24zaZVNnNQkymgRDe9i0J3J9G0Tze
jOB2IZhHYP9+/Ie2Jig47AywxD0yDS6dOIhNYdw58otYzhbAoyZcy1DieV/Xr2a/
+166Ips6fhoUDM1fhbAugzJGXb4yrvdFieKxT+VAZZTTFQUfmo7Ewz9yf2NpY9bi
PzkHdKYWj3AeCv9A+4xTuNVFgE9SFM42puHxr/mRR2Jy97vkfberrSy7mBy4gWON
BJJC7mHkzWp6W4CroDXw5LcYdJ7dQa+kEuTkJSe37Oc8V6TESGkgDls33N5hHHZ7
db2aT5jBYgcdOWu55snnN+PAtVYX1DuJf6W0fnMVkRPV7N+S1paWv/as2+dxoEOh
Q5zOhsyKSdWeIoD61oeRzkIqIuxpiq/cWoKTQR0EGkdpXn6CSMBF0sRglMSG04Jm
b/LBGTBO0kMt1QAsL73ZW/gxZBrdVl4pMNBdHkItYkZODiAGd2tJ8hjiGvrH9fH/
PCYCWi1c0ee4snTso1j3c7Fiw2T829TSiYHLBxx7A02MoGuHaI4+xdKdKFj/pIq9
YZsO4Esy/8CAJurYrliOiVDA+na1r9vo7g1nBGvwxJWrH63KcSsTw+TX0fzBiJgr
5pL47hwVLn/SjFWFMOz4DK5hHv98QvHlLvQR9xI2WGssLbEijnBOBlvJQ36mOKNb
HgPOG+5AHHULxmNxHhG2sSgOeLi1jNw+KSnGSF5HwMMcwWggcjuAt2fwZOStj7eX
ptgjpCzaMQR+CjF4zuwKYzUPgfhXaKbiArSfpLZgou/lNsbjVg5Z9FkQkrUebNYO
M0RDYC/U6osGHHSlN8zN7+YNrJ1Rxa5gBA7o4IVgC+v5zLIoit3uO8GawtzuheI8
mHxPBZNyVLI1aMc9927oUoFDFCJ1qVNU/qMHWewBLux2R2C1VA+S5YkpYyYZE7nS
ByfjvWmvGyTg5p3Pkr99iPisc3O6OarEuCL80dCy0YNMSIpOWZs3yYJriAJ4ca1E
Uz84z9UWAxV7aesSkGuWV2gSGZswiHP+aV7C7nSj0IikQLOZi1MrrporlqTJxwEk
hv5ckR1O9JbH4WTjOtC/wH95B4u/c1nAnuAWPdVEgCqrLLShdi+FzeJ9J2qPYsjv
UnrJW2hBRYmubjBhaariQKTh12Hb4D+KrZ1FnMyGGEX40jCxOTO/ldmDD22Loa6R
Jq9r+1tJiacmPNLsP7LmX0+Ar8TGSmjUOpx/uB/yWR5b8qsgyCXL9FV22Q17wMcC
sznm68EGc97erHzNsmDeQc81UM4gtHnMFw9gyutFVVw0QuMrtAzhkmPj8Rb+H9wU
nKZCo6I32xELYc0PgIco7vTdYkHRpeTzZHwIuFvFuyXlL9hmTi9WznHHn384QyFN
4r71a9VOp+qyHcRZnJDl7GAELy6KWSgGggFqCgrHVuQA95pZ1uWogfZVPPP8QcDY
Ng1Se+5adApSo9sTniYvBty+nFiT+rn3ul7+JxRIxJ+fFW5C3L0gbyybqn+uLZLM
9DD0Ez0T4DrJMu+oSWWd4gHhb7vKNWSi2V1qPqJjLmZBnUyopsRcP2g+fbVU7Myv
HufAc/q1a/nkEltf65Dvr5q/Jyun53fvkqnnR2osPndrUoU/jWoDIA8oD8qOdFhd
RHUknCob8mMQztw/QgndMDa6MgqojDjwUp3JWMTuiA/NsZiDeaklrFezwk8xm8x9
80a1D3S4V8W3mLb7ANWtKCY3NQoUbU3F40xol5PkMUW+BK4I59iYLAo2Duo4yQDC
B8uU/KDEqV72ie/Twg4wOGtjTUJqYLCNHwETtLxq2OYFR9uUKER+YQhoQ6B08gju
N0mccCuER6fie2dDz4uoMmrm/TEMxJ/AlAibDBTJPpzC26IyvOPwp77bCqycu507
/BGPFxxrt4SOGLjLPCaAE+W7lMx6sOx8hOmrQ33cerr34/QosRaiQNYgOb1wA61y
gF15T2TcHmPs6zyOBwTSessRNp6x4q6KtbEjdTEyhutR2dCUTv55cfok9VEEvTE5
vPoEuJALimil1bZmeo3VlRLOzVXOLSQiVlKGPLPQxM54DiTC4mTU9hkmH6GpKj29
2qUKxCXBYe3AJu80j8ZAKszFRjGDmJBvh2R+OshkDx+wFE945/G1ocQypwFBQrUq
EYEhbkhxPSQXUQ7cKXgdsP9nZpvvDnqcnanJcE4mBQg+hLvV0xoD1aEomEZgB+Ju
XbuPa4sQEBDeVS+Mbqa9J2A1wlHi32LLp30j/2hEOHXOoAYlymb/NZIc/+BhnZta
T3jYdQrtDDgqASZ6P9DMas3pLYS8c0VGwlpPsr+vGUl0WDxKvXs9BsWHHW4hNYKy
/y4Hf7kdmDF+8bH5x4XTv9YcfYb38ac/1KBIvjwiDoLc2Tyr0HxtaTNhzlHIsifi
Ds5n5CvIJDa525RIsn4vfLGlPuvTQX//o/RwvNRqfYwATZbDqB+ko6Ma9E5KSNl2
Egf67N50H/1NTgk/EjT4Qtz1ykrI1culLBztfP5WRykUJgemoDBxP+B8sQqybDt9
Si9BhxX7Pf9h6jAX7O8jMKLVRNlUWFvdXT4f5ngFzTApkv+O+58EJkOoYyr8O2Km
+73SnSmarogbAxZJwaXH4Kb7HxttaN1MJxV2dM/O/Hqqg3R4tYon3/H7zq339c6L
yDA4OP0ICtQgY1XfduhHxVcdn3yADWbi/x6S/w1MVCdkxUGLeeQjpmL7Zkp7DuH6
nsaUKspk4DMATTX8eKatwsuvuU/Vk5nARPfiq9FSL4la/cFTbmuUIB8sUyHVJwfr
ipvBOZRMDTApXXPg5qI/OL2DjrAUwHdNzou+vROwy9v5g1q0oLWhkeJM8ekmugmi
vFNk92jwHYqeyS3hWTddlaKAeKBsi0QeumX3FKse6XA7gdzTzoEMPkd12Ijh/mfW
anR2rFC1dYHF6CYwOi8qpEj+d5NU2sZzrT7Vz1eOSSqwTsKiTAaHOkC0SK6gGEng
BsGBj012f0DRIHs+wQ4J1zf+yFPYyc+DhrruXmMn9dMmKR+1Bh97lfeoRjxPjXcl
A1UIK+opyVFKOmq/vJvSLpNvEfhhAdgnUYSs8TW3MF6OXMJbpdOJEN4koTzejHwY
iWVMWZhTcA4EBPQGlEtHm6uvfXkeLmCM81owbzRccxGOKi4VYkdaiqSpe5YQE4u8
oP7xv9QZHgai3fGs8BF5v5iBylWwdO7sle6wTjdXcH1QtYD/5oqBRKRSqyXAr/6W
h5qROm3INJPC5WbDoCVsZGys8FLiTW9Uj92ArQCkl36qqCzD1A7MWe6WsoYwOe1X
VYXGQcKp7j1jwYZGBf3c6vQzZsJJ6hFUtV2/VkirJlTqk9x3kskYsng8gvgYAJHv
oOnUooDe9h+uUtujzPhOz13OmKO5SBrcYZXnZdlJaGO/HXdkX1Yg89N7fn9QIx1f
gGCBP2SslYyIhtdmqynxQaKP4nmfOXSVnZBl8X3RB5IExwBZwTyJImDz4V2Q5kQl
6Ro9HzsF5XVoExXDOJrCNtK3DgzYDI1xMKHtrIcsG5knE9W1Q286A5wD/0y+hArU
hTBgidFeJsnV5zDlI7zoSNvvCuBVDWaBFfcmbTVsEhRsVgYTimpyd8yQFbI9Ji3x
1QwJbnqxe1NZaDOKCgsl0NxYhRQu2M9JEdQuq4lHI7a9rV88lCaRw+d8w5SCSJuw
QbNAG/eC1VrgU+T2WbzEavRMqBzJqNB/6AdAk8uu6wQmqlweEhQ2t/m9BZXZ9P2c
uslg4bXOigmlPwPCr6gPj66q8pMXrTofVrrzGWEDmJqcJIBEpxlEn9VYgvYoZnxa
NWMqgr7B3WnowoIuHt4yduMY5gniII0bzyxypS6QZpK8/sEuCspPNoJZTUGBXJFi
Zob9hbORdlgQOl9FuFf2wqVntcsIukDMOWJqrakgBnWoSBVUfg4vwR9bNwl0ygMn
RuWpvrY/WYE5kVgOQyL4Gim9z2aKTHvEqUs8f9OivupXk8flC+uZOI1x+JzI6ddn
+sR4RqZRJzhI/YqPOCXBxRpMmzZ3PnuPSed+SZbK5gZGr4x6HN7wNTMh9IbanXAC
mYaAm8pFXheWFkh02V7b2e/bpbG7ZG0p87I2r+FitJQUgoZb+UShspXkNRc7qBON
TI4lErOWLM3V7ek4q5a5HcW9As32eLp0fvzDTr1GL4huhaUKOG4EZEDDWyoOED+4
kQPCuacNf5Ed1QV3b00pGx6qUYVUlOJ2y5MhZ/z9+lhEQw5BYKkIoY6ih9psSAAd
g9THS6JuQPW2TzYiR+Me6rwgQqOEHKBpdk8MWKuDaWKdJ47t/hzd9TeoNgrQW/qj
8nTTfdhLXsGuUdTtDxudkshd34tkaZ5COjnEVzpCX1Nk8QXJ/xUcv6p2xln0A5iu
BMS/BWzezxnVKEZVI0ELegmjyt27XtGyReDo1lHx51BvYhp1P7SmHk6ddn15qQKP
2JQlK2L0l4MI2Umi2bFEThJuCXr5r3WogbPn6IvCBQjuXZETAZYOlol8wggjw0gY
STyrBHafb/NggL2udZlG46yXWT/+SU4iYJyFRfMOi8rWFbTxj8ONuqM7A2OxFQ+E
7MM+lMnX2SUlo8mCiw5hUWXQOkJGrxUCMGhmIWXY7LDwhSS02Qn3vdk64qPz/fvm
m403x3JkKElOhws0nPOozjTgBaHjNusH81V+vYRTArxeqrNSIqtLP+04j7DgNoQh
enkjZ6ZNEtTK5R4DKM94Yw/YjCTDFmdzJf6d68Pb9SMEP5uBXiwd/1Fy1CM2UUSP
duwGZuCzOpVNgbXK6p7Cm1iMWQgwpm/8YnM11UoDo3KW4NuT+YgdTZ86OdZjH/sY
MNujMBeb+DcXQxHP2of+nXlRzAYZ/52Ee1JNOR+Wjzt8IF/EyU4uz9Ed8N8c9R0o
rSxCeH7hRLdToXhX1HS1l1kSgl3xGCnQ1l73tq1vMoZuXrqZiA5mfEPo+UEcRZdK
s1MEtRtq0VG2z9R11AQyPLO9eP/b2qr0acIDXI4Cy3lzXvBiQgWym8KtZan+kWfc
gnuD38lDFBSeT3YsHXW/l5Z+o9+p9NxUT4KY0Ldgt3vRBw7THx6gd4oEmF2mNytO
pXS/UkXWaXaGs/buFRmy1R/pvHtCZuVFYsVSBEY/bw+U/hwJ5uwfgQeRaGuClVwE
KZlT6VN8py+ac84H7QubUTRj8TMUM3YEtCM5BLEBr3T5Xfs4pCsfHft5ZkXsfaTE
b7vlzWWi6MN9kNhNNM0O7aBL4cJPAVKaYv8tLVjPG7/5XmndxmPBb8/VF8L5C8Wd
yRXnmh4HS9zqn9voJHCKfBSa2GENqKRXOOcIyGw+J9XhonNHDUkgiWb2iPrcKbau
fjUIfGEPdbAAJh7y+bQziQs92IIiACEspY3tY74FrGWaaV6u+L+c+Irj51RZrWpw
mCDdpFBN69rTJdpw4GUGyB4HD3ABVsNKApTeD1784B/1NWCeuquw5y6E7KRULq14
R11atWeFzd0EGeFafqNzxu1rfH7tI4RMWTdjGWe6CNfZpeemY32tm6Sg5IzSyCLO
HWoLM6wf7Ge/oGWACoviTMFgrvP1MojcgW4oOxjA48TAjxsGrscJMRwbStLLBMbL
nVaao+kq9S2TOTfBt4LHjTi6vJKIQBxNesdyK1BEo3vNyZCM2Njkabq4GS1mxW3w
eQEeHNjQl30rCEaRlDaTifi0nsGiUcoKy+PQJ5KphOMUA5M+2vZjzK0YTeM01Nuc
oMlTSnUkPa/hrNORofpsil8EpzwSZwRoHGFTa+MjXPvdvSSBHhK30cYXGFNaz+bg
enupTD5qVAMaP8N3jjTW1YvmsCt9/YqpSK2a4kOnJUMmRWkGdPSAUs1XfQEFzHI9
/FAIFB7LducoC4wPtCYb49+D06FQup+uYJFjifBn5IFA/JwFEbFPeUCqvYimUScb
amANLpbdCwUaOzHu4EIK77bY5DkxBnotaw0Vd6ZeHKlyOoe+6sHkca83ViLFKRvf
76dLXjP8K9KFCJa0K+R2uiyWeYDPZTC82BDvn0tvp+a1IrhhsW58u5DkqMxyZmkA
Wi14gcm3vfBwlo17J2TnHKWZ9ApIHnM77a2D4rgg8TQfurJW7de+gK/6/95Ejtfi
xJi+Q8AjTyLPlqrT4xLGDG9XOQjJbeERc9EnXuMMkX+2j19Tw/fZ5/9YaLSUt2q5
c2HsNzpqlIFsEJk/wUr3oI7sY4bveB+qanO7IEbTUVoOLwvzzZhsYtx2TIrh1m4r
C4c+x9BygO9TP/qneRBDY3DCEKpulQRoJD7OF0o184vDl2udvKcHqRfHMNOW/i/q
uVdPZVsxXrGH15ovDdINlfMGqHO1afAgUuFe8c9BFAFNGwTEPykVSGu2/dXs0njo
zNVPk9TVj/adN4pQZeYUM1SiVnzznwqjInVcSx3lbJsXhzSwu2q5QqU+Ipm+vF/T
ZWa9iQ/zuw8d/cWnQ2NVud2CAMNVG7VNwziRXc5QuzbK3gWVK3DYE79KH+vGxoZT
rIZz3/QZNYvo8wSU8CjMJ9CKKG4YIpo4tz+A3JHqDEDHaD+AD1l2w7CqzmPTbuvv
B1mlEjOL71OLAFF8+CNj06dd5jwNCAps4AhC82fyCY060qmwIZfnG4ohvOptI44u
ccCH56IlYu1ZbX7l5+0d2nKr5pzsEucnHqh9+aErllfnU0kHSuQd5oTq2PQ1YhMe
4Tj04BjDE8D+nS9E0GCYjpXyfEkIyEw2wotBgW8EP2UG25tMg2WvdfZ5f8V2WLnf
ro3DzTqJOgYeL6Dm64sn3mdz9zdP137npQ0Kfj4nmgHQzAYhvxPhP+SRVYz5PDLF
32KRUiz/WvjIJsf9gmyiQ9UKNL0NPNtbAsOaYWeKlw9MDCZPSJ9qXNQks7wtMCU7
SdvWXgj9BpzXroltlAfMZOa1+lA6LN2Gs1jO61EwWMhARbcRmKvYFK12ccaYA7HV
dQQXh+Y9qJA+Jv3lXJOog0dvegq8TZ7nki+68jpRB1okLFO0eaem6F3pmXQ9zcot
VvPwlQtoE+CivaiKtssDezj9CKNxJoDb6V6MFGgbGdehbtH0TRP0yaYo/+C6tyaN
FRtG+f9oclw6VuNjvJvWSQaFVQ81rF3YSM9CO5p62MKGtdEr0GlJfx1mpSHV4YFr
qNpPYax2p+sXShr1ppy7qo+NSqHLLJvE8phPlryLVOwoPUkTiOJ03dAJMh90ac2d
a0E8Qy1ZbUeV1n/mpoH3CGnPQAE4PNMkK0M7JSYGvKOISyBA/yBtbHjBbFiVGTt1
vddzn3AErhZ9Sir5zjNIqtt3VjXEhdsmQ0FX/3Z/zrQB25vAmQ/HYU+FhgHq0qkl
VzSi8Jy9/ogm9swP+AloRW61com+0jIIKvXy3TElaOnrelGiGns0+FWbryYrr6xH
swcZDbKvs5Gc9UEC+cNsGgAGdUW6/Iv7db/r4qqiqYkjd/XMuqQNpRBQqbO4tUbf
OT0vfQnNP1KWYmgTMsV1LIwYy4jg6xw8YcHpH39fd/Ui8btk2cKR0CG45/7n16PF
XjTIiLst57Lgx2fNWk1Iy3tCgGGNpLkyMAFZyKnywRhmFQTTrMWOPDgnnlWAvQ3k
G8Z82rp2jd6xYucxhihGdjjsDlA9PBDrux2qyJKZJDRfolGFOZbSAXwCXrDUURiY
UojQGBAL2p6F4VNfqQ6Iczqriq5FkoPQQa55M3rkLCZyLsz43T9k/39EL9OtGSYA
5NjdpowTh+1zvGTTjabVeDopECvxgm9JottZ5VxgN04aKi4KsnVGgpmHj8XBT71W
PWoO0EBYmMIqvfb6YiAo9mYlB1PZytV9KiQoOGKCvDbOIPst4U3neSUZczIedR3m
shEZtsUL6/HfiRCtbjCQmeZdhxG45nJTNV+ke22hTtSOdDh9uk5z0OISGhEWOoCD
Visg9HjSsfIy8QzKj5MbrxcD4Rr1UlvMy6d/cKjluI1e/toB4aEMy9h6HpUZ7qqG
0DsExHWRLW62EzmvPwRU//PD63QgzAHZNi2N25g28LIos/OCGlouNHKObnvfG7YR
a3i/euITuf20LClxQcnF1uJgmSI/Stpc201dU2MZWdYZHyKRd92/zxB4s2V0+wVb
VQDq7+qMClwHx60Af5y9Zo87nUK5zfKVTI9euo2BZ2gmrA9nqeMFb7wq2hJ6Vxo4
LbP8CgXeaQHfHgumHADnL+H+VRYNb04ZiEQeSzH4U70rSEiK/o4uoAJg12tgCiFl
rz5VWrVDNpAiQlFDQLv7quwLPucsUL7s2mj8jX1dwiUV0KP3aCvf/SOMU4IVU/gk
gh8CQ4aTAwylhQxF1lPWjL2/qEPDlgTHj2HE60XB0/Z7ytPnZcBekatwKWgn+s0D
1wKsu4xEcag4c9Xc51TAiCXzlAI7qT6ieAWoAMC24BvZnLx0iqsWBfRm3H2efA+A
gs8FSWaeGcYw8AcJQK120tf2XHK4rsylQ1c/qVjkPKB/2WOTISS87VYlL7cD6tyu
wKxaMhyM6krR8ZyvGNuJwUF6/MLviclDWPQx//n4Emr+Qjfba4Xoga9fZZAPMQTK
cggf8RpTS0WC6yE9UrZ3Bfr0qUOKqOagallTQKmwYPSrXSMpq3mHaAYU4ciZc7Oc
Wn2K4uHV+RSTfFA3uR9fm9zUOcu4yNWPsbQ0VdesJ4eSlYRmgYvJThd+w0P2RXpr
3TQNuw3dHJh2xYgxzG5qqBfKlo4U/EmgW7B6k/V0zlbTKV3xS/x8T4kH13WKPLo+
FD7nWpRqe+SoH4/dFzWtTf000CseB0YPXpKrgiohOPGEi3QZ2c1BZaJBm+xiZMF5
0c8LWfjYXJiGuUei1c/ZOaB3EKFyNFphHaOyGX628FnbJH1t1ZwoRUupc6Z3Zejo
qTNlW5jzzpR25qzYaNTy7F4biXLDMgnom1hmRfKL85GX1gLtzsZs5Ze3XDXMLpeV
AKUPJ2fBTuX/ceorAh75N0rBDe/d1H8b/O4Ioi3r2lkLFBi2oo9vb4x8BWv938mB
f3pGaqTrKDiYZFose+VpMKudyN0A9nuq1TI4BfhpWN3FdFgW/CX3CWdzgHhtochw
Xt1ONyppnBnwW0F8bRgTEnjvc0oHnb3f2yTM1QB4HPCT0lULLtJRfWA69Lac88Q8
mUiBJGqae+ndvLIF4gZQ6KrheraUGd0IOhfH6YEH0qHg3AWTb47BEm+M/43losI6
SEY/2ksev613BBTb6UkHTcTVXX0p939bsn6ntoH9dVWq3OodnnQ2gGNfPfKcVYxj
ZFAevIQ9mKlqzZwV4r8bf0t9Tqt6hA8zkRkWRNHK54Xr9W2wbUXmA021XzgjnkYR
B9XWAWj+WFQnJ2ic2c2Wj0oDW33JqtlOtWGY+dUtSzno57QkuI99ncrdooE91Vu9
pVgQyElTnJrsuvO3z7VaITt0RnJAlZhMPp/r8HQslhkmTn0FkoRU1pMrFa8pwZYv
ZeKk9MorNxI7p8Vwbiv79l2ypJMKKpFHf6GGAdwk+JaW27/7NKJjTbKnSiQCQmze
gOBoAFdppcsGjz1OWvTq1ZqfML+h9Rg4ucgnQQXGfp52qmoWNKh8nxM3Wr3z6eZG
MSPSfGlr17xFDi5yoWdcDufQtFYf7Nb8+/72p6by7aI2j2jkhxAU+LUzkYzq6iY3
fmYE2PjFd9D04jlwfGzGMRp1cN3pTGiiN1CdTqXXm/5PvVPYWM6yEee3Nox1l5u3
6UXQa1LIpMQzLAQFCiI0PxfQK8kZ6Ci0Exj4anq705o1rA/vI9/rp+3XMhOyzPdo
75d83TM9zE9S7aS5H/CNpIxbw8gtP2VW2tS2BVYXw0iZnmBTkROtW5uSa92xp7ny
lC6XeFcq39UtFRKtzmybaJhlLn/5hYnqucBQqK3Jl8mKjsvdVdKDrpUwaC2Vg8pO
BrUjq8gOPFtXwNPtHZjXvbSj1O1iYifaD8J3prlLEF2kheNczn1EC89+7GshZYqB
KoGvcHTOKgYNUTjMzJWd6ospKWawBflHTlcn2tqtF1zIbu9kKFejKXgpQCEX/Uv+
JI0inOtheXiU8eVjxyv/5k+TNDQdR2WosROabjBIepFLeNO6rhcisinNpXsycLgt
x84i9aGEcgNjK3oBnWH1blpBmyKxsAAcXrRWQkl8YQhRe9Kbxeh3aSWQWip9rA3H
JQytW+fpsItRALU7yK94loi3tAhetgQKZj2+pVr9a8SP1p/lwRkxGANCS2arQhT1
iN0gZwDTwYKf2/JSD+Ptgewp4rewBTD+S+rGMEo2ztuA5yZsJ8HTzfF2uiEvdAwA
tmyelSqVOIln3KN2TUjII8D3WOKORqRK83CIoWHgSUdUSyBL5mTlcdse18cjMlFy
/eUDoozH5dII/wSwx1OXUFF2RVP5YUuSEifZbOeoz3OvmB7EGR64aOSaWcOtL6XG
m3oZ6oEsRkEHj/0ZkCERLozoJS0xfcyU4mtkaGT54qIH8NHPAgXhHR1M4HH1UEZC
Fi9UgNHzvfAj1j1+H6F5tX48YDUgl9EXK7BS8mqiLyF0zICVaZKQJ5MmThe5huqY
unjP6ucCwba6ZLSSTPbS0PvnFQji52/xxPwLIxhLiCn4zsXNaghQip6jIP1AI3Ms
ZvSYQiBIhibxvOUrAzMIoVkTqr24ORKqQg2EdDkNzebIgLNbOwHIUf7+d9q7cqyI
i7XnCtjkSeBfYaWAXnAf/oZilA/pA/c8ZLEn9K/Kex68myVI8uSDRJjIWOoO5p0A
7tYwDi0RQlXkZane/9fkXNcTL65R3bHtiR1YnWQXlBj6P5NbyxW6ZtxrOJWrF4aD
bS0R7utl7QQASmpfVsLQbLF2FNTkLdVhKM+eXXepZvLFZpGszB433XAzbhqROfrB
UFOcnWHg/zWZL3FozR7utGN9V9Ra0AzhLvTlIC6TxqweXW+GkB8EVysk74KNuD7Q
`protect end_protected