`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11040 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMWORzZC7bo0toZS2Zods6Xs
yljw+BvqICQb54hGe2JGpBpbsgrlUz60qXw5n7sklfD02cg8zmM0F57jsxk8iaTC
SUfZYBylCx4/riR/9qEv18cNz5O3Eb13hGxOFCzG2de+p9kcXgrEPlaeZjc8ykXO
YxNstnyESvRYXGP5rq7ez1sjiZx6t1A4h6RUdDBkWGcYlWB5saxgSUhn5rBenKN8
6saPacXwClFPjSzOaq5R/pNxFruiQIMqBtVQH8dLQUV+Uro4eFdlu5FH/1KO2Pdr
LI8KzHILAUvuzcS1YC/rdpEOskfToGanv0WBZGQegZuEBV66e5CrIO979F+skNGu
HHfUAIrKKVdTc+eMUawFWis1F/04+DpR4yK+eUZpBXL47YNBqXlvrtLkmoqCaqWl
fhFcNqoeJR2qIcWIWUL9K9oX41+651CWD/vZdU/CdrXYKuIpzsWldlrTsVnjqqmO
Y+c9UtWp47Q0qpBnBSelDj5fCoCs3VBz5NYq46h+Semer7UcQ8jfD1p74zN4G7yO
8yE74Dntn0AKctbFDZY24mh/vuDYAdzXKs1IubKCcbPqdahp0HecgrpZDQyVzd/w
F7S2e4Pf01HX3HqhnA0xUgSU4b2/2FyS5U9CjYU+6HDh0E3H40MzYKJtsiwN6wOQ
dnSiLsD7NepPxqIZDVRwIUHxnYXj0O2mBbNHDKm+cdFvkaYcxqRej2QXY/GJQMox
LkLdLU2u1m6u2GclzeUmnHJzbL9m9FuZ7s7hUIUcNmR50clbAZYklFy5I6x83w12
eFEudnyX2kTVaVVFSFxv2SuwwvzDLrWp4DtDu/QhvcdzSnBbjl8xco1cdWin7sU1
qE33K+SvsHmLSc/WnbgoSI2P+elv1mKh2LirzZG8xOX7cWJ+TkBrEVmzx9F1Mdaj
l7zi9epjLmkMJSCsXql5nOtNq5aT3D/OtaZXccZgmpQ35y4Dig4ermNsMpeEjy4i
ZDzfUDclWHDJRQMx6zD4GC0hsQIJEpRsMc2zqgp+vRgeBVz1ua/aZVX0VbBYeUjW
uDkRfrI7u5T8Jk1bxhPe9f254A5QZd1GUAgah82CqPm0BcR4i0DyrbJvjWxUyKoa
ABKqxm6WkSpeSKiGSlKbjqBSKZrwrUgBymMxj17wVLM2yRi37D5dB86so4Dj3NXi
0ZBYVf3gG1xgHYucecbxl05XrpoBfrA43ET1TY6g4CKIO1vM5zKgCEOhNm0YHfAu
TGbqdtZ/+W7HctH+bAoiXCClmOUYbZHFOvGZbaNZIeZDQMBvmEPfDan8ggFSazna
YgnDQrUy3PQFhs10PZvw855Wn1wVmeDN6O5u4Zw7uABdsP0OwPPe2Z00Hw0Bt0fV
ypovV1AanhxoM8sLyr9Bv94SQ9Htt6coHSe9ZNV28RRQhClIPwnw1MILJBMZ3Wzo
T3m/lXrSGR4T4hK25fcCG/2HezT3j2nUfdZPfQVxHzvDpW/5BYbuYAuhFWdu55xB
81hlxHzUqC5m3wuqtwJAlGiPnAWCIAKmXLiRm7mZIDFD4gPz9B6SFjEhkhDMkjVD
IM+xaPdn/LwWqKcLyYpk7jDnF+d/9vS4NczSRY3dgO7xaOoFTR84CqGOZHAAeAqe
ZTbOu6oWReWnVLsPd9dk7bmkPd1q+1EY4otjnzAHiw2T83BGGk9xUyF212jnf+yu
1ReG2cQKjKKDjqtP4pBoyEK+zM72eAfdw8CTHfdoS3jbqGPM5PR78cLKKKA4IIbP
o4MM9ozmfGtgn3voU1sNp1znJSVinOeIapCsz46KMY/l49h+IGUtMHb6y26ISwnv
8GLrBhopMLrYC7i2/HL1KG12L2G9GxSJgJeZvL5+PxEi8sfLFt8uqcqZnZjSkT3e
r3RcsIy/EjAR0/EJNOQaQ71qwwfWwu1fwjfqr4ksLixXmAL45xinv8GOr2sij87i
FGpRvzO93Omn1k3vdFs3h43ikFREjWv1VrTNNsmZInPr6MrRT65d+md5g/1dEiRc
zWmjuo53wPNH6VWiMCXQBk/MY00LOTD5YPfhhRVTCzgbOgekmLv2wa5zfE0BGv/Z
g6Stm8j4SXiV30v1jRzxfN0X7C8VJibHZ2SB4TJ5MFOjoAg7hkQKYj2udG50pSvg
4xqNKPFb0voXvvClbcqH1KY1BiGz8y5wX5trkPL8quvU9VnSsNMQENujK33chW/0
1tdhvMW4dqW91/Jb9LBJwMUlwa5p4wj29GUMYouYviJjkpEoP1+oXNilGXqLoPT+
87XaN+Ol1NOmlllN1QBuKXp3/KVDzR4oMtiIgAv2mM3gOqhqJp5+Ks2kftMTKRQi
0Pba/ucAVu1aMh7l4erHHpZXrdoCJxaFB9F1hH6leBIy+ai1C2kt+VBf7woQ+an+
cTieFGXS0vBdc02+hCibSGZWTHMtD62u6MBWrDLtNvqKLZLaS5BR7QaLb/mVvXBV
32N0A3OZEd+2W2ieeloG/Tmpe5TkPCwH1S4zmQXWu0wFFamD/h8JzIu7mp0/4kp0
9ShPUVdBdYTN59oTeHwApQnRrKs0/EYA41yERTOV8bH7mVld+ct1T3I88u6H661v
qmnLs+4NPMCaSJUoPg6doVevyqRiUe0rByYU903LbVilD878ptisDJQbXaS1skiF
Fc4bBsinoj5VXTan6zLlI86HQWhwh3I3+ZhbJAhQLBrISoa4CxoW/xbz9QinmHMv
vDUeQtDrBtDa3OYku2KU4eh1rgTf7baeouS6RcUZj9HVnwsKkzCcGPCpuGE2LW3d
VtkrUkHnx+A+w0334xtfHjCk+NeD5czrVQyQPfHrJ9qSbpk6kI1Sa/b7RoNb9UrX
bGNM/1yY/sIwENITlcvBSpD0Ov0ZkGY8WyPfsPSCvdw7NKqZn8f+E67cv0YBUEcZ
LdSxkylUfD1QFwiO3WvnP6ybP33cwB/iXYOaUM1V2PDwvmsNVFjpGQ1TUDpNXA2T
pvc0TwHiktT2l4k/b9K3E528ioy8ZeVVJPpdzizek0ExGFjQv/dOvZq9VRl6XRMN
76hw+0hDyuMK9I18GeJTa9hDvyXqGmLbGBPMgy9QdeurNyo1LU1AXRnsx5Z9AMj7
hnhoBBR78q1OS1n8d1CcmxpkKOz459mRCqeeV1FcgE8ZYDutLWPSbSyI1ZlfLkK8
YNiedfMPzLI21qEXyTrr4IqNWgzmloJ7TP3XBJdieiPb6odEnaNRxZ2ToQ/RAADw
jojWDoGXdai5rsRzdCTDiE487KlREHwKnORszwBJsy4E0EbiZyz6u8TlF4L/Iv4i
q08AaFji1lHswYVlpYCRvVT+nT6qmgRydxrs+PIhAyZieOpCE3m2/KMldbSK6r5n
Db7ByQxLocN9Ov7d6rVtnKqjM4quBNwLDRL5yK67xUYBFuPXBx4LllPIPOdOPKX0
hNvbjMlAcP8mA/9juzvIm+zQ2TAKZomUBI2kWlqXGmmZY/2iQRHiqwPB2lY8hgET
p5Qk3Q8o0cAkZO16dDp/aJqiTqedZWHd0mmAtKYqV7xNibrNGVPniKl6cBSlfKTi
QibnHDs0+9gAvzy+lRg6PnvjpNy2rnAiS0M1LgG2jb6pJWqkvrTcIZx4313VT/up
qH/do5Xw1CfyUEBdFEFNKOVVJUl9a9W0o7XRZiu1cD3akWmluTr/B6TCFZv5eql9
A8f8Z2xgNCEp+j+xW84xZ6VG9e51PJV4HGSt8PbyMv+h0B4jaiqBqJCj12+zj9la
D9w+YnebGJTttBFJsWnw8Kdh+QIvnwOWAkzVI5vzhtmxlVPlsEvZru3ecXm10g+u
i9QQ3COOVY7lJOHccn58BkP2L2lY6M9RB8E2PpPPkoSHl7usrPwuftoZ3nm92qo3
8UWCTXHGmPJRNO616pr7TFxwhYOdwfj3MHjDeX4Nmrc0oa31LuGpNzB/bFt9R1kB
ZbICvipGkQI46gzzELCuH1hIkAm3Z7vuxyWKLMWBq+2QIWfulfOMskPm+A6Ju7Mr
B0EJ2mZCUyyUCo1r0p6h8etic2sozG0Az0CiTGCjDgpMIAfb7KjliMC3FSTdLkiP
64UWL4/RGZJ3w3qlU604M/Zsqme4wQHoX1Q/OIpdyYJWFDZCmLTJzvSGRtevWmY0
7kZRpFeJOvXR7GBpC2t7Rj3CiSeBHzo2sQAsrPjZfMrBSpGtCSfp55kzPCvNOF2+
jEAJUw2DEFmItYtHnMa44m5XoYoJyupt4KvwF9sP+0vhdE6/mMqzTgTmdCwFIdGq
7INp/U4SCxbk+UigFJmOvgV8S43mt6kbo0HoeQYkognzwwCBfpkoPLJ1EYEbIPzp
vPqKHUPegeDzulcVw19BRqoyXSgDc/zAZWnGO7SCbQaI1l+JB+LjoYX6vQaUWUgb
ttpFqV675op2tfotj9/tA+lm58dP9YagA3a0zFEcQLF6Dd1PNkqYQZ5aj2PBhkD/
nipwsvVHmO1SzMRHDMCMEWhIe8PMuq4pHZJ8f3TbDzICV4RqfM8LjfIhpUgl+sF8
YaPPOPbhzsyGDmybbEz7QSU1WvuxDNdh8QTSf02ND7rdtTKbKuo02LEoXdPBcMDn
QkohYseqAR/1O2s9d0zQr54CxQveu9S7XAXbeDYbmR6vULZmfucgmzXHwABqVW0+
3pNdGh0dujVQ+VQewqmpvfrazdcwwQZq9dlMwTRKP/S/Xw6cBjSTvGWZLjPnHr72
E6b2M4f+EX7/iX4nGAOcWBH13/0rvRPRQrc/E+EC21p1YRCPd/uzkAKsdFkmpTgK
MqjHnI888cqP/gyCdGFkg4eUMOoVUmwgftNn4u5uhXGCHOoFgY1rTeutnRrPygQY
pWbSUztkk1KIhJ30EW9FuZ2p4o5l67PzqnYod52INxuu2tUHYPKwqSqKJsKT2G/q
2dv+R+mUck6arUNM/Y5vEICIDQMUIrRQQHuR/ELVsK0bMFxKFkPTUSMFS5OboU0E
4/Cxu5qXNIta25az2HSp8gzCjcpwRzLceQL5bbsfWU7E6Jo12T4a8xuBYWEgj74w
YoDQUMCr6ACPno5hvl2aUDf/x9yCaH10oLZ4m52mpFAkLjLKacK3mcMI87E1LIP4
dlwB4pQ+H0dwaqOLoE2+eewCai3pH3PHB4xY+Ox2WYOhziUahsI0FwLGZnij65QE
eS8n6CWvWXIwSVDYkIOEyl9oUz0eQI3KfbOJZmnmQbnYue6O/hyEk6wBjdRSsd6f
f5jSz75KzFoI4OaWbNeIW+pChC1ZZqksMxTfgsM6er11Y7we00mjMO86Srx6YeFy
QaRAT7Hz3B7bh4MgCsBKiW1hfWzUgBFAi/s/ljYnX362SdcvEd5w+DeV8UjAtFWX
mQ5CXe2bl6eVLmWrYJd0NhIJ998oUYMlth4UBlrTmdZ2jU7ZmK8XvG2fEUlSygR3
tgdwqr9Dg5T6vbxJhAe03XOlW+n09t3SIL1tOkXmsLOg/gi3TJP9CTkjvFUqM4hb
CbyYAHREGL2unbJSxbxcz3lH2v8PNUBdsXzk+DCi+J6ykmOlUhPtlRlWwMxn8uhR
2uf/i/SIlPCgnmqSjWVuW/hnu6uL72SFbF1XU74+qY16X+T7jf+2vPnVzfpEfFgr
tI7yHZKUO/wRSwbdKHcqU+1KiOa2SGJx8OgluGa67JfwDopuk69YsQxJCw6QSznY
+xF/QhjpYz3ETZ8fQ74jrcmQn0183Hdk9VFIPwl9bdKIDokVrgC77iclbTU5sB10
ioYTKrLaDE8efw0p/zc+IfQakGrVAaoUSluTwtCfnBRC9HF6aSNE7jOnqophsP4Y
hyJGFesC1eQZzE/EaN3Ou5beuO8WXmQqRx5WYVxaLwt5vyTfBD351353AT2P1WEJ
4tRo6wAlrhD1y9X9oV6BhqFzWkC/ChGZKR0Yt+UY+VfgPEJvxWihgs+gS97p2tfx
DqQVkTzLd7+WCVSDEqzW4Tu6F38Qu78cWd+jopueSCmiyUj9790R9X8kR+Ej3ebS
+kz4Sq8XtWhCXWzeMJ7JXh8rVcuy2ZZH/scYnDqKzvlJKYhdomnV2Pyz+XXxfIk3
yYS5sgVtxUQwd68iFhNyvo+5gffGZCNu7tmBh8QyrBYAsClYgIYDunKdnH7WffBA
og5lVtI3PaqkfiVHR2ss8ytJF/clXVrVH+rqarVeTo30Ja+gBqh1uraI56EnWEnW
cOKcWodRTso0LRxy3naJf00k3qVhPaE3iCvRqGsFoTDE1PYpbfNNib0iyvS82n/2
itIG9WhIWszlySer7TLNY6KHnP0n9R28lnTMMUq8qprGPr6qHTA9B7Goy7Sl/y3E
P5wHs68TMcWbK1owNxkt3pCa3EfXHdPBTq+Ks9+MGZJ4ZFfZYbIpVbTCM6mj/B8V
qVHt4uGWgt4OP9taKSJ+78OAOVeDrSB/EADi2DOmu1pS2w64CPhrjhC/AXM9/h3x
D7s42F5Ncvv0kBBebBt/TZrHQ7OOpp0pcnbT3y7S8r6llS/I4XuhoUgzCfMjORl0
wcbD5pDIGijI07oBKbucO9cM7B2uETCncZeTsqJ42jR9o6HSz9IrNKijtHw/Q7lR
XDcswhLvPr+yY3r7uNsqBkaLHgBa/RJfYiB/wdKFoBLvmFdTSGCgJOykLXjthxfV
25Hl3pZ1eDWtEOdFvdHFQHSOBvmnNi+BZQGtzbbyu0IbuqLpDDsqykIBuXl5UlwV
c6YFbeonIfvPKVt/TYjdZ1SAZ/yY2+SLM+r9NsRgaGEZwrB8EZtaOmUm4iUTAZTH
PVmkcSWgjcuWBzS4y1f6LmRywlwe8cHZbgh3si+k8Sy+mLBG6wFvRbtvtfnt1Jfa
5x7UwRKaLeHT6C2epCoKTtjpSGKH+KpvldjU2rGnG1WrIU/CUnoy8m4oftvyz2xg
UHS2RZ4S9UWfdU/iqZ+irrt0fZ6aQ5ZddEiCurHoqfHazdjXeTPM2TIQIaa+l+hS
hq6Ak6ru5eNSI9prf0ujH6ZliWUntn1cK48mFMIdIRGdecsSJzmNKxFxa/MgQ7lJ
llTAUUS+j/fIphjQlnp4wTX18TJtyZukEjfQalje/L1P88gg3d/Dl44S8uteDWF+
dpbTzVAWwQq2XZBPOTio/LIvYhtgp8t9ZoZ7U55ZwaPvgt9iPRLGhX0lucjdm/MG
ATDM3wRclrmtN1z084nLclz1O+rmvzoUq+SdgVjsrxNqwh6CbQTp0nxtDK7mIxmu
wiJZu6/TYDswCJwCckivzaULgSrd6BvLoVyxo2nQlDI/hy3OtQN0t2WhcDULDFqC
Yh093RrRJ6KbLtWSNiGcLg2ZzeAhOEYwGug7IjSPQcHkYA7ER00h81euIXcDC5mb
bFiO9AX9LMnsLd91yQo1zk9W7ca0NSKVD1jMpWDNJCTnnpufXNCMTbjR38tSaiOz
z+fQoTaYDcj7xkNOwbGxoGXmjHLYMBK4FdRi7JXTPgaeo3soZ1mxqDSBSrR9PdY7
6Td1MT6x+t6NZneYlm8i38T0ZuT8Ombh8aOt6Gq8pP/abAkKYOZii8+mTyy6Ntrk
XZ1F9rst65L198McCtr/gA025H58rc33yVp++1vtFAopHo6gCrwpeW7haYAmOkox
HYhdIf9t/5BKiGOnopYkKNk1vJwBtazNBvlgaxRh5xRd49cJRnZyiHW8IaxwgJ7P
QoAQCxDF1yIahpdRDqs3Jf0bKOeEFpZ8gIMQbTEnqd5/blUOnA626y0fZKt+IRiI
eUQT3bW/TL0+0wCgBb2kaRQwKKbI/psak9Z67aZW46NUcaWrIudEhAreJIYxl1u+
U9OZii9Dd20dKyqo5p4wuVjCrHq3W9O1lYmiE0nvKk7gEC9mh5hmCa7ntgOZdCNA
gNXwbzSmcwd9Y7qUbWI0CR0BAGApSA4P2ajQokL/KFEWflNCxYytGbuJ1Y7AKc85
zX3JKuHpn/hhW/h7X7qDjjcxLVU0eviqzKR+gCfx6h8sAUNnCUuVVmiK2qLMB5pY
+XAx7AKlTFer2Yc7E3JqF9EwzmiJHBAQxKsLWuCF5OljyXeV/jbSzuMv+30SQesj
ahmXbRnX0KP4JYuTVWyTOqoaq3b6uuUQGUn6Wbstk6CQtfnHZ4kxLI3PiNmgC75e
QaG35IdJXN8PMCAIr/cevhnbyl05T5KTgokupcnyfFbIP6rT03CkAO7ElCUzAPyF
8IzaWgQF7dGbKOVPxXyCNMoopW33YWC9SIA6nBcMOQxxz/ZCPN+KPvggGf3PmgUE
exwjwF6T0Ii46aDeNHJC3krrnI+ddGaHoy7DIxjQ8WmPtvcLtG/jbQqxdvjIDXtQ
+pQq85dzJ/b7PlL6YL2F3/KME6zX/nVpLTgxp2DjhgZ2Zd0wKhc4m6fbUhDzfizq
+HYf8VFOGjpyG/bWqj+OrqZN10uPpo+js3nE/KgFvGYm0/Yl1bTlLT5XrCoY0rtY
WRW+qrGBvzXo0hx+qDN+BbJlw5LLG25QczZH8h2rSpZ6i2VRPME2l9SPZRJwRupG
o1Kybzi5Xpfswf4kx+wZpyDS9kRPHsWPnX5xM1QpiS04trSb4ykvu/9bjO2APuW+
ZMIvdqC0RwvTvRCoSgS6lhuGKipYLvsWnWsPVc20+D+1NyLk4AWUB0sEAjHCQXRi
Ba3bNf5sFC1m3TZPXaKVgrWdQ90fZPWHsEv2OjW4yynvwDlKiTygnbPDk8bGKPwJ
TCkRqkRJuaCg6UIZ6B4x1a7RomnfGgh880UnmcY9if61s+2GwYSJik6kbBN/xQnr
BYuC2482RhyEM7qIJi308cOgxMJZmLCP+7ArHLFeevCfJBI2iNrIb2uJaoypCs3q
9FjQIfn2IBQtefCzdfKeXDHmIX+KUOUMGXPVYjLx0isrrmWPgCqwIdfpstbDHW9z
PGSc0kkAh3GnO0f250jsvikR6CL5AL+6Qp1aia/a4mMemyA1XejjCNmBNI2Qfi7/
0PSfRTuSDxeLoFN7qOXDMC4XJfUyE/Kqgyop4k5h8WRBzURhz2tDFcXex0wv0Roe
zfqmy5tfNmA/sntv2FP9o5O57N+4lSKYPgbTPc9lmMQUkyF7+2izB2fah5egjfyo
FRjIyoPQUXBo3SWq6KYPZQa4SIduMyssd89Iynn8snsEbO0b42CiNBiKcbm5ubmN
VfdQO9HFJ6MOrep7GfKd8CigV05kkkDJxkuYWckJ1F/CZgvJxlDkvLxV2Mc24/oP
DlxQe31/VRZ5qx7BQZ9LVLjpvJLCp4xv8tbpQzl9JYUscNWqaRU66TsY+Cbzy8WQ
Jhq3ks5duS8dIkDq1an8lBRR6vF3tiug1gm8FjPiBWlLFumpcPnkHeddRcpT8srN
CXkS2bfB4duiAu3qVMWSYRtv6vyJQYLjRQFOV+pZ6IywVwi5t8nxq2bjvQIC2IcO
4MrK2A/13s9k2sCYC50JqFq819uMqgI5RuE4nEbV2HxPQJWWlRDPq55NhOEWEitq
lZHrKaz24IpJczccUwze5014hQe3PjAJps+J1h3PvNwDsRA1DBMBi19uI9usvQT1
tHhkW8FRb6C2j3aW60tl8PfGwRH7MgfzSh0xbtSgxRli1T4jLjK5lkG49J9pkkaR
vbQP/+2MbXNSaOfY7G6nCs3uKLp544whew9Xpy1D0s6rqNjNyD8y47NW+LP5Rrhg
fKirvfz6hngNyw13iwtxy8QDwkeePVHzYuoeI9Qn5Ktj1Rx4beplsGHEUotx7/Vf
0QEMecqyienUxQB7ytwEes6l9vSwU3N8EJU16iybapxsI70MvRVuPe2kQzWNxlGA
8ZtFBhM4hSnc/V5zhzEdGAqLuxLv3nWQiPAuFWt3MBRtnJ8cD3T654bppaydHdxw
U26jYyemSHh2zjNCeoPIMND204qmwpmnQucw4d57dSRpwOL/R1lMy5jDh3SP0N57
yvZSIFuSLXDCsFb73OdZpRZepO8HV/EwO2Q2u7c2Cy6cBEXEQ2+I2KWNyqUkHw9X
GRKvLHHMkSekA0lbBw4pqSyZ43NWpOZT23okqWbUUSA5azP+VfZoqzS2Bz4/STF3
YCEGciJp+Z8DT+QTxVixkTqQC8O0SgFWf8Lar3ts0U/FddoguZh7s6gXG75zbi0G
bFg7s5KH3rMzacqZiUKyKCk43XZPlZ6mqVD+XkbtEzaTr+D4SYbOzL8hjKaGkIDR
05jHrkJ1I9CWuEDBDCwHECuuGn79O9HUZgkDp8HQtr0E8sNA7xJ3pzUbPiUhmSIq
g1XCaaE9ZQEUBox2jqcWP2hyFCYI47H1+gn0xWLaQndo3WMbXyiyYKBQ304P5wLL
De0fwEIo1XZ+sVkj6g9i1ExXk+9XEL9cpRmdG/05q+7jI9Qk9FvG5gNl/PObl25L
xpRidEh5l3jIFggSA7tqQo9SX7KQn/mlS18fJSdb3cFh6PCjQnYFKH55r/taOCvi
uh2pwmhI/QETGktzD54LltksiJRbC6iMf4hwIsrzMKgeFMtF/mtWIy1cFhcvFsgR
kpZHiWMm29C2hO5W6PgpFYmZ6eAlAYM38ZwOHKG3ekTqzyISbTKrTjdR5GqxUwPx
nNdVhcN+g7A9KWfZIAqtiI2IIzhksaMoq49QngxHkF6XunE/RwjKzILtPDyvAuLW
dWB2EPblbvFaNhh5Cb6oShJc+AL1ej6ufb4QTZaG3CFqB2UTPyHppn8l0SEOaIGB
f1j0fo9R6GMNyvlWyLn0okT8U/Bi+23XQsLitX5yuoch9XCTJzD4jPqbTw6NLeQU
ul4fy8Z4xopKa2Tbk7bJXa8YVgZ3Tfaar3dITtnqeQb0wndw6L2kjycQJMTkucE6
SxCJYh3voIQLuya2D4d+TnBQ/dOwWs811sPjmqO6QQeYyVFpHax1vD3u894P1v1a
c5KbJgMgpYvWDsNLAcwYf1x86im0Ut9DtVLgA21+GWMF6SbWu4JrV8aB4ExZNqGF
BStxHN5edY0PhO8sLoxoO35bYZw8Xg91qiXH7NJq7tLdKAqCwbi7h+t0oIXinuVZ
Af/wqquLGfdH2A5WWfSiob61jHPzDiRO2X7gSOHzzwcYlRDtlnRQCpQfd0feWRBC
DjDVfLFbZnRWh8eRXwYI1LFmHKcz0/T1Ssy6hqCor8/mbk7d8l6wUP79bsFmhaOH
fX2WcaCzGOya7Tt7PXKMbWgi6SFb/kpNMmdOiYqm5pEy480yUx7w3JZUyonpUwZb
HSAoBWjJ7PZWmD2tSHvrbZ5JyNZ7EmQy4vHfyMmybjQf5wFQXaTcuLY4b/v8ThwQ
4Tb96MzqAohO6RH5/XOzLi2q7BCW8J0M+AiBD8PTyBRZZ7SHu0rPidQcskxJJO59
S5naYpgQGQ912ASO5jqFF/MbZjupUWdT9Hbec9tLlrGQ7E0bBWGn2HZ+xxNZeYa+
Hn6YP+Xyv7u3DS4O4vFFl09GSyF9jdyXEXcBNc5Re0sKRxWjHNpo4y+0RUswChHE
fcz66RJpY3W3sGx1FYqFU1n+gc0kRw9pSqBUQToufeJPHTnH8zHSEGmt8nFDJl8e
nrTIXNIkxNMszVaWl8oaGNEJgPuL7Hxs3SpN81oyJtNZ32EvEqkXLvYoCkeNAcva
E99nMMWLy88BPbCRfgfVqvYj6siLJPfHYlYytTUgQnUZebPrmUW70Jrr+8CMMPA1
72EnsfXsMV4SE/Da+Gw31MnL4pz0DlJuA993gzzFFVE4GdJna4TeORzh3hcYNNSx
wL2jl45h07JJIBDTG30WVKepdiQL8V6/nphvS9VPJM1hwelqm0nLCGO3pk76GaIY
gMH9IUmyVBOVQVYHC1yR8/LnX8shXfZS7qR5CUEBOLifeRb+mu+ODclGpEBHXFba
s8BLGWGxbGwnkXpHsJBZt2vnc3dxtp/erkMoz0sTdq07FHwGfizBOQuIS08chx1C
pZbpDpJrQNbAniKZ37fMXK1Swi68A02k4Q5lzgMiqybXKSwVhAK4Qhs0fXSbXZ+l
8Pcsu0NoAU3Ii4wg4QlGjGjTRiQgBgNNMc3B6BZ4jQe7OIZ7Ypaz+oualEXa9LLn
utOf+SAhhEuPofXVXiFa8BV8MQX5mBbOGu+jD8l3cwsZVFGvikeV7e8Cr7oCu4YT
RRP3k8YHiS6knSwwtsq5KWaT8G4Cm+WBe8AuDIla++j4fDQFOXdElAfBWUR0BdFM
4steEVWtIE+Kb6C15bRFgCxuL4vcOSg3EdXEv9nOlq9zaXIZu5ZWQmZZU1cRwig8
amhn/F+rQzdxdr7/PqTYpEfg8tFHUyd0kHA4OypE1zVuM5E876aZGFOp5pMyGoWy
09axocoRfyWx3HhHme5QyIT2B5RvMr7eSWWytSqyDcaGhmTA7q13X4jM5Hyw+/b9
0QvvF6b1g0Z8qr9jhpe+/UBedjMFqyC2wvfPD7wv55Iwni9I02xjSXQVf32c8hIU
5Dmz6MJtpAQsiPypUGdQk2i/7c+GoJdI+wQ9Zgd+G7yFUIU9YgNNjwS3z9jeo8gl
MO9a4hmRv9fSgJP3iyl8HswShDY3X/hU0M5URzeal8PTiRg/JnaTbAa6Jas3OIBJ
hd3J73MXr7O/ACRPySjRmyBcsycMEeCAfL76L66zUJP0AmwL6WRxsbRuJFVCNZrd
cVIfzptmBL+aOmw47o7Ndy/RjjTGBOyO9F89GJ9aiYtobIGoTa/6zj8lCQCEpumT
YVBhQb3SsgZjlJPlNPehczUFacJZVQhafgeFN76AjytryFksjvgWIqBk2g3xY4Bh
8miP26PXYvULpeqqEFYkigkMH7tigYL5PMgEk+vQ7Do37+MdnfTSy0gPsDPUWdEI
meCJ9r0F3HL7/KW6+I8HEowibb5hxDRV0b4JgWyFivl448P8nGM4UlP1aznofmdO
luZSUj5v6+pD8a5Sg260tEqtESffefTDqa7oUdeT3u5/LP8Zxx4hTCvtUnMFM8Nk
QtpBJv66+1hCxip3aRfPDcEpBcnPBUfuaEFxS2k7zNiOU6VCmYzfjAM4EhE9Fw6Z
KiMdE5Xx3Mwrqbg9PqccCkQgfkbgJHbt/qo0/NGO5/XOrc9WOLJzSXl+uWMWB0gy
7cyqiDA8VG4tLLDGHCEjnL7Tsmj0Xj0Lgf9ScPyXPYTlKfSQu5ASVG1OTcA8rKie
FdltpVFhsLIuf//jY4E7/3KEMUvaE/fZ/A6M55Y0XyGhQkru91Lu6H29R82mQF85
OzTsqvQpdHMLYV5p6w2suI0qUWZuLaHYwOhe1PHux/Y6OjmKT8LLnj7MWBDItm5C
J0pwhb8sAuvCLhDeeVpJgMsbBQAtawkXj6AF6Pz1adKxdVSv8eECAXgSGXC+uxXN
dKJgTBTZK5osz0uJG+DRo0AdedV/2hMgpK8Pd+a8rQCSr09DQ/ApXSqteLXby7qZ
hH+7ji0U11YmDZetNVmAbQ63uhJ42Duo3rLi6TDcY26oh9qUzXCz4c5wHaM9STZj
dNgWbPlkeFp7LGYE9tynv4+0QvBeK4JcBtRmSvhqZwzOxH4ivRDdcVmaJ1n60Ca5
+IM3RNEr+M8WxjIGDVgh8jZKeCJMvTAspFu5VGXOJA/mPjH0zmhuqGEIC6WBC01C
wipSNM1lJ50B1UJ2MXUpojJB1zFvkEYlNmwqTOG3W0oE0FpEnxFHpGhzgh4an+jD
jXYjJ4sJzstoM4i2yAdOK86zmgRfiEkJvkjecJDJfilF4+gsMFmBRPsTCJqg5DQL
mJvOSnKk207MA80fjLuJUE354iG3gbwb0ZRbenVXaVAJ6N/7L1Isds40EE6QILkQ
Aj3vY/Mo7AL8aAlzbOztTDW6tKArzTOvoaiUeHBUFc92JE5Qpaz3zghAgKsXPwwo
tKithYxHIOWpkrnZZmg+JzdGOTtov1LolSYdqGVf12oP2AolfywV0Zcpm8j1g2iY
+Jp8jUuBdjBbpZxLlL/ygySyZPx59IUhtwuYkVL8FEjzbqaYvNnxHo6cxJAL/r5t
O5ZUxlBhf2mQZKUaaDuEy3mPNEtQn5Lfv2J3s+a+t4ldYch0ffPzRbz/FwkyEK7C
Jif50CuulqLD8HWO0uDTKPaWsiPxb7bROR9bBYGRU+x6PowwI5zHtGJB+QZD4cl5
23Y6gfVLw9B6lY1jq2HV0ZlrL442/bm0RG6VSf1XlNci8mB1vlBv9zDhN+OQ5jvt
0zfcMk69Guzzn2BLSwNknz8TcWzPz6SXygFpoQr58TnxEstCUrZwU+mFPEZ4py/3
z7jORV1pZX8aeMH3ZFSI9wQgXf0fE87Iaf9I5rOBs7kEMjRKJUfwt4kXE/5j2b/L
AcLxUD5MN4ZcmCv74cfaS+Zs4+k9ii9cx7mLZ2gmkTZdcnSrDmtFb17NZ/l4ojCu
kQ06LbT6jX5t6qur2xEbSnzqQ+apiSNVNewwch1MNk/i6wsZ2PGiG6mmZ4CuIMuQ
meDdPA2q2uwTzXJOA6CoG0CtCReBqM1GKg7uppSXGXNHLSavG3ZxlpkSHEcfBVXL
WFfn+YURjV8/MW80BWt21ziNnOvGhjeRYqGkGdAG2G8KTLPKlfkHqwkUzwX3ZFPB
IaTw4YF1y+fogpyBOlrjGszqBxzbYGNvUSJbWBgA8LsxxStGje+AMGFhN1PVMuIm
8BbMpKkHb2vptg60y6OkcQfkeoCgXnr+pk3rnWm9qQ4e3fAQ3Ie2fHFr7QemH08n
`protect end_protected