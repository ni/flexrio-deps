`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1952 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
yuiAF2djpiMVQLjverTUdL2/04J95FrIXpCK0CkYwhFrFKQbFuht4zv4bPTWb7+I
2NYgbqNWES1mZuozrp0/1weIL3qQmL1ObjKseHgC7tk6Qy0yxiX8UMI9YIJ0cY5x
0TE8qRvWqyhQSUXO+6YcGoVDzY7NhN0SLyqk8Dp7nZJtKFs2BBKhDmUdidbmaL9L
eWhIRDuF1ltAU+lwZBduj1cx0X4ylvGY4Nos6L74yx5HjmVGAPdLNYZ7o4AIF93y
dg3fprgL+weCm1eZa6AHfts01htSzclKOn5s9BLv/GwfleIEHsFNphso6rvpcg9a
EB4TjEZFWi8aYfZ5B6HBjlPL3M5eiI5Xu91/YdBEabhMf3gAPqyWXNnq7+F1XWVk
zkZu9sQ4aV6b9g7eWx33hnEchpj7C1HU0coABcQlF9mkVQJ37x13t+a7AXlJaI+q
khCXhn/dhXzLf4sye3pPeVm4quFAVKoBUV9d/NHwufkSS++HYyxb7KW3u4epmVLp
8UtViWraEj9YdsSavCL1TRbq8CF99iUS405/G1VFBXZ2SMSCKfO+JywHsOYregMh
r7TbDT/erf3PPiqVLjRMGCOQNh75SAIO0vDWRNTJTdAPDsNNYjNtL7EaOGB/2ZDc
X+hOV6HoHuzUsbzWVHT+ucNYMg5VearsE4Dow4Ya6DF2ghuYqeDEblgYj0Yj/516
8o86ZxQw9+eltKBzpxXY71rBeWc51e+i8elcabs5wZsdlT0wrD1cRv0XYCkC8ZO7
A2iOCouUDB6RYfcC4M8ia5LX0UIOzeTacyYheQKMoMTFdXLIxl0I3P59PEdjcSbk
Pwtj05/q0KtUu3XgB+HPajhMhzNeN3o8IQD77+CVCL7YRJsLnppw3F61nmOj3hxu
7UqYtou9tAQzyGbHFxIePk/s1qewMnnASVyneFNUJC/wFvZ2yCwVzHWmmAsgaupq
Q6bt7R2nQ7TSIsL3ZsgjhlRL7qNoSd+1VfUx2f6A7JgWHb/6dB7KMU8tmEJI/PLw
t9NMuvP5PMssnE+C1AoLTvzkLIOrNH2wtDIhk9Dts96RxhSe71XzMLsdQct4d8sq
YUlFFPs/M8hhnRYzA13VUKKtYSKd9iajOirLQw/rPAs8NaThSbmbJ3eoR1+3eszm
fXlst9DCtVC4MtXOKggSMQvSmxp0u+liZVxIaDlh/c65vyfy2GHcrJxpc4pDaDfs
+LrE8dhJnwk0Cp6NQTwCvxpRxRDuYQ76Gl6azKcnnD/NtimmLGSI+7venIJ2JtYX
FdkxcXo83PdcJKq0oBXQ/pSOLNZIYgosiJc7laEqvT3yGMAQxSdzG04jxADPlDH8
fnVfBxk4tt9Lw//QxLL5EUgD/emqdaN3a7vkY3AzZGgYmKoIwz/Q6UG1fGzuqPTj
ksyjmJgnxKZMSvY6LwQ/NAOn+B+Y3nGtqCmVw8SeijrvwpD/T7uGNPg056ie44bx
C0IB8cADG6OqNhjyJ4SgyTMAeVjFYNoSuasgdpcydTgVZDMPvt2qjKNO0H2kSuad
gqqdToMmKrdww3PqFlrw48dBRa9V1JzWuQLn48nj6oXV2h2sQokgtu6fYp9KuxNY
I7265pTrLHqTVUGcgL8tyLPX6yh1udSc2AAJ2R/pWFIht285uvydF3a6aTj3pimQ
IsJtb1c2NM4catZEAIy7B1Z9b7LPXloXVUw4Ew+Kst+JXaJ5gvQUjB6CxG7fll1W
VWI7zaIS0ES9f5jQBexJ+g3xjrpQy97k3tUVSxvpIP4WOhpOE4Lt6eF0lM359Me1
Zt37psYjSKfc2/tf37f2TFuCotgTFIghdprkmDV6IDBc/VwoiimdkemKl46iNW+v
4DSdnbD2xZUviOrGjGYGT+z8nahLvYcOfelfzMgGqZ5zWkBYfhUzEBcSfAMiPuBZ
8tSNHfL2vr4qMFYxfHHlVXJIoPUj3ZHHY7AShCTyR9osF1sUoqDOPq1KQHJJq1WJ
yzf5ZPHzVWwzGLDCRKP8ecx4pe9pCEuEaI5KTblxma1I4t6IjHOPSg4yyP4XF3gv
Q3m+elLpG01+iK1s45h6dtyBc/Zxs2gTCul/hIgoEu4HeeynUC+eBAl61YWRkrXB
lKKfODztDGZX/hP/kXKF7zCfsxRIyT6d0BxLq38K3aAySVV2Egjnur/hWtJWwfJz
2Z3KzKuRYd8Omd8bfh+8FZ4UMbQvTbZXK2G/whMgMoBVXHbnSWoyTQzW1knN4JHI
oCxH7BK3AwaDSjX14k4c4khcCIDBa8PCT92hw2EM/tUG3vxdBEIL/1R6kM/c09A2
DmVEKRQ55uLiFxOBgRzSp7d4pS1BGGhbNopupdL/Ud5cqkAFBDZDm5n3AOLyV9Zy
r5hkJf6XxDHNZrygDBlolPeGC6xioHVveNGF+Nztyw+XrL3a4c9AxhOSIoHSZPwY
ZZMmR9RD7Oh44HpQ7mxp94RgvsfD/Ikka+F8evtdIro=
`protect end_protected