`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11232 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
1z1b9VGiiW9Gp7THxpOgEbxcckaEJrZm8yE0Y9Z3eUsOWW7oCujLlSwKgvwT9oE0
HsXnhzme6HFdX2/PKzJ/7mvATeaMp7/u4NF2GZEA9cIcGedC62IHchaD1FL1e3Nn
4PMGRxgXNkXnSgd9at+ihI65HuZ2JGV/DIKqGK2nM6pakOrX6QN2qr/PmskqFtvq
C2SwZVNT+5tzWPT/WMW3/rDTmz6hj/KvCASsSL/3+55e9vj9dfhTA4aHRasBKfYy
DG0NNvquvwbF1BgfU0Bhr7EQJFAWcJv+SI1ZvaF2EmTiBDMmZrrC3Dmpc6SKlklC
JleeVeyWz3uUUttVOygdK6Q431ZAnlr55d27iuHV8dvjH1ZLpDMFv4Y4hHUp50/a
hQUGKTY+XJjwiQ+5KwKiT1NIdxf26z2lZgxIfhHFbn77tYb90vd10DkS+9Ddvaww
nFxqfico5+zKXL/gdXCfud1GLxiL7OyCQt87TGst2bPMKXTvpZNL9q0Y2oSTZXni
NqFMJot4SG8WsxP+x0Pq1p0rqX0vQMlprINkGD1eiZpPS5EXl8p3bVPvP05VnxPG
AR/UN2kPJEQeW0nk2nXYrYRfuXVucrHqm2Cg54MGoIOat/LE/f1AQ7tsvxs7TVZJ
VW9wRNCZOwNMEePrSc8vHz76i/OXlAtnSlCTf9qyQjexxXxD1zHa71Mti6KX9mKu
7cbVhycI3GXcxOOnI9BU9khOUeHENVxP7w68hW0dPKL/AfV3eiUMv+I2tDUB0XZb
uNbqTNSf3OGtBQMUxaxg6DUIXUQ51dce+c7XNbwRqeaongzTX6gbPV35mUMtDiEB
1grcqv0xvcsDR73qtpdMWdAR9bS3CinElXqXQp8uRSNu3FkGM/iPRuSG+xNw8jM8
udcmH+IwzEf84geJ+Ow3x9klWvu3N7szV8Sg6glG2WKxiVoQtWkwOs0qWlwlIo4y
+wlGYeE+orSSaDCkRKVaynJEod9qVFTddvKOYHl2jCja004DEjdzsQ2GD0eyzHyQ
ZcrzDLZTVWHfZeznvEJIimlg0l7mo0/nuKAJQllB07qkT5NxK7VrVo3n8qDAkU+o
sHRQjMPmySYILpJ7O+ru8xbkIlJsVL96r+2AXe2l9/rTlVcmczyyKYNe2nlOpfw/
kFOG1ZoG3D14TC1IEkttPpX9TEsgtd5yyzBBMBaka9ARoBZTnHCONhtsdRkXeusk
JrJv+3ArdFQC11AXOfMUv7zopSdpj/vbw/uE3rQhaY+KPM5/HPJE/HV+M80DuEdw
7fsWZO5dK0UGJaVA9ohSmjYRrGR8Tz7N6OZUp12Xa4VHlXQaYYAJ7j4rIDjH7YSA
5eUCa3WtiIkz9XAC2tFnL4ZlWotwUYa+FUUFZtEjT874CRHOaeyycRKh9icY/pDL
aYS2blDdriCTNO9bpYV4cqRR9Lvwo2ES7uuPYKCSjELnnf3wIYznBzTzogWPwRat
Y38lHz5zwVkOI5MelMk2W03DJie3kn4MEnTTyzRuinAi3I6SW5GNuugvlwVAry2D
pu2alfWkqxp4wGlLr1xKCrUfHb97gYGiUKKcqKIlgP//o/KRwgJq1OSsGTxDuGGc
kPzTWGgLqzAOCAqNd6pvRGfmuRdJVA/w4bPmOFVXAY0Jjx4UwvN24GYkD+EtV6wd
bXt5mHwrBdqYLjer1q2foOq01D5SfYOb/1rjT0YaH/4Er5cd7huOoeMUa/aOdnxA
937cO/llEWV3WXeD3XqecvNnky9tJvjShaB2boOi47wcGyyUyQdq5Ct79D7noHio
R2BO0xiaTWW/y3yqxDPsXprhKfaYIWaQAPJ3IYmAimozJh7PAp96iRD6HZ29K8bs
gZMuxB/eSaKfzVe7iuB5KauUNsVpEd7KtQTR2eM1ypIGfHL9MB2pGrhbglC+xyq+
x37BsrlwPNfvi/MuyoQ/1QGRCyyZk8EFx47C1M4mXoVLpWaJ8qI89wunT1fcQa4O
CtJ6mjdmwX8xo1jL4nfMGtoMGUfc5BLY8D7o9kmslyONBm5V5vo9KuDHNql4BcY9
eIRf79CmO8SCdDC0DQYEHxRPz+Cpo5XeGR1KxRE++11SchiRfdW1Tp6a2+j/5do6
N6Ru/NRpL+n/EG7AMig1Cwg4X1mAAWrRcFDCFbX1Pz9+B85jI8Ega0ZC3ekCn8wO
7g7XiUrPXv4Bw3X1t1/6SHg7JH6W1li110RsnT2rd7fr3QAf+yI7QILV21Xv9P/p
dZas2DWcjiWGvi5iyoe1ejrN4hty8Rs/cSS8BuelPi4jbEw63S/CQSbDPQc5l9ol
wSGOSaJIZlQ4m/w2dJJererfQnPw964Da7pdavLR44o4oXAkv5pwKTNpVEUqfHjt
bMOfMbgeXzBzheZj24jUueYMWUus7TvdOWPVcKr/nso4It9Hvq3XF0n0WK/vnI2u
xWknH7RSk1PFRuzMYp4wRg4DdqAv3nxO1eqQqfp9Ga1mYXf8yE4Y/xGGmt/1G5h7
78smhQ85Gag3Xq/gZnfy2UWiKEORsp75WSk+fVwkO0ObSuBjIG0SxypdlM37w3Qv
UcFm+xQOKPWyFqr56b1HXHpetBR/wbH3arDEu2R0D7pLzpGXgWWoepwr4QXxBp8K
i6uRETqCYQpkavnhWNxqhscqNZPLMgluYURp61vJiFWadbJc/RbtGD+McICGj/tw
e9St0LkV85wN1QU+wTMUjh3nIOSEDPOu01w91p9UQwh673uT0rncSZPruvgWgrIl
DHoVVHLNoXQTdwX7D220vM1UngBOH8uibA1fN/5jd096+Ik1WyFGXyY540MyNWOV
4av+8/ZfxRMHtf+3eLGmrgZhTY1TvrLIH+k+yOe6L8ipnYnC4vaNNJrO+NdizM3w
K2B9Y6GXZCwLGJSZHq4E+rqypWrxwC4NCrqgO+E++NgbJBqg8R2hkVwgLQYvjdWF
jWY+mmuT/VF+ONtOJ7bTqf4L8r272Ev7IM2HsTBO37UoebCwKeszNDdZuSKVvZE5
f3l3uDf1h6Bv09Cv2l2Wfe9MGyov/niRzp7CFCm0Eo8RuEj3TujZKzW/faIb4/0S
jixFHGeb0mvEJ7ABg8ikQ8ZoZErr+iNourGa7jHL/YwTzekBqP5IMNlcYil/tadN
PMX2bhoAiLRJXksMJkQsMsA6b9tFGNJh4MmdzIEpjptJoviziFC2kL8Hkrs7dSHc
9GDY2Iu4P5qPjGMMZtEmgrECh1zTEqDBh3QQwdnqbhLqB87gh87Fn4LVPac+ZXxm
d7SCfRrPbQdAzOWYq3IPXOx9CayFq4cR2AbpcaS98Nghn/cyfYPFVOTayzqv32i3
utY9HXaowb2rf7cz3ZKcIS9gO93kBlnaV9QLkc3rl6rmd4wl3sVcSIL4/FWAgWSv
wmJyAuMXWYFf1KJuGD8Odk0YxhyjXGD4gT2JZyn8oHTHJ3AVLV/Ie7I3jeQ6pYa5
dngbKzO/5zwLwYg8MHhKLoBsnICV36kVhJbUSW5L/BpzR4YB5XVq5JtltBBBBD0R
BcHYhy9aMxFzWgr52xvsi7jdk6yzIwHKPYXEjDy0ag3tOS8sh8OYYSsykUGi2Bbo
uTJhKrQaomrUsmqiDLZ7IntruMsMXZAdOYXuRdeQfxg2KYlgHRtYBIjjYx9v6jpK
F9r4lF+Ylk+6BHDmjETMjSxAElNBKVBkbp1vfj06TUw0mX2hnfoOR+1t6uvrPuh7
mPpkG/ewddrZr8dFMETLIKQH9QKmNY8QXrJRz6SpnTA7cNWxDAlaLlWCOqD7uum0
NhpyGF/DdSrWi6yozZRlYrXcdT6I4WjkMyS5ADz7AnJGLERu0U5Kth7Vkn2nX0Kw
V5SA2aI9W8wEz8cbqS5GjYcItHif2+gsmSiymO+gAb8FXaO+LzUj9o3OSzYi1UP8
vNolmhdyeGGGdzY5WhUSYjFwpaVO3UbfeQi0o7t01P/8b0aQBnzUEP5Zh+xHHxuE
EVwBMaBmDksFaYszy1vfHhT1NoRkpbnXNku3IA7P1nGHoDCCKWRBjqwzlcuVLoYR
Se6Uyp7rqbrK/R/7aLby3zl7MDCFw8j8aTqQHmPBQJ6jdfsAgU1G555NwbVxi6xL
svgQ/3OYxQFmiEAJbv6S6w4NrFW8Bz6VXuKIFijLKTRKnHs7gMsxLPcuqlzzXi17
EDr3CjChwueFW5GAjnBuWd5Wawn7RLnSE0mdC35OzfcpRbs58GasAaIxhFh2MreH
kfKtMPRuY6vcbC3GbJk/XNvp7osExPMc64gnMAIkAY89j2eR9tC4hOBIm3dSd+dO
S08/QEjqNjNh8KbQZ5TrSCdK5I8YglMYhoH8GKUhICoWGwP1/wO1xzJ/LVz9d4pi
8/WDblipFTLcG4a8VnsXxTBH+pLceoQWTRDrbHfIOd+ixCXr89FZc6zy0d9yT3mj
FJk73twHa1RK7noljJiup+2YGyBkRVqND7fSbgdT+EizHGvZjlYuCArPKljMuu65
pHNNE875ADecnSDwt4LWmdJmDJXUd3RmIrloap7Ix9DX0wm5vJkN3xdawueWAtMh
JGlwYqFnhWANSXMKlbTrzeQB0pVRFIt3GcyNc7IDJc9e2ZEJf70SiJCfz4X7BLO3
QkBD9uXf4nHO/AZqIzHrMhVrQn2LVBrvCVr9EMF5j4qVw9SlH8MMIGUmqzOxymeM
g8IAddDsRUGyfPNU66t2i4N2vtK5LcyOFAAtqJ8sKbdh/xVMIPHTiE7Uaw+XhV8K
B2W251jN8noRp2KbMhQurEL+hpPPG40KIpcRIiBcio81/koHxsVFuOyklGTTcGpA
M4a1g0otrWmK0Nj3mgIFPmUE1eVaQc6xNz7LwN7wgzD5W2BSq3DHHb+CLx3rOY42
ltXY2qUVzuLV68X1Bb9Y6bJNABzod+suUnazuyDmtdmRoQvKC0B5oHHIdW3dmpdC
XQ8bmhIw/wzyTR6t/wAHQMS3NokesHJN5M0Ozrvt4KPoXtJugGcqj4JJxapoSpy7
kbF1FwtDoexQ/aqdLxucThwooVmN+QtqEhR+NFHu0WCOs9ZfJMh9Sc3t3TNDpS65
1D13e067GJYKifTdrh+5IedOBaJjeF6VCd5OU70dyyHraWLb4RDEaXzHB51zW0K2
flSzgzSFGnZ3Exo11d2wFXO/Ko6FgJIxlzppK6h3ce6A6d5frPwt9Fm2TCzlf9YM
O444jjy1qXNIlduwIOLwMRn8c7LpezfgY1ezuHzjmXK9ilEwR2Bnks6DG0JUZgFm
LAs9wUHHgka8I9QVShS0K4nl2OstZL+/4gGKEIvqWRNmOUSUQFoA+mK8dOwHoNAX
Gbh18alrv58St6WX8mxWNU8xJV4SWITgWLy4vVTalIxLdnLiMkpd6HszNOoWQB5t
PMVlkCx45ZwyXQXzl9EWkd82SjUbZZQZe4shXkfB/qH3KzKzCDnr8uwdVmdcLUYz
pGoNZZrtdgcm0EBeN6RMdgR8DzWlRi2J20wcDhZTa//ZiZhucllhQ/R0IqmP4cf1
npVShcITOsuy0FMD+HpUyaIPi1gz96yNzWHWWxa7mEGT6RaBh0qlli22brz1+OlB
yasxKOXU1D/pLiGpc4orufSab1uiFZSER8dZf4JAhkAPnfoROd/834DMkZdt9jdv
0VjY1oLrG4OEFVJsfssdJGxsTSr5v2cq2zIZgbFEAy2roqka+PbM8tfPUJWSTt2S
mvsIZQoiW/io3s0xZmqDpTC2pvJczQf6PbElvtSv4XdFUQhazUZUjihW5/4uKT43
OG7yBv/5K1YSr+gNUmvAq91WHLPSQAGMe8mCYzZ6YdVvZsHp44tVsMDsXImvjvhO
KGcvbefCZCIFC3Gk2BRYXEFT+b9PDa4T6z906LBuZjX0QOQKrPIMfScTht+q8Hb9
HyCY/axlQrlQhisFi02R17BX73/yCYDWVySV6W0OErgXbzXLXYibMaTyWYsEbX3W
Dt4iwG//ayaTn/2PNyIHL2PG5zb+M93RRQ1e9h8oHfmhIjmHx53IScKfYtUqd5wa
GUUmRQVOuuieVP3P6gHeLKC95USM/8OamIF0z5JZOBBHUt6QzFnpq4hIIO9nd1Na
iskdh8gYmvqiFaBcv4D0GMKgfxr6FcTWMwAC1EeiVljwAc7ESeLGdnJ6Fj9z/UgX
GzJjFUYbzPuhLGF7JdnkSmuQIlf8BHvH8Of+h0gzUR3WiFSp8cYylAA0WI6ZLLI4
84srCSJ+FZ66pyyeYJpiEMhy0wkzj5Q2YBWE9YHeWZOgx/G/EfnDHAMLPCZClDNQ
jxOPTM7yAWIr2eiBbFxVKgjanU6YS4MnPhNHoKmIwrcMCe3S4sZm7Kq41pKLwKXb
BJDpcvHsrK2KM8QuRQ7ZZuCsuhGZ2f0FSldctsuNmqYiJByOdWBjl48V77z9iEcu
YgZpGnBvJ5s5y0ySmAFgULU3IX2ew5NPVbmtJHKT6taMmgP8IkH0RpgEe6wlEOZc
fpxX9SjFAgZngzuovf/eknqZcbl6VqsXxrd7X6nM89d7mYibAJRF/V55NeGqZ/Gc
B8LoIG/F3/IagGXjyJI8YGdv+ezpupKAk8l9MEiV3tWH0A5TsfJkDpaTs4kL8DuO
DIuyCX0kMKL2qZA1ppQOttbyVabHKFHBW3lfZBOTsarvuVSUFTyUs8LZyZxmTGAW
d+V3csIqRD96/2BrPLAbpdN6pgkib+wt5u5I3U1M39OXrR3mDd/KrDfvvu8D1j4U
f7/qa/TTmKDVFeJDzOmMKO/0aGYHEkwEUtFPdBSUvLeLUCbE6qQh46eYc+1jxIrw
Ru3/I0/MHnJzfsNyFnynIdPph6hZnk8BUKEsG076uBWxJPjP8nDeIMw40TIEkCbb
jUBX1VmUBcd9AyySY3ugMbErjidu46S2lv9bnS552iUaRj95x37W9XgCqYKpcurE
AKk7HWN0Nj4L4myakS6sjepIctpWfO3imYmfxQYwhnxm/GMqcS+ahUroPovZqzq0
G+HvrqSgienzk7cGvon/Bm2w+RNxuQZo6uuagpXyz9u8u+u1hBVJOoHqM8LxIQuh
NmscEQfBrpSVu2QPtVi0pYMb1+KZf0CsaFZl37i5BObfJ2G39z2NdQqIdqxmFoax
cpNEsjmLGOOI6cMVWPcGlpnWjzHweWp0mP6PSuVhjYaIHS8GBoBmoe79MAqHVsab
+kqQkGr5JIaxJ88w8QbC7gKCkIu8AwzjCrhp8uzAg90JcwoCYAegEEZpBXFaGrWN
YxjwdY9dWsfdkS6xBsy94k9aN1rDlcrA1a0h0GW1DNx1XV/86ATainbN3ARkK8HC
rg8uXKdTD1R9fsVv/zPujw8LJV3CKdMQ+B23dxYWeqn78v/utIU0BzgGNkZRFhGq
lvjoe5qL5EG+TGoCcDUbhs3mqCKgvshdU99Qc3yxzp4vX89iDk+4hNwZxyeK+wnH
DUPNW5lWevL61fBum5XayBFVKNf0CUjCqS6gJtebRmGA3pVgh9R4UXVhce8Gt2A6
obIgenJb0mV+7KvdeVImuKUPPYD9X474rjB9mAuuRhe4BXDv4Qz0A95MqgD5TW8l
g53w7RYCI0T5V8NUgzyAGi7we9ZXEPEPYINGkHgodrfoGmveQJ1lhexsFpTgRGPR
UqV7HNqKXIhBYsDkbJw56YeCDQXdiqKudYKcVPI6NHXr6pLEojHHgisXhzT1jzR8
6WFZQmtPceoIPwRrQJx6p9rm+BzypIxEHEUhR1BCDiFefuu5Jt4VNb52lt9Kb+VK
o+AqPRRA2Q5Ao3vbp8KIqUPzhEmkpu2En09/A7gvdzePfVD38E1cOeW0vOqjtbGh
Hy8hHHEz+1nKQwTPut0P4O+FKK/r9jPcM7dNf4uDhOqLTI3IboDWz4a0U1CT1sNr
bH6dmGVmnHt94zaqoha1G3wmqZs+pWpuW7knJw39S4DjoccV2bAP6ETFpftqyd7q
nT9ZtNOIYniAt13zsMrc8tOdBFGPoQFHykbX1lATzWUsLHP3Y8UE4arfFAiKcKwW
kkidws87NoTMYCUMnb1A++8/WFK43LzLuiW1bdpO5LKf0YqpAM54nPEaeW/UPeQC
ugZOfdQpF4Tia6TFAENa5hVAaYEbwhhr6+AJN9GKeFnhFdqiD7ZmoIFYtRB5UaHD
SLXbkFxU5g8o8TMGRiYluNVh7TZx1eoghLsJPt3vIja4RYmkK0l+oKkY9ZPYsOF3
QH9kTfrDfhqrshGpCGOZYgzQljLMBdpwwpgA3LeAKiV+w/y5l1Ho3A4EK/vnh7sD
1mRSE1GcooJ3VFAs5+8mvOdUUPN16d+M/UplIcoX0lSn66c6vhs3dGRgq69TC4MY
ZkmIZYGEL6qe4vmV4a2phR1mbht/p1fPTWQkh/4msxL8QogJdWKQNDl34Iy7UCyY
e/yHcQLmBb3P3j+8js3Dax5F9VjbzmeIxpZzRNNypPI5Jfvjzihc9UeDiiBNnxQp
e0RqxvcHPDvN6IpyF20tx3yYTO7cQ4OvYYP3mOXbVQDHqMa1SzyvTkew+Yh9i4PX
jWxFV1zW6MuWfKQl7pbvXFsznRlrxyrHIJO6ia3Td1v1s77gBjAK70qU8umG/owZ
7dVAAqYxGbNzAyjymmjaf1uok8vp1MYcCqv95tBBnAwwizRnecjp51DzUYW1/vLF
I3veuN73vDhJyr2nr+Texq/+TbWqzRj3HDWebrGcTCpB+/PV+VLdjOU0Ft5wY81n
qxHA/q/4cbnUn/EGaTey21+JGaDlgrgD03hREN7N4JOB3xbCmspuA2kHB77TGexz
KpQGsRxCNjXAtHQ5FQaYkqT0dn8LaW/c6jtPghQLOuiBL78feionRXz0hirF6JRl
ju6bj1h5JMdHm6pspFyQb1ORdLIzA0yfNkU0wTEG0LVLajLi+Gkms9Vbw43z+6yu
4ULFCLExKY4AGl0IYdiWGtdS929fUHzo0u7+MobSiHkIKfsLr5y+4g0SLka2Ikcf
3jMRM3luASSLtzS36W9PNZT9pw89+2wb88TQm5H+BZga5YSWX4PK8uzRMrcn8pb2
+jWnQraWKQq2vKQMOc2e14JWIp+TJrs5Q9Ha7bG0VCa6/H4GTX0rxGb2Gy4px0di
bM/pXn75KRVYDKxCJ5DlVzPhTD89mL+aM3rurjV4u+xeAo5lMc1fmoORN+aQSSiM
GbktalJ87xwm575Etzh4hRU1G/vb1M34aOKNPAEwsPeUudt09SpOAHqZaSs136Nt
FvIL1T4Ub/J7vHUrf19zi4qCZrlvxz3U7OeTK/klG4OSFdRcisM3dBxpfDOyVkOx
2SQC6l3+4/0ZfjlpFj8e+Kfa0NLQ7d6xG6A41JZ7jN6T4KAEdq2zlfnqr0GG2sgK
JT8ersCUOyULmCav8gF6oBnQ84rxTGx2SP6sspHQGLmG/i50NX+OEuDOZmHtotGO
DYghqAfmkwezLNWrpsKTYEMYVMYXPP264TnLW6PXIJ/OSBkraWKQl61ulHQWs0Ox
ju25MrXFlxmXDG4k7CdWfiQEyKB4V5axwaVF8Ru0nSm0vYBx1Askxhx1yEjXsUKs
7776AKZE5QB+LyTApirwg/c5d8ULMT9l6zX3iUOhD2oSHzIzLpVUAL21rQYAAnjJ
Tr3hIL5F6DNGAcstvHbJUSgLDVeKNLqVcn2a6C5raSZ6NXjQ/rul0qWKBi5eK+6m
x6BjntRBP9jzY7N9jcraFEgbdgaTevmakq7EN/KGw7bpt/iX6iaBu4/bGmd5OY7r
X9/3oZVGJdv98qbxIxh8SR7kZrzA4+yppai3fjR1n78LVTIykXX5C+exrJiiJ3KR
sXzPtVbkAKagxS5scXgt0VEnb3NshLZNje4v/AVJ/45PWy1nDGQALTbYVNZfN/9B
vAd8d9V6kplJ8fRuRqLk3vVTGhWuA2cfikZtzb5Yl4FHLiTNMvjVItZ6zgSEcI2p
CGJeMywZLlYC3I1rKzxxX1OGJYcoVWNhTNTmghlwb2e8SJwQ9fIomgK+piYkPzV4
bPCTKzTY0ip+9z3tPIfqQzb+26WaLaesecsmMD1Q6oPWzfLuECmfjZo4VNxbuczb
MjBjs/5w0KOqsSH20/u5BhjEjxyhJn5fQcLTwVf43QaEPq4mRNWHKWCXWVHGw0RA
dCzO9qoUlIcHmXwUUCsbpE2RJRce28+VgZ6NWvvsJT1wlPxJXDMxcKcgK5vISy84
HsbWWLPkOuJRbS6ARLpozzR0nc8NbAiArwwC3Prfa1fYWLenqUX6VQOaCtRFwdYr
/IwmPhCDpKCB5RRG9xNJdoTrE/KENeaRb69JskPOR1/X4I3pXy3l6eRB7C3kPhoi
tg27F12/K6uVmbVbRt0KucTWZUJb3M0kZQQhDn1zsDWRkurY7HDM1X9VL+wYZWUX
nLSChPwSaOPbVKt5MEbKrnWL4cF5Vj9HXBghS+y9lhRktc6deN2Kp26lmAD0NM1q
fBixQANwBAzDyroBZ4EY0owYbzz0bEs4WO5jSlkm3FjMGjQt7RzdXASU7I2ba/7t
22F3KgBQRoy/1B731KPb2YNQDGRt0/zyENTuuYtFzBNw/lZbBesumjLOn529lhp2
BQDwwSIt91F6DdhWmyJAZfg3Cpqls0Ad74om6epYxtZyn3WDkax9PsArLERONjRX
32pdlviTC3Kw30Unjp5R7MQrSBC7mX6pJJDOaRS+oIF918QjNLFjhM1s1aUQARAN
BksxJAasPYalYVgM8fN4M03J8PSqh3c0vPtFjoGQnQvWXk3HDjrmxBfCrOCZ9ov1
8x8Umsa5d59xBwdikee/G1puDXqgkEvH5YJOEi2jwg6PnRvQgTrivtpcyFWGOU94
PN7GVeoDDtjkyoPM88hK50oLyDxFcSaL4LIe5t7IcRT4CMC8rBZhyQ/HMMvNJSfW
eNEo7ABTKR7JRpNZbQnKD5OLI33lcmvS19PGVZZghPKMKmoEB7wlZckI2CQDn1wn
dcouVbmshCbMGrzpRWX5WVFNe3+3U91IdFoJdj2LOgbE6E0N13UVmRgZRbAMHoBC
HFpqrrcJrPsLceZ+6XA1pkFv8lIR3yO8PFefAEeQX4B70rqkEfaJXexsuZ01tsWn
wh+SpMvL4hJ3zUdi5OZDSIP2oPNDMNRf0ndW9tWoYBnJoJ3w/4lTo/urfndEOQI8
G6Za8VZ4kCTME+pRLjVCNCRM1z1FLlLM7IKdn1yUugvdmusjnjIDPhEUR/dRiKjr
A0vtTclP9vvRfvUmjgmY1/ZhpIeziJmts1niAcg+150n0b+K4T+sN7m5y4H5C/YV
5YJD7i8+Al3xRIHa8QQiGrgMbsAzIc+ZQUMg6gMGF2hFbv3pjkfg4n9ST/oDqrBD
qQvx4BMCN9q3PYBBjvknSpDf7/o2/WLvMva61Do/13d1tGWnTa9TMqEQUzPwRECw
TGMDFAaf/HtX5OGkgM+Ya2rWB2sZs1JgfFsT9LWSuCBF0Z1fFQ4iw6S1t8+rYDLM
qVDDOWUpDxZq461/pji+5bi65ysGAP8HYufJWvLw1ZYUW6Dnmdcx1rqG/USmKmd9
c0D1LZHmOaWcQZantlu19tCgZNaxeQ9iOnPkXk8G2Jk/duNfJ/g/Tl+dDr/EN+36
JrcDfGlWVBWCLEq5ajiYAlJVqK+Ducho1DFil2B1JOe0cb+br+cwWgIoANIXlsBI
SoP3K2GB88ZQd+tJ59KleaDK3CJC5jWGm0fdL3GFlhfauVP1n9G8D9EkJtPsnDAM
sROsGorMw++sMWx4V39sJCbX4PMtyA7JIiTRhIJJzbxcQwN2zBPc5wWCqjn0mLnM
eEkCEgb6mg8UFZ9OVKP2ecpsd3mDMIxuccpwdTrHQWa1D6WkZMPrLV2eObBtq9sz
q1w4RD0z1bYXbdPzArwa+om5BXjBg6p4CMKG8bhEduODVaSCuFIfRKnJ8/nTviI4
SjH3EfIFOITheNHVsgDLVpgT895e82GDRHWy/xNodPEdW+/fEeRQ6i1Fpv5yBVfp
Gzt+Q8wgT0R9RMtUHpJYUcJZuZIT4RyzNkXMS6NyHU15U5r0ekrGO48qkHRJ4tc1
Np7oI562nxIJRS4LENDiXJ6GuDtIs1geXB849rDYg+Nl44c4v193mkHHvRWxSj6g
AakyI0xISVYANoAh89hw8OG8a8dLKUt/3gBQRNu1TxCR+eNOtor3EfJuZzLJaX5y
UG2bd+3pKu+xU9kAlhNB4gUQVpSwmsi2PVLUyvvVxGjfi3TYxphNEC74efxThFuv
wQDY6ciZLcP/ie6K311K2F2pCM9kqDLGgSaCIIubztJ1ecVWr8NVrDKgQFMEO9nI
AB+ZiJZ7VuwAqEpeVJ76JrKpIZbESiZzH+IIUKuh+Vfd3ZA/Y5VnfXsnlTFLhdHR
Pr6KgXRAkSWuFLqwmj12qL+WBt+bJwj7zLCcTVv5RV1PdEyW0WJnCIw64fpL5VrZ
tXoCDhVwbF50eSKe2DOp6s61G7GMOtMziCT+bjtMC+rpL6QsKSIUg24qWNKfNJDt
d/POZXXYLRj0FVcnZ8i0mHUwxOHGMKotiXQKzQljFS6l3K1UewrRMM4RRXvAkK2V
5vKdSKJxgqzOs+JNjFTYtrVtb19cwYbozKlAkuvtvYcRnG6o01xqeLArNSl5OaBW
LPSASdZemFpgL/7k7MhtEaKagb3IJXzSqG8bdmpA/nAYaDzQNAmG4HImlsgsNOoA
2WJ4tQa8Ss1eUxwMa7vEgrO3MVx7nhwKY8qT9hwoqQh70mSyw8ATR18qm7ZRplJa
xgtKvQvzhxdJFN37HVYG2st5WufxuN60z6UihJrrgpLNxoiuetWrhz2aSiZAwO0a
0OAyUht2q14SVX2O9/1hMuLWi6Dmlt92tCn4Tj+DPKJBYQX0TR0nGcnfTS7QBWHA
sJX8ztgjZNg4eS2QVmRQORy+Oq03HonWOJUPR5cUiLcM1Rxo+nPC6NKh7vq+OxLZ
0sU9/B8aRRSROtcUP7ogu9855O+amX2dOaAJepgsiKTiqjtzITKZogBgtS6zFwMM
qIaF+c6t9x7csBRKrmWgyPvQhHaZosgsKL51a7hnuqgShemWmkSQFnvSHCB3uDJv
pSTapjmWpnnyVfIEyFk8lbhB0NVlgUspevnuOqVKA4L2uw6C8FS7utkwSM/UowIu
NG0bEAt9Qjf0Tnk3dW7EDtfUMRYPGrBEU0Boc4i5SuMhtOoERciQxIb9UzzP+hRT
nSZmd7ug9II0wMogyiCY4LcyerC0vG5emi+j/uq77KYRNUS1LiT4l09NrMqDdBoI
K6YaMeaM53sUJdqDJjdvr9/L0y7kxV8MX6KrWXUMdK4bX21qI4ue+dki7Lhcbyoy
3VSSlQp0KWk/NqNaBtOuSybKzHGXEovL+2FIRe7xEcqUNn0MApHBIH+uEkAqDm0b
PE7RONc0ymmEC7Blk48DlV9ge7RapjAscvGQ6DdCrI6hFNG3EwkjykFTJQtNX3PE
qaJ4rGRmkFuioKo6hou+BNz+P0pWN908mpsrJ8DILckpVw3janddwdBSsauTAbnv
DyHsqMCUAjuM1F2/4fq7vDbr3jZ2C+pE2yQLlO5WbDtY0FzXRFF48aSb+GlcDxRt
A68A9EYl4kDWu417+t/5HMihPt3J5j3Y4G6xklxyswkc6x4WNFLRVLjX1jnaBbxG
+hBx0okZy0BIH0SwyChcIjBnP62Oc6yld+bBpbJ+C/kXAHeYClakwUkhafy2ap8G
/5mou+X3eb3ajtkQxwOQv41KmnmPM+XRi8eaWXeI8K4JdavnQnriRz2LrvUlzv1j
FnchtRM/mfQUFUTwkfov0sDGfz0wDEY1isZN3s9nNUicTDI1lwSlMURpC3YJIf3Q
TXgeOjJQM5xcbDzHK7NPwd9bssF3nrP9H/9tsl6seftdQ8pGe+9YIsTWN7ZpD4LQ
fIE/4hYJU0j47qDPP8EtpfHIsHBU+3XhQOJ8n6ljofGqj1qx39KBMDISaJGLExx5
s7pF8N7NmrAZrC4vXe635uAf2cdGVlq9wqeus3qcDprXJePHMytNodZtzmPBtYWR
gCpdr4m39sJVPhf+uvXE9k8RyzZVL9c9FJxlPEaNFd3Y8pJ28FBgM/22yB9snja8
7Xqwu1ZnBrbShDpcIjhx7AY0j3z1QaUVxs421NuvK58LCfl+DsZRNbt4rQ5JLgRX
PK1iwAwY3iBwbzz44gLyelEQNj8n+6q1ciw2sEdio5l6vqg74tymxvzBO3iK3d5G
M0EAc5CYEvbDxI1w29ukeg7/S6nS97WcbuSNQ8M/oItKT+NgGphWhoX6SmRqA+cF
rJk9Oi/F+l0d0KI0jDUyIxLMXZEqRqnl7mpknqWRYqvilRx/EHUJ/bQwtLy1eGNz
EMFwZ+c0q3/M+nQztcTu11/2Ly9wqGA/Ey41FcpAiHMWpnJOl3Jagv7MIjgbzcjT
SbZxzx2FhrtLz5tMUlsaeF0PS/RU/0h/CHGcMLXnBryyrVIuoG44a1s3J4dXA1VC
oXYnxgCXMQ6C9+MYdAX6EqVNkTAGpWBY5g/muYu4tKECdsmmsyBOv1FlNq7fkdcA
0EDkIMNH+1PFieokzIIWx7iLG7gROq+LkbgoA/SYjhizMmRufKHiTTjWNWrU2hLh
RgjQQVwDb/kkzdJbqvDTiUBw3GHU4Nvqa9i80V4SAUZSJiAq1/tf3wQ1/Zav8f/1
5sb3q0iE85nYoA7pL5nRcCbB09pao2SgX5PdIhEXaUTErDuUczRGAHEADFVg2kcl
D6Uq2ArI5F5XIe/uJWF3h9Cd4ZBlLxfPk8mbrdT57ZgEmyAFbygKluRgBD3m6WyT
DN43vT7s7CJpHFFgcB0WBmwj07Tazb5iNQKkCpLHFtM5tZ9vbQTzPzhhTb900izj
`protect end_protected