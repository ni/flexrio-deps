`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6272 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1wB2ShNYedzmkmBWjqK4Mg3
8iDfXbv5M0vDNkp8sRs0MIdGNHczGwwUkQJSZju64c83JtNlj8lbVu/mwVHcKXTP
+03nFcvGYD+Wpd1O27PkKGMBLXkn33Ag7OwOdVPjWP4y2hWeff7REzp2BXwC4eKq
PHcDjyTP3K4z6sJdYlOwzamNL30nDS3GxWAsyh8ktrfWf8wKmkgDW8ZSBt9q8Tcb
PIghUTSeKIbxGpgp1H8glBItiGxtwBUZOjcsXV+ieWftsgxPWdSe7n8jnV0k/bZz
ElBm1rIEAu7m3LZsrzoLFVPWfv+Q9PpPCW3gSnbGqyWvrPLeT4BeifEjnq5sY7rY
JfQyQANS//7efN480LWQmyjoHIkhSN3hr+OdRU74niE10t2o13jJj6E5QEdLxQi7
UhdAmaSmF+u9gEL0qkWvLBU68e28dPxy4aIa6XR1MbgDyQoWD39vhsAXiOGKOlJA
Bwf0EdMUicAWgVCxDoQED/5rWKozY11577FDCnYkxjqCr7Q2PVEHWtR+Epsfh1K2
dZ3dTpX45Vi/oa/hgUHfY2hxKBiVrU70nvwjcYU3prf3jEYiGzCNXgwoGyFbJQY7
IMBAdtYtHfa/Q5ByHh6aMTijarC97Bnap3EbIOwXcAp9KeHe2PfRca0GDp3tV5xv
Qzr8vdaq7ypJvsJ0r3+9w7WKVdA79/RNUJSUSt8Zzk47yI+bdqU260zy30aJsWEh
wCD3Dn9mo9f9n5RGg24OEUvWYqWQ6TxRioxXzlIum5OIyFzmxOS40IhbtloymufJ
dd49i4tRMcDTmbYKVt+zaaX6huNlzGvOn4SgtSeY6N1ro+z1FSyW8phlCjCga/1O
TUvBFdHKkqZQbWxUClQq7H21fX81bYZkFozZf9VTigcgpWtE55zNZ0GY9Y9CqHyj
txOd3Ko0oBdT6j1gE6/sh0NDWRXMU6OZ0wUt/rQp1Z5VFQ4FWbGVUT+C+DChZa1N
B6xP9cvYTC2IGfWtSPkJ9LRZLMGBCb0adX7Qj5ewmSPpqMNhU4sLCPUCyNTVH9sY
S/kxD85O91zU3HoJbTHt0Uee0+pRyjgg9m7uGNCRgTcb27jc/4boy8uZQ33NtbNL
TDGIf9FRRBUfUMktB29/yJDp0UUxyApXT0Fp0oM2rUz/hatQXdgE0OiVTvCRp52Y
4PaTEgz6gfzcdT88++ECUkzlWVUauW8/e6hxe/9kLAIwm6yMujDL5QS/Jx5cgGeZ
R2RrNWy5ZI6l56GMjrrbWcxrGUQrVejTlSaWrOgkYz6M6bT1NnezEDkPGPTfbU56
G8ezadZvu1S2JQ1pOe9a1CePSjeqHKRQr5Av1sdVggjb0G7swtI2Ofom1bWT8xzX
7NQ268p061DtbtnDhlzh8hR96IuI81xpN2QK7s2yQrmt+ucuVeTxAmWarU4jOKLY
wE/0MzSMZ0gG5BeoT4SiRY8g4F30jgrhYzz7gBdysz2hKc826BX7hb79iB+N+R+5
3Q9ktrFY9rYH755+7PwYeNq/zIWEc8xvZkf7Y9JMF8UvQ6sS3TuLdbg+j1Jik70/
PX42m7iSoLi58IMbVlm3iP5DDQhfbzlQ2I5QIjJTa9MArMt3PXl++aSkuN2qBJ3x
+8TpgNDvEeFRjSo4YsSEMC7bfbD+7n9dSNXgk0HQouuaCh74jWP9teFUKEVjfyIs
WS2sI73ykuhA/sDE/Yyda1rMiZ3m1FsD56tSSWeSm03K2uh7v4kz4JoYT1ij23Y1
lcbCsUC9qqVXn/9SivgZ0REyrbHmj3o+I5KZhlZlqT6ymbNedAtFQwheZcTIxeJL
abDwCgkDeiZSgtXnqsBCuH6weiHUisPNL/krJv3OG3t8mOqXjUSsp+2OIovHUfza
L94Z8E3ExfxjI4sKif5qsgES2EjN7nXcKhAtou4Vj9OSFLWu70jJOe+NTbCEJXKI
ECFOyPefBFoTtuemDigfpAfYTTf8V5ZOtgZVzttc665R0pNz315wmv5JboW89i6w
eZzw3Tpg4kiizprRghbYad8s7qX6jfJHA5n8wv1qBjqmjuye0XcGgNpz8e/ePsBN
Nw1G44CgnX4FWQAHoNyecUqEhVQtQuugcK8Nu0sDP5zwRYKgpXHUbKtuE6y8CCDb
WL8aYGmqTdx0ssuz9AVOdMEBTg0WcrzD7FH9MrwkAaRCxv2LP6LlAx8Ts0zstkLd
YZ4Y5mLIl7ewT+gxMXQINry51QYntOEztinbSSLo9MOoi4men/lNGbiOOclGSUGF
9JGRIKLT9JgA1XIGLWRufYLnqB6ZWbcnOgS+lz6twusZEfpn8xmG6XfgIL1qfbnv
hGWiLNKZWv4DDetEkI9vM3+XTJS8r+J9Ij0vtrfu373dXoU/z3RHcPNqyLMMuaUA
iVJ6i93BV2oLGVRZkBuwlkPl4W6J6eifOvaRCcE6YbBF9hPHZWW7hXmmyqAcM77Q
XoUg4Z2QSGfsIYSugBIS96fctPeSjdKxJJ7VtIkwE9CUUkzFAWMal+uuXlDN55O3
L/PBlk+XoQQ1qh4lCAaPo02BSe/nh6E6NstQjZ/kOuoTtZOTvGVSZcm4E8Wdk0fq
jeU0gxGkiryzjnTi25DXNvs3R5X8gsMGrjP95+GbwSdrfD/CQUjukpOnCe07Uxho
t/BkcxlBtsbnCuI/yHEEfguG+dTRaAB/zWwK54oAj5yJK7pwernJBPiPJH1repH3
22KK6xynVRDmviiwUrQDf/213fC2D8NaaLWqhGrPjJY+97Yw7nMd7qXmRDIEiafQ
36QbimlXji3h6Kgv93brATflzWzwr+P/9k2hXu3WfjNZb+s7wKJ+bK03CpjY//P8
BoRSCrTww9MBFdMFhNh4iHqb9GIKzqbkLcbGg/hN4yEC1CgTL1lnAg7uo7Bt5aNC
jOMYerzzuYKxoTWfr616LJb4lnlGrk7qizMWqqSe703L1OYhUIrX/MJ/uMNm7Mk9
enj5q/zXNk3WIRpjxAh5pIMvI7/yhU6UkNpGI7oVCePRu4WEd4rOvCtpdvN1f7xq
kOYaiKMXOWSL6m9jlHczsUPXM9eej5H0anBL2Zzs8MkfRczVXbWTYcg243APgURj
gvT/JFLXJcui2xppwtMrVRD6clnmbtuiYymyoWLVbpKcqjG4aR2fi4VHU0VmDTEh
uGtwOT6u7gTBKRCp+Zoly80gLm7dDlhdHe6cN14grneiAP3aI9yJGqhcO5Us0qvp
LPmXDeygKXmE2Z09YEXnNRUex9r9qJ9fZtNgoYXdd3aqcaR9e/fmCQ/i+SKgiNSm
BeQTgiB2AV04GwaZXJbICHOQVKp6d40nHrJ8LS35W+/HL+NCv1AbU0Wpz+WUkhBd
GG9NjnmAuL/SBNp36H2N/1eLg6HuTMTgz35pukwBCh7RfM7GJ36H/cZL4UbZ1xXk
z+jOPWmyofNDeGRyHDr+qWkub5FjMu9eMLW1k+366wBH1fDb7NT0mE3EdIaZ18cp
qoCX7oSDMBfTIjZrhGmE8811gMf22Qb0BzRQcvAgm5RYFDalCxe99yeuNggo9Gi5
Cbdswf4BEVbZGQZBCAm6k0QKk9flJ3cGF/lPsT40Zu61b0G+vKXAdBu8nYdYLGPy
pYKi5b2basYOytmqPLY4wI+TuuV9gKloait/p6QN8LUdXv4fZ2KEh/knr9gHqjBE
QkMipNcWca75SdbA7uMwXwKokTNrecuIaHGw8OZS6a7IWVTvEzYc4vOtuEgx5jDf
jUPCsgoczvS+t+Q9eI1tqWncxpuMVpqFPTYj0wMocKo9PmICFeMvmPgu5bTqSfPt
GDUlGZ9MEM6Lasnqht7fUv6UuOgM0aJIlYXzK73PpBqmpicfFO6QoKVGonlTW4nI
/xxWgBWZ4/QTp2e+mjP+v0BGrCeFT5j4v8kfHFSto4Y72npHsJpHqPvIALQxWnUh
6USyCdcivPLKvfDFIpKZxHeMyHKPnOFObSBIgGmRLx52/ByuV+ABmexHGqontdQD
aOIaLFApQJTIMWPWnyuFuzRKks+rAox/v5MVTx4frmshsrgcyT4sauj9Y7PlCJNJ
ekuEqphbuT2qmkteLT/CzLV3aQXPaJNh99RIFB70XBtjxb82nxxFs365g73tm76g
m1/+cNRhzSJMkK1zylSUjm8GkPxdz63kMg5mq6aKU0bq89rtOEUddvoERt90cZNl
zae88QM+v79jfbeYB/x9ov7DxsOgbfIFwHWo/P4scJqXrdbSrn3XelAD656IIboL
GFfCXD+NoTQU6q8FrTVg9P0MVgJYXvxmoH9bsepBgVDQZgNvhSJXw3x8FRPPSGKG
mWhmFfTLDxiT40+lfKn8Go2RLwS8micKDPGPCcKhqLoIF63Wp02gPLV2s7uzl9vm
YrsTDc5bQpgtqkC6lizbLG8Mjx6p7JaQf3RXFmMwBwx7Cj/qjv94YBNLsNEJtwJH
dL3VejrRZvISz6bUAZyj/iUfsA+ulHmhNPDFvrRjndW5B1R9rYbdjCgQfFgPfImi
qizr0Jji9A08fxr1h9odtY5vcAXXokilSz0cIOSVYpGLzagyVCGvDitjWgbb3Mmz
oMR1gXRRhsOxRtREIgpWR9nqGojSiHEiCtdVUxiEA5Qa2Ho9ki4KSICfALnjEu51
Nst6nMIOlFzyWivIyYU4e7pQo80uGrLMmzJEkK6YiC4t6zdvrfnXNRa9Za0tbyfB
v80nhw2QAJGMiTvmdtlg5NaSmx6FS76SLIPilR8nvEiRMIkzak4enqBfKvgVChPH
xkwelbyZZ/LBhOX2SJ9o+fK2Q9N3Qkjryaix/H8R8Gp6v/snoHwJArhbBrN5Uc76
jgMjJKO1Dapl436qUd0xgDnHYRmaaqKYeeY9bOoO+oo52z/OJqSSaOjd3MeqwnK/
1A6xsKABnP/SjF1c8LCGS91/5iVheG0Wu6KcDWmMyrNV+5oZty6xBGJqH4PA+0mZ
6g65kjy/ASnM3hXvveiPBYcX571+cNoNTd2M6LJcUqZl900CS9Hszwi9Go2fv4Qn
DKom0gharV4ABYfMCvPu7+ANujeZDImdXn1mKFV8ZQ5enNw1YYJTRyPw2ALjZ0X4
JGahGyaOJ3+Cej/pFatO/uu19GGRpUJTWJfPfFJM3bhekkbN73ezfHug4B5s4xea
zOn2tUEqGEYlrzNTP4dvkm2Iog6P+keFJ3PQpOXzHz56BBQp/jQwrfDju0f2L+UF
AkRqK6MBj5LPjWg7xl7a+yqsfdkiCSpMur4QP+/d9oUukTHDOhzRp5SorE61vGiF
ebnqdCo801S1TuZzmGZ4OrBT1sdo5iACmjx1jdLVF+XZBT0M/8BWFxJoLKJroU6T
8IzaFk3Aynl8ppRMY/i/8ifLDFkSdYSilAjrKwShQjWBFTsRngamFpo0xLbd7bjE
5F+dYyv/ufXuqXKjPGJYL8eMp+imFIR3/O0L2tZkFWviFwycFFzXeIBdR5H0KgSm
I5c9x9YxcsX/KlS3fVyZ7lQGd0RXbnyi9Efix9A4U5qvHOXPUMLUDxXIE9olLjnP
rfV/zm7lzYa4m/+objlPLAtRp1G+ILH2D/1iPur+vPOYsfBmQvpl4QoUTjc7iZqm
No4V6fsxmAfFl9OgHgHJJ78g5q7cS/1ymgn0ojtYgC5x7IDMWGd4dxyF/4lijhwN
Jz7jPf7mnUjSLU+r/yH7VXZODCvLF4teR3YRMpYtrMPB1wdMBtcaxGxX1dY3kw3s
2WpJPwMb/3NGmLm6u6qunx/FP7UZ6dDAXrgN2KPLHOqvq8tmDy4/XLWTZ/xRyU+O
1+I59YVcK+5rLU1d5B8msFnqJ5QAhDVfF9dU2eK6EZ7Ibs7KuvnsNaWjhKBMx09b
5Cth6smgqG9PW8gXnXIJQ3HNryewQs0H4YeCJZn+0qkIyIguQ1Aaf6uqd/2La5V/
TP0fsQfUM4DMSsG8IJ60Fc3zjYi9ZCjEFR3WYMRCj8hI97eBnt7SiIq2gKFREfUa
2EInqDFl5thyLYOD+Y2bjEn1aUVWQN2P+zBjbU3HanOgzyxgez/eAhSjP9NH8Cz3
3esfIaLHFKfo/7ZEOTw5eTbSN5MXqq405yZ1pO98cToSWaFBFv6feaHLQQlop5x4
8q7iy4lAEXcYr40/pcE9VDESzDdQIByzMumHICVHzVowcKn14NjmZ8RCkmBOlU6p
t8vTJl8aVceIWEBW+ZpxurrZ+KqDy8RqDLxbnlSGb0lBoXROR4xHKKMLc59jh9rA
lIHiKbqweMaXYX7ExG3VnlFx+dj9b755/EwowiRWogjNygs9aDgMOx6X1SLTGliR
QnLQBE8kxas+LiIHB2wzNhgv9Px9dsrROnosPOh7T9YS+ZL9tJGM6rNgz5p/KW1H
TBu1eRV6c0iC15JWkZCA4cSrNvD9t+SoQoYYiVCUVueW6uCA9E5XMbbQdwCAZBW+
VT7mSTGygY0b+EhMr6O4/dWV1o2orVnWDDTr+Xjr7qi8u5xVAEfTMcwOEF3dOf7J
LO0kffRgjXIEejmglURtfi8Hjc8Cy64wsXTfNIGkMPqMfii7wsjMu9wlRLGeQ8rz
+LdeVA3kY0NoS15MYMGwnnIyWNsGMjT02SrJntwtTRrRRmswyIXh6H6PZg4x+frl
Fp589Tl9O5k8fjjUGHdmfTjtviaqvn2LR8g50PowLfZcvfDmQ8MFRQN3uqiCJwJV
xr2K9hu3Az8ZdQXOJdHQxmN7DO3hBRJbvO7Ckb39BwjO9KG8m23hV/cHUhiJTMcd
qJ9EvTI8R4ExOr2ixRm+o1T9wCj+PZ51ZN3vw5dpnx5hVXeqTtGCpQwYkUpJJ4S7
OYn2s89vNH6sMFJSYCrPiSW1/lJkIjXReY8IplbpI6DEuSZaQkSGm7Goo13gNOCM
ZnBZuWcX+FdSfSFlME7e2ipRpAO/0DEBiDbkndEFAdqAR9dtH7hcIqP8LNwzitO9
3iIWHwm/izM/eaFiWV4oxvqYlm4H+TVuPGfCwMyoQMbdo7PRql2aZrCtxdXQ4Uxv
YMSjJdbOmOQJIRUL9wJGnxJ2dL9QB50CpuzY9zuXzU0gRjxgLjQysy74qIDWiSgx
iswumlorioeSg3lRtPz5xVXPzkEYUYSVM95OEN9pNTvnz77dsIBk23ZYKnW8XGTi
nJ9HXTZpKU4xu2xAJhCTbHN2NDjCWBnIEsl+AGb9ua/JL9PLWrd5xLEVWnSd9dYo
98jqZ/VtPxUNU8vRTYhvFeZr93hGeqn4ppYdfdW+ZRExZpwx1P5JNiGU1o8xDhwm
bhQyAN1e2utdAtFO53WhqavizP2Hl5pX+iiOKiiX3OrNyrqs2j9oD3Sj0rM2p+uy
TO7eD61hgRkYjHjUPFpfDnNCH5DPxe5GcfF78fEJet8+XNp8FdT6n6Pg8b3qgpS2
IvUjFdqt7z6RZeUsILhYrXCIx4VbFcqEloSsx93iu9MDiL8NzCBDiKCxM/mIqZ9t
gmdRyEfDoWXDqdeWvycZslfNyUgCxWMmobLawB5QhU0cTZ2HI3Jc389R03im8WG+
Bu0YWLDNWLtg1fsuE5xPh56uB8YvVhMj/HVWkIFsLMAZrclpPJbNTY7tq9BU0gAl
MRmvH1fGV8v0KFBFwxsReRmswAp+BNbnEt9SNoh3eQKJCKF9GwoY/Z0tE5hYRjK4
XYLPZTev9Luc+oG3/ODj7U+N3robQElOtfi8nvnJKbs/d19Xp8KD8YanFhHsd3yX
qJmB7BwuaEnQtG2lbkRvX+RNHkzNZX1Q7ftdKQ4Qfe8sVhxwn5u//+RQj35U1iMA
Z3n+krgmrUSAwHTPZVVVQjkYNJALwLgOOmBWGsGihS2xh8pyjdUXkIC7fA6++xCE
OrN4wIMxNOJcc6Z4bl9gZGVj98siuTV/tSdJH420SuifQuC6OAjlHy6/2yFqIgEm
4DETgwYIUclAC6EXYCbGuUPDdiT83is15ODJOeCrCU2n1HdSm46HG1ju1s39PbL8
AzGEu0s8f6E589DVS3ECrw4NX7C4Nc6bwaSvUi3LSBwV6ciuCmRu0FQLkswrOL9C
cOqklPnUQp03z1WiJIB4o5qdgXEAHlfmmY6SL/rVw9DTmHkK+I8yRCbwTkWsFD7u
6vtjg0OKE3rv14194+vWw3Et9gHiGxibzuORj7NPh91RPPl6URb+z4iLTYAa+QYO
bqOc1UGOip3231hOa9VBrFtqvGNXsASlw4lKw0Mwn7BnhzdqjG6U1hzOlgavgE4u
C7e4ZL3BTAVZy58L9NhYboSKCx2ozxtYBHodFmJmGl0=
`protect end_protected