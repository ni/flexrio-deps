`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
YATj3kULTF7Ty4ORuRfFpnT6YIk4rUPRrM74bVTnc4GjdV8oSnW5PtQkMCLOi558
1V+/wvDfc3y0Z8//ksX8sZm3JZWtrxUppw8c14g9Y7owiwp+JumRtO1zuk5xFbe3
0MMnIxxoTKLhyRJtAxElG8sbx8N21OWDGiOk0Xyd5CqAmk9dcOIbxzMjW/wndBXi
maijUdqS+5KiRCM9+Gsp6k/iEAa2LnYTt4WtjkmDD1P5jZKsiMgFck8WOqLymplZ
ml3TTfn1UlLNm/+zD3SFGP0kABAiUT8NK2xBPQ5UzQ6sMFPd/np8iUZ5u4QLTWOZ
hTrU9OSX7lOvRUo8pJ9vPg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="BzW6NOo8eyBw+CxsNNo4wIDxODIsVe0ft0K5tGuSUZw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
DhjJh9S2BY18dG77XPz3hsiSQ73+w0XqfJhD+f+lIDHHVjOB7CfC8ieNRTexgzn1
5W+qoqOEwenoVQtit9u3XViXJSRJ0wfUC5a9axblRNyD2mUbyfH9+f59nWqGkVOh
ieHxkA/DPprM70F3APxk51m7/gNSLICSvbONgLGndWc=
`protect rights_digest_method = "sha256"
`protect end_toolblock="L7NTNW/5Dqy+2kJZXKczEa3js87UJ8H00YWI+92sDHA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 35344 )
`protect data_block
6eHODtGLmq6ccbB074dgNWpdzW45i5jL0Nzx5wwM+RA0eeOHXxEV143NNyQGmZjT
bzHAi/6AyRCB4X9z0c4MjyrZE8GF4crbMH4T59xFHqVrQ4zXCea5w0kG5yvHgpKo
qe8DCPhYAB9sqzbPdPbHVr2F/kFA3FTLRg18wUUtS/EuxqK7HMqb2FV6b6xPZHkM
EqAvnozHomJ90Q7WSwacK4auBjMm5SyBmkNbskZ1sbRtKnj8tTIqUre9T0Y5Sz+g
TWsfHs9HDqUJUD6YT+Fp/cSTxmG22e95vT7Nm8y7J8z7SPp3mDG2tgb8uV7NrOVe
RORp/ucg09LFSosvIxZHJDA3FMV56ewfH7JmkL81pRmTrto63O3aPWND0fkXfE1k
4zEojVLp+eMKzmtoTNg9CBuPslb11zgt8fGKJvYINciKhyQd6Iyqpuzn+7z8sc+j
vIUMKpmP1tzniLGX/B5UCLfFHPz3evj+AT6B+m0jsN8glSR6G2uWayUISHPMZMOT
wAiq75NGZe1vtW6UIZzV1KmtD1WzuFXS0c1/YyJQztGh1b4wlcFL4+ywUWnQvpqs
yRjwJ8TWzAyjeq7r0kgzBeFzgu/y7+Wi3FHvrvyrMPIWvMP9bAw45LSjUwAO+VLu
lgHWsLREzGvXMSKfXUP3VZFrixFvXMIfku5zGECTwAYVhFL9eiEQpGMW2/BwqH7i
eozITI804lnRALB7YoS0hDv3lOdyXLOg3jOdA/GHTMIim/h1T7pWwSjadtOi3vIk
evbx2rm0dbeHI+uqnMBCDhi0His+4wzNAlfq2Scwk9o8t9IZZpNtDuK6U18C5j4F
3F+8p0EL0PkTmxi3YfzLBMHTiLXTjdMPXGL89bL8JuiGlGz0mSj55OMqnD1JRdJ6
2jOksIDb8iGy5uVrGcnmHxpdzNxxKTia5ihw/uGZtJsPWzNcIY9zPe8rE6sSz222
P/BwOYpd5JRVgTUpUhvhZTi+o7Xbo9U5518rl6dE7o9ZpGVnnG4i/GWxGtN1qkDw
gydz+scY8rWk35SOT+CyqF4U55Nw3nydGnhh+hUdugTNLGkHhDTUEsn0vGauPAWC
H3UYMzOxFk4QmPgAX2XwzkkiHcH+fB/y/LL6beJn/zFS/it4/ezDoSgXueyrQuh+
0GZUdCYSaNPgsxLaJTuXIL/S36QT/sh6sOquH1T/E1yJbwExkfgzcmSB0T6wTou+
yphMgfOxcc8tIO0c32R/14Qi/Wjxzbb72LM2+UbqdS0jnFfHvVTGDeKSEwx1C1tZ
IFUJfeU9O4NeXxdxHvX1m4DCIxfX3Y8OxJa2eUIzVhwCWsmbjvnL6Ib8P4MedPcO
WqTp6gvNMwKE57S5bRIdIJJV4ahcI2Z4YMsJTQOYcpvD3+FjsDZEI/+LZdioYGk+
mqXXm7Q2JAOAv1I5O/20/Iv45/urS1Y4cEYsDbdiITrGXK1aY/Y6L27kzRGWB5Xi
YmspXrdeAnC/NvIrECjIGIMdDYc95gBRJiJ0L4dKDD/vhj84Jt3J0F1tQPAy1UZI
fh+eog8Ijoq5HGVzgQotaclMDZqjdjL9VBksp8sZ/4f/2rEPLylHctyBxnI0WFQw
fbAlYb6CZ+YW4Tq4s1Cs+3aDTwiON6N+vLhNC7GM54eyDUSggCX/ncaTDVW2Ubln
eqvWPSkDfKToEhgq3dltGWbAKPQIxrTpkdmYL2Dg9ofU1eNiDytDEs4ZeSNBQ4n9
AQksTFU4cqq2yxz9JMNmLTcuhsoRJFY5RUggQG4NeSZKcu0kaurUqQoQfoQ73PN2
yNUqqDecAiyDUJhxlq0gcLuwRQwmZ8znfTPuzpgN6A8Gy0NtCQ2BDxxOyEebK/S3
6y8XnfnLsPGxYNSHwe1rPEs4xCpvW4hfBwaqkXgphafPtRHBRRUIkEf1WY6CyYlc
l7/lYOm2BYwNwwCh63wxToK/vOdsbFnK85aPN4wC6pBhWM7sxnqic8oX7hxjDBxS
sxoMZ8BN+7bZJdEjXLCvUMJhbnMXI1fDdXE8ECRgps+rT5x7+Px06irS6RkHdlao
xIHjJgz7rUayvfi9Hk57X+IsOsytehpmS2xHiqFT40LANBWrSaF+CENwOwFpniyG
ec0xuXqRUpHtBesjpwME4JH+AT34eepurJK0CwcZQAR7KBld2yA3lV5cuMIwZvLB
4GpOKyvbcPLskq+Ujm3w6KPIYHHFQzOgDq0/eAJWx96SfsT3OZ+syuzkbNbD4g3f
jHLQOqEx0WdpH59HIhLDQRqXpyE4pDoauSGs2laA/7ENRa8nSTEEDv2aV7PzBr+/
tYTp4Mz1qKGaEmZOmNmSiGDxWmqzUPjIOhm0VdTYiT28LbofFjdzvCfOeY+M1pDQ
IfVp6VEMa+8J29Jg1iDi+w6/jC9+QrOUBioQdpR7HvEfFRCXNIi8atwJaNsh+71U
wVwMweOjpSJfK96ZEMtUfbcCB0oQMlx6vL4erK0sSQhWTiLtRvPWipbpwR/09vHq
yRQGRKRma7FLOJjCHWYzbCjXXNoUrweca4wG29v7VtdO6zHbjsdJd6OJ0dRZTtdX
sRBJbz7SCU0HEBq/8az9oPrmYVXztHcNGUZsmuv669n+4L8eootTYRjdwIQpvZ46
zQRrA92So0whyE6OphkEnV4wzzS/zH51f+OXlSCCqPKkSwu59ZvpNyAzBWJJp5b5
T2E5ksL1MB/vBQ96WiG245j8KflJosI4B2JsEWJNRBaUuCmudYeVC8jT5qlV3Gs2
bmzKWGyVIQov6sZtBu3BJ60hpzTuEinQmlumX8IGIZsQijy2ydEdmg09nuIIumcA
qMQWnEaRDsfgR9pl+W3NVLMRwz1u9Ekoulnj5DICcSNef2F6KyqVGXlkUofWBntZ
ARyL6m9e6tIKHwYudu6T3+k2tcjRfJtGp5UP2C8bz8MDfnGYABVOvPGzOP556Yu9
DGDAd4LqaBApj5EspS+bye8QdQ99NefPuHeeciwa0CIbmckntnyfWNGCfN8/BT4h
kC6mZUJlptbajkZPi0Q8GqpyD9Y1Q2LyfUKoA7OzHsfa0/OE+uwofWjiJfIH32tK
bXjxJaJY8h5w6MCh82AkAxWP7Vr+MU7t491mRH5IQfN9NClx08Mm2jq9obxcbja4
5wGp9n3kcH187SB80HGs8dIkkYoQsMJYCQ1OgioaKE8mJFRIu1Sp4vXFHQlEGL8z
ckcUi13OczfeasE44EIKiZXZwEALcEclF7TLB+cffxqaN/ZKx0nUnUEtgj/RI2QG
H/ReQ4XegMGLbKkIf2Ml4SCxeU6XEqUNAouHsNF6lW9/vPO+ppi2Ajo+RvR3Bl/J
ChzGkK95s7lfuUdBl8EKbLl5INkJabFpCGwj/kHpcrX2xl4SaBxOoHa1dR+VIVR5
wumBxYSAHaC86M1WrHepEYlcXOMRHx0VZPdAcrFnaau/U7wxf8f/dvyjzn4THRdR
fJpI6uXck4PisrlVchVsi2nCAqDlZ9k8Fwhb//xM4PV3VM+YgPGS6aay70P4Mgft
jSLrYujMMM3VfLHlMKUKKIx6QvhJ15DbIaeGs9l/A8/phTbuHUb6GZ4XlBhlOpQx
RsKMMpyaCQlRSuLGRsdmx52pB7eX3qFtpyZ8JIwI+Z4hbz6OP6gGMQrlDhj1wNzj
+JOed9g9dm3QAm0rKmITyoIyZD9YZJJpfCwZ8cK17TaUjuIy6eeM5q4tCM7RMaVK
zzgO1l8zrpH3EN6ebLX1ickWbiE0c+eoxMylHuvCo0Ip218WLiXLdiKWd+EIWqkX
FCpuHm2CPwAGhIKmzzqeL17L6vHHmAbMqjyVXu6KYddQZ7yp9Xx1W5f7J9ooh/uQ
huJzanzIPNG62GpupXTJAQkgyI9sovz8Vuj769RQTIizviKZGxSW+X8cfTZixCBq
LDh+H8TaUNqvFzks2pZllPScIRo1AObgt+vLu7xmlwvnqD5d5b8KwWG0zBFisyOP
aDja5bYvDnhP6Rptd3oGE6CNz3xZUNAfXqSmI4qpZJhBMar12kB/Vy9tuR33pNmx
VTqkXIYT9AmkeC505plcR9rRis3n11eccfTa8+CGajYRafM/99aM69q1tw7gdWNb
rXtkPahV9b9lY5KeyI+t3avRO6yc+n44Gp7FcSBotFgzLHyE7/k1+qcHZE95x3Gu
XByqbKuvi0gF06lACXrCig8bZ49LIE4SdNKkIl2+heBPLmpwq5ySr2ADv8l0Xp8j
WN7Az0+LY+PMQpqNrw6B7DCh27Q10n8fYcZVTt1YaDG4352k2Cw/HdPOGfh8hgNK
S+/CI17D72NGMyDpmGZj/iac7HKz2OU+1A/YCC4B7srNy4Pmp3GkghONLoJbkYnN
tVOvFhM6VKkTvh75IqtWnpkr6e1uWSpzxqqT6O5XO5InQWsAXQAF55xH9l4JadYm
JqMn+TNbpOcNKU4XaM+e3XSl86YPeGM+5/tN0H9fdOgi6QHLZrpdEvV3xP9xtGCr
D+KsJZlpTlwBtG6utgSvcR8pfWTzZZLpFhqq2gGnOSrrLIoYo2tgFa48cCg4l9mi
5vXaYiqLU6RzrujH281TU4aGHeAHtLOOYNaOrBsVgnT/KyXeaQ4QiKvV+vTAK9LU
YRqkJR492Dvog3db9K0MN5/eKO1j0KbENe92edvshX0k5Nx21TEjC5jIG9afW1k5
ZsJSjUQBRiFWzujP+Fo9ukuezcn9NAXFUs+jinbDxrX/6FmdHH1VbIwTEJ+63oti
IVoIGe/ZkU/Zy2oGa0RSQNg3oI7Rx0YtsARSGkWlu7XgsSAZ11DEg7XAjjLSOxr4
VcajGdToz+7mVBqxa5mYek4yqbIxPylfgN4kHJBMBItcEkITqxGRici/3/WFZiK/
mSur3IytaDEGb+vZl1Q6IdcEFrWrA2VgZ/j6YtvyLYgMM+BUPkl/2WXZnz4u0IjM
/c65Co5Jo8kLJmKvVFyV2OeTkeUEC37Nlwz8+w1ud1lHsbUTGyKqBIMM/m+tzCGt
jzCQVv41IHHDy0MKP3xcjBbPSioGzcU8cpGEwcJv6TWh1qLPHptr24G3BPuQ2tXv
nkyV9Q6aOA1bGwoP5sxndgMoxpvXUsiLloWwkKNlkW8+AJqg3eNKsH/1t99QErIc
FD6tThJ+ejProHO/sXBh3IHLiqm4QKajvrLKU7hMgvJi8XZ0Rl4BV/ply393gTc8
s3dmxf5iuXLyqcMQjeoYjkn0BeF/kWX0dlN6+C6FSWxbJ3K46jblHeSvVBfjVEUz
JVc+nSFUfJDe8GCS1UuwiwfFY2MICe+aMuIA6qzP2AUzcT0vDj/vqMcEg4pAHGEc
6A1i9tYMxtdJpSVWhSea5JUV7FME2/oV7XMmC0ozA5fHk0ICZsqaazmzcB+JXMZK
6sBY1XBWvbylx4EQgXYVe9B5QwNlV8cU4/CJyFYyrgt6EgF/J9p6VUn7cBBrwfww
3ZTxXO/3wmYCzTRLeGFHgbnv//MJvmE5NfF7+MVCzUvdATiBSqM2BzlrIHj8rQpi
sOT6ImCVqEmnMgEWA+hxIElE4KLnXn/kK/ZyXByczGn5zCzb3cRtGROVpq6EjzNO
0jHwxzbahMkUR6wu3+9J7GoKzXLPpqg3AqgNY9gLr/EWGyompFUr7B8W2HzJ3DO1
kBKuHVwtVmfQtL1OZuf2gkW6ffU7kNzZcej4Ja3p9L8RJBspLx3P764cU5iiNrpH
EPZEKTQREzTUMHYpO/n31JlOYqdu+j9s8mi2yEKBsvcaRsIQQ1YVRXrtDczRidOj
fQrsiB3wbZhvZouHaCZPMv67Q18uUgKHr4vqRsqotjBI3MR0/s+8ccxlw6FV9SHM
wK8ymOxjaB2ZsF0HbhoP3BtVhDhqiLytbDLYBB9Ymwg6J46BlZYGgiDzpPRgWDs/
/aaJbXOF1owx9b/uCXvLSs3tyx2DsaOPr+461IBgT5oHxpI8NHawbH1MwPYG1nob
kjSdMNq4bim5b4tvd2eUPFMgSQF1s2oguWAgBKihkYjGFl/QRDHZOaRAyNJRf4gq
yZLHvYyx9NQmc2APDO+3cEB7OLTANdg+JP4ogu+fu5duT78jyqIlIqL5gchrpwEc
JQodYijtXbfxOdyu0EPAY5+kYrb0KYtGbssaci3fRCNdfa8dVkDIFOCbVpnkJ5EN
WHMnEWYqRyRPgNsx4s6FA0skN8040wAmEBym6dItRYn9xVYsin9/1+A2ekz6rhB7
Myp19XInicZibC9pxkyn4SP2yZ3UDTb+ks+SPLmBgm73VZsE7W+TPsz7Vd8hT44v
ltX1xjrPhBSjIYeWEnQB4PcFdbAlRxuu3w1UKENl5jtIGY79QJqbVtKpBfFJ6rV8
fqchHJNFdhly2//8pYv0Xw2kOvmzHleziUU1h6w3Co0KR1HA83ZI3c5+W+jEkgQi
jqBv5QS0znaJjO6/eI3gly7kxlbOmbF2AZKmCTg+UtWuJHzeHl9lbZCUux7QhNjH
8vrsE9US89yxTEHspMeL0VaLCfjm9JVEF/Ettsw7Sjkuj5HwlkVdxQLfMxQ3VLf3
XkseRdC7AUF0CYNCb6R3kgR2IF5EC2jGRSYekIZiWPa60I/AIXplb5bYTDWc8YFt
nl3wydT/JrHgPD3X8VIBn3CD214t87x1sEko12fQhCPlOMPp6L/VwVlKSxZQOFD+
6qCp3zBlTqFq+6N6rc8mLcfQxseu0nheVP4y6t9NBVy4CO2HP1Z1IjqI7qOZjpAe
YkTC2YwmU8FzBliG4THQXMjdhoCTp9KEuCR534965FhqE02VVY8hIWljTsJQR0YD
+HWIJJWV+7eUHZwe/DkQUBmMehfam2X3wqmr99fiGfoQpCrNnaU7cK5QZDMfGbUx
sieR9dddOtEgjPULZJgDl4IezV8GYg6dFQeOSFOiVpLFbmBsq/wO/gTo6qlGfRqT
De2ka4pFCM/mfOAJBuIwBoM2Q7dKIssEfDy11xLHCvD1EFls8dFlQbD+Ty2lPN3T
MAqUkG34kWgyXKv5AKQbO5QgD0bZzHBxexFPhAjqnLCGqsIyu7L3e1RhohptX78C
GegsCPCoZqoPxKr82NhyXw/hi3UhKWy/f2u1NFFenIcuj37ETxJ6Iu1gvb0C8rKx
rJoOHBd5pNDEbO4FFxYsGlFLm5C2V3Xz3azgAAWe622VUHN/bd0fMfzjmqZeNJRP
psnLf5ftWvmY44fdWWj+7AbFNelu+fsiMafrzlFeEPrs8RN/ydFNwez39xcUVotk
kfwk9OsaG1oMvB7SlZwN6n3l+AjsSMCeOPLtzHmR/wiWDppKL5C6GI5a6DzsogXq
Z3u+ACuEMmFnNl5uhiN3HsGTAm/DUXhk2Gj4FFKTPWM4glJcgHIYYFac2yAVqkz3
IgUHhnSD3ZDJfLcvGxgpIYjbgM8xZ0umcUhodo3BXuxwlJJNqcE9DwEyxSiXC2P9
BzzVVEb7kFb/A2WhMz3TSmGMenE/H8pMJk8eA/gEcmg2R8zfVXi1eVavOF96Q/IO
Hkw92sCUbUMAIRZqgVKwV/Cx/qCs8ppTLUyl4dyR/NxuOnblU24wwY8Ufp420yAZ
tcPVxGeQ4kuyE1tw138cz0DPSN9kyKV9cWkaJ0g8831tBPMvJ8LtjecElYkAOb0t
PC7UxXXa1kzYJ8xQyrUbDZl+Pv50Gk2xt4/iq3WIxuTKwwxVCamAOu3HyubltPj7
WMOPO2L7JHVOuJefoV6isdU0i22QIRtq4UBV5C73IhSjIObevEq3tZIT3RIlNrRF
2VOLt3aTOT/0VZgkk68Wmj0DeoIgX7dwkuxDLMgF9AB8wfT5AyYtUZfcTqzbTuVc
8eHcqxUiJ771DipVV5Fvp/lTUlmobujOz52QVdADqI6PZ1SKNuwlCiSNZUqjJA88
GUFVBXRyYNjJn5FHjcTMFVIEkvYSxfEpE3HYs0BbYwmtrPiMZWEYXwu/QI1gBYNJ
/aVKzUvZ91l0hSLbS5tZqw8OdARgM52dfUXpWwKD+N1O3t+i+PWaJauWpjs59D7Q
1DszNY6Ho9usaw7Z1Y6hY38dJCEN6XSgAVAK7Ws1d3eV/Pk/qNtOVBAfYWagNDb0
20I0RqGjjcYvSb4LF+VIODKf4sWNsPj9YXaAdvX2JGv0zzByibH02NK+mdTX0qhA
G1k5uKVS4YtF33B1D2RgnMbxRj3+VemgOphM2qctjj9EPlfVjjTxypK5R6YurgUP
5v0kOKg+jGraNmb49x/MmZCdYLWIW5JznxakdQDcSbCef5zFfaCmJBpvkj9qgdER
LR1zBkVJd3JjDTa6oBWloUrgK8JORhB0e4wkVYzm9AwVA9kVK4VoDl+zxImYh7FJ
Rc3bk1MufjczTME1DsDkkeNJ9mDRbFAS1efZvqrHZjIr+IWZdASmpVYacTEzq/Sf
3Da3OnzDDIZmnSmYBr/dfTpaPZsBWclpE40UtdeEcpBrEklsRWvnRheUuu7r0jBb
pvx/AWObLmsaoaWBwZxsFYjdH91efr3nM4KB7EaDIlt5ypZyxaJQeVJcKGnLAkJ4
0qJSTgr4oi1E+LZX4xYQ8GAKuoVuONKc7Zxi53rOKZ3nfo4pYhalC/eRiYZWeK25
JNuVJAoP9Xl6pD8H7gz2Zt1/G5/d8qhaZGQg/r2c457biqnCkKDIXoSWWlbOzs93
y6CnvrzmA2FPIBwUc8Q6QcM+gS3CbC0mazK69VBlNfQZSMcGG7jzpb1JGkVnzv2q
Ydwp19Anf9buAc8ofV51uEFwTbAYs6VZfUndWC23jerSDXP54iSR4RPtyC1cPW97
ViAX8RbdqHoNMaIb9xro3r8czfzA7PSH9ntIv+L/hLxVgdS1kZ4XGwHqsqNwzibz
recTwlmx/uPdBSfQbnj/YgXHpnjGyUmHiCAb0xdBC7xIN8di/7xj+dccBcPrmY2S
6H30AtwL1L3XnjsjkB3mksjVX/6ojx4V05UaiMC3woiS8PO/206C8G5YKo2ik59E
lj4BCVdiHyCryMxtxDg+kRVT72VN9fHl0yeJaXBqdv5lhy6JWN9snZpRGAsL6uVP
UVq1QZfmGtAjhZgAhKjEd1GqIrc/rG9AvE0CUiLEyPgneMMnHQj4XXgMbDsBjInZ
PCPk8vuK35mb/88WyTvbVrNC00bWhYI3aQdtLPKGfiXu+soX8KQKRPZEBYsoGiME
QLBDjy7thoZxOqtvgQ4LDY83HEHtCjY7a7DxWmoybWdlak94SlVNm0fAcx4CxOUa
xaOP3qCalVGmSMupTAqf3BA8uZJ03zVXlJal22qfuGAUCkXKiB+s7wBYdg0wnFpJ
ICfA2NQDoPfdQhjulh8Pe4FGxTShGflERVgK+rH8Jg8zIpE/bI5UNVb9upjsmhuB
+IbvYnnLjFMd0o4StKnrJ9ZXRW/BOE66PmceXHbjbHnPJgaxhM60fIicGVJCEGIQ
9GlW4I/DF+T1JJdI/wXWJBpJm6kdD8IMWM+ETzydtaCfwzA50zayj7D+k7coHZyJ
m79QV6HcwuF4bI3qNp1+1lEWY8hAC3oqtVUfQBhkG3JctnbdaFb16VzV+bJqJIxj
wYPCXT2rveMOahfpEiFSvsxYvEyomycdw3zCjawfib+aUuRqUyfRbCIALR2KDHw0
5UG9/ZbPDR/fZporzpnafiQkVQ1PLugQGdekPqwb0dauBpHIZ05U49cmMwc16bkE
e0hLxrJfH4PJtrzghReqFG8Ab22Z9Pnq9KNCA2HSK0PqbeLNvRtiPc2Ao8OKsUFY
EM0t5MEodRy3IKa6bh9eo3Q0BU8Iuxb7YO56Ax+sWUiC+5s3kbZUUySBe+zQbhcK
SdwwcRIzrSND6YmYOk2OhHSe8URllGrXUdebXj+/OlECW1Qoz1Mcuz9cov5PQjfA
xHfiHnXHHJvAyiztGPXQksoOSAshHbyekQ9Wn4RRWR9X1I07ZI4pDj/j8toYAmBy
Ed6vPnRkwfb5kXfjd1t91v6SYssPotImxmGEXOisdbYtVieMB6o/eSggtg+0KKMN
fMMTxJvfEUCKSzwZaDrGvIgxjnqZpt6GuN30wxucLopzNRR+xmsII5F6UVMl6S/l
DJ2FYOwmGnqFGBoR5Tso/PyIcz8Hpdxq3FY6RlJrtOMgNpGizP0HNyLmg6S7jzJW
t4XOdAzmjAB1Y22LgYUfq96r2M5gGiw8VEsVy7cuqXgiWTvPchVvaSY5rg6cUqeV
g2SnZ3F597CYJH3V/UEUYy5YxwwWqpI7LmXiGYLutD+yyA6dy65ltRAbxYQ1nqzH
IlsT2sj0uhGnF29NycIJPkjiZPtgtTqgj6dG0HWoxeE44gdnZxXA4WHrf7wQHi+D
6OJOl8iK7thCMwrA1T8b4lb/1NiaImG+FCDE/ROBQF2W3OFK1jRLE9KKMMcnqwev
OsL14Q6JpNMjuUZBOf45nDHRR2Q2FNUJ/e9CGks6q0OfFGI9KUynmfq9P98wmw3I
dAo4FZ+Ewz3dUxnggy8XljfCCkRH6B+Y6LdtOuX0wAEIIN1GLN41OOtlKIaB9hGX
wQWBab6vMzNmIJXt6Gl+yIGjfdWwBo4zvVyQ18DR8TD1ee0PK5WjfvVNTiB9ThRm
B6oycLjeeMiErnGd9bOO9/FzhypoxQoJ2IqjdYpDTrex13AJNtjL9y5J2ig44Zrt
NngCjMUD0P780Cb5bmPlGuaSqn8EUGuYuSZPM6CvbTrHhqpy9QNPS7Vo2+Q0JFMX
l9BHC3F51GPeGeuI7RrTr1qSq4d0eIH+7rDNg7KLf3jYiH+4ep3yj6HNhcmPrVJx
nr8XqHZY0Ob7q1n60Y7uNCL6uC8x1rozOiMYYzGlGTBHtnL9vgJ7nd08cOQJ3vJH
MTCAFDoT9CgvHSBOOv6HGnMXHh3w/RAlz1GG/F3hLhjspkqiLbNcO/KexS3rnpND
8D6+JiO/BdMOQrgsNcQu2UFrbCii7/GpNCjuXAPPubaHXezYNxRpym1439HtDgxD
w6p77d+fg+SdqzX++RABhYymj+EQevFPa2XU4+LvMAI91u4DJQezmi57Zr8xjbTF
g9PlEMnvrjhv0tIt7BG4dHANr2aEobSU+l4RWsf3wUSzmVns7i9nIX2rGgs/pjwC
YNOlfAZOgbF1ClQh2206N1BRw3VEsNMPyj0SF/NptK/j4GopJWPLbpQw5900GqVw
gCclfN1t2tFYJIsSAaoCXsm5CYO5WbAqnvrVeD31o1E9Mg0pXYJVU3Jlk8v5Mwip
VYVE2wgfFFxkSXnO3OetXruQX6ybVqLV+ZqYG/TlY6jz85LGdUDyvBfk4RHVJBtJ
wCB5dOHwyEfLVWl5j/3rX3Lbhhl0khkVuzbhal14wPBTZMf0RHsAdIyz1YOmnlox
7jrp+ecivjcNjYyWLeV8ggyILbHa+CylIX4G16bG8EMz7H2vN8xSILPGAkyStWmn
88bUNUD0cGeO8rlCMKczSU9t2+EHsJIB2jAgSWmj/m6c5qdZ7cRn6QZ+sLfShzjz
qVLi4kkyg6Ogp7Y+beEfDdISWbVqV2hdY4sESwknwTElp/1iT8yq6FI+euKMYreX
p+Mrcxu3zzVHGe7A0pB+x3Uu7qwSnYHc7oRczNgg4DMlk9POHRLbV+lOKop9yiyJ
3lN87AHhWdg+cZ78TmWBe9aYCCmXGQxCC4k45fVuKBX7nKbqRSr5ZMZT9nc3gQYk
NLkZLXtKBnMitOuk8VnYzIsOaH3g13STxpCc9xRFmWfTomWQ0mNUq2TcBowcrS5j
3m2NIJMfhK7GcorLasuD/th7UdJmMGHq2IhYbLtA1qxZ6LphV5wdtSPShd21kl8L
s57s6v01a+G1bqv5rwuj2zHpfr7nc9ul/dRQM6EvhlODFxZsFvSed64OWsFWMOGt
/dHtqAQoawu5MSUJ4as91AnFnkCoSBh7FrdIkUppNKMO7EPgBnxgl89GIGbkY0U7
9bkCSvrgiCdznK1PYoIynDDhZHBu93vku6lsS9BfiIjMmaQjFSMM/TvMr0JN6zoO
Ifowfvbnf0ZyLmPSJqRUk4zEd4M3etgL8AVK3Ey5X/LnHvbUHsepTmFZWN4ewXaT
FIKB7FDzfeQbSmfIMiHCv9ng9uAWrZYu2Iq56bBMD4Q+WC9d/I2b+rpLxRT6lhCc
/GEA99MLrq6SpmOByCg4DUnx5lyx62+PMc+eA32DTMiDGMFw+9S8sri14KXrlHlE
KROzSNcXQqQaiRsCFzylPpADxnXYLqsV15l8FEVXUIpZG1nW3x3Laasut1RcVytI
DvDmTIj56J1tprrYmL5/lIWNR7elD/kkVWsGPvWTpyyBklx2qs8VBzsoXrLi6OyI
TS2xsu052sW65MHIQ8EKbZlqHs3gK+LsHc+1MkN2HZIvNBT1SB7b/jwMJPoepVRi
u9Dam06dA5ML3UpJGMzDaXpcBpcGjFfXmFxKrL95gswJWfCxBAM4PZV2uQhqTe2D
RrBRegXc/U5HPdyHLe48V+wGfCEJUW/80OFcPpNJIIh/zW4FYSAAgSWiDlBGHZSq
4EwHOgyAuyzsHPw+ou+7VJ09VaGruZetUwaWPcf8FnxtmOMHC1+ePvq9oIuGKlzq
gQ9bMBvHhTHYKdnFa4hnV/SryusNjDnC1ZabJb/1SuPWcn50YwJdQcfRjd2+FhA/
TFxD6mCZfA+pA5jYtdpwEAVibVP/AeaVwZmd/Fur1hdrwCGms7W3E1TxkoPgqmGD
CSbjg1JCnrdZZNVL06+4K8Y7WsE/fD+8fL2beeLXtOC4AjYPUTYi1YPQmfs10QZ/
UDhdTAzjtcq96aG9fqGIEZTyHcUnTRC4PnalOfULxxNNNsWpzl78p/XX+b8pXzmC
DKh6iL4yvFx9iEN/WFjG6IXRmPMj7ev9k2Fk1It8maul+Ya4Tba/BrDyq7SVlsnJ
xCzOKmN0FrhZw+RqQrAgV8ziK53GvOraVZjdHn+LImUeplWE6kJOMrcXDJyfsZl9
nIH/mnAJfnA+WsZlM0xCMEmvNgUwvfIeTB7lSIBNuA0KwzXiHZAeFhg3J4M/AACY
JOhkAYtM/DjpUamN3medwtAX3HxJa01tuQHKHhsECF/fAzcFFwbm0CzrYXXkVC3l
u+A0CsBlg/sB0SiXZp7laZzmSeIO5jVcy5ZNDb7T/wcEZ3XD6ReGIxSaIzOqxaLT
GIC3xhLqtHhzwlZoreeHVl2/Hl8nwpXoQfyRk6NJXmVYMl2iR5302In5IG5vZF5K
P11OfN77Vi+zF8npLV4pKugsRUhjlqm1cTRNILy+2gqljGMJFe3dAZoUDXH5eJ1L
wfEBVqvQot43PYYE7NqYDzDvcm7JPyDCKX1zCM6mEbU3rTpN3pvKs/RuHHMfqh0X
mERmEhLVpGj6pIZPaeBgb+dsDnGYv8DtmBBVLsw4myBNh56+rtOf1mgIzOwDrKTG
X4VlHvpdjVawVJpcCMxSM9bNoh0ywlj//OLj/6DcL04v5cKOHY9yBoTffAEH4/gz
yHzyV/F5HX27gMA8UY7EmIMOwS83CYOJkFk1qlB6m+XCTi3cs4pSbh7W5PitiKlI
hj9P/3Q+3i5Ma4MxCsD3Mbj9xluR3oJRQy8UDhUQFx38n7RvYrPTMkfJEardGu6W
h9DQrETtpqhL5joY6ShKP+XL+4XNdYmH2/h/GnQmX9Iuo234Bxjrix64ma4Ih3ja
DFRHXRtF8L/aNUWNnMLvS3LKJx7wYWi/M6iEV4BBXXvRa87Ou8uNXbfHsdwiIVzC
Zq2aBTmG5bDWhTr99+MRU/fsmdJoCMaqyfoyW2DIWGYMzRpoX3etdEB+2FWntyeC
ZH1cgIFF63ldT2PPljCq7VFtV9JrkNKerJ5cI3k6pXFstbmQzhnqBm9s5+8bXHUM
OIyqDjmMxk/DJ0ThYPrgQH/BKpFvq/CICDBd4QAvYyDbrKCd53S0Q+aGbxby/9BY
F2JpWBxUeNrH15XRSaIWlAz++VsEAkcX7LYoMkJaX/6VkBDVwbopk2car2UxCJ+K
9q1utobPI0R/onVKLlonpy7CJAGDeE++dTeWF7/ZcWM66aV+Dryw511q4zAdamCZ
aannOibdQu6XjUw1pVdlcY3GgsnBYpB95vg38fieAAzMteJrQzHZPpqugzGlyEar
eKJuZzyeM6y+igo2wctWtZfSNA+6PlhrSPi3rxsWh4Z/RfjUAwtDveQMtvLqOgZF
KWrugDt8l2z3O19GnzftqD1ZVuIrjSLmyb6G/Il03l0gQwHRkxdPAKU66sWdDf5U
Zlnv0Uha5jk+j0v91O0TJRNJRY4qNjE823ZO74ApsUki45LV9D+e5P0/ZODoo/A6
MeZEUSxc8vrajVx6WeZz3lykXFgYbR7n+8T11EClkWJS0ta4Z/JvnbNW9SdjVEH7
tx7sWKGL++3U8o6LYbwT/T5g+vWsd6JOWfL/i1gpB+cDs5KTWaLQtHOcroKvpKZ8
CLzRIOciWh3eciHxq4eo5hKjOhvTiSrGmhfbNYb56WWmrtNoZG1k4MBlIMEBOPIn
7BLi3RtCKj5fahvgve1bXx0pnM+qB5PdBBqg9O350qC5wQOvTx/ZwbxI9AQmR4MV
vbIzaKWAPUu7ihDEdUWquHf7r3nLtH9HHGvbj76ULDoIy14mb6oGqIH5y807TSxJ
2d8J3tV5KpUCBrHRF+LXrkJfgMS0rMqmpr9PClgwl5BoS/6Ks/BOOLvJ5GV/5H32
AqqwKCuGB+sZotS4P96S1OkMtexrlTxBZ77ltAGgStlsR798jIFDAQvn+55QAKom
Gc2typmZltLlEGh7GaClR1HL2YwqwxA5d5N1rzZ1njcFBpbsKLtX+UnGYgTRiUjQ
D71IlCzOxYnWwv4LIsbQiob+ZL+Z+Fl1odTWVqgybTK5DmvMOaJLZUdKiVMHuu6b
33+Ir5dvHzwSPzsH4zQn3NuteggtpqMZ9IQPCbMNknFCrQvKCAuNpUh/HKsqw1HB
xAHLMJ1zCOHXV3Tr3D5hCmbNZzU6DYAs5ceEEHjH+tkjQYCz2E+ZYqWwoSSll6V+
cW7zWeQKb2nklSqa4wXUUDBlRFRgCmE1TOmuVg87+tAG8g4effPcJHyZYidCqJKW
kvjYOThBSkHEtSpcufYRRZjd3Y5QpSblP3Tm3GLnLtOIXjLYep7MFYCs9kSTLw7u
uTlJEtAXpIGui41cXzJ/cWgL9jHtESE7orSAMYST5zqxLpJvwcqR6xEpim9WYpia
a/6qRZU7soxz7F7xrwoVJcNQ8eiwFX8JJSbNz/bWUtvMFQSwPWGeiYNw/SVUKeO8
l9U8aFzv1v9hKYwVH411yZcH3DlNgv5NMHqoX24xIrI2AX2nZUu6GuqURpBAzz8A
NdHdBwBufC2ilJTZ9gY0Coh8KMzjBiew/i2Jjbdvf1Cq40ZYFO+y23KUizZaAyCX
V6jxFD+InzWgQ4kLXYGwLUDeI7KLiF+NUZkeRJEdgFuPx+y5D5WnylggyvjNtAR2
dKnzucYSAlE6INOIisPPo8wDXHUPSeSSDeHrkqOBTAebtv3mhl8r7XvVVbiRe2Cd
Ff38KRemcBq5zn0x1duTfbBN+hlPnAWIeiZ/helH32ORxe9V/4iq1LArFfSgnARu
9feceC3uVPiBZ3F3888oTwyM5MTLljHLrsZ3XassYujsydnA2fH7/IC+fkh5hfsr
47xAEBz7GfZdthkN9XbZcW8oBp2f2xXejtV7JRtOyDbsNm6dkJmYSRlz766o/eLH
9ZByTUBmrX3DrxhBdMr3S008nW/C3m1aijyZ9PPVjdbFmZdtyuwECHTY2f2w2lpp
PWX1XbU5RZ5W4XkK0uLXOsWAN4l2dcdQ/3robysjIkiN5YuInfP8SnVheF+91Qx3
NdNbXg2DZcpJLuHc+wtHqeAkZNbu9XDiGmI+IPvvWiAq18+QJHQhllcBKkDuaOW5
kLjm7pGOKJ8AQ5NQ7bu5B8YDXmhbcNgvCzEK+DrrJJIVb++ftQBO9XJV7RXbO9NL
hpQVQIJHaBG7tLU4h+37sm9ZBgAdah+kYohJyTnN6ZIvlZjStIzD+Fw4o/piR+6Q
hPGAWPuWxEdKCeTsOvgIGOecesNCZGAuUAEJMgD1HwmIkfbujqaVgrnASP4HEUST
vd94Pn3PIZ0UUyaSH/0eQugj2SOBWn3M49KNLbFx001MxCF+Lc7ThPDaTUxWUq3p
nJKAeNtn+UBCT0nm0kIU2x6oV/L52onOWhIAeqkg55kG1piykkJRGw4pUdBEh8bo
jGLWGqesNkqXrepqJEhkkCmPTZ1bC0tLrUWfU4ZQ8JOgqhOHZIUoDcMjXVZPLvE2
L0C1mmegXyziCpQ2PAuGNZER6gdo3rH8ad1QXlhom6ceAlRFf2y/PUshN8Xo8zVP
b/yncl1X0BOlwl6wEccm2o8aho/3mOLb7nmdI6euGMjxZnHlromqNBq6K30PFqpK
FAlngyFCN0Cgpo+ugomiOaHRoi4yImaDeEs2p9RiNqUyyK5+8j+gqq4WpQnyGX6g
VYnQqVXx+V36JRZfVj+SEpr+qfmpdvzr4vi/wPxcleTWxRxT3JHULS+o4sEFjk1y
09YdWnuh4obuHj1KxYSCR9v3rymnlojOHEGhuTirzQeBRzLD8e0Qz/MUlBLPXENY
V+Sf58sz8L0g3sglk8Ljs6UE8Yi8Yzgo4MwZgTk20J8SiHuFlXGMlHVJA4qcK7qr
BvTlmzFnQS0l9iUOxoO5b06L8i6cwzwoU8XXvB3uovuF22CCaLbtOzBeqPOWUsoC
3gruzgFqjFzjCOCHZqMfz6tFeYBskPSLSJbuMghRoiLh+wUu87mex+GHW8wZ1G2y
QJy0BlzuqBF0lZJaTq23cJw89xb7B32h5wImPXK4QOb2lYUvJb8D6ajV3Qut9LOj
tpI17pbhy7PAdQ+5Rmg04oT+gek3AskPxfZKha61GOlwEJF+X8492gR5RqMzAeXG
FP1qH36IyrD8dATEYRzknqVS1vPSTgxm7zSjWExZCfRuU+lhlEmYqw/8zf7AXL+F
vub+XB8+c2OeZZc1Lh6wg64slQkIEoaxZQUO1TS75+wDzobDKMkfVFIQq6N0qele
vAwnn87WJCAi7voXp4VmsjT8A6JIbQhA+W/pN8c/Ns6YTi5bj7mx3Po0GpChaS3r
bv+ZOuhJZPdOPWtBMZdFLgzr1j7F2QIX0ovy6P9TuFvt0FGhoL3CqKeoPniaFuCI
l+RzCtdLp2q5Ru3lleRNCLgzS4JMhw162ZgThhAGeKpPU/Axms96jbcDHNCl4EAr
saoU9YfTGa0ccsdzPj0Hv5SIdAMSw51KnnoUKNs4Xr5n3wgo19tB87g99prdYkKE
hJTgNqW0ptNukPt/ErKL7KnGZZ23a2iXPC1fXS8K5dUZWOQzodhUgwQtEaHeGEFy
4v0NHcK5dDwofkozZT+jGa0oYrEuBRGGpaNqMe89skDMKWgsxKdJjVTIhWY1AmgD
csjkDgTn4ApxK2noS8fduJ8kBA5x6EuXfN/HyCJ612MX+EvyQzw0uwUJpRUG2q9Y
Hafm45czZ3k6nGPAbE4wjkTHn4yY2JJBJMMzh/9NhCiCVGjzEjNMLMwGQi4c0RDh
bZgCG64XvW+n3imkGExVtfLEUd4JaZ0624FJaH1qxjqbDMM3OfvP1X3OL7R2zC8D
Jdo1u8pFEXRGrWa+/1nZzSekL655xSuUgh6hv9spWT75neCktCgmf+I5oJur+cso
t4+lvPm24uU2wzYrn6eTlgym4MM0yZSRqwiMRRp8ARuGLBVUWljMy9FPnHLNEWH9
Dk4XG0tD7BGT+8oBjl+IWMF9+1GrRPHbUS1Tjh4h4fkVo2NOTjSUJElamD8rKdsm
KurAL8x6VRVofn4T9+Fh/1MyRLbsYrxMgnZv/0UQmiYtt7mzo5EFpswju1DqUILK
4bl+rhEms6qTsIbAhHTeW5+QJky81KPE8+BsGk8VOV8P9iMJGPiPNFlvWz0ev98p
eMi/Wc6SfIzVvDPYB2HmStJEXpHKewMPcUTGkDNz6e7dsKNc/YG1qSXENrilTrfr
q80VSkEzj1gx+j/nTk47VEFpqdcboIyvpJk0OC3oaGObh7JTD9D2QDY7VethkRzl
eL4NbWbvzJHRwjS8gAgWWPb3O8ro8RfKk3M4EqM1w/+ic9WJGNeagjFthmAgFc94
uyoviG/mtyagjgY6XGnZiB4P/dzi0Bw5T25jS/HqFGPB1qxubkuyOp/AvvKRpg6/
wT3Khk4IdOBGDI+ccz3JavUdih/jLvv+bBEELxl2UX7LRvbljzjcX/qRabEEz0sw
tkXyXRgiA5KmkDvFFbXWyVqXr/Mmt31SAk2UwcE+xaFsynst+dPrF/TPnP8NKJlV
zFAlm6pvi5Kr6Au2gxH54HjqHKfU+Gj/HrF9iIwMwWeXPBgwAvIwZ3nq7iNFzgJy
NJ+Fn6B6Q3EnYOSJZbORqm7ztSXtH5RI7uyj5lp7L0C7XF/BwXdQJmsUGM7HEWtf
CTiD28bMkzOeZ/6ySellrL7jrdQx0demteN+7rQ4Z2gcmoIYO+bBZ1F47IXYEafQ
sdUCSBmi0tW1sgkqeLKjGGuspUwmzT7B0c5nDKtDh7o6V0DtK3K9mXzjD1toCiaY
HiNYj6VdA5JF4XkB5/2Sbadgo2IgmfTX5Izdejga430LKKwaVSLnS5r86Dkgribt
jq4A/X4G374o2WMRd+o/7sf3OWOhLAP9C+lxc1YP8t3IM7ElCc8G6woChbPFGKz1
mJempzpomdeTm6C1Km17tzYuPcZmyweJlPFMKYbKmYcfEzLrA4jgwe02aovFLFdn
yereRFqwIuE61BUYaOtVYaqZD3aKiAwNNMPX+C1B9tEO++1TnKfwMDl/XrVBC+Hx
IG/OrcU5LAb5ZucVTA0JdXcvezNOeEwDgulY4yvuKHgrVKWFUo1HpqnBO/e7Ihhx
9G4fNbGXqM4GpZ170bzxA5jioAk29YleFLM85a9vD0aVlwW8lYj2kCHFzUjceHHx
Xtw4TC+FWStf4I/WmTrEM4z/5DabUvCwBt2G3iZHQPFGQDGzc3H/hVAr/HJTkUzp
V8ISBedmDqvzz8rsJojVzzg31rX7R1hVJvN4YOtOMoqo1w8ivxttlTCyeamk+vOm
M2bkBm1yGnl4eNmE/T5uJPtGUdxeFcJeeU9u/PTh6ZHo7EIf7SfVGoSiMSyvKZww
Ehyvr0rA9X5CNC4XQK4nc8u1t53W90K3LQfhFMOfBiwhhdJ9nYwmIXZapxZVcM6E
B7iwwlgwU1c0bn0ZJVQJ0AclvofTySRCREPg2RW/sJhnHbYkbvvD35fm+7oqYBnk
NJQTYU+oABmd25QpwWit72C46HWIHiCQxxdKzmPmx0EI4a5gi2RkG3iyoCjzGh1u
nVBfyRCFCupzrONtRy8PRLZMRVWOUrgAdd0A1uULkQMxUlo+bMsrLcGtWT2W5T1N
RZJgIO9X98vRtHspaf9y6ULqze1AZiz3wq6hVxGabAjO3mo9DM5vQBviCiAyKJxk
/nFHkWYeUKdNUsIUfecAtDNGS1SOPN2MVxeM266rrbT9lcKD7ZKUuEjAey7k+q//
myUIDUNYwCp+qUdmmDgfizcbqWqJdVtXAz8NpYzGim19aTFHatpwXfVU8ffrEc+O
v5jDC80ITjSrZSCUKBkD8+5kVC8s1NhihUVC4NDUqXMOEYMntlDPn42oR74H/nCt
128PK1Ci2abuDZrh3Neg37QK8p+hZwsQ4+XtfeiCUDQZbpGv2kk0+FfpEi2fEtGO
0nFL1hnaXqqfA5ZsjjmkWAny3oB/p/DYA24iGYUbuvgxHM90rWsJ5JEkd0JnNWnY
zKhzo3qVC/zHPZuGmxeQUKu0xoBdiQqJWb8GlodlNRccMMt2X8pzQ3LJxEF/8MQb
WLnlJ8gMWtIvrpOHqAj+3aWJoPVqdC56Pk+zRLP9RgzCy1hWdYPowtUKFWMrz2LK
ddtXIZ1jijquWbwQJuBPOfh0w3QIBPudPkfCo122yYSx4Jihan8VQ9KOAUWQdeBI
DPw2u255MFGA117ytmaUhFsJOISDGBLVEede9oQLoLXVmpjiAcA146I8x8XSS4Ns
2j9DCi99RlElTgWrlCvAKRBz0KIT3FrC1PkiCiTRjngSCgjwENT66DZQ300qqxFo
aeljzfFGyT1zD+UpYoX8BPKgDZ8B6URrlUdtsRuqJFOpG9rP4n87EQdfHn4wArCO
uFH1yP8ozvGk7IFMZ0B7NKtW2fhjN2I8N20RdD/mwTKdWVfI2x/+mZ/mKjp6O/3Y
CLoXgDxUWb403lFAQswkE1JtfvOGpR3ZYXcUksnnSoBn6MHTtnxOrldXDDOFKpww
BYnEgZXfW1t+6dVN3sYu3D5CQM4a72/ZOow1oj+oI6CC0BikG0/5Qq+1VisrT/Uq
ynbus5fQS3bdtEYunVNc+1qjwMRRQ3RWuWiiweJxoMiZh04QwYfGBqE5tyGvhznQ
oETOqy+XPY9Eat9t6abj/Kgef9jmhV13OVDPFEAeXnOsD+1rXBvhz5vN9Nh2Kh3y
PrU4YfM4S+LjykAQWWuBXBbXu0jDQb3JwCHMfd22z8pwN83qjf95MtP3KpDhwDBg
yLgyGP0eMlMVxlcs4ha2SCjGb2SZGAqR6T1r6qjapybqsVT/+vWw8c6s9KQl0/Gr
GOvSJ+KUAaB7udD39+JN6ldrx3nnoRaGmCh2CDh6CWkUrgwMpnY0LQEUlholNunc
TmQVQm3zDWD+mwzR3OqJWlNu1/PnJJcY7ynuiuc4AoSHeZ8Qb0pBI505gWbtZd9C
P3ntfMocn/n4oF7YIuH3DiHQ2YDBMwzGEBQuN8z1C4D0STDX0v+gIQyQ9ljTIn84
+iuxrsYUwXC2ztQdGcIsbvsCDAj62kZ+r+tBgViyFIW1upGzLtz/Uof2O6j6ByT8
/5TNkPl7O/4ILvz9nH1tXZF2KkSC0lSicr3e7aTW/JTHlzDS73BiQmD3wkE7RZAd
u0quskO//3fkrpJfPzYhkGw7m8TpX7yT9volKM2U72tPJ5O16H86mnjPvO57Lhfx
xceqFRtniQzOmksnq5SvCEcegKPHL6nr5bg3doc/Sf7rF9FGyr15yz0UlM+sRp6n
3VQOh+m1BuuspYZkSdgfjgM3iIpmXgd/IoW7wrOCqXo/mwyZWLQ/Y7ZzFGWa20fK
s2FeuReGHUZco/zwoSuocLahFQuJ850qCLkYUiTeDNTzvggqVXNngflIDC9IWC6H
HWmWzS2BDFRt1ks2BytZG8FlMiQ14EkTxBSCthNydgqUIxwXcsRemwkPKoYxolam
skqnpUYhB7tl7rmgwUvE2o03xk1iBHhku+BTz9YdZq+n/F7NmkZficRQMzMiyEk2
oYW6/5h1AZYTk5FyhLlN2U+DgApIpSjI59QSu+nfrjEeUcXFds53Ph1l75N0mrM6
V8/hc9cXTdeEt+osgQRFIvedSHnxsPtxLvZieZu3XCqA04S/jEHOzK6svMMq0knn
w5c4WUIyq/aGmzP7dqRGix4g4O5bxRIaHRC5Uiwrav1fv9p9/cYgeOA65nf4XCuV
gaoWeIE5Awc7x1BSC7WiL2koT1myFuQIoTBKEbjwcWu1tB1MeF9ZGwhQ92/z5Bsa
CB7hJacOlHDnGjOpqVsEQrrjlcN6cIfSYB4R4bCDfVxuJ8EWmDd1ZIpi+POogxsr
baJ9qkErZSuwnsdmw3Cbky0qWVOEOKZRzWDRNI+TPoa6ZaFQ02wTBiF9tBazuM5M
/yMyKKsYk8TUkxv2XhS0Uz7zIJmfewqhTyBgj7zMQUOe+msZOdXu+sNEDvO3eCX4
/RwnIC6WKHZy65QDBw4T/Bi0ufGiXdhNeByyRxgErzOkJbNAcjSPiATN9C286YRo
T0vE9mPJqbawVxioA3YF1DMD0RoZGMO286FHb4JdsT5YltPBIc2/iF+ZlYWAZ60k
i9s2EdoES1ugZiWj+V2wvfLC2GCu+pmVYbzJPGzXqSsYSyuv77CneFu7t4Djd16a
3lpw939LVp96mWdnkPczjqVGukOpTfMmgI0IHiQHhG8fop3/G2XmxmQR6oDRAKeJ
J+VIY/lY8b1klUpj7ctdSPtvp3UP5duqTM0F3uVAs5jYBp0yoce8XCu+teuLwwsV
enL6WNUsqc/sAGdW3X6a1UUCQYb09KIc0Ap/UXuGPn2nGZWDcfWqPGiBpNgA04Bp
y8kaQ33pJGzbnjimQ4dG3Y7CkN9KbfNSyBvJ729DI6LhwMA5f8H+qujQt2qxXEtZ
vLV4ztRKvOt/stR30t1DSCzylX9XcCUNO4ajdRxcV5Otp8p99pSM/VHhguw/9qNR
b5SpDyuil357oZj8FCGaRsD01EJCGA7SpLyOCtqDeCVaBQIshNtkpjHK7W3xTYxC
5PtQe25BQqh+D25GBg6KUGv6D6yUuuEKjUYpmiy+Xw+SdJBvU7l/MlZhB3J+0ew6
yVwpAT6zXd/psNxcwITBa+BqixhM4cy5ARZk5pTFv1A3c/qjSV52HclU/XdPWSZm
KQE1aZ8bSAWcNM25Nay1guHON03QzGl44fYBZwZjUuHxlVIyRUE1Co3VncILAhY8
1IkTBQSrTjJdt5lYqmVzA/QQCy8Zq9WKKlOxaKtA7yLyZNFaxxxv6U1xspv5RSJo
YVkLFlx+9xBg/LD5P5s6fDzjbP6/BMT9lrtF/dZ7XzhDMOVcgFMAzcoZz8PshnI1
nVunfN6S19k3vzxo8+irLjLYQ1BCqdxVncPMJE2cxuzTf+w//y03XOnJS/ubaFya
LTkFKICDfzjrUjtCGxhO31Hv1/QA96Sj4SbZoem66nyGmctXz3WduKW8fdzEITFD
0/nqgDe/Wque2byDHSig098p+xwB36edLqO4OYIWHZS2MUvWBatCYjTGM+WXX6hu
ZAvfGQwD4iDpUgWwuMi3IegEN9fYyJCO6qw/FXzeTLu/1JD9u2BpWUrKGVcUksEk
Tt5ey3/tTPrFIVkpP1C0leLcvJJJtcK3W4BndJqZQnXh93ZuiqnOpvZMKFtjN8Cw
DD6cpQyeHCe3YM9fN72GH7KrwhBuTJXBp9MKmyyJTZULnMPegdIsKy/Va1NxNToy
Y2SQqcelUapHJ4OuoSzA5gk+fd0NI/vZkyUZHYuJzC/wc+X78arnG0ieAWj/AHpp
JB3WjSLqKrQn23GSMCp3/RUrgJqTwbdyl66T6nGhUxvuyDhmHHcKaxkR61QQUWfE
IoHniVYfhNzUyxo7+foFQXox25BEhdX3pgM8hheqtiv8cnec8SNNQ/aoQrPojRoS
QLBQYgFB3zT84ymsJGDTKsdz2tWZef7OvCA1SMSd4LsUmZ78Kp1Tw4vMxuCeCOgr
pWTgiMAAJNgvPxDKptt8phqilKjVTthIy5kwkaDLNU3B3eDg/ZMve02o7rQIlCFN
QtY8pZ30A/DiVkYHZTnlkF/QWFL6f6ccN//EC+K+sHwjQx4LqN9EhTCvMIHWK2oo
6UC28ETanXjlre1+QantUOaUzXM4zNxqW6CVOOj6xM3HKp7JfKLpXXvmzxudxGrt
q1bfZBCsMjSSVg2fba/KZqWNKbh96SoR/RqALNFRBPXUeSDec6gGXDcJBjRGLNTx
iZdKNjr5UHgp4t9l0QENdd1SIZvFq8RbmfDl8tGj5WfV172KRZkczAKdyGHAyobq
PvGhUgQFAp9MhI+DTS3MT8FJXPFWbS5DH56IoEe534f/c4aB7CTl8ytwnbntgzZQ
c8p9HnUgb0bc7E05+af+RDikJdIjh0/2amwbPHspnlyJUiGik8J4W+xReYQ9q8Ly
cZHGDFYotgIZU+FnbPQ/7fVP/4sO44BlBt5dsFYIT5c40s9S5mbl2Yn98Tpma08N
z4oDr2zA4GlbDcSGVDLJ/q5XK0bGKQdR8j7k3T4bLtX6C3JFA8gEvprTsKmxA+4k
kogHApcGAxPlWyK69eOS8FC2PKuzGAHNSYaM65wmXOkrzu+Vt7p8FS9jyuKNv/3/
u7AmmKpoUizVTd9/2tAue1eZgiYQq55pFyVaOv4qSan8qcSQuKr1+h3wakRxe7hb
+pfzSiaiotFVUKvToppho0QtmMIK43e7RCyRz+J7+q4U9V6y6KV8jNpXKDmAao3L
jNO6bRWz8JL5SxKWqFqsC7oyU9ilR4GIiXz6plyCw3CAVQ0ZmxNiv7QilG6mjr9a
eVNg0RKgkXVv8+aPrBGcmChykXlIGLHgTI2RbbwnvzeRuo9Js/CI+3eOkxlgcVdl
v2iZsl8WkHIE6TRLd8FR7QYf1/AHVO5El0xmSILhsO7rB3aCiM/Bw3QImwPuBNz2
mk0UrXxzCT6BGMfk0F+pvocaQB5guQODuc4aAdowltAlfv9XELiR5gD76PznwVUB
fkuebKUlnbS2C9FG/jI2zvCzo3pFpNryWkY8xMG68AJoOmYDPRidxfVjfdiF1+XP
msidZSLEd8QXi/Om3oIOj5vvyLBQheSzIMBHcTtAHpC/n6yGDEtPiAPd253/jZQV
r6yIEHgRdvMwmZSOg/CExYCmVI8pPyh8EfPmFPImBTQGW1SId5hjrx3btMD5r/Kf
SNqtMFH2+lrj254odXWBgKVxlSTzrXgUEV2XXGmibnAI5zODGTlBEVj2lUXUx0WD
bY1aPo+qUIKd15cFBYrIqdqyH4B2WH8nPmrRhhbTg9xsHh8ju0mj2hdUZj3/cF71
i2NGiKR2wMgbACVjF8kq6BgKo4przcRgyYk9bh3kGA02/ZP9hJQnqUfL8NvRL+Zf
oF+cWBBoP1lp9Rsqj16GtJDyvqvXlEszgx+h+hFOIsOuWZYvWRsGTG7ig/UevxlZ
vOtk/AfnjEytA9SbLjXW6MJct//wB5cplt7cwRvkWth3IaOZqw31KGKcFBhFAiQL
Y2MxWkay1P+1+fXKGOrOKWGQE88XDsAOtkfRf1EmYWsX7uxCU5eWkC77BQURGU45
JZWy9PGZbg1oVu9crvb5SDo4ZGYKbkfEjyU1+wZmQ8zvTLWVyL4zwtQcoQ/4TXVT
+fzFhv1/cAoyWPtI3DFP7FNT17zjaSSvRcqKFrPvwiSIXZmpLj8qDv4jCnzEyo9b
nkF3KMlV/Bu4mLoitZhkndGfWePh26tcymNcTf8Anhs/aKKmFeCT+KsnQD+Kjc1i
wUd/kBITcWpT+YEAcyChVi+f2O7fI+MkKhO8JmJXBnwBu2wzBOEbl3K1zmRYJiDA
m0QSljKTQlG2XBYs1pf+1K6j9DVvcN6SksXfvU/prTNsRXhKnyOHUMVFQkL8lErp
Q1M/bhtDILuT1vTv20m9/JNJKI2Q47mNZY9bHBxjaEuJLABpWF15ddmjJJVDPxcr
QyDgkyObKHp4/uNasKhIXUSeYPooyU6M7Xstqe905Ml02S08idu9bnQlmfOFi27J
qf+WMiulnd2xUhEuGY0j66MwZkSeUJ+KQtK5U911p4LVRLzYGLioz40CLSDMX3hZ
kPssJ1q/S775WfX31X4seQ1ZU1QzklCJbZuEqvACScIdq2xMVc0JtSspgDiBcoVr
N7bTAQPlFAGbLy+j/kZCXVLHYlB4gokmfp5SxHu+XTJdzETcPxAeI++tyb78Kzra
Mq4p9GZbmf2ELDgDbrOGT7OrhCfmHJiZ2mmvklgt9EpRLshBnxCDae+WZup3J4kZ
B1Q5DmLUUMPv0+heHYMWUITI5j7ZqLNd4X6sCiWpKyUQAwNAzIrCTtKyzkCt5sCf
uTvhhs2n88tZnfwtLonRRNR3QvDI1JS2elDrjIMOfs6nYjnJEPGQ4PZQw37EM91D
Eye75Uvhc0wOieyF41elO+8oq9G5QhZ792QwBWS63Oe2K+t74dPGbSy/GMEvsb58
J1yQmYn1IjR5paXZ8XuAea8Ab7Ec/o9YQluABxJHKNtYDC7U7bq48sROce5RHlgL
SeZHVWB9/nCvwnMLWKR08KOHqoAfxooPzYsBa/I5C8q0VP1YY2tvPJt1rwW8g0lP
5d/uLAazpihfyqXc/WrAdKhhJ6AOxvSmg1r4CMi5hotTikkxc8NIhqNU/0UjVCBQ
6IGcmAVNqaux9XSEibaBF8e0tj1puKUijtXzfBJW8p1tVR7trrnl1r5nA1MnuJeY
ld2SVnXaxG3RcQgH/JtNMf2IySBKOrH0+9J8CFExgWsrS2WrX2tz6JwHbxbtEyHa
VaHNoX6wiMUlCq+AkDSjBTWt5od/3AL0jWabTorrkDHv2Fs5bwwkk+c49YFTrhit
yaWOc9SeatwxkjZf2IZZQLItQXph62nvOFlYSpVNt8b/G333vmBmFUuuGjvW1RA0
jwI1iY6q0AwiwpfPIh18WKDkid8iWB9bo6xrykO9aNELSgOad9Ilolg1CNSYTtZq
2+FUNZapcqqKwV6/dCNxNVzHanV9Ny25Dl9VUbAmmN5aQGiay732e3M0UBq4+zGM
14fuhWAfBTfFyISL6m8n5n5RwsyQcFo7whBOjwsUMQWlKZU2GNCUMNw3fz0TaRcU
Uam0AslUJJKPl1oGVDFH00LylX13GfjbcJF5fZY9KjdzdfeOvrietmWkOMjiTQ5t
0zyXnfYyWYb8JgZAQo+sEdTAjkiY9G3cZUxBg6zQGIEKXx9T8+nAgGKL42z2ZRem
zJUnZQpijDkYdI3AwbPxW2HVRdvVTzXRfyaZyCfyWj8sm59D6+BEJeH2drfkYfBA
beXZlkMLrlyGTt+KTKaNcvHpWemv3egVaWD2qnOAvBDRGreRzkKp54k8YuX5zcfS
o5JKBJopReeFFIUGK+vj0vigUdW90xpHIeFFgMAWy9PueU3LsRVhuAbqCJ+p630G
KsbwHecQU7YvrkpevGsdS4IYuknaM4CpA2+blY4jMxZ+LJavWMQH6nfYyXzSISkQ
WjTxh2+1UBhevlssNFM9R5N2l5J6BrSQ3ioVF+gq3cdqT6OSpYExOcbung3jzkCP
CehtQMByBVWH5Z6QiFv43la8j8ux+MSiYUeom9KZdQxtFS7U9skL6mbjSt/97REb
hl61QPVHJUbnqH3ZGEHv8tCmqOgSzNMfv0tZsKMMWsxABdbf7ArbO2/QxDNWgiPS
JZaiM1nxhWQPjlq93CrkeY/A0xx7qRqcl84l0jear5Tk4j8AVnnt8YeBo1enDZln
B/A3/cvBRTxfGpuLcFlQFr6yUo42/jEzGVFQvx34aXHuLoHWHhgntl7CyNoJmlkv
YV63jYwZKxoDRVyrJFgvhjReYN2aRucZPiC8gzma9Bzv+6KfpHdZJ7Q6qi9L4w4a
eLF3Xp1ew0hwr5KeAnG0IdRbY2GNhEVKVzi3au80+EcczurdCLLeYG0bWrfuK303
SkdjqRhSXyydwcn1YG2NR60+pAzVCVIHFdeBmAnGf6tO2EQolmBcLLFkyZB/RUc4
BLtpN5QWOW8Yh5Lq81Cg17gRL0NP4e+yJYKiDNXqXeMgGuc0E24U6B5sTTBXcDCc
2urApoANwcl7EU8YW7frvXGiVQjp/z3ip2S6mFZsnrw5VPL7/39z2FDBEGg8gbuu
kxEy4W475EQzT7YLbTJauPPZf1H7/N8QvtwuAk1pNpVk3tZW3wfgkltg9zpTcjmh
kML5++2eU+GZssPG/zSZ24mOrt2/wg9gFrLGbG/mkr0rdrMoiANKwMGmyG8s5R2U
EkuP4W/9WVoiixA3wXYdL79zsDctCqoDeSJSgBBdfMmm+OXmtyZv2V1EmTu4MoBE
Ba1m3317xmBhLVNLyuOer68N1RYbtPfFSbqxx9yucqp2p8BX3CzJ7juuNk1AJyWy
ungUgmedfE5e0uMfKMIXE3e37g+IRdhk3G7pckHJhO0n0NRHsTfFAoB+jgqDYY2K
ygUzSUx+zsLVZxZ2By9kXILNNJfnN8WP+Mh6WlhpjhaOXwRzRs98Jo29N9nFTmJn
PVTW4d52UuQtBJYYj5tzMv/RDmDetn/Ab0fDKbCZ8btGrAJNasRuIrGrU5EiqaJb
omqxnbynAvy11gOBhMvbVvQn/w2r2rCiooNNNlgiJIFG/cRxleobDHgJu2+UWzTI
I4Itg8CP/Fz5RYkLRfm3tedRoLkKfLRjzeQSHi8j5sHzbOL/lfDQf5E15Uqiv9zt
mLVauknwI1hPE6gjn0OAtOQZgq9aK3gD2OCg5KTb5JYs3Ympd0YIGWWa5Y7ILMRB
c0hhQfj91uP560lx4fdo8uWdgMFBEm9cntNkpHFW5zHbJcXNcau9zaMnMOEmYidh
jonC90UhPRdGXbw3gvAUgMz2Dl5PZwunDV4Mav3PCOIINaDhxq5/psN9HU+BngI4
7ee7CvKbY+k7D6Cv0C1T49aPGsr/zLIdRpPhlNGbH53BB0WFsgqDwM9v6wvU1+Kw
WqYyfP2magQCAW8Md92XpNlpU13wG7hBzeVqrlZeKBmoaTAYPA/OH/hao8IBkMf4
eZbiqYglVea6sfX9pZH+SQr+3WorIaHcZqbF0qZvG5iSiWqhhzMN4H85snfIdm50
48I/ci3nH0PX9yCMU38WIyKtKofEf90ivB81rtsGllJET35TpYNG9WbAk9rI50g1
4s7/+Dflhil5V5CcFPUviJEbTVLuPMSMmWJ/kwRltOpGCs8UUGfLOKCrVCtyVUql
q1236M3be64+2rGgWqjQMoqyozPYSo/r8o1eRu4gDyQXsYG1o3dnpIU3+GfhQd1Q
+2leyJcLfA+I/JJ/OEnXRa3RBeG9TCEf1HqdX6FL1Zc28tbDIA3Xs1O7e8fPYCf2
LHkLWChFH+TxUm1A0XIkIM/gb8TLxWtWwacXZhx+CzKAGnGVrBozLP/Lp3tgugVK
39nIVtNjEOyxBFyjMxrF+TP32mEthkFEmQic5hE17D1uwT2TZboQ0putyLLR6it6
Hgj0T/dPSRc1WsqeAiSANE9wbcmhtzZ4fqekvfCxckKD9COX5aO++h0fqYt//DmW
Iih7pnVI6pfbH1juYsXhdsssDuJIA7vMWCp9Cc9iIg3RFd9P+18l15l7HgG2W3Vf
FDXbk++nrpPEyuiGKIqyVxWDi2vVd3Pjoaqbxmz8htQ4rZ0dqToHCCx3MQ5S1sxX
CioxJ5o4GZ7FEtW31JyWF8nPokE1Z7KuCarfpf9Mztm0moEYUMdEHulvXy+ixWqn
VVnKSQTa8NJvxVtm8gJBiKNAIetgXv/KC9vK2SIX193HvYYDH7FtFUvxmZlZjTVN
q+INrZrkQ0G+IywWs0VJwMATBlgbfOJJcDEcihLYtICrIRIGgsmDQ3rJNlWVTuGz
ObJ82MeHlLfWRGwogjP1ozfkz36GKhrz9v07jaVd5xMfLQWyB5c27UaAII32x1qd
veDvHBZiMFamh/U6CD7iOkdvqetD1qGau/vkQ0uVhtnukKvA5wiSnxZ8k/SlqesX
TCSXJvG9h/q5Kh3i3erdfeXax/ML9oL801PLob5waZ2fkLsywrPBMAeMv//oQYiW
UQPP++tp/YobwP+NPe0gbV8mOBh70oInZm5VC8CEuYLHauwUiP9fu7Ys9OAoNdtJ
nW8rqAjofv+onmSsRy6sR13sykHKL6DtBZhX5FzF9VK4VnSEQ8z/XrgpHiaEpzPH
g4aaZfUMFF6K221ystdIDG6HslmK1wSxsb9obVTHkV9rKHvvsjSsJtVLiWKeHl0y
iVv+QZqI/+33iaSQI0lVT43qtfKysGTk7Nscsi6z11JZQjH9JUwFsm+bSfZ7eCln
PRYJ6pcrcXfz3Vc3oVvcveLDXavkgy+Bt8X+P0Gn+tzRAphJ6BmeMExStk8+SVEX
uFc5dXP7tTB8WqnHS4uHt8cDrQjJMnTjMszOuWkwxYAbtdZ3UC1FEmUH1R6uU4b2
KFa0duf0j+yObuGhKgqjs5N+WFFQYfX1jJNLeDJELQJq+63Ax6nT5SKJ3CMev4j1
7SqtBoVtIOMGm2oNawaegEAtz8+GLboRTnYgwMRkqFM/GHFtapyVvWfMD3SQmI41
wihT4y8GMdsaZAB8uxEiHOFjQWdTRpD8BbBzT1YQjlLvt3MlYs9y9H6xDkfMY7wc
UF/vDBjHw4yHi714vBfxD9iAzatsO7YM4nHJQff8HQUjqYc4zeQWFd2Cxg74guiu
u+Dgsz/QhXsaS/yqrwFtOymuV2jKs2aRqtgQY9LFcDvNOSJi0fB/9fJ3lll2cA1T
TAQ0vDmx7GYyn3YybpB0X0SNEpjIeaq9h2snJld/HGq5tV6ji4Lop8ByQZRqHliD
gDg+zkV2PVIQvzPkYl89LjA/E8wBgOWHv2vjVliohOOl2+E0+OIuy66rUi5Dap+W
ttSr1W8KjkvBCWIoM+hYfnunXFHdMEORR50+tvrYkHS4v/akL7xF+0WkKn8Z5TYT
Gl6/NniE2XlFE6sid8O5OlhKxwi2ywfp65PJMGbcGsWF/SNJqOTE0yk8NZSbA/C1
BH/GF287cW6nqPtf4nh+A2e0hsSfsc/yKRHDs1LRMPWcUgaxDQgbmYoVWpXgmDig
XAx0FQDeic3qKnNJLN8+LW1Na9bSHpxg+qHHi3QbLt1TU2feDyM2LW/R3H+qpPLY
+zXvL5itHca+OB7F2Lcmu0pSUndXHtP7K4g9SfN8jPTRoK8mj3CCoiTFyU40ma/7
J23a9sHU6y3AJYqgrNzHRXAx/WHA5C5zM80a3WcdwbwgeppkHfSia1G4VRRDkSYn
tBq8tROl2gxDCn1z9ucsoEeDga/eF3HrAZarY34KQuIDFNg6pjUnVNM0dwmYYIjo
usCHvmeksneiUPcYU1kG6IaPWFJmHvSBc7RKcAXa3Iab+Pg7gkZeX7DvcW/J675v
4pWKmkgtZkL/xjrr50cR5DgHq2+6BdaUhGzvO1tNkBk1ImlYQ6rZu3b3cZm9eeGD
OZrqsyrBtZdVgTGdOgwhutd8lJ6XFYwndc7vnJDqQpRbyjRl96l9Wkt7N1DE7J3w
/WZebdqb/Uq2fQ6fCVqVlLr1PnFy0TMvXZqF5JeiS6G+zJ0KNN+QtEJoPH4ejTcn
e3M4EqtKl7hW0EOelTWIoR1To7EPbcz7Blttwu/Dj4XVyQR3V8e7Ser5QL99DBlD
td+efltknNCqDMQ+3EiEYT20Hi1r8eGJlninyDTNfYM4n0xOgHOSE+aBTaAp83In
/CpWdA5a517Ph8fvLuHNlEu+hY6wy5iKFOlPAw6hBkOLiYP1j7UVVuNkY5Kotk4d
8sk9hURyU6HKb8beWJeGrqHCc/qKAqDR9J+fF5RejrCO7KS+BFz9KFVeMs2djFOY
RoueRr2kh7dbU0qcw35QIB+TF12OJzwcD0eBMsxVbigtUzfFRtPGseJ9MqJQLiIL
BPLHSslFmqq9XkgSdCYsBJR3rTTy6p7e3pUpzcPQIybDuYaHM03SidMLzx11NGYV
w/GzQ1O3BZ6IrOJQBSnznvzVP6kJ2P4OFJmiP25nxIYHLtBUIhkgBP1WqJ6oZQrS
heayj+Vajuh+zM1cwxiP9a30GWQDAXxN6Hpm8319xuI6N3v/afRD2k78Xja32WV5
5jKHenw+hUv4w2/SIiZhyffTlZ9mWs/nInKUwimXIuVzmqmEXfCnEEbjlxy5U/pT
rpaoRWzioKc9nSgMB+yl9rYvMhFQtPNiJ9doyOutOYiQ4TpjroZbSTSfb8vUv3PK
MRWwjj3ZX2BHVMRwojNBCCVBzT1shcdRqv/EuQ+e/vPQ9E7KQ/7lCd0Swvx2SZTH
MMuh6z0tva1UDIBccTPMiXLzJOEid1WK/6CiVygC8l5y1s+8fTvr/TBYvZ3DZ/h9
hs5XtOjDbvMRzGTeNQUsIu4qYGnxL5/7nkBN5jzx3CJCjfnyF+4/ZnTSRWtRdMFV
G9F5IjMZQmZDuAD6gQY+ucK4XMX6D5G9EsNpnftd+qHGzFwsZE0VZDN3SkNkZWDW
qSrjSgaoFp4AT9HvEweaP9Pu74/juHXJufsRJ7sLmjzqwigtaMQrgSUnXuvECIQw
Lx27I1xpXIwp0eR5gsjcSPAXAjymJhoBoPcjGXLfzjlSPe/FICAW20SbIvpATreO
EZpoSChdfoczIzQgi8oIIhkCYms213oHJpfJcRHZHWJfQlpUIIVJbnOSFMmugY1i
X2uuqGOUOmySeR3WuhqP7vncFft/mVkydFCQVv8f5nFCJqSSndCSmdVCJJ8DDPjZ
7z3FC3bSCNeYJG8ziQ6GD6xQa5aYPtM72IzvQi3E1u40XaLXi0HJO42JEQ4sJVms
0nzoEC+pi6zJ7L2AIiBHIrKVCJhqIZSYBqBbRzSQGJaJ0fn/c5tAfS+Tg5kegqpx
D6nFQZSjzzm3FkEV2Riwv2NzNkGbOLhvb+TGJLw7rdDowCpjv96RjkQrq523lj+0
dipfsXHPTGtqHMyhj/IBJp/3fm7/twdJDFywXNUrFWg4NF/Gcwy7gjoG003DEp46
oVVnh+07oZVeXEJCqa6NVILYJQuGwf70Ad1uu1laG+jsNJnKw1ICsMFyRi3LeZBp
wOEF4IMsftjZHrJNRDinGyzg44UudIShHSuP4OF0y2HuEfQm+IQ/ssstk46ENSLP
MpNY6p7qa09jEvj0Bzg1AOOVJmfARjKXgNyQ33seMoWAYa3Re4JErDeMlN+7HjHL
86ZdknoRZtp0NndrTS8/QEQDY3jqfVG1xBWrffK3iKY71abWOBOnih/IlxX7bfw7
NNMggifmTWSPu8gHL6B+/P/3hom4vYK8Foc/QafP8NYMlppyz37+nGK34aHSGx/U
Xj/i9MKSc2f9PGcpB0tRgpCxDagi9jb2TbW3IKBSQwNYvbqmaWlht9aaEnof0Dfn
VjZ/5Edb0dFTyhrsZmteXnmXXJyAuvDRtyIY6v6k9RHVmP0Yl+lCK2OCHuwPUbM0
YXHiy2+vah9kdOr/K6Gyd7tRtz2Hu/xUWVDQO27k6iwmX03fYA7OFy5eg2tNBol/
MLEX+vQ02TB7f422MGoCqOFNIIcmVLaqMVmyTH5qep0mxw92w+fTs1inK8faliPW
I50EYl0m79zqt6HjH2SQemBrAvpxQgBqSBpqYQhGInJqlAE3AXPQk3P8PyUsS+nv
hkX+JfD44mtMhTmo3a+BsDwdyxuYmTtMmFyTXqYG6+L+n2/jSgwrcmznZD+cc/PK
hiwJUpSyGtpJDGjDhhlLsdfn/SdHejLPJqRy8yJ7cxa64oAafV1wDr13pSDcWc/y
OJQ4S9Kt+DZrvgBBUuangQaAqG8YRiCA+mOTzOxhPAdtBij8XeQEQn9nPfvjy5WC
6EFuld4mpUyJCCr7S7QKmwApcxbSFd2DeudjDbpqU15IKHd7COljY9ivuMnHid97
bFM/isrIvho6UsDqMLSiWRP92HLgAATolx2SndOJEj6hnHa7Wizr8QMDu2y2f140
4QXgZFxaS5fOEu/PDGyHYLt1NukInmkroaUIwA5IpWvEkft8HwRWxLaQkkpCnjBP
JNzzunQtwX304AQriv+2dxq1fq3PV4opSKIl3vpRCnvb+F5Z0yry+0Ecq4vC8HLC
x3xnrcAXiIyVEAxo1sR+jhC7o3FZaTSEAZLXPcEdX0KgESlVFg64lBJPnCQlGlBg
V7WECU1nezxyig3qBbMO2K+ktjOWU1jvGvzXbgTSIL+dfhZRc55+gKyeScJYRjI3
4y1Lixpdp9AkJqNzWzXwE9XUpqxyQVIZMo7mpe5APu5xH3t6i7Yxuh94HoYXCr3S
1MK+qK3QlUIj9i5k3VB9DwNR+SEHPwrgnNnqGrZH4o9tsGExiYgZG9pR37W+uWGV
juWVUN1qbvZ62cPsdsWY7vcsUpp43ECYZYG9cuPTNS7mP5vMZBbD17i0kFXjcJuz
HEqoaAYzycOvPh3QE51CtQJ6M8CB7dk4K/ssTVv0wTWzdc/Lf5iU62M5WKhlKKBU
nwimMZwUi1oZAX8pPXe+v6CQc6vvjCyYfKhxinYymfb5Zky/9HGFXCPWBqVPoYMw
F/WXmYryapA/Y3Q5sCwL4Qtj3b2qDUXi7c4+0F4E2ApmMcfwlAZ0lt6f34F+Ls64
Zphv4qQEKl1Q/nrrSSEmQg4aZa/K/mMhyyvk1JBa0jL4ZDplPl9mlduyKA5/EI8F
0UroJYw1Sef4/XwaK7hfdKVOEY6PC8uQVy4JhiHvv4oUuA0VYDtLQXqwJvXl7Iol
5jdnRVTbQB3hJed4CSs+PSNh5Eui0nIXM64dG0l8kJXK6E88YMH1xIRq3Pv0ja2P
r6ATyHhsvp1MMFIUj8bSd6Q+vJSg6W5d4D9qFPfvOu3Wi9dik414Ppcex4Qac2m1
n/581G2B1VseYvWIXnvR8+e3uquChCaqxxaStJ6dQPB/AsWPB8gR+WEQHfnhf1n6
80aQyEtB4XU//ufTtMBew25ttAUdvm/KxcIKgl4GZuXa5l70FWQJ4Ai+Y8el3jiv
XmvZTN7h8T2Ec3z2r3I33sb9iKLS4sfpB7HNHZcSLlTsriD4uLXsPkxKLYE+i9q9
4IV8bq7gFUYTILEZebrYd+svjgzbYvObf5OvREHSbdc1kd9xJ23SpDvM2FX6rxEF
1drACTAzQII7tu+xaIrQ2u7H7nbz63IaImYNIDSsQcuZpqua9OtP64S37WRGS/e8
dm3TmOR1QSPjYbYn1P744jeHF8nDPBRfXf435ZCUzgsMmEHJc0lBOxZ9WdjHcG+m
kencHzAhvCS8AhN9gQBCUiIlOGT7z0IzhRXD0e/Iw+Cbpv1s0hbiX7tWnUF514Xa
kDkfCyDFpXUXYututD6czRUPDxPHslCk4z07O7ov28Kaa4gVDi1JlaWU9In157J9
qjrwxI5cr20cZzK2RPta48kodQIbpPHAtK4582Eto63beECYFy6S5bGdxcG+Yjlq
X+DH6fYwp5MAeeqk+/lBzhUBSLKkHRVKTYzKNMKJQzwCENDXA0Lmwo6qQLI0qoYc
LTGMymPAwRdOCA54U/WFPGJJs00KPdyG0Tl+wr6ztQ2gz16E+o+1ps9swmIiItbx
YcsyWr9gkLr9unwSciOCnrk+Tkz3nIff/GZLLtUux+NIRu4fx8q3o+MreJCpFLuR
6xOJnBJEqGzVWmuLpPpPzNls0CGUiT6Rd7D5nx2vqzBcid5VhYDvE/bpI0osQtTK
+f5xi1Q8RkW1t3tPNQWKXrmrXhSDOfzWrFTGkaoHZyJlP4m0uhvYicwKsRYWOySD
MLVCFEtzNlbou5TRe9QNwtzc/yFxLxU3KY1ya7LgXQebaQfn542NZ6+9ZjFBbczJ
RaL45AdHh1KFZxQV+UVKTRL3iL0DlRzQ7uyI8tE29eyso8isQY3qWgas5MGXjQEK
qxSxhp3xnBwxNyik86QAKYdXeKlI2U6Qk61T1tJ5NTD3mj9zc+pDd1eCFMUNG1S5
qvEDGMxbM+13wdtMQVT6bmfdGa3Ygb5Ebg5jKblBkRcGcRQ0vluvLJfguoEq0EZ0
fL0B4mb6QwF4Xet7yKIOeb82MN3R6npmtFkCmxZKAj053PkkC/7XGobeBxoB3Wlx
53rl8us7hYAAU2SLOxuafHiuvydWeTPuoQekpyvjsFkOAR2lSg+b+Ra6Mg6TYDms
lkDcFXcySeOxEPTV2Mofo4TnOc6VPAVx91MFiQGNThnW5rGQW6EyJPNCsI4YKcZB
zDwzRtlfNQAyQk63sh5BA391UngRcIj+WBCe/oM7KDpS+NgrJQwvHAH8ZKmRdofP
/1ltdJ9fZURq4+3GXz7Sz2JYw1xkgYICePJiztNlxRlUVZpRd5ol0dwH8AREB5qn
2tK+9ZH0Uk0n21tPVkktkrWD7jz0GgO+e4IuT1bBqrcRgTKpXoA26yJwwSeKwd7Q
TkaSljs2WYllhwlHdhCyI5nS9JVDzYRNow6OsGcjAn/wInYksi/41ur80xiIcrne
4lZ2kfb4+rN89Ya9U/eZWVjRWqvNVL10USKrCMc7Br106eTe4gVOpgNsFH66Q9ZM
7Q0Natd8RnySgKdT5Hu/R6EqXwyJKr3cfvbRlhHY0GM7+SMiSX7GladdHVPD9SlV
mLskTQo9fb1zAjyUrAjHetf4vT9Z2HmM694zxroU9cOQTJ6+ytoXH8eqkpYTgAEG
RK9nI/ojottEtF55XkoPZTmCvfHRBte/dQZWugn6GvE9rQaPoww+CkNeCQhufvpH
YPuaQVf9fSmTT+xvw8WNOzma1XFb8Ck0oyXixA7vi7QfFS0h/Hml2Puoj/Ac36T9
Nzr3mfB6d5OfUH7vKjxoA274DqI1+8IF4910iAWxVCVfyowAb3yeJMW//k+gZXM2
pbrrd7saZ5U7xXH3FFyDz3+ihhn/MZVEgMITvA8k3M6gmAwUKuUV0Mv5G/VVu7kf
oCXe7gMXFct8owpO9yJanxFJ30VkOIMq+qBNdCiOO+Wf9KfoAwEup5O00cEpIFKg
/SR8u4WAIwcnke8hcYK1+dKU7Ui5fPchdeEAbLwyn+FBP+P/rFJ8id05VRf5evrR
JBNeVfyLRfvn+QalNGMFJLzw+I/zMkv7vpwhFrzobw558Y8RRvedGZnHNjfb+zBS
Tju3YdWP7w56K20K4/8bDvJ3ogDeKNfj+3PNRq1SOdrDLDBwCvEwMX8/nNEPENuD
hQp15f1/wryOZZ74dpjOeA3+Ziul+I7rEhjPFHEjBmTtXiV2xGPn4KG9/j3iIsZh
k7d18/SJk//JvMCwA07FZzQeXqIfJjLZk3nF9R2tS5QQh0eSjETg+7f5OrRebSnO
34olYjUDFERU4QojWSKnTup+vIrk/7TfwGMOja/cQnjzqh/Rvfzq4TbViWX2ZHmc
QUgakPTNTrx1zMC3e8/KzkVTjzIm8I48Q2HGJQIzNy6jOkfcnzoyGDeu/hCGmrdI
g+UyZtnsEbwiqiWY1daskxVS+LdJZAYUC65I109UzpfykLw6Wsvp2xEqJjZNwa5Q
ymhpdKv9B6yGLdmC0Pw+EGYindyQeWxDfMlO9OmOC9LZPGmMEb5O6pFHgnOpOJLf
4tJVHQ3++HJom0lEKOvYJPRzbP3wZlaoZhfKVPlXKkiiwv1i6E9/BJ+YH1m+a9Li
Wpd5h3YjzMcAFuwfVXqHwA/PsZY8By0yLvrbY1MWrW2R/jpZMBlc6zAbIIP8WX8M
Gb388V93NVNbBueRNILGjYHvHCLsBfQw/zNcFy9zNea01nSEo6Db9okfc4VtrbCr
hqhjrwUEaHZaVIsMikrJ5THmqOp/m4ONyITk4z+qnbA8BX1xY2Fg/6SohJTRnSIl
AXdjWu4OkvdM/bq9wF1Mxm7vds04UlY2NIwTLm9Ow0TGRbVfetGeYOBNp7PK6gM6
Ssu6A9Wl7UmnDHZwRoWgn9LghfNQRxPV2GytN9diZXLLvxAp0NSn1OP3WQxcP5K5
trpAoYvsg+Bj+idKzWmIfAei46JpJCgtY0tQckQoTMqUGvZQat40w+6RFoHVXG5y
wUebeSW91hNZkBfsWbauhPKaLr2VvJrKc4D/CIoHMaotZP+dqcOnzjFFiUEqffMl
q+V3WQHK8YkUedFTP9CqiPMOl95MdpGgKgqizozxRq9n0AQdcpFH4LoagD8QP6GB
JmEyy2LuY2e7MnrWMSyfwZtEyld/3wzHUgCB+HhraPhnuM4OXFUlcPVMvL/Je/5t
yB8GisPSUY2Ke4R7T1+AyI3EbOAnFYhLDMVBwdDQP4yLOHmLqzCRVXucmp2l9iNa
A2z7egHX4LUB/PUzJlNsyozIp+QG8LNUPDMxbn83YIZZe8trX07pp2GVmgRKtF+4
rpt0U5mV5VCJ+dBnQeZ4OsGodqlR4YZsM8KY0t79NQFuWQOaLg4WcIpP3o35D5Th
qfZp0q5PUCDgUI/SJy+Av0lSog/5fnRX2mGTjbwIvS5/rHXPWn8nJbxxj2DyLKEz
b87LO4x32kBZRYkV93u8ldHBsMhnSJ/Wjan5EsEynZrLhw85COHuMKq7vyjctt1F
TAgNAekEuMjnQs7TNTYY9aLls/LE23tedxnsFSJMiznV9myL5qs3dkL1xqUsb647
3ITwnbTR2Kyre+sG0P5EahQqsE1DB8zdaC7KmfXtg4NCHfczh9jGYO0YQxCCByux
Fe8s3zdrsyFuK8wmcrvb2acXheVM08BUHSN75GZzRkR3jhFeO7MHoCRvugIP3d8/
FXOT0RgmVch+mEWL21g+1TBfCFerDNQmMxTFGetlG3wtnX8HaAHC1kOWIuhq1jCD
BMVTJDGIOlHKS7lpuduP1kVi5lfnbyZfm33y+4ZL7loWi55a9yUd/6i6BslnRreP
js1BPVbb6D/zYuZYTUxlVHRSC8kWcQLzLYlm/vBvyVSO/p/jYPFemtnmDGqsa3Mc
OBT6mpTJqg1p5Qwu7URhtDMYIvLhi9SOv4t3ICFkKIvZAsanInT7ojHgI8EMhtaT
Mj4s/Bou0tR7QDGpi/OXRCtEY8rlm4Syy9GQyjaEsaiAzur3hdsyU70ORsNJltMm
bJFFOKeISZJqIeHkTDNaIzSv+1jbbt9PgkWl6np16avCJTq+I8ENVwNiGY6mxOHg
u0Br7bg7c3Kh2EyZM/jf0zUGchjFncTQr2/v9DoS4V73wbwWuvL+pP+9XpoaUgvm
ygddW9zKfdXzxYegIx4e5iEt9AL6wBIIn2rp180LqX326eNSauxsXicmVd5rDRPe
LeVeR/6i5XFggQYWVWibOPneJfMF64Jz8VWKGFG2t7mN9hX9C14eVGP83e4FBHrg
1O4XWtLulJLKAZR2kjmFBvbAu4TAdZiHnTwmz7SNu70gGmoKxev/Yp08RCYdt2Gy
N0mfN2VbV+Fnfx1YvgpO0ZhCnCZp6VxQKzZPSpC9cUQl0staue2rl/uN+tXLYHKR
dkYzjfrqC7vtfY4oTclhdTr1YA7IRTPIL6BNkjIzPbGWK67E7EasJDEb75KSTRTy
kb8HPh/+9qOKIACmsuzjZN3mGD35W4NjchgRQ6e9ii5B51tE9uFH/cgcFhYCnoio
uaDQWq7kBCBxCNjiMqaNIWQmLHDbh8SZ/GRpqzCNTeTAuWXVWvC/jGz+2z29z5Pl
3YerDG75iPGog/mp5+DxyM9fDIL+1WpcI9ofmhUZfDyohciVT9I50oYvf7ErtMZu
2Jj30UM2CbzQYFAKno1LW7sznLjKqgSpSy9aoQnGQFbMsZOAutaZdJ8BHKtg4nO9
T+6qk4pYKurAwBK3F2l5XUB92H45w9DYP095Cvq+rJcKBurmrhBVYd1/T3b7To99
ZaGtWY9z0YxnfPhqTgVSJIBEdPIl6lF9FzqmfEQGygHKPyjTRcNjmkfAgNVNDfjX
lnKUdmA3pHfNuR+czu3RG3jlVYkdC2Bi459aqQsambCUt38adiT/Rc+tuGY9FwGs
Ys2YCDNcQZC11PxwZXLG8KHwKpC2U8S7rTkCCOKoHqfU2ezD4JNWK6EAghI7fKEM
zI4Z/8HSMEfDiv2fkUH0Kn1CNruwdecZA8VWINWp/rGHldNjzfhT/+17i7wUZ+jR
k36xdvpov8Z54KQobZ1OWkXvzWvmHRH/DbT5IUaayGbRYBtsr9dis65EIL4vpYBW
g0oSFHz/pU3rQK25/Q0mEF1A3A92pTz5jUGeZSqAmhC6RKGmpcFiuYJK3LMpRIjt
iWeTX2ALdpB8bJbSwk+8NaRrAnlSYO3D1d001bAjr+GHXe0FiBeaDpXjjVdys/e+
XWYsjR2sFKMrPgq4cVzItGUIQCqAz1e7UPnHJSVtEnX/4TA2D5CLqE7yZv2AIB9M
qmvzNxwrmwto9OYZDEiuRF3pc1VzZaUzSLBKRUMiWp0LafhQ1qQ7R7FNNx45tHPV
n2P8oTt7C+JRid+r5YE1vtNjORcqC2APLnSDK2EvWhpsb12/jc4PcKpFx0QnE6DH
/nbjiv7lfQUSNpEBekVwpVEPuXdbct2qu3uLAcxeBwrXJlqNYVDtwpviaJVO2jcX
4MYKw3PoGSALviBmCxxvd2WiAVnYf6fxo6LI3ti/1HHayj3++IGytvZBuLSz/sCZ
Chv7KKYWjUviYE7pbjHjPfX1kIm53Uovv61yFJX25rboh19qG5TuUBq1D+IJWm0E
2ICYfx0M2ljqpsNN4nnOPrYk4Fhi1Xrqqa6jwP1/ZjxF2SD4+OV4kYU+9nXshXnA
O8WBC4Vyb39tTK4igKbWNhAYq/yWjho8ehava0Hcx18j10vG9OgmxbqLF8fDf1nL
/y8AXkmzZBmKqZ7TkjMHx0pAufJGRw6XzS3pXCZFnS2UVeUVcwyf/3NzxOzkg7/d
O2+4qW+dzZwvtHnNSE9z5Lng/frC+CMeNKg+gRUZz+SsJZ564i7ccifHf7g0erao
p7bGDefNsaGvih+WX0TOsZSwvyrwYT5frTQ2NO6anTv4ZgMGKi2L68EcLxnVHU+Z
Tbd/VpAu0QTQF65vJqIiA3C7VmHHCFjl+Iar+09hEVaoz63UXJzkurqpyYCys9ty
16wuTSAsX/eLIIjTdkNvsK8GiumpsUq3y72CPv0bsHf08+jqjq/M5kufcDWTD3m3
3U9/ABeAGRf7EENR0zKWrwURq7aNS86xJaWxbrh9Kl5mJuf+0pt6b2n1M0ML7bjs
/GNO8qO4GaeU9kZWjLYF54CoggOpPNf6TPGPaKSTrBezuKuLzBNAG7/eWos7uy3z
OB2uTJ30+7JAyWiNs0LQt9pDsiOTbHqhdZnPJxrgntWKJ0/YmusqpzlEuKZ+6kOe
/AoWLlDvvtXSYHQD9aSb3KqiuuPbtEXIvihoucEoFn5SWyLAr+W76zZ9+gLj4OGM
0UtgeAy+JMQa4cXLYgU8pmzv/nwIrJX5kWwX22DIB6JTvaUjIkUWHHcVInZ+ukJr
Mc66nqGtkJEOxRGf9NmtCO29DKruBAI/Hpw+qeZa0kuuTNRDpHBUIVsfQBYkMImg
mrlN3VpRxcVQnMmy4Ti08uTgVvX+HftQXKn4YC4Bhmn2G/AFIMXC1uYmTV8D6rNj
H8EGxSW7AkLzWQhUsoYaBNAkE7//irvTNFv3OSXzYwaxHlp76O9ctsnfm9B1XISz
DMIV5kVBtIgyDMt0q96FW6OE3s+H22MxvcqDMeZ+3GhGuxeLHGSlAv03mEdmpJFM
/+ffAMG/EeDZ3bx0F9EWov6SxXEFGyPRZXPSTvRJLQmBTsOJBCNYEotYsKaOFpMR
EA+sQQyrRfoAniw+btgE8fi7/ig5/iCG4YIV15sECqc3bwltyJlLYLR3dcTTkJXF
86BGBsIMZyEdeKE3ZbDBDCCeL8XMtPtyYjnaMbGJmbDRysKV/gD9Lt0ysoPz1FTD
/ojIf9fHvxJzeO+9wzhTRpu1heVIo68nomi/lF+LaPV71l4yaMrvazOgtiqDpFAy
+8dEpKmM4lqXdIifSahWiSKbszp38+ISun1P5BTz7RnIqAr8ZRZ90FMR0/G7QCOW
YvwzL3ILhKrTyrtUW6IgvGqlOEvS3G+H2rWT/ZTDM9N4IUZRUZiUlreiid8XvO7O
qdpmD3ffeL7f/bVkhYXdj89WMRXB4xskFepzmYSIMksJnyZ/rm2z7jLfnduYDmmz
6TV8hr4Ok9bmWGPTLAvH0xaNzsQnCKPH4xcGOdN873Zg+fGLjP32ueVlMYG1W/FZ
DSUAKIyr1rm5PlDZ5S+uYTPazrMSZAM9xvTEBGz9rfiGTbnBfNz7zjaZ/pbKem5U
W8AUCqUcFJJESbAW2rIJMxUczogiAUe1Q4Ki5aHMsscH8fA9sH8SJJ/fwaMNr6jY
mPNZIZ7AhZfPHy0xBiHhNB9kfzP/gjRm4lVbe/QkfoQ/BL+WxO+kvWXLpQlCEEsF
B+2spXFP5f5tWu9SogzTJqABp//UENrbu3J4CBku+xdguhvh9FytFmhlkBeKUoUK
g86cJiNFpVTSCrRM2lH2O8D7QwLgcBMSe7vHkmUOJvR2qCPfXTzZVdYJGfl484vb
KWi5hNGJr2iYe5ZCmc7mfyB6XsQ/FL/dH1A/eoocQrhMlTYIPRp2tApAZIjX2nX7
la3+0egWJ00TsQiQk5YWtZ9ThKOYMJ8SYtYZ7OnCeXDBNH282uOXUlnkGZEvxwUK
dQRLO4B7NMSl2T+LDcAFFPinsC67/FfVpmJqUlgHfP5IR4KYKfaWraSyalt5/k/R
WmejczXDmz2LDrzvO+mQz/XnzS2jNWe0ZvsTB1B/lhL4Cxk4drzDcbIv0slLABiq
k824EzQYnIqTWOKFZYop0ZpcFxhpK7X5Y/nDXGG8Qll2M5EGnTnIyFN6e5Q/K67d
IlWT5s2mMsyqJXl4HHDCpy38V+mxU2XHJj+oJr/Qj/zkL6ss3pQfNDBfA3GEoVGV
ssVCQ9QOZK1hDpweyvTO9c1JuOOS4XlmIu6AnVDjK50aibKicCikI52O8T1aNJqz
J7V+PgtCHjtffxxi1Y242wRTLO6xuiB6CvBFFEGsm9FOk8nJE+ocakiYeDA8YyIm
lGDLy0YXdcpSRkZupFzpQ7XBqMXgkwl4JogdeqatdWmwdDDLLUozyZNbUyKDVmjn
YlhSRBSnY/anV8vcNsBBNjoTtBAQ4PLRcGXLI5ZygpumVuhMoqX3L5d3PQU9lC0y
ggpKSCpQ43GxxoPLh+appu0Ok82+FuW11I+Ieh2RSCccK+6WhxWFYTIk0iwUjG9N
58W/cnsgezDPDw2q8O2kLCGrIRkwstE+DVZ6plVVbFxB1L17P6+gELZ/a9XFw+Y+
uDdamPcjDDpDQ2IS/IJ/tkpKvkQF8hb6/0ChFzQGA/yhk9h9as/Cn2N9RjMd7ryf
H3kJneTY+v5W5LK813hmAuihmsm7kuizJd6iq9Xel3gpRPPTKVdbCBSd9HDltM2o
audTgGURRWgK65v3VafPqN28PzMT1z9qlk41yRQ0+SWCkXYcSGAqknlEalshQCiN
/yCkJwHwN4ysj8ecU0p7VxXJEqB2A+xIs4AU51ox+rXile8017JxP4YynMY+8rUx
ZczHByVa6YEqX32rNGB96TIl3SRDQA6SojKChox7RHs/wDIzA1LBdP5F4TSoBVa3
ovPbiq729pUVJ3dlB8t+4lpQTdxCa4qBzCQwU/WeUKzMh4zEduUC0+eycW15V3gz
Uohpan+muTRe6IhI9lH1W5FhShzr7tOvmxXNX+PJnL4fIHJw/MWRWQIYAbV/f6p2
KFucBJaKAluy33MWbfxAxL6OzY2448UUXpF+MiCNpMyAHyQTPkfMLcBj2o/VVSNc
By44wH6WVnFwqF39vvWfsujrhZGV4CxKSkBJMsuUiooRxHCoPTJR9hJlv2vpZN/7
tsc443NAjjeUHLlDsWX3kAWZzrCxIL4Lsr+E567ser04TEUVKMr/HcPvdYBfSS+f
U0QjSOusWxHPsJYEfL5Ij9dezyWAEJFVSTpm2lQMiF1dzs0AurNdncJlmfYoECr9
BWJyi/rjl1GSphqzQMerKlPjbtMr6Ih1Y19eIZJ2CPUbbWA8crYnwKN5Zq1E9kKm
07tLkZrAPBKpWIoakiU+1NXVigjc4t/zdQ5pRxDWtLr9+B95bglptFA2j3OS5TDm
mEfbjltPpNGV4Zg2rnLqHqZYO9ilUwvjv77KmT0836hY4wtBY22HKunZWQ70+sWg
Mv0taZ6yJ4BeRionHqLxSMAO4bZ956WEzhIj1QuQBUYfG9eV8l3x05FbaHtoNBei
r/Sv0F1gaPdf0cmCvxcy9LVjP3wLN6EQKKEUSG5Oas5IvBbZ/tqxG4oroDReUVVJ
yl1oiuRKsGHG3IWHvmOHRRVBGwpkY8b2SuaIUyP4k2lyrACAlmNg09Cix7pbvlbZ
fWymQdj/byCp+Fyh5QG1lNRGbVYRd2kOJ0Cvmgo3YYzZuD2TTb1gyyru8Giiz6at
nZa5ZrPRnxdyXUSV0HvbFNMnO3pc5BNjEGpAXmsI11rT4w6a/VtLEJO9z4KdfVBh
3O/j0hfizYS9GMw36wvYFEghtk4qeXaacaijAdAIGXjGaHWxtkvBwQf480F8w57+
wCuJ5hFwgzxE1bCPBzmMxWvM4sVBtVTeWJU8U3q3Xs6VFhpouzrEfLhVd5pyUyMT
CQxQwtHd6CEt4CUto6JP8ahfYjiEZqp5IbWPmODwDD+DMOT8eVZfPXsNlpYFD6/c
MQfjXGbqVTHbJ/nRHvW8xbByIv0K3bwnrRNWxevAh/RJp7q2iqAKWX8yeeYAuUq+
8OPjzZCR2/+pF38PUcral+hNN9gdlKi4l6P2dmMaGfmUKhdU+bThmfPnreSzIZHS
5sAdHh3H8r3A/dAmjMTDyLckVtPNQghsb8RilthQEMRrNZmDSwH0ZFWtBGDhd/7E
91BHzSEstDWakJ8hPtj+MCM7sULWuwbjl8rbWkOfSc9p+ZvZANvl0i37tf/IMKF9
te/lYrYh4muCCvMK+vi4Pd3FDFN2mhInmDTv8KAZ0+F3HyEEtjKbgWJovMHYVuWR
VpLsIPk3HLpVTOo28SwIXsF+xXjnQEUGG2Q7fYd6tF0QntI7Wk6LHit4qbjFgq8x
KxjHFOydlWFAIrBraHgot8NCKaxD0Pu6HRSpTMarN8LkqQAv3GNdv3SOEnlMxhkm
7gglzOqst/gRPxiOP9joyndoVCONhDrpXd8s2Yr+Pja5TiD26D0dvU1glEaGWgaX
PbS2vzIcmGpuQRhTHZrKIctv4IQKdKc5425yjypIjQAWwFKZL/nRDdHgk6HKX0i1
m/coNrnD4lWGrrfR1QwREAJx5RrlCOzbcops7+FltgCYAjYWGZY+yBNuZtTYlVOh
zYp+C9bNV/T4rFgJsBI6V5ZmyxktuvSrzyZfjIYYugcFac9bzhfpwH7PDta4Nhjp
Gv3NG7AplDnJHUDSWdwkDvsuYaCFR5PZ2sQAV50Vi6EiB8uhw7Nmic6DYxzhmC5s
8at9BnN2NCN+ao8/ijPtbHm6nhj+GHyrCz5v8s+8+hH99k++rjRTSCyuROT7KUCf
uL4jO2P4TJzpgP6k/UKQ2zf5dbFScWO7sjg8i3iuRmAEIglRNWOnnLRuzjju/1pK
tXMpsZqs0KgtTajwYgv6mKtwsGvDkL16NRA8fNHhcss79PA43NRJ60tDNETNTheC
EvUUlAM2xGERngGNX/O0yEDZItVjYoVD0rKE7lZ9+8i08z6Q1OoecHUEHBPw14PK
07hDH3vgOEo84Yi7ecU6s3qn2SggkiKXvsFvLEKiy/mlTI64fz1S3hSIEzcnMxS3
rv3RlWCdEZgNF0D2xTOLOY1w0bMyd20RPS82VkV9yoB2Xkianx+DlAoq4DUOROOE
dmaFgzN10p+p5l0aqK4HwosvM6aJxTRiCknm1kiIscQGLUq2vW1XwJkhVP3AbWPu
D6qIt8EsPSTQKiQGXMhONANYpkwWHuETiygAsoKCIBlrEl1qtBDUveXJthdaLf+M
JRQKuC5gi76/coCShbYdFei3QxjhpirEgKGWrUOUIG9wDxW4QxFxfberD4sqsvRQ
+nSiN3aAN/13addDX4kAD9rgWn0f3IHB8KHK1rNzSvQgWxoW0F5/teXsxqurFu4U
S9vG1wOlMwTZizSRWW4+R0sDkj6OtaKPzwa0SWjSlxWDewOMMAQp3IvK6rAMLCEz
2k57QtIMbvxHPi42wy3bPU9efboegGGutdIkXyHk98TbsT6PlBxaDlrHG+/disWg
Wpn32AS4LwpwVPhHzvY8kadR1ruFy4XJMoliGzlR0d2LwNgrsv05N5Zc+rD8iKOA
A4RKOv/+Ao/n/uP8lQO1lpbvoB4EgI+4wboP5txt5aYrrLzWx776mh1m+4OqH5qn
Oo6quQ+h9CHKJLHAFG+FpM+l/4m0JZNE+0RR99UPWsUh0o9vT7dEzuFON0CdMhbu
cjhdC1UU5a4nBbCPIDw5HX4OyCh7BhKdCQrVSvXm/DRI5c2nXdcrjhIQ2zULpEEs
snLiGAmVzXrcyt3alz0wJeaBxhY3OS4CTkgAAqrXPqOzestV76iQgKw90LVn3bkM
FxaeZcxzFEfly9F3UzDH0B5Yx98wZopGKhQqK3Xd9fuV3g4yC+0znEw0Y8Yx1VKN
ox9Uibwmm5Bd8UPb6uoFfayOAgKhfI9s6c34T6dudWwmTGbCz8OTN8gE3GG8ffuq
cikZBdJ1CY0vbKMF26kTUwMCKLIW/UeyxMcgE5yMJwQXVH6N4CEPPRu+JvHlaG1Y
mOhI3aD9A78JmByLtuCCWbHX5tvJxnvuVtquM6QI70SHtzJV8Ng5C8cYfyFLSAW2
4D8/V72Ii7wbPyr79zK1TBQEnKvEVskZPQptDUNniic5fWCuyCVGGfqJNIt38+r3
29PkLXD6q9W1B2g6n9C87W2OQSQ+5yFxqfSy6GkKYX2u3z5hf0PK/+0jn5wKwGw4
eIZ3FNyqA76rn92bWPuufqdyqLwhCf7A5Kv3OOk6zCrt4H4ChVnZSD6LpKIOJkXh
T9d0SSz//D+GKLpVvylm5CJlaYpi+jK0psD+WE4dspKzOwx0ad4+BanKZU5v+v5i
B142twv7J/BJkNbl1LUqahAtxqcg6NAK2sAKT+/BPKOL/p/mmfjyY+Bdl8XDCJ2s
+HrXGV1QSeOEoCbsrXgMcShvzxpX3tkCNaEXM853WebrkpNplu1ctDMNyN6UeUOJ
8QbKO2qiHYlltUMDmiJDOy2MsWW3jS0ATgPoEzp78lZmrOZhocgBAiyw0227oyBY
DC+YNbLKv1+NmZvoQpn+eXcQBd32nEFe1HZnUyM5/cYsOcN+8htfFdQTsFiEWnwN
APdtdWjYO2k3IzWG/Q2cJe+VpOlshzKySUIr3mwNDNqlLXKPb0V898gNSKxMbX+T
LqWpI8QnAbgSrizqfxBfnRAhnYwQs8ecxSC6Uve6639dPtF0SvjRNFErAG+wW1Lx
y5GgjaObiqFNEJnEYkWvYh/Xvgm3gMGIiQRkoMzJlUJWyOX5xZwnc/1SOw1Uz+fg
HNAFuzRZjMOkvY2yWiVlLEJbXMSZzLtzzQ7wlt7MZzN0eH/6w8S0hVpA2XakE5v3
tFi/BCIwicqinwVPD8Pnur8KONA6pJjqwBVE2/kDBpAw/xGKXVuxA29AGfyjK4QU
fcJRooIrR0y58H0dlrFpZVthylwhFG0224G4C6apCP8Cfs7ERXqleZxzFK9Mfuq+
rdVHn8ZQRjyRnTzY9Wamjv5Ukr+xl+bucrdi6HjlEdsOI7VnFL/lzdDdiSCSSOxE
ScHsyXrgjyIP6yGTDqSjwKAlbNmzfIQrmxgqPRkF3vhmsq5G15wIzpLnmTFTaCqw
0dSXmQqcRXYPGzZwIH50rQ==
`protect end_protected