`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2096 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
XDmUU01KuyTGZ0KfD/yCUyVbZF2+vZziyxzrJzdkZN1oYbu1vqDjhWF1+69ekpgc
Fs/22vVrniajSrpqSiLtfNKC6Vj+bdhCQsc5iq8ifBLJpEvNmMuR/Pt8U92eJ4vH
IIr9FxVIEN3QC7C3hQFo5B2ziNq6Q2cimZuN8QWXurS/pAgwEtUAyqTz+qgOo/zr
kjs5Etdk47eZ0yA7YCj8cMt6wEv9HZtQSSBQn5+iizlAX1Ykw1ycMLL75zOqFLa9
jTUJElmWCoX575I+UzAfhDitxSlCtbRg20cbUDiqfO/D2pIRIgKCvEXUCm3295Mn
ynpav9VVjuZgjpqkKFxXjCipMO+5kGlpwNlC1+sw5AuQJdFADr369DyJsEYvrEs2
kdpRbR06DWsnistYVsMOOk9pofsLcGFP76UYLzYL2bvk0J754a1qF8j/7PnV0Au5
spnAakYsMa0k7C8Dexxq8JI7ZI3/dPB9hzTTLqICjww82pGtgfWZVmpEoDpYqoqI
NnLs07IprDdd/G5hS/Oz5Us4XRAUgMllLwck8yasFLe9xClzdp59wXygVz59o3YI
bJLFUXI2qa2XZEA6Tufzxlkby/I20cqcy1uoQDmNXltUxSFkaQ5QKoACiUqfi8St
ZsI3LXMwycqz8d//WuoqDSbDuvs3tq8HzR6vyX5cvIhwWTtW17E2wucgUDjvTuI8
5Sq95PbWLHEryshWj6m3isb+jLRO+CYKQJg5ilgXt3Tl1zV9h65vOjmkWxyKYIN7
6N1hZDpmA9tTbb8CAsFgLh+ZlaAOlOeFogML+zGD+KUl+4Nx3tHCDvlxOF1sB2yN
6U6/UCXItWll7QFGMLpyUaiuTUenLzfNUvZebMreDVAuLKR/lwkRtCIwv7yRuJ0R
YzjQ9ETvk3AjofGMI/t/U/IP1mxLvSXjg08ck5fyehLFINoxOQPQg+z7Ww8nJ07i
iX7rMpnxwic8VUzrxl+n1l72q06S+xli5m+jcDcIO+0ABtH2Nu/rcjqN+IhkdGpp
r2Dtx1/pftJgYDwvylCdEBMG7gm+v1BeRkNIFR98LdozL42pxFbU70KfITilYT+x
ynq1MnP77NH6tmwaSM7ZQpL0nTizjCZO+4MX9p9ZlRjr2D0BvY8tap4FGr96rDyx
sE6vyjUVr8FR3zqd9rRfx6BRCIbgI5XlohFhESg/hxzdJh/tYW/q58FHOOcCJQWI
DUhl9t8iwGcIvnhVuTfMtDE0gzZLqeZDAQTNuJA1fdXVa/BlZ0i3Mw4swIKL1TNs
IOVZKSGyxfAJbrAglq+52UQWyC1RsdiHcWZkHDqgEhecRFMrathB4YjGhLhNHiUR
LAWNbeOKBiR6Rh4WhUjSsqFtOxNdO1w1PJNnrHRbH+LfNdgaHjE4y4WiFzS59VbA
r6JCwBGUpPV3osnvomdWZTDLztDYspOxX2JEt1HWon+7m4ulb61nu67xFE88tovK
IoWH/2AxwgHynUylxq5GWLjoCn8rczbm+22oJs6yRzew/jkgGmXfJc+V6YUjKEX3
7VhhWyw1wW4fd0UXclLSgJHvqIXoGlC999Hf5+SzxaKLLzg3Q8v2XchPY3SIyKHu
d+v9EChNmMAJw+5zmkAEJKb+4M0SHk4oNGvA72NPo1Dtgaq6d2BkogDaUdTwv+bJ
8wqUoQCIeV5USZHrfJa3m3DZG+bqTjrNwMDhZTuEJk+b1tfdq8dmUJZWYp5F23XG
1oili7yTK0hlZ8rkCGGlDUrm36JkmYZdW9FfS4NOjoWtaAHZv6yf5M/UaGBJqu62
5TBGJxNUTmwWQM0Wb30g/M68mGH4SIP4zMTpETF++/m1YdJ4uv5g6s+FsazJbbdn
YBVnnyTtaGcEgDamxXo5E1MpQ7aMx62wAr/BFfN8QGa9lXC/iyjLf9aFZn4SNRJC
LCTjf2JVx1et4X0wObXfr62R7YKcCmOrKRd3fQGBcPPmoRopZiT9D5iBOdaqV2an
z0qCTUzrOhaDgUHJ2F6zCNSK08CR87UCBLptsNThGXf19OmRsv5Yy9e1Jz6zGihx
+FERmi5jPsr+5T3jpy8dKH6zbAnzNRn1yf56LEc4gaMPSC1KRymXmxvGaBQPURYy
0RIGyQxV142kjaiJlb02WcBOA+gGr3H4p3RWtiicpF/2ZQtaBbk06YZ6O8x8eQXT
giDXPv1Oo2DCh6NDS/12/AzHmcQ/ZwBcc1s8I/w++d25JgP6CTRPoRryCky6Uj46
ka7SJLm+fZTUqseE2GVi3pmEdmTtQDDLsIBrih4GmMAI8Mf8ccaZlph8Zzy1NfE2
3BmDsVQZdVqubEPJy2KTD6ONBVMDtMxMRgNe6h13ekholWvlEu6b+dWjMpjV1qvu
ubo8vNoAv7mdIaW52kNB2IsuUYstQ68FdwkEf638VAXRy6a1HJ+RfWF+FslTjH98
BE74MyyBI0GZzwlo4HE9ewXpETVgRe7fN9yvwuSjduTpy0Y+oGhFVe68aQ09/YYi
H30KWWQ01XVCxMs5FBN2nbmdmInfvHnAS4hn2Y19oQ9uNMG4X2YUoYrmARfl61h1
3VsfuTEA8jNS6UhODSHwQNqEpAH3S/QtceOa2epZisy8K9JXbWHWnBwGOrKLKDvz
3K7tfSPxdJpk/Ph2Ll/yLAkARutgdGQ6+wMgAJXSvu4=
`protect end_protected