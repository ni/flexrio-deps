`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
YATj3kULTF7Ty4ORuRfFpnT6YIk4rUPRrM74bVTnc4GjdV8oSnW5PtQkMCLOi558
1V+/wvDfc3y0Z8//ksX8sZm3JZWtrxUppw8c14g9Y7owiwp+JumRtO1zuk5xFbe3
0MMnIxxoTKLhyRJtAxElG8sbx8N21OWDGiOk0Xyd5CqAmk9dcOIbxzMjW/wndBXi
maijUdqS+5KiRCM9+Gsp6k/iEAa2LnYTt4WtjkmDD1P5jZKsiMgFck8WOqLymplZ
ml3TTfn1UlLNm/+zD3SFGP0kABAiUT8NK2xBPQ5UzQ6sMFPd/np8iUZ5u4QLTWOZ
hTrU9OSX7lOvRUo8pJ9vPg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="BzW6NOo8eyBw+CxsNNo4wIDxODIsVe0ft0K5tGuSUZw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
DhjJh9S2BY18dG77XPz3hsiSQ73+w0XqfJhD+f+lIDHHVjOB7CfC8ieNRTexgzn1
5W+qoqOEwenoVQtit9u3XViXJSRJ0wfUC5a9axblRNyD2mUbyfH9+f59nWqGkVOh
ieHxkA/DPprM70F3APxk51m7/gNSLICSvbONgLGndWc=
`protect rights_digest_method = "sha256"
`protect end_toolblock="L7NTNW/5Dqy+2kJZXKczEa3js87UJ8H00YWI+92sDHA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 61520 )
`protect data_block
6eHODtGLmq6ccbB074dgNWpdzW45i5jL0Nzx5wwM+RA0eeOHXxEV143NNyQGmZjT
bzHAi/6AyRCB4X9z0c4MjyrZE8GF4crbMH4T59xFHqVrQ4zXCea5w0kG5yvHgpKo
rwIIbW7Xn0p+GsC0S8TZElSDgaJgFE8KNc9RSw8/29bzvpe9Nh3CbY2WyYxW03GF
sMHAgPvjhCxXQFste/yfZdW82Ny9e6q9jj9hGIOXhaEJbJVKxJuKAQ6m64ttNGKI
ZCMF//kWl8w5d+LQYvvRplp85ek0L4o8TvZV8oi8BZdx2GOsImFUr8YplDKoh39F
tQn9cNSzKHL3l43jYkuWk8IMIRepun9N51E/kTPKTlz5YXSMILmHE2LeZV2YIHo+
4aO54Bal52wqpY7T6N+EGjljmt4OLUYrhRHEQ6qSIZHG/M5kyJqO7F0q2hhYEL5b
61CPRm92sZpb3sVGJDactPPp7Yqtg6Gld2Nl9eMQUZ9WYJGsOkfdfjs974XF1lJb
vunVsF8nwamLv21l6lNuPjRo0XTStua6u2FTM7I8B6PQHclaaMJ1em91+33ImJL5
QNJeOQRJzhcmyTrR008ofZB1Lih1FiU6U3KePC9rZosMiF/KZxIQ9uYbWoVCXBeE
UAN7O2c5a/MEcUbLa5lS/RXcXtI+zsoNRG6fjAz6fsFuYrgyAvLv96Zb+aKJZrT7
RvTZlxoUNCdv5l1PXJseudlIWjru0vJph9pDphmIcXvyQfsQstrFfpNamEVi5OAC
HJZF6LShfkZDK24Fr/WZP9K9EhHSMKxeKwz6Q0KBMXeOjvuBVdAf/3dxkTmywFQi
WXjwPs37I51/srLx36KmbrW9FhsEC5tE23dFPZoBQ+uzKbkZRUWALguUkXlOYRdq
xpVQtqw5v0wqtUJrFnPXpzlx71c07tgh2D0skzM/XnlqyKr+2mNNvrsSYDJXCZuP
QehPKSbJTt2XVNuoKT6eBV51XJjrI95S9SR0zWImjVQRcX6DzuEyOiLFZlNjDuzs
n3JcGPUX/Dq9HjbDEISq3aOTAN3NQGiFs6mx5Qy2Xyfuh+PlXR87wTQDAoh83aZb
pKEYDaJDdNntUiknTvff3cMjS0+5idSzp40wb0HsXm8aP7Z4FqOb+5kLhqsESiRK
zKIrQ4s1b/LT0xMClDcNcwL474OImlYhh4vh2lGNfSjgukYb0jyA/OYliAOvE8zz
tjfjBmZUrx+1hpWSIu1GtbcGLKcdAdBz4BA+ZEXi4JWoqseWjXQVEtZNFuLcmZLD
CqNF36tOkcFDlGHg9s4Zb3Udeg1NjD/0zt6D3S7UR/bzgPdmbJq2B+MyBRU2l5e5
Oxcx9jeAVXTshgQErKp3Zbo8L+OaSbxFLFFofvwG06wY+3CbVoF5lgVIJ4hoGwnC
F2+EmHAOvLmCZz5e2qoEjbLT/xdbGHcp/eHWhDE+2mx2ZV6Is55xPvhX/SeeohUM
5i1KwyV5g+JYuPIlqO4sI/zQiW9RajaqixAY5PDJa0cyDjXmSeKBKTGiSn6YIuRo
2ISSZK241U0XVvyFbcX+XdY+9ISz0KL7n6ff71Cpm2GrSTIn/Q2+CsoaRBechcF+
sTEYNtqIRPFr6yjIHITiLtQD/koTrqcFaWhqZOY/75HqQMabiLypBBw9Ft3j1H6H
oOcdkV9c7c8TeSRBLDAFDzmm8zj2+aG5GVpeMQtWkt/MI1zleiaXj9zmwBpTldZ6
I66DdCqesHa8wyC3/nfMEy9MH30xyTk7tW8ESmvcBHkyOEgyWzmtHPjHXsB+/v0x
m5KW7ZmUirHbhqHyxGg3sClyvxKGstG+UqZANkp7KzCEir6U+A7ZaLs+HTOiZ09M
2K8GxHaB/9eGYVyX6JDGadLVfGyLGrHdpkPQADWnDOEmysRMcsgbAKGyZ8iU0Xd7
d4BjGlDpTb0U5qLOPkgevXn0Na+5Sq2q0jkrGeDifw/c8vU1Fo2d4EY+Lg7KXTzj
gprpOxRWGXvdyQqp9/aiaXcrmCKfRAlq3U2TEM1K7PNgIyzjuz/r6Sy/iA7Cihaf
D3Q359m3a9Yv2vFhoLFkNYsaYRCAs5dHx7RCc4Rq0j7LeJb9tZTH2ODJfSwbGq7H
sPpSNHiJREhyMqOnr9ChuryqycQdsoLqORtSunB6oJFk5FdYg6IabmCZ7O6EGdQT
dWitO7w5hIysbtYMg1ru/TAo2YVMy210tkVoybwFru5xGBxUdgE+zKubhAR8HRd0
1DL8CnjEXAediGINMb2OOojtzDNIrAdlxo4s7ezxT9E9lNepHEYoKbkTHZRjVVxg
BlRKpop+CqlI++h6GL/iPlapOQv9IJ0ZegLdua3NgkT3oVK9Fm2LkosW7lHxd2zx
ESeUV0wjL8xzT2N7515wsf3id6PiNesrYDT45srJ6cPWmOAyUwQFA01gDG53D5wH
L6GYEsNk5bxbn0FqVkFa9iYWN7E/o/NEXKKMNqawRmOVKhJDLxGflkoKMHh17pH6
ILKsIewT2eQkHUW8bZRM+ZlkMgdyIt7fpgTZzZafP8JdcTUSaMc+HPsLWtoRb9Te
1/Um71PktGNkTxWJcFTrBvpV7HnhFrts/ra13dDX5hmebdpaosS8H6w5ZRcCuDdb
DxiSKIxGr/2zHcBMsAXPJNDdaNuxKYe/sfcXvpeJAbSpzcsPwsp5VrV5dwGhMNL6
aA7DeAG8/JxcBbFbJSg+QfKFjfWO48SbykQMrbJfxFQ8y3wsV7I1PMGWVxCUGYcU
jZdq9vwHYhBi75w/0shhwfywzW9OH2JB8TjXGYAbaXc8ZbJCRde+5j9LxWdLBM6T
vNTGTX7AeQl9+EucC4z7GGu9rgYXu8US7NJ4JnjLx/k8yWuVWgMrgwILuXShvFCm
lFnWB8ionlZHzHCnxqlyWS1U1GnVXmdf2EP8+DMYcUrVUoki2NxoAj7tgimSXWdh
Yu4Gc2U7gRIjNbU2WgBKS7WH3dTp2sBoE6sxh8pU/zmVjzJRu6owft9oNVhjI6Tm
nbBuoaG6V2Zrqy/QgpMJMqIL109U+HyU5x0OwpWlKUCx7qZlX8fY1XXhDf/EGOS0
FYq2g7/8GziQIAYvbWQYNV8p5tZoehNIZE7xG5JX/I3bdI0jn1rPPwJNWh2bXxMP
+OvdWlaDWr9zayEjsZ7dLhCzw8YkR1ekSP33hGWYdEnLsbyNWQgQEPUxdBBOU2ct
bFTNz5iGeYA0n8ySC4eWiK1pwRN5B7cDurHKEe/qT3VqUomqLamykjjXqHN+IJAz
DbUipFpzLHknugB7UlP5uBMaLrxBPV+jCTEhohYwhaeqJ6tsBih2fh8YrPRvgAK2
AX9x3nEcu3zp2GnEeP5BtJqlCfH+oXjOMzE0ulOaZtskB5/Qgj8qQIyDbelW912M
1OkUm0TMSwitekZhyyFQgRcr5co2J2ZsrpaFNJytNh2yDDaJJ9mkkcgLSYsYmeU+
4z8I2QYIICa6PDkQtR+sDhvquip1t8RPoEi5QECzglLxEtp2t9CcBvxzEXlX1c/U
fzbgQNjd7pX1qEOm/ydY+N4x0eZGzy4R567t08IG72Flwu5etn8OrT2w5q03vzFi
MeFHBPC/EMkwkSiLGTgcmPUHL+2xBgKmZOTfUfqG2qIWPF59WdH4K3Uzo/xwY2yE
VUi/xpdNo3OiZ5o6OiQk2h/QA3nuKlqLQohsPVw6AjWphMwxORVXoeh6AOD5YipC
DSLibZBa2OssLrfp9zeAN2/2x5pfaw4YNM4vfXk763ryIY5AdLckQNEfxBPnaVFh
AWMGaoArkQHdFMt+WjXPInnv5YYImD99DOVQt4YY2ZSwqJ7nH42/kJ4rxcI4waSD
caImGaXRwfvFevUi55TzFqOD7RmwlvfkJmvObz8ioZjLXAKGo+q4VX6IuM/3JCZ6
aGpPfoqDYGxciC3nA6NLVx5P0wWm4DiNDOue0BeaaE7jF8uRse+YI59mi9fLAwlg
AudcMvj+ugc2KGoIYfL2LGAgi9C2Zhj4S41EVTp4pbwgbnqyFRiUng5Ldhp++oaN
PVuWN+E7x0/BlXeyncba6cNpaqp7gK+155oLzxqeVmpcf+1jAG3wOspobeGmhaTg
5Spri5dOcJcb41fpzM8b4AWmiRpxJzYqUU4Ex2LcWai8gBudBXUkxMIbiwYNr3Xy
Ffd8xU8fP9mKWGE1xy+U9KIDUnsQsNuxt2KY/+S+74qSHi98ee7cBzw8sLA/U+5i
ZxN/cw7h6dA3FsKeFcWkQvrrYihO1bp0vHeJdnx+cBfS246RiVByKaSsgznCsL68
oPuxgUqjDL3G78nDX9Bd84kHbClwCO1lmNge7Eg4oOD0h56LtXb28avxSHfTnP5b
1ANTWCYgu6g8pk1mht087tOH3vitlSgs3okP/DFWCBq+IwyNL0/1iMyYghM0oBm+
u7Qxi88BvwbiF6xRdBs6neYMSwjYqsrlHU3ZTkjPy1kyi9uZa32WwBIPeBBmXSrO
StW7pgxz534f+WoNL96jhzJPNSfPqaZAlAcgKSsyO7O91OOqFSGNsapOXI6KpcHH
iblvKoDwRD6ktNjMyTNDyRta9YeEgb/Rj/E0xv5muwjBs/z0WE1fRozN7tinNI0Q
g/vkYWxb6LgbZskBjt561ezXzROG+5qpC4CaMMZJvB/lEPfL46+SkF+I8tBy39gd
ojCXT1P1XTJRBWmaldLocbnbrAGvVhExj4S+8TIg1vgscHbpom9TUlm+7fwtsjbC
+z+r5vf0LyPBcytfQGA7KxyE0nHyiqMRAYbuGg1VyWBQrSvBi69Sj4Bfg515TL7u
waz2QZQ/GKR4HR8mOHy6/9sObj+lAYhVyJcxD78YewI2yo0NmU7Ft/lZJ/SXjVzW
MsziVr3Z5OMflogcJh/Sg/TWrorq8hqd7Po1dDfvvzrGjUqgzoAuaKFvQKd7jk8l
sHn2eJ7g5giINBVzv8xW2br0GIQVqjyi+k0y2ROvuxzgBgmdUc13HavuxzN2cj7t
2ZXr9kGXhgUJikLZi0KcxWhyq0wTM7iAtc+qq8rANd+q5+i8Qyz1WzqEABQvp4WT
OtM1mehx+k+p/OF+VuxJIL/Ha9vtKrMehHxg4GWCBFDTMzhqKrSf6u5tgBFW8Uz0
JLpjfdtNjhbebv1hfdhSSjPTlRiMJ7lE29PAe7FWVe1TjwkiEsvCUuJGVvUY+mRT
kiQBBwy63ZCcKGrq11//VN2YyFHejpsNGNd6R9HwHrC0kEqmtwJUpOvgV0U8/4Vo
Uf/FD3XPHiN/IduDG6lf57I/I4wdRL9ho+9uJtHXAyiKd6/YO2LGVtzUQks8fuN8
omYlAU0NKETMtDCzBhQSNMyJQjyxX8tAsaw9UCdKv9vRu6OLj5Dk8psqPG86X+Rn
Vu25HtWoRoU3rwJ5Bd5bFjjhBlcgS3ba6tYkPANuttW2+LUP5iOU5I7QwkoMqD8K
7RFQVzxm9QKc9lp4hRBnvp0hjUfsHIpilGjrhjvqUp+dVePsBOjA/5cUybQQ7R2t
F5aP3lMnlBXdS6yJhmH8B5HKtnpScxjWGM3ecx8/RNRp1+uLrvglVJclYZq7oT/q
tUnb51HICvT42zUhk/IzeRFNRbU2Lh76YUa6ZYWsdJPvDjOU3u3J5RJMsJB3rZBA
tNd4aMV39e+awhNPo5R7LgDMy9OhkAwnD0X0ol9SPsHU7Rzcv87kp2AeR5uPss7e
49LONAsdusYFG2C4OdWy5/StDJ7RxgCe8YzPQP3Ne14OE+EY+bwQ7MoSq45v+kOq
4csahoz4Gklqxjm4GDcQicD1BLzSLG6Gv7VY8WgN0I+z/QhuegTBSVo7XdMxGnsH
Vopu6SM3Xohm7haPBmb2Dnvw2VzS8PnEKw/GB+e7s7mcV8nRVAHeYYemfcK45w7h
PYkALk43JjtC4XE3gTVg7X8EL9XyR2QSVnN3h60/1h9XZ+vaYvhbE/E+iHXhOAh5
j4gTgZh1RiEYf7NVAVnNR4POWdzBuKLs5noJ4UHT6S9FZfgFg9oL+31wxpdSNwoo
NLuTzyW+PCn7LBdyuSxDVjSyK9eJyoayotUuQhDXlHevyDOQVCmwDYaseMXDV1jT
yDqp9K+kzIth3pK17pnI5A5RFPNpjuLltMQbsj2UKLTfZx+4x0EiSH8W1GWSo64O
Ye6xEWnS+33VZYzwtP7I0iqCt/x0bvEGpYWjqxnnnzOsDO/jKvTVCRkunTDpTghm
OOxpn6prHrbHwsGIgwSdkQxKq9jzayh/Y5nzsHOVOawVoG9iJpDlPqiCKoyi8J2y
g4rtVN/vIh4TA/sJmgz8w2jE06Q3Vc8Gx+87cMt8Pc5G6FMtuClUgwXkeuE9gJ10
e2xZ93D/ozOtTMaUFjEZooRSaXzKkDU4rMGdHIkgxbNP+K5q7GiOPRawT1OJSH5b
Arx73keN1GUnrCyfF8LGx+31JF7UzuS1SRDQOU6HYM9VA4vR7nLmes9ZOpd3cWEJ
rBuSZOxB5wwx95jEd9qH5XQYWOR7OQie2Xt12jow1+BNUKPz5DgJrDrvlo8c06Rv
v83m+D3ZDGf+rN5apFD4SyIf3385SJ39zzMDtKaOsT8NN4acbKatBCHhuI4K0qev
+TvzoJ7NglwDPsUNq/G5jzrb1kbMAQz1+kL3wIqo5m1phuLTDasNVd06lSjsPoBe
0NAarpOMRx+Snky8lsmJpdnlovHJwoVknsIciweTa0ZKpOIBl+BWikzpnJT3NvAh
c7f5DHITHIVK1c+fLTkb91MbHnEKiA3mwDCu8FN0CSHKd8Hzyag4Fom0+PXdtXkA
2IoO+3y3WhwMjEF4gnBSJ5maOSH95TdB/n1A8WOmmLPfhTUk+zCyMpfXk++PCli9
HoedcPBjV9MzQ4iH5TImILYEYqDZ3FCwLK2yotOk91wGahD1erwIkfcZa2lM5cQg
+5bHnvWGeSGnwfw+7Ps56kqWcX+xTPFsvTxK1t5Q+NALMTjZtj6muTwg7fj+RwOx
E+z7M76nTGrTVXguncyO5NmagrLvFIV0Xopjiim5wHECstsPWFywS+vx5/qp8+Xu
+B6TocRrADkZ5lUgwwrianUCl1x1dDMjPSUah8LH5arWVo7H/ODe/X2UZSQWdFTf
jpXqs3dPf/bMoVlO8YW+v7IoKlzMQNXXkzr03DUBgjsUPN35qsbGD54XyBFGTG9D
ZYFe4mFGhQ2J/19lVdJ6zs0PLidNzxwKbSlLQNFkMKWx4errygshAULvHsRWRRro
t/2r90lcs2gA8lZ9FTJSA8+zd/pK8FnOpKKiSX6QdnlVABO7f5fBnT5cPBg3pwP4
6dy6w38f69zg9xLrWLGYcN+nrxsVHdUsaV0an9EiHftg43IgBdv6yypxV+lQFXaJ
4p/DFXYLQNXM9P7nBZMrVvX0ePL+yscC1u8cx9TVKJDhWwDdbU1c/yGmNUINhL42
D3TblL1vyHLoZxU314iOp78nFMo3lVC5r+BAtir6YKwxKTTZuSb9dn4pdBZXGb5/
pmPs4rPa7v84KO0Fqd0tLRCxfK1MXm8l8WebcFi0ZBH1+VRUgxHMnEfXkfSHJvIF
UyZ5+Bz91NWwhN4DjUHn8NFfIUJ8XYHt9iMtzhdCqeM4JlqiBr2KBfIgespgj8Ph
iQgRskR4HvqQskDwKWw148Z9IfFbrMNQIhOG3gwEWBlD/1wgSZvCaixMS5kRJQzh
k0caS/L22uBwRPs8u1LXDCS8zkX0neVN8q6vj6gmrJmUdSv74bgZXEYOqvxtpDlN
mbmYNMiytFCTx+UdgwaHl8pFc3rIUZDTfk/IZ9wFErr/5StvNS/eUJksdeVoygBu
2GLQxoJ/rvV4BakgetoLNmbM/QFyiEED2xqkTs8vCNnkvOI2bpf9TFNVs64vBkCK
ivtDnLeErSeCqynwATuzQpAA75tdyFwVta1T5WGsWJTHAaJgRHuuixW848HOXtPC
07UmGFqrvTWAbzrvm8/UBU0mex1YBnu/tVUY2QsqQLemBAx2GrQgdAa6xLbR6qrf
TZvE9HFw6pyhaRCQHF7zhxc/CjbTNTSMDWkEcXSmzGk3bgajjByW+gKG/D2mmMDw
W2Mjy3jNa6H3rmYiz2LRwCT/zrxYL6Uv1v5vjRg4SVwLa56lMHwOprfAQzzqzHr7
myvbudY8FqaJinusHCJEczmuC0BdvieIoNksGzCXsZXTUGDPsRvvjxRm/0S7aRD4
5MG98uKltLOPPsrABU4k7OlrZooq9RikL67ArcUPeTq6XuYR+ZMKfDb2R54AXW+x
XMWUsrpl5BGGeJzvjF2tRRJL02chGKP6yqWuS9i0JqYvB0YYFKygA4XmPGWNfv6w
i1IOAGTE1cAxECuf6ltMJZ4Yf6QuYpGWg5dmwwPX42RGd/TLgq1rAr8NqSanw1Dx
qd57BZSqOfMRbtU6RId6/5tM8hQVwGwTOQINZBgB+qAxBGcGWKQ9TuWfqBViG+yF
ZqtcEvSWxwGABRrBunoVTu1/IhfYMu/MGy7pLYVkSnosaydxnLpcV9+kyul0sqOs
2KnYyNvUtHLm3xHUAU59uiRn18KE4ka2ayGnRUZa1HKpQXVfQ5SYJnPLc/C/7Ebc
Te3eLdFAkxFi3tQnIEBLLRTcih5N7mSx9PWPReI7yxFr5FUUVxdE9+t0grUnNiiQ
H39/deru8pU+TW9wOOjbsFjLhk6bHBLLbyW2FTfI5NJ3qulE9D3CzK5WzdP0c0kq
tmXetsKC3qfSkz9szS75ZQvmhEQ402YJHMLNKGGK4POHi/FN02pJ/Zeb/f5FLf6d
YaISiSkFF6Wsyna3O1wRbufO64jczXsk+dikOMa53UJ8noPFUiCJY9Eesb1OqfBa
O/DQMldixAwSxmrZ9gowrZMbPSji4k9sh1axTOv817KRMs3fKvS3mFqe4g4j5qn1
fDleZZYI2Xpn7a4cP7N8Z04aIEAqLpYSfaCn2wDXDBzBQ8QzJMYLQ+aG3WUNn/6m
o9XgsalCs4tdY7Cq69FzV/+doVKys6wCLu7e9BzOCFkpWdKfqcTDqfDVSBtd/7YX
F11+RwMrXPKuyYu/IsPz854skO2s2ZAyYQJSGM8lPAXG9PO1DDWyEj1lx7egeKKj
6H6r8093s8A5RBUH+sXfNCj3eYkp1glVh2X9ysCV048+TlMUt3vHQ9azsge5703c
bfCDMJaYHstfh7DU4yIxnDZ8KUAGopSLMJRAqHCJbf1Dqw2PufjP1tETXyPoRvkk
ylWYpnrYNwFOUpsIGDmr2tfGgpHOQC+MUbmV16Gdohbe5UlSkZKqD09aHubWL98N
wI8QVlmEqwpOufSLp/93eIafH+zm03bZn+fsURQcYsz9EzPY0axPKNcOKV1rMYyn
au0q6A0n1Wv21FX8jFbEeWki9iRM5eoYClob7PHgbO+rczo/jVsUjhtQEq9W2Xa1
uRX/QX8bk5gD6M+ZC4am/IDAJLdeTx2D1g+my71tkIj3VAYW02w+YdXQIplVKZKl
Sx/M+84chfh5bueo2q7298PFc3JLtnbeCJMLrlF8MTGgAbmMQZUIK7FvWJUwowfm
SJwtq2ZyH6qoorRO50PZ2JdvkCbCEIZO2/NEBsHx+UGDc21sr+FW69WqZMr12lX0
eR4OpFjKiPJoYn5lDrVtc+zaGLty+G208xEILdiYrNCB/vKb5S8w4oDBOWcnftWr
SafBp5111I5Vegz+ZZGIRNqi5l8lWpmsWGbrLlDYV1EboVLGKLxspSm9qRPQgrIL
56NEK0LAGNn1la6UuOajejCeauUR3LYgdA66pBpEfWiAbT/+BuPEb4x4MBwdZ1D9
YzLJnZ6ucy5e255EC0KOSLzq+Adzi6+jtCLcPOHS3lm0wiaSDpKZadDlwje+i4XA
8cFYHQ3MaTFQF26pwJOLBDKpNvYHPF8Ujlvmha7W+++5DhoOy7C+9YTzEs/IBWty
9D/0iFGleSbY9BCISRTtRLnLlDP4F+PWXfqcrAviwfKU6gb3WrDyuYvwYRKBczMH
uin4R345no02JWN2ljrHV+4iCgVI5T07pE3+2d++VVm/TdVb4FfSq/HzIsWyptIe
hR5fj4QYDwhIKigSoxHbnm/TzEwy5eXfVlMixdQBuiVgbtuhT0x5DhgZvyBeRoJL
Ss2ST/xUO/t/S37eIpRPUOGUPO+CFgcF/FDg4CBMdzESlZdwK8r942mKVAqKDoHo
6V1uMRxnaSkXz+CPo3J3WFoJsmX4wu6qbuh/tpzVfym3RoJVSo3J3BBRmubinoLh
APjSq4Ce3bIxSguz8kbDLR3XIGLqJG7tbT2tSIgTAgK+qonYwrmlpVfUvqjNXw8S
MB2W6Ouz7USR8ByXHm9VZZOiBzGBemwjGl5BCuws49VSVl6IP96JVSIozkFH3fbv
EqCXeUSbDiiNdWYHLwphzn4d+6xVu140qxiaAyP8xDSY5ucd0S7hJR4DExRPhVDz
sDO3fjUCovjxK4bigSZ/t3ZMLuXTwUN/QTud5Gi0PozdgDjKFnLFqoB3XrT003yY
2BCfwdPD1l5tmuAtFkY5PAD1daV6yfmCowr+LpmAglVWbZPA3sG4bv6sz2X8Fh9o
S2f7SiZVHf6jBxB/VdiYr1zZfrG8jV8xKncOc/G9kiPEpTmwTW95JuoqkLeS08eg
PjqckTM9+piFf+v3zz44tltJ78lx3umtdIGLD8TIWCu5ZJ+EWTU0+h0oUdAXAt4Y
LQkwQ5phtjS0aQIXLsNQyTVbTJQDOUXeyzkrn2CAmxYe91M/swGFKtlBGthrKGed
FCsMIRYfHjNj5xCyqdr3gas7WVgVq1iIh1NSgu3caHU4yFlHCaFzecIJ1wCdWILY
jBOPPBMUaSlHODXpwT3Mk30uvwGxZFhOvK5kxKl7pOrNGz7/A5T227PHIYunrpQi
H9Lnwr/pwWULNhoBKVvrkf7IsbJCbfvmCW0M8XbUCIUBKgPk+SufpvIikKsD/sS8
7ExJlr1KY0BbqrwNGzQSTuOo/OE/uNhdBg7WIp9SjdtKXTjCifEi4gD71W0/2O8Z
BrYo9FGl2+Gg3sP3832506YEFNjFw+Cr4+1O9ZkB4SbL89pT+IsfumUSGlLj7/ks
cjLMXXaVCRxq70kHVciI+J0Ym3t7o/u2QL3J/ozSzEfTgdzPuzJDQpUqbJuS2QEb
SPLIMo90Ubkx921M9oma3MygdyK5ve6twOYcxRGCEdQLBasrCFGtiElI+6j0w05l
R1/BIka1O8nHtX/Fnjkkth837fWBuAR2ihQYcBkPlRZINrkUQXB6lv0GHQwxrSb1
h1eUJ+h0dNHYn/PQy2n88G4BvcT8nIhLFneyMJoIhAuDHHpmTkTL9FJOEIeLsBr9
mqgFIBlSBp48AtYvFwWR5AkJq7b1dFxyq/1Jth2yu5VI+ibIyHIq/vfBDld/iSvx
5aI4MpkkWEjkDlqf92bRuqzyxGJIrfWq7hPh8563FHFlEPSwhbrdflB9VPRluyQr
Ygn7Hhe1EmZy6K0HZUmbcdj94AvbdEwLAhi7Ay/XhXDs5c0jmLReHtBHemaKUpvs
dY0PMikfa56NHyOxYH+TUSfj7ezL+emU02aRYO3sEjVIPtMkCbblvkQoRVAyFdD7
fhphVhV2xTpaLaMua5PZF2ia+E8T4vw/wwEC49IIao8vuuCMFzByR9xIBRT5oqvm
P1LiTHNQ2mrqQ1Qu4e8HhQjTV4DTkY1bZXFH6ko+wjadVrQbCgXYeooscmMj9jAJ
tkKPLKMDi/bitWxAtm78tuia40FXe8MEWWD31Ye0bSDo4DoKmEQMsJ0xUZOG6uMF
tyOx4f4rIM6BvXVuq2SiKkiO5N/ZrAjpsDScGR/UPRRdbUFjJ1nG/xfGhNUBNijz
B42J0yfxFF/owhabOPoGMad2cCbaBHbvYcoRsmbZMb38bHp951QM++I8U/6DttPa
Jz/y8FDgDSWkQW1a54A7vjk3nq8dxYnN+QkyCzVJMyjA1X5Vuo0DmTH20XJKwJCH
wV4QCD9qroYZlG8F7viegzz51yQuwCyMZIQIvB9eHfGXB0pQMBnfJeViZnqJU27/
F1G0q2tflGbjRpGVEWcxH0Stg8fMRnfv9WPJJjq2GzctComSq+TkVKe5BoWEeOG4
PinVerIbx0LFpje5VjrlJ6klVQQ/qBID/Dn29h9NkeObnx+ELzdSgMSHDHqLVWCg
2RvT682+XEWFASTyRc0xeIBpgShI9mgQvXkf8IiEY1oSVmZN1+h+36ECajk2WTDS
zT8m6zP1/plVjCLnvGuvzfttiASAL8QOR49GStjrAy0cI/DnpwMIATUw6yJj35R3
/Aes3OoHzpqp9bREqChheuUT6vLuZhIyuqIOoCAOVI60v4zubknnzc2Q5Pl9Lzqs
M55oON5AiliniyCAUwl7xoPxSbSgjvoWwXxBejv3TO1kqfhwM4R/CnHdT0ydT5Rq
GsTLAI2wbE/pqx8nhQnLArq0jYNFUwCRXdAR/VakNysniJV/IVnhOrlxiX0gdeNM
WKVZBFcXsCF0wtVUjtKMSTpGBmWfg9RalPKGFWAhAD0X09jw8mfOWm3+qz2Poq1D
1wGHc5aoJX7onOVb1z/uFWgwFqLoATeNyJBd4zcm66Cll1wD8rbVMFTtUDg+O5MY
gSyMeNok9onoFK3sJiLoSy+9MUTQNL481jJUbjyk9Cj9C2sAGrUKWkf4KKW/PiI1
7dcYZzhesaUZGAlU8mm0F0At4XKySqIm+0QTJFjl7vXIu/z3aUsKgcul2rYPWYAD
aiE/I/hi/lPprVcEhAbBrHEmmR9xhCax+1913PtprurhU/+f9wB5OyUCLYuebTk4
sl+73ht0gf8EFIE02PsrgJIL6khNioRqZF7p6wb0VhKW2DmBJ3K+NsRfUrdIfq6s
cmA6vwzwaJKIkPo6tmuLpidZ0oRuGZ2540DqVgJ17aKC9Xv7rvQvXEJGOuQZ32bI
6lXqNYsqQ7TuuhOV/O8K8svWOf1Q5zNzz+F6dxQt9YstQlk+KkqhYeo9CwZxV1VO
2MnYP+HxlQ7t92U8Pd1Wjn3WDUCxcTny9MnTxD0wRoPcuysZQiiu/Jhvl9GPcTGv
iobHMCa4j/7GZkiyKqKpxAGBYrPVT7rcdaeluN2WzU5jrnoNOnTdcNuHCx7/5ktp
XSPZCLZcnr+cxx5dxsHtJpJDTiy0xPtIkhYFHeNNMSbJMFNIck7wUeX4HvVROoVP
XbUG/vRJe/JvGhrZQbih+dsApMLKvwrjiu2vmu+N2nNkkPZyg0BqCZriJztCq5tS
n4H6TqKXe5fKZKB+zF10MoujARBUlhaI7YAw3I4L/FYdA+d99YP9/uM321BczfA7
kfPx/Guv8QBn8OrWWApCPKNxVVcUF+Q7iHA4soUhkqjrFq0zvtadxQlIvu7zAxsy
GrUk9/8NsasmEXws8ZFMhz5Kt49HWhmshQJ7bP1F7/mxZTOuTGv2+h8KYf8O7S0d
AxTGgBsbRm9GK4Vz/UOnvZJ/5kLNS+kk/LhpJLaRT8AyqRmsPOmhHIVp4d5vGXgs
TrYvwqlf8qiMw+OaoJxvKwGLXgAYtU4oxSPot/afT8xckkVFeGlH94UUSF+Lw8Jg
gGXOFc5exDprFY+nUkYDhxcwumyE4E4iY78ENDHWEqMHVNyt+o4JePl7pS/GsnVV
XijN5j8ssTyDB0x50xzvjDcfuagak0/6U8zkGuNziYPmaG3jZRmGmWeZvPVM02kU
tYInljCOixOx8VJGLHfPSo4Eqn3+RTrdoq37yv6PolmskscBAcx1b2VL44ABqe/y
23P/BWRiMhwXS/sY+VdNtngP2iggE6GZqU1D0b4hjk1kVN6GAk10MO9ZwrPnGRIB
w6llhTCcberFrZvslxVC6EbvP6YgLdPrMSeZ45Fw3toasZxqzPvajX0Ox8Vqw1up
blleNWAm6yOiWMdh/TLNiAsyPDo77MaRSccU9abzjXfnPSabzg/vgbcjw2ktkWPf
0Pt3VFdSwEIPr8tJsuBFteYKrF03MRQwDOIu2czRCcKW85NFcCwLVvhm/7lI7OUC
pHJeM5QN4JUmTPwROcohThe4AiaCNUIVeQprSa62sMcNZGZFP7ZFpxH9B2X66tt1
sGJL5j55nuBOX7cMEfRtCe3P8YtGG3f7VPfH56k5X/j2ZbfIzLy4e59L2j0XbyBq
14bg2NFQxwZk7tmUHYl3IqIdtMYuYvU/tk0RSG6HPmFF0HA31g4kGI9NuyjOjgoa
8HYeN5lyz4xlgwwqSRToow1B6azWzJYLyHFb7Aobaff7ZwvYVimoML4QLaXqPVjm
/kREDh+nQB26va24nWa48NJFKQuVbND5VmLzjaQzc8+tslTzecZYQsLNntvrQvMI
2xDLkOFxKHs0o35DGoTYL/wqFfo5CTO8wlkUFHiA3xa6hDOm7PiSM187YOTVXS/9
5nAhLycsWSrqL8VEXDqAw0dnUSnpsTsTADU6YvYAbRiBzPlI9J5ErAttPf/g8hy+
PIhjNdxSG7/jjBUYLM+5Lp/kqIviHc9fHiUHQYMGIqUSde1qzLuihpCK5yyJ45E/
SevBZjzuwLCxub0sdEBx6c5Vn+dfZfb7BhSrZ420YmWE0ikZkk17ibFO50GQEST/
o5DA0b5ZcZjzkkIuSTxJG/7mGJTYnf09kmyA6aRwyOsn7TKxCHrZ50GMhYxQBgmi
yNgDkNCB8LfM0b0/nwI3RGWFmB5q1V8wNW6fw1kYXysKMiLBjVeiVIodh2CWutMS
vwseOdkxeqCjpEO9+aNo+EJcuV8ODFhNrrkdU5FD/6I62Emtp1e/Ec82YV3bOpQ0
No/mmLdefbrCZGJv9npm+JYdC2UDDWPxo/I52OenEx44wpHUoZzmyhZIRxDzavgy
06RcGv3st3XjK4lyy/pZDnuA4Q5+Y3FUBrt+h0hwoGzCAhXXb7KQfEAKeecyVmet
LLh5hrMpRu9E8aygAlmoh4wWecv83QZdCJFwyJtWyoiEe7bPZxMlyjASfaSssbYl
StYvz5VwCUOqMYRSmxB/zyNkVoy9jEwDe2uyveTl8XQekPWhNDSPq1UW6cDXxHyv
lItRr57pxSvPv17nPkMUyzbmtenL0fR+1rXxnxeQxWJ0Wf7kawGyHpdWy2EwxTjs
6LpW+X8SrVqn9aDRLT9Sq8MCLCeFwGlm8//JY3ZOWX9uS8M1/u5+l1LCWDgg0Qp9
wE7gqxyGX+jXRNCi8EjGfWu+UZSWVmbK1v64n/RKgDOeEplyDjOAqCJKgC6SpUFb
IpfSwmcKIID7Y4zUe/joki+Dn+HtieP5wyKC229fLcRap/R1sIWVWjjjCZ8krRO+
7oihC2eZ4Pp/DwvY/o6nxdpmN0b+ZSOTMZr4CuMslMtm7niPbiqojO6zY1J37KAo
mo2pPWyf+Oi+0UUvUwXODtQDYvB3w/D8rMYO2FCux8bN0B0p6/mGh+gq41SRpVRw
D47RrgGWphtGtYUpxDGtUyx9uL5cPPPqcHjiOycD8qf99D+hqmm295aKTBwB33gr
fpfRA/PizdLt84l7PTjDaUDwuJa+RL80tlsU3SpuRYak9/fg53TtbGdGnUAJHs/2
XsfZmjZJwXidbyGpbULFdFYFpsuDYismiArVookJg2w+iZPglJLp5n9Q0+6GbZrt
T49oYgGf5fxsPh+PoGEi3m1xAU25d2JHXFfmPapweYOXNQJzXyWHVmfSeeSzBYpx
78+Xe9NUA6Fs+dNiPUZ5JUWktN8PrqMFMERKaoQOigc1w4LQ2Tv4NqiFDKbxu+OL
jBm1S6Ui7ib0iOSFgVbN52K1sFnkRXb9mv4TEGckrp9JMJDPxU4DRuksEKNvPJQS
TMgB4ddBT0N/P1T+ntdyEInSJymIYd+W3kayr/XVJNx6Tre0kI6zf8OhMaZ4O8Rz
+eqtbHo3C6B6Y38SqksCH1WMonhKfKOk2J6RMyzAOfVeZ4cv21JqO9qL+JmHbnkU
WrTfSx4P0EbJ+J+fOsl2qnlDPsEUToPCQe6jfDqtNFzCbaATqeZIOdSSS6te2zr4
dGlvld04QR9FzH/87BYXgGFaAEQYLG7yZCcG9k+EnOCJB5nnp5BHiu6SpvQZiK+v
FDBKEbQhu1aYAL7EgV9DAznuYC9Bi11fQkZRZ+HhLBS8hRa7+fZv/Btz0OrIA8IC
MFl0c6HHi6fc0KL0mYidYXYd002PcKTdTFXIjiFLBbqYKE5WaWJKn4zXlSLnGxxr
+3KJuKw+OIbH4aFnFuP6yLwKE9g+kCbSN8lluXlYPaXwfcJKSyTEsSz/MLTpo628
Pkp3RMHeCpALaEktiIrWQUYAcsQcUe+m/4E/Q/ZTq6+uHXor17KOVh+pBgi0bjKs
6+uPPooI+EZU/Xr5op1miAlkbfp3qxxHBcNpx+AfKB4T+xg9eBXKnkmrf3/AVXYh
7UR+bim0ekKAZlNJTZxtmNYiS1FHEuMoX/igaPUDwy+gnDIt/Up/DavTVaZQ51fE
Qv+URaav2B7LjEjOM2nWLuKcozdLSKI7M6v553Sgu9f/VycNffetR/dgMmaGE2aa
a3NY4DWKv4zxbSpbx+Ae2sBYE9G9EcCY3LHw02Ie2QfELZ4coF2MjlHmITSLqXNj
gsLdVZdajmKVpPsR5CNygQQ51JVd+r1puTez6WJnrl0J7ApUOugJmoF69JgJLNZZ
EVuV7WbvdtNvgxBi/S+fgO+jYT6dhTDw9cgYN/Xw3+63JvdulRwI9z9WxAbMqGay
5529u/7su/7xozxC34sNI9Z/sXA2p24LD9Uj2OTrDGJYZe2otqw1x2yALRwlWvmR
R3vFqN/LC+LqQlqvyzp7kPopuub+AJwuMPEKiyhu7wYsHWZv6mSVy04OQXj7Geb/
XxyPI09P2ehdrO6z+D5iLp21LPRfDSd+pzOKJO7Z5UALkq1W+88boJzRkY38vRxy
4mdax0SodE0b5DiVaV7/mwuFu9g/DLH7e26EVwsXIMH+elU7fXiVDIV5OVHDtoAM
V5X2LOVAFQthUTKVDLxYKHJ77xCMW9PTmdIGUSj1kxlIVc2BCFN58Ak2wj8z/85w
hOMcFhemZH0nWb00AsGLP56X3yfgxGZ3X1CnsncvJunPqWIkeuh0JMy13DM/X6h0
iVjLyRfQz7oiKWTR87AbZeszTNUaF9aLz14hmpa6VP2HtXhm6JiqJ/k9J/TLRfmE
v3Z76ZoHmMN66IrW0kzSWg/ehoLcNHi1HrR/mDDfLDMuOUkNPP1a1RkqByrhqK6V
RFXRk8XhO5g7yAePNjuTAb94z1Ae8ve+3U+ibMbqQFuq6n2GvKk0LMABqMKgXSSO
+RWu+4fzYICOHjMiAXo/3TOn8KDEVpRYDe8103cJ1G/dqqCPkSjoK21q7xNilek+
8iH4GOuwFrq+puwbC4xMOlpgzI1Slxv4XgotuWVtl7T/9wxwd3IkbJUAupJBYXgJ
oCJgloDjvqKlxGSVxHgND5LDFpdMN0yGxFNuSsXDjIJdPOpqMTBR0O+n8GHt128I
uVmP3ufAC4PwSoOHVtuUAyzP3syvxX+apLh47oN0KRPXSUTwvtGz9hFwnO8fmGMh
WWNA+bXvRoUXEc4D0bE6DemQaB6Awxh32/kKSwMK2F7tPNwdhuJlpnhnnP6kMhJt
m6Xc5LHpsEmVpWzixTCEH/l06bDPzMPAcjmGaPyjRR3Pv3R1JkghFQaXkFtxfcf7
k9ZyWdaad6xIs2OGRpQy1DYdFF2ZD0NY/Stph4as3K4iAnm2G+HZ+xbEPb2hYaRV
sEP2SVuGy5iXUuaKYNQnG2jc1Nbkl6dPzTvwYtMOyT8ozpb9OyTKr1/dWTmEcTxy
c9SI2VIKLXzAeI+mzYyFKgA1pLGuE2nDASB2QNs+up67HeJLgrBOyxaSj9OPAOHe
7G6kpI6jE5hKCFvMugQBpYJmu+mqVyvEq36am/kzyyB+VxWZ8bJ8h1GiZ1yEmCnr
y7OwcB9nJxD7XuZY7zxp2cq4AlRgqt3Bq8XZXd9jdS3nfJVkU9nCTR+/2ZRMOEWY
LEyFqMP7DbWSMjIZrXsBPbUoujbsodwlHN0MToI4F2VVTePqbwDDeOGwdPmcJwfZ
JaVaDZCAhnPwzGgOJSknlcqycjvTnDyDr3gkQ/km1wXIitg/xf0amgkm6fhPYvpp
jL+Q76n1c2Xigj99FBfEiZHQXvGjubI4w3zOJPg5f4xgYmIMKXmZpNAdId3jXh54
bt9IQAzglG4xKr5cbKCJnikjGuxJkV/2YqK9Sh9ALuXZ3b63B5+usd8VUJRyG0iG
htvtYFFmlfnBCrjhSR64OF8RvLwr+E2byVQ+UKvZSwOkow1gzfHOzZKSEViVBMwo
Vu1cAxkX8kCEoj67h/s+RVlXMKLKzPYAejuIfO+O5vQ39LVW5ZTMXtXu4TnIfIS0
bVkDbGFMjCDE3By8O4u2Kne4eJVMmJPWx83DG9cOPZ4OlckGPAXawOnPZBCagkNx
/aC2DnYoAGgGdwVKmIVYnzk0uYBQOFSqPG7dDO13aYtmEStE0ar8SArrw1LVZsLG
/YZpjakDExAha9WEB+0KWzaAiQEB3jc+LU9XqptcvfQPN/fyxjWvIUA3C9t+XY8t
LltiyBltgIz3lhAYwYCOim4MFGcbJLatDcAx+9Mt7sYdRFAIN+nwmxnECK/SIh/I
WW6vz/Hfw/sGB1lSBw0Vt/VPGt6FRVcoMVJ++H/IUwCdmraRwoURSK3ysZHhUON7
seiOFte4qnmIHypPMCoiw72xyVxHZfHtRrbedSojvdseoyluu9TRUUYU5j4nT6bt
4yR+N5V1RuUGlYB742KiT8o2h6KZQsL32CoQxAqf03UL+bnB2W4Aqhzxp9NAy029
bHLU4Xlyod6fTSxXMs+yeO7exKRsV2cP62QYfJkCxs+Yh9TUu/OAXxVraZuI7CTx
NiZRhme39PIN58kxzkEk99cKVLnsfeyBkAvTOzYlbBf47yFu55dzXBmmeVSAJtbQ
t8HW7rg0BEARIBTfY8v1HDXwSO94fQPJb4eCtIkwmZ6ErnfCo1CDJfKV4ETU9mlx
14PQHQJfa/3qONo1oGUz6/oLHMCtu7LJjYRVm/Z4i0IVEs1tBGpscAhmPDolc3Bh
RNTEQSeCtK47gTpDwNZyEP8ZhHrS9/KqCCTxt1Xx8XYPmrIwhL4oYXRN1t8gWIHa
D/UB95lP37/ylIPdGExihn8+A7iG118t7iJvk5gKMxaXAcaTbGoNaDdySFFXP1CI
WTF0mvSA+W2UzPaKMapCY1vWYre9Sg9F+Uyz+O/sLQi74zmOgjb9v/nYq2dTer6Z
VH8bAsuWuGppicMWkwPjaoBxBJI0qjTwh9vTFDJgxfTCRYDcQvEeuZqdw+s+wmIX
I+9LV42nQ30ySwzqF/+3+CZlf26ng13C/Cia1lmffUw+UhkuW56CTzeHXpaRnfL4
7HGb+rst1j66u0Qk3W1iA6+87k2FqYK4TylB9R47n+uxDJI9wdZzuheLUlCnlLyA
AMSuyGMy+YL52bkm+eLPTlTZuNVf8gjHGeRZqCEEqgRLiWv86CNPjlYeUey1tqyU
vBcMXqJep1CG4rEtyjl86zazQ44GMkSESu6Aym2P08F2R/n3R3K3c8C5jCRBUyfD
G+zxOi9/Mntijzm5mCrg9aYU1iBqC+O/pp22Yl762i/qERhhlDeihHCpKpI0yGrd
A5CneK1UyvbQHkzepM9big4aLY3oh8mYdl+BJqxyOeyvzh7U2YQxa8QqO7dRada+
R5bpdcKe/0crTQbYhxK5KNDRbZ5yP05d8o95KzeT4nupe9sBIUl/1aUKVdeGuA5Y
C4BbOK+nzikOTVOIiwT2uEM7Fp7oOrOzZqWY71n/UvWqpBJmM3xCKn2IeLbN4Cyj
AiYsRdzhSQCG/O3t6ATdB+eWLc05hsK+fR62NQfnLLjYKLu4B4+zKYHa6x0yTki2
Do+Fr6Ha6YEMKJlJLihnRjypg9QLqPe8AAOtRut4x7n3HLVZi6vNF0WOnlmUSTR0
EN2AfAuG5ys1Hinb69/8I8h1ND+c7y5NEaff1z3UXt03x+ZEGeOPd35vaLalzJHX
Iz6AlkkHZQJf7/l3nseKtxZ9ej2km473AeeBr3oinpYJy7HqvgYhivLG9kz6p7I1
7j7parUTnK9jQgZ0MEsbDMl2GyRTnxWKSHv5h3wmUWIfwlXctYuTJ/jaMY9HoE0s
oQJHxECL7J9eHLvobzRf/mae0EwkBxbII6quOOOLQ0yOBBF/r0x0nOPflFium+3S
NL3nEZvFy3g9x3Z1WF04p9zUW8rn7nqmVL5A4Q9TLu0J2Zocuw+cmVjMtc0lEU0V
f6T6Ul2F/uvB98V6MoL9grrFe9sBRxYY6csEpHRiX6G8Om8ZLrVgZXzJVtwrYP/K
V695Yn0NiIx8eATFC2gB/xF+3j4mFXE2b3Ch4eklWXSJuqByiJEnyzvgtI7bd5tW
ntNLKzKAccng+lM4lJr1ENXP9yB2LRsQtS3/UXmbwgtbFg3hixUGtfx1gTCJSYY5
gGPc0TYiF8/goos9VPg9r36ja6Hoi8rDSEf45lzgHD6lLGHBKA1cGFjPNUxkkEZ9
8QMzBVvOzoDhthluMPkOHzprNBoUjQX9i/cGRqUIFMlKgt5sV6CWqOwtHkCX8rec
0TO4PODL8Yi6/5cILzIPxbHXBFMGxkeKECTRE1lBAstSiMLyJmZyC+KvdYrljRpk
htISea+jLQnnS3t5n/ipI3enkI6j3QXr471KpPMX7r8Ue+z3e5RzzJAGr5BMlOSQ
JcweDal3zj9MAC1Vje/6S7NWth6GG8NWMY59RswgC+pGqHoz7orwcuavg5E6G5ev
9qSanar1vxuA9keZYiwYxNFBdwDeUBDmlEX2vx2hAlRU89XcoatA64IVt4Oi+u57
4djaGJVVkUui0f9hMTkA8qSzUfWlVqJvu0VsOoA6yqVuFsklWvt1kaCe3y4FZc9D
RlTjLdVUl+XkCuhmbQdnH99fNBmYk9w5BpRxghU7EzmBo09RsBpZOWtTSfjiIfhu
Iowxl8CbOlneAhEbnIWrjmAT5QpqheOTZ2/BFbBhGwQJKaF2AM9TpmkYybgR8FAX
HQTM1ja8U1YwrxTHeTTJEojltJvZjzaoaNsixIiF7hGT6DAYQX+DUsExcm8m5ASm
6NzEc0z6Wo3SfAnqvXH7fMq6Pw9pZ7xGMOszzK728XNRbK6sjrqjbXf6c9i+fWTW
La8q3hj0uOPmbadxu39PzEZKeSqHDDy9+5HnSirEO34IFldel+XpZjl18XFNkiJO
qY4WZmp/LaBSFWCavMsoH1bwSfHXCqGNsP19626YfnwuEM9UWU1LBsERwAxyFf2o
bdiEocpoac2xIOyRb85P4aj5MoN6zaJOeO6c+IWlDfm7SpkRSTwCsMeYAAvyIrQX
SmpacfdpNbtfAMERgGOePxYwKa6xCCm5GDIdKypdaGuZGumXZExGMVASXRkYVqNK
cqaMwuepCXInaoeK0yhSoxTDPsFHE8FbFClsS459QkOLIWM+N005cvVdpO36fiUU
c9kgskskp/fq2g0mHzh/k2JiA23fxQnCTpwkpAmi+cpPS5r6Qs1iynUjzsjMStmI
kZolpcPTzsv+NUu4ZxfiiLFLfygFqpLZcZIaMLKE06DmkaekLEXUSrROrBbjUC7w
XYR6Pans5aRX3eZW+GIEJJkXmebPNyxC16Da9BzVgGeihrSa/9FTTBNlfI89qksS
EJ0Vz1RCM583XVMltYT1QS5i9yjQphHxg9lHgkAhmyEh84LVXnl4M9wCDAiMT0rw
+JZDJdHRaFT1i5cIUX1oYI8gd91Uf3CxmIswqiVPXZkVjlQ6oGmMqUQOojHg7qMc
MItiM0OqkM7XXNvO1DjXPF31jms3cTtRiwowAINUQg0YLZTwdfQv7TxAuz65lzY5
bursaWRPJp8n/hb3oi0cZfvcAbDj04gPayL2HEEw8AR6OCxec48jYXbQT0RsGxLJ
HpYOZjYC7FQbsO2fVdZxiVCkb7EMKJnVcsZdisv5vhfkYWazobRQONPDxk5/6nxs
NhZb2LC8zep7Jb2FPpsmvsqwDySgRPpZalxo7XaNxXn8q0ZW1J5oiFAsdaJ9o/TM
227iqV8z75Mf/70BoWOb83G+CudCj9n63OSsST2KSUfxo46xEZklpoZ/njr0hYAI
KIsGHB2LOyIpUeCiYW2FMd0qFIagDWgeYy1BKfoWc2t8OFdXMkXr7l58IEn4iNis
7t6hTZhwEX3vP7NpK/v7cck6HOzKLW3OOxGhA6+LrMQ919ZeTCi3Y3jztuLTjbBB
Zn5FtXhuLsLIGXlyOaODEDhfz+peoJM4k3aJetFJWPbWAq0a/ToMwqEfIqSlZv/b
1+rgE13Y7ouXFUbbbR4UNSqaGgMdDA1ruI44IQAepaWaWWurJO6EE3N9+C+SvAJt
wpSs+aigO9aGdcUdNmcdzlgLTQrMGMoq9krEouTFglMp6w9x8B8P+Frqc+hvUldx
gXbOPLColzQ75Uy0Fv3jZ+T5JiV7Wd6MA9cThmzsM42AzolbO1LgdBzVymyEqpkf
SYLqSDR+jgj1uHrFuSUzrizoakAO3/pA6Ga/EapcztQxaKzLlf/gRQx8wcy5Ca5C
tByPmut6lKkVltdMhhiasCUI4PtW/4bNPkU7GhJDgGelYecxdhhNmyonvkQDWtdm
JWvRZFu9mXQ+udiUm9p2V9+zS6YlvKKrfowxs4W0X1Xa/1qBKe0P8jOU3xIq0dqf
VJMF5i3fgGeGEOnjcW2iXRm2vQlkRKh9c+wIwnrtviwaOOSbI2fJikWP8uLywgX9
TioKGG6Lcj6tiSZg/j2R/QZ/zYGFLqMBZKh1/08HYpEgvbmOV5r4LloQRV/2jW6v
2RcepLQpOygJdLiCQgvc+18omlIjNJG2OouGaXkA/QlFRJygCR49jd9NaNePv68V
oJct2Ed8eronhxb1UjIvoc+dboAT/Q3TmCUIPnUVSYewtIicJNhq4P0eSJYINvuh
iBu75u27LTvKJHcisfGsnOld1SXlVd4OPjdN7sM1WP+cs07BGaLmwthetTSlXYWB
Riycl6r8L3C5cb9Ma/pCFfwz9llShmV93AhoI6PheqRMFpctXSgMtER+1tJWyR7G
8SuS/Sb8PWUyvinixrkKZssnV09s4nt2r4t/gql6y6B290Lu6KBgw8aevT01nL9X
QpUX1XU288ia9b33klSGqsr55h9OSE2k6NDVFwnERMDkPXFtNzOZhYqrPzfvzya1
vfWXaklQHnM8FgLuyUq/Ck+qsMtHyBnADHeFOFNc3UaXrX730ZYbYyyR/Bn2l+sa
bu1GqK2Ey0SDSiilflerPE2HmxA31fYE7uawv1rHCoSezt0aTHX/2bvjPaOg4pla
nnvBFWFZ+5yNE4Of94bSNy+9Xt8ra4JrRwtF1+21dO5U7SbmwmKHCZX8LP4KnuS/
Kgw1vMGmlafJCY20YaE94KOM19y/b+KLXmJY+Qi5ldxYvFNoNwQKF5k7iySasGRP
Nl7TVWmIfihFtgg/b15YHqscQIdWSNGlBSqzLXQ3pyMhDJJcUEdlf1y8WeJGvUoN
y874ueLJ8Ip3q80nGOteY6bRrdOC68r5pOOwajiaNYts+k2Fz/WqFqgz2uj64hzT
rXQi3cW/cMRBYd+RXoNcEHrV6rbZrJAssuDHKDm/rNIH1aSDnmIG3mpfMttt3wed
vfqfARlexcpsH5QR0Tc8samUK/EcKcRT7lt9mxgghVj2yPi2+gpOHKQ7FWUSYaqk
5lT2b/HRNX5J0l4Zyp1ZMxxzESVOHyR7nFdY5ZNJAM7V84CoQLPj5PaBXkex+zsv
0LBbRE1IvCs7AS3saYK7pN5zES2gMnusDe5nYnIhD88YEgmnObFf5dFssQZPGYGW
a9qSVXEgH9LtT64uPn4zisxCoAS4MvVMBXlPIrUqximabyMl36/1RVMLAQSiK0K2
hZ17qkef8tWs459rz+pq6gUIO98bY7v356h6m18sMLvchul/NflBIzqf/96GOtg5
1Lt2TvyL9Qoh1y97pW/Wn5ExquSYec0sMDmECexYhTWTrq2W3MoV8yDyO6VrRZqt
pSOaAP1hb8yvBnh3pdePd26XK/EZWMMu8aPb0x1MOi0Beuu1kg6GP23oEBv69oMT
4g9uGmP+84kvBxe0yuBdnahrCoG1y1fLFyz1s5jkA14/B93f0dvwut7IkYkNUkGD
LoyBgI3kxZm2MiIs4FiWyhx1/5D+XwYSdiAIkiPK+9p/5n96evXEj5UZ6AMXRUw7
eFxuEA9rrbyPYesrk4SdLAqUXAMJdGPTsB4qVS9E2DSIQzfwmhdkeoPA22gfbNFc
wERawiL63GRTHrRCQPSH/EC6xrFWUCBCJDCbtj4Y8W/bXV47w0YY41n9nTvkHnTS
DShYIlCCbLoH+4O3HEFNpYak2mx7WN+GJexbrUqvQtd5p8GtuH8EocUWBqi6JN65
/rsy133Pq3WflTcqV+E0iMivs5znKLodEoat20OQ0Xh3bRZedK/1mNTl9X5Q95Ha
hpUbCHWCHKfVw+m3gSkteRLrAeih/0YzUNktn9N3/R4oSR61Ecb8lDpa+bPmlmsY
7deMZdJ1AdAmiBbkrF/lZKJ69pq/bJk1fmWuinvlLMCccUH1IcvharFeYTe2v2yE
B7KAHVY/fNFXp+etkmnA0oYD0QjcDEafioFpGcBvMP/MRzZb0HLApyxGGa7IdHRO
yYMHB6dQbxTBIQCSttFibmAj6KPBCiO1kzL8G2XVWsUBqh0iwwEk+g/AxAWX/sY8
voSFf1SVm8Nj/HSVWbZAfMHRUtrmtIHBwjG5D4YCUTx1TcZ6mR2Ar/44i0dqes3W
Hc6Vr3hLb3a+J6Zn7htow7PJqZh4tu2lmgY+kcGwaSUhot26p+Zzi6dyxzazgTus
iMiodwBU6ouQRkMiILZAm0P5OQgihJ36BdPVsm10swUyr8bjvmWFftsw6le7KrXC
ZMKzoIp058DNtlSzeG4FTJlntWazf4fsAEx7zM7/ZiXP8+z9gPEfDOZh1X8dsNaj
yoBFK8vH9UqwkvR4MM/ha0bdSTaMVlo9vTHK7nBYg0O+kNT4FEHIHWEwf42atlL1
7VweY77HIET2VnfaOFocIQ9QFQI+FBzSlW0TPFuJSsNiLA05yYIB+fcz0wYepTpZ
/TBbaSoznYz4PYY9lLqrwu1f5WQ7VKVQB/EUm1CgLlK2XDSyXCWtVLdpLCLSnaSz
mTEgVU8u/gAEmsKspDToMIHXhlBLH8nxNyh44Ks8k1gdZ/Qavyosq0AvaJ0x/qzT
1cj6me2QgVbn19I5k1NElO44wPCAIXlnj1xxal8m/HvX6GK4LmWlSgz97mzv26YE
X03518Z9Arpj1CG+zs9DEa+Sj6NHC+IF6VEGoxrP2vFTX1TkmbByGW1r09QS4EMb
tQhrXjVmFlgbM2C9BEVEbG6d/fR7S5HpDn2e85F+HQwVEZf+pzPrBtv0ptfY/aS2
IqeMmEmxUaMppjXw4WLIJ7jROwpm+pAgNIaW3d/VGp+H9t0osV5a+05AoJ97Mp+x
q58gAAx5VKhSatVTvfQi8m8ypgx4bumAZga2wHMuO8qMX61w0oo6B8FcYCBB/0B9
yUmEyC0Vod9eRlmiU7deQ5OEQGtWONXDDt+US7D+5N+TucGcsWc85tWyOYZkK3sS
7/C1ezTzPgpf2s4rnm9tGDbqwzIw7KC1oWWH51w6m5LjU1Oa5oJVWnfJmOsrexU7
hkK50Icdro6PGHz9GDUAvJWlwQYv7ECItlYERhmG025s3203YdHli5p4LNtKNOjS
NsatGI5KjP5INYj/ngsVxEiRWfa9c6JSJxtwTY6tuhUJ5Fsi9M9TPEKKsNIuXUx8
jkKp8tDTeT27ZbMfyim9uPrr1gRMjwD+9XLPSPM2b4uwnbjGvFMjqqkOuMorb6Zm
SNYTEQxb92tU58pj8Xql1JN84cjAdrZCrr0MIlayIYujfKqML2Us9xyHkKgGBU3B
NibW+eo9r6vJmtyDOCHWmNsPF72Y/eM6cCQGJe8KH0ewS5MEI1kGAqnfQsFy8qKg
J19Aflp1pWwNdLDYJnYHFI2kaZ5Zdb5n8lveEOD2RMPYHrdayybi8knmHIupFxNq
u/ZEf3ySmV0cIGPkjOA4IR/0PbCPsuL1IHBuvYHkBPhG3YAwkfYGLiUq9rq6Bb3h
4SOKbt2o3sWY1TmRHyAXTMuFxAquS7idDal2X05lyQ4PTidpFSKX6Ugep3pZqvAC
lc1T4quO/mVytb+7jC7K3ZF2nUz459ZQTtlbiolRF/s6rqcw6GKwQ5k+5lShie1b
+qlEZ38fWwvDLZxsE1HREV6d0Bu8c1mLapXK6aO9e4n1moRku/Gc1ipkhxk/9whA
hJnKPpiLIeGOiV8pGRaHoPmYTKQqnodngqwrb2WUAH9Q9AtydagZPlXmDFkKAmAp
N5aFTd4Eid7kgDWieq3KYxztwCDqcpMCzvCvJYRKQJSWGuVTr2I7A+fJySxYmxXZ
NAHJ+seEE9OyA+rzg8HrS/FR7ko8PoBB1DT5sDUQ7J/f5d1n0buB0W6oLTiCVg4y
Kax6FGp245We+3RgtPnuqwYh70cjkfFY+BFs1uCVodNz6YzTGFcXWEp+K2/1LSnl
otY2QwWsb10j4PsMpJuLb7tCxsa3ZER6AK35jPl0KPOugwcRyT7cN5CUkMY88zXC
o10Ej7pbHJKd6hsJJaYBFBn4RS89Mw0kNO/U4C8ufwT45JeWQmpHJVan+veskbcZ
sv4tq9FVBRdsAo43YpS5AD2psQjoSJU39NNMqUUhq6ZKTN2njrT3xd4++w0FVRZq
ke0bYFBta9FZ8ztrHsPrrY9JHK2liHQFr6516lKrxZlrkWhOE4euQUnYRVJWWyBD
TPbNJ2I1+bEvIsaD1161o6oYPX748HXzcyOsXKhiLdmUqkYpFsaSsb/by1M3I37N
mOUxTsv0XH0s7hT5hNFvRrl3nLPpUaebgV5386uoIyzhwsIMseqcKZI0jRvSvKPA
fmxUvd3Qmr5abLXkPKMFIJ4nLB0e88HedWHLsRZpzS+CV7KH7mj6aEgCa1VD7iaZ
8+KqAbuG1JwGvW2zZ03nX+fe9NrjjlJs4vZ8ZdUOCjMcFV1EeoyIAstDJZjwKV2e
l9h1U4wztyL8R9O9e/mNcJuvhgaI6CiUZcOI9uZDDGyQMSjbBfz8rxphkaM6eJy6
9G+GZC6cNb0jUvcJ2zvdJ4LWD/M3m4N19yWwsdDWadLjoTcWeLSie8itn83xzfaP
zuR7Dxk6jXBFrGxbO0cC5D/yyZ3e/8U5BIoSv4XiAWyAWT/BjbMoOgTYbKYCiQTP
lsHGTHa3OL5a9oc/T/dzDeEVmCejPMbfyKVxRA6gNQE+8F/xQd5aU1hFxpWeTzGV
qE36Du37FA8ToGohE8GloKvzl1Z6vQhY6/BLLi8j6MQw4CHp4t5EI5Xi23vOJwGt
Tk6C18Eq9TvNQ8v377kMS/SkNRdKVbzsCydyMylSQVt3IN9LWefVq+y+fcqoaWqV
iX0lYMqy4b+hFHIlMDrAwywhETa1MtceurKH1/GVV0N659PcAkHsq0JxffG1AHg1
xbg2UaIzAT/HJgwrw4Y/HZ2uluyxrRUhU0tO4ovFM1y1ACADqC/zdJ+yH9RlmjKF
d0qq8wuWYaoZg4iROHPJ7efiYRYaCE700PNHQbIPYtMfJ2TPlrvUHKqtkiDnsw/P
D/ROwpwjiNVsF+8r+Rl1oaOV1WttWiyr2WQXeFjfAnE1IiMstlqR574Q77EQ3UBX
UWfiwVUzitDI8unmnU9aeTRoxEt+QlGF+l74/NiHDNa/DOPrXcNq2q6c6kchI6DZ
NjD4YPJb46vwaVNCrSKskRCEVqSfT9BHizLB/naoqAembaF/Xv2D5D/1SPqLvm3U
vkph+OCecgxcnEQ2GGOsKNlPTZsAbCkreHcgJbVvDTF2hZ1YBZWk+8Gg7SfFuVad
zgDQEZ8Ztq4AF6HTByki0wbB0ccvUhbQ8wnukNdBnFr3fEFwLjuP9u3v6XmjanoU
Z3rds5gBVIV+4B1KytVc9nE+55KqGI8WNNnWNP6+R1Kx+Qk/SAnYO7Fv099n3gOG
ze1ndAJBE1MDqTTHVTlDNpl7C9+QEoA7iCharNTsJkiQmRv6lMZmWm+5k7YL10oY
6GBMkQev8RzsPf3ddRtLoxiZb1s4RIC5M9+ScM2I6h7YgJ1Nl7eqaf/Ew8a16Fyi
bNDjy5+k3Ubc3yOUspsxRg/XeRfrgS4OcEeyCC+Uza7hBmzedk9jp54/fSip9h56
oLpAIHW7P0TUc0o+rceZAGuNXawcOM45eKdJydnsqc01k/JdCDY+hhIPTZr5sNWQ
B3fTDx9nSZq/0aWkPLMUqiTU/78x+0jmfO54Oz9sxGoGvBEVNaCy/8X7woTXbPcx
hYw38AnyqZOTyiwXDm0sBJbt2zrfgDVHsNuvec88zHijqQIkK3/NHutvwDWU5q7C
82mMUW2W7T/zsbTI7LMDShsO+tG52ugE6EXIM945Nt1p9USsQwc4mwgJVZGiaDkE
ZaAXw1kn0H1WoEFbUm+VJXXrCRk8wPRTTr9Ry4gD+F8SPRVH4MCWwXiTV2iz1Xrg
yQPJqX436bN4PgZ8XIO4C8u1cfdLt+QrVhqtXZIU8QgboOOaJcHVzwloQz5b7Ce6
cJZnr55x6mWRr4T1AYiMOc8cwefAh4a/NIP7mPNiu4spgHf9eWQH9zGhE45ZkUx6
dbypIoMSscr1hitWQLs3sRlYvNkNIP2YFfecgAFzt92Kk846QsEJKBpr2JHRa9mT
poCRsoggLN/fhjFMsVA/f8twpMpUywso/moUdnAi7705grH0KNsd9GE6w4Aqf/Q1
HbHyiS8Lzf08h1eHAWwWZUpbPvt2pkhuigQB27v/CaqAMqVord57fUjqqtyEcR8I
cWWrHmVYGKg/FSruf/XQ71VUmtpeu55IZr3gsUV3SPz6R9N3CF7KisR+1TSIgq9H
FBuCr2BAComMGPkVxIsuCrZ0V0tF+eExkUNMoFdlBXSoG9pI9mwurGlu+onaX6lX
KaCR+OIFFYb/h7vA+zsfdjVSSoYmmpmX2vc2lnoTX6RQDWyxqp8nkZaCsANp1bqd
FIpLjXhpn5VoWnJtCm9DyLyX7JTCuWMJGRSqvepdRyZCbjChQISfyWfBymMDeDKI
2CCFYz6b3jWd8z5MHbwTK3Dw284a5f/6k/ykOldYqVcvrK84fXpJ9xxb0mwgpm8Z
URyPKYbTiLwmvnDxYBuVMn0f66TW+8M2TokV7jlEoRbIVnq+r7gt2Baor0lY4Wuj
AECTZsNGmKDZN1sVmsKhxf5M9NliurSIQBgEes6RKxDFYF0uidvcXOm0vfERYx3Z
JBps2NreRu778x/h/3Y4o6fZ5fBueUC3Wl31E+erLofprUEC0d7yiThWchddFaoL
KgIN6/+2CpRj4Adq3SyNTze6qXt0jJaYMl6PwCksmCJVkg1QrYNU4KvFvMpNtxdY
ShNNyL0O8KAWCBHnQxW0ImVaFQL44M6XuXwicw9igUEeJC65HyYqeZTWIf5qyb1V
iNE5kj0Ql+ODoO8rssO5PrCEF1N9yoZ7eQl4zPKDlijnK/NZJt9DTA+Qrf3tV7hG
AW6qEB5cEl37oyCDeGjDuofYlLb2zUGWIVGfRTX2SAZLaUjxnHfJaKBzM5Sw2Jdn
T827lLbO7iJeDZ1dEZppEU14o+0vKnK4NE/Q5dCqNUhIosDpanpjwZrEA7E5FOlM
rfgUJ6Om9iRWWWQnmrgIcejxhNI71fWiOwcM7J7kqEHO0SSxqUV0ln+3/Ju9B49N
Rv0O1nAGQHDFRu+D/gXTlMLkSs3ou2fMG96EUyJFk+ksaBtpuaJpWLVl2sqAWQ6L
QodDIcw9kkPTmzFYDC0opHpnAVccqmLfQdN1fNQc11If/yb2IIfasO+wqDrswp8x
3CR3suDnRcrOrO3CovnDITxJ0xQqrOgyLar+VKWyMy+05tlWHL133Y9Y6FqBf0is
LCyCq2K47QXdta6kaCyRI3Egzjb6l9Efagdn8ccgndZoGHzMOu7YHSEhQZtSHVZZ
5V/M28vGIv3z1yhH76QC+x/6ejCVV3GqLYX7xDmgW9cenY1fKOnUizThTh7zKhPx
9gQNhPxzJUl2EqXAmCeFIWGHJMBl6IoG7r3GLKNm57my5i6fV/jdEkrpHOtJEqke
0uLEIYzFWbxY4x4uRX+cMev26ftQBn7RgpE8hJK2JXBvfRcnL/eZdDKcGok3Eaxf
ubp8Gt+AqR+jkTAT3UYva/Ar76SJMgKzOXoVk+vnLZsfyVotC0c9QGQ3vBjVqQ/P
aB0wFHBYgMSAbMC+sxB00yEgNwE1sFsybufibSviY4u14rPFC3BhtQQsCmfC2JVi
x1kaKwMF1op1knqfEG0zGQoomuy6sf6Ah0dNJ6j8SW0zssJGr9szqZW6ke7K1Q+O
LvxxBbLb8CQhwRtIpLQsvVp+cotGLgQE80TfnHv7wmaQVTDZYkeMFZcvyZJ1sN6m
1oWVqfcs1hyee+9YJJ7yOayzrHhtfV833UKuXIiJH/13YjsPUp5Qj2tc+zDPSzcR
PH5pLcmlc4P+HSBk4I8btgB2pXv1FwP5Fg5n92PQ3LNfgyKCLlWJ6n6DlxcLHZ8k
RMZ0vwTXmXU3oALsN8PV08MYtCcLJwOPHkiX8reVxOvGFzkJigF4l48om6mgnctC
CiA2MammMe1hKX/dakFM+R2qp3u6gMiAhCJ1kxyip1j5BJS08/VooKsL8ULSSkXh
J4U0zwQF7fb+hjUfpxD4mcA6WYN81/Fcp3CoN59ggFc1SrxrZkPCtGqk+m1q6Ter
1j7ufuX0LDNy4FfI4SiAK5pAcPECvq56mEIppOLkRKjQNarCgekptbfu81rB7hQE
uTm6fO2cnSeElzaWuyZtIU1UiRTdwbqXIe5Ltitsw93uZyukriHwcqZDQ/Zv0z1C
XrVCO0robvCIXm4b6bPDUkocb1SHCvWR9xA8EG12pVlQ99r1OqVcfO0+V3XH2b8g
NUCnnwPkOSW/OiZpVUwC+1ZcuttQxOeyjhKo35U5peecjDIIhLNh2A1beKASsTdk
AcCeNnVsAkfWtiMuBmx3u7st4zw0JUYh4RAeRSfSCCOa2dwoyCjW9Wc4J6Iy/fmh
pyqBBrnnEYS+a6u0qQfGvDrJMDv9U73GWykOmHCLgnVTIdBD8oEAch33sXEFVFai
IP8sCmbgsV4wdC9AQoFoDMf6clUhGs4pMBRoLui+3UbKka3xvgbMKZe4nv+aPJzr
Abn0CCCX+Y4ff6eXNp3OR24cq/EpVoym0crh0wRGUHg0WJuKsTeKXLh89638fj9h
gHHPJ5DidmcW15S1aWYmF3ATLK33JM1Ua6tRBYWtwhSKty7OahHfoa91FBfQ4Qff
nZhnHhIWOE4UYQhF2Q4CuVO+WV8MhUTEHYF38cdaGrfZiSb+ki/VWMJcdj0uFDEv
dowbfjgv8tnVqA9IWXW8hwZlCyLbLPIS8rglEyij+AI662XxP3FTrtAqRZ13z8GH
wqMsxiwx47yOxfVGYR5IkcBf1E6R6HTF0BaTnzYyLsBtFBJ0XL8lnMsrpiCalF+s
PkgCczzacH0yhFECRJ/eIWgtKreKsCzmQW4Eb/nk8hLP2lD7U1HWfI/vtUAtPRjq
vG4KcxKX/dolWHskxgr8CP3Bzj0zUSLRmYn/+awEoM8UeWgLCr8lB/RJPvM44dZR
dDdxemePzOeAWtRv272Was9FI5APjX/y2NPO/Lw15cLzvrat95zRxp2Uehyf83i0
RpZlcTeEUxIVBAXfw3BP24J6kMJgqSl1qEoskI5WAxilKSZRlHVS7byYKkTA8LYQ
5fDTBt/NkvFfHuUEp7eDI8OTw6EIIbCMEm+4GxmwfssbW63yWii+lQIHqpyoIcMg
/22a8FKpXpk4ECjezCthLXTGNDFPmrnhrsE4tR77UIO4PZdqUeXlr81zoxCUs8zQ
eYldXBjS7Hl/UFQJ+fhNSDxaIBD6e4+Nhp+QHrxJV1yZbnxX+Zk+bGVg6M6LIWDT
aajem7PA0tvdG8RrW77LOvAEo6pc7+++2pYAQ6ocOBs7pGSpihMX+m9FdmbaACvM
E0CFw95o1PbMBGmCdJhfe4uKfPjuJiGPW2gnxkGIpayF1Y+o9nlbNU2aF4heJdLD
QaGuoY9TggAb5s+RNtQuO37HcgPEM5RViOEo9CBkv79I/QHpeDBKLic505q+t+FI
G9oEvNwrrgUTtVPJolQvgRhvyaDjwzaayDX+sp+tfuahYH/QRxz9oVcPDCl5x202
G6pcOPOiGZSLy9aJ7lj7maePKxEFAV88f+uMRA4YFvhtKzlGyNIDaY0LnSRCAzYt
2Mo96/wbicIqUMU+3Znu7ubVzwK6LHDPgYRRWutQI8ObMXrkNthf7ZVRhUytAsHO
AemQ0VZ/DILihIaj8Vbrt8cF71swPk025p+Zh/J50vcE7P0WmXwb1L40xkMJExY6
Y9KQ7455CXSRADCPr/vytGiofOGXH8sIRPT7qvpAPaMGCCyZxPX2pF9KguYXBbBh
yb63MB0ALa/18OG7NSFG72QIjxfq7cKcGZMMmgRteiwVuhj3EW+7Fe43J3imo/Pt
qYQcEa8qZ0vnpsDTx8ADLUDV1ZJfn0XCeI3HQKPaVOc2Qu1GQADPWqLWXwqKDVPl
zw8oTkry+YnGL8Z4QFLF79UDeoo5/hYg+wjDs0hdCM1y1LmBKDjq4E2aPacRrjlr
dRXkPmVaHtB4khQtta4Aqk8s2ItdviiWFwJGQAgo58WS1B93ShtBA2J/RHhx7Qhb
u6HgveFlcadgY+c8QzNyAiaO+cM7+2e08Piz3lBj8/8jmUxQhaS2pCg+51aJ5GyX
70zhR8QBOSKteO+YuQ7eWTq5Ey1lJ+2eDTY4S5Sz9lxqeGzn5mdWO2Z4J6/xV5+H
iN7JgJC90CTXPn710v9AFpXtggm7loXdWQiBFWmpp6lSW8ug2vZUEZYXUGqsCIjx
BLudSIQt8qrRdkkQVF+4/E3sDPIvkC0JB9UMTbNFKqYX43GAuhEzBNAtoKI7DdTP
PmQzVF65sp6FB8m2OZNI8D1QLx9Z9Aj0l4y3WkkszMNTSnYwoNBn2oHkRzN8np6N
H7b/LP9s4vD/sKCgaj1TzhUU69gMuFfOLhJqU28sHXTRVhRB0nflBTvoh4+olT/Y
Mnjz/FcSkt2yFxzwr9l062jW9y9g6TkSp1yqfmHuoSlKb+Bp2NHzJU9E42SKB4S3
hSe3rXO1yfsh6MRxItzISY2HXkNPzJPrMoVukQO5kNgtm9MlgZrYNKqI5/bbg1NV
3FELk7xx8uMy7t+zbghBAczP92a3qRc+ENYhNJAMy7zxAnPzxVcWttXz94Ye9cxO
Dio8rZEvC1AbKBm3fQHLIR895XTgESpkZ0b/J7RJuT/ztZDxy/8pTb1PCYLyy7I9
VwUIdVkJ39vvsX37WuOdI2oRmQmjkHLTdBgFOT9ZuHf/N3BS2VQwmZ4gVgaH+9Iv
Ui/GUHHd5elHh1tsVj4flksvRANojMwOU9l4cKBe+5VtggNv+7vdN9oQURiM/9vP
ZCs7I0Nwb7s42UMvQCPCQqMREcfn6niWFLqAa911DZ0bFATM2881hUtpnsh4vK6/
+9VuP4lwBKJonTaHFKF9mnM9vXWyD+Xo/aH+zhH54o20mKiLNN9aH+PV7iiMT6Eh
JozkXQW5wTIfWUAr2YzWh6jC5qGQvGnTBPhlo993bVuvAOSJHjSZv5Dp2RoVaIzF
ORe3n/S/eIo6wglX+1HBWoHHESEXo/DTSiaBrXsiHIgt305uDfOtG8OVPdc+AzWJ
3nZNdjt2FgJ6HUvYy4ZuHyQ4MjUwVYC7in6Z0GkiDq2EeeCTY163hyTscfXW9esT
viuvgk/EnAiISGhrO+g7WWbvuzt++ddqYVS9avb1RmriiybYt6v5g7kZr0B4KKer
Qo9zlE+SOt8Oeh03Xy0uZ1BdPaUOgyyXd+/K1Njr7N3UFmCgRdl5adgS/EmeTXF1
mTjrKRI5WZgs3kveSjACGHMbWwED5508Vc9Wkei3QqDa0qHaZSgUW3hOgSp6PbDI
wM9LhusWv8rtdaKn92VUhuvSFJ39f6o5EY3VDGbV17bd1xMjJYS0AJEUvlSDqNFl
w/cLVysfk+hADDEYUpnubyx6vr7kEpOfHu94laZPgllLlF8bN9YpdD2P2u1I/+jB
9Jj4NEwr4UbGlbKKELoidlA1nYcqE8jv4PHBl+3JAmb8UkOMHBq5+aZBLFwPe+1L
nenBMfdjgHEwhVaW9CV77AqRQq3++rq9mz13p40lis9gN1e4rD3Ce1iXoU2KkICc
iCZRd4ukA0SiJil72HWNXKcKHmwnVfUaPbCcqZkeQ10D3QJqgUuPra4kmXOBkLDP
0D9N/SB/RuxWaQSsCNuhtqkLLZ28OeknMPX7qa5Psxm6vOEWfqq3ewM1HmqSTD2a
g5EEbbh/KmojTfcCRjgRgjWnjA1zyjK/UZ41EF6SUyIw6i2e0enz3MWKlbYEgCpQ
gsrHYTYr7yHiHiY8zsCjGmlGdCnH3Y/sI8ui1xDOo7ITV73ppDbVRyGRLqnwz9Ji
bZ73oGgQP3afAI/pKGtoAeRfOawpG0XKr3vxPaTGmh236gWxRl6XlRl/ZkJcbBhx
bwfIRDv5XPAAkuPhjAWB0JVVaNlAw7Lg+er2IeqFCotlgMMbTz9qQH+YDTfjKNE6
B5UlMNLuEce3raVWitYdMrGjeKIGYlgA6PLN/nEawB8vGcrecUE3x4nOU++Dk/Ka
uEjMpgtnvlogsEK1nnXKMdvDxC0o98K2ELZLhXlx68k0VcXHxIFh+pNPdxj/uT7b
aABhF96NB/Wey7KgcdFqDJjTidrZLwbdGBjyRbvq+4GM+5bYIOMfDO0E1IbUd/B7
OUgQgnHKjb2XsiWrOLStsvdHDVdWg8Ntya9KgpkH8YGPQcO5MQGzX6qJ+7YK+2z0
GAnuXhC4ttL6MzympL3FtPtmMEFME50sY65F6MiigIuBHX2WeOeavq0sQhBrODTl
sSjNTMPzkfpZPcL9iUGxRi3ir0U+DZ7pHxoUmsexA2FAj1R8oolw5BaCIrjEfxNr
Ly+xEe1TfegejXQ3Hlms9pOT4HeRO8RerARe52RaGwj6Xod9ZRVRbahT2onCJjci
poSWuN7l711bLZfAxCtHU/LWXJf4C8K20x/iT/J4N19tppDoiQjrSjgCEM0Svp2z
SqEawvZTQYFBlm2eD9ohqrtsizxIVLb69Bt7wokSZ6bi+Y30Wakha4E1BynuKe/C
LitJvWMG/9ue2heHeAZTvWsVMIbQ5peal7ocQiWCOkcJq9LJyledC5bqWZN36oOS
2izE+zxW8oVJA7EtkbND9Sz9r3yxIr3ARhmup3GWSOAXQllXA1CffCtisFYE8mi+
az+prwEGuySFrJGnaG3l0oKTFvPnFzXXTkAZe8j+rvsQnXpz2DeBfgkQysMKe0Uo
KIjMi+56e5I2rDInlXIgO9c1YpO7zXd3ndUFuLjWlCm5x3IFIhAJhgs+LfHZZqmM
Nqa/AMCiqjEoEHGiJRebvtTwjD+6/ZvrWrZs+olzZRN4EbE31WBw7HNnF0QxzXLK
nUnvnHWiSm67G33uOLrZkbuUwFGHuOC11P9L9Ns+0q8UDn7R1nVguFgrbQTjnmSE
g4JRir6jKV5RjSFmRVakHjreN8WMDiz1tf/+7r2iHPFoYYq8RzTb2bM6UhPNcJMd
w0ufv124NBL5hFPWh5er3Bb5bglNm2ppMFXJZW75ULSYu6qW5aejL79wYCBFZMhb
1E/v6emdzBkcV9J9tG0c7ZaXyVzIgHu/zn4iQptpxeg6X/yxFhNtx66qRksGKVxt
EvuAamRPAehLz0KBpBF11+ta0w2tDzx9I2boVHFczPhAnuvq8b8g9gLfBPIP9cZO
CXjYyrvMQ0m9uI+HCflhxzRTSyo27q9nHs57igiNn0PCJ4hETOWxrhnUuYf46Y+K
2SkcAYGisuQPUM9h/5nMjoxQIkQTgNu1nnL5enPb8Jof7jxLQZFUBrRL6IeeoLqE
Iz1u17C2YTuGOASvNCNIJ15Js3C50D9MXH8JDFegZ8oGv3nD+7m12dVXaUElE8pC
ZcTaF8NYGWIG2/1jzR4JvEG+3J+l//WGh8Vws/kjXR7z9iySbzvTnPBHIr8Z4ZQR
I83z1j9hMJxJohMtvhq5qreVScVtl5T7cw0mALejA7JCfFK1q2JFIYw0p541Ll19
TBHabN1k+05Rn2ZCxGq4baz+R93YuyR/2CTaCqeB2xipewmyLswz5ABafinEaper
fqPdfpInLTltiatxEo2RN151RI3MD0iLw+ThgWvyfm2hGjvKX6GlQnE5DOdNQi8M
ZWDpY0zejdSqLmci6GjrttCG9zSzP32BZ+NDCNNiBbFEWE1Ykx2Tnl8NSIZMMnHR
Sc48J92RxHG8mg74RDtiFnUZEl4lABh4vJ5xmfFbHBFUwMTmAM8FjFiUMALddjtP
HUWPcwyiaFf80UhgUI/dzB/GaTckqrIv0E6LyRQu7VvD7L/JYdEC16CSTPgFAYu8
mJFtRTiqVTw6dciJLX9REq430f2s1AelNbfTrzjvDskoMdrvo2kMNmrRcOhUs9Je
fdEYzpE2QC3bf/15xnE4IGujtYbn/kvdxqPGwocPmAKGiGQrCF5ox16rbXTMI/Ny
51TerFMCuEJlmfNdRjcfKyrp/X6WCoft3s3woXUErozQ3bwSF/3RCpbgGq/JhhlW
HGvekQKKoAAAFeM8tBgXdNSQzktJARqVtY2rJy4Isu0ANu+285dqPT7Kn1woS7kj
R8kig6Hmugg5lBmN3NlVv3d6knfrA4x1eTTYbpJBUSPEr7cDdYYKBOIfqwhDWBQX
DA+W5Qb13ga61vKXYAu20gFOSOr4xcafQXmUrB2ampAaSBlcfQofOSYmF7LNoBUR
kchgeTyK75UPVYVE1OAhnlScHN4n7xklJUjwG8sEBdUz69BVD/mYl6w2P/3+gKok
U0SGiVyWipMdTK+cXMK+dImUY/gI5hYXUboZfzySTneMZWQukIoMPA98kiktNBR1
ZHxx/mKTykQ1BKTZKBez5ohaQIYrlWnR3J6l6qhjB9hwZsvzuakB/PtpYLPDauv/
9r29EU2qUel8u/cRJoLRJYP4Q96yhOkHViZA/smoiO4ZhgRQ/At1GX+N6ODXbfp1
i2Ady2WlgENRl5XC5LCMGu29i3/Wk5WLF+NYDRfXvNqk9A39GnjjpSDrAscpBJD3
FU6umVJd7X3L2szeXMsN988I15YmKMesZgQvj1C5YsjB4c1pFVMIv36IMzi9MP7Y
71er/8xe7dOXtNKDju6y62QRJKEdigaZAjS+7CCdTkT4/EeiobnZhJqWCxlB9H5W
j0jpjVR8Kc6S7xkj/D93/dEZK/e3lwraH3XjAPi3ptldOdL1SZP6mwtqhO9s7OJ5
ycYdAVJP2kiTaESXiL2Hjcb/vZNNoGsTsXju9Y4Zy0VYWxvqkf7DfwTvXyIQV5Cc
17qHzIbjPFNLqYsFmXX28XOo/Fy/oTUNDvObx6CXKtbF7ZNYT9zb3Cr2qOHAMR41
nvjxHwG8IoyT77C9Z7GcdVfqDcSDYjsq6pVOKwCnEA8tfAkKJm2gwuhuMZj54KVg
VXKwI9SP4/SRZRx0o1AASs+4Z/urXyhz3xRl7Q3nvwShHzj+DVgvNOL963fkSqVS
MEmWd6I4IjHpBtSC/yPwctH3dwEBnpVGUn+Y+qIJLo42sRC35T3RjSIxShd5Cfdw
ULotBqcoAAeBITbvHKEaChbagBOaBbzoOJJLUUSKB5efUz0j65Tfyy2piVJXUo0Y
R/60dXfVqWmdDEZBj5ItxZ9Uz9A2rmsORsCUs/txBPcWqGKmQGHJQwbbzUygiZgv
S2nIU/O/GNiaWxaonkgd4ncJ308diZvTgx03MvKbZiCdF230IL+/EdZC654xxvJE
OajrRA8ACFV7qQewdlq/VayzJ2usW09UIPF10cvYxCRnhdm3rCLjO0AvEPVch2Gg
Pm77mBvnMgbmV3s5Y2P/FPvg1nbgYvXjviIxTyEUtTZbtHMAYX3oOoXbvqAltXoQ
lM+DuyWp9Du9lYvyUhmitYML6JCRKIw8axx++bzii+RZKRJW4KSjnZq+UdgVXDRH
9M0l5u5cN8Qs0MN83vDUYA61qhp2C5uQbqo+hKIxQ+rvnPDrjPmxPjEHKzdPh96Z
kmL5feKbTGi3gpdIi6/4DrjUGI3KIxqpxgNUpCmROqq52suvDj1BUmZXMn5UXQoY
5ASL0oSzNsuDUU07zao09NTdbBTAhefOGeRvLaZ3r3+zI/2k3RKrE1D9nvosTcj5
E5S1ahTz4p2p/DBc+D5xah+l/kyxvud/VpKwvFsr9+Cy5ezd+gLGone+tcsvN9eo
I0po79WMDOdLG8sjBVsfWXnU31cadVSZWhTSK9LhlA7UKoJGbXxIz01KFmyaTHR7
Y36lrP1BulYMNvLnofqSB4xw89tj8DVcjfUkM1uOuqJ8go7NZ/tolReTSpPAF8Z2
BYBBCqT8De0pcdEmXU/LsLkLQk/mS+rsLYPlHxEjNztb1ZAfMeUFh+1clfRbJVCh
zbksQvY1EHyALsEEDp4AMErLcvuCK8abxeEyRs8slPExGd8ZLEVbL3eidx8jHz19
Jdv81FeMKrbmRQGUJLpcsW3YqKcpYfjgfteNJCQF3GL8ld3bYY45LXDmq+blZ+Wx
oUHIbOEk9gVOuRWVbbQf+IPCNUe+M1HNUmghA0WU+fEptmgUcda3lAXb9p3OK6WX
vb+Umd/3oZv/+dHhAR2VgYepKxdPwXFDs5VROwTMfKlROvF0Nd+GW8iRxOf8kodo
kOOg7qkhZo377KbmhXMUaYdmC78fb5jWmpAXfZgwJU4g7KolQPBN4SiFLqwzrkW8
SmdvCEw4DCxTuNDEkB8OelbyWuS57UXHMFp+nYJ1NC6MQHALGSXPAs9UhcBnESpQ
Gj4sGCfePte5BwsudDL0q05S3uXO/HDYrYyNQJ26z12gkPEcFsVv4L/IjMN3/Ddh
yfEVrjjtLe+kC8UP7LEvU7WC7SlVSh3b/qFFG31kBBiyqtENe6/0VQzcZV/txV65
622qPe6DaiF6V5RRuPGeszi9tIJf9bEyxV4m+WY8kLbCwlUkuFeRvMlzFnQiDSGt
mWPwL2rWqy/ptedRldvzmI5v93Ekmd11f/hLGCO+MpvOVxxWITOSCHK3ArYZayKr
Er6O9me6YTXkkeF4H0rG6BW1NocGia+LPlh+T+l3X8rEaS4830rAHXPIOZcdhu91
R2lgYqbIylqaZ8ZGKhl4LSeylHvzYB7BPk8V93f4HMW311FRzPWzUR3FqcT9cKCn
If5wT8tx7zIB7OyEWwYEwpQxckNao8UQeZXnZpkHGlBBGFBHzZYyABfjj4HDaOiO
//jtGQw47jGw6sNT7uXB1jB5//kju31Xk1U6tE2wro+jatn1ArBxIip3nBq8lz/5
oktccR30/LBTSWqKuaHeVVHpvJFEU4XuRBggW3kN5acgcwzAtpL3nxeTC8RwIPUV
noO2WMcov8/pdEEOUdw1aUo8OT1j9wt2Pe7gdxCQWUZp0PG9xh15kKNUrOYwR6m+
5ex72XEWCWDAFE/EQg1j5UR5GzeK+8wEE+HJIALl91IIIKmNud8ksEWAlWzg3YFg
JL+pSJ9+AKwKgE8UoyYwwyCCRwhUCoV7bM2AEDaJVb1y3nuupyZlBhjyQ55j1drK
5kUjK2PI3C2EnoLRE4S92PLyn9IwO4v1Zesf4mloHHGte9k9rsnbYSFhy0tniXXP
WbmxE92Zcab+H1egrO3b9x569M430W/3Q+TI6xfq1YIR0wz7vG+77Ku4EKVpDbO7
JG5FUV8Mr60HuYPHEtdPBY0tBPOKpWrhs7pmwawCkM5iK3kYXjU0JthsUHtKZdmk
fEshKMYRAQAqYc+n1zX1Jty+FZf5ose+Ty3PPwaUVru2HSlIiwFkwd967COTNpuf
3Ss4OiNO+WVUkCZb7jga1QnD9PWt6B2c4D6weUVJayouFu6o+NOWCCfPQf8j3Pow
8N8G336qBqR49EDlwfF8r7MmlJYgBAqc06x6i91uRpd+yHZixyGwuKl303BuytS9
AC+ycAdwvCBoGnaxVfWIvLlZFCoaYw3pvPfazapiP4TzSYKhkCljyqTeV5YNYw2c
53E4zMmuBxKFa46n43ZpGuxW6sdtlTI5AxjnpC3j/kfOOPeod0nzodZ/Rusu5B5e
32Ae8Lm9NeNmBX/9cbbtZ8xXjdL+f4IrMQg/4Kt4qCfUZnetOqoTWKyvmnqmmThv
89QR1rcfmVCuucrsSG9pG/KU0P1SY4b28JGzsbo4Xh0n/OqmSS0dCPgnC3v8x6+C
x6xAbcbN8cjcXfDAaZXTntc2EXo0BkjWKRMjUSwAkipMBShbsxWRfGyT79+kBPsI
EdjGI7zlnjOFMQU8Ow53deZqGLI/cJN0yi71foncbA3vWFQ7SbKnG7nd+LU3qQXi
/oKfWfi9IRSJwZvF/7bvnLPZsa7cCsWkEdcrhDdXe21EuxYhGojDle0yCidEN9Ih
V0eUZn0pEjFYY/DXrYsTnYdagD/w0TdNRR1LDLYkIaUIVfkdy4/ekqa2DzsIzyDw
6d2wIdRMqFJY8LWRQWP2pK37noDk1B2I0ZXNR31DOqX5P5QTj5yq3NxmuyoHqMO4
yGoog1tDnd/Lti7zk5oerNx9DZOIuVMVJ1ILwj9YGv7nDIxTHa4mklOK+wY7e6JI
HUXvtwzRRU98kaYOjpS3CHYXKHkv8xgVEdz5AFXmrKvPugrKFYBbRaO9T9ROHRPq
qe+Ne3wsl9SOQ2sm2RJ4Hyp4pXdryQ64/D46o1IeDeRKogWCKBXTcNfjruI9xffa
bxlAKxR3bQBY0L7Eztizm+UKMd607VN2GPkFGVQANSiIgdbcTypl4OyQhiBQewPl
8i0/LNJaAHtRVMpgxRdCRc0y+gFDA6rDzAP3rLHpHmdSDC0bY/F/+VhHBQP5sUCC
+0/+jQQ3qQx1vTxN+xxDWODvQL7dt8JzfddIv962HYjpSY03y/dqsYX2UcZNAbop
GwkNXCpvzWdz5Cpk8fgguM77KzoV/+JfyZLOTgJNS5Y2vkGh0XjSi9senGN6mx1A
Nk2bnSa9iZy45mT0Za9eAOW3RVyhAKmjhyR6DSqGaGKY11a00cXOsEf9jenT0JTb
x/fVy7orY8L/Lpd+7Cfd+2Gnf94zs1kDKdfkHhyIT2ag2xLVcAzQktSjWjqzx0IJ
ptgZ62tvZ+61E441wxdligfKO8BZmDD7s8H7EYNJnn1XUr5DpvBZrJn7Xa4JQJdK
VwPRpMq28BdD/OYSk09Hl3ItMNGDZUZ9g2FSo7PYesCDeVHKO0ztQsGqyR1EIb40
V7xY5Y1vHze41uJqYBGV3WELvJ91QMOGpbXC74drpUNusyjjrBzOwm5XhMgJjkR5
neqAhtBHGXyObddWctpwNypOImvItciJhHGH5WNTV0GXoA3Kf09fFDDMMQAA5lN9
kW54nfLPLLYpTNcWal/7tevnYIayZ+yeI2jOP0DKYF4VleAjQhPr3lRDmdy5se7V
TQiVjbK4JAnd7Y7dDFWYWpRIFARrEN62IuHeUNiiq89qdRwh6MczFEjn2E16J+R7
cfZUiOMP85xQdtdG4yUdBKP1Rvrm4hwg/zUr/xbUy5jFF4aSJNPEcX1g6ZtKiv55
uCf0fcEFeNFujICDdVOLOWrdQNREs15OjdHuAnrEuP9Nr2OUCrh8/xi5mJoc2YI6
kEDJzirebBnyCtQ4y3U9KvpvaWNAAhYXjgWTRJbOyPYj6dHyQ6I9kaXLfJpwsU//
uBJfHYWjsLBo461PhI8jFC9Jfc2kYS1Z5AiDAzdM7dtHqTWoqDatTf07wt4+X+LK
ObMYrDO56Gpe2WpfZracLrDJg1I+CuFBwhzwN4Xz5vW9JPj/Xj7n3hDlWI3JmVA2
r4Z9bqdhJLkWh0IhN1/SmjyZyw5cxKUanVdx4ADOViCLmDciLfOuCEKf3kP1mws8
ZfJFbHfAMfoBn6NawKX5sBp1er3Uft8Pjco3c5E8Z8OtWVxQ+23ivGvxY6eQiCCE
pWveW+mbkkFx8pt4fk9ebvmaqSJ6lhj+/ec8yd8vINA7RhPC2C2sFXn5aHjJlAwX
Vc5dXUO7GrDK1atqi2viQsYkQ4qwmF0ECyLenTJuAV+UiEpAUeGtRInL/WUxFjAW
mGQsKUJfupgnkOmbKBHjwUs66v+nwWZoUukK5ZdlHlw/N/gZ2INE9JT5RROFtkFN
3zEDeqNxVt2nQ9KBeq/5U1tqFuebNzdsfDtadyRJRC0xLAqU8wl2UKpFb/E+emad
dxulFOLWGEGdceRC3XAvzOoO/0oMIJWuWvmRrbSCU8t1/WG/QyFWJt3o6kYoPAGw
z92n2vG7jAhYmHk0qG2pXS5+ea4RjnIKBkYLVzhLFgmbxI5D8Jg54IDiaW59saa1
d/fzjP7js6ZkvBnbO0W6yAGS4NqHMP2yDsvt+fbyVg2vPdfIXjPTLH2qXaFipoyz
f+bYAfHjxzgMyqWt4NB9EY7vVrcfgBQAt6PHnGpTXm8CRKHeEv/K/4jYVhWRMfyA
98XfAe5Z658kVTUmASjQ1ZBbxy87JQd/sGEpg7J3dkD2i+nRrdC8VH+ATauQ29Ha
QP4d881rlLD9Is8EDpuOcFEq3/AS2ksh9SH28Q9jf8QuYSAlEWSaeDkTBwf+o41w
DyPm4IuLzKoSaPgtzag6+MtK57Gq376/1Q6sSdjsGbKfz9kOh9FXJhA1YOOz2QmB
WuBdLTyCt44o7h7w/4Q8AiADDyzlhsQNkiLRZaqCeGXj36wMeyWkHGycrcCG0lEJ
sAHpADhlXlgtlx90NxPSXFSFgK7/bjk/LDmMDtbN2pAA3yehOm9fsRN1bgTp0whK
0tSdPkSA2ey2coseF+HRPHAm9i75/v/sqlTO87SoIcgWDlH2NpiAIW4rYmOYMH+f
sK5nzYKN0D1/hqkn+JTrGm6364+PgIzw2QHetIGmS0+fszzdbMKzxMKDrnr2oXVr
xCRHxMoEqUdh0PB2jIm5UyRqySWM5c9jUm/XyfK4GVtJbesVYDtGZ0V8Zs/1LBPU
BwF/uDVk0awABt8I3Pv+WfaDgcujYrC311WyUEPR9ulzGl1/3pTnVfRBGRSdd9U8
vbWFT4vOV4QdExVpjRrtf+ZfnK7QcIqT0z+M5njFd8D/YOZQAvPl+Em5+VM0itdv
XFN2elPdqsE0aKMs7ke/MMc8qmWgGktFu+qdmTAsHZ9YAVyp7uVpgCkOE79/3N8N
PbEwRwjZJniTG0NRN81AqkJku6HWge/a8nAp5J/WxINWkRo9Q0qMku6fdoiDIDFs
hJaXiThrQFLC4pxsH71pNmVcg3ddEcHPSA2y8DTp+TvGKIOqW5ga4biCBSrsUkk0
vy1vvReY9eeLsW9NRTOvxbnKjKoHUEeBZZcOhnXQlahihnn4ghfrxBTNNq8zNPOk
qXQjMikM53XIJRlxOe7e4CAq307HY6y/INJOxxV9poR1/Tu2HlgBucaPvkinkEyV
sNKUTzZcvX/zEblsjInH0T6q9og3k+a0oGwNHMkmt/esBz+oY6c+/cNztoBA6W5P
MyVk+x8DboW+eCyKhkNz69UGc1ljBj3uG0fOaSyTIOuytL2IGIu5JV59gB6L1lwE
n+g9SxGP/apgtBHgjwqptvh557zt3uVrLWqgLoR3mjoKuq1JDBhXmgfuQZRYEsT+
DZJxjN2U/iC358ouBDGAZ9tFzFAiHr1ggzWMD1lmSCPtzNQP/SIQNZ7JXSl09p7m
or+jIh3aOe6JdF/JJnkfSWpCyyz/4cFxbDhlU12/6m8/KcnSGBVMCUUZSJwsyiAY
j8T0voD9Ni8U+1gu/zMxx6ZJkDfb98wfHh9tEnr+CR0yFr8TRtoqaydsEj0WsrjJ
FNVGHX4a37XzeUb8De/xHqKwWc1zQufUu34sn/024EqT4+3BIYGVectPHhfpQEPZ
eHaFDWVCOCdvEcVNIMp9LrEUgYdBeE1Q3EiGHQNZOu/Lb7Q9bs5fVXKFW3v17ILw
KrqtVO3PMYC1i0D7dAN02W9izqLfq6xp+Go+o9DEhbCs627Fs9PRxeQlCn6mWOvT
KIMxwFgQ4LrHmL6a08OqtQmfXAW53mruTGzDFYwNjh8xZH4vSxI/kRBfZhNjLgPY
oSXrgRH9m1PDlezZCQ58LulRIVYtIp7VIT+P2NK+1LjCbq/DBfGlqzQItzpYKZRI
PttEUWbWJNWVwd9PUP9ds8rP/RIMiFMtQg6vVoj0sgJKFDLayIImHESzXtV+vmgY
G3ZAv10IXd5Tq20dioXLRkIM1fRwpf+7nE8TucBNMgcxqzdJCHboFfI1+DH6PaTC
FsaetPUGwPtpu3HbyjihO9FeSzVaVsSMjCu/0CBOWSohOBjaHmr5NtYY80FYfGvs
rHmjSCTZXqaCwsUB3WgXJHh6iqLTiftrHN7BTFB+jJRg83DEhowzjIWT7SMemh0L
+G6YLec7gHzsNR9ulqjsrAqcm9ehhpIbwECxNCgLMRA97Y4Tja2vbK/X9z0WB02w
ml27Jqcvld423ZCNGr/f5ny/etIcNflvCTndet4z1BCNbHEga6YFCXY4tt574hv1
wnOgraPciqEO9yVwDOY8fXDyU/1wC9MlRR8Pyllx+UeC/98FEBRsovibVOELknlm
pnAyeSUQ+fmkT2WrhfacsndgSIBvoDklNwNR1VAywF8sDUpx2lkP0tkKNCY5Iz18
3ylqCTbPVbKFZt2NYRWvZtk31H8VRvhRKhZQ6LIKTeer36RD9xRJEtx6AI8juQQt
O8G6HJzGf0B7MYnsMOQI8Wdd6hH7zisltdUQUbwiaRUyTv3bZb0QfFQr843umSmA
om4itxu0YMMwMOYa11XFnWUfNFhMbDJkf2znjIHzsmXdGejfIjnr6Xs9dL3Aq+T4
MYW9rnaoFYRMmbwok6UH+bXQeEx1DVj5dzdg2OQo8ut+5gmI51iSvH2skWLMP6pl
V7JtmDN8VzK8PMgnAiIWk6Vw6/EQ9amf+vD5kgNLnXRDiBSGmUlj/2oWDNw6YvN+
5J4FYEQLR/jyZKgVCA4jWp+XnNu44CBc6ZIwQybcvmYOk3JmJaV269AExofXtVvJ
PdBXaEZ1s5Q0zlw97SlyHeLooNnAWgNM++fF3PVPKjVwlvAifHTL4mwf9RYQ9z3b
/uDj6oWr3OyykYymGba0igHrUxwpDpU4IDGUPZyWGEUhNSaUYx2TkXIhYowPYy5S
TJ8T/gq+/BBKTjgqM2PokvDiVLtAytVewPYJySLjxKrzFM+znTEhux4cfDQQtwyQ
2f3oKorEy3fVGc21kJ7DHVkyHrzp2/Ao2gcGzoi10x6717308KX1h4amaW+FZ4ZB
/KHtoV2offULHzm9s48xIr5lYzmFnTeAfz2Ab8gNytIzHTkPVSKF2GQ/CTvmf+bB
vkeV6wZ2En3G7R6MzcP6Td2XzEvKzaRToiE9xoundO8FEKhuB/BcZnA7TM7FLvBS
ardSaHueJg57RVLIs6D/U4g2wqfYilKgeeKP0KZq3FwtowzxquIgcqlPVdCDKt3g
tNkIrtGzHJgGozyor4um7pPUTEfOHL9X/5KKtwHV8JYN7vtGlTbpF9L5XI3F10hb
Tms7470cPT0phtT+C7nu/fEUOqsVVk8W+LD2riOqz0FA9AhzmzP+aOQfCCU+MO8L
s6p+t3RX734utXIrbVg6L8xff5I04ueF17tHG9UAW5Idk3ljbIZk5caXtwZa37r8
mhrD92M0VV5C4W/gVko41hEdRhsaaM7Bqq/x5p/Gc7KjsTxAayztPDDrvwPMO7Ga
dzOsi9/My8tbKIfk9qblTy/HasM90QDNaTOshxkdUBkxBmImkg0/m7HSLEnnrGZD
QRcTqfbqtmw9D07y+hSACYxAWhoW3wSGJy0EswUbSNOybUNlwBfMhwO1suDL1zc6
XaI39sImqE7MmHJUeuUBdkTWguahL8Dwxq+/BBTDmYbMpgKy8jWcCetnbA84PbeQ
LA/mLFtSM+KUSrgaULRBL6LtbY4Z1OXwKC3ro93eGVGQGmy9H2FOGQ8mVn1Ofpyb
LEMJEbRN5/JLS5oFvQteaXCW1foXBvIVV6WvGqcKRoyr7FNz/iQVJFK18BnFsbvz
exD0pNR+sIWfYWYaIFVAxc/5SD8yE7Mw0/tLHUccvJBKaCPqyYeJeSreSBDEMlhp
B5UuijP561f4cWMTc4ZiB6SOWgP9G2iqxVQhFErIN/zIM57UHBFjGg85+MPPSqvN
alhIB9/FfbuC3/ltHERzbTjVc35/VM37EaSnTkeIr+RJJMyeCVsLrjCtgad8R3Er
sa7qBx/ha2pck3Rv9E1eRdomx8prtntshuwHCEw1zEnTe9pw6yLGDmklYcTjjggs
QWL0I0l4gtl+c1urjqEoxUfN15co/tgYuL2OBgW4qVb3n4JQ7K2YDdUhAnAjgDB6
CcIf9Du7dpuMUBSlYfzaP//s1Ox114NvtBBV2/HKJRYwEbrYwfialEI/58nRKX4R
JP9/NGtJAICyet26Dup9axqmbQ8L22mMSwHZy7tPrQDJl7JGlgRMshbJZwqkbTGD
D9rwozrVIqi5iI7g56DVM7P2pPZTJ2S8NlID5QAgFPIT24StG8oJj29fbNybM1BZ
bktE28DJ7/dWq5h+8mhuXRTYhQPyVWYTp2bB7Jl1QH77g9P37RFK1RfQka0pmG1h
GXBhNp5b7T9A8LD8AxS+SwUtdoMY/3kKVJ6HsOg8rjn+OJOBIBZ5whbm09FMOhfj
70ygmAqc+l6cpQT75t5E6PIJIU075n59RTKSQdTVY6y0J0NeH276EijqKsa2RYoz
6QoUt0kG7Hczl1nA4mgFY3fE5bb4nm9ms/2Ki3oTlYd/SVPIJ9LD4hGrwrUq+tH4
5Lq345qRYYpDiwy7SjN9vi5emykgJwPWLKEyEofxPz9SCF08eztRFn8KtaP9kx7L
iHJIEuODg0CX8EQbqFRvhfplb83o7NWlHpg7ZIIJm9AYBJLYzQ6no7GLiI8Rf66w
6Ivk+5lKT+rNEs0y1aSm/7Nf7zX8oHcwoX6Isw1UvgAzI9TUrfUKJ+3qPVFNLX2v
rL0SPn3XNbGohQuj94Czj1ci5mVb47IWZg/IW3TvOxsRcNC6yLpdoZec+l2FFqxw
3q+gcnRMAKaLPOsrZaD0xkwvkbViiyUqu4wSSzQPpKZZPoyI+Yf2SbiDlKGlGdx1
iVHExovXZNBSvq32XmuSbVJKCCCDK3BgCcikSiDHuwTl3LPm7Or8OZv5nXb7Az9P
MG5qHAsZgBmv/8TKfTMGvI0Y++/hvOC5a/zTwrQO2o4NMQrQNYGVo2jgjDQ1rQZh
j7vS4BRc7xdv41bxD2Km7Sx3VanAmRjGqKsHLzD6Tp8ziQeNzgxQ9klI6tid3TtZ
C4tVkfOYZiSTE7Cg6e59hlhFKD5vvvmwJrvlysWIVovt8gImxXQyUjYvRMAPH2mS
RgjAndkpnvychoq0KLcDtQjEuyb3DmB/N01mdPoEbIVfGag/2cQmod37fg4b9AoU
DA9oO2m1eOv8xn0cWum/3TfFXaIA/qmxlscxSUGCfqmrerz4zzdBqrNxq6IYhuW/
6tZLHgcJqXBTL3ljWJhvizZnZZ8OK03On0Hh0F4Y55LFrqscIja7qpK8KWAYM3ey
TM7Fse4P+ktIY/Zq6A17Eafes2vNpUQ+PR9klcWMZCdjSchG7VRG/+bzDlWZJqU2
3GABCrGl7ujag8VInpP8qsVlhZM9EYtRJUrIAsnI8ZwJzFLkLcySPyyt3k2XymuC
XRfiY+h8SQAGtjOdUFqr2/xz2uEIMhbiw0hgFupuyRhyzHk9aXl0ik1aTHLR4f36
KUeaZFWgPC5IjL9EuS4NClxWT22WIkMgkCgCWtrSOAsMGebj5WEifb75+wpVEZf1
3oT0KC3f4fem2teM8yZkRA0qXLtgvZavuvODtdR4RnbBMZOPwjL//524+ms4fvda
eDcpNR0Jfby9f3ybCxeyeCr/cL9oZ+DtyYgbVha65OAK2QVWLGUe8z6NWQy+6M5X
betfPMp9VAhYTYBPCtkM/G4MIEEgES12pOBtUiqcsR+F82WFZUHGpY7PoJfUjGeD
I9qqOP4AdR0Ep7HMdAE0esN4LkHnMwoYvCxHrfcXGD7+TTl0sQdl9mXsS/6hbD13
nu92vBzIn5Pu9QLpgW3PU0vtJ/PGLVJgqpMGSDYX5ysA++xZThefT0C40mhH99RG
ZQL4VVX0ileOHIWEG/N6uU08hmQAN67xw6cnZU3UgjHvGZmm/io/AM1l+/vQvAwT
KyUxV6NpxbCAFHDpNNL2ahxalv1Y7zIPQgHY+AN5+PeJgeADCpOZs+ZiOFZMIbi1
U9POe89vmjAowPoDjsieICH2eZQeQIV33f/XcI3h8+xUlAzQPkJBUH/eHytouGR6
jpW8heM4eDmtXNPr4I2v3M82rOHKjV5EE8DOrKXUROhyAvu7GTnu4MSqUGcLFVCf
o5qOlAaNW+LD4lwYUyXB0YrJ2Tv2qcvBDHm1wS7Cbg1UBnkYWKxhNjNnJeEgGgSE
xg3dFJxKnxPP0op/CraT3O40SHbeHCwke8H9Gyt074qTe1e2dd2H5EfEJVBxkx0x
eJCPsNGbC9dGH1mNbszo9VpXkGSXvaDtzWQENNQnjl35bVfMO9CFv54EK5PFOg3/
2gdUSDMI6Im51ExVx4O1eV+1c3V9BWUboMY46v/UnLziRapSYEQ/74M+KLbJQJl5
WRdkTwBj2fJGxb3gAnHu5js5K1d1zv4xxxqgSqMg9HhNkQXoNVuBnRJx3GX1Csqb
ho42K7jGOj93yi/kvDxUI+T5FoNvdgNkK3EMzS06MZhwiZLeCHSgT8DwiVkrfUsJ
dfLxlaoWJDH0el9sDPefK3nF8LsSnu0Pw3NWSCs1cUcQINxY3ZLs7lfi7W/9JVDG
bBglsRmQnmzCOOdN0Xc+bNs232P7AKGjlSreQ1XkUv0XB6ApTJaNlVOCkpjbYVz9
PDmf8+nCo9uQ846sUNvH6Fd/jXHG+kSZiFL4VlJkzfak+lSauBtHXEnaGBkTqO3d
4PX6Grtz3T09RzyP5GcdVohBrNAprkB36W9KuVnfum+Gian1JGGqBp/D5dGj/btn
9cSX/SVXoKXhkZ13cUgB15GFTS41BLCBOdszdzHSVaWoXldmaAJmn+gKPEKEZx5t
wti6csWxgQ94he7QE7eQ8e8v2K5h4pUSA0v2LRyYzDQYynyZ8t7IpgzO94oLLzyo
zgaPCWYpgCGDIvVnFhIuc/07+NCh4T/oLYxMkCOwetkQ18K1I47YSvNGXafdRIKk
wri+eZ9AnDjTJu6kXOmXL/0nTtsB7N81PFZqMEu4juvzEjRcusu8TgDh61HTqW9F
CCP4MvCDB82JiULDCTFUrjKx1v+J69+Jp/296rbKJqQzCi/L4J07nlS2hbQQK3sK
3xpU4etPCOk9Wfd/St4T1w+0qAvmVxMJyAjYcevGLczhsof2zZtTiMUc6sUxj9y3
io4A3UEU0r8jdZ7pCHR2q9MfOJNKiy12DvuP6+XIHbghzDW9cZ7P+ZQNgu2s8dTY
0rX6KJFiL9od9z5EauLUo03m9wJ568F9oYj8n1vGXoZkj0A9mV9xWBFkeCVI/xg6
ZlSzNMM5GG6cOk8I58E9pLFDR0O1homCHGHp8jAuilkExUXsqpsQDdyktXPKl5dE
10yKFfJvHpQLH5bvvoTsdaGHI8xOx90Bi0pr/6Apw5SWDchZkrh9zeY72VkUKfBX
JUlmTBue224wlsJt62yfPvIDUHViRhIGSfIRBI8EirqWwc05eKa8sk8bldeoDEpi
bHG2lzQotZyoo0+w2FGxs76VwJ4dWqhHNZzlyEIUXJyrU3iQm606ttK5sxlcFe2m
5+97aA7VMAKqF15QE51e/aG61Jk0Q/vs2OHDR3RsAnHg1wzgQSmcy8ZisWqH8UAI
0T9ik4Ld+87KJI6ig//aiwDqOnBIAyVqSyBoZrPuUzcKb460pqYbT+Dinq6hun4G
XsM0X01uQNm1oTxzxP8uPBZW6dIte/9hgdP9o4Qadul/9Su8Dk88awztqNm0iL6t
ce6zuglIWLAX2HoWB3nU3N1voN9xg2vGlYF0kIXfYoLLepSTCJElEisyd/z8O3tV
hYTtbqHz+8RiYs13Q0GdzW1PYNuQGT75S077sV933J57suYJEIEmTh6uynkhQ2is
aOmIeamrg79lpIpEQPIGx+jLd3IH+OrOCfk/jpbPnIfjoYPeYQ+3BFfUGG9rzqwI
DlMbi0mi1eSYd84H9JPZ+PWJBW9hVQuX9XlX2pX65+5vf+vJIKjpdrrK6DDvonc/
hghZxbb8j28mJ/6itnn12rgqL6gH7yUboxFgeAnghRx1JAO3syk8pufkyfllDXg+
+QPWR26uY3PhcZ3vAZO4QOsGjh2J89/7mjoQXWRpSS8aVEtwl2MNZEOok9beQY6/
x7pbbxSgQ7lrLDb7B26XaEcqmrWXUTrcOC8zCc1sAD7sVZ/FBFy2s2i+HYau35tn
pv5WiI6pkMJE7yoqs15CDqO3MCGKvuzWJXV/DR1RRGTTg5PqTfXnTg9+PoM27OiF
Vhm/ocZUAo+ydosu5ZuFbmZRQb7shJIMVdp1UqRgncmAj+3SatmblPo/TAbLjUQl
jE/468XRm7gYypN1rwskXjkZcf/DKHBgnhzVw1Ewt0oqQ065eRBqKsXwi1EodEWg
VIyAcwuD3G2+ft9hefXNPiCP9BUl2dv0uz4f7Fwxtkhp/Q4f+KtjlxRH/4JoeBIo
86VrU32qQ5k2OMryJH5ijrILQbB8QBASTy/qHAxLFHknVKBH80+9pigTNM8vH1HY
KRaSxgA12ZHNCiWiulgD7mvPBOrSXlEzcwiqN8PFc0JzJn+JHdzJvGJm1tKvwwoZ
TfroUIIB8Bv71R4hss6GRToDu3qnsA1shOKH3lBFT2FI24ZDnpewfiJXRGIOfApp
4gKLkBUKuCSiLWNB0WEl5OtzSyGoQzp7BJOs1W8j9wmVaaootKuURBShuPYw1T05
XRtz2+lEMA/5c4JtgnxbcW0/5OMiHUpEl//M2f8R3t4lceTmRrb19qQzPN4nVJei
NF4TcJcYgwK/MZK8kgWRW//vl91bUPO/qQfvMdH4wZx56TfYLgg3r0siMcZXghnX
Pm5mCKyZSUfzaIL8t9nCIJWkctTaZk+ddqQQjxSQa+z3U4r60fPeV6amj/gR30Kt
rWP0dYGVAyTIGoEm6WDwbsNlAp9rzGFZ9PPDRAgeX2uZYO+mIiqGRtMqJFZXbUOO
6FZZHPdTBBMKs3O9Fr938Yvcv31/fQPkoH4xGDEBdA1uy1WhA3mIZrKVTazXjuPj
s1admADVGra6WjtGMm295SzL4IHdwYpKz3NBhwEde0UkiojjWFI8gng+5hdROfam
IAie2uKnp/ZvG/FZwWg5i/fJK1Q5/lS0xJhwOCWwW0Ch5kg6xHJ1PDi6veiv2AjI
ePCa/J6lWReXH3DEGBVEv7LUzSNoJ+9wY9luAbyIJ9azBnNZvH6ojb+qU5rpBM8/
4uUhR34h3piZUCif+tNKL3slEIy31Cu5CdPv0ejWp2rwei5Hm+mlxZlgLhlIvsSt
RI5466tZt6mlV+bwVUWv9MACBf1TY776L88lhtvZHmXJiaOP8hgzSaEWazq8iLl5
GeyJiSuojx5VsYw47ZjIzuYXJCDTtbGa4RwQoHmESFt5TidqqLsfSqpw3cdANuBH
WTJXXMolWrTCDQ+rIJTUGGUTx8tahyJ4QcXEWRbBXglf1V/pPzd5adA5yesn8HhY
zbW/s5wzHmkaoCxFp2U4b8arMOYwcvrppmqqSopmiOWuzprJFhC+I7m+2mpNbhiQ
FW7MeKnTF0inOn5mOz15xbkg0gxf5o7au8zlqueIwnq9Bu3/SwqQpgeZ1C/lHObF
woKgIuLdb6DD5QOoAv9TA2xjiP86fPrL54UDrRAcix7aCHqCLNHXZhTqgTxOrTL3
wT5YaAqyxEB34H3Go68LoOGrtSvvcYNiA06w1AxnhdcorJxk133uAYsL+Tt6nYK3
HPCMSqRjRCfow82LvDItF1uX8nHQvIunmnZ2MmKoMQjj67JD3PxbJcug3AEI5CgZ
OXcShYmE/vimgY4piIqsirt9zxhoG2riLZ+Ki7yDbTM4JPjNafRnK+Q+7kOuzQK3
T+66BKiEC/XBe8PfTtGA63OEBXcxt4g308ocpgYpYS2BBcAqfYVD9uEdTvn0JJZ1
W8scOqYLn2M8Js+kSiAGoLM75bXJy3Y/PUI5Y7EcKTc1ZhHcTJHvEAvncu7h1858
abft4IivfzJDygEVLQPCXcuiCKAfbk8NjW665kd4pJYsAHLNFTIa1mydKfGh2vcT
XMgyWngn/dVYKLIQhUHbSich+lG8R7Z5LxqEnnj/8EC9qNJD9T+7Vrt0E702UgrP
LO1le5N1Z36igP3BRICaPFPXkFgLsvryb8S6yFGNZjOyHtncMObCG6r002mqzW6K
oK02HBpihsgFPlh1KgMIxCzJn3dvB6jwEmGsZUF97kRdVuUN0CbofNFJjXMEDtGA
ns5cVr1QqNIWC2SpppNVz7dIaqHJIAl2Yt+3FrAh5QF87DQccFlLp9//TFFq0JWx
b/9x+RZmYNElfm+giMe++cx/m4OB0PsmDPDY1CpF2dLtVllZtlbpZ9ZoHg4soQe7
gev2+xOxcQDE+zHiQQ2OORUE3zv36MsV0VEhdU3omz0tYEbfbJx0F73kUA2nf6JL
gy2TRjCP2y+dfXDA/V4hvqaj2KuMyGLMacksF9J4VbA9b1j8McbP/E8ZmSsX9S/M
YCOEZcKdVh8AmNOLzANX24dKBPnG+66JcAgAkiM2eN80MmfY+oaiXCJePBvccXq3
BfVH8JKKUY1AXxcFfrB6tse22aZxjmGp/KJepSLbWoHpVGlcaw2faNOfYflbPZYt
v4mcYWw5ye/1rM+yEIK3AZPp/CW0gWJVNEM+O1giabIClOaDouirZ6N9QPt3qSYW
quy5vjFmIQWkfzrwRpXH/PGlfPThdj+2jyX9AhVOwhX+DlTpcYUUL0xrpkNgB4c6
HtzYYg/rR6VrnPyf4CZRrp69YH7sXlOc59sxcec3N0jYTtO55JjerVZUahZ+/2q8
x5ZBW8G2+2FutoKbsY81WZlPTEQr1leAz8KZ06cp79d3eqg3vzhwKlevsxwRsdMK
1nVW5mhuO8iDQO6fUFJl+66WYpkIIwLaHBeleDOt47drTPEYP4cgz8fxkC1w7B1p
9VD5cghMQ/WgZIalE8XvijWZ5KKX84Ur3ywrBkPYZiMAbWF3OEtPmHTS6agbkDUZ
wrHh/lXbq6R7DjhWx4AH3oVlSXlzAvTJf4feVhCvpGlJzcJWbkJoywq3rn9+4V0Q
5BamyqfNvhCvSMf/++kFPBfro9J7qKvqH5t0GD9n3aMvAhUOsrgr1pHKNlfSayUl
uOMhKqzC6aqIg+PeIxlFX7VHyvaB3EjpHYtYWSTGxrHE9+OrfOl5h9szTugQVBhm
zIYjvJQDwz23vIchhF4FctadgD7symn2ErMbq/Bdc+x4EEkAn+2dP1+5EA4Je10S
YiUbaAtSWDWUvI9YUtGu/zVTd7x9x1Wj00qH7YdZD6sSvQuLaSYd6Us5O2I4atNW
zmUuU6GRH7tnu2CCil/Qo8F8g6jwG6yrPwbSW97ZgZKRswYBpky9R8uFP6Xj5I58
qodw5tsEg1ZTF98y/iHi6RnCMX1OuNMU/AkxE9T3b1YmfSmQYkulSZGwvKXnUTX4
RUerbwy8yDoOpotC4XjVI7d/XV64UP7uq9hbAN36tnAEA01fGerrRKJPXghtzcn0
TdXKU2xqroyc+5GSn0afvj6TgPEEOLogz46anb2WT+BEhEpDgf8poZtxHOY26MEa
PKnzNHayJpe8kJnJPEb2++JBzTP83C+YnKqeks6WJoEut8Sn/Etx7AQBtyR0M993
KgxnyJ06rn24IicqmZ8JRGpEipvV+2+yIagd3EbPxIhOUlaG4d8D54u5z6px/2sT
yhkkR+UlpAGknF9yo4qY+AsY8PtQoMuNw2bAkvV177v8gVLFJpyRvAt/63FAHl4D
R0Gvp/qURWrjy9kaKFprgoKLqJI10sNIRiY3NrzpG0WKSVkd7B3dbWk6UsakixRk
MB9/AkUzl0+Hep9YCKqRm8F3LuDmfZNDjI2oHY9Hj39OeQ9g6xJw3BZlDMuzVrWS
nBX5mswhMP3co1DTnst8hfiSS8OmvYM1D0XlBGMp9C+lavz/seAhw+mCpJmVFakW
MWeexwCvZvKCrHZnn2zElN1xxzeKMjKQM34HR6HjIksgiy03XuCFna4H/Fj+X6+b
s3oqwMFif70+UvN7AOOgUryRX6v/j7LtqYAKomDzTtOqFXx/aiGuI9i8pQY2pLnm
u8/orNWPgRviiqU1Y4PFXCpgVSLQ8Wn1C1NLEjtq3EyXdyT1/NZMhrsuiGi6vG+w
eaVl+fE21khLQJXOC39uN+ExP2VhDqjWO3VWQ+NxrYSBEvRgFI71xTFSSpN4bGN8
c7cBhpTyUrub5Y/n0p79MEEv6PCYtzIQeqhAYFuNvP5sHR4YkPF73FT0VbeFasn9
g7O9gy1Xw5pjXw+Kx6Ym3sRT70s88rsQnKlGGRbHGH0jEoiYanqLl0yikox8YH6+
6woi3BzWjq8IK6l4WsdRh3rJEuqM+D71cB43+XleqSCye/AD2YESYtr9MhvRxxq2
Q80UpObhYvGYUAnRWfqchAAgUqAbUzCFrxYNrSsSVCIToglcCVuwO3ZhzHait9AQ
xqrDmQJ3HlPIeQGHQ60bpR0z6JYeq09ove0JvA4adWJsUZQ90LdtG5bur6xiKlZJ
jJt10o0mL82LpyGT2gl52VLLRtKzASHeom8EZjGHsiCFzKsy9nWcoqYKzHeE8fCH
YmvqT7wTP7+hBIMiPDYQrsxH1Zy/TbaZyW1cIUXObYeAMyjHcUQl6aCRXU4v/RXP
mmjObvJ16yJRwV5hIZ+2R6mxBTcg1cb5Dyr0t2K+dTrBVDry89Ex4SZ/nx6JZQlJ
E/kq6ETAS5xs96XSkg3sVRezRdnSdhZgzm+mFX8KdyP4Pem0j1S3mX18k72f2wXl
4XLpMgMty5lK3eQO//AcTp9tP5q56FpAcZ7raoUXreNq6Ab/7Y+e6Hb6LTkGlxGu
DWD+wecaPMkGgQ/GZsxxcJGTXnGz+xvQ4Nynqvn5/Xko0p5ZCbbqyClACQnj/qbO
DkBibNLaVnNelrDFufOlE5DJDJkdAffoSMmpFshJsdB5BahBmjlV+7wEKA/tUvGa
yCBVrLka4jfIoLdTOtIb6HSbwuOjpCBsCSNDI3KOyMz0nhspFZS9+TmYRPhhZ54e
+iTbdFBHFIYAIz035MCN9jNvKzyx9GgyQ5YaRipAanjNjcn1EOsY84L+Y6KF/FKX
jAu1mCsZ/sqCVZabbnJoV07t/kUGmG5ZnP4Ac3CJqPQKT7tVl9aEaaowWV2B7rnR
Bip3HEmDf+LQ2DIexpHFFvyhZcEeOUL3ff5/6JqmtX2uPqMpaIL4jgiYAx/bsrZz
Ukn8ckVV8NcEZvJO9kKqQrIgM8xfqtMKZAPNj+QfSU2O2jMT8KB9qvHKSHnfgUyu
T8/ujem3GHKbuQWOdJlMDUXkkZ1hcpUcat06MJXXODPRgLsaPGrZxC9jFfxhp7mQ
pVAxSkJjMiepFz4WdYMt3ifocfYwKuogv+Qr8yWWlxc4lXwHSUn2KNrLqNWlp1Rz
feHQWQunuw5qwe7UXcnXsIYw2ADPwz/Qc2jc0NRVvkFVz3HomZW8U9GZZQlaIUPk
pTj6tH7NziMKkhzMsebOFR6YJu2NBexiKdy05V5A2JHhtxMH3L/ZUERWAg4/vg5x
UoPaip7CYR04cB3pBk0RG6oHLAQdlgORQTnN6+oKiLtwJVt4b0iArYZJIB60bIJT
INB8Tv5fPNLJyWupOlekfr1PgneMdElddE7NIHJ6NDkrrmRvilVCnrGOF+EwO8k7
GtRnAx3ZPhTNGbDd6/z/LtcVbObRs58+SPbSVDjVgmJ4qeZ3FFPb4ykvuay6Pv9V
jPmS84oR8WACS03TP3R35FLWsiAodhEAJkKtNq9rE+T0zeP/PnPWCnfLQmIHzo6L
I8bx1KPqfweqVIMWeGU7k2pqhmRMwulEn46YNrxDObUhF+NNWyKm+nkEzElJ7V3J
b5leZkFQQlLCtAlM4ZN/p4PwrT52uG3+nQDzo5b/qUDBWonUA92nHu70Pgw72DHO
+tDc/5uWwKOoE8VJONCMyHuAg1CCXiB7AiLeQqkkC6AArTzeUKKewjyRw4lWxVIp
SrK3DvRtBHNvrDC/L9Xm34l/6kRwTwzzL2YUIndTyfXt2uyvOr+gaCnyaZ1A/jmE
rBs7ErXoP4bGGJ330GxXvdk/adqXT4unlGE6i3+j7h7GdRq/qzTp5owOwaREFxFD
PZT545hfnBEFikIEtFgfoeHm+FwJ1Vf4dqnikWB9h6jxe+dgPOO9/V8qsIaYIKqu
WSN7PKruKWPOciSgY1zq7LRQHzpp5sr5IKyG9uCKyItZvDWRgsNuAkED6XSRGhnZ
hyeyR9Y8RyQj3enL8XcqOLhpbvBTUaxHVrVuTyBh3+5F91/2YA+MWzxV6qvP1jBX
lZDR05argS4wUrGcU5sKP6Ro0C+hWuoIC24JLEU1cTW7IcQYhiBuabmIApqry1E5
MoocaQt3fN1rMayfNzMC88LBp32+pLCivSU7nHuVJWIlOSKNHeySl5ueBZ+GuW3m
cc3WYJRhdgFW/SbcLNvBOo2ga8dM8OZh6/kpSa3nyr7hwBuX/d771NRDGyyeii7g
hqKh50qghzjB+C4EryYaM18ulMrCsjkdHjTQ7Z7av1mC6HYi2g12pqhIeGKGT58n
LM5NvSCx3ayKFu4CSy070LrnMtMJGDuVNJ4Scw+qeFqYpKNogGgOYCxhHyEzRlvL
WOtt06FULurMTWX8izvS9orBxavG3y47shWLQBUq8fovM6ak5x3yC6REymwfX4Gn
akMYKCOlsjmh/CdzQ9L6Kzj9uPHk6byISajRdfmNBfRYCzu7N4Je2I9Ti+AY5gPY
7BtsCeMmE5cHZ/Zf9yrg7mD8RlZlMGWrA1jehK23Dq1+MNB4z19PAMK4TxoTh4or
bi15Tt9vm2YV5S5+Nk3FVbbDyBr1FHK1w5vb8flZ5iIKBljYbdQbex6dj32dVX0O
FTm0OKmnnH/GsADj7c+CVvuwWvoMcE0Oc8r7uNUIASJoDpNGSykWqzLjhQP4M9zS
dtFCOAVFt17xMEcjBGj0zvo8kW3hQ64XVj/hpHlYcmzVO9j7Ai+/rH0hW0TQa6bX
JypwblOU8RPdDr10vuQeKm05LJeajaFJIpmCR1rFurEeub052w/sUe3/VL//Xcmq
QpkdanRaR9qBFzDlr4Ruu+RStduc9AW0j4li2A5mkeXEHeHHr1rVv3CwMEgkzS8s
e8D1XlAUt9rg1EbJAsgU6ez7ws/FD6wVS9W/qAp1CtX8JJK1DKlsI0JbpSKjSzYR
w5pe2v7sJSJuwz6FHsD+xfaUCDSdXVHTKaGQJJdd6VdCdgRvROnS3YZkAmz2n8Dt
qwxsORkTBm3awjVTS/riN3gsKAmlX43cSANR/h9WqOosHUPwlMz5tNzDL7RwNM/R
ELUgZyx1Q7fgStZ9QGdSxEfo8u+/WlWV5u3lRJdyAQ+MsAGPDLJ3oDnyUI8YkyVv
iwwMKGbM0xYVmB/X1ARDj6D3ZPLFmQH7ojAFupH7A9A96gnLZRAsI7AO+f0dnQLf
ZadRrDP4o3INYTOUMP/H1p8TnGLEJc4tUWCGCp2DgwoBFrHK4/W6f/CgHfWfH2pZ
aDAmA3mt5xfF3FeRQaQDM1WBrca9Nw/BN3UPeHaF76bf3W6wYHpoVM653ek0Qm3b
WXGLDTPrjKHv2lQs37PUaGDMMu61b9Kh7xub0Bgtgi/qQLrwp0vt84kvkEQVHfuJ
cO8er7QQy1np/8SQWtG3YEYOIfFd59V7eDKsta+2Xq8BJY6W5Wncrs72V4UbznTM
XvHlyeFAl2fVC7cCh4njve/SW9pSX/3XkYcTRTl/o4dQ6x/mvrwdlBQ785QCfX4q
tXLQpORIgqSunfjcz6ke1sVjKURaJX28iq5rKLRuaZ9QF6Mv8IhjiX7XtRcdfL/i
CqAetOsOvUPX69hKiqnj5NtCT8VfLIHaZN7M0HlsvjQdH+SMbfh0ISYy3q38PmpS
Y3npPtMpP/pek+dxhzMEd3o6+9nyRx5UKKpeNoyBWvvujum1Op01Q38nin0wSF9s
EfHcJezd2EJl8PWyhvp6dS9brShzv8FsuBgBMMOtlNvty4a0bs0d0qR3NGHhhkES
jst4hAq+CgeT9AY7uH6PlETwjMuK8g1Qyt3GXbOqmml7xFtvQlJENBsPgCPo0bs+
8/3Z6XIiFaV89YZ1ECBNoOGynRKiQRaMlBJd8nhUbJBjfotn0jC/ge9S7kozFHNe
fNUsWbgt4CpYNPsRNUYb9Y9e01uTxo82fQqROAM6wzj0uhah/7smEvsDXkvGoXSi
d3rLC6tlLlfYPDwCVHhXFeM2cspL4Rh7+1S73+LqQkqg3I3XiuD7HKXb8ECvq1D/
FOd7tdlqv0T9ZUsuExhUfq8WDRC/lI4kstMOEryKLOKRGC93uufo/69el7vhSx5+
zJr7Xb1rcKp4TdYyvqNDrwAWsa7Wh7IAE1aZ4OGlWe15OZRCbOHuCG4xY9CM9Gtl
bFR2i1/AnPEl2FibzN201KC40BJ+rNflwzPI9eglZcBt6NM3QKAQijQNRxCD054f
lI9ALEOAffffLbb6wEegvP4CayW9lK0+0ucsUNck9h3v6euCsbaq7YFVQOZGIJSX
zHqRiy9d6txqHLYdkB0kGS/Uamcr0CrSNm2D6YhKT6QdxS1eqjz1A9afZJbHFIIS
Cl7cPZ2b6pe7A+e3uWhYlUVi3NPR7sKfRibeboBS42HWVaKEVyDl+ycVIjHqAZ+f
cMNFg4/XCrQJF9UfDKEw4/4A48cAn5CWnuotKjhiIdmxPjsXC+f/x6Utf7XI5pcI
VBC0I6EIzEBsbTFkyYEJUwR+zVe0lviiFRvsESwD4A9VJUHoYXsiSsS2gnRdAaB1
PnRqaPwtr/oMDnh4bfI1N5+djgAYWrMKxaOwWNyKGBGXFLe8WtUaEp06RaPDyPvX
+8H5zHuW7AWm6c0RkOI7CEl7CADyGXVhlDJprFhNQtm5akcWki1Rwz0F4B2ksUdp
V7NmLNhoFJh+j2WwxD2a6svOTFMOb+ZDVG5Or/tKbyE563UNwfLiAjmuklJ35BT4
tstY5m4E64xaxQqWVjDZhpV6Ye4qzIS1BjvfPatW46bIboW33XmytRXa+540vAto
gONQMy0eSAZ9GyAabc6KkEUDZAaCZ/u6hcdWJHPZK5W9HdYdY+/oVT8iVb5DVf++
pIl7wuMRWl1HnDJPLXHFyDFokmvKxJRurvXpDwVb3TmjMgs7WPPXOjcG5O9kXaVj
8t5NNFZR/67HHQdWk+I9i7DkiYc9Q6klmcnnD//rW5QU5UrS2nrZE2fP+vtU85sJ
Pojk3MYqDviEMT3w2IVlkEC4D5zu25tWXVEQK48A3zF0b7fgv9i4vNggbuR46R2d
RheDxnaVYh1Zeio2XtmWbJ9z0NPL6J2SdAt+b7zf/yh9IpzHjupfQSJdynSEK1/a
A0DAcxqzlaeAhXufRIDpoy1xAF2SIMnGmn9aGALPjsP4MO38oJlFaLnh9obv4fci
TnmkE4FsATn7n+vA8AkCZgSg21xSzFZq7cx7XEe085D4SNTjY42sL+JDpxZXxLUM
+SVXSUKGCO8ftnpiqgtCZY1isa0ChF+vjqO/bi++3Lb3nFCWwsN9s6fesalA+Kgi
v8HYCY1TkUnk7jx4jW94mwcs+BvclpLqJ+yrzjxomLU1cgnHZb3HYZZz3itZNHBB
m0ib8Cmq4lHBdZeT1u+bsHRn7zGreS2fiWxGqmrXBAMrFB40scSYIn2crBB2cHQ8
Ehnw8Dm4moLyTg1P4695eFyegTeQorQ+k6t5ANyyJFiIGiRlEowIP6SsZfRlcYsG
WQ1ZPC+r37DOnvRWGSL9DFt8jMGHYu3pS+x99whRDdtuTFhhjOM2r8EaidxwaVdw
HLK4Jt2TnUL9E0U10WUbw9p89GH8zbdlxgg5D+8h47/zSZDo2bMNNx+sm5NuFI55
PUBQTYPR+X/YTXtT8BkNqP0AwH9q/vk+kvZeYsIDKTGe7uqQgBlnZDPky0tSVp67
6kLUtcdVR7EIkbv++TeuUjCm8tE8tSuxdgPjsvHBFo5v3VMXQQ61yRazg0mPQrzL
94uJf6R0m8Zx0gev5cy17yyV4Ao1z8mL7R59wn580dKn8GuAkmjLf3tmlhSwxadQ
QIlDczQq7jAAoC6hoXvmuxYgqUshqw3ZajRuMjH2aeeKS97wmcoq31yupvFCjLxV
fGZBl/Qd4t0brIE5RrOlkZFbc9CaoJ9CaHehxqky7SyNXoLHFvLKas4c8Go2VKjd
zO4H0ygndA7KRcy2gefGHICFhKF8MKbHPBvVSnAUY7eI4aQgdpCPBZjjFxRm7F3l
rfkrUv6ilIy+86knSL/E7EwWvwFmTafSL/cnBa73ktocKSx9VnM+FEi9YjmF6lP1
xDcSdt/Dqkgpx2p27sqQpyw5u4YFt9YCER47gkfYlmYHmXrKImuupDIyNoHIk52B
03rJWk8CcJxo5/IaapKsc2F0GDxPXy6NSAjuUuhGVZjPUCMbREQvoK2fmZm2O/ha
ZiG7IPdSo/FgBODUuEGlnfjVhG3qO79d8GX5iFQyCdebCqB//JpqySeINwT+Wcsr
nmry5bFcOq/7VD6tEwSDFBko9Uyc9oz4FYtRxnTj8SNgI//6bmjm5SEmWMng6I9Z
udqI4jRsAEqyNkpM1CcPBZBjDat1a0ZecfOddJpmKU8qGkqw3ZJEnww/p0mEh2Vn
35CzdAhqBjQmFBjpN5vIIUN9HGS09SK3ruD4BQEvyjNrfvgTQ5G9EGAi0ZhhnTYe
kwkXjRse8apiDJ73yN39BS3CXuaGm3RpfU6pXtUyjX9Gd6Pm3iilE78zXUwh1n+w
Rwqxxoy19jOXpB2GC5qY8j9jFZuRS2QQSQaGrJXcqOcG2aOk4vU7J/yl7mKZs4lY
dx/ULatxnOxuiEjdxAdn9HMsPgm1dRAGD94YXWCF1DqvGAfdthRfBCyv4e1lidfl
1MuBNpHlSaEnro84LHWIEjZ9o3OFLsVtvQAzJA2PxWSBAhP1RaiQRmsvl770op6d
vFH7GWnDIv3OFOD8GAaGjZuXsT7zUNoGkaqalftsBhA3fTr1dzP/8RLbST+bPKL5
JitFI1L3ZgIw5omXSOTiw1LaREayci9Bx+FISQxEowmeAmoApoW9SQ3cihG3viZx
3O+iFWytQsVdYQ0RbYU+lH3vi8wKX4tFxZtA7U9YX/0GTxaeAml5eHP816BEaJ4P
J7fY945V1fAgIJ5Cky4BuBdRPewuaTKD9CeR8E7QGrFaqsWG51foLgOUyTXTJZXt
xQcROrQvLtCqw/Rz+wqTriu06yK6PYXzaDieGTJb3M9nCGtykealYnTWzLLQ2I/j
Ogr58CPFA2Z7SqD4H1yAfti982ubd9RJFv1ltV0pE316we4mTKxWSy52dZw1FVvk
Kip2nxJeAqQsyVdXFbC9A+noXAHQ3VMYiTIAB96eIyXHnx/YEQk007ZDrZXDvAqJ
KSoGhS/UtE8S5u+3KLY+FMsZiBRiwie+VxSWxCyxEZ4AIdhCJ+jpnki272BJ8C6r
i3/yrkm6qwKohNMnLgW3VUiKCcsBcsaC23gjjtHUzuVll/nUC+L9MqzTEUwSfE70
CnVUoKDseLDX3pf4bcAAK4b0RtDiCie36Av2iwU2Ffqcs74hdlXVpnWTU065AjDv
+6DggqK2JtrWTxXLDLwFwhXKF0LWQOt7lKPaSvEpPW1fLBNG8Zzug031nFROzcIE
GjrR+Uc8owPiFJtLR7/p8Xxu/gMCNIqXLUm7DrMhNk/y3mwMYqc3Xs921ZRM1/OR
SJf+bbPs5O1gs/liFrjWlxEIPpw6ObB6rLo5vMmlwMI8TALBLzuUHh1inD3shLDt
p9ORx8WZDM8Px7/HgVMGnqfjFgs9SF4z/pvjpI3CDxRO11F4GF0vhXR5THLEa1fQ
rNXsJWZ6xtKpuHBZasXWksM75v5FJJA/PALM+5EFHvkhSRIf7HM3PmN8ErHasBsj
2IZdpLPa4XjH50MRQ77fmaVsxNVBcQJLsp+B7tjMQbfN5qGpGA/zQ8+ENrI4Es6g
CEOFhQcvSDXRVpkmgSqPJdtdXBjzLWM29TTcEfzQUlHs80bFZLpvVrHoptAsntbC
1/euyi23GloFLBt7Oqmxjir2T1SIpHbn3GZUzGDxyZ/KVtNdZhwHGzCM9f0Y3iYR
DiAYg91zBNdAsaAwIA2KBHz/bVXKT9E4ozrJVP9ocD3joKpiHZPeuSN/f1XslcM4
rDg/tcA632o7fbLltaFxW8pQvFeWBuQw0dT+sdvI05LXX8uLjC9UYb/Ez2XwYKOf
lSMPOyp81vXJVajm7O80SWl418XVEYrki46uqtCNkUZA8rtQ2p2mZhWJTI57qDrb
SQVRplusXC5SRAxUXWuPV/rLAgLQxYCYJfUII1qQ4DvezoJJVrzG5eTv5YqbeNCs
qxHyTuSXDs+LiVCBuD1nip4HXnDuFKxQVpVMOzVTJ6KTdFe/Ao84G1QEIfa3lXhK
wpyFSZ2nOXZGuALch7IpR7sX+9DwHyPAGabj6YveItymVP5SiCVQwvZkxLryEEB6
4sToY10vH2V8/XIt7o8BfD7w04DLWlvU3vKofZ/sBNVMz2rQ/kOd7BjWUqow7r2B
dzR1vAS/3sA/rpocLzQ2j5yjP+syTD3sCg7HExWSk5uzV0/JGIJKofyFLR+sZtkk
qDiVA/kd49DyWiJUcESov/Id9WOn24GI6yaPb/Ha62uwv548aMdY2cPvtG/jDVQL
7xTG3SRw0Nk/q/9/A128+PjJy28aS5iBv5sAjXzVt8tRBJ1LwddtrzEz4Gdu5Kl7
MGblKFy4k6e5ZBCVoCJGrr3KohzPlU4sbtPH/8frxBhg6mTTfInco3Yqg/syiG//
0uL/g5Ns0dV9OG9BREXtUxFxqRFLxJt8QBSeLC6rhah+bbqwr4kd+GeuItRkuAyK
1j2adADADlaj9tSMHgd2mNBYbTVzNjkyGG4KtTHasq4QADpqIC+bDjdpHa2tX6C9
jHkJxeXmVHe84tmVIm4bdgNeteGx2DX804EjSgk5NwRUIk9BqWqNoGpCjF9SfFSs
JxhFHc7aqMB+r83Q92zzNpG2RII1wTWMSildgQY44ifEwS8ZD+I2t2vkY/O7bHUz
IOmWAJ9Qm9gkzHLQoMwDRUP2Yeb2EMBHFsbJxLAt6+Ydd86yY7caMKBM96edMhaa
sU3SXFBqmL9vs2LIy4BLBQNu80yqhSUTlnWdu3kZI0REB4TYqvePXj5hbef7cAyk
vZZMm2PZUBQ6TEnDx1ts5uXEdG0yRG2dQoODAuotE+amvlXsvl4pwDtfaL54X3se
dBQi0OhbX8aE8HxZWJGZTKBPRYi3do0uzvLB8Sz81IaU/5JYOquQMn/3ndW8vGAc
zAcsv5RxQPilmmIUPSxV8WsyW6/2LPl1O8PjQ5uCtzE7sZk+UrW309JkvH/isNGf
3saeb8DCaMG642S5ilZoTvct1nx5K1iVngzQN5Odk7rzhq1BWzCw5Mk7XpAhSWQr
0hjVxaGqcbXBPaGHFBcWx063/4qF7Q2ryKDpR91Rr40hikpIvIc1j2UYbYQR7Tta
funzBGLrVoBjVj8KVE90rMc6XCugJ6xGMITXrZ6pLpbFbXrvV8Vx2a78jc3lpqev
l5i9kwaCON+6HzR+4WYTV+FO+aaTyaN0qT3aoWu3OjY6ZGdp+giaigEq0Gw7ED7Z
CS7TyQomB7u4QRthdro64E9o81gn+GLrhpm7/QKkVzyckTSQPYo7dM9s5z9DviWB
EeFz0MiuZbxogW+A9XL5+9b9w6rW2bAbqTPYYOyykk1SzwhuvjW7Cy/yZDF35YXQ
biWhbqUnkbSR0kArG4btdcjJ7NEsvCtzqfTsGzJSGedQFDy5Ax5sPHslvAxQvsEo
15dC0A3SL9qAJA4pMMs6LHhODctKLVFvu+9n2+kwruvY9WQ+vTA8K+bnsYAHgEtt
C1DPUtprzruzEJB61ucrE0bXJLDZ1EbXYB9U8hvrXnPY9RO1lLtaYzhE/RkHJCEp
s80ueRU1/OnwrKnrPjPf0x35z8wDkmWiKAlTv1I9d5/AtqdwWHANEb74dzw9oMIZ
pE+Phbut8ZMuGcnYbRI1OZTN9Mt3DUfW2+MtFDygFsFc8r28/cXF2GBOvmJmiwun
68Xc90ieF5/Vji+gI4s0LpJwC3Bqu54xuZJ2dz577Cd/D1YzRUvqLvvH8hRhAJof
SwLuP69vv2rj5/Dz5pV5wK7yrT+3819NVnQ7CSejO3qM/ymD1ypY+6sv4ZCUsUI9
fY3RgAmxZT36t0I+DYT5lmZBzYqO3s/KF8YZkaimGU3EtMWee5LTrcZ6fa2o0TtQ
Al9zY6c0lVb7oVwyd8NV/GM/Vr91qvCB+CkeehvIZZT5+1IS+ksEGCUHC78oLMC8
2gxSoGn829+pGWoEqicio+HWOPQAOo8cQiDjBdgwjWqOtHoQN9/UjmYR/XHqIMNF
QvPnrD7TNqZs42k6+voxU1ZDO/mOrB8ZAOFpN0iIgKyXPnfmnIAfvNyqgn7v8EIe
sLwmbxnDMLeAgzpyPhIB5avUWz0TqVDwHLOSwkEsji0jp0p2jT7tvG5l2PtUeZci
nJqcQTj6WUwX5asYUBqkaDXdwoWfoRx5RqwIW9LImIfJAvhrZoBbqQwgPCPDuHiB
Sqc4RyXQ7DgvD5UCepoEGrixkWFgUJ0gGBWzlmeMDqbN8hK1ivdVi8dGfaxX+LGu
gjAZupA4w69VHn7NL5Ku5QSgbcSR+mPrasPphIpMpOM2wknpuUkN87HszsjEfJEX
+QQtOAJjIgfklSd/gWxOwyo2AGWUG7lntxMWGQCGkqRfU07gG4mKugnnQOTvWk5Q
+ixxPwiM4qo0qdORQF6374reXJ0EevjQSeLrVMMpkd60X6fl6FCYv63iJM+SHddw
jmbdnJS/3vIW8KMimvkMy4Lzq5dYGsf2hYbBDPrlsCyR24xACj/zkuO9CW1WhkrW
jfiSwk/gP4aO2ts3ep3xlSIqkFGbdcR4AjhD7c3hAbTUl7Bh0Fl2R7WejLIdWxdx
HF4WAZx5M3noW8nK+gUgfRQc5UYN4G3UQ837uekmy9zy89xgSBcrorjGHuxqvEj1
kHKAMLODAIw6pHDqyxtCGKSRytFNUAN2Og3YT6RB8Ytjhbtg6xYEeRLHJwDWXben
fx+Hv80zDQmy4i2cxKkmo/fJLSrJlTh20UQOhcgfIfSydcGn67h6UkoKgGP62eZv
9LqcFyyag9cl5MVinlaY0cenOnNOGBX6XMtGpZQu4eXvUJl6I/PtxUnriHuJU6Hz
ciXRWbROEBW6puvA8KCMPp7e8tWAL9w8hd3ZgV97oPy1wg2jVolI+Pkpmr8E2Koc
Ayno76fBwcXq+Xk5vo1Il1jbWWkmZX+iiwcsJXJB9Vy5PgDEKlIe6vLU44HXzTKT
Rl7d7eJhKhlSLD+IIaM6Lh7vdE0LKzQFmfHvyTJKqqc/OFEgy8gFaApkW3SZt4vQ
JrUZK0J5OtfACQ/tT4JXQfgc7G0jPtHOg0kpaL7uyhgBQGcaetumNbZZ2cgFTkNW
vD24a+noSh1C/9RxhKYnM9Nxn++qUZ+U0I0lKDwU4Fk4hz+zSiH5n/TWleP31etk
v0hYpyNfiRBciRMWVXYUxLSvteklV5OrzlHr3Zt1y+AZ1gQVq/KJz6mhfNpO4LcX
QMNJ4evmN1k0VQOfglyC7fc/mKwX9jY3bKplJ2ZWg29++AGonn8GfbTz8HL0XaGN
LGgICZprhjd2Vp+HKA0n1b79CClFyEdYw6XFWfR8uBJ0c410/Q9GBUxZ52ZBn6lc
bXmgLZDL3bh1jRmuvflz4tYH4SaqjYRfW+2IwEQocPct3L3jFDQJ6Ngcp4XE5WE4
/pzKLTY0etBCx9/33OyLbUsV3s9VB8DtsuFD2dQGutiqazMep/ZKizMtC3ZzWk4m
ZONUmE/qmIw+lxsjxMBNtRpndrss5PDaCHlyrViYvca5mwoVzH+yqWyfssITGP3z
2IYdK06BJXcKWwOHLfi46Bo5laZvfEhyWbdabeKw6KyyHe7DqOlswNRl9n93YW2e
g6LaJzusMLKiNlVpVPvIUZUa7QCzbQ3ad0POj2SzCJk2NRlL0KniR5nW9PjvTDMw
lENLUcxY3nv1jPKT+pLDLvexzutscwsMAVClcpfIPz16IlU28GnjlbCLGgvBfcJe
cFt6K5eAkTxHcz5/+tUrH89AFTl396v1agU9U/RURvGDTrzpVE09laIj/3ttwT70
QiILezE+pYG3EyviVJHd94OGzT64ccVSOU8uOLIlteq4RP4+JbC5N27QUKQCHunh
keli6WsxpeyRSIsyknIfryDM9sQ1o81c1Bu4mZ0IkzYQixvSj7W5eRLlp7byCEbd
cbgXam7jX0gSlm/iMJkYACngiy8vFvbykU3XKj64jl5UBusv7+Bd0arVx5Z143mU
zxo7syjaC841WAk64MQ7GUgVCXAoIyEzjlcOYSX1BpdAnp/lfJfWtmOr+5/lweY4
G1+D2cczv8PQssZnr1FAIxfpV1SaivsR63r9mzUEYvwmi8Hge1kBhjVNP9EBkKWL
h8nlvn9J+7BwsduKsNZWf8XyXHay+C//W6toYmaDCBsRZDKI11zE17UaywWQMmI8
c8qytDNOCm6GGZ6sg7sThTPpVbmiCTa1QlOqXjetYemWt6YbLV9Uct6FesTJ23Xe
ck1vPli+VG6KbpqcKwWwrinTK2cxzXlqUXqDMMgBUXjT26MYQFgUhUGvQe3AP38L
g1GvvYlNgkluaAw3VUapPlTfWD49aMGPYyXRkzlIxrtj+ddl2EV50jFr7mZ5iiVc
/ba47v94EfvLLaYa91dIdUG1bzp7twJm2DKvRsXnHFxX4YC2M9Vnzt0Zz1mjt/Ff
Xn6wGAswx14gdoRd1vfb+v9N4Icv8fLeM9dzdcUjQu8ZWMH4xLhGBKdAteAY/9PR
KfvVKewUcJgYpEctl7QDPB2Z5RCRJKRY+80N8bWLYFxT4AI4UhME1qyG8TyfU6WZ
MuqzRiDstN2IkosnlMhGxi2cz2mmRZrhRAZDalItrqgfF60MvJmrtQiQlG9bwnTe
0M2w8JZyN4NpBPellLnOWcN0NHCCMinYnm2yUOzaIWUsT7ACxnx+0Fp/hyVCc/5/
C+ISqTmcE+tD3cYb1YScawsFdEEYzgIaU/1zyM9UC1bXz/CjhL/v+AV31oYVq0Lx
HD1or7DEVDBW7o1UpUup3jUBNUbSZeQfc3NTODcSBPDROcXuWUJwAFuG+L46OYCd
yAFFMPJLnpUlLob53rFLXVTUoIwwVR+ZwvCM0JSCU0kiNlO425hF8v/vcDlUAAvk
gwr/lxnIxRw5bT6uHaqGSffMQIC6WJSyqkbhRdNWlrO8pat8XX7+rhaUnf9po8G7
njK9zZn0Rn4bhFofdypj7dZUX0wrWRLg6+ygmzp9sEtZfAC4TbZag8tHt0Wk3ThJ
pjpeJbBXuU8+kdIgxf1py3594IAY2gbU7VjFa4UNgqCkrbWQJMIz9A79fmrPNI82
eN/EoasN0D2IkjAEjBqnz7SIiM5tQzZkPNDcTZORlcSFEnaV2JA4a3x4gVV4Plx4
lJkTs7a0EptyohXfD2or+eT+qHmEYtIIL0JyB8sUm110aAKdqp41UnlrA6PWjGgd
aF50Wbq+vpwr/vgWsRrdBilCM2wCTRAnnHpWPIoCzUm3FQlQB9P0uS6ZRWXWecqZ
bPtf6L/sVm1LddRxR/vEaVXPYz0ChrPc5puUdRMQGQjT3CQNndSQj6kOeT0V2NCB
iJownfrA43Urq6UeRj7Obrvtr8RoEEYTgWdi3Nsqym3p7tqaG1ShkzVuXoSHHn4o
jSj9K7GIdt/iPW/BYYpXMmHRQXV/zMGLnBXwsNFfhiucDBh/PW/Wn026MjXeMDu2
nZ0Aja2vORqMkS9RZbqVb3x65d2r22cwfEPDMuBxJQxJtnE1nZK+ivNLA0OGhtZe
wc6v6YTNCALpkQUBCE+LtILzOvkbRi0dWYfkdaNyDItUkxUIkAaka1ue1gQbpEJk
eKMjUvQQF5GtwgfNzsq080/U5kkaIFQ3hgxn7t3d9jmPrCezuTxfswXDURcJzfG6
F2igtAhXPbRGAL4DHvhATJQNeAcj5W73T5nCnHDpiUL3h7JabBFlPzdpfYdgOgcB
XaTmrcSSIIsS3M018vQEJTaInz4EE2RaZG/RX8xTGad1Ih3QF7JBV3205Xl9ol5S
znMXgdhYBTVAuyyn8ywO1l6wHkjU07KQ2faO2otj4y8EyrRO6hPxMGJJaPSh2dQU
PXlrAJ36LumJP3PxTrPPMWvuT3fWI5ABgeAunwpqQ6s+/qrF8krdobhJ+aFub+JC
bYtwohuhZsPPSKXZHeX/Nt8xexmBoyiKJoeUhdD7dW6MYPbbWJ7zbZfxRYzZohrj
VUUBnGB254qboWX7D7Nal9XMXzE8/lIvm+Ifq5n4AceHFVimLlis3pUWqAiYp9Hx
CNTtaCcvUnZ3g1yYl7SJfWBwOuXh+vMsNm5x1vPuIGCz4OPPam1ui7r/CuNR0T8W
cyOo3OGU1NfTKH76t/7FaWe6ae6JWN/mw78eSBdFjHq+t2jop/0afmd0gf7I57l3
9jZ82YINvmr2CPffVGLA0eCkmCj9CGiWUBWcYoOJKY0nC32xlE3TBzIhDte3/H3r
FR2kO17m182sJmbRbHEzQkXTxp0zzMtrjogrVTEcPA4+6Xu2Movq/n1Lzc0U63sz
VIcVN97EkkitkIAaGnfqpxlQuZtngebLh0PNaoeKgyxD0FmdtWAErUbLBvevJ72E
TWY4m+y/0OvGpXlVTqiuLflohZf0Hr25kRbVVZlUJxQtf1w70BbUNLaUo1HEzraD
+UZNNMBbWrnffb0WaWn3egk0WCDGEBIIGSw7UVkKDH0PztjflRW/dZz4ppScqeWD
ADqulehPPVhqSFXZrPp/fFkYA6n66SS2+E7fDDbCmZRoKeZpB6utl5PZ6XXoD2Ik
HHzZ1ETwAlkxEnkopbPjqr1JR4ZXUAJhvT29dd3n/r3CuYWFmU/RYa5y6NvOqhsk
CiG+ef19SyhPM4Yco5wFvGyk0vlaodJHm/FuSQWiAVfE8DqHFhetOna3EDPEe5xb
GaZ8cAut+fKdwdVXhRjzIAbYt2SiiqSV6jaiJ8VTV/S9dkQQShE5k3aAb/eJKToq
FpIsKr7Uai0OSOfQIEVnrYB0jaWXKCwY5kFMGsY0euQmclZ7reOmtxCwTWo7vLT4
NOZCrbr9Yy4bY6t5m4LoQAjX+cEaE6x6SuF6thwiLiHLLrtasLf3fggrm5cuQEJS
m2eQS5iRr5oFxTwyEVXOtEr+3rS9G8WQsewWlhAnE+2bjCp9VpxXxrXWEeaWKiaV
w8ovrUT/vMuRUhCQcoQtYUZAXk6BiaCHmMfwhut705RiB10derRd40bqTKtIEyoY
Ok6s4uW0J5qLd06zUvbbXRRTWFORb153myDa8Z17nmO3iJivVlK9R8MlduCB11MN
P3450flCO/fu2uhAY/RzMWaXNNIRMRWLPUCOoDHPf5ic94tfhVBIv663QLKU6FgX
cYSpEcPKfPUEE5Zf95gZNP49WZ95N6VSzkd28lOLctNn3psu/d4Oc6qVjVkT3fw3
5gEq70orPQ+60hcQfbJZ8Ka6tFeTDsB+xz3b1FWxbdUm387mU5az1J6BnaqyJ0kL
ITo8JeLMh1Xrswh9kS2P8rdr6mvN2jSvaavwaWiQ3P43nFOb9QcsQREzrC5yKHSg
fpca2Yt+3oC0ncxdoarRoY7xf6LpV5MXe8V/n9CE9hawbCUYS3iqtVaTg5Mc/4+o
533GsFgWLUWHlvtNYMetsXgVfZ0l/d+HZS31rISIzRmPwTWSQ2qROKxivXL9zJN5
2cNmWIaogzyK4uKwhcVQy+T7KGqp1i74sbYFvAzXZh0l7ScbohSDKcTIkG1xPPFG
xEb7qabCVvrAzP6jr2HDlal6DI1179biYiQyicQlNC9B0ZOgwtislE2+dN/UpLgx
4Y8XZNOAjLxTUwH3hZqijZUybRB+WS35NHWt/2dtVrT2wqyrOOWbA9q65l7oJ2K4
sdvj79aUl1+ttwVlDpRWzLvfB5bl+Ihuep7gWiXunEZoS4VHWtlmlM7xjK89hxf4
14LQkyiOIFrGm45zUq/E1Nx7EuXQAh6rw9Dsv3Dg9Nx9PduBkc6u8+pD5up9BaC9
pHW0bR+1UTqfZmXFAi/1T1wbMvn82mkDavEQIvcQ1DSdJjQ61Mc4WcWNtZYPyR6/
ZRSCwhZ+GeuT9Khl0Etb4TgoPwmqxvGnmTgA3OpH254qaIkFUdkoFEPKLq1UM+py
K5p74urle0GTqFpLoPz9IcQoCrKT7ACfeRXHyvGL2R/u4Fj6L1mu/6ABJANVJEgh
bbeLIKXe4TAdQd0E/CVLyzzIUkm5OmcCbarwH4In415HwApWRtF3ZWTiism/USnJ
RwYjEKZNaS98hlu0r5YCcvPjwcsoM4i/FZg9pvS+mEKaKPLfrArvmQarfh6Eqgwz
rFYKfcp9ef34KkPAxuJPqqhPxUHj1DbJOqBHYJGMJxuV+62qfwGTYbsYEoz+QFoz
IwHPHfvPbZnqyRM5g+iZ7oEc3pw3xMpjyfSk0SFjKg6uxM5C40tW0LAAzhTIoKy3
LhlfnVuifdZrC4WNNiBGVnG8UXSOvRInHsbG4UWNRYlJVtYhCPswCuW0opZcYsDg
g/vAHa0xaDXzPJ8vcU8mr82FhOXYqxQ+ji/hLbCZ2FVYabxObSTUGmTQejk25scR
kyUKP0qbPtE3Yc4FG4N82poA4gFZVZS95uJGDW55to/Yba0S/X90eZhtnVX2Qzey
4TjMvyGt1Sil+0paiuAJKKgkmwxAQaG/lXSJjP4aOcdVOm225IYOeFbwfdGM91xk
e8bHbc+XTzaA29E9+U/wIbYiNk7OsomU1l0hFto/aAAwvTnfTV/n/U++9ewwS0pv
RpF1cV/NWPf7p8aEi8R3KZEiR9yyXv8DlsZJC0z6vOt0qK2JUCaRsTnHxH5E0pTZ
tLE420DiDPOvUU2eDX1Hzk4R7NCscw1iqB10OisQ/u0MCwL/g3v8BJtUMo4OAmkM
rpe7Trx9tmmYnWCeudI0cRYH+aShrovgweY2YAHSt6dd1wXj6wWs3Jx/5+QN3Nzy
xxud6O6BHL7YquMYtFCovZe5gFRg1y3XhU0UKkqkWqoQNOBUs2yulsHv6mvDehKA
1jUHJtGWrOr3dO4mAO9Ggcp45dokT17nVxH5f9dO+5dUB8+X7J9zsnFgGVeod9LT
lfJlgH+w4GvX8oU0D7Z+7h0Z69L9vZMZx3GRQcnRvJXhqoABDqqQpUEcH5QSEhQl
4XTCBZA14SvwfQEkue9xqvjoa1ZX6zZRPhNE2hPkBqeebmg946M62TJPJQzf9o/D
dppHsuchDNjvBi46lZFaG82izsn8eB2VayAuvUyRW/OIBw3gisOIF9N5IL/AZKUC
LMzMt0hd2Fu4hwJ3gyfi8fLbPX8gGfwVPMTpfMpa4HHYh8WwzHU7Tvz9x/V+cfWi
yNUDtv6F3zbBb8ro5DuyaR2mhD1LWT1SaUCv/4tqKwnPlr7jXKwYV3qwHhrjlOSr
gOgEOv6mIgYSzjQ9JH10UPdxbXIVrCOgQLg8BJa8/2y7o18l2y9KjusGa57tr/lL
R8V07H/PNVDlNt61KtubQBktVykKPIQHZzQdHNpNRHpT0X9JKu0pVPgAmugYRbo+
5lbnLIUU6WUAliqXH4sp5Z76ejVp6h0gBxHvkRnEHNNhra1U0bi8YzCBUv9WcIYs
JXCHwC0etJ6U0EghvyDDiKrnx1Ew46n+LUagzY9go5wRmHEmrzrRt4jQXEmMyAgp
qfa8mwjsD+xCpM+NdOikDcnpy8BTrdtJX5M/KAcd11dmhK9QykzgT7NnG+GRZzAd
l3d/EisK5/p9SVcO+SBGYvRu6GY+lgwgnJWMqPol+U5c835anJnRx1BFEt4xYYHe
J6XjajABMOhKiUUFzV0JIcvSV/xiPk3n0YTXlAr/QrEtk5fYIfJzNi18RNSZ3VbY
smPg3cZmFu46zzDFeo6ILSMD1n5bY8qV32xeG3itN5foqZ2zxqkcLkyoDyOqKWvh
3/R76oYVBXUHrTbo9B3bBEydzATQeQ42dQ0w6Vy49dCsOYJoCP46Mx6T3aF+QpVi
faslPi6M91iq1AXUW5Lm1n37hkMJc7B9AfdJnL85Z9f7Rlbth2B1HPAG6JeBucCY
PJg9kZ8GPG0rBTeGUALM32yeyc8yGZFh01DsY2VrZLKDeIgsF818GCSMW9O797LJ
ZblJS6OI3ux1lKjFz2xoyb6k68zHeaeabuAT3qHh7Y7+CYTmMJ47HWhM6Y5cW8JJ
Hnm0fEcsys0KCRS9AwP+E3p6KDwvTHkucKUbVOM3yvprHRhni4ioG8LKZaEQ6Yyu
WJ4KyoYzYjR9UoUJ2ddVcGoGyMQYzG4cLQ6Vd4rU1dxWPwpxA9yTaspPcriirtmE
vm2/iU1WtRFuzQV0ZgEhgvV6T0BvLBYkJkQ39yIPXpu6v4gzVqXuNJyTybnwTENq
As3aXD9aoguVCBW87l4UuvKIuPAvhWltAFfs2BxIrFgCOXfl+iu/1oHtresQQCiN
5pbOP6WIx21yFzE0HSBswaQ7iCOQppyguyWo3G8Ly+zTELIldQmJHeWtWpCVjX0c
zNgPRk4yM0aKgiKKFcVGm7tl4DIxS+jeqSpV3FwRuPW2l600IuUKuPCHEEJ1lcfD
BoJJpuFRSNlr1NsTkp1x+83ab6Om21z/ygOhx6v0t2IueJrb98TuBQy8YQE8zO8M
/n5druqrWLtxH2FJR7FnPv9pV0CoEdfmY/bzZkyYnIePGkseDzUU/2n0keSDLsRp
oqzKiSS0iPtsxfSsiQ1qMtCxOXiPelmkZbgXqXaRyvgn+XhHK9LdjBneGKTUPLTd
qoqzq3Afk17eHs58o6ekw6x/G6nSaEKnFg4yJ4ahzkymb9khDUgi9L8N7stbUzFg
S8gVf6beVN6GmJhob6fSoI+rIQOrSjGRnHWzLKqccpk/Y/4oisU5fM9p6lT11Ei8
+Ge6uYIi3SlC5WR1rDHoVU1laIGryHAVT+XYB7uY6MJr5S99K3mE1VJIR/ZL61zu
VSRwtzUE7giLbMELQYgoq9zXtBtzOZvuJ4GJ0IV3U8gBll8kKeH0ylQcuP3Nrfx9
KFYsigD78F0BbgjVKA0cuKshJkOr5ZYCzY7Hs+rkKEl621cLoU6IsCk539fvShlC
q+4pi0YvnIvvoNo2E9pXf3Sv+4G8hc6E+I2s3aE0HOwODr4GSlFyk/6y9WIiJK04
GlyD9VHiBuTzxbL5WYd56Q2WRQypGECqQM5iCmS6FndEMPuAbGyBUjVysC58W4D/
o02zVQwq4uKQEGgEyUhBGO9MpxNOTQ4E4T8Ync147y8NqUTCm/I5ZmDMeDbg5/uO
zZSUxrTq4g5CCWHXVRB04NLQq66SdGZ3LmI41AXy6FgQtZmfE1lhdui42ySl22Gc
Wl+t7PIKpWbQoWpil0/XilCttwP+vjjfuN8OFOZUQst6cRIXCh0PkOrtQC3jtlpB
XKwazVVQURP/psNIOOEGmINtyD2J2BWCmXJTnCftWZniHhQiP5mdWODmOq4ODpim
fZFnGlbWkOPP5EsSmyiOzUPX69urH6gz2dAjNK936X737quv7k6hykH+ijdZptLc
uYUWubRpZ+HqIONMFORyIPntkCFwRO6NnG8hb7yhMrSUlHltAAhtHdeebbvzoCzo
HYZdIH9QlxF9ihsdoC4L5311TWH4ePK1A3OeIeGgDznkYZg+6M2QKIDK2OzsDKff
AuGKwpWGJGIoTaM4q1JcIj/OG6Ql3ivhJws8c8+6AwrWzWHor4r9tJ0VFykgAt2P
esjPKTwVPXUzoN9CgMOn3+r1xYp7fuZEBACSGaaG6FEoKMkylmVYBZxg6shKEGRY
tSycSuz2KSogQ3e5bFUOnv+KlZ/aAD3ALnIGX+lX5WudRfT3ORhB3D559rLbOyQ1
ryvG3D6sFTu/aYY1DsGOmU9KxDs0dKyLKJ9RDUQcMD+sVdDysvW/Fi7NXM4bTCBP
/CrnqQAVmPW4OnZnR8BnDH2db4wZQpePzp/VfcJcRUFvYJW8SiUt9rvBj58XRHa9
edwMI6UXylh/o2UqPcTSTCsO19495X6PWCYpHsYBmnt97TfvnccsyJSrmcgGbHZQ
X5CKgf9/ngZmRMCEuaTRGRVw0rsHFJ/BjcrjHR1nqjtlEoW7wrikUNrGp5Ui4Fsa
iS4gkXQ9Xw9hTlKDPk/xbeli8dAjVsKJaiOOaMRoNST2q5vi1ION5ChXC1lsulB5
13gcPTmBTOzvbXBj8yecZ3O3X/I38iwOrvBCV8pPqz1Du8e1cXNxu8ywokJcdpTh
zgebcZ1wX7MAp/gmyik7L+uE7TUWgYp2hYFKQJwemxS2QdDFcfW031ApHXtvOV6Y
O6Puki6YNdL7u0SDFR9pZhy0KivXCvD3Aaw0DJpzOoEDPD8+ajLux/+j9YnV4dCZ
T/5C4XuY3ZPiBgCN2uXc1lFD+5IhsIJej8YZ37uGEjq9dnrLn5nZYJm4IeQuEUJ8
ZmqtDqBz+CKDi9D/mjw3f00XsQ7hvMgSh1a0hguJb5qh/NrO1LvEppC288aKo6iq
IDarsuSNty8f4f6n83/6OiRGBzUnyEtWxmORnR7GMChSx8nUe6qmJ+m/H67rO5Pf
qlOIU0YprdeTXa+yqnkEEUzAk/eJbzHF7bIGdrJ1tAXzAKmZxF3lCC1QC1qkG6m4
6fLPRKdU7LBnV0M72SGz+NUzJYFn24/d6XUwOO7GBcYnkn5bpvk713RBXgMp1iL7
bwYVUig2WQVS6LeBbN/fiybZUURcz2MrXENtHYMNkv/YyC1LW5goG7AVVRg+7reZ
Q6xKicp4lbz0xxT7SebYuhx/KRP+Yv7XbYasKSk8GaCWqmSsFlNxWkI+tgsxzmvy
o+YpzWes2FXhbIoIXN1atHGCzXA8zKpScgXImIkcWUst1jhhofyg62dYTxTYk4X9
qNagmb8dcptaKlkByR9TZ8Ogzwb2C7DtzlfA5Rfhi/1Xg3qcPYy0M/2WQHXqbN1W
orRu8oaSkm/4OvRY50nX1LdjbCEAh1ORvbSoS8590N+supvcLX7JhxW+c24X6kPP
uQ9zgjmxkDvvB0VOIOueYV44zFrq1HDrFqd+RPtHbTBKel3ixu2xvBiUPFmufyub
iCvmzYpYgSrQuA34hEYC2xkLJfv1Rl3vec4R0/dGvvcccMB0p7oUCznWVmK/Y8CQ
c2k23RmpNFrS8g1TchsLBQE3i3dLBWnrsCaJGPVafgCGO8R0WQRe3RSRkdT+0mkg
YYEReyTOkbI1dF2dQAvamq1+zj/XaTNgb5P88VbKGtgYrdvoW3IZBy7RgLxsWNoe
NaBjBbjjV3hPqiUxhqKtFb/gRx0nuorIS/5OZAZCtoCUDI8e24RuvlagY8wkCmdU
w8IUvtdR3WmaKRG4cEhOIQH+uVosos8txdlUEieLl96SpDdLhGIIQqtV/D7UC7IQ
aZqUbFQhqz0TQiwUZWux1TvtlIVMDPbBWoRX+D/TQx0GbXKCPPQ6oe+Rjjf4GmaB
z8kQHiiMWu1NiGV/wENoxKj3rELPkNmMQdVsXoNDH1v7TDWygCS3dItJPvLGs4Cp
Cdz7stO3GYNt3Zq/eLHfNXH/mO09cYsSfTmZhVZLb+zqUyM+hI7V1g0gRldaktul
6IxTamDB6BX0OxBzsLuw7f7mwwMRigEltztynWZiyd5PWjK08EwA2d/7PZLzmEmE
9vfvOgCTrL+ymfvFhjIL9kWoNxR1WMmkBzmwYoN34DhfIKwGCFzZ8R35DNLCJ3Ky
r/zI+tYf/GV9qJ0C8J8ZteNyTbvKgjd/maEB6KqyRzocOByAG1eW6df3SVEc57Tn
JkfPTGUxm7STtO7KhIpv+blbmXlO9QRtNYLNstNbQe9Fqrs87chfamxcTpcFOe71
czIN0o7dj9zuaDS/IAhfjIs0Bay6cyWovuaWYCKML9z8m1DntQekdtWd/ioU19Ui
1XoQqc9PJRU1IjnJngiFjD2OWwJWaiz/Rq3J+Ktjmn95YpUz+Qsw32feluPUG1fX
kYJBRNTE9eyME/xFDymnzjMzj2U8vDqzWLWaRq9Lxf4Ypv+o8UNji1TzKdJbZSOd
fRAhyxuVnk/rOR1+ED3SInr1laoxzk7iO6W1nPkO7CeCBLx37tFdB8k7TMWpe2bj
IXgYnLVJ+5sd0W4JBIIX7Gd3ENHH4NubyHbGCfv/njMZgH4wcC6G0HmNJuPx3cKK
DqdCoY74rtpTm5IV9CRO4Do2+l5PEwCbucyLgEa0lRTj1mYttijXq9HvU+EWvzku
piC15EzHdvbrjgKusrfGvYfXfhmpfj06OZEjTJRbZ1lF8jumU+qUO9C0yrbuYpRU
+YpcbKM6wFeaU74UH0Ea/wNKif2nVmQP0L5smXt1HKieoRbPHEdyz9czvhTQJacu
IoaADjdCRL5r2HW75Ual/OYgJQJJrK1+KAetQlqAvtOfFYiGolJOnr1FXuPuHzuV
HMiAWM6/aDG5sHheXgK7ZbJMZZrPbaJ/L5jgksoOZFfwkkTTgAyDRPzmYQX+zEWB
F1XTIIehYIkRDsUzaqZTnMoWwEuIDoTE0NcE4U81WdLfD2CC2olrHlBTHc6EEwaI
1h+Rqq7KutH8moRkQFuEX069xXR1yKraCTZf7tP1KmtbEnru4zo35Iied8+Lgo/9
XNXbIIXw4DSrPkO5HUuHXzLQMoej3eOqeh/qiwGHxCTHWfInMic5j/qLDmjbwLpG
4RK8p48Y6WtcLrCMBMApcn6g9i5eyyzC1/HoRuOowHKT+Y06h/Egn5r6d6+gs9JA
4zJBDSFJewlN0txZkVPJwom4AmvhFdyjd9cuaujLh/q/yBKmCFo3ZjOEdeFp/TtP
u4ehufTw+sCPxoI6nqcb4HtxK0Cw0RoxCKLfvtJWReDBYxMGJAuAy9cIoU6tcMYJ
sK2fI7rmG960p8SFZdUqhBB/hJvHwIoh51M7mUFcSGzfhgh4EYDFxC+Y+opluMhP
S0p4+IeD0fMvxvDgMjQ8C/TWd8Ss13iKzFIDn1Jjb6SJd5oQ9uuF+nCr3Mzimxxg
EhhiFlUEllp3Xrz0hEFi+Y5E/u9h+BHullF17mfEx47n00cBGAxQ1r2xXn+qZsUP
lN/39LfS57wqudcd5AUFzssnSzWi8OKIhQP/p8alcLEO6doZHLc4eMDXplVJ/kr9
H7BhNPCdYRYev3BEDI3NMSuQNO0MT8vv7JzDlQIne/erfkylHr60svIew0BvmbjG
T+slrherLpGy92L0xzFPXUrn/6/M7kqKt+h3mC5spBAMzixvm0ePZu3SiunEr8om
Mhi0zOJlwnoxeFgsLCUWyqsElT2u7Jeaxr0du0pAx00f0bbP7pzO+x+PI9vxlBAB
p1wbJXIM5sP3BU0vpWJ9AIvXwIhita4FD3JTl/My27XjqbJR1qXng20JKVh7XMYS
bY3SX495kuSq8ojn5tXb4CgRzrC3FBhhF0osFKHBUeEUDCmAX/7ojrBzcezygrUD
YDAYxU+uWvoPpUchuu5ej4c+6qHw7x4FTHcJ3Cw5f3E31oPvIbk4DDRoWyt62Ke3
D1GM4n/Kg+PhgIHqSl7Bs3KSXWOYVxStkEdkvl+BnuRIkY7P8Q8HDiVCdN6tXqgK
SkJ5IYJzbTMSHOQbhfZ5U7aRiV8zN/nrclb8H9tBxu6lTbCccEMNWD3Yg+Yhy0YC
RYCpwz2TRltyNMNv1x4XbQa1At3g1J8OpObkRjo9Kfu/xwrsxv7dRNheQ1UkRAyh
ipgVrSwJPka5HSHOvVtnlt8iGuTHZaJUhNlOBseh6R5Xhv4tmeFkCUWOJjD7hEsp
6duzb1P1SNwwC4AVTqHhwIqztyZYy3Uux06U8van+41g4mWX7MqVORbFJecEAGJX
WfuRTBaRFqaH2WYuafUZqeM9sKFPtyrERTw0XYjpkgXoKu6kPJSPttzpqpPfCCoG
OXZc3fBbuuAt0EBSryb774jmTJqMmZw4sXykfsEFOv9PtsGXxURl/+l0ZA5xns5R
+IxLzy+Bkczm8DqcWVbCRw19nvNvqBLM8MidUPWUV/n+34p6+uLQeDkdVurIVTOO
HsoGbpCRSVw/PG98RXcs2koSJRFUXoXIX1RgZsqpr4TiWcWkhPOEsN9q4Nw76v3X
2OvDaUqzql38p6bHUyHKTqeONqAx/kX5tD563jhSaNKbhuD+fVHVF8Z5lh5RQaia
50NbLzejqVcdk0wmP9EPDGPAK6xCfGNDvlGWBX0R1CdD+awQcU1tPm9nLm7HkjUC
bYGvnec8b9iONCaXbi0U3nsEHKqXkdVB7zYWM+zGHYVnl1ft6qg5gFsaFTBxQFAm
QPi4yD+3PflZo20R040dKrx5EZ+x47Wx4BBNiZ++HGE/1X0CA07N9wcsbN70i7TZ
btASowbPfQL0d3DWLnOM9DrD9f3k3tRzMKI1PC+PysYOsDWJpvlPVHnASLh5K6LL
9oFhnPS+4JUfnentTzBY8gU/lTqVwGOSxJviDDwueBqRFfE4Kx+QkNp51+t5siNA
kU1C2n/tjBbplauPyxrRiemVnrqhUNZnGHOvLHANmtGRG4W5UvLITGhAu/zhlfx7
8Csv4znFmAxvP95Th7ZioNOHkmNqLbh0fsZ7CbMNT6f12XSrhWjFo00KkkkPXpF8
bFnp6FS9nuRIvggZ/G3fd/1iWXC4QkUTYC2Ji4IXvpg+3w7lo4OcmLpcRhVf2CpA
mEajU8KZzG3KUdLAE7yYTHeISI7AnaLA841IOyV8GmbN9EwTbAo8z/lg/AIoZNMf
kF6Bg15Esf1X8zJxvM5HtGdrvqnZIsPGhA9bBNF9njBCguPufCsZjizwTLnkBIOu
Temlk1KAm177U20+JjoBoDhzbg+jfod1WOga/ecCY+X6RGtVTkc+sMC0y++oE7tw
uuFb6sm0wJ77v89v6Yrat0JyB9LSKxboHhtRjcezqitwR0J1RTV0GjJFZ36lTrj5
Ox2hQA+bKVb1e9ZAQpk+3ApXAn8UBXYZQZIizriT9vClSX+e9z9jnrn+Zf9dfhSa
OTUk1OFFYex9o9wOLelsw9/Iv8CSGxpfeaJ9W46w+N1ZJWRk2oDAcvI4AgkSJ6Kb
8Oz/8lUiW5H6mw19Y2uufWibAeQXT10Ar9bf7+x9yifFrhCCD41JkGlZ4GgIlH8m
sog6W2RypLmOBVTGzF38pgI/SC09RToPEl676V4zyRdAyvFjvszArk+06xtVHRji
5+F7o8dKGp2Lii9NxnFd07Y7xYc7FD8tuUKO8Ww/IiQVJUQWBEpQM1YIeuC2b7SR
I3vlyc2xbFjQfBIMYzgLCcanh5YH5ceacObv8cFluSaZZJwPla/K6H38Cx4Th8Ip
lxtqDFg6Hm/iz90iGGuAeTJdvkHfyPzt5OuhDjArNvLn56+YBtYM3vvrZ2mrslcI
sN65CXRuosKlrUhzNrvPSvhtIC2LgZPNEqYt3OwwyQluXcqzabUSvrs4JHLq9GOX
naHO0HC5XOunaf5WLtnGyUIOTMXr2s5G7/3FgB01isVK5jceD2arED43YNrSoCXo
pn4mIO/+RtwS6ebkuB520Ulm8rjLe/X0kBGr2BddYSw/Ec8APAIjTQf+QJoLVAWF
3mn6sauMFWIunM1dubUGmhWgH2Jbza3JET0I+MdxjGSa907+ZwNqqA09mJbnT3XF
w/LEno1KQCiw225Miv1gLpDQPRDWbYEY3iszj2sZOhmQp4id7s4U6Bk+K1wtauUH
8sj6dZ/OeBj+9qCHn2y6rbLOng2kY1lTHwxLmY31QgOu8Zt0r92MDKUto7Y4YJod
LoeSJlXBORm8HBkKzE7ippIzIHv+d9FJXmkCGvBdNpQ6UkuNUdzsNmR4gufX+4bX
FjN9n5aJ1aMmr9+qJrvRxPn6GMWvGgzrTIeN1plFerGwd99wXpReyP286j35PCzE
h2BAVc6YsT632mlz7Z10ZCKare7CM1L+5a8oNswu/YksDifSqFr7X+lKjvWU149s
jjkFaq+5IcM2uq6zDFxSHBvyzArNMSOB3YQXdrLJHfHwHfAH3cfk531NSeI4AGf8
VI0Cp41gNar1I2YZErgIeI/9dV2/F5d9nboXtO0MZP38/Y0ZtYh+nop2rxv02+44
oxyRWjxNvvLHhW9Sljh//rrNX1ORwozVX6ziCuW42QjsVBl8o3clHbKvMqaD0/7C
NRLKuG2mVCHjcfyu/ObwlwHKyEGKNaRUa+bdfhBZH1tS+nfrHUVvsDCBNJ32srcY
hw+QSiSh4/jKzS4zW1mqbRgvV6h+bIFAhct9QUaSyvX1fdkPrR04lA7/9aVeOUqQ
I+mlJM/TNz7yWEg/BHGzCNCe/rFWM30PibTeiRADOnOV6zavWgeg/vnaLvxbFYos
CNk8hNVHStslYSqeWGCwtTBLIkZ7HEvYljfgDJtsiw7qT/QlcDfvtR6+rNuJXm6G
n2bQSjPvTkyGT3lQHXkJEOuLhK+hTMnn8vrE/U2JV3zDqt4BNP+0JxVQXkQn4DFt
tf7oW7KeHeKvG+vtU5m7n8Tty64u8gxRP1g4QKXxI+KuXHx5/JeSzUx0VU16l7oY
7+0TBfie1sskQyoZ+sZXcC1pWp+Oyx3I5pxO2k/asnUjkB4TLjgElBlAs/nGRMHR
0WpgLwzWBpMqbD6RIiLj9md4cgwd/BwxP786bFwqwmdDmlcibGPA8Ud9AYnZXcpx
yJD4N0tqgikx9ZEQchCjs2TlD5ZTmEtCJSb8yYkKyHjSO8odtd06EikOr15FgCgJ
eq7RvRVta4qGp7CcvY5JdkaZRDsukFA2lKobY2J2TldT+k1aYNjEiFJCPh+ATkis
eavDAh3GzP6me8+Wzw7whqcX/9PzH+qxy7owf3aUdlFoV7lI+RCivK1umXOsKQ8V
9+oznakBCOsNwCEMhNaLPA2Wk8TUDYzlB9d0KtRBZ+fWx6bV14wdYtRRnXERyai2
R+BTicoldd3KANeGDw4EbBI8a0O41zEKvXy+ozooVmQaDbmoeHxejl0/E2uo9lEC
hGpH4RTCSfGOHWG5X0K2p2uPSOLzoVnjG19/PJJDrg7SPUzVhFJxaCuhupjF/AtQ
Mqgkep+RrPsEmBI/h9UXSwBrSV+iXDyTJ5HIrxRxmwu3ppR9CcGF/bcTrRKWeje4
7mkyDfgmRsMrpNdvGWqO1WFI6sMLtVdUMHPDEWx7ulWUo6pAMbEKze7s7HqXi3AR
KTuVAmqSY+c2L8eGheUTiciMiPMkrZvTuH8/Gdjz2p1KdJjukZfn5jQip5SCkDmE
sRVpTsd1kYlLxDirJqv3KqIUA0zQCLWDwCNF2SbM7PBGPC6QHSuHsQz8I67iZKbI
RH6EXY4QO/d7zEwXyAiinK6F/xBVz0p3z/qciiuzTiI=
`protect end_protected