`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
hVdJHWSfELCmA4ds+csnOQAALbB3ps7EiTSHEDd//nts1r+JQrRE4d3bDPRJpiX2
Sl8d+xAK9BIi4i+3ruAzYvB6kuD7r+gs02Jsvd/1kn7JYK4xBxCjtdDFjVHOTEl1
sSh1oNiYUwLuwR1yKfP+xBhqxD2Dv6pCKhH1NdGilpJQ6cvivGkSunAu0tzP76T0
4x1pB179E7uIeRplfHWX03KzEBF+eVtfgXVp2W1BGjfAe43y1pCvNYZOh1+TY62g
EgAFgbo7pAujZxZy/YSiZjUr2mGp7o83qMXyusx8+rQ41D3X6rxfuP0RiId2pOpC
6oq5Dfkx04a1dk4s8w8cVg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="Sm9DkM+kBxuxXCFA+l3fFkxuSWV4xqRc4Nn7Ji3ukao="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
m2emGBqRy4AuduN4dffN8194qYvc9UXRqiQc56IrQYMiIVQPyh59I8SYabcDdspI
7AFHnvKD5YaF6tQfxWm+mlcmMEk2Y//aUjxeiGGs+RkKgbHitJF/K7nqg1dmKvDg
a/GaBCq4Bqh0EehlN4ntP5HxM4qcvSfh5m/Coe3drc4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uG91daMWA1mGkhgP3oZKMYye3UAomMWgG80HuuXg2E0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 27696 )
`protect data_block
c9NqBF2D1wSep1rW7utzHsk2j40aow1MnrccxUTvKej2Q1cyeDDbgAml4eTSXI8z
QYgCADtWi7S8BeChdv4B2VxKcS7CMq/DaQrOy1MKTfT0ctZFMgnfJn1i3L7BUl/I
j9FpoH99wcKG2QKUQxXH/giA/GS1rc/f9GN27YZWtTl+KnoqBaXQpHIcQJ5e7xoW
qb6WYC+bKE3r4bBpA2iEgtf6KRzpRScHPr3fSKJm3s/lHul15Zx/HOoI40yOedSK
N6hVrbRS5dLA7Di01ZAZyeqID9Xm5cSoUqeY7R4sGBBAuxJpc1T7n/s+6hKf7VF5
iPnLLDiKvNmh0WQSr7vW3llVaqGQ/KHOMHD0Dp5WSb+Tm+OihuDK6P07/b1eSgCK
s49AHTb33U8TbxUdYbdLXuE3b0sqDTigLGM55X6IcjuBFAAVDL50He2v0VMHSxw+
1u6hMoZ4Ekk20Cau4RLDwhOQdvVLUUaqRgYVjbiqZCScObE2TSILRux7CCxTx008
ugXUUnB/vywpYbz8VxE5mxa0SJSgs22dyiPjIp/7FBLBiLuee9PTqFEQMobkZzFf
vgEFUZS9MBjwGNZjQmqbIZT6Zk8HRZGwYLNORrjXejk4talu6utlj/FTx4/OfDUn
HftezfG43N1uVVT+wjvmFrgaXU9nTGHlrMpO/lZ1LBlJwylQsmJGxdJ5PI1aDltP
z4NHY1mZd2cKhzHrhSLr5NgFPXurtgMHKRmPmOnQqHdnWUIRs2qC+EJIqJGsiw1a
PhDxA0BLNsc/xrWXO50YOZqGnaTUYMmFf8V2OYs9nJlGiv7pO//qxZ5Dq2w+S4K8
XlRmbeahMabUER7V9/CDk+JWwab/LBjL5H4atj990acGy8YNopJpzh5lVk9HAS0c
uEAFKWIDnSZni1JQkdMe2MTQuUxESxvzu2xNH8SZ3hm+ecxLzoTD7hiDwuC7+v7q
xMS9SHyeRhEToz9dz/IAsQYzB2CtNy3SvxloNsN0inkj0JMoWBJm5n10AGFaPZdE
8pYBq1i/+PnEeTpMjIVYcjh7OK3FqQeUoIIcmRu8MshHY1HqEaBrgwd8gCgBjoiZ
xezi5PwfNzcCDvVRU0EWPkFa5jQs7QM3w4ZfLAmQ8Bpo0i/MAEsQp3lEjhvveh+g
zN7PkGmO12+zfigv9MASR4+2NbtSPk4boJOUuenn8c1+4wOjHahkD3Jo/UcbUBYi
QI2pkkJdq0TAQzAJdxdflNXnWyZngHa264U0qEFTrImsdmJwnBU+7QEheDgVhlqG
UsAcyNjY4AsY+ZBSMplVzBDdVj4kDTWXPypEnAE0Pi1gqQN+fxPyqWqibvpanksA
MzcP2aPWtjQpXknDHwKm4WxU72uQjRhqBSmqXAIu6MoPmoLgImjIPGlcsZBkpt4/
3PFNZa6OQl2nrbVHfmWItdL56/uPvuShXvBku+AEDm/+u71IWoUNY7fjCIhP9PLT
xfAx7tFuUkuIgmltMFwqqS5x3MeafMPzNjBczCNDyHW/cb+uxvTR7dXHRF/QW7+z
rjzUH2nfRG6aFlEr9AQzfcqxOR4MbzY0QsAzLgLNOWks7cwFjxgcV7tSwmjK0A77
q5cdMiiTz4+4nkrZL4mxFQAE9P3yaL0pcC+FACZhk2U1E4J8uTFwSiW6XIjTFNzZ
/CmYPMm8TRkzb7yw9GqfC8U522hS5uhRJytjjHXbzuizpgmktq7HS+IM9XiDsQWg
tyz6ZumLFWxk4rgcSGVl7qgIvxgC5BOKnD1J58zdRsapWdolMgP97Z3aGIyVCQvU
XQa6mfN/2trjUN1b3bC/HXMW7zCM0gsYe5wuEKQUgJHxjethMH6EQR7gVZ3N5oz6
TR1a14x71AVFjh+UozYDucV5rISUkWj4dgMIpLeWVrjscfRiyH6btJe7HTja/voq
Rtma7NcL5EpCWF1hDUZu3Fp/SZsK0Lia5o35YmWV3VwoGshCZ3uUbunZHS0dYrYr
z67fx9VQN4/hRbJhTE6lfBFI83Ircq1EgmjelsMFrnLuqBwh/PeWoHaAjxaUX5XL
OkpLqjrCfhupm/hPgSN8+9y1gXSett3FVzqQQ1PhbgKmfh1U85ETK1Bz+lqAs0Od
K7x6j2d3qlhCxUmiTYbRMX89sMJhh5AA60IeBFX+j27cxO0p8r6VB2AKjV1IpFkd
vkT8eu27ZdeZRuinDeAwYk1fgBhg3nQob5dSDM4QIe/TLLAwBstWEc0iHDNP2Jkt
XFaRQhyk4yGs2bgNePLDWK7GTDcm2UsmG+5K6S17+QOStFeS3kdxycfDrIO0rdS0
lEyr9PnZFcRaiw4kLy2/yeL3ykpGkwZcGSRNh4kxMLTxo80ukpIFv13wqJSqyn2R
V5f9OvmLmgCnODTqqsqLHXT27aPcplYIa7N9Yo1rKvnmKTeNrJHloEqf2GyejBh3
+K2wcUjtxbq4OVcTguvx7UaHCKFzUxiSnkSZGEqfX+b4q2TdUeh2LK5KsOYaqmg2
2NDhWGv7LVS5dLniq79HuDyiQcJ/6oA9ZX+YwV4Rrbft/GHGFJDW6QgHaC+bGTT7
nS3cOW+j7X4BbokKv3LLFWp7//uJ52p01Z/IIO46yOn3SITPfxCXsOPidHNylMe6
dRs7n5rRFZUcMwzUcYZwoFWqZ6TVL0QmtBcsHCOhKT45h3COyhcBqZgAEMGBvlfv
KwXsDsnbt8bxrJ9dIfUhsJDYIkM+TQb6Q9k0m7bWOtxYqJp7FY0bJ/SEiJt3vCeV
SzQoXrVx9TGBQTei64fc59Srvmv9HCtm650kkcRopEzyTum02q2a9P7yVlPiTPg2
3i6XiZRPCRUXpk2a4U5S9C9C7hIRvuCK72oqpo/lHiwaXKBpBg3Rp+AnqUavgeub
9oFL5TXmj3lMmguyTF1s9FsC47oCD/bVNflaCGvSxvwe5gS1WV9/a+4yjuRX0QfL
h9Fjria36oPIEbRWu5EbsrkqJdzxiPenVna0A9aAAmtxZTSFvcfg7RSa0Jpdkz9p
r7HLCDmbByAed6S1TDVjs+YwP6npqqy0YAwv8BAz+QB0iIi31URPIe+fZ8ajRNZ9
RHgAvbzU9VISn2p8Jmv4MRVmf6WDKM2vECOy+PiDLubBxmCj3dtqQJZKJNiiAdvo
+rc5yW7D8909xS2QAwu2WlrOAp4fNklSg3Afdv+/Gvtgg9UKBvz36JRWeF6ORR9C
ba+ex6qW9qR6PsFdpzUcQmbaDMsJEdXIvr4Dv4a/uNTKkJQB2Ed5/lFlH3waVaHK
lj7hTwZPOaaVfftcg7p22nv3Q+SqEoKPjQnHVIRxs9UjoJwQbEG4ijmZPKunRSCY
pOqIxWZjKzbEOfKPygm59wf5sLNuciwbsSKdNE0OQKKiSYT+9KLhzejusPE54aKr
JrHWACAy+9GyR1EX21Uaqa2PnmF1m3rgzv3YP3Zg4QAhoSZi/czCQfJwCocQ1vIT
9KmVABpFNDK4MgkKyvF/aFvM5csQkoFy9AFBuRRYuK+d5MU96bpe2VoZxmeFXlRQ
SQspCEQBmZ0NEdD7Vqf1r8QFzC3eIUW71DfnQQu5w8zWNnAlpJgxk1Q4OrKr862x
/yYA8gtSoZ67IMM4ov/TEh7KdezQY5YX2Uub5IjZprNb0S5PZuleIdNSHhJJnpdo
zyBv+cxlVper5AWUWnCjlyQxwGdvP41lPXSpubKix2gvTuT4rPm3o7vTJdZVQg5e
sbhgETqSlyLn5HbA0EweRAuEI7Pi9MWID3KqE9jjkciUTo3N5LHF9m3LMxrU3gh3
HgAwCTlz0lYcSJfRk54ymEWSvOv+5HFfdziVXGhDoxE/Q3j5yBLPBasywcSReZV/
W/vscBoZft9f9Vux+w/zndkSvhZ2V3xVh0sKi895XmhwzHa8dy+EwUPEKjPVVWeS
5v9HALHr9LVIsIDP4Qj04+D1LJJSCeQd4s6xGCly3RD7GTEQMkvKScOREhsF/pA5
f35ugZ3rfAjT583Rv3ITleeRijpE+pDOWreX4R4w9+zewqEbW1KBUjMIQO+SkkoW
oLpEsOBLokZ8ThXeHl0Gaqy/sVi3a42Utq76IOH2T9M0hrZSdXW2nez7SWW/+CNq
hL3azfop1Ey60NVw52iWEqeHZ0J0NNtq2wppaLlHONNJBZAlnlBNQ48MvkMRIm6p
1Tj9ZFCmyGEFJ6NdPYQnmjUhE21B2C41UrQHLiEbO6Hcp138sJZFLaawovn0Dd9K
72AZ2rDm8esd5QZH0xN22fTDmzjSMrz0oaLO/nYC1bMRvJnh5/rGo5JMNPt9f02e
iGo6cO6/dkLhn6jHSfcDb5n3DU425L+RPzptquCB5PzaijBQ770eLr2KGG9gSJeZ
b+gSjI5xhdNq+8w13+8NDfe1oemM7jrgkbkvs0bDIlQZQPnfTQgKkmHKmlRLSZKh
dWcyNkyMpMNRmgJhJCXP8U3x5+4KM5u2t8keHi1GhZD1054XJWlQkaDP0j695llc
Re4RZo9mVmQ5zBwiRcB9OaSygIiE9nkAbUwTyv1tlMen1TzBwgDg9Bgl3LVZ5kpb
S0JjA3hW/bxr2jpjo7DUgANoSxKdg7cPwqzFj9aLwXIQm5ynMT5nbqnOznrUU1DX
bBt7Pwdm8KFptyutt/omj55ZsvDjkWi/8MlfosUdRy61ZqrHbtfY2zEnF3Etq0fk
D9KJdOJZKiMjXOVTDjGCizZ9qK1qNqkvbOKZWYRXaEKqkGOfslvp58ZmoQRA0W4G
SL8rY/qmv3QCmGvkDesiNqxtT4aTBPh2M3CuIXV2YGm8hx31IIMtx2Y6M7gDYXfT
m9j2U/0clIccuCksEHpo/FSj+M6xHzdYSueABTGkxc+82L6ErhWgC2Vax5Z9gAUZ
bfQkIqFfpd+D0OzVUvBbdTqkbYAt5a2giPR9ODEDiUIhiYFYun834O7jAfM9imFy
E5oevKegVcjZ+rVig73zXaTHJQmxHL0ipH3Brnk/Pb42Ig71vL0E27avO7dXcg5V
cc9ElNgipsV8GJeiReTTLc0qDR90UtWGgKpaClswGUUpie/I0FCRUzE4hlCmCNLd
Nre12r8Oz46x+0E56lTFKuF51MApSmeWZQqltDDuv4H234AcQLuxuHw3rbd9Qw80
yB7jBs6j6PWVsGQV3zbeKV2zDZhDW8AP9BfV6KfvSQP9PxvicePK+6tYbrIq3i7m
9YZbMES8UJ1wwvHMT+FUe5ofjibAJvbEuJO6Z8WtkvNeorHauG9Pxd5sFkjNPOXF
IjF8k+VzsHz9N6m3GJ33BPm53nDSyCFODTRSiXBy7s8ThXE5Sg/WAp8jZ6RqulKH
Cr1zm2aOZmBXboEg3JrfBBYn3/td4+HLAhvxdGmLDqvvF6ukChgTGkDVWUa46S00
OTH42Ca2av5FoLNxms4vdEfRvSwim5kw6mf3GcCkNBJmgwXwJrvV/YqwieRBMyMF
7a/baFIvaBk8TBj7Pb4hQEixOtrv+/jMe2JacxJ6qwmOTer1e1ZtAuMrx2sXNJrE
K36qUx5q3RJ/HXjant8wvv6ZuzNltz0k9m4rXsyQ5ZLpXvgubZN08uksI+X3Zy3E
+0Kmwp3GPAauCXNt0zLp/oZq1dwi3Sk05b3LyGJagrMkHrt6maJqu9Ob6npbesm8
zwBqWXM1Sz/osrjXmzVOcKRUWdmmXVwWtzoE/4arIE0PSphqpIzaf9TNzsQ7cgU+
DSoQSzipSfL1jtaXRkvUqrw86sLdK5dDxZLb51tRREW/+lNKE5/hVuQZMgrF21Rf
QP8uc7MoJhpJXT/IZOBeWqif9uN/05jQgazeNJnyZ008lxNtMY62uWIv1ws+aE7b
NLhFrOK3ou+OvGk6lOUu9TwfBP6eRiaTCLKNmmihZOcEoftKTkCvJpZuncBn0pUz
OJJRkGOv0q4omKR/825KXpNzgAtA0kr8wqpdnzA5vwU1Wns4dHgzoGq4ea2x8HXf
LzsptLZbAXkU/sIqm7lqlHrLGb8ZOv8+vb9OiA4D+oDLZHgHzWQFmduCuE121p7x
UuPlh/wmMJ4cjhNmjbMFscBdk6Mvt2RPuIkBBOs7VO2VdDJIE/LXR1y/yi3y+KY1
V0BoubzC+0BvjndaicccOTf3G5MLa0LSgtXK47vvVx7n51YYjTry5HYJuhI0AuBg
CCetG8TpNcGbCZZADeNKgZfA4CaM3SRRiff+zKwPRKQ7oeKa4Vm4Mhqlmftj3zQ5
/pBvK7KHnSG4cBQQpN9Fux+cVyKXfvkGTvk5SqqQW5XjgEPMDo0mZy8+lLFDC23B
DEd4y5NZgQl2ss+pTeepnr6QEckKop7LawAIYALoI5dPrSd8zQOCpD5FDkaiGDKA
qRhsdLlQ20aFFRsQG96JYeG5sZkGAaN9oXP7Cf+b8GRJzQonTR5kZ8OxuFGOYAQE
vtl3hbDRFxsPK0trtv9dZP+ilKWgendgtRZHdxj5NgPVF/ZB3zFXkXHljvOqyb01
eN229S2L7+zPTcBUL6quFMd1orTyFm60Gqx0c1yaXUabB7zcy49R/NN/+IqBeSj9
AQBLH9WZ/4nIdbJP2rIHqPRHk7FbliLxF1XD41LBpQ393YsuCxxaT0vpF8jPGILn
f/Wh4z836clAut/D0qu4l25eyYYLy5WSRBaD3HXZMU4A+U+jIEC+L3qmNLAJtere
YlDbd+/rf6BLkc5GHJRA2hZ5ErPd6YfyxgmXfMA+8QmyEOn4FBX2BhtxK2PrJgGT
EpBYwvz3hIiqUpoAPTFYjfdhEyFhHAv+gwnR5/Xujxic/UXGJkQwF8imZY3dLmNu
fF4wWoPBl7/zEC6tWJevEhP8whOo33ujYnp2fRbuaHN8BcGLF6VTQymgMpiRI8N0
LA6m/2wFQMwCyBobkNPLJppWOBauuhA3G/UtRu4T4XjBNLHPKSDmADvG820RvzMV
uuOf2lsPYoKQ3x6DHbpkqbrNw0u/u6juygYTKVxAGQTne/2qBUoI6phi3+nrfKmk
OWp6Gytg7fS4KnaVZh5vfwjCfQ+y+V/r0UdHtPv/RPFYC5aAJb6I4ZEEXwBQ3FU+
gYW5MFiYcjLEAnYY/iwNGtvavKUSOd5R4bEeQoV+VO+aTgjijdzIVaukDyO7FpVL
OJsxyMqK4+/aFYR10yZK70RvRK74sKDYohmmaQj7u7B1VRsUTll8eYNJyIM9yiuy
NhChCHADEyyKLrIvvg6Hk70CT6ipk3JlZ4kXyV/gGcMQu7f8WNyHJIKuUaOd6kmJ
iRGKuWxyAGWnjXFJys1CiHdameEDmmxe8nZ68yp9WS8n4oLDPo2yPKfeYlAzM5xf
KcgQY3fnEG/7dorjh7qcei4/SxdYLp+imi6w2YJ8jXFynF6CzDmHX9fbb5XY33Kl
8YcQFmwZ/qKuBeVNW98t2AyMIVUjDFyle6iRoZxAqeB1MgAVsnCysYYbfg04TGmg
MKzJyh71q3ezo7glef4V9zZUB1c+y0X3iUUoVJf+VX0+0m7bLgiw2C+IyRG6W68G
O2tkB2BkWJZFV/F1jnH1BU1ZaH+WjgUmMDGNg87iv8WSiR4WpK43ZPR1RnEIPyCq
Lh+C5nQ18wDBb3Ocpj/xHot0OJhEQKxdy6cTnFzD4xe1fJCS/sffs2V+F4IJ+sgJ
5oz7rRUy/b+ACfy7GX0M2D1C4PQIt/orbU7NvA0r05ttEZ3Yb+fNPiS95Ug/1LAg
9sd0b2lZ+E9Y26MTj9AX3a39lFFaQ8/M2HK827mJ0BBINSTUcIIEuj7YESMNaj2M
w/CxMp8arrTUtPC3X/kpxMHbr4juAzFHCiyfAIq1SgGQCOMNC2k8EqDQV6hZ7bE4
oZkru572hlbGgh9KGFwN/Ue2QTK+1kmC5/x7suoNry4ciLECfEjXcTP15ljmi0Tb
gDxhsBYHFwFtfpHh9RGYNDYPDAangBDXgf6dnFAxgMdUNdqScxAFB1kT9OTylzl8
a5ykQs75nMeNCSuXKdgRpW9zVwvElyb6DOHDcNHkQvM1GKGyOZFI0CohMeWVCqzp
d7L7OOhiG4Pmq3X3YZYazDedPsTq6n3G/mpfJ94ygMDQin1tfVoB0Sq4ipDB+6/k
qdT4a4uyqn1YxVOVcmZdrxkW4nNgxYKUkMwO44Ds+djfsKCHtEJIX46jrYf7yD2E
rHhNOkFfaVyp5sfaoYeJVnpioB3vQiVwHNnzcZqkYYzItTbZAeHcba9AkJGOA1xQ
R1Yfn4LRLDXtMhbGSW1ygBKFhMbl22meCZhyKI9zi1f0ET9PaVD/FBmZZ1tjHckc
V4W+bWt+EHcrrg7sMppsqtuZniTIv3Abse6kC5Zck5HntzLdPGNyV7rfQ1ND1Ccr
dy4QpsyRyOgCyIDRVUUT2JLczi7JGDS4Kur/q9KwmX8htInAUt7d0U7GEdafFFXt
ObEmCNvcncH4NvfPrcrYLOgDxWTP2QAj0h5jt21Tsdf4O1334Jdegtb9ijgCdJQm
4X6ZEqlRn2uyMyQxf5IhfNMjwIvx+F20VukWdEmqNfz52y9v3QI/ZgtbASd9Kqsp
J+9UQ32QBUcYr16bmu86EUBlaksTk8Up82O16PC8LSdeipMLfZj4It3kcTPRLYrK
vECJyEN9Sg1ZwUCeixIuc5Trw2qryIJLEQfqavXmhses7WUYR1goDhYEW50tvT5N
NRx1XerT1caKyVplkO04GUuIdWEyxNje6iY62m801oMC117yEGXxroLNMb1/nxB+
K6Wvkthjua1qjuu3SByaHYANCGaMcdc9hBySSyS2imnkqJ1Sbo+LSVBjz/xlvBeI
6MC2TwJI4quxuq9RHRl3QQe+N94WUzDE8DSRi82nxZS2WCieJytpfeO+NUpyf1y5
Bb8JtdmfNhTXK5NqsaY0Idu3yMD6qgIuf2lc7DmKezgw1qLpEyXiNva22n/s/DQK
ILyBSlM4lOEzmYQyyyiSs4Uq/n4kAP6InDStS1/UgEcoRWPu9Yy5qRLtxpKOPS5T
v3u/63RVuQFe4gucUSf+w0CKulfW/GR1CE1nyFK9j1eBO/IRf0rGjwe8URfV3n9F
Hq/01ZXVoxdpK+h3WmzHwBKyjnrvkm6tquHwt/5PyoRk767IFBDoNW6ZYtmaXZxO
8+yLHqZQqgLlTeozusPwxSG3M+Bz+9qeGQ5F0zZqJlyoku262p6R3Ull73DlJR2U
X1s58GMdjuVc5xd58+UOlXYHwYWUDbq6io1FBoJDOkf3gGZeAGCNWR5U9ecdCkiS
gxmqWmrqGtqH0ar6r/osu2fpKnfEceiB7QO4fFjj38uXXj6oJtAuuBxjilWxrBpf
ynyozXt6EsgFweYNmhwTULd36fUc9weHvfeDWo0TnklMAz7ZeIIROXioctZGUBop
3RvTUK2+ZjWxHm/zHESZvIbOwrQ7MjHjRBAW18eJdJBY+joIocR/aWBLMBkzyBS/
qnIPRhTG1tlu2lxhHHgMnc1s15dRi3vSPFB2GHfzLr2S6ONqcSI7CcEZfgpkTY6z
VOTbQDH23AkhCbAVsynfOK/soq4pVA/qPbVsrDn1HPb6JfwDAFHoN9gAYL8tyI26
HNCqvGX6Lxw7TnhT3fopFj1Zn0GkPyhbhfeVz7t/qBBhioI1KKHIJdwyMpmVU6ND
I8MJuYsE0cMomdKj+dzBnR6JtgjJRVZas+93LKf1XFropyEdO/vBDqRd6QuRkRb0
FmsCnNp8M4xEb4CFGKKefA/tqVCuqTd/wwn2dG05P0AkbYvgIBe7YgpnZbJITFJA
flTWqpGf5d/1zCfParIwN8D3auS4lGAiiFjU32EIimJ6zAPo21zf9FkQ/OhhYuRr
PH5aFnS4YIuS72HU52j5tRFSe9lGRB1W99yCsrGZmXDAhwnRUR7FXKMnyq5i8tbr
NGqAylhM8Tqa1Mmx4GMAEqv5QaaEHHOv+OLR4Lwl6HQ8jfYY6w+3Zn9LlRLtFNj2
z4E/uJ/M3lbGJFfKvghDj5yBQzPoiDbOP2mTvbBSuRjHn8jEoNaXMklpICmao9Va
nM2SmpmW7LYwD0M/RHGI7sSaK/F+rx1C7ExEB7zp+VImSzts5yIrGJb2clJXZCs3
+3EljGB3VX3cC16tk78Sh5WE9JEuMpMVNqbhThwK/6OS4Pm1RjADP/+U+NErySpl
FJyaja6ZAACPyJitSqj5V/DMSc12y+c0ZQzwHcg1Qy9PqtUFUSnxMG0TA6apDYb2
tEFdE293c4JsNj7a2kymu8M5LqSp5W+SXgZgHi90JtbiDznMqfrrLFuR8rbwGgQS
LgPz3Gmdq2tL6CPFzFc8bzUl+VrXbQ1+x0hNr0c/1NrKmJYGfldCsUvaHENObHvs
xqNX/zVineTGh8xWOtirZRNJF3tZd4Gzino6T+0yLA0hidbk1fyr6s1yX2McJiVc
3s408xTN6wZLunYVqa+UNbnT9E7hekPZn6I6/tXGXW8SRST5U/Ms0e7s47Rf7FcT
47qc3gx3i1EyE8dN9OXjXuxsOUNCvywKXv7ZinHftag8vfBYVED3kiVl49aj1095
QtvUo1TA9S1JSJLerMMv3/LmOCDfjF0YV4GuN3hZPltNUah7H6gfzdLX/30QmeW9
Q66a59nAxm+4uD715EuQ8B/jFPPMQWd2UgU25W8UIUMQqSWEGOKx0yAFHtzvKE7A
FNvDHZkfVikuse3bxjsU0V11uh6c+H/UTDV5tZR+Wth5kJMZh8VyEJQeK0erTgjZ
k7O5quj5HgdHEGpkrcgdfUcWdDWgIxenfQGdC54CjocB4CzNxSgvB8VLT20Fz2sd
PDtytk/HL+LAwE6kI8g1ItaC80FP4/d+Bs6tnLpeceojYNahyEjPcDTSEYYA4Ebx
FOvh4flW+JsbLtQANfYx7v+Hp2fM3mChHdbOFnytkQiZ3BKTAOwOlkP53Ue47fuF
rVEGSMM15Qaia1wSy6vrVUcoGwi0siLqeF2EMiusYPofrXXwvvshN18+lIo65jvB
gQR/C5cinBREDUdyrY26Ps6buBTISJLp/WBKOWDd/wY1boXQSJS/T9wy4AglbFho
EpIia3dFqSC5rShTvnfluHXy3FDFonSe1+um1r5mHNI/WTXQ/2NhgfFaLQnhfA9Z
dD1cOsyJUyy0Ew0s+5vKtvi1Gns9WJFzqBehm7Jh0wX5chDZ1P/bVlzcLY3Fqi2m
pMsSIE9sH8P1/pFPC0a9rN8Ozg+y+XfdtScOySeA2hbMGjnoOj8FQnVirRpYyF93
FUwrTgw2MgS9HrvcyXyQ9VRZEddv+ubmXNq9izjbQGLYMMqZiymSrbxLZnmMMwD/
qQ1oftPCHrAFLOVKcu13wLRU4qMkkHhzC3uG0h6yeCWa+Lukitd7/ADxH38127Wf
A4BxBBSAKjjpx7lnBIQMRQWmSJCC/ggsf4Db/y1UfYukN+l39znFuzxzu/peyW6o
UBT5DNHTqjVn6e3k1boRfvuzE/Fz8g/m9nJfX4Qg/rs0biszGxpJJVjHJ8w0SWm0
yVp0jSejCeAGKwRUp5Lem6wTti4I3in8dRUhkUjhVYfUaCjxGT2tLo9fOeSYocMN
lt9w/JBTQ7WyMsG+8eKACEoWz3ED8LTzv/jrXRpJBLo8ljZWlpQC/xhGYVanL5V3
ijbSe2m2DqNlPwuoSs8I+S5m0dhEW0krKGrPk85TLKCKri4F0h4CbYnSUI7CFS02
T1KYdZ++/RnSRHvDLeTXaXcXoDBujaIYVcOmsVJNViIVGSxHmQMgyYwDIDMmqZVy
y1miyUAf0Id7d2UEXjmiJyODyuZAHiwrgiAyyvhqMdSbLBfIn1fLKdEIHGB/BY/S
uUSK3V8YQ6boEyj+r6p0bbs1ah+Q412Zg90yZm1vnNnQhcj56aiwKry+sX2XQFJO
cBouFD/TZDdc5HUt5Ndt5dHdVa3sFtHldzg2GDyUwz+k6JX5dwEj9TiwjgNmdX9s
HwBdyCgicevhf6FLjCj1K6AzTTTy5Wwd9LGZfhSpgfndZ9KexnflA2dVo6trOcbx
IjjXCM62msw458bdHN8QZ4Bls6c8cSWXm+4FESpDIkGzPrxN+EBUZe/0kAQwFYKH
evi/2NqDGifzNnPFhGxPMUzzC6BGFStfY1IfgYx1TTctXWSCRQUzvOkSp9ds8q97
W3+ZRbA47PvZXz8uMiVmHqIxj57wWaCYMC63aQgYWusrS4Clg+vNZKFQrQufoVxw
yFCrup2niH5kN8ekkO0pdwiPk1BadvAzxGA6UskQUjpAwFVwfdjgwu3VD5RAe5M5
wzKjggfdAKb83IdYNNg8408bMXR3gdMSp4lZ4h3q4XW6oK6U1Qgk80H3Q0dcTZ5m
8cGsnUE+LWy1y0Oyo3SOcgr9zp+1GpjazyQGTOK9+z7y3DWr+8oEnWA18fziGf1q
o271Lz0oceGfCvPFyFAfWa6/WZry2WLUO8s6m67mAM0nSImBmNH345fJWuzyA73a
ANNF/1XTUJNtm8UzgEbeIw58UMVYQuBY6CGYJUly5v/Uv1MHrh4/mVILgQeto7x/
D4aCiVIPQHiiRC26lrMM4y+gWYJ34pylrIv+TM3w/YOR1WwhWw5DPUKryCx5FnEg
HFCwX1Cft1vP8w8Tr39tXfZYK4+EIJazZY3d5+1xDZCvluW6r55lhc4hLDP6PGY9
+eBYXfDGEer04SZMapFSXuNEKWht02VedVh4T9Aat9YRv58u0aurrjDIsM+AAn8q
bDpHWwg/4BIFpiDJPD5uxQQ8CiqUlMJL/IhBazm6XHGQQMZFhx/cMT+bVqOQvpQ9
vuWsv6KEwB6ExeZb0xkTqW2ECJWGtBeB9VSl9p9TlCv2ZHk5porAuje23UimmQbx
pEQqU519zv30leNH3iDXoEhkRMg9DiPc4XYzAOvc0A9o8eXJ5+id3mMc32d/rTah
wCbSKMK1BvzXRdxsevTcB2dS3SYWxWLzWB58XMAd3uD5E3SJnqkVn3pZNN4XkXTF
H+pr9WUzt4rUkT1DV/GUC3INsr4a3G8x2wLbs4yKia6v50LDJxgkbg8/lSJ/eLfM
rJPdhwP5OOWnV2S0YXfeWs8ndp47JwRKtq+uWyE92Da6lmTRLVom1FN0lILRFAOC
rHAOjnQA8fxwXFMRsNe8pQ2XUsL/uNRTD3eyqGw1wFoynHdYbhJ98zeJos/SE3ak
udeWhoc27v7M2HY1INHScEl4+ZGPDyjcvIigt+wctHO1iSTENU2Rn6vgf6tT66lY
et0ILEGPezS84bSSYitMZkOAdZXUC/FlijJT+ErBPbxa2wBGYMGG4h4zKMqtVubl
/DSSyA8hH8osokuG4T1Qy6PRn5FDbwKA4b6wGMyx8NePTnysTpnkLRsIaY65X1lg
7csjXJ0Zrs4N206E1jP1lmN3XPOynMNoJrSerCk2RCjxjKhW1nYkoMOMR/xlT0wo
K66db+NBlm4tUYaxNJjPYGUbPINn3S6Hri6KDQDDAgQ1lA0f2foPyc7YAGEshmHY
jpZ70K0s8SHUIPw+TO/VibWeyNtjYaZrVj2ErF15k9Cy5hD3qNGaxW6VDfpKpLKo
jFiB4CDmA9aqq4sbHGqJFrrsU7zCc+E0PDxv9ANnBEpNR3FnE020bOrVgeMvdDDj
k3s+RtAWgAdglZTwhybu9BZkdK4xEfwIM5Z34nD4utJL705UopbuKb2cocYwdTrh
zyPS94bgyMtHxM+yHn78HuaUkzMG1dCt3H64dQlEdW9ZiU31JoL2cwaENxf4GRXr
Qe+IO7VTx6qgQrRGeuKNUOzeKdbS5Di2WWzImpEyQvtMbNDRtd9dSo2lcRFImqxC
q8J39shuCMZFTACId9kHVcp8LhJN6HbT9y9FDjv1pUtDFUYb6/5LBW5d8xzFpqmp
E/y53AEa0Vfxp1+6AP/MHavcWyGrl5fuPFPmuJXoDJSHNGOGWcBoHkQWEF460yeG
gmuHZo7mi3l1rJf3RwQ90gcJcay65k3xd7lkphpDnZ6qsmN8+zVEMwI5nfCrk/t0
7y7Jq31ZdFFg5Qz+QktRMQGLWRm3pis6piLvkLktM5LstIt6xgFO3pkpaqDrQlRW
RO+zkRt5J8ZEg35eRstDmdMZAUK2iEobhEYShIIQxDPXZjnY6lEV7/xxALCkcZvG
rThsokTmopr5SfPbXPFasoGpVcWNaJ34DpEwXowxe724ckNKSISGMoXCUqw2Aku4
lmoYjhQEkBmSzOOuaTa5KRFbai9yrl9xlI6c1caCZ/hA5YYyRyu8wtYovR8oZJf8
4ndg4lf0m78GwjSW2q0mkNfXlA8c1olqJbJp5TQT3rpTL9ih3upI9HFRKoNwijjg
x3heOPnRww6fbpAw6XiyFvAoVftEkckddXw75Thig7jI/4BJd7FYtFcww/rihT8z
3FBq3SJwQS7a4DDYCzynRtGANOcL6dOVEucg2HZhwp5wXx9qM1ZWLekKv8g8z+oT
Mt6GHMjjN1N4v92MkBsWp1l/plcxxn5IyupvP0cAXxzZAY1HvzJvBBqrwSrkdaBX
v2mq0Z351E8/5e7XJp/BuafMp5GBri9teDesZBngElVjgUWq05qTmN2HIMXPxf0H
BM+WZGzwIUrM77hHN30GfOr2S3kVMN+Nwz6XO6MoC6BJCtZSJgRDfsW3TWpAOqTQ
E7Wv+8qk3kp+RLDJIqwkgpjHoGJTeST9kUebAiKIQKJ/7ZVQ6oEqSM29Q6SzJ0Fr
tnytIE/5HcDeNNOQE/mV67UU9AcgCQTpWI0d1G1AJXHVz3Wn+pGeX56WgGB7JIQt
3bjcG36zAnnenl+3AZ+BzzNiqjmaG4BsXSPoTebMsb5BJPZUuOajCmdXo0BOKmcN
GuWy9dsEdccscM0Y6nV7i0Bl0uI+yDCOcfHDWZeMHAttW4rtMdHCHRGchPWv146I
oYDmWukiTt+tTxYWZkhsIMR5+rN4Wh2Cl9DmLcsv21K1G6ZIf1WLHGzTs50U2mMg
C/Fs2OzuM10uPPJ3+W6ZPgKOVLNgmsDX0e5a5/Cia1ilpFgMLiPPE0Ep8IAVmf60
vIyIgKG8j0hR8CuIciHdtlZ+XZqDG//M4R6zCiz2cF1S7s/V4pXNWKL2SsK2iWDH
cvqBjRLbKdObGt1/mg7nlwccQopr5/XQPOzGN4MEukZIoT+0u94GthdUoHxGiHSB
CtVFDMFc3w5dVRiknzKEZGNORH3gjPStog+0DYcgpn08veC7mhsWOeJrjjn4LOoT
IL6hQYIg7JuU6gslSgMb4Y37XbDZ7sGdz+CdsN8GyDGZukGt3ZREbh7ixF4sVCXX
3jDBb15NUzYacJ9EDLzZIn3V904bBaRmaC8h4XNxJvu6xEp6cHCToCl5gNW4zMFm
EW3NB86R6j9/YnfNo3pxiiJ+h0zmMe7GHnxdpygL99S9bYJFBmbct5qiAtpRPlE/
pmxavyx5QJNsbYKy4JpOYTgXRQWIn2L1cyuIuNk0CFNU6t79TNsm7YijTsyipG6G
9okpda1bHdYtOBYgYJ60mb42plIAFvZ/H8ZNLkjLwrD8ezaSitnJEByzCpLlhGLR
xn3IX7BCAGOoawaqlolWQf521qK4MyS8wvqk5I9cewR4m4HLJoJAuogJunsG0OdV
RQJLAWAbGFQ/UpQlH2cyZkg1ji/fnGAimHgn3rJIq47LiURtVlv2ZBPeL04XNtIV
hqtMqBvoyYTuL7598ZJJhONRs+S9Rw/WHaf9171Gzfk12quJv/epKbJcujLmf81e
kZGi4sN3vVVBvsf1fwZ5zS/V8IMg+UGuUCmtdU8+izhR9/81FTvKrRV3WUel3qBT
+P1+r1mb05ioigI5QYuLpNBhx1Stzmx1czH/JF5Vlqsh0A6xMGnjWkWjDQcmGeD6
pOn1bZd3g8gdG9OynWUDQvyS2DHjukg/7stddpGIaKCvc4BiQE3kTvuNIGd9gQg+
6jWgCN7GQ/6HEewjpzvkXodzlM9+mIEdD8VRztjDNqhZKIDSSZxP3RGpFjoKcmUV
QUrd/ggF76x6wB9GNvoTceNSWb0x9NF7hA0B/pb+4ozByGPq9n5YVSXBy8YIXUM5
wpoA4KE5VWvt5H5d1Oqcr/cMgwUz2OrYwVAoWY6QqR5mFz/KzV1aV62YPWYJVMte
cNew/xUrNnexFZaqLfLfsYQAG2bsNSOWQhNRkfUhAzoDny2Pu8uHK+uPeDmbHy3B
jsgH6wGzcwtiSlKIwDfeIncGN+A21zsk9HgXD7iRLsIE3WBh0PWq9SAEw4TSBQql
ylqal7hwZJaLAwOg+AZ6L5uQEjIqxsDD2SvI7n85oZQQ0ntbhaTdR4bUIVuwlRoS
svsEidfXN20IhZgaGSaHKA+GUC3q6jDLL9ToA7d4ysKHtfqLaUvr46Ygs9bBGH2S
tI0+MaJwa/SRMETP5jYMioJwIhfq6liN1uR0dxcmFzh9fpjReK9praKay4Nrg2eB
4bEBhhA9P8kW4DxDt84qRIC9WS2e+qn1OPkEN8UuwBodrmUyyaFelp5YPKCJgwfN
LNtR+NL4oTx08nrrO5/v8dkDELVP7u40Ai87KMgwgsk6qdts+SafWjtCiFL56Ebh
bbElsDInQ3g/WyDjcVxX4cE4MbfTg40OoZiXIWwnXBublO2UDPs2nMUThH+MbT06
ZOLEF9+001Nmw/JlSsM3mVyVXsLYlhmhFC9KJSazK/pBwGVz65SmAoJtDDm4hCZN
e9YwzVKBLStyF+xIiZOG1mIiI/Q1r2fK0sESBnfmWoZE7CxDszBpxo3wSaqyeuBa
e7LuqtA37zbO+PrpjbA6IaOrw2mttg/BsKeNVDLtte6n+iNJk16k+xeU/jQvbz/q
yFsZ/7k1m0gK4wXp0dKf+cyUEolPzNQsujhyTF/m6vHYPG5TGguRIjoGlkiXtNrX
UJD75xmV/qu5NvMdWD+qZdc+fT4u10/hpepCIZc5Ui69FzAr8bj2gIQWHRU6Orzh
Wddmgd2ix+Xt5YtzMDwNoUo1Iz2bU7itnF1gByehjjGnXBGqBzrbaBdkOdkIiOUY
GxrxKLOM3hi9Zv+eQQAURSm6JGLx/WpI9XmK1Ub+fn33uuL4hcXN+e9j1rO7ZGoc
4PrmfVpS4FI3zV2yDbtIfjPG3NsgkdVOD3onzY8TPGooiVy2MeNWaAAI2m8HOI6b
Vy90GJ4Tf1NRQwBOQ8vvfabRuR2Hqn52VsWoSsXMHO1I6dHvA6j11UVsA/xkazeL
LbR5+fIFf6uZvGKZpWN2CVAQ/fYTJ6ckluupD2NLVGFOJhi42q9fHMvujkhPdt+E
SKt8D/5EZ1kxm6jZ+24/2jI1mo5qpbXwc0IICXXa99rX8cgdu5f0i0qT74yL6rj6
GO61H1oaKMxr/OJdCbwOPf7KxHsZD6pm6b7fq6XaQ66kYfdafGIEGsW//3MhAiqN
f/PGTYp9Ijkdy5XkkwoFjN6k94FdGNhojHisu7a8x4IxrMo1gNwkyQba7AgWP9w0
adu7bcqJkp14CeKxgDHOBpKFE3kbcrL6OW4WlE0a2O+iNmj7lNESmXZzLTVB87Gb
8uXUb1N5EpEE2Gm/cQBwWFdgXGeOpl67kdGkSIuZFFUW86SUIKi5VnQ+/lbdRd2g
/n7za4nW7baz5zr2bQrJ+4tY/5nBn7Z0VKTE0S6FeoiOXJHecXnu5Z5v8GUcXRQZ
g2Yj9+cQxN4ztjA5K8frlE/8HY+5t4TQwKjkpAWQkLZHoDNlo/Pxeqt5NLsTpIBv
nOpJFUE/jHaUXKd7SKgkLclTNEzdDZEVT7QS1WB/MhJVKj+tRs8mAlL5lf8TcWIt
b81288bHORrJBE4VmeS1Nf+EZ3ytl52ea+fOllsAWCwqh7rmHPGgEZ3FfZD7fP20
deLbfIjHXZETDkU1KKACzUtKReIGRBUeh58zKH8qgrQOFQSJPOBqzdCJTQi3Wj57
gH/Zc6mcX4UXeI9k62tFtiWGUMenNaVc7t9ECg4owJLQeaL8vcA4cBbDwlrrKHie
HrbMtljdwW5DbDyxzipAVw3BKjCIee2BTgyt6zbO1yR8dY3WeWyG2KHasAFfZsNb
IlrYtdAMAtoRZwEB/INjrJhR195F7gMJXmrVKb7CvoOpqtTUtLpAq068xvvEd6Xy
4J7DdWKHPI9JUZ8L5xqdtLrVPWa5bUl6EJr4jwbUvMd+qew1c3aydNfa316yNhAB
oal0dLXY77Q48lRJ6dDuacMR7t2YP0c4ad34zlRuT54V5oOWPP+g0qkQBmJF/MIp
jHj2aLmt+m+m3ZzevgxKF2ZdPqy2QPpfIG3MEhFuR18ZkDaqzaIl8pVG7HbRDZBE
qrfAocyJ8M4TQZAD8ssOMclXwUedgUGTU+qowB4Y2nI2PRcdlfcid7TTOxL7H6a3
GZibQCm7GWDqzCl6ficE6UKtTesLFZIomIZYjL6Ets8hcAmMnt5vL+UuZ6qp8El0
NiL5C0UtRieZJVXEf77csegLi11rqdOW9aXz3x7m4hZW0afsLeTMxi367raS9/Ii
Z4XkWkaCuN3wRHPvGNxaCSAvqF97z2lm4YaMUU9wOtpNyhW8e3GfsCPxI5hvTbfb
5yiRH53KnlArXN9pI9lc17mkMjWouHPA1moW2MI481UvFZ/xG4UUpUGykQuKKQQ1
cVrC4Vm0jtN/gmVWy3qsSYiMH8VTVggT8ogU8JwL8oIWN80HJ8M5UpcVzYpI0m2B
EI7sbsGUzujvSbvPbK+80NRrKSPgFu4wbpJ0v50WSrq6USfdthx7S9JziIexyb5u
LudH3FR62enxb/mehgoZRF5BBS2c/1oIdi963yaWItMci4Zto4qV5P4yh7k0Hoki
3lad+rWbltUqald4AncTUToYnM27UliciQIAP6lrY9gzQgCUYlj3stg+vxM+wsK2
qH99ljgSzScpl1IB8/OmWw3RuHtA6yD9D56KLZ7bCm3h5zeSokQw82M+kmWX0tCL
+fkPxjXUsmLBPgwvXN/7Ylba75oHK/rzUGFymDtYvviZBCMK+zC8YTKh1OwIq28c
0442nL+SqtE83uxplvxiCmnwWDLhNbbbfUZ23/aee2wzfdt+grlRaNvcbED9aY4b
PSle+0CZGGBuKrYSB3RQhZxeKAWrRao91LrKjU65HKakOom80DZqqkhlDnvECfTu
sZLbZI3PHM2UrOGu4tc8CgyhTsULtrdRFSdQEuman5CqUp4/7QqL7rasKdrjl/Ld
Uo385sbQontMCHKH/AIsK3dso7BPv+ptQJL0fM3rPdhAggxYvo8ll5zDk+BxzkAb
PLP/hyTieieYqs8EU5JgvjSHF0m88PalTvH+I5j2mJ2I5k6DtcTJr/QJ92ZPcfNw
Il1jWg2CVgpzRvJfYz7cGoruCpUKvs9EKbRUqd70VmUMMqt4j0y9oxf+fW2QOBWw
YLZ1nEDS6zN/JsIMM5a+tGiWFjuFb7zrRvqmO2t0wLhAnDKBdXxsPzO/AtfutyzN
qtpA5BJIJRnAcB9bPawUyi7wAKciB4ABXphaQp/+4iovgFYwZTVZ2Vk40evRxRHM
KRYdMSxt9hTfBFGz6el2VQCfKgxMsa+dl2RIBudNTFfz6eevFismbTJtkxUBSd3A
61lxTRkhMlSCaZACmMSksXozb9Ae3pIZZran7e234j3Jz9CiWNg9ZHWOr3CUU+0m
/PpibPDdEu9dZbOz1MmgepK4ZSKaCT3i7He8Vw2VxJ/8joFxdqmsDX+n5Nag+p9u
QOQHME1oojbWvGDnUux1bXeRKUMdcniOt+TPk1tvmSpt5V2GYfN9ZgBVUCmiJWpY
elwCVZCS4BJ8h0VN+VrnwASywBSGyiW+uPc6BTBwaXra3wU+kwP3/sNOeCKvQp3h
7DAqRvgBzCa7EQ85MeBRO3XQFD7oXZyUhIqq3HgRJICil6hZ8RYhi6iXcvg+d1LW
GcyAqWk6p4D4oJaKDQUifl2KcHApvNKnP739zVLoIDgsBLcVk9sotP/FtQcdmkxL
SUekoS+WTn9I5dz+6xPcq2yVmje1hwZVewtE0eT5qWPX4HHIK5SdRgksCgYnWBNq
tNtRxp2K6r3s4mw/nq5iu2bR1qldPlZJ9d3vQnb6IK57wpccX2CMR+yqMBOq7OPo
f+RMeT2IJ3InmRUv6CgFVn/1yS0uT0bWMZaSyasitvpOVoMhnyoiXZAHLQnhIONX
22gIYO3NCi9izMNX2MloCHCJW9jWIxh+eAj6h9G7P1VQFA3xR2Vmz+coKk1XKk6L
VJ/HlUCCgZ7NIaHapLyP2nQPc2MEhTtscGLMQEJNC6i0TuKU+lj5VnsL4wa5bwWB
cEDvzzVW6LLibwH8PXnLV5rWRy4TgAtEK8y3cK4vGMy1GdunNbmLFOC/y2zYAoIB
imF58Jv9boSbUa1XxZgREGTOZe2HWWwH05pyQiWl+ttNTcH69fm3tZ175l/+Vv/z
m7BCP1ZcBW5BKAuVzehTv795VcblBYExxxiFhrJGu0RIlZZOuG2rEGuuHveNjkso
yjjPriaQHD9gh6ivWBNDuuudytqtxF6tgafrCk8leKgZEBwpMVQ0gPNkT2ctNH6G
+4Ry1VxAWnHs9h1vgY4QkX/S4bwbPWCmvg6iHgmQrSYqiN9w9doiXloQP4cCmCHH
fhzSADCHkYmbedZsQRVDT7FlrZox95rrdgKjCQVZtqO7qjhA+TPOrjqCP09FmeWq
r7YLt5XY169sYzYf7vyNb+7ZQQxBovdLa2qPpS9RXyes3uvKtYxuKWipMvBKyZ7g
EJG+/X9b5o4gS9q7/XAQZG4AXD5diafGqYU/NKKQpuunB5hjt+jqWI9Y4PuCx/Rm
QDFw+hJ19Ujb+FDsAQgITg2aDHMbi8L0g6qYqoGHM5w/fn7JH/wyVfGPV8cZdDeE
KhtwQRDXd7F/XSXgGWWideLm4lmCMvUV8S/US3dkOJhuJTwWulGxilHdcHp4vA46
NnoKkMfMkRIT3JFPOpOdGlnVWLfQMg9UnDgWk349QYHuxBy6s3kAnAHUF3qG7Q2S
bbDAihI82i2vsSsU/2M1VKgVJR5fQyNuuZ3Kj6VCIfC+W5lJo2pTic1P3Hmd7hKW
+W4e4MJxV5EkR6ymJADa/SiANvGXUdkYd6atLwU24hSE2zRPCUzebW9LECABEz8n
XpCQ1PqRnJcVZU7k0pTMq4eUqvk93F2gr7dMv6CHZJs7AmHbQfcGwsF94GqujBfh
Iw0pSZkzEAubDIgLjBzjoGaHImiVf95aEt6jgGPoEEpPZW2T25ZEm2er+YIPo3fs
s2y9DBl5aH4XXtBDL6yXDa88EF+0QifKiIhJlx+mlrCa5ZsTg9iF9hkMonyhudyo
F0YpWN/wr8B8BUFx4D6/0MIQ/AqA7OJ6vdV9hQcUATCrymm6Yr7Cy+hYcbX5252n
U/Ir83NV3NQrSQb+52VgVtNFYmzdIFOPDfxTiXlVLGc3cQEV6l1NBtQs53eWFhBP
mcEItyD8a2m+q3pk3L2sK9Xfb1a3D0ZKW0MSnrNWOUYCktjGFjcaYzG6hzmIIyuw
IqOijOQjSldxuAPLidldBvrmMmm+FYjk7p8W2PvJl15tfV/gsQsmmzPtQmqX9DSa
quO2t7afRYe3mkFoe9c6Rlg87Ntl9L89NuN+jmbC/czXWbV1mDrS8erdIDkBG/RM
pHvmJ2mTMFsQKmO+MeVU5fqN6G6F3fY/24bXlz/ckAUpfEGnS2LX6iBFhtgzydrT
xX5CO82rFX1HERw37NN2Tqa9nypsWWzNR0fI+Ra1PDlTSWDtl4PvBDz1kOCfigwL
Wu9ihFVSy/DKFAeyTX4p35nLE9B4nH0MpV+6UtFY/udo+AZV0asjhD7YP+COVWb9
qI1bOaF8OeTQ5ylAEt9eNKTi3himedmtcnbXNgBp7njMAwFQeqM3jfwDp86KJAvV
SgTwVNtNpbNBdN1J4F1KcfzZF3nRIkNNgudaPR+yw14EVS5zrcJ7JO1uObMP9Jo9
5ZfnbINvEToTZjMtPftTOh0pge60/i1Ts3udiU9GJssBovfNwlWAq4OlfTOLBItL
I1KEQgYMSy8/X8fJhfyvqZjML4Ac9XhZkBlQ3kICmMyL+LSTIbV7NR39Z474elEC
KUQG2hyg/JAj6uB2fJ4GWeaJgRMDrqsi/neYHJWCynn9DmqnJNzwEkn37nm+Zt4g
h8hM1ITXzzL50tPk0tXDi4LL3+6bjbbpo3s9BZ3543NXK++D9tH1kP5zrAeusd2c
qY7QDhkQgTn0+pc/GoHhz9Ev/zTipt7GjTGJT6tpvGYBVeebEpACKu4paP/sCVS5
7uaecMvREyyDKwLgd4XGvO7ijOJe6/swLtyd8fB3df7JAW2n/CJ4yaGFX/Vysc8/
XqJDV+PdiBGlOAdxNLygjLP1QL0sks79K8M6q1736560sNVqyDjxIcnhjTkshiiE
V9C/2TLPoH+gb05KzhAjlWVF+EOGknvVRn6ZmEVO+vVYJ4zhbPU59FCZeCvjUWIe
52Hvj/vRp7YuVhe3AuyTi9LM7n//gErJHOO/6jG5M1KyYWTZwCBLfbWAp/9WQtuO
+f05U9ECMNauY/xno+6LJZbcZ1i/Qw/ZYEVrscCcDClUrSAM/jS3z+IJ+SrIZl+B
O4pGTyNbZ4DVaVXC24jDIIukT7d+5QbY6j51NtfVeT/pJWbfbtIQYvw/Yo2pft8s
s0dQ2Sy0fjmyZnPG8hZydmdAJi4oi2U1rduPSVJcr/6t1VAXMwVXopKTSoe8GRlM
d/ltO1wDMc3ZWNLbQ4C0yZX4zVg6Zmhr8T8ZlLLzHWu1Ub+CydOx3+AFEoYHt4CS
AMctEj7qBofxGIwmk/L4orldSgvdzdvX6lFd+H1E1siTZwuw4JJXa5VzSt+2WU94
T622aZ0YGyzEBETEq5vomtJdBj1McgF42N7R6Xkt428x9V89YaSArN7C1MZqGX44
p6r6ZlBW+jZ/WxLTaEPsS2eozLqEcrMh23B6YTjZtIypsUhxu/bKGKxZutCpKpow
y830WMJDIkZJTMJktVxuqZ0Jl/GWYKROlFe+OYcIKGTe3V89RobbypRWLC73OXcu
fVpx13mB5UBdVeB1EMJyMVvTG8q1+YfWcMtv4HgKUP5pQKB0yqVC0mmCb7KTdWme
U0KYWwN20oitVU/jcc1SSj9Mf7ajDb2Bu8eTiuOIK5ROj58sHqavRU/WXyfbzGBy
JjCKaFwu42Z2s+jBZOWvSLXqdL8ohW4Pb4Ox8oaIpseBp44WEw+KoBG6REPpPSM3
zE9SWRXPEghsWcrEtWqizIYk4k7y8KqC7hww0xsEPVDB6i68Vz+mS2tl3w2aZvX+
VVPQlXdcbNric+VKi/Fwk4S11oyZ8JCTKvdkJ5OJR729jf6b7td2wcTgGTzSs10w
e5lAePXxEpmdoFZcVZ7ldYbVLYGKMGTZ+T1SzU1x8kvNr9ZGPq5OZ6JXYWHqmwTq
YNbIu+JP9E9uhe+RMah/SxmsqtkyifSi6q3MKuNv0TudSbw0DqYsBDsAX5w4EsB6
yFiaJyhX1D89+df+XzGTUHtL06sRcAuwRA9Bdfr7/UJ7UZWqnTzxOQqI2249mU90
gcSLJqW1PyQBGY7XCUJsFxQiJ7C/4Ei7rpqk1OiK9nghD2QxawpqKX4JMX3ecLx0
hdz4hOcm4Kodo3LZJrKVI0GO+ch+QXz34iYCF0QjTw7yOTgNavvG9hcKy6xwyGGw
UDwhJApcKh2cTaBUX73bMa0fhHk2fdTCaMUEe7qk61/hwGSVe3tTmrPq4L7kA0AQ
6gQSrw/lFclMI7/mOetJGFukt6Qk8ApvZtCx75uszYmeFiHhYmYhSv3XZZ7MOzRw
9rZPTE7spD8GTJrGOp6W948tDFU0Zx6dDY3kFrVd2oXIPQZzmGSECW7MmyIUmJLN
XLyxUXHIMSJG/KQHls9TTfVye2voLbgdKhfcnP2qImhd+9/KK4e6W6R+fa48JHDX
eZCsjTtIbVuZA2OzS3KpqGoXupZ+4kULJG+jnPlsTTbNgwh1ivOW1knlqOW/XLPa
79qJc2Jq6ZOw0Ex/qdq1sx+4bseFfJV5Abk1wMZctnIdn5Bp9U0PPTHPdmrdJjl1
OYNtH0ka3XX/HI4rdWyoVnDi4qcyeejF6ydO6OQxZn6pgvSrKzCfRU29XepC8d9L
D95Y4WXC/LZKPeoaD+Vi1jCzeeeMSHWvgx36rYcKo/1umKh59U92xCILxv57FAXt
SLEd7uqYLKmUx6xPoFhvMBLzAkNu+38uNTxyPY0u+PXfdSdTvC9RChbdvezVhO4V
RJTGZa0Ti73nPiXrCf9YOspPNZF2e1Yl27N4x6fOHoShW5uHt2SVFM/GVl4gL+ZR
mAcn3O8dWV/azdATskfEYFN35XoAePvwmz4BGgTBNgMhukr8j+cm/jlcm82zgp0e
ZlwlK0kW3s+qVLL3tuCg8o5AhgQxyl1s4TEucLtAo0UXzP5CTqTQGeE5ngDaCGe/
/qfbhAIbnSSnhvOIDV+wq/5RYagSado49tm9gxH+HE6Awo1rSrHBcUM9AeNiZQcj
J2mQ25eqPedKtE6P8PFEIDMITsf5DKA2XNmQvl89Ky1hGxJ3+JozmiSgAt+TLTX4
7HnnGi81dLR69qqHjgfZC1QUO/YlPxipL53oWXPbe1yDA+SUKWdXaqjgaaJbc04K
ySW0HBEZ6BGG8ZhrNE7d0v/mo0ie5+DU09JGbQ9jyYj3L+PDkRuPjLirW8B9AZKe
9WJl/rvaFlmq2jNj6/EzKwzcrU9KW6Awa5jNn/ohi/hbMWrcZCMm3Z3it38hF2ME
1PRjMY9QdYkxjNXJLQ/vBWAdSCdph8X56YMZS556rjBonExy08rvNnwPQPJzFFIJ
H58I/ZI/lmVAC3LTCm+sQRTcIfMlhEnu53u+137Q09dhvZ45Rjvw8wR+3JkWF+Sd
SoNrdvY4zs8ip95nhnPeEc5MMbYGyreFWl0Go+8QA2ferB8ouuYkECL0gCTNKNrM
OFgJKWwzAeIKqAkND2fOoD3A9ZMMhdKzFpRogxK4Bb/FKB+xnGgCAwPODjDZ6YgC
OJdMSF8duJG743lgs2RQ7u5wKK9m3APFQfn986/VHbeuCCmGzTruWmvs32iSR3dF
PcJ4UdyGe9rYjUAD8CRYvKHoFZRn1IzmoaMPrfzDHXAQbFnVOGN6wsD87uw5rVIf
DOZsx43ztK1xmgMuE5TZAOg6BpEYTJPSf+ZxJn+vu2XlorV0VHzYe2N/mX7m2tJs
UlgO+ZJVKlvdPtKIHklV37XBU71CDD4lBKCv/drn/GJCxrNDKSrdT0gXKeeP+qTF
O+DRfN88vdrbOQIdwHVZc0Kbi5T98+arjKjLr+pQ0xY9FTPjeRH8rngkfo/y0oBE
J6hBjI5LxHOLjjqUMd4fCy04Omin/k2KchM9WKFr1+VmpTmP8fdxHBA0fK/QJyTb
2nO4ioC3FqHVfRrf+rZHcqHN1O8fU37vdEDXyRYdWxPqGMXc++P+jp/1GHgvxya5
mHbOQRU6aoyzteRvGbVaEIf05vtomK97/EKK+U5eSRYerBaDU6LRIi9az3WPuigy
B8+VbeyW3Y5b84i0cbmBe8d/o40HkYVhdkK20PKToCIsWFq/ygPv2TBCp8m8FhfI
GDLUspLRVJCYeSfzULEww5b/sGR0/oCkf2E2pL3dIdXIP+MlaxFT9wV7a55Mkk9r
sdh9NrYJ3i0mNavMHKQLEIuaxUgQQLhlGuvA/eELDPOiEzfN+v8Mb6XIC9mL3iBX
7wQX5rXqa7UVOpbVTpqe/Z8vqJE76Tvg1xmFVrj4uqKKmz0OVKPQKSr6Q63X9wjg
h76Sm0etsVqT0gjRcComMImR39QVuNix0S1Zl0B3W4xk61vpBaw4eRh8P25oEy79
ZehtTU9peroWLzGkTyUgIFJTcDRBdUSSg9j/j3rS36Vsy07fm8L+aajFaZyioXpS
UMmAhklaMSRRrrw/7kX0CfPb5S9LIltEQWjM+AatnEZsOvVy4eB3GvRIbIdwK5MC
96/FSkwTm2sWDACffP9Rb5BSvPiBVhDEIJI89hLsmYBEwHq8ZF7W317THVll+USC
4D2Nh5BbhdgBLZ4nTxju7UFDJPf7z0VgkfA+Ljqkmc/Q9Y5Gf1OR1E2Dqpj/5n/m
ufWQFrBwdxWtZpJfK+y0GWh5bfiiyGzC09SOFDW7vJX3g+BGRs4TIkmOESf75f89
GaXo1Yqo0H4lbGj/VfkKIfHK2XJ3Em6ja9r5dSM3hY2AnSuOXmSaoQh/cwQnaqkI
ruQlUIdg0NOKhWtdg/QOEbA3V3iP9cBt1ORK/GHFMYvHfQC/VBFqFHDMZLaIUw4i
t4I5THfpHPimGuTgnCt7VIRh1lYd8uwyiZdn4RlbxpHopRDfnVc7mfqt2quCPfkN
rAx3vZ+J4p0VV5oDUeg2jr9HHUDlFdHy+J6vnHD2KDlWir48I4ukG0dw33ueq3E1
Qp1Cd7LIF9VBAjqbb5Mf1jiUEdg3YxRBIVW9L+/8Pg1yL8ZzVFfEXbGeaw4MlUQn
gZdYErNi5Dk5BNgQoSXsVuxrCWI25koFJfT+pVXX1EAlCYog4fXLm/8h/Mpu6GLM
mABRzWHz5CBpWdu2NyVcz+CKSN6Tba6yCLucuvJpUZvGSkMcSpVXyXPbfJSlSkWb
+thx/wq0x0YB9Cm8jcZcVpA/RrrAngIwkmH6j86NKF/YMk18PylUadppoN+IpmI3
XiUfoFx4rRJLUeZ+ZqTHD7coaNCBC3DMryZfKKI16E2qoTChH9JiWWHE/Prgfqm3
XopMibVFQnCtA8ElwA/xqyAOcLaq81fmfrVCLvbBkEsf/F2/m/KI5JHuYeo27jsh
iFOcSr2G6QYRXBeh9Jt9ihuPMThQlhYb7x2RME6sCI1Meyw0n5/7uYwvY/SPkrjX
kyvU4PHfLqUanQUmX2Twv1+sfEOH1G8yZN1s05FygORrZxrJwAv+spYXI//8007N
YYpPKzthjCc74xHChEfSfes1Q3zY0Ell2K+hXLRE0ZQhzLUmPms7g/tOKgrvzqiA
pu7BhJPY3ubUA4IesjzZzzmZ9tvQiSCzJLv7DSck732+NBLMzxC7+iohiltBNlKe
d1ilxtE61dpFEaQlzHX6HKzoqq0iT5FiBf09dt2HnmcfvqfcVHbFH1tqqheS26G0
JJgzjf8c3FNPYNP4+dTy78eeiDlkZpppOCToiEdPI+8HvQNjNfj29adsoR7g/boC
Np2UvlkdCgsVEGg7teXdjD7FW5QQaF8VOUaKLD8OtPzjlkbsPKNH3Fsl/5eT0SWO
cmRqKe8v5UYEgopijO0zNSObuG9VKiAbyvrTR/UCFxuSbQ3CUw95K0DDjTDtPvlQ
j99koBp+fL7HZc1rBQ2G2r9hXsYXTJtyBPfX+E/t0PMIIVzSJJrJZwP9UQwk2AHF
FaCBEkORe6qmG4Jfj6/FeIffX5IAcsOkK9fOqgFGIP9hBLcJMYlQcC4w8rPWYw1b
m0iy+qK/ePJZqxHE7RmsrvQ97UlXcvwigRYim+oif3H/kfJxZjIyjuOOPQACCAus
1fbtUR9qjwF/I6b+UQYqRBZx9FAIAKyI7i7TbgzApBvJqtmki3SL4/+IMB127zDY
N5PMbxBwU828DjndUUIv147DhQ+00A0ESYuez5vQK1tuRM8f0lOWHIj5AUlcF4jy
Jm/SQTu3QmuYdzMVQDGrOJsieeX5WKDwu6NhH2dIyBokNkzUmr0Ohy0CMkvypfST
KMmOCPHXQpm+sF9mivuKAzdPQEKJBZW0B3P13SuKP+cRoAaJVCny5s+mSWsalwVD
/iniKV/sC75aQf5QHKdSZ4Xkg/ioaKivC9mu/pIWYrPizW1+tX35TfYPj9fxxZCH
umSrQItm+J6/SFicWjIzkL6Oao0Dd5zqIoN+vi76uuhpbr9jg412lZ+UDy6Ob61H
0QNSP5iWe9kiUEou3XZg4XKSqcCb/tvt6X+bkZfqq9HZIXLzBfQbmC4eOm67XoUU
ErfoHgdMLP246qr6H9z8x6AHOlSM4xgITGiCc/60YolRfKIXu4nYFjWacSb6ynx7
Db0XTidC89kU0xh+y1JKhtXjbKXio6VNQnhzFBChddsD5iTH1d++VS8uvbjD72MO
Lnt5t/pcmoPpWz5htUhsR78avPbw/JQZTUJ9wJzvFIPml2tjr1jO/MOq6hF22n+G
QKEsrNRas5oZCEPE/UF0H/+i9Ra9mLAlg2heZPjIePgfXCrIaxnGDaxH+dJNTi2W
nJ1uuIYTclTFt4vhO1XLmcMpyUkhTIrtgNJoN8bGGaSJc/xFmvOMhYXVgXoRIuZx
j6Y7PIKkeMmofbyw03P1FL9Ciwj5YZhfHJipMsiTccZx84uRVcQH2gjIufrwm7E1
S4qLa178z+++zjYpEz3Dg02yHYwtpXCrOir5cNqvla+OMOUvAXVgBbWlQP5o61Yc
Ta92bVJP5kag7bwnl789PSilYOh8sfOT4w1vbbCg9i6YiCx95GafVwFUw1me/0WL
gq9G0/KB+LT7Ybbp1nJLbiyoYdrLMS+BHEkDucEc4cJvv+oWjFvi57rwowNUf/68
AkmgcGanOePe+Rw+HQP873rCfXyHZCPn432CwSiO3ijZGMNbPiCZcwXKVELcLi8R
yKNT+ncJCNBVEJKs9TLfZYVlEAmbTPG2BZ+TEcZg8cyLAUo4sYTXPoweFKi7zbEx
Qu5yNoMfW3zPyrMaVZ9cYfuvGKUQrl+XX8mX4tIvqBFHyy/aanAjbcwZ2wmTtR46
jOpKOzxxcj8h8uBkH394utSMMUUcp6Xp0Q/XkWxn48Zjf18om3EYPnEDiP3ySMLZ
jjCmb1vNxciwzJuSwBRsZGl8ANDG9BBf9MQUg2WQyR7zRQdyzbp/+WJo2Swzec0r
uljiPGZvvUz8FuHE939sLsPMDem+VJ2q2IkcV8nFEhXy7FybBCDkHmNQv087gDjJ
kvQDmHprs9gXWxHROqXdsyPWqoMLb+ZDJl4Esx3JbbUGRb5UK8hIGyQizpePk8DN
yTetv5iMutsciGngeZVYtZq70GOBucU8OqqGfKmiX4MUEA9o2FcYXldZZSnqwXrD
6KU15JxFOtlTjR/fr+BgE9H7D81A8TSMk0OstIMKyvrvO/Zk4hhTvFx1sB7smo2h
ndQQj7MarFJ2mBWdK+A80J/4qgPifavkoDC8HuWIXy6Y0ENP6wtpJn0Mmi1bP9FK
KZ2zlt/QOU0fznEAzZEONsTT9Kzq3MJ5j9+1jhGw/5DFeT30HMwv8JFwyGVV7JLQ
nfz0PCef4DD2+1ETKj9/fJfUIX8EIWYSmrnb28p9oygrKoCnpNzXVK8/k2IyLAT8
kDVEHiJ1iYR7oilRDyn3e24nwb7qp1S6Em3I5cKyHoQfi9MdYh+UMc6lneKnGFak
sdBVCqn9NZni6llC1D9nk6jfCUJDve/I+em+CSvFkfHEmOoh7sygUq2kVIVmwTUu
tfr7dPHyHwruq9U7oazNKInNvLLFuvPjm1Gf3lDFddDw+cn/2+4mKOfQIf+SedZH
LhyiBnJkYGCX8RCf9XcD4dukaAggR0T1/eFq2DcQfC9KhzwOss21/i0kRAO2wvww
w9urFUuD0wTIRvwP67sc9WQWzNODFnHh6noHYrRIlK49F2cxlganlWi/FghbVUpv
kZWWh4TZGSnYQNnaGjCbqTQnt3j/qusfWhbnxpcbMc2kNSUOD16r3FYQHq/2XUsk
mY/x6zQRwTVozbpYs0iofTX/e2AKvMQWVMIRJEleivXKNrIfPAqhAs3Fh9hIjlnq
4A9LhHM2hrXRR+aAqir+Vi+Nf/tjtYJ8tLFSRWlCqCJFRCoRAU01u1Ug8VLGrZBh
+TVsyxcxMXboOtxg4UbCi7PVU3UBc2qOG7H/3vQmxHYppb2t5NGaAVuBl35ISjAN
jigXRBoMz5814bfp/IYv7/7S7da15cwRitoLgPpo4nxzAGO+lSiCuIez+ZWuHvNm
E28IPRuqRoM2UwAXPWUjmEiE9Env1+TywH/10gfcfeToeyI+cj5m6mzY7ykRkuJa
t1h6FPzrLyUxQxb8ME0538XlaFat7VrLr3SQCDrH+7HotHwS0EjlOo6yLLCAyGLJ
EUkllvAnIFaqMH2RHBuH3vObnTM5DSf4cIplN0kQUsp+hdxUu/vijfhbBtU39O+3
7a1JE2CQZ3ALj69yHAhvCLfg2QAb21i6jcDFJPwU10EEjQvB9VvMfaVkyvvAxKyV
JI70p2bCcAOEJQY0F71Ux/0rB0drqTJ/B17RQLQeqSu0i0Ks8PFvebzmOzKWtAkw
SQrtmCOdtCwwGZlXiFAI/uqHMfyxS57OzthvfDTa0ZIyAYo3Yda9CyDO43GvoUPI
F7SRA2Og7vDbn+adRMiwcI4SQEgcJFPyM2KVeVk9RniHXUhPlYD5sTQg+KwJBdG1
BzTpr6/Xpd83CeOq8kuzQPCb9xU0TRzqtkgd23gzxYTmTbQOe5DvFB6jrmSp9YA0
MbD8vYuIFIEcexTHLjfLOotGewpPr7S9IC8xQyNuFD9XLNhLWwz7CgjB4hTt8T5a
w/x72GdKK4YQ+K2uylaEYx/x2w8AUP0ngL6cDhJvuHvsIYR9HIePvuKTJHLbCQ4o
RkqgVvQpqJs/1eCQs7tikaV4+4nDaU3krtb8QhuTu5UZQbRbtMjbBxlENXbdHBib
7dDw6g/CKyDkNFqDkzZCDVdmhMlLUO8lVXTzuGcYrggLA2fzjkalIqHXmJRPF2rz
DZqtyGQRPWTUukq7uhmaK/xxbyZc3MA//h4+gKstitp5QjkgvpkNnYv8bXdBPKdk
TfOABJQy5aXDsjJm9WuniZwxfM0o7kaZotTXK5wGF54JT4rVnNbyNH3jNv3HVqZp
2FJrwDIP88UnVf21SNzFBPbcwd2nOtbI6JtElH3oDDuu0rnIJ3p8Shmmea+SYUpZ
UAR2rVgVi4R3gZqVvnuBmt+hPkpB+PyQiB0hRQphpqbzBMRkiEO6UKpt/xZ3GIaf
kjwt50lvU2NGVgrA0o9bG8KvZ3/nQhxpTXmHB1uLgZt+aoMcmby8glfjPhwNLNH5
Da7RFxOojoFbtTUaw3t8DJSgjJ5j1O2sJX76ixoejOwH0hVqXg8zWbNUuMZsL/S1
WiigyzqMo99cKoa5MmGYw5duUbddW5ACgTK2OmEc/GrKPE83Ay/Ch4yTPyNi3dRt
TmP9lrvo30IrGbPzJpABQz0kbRkzDV0ymRpcKIGshyWdFfv+VSpRA/yzrZppVIZy
C9VLvFqQdwRQW1IYr9x9dwLRyxqF/nfSYD4kHrUCQc02pWZ4K70rBMxLyDlu9bTx
kXReUgc/UKioB1LAevga//ExQ26wE1TtcuUuB2PZ+/VrRhe7qxSFRMYKSLspgd6z
eXoVCHtMEl8jDDaKgee4vu462YGAn+E1PZWoxo5fzH6NatKoMojzOe4TamPehNeN
WbgUj7Y7q0kByYiFVGwREUdy3z2SnWPnHsccJlhBAx+bjQkGmrF4OJ1hCAYOP2wh
RGFNo24LqAZN0CYYxsNGWWhf1sQgdGhOzpFeVkG0sL/wxKRojTCHn1+XLzVOxDaq
rJ1mLkXzxV9Pbxxq4RaPOkowueghIVlIthLpvm+lGKGsuzg+uwKok3SmuOto1puL
YyXMZGHBQxG9+VajsLCNhHsK87wodAqJ3ab1Tl3GZ0pryq9j8chndv3gEtDwTslE
ODRmU4t6l1CFfIPgsJ6Ift+GNtJMtbeAZ9tI8ej6tur4DI8YYM1WbUUGdAws4lA1
Tz1l8FUwo06hHP74j7GtyqKzsjvqwD+ZW0Oci87BAnlSu09ymGaRvj3t/Sq9ZJCH
ylmWuXoJ0sRl2pck/XdL1ETJQfVFTvyX49DB/53Qw3hsriA/InwB7F3mgE/2uBlD
kIUQCvov7XRpND5h6IQ/88NS3BIhlAu0h6J9PCQuK4h0mxkWR/7k4zx98dmtDopW
bBblgUxptwchkHv+8178i1k9FNNtCIPKzVNhKZGCohDfaQL5PeUiI7uGxHV1F36T
rIc7P6U+EAcTeZaxJdOcF4XdKmuOapkE/G4DRfCHgOPZpI/6Ixv2ussgTKnC3Mjv
RUwXWgDpvO5eCQ/LOtC+HBugUDFGL5YU+UADGNjR2oS1gw4ddjkyiBE6n3HVeeHx
c5/wCPZ3uE2TTrHnym7YQRBrr4FwgmTqamBrvKhmrLzrTZO9wEdVTEaf26Py2rea
hQJznzSYayRHm0YZJ1NtoTiW1iM3wOs47pRg83y/hbaxG7DEO/y/KV6j49Lip95L
SFd9TloSB8/mJa4Mgn8erRUBEnesVK6XCsqbVAq8xABsNt83dwS43BXLTNoqsH0i
CSAQjHUMPm8q+7k9metqTXctLCSHzUK6H5edTCGJBZ3EA7T3bQxNfwnMUwVSrIyZ
mnlui0WlFdSXl7o9BCApB7eph9gIASNe1SzGLbFRhdzYNT91FkWCKxs858QD8VYZ
nbzBTToaPbi5LOWmAWts+aAgbbLFioV6mzAXXijjDWldE07z1jczG3SeCngwJq2Q
skw1quI+usKRka9jHnrw0QsrzwOC9akqWEToL13zM7dkm/ODCeVK3GsJXJ3gUQzp
DmKDtDPFZ6XGvHPCXJXKcbmHm8PSIEphx7LXPPP9v9h+/8VWVlwS2uPf2UExRaRT
oJzvIwYksGtn0CgVwDNXuBDmF3oe3REgbII7GX1HStUfKIJXWAe3kCP0sCV+5SPR
7y+05Tf0s0fKyEJId+IJyVB5TUjItgrCfg0XHdn5LgoTodarQ0/BKTTrCTqS23jM
Qth77EbGczt96pIF2gExpSJTKw8WNqCwxWuYOMfJKNwihuAc9gJ3dVFR6PFP9vcV
dXTdyl+xL67D52HINY1Km74+VWMaK3I3wJF49ELrfkJllF+y99+exAXHrTXtPlMK
6Z9LIBE7MUWPQmVS+Ie6f8yZ4X/jzqhzm0cDT6B3fdLTBWSLmw/FemJ9U7YoggiA
C+dKGIUdEK4MhtiNAqRKupWIZ/c2H5wTjX2mzfTi0QUoc1AIFkKnMbFZeWZZP2mg
d3uXxRn6SOFsvE2stdyFjhFfnmsnEOyrRE1QuZRzKT2mJd67jQRj/EWXnvP5whPd
uuwX350SRVlC26LNDkMsiVQGEyBmYpDeeR6eB8v1z0mROMC6K0WdhzcNUKEMHXH4
z5ymqa5C6lCRGMxwmj5xFveQ8jM/b9KPHJWf7nxBCwAoMRTFC3EfFaeBwB7WeCf/
IQCQ4CAZSaFncvjI5AffC90QwgQmas/dbvSRutmtp/tEMbVVQ5j6kdg9lEYavRA3
rRWlH+F4Y6giJMm7iCYvlRpKSokpHaW+lWSSlEXVW+DgnRY/mqoEkQhEe3jqHuMQ
NRUGkNuYS+5LZMnM3T9OoufqBp88WdrnTffp1WOrzkIbns7mRGVeAIaxWj9DGJql
jLf0XymN5okpOAeIPERzNFgnSrNrwkO1iH1U1ppR0DrVB74ZalFFuiC6bi7BLcOM
Yz4pndFoflGIYbE28lSjqsPTZKXtannaJIw5fXYvxe8vms7+IBWUncxBj6aMnoae
o7HSDkgf0RwQrpljTNh35RqbmWf3U0oKwolUn9oT1JCTlu39+PTKmCnGxrZnP9po
GlNiPa6CW6e1sk9+FEGLVFQgPZgF8Own+S0NvYSOdBPXwdo+xlR12pYobq0tzQMp
hipzdmbcW3psyDUFd/sP8IFz+uksVSJ6j/S1dYVqBVQPJnicWi11/ZyIL3aqlcxo
+xM77gZ1TKHYQgAIOwtPnPV+DUmQ48YK7wGFSFN7jmMmVQt3J+H3tVjhYoz9KHTx
6sETmo0ax3qA7iTxjBtiA7ncik9PlHhUY3+jr3z+Mzo+1JLN2xRVuISx3NopWnKo
4X+M2Qakc4DKAV3r+/cKuTDDHwyOZ7EXCAqBRnOtZ4um7/bgST3j73b32ziG0w6x
OkZt8rLDCpxIXtyEnmEUTczilHeeysGEpqup7L9HAKCVA4fiUZrDVeov1IF8zN1b
OtmHWf3ctvqDRJJ2Z6rFVzlQ9uOkkOjUrPmTF1OckWc1vwdcN+zWlPKvIcEahwNp
RivYeQiPg9WFDqVXyKMockEZ8elLwUn0e4JJjLLUI7thePDRHSMImer+UeLzAmLi
j9kJbqC/d/bPn+zO+mMzmO/9Dl9/7VIDxTtpRTtI9hPweWZCLzSQVwzj/k4CWCZ/
w+l53e2iWFEZ/5Yy9l8z2JOoAEeDGfTJ79cuFJ86Gb4DADoA6NDSbwEJFE2aqz1o
OGoVz+ZPdpaGU2H+1uAq1WagdpiIa/17p098LW9PL7LPfA3gndGNmfbuEWXLTuN2
zhnwNqjwF6C+nHU66vNHuEklnOhRV74lkUFTm/BK5wgVCKt9Rk+O++kLhu4NyI56
J/RWlfbLBmlXinCToR5xtxqGV8qd9kDVWBgWZ8y0W8TmLA6H6teVLj6OC//tYQam
rPGIl3eTkhiaGsj2MkiO+hvm8NuQrXn9pRNQRoXSEyM/lHFbkn3swkgGHAYwv5Fr
USyySnOwJYTzTCVxjyUQ+y/62NYFOGUqKFtA0vkAMck/le978Bfpn871aB0i6Bv0
eB9MjpMv4VxtGUwkduDtFtNuwo8PJIqj06brJFjx9tQWB5vtfYKSQ5SfRc066rM8
eJuRC4JIgJLsOYKEqoqO7522DhniRSV5NZ7aHx0EWGp43dM7vOBzrf8mQg+yHx4A
NFpPQp6hVT6ZXf1zLpZivGRYa1eOLqOgg9WTy88C4BIXmsyUKtaKhPLGZc0RuTqt
Vc1u/nva5XVGYgUSCPqlA1EmuxXu1cygCX/ZSQL6lWKYnKAgUlRwW6euhU/MU42g
2MwZNutXoDwx5nUPWZrzor00NPuc5JThlMOohwUBZfQF+/JzQ9lAslFdk/6NE7zx
K0zeYxr6a0dUPIN/4HfWApm4FZMDT/2UZ6YvoKW4YeMuu1N437YJlA7t9DWCekGO
boyLjESh+cEYnXb2W9gDncp8G45TUK8ido+oa3Dy/sWz+7MmJLT/fkVB8pAoqjJV
ewkJwlClwsKKvaTNKlt69ojJjVtSBHliUeuzsf6UORcQiWUeUTZYFJmhb2AI+Y3x
Q5llzDuzYZX2VMELswOUPHxsO6jgcAnCFlsCIV4ZwSMz7i4yXvmCxh98GlxiQNBZ
IQBIPWmFQE8kYI+83tLXDttDD/isqzoZho9lnx4IKQTLXwADGz94IZ1eejBw3bAY
1IcRsG6eKiJMnJsFZCMZAWuuog4kc2wRL48OqMswVFLHpod3upYrS042xeJvpHhc
VD8Xp/L6l5CsvZDHXzS2h0oE9p3ETRfVfsyCji2ntZ0QfwAagly/doGQKkVtK9b+
mo8NQIfTdzUxAMCliItkQruKMSyAl2fpuKQsYA9y9YyUfHln64E1SGpat3JMXadH
3D9/xsWQHzJQm9npg7ZJc7equPh6w+OjfjxfZRLWaSN59+4+a8V+Bf2U8vo+nITw
TASr+pdew4fhdh1zR9PvGWTFlOVH08sM2Aek4w44SEDUerXMvXMJ0MnSIAv6FjWr
G45IMEJiLXmKCPcNaCQrXgWR7f4BinLwnKmYiPkoF4KEefngPDh3LygJ4lyp7ali
L6TxRPQYL14QDkL4EcejftN5qsGTfdxaok5vca6bvTAelCHcLiRuzVNA6ra2/Pg9
Aqsmi2Bnd0xSVs1g8gMgL+kuycFOPo8zBU5taTmnGsidcSSA1zeSJXbr4LxDmA+S
Y7zeCZD9/MQPGjkNgY4BKvBkO1rN80o+BjI0t3P0yRESzhS3sImAKiMG0iCWLv3u
IRJrcOuN7LZL1TVlcUuJF1lautmjoFAe09AUu08pZIiGYToGU9On5HwdA4ecPPQq
AhKyyA1mechkuchRZkvT+6vuVJQfxQJmgmfVbrPRq9Ivd+LALVcmARIQXNpZRAgG
UYCMfqnB+DJ0MthQPJYXdMRfKAE8Shq4FyCnPVF8GslC5vaJqx49higzGknSduV9
jtPirFOj/5hm6smVA6FttAsahty0nMCkzXfRUIv+5DPFxVLt4M6DYSWn1vLw5o72
Ky7pg+8slZJFEUi8nu+LkoxlZxhjGc3HqGBgdBUDe8OaroPqI/8fiXn5V/tXcU0V
BLFFSueZ1g6bt+AtA8BMnrYZuCGrA0Jaqm4srhdeKLxfJ6YAyjAi0gJAofXep8dz
LdihLc7wTjm83Z6h7+1u7hR+YvZusaYRSBc7jbu8QBV9OsaIddklEyHBnodgkL4l
7n/rt/fesqjY6DK5pVfnfuv7D5ye9jV9j1Xi+Lk2rswjsIOSI8qlHM50tInooywl
C7MZyxpfKCrMR3orLP2PxXI/fjZ0/eQ/ORTSbWdrnhzc2FRoRm0EumRXXoAxml5M
3Amt+O7w+CMiHxhH5J/RDlrhPyEEVmmlIW9sEErb1chHk6UfYr87QnW09sbGC5i1
8sm61bELNAQX272lLLNvVncYa/0664wvN3BR6x80ctlmhlPgULWj91QaWyk2ysbQ
2syt9ju88eqNu93ulRtNm0+oXmOqCB3nWjzFoaySCWe9RsLbH41ayTmOXV9mMQrO
B3hAy6U7bTcKjZG4XYBYK375osusjmchPZnvRBE2wvadWxfs94recoTQhd7LA9r1
XebFfFeLTFqDy1W0afoI4a8QefIICsuWdIFHPhWzCfnaknf5VEiPxsuYDBIIkJXj
cFQtCSAVeTru+8/m8a2ZQNJVCsw5br2dlZD6/M064QSes8eQ4tqt8TmHP6kk9AKt
erOA9X5aDsMRTAJhCcKMXeXz0TIwivt4O3Cocb+L9tY1prWsKoUceVUfx8NiRJig
is72y7EkZ2O6gklA5818qGZMhOpTS8B3f9FO9E/9+yZXLm5gVYAFRnR68HxPwkts
VT7jlCpnVXyj7ysoth5v2WAcYRtkOrKlrhZUaEAanYpP4AfUyoz3ozvpGyIK8W0Y
14hi1yTkJRBShh6KznIKvVrGZYogBCPP23BKliDVeowJXDaYMzP2lFcrkEUo611B
`protect end_protected