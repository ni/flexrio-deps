`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
j9eMmSPGcKCWAR9PvkqZ1R001FU8QKTyJzFqNLn+qur6INyYDE1AI8LWcxAzfnTc
IpZG7ua3uuk5/kQKKQx8ZIPLfmv6H3t3eWjki8YIAtY/d5E7Gq8Z5mNxMYRzGGTg
TCMm6oOrOTVYlCXHE0X9AW696Z7UGfWirVibl8hs19hrFdeZKGiGht4r09vHR+Gl
FQQmSObM5aSK5wu5KOrK5ZUKGHyBhjnIQO5NnittDjOwxV/57nHVg0pdG6JUqyvm
tEgmCY36RCMRGWN7sekPtNHjqpZkmYrVX1T9QF3h73+8ZekZYd2xY2hpHHGYYeWA
t3+Fmb/6NUmoP8+Pt2hI6g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="wX+NBVcG/A5ruHK3pkDqG8ZVPdOz9TJPJ5saXZYSeQ4="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
j/hqWUoxjK88VtH4QmjIrexFOSwtsLKOZ/LCP4cmrqgzmR/e71apdtoL+o8nlfy6
eZxDZMmrZmJGoazz2oK6kz7xJU85UCwNc4cxAsVxNdCP19vZxph/nCYZQ9lUFkLH
uLBkOeFP15CD3jG5/dp945fHP13J9SzB/L9PWvDC/gY=
`protect rights_digest_method = "sha256"
`protect end_toolblock="sqDZkaglKf+bDjC7VKm3lOELrT2Jlynh4UhPg2J0Q70="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 55056 )
`protect data_block
f9kZDbPp4NLiAOFOgATj9W35i3s4a7wbt9jeHjHVcJxMoXY8rb8laqS5bNUhXGW/
MOc7UNc1VwolqhkS7G27SLamkGClZZtXSbRcN1N+5kZpEaBEj1343vVznnU2Dre/
WS9HsWPXe5g0wH0AJA0FuMwn1XqDwa0faTwv+9s4qMICs1fzJixbHut7car9Ywc1
+XgDHgrGRva2JAzaQnf3sYpNoRGdcRFA/OcLIwSMcgAGb8EfP34a2dC2DE+RC2VQ
MII/4zjLmDLBbyoQjQeliWFZxpavn+9zvdKvPzJGjr7t4+tMuJeY0ShA/uB3lmas
0vGxyaH+ZYLNQjEpc86B1RezQMZiTdeNq0UeZwbJsi4vxfsoZJWHbYQ/x6mL0rc2
+vmo2n6SOiatLuAkXKcZ+AzJ0aTAflqOBlT/OKElGl1vJRxOwmqVSmmYgtbOiaT+
leaY7MtzWoBULeud1DlvfuMXofPVaHCU9n/kpljN4+PJQO+Hz33IQdlFHNlYsxsK
Tn6iu6jol9JTadhKyycfpZnD8mb3NkjCHNoBXvy7MP518FoQjj/aYm/busyg+U3I
rdLqjgXrVq9Plizgmj47joRPwg03TfzurgjGM8wN5GoRCD5qStcdIDHOYQx6Ultf
M5q1utEnvq+EZRI5Any80NLgu9l1SFaCt392lfay+V+UstuGMq0YwIYa6HvBzKoX
wlibMBZQsD4vnkE3TSd73cBJ57BB/X8WT5Gc/b07YVdoVRv/DpKaQ9r6VLO2ekQA
eD3TfPmTOM6bpoJnOwwNxpJ04xrgKgC3Dj6F/5SsxKNE+udoogqsrzPozeXYkB0N
UduUEaxGnCuGeDW6Z8z0RdAr9uer9ohqQG1iRgE1woctx96GzzzNgTnhneukIo6E
AeN3I1vS+6FwDngOEoyxTXoqD7qh71Mq9syKEVZfyGksslwdUitDEsMtoudq+8WL
edOyDJmgn2xZq33HZLzsmcje2BtF/Nkx7H05C0HQwS5bdqB6KxQNcDSZ6Nqwwpbq
dxMWA4kFBg46amCLQaXFNBhdnLcgDKPeo4DgsknwiAb4GilJND+syl6NUkwo4S4i
/PDtFcXR+2++ccqRoq/o64USYTLeKx0aWvHySje6PjQv1xnRwcsJbUTvK9cnyyi6
0KOLbf/dqbNFbpYB/yKEcDeJ5mTkTelm1kq1PvLy6Aw0ue1FbtaJdDAyMEd8YSDr
S1j+Vg682Psy/mCwxDwwiiYG4OOZAQsC5Kc8AaLQlmlQxta0r1N8b865rdpSiDlg
eEKhrtYBFmk373UJbxRVaL0FKpbXWw/Etz9taicv1UiKlOVC6O5f1TwRtWBiAfkK
Se1F+Ik//TQBG9oeWC6n5GCVREGdN502BhY1tMCj3uDKOLZyWEE+mDyP17WRUNHl
maFcSovymrhbm4yODjSDT1+BcFLavhGv/Tc7OIjo1q3ukoCPwA7yrth9ERFe4x/j
Q9UPT+MuAMoY5jDEf1KOoGx/+M7yPNNBdiorBF9QHaK37fSBwW9bZxkVE5BsKKzb
nRKFrHugKKFFhkOUEIXvqvg3UvmVJX/qzV++dVbxOhnH3q1lFgD+lii524iwwKch
dJkzfYbsQv2BIsmy+fvJCseh8eaAtkKahUs1MBEartNJCgb+n5IELinU63Rw1BeD
2/qvFufMx6d6GhiASX/ei4brUQdU6vgrajP2Vqp7HJSho+ZKD83fOHSiRcxmq7Dj
Wm0yMYbEB9el9KbTuH/2n1MUNvTvLA7/oBdE+JRfjqmuFnO+LlITRKj7PKyyfqpg
b5lhRgpxeAqr4y1BdWwn3Woq8rWmycUtmIWfuYXC1PNLzDDi5f2tbi5DHz+ovgwS
XZxWDCbpgoDjomBoxE8SN5sLb0S/P34OaHoluBQk3T4ihfnXIXuLImWOJ1tLFHi5
eIUUATXPzNbN2l6mX42S2Dhlzhe8efOEaR2hPGW6RzDjCBzF8mG3lm2xf3TslzPx
125umWn4dERu4dmoeQFzjhtUFoQijVllw/5Of03nc2PLit+HymmicdAfCrN37KR7
OXKzcgrk08Q27NBOJDE7AXqqhdOnqoXbjScO0zeP4LZ38IM2h71bBuAgIoAPPqFc
zoUi1quPlIHGLuxEPdVdc951bEQ4VD8CrkIFXqIgolYtAFCb/hfLDvSJMcbU1gka
LbsSq6TsMoyWI/OFDG6gXipb37xl7taD1cub0hdkc+MJJX+Y85k7lul2uVPRZYiW
hp0UT7HXt4zjl2RjTQ2M46k16D+T7SasveYfghCjz90sxPtct6kNglaNG/XshDDs
yjhWeJ+rDdntIfEpOVzL/FzrzvcZGApvwjznI4reS34hU8lCSm/m9etsFUDaokXt
hm7OtIuIi3HrQG33+JVB8zSUVNZO3Q9rOLWnEMDAFCasNitZ1s+igleyWKcc3ApL
kqsix8ztwGSd2ssC2vX7axrPwIckGIWGKo8imzUFIMt0i7EorPO+GHMTpxTzIbQb
QTlTJgnAjbn10M8PwyC6rtLNTHrFJzx+igUG6ynRg5w9sYkaXJTD2G9q9xVSZW4V
/u4m5dmzDEPaOx6pyx+wjn/jtZSb5FJKdM2AGniVTjpovKTuYlGEjysqeIwAc042
/YGXFBOrpm5ELIAYTSHSycfdWgeTjTszIxb5xiuIIh5VcJKP8ErwddMYgP+EG5RX
6wU7AVBwEgC9DWlwB7Qil6+ZOVcXE9L3PZwSPcnJDI3ahjNGFqyG1r8PFIOyfpOR
HQfDjm9xuP0b4nm3aMjVa4ky8Xq6yOjNVcukYSdsDvqO2CY2Hw+4TqCITtvSmcgO
cKeIzpGtqGtzeg0BdLgLRKrxzx5DJC1Zv/DTj2esv4F2onzFD6Eqggf5XDSeSkDa
6r5yUugCQpuvBwPPG5RT7A3BzBWnZNgwrGQScfvoAKZD89Vs7CwRwn2uzKhsVotj
AxEMtH8Kk12KMWjwN6SXPz2ND08yIfcSgZwGz2/7PUElHgXEgPP75tG0d+rBS4td
TecMi00rGwjLc4wnsp+zrUj/M0QBL6pdDRE5S/2Ngg2DPgwuAkynj2iOUTWkmwFc
VhMUhVQ3+Q2teOWyIGBbPdovrZ+yNqzsgmonE66K1HpfC36kJZ3iSqb/lD3gcGie
ftja5frFSOh8e07RHc7yt6SwE1xdCcuz4/huqnJiFqblXHAdz2DP5hSJh6Alca4c
fRZSbccLdO+grUpQ7y/ItbqWAHgA6TkCptPSFwEVrgxDKwdUd9FnjUVSWjgOb8Pa
57pdLOni2PAO6j1c/KE56Ae8PaJkbifOw0X1/6n3Zq882aku1HNOEu3DnG56Clm3
jYm4rbpXF8hppPv02+D9YMc3QJsI2ASYWAlIGELTsWhmO9Pym8uEGvIuTLUx6fsH
vt7xwzRkwR/mUo7Nz+sH1KVXIRve56GEdMaqCI+RtlY/IQVeKieADsVVvuwXaBFR
+LHJMMrAAwAy2FTnJkEqcnkMmI28ORHx8yM0OZWENxCLe/g08GlXf4U9nVUhPZvV
R1HMNdgzNhVBAkjep/irQXGq1hluIXPmzWdJ2L+RT+/Dd6sM2GarxqniPpb3H1Bh
Crpb3Buaxq62+qQo8vS79dbmTajn0zxJJNj589S3zEHp+B2GX5Ofd8U6yZ5FNOFz
7ahPits/zGM2xiAQoxKGMqTo90gP1JIBWfHe+WXI9XE2biSqwKmvsXdgknlTaQUc
4R7Ke5RR9QaLZgHO0WyUii2vSuzO52FvIc0gvpToR34SSU0tsgiIsDHVvdC4TEME
Uk8dmwnYfwOwJrTYvnOEX4dhnO2RAZ+lbJv/QC+5LtBLeoeVZXxmNI5hM7UBd591
0yzyrVxrYr2LnIHSAYFp30XVqC6YtaAxomXeaKyFZJOqCiNVAZj8s0VxejAVizfp
5itvqdb1JWKkI7R0hbh/VaLLSPAnAK81WLklqjYvnzEIyixCT0IS0p2gCcrzn5ua
rpyAL4zTRHHXA2A8R4k0Op1SfQv59DCdxCtu+XwtkJA5rSiMcTXjsqpFKHTR5F8B
FkNx4VTYlRS6fnWiWo8m715O/2gwoN0lmAGIL+lEUMeR7P6eSM1kqflHb9KExE+S
Y8jaltvpQh9bilUO6YxJHbEnopyxOJcpIcEyyF0HpGVLHTLz+dgJzMHrv1nununP
OzlYCn68lcScqyNi79B+H8PkYQKUcX0KSV7v8BHz4Pc5t2MrqW+ObnBR4oXeur3B
N3DGE7jyPRXgN1k7j8hERbBFI5y5FXuENWL2h4cV1CDijevDiBc54cUHUYthcaxJ
jA7VD4XbBTtwAlSYAdKRHSpNCLYxJckbX6F+glVbBG5NQ8Q6w/LkDvgdvLRjpBGG
6VAcxWqjWIx8vptqv4WLdHCNU3e7GdOpcvvQ9DaQYbK3fTbzGyaWGBwRouNSMa32
tPg5Bhp/6LpKQrnopjTZuXXlr5qeap/FMtIagFzhtz8QioPrhg8hm1sBH5xyO8HG
Vjvqs+YXlj3X6wowuVnz3pkqhcy0GLa5CMrHJfr0FAzA4HyEscw6yhFAWXAbq2Y9
XhMXRkWBSmsk07rm+iwj4eLMtBrb0k28MVptEySDWM1yAbCm2BOAgEWtQK2J75tO
pStkbMCHqzCB2aAOv2Z16pHP6S/GLkIeHF5jDhStH2iaUt+bHQ1wx2Ny68pQX11j
ArOK11P+sr1UzA8B3hhcpzugYKragrOi42JXlqQXZ9I6Lq2VkKW/FW2lWmN01t1D
H0JEHzzV7tWuOTtOelpl8d4oer4Pnke1cxY5Z3BzGxp7Jdmcvo0En3sy983ov0B3
kwK8dCrczqVdHCwcF/Ja2kUBRV1m7ZCHePlb3wDoWqS8iYO+jhpkF9Li8ScUNOla
rhSRjevoutoNb8Iz2Hl3UcXe9VJErmrQvr6EK7Yi9AxpS8flRrWsJMCzp0WIilH0
KQrT9ffFmcrnoPDK/r38pA35j/+Fum1BG3juxbwpCQMaHxwzsrTgYAyKj0DycIIT
vBkDK6tdzj//npilTuP3vU4TskUKPH8Jti/j9hhUOkN3a+6qQj1cGneUeCjsKbAl
XjVwCWGeRQ0dFKfxxQ0oMGYil4CdvlxjnhOiQQlzSHfkdHSmvxHivLFUJf1z0ePi
mRr24C6U9Zi0aH0oAF7C9CS8fDD5aoUJegebUJVG0SXQU5TsObGTsk4ulNGgQzBs
0W+r9XBpVf5TTfehBi+42JsQeJdyB68QtZhP7mV9NZc1xG7WRAk/GftB4385+9cK
UMuQ052xApymUdUS2CSKuyobh9Puofrc7yatAA+rkam1UMy85hZP/IGua16hh+jY
KAtFmbljcsTY5qE2J22iA+jF/vhYgO6K4AYda1AfD9qS4BXfArNs3e2SGniC5eT6
9Woo7X7q9aWpLHpdgIioubWfX8sn8oqc8JWeau951F2JkxJPbCDPuZLVWRLut0OP
6VPVPbPx+1XH7hJTH6B1G7JKxQSEfD6t3B8LsoZ0W0W1zHGSxRDI/+gzEDuWxfWa
Dy1X65IBheFNZkkODzQA3bzjUIhvpi6HMY1YhjIVcRLXrg/C05/ZdOqiT9ZG/Csa
LCC2NYo5V31oAO11DGGSfWvCXsqGoKMzTgrWc7Xrm4KPVwZIcL4vJOSteFHRBShq
x4yWqLHEAd/oBY7eSn1mUl/e3J7oi5lkKr0x1cbjx9D51WMf0wAmruQYbhNrmoYu
CcTq3wewnP4wM3/K0Sf/sNbg0idv85IP+1T0456GXMR30onOVgPFCVkJSMA0zS1d
NwU8PV4Fe19UQi5p52rB25zQGqnr6+T/55IiDyFidz6hQN5BEb/e2xaaB2YfDaf4
aWrcobdgfIfsuZY4vnAJZV52naJIwCcl1to58+4bx+PyC2z1TyEYMwdrvdw/UsEh
0q+pDmqqB6Gx2IdAupXTRBssIo+vp2DBWgbhOA3/Mo7OoQNGar0DnvYQ6QrK5evl
djyjrikN7nH7bSKFGae8aTiufb/Sqa5mkNZY/cq1vp/EsZMa2Xx/UxUMrvJ2lAth
8N3EZMdpKU2U8+APKVrxAXgqmspl3+0iQd1Y7ycMcC1EvxO/HWNgc3UiIjc3ZAFz
jEt5/wFJAJiZfUVBZj/sl0D6RH5wkDnv6lWW8Er6xsQ/BJxbmH1or7W3q4kaPaNw
kZNuGJfSov6Nw1l5z8Xa9LtEQpTd9MV0GUNF1QAqWF9QGxjzyTZU3G1mAVK+MuIU
FGoJSEBW+otE9YLcWuGZjEhcEI/luRUEQbAAMdJxxN5KLL8X7P7gBDNvdZSy5OpX
+lAT36nYiaHucNl4/qb0LQnqC11kL7U/mbZAKMmzKUfBuoSTa/rGgkx7WrjgxtwS
lvcdpoonzSRo63I3jvYN9k7ZkoVTFELpa99OI0vX9EeKo5pKdoWSyQECpdr4N/8+
ChiFnNbIuoAgIK0GmKCrgsmYgYehiL5Mp/2CuLRFzH/Qu32OJpNResva6nWtb7Qz
LqFSmuVmULYUcDzUzQTWC+4R2TQpgsIZ6ZE/2O23ZDRIzdir1j5cwyFfXFfvAUvb
c4IuP5jRzcmU8f72fBtiC8u0Ecb5IPDiP77zLZgty9S4rCag0yG8KV9XcIOl3LEN
h8FRFdb07SB5nHNj8lvbF9vtUMjelAYUzvZZK9I1afYb6A73yoBlDmCdTrlmkMtj
bYjG0AdNleUUKDwCz4YcUIeY43aNm3V41LPSOUTZVoc0BhpGCwqwGCHX1RHW8ZA7
oWGy5ShWbPc4QpX8weoJgrXw9BJEFFsybmKnXQnD+MFj+3sZqP9JAV8kFaU+MutH
nQ78FUnCkpQeZzGTMK6i1its1c6Kq7vIRgYt8fqW7OSWk+asB51THQKtKN7L8Aqs
w16BkIp8zMF2JPz7baga74oIQONZJwYQQBpsi+3+Y2iDgQwJ3jSzPslNJ+e4RHO3
h7Rbn+E+vKyWhoq7CwbWqNoxuBel93391p8YhowmTd+xIBbyq/xp85mDV8p/03hA
ZXp1DVP3kXesBG6gL75Djz2PXvxVIuKJywhwHVnKgYKI0r66WMJCw3x2qrPkCorB
+QFPzHSBV7siYtIvdB2g1baqJRZ3DR7zI62Uu01SwR7kpLbj6qfDFygw9Zfbr8Ne
Prmrxe3rai1/7TpF57ZSMM2BZVg6E9CyfDH2PvSGtX3KkiKfPm2tQ8lIJF/IViJV
1uwqOyW+2EaRxJYw+SLQjb5CdONc8PPWXGIuaco3OtpbYp6WpFr8Bu5YM9agxWEa
VkGYmqsZFyPs/xqW8LQqTj1HD1sQt3EjtW+IX0u8mFJ0CXemusX+7s3aO+ksOdhy
Rg719VAwnbUOuNyPuKqM4YIbTBVtj76DVBAnPKsAab5egFNi5yP0ZdRuyX217ycR
ieL0yBZuRG7JpnFPcL4s3uKauAAhw5MpjWem2p2S/FSmJHA9Du4WhS1SqJkE/Xia
Nj1ry7sYonMv1EHEYWIbA3syM2sqSnqR9KW+E9opwf95LznCpS1Hr5HCgIaYP49i
eztwI/72wslLFvqgRZyw+vJ6AsYb/ffaSSAz9b+N8uyk6vIj2A1wPJYR59rMwBTb
+N1n+T2BecqB/ZteBmvu5ryIA+fdZmG0xrfjAJKAoDVo42uOSv6mgDsRts6U4uiF
/JYgwulN1p7ZgjgLVjiN0rmcmY8jM+FdRSEeGfzQ/yBd8vimUOSWdDXnmpBEx0x0
AAPPDmgrSVYmrwyMsTKTFJ5dc0cnW077QSaR33ZNbyuKiVcRqE8EDvbpaRr9Ey9W
dAArrvIen7WN2RM5N2J3k3xMJQ1/Zm7uHE/dBcdqU2vQYL+WtOSIo6o2vb/69mcO
P/QjRTxs8v+aHy40ER0owymIxmOER4RNXM64ohoXKeA3EHRnH+/j9iMBODGxHDuz
mQOXirFNeOg4uCAUoT5MFEC13d9mtDpxpD2D5fCAFUU2OWIvCPwqhdTSp/2BmDVG
tyOAvxqa4xLWg1F8X7NuC5CtK2qGFmXROKfNSxAlsI2B84+GxdCuyc7ZzOdUA+JR
yIPW7gHvEduAYMecdYNJ02+/mARwXTOuF+h8aiHK4w33o28fU884HM6VzZmUUMzY
NMKYJfS77proJZHG1bAG84BKZghiuhyaHaOtFMHyHyFpfm4IWDiGS8Ze3/NzM/Eo
FjYtu6ZuLvo5PXVL/G0NHX3aQbijh+DpyvEhD5xrVST+3LRzVu71vM9wTDZ6cBXL
jAN+ZOB9/16o1x2UCg08+Xis4FZTfga83hC0jWorLTOno8CVLKn/ejOkT+Ox5GsB
3N5a5gmrQWAG2y9DqD9PJASBh1g3forX3Dck7jTzVJqohSQwDyyGRNRBJnTqHEq4
R4N31kHtNgpU++dgUFpzuZUUbBiZSmwREd6+KquCHunUsg6CRZE9GtYBGMhO/paZ
kjX2bMxCBCz8TSBiQcj7d6OcfUH7NUHe6kUjSi00rjgk5VWMW4xjaaapD3W+yvy7
CzCrQdQFGOUYxz0+355caA3WhfUQO3r4+xcfLmH06AuBqZN74AFvodbhIhIwjod6
wGs+Gw6q6CLPw/paVfWGrU9TtTPF49ROeT5NJmwj0LdehkfbflWOHQTnYzfWNMQM
ycqvXx3q0G24VaOU1gr4UbMcY/JdpXWYwJBgUGLMO62bolLblkdphXqpfU3CGtiE
zslrXizjNIixe+kI53ILTSClUF4U4wvDzuWiGyZPgBQq74DZeA0JQ/KitSek+fDq
HVyXP7Oob5tqZ2skNbQMAVtd5gQ7kO4LoZ3+4rKiGsxAxzqaqA5PI85bH5l8TC+T
57yG5hZLH97SdMOLSFKN90hskUssPddKWZigYO12Q1d/4S+EKnTY8SCk7HrVkalK
wzZcu1Al9D/khtbX3yX6RiVjXlbz01bITsfXFTqtIpoeFGQQU6ydLZXSVgqA/Dqo
KhX8f7akrSoluuly0M25waH23MTLyagwnf6qceyy9u0rvjBVJ+mrgn9bYJXO+DoJ
hzsuBMRqb2X/wFIp8fXay7rc52Fq7jyg+3TjX+RFoSGrrrhMh4MynL7RWa0zi5iN
+BFG3WEqDVt6eNfwANpPMMmlaKbBhKSXpOJtH47sofnAVA2bfahkujtJLgtLsWsf
/E8NLpKfvR5XyfHwIWkQt/4KvvgXPSaW7T+mz0VKiA32p84uZUn1e+hurvCMTkQU
yPnTu8qLfLX4oeiUQV4o5G1l9xFqs8N/cHvyhCwZbj02XPQ3llHFK8IsPPcsGn/w
co4v2s6lFKm34nx3htrwdXnCvoifGjg/MMttgcE1ZCQcTzuiZlegLwVUAyYKj9Ab
KxIbkuVKsPIV7Oj4m48IlF2h+9kviR7rZvywHFPOZ/fy4fXFipfTHjFojDm2O+ha
r3HbvlM/LPma+n8B8gzXx6KhwG1NCE/ktsV/zF8UYn7etpYbC9SsfNInqXZXy2uX
VFHkNTyEEa+W9rIshi2CKeuuZAfKZGhfj/GxvPLXM+8xd08IS5PY4nOT7tu/TaAi
EVTZezJsAYRJcLEP0yGy2aLOlousQWmfTea7vO9OOkJeeCn63LGfPmip439plQgp
CJFkKA0/kcXD+kxbax4m5q750I4lMT/Jbet4R+dL3tFt+TH0ArWGO0/BKCc+eis3
JuSjfsVwkCLZBe7fgBPSe2TKrLMjzwguPpatuEbRKz8LAfaM/35dxKTfzRSoz4kn
KpAgmE9BOFIzNJ3LckiVP0x4Z36nb81lM/5+t4+b70UuKtHpKvMXF//yy1OUVlTy
6tkbCRAtWk8M/oHVAQ0+yOAAof49r5kAnQjkta4Mj1PyYcF59MPt2LfWS6uPYnVE
K6K/8/KVSkcH56s2NEVZCLi1vA1+6am/E/cLY5wppvaZX+6SGTiUDkI0eUcwjHnN
g2QgC7CVRcW6LLQlkR1HtQJ8l+3BNSBl+hjY45WwrMbT6wO69GhSo4dnFLr8lYxK
tJfIuY56mvBL68sxWZ8EazBSGjJzW9VxsVbaZQGVm+Vt1vY5gAunwd+F+MdHDUl1
w2HutWvN8cXsDVd928To3wEWD3Djjz3slwEGJCPCmarK2SjUVKEbdGExPkXrsWug
/7wmX6m/CFmIXFMV+UXxJmhc9p6OitZUfFNLjZrSkdOX/ePmqhilnBLDlJNqA/gQ
ff5XZwo4miZRu6KLrQwGBn75DmV5WUgJPXnAJygfwFiWpRADhOwWcnaEbRagsrIR
RJ+o9MI3MsyDWSJU6cWql64OHg23wZFjZpU8QlkPtJDg4nI1A4p/14ug3VTT7GzG
dmIz2whqCR+9IBuh0u5s7xW9fj0UxKLcnYZScg+TRfGPGI/ty81rMp53fxPhafZA
O+GUETda2vAMA8mQp9+W6Zh64uF4uGvePX99fQ8LXp7EhP2SnuRJd3kRMiIXamcq
ajtDS0rpCqcVFhQWEdkQTzW2Abnt0S2cZDpsYPjlowp9/BWjSEUqan+AjFXkZmSc
TmujcM2QDvnhmufYpmWr3b9OnitxJaK88UpmLVI83KhHwCE/1eihMUC7UpoiWb2Q
JLrb0XgjivPNqfwUP1tldqB0IDR2r+VATFxwdHVXtoXVNwIpnZWxUX0B5QsKS5+d
I/BHq5YtbgVYKu14mv8+TSg3yQpzmZjRLtgpXcSsgOB/luRLnC8B3uxscRCYLHhz
gmYnXfsygQGRC/CsB3Hlx87G0oBHSo7gZecROcoGLZ4SD7UHzB0oFdnsmxDj+DYx
O1szGURB322gTPWDb+6sfZRGx9hELbXbyFMH7ERrhyjR9ZExjQ7r7gbXO3ETHSF4
coFIQgWgO1F1B34hwjXnKVPneopq1b0ftFed5puI0s9cTBsm8duUmbW6yr5jibH5
jz2DslnYKvBBOHL3XpPwPMdz/o9epoqY+UuSb6QbzNf9Sgi+ajRHfm/j7D7uhX6E
TMQBsbO8PVGxPWnWNpqzu9ao7hliKaHzl9KQqYLoLTyJOX5NAGJLO7Skhh6E44AV
tfhEAFrni/9+jwdTrkcEG1smFuxQUrSQ9WB3vOC9GsyS45hWQh/BQlhHHF9wjneG
+bd2EsR6R+FfeoPf5Pwer5V4H77Ko7LvmPJBZYKZEr6+d7taolsrI3c1vJE55DfA
MsL6YYSS7dZdcTKjSXoTJj5gxNRVLgfzonVtdY0lNocUtvABM58EElca5hn/Sp5a
o1B2GARrdnG49LHQsllQ7aCLnCEwwyYkOg2uz9/uDAK8vXT1WxWKVaQAGtdjet3v
QdR7MHbhEGd7I/6RZUJbDTQ51JMsmD6nFeucwa7Bn0l1tfCSrM/SSxRF9lH1Y8HX
7J76MLG5Dm/3um6jn9Y/oqtbZuGlWV+5SrWtUYif8YKHzMh/Za5hYr6yjm56sJqY
mqyZk3uDdv7yyNrpXG85wYVN/Tq+eacQjzUlJzRMtTeEIJWWyqKTPLq3RZPSCRBM
AuCCTfOEf70KW7SjZxl80oQwkS4zoM6NynNv7YYh1qTj+RByZDaH0QMbbqVQDebW
lMwcDqryfnai/9LrBgeMHghPiLzYnfNQGTOmvGqyQUyUmbrA8w2G5R0pIogQWzlH
kW5+NuI8h9mdus1Uc1jDEkhQ7Mc4+LqTpkm3aHBLrllGVJv+wQN9MRiPK6ISz6Ko
ypAM1iEppZ19MPql7R2ztFqyO2CKcGCjjCsf8LCtrljMkrhpcwyHWvI8cZMngyCg
sxQ6SkiAk3ZeI2/whLxlIJE/IJQfS7T++hw1QzhHNgBOKQKeKaq4VyGsskBcCO6o
5c9DetSlX+7zjJtzxlDZnPRPPT7cpEQmv/DqPXtQVbXjLJ3H8Mh/kuRXjDCBJpzc
pBe6iiOo1Az6iuxWI/RdI6aiCIUilx9r1T2/p71mAU1Y7jfyh2924tWSwYM25p0k
i1Ky4EO4BDm4tWRgxpuUFFVzs8HP2QH0ykwuGD3qRlvAj2K/GMjMcc/+bUOqN7Xe
EMl5PkYrIcAUmYKZZzTLALx0VaISNYFpGx5ThNSAwwMYqRXMQ24CZCTf26Xtda2N
Hp31Dlrrp8wg0D862aKzfZDzMQlYhfEbCc6xG+R4JPrXzVpLyyt0vIQ3XnXLo7ex
/XFideD00ffFTlZ3/FNunEhZRIKLemGxsBh4Rtoafz2N4kZIf690hecuwI7nH0cE
pI2DCkp/BhsTDIP4FfFSOMYuKndrF5BbNEuYH6/IH2vf/9wMQs3/A+7beFWjdbup
xwCXPoipkWIt5eBgMYSdakZeqDtyfY137Uq/9XNskstndR1B8Tl/5X8I7h50fnaj
iGuqQo7JBTy+V6C29g+QC10dDOJbPM3aNpiTpUKXyWoVdzjPmuGYTYW4w/L2l/vV
lgv0v+CpFTO8uchayQs3WQPOSHiCBm81bWeRa0XwhORgrjTwtKwq9jaIGwLiUj/3
9nSYvtyZwWAeh6siOw014QiYWIJoCbNqnX1AkNcEWf0H8If5H0MmbApz2B4+KK7a
jKIlZ2BnzYxQOfDYKkRApGSFS1wpN3LKrGuAE/QhG4r4+k5CobS4hqL8pB4E7VdZ
zs8soFW2OYSHFluP0jljvy2VeBIc8hsE+rbGU52ESJYZ6wS6RGE8A8GrLhbi4y6X
ZfLTykfH/Uc+FJPl4ig4mS5o49aKzdojllhzpSQWZaLa6mC/ulqjForXnyqiqyUd
h2a8Xy9nzOrxAobJx8zZxwD/w8nH/EG1dZlk3mCjGoJYhTVdfJPhNvvDuzcNbLuj
DGy9NvD5yvFkBFQI4nPLDFSf359GCXg8TXqVa/eF2zMkQSp48u6yo9CGFfMZHyPs
e71hrx9PMyP9p5fUKXeq4kDC9rIzVyd5DsLjO5sLnhIPu/nU+bRpG3hNbKZkvV3G
VunEhmVY/KyJn5JTaM42PMkvOdo2GAZAF4sjLmQG4kb7IYxCP5ZXEBDrqco3qnt5
REopVkEvXKdfC8/el4IHiz3c8Qr1uU5/8ZyCZmnO6b6jzzCqUnE0qWONgHx0CfSP
rnN1Emf5j3OtDq/b7cW9kDL4xBh1fJYPPQObSHabLzwNTxE/brPy//QoPIS/2aLW
GnjVOmVN3G5N2hFZT6N3dYxrgfFYEk+ISpeAdOQusKkWMSOIb7Hg2CPoTLDny9eF
V+xK5jC69oIATpbv5eC+JJYudoqEN0+HeIr0ezZGXYRcoPZtvHQMSCg6okjJ3dtc
9I6MS0TxvOaZzsrsksas8PPwaJZZfTPwT//zkqmrIE6e17m3Q5sSqMz+HDpqofzU
HHv1B7ildqdR7Qe2gKTmlqlpdYphxSjx8B7aBWL82OhtwDb+0NtCcleV2Nyiaz7z
hF3RFpcMxEjPXYJiOekndGm2Sx6f2jSf3UPULJTOR2u6LGYbQuOX8pRl895EP9aw
mYRBt5pueBakzbWvv2lBSS/g68MtKkA8RPQz6Maykzt3e4DWkWm3ehSKw1XimAiw
ABbWvKz5k8aRa/OUZbW53SKD3sfIzO/yxXciC+iYxHV2Yqt/vYrUlRGJARJ1gcqE
j6wvPYTSSY0VUy5RnuPPYG7xIFYRTRtNqukf7tVoJ9vU0bEfjfROBWJz9arQESWl
B69eeCfPEjEz7BzSBLn4CkHQ3XVXPlMemTxa9rkw7gVVmuld2kfRHJwolaXGV9EY
Xw9w1LfwAIlmJzrftyJQdd0fyRwVn7RBLHDOq9hTnJnklgfwf2iUBHcDqm2t+eKq
I02iG1sQAhUBD+10W40aQqNgImYfR6/FJyksMHtEfuzR6jIodGJLG871gH7O926l
zdp2qR3pFsYJ9wj+FKW9kgaOKd++PLSCKZip5SXIL6tjSxoCT2j3/wqQK95cHhhS
RW1GmRBGTudx9hquJRblALGXkLaMcr1Pe5eiF8UUPmqbHeFxPSqCbGqukJw0yKMm
hggvnFk0rISofX2ONeoW9RcTNaR9nNJtIh850zbw0jjWnPQmKdzGq3ekM/0AE7bN
I0HjY6VlSjdhrFQHFVC4wZ2v7UiE5Vutsbkosu8b5Yp6zI3f+FL2y5DG5p0B1O/n
DkGrx9aqkxAKrwd09Qw/9aa3rV3iyEjtqDndyWJanTGKPmYj4c6FUN/GxMm0qRNW
ww5+Tf4bRfvUOte09J34aBPpifey8sAnRXxRgSlvoSuMFP3pO4SwIDD6YY5rhCxr
EsfewzcLVw82YmpN3FYjccaLMGwZJw9zAJdwkzCYdxXtmBxwFszDdPYS5Pvm5Ara
lfzWMN7q2T7ptGp5exJJoUgdQgi/Qf8A9jF1iSurX7Gi8Zne+nSxuY9bio7/r2iG
twjo6rEiQBO719/GvRQXyksA8YeNqvuikH4gWCCZmDakpWmjWlv/nLrvjDbOcU2S
jXYhkxg594uTwcvZmBdPcp1kXm+RU8B/rd7xohhYrWGpl5O7GJ7nYR63oZPiCXY3
VjkbU4CrkZPfLx2+uBkgrvNq3ImIkqZJLnmKGAwgTGdxJOi4SrHjCR4Kdg2I8ECz
uzGW/o3K8FoNrNmebjeE4TOufgZTUoeky3FGNpnGC7yCX4WpeKJHcIVoWIOqYtMU
EBBc+BbbZCB684VCh4hbL7ZWFvu/UBgcc7PUR2mHGZUmWHVQEYSASXF9Qdgbt0R6
HsbJAO3PPVhfw6I5uhzuQVduI+tm9e0aXfdF3+et0LrTsZFsmBjjUlq1Wy+uH5uX
wSWwIws9LxOE/vu/lNoYjnb7Ln6wMt9vtAE4M18viZm9y1CFxOUK+/OUtY0iNB7C
TkQgR6LZypj5gxExfpKUp8D9s2o5/1mY0atQjfAo69EQeF4KdCRhvPx+7rlYVwPE
xA8zgnZYPV2p0wT50ZufW5wKpm9Y9VOe47f49cD7g20wMO+gkhgVdF2nUhtFiOBr
HC2Z0piJBi3E2z09GwsJKCJXxUFYPM5Oxdg+9cRoxTABGhjL7IoiHMxIU/IUB7O8
mIMlatNdJHIhbJDaMKvH4rOby5xSuGMBhvlzy1qg6uWZET534PGw0bBD2Zq/APuJ
BLLoZUtWZUcK71blLG2ZiR5y5hLjxdYuvp9Z5MN9Cg1MjZdLu7JFg65kjAFpOFSR
nWLKTlY/99jj9jyg0TwGUnyo7QY7nr/QHC2PmIBNPrzou6ZgM5BNqvrKSjQxy45V
Dkh9ZArIpG8d4RZgGGcFo7HqK5jLR9HD7j7lNcXGocXP97wLWDVa0b6+kdLxmrm5
6bt5SOT93hPh/hfzVr4laENkCDXnXhoqkVoGga91QCw4nu97U7ABIijKkd6pxXfN
+xF87FknFEcv0JGVDHtVqEAet1bnn1SwgWXzHkZAlZAMt3VyVda5kLsQ4X+Sbmb9
G1OKQJXwkfgvYsyZTRIk8AF1MaiPP0mn20zuKBJmkdA9ir3mmN6LedcF1gIRvV1a
2cc5EnMzXYLyJyjiZfzFs/Wq9Vq64O4H/yGvNGXezYKIHFV29GSPLhhplCUbDuwj
kovTpPX2rwJrS0fctx/dXLR3al52j/wXtJ+70Od0s+N4lmBXAxDOY5TCTan6klot
5V9BsTFmwd70Nl40cWi7XaqmNXVBrghv4YIW0ZOAqtz9TIsuJ1oDwWBlFp7iahZB
qrkpiKCjBsO8KdhOYR5yVcqQZzSz/nJpVIUNJu7xGVgt/+bs8kmxWLcTX7HhwFND
9xVP0PT+FfBf1Wr2iSeQDvlKUdFQ11k4GEy5kla6EGA0rKGf8UxIUOJ98tY3+Wr6
wd42vEgQBE8/nwTtSO2+Ef7sODoW+gsc4Hvj4gsfG9x7Nbt6HGP2FY48x5hgps2I
zK4o8yqbQMcIdFzWXlxh8v5lJqn9JEFdqJqzvWhB3ngrOj8nYz6DMA/W5Rg1bR/8
SQkbtKFuSca/bTY/9iX5e7jpgR6FWWeX7Q1vn1onQ6lRf8rC28pWN6ybs4B+9d26
/FB2qcGB9MpGadcYKukNznwlw6iH+sCS5aylT2g0ZZ/enyr/DRcDFM9SQ9DnP66K
g9D7KW6Q253zg/BJfl/Zv0cXFJBAGOQSaHytcR7DvbYgq8oDyt7tD6gkyQANPTJI
UjfhMK+joOEZiEt2IRd3eqMSxiNpVNgdoJqZnWA2qRlB3r4bzLleUx6R/cHP4REW
DkoQLZwIT3dvITyvMJFp8G11ftht9wFyzvF5Wx5pLhW+nfnBnSklT3iioaerUAwh
WLv/3FMLvmDCChd8WQK2ngD/aBOkuFcwPThksE0dJw/0SeUqsgrIkd/3TPl2HR8j
0x7fYRonuynmkYUEHWu7+sk8seqE38pN4HwOBnc+QpuoT9ebaYqI5p2YhTCoNnLX
592M9alvN/yd6w3upRRj8WSdMUOQSnUMHkJKTH2d40z/wfwykB9zyHP+QaDdyUPJ
3erNPSH5ppGgE+rZZ3CbCbRz2vHuEztw4KgahzQpOkuqsTmc5ZvQLJ5hqjfX0MYQ
96n+DKaxCHT11+buaUwlT697/8yTTk+zijzHeKgs0qNqIexMYknifiiiqvxACfCV
k3fmbkhxFS+A3ck4j9S2LP+ZH9cxGM8MESRdtdXWKX73IeRfqbsYw8lzOIREs+7Q
7M6QZCUpV/WkEOMxVBfJ05MMWn8KFWwxLw7/EWlcF7HMUT3SZenU8cnz71hPQn/+
Sl7GXHzmD+USqnRJpg4cdeGRp8EMVh+udv9Dli5Db+sZjPXGpVEZk7n5LKlPNrdX
4HMvwwMQPbuD7q7y3d1O8LC6c5Bnu6u2oSIZvDjmlROZNCxs0zJwXOVoiqQMSdRC
3W5HvbUcbqGcd5gN3A284azqbWbK98M1edH0wFtFB6PIUCWqOOexKnU+AxzRNBY7
GB9vkiuJ+jrwGbdXILsjts0XRhTlnM7f5yyGcw6OCXYTiN5kQ6XOHKprbVdgCR98
WaZRCeXpwSRA1aWPeOkmlaLMRjTbtKW5BJ+8FZzSwVB1vOWOqLR27mD6AYCDHUeh
F2vTXX2Wbd7zueFSXv6vmeC8xjk1X54gVNecdifZ5PKkKI/v00G17EkOHHPCWqIt
BHxubbQtH5irpHACTrzKNC0OuNz7lg/aqUu52ESTkgBspKNI/WmJYU3CNPEPCEpG
f2mTvyiR9dQdNTkki23ip5RtmPwVel4uPE9QWVVuGSgBXYlXDYE7pm0r4ai8ltTs
blbTbvv5oEiZbrBiY9rWI+TtTm52BijKlRSevs+C9eekFRx4/xte2mxeY9IZYNDE
zK4nVNws2Lx2WL3CgU4RKh8dNPOvhxPUH0HCa5/xlJa/JECKOf1RcTRZh0nZq0QN
1uAGwplfT+DA0DCihhPIFBXwSCO7SVM0fLBe3bbTdi6TCZ4YXzxxnEjGO/U7xczj
iQ6jtrpT7ysZj7ZsJ5lq/i6Nic53/uWSTpB+LeCdhufx31YQ7xbkiBLMXQcbjwBh
JVgIvNsMyHt3YsULvkcOxdCl9B1U+Xf+cpJQKHG+tgk2t7Mukat2kBkEzvIjrfwv
zUKvUMZXeVLz8wTe1MMqSUjvYGeGxTF3EBYUdGfNTIsJYt6MuDT3FbDjjKyUi0vY
f4kIp/4wuv5TNt3tTLwVvNJ0FIvjvG6RxujNg0Q7B67MqQPbz2hbbOpLLVJweM/i
RmTijdiXJFrnRMP7sF/ps3YN8eXQJuO8Wi8Bey86yk3GICSbU1O0WdYtFN5cK8Cz
bxHy/YsTHWBLGl0j2p2F1/AxlnhfBaA8VgDGvLobkhPyF45TbeiSe86tqiJhBZ0h
b33uAZXnEeQZLjxI5WmqhWdkuk61HAOc60PVfHKoYYvQsNf6LDl881g9SuIBgnJl
YwG2DGeINpzqM+yTgRnDaKG906+j4K/IcMoYp14Di80JEbjYjCIhA4HESrlsseVt
GjeRE9WOpDUMxWatw7Va4zD+bN1jVcfs1joQclY3GunZ5DXLbaTDOwtw8yqYmXeB
ECnEy9pRkaq9dMcyhGbhlkH9sCuSBlQlbTp0GXQxk8Bm1AjMVZF7gf6A2oNx7fPc
EZGDcF4XVCwSFQX4cymhQD02nrd73iY6NKZlBHcIHTG1S4Ce5dl9fvtK5zjjaOH0
0/z2LOFvR0u60wMGM0SLkGEJCl/zdsI3S5iHwSA1iklgBHSJa1Q4phlBf1mVksC0
ZvcME++I9MhT1TVNxGvyHutdPb6+QV7k2Uf+f9DhKPtPcx7t6VEnM6Lu6n/9Ib39
gMVT4OjnZa4ubAL2FrNWK3hkqqvJs6kTvO5amONfkFWrk0/XzCrkePLWP0OI9TFX
O2YSw/9UsbfEo7eyoYWYb2r7rUB6tCYOGjD8b0SshhLY3PwEnOkm8Co1XXKBXtpW
Ru91YSGxED8xG02dfrjXr9cFnA8dFqkpeYKbmkrpLyN8Tqw3C2hCXE90i9ZZ1NVm
/ymXk5/TYvdK8jUAWl0xSnkzCm4155enSn/WJi0QeLmgl4U/OmimRclz2oXSd22A
v42Zfj11B9hyjemuRyMusaUk7J82Xeqpotwp9cnBJn/8NOG4m3NkZ9hFt0QQUiPn
aR1KydQ8UOVVCgk3YVnSCCLpLQkuSW4YS6HpelBiMLK1il56mljgnZg2vvValL9b
CwxTzIqyOUd9T6dbvQHbWURRVshhNLblBxfkKHBc/qtaQDf4P8PM34CTqkNU00sc
a+4sjPYhrc0johkbmFgnNHjGlrJg89MbHhDVZD3qRSEoR9BoKD6hP8HYI2af5YL2
19H1qvrR4stQAT8WhEYRtQJS1HKT/6COxvu4YgOE+bA5EhT8770tS9tWpBwVz7mN
OhLkDf8eoM/n6aEEMgQkwUBUdkIshWV//LdECpqU/FLVIUvFN8f9vVbX1RuFKQyD
hFerAXIH9/xiBat/r8FEzKTiZ8aCm8g0T4tbVDaJ3HASPtcwWs6yGauWHbSzjywn
FRfyJHibyDtdAdHP3eXM48jlQAF5BgxW1j6tAHaKz5tEDuTZuEBag+lhtyo1trHN
9BYDO5EHPiEVlS1WLoR2btSouggH6oqjXX0QLJLuEYV/vCBZa1gc2OU7ZGqjaQcw
Q7l0FcNraPT8lCyueMACsXggr+uuSSU6peHkJJpF6TmrkSIRUeyPWa7rVZ53xLV6
YRUtxezi3s8slmDcBZJway8or3EyrsDsrCVN/TtTsWS7I8oPwTDEaFUb50Csyrfw
O9VhVnxDe7IWvFIp9QZGjX+rMVG6KOg9Su7vNqgd/ze/pfszQX0BQloUTGqazO3y
Mtwkl2Ok3k3BmSPqlgedRI/Mxq8cdPjkeNtL6hG94imtPfkK0WUjbgzdCKBf+MZX
DiPeJ2PsGZbDxroMu1jGBzBhuV8lC6p5W139nbJ4ben9B0Z2ZLkGfsMxgvyu8FYZ
2e4O46LO598igjjZjLzZ72TCpiSJfF63It8lHWBr/RipGHDhm/5z8Yo9odszEzrJ
XLezsCv6h+hxALJlG5EDtVjFJOiCCDvD7ngCnoI741wlY6Ug2clNLbT4TjZG+W3N
oQ2spKFpUgJJ8Ad371p2N9Er3qYSpaGM2/9rUBGoAPdDugI/zcEYMhYu5yZo0tHp
DDdwy+Sk76AcCdHD6b51Zm22u+bY8QGNUT9fswBOh+p/1riQr1+vGbfOcj5Tz2ku
fdgFp/hAr45qe0g/4Sj2myHlGJQdXakxvbxCCmBMVgtw4r+N1uvvh3aMJ3FdcX7s
nFadUalZXMrYIS5dsvp7DH+ERSej4M3FdH135ZEKEC/R3oYMZiYvP+Bf4JroFV0o
sLmrpF4MmDuKXbjgoECb/qJD4qCauM4WpmARQqZ5A7cVz2QLF0pMH9K64uqNG5cw
0/jvRSNkg8aC3+NpEgJmPFtPMjoRE5GyIRglYu3l+JaF6jrv8y57XxTurv08yUjE
sHSWFxEvuvpzcFSeDNcQSVl98CQBMsF4Qdbxpe9k0GaXqPdblMS/8oxYV/mydLSC
vnPF0KrT7DagV+mMUlrJl4JXTq8EyLm8PuII9obfC1DC0aVsimoHQnOQJX6fivEh
ByE+MLq/KQrGnp2GaYbIF1d4LlrzaT5VH3ttTMB3M3iA5BpELPea9Rqzhpt4/3aa
2O956BlN63zPwWkeJWuMuAwBW8MjNHqWB14lke2iQgkzbUp2sJvXOb3KIkGQZ9ZR
mhMCDR1RUpLqlYSj+51YJo2EnHE/T4erqRmjz1jpHaW3OTScnqgMGtAkjEeD/zeN
1vTk0VPbBS10HK4EHU+VqNY0ocaxhrfbOOqKZs2QeSj5ICvreKye94DeMRqbh/HZ
vEOOGBqx3f5SCXgW2JNuhB0rzUuFgGgae5mh9TszAE5/+lOOCoam8gZ8wFce2R97
cx0CBgi6vkF/VcTdd1dy0cj0Acn5deL2YHVoc8z9uIVPK1xx2DD3pWyufpIwxQCY
uGag+6eR9tc6dIeVbSANb77v2Hkjy5UCcpqYTaWJr2pdj70AhF3wBjkTzp2zmpiD
VEz03p6hJG+F67N+c8WIRwpdv7+1qZ2WJ3CFkjHbmVPUesLjYJXLTnxM8f4duWZS
R+7W9DDpAn0b+/iT6pYlgn33k2ctzMzaLbk8CaCt3KLvR9pAN3RWWTazrYKfO11W
8n0dk5KQlgpneXEZncRw6EPi7YfsskeiMl2chzkFZ6dl4/dE6IlGCr8OnX1pAGj2
QgsfDlAs5Ac7sF7PLELxTYxKOU4bQA1vypEdHPdmEOKYonApfm0drGYkr5M6tWIl
Cie4oPqHgfaC8Iyz+80jqzb6TYV5Ek8WcD5EhAye9M3pHfOzUzMnm4t07azY3QGQ
3VIWEit9AHpo/E8LOMh4jkWbch3+IsgZEH/IXEnr02ngb9sL9O5xxOgxKuHzF36o
RsKu4VydHG36fgnLL4aSeQ9dJ+cBMMqHfve7BPWHAIcaIOUHZo4IUCGkmEmGO5Ec
6XS2AFJmal3gYdttWx3UZbmhhSV6gZdJ1u/aIznf7vZXF+S3N48ANpSNJynFOWG2
lwRhxMvJDYP5FyhVLcyLT/oSXaQgqUFAUkLjP4rmsEFoXAZiraYJRivZLPdfIyiK
7S9PkMdyDC5rXYxTpjfF8zKYmjSWtcT9mkbk/nicrvnDwuawBONyvAwL5HUm3Ww5
Sj1Tn4t4hD+hKZeD7R6qeBtMmCAxRKuTdjZEUQAjZNhCK3tB3GUasCu9aUuLGnhq
Ei6hAMyBcN94rRF+taMGaxLvWSNt3vaM7q2kjJ1yjKPH8fpTKTqBnETwDW+PmEZf
jTkARwdjjML96y4Au6dKB1eJZfx4k6jIqaTUuEKlk+2yuLytZiOhfojBCGxQnA0e
gnIp62eA1j1IDDpXkOfNnu4vl61iJQDG7u53kiZXuIPpzQ8lh456h8C8p2mzuH0o
P9fCqDHfCrcq7KdPicfmEgsG5j/QB8a+Uwx1zwe6gHijUT8sU2Q1GucIVZHfPU3V
gnH8qFR8JgLy80sB0idTNaQKstFRmQ9PdvTBIXZOgxxcFrgL1sNMedqF5ki/VRNC
z/EwLhKnVrX89CdhOA4gzNjAMhubamMXE/+YUaJr7dXft8W7tpetvx/X2a1Tk4HL
yqdO8D34HxZtvcX+ZqpLKW9qtiEVeQmCqZcjCii2EqgZ/u0FSW5+rlApbIbJoBoL
m+nmWWlvcnyNwaV2+2LRtgVNP9PkEHyY2JrSpXU7hGNzbFs1F42X/r/DGPS3Xbgc
0K6EWBbwmU0ZBhJVXbaCNxjgVaTAPVefa5Fo52NyEK7qLV1/MWUha5tOynPw2Mj2
e9tnolusXFf38cMZjSOX42ukjvNHASRzIa3FQwPY718+QET6Mig0NV16X6S43xBy
qiooxhEQB9JxMyPgLF4WREplqEQY/cPCBKaZHeHQyBEWAPAdSIXP90swnLYQzPz2
zJ5zabyWlQdmys3hfWTY60P1N+QIGPJjJQmIQhJh+Furd3cUDxdVpbs3gOEEftib
pCppxlK1ebyiRy/n+JOy0tN1y08UQS6dutpT49ypBfLea1GPSpDLFF9liX3DMTG8
sTyXSdl8CieVDlm59wro+A6TWGHpkteGNLDbXBOtxL6nY/UW0s2on+3ffynDSYtf
XrnNss+qJiedPriF7vadPU7CNeH1ihq/BOd3mSvUKpFjNiJSwxJ+kJcRCC/2CiVV
ft8hT5Q+oSbfNMYDMuoECnuQud2u6TWM7LtwBvEl4SxxdVN0jAvkjM8jAmRFDna6
SEN8k+zO8+ZdKquHgoGeYf98UMXfPIQrq5WI0UHFtX/oVOaVZ2JPjly3BGGHN5jV
2OydA7dqhtpazxVaVTCXexpRHrKWkMqH0ni2bZX1xE5Z/iwWfAIy103pOwjBy5hj
nwt1wd2+t3VZVA3UmJYpZL9UThU6gSzwmE2GL0d498YhsyhptOKXYypqoQWe9IJX
AfjR9Fbl+tSD7Zup/9/FwTKxY/50uFQmdz5OIaM27syZlU7/Se+D/3/j+0X5YGsU
Rv1ka5BL/zpHi5HLkbNlH5LxyQhw8KuFoushfeNyDvRNOmvCi+YjoBVfGX23FTuA
nCAwCHEbXOTf1kMNyt9a/unt7CT5LObTQoHcbsuQERbajerKF0HAma3QIiNxNJq+
qRcEPjwBfwDWWQHmXCLHTgZbu1ir16rUwGPbKUS4B2hlXnd71CjgTriRutVO27JA
XMJ4+nI5++nNBN/25y/ETh3+TwBMpvJN3+miIg3nRY24jm+x8H01CmoqPsR3/A89
EKY5fc1UKDzKyPfpdUTqFC1sgDC/0Hrf9IayjNPR2I5tNyzIwZRKfr7LqJuTxMcY
va0e8r9zpoogvt0qAArgmj1qGA7xr1tSVQTVRrafhvCnoQF/SbJucrpJo6nYaSY5
MtB391ZqS7CxMDgWp0dcAWqRMwCGy3tCcXDnvR4buYkRwKa+pNjoeW1uUouB7wJ+
dhkQXHePjro7BzUshKHKzuQQRr5Hxiv6jP+A/NweE99LcEEfsN9u8kBNlZZWVkFg
gNzOgQjoZrjmZbXr2aHk/sDABLCgC2v4g1iNRNooQ25Y5bvWZQXKB1Rja88nldzE
56ae+Ew0Uu+pe9cAyMwRMtjLAGSwRO9nSRR9WPhJG93pqueK24k2NIyf8VgUsJ4c
Qy2eUF/mGrExcpn0TW4WHAzkcocozGGl6bycu3Ks2zwtd3NTLW2SwBXkjVl2OwpE
X8gYzd48/BcSOmK9hI5dxLwhP/ZV+NNR6qVCUNq6DpWcPleYK/sAFvXe1qvjJT1e
ljuSC3LiHf3y11xdqePdnjKRwYdee6FaQ1GEbvoG1iu72vCqnfz6RPaFT7oAnLjR
jT2Yz+9xbo7P5xMKZE72NUlIhqjIoRoK7T/7Aiu/M72gyosObvljrOAq5Jzh8dMh
SPnlssJX22pXW5ZuuuYcenCeRkSkmqV98Xb3f9kPrlKIOov0+TMhL3aJS/BqUFKL
26EWgXsGbJ6Yd0Rm7NL8sK6oekoNCLX1IRFEtluqUoPOC3/z5a7va60uRRGzduWW
LTTvmXz7xvEX6tL4OFzg77YsGwxQPtrD8Hg73QV773VGRLiDdwYIMOYPaaF1vPVg
b6U9n1xcUTnCyCzilGBQJBWk1wflOkrBAtbzgJCfpz+q4ekmgAcGPOBv8w4R4GIV
hGEKV75wpNJGJdayaGNbFzbuK8j75tvX1uW2XmRSpgWo5nfU64+0il+qkrHJ7EJ2
PwbWhkbCS2XNioz/Gh38LWah3Fkd8+Cy4i9s6WR6XHzFqZZiccXziSBz0MZpf2+R
2B+QaduKxkySG5ZnFPTGLcqJnVLUz/7fdCUohqXdLdpX4QoDGtex99RW4+JUUJqb
tjch6eonLiW97OKChMq7bDcsLvnvpcUW1c+K+h9e/FJBtkU6A9jxjiSVTNkWgDef
CoBktHT/E7varac7Griytwo1PgulMofdZ9dgP1iOcDDi3VVCgbBdaOf3I9OT+YWB
UT0tYBOTiXQ1Qeby7jAwsaMGlQJJ7QfMvqifPgEop5Xa8GEjj/wB1zx0O8sC9Gae
7VELE3JIrgcIjhJr0n1El6yRKxJWB7JI/qV9bWza4zM8B6JayU6EVCXcFiucCyGT
DCFCVt7Q5vsxiEWdehtFu5coKkt6QVhwCI//2Ne1wRE2+z1JeCkEp8HrPGuvwqm1
an9KeHMyq8M3P4eoZEztCGTgppJ+FkqWhnE04Xq2WZkxOZQxfd/b6dJY+N2GnPrG
7loXddZLI8IPl13MEv2W9RneRyYR48hfdtiysUEwBuwL9kRarFWAsA35l/RPyZHF
grbcGW8PcJNYNOgPfb40GVY6OJrGFO9Lovff9vj2b5MxlaQaQtAdnSoS4cWNRgvQ
dVXrSXK9ojha40mIfs9bJSgiGPmgNGq+VrRWJZo+VgQl8DTTlLz7TiD0Nu11QAi5
rpzjGdbEz5ajCE1WfVkh1KKonjcz6BOjTGQ4v8SNsuXIVm/fSBYJDT6cMgWAbg7z
GUZd2HZd48YLEkGzgPUJsHJ0IN68gUqNM4GIXGuM4RTvPbSJS5jCKYk3BwptCLjN
yfMIgan0s9reVs1ri/jGmy385BJiG65HPwnqFvuE3t8o/kdgfx8/kHbs/XMvgQ5P
OIj0f72/EJPJJYLry3fdA+JUgbJW8VocqhFITzgeuX2osP+hVI0PSmfKK7mY9Iaa
CjGPd9BK1IAN6dz4F4inaJ+Vpdy1owyyHNeHspfKHaNiHbNvIYJ1SJ0di4KgNwFx
2NkpywJX/c4qSzbNwYpAqYo8t/MZhwbT27F3OMUuqLcNCOTZ/zaM5KHlaGnMT/v5
vAAs+KFNhp1/8rWBA17LTM3t8Hpy0LOm09bB4x0fquL4MDHY4rPuIBpw9FT0rPwY
t0P+pEkcOXxF0lo0OPnbXcYAmUbfcRVyp7gLilJZyPxp8JWn2/wK8NQP1MvKrdqn
ZGoQqTuCkbuBPCLBbRbLmfUohit0lbmPKpFzND+VE2FExx/d/yhHm2QZ5qLgXC9R
nxTR/JjOINKj57HRqBrG7LEpTYXeWOnWM/hK7ZyDb1dcc03mah7NdlAPB+oVUCqJ
UXln56luembtBRB9o/s0BVZtNx8nXTOJdKubmr/4oLSizjxpZRNuHWJmI46dzAvy
TN2utiz8pft9F1CFNy+CvKe8kRlY/0vHdoH/peB4eES2D4/lWp9tLR7NBdAjON0Z
+3y9NI9BlJQKYVtDkozCvJDEPquVN4DHxs3HDNOK62KzRRymt6ZRnObQ5vBAXVhI
vtA/X2KeKk8D26lGCHFtXgD6EJVrRWifeuzTswY7ZzGzjoWP5zrT0zVem6SkJ4Uv
vaiaAnWrmV0wY4M6fGT4NOQq2qACnEuO7Rr5+W2UV/XGzwEzv7sRW7/O+Mgwe1ts
cO5UfE7fCTFURC9/UgYB8GAnaWdN0o16NODMsqlNrrW85Wg/O1KY8pEXJCTfYhlL
SnQ0CMY4ujj/g2MVNN+50oy8mu7LwqTfMIomn8dZNg5nAEaHZHTqmcoHzDmin8CO
BCRTA/Knzib/hpZhL015G5/QTvCaBJgJCTdjH5TMVW1epygQgI22nWB0FsTxbuO7
F3hvX9WqoG6ANdSfRSO1ZrEZBdQxWrJ4eWQhDSs/MVn7yBhCDbLJKfJ8B8rQUMyN
rMTr1Baog3GZyFoxLGr0Lwo4RDN92vfc71oQc0g6an6D9V0aUq4nI40AMEv3EAPD
taofUltKPdZNpfvLjMz2i6G4qbMgca3W1vGl9X7ZtVp1d2tCl3sgf/5/B49MjQqN
9F4ga0iBksp/JkXywsL5ZoIq9T1n2XioA67JHecm1kROlPqHeJxz1XQc5AeZkxWt
wxa+uyzL3sMID8GszlcVZp5Oy4dQjKvJ4lU1VGYzigqAlWW0u+XZaG7U3Yy53xgQ
n+o8OAXQKFCgeZ/EMTLbuU//hNcFH4bw7QCfytiRLgnY//tgEZLo88cvugX6LkSl
+XnmtVCAD52FDhlr1wR/2e31O41o9IxQEfcdJzKl1Ljw1DFJTx8OJ1+QqvdwZdYq
96zlpcBpQTbqzOaEsLyR1L/g/5qSe3XunM2t/+o/joZzcsOD7e/X7w+7mdQpVW8I
SUa3mdi2X94XF40Cyy2lqvqsq3o+xjoQr2+NPDbcrTudAHdJqiOLuCnSOsnho+mN
8dNaCm8rbi5N78rh0qBG6GCFPJkdLqdVNcBtWki5OfJY1jciqa8pUdJLI6Lc8MhX
GI5egUD1QBbQpL7uSO9uK3lvt8J8y9jVm/pUKkWMVtrWEBtA4aCSzc5COO6ckkM/
3B7WErobMsDGifVm3Ow2lDtmQzirWJfZ7PFuuusZm8XnwI+FYu6L2njlffeSO3s2
KoFjHpV6mSfwYhzbZYtJk8xHx+BrZahWzWQ4PLSAZKclfV46M4fRN61jeMFi1pOH
Ha+xUGo67htgEVtS2u9ip0aHFAGK3VU+oO0YygAcQBnA0gs8VF60uDKfI6LlBBSr
ZC5pwpYpUlQNqysvNqHjfcQrUzt5RNBcvHAJe3KEw076+wSTSYpF0PxMofFHaA+m
PfsDuNZJpg4rzS2kYPpMpf3RqGPgvN23C3+uLsDNwFMuEopzGD3e0yY2BH0N4Mey
xEtTP1RyHglK5Uvu1ai2NUa6MrEKhbDpiMu7raJKGf9xl75bxESHZh/3kIZYZ177
smLCVQwnq0ybNuaqyNbbVc0J2PGzJQn1i2/d4lEYy5wgrbkvufeOg7+Ay4Xxi05D
Hu8DLOvDFeRihM88W6UJDHO9xd/nYCR/Bfg0eNDOd1EoaFG0IhQyIGqp3fqFnyAQ
BCXchanwua/d4NFD8iBBxzM+gh+hKhFysA8fFVNcjv4yZKOkhXI+lyeR//Go6IZf
KKY0im10OuTYU7bWMV403e91q5DQs15k67xx8EysjLOgzoetOdjdO4E+6RH58FHY
QM+pLvAMXQuPM+B359fdt0dAaa4YvQWsxbps5Fc8VusvTWHwbsmASjj2SwYnfJ7O
MaWptdGmkHOtuyqbdKS+LTMs3+hfrNTL7NOcivtsKJlcsNLmR03l0GvgQ3BvulGU
8aGGCTKLfG3Utjy9JdUOc57mn+xgvOrqyRPCRM680MIN8rk8XRzDoq8dwBw+Cy1W
1v1MHfVoaBAUrCemG0qn0KLOAzU+kM2ioIjN8Z0vYpLxepQ9d7wgCJoDpwCfw2FY
rQblRilaP/TS1LNEP/E5Ogyikj5eCyr34Ee/lpDhbp4d6D7/ZGWEAZ+yrFEcbd/U
pRae/vdz/3UOpZnOs0LNJ3Q5KGx1VLfC/iZXBtNZfFmLepLowi1cFOBbfoOUJrvI
XgyXfDpWvAyit5vbTEezjBYQ+ZAyrnRRD518M195OPWoX4uJX/yxrBo7zvfAIK9y
FvOgsVYmPTAPO+EQXlQq0Y561tpUoJiuad7o5GPd2YJZJnZxIPAV96T4Gz0+Tu79
tltgHenBL4JUNhVD2XAfimouDYagxpkJIN9rhwLp52yF+I1YHSTeMgKIgLzrp82t
y9A9yi/NUuj9562+DgXWyMypocOObOUIWZiPRgAglBhN8NLjJSSzsXjkBbMt3tM5
Tn3wBILMBVGtCMWgilIm2ngTqu1pANaeD4CxQmI8tQXNoI3zyLbo+r2CU3odIzyF
hBBcMSqisL2w/ZffbxRHW82EkcyKc3v/aTFbAWOK8rszB28bq15NLRXXnuFjNmJk
W6Xm/tkSGTM4YymD1S4XNbzwNjGnFzU8kvnOzN0AFPWbPMO9Mnax4Su1V3LsOr4P
mnlkgZ26nrnPQ0s/FfbtpIf/G7NzZgGJzoAjAP570PC5iq8iBiFfPGKqk488J2kl
tgzLxJc3xZNHX1sMZFXF9AG+OE1hqYWfNhBdSxhYUd/+RAWqxJTl7zs1SqaYvkls
VBQMbiScSOd0XD4DN8iffBjUz1L9RbPmeWFpRDww0Fii5vLpI9zLyPPr5p+y5lFF
JZSu5Y9zP2FrLh5zRKY8E6Z/I+tIl6r1d1fhLHtNBOfyMjUwYY6VLSpmQLm7pQBo
loO9oG3LOwkVx7pnKepbsbJuGSxRZQMkop0F/iEF/+wmG0OSG/02uAPeivQoVxxQ
68N4DWAwpGuA31+6wWisHWd5CHLhxL+Elhn0a2BviZXbMThbDwE3LaClLgP8Edag
qWFoWa1c1IHbWqJkMw8hCW5ppW6qpV4wFxKO/br3ZOftfhE/QbgapwLvuYmJOgJZ
Ow8lfkSHsEmGm7VnGk7mKntH6HTYVmTLQiZd1YHEVinNKTWAxRy/70vo88Jfw83w
kYq5B57Iy5yP77QiRoEcxbDn73pmFtlOtDKCxbsxU8FLieOFj1vUwHeftyAPNwD1
F98gKXq3YlePNQSikgMkdKmevncikNoxHL+oO2azH369G13vdzWLckHgLmqYvWF6
4VDIEA1rlfLeNpa45SL2k15bDhKM/+7MYyUWllnaDtrCQjimvG2sLltbXkdtd3t8
F4BlorwDPypLQ7Z8YcLy4q5ue8hUoBdH7lo8/7BJRc1zUAlRS4RvPE//+Q5nRFxk
bPzLXufHtCzYllJL/CluP4lBLXQysTyAEARjVfEu1mjKb5zXcgJAUowLNlCkOja+
2yFZY/hOaKQOLHdN//lo+XIz2AGyaXOzHaJKfYAvCQ7zDxTgsrQL9Ei3x13NSK4L
j8GVt4qe5pVnyNjFdL4giStIdUYCWY9aGhWPXfzNIb0CcX8U345BsXKgg0eSk5QH
qqUFlwrns4HfLwfDuiF48o3wus6x892SorM+PDKlWq/fbD6Ol1NZFnHT2vfjEJfX
ZJN2BQ5cB/vQAwPr69HxIyymmjHpSm4BuFxbFSoGqBvGKnB/5xRXypIitJJ1CKyH
w64HrUerI4Pgkzjb1+15FSdzmKM1RRyaPlgem9OdKYDIuMuPF+L6t1qU8KXTn4F2
vNPSiwy78Vfddey4GZIMnqGEVNcH+50kFkq2grggn1oWR4vfMJvvQuWnaCs44+Uv
R7sks1sC/zbTgYTJUz1DBQqh1JNK+3cf19Kw2tnbT/tQoy/bLD3gP3M4fJmozYo/
QcsVuUzAzu0GP95+NZ+hbyWABEx/xvqpomDpXHFSXdtNrKj1iTsEGBrBbO9FRJ1w
hBcSRNH8Y5GPZDLgX3Ovn0PJLebqIikhRTN7O5sF7KQrgAQuzNjWfm9balxUFboZ
2ybMgC8R1FIXYzCa2POdeWCo4WjmGgMt02Fi1yHZiFZYPso7iDfjq8SjEq7Yl1BC
Gkwul7ARtgWHGoAVgpotmzbGSlp5VUszDjf1I+J4izj5wR10znVelptzbJ+aHnJW
FuEnRHRJ8b5z0OEyWCYMLq47an63ZAomjv3sxjr5i2MNBiAOuS74Rmwi4syM2HIE
uX8vI5eEIBOA7R8TCEtBF1bZ81OJcYDtOPhDZCITCBgyp228oxhWQZbyNLdA3RI6
eag6VwjQqPDN5FOMBL3R/js7gqSDiTAwqmWZOT3qP5BqB7e7nOlsmEqP0w6LsfNk
58Somi9Xcs0C6RkFChclV2trcweiR3UbxEn6G+MMr+rNcmrxjPTeGIMUToZGgfC3
4U52PKl4qZuuWOljstHK35E1rCcPh0FBt3CliZy65CUGZAWbU8gUGj9Dnnnx6TUw
g3VdBBDbvrsk0JuhU4yiFH48vNPp0h8rcNU6JnwrNLxyA6AMUiqlhkZyNLLa05uf
PocHju2POq5BQvTJrhzvzwmb8BKAuo+iQH7m0g98RaQPs0L9UO6c3JVy5+FRCYR6
E51/48pgDT3EphTs53iov22hsE9NAU6infJ9bfAW7GM3YwgOeF5pe1dPh43hizHf
NINFX2GCxzwW8nLci5aEKOv+OSzrKcG0CeFSLVWHHXOIGryyJ8GegENKdU3skfVW
kD86ju6Bcq9Ysu7W5npNTT9YYhW4rNsyNvJ5IH9xRcBtKQ14RgFgls49p8lMo1BQ
P1rXFSrsyGzxHiUtjjNGOLVV7EhRJcic8shtt+y09NGkthGop2yN45MlBAsUrG7F
2sSRGtl5mpOoXcji3aGw4JT2V2GVTR9WtwInfOaQ2MrqM4Q+DqlqeW3kzvlRIrnc
WHF9KKr35iXKu1JyXQhJlTCySO4+MNjjZLJJfXxhfipr00xzhTS//gnAeCXL09qx
IwVNOFm/B/orE5Pe4/m+j6e/Zm8v5/Rzl1+UpJG1eDEmevuCGeoj03e+UsB4VdUY
x4wzkKlZ3EhlsZ3r9twrCopbudMiJuZ0YFRzaGmSFrTjhAntQZpAfUAZlExSqmJu
zEHXA0sY2WnSBHhy3oMbcQ7NRv8V+QDUBhGYlz+s5G4ej4C8eaRvJ1LqGLNlhyB3
pSLMSq7DmgE973xlkcPpmtfpEfDX6Znjyx56HsHiMa9ETQHMLc1HxzqVfFqwISkp
aI/J3fYjPNo/n1Ff7tfQDbRyml/UY7X2oXoGY/BNh1V1FPCXbSMCERdkOcJ8d1Gz
YTSBYqtS/7ZFkuaMW+PcqBYSCf3mqhtvXp8Nq2vjaX2hNI6IpCixb4GAc3aTFa2T
IRHbzwWH58esqr8kZygBtXsaFO2sneHo9jIhDNPwxQqkdDfaGnYBEAKaDpB0H0OZ
DbBfziYVurUvL9FxdBV1haoBdWPIpfyXxJGXWTFod8uuZ7kMi/MiGJHuwjzY6UPd
mekT5+t2hSwUGxH8KvI9+fImvvuY33wEvxYdPvFdNj5n8vvQWvO2Ftpvnbqfekiz
brx07DXL0x/jBhAdrgVCkv2L2rPw0SBn+JB6uakXe6s7dmkb4j7vJV4j5/5Yn9qj
Ywi1On9wivV+yIn+8NQw6uBr2rCNTn9/bHJsG/cJbKbjrpX07DWAqK+68ZNPaAl1
+ASN+vLJlrXmYJe2dypzRgb5eKx57r0OtrcjDbm/u5cOx1JfJqCwffkFGRoqgDY9
ejuJiAfcp/xRVjg61fCgalGidU6JFu66f+nnHeQacWng+71aAw368S3t0vPkGyQH
NScd0d6mBktJcYkAazJGM9Lnh4qi7D5a7VIm+lq2khroudPEf2kj8oc7I3dfXDtc
GLln1coPFiOqqkASmihb2Iy4mK/103iAur1Js+TvidGsMUc8mTfkwWZXg0FrEQ/X
Kvyz7E1ThwHBoDQmDKoKww8AAGh1ngi4kwN4dPmEyGN68g/AAtkRh754Nn1Os7WR
kA7r7uxEzc1TcgfTWB9dmE6rlYm2lZOZWZ8RM30JmU+DDG7TiId0plPVvwVPe5TC
lVw8Dm2zgW2QrwcJIVdBjqLhMVyZnL21y0V53hDZF/JTbDoielZX2FpWJljzL8qI
ncYpCF8u5xTE3UsCZ9oeTGdkvi7VflVj5/5sNjmISrxl+yA7tnVnopKvBEL8HZR+
78Dxt6ICmbGN3honvlHIHU7EnzCh2MRAcES11a4XzSA9a7u/g7Hnp8Q8h93nAsBP
PV+ypmLfcyalxzwMeeWPXPMI2FZkGuFlXcXMK08y09cKfV4SSceFtlGEhO9dV2OU
324IkEZ7MHmo7XuX+P/w4iEt1CltjKS6I9Vm+83aO39qLBipolcPtrxBM8B9axCP
1L40H9rZ1X4GxL9lM7MmBjLS6PLBIIfX6K6NAsiIFXLLMVOSbL8BA38fq27OcFaD
eX6fditWZzR4flU38731bOTIxx6A/KOhLmAnSTI7VOyd6810Id/8hXxpXLKMc0w3
EkHNPj13O3+iAVoQGGgxjYwzvp/pDmaCOszt+V+rWJNofMa4THFiIup4CZ7AY9EL
sm+urhROFt/xIT0DPPwnU+3+m+YV+x1qaSR6w5E/1GfBQsZE0Bw5hSWQ5NB19Qx1
zB2PP8MsRh2AWd9nA0dVH75u2ISZmQOLcGeUhCie7aPJK5KA0aUAfD6RZIbMh4NO
O5/W0jPnmvFCx+C+uZkC32ivyWcrV1RbBCcEntMPXBYZXsSfoXgKQfnVBaOT3cye
7mRFwnWHD8zcmCAViMJ57Wu9COr9MLZocU1WgGZ49uz4w2CDLFgiUvMcwJH4NPI8
vInZzzz93Ju5qqX/SdrOxiyWKPnafPfLPW00soWUQxCA8gbVtzdctOv0XolyRgev
XeR4PyoYHM4CBeY+mv5Wv9XOtb1Cq54rt5g4/EyiO5FOsJxRyk6YiSFdtIVr6OkU
lbLuJEv0dUE48qxlQLAe1hHUF7QTzD+mQhFML/M0HYKFSrQrvMuRpBnhUgfuMgJY
s7+kxlmGzgxoW9MGekC8KoFmYaaHUnGGXf40no0PTY1PUgIbeL2VXyqbZYZSjSAs
cYfBNf+lf+mrCnZtdS4FkZd3X1wiwEQmQrgPydwXB5jIAmMYHS10QqZUG0iG9SC2
1R/r9KlrwhC7NQvn1cz16JZ4h64dl/f4DpjViI6BRsQtM1Ep7Ov44c2NiZT3EgvM
I3yrmlnY/mf/M/Q1P4FcUMXuFiuOOajwuRIeSXZffjPd48U2Oaeb0HYIMYOnuyZE
JNZ3qFwBPAYgLvcUqbyeuIow+dh3cXGVOszg80j8GXx9TwL7yu3d3tSWLQMqdgsy
4x7IOip7OD8DHZiKak1VApwpXKdREJcY2rlzQYpAMZDJe6DKoDBVhWZF1DhTdyuR
cEjGwWGy/6KUUgjIt6IXWAPxJWGxdJ8aXnr7PKvqZl6wlOHKvPmvc9F8HERI7ayb
IbTKV8GYsqbIKri9mhqNpq7pkzQMEAqbft2i+Gkic55IXdjcE6yD1lKBqHShJqNf
BYewuSQJGZL/nNURnp5R4emCKHEVDHDKwixLb65bJHUZ+Dy21P/EPTuFVf4vlOhG
g34h84zzJ8u1/fUooXwhZCTEqT7PjNwkmRhQSuiSt4gPZGhnBWPdyPkTudPEGYNm
+f3WkR2kKWulMSSBE7hDf1cTg7lpxDqq7jcXPQRFdhBe6rSQMBwI4SnA85cRjFMu
FhcsU6AQqdgplfxbfhhUmqCgjc5z3MVKX1HAgZ7N77FwaPrqGHLCERTS2kJWF0vO
/aKZrUqVniUkaysYpvJ2cHppT6xuBQHBPUgSwGsmA11oyXTTDUUHV5MzfWjrcCPq
Dv064iZRt6MYIB7BCNdivphufroqAnFOmyvYfwA7vohkX/R5YfJx/jtYX00tNNlB
+0j9TIzL3PhjPp4ocyEsapJuY4z5hHZmwdNfSSKI03QYFCyzFqFzjZhfiSO/hEgD
ZxzSc/GvWKetvR4fCgeGDKRYI8o8O0nO2/dH2VLFe5SL+sDLmn/ScDn6yo5WtCB+
/lj9xvSLVGJlkehnar/ySBifBHYVp20/lsStKJBa5mrSkuWdjh0HFTyjjTd6LZTs
HWtrNhsXHfEejSrXNhok4US2CMhZP7vBuiiqEu7JhUkAw6s92UniVaCJNe6krsdE
7cAuX2GSSitfjCkDq2d9unZeLxRbuxG6LXEdjlx8pttuR+2fRpSfdMvYvWi++TAX
tSMqU0YKcZerzfbAbl6jRa457Ls0bJImigJ3hHcX/uK5bn6i9olxQ+5NgGBUzRuj
k8byL63bxtY2T4jEktC4TkQLlAVOPYiCKpuQJY85akwsCwpzYB6udqIe8favbZRR
MhUCweX2+G4hjRluazMet2p7DcbpWPyZ0zFa34GHfthcMnKdBi3udtQVWn7wLheS
hJqjOQ/z/bxK/sWlXhTejf2dx539Y2CSIlG2C3vXNlEXJBz/s8fsjmGzOhLnef/1
lUeuWDLIFBhLtagiVIttltuS3KtaCtWwVwjmQUtgVGKotNHpotXdLPH/GKu46u+n
TDfFuXJxOBNszXmzgPTPXopbjAc+08R0lM0YydlrRDLQRxpf/U89N4itfcVTpKXQ
nJiRd/rL+Ydad+SKfkKdLU3roD8vE9i6uge+KQGxjciw8SvrSaLtEKoda9/F3IvG
GY2mq3BMRwgJPfFnidOxhCHe7cgACHqh2RGAapq6ge/EJ9npHmaH5+N7fvGM/h9C
nP+iwMBi59ZnJLc50eBA7h/Y0zcBS3mfvji8h9+o2Li3F3vjH8zrL/6wJSXBodrj
JI+Dspk6XuPuvRnLrA8a1cMGhkIyAOcD5kH8rM7zQYPL5rqmLoOkLxeOvbv/mqWq
XwvnWOGHUtfyNyXt3WoHzI4bFltzmBT95wyYqO7dy7ot2eVfSuIFgT3JOJOlMiCZ
+p/U5KmkovxIrGtS2Opvh+uwqmiIIFc4uM/+zioo0evEaVA8lSxta9Xu2WaY1t4V
UZmnNrr9o/lu07zpG+kpBOk3w3CBUlO7F9jaIhKlLzpGKv9ku60aSUEK/zmSZR98
x/rgWm1tX/n5Ek2onmaGRAe9+02Y/Q7PSITnmGbe5O63mYTkqpL4knzK1Rb8AVIt
xc0ILJf2UfkoIAGiw3BmtiueBWXI1R9L5P7sREG2F2W4C/ZCoI4C75OhxIHzl0Sd
0w2MHQwkVfYYpwP0/8pAWUtzQJ0pQ1dbYKqRsTbr3+N4tUNWD76CYDgnBcYGuIpk
sdudOOrPpIwJRzn/bmIp41JrhtCZ7iMvJ7+R0zg7yhe+5NQuNjhzlCl3NTVuo4V9
IK6Htec2KJgvpFT7yW0MAk34loeoZTtUaw9WXWLsxgsv7enDipv34fO+XLzVzGrX
DAWTTs40o3Hu2H/dyUcYbIVphdVP7/8VYyMWJHoJQOfM8zhYHrCL6yfhQHqaefh7
xQHX8RuHqpchn8vV6PQpSF6HA4wSi1TEAFDEbsQmH0NI7TrhaI03ofwWnelzthUB
P39SVIrSnSqXIE/9H/hiTaB1w5NGNkGaZwTNSCBSRxvAjGjbr37AUuQdt7dHFFHG
OOccXyRjKyUDynh8eIdw8alsMR0O5RuOs21KuO6U08TrHaVpCrdUb7VcfCUm18r3
3YNKdatZ6xOmZII+wC8ImO/GnxRX6stwClANsKtk/au+p/4d2stQ+HYXAWE5ikur
x16LtGqFVoAQQrpeguw6eljO/kpCT6/+JIMWXgUACR5UhQR9tnsGwa/jaCYF9L1E
AmmXSD2p4R/2WPQLaHRvd4vODZM+N2g/tujfZ6dyxzJSY4eu+ZPvZNDcowC+x4nI
AO3LHOaiOnvpiWdMQoLYIHkQwEOH9c3aAUSuGQpRypT6fTyIs9S7pd1OmBVJPlmH
X4i6aBgurbmYDRZDU43Pueirey2Gp4LhVDNrAbexH+mbDVvf3HCX+unbGEAnExfl
00gN5/AXL9ojx7q1C7afUVWLeiKVng8me5zXxUD2wA1skrPMEB5tdP8RpntEUbjv
tKYd1Jr/+Q4PoDetGrE1NBAo4OUbQsdNoxvLHR16S9Q4XodtnwboWL6rmcCDlQsa
Z181mIiXy/OzbFd+fyCBDtzXAMr0Fgd3CwYZpOSeQ0FS4Rtf4p6Mwzfd+lGbLOcq
HmTAIpD1QujqqBjLmf71yIYPhrvxnda28WnEf77nj4JQMXbXEWTbJPCeFBdoUcyM
vH3VjnfLLz2WJ4YbgC7VsvvUBBo6DS56jfoft5UJRNKIXwtWwgNRl1b9OJuySDap
8CElv7AzM3BYgoi3cSeepovrWEw9OI02JCOGjXEC1mn5oTtGPI/POmRnY4LldKiw
WrSbCbBHlvmJCHDjhPbz7sjfCL7d41RtoNrTZmy5xAJymYqaQBajKdRUYI6JNQjZ
mchQeipyDbpv9JlxsH+OiVosPMX229GkgpBwjnqc9x7PAhwyS0Zn6GprTuMYpw4X
Xfr3HctS1I0V6uihzd/0/7nryKn3BcU4Rv1HWQ+fq9kRyVCDqV9uYeT53XlvozuL
N8UY09AD7SuubtdmBdepVSJB8uv/C90RB6aupR7mGkt2k7SEcyJT/WARqbj6CVtz
Jn6ZBwSnKJYHppZnNRcRNBuWll4xG6gO2t2XMjUFpzS5EzZuQriDTL8HMmv8HTiy
3RqWoUrf60DfuwSICPHjs9pPPWkEWtZ2B5Qg1EVffrg7bbXaJp2lpv8UsxS1eds1
aK9VZUEw1knLlH8w/4XTzgps53yexHbXqeaJ/ku+cFVZrwWR8BVvPemn1TP/BtHQ
fDUfs69wWUzBOz4787YjjLkY00sTEukxQO9UQLnZfAuUtBOTdL0JRAC/TYoNETV7
fnKlXSQH0YCHzuNoHMCOpUx0gde6Q2arUx49G6U4tsHdszs5znh1boS4Qcxq7E6u
8JX0UrN0zd3wh8m0WHmsQXKUv+dEGPgF9KvkIOSjQwnmDoQUb24xFDQhPTl6VAOp
PHTNHwsmOH5MTiCMILWUa+Od/Vnq4r3BhsgWX5c60EvW2lviz9K5yyXEGA9Hd+HA
eGLx3ynpxg0K0GqVhQdgPz2Xrjx5KsOObkUsJrBlZt1DSFuaf2+Cv+196xhWWzQ4
NAyqX9hGenGJLhmU0O8Hk7JOsPcrjFZkGYPJfdItf0KFaG5olFAifzwgAjES8BSa
N+S+NXpnrTAdvfk9CH+S4N0VWBZFun8HT12p07YXt47sRIRxJkLjXeanWFWIFyo9
CzIGyvaIXb8lPbEWBWuC7kw/7YA2M6QKdcj9/vtw43t38clqnEEG11dDvbnEGuxa
RXEA2M7rKaYc9n0DwPKmTASs4BcwaHT+jwlVhtZdfAFTNaVpKlco4FM92cwf1dmo
QIYZ1V0qJ+RoSYmY1Z85qhuKbXaU9NHUdQ5wTnWVSs34IG2ProSeQhQLdWDxZIm3
Vr8RgUBV8JaVTdj8/EkX1bbY8H3tei5FDxEC3RWz6p0y8iYMaUCVBIYTnCfaQDmi
htvDExwJgG6+T5ihviPD23tVF099/6Eq8Udj8s8KOzO/wgZ21fAaJmxD0jcl9vCQ
nENtPwZ/QNJrRL7uh3KqdC8PMvDs/r6P17IHkRUbgsUu0K3KwOhXTlYSLGvc0dfG
WO7BpbLb3IvozRVWGmAzOT104AZslMQ7m2vDMaezr5h4zGiKpqhu5rfeDwKXL0mk
Brc9mCcWwBaVIhquMY9pztINUTcMQU/ndu5WOfls4roZZzYpzlOt0zW9yApDbbu8
y5H9F3YfaOly72xCHBI+hoSd2p6IqhDuwhmDh+/xsOj6fra4tZbTP6s5mHjidVrt
xFRSr6hYvQzQKoywWiZQwV+an/K9iZ+VpJhY0P45MToorH6DfPL+lAJkYkYYfbAH
YoNcAbokUU9FKLSUMRK/Rw2dDFkeheYn57XHA46gGKoe6WY9Zke5joH6OliND6WW
HeqVLJJxy08NEzXMI6+jOUi5pvtq2pi66zXuD0CVvAOkNccNBEx4sP0PNVzsxgvl
MY9nDpvXVDWRFBQ/UuxLQtOd42kJgafSsYP6SGdzik9HFwOz3ehBprW9NnA0mG7q
oeqkmNaG6xz9Kl837KovVblU23o2YMl4aiCbwnUdFSxkKxHfOpTAm3VJz6SigsVN
L50GWpCxkCfIPzEB3ApVo0wi7/ehw4CRFPJFrTM66NhFpPuw4SlrHuEsPFgehd7U
mcZLewZEh8BQ85Ga9Ky9u/qTT8brhV7CHJ06hnWbm1oulDkymwMC39MXz/HBuWF/
RZ+sGfUu8tIyqUKc8SQlt692UKb/Lpevfzsd2gyI7YeSQsZsd4nsjs4HEx51ELWm
up5agt1wiKJkbUGsgaxgIq4r0aKBiMruZRN/BT7b94J55LrtcUyD2GzOtKw+9aFd
2kfeAVYjXse32LR5FBMcL2N0m5XrPjTAoe9biYMCNP7XAH/2WYG/Fh4m1LCtjmXc
nQbIx+rzSvjhawFQk34X+KBRIN7L4GBlOaljySQpC3nGJoN+l0ePUubryJE7bPjM
Dy74/7yuLUc1wpapF4jkWnd4N3ae5wweVoRkM1I9x1ieHBUyl2jy1z/g1HUUy6qK
eye57eVP4a6HN3PgH7HOpE61jSHKRS/4HzLrY4JfJrJfMy9Pvg2x+dKbORrlTmeS
kuv2jxemryICcfRvxM135BciFneSAsMm8pGSk2Tu6XL0v/+eTjm4x2oZIY/XkwYr
V0IVC/PjBR+Dqh96zk7O9U082sh4qR4EaC5namZzSNKCM9tFFwPcPW6JHzIaxNup
9ztW7YIaPw+8jYf37B71Pst+eY6rBbWx68Zfka40mOW0t4Wh8xgPZqkBieMg+DOA
RKETDizbl0uHyCCj+leCynynsfoWe9VZlbmGJwaD35gKpzTa6xmvg3W2NHgUpICi
hiPHOzWjRYEwkhpv+mIndItOIzpC3VW+w1ZezgHc6URBWRDBNoGMGeFIG7lXMfvB
cTRmcTqmI7dTcDZnKVHxUm5GZn+X4IWdMNrtqq2RFhxu9BWjA/DtE48bto4Pr24Q
hvwaf7z63SqOJMOZRUpum/OzlC/50vhDttqHfbNE5fMH9hTKVuNGgq0u2yh/jcMN
PDXNH5KEwZbwkoIFh8rZBE/s95vUTR5o1WO2CBe/l0lmlICFwcCy/fzqBFDQMn9j
E5gLEMdivTCM6E7MVxagH2tHi9N6GpBseXY5S0AqK6G0nyPEl0vcK6WWC/OlhhGq
vJyhvgxQcF+/xfbosYa36bPb/fzg/KyWiUFpdYGtGuOcc0c789RxbreK6Om4Mhtr
E6ZuLxgLG0FgcPk2jq6NpGZ5RnKc/TJGAspquUl0wjZay3Lir9RBmjll5PDXcC12
YId3jnT+XwC6Aav8yzLWSnNf374HmSYlauJieTjp2/zh89xGROh/2Uc4vzVzBk8N
wMccw8so+0pED5a0KTs/rzFBXjk6gKUqZSJTmOom+w8IGwvVapO/RwIWF/e/W126
sfa+1nswIzWrre//AhZjAlxd2xgNNZOrEpmfNbV8AOB0NC8RstDoI55x9uuVBKyE
FZOv+mtpRzzuyRKJTc/LSHW0dubWLggdPjTjy6tAA1NS+6hzM9YJTLmsmEM0mR4w
jYwLgMIJ8ExBw18xxy79VOq0D8prghW1l/vJjskwQOvAJJB8POhx5T2QJwH4ZLpJ
9kmnU5bscVCplTeaaBJMcFp3f6RE9Vo3LLkgCgUohrCvOC+PD711SHAOCRxnJMRW
KYGuxeIQsCYnngVX7326Y1YLU4MFFwaq+4dTdE3mhoyXq9CdTACVhiy73BjdmNER
a9omcQxGhxM2E40wqYCvD4J32uiNrUfZbTCRprONGsK2vKg947ivo1jwsFN22F7E
KfRg9qAXy35BqgxKRmqcTNf+kGF6wa95a85i9U4L5VuuSANL8Y1Y7Pj3uLpkIbzu
iM7AdmpyY9r1gjUKxXWwIaAfGFXiMTijihs8cwM4NyU4wkawVQRwU38Act/7y+qU
f1GaamYALTcdCkkQp0XdXHGic+jAFEb2U/0Oi4PY3t9H5+gW4dwreJhZWA7lyCo9
6s4fE1NyKjlsgIE+tJDYQjf/SbxkuJ9FX1HNhBP60r9/Xq1BiXNzK+936uLtSF7W
7iXie40hq2dYU6H57akGtRaev+uwvzPJu1U/W7ZPCWTjrDESyExZZDxnNU+oWbnC
YqQNOOIJJ8LNMSxIG6IGeWTfEUSOHB5E5cCsNVg8pVTbRG7bETBwKUktVcWWkp9U
rrVk9p+6SH1vZNrJeYdLRKy8lK2EVQ5mMw1g1NrMVMsWRqdrxOu4C/vUKL0XbTRl
31w8PxcfhGga07ZH34Vt5kkpdI6wP0sKHQM7+d/m3HOquWVu3wXXb1O8MxV+PA3z
iBbaopqdoiNEaVug4/3YaEmSCDpd3lN8qwFzKSBgSuhEUngbeRSpq4as7vSrEI9X
9vc+Tgh+MUvhkO3HigIEc/vNi/hFZ2fPUCGRJ+WLFFp5DiBSBB+W5q0+nuXI7/qw
E4dnqhgLDmsn0NCTKQ7KEqriVXr9ZULEaAWLMC6JwwgJVUB0nnLcOstOrca1twUd
gcvBUObXrezkL9K8sSrOC1XBVCKgGa23UqZw+LZ9EN+hUHiJ3DndQPOkShUoccNr
U7HsXODVfvSCQlhP7phDewuq+XmXVLJGW3Zy/KIEHqq72k/w/t3HSVhTFvsjbm/l
64txoYhYFjP9QJkZRxlGugGLrUM8pXWk0iXdeBlRgE0Fjm9ZFQLjTDH5fy08Mp2Y
AClPbTLG7ZzIW7mRKdzVk/z/ckyAch9C7VoOYlOHq/Vb8hRHQ3Pwqekhdqwwz5cu
H15FXs4SY1vdtYsQeoY1AfFP7q2+sH2JWJX+levYAm2MMivm0KasvanP1jkBAFO6
F9Fc6d1OltpgfVYFomFijSUj8Ac3cY2ZTZ5BGfTPsG03ttA6l0GUOPJmZa3dZIVV
Kdg1N47/OgKyUOFtQpbHT9Ud7tun8AdkU+VuTdDxl727Qu0zooEWEqfwUHTnZ/D8
PF8sdhYRzxf/YZ/0tUNqR3cT7DmayO/mgGrXzYVF6AwrUv94wpK2tLzX2w1Kgrol
XFCoz9UcEslpgciLoS6yctJewf5Wkbb0m2L4b/i+fA4jZDx7XD9vXLqcJEUS9OPP
ga3mQwjhPX656eeQjfQXmrSr/BTYsQh9M2zys2DNnYL1h71V1SLGZBz89vFutU19
aPCORQCwa+OZcReo8cuiRSC07+W4VzzYrfeE871xOxfIYO1fKMYDlrhfTXfCfyhn
5D5WajGV5GD46BcpD6tG0vXGRN/tXYpIOKranv6KXEzL9J1IzxwAsRWSxPkE/Kw9
wTBUJrGmbmC5NXfToJPxHhqWFWzm6MwaGRE3urRadwAQkraX6+5Sd77FEN/cpptM
GGERdwpS+D3uaVUWoTfdPTp/2CkkMBoNE1dm52mGfOqV6w7TSLMj7F+Kj5ozBW4p
kdRO+mqNEroWyqfFYLH3fcZ2sn1baUfYo0kEbDYtr4wcOQ572VQC93raUv3Io5ms
BLR+hNlebh4CEOH3GcQMZdlYGeuFg8VRfzGTPXwfdECseieYngqh2gLNetw1/Gcs
49KlHXtxPJFC3rnOH+lF/8NEvvqi+8XIbOpBxX3qe4o2vRzqGDgDEsrllPa2RmMU
YQXn1ubs3TS9BHfKlimir0CCwf8upVH9vxdieej6MXnZB+XsjNi1nbc9OKicQis2
+ZSfKnhsoEmCRXQIcUydTJVmgYuuJZ+iEE07wTNBIXEHmdttr1LuDQ5z5eF63kTG
9ssK5k2tBrF6jMOyYu2B2RmTtZFlWyVM8jSXXHhvNQgSu1TkztJpcbWFGs2aJ7aF
ipY7o1C9FCcfNj/fpT1dwIydt3NjHNWdbFsNcsoRX95enOk3/B1KGlFR4WRmLlOS
5se3f6Y0slvAGCkeeg9VA9QMdyIJgH6eRGN2B1VVxxEo9uloM5Stafr5VPg3grSE
0YCuqthQ/4rXhWHSAVdyFIxQ+ztQtjFE2tUm/CiJPzUJYgEv1Ptf8Ohjsh9eh5Zw
gz6cXRhSX7NAxFhH+EmNbAsQv61HkHXngSGoR/qNdWOW+F48LtMafE0SV2KwsxRj
wIAexhf3mbDQHCaZ1nFUVsmlbB7dHkWBnrc7IsRod59B84H8uwJL/xX3ShjxYQ4W
UeG4qBxKj4uJ26BjEGuBJ99lq53jEOglYM2yuRFEHibmcQJjyIcsIRsJl+4jVab/
/G2LDg2HaNNAh839fybZ5FGuHllwEzM9YhyFfmaseS8wo0thZW5piGw713ekLgUY
Suvxc7ca16W/E/Dn9N/fStBYP7ASWIWKAUk41X/NdC7b9OB4IbUzj6d4gH3kT4Q3
1uNENAvem7w1mJnk6WSvYSsU0kJh2Qf1opCIDFrfFlpYqOJcb3Yv8Cf8Y/7c9qKS
MyrNCjmcKbbejtLnOK5IMeOdkMAgOaLRFFBNWnaVOqgxC3YbxzPyxwEcpNnS9jPM
bUsoopMsuOpMF0raBc70cyLv2m7zGHS74iL5ICjOWE80uxQnlAcfyfld0VYJ92Mz
hMwRCnxw7IRnbTaT3hjfa8RQpK/UN9730CH2CKCEsvxU1DHBJEjxu3ZubdjmzZ9A
OzJmXHiZlXWDcGNRJWq281tO2C4eh5qoMVxUHrrlmEdlwKdH75khmWKePTzKFr7i
3dgqbrSpHmZUa7pZqi0WxGDH2l/Nf/upwxphKlowq6ieqEAT85fhO4bGt+u26SQf
X+tStOsRJlbv4GuCv53SDmu89d6ixve7c0Vaoc/dcLCo5yhATgY7rGbdvyWJ9zYq
+q7fA1vfXPHkx57ZAF9jD23E1tJuejc0Ue8jZqVb3po0JQOVAsy/FrlcO25kxG7M
rIPCzlvYz2wuSOo6XOVSoK/lJV671jBO5/a90jJpUVebLNcD6coQh6e3EKewmCoy
KzSzu2+EjAyqIhJ5ZC93BNrCLUfVS0GbbrM9/HwRLUI4yTiWnizGceNVe4SccW10
ClWeE61G4u9Ok2xml09IPR4XabWkwFOScrnthczb+8HSyEFMsi8Z/mW1IypSqw2R
83fazhBNztWkE/TmYxRfUExRWKu67SLeHuMpJ/LklsvI7yYOyEMgZmUwuHk+MBG5
i6rE5mKFEddGhVzlEPHmM+cxjWy9Vlpv8tMYIY2wZ24b8+k074jkV8GwV++oIRN6
SKKb0dxXyzA70LzmdV7onwjc8+9Y1TVdXX+nKV2gMi9kYgY+hmfxvtwe/wTWzw4/
ll23r5qBXhDPfgsiCletzDq6LB9sX+iO/qW9CkYRwMW2Onl7+FZsCVI1PqghuxmG
/U5ug3leL28t1c9ezlnsjvLBzRApIm4UvYz5PrKLzpwpXnVl2X/NOi4YpusOxzY5
d32yLmxs9ASIUTU8uG1mEhHC66VU/OVzofDubVloJSFCgx/RhY/k/08SzbycR24U
hUbaUWM2tdky1u1AlJ0DTXNDEYPDyqCrpSutPlQuFQg2a4IqK+qK5OdeS6iwZgJH
w1zzJGusD+zA5y2KUKtxo81Mx4DquQbP6okxpFHwa+mk6IRND70g0wi0Hsef3Z/E
zW2WBKfX4+2GOGl7YpKMYJb936BZ646OuVgYVo2SXtZH2tT8PF/3Fh0SYLiJUt0Y
hoBNsvzZWX4++4NUJm6XxMe3wGhxSI0Cy+fVERQoQ9YZNtIZ42qoqohNj4/az57M
FCqQ0qBuAiw2Ivl9S6TIJ1uDmlZW3UU1WjqukuqI3x4/Xph+iwGSWsr/S1xb1pRk
y+jgujVNRD3q62dA0dcTYXMQs66d9JBtVtXGuzyKjQTCZNS7TNfmU04D0BgYDlRB
sJpXa71zSvx/LLEO9edqDmOzt8RLKnsI/Bl1HB4tISjCtzpVFM45VNlwwnEExET1
v04vJ66VZYkhbbGhXYcdbONolNN6OCbsdK+FPYQ+tJ8y/xtO7qisjOlGGf5BVYEj
feuVS0CXQ9H9xMsWW2FYV1yLYMHbBHnC3d0kvgiz8a7hFK3VF+fxwBlOhJ4fnYbc
UMxYX6iXTu5F/fXgPilUyRcpapovNNck7Kt+zhRG9siqLipknubMLpkKoK6o/lQa
PpiuaC0LMb/rINx+LenU1FYcue2ZnB7s5Gk61QE7DG0SAnhXvPL5A6TtPThDSXHC
/lTssk+Xph3XYNzTA3DiKsyznXFNey0nD/YOW2Ynz3iSh2XxoCwXp8YSIG56uRjP
OXUo65QO2eqyffEAM5+7GJZzyP8Qmp/mn/VH6MIz/6I2ZZtUudjqsbJYEEIqOU/g
Y3Zv6uDJxIDfd5DXGeONHLYtE4Ap0GQjbKVU9Sc0HKLB2uqL0KhQ2qeTXVkW/6tO
Mb3cXUckr8LAWpPUZzsUvgB41zHKKAaOKEQHUdILULOYme7K0TXa5biA+TuTzntV
U+sq7hV0AHrcewagPzXzHy3EYaU9Uvuft/i3d0PO1F0o1Gh04rTun3ZYFBNJsfxS
WGMmVfAQaHKPczmYDQ1TUeb+oqwOBeAj33STR9qOoR2TjzQaXJGnmkSvvwl+wsSU
h4Sc2PvMK76+IMU1qeGrAcmoeS3QZFhllDidaQuN9nOiX2HCmzFJBIwePmSRwD4b
qB5aW3RyTyq9xTUM+GTSpQZrDKVm8ZZDtAM9ukQpygRsaILHqzEDOBCyWA1gfN5R
wUE/qgGrcd+Af8B/bk/fiq+KDQBkysELeOFjHo8kEnkWw6fsF7NLRFhLJzXIe4iF
KUuE8B2Opwe6R17anbVkhmBFhIP1AdwAOMZ4ESFSiW32nNdyYAJYrgyHxZ+/co+7
K944XHd5mWQw3krSGzoSqd53AJWVHr2esAsADaGxuGxqrapXH1J4SugEu4v/VeCs
aMR/xx3QUuQZfuQIdhNUMAgIuAWWuEpykHK0VAYITOqv6E/q1icHdK0/xj8GrFue
yqzKOgj4e+7xoDPFsOykAoXkCrlmcahXW+bgTf4FZZ863OhTQrLfTRQDKnUbPzwJ
Xo4wtlPGgH7UllMpa5So9dypoLPJbCmq5w9R5PXVXfuhclhx0ce9r2rsZT/bTN+a
2WEoEmeH8m85xKDXLXFyR9epXlgYI59QlBO5rsOxXxnXp9eOmOUFz3HGpsGOhajw
Xfgrxw4f9xdXvQBwdZ1d0sigjC4VPV3zkNwBm5eeOI18DsA3yzGJfQ89/7g4dVZs
dSnwfiau2gEykAgiGy+R3r/mZC01Aq/zki/YXesBJzqP3TG3JIyuMiSVUCx6aNRd
6Mk2ad5IL4S0zXZq3+O1WTqsBtyPlg9csvcNVLspXt60CScBnfZ2py+Rw13qYolE
qxkmvyIOBSNcCy4NJ9vDOCmAHKFUt2igyOX0IPLrN+/Hc7zWr5Ontb9Z+1Vc6NCt
41wJHkdQ4M6bgraVVDREg4c0EML0SeE/Femv/UBYIyIODwjABA+VEdpFzfD0Lx59
gMrDRQdak1O6NLHErjg+r2Yso/IlSvat2gwVDx0OXD+Yc3QkrPqrpt/8sWEKauOi
rOJnMI3B5sbgWBpIVCYoL4fyGsxF8muRvgHE24Tqe38gLuamKGk8cfgi3bK83I7Z
fFkpq/122rlN434ZFXRBnhif91aAowhD2kYb58qQqsAy/CBlJlvF4SaIlItlWmBX
JGl+JLTmOF+Dt4dZ9LuV2SrH5fLzq/D0yplePtvki/xjBGuFzr7oz3kG+BN7BopK
UIPU+/jk51NgRJXZk/qXOSq+pmK2oB1FU+fccbe/bQMAJ4yAuvojZ9EY36EJUFZu
wVtK29DqQ2WpNYLDR89f0Sn0XPFXcGJZrJ+eBMEoeG/FkAeuUG0p+5S4CI5p2l7j
mP13JvGOk/DT3ZnAHSHeY8VSSneJOr/cTTOBJWj0G1F6EunmLsd7fegmZ0on79p7
e1je8dyC1x2kHrZw03H/M/AAeZkWkroB77x6TwcGHX5qDFHW9ilIUI8HmQyH+bKC
CgnAIefSj4ypgyjiRiefguxTngWM1Gcd+LM20kLpJP4g9dYR9tvww/nnupIlpqC8
TDunGbechW/9syZHhLXj6ax4IvLOmgusj7qKwj4hOZl8BShCLR4QFX0lB4t/LUYS
fQEBQnuf/BZxWnsM9D3Wy5AO3Ok/5JWRPm2bxJw5SADhP/9UxohmrlQzCW5/mhZN
7CzgKmn3brGtDpVK6WqiUAaSd35P36PSx3rU4JZBQF5QNMbB4kp78nsEPsqZBFzp
9vx7VwY8yvsVRF3VgJ4CZeCveoErzhFVzpVsE/M/5qrcIzLwPyuBkxlxhLArE4zU
/hZj34VGm+aC29CT1IZNe/EcAlpqaRZF8P5doJ5MkLe/3LUgpc3QyrUUw7n3KuTU
DUVq6WtR/BwBYxgTwEn5kub9vkJ+ZE9visiciDVxZGLntSoiVc84F2Vgh9X3fv0r
qIBZ49h/gDBoGB6fBk2eiMRqHATCstZQ1mNhdFz2waXsgsp0VfgTPcSASel4FTmB
pGKvFWNdMz9DR8A6cLS3DR7hf2epevxhtZY6tnltIeLKUTUxK3SXEr7hWWNgTn/u
STNyheugtXdx/zJl5VuF3EPqED0PS8LJHSiEy1PT8mrfzjdmFeQ35MxQb9vaS9WJ
PVbHbLriSKk6jYarcQYwVBaz0LqN8MDWGAVcgT5pqvtxlBb4mUIJrEgimNZwpEy5
iTMuP5+AZz0IBMDaSwIG0khXWbWgCXVOpfwrNzuykM6uwvXODDkFi6RWUonsF4C7
JSh2kIuTShlrja3kh3FgAP59X0/dW1SnLpI2eVGRJMj4B9tTzK6TOnfDkossj5VO
V7V2buyGwJS72Wv7Xg6DldCGwC5wF39u2YVy5ptekBnZi6NzJSVi2XZy/cfjXAob
JFu+tVD+Bc7xKlsOb3Nt9dU/qyOdVuZKmmz2vvFEGpgrNGywqxkHKTn4STcQgGMU
YYY4ShwkcbBwtVgCKzn5N5jHuuTznWNp9VdUdUu9t0QmUG+OUF9qxtfC85sDBcll
vE7z3tKEslUgZyXf2gmbVBX1BiRzSEkSB/1KznbPqrHG51+LGlLwXDLJ8ehG6s1J
PwJ1WOufXQnt1Sj3+kTJosPSVfXlycNbl2c7XvRPcUaqqvi3Qdc+dvakmMZxE28H
re/5LqNAeK0xpUXQtONv5E6Ya4iJ0RPZzmeYjhrMAM6Qw4n29dZ42eFdouAw5j16
+UwaUKzxzUR9eskc4geBIlC5MNDNHSNBozynw0zyN1SStwD2WhdOZUhGG1ZWR+Xu
sR7yzeB2PJW/ZWIGAcrPyodK9qw10UG6el9EEkLjkimDGP9gTPIoLDM4gfogY7yo
BhHb5vAeeXMCsKelVXvkthQoYXgCwOOY0tEZFD99dkDfJ6tgxpi9cpMUVaSmQqHg
0JwTQAhrtmwiRfILN6Mo2HDmk9IQ40Qblv3nAPaMOD6NIvGSXK8Fgm2TWDRS39Da
vSrSvNyg4wRZO4Rl7cyePTJqV7a1tI/4YEkW0RvkqojD0INX763vJuJtdW0dSZgC
5+e/0M0vPrPArpAXbu+rHYOVP0Sh+RFqeHLYYRMimAYT38xeiAJ0ZpYe/lGiQ/TO
fKwhVv3SlkTZC8pcPSfQqNckyZ+rXcYdCL6iXIdtXQMCGQrEsF6sI+2KLDfsxKs6
FbLZMhahInSLa4fPbI9tn188r4bh3Zk163R66zQ3Xw4Bodkz8fdJg2XAXG8sYnvu
BCwfOdUZim5AIZtazUyDS3uliKUgZd5aQTvHuL7Tb70wgdAa3XQQvp+xibTBnbe+
7EKXb0TMzeFZqA0pfqh2Fb8b1EZ50ce5BpGMrI0BaJpMj2jjc+DuA4I+DxpYuKq2
s6OO8j39Y3zZTQb6dp7T2Gj+TKo+rdPkX3riJShrYxUnTMDg/VexBAkHMRxk/vT/
O+IpqhLudUsw40b8ObHKpvd4Uusp791Uhfpg4nA1s3tOfxXAV34L7Rf3sC0sRma+
Dogq7O61cnbXRId/Vy6R820iQWwTL5+YsGw0cZXnObl1lHqiouXvOXaQX3ekljDH
71De19hLvhFLpu4cwe0ZpThMVTvSdDeZLh/D+8Z1O4J113jriDpo9ByUlrMIcfae
l4rLIAZ9DLJ8S6xxpnsZ6kFWChtXqdjUQKyI69W0KxZax7B/hrlpNeBJRxslyn/M
JcQMQtN/K2POueHHJl2gAXWkODQmslO2J9pkkSp4USsTyRJCFM62I6wDTFW8Ac3J
+zLsIPG5tjsuKDzR2BwlK0PGKCdC+rE464QfRh8bwcmPJM3KuXsEOsTwrIJ9G3RM
8VFT9NHMgWoUHA8qc2KQQijQL9XB6NCCZ5aLoLGYXvsfSMJldb9Z3zlWdYi0//7b
2AO6jSaUb1ScSzsF8REnwM55QS2mBI1FlCODg5eoieckGIFCRGUM1kJ2Xne8ZRfC
bUme5ciqaLpmulufvf+QzqNultPlKpvi2aEg6i4h9ds4BpqaXADzZJZYGCk6Lln8
mJMVtA9VF53OQmtRu+RgxyWGvbu6o8c0eEz9pibHMoO1/rhHYPh/67d8tdRoc2EC
M59hxDbckiUYCDFKiruxWdtCNsgMsT05hroPoFNHanXfpN6TAZmgPMvAhgNYRStF
sH+pvi2Nl1ylkfhZitAYuYIxNn4yNqrMlXK6IS9UIgXbnDvdWAFinh1NiD9NrIjX
ilzkgMCFphNPMaT6UpDDhDKSB8Vkd9rhO28bG/LGde6dqu7PV4PYwdpgQsz5SgFS
t7tuHYy9NJt45rIUWXhqDZY4UFSAzXSoCyjTJxrSK8z9VpPO24NRb5peTEpRuJUh
rVS2fLaC080YMBXbGrJIo1+CTkYOsVdgoS3XGeCIMLVNYyLdSy7fcEwA8ZN60Uqy
E+7aXSsDRubdtkk8ANEYGeI6ltjk8R3J8PmWCKPkkMUsd6wFb0QW8WdChlL2QBMQ
2IE3Ei8VWzhvJDBrth676/pF+CqqdhsNMc2tQ9jZWGQkFF++tD4hA1sOwsVPQgjV
qRqUmBvPXgOQWX77bdZzmQToNtIiceB6qIfxeevht5soqSZGz/5Uy79L3HfRZTwU
hbXrhzMVGNd0B4L0bwqvQb9OcBPS9lURr4KHoy+LQ5adxF8uCQIzpVpnpuDLDeGn
NEvuED6AqZwls73h1ipSFSNi721PjWatm8AqUGHitc1WGRZMSWkAUsz8nhuFQ01m
wZmLmyzgbl603lYlkl9MT9FkSJyM0WWmSTMPk/NMpErd+uahm+qah4mlm10ksRbH
90mQYOuzeOJU2rGioMWoKIQA/t0OBJaTKYgnIj3YVgkJ9PIgdxId3PzJaLDKLMH+
3Efwats328DObQ2gJaTv5emAlVkq9nj1Q6mAfcXOUuBz+iEZN+JnrfjlVTf+c68p
FJMemBlNiF8e/qNQddWFNUee5aW1ir1zloHq03yNPppg7FtWdWpEmcdXiVRH5e/Q
b0Lt/6IfzmzJtxrSWsxodiK8MoJCJgQEp0oO3HtYaPk9Mze1m4RjgRaqXlg0EQEW
R3IZfW/eilnfeJMqBCunYrGk69Cy9oFBJGG/S9Yfv9rKtv6hP1OjRAQhl6sOY6be
wQ/8A0wrJuNb7k6sSV2j05A9BpPN/+7hMfVSev+RwjLumkoxby/AiV6mIL1b/vWi
sYU3dNbf9eEP5lKgkKclqKm/NQET8lMlXnnuM/45NcWkHg6m0dYmNX7AAIJXXDfY
rbyzJy4NEPCY74mpGzVcs96e7CfbtTNokOIILGv5yLwJtQoT/E6c2UiTYOvYHw9e
TsX6O6GpQI0mCDh8HEJsTi3wQm2IKi+kD0RZO4j0QMShNahf3GLoLokXUe4NIXNn
T9R7z/7PTX89vtYxxq2govhX3DGFeyn95SCz3rh7FNECLM0dIYRt/MVjw2zPaBP9
91Fr3lseYM+L+vK9RO+4/qm8ReOJWvOcGrnwsnKHayrmjyTGRmTbomlH3lkY5EO/
I7FI5J5dmELvgBBRyBjO4R3/E7Guel3zChL+AoENJPLuubMlu1Ts/xJne7msZA7s
mmRPD/1OleHiQ46P7/x5erdyq3+JylgBBM7PuRQU3CeupI86Hmo90mYksK/gQmpe
ZadiGLNXSpSgnJkfA+U4pJK/YLT3IXJAjGe5kUIUSX1S/ygp5pEvFwAJEra1v7u8
EjBDDUWGzomIsu/2r9m/KRWDmFwZ25ofcivgLPuRdXvzJTsuIVUX27eJuOWX4S1L
aZrnrbukjyEdiwwjMGxSa0wP+fFKnypnJHf/1W9KcmN72Yv1fY8SPzm6YMYzC/nH
vumWup8gqgB0fbYEU9kxiMarwSQw7jaqzNYs0BQmKw0Hwsokcc+SWbKkwfHwfpwz
H0bydE7pQG1DPHIZeqr9IA9PlkuC+lgum4+r5hTyli0O+LLbQJV23tchCuOLyw7u
HBWRUCwJcKt3RgL0scDTIdk4IAvX+vMflKhCcfhuwmkfwar5kMaDKyG2nNhmZj4J
I6ANtrZ0jJtsdFJ88ZE09rYvadbMsvzHKubpDOFV6+CDB3vkPEWSu5msapdAUwR2
5ZYsC46xx29a3CFu1oHszKie8JV8+Js30Tk8qNS4VpMYAPsjAEGI/jkNaRO0oiiY
FCBoE/FRxfTxA7bWNPs65NqHQ05HDB892p52Yi72TJYQuMot0/qa8dG10N1zLngC
B8n0b8DrgBFGKu8Oo2vSgQju1OjXZYCHW69mo0baW+s/Bgu1U4yTTCKbFc9mCp/N
I06r2/dJ+6PRHPOvHknHSpW8Sr5K9ZHj21ArGzLxBjPp7Yg6mA5A0YAWkD4Sb/jQ
B5iEJ1J/1+ChtAbEy1GmjycsSAP9fRf8dd+fVMlYoymGtZZfYdJQYIrk2vp0YTRy
x1cT/XEw95m19WDt1MXzmdSOThHE7WeG5WTq+d1h43FvE5QNSH3yBIbba9XvMzX4
9UDUPiJgXz8zARndPjDPOBJkNnbnXY9PzeslLfNWJ0x10SFubvEmDwyGx1hpIbBg
NO1jCWBUo5yrT/eONC5+0FLi3M3ksAytFyHC/T8DteUetWAbFCD0mJ/8U/ZeG0bq
rBVCinySO5HLtzE1PqBL1Y/+Q33JIukkhipx9CjPLEeWKRrJl2h27ce9XYVJmhCx
/KpEAAyEFD3xa6G9mgZe0yjRxOrCbSZAvIfkNZjznxUSPA06O2sw8xYWdO/2C92l
Br4BAYmeJlc9bTTPtHKX0hCwV0OGApbl5eszql21PiKod8nZcQQtNMkFOxaAJrdl
DNdaew+nGCz2piURQbd5OB9WCGmHyU8rsHNSgpAenu+LlIEj6WZPZfDVDYNczNPx
HDSnWkOeBNvG/t0OaWO/OpxczzTyioYZKDtgm/A6lZgrRGcBYgLDrg62JD58jMtN
8oY+USTLz7ggX+7AkMPQ/PEOc/fDq/l+npEWvWlQSk1r2WGzAIyYlY/x5YwhZMM4
nTIJ3V2/4JhcXI9/6tPOM8bd+zDAb8qvKOHlJLC7YrSE7Ukcd9evqBGdzkb81AId
r6ahBxPemdhXO1+ekemCO0JWLabSExEAFbd4GoxnTKtksbHW09hZJVXnQSPZIRMu
I/tKYQfVCxajMnWOnZctceLg+oDXZ2zcbnzJku6oDJHBqV/SRnhD+GOUtoyr0/vn
6hbFsVcPnmts6Pi2iiwIK7CD7QEaoZ9cEFxB0i5gKE+MFqjM8H/8BfVh/F3NyoVt
ETJqAWH95vku5JSOx43vMQpVo8gkTpX5G8BtjmDSVHUiXmitoJwF7pu2qTGY98ta
Mv3VwnX6HmDH8LZW/uc/C+ddYYrrX7ola5P6Xup9Ah4QXOpTSDntL0eLeI9FXxDr
d8AQ+xqFGoDcLLfa5D8tV9KRkblVh8nnJ06fImsn4dkb1KAFU1eLFX+94xA6msGu
Qut6eycYdYpoJb6oZOfmo8zKvqmoi2IoINoSbkXazqZ32MzskGOf9mVKG/2OLiPv
CTLrtieVWPjDD8tEfj6GfBAjbRvrIXBOrt/rXPasgx3SlJV/ufztHdLsMH2DsSPV
K/QcGv7aF5Gy62cIKzH5wZvWJfONmK0RyJEPg825jiU7zD1k4xXdFi4kkY2uib49
fsfaWinIkuq752pqM8ZbLvtiwhe1wJnDO+26vD++rpuVQd800aMqZmzoWxWLl+i0
0lPsFbPMYCRJLXFpzdx3x6GCbRG0PGHRY3AoMJGub9X8u23mgaV6Wd88CnyVuxV2
eE9Esq1TPNbJxcUMGAQml695JoZx6gElajj9zBxAdiLknA9uEJxuKxwUHwKNidEy
dFarvuJs00himnvJl7tGveDQhQbFugA57oKaJ460SzR9IluBjmtOdPrrikj+VVo5
Cf7WheGSK3DDg0M1CLXq5Kwq5KOL4qALXM7e1bdOZjVapripGsi+ar5p2HsQDq/g
peXmNXDahYm5ua4kku88dHCT8cj/DS41IkG7skKIDBcWqfz9nG7kBgJE60djwxRd
l/X3kmy8DA+U6zWMMH77gpBojldv8tgl4uQpFu7AQn6zB7ditG5zvr32GnEd3SgF
t/optD8TMou+sgKzgswEQprghxu4D3J9KOpqu2n7/wROCOjWneMx45fgvmL3Xf02
Tt630WAubpAe/KEGf/SudJCZFn1A84eyOuRy0ISRvE2w0gsTR9mCGMREBw3xLAum
7rpZIUHN8m00XjU2rCnURW+V1Hxm+v9+hBeOD96vUoJNRjPyd59sQ9OvKAbbz4Hx
sfe9OShJpAFLmJ+f3mz5/b+CjDO21WJVtUxS/NzfGhoEjoZ644FNaXZUR1oir0az
PP/mPD9Oxqkc6RJjy7a6tk2kZCHKmIQmnmrdKYvDMmi9UwYNgAPCgK2hTJcfOviS
Gx4fC/AaAE9EFiDlFIEjDSZ/Ab/d7+1/Clw2cpcwfYeVzQ/Vn4fsI8bBqQmDJKFj
L2A/vpCC2uBjJg7MXMkYfLJgSvHhXyxEw/MSfYGDQxeZmSH0Bi/j9q2zsZ5Fd8xm
BOB+K4f/shrRzhgpqsTNtObkXR9PmRUFanvj6ahhu8yIwturYm65+GACqOdi6Jy4
oRxCrb0tTNaAOYt/lugh4fTIeuIb0okyNwplFKs0iNj0SLh1/lpsp5yaIpewtNkV
LR/lK6+ATZmuDQGyTu7AJSWH8XIAVx4/sHWnXYja449MymINWjn30E0xNU0xHlXv
d00C3LbClBW/UjPwIZcXaEqhEk6Xf0+D6yrF/DcYycwOiF61lTjoRQckvoqfCGR2
d+v+ERwcfL/IrC+1SqZuY1m190e4ZuKJAN8FXyXzn7tTLfwsDteDiX1LqgdgRvhV
7IPljJrTB2CRSTYugdXS73/2dhT/OaHsRxkVIW/67zzGzqofqmw8f8YDS/1e+wyJ
7EbtQR0WJCUxM9nhxaWLwd6pO0ZgrFRhMQi3VYH62NZ+QNAZx/56+IwECofxvbka
uBnlaV1NzFVTz6HL5JnL4/bnDepFwy2ua0j8zMH5XKW81UX15EFUUSZKqc/9y+x0
i47rttz4vCim92lGcOA4Cw5c2ivqu6SCc+UeQv66WEt96wqgTzZRDquX9vTxUSDC
GHDeTCoNEV93hVzUZNKm5Spnmngya8u3hWtKblP76WxuOC2B0bfD91FED/sZhyUQ
5kQuGKkrzL8NB+0lu3ZIlEYA1THwOrb7iDwseQnI4BDz9JgHFf3g0JVZucGgfvBh
wFYviTN7e4kvS2RxqGJYXa1ld3I6Ad5BwuK3eJmtzkjwNRklOGogvb2OpBb8We+7
NVfTID30uPNB2ywAvKt3HjjH1r7MFl3+yqxz+vGBzQgUrPg1iEMrtH42/wCYkRtB
cdR1rOsPKLCAXQED1KW6ovGKVkkB30BKHKym6MlRAYgvvbmc0PPDRXUAg1KHeOSG
3z+yl2ciztJHyiTu9SZtJvyAXgNDAyId9e/FmUA2qiBMF8yiOxYfTVTKTP8sijd9
dnWTZlsYxBmq6MER5UINVGVtVAEPaW+iXyhbLTcH/4jjRhmMh3FMgibsxDqCgBty
8ikKuzzuTS3tHlfl+f5mpqJJhh7OXI/nDpykT2ljqkj093ZyHNnRE52UHJvOQrnI
flBMcfkdjB+gSwONu9CzTH6J14aXV3LkwI7E9X3Mh1uMn5CcMgCWE75e92lr3lAl
Rp+qXTgmVTkAeOKcYscJ6ag5CkUa7sAWO6fafLqKWbtks2FLAcWhY6PIixHgxN5u
Nw2OlAUoik+GOJ6Ju6h7IEzBc9YOfJnMThnTACTFSIQAFy1441V3CqEL+8KApigs
5Kdu5LLpDAcIIBLSjz61h0SLfN87lgPoa8h7kOF0rKuOcgorB6IrQ1bqEQ/rxZD3
SsMiRK0Lp5JxZVNgfVkTH6PxPRdd4O6KK08hS+/3FStksqqM95PvdYuQgDJ72vbK
qZZ8eBQs8ZBZwLqNrQZn8fxlCu3H4R8s//LfSTsl+5PUDuYFKNq0vCp8DoP1vMxX
PZZdfeEIlBkV6wToZ6bFBRn58LRUfZU281JRzngnPWmohE2Gswpy5Rrz7NmyeN6v
o0YT5LBxHk7y1oqlFsFEKFJw/Qh4TAN4wLAWSSQqob+dNHvX3UXsL1l6T1At+bFT
2e5Dj2zXqTJbxzRsybaNUpA4W+Ha0jaqlExWoz14UZjgNN4WYj4aqZkRUjdPSP09
7qpOx/FreoZzNiTpsCL+FIToaTmItGyqqIT2pXjrt9w+eWYrZIT4Tt0fwm/kVNcM
Xk0LNu2Iq2vkSdQzkFVXpnoT3hQcSSFs8Kr6MFW+Ixz/lFRu1Z0LgxBnA96y+eXa
mzqZLkkNT4EvdFRWPH0cpsGswZ0z6uOEXbXrfjN+e7SP+GXbbahpHaiVc58/wyr6
3+FcgYQDjixTNOi4X/xrKZ8wp0yn4Uu1nCj+L+bgfYUWuje3X67PG8U5ve/gvak4
xwYRnEFzgZMq2uQjMpliuwKvfrxLj1yAgt929Ce+PCMa9NMIYfmTyA5z3lB7dcx2
j09ZRmJkdDi41RafnOxUjuzLTZjLVPgXNPgnuL87IGkUi3KloVlCThlK+H1+YP2O
v7iVx0147h/4YfZrm6rrPeG1RBkvZLHga2M4szqPTJCzftWySePU7eAeQfgCfMlG
h18sSUewkw5SP0TlcPfiaFuYTCR6/71nha43uf6KY2zgNeQJDaItuRDzATWZrsl1
lgQj6MCnQwDRIB3mKia+CfqcvtILyIrw9E4+0Ji1bcqJnYUqBN/RJ2iSYiZ9BYE1
eN8v5yy3cRYtClCai2FkIpUVuRrnWlC3Yx3IRz2PE3KqJD226hVVEqjv/N/Ddhna
baD3S2Kk/ugGVgYJHmALJyFFek3ZWt0Yv8kyvmApl+q36CghlEtTtaKQbUlcynLK
uyQ4+BOc22UKruKv9z4IpX7vNi7FO8q8JTHu29AqOcWhfWuFpf3WCtiQt5ChpvKk
mHQF7jZTcDswPPKvXZ/vzMeF//Ccv5OcpOviKGRadmhY9VHE0rHxfZFLuTFtmT00
BPDyc42cFkauKf7P0YgAez1ZABpDb32SpS5p6X/VzanLNAbptheCMGystbJ/uHRb
FGPdL60sqVS4SEePjQN1SJra0Ma97E7oRsZ7+6V3w9XyKfrkh1tmwGun631t91ry
3JKHtlvgIPXy3sRRB9km9BIgqa8F4Kp+FJheRARCY7FbtGgsxJ7G7d5sqKvZ7eq/
zV+p/2NicWjSZ/cawKtLrtXsQWedRXMVvKHpdWId5pHdS/elvdaWTMzIKKChcqK7
2gxBAIunVKE4qVaV3PCGi+17R4A5zvSnHUwKMhVU/miI9Z3HpniOIyh3x02PfQ7p
f9QPVLeWFAW1OR6NycklhFVlyx6k/D1LKGHUcrpd5DfwSg4DXU9fFgG0l8dtbHoI
NXo4wEXpvo2fQmOFsT9Z7PistJeQbCPhdF3tdig0bwEmui85Y9mZRGmKIVtxaOtN
KTssZb6j5EGDZyRn4CWkYmXrte5medjxgJPkwbnxu9YwwaM3WvGQdvmuMcpxnI38
nIz24ENJLsnKyzAeNNMitx/r2Wu46hA2OmxgR9/A8YaWr9o1tBh02Skw0hzbIrjA
w7vpttLrV7jGlYQgO1fGNeYRKymRVYIIz0jXSdw6i9711DkjAkWYU41byBqgcJy0
96Xtdgf3jGeXhSJM9A1OXrhtjhagtZMjgYk+BGQVr0W6ZLB0TDJ5J1/RjjIFZn4c
iXzFOOSQ9ZMzCW8MEo6IcJ4y4puZpgk5PEdPGRsWpso7eDzqNuHrsxngX3MYjOQU
YCKzsC3zNc94sGji7utPt/PMgPjV4oagxpUFuzgwkUJVbiLmBQJ0Nn/XO0Gmv2Ko
AZVIZRfRtIk2MBliRENtr67UZpbOrXn7oYWYpf2n2REInM+pCJJgRlFE99tmXYcp
c614nCXW7BMzdcIZTD2KZNWepLwV7UsWmEenx2qGHLWyoyRM1+yngpQV87y4mS+9
vdOlDBq175o/5xJzQ8H0YrRn3bauy5XGihP7qTDbtMSgObVIa/MV/9bO71mCSZpf
lzd4MKj6mQn9dITwN7T608gBWzz3A5Pd0XIn3zy0qiXYi3npQSU7MEk+dgELTjzW
D7106DAds62BrFVxmU1JmJsnFGk4MXEtMfy4zZxzg2OEw1Q/3/AZA+hL3KS35P8/
OogfRH6dPGbXMW0LlrNATrnTBYlPgWhD6WSw8vFgBdHd3fJBr9hxzLxJX9yqDzSZ
hITWWYe2kckc2u1exkElRHx61aOpqpTJiCR/xsGt1rcxyNzKOP+PPdBlauvrUiW7
O6pVTbZcMk1preYBjQ1I8z+XQbcyiyDG4NkoKIq73H7cBxYsBeRJeA0GYSSDgoyU
IH3J+TvrWR9j02B3gH9GBSKxRn7T/8I7NCqdppCq55AYcaSMA5v7swj6tmRef24t
MmHYW8ACnCV1vMPNeS3eum2DPaMMH+u27FeIm8B40rU3n+uJ7+DF0JRMRCMRV+Bs
E5/Qq0NyOOyrlgG27ZLDR6ifjEcXNr42NpddvPxW8CiT473mibsqevx+ImJsZhdg
FcWEytZKAFHc4RU05DCoZ+IA9Dq/J8LQv16PYZy5aGG8dIB3HldIrlxQCiypzY9h
Je2BRQmbjb1QWLKXYN/syUsljCvxBTsfCMh17RVXI0276Hb19WYzkagWYXNN+IyR
QlXeNBs+pOHN0pSWvk2i9xxHdyUe8bXZvK59ioRfqmHTb57PHrQn8OmiDwgG7xp+
Es5OoJsb0yH+A0wWdF6+xrpKUkZHLVIyPKlo/GPsTRrvGluSw3OOej7rNToM+FS3
Kv4hWb4H5RHqCp7j1yqIu9ROhfFtBi/izyVPZEfAg4IB9J0W2dy7+tiR9aRnrC/D
DjoMx1AFIsL/UOZzZKp0SIqCjZ1oOOWXfsqf7ChEIF3PdW3wPVn7+LPVpbtoQxiM
H4WbbLjRMSoB4dN72iPk0aC1i7xOTj5kJCZaw0ooGwQ2McAcTGQ79QavNpW6pMwH
8WYI/Qmdo7OSoPlOM5UPCaNlby47qaKVRxWs8E0qdWFgSU68C14ueiLcHPWMKK5m
87hUid1Ygj0rNaCSV91tWALj/LDws9bgyNVb6e7SLyuIz4iu+afjX1x0XdP0VeKD
epTqQQWZTz5fMKmxZpkua62J+K2H+lbyq9vAgctQQ+ijkSHhS/9n6l/LHaPfluPD
4W/hAKQu4D8VjkJlqh7PLau54kNft5Pdz2ilGhSz/+GCnAIvWsXmlz9GmzBg2Tl9
1LL2Re4tZkjijClzXHB3ZXpGu+tXrhGTI9t3MRNSU/H9M3me+HtY0EPLFdT8Wu66
LVauTdmeJTfWcu46Y+Zg5j8cB81fld5BvPLaTtGqHKMTHhcMHzURcWJJlawGW0h3
eBbuWMRDwdfbdkFBHfVWCtO0OZHhrIJxPDuAFCsUF3dfJ1nZso6e4idOiHntAQt6
lxXy8AtK/JMnMGZhfWNmMSpAldUaZjJE4/U0Vyt/ffv92D4lPMCvhCpmnbnMqkf+
5JCLQ0m/KDz8FJwC+fnKiv6ve5+OUviFoOtYTqUYMiMeWBVmoI23Pz/ST7MwczMF
scXrvI0wdgpnZi+Yy+48ridP/T6hp96EignpzdYnpSVphQZK90o0O+YU9Qzbs+wp
K7uct7e0oxlm5rQcKX1pwOLyUx2ioZ2z6aunI31ogV305/FChecJhfjPaZLaklsj
Q0TsJiL2iUpdILDPdUHu1JmRxlfexhRbICEfxPjB+AGDW1as7EUT2aFbionji47J
WhEu4BYZLD24ZVfGJiwn6F9sQfwWiSqgF/uSjUh0NbLbh8fKUb+9yYKoaxw7IE9l
hXtiaEEn3V91PfQRSJo3f4dxNQo3RDvd79jkIEzfTS47un3dvztg3RAHqaa7weAZ
ZMl8nNQiSeEbFv7nIb0dZLBQVKPjA1539sfwbNdIADCGiC1pdi6CJSCOI8dJvYYp
k+h3f6S3mI6WDTqa+KZT1DCB2suKXwC7KCaN2aqgFN8nzKWETGuYBK1p4bJ4OH4R
hZnY+L3FZW/Q3XzAjmt/kg6UtXOWn1x0qPPZ0HrLT2Egq2DU0q4dm9sbkpJaI+xn
Z/tWJU4Tw8mpVhaVXo6Kc042KPMIp2voxi8YjG/JlrOahgb4nlwnjZWWSjcWM+/w
Z2fHWelIHAD4aYpx1FY7L7DPkaQywCpCeHzjcghel9M9XzQTurK5d/ORKt6w04NV
6ozsDgtykxW0OqsLLn7DCeCej4ub85+Btwxh8sYrFi7/dv0wKpjlg+Xb9YPmUH68
W52zHpzE5m61Jp0W7G1kyFp5XumKdgj8wqoR4hItIK+IdsxHibkhN0T87R5zUXYe
11ciYcZwRAaOqP6tyh6TBTxMXvIrIq7kqCP35J4wxXKidUd4Eku0o/6lvUObwzXq
2wNjVnKmgFqKDWsJt5VM5gCZZEwBoymD8OQBT0EiDvaJP3vR3pHub8cDWgkwsbot
sqNJxxZZAggKVyI7EyOg3pPkr1Cu/zV17Eijv9DtEVQIkV4NyCtFVEpl6c8RKUcI
3kWU0l6aQhxGcYw3IUt1IBM31Kr258yRQjUR3PSN+9hf8gsNKSeEKDXI7LmCCQFH
2JPnYPEKl0JtLwXYO9WS43L1A0FGpoGnwRamlvqCL3qFhCxTY4GR8PCmUvQXJdR9
evkPFn9bDQXy5VUcUS4hdnna4dbE/uS5f3DCy718CeM+KRUEUzXRjw3tgv7l6hY2
H7jg6FID92WIn4MPuE4aOgrC/uHIsn8bG0scM7kmsNFXp5yGc9+l6lvbV+DsIPvl
m0Xb0AEP9TE5I38ylvA+b3BTZ/xx1/Sr3fdG1i7SvIE29xZIUxLeqDGw0bybdIUj
pext9RtvWjIbSRmKKQi1ocLgxv0Bi9VtXAHVDoxR/KzISt4Ds6tce286tAOsSnQw
qAVLENKqyfx86TSzeACrtAhXbmZBaVEu0HoW98HeTaclZeIxTM/OeVzLMMiGlIyx
/b6Gv23JF/dXXlnf5Abmo+/8Ksxo0qS8g5oneQuuUpaApZMSqMla8HqE19TkEV8s
RGvtxqfSm6jc03ESQtBlltkHki1xEyelF6K2cFSB56+1sbAIhR4l7J1ZkxPCwciQ
JzzhWCwikDx+HKrO0h35yAE4YHhWg0r00uONpxKpnb0IkQrVny6ovaQtpepTsE4z
lRiUFLWzHnIyXuejT2QApZvTw8x7+7xqIsPP2i9cLY+3TvZiS4Kb4+bHUz8xiM6G
/GLDwliwcYef1u/z97Q+QpMZBQO0gKYBZwNW0xYdyl6UZ1jtqiUQDl24ufQaJPgh
ZPX7TeEj3kWeSP4N0XYKc+v2yBlpLv/YvQdgBe+TR1w6gulECBk7cFQmN4EO49pm
4DtQ5/uZJ/SSI008Yo0rKEWJ8HpZxIAMDR3QPkZUzOMgCZJqCfWVH5P1CZGtaSeF
/266Mx45XSSq2M/5vtrLFQFEhQshUH7dlPUvw+uJjfJi8AzMSEuJIzEZG0gU/1kY
OKRAEpJWqY2H70sduB6SLae7uniiC8RRQqpb4trETnKN9rnPVKHOGOKIwr8PzMza
FK1MLdF/b0+7D+fr4bN6pgoyzspzHZnjiQyxFP/dAzahfQ/VW3Ae5dIVOFECDBkR
KtUAZLLXpSKdoUvCRCBe4OxBqrCHQRNvrY5LtoayNe1tJFPdxK9eH41ot4J/QZtt
j2mOGQK93Egz7uxceUN62IX3Hs/H32m6QZHwkjBLeqJYqhCIY+I6jLNX+vpTynQT
HzF1ffPiXSos886jDm+ic2P1QXDKxMMy0rO8FFby3FziU2B0OGQ01GT2jQcqI0T5
zQehFATuAQdbS0weYPW2C4nsdO8DIsLFS71UXGzUmfAQoRPdx5RldHG53b2Iy1vD
tHziWRiilzQSeevIDVTKCjYHw+SFoC2PAKTH3cQjq8RdyqTUA2Ys3Ii+aJOndTyG
Vw9RmeeSsZIn5enxSWNko9358r9bATfUEhhlDYVm3bmr+vfO1ZNw/fmFuIzbYnAK
9i0DrDG4LzjvbtMGaWLvl5aC4jbbIvhE/4ZzOYb+EJt4CfwpwyX06TgKU1zwUlVp
bf/lp2d61jPArF3uVbd4KpftFAugL7L1Yct5yFZdJsfgwm5QbENpT4FRq7qBoUaE
oHX1+l0WTxusfDfiMWV6Jymqj6Feh4QYBbgTwpKg8anTiXxG9fFe0Hby2BUeD1jb
VCntZ2T8Mq7Kn675SyU5Ug2tzZB298htzIKMeV3heXxeY0xuQaWDa1CAEN8KTAOO
mpm86gfZ/arOarCQFDK4ZdwKF7GuXkkRCTugu3dWvVc7KDI+LVnMYdm9b5Je9a+B
7Dhi+cfteSomoGcPW2CmoaVlYjIY1Fh8O8rDQlCb9D6yY459XBLm8wbmfnR5TbLS
Fi8GSD5smCb9cDvsGBnPDTE80FEzTycppC4XrE0DcjxvYYZV3sLYzZ02l7ZwVGYS
EbH9aLMSe18uxQlBUHQnZkUq9q1eZTubDyxQ14yZILZ5sA7K7hyKfkAC/EiqxoMR
Tap46EAhGvay6BfnPzRKT/bTT8kImJWsYirZM61kuO3qGpcdb8U6ybKG2yry7m6/
7rA7GKYuHFU0hUhTxAM/Zl6u/3t+Ep249bsnWUsH1f4vCho1XNmZjt3GSiboYojq
e4W9kXwLlWBDzt8OEx0Tt4cTkYEuJvpaupOx5U2/EAMN3oE/PlwUwRoAZ1ccopHN
NIbhHhrJ4HGlOURnF1NOBiTeMvhZ7z4RqOAfYKWTYrc0+5SUgfxEMNqF5DjSkTwo
+N+uE27KEvdlBL50J1VLbbSldUFzNGQKlllVj/1c2YzLzu+sNkEmRUfk2Y/X1MBi
lA3rHUetijzQXcWIGennlNGeL390nO5JJUQIkzZLgnJXI4fKvV4Esg17hG5+fNft
PvzKP0t5u2/Jx7pjJQw+iJ+Ybzj+qZDGSI3i4ESG2vMQstYa2orRG6KT6n9V5sri
15Tgwjep9TZ2Y6Pg5sbfw6C/yOHG6aDrfgAMWh/B7/7w0nw6nD0TvbuG9pEZ8Fhz
M6XfnVleGhZnOdyGzpFQ84DE2GWVgfRFTl6HptxeHhSEQG/wVXhLFKACGyxE57Z7
iGiTHW5kNuSGYkLPY1GFfGb5y/Dpjjc2QmKWnigD2Wi2rmNW5zhBTQQ/hwpKEeur
eYe9HtwOpyZZSXtGesC5YLzwLW0nUw0dTLB4ZbTfV6Nq2AFgF4QfevHQa8tTP9vf
DvMIdMTQRnbeoxCAqEyTGW7x9TexqHm5Gf9M1TUuuetD0UVeeG+En9z2fy+Stqu7
P+t1rZtxqk1Efyq2agvoy1IBolT6iUmptvcL8eNNhPAcDwbHrr4SIbrfTdJHQF3D
YPu42bqSOy6InhQgAcvZxIhwYsDM3nTdI4KanwK0iFx+WIkVl3XqUxi3yYc1ixAE
ssj9C1nRlULQCcYOPSAviX6ju2SKEoy7bJ3GvXzEeA3QQNEFqqbxEq7DgOXH7Kb6
FiGG5Nf1ouK3muheOytIXO7hD2XvUSMQrhSsUNKF3f7oP14UimLGfPOk8UWa4xdx
aAuE6P/hxlo0Cy1KGjSjoUKvdk/0F3LMtPdUOy0XDHMJVUOABkmU8FGmYyXODnSw
cJ1XFhBZaut2R4pA9scClZnbCtjMPi9ESwwD2ywd2QKoVLFWP2ICL5gkHZLL0h0Y
vgeeuu0Q2dk12V/kcY+VhVBPvAfk9IXJaRhGTtlJ83kDzolapHMMlwWXQAs1m8ed
oYEq4IMHkEjZZZaPGRH7/5Pwlb/FUSZiz0P4ZKD3aUkr4hcGxIq50Rdj0rHkfwOE
ZDpomuNKTw24k5GTc2EX/hMQOHMcU0dm0aFEyGRrvPZZsJu2BR7bI75I+rAE3f/z
iL9y1AKOmO/O1X29PnFV0Y4PC7WzYfBUybVZgTNrpm49u0j6Q/5TfCVm7BCoxWJK
TwcMNeFypgDgv/LoJ6i+Sn1pf2zinb79bqYmeEQweQelrBfX+S7CPjs12IzX4EYr
4BWLItFW6m87hmvaKQ62VvZ/8OeqHs+BmMtfpOY7ia74be3iJKitFYRzGTn60Iyu
/1pvAObLEQY3tqtVlYhNx+d0175tKGrXlVcTQXYeDs0VgrbE0slgv/6lqLPiNyDd
r2z8Uk3PmDaPltT5GLdeIttlPZzYRXnYpn9Q5hanFrwj8DqJnhXWNWWv2maYguF6
X+7r8/iaBa2MaYOZKf1ZvDMVd+gEQos4JQj+TCu/Elr7G6FPkYCFf1zfTd4wwfi4
EvI3Y+s/9ZkEhTd/qYjWOldtJFJFJRVuokoCk8MhhlVfGvQwtSv/bnHAP8zDk1ZP
ipcddYrk2eCj7PXJFiz/r7F8xPbC0exeNJgAkYds1bNp0UHd3BdPRR8ocjmy3TmJ
KTOmxK/pRnE1S2vwLjiBZtyJ4f2bwGsq6eVsX7zP9QjlyBzq4YReLbAPAvnZzDBl
rpPhYP9/lUc5jPyEjB8PhYKwbqHJ3wLpcmwFsQxxcJCjUCANVkRKkHiChbeO5rto
9ufq0r73GldAbFK+wtNpea/Sqxix8cv5wcE3r0xiFf5pqZz9E3eqHHcwtrAB9R7s
CYHyM28S8P0myNV1FKIRM4CNJC+0DwHkLwqTgxZ5TdR/yzn9o3JyZQlbpgTomzpd
E/tjlMPd/HeS8+7lMKtvb2klAwHi0d+Ce2XWH6B8ZFyuOlN9wrDF/e8V39VWLpRR
Ia+yZ4d70jm92CQ1YQBeEHg8W70VEmtheYCeDJtFC5Nqa8ZejJh3o2ylaPsuDyel
oCgHUdRFmHFazOdo+LWSlgpO7ufa2z3jd/Qp2a0O1hngh0KStp8rt38KddTSv0IY
XKFETGftQYGIp9YVTl9guoLz7V+XEM7ndb8WMtNtrlwfrjMPMevPD1XVP64b7NUC
B9/ShfxtmU/6cvE2MxKlL3LFlcJ8z1Xm8FbKrHzT56BH2ZXvwgmuY/Wc07nltI7f
XA4aOldQjzMQ/qPYgE6Vn1mtrhiLOPo6ocE3y/HOiRc0yfYJ8XaOCatI1OAKZ8wc
SuXBgRKlUAMTMScroNzQVtWoVuhlXc1xtJNQWJT9RfsY+gD98TamvJ4NiEykNspo
7Og+ZPeS93WqHljMxcN5gK4Wyh1/aUeHslTuFfm7WjX23wAn7Cp/RXO8plUPsAu1
G96GSvjLvGtTQqV08DuGSLCRTlslm+fur887osEwdigtmgYGKCdGY42wnUHE3qCz
fzhVsEGo/zs/M4cLniVUR5i6juwPHN16foJjN8qoMtLQlhERBBgXBMemfaeWNnup
FWLcXMNhp/gJvT84t1lapM5dKHWJ+K8qH16OGvLnon/nBDqjGQHOB2W50uBJ5/JY
ZR4ZwgX+lRxcbiLOea/6VQz3D3yH/T5VDWtYS/Nr00smeGhmPULVudrQlUHiGcbD
PUW2d7jLQC+HdDBrkU9cX7rxPo69MnNwq6a3Tb6sUwxYt19tbY/DPyPcLUnYigyi
xBLJi77G2AVTWjFylRqVj7G2tsZ7QNwup6oUpk2uJIdB/rd/vZKNevCtdc51y6q0
Bnl45dlCMnrMShkRO7u4iAxllnlpSb6Ls3OnLBoDR6FG+aM8hzCX57aQ/l7lh0m2
LlPhWV5sqpZx0sisUwKKjZBSvoCktDT6mdp/tJ2RSPT2drdk7v9g2iJFcJkHf7ZD
jPbCmStONBEV9xtvnCvdjQqBH/4n8TL9nEf5Nv2jntPC1W7/bJdbadSLwKnylCo3
aB3UQ1Sg16rcsoPgUQqmP+6sKf1FA2k+lHRNf9mDMSbauxjUn4CGgSyQPabyZZb6
Ej5PV9XZwG05hb2Dymq6g1TNG7+A2I5i1i4o7z+xLPuoWPWptE0tA3gzGn3mgTuA
kQaV3Ef/NOfvc9os3An+IrMbKASfOC1WwVHQB70skl09POx4znfpCMdjgpGxCle1
O9WT/Gc0T5JqRDZmsMdpsh37XXF1rnPe9tnqXRdLwrkXotDW4x7fAplEPAAzA1HW
OTYSbwwwXBSJyV2elgF/B+P/EKiqXhp34LYKR9jZXBye1zvI6uqm1QwG2JCMG61a
At1/OrT/lfFvSluUoiQZCUFQuRc6ev8CRh7Sv8B5SSyCUs27w28j4jR1bIcRgVdS
ykM3KzQoMwk+MO7R9k2ur9vYC9DOuRnM5X+xlVddue8b7XrxB/YkYLWV1l7gVEEI
lWh2z2rYeDdhar4QdTWCYpuAlzdeaypdrKb+9RcW2EmjpmAXXS8XCph1t10J9epi
zc0WfyG2JTwO9zo0PX7FL907EQkCkLCYCqEV788H5BdT0wKOT4uIccXu0hn2PP0I
j9EhPn0h74YWjaK6AClM2p4dUNvcEdjhDiM/mvO29LLEopB1FzHKj4idHxmrXD6c
9HZIwoPwcN7Qtbd6ooKG+j3+ypur/7t9+y7/JweeYMGkKa+QCHrvbaJpCLlF1Xuo
9PeA/EP4OTr3j0RsJ9lUq8mvD4lt1pwJncsUPFW5/A7B2WmrXqj+xdmrZGbxZwjq
iiXC42Zjd8rn9bVFGjpjY3pYkPdtkjv9g3nhzx97uPIAhyOmcGnrqUPxWKojQhW7
3snFSR5MyUygw9cz5OOC9uukmsek6ronEISSaTZIkC46zQIcoa17VBAl4kp3Gngu
PyHqWvHbVldIJ3qiCNHm8QFZA4PqSsvM4mYB0RE9i4ptjOihRu1qvWl05X4PwJVT
kgVegnwvj7aUUYAJjf+MrwVG8WDSagmqfXEFNqWJN7vXzTH29GsRhXpY1JU+okzT
Ph0rFzeifsXk6iL9L7uJN9UrJ4NchpQJUFKv+nNHSb3j8HOpNk0dVdQhVhyt/zMN
yA3yDOkF65fwNsMOD6Z1XkXQOJl8Jtbc6ZUy1mWlESAX5s3aIsbH0WWwDsc1aLs8
RfsjQTligt32aJevAfoPP0Nzs+A8HJT+wAkQvQDSxhs7Sn/RhBWbAAOoq2h3VSpw
aUwo0frvyyS3gOBdPmvR3noYk1317DeB5L5WeyYVHVU8U9GzR4uezy08XbboGYy7
XGTdkDpGWy+Y3y4WTfc2rDn4Ihu60jNEC/BUXqHlNpISCywMj4lJHa71URwUjZMc
KMtMtjyKi2cEEsKFJVhYybsLFCFl3eWhSbF319UrRkWh8eNFry6esnLytUAjMvHY
4mZec6/7bcYuVt89EI+p20dyfiOBixtj+amGaB26hA0FJ0it3khyPu5YywAL5IG3
nsmLP01naHnbArkPt9uBIqEh/GFT4KTfSSTKiM4RNwS/XRO73bGpGn0wmu2RhR3w
b+Io6cKX9U9MKDFZuujBMhWMtcv6srfZUiEkV1DmnfqtW9eGvC/0fAGUTDCZrsSw
AccTjd3XyKhE2vsel3S/FMDJr4FUiBOuC1fbch4SH/n8jKcEDmR2J+GqxHtA7S1N
49sRsQcpW7wo/ATbXdW6IyUvqs4ZfKV1qd2DbnJqlTbn5JBTmeK2aRWFe+B/oXkL
K/aDgztJu3KetHL1Se/DY5DMjLM5AkL1wbhsfjKD35I6rZg9AkgLCi4RxAfElUNq
ak2rWWc+/R2N5H+zB66tOoU1zigkGFAYzUHy/M/AeGAIvCI1BcXkd8bfNWrCjWZQ
guG0iPvHv/9tdUaXH1sQyMJ6TdN3vjDm5/RTVGYZLtu1K/IUrG4E8pKP9TR8jCHw
qMifI1mo8OQJ4rfQujMDtL/xWcWqfrILljRsCttEyfAiY9g0DCc9B9fHaMvcm6JC
sXq8ADyNXfaVg5LhPT3qJfretYrLwGMB4ycwJhkPl81HoQ9m9qGCsNz/dnWB3+jx
xMOxecyTczvwwwPN+9OhqhIOmWpJxlR9rsFEkHxks1dbk0GO7DjP/wyW66uBh7In
j1fyKZzVouRz98ZTtXrBzwuhzDK1s+SeCJUuat3PyaFxZ/AO6fVpXTl8/yOkqk1N
g3cejYdfXVrV0LCug3O/1Ul6hPOX+21mNXBASZb4j5a1EehuD58VjTzzCpPkt3Yi
LKky4McAuFUq2KrBIhonmVB+9f6UwSb53v0FHwQceHRKPvYO3zNUeALgZXuC1mgG
zC5U/vT+Q0My8pshJi25bkQz6TFy9F2jCW3oHv0wRupRcHr6bdWS/ePRubXOyvf0
HUNhv9rRP0Rbeua0jVHmkNXnjvaWPsgzmZju6xAU8IYccYwzrm9bvJ/0/Xc3cldJ
SFlUc6HNj4GvPZtdCjj/VpSHp+iKUtUGwRVV4GCUsOI+e2b1cDxBZUQYD24iA4L2
n/ualuwyWWVvFHRm2d/bfqWkLL0U0+vbSTapmCQQx8+8lWMJ2fH7l756mItbogXs
oxPIr9xS7A0m7UoqjVRRPasfh6TzABcQh4VM6/qDRmxZ6rysQPJmbyGhN0xEvgG5
UUzGJCefUFAkAcXpgSz54kzpvXj1TVj0vyiKN5LYQGoeJEIXTw2/lKr9zmcQhHPX
Mz27UNVRksz+cHorjT/DQ48RD3wYaUPEWxL2Ec7DtMBMwjezldXRbalwuNSeWOAe
kjPtK/plOA/Q+XJTFC6qGaU0FBdHDpvSCE9p40NKLd7mrYzXld26Y3cHKuzioZxq
pMjGrDzSyYRZqabU5L7pDudXpgBmPByGL2/nnqRTl1Zq4vZvwpTKsDINXkAmNxHm
E+Bm6V3nnSC+Zm0UZIdnA2p682GyjL4piySuNM3tS/spwiRehXws34skxlUXg6iT
N+tA4mPXDwO/t9WtbvUiT/jDjERzVIkssGP2VyYnS0dCUHiY6aFqUreAnQwvZBPA
AZfrGJP35byV5GQ0tDFqZcPq1Ol0Vp0X9l57pWDENqrPyNmwPLgejnUMboTFjadd
P2qeKPLcrWY50ppT8W+EmpWdaYHE2nzhOk8DHeL/glVOhzDadWToT1wqK0Ta+zM2
VPHHJFNfBnJug7s0DfNo3rwzgdTcvWffDYBwLxv8pl9TThz9jkMlQZe83nXqvdBn
iEaOg24a7CZgTE4pU+/RMj4Zc8kw7B1yPIgsRqGi9g55OGQDniiAAhukN5/ce3Bc
bJyykjigkU7F3SPz41NSMsOF7Y7KtR0AqiRQw7eg9JMabx0LFvRuju6bylqmtlSD
0djL/tBC0D1cDcNOBSJY7kXlcwi8a5W3YLy2qaj1Pf+l/Z/S5YQEqpbM6BHJPR8X
8pXil9o/Q1YvHw7owKHVHeJf1VoesJ8bn5YelmyE4teoQNKUcWHekqlcUTylzn88
tqAhamAQt87+dcnD45tkqirrG+s4xXgy6D/LZaDFxbzLO5wbnGMbFeYBkXdNxbdh
5IF6DYKEFPDAEiCSgZ7nlz93Mi+lhNRHcWSvQECuGXWEVex58+D2jBAabgI3F/0U
0wJBwNzVT0bqZBM1pZU3cQeirxqKnbAp3vNX+oeYEI/UpcF4ZWT74A+FvLHaZXuS
TFkcMQOpKvG6ZqO3RSb6+RGqaHOoqUaHzamQZ8lPUjYf4m6kAN45vgvRzQW4Tk3M
uVIkeAmE47JrZxE2VMD8p46hWg7BSiaxbQsNnQJGRc2bhkIgdmk1oI+yrB5b5sBy
zQyc2DRlYnbUmzqxLAtdgJTR/tlzBUubkD4HeNxbGL8hUvzr5MxIoSqcFx+66z3D
n1dd/Gh1GFr8THLM+zHgoU5qLmEspbZgStNn9eba9UNaZch3arjYJrwcwFW3CIOK
9+nElmLdiVgSercyUAKcYa/dcE6VCk6WbuZzOUNpSZ7kUT5iZB3bOfxryI2u8kCh
iTCi9m7cP0hU/Bhav8wfeyjr9IfBpWCZ7kqysEedC628YIckwwRNSvl5LbeSZ51u
tXXm3IGG7mAVep9jC9MEyAlh2Pz3A2B/u15pj/r8kD8AScbJ67DCazGGIobe9MXV
aRtp9wfsChlGNZgIZ+CLt8dyMAqVKtW33QbQfbuFGgeV3scERQ1Elrn5J05WFBDv
yuR5mEhdJ9tnZnpkZnBJjBmNG2wyyvHPQVSN67sPid2fpimoIG7qeshEHyEjfwXs
DXv9/oIBOrwyAm7d8xwCAYYihtPQoxBtMuLJYTfmSXXMnig8xJFXL+ecN4QbpRtb
C+0Dn+UR5195F2JoyCDVuR2C4mputk/lXDrqND5Nh354od9Kxwk9Jv0eRQtbI55M
+7teCpgsVy1UEAafnHANhHFplKZZHP/K0ya8AhPvOgGqo/A0ljhsAOoo47l8+6UK
fbnJ8eaEt6B3FGBz7bD76bZxBhe1Evj/x7WHufZvvCyT/f13Ib8CWcOIyujr8cAV
E4Y56yhTypfVtfs/I1Zjpeg5av/r32do3Ws8ANorp5cns+UwOSedlsTEaOAPOlWq
3OkN7LfleYj4KhxTo+f5EZ/UbPBaLuT+NlkmxZZBM/NsiEO3XqO0CrzC0GYhpxFx
uyxrbqmiiZYMoYhobj1v2N41/Q0yn8P0BG1duirUE9+71x0/5LvWaRx/kvLztZVh
6IEyGeITuEBUvBLtFovRd5zJtL77p1fH5tqEOWpxWUjrnp/+Stz8zDCuWKv/Af/k
kL+OS051ji+oDrOWd0vlnuJzch9FgIxCpubU5tWBrDpCHxrlgRTx9Xrn9Hp0KvWT
FNqluiI5fHah/ZJAxheF8zkGTPWHiPIaUPduKALgQMSNDxlI5XBaUOg5KQ4rztma
R1ox/o/7r3bkGcH5gtZgrccbK1SOvLAiahv+26F7hIwPNb8CQlen08OyKEBKROuB
N5cmAsA6biT/jBvXEAwQ8TRqD1Pd3eE2n0dVGEY7luLza3GXHk6c0kcBnbpJtoOf
vxU4Tl++G7JaGO0Fhtp1Npep3R3EREfk0E6DpoWCn3VJPTvFvvXu+IJPRrbo3STf
XhCTmzmFyWVPmMwUi4moXCxWiD447MJ04iMMsvRp308mLEpFXtbhuiST07UihJ3J
dzV1DliE68LjixcMldaFpLjMvwbzOeIvLWE0tHZlK+SAW8ITP/SgDm/wKu7x++/m
TU8Fgb6+C4My3Y+7rfNfo47Txjd/14R5KP3imZqM+FyymhfKpogLtionsWBqwoRu
h3sWTs+4TNXKRhA5x5A1QsxZmfKgMcItkAEXAtiz1kTCtp4hkP8yzpmL9giIYUH6
iRlYA8l5iWkgc52UK0+nvbnVU/VaHu/NrmP9dEqtYMop3lLgDD/uG7CXx63VbEvW
4XMcGAnyQ/tPZphOW3FlWpu6uz85Lm0OVJ5yw+ZIo5l59JqbJwRX79V3douCWMbH
6tscTNTewsFWfX/m9qm1HZVOQXni1usD0QIz7NUW51r1t6Oi4wcsjbifcFwlpZxp
BwhVQ7BXLXXiA/8UUi+umHT51SLNHzzzxFQfCPXPXo3cHQL9N22bzt2UbMCLYCA0
+RDmJGw2wQOUe1YjC05K7DLNIXVnfMGBpe/FGp4Dhkz2orgaZVToFzS9yrfqhBcl
f/4C6kaO+khXxxE20M1qOqHofW+wTB2o3ikxxJy9/X9uLvJsA821m67qmZTkS7V3
fAHCanb1wieYE9BrLMAQN1xyfMJfYfG4L/ZKZSbDPNtWmRcc6vXDYwlzbarj7kA8
QSZQljMv3AhFhP3k8KH5Xae53SRi8dCYkP6tVHwCx4n6ZGoaN/HUF3KID1+CactT
MNK7a1uMoG/g+1DN8I6jS6g07RWbnlY8oPM2Pj1U/fE6vbGGAcIL6u2bQhu28EYC
JkR8li7h7kpWyPc/wu+sj9F57chymIaIk3n4WW2G2cSbKwq8cKfGn+qLVX61b5do
k4avSPDNTz+Uv6FOpB5xOchIIAmPGzRF5NHMIrGTeLwTzmV1/5yfU/mk5oVpUfJc
xHL9W+Scb/pZ/EbY/PjIfxE/0DUlxgZr7t3idXDSsdSHHdTczfNIbS0NhrDH1R89
4wQ41HUrmUMmdKzStPt980uWoyuNOVUX1H55YDZRmR8RYxp9ngXBCSgMiPYwTMPU
tPzMyfP/+faRyyLrws1X2/AldxL/ii3PP3nb8a+MrFr64ewAfu7vNLjiu9QpOEYj
ET/BuPj8Yu0OgmIz3X19aE0jBhu03aIPrIdT/W4gqw9D1IQ0LUsy/uISkx77CHH8
PR1/xX9XDWxP8PuBIUvRzEcQJzhkJxb/W///HprwLtXcE4yFxPodHvPjPWkbqIMV
p3ej6nIbcUkolv+ZTXZ/I4i/ZDExdxG/jnuKZ8aJkYXzYzWy/5PuiJD4R7Bp2bXE
6EQ/afbPyTTBBjQovVW7iVWzzJ4/5/i7RQ9QavHFnJRJTJl8hAxYdTfDh1UQ2Owk
92BYQtykBVv+YT2YlXPwj1jnjR5yU8Z8C5nrcMOeCtX7GW+krYMVUA/qUVcgqCp4
U1Jcr4cyrZtqbDpmCJwKZrCwi0Elp4wtq+ROUYtDP1uIs5Fug7gEdCRHEa9Ukj5t
2an7IwVC82fTcblH2ab8ht7e9fFqW/SStTn7+GL6cfSlPU754s5dlJurKdbRewM5
4xmxlyUNiVG63Hs/Lkfp6MuxxrKVmWP6psqwEGETYouOyJOfNfcNFJ7PAhJND7La
EPHNfuxCcjdjDXDaTLp0h7UU86R6KK2tDL7/bi1hzfSofHePZ95yBeQZtGycstVx
yBJK0klOMw//2UOJVv8VS4PJtLutw0zzWDffEgmHT0mLHa//2m6rOl/4c2g/VGl0
MJD4uvfww3bODBqHGcRu/EypQmYaaF1/eMSE7ZLZobw/6TseiSfbD2CiLuvqVeym
3CuhA03phFWUTdkoap2P273E3VEzukrhvkbxvCH+o0KkAVJsXXelpeiPiE5YdJmn
9j9w7EKtkuzx7XvnkeZY7J8A6ugvBTCRIVTsHShGf9a7wdMuMoe6m99Xb3DjFBYl
g+43C5tHimeRjB9rqYiPufPw+4sMtuPxRGZqUj/idgioxFCg8FZs6JguqWt7l5Ke
/KEiNDAjzoJu/dut27ZJbSz17zg8uJvDzLRupe9TJzYSP0XZ3gy0T0dd7ugCQzF9
Tba2zOpluerzs3adUwWQQJSO7EGpoemQf1DDsuq0/nGJFl7XcZsbPJUdjO+sgKro
VcmpnS8DrBTx3B8dRbv+glrxRtXB9iWK8kRDBL2tdnMk5p/R9VMDaksQ7rxeUoc3
W1otaBQ+PCPncJGyGhq3udeQwfb+DVdB9UujzfDo0lHyKYj//AqwS4z35w1rU6uO
6xl72S0LRsqe6QmtjJP9kNsMLXaJlCvYA3KyV510KIPjqg+rkUHin91oAnfPXMdd
/dsGZIdqaELywvScXygerP8lvis6zjim2DLlfXcCB7VTM8B0Gh3ChL+3xxmrdH0F
oll+zuQA7TjeJMM5Esi7af6h6COPCeXePM23XAhtZC4siY0yZZtq3C3+UPDRTS2S
lZ37gLniPBV3inZv/nSoZvOMExyT5MyCjSjGvVz0uqZrHRsvkNpcGd9YsLSov3vg
fse1R0H3fP/QGNagRBxXJ9N/M5r5Axe2rio5G8j51GVszuhVCpRf05pCHNC775Hv
Tn1kxj9oWathznC4ibCYV5Rcry4Fn95jdj1hlxrg08QYvJ4xn8BUUgOHYivSNVh2
1JLprr0cWQcmEeayCkbIrXf8Kk21XzHcS8u58YoJXMWnQWYq7VO5de555fS0lmt0
srDUFOZBJPKNFhDXIuCPY6wsyib+MSoqqPSv0Y1dM7CrFOmYULEnrac8xS1Mm2Mo
bqh+fuFOxp5AYi9s813bUA4j44MtVUP3UFCNQWkBlaHi0Wc/UlTu6qTYDnoZGXuu
s3F1OgMhL3hMPDSSKHjBg/ipusd0TR2NE+ZzP9+y6EeHpxGp6pQoXrZLdCwzoiQ3
g93mF3+MYZMmrlY8QKikx47PMfFLeJK31lENosiugQBcqxrpERko+DC7ZxI9QDd+
/ccmPWMmcqC/Bby1GrL+HY9BoIcwltU+EZPkp8LKLiICzsRqW5XjY41KwW8IwKrH
KfqW5R7JKb4/z9C0HMFSAW7woVZjEdwUydXOk3DH9y1L1OvvKMcBlWt0xxiduWGi
p35QM/i5wSxnIcnJVfcc4vPWG7dtAIkAZ/XHFDU4kRVqYQjaMxKKKLkbua6JWGEX
YaccZY7TBqnWmiNGO+uFxf8eWeORiwRojIct7Ga2nNLrJE3Ox9LeX1Aai+uRjfQb
tuJP2mleTtM/n+MTIJ+leb5eErpKGncZ0QUEI3NA/pCp0wfPvNmvEuea3Y4A5pTJ
4WMfhWR//LVUpm+KEQTkbliicrQAZVgpV9cuIqZ+0UP82sceUY7GjEj+962CJB78
DiBkaHk++73KwjPDxa98QDooC0pyk1LXZaM4aek8BKYnQic+zwmAArkMN5R0KccV
KkLczcKXTkfMCcPO5VME+GxhHqDDP2wND03ZxXKgA74/tn4O8roniVVdVZhxZJ4U
Tay998H1JfR7iTU7lP9kFZjAHf5qpT7357vZ98sSJZt8ce9mDsW971YrFTu3i3+X
oogPmcB9IduR+X2O6zSJ7vKF6QNS1PtKXUCzPIovtHRWoBzV+DWRb7U4JRHw4/nb
nxjkU1EU8+sQxPgNhqvrCuw+kMVrWvLTkViK+rDMWweOOI2Unr9Y7tMH0KKC5vyF
C1yXlgq6VQulCivIRyY97VDXuIrCXms2zsL4adI4DFKHukNctFSvjEpSz0WGZlRd
f7K2tgj3FWF0Mxk9Nj+AorZJfcdMkqVz81d9mKWzPl3Th5M0t35d7NAO+eL4wNzP
vK9WGDaY0Pqk13TG/SxvZFeQnmnya7FyYGqWyWuyQ9Dpuu1svLs0XXPS+2Mp2r77
+z7mkWcZy80DfkPKJ08UpSZKhQ7cK1ywczgGObVeoyWqiiMnbzlv9LPUQa9Pyi/+
KeZig0FOH/n+NG+2R0aAmv++I7YGVFx2Au1XSbKvl8/UOCkROKGtHp7wqwz/bRi4
3Px1xRaC0vXOPIaqaLOjqCuO1X4gbDX3c9dd/ukkM4FgIepseeghLq8UoWQIr0ow
UgIc56ofWw7fH4KDzbmRAV7ZSa1YsBFQc3ATFabCpZNkBgxodLi/jECf0betOSg5
B6C0A4oGdDnfnohiKPy7zFTROOrXrszWNjPp/mUspYMxSTGZk1T5BMk6YmIFIm/k
LneQpAowo2b/gsrSqu49VEv/sitIKyRkr9zcC0/qV7/pB+0sqm6OksMhAY7fIcSe
8WDI1GInekZis9ZXDbv1kq9IsRBCR5wb0Bcam1MqJrgusu7ZnTFidL0kVU3Mge4r
SFbuq+zSu9yVOnrDyFSvmHqrhaHW4b8CvzhHGVK9SMS7i0yezpw4ac0Kc4xWdZgi
gqk+YOtsG0vcdgQlvPzGB4NqNGlnazI5yQpKF18up/803+M4akoeBzzvTCHJ8ghk
JhTkwZQltRIqlPgBPD3Jg+DayLQG5WhYkFFJUBpLeMMcJJLDwR7Q409SukYEys0H
4LaBulllW+RrHsOT8uQAhTpvFyu+LC+o97fzZpHlE4uugXCncbgM/IUDwdidZzW7
EDm7+uLsfu9u8PQKYZNvPBrzxraF1y2mDCuHZON7l6hYiVQte9p2bFJF6co5EmZY
Lphwd5WrEIZjtP6pvzr7teVlV6kyIxGxzKmzvnTIrr1R7Db4LjxUyjJx9T4fla6f
4QZ2YZv6gUZd9rVZHbxEBd8JDoPqfHEKQQjlzNMrl8khYHb/uUZxL/nefQH1ToWY
elk7msNCy2pL1PPZaGSKH+R3nv20eEzD5ODp7/9ofP02I33LD4qh+hz5YCYnkuyo
gCu52N4Z6/wAG4TiaMYqPeMJ8e/b5TpHNY8nmP1rU+LLTpLq8kdHumXb91vjwNo1
M8GAG/NsfuEThrSYltJdvftWijQGeYPejkhnwhxNZYpmECZHxs5a4wahQqdEALx/
/HPeU2fF9nyNUhUqtXzb6E5F3E9zrx8F9tsqwApuabST2sJ3o6mo5V6qNW0SpNvT
E+poePP8K9ihy0nmLXzPEGUOHP/b49IwE/XIvFTCybZNc2Lp/43D2LPyDlsDFMhn
dYWjtl46s1gH53wDlt6819gZUJSFcnSDZD7jFluLko/iXw8tmyFnixio56RIM1aE
K9heoWEpRFT+8+W+MyN4AUCouhQvEVADlNAtq4oXMBFkUxDH6DjbvhiBSCY4DGaB
q8ctZ4Qae1ZfpypX91Vgl21ZVzcdr/L3olasU2Y1fVm6cNV5w148PKpxI1fRH5h/
`protect end_protected