`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11040 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nn7oC/bbltaB6y9f4wbJdgh
0G6WvBg4Flfb54G2gjKn24X2rlpeAdI4EpnLyqUdCLItuov09Rw9FfW+WOIeTVo5
hszs52IJf5P0hALUf/npW1yBqksV2uMUIknrR3YmjFFELMGH6mtAPcya/8LDqoTU
+NyCVPLPiKgSvQx7cT5i5s0IecABDtv/gnqdezKG8/nrPyc2uERqZb8UR2a1OzRP
jFBQ9e2U6DOaRGZ6XCPp43cIh8OwSdZ18Py49PJ1XdBD+I0EYecEtQZGbM4w7ydA
q9i9nstyjp1JC6zUVTN4I1FDmUrifIwLnIFgu7IzXE1jbg4awDPCZ/6nA0mKD1Wp
5IY1BvJsEEDOrmJJyDVvS4UPboRkVD4qjQ0BZBdqEqAo9/9ly2sfpL6lPLtDzI+f
tvCZBNUyswRu/R1Z2a0ocG4jeemBPJ9nq3xLtpuUws2QN4+EDeffIYPMZ+3neMZ0
5qev0NYLnrxqp9ZlqVFsZIK309lEA8vBTS1pc2umlwGVMBaFqR6/SxIirPaAj8Fg
I775jqgoPPqQzRZvSdkg2re8OopH88Cm2/VzGWD7w/yoAg+aduAnN2MjuMb/dAzP
fRtZeKlq9RYwVdku1QCfIC9/LnRwP7GflID8YKjFEYyiuhc7rtk7ujpFQ+107Y9F
3jtUQ1QVTeEMMsvtC7HBWCf67Khuk2AhJqMuIsf4+/BVhPYTHE7RGhmvgOHJ5NRN
qCykc9jRkLK1M/p23IzeT/MkaUcshK7ZYpurzohEoMx+qgojbS75o1iJFq7OPVC6
PZ4LSGmAhB7RM6HM4NrJq//jBNdcWi+p4pSDPNq1FfErBVkaIjuxWZHWLZWiLZ6I
SsA0ksGP4C1PDpSbKxBwetb8UcDCMsOh+ptCEmwEL4on2GdDjK3tFEfJVKhOjVpg
vqdSgHkFCsdzbb2A69TApG6OMROS4YzTlF4BUR2LWL79kq7YsQ/eSoEwCZqn68HW
iyeON5DsUrgzOTpKHvwrFjSybMVEyd4Rc+Su07FRCwzzm5eqkZvj/vj07W976VZ8
HwWUTKaxsifInCbOqiTdjfmj1sk3pdirK1kvFbQdGBwD69LbgZ9Ot0ArpkKa0G5E
ErJzE8GR8Mnf4PN2BpqsSuQylKW8mG7J4aMKBoAOwq3ayd23gh/+z0SgYNeiCrVO
FJil4fZi/+QlAMvBE92ZM6E5nI4GPeGsJ5IFlhkau39q0KlnMin4hBObWAO4iL3N
/3LV3AiO4WEIE0jHOfe4teICThbKZtRdR9vGe7T+NLNFLRj/oqnoHy9B/vfX9vhK
UAiekrYwaSwmssDdCCoyhW2C66R25wltPmjVTBcHiGkKu96K9gpjERVd11i6YuuD
wEPG5X4GIe7S3OqkrYxFyvl6zag5rLRieYLSTEq2Cbv+0MThb2TzhxyNzhew4Kc+
mta+M2gHXYO8JRPAqdWyZwKpj9vZlvlRzCeVlxY0igJD5D6uwJxqKnvYGRO1RwQ0
Bkf/TqPpfPRDGRg6k7GS9l9ATNMr660c4rhklsw3zrAOQGm2AWHBXSUxeL9I1Bm+
lVhgTNhwBfgvooR+Gp/3VwelfCwp0YLWxCje3KLhJ17jCmAytDEO1DnKIzoSxsEu
fBQQFHFLJkQcgBTxtOJCx08Ix+0kQ7qqvAOKz8vOewu8jr2EMdsV+qy+qzwVm7UV
ULTux3uuXDj1qjDEK+GnrHYTWOA3mUI0/tjyjstHaBU/nLxYA1O0t2R5g1z2HeXn
w0LVtViaxc1A0PsauPD8A/CUzdf5NEDlJY0mfJhesQoGbEXt97eq5jpo9suDGpIv
rpE7qxk8+E3el7R5n0a0rrSLIZbx7f/ZWr1zGBsPc+LW5zHupzX89cJjqDNSMoGE
DTNzUfkESwp2qnP37qgWywR5YnuLpT+y7J4JDxkFnS0QBGc0YbnoRaYdm8oOrHe0
K85a78m9tUCEcwL9UiYZQULu0zr+JlcDZ4qtacsBXayIiExyDr2SRCokm7VMRXgk
V1tBqjVO51U82ERgzq6aNeBfufoNlHdZBke66NCIFtz9/6n8MxymltL54vzb3OzE
ZZslgHPwQNthfD5Hr4B+E4w3cgkNa0Soqsd76i/OieWcJWble75XRtBbOJyqZ/nT
SBahUh4jvwMrdrcOu+9vY6Jye4oGbaC9qrPkwsLMNf2M9Vrg0dRFvd+x3EzzopSo
CXhQftnJXOxrsMZkX+GbFz7/vjJHlB6yne3puFGFws8a/t3I09bg3YuHgKfZ48qt
LrwNQFWtHLpVCHM+iO6tC2rJWMHF+Px+EqqxmxkP6AN0D7LW2NJC8NqIFlgobcvQ
DH5E/Knw2GQNrd4PTbWvI+ViWL1XFXm5ig/bol8rutPqilVeFLKmCee3XV7hWasZ
vRa4tzubhazhsgvIuJNB18JOfqZLUnO0HzjTT4m6r+v/iq8opEuq0h+Z/Tp1wAJc
RHQD3fFzDK3OkSALqHD7ckzmYQwA3Td63tezrNRiYUmhHDkMWNLZsPK42mV2KqA8
v5wYen+zEHLi4QD/zFLGiABh/9Evs7eLHDUv4BEBx9XxOKswsd36XVts3Cc6+Lgx
/W8X7Qk+jSRbkmW958zU/3/44wsnA/wEd76uIAQYSYdbhQQbOSRA5BbGUbIBXHcr
B+ZW5Ku8nv8o+eQmxKemMVNxhb2iogRaNJDErBN+CgSDlWQRNj4Qah600vwqUKPz
Sn8lwM57r4xUEbOaWGOnWn9bcuNGlyMpCxoHzB+xZSWBPhvrsDTCGOjECxxqxPG7
48GatcpgKXP0abXYfC8t14gTey1FbXnNgQZvAPHWi69D52m/GgfhYfKsT50d/JCO
xzfVwTl2UaA1NPth1Ry0VP0Nrfsaib2DnBwQS97BGnlH3dulN0lkI+J8C8tWtiRU
D8tLP8rRM7osiCYynSUqQrx0mH4zEDFKM8N18461zagzYiqVUNLn8XqJeaVhGxWc
eQnL12Si5fPJQjx6AeXtK4hcK4MQdJRtfqfAapqSu3xocMWyiK0qHU7JZNbmySnu
NIfbRuvMNW//2QVuXmMNGre07ECGRhdD8oTZ0QtUXjxWnDl8Md8/pljA1IzlxnJo
YWW5LRYmuZ8GKfhzTtIaGBzL4VTTPnyu/3eN8uyfLj7fXTnlqcKBebnFUQm8JRzJ
W5z0XYeUj+mOSExm4At3dz2EXcU3Wmss0XvB+n+rL2I2fZzMXl4arRMqkorRDFMc
3VPYrEnfhLuadgFVC8jkyvVgrfZDi5aFzzxoFbEDY7Z6p7yvPyUSNSjTLBwhn3n3
UFiYdCymNvm5wnX1OlIYXR+hYXAZJlHfjojSV5Hz5XwbziNyYi5fTdrbidqMEdTg
+qqg2p9XiHljhTmRFY/aB7OOzGE0tah9twp9uMqN62Gsqy7uBcGhgu8sgdddf6px
JVV/b2AIEOr8vmP4JQXdENhKsP4HU+VFeL0zT8C+s5WLcmx/hwW+eRV40byRrHRi
IGEklFX/05ZRZ7eEHE2rgtFjEDiDart+108EKxfWeE9gNlQ1OdeA+WObXwCj4t9s
S2SZsed0GyEDh5TFGc0JkBbC3hNnWXKXKCqSY9pGHAzPzx0Eu+63ZNSY0KtYD0px
Eh4ZP1upFE/ukiRBlRILfkExPgI4NHPAQRSCfmAgDZox4sh82n4Th3IIkGlOpRwP
3EIfcda8YUKyLhlm6fYkanxImXaL9BLidWDsyT9y0L7mafQ6IHTd9pPFVtrdXTAA
XEvXWD0YT/eoeVHNF418w+SOSPXxgFLJoEE4U9LhHF9OjKdNCjQ1t8kCksnD67Oa
K9VjbQAgvTK2o2/9DKpiYwlFsQd+i2LmyphciTb2VtQY8DKVGF4IVI/jK1+z6E78
vEZhKEdcjuYlOY14UR6B4RTuSLHTagAca/PZaks3zYmS15p9ArrHNaqtj6ITjAq4
Z/Gfas4C8FCFKcqkKYXWXkH3Lh2yiaCauNR+5JD7jsMWpsDxA0FJDWDNISfURZ6V
3tbcG5mx1dhW5kbkXA20qxfqI64rPQ2a1sO0n1UzDpKIcjSBg1uV4uXWR15M7OEi
KrWHkUCSgcegNWT/lyCBw2guP/Gieh5tNvpmEjZu0mQktYArvtn8rz4RL73/Wxm3
L67uALprC4kAd308JxkBrc4Dknpyl8iMvvy3cGshsrOc0W5cFRlaPK6gBeGFyxVS
WXsOSt/XtDplzPCAVxjv/gyVno6HUpFaJ933ZPLK2CTLaGZsZxKAarYSZM7j7x6B
cawaj1n5/pmWuMN8wlu0arCYP0lmIzgWyYh/XODP3NPGmf6mSwDEW8QtaZG020Zl
U9MO36G9nJ60l+yh/3SU+QPfYlEUSFN1PkblVWEXk1RKl3UWA3YtUZjoXo9vFI62
CqXWrzL5m9k6PcoQ0pSHiDZtadvBXNranvcNwwUspyqlk/mYD0//LW9Bz5GueldP
ZBaFoiaLlMkVYVp8QByELRkA580Cl4CABOsO8Jw2u13iJrEDsL9+AuWkdXAeKBnp
pmCBsq1Bk3ez1c/CPPr3IjpxHEV2yTiBFm4XmDFoU7IrfDbBTzTXgWYB/CwBCWUC
pbFMQPl1X431WEe1GHQErA3A2qaQGkJmSN253ghTmEbj/YAUcPx95Quokk44sc5D
wZ3o9n84qYK9gc7KYXlX2stpGGGpHq5/2LZRAdSC75JozOgxLN/XTWBWd+814U6Q
ChYYAL3HRbSMIUIgBwe/MNikMDEc/Afcn58c6ms3phNNJlP6yBJC4sIriJa1D7h0
N5SMOJo0mB/d5AOG0CDYPHv4aGW+kG9cnVJW5f0GrQvSGBBj3G51se2qYbYSpVHF
aeKwBaRAgGs/HZMTPwo2PMq+gw7os9f+6jCcYffj++i4wHi0SUQTiv1WuRS5n4bH
yYx1TU+5gv4hASiKyMZOU1PoDrUikHn4DnZXjBJK57ykkBpdHKkmr/YLflO4SjOO
bQEeBAt+swD6kFquanvzwzbZPehRex8oos6ITZ+BiatwEBrvJrLxsiVwYKTbxON3
meCDm9KZEEzlNs6j/uLDgnHWNgwS1pk0y9Kbs4vsH4u6wl38svImNifSy86iSFKO
2YSYYYImh0i6Ppzz4G2e8GPofVv2/Wa3eL5QARv+cemExNB//6Uaf4AShFkJLQUk
HyvbUOUaQtl4mm2vqPFQbqZdrY06vX6UNDzThAv40S7DXJYN1HKumExL2FkWIpM4
SCAXVZ157RaUJ1UEqqOsophYaqWqZ1TY5By9S2DsICrHq61lflrtLVpQ284NgrMJ
KW1EpNJrqyPqx5j531OI30WbYpPasgTklc32wQqAtXhrBwRnth+UUuIL/dwDc8cF
Gwkk8nrb+6Eg2FABhbzpEYLzJONc3mzcWWh92CBvgpheSOwqY2jv6ND31UKRyh9w
owyg7WOZTIovUa+CkmxVb2Vstt/Z35L85k+KK2HswjgFmlKnn0SjQjsiZu2iXqke
2/Ux77c/ThaZzcl4OyX5IZgADDuh0ZZDJ84GMXlD0v8tooCiUiOU11WAfFKpx2kt
EWS6P4T4Ys2lP2vTOktFxN4U4fDxTNU0qiMn7MF1gpDb/2sB2EaUBwLxj2boWWX5
g5+Y7+64ChcZZb4vtFFmyLAevYbaxbN2tuJLDxqotKImz8C+cLwGYALZqzQczVen
iaBPIGr8THVCb9fWCkmevNT6ocTF4YoPuOqA8RKPCkfpoX9YxYPCCD5nO3B6r7In
761ojcv1P76bZ7Y8/dy+5OVdYE7xUmiNqSe2TjpbfEKc+BsyuyOswGhg/2XxNjX3
65BbnaDEtlOqOMxIvbIQ2LlMzCU5IHrEuidOO7L9KPDod51lmqwa4Qoc1WsYB372
ncE8LlaNQie/B6es0VWacWU9Jn/n1q53i1TDXEkqy+lpcJHCSNhrYkRLVwBGaGaS
1s8F1e3DUonaMyQ6jRPEUDrip8gcxZ6V5RfxcRsw3+RQtGlPQa2HxzspKmlCDZu3
DCg5IxNQkSNWqOVFXUBkgcMaOUBJntvr/C9GmydpNzyWviQFc46F2ObMi01L3nYM
YwmuD7PsAjc2cQyICi0wgs85//pm8xLCIRZlWimz0LJCMNNxhktik7sIZ4wFJxKu
+doBubij03+wMWRQ356uW0NiBj8aUf5vHUshNuz//lsAWwZkDhBvQR6yeUQAe0Xj
tlwZWOADd/5zh6/nhfSyj1mSK+PoBjdsMSatIb566czgAeKlqWH8pseDmyldwb7K
/oJsHzFlwIXbVacTaylGyoeH1r64qB95/q9tIGB4io1qQ5ZFpc9BzSCkB90tZSsb
TSZAkOnskgvCouq1W5QCXFFB8TbWmSQI8rzhikjCeGrWA5vQpHtXl8+at3K9/s+m
WOrYuzn+bf7pSTIfH/FuBP/W2gF+K+vK7r+iELY4JvTlHXTUSJ9w4rY6ReK2rm89
hDexM2tRT1hA6a9Sw7uAroTXLY8CzsM0XtyebEnMErCfYeEPRKNmJ+P5WiSnEYFr
AbYj6kAvJdbb/UvdDPB4mIDd8ElnYJ3LH0Ahn0k5rsxlBwSfc4bZRlHzJCN5b2/G
7Pv2PNEioTz5pI1xi7USdANkI+X9v7bq5DoqCB+hFhrWzd2GPKmOMW5pNxr65BXc
/qeVWQQgC5pGGBDNr3KXFpQ4PF/RQuFV+7qih+0/Acd9/e0uu8p0n+K712a9v1nO
SGDQlq9ILSuGo0OUxPwH2lkwyFttZ7rmuYMH+fpBAY2+IBnwzsRVnv6TwNqiZfgc
IEZDSZQg+8VlRCNiS9K8xGoYZK7rPq+yhuOllMfxiwBs27RXFH4q0j68dE3fx/jx
TyWu8S/1H4k58J+EfE3H+qEuuPqDLqo9zBdkpGoObldEocJiS/uN+9f4w4Rmxd10
4uUxzppiJMYay2rCxSDzVkqViqlOmh4yog/8yQHgquJdwrmVBYHyiavZjplsqilb
GRpfubFy2nrUQhqjEw+I9yD/mj6kygjGUL7C9LEZ/9IlKMuxTccIE406SrUn5TmJ
cykc/uqKfC59Pyo3OAcbhPvCHAGxAM+IQ2BMHzDo8sVfybbFweqrIz0xwspPlF2B
0V/T+/SPojR8cW6vxBTDMbW2Eyrbb1VhAp5Lh8vzaIaIq8o9RM2Znrhv9uuCM2RR
qMmFYg5e3L1RxIoG5u8VoqnH1eY8D/d+5DyHQ5+cW6LtIc26wH4JDZFl7ChKAMQ9
Ul77lBhHD3ezRgAArfxz4UywCZwyN4w64xnsSXeL7aSUlhgUmVlWigCpcrCOE7bK
zIlyiIC5jVm+ONmZbTovwAQuEx5CRP9DnKewoIXqyUileVX6DTtPgRLYkubi1kYK
vuZn4VF1YcJOOsRETuL4A+XoqQw7RxlwS+txh9RbKw5wujbOHwK1iUhxnKAzd6Bw
BrtSuoWqdBmhj4e5PSS+gxZBwe91U/ediZk7MhCzrmeZu8gLkitUuV9TrnBirgcl
A/DxCcRS8w5kH3wbDm/U1JPkKCpZI4ZT7goWXg6Z3DVxDfodtG14TleLXnx+Q57z
8HzwD7LUGcDEcWOVCtidt/hn19xtj5Cx3VrbxTdNAxshaMRvMKRV6ZK0h6sbELCA
TiFdtDGOV4TY6AI7oSalxOP4xO1bpY2EhIZ86k7aM+MwaMI7d8NTc9sZa9lbfgww
kyLcWmP/W+nRWRQNQA5SLf4vytce9iYxHc55JCrn8FxIuVeHCRtrrnpc+jwpts6v
yq0VS/K6JBrtgfZnClv4+wuuWAgcgOgv0gQV0UZudcZlduF+oh3xcgDwwt4vo6GE
BnP8bJTkKvEMP0XIYx3g3A9sVMPeoKVcBkSrwVgf11//LY1xoPGYKbNsoY1YDSuf
hwMOiwFYDcncPVsa9+azjGHAHCLgzGCTy8Ym0Frbkl2AIS5kx2tHDczLuOiDzxOt
Ux+QWEMcOHGnAixaRgvsW1fwU8E7+uCUOCdrY82jMQCOt0PKOtnpdTo1OJfnU9iK
oDI+LP4uDr/dLelT1Ml6ac69AqgKZoZCLRgj/mn0BHwUEkYoPp6NUbPzmmRcMBwQ
vjf2oeqrufsSeeeBX7WJ2HTQ0HmrxqgAPNs6NpXBzptBHH+Ez7fCA1KXgN5EgSEb
+I0vyhSnSnFVWfIr/ylpUDLe682NhUkWrzwYr6DKQkS9SB9vGmQX2icbzLS5JAvx
wx6zUODoJ9RPnIl9BOGCtW2ST10Zur/oI9jBjxBa885TUn/exqADW218LsPkN9g7
XxSc6UHSTXO1wkDORzucUrme00kwRrQbXFDqsPdQ7INYy+u7j3lMgEvRCSJ0LyJk
ie5UU3ayEkqsQzt41bOobRXwCJy7Z6E0Sm5Fisc79258vMOJdwKaftqs8OHpGGDi
uv782q1pSIAiFpXj5UP9GHnbvDwqU/iaUVwbuGfX9kxSa7wM8uPpV84v6hFu3nAz
U7Bstsijby1ycTuOYh3YOfAc/4mb9R+Yz4Ouj1xw+tYPhGcJ68TSWhLgtorIu1H8
M9IzM2ijoOjPVlVZJHZT/BKuOdkBjvEt7FwuF0gClV8pyvaQqf+vsrya9ubJo+a8
EzRCZZIai34AIThdm8yH68aIZ+TjD9AFZ5XjfJJOk+dLVQftjShrpV6X1ahgZf9C
r4P/UZu40p9HpXTS5ZovO+VfvxmGeRYu+IRUOkiKNgNy+WFuOOVe/gwpvw2F7ZhK
ZoKNcEFuw1YcSW8B4HF3fC5PF0c15DWqZ2VhtTOxOFB8Z73928KrSNw8TkPgb4RU
uGm6pDYrUEVy7zs+YDXAMfBi4GIMo8tfI/BlokDwKwwolG/rQO8E06NfkAWCr3NU
QQheYHqgtmuJP5sHxm1qTx09TDcTuxW5AeIgDcie+ucfUsuowq50GeXxqbJdfCGV
n+8sKue3YGmvzkNIeuMcNtXAqyip4JkKuvmpkWxZkGfiTDfwS/ByCxdgvl1btlM4
1dTlmw4xKYV4H5ljP1TflAx21EbVVIRNVHc4tb62/bGUj7PYxB6nnZu8dKPO1s79
NIjvWKFaX2EhnUN6OGc/ZW1ofB0w0X/2kgJ7TqPPzL0mzuqKFhPig96SzwoS8zVI
EVVR4Oi4lNWMjRGWSPWT/ccbZ31MM4rQe+pipJ9vXze48g230skIB3zXt7kJxDhY
ykFfuYVWUYQvmmAhLugRV1UvhTPqysMJI8XUKc6odPMd73ux2UjxfmZ0VYY1T2NB
5Ek9F8WoHC2fetqbXRey0O5bK4iTv6fFnJuEdDWG+PPagarY98cE7OOn6rbFrQtp
m0Dtg7XQFJDydmo2XXdu7kjq/V0fDhBnesoVNkYaU/EwQhSRv20rPQ3pT/P8BXOh
Avx5lLlxBByFVdfVsiv1gM5taAc2oRLJRVGJBt0xwwuX9ArSuCGukSKPCZRC0JPe
90FL5p5rLgdXKZLJLdW1vsBVPSI9X3VYcb4gSAtoFZeWT2ipfHKsj09KCz/kogwL
rSJHC0+ErylmEDqjhJMimPvZVRuKkWoRdUBRRfCndMYxJDZM8gdn+6tawP+F0K/Z
dzy2k25T4u4YcojI0BM/K54zdwzR49rtHBWjxpVCgN+ycFKKwifAtIWu41sKYtQj
OyoVqnmdcz/KadA1zKQQP/4HyU5eK7BWy9gNBSqa37EsypBLS8IICK14CxC6rcZW
GizGs6JILhlmNACQRct41WQYSo1icCqETWU0SVCH8wXLOn+n8R9z6ip+hHLmZmPM
5D8ipBb8aVFzY+f0Wq9AFSGHccn67W3GvwI0t7MGPgZjvGTT+jWA4VWEG+j6xQHb
5/83CflvWzeD9SX7KZJe1SR1PCgTZTgX/hNBzRPYlYinQfTuAQh4eWcNoprU6CwP
rvqlopoUxXSrbWQ/qOFX/270JL/e2VZmtafFKyVzGRKzL6dTGXQag5iKL2Fixmq9
GPdCrY9LoMXv14zp5sRLkW5fVBay0RGJK+TD0iQh9/2YIJjZaR4BbLwBFj0TotUh
t2v1vp/qRp26kD4FxW2NGzIwPtxinUVl0moz/Du2H8G82dFqAEpckKe60c0EtS7V
1XPs47mlsDh6MFAUuDO/hbgsmknIQ3qLu0ssnlIaMfphwfhyzBCbdaMnnrcmUiHq
G80tQtQw1xA+a50if2UiYmwKmidAQEfgqJm45bS4vo/NZUS6xvMYXceeV15KLgy7
+b115w99xWazsB1QS5k3d7Xv5R8n/HqEvRnKlk1scJZzV4lEXD7tJmXXNFxZJ1iH
nT5hQvyvnGAQSXPNs7JCL1zkdXZ6FUuHKoG2nt8y6aTkLIHaoCL7v+xAwTH1+eDx
7e1XaYcqUb3BTyt46DCOEFaHDtE8i3m/WxE+BqUo2dOQKoVJsXqnn/WrSnllY5dL
LSQFs0nqRNed5vTWEI7dt4XPtr0EE030By0MiCIfQkz+QLch6+XhjfrG1SLK5/X7
UMkZLvb8FiHYOUfLoB7xi5upSncgKSGxIhj6pF94hKKdlGABbz7SOQyMTJgzFlJj
R4/hl8pX2dFAvH6Gi/fd/OZpCIs6uZRvQIMksWeeKqapMboHGI00y2vqlH0MLPRD
jHJmAD3gf03SSBCBXoUALbeVwb6YFDx0wczHVLmUb9gzLeeS8cC9Zd6v/vFXCkZf
/mwS/iesWhUs6xeuk3SJOIMRbxGKA4HEY8StfXD5JR9kVq8NW6CuuYT+D5/YAUAh
GG7OeihzSYxhKls26chgfQy/pmMR4Mm58EjbM10NxvR1pYt6shPTghlfwWFlhJiW
xQbm0Q6+xULZhuPtUDOv43/OPcaWs6aQ8+LSap3uvQSkur21oe21DEzNb5s/l9P8
HJ6gP1/1iAQ+3Suk/6jb6MFCWxwMhbzhSQPNiAKtGQWH2/B8YMYREu+3yzHJsAoP
+39Zs5McNDLIfXMY2kgkyDIuWF9Pxx5kgRg3dwUKpNBAXs24j4wgqgFcWXlV/TP7
F9e9/xULJJYpLCQsrJx4aLEPvn62vhKEm+6t47uxDgodVCsZIoiXcjuh4KbV/eQ9
xfvoCDESgkftlUi+WGT/XmMAl7x7BZD0dYiZqAG1f1P7FMNRoxv28JNhWJkp6YD3
/gUvdQ0pHZroaH29a+OwOuHW5yj8ttcNdlAD8mDYvdPyafM0h8HkknKzc6ta2px9
3L5db30MYY+pEyV2JvEgs6IH8Am+tuB5pH/W1ARYSkI1CCQCzlUPkg37Nf23jcSw
lZOj5f34LgK6LeyAVqmztLXpj8GK47ifjIOkg0uETUR6cdPqr8u0Eph2GuQC0YUJ
iEXFQgswTbXTyy0zdYM3qntU43JXpwC1S7BaKuR04ehMLaif89sWFqkZ1voLrmX3
PdvSnZPmZa2/Q1VLe8CiRnxipE27IBF2AxejwrQcb6sgvrZa44KH+INk4zzymwyX
JG6Vcljlga4f7rfi5CTx/IQk0iJQ7RedcgqrXtkNikazGTXCwF2ehksPSdodnpGi
z40tBbmKgz16zjt/bjapwSP/igHl0si0tKquY7q6Mex07k0Ei5YaR9lAAKe/DSb+
FD5i9bMLZ7QtaSmotNi8fS1zn9XX+IoXg7L77uL8niKHeN2CTZRUC6/ndCPp0ZdK
a4brMkkqiRA1G9rwCde5oM3gnrpIG4XS7cuuU4UpOr9XPg5ec6s0u73Ak0N48yzE
TiLi4N/cQxCdPIAchiwwCb0Zm6wNH+gQCnEc+Io3L/XQ1BAx+RAXkjc2i7JP+HuJ
j1wqYCGvl1kYzp0ir9tgCakCsczNKvo2l8CgGx9e60iz1ULetKLOfYiMSlbZtWox
cvosuWjTAGYEkSfG4mhXQ5pUH4twa/VjLeRgoQfuqCXIacXIwnScYYDCvA1LdN5k
+nkiin9TGZ1JmAytv3hD8FCMfUwAD1UlpkP6rZxLkZNuaQyefC54SWYfP/5fJFl1
qHIz7We94IFC5qX1sUv/XqNmeYdGMfBCfa3CrhoTt/DzM+SrY4KzqgU2I9IeAUv7
UfrveqmYTca4nNmyxohq+Dyx0wWHX214fesujXMiptm6SfC1Z2OVV55ezCeTKYsZ
wJQxY2Rcw/pftPCLN4b4g0cut9KQsz8qFdnySliVOwadDtWV3ZUvtStCO3clvTyC
5qzZN4uxNvJ7mhthVshHLkZkJDWSxhsTZmVHQJDomf3DAgZl/4igrGR/e3JL13gl
j6voElu27/PzJMu1KQtSanISfYhqKDWSwanPe/Ke48VuOrWXvXZL0qnMDk7PQ6IT
OaK4V/zYV1Uwvyi3l5mbV/zWS12JWX8ThouSl0TRsiwzsvGa5SHPr2Sbn4wGQ+qC
NqHWN+9J4i5UnmG/D7RjtEb5AFlV9LFHeg3MmcN145W+yS1v70CohEnEKQ2qw8CC
vUlL3LB24qlTbDqFL1nlkXLg9a8f8so7zc+LShMNPAfhr+hHhoNiKQdNcNh/NEHl
OYHV3IMC9YuluHUc2GiBzDT+0/OiQ+/5TdfKj4cYTGw14WQdSOqUw4x5tpqZFjHH
Zt9y2yLfz+dwBn8jDPuKCnTriZgaOp5E6al7HxBzazvLfYAJOJd7fFgQd4MwiCvp
ZgSAPtPt+isRoG0PXmm9dEC8IC1WBA3zozWifgzdaoAVWz4KLbwAsGBnyU6IFNKZ
a1gE8N3HNMPfJRG1LYdUP34Ur14Tdf9UgW01jT3yGfdUpy1gPGI5WzsbeonRQGES
QpYJ2RxI1GkBF1Ox4Frx3bN4uVQEI8h9AJLcQx+Z/D/l/W/1Y5ieLNODm0eI4mfn
ww5IBU4iY3ffQw8lLsr1ne70KuBEaQw70XDMBPsuufkGD76P1N4vriSY9qNhgWMY
3v2Lf0w5x8Ezyoe1ZGZ2qOrbNTt+urNDZsOCWAK9VR4S5ca7mdQgIdK4wQKzGD2M
kcM4dcKfZP5t2FX2NRvn6YAzbnF3/OzsQ4u/doxUWT06J6OE0aC89mwB0BloUdFk
pE9AtFQNiHY0llqD2q1ToZRn/zvFwEErSLH3Mm4P7KOuG4MPtnDnIC7KPisH8FGM
O0BP1tdWN3hc8fzFRy7K3NLRq9dqUG7YhjPspFIhK43q0kBZ0jpdZaY47p9btBfa
dcznNUAfY3esqxUXp0/kY6R7SbaSD7ipR2DcHJEr7fXTOXC/lBqSFx6Zhxvym804
i2HBg7iavIWaYS79curPyR1+gIYKUAV5UmjmbzjyX6aTSoF2fV10JI3WpoI49RrD
M0q/tW8IjVjB6lWQsKmB3xJq5Jv9wFlu4T/FohLU0ZEOGmIaudKfBvPnd7wI5Ntg
BLZV6FbZ/168DinoYkxTT1ulDbHWU0BeIB4v7czDcmmtx1cAdCWvcAiY3bW7Ms5N
l349/F3bjeFRo1BIGpv6vPYCjVOKZisAHdQJ6J+/KcVay3iH4X5ynpfl8As2oVF4
ghylKT6PJZu2inNVOS9wRvYaBJl0ICRp0ht1C0h3bEMMdNXKEPSLWWrcqriQO2Og
Rb5UBeDLG+ZJ5mIapulGSdTEzxBmMcNCpy6R3od01uEXAv+M2PcywsvuS4+7EnKZ
5PvB3V8ZWAywSP0la+uOoZvvlAQXRtEXEK2NGNf13NeupMZ2J3eUwayLPPqd8KKx
hwRT84ZPr7Hf+CP58sfotEMpCs9K60SZO8CeV01CQSUcZ53dieNSR3PfmxbvhC1v
l+sbJ9fqgN2NXMFjZmm1nBziyc9YiSS1YIUYMGjhcVgC4CGcRAPtXcDsu26SiMXR
Hcw8JqOEjga6oOLPKN32bJoT2BbnxenKmT9wdnniriXuN2zhFSJaxqPLIQWvG9g+
WYkmTXlXyUugnWzLLkWo9jaB3P/Myt5O95IvkHjru90Kwu638jAaPphWI5EG6IcD
30nldRvWXTs4IspHc+9gkLmyvE/+X6RhYo8f7zfxeoP182AFj66as1Pgl25nprm+
y8zWONQAAgcSnlSHTJ1IrOgW0kA1FnvGWmkcEXiBh5P7fCEPy/fw3P3dnXvi1+qB
VhfsMiD4vnmuHN8saUcwXA1hERwBBNt+i5dx39xhw1gE2Wg2m3KH1oWud4cPDkiD
2Xf8IMLo1DXYjcQ+AlH2GOSZWjXNYKyimnMYNKzCX1qq4orpNi0OiIhv/vn2tYnp
RywQ6WximGEAsYOOjzY9lEMCPxeT8xmOuuX0T4eWJj7W19NEkagyJMHGEqZd+pjf
dDaEiZtcIey1DLZLEYeGIWRkeLgpvrFN81k/154mWoWgJyp9X62E44L3GwT1RE4Y
R+6gW5X698odWrDoTo2U6cuNpcLjdRwAUc8AwwZQ3uJSYeizOJck4HmBvuuLGuoA
sMW16YCDA/RSk89t5fJEWlRI9a0jxDKonC2dZEjzwOc4uATlb7r3FKSWPwCY1nT0
2Fw4+uWYgbJYYbSlNv9T3qLBmSFMVrfYTBZrAXUqSOmVcWR4HSBlZuABwj11arBb
wc96hWXrQWcogevgSaXe2lg9FMFhjiQEvnZWttZZ6Pmws3ndKy5oelpjqw4TRAN4
LaWAeNSh5h/dmZC2E4bzPPm87cZ1RAW8FKLZ4OxzAVQgabYRbElHBvu4gYFomvIl
RCknC1VWMAbHWsoY+obfHYsZkO8MgzyJ1E7EI9x5MXck5O2jKMiq5EPohtCN9zKf
YAPkq7bdk55M8hpYsudqqlhnCf4/5yca7DTYqONn9Xz/ceXy1zvmT4WSlSmOhvln
`protect end_protected