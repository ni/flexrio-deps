`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2688 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
vAIFc5b9WPJ19N59E8is2hvFpXlGt1SqCBlQRtPM+lGRcT/lPDnqoAQ01iDgYm+p
QFKEePZRdqHfiWnDxXXJdnVqP6fKSGRFL9wDooeO9EEnHqre5zjecugCzXiXpZxt
B+tHzq7uyMK+46WjYg8twgj8UeepnX+SXD7E3GAmm6DbAMe56UepO9ErLZxsfGqa
pdBcWztq57xs6CoQ3fePxmRP7F9gFPpWWiV7fpSrOXCUVlvT1vhrmMwRCmkyAn9z
Ur3qbZHk8aYI+AeEGuVRG1+0QkYVZa815Nykat1eQdSC3HB9f4EXzRDLZvHZtlAe
XN+MxLQxZzIU4EtqvY/RkQG9DSzMX2cDCnq4bkAM5HVe1Lwf/hq1nD8FB0/5Ep5n
Or73d5pkDaYlJJ/EDtHiXG0JRbXsDM+QTzEgLDltwN6lL1yndZlJ5dqOx68KjvfI
eBUHyQQjRV3e0xiisjaoC4Yu06jaL9er1HOlyT/XnLoI2GHVqqupEZ1N+Urb9lii
D1j0UMYafgktZDzY2GoGqYT49Bg80YVjJFqAKKnSfDheHNthnfGeepi5GvtUqZoK
/wadncejqzSrbhhgGR2KDRzkH9A8V6yJ9amRBBt5aFHj+dcJ6bo/5ymmwv4JpwVh
u/Lk79GRBf8zh2MIIA1Dq5D1qgm9wV+XcBKpbNblYNj63PviKmj/Ppi5InLf3HZ0
ZW66220AMPeDt8VpiPIAPjm39xoj8F7V09CjwSfw6zythBIxVdptcVfOvbszUgR0
UaZtl40ockcJlPcwdrLqO+HI8FTtm2O8pUy2WuHK88kyjFuQX8+2+vBifK+dEShq
rv9bgNamaiKX5UHp63gtCh5vpN6FoUOx50mxJLmzPHTUVHV2k1PW86k5X1NkvByu
DM1Yph636R+ac1UKJUyl1bO9JjTqp1TkrUgLM6mnoSCamR00a2llnWSL+WSYh6Fn
jFQAxlk93R9ekPeA4OeoZKVORjlm0s/uuovG1ts/PgDLXnQ3qtrL0PRejELYH2Ew
5n1ioGtr5GkAyrMvifLLETfdoeUiPcLw8iWRjQmdHguedScmA9fwLr7H4S9akDbW
TLY0bzvqzJGybli4OvywprhoqhVrcsErVkLxvNYC6D04swoQo7Z/q2+E3M4tlb6e
ml4JAyBWpUP459s/6gbgfAogplN8YlQysGi00tHQtiJMtOzQTziUAHO1Uyi2Zz7S
52O7gK4vLvPyeW0FrL12gSXQv9O7UyEcMzlB+GJZIH8dxcVPtUqdOF0uoSY51l9a
ETaOqSlQYtZnb0dwq9Af4ujvwjkOXTEVnzxM4DX3/JjLc3rWTaSLYlqcF1Jjqxvn
FlhQ7YcP2/OYOj639iCh1L2xtu1wgQlOkojCl2PlnKG2aytNrAoDeLMRVxI6V+sO
c3wmguQWY9AoH18Qa3hJKDc0nkx4aBmojrcObdxqM03FR2Tors6mfGmQmB+vPXah
udVU6k49Y5W2wmLPsSs0QYxbBIWoo8XEO8TCoSHLNKLKmFFKqEO1+/Ci+X832tVd
KSWIYhNUPTbDxOFsdIupLOQ6BBzpuAfePo87eqSoaA/gchOcyeq+sCDiTG+kJ/mu
nOWHhVqOW+2hH74Xhtg+v8eS0PVz/l1Nqn4gNEmJxbPxoxB7N9PjGYaJ7mDhohtw
V5cMfeA6yGa4LcCF1+a7X5gQHdbspBFUoHt2k3x+3spnym7Fx9jhhXhiWcKkPG8y
4NK1t20eaUv37A3HNqqvVl9qWcEufnHsSryU81qZU+K67t1djfTUc7hSX3hdClgn
MD7+A4s0Rj6AXo/zEpXrDRBtGrUuYih1jt8cDyVnj8ivv1XCHna73GTzFUlV1w2w
msIY1Jx/nwQgYoYKeOlEy3n0bDYZW4o2lfCS3ocF2jfzdD2POWAgwHCTKWtASTYt
NQH2vwJTX0a6sIqHML+Cb7P8Jwe6eIIo85aUhrmj1/Tsr3UpZ0mPSJ7k3yOO/M5o
INRBAn1xaH/o8rxKF3COvysiIrrk0E6l6eS//IzvdsvmsPJ8CEsTFoz4WI4UgzfC
XEak3Pq3/1jcgJEa8AuRPBaCNndWW+CULH8DI0ENqTqlio4yLCtgZ9cwAh/YmH9a
a3QZBIxch1dv9GygSFvcs95ekANh3kExdYGRU3gOoI4EJ/op+FdsHlmxCUWhB6pS
UN9VDOoIK+k4y8u34cuOc3JpjruhXvzEgBZYlo5jbo16e2/BS4uNXlag+6DQNbm1
7Zj5CdXUCAR/ph9Xj79rff7uVz9ml0UPb9H6ZzjDtA6NXVQdslxwTFHZC5aRahlp
RtYdaMTKNDzu2BYc2294CoMjsyZxntWPRvLec0hs5cMyKmAmY8KfrMWwAvyevWMU
j3OERbYZZgB6Z21ifbKAvo9xeLPbAeTOpZ4y8MOHszR8ilm2+VPzWWjY96II7OdO
oLnDVtrCdaJHi1yeRRukTsAKVuth1VJuG00Nim2T5ySPBYKyr9HfCWZ2FhV8hMFn
ZjQR6+evrsqga7A5B3CTWyEZk18XMOEu7GTDzQeK/NOI1gciKvtLHLa9tmBwEfYi
eMUSLgWY4OHFmk/ufLJzE7Tlru6P2/XNtK0c65oNPAQ8te7ryS1+WpBqZ+sKVwyw
v+UkMnwxB8cKB3Qvm42QfOQ1zdQMCxQ7cKfbd6HgD5/7M3cGqaZ2oTIrMx9SYBtF
mlg8sk2csrwmAvuKQ+GkOo/R/+SDkWFk8IIQ6PzO/fMDSEYqbuceSWGMAFbGKmPR
tL7eGpHuOAkejfEMP2Z06dHEe/YDtqQ9aCdoolEu1twrpMcyQQ9Zf/HPPGkBcXtt
OssxZ87acQagZC+oac9mxN85OxNXW4I2fgVv82+f8nOVha0z2k8hGI+v/u2FdbwH
WlngK6n2ow7DVCoiJs95K++XOPvCWoujBcGLAKC0zAFL+suLyPhS+ULX4chR3YJN
rLhORBpxDYvJkrv84GCNH5df4AvPdhfbKkiv1yfgB8NPxcPwPgOrsLk1CQrUGEh9
Sch+BK1ovMP6Jfkh1uq7YH+C3APk7NJ5017wTuHZvRrRgBONS5I/i06m0qbleoam
CqkHRGN4hza5d5bBtad5nZ1a/c1JDpgodY/L8FWTlCskujODZGQJf5ItGGgV+1Td
MmpVu8xFSJtXOCbsXfQ/B24puM+TlxA25GKaOEU4cRQJxWxl3OW29/dbiX30Etre
6AjANgFQku9n1LChJTYSsh+2oth3iZfe70MpeiyumZ4RUqmdmtq7XA0zDNPwcmrQ
m6/9VAn2/6beuTAYfklTrJA9ubOhysBNIVWX2SZGs2GBd4flX7D6cSfYl1WWwIe3
6EeuC2isN8VR9VpYbdNfPnRgnvYnapRLC6vYNpRWItYBoc6c/PJu26HecU3ZnbwL
ckdAYFtJowHC307/M0zkyFX5j5Vn1dqmbg+6iwO7TWit9+NcH9g5uN4XpEa9w5u7
`protect end_protected