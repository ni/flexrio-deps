`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Jm2uGAVYfY7w9Y5qKstopObZuZAEY3b/Io3MSEcWLhjjnKulVhCBBYAEQrAzzGsT
vMbffkdZgjdXQUg8jOLJXSHZ0Dgbnob2vlppjZs3bgyHCF7MoJ35E+LOsaLimUA7
hlqStcK49hR1hdeBPr/OwfT3UeVrRtQyq0eJXQ1UksinX1G9Pz3/CmcGfTZ/C72x
p9icpt0bkY4/1I4GBvNCsA6FFKH947JqH27OPACiQQRW/K7JToQn+1uhWr3LA1od
lbVrWu8PdZi7zW9gK3jiW5GaPjwbYQGqeGFs3bTKBILjb7sYHxfxw7eDLVMAIu5D
W+OTIN4JiHiE1gCnNEvkSQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="pm+c2fYA/4JT1uhlJGVUubML8hZi8lME4xPobg/m8uM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
nBaXksR//iZ9fraC7WMJWWSrjqRXHxmM1Y0+KKN3b10NElDzVNMlR76DLrcnamFd
2n7uzsxWqhhJR5LBl98SXO3Y90J6BMbw+OBG/MFM/zUulxh2Si5YK5G9GCrG9gvZ
5JomxuZFDu9CzlWGTuRUt6FsE4Lr6sOL1P+hraQDpMk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="M8TXDiNa0BVMX1P60yIvW2WA9jKGGy8GtbuPknDnC9I="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 57664 )
`protect data_block
/5TNZvs8Nu0G+mfp7M8H+iVAGG3Mh5DYZ0Gn3rRNhV8b5CcJKgjQajrRoGl/gSxp
rBAhtT8Vd5eelHgtvBjpvFBA/EBUrRH6CG6pqRt9r2qUDt4UernbZbxC3BC14KYF
RNY2BMuh1OsxGQlxRGFb7uIlsh+dEdX7wN4HQ808wWVdKgPEZtzcNrAxF8KIWBBZ
CGco7wwsfDBMtt++k3kihE8VzAxrU2zVmAATPcBli2wRJDBAbWWhSusJssk6D+qw
Fp80njtNSa1Z3jGfG8y19f2gih1EIyapzV5eI/qzJPNOPxb5IXBUukC8nchcUjar
cNubWwKs3SKebctrUW+vRg+CpttOJp6Q7RV0+K/TVFhQ2KHNEoc1YRdBRlJS3EsL
sYqglexxE+fhLH5OTM8pOM7uAyLzLnbRG2ztqqTyPFgPz7Q7LnHSEPav0omkuavu
j/4PgLPrfnszlSFJipXmsnEfhhZwJSuSTpjyECRu/q1I5dVZvgoLGZB7TcreSBJk
5rcMd0FitzuDHmhIIrzNldCrncnHwvddks1SlFbJ+h2GQ3e8/k5EV/XReEYWsqZD
ZYSJ4Iq/Vh8MA70AKvNiavAkx8M/4KcNaskYms+VSGcQyzp+SE7wywIN7bchMxqw
0DMXKCAeQTN1wGxqO6w6eu1M3EwNPZY2bQ61uRYuSlBMqYKSZfcWFGB+i6xTfdB9
gvPCn7OyyqhvPxfNzftBUveA6LM0jgkAi5EmRwp1w70iS4cM3Gnqzs8MbZW751bs
pD229hFFxyNCu7pwj23sDT7/Vx3TORkIpXIHLO072M7/UPFQhZuDbZ7UvsKHxGyV
xsqsbKbUfCjwzV6IzwixdVS3D3iAXup3Ovapog6JiNj2J4gyCx34N4ad5ylIcWKp
+TL0hc1mMkDqOeZjqBJraiX4Rscvzq4nut0v5Y3F+JyGZCFtIEaH5EbREwYPxDOS
NBY/04RpsA7pFENDoTycGR90OJ017QXoOb0SS4qIQt/D9+a4XO3bzrYRxgNDQ6Dw
xVQLmQdGWxT4+BYZnKTYfgRZkK9xWahxRlfI4TMRsPSEIP2mWZJqhmRNHdTlPjI2
/yKb3LW0Cvamj3KIbjUewwu+nvvlmeCfB+yTucj8HLior5e7wCgTcQUweG5YoxiJ
PXTy7JSVAYri6lEJxfRURO+/Xmey2TIDXt0M1koN3T53U/xgNJYqqlOsixpbdMFI
o6+sAyk0o6bO+rGetMF1kXBTWJMtfleAsZ1HnWnRhovBj1n06uv4NpLM3cSm1o3K
CJuT02SSa7QW9np/F3b+urFvygpjFw8z7wRJwssBLlkx0yMhxdG/JBNWkA3eANTT
oZFIWDGRRFczlYoM1YSZ14d3omR/WUzyQeU6NfBjEAzeeftzhJP1l9KkulqkjSUv
pOuGc7anLDHcwpLhYh0rmsWn2JKo+BhWWb9FYcKMXVCmHNF/cyFVvvLbdgWpoMd/
SIbrMpk9PEdj+Pf2skS74EWan1nfo3zqHjoWZ/UhkQfgVkeii+VBzXC5j17i0402
58yqaoi/a929Ovp8u4f4b6pNyr3H/xUu2YIpJWkZjbvUEUZYxnkrMgBEaQDctMO3
IbjxWKSeIKyuYT3uUUTm9P3TbrEfToSN9QAFnjlAlAwZDBfzHFbH9yNrOqnwxqpg
C0K6tuClPfIb6jnxnZy16CFlDSFOL4EQbmCFmWnfwhdfQSK5/m4qyJUkx0H+MIRq
MmsniRnjYVe3p6L5yGvgPEUAH1lQTpV4GSvkaO+YF9/l5sjrRDGHPmyxsvAMNAcq
y6fzmTPdX8nYs7v2EuVRY8xqUsMv5meTTrBwctyic3F3Mw2TkVLFQz8LhbrffZWW
TgiFrr9wYfTZM+UtMFaev4L+0CY5ujeML6luGFNNZ8963+eiCLsKBFP29Fgn92Cz
jbzg3gNMIsUE1UaUi3YNO+74ufvW+c6RVyn5wah0S9/lJAgLrzqwUqL+LzD2YWcy
Q+EHq2un4Kq2b7eG1vQBt+PG99aiRkFZ4cODkBMd3j5zeKyX2LolIBc221mSKFLl
4oupF3uhMvqaaeQRprGrKOqolCt/TvqJLTvxKDFi0ahR01x+6GIZwHTmQL6YeTqc
K/86oaNqgFe/eNO1BTJPSbze/znatLW+q9BCz0szbuKLQa5Cznknw88ZIiDwHgjZ
Z5h4I16Y3+/CwA8D6/cyRTY7OfnjOZYLE3rKhj8iO0uNWWobSUXtLmayb0MQJKiI
+UaruyA/5ZaE1ofJd4gl1zXXuq9oa60XX7vyku6R7Qs7FxeCu8rzV5l95G+eAaVg
C3ba/96wTCEO7a4EC28ATyWbV5BT46smH8IGZti42qyfzpUr91+o8VcTA0e5PuZj
0uqvyRG4F0mR7o7cnlCuf1zNJdOF+KDkGS27rMd8V0AaJjFBgnM8lBLm0YXvOVRM
N6v2u2eLqWv3qC07D+okYwWatrvjieO5uR/8/JrBPCJK/BHmFR6vFpQmEqwhM7ie
8A5sr4HsYLbciaOdQkKKN1IZaAxIvzcukR5StIK60QPB1YcQqLT2JaztTO55YjsK
CunUiml97H+/gp41QoBfLGuAcs8tOeXyEOwMlJW9ddLT7tSMAQg8M0LfYEXhc2W4
MOe59lbx/yZY9TWWrEm0h5v6hwqP9Rem1D+9mkPopg3XTjiyvG2tLaFkBPmtG8pf
qZTkn1IjAipVg0xcwDlPPJMOF03qW41voyzTKETXUBHDju+aQOXCwK3XHnK/ljae
qEJ2fqtOBi8jCQ9C2VqUEN5G0zHuLvcWGyifeVmHEMd4jwIVfIKQbCs1AA1YorG3
A9niYobvzpchZStX+1JN/bnO2g/M9ibWhNU3+lIKAYhtftZg3EWvszvjPCCStkMs
Bg3Mxefxt1kNj52kleB6Al3h2RZhHRfv653cTlMjl56USeZGVxbS4a6u0TfQCA4c
olQGpe5fmlE/Smlg5BGLOrVN6LUz19r0eJG3rsLsOLQDZEiUTh/g4SQFdH0ammpl
+jscz6boBTWl740sY3MNIJRNsN6Vj7E8/l94ZHjL5sztLzkCq56VijveXoJRY3PV
OrhMXtuH0suOYjFbLE27Q+ZwuZDyOPDhq2SGC7/Ci1SoSQtY+vij9xp1BWZdvrFl
6pySG+kSAtYRXnagLUyJyo/whzSf2F6Up1K6izdyQbOVM/Zsmr9j/44DRWmJ0Rq2
RtLuNFP3UgYS+v4VWrmVWir7OlY2tNsbxqUn79gBdNE6r0STHM8aFZf3paNt8uTm
bNWwsrdWXSg2jm9CFf7eg1wpg5DXbVrSDv4z/VHQaGVM+QZYDAFywijVzZmh2Tcv
73QCRFzLV79S13w3QIsyhiOjMyeONi6bEeTjiUnPxe8roKvkkBC+qpOBGTaANlMN
+FH2y0sAEIhzjsatkA1j/H8tqYe8Yg1QveQ+m1csH8FMYiLJOmMVZ+Ks0RT5fvxk
F06hm5VynSjoqLUlHYxbIdv4bYBak8yLBnlpzMwZY+MDkKuvq2P3J836d0JLB+JU
W+T1ueW/OyGJCxTY14ugEkgqZlD3M8m4AQRNcuh6/0YmvOpbhvPEvtZ9XX00Pzjy
FCndNqUMMXPzmPSIQk43XzRqsDIWWxaaJn7MnuJw2sV8IcT16XGac4orDlDq+B74
LvhSZ3ZjQ0i6LN3lhNIMB9huC2CnOLE3Yt+q4+tZmycAEm9gzNYb3DvRkgxVgCtj
DZonp1Szp5srEAGpfmP/Ycllvq9AmCo0hDwd6AxXveqxOKZNRk2vpeYybR6is8Z+
FxN5tHzGp2Kg0URoEs4KgdTI5XhTGv+qCtd1d11akoxLKUq/pPIbHx6MPfZWqcnY
jTEsrjdyaElB16IF7UgR8N7PtoR6AbAehWcywN+Y+YmV/dr9Fpf8Fd+TIGeNB0GL
7+eCST8ua/LJSeeC0VdURM6NGHQW4zp1mUjLcGoYAE+/q6u8fdJpc7JiNKidrhb6
j2mq5qnc4L5RGBUCGwMjHutAXtdWxbW+DaEC5NogxN5jlND3O4ZxGLngizCDuxjy
BY7s3tgaVPn8BC39R5IX6BRmNWRg2V76Xi5Kk7OTDPq5cKWVd/8F3gHcy32pqfhY
nyrSZWPQC9fVz3q7KJAO9E4msO5OGYgDMsWyvjTIEGd0mkO9BiZcEKbl51Z5osW5
jMO8sTctQ+S8ztKnfv0yA4yN0W9roJk0jFeBPoCEfbN+ePSO/SrbcbYtVSCJF30w
kHc81ZJOCl6rRHMcyW8uM1IN2RtNyYB4ilkilfN6i/PemJ8wehWtV8w47jxjybEN
33Gq586MKzAbPkHW9hZLze5Gt+eT4b51XPF+w0gS/60xGVVtfLnNeELuHt74WTYh
iJ9GDw8LNAXfJCzlbNJE+JvleWDuXz73OmFCYAAQwSI5l9N5ad+u5iD3TLb81tgA
5ARq0+stN82R/MA/ZhQmXlU62UR8MWkYUB0DwuRfV2QQT9NDLTasrVbhUwKH8xc7
i4IgLHwwR4rXL/wBT2So6XYey5pRQuDQnolptiXrmZwK5cJeCa84GzzVsbqMwp2c
xqnvg5b1Po/fiOcFbkw1r1XWo5wWtbI43h4amgPrEMfvclo2Yd/61yrbVTOZhJEf
8etHFw1D5//1D+kc/JL3L3BMZIcw+lRVUSO5zjxc9uMxDNdPCyR24AlWh2aXwCmB
z842oFai2i3EofBkO3aGz+n8ddScp+yk75lffhcyLTJxiYneiUDEX4jlncQReccn
tw8uaQtBHUOxCe2zPqkrd9s4UoIFKrAG/O8tYXQtvo72TDn5XqLmRGq2eSOfCIqu
3talNTrDsLouJwGods576UQHO/mlFIsjxxO1EPhHCprwluYD2GZxGWTVaMy1UIYz
kwb2lagrhK6/URe4TeT4/IaJi59HXcUpxjwQT+I4qeFm7gn1mJ7eh59zV2tP5OX3
z96t5WiDxmnCP45wZl902nDgSliC9BpH9o+rkDSZDLV4qdxJB8QS5A+CLBfW6IiK
j2MAGX6SP2lybnCftjrKX6zNZrs56FRswnomOCsU5LmqdAe1t8FikGXAEAj/Zupl
0X3UhBU+1vE/YADQUuWpQHwAnhtREF2QbcQ1DYic2FnuKwGslYli8u9+ZVnX7C2+
E/kBC0q/mhGD7Dn7XWej8M1UUjCzJb+SKW/tvUvypqhQ4zN1htWgq0uFp4PRXO/D
+6UbhABQtanPl7V8tSJlLfFF4jTbRaL9t9npHUI1Iw9o7JIcCngWQIORBDhdO4o4
5yVbQ91E1Tlke86qKqISzXgbWDIyLfBUHTmI7AMdCv7wqvQkMpb4bL2wjarhuhwq
BKwQAsTzMrw00Pg4nx/WXkTgWoIBNRYlCy3Bjl3G376uLyHKW0lWO9CnAkW4ANB8
5nO9BvbM7F/Y0HJdj1UEJEcwVHz6EKTZtS49Eby1tGVClaHazl7YmPnickgGVp8+
mNjm0DPmSwA7b/esD4ZDSY36XCIl2yqK3PZHCArFQnEKWCvraveQjjisUG/VKDRZ
Q61S7YgSo/2L8fKg0h+nTp186Zwwyan04xuYJOigc8NCrlyraPtFEX258uhyhzYK
2iQJW2z/5rtxWST42OF89ZELK2vr7dhRdUXfu6m7dUyVFZ7GvirPxhfTjNm202nA
tV1kZe8cBY+JazIpL5q5mzpUGxLaTXJdinepLO+1zFsTelYaAEuTMwfq/wzXV2Rs
sdVDHCi1vu4JNPhjbRAVnRWoxerDjuBPPWE08IuwiR3kITiwTxHrhEe9v0ZV8UfJ
ccMlNBV9BVYZrsGi8EOXmQF02J8BbI5Ss+L+N6AoZnCxTFXS3X+aaBEiZao3mV3c
XhHzspNaaxMk0p84mR8d2CvecL5j2suK6G/CFO/V1E+k7FGjcOZAwDbjwYsbRKS6
of8lG8RRits+hU7NpTaaPEk1U4PrA06G6ZeuPkeGVo60f8KAhKV/D1zAiLVknF1Z
J10nL9qGr9DSRvOI7VuazWnwm08qnheS43jA9qW4v0Loq3nGdMO5wjTKPJHGkTej
eRq+iZl6Ht0QWJ2W9DQTL1hGu9Wa0Grtj7ko8OkctGKO18DkFhr1YvltBHG3J3l9
PwJT45Fng4j2MkB/jwZu33MvlbdVa/sxkWUplmZ1klSPeCdyxhHcFDvjMxYUkIo4
PSXnX2+w3ks7PpbwcAT2LU3pB0IsxPsx8mEUfLAwYrGRpVdacSa3Wga4sw2/MEfJ
cvTz7A1/lEh64qYel7HIXb/8CmljVpUkoslA9lYi9AnGkuxq4ie6YyDodx4cLNsJ
PCj4hKj1AFvhk96/ALZwJuGC24vil/fRH8u6ESBEszCbivBjI8D0kX0WHqnafvCj
wyC5Yws9oZ7zo6GTqoQI4rRKqufT+iQ1R+zo46A4xhO2NPA0zzB3dIHEFlaA6NMw
2orUetTaEsQNh8oLVHn25yV4yCuo/cGGOU9vilTGsf1D3b6jje/ukGXvIZ6ze5jY
1omEguGtzjgDmLqLT9jrpx06REprq0QGmSDOxPev2CZ6fUskmlybAg9fhAXksfzK
r4mEjrrnmyCbrwkp6d0Qecg4MCcF2ME+Wdx6SsXy1ns6+ZdWgI4HD/ZbRUOl3Z2a
bOZYVfefGocmqZzLJr9lJOf8/tHR03T7sDFx7RUYZmppvjNUndBfBM/6aX3q7OuZ
XnG2ek9KQS490kWXQo74E03ZpAiA/vKeRUF7g8gp5LQs+M7JhPYbtG9zT8g9U0d2
xt+P4aiqOL6FiryOYRH+Zwt/O3lWdYLsPrsm3AJ8OANmsqSxN90DS7sTK2Wd5Ayu
CNKoz9NtxxDRgfyz8dAaR2GueEBFSsv8O280tyDkX2GkRS3ux19h7/NCywDEmz05
AeC1YN2AubQQdh5s/YbF8aSn7VR8ZttWERVAkKdhUcEFgW4nX9zbH8ws3J+avFns
KgaTjIVBnDEw+ka/M3OnGWrqtkwncvGMWItvXl6G/eaMV2xTe8G2mrHv4/Q9+R/e
gIEAlcUlNIfBJUp8J5/nXV+0hvaFBxms2CVmywlm8/dCTe3WXQZv3a1485GWOK1z
22fRQ5hyIa50sStRJ0Irx9uelsgvfiZgMtR5YYaD/Ud8LbDnTvvNWar7YHHPQw4c
PYmd3FpNRLM/aHpy+dtunOjscTpp93Ss/UdjV6HjLluFKkTjK94vuuV14FAQhpQp
Wajj1YaptlWCQsqzEqufPd00Qd3r1BRf+CmcbMEy1WPpNmt4V/pXyAdHsUG2k/eh
rHqDvJX1BDqD8HoL2PcP6NhM6nEVrKelJZhRMkjoc2G7kCje+eTRmV8kA3a9dJRL
4oHKvsaheJpbdD2KmC3VsRUd7ATCLhKc7m8E2/qAJKss7vE9t0f4YK+OH8ZWrJwh
x3aqbSJm/BMCkPeMcVmdMdpskrcRpERM63i5TkHpQyu0M/rYML86HTFhg8p4t2Vq
M6n6ddjNPYSE5w/4Qp5C2d/fSIr5G7WTO0R5xhhgHk/QM0SdkbyZFsZk+yK1+pTv
W7vJardg5WUKu3f0PWsM1lnAgDYkpc6dEPPrf6rwekzMsGMT1pmq41eyHs3LT+k9
W5SHPec1Ti65HTHYtw0jiNv3wQL9XwvnvCJ7kKFZkBWz3IQoYRG/L8qjhukR86Na
41VyjFbx9CUZodsFsfsSw0pk03X4pSq7HhMzhxvR44lzX3UO6j6jekbTnl6q9nz8
nejRKQFhS4bAPxTWdK4Vuk9dYedtaePjdYmPiK/NubeY6tszmmDXMQAci4NEKhwV
f2SffxaSY76wGf2kmDOl/8jI8CIADeJ9JxrciPaq0F6C4T9mDsreffqnQll5htCL
sVxNiJqP8bZHGRjFYE0+CbXflfQTQWCaDYseA1PphGpALAD/Fgos6TU4aTt3xjQa
Qkx3BHiJrGr/s2TRKWxP2YbiH7PTut9aCUrmf6f8tXkfqvgD3v29gStTrxz1oIAM
7OwgsQIYsVq21ZuPORHo1a9H/FlqNdlIjhsxfHQIHV3NW5MTDYmoU4i08EVZq2hr
DfOQHugwPXKsX/SU/JUqsgC3P1hvoVc2t8xz5Khx53z4fokfBobgF3Jh4a/8r7A+
Otj56iHYM22Lh7Z5i4tssO29+tIYDdKtqzxWHEfAco0G0kMsbruua/jGORZInYjv
5RkowCBS2hbVpEibnuzJE7yd+sGNsPTXpvqHNf7ku6DEFIPDzYi1VLH49SOpSdjl
WTan4+H7zihUzeRKjK4MAnaoS3ZlYoXCIMh7neNc7fhGlkHu1291YMW6Bap6M9sK
8PJ2kaH0gQL3Qa6E9wRoe3A4QWXGss/8o4FrvqwEa6xcnLDRNmr4rT7ILn/aNjQm
BE/MsN+qBIZEP/nD4eNv0GG8vfIjoemMt0U3sdB7yJse6hVXjN8W4/M7UTI+dWNB
IlmstvcmhIyjhmjEb5+f71aRrVt/ZTcRZYaQmocG2iqD0btCvSfT52q4VSEja0ab
yUr4e5UvoaPCLJX3cuo1+yxabBD1K5HEWT8+zTqzTIh1SLBfcZjei4O8qC3raoJ0
A3ksWV1quceTKmjCh4GiXuOv9qT/LKBt6O7CyRPkRLcU6HWV/+dYviVeulg0w9Ab
CHpsOUGhyXii1CAyWRAAWpAfYak4768EnvU0gptJjJT0T1KUVdZ/HdJxLQGiobWy
gX+k353yPKPE7S1/KFuc/KIQ+SlSc+v7e21Y66EzhQh6R9IcLo4nRSrSDVpThV+a
q31fbgRzkTtXShAl4DFxgkXS/AzLG6zWeKo/VwmUWhIBa8Dd2pCM4PbYIevc0Lvz
pGEpzH2Z6Rist/d86pvTSxKROmCaN6g0eXkQzwm1s/xRloEZIZ2Gn8Zg5jcLQbCV
G5DMUmI4FXFpLn5huOO7hv5QA4zv7lmbHOxnhDJ32DbtOPO67UmbNsS0zWP93c4k
QMFfHnC7BslT2TNtCIlmPc6TlfTfXHZ5uVz9uIe/O5Hjxq+DxV2wJqt1FTq8yEuF
QfKxWNIWj5XLdui1FbQdPi/O9i+jVCcFPx/QZlgjQK54TVVsRZlQIlXwnwkT6tty
HQaFrfP0rMoUCk8sM/1N6AW0yHS/d3OX/KaLM0G+KgwLpaPwILCGyIwvCfyoBTtZ
6Tr18+2hhq8lbPuIYKmJe2z6wsrxEX6NAhVijfHfs+kpoBZXm0G7tmxs7xKY/jTT
pLbaVHYIIcnT7c+D/9K6yJFlE4RGAcxVo5Ur49odlgDME6xVA74K66SZULDzvmNv
+Ju9FiAaBwWsnLuFnUqYumfokUTjBjANtHXtKWGtvQF/aKIAkGBudPxG8b9VqIog
5OpIb/M/9p39O0UNa0hDdp6kG3RnEb+6CudCRZaahx0vI6t9B4coSTssli7zF35w
q/5rSC+88sIQbcyZgN3zNZhYjyMhJj+CZcqLO8JVvqq/XaJh3OvRoJPYPG+Ncjos
p67KpBCp0zxwS8GWV0tpJOZQ6JG1fTnYnTLyHpS+wxBW0ZjepWtxQZQ/V7UGUTGM
g9EE1mPh0U768zt1PUPTxvTfsJGnWrpzrqYfOV+W1lqDv1rui9naPDtf8WX1MdD7
k7DGHh73ha9d86tVywQUOJOVo6TB+Pg46KH9MHANRt0Z2BJfrvyoWD0tqzia4qLX
jVyV4+XZ3dZvMLS0vtpGLgkdfpvilXDxCKqKVtBrVili/vS5uwsN/MRkepXZuabW
wAODhw2G/tHskzYAiPZdleEXyqnkbXnEbtd2X97SpTOmOWlxWgAeMKM2uCHGAsK1
/E+865dLyHnf7HkRiYyRMOhp6D3IMAZwNUJ5e6xSomsBSExEbXxz1++nq/3XkiDP
eaaE1z4CMQjw3tEN1MeO5ogDzpj2A0CFPTM51TSLZ2CxSPjsqpDaiHqnsN81IzIQ
ZL+Pqe3mWqstq07OTDv3sq0uJ86jU0seEFkceGFUbHeKM60ttfw3rIO3vgZ/gC1e
8pD9ZQvdpG2XYBRuJGdGGOGAVi1OeaxjZFQEqFb/FwY1O0BUO3Dbu6iiCxBBO3N2
D/Krr3G46OUHGJ871bzBDFeNVbC0FH8kEsOYVUzZTaWqg8KMHX1H87kNcqGDPfna
/yhjPgmFiEKlfhNMpbeOwejQvuO5oBJWMlZeG4xkofBNtcObHmHdNq63HF1W2Ei5
trxqJJrZG+PppXcIgBKumMMPiw0zHVP+tt/xIZQ7z5IXAhK+uTzmriA8M2WnHC5B
BiRBVQczea0BoIYAaSfPJWQycU4CHYj45HpxrWlnY7ML3GQ5EtaP9+2ag7DJyneH
NfRymDCwUhIS99dIxjRtTzveCiIojDU0dDYAxUpGbFZ00CaWN0ExVaLZ3FZM0W1V
s9iAXu7OukN1OJ3tc2x6c+UxQu8yTpWGYXJLLDm7/A4r1zhDAwlaAQinKvS8WOq+
FusX5Q39HEKKFiQsPrqqfZBwDQYLu3yuwmzcZ+j6F1HbWmUebyGkSIbJJozIN3Ev
LNIGoj/7iFaOV4WFVuNPvpzPjBzqX3Z62KRJVU5ec08riugYwDQjLy8RrdWF6XYx
0F0qEfdpnS82kA91M8RWDQYIQFCEA0rws7aMwWni6T7s7csFPvdzowIhM6crR+yj
Zx9y54Kvqui1SA6DOkxEXtE4/lJ3TUoz1WV0emWky/I1i+AyXEQbraQz0rjUSZP3
Bre0mCDCEAam7OKwMYqxB37ybIv/lmD6V5O6Q+BddvablF44kZqTd5um1TWpTdhT
tmibzN47dhpSOPqWQAPVQMuAldEJy8GrMazfDIwooMG1KIp7FPUmPcI3Vvnl80Xz
5CpXtYtqFiVaPKzk1XxeELwmNh+sCdfq09O2tpLBfy2IVlZQ+NNJ5MOz271MumeK
bjDrG7gjxm9ETG8ajHjNMPbYjvBQOMYj+es+sDEsU7AsuNRp8oUGytB2fzWWfzJI
Adf40RKpCZ3hVZ88JExXfSRswxuuSML0/RzwkDF7QJ42Q0pMxopBK32217yrmcDJ
qMUzIRw1+Ej3GdqfFxUltfYkViufv5Y3o+JgIR+/5+9QJrYkMGTGFJVuTDhtlbD1
rUKwBldOBG0OoHp2L3tBzz9cJpkINgkOKQTdBaWKY7w0GIl55H9BX59CnpsYUPOD
F0nPesbGQKjLEJD+ivfAf4VzTAaxR5i32yKm6vg5kzBk3TUzPUDtA1LgsyyhjbXM
4bMl3/0wagAD70LMH4CTNlolAM+0UaAHhpM9GNhTjfSnScNU4513KFY9EWSNZCIx
+qJCyv6mn/bnbxGthJaxomeBtS9zETOPDrwYLDKG6NTiDUI/zSyth1WzF7M/i7R1
0sLDpYqlXRUmSRylTNvAW2UrdOwu+RAiKPKAQDhwxR4FkIiX03EfJCjUA4OATkSS
WL8XKJOJnFo+1p1RVRTbCh9DmXG/2CogZj6VYbSuXJI6xoWt99ZqGzZvvf63Fe6U
C+NwIU2RfwBi45omqX5r85fOk7pa7E1SsD+X2UBeNjjY8Ns2vJ5b8SSfZhiBHV9s
NMY1fOcC6zXx66G6+CGpS/Y48LrbXp3c6cpP1ykeckM+HLXkwgTEyu+poTQkaxGX
DKh6OQ2zpYlMv3rHLeDi4ySmR380P36/bH7WlIUxMTjfGsiOOge5ifXVs7dF7bO4
6utDdYj9KZnxNxCBE+KWP1hrjfITy5TSVKjbjUD7yfe4ysVwM/MzaptSAgUp4IDC
jg0pYZxhcGkm305lwAuj79/ZHn5IJSavJVBHaZIiGDrCAl75paozAZEw1NhGxIfy
xaGz0uM25tmCWghFGSJ/h83wCnZqku+FOLWb++nfJFmhFGr1RxJhQI25hrrSicRC
bL0lNtSAmackPWUAwkIpH4Vqa2EAokLNE//3tMcrEHMV7doA2D4sRNxsR4uqZCnX
xzZPsx5A+m/unHO0hleG/B8FzrNfWt/2d0IeQkfsD2hs3NW7O2uFo2hBdfrltluf
J4hElgeLnV6VNSkPV3Si66UPA9h+r46YIbQLeLm0zmCn3PwAqqOzarjJOcYjsygP
Uut6KkU/lq9yyufmALCpoQl9+bCtWELFg141dGVZPmPaGvMgoHyyUKtezOxeemxH
mFk6TDLq/jWpOKpaQEKSlgXcMxELgbC2J6sqpsT/IrrLPgjIPJHML5p3IouJZm9M
bM4A5KLarJXH3b5GqZ7wY0HaUtejVlc3F+uMxbunqOLhVrxMwkbyYIF4+uHToQAd
HVAlCHXKkFfbsJZnVJBUPoEDMpo1BnelaZVJ7JAr31ECa/VGVWYTSQ9NNZcAhA39
RZye6uilNRNLTpbXbnkbw0TRpR+uwUE9bOz/4J+79qul/NioOfzat2aQkno2vRrp
GuaZ3z82eqhmJB0Fr1Iua5CMreniUl+2GCdZmQAvQDkhrJ3R5VvadbyvIvNQm9u5
DVNZDHavqEctL7LIJxY470bAGf5WVKm5kdKXPwQcNRsvIyRP8KxDDIRN6FvxpRRD
OaXJd/V63mU3PXa8hNKcoIDq0CjafHjZ1kmXdLURL91GmjrSWAsLCx2/XUgLsV3u
Pv4VO0At6J56Y6HxcMTLJk8NwnNtzgOTActcALFbP/+Awk0z5Rf/u9oaICkRgtbt
MuzkA9U7bOzC1q7FaOhVgNhYLuv0Kck+vFqQDG9njvbrRwTHiP1bsfMEZnd+SRNy
+ltDTVA7jUnJSDdz73NIOUoDvtXr2LBFuUxLpj8TlqSatwiQNQeDgkFWC2MV7U/U
emeaeEzfTWOQr81vzYQQk5YlaWjer+ex0yAmA7/WeVbNppxICkYNapeP+7v8PFNl
K3nohZYvjp9XxVJcAkcthqNCcRmcob7RryBFEiRyScM0jM44j3XZ9Sw26KiymyfS
bDJccq3Xt0x1kFzOIGAozVOmbQUsngE6Cd4QK3WHmyDQioL+3TuBeRHN6uYImq9q
/ZUxKJkp9PqGkQ630KtgmIUkpsrCFjFWCrzVe3vXw/DhNGdxeCFtbsqzMF33e3uQ
9DONVRFj4DmeFUUl1zf4oz9+MQX/odDHItqGbiEUclLt5Vqgzs+jUrjbVxNjRytD
tpV6FVYnn358EMHYJDbytXbl+hHLMo+djSVKU1/oM6BOjvvrpJWJN9LpsmBgzOg4
2sQe9+bWlVS3MEUrvx8lySr31Yc9c1hqJcONFUNE/HpmudmogG2sx/GTWAIaN7fc
srj2/fael18hf9bhhdxOYSGWp/u4+/5tDTLUWofmgBFzboeOGVZ6BjmAadDD73jK
7kWq2Q+4p5eSEP2DsS5e4oCoqNwiURLbvWDWNAxh2HQlLzLbPPqIlOxD1ggzrtrZ
hOwkU2uunHzEJoj65LndbyRedjxoKcbm8pCikBQT86KP83YQJwbMa3hQ4W42x7Td
UkN8+5Z0cUoMiB1051TYTCg4EmXjCGqQ+r6tjgZiQogXr5C7YXrzqXm4BbBrsL6+
TXbR7yFRvZEattJHWK8uWgzWBvHkDT3hUMI1Kd4yMFViD7xCkGHS6SEBYtaR/0tX
4cd6CTWGBEnRqgwWzrYf3vm/HIyvjNPXXDEmae5T7ijqFrZ49ePbaGASbtCnqaRa
a+1WGglBiXDH+KgKRY9R1UKbrB4n94vHr82GyX4hKH+C4bvYyVahQQzVZp0QIA+4
YjfgqMj2UibSqECP1/XZ9w6LvdX+4P8TXVR1ajB/g+0T9ZxL0yGM/d3s9V8+1s0M
DJEwQYtioEI81hOoAD08RVZAHWPWoYJ8UKPCl6u+aDnLRTmmpU0oy+O3ltG3vVYA
eSNFP89B41yEVsAiEz5sPyhzbK0xF/+/tKt1Ztu04Afggf7dpq9+BcruNFWhf9gL
qFjeYge17rKnGtnReK58/1y9wDuYyOsFbusgTKo+cgsKnndkWkfQJK0/8yP6rYGs
4glJSHkRQ0J1cHcGfSAGIp81CENBWCdWxXiA9hkVO7mxlSyG3eif+cvQYyJkKKW7
WBizdaU5YgJaoB78K6H897BJJCaIOj955VtQcsQHnYt/6sGlR24SOK4F/OHHUzlV
51IM29gWar8mJL2k8kPL/Su9tE+fYWwHrpC+YPiZ+R3CkMW04dxoSXx6tigRpqrR
DnfD6gQZmpfUsnA6JRYxtSjkC8puIg6Pnpcug23pOqypHSVF1hDMDQcG1clsPTiH
J8i120xi6qzyN9FF1Bcr9QxXXJraIXDDreMRHANE/QxQO34pYjD5ZgFVExjNhHBj
wDPOrHmVUyUkTb718Sb3lN21JR8wadcQMPlaqNyO6MFe0e4g96URScevjDNvRYYJ
n6WUJ5/6lYEy+AF2Ok8d4tKixscIao48YTbNrk47PG7LnhvT+XZmcb3rsDkNnNs8
IRB9sgDwWjzp6nvyFXglibbIj/IZkW3XiID0+JJqTG72ENGzN5hnCZo5VmPnslI7
160pi6Epa+ZIsDlUcFOrGxhbg7ez/uBIfPBFyTqhwS4uFDSmptEVNLABIkU5SUy3
WC9GtCSOjip1KWU9Hsd24kg0fsUZjH0xjc8n/s/E9JABMRkQ+UPgJG2Vd+1pKfyp
I8yyUWZypby05Q1KFeMWUVOQyZKBoEMW19yVr18F8W+1NPvTnszD85UTWIDHAd03
5qLQLC7biC3soFvPKieQ10Bhb/OfIPac0gqZVDbchk6fk7n0fTUDghSO+oMdzofP
HxtmIFn5F6PKINeObBW1ya14VUDkcfsa263pHc1EUwUQBi7DRx+7wHNykWyLDiEJ
3OQVZh7QTH5IlUVJsIQuP/cw505v0iOHL53+/WKcHXPFCrHJlm6jZe9c+Qu1kt9X
f6mYbbIjwlpVnp/KfaKbDAB3pbb+0g0ribA1+xfZDEfvHAvGCBuFVZNdCvzHXACp
YL3Fq4LhZlVu6ZGa1LFqYFPRypj/wVK4Djucox/3JndOltvAVqgukjQ7vJ83cxV6
Aia2RDuk1E3fM2TUZRpAI2rkDPAL5UPl9eE0edlHZIQB13z6vIdGvTU2hUvYQbWJ
ATxB7RheHaWTJy7hkp90S0pSGr9RQatq/iP4XoKV1QSKf7JwvaBjPmfEmyl0cXxr
aYJDDCQnkzs0ULJnFjXQ/ZSiixXEAtpx518POWUnaSkb2XIprV/VKDkKDx2X1Xg8
rX/LUv4EEFeWhLUnWj5F6pE6sFPxvAfhaCU9IepHave0jXEy6OlQKH2fBAiEZwKY
nOWx22Z3ST6EJI7ROK7gD3T8O5Sjf3pL5vDMIE+EB8pCUe0NUnGBP1dd56/hdQ8z
XBqzPjaAe9b2OEtp9/zznyouTQJbe2btLqOqjXxrSUNK3D1qqIlKODsuwlUTzZlJ
iRr355jugsuFDBg5hnvfzE5RMoSo0saPplStcC3avW3SGB/uOtrRV4+JUIKQpG2C
1fana+8f4r4RMsRTE3vDeAU+gW9zL3yGE6yUUC+2HjMHolIs9MFoA0O2IGLQ/2fO
2uYWgLjvUBq5wqIUF9iRiLcxVQR9+Pkri7MmD++oOOZMA/UFXg+Snw/VSuUYrnZJ
nHFJyVIS3agwzy+gd/VHHMlIkejO860ePoRsdctpZDG58KBgUqdVoTrFCT2csxVH
ntOSkB89jo5dmMBeO0fItXa0819FnN+4MazLRhQnzngofiT9JU7jAENEWzGfiMeH
v8YhQIwqABbUybaU+lgrIu2heSp6F+tkREOJuMJvuRnHyCw8FT5wd6KDsdtSOI7v
YTz1DtyLHm2busqUYjx0mwWUFRkx5QXMAZamLHUMXFGAoHOQYRi22DA9tdLkyhMq
3EnW4B0rEPiHgzcQoSr5kZ2rVHtHKDgTgM7clmYghwcpso+aP8phkk5f71n2JusS
ejU/rWy7GdYja34IYZIjoynEbMRW5VNh7gQKczLdvkO6TYm5AiF1KCDf1w4csVJ7
UNMgxCig0ohDecShNj0Tgf6w3P0M0rdlt2OEk9zZ85qe+/ayyeKw/Grnk/K5shoc
/Ef9TBeB1MrY94dZ9MYPSsJ61Qjuex4Bo2j6k160QiBJowLIlV4T1MN23T8JOvBO
N/KHpdaL6MgrRAw4gCUtaBadDLtlBVCa4UYkEj454YegADxHxAUX+akE7BYar2Xi
GSW1MNi8nqfBdIl723LTErmExF1g30ay/kCAwblzpnJjBrlPExnEcSmZfEBAMrCE
vlEeck/zjpf65PJvYS3T6m8nxuU7MLVye1dmFdd7j8u/Z6S5uQ1GfD2biF8fSmVm
EhRhMKOyQz6toxi19OvCH2dXp39Gvjgk2CC+NXEM1ZHxCM/VtI/p2nv64REVe9ke
gS2dnCHnpdT/48QcTIpS5sTp3qHN1F4m8f7gUlqmdY2jePu4RTHN+ekmT7FEOOLy
100roCKodVM33Detie+ZkWVkybSlsGHJLmZpoJ6i6TWiNzFHrKllORZL4q1edZu3
Y6aOcm0VIJhlSByYchaMPekcP1VCetuHYxLUH+sooSC8gSuOsNQ5ecn1ihE6K/0R
TlAJV10h4Hwn3+Vp/6sI6wnbeRbQmMnR6LD7Zg4ZNbFuiWNlF82Sd2UGt0f9J5pp
OwycAIugUYcuG+pvb2S+JiT2C6vdGbCMa5jgu8oQZB6VzxhSuyVOhkgUsm7gKG3+
31QWaEbDrFuLjGL5SbGa4RScVQftTIGDT8FImRmNu7+x2sftvldiSun3Z41kPZqn
8MjO1hCUzkHsHz4NGhRPCRuZ6Q11WpcCfeDUpnMYgGsU00HippdXVM3vDdL5K164
Hug72yq74qj/MMCponGpn1OpAhuiEKdx0ooTBw3Ix+97Pic8VZ87jxjD+rd7TQJG
Tx1wawDkW00YKT00i/3HpsjSa/b4AAkLDHSa2pymrHMLTPPpZqEc/1y+W/UR1Pcq
beCjNBYWnrHZzfwAHLinmMHxvIVtl/dwWA7/gtm3TCnG8RtC3zUbcNDMQK2LKwPO
1+7O8MGhzOJ4bXc1t+JoYhujA29j5isTnIZs8eY/P6/NL2Nv0NxiVK362bsXV++i
26pyN3SD2bCnYTZr8UcPBY43UOoTj8zpT45/uOP2Ixksa/kg1GT76g0QFpx6jpqt
5umQ7h/T0ZZFbym22a2HxPBJkHEl6o3tkaK8KdBXIk+kGQjPMMBMmEhNEs6zkwWL
qeJdsD+TSPAzWSNwZKhKL5upOaktnmvhc6gE/LDis0IUc8bAm4NwFLgMaBCfXThE
WKRpzVJuQ4KYd9GNwrUMXaLNa78xzUgHUwuAJaEbbuwijeajWcf9g9Vt9SALt3wL
UKJd/2M7q3NZFcFLAMxHZuTPfCSP8BprE+ypQs6XxpsF7i0rVfs5L1YGm+pFCG7L
plZYRuMP9e7qffOt0gs1xNUbce/c2ahkc5IiZM9Z9K0LC3KZ41WG2AqctvjsogMu
1qMeAEo9ad87nkRRr/rCu5qjR0wf9XWxOah4nBHIZhV8oM80AaGS055GwSTyldfV
Lg0wRY8Z89WY+yf8p6Z8JzYB+097pZ+YZJiJeOcxi0QqKieIvDd8fTmKP6SxLNX9
eGHS3dU1dGlut9fVdr9fR+tIOs4smn91Im6N3AUHPpUP5imvATaL6EGUpyRQsJsx
ei6iqSZ/lDwq58+t38VIITxFGfINX2S0Sd+aOriwN9GIom6R9Bxkjxb/anekVlaT
wuYoQuib28zT07t41ztfqkjozlmfvsiawoDLkzap1a2x2841ctP3n6REK26HEQYr
EYB5uR4eRwRnK+xFPzBLbGkkDxhtbGsc191plPeu2oP9ErZKYoKus8W7FAahu3OG
fD0R9hfU0q4cThZ6oNvEieQB6m15Jjfi5CVaMR2JaT+UUbT+roiJ+MVizvLP6jN9
YNNq3MWG6j4N1nx1mwu9P8UCVRPQWsuF4euFuzpUpDRtIPMcbanA+KdRFZgEShnH
G2seljyx1Fm49HfmCOdqOlkMnfWzZ4OmqoodqQU2Xzgv4Jl78PznPiGs8ZIMJ9uW
u28rpcW3yhW8LP6+79G/hdj1ekZML0BoIipMxSGkeVzp/O09onqKs8T9fqE9sgsf
0kuEzXwzVQNTjZrinXRhQNy1FWoooJWqm3qlSsDpvGYF7aRc3ACFvoarEQOmY/4I
i6sDjenn9zyLM/q84urtf7nfcovmjQwetGnTszOxtDGU3wXhfo0FTDlin0H21Av+
7kvGH/pJmgocpSA72lDqmdgI1uzCc8E9r5HJ7hdJV2XUzH03dhvbs+d88X9OZWFC
PKCXDFjWNBESWOY8Y3LkXdh4IMcZczjNqvR8aMpvehO1rjADJe6Y3OxcjXHVqhbs
dOtEHqbGteWTxs/XNMMJpM5j3ipXK8zwKsqCKX9vt8dbcBKdCH3woFxbUAm81A2h
LjBjraxs+znzRYTAaFjU446mlwovRDtLik9b7pUbzFJ/U+nhZ5bl3HgczJUNiE45
kVJABItF/ZgeltvXFW0bHsASBh6eZnDHAju/XHI/Gu+U6Mc5IWbr+nqh6XSU+J6B
uig9Ln1j1CXI4IHeZ6pjNbCdn7WEc88SLgOIOFmZTstD6ULhtnZm2JPBRRI8/hRX
nYU+1TrFkyyFi+evg1p+ptmt1W+pDPTusaIgnK2PbmiOb4rF2OiaXOUwfKDaJCg1
HuCoOwVkfEGNYcqbeDsz4cnTjgAMC1Ibxkiu2KG0oohYGApCW1PXe+attJAqDeyB
uTcxaOgKHG7tYLu1BAyBJ43Fo1ejE0KnjNfFQaKQc/ygpIk6kEnOPbwawKZb/sga
bCwQFjS4iEn8Ue6mswJk913hc1WKSwLp7+xVRXMNNefzw5xlYYScfeaq1D2SN43V
SsotRGeZXyS6BWpjwoJaXxx8D8QKRHTGnR8OyzTUHIg7j9qGwYXFijm3TDF4X6rI
ScL4cRKcqGEDe59hSJWs/GhQjc6RJMHGe0tBt6DaC1g+cH2iPIoomOydr6RfFtDz
F/l9wQDq+sOoxN5uB7bXR1L3JU43SOSw74T0SqTGUWv9zH3V6VkA+9onjZqijOdw
ttinzVDYby6bT1dcMif37olRc0f50BEEISxFJMYK5oEibc7e/UIpqZuXMGi8AOJm
kij+lHGLmJxTUZjPxoHMdIZXD9oiZ6BS626uDC85bJg5C9uOqX4YYYh7zfOs0sPx
AumNtpSE+srKA8fJvWYe7KksiE+zrCAtBKf67J7bAChSY52tVeWx904QbmYkJKiY
8Kp2q9KSY0Mk+zlFqlFUoPMi7211p3V4oS8regZJEU12MoPtmZlWZ/juVZ9ULKr6
jvoTy2VXj7IgWuij6RP7+z03wtPVVrbNsb2KTHNHSgnJluK/87zIweIYF4979y0X
CWD5nVxq3S3HEJUgHW3CFUROE7e3O/ltoliOXYmn2QmMIHXVgpu6g+wtmZTyDdtW
BuRXAb9nNOsV15ovLSYnM3c4N32VXx+ToiDJ/ywAaYgOpLWjq4h3bNbiAAuqPu+j
ulCkabc1u8n/6Gj9FbZ8ozDa0m1Pv3TAnxK9rtWFxzZyjsLBEnZ0R4afZwTpqHOv
hhOAMRnqf6jzN8DM52CTQr1mH1RSBViIsQPsrkW9LngfvDkEh24A35vDhiCEihTK
m61vB21DOczuxY4+10uI8yiYtdSxn8rSk/tP7pnvS4cHTrqOzIelaGDXMMvGXyod
T573HXGU33/d0pEkXbXtiwu4N17fvyEvE2pliFs9Lhsgmm7G692vEnR441c8khRQ
W3QTP8zee+wyLrYt8AOq8G7QfTp+Hz24bxd9KM0XN/gOGMUhrqCY1Bo4XntWYs88
LOCeMvfrwJMNWAJN2alI0MqJd3iLjXJ7GM7AGm9hgLsVhdEpg9EtM3+7L7weHC/s
aYXawWOD0fzttHmlLMu8FksHwC4ux1qfTD2slOtXDOWIVJ1XkY8nPzh8YZaBNNK9
PV1n89QL/DxLCbf1XwqAt5/JS0sDhaDQ4zBFJGzZBMdaEmoM0agyR4uskCQJ+KJH
kPS22mwOEWfT7ZgtlPqcV56c4/DK9NAfK3yiR4NyltfdOkWcGaVsCYulUIey3Xmp
FjMMdizb+UjEXxtlHsPXBo4nW1tPN2wGuygICji7vRW7eU/M9pztjzzlxyv2BGap
inwKDp1m+Qtl1xxopxXF7pG+4UALh1ES+C1QM7vn7vX9E2Bb+9ybcZcQbgJ46kKF
vre9XuDca6Jq6PjpmV+b944Mekr6P++avldcs6rvLvEoz6Fd5Li0wZsMuExy+ZJ0
ahAOp4rk7JriZidZfKFDxhub86TopNY/Uz5EIP3bDD9dbd2Zq0mYyh2PnPkaAjuy
88apLPkcTlQ1+PCRbpMBpcRG0/OsA5O7Y3cHFCgi7AgrLDztXia4Rs4ZEXOusjZt
AN2GGWjXV/0XTr+73U7ci3sEvy2pJhvkrVxkcj9bp/kGKbCGTACAPCZocEQR3XGx
gthmgaYEyHnOk+Mvsa/1kzFOWtJbPZo2ryKZXIWFiBqVgJOeKbIJlibdmTCDiSo7
+gtVUTvN0/nS3Wi8eTcMrCklRNYs8J0/NnB7Jqv/+G9idx/0olMdOeSZi9/XpKGc
8NYzHfG1mBEH/p6LKf9F8D+ybVJQEhWwJXCdQwQc3n1bAcD0PlnfSchKwImVF8MV
H61lCAHzSv/jIE4ovN8fOEjUCZHk8eqHN0lSUh7emzwYPzLI5EiwKswhNJsZrslc
pvUtAZLE5oPfZXKLqxkxurLTPFCaV2tXM2923xqo0JYSe7rxJAkWxw+cbiUHyH8p
X8DxD+T+AD4CTeAv7b20m4yQCNYJ5uiSHJRIbVlIQN4UcXCQ16Z5l8Sbcd3I6gP1
bdMa5Lso/hWH6/Of3rf+0SQ+WnOo4u1aeUTjk+NUeycyL5z3BWrz2sWIo9JTS1cM
dQI8aj1NvpqOTYl2Ng1qTjXaQBipuk2AstOyffHZbNj/Ns1MIryw/RzG30xDYgzm
pIIKL21R/xWKE0FFyrG8fRRwBszrfUSVsgecuuXtg1yv7DcBVh13SdLwSadooujF
ZdyziSPDCkoYY65sNU1/IrVreuE3fQRfhjf42pKc/XlPSfL8RMKJTSxJ6LuJfyBi
bJF7lyrRUKBeBykRi5ayR83HhDZ0dh05iXdMDOMKD0SBFHKd09DN6b1VBmDDsQxX
q/wvQqeS6qZ4yZ+mWhCcTJOIZ8L74uUP0PL8SE6LlBekMfjVMRF66LjIGz1H9Zfd
5R1+wwIWcdc8Z1HlT93Ho2CgjhCC8dJmodDQK1wwC+ad+ruv/qUnLdWKOThtjW0k
xMMKY3JuBARpIIFRZBjmFinWu9To46PmwJ5QmH3J1poOBVUoLp2tJWGFlALM3KiO
b1p+svZ2UedLPBNEjj5VZiIwpA8QZdi8Ctr3LdqC3gDlBLI3KKudSGpkD7vkAayA
WTPrPNu6XINsHuSJ9+mu4CHTppsuqC9lMiXnPaONi5kZMkg99PObebAhykXMPmvN
WhIHekoRCUVN77WChFM+6YV6xaF46x9MMWHoYRSwEeJudiWFX2ibZxEgagNhy1uE
6HRQdTpNmXEPXIu6ewneRTPtZdtM+djoYu979T37JhKtVmXgMPyRpK7NCDBmLIen
oO3WuezgnVKvSfQnRj5IAm6TDyGjv19V0qwZuzJO47yvbRFETzl1DDUTkfVUeLCk
+/QfJ/J7OWRCwJ+8drpvoQzSAWP51nPaT6MiGjzWYL0jE2NQhANsywFirASoCL0T
RapsQeN1dmbtuABP5QB/Sxv3V3An8Mj1oRME1iv/u5wW2iln2UNSJgKiNh0JLB5b
WgVqjGOjfDgNCsBtqDkLsP2m22p9V+qncjjpdtuz5dkgTk6V0AuTKutFi1T8hw/w
fI6QMdKffi1/GPWNZY1xAzb5MXhK+L0i+uIl+ezmCS2VvIABhB5wuTvlgt4Y4tpM
xOSiycUNNdFPesuOEL5vGu6CGOVF/s6ubQJwEcTi3r9Bk2r11IpfkGLbm8cRPXz8
N8L31m/bMfO3JHaoR9sH0szoO4Qf7UUOcVcUyXA4N3OqCrWz2Y0+ZRu3q7k9aSoU
YTKF+lu9xdDkowAtkGiE+Gt2hjk/RqxDP4z8PYS4QzyM5DcIvZrB7c5iI38Sfphe
Xe6IkNP3//jce0mJIy7BUP2KiKRwAbc2FAkyqXICrstxn4RQV8QQsSbj1joHtAV2
hezgwZNjITa9LF51v12zYIIcUBHBFoc0yM1T6alwgWWgAbOcqzUyWDXzXDkrirpr
Xg38EprEUFoNeiNZVNv7HzOsdcb+cwAYfyJgmjl+zWJ2Vo+lJl9aSlBrLkBsYdPB
XAvyqrttAS9hdaW0Es4d1VOesTLtk2jJTnDp3GaqGnmdX3dlCskeCGrDw+1XUmJC
M5JASjiKWzEDkMhsN1Y363xZ/ia8agU1nl/OiECbQsTekzjccPLZ/yWvDeo6wknu
IavjrpAqz2HMnFZeIxeq/ltBJu0/haaWmmYoXmQqQrFr7X8OGRguwydm2uAAjVkv
tzFTYTSi8e1TYJGHiFHfSen6rtIbD620auHseEOCHBSmUz6T/IqeVTNJhqt7gHTY
H5vrHdVcbs8TWynJ9tX6TnuniFanTWet+TY4HDjDV8SpyqJIrDlyMVWTYet+IfT6
s0HBSnA0c3Ny8jznU15JC6VKnVnIp7MBZumjx1A3p0pp6bYo6LEK5ZIzLej3l2Y1
ncDHO6vKcodmiN3CBGNeOqgbOtxlx1X9qzeyKy8pBvRmzcNbtvswqBuFW2gaO50b
8Z1A6K5bVYj1zO0qBPqKWpcKn3H5323FFurJXKn0lpYd/8404zL+4XZ7YuYz4UzS
/glqMYtS3VbnqFf2bh0QCuwpUnKidSLPA3/UhYCr4DzLVsg4BSbArgkrg8WI0OHC
uCZjB82PA6kgC5UqxmhGU/I8YGhxGk4zegO4zW8jjxwadONATy97fjH8ZKLw0I0y
lL4T9a03DeRVFIl+DvXfLH4qgx76BW7iXHgCWE/Y1B2Lc/lyuoProcu2hOaqaBwe
zmBjamIw7OoJ3wbbuZJtLabrzkHIiJLH3RlZaO1OLipQSTrhlrA13LMtFYIWbze1
Y/SllQK1pK1LqsKUOOn5/tF+iRoTeNQeTHyc0TzTGboS9sus9oIVqGR0xn5jy58l
FyUJ7H1ALhWta8+fu4hKCHEZZbUqS7ykSOdZygv0+Q/ZDLjiiRY2QStJWsr2vt0r
gcWOyBjLcLHlpV2c1AFxLstWC13Ptzk1/UOBNKwQTQOApIBf74jD9V7wX0suX07c
btuJOgvDJGbme9LDooXe3iquGzf/53Rhi21+j9WZjSkNJyw7IV/5StZGksQUpAP/
w2PJIG/Q39Kh17wu6Ocr3ddOd+hK7kO/sirG14pdg7VZHQ0S4LNEf456bI5Y1WMx
uTtXbcHdy/0ySHXMgsTlo6i38ReK5veGLhcFEIhLJmQY7rCIFE51q9Du+MG0LHqN
o78ilJDWYCimbjdWpUpwZYu33iI5dpA6DNqE5bhsZhj5T+CpbTRMM1qFHLwZSUW1
SEezh1omgAnY9egfgN3qaFvJj/XNAbnm0XzV269oA9O9PZ3OppL3owbHQnQc+HMp
tNiOHBtdWbcAocaByyriiplzRaABXd928/A2HLjO4tIO3Dhq2BBeF/RKSBnWybLH
FK8CMF2oqA5zvYHOaD3AUUAPeFd5sxJ7zzjxdugoHD1wrzv9DRDxJQ4Azhs/YvuB
srN+S7qhhuA6zMmFxcvAGdU4gjIE+aPBCei26G7tp7xG/kQQ6NZVXKsQ/ecFxVGJ
bmeqm5Di7EtdqpcYPzlOfFzuhNI+i4sJ+48ihJt5fSohznd+8diWDK1ZdqHbShLN
LvFRKzhdiiQpntHwHZAZbW/dqKQ8GafVggK40OELdTrG6rAMf/eDkvmsD+02RC7C
u9qoX7851+vRWH3xhMTprUO5GPrIVyiacDjEci8PeH8jveYRbmeoLhyBFj1aN2Dx
enFy1iwKkH7qk9m0003l70Hv/pXCccuGRZXziOM3h0OBdM5DSlMeVJ3/fzs7M7w7
ysX1L9Y6h4kZqOUSRh4eg35F1AGm4mj1yNR7N9y+m6gXUcHWQWdnDBOHw8cxyDrA
gMYG21+9AQQuWSdD/Hn5bfFleRZrlGFOr9b2Rl2zMZv6QNznl1OKuOWN9DsTq83G
9PVFW2tTjTgsSgCAjEU8RXZonqHTBfxwvUjOGLbbUBv8W1VDkpYbCBCtXvwxPC6R
SseSwlnzVkMN9YWD5MDEedLNtOk4nKzWfirtgFqzdcOhcivVN/amzPg1yCuAXJej
QFveAHD+BujTvSzq3/9xeyCUDyUOx2ql+MIllWIX1rWEBdMOpGwzjawQ8ek/FGdf
6mdEgZaKzs5L4438z6Feay3TjiBkyMwzWsWilhg9vnKT/1ye3eualLLLgNTHndft
SyLLJ7r0Tmci8dU6yZmVNjcAaPrtYy48+qIp4IOqxuz7P33yRs+51yKGPGjbeLyd
OQmcF1dioK1hyH1Dff4lyFdKJj5QbSTT6Fs1imgbIE0V/epo9RjxXJIZYX5rsOau
RYUiJ69fLpEPxnSGm2RQD+t8Ib1HFMimOKzePFyl4n2PgQsyVzTVcDNgdJaWNWWK
srDdsnbL+jfyaH5q3srH/rIUgLhqdZVl+GEs3rHOX2j0nGxWqTPEwBdOjHadEN+O
cPCWuGmERyLFJzV1uGPFtWA/LDLWcFkOjFYrHEat0kUjH1s6c7BS+ThLsHRH/lXk
CUU9+NhovQuX3lJetIdOg7ob5hIUBF8XfqPxdXrnQ4xvi/ATAI4uJuK6eXsiKjiL
7e+VC+p1LyjuULIIPfJbDq3XJFOTYpH/gmpUDtWIMgbutJjIQMB0miOe0vQX29lr
JHWowoMcIrkhgOl6BpSHPDswpF54HtKC8JP2oO23OXwQpQZcpvnPTHjPIfhtx/uo
ROkvyjwLNMzpeYbuBwtBVyJsAMsaxPavsHHk0w1EeZYUWRTTG2IYP/6ZBWEp753E
wO+wd5FrMvAEyIH4Gnz5X2hWEvlZkZTb2keqI4nBIbMEfD8fT4Jbmq0b5geBBiic
wbgpy+MAoa6cEgQJnEimoe1UtupjIkZakdc5DGGocztyJz35anXCpMOSBy7XZ3cS
jzq1z/ERGCsGbUIHIj4Ato+dPTGZ9xT1xyQcQffcjWp3yeC9g6fKQrF1evUOALcb
axkEmIcC6E13I6G+f7mWUDGes4x+pkd3kXVdAceQX10aV8UKrRfJ21zdZVgjxlwN
zYGHhFpo6C+VzztaujarsEeoYvy7CIek5NahXWndTS4qMRZKo2saxzYqJ3kkcFoZ
lItp3d0ayMftV0MyxN+kAtI1yN34q8Ea9JOIcKg7q17PO60rNYf5lytv+Z2j2z1T
uSU2qhHQ89U3HxPsSZp5J4pCQbXFvPwFNb60uwntpUjHN2UN4R0HwtCVRN2mboX5
6cRuoqgMKUz9tifYx91ciG8fSEUB1O1tOoOz7Ps80XyZcpF8EVd+qDHqIb8yDB/2
g35RzBv3bWMAzsvNeqIu+2jK25QAPoaJnZNOhcSmWvaoty2zE3UXA62+pdioxZW4
JsnjVPqu6oOCpWxjhTo0HgYl587Mkn2Hc0AXMUYQSXogRBc3WIURrX+bk3UqA31V
eGJLVxX9FTfXLUx2RuY7HhDXQqpB+NbGcm6erzU5H+CU0SBHL+dc5O+cafi5wfjE
HuqB7ULu06sqi3qzyNa+8iWbKJTIaAl5rKchDjGiwRks/Tx2MPOmvjCpKGy18AJm
K3VTP1ddi4ES21mqERp8S8wkCpndX6gTST9UyJ0+8nJgF2Oxl2i+4rtkbAsh0vLN
0jFWZ2oefWSqv4jTushVou98S98dMdJr7CEKHricKvKTT2HKt0nwid+zLP+i1ImK
b1GmhDBqb1htyZWCK9+kD9qypmnXHJPyGZ7iUEL9VVLN6o/I6FLAkuD7utHvM2a9
bPH1MNfRCVnitFHkxvU+Xu4j+z5+Lr3iEr3cuVAJ7rFQeqiWqFJznp5Xi9McIPzw
YlYYqOZj1S7skJ0dHooZc1a5fDj60HnaOHLd75k30mZcsRvJK63MiDwb9gMSq2IH
NP9rgJqimC2GLlB8xAX+v+8Jty3VDkfx94xj7kx4iqSsIUEVvf4BvUsEQkaM4bMy
txfME8rnPKSADiWq55QCUvThRf8S//Lfkpw9a5tqbBoNYLZI+xEIqOLAp9faodcC
GtL2oCmQp7R1MeopSbWqd6KnOh6jLmLXAXUv7e9dwRJuG1THuUcIS4qGXWc/h7pv
gbVENdZm4H47xAG6kFKH2v7k96CwzZiOlxLvGipgntoim+vQN+BNvIAg2kJ0O9ug
Z8zWqYNCK3gfZdON6hQnYcPsZRK1l8HDF/NqdTjYWLYHAsLBtT/+Jk4I5UeDWLc4
yBsKqPDDYHYpIipWw3oayO+Ju+yS2lcWX0IOkLV+wFxfYcjPtW6GPq5/dDMLX8rR
5iO5h80bp5x/xveSNIrHafUlYhfclXcyqU6GE6Mx160LXHAgBNMrDxnBu9vzS5yh
3BagxvlTOhjgqRbJCDzd8auqFCD8ZvpzUVmxVXPsd/FqzxHj8HaXR0OR33GTGH0y
ycapUj8wVTPR/stypzT7dTAEiusdANwDmlI5Q/3BGXRNFfzEzk0X7RFF+yoGFcsM
MO/mY/25rDuJJnfW6d0tRIPkmjAEoa8CNhequA+ZAD5ivaQECZTREwXlH8lV/icu
U7kMaJO9wamdh+86BvdhjZ5PDO5owR0ji4VKVR6N9DQxoDiWP5i+bcbTQvjmdF/K
mZtIcjai26owVMdWfS3bebnnGi5iXcA48/hJZNk+QRaZXjVj6+dAc1aTO0MIXWZZ
oyKhRxFmO1qOf/kslp9VEi+nxofpbzXHyMq912zWqwhTA9wpNbZXZIvNfwxAss4q
2TyLVzE4LX1qTi80y/HgaXYGZHaW2zrR4DpcZgb39vGb3W/G3SvQgfupJEr6SBwa
7uwdxbECStb+jDjBbEnUtBCLZ7uy4BIVbIUuFhJRmuNeDd7OI+mfKoC11nZOrQzG
GJ0wRnc+vWM3lhGn3ctwT1JxtmgPnvGihWwlwa7FHJRY6hdGqPKLfA+kAQgvx9jV
6nqCn7Gn/2koOGaUfjeuBlrGUXo8fOwL+YJULYHh+TlO3a8F3yslUNZun/7Y+bS2
arRwKG/vfTtF19Nvr4XGAPGZkChbBLwOB7UtocxPtnsL9WMPKiw1uEW0LF59z52F
kD2V9mhLY4mHJGugSSG3S7tIKwNFjazHEw4z3AZgPoxR6dhc1tfheK9n4MHBf3k8
JbXEaQeUbaxMED42/oBq7ZNpUZbtnYXa99s1kBC7NIyv6q+WWGIM70GYDnS6gC2k
p6VtJBoq2pC1xoJExXnkvd9hVC0pGQLOwSMxyMayHemcx88Hw5ahh2CxYhsTmcqB
ggVs9UttH0P6vJH+hFXl8rq8h/0DfRTFPm2E3kmzx3/EmY74Yu2JyynpGRKKQQth
mmdLzmDd+ucVUORjzYTZVo1A2ekZyoFuPjORrAk0aY5Ub/yvmNQ2BPzbOi+Fjf6p
SQXqSTX4QyMYqsqoNO1hNz6RpACB6r+C2EZ1X8y421G01uo53KsRiaJdCWwKW6Ka
YqQ4mj65zlZgpOq6/Fu02y8PNyxwDqBnlKooLXjtJ70YRm/cqF+drJzvoDT1Vnek
3fCEWnax/HBj4CrQKKvwM8hIv37P1K3b0EIMSiD9dJdyDcM+J6G5UBG3Auw09Axi
ShQZBbCqptDyLgWKXk+UVIZLa/ZwmS8GmtI7PThSODirHGPxYCamE0jZe+pMCfD4
3jana/FiCo8qs0aq/QuyWmDi6ljO4UGTZ13DvwH9SbzHlKjjFe2Rxi7AWFhjYlKh
4APVuDeDny++e+SnhY1y2oGIi+EfHWFpc/+ltQmT/W1aVWy0Y63lc/k+btqzdeCF
osjtd62wmOmHqGZfbALlvJYcBP29GxCGV+kUPGANTO2crPtJ2ztyLGA6bg9xSfQQ
Cw1nlpWrQQ40HhRzLxD7Is/PDwoUe+uPa+EY9B8wU8tqEvdu10mCGWTM4g8G0N3Q
3c+sRdjvaX+ICgVGUv3FlPrr28xmamh6OcVz3F4iQhUv+4SAtFP3PM5axSLMIQc/
7OhTYHarHnO/4ubi2rq80jpITBKe6qCTMfLBV8UL23Zw0p6qbgd9n+aT8JM2STuh
d9SY2hS3p8SGgArzbEpJgG751Sk8ZRW9wfgTh13zAWtqv5hle6r4rYicItQ5WLJj
LPFmaUnAPcmVh1HTRgv+oVQXjGxX/e1cL4cqEZMHcr6GJJCrXXIkkU3VvdirtyZS
gnVktEJ12xE5H4v4W3wXsBRTkXcno97K9AbppgVppxyzMY27SOEMIdbbGSue39pM
y7aX49/v30LLqzurdwp3cvKWHZvLENQH7QIKFutuTsbGlIgUGn5m/+GVtpxElsCz
k7eC7T1YhjRLgFUDKinAP18aYAb/QbU/VULauSENZymBmtuhAZhPKcn8zOwme/J0
yK8AeO5zIlyzDRVDryl+BPMUfa7wo6OvDCQDN2dSdfHonSaaE80B5O4VSulmS1eZ
mUmuAzKgvG2+Dh2Lhh4GBXiQzaDS4lACBuswerFLr+g0IkiM/xSHw0GYQw7NyyaL
UJu8Jaql+s/vXU5HkB4+maGQVRIiYo0As33F6nZ4Ees0zEyvc3Es3XSvV3prIpcn
wHpzGQ1jvsTw6Nk5W0wmAvUY2sTMpuCwoJTMwCaR73HCF8ZlAsFUnoEFOjpL87vC
mPAdC9ssCgtr0M3nQKIsPj/PegFrb8z+bXO5bPZotgsz1htKXQQw65RmKqEZj+Jw
BuI94fYh1W3nBxRd9z5r6QuBWMH7vsIGOxsa47J51igcOtsckbyaB03f1BrcFo3I
iaV5IQkYFY+g1DWBP48rg9P2peMPKATXVDxWDPRomjhftJL7FaqYiZl5vU3aUQuD
MRSmEYynJoCwH6f6yPErTT5+s+FJpl97aUN65elfL/Gr0dvwSc2Rmz/Vjemv+dCJ
01aX8ztiIt/JIGAGRH2ydqXhF5AJDqcosuN+KDCe/xW7prjsmi48vCwwKN5/lDIL
DTFKZllFGQwPFpLCx+TfP+GMzO249YQEalYxL7tl/3QEvF6WrxO9CunmnShvlREC
rKFWhlc/0tkCPw8DLyBYkPEGz66C/eUb6/XSoNfypaUHbpoy6zE4ieMvCVeB39j1
ET/UinBt31+E8WIutfqDpFrvD75fKK4TxgzjCJEG8HOE8kw62rnzrnH6DsN6gbv9
Wbb4rqb20aa2BSf++puoU/NLQgr5x7DGAL+Tpo7MK7WFc8DTSIG6ABlo76ZFetwa
RrfXGT67jtfXb55CM/yXNk6IjmL+ClIbZRwiAKEq7Mu/XjBcXah/BSMFI/rBJLmz
qhfo4V0aoPjGToQs43u4DhXUeAgi55X8XB85Q1VIlFMc8wES7teKk84QXtAE8AMK
/erAhaWYputbVG3ylgeaeyMy2gbRaVepohzeht+WT/MDXuwrwXfrXK9GTNH/JRXF
UYFuNYAMF3p90dfZOxSX8jQc2PxCrK956cGnxuJKZdDaYtUpr2yJMz36b5YYy9p8
k/PS1r1Zjqe4QWj9T3J4OSsI80JIuMZ5lfQb11jHROVd8sWEpeVxDrUeuEKAX9lX
XojSXEj1WBKSD05VgSeseqSj8LIBRcr0Ga85KEPX54IdJ2weI9X++Rmt+k1sxw94
4I7EsU9NXraDAA5K/7jPsYY2xg9TnpTJS/d2pOzzqkPvK4cCsYEGGS+RG93AJoNK
Ri6sgbQ/pPTE7ehB5o8EdhxB1Esc7gv+0qrm/OELjf0WVRS7SvmVNsheD2OxnJnT
QxzZ+tQ9W3HZ4qxhvA3dM4sPUkJbd+mxkHwINheTKefIu/lMWf+9An79VhVUtGe2
5F8EwKi1j+WL6iG+cETiNcdXxK5Ppxd0Iw9ronS4gtiXC28uNzT5WHXr4DH89xcu
bjb79BKVOk6NRrYQQSLO9pbaiKQXCXZzApVyUCzX4aXviDX/8eJcKHadcS4bMKzE
tJXNxlRnS3IrHZPsJDsUqXbrCqXV0vIbm5RmtjBaxPLa5h41930wmT2WzYEGMu8a
yfGviBsdcOhAjKY2j2ytg24l+U76ArQI7BNS/vT0XQx2bwAvMB9nmvOtgSTx1Uaa
5vxVrjiUDMLP8ROxNqPxGR7c9qZ3AZGsocVtabkhfCjHmXOdHQM6RlOP4W7FLDie
Qeka3sVN0p0oWpaBqA4yoTp/r8peBvajK5IPK5gImLdCsBMSCHt4w3Dt3hYH+B0N
5Z80891AO7IAWG7YVGHcOyJa8fIRQl5ftKF6agrqGLKboQS93GuGqet57pZRlIIr
iznSOtFwKsv+w4ugwKEM/kzyPy4yAtpxCs65xAhxKee4xmaZL+xcxK6VYA0vQGR1
6Xn8YNqSLHNmlGUTy9CXd/nTgNqv5BVl3dZMmsXwE2vwdkXNqAaZI2iDHya65Nh6
FdUbWKk8pRT6XPs+7JfQ0krXn7AHd2FtvMt3sjixDgRLttT0OdN1EKEKGrF0/UVG
xhMh+/QS8YjVwx48WPIxO8dnH0q0BhZm7newpKofCVMfmy+aUSFLorJ+c4mFbGsv
9COqKmJjsPckOj6+6OaGMOgsWV6qrPyBFP7BbofsluvRJ2BfWabfthpA1PzJsVWn
mhEtO5NMKUrQnsLFNY6Phyb0WQ0TRnkVwc4WY+gpAAdzFVFX6LEuJXYGovyLxaZv
HTMwGBPVEcDxMc9x6OVjalIlkdrI6weGHPr0FKtrk2t7wvnrjHpISttQFjTjmbC8
0V1pUz8WDaKN36sdKqKeqFeHoDqkU6mK3WxItam98ejo488OUQ0+8skWHfnunMXE
8IH+jDWIOsVITcwmkYAqMmszVTWDbXLn7x4FycIXZnTNjzWVWLmoY5GPn0zJ6nnq
379kvjqRjA6rmNKPN1kRiWzDheR3w9QvoyMbvKN4wKuYrpW6hTbC8YHzI4ZRRu0b
zlvSPs6KzXlfdwVoSX2CDxVZ9pJa5c5MMHtNSCcUANK+BeZ/Zzmutfnlw6jMQENt
8JSzxvHJzs1qMSxpTVRcDReMN4q4POy2VP73eXvVeq//PXfCSM6PXRI/lK+E8dZ4
bS5NDGr3ev5qlsk5jbktzmISHptBxZCL7WDFB7Ks/frpI6OE/V5k+z9JZSJtAT96
qoqzrFd57M3R3hlE6lKcys1i3Fme0COhtTKgbM7hdY+kbjGaVcsMn+whXx/+GkhW
ZgMYLR7FVxkj/9N1x4F4rmZwRGAinYSU9pCL+dJgoIMhIdUeNvgqz5CtZnIWMGDd
fUodv7aDy+6X/fyx7hTgQhEfZYVQU7SIwdLCIcaHB89o8cAqhfKWq//zAiScvpTl
jP7zP/dFzqqCMWD3dlF7PsSAILEZNGCWvryNqhagf5t7r/3NrmiBJ2QRkzct4/CK
c790G0J5McBb3Vpx2mCzevYnYjlmytx2ToIiGIyI92D9DcQ8DHAShNGRptvSoa3r
lANKGl5V4wXIGHok2o1WZHtXuGPs4TtZriERg95Kk2YcCVB5pwFodDkgKuUDedJX
m+F9ZZcQ0xALiL1kZhF0R656AOeYqy9o0gIMVvyTv1BWwg6OCbG7h2oW/cjP35Mp
dSVPKHU8K3sGh5NUBth/NQEdks4VqcdPtgVrLPJ0NkMhTH7hEU0I9WbUSoKMI4kf
nqbfTd9JO3SGmn1LKuFZnkKuJtbLHOc5pu0hDTQftk8iaTgrBv0t1O3StUTwDe6m
1KCj527ktjlkJ/DVwttdIzCtdkL4WF+dD2JxhVCEVEynXbCsOG7RWgcApyykGtSW
8RB6+pzO08KY954LLBZ5q6m3BY/Wmn538+etXeck11sFeia/l7S5RaPRw1dWnibF
JNmfb4QGrV4q6O6lcZckHS8IO7iW6SeFYHJdep1YFhH+LzftXEiNTv3mi8cO5YSn
X4T0957TRzapZJ70ZQJ/B2yPAg9oCetyIAkAcO22CQKiiy/n8+DH9tWUSiW8bCYT
HPvU5GN53He+N5hps/90bWyyeVdxOa2hSMGRsypt0OmJRdMbrn1aTzONe9LwIaP7
HPiBki1BlB6VJHo0X7MSS3WgJBesq2f8aFUqMiWYCP9j6CLZLtJx/RGzC82B3b+M
mdFWzV2b2x0699EVYfbSESZDZgKCxITpxIZLH/22leqgnIAUIto1CD3FiPjjK/eR
fHs7KIW7HqutL25yd2cBX2P1tzmUM9pHo06kE8tJrHhSLhbmnzrJt0OXX3D2VQ1Q
mvsakGWc3UjwVteEU0vYDRzihVeLDvuLrd4zkMGE9UA+S4uuyai3OM1RDBDA6syD
EnK2ceg9arvGUiBSwXZvwB5/rPEK5zdml3kAMbSa7Q9TX5F8+GYOY+VcRXKtjqDQ
o3MUpWSNPI2gXFHZ6EV5zUu9nUuDAbfTPn8vC7PirrBUDRFjqKizPNHpIarEBYGR
TNEAeyaOqQEbn8J7CA5PwtSaK42pf5z5n0W4EibWGO4+YBD9i7kjJr2NVs79C31g
X205w7anJ8Nt3wMGr+2UrbzO2VAzPnlgbgvYwaTdWrPfw3n9uLAvBQHMQA49KSDn
2fboSrwS168/r8f94ZCAarA5MmhWVTmio33rsNKPYHzCOaYkBwu5gHkBknbAURsO
jTKMI6mpPu6Ngj9R5EMV8cQ0rGLDSShDUWiiaLmU+0mlOsv3LcCcppm9222YLNYC
8CAQ7QMsuv7/ts93qYhtuTZHXstpxaT0Z9RFjZo5jK0FYms8Erbn3XhUxJ9WqEOq
aQpxA4m88cf6T7JAbAK5oyg61vLrxdiOH1L0rszsl3vReS6qHNhQc6/k1MKKZxBM
cGHvrohIeTYoEXcoyhgyJTSwTofT5m/TFP33A0q7bvkMREOcDVYfXufprz8zbvbj
ETj0e1OUu4JVRE5/Ex/efamvalqRNqRHUU3+9HWcE2ynHRpiij7QX03MLQK2Vh2z
egpWtgwSzajWCazWXC9rMiFpxQOxWA3qAZEq1ZO2b0qBf8YrLZnnrIlo3wQAhjB7
QXy9OcPEAiK1+ycmFYqxbvgaWNyH4b6FSPMRnjGPu9GRc8clqZKoU2haJrSgy4jW
MvquUSMCGxrM5OXE5aH4jU9/1lpHCHCMLp9QmKSosdT4Aq4aVOLcZu2DrSmkhEw0
aW96x8I2+xlkcNwZ9Djy+/RHMJleG/TcO7X1jS2ysbzm2GkmGa3aDOBbonoRP5Ff
D5/psJRU5IqTWgsrVcVvBnJSNyuReexIMXL7ReJkGE7IMe+FTGNGdlvxvPuAaxue
m5WxhvMovkxKMccDiaC71eUx93FY8wXrlBjc+dx9CehCIUS9eYBCnyXeNjaq52y9
y+eNqDMyqvFgzJctXNPdDY4DvSeQ/aHgLhCiaAuUMx63DmBakaiv/xAmitSWq/jR
gIlOrB33V7z1Y4UNFxA9lRRg0pJIo5p3kBagW7bPyfza/KeO9EcYqPXMZkKRaUp4
FzBlL3DESiEfHw4d6m+FXE2k4QLhSS6NNajB5J/ppkFroKJR9hkGtvjSZdvSgSPx
2NhGjOglm8GIKtEHpmnbewSdDGvMyYLQLbWjNg74oxGtbp61gomhMlrXGeNDslf5
RKnCrTve1iLoR7yl5xErmvMt0rIewJn26mtrt3FaljIGOhyB+T5apptinPTrP23O
1C84YFRTpxCG9ZmhDgGTPmCfyQBHfgHCsAyK6nt1p98jxVKajRp1O3xHHUFjnLAn
40LEdzfXMaFY8/tyoegp0B/zWbK2EBzbcEhFcqQt8upXRlhiGBLun4CFGgHG9Ukl
6yGeD/cOrXLjwPURlflzHfW9IrHYqrGYlOcaWXBWsHbdE6WZGdYelZE7XN8igLzD
AHRHTp40VfD7Dx3aAheQ/49E0ediHpdYwPYX2UsKNOPE52xkpk76dl0r9QzQ6Z1Z
HecJ49yGPU+/YsGGaz3M4PKMLwTv5+h7CiuDE+ITmsw923yyNgW5NHU+XhRAvND6
5371Q+Czxm0qG/IuG3gPYl4ngmy5C0Nuyjmf1PR583R13DYax3dHEbffFmZeGjpX
H4u2694oQSrjQIvqDlP8kKIdcgoio9YnCzpFGGD/qak3DB0ERQ97VRyhAciO3d6P
ufYtgJfumabSEKVK/IqLDrp1hOdfqjeBQzt0QS9cHqCmaxwJOUIlhenvJ1+K14YS
yDIkmKEU8S+U/tlrN8gFP/PMBsx9EhxFRYNFf+HOAs4oBY+dtd3esBncE7Pl6zkv
5PqRXSz97sr/BbMj9exypMCBJjVyNhhNSvQS/CxCHIg0SIc9piOE+vYx8k0sq5QJ
DG2ddyq5pVoKDUESZv57XjuSPWJfl/2084Ed/Ol1LQmnyuw2wTLL5yhC0ceRPkP0
P4HzhHFjwxixrt7Yj3kSdMPhhuAkIH0KXCoCMiTU8XInox4xq7DC/aCGeeXKL8JT
4sbyQSepzF/sflIxiSZJIMfz69k98rd7iOe/V0sYVIeJb7J9L+onZwI6WSe8d7XL
uXdQkpuxhJzasFRVG3yyPtAbS0jlkpSm0cpTOv6NIQnM70dNvkGhgL7lhY6n9V5v
P0CJJL1Qu5mW6Mq0pLMU2yEoxto+AQZUFox/BZPrRTDTXGLChjIvYWe92raz9noa
dDHMGwuybiS5zwjfU1Ki0Mb39AMnf1/RXd1L4E/+WQgAczE0XJBfOegN6wXxL9ZW
a41nHeIOcqAiwypQvweYpBeX/3l6XnsTe8jel9PqmVUXTQ+4BZr5Xyj/aptq1gpz
O0laZ1afh4fiMv/cG3B8vAfhQy1XJAw882u1P6idqjReppNossqgKD64lXxo9H1G
rwNt8u3692EHMV/sUu6KJbNm2/Db8iQTlqZi01A+HTDXINHde0UBJ5fnRYyMqGqd
zOoRs8dak9Mpp7bU5IuqaMJ5Hio/CVbL5imIMzew8j874D+U/oO1bdUlWHa+E6/z
A2o/H5Uw80f14rn8o8qa4yOrS4jKMKdR8QySNsTFJU1t1ZDn9zDhIUQanf4ub4tJ
VOdkpEb8n6VfjeDHLTA+X7tUyXOirH4WyfBjpzx5jbgAtsaj9FZZ+4ZfGUcR6psc
8CESGLW9H+prRpLL0QdsKMEANPIDj7IcGiuYkJlkRH3J9QKVj9G+uC3B239ft1BY
zoxubQom9SD27V2OmwiIBrX9iGRN41UiI0gc6DBAvkJxqQ4tG7w629PQruyo9o0M
TCe+3lrgp22g44N/+EQZl3srj3o8mpXDJX7bpn/6ab7P1+ZiR/xjOYOiMXnwLd98
iOr1MI6UWEL7/p11S4zMQjyKO4bftxpDWF22ZbeG+qPJjlG8TaCjvCtvEs7+au6b
8G3cT6L6kxZuLEIqUP5azQmK//NNsSvlZlWXa9+OtQtr0T9XlWR9KLCxfDbV39M/
4Xy2k6jlIx/fxNJUycLvS+k8IUJzkZEADckiylaR0iPYFP4aZ8Qo8HV4gcaWM7dB
FY8egQUn0AVfQycYaBeh/8evBb4uhi1t2lQIMD2ZfE6AQXUV6yboFFZUFrbBYkum
QVuTXX4V3bxO/28PI5k2squvuUaKUiLMmNORc1GSwONZRSaZAaZl83SKMguj/kwc
lm56hfnvwr4U/jsSqWhA6qy3KUf+oPOLeHeZNMHl1okk4JIQEBz/3gZdZWnN/SEB
3zHpsdv4Ac9+rC2uVAyS21EUkDxexIks7+jdu6nb3CaGuf80L75HSXooOZjiZobx
nIt2EPEOsXAjcoLZKyFkAnbvtOdr8gUwKQkBJrEr50+jZ7py2ovIYbAIUD7dDnL8
jab1a/mz62xBMWjElYlHxNjk8jNW4qtgcbGk6SpqLv04r2av8eh7rAuDE8bDsa+p
GeOpWTvl21Zof9hWgID5XTMtQmmRbq8Tvpz1I8ZRM0vD62CS5Ax3LMBeqHLiDGIp
rxaQ44Ex3upXz+iFQmfaWvjjrXmdyf6NsVZMpLEW5yYiegRHA/wmut5yAHuY86Kn
B+nSlXJOxb02Tvb6qLlO+WYYENxEjShVx8+28NTCVuXH2iaedAOuuJ5GR0p47gkd
bfR0EObT++tF+WX1I861slFqUb17+gq7paz8B1so7W2qZMrlxmN7qY4FJ/cpXvIV
n4fi0R/yBBuOe//IG9RIFCtirq2zLdL5Zga1jw4AKPE8SKMp5ysg098qHpxEYSi0
bGNQ9DX2llOgvu0sv4WEnQtDe2KhPrcESUa/Nb40Woumpv07IO/G5bc5FEr9D3Nf
KZ48ao9Gz2qP8/s+TD3/6aE4vKf4hPUu8zg8RQUrQU5QQYXSBdBO1MiD6GEdJeWu
CJW1X8YVE43B0qjjsmA7ajLYTKoFwlnbeGo9eMLQ+i4TSIaRLyCivjRq3kQ+S0Qa
f0Ul8eDF6W0eUr1kdaL0ZS/abOosMSiTWFTDahz5atoQeGOFL0pxgvd7Dv4NgScs
aZCQmPKECS91HJ4HIcAw0iAc2fFlH7rRP6lTbmeayKfDwmm0MAmj1PsLPs++YK3h
hFf/p0MNYJwGM1KSjmLkroi/tgOk+ye8kGSGiXUeVQOc4wD4aANmregGUd0heExm
d6AM3n17268x/og1U3xDQ/7tfcJYSOMh85e4AzUeJw6gUtu5Ik1ocp15UG8zaIgz
I4Tkt+ZcbnYvtv1m7POp+50sA0e6cbFVwocSbPMV2qHqDkI4dT48bTSBX6WY+HRY
g3fHdQfwvf/s7J1HSKhAD3MKKho7CVWQ4sFgHVeLKW1/z4c0TZSy07Wl22TrwnwC
dPU5NogujjEyJ3WJUXe5+G/uw87CBlTub3tyaA+epidaZ2WQDlD8nU1zQHvmAhoF
zW6tdQdLeN0LG0P/G8878Iav9X0WoDUAa50EcOLDE1VYukR1C3OXOuFQBKKC424A
qGo5w2VNkI/ZLzh3x9+o72o3hOOXFjNeiU31kXxwqqHI1n6n2sQgK/YvUFQWJO4G
NhP6/7KzruzJMnAXnz5jITO45gs2PeWCRpRPAhbvhm0fobh1vagcQM07zy/lK8Ak
1JJlTarQ/RYBXi7+hINRp0GUqRz2NJ/x4AP0asXJznUqGfOP6tsA/R8xX1ce60HD
rpJwcI1oJhqt5tElyDKNNOQ42jv3YBFo1rma0e/XrTk11jDWRjYIKWhURUGmWWvc
PhHQ0RhU+agZZ3pGOHRUS+Z8L4mvEe6yMiwXRdMrv2IOvNNcelarininRO+5C260
IjUg84Xl5jEL1Ax57tmBT8QJR6esdXZBXtNikSTyE8naQFcwDo4uPxM0H01369pM
+WGdKGE3JFyzOQMaMAZaNjxkNbBYbByMdSZiIZcGU5e7GwYx7vNvbkh/zzqHU4LD
NpImD3HQI0chvK4W6Y02JC6dDYUFFDNTxpagB7on0agEJnNDU6PVfWlUjujMQWhL
AtSQF0objTTa4Y6dpcBOFbxiQYlnJoFhFKQIyE0Q9A/QLhvWkNJiDW9FD61whLI1
weawbSiJzvR6C2pbi6jIHrNfpB/LJQZIOi/FWZ7DaqX9v2J+gdbvyfXavi5eDmzU
15m0pFkT/3RrpyV+qOYg3ziRXuBl6bdVFHB2V4B4RaM4rfdx/NJl8BHRlGKNIXZy
daU1Aj5lr1bperZwYz7K1adGnH/ekBka17KK4ZefZGASPYtriWBTAV0eBVCbVjBi
FBt1AIo/2+sxY2UFK1Ix2DoZ1Qv1Q+LNTjF2OUc8WwQeHEmor86Wg0q4ExdyJVN7
iRjD+4+jVthGcNTyx23hH0mcCLUlMsf4B0U3F4uw/m3jDUv3bydjvnoxRNhlyL5+
Kr09oD0dc9tfczv0ZuMx/jfpPmPEKbq07dnMAG7fcOj6fO8IT5IFyBb6+IyD3hUw
2OQWTMHfcj+QSq6ZP1YLzQIAE6yOpqPYL5u3NSAwGNGcOAL1FyeNqD7o8vhkrsRn
pJtuNGvfRw9pBtCugU9PA0Au8b1A4wSpk5tXG59i3zVUxXzeXWXW7BJ3sw7MSeIE
NubporkFiJemCQ44ZL9yLvlUdhWPeUgg9V+EQO/dJRtLxN1kg8tCzEzaPpVsLqdH
qlzDWBArY7nzSrRkuKmApUsmEN2FWxNF+lt8maxAlZV85EKCWhWEiNtlHxFZ+io8
1FBHtrzDQEy3x/vBFQ1HE48sDAGTwIh6/2sVhNxUrlnvR9Pdw3moEyG9V7sf82Pg
ILl/g22Q6Jfw0TStkyZXOQvhWRQR/Ni9tot91op8lUmb/jx490nSEApByn53p62y
kVQ8kjTFl2m7iD2GcLdO3f4T7GC/1sSw0nRUUk9k9YHXffpYgjcoPXek62v513yN
dg2NhKLQyAKo1nMXFzPa3RG4pgQLk0KEN/zADTIofseFEHEXp5fO8E610vnW2Own
Nz+4rvtzndQXSq33+9BCAb45Zt7OCVvlvSxE3a1Iwh17aO0jFmJI+nRlSKwMXvBH
ot6azUBQtqGUJBxFD2pz5kx+X0quIxf7rV4r8vmwd9cZLLs4xmRkkjZ2JL+RfEcy
UcQJnblmE/a/uKozGA93vW43Y76tMf+NVuV+qBq2YsVBMj4p9DuQUMTGTRHLk4co
M/N9kK4VmArcVoReWnwOv6WUk01FSOPtSMbXaD3AN9kXOSTSNRgyIWGPO9H5EAxW
DJFeQpfS9xKOnLAV8xthyxOqeHndZwlwfjssN33xCrGO8TriZS6Uq1uwN6yIjOSq
oHdNCrKOlEXg4kbH9HqzGc/de8xAYn0zpYWuSkbZG5+j9kPogJNZSyQubp9UjdRd
XF3aXk7HAO5oMF1U+L2xE2Gj2m/TKTy+SB9h7lBP6Ko88e+7Y+XJGSnIXJYaBj4i
XNwU5YiCifbtEjWPXubCxBlfNJb0TjNPzeUXXwFnSxFOFDPNUvue6s2apYPlnsAV
8nI+33oKdJxFMy8sUtprNP2mD5S+BtwZ1osUDV198U1a9q3Lvvu5KOREPIEXiQt5
XTGtnhvu4jB1g17l8DR+tgIcmzi0r0OKtsvmyf2dZR3BlgvYSIJDmBihzFhj2VM3
n6I2cVlnexaxCzYZT1EINtqrsSel4qb57GiQOSR+xXlM61vcHTLmvF29twNh79n0
0WS3NsXgAnImB/IhAEhDfQfc1+GFHwPg6RxlqMNumaBqEGg6EKpEEvMHKgwoB89A
qY71N16tuYtjeLLk1unxyU3OHeai/6mysa+hpHT53ttOhMBy7tieLeoAdor3NLLy
7rZnfDRQ5cLaoA/8vd2+EOIhvrii96i3F0rdTPThoH3eZsDIM0qORAxAqdV3Vcle
oOhODCOEI+Z67nZly47/DzrwhN9LwisVvpJ777ze1gD6UwzuL6fMXBs1Oq99hna6
jiS7Ods4RMEJmu0Roy8nloBkkv1wPEOa1/bPJP1BEqWPakNoMQsXzHLME6F5fkdI
+hWfsRVxHm2ooPNsEQb4Df4pim08ufHmeBUezb+b06PaaQIDrPUwmMMGwL1EIf/W
/Ucd2jjyo1MYGruEHLv7DhrxKVO+If3GqQINBQT/391Z8csHJdSo3uXBSmeZ5Z8y
PIHXbebwkW60j/j2SKXvaxk59xcNE3V3jdlcpMgC6WoNkct1LnG+vCGllS+zA5P/
GPg6AR2V0hHPWlVR5Gwrdzp5yNZzRGXwfvIrMDlynh6a+Qt7b0BiG2ThBnytE0FH
Da4a0xfPbI4Uo9hEvliMmQ5DsWiKD9ec6jCpcpwQSsDDaR/qAAd+nt9rkHC3gohK
F521TSsUqe9VmKUmasnMjdu7wBOS3fppsdDboPpg6ZVeRQWkReGZ5WUMF181ohCj
Ae4dISLag0IK0JlmmZ7JULSCioZwUAcbnxwTu+K50Kr7lACCuSrpn2MmS5jSOH/F
OuNcSxe+H9jyPhF0LIeUEMDQLOnYoTrrKwJVzfni+e2O/COFDrcBCDfTzkQDx9Kt
V89HrferOo70avWmkc+M/U/M4+ENp0/EjBn9PXym0t+iNwn8Mkv5LV1Txqtz2NH7
6/DLoWtBFB0Q7JIDknmG0iY6nYtmQwSVCSeaZq5/n8JyJajX1E9qb0HHEufGW9z5
g1H1FHORahIrFYoyvGOxJCQVm5pwJFlLoBdDMNGH8Kd+sQJkSpdJ4DJXW+T1GqZd
kiFxZc/coknz5sKvbieLo0VIwTnUAyKYR1FKDWE1Io1ztAzw3dxYQ79rS2b3Juy1
z+FA0996p6L0E8266b6SsIDpSmZgYsPTlPjE6Q8HnTsttihfgFqkCJhcvOpjPsUF
2WoJYsHoz/Fh6yNqOiUbx4iRGGgvNv08B0c7T+ktRVoKsDNp1KMKuj2qplFPllbs
WHZz9Qiy24/w9JDQBBPwwOfO9jl5pVy9v0yu1guFrJ6zkQA8uDyjrbrdhGcOpl2n
SORWHxk+MHbTPi3/DNZglGkZnLz7se1invei1XQ+Y5iOLpCn4Yy0m1ntyLvJX9DF
/vS1Tn7EQpokAY62AJIaQy6VbuG9AyU5IGw/3eBylduRcanegAQGTXNV/g+7Saaf
RykuKt4ub1FOlFphdowTJJDwdOy8SVWhC728OkzhKg6yFsGSskhYt0Qn/NPDvF3x
n8iW/wQgBAlUBFk8OekZVgibPK0iAdZTvLzZQGIgL7L0mSEGT9ElGSP7mlhCq0EP
hqo6FRML0UZf9tpZAHcdK/iuMgEOI3TOTCnjN/w60yWHNwc0gaCk5mrWx2V787qS
yJoiirWutblk3Wg9VGukPB/odk8bu9Mk6q9abndLhSOOr7QsF4wwB4c5m+6/9Xma
28/XCKbm6y4SzBxe43ag+TS2cRgOcUC0cOQ4TEvt+vmgydaKwv8w7OJpUtl/RF9U
t6KKPVxVEVkFEoUX9cJRoA/qug6BsEXUGyu9oCmiCUg9EWuT09N163KC/fvkTGfB
CnvUqXS/cxxvnJ0I3EFygYMJBogUS2XD3tyRVAYSAr9O/V0EVv5ICMGiGedGApXg
c9Vmgg4SqbwX7wQgynYXEcbHhG3e+QYyNDt2xLopjYEfOEJTYX6EuvO4DrLYQ0cH
cD5hfj3HVWxnNR5vdJhTx2nw+06BQ+Gv12hloLuYBVA/J6l9GNcxIt+1YkwuizRT
sASZVx6CZ7e3BHcO6b5ffxFGJbzWryls3O21Gls303BURI/ELSVdrxw1Cw0aIGch
SnQSpatWewdRvRPiTeQFGY+F72OdK2gHlgYL6SpJcz0hpVgFtpH0Mrixi95t04Nw
mzNU1m6JJ/nNHOaJs0CV4BQKIEkS6FuIHs5BRQ7P/fWvWG650EjqkJauLG6LTIDB
KPYSlOdeZTDHxhQvAFLP6toGfdirv3EdHymZgwIBpeN86APo2r8GsQ9b0XvlNlXy
Z2XSckekT6C6SKQk+tQ9DSZjwOdVpxYJbcBoEn6qoczIWVc1aBTsyW9fR2pmw1Dn
2opJlPP30Lm+0h7RYbDYHFO0BkTd3QoMYZpZ1n/kyVPPQE522VxWK4SlsBd0sbeO
8GsDP7hWJ86FQYEK2myIVpxuQrSPrUW9q1cVxAbrBgchHqZ7Df7NAXPQHWLPULdI
+pTs4OEfgrBH8Wjv7LhGbqLPFdKnl7qxzYzSBYFjhFg7dw+f7Fd+dNot7a6p0M73
ogSETTXdmDt8jn88AjVgOvSsZp47yZZX4YKsL1pQqWmVTraABAKQ72JYi97IQ8wF
gmjSueKrBPjYUm+tZb61bKnigZTn867+iPLdrNQNh04c8njVQcN26gF+CUEuUAz0
SSfHgCgMi4RBahp9AnTn53GvVsFnA3d6/DCW+h/Jrfol21/MWKt3QVfwQJZj1ZZ0
OCZhk+8naCKnRdZiwwc42ExQoI/v0ggNM1sher7LsIOzLWczDoJVUFiQvQSp8mTk
tkak9C31cux9ypfXlG0JQdQx4rQi8pM/JAWrqUMfL4Y4EIPNzsxf0Y0BwCz5/ds/
0QYfU3SWetoPaisrEDF4+m8yF2KdxU2DPGfUgcYC5IhtZhWxl44vn+j3ZMkLXSOV
GBO8knNeaaLQfrMHNLYI18cO5HyZdoQeaJ5gr2b/hHjmEAiOVfOcHLU8zgcS49F9
iL0ji82laFcLnjTSUDaJ1ZMX/CSgIEbggC7iq+wP/IN6FLh6p9kkQPkpnNcHpGCz
L2qTOydcGs2RR5SLgxOP810JE69xdbmHqFiZyADqYKR9Tog1co7fXvwvoKrQgLpG
W4rlXUBecSgXVopgNXhM+2npc5busUH1z51lk6D3+yk5+uxlB8NDCTM/BYXgDuN5
0klmPGUEiTHkWd/IW/B53YlQwBKC2bO+B2AiJLcfCrKQ7Atap6t63TvHIHps7b3D
myqFVy+5S6RKVffyeuVnXXpnP3dE2cHH6RVxfB8p15Yd6GPhVcQSMD8dyAvdWx6t
2/D46tqJqyX1PjZ49nr0QFU0aV9hfOHfHzydJ+ORO41Ee61UdFIhzs1Pi4WztZSU
u42LnjBtCZHWyWjeCtChj0aAR8FsjxnctPExiAE0VijuSBeDuL75v5GuX+MlWyAe
HitZ9iArIWNuvg5RTJ22VMXx6QkuTvJc60mvoMCDja2mL25FxqGhAwhZtnhHkuex
pL9vMdciQ81Fnui6iBgEkBqRs1h87crq1oORHfGknsndGTR7Go6zMLmhl48+Ywj1
ExGvX6jEng2+0cyBnXdxKl/VaFiYbW+Ejp1nM+fN5Q9jXSKxz3J+QM8Y0aun3Ivj
lYavMXr3ymPqhwQm7dNlmCGmj+vnEQ9dNM2Rq9opHIxh9fF/wr9jEyggIfHXcAKC
GpZAuvQYzuCcZSQ1ie9VAkMQODE0/nzbSFuuE56Dbv574Yqi1XeUg4CU/Q43r/QD
menXX9qx4y26c4gMCFtjGvswFtAZ5okDTtZj3rx2DWJJBHJ/1Dopqly5quooB2YG
tNzHmm0qPi/ZOY26r2RkjaEvT3+shlg8bxr80rDGH6CivHEedt6zVv9YpWXUsSr7
8FjsofO3EOoxRtltDgsUw0JoMIe687dOhauAKRQi01+07HMHjCoGWMzN3lSebk8h
PPuLVZYWIpjyLc5bnQBlNboKbJ5wCO94Bf7EKZI4Q1oWYAoRNSWtLv9Rbe83FWt8
VeJCZlRY2/iK816LPGp2VC/x9A0MoFJCalUCYAL+S2PTZOXSJizOfrfL3+vymLXJ
t7Am108DadR9Zn2sSZYuEElngCQKsUWaGvBuFD0U0vTraZzSvb1YImd9lI5TBeZs
VjEAGxKzL/0mB/qf4Nut1b/3iQ6S1OYAoDgSX78ssP/kYsss4DljjdSK8tFCLve9
iVr3tLyCk8q210v3LpFY2oHLBxmeDtzPV7Nk0NtSvxFN1X9+ldi/qLGpPxtqsqp2
mWRUUIILb+7pVbYkVXK4ncXuIADuk7i0zhF52jZmUGn8/gnOykesD9+P5a6XvB7l
PJCe1s6Iwwf1u9VYF1E12KNKGhl5rFmxgCVsOzDeNQfJZW/YicxnCQWE6TcM56T7
6OiY4VLN6MFxbqo/iRJgz4EvmX+zZZDzcc7Uj6vaY/UxSWhruaoJwD05frakMDyX
OzgA+UosfsRysgJ0Q5GTKGlS2YvYYtzcOiUpqi1FHLZTN17UrmZxs2lp3UZ6vt+Q
358gpNVRio4z/YWe17tpxYN4uACaMVA7EP4uWxw+Fd0AyPuVmwGcKALrmBasK06w
Kq3RkLIS0bgloKUQOzl9ZPE/UP1zh1ftEbURnOAKCG9TN04E5VuzdSfP5FKr2M7u
x9DXeLfe45i9dFuP/4P5lveWq4sEURImnIPyxQAxMjNaVFyDwFBimDNGFvzjMv2R
6BcACUN3SJR548WnpEPAM0dLBnPLvksrDX/D13nmSll9py82v2TXkHMfYgAjhhxU
wY7Jb18YBPtyEUlkoyPQJiImro1jCu0nj3n2C5mQh2NJ/5GB8WK4oQ0+0gc3U2q4
4OUkX5+IoejJUBZstglLiisKS/AW7O0AhIVG1iC7AOnmks9HF6ncq11MDfl43GG2
VHN37sBKd5aZz0wGEg6yOEqYKpMBbnB39I2i8TndrDdDPxC53ApzyJYb2u53f7TC
CxR7tkzQkZHCq4TrppDy7gJm2T4vy14FnLJB2yJiwvmlsiP22cLXe35jqin/hp8S
bVnM66geq606MOMoAuM4Fngn6zknMewXef5w9HXdw2Eow50PLQ8iRgkMawDIzSWd
iSdzfQJm+r6E39cCPFiIh2un9JMs0/+/a5OBZICcjudzpmhlG7DlQqSE1gl+sh4O
JDn3JSu251/lyZVFq1UuxSDugA5DCc3gLPEwh/yswPCNzsix42HMMlrDDadgcJWW
bc22lULa3DVWZIyKZRS/Knf3g7U2yCLuc40uDTnXTKEHc53uPW8SfMhWcqPGUVFM
2z+TWkILwu+G1HbzZSlnBOzZr8T7AIDA1U+Ga8aR60yWNhLF+Sxz1kdjUWzCC6l7
Du9wesJWNwD1/Je4Os+y4+x9OBGwsX0hntRhYGEz6GLtnT0D7XnqOPH4Matshfoz
PvcOTYxmUnVhu9+eUuhK6DbvABmLujXUspvcfpy5R54QZOkojQIiwENNAZI7k4yr
9eVMa9zgNH35z1lybYif6ICRIV+pA3FtBWHhXeVfOqUvIQVcu3zAsLs3WcoD1sJ6
cgxWUvk9e761Eb3/d90RcvM4bVCa2Um+LxQH7JocJ80zFtpx8VwHlYQoB9eZKk4A
SvTFkmBdp1/nPp9F0ErrhjR0Nx0KUcG13REdMBOdQVASfq81u9Nkm57zWztuIKMC
HsrYKAwIff+FDwW6adur6yRjWppaYZz11Kk+BwcIEEYd69QYg+awBWdL0EZqRtMM
XMpwIjM/tlNSlm2GRZmk7lJmB729F8Tf+fw7zRZL7WUSUBDRSmkpQhaVyDISYbZE
ruIQtL4WNCMt/+MGQ+s3SocbUomUHZu+saY6enK19REWOyHoDhQwNulfqgeqxN4y
T6MjILmw0TxpeouiwvOKm5fnFDZj6+k59VHQv8D5wjck92OCuC6lFUja7otgevNH
Tcuzg1VIp1UOBoGt8Ln6xBksrNL5ZrpjlCZXXvaxmY+4OHNkXVT5XDZ4eeZhX4Zi
hBkbYukDyNC/Ujc358PNrEI4yy3NwEqY3p9Jry2RRAEhwb3bn+TmuVbYPdSKLESd
H8X1AXwnsXOQ49tH5n3+a6+X534f6I52LNhUfnm6yJz7Ab3D4paRz+RpmEUWr7Rg
tWwnX6eT35KLOAASE9KVgtUUFido7Xld/7F19D6rXI4qzmd5OX7mbyj+px00A2mD
1CPGYTPF8VfDeuQoTpNgrmGdeyE/F7kkrLnKPYhe2xkWbZuitbcl+2QqDuUOPXbW
GEQ+Fbnjglnpe3bmPFrbAiK9h8vDq+wAQBpf95dw4Up2wfS308bf5cfsfOWkYvVW
F70XH5znY8NuXmZ/iJF6gNXGlMhMRzvcE4m6//JVZ04RS4YA8IzXrY6Xd2Hqku1y
+vbB7g7PuT+hHF0IyykM6psBqM0xCJBdxuqziWM/KRJGQKGRcuFFjrBZbVH4bhuI
f2NrSQMvYsz75LkUezIs9OTID0EsqhUStLBdj0ZwFosE0u8PZd0TeEGYpNLtE1w4
jM3pXPC8mITY1BUQbQ3uXL2uwYgBlWMYnc+UHNXuuLC+Rq//p+D4STFeQagl/vAT
3OMGd3AvbG24CnuiyhLoldsEipozZSjpFHmAkETjY2+sa+gcePLcWiQW4qo3P1lm
aB7RTYGH7mM7VzZpmFFFAtlO6bnDlVKjHnAAbYTS7BqV328oDXkJ46MBi+ylin/T
taN1B9wP1n/wrJz2KOL4TbsQtPFM1aiWFGXdvUM8vU7xSJ1B9dUGDmwucGTI0sgL
WwnBIQPOByBpLvBnsJTFmlnDBjYL5BQl9zvscLgGbSk4rYTCRFfqiLHJkNWzfNGx
fH9mge486oBjaN4VeqQuSjIEuqmw8rGbJB36h7hpRQJeRZ48mJxMiQeTetIrQxpp
HysrbLsvWM6lSz69jVHiz2L1VvmQUOe9TOh+1n2VbHWqBr86lOvafePrkQJfITqc
xbH0O5dN/iejKzrWlvZelQR/+TZcgpNrPi+2p4UHcd+amsxIUwL/Gw7olFkPgPKX
tWW7G/CRrwAkjmELSfJ1DdFynyQRXkkkf9/nXJn/PvEdUY+0JTl9jf2LuyPoCC0l
jpvoYHUwFdyN4vlPQXH27+nN3+fmK4PuWBriUhOmHKKOGpBN0OzJ62tAC4AvC9vx
QqpfhrMh2FZtEkO6SwFDxmSPwWntJkxvt+zQ3klxGuYbsvJ5K94HD21Sh1KNQ8zA
g7lSegege0x4oitJamqqkBqum3aEEtKrpOP+DgVzJ7u7AsU8Xk61LzyDoASsqbU1
yDvFUfZKwCGUy1hl8V4UBGhlHX9yl8zHdAszQlLFc5KXnuErhddf8bBk/FudizIt
MEGekopYZEpjwKu0Vggvvgbw0BP6xz/+qwKNmabq55rVL1YXsE07h5zFT5NLuTFF
I7gdbTSQQs0yz37pDS32kJLBkjJWvcbb1+CwlWPBADVlg+VqZGtCOrlEgKkKIe3m
eGrQ9BcVcKGGoeTYjXje0yxjhFAmUBAxIffXJ5HAHCvl4ftdva2I+qCZJTNLtzZ+
aRoahoH/ao+vooBK36EDLev5wQcaPCKdT7k6/LMirGsw6BCzUl54S/MCHuWxq6jS
AsZb2uDxWXKQtIaQ6dgu6d+ekmHgLEBXk/4RgBlCh+EfNrSlV2IAfMVQAo20tzfG
/K0FmDHyCY0zX19bZEBIQAGUgWxQ/xeD8V/s+xXSauI23JTsO2X2OPQNGpocxhbX
nueg4Op+gmYwSMOlrk344sqlnB/71lsaePKOsyCRnPcUm1/BnYsl580gYkPM5FKS
fSZZ8rCj8eX6if5KXwM4fGYyADa/GQ8bN4a5BH+wIOq41cgKqJEYEkQo3BcfwBF9
XUizkVE16bQjh9ilLbgTIR8zAYC/1fe8Yh19m3DDRlRjKJ4rfYKrvHQjdtWQeyAq
wh5h+Nd7C9Vbsm0LhazkHOIPh2EPKn9J2vQW14YzOl+OxLlBp5IBvZIFR4hipZs0
vBv/H27wEOzwQoZvoiArj8aa/q3U34pIVNynkfKSEQm/hrWJQ9A8+lA1z27slGSn
cSO2nAkdzXqHEXWY8wMrXgahWsXXiANHHJITp7r++51KHLV9l2JM915Nypyjx2np
XZfXwL+NyN1NuDXDYzM8TewNaI1iCd6NUhfVbpNXTtMGtHb1SbMr8Ut3Vo1sTCTe
VXNhCQDfHNHbjQJ0i6FfUf+zcA2mz93tEuaVgIoVjh8dsRNM12SqfdUMjMabTv3r
lNXVZsN1GY9ZxKK9L+/PEIA7r9NlsbO5m8iYceOIUOeJYuO0KjlzP/EEe4IHdktj
79ZGqicX0gZqxV/jaIC28BgEYBdC9gENYgdDutKSosxjPykeeHHhcNx+TIJSI645
ppynFMNlI92CeHEGi7PU7ZRVV5ulNXMZl+/QiGm/TL1t/yASh+ktcFWrFVkb0A3u
jinyTsmuzSM9Su7nF2n3tCSaxCpm6Jyu59WkZeTdB4dJnUc+sS+ap0lBdwTzliH3
Ve/nvR25nXyu03+3weL+42jnCU4B9u94PZxPS1YP+Ks7+AvMW+MUw3MyvZHETe+t
mDP8hxvfpIc8sN6Rqp54GZdoYnOzbLFtTAKV6/fa+/fNeRrZ8bfHBGsRPQ2gvzm3
LaUzwZpnfKrYhBeW6aEAlX+G37TNThHFc9nVJzXhC5ANy32Tc3xYAYZq3dLet/sH
58lP7JWnvVndWpc540ParFo2PNusFlPek9dnDXoM2NOo+BE1z2/FdTc+tx4ZK+0N
VLJ3VSmiQXqGQ53GkkZFCPyxcN7xnRdZjTy7WnbUOwGLCrw2yurXr/sAh6tMPeXf
4HXZZpV5NUlSEB56DpE64MT9IzLJKGaJRpiVEssWz9f4YEDU3XOd6G9+uqpkTeIf
9oESZmZyLoTaectbI0il4bFnkOXPvVSxh4RozS04azxI+NCN5U/Cr1GH2iVtr2E6
v2TFze/7F6SDyANQGBg7pxMtrOiSZacZozQVsnKgJVQLt2IqJ3CM4VqgwH0cCdjV
6MTA73uKHOjG29irICZurY+rPFYHOlZBaUfnsmX0TQsjayGU4MnjYyqQ7fEuI4pL
HA8fPI5WU/2NQkCuaNfSQA1KbX9lpvTEjDfOQlr99g6mZAvl+NWV/BrerpNzM24x
uT4oTZY/lytRQiwQXyBuQaIhvh0/oMJc06JMSbniDlLEFwXFXP/i71EqT2aQ1ZYW
Y6wV5ff9L+Ehw47Q7vumZLoqYgwWzphlUWWOJo0/akwLXQtkv7/BZGWaj3Pl00W5
HJK0VaHefRSr86gPt3DA65dq2IMA/KrMGbwyi9a9KuvJWmLlGsU5pdMZqQCJhC2B
wVAoGAeldmnBA9vzSiBHvoBaCoVDUT8FmLCnxMhrtt3fMyLkNDr1wSc7M2LpN4oa
GPCriyKjiqbOdhWJF4GV27Hmlu1ycuuIhLgp0NUsCJI2+hoKn9wrvs5AJXQ+BRsd
XalsZT1qr+QJqO5CcZSJTnaHW/Plwkdap/PKe9vnq8nYFahkbVfYrKBdSOZ0bBQ/
QLV0k97ZHyXRWj4hZs0KmSQj2iW9ETg/pEQovYMC4WETYUnFmNCNgfxFAw1eCehZ
7gyMgCLAnWF+yVHIGDhbAL2lmwsGnSyiswttMq8YblhJSv/hwmitjcZIzkw7seS0
QLuDFwlcZ/BKn64mSuxl4rOD5Z+6neroNNzWgJlzgA+nCm5TOpIuVAWzddFqPmJk
jIWOeOrZwK0Khf1DshtrhsE6Dmx14Qnzvfq/Z+rAXW6mBaJEixJYQzlMRbHIZj8l
2Br0Do7RiJPRP7fAAzEMGF+6aZNIhvdJyT2pIfKWKr12H/3GumLBSUxzwEo628DT
L6Ea84ddzLAY5CZXaaii7KHyRQKJmyubjDyBPYwYIVcQNIhf2q4FRG0ZI0enIjGC
gCK545idprLCAHTRXA3pmH3tuLwhJPYiIdA+xaAydHbtvNYrGQtLOTZ5Q0yOvD6P
QtvYfiz8dV8FjbAxEeT7MKdjBAWRHU2MW0+2rDldJsacezy+aIdKoYAzt6KmZKEm
zbxT7gpplljIOSmIk5ZBCnc/p9vmyTWTBeTqXjp9/UtYNfvAM7BQab7HFeK2NGdI
HCKFFE/iPm2/7Q3mUkrKBqaV6WMnTlPOponEFu9MbcvWxkZlEBdsV+kbEZj2h79F
eIT3LIXXpwLIvF0Vkv3TYqc+UvqmwWUyBZCSVi768CBzkt9Om8IZkRPnD289kUw0
s2SXdGkWfK0/GMA8MDP16DMEH0pfMX/lqnvLS0tWQmsBKKkdZqZpt97MEyYaZ1xM
BKBigLZAcuw2iIFtM1uUPdkdYPtkkiB8qg2tyRnQSC5o0pwWPtVnhXLaP0pzyL5Z
Q8cP7Gl5imP05GOW39jKxYSKBbc/zTf6EhbG7qz45/wu7HwEnxn/d7yMiIgbeXez
e9C/V/Mh4xgml0a3Sx6ZJ1e/vy/WJ3pBlDktmjJzn1xTdOkKqBx3dDJvzWvkG8di
6qo8E0Y/tsx3vWv5+9H8QZfsGeNdaf7W/YzvFCtf8edRzPJ9s+mZjs3rJ9XecNbX
jd2PIyinqDDu5T/N8aqBVCFHVxS2zTzz8SiId1Qy6uqoIJBLkcHwa5yC1za680rK
WBhJyTGu4ms3t0YyNTu7PIwJ3xNJoitr33wSrAeRWHOFlv8NsAi6aA6o5SXA+GbW
arOj9aOU+lAdJ4olOH03u/hcN6pGjENJs6hxLZ8rd+PbQH56kwVgajn3xuY7M970
PvySPruwYpeIW+q4VAR9YqGtayTuT1W+OZFny6g9RdjNzhop13nvcx9qQqBoofq7
pwB2FHoEWXEo4TQsn1GsQQM4P1q8sR4XUHY6xjjSTIA/5oGUlqgoMjULL08CYxdA
aHsXw+PDyymd5+pigyGjGz6sTi1ax8VGiNXs6DYNJj6dX0kSbXZCfloqXQltL/+n
v40Ws48plRbDg7PEAdCq87vr1eI7SmocIHgG4rFznaL3G9tvn3VtxAAp3yOHNOEK
4v/LoShcBI4uBO7SjRwyWbIVyqUSIy8UFyKJ4vSG/BeguF5ZF29JJLs5tfTYMhMy
19RXIpIEH98RzExZiXUIbjdgajbOywfE/E1+2KBob2/Nc7vzF3cgOw2O189xs9OD
IUsqQ0E3IH6n91T8x5GqyVcKsSy9UB0Soq85rTbrFZazb8Wetfdu4BxR3iEYITx0
7KvWqSuiZ/TQ16uKRvMrA1dfGBsRwDnT6MQ5eMJPFu2O4+T0Cht8hl5LM6FyLtGQ
D6m3MdV9JDaAusdVn6iO3f0MCPzBzTEa6o1523aV2aQLx21iQBfMKU6fvA7Yp26l
uMFbr5Uj5b+fidnoHvqwo94ApNfJRm8ouAmO/QZwZKrDuqsAZCmIJ7e0BuJz8bHO
K5VqlhrWTTPSdA33NJBDq4Dd9gEoi9BqlRunCOAC5e8wxCvXGcpWPsrz+vLl9oqk
pCJX9zdfmfaHn+gktjEeSbaxN6WlvkQYiEbAlIh4V2nkHREhM9qfF4R4A7CyCuC3
8/KQqzhRhpe3th9tayU/Y1ZMm2J16kvU8gEEhvyhUaY8hNEV3zM4wuk0THEJjWyv
PayFYRPkIJPzbJBcZYidI+lyfw/vRIH2OCUzzeFKj3eXYW/Z3lSyC7DW2JANU65H
Ew/3DMBPuByUo3bu42yYftWA12BhJnGhNj+P63wNPBYSXO+w3b+rZM96KZrkBvrq
7OF+hrpn3X8RarREZMa2h/5ysxN29F5rFhZlzFN56MVg+zb5PJIAfWo0GiCe46Yn
Vk6nBTBoictNcH4FD8EtE7FHUIPwhsyIWFfvBHV5paX/77AxehKj3QlMe9d6A1Ae
ADbrtsR2dU7XAYt4wTT6aK2hDbX1n/mjtb6k2kPYxGgrYEAxLwqVHmz7UCtx6VHr
XqXBACANXCf6jstmcQJQVbEQslN0ZVqEN5GiyJX8BjkC+deKScuI9pxjMIIEqopE
+iBEj6bNJNh9GNwy7Pp7VoHgcT+wm1+HQiFRFoh6DZHxYOS4zECNetWG7lA6K6Wb
rY6K9R0mF+rqar9mbDeuyqYzFSEPGgzPZAVOQV1CgoYNdu8IljwtuNzeNY71qC+a
kGflpPWsBd+FYc196YO6xcoxUp6unwaZA1FhfSC+H9g6sDqpMb6IK+LTkbnIBpv1
7M83H+IEX5GL0LwynSiZX/WhC7mAUvHWcDS48lm+X3AQvfQiqVkWRxM/mgPf8Tlp
Qmbiq2LStl5h2ydAkqrFT7Xv/KbGdreaNX6PXqK6/iRefi5Cu/+tLSUKvc3IoaKj
k3MrX5lX90AmvToRBwWukexV3C+D2Q0XwDDrdiqLlHKCx6epMQfWl/PPvxXQpDEJ
+O678hbVJE7/h14fxLg4tJdLswugKeEVOWXv12WFAv88GxFt6s41Z9vGr2DzeaLd
+6Cp4qRi9eMQqr6nRQqbcp7AC5LPrSOBid2uakdL1M+XaqRMq9u/eWLPScZoyDwj
RVgOiu5NK7h3FeWnO7lf5yHtOsBc2wtqtRs3iS7J5gfvL+L3qdLwsT8I3DZ5zSVD
KLSDeXZ5lEohvyGdR/HDL0lyipSDpFxO7HWRWy1kHs1tWEheuKu+OAtcX714x388
TD3OF17ArgHuiJKDU0uGgb6cGYfTg2X5tE9V2pRm2U5h4IwUAiwQNRUB99a1YVZp
9/4Y/Pv+N2icUDu4tiKFQ6tPjH4TnFK4N1QQqWmjpCu3cooULH1jAqvYNZLjFZ/2
Uf7wFhscptuNZMMNNiD0XcIPQRp/uXwANCyLIr2AvQwW/5fPt5puHwJkxLb3d14J
St0Wxm2gxD3CD2JWV+82ZfHLnlDGx0easoiOBuRZoMzFqiahrm9o9sTVl4UYHqHu
45JHxKIr0Cjc2N0kwfZ60zHPtLL9DlvEkQVrLEAudDPavaEVJBv/JiyiE4yP5Nj0
mwPCVhovm5edYFF/YE03wnRv1BM89Ak52it7HsUl423Rb2emBdStPQ+ob+GeMNoC
RVmuILyLMuF+6dSls+ywLX6wNELB/VEiBJV3cxLEi7nBquj3YzIHw0sxI+RdEgFD
7wqdpjcCiEBU82rJEp7kpfejovNYcF1EjPSw37koEfX8pC6jjwJQHwWNq1DWjHM3
BTRzVS3fmNRLGqeoO/dnbdZizgENT+PsslI7sj5GDqQwHGGGXbfwx4euoRb5OZq5
7ZdQZ9u6jwbcacKhonYDlD0SoUFaSVg69zpVVVEk7HytOf78mMOKpSq6Iy2Cj3T5
oTbaBCkg/Mgz5WUNDJcn4yJs2Yv0A+IJyT3E+ZyMCMG7+aFD6t9HryslWDDY9mx6
uT5TujROrPNCf8pOASraj2w5UZNFCJ7A6wjg1KuBpLDG8o9Gcqf9+wwmJOmbwssI
NkEahmr4OW7IPJ+viunWzGp36db2xBig5ehQYU6OliaeZtO/k7wSyx1FFx/AJGkV
czT3PI0IJ52vPszmd4NvSmqsEcxzntDYosVh5Opr5vO2UKsrAB7pIibE2MqWE0Wm
y6FBRT2SesbASmpcwFiai/riNYNnn0Xb4i0u0mL10QTMvjtApZD3YqdNL2+w94cs
W6XvEwGvEiML5ovTplIvJFheAX+jck4Nuc2uGgdjHT11xeDJ+fw1FTMDtwVaPhco
5EtIBTGMoQR58YonI7eLDF0zagR/gcFAzsuqJ4IlbE5O1I9nVwB/ZJmz0Ta/UcKp
m7B8mHlTjTlv/VI6jS8YFzAEpDMbnWqwM84pz9Rsy0OO8jZhAu9vMJBsL1q1EfTf
naTn1QBZ3IdUSMFeJa4NmOJw4//40NISE/OtIxlaJcH/s5/HLGtZwtC0vFQxDoAP
c8tSd8jjUMD+DAjEtkcqmLEit3RQHmeiJxyyCSMP0eoVGkkXjybY1mTguzYRSe/e
USK0r05FVny9Fw7Dp6On5MSI9FcF747bwG/rjOhWaLGA/Dc+6NaK6B/1CnKuftz8
xPAmJSwBysxIaQPevqCG/J11JfllN9eLUeJgRVYjLXVqxPlCEL3Sk/sEDG/tkAur
KNhdp4tNyYY5nI4aP1xuJaJhojUeNPN8XEP2HALhvFZZ3R9JxrAT8ruZUjWGoMfd
6QHR0GyF3CXIc01xb0be9aJsIhoeQTnWCRa3XeN4eHxEOfuzDS/B9launouxIo+X
Ck1iAlgUWN0Y/vvZJqGEWFJpiRZsIVXx6YyyEoXqnqcs+ObU4YA/g9FtAMZ0O3Qr
zFkMfOTOCMJ8X81uNF2ukCr3tH9TpoXiukT62rNz2nYrq+6dTwtRt0O6CUMtZce6
NmyJCaCT7zJm3b4H/jSK6RCDhoveqGO4q1SveN4mE/BNTIY+J6qgUe8QCQa+/Tdw
A3QYh4X9farbwpwZVkJZmlktpq7AvE+UR1irbXFVh7oaGLbeZgp3grqjJNFQ3tUI
VwqhbN3evlqjKfXZQKWUjcTD9ys7mHEQN/6rVHOkR6wRq/XPojGX5ncISEl5siit
NfGrOztZwhZuyymlpn4FEnAtQa2elf3lq4Eai51y32kjlbR1/NS+dRPanG1hrAAj
hblXSA2tNMVzImpFaPYMzS4RVj2raMhCkQ6vb+NY4P9qouwawOOE3CrVAM5R/DJ/
SPuOU3oBgv7XxNrsZTE44F3wUmafe9bg7kt8tFrATqWvGgUFjlnrcKfwf/KalLF0
RjQOB9eRcrREroVtajx3+LSYyFjE2YTWUrWCUs24OtXNpWwM9zMDqcXRQbGVhkVu
6QuE+aN5B1d4xXpnZ8DYmY2teLcjRSnWnProv1R72S203byPv/GllIUA5BvcT2Dh
kRrzRnQtRn9y4fIE/9SiCs2JRBlyLqnSodEdO0c3SUTSbA0t+WxKwggx8MvNFzYd
oSpDX8aQOv8ayXeSes08rHaiPbH8e+Wosx++B+Xb4+tM1y+VR/fPjQPjIHQUXMKo
OMG2HcuMkB031ee2U6liYxjCwpklCiRGPZahvJvuk5BWRqEjm+WZFEKtM+2OPmZu
9t/MwfCWh4rAH6U64HOha8gzemn4sYMEkgMANToYIovS/kHS28rTqmrhu0gRdWi1
MJkmOcsetb2KRSTF9741AJ6Sa5prpMA4skNmCRWhpkE7SSpsJ+3oV4h03aDpjRt3
SJ46lqKHI67n0c8cMBJjGC9mSRYOFxu8q/SM0poMbaFzlp/V3xD9Zdw5ID6Xv/kH
md1UeMy1oE9woofNIG3nOy1jDPO4+ALNoPvX7egOfhEsYoXgIEaCqaWc1RwOglJC
R5dnMGi/F1ZClHp/ZtigaZdliIZQ7q4x7nxDuvAHz9S0eJoIDeUMfC8lgQ0MEKup
tiy67K915xwHCRTWZ+7laUmp3wpnQ2f6xvxzAaLNHJ+8jwFepBy26jVJi9OfP9of
JkODN+TwW4//PwT82jSxMUl2CVNhSAcZwd+2VbV3nmR68Ql+W7D2bF5ZzyjhT/e5
AlxQXK66nuo7OrDtq3lWqHJklL5aVwIernAvkCPvnJFRqYXPv9iqHgcgVy5fEZVo
IquThgVvrx0Ase47Hm+CdVO4xxY9MVAq/Xv079K+Fi+Tfgz3gEcGqFonpdhGWA5N
LbHZC5Nh+iyumkvezSVndOPrMyfF3OgaVECH4t/2VEPuljJr8eYF2eTF7QDlzRXA
QR2RaV40JaumRPS+KTNVXfnwrqqgnoyeR7koxpY2bRi10oqpFHA45GFi1qonb3TQ
ZMdxS2KH11d+xzonpQPJnmH01TREGLwrzXImzowSjk3Ujg4J6WHeuvuaXIjW2laf
/x+tJQ9JNsMygW48kFdoyGSBouwgr1mpYd9JkK/3cIuIgzvc1XUEg9XyXf8+evNx
yX7X9s5X/FUXLQxJVt8T6ERemwL3lmoWyqbJ8nbdASYrmJbP0T+DFiErybS8tQaq
wsbypVAr95u5rYdo8fY6Qunwwkj4EMWMtFE3rn7OMv9+Q5kzy98BGNmOmyHaCe+2
lVLyacmpWNX9Fhz12rK6OCWwi7ieqGhVdv6ehrIWp0ZwgELPqY0816rIiw67L930
gq5yA2n5/iDbdW1PUcb1HNnJr+GZqGXOmvIbuKMrFyHQsRJxwJ4TrbcYXY8D8E+W
40hwutDK/shtMNHGbeKTvO0JvtGTtWGYnAVWUvlWQGxZUjvXbYfHElgAKuPKCbEb
Cymj8zhKxCrl93YyDZnk2k87VHkFF2h0m2FODaHou6OWJK5lPdN6c4RwYXQkZlDs
pAskd8myyQPy8nbiE+5Zn/5fYbiS6I1tUCYcB7LVBkwr0TaNmigSePylnY6iYvmr
veoE/t6lpJXBItgImcSB5YmDlosqiq8hqSvjffzmcFwtG+UGq+g3fbmlclQxtSbW
yLun5j4SjYWs1bxpUt0wyVk3WeATItWA73wKlfJOkGWM+ZWXjlUXiNnmzj/5keJg
PJuymr3YgZaBUaj1M2Lw187EHYmpJUM7SXiMq2vr2wQ4zf+GB31qySzSbw9rBK3x
G71961mvKk+SJJAD0RBw2/KnOdChWQKE6+l5zAxSa+hxPNU7Gyid3UHWWu3vIvS4
0fmhKA6Bo9AvutHh42JdDgW7nPPTBAlpTsi3OePOZpPzRmIVmQs7+eWB6rTDtcWd
dwa+hTD+1V0IZQ3kpcP8mXc7BTJbtHgHgbUxh4S7ONMPl43Se0H5HBGpHMlzfxE2
Y9PVuAF17kqze/T28/0bBmfCn5Obj4vkm9BwnCtt7+xRFxrJIcnjoEIy+GwhTQ+K
NAhOkxWSLN+B4+f2A2/w1plSBm9SE3vuOtFJcW7UqhEH2lFDUjy/cinEItv+UxPT
8X9vK9Q6Wbsq8VQ/lPhV+UFS4FK5zr/Uityu95rtmJI01V0E+TJALzKiSMKC84h4
G+VtFl5p7uBYSoSnDLYKVCUqHfqyw9Oizjq3jLvsfsLEsNcLelPRqr/WyvxRL5jm
fx9K4ozQVce4Rse5vvhO9rc0msNJZBaeJ7KC8DwS6R1TExwk305HcXmAXQog23zP
aB9xuG+Zxhc/qu3X7gJ7Dbm1DOm1V2nyokajFhF/lSC3BMZZ9PE768HoLq/Ga1aS
XeGxeD+JHfuNQFhc/FDvHl6mscLkWA9WiQQL62VWTwHCIgR9+mZ17PZf/tnVwSSq
nrxT0fvPm9SLZEXr4Q1ektslt9TyYzyfJq4VDmmFFeOJ5avyL1hmowuFiRuWi0e1
atO4TY2HM+1LnYKqTBD3dbFI9T231KybG+QKyWXLxK15GRAJkFdXcNO/PBMPgTzG
RlDW3fCS7qBIRMlXzglAwBHsmDaLzLj5aUZK+6GeiSRu51b5MRmTwHitP7tuiHC7
xQY4jxyAi1TyWdRoyp4/UMIxZKjIAUEQj91p6S0XctjwL5cdL7ixABXHD0fFEHnQ
ykY9AzBB1eCU3ydX17UChC8+Sz5NqezChs+FkqhhRlSPLqmz11gwyxdUY+facssN
OqpJr4eg1j3eBR5gHjFgY2x0UWVBiH5KZPmw4MP/wzHA+m6yaazDCgWiNQRjXrig
2mwqj/VEi9mktq6EPJTL7XKatFA00aGbVQ2Syqex6DwS//RrfkvdQIBDUu4gCENn
ZoYw/z4Whx7XFx8WHOdC752TGZdfgfG5B2njbHDbhVIELmUQDBdCkdDVwoCCGp7x
9vNew0uFXMAiuzx9Kxj84eFX9p3K1Wq0oP//OJiVjFQhUI4W9pyyrP/aLqeKVmeQ
p9ZodwQivMD6rwyeCy6RRdDC0DEHjT9GWrjy1LAMGWomEJYQXcEwb2KrORrOxQV+
9S051frMXlm2WyNnrRw1BwKGTexfhwyJm9q/Vg+m3cRTM5AGrvqP0372loJiyOZy
jDd/lYvWjOdtKtfVdVoDACj91Id7Qg62ElG3KXj0Ypw/XzPmQNPNb+JCILqg5LF+
KK4+JlbEz5pgh6oYTr4JGbKOs87PhNGVx7E9fxOUbQ1ei6mawT/40xIbIr3J2S61
+HuOIc2cV3gK/Y6U7cuIcYY+WWwYt1wjmboGIVZpM6dj9CYNxFCe2Vpqx5V6RKx0
mBZVr/KCGn26WNkGjWGhjDTF9xww/HuTv3xgZlTe/YCxL9zVFDLspuetu+/PiMvA
t+stUWARj/M05AtHieDg7EVEqQ14cQm0mEMjf4u1FAGAsGCmZ9nz0ZfzlT1f+BfR
0qaE0S1RF2oCrlx6XFA9RPRnFyBiJ/BcNsIJd+wud3P6HfvLyG/hNuOpJcDBMeN3
bJZvEFxtEmvAUER2DJgdByao8tX1wCw772e/20JrE68iwMTsieu4NhEM4v4SS2jg
L2rqVcLahLRCXOqNQ2bnXdUcanN2h430ofKRWoo8R6oRj0QSt7inyxIZ03U2Lufh
bV5sv6LWQvgkle+kLlHZl4xtMz66em+PIL1D78/JdLosEc7UpganWkLEdsZP5FZe
73eSQUoLpMANjkqBQfsccqshIx1u1BjApS7M1QIempFtxeq352gj1y3ZIEAkfTe5
TUaAVbB/AztPlZIW9EvLsuQdK69JgtV5OsuR86aN11A77xPPjRMp+JbIFk7l1toS
0pLVVHcTK3txFf88AllRZihRB/Tq6qhlhRsBVNcahLRSegYg5BCYhcUQgOrRoVIw
RBex/64TaE0VwaPiNiYFzGaKyiZLjJ1vCTSCXOvk7BziSAtmho/ZcloBTMHPWR6/
65bkHSxaQdmJobX2fX8x+0SambyZ+EJIykc5Xq5pffsQjIACTFDTZcP3YDvD8WQa
EbKyLr185eNcVDA/q+sFFuGoZqdETE16wVklNO//NdUCTabo8pmptgp4BM6uYQ90
cWoSB0b7Crm3kZn5HX9HaHDJo/JhSbNSIZiP1iTIoiI1+pfq1khOR6mST6o/WqBg
nOLVD35jWGSUx16GwUhoRuedEqgb074IHEX6SYOcqHMogVW8gae9mwjTx5EDhjhS
9Wi+Ibmy+wcb5P98bbjsRb5le9SX7msFw16ywk7ZH/TBWOG5KD8kb8GmaJsiaBf0
B6DVUfRsLJIZ32P5aUOBdtAbQbgDIDvAlMXS5lInk4U8Do755NJoqcmcyL2OKyRE
trRro6u11Z7aafeQUVtzTk4ombYTVe7NHSaXS3xPvTwZFyOIhZJpmIeq6cTyKRSv
HR5+jRC7jUm39PdiroWRdFEL+ntdC/YZg45cCgfWpaBTD+0sG/ILlSENeg522Gfy
UuzNmYSktx9OTIT6YLwbhVICmhjUoXpPlc/aIBiJzHRNL+JFMdpbC00y3zmkYLqF
ITSACUpTMwHATScI2KRjTheub0bGdv82e3mtgSqfsWkG2mXQzWpat5n3gGXQMf7F
v9nYYbAmnBlbBVaVRzF9V8oZqFHHtmHz0L3NusRUaZDlCzOZ4AWAjczNpuEM9aWJ
7QxABNmhLKaD1vYMsuPNtqw775NLYL3Xp9RypEOV9aBtJ1lfHE/9b6jhbpv1xYvR
Tel8PioYzi+d9PuU8P7zUYvAT/eK+bjO6Bue0dVI0mEB3p6tzude5AqTTHcF5tdH
Fu7IhY/32OK5t1bp8GK/ldgvLxYYbH2vji5DwW2LBKcaRjUt3LlWnrZZAFDCq28c
6T/jGWcyS2end16RbjjVv+SJtxA3QgsYGcG2FvOoo0g/cvtGzxRvNEUXGgy51LiX
7s6WPA4aO9NKG+sq//mfbm4n2BQsuLDaV9oSsjs+ruYRKNwyzVSf5wj+lZ5N6YUL
9VEfEFUOoIo7F4/1Y/HDIQrFk0ybyimSTD0LLtZaWAmk3m9vwQ6me0V5GAgNrRlQ
gvV1pbg/iKF/z6ge78SEvJLyQjt0vzq1ZczJTFRc7jfLf8yyK4tqOZC7RogbfMg6
ofm0WK0pp+uze41JxNiK4OUnReOp412fl1YBhYmN9qCQg4FVBNeZwQymaL02h2pm
HWKgwE8N8rjXQunLHR5o12PoVN/0VTUXfMwRPXLa788hHq+I3Ha+chjOJzEyYhYp
QShxAirWAvoyyMtI4z71un9jRpzk4uPgJfHrr20etNG70JfzqIGpgkCPNUNr6o9K
PWgbfwtWVB1Tq9jvuGl/zZb+nKoiWL3S4N6eaGQ4n6wye+dkKaa/l3mD5Iihae8J
8jNZNTxs3PYKfmzu1encuBU0/27fwWfP6Xt66Jckima08+XjEH9lSh5w24MbC/dS
PcdXshDln7Ni3qtkOuytK3WHmyQsa+3CyFeQqv1jkhMJ4pk69AbplT9WpJzKgXKK
89S6sEoptRhwypSK9bPDfEFX4s8gBV5HPrgUGanPxUPkWKgHF6W/+dqGMAS4kAEV
Zs8/uzyP7H0Fk3LjR7k93KwYTFUQrwi7Kg3Rx6KQq0DkIvP+XrsJ1f2AAmipyyUj
ovpNGNk7qyDRZBVUNf6FFMtdlwYUeFEF0pBuE9WBSjmYChOU1epI65fBb20U/oUI
l/+ps7Pa+mGMUa05XAXsSSX3uBM/ILGbNH0b+7mdNlDzioUXY44HGCN5I2Sm4A3K
Sjm0bXOR0PSkEQNnovqaPyLwjFky5fXIeNed9ssbXuc9CBlqxSRKa8ef/MMcuD4h
ZLjGTD9DHvlh10hLCp6NMN4ZUxh1oiMMU5RCVaTyRLtKzjNf0t0Qd41cNbbmf4ZY
a7Ezd6UBdXG/r9EDUidILAgEzkYcpvrcDWd3B74jUP7B5fNqnSo0jpph3tKWUQzS
yD7CpXoQbT2M1+6r9eltIZAyWMIcAlA2w7SGp8X0kINZH7pwKoLT91L+pZ0hLGMU
dmQm6lmCoxRnBKlbx1jVl2oPmr0egrVNY/2rdsKUoLHPFUOfxHQ0SlPYH0rq57xT
vHtZVaimowEj/xMji/oNi9zoVpDw/GAgmkFamz7aK64fthOIGJf1zvNs78o6geHi
L7et/HktHou2oZkrduPfGcngxUuyXDRsqpXVPFlo222CAK9VvxTLNRqrnuXFOWN7
HLhuPbMF/MfKVAd49JIz8qRDXTE8ZArfdKrrXeMJx6cSC0w+AVVZVrVhVljAu1zb
flAjUmIRX/84N5yCqSqGmK9ZtvJl6qPcfoRnouSB4pOlizrlyTAsFeWZhw34nqlM
aPLGh0xy9XI2Hk8l5R1rr5r6FIYxmq0LsCqe2kMnzJLg3ScBklYmEx/weiCin6ig
pRbhwsz9OulQ5Z0jcUuQAl6nU+fIf1bOkwSf7WwzpzdBY5RTLfVOJYIEpT5v6SAU
exmUJGoWAL1t9oejrnx5AkC113nJYOTAl2KmFvbg69qdwzkjUwy2WPHerR9YOo6U
g9P1Tbs6s86AZ3dm1FgBMnq7MN4Z/91UhY093mujvm+4ZA/Rd2C7T9GpwljVLR8w
YKBHCdEwZS3IWJ52C9YozJGCVYakoCNFjcegPpt7+vkKS5XJ7VZsACI17qeoHhsU
32Q2kyUGvQ05FBH9HIH4MhAM1JRbkJwcXVaqXhXzGXuGGmf5sC8/YWJ6StcIpkGn
yNbi1E0LS7KQOmlUE5d8poALJ3mvUIJIHVV8BtnCNGU2Y+bOkCdcZdHGTPW0/xGP
NkETV0XaeUr9RLXkE9AWlY16BzrFprC7qnmzTCr27U79h/di4xTzmkNz5yhDr5Qx
dd+k7o3hrmad7M3U+Wm+HWpfGU0O4oKQdf00Wc7iWVqZeQl5EAaW/Ts7THNxIIEY
EiFhoaOBWF/UxOfPgdyIU9H6BqhOAym+7rcnDQYgiakoPLZ37WfIwv5OA/bkYw6x
kg6Vs+sGsIXz1FdoIirAM6ZN8nBclYjUbQcTnR+36XEkfYd5Qe7Nym+OZHqdVbQu
WroVHCCcm7FfH1cjTLX6pcSODgb3kqiu6Tfm3yoMZ9rufDxVDqcv5Tf1h8rVvIdo
3EGEf6P0pakmB1QYuZcor40GVthXfp6rqMk6fj3lFJA1lqsG4IAH+SAIGfiHCVR6
iilmDXIbLeXvwKT+PYtqLBolF4EQj09NCnGn/alaxys/hi+IENScmSDCl3FIQza7
hWwJiC6KEgFnN3UC9VddRvTaoLjytKGKe0Yio1hIylX0/pmCC5yjO2WwxZqHLgnR
bUGvg1O1O/6I6OlFnBZ35R71DSTXU75IT+pamt2vwvnJ4knNt2+IWzpG7345gboV
VSM6jGuDf9I5kTluEqjZtjbBZF6bqiHZeMan6LmHHdwaAF4hfCKjgf8UemcygGB9
MS7YhS23dJaa6tnfsrFJdGXbTmTSNocDs51hsH5ldUWiUtpkE9eXZOAfpJ9IITg0
86dFKWscWcHMYsEkMDMe0EO5hl9F36RnLkhyV8p38Ls48H/YYsLi05NnEZ9vocon
HpTcFGrNFmcm42ihss/AtMdztI4xposv3z02PE7Vb3t4zjCUUSdkg6H48qogS9IJ
eE5NFIfKRTK1UmlD9/n9gZKB3hz5NBnsbKG4f2XuDyIBtDk4QjYgwhwnoCRPm7Yl
eec+WxG4OgglN57GpV8PyPAD/DL8abetLYda2aC5Ga8duKuB0Pzgg1NcdluKDR6v
MrsPM4HJKYXJ3uevgoTartm3tfQctBKPtUdoFetEoPi49NP2y6nLoTBIhKaKjdmI
n7eeYKuhFHT+CmRB36ivB3oK4ADFhyZP1XYvc18oD72kz7sgve2cqhjc41DeUy/V
RdKWqAvk82LxwpX8Jfgvr52DBCVUK91piz7p8qmjTby2XTN92ZSlijBSo4Z5heaJ
5xE4502Yar1EGiql3cvbd1W/AUmCpTOPGs1aPuPlOe5npoTpVrGVdOEJ75UQDYh3
KC2uzVt3nCZZ+Ou0U8B81bwfguJ9acCTPy2FkFO7BlsdZ2arZqa2LJTkwQDi9jmN
CT/Zq3i+wxLqFynCnLGPQhXdswFj4oc+fNkEAWaUcQKWY/nuyEhOMJWOIyOaw7bS
u12YOv5NrkTKWKdlsAkI1gEryetbWDXgXChnXJ7PYYRG/BA0hgKe8o68epedodZH
UM3XcLuF+nBZml4Edgy6sFPLTDA4m/stDZqy33xLcaOidRQEzKi4mC5thH/mS7qd
R52Ft5R0cfqtzjDd27XsJOX9FbSLpghLDJnMTcWAKdz2jdSExZKn52SHaQAAmbx3
gKy3qn+cM6Ewon5D3n5qKMV1AkfBpV7Y10lQ8rUKKjfn/toHK7y5BYnLfUaaqSro
dDNXSbxbfuV5od8tLl5VR5Y3pKpLsDT1+Kx+RPrwxPmjNAItzMHxuBdqIuA2a/JZ
WLasyi98qhkplszOnZDCJoUAG+VBnYj/WeLOFFyzdXi5KB62rPWYSTjceraEGEm7
CrQMgAo4PtvTjpNZPBFDV7xJRgisZ0xTYEZ9ionaD8wQY8qO8D2DButk3JazRuE8
necjTM7C4uIRFcUVUl3edrCifeEmOddlcko3/ossQR6HAOJfyIF3YuUlW8dPL6ad
HlTOpNOhJJxdN40cF385YU3XRWqZ1sxNxlGsYS/uBTSj5JfM6OyjBmcoYRrwA43t
WFBE9fuh8TC/nsmyiNJ6jRGj/OpN2SMp9Jqkz+TPirn/Ib3Vc271inHj5y7FPPkZ
wPYarMoI12cezMC7EbSka+2pZRuj6TGSokwIi8M6HnQBRGfm2cQaH+tyVERNF0r4
Khwl/Ah3K8CdsPi4vk5wHrId/oUS5XkjCZDeYcBo/DOWnd3ZV3WDSNlnZv3WxrmB
BC5DmuoEulGpA1OYhBliKmatdHWLH0jg79CG140YKM8EWXQYPC4QSfmoIUTCsuZH
TF+ZcL7Z9eSxW1bMoStW8YXo62YaPIWZmjfvRl+SLJHp1msTl2Yn+gLLlv9lBxzB
PrxmsH95J32YRGYjcmKPcumtorVYtZOWSmpf3s+vb7RY2yBkYH28F0402m5KG7bF
WjQsQs60Z3NNYExJNbYeFA8dPiVBoNBoS7/h+nTmtzbDn/r97gylUM4VqK5dywN0
uNsMBL+464lpPbkdX9McmkreuqxNnbF4Y/wUPGt0NnEWf1uC/Hq+svaLnBD1dVt+
EirFHFdPw+dxzKbL59+QbjuP/Ub9tacrdN8zWzgY4j8qWDKFrgFFqARS3KGSyiMT
tZKjI0ceQHnzDIMxkCw30N1QKp37RoJVXDRMTZ9pRIwLp8TYuNWkqagpGXwFzKqq
GkzcE72hy9va7WkiYJ8Few1tVpwc4HLoYCQybeD/oH2j/sXBGGj/T9YUDM1NtG1o
ld6zjUblFuegIQzW/91a35dcLVEsUl/clr4YOMCx9Lu8cMMRLTt2INz3K8VkRN9B
Sw9K6ylQx27IS7m9eVa5XumwHQ7nCQDl5NqX05pncqJ7+RmggZ+54upAXK6S3VLN
PKa1nWxP2V10G1FK3ST1TwHGshFR0dngfDauIGppKVH1LyyWdGZHEkaH+GgvuHk0
eJ4V3nM2b51fa593fctjhhH2NdF+XHsY1G0+nx4s1O7ZC/6PoedAzeL0vifNJdPj
PWTj6e0dtksNw2sRYutyVhS0b4jaFAUUSqyo8guNoRMh5Ev9Y8NQ6YMvkMwrjTde
25DUkkvYs5Zp3BSyYaQw5u5vN1TmzTg7RykMiuNQ/xpcFIWCflPME7GdQk0wScOd
Vvc2y5Kag1ecNIo3ZXqsQjbs/DauTC3tqJZBGcot67SQC96AnJU1XtDCQezdXXRz
kopVD7LQ5Alye8GhPaDxQS/cJDJkBdU8uvycYNyUhu61r3yVKO8TACCdEs584KuJ
u+7LjySYqKl75k5ruShCoKaTEdOGqsqfH59js/4lHZ14ndNNN39jxfncREqvPS5S
+PpPx+11QeZI/VXQqpHkUAR2qcxpV1kJOepd4QEwcGiScuaND5XEB0S/jacaN7tZ
PEAuCObHwrYETMWxyizJsmsO2fkV7HTInuP9X6Z0jZ9/V1Rvcktj91Q9/7TKOFl1
uKb45mW5O62U8UihvSvw9sKUPmODJn+zKhT95i2/tQ5CIJmIjVlLVellyfO4OkMF
e9e6pqRr/YQf4VTPNOTlW9YY2AkFJcjlj84RS0YyL92rrPaCE1lC++NzF2svngye
bm9fyBFz5913aIHlAbrSbPtAFKuHiC+XbX/XpT4czYxhz7jMB3iYCLyPC5jTCW1l
xnw6vRJWbts2trQ/sjnj3ozHjBo3/46QE5P/vUzta+rYy/o14k01wm7vJMP4bnpe
PHIVJUqc4LJrqKeMMMG+JyBAs6ScgTSYblLYLZBB9OTW16x5VZbvwAXHpW7p7/GD
0sVQF1nCNs3H0aeQ5cEoG+FbPpHpAGqWJ8fhscqPox+OQzW1ei+FDHtyKiMNcnwj
gmtXjigh824yjGr7r3bMxYwWuAGccFfUL/gGLwQEwOnyX9Tvrm08tXar3Va1aki7
D4ADc8Lx2jMCwPaeR7vWWjW1oaV4LdfDCBhrsYeNlh5j4LlhiDSXuj7jOw561Utg
IDCq2X0UBMTkCFMmvhhtMwAyNJM/tTZdoRRc35FGd6R5kpbpnRRohWmvy9Vsqu5y
tgomcKfxrVwo+Se+diTm4Me7HuL948xNJFrN3+VZRYt87KU5sUDUWAVkl9iy2foQ
QAar6gXp6fVojDm/GE0Q154aTWvTRYAbDcxRhqIpBrB30Hq5iZfH1iWWFM3wVizR
ur5moFCT0rXJgjso7gZYKE2y8557RtwYjV5OpbSN66ig0N4lumYkqUUJj0I0J9+2
Osg4mLp0xmvU4CdmKs82WeWm+Ec3U1VndfbHikYfBZjLfX6lOEXupOPHpoaGfhDU
QKvJiInAOb4vrrasU51qD6+CvtJFNavsiAxdZ6NjCXFEW8HjrEDVTI7Nt1MGh6Mk
Vvs1So6nwZ39E8WwCKJM1iF3P94FvLvBMCXV62yRleSjSHLXbqECDCXXQwL9MHkd
SRYsVWkKCjx7sphffk7taQdVW7A58bcWiZj4JxkY0Gh78vLN3k3ZCgVkMQnMmCMZ
9lyKoBIGb5m7mkuqb36HusklkMK5N+UUtb3EYjx1WtGwj/elDiV2QjunaRFbcDgn
cH+UhbBgxBeRmhhLOCvCyx28BqxrOY56jT0TqaZ7cCs8OVwUCRIfUTOQuaxROGTh
d3YGoS3CewW/ebGCsopdFijJG7J4ULyUf26nUAiz3uaQXJa3pZuWyGcHhWN308u6
vkaMXhyR0INn0dxaIks5uUrxMW9t9eqYlTLO+nBhWEqoQxpx7oa+RVy/Tpow1LE5
ICRcRhKhNiZ9PEuU3VgYG4Mwx/KouhoP45iFP4wdZcP1V1AYFP23oBqprFI9wo08
cP83Bu6IV25KjKy/8xAYyW246jciy2rEzPlb0ZdUjS/XXzFutV7azEQ0Kn4BbovL
/N8xGuCzg1gCpFDPMzlt9kdng5A5HuqQsUAj8P0faiSm7n6FK1KfgZauDB2QfU13
yV5tMzQXuzRUEaCvIjuKbY4Z/tK1iiKuLCGhNSzGQlMijAu7TFGJI5xKAiaSjjG4
uzr2iTqV2t+qP9onYL7lmnIkIy+3Y0rpdiopZE4tGiv7T6Tp0I8non/WL35tjMNO
LpQWycaSdOt13JaHOwjgtif3ZJr+9Gh44J5Andah6I6BDMtiVMceI/umDVTQwpLd
MVFz3ri2en8nLzPjPC0TVByqTymXjOSef4OKPEuVsmS7/iRk+wrIAfVnq3g65io9
OeDmk/Y6wcl4OrNP62Pb5Nc5af2MZ5Z9e7QYYWKVhiO/7Kd1/ikzJYrozE8He+Dg
9Mox6hRvTgElpE3Zj4O93gcs1FvaB3CkRNcNzFEpJu/X7/D/+S4xRSx7QLldRIAr
ufg4H6JEy4vUW5qS935C0LNTFRuj2iLmdie1sE4C/QV5ptXLyxZRzz1KPPKHr33g
KgSnTAa0BF1bwbVGQC4Bx/ORnRmF1KymCa8Km5YFioUoj3Bmh8XXgsKG6fn6DY8h
3VC/1o5q2/MrjcBp/U02zZRWU/HdyJplu3eD7MxfLR12QFomABHM0ktC/hR8UozY
F2MgYUy6AeaoukJ9CQlptiI3YsGYopT/Wy5SJf8jSHvB0vVdns0YHt/g94XyihKG
69dYMrwdMqF4WLb+GjGoFpTkd40MZG6l/ZFnxERQeHUcoGZsBa777PeAkQkaYtR8
czpD4cvEs3c93henmdDD/66a8RiYExopfCERoRKR6FIKJsXoS/+yDGDzXwiiWPdk
S8SAJFeDQycXCVwkeNGzDNafkWFHdg12RFebsWqONpjysZE5EmsOqYJ6n5RWaMGz
0tJPHoy39JsVkNg12QPLKW1tIItr4zpiktpGdGOILKAqQBiLBwGgYXX3KzoHWb2z
8KGp//AD9v7pBFDHT+UZDuphUaId97JWQt70A2QnHud9PMBUm2fSQvLsMW+aKwih
HRD4s8zEtmIPyd34gx7GXmpK/Ye75Re1liRvnJhxc4oojDiwZvXvOelzuX67869Z
SxgQc5kazgLKNqqRy7e1kCPHi+QSoDlQehcLSC1lhFhZSkutBLYcQ4qmAVT5wGG7
pK1IcAAiZH0gs10iR2JL/zPTnWIpGfTp6cmot07fmQxrLLH8UWJiEFZbn2X+7lI5
X7sJEjEbrInBm1GGvzh1TIqm5cwf38FXbOQfFORV/MhOyRPCW9u9kHlfwHJt051n
D+FRelIohJALaxg5MeFs29XfdNJ+HOhLGfVqyg6Ejlxo63kePmghS7J03faIeFIK
C741Q5bu8I2jBEYcNVN9oYTF59YfV4IWxXMBpdMdO74ddtjE4+qd2XFQoG70S49f
vg7iMxhkaLcz+aP2w64CKrTa7XnTC3QAgOfFGthqeqcp6TIQ1Pn3vFxQNKyKfgZK
PkrWHXt2utWw2g9f6uk0X4YIGwCXOrdh6CU2zkuMA0nAm/R75WxxaNPIZhmI9Had
Cma4oFoANgTr2NErm/LdxS+7iv+uUuOs5Awi+N7BEeEDMxDG356T7hd+jreSG6Fr
VxAotdGYJUM5jzoBG3jHoHXMaXx+IozuGw1EKaNE1ZfoWo6vMvsw/4qBP4vCq8HP
2LloSxwIjhBC1z6pLn+uBE7pAafZPIpNJ2JHitGqB6ZIsZlJUeOszRHlptVy7Ix3
kkRiGsW35BE/tmblMylFpCLw523Rt/xeBTx4mU6xIMQgnco3qkdyBVps4EvFj+t4
KTqNByOiSKrh4naZ1YsRHaVusxVf9gdSa6QcCz9/y0hhjW/sUKWTuQvpdsaObB/9
m5HY0jfoyV1hwhmVRr9nkiRvX30UyJojn+81bxYI2sZYYGlyIRUrAUPWwcijLIKD
CzB7Y352fnWWz0kueUGdmnZ7R9lT8mjnsKbG+SFvtJC4IFlFuxjREDn0LTLa4MyR
6XrTMsrWgSMfMCkZKdk5Tn9acuw+M35j9uW6QzUbYCkdmvT2p1jsL3VQbOErruaR
/8u3cTbUa7jZRB80+HDarV7AQpL8mQTNTRQd4EW28XizPNYnWBwVwKJ2kYsDp9bv
qcqbSL0FxlbxzGNnTP0dhOc+oryIGEM2aBnRpdHxPLdYK/RgYrNH3HjHJhzRmTrb
r0CtvnQ5WgY8Yp1IrHMp8FMQrsolmxUiV4ZPMZ+TUlCgAm4o20gNNcIL3qltedCD
F03YcgMqMYQi958wjYm5T+S1yHLAA22ZRRnGiib73dJOIj4ZYUhKYPa2GxYZZj+7
9cKMKwnLkrI32BUlyYNGgVUVsO9MKI5O5iSHEEC0ebvfM7bYv5bBJV0j0ozpIScq
BWdDfL0h9v41jy7M31ageIHzn736VBtGh4MfpgSxe4l1fLw14GsafdalQnejbkG0
ubVbAccdyPxCMxUumvI5ffmnYND9xoXVx0IpNcna/msCaDwO4JjaleE9e5XUWkhl
LVLjTr5LuWgmZSctNPy8Tmbj6nx1xyyPx3yxEVs73lxpZ8UV0gE7zPMHPaNNOReO
7bP3Ad4w3SF/U4iHX1pSWjmL4Ola8wIW/Boa/bQySoN8wf8X9FLvfeQIhm5VzrZ2
7o7TtFdk+r35o+MJqlQQdqtYzenuL/NZ/tXD+HrpdvlhM0GLIoBA8G7uD5NDnTkK
hwCbmwOWZ9nLSqkHq2r0G731e9gD4KrO2B7W3m0iJul/w63/EuwWR1/8VfdBuXXf
D2Qu44Q0z8gF1RwoJQTKgeLHhGGoI68QmE9Pnf/B5wJAOA8uM9oKDGGzx5nbU2dx
AZXAl1VckWbaiC2phHL7zQW4FGYBk/Q0Q8UWJu1Q3B2hP2tR62P0t/+qrqE9glxu
YJW12+TsVamFjd23Wm5RplJCM9TMX3gsdYgbTe8U8FNMhSBYplYTahbF0ruox8Jd
69ZPoStytrLnDrsLeza2J/DHIoZFzRxKc5odHc1gk+WTgm+bHhKHTgJI/pAFVtbq
1KLdF8pWJpC2oQGcy3kGRDruoXJr+Uu25aA02rHZMKpVf2FavMLoeuezcmQdidDs
ITMpvQub1rfwc1xl7LUF2ZdBdyHhCIO+d4rcvoxhWUfTJcA/oKY3ZGwrdh8y0JhL
Iosoh05yPWvljIsgN2dadR7mVxQQaP3pa9D+iGEecM6fvt69zNChHRjgMqtHunyW
oNjazoB1KKRfiOoGDE+3x/uTqa6Asxe/UKC+TN4Z9+QwXBrPOsXouv5NBMmDp7+J
X3lOyIaBWFz4WWEha7QbD9NlKmcQGJYmmZLBPBiFBW46IxDADAwab0PtvH45EdcT
jCrDBzrWBU7o0pMgvaXwbhjqQCy3/0sQM51iKQIxex+TRZ91WsiG4I0j6d0Uv0mc
GySudgdFWnMzVtAlkBC6QCpinl+h0cJMYGv4Nf8k6gimOh0wZuVznw0j5yv5Pxtg
IeQ7N+srWx7SF2Pd1hixLxqwHr8jhKnS9TqQeYXVAaI2pfpKZ0vexlu7mHOfytKJ
uGSeNTX4YQv/t0S/iODyZThnk+VNUq+69VcSeph04xpqk0IJwgYGW0BFwpn+dPfi
gkgbj/S9wQKmjFupjHaMbm6RBPxyur2F82pN2AzXoK+FUNhw1+0Do7v8FX719E/r
sT8IXAdu7rA8BVw0wG7pE2SqX0vD9G7270djGbnSD1SYWqQI8ngSz2HEa3ClEIu4
KXH63OSQhgq0+fKr8uss6NJNRhvmHgJ3w0EE9LRgXc+YMG0gi/n0QHcK4ENnlcE9
WPVKUriEcbfgiCWr+44QSCdU8lxt46SFUpgQpAqg60sQ0fnEsUGp/vWa57p9RVPD
uCdzN1xT5YsaJs4eVjm9RauyhpbygxFDaySbfbtiStRl8XBh9Atq9BxHlrmPS46T
5YfFtR6d2afK9DvIVctZmIMINaaZ9Tklo3nE0nXpVAQ8MbZOYZAnz1j/DslL3J3Y
WTEECEWT6loSj3TcqbsL3swEQcO8u20/Tr+zejHlR/UEX1DYRZEyR/ThANIlG6qS
6jSaVZhul8iMOT4UsHHU7E02dk5UV05uHTbylFsY3G3qR1P+8SGSPe89yPUu6kTc
NgYxyaE2O6otsRkrAheNrqPWSP7u5TRBgnXHBk9JsDmRnr6FDorua+leMa0mcgGZ
iDjr3cNR42sk5haPqGkDMm5IXxxIs2r8Pg6d6uBJf28CyKlMTsZgDF+r/GIfN5NA
An+k1TaI7ppAIIkTcwgJMfEFP3c9XKQdvvH9N7i/nY/zJM1/2eUOy9lJ8bGm57kQ
sO6Ct5yRQzflWlIPRtbwRTMvfzFDCtlxLLGaVxZ9gLQ/44Abk6wNfnrJRlLt3OTP
biD4qvuSMsEXh4Z1bLkTMPO2dI0T+8wIAMSyTRVIsZsM5cQpp0+VgZs4BxqATBDX
736q+tf8jzp2UgoGmYBIOjOMDX2Im3K7fQ76fg5Ke7l/FpJ3pmY1EkSJmHEy3bif
rwGgRC/WTLRLJAUrHQ7LRKcFSExxESZR7xYTBHx+Vra2O/9lfbQczgioQn8wMDF/
Jz9+vPf1AEOtyva2ez5usQSeOo3puqmrpogBjvmq605Qv8Jznpsn+JsKQCKCoHs0
rJGadYffBjz6o47usOKysaSBDd7Bk4qpQguq4diP6LdYF5zCvJ/a06M6LCD2nwtA
aY0Qxtet+C5TUTW1ySfim/OD5emWand/27cYw7Z9YrY+FuHjU2Bgtwf0KT1LNQK1
odNuP7B75fxBGNFpFPY6FVG9cOlmZG7k0SASYFRbD1aSCVSMzKhVPst0aUAQu8QJ
2ZvtwGCbIxPnpKy/UgBVvlx6R3iO6P2SNmRuPpaiZpJxIZzf/XBnjSDzg6S7Gknv
jzjehL+f4/STXIDBesJ7GuMbgdNEDkd7cc4kKHRJ3c33O3pJFLstrrsC3BZVIxT6
aqDwOimrRilhz4Z6CF/Uuo3vqMhJ67tie1v6TKjjE2tdT3kvNG9ygEoTbL8MWgU+
w+AUEtqGEZLoytEukYX0oCqOZPhini5yG5/xt0puITxNakvW+ERpl4K5qPySILTe
pJC3KHjjcGPF1zc5sSnXZgqrxe1lvlBC3WX1YKh9UCN//5kyP9uH+5BCTv+zep5V
mF4ij6fEoI3bXiWiOVHuQlL+yNpSCDQ9kq0VUUjN/x8kpqjFheG0T8OnTfqfAW8R
qmbtbF8CvNKUgFV2SImKm27h25p76DeIo0ksP7ILlJk3rJEfgcuA3uBhIaVv83uC
RGKAnZj9GoKl+s8BeV4UZ99PEkb8ksfXtmIHBZg6wdmdemwhYbyy+3mx2az1ZStb
VJv7CRUV2k0FROWKp7cdRIZ1zaR/1XGp6XKvs/vBvkmG+I8CIQpwUZuONbY2U5gQ
/rteEFfQ70vis/kWEJDdR0MHHENpLToXuU8Ewx3lTtoSSbfqkg3uZXMZRNueqthf
wkQltFNzDxE5E0VRQEoh7gpdGt89Fp0mm54z70RizLEg8AKOesjKPMawt2jI/oFQ
l1k5HMThBSGC9y91nz+vMk0yrAUmEv7VVEwB9UBEcSlclT3262FDTx5iGglkOStW
jcgQ6/EHcwlM/WDeLtHLhrsYvPlCqtfg4pN9OiePyVYi0JSmD5C/XsDUMEvOeKQF
X4obwW9gecnkBA55HuUZpz31aFeWPJ0VnRh/Qs70i5rdMzRQ4jFrpTneVYjkOzp1
9a1/oG9//hLj4QYJQPS42O7KhloyaD5H99CMS9BgdkQuoAMbcW9H5356tDEw/vjQ
eKYSmQwGog5lHgoGmOZILb2MkM5y1MvJxgFVc0VIi/bP6mJ5btTegtwTz847IqdC
FyjQkbNfTVyEfV5BiAsoD1vfRh40/dvxCh3ft9/izjG1HR3HTMnVbtIUcjgvMUJ3
aoIiIIOgHosiz6yIYSF3FKDr8Pl2HsQat9/D2zmlbxUjl9PJZyXhBq6examydIpP
G9iS+JIbbvipi9F8fkK0dvO/jtQfHUN8ELD8LwHnwc2+dopE5hzZ2lJl/IQlWzMb
uABDEIwi1Wvr9YJA+Ax0z0wFDY6BYMyOULpn1RaLA4InRR9c8iicjhWeqmenlVKN
i0TNHS3MpD3qxgkYr7CauRq6ll3BD2aasKfItZp2fwjxH+I5N+DebzQhXXe6ezny
ytlLicobK18kqBxsPzF+Z3jONQyCO+TtVpzCYnrYNuqEHYgDlO421jvmvOscRDvO
r9UrTND2Ntge6q/uSIyv39uTsjr4qKtNCcRXfSmETyMG46Q1klhoCEOoHySD/zcp
zAxpmBXNH+xV1UStY/lLmc3cQTOk+MdLQ1BqyUrakIdmybOKW4uBRXsCAUr+oT5N
zFVpBkR2DPZa+eDTzd5rAMSdHRkYWSuNQfNT4zBKK8WkEbYGj2n4pR/IIrN7CXM0
fZpxEuf1P7o1F0XbssI3C3Ws/Y0WtjsUjmaQ3qPcr5Esz7k2ht2EDolAm3d8m9n9
SVWg40TFgCPlpF7dWPrCJ6W7ElFIGOL77BBO2J+qpMif1Cz9NEUybdKqahR/COd0
4xGQEeqKdX+8e+LN8KfBVUyqa+I7G9KPW0ZN30p/xH5iPueX1Mci4PPTbJIYXu7t
wo0850Dgd7tsseMXggyziItJjiZGl4VPFk7rykeab/rxC0GU3OUpRV3aDv8CrBYa
sU1Sv1aveNvrZTCTyyxuzO9v5DkBj06QJVj5ztzT4ZBxaKwX4iBABEdmLH2cPhD+
q12Ev9jX4uEv/tB3/dORl0sDLxVZLYtsHZDpJjmxNeLmj4byKkcIl2fZsHyF0v8v
0l/0OsYkmiidPEU9vxiYVK2IYdcNpVI4TpDDSuROb3qwfQX07DYAs7Kem1UAH8qf
zgnzJhIMubpsA2/FjDViaTl29CFU+GNMj8ZOReCCO/keI5/vv3TDYjSd5rq10Z1b
oj7tu9qUxe1MHZCqq1D8CiwGH7NldbIP0uL9VxRMAemqDJ1Hi+ArRgdxBfXbx+r0
Furf6Ht72+IYH8ARkBMc5yHTIB/FKH5pGnkf1FVn46FTQ0BmhSwuJ/QPIps1DGv6
N+b3Mc7Dbfbjy9Mr0rAj7HHoSFr7JkZPONnJuLD2oOzPQrD7HVW1zb6b5FxrP9EQ
PEHFAATKjYBLRbkvSxgxIZa0aCl86XOlZiSbdvxaGjxfZwnXbdOPF6xMTzX9114d
ObcoLIwOmfuMNjJZ8rYOtmnTyBRlTeSIw1A6bRJ7cbzMT5OHnQI6/runjL2awhrA
bstTrXOEZZgZ1CoRlXTYPNeJC24bl4k5fI79xvqV3WsIpO5rYdVNzxonM/llHeAn
aKnP4J6qW5mWDg8nbkWCAtV2Kpk/NFmi8CeoIQ5yuiVQTD4Tvgut26ZbYL82wcsX
JrtYEzS/gaXrJSmB+DsB6+7bRb81V6LpSwrQpEbx5Fm1Ei6LF1ms7lUQjwEyLGmS
WQ9GtPQzqqcT35/nuvundy/AabjT9uXVdmBKNpJ8eqRsiY8mbJNGGZjyaqN0LTi0
xWQ1GIgzWJaqpcHe8mYFrmFV8b5dl6XycqJ2U8oRhls2zEDoraw32rT2E0kmqPk+
2wHL04BC5jIHcRLww35G35lvT49088OlLU5oYEjhdt3NrYeXgU9J/7CHJJyS+dkP
N9lvGME5x5kLysoa+S46AGF+dQPQMy8UOehO1PkTsCHADUNkQQs2z4AW6wGHyF3f
3Umx5neyhdwNzsyxyAdo773JobMAQbzQqFXyeFtiu96vXd6CbPW/2alBPMVY/hhH
oGHJrUTv5a4JHNAeT1BE4qHO4/NpPUdghDhGM1s1n5A5pvD99+2QYl++X7FxYTn9
oKbdIhd3soHFjMN1l0RAOcBs1LWS2A/N8cVx3cONaT5IlEjCearqE53bHBiMlVXm
DSwcl4u73JNblIt/84KPFIpxM6L6te6PLEPaRGH+9/1+9KvpDt3SckiWqZ5muwPR
lh+68ltgBuBc455zfVa+KWyFjcVsR9vuhgOrDbIQfORpD/ATyKF4SO01XNM2fz7F
f1l487HiAcVpHGVnIY3zavRlTxKfSRXuVREeyS719UcgALGYvRtAuIgl39pE9oNH
Kzhi28UrQ1OcWxDEos/Do21KDLmfzoSg6j/R1WFrKzXmuUYdiqK10DAJN30AzmRT
PtkUKDPv6bXFVs+WTH9654kMKChHu00KMyNRnRl/atalQe67uNZxH5gJmY4Iv9SE
Un6ouTCzA1h/Su+zkgbKX9AhFHhB+pWfJV79RMEQmLbc/8wfq4aixFW6JSMMXcoi
BvmOJeU3dEk+3KvOVcYJ6mhoHXelygMyBuUTmqvHUqlyV6sy3rTtLWTfWycVYOLN
1XFtBysi8tGieS1lWrfpU8ei5BQrDsCcU6u0wxkdINRbu4UY91Wfg7wSOUKxRDCM
yAP17dB18vRf4h0fpkCaRTQkISWA3wEpdzXD0UC6LLfJ2tC7ayv45V3MX7v8CDdP
ZO/gIb7niTFFJE6tZFvuqAFr5cRrIxe3wYGBJ3xcytiQfGaNXaPwoeKYjUOgGauc
gRFRKHV82Lvo32zH8sv/6LHiwdU/OLkPPwPFAn1sQ3TKGTA7HzKV4ifPFDcXqec+
BY9JmZopKMUjFJh05K9Qm+2oT0wezkEBf2RFWLpkyS2bs8JYTkFcyPsHO7gXopzT
Tm/OCSB7qv1zwVm38arivuOYMVNl5S6Vkz2zWtey/zrd+DAvnL+85jVyLXr1o0ID
6IrI3xbpih4dNm5SwdibmjSWL8kelkhEtSL/n5Ker3i7Hl2JQfS4SeuszwjPtU7U
ENsm1nD/WJheCmSFpQPNqdjzAv6G7uIcojofiVIS8LxtndpFdS6L2o7Ia7AHlEBk
IVVaRr7LmViepswZL3SwIetno219tDTiKoP8af3X0CIhNouJZmcXj4iqBDqizjF5
WTdXKknvplf5vflB+vuhC6PMoAU/X4BSi6/iLuSy+RP8apBVxZEJm55TN9aat61n
2oASZUABLNh3qOgma3SC/74vOvoJGRQINCiF4oU3tnfd87aX/JoDFr/goJMzIXCH
ojoKaZBRgE+fkJWghJNCGK/WyjgyZfPJO087lPt9MnR7vjurpECvFGasaSgd4m+Y
zoHfdTOzQvqL8eJ51MR60DXCtxSpCv0LxWVlry6obYF67Kf4iJzof/McZCw54qTy
5MHCMqwuhL6s1cJuZ1yt8hPW5biT+R+FgK+QBMldKN5xQOEobJxX0fL+D4af0/jW
uGLtk/5nkArtEfFSuTprSydQMSl1Av/A6wwZX1FtcVgeWBdBcrtgOD5kePwDmurp
/KN/hZ6lRM2rEexkn5n717Yf5IE100QFoYmVzTuulhi4sDHtftaMEW32pG35d1A0
ci255/KKrF8OF3DK2e4e8c9iUHFzOv8WlV86sin+XJrgpJbCbJQSDOh5OMdo9ezA
zlCm8Cq2UF63rNvb+slwsM6iL5FaL+Tp6feWUvZwewdvRNn+mdVY4rrAYLXOCH4T
M/f2m8Z06hj1LNsab+85Y0cY5q9R5l9Wjc3Bj2CUfY/4SdJxpL/h/urbhzjbdhhi
fN8KBgo1dZ+FZyIjOpbLFmTMq+n6gTq5VXqY1mGMpkmHsKX17BVsWqZ+234ZLf38
EBt4szUec6YP2u/uG3h6ha67PxgyMvyZNjIBbDC11D83+8fe2MkEO3LMcPN+I0WR
/IIvEK3dkIrG85T99ArUhYc+LqEHtDW8LlUHe9IfgXS6koPbLykTZnx4vT2uajfK
ARQVy3epGZ3MpP4oYJFQHmkrQHwqJBswIwazMIcaxB0f0WWjqPDgJM03PmgvjNi9
OHK1bbu7bDIToPqxtsASDIC4Eku5nOQQuygSAG4xxn2pujGCc1zcf1G2bqj/2RNc
LqKfEziqmfx2vOoIjKrvPKjZBf3CWB6GpbjcLfzM4Ml4ff6MdMlfLSWKnbgGOfnC
ZGENddKINispVbvCi1X51ap1ZeXhIi69D916qFOj+ZENco/H9m6PtGWyfFQeSJL4
W/bSNbfnpYgOyKVswu4BXCKuWT4uBPcTjIP9BVacsD4IMRMLZ8yY6EfClpdqQ/Nu
KPzo9RJSdSuo4qEoEym4Z+tHejgC3v8TWnr9dPwmuQbZtCbaNaqb2KHzyeAXwe9V
lYUnMHhdjUMIAmGdtu1lT2cYUCQe63j8djTiLJacIq7SiqgkLLmVP7sJ4o8QH7gU
ws7ZdkKeXkaYHvXGFWArk0/FCrTsTubEYP4l3xKRl66XYt3qx9Zv1ZLIsSwvKWiv
cvP52TZlXrmO3FFA08wskBA3l9ivR8Is3lrSG8iUTiP60E/CiFfLEDYBMEr5ZuWq
yB34kdjqFUTXZBkXSm3J0PlRmgPz4oMv0sH9uvFWtX7iD7jcU+ABJRyDvTPcLP4I
721us4C0L6/i8PCDqkdRNOz5oGeRq19hQskhfe7spoAIW1IoIcln7D6CiKj/BFhS
jI0sAiTu/FQoHOdvrhnwvy7GlOuGN10kWyzwpv0L4QVQNS6mGcUvPWip6WgDeLQs
WvkgoyRJftPFepXDPs1COHcfb13CKQTRYTcKGxSbcSWLqtB3O1+cbQthaLyGEXQQ
Ci6nL5ouKZz5PuRxGfdIFyco0Cxg4Ho9aX4CEcbFzQZpFDH3QGEmiNjQLNtA9Dxv
CLSGg5fNbd6DcM3nocjXhm2xNJEWhKadP//S5cSd0phtwV/UZhi2AIaishbmwkf0
ao3miQseq4S+gt8KYims2c56SoUxCYF65QdPizEZ9+KzN9qrhru5NKx68BP25glD
lwDeuanknnJqsKUSMKQ3Z3R3vk2Pk2kxBjienNohPxvrDp8uIagDkaGSjthTGPxW
jicwbmyH4oOMywE0oC1X7IIzr7+4Za0U1WHHlU7hnqC1ATm5c+aka3PaZmAtDs/g
4ij12EPpDrOThIQ0pjYw25cuRNSflgtzMU9d7QL/xh6GxA4fFcf1nwuffzx8ybye
tOpAVGmhgSt5eKxX7c94K2fFXFBJxLtXvbRxCmmCeAB9S8ygOfaqmmdDnkidSQPL
86S08Kb9ef4sPoeNmHcA6aC1bVvVWrOOLEpuw3xKOvrMiNHmGRuzrNT30sRraJOT
cROAQmYIzWe27wzKn7urBoSe1hFr/CGo40+Nq+WPgRkA2pOGvmDv2g1FcDMYoL96
ZyNtSF870ThsmwDh0aYsx5Insc1I0TXpk593KxEQUWONF3Fc/Fr+AhqaBywdgaSk
mHTfgyftqlABLsLKVy0skLHJpgi6Gw9NuzKAGfzIjD8rOjKgGQRqRcl4e10FTe/I
6M59Uh+1+GCFNxaYI294LT+WOHQNzz6XlDNvf0kzmgDz+wLK2M7Qb2aeGxIGsQ4/
Ss4UOvSEfMcJnLIIdO9OIcZp+7KwMnhXIMTnOP4L+Ry58TsH7GSdxvUB5nFzmn+h
bAMcW6Qdl2rO7tBdvOBlQhdkv4QX7Zsu0e7T7lq4cYNR4EifDkf+EjJtCHvNur3W
FhS/2vfTzaS+AVsytjI6leSQCwXAiLMy3U2Y//8bDzCoSRJFpmZ7O1+YGinxEyhV
1wqQ2BzAeD+eeMwuCHl0q/gXFvgsGMEywM0Uw/OR65bht6I7vbxA5nf0qmgR7qhI
bWWkPdMoubf2akmisb0IoPBMws/7MS5VmI8ikCdThd6fib31K0uJ6E/2SZSRpqvU
gbgx4fDvyZygZI8RGgz/EsYILCtnLYCH2RtjFfhdm9CCme84+xtd9KfQ2h/Wz0VR
HGJAOPZ+i+yVlcoDFpZd2YFC09XnTMDKue+pkthUpdmqBy3AZaRamKKcJHBkAxNJ
ad2j+RsWKxgaCw0rKRtx57QiYKbKsOAhVQXW+Y9g+v3cpyGAobMxqKYIhiJs7kqc
KqBlIUjJk+m6noOqHHZKZQ==
`protect end_protected