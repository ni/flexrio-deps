`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8496 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
/GMbQK29Y+AAYqzOrLs1aXtofNDQzja9NaCJV9U+TSYIyCYjubxSSFgTHi6BMvfk
vMX+zY/oum85alqOnLzQzl52M+zSKzVtDoT9vopDmBJoM0DMjz+jgXFnQ1lfSRR0
4OknDEslfcbR/TnlyO/GleP7OkCqRuxkUVALpqKLhJAzEu4kJIa3/WVbBaRxZaQE
90jNkVdcUcgXSgiiM2/OIQzIgdQAzj6tj3HoSq4Bhik1Fta+DQuT6rZvj3xKyIUw
0PKx+lfqbez4EFbK4qls9VWl1g5jBIG66bFh9ufG6H1sWWzBNaiFi8H8UPiDheN/
PSWF1iOfSRXRUMxeuzEGFz0pUwnvxaGDaOm1e23lTHWskZ4pTii4nPBWCGuEgq1I
UoYl3PX+L+/fG/6NawuYg57wW7NFYAtJ66nfxDVohsN+UAZv+cQMnaklalVGWXnj
HmiXEA3gs7kmK4vk8gh1htq5Jo5oeWVBTX72ErhgaFfKYS3J0CC6/DYhrj9XxD4o
i9rFfXoQCKdO21BuDV1Yqr1qeYCj0nUuUf36/H6TflGUPQb3CvmubOYMf63fXFQX
7khf4qxuq3+FkY5J6d2okv+0PVd1U4pMt65mo6btbJeVuZO2EkeR8GXI85h5oq23
vgNSicmJcj+5GQf2FXqyANc3yJoUYmq+LMe3kpsiIWpG/WkJdsmSE4+XFCpSJJfQ
OLRzGNA/Zx1ejYzhCLc+OQo1rzwzoGNzKS5seIw8FWUD52hT5dZ1wXiG+8+DTFLB
Tl3SMbBNhHfEHlvf9Y7Qn/kuJn3U+bqUYQMy4LN/ByCISJ5kF0+RhtTRAG6Vlcno
/UwTeBFVQ8ZrH/OQH2GvX6HPmfHMFrvuQ/zFIZG91f1FltgnB6JqRRDwe7+HMLcY
InWWaJKoTqyMNE42/M2OLSDYhp2a797yPzZSQLNbPaoZO5vi79X5Ysbb0UqeiLEO
BaiTjbzmHKG+6gyGqqIa4yZHnaleeWf7DoCe3ZD74W6THWZBG3cekAc/XoDozPiW
POCHLwF7ljgldBkPRONlJoLVPMeq0dWXklYaxRxrvBwOH7ECL4jEQyAYZWMmySo/
3dk9C53XjJHBn9UUXOeXa8xpMKDywpZY7MuwRILu4bwuc77jDkdUcWzFt7RqCDgB
bOrfyMYoL4PhvqbloN5+rVPAA/znQFBHiLQxjo3hibD2AJoPgIfN6k6r2bdXqnaf
wGb+pMwkShVisj8fzyGpjkfAceKiE8UzdD1BeJ/tr/1Kla5ExMSMyN3r/y/lggP7
NN2wrel7LqLj2dbTQcQpnlHU3M0iTaswS7ySw2D9By6IdxonPOtsXOFbkY1RfMdo
/xCOSfOPPFE/yc8y7kgBMM/L0/5cF4nlovQG1svalOkq19b4FJ+brPxadUKgbjWJ
zCS4w05vVfbIRJKByastCf6FIgMXti49pJxvMqerRsghFxocC/JKqV8dtWKvbcAI
qpGlsASZhikSja5MVMdMkORjUvKZzFKgCskZrbwPeOqH3KDcAuopHjjOn4lUBZ2Q
8djdRiaQAmI3nyX4o3EJcSKyK9ZEDPG5wOKSOYqOtkIFluwkFiq60h6CuRJdnj1l
e9OaTkZRyODwqt+Ob9V2K/ODfAMmn3SGEtjn8fa+esRk4PXXAqrzXaQOFIbwCbjj
fAtcZMV+cZZtDGU0Okz8PhMC+NJ+eqQgvkzF9JnI7AauLwINXF5PEy+mtNxgqjuh
F9BN1ATFh74TUo5IbzihQUXeYPhWRc4h+ec3BZAvcAaSlURxTmyDCVj/9lMxnIH8
tdDtgwtHqUM5rgw1kvt/vBz/wWMEzyQE8+E70uGBWnkx/TyFJrae9X5DaJSmZzIM
5kkkKPW+YZwBYqKec1rIJnMAayiCh7h9zFCYGeI0Krq0ICycSuHi8vQ80aUqA2WY
zWYpDiAzu9kULERUwk/uD+pxq1qbp7swyrdaw/YGu9BLhtNzqDuAghtJ973X4PC0
hWSNc09BN9mIMHhxO4Az1G9IJTZKeTVFSa0hra2KyHQX8rJoXJ/y4Cm3uymWIKeD
BMS/Weh3VKRE+pS0a4AaOayNWZXrkVPi2oVMO4uX29NUhnMnfJ57VSgn5dplyhA6
GU/pDRcAL1qnQFPDldoHAoLrhqaMWdAZDfocaEsPbeLhDQI0pvUrbTIVl9LH26P5
nJq93t4MGYZsmByGV7OA7fRnocsjQzMYIilVu912BkOf8LUxH8eS/07/8OJD0MYa
GJGcj09luqsIlGALK9sAJjKEZRVITLlLz1iI7d+qdiTzIhfp1T/5f9zoLu0ddp+C
ZF7XsgSWA3k+m5jBVCX1dcisNKfFtewVO2pJF9j/yCh7aiNrrzYqUqmpT9HKNauq
MOubieZdlwQ+eHgS8B0j4xu0KGkVcTcY7b5Ll3jnCK/r7nzc8a6awvc9d7TC4LZ0
peRV8vltf1A4hVjzLM2Hxf8Y2EEU+0k5adWWK0821wuK3n98YzpWZhHTD7T3jhTB
ZkuDUOKs0zkOCfmzBHgE8VzXaOiwIPialqAL2oND1YtPUQXSORDmWM4/pwUNyzr1
49sm2rZqZNQ07wTlduQZX7zs0hcvVTMI3OicEwzjs8VZw+/lcUzljhv0OodKA1MX
EDs56chhzD1XdhMtXgtjrRzjlrbC6VqzM+iBKVmIHYdECrG2JvuLOaIQHpzFe8fG
viMJkXK4qn8SnMkiOle3gGaQmoNrSb8afUf0C0AEHeVAY6dpFiy4qdEwZHIDUBhd
OVYBGANlrmVwFIPgjjK4DoKzt7jsHueeVO4odMxMADimaXpmVc8a4MzWwAwThTxb
srQWbW9tsU7CQ7Lc+inP5HMMd06hmcDw2w23RFu3TW/hdB93PWn+wHii6hx4YtwA
m7gryoSWTx1dwZdwwTGMOkmZt70iMQmdLb9p3LZqkhL/jbLXuczimhP3Nol97a8N
BJmXDRopIEqVWAD0cWMko4Ld857KspiTUkFxTR4Oi4TbXY5Pb1MmE7AeiMDIHQLY
51xYo2UtaM93pfzGSxE1tqq3Wg30KXBE19jIh8L1RCZuVugTKrLBLCqmwL3OO96x
c0wP0UIaGOabKHMnJlo7VHo969BLiOoptWAu6c+993D64UvWf6Co8tnIS+ycspl/
p+QMggHQapW7/LR2PnUMB4PmweVtY4rHXoOoEU0tpvFi4RzCtKl+1utUQppBSkbm
G1O7QO131jQeJLHD3ETs9ZtsC2mFvYvas3Uf9ziyU1fc27mx3vFlXcsM+0aBAs56
v5/tDLJUQwTusCnkhguT8rozxIf1u/kw9hz48PiOteFHX5gmCB7lrDADOKqs6r4x
0NBJiY/hUVOdHYoru3JVvvHOMqI7JS2vFawIW4/481whxJUSPH0CjZh03v144zTO
rLedmkuZITP7RK5pjwGon8PgScE64dgeaoOsxG/whxuK0VdgXOkj6ss0AAlpNjvC
XYOPPJOaZLcBYnqUA45uaudt7gavrwJa+/Mz1WyssORK3dwvguJnHvVUwhOm3xGe
GpZ/4ASAZ5H2x988Ne78YlUn7U+q/8Xzr3Q0/P/ycdFiuXE3Yhb/KgwZrnT8KUGS
z3FTC1WVOTa6pmjJAZ67d8p4ncxAu6Amj06Xv4Mx7av25JPMHfPOz7yK4Gs8AcOx
wsOY+3Me17dl6v7PHSkHTcxgBgo7zavc/Bt/b5EG6TLBLPO7wIIAZl10EAyy7S09
ihG1NbieHmPByHV0hVaeIPCpfHOocJpAKZGjS9m5dBk/4RIcSToluZeCrrphd17m
TsMd5cmfydkSnx9W5G2vVhChMPwY7GuPvxYrJLcJ8XauLKXb/hyu92eDT28tStDW
EutBrPZsu4bPCUfx7GNEbJuLpGAL6USUDq55HhYJ4EUiLUZmILwHztW9KRsetCPr
GeKKKH5PFgDgHplRPmjhYmK68bXGH/duKwD3Y0Z1e9dm6AaWN8qpUgDt8vHO0wUn
NfNBsipohSz4SogN/UesDQcvdUavSljNkHbYhzPLbjfUC1YIRGmqKFQuAJjKYFfl
Ci4s3qGjXuQ4rZf5SwjVbA36II+RPtGED9sA8bTN+3MhPx/J5Cr1a5qMdKGgUzdu
nrRM9kbFXYewgDJUOa0ypyscgWdv0l1TcZKRP2Ull0tKmkjoITLQP4vY1Tb+jrov
aYol6yNn1eMQ/S1cwMDaSkHRPkObj5sJi4bqTj0KFcS9XazMXl+0t2rQjP2egHoP
mrr64cg1Y2RS95NyR+yMB1zMRZY8G3ZlSBNz6A17uRAZ/ddyZutWgj5sV4T6aup+
BeObhPeX3kLMtUI4TiM7IfZEsVjNeaaamHlMbQat7g3AN0UIX929gcbvnRQLh48V
pYlR4nyKrS48lKgkfDisNpJzggUKI2ifBObbgLiTi4fdyCgxNFkuUvYcsEMif4hG
tM5swdfuG9/7fN24gu8aHEWeXBTCCSZTqiHWTrmyys8wzi/WqCEqKOyh2HWULwyh
hWt67Jm9OQMMC83oKZrKRImMmqgJurVHVAv7uqiNXruTzH1CjLj83nXR+in6KU3T
i+l+CMRqBSgHiw2FtavVgfyPtk565BpxJZMhV7lq9vox3g8LacJweaAOVtTDQ+vf
TwMk6Ht3OYD2k9gRKbiwDTGCGeYTF6mbsrd/IKBBmcQzX/43Xlq3a+jNxR0ssu71
kqQ5c34wy1oyB12BURt12heHsP7szCCdtDUCo4fg2vdbfoFO1NfHNml1sxge/D/A
Og6M5grxcrgNwyUIFZdBAJG6nTm7vk1xxuG+k16jRoR1vNY6iXORxZXjhI3WVzUn
f/8AGSld+N5T9aKIE/Vby9V71HVhO5c4bQDhYUXsJNhnm2EHtuWhJ44IRV4FRAGv
GwIcEPFBrszgz7IUuVjlYVv903mMCXjKyMu433he14cTAigzmaOKWI3rNDD9eJqz
Yzp/pdB/OxIm4uSludi66J5VbR6c1fdBYc9/Tgq02auays3WfJfNBfj3YD2IlHX6
fIVPvwllvj4EFwU6bz29YTnpPjphw+YrkKEr1HhEcwI6hpNG25w5QmHPdHwCTtgP
3VH08D9+PUqbbqrvGpF/ErdvsU8MNtmLVoveTaJmuMltBd/yRH+rKydOYMUyXPQS
4vJGG4pMfA+i1oPlhQSrzvCY1cJYwebs56dW9w1jZQddwZzgpHRPjch4nBFAUq5q
RFHcpVm2G2Hv+T7fa7EUGYTWaoecJ+eYBfJ/9xXXGvI6gVJUqub0qrSyCZA2VsbP
lWVwb9E+23HUY5PiWA+Cp4VCTYe2hFtgGsK9HYEs7raXd1OHVtu1AUJaykrHJUYO
ib2zx3eoUOfx3FCIZOj26vsQufpStG2gmeY33hcyUthtzbFqoSp0xEDH0N9jSwjW
VCBUW3nFzvfbUDrZniM1vxANbThoZeDlXiexVBuWS5UsdT5s99fesu9g2dr1jSkS
Av9suSYs1nPffOIIvsq+tPddWtYNyhubaPZFvy2IM7EeEk2CQ0JetX0cr/p6xzcA
5xJG8PDwfGq6GuY1dnp9pldbizgjB5O3+pSZwIqxGf7mW5ZrSmi58cJWf19ZRPq/
wpVmCGFbYOxohn7DFrI842baEcSHo8Cy6i3VIposzOAJ7TfjjnJQxY7QzKHENeRI
nWXRQ4A2mHhIaVgRvN5r5/CBUvo9Ex+xhmxfa/H1s5JxugB+pjenGvUg0phDTE93
T+wQshgy+uyqJ8EDQLP8AgU1ME7rvkEw8ijbCVTI8qUirHtJwHsyL5Q7cGHhL30C
EbM2fWQ1MD/1jusaIhN4eJN3vVhhB8OAJOigWfNIKV1vfYkWbRDE5pFnD924Q4dv
wC2+BmLyyKKdMG8owTwqRni5+hVAhIhpuv4N1Q5pLwtTQJ9VjTSz77KZ/jA0lttq
qAHQuBuWkGiSb+8wFKh5fIAIGuT45Hhbm5nxt0YmMLl9O57p3sH1+kbuVVimP+zH
v+WJqA9S4ofIJ+KaMxTvU8SVe8jAFuLG62Yo6A3OxsOYYQCAGn8Lp3/6FjNxm2VI
OfDN/W0MpLxTHEYxRMQY3GYwJtwcLx81KjSA2DbW8VFuW1KQLr61Rkzz3jiWWEbA
OCxBjZOOQM94cjoQ6i3jAr6gnkwQRJvbYrGZTgn4Ol+9XmkNVUNW8sk9kBNgnIVU
cUFV0/MiU2JKvJy1JEEcUloL1VD5k+NMRhm9c0Dc3TPURkMG2VbBgNF2o0w62nYx
J72mjh6wVzk6wD3ToI6n7yRltOr+XJCv0oXJCJyY7EQ5LsTkJsfd7d5MD+qJCviu
GSOBlnbe2rjxE+tZgXrxXA+5GVjjp9aI19yU+ZxwJL3YIhfT1WH/LV0hTjybx9ER
AnK9EYzM0XyaCsK+K6fX6WUw34/2n3A5mV+oPO1XM0/bEVptflpZ1FXx1BlGRCWT
bKETAelQij2uwJxntj8bNlUfOAtml2GD5+j6vQ4VSyCzr0ajMOex+ddCsfNLUdg7
sBHUYnCC4tg8nYOA+mD/tlSc1g89J1rOUI2oBB6qVJmvvy+oRVAtthxhhXhMDU4H
nensbCYzKfI7mNhxN5E9qhmlSuWTTD3BOa/ESy4V3aGQhiZgPU40WeSCzpE4yWy/
vp4z3W/pkjylidTERk5SlVSeqxJzNYuRzgUcwQ1i90oOGRtINdDNNYEOE0eFBt3X
skymgYBrsyXtgA6T5OdUB+ta3gl8gAIEnch9wR3sSgZYzy8W7YhvhPV3gV5GSajN
1fVFHdnBVixsHA6jNNkt4ozaOcMAqnaz8SYT0StI1WjqZGPTwCjAz4N0oo/CfiVP
d/1DDlJ5BVyx5KHwD2SunjSqN2H9pmyt7Iwvo6ZiOIuJk87nNWxFhYzGQnVgke2s
zLsWyQlpO9y19Gnhpk95omCrD61Cr15ujcgEhhbUMQ1w2TDaSgcmFmcl0KE4YGjH
BXFZZ1LqewV+B6RYfLGIV0FaIs5D/5aIVcZybDDJ48LaLf7qGUYwZzOdJinss5I5
8sgIeOEZoeAL8fm/Zk9A+np6GQIysDl5rztCKdCzZuNyq7j/vGXWl6ud3TVuCDPs
uJa+dkZ5gi8b/JVBI7PXHJN6bx6ku1x1pR8NXBxjGKXCaSK28iN7XV4xJmlX+vQt
YKvSJSO5pcNCMPDj9s9XYHDYkH9ImDn0m2gcUzz0u5WBJ6avCS+rolHi6uldfOwa
JmlmU2iHemhRs9g7Qsr5vpaTmnKfcLAqfNjismOyUrEGqfjnDvn2G3gkkwkXUCfC
HpdsHmbWyqq2o5dy4XuFYNud4Gq9e+M/2V8voLZkmsrgkxKO4bUFgETtG59jOQB1
I9nw9rPnSiZRyLITa8BIvHYz8h68K/WDvthZSEr+hPF6xO8O5PJzcmKKTQ1YKKAP
064CJSMz/9288ZLIqrgX705kedLMdDm620O+8QeweePkeB/FbQ4kDDOarYm/ScIq
3h4PHlwnFzJI15AkoAc8WP8Ba+dXp6yFT/YLCe1hdd/+2SfcdWuK8iKmAOBOE4K0
OU12lBw7YUdP1ahSBoVcT/l+FKTOaWnjwv3o5Y9jmx4VtuCjzFK2lOSUxDOY2+1Y
XkDREumwsGDMxa8ZOfQSGdLoX/mS3wSCEz+JNk9yxToaHcrda/X1LWRJ+bAQjf4t
Ucd18ByV+03az4wsKuzSQUZCzU/bmv4F8RzpUMqggS8KUn/J/rYZ/qQcvlOPP/lF
Pqg1pAVgn5UnSQIM5Dhb9G9UqdeMyiDwrkj8x9R3l+8AuEdn+4BhNhWnKor2znS1
7W4GLNUbHRkS//hQ0hsbiboKFlnxtQaGpchsEdpBpmZjQp1RPC/qEay9Az7tciJf
W6otIUDRuDDvQCvDP7ItLTZxgzrjGRO9M6TPojuoed28mF3yzfCW+1O2nsdHaXH2
7USOjPb3NXO3M1MCFGht5Dg227uqCts9uyNzPC5t0KPMghKPvUOgJCJL0lKh/rax
x+BC3VgCkpjmXVEdsOPltNjwCY1hUOlNZObX6IUMQAFIlgwwda3dgkUZqiMPjtfE
KRiLGBpGtVg2ELQSXGU4CaJMT/v8D9opob5MKTGZ0sz+GY7kJeXGUTRZz2VjlKM4
vkS1qflXffc04IjmZBYleHeOYu6mcgrO0e42h3mZAAQamVmkkcIvr41KgrtOs14b
qz8nA04G1ps0JXUeq+AbbF9G4gcBVhj31b48BRgTJL+5Ez0ysbfqgRioSp3r8ihL
t392FKetlNpCzrR2Luw1uAlK64gtadevzMWd7Yh24GUjsl6HzH6M8TZAmzVnOATd
oX0q+fA89Gg46LIfitf1cHqxG/i4ulOpkp093MIQUAVfI1tGeyOe7EdOcJyHvKPt
jWOKP5TezEZ/rxhlbrxL6P0Yi37rTfRGqgbWgs/pp2YDkmzQU9cEPgc2M7c6jruV
6Ky94PPn4m0FXf0kqHnTPQw+u66RvE23PhO3VZpXShg3APIYz6MZSFKmv2OzvONX
efXkLntR7NT4kJCx8rhTmkm+uPsJxPTn8VdTLRhxw2lYo/qa3+5oWB35dv/l0C7H
tSXvEjBWEf/Zfx5bKQ2RALX/V2nQiYn8jn9QXeWCb/cCaTwSOrWYno/q6uJr7i6C
qFo8zrafncq/pjFmuwjxcBnrvNc0EyhtYMkn8NlRsJTTydN400rC7+8bBEOYT70J
muUq6/5gajV2ciDeg18OdtTbQ3UPcfLIJn78kZXXF5F4/x2LiMCLCT3ln40spuzZ
gDz1++fHq2zHuMevzMLPcr+iQzd12mgaVNMLkpGBX4M1WPdQe4ZKViKETYwoVsCL
C9lxd3MAqycaTRI70/nZdqh1c4JmM1PB0FW2wE9s3ivuVhmbS1llIgD+Uuo2WVis
D4P9E4RZeOEubwaZdRJSJD3AqbE9T+y9PPnEb0wwWCyCVyYscCnLMccZHI82PVb3
Io8L73F58KKMvbkp7zBbHHK49rnonTANzgrPHaciyBXKQ3MsGJJitKapCj9xRcbH
TrMHaD7ZQ9hJGrq7eV5T3n5gh3YuWACf6Hf5bkK45nh0lY3zE0/Guq2r4lAdpIbq
Tvdo7xAjWpo27ueq3I3thwYzQKPWnSKZGzKoVH2aXcpoDaf6C+28+pggjvZYY9BQ
l1VrfeqWjW7JDN1ZiQIuXQzPdJQQZ7ZbBT0FQQ2UnxekMt1vUGEiYQX6WUZcZb5a
/wCoHL7wkW5S/fwKx1vZTPlzGmabWC9zr+XKu6LMloYebY6oZXjoJBWrtv8YLM/y
85B9d2fEyoRgOnGtcxQ/1D4z3nh4bqNHuLTA2I7EkaTvUl03F7qRx1QrPKPSUp/8
f1lVZxkSLMl1oEnwNdc+5bZo3SJ9ZGDrpk9rZdQ1+DqIgvYqohgWPmRYviKnbSXy
P8bso7chfUyp1LvPMZ30t0fwiAL2Jj+WI3Ut9NRQ+ZgMk6+jqZHZc2qZcsBDIIr0
JJxbvOiVO5hEk6574IkGS5mFyf59NPw6On8lisU0fb5C8FVyAMQPVWD+9H+H0aeB
68DVfNpa3cCO8VSdbW5ZrtWvqVU4gdM0FtQdVM6dDRiJBUVqke8EbtJQc3ySn9M/
RODBWwW1x9CyT046+Z4qBQRg6hEmDZfH/Il0rg0MS4bB13vzc4EKWFe8OixgvZRa
IITngZBtTC/8rX4zDayHpivZfFiATRc0PDXEfuPrmD8tQPXsUJBkb7gtVZIfaL1A
o2+cRWH4nyee4CZ2dYEbOGweZXogdMT+/gUkec3YeR/SdP8ORlZ4xQbYLvTHd1ry
Tl5edDGJpOLsgFlVDwcrSkm9hGw19w6LC3NhxFTaaIeojnFSMy2iPdNEbYwnfT5E
feJCAYKebp4VlyqcXml5oliv7D4zySRfy0HKyt3mpOr/WfG0Zkc01L/mQNXr4U0I
IY+buA2kYUgMAU3bSJOAL+VN1A5G44KjzTqKyPcMBGbTkbwg5bnEcZIX7tNwll8X
hrBNrOou98WQjFzpMAB0U2Z5xZaTZFDjrIFIE+v/ZXGtO6LUP98eEAN7sFq3c+D7
IJwc/lAG6GOlmIER2B0EkDY8T8d5UM7K5sVgFZfwclIj3Mu4bRZwbbhVHbxSmNiZ
6HfehQth84xzpclX2GnQYn6lDd/oGbRzL/KZvbrLvXknWRC7r8nmmk62Hkg2Fj6R
rM0m7evxQoYzBo3DF/DHzb6RBBwuUeqAyLQRwoE5x5uP3RkrpbL7oobdmgoaXG3g
qSHBEwWbIVVMAg+HD2Y+owwU4rvzJk9HAzQAP8W27Ke1QzFNZS9lFSU8c+xvABg+
24NvoJzaecSVNRUHYxeoFmHPwuml8B25gmSu56a7LSg7fo/fdzmgXUPx7RffX7tL
zFuHWWmmsd580CXTT9dL06g0CSHfQMlZWxv/w2XKrLvup1iHP/ZkYQtf4cf89naZ
XJHv3GRnDfNJoL2zs7bqbmB9KJpn+TiRHZatZt/HlVfMs+jLR9i9vaxlN5+uPAAH
Euiw8+BTEKFCvshD80xeCNi1igMsVNY+PdrDIe37lRp4X3lz2tb6ObYUgBACWPgL
M5RLaZlLxzhVOyuRg780BbO/CfvRRVybw6sqpoiQjsAs8CRCfMWREidz2XyTwFge
U4F8PVYOXIZHDpfy7d4Zf9ec2nfhU2As3BNat2DWx25WVco56fVPKhX8gtM5nA9L
A3pztB4iYsXjdJ+kDVwHFJuSZeG3ysqGqgMZfkEXbp9rnJHFzZQIKRROhsocGgSj
b7o+gQWDw1nqIa2FPB3F+x1hXmNYuu1HMKLn3KMfEO0B+ISpSfPMEixmx4mm3zml
jRKpl6+E2zSgApfeqhgmBAL3PYMyTwQ8nhGJFvq72iuSzdxDEgyz5ROicv7/vMnA
zGH4CsUR/W5frvc3lOi/1Bt6jEGFkdW20P30DFG8E5lUDrbFxIix1Oo7vCfYu60C
yKTxYO4WOtt98qOMv2pPzmuCVty2gOsrRBE0MhYZm4GUYh4hrr0E5uKqAyueVRDw
hftRCAJbsd1StR4aqBu/LM55twv9fFi+NgFqAglFgFDyFFKMbxPBKm/w9OEkcNaP
VnJ3oewQ21Gq1EoY+MhITMhgUjb+9wtVL7KtKn/EjbyqIw4la7sJIRksa0RFNc/K
QYPwA372zbTQrgx9WW5VoOd9jJsOpmPZjGw6ZXqTiUMWCctWiKSFb4J5PxkcqnTz
q0fga8sL5ZZOtGzQVRvr5i6YARxlVYjV5bOYPBJZKSOhzNoKc1jQh//JDqAkhPNn
`protect end_protected