`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6656 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
ki93Foj5FzFLQL1TyB6Fq1mfn0qvDBe8ivBeOj6+4hcHilDFjQn8DgKkxWZpvTSv
nXNjUuQ2c4yle7BAywXCU25qrOxJIhlLr5gvHTSMPUf850evv4I8QEDJpHjfdROp
RAjZ82Pr5aRcYrglGJ8frXMJNQ2JY6P60Q3i8pFA0h8vEEkhaGQaH2vNRwdp5LH/
Bdm9jOHJR2zYshN7RbJQYNvGvjPzXmIaGe6US4nVvD2twKTJcd4hRQUW0R7MevJR
Dv0RJEFoZZ2yFn6up67aG/dV12IriQIveZafav2z/+YgOnnzRIGGcWfsBGt3AFcK
w5V3kZzPWkGLB9hTef5OfFcA0xrcqiYpiGOsZfBPGRw6v1mDGdziZHalGjBLdubE
W10OTaM4Uowe6OvL+pCWjGUjsxGKnp/em6czyieYorKxzf8xl2fLJwnQIjcXv89D
ixBKJBppwneORHQMsoq7xvanPw9aco8MmPIi+YSEbamy240oqY4xJ6udlc339umP
ntv9klSsDlr887B12p8iu644HTYwbEOzG4fyi6B6rkJNEy99vR7owOdoE4irSWlL
O9LmmaW4bvBmTTFhkcVnj+i62XM7hlOxlKHvojWhXC6anDtFqc8tc12eSSCeBLgk
nLb6HAOdLyxRXFAN/2HagVHe8TMXttwzGL+L4FADUYNz3+ZFQqQkQ+WmSUGetDGP
s8TMaWj2DKHMnmbKYVqI17sjMLr7QmqzcTfEZLw01Q9Z20d7u0SB8Nl41Y1Qyx4a
7z9/hHz8sx5FQyolmt2Lp5Z5aKia8ZztMTh1ZGYHvBoPrb5M31/5QV606X3qbSbb
OqAu/1R9GHqRJ8g9tljIlHiSZFJjeOIajq99lPr9t5BpAL8+cYo268v5M3X4HZrC
DbGVfOeMJ+3WD76UI6l9w9FueWrITJ+lpr/saB+4nVLYS6AnLs2noCFj6T70Txwi
/ptpAiEr5J4ge3kzMIee1w+Sd9aQQ8fM28MttNrVhFo07ua6nHtM/gi6Y/Fh/hmg
ksgyJGdp1GNPnFWP5d5JJH6Ghng+mys1XGxadCLnocdNGhb9d3tKYi1wxMbfVQqX
6wA0e40sA7U5LYDqHxqIJo6NOOxrCDQ+ezMtmUS0SGClV9mngoaUjk/DehyZ0RNd
KteMfonw44syOgrjlOzaprvVr4yhwVuGkws5iy+mof9QZCFoYlLBMnPGgOqnFKNS
JmVV1QOny+UzM9ywfuJlrG0eIfUCak/Zfxy/TmnOrsN7px+oPMCXvjKg3ih0FzJB
iNZFC6i6+uOXtzaSGQ/gE9HUMG2g/0tcEaaE+WgrFJ7ZKejWgoWO4qRARrN4n7M4
Ap6q5lOLP1RA9qY46Ht88GC8AQO+UcOLDxpoO2gIGxLb+v9DPiqVTpc83z7nZeh8
Owqw/hVU/UsFNbSx+2RkqlSpJw7Eqp8a2uY7yQvxpqK/LKcPI/QXaLWmQDAEYtPs
mNMGvGib4TcQMc5j52RxmQSBi50Gex1iOK/t+mmIVqNndezENG3TYSeFc0O8U+aW
aDXd59OeY8fASw315gSq7pLNPQIOn+nMOpKHurbq70NENWU/yP9JffXK+q8Q83v3
kKG1671pl4tjoYtCJtBec+tQXgeFLTp/xQVhhGxtknjHSdqU0Anec4bvHDcj/FAF
Xys+lO5SxRy6f/nv+h13aaZrhhFQNfwFlH2AqF4nAGUR7SKCbz4vQg3GAVU5xxMd
ps69YJYUQpw1NumUChlomDejhmqI7p4gkSbeJaMUkX9y1pMYWVlnvjrIvv1GBKkh
KaId2kUQmdEWTm4RQa+JCitqsNv0t7QqZr4LBLoP1gGKlRHaDx20UI6niYro/fUL
v6+G3F/N1WA4cGjd7TthnhKkQ5rTT8TNsHMO9qnRIxS/06hVFQGnUwXRvErFrGix
eydwcuSRAbxlb+IoG6eNmLcORYZv6F2r36gGlhnrttuP0OY1D3f+ZQNo8eYRJDqc
gE3bYGagZNgpz99B1x/4XqT1d8IBWC4bkBS+m/6Hja6bNQvoyzoE1qfelTXkKRBe
74sWzpQksJ2gtiDT+JyaEJtqCyA96cU/9WrTMTWtplz4fZGzt5lET4h7RrbRZ9QO
7ngk0ytCmfTDZ4ZW3h+mNQhixljngIh1NHCzErf3IvhmjZMJVofSgkZbYgFoGHAg
h2mzX7nB3pa5+7ffW6Fz4yJpIsfxY7yZq12Dg9kJ/+cyURK5dUp1uaDpWj0myusv
kXE7Wi0Bfh2DxpGOFPCutBbeBDIupBRZoy8eIwTTvYAA8H8BUmADv8M8xw48y5sa
6zrgDU16zrxMcfuPhpVSP2th0eJvoaSd06WOoBSzAkWR7oaVvsT1diah/OaKnnc6
RR3w9L5A+mCyzNsoPUvtvl+DOL6wywnLySdFB5GrAVUlMsigCHAz7DpJTPLtjpbH
AVNt3lqQoxrpOUTfy+nUcYZ89S7Kr9d1ZwAzVDFIz6mIz8LpE2WIAXBBxwf7A98Y
j688PP8t/MajTDKUI/JR0BiUzrQlUGuVU5/QaeeghoKfUth5VXpplKcWVNgg0ngV
K0veaZp7HCXTiVHmvpooFYtHh3CfJ8Pr3k7euyxxlTXRDtjwS2GppJ6RrgXbZRky
lc+Nqr/APL/rAS6w16ujZj7OHFCK0C5EAs53RVz372rfBFiitW+0I+ggJRZy9+YG
UmoFXZFA7P1r70RFqX2zjXZsvTzfTZKusX+G9ARWs3l0K/UKqN5NgzH0fhWM/TXh
Mga1WhfAKMH2zU+IoOcvusJfPsBG9miIZxLMVRcY8qn7Mq6+XGtiUiFjAeDvm9IE
73w7B767gLKbkkFLohMFwjCfeFPmBnhCuUR4MKahnhSCKxr1DIR8JGxtLiqBa6qY
Kz2s3EWsD86n9dCNrJgmqqFC3Uc61+Fodd8/azdluPUbxuqVoTzqAtQGuMIp0wbV
wce9idlg27IWppH7V3oNUM9qYEGIAiJekiWuyc/8Yc9MkKBGmy1aJSrd0d9M7VCP
KnxTT91kmwFdvS7vPhAdNn350YRh/sSGagbvpQj/wBGa81//FRaYZJPJ7YrrMAu7
Z/AjBSnsFgUv0Q22ibK1dp+GahGz4NnsA+v2xxuJEWte19+kgFFyVN3WJO48za+I
hqZh8j5FJlq81HXtvhBRB4iInyEFVnJvcqyoA/qbSQRDoY9qYXDcaqPIm7lbJZIr
AU7JjbVgoG2vthMWDam5gWrtSjodmSzYMZdsifXMhxh/Exo2brpgUmr9rXEkToju
tKs8XP9BsfQMhDWtA4qI1t8zE5whOpynnF5FEl0aITAFU5YQCHL+1pB89xgc2gE/
1P0pRSlEIIjquheOqH5JsUhaghZTzbPwCtGHODft8KohEtrn2d/yKsdsjEUC5acN
NXIL5c9pqQ7Q5+FZPKG5uulUgeXyHynqVYZtMbqAMJ+G1IOlzWlFkP0Vpk3IIpUE
2FPJdws4bJB9ImKQ7pLBUlXl9Ehxo8FXts+pVLrTNUMaESnsawaVrRfqZsB0CtDW
Q+cIRWIoao25oJnMptlp8C6p810iwrxNw3XwotUcGLGkgDispwjQaZFOWfQ75HsD
KJzFSz6NuWIsBsxO7St75IK5ylZxY+MMB9AStUwP9yiIbFGZd0byiqG1gWJEwoxY
iQ72vmAd1kx7/oie945zQ8s4TRZS9xvEqVsV64CkT+eJmPgwD/qibSVH3kTREC7+
QlT9Oh39GKzX1op39Cg9+z8FldqeQxnMdPQzx7arYysLaQAcpePfz8vGjBVNy+tM
ucY2vxCbL1Qv7zZ8D6DYxxxc/PDMTN/BEZ5aynBcNuXq48cuoWmxVsUkB6uazxjc
SWLQcJCUcrogTk4CYstSn0Bby1NwiteBGukCnjJafppwD9X97VBhk+fBqiSH+hon
DYyBii9c/ditF2bnIv4tI7GgmJT/TtM9Wt4YGQ4fjt/rEg1AKpkCsdC+oxNo5X42
KD+ZLBaHTe70aaLXNM/vXNRfnkdH9yPysbEiiWQWICSo6RJWzGm/wo/wm85ezUS3
SrOE2T5zoP52GtXX4458JRwH2UvCEOOg8grnCzRQTjZAqOe8HtX7ao5+Xa55ColT
jUWlRHKwqHdPn4M8guFKtgRWpV56YDtG1dk4Gv4k5hyrgDmoM4voltZ3IdyQZQfl
C6p2uKrwJAYdtKfVh9eiWdBQ6Rxhk3At+avTEY/buCGIkv9Fam5E5XtkR1MKC4tR
Ron9AKaGENb0YY4IPYW7jeLOUGs+izp2rlOQzgqMU2EwcPz8nlAdMBL1MnPaqFCA
hLYm32GIA2/ztPVQmWbZSTt0KOQfidYRgTD0hllt90Vpp6P7zmEoK4+ebL5VtifM
Db6rhKdSeiD9HhHjlneJpl3Xd30/5OmXAwZwlIrbUcXwXFbFp7ZFATDDZQmvhhHc
gxJDAVOh0rIYT76BalZpak67upxZ/2vEOIGQIBZC8Am4wys79W69AJKbN+Yiptmk
95NVdBuRIkZ0vFKYU1QnOrXq4lNGU+3/tFgkEXHJTBDgfHctvw218uZK8T5w8bma
FuVDmB83h31tvWmUiPQ5YItZUnAgbh4D8eKwMLnDiBrI4nP5/FxrRkIvZs68N4bz
ggNvqeqlnUhjdKvwYdNL6TPDTR40SMiHfCn3J+rlmFszXedOGIvQbOZX/4/xJNiy
kVoaQ55O0GDsoe+RccVUfC2IQJn1+vOmAmOX+RuZxYWIrT+u3ZuS+lYq2lRZurgQ
xf6TKtEHdwyJlUM2PLHG8yczL0/dLdUKwgSsmONRT4/ERWO7YAhaDsfLMVeZpDru
V8l5GiwrldJs/A7pRdhmioqtZ+lnR2KnjdGRwsQJ/ctOjinLjQAMXL29sNOg1ROT
rGz4AAlr0J1Sdt1Ysrz4ximJpEruzJmJdSL5X0WmzQS6VKJtx/wh5rR/7RYBeYiU
HHxIZRhnt3+m8eM6pH0/0g/MAVYG4WGMqULYJFOuHq5xm++8C3JWA8hjcd9C5LYn
MRuW4EJoVU8uRjXdY00ZyN2PaiLCSw4LLz7gJDWFYqRtKkrLPxy2oVQ4Ggm9z2VH
HQ4Vfxg/ofLWQj5XfdIr5He+8Wv3ukMcVfdgV8whvT2j836N491arqj2WJagUCG8
0tXtCWub0uRWe7vnd7370vgO/+lvsHewgNaKF7p74I4/vZCayrEsvYxxf+x0P92D
lHN/MMNh3srzFABIoDCfZ++i7syWKaDHj3NpSluCqkasR2c0VcGHg/P6IYtejvWK
bwUAVAEIgmWyeUZc4whHSjCz54K7WQxb/sw2pi0niTY3gfuq2j7sSMGUH0ct4mq6
B8w8bOkM1sr3rYbQPk6blsLl/eWHrcLNmFWkdJbU7NywDfVBna7ImsxpcGJjPVSv
S/OzctBVZKvqIOLv28H++Mo7yW0k5G+Ca0q+S+DHv7cQ+jAx7Y4Yf2I1GHeAFnF0
LNqWGIjHPl/+hS2kRKD/bXVwtKcEfmEsvXlfQ1qaQEGzZmwI0SnOlpWD2T9URjKT
GS2UacpjAaNVN5Q9keDReCHuHVe6ZU3i79CYRaO+aPG8AcckGFPRyra9moZqLU/G
6AbWCtUDMJjqYO6h4ra2R3aighLoUmcew94ucc3gNPSu9p3h+MCwlmWv0E97BHjL
XlwCO0KnATDXgR1kUb3WMVFmmFsD3SedOOKtQz4xmnBHmj2D+NHPD6o0O3XIvqXZ
WD3CdPOMuVY0+kjkUd7R6ZeSFwk9+OFdsF+f8vtQeTlYmBfvd81eTrstJTZl/QYR
ZA7Ge60N+WQJwBHBFEGOCtvhAaGCAf/+1OeGa0F/UTfJEowP9bfCODn6FT2GPKmZ
9f3OnKrx5mVyfHnhVGqW2SxRLkIs088VSideNnyarTUz5L+B4XhSrrSg5pnavDK7
P6bNvJrXXDY8ZimMNbKPQLN+iJEOl+5YdqE7bkzbb92tI48ZzM9ukqUg+5g8Y4lj
gQn1JJUTk2+KmhT8OBdjzWFURmhvtokCwXk7IoJPCPsgRPhlT+/WmRtn0JiYofE0
DCSz7TfG4yKAimF5JLLeGktCBq0XulLf+pKmpIiEOzW2MwoIiUau0ji5Gaou5ySP
7EWw55Z+3vvUogkANxqTpx1QoscKI1V4QW73E+0fDKhC7JLIG6cZudxY80o+MeX7
QxAvFqqO9DeGNTOzU6yHrbq7X0yqtMn9C7hkw9hZBXv9QwJZ8X4QjPL6y8rpEcvZ
KqCvpfOPkhnwUqKzTFf+Joa95O1hiSOyzm5EPlOSYP5GjjYOZXyoULYaK5FEFz6r
M9xsaj2IGa+YwT3Gv7yIusPOH1k5jTlwZ9Emo58Sayu6lDJ+E49/0GL3DgDmpDJx
63n5W1J+m4xFrCB4K05DAd1+ok7hcoObfLvVk1NKadWJ8gg8coh8toysUaerjAqP
jwdQhtpOJqere0lAS5Q3yc0wB90r5d9tQvuRjq7P8Xop4Dzw7bPr51zkdwpIBBKO
1CrMO/l/fy5cJAaid+FInkA8XOPggB5iKxXgRPAjBBTxRlbcx6MIjyzhJYMGPOoK
mJnUW981zt11YRg1darbkFJNy9hORsMur8vKkx3VyFOK6fTdcA66upssRA4+bFid
N6fACjFKOq5NMhay2lx1FzOj/NWdLBPJs+Sz8u+l1Bvo70YmRXAf36yhsd9Og472
sxYX4/zAxrYguyei71fmbUVcZPQq28J51Bokv45SeAxh/+CHHj7tSz/AOAWlHfGI
SKJCdamAV5b8d2hVYAbGEMKrRnbFmw2LR8ArLW7wFTjgTQW4+vclvqW/94aizx1k
PVFkioczJRfLGAHu+DnJSxHHlNDFkrIucoy/KDGL4Szwcd7Y8KC1WlOSRXYVBIxK
kB0b68W/CwrFN3IQ1u11GxurhTZHZFYaVW7qoFc3OmuIvJkJ0XLay6ULXunsJNrX
erSTp8uN22TSp6QsUPsREJpccyTDJ8SGuxJXG6fm2g61mJ+AJT8FRcJjm0QnaMLA
IYFdLBg0Q52ZwNwXos/XnV7QGPVbsUSU59/006ObeTPcli3g03gyGu/02861Yc4d
gwoy/2rlunKxXLVz1ejmEUwTqpsPua1GM8RhwFEDeVIlNoU+Qy0J6FgryYhuTQXz
d8hRRCkMqVYSXEZTfUabLlvMNmnntqBdS+2NvO3MhOhrXFmKryHi01KJh+V5myn7
L9hwQAKW0LKZsmO1gk2zVbU0haxb0u4LpLaHcjUGjRlUWEudlKjJyK6jnZBXehki
wYzlfd7umOm170Mf1DhqWPaP8kHIIDQUGq/Gi2oig+UusyR4aC7Aw6oFsWD++T/J
4mCKjihyKTkepMijGfKemZr66MhpToRhOEWY0nRi1BwjUhEemG/1ITlMkOih54zl
tLDKv/6wQkKGLHn+gI48TbPbTDHtThVTkYB/tHoiEMuTzKvN832wRm/e03NChXnO
HdbfCrZO6JXL6Ygti0UknqweIuaVF1lNONm2nNZoJBIjbZpm4BIwXIoYh/WtCket
aGcHOjVTSNRiTMHuyatm02k4YusVVu9XqVHHKvcBZNRv5tfosGmK0GoWSDarI3QU
NEHM5ZwZiq0Crbpt+3yXpjOl+xXLL8voe0sg5EPSVGAgnf9nSSCKN8pYRLOGsbGZ
GzaBw/K1ZQ4Gz1ZyxXkv/bjUtf5a68PlmWxBUrhRyS97Filw0MBSXTTmB9bWNPpi
Bd2ESgSnkzg0kKp7SwDTVRKFJqlUki0eJEPQTKUSPuPv4IjRLKwVTsj1pdN+Wv+y
8J07UUntPLhu3hB7Av1WhD/Ga1seUsSoz0DeHPrjMScDBY2hn09maeG0wLgxQ/Ah
WIoYLqq1TuKDPSxczninih5rxN4A+H2aVNfbWWVOGz72qYWQ2wEN50t9HIyOwpyJ
zC6VEAOxs3MDYDgXAqcV9cGFv//3IGTqtJl9WY3vZyVol/wRgb75Bm7NbniGjZvo
iB2jXaF2ALi4+TUDqwhZmk963S8ElAB+S3gyUQBf8zgPPpeVZmOpMmb9y1KyeKIh
VG16xUrfWQUFFimPqk5LSEc1qx/LTU4Gic+nHB6GC5Ok+aJqW+baQPDMYeg/MGQ4
VDdfd8RhsQ3dKMSB1fo2gxMLOx97uXrMhFhvuh0Bem90YsFlW3OXquLmp9rbRJeD
P5YnjcHtCo2SkW3xhBv7gNqpzBiUcEUliVk4WUe5yuk1sbmjkXUJJB75JDti9O/c
ltSJTCfArnyK6pERmfQZDB91h8EZiz7hwdqj6sDCjtCCagkt3suFv6UqnyDCw5X2
9PIKf1j3z/jBOQO4Xdfd6MeH88LAKAdtw5+6a/CHghLZhbq5CasEkHYf8zmrRhjs
HcTizvehJMtwAzhX6q+ttnAcEXGJgZHGLaCiBN2HpIAWxXMRXf6121KGHdJmJ87F
GcH4apdL3ll7YEAp34RoTn5wvI96FaqtH5V9GdLHkuncWrdz8bUeAsasDZ0bskBI
sypuGAHnMOWBTX3FvEMMf7IfRuXjle0zcwHHeV5yrcpfUcBBWdrx83u8EgWn9Njs
1GKgBXPTmxdgdkIszTMT+aHR86C6fxBKmWroJtfZ+jf6ScNYkHQJx+VPbrXEtkP2
70qBniWzdXzMlODwQjlxkIN3WjBMvDfdMhqxE2onAGs8muNGyPINMuhwgqZSQlKO
p7nCtVI5+acfGRwm7omuyOA1CJSfyB9J+pVVOG2SQ707Dtu0kO8s5a2nwv5DuPnL
F81BS3GwGH1LLBtZoWeQs+WThwxayJ+XIETMG4fyRKs=
`protect end_protected