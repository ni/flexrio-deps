`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4128 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
CRVGrXj3LNIgA7Z8dvGgacR37c75aQt9423YJL1xAplupVIlSo+VLjTm3puwEqWC
MmkyEdK3y3RoU3ns17dnUSXzlFbq6HAN6JQEssqdV2p9uP0QxaCqD6XNDhalTOmO
HPPHMKrwxrqYJ14GNeAYXkRrHly2Onzeq4FkVwLDw5nGbrSNaaaPkfyvKfT+iCB6
lclm6J1ykJS0lgZ92qe0ZTG40tgazon9Pm586jJVus91/oUX0SlR+lrwQ0eYsTJn
ZouYG5Yxjaihk7Ruls5jIoIPtV/uo0FccskcZkJy+w3ERzjqH4JzF9qACktT9OKy
9bmDKUEj4Rz1xMBW0naOuESxvuc4hf00Wq2PF/Cgl9uYss1KmAJshZ8+wJ4MP6dk
s7D0TwehFHVEApgzvJ9HKihAO1piCAm1leMfmG3LHgVGFb05oZ28M6Lt4nu4T7bi
G4bYqVTAnztGerHxlqecYd5xNOWgkNi8M6h1Bc+DlqX30omy+MLcLb2XB7SOnDDy
4AgIC4EimpTy9IByd0eDift6y4kZUCpOcF3e7Hxpv5g8iGxAZ/BZF4Wp5gerMph1
3l80+Q5XTGVv6Im8rUErAb/n1LSho7cMP3xw0WSRrvxdTYEPhNbZOWWPq7rXFUgd
6W0YkDF12IqZur4Hup4wwo0jqCUEcgStYAPdm9xb+hm/kWP++JUmSeeGDVTEgWwf
SYYD47shjdONfbpImMQ+1KcHL2dREshj9E7jU+OtuF2F/MA12T+ofyAMjHmZq/Yz
tk1cQm9Jtl+t39btkzagf3VAtMEUutelvBkXr5DaCl1fJWl01yZmMntaDRf5F+Tj
NDRxP+8LolzfiiNoLbAxbkD8tknAL1ktAjIIEKijxpNKYw8IVqP0JiIcDl04J03C
hbWA7aGldX4TbBu8g85iiq5+GmEe4UwYydaXpO1YpNFIaSTvGcsviG84Pi1rzNaF
jG/5u4w2YAhAb4FEqxJhYhAnpEv57ryUi29jLLFMPbiUc9x3oHewdFjVkxBt43sz
TmMEmYIdsMjj0mgxxRZGLwloYbB3SwYiHHrwnRVRTZn18+qRJNlROx73CxxbgPYb
gJ4XSpAhcO9kSxgjNBw8QGD8L7aJrG8aviVP/FOJqeFzcjymsd1Ir8o1QxERQUG3
B2RNk9zOzC+gRjqUO8QNDR1di7WeM7jsRq+U2oPmzjPfbGb0emNZYGORfFlI7LuA
Z5MsnX/4GNe7zJFA20DHO/ctiBjoYb8ydp60aadFCU9Wx5LxWFbKZxNiOvDvqFCy
rYQHEVPCVV4zRcLEpNKGJS1h5dGc2GobUHfbefH9xq4P4DbiF6pfip6fMPHqvmlj
FI/QDeL/XT1ZAY2QQYnLe0mk2y82obyENaKPa8WW0osqFYO85RUZbTj1o/R/UOeX
kGkn67VsUZ4BGH29xarq5uns5021K7VPTpe2w6oD5vED6ODVARd1ct/MeIlzMaGb
umL4NlDqmsdR0LkuWOCGDEJ+/uRVSp34HeoFHG//y3jh6+Jk5CRS7MZYQelBlTVz
stbh7GJe0rxQsycn8iGlC3rjD2gTZNISl2h6MV4BXwYKEHxGy5wL5f0v3rj5f6LB
AlofRByVBMRlgdK6J4wjnpu4OLETSRGcZKNF8kcoOluJMmPkR1tmp+t5X1KaNCH7
FzZ2XHZBNvfDOudfcISgGTdx0YGNICpmlxJ29mC5xCL3oPYQYDFy5cbJZ8MMDLAY
tYZiSvRLPlRq3T+2TwybX+cJrqrKAtKByMEGnfvf2xW1TiuSaEQItnKO/+Lxf+m2
baptIQX6JXIS9lptfDbrbsuN7r509YQSpXtegePz+kOEOvOQz72bfr4PHs/p6Hjm
ohNix4ytT0i3SW1OtrwcvT7S9wcWrnt4ExsS+hXYbQNvjblfHa/VomEQOn3wXFEV
yRvx8ooB8u+tRLY8kWNmigXeUFlgPGK8YfraI+R9tMpZUbnQ2zq42TQY0pQ77/31
YOb1w9a4ra5f8OwN4RNtTBDuITUS8DkGV8i0uwJj/04NA/YHQvwF97BexE4owS+y
yE9AVqzOa10fv0k7IQlt8MGvOIfMyqjWGk9KC8fMh4vvw3gkMO66BxoAalbEISEz
QpZvitcH/cDMzrxRuFvzks0o0v6SIFrBL4C6II3XMUm9j2WV1Vdt8GCkqzTq4fM7
f3Tb3E6gGZ0a7LL2i6MoL6o9C4SzZtXfiGLXL49LsL9jFdhrYQSJIpnYwvPAr8u8
MqWd8hPEhmAxiyeItq+tU6SIoqLjD0vCjfVzSYESVIs9YudS5CMGa5ZIhyPQXjky
v8fvlw5D532GbkL+4U2jYSn6jQ1UA2h5zv8VfYuKc67/5o3toJjjKyuSCZCdNeCs
za3OPnUpOXx+GJ6VfSTxrZS1nn63RMMEtdGo8ztSBkjEBlY8ICVfUJF5jkGcQPIm
1x8IjWLU+ITSvlnTUlFC3kOsDE7Vx3wjya4HCQ2jFs/+tZwA5cZ4y+tykCmGB/6O
2WY5DgYx6v1zDMtQ05aqfd6FRFPGkX3h7AgO6dOyCF7ckGohsA7+pA5Tf+v6rMrQ
Ix3naszSNyc/sJ58vydsTuMse+G0OwcuiIEsLspVRrfGa+GwNI9BKF1+JSWAXUj/
wOI3TE5ku6RIua//0j38LOy2D8fIfNsXgFCSMRKRNh/aPbRyzdN0g0eifkMzv7SV
KXf3eh8yF/NJP77vdkZj9Znjdn6BudO0NaNy8j7KbE90eWJroVYjw37ytaDGtw00
j5281ZqbMv/s8+ffYYuWZWLpq5+wdTFB9iGH150nwr5z6bFTWU+gZUTXHBh2MfKZ
ulpjGFpRTdIQ+vf8xHJ49+aSVtwP1wj5NaVMvQ+bhf8Rscek973XkRg4NbNZ8FX2
Zv1Jsas7pDj/MU45YbA/tyJ6XmdT8ztkUUUqrnAulxUKO59AT+zHPImW6xiyj7rQ
r/PP4Slaj4f2nQNLCdYEbc5pb61rSf0Gu0Si2hI4Ikum6yltekiJzR2AtoxxPj91
yTiDFda6fpKcG+d37aOs5T7kLcUGzzVCwHvnp3Ic+92YhC9paryjE8zcSm7IpiGh
TXVTa9R9/DUQGTSn9l/JQuWtctnDjjft1G0e0YFCvs5++zDhyaEY9OqTXT39u2gO
/Cu8zdboGvhb3EdVbHdhFiHCf9eDb2dNWPdjXB12o/TSmG5haOHFUbxAMLOVCKhs
NS36JGT3iRcO3vA8PevPTXdHTgRj9r0o+WVE7mXRQalnTPARXnbG/+Md53rUk5xW
oPtxlfiicvw2BTkldLH4ssVZE6/hEaZ9Kj61KNxCl7Oiy/Av0xbwi9+/TWo81OR5
IONZSdcFuDvvRe+CjocJ2jjtwEJcXvtpiANvTlpyNuAag2Zlo45PsVL1z6zRm08D
n5YPoeyHnTmvbwBPlKicOwzydZhTB8edIjElax4uPzWSUMdbmSh9y6NoTqc5EEil
1u5h1Y7ACFA4DXpiXVCMJbSP4OTugFVuveinnWz5KBrjViwI9+VeAalWKyHctgqk
I8nHBcftkpUsMRIMQB3cO9s3NJIWEsgoukI8j4VK8veXnMK9nnWN2PwhCpdDcAah
ee6vAS14fQNoDo5e1rATmJX5bcnBRI3Tk5LZJG18PFDG47hi7LUdhSXz2OhjUU4+
kW+H+TYYSP4R7VBxhGBxXSI7U4iHSVGR01lRlwnbaAUdd+TEMEeWLRWrYitKg7o6
tNTEREs7wnKO5o+tGlB19rzEvNYXsvtzA/eksk76VH7q5oxaD54rj+/ZlEnHM+bv
V6T14luyQDcPQeRt9uLfiPCbad+zP3oLDK48AaZXakPFHjOC+p2/T+X6yedtyJpM
3H5UlNjuHK7CQiVu/1rCXdaNjv2bh0i9QEpg0V7dCoCBlZiNB+R39MW+Sm7xpvWz
Kfgp5l/BGWFyryyvzi3HIWjyAHCCEa3EXGnOwMWNJznVLiKFQv4CkS6vh3xl/JvX
XmGe4Svowi9/inK4YJhyGCxpNGKraHyf3WWw3VMXrhGu+8usLSsjRHhk3XI/yDBV
5wjvfoUZ2HWkWSqQ0uNoRq5ntaqdGq0yMYrKIUSEXZ6m8/syGfuAuBHpILPYjCE5
UYnAQEjwZmTUZNNuqc6TBofuLSY/Q4qSmwBa0ODYC6lf7nzeu1evN1k4JGlNYvG1
z9wAvHDaD7mHO/ivUQeNWU2orqi2ksARrkppLnvDxSqkJJNrxd9fjXDt09/4dLZS
YcPFBO5byVk6CNvDkD71gfITt3Vnv1O/ZzqCkpGYEMtJ3rHQJ6lUA3mys9Uvmj90
m3Mu3GlNGfuvbjuzb210r+9JwjdfPI2WTV4lUcnDzIDVrLk01gg6dgeL4POPho8x
P+85zb1k06owUUoiOIY1rmMfmIOn620Hq9QLkSJgkDi1kxqNsISa4Mi8i56TmBQg
W9RjEwwHO9ZmpHJpT2VTkw36V3qZhrhBb/rJqvx+OgMwvkXfRfWpOIxv438MiuCJ
JVee5AD3JqSUeyklCLjM2TfjjKro5h4lsggmijq47B8tZI0m1ManmelLBlZnW5o4
Ny1aqqqLEHkti0AiaMIdaAUXfV1d+qCvtn3X8ii9GdJj/TFDhvnLfRPMPR98QDDM
gkaf5PNFhyJaqnT59gyj3NDGa8501vuUrRbdwmJ/T1Yqa5d+1eDeG97ReszozGq/
4tDpMjcEjToGKAJwtVlBv/aciZ1WAWOzOpiGmFhVV2k1Q1mRpT3eY6CBoA3jmtCj
uW3m0s2+oR9GXUqgBAq0UsVOe+mUI0vgU3lC9U3v8uETnEK9qWFV36uM7MXVEt7p
SWTfCV2zW32cV/pArKqb2K0culCfGAmji8xuRbFPhGSzjMR7rxuSld26r9uBv4KQ
yKt4iUoGYFYeyHltE43ZYUmrJCxL+HUXpxP8C8YBTQij/buzQv5tVRoRcsKLc5tg
Yv1AlDxkgbQZ7Gj4+hfjYVZUwcaeNanEphAF7H68BMLm5aZzMw4eCcbmYORzJuG0
VpNW/KaMvzwaG/xN4B4h4SrL6uJH5F+vvRpm5CewBzZNv1lIdIGWIr+gzZteioXm
4M+l06HsZLfORiTkoobCsBWuuxC7fBoSap77V+E+MG2zhuei7qd7yQplMWEhwa9C
VpD7p81uox68AyCgHwi7WredJI6SgxGP5CeyyiNqzRMT396gOASbEvS8+40kxiDW
ijdDc3T3gINiiU29w+hDTwGTxMSoaorpQSnOiaAwnoy074pi0xDOvEz97+xPfkBQ
0TbBWg+3sq956NTggXCZTDTj0T4A73Kx2NMLxfIbmHhIDXb7azqeOkVarxukuMae
jEaupDeA8h5DN0PJLlg+z8OWnYeiehsdc+cjRn/JtxsMImQXYikVjexAEAg/jfj8
`protect end_protected