`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24224 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
Ju3IpcJpVj/VshHyynUPTOEpOOFM9TWog5695c/TI/jU8JfEYrX6IaW7OJ0I86Vx
SbCEYJqlmAg1xEEbm6ckdTuJ1Gk5ALe9u2OC/ADJK7sykP/ZGOPL9zd3FWv9rnBK
lPwAGmSdmCPVTaNJl1GyGHmPVCqw6OtfzLpZZQ6hXycDLvBGjBz2/X8J+pm5ybTK
mnYFO3YxLdPH1eWxvNUJ3KJ7kf1SH11JokLBKfqciXbZkQi/+QSQE1Hd8Q53eFRe
zRLG7ogJSIBLZxZcfFVVK+PTDuETyjG6FUzYNGIlUYOxSfzjQR4gEABlgpLBqrf9
YLPJmjaARDXto5qYS/TB0HNGV80a9sCsv9733zJHnSsnH9NAxLZPYmq3CRjNOsoY
WI/EWpY0dQGYNfzuwQdX7yB+OK58EEni6UbeO/Al+wvGn35Tc0/UIT4cPZ+UD0uu
Sc4+Sa8fiHhM+ZqVDrc/HcSSl/AFHIDwCdV1Z600u+usrEOp1PVG29HOeTubJSBd
aj/ANq2tlJe1LqUC+TIy5K1tJ972oPV6Jdgo9Qdt2qV0DCL4OfCgd2IKMijZ11mC
Y+l6NiGgO6TU0rmR4y1PmpNh8c0RYDU5JT4uRnTuf44qL/yKc/sHxYuGUfZrtpU/
51AuzHDKJi2UVwfxrMS7h1zp0H8fBwb9i97TgIb9o9Qw+TVP1tgLg9Z1hJ578kZn
gBikhV9HUXXAFrVCokGOsrAKI++8Y6WXQdB5xHH1Pb9RDnoKOMWjTLnQ7rgtKCDq
rwZVMkPdfAUhWvB93FvYSA0qGenEDWwGqwvB5j6e4jmXj+rRTTFYK3O4+cz7AnqE
x7ixz/dnafAmDDNGm+ljOwktB2ONbau+KcVwD2ckUQvjE2z1KyLNDVlwqo4a+0Nv
Xoq1pe4kCeR3VO2XXMrWiTiGhtRhdiYjLQCLkGtEkRmtGYKyg8O/azPKUV/E60on
hWPvs5oVao6dzEje8DmKPhvzwnViXTAcE/0w/19xHGKVBHig815tL4HPdNa8+hT+
x9+MTM7IqW7KDwyWCp5x4NlYgLlg+c7HGQPjyWahF6IdyTTp3Ib7ziDPSinuQJ7B
AdkqBUXddr4k+TISOaSFVVgrKpxG1BOT6x2YtDWBpGGkMbQck39SJPWQgUbJfrYs
Ry22LcPc2eoEISZBo/38s8p/pTuy+Oe2VsABUKrX0arhRuMUo7RzxRkXTkDcQMWK
XSGDDzjVHfX43U0aGp5CXd3v0xj8ZAR+66T9X1FDtBsa8mSaHsGfV8fNC0BP57Jn
wuwwlbhiBTUQXeDL+H9FoH2MqQm9cRrIBKw3XYZ6zIAluFshQ0de02sLM20Ux0Ym
yaVuwvLJczS8dnV5nReEN96RcXvPtDbpJroetnmwyQHZ9YZgfZJwFT1vuNMKut0e
VKg0h0qoLz0Kum+ULIq/1u8XdrgoKQaQ+/5k1UUTh+ed+VXlXQpZeTa07aa3pxs9
IHZuT7KXOjoR3GoYqUAhEd/OAKh8adxfkkhvfl75SFgjSQRtzENvNd6X9xMPToIl
tMDv+LnsLFl9QiScud5nMlOP8fxSaKeepRecagZYyoHi9HaXsaQ91QXz883nxO3p
Evg3GE48Qjv1vtvweAxWAMb+DmjReCoalYxXQCOF6L2LO3VBflnZ+IyMcy12554v
uzvhQk1k+sLTqjHC6L5Dik4fQ5wUV3sue2hYRiWN/WHpm2M4I4ldIfmGSCB++B4x
n/LnsBDHHq00cl6LFoeAOOA+zXdfVfjjmlghDd+OSfQB7mEQLfdUX8knGW4HvJVj
wnz8nbGnxyJqo9hI+cn5lVo+Vgi5f0c5J+37mGVrW57WCFqJY7k73Z7FODSEJlxj
yVOyaSiluhu1FFDaGP390K0nBjssQspwsgjlqh+SQqlwQoHviL+HStmwnMJAGbwF
hIvQyvFYMH7h731Wi5nmcvqC5AD7DHUCEub8Faf5yvzJqrp+/uWprSMbPHqNVkOQ
WZveW1zzTsNN/M3dlfGAV/9yeLxAdLFl6ah3NYpWBYlYz+tFPv0WN8wa76HbkN7X
rU7zLPp+U7JJqe50heuqZKmh9INR+Ry7pr8aY7EXwWE+bOlYrV7oZrnduQzbuQYT
RMugE8LsZLg0TEiTSqm3H0mGaDGXCP3Gkj4/8L9Io8UQOpG62GURe66tgxnyIuz4
+4iXSEiSrDRqdo6oZhCrfXDAklxWlMq64gx9O8nLMiylkIpGPzA9iF2BqmN8uT6M
TQe7iFQgUXHN440riw+9L3K44XUkYXNJddprc/ZW+C/6caI7YFvS6Wuyai83d3bK
DirKlbXqfudOk/+ACHLEBkvI5+usjQmEnPsUcQgy9PAYvFPZJYuy5MaEOXGKPzP7
Ipi0x8xnu8wH0KQdeuc7MZj8y1efWgaRgjOzniCk9NKEEqSdcrgBHZAlmZErc6tN
K1WrIPol8g752EsRzUegNyKlmNj64xiHb4mqzG9VhA3E1mF+xMi7axqm/ML9X1nz
zWlsQz1hqcEA3dUPOl0Zkc7PVA1EyJ1oy7M0Mk51lwX65Fsfu3W4bQpQ48TwjaA5
mrPeBycBHZdWbLyRo9IOwTR9R17aOSCOMM0u6AQDTjAd9/YujOTQS2hlb8rhbNFC
qcaGUCLSKSIHTL99OWSl14gHaRPmhTC/qi5g/wV3hInF0dXLnKz/WPOsoOFRCJyN
70F5UUIg3kaSiNHrlkIXIbHB6JeUw5GQ7VtoTR7oLT75vvbGtO8cOIbDkO5i01UW
HlaZPWaSF5KEfvsddbvgFKRw8EHhrnSyfnYT5SVXAZhup94obIOgY38S+Z1k/7xE
2VzjDWAA/02wF8BlnZcnfaQqXOWzKoEIwHEpc96h0n7RENyJn3sHgiXhXzEk2uEu
vXkUyT/DsYHoJsnvrWxGzp7/4UY1z8xz696wrQ57e68/oaWIldbTZte23wkBfHL4
m7PPoCE7Hurryk1EuhNWKUBL5DdRD0iBq4MLLnwGaZ9B4GnD11txbpfsBP8K15kN
XcTbeuQAJgTXCp2AxL045bKjo89E2dXlD+odWjmHqyZYQYpIAKNv28hOF6K9VHxA
x2+9JLxOKps8bY4vEQMZRmd7aOoxS3OmEbIHnH5BaUtpgm+D+KiZ2uOiO4x0Z+eD
pphRTVTqR4g2ZcDFM6Bi6mWvCME/qteFyk8CSj3GED2jVx5wdVMQCIsWsARfcYTl
uTOGKRL7AIn+KZtwM69A0wMr+XqLj25CvpXWjy3hXwH2CC0au/wmEcd0DkpD8Bco
amtMYp0PnKJSuFWC+3A7plFYHulKoA9NqkeU2umOJ3nGz3DfbjZ+0IZf0Fez3X0C
F6nh9vd9tPxRTEMWTf3ycKsoQELIEBlhMlBvJ8f3gus2iohHAHrQK9+zI3LsKCmx
CgknV5tG3XMdZIYVvw45ZXQrVWNarsdqvo9bS2EAnUMKkc30KcwsDlQFRwgx8lYc
9QDYS59qnF74hQeqtbCyxUR3mSg+H/iVy1FRAuqA+tqIowhYqvRHCJyUfHJQjT4B
ux1LKmEvRc4wjTUtw8oobFPJH7vtgcDOsPXxs9K+SYtqdzeOkPg6eqe7LxOcX/kH
EZ5D2DGnAG4nfJe1y+U17jwOhicqCWIt8e6Cf0B77kCbZRKYzlJ+OT6ZlEs3Zi/o
uKdzua1IOJ3exUh/Ws++yhX3sfzgqeTyYL1NCl7mydfC9c4OxxCRIRoXFr8hP1mr
GOtCPfUQTMUk58M+s/qB9ka7unwzMNSVA2LBsOd4mLLbCd7zLWMdIpB3mj5GTOxJ
tiUfxXPonXhiJsIjBw7UrpoxnZdgLriOSx/M2WfgZH8XjkYKv4Nn3yeqtdn+aUnw
Cg4dNcXxKdeNXjaRKx/AaYgDTEofhyJwOlQjEYLAEsCWGHc+MyLqd3X2pZI5Yeu/
BpuEX143++8Jbq4/kQjA3g8mXEK1wQCLuRKMaS55i3AXMqSntG2n+8g+MdD7lIEe
qm/TcgrOERCTeHNw9DLz8fXMr0tDirHGMpbCoH+u5DqTAd0WvUYb8oY9gDdtfwaK
S9PfefHdEFvs8auFJvTa8OFi/anAuvrOrvdR97zRC5EN2pITLRonWobmqndmXoOo
dQ2rgKMuu7QM9d+cm0ZEZHvIHtfwfwj5I5YhYdMgxUdVmgSut3AOcHLIihjK5Qs+
rYQeRMjU9WXodHLmQ1rB2khtGb3fw4M7/97pda1m7EGIQJzyBCAVGuFMf6TYfoLW
TEz4uSekK0VuoqiCGbOYfOvO4RQF0Pmy0S6vhfFfAzsbLrCPGEZ5YK0yJo/IjUdN
EPiqTk4rhaWDhSE8Azy3u8gcuTo8g8EssUrhXkCROhhDVTHLpHqritYKidBer7L1
5yo9qA43BZi6DbtDxXQhEFrjPt5nCzhwjJeZMenU9v4icvGcYJSf6AJ3sn6W0l3U
tFQrt3fIpbQmlPAQl8s0AoI2nWAshTmW3wRyiGOS3Hnwt1XGvU2g9yEwgme7SSiS
A+wBaelWq6PtO3ZrPSqvTH99KUVYfJHLnx9fDh4tAA2ZcVy5RDw8mkGHLuOsRJXJ
w8jiAGukfwSoEbNUCTTOqCtutu6FPC1pJoV+0tQi/43SYB3J3COncjoNpUXOjdoh
wuFDtY8YmcO7OK7Fg7QMZEtDvybtm7WymZXw0aOZmeOU/yZH3kRqJsro3i0w+4of
JQmkpfw77QBx7ieYJVSUo6NL/Kzy7NLFX2ZHlEdibhiy3VpeMWrXmehFUxmFH5B2
9xNe2JxHLpHErxjNW1I8DK+4FJuzEoDp87wPR7q3VgFu48feVeFTbfvFC9a7IEjk
7ISaDgTXhAULw2+fRmHDN9/oE3FEb25g/xyPLg6vZTA77leH8g8t/+RqyDDzH6oU
EaJO8TvfcCdnX41wQV4p6L1NV6fopa9hod8G387MbxNBnpM6oMNDPalW6gI2Yudq
dmHROTQ29sO/52ZL8aEd2EB+8gHIWwyELtrVagZ3Vzh0DKx1w5JHSbbg48/KL0VI
vShqpNLD4NSJvLFtkB5ZHiHnUkKsgR2Iucb9r09ncm45jlRAV95w7pydPjjpAdyT
NXasa7ITX111gQVRHrGJVMo9g1/w1DcGgCdpVaPuT8Bz0FYz3D/jDzINWCWFKUBw
q7AckT7L0VXsVirzpm20kbTBxmijLkQWbMFZ5Op3e0ce6nDDYvqWp/KzifoEZAli
qnJOZY1IVy0NdACje/o7fSSfy4sZN7KucGIpB6Dk0UVGin9/1/YhXgJwXQXv7hr6
4R16dDKIJofRCwZI2KdNPdDdAZMRdprchiHwgab77/mo1PNpBL1qyhXo1OCfDZuR
kOu/RQl7COcZP6kmS5ATvDGeO/LgleemyWOcEkzU6bRtxcTldRYMVNGMbkWSScPD
+jaMu/dphi6EYZUHVBPveiFQWRgSvMXPEGKF1jrKOEz0+AmL1TDtluWonVrvRxDb
AJzL7Hg865LI9b/4QXk7b8hGGAR8L6KXq2POHJhUXqB1KosD3ZhWa/pu9GDlFeq5
ciewKP/GWg4IzA4C/UoWm5vRhCTgPyojhcfBOA8xXspY83TZAn/kJi5+w71I0Tx1
O1qfNgptKyXsPuH9x3IsFb6s6Lhx+ghVcnOSh9lPKG446GzydM5k6Ttu/Y0YgkPw
y/fdxLhstty5pY4Bteez3TWXIK5h8+lO7IRsCWse2UPfCKIu+fHbO8+M1lCXFfDk
XtbXpUxn1nvxs/TzqWuHmRv+A1VXFRfPtEC17LN1dZN0ShpWJ5rCPck6JHvcwOSo
cOTsoIGaBSSklwhIX7qJiPriBVo4JyIMSe8AO6z8SwnLOtitmySOrZmLm971JvH9
DeTBoU84iSj1QrEy1DfxOO7lHP8lwsh0tF3dN8gEBRJwNI7/lpbK8GkIaEwIErBh
0D5okisA0m97a4I2HXO/oTRCphpKAXhpqtPcgO3rCMU5DfZ6ox0dE3n0BiG4lzKf
Bi/w4V89g6GrVoDbszf6aapAen3R5SNJNlptBwiAMtlHUSPgZ72vu0XxwL/wSCrY
8yEGCaJd7Y9P7VwDpBP3pgNwACqi25M1oOLPXs/cRbxi5ZL6d0/2B6WjAoMc7D0k
Gs5bn3wJqSoKEbWCmSpUrCtMgQPbhcsDnf/kxJQobKZPb0Iwk/MwaZCo5rGs/GQy
68O5/T1BkZC7Q9vogD6nJQzLOqXkDq3s1JUFIwYOhYLgeoDBqaTHLUbPqTs2AKYy
47AbYtWQg8PvP7unfKarrnGQh+eWzCw50vLS1pu3P39tAEtcPueQsjAJwqMFjEEC
eav81gjRs/rD0Oa6pKymq5u7KWi5rz07V0koBruzk1YBUK8KVGh/RNiyny1x7eC3
/Tr5O5Zdl/Vd012jMKyuSlhVNqwUvS7EOAPqrWiqDM74dAZ9Anh7wE5oiEhqQXgY
E+Phi7SE8F8wxoKK1ykKN40ire6bDrR8eFWaDprbOIY7PbS+KTotjpiyitXUGufI
9TxNVmAv+ISVdgzCs2jXXL4pECuf4eoAzAxD2lgjLplA6YDUk4rMzbKTcZ8EWMty
koH+StqP0QBslvWb0KjfCEPIXrTbynft0WLQ8FjYHqbuV/YMYFZj10dph/TUhQ4p
gZXz944Ishgg8zeUzrQn7cyFjWSLNvum1P6x0l/PASFDdm8CBrAYdKFYSAzXxYoR
2YcmoLjbpir1t6+Q4mCLXuPtcr7RZE/Ga97J8OBxWcjYSdD3C8yUE5GGBZN8PVCP
n0tJRgIDwN2M3GQrfVxrN7vsq75TR/z9HJ1QAltmo6KE52BXreEqLaOCXPKN8UzL
9MuEqhzlB002r138gz0l820elW6MFLjx7uOzcnNyvOQnsA3ckQBVaKTjwFMsWfvq
wTVIlXGs/W60FqKGAP/1wWofxWUCem5IucZduZzTfc5PIZdsb2IZw86ySHVFRHNz
sRrh+COjqlJLNg7uTvtfJONPWvHS1EXjHkWsyHOwEHnfxMZZJV2sBf9PVYBfPemq
wEQbiclQMn1fUU92VN8OTbtHZnVjH4rcX6KwMoXwg70es3Oxzal1hwFyuovY5uDG
qGGwN8jDHknTEFWD25lwPpkkDDUXGGCmS9gqJ4/PPS2JB18dlCZ28ikuuxNOVj7s
asbk3SxSSNB6+Ex5M2aMqnldmx3s/aoh1NHvzOXC548EW2a/FA9n9fjh9CCp4rAR
WGRAQyNxcpzYg4lR9KyGp7d1aarTZXvMIcPtZEkqs/wihFoz6vyiHXP0OGJk3geY
IGVrPlVXr5on7lZ79Fz3wTTJw7P34T1aCwWm3dufNWtbkNRZyIQZkpqFOydt2U4O
53MQ/dr+a7Q3h9D+qWBuwIow/RsJHUGOc0buSrEWkAzexLnKb3xrd0iHykHKj5Fk
N0Mf2J4WKSU8dZm9dus/hQVX9bYNEe2mhgCUSiUZUqsjkDX+fWUM2RL7GtJlIy6Z
LMrxXwgN6r2J92yP0MVMP1PlqUZjN6zH/QzmVjzLY918RWRHTfOkak4Kf/kgsMdY
Bv6ziY/CDjmZ4n9ey3x6Kxjo3E2CdJnb8pBt/8D+6V0ECw/oWXJLxlyNyk12Lt26
0K/w8lkyIqQ0/02YGgQz8WZsxJ7CYRkBkAgzcapLfVQfn+jgxS4CqbBjADxYrAvr
CuM2rRJh2ysZiubknIsKyoksHSI/5sZ8dDOPeHLy/i7MFDAH34z+6ERrN/3otUKJ
RO9UzQ/KnQKbgJlK4LoSTZuz5x2O55aI1AGj+q9Uf/dQjzAZRhy2mqCIDQBK8Cdr
0kwtK2Jcv+eA3lMOzrWWGIKQhQcTaRQB0C1YZy9mBuyiuNrWpaImKMJgWPgprd73
G3PrHy4DB4SGOoH83WFdTp346tlL24tPYwFxTkMPJ55psGeo9UsFCyn25aCYg17d
REDwJj+hmK8rabLMn9q3vwjnnMT0PnCyaoztg/XaQJh8cDCh/jDzKYIER6yrBwCK
RvHb4GD0SM7TxVyRf9tP9bwe0rsidK97EN0U68HTqP5Di7lDwX5iAjIlDk70cO3w
6onNfmk8Ly3DrIKGTO6wQwb2zLXNjF8SUF4osng8W2Go9yrF4Ph664UCzHIPxKTy
djwOZp/ZhJtPRJsrpxbuZYlqtC+sEchsj3H+lQRLH0aDr8KvDjKd0G3MI41wX77W
cJhnV4CSJOpYaUfHorln46LdzlqBZiT1IMCFTN8rORlv6QUD/bqri1zqxdt3qxQo
9fMqwytSZFbTWR0xjrVAE/cxKaDLGL8xREde5CVPmXV4RVpj7QmSAtMs87y63j3u
FwfgWPsVRsjZKi3X/mnKjtUrQrtHeXoC53tcSMyCJMxZeSvgkuLRGx+iEKWUmbyy
ZwjGSr0dLt+FHmSkqyIUb2xIXko8wmaGmHYKJhk7jfvNMqsLCXmqEnIFTwmyd+sh
MmFZTuZExzGMeixp80PZsGJWm2gO8tgPH4Is8cnqo3wq2ZkoBJ9c0n+gRpvwe8sV
rncXWx6l6t3VAhwK6baC4YJxcEJjdzdKs5yAjPumi0pxJVy4KSLpKqexSYP7DQQ1
StNKqLHCAoZePsKJJnfSkUkn11LX4k1Bkzk/joAebhB3ZHHmRT8L2f84CV+INnRI
F4ToT8RwsKVZZhOPqeLcGcKW6a1PlbqqjjGtC86bUPV3y+XzooC1/jU7+GH5nneV
35Uly5pG8MguLaKLYkFGzPh8gyzA2wa4g/DzyaP+b+opUQqbRUR/6zVclLbnaGfE
652J04/LSWFHK/XvWKC7mUZFck9cBSDdV/YVY6hK747ZmOHBzPafQ7mTNNVnc3Y8
Yo81cYlPNx2G1BYkoH2u7eQRxtHAlHGI3/jqDS5op6d+nRWMZ7txM8Yd0uVhLJxk
8R8gdP49wmUfIP9KPAkcFJlfWcIC5kMO6S23vurPQ2UoT/8PObhPa8Rf/9YvVHwW
JLqCUkHtXFy8W/rx/LWKsTQEHiv62adYKUsMHSBI1n6L4ALbvAzYyqT04KRk1CJH
oFkAzo4Jfl2itpARvxOk233BDBBgKq2MwWBZMrIaXl2E6tCE6hGpuBFskQ9wLN69
+DVmhYCJKY20TzehceQYPyamY0BgQyugkyMpSsMnR+fnt5caaVgvBRj4pnVmwEar
blp+7SVqn2x1lc2PGyeAoZ/uxval0GJJT7yydd6Sz2XMhOS2eEIrj3tV9eUMOuas
/k9eiQB7vU8GsuY03lAnphMwzlGfYh1mEWRzErh3EPwqCK+zWKWWt/jZhD+Bi3Hw
U4fyvY8jJ5XQoF61y3xCULC8tEU+2/cdB5zjj5Eg7Ugkv//Vf77CPO6FPylRlnPC
72WHdcA4rBNigvX/a4pNYiUp5gd/YKoQ6kKvuDwy6ER+Pp7GTIVtVz+KI35yIDdr
TxKgXm7UYQbcNSYFh4u2YdOKzTqmjIDCa0fAhzMReH3aR6iqu+n323dGhvJmOHtn
7DJrK4Ly2WZxDfaDnGs7wQswtJRqWqfIwrGwbFwfplkN8WdluI0ZiNsvt5d6aUX8
n79fAnD5Ni38vuS4OnaNJZtOvmNrD6hd0rCDovJrXM3qmaY+TdqTx4KAQ2gHdwc2
ce9xoqss2twx5tE4qGTd0OYeL3Z9SzsnTJ8iY80EUxJTaL5CaqUgQa7ByWmLhRRp
Y9fldiFnrQkc3l1Ec71ZaCoMgmfPmGVcAiz07kJNTZMqHLLjwQUO3q4hM07L3+oa
zHz0R+XNlVz9Ys8j3GN/yJB19EkdkpEPX/C+okqVZ+4YaQoIpHZFwFTyE+1/UkpN
fLC2Nep6OgAimiQyl4+WIwE79bovFY4SRZm1dgFRv/g8jBNx18EkjQh6JGlfWtmQ
fvV2NSm80Z31OYlxEVi18eveFxZurE54YCdYgIGey2rXyPuQBbOGjPU2XhNfZF2D
prJukZXUSo0Y+mIfQoRW+uN5+L0DqCLiOstvOH7wEs340Nlq93PrIevnpJjMAHZZ
e90F70tEAX9nr8eKC+wLoCxngEtlR6UlBhVwT4gDKh24z/Ykyt4aQ9rBi6qViqi6
TDT6IabKwFwLP4K+CqpGiZOc5UQ4H2ox+Hm0+xBioiix4zc1ECVnDL0eF+8PxGYN
6C7PG5Q/gFvP7/OC+QCz4zK1F8LKIplN1FJoNeA1qsghIBPRezNn1syshhW5Jyf9
ksw/NiXSYXlw8Xw9qND1LX0WSYCENoBUDCfywajDdZhN9BcHVnCuLOwJUJ4f9Inc
CM0SERD4BDr567DDURKWzVPkHogLfoBnYu8Ddbn++7jZlhbQr2JGidbA2PbZ90kI
BwRF4Y7DQ99F5M2hymzfN4hMfqyKRtQlaikGG+57X6Jqy/t0znLbLI1OqnpV2N7o
bpeZ8soH+9oZ6dWO8cLLvIgcSDmLz4ngwH4s6pZtkdbMLu36D1d/djro2mew0qP5
J2+zeOpALyvonqJwipsBjHJ5tUmdFzLnIayJIxlQg0NqTA7rJdQC+TOldj/8mPCy
1hygvXQ11OWvSP1iSDkuKyCa7Zs8QWD272Qbl+LAxiBLk01I4IX0BVin/XT9S2TD
fSlUbdHjm/S7V42pyrNhZz4bvnvlU/bN6tx1qt0e16uzyTr9j4CELOHaXALQVSpd
pcb2Qwptloc05Srbmx/2lvu+EetLNi1+m4482Uee/YRC61GgpUgHvnjMrptnCaSA
ZqddadcuIwBnNa0DB+RjdLWmE8kImRGEs4UNEtuTYrnMF+GK+dJt55DghZNmDHmL
jpzR8bm1X9CPvj68rk5hdKRsJjlNRHV8phD0ai+ItD1HdBPBPfoi7a5d85sA5bT7
uETQssjUe/621EuUnIsBR9P35/O0odKk6vlWsXNmj3UbrL1om3bp819XW86/NVs8
8449qH/5ZPtaMedO6BPu7tSExwvrIWeMMo5B32Ze0MG4aBVmICNeAO58Elt6dbkd
RObRB8uzyGNgIWlUGYGMEmHJxKvYq4u2pxf/bXblIzUb9qqB1iqBWLpg10s/iPSE
bKJEquMlKtfi93s1UTipnMZnpxd2z704IUFk/srX2fcP7f0diE5yS4x+Wp0zwYZo
GYUpSz1qBIiyhLeLI3uXwsl7MN0H5L32qWXEyqWBTzoOgsuxq4aYtUHjLw+qFxI/
WhQekdjlxwXbOt3a3yGkPV3pSkc1cx56BEzklJqOcs7NaHKW4rA7PLV+ZiB9LiUB
hrlPUnXlr4kwbKQaU8TPnYWYkTFVtDBp1JTaOnf1Q0teAddGqVypcRz512rLGaMR
XoDxzDu4HdzGg7DhvPeA+cqRk8hTKOXzKWa8JsXC7LPrqIumhOD+jlv9XhQ35SE5
k2PItgvlJKvOEI7Dy9nzWBRGftphHp3tsB/nXEXaKEMCsZI4ZuoaSXOR72GQj53b
bZGVjFa1ic8yHYvFNnRShSIObarUxRHMlkPjliYRZZ4hV+BQq0LzASkeutoHx5cT
J5AOiLfwssUaciEqVRToKuXCHQalcTqUoefzMOnMz8L0mXxA4pR+2vNyGRfl9XYr
D1V03DitPCPT9KFcP0k0xEOjDCkIXyC95RJ3KMFuMv/ZU+MTL7Q3YDhpggkFaGYb
85LlSJ8KGK4kdyrY/NRKNSMlQ4a+glopkDC1Rrp/hDmngMIgyAdakgV9UoEsf8BX
rpwp27nQnIPuvgWPYq1gue2Joe6GAo92341k4nT671VUVAkULJAFlgOflJ+0ywta
zBZ9flFILAZFJ3n2n46bFloXeU8js/N2GafhZoUTOmO9tBmTfzLmLLEzU8JEN/X8
8Z4x5b9srKvFXJKEiRrJFUQXKxxVbo1yp8SLlLz91C3PpV2q1rNVdrAqrfMqNSEr
rRfjcomwBDwfPprA7+AOP3swUn+ATn2U+NmEaxZU9UC0wI3WUNsjaLgwleAHCvRG
avSDO/9GFyC+miT0unlnUPzLZjVzm/YC4dZG7W3LvJbB6tR5b/ZgxwE57l1yjoTG
cLrU+VhG0C3IMPkuU1g+8Brqi06aZPixEHSrmREFffnvE4rS2O37FNNqoyXemGxD
HPdPnlkcHvUWV6SIvPk9Rz9VdylXftBqr6FcfiuEE5lGbfUUdJa5RBRiENPn9mOV
h/d+W+cwPWyYhDK5SAvRu3618q5Cfq4+Y9VEvsiabfespLGEUBGyKDRISCDqv6uO
WGDiSd+KbJx/eydmtcjTTcy63FNVpBG0wxDmP+koXT6vsQqMoAIq/6LDMX3tuy37
d+JsNqh0qTxgQ97xGuI1u/2hPxdEllGVPSkeEHvajsr2j+nQvl/Zh0l8zjxxmxjL
8j0r7XbsqZ8HtDSnCvoIOSl29cfF9ij7WP3i7678ttT5lr8iJtvWS2CrmE22vVBW
pvMl+RbjNBY3rqvfboHuLm3y+H1cWQrJu0EiMEPV7Vk6LxKQMtE3o7tXHVcToTTl
vLYohBrEutcAmwV9cL8+tJn831c1KnJzvUTzncB+8XH1z0lNgWFu8uJLmhpTgNus
SpwPEhdoxJ3hJjYD5M/oLLPhNy0uj+sgoztXvqNZ9NxX+U0v+fcCziHp4VLt+I8o
y2ljIn+DFl+j+SB4QKukcquqMoxyeKRvLHspLP68ArKoRlHHvTDcgM+EfEkl8j5f
7Oyrj0diegNmY32scbEeWu4nWKc4e+a53flPw0i6S+1TQ7QElBUgzzbsxOPUbdI8
1uUZS5TfEyJc3gLgn/Rx+AhEdeyc3DfMSpgR/vG5sOeEVU09Su0bTu0OZZMfRMb5
7w5d2AkOBbuzqaHFzkyE2U2f4l1I3fu1LSWrSVS9b/WQ99eBOuJn+chCHVBF0aKx
sWWKxxzD8EQ63JzOMfrRMA13vE/bFLqjKeIPluLSSq0pYNXsWE5ZbGQqmo18O/oq
CFaOxLjtt/RJG4TbZOLrXdjUPPRHGYp+Fw27v+DfGXmu8ZB1P2nk14zg+3f+HiuE
rKmf0LkNUPiR+DsFSRlZI514EeaeV79j2g0wPCprR6X1DxqXOThEVxEbb7BolNDO
H1fvYeNNstJAqG4mdEUUjya+Eqc5o2AWIFEd0s5xjYmxZofXUHZVSZZj54k0sQn1
oJxvMAahMpPs6MfRMKQoavKNU5DbKxc/EJblP1uBQRddlq6kgB+GL/SKxPXNGC09
O4ppWGadcNQK2DdZ/W2EfKNEiwgGm/WujRStlDQ5dzAMZyb8p5cGeh7X7kKg+w0c
n89bmk340uA0EGzj40VFfqu0i/PWLSEtizOjIndBt8zcpRH0V4koBWMYqF8mNPRV
E9kpJKzFcWEhLnItd0zr2U91GIRXAngsHuXFxbBDD8Q9UvpO5l34J+mDGLBurTfT
6Zn8Eq0juq1XfsIUfvMAg8qe1uR57qbqXZlTX4238I+I/EDuedjbvvhytWV1+cER
j2iAu/+ybfwTRHqyowARAd1XSGden2uZoXcitJnQL/ibg9GYiwsvmYQzHGAzPJjm
A+YNPnnF5MdIKnUyTqm/POJ/prQZZYyMW9zIIYqeG04cDuQDJMLaua6WDj0fqtQP
GjIg7dEVIbjqiRmeqr80Wn5mHI9jqHx4WBa81viuqfzh8gwgnOhrcEPjHxO0umMj
B+JY3eNZjjfa2wDk1PBhwwbdaqw7uNlj6+0XdHoYzIiHhaJ3j1LjsfX9d0QYqT25
IXVwWCSu4e+osI2ydjjwpsJEqeBsU6jijcl70UPKkPcbBrW6uT3/loz/w3fl03n5
BKc/+nPfz8YGew5pWyAKJSDwq8mIfz5ta5bdc68a7EhybXn1hZNLIrNzg01RrO5e
tf4sTU86Ezq1MWDhRvr7cfUssoUKukpCoOZ6qXgGxdQbc7lMXST3I2+wgW/m389Y
0+gVHj1bW4ghHUJtVlNE91Tg1965Q1Sa8zvVY7WxvDov/vwlvUbAKFU9DTWARowv
1yz68ydQce2CQ+AkygM0OxpIdhrE4qxUeEJAOs/T7zg4bYouF6qX6/HdXqVbh5HP
a3ye+EgXZihPgsOJpU7o62yYj1bYDuKWcnNLZ2iEeeuqenloVhEmNwwWGXZzoWMN
18oPCmiHvx571c36WgJ9atsPEbLjXrTk/4mQYWEgy321/5ZE6im3Tx6z8K6S//Js
S0OPzRlZdPCL58OnujjGDB49+8JDDB0BOxZSFZCAM9YKGRJxOxP3+AHQ31agn+ru
mZkJF/1MwFd6/lWieKKBOVET6ZGlkhnNx5yKotriS1R6n5pWv5nE0T1nkYC+RgVE
/Y1SjNbYj+jZuIm9zUSSUBNoHrE6cwbHZMvtHUlQDaZOoxhzeFKcsEwn8jFmB20f
BotlAaTAQFBTRvdXIxdYuMHclu9ghpdIeOi1VD203dokJnZ7Mb//k9ohSkRAAKXh
w3THQb//f3KcvRRffG2RYHvhwd9KUOK7dIG89A0J5W2Xnwzu42cDsOoLjNMARmQZ
cZNE/IxQivKJeKfH1rCnJp/6QMUVNYNPk1S8Ed1//JsuOjP21tBnhJPj2M3kGNvU
qx1wh8w4+n80w5Q8CqBmwOJOvGiVmNX+dsOmps6dU+3uwBF2S1DYDZ+UIfQ3uPj8
iVAJ5EesLWclJ+wSbozUP8ElfLViUlAEDZ09FUoYmDz+FdKGCEpQXTrAZDFtA6eu
eOseLRg4c9Ifugf8d8RSE1WRL6MRcqnl0y67zbf70SF8pxBWfkAW3iUJgqIsEECl
veYHebpOr6c3FbKWcyQDNDxTiJ/jBbA6O0t4vccGBR3UcD7wUsqZExlTA5V5aNvN
o9VYDfZXdujc5HlGQO4req/GHlSoK4VxJTwik6tJ8EmQNSKfefajhkmSae9IymWK
19/PXpaWAYAUVzDVCWYitczl3MkQIUzP7mXSSLrH5tmyzsTxMpouK7st9thGj4M6
QITwdBRPKODq85yd/trG2M0MPdjyP060MnHj08WieQRFbvSAifBI7GKQZ+UGPE5t
fhWX8UB/pfvGG7J8u9g7nXvja60WPgEId1YZNKo2wN/1wWKySiB5wbCIUPfy7KPC
nvK+Bf8nedmnGBFGROSi8r3KPH0CCEetrHDqYP1R2p5KE2E+GnTx3UnV6+8ABN5r
RJmTV+PFsDNECACngUFYlCO4LUP6uGMkm0InWkQgOMOms6OaFLU9TXcUkkysJ+nR
l5axVhCmf741pGMyDtvlJG7wGW8y8cXNV26imCP7CUtkPtyn6GmS49v8YE+IlYZX
yauWrfUG7RaJo5UALKHcaOX0tbA3gw2jJcON/CRAgvN+mZCzphjlUuimlNS5XKTa
Q49D9c7wsCgNnSZSYeoTfZ8b0/SG+gtDK7u2Nzcsh92ju5Oc/mBcT16L0BvZCcOG
7PwqEt5ct9F9bHoIgIWNfdOAOg9oNWrId4z9DK+s+BdyydcjVkQdu+iIR+NDlbIr
lZkxguUEUxWCUXRlBLFvs70BwEt9b4nSwahZIGHKbFPUv62Id8RZ/wiiHU0JGRtS
A3fbhLHKYdRefos22rJZRGAFMEIXxTgSAEXb0NzroeU7m1k72coHUkCEMxH94Zrb
JjhTTy3Tjutu8A7K1nSAYK0ms3qXgesS624MWD4IgZQCPEVPgPxPFNhDmCwg1Te0
emx6kDZn3Nd/uokC8rm3gDciLD6FN2DurWVWFt8KpMf0mgj6v5T1mUgstLxAmFRf
+2IX4Ee/F7rokiDuf3VAyMPkrU16kZUbFxWaUaXiSm9oc2okuhta1gqeLPeRM7od
/8O8VQHv46gqpOnVeBSYoaDlhCYZ0pDu+cXJ3scvAqPVMwF62vVCjk2jfROpNv/g
wabq8IhdWO57qgNCYg+Sc5MyHaQgN5chMXY8/Kds56R8OCRhGreW2dA7FVQmwiR8
xQ+EFrnEnyj/JXqYTtWztt5kOnmtanlz7MClpy78RyEYhqWLPyU6z8FDSXHsBimY
xD5x7jBcSoWb+eyy4F/DeZt/IKgWU5CncNMyW8v6z//rP3XtcCesk4C5ym11bsfh
/2rJhfb21fRNXpYd1y2uPtmIlnYaiNiDvgeouSFr7PyQ9BRkMJ8ow3LIG2ZW3dMA
s84VreeV/op1qySHBqXe6VamDPGDHlw8SBswm5te9rtFLSkPf7MqJlnbi4tIMgwu
MSzsgA3I3Iwdf08iVX6MVlLSoVm1rA5HEqjFQDLd0/KcKYJHI9fOjjJu1fp1cZPp
X1OnliJpGZtWg1yzytVJKAlr/OfBfQVXkru3cYSu0AIWT3xAT05T6trgP3RTfv+9
xj9vFuefuD4VvgBBtWL+W/RqmzNCV1Thurw2tT0y+7ct9N05McX8Ib0LPgMjw1ps
flmDmAXkMVjPWdmsF2Ty4TaXOD8a2xagS/Ca9gyFDrdRp7FW4il4GxnJQWlsRzJs
Vz32GR1wy8oMwai1eF3hDLSDy/5NvZs4RtnjIDWVZdHY/8hR5RBArqJA2H/ZgNEo
cTPjbO/sweNPLW1mwC0bx4V+QlvOdmQXpZgBYz11WD6Z+R5yR+NZCqUPBGrsZUoF
0m8MtKNuqM9f63W2GqgGR1PMnsDRU+YpVs4oF3zvuSPBqOTd9Sorlmq69bziMetr
OTo5limcL0ANs9TtXsbeaNjaZrXRdVNAnQDo1Psu5x76nc+VwkFMEi/Z7merK+kg
T5TAwpIpYQLkW6xso+hoOGERx4eTSEDUR55WWUsRmWGypVwySZSmFTeZneA49hJy
iO7NcYlPhItnR/zc1E2rvJLsVPzSI6CfiteuOpOQ/pYZvEn80UW9l2bAJvJ/PiEY
Kx9ZCMJuIRCIq3s4UUXgxKuxiiJ5q+o+7m+fDU13suJudCZYU/CR7Njrcu9TiIw3
7e0ZFZ6oAmP9O37eZko3Hig/rHYD+C7Qt3mUTuWqeg0IbK0K/CAxxaGGSjt2aJyF
0Lb22TophLn0mG0dOjay4Wva85NmjdxIzbBE8+UELBU+DI61iGza+oRNNQjrigiV
sEzOafBoR0vwf4uYD13vejdLfb8HAKkipsc2rxmJS7Ub9RedPTxZKC2nY663QUoQ
/voSpli3Rmbp0HYp5S49xPeAIsZ52yssJoTXAVSR5U3Q7PjLMxxn5vBk+p24ZBP3
eaDyOk71UMv9s6hPm1U+OcLSj0W3yA94NHbHPyU4MhCaNdXR0hpRMXQwQcuSrefd
k/BTidF+SGruCfOtJS6S0KNBoMJ8a8oKZtdg32skaAWzBqtOsBm0h9HmR7Sy2qgs
tUe97gLhWfz7Kl2/F1wzjPbOu1WuWgr4r/FcfXwBtji/OWXYmFClkCNA9g115NRJ
f9C/NeKrllIhtPhzU4dR4/NzC1jLUpAChLtZsMKZz7hMEFSlNGoRA72wRTA359/8
2i8qeMc4H2U4eLxCgQm/nrjnRwgFVVLRuSpudMjFUa//pRFtyWFsqyF3Uk3om48S
z5BJ061tfIYdRU16ymiS3z+kXWyspVUg8XKwjIi1/xSBZ1buDoLHzuEOk2QpK/A/
vPqJVfyhAFG+Y3sw/EkjQPAdUoZo+9TLwrPiGBL4d1FQK6jD0eFbUHihh6QZ3dU6
VWEkq0rsGxb3XIeJCLqdI3ksIUze91ioEkVWVD3N5/19XnApsSSEqzQRtnOzvN5I
hKe0uQ//jCpbW2pEVQLDxvJ1gN1kNLRdoAk+5zx9MbC1xZIMoWYhKO3PrpIA1rwx
kFZ/BoV2uDAZg9WPSYvTDzY81oVy49jZZ5H8a7PMd3a3D1T07DTJZARhEsZtbOJI
NYVtnNPoxYhQImzDvpIB/B72vSXv1trSjef/VJhB3dycWo7nqcY+EOPAA1DUuBI+
a1kh+32WwcYKQpvogMnb9+o3Gj+5BuVT3khOWskNwUprgBoZX9JilMihZAnh+EPH
jhClJHOKqd3N7xdsLzsARxAns5ZUkcAci9G07fagrT2lvyZbab9DSoxDvtEYLfaS
Qz5U7uP3ib+YFOF6TrvGW+cteOVxC3XMRu1wfKT3N6YNVWiBuLLDKhk2AQ7A8xnz
Fm5mumHN1VQU4ClhAsW2uc0IpBpaNZiYqwCS37NIlFLbpVtd53S7JwHwHno6Qq6c
1cqaLF8I395V5fCiCmVk4izi1wo8nyQTENy0WfAlt+SAbNaQjSfDCJ9VNeQ6Fp6r
7FLdi6Gb2PtbUY1Uyx7LFsCWlAOCh6uUiEOUqQbVxErNYDK1QqIiqme/C1MjBK+D
mTufixgHE0EOSGkEkPx8jfPVI+XdiXtI+hzMfyJtHy3f1s4ILIhylCIND7UCZrZz
sXlx127yMTL0Din2xjU107xV7buCkSd6UthOIMraRg/H1frZg4mnOhOsOcWn+k2s
zkjeWtYgqyGolOn4/k8VR7uyiXzaiyUH9yi+q6HaA4wg0662r3KWEqSfCOZqvulU
ly7xubdTnE1qifizM03LwruOWsLSGLU7fvXYCldYTo6f2HjhVLMd714opYVrNk6d
SC3qU3Tm86DfyGi1ICFkJ9th0HtzRiCRD4KU6FS1Sou/yEDm6+iuWV/k4V64hMSS
8ys2wH+duozC2qFAYt8UKXYl+9a/q5sZydsGY9jYEVttbRlWwlcIPZFfxAF8TH+B
6PBPaJNeIqXENBgfjwkiLUX7KvCyKZ61t+uEbWFmv9ubXEV9BvhFJ9dPbSNi4n5H
bWYZHC6gZe2MG3d0YdmTQSN2qTQFP/b7EKqyKKTtnJNHgi0g+rA0YlRtXkC/Ai5j
VPCiOmPtgjxn/z3Lj+T0nbGa3Qhtx2i7iKOycMsbchjLRrn9N4xtJpdaV3tYJD4/
xbOXy2qm9lwvsXxgfYWybLKDKISK8XF2BIXZ22sZxP5nGyaGPRXQ+utUaI4t9dTy
MOx/cw/CCD/H0JZyVQigc1iZXBT84mHqPIzY+m17R3SsXQQ0Y9v/a6mAwZkYngGY
eGPQyFjOydqTS4pJc4ArMpMjrMjaJYpAES2l/hYlXMa0RCjDqWBddv1ZYJDF5yQ+
c+W0MWF6dQ9FZfarAfXg9DEJm3CQbC2MYxUItkfWAm/zcpvPY7Uyb/zOJDqEnRUR
Ns54ML07k5aiYnOQh4NxqsNXY1Dyrt/8C9wFxznBtScWTiD3V0wEf7wjwex1TjiQ
HdEJvy1cmsZa/zsXu7fJIYioHa9GCQm0RF7Oa5ULJIIn2db08cW8OPfIveHekJhm
3jifPNDpsnJ8YJYqldAA0FvPow4rr5EWe8HFEaIzv5fQVD0Ugg27o2LYb+V3FjSz
WkdxXeDcK5lwUVSbuaaiCUGNzmwP3Xk3ZjgerArgUPdV9bCJ1geanXjfQUp16nfb
EMsHFTYQLDFiBm8Uu5FFyKzmEXDq99BpQNFYXJF8pIWX1dUzwWgRcdsbSZr/4Qqk
5QtA8857L2f92wOgjdMjBLUtmD/RPHj/wuERqlJv06AQW9fcWYb7lqrMjdnvuUEx
3TQGUW+I9Qmt4TmL3MNPdoiA6Hl0RwH+guLhhTp0zEhewjNS2puxRuQoyL8vaKr9
9GwV0VinnDIC2qPur/l3hwbKir+b5KddCTc2FccVg9VnWMb9pWAvNV68zNrTSwXq
sw1ALtNcStOgmbT9sMW0LhxHfQ007TVtCKLspY9OlhP95KoKqKzQFqLQFrQeA4d2
CnzOWbe9VeF17pr4a1FQebj63EomeZvsNLeCql/BJPvUnRPgFnLTk08SqvSW/Y94
59MoiQLMWjFz53ToAXbBX4oeCdbvA5dgQVtcoWiQ/0E6I7h4QsYOgmm154xxMh5r
z807bsUteFVytosTUaMEaS8bYseITn/t2zz3zTtUpI4YIgTx4LM14pLPoXaT8xRH
ZS3E3+Ia502CTq4/dfyDFtKmP2zrKZgm2ZKzqtwj46Z14zGt0zq7FhzUt+PfS6hy
BrhIpFIJwXWP731yQuyFdCSrh3ZvTbIyz2QRPx2/dDqfGk8mYHVByB65PBef09iD
UyXFvehByENthBRvfPzpus7SToqfLLXtr+dNaWQiwWYYZQA5B4Pm99UdfCfAjEyF
kFIrgiSA/0qUoV2zc1AyFApFnwCtqfqmvOv7iC5AvvVRnTAvEnAmcKZNEflfv5u/
doQvTiwI8mpynJbiykX9m32OqnRjsjJ/+Ayaeifdn6u5IAsjDcJTvNmhYXOqkQM6
VPqf7NTDRnQWdo5t3YJVK/jR4zVLrO7EFaNCfmQFHOIt+hLJYo8vMoi5o/be6RUz
ikDXgXnMh1o0Xzpl9e/eRlrXqUK4WoksH4MCQkahoeU6vi8sY6AXQIqCOYsFq7Fq
qYvmz/m+eND/uHf9oAFqiFofy1T9bvz0QP488o8VNfTQQyy5OGuueMc2QLoQNf+E
UtWZJiMfaVtUj/el4kBMKdtrjU6Ym+V+yQujVniG3ncOd+X9LfdVB7FECJD8gmwZ
lwNOTs9W2ICy3tBfJtWDE3t0YIEJ24PAHINwKWsO+E9pEZTNqRZScryrIXLTeF8t
HVnwZAihN084xF7+JKWwzMqI5OwoAYNy+OhZMqtCxMyzQ0nTG2gn0YEPIqLgNSu2
aSja7sWY2GU9aNnRXbtXnKG+cQ17Q2dkaYvA2fIHDTYm71pgeEUb2hdswXdmmLkp
7RVepUrOfVMbIUJMye1a6PxG5cmTbGVmbUiR5QLMRVdHuEXvkkUitm31Bkw6qpps
o6Bfil1FW05TNPdrTTZmf9wFQIYqwsLEA142+Vkp/GAQUNhaVhjaQ8Bn2oUAZkdF
iIs4P9p9O+P9LIbpLspIDdPEVBxi3jz76eG2C33dHxQpaGV/XlrWsZ2HShRWNCWt
v2aZTALTlAARyzscvKWviIyZAQoUhPlTQpDZxI843l58XknXkm5rCeCyNn7naizC
+uX+fhUO1aLtMC6q8CNeyz8VY0PByQtrLvtg+NPHtGjw/VyUNaqsYqoF6N8UAM7B
1+dMLsP0Z8/V8S92Vmte74zY/Y4juc5XkVfHPJ4HPg9fJDUvjBsS7jIDklhyfFTT
mYwa/AESBkEECW+1tE5cRy0ztFTU9JYoDol73oMldIKIV/N989hvHU3JCmhKATO4
/SiXDfb4FNyomON6YnIIVYZAgq/WsLxKNJNwgFGxcSjdOPe6E9K9ZIUYapfUq84m
ZJylWnPRcSnR021meXpAzEp0aistMq1MJgd/ndBDrEq38wn6tI8+eWV3cp6q1ayq
0TFI9WhaXmsRgKL2s4snQWC/XK4sgSd5zUlvatFLWGeLTWrxzZxfTAJksRHB1tff
1vfoNgu/sqBpcjleUFROcFf4fvIGboacBgbMfunlHn+hQv7a2vrQLW1spVidN6kR
LQiZ2EH1k0cTg74KHH+fn5F738TtVzALuSHMjNCpb7vyZz2OKLMSMMF3PIgG/odv
FSX3yS2zujroqRRZ8bm3+FLUH01r7ETihwwvvfY0eLloOuBb3YDft1/MsvSpqCNB
6YYL8G21CS7SLqzje2kbnDW5ao/cq+2vfCSH0AsQ3N6VIZxXQWNEZPlqkI5QeiyY
Nd1JCRAQ+jce5EW0DdbFKqR4hcYqAr3rOis227mZ+j8SgTsE5jzbOGV1y/P6aBnH
gO7sa6W2H33Wln3IVy7Ydvt7JN0J3IqbUtr3TS9ZjcsQ8/gpveCJx/NEl7YqIfpt
WzdIqTS87gVCp3OhHqv/G2WeG+YKW+hip7K2sF3mZYQ0Sb6nq4BOL+DVidfRbo6x
YszvqwdsRxqDqZWGExtZIGtqIvF/9w3cCXyLQMO4nPwFoUlv1jcRbtqLzLw8E8tF
l9RXRNSvgTNnhhtw7uVRb3UQ8PnisxPL2AvItMz6o7+VsAoi8/llLhHlAokECX73
vDl1KOoTgle/BVIra4Z6+7GNPJunvSRKCXMIwRNbsyYaWjONUf+oWE0sxkQRPAfr
Esf5MnFcpwZGFSB4fSVN6nwMhADvYTixGu7Flxto1vqOgva6uuqktpX39+FGZh1G
iOGW8As+XhXR6/yzJwBo3Fj9Q+Zg5+7x7OTQqb0ctrizN5BbXpfZe5RjGzkHYQLp
3qHVifJ7k4GHTEr8PYsccy3Nouz5ylXmzDTNIDD8Arzx75NSRYm47gaLXTrLarkK
FrbznkmRA5v0M+uHbZxLojDjr02UMB4Pr8tm7JmO+CODqQL6iBuRu4Q+trML+HOD
c8Bbfo7Bb9vgl7MQ8gjeZnbXfbyGqhS02hI2rI1EjJoThvYU1GnvRqekhxu2CI8W
bRUettOu5JUp1tFQaEfbEAOXOzbkRn/gQhhGrOuD/o9oLN0Y8tPUBsseQ8Cyls6v
Coht8czpq0OZOvDs670NPSuck0oxJSaOrQmN0wLPE8iVK6zRNSdP0g1wWyFU6ylL
Hv3YdQwTCAYXBhEwVWhumSnNg1n55+G/PUwQJFNxNi6hRtFGGl2H+DWAXM0+pBnD
LE87RamN0G32VX4BVCyeOGRG13+jTzerE6HNTNNVeijvBcK4AZNx5Eq1Trei7wlk
DVMaWO8bwGCmn2WqwDOsS6Hi7z7l03VjSimlrsc+PjhP40QIOLxzSB9AmWWnicG0
+reYh4JHOPVBDkofySiS1ZnMr4C1Hqc6N85cr0bsyR8P0b4VLh3LgKH7F6ZOUovI
8dGu8AtzEJhJMvUfdmxxEnaO257EBervoQMz70Zg68RQkfakAkid22OjcBRvN1Jl
rQqe39MsACa6QlNXzO2Mdz3rZ04NoPSkyaMFUDEYhVIUJi3WxJZrjEuvnw2MsULG
HNNaxhtitkDJqxnYTVFyrhC8wOwWYSejbsOpNBnwQKCO/J9XCH91Kbezloov/oQ8
vAuW0TK/da3nOdg/mUg5izA5smJ+WSTZHnwvtrqTw4rNQ4I374THPt2Z9u8Mp4p5
3NlmjdkW04lX5fAQQb4+yTpN69dk0jQ/Yus5Xzbo/tMFHb+uZITqlIiT/f07zz2l
C9jxhfME3s0GGYNWB0+6VQeeQ1RrbfYtP2+5lgWzjJ1fMIfXo2uBBVfuSW5133s0
CVw0JyrMoRNMYBuOC0FwLJiMwjnaRdumywT53rfK12OyCwxp5QNwslCqbIGGsQIf
N9fWH5pT3ci+9oTkZ2/O3EuRKMvts5RCl56qSDnxi58kHR0W/5D1I5T6bMWL8O6t
YUsnKBno1O5SwZfBwc40ipMnq1OUkzbEMyZk9bMortERcwRhjk82V5WMpNBg4qiY
eacHhfqKwAxltOZgJpCqy8+07bcPkQ9Fj6J4HiJDyu4u+lPHsocb4Cy7RNx3YxOG
gWRzt9MkefRqgqTeV0PM74N0pAh3rOJDsNjo2uYRlrz6JvpKeZ5FRX+dkUV+b1t9
ediir9voDVdQ22wLlaV68DpinrZa9u9n8N5BIhm9YCW12K2fcFGv+Tlb6DQdykCs
IGLCFO2jC78/7+/bJnvY8HALhUY1tR0M1D7/XgA8qyhFKT4JUhrPmnA1gsh+IceV
EOhInbLt0tjutN/hfbZEMik21XIUGcOpAe4v+td8LDa3KHfLLKMML1xQJNo4RyaW
8RicMWbAqObMHlZh6lMPJC1I+BaFVsVBKWy+KY8g0Fq0rJQGosFlOi/HZ2jJhqsa
Y+nW8Z5ilqog2YfLmd3tF5yDmEMkBsMTPVQeabHt1QfnlV+zQlaF4snfYZ4X23LH
QrvlyWGApTXunnBG6wFTMv6f3422/mF+OrYEpLWyeS7SUZ14Wed+8mURc2sXFQ1M
PgneYfcFx8RoVIC8TQDZhaRn0KWKt3x8menndQRkg52ynPtWPyFuc14S47bTRML8
98E+r4PkSAhdHqLuk1uS2IIccoimUkCSHksfPCl9w3zgCnfHj/XmPqnvtxGEcy/8
QFJQrm6bQik3n7x6wkb1gP5jkek1EUh/VQ0QM2oN7Vj8Jp3WeHZ/OnkdXyRkbHB4
QE/UUd29yXfLFl8lm0GTOgFz/rWpOUX0ZsVRWBP4SCGaLBQex5wilQDS49Asb44M
EQU/V64KajG6lKzps168IVyMHwDczbziZ2YkiPt4WZUak1EzZKrgLxAWA0gZeVCJ
rSP0MW4w+f14kkodj0WQiEBVYIQE23CrgN8JJFy0k/NNDMrNe2CbsQebQuqPK75f
AmyzNd6mJPJYQFHW8v6JdDO5plXPQCDOA0YdoDJ1HJnew2jSePC+gbVeKhFyuZju
HExkGeYrcrnYAZMIwxxJ2PyAHZlroXaedsMSZnJBkSD+uh5GLn3UrXFK71wP0Ey2
tphAp+ulJPk782hPC341JnP7RB4eavtV+iJNyHzxm+EO01D38Hex7AhopYIuBi0h
FhaBRyu0Xwoo1p69aMe1hYFDxNIWwE54vV588N8UMrchqGErTBPTr1Qy8ZW+Y7Fc
9huEJxSFrJcIlpjvp4LesJOxD7CIzlKd6xs5z1xa/URcRtlhdNFcrJcDzalwsXwm
gyngw2Ez2f0FhreU8GAXywFTuimWLfGVsdLfSSrddySUtPreqiKNdJZEjQPJYlYy
IzSVax4joVNPSEiCP+VkDMn/vGfaZscSdap+B0ffzBjL9q50YCztMikn0oz9p5b8
fz/TCACWMIKg+mwzTWyIX1H29p+KH9s6JK2cGV8gqbAVmnSrNvW2JC9AK3I7IIjm
48Pnc/yYVcopRzq1ZW6QenV36etdaF8ljqjPI/X4zQL4y2gRcQoTxLOVTcXO4ru2
ZnsWs4rgg1MoFrh2lOaBpM606+YuD/P64+ZENzRRWqOMyQqNoCJEwn9Iwzr+CfY6
/mvFPwuwLu6thMKUt3UiilGhHiDSIGWxoD9/6wIZigzd2jgyqhIlPYQ5RTXSt93C
FBnwIBAuYsetrWGMhIpNm+1D+zk7TcLBUzcVNaYIWqrRRh7EdLGQDK0I/APcAQWs
52miCkytbEOCOWRXqMh12ELVBPtRpNowra3JmwZfQpxdlMbdc0VRI8Fypn8paBoy
NSNv1TBRu5dbg2TWXbynqGam91ZeDygTbYWDEelxvOl0exPJvSJ1Tem2rRaorPts
GGm1txHq+LTZDj1zeEMEoOM+DfxqU7s9DPQ1A8htTKJOloY9W5p4zA/Vs9bk5WdW
ID6CnGhxOg1O+w6e3gHthFTrNY/YkgeC9LI+2DB34O4X+0jxbGT0egvj9s2//uor
D1TiEW/XNskUxAvD5qvKuOHHC66zUzsMH0q4sPmfIKabiWnGtYCXnXUp6C8aReGY
5EUbBWW+wzS9cgx6oHA95ffQj1cfivwRqXyHxV2RH2OhllHNRJMBPDBkVdgHHfYd
vCtpBrBp1Q0PdLakD2IgMSAmYqVj0gRHqozIxX14hKM2DYtqJ3eVjSPEIA4TiLgM
tgfOBN3GQXUqX7TDOPuNd3T5R8jD3bLi7K2bkc+vrHlxwPKzcC4+Q/UMmeK3x7LC
pZGnby7UslZ57xrdYscSC/sFZEnbv/j5RDeAfOs5wVlHA58GAXVToXE/SSvX7hpu
BocXEOtG1OhOzHvj1+OdCoDdLZ0DlU4o1CI+Dxpl/NKqwqKC7i/2DSSfPCW6QUpn
dWtA72meop+b+XLPjU+OCi+BC104DQ2/NZuBAF3RSe67S1TztiC/8KIiBC2bUwCi
gKzrdxj4SkMlMdHjAhiiuKU4sJNTkVShOSnq+RQnpH7dSOZBIA2irDbv6pZF20wI
3OQmyd/2VsmXUJaA4WA+uTkSKJmz0pitk/T7WijiOT+MpMWqvVgPWlTj5bsHVhrl
4d/QYOmpHDg9M/+bgo2X31HCcfgLctlk544fCShwSGMI6ZOSQiqIxdvQEVr9ud1B
YoYtaUbIiOUK+d4hlyLm6RKdBQtNkQdpkvfYUZxbD9DcJlKj0xOCzwX10wRhCoTJ
Yz8sVEIm49yUd9GfPF4HcZuASqIxAt2XoPQWJpUnM7ilj2DmdWhQfvDB/KpoqHAU
IYi6JvcwnembNQage8ZkxzPXHYAHUEGI/2PvKi/3jF4BB2tZH/mgISStSVu3WClh
DKuM/RJK/E2OdX2jvpYY1C3vCQ62f5s62wOJxIf5+N248IsacLR08uhEAgRhG+KW
xqjirhq7O0+1p3leInHg/3xIlOzOYgDIOl0rTWBePh+EvQ/kyO590D9XjUsOovyX
WMWt67c+aeO2xQ76m68N3aK9hImLYJ5x1LXD6exo3tBUS3OVIFe9L0VC4FH7rN7j
hKDvayi02QPYcmDUmLCC98AXlw/LOtOnsdjTjdYsaHrx8GWK4jPo9g4D3lTowqb0
CJqY4Zhl/9FbFy0q5YjGDJzABGRebjraWU3X3XRDll+fb4mM/ELJGsJgXONy8TkJ
jxiRADED1iwgMe8gPUlstn0zahpPg1karK5iEWOsIIMMhSrkhm32QcMRXJYD4EIp
ExC8NKDJf5vhp0VWn2Vx3WXV9fRqJejs71UTFv+kiB9hlVhRhVd/nBx+tMeHLn4R
NcUqKZDnf8QJF90NlDNXeykZ+8X14xAVP2C0NhNQzPPyrPoF0zgXWNGP8TgimZ4h
IBacW2Q7muB59RIUMBVsS95iuw866ssIyrOpsWmrIsez8TfLwFsX51C0DyCGDjAw
kmgcfrQKuxB+sbkGLMNmXVJ2SRAKmWWpF5Xu3Mmr5U25KS1j28wzkkxCDlEIKKrR
db8tZS90vIx7tYtwCX10FDv/hE5CdvulxzBz5k1CCN6471n2M7PEqOMOc7ReNSnA
cSQuKfXYSIPyVlXG6rNZe62IhOoFit0GS0P1zoV61anM/SqOH5cpEEhxmNhH2FH1
aBsd+ObRDaMfpoqD+qwVDYQOyOuSttg6KeLD0z1+7lb7uVPTuVA2bXiThLubHZ/8
YxpxrxypndDFKihc81Q7rz2JvDkcm852MStZmoTd6ONLUEi9S/CoHQPlW19wbbRO
wjGBC8jVF1m0HXUjsehOOV11RfLIYUctyf/hZx1lmOQ9vdCWiher3RPbTNicoHNw
5UBabYnzIs5pMAyECDkZ4s5XkmF7qmAYFPnqltLfRO5kTtgDIh+4jwVAS5WTX4F3
m571k4zHaUSvcumpQpWJ/2AgBFFN1h90r/CfcY5wOzygLtgp5UzmwF/3zKoZGjGx
csJdE+K+dsQAPVPE/zPPUgNqK6WBue5FfR5CPu8TTuNNv4R+pqPJcAMRfeSibfEK
zzCSFB1RJGSu29GIGn+2EZo9k743/97BaWYEExIWGG5Wm0tEqEVbwmDMK/jCjCub
5M/vbNQ5X9VDXntKnCnL6MPKyL2P0ptUDmqSx2C8iGXMNNzEirgnf1MSba2dvLfz
yOz/T9ctmBLdz7CvXNUyUNTO6TkDHHXRcpmYSkfCzsSuZ3QZ0VkfYQ0XMY34n28C
v4iysfZ5/KU5a2xmxLzi7+kUtHHSPi6qnW/iyNG9+QimoHRt6/nY/OO2iuvxugts
j8IM3Jq41Hx0h0KmUwRIXBS+pf7082BqizOQXWjhdln+0KdBU1Wf5qgz4hsXO5wZ
oax8AiwCvBIQO/6Yg/WFWg7Oo+Vhf47Oq873+KDZmny9166x1hxfd/NMDC1rV9ug
Yw9RlvttAkhTMRbSesSQj8Dir8XC3Me9Bet3ME0dlOqPpAtVL/o9uZd0ysftQugD
PWPX1FfgMnSifnczXcWJXcouPxrmUYwUs1lmxjAO8ASPbLWF9ZB8syFCC+emW1M8
HHqY+XcYUu0yTNcE7y5x3OVzJfv0C9eLf5TOusaDI0qkDQ5jHZ3EhjUQmSFfAx/j
8/Ikt+9n7HkwFykxy8XYaTjJAqzRgk0CgqodHx6K8r8MP3tKPradh0y36UgP7Brn
9j+mfRnE/oLxjezPJg6w1pEsG8wgJbUYPiGKg+ok8nZiuTCVxB9rch6iNNDOtEZK
nC2ztO4HpP2a7K43JxqzcFADE9o4BRrF2FbgyhmeZChH3hl70M+rWH3SoEJ7Dexz
g/dP6GtbQ4hjX7a8K7cVFok3Z1ml6fwhBFwp4U4Nm7oENgeus3JmmCFY2yopC9jB
BI5uOCfe4FqhXs2VeRdktmOVNYCMseOuWqA1lyw7RygRiAWKBR0vEiXxfcwwkDER
oAIJO7vJCk9QaG24vnLEnE0atOBg0b149pObFWKYogizW6SLUFm/DBZodmisRvZu
hFHQC/4hPdFpx9E/2Ek5uJp+WJHwpyrNmRj4wpg7tNqv5croyKpLgL8gAr8GpDGb
cp8wAYMZIagh5fWmGI0USEixssqCDHf2Ir1CVzYDxMW4ryFP84utTn6R3nTkddRD
7M8ilHywfSu4cq5eUgZpvmsIztLvpX9YukznILPX70ps1B3C4o01Kx6/vb2AQap5
CjmJtuES3wYS6zPW4mjkuVy3Ma93q1pXEhspwKUw7CNUyvlaM+woHsid+356SCg+
7vuUBaXaCXkwvcRRhky3dKY/gkqel5yCAor8yXx0i/t0OGUJ3kCtEwVib3WkyX9y
ZoUya0Bkkov5ejmgKcNwd1m9zzhtJ5wBhi6g+pn0B0s9PvD/Xf4yJn+EHUcmGqZ+
AU2b+MTGAUYCJoe9gr3+mZpOhJfOH6VMTc0mAmUlhr0hieswESSOzx7HW6NgH/EA
Rui8QcQ2bQjA38yelW+JCduouBtS5igaULLazvXNH/CbqqULf8bvxfQV9lT2JIUt
mA0zCISjOlBdd2PqTR4QDNH9TbL6OJQ98PKvWo7/cCOJcboPCA4CL2QgnOTXGpXH
tO2jYAxhZHEi24CtZkoGW4pZy5X4PsqZAdC/Y3uFnXtR4Y+A3I7DoDZKsrHxNrfx
N3KFZWy2Ulqw1SysDa0YT8RrwIx3KoiZFEgGqdyypASQf0P0xtPBuTmu1Fk+hxkl
Q78Cj+j/Jk7mPhXIFTIA/fojyMVYcnK4d+suMZ4M8B2ASYxy1hRSoWyhKNnQZJxh
chWZ0/3+dSrx1f/mvfqzW90+bnRy3uYINmEYAQ8I1RkyqB/+AeV6Yo0Ef0yFqy4D
SHYrCVZtNtanf6xsCwyQYNPOwlKgg9J7DqkGNCSWhPHW+zDfbv3DdIjETHm87uGg
gdddsp82wgXE5pIgkgEd8RRfx9OJAsc9SCU+CvlsjlEguEDZTwXxp45wq/fFab2z
LOW/CB40aOAIVk+V1fjTClKSRO0FvsCBS/KuoW31durDsFlap2Xo9Elxbu158g72
+hbecHACiiuaTNZwKuIC0ccK0HwpJgV34NE/7ECklXuJvV0N9fOLh9cJWkdQdx7z
fOAbzlV8zzJt7kOOnZr4b2o9gInt3XRXokM431HVFQ7c9MXY4rJ0G0RdLsVBq0DR
pRT9Aa0Qiuov/PjXbwciRlxL8l94mYa7yFU16R9oyoJnVT5SIjADJQo7hNJHQw6E
/f5T9U8tOZd1pW4iAPhtCB5++weGxini32/pnjDxnXJFL7PaL2/jPg7+YskYJG3u
t0BKnpTHgZVhEVAPvBa9VDgP94TdlDxt+tPfFS1K8+elA8vIalwV1YhAkdby5rXK
4cMVD0RnOys8fRtGp3B4EYvDVS3Jk/h6flNThIkOTmES2USNQYsT6md9UuvLvdpE
Emo+ODm2EliSSZc64SnUAPLyqD4yh08whItMesA8otSutFrhntBDChV67pfZOxrX
/IQkTRm+MCndypI/ATWjI7E2G0kFYg6abpTBjmX+tfNX9S0ZT+lFhABxOEm60yHS
rV6knhkJlbFnMVV576khaiTqL4hWdeJRHtHXCciwuNJrFPXTunOWFpGCgqkiJuMR
9i9wfsjySOZMtkMIzsBOKYHVV3uEIbWZFORwniZ1SqukILAkoK5BSYxUy68S2kFd
Hg+1pLbA4vvZggBWV920ONhrHh8POXC9+L8/QCuUnD4tKiBqlam4Zo7N775PxjTt
jWce4RR1MQAUcAwO0Qh/OzANLfuMpopG2w5ddSVxnAKNihnLgoCRCHmSqlOKkeng
43e6LALhygI3mNwf2zarnVg+oMHYRdu/WoWaKMq7opAL0gHlKnrOtuV95LpiSEbq
FGuRJZdrVVBDahOQvZGgXpf/pKrhKqIdxlsZ4zZBgVmE3IndIvW397WaPs+ldzPs
zHxcknGYU7FFKPrBm6FBZWcLo3J0oe1JwzmA5inHJpZUEjj3cY2YXbeeZB/UM1vO
4wGkvwDZ4K7TTX5gn4re+QwslfZyLrIWJGwGHlEcMtPnVf19/LmfEkxVgxK7KSE6
hJR4nMPUBQrhS2LiFLxbxS6pmlJ65jxXbVxaZmoxLNwbwbUl7qdhnWC5dHpxsKC1
hZzatLeDYV9Tad7ugW9ZlhGXhry3+lcBP72SD4vPEK1Tya7bNLU5nHZOWbkJ92ar
N6bhM1mQPBiaghTxb7Gu48zGtx+YzP649M8kcuEAzLIz2hTfRO+9wYmr9ohYPxlu
wqCtrpJHW/KQjyH4xb7N7EfWsRfMhqneRrMMi5RbBy+jSCdqk7r1N2svKB5rLBJu
szYqvllX60oehq65tza040+dogfa/y8d79t48a5rS8yFSZoC0F2CSQ9sBvIto239
1jYX9okxZ/J6BXqkItqgIqGyljjmRnhz6Lhie9gkpMSiKpBFQqZt3W3WGt3NlKlH
qDSVugcDWNhBCg2xX6xGdM8tVaRPdriILKmPs9ekCbiUNpz+nrniZ+hZAptPrJ4Y
XspOqMfZdyJ+8VbZsyYkwH5hegpZui7wrrqwfsipLpOn4AXBErLxdUjv0ZtmfaV2
pUtSwVq1EYxKe6/KAqQLkF9MHUewwhywLsF13IYzt/Yn1SigCZPtsfcG0jRmOTH+
zrYMvX8feOU2OxAIQck1lL+gaVYK1A5eZlDR5H1D5T0N1x3z19+4XllZU9Mrd+j0
0TvXaJkiVBMt42BOY3qC/Kwt6VLh4a+HE2pZbfQCSkKaMa30AkgwMiCHNYJkDWuE
6Jyky5o7QxJyfDtWaLih0Y953/Nsk8HSqAu6CA06ZGrECGWvEqjTDiPvvZnZZGRe
/16xRLmwKZ83V8mx/PBd3sF3ZOa+FejGhc9g5MRCrjs6D3VPy7qvxgCx0rSuoqQz
qBNxbjHADhEZEjHfrZnr8B8Z3MiXSC8+JcSFl/lips7qGqFM1Ek7JrjFZtG5boYl
h8pa28PwYkEhqRySE469O/wLCKCuq5t1gnJPHl+JofcHuWXEHHjGwshkLxYGZQWR
IXvpIwuaLFzvPxvuKa/EH1E/Rdm33TKfKNWd2OgioBEMKD/NCl1i2kEhcs8Y+k6u
kSpnPr76BrvwsN9YBhjrTUX05nUMKIlmF8ydXFJ8VoQpz3fT+fEq7/FM+OxU4sDa
jXW+0uYMkKn0Ccf+cUjWUOJXQXuZFrWRIZJPu5n3HFgVK+MpLnNfFah4NAk1nePg
07FJABRXKuV/DcT7aKf65LpISVOEhodKOubDzkBUk4/VZ6DITSAWiaKGcRrKi8TT
4ziItjE5NFmDX9tbCQg4tLpvnz8XwNX6FkNa6MBSY6sWE3MNPplpoa5frEeXJm+l
GP2AFj18t98saIROIZukq9/NsdeKp+Q30MLcVGbjp7PMRDz4K+1JSPiSl2h27yM6
Qr0zFk4KzyxUHqBinQyglXU2xH00tDhHybu9CR+e4bqdcyvse7uuVhOsFF/zLweg
D1qZZKz9u5z2G1R4A07/hppnViD98bYlLI9/2RB0230Aobdk3rOcSEGUvVeGu4hF
HDH4VfqbGWh1PVlB/KsANUVcPu1ClHRajFmFgrsPZAmcmOyCO1ykhukJ//8gz5QC
FX0oKkbymUVpfhqEehUdhOK491utF/c5utw2bmcQgN/G5fH4U74rBsVZeuA2hslU
Rpp0tnFrzFCPFkq2hZW8qkz/1mH6/8cRMA8FV77HxU4qIIh5FwXNjcXYn8rwTiyX
d8XcywUkvTQsm4cXTy+LVkyKZ9CVitvnFSAqyMlN5kJrZVmZrVmTQlq+DPK3J79m
1AUg+cCCgZq5m881axnNfMY++3lygLfcJJZrQ2denU4pwIs7X6AM2SmnSXbyRebS
gfVS/h4iBrPSlSaaswzT8W/GfCg9D5ftGOeoJhh3kFsP3GyyfwUbmkdOrYFvkkAW
jlNPo5XPAHSB5RUm6a6m/a/sVc8hdmVjUlfcr5Bho1WhgYM422g33JbbBkJ9LUP8
fZG3+RKXiHyT1JsBqn7FeRAEeKdFY1fUJX4E2dx4qNm0qMl9TsVp85cAzo1MNpis
L3CyjT+Oy6BcnZjkS+nLvdpo1UUhT4uHoxzaZbk6stGAH8TzvatX1s4wUoxXG/kB
O3iGQZsI3hg7HEI9EAUuZPattgBFhrKNvrC2ejBYaMLpAgf7gmGBrmVEAuW3rzOv
aJGINGRJg1NqftA3eZTyvONNBbu6Og91M7y3OyS5zlahmLqOuJs4q04Ts4FFYOez
wl3jRuPJTkTz8TrUnk7PzLy5D3jDh8qcArbWDis5sAxUUs7XEqQJNPIyWhOWjfyX
myHizd4SOn1uMmeKMGVzvHbHN4QJnJI0HZPd4/Za2Ik=
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24224 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
lmOQgIOM5jiJrGbWpsW/8s2WYtKCWHeWK6lW2Yq6jSWQU81uvxzjiZpqW4gDFNWH
l5LiKWeeCfeOwueWpJfOBSvqgDuBM9sl3TMjptghxMOgzUGgdpBsVSpBSTF7mIdt
67FdSpsToUu/+rDyx3cFPJdJGOlb9nAkKgmXh5+SJ8Fkrpr8msW8qqekAvqpH0S8
A8KqWGM0SpIwq/hA89JHa4AFB0jFQ9emx0W2Zld0b8KXRog+sM+lL40S+qsJFSRa
Tq7f6aPQKGsw2I+u/nw08jPC1cdkt7lrDmnWTYGCtF2di92FxAqj7mZFm9yS4Fwx
FE8nHO4LpVDfOpHV2WyxhjlRfPgPtGwB9UPrSB2O1+mosolPMggZ0t4Hst3vexjq
Y4LKBMYzPY7aOABD6AQspMicOs6d61Cg7+iVmIUg2wZLCmfdzgEgbBHof6gSvXIJ
C4Hlhs0adObmSYUF7iFxxDjj3weVJoE6ZD5/thFl+jvp3n5arPWU2Y8EofXWETkp
kR2zoaxfFI2J2H/zXuuhHxMgL/Hdy6U9AV3uKlmkczLQH4fvaJh8v+Fr3WDD1DJ7
ws4KwogpzvTyZNglDw9ujm5qf3VJYjb+Dw8shKivHU+Sj2vRhJIw5a4wh5h/RgWd
5Ipu7ZINawW70kL07q2jfsH//9MDYRF8KfR1LllzvQMnclNIqQbB2prQ1QpM2O/a
3o8viOYzAVSSTbYHsXUjNSF4ODLmfSU3rC9YGuCmLvvT+RgTTI3+LRmfg7H8xuM7
FaXTd1yxTWvADjseGMawqnJXvrAD9fo6guMcc8xnXWttHnyTOFXLJVSLpIMdHThU
Kau/als5Z4UMY2t3s0+cVxR6UTlke/dnyr8Rzau1sAUGfjj8ftr02luuGxXmDcWb
1Wr8yBrLUxoH5oNiKDiJmPQkBajOOVBgy62InyIQ3tulALfPL6vn7M93xDcaBZjm
Mh8C4tIWYpniDvwpD0W4VAdnAm659+Sxvyy3uqh1BS5Wxf+nv8QudIM2EfT1por3
QmFdH0qI84mxxdcYyBr3lTKw4yZSi+hfj7QVCOlOamnkoq8bnk5CSfZc9LYdbEIo
y/F4VgrlRdwAVydBXTV2Q/clIpONlJAogE+FtFlHaFhKhoLYlmDdjdtOiHNlXUWP
e7EQN7BSBunYJMvy9+gDzxTCBV8TvJCqFLIBfyknSpoO6hR+Ovo6M/r8KFs8vvhX
NvWTxl0OHhv/fBqjJpv8WNprl58S0z4wrhKg1HBlPI72e/NOduQh8Nxqnjs8CAr2
sF2CCQHRVdCmB6pI/k0YTyIEAWuDE2bccvZRqqlzBSPzteHB3eM2KTgdJY/i6jnw
UeuHpsgTk2VuVBhXSM58phn7/ut+VDPOwlNs4S+rqr3UlcwKNYrj2EHOFcMASGS7
VEWm6vQNbxe9R0KVeEbbZ6iijyTI3eEKwxilnG7xSUcc3vRcmKnzhQOkWt0G2PW+
f8AWgX1pO/u8AqBTrBZ+CsIvESmVTzXhNNrWCQQ5uVZRTMPWHvVhsYuszWH2Ms/e
bcjveGAKOhnzGxaVtas/m5excjwQzopm3FWeaSzm7ZdQU/Iwn0eBV6+Cu8zRjwqb
Pt08tHL9FjiF91fj2lgWCeKaVEmIWApdRdIby3kKMZqFJwIwe5n6QRO44vD/aEyR
E4cXeHaTM2ZgxJf2YD6IwGTBd40pJygXSmREY6oQsOHMS2LjljoAC2dQ+AOdEV8I
O+TVk2wxznrLYYwAbdPbLRPDX80y34D92e0/e4A5S6SQxHj9Bn9uE8x+8Y7OVdKR
Y63rP7lkf2jxhL/zP7LhRKfvA2f9XTi5LzGElW5r9zhysvL2HdX1FBKPQ/xlqx6R
IkL+R9nAQ1zlThlxMdhCHdT9QKByXtwBt8Zp+k30Uh/EjRxZaegf7FqFrviJh5ol
vlqFd5y3wu66vtzOQpifvcUGG86IQmRixyjZ34yrGNqWEkU2EdZRdRpRR1srU+P9
oROb1qvSLX2EvzX8R5GvesfImved3dO2uhTe5UidytJfiGtKK+oAT2IqKS9B/Jy0
8bnPV8xMPsxv4nq2PEAHkKj0CWSQT61eflzImTtw0g755lz9oYfV6XgYm/NIP09F
c/4gD6yvkjkCEd0SUXHZrGvQbB7QkGMeJ3BpsiI3SA9J+UXZqQxOwxSYKEXUqwyp
C/SZXCalfSEbRcsK6UWw8Q2oPnuzqkClRpFYg2u/msPoiAW3Q9puMOJQmyvoln/+
j3sKpdbiu5Tzkv4OyRv23SCHke76PmDXkeC6lV3s12/FE4WpLwt2RegxQusDQQWn
+FFo+7RwZUQ7Un4AWEPqJX3XujHvUwE9cmf+bbv++C69go5dggte1ePRIRzRCpC9
fhuxfUR1dVIdQdTwuYGf0ZwrD5iUp69wckoqxPO/O+G3DFE8ZsmJhL4QDtQ3QASW
DyG/kG1JHuuaEYPFiLVOvlcn5h7/ShoS2SLC2JqsfJlrRTRuu4avHv6CKpzhMsW3
nCk+/lYNobmE3bGaWEVpf3/2hmL0zSE5N7fUUcm2UDd3WWkPTwcIw12uFBaoBq1P
ePLIXNxZ1OQXFlflHFXpVghy6UaXyS8WkMNKZSWohK1SeYZU8HvAxy4QoHi4gCfx
RiptOXlzUQGTW36HPjHEMAfA27Pe5Qb2fNdsk9tgI+7twk3F68D/kdmm6fXlzKNZ
h3+952RvkW45uC3ruCh5t2vsUThkVBzR9CULiJKgFFAsvb/zxPfK/yz0SNkGE18c
azifeJOGmOwoq39eDtN/oc/qBu4GI9d78+b+QTOBcS8Tr8YapNirnesV3yomURwF
Ipw8WvKKIfgG6XuiJsvOHPT2NqQIXU41kUxxpZBzFMDNa9SwUguzqSp/3WrV1WZW
kOYBPlLe8N2CRi1t5WCQrTA+1p4DqSZiGQwhReKwaZjAdt10Lh52yAsgP9RfSDKx
FNg+Hmh4oXAJO781SMjO1QrZa3tOtQxy+LHekiccbsBhBTUMXXmlBb84azr7tYd3
gEOQumDfDnVSG2QwYYql2NZrSZrzh2IC/wpegpIJo3F2M4V545KTj8OfQD8ucALt
TLwCWR6XslLd0vio3FUWB0MAlLd2ImEUt/XlLqLWRsYY9MnOXNetyXAUhFz/J9Uz
mgmkkzISTRNmwkXxxN/jjR3/7CXX5IpxnU3umqxWM8JdH0jrR9KaL7Eomhoyjc73
jNv80UOklWZ4RRIAbymwO/bvHxuZ89S0KubyrAfEA7sCorB6nliA8LIIZUa6q9u1
sBkKc3ZrBA0cxDEZWKFdZqXaPR/sQLQTPG/n8XNiCcldh7l7k8ySlRQ4DcE8iht8
somlf1iin3LXwgrfPoEU7ZXw8ZQURLUs50OT6jD8STWILrRTFKfNnRNPyNcWM5Cp
y2CR99ElrM0ZXnkxp4mhbQpdVItRjTG/7AvSjqJBtCxjEgJVsZJtGp6c9Dzx1BFv
5Oxc7u+xO3fhYvgyiIymzNGQfztEl619qMeYl0XzRUjtD4Yr01Ut6QiUmWuOS0nf
mZfcKTj++X6iceB+qxQ2rdfMMwCZ5vj69//YsCZINRlhCjkRJxnAy+TUcurwd9Ut
iwVqPDlyl06GNOjXRan8CRhUlLecv3EU1URy02Fx4cWddd1lsQTJNy3WIYy3i7U8
DEeWvCCFJqkBPdb1jNnJJFzfNKBngo9XmZ0+s6Ts7BzUsRgasACkfirHf9hxxMWZ
ZnNkWfkN13k+Ik6ejm1yhBME+gI0AUAOgSuC5r7NFs3aI10hb5A5WNPzOjyqMYLR
y7ulvtRkiOZ4sclVduo13UFwtP5awFl3R+AORVV48XwgeKFjs421xzRHm+ndK5lP
LegDg/TURtIog3JKRkZ0+XigXxk/TFlK6tG2xynUcZROdQEh5MvZT6+DHQwfywc+
9pgPyo91GKr/ZZvA5c6lo+dTK5aTTWGGb9kcrUWfRETs+1lfBcBq2QqvGqgt0kxU
b5MQ9wHar38b1tQAdbFrWa/jtdAF1pUgbpjfHfK+sLf9yqSdHoZNDfu/ZJQEtzIA
nTC7xDBnc8CsrTI2DLxsEpcIOzbHF4438XL/kyn1997UR6tqIcL5A2wbbm4DATqo
tlMZHxskWoOjm0nacpcLuuFT6kaAoi88WdV18PeEsXeOHzwQlzPdKofAsyrgQi5/
DRDfZbl1PBZNkyRD+snOBmd+7a8hrKAsOlSuXsBKRV0JiwuIcU0bqqZ+FdV/2qc3
rEDSV0hqkr/kYoj72VsN2tt1aaFPV2ZJNzZ+Jh0KK+z9e+PyQp2Xx4BGSLy+kOcz
+4rgBVRDeTdynjoB8oSajLprnrqs/wQD7XUWZvUzz+ZOhuKni7vdkzEHDQtC4Bjo
iO+32zbsUz8ZunQbcJrSqvqIB/Izu2MCeFZODWVk+Udhpo+Ysem+pQQQfAmQgrVG
7qVxRa3MBURyPKnUMgi20ArndHGjr1K7eY5uSJZokJYef4zIFYd/Ze6jwI/AAvBV
hFHVwv+q1ZPPhqWvfvPQlhqpCppdLEX1V1EXIJLZPnqJSvauRBCrb2NXj0E81u9n
UFUVACZj2l5/gDnR/ZaVovsuyxZrwLI2HewB7Wa6R0mc829lrMn1H2fH4HXJw/b6
FvpaaqxjHZOLAUnOFyVkrbMfOQVYyPZLaKNZnGTAEahFbL8tOvdzBRn/hfUxL5qp
B/OcXe7oJ+S6YmMR3hlojtYI94sN2RpcqHWmNW9cbtojQ9uSnRaPAWg3/FNdNvzm
A/YgjDq6vaAPETOFZ/kSLwdrD5UYO8Y5dd/fHAwPrLWaosIpaPxUo4rqbZ1uAohF
Vja8F8aG7bO2/ubcX5jz/dn+FxNu5Y3SQo1VJO/UV4pC55Wb/ueByioN3KC5v9gq
Ka9p2jG5okV6FJ2s7CvvNOSdsRKwd+XehqYkOImFi/qvEZ+C/YuczxeEsOjleogL
yMRvvMohO/UbLUlY/1Eu6X29iQccl9fvHuyCCbLDolCEIRF/GTwUuDVIFY/7Fnwd
Ux4UAYdYKsQI5bDOUk2sD72X10JLZeXAGVmbnDb4h2EPXMst27jhHMd2BdaVBph+
BF8Iefu3Gh2wOPAdk4xM74tZ7gG+LBVqkOfLG01Fc5BHmie7NpxBaKGbii4uifAb
FNOrVecdqMzy7v28EF30wuyPsDUh6Mwt7FSYfix+fkHEIEcCpxHJ9YwFRRJoTIA9
DJ4UFf9N1NQeFw+3a3OX2xREZGe16uwZgkS1fDK4q77yxGrqLCRruM00L2rYvD6Z
PLiylPTAH9QIKYz86vudXfdM8WUaPIQmrTusKMu7owsIvHokojszg9z/shitgj4N
zrNdmoah0Z++YZi3orizwNa1ePr5GVPg+UJNiM8ucDQPky6/yRe564aRxLqRnjwb
Mi/VgTYGdtmGtR2JhniT+7GTYu3qiL/qgp9adrFy9TGR93N01oQlawal110nXe4c
kaluB3jzyR21LRglibS5posLhAScsFrCPx6OEDHW2dxirZsS/uP0VU/zLMxQgAbZ
2UwR/N6bEpI1GXP4LNZilZQi32FxBimCfrFZud13byNona1XI//5/ZuTV4WXDFYD
cc4uLPHXHC7C0Sm+BchOaFJavMEJ5PJ4jXqkYgPbP69ac8FDZP8XZLKso4jOoPTf
BWeortTHiVFdUXVSafxlZqmxrlY55c9pV8CixeUswUfaeJieeJn+CBKq686WOk82
e9nyUJK/fwD7u87M1Xu4O4cPMdmnHBzxOQcY28CRkUA1RKmX+p8AOMf6w2fJzW2b
7ROagRV7eCfb/RYwn8kanr373/7/rcDwXlMT0g/WdkJa2OBD2VnpbMVI0V2qtEb8
O+YZDvqxBH9l5NxTOAaKTFb/KJ+YPt08O4Mvl2NYKe1nB4HoLj5ztiMe8G6cvaHA
M05bSftNCsCdWh7S1Mo0+EEzes3wcKxFR5ySfY9XOJrIaCCGTIqwksqNVg4zFbzr
gqk1Bb1/+OnwB7p41pJ1mIjAZGEc9OT6dCE+lCP6SwfAEW4trDEMHac93g923d0v
xB+eSvn2pgYVG6R2c87FFmS9isy41oJ+M1CBqStLUrQL4HJMoscYhdLDhDg03aqS
6b97cnrZgTL+oPAwrrUh8W7oHciH9DJoTpR1cmAKaGDZq7jSMVHly3uSmbY71zuw
XLsEE4AD61zSUw1MiJic4nrH2jZBT4zBe2D2nLLsSWhLa+b0aF28ZUKgsZwcZN+b
tFxb6y4w+VZLk1sx+1QaRruhmQXBlY1XnXSPCqeGpnLkYZpz1QaJbfM2wgak/vHj
chs8ciTAS8ULNlfzav2G/ftd44ucO1ICs9hByYQXUH9Y+R+8tveVHkq31g8Knp73
Oo27hk3yqYnsfMPwKaerAHFjSuVBZA60/T4LM6ocgxZD8o2c6/IHsK6xTb8OgU43
UkywHrO1yX7AZc3f6JL5kjLulXoo5DI5wKYrDjzrYY4UaAX+JxXfGVj3/8rXxfRX
gXaFgm0Kwk29aO6uQBTZ6T/D7dxWJtg+rTzUWH7GIT8F44FDw5UV35i7T+Za+uDC
goH/pyAW1ZCG18eRhxH+iT72cove8Ah+tnNKbj8Er/n4sRlpBWkVwMBVqY6EO98Z
jrl+KiNWcRgD5A8e/OIzT+1hTkE8ph375aquasKNAABurlEcZifS3+99d32fm7w/
Vx4Tjuw6uph/fePBdxLObIyeqIeYepc2AYaQu/HZYInRDVEiY2jin/NI8Ip9JrJO
38VaIMkuC/n/41CtB25bNRumXU3ZLUQNA1wLP42PuSLgIU3dg3W51lc2vUComBTO
gR/kZ8j7PNT0ghWIa+cY7vVAcwr9LxMJ8posud6rq2uru9rXP30tgC1pJY0gljAA
wIrz9AhMulmmebfvuyno+slK2h2HKsujRGa9piZtxAScPzeKcBTeqEyacTvJ/m3/
d0BLWcwyn8dq5I7v2hnV3tORy36PfKmfvE+PllkhLn/g9Uq/LcY5B4goO9mAS5ZQ
cox89j40a+6KjbiNUABA6H1ms2+VWA9V7pdq8nPwAd2q18aJwFORlpq1VMLPXrfI
esdO0O15/Z3/ElnK5OoIA5L0E2brJrRv/rT7geOxM4tBDZW8LzVs6GWqN7xETqDl
4QOjM751u7/6QAstwGaApPqvNtH5BxAaGFbeIJEq5cq6PhSI7q9zR93sjW37d2o2
KLkgKxr/cZxdKEAovY3/GBF7N7IpGjxRoF3y+amgm4YzqlWcA+LITlVFm/kOTu82
Gf2ekAK7APcCtlJR12sFU7Wk99VXIB/HSMZ1Tj58o9BT+00C0W2XEUVPLfErtyiB
X1aaEYCEtbibFXevCkfscP7WY7JwKHw2XwnUZADhT7eakgHcOehIvxx/eoBa575h
dwq/ItaSpqut5/roV5z0lF0WG9YfB3P8KmzYeRFmTvM3TF28oQZcvFTA7SGNW/1o
pfR9xEgJ7wMgo3ncj780j9Xw73RBRirxOQvjR0xXe8OjTu3ssppHz9HNTZbXOQND
utj0npvDjjOtOl5/YFYPF2N8pCkH/qZJbdjR24HtJX+BtrdOMaMNq5ow/pzRtIKj
TLxDS45PjoWQHKSapCJ2eYS4mgAxc26STaCQKrm0hgupmhuL5wQ69wya17Gl65Pf
gYdCn73YgnisP7CBHVC8xX6y5kVxoBfHJSugBiYVpG6z0YPm38IS6j+YytoKup5y
EU83j+kawQkfApEAX9rzfmmUb3cENgVqDvh4zG4NPRg7MGg+9YiaWwLfBNfuRUSF
28Rfbkgj4yHyEIbglkF3Jbcowcx+j2qg0unjSEHLbopn9LA4l1Ui5+r2LKzCGPEB
02whttWwg35zMYw48SJdPEomaFHzOCZ2esfAKXpK6ZGnu/+rHHC14ADlEINBNjqP
Rt5J4+nGtIT3pvEOC1WM/e4C4xuTKEgqG3XhJRazu4ayzOuD34w/jOS1JLG95c1H
RB9OQVm9VyvkThNEsLHGiqPMpFlJiaTLSJX5vFpEF3/cH9+f+ATLQb363FlJHGM/
heoksVaZivfoayD7bPKhUKEtla+0YRHR47rJ/fVryY5NvRh2RCnc4aFXl6hUfbQt
9lWRQxwfUrDE7W43B4yeRZkNCvELl/FDmqNWjpcx3uNZ6uEBh04uIpjwC9jlBvE3
TMJbqigdG/ZGCjtKyzHGs59ayEg68k/6jJZCpKo0/yQdZ+C+TGwyM89O8KNQiSXe
Gph0w0YyIn/a2Suy80U2sVINOB1MwbTbSdw85dz184FtxYncm02UyVOPBVgRLb7E
1eigGq9bI9I532sgy3FQyuCnyquucDu+R1MF+uyi4ZFECjIF1Kk8R4cTOafsG0bL
iCP0SOVR2V5c6v54BPfKjMry9Deja16oWPunOaf+9R1YSR5jnwc4Vvb1dbrW89rK
ls4c+ma583HEDtBnFL6+Q/Pt7XXkozTDcOhpnJUoq6B1aMNHPQLk9VtX6Me0OYiu
Woxjab1A7JOfPT8HxF2i9fa1xKeqosANDHeNvc9j0GjuKiXqmjJLFv2rNadBhWE3
4Kep+iZ8aXolTsr3LqaNbjRF5Jl+knSO4ufU6DnWwE1Pt14nFZteuu80B2DEFHqg
NTtlJ+UO3zmrPGya/xGgYCvaJL7kd54YAdphH356c3sYutafsTpRWIu7/zkD49tu
Ol51n6RGVDKHX2LMx5yy5AsbxWYrBg6aZnn14fyJmu2iO/Hj9QJ/siGE78UCavUO
rXgwb4hpXHPrvIKK+un45jgsilTZvU07E3IdegGTXIOovM6i9R/N9WySu1bJ0xha
4bkkVVuyBG/84K3zXIPS4/x/SWtYNtAjZZ+qCN+xOsf/S+9QwK2UykPpgYNerEQe
60Xcv24BFnS0NV57rMYIB50o6Pq3iymb93a+/adeyzX40nvnLnK2kHZctItWSo8x
CjdWyqJk39pf1Qn9wlY8z7mhvBZIm9b4F8zsuasI97icgwBWgiEMmEMQulpz9pH/
+pZqKvvDVsxNZa59P7eI/3DL8yht6bKMaR838kwsNk++Cs8W9Dd3xg/IhZgjFxc8
uIPfRPHgDdybSCAAFrhhqYyO34olcjdO9mxLc9LF50MX3MCapWjd2RNltIjs+1fE
6CvEL2h3gIVA8Fj8b0wPsr6OOXSg16R+2V1OkW0TsTS7yepwhHINyirCogsp1oIz
wRgOWtCpot5g6LbUf17etDLGmUYuuljuHtz5UXDDO01e/0cVS3uufW3XbQbzetsL
a9A17X9H/wa+Wz3RvD2Pns5rwKAoaSUB84jvtIPvhdMyz/euGqSd+9B8YeCcpkXS
m71dl5V12aJgCtqwRHahJMwQWAs5k+pBN1oxmAuQHKTqS1/+BxiWnY6ePA1JkFQm
UTfP12RFKcFekKEHPcXjJmvkjRFadJKn5ZwgD0rgGjtOIjYgyn40e1Oxr+r0Xgsi
axSVBtyEbHBIADgpIsyt0mwM/K44gmmTQzrLDGBUkCw9pYSwQ0rzdbJxMdrpxq0Y
6JI8/EDpFeQcsrEFXikC85ahniSkt28Mfro7eqSK1vcAoTvs5aqgzXff6TR57MUT
YEm0A4Jk5+lMK7YJQ7kLOHhP7IlvRf/h9gzZBK3mUlEAgsbD3amvb+idvZVIM6jA
C89jTKfBkh3/lWZUKetETXqtJWvhPgQ2Jg8d4I9b8CsgufcV8SXO3kydos5BU4UT
25RQ4GtbqOZrJEPIJisfNSCmMWSDItNxaWrvq/65J+Ht+DTCp8nAKrECamLYzc6k
0qHF8j8e3P//SB0FL/idEL8DOkIro4C9YzFe2j7pwR63rvGDDFa3N/AaSMv5wklW
pp6B0APIiZiwLVDxAkACzeQ8yg4GE5JC1VQgnUj6e12JLm285L/c4LNQ0+rDq3p5
yImkhuskhtK6s7scSsBE5sadrhAAWsJy0acqs3LMzH630x4K240AwZhrUw8vaQH/
+DVSPzshQxVllpNf6mcwh6DaRFEz+b8nE+CtlrJl1ME69QHJNBABtXW7vY/zzsJo
qmf0+iSSONw2HnBpELvCz2ZwQZrCjMMvtPfE6be9rlWlg9HTQwkzbJM2oygg9i0H
LH4y8VhG618oh++r54Yttsq7SYXr/xCEe4omCBLYJDGqZnhzHkt64LOQ5GVMuViD
7E2jRj3kglQ0wiDlEDd/NGMbojnf2gXfVn9KdQIjovKbxNQJ3zbms/lrGZNdugoq
K0HfaascTmRxRgoO/WbA7YMmfOB0qFj07gQPAV3RZcruxjcHwRForH4DYrWYnVbH
HmtcOjRIf01Bf/UDNCw4TEfEqcci85a+S/LVmXtKpaS+57venk+U7D2cFLOORFoT
bsFmA6OXQr37ZIX7Umk1bORdTr7d1oEMN0/zOw427xYXpc38q0hBxYzULlinqdPH
vzchYWe08HLov5nskt9+kp4jMYXrR59So6t0gFDKKJayAvRlcgYeQkOi3Ju/cmFD
niF95bDKNFH3xc5rNmujhDSB/q69vFGf+LWiOXOLf2v2u4iFWDzeC/IKW4VV/89O
8cv1ahdpJFA91ta6mocczCKmrnPiTkbI//t0lL7e6AqvkKv0sygsx6giw+iWKdXY
WBCpSNzS+7vzWy7eUEm/0S3ohkDdKTqMwCzKM0i5lhQJ2dZ1cV75k2/4J51tRJP+
qc3YCLnVIaNiodMYML99FNAr3W52ELqKoO68WGeJ86YBgkRe1zPZScWQDartwUd7
i1P9VqL4lRyuC/NFiB+OVpanJjvHhVYcoqXuiB9YhcwV1Oc63aMUcC1oMa+8etFa
IwMJe4uxHV8Sq8hqEfGDL67F8qNMU+1o12ZwSW1URW4fhzsKjIM01voJMlGu6KzS
G0wzzs+04rjKUlX9D/KHoPE73F8CJMPblRpLbuQ0BIVSIKilp0bHL5RFooyzjRTz
SbfUU2pLeZmi2+sR6/kmpJ49BuYS4c3+3mdaKGOfr/S4R84FUmRCB3gsxcXVMe2c
9Y8kW/rlvNFgq37rvY+evJ4UPVFPFAVS9Hse20QQl/nz4dg36LA84yz+F1a9Lc6b
Y1sGOK2lV246dQAmcmVAT3pC4fXDmvbFnt49ELzEGjGk54vIwJj+q5PtcTGDD5Ke
h0g13QkL5YVnQV3y9nfLuv7tn0TNJQM2DMoOU1S/wbq1ioU4YhjiT55NXaXF9vOV
CgM5y7ULEWwRRuAqt88fLfAE4UabQ528wLt0ahXwUvlCEys92HJ5wNsn4ca/khLA
YmJPpbGjkI/mYzsIajZGwJ49aO2J/Y12kNLrjbh3pID8HZhxqzHvvgqbLpe39yNj
qgEy7BsH9QdWgcjRhXPIBr2Nyhaw7USq9gKTVSK0bqeOEwnJ2RlVLKAgh+PAi7hj
3bRMM3Pi61RIwnXCpFQlovHNFkauUVJyBkSVBzAv0nm5NcEfCBLiFgnJmUfIOv5b
UzhN1ay/pkkp2+P52Xn9lL+ocjXk1wXQiYZoTOhTGVLqHBXsp3m/YL6eblPp3Mr3
73QQ79i4NCiged8uxIFzB2PzJhMi2xvCIRpgVcGsW2DyhgQG+Mkg/C9LAGUDh0ZY
HbU/lSeHaLfMK1vSD4Ln6nDoHcbHvxP7LyYNgQ+r2fg2wpUOKO4oL2QVm4xBql0x
3LC6WIgtfUOyH2OmkhilKku1JcP2wuzNSJg9BaxhmIPWCdQsriy4ZX0IrvKB4qNB
gKs37M2feF2uNlbuha0E/tNdS0+aez54mtjE4CrgBUk5A7/CTH/w1NllQhKIEbfj
JTf0v4/4E4oeFnpXO+YB7WoksdF+vGGMwFHyoPu7Nk9GDeff2raJRr0y9qH9ytaN
FCw+u5SF7l1Z0aVCxQtPZqi/6/Y+Uu2dG/C++8qWXMxWyfPflhPEH3x3sfJWIZam
ya0rLuwPGyw16ZzSWrThbegTqqGBro0rA2BQs3rVwfuacSr8L45TYVjSGzoNQ/a8
8TLXtTp5jFgfJrelWq33QlVSynDfMtXdNwqk5BZYu3JO8H6KqIG256MCv0lFuh5Y
YQfQzJvYe3DWODym9g3Xc8Eik5Dq0C7FyS5TXmB6AMRhrTMMpUzLZ2WH9BzlOw0E
7F98lP4Vj6PmW5W9sOW56xEKdxFQRK8EcaD5i3AeLvgr12G+n25YoutNyKklY/+a
1f1GXio0TRXQxINJ5OXuEgVgpuyz8gpUVzQYjkq1LPL3SqCXCDwW/PgYUBzJ69F8
9P2nyUSgAT4GNYFKCODz8z1ez9v1g/Pth0YANh7Enb1TmjvibdjgLCwUE1l3Ya0M
VHuEVTo+1aCVD7gzVTrwVwVjK5g4AdBNWKSqq+qZ6ND9ih7vdjSLayZjVcvEHMBg
zZRQkOYV8DYDNUfe9uQ8SCYze8atfq2UI63pTg0U087gfVPc/03Cx6YOVakuFe2O
A++w9w53I3NU8NYJwDImSSsUp8m2SKP/gmOKokVTOcNl4oP4UeJVIC7nqlGDzwaB
1NX9EVTnDCrbVQE3PneZUYCmw5hykKzsZ+YDgqqzKnLt2b/peAjahelsdIBZWgtR
32vqyEOb6uOGk9j6aSnpPFuT8eUIFi03W39/l94hzz0Ab/5ass/r9TWFo4V0DCCx
/hARkCie44mw+T+j0/12Wxw7xo5Ka6g0vSQ9ygO4zAokGxOL6E+q6yGLZEsIyBn2
1EmuW14X9M+WfZwaKr1hzezdB92ugqywrAuJA1IhnLxfcSa/fBdOMkCtdp+S5ZeJ
U+nYIHjWMKzbgdLYeCqEZXnRonZH5y2dv/YaYSdfYGtTZLFDBqKn3ZgUYjlwXMXf
hS2VO8kV7ahlXow1lgRI3wjNaqd+K/wbXCCpmX8dThR/l/ddmF4375FdzEMb406v
pCRhOoBea8WD+DSZga2VgeMUyT/ZXBYW9QPjFwaPZP8qR+wKpAOz1PJ8i3Rwz+B/
FuPLWJH6Y79W+pHSgt3uV/UQ5YeVNlvKYWw7pqWYjqbwzvW9KAQRxti/Cdjnvsjj
ThDtq7ZzzQOERWnWbuF5V09dnTPhTR2nR+BqQqIxITfWg4HphAewNHSANazpKPXu
7KJDis4iopqQgNzCnOcbNPumeF3OV0eA0ITa8cPTb2BOy+8TkY/vZQDBuLVTdKQW
7mhix1D2sXQ3E04cAAOeqfEsElIcciFMSfyS9L3E+8KTthi8hHlmhKtuWSlXeqrI
5zF5iKoUvWAE4KVDDSSA64CteEdFW1CKapJFwYPxV3+9f7ivcyQoKiQM7Q1KGUwZ
LDysNLt0/iWYKjzRhx/0OWmSTR0H6DXbbA5lag1dECcvwGFvI9vcqeGrVr7ZT1HD
ebutDeHg9w81vG1JPK2R7XlR21XAYmPTZFKK7JypBz2mGAKIkUXKPBdbGrV8Mk/6
qZx7S9TRAYidi7TrceuAzj/moMIbuYPwjs/auDMIePuRgbyD9nREn+Yd/J3ZnU8t
u7kqsKK/xHMSnrgOUOB+ZpB8fEVK7E1Q0nuFqxsWCfoT1mXCa5PzoUVHhoA1gzRr
fe+pHcUol3XvlEdz/erpj9xujuIbYKSrBesBSqi20+Gal1/zmXZW8DYY0+Dl24P0
L99bGjy7X0YEQhZHDnBIBEGElHxblVnzm5gvnppxXvpZG65kmg/f+xT/trKqy+qa
0bJZMVAS0ofzelGWayFK54q2ZddPokRCtwonif3Yw3/fPlA1bKjI6wkSApzDBezG
zFijb5Z7IAbATjNcl60CIkcFfsBbvEKOYv7+ldciYp1Fp31QnqMPIa9zReBfb51G
Loe/tY1ZdunjMaGbT9+UGG5CmxVFYV0FLChhk+1XMfH9RJqPIlPONJbIVGj9oLYG
xNgCzPh0X0PgAgsoEIGhg0EqWZLWsTxY/5utHqCJL/A2ZucSKOojVszyR5MLFjxr
VUHIY4qGE7BKQAaKXR1+xq4x1DujEkDZeNg+IQXr4RJ0Dh4KYS4VoglUTNegGZ4e
9kcVvgDMgNRX6HBiNkajJuECq/Jw6cc2Uho7dQKo9MEEL8ZvAxkQcG7j+ANBeHYA
VCvfIDICREYl7naVASPh4mTh9S7xiVeRL20YxqFBGAzX9oYXNY9JO/MoIpo0LIcs
v053Y5pVM6v6yJwApIm0t3pEoz26v1CzUr7CLV/fK2RsBtrwBMq9OCBT40zAqQFt
tr2y6FyTkGd9fsCRoBi0eqD2jRukJXGBaQUwK8eNZSqMIYnHZrp6OAuNou/snm6V
iUcn5NApyH8Jdy7ZGAgMw3pHzFpaC4Y1Ijib2nBTVWx23hqokAdWHERY1d6ihDWE
57Osa8mcdduHZm1lxg3osIssQRVYMGAoerstAQ72nIyu2pPfplO6iFiVz9TmL7/+
hp54U8FuV8PelGFASzynEUK/6rKow24ayr6tyL7DB2n5EPdPghYqgU1l+q3d1/ZE
By1N+xWHpTvxYP6FapOcNC+sCuIquhLA6ObyGDu9Q+Tk1x4yGPJjG9V3bOd/NrZg
17TayN+U3BB8UKHppI5kDP1oWxxz7eAp4TEbpE8oL+IZ0++FKT3PkXZhdJ/NZlW4
d/ZxUwXp2qYBZRnMPOHXFE9MFcDC1gqyFWR273TAdeoXPcA0nI5OOotXAv3Sejof
CM6nsMeTGR2vk2LXSg5A9IVVxANxQzFsJOZdF+sQvlzuhbb0bmEYLu9keac2YMzs
1QhJXqI1NyrJEBC3WnynE99AXFhotNJJkuSBg9phOOTAlLzvdoDp+X93jh7IePIZ
ZPH9Dm7jB9LNOiSfkkOC4tDzE2krkXFp4oYFHRySBtGmjUT8fiAA+J/DQmjpl9SI
BohZYEbJ4MVgx9rwg9Rn9naswt/oO72iCUZtxewfvYLweqkm+YQQ3/h4nQC2J/eG
92QtgxQ9HtQ2AIR4RjbSuo4pq6wmAkZzzA3LbmhZjQV83eIGf5GrcmWc+ACZjMvh
r4E7WYlSAB2y8ZUXfjs2xOMGGgXLLnTD1Cd4QjbrtWrdadsujs8Dhqw2qIvaqCyE
mlPjPrqL7cNdU+oHdNqOVc/qKeMUDhXg3ZdeIh0ACa6aG4+20W7sIW5HNkcggTA9
dvx8wmVRgFTuXTzU9CtY4KVdQpVGcHcfAxpybM0l1UCRw54eFHqVWzjjpKm4SfYT
cgi5OgyJUDL+vV2s1wgdIM1SsyLDtnJ228oxDxBDD8F1e2vMW9fH4tGtKrCmnhyJ
NZC02owS4Mg0RdABkH1/rxILanUdjGBu3EF8cb+TVtOjMrLdMIFT5XQvxQzEpZqJ
/cSAHY0/UyhGXbSoQnWo9YDidNPZpzJLVrodG7fZHWAcb9QXhkB5d1dM6a/dBn6L
aXWFfLQDgDPXGPtoZ56ZOEpUT1+GpbaahwC40WN4CxlE/Hiy3VaPpFjK2mhpXRmV
fZgdcY/5HaodmYfflOwjIsc13dEHCOxgLPm0aFTUb2YDtq4BSxvvVFlAHyj/1Omh
mtQrcH1gTWY668AgyD2MkzAu6zxmPgt46HX79HL/IaR2qRRVjoltm7kn9AbcVmjq
cgPeZhNzHrnIVAA+g8VN30uL/j5qJBKDi6U/OqI5LVs/ENeixwgfZNKVac34nWAM
LQ80r0qJQm2BeqgSaVX5Va+sJw7lbMUQV/csRq5RjLOWcycCQsrUA5hh3L/buP5b
FqwtupTBN2nfQ6X/BwYcrl+95oPRdkai2ubAWEGthCWbewfPSUxaQqzWB/6Ye5XB
tXC0xxqusa5LD2LIcl0QGsXBzpfm1sArwxoPc7CpiLWKD0IXoGGfBXNV1EDeuUdf
M/bHe/8H9EFbGxpriPLQZXfjCRoFwGAj3YbGR9TmqNeSq0LxMgcbQEvHfTUR5XRE
bdATViDW1lbkNkAFwl0ldUhpFtxUew9Pyqj/ylI+EYl9MRyy8Oo5SIW4bksRtKH3
V6FCcTEYJz+FNYl1TijjvjS2CyEc73sV7oEfVfWa/IWfR/tI3Z8EeZwKLhEo5SAg
qsVfSMkwLGv8JqfsMNVXG3vgKcrAWngBTrtB/r2wGJrRTYUYzseBBOMVv5ORrH42
fy48VC7a6X8xi9kH2da4fHObbwyeeKqutpjthJXRdXgt3s16RRva0SlYg5rxynVS
fPY/48FSEwZSNfdiU4hN2KTO4l0D6JOaM3FH3KkEgucdSe1UNN2CHRpfzSQN5a7y
Ih3aHFGLcHLQ/KiwEXto5ZqbDJynx3mWvOmV9Y1NmePly+7kdi3zih1wS83e3hXO
xkmIiPaa2ZbMl5omp0LsZ3O0hVUv/FGgfBnwO0a9y4b3e2cHo0l3RZfV7BkAlh3l
DXbzL3E+OmHDqiJK70924gseTjTZNgBGSlSqB28UmYNWokqQnRZC0CYw53LCpQYr
PxRoleXf2e4DlAX9W+QwAKpnHO3xewz0qMffdaNI7dOhaZMdbwCLFXqRhcsFld+2
G8BB0lBHnpUCKhKs9Xb0KTmn6poOJ5W/ZkJFseG5KoeP3VhPS678IJY4Q70t9vV/
PthMuQxascFufC1FYUwAGQKg6IsON1kbhy/Xf7MYMjKh8mH2E7QPl9XiLs79ml0J
mlnyYz28o4VoQnAp9Ih4DoAlr3wzkyHxq9KPiXedA2PYmonD/GjlRxnAz7Z1ntdj
Jm9y9wz0FOTy2NEFEUYXm7bP2eG536Zw3T0JIIZBEVcFMIveDQUUDX4OtAvFCM+Q
NZPpteH1mbRKAzVL2fEi8xxBTDlQ3iEtaNNUPy8qcA9VqeQqQQdc9p88QAVZdn/+
WPNmPMQgrAFOx2BKSHCijbkgyLRUMcEzAlU0Um8naKv1I7q/zf4luR6uni9wchp5
VQlQ2/W5MbtlNuZOzAE8cTY3g6Pp2fVnVqDmka7rPWU3ybS1Tu7bhnWD3hKYTVSU
GgKw5pfSwUPIoG5U5idvumHW9WJRMHlcS9PpKBpENeYTxXb9IUH6cEf8/mgj2Ws3
c0SPdGxZX89diTNQTymYBrkk71+yQ00Rs43Oq8YzB3+QfmsR4SP4EwgyT/mWAwoK
ojnarWTjfSVOUl1jDxJcy5CudYuf+i3Uy10zGMvFcFo0aIMAOUc9fG5fbecS/TDp
edUuvG3AllNWh8v21Wg2MCSErNBiNao1u+F4VO5S6mI5r5e6jijxpu83AQAWkNzm
DcX4rCyVdYejO0+fKHWc6b9lYwXjP2H3nxv2j72MjLzeLZBEEYw7b+hW5tRwYkU4
Dx4k1LvW9CiGuRctcDI1iyaED89SYAxbCwxwV7X0nwA4tXqcmV9MP6qqr2NXwd5g
juFZ0ETdwc2Rkp5ISWGpQfTRfWF0snhpZXOrBk+3hWAa+bTDW9bIs8U1q9sF2Pmv
w0lvB1ZVl2oPEa8W2wdpL644hRihMF6Pj+85xAl1UG0B6uvKb/GgBshQyXINltV9
Fg0f8hBvxVXJRoWT3YAovUB+DNCPsH8PP9W9FDtreObkVndmhNyy3xByy/fcqkXf
sZWc1iqT9Wr1R2pho8pS8t/mUouyDGnYJGVBFAohsBa1VqHTID/rQB82TAG36VVC
zvEvNL0/p3RH+48nzXJ6fakCzfRLNZvedMYMA9sW3u+BD1bIc0/vmtMaTiHX8Q+A
Qs+w7qi69wv9R/pm8nb56mN2+JXjfMBizyIpSd4N7s68m9dLTITlLdftvCl6dtQl
bcYAR2BEa7gD5oMu4WbjlX6XBLnDY77sZZHv28aB7y12iwX7hLEjGPP0goFcig3b
XATGFXvFtVvlwx4woTcmhemkYqPlw7TY/dPGkAzesic/Bc/OVRssAqYa/rUkXcHi
Jg2kEN8XzuzAwmJwhaQjbk2akRQNDEpHhR6X4IoA9dKY2N0yGZUgCxU3/yGl6LQt
WPRLbebCfIpGvXdVunL7Agb+qClWkodAN8dtVrxAf3dsYxRWTy6zC8urfWPy/iEF
wo9kItjZs6Mt6KWP1Eq0YdmCyfV0Yvv7RdTTBZvLo+pnrhQOjo1imAbP9X2xHuQT
Pb+CXMGnn+/quA03uZTLU3WBSxQq+SXERafsn9y5Jrvz0V2yyaz/HoIivqvf7wxP
ztSX3xW1A7RFXbwmvZz9E1YeZPnQOR3taDa4uf6tlpm1KoohhGEtZ1uhrz6q2AP9
8z3JV5qMmDC4mKAKbZnCwHk4MpZWqSxExz8pqrHJcIj9f49Y40DILok2T1SspT/G
dTtD5e6jRGr4Mjx9puGOzdl1PViCV28gT0GAbvpQPzadVlNxnOE4OJFoUcKjVqNB
HX94rDesLNHfPzip6jBmYuYQO7yZdMKg92570nCq5n15T6i9Im5iI41PmwGImbWl
YMponeNWrLSSxUgHFR+KNb5LgVAnEjpd6UDYc/wZvQ0r6RZBVqVw0cqZuViNyjrQ
S7H5tmxRxofJWhtsb/zVsBADAEoeDsdG8evuzgbnZvgJNhTGWdQy6yXOnme0PgQE
vWq3h6UdTX8lnvWKYs219JYjF3ZvnaGJFU5+Ku7ZktHoGj8UG/IcYE2n83C+yOd5
oGcGsRD5b7E9qyibhqHTJEqmUMudC9ylKmvAAt3rE8XiNeC6FIh/X1yB/qVpwZfh
u+gImDm5UCpMf+F157MsS0QItekWjDXjWvcKBpYMRyKWgI9cIX3vlvwKz7w8ox1k
g+c9csqKHenZrqbnBWOCZEcisVKl+vuNEhQbqufibOzc/srm/4sxaARZXwVoXX2j
AQ7xCcRrTVbz6GxIiKthDW5ejmCaF9nWJEEhx5U50C852Qgl2x8F/uwLKxOU60x4
qxVeLWtn2Eh8/9ialy9YcER5qvE/n1nvTO0cSh4jgZysUYvJqn7K/PpxxDWoEtU5
fDUO4Koeb7Gf7ouSUyL9/xdUaNA/amlAo6V7ItHvl1mHePoPGTnCCsplN+unfcJc
7GleE0zJOnCG7Rc3OlJRoGC2oyqCFqjhlwZy0v8n8UWRiMQLkdNLzJ2JWCJWNJfg
4oIFM1t/+jfmNnxXrqycHG1kYpC2H+WScozl+jKlCNXtEUFRErvxUFQAYgJE5yFa
HXlUi1zQVlWq8Yb1JJEd2meyuJNt+VgTvw2LtwjRVsi5cNJK2Sg4vX/DjCVWsPj4
ZhMx4HfQb+Iu7xTBzlhrI77eJGg0d4xvPl5K9NQyAlt/PuxaynnNIpStftGT97p+
cR2Li4FnFHiTRzstNmkJj0CexOOrNK9z/jv75USPsPmB3iuwFQWOm31lV0Ic+L6q
1orkwBmIu+/FLbpPqu4VeAHncSG/qYI94kpzp5KWG2hAulgSJjpyGIo0LDJcvClI
iDIj60LGznFaqv1d7ZaH5wtGTolLuZ3k52XynDlVlep9GAwhKJ/DfW5Tg/VOcUMc
Vot+jHxAhlf+w3RRMeNnIEaSTrWBdVdwl6SWJQDqJk+PhEtadcJOovHPi6bjGxXB
7kBcjv9PgHCFsXHfVbHxkylJc7hedrFQV+q9l64iiLRBCoIFWPJEJZODtbT882yk
NLyXbScVat0jAJLJ9fuhmkGW4D/5ktKs2M02rL5Y4pRKpco6a1UK6X5wUhqjxtZJ
70//6rTIdxo3OM9QSDKpBoHYiegAih9sFQw7Ec7JJlWxdNQPIRcii3b0J3Tw5Cx7
HE8LVt4Db3VEzcu0Em3CcoB5ZAOMW+jgElcXUMFoyBIU/3+KKW08AwY60ZinzuDT
wL+qaaQRNsRsmmsyE2Sl1QlLhraGJDpY2F3zuwVdggQCYmsJ+c9zV/DQvhiZG97d
+059HRQGg4k45SbZBGXCDnHccpnJ4N3zFh35tGvw4EtgHqo48zfwub4AAvZJP3DI
VMeIEjPeDqbKlx9/rOAqWuf3sWE1xRZE09y4heJjPxmjrGKp9bRc1BI5a7fxx93K
Avj1PsmWke6ZQu+eJGptltpTBsAWLndE+qexshvQQfQQADB/m9jL5FOCJfPIqAUG
80n14PwfXwgFgzi8HsuDDOALNKq+fgTJhlqAORURVbEFjoQatHO2cybW1vqIiS6G
RZWDBmiP9RNC4lDQlh5TiaIBteti84yJLqD1QzgvpJekOP9VtEnlN3sEeL7a9Tm0
jmSVXQwdb2peWzoA5JUQtY6Ns7QI686ybWHoEKX6VV4+z07kjqAll8mgRn4F4jGs
1K5xsyWb3PT7uLPS7jdWgxqf1qGDS2oFTSXXYxmPz/cKruEHFbCuLMuYGDgwOIz6
8fcJ7PxXdWd9NreDx1xE/RUqVFfpC1hnwz+qanF5paBgI7UdNHvVrDk27rQtRxBK
aSsTL9ZbgBLqZJeCwVDduZnm1UGSp3bbPetYeMna451vkLkGPSqDVnonL+Cpj9do
ctW7NtdVHqe/k0r4JvwnBwe0wMlhWAgWAviduQN9q2Nq5f5bGQbbNMOJHuocwtlE
i8LZnllZO60GrVClKXlBE3oaKKahznVYPyfZqfCzEramI8Mus4jirDes3GqUForN
nF6f56GHIQOcXCOeenKouRULplQpDJ+IFyLL9YeUh2nnDOz9pTMyUCe21QY7I4Dg
cgO0gOKP6OcQJCrh61SLIwtdq1vjn9xngUcvujwGv42pn8n1bei4TOaP3Pf/u+W0
cDkuTxUwqNiWUUF2b/ebyaV7i8S85mpeCKTJn0ZGhHQFoJo6+RbKiEK/rK8wRlMu
JnvlHvImndTg3axDYIvs+dD3ACLFMjQaDcgqOfKIyh0canYXJOZpdhC1cA0Lp/Vp
T3VNcmL6Vk5fLCxonDTcgQNTXZuH1mOPMSOIKlStvOhyqsgtSN+OTg2EPMAj2+Pp
qscXTNQkj1zjNEwofxHCrSMablVyNty0eMQf1c8N/JncqpRIieVWVZkQN6adl4gM
0iouyJb4ohfkcl65OewcH1b4I9VxeTXX3x2Mzh2Bz5Kivx2YOQJ52qu/bSYLCNbG
X+RyRY+tSLpH2b/TU/qhRAw4mh4LUDCXvcIyLmF2qtr+wgIeSlONBjDyIs+ka3O7
gAx4f7nl9BVJ9IsEf1EJTBCNyUQFZOFNFBSlVI/ZPDxpnJHjWyjoGnnQrV7AJlvp
i/0So8T1NMkPGPASqMsp9oLIYAO7A1Jc+jZwz2fv1QVyznwrOz7KdKNBBNhig+fU
XoijHEYI6IfPVU+B5UXyhI0iArRdpzWuzBy/lJYG/xXQdMZDSyhc97I6XjO/95rD
o6aRH8V7/M1Ty47aFgc83URvzxk22z51r33pd+qRBAfiIBBWzpR1o1QRNhCuGLNo
OigSegzDqK5bHtTME1OVxCvss4EJEjzOViM7xNvJjt0LVQZxxGJ3C5369zFKGuk5
IWKS8OgdKSzmTJDcBLhupQFTBZ85xhvFMvV3XWhM+8oGDGQ5B/rvqsEU4UKgcMSu
Hb5wOAEPtxolYbk/5BTr0H3aFzttrCX1pbekmeD+90FpE7Dbx5rK1FfQyUOTdxJA
hbqHhIVjbqkr2B8Ae/e2OBWOeHnH1Xft94hJ60cNDkwFBEl3KlyktzVwZavQm8Ap
tbGr7fTucG6+qdZx6Q7Otptm9Nmm815cgXFPMDVpjl3fcAB9TTJJSt/pBnrkYJmm
BMR2dDHprMjKI8J6rciCy7lUoMVx8HJEwD8RdKbEVWd+s/0Hbo5n60siHitSdtWr
Mfx6nP0a2ygU/+1jWJyjct++GBa4RzcZOOVCe9q723mkNrNJoKPwFtKw9iovPXKb
GRHJy6L0zcsj0/2aFVFtr2Avvxc9miLS2vGzSSdEETEVW7sYVSQKmXof9+vUEFJy
QHE+vhkPuv7PbPWks5t7DA6QQLfdtqhZ4xwgH6AbWFQONAcLJhGIC0mXWQ7l1bxY
9MQ1WJLxOBW6ZmaKh2Zt07Q6C+seZpmxt88EAMuLOo+qaIY47Fb7IyIx0rYt64Ud
e8H8VlK6CHma+oRHJsZ8kMP3Ou7d8PbYwkpFia/qsZMBAyHTQaaleDY8NO+uNuiw
mTP4+wFqQM/udU4Iz5NHEEVwTt3bW/Gu7yBEExcaKXJ8u9QgbtbCDoZoy1Ew9yCM
lgb/CokAk7egSOJ6Gcz+IsXlCuR3jQiz4wXzM+8A7Zo3LbwDQmETwlj+f+aHAAHt
Qx1RADcpmUMj3i6OSiqDeM7YH7ob7WBUkX6GOjdOI99tHl3bfR5rlihHHoK7zoNC
kHw47upXkGBObAnwbkiqU1iJNjwznUPRXq4PUoVpyzFAESNIFWEwgufbGyI+JKem
o5Cr8AQ6n32vDClwNDiDrK6r3dnwYx7mJfc1RHewuc2SndZImyQEqRlXWYmE8k8o
eQIkX3Zjm1E1P1NGcoHwgaelnSrE5hwXvl+H8lLs2o3xrtycER/ShEJfKKwule/j
dgBDSPmdmwzyYsSe6haZigCZVhf2Hk1QfV0rguv7RrxBdW+E/yTaj3JnkGnHWPri
MJo78RvGCghsQZaZ7PKU1WOB13DRm827OJyJi5cufgUatOTypWnFYEJI94HJm+wx
GrQoNBJZpuwn/+/8ndj6wKADK6G1I/2RxxG4qncKvcBIDL+g6/PsKd6dJ5gbRxAu
Pbg5fSHSFysbisb4vM0rYOaOIWvVrRGvQrXgxJ809DDtK/kAVmzaZpiN6YZWSpWU
0sWrwereZQp/4glL1JzCbLXN8CMspsiuDFSGdnwqLl2Gfe98Uz2cV0CdaMiwSxh5
vZNCSaeo7nk/asx1iYvLCwpvGdnFu5rOnx5G+SQEUUHLyBA+ygE+5T4PEPzP3x0F
oswf/EvcSVjloUHNkkLPhLiuxcRvoZMgyiulR8iSA94dmPlaFoG9EGkIHgeGvZtj
72WVfiyk/t40E1+TShnzzR1Yl+jye1QaY3UTdh1XcBS4vguTTkDMvOT4MV7V9SoI
JK7/3oTSr/e9MCv4O3gV8KHSUY6vvLuVu88wJe6uNSS7OA2P9cHH1CglxtcIGpW6
0DTUmxtDHD7DoVS98FJs9K9wnII0DCukSgnHBK6RKkOj4M80QydR1RLwE9+bxjqq
yIqvHKAAN4GfTuRzISyAuLvVolGCTlgYFFhEZbbjL9KZJd/IcueRBHHmOqClkEo2
L2RU7SFayntrSAAeliP5rCPvDZpkDx2XrSVvDB6LeCYCxEE7WiAxUdn3HXnnu5Av
AbHgmGgzGcko43Y82YooWDjCIkOekvk9xfyRIimGy+TGlZQmCqMGtkpM3gYu1Vxz
nVenq8dSijSr5cLiJCpoqc1yQ2UPEtHeXPHafgSz3gYEfJJXSFhqOA9ekT9h7y0b
ZgEWJYu8P5V1yi2REl0MPx3ERuzoCwi4xlIWwqa73Ld9RzqdU6zMwjBc5U59xVdG
uJd18ltWCb7LYTnQyhukrkhnqp0yEfe9fKRcDPxFL29yMOtscp66jjN3mIKduBk6
XQYsa5ufBW+yn9IT7lZe6XSl8fvfwchkAWEmbK/tafNZSB/wVGO5QKWud2GWLESX
GzsvRpTZPiAodAN0anvMi4X49UWqKohasi6HkCmZDts948OR2dlgrV+jwrDOjtNt
ukYw9Of+zlPtVr/f6MtBFxLGHNMvurx3kDVXshDBAETdPOi7PPqNgu1OQmtdxvXl
F2mlY4CwKnSJxfgouWPGQEPaP10P3urEV69bG/Su0+ndgDdsbBNYPJob0d5ZpksE
Ks9jxiuXegbCOTO7jnU4/W7r5JZUUkSg5IUTyuNhH9pJxugo9Fj3QWT5z0Zzw6VY
9lXAuebBLsTqvg4QckcVmcaYjQqI9s/3BZqmzK/cyc2fNfEqayVtsyI3emux1OP+
AeXsmdSyH/p61nyzxSyDHtoEAxbInEVhLmqK/EoA//05Lr9tTV0+cVbGKHl06bWT
UG79I6+7L1AYAnsTyQ7Q9qnwNlmRse+H6KiXO6/1waqt8MQAkNFI6Q1kTbXc+rUG
jreh6IofTcvqXIE8eqAgb6Or53bHop/GBy98hcykzNfDZ2OhoXD7HTew7fJmq+Sn
4cUq7Qz7lV1DrP+yNtvVqoo9A6+jY5Or7H3k4S9nf4QfYJVcP9K/eN6tGNWLIyXh
iZk/RobCnFlVg5nErDFzg6rPcI9pArrmw6RYeVsK9IcGllZ3bwmM2eyGvMhXI6O3
j6qDsoxGEu2agSMzKRAYD8r57sV7u6kF8Mke/HVCRrEMe4t5U4TB8HSWfHIJTVEl
SuN0ir8Z4nAUnX7bS29P+RadyYv6z5ije5wDPBKbVLeQsamdS/09tiUC93VFYgkU
M9UkKvXOMAX2tbtfb42PYLRu59r4SoEZ+AXbg70Cx+EzK+Fn+xRCalaFM80UKmLA
+8vfv2zKswMkDwMsTsB8FQ7eR8fdEWxlGR+h42/neuS6dxLpi8p9IMZk/CV8PUEX
IdOCxTZ8GKEKkHhD7HcH13Ga7i2wBXf/CyLrrgD6Rg4v1ZUQ2RdXEA/GNoFpl04H
REGutG060ERSjlELojX8W7wNGHL+QhMpDcB0kQ+lyE0n5FiBA9IqXjX9CmQWjhox
sNhYRApQNhFwwZmspLfxMtrSgm+gmXhPnLU8WN6tgGJTq1GEyukYlJiiTTSz9pGh
I3Gyo//cHT1c5vtaNConLNFkJybiylgP3aZRtjF+ul1AdlNA9dkHPVOEsCBf8/NM
E487YxL8ftmxZr6SxFrd4kRTWaVmYqfMlk3weI3sdy6mW2lyU88hZ5PcpNjzfx4H
dSTy3/IilteTGhxoq/OWy5gg8Pp4qvgmDMg6NzGwrsVUB47FY7JZN49HzRTGNMZl
sj8quVZyYPwXZGfFN/lPnPXM2fbrKnKmBXn9DYd1fUJGhNLRY4/tYuK0r6F4R6Dn
hHQ4y33g1163JMIdlo9nJPfbX1RybaeDoZ4gosl4MnC168QljqIPO7zMuSWYHsov
KiEo6yINxBJhp1djDuKgkF5PVeVyflW88/YcKt6W3ahCISFlJX4SU32ux2dS1Whs
OFl2g35vN6SfNKG2Cg/Cb813lKco0S52rsSxBJHEeQKrFhKfSUofm555rnvPzqVa
iLsuDUm+2Sgcpukrda8tIwLV5vdSDYZQGlchY5f/L6EkPuDARtX2OzFvKaUqzNYS
NKuivvO3jfK9oOFrOC3wYyQGDnfIsVt6C3LPttTvchmRqkEPzLXAHBVv1IepEuYT
vKXsGt373jS+vEwb0ZQd/V3VKh5kzqPcyeWieNDtOpobLtGG5RYwpJM15aP6BehX
XrHTylbitB+34xyekAwXI9AcosusL/DpozxuPNW/E06s6kfdnZuolVpC3O89j7py
pmx4i9ZJJyTjbOQwOEJAkPByGccLqArfdYii4WEGd0aDExtwctv/kI2wFkttztp7
8mO0FSTZ0F2X/GRDtbcBUQSt/zY5lS35zzDf2yzahimk7AGF0s3EzUS/cn7W6cNw
SQJ7P5ZnRjl8JYe9w7UqvauCzH281VZP6TORrfgs7syauAFVCnuuRkrX8kEz8hyN
v2ZYZgLjNViZtjDKqomCIycsYgDr2JBfwCWl7IkzUctxMIQtY/+EN4gQAkCUUhbe
5hRUo0oed5ecgTqt5EAtM8hLX5b/xxJeD1govyXWapTyJeMS4WUIR3z9oYPzFWpl
phuKzeEUMNj7nxp/8owRHhvh757yhD3H9STNK31XoHnXo+iV67W1gCGyKa+lO0eN
ovQyRBwqMOHeHNAb+0gmOy8FBOVGW8kUe7Ohwwui76A9BhRlX8JvpobxlGA9Wp67
JoljOt+ZkfNkdeZHhyCQsilg8xak/5w8llIOXbQZKhyxS7CS+T2OXFHjpBfD3GPd
ozkx70HHUTsHk0/lzYmxLSbM1Ph4y2BqFnySYHvOp1CJHgeKm63/ng1tj1u8bKRg
PA7LLwwvI9Swt1xR9mAGRHBKC/hSCX3lPKVB0v1lk64OWDCio6i8XQcySUlrbtHg
Z0OGzpnZujKPQAlWDHv9oTqitUapTknjLmKLSK8zo2OWgri4+p74wFtE3hWlRT0m
rcIEq8EYp9JONZeJj49JbwyaLirSM+KTQerRPrLVNvZ2CQSFoAnlyi8O4B2Ji2yK
lsvDRh3nK/aknUrp/3ufL3C6pekt3ZLmBv7SG3Rb+i+OmXLkceWKzusEfZ6650tj
Aq875Wrsy2SVNBD5rEZ7RUZ4rhYTVyRvt78GwDKUYCRM5dBO7gU5y5yekHeSmJKJ
kFFVziDfd8CJdVCdtVbQ1iEQz17+bylLeydxLKKX3wkPhIFEYOG+pXMl+9Vcw7M6
dYKqvgVH0MMNmmtRYFenp6UF1tel1ZUBKS29HKIpL2cqPny2GWHUchwFm7zwV5Ni
NIWWtVZsGlpu7fFNgKdXNYluq5oKkexrqK7R4aIPLYVWnfWrjmnb/eJwhv24RCPR
UZ2ULXx9JJ3pbAU3p6Nqw/xz4uJXwxBSXRTcKD5XroYsmfKQeVZdRLNPfU69GIqQ
2x269qd9OwefDDILjyKVrfiApkEZ82+GaTXPdaLE5U7DafG0rgeskKbne/+VV14L
tuE5en8QJsu9H0Enik2/UyZPwBKixfaQe9LmThAbPhoT+IcagXfGKzo7rck0orHe
aXeSvaBnQDpUjBcLgah4kOmnfUDKtJ3WsIhZy3liurcWFed5VVSWD0iMV6IymBJi
aQXCrRTUXn7HRNpj02fmnEKChbem31N040KpqomWT+S6lmou1nwqsL3uUIJ/GYT/
yC2BQB+ytJyXXfXqTo5vljhhrHMOJ7hi6rdH0G5IwwoujshNGNJFy3uqHEPYql2a
HOwYNZM0EW60MitUHjgFJHD91gf+1QmMr913FEK0jYUiXHbvOmwp6MQXg+M/ArLY
keiqLkM3QwN1TsCu5yRTrAGk6GHoD69DJMAxBp+pH7cdCjXIC2dsiOWWAlIs2Xtj
zprro5WqEsxrjWO+mBYmF5l7PAQBMyw0lw8D5KFD1dC5jM2LaCgcajZ8OewIg8GM
tVKjkIc6AACq6piHt6ATgvwx4bAbWNurpTv51TYeSGGq1kCXsIWds/YROgtSZJKr
Jaz7JZ7kXW2ka9bBOFdRUkMzqIhyXwx8uW4AwIQS5FoWT4VEr/OrSZRwmhg2tZW1
foMFMFnT4kRgooH/CMoOr2eYCXbFVE9QjwsSNIvFEI6ZbRA3MP2Vfq8mJcGR4oWM
Fl9zXBhzGfzWvFlbAfQlA/0c6xrMbdI/MINtrl0pmnE2dSaD2LDsZLIIEoy3zLHi
LTNXQjvN5uOXgDjApVbqQU5k9jG/0j1LHqXQDvDl9vEuq5+EBUg7GcInqLIAZYWl
qe1NSk+7z8mISQYvOcYquPULoXPiy+WDm65rR4bOV/YFDEqNAiPMNVhFs/eIwCHh
/CWOV6cas+QlhwPkvB5u9y7/f+m18RVapAowUqZOAgqUUpsqVGEspdtTkj6ActNZ
7nAO0qjgaGl2Tf2tXuuokApM8DBaIeK7gfk8KSHFI2Nvqi/fgD7WEe8zdb56Zaqf
V6ChIDxVFuEhNTWAlDanqhxVSjUyejfoPnIU5/jOMbBAD3ByF375r/MZE/0fRRjm
2h1fnVXdbipok1zkMrQEQ4N8daZZ4HjUXS1XFBfYLOdTb2my/SsyugmbxcO+Ot3Z
SOJ5UxPYbvr5zfl5j5fgyc1b6j7H+Mi+D471+pMsHy/vqHFiFE+adzqixIASSAI9
+f05CR0Ar2JxNO+B7hrOUotmHSlIGz6pllSyvXRE2v8c/S5t8qA0ymk8uKG37+A5
xtZ4R8KFJOeOAqN/eQPhY0tpgWLMrPXbRFaeXoA4ScTz9Nfjaapjl60s51ueaCwx
OoA2fYPaiY+YP5OC2r+W1/kqs3I70p0/g8v/5VMQR0yLYD8cjD/dp9aK9bq4uNoP
qkTt4RvYAq1E1wcb6XHTxFM2btrQxvT6F5LjYtvDvUIpH0W1cjPiHRecXRVyUPQy
2jtP2WyvydqZE6ab/xhZoKWbDWLHM16tIEIhckpIKHc5Oq2tJZxiAYsNA/FCk4MQ
xSqQIhIj0NQS6B9RZq5yf8nYTtezv9WYV/PD8FZYiu4Af914wBvOhZQB7aHM7uXY
JUgfHHKWDd27iV7XEl7PbErE/Qe/ADK7jkNEpyU4njgxUdx8EWg7wUMfRTlatWjT
hwkF60UCXRmsLByr+QT6ypLlyv0Jt/V1lkj4LBh9xbY5idwAoby6zHjsUJW/w3Ab
azpgXkRi67imUuoz4xnyGMvRstb2cDQpIUwMENrDv9n52O3GcHDyyB+JP1X2Ko8P
DcbLh5+yys4uQy7+Ebg0gXypbFWai17hf7GC/nE+wguwGqPAfqD2P1EGvOh6xyTL
mcwyT3R09iepuRaIlktd38EdSzGPGxlRF3+iUGzXiBsUSgAy92Q3CnzmR6rIlz6g
ElF5684a6kCbBCEuDt+VTnb7bVwd4PoKp7Edzxnb8n/tCgvmmXZCkPrxHwRZjRMS
HE7E/QtlbgGgV+Dosgi0AuAvN5EyG3matjpPttFisGNzc+t0tISgT+b/WWse4A0B
ROyKmmFtbl9BTT1vS5AdFuY8o6Pa6MR2Bjj7wPQ62mwBYS7g2q/nOWIG32brxTvh
hLQv3VdySrSnuu72sEtHGelKw5oLVVPiI0GPeoc1YTcoMIFWj1DspcPBIdgpJAF8
24s/3/HQk09t1jm7dchXKsgd1vEE3XgmMdMZWlpLS4n8oFxrZS7evAkEQvzRTjos
QqXSlyQnIh3v/PQKU1qfkYsmaJkS0iiwRZ7b5G4rJHmHUPGgultHzdQkkDImSi25
Ta5Kef2LXApVc7+m5SUKnZv/G7UqYz9de3+TKiXx3Yn+IgAPuabXeqwArb/vDa79
5SF38Yk1sbDxp3hxM6O1oEI0FFvbmhp5Om7WK5DPO3XA24+rDu/KVU8650pS3KDZ
HBRZ7E/UKBiysEXgWHFgEzOvheJEr2oaD2gjVj8CnpLO3B5F036nMCxGaNZ7nYRS
W/200u5Sm/YEaDvQG5RYpHoAMpo3aG9FVgy/z0NL+nThh+FT//d8XQ9fV61Tneei
A9c7EwqSPksjpCmS7bCrc6PsPQCuTdwgOyPN3J5GH/9GH63oMpkg0L8mZ30wpe/3
q9tyKdlThb4BMn4K3kvFCWA1I3fh8b1oQ6LnATyZsUsI40Mhe2H5hfx+WH1m+Gfm
Zsw8y8p9aKc+QPNAPr+kbjZPuypTyjLToCHyomWwvTw2P+CTcmrDEHjCoa0kLIwf
DBxxXEETKxalBNCVF3I5EdrKPK9STYqwq9o9BCcRxvc+sfk1lD5Mm9HkHQ9tvA3U
VoE4oy6MYwLHMzC8/GhxgaBrAirYxdKbR1ocOQfFXb4vQQ8M0y1G63yhJiZ4D2R/
NH+WP4NPJtDqzoPNBdil6zfrxGHDpgVqEHc4vjcjiK6OhxMXryD2Ylcqd50IVSY+
r95dKrhjdVvALzE2FYnEjE6GQg06fbTuGT1BtEX/EE9CW7aSIgdqmdQlxyDL02GO
n0c5ifTC1EnfBenrFYStjL3MAllntGMd8uPBcEXz1TTzhdx7OfMBzb2CYPIPaqXZ
t3qBRBlAXRPxp4qNzs7VOQky/F+qjern1GnyRJPsaq2nWFqNGdKHw1IcbjvV7FBD
rnDJxpiZbHfb7ngK3+vthlcL/9+Fd2HQR03NuTxhLlcSd/CeXqpkcVysLZswcvHw
zorhQ+OAFiWOs9UvMeSKxGxLGMOqElIVk68B1brQM6X/d7XCtxfSEIKey2PwqFLt
pXEw+pSb6Sd8dffxyEw4IveLPpTxg22AnzOR0dkzjuVOuhC6rrtc/i/ZpChbiO6A
mpDWt38suZtEL3n9+xjl76VXFwJyLVKTRDCQQ1rnfrQEaVmwKXGOIZpoqP6IyCIm
FQzLBSjCRuo/LSfr81qgbnv1Eyrzlhx8AqVGL8joOOhk30japle9VhteFi/UNJUv
N/ur4hj7lvMOpfaC7qZwUcLz0uayy18GzHO7cX+qMbKpyXIaLuQ6qXXw84qTZ53z
R8i9AR2JTDS/OMrKLnpaXdciSSXH/8ZU4/sZpgRab5l6QXc3sH10L81zlWoOAEaq
VGy7YsGmk2DvbXu2JO/rZP/iSPm0tJ/2l9m0crT66V/gVZ/lryweUZibEUnUfgPb
/J5k8jt9jBIX0zmp2Uv3K75bFq4H/nWdCyZLyKRslOgoW9DnEJP2gcN7o0rpGPfW
2lJ4TtGwjRO2gwP2oML28T95oudimClalZRP5m+9Q/aikVW6/0fnufYryhUbo+Pr
cd1OCsM03/kt5/GItfd3FwavXcVXAbnX13Ofj5Cetrd1yUxTUmmaV4C6qryRbO+r
ozPnk8f16bWIUp0XSxSOD3pBSTx/+F+gqCpA7itnjSIeR2q+qxtmMZ7MHD93Wg+H
hoXYMWGP9uzEUGUCkyp09ys/WsCB5pEOurt1Wu3VkG4F7RDmLci/Xf/2nu3xyrbT
/bERNrjAcjd6BjqbDm/i6d8DgVsdCFrRQkDBNi4TGpiSi6wYi8/UIzRrDDtlZ5Uf
nyQ2kTfKdiIdAXgEZKy4Qt9k+soyXRgIZpJLi0zgbPp0hedTLlbcnOJDwh7gR337
qH3cOGD+mzLFuB4hZT8azgJG0aw+owzC2P4KNQpBKjqfDGkLLbKYarVegjYGf9Uq
Alm/hnXmd+OnPiXhUm4b2VT36Vttu6LxsN+IbzOcyHAqJ/ur2/4IO5NOJTSFJbS+
yeJSSkEbGhL+qnz5iS42rK6RbmHkM0mSWmDkRNJvSudpLqOfC9NnepHMLhEzMc+i
6o4PRGsNxuS+Cu++0VLUhkbmbjvO3wp88XjkyiSTyoMD2k8jHCliaFGEh138ImMJ
JxOMSSZ4CS+8+vvAEcwQol80J9KfqcZtF0dPppSIQBbN6dfCwQqtAsMnhWKy1HVK
fqgx6qoAryMOKLUwJ+aysrxEUNuEgKN9A8++Xj3cs8eX88fO9RcGK0JXLwMRHo2W
A7J1vWpeZ+ZmdOALV9RfZNdJB9H194XYhpZap3+dTeWX7pJJhH7SWJz4bXfME2bq
EZYcp8+L7Kks2vRMLWPME1Bvy2HIXWRUBxYbrK8MHYr1MjiM968m61mF1pwyW9MP
x5IwV+HSsIQxTb+QUryfI/cu4BmPotUcdtUpjYqbF10BhGMe32VtbQfO5tAB9wFA
9pwjEpNzefCyvA2RgRCPatqXNV+aTStZOqUbPnS06AsHVl7S613tBABKJ2NAOIpi
N75eflIz4IhT7URsv1M9OMmfxvb/27MbjdH6Yjk4aO0QzdY8AMbI+F4B5Ry5OPFq
1P2Kr7cVxdrem7x9QQ8y8a9m8jiBKuuvIXpkA/yl2P3FJ9lS+BgoQlDnZfcDondG
Q8/Jabl39kgEFaDDDES/AxYYnCulVfymLsCuNlvvuRbvOzPjsECZVLwFrgdC1nBx
IqcBsXYQZ+2SwZ3Xh6v8LJm0+91looswsZ8Z/pryoHIeEZVvr5D9JU+boy/DW8Cl
7s6eF0TU1aoXh5VWCe04MpTNk9ezZUn2ueSLd4Su3PKaFGNVPpZm4u8t4INCC/Mj
PN2YV3OfFYgK8D9Lb7P6IMMIalPSRbvhY+k1P9lcSLrgNc2UELCFB+ycOFb8z8Uy
cqT6tOaWKpdSk1XbMfCNPlGYG1Ka+ntxBWz8xLchHjnwoh5nzWAmVYJDMLS+yQj9
vNTUjRTxSFF2vmZecObjXEaH4WGz6ac9vvRiJrywzVAfvoOydeOYmr8sZlsRs6gf
CJKh5AoDZL1a7cCz82qn53t+iGRfRq3LJLsweN2IveMJp0VVMm/OD9gMGlkuzsDT
R6LO0EadfTwJVcoGzVmrleCmVo6kcHm7MhC7MiN9t7yRQ0nTfG/PN1ifYjFuNfFl
QQfPciJOSlQHvEFjDG1yEKNFPptkEcD2EYYbjK9lMreigp11R8BIcj10XdWwcKq4
0frrC1j8yE2W2iDLNEsPE0HbJSOJijoHoBKfusBv+HWrLTSH7T1iVV17Vaz072eM
nd6Za7bSZPISlTemew8bsAjHdvqvT+fATabucDyTmfFa1LTnuUgqPCzp4lEBst3D
GvmlPx4euUlyQ8ODBzvC8cgfEXIhNik7qwULMPMspFQFZy+gG8IN6Q24EH4BG+lL
Tiofz1hLrK/JKLCGtYESxTYJy2B37ML4nVxQz2U7du7fQW55EigNTcHsnsa4T9Dm
JWW41vRLnTsAkGtB7V3kxI3tAj+NSKb3QJ9otbLeoicCLcUl6Ca0AHmtbIS++70w
KeqXzTA1aXT1cMH3h4Bnyj7qhjaAKIHb4vftNFALWXyo+ELt/ehsoYjoxNKBa1pu
vm5OhGjPbd7hweF3ZM1b+pXHyVS/NGEdKLKxd9ppU3+mDkrZa+PHBAyxJp7Xpz74
QomR3cbxUPO3JbbOFhO2NClYefR9gPtMMlIpe97k6AboqI32ZgCO0xGVXEuUgfjs
hDT/JZU7A1aJ+6ZKXyPCjvAaDm2oqHeNMh/6wVPSKXA=
>>>>>>> main
`protect end_protected