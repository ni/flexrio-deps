`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 19632 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRvSzIdqqwO5JLOHm2ufP7Er1fodAbHG0kpDIIj4Ba9VK
F4W01eowefxcxYxcjE1xNGJzw359TyO6XR2J2XH/Uq7Bur4R3JNQkNRc561sw494
rB19sKDcKwEWksqlMLi5A0rnpgt8hRjGFhtxwKDRDo8PZ6cJr9BNlMbK4GpRw94P
YqRYgTMs4x9fr3oe9xE1ejiUAm3lQ6AGcXQ5qlhaUT8Hyy29FG795wQSh2cKpD+K
A6pDVjz4rtDWdatnJqsB06FKQOmD4Kj0ush6MGPk/t/iWadjlGxAFsLsyVgnKUfU
PWLP4Or0tznOFUrbrMN0EMQKGUHMPyw3x6FoFrcw2GFuWlCT9hcQpi1Gr4Gl/Uqz
cuYZKQ7DQ0ZYdd2kpScWKaUfpoLrA0fTAeE6/FMKkNip/xun0Igc7qCFQqtyWOTj
W8EE67QWkQEPOtSH+uNzfJXB3WtnWsSI9WKHJ9TwNDGzL4J/GCIjDn0N38YMFLAz
RTLaUvHAKnwTvlYF88hH8a85vRwxU0+3OKQX/uvbXd2uZjMPg2nUU8BCgtYsYyJC
eFap6dXSRxBLXyTH5cHieKrQVyuOEakDnxFaFqZ+qS6FLSFFlFHhrto5z8KdpjuO
eUpQs2AJyzrcdffBYrwwDuw+t0juekF4bSp7PI1AwE2c73KL2/6YM9J5YWWoAhMm
O6G5wTXzkTNDHi7lRmNdG5xO/yYCNl/LkF8uN4/a4y8OyfIaBIp9ARclT2tiS1Si
jyaGy/IwX6hopdtf9gSM24+pc+0b8YV+yFG6JAEKbLj679oCs6r67CR606YKvMHg
fjY9Ze7SFFvkyOa/bed7xInnbL9WaEiNSOGWBtItiEYfDIz5SLYZFfkV8j84O+v3
kzSI950CyAU2a3t6gFxSIuMagYXqWEECEMIdOAlD7oicJMyRr6PojIrUwA8DoaDf
ciyXZ1GVbJvj4WMCaiHUpuZKTlwY+lcsYnaKnkPhdcr0pWIHMq+EaDSrJbBRoGLm
dZQRPuInY7ewjib0uUQkTG1tWD+jfy5X94uphC1n2FHVnzysLvV6pv/jpozPIlSR
8pQ5N5bvBQWgu7MSNL64usHMvNWFsJpA2Ck/+zPOST9D4EICXpQ4ChLueu6HYdeA
GZ/pwpvreEZSGkf/oT9RwLVP22yyOG67es/BOxBbk5IGlqmWdy0xS61nfKdWyM12
hjIv3StL5nim2ah57am/QRy694DMwCqz8rtfhsiHUPwLxvtr2XoNDFy0cNvWSlYv
9b4LuFcBb03q/hpzf++bMggfNEGQBX7Frpdi3HWN8Hs8i5rlg4kyH0P1Tvi+be4x
3aaXhV+Il6HAPI6anVqfXa+L+i3WYs47psTzYAdajKLtKe8AeXjI2HTG3GEMKPsi
tH5h6O87eLeCJFY7DtM3NrDAhSRlDbYuo8Y7noEftD4wUDtsUkkupbgN5QdOgscT
z5OT4V81/xRWgSNJC8sgIU5VsMmdwVE+OojpiISX9V7kZYDHBcf6AVGv5/dmP3XM
++e9gE0gVQNqtzR7jwwdybAaT8p3nsEjU0yLnSczX4VpY+MiASbuFbMhojpm+4DT
a6zWy4UtSXFOGCmQh5zZA2nZvJk7+IqyOCBayIhYw8stRJ8VrbowCK+QhcZ6PM2K
Hm6ImhPVg1SO1Om60IEu6/COLfVZDUVLPoOFjh+yzc37k5GZ41tMnX1wsLt25xWV
cLjfl2CYHd0fcAqpKoTB5VnF5dA4/D4ll6mLI9ufM7N9kiKOtbUk127UW/4p0vlx
pGYBb/Evr+qFujjB2yW7Xj8qbGAreI/mb04TgiVm7RqDRfoVRQD95kmddv1YJa2x
gyEQVx0W8UYhyWrPj+9NZ6HnRP/V2wpq7ep+Lv53qQlarJTV1g02piX0/NH9kmMT
lMEaPxhNLQnXxpRxhf3RX3uYfIQkH2cTRq8HSlttTdWEegiXV6xIkULJXBle2+f7
278uro1H3GQrtfxFUaHBk2LdLKGOJ0cMJvMsrpzzmzVoBF8oaw5NNvU+0Asi29wF
GDEtha4zNn3Lgj4DNWP9PzxIGAE7ZrNObd8tso2vv/oQnuakIMa8CiVa8ml9KaTB
C5zUug9uCTAVGQV+Seay94ZPX32peSw7XLvGszY4erRrMjya3+FRuRLr27sfDfC8
nydAVC2Lkkapt4mYvcQ7kGeBkJy5tJydTuyhQEXaus8WJ7pyM1DQOZ7t+d5M14v5
N6yVuh+T5UMNb4hoTurOmC+y78SZ0SBRTRoONfjQwPWwlvihsUi0RbWR1g0q6e9x
DUJ7e7s2G34IZzavd6JiA1C0iQ7J+gGriFfOLojuBZ+BF5zUyTgyRRUAGmIbggdg
WNN7PhLXtAr+7EzaDP46Lf5oI7AtJn4eshu9UHKo8lMn9GcJgR5I17Xn7uBYeEdX
Tc+IJxRHq4JhwL4D52BMNrYbT8Oie7cXW4Vr3PNyNIuM66EC+v3ojp91LmCFJEpR
BI2LFB/CAX3BVFOJq8dKEcMlogSBAU4D49yGCtREoPOO6z+ukHUGjwZm9cVydVNM
VdWRB+QPVPz4bRVVbP0JuvUhfUeo0wY+r8zkGzjK+FRJy+O+cwTC2GKgzhug4GR3
nmE3rNAR9rXkTS+qqcfKcElAn5lv67c4mK0+QAMAgv0sfbxkLuP3rbGCgOZN+qCz
Kf1eyhYNj2579ZNxM8IvC6Usg6eJ4mfPx6oia421qcHkqw/Ib2GBUdtcGBxmUXHX
fCbhm11hVCc2so+MUD4lr7bwxhI4tpD1fHW0ANZWoxUbgae3A8ENe714fbWWD3eb
T5HcYL+1wB0srNDHa/GVUxG7CO9ALWcEeGAwaMMoPo92sfdXMEFFnBW/Y4PxqKFi
4J4RA7Ocw5LVTHPMi59f5Shbbh1a5vPAg1AlH+PGWxzsHHnGnKBsMCId0f+LNbU4
qzdIm3EhiS7Vl8PK/EM46AwrZ5AiN3RpgwyQ0lQ9R0QlaPzkhHvj+Y31UXmLRQGp
onHZUBQhORuYoy2YsItYMRLaXiO5k1UV3GFR06br8rjOCxGCo7m4r0LwUtSIhEkZ
LIimCIWQQTyHUzHXKs4WlmBgUxw1rI/yZPCmBz+dkfeA9gM3nrVYE1rSwxB/55Z6
bFBDcGEGibpgBFemx2BMlvL+WzX1gcC0WBeO4wt1YE5r5Oe8qtzS9pnMYYtVXg5G
aZOOja5Qo63+mVqiA/h+sThegR9QHFdOzBJ1e/hQNPNLVf08ExCz4sT3zF6b+csE
QDCeq3Prctjqb8RfZYeFz3qGg/5ZCGsDdhWbkAUOFJ88CUM/CZEBCVz9WLXeoIQS
fWAHeH8scT/nkzDqva+jt/cjjO7J0dD26EjSoPkOPrb9jV0skOyeSXznWpnXf+Vy
O+XklHP0H1AeVFRFmE2X82RGK2sSgMC1VNXO7TMed6MnViEsFWJRS51DuIwKoC0b
slq5w4n1G9xqTmtNil6/Fj7WOfBqP32GfQGPkHTQRoj/1pBqFboyCqnfLGnBaAvH
YPuwnFI6+FQyUQ8WvzYBB3LP2BaW9vmCNUpyd5ge2mBHIarAij4gs+QQ7xLJvYr1
LNhdyS07IWWjPyCGlJjni7md10cUnSKxzblGBpI+Y8BG8N+nBSdiwJ9AuR+vXNww
9yn5qXKT6Nu7DFcLhlDDdeo3fpz2iaLdk0EVCKd9iDSDORXcjec0ZVD8uKWIscbY
gMRh2kSp0HzxFXFklvfh27SJowF0NQ4tRkwe4jRm0ro1nX9jRV6ifQrWbQDjV0G/
qsifIVyTWDkkIFomuH4+FrlcbgRtYSjm9klKDhqaDKCaKHIB5X0VPzBJKbSg/bIs
LibnnD2hXt4GLFTPvgdUVOajJGrXtIs27hhp4OpWxMlEeCrga39xnK8t+eImeN0c
aoID3geXc96Jwp+p2rnkF7+IQvuxNIBvWQnfbzItB8K91MkoNopn6bVNMboebFe9
A6uW5bEBhG+2ROW79Rj9dZlh9r+8Yd1lLQDItFGOc6Y/OZUopibBdoDpS+u6OwhF
7x8W3qKzg9sPD0sLwiBRF7r8tBphvO76P6nNkL4QkrWsVlRjg9uLscpkniOjpPH2
9uyGlgfWZ73Wy8wg28HNUf2N/ltKWLtS0TqrD5QE1xdKeFCJvhHV8qAsPpPsqvw6
u9M5NtodnbBH5dTp96QKS/Bd9/VBfxDT3+Nh5jBFmqXwKlVzHsm6TtQJSdf1XAN1
BoiOtd8Px2xpbkT0SIQV+VAq65pq924RPQmtFhkEfjsfCK4E/TBFwLAVHJusogrO
mCl8yfLw0Y4yIoeVTzZLjEtR22X/7Q9OW7rw0sqU0bYxUJWDeozs0ifWpEDmKELZ
uE/P88JMln4OwPiohgeiQZOEBdKbIbDyPPnh2TZqMb8WmoUOaTej/NmmuG5Szj4i
916oVPxXr4/HJBKmrEU1aZFbGulo4paPQi98BMlIs7Ihg9aX7SumFRRAL5ndpxlx
+itbD1IX+PD0Q1KQ8MpSItEI3pB4dme/DlvgNzVYtsw6p2GS0/I1fqBxNGNgDt8z
Av/EVnM59vhAFLUrfya0pi7AI3/RZDqyZmtkxfevqOnQq5uklThAzT5a+qvk5PBC
GfFUd1vPixg2Da8lvo6zjyfieh9b+3d/3ek3oS9FZB7BFsNSdh4HbxKizYUKKZlp
w7TYIXl9MiHfLXveh60W2H188KXK/jff65/9t6y9KxE/jbTas/HkDzDKfimTnVLU
gK7oV5cUF/eIx8hWjRVWDI6GadbeKUVAQFj/YHK4tAvK/VKmu+ssFL/tiGxu7Kyb
RuH5UUFRsQ5eEY+je9eTZFTjboY1z/YuXpV5VgP0TlcowVTsy3KDSH5M/XQ7juvH
JwD/JoFLbUBdQx0WxjQWyEcIbop3xC7s+TlUaeXvD62kAwZxEI8ht/hzbKy/N89I
5+Q9KqWntuvGBrkBw2a8FwFzD8zNdcP3YmLD5R+VEOmSNt6WSNjdsHaa6nKnmmSv
U0x9q/xE4eByiHuXnO5wALxNd2Aq+Om4lZ8Te0RpXveo4eiFmK2rRpiBb2308Zcj
CBTXZj4ysJ63624Y9B8O4wuZ9zoka7LJ+eoC6UNfme++4ddBfM/VlYE3G4ugpu/0
lMh/1rd033CfacS2/LKZGWXYPhCjwaUhGB9QZk8o7TXKIN2BqQB6elVpQuqbEQwr
GgIDcG5GzJQKx/DRENwUclTYiOO03dBVqxq4ByWUraZMk3prJCAH0dv8/rHgs8tT
LE5wRCHGDZNQ+t2o24ALlehbk6o7vBhJRDskB+iA/yzQf3QRb5NvAvBthJt6zwLo
EgP6ZfNqtWhXXr5dVhH7+maxJ8a5dKY7x+tlPPRcEShlOYYHKXxg5Ge3KzJn2ae9
hxgYXgWp77WvXMBLK7foBdJMcpCK4+hzdOMU0iNvLDnHs/oXKQEQnWhFRL35IQ5B
oCl9R8JHRKgH5hVHBtXIX3WhydWcrWAXqs/5OB854KvWVkc2bY/uBqDAr3ZlxySo
zOQK/06uNYWieEL43l6st52TZJkhPZvbo7YDwtiSTiOHMcv/F1RdYMjOO+6XEbpb
OwDchmUz9vsdnn23ijpO4Jap+9R/x9jbuPyPwKXvrsb6WxxgGa6xcRzkJLYtZr4e
EC8IIByxQSb12kkpINoZQSiv08dVEqAxqhqIi8bklcX4aT/vakGjSnK2KbrKyGvJ
ubbh1N6WlBHEeFhgYvdqj7o1yPkgW8r/bDA3n4dDfwjbINNYJGrJWfggpTC+TxfL
5BsxOeq65kw7+hL2CXptqYTpcH4acXsQsV77YEAql9DI1RcRzdcGBR8yai4cpR1Z
IQPFrwbCDDjQuTtFDZU7LmHbqtGYIBj3gtmRnne+T5sc4HbKlzTuFavBThBobv+S
q8w6mWBJSOpckdyKbjB162PQsrSAtYPwWqnSh83N/k8DrfcP2D9MIZzliC4P+2VH
hz/gM8TJRrJ+AzEtY3LXaMaCjemzh09du8/9QpHgrxaip1yy4v+9GxItMeBS5xcW
lGV2mgILi2yOeQh+Z+UeQXgRiSq+zyDBkcCDXwMwLX4YCswznCs5P2pU4qIHTkyT
J0sXbSrsZZUKB3i8yW1fILmhNq5WQila5Vv+lhtFHar5m2PRLSKcGnzwCWP6XFLc
2tMZzWEWB70xRNIi1Sx9KQj5gK6a3qatNQDV1nmg427ey7t5kws8PFQ2RtPKksWk
FjMvi9In9V7mcNtdASYlB3jIh26tpqV0Hqs76ZEv+NYskGr1BViqzTTuCRiLpKJx
8x/PslPr9f3zVYYtFZTaTYay4cD81sJWNtS1TgLb+BhUVNDT6UWw6AJvBz0dwl2Z
x0CitlJa+5+ysyt7UP8D9/YF2Xcb9584Lxt7CpI4KrFCjqDLbNk7IkVO2wo/ESSb
+2T7shjQ63NpnU6KV5iyrg02FIlpd5piC9H5uyf7an28pQz3kX6Cn02UOWUMdvqG
BOxI+Fq0B2fLjNv5jPaabBCd2X57P9/YRx0lKCfme02AJhirO+atAJ24Otaz+LOq
zaU3koXnVYmw9O4B285QugoyUPFR/ZZVgqn4PuAkbfcIojArdw8VMx31/8Cd5kSs
0IzMmjImN37b0MBiFSVt7QGVEBF/N4P+5T6mMWtcVqw38jQYDdrl7Jr8ELLMtJXh
uzL9KpGEc5UsykXwIzOQQZA1unsFgAEU97RX71DtVpTPbzm80Yhz5bz0JSH+eM6r
EccaHeyuJI8jfi3SqAZ642xJlRCz5Pf3cAIl5y1WyKXWIA6BF8/Ukhe/sDA8738e
n6ieYeFV/fpsF0uPYAlKZ11Eh0MHz2kTZI0iRtxKSWvwkXzJuRbSZcvjT1gC74A+
DVaQVK+6l7NUoAOM4M1mAU058pd/HaEycYwnpE/gai5Bbl07x12+x+YQr9DT8fMI
KOzZq+zy+Wlt4QMCnBS3xaUqYLPTLr0CXalpunQrPDZgA37G0uCCyn0MYEhjfTn3
qnzW4xAhPD5ezrvuwZrU5TZP26owHpDzOhmzYCfGY5/LPwMeqfgPG1Ni8zvIOgfO
0fLNSkwHGgfzwLpKnghE2ys9hM42Pxae2MjTyofFvys5qi8gvaNLUc67L/e6tLHW
mGOAXCaEEbo28v19laM2w3UvTZlJh4+HDrPWJVX3SgC1P26oPYVuTyRvYW2HfH/1
DXg55eOVkHjCMw9HKvxhWuEa0k/f9jOYkj2ZuUxDTQhSXKVJ1ONs9pwGbxYB+nTR
7rpRwoP3oURX7ozssF29zuOTuYDjhZGTxolfczQEL3D6lokobZDPKV3p54SI5McC
TmGbo/+MiZySTYYSAKmeRiSlUr3IKucgS/F6YM+/nvGnpEJim1ifls2TBfnrbVt5
IBXidHe/RHAWXb09DvD/X9qnHXmjGVmz3wnxtaYQoXQ5FG6gYjxUzLLtcU+iKOBl
9B1xLJudL/l37mw8f7zNgdu0B+CbORquSEONwtVU2kdeShLdEDq73hB883tVsyv1
fGOV/w5KHL8egjMp7niZPZR911aT6DufQYxbEXeZyQj/YesqrlTBVVXZZbo5CiBa
bHooUoTSofSf7/GIx8UX/iAtESt3t3lZJqqDxTfZs4GUimvjemH/KnfFcYAkKXLZ
WOg0I9VOw6vOt4aNE3lwG2ag+SHfTM9kYFI3UM2yvboKBpAjGD1bedCvvcsEXbB7
Fcv9dlwQeKJpMWKrlaWBYjGp6JEBLJx0Kmgl455oEhYUxgiigqL+Ri1ja7ku6IWF
5SIePV1eEa4X7gpXA9cNnfpnBvE8TwSLohZSLozDaAEo7pMQEvNWgLizMNwTRm4a
OUWCplVBLElAi3aPse7IFTWpetR84RKBZ1+t991XRy6Gb1wJaVMo6qnUxAFvqpkK
IsqUWk782pv8S4unvZOtSNg0NIpJV0UpbVfwUYQg37OfchmB9Z0Wnkk6FNq7jk1z
ZPmm2SGL0DFVKoOQEfGKlRj7X8nF+hj6tbwVKxE2dUIEvbTvFNoWPxczvBYN6GGo
3z6Mde1Z+wjRdx+BcBu+2ilVSKJouXFhUuV2vP8rGYX6KaBYamZH+fLxvrc/LmKX
RsbzdE32go/9FCVNMRCMZfR34hr/W3grYlTtxO7pDFjafljJBM3VImk39q/y5D5O
5DH+zDNmR+FVH8yHq1D6LbA2oWYlIDC0dtM/3y5HGOQVY3pFFy+KZQmIV8n0A1ng
OCp2/IG9LC4fzRzAnr8EgIDDBXw4+u6vrkPUXSmfqZznhOE84zHcD16IBYd1GaQe
dvajIr89qLPC7Zzbebd/IPzJ2iOC1QTVHGeyVlWjYCx6ijqN7UPHOqtp79l2kbSd
G4kP7t14VN67vo+Que5EQhd7Jv4st71R8TduhArLKEeiJFdHbbKHgL8UJQMr3h0f
f6GS8jsjwHmcgb7q/iTVTr/FUiFKUtMMT3iPRN707886Hg8SLJ5WwIPMP/wOYXYh
V2fCRgjdLSYH4008qC06GhL7rlWdvzuuKqIAnM2jrJ0UE1Ej65dSV2h1yfH9vCWY
tHo6mNe6iAKGIZNp7d+svpO1ylgoOp12B8ULyLLe7aECr37gZfz9rulEOXIgMAxR
e8UE8Hk378Wsu7wY/qkK/Cc9Lf7z9ZdpVkh7u/pazB/Ew3vjqq1/MhKOnUEX4XFw
T75QDY1UmD+S/2YLsqQZr91VLZb05haIjB0KfqCQwPG4TdlXlm56ZA2haL6Bpok1
vsv4tMtMnZIpCOreavN5i6E2g6fKYQCQuwRNReCJUlUq7qn8FYpw8NRS75ioKROp
98MSvRkwH5IjflbNi/BEIpoJSELv7pdoyJz/A5xjTibVIHOEnWkLIXiiM+jZzkoz
bTsSUSwXsfPHogT9X6GxJEHmaw2tN9ZeEWE7gYM9OP+WrWzkzMmZT5PXIR2VqIKt
8iBxphiunZUYL3UBCmmZTKwI4twI/8E5TW7F5WY1RSmzOhdRjRkWOFJi5STgAVet
h8s0v1I3SKSa9sJE3vYHtvYbPjY1jXVvlY0PohbB9NQAS7rcopbBhcs5vjaoAN82
j27j5ofIiBn0TQRukDmWf79YvCdJINXx4mLIYtHR8tqBBS1A8ixjMU21I91HBayz
54UvcBC0StBz3SdVwDd5Hp+DVYlfoWxg2ac4mR/Og150jEY1grYFoH5v38q4kgv1
WpdcQXWaG+bFDY3qOd5nejGxVe/Q4sDr86rtguaVkPRWEv0QYCtnnykR4qZE9xIX
zgnNMQiDRxINepe1xGwpC6LhnDqP1+HNbMt/20Tw6jx3d6ZYkcs54sWfObvfHlFj
odATjp4CPKT/Qupa1dhv4yYr38e2Q/CvAGDtSdzKzMuQrVgskdtuNuLF0F0DIXqJ
zqFLNxKtubcIHFkUB/Akr30BjGewDi6iV2UK2Yu/2wKVG+t5oEO77bqHrvLKQS73
IEPcuGloLaKBCQlX4OmHp7km3tN5tkDwBVvqlWyWyOPSj7CLdIiGkHz5iL5yTHFO
w2LD8g/xCvT/m8z/FTNv6cbQxN0QDYXAp/fuUkFZmiopQErs4ZsUD8UFA3wzvLzM
EJwut7gBa4KgFLOuYRKtvP/wsaja0qHg6XLcLeUvLDMxaOLxl9Kemkf5zRj1g5qg
fw0EYBeVVfYFkRbscruLlKT+5m1xYVpl5y58bczb78q++a3n1owZJxLlh3FmTw2N
Mb87awI/3jKvIrmszEijQ72k9EvqA7S9KSPogBeTjXB1USCE+EwJOX7CIeQtYWWT
5A9t/zs9Bzl/WP/llxN6tKo9WkqM066Z305jmAIRuhWdCPS22TLiW/2nTzUZysJS
CASnQ66nKx2liDdQCZ75JYSfJEdMYOomxq8/HzYYZyhlPExHAznUcc4A+O3z3MZ0
avw4uF1y9/sCc+l1OnsgKjDElUcQU4JByIvRr6L0mwlTdF1v/6vNIE+BFKd8K0Wu
t/gS6QksRpuHTMrNDECdJzQt8snHXfF2u0Wu+Mmm25pOFT8kzei3b7RY+eTsinUz
B+OebRbsSSW5G2/LtmdEr1k05+rJcbhjP6iZcGO/8FPko01K3XSwrD4Z/Flv7oxm
5lLN2sBlKPxEZ83+ewWgl9ztX8Ltm14SVRFuuK1Ycu99ZL6EWz/9CZqIQxsUk0ab
iz5PWz6F4Iyh05ttieTrtkcePDqxwXNRViCOV4HHI3PPzYcbJib53msMi/qOKvhz
72RVmTQCAmqJLLwW8UoClUPlp3uCTVX7MXN8O+Y6FUfBK73TQJwLDPk1KIaZQQXr
oUuR1+eOwi6Mm4EsPvyMvUk+Ng+OR3sCZPOfPSf5VtNj29AyPXy7qxaIbpc7AsrB
9fMc2OKTfd1AK14/OLt6EZuBT8mM8Zpqpg5aFqKvYgGEZ20FVN0Tgljj3D9I/KHw
IMOy/sfV7kalncUyvKLq4K/EHM21XGznEvTk0ZFE74Imfz551YkaZbm9K5W9xKBh
qZ95bRgNAXJ0Bw7oJGRWQmNK9yw5LvxcrDwOx/UP0UTI9F/HtFRfqSsasXU6YWoP
gI0RU0Jtmulqz5acHmrf1ZPPin9+oh2i6qpKR6km4tq+CZ1y/NP88rsCza3b+RWn
sI9Ue4zWm09mumklQ3qlk1l9YP0LqY0k7sZyEXwKzmgOeMr0hCtIHoMCCNArEsTk
TBTmyzfYSougOoc/6I4jVMEHmLKJYBktJpgj7/UC0MgB4wSgnPFM4gC7ouX5PAXO
OXpYFoKO6Pu0ZmQZpuRSRFgujkGxz6EBtd0cwS7uVZo/8P+P9Q/3U/ppPgPeNGmh
Cm4VnEDRRyPDbNbAXz4OVMtM/Zip+Dr5o+Nw74sJ4t4I5PHW4UpMyiFOU+g1gyy0
4qwj5iD0I0MpfIA3OfA3l8YbhXFwHEOzWmTShNG669SeeTeKD0laPpXr/TNshXLH
W5//OpNS3p+S/2o2S2LAmZa1buW+BWSEcn4Eva2BP6EcxdmYIpYuAAy53Y4zZEb/
HJuN6lO6atbEzwyxNkdMESwSdvZk3YmJIcogoTK3OLbqhG+ZEX3AzqfO9hW5LFGs
wGetXNuQH0fRWujU0/TfA8FdCXSwbb5ioO1ulsfSQCy9t48dJrVjd3UhrbfUhpq5
zSD39KyjIK4vD0a/ApSp6t34ZmkFGwEcn0NyWvg71U7hYGcwU3+zk1CdlgNgKjZX
sS0wV9wZ7zOQosDL2uAVbJ5xJfCnYHRulKBBFR3IS70+2lZtNSoh0PoJDzNjwsau
QZelKmuFsKLX1Z2X5hKnZ4Pz2BFBnoGZd/niHQJXEqt6FtAOB5pi4BKdD/Z9cDCY
+xCmpQL4iSVYHlLeXGOhkhsWfuVs2n+WBoX0nNv3qrfay4C0Une9cZR82WhQ0qRL
6WcQFSHGVQoRMEth2ZRYMBObDeyBMxii5lGDveaFjzEY2xim1Jix6yXM61BAgnbZ
zFI5b1UjZzmRHDUIfxvGhsCBndBGJZ9h3kCY4vclUxZpRtMnFxygQ48dYHeo2cB8
GYcWTSWQ16/KLHrvDxKGlbwVoK91t5qKocFanKXYMBrPyz6ooPUf+IMOX8vjb11u
mP7FzZxI9Hs7DIV7ZrdBNGy2TCkfndtY8Ah1Nn+av4E3IcoZpUYpphwVa+CfR7hs
g4xdnqgW9/DwbrfMaJHWPy18LpLDHqznZhzByN5QLHBTi/wJtjqPUqqBVEJba73Z
i7xm7Wktgd5MtvSlOcmIJIJmiVE6rI0SfSqxwILaXXCtjAW7MtnS6R3nUG1pp+PR
oetl1ZVaWr8F57ntUFQpy2PMnskwbpaxfjDf2eDTCqi5LHWBFMmjG73rK/UVlr3I
vUA+LN0UZN6DwenbHjgk90Yp/9ivf+YVSzqabaN0ZXlbt8L8AZKfUh240Qugeduo
J6jhbunvOJzdQ6aATt0+PGqh/b/2GJQbkdvz14lJKgLKLRbk4Lr8hj6viP5iWc57
UnXFn50O2tzd7c9OShl/T75pOJLMY11flYG7KgGzT6O9BB16hoD1a101yA+gitOZ
/isjWAmhleCCrhG9dNSFfrGCIROHB91khK627taPOE1/RPcU1m9eZ3WDNDnEvBDp
Mmja3xG4F4ET59BjOhwQDOgVh5smPlfShQSvT93J+mybm3dGVvRDgFrWfXyvell+
XGoVwB6fClGitjvdr/wFu5Y7CVH9+H4f4LQJ8yAxPzFr5Zo486Fbc0Ks1s6Bol7J
2tSJey4kq6IIo+siJLPYsIBuMPS4KkuvelNrUlRBw0Gsb7hWITU4J0EzEtLK7Hux
nxeG84yr95cEiZGfUd89FgMQmVBftvHCtdIeUZHH/3S86NsnheQjsdNYzK9r0V7i
RnPpg7I0AHri/yFQSlQFsySl1XuQUMUy3lqGv6fDgmoIPeZR3yJo7TfipY/j/wn2
ORngGWl8vpO8p268JKyxza1tSxtFh/Yv1syfx4hisuBPpLS2WMFrd8FCri7qn27F
ZiPIeWS/9WUEQsBpMSfbA6jo7YEmplRXUg/bNDIefN7Ku1CGkE9pF+svaFmGEBCe
yPtCq2MXASNnQRnDgszmG5qgzTxCpYbvN5XXYRjFuSB/cnNo8k9cm8wINnvGpwjf
73oq0IRjqd/3hXPJgOvHvjz3qMUaBFX1FC+FNggarYbT/TUYe/UqgwHc7kD5PSV6
IzmNps/ihLK7/PJiH1oWC0H4AgQgzfCWVrpdOqZlJQGVPAf6DxtgcfRIf1C5WGbQ
BrdAn60fwiR6r+5To1qTNburhbe2q+nvmLrkjmdCuyM16Y8fAWnUXa1feYjVtWfH
YquLYHA2d0hQRWTjV8fk0g08BicIGhW8n35jgAT+lZrTag2i6Qv2pscwsQv2IpiB
TeEbLesqqm/FEb8/Ho/qt8VzODozn4BFq8FQuKJzjnXJtZUa96KoPKeX1PC4Et0/
c2I3srZBF7Dk4qFTFbyY0p3wxP/8FfQALPikuaVoXBy6lLvwlFaRfyZMro08rT48
w3fGCV4C6d+fHOcQYGf2GHnIU3B5SM+D1EaTj6QGY1OGhOlulQQzgBfUi7wNQySi
VU+YlacI+aYvCH3Ia2RRLMnvgKasE2YpcFZv+ooPE/CzUhmRSp0ZL6ZGVQqgr8R7
1d+h1D/zA0a/0yvZuo58uB2bpb2g3pY4AcCqLIrErqEnlHTpa+Qwm8vIOMAnaULw
ev4iC18sSA7QGvz29SOY9y6cFqnx739mvoG+jTxbppFEaX8i+KvDeNas6pgONo1C
Dq3ndyv5T4HfAJRG2RkrIVzUokjcVPoDt4Dp8/H7jviVbqhwFHARC/d5llMELLNl
u9d1nVSyC1s8JCpExr2CbEIS1aF7jsZIpVGTBASQSFVrj9IwG2BTScbthV7j1Ru/
STF//44iuzOiLaf4Dk3c1lDnnPKdyVt3o7Sg7rEhLE42Qq/pV0S8VxHw27/9gDsk
G+ZOivL0zacNny3a3U6EsTaEl2VV5QS7LTE9wSbx/q3KJ34NBJ2DGqQA+sAO/NhF
J4UCk07z9Rh4Bk00zNNj36Cro8gj7hnqe2mmTE100jh6vZp8U7KDjI5doSx0Hwbs
5Ok7v+4GLDneGfV69q25iG2dt55AEYnX6ariy9XNtke/k3V0nOAQ7ywgqwaUQnff
6BNZcr7Dk1pOLBjcEfzzNiRf0HlJdIuOn7rxDfRSNa5ApidYQx96wSGccYNUCis1
eyQKGwK7M0lAzFO5YvKN6aGO5ll9+iow8IfuXGfOeCxZdBtOHJiRw6CShIb7rmNb
DSee1+iTRbr09dsydmmilV/awA2ggKGQJ5Urw0nhaB1VCtjOsCm5hGzoOg/zIax/
WeMKJth3s5apQaJ4AlXnE2E8Ig75cMdjLYYenYR/bEmR8T4V43TSJYrk45wdqL/c
NCVykL22u5zczvasUA4qJq5cVC6RhjcIhKM2jq6KMGFqaOKmltFt+oGLUiKv9aUo
6mKb0TLZYLaY5CxvBX+ab0XnX7gNlZzeEvCbY3EuEbSzSH7Li+E45k6xlk7drAaH
8eGr6PomkB0egU8s6a50eRrUPIENWYOT2RjQaTNy73AlOgPMNHT3k0xYSVDaPcTu
Sa6PW6YGKLn0oh8f4mjor9eVrZ/nN5byooUREw5ji00nkqMy05VIaYl5qiiY3Qph
7f5NvnOUHj1Uwr4RT6vae9JbL72OGXf0BdCIwuVrX4aNWTBLIe+TPVi+sEt9cSAz
gEtaLZ35IlN+XcdpUHie9LHiITeg/irwmUW/wy6UClgt9WkBNCNZIxfx5l0M1rcZ
8uqcv3id8Rt2pBnXFsVuyK5bc4liHyGknxKMKbrBXbLYkznhjmtt7CUuTHaJbYTF
UeU/ZCrgBvHmbosIw0YlNCuocnvwZdrQjV4QsUTV/zH2EJK76KHBU7jYu5j+aLJd
5ij788yeLGt8gu1Q5wQV1d5pJm5vAB6W2uWcGVKO2ETKhp8slkiyfdz+/mE/L68B
XXZNAMnDS1l8mEum2uvQ+DrUFWZx/2wfGnufS/BoJrPM+UARX7SsLmg+yEDpHB42
j2IZx2HMD6ArnO4xHm6yASIH6tv7VG60Bg88yluJGMl60PPc/bH5TC6mCozVYJjS
dd+zrKX77cyAVGrgHStOrouYPlGYlPW3PcEOEwAzIm+9Bafv+5ZL7kBnR2qLbW0s
cgaGfRgtBkjg6gcDpN0QPuUDyXZQcHGx3i5uwALI/P1eRWDcjJP/LU9+GJx64f+C
+3X8x4x4s+0PMISOu1SLuCsQnFpLGmPgYRmv3cWztj3Jd4jFUno3oH5qGXa1I0uU
6EKVVbvD9ZoXQxZqwxfOpwkusFEZuQ38KA2tM5Pu9hMfsjQkkCJ0AUHMugxfOQBJ
hoME4Tbe5csvFi5q84xVMGz6TzfWIdFe72ySS5Ws09T7B1bJXbJQz4aikL4i1fb/
ma/YYLZObzMHffccvb55SsbanLXpZy9LAtmq0g1bNAsPhdvvxS3FUOue0f/C0To/
gGrQRJqtSDIUVq/9TQNEI4OU5KDs4U63Ri2QjnJGRnt1OCh6UiYh9NRtp4nxd5zU
/v5jJZ/VoNnDTNZTTh6Hh+efi1NSWyNvDeq7qg2D66MPCkwG1mByZxgJIDbTuLCF
7MNQZROEdHbaBAzzsdOmr1RT+Q8ktLaBmVZ7nD9XuSpLxS6kCeZMATx2Pf5XSnIC
BWKCATUhdsXFF9MY62vXw0wAwfjRSExXB6LKExdo9801Xhy7lmj0zcWmcFjDooU2
7I5d9IKJHrV1qHGlqBYr1IEwPDSkr6FzuMgzH24q7rMnMv2tR5Vx89jxa+o6apR4
7ISJpkZUo44NnLAsMzUuUcs4+Z1edIAIgN9AhzOeW7mItL6SLSYY9MMq7me24LQ2
ZayvvyaHFJaorJZPKU26rcBrAOqWif+kU7EM7YF4xHU5IUMx1qQ9mzHFYjtDGRUZ
UIKNNOoGWspD3DPJZ26vEdDQUN1ckWh9m0QJ+l5Erm0oHYMIINcB0JcxTxVc9lJA
eYtTrUqtZwRlK9uv2eYr/w6PVe8/OUNGsntP960tAX5qEXakLGOkaqS5UHzXJ2g4
cVlJru9kHBGswcDSeo+PBHTOwvjOLtNFn/hSu53tyAuWpzdLvMJmPU1G+lUiUbnl
l2owjQOfj3k0dO4jrR8Z+w84qgx+cEtRxkNgzIcg/H5NyvOziur7bqhjIOIMyE9m
avp6xGS4/tIz86Zrt+ERB6IK+vGhzjqamO5DNXBnar6wpQe87CPIWiEN04uwv4GX
dU1XDuSq7igtN23HZ7R5CmRU6pyBThuI0qddYCJGExaj+yNFZdrFdAYczElmM1zW
afKgtpJo3w7Pu73AIdgoq+TOkSaymGkYJVs8+CsIKhUsYPMWcrKwiMUGKnmUUwrk
vbOxHfxlOGyMXZimM+CYgcY/cpR7Mw2cthZprATWY7p3dWfKH8yER8BPCNB7Jn44
0X2Xv5R+8j2knDC38xN6ntStCX3S4wB4ee29JAW+JimrNvH/QdNsQfzs2bOxIlOF
oB5SDGZs+K2y6nvpejUOXTkbBJ3F2aACvw8Nfq0P2I/XziGpJZNUYpef1Ux+cbX7
H4y6SF6ZJmI1e6+wnxZQW5DSCYkkWz9ZFKmPC+d34Ux/oZEu1poMlzVceSZLMhzE
upKC3ypYUva9xyGdDdK49w2LeseZpUsXsFbgUFpuw0FPUyzrXEGGojWi6r2x1zBv
R13qFJ7kLP3Lt4dnM0jM9m22k9x3h09b5tagHvkPEUnlxdf8+Q2Wt38dZQy8JEkN
ckLtNOOXASrlBGchyoEdXXsudDdlpH+vqkMBqyepkb98WfiiaYcvB1dhwahZzfca
EZA3bXG9DINg1z+PmU7f/xVGVEWNUKW41tSwJyety2PVb5lRETtc9Gy2U4mAx+E0
0+c9pvUqzQxNolhbncXJChqnCBWl7qtIAJskQB6NWRSGUczpajeYo8gABU/lPNMO
SGPdUEnTldQEYW2HTObaS63ktWReJT1acb7e9Q/5GDsCWsKs6R1mkDKWSw/YRpDF
TkEC3CAUHBm6lu2StW/D5bHAwntpCCcULTVslT+JLHeLnWXLL7QA0jde6O/p9+TT
xrdIMbk3QAJ2NQ06kxzUgWiibNq7JatOU+AD/yflVPiPzBeYDBOnuUMSAofWGqlI
MKoKlvb3IebqQJmBOEgpp4/owzfEZg7gjo7qhO4ikbzd6j+qr/C7JdJ1YbD0uay2
KTX1Mp+6jHpCMc2+E5Sv6d89jzLr3MPPShzUpuN8DMtFZHO/BURJVoIWVR3uquwl
IOyjus9d7Ud1APtWQVLVDXv9FXXhqsYonTcw5MfsETbs4wUwDi7P0zhSoJ4+04AL
MU5a12vw7ZdDq6/H54rXJc2axWB/MCzrKHpHIHuyvNtQHQ4nqcdAWtFSkwgedTDL
ADILE3ZVQR8Ztt/IeZ8Us961GSKLBW2iUtEWJGlsCpODbEEZATcqQWxOKJrcPr0H
dkPjO0ANMdXO+MX5bDe913PkdUYKAcvCI9vZcn3pUplmecWjmCEUF9TVsWyRoO9D
u0eFWnrco4hV8m9jOCveEc1VB+jmlqqOCfk81xKw4Y+3SgAZN+Vuig6xCkleWgtM
E3Kuk6IcPLZNhdsExLT6uCk4FgGVEwafzr2IP98lei1oKcq2s/5Hmqq6i8BCGyg1
AlEImDT393SqUOCZ8nUaw6aInU0o4q1euJBqQfgmMNe4RmRI44Dd2xbHsJTU9eEn
V4zmeGetJuR11W4DgRPjWvFaVi9wcbNxSUW2cqpCWJ2BlzLoizc0Q28VBGb0fABe
DXjy8PoDkse2Qc5AtNnGYe3rFhbnBZU3TKvsAaLyj7ceXnWrzuDwkrLQLLA0GN73
5Krs7ZvWlOJ7iXDX+k150TPdUrP/Io6wsceWIj+yLBXcLg0+XGUda/VXinaAP9Vb
Tyfs28VYLIVtk2sucAPtEfYWkbw+JibU8P8afxx/0iVEnF/ssOlM2QuN2E0feKCX
FUYqF9oIL6PlxHoSMkryZw9Yxbieqw1KQIEGRrdl+TkG6wFbWS4WVBNPIuQmn8Tf
JBs9uYduI//AhyqJlqi2yY5OcPVISbIXmmRchxqq4+TCEhsWdjiDkhFtik3dBy3v
B69u/X7WIHW0fm2pjNa2lqZvlwg/0Nv2WO24poivE1Re4vNm3DQzgepNDoGqrCUw
ZsOfj6dcRIthD7Sg314tfon7q4HSI9xErIYdkcEyhIiCd31t3sS+MQLHqpqOVG6q
Z1g/zBNxGE+iFYKr/mIE8jEAWqB9HFD/kIZmgeDKi41YlYF2aE0lMJMNsfvbDI4M
pJXhG4k9ibwMRAKioWbn3cLWce9w1PRvtiG8dw34sk4ztFYL0yiVN30h0v79OGrH
mU3pIzgrHw2YTcs/b5FdE4ht1YVupBTWlFQ8sEbyIcRx0lXZWQeeiEnApmVqwVVL
6c3t0u36BUQZdheTw3r6ubcERkj48hOd8t1iBlSowOudH8M7QhpomZXv7i+RcFLr
sKDW3osssHewBqDmnXYKpAs4Xp6LWN1V1qx6Fqq4Ip2maBZ8Fwkj5gAY7A4oQkRe
tlHoTXjqePvCX+n8+FrB6Pa9MyP1LsMgldopdWnpEs4IatIigHLgibm2ILXqN8GG
BEAuWEd62r9QCWBgdtSy4CX9UmYmm9jHsHI+b5J9bUo2d7VuV9Kb52vG05c4/7nV
DQsPE/1oTLSeeu/0nvOAKWv+gnf/TRibZXtjw/ueJWeRFwnLNdeMddMpXiKo9YnE
9w326GXxPRgM7n2xmsFHP8Pi1qjd2MhCSPeJYRjZFiU3CD4c32aDfp+hcKbvj+f+
pA2RvB0Qy5fKw1utzTQrajULBMqx3vfurEUOfnmNtFNnLbcs5LhFeJOcu6/NYcxG
x2F+cC5zCBx2hOdUrmWq8sEh1YQGHOkbA1AwhE4dYsHEVyurLRsEw8ERtz5WMPSg
W9lyGHnoY4ESjmsgb9OlOA9800C36JoLuSaLDZvs1+RJVesEeMP8FhG8X7PZNAuf
LxbxUxQox9znvx/jes68VVTU8YYi85cIs/GWsn7+El5ptJZR7SQs5pbSENM6nS2Z
od3ikZ2E4lPK5C7wyJ5ZLntiUAU6V1GbcxLeNsx/ZtiMxfMV9XvcNGdBgscsUXpy
tB8H1agnSnfvNwWFbI56G6SKHpCEZ+VtAElVlIgyeDxgDyW42Klrmmf076bVPdZz
S9EvDn6GPxTrSJMPWSyRBhR0aExqpiWmTDUIb6ie6mPWgBakOz0yExaHLRXiwL4Z
7TKqUzZHjblswDHeeQcOQFb4g+4xHsIx7utOeRYHwRvKyL4Acjm5kdQ45mhMT0l7
W3sAGYVNyMRJlPJtyblEGzFNAuV5Ow3Cagoh9VQ1GMvP69NB/cP8/MCHHYUgeLwU
TNtYxn9LUUWxAfmSxIN0r78YqMs/+tDGJFkMX9/xTwASULdIo3vnC3AbEqMWySyc
NoTsBfLhm9BEmOexOVyF6w66sMe3dR7D0u1y/Tx3XenBAJGV+W5JVKZwMgXBZxb7
8IiMSujHgLYgbNb04iwftUDjvong2Bmuoxs82scuKA8T/3oVV2Fg4ETU0M/UuRmO
tN1+EhH/jEslfaS/h190CrQomPuG1n0KuJ29y66Hwlmc0J5t8L+00xIeKAnv2UF2
FYO35E1NHkZ6peHYmBTsqiSIzXJvCpzQGHuiVNV4aFHpFrFCc/EIG5O7bGv/Yi4U
Ibt94kM/mJz33b/kSHK+cEEpiqYKrMl0HsiYC0L4CqDgnWGOHWmVGn7sKDfLJy4d
lo2u83quGdKZWA+MVbk9KnK43qYQSqeQjm/iWUUj1B0ryvU28j5FWri8lAgyKa4G
2G1wnDlK4vaYzXQRhsuXFByeFybXcYaaYYDnzuSzCjA/g9Mnzsx0iDO1rZA1xYN2
i7tr850WLyY2qPEk+VuEqM7zNEWJQd94HmoHIiLldljT5rQi2gES2glIsPYdFmhf
D8xV/MIr4iqe//ddQPU3phV3TvBZi3vIIdMjH7Zoh+8FJ36pMaZE/l93VjZk35wa
w7B0J4WhO0R8ySozMK8UqDpnQkE2G7MFLSUVmHwtbiEYSet5VC7foDwQE2UazWDz
snHvhunKPrPnPmc9KTJCWmilnPeUTCln2SZ0LKPuOY8f9p+58j0fj20Q6Ly6SrLe
B+x6qPy4AQt8RsC0HNhTuLTXws7RFl0Lv74znRsj5bh1bkkhWNtAElhVPy1AtMVv
urFhFnWvdVQxsJz+XR9b/lxsbS875Gta6EGgmXGFHWjEApnXHSeOVw2yq0ybQ5Cp
bc9e/3o+tTqwlLTbxTU++ASCGrLUn6vLfjcOl94NuwcTDjGW5IrviLA4VPhK5eLH
FedGERvbksmB128LFTotW1qW++v6mhtePXOeNb4HB24HhVJZ4BFUzcg9UK6IQvBt
ibA8eYsflRL9Tkt2issXEBV3VsuhW/ARXgPNdXJZXcZC4evaKhoijxtaEG5a7L6V
jV3uDPIyrLcZGHN0XFRSGsMndaubV6ot2fjdWDWFlKDqY8bkxbfIRjwPKY9uvErC
x2k7Z94QkjB8nXxwnRq+8Js271/7dzcSlrVIUoB4QWuvt5ZtcpI+C1lKbLRyEfEF
MhPUNLPsCqA+5uCjaQW80/TKHU9byHsX4ChB14F+98vriNkZv/XztZz7BfiFQ6as
bAWrXCPwuykGFWn/ekI361CQZL7zZhp8jr2buxHD1waGsSSFDNkY19DZ3q7CdUeW
agvou7+V0BpSwX6+4jYK5hbccwfHOsqsJLRhsEysQOJM+OkT7RGvSfz8ojGtBDF0
jzN3zhnEO33OHNpFi/A1qGVtUKrMMhpXVi2NCOg55cRMXsNu5BQUM71QTeLoxt3t
5pKCvQLJ/Le/UgwT6NhdHw+j6AVpzgyx6LKogDe7ol8TPfZs5Lva9LqUcajJ38rM
Mo9tmDqBQWRCLZl9lwOMagU+T1pIfdSInFJveL/mPM9iM79WJ9AL/+FaPaBGL7v9
r9AdOyaUobNniAOAG0qXvbesqKmfvFPKmZxEqGDzgbM09YTfUvYg7b5xMg7bF+3h
97uSOF1Dedv6fZDeE5315ZVOjS7Pn8LssqKKLtuS+bSaF4GoeIzLG4cYg1X17TYI
+5+3poH8RoVIC9rahOo5Ep+c3Ebwax7NSxhvUQIyJyb8pvR+0h/8Rs1a188NxMDC
brD4QeE5jDfLFU2QbpJHDzdHz/cR2skySIK1h1kkiCBiMyM1xgYEvsTKoWB4xgYX
XE0ND3+GCwEL0a5UsS7hHp/4UbgQ7cYXptoXelBEl5G+Ninun1Qqf3zX27rc0e3G
ZosOw3CKi21QOLxKTc3XJt262UEuUbgyX7+JY38Z6ukLzFAeZqAGksbcUbcWx9hi
2fyVu/pcxtKVwgjgNOSyEPJDR+nWsUJPmYdEV7m+Z8HHY7Yxcsdffuimo5YNxYjx
LpxrCYb9gWGXvF/n3RYOTdItmjulgcqa+qjyznLAXV+XCAOY3UiEju3EtzsXSpLo
E6sFQkphDH9w3uX5fWKM+vmC0c8u/5vrkBmjZc0bj8j841n6mfTuqvc/stPIgaoB
pb45MNtR0QK8HcCeXygi9I1y0ysOzMV5yVQI49rsAQ9IIfI9Mdr3vi53pBnVXWAC
e1dBKBibiC5pQvcIuUDBQ/IbTfpLbMqQcMmwtGyyyCRAQcpZIY9IdnY3MdHlMx9S
GTSrwnhXrvPS+tk++fRf4lsSCsZFgyfL2P+7QaxGRJLk0cKndKwWQYQ5PbCoeWSM
uOfBVJ1fKKg7/3n4nqg0ddB6AEsk0coWFGn5lYFpSXfDWqXUgPiw/sOhSxqxgLyc
BDVIu6koQuxxq/zcbZrhJLH9uVx/FinGsppWhpDzvhn3SsPMKxfNelxQDkcQUdmz
biep7FhEUBWH8X60Ol+Wn++IYyG99cCR4aTC+5zcuSFop2K7NewkGQn8fuwW7FRh
Z+2sUiRcydpRFbNzuiuBiW3nKc/AlcSmOaVGyXrbxcoCDWcBl46bV46Rqvowug8A
Fgqu3lWOoVifNQ0VFUEwTf0ql+EIxcUOM4oSGEZzM81GGilv176H2xpQP+9h99Nb
QpHKCfyrRPNf5bnnCcAwLl5ZbkXY8j1r3v92BXyF83Q24JRZdq2UfzYoBal+XmGe
ZTROEEllrGsckXUYqr8lVWVHrSalrZQ1iQ887lOMHrxXDGx8yrFtU5IZTzZhAll9
ITs1PbIp55Zmw9oacAKoyTTgqbp1Ggi7xnNe9yPY98XtC7a9ECXRQkV1rbsmhUDR
In9a/uJchF2MEOf4IqtFZqJ3wW9DaIMJMY0h8ePFwM09Ya31qpstXHlnEwKtuNTD
eOdXrzXZoPH8R0v229EQpulHre17SqS78xortAC4WFVdRuj+O+TDODigPC/MU4vc
X2oWLQjnf/w14p8SyfB1BnjwlkrxMuozMzmDAhjX2TUJ8D8jpQddksPf3nN51q5r
ORWDfPpqNSKG2fmqzr7MuWuAx1fNlUhTsIwmMS2UdCZ6S5phzPbVT9hj0we5WJN2
ZEF9PD/b7VZ5fhujXUkE5LkLt16+6/BtVGLxSVNqmcWA99BJ9zvA28oqKDXVnh0c
WuVGOoqWU6Gd8BvsqUDQF5Tq4JfQYtkAOWY6/pIOH1i460cVkiz4OsDGD390dOyD
x4CsyGNEG5zMWRWxh5CbsJZnwG6/Aegp3s57kL7t/7XXffZgkF1Z+PVeKtIAqCbl
P7FcVEODiolOycYWTynUvhkuKnKc88X5WfLdMzCzhiObIep/I347Kqnl95xdh8Gk
UmFgEbKh1zUczPZqbHDdcMqi90xSebyRKhQVHIbN27Kyjc5FVpzRk6mVq5LBLNcx
tHAo8GRJf/Xaai9DayANv48pg/3glWd+uB3zUXL1uc9awrtkbHJZy6G9yoXZcy/1
sdOgOwI2XpY0+DAuLCPN/+m6PFcHir6wOJ9/301wfHIOk8Qrix7mH7OxLTh0y8cm
SmjON8+y3rzli8Kls6zWqDkbp6o10/jeqKbQ8TJ9DykkN38z5qztmELYcdjkIHZS
Lkid4+NOT2VmbnuBN+m7iX4STNVnIuxt5MWivSj31X58wd3+4nD8Ssnrt7kyRwu5
Tr5wQIQJUMIXY1IQisIj7ny0in9lt0VqGPxXUADfoBIDqF3b1E/ZS24ZWaPJqd56
t6FYjEhrb/iX7D4CrDN/TUF8zmh96QJgLRqpkdC0vr1p5E29LR6g7O/R3XGSKQah
o/S1cNWUVMG70UuA6uI6P37m5hp9VmI4STT3pWR5ohIapmyH6Lzda6W1ACr2WOmz
DHNuDCpI/a8qFSfy/5X5rIOMsToEHMPoQkN0QrwipybHKCCmZlJ5cvcbeLTTydCK
wQ+TLMjLQP9RhSaF0xrlB70aBGwvUvQarKOGpai+n4jI63Z+HD5htDTfHZHACkVs
CSw14rlKG3X6dGOFhXpmpdJsTnWCdtwTQIWTd+l27WNjD4oiz8kM5nSTsUmtEvn8
Lqj11bH1JXM2FAv7ShA7asBUC7a5UhZC0SPlf4TOG2MgXfotC2raJqBpu5G9M/L9
zdiDnzbEAm92Pz8QyTEOZKG/xYLy5wdw0MWcXTo9A8jHrlrpvMlAtrT7nKVJyqZ9
FvrTkL7ktWWavOmH3xrdpS/4TJDOW9pR/QctKeztWjYkWqaSfbBcxs6gOHgHCp1a
wDf4K8qOLupCL+GbxSO/TA1WMsRGc9DBm7ReCYi21mGcLj9v7+vp5Z9G+qF4bBIf
CqhDI1XlCycPYXBASRG04GvmMtpgQ4H+BDDEfBD4eiiWdBMeTNnCK64Odg7xQYZW
TAUq/EPk0ScilgMGAUea4qH2QAMdlUkjDU1xQIzEqeG4FPu8rgSm1DN1MIgQa8f1
BG3u5L6zOjPTnCDb4doRk9QFkZ9Or3Nq3yNDX2LDU2YVkXwyEeuSScnc63PsA+dr
0buOBiBmf63nQ1ayAH5Az2C/QUHw+undijAh8j5mLuiwXUAEJZzkE/GVBRdIGf72
h5tS9A5gtgnKyRpkZr3X3vdDMSwY5mn0bhW+I5+aUT7Hi3BURJq2Il7S1V+13RUB
KHtJhyj3t5M2dJJzYDjhe+9UK1yzsKLU0gNadSntLjY9jTjP0XvwlpU1mImkXtN1
PDAQ7PBrNN5bHIEiPijeaQVMiNZLNuVhWfeGZWyd88pD1PSOKQ5jKy1m85RRWfKW
wc0ACcXfhtqucHuG/IDXRUq6Or7j7kX7Tni7rjcedWbG/ZBk1axFsoYEmzt8UMeA
3X3yfBtommZuM6GrSUnXSEu+m0ZiVAwMpsZTmytPCcGtb/SD+m5sR8sJiWmlqzIH
oIi0LoXklVK3VkYHCpMsJbBp2KtA/z7wu239nP/YkL9F/vMvKFYMtk586mUqyyrL
BCicY2mn6ccg7Gld4Ylmhl8BoVHBQy61urbjGvofNHubtxpbPTDvldVBqP27926k
YdYGsY9zlZNxFCwwWSoZ+eCk7He6JfIc0kslK3wP1WwzWBk5Yma3FRCVednyl8Zq
YdTgX8GyF4dZAcpZfsAIe2lq6CC7i8VG4T9ujAvRYGAhPEFevw+0O1xbD6SgR0PT
ZmfaNeE6WLjV84z3StLbXFFWpXnjk54PDO5MsXRsbWoi8MjmxJQA72032u+mxhVA
oJaEF6J6ll0SEk5PdciV82l0k35SUQzdPDm019MGVtVsqzqiJXehoN2QlzShUKtU
otl/DHGqdB16HsRflROWQlMASyP9oVX3XTs3p+ZE69gXp8Q1lhJQScDmIEx4Asj2
XyxatB+AKOnvy0GS47TzwhuErRDxGrdQ2sazyQZ5txtbN37aOgDQThpxnmfX3CMH
y2sur3AEkdnBvCMaR9QPixXA0Aa+WxyJFcmltFsyCokF9VzOAuFHXH7WTH38Y9FZ
fdzCxh/TcUGuOvtH/LDrwDOywjVoki0U9d5keUMUdYeSnueARswtqbL0gtvyGrzg
OVn32pv01OzuwuEVSNZ3XXYpMRaQW4BURQyI+thZa8MZBEqypFaWEyoLvLjv7RVa
M9XAJBtMXsMW7+ySrlQ00zYTQwkb1ZLQ2zSo4CKjWAbe5vvzULqkaXO+Qto0BHmV
5Dxb/G4QUVyVHMpVnwENBGT8ZRM6Z9wBVZwD0A7IA+8TEgRbCFBvFSPeh8BiWcsc
Rxz3koK5aAwnegybun3noKAB5A+O9OAAyQZ3hv2e1OMNFNQ5wpHNo3MfvmoGPjB8
z8Hyu5cEY+fp1vIef2Qk6kgMEJWi2Odum8KOrtEwyn3bmydz8fpKkUsDgSoODD2f
b7i2G5tqGyIaZIDL9X2JawyyODry/faWDENC+IlwNsiM5iNdmevkvZmxXLf14nQ0
eTUX4cFA/mJx8E+QakVZrl4HG7rrioJo2vEel3xm8zWJhPA5uIG95ZGrVfRiwQsA
Mdygxv/IUn3h07NSzsb89yuuGYVl/D2M/hIu+5BfsSb8k49nYsbo6ZoZBcf9K84O
PfNREWA9rSb16nM3poCRUyp2yQwPqRt7U1iiu4bYGgb+WSz9SeNA+PtAtUmxALjN
0kjlQnb6h/ehR+1PMc6HQyw58/I9ms9D06LaaxPO9v9MfFqmceRML2qAHnFPDFEL
JKAI7V/GaZcOOGVag7ZGgC8C9oxkCyvl3I/rFHMA6wugWAQXhL5v1Btyfq6c34pz
A6NSJ1dDd/TFLkdnB5w6j3DIGZx5/6HxEBluBST3FWGFW3fk5wJXTCwDrv3m2Ykk
Tdk78OGqNPp76qJygNLQuhHQ6bPhZxrHQAJJ3M/tl+9Ek3E3jlc81X7rrEWci8eP
IDiobQnsKA1zVpatt0r5oSeTd4V8ekMlZF6mI9NUe0o8rBUvXpUbwnvE7QvjPnOV
EMs7mLRq9GxjGiysJ1GAgZoghqJfhhRyfD4v9uSQ9SOgsUMpvgVHBWZTrkwIZTGe
vb6wJ1m1Hwabr/oby2w5P0HLuk4+5nzTB4wPnAI7got772uD0H3FRO3gP+wiQJTX
RbfAwUvebDyv/qxKLq16xmQE9hYwQ97IFq14Rx+UKu9eqNzeltbXdV2mXNk9OPmZ
ATN4gSYfHW2aDbNsOfJF05bg2sPF8yggLwiUWNGZHxyu/9QqSFH8Mx34KSPjTqkR
VgqGjhlP4shjvncDjqg3TOoEm34xQPbcVSKuYF/eR8eP6sEp8lZOh/BA3it+xrv1
t386I1OeYZrkqpcjd8y2sO4ULe/BZ9M5GJ3hPjB9H0bCrJtVyi9PYS5pMuNyvswO
uigxlDZop4ou7xpumjCNPLZ/4muAbAYZhDHFj7OUQKmGPT0USSm3thjMTrpCLfYu
sPo7WEw4D/D0MwM5vPiG00DUW45A96UZz9iCIm3itVAMDlEdu6Omk0R7nAoupw2i
PJ33D3FisGY9tMxXG6ZfPAw666Bcmmvp3KQN5heQOVJ4yJoRlYt3NoznOPmJi9Bj
A2jY3S7FQSd3NG+yxDr0hbmh9jAhNQQgouK4U8mjCINAOVSCV7gL30I8K+CO42nF
cUbcTjcIhDhWDjIMpwL9HbsXFA65Ub+Qs/IAG9E8JL2dfyAtZaLJ1G9yJvG7ahAS
hW3jA97uqs1s56dafQ+ES3bxRggJCtsj4FNb1DXVfgMW3iUIY7IzxKY+piE34i95
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 19632 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
/GMbQK29Y+AAYqzOrLs1aXtofNDQzja9NaCJV9U+TSbKpdTpng3gUBS73R8IpaY/
uJd6DxaKj4bR5fMutiyS0BCSrMoVDGC4TbfoIJwGJpg8i6RVbgZgg++6Sp8/ewCX
oCYLY+VTahpLpqfNDsIUsaI0p0D+cqcb5jALXavdSquBs0GZYTGokWA85RcNNSi0
+ceCszgl9GiqGbZOVjo4qTqh35nQb0vSyM036qHgB00RkUbFGtMNMDNBWeo5t+O1
DLSIEn9UZ/uL0jExJ62I6SfeOsd+Bq3U8oBF68jwtw1cTUjBSEHwBIiZNvVIRrLn
1c3hQAjtTtYpE99LzYpq9QwNeOYDPArsmKAihKY84bbWMvyWJISuHnsHxF/Ipv2Y
gWucmxm8MwPetHtTdFGSVJyydZwuC3EwWyPMZVy5vFSRDt5ma6Vy09aCK2FMB8ky
6JPzMHmIKvXwBcdyJCbSiwVm+W1g8xOBatI4F+FYH+XPxWMMzmmj0SXmc4vgUboY
xegVKx6FQCFqi33i3+SJCzNQDf12+W2pSvJOCSNBrOrTnWJ4VQU6CLLo+SQBXDFe
l9b+kqsLPPTF7LjrApsVhnZGWdMuBMB88GCWzhqUJNiBMWk6gR+WP62zQUJJaeiO
WP/G8pYKDzJYhM2sccz7Dyc6NVsDkLgDfLNO6U8DoNtxIz0E40cQ31ALSScB0qVp
SDQpDArkS51CsUToGG4QtRtwcnOD35LH5DFd2X7rn+0donE/A2ZeNIfQ4S5HFFCl
h6nfM57kuMQCNb5uaQCuEZcYHg8f+ZMuSEEqqDyFynwV5pjGPpTpt846NxzIcXWe
MRxvyleVKSUcAPlYhiuMkCetsr28OeJSOvsPMk5n6oKB8OpZs7Z5fCUqFr7C/b7l
74LG1IHi4dNVENt5mJBOBWy7F1Un9FuaE4FD/Od+HqagYuf1nWJMqOEU8e1Qteqp
rR+Chi/H5lv/p5sQWAkcB1Vu7t/SVQVcItpuDornmtEjUssknRdQIvV+gbkI+y/D
9zDNpPmtj90EqPEs577a29VVFnm+nNFRmf22eDub8VuTpWOdWwepaoAKf9S95giO
BCsxrvq8aun71U1xT7dF2Kkx3P3/hPYhdDhCywlbC3pYjOeSotI8wtLBzx4H5bvx
AdH6DNN3Er8BDkFqmN4+ntXNmfIOmLj+T/9i/sjTtEZiAfg9ZspBkGY1IfLj2RmY
Bq+2gM/ptI2BVsMC3TRA7RiYCbKxo1HBN3bzUbE2HCJrs33F12zv9aCU/hhwMqhl
mAyL530EFlZAeteVbXCHGzElKfTzvpum9OLmw2smfhBiOveCtp6WBggr3E/QGoCU
pBeyu0f+XYxyxX7WFEqFtRdvMgR1OUGI1J+C1O92bOxoCyxJxS9wFoPRLZXkkilF
NYSQb3FCQNJn6Y1MYPLL+9ZXXqvFVx3Euive7ZqdSF0VkUfRQNZ9A6qu4UeiO8+7
YIBxDY0DobsCH6yopyzYOVReg4whWd+Y+6UPyvCOBjekqVE3kWnhwC4pA/LlfFVn
n1coRUHbIwy4XjJpBsDx8V5Bt95tjH75jOEkL+Sb9VXTz5VePC+Lxb2tdAgLu8Lb
VP6iW32Ve2DAgD5jzleOMBFTCSzYc5jfpgLD4LKFn6EYGjVIWmjTgOJuTh3LYo/5
DVVKlfj/Owi9iTHkj17mUuAxTEgZDzHk0elwsT10NusNflmEqI+6LuR/LnsUqNTD
dXLIKMqUx/ombgribmCsjkUCLhq2v8UcUklYkjzR+6dcMpakDP1XiqJ4Te13pi6B
jM3FDm3valgoMb29GGVzjfN2CQ/T/Juw0gCFO0MHW7xFbZ2WhiSWXCCC//r0X2tn
Fb2lf+dr7dWfz427AK4L8GSPpuTY9I/4x6AMA4+hnzSVOpxCQMRZtOfOKf5qRepo
9/uOCOccZuK+vjA7fM6DYO7tieSVGoRtNlKMhbyE2UdcC3MfZCgzgFwJQ4wjqGiF
7OVaam6FxS0m5XxPMmqFJ6Rl5e6vxlNp8mcP+LwsgdHt0biUrXZHwqB/wMQfTgZl
MAPib4HR9cYuS1ueXqobD8Q4DAgvhCyRF4WlqIOXdCS8gFnHdzHAAi8RMR6qvcWt
JnsWtdeXoN9i2LSzrdsOhbEcckEnEkLLcTzmarayLiRw+694ryXwvyx7IY6Glyj9
OOnFSYy3QEvu9QTzufoncqF2389TprfN0j7IpCOK1pSKErDP7qHQG5rYHcCtry6N
ChqArJgOQ7lc4nYbrsPTtAkHKTFWpPcFzLu/5xm9It80AB9liookw+Sz9l7LvXT0
5KsCrFDQLgAzwqV9Ue6Kh4FTxy6x6coLfxz48bvHpOYbptu6QPvOGzcNt+1vsnXy
ZnnS3/98Gs6zlpWpqAkvM8KJM+hUxRuFz9K0HbauhSGuYCOKlmKngWz/CuQfv+Qk
to7+S82corWJgC3ppKzDLAt6BjbYYN0Ns6117ae1mQSq0jEfVQ7kRFxt2MJsTZsb
gcb+gDPF1TKo/7oJMzlZ45HBtdcvNuyjeywlcMkZgJ6JX2L1wwKqGvfAjABLiLoa
AnzAWwKupP4mB6O3+HhP+PclQ9cd9rqbm9VLIsLKUJgLmyFUcUAk0oE32wwTSKgo
xtv7Y5ATPuvYNpzG8WrscXyXuu8cdHIyQI/lUdgLIXHfuLcgDwou01Y+TM8U3w5U
nPW73BqiMVmcf8yi5WbuH0+ZpKmZWBjKefoJdSOGhnXAEe4aEVDFyTo8rXbNS0zU
2LfZU5uIiEtVh6y0ycED37Y6Kwnbc30Zt8en7qRKfKsUx/Jc032sWJGntepJQMCM
Fw/ezw9tzClyh0Xv58ACW3jSduIlkVFz89owu9jwMqUos4G6noX1+5q7AiBIxw8g
bkhkjG8cRG948rBQuzn7fe91s54dR8188rGJJ8BprDMFVN+SVRctQtiXRuK4R3Gl
ZG1KtOI6xXZhsMBog6yQ44oIlz3J71fLu3ei7vvMb7MXkY6msydQ7kGuGxDaiEpZ
6QhM8yqN2qMO8PN8JLD9ys8+djw1axMlLP37dI42BWeyVUSjhXQoH0UPTcw2McdS
CmY/b7Ac/8TMvjeNO96s9ero2LLvHdmAjclBDNc1WTD8tygAJeYibcoNvPnCPuXO
kvIK/s/xW1CcM6i8Ehh6MB974eCU3lhKKgM42Tzuewf378XvBX4Q+i/yNQ3sLyI5
EzE01uLLou0lD2XtZxyHsybabErAQL8F9cWKHoiz/n46TQoWfbe4xqUiKnUPmYIW
epNVr861NRdNPTsEvc88jPkBzYaTcjpV+3UP54OqLoiHaLPqPzS/IEdiWYr3kx/Z
m8VQHRDbjRz/UyB5fqLUeu3cAHvfb+FXGsAULDk7ML29QevAQDUPX934kMHDf3yg
qq91wAxGJDDlHaeucal0xKXFQRaOPTWKaLPrCiBvXWAOkdYrZk7yh+C7g7wlHTkO
p151D3znyv7YwOeS0flynbuBECbjj0Jk0ZhNE2eU5hTPs5zjBm8rJJL83dETRDln
7lHV19Xvoq8XRmTDeadX3D9BA+Vbo4UAznQw/3T7K3PQjrXkf9dU64QNy+VDDo7w
I5fALkqFvIHtYZI6JmjrOICnWwzo00QAgFpLfAWRoCBgZp0fqFpbCHriOcsRC0/5
/4O8qDZ2Q/s6m6Slc1jqgerLtaTpT2KYyrP4DtbNrGxjbm608xuIusEx2PdUbz/M
ctt4PnmyHVbRyDxYPx89q728aS6/icJCt0NiSVaxzqKb2DUh2cdjGDlb5GEurszh
lp+u5I5Emhz+uIhUA91CWNdGFoiFerofzJXUs8tjlbrJRku/t0Yi3WKy4ouCpQa2
eDNRzh66VqxT6UR38KwNboZBiZUXEelVI2qJhNMfvpdlW3tDtIh5EvdVant6UvOJ
FSWIdXv3P8z4NT14TYF4t5D/d/RcynQYqbYRNdQeCtoMuT+Fi4Lt1RjANiJlhUDO
7TGoDwwfddYMCqWitPt2UdNDNltdscB4xf4LJxnLFMhr2f+Q6KFa8eZjnQnjPTy0
t6d5VLCMyl/cVSWm7WaFxsT4XRBJnIZDd9e9vml5TQnR2G0xl+C1rqYA/LQ24YIV
31sSzBcTkQekX73Duz7SHftKVAISSmBBrFwlT+8wp1c4COjDkaKR/ZjtBxDPk21l
MlYXH8gkH1l7Lw/oCxKgC9A7tgYwEh0lwwc5hAFxt9fBlr88s78Erb/uEg48AFMB
i+AY1tzfpweTEnZDMTgAaa7bkdktSSMJxZ+Gmgjh6EnOKWBIe3UspLVeIviQWcTD
dTZNp2aF+NKhOQmBh9z7SUVJFGn7YPDFMhnf6EdprRnXeBDubcBYykUACii1u9HV
2boh6wH/y33xTMLISzvn8bRnCEjhQmw471czIEZIHAmwXXouFAhYPD07RlSt5HZA
rQTHvrot3icIftiIzOd/FRuDJfjokrJbe8+w2h9j703j47Fz9vYbFB8RXQGQKCHp
RVYigqkmq29IVUj7OO9bnZtqy0LTc57frZvbp/wFJrEqPYWeLSp3B3TvJjcf688p
jP5kIJ/88IMDquoGfrXfXMRvf3p5nXqL9vkyxZSiV/h/K02a7ZMO8wm5egi34FCb
riH/T5pIyYdGqbYI614TSHzAV52HCJ+spNm9pfrJEmQsfsgt/3NUKTah/AXXNKzu
1W7+SKKhrBrfjE8MFC5xKg2CfYsZBopIbnu2gE5dOlBD11cBhzYgaZHT/ECa5cJ3
h2m3dkx2++w+SoLUi4y6SZe6zXuXiXPsO2I+hr7lj/2JO+u5wAZcmh+bCo3U4rup
GI2iGIrUelWa89i7xYFnju8Ui/pv1Mj+dF22JoyNfzvk1G/BG6x6dE3PbXCgoADI
4+DbF07xqdve8wOELEfsqjh93bhKDizaTz0p/RiNyECSBD+4oIN9lkpFqF5ze+yA
XtQcRSVLWTskTKAMwEA9G9u2IqtL5Pv65IT/XpM4tPHHgUAzQ4devvw25JyVoXOv
X39tjdlwBxOb+PeuR49IQLBOYrdS0ANRwacz21P12WkIHxdhkgUU/V5piQis3Fmg
AcDcUvh2CFk6lSUQTgJTNfRPECyE5Ln86QVGW2wCieHdPNdJl1dUKvIoKqryfTQU
oQXkjii3iS1JOjd4s2nAGF38uvjdjT3pKsrzrnzRLiPUaAzVEvWTAWlGBpenRriP
yK31pbh835zxNStAHXTvkh6gX/nvviqdmv0aomoQgcUG3eZVKPBp052BpZwktu1R
9PLPz7/wK7UKNyYh7xZM2O7peBPDYmAnes7/CRbnaF7gR3BSSKAtBknLgeTmIXd2
LJYTpdRvbf36n78Qje8rn3bwvqfTwgExIvFyTYircoDIEkt90GLDdYf1anQc3ZsA
QJTN9niEUxglM9tgmLuEhNMexnREUkvOHweVNcC61oWfZfXqkcrIEqjCzcvZ2Jdo
e+xNRrRmIcyZmQVrG4Q83HIA3Mi9QYCzowSs9utmR+m+zejKI2y5kol1qbOhvUjO
I+kXQ/8gKtHQ1ixk+wqxNuyw/QsAu18VJOFmKli8/oB+xDcapXbbI2XDFYe+eTwS
t/+uwCGxcmHzYSDC/UDt9O7MThSogy6KOZbtxyYvZc9kSZsKOAawN7gSFaPfFrua
9Ht0Vz+ZQ+ancpuyATiY4fWpmnJT6TtiyIZejrD/XUJi0g719mh2tKmIHSSpgbiL
UZYo7pnR+jyO3Qnih2qXJ9dVh+FcVafbLnBgNUn6r4FPvt1apqSFT46nAqmVqEGg
DFc+WaxhJdSR/dWQ9A81AUEKsNir97bsG8sz8ao+jUxv/3Bhp/T57a2RwbOAN1ow
SHtlwN8oTfKm3v2XhnZouI+kts54sBGL9xa86gwS9bxl0meolEwoQ6KTuPFaCwW9
yRyh9l87xk9+dgZSTF+jrMzPot+2XeoYqR8Wo5O/zwtoKjzdm5sLhcXPkEId95DO
52h5uz20zmhhbY1SuYnlO4wnPxuCDtVIiXN0mb71aygLbxHLAgwirp1nVCyYkpv3
MyDP4jZjlyk1i/VGxSW1IKCiOTgdXUN9mDDIGB1s7q+7QFk4PPy2G8scWKYuNAqw
f6350XuOesnBQSKvmaE0eS+eWUscaBh1llbJFtordPsFL9nIBdOUwXVWNZAVZxxK
kqA2fOK7zGVbssnGGH4GFddpEewWvPBxdGGSm9S3jG8y36aHgL6CnuxSBh5cWHh3
iVLD2eWUYrAKbZltY9WoFRb5s/QrX+yeI4k6w3HS4KnkB0Pq5KXiwSa9ll/lM2+t
GqAW0htf/Hzn58ORj5QzbbW4H7VkM/c3RbKM4M3mRUGx9FBdBEWiu8UJ1oturDGK
fMylQaLHrfCCfaE0WCJA+7gysqY8vmAsV1p09CYO/7CuNDGpomj5ZThHEpSE8Ejx
X4Fmz/VdaSYih8Da4wG1XfJbEg4/0yVw1ag3m/tCnMvOylFIbrZjq9zK8wUns99z
mhH3Nu90KJpws073eTtcFVF6sCQiD7Q4brdxOvzCPhQDg6R895afhbLflD9SJ39R
/c2ADSgQdA1YwHxDhjfEm5n5bkC0puco6DR521RZ75RWPtTWPfVewjNsBRyOD1vY
1eMP3JtRC/8G7nBcD5iWw7WWsxOUOhEU0mrDjzj4y3R6TQQapqtWcOoBvKpPe+WR
qX0rEQ4Y6AL57tA5qe16S6N1TDaGy4Bz/TdgeGepMFG7cpYoQIUZcAdKa8YlvKeQ
20q60tCtX9O/lYovJ8O66PeJwT5JGbwx5yaExrtB0iPjjOB8VP3/AMbJiC7mkNPL
InxvsapxRXx9D8jeFZPhp9lLdF0hVDfoeF+JPGCZgCcqX52y5cEO92jmwSSaOB10
IsSimRx8uXYJdjCzLXZUwmVxb9zFhl0roPRSzuS18xVVOiiUG7AT/ao5pQksa1JZ
AtyBoKiCG1NoXoy4budSH44lIuYK5EdDFkwDo1EjlG7nMa3d3vWGgUGK3Trmp0qP
CPKQYaFdYsBddQgg8bdTsRzkJsEyv/2rrj8wm1SWiC6YMOuwm859kd3yycivwOBr
H14cLmmJkwUXGC/H0PaHKBi2lvsbqMdPzGLE3FQcRd1WKRuiul/xp7EaV7h5O+s0
RTuIrNo5h2WSLBTJFcdv5KjL5i6I+jVKZ7nJzprcsASPhmMIoW8abQrl5uymtNib
o2KdPnpLFGlK1l/yHzGrzvfOy7H8WqD8r8t0Wg9kC5SjFaqw8T/8mJIi8pPy5nC4
5vWqlk6ergIup3u5HJ8fLtsunFBSQBSbzq+Dc1zUxIREvlEQbBuSr9iZMfac1vR9
g6VSmjH7nZ2yvMtmtpoqnRH31CViK6vvjdH04OW7Woc1fZB1Umq3V83uB/fTwjhb
qAtiFYL6tfblnVO0VY0eJov+n0jiLKfm23tCOdV2g0U4+p/5VZG1jBffO83WOaba
x0e/5EKwYzjO20aL23qBt0fssuq5snqbzmkAz08MYz7oTAgROM7HT1hzCsXeN7eu
NdsdFKxPPY1JcLTGuqP3TqufPwCti4xzv/fEvO8ibq0pP33GUyO1WDi9ziC3vWoa
0eWlUNd+n8n8qtdGT9DpKUf4XkSrWxBgS2oahcIhIQGgBcvtnDwJ24N/r3PuI60T
eOQ16sIQgiGlYuVwFGpK4eJ29ui1WA9olFfVYv1ek8CHkRF6spxSvLwUQwwHcwuv
B+IPbGXB2Lx6sbueW4gfEzAydMqw160RfYSKOXFpyCxl2q7rSZW1Buj7wAA0MyXu
pWvISdPNkcG5gmInEl6y1q7iveb9MK9iHi8KGoYIrrktPnRQ27ZNpNMz4s71SY68
priBTiTZrBsxCQQql9o6qYQ3XlUP9YsSseCLAYWKEOTgctqSPtTjgHlA9ZUoRN0w
pXWNwh31c9IBxRVIYIvBaS0E3V2RfPt9gucLPavyF0hatsL4tM0khOLkrKLBmvFA
L9dw1auCFKMgwKWOgPu6Dma5G4fiVuzL51AqIIBoUOqxrKhsJJect4U2YuHVHgOv
hVnQjvQcFn3du6w2fM0oTDfxXjp58rlWEd5/GiVsGs/49VdMBUqME3L12fI2zP6Q
hNBPbgzUEc7X9Ut9FVREeEbe9FRTb6eQjKEvJHqjT2BsFHwoWKXpiONfzOTa5x2s
irnks3cHyJP+8GGfRQKMr+y2Xfy4aTo+Ma83SsHa1JdkC09LYffLkMLt3CymEbel
tFvOqK7FEgAR1oW++dpEZc1MfiCgA3RX3dDP7s9JNFfbcuZLHxmiYCfjjyAoA7Hd
Ek9zZTCLqJGKrOeq11kPYDqWJzg3jMoD2CBPAqTZCKvm/lnIUxDdsqjbkquF8MlW
oiBqJXi2YNZx+AnglG7NU2uOEKeABR2jpJhL/Fn7NV+0dHjqUz5qGPl4ShTjhBww
wHjPm9yX9vtaNFs77POjrcTX+wjMYwdN18FUsehxL8r4LMlNyocY5X29+oo7Akz3
e3w6tuLaNwzXW8oIQgRH6u7AXmLcSxM1x2VO/5GD32zUo7iA/P6srnr1QGbNiyC/
Y4ej4VYX9UA6Z4Zb5HVLybbGdJQ4KjeVin1JOCF0wueAhLwIEtRKQswDt80aKQ3l
100Ri7ElbETD57xBOztjOmyQrev3YueC3qgPNs6HcCJx4PmFgDNhabMWHkDeI252
nnjqkOvibaIpMEjc8BsG3RLmFsn/iSdn3mdswoYlsVmcgmqVKrFjmpiPb38VCrWv
/OoKoA4pupIDCqWJ6dsnppmfBZHMhSdDb5saassqbrGjhw+rIQNKLF2NRhrad/Np
760InpNzQ9q6N8O+T+/kauzb+2c3vi0Obbrf5fjPIM5IZbkYk/IxtNL3g7Tzp9tQ
W249B2T24Y4vRmyvQq1DH5AXtX5R/LEFONGKJQc0AMSEQsR14PIlxnZaJfLxlETC
4Q0KtKbYrrXdlml2HpiiMU7EvyPts47TMOAaEZrSpiFtjnt27yKrngovBva2u18T
02WLBasPaSieGx+13WMlJVDNKEqEok8DQ2MmZH7ypEYc7aYBJEOr+jfODlxp4T7d
5LniRMlbQv2s752Cdrx2/kJxfd7wX2GMZ+tS2l/GHZMJB6yJwCy7+j7FYPVS+A29
GqiEBvLza1tzN8mtlmS+XjQIpqTsTnAU9HT6RqS6X33nig9gVgmFykeeOFACOCOC
ZgWdnlpzdvV0iVFhFWs+OHNz/tP/MyWPWVdx3fKatyKISMHED0pCL+ZtjBfkjHiB
Fmj1LwvtRrnWtVkKacZFwsOyB5xs/saOvU9CT/k7QtYEOT5qgaZF0nTarGkbMePL
bG+BXHzVHfV9R4kFMtpNbU/Te0xZO9/+/nQzmFx2+IdlEwkUBzdKFKYxHhRlfhtM
02XfieDkTaP7F5GNmHgNODZtxEqUVPGdEn78ttwFAzeO7U4aMcvTUT98dIQ8N1zI
YFR81+B0dI2uC7m105coojZi2AuSnKoHPVn1/0uIKGi0AxgPx6GH3vSRBV4XOL5T
wskq2chq//wHvHo+JpYGBbHMKef3q886zaLPBaXEs7gYlOOCHcvldSPD6kvde4XW
LStC3hDup9LH5U3X0JUVLZHVIKrmLJqU3u/FXr9zgU1VApi7+OhztAKWzBpzy1ys
9Rao9i2gjIFrr8NR9uO+W52v8IUe7FocO+J94rz5/I7kI6rww4sQaN+M0kEpZbg4
3/bYibaJ47GCAkw+JAHSLSyta01g8lg9F6RxgK2CNeqJHfhGcZOrSE+sZyKxH1wV
x5UUfQ+33nopChaiNz12fpYinrKf7hJ1kDen19RqQASdwPmOODVvMEPrJKYRSno4
Hxh9tIsl8zx+Xv2hMMhQoS0aQOg0RRmN7Ab7hYw16tsLF0Vt2qtbMVT8ymsQZG+O
JnT4ntJmnFuAKi3/YYx10PmQlXxdVNRd2ujVwt2I2SxaBd75CPw8V+8+YAuvNzWU
aPrbj+oW69VvPLCx+dLPkr3F2GA+1Qses3jh0DHwJ5A77yOecBI+e/3kq3ZTAJ8Y
wMpGIq+ukO1Sab/1y3yuverHZT4o3LejbIYcS7gADhAbcKZP/Zbdg+HQAq/QobJ+
emY6KukRZfgkX1mOLNWWlDJYBR8hL14ZspkRuLmVu6u8WR/X+RXnhWCiJ0l3bYHS
rXCWTVA41k+HeaCPupXVrUznbjnMt9/jcgjqks6bDWHUMui9UZtHs1LFl98y15uB
iV5LQ8HfVfBNIYv54bOWpliE9XkBr9ulp2h0xfQL8Lw6lL+dlodyHgYpF3pODSNA
Z8PR72HaCRSc1DtmCU214GFnw+lb3ciLDa6Xleo7d4jxXxWk2jZ2i9zjjnG+uwCp
aPpAFepL1JRlDNa3i0Ce3Z9jic/1aNTHjztSMDc1QX5Y0mp7c0rzUdKtjQ9wV+9m
d7+B5UqoQ9PZQakqmigVDDm3O6qnT+cdcDrHUIr1PmUAPFs9wqxGumfqP5ihVlWk
yGdx3OpnOFM/p5tOc+pW2chsUBNyi++QzV2LA+JAklVCE4WWgji8aICp/pXD5/y6
hQjaQ6XckVrin3QrW4ze42oe1+vFtvwPnduF0c8/c7LaHzRjGjx/STT+wcbz8EdC
Pf4NnkQ6yhy94gPUvbkTpmV8wORcTKE4RYMYRPD83Go/YM04ntLKuBjpdQVjj3G3
B4lUiMhjcq+C2iI4/jI3KWeioYXrSk/SXGcYzMOtUOBOasoy4fNYcRXwAJq2Qj2S
zNrZbJML3992MFzJp6X8farYewfjGd8X9rGCfCGrFcdG6+jH/OgXTG1Ofdh/HP9i
b07iE/NtM3Z8bPYlMGANvp9C/lsUicSiO5I4E6TDblZn1RccXNnFvm3yka2bp0Ik
DtqbdollxCjZqB8npgZC7O85pMyscRlRQTXM7trgXsW5Er7OAlcgzRItvM3n8i/N
yiUETRXLKlm2oK3nwHxHJ1zToVg/bSfi2/27ahKAmEnHLnUj1LlzjUsrXDanXP8u
Kg9gTbfTrIj3fn8P2Z41x4nMKLls1ZFHTlPRtag2Nzpioqb5BWD+26bBGTw0Mkfu
oK8DXv1qJqcJ1Mo1wvlDgy7tzsuA4bWHMHVN89W8O/9+VT5W25LcLdXS6wjFNhw9
HtF22QcmvdqLC6t9/YEC/XvImwdruYUlpvG9w1UBWLAGdNH2gKESOTz1tPAzCI/d
VMOolQY/i/mNpA3VVFYW2uC/aRnpIhob2fqCGRC0hdBjOVteHvGXvoRY4W4cTKDP
TxQxaQAPUaLJ8C4DC1zMBwNm2dfeKV4aB5Ktvhx0f73MVud7h8+3lbJvUQxJfWa0
Va4anf7/f++7/NstafZKaf7Fj7yJsA1wHafauWAMLJ2jMOqZY5I9DdQ7WkuUxXdC
aDV1U2U1njyKSJ471J+t/z7zAMTfC8rRmBFMeM9wYcILepRol8usQ9pecxbPG+Oi
V1RGfXS1JhHYD6+yX/VQJGze6AxMC12Ld2TEIlZMPAPa+s9i4UFc29wnrcTel4vd
CJSkGbHlHl0iLfAxctfzabmilPi+N+WcqlqyqYITItKiLMrYTHOSx86cGgfZ/VNs
cJQl4GkrcKB2A2BtGOwhfLLLVSWgcOgjUO13C77cpiY6/6nsPPqawqof7jnKSFcS
U0QRF72zP1vntx1uVSuB16BCV06r07vKsF79wBCu+K97/afrkzh2jKSznte+xxcg
nMD/4XTYxaSF7piOnaHuJaBYyIwcJ914ZHL8+ef5xPAGhQf+s5oJ40VEsBaI7HS0
V+FhGYd8+8xxQdDA8cg/J+0ftz7HkHP0IxfRNlRts+/LqPVdc6WEV7U1eVjn5mIJ
MhRiCIfePVr8f86REORdcfqPD2L87kIl3Rbl/23s5B+9BiCk9yqWyDknAZKs0cxf
dBDX0eu2kFgrs0f+iHFzNoTibYkw1P14KcLnkaeYKMh6aTkOR2RBDDjG5fBZzheV
BILMY7eC+9uPMm5XkVm4NkHwM2WVcXMrBxSLMWVSKucmlyXFH3fcJ6qeXDN2Xy0r
jLhM7rF4nUx9vVE0Mbbi+AkR1iqrZDxVl9gM9+CAlxv/oSEMNQml6LBgxdNGE31d
ybn/PyJFRA96YzdwgK+xR409Y7sAjMn3WqPSXQJhGB+BUPp+xKjnxPWlgYAoobYf
dIVmyL7mIfzka75tkEHRoHg1bXd8yh0RA+niGJKpohxsU9XkvSvOzVhIfSb7mRPL
AvmtejG8PdUXbCJRwMPVb4EFs3WqgWddMIfT7fGqXJVXCF9PbBJe/Qbvp0AHBeDP
r2Raz+VA5Q+LPdokwKrHf3ZDB0fdfBMCQT5xiqARX5ljzPS2r+780qy5vN78x11x
VR+SuSK0nThISxvcGPKMiVTw2Rt1S373eFsjRTwItqugqscdZs8NShan2XG4bBry
m/rCFmArsv7fdxeJXBNL0nlpqGsMrd8piLl65flEAFl6tn30yNTaMagVrE9V3cRL
Wfv4I1TuEdA+kF0oqFc9yH96cHj6reWFr/VUVwzoC+shbW3w2MtafRiX5PFp2Wdr
SyD4x3zMPEyP6F24YtvwXM7rIdmgm61HNHd02fXgAeBUYMEw9wdrguFQXR2F/pEY
KyRoahNUj/mf92J4a1nG1A+on7+b91bmsoA6hLGy7MolONlI9YEDyNNn5ic11yxT
g5yk1/AZ8uFKWI5Gl9+YfbRWdViBbSkrJCapIPyZkXHt2+fviEsgow34dl1b6m+K
UAetZQ6ZzR9/Ru7OMWUhmbR5gYCLrrDvWkxbXonioqFXV3TJIcUraM5i6zihg4oT
M7Z3J86sreXA4DHLymztTFiCJbEmPQr0lSBvIXfwCgy7r5UXn4m5ieBi9FfhM4FH
HCjUaG3Nyf46UM6tT+8Cxdc4i/SZXFqz/xUR0FZsKDTX9XRJlzl1HGXCSdZf/16x
l7ZcRQizAIB+mEw2tYBdbpkfLigtbTD49Z9L3rkvqo8MMe6TjmkNeGaasW1c3HKl
Kdb0+ooadkYeRyJiC7dXvJ3hl91E9THDy0KDweD4DldzowvgDvGBAHsZgG6FzcfH
Zpi6Sulbwek0p23awaL2F+OgxEBN0csSHNNGyO4Mn51lPup44bnHGG4JlIy6l9Of
pB/rq0qghOjANKwqOSzqvyb+dyg1Z22yEHHjaNY2f+imvq2ZKoF5D9CVaZhCUZAG
vtXuAdHxDROFKk7bJ5tfT0Zxl9RSckZUhKnVkVlFyGJBrOWa5Q6tMCLfU1Yb8fKf
uk029IWEWyU6AGILmpvhQ5NIQWEEvgsbI+enybKax9jIvaaWn0cxNrvG1miyCCI8
FkER51Mez4xBfa15iAKNTV9xBW6+yuLVKYiymNQirNqDAreTq4lZI6b128PX/e8s
5X+mFTYmXfb8COdHJvF19bCw1iWt7vufk86MdyLrZ2xeuVFC1OunLNxnOTMrfnWZ
UzxNoka+oWN2mMlwUM3MdJiS8WK3phgzvUZY63boj9nJ/LLFCwrJpfANO2F2XWlL
kM6e69mzysJ/n83M3LG4B8r17thzd4cny/qPKhj+wfmo+IJi7zI9aUYCNfol1w8z
j+zzZxcaK4DISVD1MX71PCuYpwzIAZraxxbXKU/AYcEZGJxHSoDImyhTB5xEgrg0
qP4WI7FURfZj3JqwsWdkNsevIpIyA7zLGo7zynrhgw8x27Z+8CsAesVy/nIRK8Ok
xQYfs96RZSqKOCDyL/NdoLu8qUST/QvAlRWpwY/+qyYtIHYZ1FQr/Epk7qUpvSc+
KoHQ001gmel2vjRmxaAfbUO+Abmkpg5kPGYxwovIO9NHB595AsDjAn2pONFIy//1
tAjK6QMzOqtNMxOFRR+DCThzjlnmSi532YCaEozVUU5AXPZmnl1IA1xkjbmEzxLW
ikWPz3Xzltsb1vAv20YuQMcSO3wUrlHw3TqFkt2TaB/4cRgOnBgmNZKcBtK5kzPO
nzCbBGTD6/Byuc3ADEHwEuh4SJOFskd56BxLSWbZrJvHHjraE33rJ/Lrv/Jms1a3
LXZyrZV8zyGp4/nrZNVPYhRZ+77FtX2EtjHVu9TrNeR/nqmcoL4eAM4DNba3ggdO
+U53ibzJrvuhcX0gHbb3sgLQL8KLaoNzNyh/04QkCSNaU11XLeTaNdoGhaEOIA2+
jyREEOrpAGJB96zs5lWe1FVxWHzBGSpkI27BT7gOEqHZOSuKbFpRYK4G5Y7a1Tor
uQkI57qidRQ7BN3V28svIqYx95N1fwo6FxpbZjHmXR7TM+QTeLyEisEG6YVIsDA2
egTJgYcS869Ikuroc52YKxqaWCq6D7KWcs24hTU/Z1pT01CnByie80wJOotdz6ro
9WHKFVwpwVv5p+X6mjA2o3LtFw8NZGlMT0arJ1TQ/9pYjqzipNInyD4OAUAglCje
EH4D034f6oz/v69kzFY1DXSuiKee6A7tC2/jX4dEs2P65eqSVRhEyKUIOZW2sjuK
+mObgSLcgb6IBTvfbsIb4cqt/E6xexKlm76e3ZiAjuslbgAAKwLtqci5laQ8qjQO
YeBvzIps+66JYE+HuGxW2bD5Np5pp1GbFgkYOm8/uxY7uIULVQH/fYcpeBbSjVt5
OKdMyJ7b/xYTghmNEEXEBTfmNYTMqbztNQkvZtb7mFbxu89o6PCvTIsTOFYwb/Vy
9BogpGP91bsSmsWvFH87ctel2gc6zopHTE8SsPiqfHtXZMiECmiymgFwimcgwEpc
UHRWXUqqf2dvHcsxizlC5oezSkoHN5GiWlUwoA99hJiilwDSpFTpXArpo4jO6ipE
9nr9jPachZVAo5VWA0ifj8CMtsEcfERir2ir4XrtpxArXZFtgnNt0y2hJg5HOstv
VdgVOUMKgijYzL3CxvYJP2nPRfCZhEEeHbh/YlwjFEID6NpGT8sSnlgjFvpLg+jG
3m1828epUFxPQ86GWIzssDZckOkwew7nrAhGNWqOb0on5Xj8QDM8BP2M+B2rEaaT
pQdYL15eMwa+hnE7kZi6kDeGHkatDLvK//ncHeELEUH+TlEIrBCdmZdZB0XoEt3L
vuP2FXQWRmjZk84v2hdn23g+25tvIS5MyIcT93XCigsytcMY/FTQ0JhORfJCHNV6
eydvszMNdhgNqpy6sMUnfvlmehkiLD4MwWKyqCBSoJwJJ5oqbub05ZZQ5F+DPkK9
DApGPYYq3sWFK0RnHD7r3FhiLeKtehKQx+fkSnMfRuwBI9m5jRhn+NJvgKsPj6r3
VOMqDngbIhq2or8u8DVNHTBqNDSh348E0GARZVkAJbMKlvEJUotM19E0WEKAxgWY
3tmJRrUKpHzCsKqfGNI7w5W9otAchQgUySkN/dGAv1RppN602PyksT0Q5rCx++f5
5fvGSxWLtVIWdpBQCsvJDbi8pnp6MTUnM+b67ut7b52UZp+dmh5OwkabKkiBPcIn
+Ki4GsX8QV2TqpO2K3sgtsEOTpVrNpw8piqNba8KnCLR5k4TnekWggDbxVD0Iihi
3y2rRr9HvW+EBI3APJpN3/xblN0PA/F7FuEWTqtQGjssbC0OQlBRBI5/tSl64HkZ
BAdJouq5aG3H+3H980VH/Qld6GG+fbuHTtUL0t1Nj90TJIY1Xg5kJubla/HoQIZJ
m0bXnF+QS019KoV78iIGzhIRZEkiyp4cbUSyXU13jKm8iCtKdKFSAY6Ajb+29Qut
1/Wl8RzFwm9i8Tn+O5sqaSeSwzofAcf7onfFiSzZJxurIJHEQpPf47nlYZCqFNca
kAZygFyTNWsKhFFbmjq1DXv656FPh1jAww8ISjbBUN9pCTl22vVqqN/MK9UfJwIy
hD3gxlmQHh9aisUBLZ+Z4PDZkcsNRWT8DYjGXUCoGNo+nqnP49HqlKLl8c6kLAPY
m3xehOMvVgiJ7XFXYyXHSN/dHaOLTGqxBhnFkYDlLZDKZO8pUEk6RhOMl8EFbfEb
zRPd3WUp39IK4jSYRPdJxKWmxOTou4qSQFe27cS1dKFPj3IiCUryH9LyI4kkcf/R
Zll0K6EIN8mgbCGn1xYzrxDNO8bZH8G183+AKUSp8i5NWYNyS9B4IyVwtIuSkI+o
qlW+HHRAt0pOD+WGFNvRwziA8zQMGjZC3dxNGtxWp4iENpWGiN2ff5fqhyocS4CG
5PgUuVU+wQcn7y4J3srFQXnYXZePr3p8eyeqnHOpWcGrCGA4ecEe6fgQ0tbw10HU
kxgx0pPlfr4y8v4/Ywm1t8xGPGoPByK/WETKYHZHzlaExfuUlW1OFQeHUbT3PrqW
ayH1+ynVNel+fEwRNNVkbG41Aw7Vrci36X4vPmYwfqKFRwtrzeQZTeGTRydupOza
/99YieU9Mm5hkoDU1eQLSLhM8nhRnUzysegBv7FvPzhoBMcebBz2DDzx9O1Yq5ny
STak8ZHc7mRQ16nZqqgG7VeIiwif04vRiRtUM+MYW8Sza8x5WE/Sf7dKF5iW6cO5
fJLvOEO1924hA1mpuPa+gksuBCTrvPbZpfmhKjOmbyPw+Mr9pYxlp5iMJHG5Dhj7
puIpQWLoy+FDA9EoTzTQ2EQnqdoCGOVHruGxQjQ2qMdkpoY7sHlzrxrdCoN0EZdA
BZH9zr62hHERjFmXQ21Kc2uJyNTK5Qsv8w0RKZlyIL0BeClB8ipvfQ1lRfrcSLEe
FXMTv9/ctbw4j3SQtR8POcn2c2q/6WFdofb+PsDNhEnBG+LpY3q02fUZ3QiS4BDK
PQrzJ/Nyk9Gc43Sgu5bftfklTlIfZq8czB7uIQ2+0NrHyMHSWe/RVtF3wDB6w+DK
0Pe5ualNr8CXorQdq5jdEhBls3uqq02hblbV4xvUpDGck1LwqaIn/8BFuYmdsNH/
/cGBwD2mz43GdZZaXwZfRLgvmi7GVzsiZrgWUWI1Xq3hDND2Z4R4mYzDEjLgvuJp
Bg5EQtzidna7c9FtP0xSzJZ4yZn+8kGYYpBlxDYMtBUazref9q+Opli5cXu3Zk20
Oe5BboYfM0wELsXBuZ97xG6xORYszGbzmR0DsfO6jFvxnX3bCbMJGwmi4P69HAca
u/1Ad7X6y7BGWlfHz6X480/KOegKvh/U/naKJkpQ7nZVf9c+SBakWDgi9oGnpRS4
xaj8jQnlwxzNvUO9ARJIHVUKVD5PRcCi5lGduiMtbf6vEiLkZAfNEBGDe8j4rALf
WVzmY8c56qrB6rkBhs8s9dOQurHCIHMmXz8ic2UT2sO1/lLvVnPRtT1UIkR1o4QE
hiutjgNk0FlVHn7sWLfTrndEBpcfUF+zgd745zj/ec5v339wYq2qXfpIMpkDeSjb
2k6a0LloO/sjGqaaIYeMyiY3s+Rf7vV+z9mkyGGWvlX9p3706ixAiAqokUYJ5vjO
d5viNt2dm2EaH+n1Oa+52O+AyrhG/U2kF3Z9Odi7qxLoGWWkXnevZDetFeS6GSIY
EoceNUrDNePRQNaSvum/vyl6oJZMu9x+tOSWbiKQyc313+6yy3sOlrPoT0zkVafS
zUSL7EeBspahlzM4G/FjqrHB3Rt+/nmMWsNYS/9SNEajiK1yIncnpUDpXIjMHgas
QjwmLuXeml5H3u5hlwvjI4htuZCYsbwLAePjy3J+gYeYSOC6ngSqh+ldh1zwVv/u
CLBqSScBOOncd/+02E2Tf+ZzcoaNISZWYV02eQjR0T8dgO72rWt/Vib22Sz7247Q
zh0H8oIRIviQ6HUTjxqgl51xKe/WnNqe66i0AyJmh6w2q/ftzlxWa6sMwvwceD/9
9QggEvIcHpXnR+lu6lU+adRO4fhIPLfbY0o2Hxwua+oO/E1AwxJTtIBvXDmTUH1C
LYOymj0Ud6aRfunTIq60eKxfLuu70RQX14Bce/8i+T97/Cabi9XGi9hXXIgL2KXH
68w/H/Wb0VVrz7tm0lbh/IzPeETWPdqLUa+T5CVQgzRFLfcBMxmzpR84vIO/cP1i
8CTZV2BBYT9k7THI1N0YssVVij6JeAl6YuQfeLU554h0VmYfzIf7+kyuIyHCYTGg
l1lneAkDZfjJZz8hKyYzNygPEJizvakiIiKJ4DnMc7g2sND99UOsB0uA7ozGFRQK
B4ZVgzr2JaWL78mJuJdI4RQspYlzYjKII2mSqnkCuvVcmKpSqRHkTf/o6hU2bmKZ
DSS3zcxAEsBAuLbmPDR2Sz2GjZFFOC5S0a5SSsAG56k4FFSzIgpTY0qZDFGJvBc3
ula2apik8L2qrEDjt6EmZYU7fdfwBF8hOv6SwrssmfI05ODt7eGCvBsopNDcOps6
8pgtCXpRfNzG6ltu6H8QzAeHH/xbdivZmGzqnDFOJkDM8tysIgKU6Ne9DbIli1j1
HZJuzoxSRXPYj5DK4xfDwc92ClUnIoUYx7fuhwYFoveYXUs0E4/J2jVsekRR8juU
dawchppv4mkng5H2IPZ8dD2pL0Neb79drvTI1qprxNw+4cc0VeciHjQJ4x+M+Rmu
1ICDAKObmJkgBKExT5vrfSMTBJptipy/gtDZaqGOB7GHeF/JR34zdVSEwTDYKbg9
xrhfnpFugl8YpsumfCKb4oaqv5zu25Kk2TJjnizR3eY3AtwdFw+o7LGb9ESVMlyu
sItpvp3XfpRGfn2t68N1G2JUCyikBR/2MiVGZg9vIcZb8KJSatc2eAXqySAgwJ4D
IP/PKhhYxU7z25p0GB9Sz54G8lN4h7HUKA4ANrB+hk7OYI/a+fvqyIKH6FcE5IEs
ZUbyngyg/rWhCIG5sVbAArI+18ZGZYKBCL7IrNjRwJewfn8LVunr2L+JBkKx/8EQ
esnTZgEnDLGRK5Lyz7lJGtFSpHrtzNkbTP8sq3xhZ1Xfmxfr8EObtH0XRoqH7An7
ZqS73UBw0MK/kxeRirMdAtO9qa9D4AWK8H9G3NCEOx37mZZX2jOWd6IjRT6nWkM/
FlirapK+QZpTIKlkRluc/uZa2LbnBKrxZWUX+Z3ukhJ8Up1k6HScW2Csv5FQwWZZ
aMepAhSBvvuJxBlR5n7it038P5pVKzvjfxVdSGS8P0JVq7dFttO22IwA1dR3NMcA
2x6PsSzjFNXft0wa/36NMW5zNZkQ8STvOCJy0Wwy2FHPkoLISh557aTRqy5NvU1d
G7yy1J7AQs2J1eQFt6NTC2Yo84JVkczWxTydKvGRjVyLyobw0m19tjNjnfa5D/NG
2E5+T+pLJxbFPAuK0ZgjzSeF6DtldfF4voOp7M1QK0pC6pbBjdds8b9sFinAN3Aw
OncHg7qAQw+EjAkrpGBG7uYbZtmZ87hoXm8sGenSzC7GyMhNL/L650Ps2LYpUakZ
F8ln9uwbEuIzY6+gZBls9eijbwBZpuDw/tRtHOj82hTJH8Yo2geYbAbSetX6BB6d
WxB8opV4GIgRd6cVxQKoEKr91wVl6ZVPsgnuIJGF+N2Ib8x0QiXc5f7ECEaF4UOS
6mSbum/PH1Qq81s0i9Y5iskspYpP3nrJPdm3oeNM2PqRn1D86TW96NYyeMJXl/Jk
m/Cf8Uw4RuwwHdEuw/vh2ljbo5AjoK7rdThBOsUeJJu1om0ZXTtXvr2llNVX1i/p
QT/BUEYZ8rraBwIsMcAoHg9yxK5G1tBaOYtpojQpgDF20u+wRU5gMA/Vq1jG/Kv7
ybdCufmZB+8PFRc8fAytixSXF2qjucHfNGI8WqiMK3V3YtrsxMLa3Xk0Wa4R5mG6
kgiYFYHDLLTD47/uOL/ctZ39FQfXui13/xmY0eFObHQPsFuPOZD7UJktZhbfxNih
hxmak0VhfwhcrzgakdFk4tD+81J3+CCNXSN6kunrMnhaLfOb94KtJ0QeNiR56CmD
i6m6PIFPfFri6X08UczASC8VDeNkAk78as9jTCGEdSxlGy9OB/OgfGcECfsr2Fq0
YmVUmk5IvGSVdbwK73Hkxjf+1UsxlHu7j0572F9o+fq0/Soskrm2CIv93N19BORw
wGt7cp5S8zfMNKjDdPN2fhyms4aofCZQWhvdNckpcyO0A9wHXfKmnwOPxlBewj/e
p8xCnT2oI9wFS3nnpLc+JJ1DaKOaK0JSnvLCJpwTjG5unN1JIhwRjg+UcxGME+Br
yRjAHVpg/LURVwoERz+oS+6AuFn+6fpzBI2rBmql1cY2ggKD19BdkLYLPSbDTw8l
LULZHMNX0vav1EiF4KYZFmcZt+OZ5VkKAj/XrWhIzT1o+k4LWqPx2UqhYchGzbsf
zFCuzUZ23uJCMxyIzhvSBi/Obb4zxEjAZelRCV8FS1DmlTe7WNruH+wtCprapmHa
4vJeeadgq4+Asav+PrkdwOObODG/86UDRnhviDfNPXIe1i40yY98rFQMITrPoAPd
ld6Q9eLU4pB5rdBVvF4b3Yt2XU6L9i6cxfRZOi0eDLorH6WI6qlgOSBFJmgakj9f
VNyfIz2DGambgWFKmQzvEy8ifYT1YzU9+GF8nkLt4BB2C8ImcJgnmFn+o5sK7zve
67u9S34Aw/qYitoRH0PVE/eQ6SsuoKaNWFXolXmLbiBcSmsBnNTCf8ds8nULj3gD
p8xzU9GS2O3+5n9x17z5pjfdjzKNxy0r5ekCIFQpd0hpVNoHL8l8O7Niq85ya4em
TtQOoEjJ84anxTHJ6tMeYVW+Z9u31Uzb1JX9FT3oWR8ey3hieJNTHDYEOKlR43VU
A2F9lNeXFnpj0vOBy5DtXjtsHPr5HTNMcmOo6p/PVmsKPwBeSGj3dt+skyOlIlL6
RB4m4hmmztQFy9oe5bxzlvzMg3ADWYNFLJbOoQOwhYs92LOBu826Q0wLjNR7kt1K
3j160i/WXUm2kEjBhXID3VxCgq9ncb7ZQ2hoqyWOGNS7HQtZMAyUjjLapFlAfWya
cgN1i0ceriOVKV3+TtexT1Fo80USYBYn7PaMmnOzBxMwsRlu6FtAYmMz4ZReSo6z
X2lSsjwFSZgwZvWD5o8trbDUrL8mv2kXUbz38obWIiQJtTJMc2BywuQ25gWJiCaQ
/+cnlABoRfigOmo8gDjbAXAGRDxQ3Vm9mreTisQVB9xi/jyPr3rmmR+LZxqs+Itn
PB42twoAeTFCZ5wHJO3Q2FbNsdFifIkax9IQiL/A4FiVmRo5vp8NFwsKv54WERDQ
GdyQ6TXur4KCqmos2n4Oali7KoGdSxxeQmYdf56tTfqL6V/jt2rVMwqaN8dj7vMA
FtoY36nyXQyPKzxNp5nvimss+d201ejOV6eXybSW9wTardEN8CqwnmLptkDZ5Jn4
in6DU781b39ZMfk3IYahA9ONyM4FQpN6V8YlgfJsKR8+E9vCbUeSqLhNN1x3I5PE
6kLvgdnSHcOegOaLX8OGsyveHBRB5W5S/un3OCmt4rtRzAatMhMc8vh4ExYlkfaJ
pUfczIGjqOUaOqYBTBDo+rkVN8qC7AnzYTBbNzZ2b3Mc4GxuwYYU7rw25iF8VtaH
dTMw1PjZHjTUuhi5WyxH48/r89lEWItAtSrLFP1QjLlV5n+KQnTFqDn2y0ujNsf+
BYt6XcCbgxTfDATwxxrmhIF5Epw/pE3a31NpVOcRCGHYAhJHCJ2E4LW3yClLf2dR
lmWQjAFaqyEXbTrOhaQd9wifNaCrbN1M94LR1d80i+TBtoLniWvOZlqAA131xNjF
AE4z4LKmXlm8JfLT4eZmjhrwen3jtDd+hZq4Iv3b/7K8tv0nSCvCZVZenqsQN5Mh
cGyv0wRYyPjuK8ngxePllQ/G31CQBYOuc3TT1UZoljMaFDV1mvfnQ35Iw997nM71
3HqoL5D9wQ3NCHWWGRVH3ykoN4+wc1njWqcxEjRLrBe3hSqcMoQDhFkXnS1tlZUm
SZeHGNyHZ45RI1oxtOOHMR0UOM8/gbxyW3FIB+nF0LtdKBcInAkQ5tMNM+SpQChx
Ry9EmvxzI7pJSPvuC7jVZK0KbRiAg6Dlbfprsnib4lEPqGPCABkuKg/AVO4wyBti
OqkMDnR2BDVs765KBXByraYTkUeSZ4QY1VEHzNJ/abPtyHrz/nPjRCuOlOuF9DYm
1jHGD44pnlHuMJYHbCubTBMkku/vlI6lm04JmuxHyOnphU68g4/WngzPtAB/CU79
ALui1nzBCNzfaBqpcGI8qLmFIT8G7OPlyYw4W2y/osx9yr0iOa5TG9Zjx23FnC+m
xa8XrUhc6+J4XWH8NGz3YiEszLcpYtTJhqQVyX2KM4F71ZouHedtgWfUNdqzlszn
BRNLMgg878bvLoifEkEygdj1bh12BQRvsPgqedWlDzPo5FMbe3woKM/ibUX2tBLE
sSKpLjTSiOhWJUZENvdVynCQOtcFVHiUD94o4qV5Ybbs/OCcHIeRjsiFbkzfj2ea
Cvg6QIZiHpFTexZ+Yax0zcQIJk1IJ4lGSxuaKNHT+KbhVw7nOCS83r4x3cxWz6LX
xCmCg5y9ePcxeFTvZdCwBYeo6KGC7hYHl8zJkdyNeS88wFuPy8qwNNZ6S2CvGU/e
69TLTk7vXf+qU1YVIPkb0KGQjGa+t91WM0lFGMn80zR/7eybFeqUW7HRFqhsQ6RC
oUe/BTuXZXZfyitzcrawHVjxpOiVX8Q4fowqkK44XtDyvwkW5fJiB6Pd+pQq3jjm
5LdVkA1bB51SMO/648YlJ9VzulsFqaYoUrGg9Nsg9hLeVk7cAYb8lQL96QczVGkc
j6wwow+E6/I50i7OEloyacKiJJAAhK85+HC7Kjd/NZAKGRgx79fBH7M+qj1FFnnc
n4zRETFHZPJ0lqPsoKCtwGKhmbfwFCUUc7so3fkXqNGQRTXlY9XdQO4qM9kO5key
WGHKUYIF27MY+frEjWuNHgnZka6b29ahtbWD/37X8EiCIkqDZBCWPbLWdz85iBGD
QdV8LrUGzE4QYt7YZPzv7wOUZ7evgtgscQhXYE/Bb1IBsnNsZNfl3aTngpgT1Zeo
GJj8KOO4C797LFuuTy7knh7GUlBKfToIDo3Xohogkqn2j0fODE/1qPpXSV8BuSjp
Cy4VzjFzKFlj7F+e+MxLhd+CowWfcZVVhVx6A2fDgu78R+pFoKRPBgbJ+HdaLTfk
5uXV3pAw116T5XJCfuFwScDyQSrl4+xpbgnRLDOmVSSwYiD97yooAF7/td6G33jx
iGMCCHop06D5oV/M9NY82/c53HiumFN7+qlqa9tivVh3xl0SQwvUxPpZkjFZdBr6
ZSDOHq0cmoBqGxOH2k4Vyl2shrgXgLknGWvHObsi/ObbBRudCJ9Cs6t/DMDPXkI4
GZywgz9q0KgttgqTC8zLXl+k1YDXiQMzw33Thxfg0h7/PhXFVUT+QijbdJy7Lzg7
aqS9JagS59IwHG9nOUfxYOCk9lOi0R8h6kgx/FjTo2FpOMR4w8tyLrh2eFwmcB2B
wk8j9cPIHn65t+EwntVx3DdAgIm+vrK6RfNZ5KhNuav5wWXPWCcwdt4X2Ug2Ndzn
vcNeG5P9MqRWCxF2tPUQlJKCdlX2Z0WYZnsExkMVcH9Q2hcCUbXRiH2du5jVbrrS
oP8xgPlhILW/KrNYE8ZFMbg+wztljLvchYsGf0cutSE+av1+zj7MJqFPZLdjzgfh
F6YtxkFBePrGNqvaGMmtt0Pqp7XF3D9KgwVCT4VBkehWHMqVNq2W8wV6C8ECr/6r
UX5ZtTPlQ2raCFNFJVuAayMX/qc59/uOAo7bPZXK2FFegdAsfW+scHWAo2wOvJ5J
3xgmxrd0lwaGUf7Vj94upovBa7QcK25zl1jyfr7AaJnvdl4zrMoiNBel435PVrZT
t2dMCm0L5RZBwOyMeEtAoM0x5x6TkgcD46E8VshnFp1OFwK7JXQp6LPfCjmSvZDz
4X62r1asC29MhcDMhBQ88kex1Ec+6/SBgslgnIn1eurGChs7+fgERJMhgtpaVQR/
UXDBO1u2NleUpIzguiCk1AcRt7D6h11NNb6tT5LDIfj5rS4moYCEjcnd6CeSQKw0
XW6SOF4YdLInylkoe+WMCHasoKec6MZ6MlC+u72zIi08ABInoHT6m2XP0jXH/4eP
z4txwanG4S0cdhEE+qb6GGrGLwVdhnWSi5v6GtIGOEl4lo+ZT3JYg/JuYZ5NvuNb
QgqGNCgYKaFl8+k4FzJGg3ZloWfadK+iPm+eoU6bDGJrW3/J+B9fB28vA6Fwr3Y9
qpUyh4vxXjbFNPakz/vxWPvhwHSqCWcosWjXAvyzXp9KxYX4Yp7/Ysot8WQBKDnz
MW20Fi1OIrB8FQh3dwNQTUO8GODFFoGkFgEDTGcnLEJJ69ercOIqF2LmxmlXuMvE
ldVtNa90oJds/m4Tya5q0hHlrpaEp6MujOt/A3QuO+EQdPapIlgnQRbY9uM/eHj0
Hh1j9vQ67+ZEhhUo3mTEnlDXktEl2QPAJU0eTLH1pEUQq29c7JX0/5XSRNFnVQL5
K2zSidVcdCr+U9Cw5x9FwuDdrDp9ivGcyvo6SxwcshKicADjmXRY8kReqk9Pm2Wp
R1Y18rWeka8PMHWcau0cn+c6Il6qIO67vYA8kW4K9+HQExq5t2y8dUq//4zhaMFy
w/7QKR2+NAg887YrRIO7zndPQ0L7Vt1Fqe1YPgDuJRtt34lYTgYL8b//v90+0DLc
e3yKqO0qk6HyMXxnvNFZdPMuoWhcZsQrZ3W2DVVj6eC2V8AT5Fn37P7tBPE9PTHe
vU41t7sPndgjoziiOLbsI5U3NdYSXIhMFahAaYfubwdVEUecpI3ydVDQYYDC1Wsf
UjSgReJS3SkUN9xmgsZdPZ9KNzPLomrOYxNIeSn27rfX8WUw4dKW9TnIqiS8GLcM
7riTtZnjQaiMzpzEVaE24/2cLTDJVjrTJAmydTdLG8MVixr/u0Z03Ry2z+YHOvJS
7nWu0UoPlzch6Nszs50I4xRitsnC5UybVqBgvosK/sqqKCJxoTAt2wK4569uwmhb
LPRozr7o8fKMplNmXUcd+zzimXxdKKd1SkmBwsvOCgHBOb7pDW009QFcPfSgP3nU
IHILvSnakMw3WKFAMJgUFFe4whkYef6ULCds9a+Z6MHHb1Y77mAKtNPyvQiCZwXD
q0uwna3WDBwAPXvPPy/S2o5h/JqnvstBCcNgCbXb8gWhyDP6I43MZiXHQVBYM/uL
RdaTgJqmggDnP9Peftijh544NC8AHZGke1dMWFqOB6/X6UVJKmWAqdLMFmwihTl9
I+UI5W/SIAB1R9UPrVo7G4H02+oeEuRidGN0KB6QvR9N5hkVD3x/cCTo9UlYmq/V
7GrS8plgC16MuwphGfq1GcRPckwmpaknhX+VpI8aubhIncUgTSdqcQv7ptUN9c8A
JSO/NSGV+WeVKkJPBZa0hugd5xMeaQqvsfm0eFH8/HHK6LHqfLE6CalfX91SFCak
LKLit+rJWS/nfJ4YF/Jk7yPNYatvfP0FhWdaTQtjn9l9LTFlYwhqqCMcm/gp92zD
ASs+fSFSCq9GkPzw1De8Q7I+tSUGEM+OfM8booAT655O3Xg1zOV+7wPNpCInT9FO
GEBpzZjIqhsp9AeQDqbC8z7hAB4c5yGFDVD3LaBaBmeRF8eVw7vgI51UdMVwyadn
Ye9f9Fx7fFWzxr0yLgzKWWdWlT5LHO/vcz4p/+3iKbCfCNBVuxuCxYoPfaiwwglI
R5CqIvTLL0YeV1q8qtTwWe3EFE4uNKyp18Gn/klycvSCuMuM2+5jywBo44GUgT8p
C+8HFvQRcmCsI/KzjdIo905odj0byus7aLUph50LVk+xkbEqFfUU3MCOJAhslbcU
+6vxsVPfFVpqXdCf9BAbEz3GjJ7J3ez24kv7WnCvkxJaU46HbMpc474S8zOayMmw
uu3llI7qhyApvP3n9zqOxLh50oh0GaFx02sWv40m96bs2hzRbd3P2D8IV6VsOj7+
DDx1ozMKL1ksAwOAAL7H/I8hxiLtFXx2UA1aHorV9iG9VWwzB9VvMkxR4tNmgYku
q+a0E6cvSm7ZmFH2k8f2LFSE+ycHG62H817gRCDwfWrevlKY/5ZBAAxFt+bH/Vla
FKE5OMlfiFtIWYQs/5WcOcXWIn08V9/PF4/Lx50eiIf5YFs/YMXUz01luQAoRJ3L
0VjRj+AXcYAXz/JqnLaVoMacskvko50mIjBF8OH3Aoyqy/8NhNWm1gXgHoX93/Kl
LNeXMib4r+0VXxc3ZvnNygvXxpKnKNgT1gcuhDo7/VFl8RcqVLLShMZuJ+x2LVH6
>>>>>>> main
`protect end_protected