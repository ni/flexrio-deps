`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5040 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
ky4SiZwRIlZeVC0EoaoEA51p+crL/avqNwYfM3U4xdCNGxC6UpjvGRXqyasCAA8J
fzc7I14RgwGEOECfBF0fc2X+TY3HelGJAyG/peXnffcRQTQ5FKCzudW6yrMuRfxi
6/jS7JuPg+kguaTE3EYinpViaZEMEtrAk6oUaLhAVARmOEF0b2kwuBY/w+GNhjaG
CvjrVUk1geLmOEIhes3J9WEpBnQTo5Zky/RkFPco19TZvqdbNs8SHSl7wVcLs1rE
uKsFpdC4MWX/ZYSmIvQ1E/6L3gIwrCYlIMlQ+sUxya2GLZGMenXLsVdLE0/Z3FpE
OoyeUsdhzXx65vRRdgYfsUx0vBx4Na/4/PhTZ8Ev5EClJcLwL8eDNmhHzzjWPlQ0
51CEE5axO7klqbd4RtbwD58tJAoru6Cd3Rqlio1aHrk+jTGgH3olG0R2cRWXsgQm
rqyCQKj4cUEGuZDENtv49JAwr6ykDwDzmG30x73fOkc4g2se+Rat9odPCs27sZ3H
VH4BD4nkMuEol9YcbwE9TgzicA4QUbo0Ni6Jo/fap/ce42m/cuYfTJsU9eqnF06k
TIW7mnJFHfkWOlsFs782TVIcEnXDL+2UoukTpxKwj/lNmgnT8L1p+RgRU5k0oIwR
LVpy97JiJZ68XtiFF/duGtCV1S3GXKdnz+FVUgLgQlLJzM9KEy1yyN6SY6VKIkWE
5sXvbiZATQhsSCQgPC+MBAdrpfuicv3f1BdYnWTnlM2PsFy3REzvG6OssdPAn+tn
xYH/kN0bDFzR73obwLh+pVEgb3a6TvyKndcPm8GpauKNymKCt+yobNOXrHNqCxAZ
Q880lnOFFH7n8KwzgRGemkG+Ky6iI3XlO+4bIAbY8KXoPHBMOe2GggA0XkcUpYXV
J4oPHmBillxLTDGKoDErbXZOaFdh81RbS37CvL638aAGYSbt+h/Fpy73/B74+T42
kCJW0h59COkOE1QRW16rdCB5xksouVD7NHf/aLvCBaVWwmq/BtN0GzUlMCp4RFKs
cwEUYD2K/MB+0uw44xNqc65WtYG5rEvSK/qGaDV5GDLMXxjDgYHrxJuJhu7t4y8U
RQA6MxLSL/XUdvQd1gKax00jXJbubr+GcpIkaREL1Fjx2iXpLnly8+E8op8As1T1
gaHfAv9w/1ErsuYe9GjsRHvcpjgNN6poKQe5uOQ2GhQInjRpFiAtooFXxEVbgpy1
rUxA+lkNzyrP3OZcVv3AJVLZ2NuvYV19OyhA4XhdMopvMO/gIzBkTK5Chy2MEBAa
J0xyOtoZMs4lm8ZUbLX9kpdkPzf6UgK7L9AgIWzMQutyBwOYUo3rOlVByN1kIHyA
zGe99gXnW3GbjTsRy1vu2LeiMMY9Jh5XG0FwENdXeqqtqS8z4IgFuxW9rroCLVbt
QOVtpPHHVIMtKbTumx5qWCTdC8bsVDeHoWxRN4ozZyI+guc5gns8+aDGaQiRo8H+
7ofitEyw2dcqgt843aT4+rEyURlxY5KtlTRjPjYKVhvHsRXv5GcgyYmlMg8BTh7x
aW6LOkcPjjOa/esQ3CC1s1XnFSNuDu0xpzTQWfzzmAmjUEdVbRf/AdRxObR4zFvy
MX1PFyXBtxfKdTma+Ur2Wn57/wtvhT7tmimaFgGpPQBXoRVJyiUTYTRK3F0UltiR
5oRbIOkqfGQzvE21Lj+fZNu+Dy5IX8MhHh/l9pCLwjkdkfn0RwuqxmNC4uhy2w8J
KNCqlkru/r4LLZqxTL9f1e8D/YZmXocjRQ7retPahaD+q9tqNxnm+VBYP4eVdQCT
oWvAueOwSYS08kf2PO/iZj4vzMuT31ENJ3L7ORMJ0r8SUqR8/8k/ODx6d0EHKKSa
RIs95n1cOL4QCVmd9gBceZhPfYeJDMIin6BwYQ+EeDmHc+4Jw7ix00T/Rq6hEBnt
orhupjBtTUDWbMynZ0uXp/fB0DFaLdBet/R4KVBbnRHVuRBR3P5KTVZisrxiIJjE
p4+jpR2KkMMYldgvKEcKDOtCd8Yri2j6ufwTscL6K8onq43wW0KFFw7g0NhXP5B2
9fj9vgfpXuyKCSguEyPitQZ5K5Z8YeJtU6c59mv2AL6yLf0SWUyAIkO86U/uVHGh
4aa7NXCGLZHQyarn1+DiNduuZg/O5k7IPS1jdho//HfPF1wyCUchDr7AigQe9KOu
P7If17rryzZlTahMmDu+/2Mn6MLuULQkXMtCtI+fao7qHdr2pCj5AxCh+wqEDG23
lzjJlCReQYyCHMPLrvBSzudGUC/Y3jU+JGzs0lT90fLZjiaovsOAJw1emU0Cjwzx
JcZU0Tw2sPiQmavlXaf1+VuOrZZ/94SKYWeQL/ofbzeEeyiCCbQRZ0nLmz5n/L2A
8J4lS/Klz8lQBWw4bS7Bet5lkL3CGjlI23lURs3hjUP6ekSEb5LWQnrTw93QTEXp
NdF62fKUshbv1jsJiZ++AS7UHqCtfBSYKi5rpCBp6CIJyB7p1L7IiQnRLec4itGM
YBV8rpyvul3NLZ/oi+LIzjXgwj7GyQVjqBFiAG9+wv7bYmmH/xgpNv0AcOuge9ii
4/X5VZbKHaLqixa+hVJ4DPKW3sIhhGHbMqHO1OuUpYMp890Ohbf+35uCRI/WBOcS
LcovXSwZSTZfPksRVof1EQzHzXJ2k6rh9rVea52MxEOjqHB1y2GZKIk3mAzqQSen
6PEEL/RsqU68e558SzTJzFpn6MIuD4umxjCBwPLbAyoxBXNPzs4MoCc2SuaXPMr6
CrVTWRrh8w3JVvuY+/WAT4VnO4/MdcwQGVvsbvjzHzWRCPj3gSoG5eHepSho7IAw
xwR5mZV+VvOGDxKlpIbzrPkn6nqQMlNvFsWs8ZxBiCixhnYHA+s9V+m15l4OV2fT
rrUqkvig6KBI+/udydtyeC5o93gxaOfAmDe0mje5pFUsqmDLok1r1XfZW8Knlvrp
6r8rT5c+bgsHkwJ5aXSkEwblFhbLKeY/T/LqW6WCu8tSGVMqCy4fuCeG1Pinu04K
e0oCtsS/723+3KSbj0c9tCqQ+wJia0KfE4GFPXPMHYr0AAacq3ZKIGTo5Fk9vmyV
ApStigGGDrKIraHwVTeb5QFpwS8wYCdN9p5gYRQh5+zBbL1gMtWq62/xRiY0WR7R
0Q1oKkv1JLiQimPAgGdDIh5+mDGesVlWadAmdmVKEel29/4Y1gcubHm+LHyvkyul
aG+UK3QnDlIky634Rd8QanSSzg6qcxjDhS6S6uKfrmROJ71awYd0X0HwCPGQ5guG
zi6KBoSox1o0RL/BWeUHdiLzc7mQjWMzNmYRAYDlT+gMwrv0fdzvBXXpdong7Y2m
4K4MgC1F78XVpZ+aH1UObb/HQDNF9suYso0pErMaKeYf0oxE7cse4LMJ+BiSoF1z
kobFpaFjhKZL05xoM1b1rZyBVZM0mVlIgr87q9QedN3tlzN0bJNkg8ZP0To4Aooa
mWNArYCqBR9f0IsA0i+SYhHe3Td0UdySxYWe2bxplla+/NE2Wp1cruIsNJ4P4pZw
7acHNx18xL9mDBdc38M0lTnGfT9CsckrMTRs6+vmFFlpED+Q2hs+OHkj8KKczJwr
WPmAK//Cm39nmap75/xlHI0jSwc4j/ZVkkECYsDdYQ77PK+fgCdDc++Vy86GYHF3
ToE5D3tCnIoJpBnV0kRNoid7dqNzcy0pEG0NY+4hDV0Cgsw5Bx10PPrM81lUbCK3
L0ooqjDchNnttDZ0H1ORCi4sfYBRZCEmiTzQCPT7k3pOa7dB6zZHbAWNCEG9tafG
aVfcipe6uhMExu6vWgyiU4RICK+OWaQ0W3gRwRp8mc/BcKGJpFo/J8sA+Y5dzhlV
9SEgeAThuPJ1JEUdymEj1b3TAUYjM4SAeMf+hTDUwC2+6o7VDd7u1nXQOT8+9dtg
EZPu97CgeI6uHLbef47UeUquz7APk8SURqA4BlvQBQdKsx1Tks7rA6tcqyawcJ9g
GMPqirqHygy9Tn+XwCnthnhWTWfiwaIYByZ4nGkkgNdHfoQmYExO9BrmUf1BdR7N
i3IcV9rYa6Z7Yrb37wKx58x/qfG2ni3GVjx88wbopGaNPZ/ul4cjd3IiPfHweZzX
xTL3jNY1J3Ri0O4IE/z19paqI15T8Ue+Y4MqssgHSdOPDEo2tCENz92mJcCz//5q
bmkavbXi0G3T6VEnVgI1UaA323XJgAbHbeztwh9j1O+VL8HzCRuGMDMfuZlu5Sy7
Y+e+/e3gwvwQr1Jq+b6cCO5ctO1r2LizHwGiZ37t+dy64TdWQ59GlbuPhrh0/z2O
pGkRr3L+j0K/jve5Sc5QGBDPiobOAlXnSJQbZ8pFriJB65DnHV9Y+rgNX+PCnHx1
dkFJVUlMSi/XkE+9ZWu7lM2/az/FICodskWAqkaWo+27R+tLNCiI3H/RrL7f3By4
6XNZih1Be0REKQc0jqGKGl3ez01EGMvMua2kfNb+yjPNC7E6Dd6OH6ick97N5fxu
0KaDtxjy3aWbxJ7jRgazrshTP7tJ0nid//Fi44o4CUKXrAewzI3uN4XV1UuPiFz3
Gb/Q+k8zwoK2R5K+FTroVVJ6+WSWLvDrTmwoC08raKa1+cw+txofVSQWblWnmdvN
fJC3EPTFRJ757UoR3tR8KJwydP7nO3dP3nkpdkv5wtwknpbiRKxHL+CZpCkX+xSz
LeXbe5AlBeO/Q0AASLSF5y0LYfmybSLjwcraRqu6W7SUf/b//QpJxge0CVZMnVJm
7MURgaXqcY3E13tB60rieZQYQ1rFulN5bYZ6Fo8YX5hNrcVLdaTNmvCPhQWgw744
6XrkQQUOJuH11cX+W09Xe48RFdLjbJAz/vwrq+AAXKetX7FrZ+8DGGUELq3iCO2q
9W4YFj3x3QaFfy1LLm/SNH+MaLJJABV2SdMcn+T1FXbA/HYDLUmktCOGgf8/NrBy
j0rMtPtzsaoScjwVnGy/B3C62BrMmYNJbC17tllBYNbk1HA7sFLv5XC5FHPJ+6E2
mV5XwRaG+wx1rVXRrUsaem09W98HxWQGSDDSon0uO2OXyi9nYZc4ClJbFXDcS0nL
1Pl+OkdBD4QfoyQ+MgokXbHKBakwIOggDstH1yIM2ETWMHhlf0rFKcmKOhhZLhxZ
uDRfJIORbE7duBW/h+PjFvL7oCvooTFq4V+OjD37DiVgN7mZuSp+4I39V3CY7Y2S
Yb/Uzwr86Vl2B6jI4Jo0RcLRlRYZRBnMtJQqDat9RiucSl3bmk5LimRMk/1n3hCT
+y/l8+CIHV8LBQ8BqnHmqYQ8PIMIxSaza+SyVcVORHsT7B7jna/2yATUpLllE4Bv
mlYNcFLEShNGRvEQd1/Yv/FPG6rWaBYDOhfpMsUprE9dPyTT3pe1DFIMsfQjHtdz
rokefVrSIBWeCnilHyfd7QZtIDyMuygKtGKyViRzLDKby63O6yDHynsEIh3Fe13L
yVF7GwAUf7TnD47epT1ztbYb708ZJI5nAiKQwbikrDT2G7j9YCLpyE9cbq37xKWF
s2tGbj6fRusF6ImVSL3zF0utsnCv+aCrRLjzfeGt04ioHJS29jjA2guRXRtDvH6x
yR0zGBF8h5R9GrZRu21hCyoswjCl+I+Sw7k6aeEMzfHv5QNfqoikk0pJ7oSnF4b4
SQm08EsuVZ8cCM/9kFrrG2INnxgz21mZaHRQaT+Er2pMhY8DobHkYNIUHTRjx5zs
OQU83jJ/NrbLN5AYVFsO0y/7zpHCPKWd+P9qUkfCb4ima9nsifvQ9PkO7efUXFow
QtOPuRkwQZr1YzWW6HBnvubhoh5ttd0HA8hXrm9j/NPNSht+H06Iae7NyNIdQSAx
CaFTTRrheRSxqUmMjyXnMgmyWGridkm+mfnZrOmGFwMhH+UGOXE+edm4IS3ct9Xi
ZBT/Y3JTYyQgUOU0g3AOnzsLmD0OPszZatQs/VCly88AOqpsfaDcyl5uW9M9KH0H
hJcIEs90iYZpeKYMC8QEEkW1cVKZim+l8tv3oZxn5Oay6fWKeUgtlHm2UOEqjIm5
vlkW1FsZXSdL0Ro6Xprp99AS9+vbRMPL68AE+ie8qzWZSKcynp1KLxiOTLlDFkvX
lCXJF04Mn8R9sS6GviCSvsVHpIvb2xIuPWtvrRl6dkn4L0Hjl2QXy3NCuOQCoTfj
nbmN99EqBfqh6OnSdMQ0DODNbKe5Cr7WuFjoLGRe8bpCTz2NTE3Ixn2IJqPuOG6I
GIkpv2Xie8lri52n+tmXhTBsGtdLEyxzBJ8+fhyQiOcuVunJ/YSITEu3gaXhIMpE
7QZcwek98bD8inysOoTW/k1IPdDCUXrybbRP/U4ycOlHoWpo8z1/6lVNDGGs9aO0
SlPRKBOp0jqCb0bvLgUUVwzoibJv2C/OoHRlU0WbAOhNSu3GDPgksRrL3MQSYO6+
NAYZz4SpmoI+/KdgU2bZ4zay3Y8iFuXBw1eAAZEDCtyWuk0Tj//s35WamA+OkH+L
aSVy9yiJnGt+Xgb1z2+g4KLNH6g3k6Ox7vU6l7dvpNml+c0ejmFXIAh2/8DUPZI6
qS3wnRHJsDi6kI1C6Za5X9PRN6bHVBR60s8GbQ0aBTOLgpCUgYhIcmV27DP0jBgW
`protect end_protected