`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2992 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
JqcB4Dlx24+2+JyzNOorx2j8IsHamZt1VvflUO2HjTZ9m6EuUhmqoM9+ZjhjiS2Z
d+kfrjQclzgYNfDoBtSluSFoT4Cxzv0/n4O5TH4DTQOBPJ8lrAILaKsDmyG3usN2
MZQtDfdxDp72vP6eeMPeEjEEuoZTpMepA+lXHyajUt/hEqrVcIJbb6EUrjfvGRVe
Z4/7VEziblfS6FB6rPoZ1fWBVWsLqZzFFsJCINmFm6yH4psgvnOaI9nEc5E7OJUS
6ekTgjYebc3XRSAmtxgs/6WpSMYETHcPn6B0gkWXTmwtyTKyveHHmKOKyNQ/HFcR
lMskgJes30jpPDDELE/gitMkPqEVtxK4eljyx+XG+JMLmTofr4zOyrsdkerW6YBu
cJwNVb0klJuqA++nScMM8emY6X+7nJ3q46XuAYWn9Go1ezHGb/re5+eKjRDLgwwK
Iwlp0hpXP/cUr4U5QVle8y1wOcNC9caMTljws1NCesxPXDy/qsC1EKusEAL0u8nq
JuNfZccrbWIZCnpdbT4br5JaUtQ46Zj5tKUQDPaX+Cw1Nvq4Hoo4CSUJn5beJY0O
v/NL0yHSFJ1frp+fzglVpnv+A8kbgSX3eINeMd68/RIu51j2srgZNM08R80IV1kM
+5qK+Ufnw+F8v4xAR7LBSe9Hi8WCpPtZxnIO54iSQo/4RNFpofX29DL/9aytPh+A
szhrDwc7SFRdXk3ueP+OyKSw0NzANNv9HdjXC/NESUJZDnXvRXRB8MPab7qNmLM5
l24BC6d99xhIO2gIS7dPfskManXUhIsDLwUPioeTh6kmWGhlab59hEgWRnOX1ypG
F4GqaQJ8X2LicblBtgeBg1xwLEtE/f7AV8EcAcx4qJIl2EJ6PuL8f64Ahpa7pjVk
5wmYEAUYD6vOuc5OQM/F1NPBSrCk5RTAV9rxnmuM/39WL0l30FfxZ3HsS2sUGEDc
+EKWp1Tommay9QcIv4tk90pofv2g65jJgUyDYuckG0nluyIFtzdsIKJiP/BKFcUm
GtikBXjHJ3la2fGDkVJg/6T3Z4vgPOoAZhdiY9XsgJSorb/JjZ8nDfHAIIm2PpjW
4BPDyxDBqJYuv9WjKkjE/5CdSuyeN2pE0I+w7HJCIkhSOX6316ZFTOq2Td2KBdv8
73N96z26A2PvP3ja4ZuiSG0VDQAZmUSHn4yEuJ3QnLVQwye1i9vkb+95QeYyGsBg
Eeu78CsC6y90vOrVlCuCV0YzFC7jxPMM/ZYCwtAgTpkSTsVbj+p30A24KvEbEtTx
2hNFKxD5XX71yZD6B2zZLDohIjdnZURx45XDo9Jvrx7hOScXnAOxLjyCEx7yizyR
H6ClTlcpekcV9txVb3GrDM7VvQRNrH1qOT5tHvI3NDtYYzRmalDrJTlVS0AtgGQM
qfLunTp6eh9vNLUUuM4HRDozq0HiecSFlVwAFcEZLDB/r3QWDaGkQCqW02fHlniI
Nx74GV2O9sv50NzpB/ZYgQKNn6APQ/ea1ATB5k3dF+gWQxBDUSzqy8PAnyJQwgrk
vuZFB3u4gN6N7TrWpRjW6enVFZGJjZuoFgeR7p0GdfKenJdlCayc1w6Da5q/Ie3h
8M4seHrkWEE/3Y4wNHLylyoW0wQ1wxun0oX7Qo/ZMtzxZPBs0HfLMbPxUQQYbnUZ
qus64IqQWkGkEihgsQjCiZ7pz8G4lwYLwrcJ2axxwKWI+gphmTGs+y1xkVVl1oJw
xVGdH2UnFA5ja1qOZyGVBcqDkSnpluf3hUMuG0MCh6tVH2v3jIJtAd9HA2j86IIF
uY9+bQF8P9f3Kh+CQ9RqccsbzBiJG3/CxXEGcTcQ+w4P4hY7RmgI8DQWP1SmKMMm
myhSrFawmzQpQjjXqt2R2zv5977A9bXmMVHKrG8Pky5jq+x/UhpDMhsHTjsv+w7v
NirZno6Ra+bEXndAzB0zkNgLTWTJMulX6PWEpWSrnTGvTDOQtCQ/gISegHCz853V
TmNop9S686zr2IAPPRaFSTqpofkh+UdSEv+EQ4Wo1XdZdHUPO+Y3evkA9EWUSeml
fH0vwqvWyP7V0oMbrIdfJ8Hvo3MhQKLOTGww3fwER1Vz6sQeSoJIEhGxiaw6gI4R
7jXiSbnFUOwyWTs0YBLBVpjAGJyPIgTBe/Pz5T/shNlyUw4vGgscUHoeOKCaHXKQ
a5ufGJ8dTedBrYhsrw+M6+2M9QuqLkxEPudWNKAWzrgp/afSskuDv0g7q6TWisdk
kS/C4Icox1VhWkfin8xH02xBvrRr7RDC8WlTB0CU1Z2oLRrM882rxAbjZ90KcbOe
ncStkzjeeH6KpwfJTe8/VAika9uAzP80K7o5mYV55W+K7NFSwNm5GvlcUOZ5DAgx
fTO6RM6if5JAxUyWOtr1dj5sAc6vPALbF6QXcHoJlZO4XlU/3fbg7czE8wNCZjdm
mTXKjhZsAaxRR1BfhNcNeUAghLyiXoBbgc9powEXoGgJLza8ZINL4cH71RNSHt6l
c3KKHCKXi0pTzAqvEZPaE3BuIdhDAvNnMbt7v14o8sntQnWQuizAlyfeGOJEnZbQ
yySWz+iDWAXatZ8c2DJQVM3W3jF0D6S734VTPJu16uzhXbXhoCDs0Hhon3olV2XS
9Xprq2qdxPQO53jrPscLME+RWn2Soj2R2p8RMHZe3VwGQ0QAx4K7V8/b1d8zKghu
+QyXpfH78nrHiriHmYCn+JGOe/y2DpTJmb4nieAZgdF0RudyEpIKZxop6APzMimL
k4ZdNVkAEmGhzJIhRyfaC3xalzTpMv24R8sLRvwYNYlzpY5FeywXVd/QvdO1gnA5
Bc0+CbgGbLFqG3zji0Jhal/sKNwEESPHg3ck7vNzqxFMpFHNe2fev/8KA90zpIzI
LdEqEfTMqrvH2h9R9uUSTd2hbC5Xwn175bgPI2gaQ+HNlW1aw0CL80K+n+VrXNze
LXVoMwSdcmWQ+PQyhcwV4iDD/DehkoeH0NQxwVK5eDlgpfGQynk7rxNy0qo5uTlH
tSBPHrnKcXQDQT7NnrZOnvflNFz0XfgrB5m/fCWammwfCsQGZM4UQC9UnlQOoLgt
ax5IgCSFEoLCjU4XrJizSq7vjf+jo9Xfn6MhB+ZLUAgehaQW8rxS/kzZUrHi7xFT
vsX1wY9BTyipOilIqnNrR+MNDbRFiqkdZSMj+dS74yvWBDoWsk7VtnD8qt4bAzQO
xbJsc2FnASAUon5uHGSlRzOMYI2skWx8bqkPysO/zZKcAyfKH+PWn7VWQewuyQfl
xd/VDsTe4TCCsPVbTUQPj3S1X8jPd+PhTvB2KmeW1E1lLW9HZ6Qe4Ukcel0Kk44E
JNB7qKZmyBwkn6evUPzSnX8r8LiFeOVWuBU3ATPKAMa7ZFYN6Lx3iPgzTaKgY57l
y7FH4ijbUOcJhrtIhjtr1w2hF+cs13M2wkae7fFUdiIE9E3dyWfwJaNCZepn04d5
10g7ap6coanNurRhfdu60LWJV+pw/GVQ3F9056OSp3lhe+fYoS6Po3e5bBCcdBwh
9IRvvONTbxRSztfk4wVc+seK2/Vx68Cqb891QRxeE+hwcEHfqIDkr4310rWgGTPl
vDOaobsxGb60SYubwSezLPjS+FmGUYO+TOSlvTokBL6D++NLfu9SeQRXGob8ao+7
ywcFgrPmpc8c1+Ie64kZGqLusYvrYOdo5arO3wVs1SyITUD0wMa653LVWTmZhjJC
ZC/pPFBd+LC+U9+efRrueofKfo8Xrz/NkHCInCA0olqK9AJp933QVBdLSqpeyycL
nJL/WCPcUnM+KwFp1XUwsM9rXf80lrwopfsYg4DdWWuwx515ffln1Bl5bkl9a5Wr
PJvKpsQxJZOWIx2cCPsyNQ==
`protect end_protected