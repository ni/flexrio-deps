`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 19632 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
TDkIdcJUWDKCGvmrQYRemHc8P+xeEMS6bKuiqBVNXMxvicmw1S9cCnZ5YhjRu6qY
yKdhFzQtCcgKowPSVYSfdY/Glcg5ys+TXIQePMx9iyjhC6Q0en/HGOPwtzYSegww
T6PVRlXL7hQKGu+C579nyvpK8JeQyY94dhAQzcXFIRwbbX76Bfh2wsNSmZveKQxY
LFF+de/vOVd/CjBe+rq5zWW+b9EhvDJfauq8xEANKD6JUGFbAL+KOg+0eGPplOFE
iIScWbDVj9JL061Dz5H4FZiS0uGR1Zn+3z5DNHD3obzIIVR9E8q2BRcS/oXN/z5E
nAbD7XFjXiN4o/9V0QNGaltdmx3PVOZqlF5z5Lwwy37EbTvRP47g4RmRMTiq2Fj+
9jq/kI6RSkRLGUt5zNKjyafDeloz5xFRAfCpfCbr7EGEweS1PcDy66S08uvtlnJW
lLcCXC1XCgVXu8jHcs184y1rNCGSpNKI8VKwyLQcgQ0sXOYmSBNS4dAiCkl/8Jry
Gh3w2uSFRJ/Db4u9ZlBfFwgP19HefL+s+msk3IH35IE8Bg54VWZo1W6UiZY333L2
uGAAnxLHCx8DKyvM8UA/M6BDg/haXIZsOSm63Tf0h78ZorKBoQOKcX2myU1/6ssp
oREkzmmogWMCwVKBRbv3BqedjY+zPyVa3QUAA9sPwSYzouoIEl6aBmx/7EGlQsw3
h1keUl2nxRWeKGF55x9vnB4iJz5smwO0vFqw6d1rWaiLxtjxLLBV1ogolMlT5DNl
nztxYtOjd+5nG58Bokb/qr6KGVWm4axgkQcwUatqu9y8fprUhWiQ5xX8xQyPgRcU
2oj+oerk0fr8Ar89Ogei3dbSom1hsGX3BZ86NKYvGuWJrrv2ykv0y6y0H7Y0v9jX
L3q81bVP69/1iFdY9anCw+HZ8oRcdX7rDGP/mfntjQ0f+DsMPawICE46gaAcwgLH
ubpkmJzIFJn3cRzLchwIkrhA79WAsDJz8St0ioXoIJOpVL8PMpV9+6DNy4ADru7H
pD6fsqNDG0jw9gzzD8wHwvV8SIjtc7Ymu2uJScB6kwBUny44myaoGOmw4paEVkLV
lo8Vbtzear/R7/f/kibWgohTmvclWFzDAabbM76KxhaNF/Jj95jnjfOrI22t4Qhz
Rpdqe8kHmlmL4CdYASllI2QCYpud50nkF1D3170Ocn7cnDmr5TFFIWloI/Fh7DqL
rL4qyH8sCOFMu4vcFmE/DnEFZ+on8XFSkUc9/2TWkGnuv/rsKuKIDx0lzX1FG8bS
a85nnzmUiCa4jt8R1bz3C71UsXOqP9//IHyvBsP1SolnRh5SxBaRkjSvrsWtiur6
X8kQrR+BH7hBnonElSqIUflFmwnATON4gB+SWlQgc91Rgu7kdv3w9aPM3DrOVtJf
BidMw9CZeqLvv297Jlo3MdqfD7wz5pyJIPFOSKqgb4KuS/LLyyfAXretUkOfU2Tp
WHuC3D0pLt/2tsvxDTW8SI2wDtyd4b0n0z3FWfMh+IUb8m6wKMVyb+YhprCqQcKR
kwOCINRI4gXHpB/E8c1yM8Ug36kju1e14bXAYiK2+ahi3kQP3s7GyClBrHEb7itd
2S1KGrGK06gSdOqM1u5n+w4CLYcj0J+Dxq1a9rJxLeqSHjnHgFeEKAbx8v+9ZEDm
nZJLYz+KOPiSWpJb2eUqVQNXcoqWDB51njenHKtcvuqSVhd0mlpeHIbw8WVY8xhY
DAiMpOlPanSV9lrrZqfRhRuuoWhA4QAP3yFcN5Yduqymu3nVZWuFx/m5oed0F47P
Wq+wX5cOIvdzHQcAFv2feoVgA/oLmwbnDrUnS/B+XgQnGvEKFvAuBLSmAwBrnlNx
ivvOrcOMs/K3sb6DYCpb0HrGC4ylckx5GvwZxN4AQJNHBj9FGUakoaTtf7h6PfyP
OzkKKpLD+lZ6Wf7921p5yl9FkBx7tVLeAOBs0j51mWqQDEuMszhyg1i5sHgET6Ax
mczm4e62QMnCgXMwXbpydIs7CgHe757KVwBxbxWm3NLmce+vGfoN7M7K9Tz20ZC7
J+6ULb/OPFVyLi+FX5WDNNwC+XiP01zuLQWEDdVeVHIiBYXOG/PG/adblJLEtTSp
YR2DoZBO7KC0WJCZbq6bo4p9fu2b602FlYwcWW19+7sI4q8ekYmkiCPOkS829wWe
14ntQYK454OWpQn9AAMYp2t4XXgl+kXD00HW7TMD2xyKX1vgYmhY7zpRlMjaiMu7
bQRTVeSKB330nGut4P1dxgc3ZeUlhGpofAB8xdSY2hqzeKZuWzqUh7RNx1Iz6eYt
AC7imbnfdvXWQAJ1fZZILSgJeTH1SDVgOLtuBsqKrP8FYPpCVTrXUuP7iU+erlMd
ZLj6yC/d1Lb0LagKbrUWusDFVXOAe6SNg+WrhX3SYIYc+DeEM6yWKBKmFB0/uX9I
OrnAnpZ+DxjWjw4Bv9jSny9kO/pWWAJm5wK8oAgxpsNl/EuXI2L+v/uRzxGsvALR
++VTmb13y+ALM4PGd9052WHKA4pv2yHFPgUqN/M+L47UUzd4pdGLy4kbQDfKqAzZ
fI1aRtkQqq12dTeT9mJ5roHty6SadxUqARDX3g3jwChjrGm2fZiRu1Yz1zY09vdu
Zw4u7eHizfJqIkSzsXIGEhL2TIkS2SblyRd3E1Pp0kYfOHAaLAnfvZyq3jZtI7Gp
oW0nELZh0+t8JSA3wateCLZruJxHm5DMQjKijoKJGDuKVfy6IIkAuHMvgev/XKAJ
fo8nRl+hUoRVzeAkZiSb9RIDiwiHTETySu+wOpNRMyLY1GfaADWILeEoe2MFNcWS
2vuIvb7ZamZOtejptVbpvM6zNl+tndRXWBFszvL7u/CoqSrHjTn01Z5D8Cwjv/vL
6mCo/i9f+R7vxYEWYti0/ZeJRaGjcSILDHxUBWJdKtI1FQpILiyj2VudqlU9uDh/
C6p8p2GERWyG+7yz8+vSgRsKWFmvmHWZW01F9Xiq8WKqzcmJjBPJffy44iSLRbsY
x31N4uhMWm92epsnsgVg6ousSPWwIEpbzVI2KbdhJ6ZwQex9s3yilZfDeOy9ccY1
ChQ7p4KLy9i9QZEHAbUQ5bYZ7+6HEXiMF6TnnuQwHJftJNedR9nnO8a1aEphnFDg
VBY467Vvjqe3sQrluGAOreOWCOKhqcfPQE7fZ4QHCWrkp7GK4FUt+ydBFFKq4+uL
Xoj29gqwyNcE2hv8l1jzVjLmkr5EecsXqaKs1lsZPuhUmmPLKMLcNekjV3iJepwP
DLGsoIMrvUQ6C5vnniqt+P4QosjY2T+B8RoqlECe5LWrgbJrBGNL+iVm9YzUXuou
81/1xmYDpMCnKKu3IOXdNQn1Fep/9DQL89a0UCsXvli5zk/q66fN7DnNCOjKhTQA
frVJQHmk09BwiouqkCuQwbjK9xtLBFAtvH7RKrTJ/KBaxihN/WvzVVIHgfmgLQ41
4zSX8I3cHezo2iDAP6UqztGzL7cJhrC2E79Kmpl0IvodJtjnVpqVOYrqIGFoOizA
xMQHyHF0n2bvp1sK8ZA2WfUNw6aQ69hCSTSJj5fRqpTzsAEMe+tyvtOqzGLGRhAy
scv5GbLlMVeDgcxLmuvi/jnqAbe8eaoEC0KF7lqdbNAPA72LrDUCy8cavaiQvudi
VJjr1CY++z63kz0DBqypuxrhQc7jpYmO2h4zEhSr7nn884DBQ0v06PegUZNoHHhV
WD0/1k3/lK4Mh/fdGD5XHH+z/JsQRHjV0PCVl3Z+hGN5HFyjXVLyF8/fUDwWN6Q8
H/2th1uOsrXQtKVtAqtRmvmumDcyZ+uhuLVi7gdiQF3IMJ74hOaF5upbQKIlgEoe
uzDDYwdglp0hbGUQyMcv7vNFu/Tg9LtSV3tExiPUrOAWaSMMYW0+w0jvy8krDQl7
el5xzjeHMzSXFGSbTMGY35OD13nMyKS4VuLDGoff5k8WbHT+6tBaWZ5PmR03y2zj
5R14EMLRpGK4ljWGr0CKduQrWS6zneAtUpqW7f7w57LLOrzjW5JTE5J8zECO7uHn
89AMfq0VhZ+FU98OPNuxX2M8zvc1/fEygR166bSojTU2E1BsbRQ959YeImm2QXi+
BOTYwYDLqIjLCa6sAvNGvHz7k3w9sXbrttmczRJfkdKA31D5QCv/W528lWvBdXMq
PnRk9Z2RRlJER7SRF9PNt1z4Pjjc4wPLh43q225RtqY36v9X1M85E2lEf4Wmv1Lx
9sXc+si0Kk3Ifd0nukzBiDUPgJBmURMYqs+yAVUGzZ4RWXZg0K/qHoYQhVo+YLVC
1RcDmrW4Vci/LH5SXGZ1xVQDuUHQ/dWK7UMgrsIsfuAv7GZBXwGlrPVmoVD9znFf
6UWfenQY2cnbO9Z57QjWlZyaA2JKBjERDPRSSWau6NVSk178uCl7N9gE1HqKMpA6
t9mT1i6PCcWvUzRc6u7K5L9r1ETgA5q2pp7hhXavm5orSCGbgPiqKjEU+mLV47FF
ve/fRuTSokrlf+uTUQJI6rxGKc6eKflKTHnfnAeWtNFK0kV7hU3FhFnzgKfZdInG
bYvsxMFP5kG76j4nj3UWhsDFUNjPsHVlBwQoYvf8aTLTngh6iXeBlZXx+Mp6sXx6
NfdthjmJP3fni0XoZRkFbMjHDHGCR6YeLpLe/etcd007WDdNZICsKe0jzphcrOFC
Wl8LFNj8EsUMxip2Z4qdP/JlQd+WhqQYq8vTXH33fdblwejuZyFRC2ywWOyJvdiW
evToY0UkQ4MouS2xoKlpg4OvDiadLqFvHnHo4i0Vm0MdpM9iOld6LJ8ACdbU7gMX
c0MarBeprHeAHK5BfPCL2/S6OVN9Dp9GVLidM+ICw+m3SV+jPnL25+af1n8E7Syy
P5CPiRgMKJlKLQnXRJ2ovZpCH3Q7wIY1AnhcXmI++JLD1XJTKMzbKzJet/S2jEQD
BCYuoqYfOrYM+YRh9LfJulKvOvhKbnUoVT1XH7W5i95NHD2NIqCerF3KGt5H/E51
k0f0889SAk/lHShpJmMAaX03P39Zb5mVNlvRNetipxXCjEznoV+90hjxwZTc494T
DQecI1dsRwQkdJE4SvOMbt2ztZ88Z2g/V9hvC4LA2v2oS0PjWUIQpLoVK8g0+b8Z
Lvfd4LdCiUR9ihNYGkz/g8UZw9qlTUNW3fqU5YiZm3Fe4HOR0dkqgBSbAOYCaB+U
58GoQ7iRRb9LvvSe8iz35LGQp+HYgYN7jfGWOb/bRXmPXStJr8gU2kf5ijIfB3/Q
9IaOntqlqwKr5XFds6pstTEksTB5Q76ywsbCIdAloHBa8E1eCe4qpSPGCunjRtbi
yGnloDMTZQj7jXS6RWG/UbQSBTsbYParEubc6LQffedTB408Qb5Iv5jcxMEVPsUw
GbKUW6T1ftD/8Nkjeia+4/BGq/mF73Dizu+lktqC/nglDF+z0qZa+O4NeRVIOmE1
hqM7RSUK3oHb56gVR9ML8V55cPVvLw6A7WOpbc1bRwT3/h7YKG9uR5Q62e6caUOt
TIwIbvJXdYbrVbgV5JosyaQGWJ0KsUNGtcYwoODWXlCgbQmKiLRlfoiKytS0ON2f
pqR1uupDHmCyAjpJc8Q0HGvd8fmQScZjL5NO7YDyqrqtg0ZcdgvITQsuUwtD83Ap
yuCTLOTNitoDOljuLAiFVSxCLnORLmJMKOWBpkA18ypqbatnjwmnOs5aozsn+P5D
YJW8xPuPN+0SIML2o0yQZkNo/VGL6KSJQ+pNietka1dhOq/a+dNFJAlkFliRpvLo
PM8qIixvIIQCeoS3xZL0pf0U2jrcgyqQayAcUeQhxdXWVQjJb8WaJd4hRaPo4zZ0
xaVV/imZEjpfPDpMaPZdO2Y3t73Z+AfLADo6j1tSonz6t32wft4xW/K89si5NU6P
v1VfG5JkpXApmD4cAZa9nAwCfMrk3/iQhSxuWdaJdG0LnWzOM4ieBGrvs4aAr5vu
17Nvb/6L8uee3+1ENpVmpT1dLik60kDexoyzLBO0Lfgr0VqBuncwffmwk1d2YP1y
Q71b/z/iKZ9oxd8TZjHkNrSfyg49eqe4RN7QXsgiUKqyyfLaoCJ4vcdvdal/6gIB
hJaavtDjNgcjuBPtx9uRF0aXojFTb1Qq/1tjjZfk169kuoXcyU6518YngcwxYS9u
Beo2PXpVrHGm9BtfeJnrzx5aWWpTMQN93O2WQG7QR30hcAb5VBgW39NYimjcKKgB
/19aYBfgEQFCT1T8WhKpm5IV7hh44i9on8JokcZVi2DHNI9utdhVBGemmXicqLFT
Ydj8SahguV2ybas2I2nFntdBfNACCFoLyYTW73glJmU82TQ9Jj5AAIBVDo1XUQIe
sAInoWpFfkd7lIdjwaQ9e6MUJ5D7M/TwGlTHLgeLQj3k+B48RpWZvsnd5tYPUAYs
Y0/ponYGRNNvIUy62S+WEKGzM93Hk3zSvkWJ37UxMhm2+/+SMvETOAyEpwGyLlRa
cus85aFf7BtGlWwveqMBtq/tJhv6ZLjHdr43nBJKfTBPUuvkqLkqeaZjLL9zEWu4
sZV2rif+7xpeRAwkGsmaVyDWuIb/2LFD7BpI8qbjZ4SPkpBFozdxjinrqdQYD4X0
v/pvTaHrtYI/rc7kl+itVDxsCjsg96CoSBBxnj4CB7cokhsTq7VlTq5gVSftlcpP
A13AhBxvlK5f7gqw0SrvWHU+VcJREEfnPwdVqJLpHI2ha6yPyhxau7NSihAeA4Mu
Z8LfOSfk0J1IokI2MtvzW84FeDeK6S0OaAQ0uFUq9LhtnB7nfipdwXxMgv1q0cSO
JiMiPTLyUKYwP3la5rPai8Sd/y3q74UueOSfqS0dhIiOe83/FB+mEiV35MvIu0D7
WWdSC16JR2eDSEesjZnUd5oE6IbPu/aErgYLfL1zJA+Vz9F8/c5N32xlrbjI4TE8
FVLpXP1wdnsMWkkFS3xgSuDCnFyYCUy9v76c7JhsZ0ZZFm3+NJohufD2mgM4jhml
NYRHbmM56N2ul+p0kQUjcIcTE5vNerPN3AKnkdHKki4ut1Ri5lrnpmX+XM/21jt+
Oor6mgJ6cLeBynEl9OJytzy5ubClc4WDz+vKXc0jtMc/XLBPvEyYLRA2Clx7Xni6
TmD3nhVWLT7ULmGNQq7CwV2VskNeNrQ9fWMMfZTVXnxnrs8aa+2IsEM2Bh0sBwc1
RA0au2BEaYhCR/QntJPnZkcfyxPv8qq513pP15Ei4XwR5TK61fRl2M7NEu5W/o+w
ZZK3AFbDoQdxA8obBN+F4hH7gxItOBIrJZSzWprg2BivqFZYxkD2uSDv150JwbuN
RkmJ7F6h740DJElreCdkntlR9z5AMTwJ5M65in+YutR4CrkarHFWxkmhNcMJAXN5
ew2Ayjba9VZaQcmq31pEmMbBCEf0wbLfKEX8bIx822t1gDdFa6dB9mpsMGzFUnoM
u/MBe3kSW3X27NPdPX67K293jFPLlKGWptGBMbze0wuSkgY3HvN2w6AfW5An7ra9
16uDNvyX2oICT7UWCsA5EqSSssFOPGZ8zu+trWyQBtS2uNnzff0c7LccZTNacyv5
dfrYw5M6DTh3xOkaE0BSGyAiBPnnZypDn+qbdHOVE2SE7uu22NXYDqB0k4cA7y0H
Q1trXquzM+wjv8L/1rquMIMKR8h2/Gb9penYz0sLS0W95TzUWqfcUWwpUXc58U4B
DCNjiNdtSVyyA3HqBp0yDUQf3U0PTu31W7cedWHWQmXkC6YI6JjfgC+A3g3TzsLP
mIlqFLqocMH+xb3TMpEzaQQvCh8R4a3hDi+uO+ALdqa2RRrjvk8hE8+HXa6GXBdD
9QnrRvO4Fdafm4HmCgDMZeyuPVA513fHcDNVTKyHHQ1tGAedEHgqC4rlHpkdH2Ci
Q7qmeB2dXMbUROMu6HWqHe9RemorSFASz4Hj2+gxAmDmEtVTgB5F89SHNNw7YEv8
OytQ9v3kG84IosSusZxIvjNjZZBBhDbLfrG57dlLiJZsmxjr53fBzzMsGkE6cMrs
/SQEZak4/huGf7KBEAUczD9kozTWxf87xYLsgnkdWHGaGzRdcvbAa+A7jJ/aMMeU
7X1cS/33LtbjjgB/tzgtuWlrdqRW5dOmuvZxUAqiHSJ8EWisdnPdmQByMXvOEf+A
mce8HKqDfGK9v5E/+GeEOIH+pBrN4CKGw7HdqbPx7Nu5yAH7gyH+lAmqr71kqMq6
1ujFoJp8VwQXPgwrBfeBANZkeMssNEXEdhDyqszSZMEQOTzqLH9qpAE9eSGY/2cK
qiJ7QWDsDW0q+5M9ByTCWWBo1sU1dEFIT8Z0JqRDgvGH+VvwgoDXhXXOimMiygEA
r8VFSeX7LhyByuCMm1qUY/Dxbnrrvn+i2JbAhyDMv8NI1sZp0bmDXgJUb2SujRUA
8FzwiwtlBIrxMAhmK1D0TSlWYoXCCzt5v7KZcpHXhOcp7RuHDaQ/S1ECwOWiMZR+
TXCinhZmHCUsFOFGFSziTCaPlpx+fTi5pT7uDnNpSXZFTOV6/N8DODGIa1cCE7V+
jk3jES2mfAzqZtbq3omgjAl8sw3fFN7TOiczzKz9eWrNWx7++F+1ziOylK1Or8Bb
d/Neg3vMy1xASWOgaK7OydYgJgSG0y/oT6Iz6r+YuGLf41aNy560zYodaP/KyUs9
Mg/r82mAUan3Ye3Pthg2kVoBWnhWf0X8YS0BCZNhjv8bilahF35sllDTI495o88r
oxQZ9fnxkMjF9ygB92yWsVVn+aR6X/wFGGQYdUAvPW0q6GhX8LsoS92aNcqjvuhV
KVP9IT4DrPQgayGk/B+45y+BESrGL6iHRg996nw984jILOklyqoWOa6g4oJLACNI
qEOD0X2hCjSGGZx2sBKSX9lr5Ledt8cF/V/cFx0WgggZ2lIG1eOvXcj9EE8Eitgd
V+ixJ9qanY0AAZLSusG1JOteGGHYMMIH9veK+NA3RNV/UGDhtPhgLjS/CPwSR1Fd
llvnpUgjCJUq3i5vhjFnS/CqdxXRypcLlFtVpOTbHMAMEsmC3j9el0BMX/MQDNGJ
cnE01/+RUZoq9A5cALQTrQ3gK5rvJ5IGHxkse6mFZQxzdYH1Wd/2JnRznbWlsVbv
c+ebQknTVEFRNoiqKxyhSpM6zmpae244ndpCVzCOJBvyIbPqgUm3PvKIDdsQofJX
LaxvRYIDDobHkXshs5hIHbJxEG3FgMAbPmBMkNwZvX2/KfEj7vU0XCrSJ/0i3DTd
ITNZGng/mJ+0PivpF3etJhhB2roHFdsvqXy/Yu50WqDk74FxnQxg4Jb6jPirHJPS
uQBHDP0f7w/lm6F8zpyDyOyF7Y12U/aPF3uSlnbQGumud8VthS+FRuGSIOXTzoov
LV+X4hTnVKfIjr2ssVjfe7+8gxfSDRjnDO4duH1jJEKCeIESfiwzcqA7VuhpVO+W
0zZgMqN1T1L+10QQnk2awzbJdXoAFgTbTUNNXVmwvdHTNPFkofOuDfnF9UYvUKGD
scELYI+TC5uQJDnrNgLrZS85NWViW4MlIXQqXgzojQnwUfh3pNG2w+cNySYya7Qg
B4tswBDo+8DvRCG7i14kLQbDyc9yTLRfifrYUtOySGLWQL9ntCAxoNrqTJTgW39m
PRCQW73XMaEOybuzBvgiRqmxSeW7+FNyS/x4mR6okkzmvRH8OoTOumNnygak1/zc
2lkIziDg+/ydhVE/uIR+HQVEkL5BF5xLg/F6rWPxoPnEN9Q+xRqQHVNdDX9cN9PN
55OyP17pnvVo/HWkFoqISwK5eZevQvZlN/Q9ieEf2hvJ1tI7TV9IVy1pfKF8F6DL
X1SZKUYoF9NuqBRIoXSqe4aE9dynWh3SjmOmQ08O1tvV5Hu6RR5AWTpvbZSSKCpe
0vGb5kpjBVOjQsoWcyQ4FX3NoSjH8//2PZ7ofHa89WmQMTh/8KWHt7gaVnajeNB3
zI4381dSbTRikudBd8nvF6ZBG0nJrAgYXKmE4Z4LBH2IuLQ1Kjy5QMx5A+LR8qw2
8ssyTGqN606c/oG/RZPTnJ1ksPTCllngJz+4WR8RHom3cbeFWG5rjd/04178ViMW
N+2P//6nnpH2ndAbQ9DkCm6iKtLxejiSSEideq/PuM3M5nAmGGjh1WNa3pPUDPAi
FIgSSI5NMifrtsRN6hBweFWAszuq497Cs9DTm/ihDFrUr3Nnz1ViC3hQZW+4f1oI
3d3VPYIU2ui4ii+e15KQ2EINOXV4NY5T1s8K6pANEqNyc3kKI3THCecYfZMCO0UD
53dvlsFJCyoFqrImR3v5vDO9bpTfi4TAx65niRIriy9n9+hThpVZDEL1M2VXq5ZQ
nWOKvx6BAgoO9IUyK5/+ghJnvqMz3DrOn6at5zUioPr+oVEkjku3rwy5fNEbYNXt
c400k4fvFbd5GDN7+/QME9JIt6JpqeSzpFIPa5NWIWwxWZhXvogRkfG8Fxny0ZsP
HgBM1VSvBRiwxxco7lqpP0e8Hz/KPuR1Np7voHz3hsrAo9HBHUKPVuJOL/ea/3Pn
E+cMs72aTjBjfdwLbIEvt5X4TizPI9b8Jbt5Np2LEFC9k9nLTMyVzokrgzOmLE6v
dDIFm5Clbl9kBSUqhHSq2nqNwKOaoT6c+8Xd+ZH8DXJ6IHSTtYXxqctw7RPjmhWy
OGkZlEroRYfRHN4oY7/IJksY//1DBP4Au7dUJlbGYkr+9p5c0J6oLi4S4gWs1Gpi
WqOQ5Dlm1q2G99QCmZE/zKF6UC5gIJWlGGzfUu1O6TvDDZc0RuxaRix+GgWIcaTV
WoeKChPFQ5xBAUk/gcJN6kCP7x9QeEJRqhPSN4t04fAUlrOY6GYj4kpr8Yd2YE4v
u+HYmW4VdVIM5MqaKFaiXaiuwD4InMWyTQlEJQS67lizt8Aq95uJcKwiL+qCfSmt
gBNMtAr8ikp/NrPfPhkXKmVccURqS9HgFV4KT6/ar/+zxix1YvmtGuN+6CKY7Lao
punT8NfAjCppfWRKNasG6PnaLFYiY1DrvlkYkQspmJFKZBMVre/4U1DRn6zA6fBI
VfY56wpS/9/l1lc70Su54mLUtmrS6V8o4rCluWh+1uP/hQEyytSE+1QdwNZwYovm
8ypG3Q/WwnwEXIqeueorghVTZz4P2Xtjbadgh2OX4eOz+oL1qsXyuti5xKBbQLYj
dH72iifJ1WatZ5ozZNsiR8CmbOIc5hG80qN0XPPXXx6cBBGW9RkQK/BGJ9AEtAZc
XKmI+ZJPlQCtz6U8JnMyVRmDindlTJGCU4MbLg7azPg+Z8UGLOfmRs+b/X3Lmq5Z
/2eKR3TDL4BqRyrZkCvVUnINWg2JIrl4eb+uv/EgKHkpuRXT+GFNn3aZ5UkUwG9z
i7dzEN5EUVdwi5hbITbRuYARQkQ8c8kT6A7qX5gxnkfKsWmhJOIadqtFz5h5Ub3w
099ryuvaqmRzIAnt1FoRxstBwB3NkzJA63KDfZU53eatk/rjdRIght8fyAosq/L4
l2vEgviGyx1CEFE1ONpdwfbFnCn0KF4USF6rblbVRZNPfUNIFGV8aI90xkXWSRto
zuV2SQkZ5iDaUL28BhuhRkU3p9DgOVJUWLkwMGPh/eGHT1kawtgc5yb8qgAzNnqf
JdBzTufmve/AfuHd5raq4ThokGcVl6W6OWaosFhUdgi4e8eh8+slduFxtFOxO4Uf
adyU5bJjFiN9JSm4exn1PtmooM8x5V26BuJgMC+EcvdMJXMb5q1S2fU8ZG7lMG/F
HzMGElMKvlI1v5hJ24nQ2jOw+Yu6CEaDE5luFSHsrlMiE1b7/ZwPBXf7QmnDTYQ/
nAOXZ0OxuZaNzp+kMKG5EL8PZhII8tPZFH3l2Lis8wq/F0mvZ5CnZ0GXOdUIF9G6
8JWu8y0tLTb0HguDf7KSTx8sIDvDO+HZvBaDemA66cRObkQR9lDjbgNhtY+sdb1/
VS8aR/XkNA0tkr0tx5K5JbxV1s26nk3Rhlt5hSCnVMKUPTQhe4lNOhnfi1vn6dTw
dHQyJObCCyEzAsKkDOSazXBprQ6tBbzZLeAFvTCgkPAXXrVvk2F7GvvPb3U8MxUi
sbY7KRpkN9PHZXrF4O9Hq0B5TfohguQiYtYkXs7I1IOn5ItS2hJ8720S3x+Voavp
eI332DMh07ul0NNhcKtBwXfLgjpZ1r8FfjZ6ikCHsbXU4zy3UeRFuzwyeGOgqMqb
kslNQIM9b9IiL+xX9/eGhOkCE+FLWEwYTw6rXi1s0airGiIEo+rO12SXgy94ccnz
VXCSqXQxFaJdqtvtTIKQvi0ihB7GmhNGb4BOiyn/nSHgHtwF9FrrPlwfEGi/2EQ+
FGOiq/hmyts4Ht4JZWotiEEbfm3iLgHSNc8W+PvXQzw/Is9kI9uEXnS+RkKYZ8VL
b2Ngtg/XYg7Rflv/MTlkXAE8qO1dVKwYdN7uiurnS1848j8opY1AYQdWsWaoka8L
ZTvr1EKc51Z9pulyap8IhzFN2u9qIekvV8a/XIG64RGPgUkw/n914Uu3Ht1Fd+94
AHi8Hq7XvWPzgxaV6lYK20G/3tbwpwYhIxu7FAjtWfPt6fwifjbk9pGs0Ad2enDg
IL4HdSelqDd4gUdN47ulILzn670sJrVYsLXO+GVO0tseQu4qeseN94sg+7zdPeHm
ZMml//yV9Ykcx7891PyDaMIo/5n1qNdB4a0htsY9ZlvCvyN+XLKEAtadAdrRZXRs
b5ZMa5j8KGhwsaBFSrsxt7t4jRUg6L6tSjmb38Z8YjoppPe2eT+v9PKcT1dh1YGG
3ciOETpd/lKzPr2E69Rj0kSya5Lk0bRV88y2BYftPhi100D3i0rmIjuYdrR70+AZ
DUYxRI2oZ5knVp4uAXa4ulfuFW19kp1ypmw/eZUOlq75NO6UfYcpk41WdVx+mlCW
mbLXge3NRmOb056pI2Vb4Y+gjA3SXQLqQsOKv/+4sKlMV7wP3vh7enAvtXHnKSV1
/wAlzTGEpneGiMYIOwXJyTLsJgtPsV8wKJrKXWGADSiX4cSzcn+UMw4cL3B7v1Eb
R5FFN7jGxnEVoXwNE9OajF8I1o1lSdVi2yQpDa/Sshkghux6zkAQJLXl199hGIMC
V3ZS4M4oYZOR1wVBklU9fWLCtJgg9OSnNc94rd5dqxvoHhnUyUDnyXz+cOjP7p9F
t9bj14P4IaPo5kZY0oyCVHBibWm5n/pvV8DsTmj12r2JHovxp8fyqP8YCBDhW+3P
PEQt3LSEns7x/fSFbuoBpe+cLxJQbD/9tNTel0EbZ8OUNodp65CB3QUkbg+16yGn
RYsD23at/Qu6Gi93Epoez/mVZOCyePL6R9zIoL+HTrzHClxmugbK4JEGV65DGgZN
Bv7X2ylEomdaGXeL2lbulo81q6+YnIgOxR+Zj9hhGzUk7VyMj6JiV6h+KVxYf/2Q
sufb/ofbi40IzoqBn1cloWFANhpPIxJh5rlCwEycIC45qXD5M6wM9iFk2hNxfWUm
czROG40c5shIxYDBJvHoh4+B0OpcYiF1ckc8kPHqVv5gqQf+XGkTJ/KTpEq5gG2I
p8MfgyP9TpxJ3KvNpCAtg0GiAdFfynPDKKTLfw2mN+1QhCYECif0ow6g5jV54tyL
BpQzJvO/8/IuVcSbPiMdojpFDy6SVg3D2Z5vKYPLxu45xB+uF1xbe48jBdEf/uix
CYe+d6+Iazo0Jdfy846+2EuUqnuw00UHWEEcUzcqHs06U0/fmilZrbfWPltMo4pE
fwozVbua20XY6m+uP0yEpRAbjYM1BSI22Tr6tAME6PcytAqSfPP+J8CVc6o5hBda
5i8KySUSw1CJvtsGn8kVyET9bl1pouZUQTDQz9RFdQY3+TpMOSYTQmCg5EBYXfzO
RLidDPdpH/CrlDukToz00a9o6nR164CfixZHji/+YcrOMHwy+qtcrH3/99c8ElD7
C5aUSCpVv4qYHJMoYpcQ+do4s01KtBk7UOr+NWgZz/C9CxEO0v5NM5wbLHlynZhH
l/XleWEGfNW/HG4QtUNTzD55g1Ffq5pEYBwvo/9XljAbnAG0HmfxG6/JqCQPLVrm
rXqgL0QH5W2gaETKszWfhGo5Jd3Xz/suOaZsQHqkKPAeaIBFZ5Qer0RGUl5cMECw
udtYWSYzhj+jt/E99qKl7V/a92fTp39WpwIgtF5ivqAi+0szMk/632dx3tN/MX9K
B76METMlYkh7SQ2dENbvc1w6/9sHIIvTeVMMvuqa3frT+PffDCOCR0oLK/OVJdS9
dU57QqrKF/RLPR4WeiuvtpfNjVWo0jriqKd4VAedBbMj5xzfhEHoYtHyNEFjpcd2
EB3dJfrMev1xzb4WPm+pRv3avAi0h1HjJkT7gMMyjrkzZXLGnlQWqwYBY3X/bees
i81NACriTIv6Yfdt0r1nphw0EuOPQ27f8UKTRqy7y5e9EmqJsCaMqktPHcaL9+bs
qWv8g+t6gbwGk29JSst5hVutqBr5hGGJ+P12l55XEegiOlJLPTXYQG9OB1iesYNY
IUav2Fe7j4VH8d0SGpF0PHMjt27tL9IbsCfj0RpV0RzO1mbTSZRxrZePjHgQ1ETR
FPAyvGi7NXLcUUuWxTCgbeyxpobBFMjSk3LbwkijbgAwC9DSRUKXokeklfOO01tG
qxS7vG4dk9qE0NzT7NEB5fnJ6rZWOi2ojyhjnSKp+uN4e/N/SHEIwLuseJOQrJg9
QJIkdFVNwyDDrte2oSXZqLld/pr701qH7jL+FoPblPM32ghpJFch2clZISo+qizo
XXUgCf7KZwWK4m5b5vWneP0ESiVWn7Qnu5G1QM1gj/mbc83z8ncDc/3UnHs/hBLA
b0fp0AhoUYMkjm+TiZUk9ilGjxvZ8vmNA+aTuBIGnTt41m8YSs9oFg/LRsTdt4a9
YKxbJJjxleuieirKede+jw0EcrGfX5i51ZUzKqOfDlJrvBC4fVTa4JKCNNhggio7
ivQaRGvydbfbLBVLFgt0MllKnQSJ2esjlCSxNrDHsXHtJUB7JD3nKXoE6gih8Yxe
/71HS916KWSi1v9OgUJnfU+9+AqZB3/em8WG8SmrSzc/CKUIU+LlPodSkHGEAGiv
I/y9Ytkb2XHnsWQB/CMbBHHgrhY2XGdkQx+g+IdIXRsK9eeNqO6ULPJpLU0b2fBN
pIONEo6jVDLFjq2WqH8JOljuX+YnINTRjs6+L1RvQQKLfr234J8TdQ6Ty3Q+otYO
J+04/FqhhZDX4Yr5Xhquc0XCqnhK2PXGuBCV4HuYLJIx4eCbsgbQEAw4LLLbYVNp
fM6zUAn1QVngeJYcKp07+cnLL6GUClcu1w++OijiFKDpQvwnK6veXdxBKgsLtjjN
gNUOo8hpcHgdfEfwz/LPulSzFUU+VVi1XJGK+AIHy9bYqR1KB/fa+Srd0txs/BIc
/scjnbB1/hgwrWwaOZ+nLuTafQYz5IEWndZgjUDOwAJll+sWoYT4/50guAgDoFxt
+toePm6Vqt/cpkrVHFz1vDHcKL6hpZf1E7MY9JOpuegfe4tCD4keuIBc0l5U6hmO
eV2L0uJcprNqCiAn0ljx8sBxcbal/ptzpP7D5U8FE6Y+KfUr/vlz9aVQYO9jZro1
T+XnLTn8anckRDF6ADGYvQMepxi4HKqqq1A2vbjYiwY4M6DEKp5bV8yW3PwMXVyT
S23rBsKMHupr0AuvsYlyiAWkR258lHMjSPMNb58P9ra0GfowZ8VmUC3ZbSC0gF7L
n2Dd/8lYtY8kEF/HQj8boYaJDvh+MpPka1r7MeN8r5jOfs5eBPrpHvWr+ICDr5Fq
05o3ImqrxsQ5fxg2CLW9cq1xUp+TauwFclv19OYEsHBfmkuE25JgsbnTRa7LIts8
Bp9nOEokpR14FSXhtXYbBlAxOeDq4NemZ/1vi3ZkVXvY7hhPw/l0hwu7psWuQsM9
9cvm7HmmU5beRGWd3owB50jfhIKAh6OkbQwalIk02aUf12wFqQv2TcKTHXYaZ33o
2ZoG+7ttxz31nRpv7w7Xwsmn89LtjzIYrctG/kvfGBWKa/ujbda9wPLWcfh3B0qR
vrhqOu0GnD+RqpvzMpVdb9HIRpk4DILxmGiUUyBxcwyvdvxyDSOaEhNat7cHw69e
ROdxzmsKLXD+Sk6zwGawjXWlvrIHC7j5UXJ5iDhc/DqGjjhqUUhV9n93Nfppd2+J
uGjtD23R98v1x80dQFpwdMn91jwcmCtQXEv8tlEQCy880nSdf80ieR9nz1tDY8uX
xqOrOAEVeA8CMeuN/kc+inPR1K7J7PZ+vGiMx4hfnA2cI5/gROPgFbe27rTTaA3k
9zCDe1UR50rI4kILnx4u6McUjpdVpgokcjtI8Q2myJg8Uy1bopSU0QqudKA3V3wa
O3BvGjaWNkpgW0CQ+iM8JgVuEk6Xxn5Ga1EcvOonWbLz4TbzlVaozUxKAJaCYOcT
SFPvWiP60sSZQxCUvxLVUBkN2rDT3qf0bSuIWl/PdSRdE2+2iDwbYeydwl9lLfTa
roEFZ3Xa7wkPi22FX3V+UvIMNAXJqNyAqUkjJVH6a19YydLEhi0FHIQatKZAqRw7
W2isRNluzbDfzsaW6c3uKU4gB1ui7tI7PtB6Q8WZQvqsfhB7b5M05At2uQWtxd4Q
/EI7O6Vn9wUkqrw9Dd+uRYnZ6JI/OcifYQAiyplhNibLVqo+kuT8v2bli8y+OiFN
AslgV4hV791EYnVfuKWLWpz9wczjOimDDOP3hAyXITDU8TZpUmYQCKarCpkSDX0j
faKTAG05PwuHjczO7NlEaiKnTxc0uLBsUqZPzaxg9CXw492loLHFM5UXeYPY9Pu3
7oUnEeVopq2YRfiw6L/slR+dxZRTWOlhqZoeSFrjXbkhm7tydF7KAllHqDp/TlRP
Flq9oqp+KrEfgBQ3um/z/FK/OnsDzRN/CXSesVObzrSjzxbyPjNFfEI6kf+ZMEBx
jaDP325xV8UJQPlwbYzasgFfkK0cb5zSuB83tS3vdSZvqAo9ur/sZ+YT9Fny3LGt
Gsn6SCZLkEe6P4GxdaIU225K4+RtSrp60uDc/pVFMTgZrYW+OBs0FxtxBvazBa6j
5Xl7OBu6uGLLNHSj+FUVH8dMhIa8INa5Ln+Xyk+SSob8YYJ5hvHhj8J21PeXstow
023sqjLxkFLPR8mPYSMaM7yMU5KHK75RzFMRTvL2zwZ0E09Go6Q8N+UYpPHIH2nD
nz+RE3z+u5vMgHmoAPC1v/UFGHfK1YEoKKpV4T39xELSRAhgPrv2zR6tVpqMZix5
fy/R700p23WqmlPkxWSETBCCMDEpYbNkgqN2FiL5WAA8xRqL+krrXd7ljewonWNu
Kw//eHqdrih2g4FAw2KFN/R3X1UmYEqk2EEmGcbEkH2uTJwnFYFGVHvGi2Dfgj3c
CXzoPBfvUdOb1JwgIB2685IstO3K+mV0ies44nQwqPNJiYq1JJ3quNOY9K34zvJT
aGBWHUwfPyrSoCGomaas27wI3enqOP2zXHIxG9Kc3zOxjZXikQdgyyggkKBEXlgD
tY3y7VXYjDZOn29AxclwYFdv4X7P83hph96/AOaJjiQzk000wDi8kyUL+rpwKKEL
YfO8XBMHELXgHSXfbHWR9J0jj+RfdNNilcyba5BNf0ZMK1f2vzP8T4dXXFpdgT3P
jducrzQUALnyBg9niwwioAGWZA3tu0hRms5pcuK0OQ9HWGAbNq0Yz/jYbY4/Ludf
1UkX/2MTBt89nl3Lj6PWtWYz5WwPbBi+Us+BTPzMoy3El7fGfuLia8RxIcw2ONHo
CMzY9LPdbZPIWeGW/LWj4cdhL0DHurxvNgwgr/gahHsb2K4a5tVR6TqtmXViwNi4
VHr8xfCiF1DdAYZuKYBw0octmOIbeAuILIk4FNK7FHeKU9eBvZkfsEEpqRDGY9S0
Ftkb2chI02d1FUR8rqXRsgVKdfkFJFjiYDaph1YwdgYQ6b9LbqMbwdbMqI98k50o
ov1Sc2MJ3WpPP4iTbHxrniqq7mdIOHIgXCr2xosaXY5q+yDG6qEA4+2yA3UeYq/6
RbTLNnEbO2uyHoVqgyJ06VbOU/JPMRpPQzUTfRwriNHCZ0UHkFlK0hGfKuC+fJKa
YKqPdd/mfnwA1v/CnBhVs5A6Op4JdGCpXFzsIFXcD99etHAOi0Gusp2kBfYrJuRk
Gw2TZUnzGXC3NN5Thd1ECThLNiGJMkuj1tDR8KFOEb7xfIu0ugNTC95AM4Q30jU9
ieRGCA5wpd2ecpwvOedToJ7PVsSiPa4HeKYzF3NTVYYUlWxtahA4qVLxCNUIiv+f
qr3WNV/bayvjArT4VrxhYkBO8/xYbH521d0HCHOiYQLaeApbps7FB69lbXmmdjE3
l/GxwO4YGUtMhr/0oabVl7GJ8V4JEEyCPDQvMmZmejDLS0cRzVYRsGWcbF8zE6ir
MfPJ3I9vupfagm5+kjcnw4r9KcFyccXZ0YdM5bxgPIs4q1YQfS6DnK5V0Wfkti/w
3PHdwYb8u02MhKm6wDg5gt07MN2JWkCKyX17pWbOiGAU+EnRDTXc8+e0Uam3DrCL
D4+F7Sr9Lu2oGbGRDH2fuh+R1eXa4pGT6MqC5j1w6gh61FVXIAhGoPgWKcr9wjc6
QBxAL8In2h2t4K2jNhdB42Wqh7WmgQ8j2nT/BVWpu4I1mqVeTzzEejQzuhXZZf+4
A2HXcPIvmSCY8Y+kUdZ+cZJf+vV9Dvea/AQQZLq8mTGoYpXxygm2pTN4MT+Je8BV
zc16tBUisfdsw/Uj8x6UnX7RHb5UeMRAWFXyaD1395dN2qXFwo32U1OmsqNT7sXb
nqVRRxhvuJj3qqOLFZOb+JvuWcx3TcgSzxNeh/BrpfFo059pWtk6K2MV2oKWJkkw
MU5moaZLUG/eBuWX7HrRiW6hCY54H+86VOyOC0DFA6lt3nFdLdemNsYrx7PB55fF
h5v8+RcRWd4RdUHyQj1BOdLtn17ksUSTQItl1hMlS6PoujeEeKoG9N5nEhX/ikJK
IpIXdChB7CmqZXVTKBwqeE8Au2IUtBCyoc57Mw2duUfU0gzEBy5QgBLBfkCCsUFs
SuVl6fH3riE1nKQhr3bKBFzvnLsCvmkqdyKkvj4ckTIUvd5ONmw6vcVvo2tjdHkq
FRXNT94XuEQOlVAlgb2QG8rd9Gtnu9eegDY4rv66F9plcWR6Jghovpgb7c1OsHph
xaZ06A7MAd1yyS9ANvYxg32EEczCxSTwLm/eEm+B4tOvCevahtw48x2LEpcdb4Bj
JIpciy2HKLUQwrOkMi5EHsY51M+XJBefbVuohEZTRDhYwa1ipAYfddFhzXFPjp1K
kckhWttRUNFKe36iaj75hNl+Cy81znEuLOz9Bw1lwJ8jpd48A8S7FRWw+aaGGzhh
v9h9qOEobe6K+o3Ns1cT7xM8Mn0f73sJcDda3c6ofL0pkLdgggdEeIZ6LKv49qi6
WuxM8Q3BSq/ycee1P8dKezqNCzK8ZmB76WEsvGCO/bH8lxD1jIHUFVNofW9vKTl4
iVAC4eB2oPy66G6JjqYmakSmZpvXkTnEW6/wBMXavjRvIi6WHQGHhwsdQatoo/k+
csH+KzgopOc0inmb3CS5KMMzXnlMWJqcQNB0FX4JtrkTvDcvJcqHoKygijjMYwzm
hq/F3iO7cTwEn0reRgYofJVoyV7RmeyaeZ/ur2KiCOLoZ3B8ifwxN69jnuu5aLQ9
2WlW4XNUJcwSpfbBoCNgFnJXxhdQRGtPM9asFxcysyxXOP/XUHZ0hm+ZCzSZDFBK
bzdcaqAzeFN6Qrjcx1Tc/9WZnCyQPHJr4m2CCDgUC+LgL0G4D1DIoRYiU7NJkVS5
WcRfRrfXb45Br1kLo4nbhnmvGi0te5E/yUAfLxfYxrr35AMHCnrY3Pys0i3JKhTr
wZb5k2X807EmRx7Yyor1FCsL83BKNjRLnEyNqsAvt4xxSvFB6Sl5niyy+U75cNcz
cZWbDXTV0LGOpWsGYrd0UhYnu4oNp/+Opls3LoO0BlcQC8dUjOMszBbk9oJXyrLg
eHYFhGQ4KWlvDVg/IvkoI0u3qMq90LdzeduwcooaIdZ3upDGvMgx+GELtK6cKRa2
Bp6iUNrtdbEMlxqih6d24wr7KC68ZQJE1I+MIX4GdhWM00JNTlvo6oGA7w2tJU9r
+qopVUFju7wRVcZ5hYrra38vRXDVEpA3VfX2yGtEhzzVG3KIkkVZhPVDmCi+no+E
7b01HFN1nN4IievJHErnRsli7XxCfqTVrLRVINKNT+d/n458rx7eMkjZCeTL8zFD
RpYLC7sFkJ9EAPyTXmOIyzUTGOyMfvWE3IBvTQTgzg+bKjqRPdZt7GWcN49GqU22
95NliNZ12QwjOliRIYPY7B7sy4E61ErFGzJ+KYe3R+c3d69G9t4Oqc+CmOwIZwJ2
R8dywVTXWB78l66Mrxk49c5lBLEUwmcfKqOZOERVqNW8F2GMw7WgsE0EHOruQrHF
km3JLHvfgv4Em34rhTu7Jp1/Mfv71Ra6Rn41JXWg+rNgXQvShMQcJHcvrEe6CnDj
hcd1GBtWlNXu+pgr1D7WkmE5kOHoznrGgpPGTULUvV1qjz2uKFa0K/Ch7Akb6dCd
PaZyc6LPi7gGS3/jEdtiFgb6KBWlcys54i+CmRO1ia5xnL3bOjAWOWuzDpfOaVWG
lj0b8P/4tsBZl/nzP+UveQqx+lI9qJ/eT5hQUFsdKXHsJb9jPr66dqVk+aXq8F3C
KQ2Hfo+beqsTAgLx0D8Fe+7TXaIBZ7lxO80rF96lvmAokfZissT5+zANozP1dCAe
0HfeylQZZlfuyH5sthyCa4GNJo3knVmRKUhbyewqHHVBYme1uzwsxmEx72GvgVEu
vit2v57wI/c5prDQxTt8ADyCYEgQknPhm7hiHRnz3hU+wLFxltfPfhyynA1zPbBN
MFWjnpr5gJuENSPNJIwPhoXfYuxWXNFtFeUjwVXKoXXxYlouDH5LGoHaIQIaKtgU
3N8/8Y1gbDUpJbtZcX8WHlf9Gfth/T4PeKCir5I9jetEia03/i2+ZCIruFw1pHLK
FhrRomlr98DpUVkoWBxZi9enLOJ7goyec6Yd54tmSlpgH34oMD1G5VxmBOwWo/WR
MA3H6mk96qtfknmm7IRWIyqRnUsP0Z87bShSeQ1ayEqW3GoEYuHEirLbtgDXAW/R
V9ONLmlWjKi4RNykTtdGg/Mv5U0qTzJnSFRJjl8bk2vvqhgIEm8BF9JEGa9giOsM
15SuEKkYU+/X8XnWY8h8551wJ+BbByMFFl5Wp63pOyrjUFaXRi1jbSreEmdtaM38
CQxcDk8KRgl48pQwsuwUXNGyWZH5H2W6HQ2Z7k3ExkYzkMB2XeBlOhXBbQLj2OkI
JKAKp0L9t3H7QIs/bsnJyKj2rEQ9tvV3MtSIvlDNy3SdMy3VKrAZRTQyx/Aq02Bh
GSaPIL3f55ApFapxJrgvRkR7KJa4IXfkKuIP9d/R27CxLtgDEPFxxedD6DuoURUw
Ig4iGuuadNrIMFk/AcRq1Uep0DpIYgnOVyp5iFpR6XOasoSFJdm/9Pp2kFoEo13r
ZlFO93w2ez9EBeJr25gJtLWuYjmcwnnvIL/NywX6q7SAQ+o97C4yMqZHWjq+lHP+
45su/W2vVZjrUFtixiuPaPlIlgSxm6MbcVz/MxYlF1NdeKVEje54YEJ/MV6TkA0H
BSTPBaAkKY96tgnUxzyXzt0TGptnzSDAEW62m/qM65dF8/r6Y2skLMKQ8CggdFV8
RGhTebVozCFZILMXUfIzdB9vSjn5Ab4RvY43KynWb0BTm9fyRKCQoWjMibP9u7+k
ZVQ+f/oZ4STLzMm52QnCd4IzK+xmG6doRuU9BQGiIkNS0Xk/hcRmUzpirAUbpOY6
LgTbUYh3PrYuHjYtuWSzNdEelrSkovGxYlhxzFUMcUBWPvNaaF4L2zARKaQ+K2+b
+I71Tjooiu1SsLXdSSA4gSbMqljDqA0lG3RGei5LsdCT3n596EhICNwHQAtfQhmF
/5hL0jho3KTLTZh2zVva68jVeGJ+H6e5YEIh8Jqi+555hVilroxzodMqfAKRYR1+
0VZRTwc7IV9ff3jqD4LDEnF3DHeaUT88z7gzdfJyv/HGnVsXrTjDOot1JnccaHzP
mDnFLhfVNOR/qX3EU+W11hCn8gmbT3rM+ViNK+l9+BIvisgfrLakOWIJYg8RQJQU
7cR/Y4aP31M06rrJVTn5uOsuyhH6IG5ueRhhBFPVCtyvo8n3Howf+Ji00QtFHukH
kZ3rk7A11jp/I5yc7rp01dr3tdiu2xXP17wKkvYj5zLuxF33iyZLsQICLnKWJhse
rWXrlxZQET/fSXvdKDdH6gtpXk7fdhqoP5aA5iBwfqEXc5V/bX66hcTzzljp8ttK
XL562DbjfU4Uya8zy4I0qxpBEmjig9So/Scs8x7GdIqb9ka+WXBFgJKYp86UAo0+
EZFmO8IcHl9tPgCtCc9zaSzpfl3XVWMNVdHlKbBJkyxmjcQmHtso70uPCuV+9oCw
rf6oe97czAfnLrhr4u0Q/3jLNu6XtWR5A1bk/y2rgk9xQygyoCnbSz/UdBwcUcky
eg1HfRhOKD7JjI3k29yrL5fF47E6kJlHM3FLJVfH2CB5fHUysuMJOU+GwYUnKQZh
inZO4qDc0mLcwj3zvClp16J01hcP2nsRsGLtx9m1qBBOufmxOJYnJJiHAFiZ/VgC
L9162UqxYkfpEBzhe0KimYaEIVkiwihKBXTZWvQLHDPMvlVZi0UVxwWnze5ShCz/
xxFmz8L2OSQ6H+Hf2VNPV42yMaY4mzmRBFZR7gYpKM91w8MrGEoRZ6uXu6HppNZD
1ia1/nW8x3D7abZ6su4kQhAGbHB27SlkMgBZ8NefsTuJb+i/YSfMBe7atW90hr47
CedJdMEopjCm/v0Keu92MPZKL/sZ4m5KOpsHnA0KnEUEhDzrN4OlC3qDYJ3i+QD0
ux4bvXqX+lJswrsOV9vXEVXyX7RwZYGWyoWJiOQM/lk9NQ2cV17BIAlWqGcro5MW
acZ8QOhvBSev2vGJgyGrfvJTRjKFLGuqLHpvPOQWn8YcRCVV6yqt+akDZtdbOHA5
9fOqzaUbwwUiV3QHXXGOd61MX9DpcHwLY+ZwKRmJNhwAQP18vAHdc+uo5C0+pQLF
XbbaPJaVTO+GtUX3D5rjbvoy5Mnr5lKMgR5H751cmYD+znRifbYI7lhx4aj6Eqbt
cfMYY7R7Mfyt+euKJM8NStsutLU08I37K+wle8+mxzcONj9i/mDqv9/NnO1MUEig
Hv1t3hAmW6wlkGg+Vj0lOwFU019u5K+8Bn8Tm7DCBO5oCF9TpTV/GCnHsKzr0FuP
c7R5kq9NT3TjwzrP+xoY4IJHr1/LqLMaIPbH5/Wc6EUVRTmPg1YCCFDz/g3if6vJ
29JfJ9IbTVCfUyzoj5EPjXEwgoFn8u4P1KAjJhj3Px+ZcbRnm5ABFz9JIX5oV8U2
aGGmlWk9a9+CMy/hXAGEijBxJ2Rd3V+J7DxiK906ys5EL2gOD/JgABP29Na45Oh4
x4BOh2BCKmOHmWOJonG//haTHPtdDJ3zgqzalPVZ8mkhxcbsXficlrl3REupfCTt
ke2dV5DVKU6DjdGrARtU6P14XYN8bCAEu9wnCvcyHayYv24HSR4bgN6x+Bo2D0bp
vUyQ13Pis8+uOSFmTHsfW1s+Th3bLVVjuP3y0XuY+v+y0CbyVMAinxY4LmbkGyda
4kBvaNXWiXZXAsM6/HVX4ZqN0repxtvS5hTFeFxrc5Qb/5CWXRYaaFV9S7c0LMSS
KJo0JqSMp+lsKpE9iCshclpd1ayoRoAkCBfC5phgMcNipbtMX+CKLixzCQrE75FD
uEQLcGGyX46eY6OwZLgI9WJmJ7neieRCe+wpbL4WDIJIxsHtI01bTB3gqd7PFffX
ZX4URk64Z8oCkDdGydW8rV3LcxFb5oi44DyPnboR2xLlZ1Lmv6osWXwntVFQLsVh
pEqaR2aArzYomCNbGt1kvPSYB62QOqJ6A1ewK84Wo4YScSPReXsn0V0qyt9pcZLu
LAL5UTAmRwlXSQO6k2qf8C4+YpumYquLBkZqAlf9SDcwRH+q5MET8YTk1I4c609D
dU8Cq8Z5qWEZVLGstDVdm9Fkiee2F5qHryCtVjAjLHXGWpiCL00oFmsDC22635Xd
/DwM5DWvQeEsA7YYuHHIf1ChgHIL7KMVoEzukds64GfbUsLUTvAyYu1SNQQHHUiW
musCPLPIZjtfmZ5ihofVb/GZ0BavxhggiuZSGprPC3ir9+h7/ge969oZJ5fkBVv+
axYUlr+2996/tN2LPDSxkbr9yTBNEn/1i/CyCN4mgxtea3rOZ/lwNXIXk5JJP1I3
WyriOA8frTTfLnf2/8TaJHi5894plNQ5yQtiGuuWyfoam3USZXGzFpVcfri8hmhx
t4tppNizDWM2n8fOOyK+upUtQSxBYNPEyrsoabAiqO34UrqLpnJhFaS5dNyw968B
YsSOzcDDC2tor43q8uwm8RUc0kjyNMohGYy8mXPW/5SLbhxrIQ/TjDRbIatBvAXn
piC7kRsCOHCmAnyroquwiHQK8Mo+LrMzNu9anNSjP0vHi4298ZKuRyl+U0vont6v
AtZsDMjYbS57AxmUt0QkRadLd/aG455+rMSkkcKcOD6sjKAstRjw/OtX/vIKd7Qd
QUUAVHL4fLh/GlayxTXa4BrdhJjn7A50F+ZbnG91kmUMBYykpZSIlPUrNT9MzCHV
oR/IA5D+xpzk09SQNgiNDQRK9Ia5HPYOUnPV92IqeGGXwgsZEDwPnWOfkKIGNlBh
0lXFp7gqZTPNwNSv8ENk5bmLXYX0QU5B9k/c80fJeMTXpGYOkZzud2nj/aaLTzg3
N/5MxAw1/CC8Q/OvFP+oQIt5eqF6y+N2/Hv/oxAEe04NhN7TqibdJF+Nz1ByzS8i
7ZDEUVztAP4rikKHaxbzi31r9FjazHamyY0KnuLJePByQuk59KAcfULSA8H/p33d
Dh/5kpVP1o6uJWkWEkAc8Ldo7ykbwGI+HCts2gbCcZpLKethFDo88UR0z8uvc51m
nRE4Jta66QC94ZOCYCBOZu7tjj8e+TniNh9h9yH9q+5jj/cb1rbnJ0QCAHbA1ROD
cVXYiEH6UvWJ/0G7A6GShPRV/nnKXc5yt//72nnmz1uxoVN4vFt/DVK7Z5AR1e+G
XCDZImGWcL6RBI/eFFsLPWrpQ9ypk+Rm5FoWCd6a9WGRsBpNLmmleCxc+pKM+/YV
cUx3sbMtZqNeUARQYQ832cRZAki2c+YeIxGLy8hImF/kye5+WL37nr1gHF+VWjbr
pFQnUtrIzbD7h+nkdwSU9tsuxLs6qLdR1Int14mxeUbLT6ljF3G/DD6wKg932z2w
xWNRJh2B1rjJTx3AU0L1DS6jiyd6c6dN70IfbWJnPPYpOXqSerKQSzD86ZfrFcLE
ZruJq+PYJs/K/nohFOnaJVSpien1SPx8DEp8J+TtctyEuE8E1nTcf1vKzEMSXrz0
nsgu8HnRO1UikB8wWpvR3T+hWh7/9mD8y0fd9QiZqe5i3VbmnvE6WMnlrBU3xKlA
oqskytmme0WSJzl4QPV9zbNieNO2AT4fV/qxAHDY+3tKkbpyAKMWYyoPf5d6yVlb
TLNxsDumWKPr9GqWr+3gSK3P40JHg6F5SCuK6N2dW/dO9PhBcdaU7gc2cZ6mJ+AN
Pue+gcuNkhjx2BIXwaZCfB5OgvAdqpM6lfvA+IQfjJos5jmQ5O7SR87KOUG9Ygyf
LeTAIDCXoWagkTOAFsx8+9I4MGlLcsEadP8TUbH+haRqxjzFQlLtdycCw4BvvUDm
IVE0IW7WfFB9NNjvZJceVmS1bOVaSywElPi4WkhTVGlBRI+5X+2UYr6GnszK8r0x
dpO4gHSstfePnObUIg884lxJ+7sajkO9WB+yQvS3A0bmmJHa84nEoniNmF3KlVsJ
hbb7MSeTlwmpj7ojfscGPXkaCfvH1yYrtHTgjwIthh6XIN1n8OXwGgQMtdWqEoHf
jzClm2GIKFi2tuBjFggGGv1mf7QfDuyxfSj9mYRti7n+OzM6DOQrHFOQG3BvL3i7
`protect end_protected