`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 21376 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmWdo24EC1SLhDeUV9o12ewQ
ulXp2xSZ5P2RSggIKJUy/anaBVTumwtXp6e/AWaEdudXt5A7c2f04Ylxf2N7bEgH
xdGb7j/934g2W77Dba55+jZH28BQPcwS4jE1P2O+NngHfLo3WV0tu3N7IujONNqx
oLfbiWvYS5QhS+dMKSKqrmZxhD2KhGeNQfX7GvqHoLGUBxXmbFGukCf8zyAEt86K
VRQktvywiLQ6HrGOkZRtBSqMzjZLaq0QPWuizLhe34S3CSqMpMIgptVxQ+rnLPOQ
3za7K0I6i7a1+4/nhB1NkXZONSCsyOONr4WqLwknPEgMpT2nowZhbR/xq+QofW7x
EnOTL0IuYG9wtroozT00CyM2DjoEc+T1Ju27fT8WumLtfBhxRoxPHKlrl8k4+2fY
0COucMEsUrRwwGQEf3NzLv48FudnNLsoAU5PA22ZojgshMqgAEECaeRgZgwqnGyh
Ne9Fi5qSZ4jwEbEj4qd/ooftUbfWW8rrNZ3lWne8asML8Knwunxr7lApxN/JDmfg
0BzmbkAoPlb/xWBm8Iz6IzyPmp89N3t3sPGzjwpzTzD5GH/9OeU6uWsUytO5Igoy
KJvFBjk1SuWQmH9lqqv9fYQcO+/WJaJkZguWmUXET7j9cdFTWqVLNDXlB1ArVJ0j
FuLTzsJd/dXKlZs7R/ry6Ryy5jLj39/mkMH5tydWA5y3PmuE/GmLBUMjW+WgD1dN
K1TQ5XlVTLag1Gcz79K14MxgPqYeLC6se/4CGHbNB0ludR95iqkqiSMwu+h41y9a
n6BYJHt5cPbuXEwXy0Vfw8IQgdA8NtYeuSWcCiIbGt2GJVffA6hSEDKTNczdwKnB
LjlvHAplYPsNfV+DWo4Z71gnMZ6NwGn1SEUiHe3asDaA3W7AbWn2J4dTLHb9NW1Y
c8ur5EUoxBvGueCcdzdPMxqPHGasReO1SEYqwHo3PifziK39Q5NU7YN7ihCTo9WN
ywIWbLR3AkyUq0MU1F1ZDdK6qW1ktdK992HLRjeggzbHzbznLE+9/w5k4i4TDDzV
560yit07nh9Z+ddXx45xyncMVjqZvMUhIa++wAZpTjXjJLX8bYHzzRRfzM2d/72B
RqGEeP/O7YV4IUB60bbcDsEU/cmnbdhxVgK+5jDhVFl6Dn9M5Y4ZqAUGWmNVNF9S
dBHN3fa743ozhUrJpvQyAaH4YkJN9q5jJnN0hcZqzV38YT5ACqpu/UnGyVdCfWA8
olEYk7OuJV0siy6Nuy9ecAKV5YaQHU8PCEDKOz0lcvrw5gqpEozG+RfBYUUAKnFo
BVuTNBOduT+xeNzLZf6I44rjh1srlOE/xYnWX4jscpfXLdYXAlvBT4427ILZxgBU
Am2DBGFNmLx27jOCSwaby5RoUDKJBsd73awBNh+xWxbSSQ3MVC8U0pKEAHYWccxM
+89miKeC+RLDvxcl4i6sUzylJ0O0Cpa5qtjDmFkyfv+wnYCZGPjc5MpclukD3++W
nk7+ItW4j+POvrVhP3RdZehqwerD0/jqMKKJqc+IZLwsUQ2+xWALZlg6iv9cz2Zy
s4YTW/QD7AZQCpCZWbp2SsV65nvw7naREcXD2SMlv+A1h9/ht0B3dtc+p4aiB2WV
OvcKkJ3W2pGOUGhI7Ymht/n7LJ0QIJIr95d1SM/8GkbCdOg+uzbNkeiBOQRfRzvh
0UM5FzNnPkS1O6jAaQenEimWRSf7mEymeqIl+Tr2jMq2rwhW0AMBkkpi8n14q8zp
u6GK+p9yliRH2unKJFLIYZzV7QxyRFSeFNBu4brHNHzbVmX0qibtcVsGq45vb/RO
609CfDAy9EnqbnPoQSPshOtg7Ux5vAspQ+OLYjb5JwI3uDy307D08egwV6M5rL0E
t/r6WW8VeaxSDjiD2bUMQkN261LKPXZY0FkufYXR86AiJbfjQacux3qaqGlVIawl
4QxgjrmiS7G6MGBMH3B/JmPCYxO7rbHwsZKCYxLRvup/IJ1Ukb7gso5zV1kOgWMx
ljvjMDxlPzN3wN3DQzFEiVD5F3Ml7sxkoCX0hHL0k3hQG+AJoY+DqiHtLAJ02zlg
q25mlBYrdVuE85nTyn9v9hSumBY6phjGtwIWmaFSnak5MyRg+lCnA43hCOPyeco7
lmdlmviYrjLl9/r34G70dfolZnwt+/vUnrYFX/Za1CTZJzTrQmGuMsi+ec9bR6NC
QbE9MHywQ+CjJEKIUz48Q/UhynOuR7YfAC7c2/C+JPRvP1gEy7y6PpUssI6LkOps
kMUIPO51MzeteT0O+HHmZxYg6ybvcFe2JIbaMpF2XKlnhPs9lkHdSdIMkOlOxgsd
6TDIAZHKGKMpwEHmqnzvMKqbU1yonOya3qrIng+Ihc6A4nIbodvY7Yjs0zeTxzmh
b6rI/YD5f4HPAviSabRQih+Tvg07EPkU1oixqYZqEJ3dx41MTkVq8+cnEvEokwZ3
4ohyrTemGcV6bPe+V3erjBGQbeNUDOI0AmD8/o4tCR6FYoNafW3CbW9PX3AAk4RQ
06V70fQcmCIXkgsENkh0HuxHS+9y/+8NJlieJWm03yNxrLh0pdCGK81W/GTP9AEg
dLjUkYFTg8W8X/QOigg29Xr2j3HTP94St0iKRuz6NdEOWObaS9nOdCMwynVrxrBy
Cer25hiOw3OUq4mVzJkCCRmGK0mmYYDrRHKfUH7BUI0xrHDZqU2ricftuyFPwn9N
zdYFZw61yQzMb3PTe7Fz2x+HfIUe2hejp7RUU8gcyLXxCgn9FHtrjZGbk6VqJtDy
CI8vrjTc10q79cCBk1vLGsaa2jG746JJg8C+FBnkOAvXZJXj6tzjMQkLK2CqTmLV
8jVMpuqwU1qvL0YESpF5OFWagcZ4XiqfdTvAfwGKwipPsLlL+RR0XcYdDML/uNz7
NFfAzHRfi7begR/Xa+G4Ttlzziv612Wz+7KsLaf5YouG/BudAi0Pk43AWC86EtFq
McCrO3bo/Qo+jiCpJEjw/WRplDKxi11GbWsgrfQberH+36PwB3AdicKA/jv7oLFl
gp6AH9VJTF5T4wn2H+9zbMUyaGDEIzfLdeHwIMJhDzBcmjCoDNtHZUCobHs4S5VY
xNKHIAPy4VZ2gY/RgGmUaq62pfdf7zy5W/wBq3ycsviuvi4F7t/KFGYmIS+k/djS
b1hwTG7u8eoL5UECwHiCrr0TastDcE0acaF8TS2cAbkR5r3jhyb91ZEHGMpclBYj
8Am6CXKouyXhBou4kYByyLmD07qTg08Qv3/EpJyrtKpHnMh5gHqKB8wni3N4Dr41
tB8f3r7LdzS8ZL8wUuMvmWKG7nlxWDmD2lT8DqaM8XToz06WYkjcl1+2SSQoLXsk
ZolayI8rz1fWqpkc3WkdbUuvL9xUFBV4DHBhhBkVD1o/QXzlw8HzKVFRuUY2d5oU
tMNC9TnG1dlcc9RgGlONrFaFc45O7wRMunEYm73cFn/hBvBjEVLStHA0qNp2TQju
7sPG4kNAjgCGgqnz5AopGgve1R8JLnW1gzCIpkd9IzjnGBeaonQDIEXpK9+mE7V1
tIlSyj0BHV1wVPs6dv6Sk25GWaRnaSTb3OV4Fa0pkqsxkpcImfN9vc/OfGdHkp06
GRbpXTC84zp7NB8d9VEFI2nsQyWyZdqFSX3pm/EUiEUCjZlZ93vj9rk6AvA3nEgO
YGZKQ5QtMJGh+RV/j2iGGgoaMU5Q43sjZbe0eV6rIOemFGFxW3lCPZ+UkJ21NK1U
VVZSkcdyyX9s26L1S4kASiSrrTnn7/b+dVh4lwnq0IWoBXtsoZ3YRvE/gNgwba4b
04kJ03o8J7WFT9kmc/mPzS9yLG86SmyLR+PFzk1Oz/VaOOgCbYvc4Taq0wPioL3n
92IrbDs1aFoVAch2qz430dPoUfHUy9TQwLEER8vw08kK/dM54ptnWZiFQbxKCT8t
kVSZGDwI4G/ACmfSwk7fFKo0xRmmW72u+xGcSilf0qB7A9ZD63J5kSb3QHhx0Ykv
8O/yBMFD+vWFmXYercQ3agzQpvcXPPO1h6xNF1+vy1eN+c/NOjkbBTGoDvkNf43v
lidtCEACo6lRjYY/z6hmjVKh3O4vsS8td9qD9Kr9o4rPefMU6VSbxadKHgyNjkMm
b6LRVmmqR0DduVfr41A/KechP4AR5tj3lVZmuABQV4h0vfy80iqvlw7tFvMDygxZ
c2ZFcx2EMrSkmRKIOkFlA3xl2S/QB2wpYxcQ8OVZ8iOhiD8K+o8LdtUt6CQ30Wzh
bETVQeDXonoTgF1H5t4xycmcoNV5yTkBtAFQi7nuREfGv5sgxnpTzW0g9D1CNFrb
KkUG0zQMJ+rQzTRddh9gICDcT6ZzRI1lu5uqq1RtptOpO8vYaFbX/ZherSJchaJ5
P6oliSv+nIv539/LMrLXDST0D1Y+3rPXjiU05aBC9PS+jcNdr5qjczYBR2KMmZJX
jN7wPxP1yfMJWi0ZSPYBvuU8DLCD05ELOg+rcNj1twkPTF9cr3gfXaspiqnhtw9z
+rVltuzVdQ01h9P+Ym3r3MjvEn0DKxCu6qGC0YDLXnY4rq7LlydNpjD0wt9HLdNd
Y05uWlUIT9lM58PTcCGYDGXskhwxyEJLZ4rOs9l3Y8+GKmTqNbWsq6UL2nhTvHtS
ov8xMw8wTBELkeBVbpgp6SbfhwxUYprnsA4iguMOHGijw4tOUgvxDKVpSFtuhTcO
APOVlqLf7ihqtUCvG5CfkXepY5QUodmQ0xmMtvXxcwrlrhtq/wmunlg11mHUS41a
8EBkFr03NruLBTXV25EwJ2AVvBmJUKeIlCw3+3NW6VgkX9iOZYsICez8F9ZSoH1m
UCHff9PnrLHZBNQckCPQCEd476epkeWr1V9U6VANAY1GKf/Cbnz2YZ4R942czkpr
Fy3adX9TRGPPqBATHZMaZzBwLemgdUbsfSHh24qFT9eTp8N04eaeWeEu1F2BGKRt
bCqa2ljxmCqZiEViZ2bCYT5YzKLdYeK+oTzcqsfT9tO/cEzJen2VxBcB1dsqqE3C
9g2FT1XNOAbIYEoL2TnXBl5yAmj3R0F5ylFEGxEBhqaZ7MSNdQvEjddgxw6hLucy
aNzXNzsQFVNq/TAg9H0HNDuNt3zIsCwNftUJ/MJP837EOuC1aY2drfJsDPE5nBe/
w/usuIK9M9SXgT1uPx68Py+YVtgv75Gm2suu09nTTtJa8DLWImLUDLQ6MHsuluOj
XotFPUDaW5LoVkRZrhSU29Da6RICP2FOX4V3OnmngLH6vCEMCsu3er4/XI95kkaR
IVcCZqz6Q8X6ucKKUg6BSIh5lF1t+M6zKFmQ3oJJeFANfCHf6qxuQZvQE75OnqRA
1UzcsuAChGeLBc2tahhOUsgC2F/CdAVzxX15lCDAX85HIA4HDrFfKN8Csqf1Nhdu
Cv1TovcLtDMs3UpYjM7y/1LyT6cp34/0UHIlbjqfgH++rIUoVyYNQtyV0FwT9g0P
U9lLFZgfpcbEjF3O5hYwY/pm/P+KGtT37iTd5r9/Kvu7bmxQQhKOsJf06yMshg4e
fZSMxktnmaWAWBlq9NEXRhctuINvCXQ5ZHliZ37BM4EX9B1f3+wRvU/YyqCYvZGJ
LJ66MvrbzSH/HBNRU6kRutGi55heX4XXfqrrsIB3F0yWV2ShtSUZNIcOaErpDFKR
YTB1aX5rYfL8IyUypn++MBwxW1dFvIFpf2qqBrKVefZfx7MZLlRoht0Kec5H7AtO
bxHot2/Etas0352CbKuUzebb+hmnoJ4/za1ziOTyLpwXk+AfJDRr5JBuXC9iGgwb
xxAhLpVW7r7xxgx8fbmDBFqIFkL7EWzXP1uHUlrfP8ZvtYub9otc2majZyCAjiVJ
fU+SgF1FQqc5Oe4JbTalhTjiWLQYZHRwrqEjICfWkAmQGY/DsZAZr2+/OcQFazWR
bl6yR1SDRwIbMdUMLDF6pK+M8momi7//mAN3z3/qS9lWIP4JaI8SDPpYA+unw8Px
aHFeq04e1Wlhb14QYXxUxZd/Z9Nzuw3+zJd4HuzzdrnEp+SOOSf0/+r9fcbdg5M8
UqRnrsyGSYVxg6/VNg7nvl4MBj3IemtIdjJEzcouvYIG7fwFVA4E9nBij5iTe8yO
mgMKXphrsCYeIQg85g3KJ9ly9nVPjz60BqA2Tj9NYXyYptxfBHByrCh5D4zKGDjy
oStYDoNvNqSK1P6cMfoyZvuMndtaa/jbaK/PhEOwfPHYH3A0fZ85jv5QTUz9y2po
CEEWkkKSZnZhQk2dYUove+mHdDIBzeyYkyqUsr9bhmzEGrnoUNxgEkk39jWsbFtZ
UCqz8UzO7Kt/TVBk8Z+6wB7ZvJclFuH2d+JR+lVRKDaAj5F2+cys/6R96EH3tH5g
Ckkg996REhBceERWm04OT53fmMXNLlmeNgAeXRGQ8/9Sl6RXmyfEG9tuk0Rf1rwp
xZ0xV1DH0FfQUMnRrYepCZmg7jbq0oIeiK0cGzzfDPeNEFDx/T5mD1RsCQ/fhVGO
41H9gHGjHzN6dJibGf+E8auAXi0d6amHtE/l7Z2zcAhxZXWBCiSiAfiTqRlrwtb5
UDTBwVbI4Uz2SJcU30yXBht+xf4DAwoZzKUoxrw5Ba7QoODdVKhq4RpW09skf/1A
4LOAWGowe6sHKe78Nj1CySaep9pEhTHMZKRR8xhvORbouGhEf6npGrwVWl2Y+cHJ
21+Oc+S9gxgdEN4up/fWbhi8kTKz7hvKLXwY+KzhQR6HftimgdO2WbbBg2SBRdN7
mNVc6KEuUyINmDrX3dN1TTJfCpwH6OEYSwYhD5rpysWVw8FYuQy4vLk8u5UXjGdw
sU4bX2hgutY0bSbpYbICgV7Xv9Pp14/hVkgqAlhFFn2QoTNswefQ4FPSPd/ocqcH
6RKuFi4oqmFqOuugo2WqhtF3OsD1DV7B5TVSaTaxFi4sU4XimdbduZ3mzyqo1Pn7
2PoKZCxKpe5B8TICDjZOoBUQ0A7lFUINaw1zZzDm2bNv+Up6AGiMFugfksUVgivI
Akwb7KejN6UBaYGb/V86WwZ54wRAj3omQCEGfiiuML9vvIG4NZXuvzHuE9Ho9cep
GQsPmUKlsUZxoPoQlf87NGYG6meEn5T0S3iy/I1qe3VgTjrMyRks3nc5FtzU57VX
FS1qLrdW12sxDDz5Xn7+YeQtOrlf3QRESuCWli/mh50aWpGFhSAIzAMK2UZaUQua
yuAYyi4pWMvvalrlTSJKX3MRTmeAJV1yxuRqdTLvU9mVRPXq62pDabNOWGHWF4AV
bCP048DBF5sGzbeiACzXsdsrA1S4Qdt3hXY7XOjST6NzKheOQetPtFJ+oCOoITQ+
UX/oBSBKxdVBU0ZFrYWiwPVC7soArZp8pO5xB9f+kKxVS8hjnbBbNiZnu3bKyBVi
pWoMPjkvRTundTYm/UR5kK3srsgF6/cWjn2fvVOLr13dZsYFmICez9n+imjmFo/F
EoNpeIAZAjRU/OlxzhoHTrfjinj6H6+OVuV9n7zkNxfW4w0Ls7/ygxu5jUo/wXjD
UoZ8eewiYJbLG8ofj10JBpADM9BjmFjItvDBonz0ZrzGWePa5nxvuEnNHmfPzY2f
spGbfZzYQyEfTY7b2bAeRBXO9ORXzSG2hM4ehSxKm0HRf3DnPMJzZjSXtrvUOMBo
IRsqAd5EWWAZ3YgEyoTW6muxlR8IoriCcOJdEWF3UaE1Ismr6T2sQsaBkpzautnu
4s0c3YpKcYMKqEcQzRnXhx7bARktikvJugiqwgs0ICOIqdNq/thPIJAVOODe54+3
9m25k7CzaHDkEAHzvK/541U09sZCsuPHhO+RJEa8hxOy444h+Fc3BNCPv3PLCiph
CWjRNrE+U0d8QplJ4dbyWm9RAkr5sIhbpEY1/4N1f2s4gau4mzG1qPooeOGEVT2z
5hXLLn3ZELnzyD39HVhZwtRoTAXmvI/y/aaYz9xJTkVc4vyLH9/tUVp7j3cfLWPk
QD1EDv76D9Qf7c8X5f+fIzma+KtXZ/CBpo5gRXHXDw3yPoVfcgAzrpkbSz/yGzRB
e9i2+TBfaz5nHeTL6oeP7o6npOumpR/U/7lI5iy9JG2597+uT/R3pm2N/SuYBtyt
IWGGGJpS2AZOThysWSoIuwkC4czuyfTrWv/ZS3B6P+3T1HoxxipcEb0C364ky4fa
tavRENBzefHjXavGFd7wR38smHKC4K1DFEu8ux6hn3guBgGSgcySnPX+XbMEUOhU
5YPVuZ4+0xtwSoSg1B0N2BSURjpp4uY9eiK86mII82NdG+SSkoMK2JNZ3QhULL5a
6oXdLvHsqm4OVa7lPalAV1PsGu6Ehvk1oh8qD1z087NQk4sG6sheBnovsPqTrfJr
A+3LNPjsjkRIPCtT4aSDf2qPvHPDli021NwqR97gMG0+lVJUL3rOtOt21Bzm95qM
+PFpAJtlOjCOkDTzET57bkaBuGCIHleotSy9O0mr/0LzNqhtkbTr82ptOkCoBhz9
V4nf8RVeSaIe56ydm9m3tKA8uGH75p1C4OiJFE+OEtv9AUZ9SQD7cqAXX8+6gH7c
Qn7m/gBuuSwTWBdkKI8XE+BAw0HhiVyhdm5AJx1V//1xniRBRjcOTneiyWQoKLkK
YcfRWEZKlg+tbBnP1qArL6KUrmUr+68CGN9tTJ0nU2VNQ77euOZ4zsTo12n2YNg7
1UCMWOzoXqHAJ/XCz4a3dE17ULoOgAMv2dpc+u7ErhbtzoA+E5xWQi2cu18nFksC
/7gn90FFWamThaab+4JuzR56pVrJooFTKTFoBs4JxoHU/iBeZIk3cq5psebN9BPw
14C+e5NrAXhiOfgFxYqtv7ZQfWDCi5RCD2fLC4Ce6WV4PA9pFFOH1u0ZHSIr7jMK
1l2T4NP+Fec3DtfUVFUsVFf5st+CnQFd7z0i4GoDENKKHpu2RVOFnhi42tZZejic
vy6S0oKcFKZQt5ACeWhZrJq9YFl+JqZ08DlyTNLpkGeEzyZc2js7Mr/rN88FEB/i
ggVppskxvvY2ByOtjDAO47uYpBsyHG+0RbfDdwKMn3/mnxyJ6J/FkRBaTQ7doBbi
qgl1W1u9tVBbcB3XG7CnX2EVkudW/k3/YbBZysCohyGnt0qvc30zHaOeHm0YHpBr
kfvm0ksb9o8or+tDDdJJrPrk2njtU5TQavKE+teMhdmmpjofKCE+16cKiq2e+E0w
0GCW1+EmMbaiHarNCWRZWKLvRdI7sX1IXt+Irr+Ww1Zfd8LEjs1ZsRJ/SHAb9jHG
P//1Ac9wNbRS1QnjnPGMAQKy+Xs+8OGHZpEDLA761kNVa5frwzo4YURPZsNDXeo6
oaMKhj8STM3ovoWWhh6W8uews02h5F0+S78uORY+hpQpCV9St29PKE1Vc9OE2OMu
qzhdARvSsNgEQesEBMZT+S9bFytYkFeZdUuC8G8LH+OUs63u6djmAwl7WwH6TvMv
P3PA17bPvjst7hXVdzzYWkoyXzbXSALFc6pukz0j6d+iBZR1oF7Qzq+i+DzGsihy
ZtvwwWyBNIdOkrjb1CKP8LENyq7e6v9povGTv+CMHvO2UFY2Pvbor6ETCC9BmxX/
XnjBiNnIDfiTio7u/coTFEuL2q2F+49b88wLAMK+4HLcnF3I98Lkcaj3aI7vRoNa
EfMnhUZdOoIr24gL+V5IwH7C2+L8XRqwI8NIFxH+8oPlO9PE3RNzpj1E4Ly5aIWq
QQkZVA5gBEjqCxmDITP4B8eBj0ruiME7v87HeEF5S66rEhdf2gJywGuwoN0BHAej
lNJLMwnyAEk3wHINMKPJq+cY85ermuMpSXhWKNxe7+dS/M0hl8SRd9CbPWoXw/TU
Be8IMGWme5/gmHQI3Mhy5eOkUKTrZapnUY1llZvS2UAL/Mkgr08uzagbMZ6sUvD3
mkAHoWRSx4z4D7m3DJW7cHdlvM4YCI/KZpsLmn9PrQHL2apxnZ7kExNb9eQ/gS0+
wq3tyS/9EqzYIhJ96M5Lx4yK2ujY7H5ws/3fm6XHbrnQBqk+maeUabNz/aKEgu2C
kf970A3cU4mk2EO37NHE4V6sZEr3MlTNnORMySPgIRDx7ST35U2fyRpBalR/C8zd
nqCtBDY2SFWVkXtgSZHA7rK8DH8vo8A4/iee3p40qi9hb7IudUWcY26Eg/Fdb6nY
pT5k//zjJizttOU3IQKuD+evSgPPBMuNmXIlfuBv0SuJD6VnvKdSsO09hZIc+aLM
gP8+1RKk6e/FA+ja9YlmySWir+I5IBaqSYb31HStolu/udlj/G7FCfUDn6iocEsF
oGkWYx6Zjk/7m3cJ9FevAEf4taH3HJbZGqnPmcWVHxI6IeILCqu74KtD31BsyIpW
1MM2cXLJPGXShWbAotDX6BaG+MNYQEw3uaaYHfTUvfA/nhKhHpFzaNbxRuY34mf3
3sMTZH9S8iyzajlGJMtdPSYLHFkKgvBEPLv3c+JGGytlIUnEMwVCm9GrV3BxfG9Y
8r0CmMrKK1Nvgk0sI5fGeHfSJVumFnfk9qyj2FFSQlEEftBUey2Nc5S6h0e+9SkG
8ZShTuoeXZKap5UGCk69buUUwsePUN9373CpkNsH9BwlIB20uu3s2iPi8iywpCJc
OeoNiijKQHk6MNcdiYSEyFoldeOcGp986/Qsrv8dNTMSV93bDRklvMPEVX8wJZuk
u8UJKxh0IjSbyOfx2cs6fI1hyurQyZYgbE1d/Be3keOuxbBRT25BqjJs9WMQepxl
UdBcLE1umtanMWZQBW7p9rYbXB6cR9dnpLaNBtEFti6A/g7qpguV82K3DhLb7ULx
MzmRJfZrEPQZcxOKf/a//yr7QP+BI5jgYmBmuWuqxu486isfmvlZdn31LdDe9/Zs
gRs2P28MwpZLrGNyyfb8EpbJtypBqtCzjCfXZa5WT/l7kZBOdapucjJskAZVtrB/
JL2XJSUTCsUsEuetG512VDec5EeqmUOxL0exNNRnPq/h/Jq00xrx93aVGQ7NhlIE
sOR890wdPgK8RzrocS49s8QAE5JBM6SpNPSfumYvajDgowdqVk2xbOheyl0LFv0e
mrHAlfigtQxi3QeGaBI1nTMNC5a+BcoIApwoEL+gpCdbglKajPBoX2j+zCQtrwFv
ikEgDAMUZCF/TaPGZ11h03yv9YZVPlJOUgZuQ1LqJCPAM2mbwFVSllYxh7Y3/wrA
MArDK74O+9TdaVX6bHms8bUDVVDd90iLyALtswKmZGde5TO9sdbBAJ+sB07H3d7V
2SkEyT5TNMkgKFFkC1HmDQX7xRPgiIcbNPwxXB8gOdL6vAtHUo5iBJRyMTFZ+SU+
91+DHr9ACjoyi/CuLCPlN8tnU/WIUjZtVj2UJdnu4nKn+wlmR+TVJ8R+BQKFEjm7
q/E6AA6di/qiOmW8MhF15z+4PcQSKVFlEPruGsGdDYPc1BvxpuBQ4UCnD/HkYZGA
sBILO21Tqgyatqgdz7Feyhoz3KQ6iZfvWvLy/EsqBTMeLCsHiQHf/nWyhtSzNMmZ
ugPULflviCaRQEJfGLNFcQsas1unii6lA9l2J8dMuKj4S7vzxRRQ7e3ZH2ipIFes
QUVBK+4g45EBewugHe1mZclopTS6AtK7UyLhwf+pQ5yf7Sy84PCmTChZlg1K7+/D
zb13xsySdJc3Ab/SPudNHr7/p/HN4H/KxEGbx3dNt5haVgIARTuW4l/kcElDo9/5
+zm7GcXhkR4bq/kTi/Gj7CIRPydxqoPMWd6I3zzhhUH+BdEA2yH2XOWHLbBnPQcT
lgwXZehhUOhHtXIiaxiKNclsL8tTe438y8Eo9PwDyemEI+u+Z35bJosTGoSgkmY7
ajQd7qWX5Hwibi0FHfUFMN9SzhIKgRbugvhe810nSPQMNIgzGfDd98spBV1IvQsH
fqPYWDgHNNYSUf3ptfL+rxMcjDCyGfyo8Ac1dFUzmKU3pawYcVR8Cs3l5ldK2X/3
iRWyO7Me/ozOWZhGJUhZrEbFQkAI2OmMolwGI/PpSv6NsX5jwvSH/wBOoTfpWLnK
LTc2u7DeAHk2JTNQIyN+Yk5Y06rqxa7sgxXiDmWWYtxSyNJPCDeDKuETBcyTriYl
+ETAwzmomOeXun63ooUkLQeKozH28ijCyOftV1qE3EUksoNfcXMJjtNkPHP/h1aw
iyQuYqvZLopouS9RbuOpgnXNdDbQsD/H67gLneUZW3Pvc58n1UXriKgVdqku/bEd
+hcm0Mb0v+Z0ZLd5dVvfLaQT8JVWrFRQaKDNLVLeOHoHf8MlLMrK0qfhrV6DFJ3G
b8DMtNGZONMYrve+RsXHq0r0IAgSXOw7VTGBF2eiNyVnHCUd1GHx8EQnSDC1UQ5p
PQrXTpJ9lJJH009s4DMMG5o8sS5oR3WA0laiSi288ujsxE/72UMEzRH1Q7qx8I1A
QvB+wzVXr9j5I0ic+WwXsFVfpR7mTBy3/hxwA3CicIlI9bF1yVcUiadZZcBhXSVP
YwnCbIDBLKdztn8GqL4IyQz6XeDPxHJAVNJ6hR6oqZZ6v470cf2ubv71cvEOHWcS
y92Mm+GEyItMzsBMgPKqZqV8F9n6bh7BfJgAXinthh6eC/JnmIYFkc6ZTMuj79s2
Lonw7Sf4bw7v+Eu/WHwmPZVFsvhGlzrEaoUBdtvXp2rTAjOFS6oah9o1MOF4HrgR
F/3N5TO0XlrprKO7kuiLK5oqkioa38WvMin237rdB9auz2RL/tYqq+uY6ptEoqyT
QqTkah7njxF9lymvIT5bfiLC+JtB8YxVOTtS9or0EiyUdOsEUert2M11TRZOHUQD
5LSUM9lkaPSliLLT7h2jNYkWSE1Twfp4hnBU1NqBY4tHYfWyDUGG/EiDpdn5vZaM
Ii85/SzI8WjycYozJ3qsVAr8EUoWUSRSaQ4+NlCbqZZEEIXXIawuuJsjmrFwwtSL
7B7UF7SNqEPFhZzgUob/x5VgSl/CQuAAsvixLwyukp7pQwyMM3hAZ2RScd0VsXUQ
v/0pWg51Q7bEyRdDLn3JbIYZUWliG+pYqVm6AClDuI7eiXwJIDeBIt7d1WJpDGQV
oIjINKAvDMzeLZSee1tZOiqNEaVfewmiAl0Z9mp80ZnpGKO7O/IhBFNdwfUbdg+c
oTVjUmJqu11jsQPdZP0zvPK3gr6w2dVA2yye5mWwPOi9e98EQgaoou1Iqib//GrZ
aztgebJQID8+YDda7YCGOvRMvhxkRsFAvoYeSHF190c+4eJNqyaoO8PC8moB5MZ2
BICpCHAWllNATCgQHVn2q7c2jKWY2iG+6b6GROd+eoeTbLdjHwGexLKYp81/OqO2
T/pb8hWOBGr3pH1NoN69wnROOGoyOfNQBu4DSJFPDuEIIZ/4NFZ4aAi5Zj/gaSJ5
+324oFSdlk4Mzv9l7NBCKw7IpoEJKZUgit+AZgU+/A2Y/sU2xb61XR2ojOMvcr+p
7vKe9Iu0cX9lc+lElPxP6vZyngI9DmXzMzpJfu/H8b+Mgy7igQle537XaVGpJjvo
8T7YAdfiHEf3xjdWIFa3K6e3IA7QpF/GO90KrjeupaXodv75ec5LlCKqXfBrsjFr
SoyDcMZMzLu3If7WkQm1p8FnmhQqOOubG7myF+osqpB9s6J03D6ZRsUrQN2wkaz7
XdhbJxGcYwLQ8Mgv/U8yHB9H27qkCoRgHeuKW1+6c3w5T7G2eqEQz8nEBI0AYBc2
TmxK7JuIpnqY8Httq0Pad8DNyqRPO7izlao8if8hFT0dsx6lwcP4NksW61zGMPmf
L3IwHTonHoW2YenGpkEOju4vpcllTq9cTxDZSrkaSR9K7exv3qRPMPH4kNUA4Tjs
skGHj8GVPkCvNloVfGJ0RDXmujt1PESWfUMNIIhaAMprR8SEmQJ6cFxAjASmbrGf
xj2SKIXGXttEDmO2wp0Vw5WDg5dyM0RoOudYs+cGRANWNP/xHqlQ+jIMUQyBDn40
VaYeNC44to184s783W+iuvHpffrCvFcDxhGrx0jRy8euAuvfw3qz21Z7/gQPW47J
fEIqmSiOd2sK9dnBfc3wqiQIestvfUkR1BZL4QSDURpnMb7D3J3o9m9YFaHyU2IQ
R6Ar8AhwyDgnkru6jxfa2u3kpAtFb5OBq0CGpPZIiVu3lEqLYKwCt9kDiNm13bZ7
IQq3PhqMgb4suOLGasvkg44A7cwoCjByX12H3VZ/jNnBV4OhaVSFVSXp5dVZEbjG
h+leSkNSnlwTKi+sWOodfJGzinwncYUkZaUa51n7rLsAjhlNhClIYOOBwp6JMJn9
RTcQR6RZwJ6z+1u92nqRiOvVQbxuzLhUXHQWo01BVTzR4e0/MF3hUU0aJJru63V5
O2LosKiuYtuoq1eY5Uw8uP5cALLTUS/bf3FGeewt+wTNziTrNmtf92J5YhL6d92J
G0c0YtkQHZNedPx5kk6P389Z/xcdGBNiv1moMOhIDyt2E9Lb4ZTZWX667ICthwYu
JUQ9Vk6LSZRzdwy23D+xd3XAK80fddLxvw6I2dgF4Ler3Y+VHCVJ80TRGb6srnUo
ExQSZTCcvJMu2zY8E22rAIt52JgLVy2HAdwSk+5fO+t1Aje1W05cDTJmniEWtSYK
9QFDbwpN45lOK4uKhEFWbgQm14BOLNgxFmfbcrsssOAOf2Vvwh/SBuUk1fHMaJap
r12fPIDfwvdzauCGrTeB4rTQyhJF7ZV3Fxm1mPZe+B9DufmFSiXBkrkTXp2xbb0U
ceeuAPXb/l2PZDoRFwFDd27a2BQbWp3PaaJJwXKQyIUif1mZBQYF8AuquXyUbVgX
lOKM+2eo0UDw3VmMyGI1y5AOiTzBZ4JimJto0+rOBJxWRnwkYv75fjiswZYBVwB2
l30uzG8CTTbUQzt6BNJk19xbyElhTNSc6jCCjgSr4wFfaz6YV4py57lxSpbiIGQH
WhMm7fkn2diD9KEA1jxgKt4zXi3LPbITD67sJL2Uk0C5EZNv32yYBBxcTuOyLzzV
LaYJ+IhFHZToZGX878jlCuH6MP3xjusfHIxY2K1NevNky49glEkoUNMBUAWJ6Dys
RhgNVtCrVjdy4tozWek3sVBFbpGOilmeO0ZaJ41um2TPrApsl76YnH68oGjKevVy
lug2PSfqvLMiPihKP6jP9Lq3uJ//Az0+YzlUc8u+R1Etk1kSAN1y6pR68m9DIgM+
/oS3GvIYtO6s277IrohivdhFv1yYzsIunfCLjt9s3p6TCCLRo5dMYnxAYtcxqe8o
rwp8gDrYwnRego7aGnD6RtjNchgj8Q16TlXpLYtEor9yIrPa5aIzndK8EBbhhoQM
aOjO6r5z+M9ppqQtsw8EY9LyI0VutkNW23jdUuO9OvHLLrs48iIyct/oH5VI9rs/
IW9Qe9O9bD919XdIaAfeti/kM1XoWEzJGAwB3+5ztMPhkGJvk3RwsunCArNLk8RY
JWKKqNH6C7hfb61AoymnADstC9Knvb7e4uv4CC6CbgDc+m1CIIbQqwG5c0pxLgpT
c2vxB4u7hRwPMrUjacUcwQ/FoNIgqyVkoMJ4JMzYK5/Su2KspsYrWUXBVAd3MeHz
u75egoB0TAmQRcyWF6fRrcrGmbOz0E752JhmSZdQ1CTRGhhsYX8dUti4ViNmHz07
DPxEkCEC56Z9Ev7AY3uIhxvg281mtrWtCjy2dl3bA9u5tHiCPLwlEdmIaD+AUjCh
HcGxFrSq0Y1J0+IpTGA2TglSvfiJA+Lx+NrveVL7Sh8Hf5EhpMCxTvdYkr1PWwi3
tTblyCXf9gFKgiqoIuAbWTEcgnW+LMoVSh5zqbioYJ/QE303Kqj1GKxNlWrrYQq2
ShWGWAogROuotKVHESwpo5CWDD4Hxm1MJt5ThXLzlgktdXjONZOmoD0db0r2sotC
hbfKd/z/0twtWwd9xYmCLE1cSwsIxzelrHR2YTcN6563HddnSqSMdCEohwUQSwbf
PJg1XC2nnR0DQrwqFs8xXDjoZVf4gJN9tyIFepi0La8RTBUcfg1m0esGTWP//opw
dE1+yQRiEXP5nzdnknBJz6Qx6anh7hVxZUfKM5unKE8LLqTi9w5cEoRJjHGRidSo
oAOchq68hzKkKeCZGLPciULGO3FrTNheRPt8HybI53qQ+eqq5kU+fQL349r+4Fv8
tmZCorrHL71T9ZuSogi0d0ue7j3a1qmBXHZbiTeEqWAysDtaap/MGIb4uOY4K1Jr
0gWtK1BPUcx3oef0rlLg0OWNDQ2X9ni8Rdxlfxd6/ZknyK0SYltC+rXhYKS8ZFgm
3DLZMo6cSHXJaY4nfe6HhrV9m+8+DWgwcH79sxp/KX9ycgHrHeU1xP248v3pJG+D
OYMm5cXf/TZYCUoaXggGzcfl4CD4rRTJ3FnmY2V8UQ6dPdmdgnn4KqIqWBxRhH3t
GYgICrn9zVQkaegYOALD4uvx03Xmj+B8gxSi5p8EgGl+svhyjDMsIDo4OoN+E0UD
ffyCOBQhzSsst5UTPGYKskHMbmFjGQ7OIxlIwhMoNw7M09zYmg76fkGRWuEWPyCn
FMhBBCjX4441HgTyz3cbZUXH3pbl8WXoUU7ljt5FjWl9Pu2d59OVj5G5/e4Nmcsg
1rOQvZQVhnUDYvzUfzx7u+NBuTtQZuj9f10l56ZOfYhobY9g2qYG4plUjgXyGJes
/1KiHUrmVFK4LTqzY0Z3HqyOkoJ+B8iWtfcOEqDyORL/pObhSRGYL9PgeOHNElli
KUGVMkrKFrs6vpj2A+ICh7mqHQY+RmSbKrZd62pcqcVYWtfZccqw7ZN6JhPmFIMj
o7Ydxmxtyfapz1A8chk1TzYBpH8ryDvl4ErYoukFz49LBCGA4It7F4HQVhGHa5P4
r+0dt/mxHMO9FYeEjhEnxRTQlQpEXe6BX8rohfl8WfVNwYIOAJyXurxbzpYchCzH
1IzU5TBbQwQaZ4QmZ8eFiJcrUEHgf3vcQ3VX+kqG7KJEjNmI35SymnMzM+3pWKNa
s37KlBxkz9L087pD9jqjKztSLXQNAzpBB0puNIb4sowKWG5LzZAdK56YJVBo4ucW
3OO+aWWHbOe90P1aN852xD/8tSushAJ2B/5h3knU0TrwL6t3FfjRSEDFv8nW4V8r
3U6Gqm1TZ0soa02rxXfBc0aUa9p1CJFBvJyCUaDyOtxuLim1hmsP8Y252y1rQ0y8
YkNWSuh5tgN0d6x4nP8xk0XHczO19xxYyX4Nuq/dhGlny4pHqL08lEiKsGJJxVuk
onxF+NCQXBCy3v0zacZzNr+ftwJqgX2ZVo+5rX0ZEDeShu0KWA7PjirlTplXcYMD
XaM7+k2cUmWnedSpGfsXIlr2CCeOcldOzNpSmXtT48oEfhiVxiYcudvnyVyMCHFa
pU0TGsvY2HueN4VS096jGH2vUF2CeakuAiap0Km1zuJPUKq1xpmr6wNIEIzNDGOe
csOF5gqxLRE52TRLCRYqMhzfR+kffjmQVxCeb/UQKuVSV/tiPS9YRgBibJVZ2XPm
T5ccga65d4vV+KFGf1hWaOKD7SQ+2QtTNdZQ9Xz28ud537pF7rZyC/iKCWr5q3o3
Mq4NVkTBp24xbA5hOTrDF8MqukxzizucUyJCZJmk1rmTMkNT4q2VIqMTfsLndtZM
lW1on0Kj7Q5zoP9HR1sBvGc4WxAA9pZ3Vr8CFtjizW2HqCuOI0sK4KUwL5aVkTK1
EUyFq3mZbvhkSOWnbslECcpcpGdwHqJaISx6KiFfwSuV+Alfc+rUjwFVI1LV2F+j
5iRm5rGxmk+5f1+lG/IwNCRS5fNMtZZ+E1cut6kRnWy09KkRlOD4L+EoslQ5aa53
n+ELiW2VrYGY5sVCr+Ngf/NUVzS5mmp43d+418BgaSCEz4HsWwnCQGORB16n1EjQ
xjpF31xt424Ys1yBIOUppt+ubSzJ467sIw3ZmQkCWANdfA7qlBlyw4E2lxfQ3tSl
SgTNPtRyp5e1v4rK5h0vBwIgoEopJXA8s6+qqRKUXP278z6nNUbpvKFohlI0tB6C
EPQDOIxkBRlq+tc42O2qofA3pCy9avNXNmbC6G33wQ23ERPtgsdahVXmazd+cTqo
aqRRNifMU5Lvs9Cj4443/v9wpkYhGJFaL4thXAJXj0PEbfJVFq3BIkP0csP0ndKe
SxWdurrfN8Nmz30jOWBV+Yfz5vu5w8hUnkC3nPojJ0ujuXWW5vc1Mt4Rxl3nOSnN
K8ZR7Jsaoh7DOE4XUYxbNAWiRQshMlz4VQI57hEROewZx9rZ5bpmRTXugHf11TYS
QJNrjrPAz1nVz6ZzlCkGgTAITVcYUitCgGFSJa5jIPSfsHhR69UHPXHynxUBlo0q
ydMqF/lWrjiTFvb+1xLTzEHWLtLPsmnurhvY65i6kiP3RgKpv1rNAFuW+N9n6vku
orqLvU1wcdfo36YNL8N6lPgyF50uzx+DAKR71yA4vHkvJHfL1u9AwhdBKJXLzrm7
+S51xpe3Z53MkAUSVttYor/fgqnPt+0K6rTZpqsxJotSxf4ERpAScPOZd+c+txD4
G9B7rq6tXwyosOVOoDaDTw8DV1YmS+AtObZvUCXhZVgkHz36NoHyWeHbQvahwL4U
ymipPexVkT0TWy9k+C+dcUjAGA5e3dBr2wYh2zwstKTmcoivgZ3PNAW3at9YA95+
S5uqlTBxwCe3AmIkPQWoR5QxxEPHrVqkY3wS7oLst1RptKl+rrMbrFIz2YPhuVXP
2MgqLsuDTRjIB0KewbrbL+OsjJDgGKF7OcsvfnCCh9R/GOuXQ6QbWbBD9tPb3GFs
TQZ4Jh2CTu0IFTpcNW7IPRhjHODPP0ppaxBphTeoSV+xIJxzR7MJNrAhg0owD0YN
C54UkVJlOFjvbBpVUr1IlNQSm/aQlp/TdIrjdsPLnUW/5PQU3pOmTOK9nmDLkF2f
4qn07rP83Tq4cVLrQ8Gvz90EPfRmJk6tQpnjoL6wjMpcRONXjBb8lJtkFIJr/3GA
EVTF31JbblMIDfKgx+IDKtX4/3NaPrkBc0fMbiAGLJd5MK4OT8t1MxAo5lEI9RqW
vVDar9UqdmFbCGHrnJJ5/Ni95YtBzfDxlxxTLDpVeKJLAxRgOU9ugaZU+dE6a20a
Azl96EStnGiQ5pXiHFXHyN9granHOgrp6nKuq/sruRUpDVbxsoijEHz1bQcfl22B
QKCj60KJxVGHMs8DpRURIPd4+r4Qfco74qt9PsvyV3LtLekkLcpmkK6go497sOkK
CakwVBv5p1D3pEyCNsbd5KdReyYmVSrVjqFELLjtw/6kK5svpdt+StCe0bULQ3aI
aXr+5nfnuGx17nX25aSOVZINQregB6SCCr2Tt0bX5D7RTRZ1U/jDsiN92oz+DaGq
P1Sh6x3wljkqWloooJQg2mW372z4eC6Mg+3l9N2gCLTVGGhEba1hgpZtVbDwIAXY
hNWhSRGhOTYPJDVKgvvCgFajukZ6TNTTlzWTQXkj34xkxrxIwzI4EKaKWOwz/2kA
JapR9RF26vexXKD4d0oPPn10cV8PQm9sLs1S3D2xmZGsVNE4A+ZNIYD8BmMR4uAg
PqU9VMeeAtWTc/+VN94hLigmNNggRfhsDRQDJ+tzoER6YlzMK9swmh0Sg+9QssOy
SpCMBwlT4sfP051pSiefWC9FlZPZTOXK41DmsiMhj2AC6UgVtrPQkm+C9EP+xa/T
0LtHte6zsjXYpGSYZaQkhWa2n+NLHLfVpaYokhR1EAenScXfMpLZihF4SiAi1i8x
Tb3vhLfIlfHTk3Nc7n/8QEdlfJVmw0HZvq5NLQNhwzRO6tTWZ+0Mkd6a+K2fjR2C
x6SlhPR/+HyKENaiCkjnDlQWuUx/qKGVVt7aSJbCjIzZPd7Ie77nLOgS/Vz4Tcp5
YXw4JhcLnhMcGwuJ+ZU32OLNvq5PFbpTSiPkpxcanLEZKx71xvbv7fe2KectWg/6
oouVDSr23zpf5oJMZSu72UpnaymiIB6zqLk44Ffj8w7Q1u4CysrzzkJ1zCJSgTGA
Cka8A7BsP6woOQAqzpTHXe+dmRNuXtgQj/7s0mTcwcTiJlWkoowet1gNqHcV5mx1
sIz8X5nwfAkCHvFm7iki64NQFgAPtnqxv8Gm8+Ea+oAw4TuRI+IDM+y5iO938XCB
ZtfYNmFfxI4sXAVbL7Bc69pjuljlupzsAn9LaaBdv3WlAw7jHxylTInOApRiwejQ
8hmgH72FVNhBQt48SkM95JYQARpXqAk+rlVQjc3y16xtt9vxW2zV6hQDqnFF6S6M
u9DC/ZU6MCs7MFDLVvjmDokHZoHUTy9P9fBmlDepmaapQRRLMietOkNwtBck1lW6
DyOSm4LVBepzT3+SnXOSQbuR3OImqsVAt1RPToMJ8sjsKyVptAnP2bAeoC9opAj/
8tbvNetwNKyD9QWG5VJLLVv13JpCAAfzL8JdV+RgnuOQmPXYLGUBnX6R2lOXJj/u
C3fE342t9ELd1mMAOdi5OcvPzCSXz2IzoCNZAdhpotrInThDVM3A/PNQQzETIVsI
eawDv7ya6vNGsWdlV+jdQ0QhMzrkFvvJZb31EHIy1LHdXGtgk5VZw/xu/9RJjbvP
GxzFcU4iLpRwTLN82ajiR5K5UnvhAzwJqPGC4bKtA76N5k7xb7AC4zEg60HZw0iA
4Rj5TZZBWmN4IhtlOB9T+bVRyCEWGy0IC2FXlj68hP+/qXywkao++pbbj51QoRBE
gSLbMp5Yo1s7V8Pp14sh/aiTq5cq0jLxVON0GSYtCOjWKRNfsvOi5306oI/C+RAs
b/NiVLBbcubJoRsedWjjT2xjAQU9Gth2RMoR/Phu8L59FJ4FimDALzRpB0RqwmNl
lAi0gEYH5rctKMWE4nyfjm7nUezm390XJIqbABPEAz5XtrYBCY9ziD9AB6DVeJnc
rebSS/7zLGfpduzCpLeRvJQs6mb2QL+SP2EaMQeB+2VT3T74p8BC2rDwdsvsSx69
kfgMb9XyYFu4/cuoaMqqEtdwIeprViLfWZKNeuImaBGhDvMmLwMaH2yYJ8ac/3jo
pR09loBMKxGFeHW4AQjbl+lKHpLNP1K/QIRxnK3PRsMpyx1yIKYN57bw2Wun+tpk
hdKX+yC7pnUQvRXgw8GmD8IRsCBq2N6NooVmub3M5riCw1MaFuMgDQnDR5kmzI0q
lUiA4/M7//BcZ4iuW6TgKEJ3AmaoYm12Ez0QZM1j0E9PIGie1wIVvosEelT9hNBG
/lCwDxM5YJj/qrv7igSXFdOjqHP+BBfIOC8S5n9wdhIZ6F51iNtF+qhgKyYpuDKp
Uhd8J7SKn88/JxiySX+s8NkTgSkL3iuxqoJLkDb9Gmd4X1kVrBQo3aVea5pacg+H
pfnOQxFCVoMwSzNt0mu31NmRqBUptuE7Ecar3+NUO5nSI/DsskWORbEKSWxKrtoF
ijUmSVKjipu2/CIUNZLZ68d0lVKWnWZE9EN5WxeDPjTu/Qxk2B4DqiKGcVlSkCA/
ZufSYLwRidNjghRYk8VbKAX6YrssAsd46E3V92hh/ikuRsxt4VD/sskxCOalfrRI
SWg4cxxmDTkR2Hq0FyCcg/K5S9GM24Ox3gpUb5fDGGMc7fL44eKhjWk56XyHU/i9
ehX/Awyf6cfAr05Absd2nUTu7s0gAMMh2BVLjsIdL26dDdqS0kRlKMbnVynX7sVh
FUXDOw3tg+GQ5HH8q3kaS1BnT8H9LPWZM1duackheJV4SLYzN62tQ7f1FD8na9LK
kBDL7bzBldAkMxFIBwNEhx7Yh/i+PTPnCSBJ0uFNnwO5d1OyCCxB+y9TzyDpA5Sk
QiBuQPnz2kztIl+AliYW8zh38IxOU6w2U+0PdLOn6G1NaJUZc/xoPVaZDTP373IN
sY+Ukc2ZiDQC1yD8PKwaX8nBnfVIKNpuoNlHcirCcW7D7TSqs8hPhicShlimSzO9
VzKMNK7wuQpadF/K2kFZDw3R6xI11SeRouZSVt9YmuIlNMENYCOaNWUmEIn3wil3
zw0hppecAYPqKYY1lqQ/OhQZPsBAreoWkbDKROdWsbd9NXeyJWo2+6DmaQSHtLoT
WaHamKau+OCi+GI22zEalUwKo+7zaX2Th+X3f5RgRe8f/UAuMYTzv9KjOcsXkfrt
dXz5xL4ZJU0md+00fXC8Ky/XSfsuvYtrcCVn3BtuLBoUhEb27ZWwfjOoMAO74yaq
eSixWGSZeZaA1TFNnJcA45v7Bo8FLfMTVbXopq2fjWpqMbSNQj11FgjQipRA92GN
JoI+bVOqLXBzt4phVCy7SRAHeHatoh7EqUxewgL/Y+5lF+FOAmrtZuf1UZ0k7Oi+
qRtjbIbQkZAc46XW5wr9wIoBxPX82Qpehi/LYoXxq71s1LkrUyAEjBfWxMMm2jZy
9wpopWBNfOLBzDCcjKzAP2umwABLLuW4smGPyY/PuYzaPwHfkpeF97Py1msqn5p9
RfNgTd/IzzNryo/AKp9I1S2EJ7qEIwdakZ7CwdNyFwyVDDNi7Lz5D6RUKCbCoFkk
LXqenWQ4+Rn47nL4du1KiChkuNE05LgQ8KaNqA1Gdu9U0Lh0SRAJo5Q43/YBPM72
1WHMPk6vWdyIiju0uhfYb2tZ91bujixYEPV92UEvjYxn/Srcc5U0Fn8Zi3QaeFR4
iG7107gWrs0t8f6L7YYtRWSYidGU3hoWOssx8ODY7VzRwiwZ+VBCAAodydoclYGy
M3Y4rdCCKsUZmdniu3O7yF9C4TfinjqQDeAzTb7iD8x8+uU3UHs7HjbO5v8xxMJ0
25365NLjCyI6zd2CnB6ak/om508XhBLchQpm/1wSmO+CelZ5ESs2eyE2pThmkFCQ
QvOTHK1LkZ5ynuYYAxAzdT0yMMQz6iQ7ZnbqNaykU02DtzdiW+ZDCZXE9ybsMsfc
9ax+IK+pqoh5uouPAXadkV9CdSfqIU2QyBeGtUxZs1c1wXhEQUzFsVXyrI4E539W
IvJjbi7o7sVkh91HTs9GnfFNiIyZVmyQ7/uBloPUIy3xpmergpKRdmwvF30L0Xlm
iXktNrGc8juRhZvLVmdOryUvq3AHzUQBMv4OnjWvwJHsBiYGkehYscjAgdGgOb9H
gKZZMLBunJP9QFdSWuytIlpFgwqArNi6waj6o/wQCqy9t34qESDkUoqR301WpeTw
nTtrXnhzKOt20wVcBQt+T32Dv1tBbeFxqmuJy0aN8o978gc28P9VqKEF7ZIcmShQ
ft5JMAKeSnmxtSA2RzCHsf6o1PCYvi0+Vx6pjiuudMq/oPPDgDBwOxa67cgoJtOe
F/xZjru2Ain9JlhuxjgF4AG5UNomOkt5/MYUZT2Ux//SSqIcPKuDNST2kY8Xyc1n
5QcE8R9V+KZkscLFq2Fnx6IizvTJlX/OnP7rcgggW1eBAUzw99apK8W2hNsAhIAe
ELVdrlq5XznuZziS8hGIUjgn7QYYTIqqlJ4HifQiAF92nPpobEJ+6MtzhIMpXZwc
3YH3CKo+O8dLSt2ZY7Bqz0txcQ4qrm8KwykWTOq00eYG19MKhv8coSl1yaJgmnrg
0fn/yDdiwA3NZ3/rdbCgxIthnGhdNvUzlqP0fCp3nudeqXvDNhK7iC0k+Prmvm/q
iHnISTBcMAHSZi4rn2Cb9mp47BQbB2X5M3zh3DCE0X3PuEXbt81hGaQYiwhDPjRL
8ETPatZns866zX6ZpDqgfxOdJl9HpVsSDGDWAs5FR3ICXe5QbrjNjLBJX7MvrTwS
E+mh8RcWhwuTxDI0IsohTMfZgaIMnRKHIgCNHtL4KGR/sVhkxdt+zBVWZ9IUvGJ7
lfyJv58YbTNWiTv8aResmHsGZ40MmbMh+pW2ZSaEOiUD2E1LG1X5tQNA2XY/vaOF
uQIkPmCs8yIx6uECKGjKODgfTzM49UpzvrQHjWxZyXg0qtf4X9bZ2kjCnMvuwfzd
9SxYM0W4wPOWi/rmrKuu6jKqqjiiA1940Y9Mjl+FZatD+MbE0Du5Adq4UqU3mJAW
0uCBmNKD459aMYn3ueYuhjLfexA4bp0E33akpEc8AntPAYfMcOUN+eZMLh1pMpkW
Jdq9B9VtVUesv8pn/sucbfwWHrirA/kYGlfuZJXTu3Eanp8lW2oaunkksxQrzu34
2+IwHdob7p2fffWzD67EdHY8S9LKvJBjeza6akcDGYKTnQjo1vylrHxeHqUUGfjY
PLeXuro7M4DGFfbgxnMxM5QHY8IECz+eFIGLZjRXBpvWPJnS5hF7rzWaGi/aFVOi
xHlOmJorqrl96ItN9gnM30/RSOggLeYtFAiBlMd8gwptyWpUR5lqYaYf6h80ZG8J
tPdFFI+0c1nvEU6njKy32HatwcTRTLk4lqo6YdsfOLTICsBs021w8n9EUiEkm3x3
v7guHWSDVc1fHUXtzc1+O2wnMJ0b7MQuXHEonRN3YQkW066yujauTXO/W7oKbbJs
dX0muLp1dNTYnJ1RmWm1yxpZC6cGh2WdevC+PI8ogXIxY333dqMm/0tD/Rj6p/t5
SZuTTa1QM4ChYyi2HYEn0Cwmqeytp20mQCy7RLEYg7r79nWEuzFCMJqlBAfQ5iP0
8rkM24qfpn/OvS+HSszQzu86eFDLR1l6P3S4lEECxIr1br8qRMknFOn6Qe+pgmaA
dbyXzN4uw29Om8kdlJy27+JiE/ng9XJ8ssuk6/esftsXmVyl/hHAbhvPRriZMk3v
nbxBeuNWvb8yVvA0CFqX4WEVt+qttfwzPClf2KAe0mrWcmWNOfIRflj4aI63wJdg
CG12d+JiSx10ML5XsIe3vAtad2zlSdOIHcqG3HeDx7LPvaeRLqWgEUIIP0r1x00G
HnEZB0GOhQaZvqieWdPTrQk0rxm7d75KEeaRGmCd00qQGVUdtfASWJsYE5050vuQ
koJPFZwNNzV+Spo9TQAL6UbtXYsnMy5I7V6+4NGl7vLLv6FAvuq6gufPHunlaQnM
RmOUKfg9h5vTlL/4lEYzQ7gUdxgWAeXPsP6N5ReyavQoi2LBtyelOaP9B0+yuC3n
X5ZaR/cUk45BjNrno6ndOrMspbgDu6gdduoX4BzlW/E5xvq58t4RwQ5NJoMalzT2
izio4gEA+x764NPJraUgLac2wJAWbqORIY3L0upFqP8LI3vGvS9AVB9OP1FtsdRb
lbbHJidTnfwvfEzoNUn0DBLyml3Q8svp59Jo2UEg1x6Z/oeTuC1K5nvEuGp7MsK9
w+bSJ6BE86XaxG0D42Zgy9o5bVQdHpxOJlyRc1b2h+bujgK4/g04zEs3Wt/qJ51F
Jg9ghWAH7UMvCjSo0kDqmirj6h5rNcce91mGx6/iiNVxWgaa7iDBbrgFXVnHi+SI
pSRhDLdEQ54mH87SmkviI4qrYMruJhniKaAtXXLAmA1TDBDhOcvas/3zmGzo/zi1
bi11qHy23hrHmtwcq0+1cRYzR4OojlupPNmyQZo7ZWQb/y9L1vGMvRNtlmzy+8GP
WTCiiqAChEhxV9XYQTivqxam822NNqM752WUI2RScaIUY5T+rek1bmSOqFTOacWh
zjDQaOFzlhOlqpyGTivrlxTOs2xg/xz+O5ThzVBL9MFGsp0eberW12YKefDIv2pk
czCBuBjv3xTD4hP1jV5CMqplh1zb3yr7G7Fbe7KJDEm2LBAztgfGV4cFdthoPxA2
ItD3/ocj4B5SkYOrXqCI2GvY3B1FZIa/bGMCh9ReXnMaIcIDadOovb6iXGVJpeUb
w7bBsdtOXW/sYayh5YmdIZq9tLch1Qx74jGoTebpeRPFy2pAmblzTjrK4IcZqgZT
cIIfRrxvlWyyb42cvSxUuDJ761c3yCuz9pWyXTn/z/Qs4Ib0t006fIwtKdjzT5nl
StF/F28CMdx5aklc6E3Y9AKaiWsLR3BnRzqxsOenxkMZNkO9SwBxo7+vrxEEewMD
RyOjzIerm5/MRl2YVP2808vJR8C4HbzBJNgFRBTrGQRE4Klwl1Fx+GhSR2Clh+tq
gKj7vv5fZa9UdgdjsrpKTDxszcasdAbodhdJmuBVhsufSD/KvflAFXZMWZA0qWXH
hXL5r0FZIIBnSfxUKiAbWZ+hkXRvEqpuHvG6RmHkk3J2AoWuWZdj4v6IGqSmWSjA
ZkTYtLTmmnGn9h8QgGz57IxmV0oDWl1wrx9mePFnkahWuis8qU/XlUq1ZJSfv3Db
/b2BTKVdJ4O/ivXRPPdudQ00Bd3WJW+YYJToXmTKk7+ThVodRcK6HguPBCD+HJfx
GXoDbCXYYNLK4RDSXtTYYIk1TZnK2ego6SFbCIFeJo/ExTsL5rgjnzkIkeqI9XKx
kiDv7wsqxID7Ql7EMtg3/5qp/s8J43aYXarBkmuI5Z1K2fp21nSRW3hUc55BygL3
a5Ns1zva0nmHnK2C34gDRE5aud/Rv6ZFd/ubzvyXRoH2sQJ8hgAdRUC3kUNMzi9X
KXmVXKnCN40lj4y/drSsSvX/22+9/8VG0hkQELTm9czsbRzwN4WJz7HxjN27ObZx
NN+TTEFGgCrfMBYp4boKxK8snvJjR9ka6D4ixEQR4KTxl3YTNL3aKPsDONYZXLjn
Z3/WdmiYdloNA0VuXtbypgcJZfm3941CVkOCf9pNhlbsYrc1rNXg6HklOKT6+VZ+
j/R4l+ugbXyUmjasIqiI4aWGHVrtxk7FLYj9+k5pFwn151npHLtIcn7TbgRTBFPm
dWggqazUHf1MZQlBjZYWK+1f0JjsSW3/+Vu/nYziuiMh2S5oJmaEWyJIYALUEC1Z
RWBH7MX7DXtLFjyi/bSTWP8NyxZXum6tmkptSzPHd1wVBPgmCc6SM1KShasD/fxk
KOrbFwQR9lfaGaO8OgNU/xtM+RRl7DNSNIl1TOGO47trfzcQz7ESHT7BkevWA4Kx
Q4PWtr3mxERaNj6tg1QmcTwBsQ0wzCHod45OsBHb6H7wKPlSh8OtnEarG8Hidn1m
XAy0HtKs6qgrqHSdVc5zcmwDjetMzHjpaU4PE7uETK/gUPvBWWFVCrC1Eh5uNDrL
Y36ahxK5WewmeAaXEoAh1LtOzmduPYfshje5QTPGoGvkdeyFIUNP4bbJNgsGVCcw
eJnGcpn02Yh4yEMiAqUK5JK2kmwWyokcsbvOGjJjdUFxUyPl1iDKPqADgbq3XVtK
k2fxcADtcYzioRvK4tDn6vtSfJtsHme1yeObA13QtIMH8ShXfiR0TrMUzS1D+bxd
nRtvXH4ymgXsAZWSLlpUzXnm1qmCnI7SLaNZeb4gYvyPamDhChWUo9DX/kKcVQ+T
VZRoo8Gx4dFOnf534Won47JhMCJTPzTPZfgOx8p7Uc+awdQFQKMBTgMkZAkIeLJj
AbTuFeuhi4QxL3YyaqrjD44Gj88UiTDejMJ+a07BVIXwKNwX2LuXfkUj6zb4+Byt
TYgfUt30IpoTpJZJ+2ywLZ6KoJAimO88UIxOS0yOR3+8Fb2Mhz7SktVHch/eaQ0S
z900ZE1y52T3uaxo2WdO/28EEZIyMMdKc77YTGj7SnYnw4OQWnTqTGBIqDtsi3ij
kTpLxfzOyjPtjyqpNVw6wZaC2rNO0KLNtugSbYvFooMTkqUAfUFZWRR8vKd7hqY9
0KlNiANhxzeU9MSe1o3j9Q3kpWMFAioyPVV5ef0dWcz/m4JKwqo++wRlLgXzUcFr
Q1uYrS8qxLfu92mZNdtcW7/HQ1Jmrp+PcsCgBlsorGO78HiEymf39pom3tOW6YRM
pWw4vK1rWGxJ0bKJmHiJSnvGjMQcZ6CwRWT4yTfLo5JhmyJRDZzSS7gWOTyrnG5p
5CxA8ZS1B8SIBQcNErRCwXSDepiZjE4TF2Aa/OimtOzkNagzjleR4WBKJKjNwxGJ
WZzQ2v9J/eqZB1fEeiyGuvlJkkIh4VidzTkck/LULmcfYOnE7VRnh8WlHDo6GfzH
fsNKTqeGvw3G2CYJCXU/HFGQCzrMHrIBVODTYD7ptdXxEdEy8O1cPBRqUFEOB1J1
D/LW0U306xLOAfJI6jDmrzERkqc84qXD4BKQI+KxeZfGKhy+08WZBiK3P5HwTEoS
CQjBCXRGzRXp/l+oIoyrg+omjiG9wYU4/2CwfoIrJPUZGil57YAIAyrcl/fdiKfA
FWv46BcVaqIFWUMcCWfOKVJMBVoQVLNuYifEh4eqRCPRKS//o+/GP5CrXOjCV2cH
Oxuf9YkkQk7Q0Nc4UbzaxHci/klwiPXQcclzsjUHc7A2rNrJXMxioudS0YORa7DX
YnLMSyn0kT6nOyDb14crEdfNF8AMSa/KoRgHfmLxiqwW29r9QLmhLaTa1mwWHvOa
ApT1wc+ThRnQEUWMu+FkDr2LAiqKhYwZyeMci+MTuEXW7huDQ1/L/XvPMmXI284k
o4HGWvwCygcMgQOiV9OGP4vUt8OVCCV3IHC5uvptu6jHaE7bXkFo1PMI9P5kQC+j
xEdpKCd/EkMfgqTpqJGTrFxlJN2XRP2kHOL3BVN3yUCT5mnCbjPYcf3J/mCg0fMI
A5IKpjF3CoRAk6cj3PsOLQ==
`protect end_protected