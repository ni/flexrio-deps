`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12064 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
DBGZtUPdvgnvgIFp6VMrQSZb0QgH/cWpY+LjT8YDInMnarETPTlIeQnA8CDQynJP
tYmCHaTZzDKuVaMowuYygl+Nwv0gMkubNO8QT+iWYiFPL/m4IRXD48SbopKnX9gr
NFvT3MJxWtA0XvxoiXpIYwFHpf0ILTEZOPfmlmBvMGXbjYV1kafA0CgWoNgwwFYK
eLirQdv85wMQSIryeeHSALG5UY/cBSxKvXNwqulIl1h+lSusEVj8hSNUsXvtePUN
RRqYIuVrMoDYXKJ+yl9paOFl/GGLP1i8TwRF3DNK1FxXikB3/GpRn55y6R0SpWzy
qmhFSGiovhO2bbmo30zo0CZCa0fpNScSEMm73LYLc0Yw7kyaVeaPGxHAAmYtXtwe
r3QxRJCV1JQoknNUpLKfxXW4vEr8ZVKJsJD4oGy72JEAcHPzy7PlABM7uz+iT+0k
uTNHLoW+tmQJypqPIo4pQKx3J4SzgGcWXTftHGNTQ6UpBUdLsqTJNf9rgvZVpv4f
RLvc4yUovsiB9i/zBn1MSIGuzAC2emGIAyALGEL4LX/lMJVulKQqY4BdVyj7jxZK
R4h0RGdc+S9KAonU5a5xWKDOT4EmCQ+/OZ9CkUrUHNJOK2rVGdGyOxoqtUp9UKp4
9yK7n9EcE8exS2udyJLI2QLNSear7NG7k98XIjXhOsmMcAyfgcDYTsha20ShKpKx
S6Q0LBlFl76mogj5cCYy0zy7ztvQ42ZBCV7O1HM8kXgBHUvztwEsLkLZPnEsc3lW
EY5PCwhpGfmv8/73X3uD80TGcKxyOpnoH/9EVv5jsyB3D97sjq0yF0W23iJ81fNV
+eMIy69Jf7KE0ZCKyHG0DGWP13G9C/Hw/kkImS0ufZIpxptEfz7U8dbIiGz92pH8
d8m9snVU9CzRA7Huto/XvqcrYxmosKlvou4aY9o0Br3pTgltYqErvkcIGgoJ1tsK
Z+jRpFE4O1e85QxUBUHXmH4kj6pOn6IdFblKEclyXTzb9tZtJ5fzafakX9EfLZ47
jdui0h6DLPjF6QMqKl6jZvwQbcec4mgUcVxQPU0+xrNQcrASGJYMyX43xlvSQtrv
zOF37hg/sfLIu4ZaITF77PymPFY/H4KzwmMIncbjixVsEopXbeRC/9nSBL/Fvlxj
LNWlFC+SQS2cf4WauzFoLWUPtZIGpWyy+Pv0JxAnHneZl8FQIk1B27rVzmD2+/nR
GtxO3rChRb5K3DhGFwHirVRFT5gw/yUsvfQwGKRFWlLYh9eGg/PhYusJ237Qx9fb
mWCnFznIh/2iLLVWSFBxiSgPPb81qRXkKgQjYi8zkF/+MPMake0bc61Fvjx22hPQ
AIfjO2vop33+yFDGJJZhIeNEwiUg39xc9XxyUu8Ko5Ci0Op+FBgK92/cp6mGYQIp
JdMAwlaXxNyn0a1xyy+k+4ChvCyXIFdRX4OD0eHkwVAOPxXEZ6fsVVL96DtGlvml
LUsKmxSiNRRN3rr1M95wjgIRFF3v5ptCUPJr1zQh0osW8CS9Lt2yz38hiFbzOpIQ
4pZuUm8CZ+HwyEgsOT5TWQPRFIC/qOtmz6sgFMykpMe4eQFeIF/8uJk3XCP2D8WB
A1yeZjmCasnxBdUgooPV8feNCkNpJPPF2bWKRAl9lPD7wktPCEI1ZXNFjBabJSoH
xvhZTn7KfG/U5AHOs4D4wyf3AchAF0T9EBaoYrh0P4V7dLNMMMntf77gczXoxPHy
cs6n8YBRHgLsxEwcxMLfNIyFGNurZypYtunmKItDhb8NWfYerOSSOIuYMDIGqh0X
vt3GichyXFFbOSKbQ/8bMPU1EliLinN0sMu/11efvbaxFujUXLJ4hkn5+6zSk9MH
LJO1YSd9zcB+2l3ToszPtkV2TjRnTTcji9m3GMmwtczZ2R9bDSbjE1d6Wii06aGz
iVOy9whr7PPNjqbcakkJKlhDZXeZVkW6Kh6YTgRAGtpkIUpqAFZguW2xrH6fwJ1s
hSd8d2I6/rxYvkvIQO5d2HNk2U6Ua4ppiWcUSzsp6TgothkrXgI6tnHSHX2VeCa3
cmDuqs6YOo1PeuxDYIZoguGLrOK/qP6X1TJ07tQvzDSSsgwbwJBb0YDY+SAH4s2c
QhFoejSXjeYUJ5xAFXq9nDo0/+S9VP812xqM6CzpIQJZiHgttQBuVafk4NEZNu0y
TANx4pirCK9jH9ly8hsIGAijiksdgidWM/R5dC1H9ilG22vPXEg7AAX48GFJ+zmy
fK/vcPzapUZk2goElGv/8+P1YqH4iGXEs2KyTnt99xlr2hx3yTM1uNpYBhVVhT+R
PF3w1Dd8E++S7btygvmWcg302YF3SQFrdC1pyqZEfetvOAe4N1IQ37z2quN7cxLs
v2teuiqbz9gHF8DZQRWq0jX/Js7gR3rQa19eY0AgUqobvU4XBdPMfQq2Mdh8jfTE
N8kNhFpCv6i3rrFxX9s+yHNpzWeG+yfeal7kyuUYlUsWskXQR+/6TmpjRa4nZIqE
HR9aoQOh7zOlNS3wMAP6kEr8/+bnDLNMqPUDlHiPzHmtkGkfxbbU9VLtchQX09VR
XO8UXyHYG/oElOvugvf7h0dmTX0HRleYSYR3+DsIEOP+jDBf3iYnKepxj3P6DXyf
Q/yKy7xtNEqoF3ohlK2oXC80Mj80i8hJttSrks8WzwF3OnA1dRbS9eBh8zMxsRjn
Gti42IqypqEk238FHmATplJ5nEOfV42gErEC7ofZokW0pzwsjBWisSF1hyzLVrHN
36+/KpRV7hS2J9cZaigaMiZYuOJlN2YOF936+52/8dGnyTeAoW4HLE12AiwgCFv2
pldNTb4Ytv1ATpZhQd2/tbTJYlbp1aW02PPCp6uT6RBv116ulcFxCzkZFPcvbKvD
io2VICrCCLQ+0WJNdQGvSEqrp5JV/6ZMwsTPxhGjcxEISmuAmuTh6SwhUWDb9wOM
ZSPPTbvpbgCaTdZHUHfJRGE6DRGP4bUJbb9hZ6RvjGngYJJwhtTxVT+EGYkGjK4G
iVclEtO0gFwiRzu+L5ZqgUglZw4dRHArHR4k1Bks902UyhKQxrcN+UDWtPxx+VQH
lBlqWpWio9YBzmq/LdPx4FEQDOsHmm3kK6yEAr9Vr99YNesvW/GWhKDIrUPWfdo3
E7wUdmurv/sJG4B7Aa2ZdbyhTxxsdMn9RJRzmWOSe4EjwttIlIcYaeAiuawEoKQD
eo4yaDO/zA/BamEc6HRpC8dVcpSL4xiMTJscjdvscjLV2eApcHRLIZJNuvG1BoVb
Y4lMqzlAuvvqor+s3wQtdwpdXfjbApSbt4nkc9kaNYYRAd17a+23pvPnPwjYKbym
YKtZrMv1fBQ4/LkZvApsRJtDNe6YaxpE8MMr7abwNSovRZMaoz/rQHfuzOZMX0Br
cnZ04kfigcfwJd+QE+BfaKHa0MuhWWChWrya0of+45/UyKD27cQepIuFtoRER9LL
hVZsl8xlzFLdSQb8q9I1hZ2hUjzqHxzg/YcbbPZHxZqv8Nk3nPQG9WZC5dKcZl1b
Mh2+jvGPTqbbuv7PZUdoK9uI7O8FvGn30LmuWGc+s9sHtxOoUQ/PiWiMIr58mKh0
XoW41wZ3lTTQRzuzdArYmsH5pgTJILfeVvzO38pjD1wwRIhBXV7HePu/kfctf0SP
bQXmRIg91+t8AeQ9L1uwjPHSoBdPESqh/ySHP5n8PtTxAsyZaahrMmg7VpzyAY88
QQD7bmML4CtwbJeTQ0pBM7huM8Sqv2EIC6PS5vxZNkwL+xEY7g3bSOPoL4hKyA/g
d9eU+fGXnEKL+fQg7EiWCm9nSfUWnyjfyIRQsV7kjbmBjsaKhPgpK7VgVIXLDfQv
4ma5m7tO8/11/wyQCCrRCohr8W8QXgOIktwn1E/xZEvoGHbxFkbXdbMdrWrRPP3v
GZBGMW6Vn5QlUZN0Q51II5e21JQPcz1TNlC+xGGIlspz/nJEzlNb4xwPcDXCIYWK
i49lkMMLOxuqlV5pPMEws1H0x1F/VbWjWIjQ4O1cXiHYngIniTYJ3hdkFE5YrO1k
RlHbJqeZBhn69fDQVqCmzTtre9BUzWt/tYEg33Zyxj8IOVY6FdR2Z5BOTDuiCBgw
GbiCqP39AFGkjdsej/MXdpcmSjflJ7MMdIr68a8+hCks6huhKJoBGn5GGzvY+tzZ
5f6DQQRG0J2n2OBJEjtzUHvLXgosCCkDl5y3BkWM0IfA1j5X/vASgWByt4/OC4Nq
fODkJRtEID/qWTIdF451Nqhn6YW5zju27M8akGrLtSAyrMuJoQV9EwbQr2a3V/xc
dEO7tU1bGnIQbbnIN+13NQR1qPFnQmx3dKFI0f/9B1dGFo/E/FEzvi7uafuVg8MA
rsH7ZmvsgTpdsDIFSXVUPCop6FNTiE9vjx5mmxf4k/swtaQVdDIu5Fzbs6qImJr9
3wd+LxXDUtZarFGekA8ushR6DKsZvjuCGc10bfsQFWX8bPWAo2pOIG16RvBWJomm
Kwui7X7hZo/OECNvkEGJV+CYpLeImHCRy9LdwW5yzigMrFDRVnVkC0cht1ZfCwY+
/cvya35Wj22TwPenjHweXftUensUEptDrbSucDAu0F/L7B9URWa/zsRNVEVWn5oO
VEYbTVX2J0RTDcVrEq7cMTWqiIlcaKkdc/3CLW6ck6AWxu7HYiwmcCVxtZ6bSm21
UPrxATf5/8Qvcr++smDBHRTladuxsdW68B1E4zEgApP59P1YkC/ZsknTYMMQEDBs
GqxmM3xLssmVMIeB8DmlKr7vmXmHza0ff19UicpddzhdmBYWx9R52iFRkvFiEEa2
uVzaem8MAX923xRpA3eZKtYj/cylSr4G/nXD3qjMuhAMMgzmD3gNLOuRGNHiFQJs
IKWdwZGpDfUehfINi2djB4QeuetcJUB5rLDvMojpN7LCOr/YcDPycb/5m0nAWWvv
RdVvgz0mMWeogbl0o3zx+yjfcEFMWPPlbAZ52CHT4jsNckL3WP05yK6yD3E7Lysm
hXwFW5MegKLVkiaRWy2kIwc4xcxfaqKznva+EjJEGkZzk4uujIGCaJuGRc2wf3JT
h+QtVn615JXMcRfYRqZ7/csRXTJmYoBla8hxZ5tkUBFE8sxnqQT6PFz5jSwbHhJz
l2BYJ7iNG4igga5lIvZ4qQ9eirF8PlAisK52ltLnn6Zb/H0KDAUlEGu7tnyRuwWh
yioAzfjBGJVbhPC3KW7lOgqPb8NPm4yysiEBHD8d7XCOOubi0NT6bXaY54YWlTVz
4J2kmejLiQ224A19MhSfnvwnRziGzROPg9T+ynopR+XTNw2B5zsi6K05TocpLeTZ
tCZmke9sPWW2Fu6Ro/ddCNMyIe84R92bRjNq/crvRnKHzSv8o4D/r5+FDShlTsOI
YBQmI+qQWZbkGUnkuDdQLGUB7tbGel+S1EcFLsDkIVgM081tkuNCQEi97VS94WmH
W4IjC6206zaOOHxp53ibpUpyVq63HuZmdCubS6rqdRjBIrlRaaUdmR8F0CTEkLAr
RG+zsSRpMzjpn5RLomgoVuFtl/YevkMUbBTX+FD3zKVEQBkOcd2SiGE+FCE/zuBm
aVvgSpfTu0uiXwSsrSXIfuDbiw2UzFgwuajXd1YZM73WwF/PTdQE9sDletYXi074
UeX1mk/FF4ySaoE7x05TkFtArTnkiV1AaQkSHJBf0HloZLx427LGCSP8s4d7ft+a
uoxo822qCJuxH7p9e9GXtJc1xlodx9mPWFaxHO4rhP4pw0C+ZhF26qCZhciBuPDf
JZcaogyib8+xKOKMDAIx2oRgvgNDQZ8CnKnpkqaEVfkNayHv2vaW0cavyg3IDH+7
krF/+V8xxaBU9mtpgPOwxgGs1F8mikQBPMNWtPhlX4IPah8e7l/Ck7oeV3tM/S3w
RuO1lkxmSXjE4JJyRpBaL8uUiGAPhiu1waArfe8mMi0B20ONj4J0Rd30iBeU9SPx
f4zGjOG6jCRMztAg4RZJiFmlRcbRnoHDEvkAlznQ7gkY2Io0DVP3fSMdapjDmqUS
iOz8+1vCBu1WAJ1+VlioFNAJF0Gb1JH4dgBwKifGzSPe0PthFEyQ+csBbsv3dl+A
Ovx9iCcKys+7b1rSnicrwKBvPaNoYEBssh6UyBt1cL1rHOS8zlW7AfqSIoT3zfWy
IKsbGugoOrYMgypSKocL3GsRvJndT6W59PYJYWccjUW8N/wn0Eo6xVdfW9xuv6ZY
Cfg3Y5vXeq1ya5gKeC0XVxd8XPRbrgipI12nwN1+4b9E+gawp3KQZQ3hLsSV0qkp
iYwHzVj0muCbF71Yly4a0oxw6YjR+G+OgJk6m4yIS9ailvHLv/8XLKcnsXrCEqqL
nq0bn4vxGRm4UYfrIHvYObeJZm1195wBnjC01EXUZYXjhiSUAUDuWnDheQ10Iowr
0aZBA7K8m6KxAUOODzpe7hZTy9HFjqNGvO49pHxduXho7Vjre1RnUk8HCQcZiQ/y
dQo5+Ag3EGC4hezDMXpsSpmsNGY7BmLoGb29oWg0fZa62qsbdp6qfB2m9C4kJLmX
B0ZCI24twj9T+77M6MEndUvhMHVqZxpp7+7e4mO3ix4vgMtuZpBccvzrD3vFWof0
tUEsv8Id54Ar/jTqHhIEfhj1AO7woA4DFbEftDZ5qlS7pdOHcbILVZNSiUwWM2cK
0Bzn8h62LNShY+TtXUd8XYvVgfmbUdKtObYsSSI+/qUpRWIFZ6ZOQUWia71ITsUv
UDzAsPNwKA9QDTACBkgaRyT96R075WvUvhYnSqOC2nj4qc4lLbMJ5uHHL4X2tBAK
OWGSv1FE15J3/agV+aWgzYIvdinguwH3c25XZmH0RQGzXXmHKMebQxWzE8JS6wJt
45zjvr1yQ5X7skoVXS8+3iR9kqmt1uYRLMptjd61UTIPUpnS58UB4ZKnB+COR+TM
7nn7B9vwBkgO5N20+BGQbWHTytdd+wodQMGyNbYS++Ld697quKb+iL0XJsz+q3vS
s7UmTjX5D/tbcOlbmjJSMs93Taf0xyIgVLpgfcWbJmFtJykIZHIt2dCZIBONbdLA
SucSGz6bimmmW+yZDAOpEOegviMsP+D8C18D8jntT0ZpMSXqCPhF3pHqjjUK9uiR
pFXUIjN64ElAoGI9/naY7lYSEBDR9b39MQp5VP6f2ep8VBEqtTjustyAUWzWZAEJ
vaKYZETdl3oeDoA22hU59YLbwZPe5BGbPmoUTs95H/Q/4hB6PfJC0wQhTzLubPO3
KdjXgqjYL1OMfGswmv4zN5F2IJfwrHeuqXl4ZoWOf2EqNx3HxmXPXArCyJBajrOu
yXvslvJD4F4iZAO8N20BpXpOKylEutdQZQdcJ26vc0VMyhF5LshbuKUGY3Y0bipZ
SBIwSBS1EmV9FlRtqQxnmGm4yxTRYw2ozcGLhL5D8F/OTmA+p+Of5I1tcDsUEvWJ
LhOpPL/5ZQ9LXOXYfaIkc/+niwdIHLt1hak9EjPAQZTNDNXEjxAuYitSubyvN9rH
U8AL1ZCi+5+LADfmvASfw/vZ0eoacOimuFixjr2rGp2d2GmfM9vcJh8DZ/y2c3Qp
sq/8JqTldCTtUsfbSl+TicQvq2k+CozN0wzoTFM5U4k2vMyBqpWOzyaQ2cqNdceh
XSO8JzBlVuo4NAlXfzzxYbo9soQBzNwkrVgikRkaGOCSB0cSufzleo+2bC9qGZb9
4KoB8aNIl9Jzqk8trZEp7UfU2QWFPfwCrkiB4pr0ey2rhMpuLj0CmL9g8X0H4Olz
P8CokSs5dYL2NB3IL5MH5K3u9Phh51lFTEP/ZI5xMwH/3UwHgNUrmTpxaDcCRYwR
qRkpUwWn8B7nF2zDEczmVqhOkaPRc4s44XeEcJhV4z/ATx8RP8ob4DD6gNII5EJj
KeWqETVzit4myEGD3XXH/Vtl1QaTpjCCbwhj01lwdFCcd2+suQT2kh8sxxYthCcb
Z2YKie7g6ZaTH6iXee2g+wk684qC+PnJSUFwLZThIG+qzKbof/BY5H73028rE17j
WIpm4P7TVwaWLEAs58MHDTqd5rmEfVjNU8y2zetOxnDez5EVT4AdgMvJWY2bTyGa
UU5efAczn1TkUF6Dz0ItFO9Lra3DRx+yEirkpeTx877Qgo2yz87qR5jBT8Y43a+E
WBzqP7EtmZKzXMhZWxNDVH7ucalIeB0wEiJgZiSgQ2/rj0JCn0Kr+LX/+X3KNGP5
DUCjmCOQG5yTgyKU8tvrbS/DBfHYbsn33DpDr7fl6mtymO8e8/nbG2JQIYzJncc4
VoESVknsTh1odPUL6LZ2kSJXJqTV/FKXNW5ZAEbwcQrv6LezOBkgT6pih736N46h
HQLcZNPwz894H+7StXLfUmx9xp798oslqfmgNMcOftWEkpYGsNjzz4SaMHgXtY/b
ErEzlyyz882mP5lCGLcO78w4t25KvWFF4Yrx2dx7RFiAFUWxjoHuJ+tj6vxyoFIW
5WKQ9fhhOhMu+HXok3xQrKRuJ/US0ZLCnYMEpN3Nxdk6w4nrZpi2uQazEgW1Gntk
202bKEJhdsicf7AKDld908QgOC7R6T1G7+RMs3fIUfAG9r/0vZ5kkAVRUb7iR3XK
bv1csHpWffTEKbHWHVJBmaZTv7MQY3YnPSeIcxq3GXNG2MZWyAk9NQxvzXVQvDey
Q17x+AbSRN7o5VTtetT0tJgnpTwRuAaufc+vI/3wUh4yJmxCt69x1hpnRl3FHf2P
lQPK7b4AO/Nnl5eCTcohARep0g8QZqgTk0lXsgvu5syfevnz24KrApsi2y0ZIfBT
lyCGhZFCYvXONdeobsFCRV7K+WlW2m/SuJsaRbGmQolo7x6oEa38kbMuawNRHUpF
P+qzYfuXG5j4g0tFenl7E9IsQqoqPK51vRavZqER9QEKe+3gjtxEzbN5wv6fpD1D
c9pEd+G5FZ8j2Hwj7HYp18vKuig8YoMR9XJAs5w6Z6tJ8ArFAWUYXVQcI0jw0PnV
/yC8eXRf2k2y0Eha4BgvDrk4Q+zikGh5gjgLHlJiv2crZcnW68bc0M+2rwPoAIdb
ef1vntkwrGZl/cftXfQ7dRN6eujiRbc+Se2W+MDo+ypa4yj7Y8tNQyeTlrX/+HO9
mevmvBReg8AZb5QVqrVJ5vzPqtMttWfCSuwZwq5A7PYEAO7iMWOdO7RL5MvCKW5d
+bxAJeg/ykOPUaupRFeTse2lnl6P9fiAEMStTexYW/n7GgBQUYsRS8mX1kgvGRF5
SnHZf1p1g5eslA/L4LzzXWFwyfJOG3M+K+du6O7Z71Y3o2rm2sIn4eGqFhXy3FTK
G6CFsmOnJHjy6DC79N/Dwqo9/xtx4SXgUtY9iB15j1O32iwuFLw8Jgom6F156eTn
sXUL9wtZbNp9tv4mgTOUaOtGeMhsCzqUn3T3GB2odxlckEEnw18lH5x9FayPtO2y
5DOl06wUSruKNAmGH67lm7jmYuSz7mOgsgvnCo7McjNkuw+dMnqlX1DWI0JFyWVw
8AOMoCCWnaG4NiKNpf579c5tFkcCM8LR7AGR1gL26YFDPDiaSNHpIwp81tmGh1+S
a5n7ZIAMrvoEGghLHaDULbL1mxH2vIFR5TpL4bOyyLu/ngkBkJ6zR9HDbKaNcIIY
9i7j8FqhrmRsCCEYJBbFeu8uKh1rrQHEE/Sg6B6rbQuV0P4ShwRkKwkwENv3p5Ti
xVmCa6NjVPBJeG52JEs6ImKaFOEyv5hiEOAobCWyl3GSn12a4pRC9kRqUd5iyvhs
W2Ak2td8iSEjaDW++G77JRqBe8O6H9RwL466sPY9pyHLkA+V47+24zIBMA901h5j
orIzISMl3Y9w5SLRdYzYOMFIG9wBXjhGAk/iv3CDEnO9kelhQplgjSCbnMhnHv5v
DZnqNLP+5Dx+Z91QE6c5z/auMT7mYqEZRTvf+x+EvB+RS6fPZ3ox6U45cJC0syZm
KZpym7GpWYcWGR5rorA9UKIR/GeAGmOgQZaQwv5yZp8SbtWQcVEwNXGiSxzdJRST
2rBgtgbsxs4U87Zvx3//5J58nz6YU82Ipn2eaNmJeD02w6s3zzMSrVTwpzZpGhpf
9v9jG/kiY+6AIcJ1WL+zgyhF6QRcgny+zaaoxZeSF8UBkST71HRiicD6RoJb59fQ
DflRT6JSv9wzEJElc0NwCp+0Jrise7zfO10qZjUIl1GbAt4dwNDgjHzDbLzG1wrL
NivWOC2QB0TeoIaSi9quKVA8AAzU5rijKD80chsgsm26+HrMZWslDCwwyyEgDkNh
hz0K+Jw9D+m5Ui/3PAQzzz4yVScgrKWHRzjlHjp5RZERs3VZfMC1rhOtLkgmT4Qp
Aqz2539tJ2jOgwvua+9ktHWyfSZicopmpB0TRc3TORfGC1rXLdlksTGdBY4AjmRE
E1q+X3LVckBJfrjkCjIWHNQlhcdKfJGhXPfTYIcdFMjdKZ+PsHVAS82Xb7wKRtpl
iCSFjPG4SiZorSa+uOq+ZESbapsoO1OK+WIO9e07T/6Q3ZpTBDLy0RwVNsG2tYfZ
qkq/wwx7NgSbRdUpsPezqc9QHVZdNhgX6Fz0d/DPFGUZsZOBknThApzVYh2uo82m
3LXO9fCrKGnb8H0bcy1Ahaz7HlahJJM3AgfreM/n6WQBA/gc7V9DYh2d6ehAafYa
BtRP23RjRNUk7Sqjyhw1G0hzD9YK0Jn1wbUzx+rh4FyvSqrYgCSZVU4Wk6q1pb/q
HKX4nY+eW2jmhI3PrAyPw7SlYxJEa4O6yEOSJ3XIgtpaiE9bQC/YlkXWqnpri7zX
CnXeug7YVVAWxeQIewtZN+2rR9YNkq0NWTBHBT2EoZsuBPwBGUsvFzBmGULN/VAL
p7kNs/wSG8F8smOXOcovjyJGRKgWK9K5AYOonKJKSNW6FExq+iyF8Vrnt1pJdVLU
1tWIqiIpU8Ib46XNxFkUbswNSbYKHg41+Ml94tT4fh5vplDAOG7cymZMzENkKSYg
sMbhcA8vU8O9lxmhlwytYaGYJ7TCxauDDV/vF3joryb/KY3C71l9WHRXxeHZPeVH
RbQ0Ry9y+WC7nxaxhAsjr/4BMVIEStkkqIIwIr4HO90bY/4/kwNJ+MVOVF8GcYQP
EsEDqGnG4k4JQV5a0CmbuFcMZB6lAm1+gasQxs5Q90XxH0ELLHfD73JOSt3h42fM
8dc1X84k1B+uJxM1MW7Xk9S1s7I7HbQwwcKiVITNaIqzZVa1Xzz+yl9MdYcgoKI+
H/h8k6CKoLPQPiYaabpMMXOvuUcMsXCvWUzLoXw/e1OfSUKvJsXCGLdZEaTNaT+S
JPzca7UrE108Ldg3ZIrrqArrqUEJTSrxQOpjABIC4q7AUiVDxIq3cUxiqDEq6tkg
g14YYf0WpUcv9f15pb/6fDOHJX5Ad6Q4lhZkSudyL2qHTzAo0OZWuQh4G+Kre+rz
bwl/vtxy7FxYm0mdkXDObVch77dV88ceWoYUJXVW7mlWN0HCRU/6U/Yul3CWkDF/
SJIY5/AZwektIkShVnciU3OdSVxSuoPx0QWB7xwiedYMlKhvTM4sF3v8im/z9eJD
+piUti4bJko47pdm8739HUXX/oIKQ60GQ/OWCko045+jjD9yPtMk9qNDHuhPcDIf
hnlnbxyc/dcVsjZsAEt+sc0d2xZgUq01/zRWcttwIhiAOrhuhI/IwXUuEIQphiM6
mES7W2rYxjFX7aJ1Rew1/OWzidRLprTDt42StQtrZ7SotcHaQp3vsWP0aydno/pY
7iEt6BaL3Sm5FOudu04Bu0fG/2CEu4pRm7ypKg0LFSTAIlIfbbS0AJJiTpEa7mgV
UsOomPP3t4AnvxM6PpXwBG8AlriwgmxQrz9NnYyq31vMBbuQQ5zgL/vsd+qFJOMp
1kO4DeOis8zKvXYahlmxfr+DPxKXuGp585Y6HR68TdUu79TPcptmEl1vA4H1QiMC
UAt4d4gkLnzNj9nyZycrKhe40BuqV6II1gwXirQgL1j/CMEwCMg0lnxIseokYcE4
IUn2zx2/nVJiTssjlrckdSel3PpAv1tcZMWXRjT2dpGuQqcowWl0yjDbIdqKQKCq
Zgz6VwAOgbRFWVIZtrxXDjiZYfAX9OS4+Im1s3GgcDZsrb/F39C03xm2rBkexfyS
+ktkp2QQk1lb280QZdexPDKi6pvSPlE2YjkJjRy2mc2XOffp/Yxmio2oTLQh7XZE
Q4Zjwzuud9JigW0PifXmXvWmHQ/sAYhgSxz4CyqcmDjfM66jg0W/sMewGNqSgsi8
Zb1evgDT2Fp2m23QkBSpR7qfSu+X+ZFTjHDUXDfYFR2v4PtMh61BnagaG1UIWwkC
Xg3YbfRR1/+z7nBlfT2+1jUVH8ALbjOjnsE0tUyNiXZYNO+rf/NtzOfFiK6Eh2ak
Hy8M4DKikrHE9wl/UZVKXW6K6Emz6wecG58kLn0zwbYjFKqKdyPn/qUH8eep6R85
Xlsb0OYuuzWjKkVTnqBivZy8nJOENCZ3A4C5oE04xc4tiYBPt646Jjp8hV1Bj+Kv
+uansDmE/C25gR0hCywQJTMvjWLjkS1stALaDK4wBT9FHBne5YevexcYs8ra5vq3
h8eXc6zWFnJtPjzQ8GOmBwcJh2mOBtb3X3ldM1JIUB8ZcoDntlOsMyLsRkNqa9gs
9HdM201TLNOjf/vRZVNXHXZXJLtQ78Lhh6wP6KY+ef4RJOZb59GB8j8E0t+pUn7U
JoF1HYNReYOfmyWsYWRDTwpV1/ZAeiaQSYg2TbxBL9o2keGXdntRMonxAE0ckll1
6iJtZoq4NS4lgYH4y/zjdeN0zN1g/hePEMEa3fts0WWpq3XZZrAxheMcy2DbsZTr
+oz0KZQtDad5fQ+WPW6QsCLmyuk+dMRf1AkR8clOzJgfLT9aGWI4jSSpJkzGC3yo
sFvdbzwY1qVWS5GylRrKkF8eo2S8saNTIYWo0v0ptHtEAvXUR8dJAMQpT6dDxmXh
p5kR6JFT+Ovz6ifAYidV6iK8EVazJVpiyYLt1NjSt9HVt/s9xr/iitmMpROfi6Qm
MBQC/JzdolW/ck98GF7UsCNJgSQC0PlKFToaTQngHOvTCVdX/mth/mV+coe1FPg7
J82j6BHl+ERhRx+TIL/93L6v6GtNqcj3Yy57qHnBI5a4bcUO9+u0cTXfxBwljnCC
cy0vpN+jswvt6FxZJd9J21Te3mlkOm5V5JctdYXISBIzzeN+m+Nk/XoLfptYUiVx
Qnnf+1gH4/dS2PgtTH/N3KtN7FX3A4uSzw8CSXM+poM6W0JsRPUK+uYBuvstgQF0
oZ1/L4Wc9Gm8KFOjwDMJy8kg1iZLwHaAKJUsXifLUZWmgd7f798V3pnPOqFjPSrO
hhbbb2s/XcY7zcB9+3/s5CHisff3j1ZShvYCY9WdYzJQYwh2qPDQ9ufEq0jkQCPa
ceuHmc1thSoZCZoUnEmZ9CMmfaXCgFGFg9cL7/st9vngZUunG1a6wMlHhJjwLkDr
huEsrGC+b034a8pDSSzzp2hoNVLjyqJ105C7X3buIjdVDam1KZ6nL2QCl/BiBAxX
b3bFJ3SWzSe9yNYDnIkRcqLYZprXSQ4i8X61jr8HekBdOdhSYbg97LKEF9H2sGC3
ila43Zqv/yw0kA54LpBn7/3xchBB02Uw4i+JSpXToWNSMCKSYFkg/fGaG+QzPbl3
eSm6xIUHLrT0wVlXJq+CGIVS+0Duwfta6WBa4W1ZWKM+xx3PDTnQH1JOHuF0Jq43
/Re4cYVylB53GiJbh1mLDS/GWj37lI8M91lfOZNad6bWGevhJIWHj/PkVnukgChf
TBrJ0ix2FWeEvgdPP3V0EJ4kntz4lnOulcUqeKU6MWw4LKyaWYPr1zbMnQjOE5O/
+29Z50VA1vrGLhyOhXLol1h6MBvKK4LrC8ymTg6Qegr+Em4ZlCJ+k4uozwUtCb4c
eqFhcnD4xPOTWvCfN2TrYfsmlAgVCzd7PgHJOfxJjvsW1u9fCd9GpOLQ0zG0b+Fr
CBLqwwiXAR/nRTyrvuKMzdbPQ3ecteYrZ+Jct3RimCRoj2krjVf63P9eoWWSNwvr
ru7luGH/7fSeEKg19DJNSe9tSklkTMWD794HYOBqvsVQYH9LNTs3wi7wlPdc1gTA
vTrsx1+GYTsN8ods0Ev7wDm9ztwQaesbBkRcrd0mO5MP4Y9xj8y2dXMRDkPbMHri
0h3lq++RuiBJObETofHnQk6h2jmjFOfmGxpK9a7fLl90Kuh/eLDR+rL8q+nSv6hn
yPlMiMf4pvbiEgOgNdKyeYPvNmCtfnARNnH/dfnaAEBLxu4lHYrqTmOvMiYZ4nJJ
lfhJMSsZawaaeaxVVqS/v6FpFXYIDykixh3SCk6DG8OzsCA+Ne1nSvh06SKdAeXw
zhx09zlFOBUIvvEso9fDN1AXgxrdLwO4YAvq0is0quEvw+VgVIFHGoFKH/5BDq7j
7aBUrrUaJ2QILdb/qT3DUeFl8O5Q54KQCRAdVXiMoj4Aa3Pwu74SdGyWB+O6q6jH
zMYHS/8Qek/RIwTC1RZLUYUMoOeFWaYLBUGNYiBQqDixGCbLNlthyoy9iLlwJtzZ
OqdSMx3it/b+ICcPI1/GQigGHnNlPTdf+g2EzsDJ8FYBJjRWySY9RzmhgJ4oc40z
XcWIkbDrXrHTKLEkABtyI1ToSkL7gVyVi21UMja9pGPrjWLwRd97O72rXFrx5AUE
ki8CozBo+kjKFR2q+JSgNwhWDqIgibpnSv1tS9G8yKvQ5BYCLNT77yBN7aBHAZGs
pM20GY5bPqBQIGY1LB8ZlumET06e++WpuYc/+ZgNQzrfpl6eCXavJ1qNbHQJec7c
RdxcBCThoDlIW90uSxhLwf22HBqP4uLtKh/6/xjhLu6GdgMpIQxEdJCKWhuB8ez6
fwjdhsvMk1a+j4KUPMo8P7luvlSgTQDi0AbbZJ6kJpBiPqIaXLF5eMINIcMIfM2U
EcqLm5bgXBxatvEn2yVrKVHbmYItLScgQ5VXgdLxsFmakl5VY4ak+MNMqQb+gx5W
Jecn8pIRb5yG+virK5MUb4U4PvumzK+NkPgtK9mT+cCiWC9hB/iyjd13FWRcoACl
5SxvR/iowNhL3SEOhtJVkCCaEDlDYeNtC7fiYhBo/GA1HlVCSyZ+vSyxalQfqv7l
rpYNc2Eq9XUVijCr4DNbHtiFgAl9onFCYH3FKIy1nd7o3L8WuxcnMJz+GTLbxWVZ
cjcYFilq05DceNAr6O6+17W32feT//LHnrsOPhwYcoW641s1TrdkLnC/py/fsD6i
BZ78gX840HfiAKdgxKcZgr3EuANzhR41veCIsl//HS58UD2OZDPrEnFNaDyx9dBy
9q0lczkJkWPzJaZqACzC8znjUqxG8T9alOaM9nOyclkuo4XQdux8iWLkExDNqR2F
iKDm90pcAoEfXEEBVTQv9ISBOASBfxLyzz0P2WGsgV30jUTwL7ZFBEAHUOnBnkRj
yNeyd0Q1/6vyHXcxkUV0H6kBqPwG5IFLqGJ6sKa6ir8fbLPr8FVcv4UslB+CVK5O
cylRiiOM95EE1HjGF5n4qRHByqWCpwrP0i9XqO2ZfF7f9lQGcpgcAUCQC/Dl9S43
FVQs7gUVodTz0e4tBjlNurU8xnJcDHMyeH/oKzfkHPJJyqJx4VhG33LSKjJyD4cu
OYqxZbiGBl3EaOOIUj8sEfn345mX0eAAcYuYFL0KqKYF9tXfkCy6LgRujgrAxk0u
f3R+Zgba74UFuxa6PpSOW+gVuXqL/ElI3kAjifVy8XubHwnHrMRbmXNS2QaPGhzY
SbnKtjNXP+5a6pIByPUmIGnpreviLy5YqoZIgxnsOUL7RosJ2FDeuTRpvtXh4Kwp
rglXtJ17Ask8L0rgpbq8bLPq8O0SZlZC/3h9QInq2q+XUI3XF5npxfKYTih9ZsSm
VxqaCBl3gcPehIgRPWaZe8AO508HwfMoL0jUrceAmixWvfKy6sMw6vU+9KUok2g2
y7t21ddlQYEDzEz+DNYXbg==
`protect end_protected