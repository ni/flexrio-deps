`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15696 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
j8CKRAvULn7NFOL9h8Ek2jHLzoCpEgRSwRgxdOGQjWNkKl8Sj3Om4QOMwRjgOH7t
91sEuzZsuTb5kS3wajX0TVIHmakZ3lYqCRRAQXjKR2j9Yr548nbLu+ZGFvy0jBEa
op64wIb5lvjX1rxDr8knEyjkN6h9Wou8thApRbB4To8IqMvqCNaZGTKaz+jagwYd
Oak+ojn7doHqQ4gVuatHNjbAVmI3Bo6/05J+fIzi5EvN/fZyi/BVPQ+0Lyj3weKa
j2Xhy+qjQ0uOOC2EypM0Bo5sk6m06pYVN992q98YAZ2sdNaqbXAQMTaQETpppTYJ
wGW8a+W4mFa6a4az9Iy0U9ycQW3xHe3rzuSg+ooTyS/VGXJ5/TlR+P5ad88+wBzN
+AsFYWt/nxyBSXbzMvvJrPew6u6WwUtKM4myBqcWbtlVLtV0nGteoNqUE6Bu367/
QHQ6T0esCTKgBOyrzxtkOad2kfRS+MTJzRSRTT0hPT5oy2NbLpe87B4gup2gebJZ
qK5ICEcm07KZxq2NNqhtN0GDrFYr0a57q5idclkCw45zF4RpMkrpYi3+UOF3M6G2
90U/044O+U5SRUZAOhg+d5V3eVhPDsNSMnfFXqoI9SNd3WG0qUGw8KKNlWewqKXS
C7XM5A2PkJK1ryqYKssa+JYcD6Q6v1CFH6J55baQR0d9W3LBHd0pnvbwW1yhhhyL
AQt1eMPIMneym2ZyQ2GHeVN/XM7KvBUiETSFBTzmRstF4JVxqsPMqY4CoidsUVVE
YfAU1RXabeyb+N0qro95wIyYAWFjYX4luAFbYH68PWzy6Gi+ERRc3/eQXFi25TH0
BrCNbDWr+mjufDllJkYbK8W8ORnYkzI0UzZP332kh8zKiygu7cqQ0Gu2YCccFBzQ
QTF8rBdZBZgRDfOydrRYdq40aMB2MZzpu9XsgyL3QNDo67gDp74/GQvzCJUutVvz
xjQ2gszlgDur8csoDYvlZAW5poWccfEMTW0fMFvzS4louxtq94NJsQM4ALtOWota
Dv7FdI2x5aUxUK0jb4rz9QyOSDTqrmK4CaUyBWcCPMIsOWcjQlJlVpnIimqNE1DF
ugGjicAVIL1Wzo6fI4sj+ALqm/GFdqfxxRl6HCU/rbyYFeeH910fXE1sloLu3kaO
Y1TUkG4urORX+4Ypg8mj4gnG0Kn9gnNXGX+XFqamCzLxtf8neVvPaJN/aIcNmHaB
ZDQCwXGk7heKNVRueN0dyjaVgXcGvsAXKOxLifbcQBW8sYz5MWD1zvf3Jonu9D4U
pD/BZSG9lCQn2K9OSBWWHToYx54RB1urErIFFYr3ceHpv3lRnoJLtUJvTSqUJe5C
PC7AH8ZKJlvDw6lxX0jlaJ+/wdQNw/wIYaiUZ334fT2Y0RpgaM3YkIdAKEtJVpIs
VPI1LJ1BBtueRG6idQTRr70CyuxWiik+6y8mAsCv1aV9Vi/1wJ45GSlv9E/S3j66
SLsqmYdhUCWoghmyrJVp4zZfoZDHSw2crw+4HqlqMxUquMRj591GdUCjk+HTFLBQ
krDPlLdk9ozXRQs/7e5JxufDgBJnHeeM45J8VTyy0JUef0TQyVrG2YRC6MxFlHqd
jI86qUdQEvAxmLYs6bOyYhQU5qVbHjnx7H0co5i8rTqDKWJoOR6Xu6zxJxcSaEMK
oI2etotkz/wRKsjzAGaV50DPoKfb4jG6/nhYbTdHdPKiRrrcVD1yhZWYba3e3weh
CZXDRAhlztFxu6TUejs8uJKGFxiYs+9Nkns4vmhQ08KquNEGKg867x7qhDMopovX
BvxxH10YqEItWBLzp9Yaii60bEfOvqHLY5WHx7aNf0DQig3qUVkWkBuzUKSSHowt
vLalRnmvm3yEkS6e2XskwmDCFoC8yjND8/tqhnNQu7DgdDoU+92jwGSjH1tf3wyX
xGHvqy4448GYJ8nSzWBCh0hBQ0tCm1oY5Di4JiJTlX20YxLbJYNw7+SczkrR6eby
cIzTl2AilVcUsGTpkbWIpM4HdZM7UC0TBiEt4vtYcNPGls1KnE4rSloDKPmE49Nx
adwDdJdQ/n3s4rQhMcDYFH30DZYN2DdbLW3+aWuf6XWCqTwLtez9ykJGMWzOfwZA
7oee/40MR6kFc+T0/EZpnhq6LhVLe1bJYbvKNsf0RO128ZgIwbS9pPuvxic6lm9H
pcDi18kyHZBpY0iczLcMEVcQ7hDvRSQq9uMd9/bkCTZ4jszD3E+yUKvY8CeExVGM
HoMSZ9/p0BRSKSQPuTH1xrYTeRMOZX8oa8mEwAtJ9FcwFazM98EgGyhJkjqt+XIb
KiYsAbK2xxGYSmc1mBYoPvq+mq3NKR+hwQO8HgZK6BkLuHJXNYWlWFK0kF3P6nqj
bXN0eokfLoWlhxgcKzhh37LFOjv8k6oHFsPzcgrvUIa1/pJhfF44veRdI5C3k+Rw
nMi4QjcIiot/IyDqb+Leyxv0TGKgIfyVm9sXKYnzgfXoWmuADW4y005a9JzVkRo3
jD0NcF680PJ0+5H4c+SpNqMZ4IKA8yHPhlzyYlzrxY+WZwjF4DjrTW0YPk6sypQy
qpUXMe+k4qQf4Y/e35eW+7o5Ssw1DFzSIsj4Cl0f6TE+L1Fgnh2bD1D1O5nc/ALr
p0Z7tkD37ecHpD/hB3xw2M2v3mAJeQ+u2vi28FboQe4sBEcKWVDxDJh7KjpOaezI
cz3sU6ox6s5XlhvupnH+0uO059DXqN7lr+R+kY7yTHZyEojUIMXYSnVdb9driGHc
PonxFT3Lel5jV8/yFZLiPB5rCL5ic1Gc1okynW9HrlH9gJDkuRSzm+sDulqLpzrl
5JiQB+QU69IuFfasN8KNCzEazggY4b4DisghL4AUzYJKeMhy4YKYhnAWsvvIayD1
6kGtfr6Mlshg9/UkYfHEZZnFuTp8umKJnKgqIkGh2Ju13eUmm3wCT59ydAjfjBQH
dLzJd6NPCU58Joy3fOK+e0S2QjTMWE8SHOqaH1yU97fQaqHHjgMEKraInXocd7d3
RzgOHaF2PukMQsYofibSQlWyhK6xmJGHYNMFp92ku4zkUIXLyqwTNS2SD2+j0vJY
ZX/q1zaAVBqhWnXLV1fZ0zjIglmAVT22SybH0Idxocaztd3CAny9FKxZZESE0dK9
4FquYNz+2j/PjZ2f02Hs4jhxD1lcGDplENPNwTNGAXNhTUbzb473/SaGuUlM4SKg
zCGOT7VKpP07tAt0peWoT/XZlomgrpniHga8lwMcJ/i30yRjve0nxXwgqFGYNgNC
AiTFS0YAEFPSSSA9MXk6nl8V+hMiQ79Zm4IJeq+CZzrHqI3DJI8HHar8Lt02LkRk
x+I8yBX78cZK8bRM0qAPrsJhHkR/kdC39hxNssGYDrrPhKkyYM7WKeEp3Ar6p7Gi
BRk6C2asW3DAfIEs4uAfoc7HFApOs2VPiLO4GtwxXNERo+wzPKzZBjbRzHl86rXz
eaen7sec0uNpLpVla2ozm6Pp+L7CkCgjGQ6jytwcjt2o/8lFXYyG6leJw/52+p93
EIGWlg8JBNIGBdtsWQ66awPVtRD9lm1USDKe1ddg0Cn0WTTGkDk2ZepSZIMDrYc4
pIlCTWerDKiwLnuMcV3qTsReAAYHupaomgZa0celbPGULRtgRCk9zjhLC+oFXOsB
v3CgT/AuQoZOvJRhfQtw+9BKoGgeflt0DIhVuGpd8tD04S7P9f5uMmhR+2cOsVg+
3VJs4iWmyCqHzLy/U6DM7e3CMTOCegdM7N9xgagyfpe6kYSJZ3CX7Z2RAuYjp8gj
lI9EhMSDePKXwQS4jMOij28HbE1YnhaqkrcQv/qnC1YaYIJMp+Gi5/RKMT+g4fDa
ymusE+ZnMw28WwqkR+pJ8CVtj0RtET5xsxNvdLhi64o3IMnrZsRuJ0EVN9RGur4X
gpKLo8JhevHdbiunQ0XfBj6lT3g1Mm9GoPY2DCCNf3ASHweeSQRs582n2PEJoHUn
JOtBAn6hiytlUb2GKJ/YbqO9r5IJlYFZwAU0DR/1b7nHF+pTdzbCntCWE35jPt+o
CET9Ag6O+w9nGtb2kv959FcANfazWSsQvEkxpwKMcQyykjGf50DMNH1kiXuT01hU
AVl7NOTKrZQzZG0+z/uCNNIqGiG0vYeqI4YwdfwQGFjZUFnytUft7ilKmVNKaIVa
k7i8w3s0D38hevVqL4PE+Q03f1r7ii5gJXJGUY+oTMYuZ7+ZD5hs9aV5VYEPYinp
H9sVcarghkO/slPfQW697IgHbzC0lxKB6Xc3WUZw6voemQy/Dlpcil+X5QozZOMg
sZH2N591xKQCF6S/p8aLFrCBYdBpDvQ0Re0Sho57mqB75BoKW8ctbHniR0H1F0Z9
XNoxqpH1xD8g9tLCgWumt+LLz+Xqb7vXvdw5MnKSdtJl3H23NrwRA7GWLTCknhDd
yb+SeLdk8KJXenlX6n8otNGKJD7hu6m180dAgakZg8k0smxiLC52FwortY/fWUV7
o3arGcYuvTJ4UlPRLXT8xPhi/mvXx4HqdTYxvGyQf2Xudpt4PRLmMN+gnMqavsVR
15DwJINVSFjXqi1hNn0UiNTRudpZqxM+wqQeKTjU8X2tsU6h03QQLIHON+Yfz/lK
bD1f5F5j7UmborypgIVbM71sccI9d7L+Rb1oh1AQXq26QJchyln8RSuXuunHDd2W
Qu0V+1LczUYX+Y3jjiLI9t+aBkB7yBHPXxc0Cg20+LeLLsif0S7CkFkWoZ++0j/Q
32xlJ64twDqFGcm1TNX9emq6KiY1uK9OfXCEOOaTsyIgmk6FFAhoRjvJyTCTy8mE
r6C5Axb4ipq6nHHboCnkIcVm6IxG8ZWg6WFfEzD2rlY5DNj1LSagsupqThGLPM6z
KVzxLxYoBg5O0z+tif08UPj1U6T3HJqsoXax0eR1XkXXEJO85GjYkjLISEmN06cu
EGR584GiVfvk+3OF5Y2H51CN5RhMzeuUnh0IHkBlXkxCgKW7K87+yYYdVWCFUJim
y0EfjLVdPZ5+kIMgND+SKe9462tmDQbK5CXLta5Q3gzZWTocrZG6kodnPmeSr+nE
mUA+WrCmBvyb5laMKSnmVuRFU0trWaT7eUUGHsPcLC/ynRn3tGE+VcXpFtIbsnGs
YVxByGEyOY3qnuYMUNCQ1sPXOEO3OoUfFdEGPGZacWwbrjNCCCytKrxHhiAKHO5z
34JfxGmoDdja3R429H6Th35494V6Iio/bB3nqdmtIEkVSM9Ib9pr95eoJlD1i2AX
infhq9nPeAfWMQnTrfdvjVyXF7VwkIOsN+JwhDIcyDuuC3qXQ0b+Q3s8J90UZZEL
WUQ52FGZ5t4wYanIK5D9UgvZQVLq+Nu2ZpnvUhioJFGYVfZphAH7NA6fr1sAzZdp
8PJ2ywLNpXF1eejQg6tkBi3iAs1eJnbl/pEXEhQTQI5esh0oleLet9VVY56gIrlk
JNF1r3helEb49L8oGqCOHVnYNqUZrtXzVvlVFDEo1uQDrbDrLqetQ2dyNfC/FKHx
vuVXu7FwfJBzkO1eWXugxHxsMnH7l5Mbo392NPAhchKoi8UBr+JcAJlVaJLaPpgn
a/Ap1pUrfMRNArP+aPPIDO5Rxr/7Onw0Gkld9OQTHAkSNm5Lu8Y1SrOCPZl5PUTk
Tul0NT41zr3CuvCWpyto4xnV67+mg3PhhNUMuz34HI4t20t1/bdrXs5Z8G7U2IKu
xBemcUvmACFfuGBQl+v+gd7xwzjHvs7TtAF8TwqvGisuDDwJ8FRS6CiHa+QoFdW4
Yb+wKlktd4KpXXZOFcXRgiqLQt2L10wiGH+Uc0G7pSGOUWCbodS3bmZSvGnSizDv
afGF6BxV7x6zmc3WXWcTxxiiQw4sESlYJBhFHS5yzO0I3xi9afHi/FD2NF7VowC4
9TRWJocfJ06s98h1FJXz2HBr+DWXXeZyc310r9Wxmvo/i9T2kJBMG2wF3otPngHQ
IlTdpKzZi63lZzgl7oG6JUjj5TVwqlttiJOUGkmnq8OBZ761EBy7ZzB2HCmOvyfN
esPLgQbgtAevWrlT8iN0LPyJHonz6qpVDvHHdNSVIiA3dV8bu0ez6CvlBy2T9/SA
Ze/y+ECviLEBv1O/j4Lzid9ekpZduQo6VqjLFi4SOTXmKCtouqAGlD4000fMTBE6
YD2dvYR8CE00L/Ef/QJMcE61W2i9s1B1dpAsbS4q/GGmO9lyvg0xJPPR1ExYCaXi
lFW+56UIMzOu/cn8hec/q6nHxfC8BmOXkshUFxObkZxjktV7EeHCKA95DuRwB0t9
nlLnauSv/UdX9GU1GaZoAh0q/akWNd/pxlmqMceAD1H2AmAxtQxm1i+foaDn88hN
HeRMl5XleRZxRHMoiFNs2VmUSNLmcdaBeKxga3X5VnlwJUgACMzKE5WV5+FZaH7A
Ucm56YVYQIN+oSw6VhdNtvcD1haJaMW6ilUz7XZIg+/EzKzGYxxi/MugnGwGCNCv
1nDIFsxb9hmy7r5CQPDWLeZ8YBchjAmpLeoKADUMCIYWrErQ7E1Wc1ZniTyN6JGp
UVVoCUa0RZHpYSk1+2P/D7Ns0ptGLsz0Anqn9s85F4a7ueHeyL0jvTa/IdL/2Kbo
8lDhvi6exXzinuBN6FsSaHDWHp+VYguTpl8Ier3rguuZ72Cktage39bS08L+6H0E
HAUSU7So0QEOTb/bX7XmlKh1BUz20+KUpIu9m6kKEU/QGrN0w08RPpdEL9w2RfM9
6xs0nIxzkmNEYf4GBRFADeoqYsYzaacz6nkZcqZNoDHnS8ijoLuHRRwFkJ7gdqTw
RVkA/RAA2dxvO6E89u4GvutwdA6hmQPUFaTn3sWrqePGBxTbAN7HFZTPFKijXOcB
dwEF+DFSZ0DsaXiR1mmLoeL2Jr5UwDAsnD4KviNJbiHu6uKOYSe13Z89A1tauPGf
oXV29j4ISY/yrcyQ8/3VcLk87GxJQYJzmLY5bBXAUe9AlNMUT4WlgwvWnbjhENtd
Aonlkh5m5EuOoHHvuZfqjy3KZ3P2YbGaXhG0DM20s5DsGkhu5uvvxml3y/7LsTVw
t3DDRyz0tVOaCvfa/z0vBsWhTlDdXpWOGFLRJOUy0ov59+i24PU7zL/GOArJmUD/
wIHgucNd3wHvyOjAVlV/tiWfNKU4nEbivskqYBgHNzo4sDuwLmb5a4dbF7j92VSD
GHJZfNucNnfXucWKbuCclN4fpT7XcFGBnQjWVFKo6lc+EDYAznGwzvxXNqIHarw1
6zo9lQPg7gJe5tX9GJhVqQJnlQjL8vpkGA6jqZgP3ggDXs343gyNLaImkoXW1a04
cjR8L8aRYIw7UTqcBWtfkecFpkMhoBB7caW5krsBwHxFONQ4vD93fK8uOKJRRrBp
MZ8eDPcfis8sUq9rP20EqpnEKf8GmusV8wJOCIODMlKM8cKfhDZaXm3FdQmNfGDo
+5XORgr9yhxOaj+zTD0q/axBdQxm0xyFTKWVDaRUrjrwx2DvD1d3iSpnK5+3xZGA
JGsNbO/LrDcNfuxGGlS31xQevzCuk61bV4V2taGtIvApj3oZ8iC+fXPU07/0w6nM
XUU74gNQ/B1FfQAODkSD6DmBMmIt1QhAP2//Iu1zB3XC5AWdcIi4GDmHtoNa4uyB
ZNgefm3qg7o7CDx9UYhAlsmBcmx2QSY19kVkmky4dAkwGB26G2dbvBaPMPdvdJB7
U/Wq/8IY3EtB7OS2QVahs6me9HSRGxYTxF8JqG73SeNknNVE0bMxbw88w4/QjjGa
8QaRg8MdengJAtAOcdUDeCwi2EcQHStkK/VjRomYrydmvJ4YWJBSrBlIbNTP4e13
DoPn8tBcRXjtApWWA6WGQODxBKEodWVbikSAUIoOk+RlegaKZxcvm1RtHRqpqntG
vRKXJO8XNEa+verYisow1XjmB5KhxbQZ0NrIHn50oqA7wVk2oswbVH04bBYMSFQ7
Qi4hiVWDNoTV6OH2hki/yN8uTSyG7Y2pEQJgskpBBKpjCAB9ZGw3hCcedV0cnBsO
Or8hZDR53PMSk8ZUP3GDKC2Ld31fiwlJokDUCmGIJq9IqeP3Yeitrru4at3WO/wa
A+rcIZlbRbV9eCrNTQVzAeke/urbzriiiPAyg2RjhWDPiBnIiti8Ai6WFByg02vR
VGLogNDIt7HDedLnxXzMzwTQ8zW7mZ9HSwZHlwHbuu42ixnraAPxVVovCyLXrvXq
Lhfmg3+9q38SGU4KTgNL+jx+RjSDmRgXpd9DJj9D2/2pvmFD9CN3jmE6zC+s+4wf
E4ZjyUX5nLYcY9xJtCqnqvXxP7Z+vp7gUY/pttxxHqHDGebD+BJPV2gzkkMs48fy
BPFvCw6/xKq2jvWnBiFpxGzgAcOYNkmQrBaQkoY3siRPeBZW5bpof0PcKd9f5ObU
Lf6yYscEDysZ36270/E2ZYw9WuSf3djTNKC9s9NUhI+QWgGLopibZl2aRLvy2fWV
G8BBqrVLIFnqhZrYl5p1zO/mKXbXNceMXeFj/CyMJQUkorC8W0UWvrGstV8m3PYp
WY7ijTvQJd1L0WwtACWfk3w8gJa0XGRgLWwCzN158uXX0RUIGlDYY6ZGwtSKdFOG
k8Gdqsfd3rloMX+AhibrDErn/vFtPH0DRsCz9XSmoql5ee8q3mRTcxAI0BCjgN4e
ZeQPGB1qWFU7QWrZPT9luXiPpUmNMWCLnV2rcbxgjaDXMVYY7KB7OYMVXBuo7Q9i
kljnzUpDH15DEOWU6i3TMWAoRvEFD7KwS7JoIHuENxCBEEHq/gzifqkhjDbe+Skt
cq8/SOIrHCLifo8NnGdWNF+JbO/d0QOkc5W+UyDIDCqUs/l859B3cBPdXsE/TuXH
g/sZtUJl+kJmoGyIkiU8YZIPJMviTy4/Y9XEmS2A1GUGXBUbltUW0IDLPZFdnHlA
by/GbQUpjsZeVJhwH/JzogvvQfhxmxpv11sIB+rQ+Bsla8wbdX8PsXH9M7png4d6
h9Tg62zm93/kEwbT8imVwgSxbJnC3Aa4qAUYOGQbPp0YcKAUBPYJ6hTvevn4I1dt
qMoRrb01GW8Qy3OfSd/Hizs9xmFHzgvPZy2DZw07UD7RQpZ8xAlOBUXeB6b1AI/F
o6SkRiUkQ8LPqX/mwFDQH1/8QVy98lBujx2/VVNF/2W+oDIj3NaBqTVOFfNb0HAE
t7TH5slNR+RTWBxAtiQYkP2uKVTny+wfpyLDSePmQimrxzy31Dv0BTl8HaYIf4gD
T82vc3/hcV5gvLtzCI4jd2ITcvQaVkfYAsQiN3I20Sfcma0rqywWXnOv9MDAugps
7Ct9GSwjoxhkldq7CGbyYTwTSTqZ3ke9AV68XgdegLE2nTzp+3+KKpIPfAec6J4Q
13JaRCLWZeJZcsD9pCypxnyGcaZaiXCg2VpV30Y68Qf7HHJsgU4TGNyQKURt67jC
Y+jhJSgZVqKMgbLmYHG3c9m2yd2GAyPP4DWRTtx+RdQkPw0DXDygiZM1BylvP453
h6uN7kf9rwkt7wVrZRYrOuqnmLZbjpmLSLaakVPWZwCIOE14m8XAIiOBYD7DZSME
L+OeR2qY+Eh2Sp3Rcklgu1XiwZXMqmSuX/vOJq8/3PptKkrWgtMW0VOk63IptOgB
eqxgiBHCmbcASgYZrnx59CI8x/wJjfEg5IsFADF+uGHsf4/LtNIbKyxulRJ+as+T
MKym54VlrbFlJpnM3F+pzTD+4eS+ULmgUItzV0Le+fNDah/pD6ssWE85nIfHgLdp
YaUvpMBZMNJmfdEwBzvlftgN6IfoWZu1lSriJUitA08i+RcmVw2r87Oj2XsBL+S5
aeyvL0v787g9T0Tsu7XQJ6YnO+Zzehfk+I0FqTTzh/k//WKpOohDx7rxvla8TKm7
kYa7Epjszjisih+2UcTTv+DQEniKEwyZZFkhoqHF0nUZ+0CzRNdlgWE/rtRfLxCq
e5IfDxUKH/vpW2BxpevfTYC3nXaqgl7vIX2bPipC7Qw5ZV5mYtYSlsWn2qGGQavz
qRHdZY+wUS72BbnrqP6zoXReNKL7X/bdoGXlWPDw6o/1ADZtUH/uetIRR1ncAwiP
r0us7uATrwmcH79KBaW6wVwa2HUfWgWyg9JXqd/0qW4i7I4w283X7ZITi/9gydW6
FViA4/FuGXSrfPkuway8AnmWa1sTm/pos0NU6PQJO+Tx4QhHhtdL8/KLLidJ8oLU
u0bI2rMcBAHS6aJ2zpM9Ce/qyBuenjTOaNe+SQDx9ADXwcrLgeoo1A5H+pSk4OHN
Ec7JtXQh/u2A23sCnmRSBgEdnX+ymJCv5Mq/oQyxOmoPIJcaBZySCl1uTouIuO40
Sf2fdhZqBD3bgiPGIz6sl48tBFQWzIZ83DX7yjFn1sDr237a/sZbYEvWSPINUenr
uMpF3YlOPpAJAbrU7YFhx/xhzBLegxapgwdJWhHBSwQh6MjKnkWoXbuQxQDZorXb
evEs3OMt6akzbquZrsMh0GW3a+fLkW1DYykZqyPPoH3jt2ii0ODVetKFhIKaXu8W
q8XWX74MQIbVwrbLf/FBONMRQP0zhnGUt8+pATEVestPboFcbpxgExjjm22J03KU
8cCbVUltE3K/ijXlV2+r+K1DVzsBnTqbEOKo06LaLnEYXdIwHM2ynVaNgFVl+ClL
i7UR6IvroQDXAji12DLL26/7VihhTnnGdJohXVyKJuOrM/SEkRBAnCftM+ERD9AW
MATjY9qLpeZT87BTEyMWEcNcw27hBSBKbNkIt9L99cr7NLTUqByLsA1LbmOAwlHi
UKDnM1Yo0L79mqzCBvjStjLmKTlg97zHzBuigREmDygvlr9uOT4zAhFI+4X45zyK
QqzQ4BBQ0jD8QsaNTJMr4+flJ10jM2NXG6sy9ocSZpxvpvEP3setB9ijm8++UBs/
gY1lQlLBRs8rPxVRL3I/+TMfhsBNUm80DMhEx2qBShnfPhSV8WhQHlIgLuNSvf/k
chn4J80Dvf+gpGkTSDhl99/KIqoo1sPVXSG7Y0tjKZdRPkyUW4s0nnGfkLuvYrwr
c5w965WuqTBYKZlyMuSENTf/tor7x+QSRzlIae7gyqTgnZ6Hp6jP8RmiNnQvFrJW
fJDEENfKwVtuMfwdr6dD7sZdX9iKLw7Cgr4O7JHZ8kAyGjJUAbxSM4DgkjVsdsO6
meGGz5r7jQ4g/WSGfJaCauazkHvlks64bgGn+N/QHIKLhc/MRgujFUX/T4Wg/Iwt
JuBGYdZIwlI7bhrrgq8Re453osUOL/u2gwKwncebu7GVouqw5pA4vxZXz+hyZfUw
lDvmfY2cfsSUxWMczGBtPsavv3nqrsXlQIyk3pF1EuPS4shmfhiV5h7UwQEzhxt6
8Cm10hi68MzGD7BeDhFXfqu2tB3UHHal/bASjr7iDpP4CZSfclnZlRiqfOTxsM2j
SKdLGexEJK2x0d4z+AUN4GwN2n16sPU+kUdnmYHjcx+PNZrqsoIb9a4TcQo9Q9aV
eLjeudH8GtCpKwNHkbWWDeiAo3x/hsMZHfbEtvEz2gWWt7OqhkrxNtDU6xy+ckRK
SzquzgHsjwEmSF4ziUMvVJYM+6XZxwN4XjsBUaKyczxSplivqHg65phezkm/6NnI
6wGSIJ0OsGxSNODk8O2TjEtUBSKPPnjP3cH+X5CvuMySiApvG2HXM42zeODmGm64
nUZQpXUTzoqKFVDlfmVUldeiAcP6rEV35u040SXLvrDGAW48wnks37Lr66J7qlSZ
ZVa/hkBZXmlUqjiVJKlUZno35wVqLrQJ6sT1IxnGcjeRzcMN+9UPQt9TjAGV/nRk
N7BA6oJwjsnlHuatSrlndzsO9cNm+4IrjY9OFcFA8cnzXG7OeKiLdZXTNBGddCzm
b3DUfncVp89HIdcpQJ1MThourZkTu2R60fobmCCyiaLOLx/GFTum8RlnSTJG0Mi8
33v6+OmfmldsYB6WRAQbWqoQXBSVvjFu1FppjuOlASgTjqfPEEbzo9MWWyiSJvvR
+JYf7fVtQTXFaacOugSXfxqFXOn8ZoNnLBjqI9v/js3OomjF0m50EhG0/uVI9rSl
JtPu4UEtxlAPbppygBcbVRM7EIUD5lV1H6+9bI5FvNtfbNO1JSof9cjv3wPtl9/p
9PY1WZSgvikd8+hhaZyAmxpy/q5y7Oml9VY8TAHikyotS50dMSdGBhhFn2YpKb3x
De1t9oudvqNeowAnqlklkuo0KpVhMxs4ioyRjq/0JI91WTQXerY+DeCKyEWYcOSD
jnZBXDtUybrIXuhosk95uueYRDIe3iOxC2EoSxBKa5ZDqX9icj/iiWGQ9EsphhJA
PgJ3FZvbbX3gz06G+1KUic1olzVVG2jgxe4zDVBWXrftHGEmnq8h0pscguOOYks/
Exu+HjS+u6vMqVWY6CQLyfp3THtTp7++ZGI/NB/aMojWHDah+mOmMKkCuiLvrkOF
AdBAVbhasBmt85VhKpmb1O1MrIEpFG/S3N2rjz869iXkPvqlOT0zYXBhm/+43UW9
X4O4Obyl0lpQ77IqEVJm8ClNW9jLEnaMzXKz7Ds7sJBKXzoV9dicZE0Hq30VL18a
VgkKTHGJrLkaMCJHGrpGWHX4oMELIzWrAFGzVQq4rYYf6wDW+qq5PxyHc1VnuWA0
lv4jmU9uQVrbGsdDvhAdLmUGizV32zpuZ5WEvuaA3F2ZyHY3MlLgbdppmZEMlYw6
BB4ryrIHjTWAKVjHRwZc9QzosVIvrJVGEAM++E1qDz7yXy8VfwDrlTaiiQL1PT/6
s8tqg2JB2AIZFDabgy6aLhhfUuR5hEnXNcjlJ5aGSNXutHFyoMHtXf2meTgpQSxp
Uu0sMzUOIbIIvkDTCW5aG7IWvYkCG7zJV+/qqO+za0QeAn8u0U3NZFAHmhE0AApn
2AYfpxiY3xNO5vEfyLxLWtx6X2ROmyMymtZI1xFBU3MUYm8MUeYL4C5cn7KUHQKG
TiCcwcVMyyVovGXeSXYCWbceuWH6hbiSrsdLCDyANLIaks7qXX/WXrjKucn4L6vj
g6sGQG8g6r9ca1R0+8Qf4FKdX2H2lUufs6Y4O44pGeHFLrLMkpYmCWD02eSZH8nB
IqQl0xVxczXkZ8EzbtiNBdMzONYm61fQjUxVhXeii7YYRcksqHk64NvJuP0str11
Mv0vhJlAO/wu1kx4m1rjGExvEgo1wz6cwOvA7nAFgmUGPNxLoSxMLkUPIkL2ZB4M
MqG1muGNx6oGkqzGDSN2Ai1/+yGi8uyYf8O+CSG7XYAwqeEa1cmQBdz9j45ni4cM
mZDsQ6R6psTEgABISfZV9sozA5Z4WAhlJKWShPzwK41Cjg6SwPZwf2ck1sawRKYw
b//FbFXqouhaN0z4156K60h9E1T6p6q3Jy69Of3jHnUK17GFWAnzmYExjOx8P7QK
FEN8rVvYwTLVGGGYHYajAOYRtSykWsjJrvv4A6iMhy6lBgn+/Cw/vmlv1mMCbaZm
ZYrjBt9hTCN0S2g1lvOgHNYe5hU39BGPECiFxcE6CG1RnUdtis4QtjQr5zH7sgWb
aObCK1Wxuj4o5HOFF1k0gZBYp9f/OTygKhaVchtZFaQTklTzfjrUJNf5F4gzaVuA
6aPgwKhgvkBY5cd5e16oN9bZGEbx0Omda+7hFq7SapG8fhTujZrWgzdDiOc1Si97
5EOBYYVpnoCWaV+sMnbbCD6SKYO8peXV7oU8RwiZa3Z8XGkUcA3g4XQ2kWKSa6ni
2Ex8mRAnm0Hb9fUc6B5jsVOFodZRT/aVXkcC0dANIN7BjWfhf0BsZziqa/cBXMlO
SJB9WeLnK1oiPwAJ4hZFcHiTKy3i3Yd1dMq97Q8nubRFcvlPkq98SrfsmoGoTNYb
9ulUR/X0e1c/W864QekYjkSRuTsdljxKW/WnOtyupM9mNUAPx9ILq/YXJOeLT5ZL
/mPlWlV0VrtoR7NWAwXAeILXYP9qtaW8ik6hY6ZdSdow6dbhvD6ppsLRN5YpgOcr
oqsmZkL/tw3j6+wPGafCZPEoUV0ru6swTJYVfMKXUDDN85QD3XbMUoZ1IpmPp48J
6GorTHzy+WfxpK21WRTcAXwI1hO+8tYqeaG2Yoe6GtrvrRaf1wiUAchJe63zOLyJ
fhZWk2gT/s69KHCgx5ewSmf4wsg4ne0W9ncmWp+QaULjPHWs8ktJLpQXPkzSIzlf
6rIg2VM1UwyMerEWq5zzM/Ks1KhVMp7UmBLFHcWOZRGYDk4zj9+uq0NDLnS8u8uU
YTI0oSEdQXM4Hi+6R3P+xIbyuUOHK29OPbiEZW8M3Q1ZkyZy/nnao5RHm0iJshSE
bG16bE8RR/GO4Qqt8c1AIFpxPdUzhRwuRvoUXIdU4kZgKnbG+Ifm9RGSZ9H1tFyw
nMzZUgiuDbUUMmbavZAGrI6W47F8JVAW3X95jeAudiEiS/jKmas+ItyPdlJUKjHJ
BbLEyn+c+VxiuboN76U7/+zZCXeT5p5UdugUQlTFtY0SoPhCAwgAp70sTqfnMwLc
01Hwe+8WrB+DWwEG8xNxbJ4lXJ+b+pcMNRORxT1CbMblxfgkGK0BX9AT0s4AX4j2
crVhIhGTLeDYvzswm4rzBLFMZCnWK+8RvwwtQTAnr2KsgSLZ483Myyf5NNYSfVf/
V+MPpvtRcx56amNW6sYc8Y7z+oZtzXbiBUS1NWIxdTsTgufKQMRwR+C5sjHa89Bh
pVTeal4OEJsaJJJD3YwP4he55KrI9MIyaqOcUQCV2srPF8HV9v90XBesq+Cwkmyj
W8QQNjG7ZojDV/oH9G5PGCbOMFi1qv68+l74ot99npcfJbT4Zw4Ed7KGrH6fJP0S
FjTTs7IctIKAx7jiglErUwD/Bxr/7KkRgK4mT5XOxw54uqgOb3EmYlz9s/kG+/0Y
yUdcJEvnApKgpwuuR4iO1ZzRs+LB4CQoE3WtgEc5YnGanJvGMgGYbNH0RzhxiBgM
3vKXxUg1DWVuAXbCWg1ifCQbkl7Bfto40RD2sGeTBOY5HprcsJqTUgTRciVP76+J
P+9Wuh+HuUGzDnS9x2oBRI/Xc26U3qfPQCqR7ivDdYcGNSF6n+I0wWtWnJEEljFL
CjikgxVTnNK5JU+cukL2B65fFjP1iKO49oHGT0lXW9RjD9H3rCRWVUvjIae9+chw
FvymV80veuDzhUt03jIT5lVXY7//wL1X5xkUIgC9BnawLGTCXOCkZwFMvxTMqnMw
TWOs98AmzFphIgYYdVfguAGnJtn7zXCE4TFM34jsQIHHan8qAQlBhSlyLfJ9BXjr
GgRfgrb2O/cYTRMIFU2yDshzF4XvartvnnTGMpNWQVBl/Xy6MI8Mj4K6afFywqDJ
esWJFO4WCTA4ucj1RpjoWo/q4OoLbH6FCJ1bn3syz0KxDOtvkiksllsUC+1sy9rq
uke+/kUPyx95r+kgsBGgJiGCNgJhJtgW/dnsV/Mbi4Z6ucfY2fK2kiY7n8QEnPFL
DsPh0zQHRVnWYXdGx5VyJkNLklcNJuWNu4PFCDZ3Mm4GBjPqZUQtWmPq4ByfehkL
7m1IyWlKkE1iJgZ0CEgpoziAMHmKv9DRbvRkXHMXPPMT+blR+a8M5tsf4RR5fFgO
gSgfCUa5lSGKWPx61t4Sy8UZi8QBL+jLQGRkbWtop73TmTCmBby65Otj7bxngSOQ
YIdTQ8J/6xfgEXZyEIIzP2LVaob8Y4PCQoL70YOwbRdvswk/mF58pNwEVB2Yv/09
Lsq17KO+dI8fOwssyRc/PEqREDClEmLc+9MyqVJULksL6xyPG9vep5p8UXCmESfY
IXhFeokiydBifHbzGbY1tr1PaDMIRK4mJcaWRxtdWAZs3Myr5HN9HCLiVWNub7aD
v3Mz536KFnrq8hQJIPNE3V9MzwJMztmio+oonYswszMzWNkGK+VHA7d2+SkfUAtt
KbWQudnGb9/RQAYGh3TO7b8HUzU/indkKDUsi4ddrbd7xuCm71I7spj//QZOxpPI
F0SoCx8jiq+mXDROu69IHefHCG/KsU1vYLdp/3UwlMHpMAvCB2CM+m+I8khbZoHh
gyLM8AqaCxEXf/T42qzfsLKAcTF53OD4wLtAKxo4/xBULNc7Up2+1oUBgfSuZFpb
FMdLViiX8wBAmyfQ21LM/ruaJ0ZLNBXqKF32en8znv9cKE5s9sQWf/s+9Ihx3QaI
+v4MbDQ1rmWAQ2MCBU7jDeaFCkcnEdFkRVdW0T4L5rOzcmLGO1fBMk5f58yx1G7O
5JnsMDr3Jloh9N+71uYqNh/ibubnTvcmbTiHpUgBRupZKLSCfPTaabuMfSJDsJFW
RltqAXx9X5viSxvv6AsNej6AEQsBYOg+t5FkRhr0MnSVvRM92WREFXsd1vP9goGD
ji+nc5G9UBfNAFs/jsi+vXGArXtsQKDQfzDj+388KVouqvt56krD7hc/7BjtwsyV
MZKR5eS1s9sJkbLS2BgazFOQvix62KF0Ylud852qEru0g4LV7wpOZM8rH9l7svZo
clacv/YfuKNX/3udsDJl20cumHHLfEDDDUPZCsJ+vkvU6I0eRUsLGFGjzKarGxi5
h90cLqvfNQIdvBSpBcBGHqJg/SW4RDhmWdDs5SeDpJNYmcwfzJqdhSAyvi2n4mo9
yv7CKkHNWJfe+kvQ5EU86Fqjugnsr6qZz5tu/PDnGXyNGUr2unk5DNWAPorSuVMY
n0FlvsaS77jWieWocx5baUnr+8VP9Omd+yxh0ISKRtYiFmga8nfIeb4tVKGclDv5
dQSsaiPnf1UAzv22mWplidWXkB0pBtMb86H5ToO3MV/MZhQ447aMcg+oWQWLOgQo
0KzQl4tnzQ/W6vI38VlYfnkLL2MpxzLFBRqsTMJTqwq5zK7nuhns4QME65/rvr1C
KxygrokEa4ONeiQL7FWscz1sn2ZnVDH4+wzCgwAxyRTCHa6WxLIFrQM0X2f8tZHo
6QUpRh3RBX5b8aOWfurjXMbir+sSX2rZh7jWS0YOcDszxX62FZPay3OMFDNhyO2M
GgGKe7ILQRdFH8ilBFJbyxTYeXfxejCYQQVLu+1yW607JX5ATPFmOR+I6iEzYbr1
/1WSs5nrDnzpEbY0iXD4euh1eoDzwen6Ls5KwtqoIybBwg8JNl1GkTdC8AlO25y/
rY1CBeXLlWo5pNnfqzlr0MqzRYPvB6mWW7JYvsW2wUQz2FPuQ97/E6CQsaxRAqhb
ZM6TcY4xnOvNYb7cifVF/Xq445Ui9bdtdgwWGHrQ0PqVKIUd4CgzwO8ETwZtxh/q
KPdczqufi+S7UkCEOA5BdrCiyWBNilqvkwQof/OE53ay3DjSQ13dEGyOGZMSpIdA
Nx2AUWpbqcya8CO3pFRy9Zkr1TjFxd/QuwdcYxObXwwlm7MklZoj5xfBDELfWO/i
h2Dq5AT0VQA/3EdKcZaoHA7Z8dS9JQRnYE841JjoRcpnZiUs6buD36w2t4JehgIP
m42NsWDsJWMg06rSw4yalfcRwn4qj1QNcAw/dDE/QkktAWldpkGj/AG8Q1rC1D7D
0NIcDwGPAafVUM1SMoxnm88TcDie0cPjzC2ltzbVqhY9NBsqxlG1fiG19wbWUJfQ
OYEkhQsl1gync/qO1ofnBa7Hm+mbe1UGpwCvPH4N8F5b0KLjJb7mKMDZfpN/plLv
/bq8WL0VxNa83EZIpxAg3DexhTN7ZBK2o4sW5agjSByvvrm6JKtl70/lzCYNF2oP
dLTx3J6mvEgIQvxJHf9Xqjafru3g2YzpXzT6O3pkYKAE9/wOhlO7hdDP/qZt/hOA
vsIZI2hIqD9Av2KudqprpyNUCETW/4Fx7+BBor0nJ/A5A9Kq5ZoMoXyQAIKTF5MT
v2FSlMNu0yH/BdmuNxbuPpfnWgozPdMuphwZvGVudEnDPjx8z3TKNrEFw/bQIVaU
mZBZey4uUvXV23l+NOhN62L0SKAdFQ6OR0Jg+zefpVx58aK7DEnbtzkAudvPJ3Do
RgIEZVkIgwbqFXVquyLNEB9a2+rn4TjV2tJ77uGMv5v4JzvloJ2yXXCvZXqRLo1p
g8QG60dNtiAG4z/1rH6Pp/7HsMtD6P3boXVB4DV9oF4rok0g4lsfcp6+G32q4Sf0
AM8j2nwm4Pm6UEf7ZYGKVfBhA1oAWV0inCxmYTC96BtIchOuHnXFJVRv5NWX7vc7
f6J3Xkz/UI4sv2tee7D3V7ES+3hhYWkrqLZnscBKRqMo7CAWPrJMRSYkDpaZS8Fu
wsfHO7lsBCpuxfaxTOBYapslqISuzwuRQUfnS5asmIIsawhwwc/yedFXz6e1pIWa
MySf4arAmneKoRsyEVltTcwgcRTDVCW663uLB/Yu/fi38We2Qw04Okdq3FVuwhu/
FFE1XWaIdJgLaRBijsaHNvd+Orp1Yh5I7kJPTXmfYTyVLTvgGacxYn6fYNxtDcun
UODDVeb7D2qAS+IIi88SpsjlIiR58hnzJEVbruxcJcjkHpjl6XrQn1c2Sdk8kZXK
dnr0iobttL94KZS6ZqYHJOgmYiUC2d9XtkdVyilkPrO2E9JQaQHdIs46aLYsmenk
lihPn1U/RWxZ6orvhJztpwPEoj+tfD7SzCqM+CsGFOclqC7dR4CSf2QYZanPd7sf
rYMRTaSkvGYucUcdSazUptRqTB4wzix+mPEQL4c3yMn6w4m+9bgg7rNdzYqC8MB0
YKvUfqlN7ZK5aPU70M1NVAeAFnom7t/zzTdLlDQ8hEvvvpDlhQbodMkQnZSmfUCt
amXUyGQiIEp+A3IuuODCTgDTCzZ0DAr97eDvt42tJVn6gFm3cC+vyppt+3UfLF3u
PZ2MTzVTqfctoBryPwqaoR7WYb6ISiEBiEV0+4vl9l9lths+0kHine/XExc+L20s
fx17lOemIBpaiCfk4GRsq39Sv9sE7GUr6/dOfTV/qLsEten8uW7V4NPmvtiR1zar
9XE9NHvMWlkHqDxRkxRQE3fBDbknw3LZ0Jiuv8NQRi0fBW4qv+Jogg7DO5QOHp2n
4esKImxFEEjaK2wt0V/adBVmvr0dXDtEoOZn1jDhl6EwdQmeSiMYA3olMk40L61a
abKhLjAGuZZ4ynBMFUM63JBn9+KqTB+cH8Z8Va67YygpGPcdVDOe7hQh5wrNTmRs
w9eGvD2Jr8DS/4xcx4WciLV0PHNU/WOfaakzThPYth7HQAN7uw6+D6ROK5j3v0RD
qxdhQ4/Z8AzxRDplMBbYvRKsssxOm6VVeLQcZjtUNpjW8H8dIS9ywe2NYnGlYwX4
bUy8AfGGAapoT8gsHWc0spbfFjkBXqpKnVAztMdc8fMhk1AriACwbLiq5JLWr5SJ
tkOW21z/ezlQctscBdRnMVFe21QV0jIwotshfHtIyeU3hsCQVD4jmJjPFONYDQi8
Uh5QC+54qIrItt/HcVoNcOQFMzzGcLBLQokkgYqfpgDDPA0WyQOJFhZ8fpwckXUh
BMOvWrePKe980HZpljmpe3O5hVCG0FO3ikHCsTugtE4k2551piPtje/Hl3rWzfwh
IGn6UYeOSE12njS7yAIGS6HCCQTICBXX2svpl/9onYolnVR/SxlM2ZXDJL0Eeand
KE1mas54oS73IOtFFYE8kpITePCfjGLsjkKpWVxtZs5lBHYMmaQQzHRVJ1UO5KsT
89HqmNH9/GbQJV+J8ZQMuGrX+rdHThk6lvrNs8gH1GyKLFsnotjN7OeGKD3t1Ffo
ud5QJMlGR2gSvFsTE/N3vt4F7iGyPTNSEpBt0x/d6xvdpXr8r2135XdhiP1u2A1x
ek4NIcRNQwV+yRdruXaZo11UOktS3EmnYjjbF0laTnah7/Ndw+7jHCWUyMlfcHqm
2V8cC0MrY43WNerykhHG0E6JxGIiMmOPjh3xlN6rftTnxI8trzA3v+94MaPTHi3y
bk0pyU9kNrH/mywApd+7fS7wj3dmRweY2sK3QyhGkxfuCwZHT/6RGkZHlEZcT9m9
YqDsufcEtew/hfl+JEoMTwoXg6et8Jhyvw2bnXuzXZjS66ssYrnwoQ5t+R7hXT+z
haCRB3mZRLI/XZ8SPBeBqWRPNxVabwGU2S/JaLdorB3umcoI0Wx8EEaSZVEMfYNJ
O9W/cZDcqNdwfqYEUc5FMdmJ1Kytt9+BlZF1KNmJgce/NYOe1Ejq0aoOhsNgPtZf
xHlXWQ7BnceLZNS4mCQCx7HDytYnoPnLeroTVODRqBIAXL73J3v1fQrHJO7eIbbT
vVwT+2fOlemi5pyHYvl5B6DOWuQK7uqvfzzoNFpeoQi5PA5sFhVdutw7UDAD7enX
rtu5S0l8rMbaVIsd1AtAGBoIzmHWnuR8gjZoXzg6VQsZZD6iexysf44DIYpqqyHB
xnB2Yte1ibgzFcXeqnR5NN/uybJoIq4mQbbImK8x+aP8xDxUGy3AbdK7i0bCLm0l
M+c20C7FDDF1KXRsbhRSPNGNXBr4Gvp14ZcDyrcFsdjXaHDKSp31XLi+W+GhrLob
f94qzu8ccO2j/ZIM7gvdzpDjJN3UsXtzvlOBXwFOwvz4KnKJQLXakHkXbmrtWtVU
tBiVx/4gWc3CiggJs5DKKsIRuNwS5RTaiiWkifnwvSsdLLbTcqqcDq/I75L/X/vc
FA+CY80r+9WVZc08eoMtJfFARqW0a5el/h2j8+RKbJ8LCs7YkiptFoSFJaf4Q2VO
GqbCncF8DsA0GMnV3Rlaxn0xpRouksCEzhyAu1ew/UXS5WkF/YubdENO8olalHKz
WFfCva8yrpJGwon4BPvaStBjoKzkaYvtO4Eap89qx8tZedgNecSh74sG58r4St+/
YUvmP71aO7ramrg+GA7zfLNXsauMtgVNTkwx/XC7vgkqWpHbgpwGTTkK9A+wvsyG
`protect end_protected