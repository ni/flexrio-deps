<<<<<<< HEAD:flexrio_deps/PcieUspG3x8TandemGtyInchwormWrapper.vhd
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23616 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
LNzla8hJ+flbI/QoCi40dQS57TBmcv71hsqdmGY9Tz3KwuWIIsVzo9mqzMam90xl
dzKXef7lZvI3ykttcgIOPI6ZyfEwqlORHnKrY5k7srD1pGUnqb8BMiHryV++h6Dp
YfbA7tOQOwerL3rV75n4b28VBZqp2Z/dfqPMuOv1hff0w1McRk/eaFNjwmWrY0aw
u2mvos1JCeZnngy0m8sQhxbtTc1eKIsrpLrT8Uc43MhmLV1eAtznwyar+BcqRqwP
6bXW8YhDY6ElRittRbXjLPWxMoYfmE0gGF7RzfjaPEe2E5lw1svxp+7Ve9daNZ9e
F2IfSPvcctE2+G+PIGDF4ihrFJsb49lWQCUFGYxU6OPoBJI6qua6DvWCJKHS0Z/7
kSa5zfND4vQ8BaKQz32/qvY/qNpeUx9enxksEE4n+62ur9eXkZxq9rNGtajZg6he
NIBdUFet3qFrQJ9Ok0vkYic/zlKWs/OHzihntxIQZb2i0vVGMrMkDc3QwcmOJSbL
wbkmTjbFxtnp8gmX7W5k/7RyZOOuaBCccsWWgAZ4u9GwcAJad6PRxGiMIAhzZF++
HxR3+/Gb1fi1Q5F4mYmBR3MHDqeQxK83DH/1iNTAKDqpsqiVsKd9sDBHFWRGN3Sk
SYgjOWwOme83YsA62YX2ZKuyqu8S4XzXGGJG76fmheqyY+dmFr9aizUmlbgfakfl
kDmnNhkdlLBAYntUkI63tJU6cQZMPkeCtbje73YS1ovKGOn+XzmlS4j8vjOjp3nf
YeuzFxvrcAxWCXV6TepENzCVmyVNg7tF55MMnayjtk8mlyG/MHs7QngN4QOWA82Q
lqVIwGJb9YUCJobq/Wg68gyP4JdTzgZrcY/n52u6/7f9ZiGrlLa93RtGOfrDDYlg
QGacp5QtTlghBPegUGKUnBvrJNwPlZ+5MPA/DxzIOlRbMf7LQeKGAiW1k36LgoEQ
cwYbXB/vXuU8T5t4E6oiImgOcPsEjIlrZXVzmzc/u0dam2sY62A0taxnI7Eis7IB
cHvbykKQTKcwMi9LmSyeN4Gr+lroQhYEwEoRtfv0vSN3Dg4AQd+utrJn8hcZEQ+H
z1e90CFEjRclVVORK9pnQ2LS+1T1t3ij/x1ydF/bt2xQRx9LfY1LwIB1pOEpjx2K
yXAqP4i4yCO/h+UqIFMfGDuAuc7H7Mh6s4T5xorafu2WW+xTTCDxKcxSbqZXsp+b
Rm6iSpAztzdH/DMFEEYJVakTWtReJshs8nfdQ8KB2hurh8bDloxIoJU63WCIbuZc
c5uuPzXel0VVSbWCGVRbWWO04Vgo+KVmpfaQPNRgZx83uLTWl+SlYUpdI876Y7UG
DrJeCtSitWEx9t+MqAQRrGMDB/2FXmP71VuCh8AtHAqjxvhMZbuiRpcyEXPu/Yju
fScNpTQu43SS95lKsa+Db8cQ1vvBPCeBNUe9CWrVZ1Lqw3QCaUmuE7mVd1Efd4+X
CUCd89dJcTAOZm38aCLM6E9/SX93meSsygA5lJvfS6UYqGoKEaIed46DZA5UnYWd
6IIZezY6vGojl8HaOa+xHpdqP8jkHiKNi5oz0E5P/CkjUFGywxtNQynoOnz8PL9a
CF2p4EkdsJv+Fo5XBJIARqq/Dj9Rhx3C3aLyjvsc6fKgWdvo0FCFz1tSwb3NWhze
CvqphvgFaKPq8GOzWnavhuQMq/imtL6XhL4deB/H3NDq/pe3AwyAwDecG3IRWaxX
VTvhWJE6CJqeN9EZOlQW5Nwx5w21mekMMrGzmZaBgfL1ET0Uc8ggShK2ps/z6o8v
oEJNSAYx7AVqev5ypOZojMErEhMzIy1p2p1IXqdTMRv/ORJFYXJ3mCPCFAph445O
PI2YCg8iK+Y4JdqUgnPlgouAN5Jn2/TuXFRwIQtmK+sW87XQ5n/3vThUSvGUGwBc
b7gkvL0CqL++hlS1mlin29qrLOy5aBYLDtvrbjTuK5/MpHISnAXxsZUK42g1KEMe
B4914xy5s7OnMIvzHy70+qkZz82lDdzDeS/0GVqlq4OohiGGtSU898mwYH2sNwgD
vRq7WHU4nLSbMiN2HVrqtJuiU1ZPpNGoNlCIOZ516a5Hs/HVMJQoPDD0shXKSAXX
tHqnH+PPhyhDFvUn/Hu3hpyu6iwC8LciekIjIMMdDE7X068mdLiWKnmyXLQowoUz
oat4ygPwqV2gp4XBvTVkARq6v6G+F5ePRn1RFfy6UUPFJ7ZUmJAkSzTMs7Skf/Xs
N1zQ5rkguVoJmR1UB4wVkhCRq3dk6VxeCyVIjvfLVeKU7XQJVMD2XvAkkSfz0huN
ZKCVfrzSlHkwU/U0ryn0cCFZF+RQn/bFXz7c40fP2evvBRQZmBMCjwNv03X6OSzo
2fiWIbsnvyeM2a1wsZEjNqb8uY3qGEF9HsKetiXuCS4Ir/MTxubAhjFEb4z8xybk
XNxyrtH76Gio+cTrH4+N7DkF2G2Nxs2Fk8EYTHsluXArPZ9t6HKMpuwPpcxj7ORV
i1TlRguOF4sbz2XDpp/QWip7GuIFlKj0sDbwtRjQdEch9ccCrYFPgHiQTIkXkf28
mgkQ1tvNQxhcrZjAngAh4zlRNnLBh9oWlKMaH6LqFuLcksV7P5YzSMfhRDgNVsi0
Z8i1xQc7y+oH1Np+fK3FWiGF6J4NlGZ3j+GFbv5J+NHqQHNF8qQ/9gIPaQyOtwfh
KzjQ4hXSNpmqFvKrUCXiAQD9vgp8Y+udUYK2o7S8czmCmnY4aplWhrGkSpF7lbgK
9L7OmX0v/dXkAaatNnQP5wsMoatC8aqllEAgkTMxCPQkTZR9I6ErxgKeVFNjrxoh
Dgb+9CAHbGP1yyKLhMV9grIX9OBeNX+ivalmw0yFqWHTKcOgWe0W/I2tYcupeOvo
12LKJy0szuPnxJi4wyHpNMnQTkq2IcV2xIIlmItw1zrrZnp9WhbUy2EKeoqa7Q61
7XiqXSyDC3V7IDdmAG26CEkT8dAl8t1KBJgHqWvYsMDJtgeRadLqV+AmX7HCXwIu
2kvGaIQ/4BWqW+cuPS01vHUL8cAcFEEl3IJ3AACXfjGQOghITKv+UdR4W9Ybdhbf
8BmbXENQxG+sEsWCBezY1ddfxbNy1Qrwl2+mGLB1SkPRBObd2gTGdSX8FOp2cAS0
/GKzYaao51ftBidprVQ2ODqSdOXbXGvcI9PHIybYDp9u3TedwvaS2jjMcry5++DW
bWdKDifFv27ADQvmF3flmXdKC2W8C3nDgAosUXS0oLrA+QlMALTq4a3f0JikY38F
0GW+Cp+v6/QkdloJJWSMSo/3+64ANK7FVeuId5jVAhMl1dxKBWNsed1ceQ/3TlDo
AKQ0Di3j98D+app+6DgY8GdN2xJ/0mS/2og6roQDKoot4rUJp0WaYjH0RLg4aO13
CWjPDoPwh5cN5YHx0ThkR4lvAcYC9M5tMlMpXrobSSX+iU2rKlGLYyyRJVnZM1ih
Lpb/I+dNQWUSdqzryFQR/r3MN0MaXBqx9h6ZfP9R60eYLib0tohzKbTngzcFFmly
TNi+HCA42y2hIMlx5wfacsJNB3nku8GQHSASrtD3mYaFdAuj7LgIrv6FEgsuTZNF
MFEX3akdV27d0uVLU2br3juf7kPV+a74rBCI9k+1AebYQ/KrcoBJEwBa2rr+oD9I
ICIeb7q2ZynhKporh05gW8qJC4jl0N8QUXFxkxKIsHSWefvk7T3wrMMl0UhsWGQe
IFmzlTwhgzq0FX4CPqQsvGCMdGAEnCL9BzyMnBogmfpN2T0IqDgp8N+2hd32HNY7
IOIAc9QbukcuwK6e/nGsXvyWtWPf16Rtxg/WUADPNjYUFB0suK2n4Zy7IWN8VqAo
DRPzAXD6GBlptX1A0MIXojdCrlLWz5g9B4h8GCH1OMHgORB4p+ZbBTzsFAi+QdYO
FRwJEv3OPfjYTtxjIXxGozP+GKQaX5JMl/p5gSd1pvzcTFeTyH3ZxmKCpVI3sDZQ
GtcoG6bvBLlRi7kxtNKEz9EYjvpev0QrUxVX5AqAKzcGO5srD9lsPU8AHkQrpbWZ
3K5FmpF0NtgDAgdq6AjwXmtsTIeMq3FIKIIIZVbFG4PPyuuxqL7DU8ErV5Q+cEVv
JNj4s2DM0UVFTlz9+sFOsaoLl3jXR3V+ZSM0U4SSlwqFH9jI5o20qrVnpLOASulO
WJlZvxJ9+8rmtohOopAVIzHsNGbITJBCr1aSd3fL00yWKGHxKWZruah3mFVmXE8Q
jJkmO3uDaGIn77jXIijktE9WuGNanMxxwUUNWCg+SqIi4QP++lGqMLxF5MSTECVl
meRG5wBayY++44cQd9b2ot3d707GWhHVW6J2pl7e52rFScLLzFMfMIZvnjr+QOg0
7papIgrq26GpuOQcOKeQzo1uy0y+0QMge5Zm+imp2MR6aDTq1rAUkB8MKVX0qF4r
vdiU4YiIJchwmCDqouRlT+MRdh/CR2yEBiUaXRUiwdntczfB4FU7QOo4tq2rFrIB
fVPJpgVoYyLnVVqVsNiIX1RC+vcsgE6jQTEHkCIwvza2LGtWc4K0iCZ3Z0Zqv4Xw
7yduHpJA7E0Wd/DVhgsghA9DFMIOiP0ZJvH58YIy98FxTDMTbUJ3XkNKULLLiHfe
9vmQ00wI6FD4d7MGXbEfMwNm8TvIG113tr9DCIvjG3mXfJZ5mSGO+NiTHhnfaXmV
LtP0kr/d/MRNlD9aGL01DJZhPDGSRQ3+Qzn/CCtOLs6GdzFKidEObFJOcGJHWrJ4
LCYkEXv8cuxQAg9tG12zwqN3qnj+jPo3yIX886QNotyyyekjdCWfPs4YH0mcM/e4
/0QXPQkIbxEJ8q7h8qhJlu4UppKRk/o8ljv0wgRA999y8NHsdOwK55m3AMlJf4Q4
0tXKAJYLTcRVsPF01x/LaDceOXUHIiu9dU0bogBJoN5pe3MQomztw6qgTlqPNQ7d
jnl0ABu26Kyk4UdtJ1bm8aC+70M39J/n8qXpkRyTg3w0ylfFyl72mlRirbVm5W3y
SZfBlq6we9vPFHWVcoMEakbeNEvq2oYtmRTcXy2Bk5zAxUA99yOooGQhvaOXLS01
dt/P3CkwPzbojl3Lom7OF+21SS9IRZlkzsWxzIuAP/neRrBpxibj8xK6AGtFIcjL
DU72ZF+1x8+FEZPg9RthH6G/lHIksiBlIXlYJZ1JkmGZ7Jpou2cEWtagOoG5w8ks
NhpjLsS15U1FrPNNcpEYYS5yGBGDUG3ijR82MYmrs/mpNBmt4s4u+NRFiGfyJwBE
BTGb9fUHH/qK+wSSQsKGfVSpLI1cQaOWV1yhwo4QtLTCFzzOPYFNYRZWKUlP3fmd
XZX4b/x/ztkCpQnhXl6ZbC7aq39cA/4nAGlTxQyXR5nDih+QLP8mxbL0TBQsVzWc
M8IoppfEmlS+Pa4YKVsPFRmE1Z52ywJkoFJbY0p9b15ngAO4mSbw0Woi4gFTuGdJ
dCYvmWue1us/d/o4ighGWFR/BGM0JDMnl0CjMpYhNyKwcYmeniFsC3BuO889O0ni
PcvXLKI7wagKMf0SqjyMk3iH9NeLaac1ipwJM23MgXeoATakmtPkhAADr5ygqPvM
knIhbiWdukh1buhRl7+EF9NBCJzQcJBP2fKru8QypopWR6yiAJSshcr0IE3+ID8p
iCJ4rj5nzFhd2rxMwkjnN3y1VzT/HMkzH+rE9kr4DcgJRobr0phKcTBB9LNzSans
Gr82KUNhyPJZ/KuqF7ZUHC1/FOFNJwaSnsnQ2ZH9njodclDtQfXVLxO/Hn/gv4I4
kuuWOrShfDJl32N8uau8mKvdEZMHNGMrNmowhdb3sBFXEyO1aNPCnVQdBF/cWrIs
SzQjrv+7orEGy2t+rYWR/9/kVgnoPTnC7UJP7wM+91CN1+Sm0aXWpL7gGmmSSKhb
SHiRI2/HDxy4fXtzyF9hW0576rD3EtFQTItmxm1y8iJzSkrHJuVydneBuSHvuBGf
b7sy/T7OZ/JfQa4SDgzBRiSIVtTGPvRTDyDygZN2ZTSXPBNsZMbLv7VpwaBuBFqO
koI0YUhNfKkG4SlNRRL5kodk8w5YAaFU51CMzQmk7GD3JWm1gGvI3v4+0idJ2Ygq
L301e4qUTZp54pgPrSKkgMGFShZ4FALuhaRm8iurII8D5ObyNgB3Q7+Gg1F5WxVi
io+NqbwuDJ9XuDTVZmjHxqjRvGPDOUNWYdc8CArIOtupZcMvU+1OuLDG3nCRDqFe
jvFfHQh71GS/ABVPylJomjzu8SS2NN4BkLt4ufQ8LIYTD6KUVvmWH2FQUJm8TOmH
jkVVdqp00MpZpC9YwADdE5THtnpf5VcAQCw+ceCcu7lEBGsNcwhfRDQjXXJt2uHj
3sGvvXaNVNX80mbGUK73yMQ+tS3uo7Zs9qURH4pBoOHen7PPhTtA+249WKlHQKhw
kDkOtNtPWoyi19m4V3jcH9rm3/gEGtaGHBD3k082KLjpzW14wraTIZIlH1ZbfNo9
8sP5dBDA2obP8pp1daQ6tpWnCOHf3rX2jHpQf7jUP5O3fBq12vyAwgYP3asQ9A0d
zhONQLBHIRH2B7d3PCeDDRJ5ZJ3cvKWHkTRr8yJVtjR58R4J0RwuRuowtCFCBndt
sA0fV0f1fwUWqRC935BycGqEpi5GC3X1pJ8D6uhfoTJRI2m8AQRTVZ5HW3MQGJhI
lp/UzpUhpRmoHQdUhKnvhWPQ9SPnXW3mgnQPe6MWEddLOr5w7fIQxwEnq7ivUT/U
xMbhYBRIlnyIk5CaZ1WMmsdugbR/pDWOzn0r8AcjiMZ1qWiXCPXUWoZSvmDB2zBo
zvPTwF2Om4t01hd0S2sYIsl676ThQv3QJgEyFLwLsz5JtyVN0rysig3RpefEEwen
r6rgZBZ41+VphBpdosn1etSyRqo0XH1F1eg/DvY/2LvFNmkQ/8vDdxsOScJf8vXE
v4cC1KBM8ktjthDJx9nqtdDNda7MbSoq8N6VSkWAiZv8f4WGAHsOmMwKqbYJaiIg
Ww4wwCHezA/CglQ+xvZCMCrhNk1Ai4aKd4YOQD6/6h9IrmeDL/4XvKKjCR0abJHw
rXvG5CAZfZWCAYSDUp+ywfG1Oo3hYKAe7qMEmipoAjnl6sTw/h1xAe9mBkGokm9s
wdLTkigNoBWm1qc2RGFuEOLXQgBLAE6EPZNy+h+K4Jt1+MbPXko2zeYGyjlOlMiq
PBXu3D0qsrUcbtJDC/Xkoe8pA3lWsZH1rgHkceOpRJLma2sVg53AaFc8RqEb+eON
kRHZ+1qqp8wCsYXKWNhCHkLtJI2rdU/K47QiavJil8vh6bpL633ybhSQ6NWlu2An
8RgobuzuhwqHh3Mzz88RXmwzaDVyikzT+mh0CBMAjFHt9pFyelK0nkcXB2lcPvNV
FA5N3apk8BrqmBPLQ/AtHNYxzJuNXl5oOt+K9qxtEomflqc4HMUodKO3ZaBnxbDO
NoW8UM8ioUlzmZK0s+6Nq+gkSmil+oNb07M69d9sKkOBNPue4pvi4BVzLkSrn8W0
19JUoOI0+OVRSVrKuglD7oXOuqOItX1w1wbv0d5ZN0ntAmdohQ+6XrlWSaErRmg0
PSSkVqMjFX7IJjJEfAAiQpINRw0Xf6ZQRDHHcQU9yJugZ7mjvpvZ3ZQDSKpSMrT7
hGCUahvgYvSI5d6uNm45rzrCsWmyGamZiwxAixnsDQ9PSDyaHHTeRIBNRMWRIB3Y
uJyNMuSjzipbu/n+7WQGZqvj8gmmaNI7myo199LNjlEVGK1dXuEMlYTPB+ACGAEy
ymfp44U0051Fm3aG3ROIf01SEzuN2CRXdW4kYFleA+ZBjCcYRGaCa9qzGYCNOGAi
R5bIFJDVO1HHWH9+x1ut25yz0QsxM4BM08+ZBBF9fNfR1BsSOaQinGVOJ9W8YliG
tb1deytMI+cpkmiBqgjGc4q0RPsNzvspG+PZl/oFQvZ1uRlyamyo0YnLCIWrHVvE
SRg0RcS+d5mkIvCIBj1LiOVZu9mevCHTp6I6DhXqoPj7RSqlU04G10Hu6TSzbUQ3
F9bHB0/4d34IJl0jG57FnauwgAExUu4rwDyTE4xmuuvqsIfQHqcQ0r6YRDmED4Ya
ov+QvipFi7BftnxI92wld7cG8aWjF1KyIvUnmkCZl/WZAm1uL9+QNsjH9YPzOGTX
jM7YHvnExDilxBEafGytsBp7E2ik/4VLLLfaghxwsw3W1dPL0lp4aCoLsPqOHNXI
2WJBgb0oc4gUFn6ugrIm2tGRuHf9EKNqrkYnU1ONFk9e056pFtaaGhPNHCWZP9EK
sG6hyQcVCSrbjeYxAqYD9zC0JO/zOKQur0DfkSWW1nwrNwEbRaV0y+36mE2ObBO8
0DMNf52BdavqJwBSb/o7D1Vtz+BhmAbp0/yyIjKeGPsIsKOGhQl6kZV0pWLFMuBd
v/reT9hfwcVIegVgaXpGJZi/gTYY8vErUdVCPLaFUdDzCu16ZKY8/AwtUQXK2I0C
q55m56O5ki0jqvFEAKqs4SsD/bcH+aupT81QqehvsOr1jnVMV+mOOXNQov0+/MAS
lcVJM8zNjsFCpkbs7PmQ1OCdX/PBL24VfaUaeW/SLs14npO5NqJ/xlB2NfXFGXJl
+gavEFAsmjAPACnOzB6Ro8g1Vd4ZaqWwvsTf9+oSEgFAG5MmApoEe7kdh3D+DoNW
Pidzh3p14MkA4czeb++xz5e1NEG9her2HBWuUgkvm6U88kgZrySRNM+ChebCQSGP
8iWW/zDpq7pYO6oD3K+rZ3nu1x0erQqnLhyvG/58ftPs65dB4ohOxJoxfWU6mM1s
DFElWokXRpJ90N8SI09Ba3MyVgzkVIwo2pjVyPaD9JM1fH3xRUm+3v6/GD5DgywP
bgJBd6bnVrEXnniqAnqnAQeVfDLUGKA3NnHD3EvbTgh2baEnN2JUZmVU2otehxOE
BZNbd2U3/Iy3xMVcZcj+9DuRnfjWmUzSjohHPtmMZUZpExjc5gF/cSVyCWuvg8/x
VjpVRlsIfV8bmnPAG2/XtE9070ARRy9Sge8b3VdXA2C2FFPxMgb5Ns9ABUAtXLhW
pKkEcX5/uWmm4JUhS1mpLWeXcMY5vz/t/DeoKLoDDkZ4IvgWV7dA/cUx6artxmP9
kYFuGX67p6ZomLW0q8HFBV682WxRUKshar1F+8vYEPsEVz2VGBznHibDE5A3MM+4
5DIlIAuSyZYrLAoRKLmv3MvZ2GuxYNugrEVfXlE5FOS9ILaWqJmilSCwpi2xiKQm
r97e/Jty4y/6hCdEJXU4u7Vby3+viNh6GHKwmQJ5bC9FfyvrnHUacDA3Sr6Byyez
D0dqpKFmqsGKc+A0dmLyT5hs6ywWTU3VTGAWNEwfkK2/XJHiL54uEuwZ+zHJQhTg
78QNKmhlc5udpEfJKiYDR5wqsQ8Gn76YdYXwV6XdeVEhOr9ukZCc7Ei9BaIPpmoZ
zv/vqwuEd8wiGsMkEe89E0aJI4RgKrg0zPWdSpbtXV0MdrnHlUv2x1DVUKCAu5RV
bBe8KzUuBwUh4nw4uPKY+E1jpoFd513O80d+dx7IVT2Bq9e096nBM4WFGzTL9XnU
ZMHdXDkNouDsLVTMA4soXg6LYHakzYP88wN2oC4prZD00+WjFjoH2BYnUfQOhDOb
MqvI71u8DbGDf31KH6rTg5cNEgfexxnKjHOiCvHqAXrrZMPJ7C35cpp9yewJVFR0
ruUsfZG14y+/sBb2rjOCL+QIGXgBFa6PKcHIiqGUdV4vzEyWex65agKi3x442bnW
m0uKsTgD81yM3zvPQ1IRPcJCbPEYqJsPy3heGC3HMfu5w6RLC/SVuWbEoZSbTou6
ha2jpauz7piFltSlGpHRrSjraPiLF7daEOGO6qBVoTTqTgcBrI/D4R423ur9gOGP
L9lXmbIHoqW9GJDwIqICxAbHjCC23sx2Rf7+rNMW/nWKTMcONRBCXbpth9W83ZeL
PyvC8NH7FdPLKxSJUqc+8aMN2CC/rc7bDza/HuKFEeejpJWsWzfmIMlA0LprgQVc
11KYo7J6gjM+oJh4Z4uDhfRhaEILVWBrdlzHtVdc0INEpOw0YSVDFC6IzuOloAFL
8LXtZOjWYR5TRnkL4kGbFPShsR1FSSGfSs+lGe/iPU7cdU5ovpFV/NfPG4jixMIl
kpOEehULSQXvj6tmPPtN62AijmClGG+6KjVTAsijnQ9y/NBRooUcYS1cmGm0xysA
WRxeWBu1WdYGQxpBgTB3/qf+n8OTkJYFrKBfZALHpLMkqv9JilTXUkI8IXpBup0l
QSXT4VNxsxsXq9kkt7GqN8SdCGFWPPKdOOMfXG97/jZZOmMMiCW02YSJnIaAj64c
CQovgP9GRaRI7GDlyPA2qtOLq2HLqUpr5iZSLUc1KZuWg1CURfIxnHn7ixfD2/uO
Q8Rr4A6r0gn7JiZp0deHSjD2J7HVBxtGt6YfOXxyC/OjaxZynvnjsrRGe5CVLZ57
vlcaYIIQGT6gkO5F0v3IgXp/8fTD9x7Tr/YSKvl+F3VHBWTuFrwcVhGKGF2P1xeW
7uz1xiyiqk05jc14kzZtC6PuHYm5BMI3HdL2P4Q78OEOCyRZXcFBG9ZfRbORM8uF
a+OiDUn9slR6C2Q7bg6TCRWrmV/0TiBX0fuDcDm6YJdZUbqcZ+9OlkGQTy5tGJoK
a5KgoHpKaLWHriQsGSfrZCJIHG75wKw8n2JByTfRWKu9c6GGrYzf9C4FHK6bGX2x
omQHv871M19zhEWfYeEzpUAAWyRrnPvO+og7/BHxRXpqotu/tsDHSJ/+5/nDdk8C
12lhdSq7xMRzGvs6Aey9+cpLStmaZwzXoBeP/JDtwBEZr/tcZHAJomu+XzHCQDhf
hmrqENmQKqQSUsZ/zfdULaAjyjsnfoerxiAAzRDCJYfwqfzybhijkE6HZ0+6YuKS
NpAb0QTuGcQe3cCaqjszKbac5fPt1FKRRUbxhhW2NxwBIJZtkF+TSVkxQYN5H0pI
XTmF1Pkgq1mEsO4LQH3dwt3ImkmK0q2o+TpNI7LDuSp1LbWGu5nmgQ/3BU4+gZLB
81hLtL2174p6dHtBCyuQ0qUP4+DAdZP1nyF6IsEUbR7IkOudXmE/RtDDy3dXt9Cs
tUFLt+KTt+m98YnDtU2YQP7VNz4TOFIjF7kZ59rkKASup/ceHBl+oGfhXWAxeJhO
0IR4rHlYi9ZkxeRhs2sKVHsy3HrPvqB3N/Y44aiGcmBwQCZ/fm735fVj+115YsJo
y0fliI+EZCgIyXwflhhU2aQTskVVq3RsGsyEuDhW1LxU6bwAsUIuwqy6G5yRE2kS
yaI5vUhtOBRxZiFJHwhgYhBaQirl4pGb7GW9ym6/ziOFM3vc08vjpkAD5QwRtTs3
IgMwbeQTt5NKkvzb/cQ3xHX+fDlQDTa4AYKkjyK3J0nl7ZeAtvDkprzVD/CBVqOw
IniG8Klka+bLcCfgX9BV7te8gYfWZLT7V0jWnsCNxF4Fh4BUCsagRsL1bLTnxzZc
ryovey8FmLGlEngCJGHTxWlvjPAJwFIpST1XbGmgNW55Zxw2jdOrtmFE2pnfFv6c
zHX5F0h3IB+E/6tBK9KCafF23ZtC+6+jPlCm69vK4tfSNktcrJt3qmrT/zEGOY9q
K6xn0Xo5T0nDrKjmMy4ZEfCOI34SwdPt7H8mfSk+1gXdIz1cDWGw+TrhOREysvN4
CPdM68FK9lXSmcLE80bGIYOQairhKGMbw9d49OtVVVOu66Vq/aBxwjaiku6xoukb
NZt+bTfPpNCm3paLPq9Gbacr0RjBdsdpoKf+lXss4ki4gUY3z3ox5ngwT4DP6omW
bnrPNGwi93RZvfeTmDmGtJ2J7YYMeHNSDT88ziN2MpCKw0dJsLJ35TbHw0Iex7Eu
6HxduVqJEEtZBCE5GZQzDpUuKuhZS+qi11KBD4wBCuADebxWSUP4chR2ABm1qGlo
fRHgfhInhO3MD5IsJOf4Dd8CiVWL8sXgbAm3uWYIYxajFtsxXjYop9hp3uwNSPJn
l3xdKOGrdFM0uPjGjSskc4u6DmWdKZE54RuFY0QfVa1yUX6UlSmd+MRvBcOXVInl
dxjm/EwNr+cn9+ZWVhvIMtPJUcj1H8zRzSgbvijf0VOz04se9MmSspmqbipFVvta
qV/L+39K1y0iWrH6Mhjnk/mWp15Ql3vBr1G3Z5J9RzbETHhK/8q4bERPeQ7PEGnd
1xLUIVh06X20ScRyH18Ez1+dN1FqoDMij5c5ZANKotbpK27FNa0bjUDibe954iFF
tPhhhHSBYAmJUPfCMtKoH37PEbUf6ov7lqw0qBB7qxuk+ai/5r8PUeme/Ag8xR7f
CE4SiaelstH0jN23Qs4QL0QSdjEGjiNh1wQaMLqFBZg9y0PrlrFQzyrqmobvjRDn
y+j8RsyJ4GqFXmqVtcmEIFTLtEPWzD+JCDOc4an9esVwfrI0O6piAYkRITY3Y7C9
qZzfGNs7Rvghl94qZxABnhuZfUmkaBhKuGa9ZLi+4PgkHy2g4MINuxXeBKfY+f3V
IwR6viOeaZ8VZcez3FtcN6LTVDrs+75zGcmV0jENP4PXF/SLSJr3VxUCBdUeDA8E
t6PqfS7xNaTD5aTPokJ95oVvtWtRZ8TAd4uKpQFmYDmoZua+jFSytcf1A//0B4b/
QEKq8u7fhCSGF5AdnsHBZ75DdY67WymV/CUKQ0TtfwF3DxzQTxE+igsrojiD6QJR
cD40R+iBaWbtZPK8iHMjURy61+I0VHYnZ9ozmxFoYaIDZnGRXJR3GQ3sgRG0Ds8u
5LSoHXzfOTM9KVkg5BNDYemG07GVIinmU/CE5qksWnLiUPAIFETqPoGKHsUmfcll
+lv/OiRcUP4PQZ4eK5DcyA66o59aEqsHG4zKbL4NEGnMBZhNXFRvcypJlZtnRuVe
xNQ/DJX+lmGZSm/mlI4ZUvRjxvFiKxTOdl12Gd03nRg6vnKJ/7QqYrymBIjp4j4h
D28g+EEw5h7bJUdLo8gdJiwbMSZuOVfeNESSf/DHJXwFoyr5KeLlsBd7GIKyniJ7
CH7jG7PoIfRvrHB2Wkdfhh1O7BfFNpA0S65xYi29rIV2YHP0pE1lfYpDIo+ZOA85
LHAsC5pXtRWCTAfMNkxhC2fcc0i9V3MLEFKF8OChu0bHlkJyrw7cgOdPKzH8DJ/p
u6gKh1DyJoAvWR02lKFzQwv5bWSUJ6mjm3Kuuc80fH6/vc98TlvOXjRsxPrWG3Hh
PElf5/a9cVZvz02ii3g+rQ1iQ5mYUPBZwFOOJwOvtLBvC3RhIYSQUOTmkVNT4vUp
N3/mYBehSO2H94kBHaRIUUC2mWA3yI6m90mL5dKcMyv6MLzqTeXA8Rr+itwCAM1j
x2MOumvIbY8NUIM6nq4bw1ElNyPtv0XzLH5yPECHYUlxpyXqfsL1cUpSyIybvgNw
qBrWK7VSdukHZyQihJ6Q+7YzvERKVqc2MSzJqLv4+Z54mMgLlj+VynR0c2c9pxf9
nGjP3uzkjFMixUJiM7PMMoEC7Y3OZYDj+a1edZqL/fEzDX7f58bxLUj+UUSVaf/+
jRhY+ghoXIivgY+Lw0i3DhfpqEC2/QjRvx4P25s0sDpf1T3pPcQyDRwTz5RYx+nN
dsZvb5aWyJcnOvcZ1aHyA3fODdMQ3dit1ufy9rhBpNSoI2PvQ68Chl0BCTmgQx5/
SZ8Zi9L/KBuR+CcqB5xWPMd1qnzhYoWkLcqgE1R5mIAMroTHsMRZtaq/mT2BTiTI
x4KK1wDxSaRlguY9pgvzycdomdrmdNR/MzYknAo4uNuXfOibFP1piNgtq6BH1UJM
NNau0pGLQhxmyuV9Fn3/rUzXbVzE4xk+FM+h7CyEbpHcQtLaRf3dNcdmn84uoG1O
bTCOGBBZ1GqGX7oEGt9hjuNnsqT5r2qS2ZiaHFab9gyxrn24k/INCI5gCEDc3wCF
7LqXlsaK52pMCcYAvci5I+aArHwQ0JEf6qeIiH2dCcJdyT8FXKbYBpmEDcVYm0Af
3Zyy1UWeqb2pPISRLEGt24QAN19vrKVWantTFafZLzoOitGoYCio4Lno9YtrfQDB
shUF00ukPSlQqn3YEFDdHEkrai2s63ZIZmR6aUaZoIHfumZ9nOWrXBsUxNeyY+5p
G3Iz/bdgkdktsAHFCwYYTGNDPnqGGJu0ojq7e/EILXn9UFmrIMujHW6VH3X2lAc9
xRiUG+qI/GQPDUhdqmLfWwSnZA5iP/rz02O/AezD0ZksPJA0sVN7+eh3a1aHWwnu
doEX3TIojmrXvdTWnxVkgQ6yjgg+/p4vaHtz5Ur0amDvP/Z0QrJ5AscPCqe9ZQA4
Ot3oyPfuJA5qX3OV3VeymoijmCe2k1xgwgTReawAsnMj04KY3OfWYoW7LPfeCVLX
THKViPmwxczAGdY61RKBbthu6JXul5V7g9rMmXn1qmSFULENy6n2NiylYxS/X9bf
oJHrJ68jT5y557kEsPPwNgNp94j1vruqwjJHZFkqQ6ZnXsUdhB4qidGm3G6Y6tsm
SO481/FtfM5Q8MZEto0QW0I0aUYjYRTn9Qs2MU0UUZ2leDG1N+S22+6i4NgOnLZO
MXdrW0KM+lOG7icYY6wZBTYQPaS0elOIPiXpzyvTzzesxtnL+oM4CPnBz2fn0NhL
PRbtZRQFRIk2dNcYecnRpXqGJf4FpYOvJa5e9yzl1CSPSsDcYGL8XCeyghsjXprh
GAnqZU2Y/bGlszZ6c93gG2XR3nrYmm/DClWbSXwD2nUEMf7Q/G+VkHSdOBsXm6nm
ihKz0a1QbbjdJKkdWU5e8OLpPZhZJq3O/+PgQ/CzqW7wn/pZxaxRTYx29ijR58JY
uMPIt5EZwqScbJf64yK4UVDjCk2HnlzGq3bgkHtx0m80HHMt2dFHcK2arjxN5R+H
+hR4iS1L8vgX7kZ2DsOGuDZDeS8peGxKrmYd+JhKukmswbBwm7dDPjZsxygZ/paa
PnzKQR5QsoGvqhUFdbKwmsd0j1Us7qoOC85TiJJtdI/kvqp4K+uW0gQQfAQroxYq
tvNSeBoKvJ97IBjlMWbHIKLUuCKtI6I3nGqeVsU1X9QPwcu16xeEGohfZqqrvSCu
ihCg0mqxzpsp60jITGjpEN/05x/nZWWTwtDrXLNgrnI9kzZ4COidmP1AJdl4yfSx
5IvQFxpH3CpBCdPvW7OfRh9K9zpuSTxzR8sRmZGd7XDkETMdV7RB8zhCNq2+G9q8
9Db0X92wbpSxIbgm8fA3S6avCSFn8VZOnKD6e3fyD7Apu13MP15wUUqcB5O7Tut8
DuFa5uWnNUjWVYo4gMFlNWReGvOrxYolB+2I8CKJyfz+WnXqd3VfF8mR/uEW+Ebl
ackENawEFneOT/yWvyBnKKueEHC9R+UGUOtJMw8YfU9mO3ZLd4t2zkNf0Iy8xa16
IebhdEkYGxD/wgde08o37tsqxY7kIgwMaSN7W4bYoGIax8gdcczKUtxMa0Ujd8tA
ieiL1Jv1GoFuKXeFgRAcaLvxtVl7wn8gPoo9wGY/KP9nSDEdC1wzpm2dJ8xzXp/b
3Hj/G2L2mRuu2CbIM4qUMZ8XsRYufIUBjnmApJvsFeQxhRThKD+XCCvYVDDeUhSp
I2Kzdifo2+T0VtMEkSsCOuSzQVWBoEIWY8DRVBYRVRuQi4pN9eBnHU0t/41x+Opn
Rs5NMRWc68yqNKEnQdjjwvERSNQZjgVpsGh56PBNpmuFI/H5IeOVVNieeN1bNsNi
loFz4PZYF6wN0cUfALUIjcfY1icfsRcW3e4b9EOcQcgP0+ZG2ke2jsDdrj51FQSh
yurIrEOZaUhrP7cmW2o5TVTsVafWF0CZvnAOl4RvsfctNyJU0GD+HZzKZnxLOmOR
b5akUw0Or6l7CahjhikB0HiHuf0f5rRTEN8iuFVeBAHOYn5TOpXC3ggw4STWniYd
mBImReAa6AzaQmW5TCXLfvRVNk1jza0byKmblfqw8iz/GpI2VYDk20za5895I7Q0
2HsQJAaDkovIELDsO+OVaTaJh+lx/LnKaQnlm01CzVocs0lzzYiptA+U7n9aUSY3
MZv63w+oiUnC+97WfZJHdXFgPrH1Equb3dcP+DPQbUmvGGOm8XKHvNHfv9/5+Ab4
egUZZ2v/v1sUKvJFmQVkb9/j6n9D0+2jkxLIfURxB3L04QHp2o1RrYfQ8mVIyxK9
uTUw4ItoL9BnSmKlmi9LaVVFUqh22pOB+Ka2UCmrLWK6O8aXM1UbeLvYPOFBbczd
Sad3GoSqf0l7CTIwXFy/924ygHGJ5dfYjYmiajlIKD6/dFahVrTG0urS+eNFs+ra
OrFHFw/zgQbPhv4tnE8lBfhkdtfzYLDon6Tz6A7JqkoC+BdealBQ2k/g0qnlRz9i
IH93aOOy5dQ0G2ywhSWfpIWmHRV6saxMTNZhpwGa6a8INcifaOv0qEMwwaF5yCMr
WQXNjxNd4L1ox8KtYroJTeMTaJnOWKP4WKZRZnRQBH8tdXteGajfU6+rMzW7wr5h
zjwbPioOSdm2J0744S4JB3asvv3pkHTdVy86q8BZkcL1onnx3QBFYc4vk13Kl1tq
PxLSpU5SAQ7V6PTziYJVdkKRaslSkiz9KpGUAVfQyvigBbEh8vwWVGfNK95wkQot
zHs2p72vJdsR/qv5dV3SE2yQ2rHeXxF98k8RKT7cyZTLZF7+gXYAIS7p8hLAAVQ/
tTdZpWkH2ZZnLAKIdKw9xOc7O8EsbH5761JYZin+C/HFEu615D3IFH/mR5729GDE
Vc2GDtPcFGIHcNWgBnLup4o0nPZu8UXV+8yDzBUcTGllGU8msAtYaxvGwh0Ca6xw
6gsuo/eewJ2EGQJHaA9l+YU5L4AlVoUXoUCJCCbjM7If42wbX7kmIIFeC8puCnC8
2bY/FoXHlFVCtLT8wXlbmdW1ivI89s+5NEHbw/anlkCOlJGFeNGmIyYVY/iuj8w9
7VK4d0BtrSFTgqMHnXlPNtWME38T9q4bgh1bEp8Jx7r3Noc4wWoghT87tdt6RvcZ
BxfoQtefg4iebTPVM2rFqoHmoo/P0H6VUO3owZSX34lioyAnYnM3t4JriVdJIMnb
2J9xtlqh8P1LxaoV0O8xRiAuA6k6ulJadzkDyDSXRJ9YVTFOfnIZerpDMgaN4coe
GDQWtcbTUZ8rH9AY/wKeyspydEZGkznXjYXoR4YJBRXpL8T3vQnQMpTIeq1K1tpd
19EI+fGmiI3F9NgnlHq3Xwr9UGHjw+qZSMWxR2rT17Fyqse8j2NZljal3BxXQV8A
hrDK9MtGAn3MVfTqko8gtWQVawwErVUt0zDUVd0bxBCCk8QWyLAOWq/WU6CSSfGA
6L8LioLrXAw958cJ+rD4RDfVcATZaY5RhIcDn8V1f2kLQ6kVuHI9uwqt+HxrPz1g
e2A7GA7AZX74u+XVOJCserDIPLYCv/FqJ47tGmvsEqGkWEhJOmEYpYY/Dek1yK+a
bX3mih33GEomyED4BDfYH6/92i/sbx70WOA8aQ6Hnx/neVAEa00gdx9aLFuC7n9h
LwDiAcWDYJKMVCjWrFWm5buwNhbkOn/wLNG0JUQh3ga59s67WAe5nEGfbV24IrmF
GAgTSLTMSO6H6kzTCkU/EEe3eRlqFq8ZaVHYo9n4TPVBpla5jCmNHTmoyLba7bdu
JR/3l7aqGD+SsxO0k8hbw0SxiINbQ49Bmn7eRW1/FjMtmP26SEn3R4QRSzwxbbJ5
9UL0bZfiqBOKd31+ZPXYHL0OHruXFh8y8u+U5y0/+SCqNFkDNNhH1oNSp+5gLxaz
wi7k1U6t5t6zMg9o9azA3Hp4lN6gcfxqoT4RRpXu8mPpO7WHC/+ZHYyJvkmzwG3Y
DfmDYt2xaKUEf7B8eTTMj/H6J0QWj15/SDE6hQvnP5hP2kVCR7yN6xcO/MT23tAS
grG4+qDSqySRnqBxFjWLQmqNbaNYXr1Xy7dsrUqCr/sf1OmhOYB4P8LZc7T2nbiH
sG6n4HVKNXbyQ3z60wNwCyWIopM12NhMENNb2yZSiJf4id+g8EpQLr7QeDL33fr5
1Rgwgpw97EZZhvNjGFxz/C7KNLihKKCAiH1pzPyDx+rvyxv4/bdEIJh2YJ9LOV5i
lGBK5uCBvgsk8lE2gD0baj8/SFqWpelCMzZmBfqg9shFGu/il4Hnlkyq5fkJhTIB
pL4/3I9Ij1jEfMjy8um28vbo3Zo/5vRDDZQ2eq44SUV3uKOmTydjVWIrDxTR+qCU
bE3CCNv8L4k2CWSG6v7Nr7+12NZWQZeWGaeK1a7bIgEJsB+QYTlRWIh3iqd4ZdZN
/rkBo0Za7T/rTRDVmqks7E/KGAeLjfniymLCYlF8pu47t+1YNMnBB/jkL8WHbxjf
UDF40ML/XZocYzdHhcZQ7MPSLLJdTmicU/wPWIHB4tYBGyHJ9Wk8VVE6LML3qXGB
aTkHTa648wWadzSZjxeRHQFrbsDS7HwKcA69pKtkPuH8sBKcgiRDOLpwtAyTtPf9
2hqimp+t2R68XJDfBEvo2kc/ikuMX8WGhqIcbdhVDOFh4+O7mNC/doMCAQWVEQ24
IejS2lZllr4px96E9dbiYTY3Ojc9DqK/Q7Dt0V8GmgR2x3mhkl2Dffz5PuCl25XM
faAFnca0rJNM5nsNDAaAlDDMKYpXVI/izfbhw04vpgNFo1o4dFT4iY8iLbhvRgnc
ZD1IDoEuxUpzZZTJnOnx93Lzp3uN4pj4jz6b1BiR3OlzQG8StfX4tcIPUkZXgxDR
eykgfHfu35Qe8DZ4+u1/Fhm+n6ZVZeX16Z3f0UDzuMaB54dFzG/AUhRjN9/WHQu9
ohmVS5+C6igcfdqoAazhkdB+jeO6DMN0Cp3iep1tAaotM6WmzRHGtDTbKCE6dYPO
ZOMxwkf5vNYoXK8rLyGFUlr8/LFLOIweZjAoQUoqfwky3KeT1x7QPuWcvV2QdzkP
ggBKUQFxH89sS9Iks0ZRCy2MzgI8ITJjyrSZgEXA8H1lDsGYMGOBCxtoQvdCIhqK
roKMy5J5QWNW4KP9G7p37EuLJW+WMcoeP35erYmdwIu9Yx78Jc/tD7vnQD4t94cf
QK9pOSJBM4Az7ohWhlz0Vr2a+3Tn02R5pjfYfjj5OM7xEHo9WA5XgBsFBfI6xpaI
hUay/jbED9oisXS8puwn9D4Ig39myrgXhqRipRShgmppDoCUjCKXekQpeqOmWci6
hwMzHjAsfBpke2Kkhz2ixxuu6xNqOfnntc8EnT+ZzGDTfXlwmA03iRW7qNfBvj35
2pw/A9XPXptRD2TDkzkgX9fI8rJ9b0aAmoDujaIweFglHnb2tFScUnMfHqX8pNpZ
aKZ0YHp/SiI062WS+psicRYVJqYxTHrachcd8gGSaQXmKONz82qXzdeDiWv9xiPd
lFip4+mP2otNzftZ2evB22Er+523BUJYp9VEr+rRJZ/LTckIsxLV8YZMdh6M3oh4
HahgrlCmI+Hav0iE/0rF/tWd+9GGKLb3nDwwED/PRMEr1la2ow9mjYM7ezn5j12X
yoUcNmzz7dQuDx1SZdS82P6/Oz8/S+7ijhTKemHz32baFDiVN8Ao4vP8Qn/xYujx
aP8wlmlYiAwzOcgwHukS/u+dZtopg6iaCmsFej5rFm7RW6lFfB3/zdKjt/Rzm7BW
omA9wYtA30b2JtIzZM0dKMlTLyq5qXFk6IR/8ekDFR+FdxU0gMkDp6YUtB1xbM6m
ajrXHVsup0nRLtDC5v4MKiTIJBuSsEoPbUqa4h6Q0hgF+nAPAzKvaG2N8vVIH1KW
9Y+D4DKg9Zbvw/BcA1mEPur4xijZWbJAjcqntG9SnBBFvL6QqmEEdF+Qqoxn3HMA
cbiGL3WOULFitbQ88rV2aQOCJUtuaduq4/vg2YMtI1kFJaeURY/K5Sa7ATGHzpHc
lqKMdDu/yi/CSewbi03abSPfYanxNMtQU+ASFREMTLpclfnYEOVz+yPhInN7+a34
CAFe9xsJxsHqImpiCLxj5UIOC3loPDWBlUJ59GJ5ewO0AeZgCvMOSc0Nn2pSfIIV
GVfH5Xe2nN+j5B3oowmR+RhsgBrPdPC4W61RJAAUG5c7cAPAlb4LyAVeXKuOttiN
PSv3ZDUuTMC75MKwNTwxUXlA9LNINpKilFSBKRJ/VTCGBbRFES0TAhJcvlqHMu5O
naG/dZJrY+qaj2HSNsWbv65569ICU8bncT2DJSld1ZRuMA0fWcfQdpJ1xQZMyN24
JWhwBTMOtjSO89XW5HWKxTzTaecEi294bmDtJ3PM+FngrAwDC3xCLrqTnkpHf5EL
W07ZFO4zgERkq9LWSioR4fKlNoBZEi38mxruJQuYb9jgQQ0guYP93hNluegyc3W2
FitQnCrdU6+4sRQEHIBgcA3+18ddcsrjSD3mzLPim5MZXD61X8ZX3jESDOm/Bs5D
T446//dboLBSkeliL1xYv5Sv3+LefoYVlVWM28/IfHlA4OXUcludMCavD1PasVWq
DcKq6BeWvx4sVs4Q7sscFX+bNccu5MOhuWeUsuDtOyGHlNBxBaJ9ouROX7jPVcHS
gpiupnRxPB0nSORI7NtKBzA9xzYZZOGgn/8adiXHF9hBcjruX5y5VEajaGGfmcAM
Uxj9xpRbnsc//jlAm/+gihG10v1W+P79bxAKPcRM7q8kXKDOMeAcvG5UmQlz0Lvr
MwLfiVTlv8bqwoZSIMN46RHUk1/ewkLuZg1SUrW0+OPvQ7yDiGDjOlpkiYAfiE0p
V9YWC92oTxJOfmBoOLpv4MBTOxrgO7NdgL1oYzGSyhtBgmkfoK5CeD+sZUvtfg96
fRD3KbLrFZPcNbl4iWd9RKpgEa5T67eNMHvVkSiVfzDOhLfMthZvCUjqws20BYtM
cfsvdVl86zCB8l2QFN0Gqv09EQOM6rA+QjUaMEf+fB6cFBmm0q1Kgr881hqE9arR
67Eh40GcFlYLuEGplnBsf54P0CtHu0QnejIwRZvmU7FOe6Xy85yvT3xjSfjKEWMV
bMnyzVgBxcB3HS2len6UDx3rO07TToGCpdw2Abf4lEO1mm1yFuqTv31iKjP8w61a
+SwxdmDYUDcd0KaW8c1XvHoUTSJwoG83thMkWYSlUdMbhL+v+axxD6etevckdalC
ZwLtYx8LIKqy+2YvczmFT98rev0VdAlr77aMPGUsTcDVkURXmt0z7zkPHWUbUAk3
jkp/lgc0nN/4YcCLrQ58366dzoJpG1PLJYrZR83BGTQK9w7fTlrAr4Ybgl9QL0ii
CtGMyv0mmnXSbnaKWe7115Dl/89ahKJR9+Tuu6CCLD5to4E0qF0DmgsB1mCCUPGT
oITRJZDOAazGDNmMa3ZxOg0JgBpXfAH5a1QcXY35vVH9IqQL8s369RHjcYRGlZJj
NX0Srqea9aUHzD8kwU1sSsgnfy5QFQ8s9g4Xt5ULglrhL6RfNyAGvwUuw+bVjvNg
CzjU2hC4dNlHCXg1d916ocWIUde6UXXH1jXLzbPARWIISEvmWNjJ+8CKUfv9+Fl0
vVo4GB2sTIJ+WdFhC5G/erSscttPqfakNXVlpvf+bdKThijl2Z6+BfBWOB+s1jqR
xuOF28vVggv9P1UFTQ1X3TV5daH3aHNjIdtXDnVmpZ4+K6yE2zh6x7uYDQQfa3fO
G5hyWPRRoNJkXF1TULLSKmZ3SiQ2mg1eFddNH8OrKR4sxGt2pHtC3PYxQA2PWCsW
HMnSJ307pUJ1n6wuUUTkmS3l2FWniZ3tF/WTV0XjLdBNQjmZ5XOW1QLzkKWtp3tr
nna1zJzhuX+FPqFnefEsBkI4as/VCvcJKcAYBq8eweegpv1jGSFbn1FNnVI+oOLc
1dju2M9i8lfSoX6aWTrq7Zd4dlMiw1RJ4HGf7d8Pawq79UPLXPl0yZQQPYZllJEs
g5kll7NG2hCTnK/ibS5ndfMErOIGNm1MndT4tKD4DtBtrvyXVwGWHHbbqR08t8o3
MCPwhJAl8T/j/7aEbLdHqR3MvlfTLJ+d+6Fs89pP4mzZYzni8TKMCnfdcE0xwq/u
F/81x/7Un39PdptWEjODLjjDuoun47yz5gksXkK1wTlm9J+8Im5ECriwKSwMmaSc
7BWwRsup+rxwwr6rl1VsOvTCdHJheh4D1NSEBvzl3kKClbj3UchtBJgEHRBeZxSz
k67J2KnCK9t+h17n0Sg1HXC0n+vUByJZsYa7RmMsU1cRTvfDMveqdG/zGFZTcNGX
DbndlDdSNW0io8AokELCluvdtAYCwfY3MTox0tkaceh7ibZUGvkKtfx8WgsVlFlG
4Km26BIkskpFoJD81CrFDrXdy1vjr6+8C4jwrO/Qa0wSN4Vc8NS4y7mEQ02ZawUQ
RX2fADC1CHaMX8e5NAeXG1eq0v+jUv8fR0P9lfV6fSxcZq41rNki9FBEfLMWlIYu
qnz2//6pa0VRd/3C7jhNTgtSXJP24XZLHT4uZ2RfvB7pi322CAkXUIpVHxThQ+Oy
7QsQM+BEWMEb7cGXkb6GoBhyeneoUEyADFQz2pqS6HQbtLQxRS5K7rs3XNq006GQ
zOKwAYEmAvoE5a9nzEuPjNRA3dPRBUEphPpYRW7DJzH92R+Fce7HcNuEV4sziKhQ
Aw00nWK9qw8bxzz1NcLizesjtELhWhk6DtD3hwEr/OcB9xurTDfc4TwrVcxvooFE
9pqXiZT7fXJQMvKGD4Q823LE5mCRgE7IptY1cdIjvYdCKTeIPBPrdzwC3FKLf5k/
wY8AoIMBwu1vTCR5qfnMRnGXS04AzycomW/ylZF1NNL5UfJ8T1xdSFgHoQqrn9Wp
S1gBGss6pnrMRtfS3YEKor3GhPirVXTqbQmQ14JmBFBvimKPfSCcq64aqdL5oOdd
fiRp0O8yE3KuxUlj4JzXO6IFaDVVv7AhhKRABcx0lDGVJjRULJyRPmiXMu4RTg/A
Aqu/q8sdy3OUVhPArdwQl4yDLWmuKiZx5P6Wu2mv6770A+oHeFfr9ugk2JWTIWGR
BRlrgzcqkjnryQmpGjGxwUeuKln8khxqAln+rsF0vvXxVwbsAlS7DteD2FRjKZtv
40sI71DMDbrFi1KYg+1REfnCnYK4/l9htMQdwRM0pqj/9dnAgQSWCTg94Allr5GR
jqx4CuxX9kiRGnqAuy1UHAXCelQIwPA3UG8bamYiWOf4A12oMS7reENuXcNWmi+a
PbXkrfWXxrf+OgR4L+12RgLzRbn2oCsYxBO74wbpOCC2gUSrnrTeJk37nLUQHAaV
O/2htNOJIwuMPW25vDqQTkUKGuU7OxqwsAOwIZh3sz6l4nfTv2PqXmn4aZ2XF0X8
nO/sOUHO3OJ1m3mdfTX+ECEQdqe833PgJKc6BY07OotauP0AGSbYP/syHbKPrLPI
PFltArtgjI3lVKYO0T0e0UnsxVQmJqZFXmOAssUK1i/NrCkPKEyxIC8yyJGM7v0p
uJmKS/c0b8WRhO6CvW3EK+mft0k5NWrcIuFSe/DkiuJ3+p/w1J8ymoZncYNYPr76
WyDjgOHH4Alq/Q8x86iClUOv+PcRQ94HKVne99Htm+ymTmoOjauwoNMz00GpXrQj
DzAwCvOQVSN7A7aCtQFuIpbcPJb6fVCkLvxhQQXYx+dMmHDmAKATsvc5xcF3cLEN
uwcfeq0JDiDvOLskke8Hw70YjrzUdnrF1L75qmvvEw6w2iJ5BUjVMpEuiKzp3Xi0
trigz1wiT4EZJfMpqGqCg6ywOf3l2rqYKFfSSiM9VQJl2/clbAD6KOTOiEkDeWgb
81M2T0xfUvMJut66YBiTGNfwcRNfMuYKAofNTZRH1pJKkI4ziou41XOm5Gf5wsbW
nIkFsrlfHJZZGFdAZV4EF0xuzPsKAfGfDg21DHhKLlKCiT4cce3X/cd/LujrKdgF
/lqRNJUsGL+cvp+TEShgsujTTRigZ3sn6210dOkvsRSfU6fq8GS7g92QSP2Min5f
9VhM39DwKF85+H/KV0uHTDBFPyfAZE2dIJZkdMKRcQ+QVjDzU0Zdmfcn4QxAEfQ5
U4KTdbAlCd2vkbunhExHiil1W2Sp1pyhocHOdC74ZK5z/TRQNZzq1r/7KfsJmN0C
ZAcgD+NS97WmqJDwoM4sXQiNu4I9q0oLPDSHuDx2uE006Dpr56gD7e7UL6kwo7IY
kD6aE8EPlstvuBoNxQRMzpYIjq4DncS0D8nFSo0vjEOBD+eDOJkaXsq15pyUdlZo
TOtH7zHkuspKsquRpHAt7l4Z6prNIhydPdrx8/f5oOXfPlXqwikHJd79NUjAMRMI
3qtQSpA1RrkmUS8nVmDqQe+ZsgJYaF+Aclp8SLLUu9eeb+HE8+tqp9Nyf7Fr974l
4HVexcgVtYBDE2bE5qVkdSE+gi7oBBGeerJlzEOJR0d+ryDVwFRhe8LEgWCnOee2
hMj80cuzkjGRlQ2ujkW2cMFP17em6qNDDVNqOCmksxFf+UIQLHecKG281o/Ce009
sNBO+ZbpgTB/mxI3mIeDYZnhESqf4Ap4fOlSv4If8/fWkQ2QjYNU8uksLXM3MUS4
+rsIa8ZeHzLWoPznAtxjGpFd6NU/LB9p7nlUkojFAkdYiq+G6XP0l1/+lKefEEKh
4wZ6Uf6Tob8h1clrhKaCYDkjpfA3caU4LKh8reFZnniz2S7Q65b86TicuXN+ofu5
TpgGy3xvly9SXi7gfCUx7pRnHdx6ZcYk7f70MtSf8YfjMjMJxoahg2rxpok583my
+YdMDimOaRo7aufq1a38vb/HeOIkXso/xxVjT8LpmUzhJy0aM38IHOoxm9tMex3M
1DicaHxWgopAh7lZ6TtgiTJhiwJbiADJjrqo3ZY6VuJCdCUgqSona964M/hFrGDS
KDmHRiVdSzyLuRy+c1HF7e/Af1mowhgHVKFxBoLAH36XKbOqkFOFavJoh2iup0qf
KxAl9jB5eCd1UcRZJSc3ccydyn728Cr/fPqxNJytNKnlJ8jP+ho5YXubvNuxVDBc
9mw+1yCmGJq78rtAifB/Kq+3IWOv7Z3usTvfzTRdhfthGzFzLPmlofa3o5MOe7Md
5orbXokX81oIsXQSH1gxtza5oMTLEEPn8sLRG8RQeM/PYVEyLPv5Jebj+nqvcN/H
PQ1FGHhRop8eOPAyaMFxBCyCKxLkw3DgCzpHsFqLj4Cz7+qV9ipRYk1KzoLs1uYo
/E+/+fzlXudDtSZOEWu0OtcBWWmUUqyGUCa1c4KAEyMXanx4p4Wh32Ut/NcMN8KI
xy8RH8GEeIB7u17LcAwRP6vnPCRWjzWCnfJV6mKupYmc7xuLLCW6AwGyg/vQ1Xkc
2qKSBP3/NQ5evVon6D7dv9Wqx3lX7SeIrpTPhYalj5Sm8dgPkQttjral5C6OysWi
Nulhi5QLcdtNQFMHdAt/vK/4m+M0B+gV3ZkVELAKSFVd32ibI4CUQMdIGXDg8oxX
HOXaHxE70z8gRjTpEQapCbDr8oXDI35Ilig5iMuvrCKUMUrJTCAk09TOb+s2rC/s
GnHqnK8h35SaozSv5n0RBhbno3DhgPTp793H5k97Lc5tb9Ugbf8hmOT+e/pyH7aN
RkLKE4vIwOyGd1lrB3jfqktmfk8emfJybWNmu+FerM+/b6cJf+Q+AfiuEQU8jxs7
Zgq7Hn3Lsw1H5z2E2avq/CrrEzd0GYO0vTcEnWK2Kb1KW7rcryGKlkaR1/elMRM3
zE4t+zOPKIZTBwYb/VyIAYXXAQ9PgnhW8rtBUJilD+oZoIO5qFP/COopJqNgUdoc
XSgYEVXpdFhOwjyr3Tmu3kNgKi8Byj+cwm/ZzS0U3uRuXMFZJWiaTroUOLTXBSUK
agg4LjiiQ/voIvwftJMXk0A8xwNydTQ5s0ocMKe1M/HllGvj7of/pMDrp+2UAENO
iM9tgnyrosaUpk3gZ2hurYo05p4iWEUlQMg8Hz8U8O8Hne+rFXEkE6ZhbT+GzT5q
kmy/nprdzAzybRNQGhCe9wdlHzmOctk0WdmNm2IXg2+cLfosHUAlo+9iYXlDfQx7
japkbTCVU+SceLJJBfkH9RygMzvO/NLK5VkBa5vwrmw5h8Q3ezDL+mkPOKouR6+v
IZlRXDok9pXJ/5ffOP9raZ1ccYMsvSnNAbHQNiQvsF2KMZQ8yZ0DcR5azksOVNno
oK2Wl9yfr/m+PCnJhpZ+LEW5af50EDhy8p6s5yig64d4NbOMATti0iKt6HCQgx+D
Ag7qGeKetzu9FW1XwS+ad180OYoJE2HFQL8FhnyfNdEk+JgWjtP8sJMYXNF9wOVj
MGO7RzHwA0x+8MaDcW/hRJrx4IjykchNaTsxoLbMKV0feV03ijg/KZdUc+Fm1mYM
7qke3lSL11tqy83cWgNPFnjoCuiwd2hbs0R2S9uREm/1M1UWZHzxLFLaSs7BzAci
Li/G1uRAdezYwHqzqb7aRRejQEi4HL40MCFgIoLTj11tSW3uWmMEFchfi/RetvLe
BkNra+BrqeQ2ReATu5COVjMu43bbHDn1EjLT9sgeOfE1UCa1v8OKLjFMmBr6RKW4
4Ikm+zH8DkvHz8ENwkPFOUzfF4rmtzdPRCR8p64ddpehd/CLp4c7pGyzQumLqZwD
00+MusoOspGx7PYh/UfAB4ywdW4lTUlkE/vBGj9M9vUH3TVdWa0MtTOMEl/shbRf
UABZC1ZxmnPzY05lRdLTqedEiilN1L70faoIdku+d+GTMDtbklxNmI9xYQyGASbb
qgjagfPMBkv38CVCPh2EMPQlK+TpiMMY8ybT3op4KqLfi9UYBfxqWCxztyZpoQBb
RC3Q0q8ZDBzK6Pm/+E1Po/c/hUOQ5Im9B9QUBiRQM30nUu+kgvjxheBFWedTvM7A
FmrfvjpnIT3Aeujm1g5Y8WKuWT6TmQcERA84v1xEDVYT2LBPTlTAmU2RPW3WOB8Y
5Fw66WWOTXIaiXSftzYE/T66UB21bkiN03vGMFVYgj6nvm3jdwsafmH0lG3kJ3h+
qD9v4GDXY/mgR5mjPI2vrkW8lX4x+QFM4y3WkOsWT0dpSsizaNXziiDQumUl3e34
dx3SVODHO05XdrBHiTjUVhdvpz+45Ih4QN2M7FTaeBmxkjQWohbDOxiCZAkCVatt
JmQAXhRxkRsdjA8KNlUmBymsh+Z45EFhhEFtGm/BMT54o3tXJk4wM3VEApXzjm+X
rPcVdnvLJA6hg4QUejqVNOzfVBYvNgAj9G7asedlkXvmf2Ei3/7vXwYXuD7Ou4h+
uJEXpcVYJaAsh9bzofHGN90vnggY5xqsTixeHvuWpvljGX4SHCS+ClZ9W1a0R8OC
Pnp0DfaoQSYsgC3MGfIZui0jXJrQA2gAfl4a9c1rxs6vsFk55Z5NdJkaDjNRthd1
THK+KXVrpL16PMnA/SZx4uk73fGDTCMbTEEjOoFTfg70mDY07ZQSxvTfhL74xQbG
6pfEdaL/9F/6ZO+h2DWGO3xSWK92ZbA2ap1e7AoKt4BlYYw5c1z3dXXNCxSoFarT
znrup37rsgLROUCVlLrVPkJsZ27NIEVNMg8XmrCjV05ZkHt39TK9w6tKpTp4Z+qf
CWF9Cw8oCt4//Wr4AS+2cSjRgXgDbUcUGmWT6fULNHRv5LkgTIAT6sGFMPa2CicG
YBRe1n3NzHOoicJCNejfTndawF2TvJixE8Bb60rtjPR7xEyveta/EPOSJA/f6EoM
fcXrh2yTQPsur07mi7+F9diR19dkV587vshbGzvImclqW02U8eG6Fn1xm7wuOWXK
Zo4Wnv2BLBpM3AGOhvqRA4MiVZkN0Nx9ODHKf7GFrcAJeI/WpBB9ro2wOSISlGUE
Jg/mT0/yNf4aZZ2eMiR+6xSwxNf1ei6v2x2QK4hWOyBVXLsYt5hNrY+KfQM+7AsG
dpqIMLkBPrrQUt4ffrQDD2odfFynBy93HxxuEgCK1PPGv80nbpMOlprINQ8BW5pe
aSlhMEZJ0ooe2WuTL8O9kiE/tbUCtcfa019aHi+D/cpKZ617f6SVE1ZCKy9wPNMp
OIV5WLbwJOs/OvpK6zGOz8uSCYGBxrs+mRDz5GXPw//9FwZ+OxRMvWv3BjFb6ijB
MOyHqJzaWqjABTcCrY/uD4STJtk0HZBTisFMlvI7vkJS0eibVYQ+tjwSi7dRjo9A
7AqgpiyK2ZRUvPQxkKKOcIPFkCxNzydhTWUFXX0OLjeCuKUIJIr3+iCXR4EK80Km
oVXD4p3m1qgu5SrO+4s4Sp7AHw3bZm/Irkk0q6qgGHM21FGOZ855LZkoQHJK2tJX
mh2QPDolY6+8CW5XgEcOEO/Z8/vKSrVwN/qib0k/6lXUZnV83ignuPbzGWmcOwP9
ecjbEhb9QM71nkc3/Q+NywS3Mejz5n9Iwqol93p32MvmDrVY264LukmmehFU+koy
n4jtIIlmzkfqGCbZRHpc54UhZaLIRwcBEKfffhZtzp+lPrhVuVxLI/bl+Lwslh5U
ze2tyI1Cqz+xvXwnG3kpRhvOfJvJq5YbrEUTFXFsy5hHl3pP/isqzBNRIQe71M5p
KXBBBhlV5y47/5iwbhwhqMuH8upLLiDGMtUD0bazmmvotCN2v4tqtizf4rTBygCz
qoJoVkJp9Yzzde1j0u4FSnhNdujkSEamMozS7mJAjJEPVjaf+Zrh4m9UmWuyni47
vgmAE+cNTBQAV1dFPrDWU3xkVC55NwTadn2rHdQ+pkXEP8aq+nGkUUbiYAlXQQSj
30EGuaKAs9Ef7JV3dhg3mEGSTKy+8zKNdfGW/0/aL44jYhLbbxoKHIG1RdV5XSyu
mq4IspoVr5SjPGl40ViBSD0T09wJXrOXg/PmQkzbg47oH23YmcC2GH8bQs/tdriW
ykl77YIXLm8S4XNF6l90zUnGMHHRmBwRBNTfKiHvRQYh1tkimN/bPWSq4Y/ASshn
EaxDfw4Gq2wZW01m1r2Ai9U8ZBk04lFMsXBCHp3n28yaTjkbFLh7se16lXyBOUhc
ieJn+9HKMj55LYzLxusJJG31x0Nsf6FlHqXq7HSZp3CDAHaTqEi80/cxTevy4nep
14exhgVfgU2UNR2v9V3dcIF4ZbjhmMTOClnYvpbpPMy8vfSbMZp4ilxopSXOwS1P
R8vY6bdnA3/FfYYSgdrVcnmZdereid/BX597+K295wapIvVYj/BQ60oMlUFd6MZK
CFJldZmDXxUAAKmNiGBABbhweTgrCjKfMeOhJaKoULtfj9oglX3qIN28qthyO2zx
jX0iQ3/iHwLA+RCgXLLU5GineWX3CGdNGTYS/4tWiZqCnldULbGQUJPgKzEYKuIS
L0jQSxAkEc+NbEv6MiNe4tS8oTySvtcIx0vxndG5lPjRfo2jffZJShsOswcFqBnK
YxAikT1NOlRkv9pr49PNGkII7o/uqlbyrvfEPAlwG/f3c57zWHTsJnK+SZP0Fgak
PrNYnTRm02a4eQjfCYGRQsoI3kI91R4VaOCHyAzHPMFFzUHbcYWj0qRvd29olITv
Ye5fljnwGa1Lyse5UXDe0dOxx+5PvWg8RWmfk4ZVses3zSCkz2LDvYd8gsJA28IN
f6SARNh0J0rNWkTGWuM6H0flZxmlNz8DU2npld2V/iYNeBNmbfxC6i6RtrAYrtLn
VXe4zh+oXqrCV05mdrTfDqVnFxJz2Ip2AevPvesuwIxySAGuYRja3IQpdd7u/ttM
C33/35PRsazuqa+5cPMNAxoGQB0Gk7uLO8rE1XgoIuoKUZHpSMzsZY3dIw0JYM6l
Jq2U5cneLkE2ui5/rba75/81szQ0dqK9QsfzPIfyeCDlzr8RjdSY943FeG6BWn6g
KiRFnw9bj1NndnI0QMRtR1bTP++zZU8ugzm9IxM4xQAidC+8cCAIulg/KdXm99Pe
f2zhJ94LlreqJUvAAOk03dhdrGAUxBCNvbz9R428jSvONhjCra59SlL6VEseN9f2
3aLGARZwouAKsVe8uXRVWRdZ1Ue+NbFblLOqPtn3Hov7NbzWG7o3mxBob67fAS79
kHTl48I2N7B2085Hf/BPC6Q2kboRiJuf8dDCZncv71rqttzJ74j3BpgZRUANN/MJ
NzG1bJGHTMZeRfR6s4mWumT1ltEjAPB38i0LWpGCdKfNh6EH2Mkn2YVQeTewCZ1R
GwztubnnfGFfxRGviV41FarAbbWqYH8ajjArllsmDbjRYdm7KrPIDmux2up2GB1d
Aq6ugSqVeE+HflsNFHrNiRypR+I+m8wq5AWxGhqAuH4HATFuMU0KFX3OVqwVIsi9
cIipBO7XHhTuSzpkS0OFU92+wK/dMwklpLhhzALnf3/a6QzTza9SwBBYwVbeJQ40
aSe/wBiuwwNLiXVDGN0ZLhQceIxtDrDkN31gOHQtfVhu+kyqe374pVYu4vb0QOcn
+KzWbZzAuDwsbzzn4Okv0JQSG0RXN7kkGlJKzhMAUr6hsxB233VIw9zqiaylrFNc
uZm2dt4GZlpap5KJUCnActUB1CdLfbzRrQ1Ix5O9cY5cv1GDjb5rRr1TaFZb86OC
DESGT3pHZQPS5riArrsDM6aNXVygtTxu7g6H+reEN6LsZpJBSaKNFjti6GIBeDCI
++xh87EX2yOULoCN9p1YcllM+b/Wx3yEQWwlE7zbjtTMJHOAzSopa+ludDDm+amo
xGDD6hOh+zmHu1sdRLk/+nQX+NnlyEVpWgP9CP/L/cyAixc14LgyR6KhyRHkRn0h
HBM8+NLGkJ+pRyyP4vkyBj+q8YzKuusxxjavdW7QdtlYyxI8R5OMeR46YRpP2VSe
UCaQ+Yw7KUJbFoYVi1XjN3mwHYhoRhjxR0HZHvGJtTdlN5I6TSMYwtgo1tAYiygm
Zh8ZQGKoky4+tSyexSJTmDz7GN6WwEF+RWbKojH+Fomz/u9McWSbU3NfZUNOxio3
LNASjX2hrvMap/7IMrYUH95lvLq8vfgZFCM3GTrPqObKxaAE6XRDt8heFCXIt1e/
iFWXtCWzIlnUu7I1eUWh0hfq9J/tfEaK/rUYy2r4ru+S4w2xr8nyDm6Mh9NiITIj
baMFXIqHhQR7AtC/AKaIzuAWqo3jRuL7J/M9wGhKLy86yv9+4IVx8Pexd89V9UcS
39B8VKoS9jiT1VOYCFS9i9rDVZE5UMc61rmjidQw3MgTIHrWkYm2TH4qq+SjKfOD
BvnERn0xWvWPNj5ylcZV7Sap0xo3KU7PMlRUNdEJW0bwBuG6kTasSODDvmhgSZPG
y9CVs9VDoUhqCvrQnJ31uR7z+K/Y33nuylt3l4yR/Co1UGMwZdjkHIVYLnHTyDYD
s8RbKHHopFl3Sl/hS2fvsGxmY8vkeIuU24UZX/q9lYAfqbqlwyXgLlkSMfYGDFh/
YV6i87UadDbX3Kb3Ik10R2LHHzovI8ewdIn9bjHb8XbIF0/lNRnDBudHm2CCBblG
ttkuZJ24KXDdRa7qgx0aUtCHvhZsfXVz1hgo/jXZttUSNOY+wWPRYZAHvQqtkmWr
=======
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23616 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
0DfQnd5hIAXb2OPobVGJo+z+/IbfxvW8dMGIcptpCG4dKziowNKU4uGneXQOi+sK
xEaoc7WDcegBHnt3ogGBgnLMWf5jN0yWRVyCGxIgsO6+HyVEJugybJNPuTy/R/zR
WaTKYtpriHgLEi9V9Yvw7YNlsZvPgt5PkblFexJGudR5PzUMRie/LGEhYalYCLCe
h27q91C+OhRTpW0FITnXRbrOc7kEc4jO5PV2mIt//vOCWGCOkP+1/alExhRHdMWh
Fs8ofQVy69v3iW/jOvXcG2RHoowPb5M+5GOBinVYiUZ72lSAFzVYDwrezo06dPIq
XlMRJIkzgo3Yyotl5sv0wF9upved0GB0ojPj4vXeGCZpt97Ieqp46fF0xIhOQQWU
HVKr007lW0nffUAnQc8Bd+xtAbCvWPSR6+IxJ2F9JO9PfM5lndi754sKiOUQ7RkC
XPy/shal/TWtfyRXWQom+fq7WU12YYKvJ7x32UmVE8JQeOe6Csf9lMizNPRX9oQa
LYzkNlOMEVg/L8vkRgeIvcEQO9JCg9xMC9x2hu8ropMfL0NLChf0xG6BzCXCzuWd
HG+zTHyfdINZ5qiX6et2qkAZ+TJNdqmhP4BnXC43wLu3yR3m6xWNnQNxl8oIjmUp
j+xhG8pivV9QIBEs1M1HfMIos3CQbGG8MROZiXZAP4fgT9OU9UXXwQetSyndeUAn
40m9PPwoyufCTiuhL1VCtWHZ4myqWCPUhqvaUCFUuG0coiDk8hrzau1PkGeYwKR8
OVElPK71SXuXKlxEnDU8UbCWm9Xf5daAZQbV15ZQzguIUP+6++VhxJNJNsUYn4IM
AEzW5HKlE8OL6yRr29MnadWJMyDfA5lhFPWcgLkuxP/zpvdi6jrp+e6gG0vZ+VQz
4Tyo9OEKTmraqlh8J40XRLfTfWHbMic1X81VL7N4hlY1Xtr2A1pIxfg419yXSjDz
bFj3Bh5XI2Q71yUn4Xd1/rziTY+PqZfmL8MxtBF9zyTN+mtEIpDOLqruhS4h5Lk2
3Ot6JCEvJn5cuhLtrHCD8GNmn//OLr5V21kbcaU4j+DSlFtHbR5TtFSaKrVcOxJK
hbL+7QQxMNBIPrIhEF3UY88Wl4324omPaVV0crPMDzykHsdkv9/lFEdIU7LHbMLu
paIcrQhLxXrYlVtQjAZRXTT4vEbFCmEp1z0xjuVUV96JEpljDZQzV1HPuLyi/utK
kTHzVw7S0z1JiY8ngklnCmGIQ/JSNM014l4H6iVhATRGRtn8qh1NCCUyMNDld0Wr
2j/AKlCE17GiPYenXk4gv5s/Ob80xmsr6Qx7vLc+T0fmbzVg59MzrWuUsF2rfog6
dDxzVcbJqPG4n6oHv+wXxWHvxLJ9ht8tH25j/QMLKB3B/0Dbwi6qQBPyjW9FtB7I
BL55v4lqWVJzkL7tEyk5CTn8ILerG9xncqA1sdyqIHLcz8/KymdnG8PMpomB8gqB
kfO7A21bmCxzESJBydKRe1oFwNLB9qtSkyEP1AfVJbO6IGLstZRc1bo3DYYjrAO0
XqRmsxW8fUpz01c+eTvy9LIzaYZNrrV4UWM/gLR03uiKIUNtOFvsJT/z7AGYV+4Q
vcqY6baxnquYwjfc6AkjjjgOA5FjdpuL2m+yDlRgw+ocrmLEbyd9loP1WHBIpQ+n
7ANev81+aCAV1lqXSssvYS5bfKldPE5sfq1Iu9gs7jKprGQ/yFAEO6LL5drAoRur
EXp4OKjEvUGaBYEWvqcLXR0s5psdNSta0OaGkLt5eXiq7gNhFkZjqmIusmsZztMM
cmgqYBZq1aLvgilFMfB6FAs2IdJQGjbQAjkNkLTBw5vDi+I2zEHkIdlDQVsLY4Pu
WuZNgTR+d/VuehRrsPffjdj6xEUDohH4VC3PHku01lTEDVG9Go5r+SdwVZeel0gh
xIUak87NxDdvCIN+CX0wUz4vyx0ZBExsjgNx033u9DUdGwi9GzOQjHcK3FymUbjj
rpc9JghTUlU+JUTYACE/5Cv9xBEXpnRg3v0gP5zuO7ElbawCEnWx4JrHcZoitQTR
h2gcOYz9xgXK644VRL75y+lA/G1/xP6Hml0m++RS8MMA6QRDphXrDreAsUTVKC3b
SB2LyyXxftbXUz0rXW/JkOUKaMueIKhA6hK3TuEWvneJQewVDACF6q2QfpusGi8D
+85EktpKhD7L3yBuRmVbZ27ZXuoYTC20aKFSTBPChteziMLup9pddvuYgiqpdtvA
CPGMF3kqchkiHPF1VfrNPTEMMofbwst2urXDN+rRaAMEHTx2Z9jBgqhrvEPltprm
UU+mky1z8/rSLwiU9q/tMa6qecmJzd4v+pSvH+TX06Dw2G4jtj7G/HF/tACe8ad2
HlAXAS/welBlcM3DJc+ZjRQ9/wYkHqjBVWurgvnQ67X/+z/amJbIzPbn28jhgFEi
rGpXuvsU6it1k+5hz5yytBh6RvybVR18A6SYiD5bO/b/c7frB4YqG9jfEFi9nLV8
YJKGmh0U57QOALac2N0lLZJXKKnIvASFNkzLKS6ZWLnpW+Ri2Lap0IosGk/PmQqv
BgdcLO6gjmsu06jZxMuPoPO/57RecAZBJd+stKJU/bXp005M//QNDhv7FfmnC46H
52P/A/jkhfvjoe6m5L5zBveLaLUqbqdbLYrbE5abxmvFTFSQE6ii0TMMkiCwGonp
UXRRKylT1bPrNDC8UTWL785Ai2DHLLgYosHOxTzRMcq05RsxFnE8Yi4E57C8I1aD
vy6A9ysw+60f4A0qnRwkkl2fYdlSLkjarc/ZVcNGyHi/wphr6a3YQGwZW2ftKSbe
QOdR7ab34aA6xd/deNZ3FqSu8xRyePwd89XkXAGfbj/ZKVeIEI+QnTwRfFOn1GzO
fA5RIoP9TvU4lOiPkY/H5NTknW8LQBEWMkzdfUzY8OqJkromWQ01f3b1JCXI6LT+
TNgFD+QDlfnMGleWqGxFaHfgWP/htP95/QFDvtG0bLddPnIuCjqikOnhKvL7bOE1
2MCjfzurGiUSwaPtoxWlsQ0iF3DjQIHgwAdSxUt4CqX6hwbVZv67KFSNOMS08t+/
xY1X8w3QZM4uTz4NYxyzH27K4gDTvQvG5HukDqCOHBsSlLlax6ax/nW0tPjn0eqB
USJ/HY/R0/0lyOsE++KUVfi0dmpj3Hz8eLiW8eiO9offGO0wsW7FT3hRk/tyy0F8
3KSM4gwOStuzvIgVtldpHLMMU9WOns8NZBCDirrwHgJ7XY/1b1r+fRPF3l6m74SD
0ylklfj5OxiDMEzPfoYW3+0lthsM+4MsbwlfLbscsyzQzjeZSFE+bnGmYW2DTEA/
4qAO7tXrGGPmEZcrOGuJ83sX5VjgjW4X26VsnI9IyMvRW5B563EQEKIBnk5g84eA
dP4zwcr3oKGpWlUlEQ8gwBLVEImKk1LXmN9ZnmYSmkVHDID6/k/bFRGP994nRo+X
lIO0GIHwWeg1tfTqiUjxU5ML7eOA8uBsv81BNs2nkog65p7lmvTzd6y9MtmeWQ0Q
SJVbg++mK09eqABrY4p7md1llcCEUNQOEQIWcXPRzgRzwe6ceFsg2oM80bUebquH
FMlew5Hh3xW5gd0ydRe6ls6dQ06ejCdepTBJcCdezVBPnH/H8F0W2fmFMwXNBUs2
ruwpnbgeMV01kD/KqDvWuTDzFeAgu9J+d6WkdcJQW/XYlf17aSfzzpBdaETf6LiQ
2jKQb980UnOaBPFCLE4Ow2c6VNu/YpEHwOTLMbQIr8ZEE0vCtqIPTZQVF14Ogi75
P+XKa6ny+M55dmxTFHhBZcfsCaeTaX5wh/G7nNImNEsZSi1edMWwume5CVNuhEK2
dDiy8wt106AiVAWk3TOTAkYxcG3jnGSa3Wg2Jjga+aY+YOaB0slPKAw2G9wcioIP
PaCyPtkWI8p3VHW+3xuVYRzfcHqnpiPTzD6jXOaTfp0TzME/RO+P5/reP1NWpQnU
tCT6TT0YvRKr/1X+J5FmxOTTSRJ8EPQ7VZUfTm2EWXmELfmE4IvV/xUXRDpKjm4s
xqVrbK3ape/P6rdBPuTO+juViCXdNgB9mU+bCMJ59GFzafEsRDsXRrvqoDky7QNp
6l4jadCbWkJsbDiREjfFnXtdy98fH/bfPLUVet6zgg28JH3cwjukGxtvmV6MDZbr
ORTcMkNC0rEyYOP+iGRQ/aO04CamZtw7SXSgQMpnQzIQwRY+QxM4HlAUXjAPOI36
NGWVHnDip0pnSwfbEEbQNrBmZagyl31DuE8qZ8e69eHdBbzT4pheyEkDPTxA5nlI
V8ijT3UFhN1Y9aSmO7OhHNY9IO5x5KXqoT63AOUNn1XsK9M+vfk941kcBRF92SNE
6AM3ZUfJEzmxi3HkiSpjnyYnw66YnzEhz/uKtZvlY0xKQIaAoraXqJtbfCh15kED
09ariz7zesoxapWzoYvhz7SbKdllvhU3cXzbAAg2cTo1L/D4iLp9EFB987oi9/hy
nR+WZVtnTikho1OLypgkqYx/zFaRyXLbprnnvPLQseoGT2c1J6dMBfvxlA+Ylfa5
48MtuMQi35FBrS9Hzs2OvjYuUSf9iTC6kPrYRAmroMPcZAtGKS4MNqVVrMDcGxQW
fOw9osCptpC/PfkFzO625h7amr+LF94ytkKlxJ/CIVK3TJ6SiEhIk25GsQWVZfVu
8eXVH7oAb08D5JhV6XS21dIxwtEMr+J/eRvuHyQmlu97wt84qo19siHbjc4EyeI+
omZwSgULhRDWbgvhECg5sFTxRLtjquaTEEmdEadgzQRexkAzYzMFv2VaKvqKV6CS
UaxT8AafYlhB8MS1OVhh8ulFwjDcX719hYxk3aqJWUAUoxge8vuSZA4f+gMOf36x
9lUN+B+sP6by/XclTSjyTehu/tyxuXv42xl/eOS064JcWEOsEkrIsI8sco5PcHqI
h57dxYl6Ct91K+vluTF0D4fgDTI0L6/iwlzq+JzDbprD5Hs0Kl68U/aQkg0bBl5h
zqixENdjBWP4lQVmkfpoiW0c9bhL+NDJzIpZjgNYqlwCDHOBiX/rWMoPzKGi2l/y
DBB+GQOdcKRRhHPpyLu/CNvyvx0D3o4tBZxvJ+Rxf1vEUj25WXELp2W6Zh5YPOQl
Iaql8SM56HTAjvUHPs2OKhuBgtXYWLBOUulBFuKkwfyM0MCUqLLyNndnL3aGOHSj
ixKUsU3+nABPyW5lOHwGaaYHeA53Nk48SIIDHsSybftBPAPvTDRxEA54gqgBg/4b
y+LJ1AB5ZaRH0UvEcPUTd1u+Di1cklH4gFy5AXJLUB1u94jovOFeqDpbNiqBij7v
2SJvCv/MJtCytgSwJs3Uig3x/moeMzJfL6QBD5ToDYAXMj4poNJGOhAGgzT4Uwb6
pdeziWyMG+df6u8+pzYDQd8wSxP1E02bGM314u38WQHrA7tcm/Si6ibBHR46ejQN
llQxmqvrSaT846QEzm/sS6MstgMjO9iY7I15te/rtOvgsFM2ZFMt3mWlx6frwojq
n/vr6Lxx+d1RH32mdByZyNARzgzM9hkgVq1DUleB9eoKzKBBysgpghaEyQtUaka/
p0bgtCMBDSYohtxodye/LzX6e7OojpzQHS6Soe2Yohn7pmsmFUY/ypHhs0/nZ6n8
PF8wmCu0bIrJSB9ktMCWdK+ZGRFjKDPc7F1Fpf/a4kwWLh433rguj9eZcOv2x+Mi
Mc8Hpbmlq87rD+pxslrrNloX2iytNsz/p6dswqNucmz7WJdZDUHoubLreld1DpcS
Sq2x0YIz+DkidytrJRMp9UnQCoVJoQx7edKjYKpyaQ+p2PuQ5tTmZNQkinO9le3T
YvgojK+SK0jnGzUfOz3dpyeq1UMx/nDl+1LTdPYbXYqp/oSSmtof5oE6BihKIf4y
J2RTCtr0ArGVdhliRg+LZYZTkx9LmeCiOK7KGU7Wrngg69IdTXhytr13koEQfKi1
GKhJasE+q5VuAWVpj7TMGqf0K7mGISd0+OHe9Ri9XiZ8AOo3Alwm/9edIOHaUdMo
7LA9gYNcxV63abyMMY5UVbn/IfkPBANIbAbP7MAlmP+ilx8XIZfKoEoyRr9Ieurl
glUSlgmLVlrXvC1UB5tq1ziehlEjEFXj3UnyyyGVmMFMA/eIc2Cpfvot+TD7s48J
9D1O8ldIquInTN9+SnMxPaU+08LrZL3ig8A2ADQGtUmuLENGk9LoLbxkVIFg0+L2
ERygtBTWomWL+AitThTnZMj8DUYJm5eVnz/s2R+Te6tuHkIwHVGk0cElDLGu7X3s
A9dHCA2xtn8SwykhVQCLgd7zDXc667ynP06vPd2KMQbFAFVIoUBjC7zX5v87d0PG
6PuiZPTFxeGiMIMcCjAiaAK7nG1flDZeMp4X1LoIPpME4Ry3Ve13TiiSsKeJkKED
R+Lup/yv2u6LGN2pwPQWGgk5ukjvLAE/Zr+uU4eLFUsuArvr7xlbGj9zGauWu1HR
2nt5EbwYX7PxzDGDhWkUAoZYV5Gj8ZwtOPBTa8y7rd3pGtVVCwAidWQ+Dg3SPqt3
mb3C3xhvq2TrdwttYPL9trYbCilXMzRyw1pNiUlliqTERMMBE2+yGaWaVa2HJ1Z+
rNGx4aqQNuVtbrs5eFDMY06H4S6W52gaJtco+srsbfh+yBbhX3amN4wd5EozEQxZ
6ZlFu5vswPHLlRlhnd8x9KRiNPI3zq7vSpq20R94QlTbykS9W9++/WOn9pM6dv0O
y2/4Tr1ZK+0ghjOnOQL+B4dY0Ifyq+6ItmKFVChDKXYF1jNBFEP1/jra4PENf8Zo
czqOaJwFN/kfyp0Y3RXdCCVtmmoWYH5r72uItThLPUoMxj+MT+b8pryDdcujwx5I
Z+l9KtNrOkYddBJJKpPnZtO9Ezr/KLo2veOZ1/bXz1jGIDQznlJdHdGgutAGVgfj
a7XfwXPdiM0KGTtnml8lUl8NESTRJAbI1JvcQULazGwWamTHeeB+fLfHx9bEYayW
keIJOLpTgFlu0DMq+UwmAjaQBfa2NW3pGEjdDijQNngepGyYvRZ+52CD30mw9QEY
vq9fJHrRE2KSKuyzx/h4ynWlVNRFRAC+9EbxYmUsCm7cR3TShPcGlrJFYJ2tN7zi
grsutGSSkQPVptcG6sVqFuGCr02THufwj3uLfDnqqCRNG8S+1yOSuZtJZ+9/CUUg
ClPuILIWyacNAD00QLGH+BmuVSh8d4t1t+53DcwyPdwhIrl+o7TakGRvtZ8I73qf
ecMWdcTpHD4ZbtN83rI0qI46jjsh/yglOXTJwxJboGU4VD6rpVIx27WQshODtHou
9Hx36kiLfq5tETAIa+BfMRkNc5fcwaSKy6tdqrqEmp/m1NPXtVZKaGDukJxB/AMQ
R20r/A9bfJ1dAXDhnJlnDHtQok8nd3iUkaFaOlbe4tWVlVLbfjL9dfBfpLvX5jCP
5jaCUMa7xS9Yte2f4nM7ubAPXk4dv+4B3tYFW/Wrf0BVo5ZJqqP29huvef7xXA5o
vhQ/Buj23JQExGBrGMb0w5McVdC6PGAUv5XLMaUMroE3iwCLj2gtUdIDTZkdiJSj
iDivrAZsqG6qjEePquV3iQZVD5w8e6isHhVug++6o3fiF+99uOeGCvlway575obl
Q8Lc+gtL6pgD0XBxCQsbSVab99KCRaBYOkq1RPHy5a70gBkvhQ/4GELaZMFinSQc
2T0A9+hBDM5ZRoGlMGRMy2loYK0ApARJfP8S6wRwHncO7gyiRWTaQdbI+9VNn+i1
j+M1LcgH+brrnDmR9jTawEVdz94ize82kYuASK2oZZ3bU8/UrW7TDqPpCcz7ME+R
6QQq4BQcQHscZHmy+tpzGuoV4UKv9wCbKmac6BlOW0amfIPJniBJgMVG1AwxlJOa
cnP5V368Wo9t7tHMpxJMqsQPNuA2h1R+xWSe7p7czv1USvaijEjtqYgDTWkolCrE
859ExgX52AEDGjDrtIC5KkEmCPcUJnjc2qGYsXmVoatKs7nxuNue6acCCua7TKDs
2ponJ5M0risoHKmI6o1OceeONtoaKVP+aN/IHbym9LjckTngYIEBmUdnv5jr1SWU
1GBXubkpwot6HEWAttebEU7X1t1KnANP8xrhiKYhHlnp+crYNTCu/HLm98vDIip2
H5OOf3Q1xuelo+dTJ78KCxybjEGh4NcugKNpYQ9UyJqhwCYn2jozamxDUGSqbtDn
FT2Z/uFiIBE59jr6tnCnZOJFfJWilOhhD7avXHSLQCO89YjPpovLq4kyi8s0NU7I
AhNMZZXWOsm80flSog7Y0LGWb6xYx5JUPTWWiED25ykuHZBtls00QppGmjVGk8TX
kXcAyPJ3LG8sQoiK/clRbEUriEoUSTQI30ld801a14/xdPqD9cKH1fRXQ7RUX+ZW
yCFFYGLvNbt/rsCWbWnXqpkRZwvEMrue028+DPxzRvTfg1JnMiFqYaZnO93fY6s4
JleHWK9sDi5ZTH43AH7kINBxXvGjxkxNHaB8dA6VBIjU+AhCzEQ3xhNzkl16+inW
7k3R2Ocm5gQIGjowbOgv6sCVEJX/Lxp7Yv58VoTayU9Re54dbErus+rMMuZwsD7k
bHybckOEGqVHlmvzHo7pY2w1sV5zdU5ngk/4NgeCdtwWMKz1nbNqFPUUAt+HCS5L
C/C62Qv4ZN5FMatjCIJKhv+2qqB6ImqUEhCInoF0yNkjZYWczgIwhmnyFhcCgA10
8yTSsvW535Ts4hAR0veAvalPxFha7BkNZpDaGr/1rP/Vjp+rnEdYzBTBAe7nMIiF
6Ik+6u3hHZUq7Qe3a+8qvNstwoa4KWPe8KhqcOUFbeqTIwaAf4cFaSazfxgrCMxl
9hJfTB+t/90PGTL2kcoPkXBFXjAMed7uSGy9tYhd4h9/uIVd+L2oO8A51AHmn5l6
3J++ZZL5ZXkY9junQyC1PL+Sxziu/dPVU7w+1DVMxMf1hZx/cULeSsNsvCmtve1L
pc7w0e9minuGFnlmqd8K/et2QCP7qiup5m1FM1EbBS/yznYjiZvv6/1GYF4WFzpi
ZKMks8l9i+Iv1NCLAU95Yq6WTaw3U6i06CBy8F+bofnOcv/A5/4YFcpmQDnkBeig
SrjzXpSMO1bNdA8Dm+hr3U5Dpba9ZACjVQ0I/bTgHIa+/7HFlqBn0lzc0+cOkizF
GwiyA8flAWDAdISyI2kWHBmneVYM6FRKzCCkv9V8aLxWuoNQXoLA6q3gHCZqaN2b
muGDpBhcn4ucQVYnssWTcl37fQ0PJPpy3zb1poodILvzx0YbMhSMQhetXAkD6l00
ZT5KzdxdCH0BRTEUvtp+l8nWxzcgnay/0RPUbOTb7PJX8YE/u3+bFrl3Ots0GqNO
DO47CKsYTJcAFhJGQCjo2b/qP/D5v9ANf1B2tdNyUCpGA7Gna8gWWjDTjlTUzsfD
iJWcarTuijJ1R1y3eyjTlosTKWLmo+NrxSR5G+6VJTnxScSTgYuqGd6BIv0e7uXV
gXKtSbpYe9WZ1FDvsH4tpYQiCmUvTL+9+mAQbTswL5O4E2C58eC/VatcpZ9vaUs9
KrG0ckj26+AEp0vt5yJKJ9AhrsCkDL0xBa1ztcuTEmXzVffdRmfwHePM+rFU/EtM
mGJ60C584npWuv70bECq3bPS/f05bPbL7WiHLL4ImQNoup8T4p3HUDvbJY1k2ZXK
A7zL11vTzBorkaI3Khufz4HeEeZE1dmMu1StCYokYgHhsQCwNN1i3TV7IXwpT66N
/F5iv63g/DYiW+/XX5Vw46WjWObdidtUHfDoYAgsgpikm/a5BAVlAFgx7Yit1RDY
cWbrOWuPkB5x4trpPj/1oifh3f0JTM7saHnOZzIjjp6wwZLOfnm/8sY/ejj/n2+Z
gMJY5XkvbyWatFmQuDooj1OAcH22lyKZOIDSWlN97PGpACvyEvEmLcLmtpI3Heac
bHWaABhZvlKIqs2RC/rJRYUUcgHpVsY4WZYgUGn3zlniYDQI9WrXpQ0Elc3PPiBG
H8nGfin31lx0YmX0iOuF1FyT7/CDchlwuq+K4IIOSlBOyfV01OfEacWJqO07Ftj6
ytZN1v8t2fP7640agux2PNoSMV7UxQX6fWwE783YmHlkGccnprCBOkqI+obzwxo+
hXz7h5fr9jnynXfDsieS4Cw08knxoXymZjCNmpfysP8skjsv76D5+pVXkCnSa1ih
InujR6alCf/l0Ai2XTJzWMGs/ofCk3m1fPw9ulzHnPs1Gdj+Q7g5B+H6gn9KN2KC
zvgt9vmRIIvb3Thkmg0lKCDmre2PKK1w1osgsFTvwA1sLxRaELxQSgOvwE3HWWBs
H+XRXTIwn1GoD+psqRhfa5dz6H6UhHRmNBkBQv7IOpAxSSWA5mZrnBjx27/j9ZCk
lziBdRK8F854hYDKxIubuhngr+oLVb17xuYq6M/QkUtfRZhMWpWyVroOPzEG1fLN
U6+Yweh24qTcgHR0+/G9dOIaLblPcsT1UMLFkyFHVwkOqIDB0NMdJsSVVqxr9i3e
MyDlrMy9XxdVYOj99hUEFZPSf67+NjPW6OXAJpC+YjE48SmaV2tKcgs16Mo04Wvw
Rpa3XvlfqlojaADuQWoi20/GAuAU2AGApch/6hh3jAob0CZ969J0qhPXv4VHl8MI
8YCSnCxT73y+6BjLEPHSKEjjZYivU9pKJlEm08RaYEmhExODWxYTrHZ1BqPRGJaJ
0L4StjV+pP3EYCZrLW+TnrA6e7msSlqXPkWE/rSroXJ4cm8/eGzZIFCb2fTRgl/8
+GSfjKe+KW6rohZ+4HVwTodE5Izero0NMP54wWArJSk4k1OuLjqCqp9bFtFne2uY
yEq0R30TD/+/Zb96CnNqtlnJgnSrlFcbNJYLN7JivuymLXE33hejoanjMzDvzguY
ZjsBGDvAWvJ9OIEw90SjTtIRyrao7WVI3Z+jFXSBef+Ni7oKI3QSobbclA1HagjZ
O2PWK4O5m3jgMty9yJnTfQWR1mmvCHeh4uIG+u7yRucUbOzhPbJVyhTh2MaoOa75
XT4J1QkLAKctARO6Cmd6E4LfMkZf5c1jpVWyKHqMzrS4p1DVuwt1/QPDkVGid+in
QYcZanoNbhL8VnrQ622iz8clQXwnofuWzhlZJQpm6LMmO36NkfDy0pyDMqk7lwFU
n4lopZwDba4Vf0JbvOatqoFeQ9XjH4CKbbAceDH7LJkJdI7wMfBLPhKIIdEHondG
I9NuQDggccGpjxVFcjSgMGVR+mncCG9SqT/NLAUh9rzmFg1IEBxQAHfk/HpfvQeD
XhVLKTDAgsgCRVNiHK3RKgsV7bOgDxTx6d+gF703qer1u8mjbdp6JOSpQKd/K9M7
QQmB3njsh2UVEN3DllmSxzVKwKtUE4t29Md4/+BA9UXqDhhYRoH8hebrocitkA9h
4OSJc+19GQ0YTDkFQLo1cOx4FDen7BDyG4CN1LNjWoC22ZE2RtCKGiBMZW/P5CI3
jpEIJaSh8ycCZ1QPg4auUEaXnKfb0IAntdDXnjhvnF0lwJRAz46pLvF5WUT3zk0k
EeXs+GcOXCPc47Og1DnCBrdkO+pjXn1itAHclT2lyd2E7doBC7OO49eiqCvNfNrO
gQDSXYzqwttR83UCgswQYrT0p8JwzmQSFdnMeOhN51rNiQv5icFRm49MWcXTCRqC
RPxGZXwN3KQLsXEUtuqE1EefcI/NGGVUg/vkLea3Wd0c6YbCuemYBu6E13OQkyO8
K8f9rKc2kwd7RxrBGia3AkkJt6ZeyeJvbrxHNMEzyuaToOTfYEWUatRrNQ+Shjin
lIqBN9pz4dyLFLaLVN3vi6HCl46JMO0gHTLYnghdWA7UgNlczoQc9d1fNoV0uisY
WOrB7+ypy3L8ep07jBveK2gWjvtgt23wKKBM5xwourjOkbpuwrl2RSR3HtVZB7kb
mm3H0K4fs0WdEs0MdtZkesvdN8cLN9n6WuY52TQzi8l7XyyT8Qn4LU16Pf0LEBXK
sqEdK5nhdzD4mVJYTbZookOQy1RNDp3I7j9caox37a0LCEkkSoLlCf6lAHa8HqYK
vbGMU7xfZX1Hfgnk622WBmDYyJYEeIQNc1ARtOK1joPYCPZqOBV8cOM9KQsmC83l
zuUU0Ygq8Gpja/Cgwot5LDSrsqh3MXQ4mpbzcLPOV54k9NebSWe5FS3McKtxkLb9
83d+NVpMYwSjJw0g2p+zkQLRkOWZG89h8jKGFDRqiZdDJi6GVjhVO8YIdLEwelwS
PVqCxTQ5jLmLpB5EJiIpBIVTDwg6CV5QeOmSyXLMyEeO2ygMfTN/ebjG3ORWY3Ut
KIthQsM7jcxxUeCikIkhyBCommuKPJDm0t5cOjV4KABGUNI/8dmHyFkdeK05bwic
7LF1kx7Tic1LugFO6nsjpszzm1YSks+sHO5vp3qlTJAnOo0J3doboEhlc+H5GgWQ
4erxsIJ25cWZaMdThUCSaOeX2XfLB6Kmn0xa0a641uN4gtGKktPC3pRqM/Ev2gfZ
/TjYC+HDYo48cTaEyYpLSOBhrbrQztIsjaw/jLxgMJT0nlaAf3gHn3m13l8/S2cu
JCHF1tOP05mTiEuWw9RXSKZc33QkmM5G6U056qX5SZ9/vgpEU/HG+MH2rAoFEeZL
PFNSK/RpUjNUxIdk2tH5zVNwAMjfcpT99UYaY/4G4cpgKNBaTowTCjop0TKIX/D/
FB9iSodAPDDb3AA5SeLgIws0OTPQ6mvRUT4FtNnF7Wiu3CZ6bwchdB/1QSyVfQ4G
u9yN0qCfDYAQ46Hdmth2NPgggQCjRF0tkNmMH5cLNtGXOyugm35ML+Q8r90dB80N
NHABE6v7WX+u0Udor79bLHT0DXNFzr4YbeM6H/C5cM4AYC1yd/3g1nbZyI8IRbDM
OcEn37pgTg/pHZU8B8fFpmScjLBdIzQ0/NMOSlB0nYq/i1un5Hyxl6ZS+3w8i4m/
WDOARm2YPamWfH1W6qyQzZUQrh8fhk2vgx6/f1pmdEeesYJM0V+blhiU3pVdgXhp
DfUyeSWFrSOTF3N4E161TJzNSbE8jJb9T7z1NJs/limA1MScMZCBLHzredUftFai
RtzMy6svwGacjnj1qLZIZMUwrX/qUahhMk3AdyxrnGCbGH9EW/X8sajvDdQgDcBT
8c7MTZ2Z6eBR41bNEFEtK9/RfHQse3eAYNnAviKCkTCnttfnPxN8A/9xl6vEI5jj
4okzt+ct3c1BQZZOpBFMvmvZMi+nWYFbMk2KelZyoFboUu6RtQiXIyzUJhllS8se
xJb6Y5oexwE04SsdU6iSFbWzzEItAVbOuL9ANHyQUwE3EmGKBB52DiBCd7gPbsUq
DmIx7TOIIyT/VDNfipJ9ptWlR84RJbatMy3IftBOQD4l7/FDS5sDa64YOuI57XC2
oFu1MX4s3c2ewhAfV21bm7J8beSiPK6w5pZ0zg8cag4BKICW1WR/Ku6zKcOlKiXU
e/MsIPURD7W2BlDVl8dSaWA9ye8MMr0Jekw2beYNROZpfGxPRhViHUjWZm5420EI
8pYNcCq8B9AKDlQiswAGx+7cGs7z+nqQuim9jRyMoQ4tCCujNNayARd5gojjgvk6
KNpuPOtfO2UVvfXuPzDQJSIatmF5muhbBVtMXOm2vcXRTh1ZjH1NPd5x2as52x89
9xlrkb2xZ9bRO4F+JHfnHncysZF/kraYZk0mEtfpY19mZoan39iYJXDwkfVWoQp4
PQxbCiTspE2tK42WtSbXvCQYn+Etzx1qg6J9n1mbaRWGDtrtJEk1kkqs9U7z11qp
isI5hJ3TehL1pWZzbZR1csbHMzcMugxVEBOKQpPXikdwUB6/KwTgzsOzWMOvb7sF
CbuDUCuAPtklvjOnUQewvnLlNbLc48ihMx0zqdZMBmlIdZCfNJSxiRAvjDv1uryc
dE/WmmD1v3XO9GaAz9SMw1kEBT9eMH5q7wwMH/r8/g6nqrTPOkLHhMS9RCWTaVwX
ytlYVIRZEcJeJV6bwXGyl6KGFSCfrd3+mO9rkSuBHULcmzShxykSrdg0U2Gwl4Bz
xd05kbPRzm6T3kiZ09RMlBNjtgJPw/yurFjXpZWfBiXUdVrnZGo10sRv6aYLYOHh
5lnlgq3hVOsS0jB1+R+bgUBjU+H8UDDSOCscwn8ik7PtACOvAkDsKwv86MgTRtrW
t1m0bro8268v1RzjJiFOWpKXi1tGjMucSnYkS+vNLTWEBiqcptu6HdVgOfn0kR6o
3zowuvZ4vcrdSsLUJCiRSYoa80++vd9uRecgLwrNIZ5+3Dh3mZNA8co6yY7raNVu
3xo1c4/VW/+ccxCYaZ1ExfbBqHit5f8eilWj1ZWNL06V+UhcYEGH7m3aqdwX3Rl5
kJd4a3cZJHdvfIZ6+vn0/L8uYvBjZ/GsXRs0cG4Lyt3j9RoCU+4H2sLzjVvkJRqS
nFaSCQdJYXYixYpRDohEMLkm9p+R2DNXhVwsq4f/M1VRfXKc5H116eTknBpvPoha
yPbUnxHQGyFhMUQ4hlR2EifWW3pgw148c+ZtsfAKGbT19oL5UoNz7S1uAHmatrbk
6Ki66bgV70m4uDvWAdQV+UxjjoqfkuHTxPlcM4JMoPKKlzb+KTsdNoAn46Yevs50
uoMFi9eOiDvLsjiQ62+A7YkFCGDggF3bbQUfE23YZ72WSEr+pDqXwei+wXL6rNAT
mx0ugT+AG0PpLKClUwpI4wj5y0xLXEg3SGlpETXs/gKJkEhLFVGyW8jjy4r/BmVI
6EQHjjtnlTI/3pp0hORQSkdwjmi/ckHGmfyiZZQ2Z75k2qNIzq0Ivd6FkwOWfWYs
x5lh+42Rfk+FBJcZERlPPRzMgJ1ipcbl5X9HFZHld5PKRUnde9Hc9h5g4kIS1Ni9
RP0vWd+4pflJ4H0ObmYF6YgNjBCYezjQUdw1m9pla2nK+tDae5HaQ9MWe7n1bPHp
+n7T/18UKTW2TOiXD40SC6okTEWXL2gQH7gyklDlRwAKlR+Gmfz/Ox8D8hW0GP2+
9aHJ8cmewDHJIEjt4kdmyP7wao91jF1MPPGB3uBQgTLfHB17B7MAOCSGXssmh1rB
PIhpG3gIhZ1/DYmqljOdy6MS9i0MqG6UL5a4960Pp2pP/u7btEf4yaZxUnXN6PgI
8capUXnHfkLgC9tZcQCgFdkiVBNZ1se39gSDQZs9uTjri52PZJ/ZK+i+FD+GAd3o
fzoJIp11IZBX/0cEDoqT6fKqYbsjzwYkqWYxqoW1AWRREvuRUNVjjDDuJV+G+6AT
8sLY8FSKuY03SLVMWcGkkLT8lFI0+9N/ocvst2pOwW5rgglnYLj9QmWj0q9Xdrnz
qB3YdgOHeNGrkmYbUjEQs/QiG5N89tHqUQ5GfSp7+dhv5JzXGGpcyCL3a+7120sp
p7FblLNh7LGfNlP1MkjpPj3/0BPD3HLJDKr4+pqegojhzZcpN1mSwVGv2tKHJKlP
XWG5ly5ueS4jU8CDgDeBgmHH+ZWahzfYvm6PJF5jXO7D3JIbbSZYFF6u5CvPOxeS
0zfWADnQq29k4jCfPk7UDZmH652IWgkDnuRa7O88S1i/wt8IEqmfDj+XYKlIT/HO
46g8k/J1mV8C5lBW2yxQ9BnKi6SNHJY1cXnWK0JmkNB/rxj0aIL9Q3LfTEtE2wm6
0CiMKJjnVrHPPzlYH+5JHce0qOiPb3QiHfzzGJVyP08l/nypEDx5ef+jWY9NjUP3
TfYU8o1NQQj+askWEkWRUjSOlZwM71cZWWXpGCp4+0z1B+3BZ+jvCCzqtABl0Hvh
Hw6hbYmWOUKvT7D34IxikUcs3jwQEIrd9e0SBi1lNcvhsrYqYUoBLzdNYK+aJoRV
KqaiIC3+N9IkXIBgHBpPOfhneF30ShODhBjJmHrbsfHn4i798cnZbjR2zc2142qS
w70DtopShSTytHTaTTAaqIB9reL/xAg+4nVeG9G4jOZeLSDAOellxkug/+lD19c5
s0pY7HOXgiq2F4X0HPGp+Ks9YalD6yDcUpdPk/FJiHWzYCzcCplN/NHSmQZAM74S
+CxzLE+Cvdy5A16n+RkBTGrGdLOnp9/NrSHQYZcJ+/enueOLJ54wqyXsHnCgP7ys
xjMEqQjIz/33Vq0icVgMquled8QgqRetKMqG5rzIWK0Le25RF5tKoZyhdPbPM6yb
aL4p1c8/l5AbfByhhR9Na7riP2KbzlUWnF6qj7uFg7f/daohiwHboeu6OK9XNmzb
S0KKMrTZZiK9uRjmLnzDwYCKLrIaBTP5jNdgyXj11z1yv8PBixlfXKjQOVfFEOkQ
pepkY+l55DZCnkYqrhl4GaIXs3W1hVEZlw96YBvbYt6x5z9stsdilE03u7dAjH6i
PVGgeJfXeIejYaFcGwpDA+BLItTf6UfuBMDLt3pUM57yPTik84NsyDf0nFICWEtw
uPjjrujhK5zC4viN5xor0jvN3Ae/Jil1Q+v9gT+PsVvG1URLV9L9JgrvZVNDyBR6
BRUOYPsx/3Dyka6aVcz1lzGlmoQ4AkdynpkmX0NFJG7uCsltvIfXUuDvgsReC/kp
rO5KTG/eyN7SQXbjBhD3cEIIIEDhuDi6gfzmCYuhCUIM0Ap5V7sUC2u4sDGS/PTZ
4yjItDRfdtVxD7ilIUgb3kUDW8Hm5TUQlNDmPycYVFHNkVWiFxvRCNWfGuOY4VUq
ELAAF93msW50xS2DmJrJ7uYHPt51FKRlvVGhnahaOqDF28n+7xRNjcLKQGTOt1s4
DqhyYfnzLXy04923CrGWH4sAwzYo/cxP9Zc4YOmtXud6yag1iVK5odYz/gmnYkKj
JcTyxXKk9x+WG+BekDlrcGySueQJrX0EeB5xkkqhHr7SPk4clqXMJqpEeA8bfzvu
gkXcHKUNUSQUVVPa38hJGmXsARQmlYs/Bn2OL8O43aeeCC/iDHbjh1uCOoUWyuZA
2yrBUEVF79BXooVj3fFMJcMrWieSl55551f3RdIhgG3Mxd3e9MLwyoeML2f6uLS3
mDU8vM5yLWvVXDqFe35ZJgBD3nKS5F2u8/bitOFaiKy/KQ0ZHVmhTEyU6KWg4jD4
or20/BjtIwVvUTwINVkBPmy74/u9hGPf0jPxKqFmZkbPU7tzMuff90EMHn9KXqGX
cu1LX2in+kAvV21Pa4RoBAZBzkV8+xeRU0scx4Cp3WFJd4GQJydp66+tWhZhFcMV
fOZIh7kzdBi+YrR/gxmuOvYYO04BvbskbQKYmcr+PBX/Vo2bwkmue2G94+jpXjoW
si3/nVXXfy8GeUWsGcy488VKz2NsI3fHkSLhHhT+KZOoyNNhPRGNe8bxHGYJ4xBR
0C5WurBYw9ybWZ9bF+rPcx4XEa2tgW9bc+jjRKx7bn0Q/03WBn3ta+Fgmmp+aLwR
+lf4cu3HgluITdsS5zojqTGreoy70Dzc24qMHLkyZ0duH86tV9uddW01Q3Ii5sDO
Vv2D+I8PVFiqbch+IgWFBIJMQyOpez1E+77dMzXSUm6ckbLVcpAGmW/oj2MkjVJ0
Q2OcD4DwAiUd+aROBT19FbPKqzKrpC6UyCUiRuDR+OeNqNB4WrlwFU9sj2U4eyvu
9Wx0K3LpRf49tVyY8FGFxxWBfWnyNL+v0aBe4ILc9q3cuDIqBh7ZHHP+am6ukXaz
Zdd/SlMKj4XVrJHaIVYyYOL78R5W6SATGWq/HCUbkFxaYuQ6vhSOIQ4Kce3qAZhC
lluZbHA+4vaQLnCflvxJLvFEYMpHknBWXHn9V7qPQk4DZQPANhRo0scTNLQ4I0kd
2x/WFVwCSnVb+35g1dnTllTDghOMckqq58qrD1pnpJ2LWcYy/7CTDhAE55JYHueb
V1EghCdAhBydX30hqHKuSebpQNTX4ElVmuqDJxqA1HmlaOoFwPxmxCsctoi4iwH6
dFawZSSqcY8tp0C1IH8FwdddWb8XJ6JXaAaCuPEQp6wg8zrokNJKA+7chsWA98Fr
33TwwFcT4w2ujNn5C4urR3w0opfMePzFu5APHaLt2XdKxBcHa1mUncXfqhgEZaWu
6I1Etw0GeuHczLA28o3tE9ikU/e2CNPijlb8/O8Z//p3dzV73530KsK5j2048PcV
BggynrB65YHrCwAsddyeIfpvFlmsVIkCxgN1F0DmbER19e1+KyIP3x3ewVO5c8il
1yy49Rz4eu1Ep6xvDnS5BLgc9NShKKJyDgYTyHuYJF/zXpU279cWTlpV20FRRaYE
21QKc6sZ/IZ/INO1muO2vWbE2qjOlOL4ZfEOugLNlc/P/AcqxfsAibdTbdErf1/L
/O5XZftk5G+q00sayWtfP502oBwF/ifRe47d76inkn/IGSX8ehKdxGTrWpGzBH/e
eGNTvX27DUj/dOn93aIv89TbI+El6nJnrqlSsF1ARXfQEgWqFBXyy7bTvUsvNEM3
jac9FNAWC+IX7jD7pAIcct1ICq3JI2+K3/qiZ8t4XJ57sLD3YSVgD5D3l8y42ckZ
svnmetFxfTOA7/9knTQYRrjQAqi4gvD0k1YcDj40fqyqtFyWQ1RRz56yRVuLX0Sd
CD3McYMijnrv4Lp7HhWPn7JGrivYpeZ+neGGDTrsDWW2hpKGE3hRs5otgt6yNBTQ
6evLSlbbmiV9ZmjuNFJ88Lw+TNRmP+5nmRDRe17ZQd2KWcNQUoljipqWfjSyYhVX
x4a69Y3i/64orqxSPdIuuWWOftaq6dUwGOulWrhWXNtFXSDqrYMIMJBA6xJEYY/U
9YqGHVPcZbW1TLXDLG6poAiESqnNHbAj6BtcHadp5ap3eJ8Vxo4wal6OL6MJ05vX
02SvZrIt7R/+jMkR6QZbvSuTtfXtGgK9CRasGfQ0ZX2+u0oQImMeV5lViy4a1k5l
wW43L9w0lN03jfPBCTjx7lAeXsnCpdAtoVAv+COqN26V+6e10jFOryX5/bPXxarO
/GA1h3sXvswoG77N4dflfTiLfQ3sa/FJOwIfuo5J+0Eg0aT50wEDc2bU5gz7C0Dy
vBKXrZ2cKNc1PS4uHQzOQtzf4VvCs3v2iV8g5Tyx/Gc9sJ9iyeIPUhMqo5vzAdbD
4myli1NtOVgHIwOtPtEfQEtukc9bqw+SHtNamP6oFZZ81xoSaycqAh5QsrezwEsX
UnbxGX6TOmwCgxTkM5Vf5nGTG1+jr2m17+fq3NxndnwEI5GXwMjaCcdn0WVcqR2f
RcPVYCNTlfn/wwYoT+P4zTWGOSpeRT/o80169aPXwHwpkhYgO3l9a9SFFwLiW7KY
PvbWBewPZPSJQFEnLrw6hy2WDHBNsYWtTYJVTyfNfq3Cr+1hM5/5gBiByZ4v8t/h
jJFLTMzPHDih0RGVN+VzadMNLuNwAmEWHoo2EtJqkLLe7Ixccrb2KNx2ihm0ZtKE
n7Ky+FNG04gTfOUOFqBUot/C03q4xcrVTpxuyrsOLG4L8jQXZdvo0zaxx5ybz8Dp
+Zdi9Co5UsEWc5ADFJvkOCQlSp0NSYRepiAJztFKSDdbF40QGKeft8Z9XEouNIgH
yAx44M1C12wsUlVm4063SYyOtf9+gsVcArCj8LTxVca2q+nLP6/o9pOi/9B25PeG
P62hUX9Gv0w/qd269FygedzBcMM6Kt+ddVcEXPCJB9PeIUwLPeej2rlH3ZHg2g4A
tsvMPyFAGCq2mcmlIJS/yxYOowL1rFPQIpo2JVAkAfhk3dCt5zbpMck++UuY1/jG
6qQHjxtMJGhw7fN28ob4GuA8dWehHk8a35wkfyV6NkaWeNLxgvNbEF7zmFrCiH11
v4BM4FzUEWeoDyofH061kWtoYJg8Fr6du40P7fprOyw6LN1WwcgqsyetgrCRFdMG
LPnEvh9Sz1lP2gWzg/24eZMJUAApFOh7qXEVFVW7MPxo2Mvg/2bVpJ1VKcvoMAi4
UMsdFjThSZAjG5Yi8NJN3FWDWbjHrKOCy6GAVng8wpG1gusHvhmS06RvJ4KCz/VM
H2n9fZ2mwjEU8wgRpU0fMU16Tn6A/yftZJqAP7C0NA+eiBQvDADop4P8Bnx4IaWA
XFyY9vxQA0778zJtzRxlSmRTQYKf/BYawQyJBRWbCb00Us7XGdaSdy680YuvAUs8
ebhdZrLJogIS3hH398bekXZxFGG9undcFwmb2GFgOt49U+Qz2KEU/VZ0cOXXckv6
/cTvz8E7N3/WH/MxuISCmnM/CwoXdbnlC6Cp+lk2SLnwh7C69VZlgnIOMdzGmEw4
tqRqWAoKR4N1c6AOM60wvj66/+F28kj4q7SlqMSs/lEW/5dm5Q+G8w59MMxdFHTQ
Ecf8aMF3BQ8tcDfpxHGm+YdcHQH5CgfgDRCvZBwAC9093L3/YycEABKe3a/GV8Pn
EG2EdD7J6kYfJRkAy1CHfaXgJ0nchF1o3jyzXcFPhleghYttzCdo46EVm8hoTtiF
NLJHViG7bin6Nkc/qjHYZKzXUU2thkd4cgcWn4LT8kFI6q5y/AMric4z1Z6vegSb
n1C0cVAsGFc4KnKmOvsUG1eoCp7nS/A/h/BUgkD01hfUtiPvdbczKhd4yqqxxDFa
0X+DelagM33/xs5qk3ZnqrZahc82zo55hkiNPrOUbnLrVFu8BTgrZpBUSDntu3Ek
8J6lkhYCgjrwaeA4CPrQzZ5R9Ey6PfHe4uexMpdKa5FGpw1ETahzwpgv7EOwp4OX
mvyVOmrSR6vnjKnHFmP7GnNDX1PbwiIzQdK9N0IoqHGyr0avmqWyexhy87i2SB3a
fOv1ILZu5WW9QHslSclQLdDlVcZ0VRLHG2/54ozHdaXcn9XRkIKNDFIZs2ml+Ia8
EFVkGX5uOeh/gZI9enXpxOIECfF8JCvI8wY3yhsDRVxI9dDx4ygA+oO8CJm8aRck
BKIF/nvZcTk46VksrqGoITaQejXQel+WBHuPgg3Kd88+M3IeFc4msSMS2aOpdpZQ
UMTVeVBzlQjljy7L8bXjVmBLzpPEEWltD6vt/t6iGB3ppdmveV4m9FSde8Pra5Yg
chXhAIX+VIr80StxJYdL1iZgh0PthxpsL3TUlbtvSktqHX29DoeTFWliUx4L6/yG
TcLUN0WdzDrJ9I1GXFTgZzEpwkjDNV4WB8cRNd54drHzjLlIb6fvV8KWe5zEYaeB
iROn7Kf7Lh11AUfimmBRtZMPzH8HvvhVm8l3+F7h1JtwHxscWRC6SL2Sp3h6RSFE
woiWsignMXDdLpczlwVXaGKFlbymn12EPGpSDD2fBLPuC6rKGrXo/Om+4lpKSHy8
15HIbBzmoefDNsh3p44vfgETx7QE6mepX3lklq7vn0Jo+FN17kJmzd++zUMCgSqA
smHlG01zfXF4TGBERse97Z1Wj41KJhFslYnUO5EfeKwnWPHy7RY+sBX9Z8Q8XObb
nclfb8ciPjvsP4RmmyhYCN+iWspMwCKGf//N86yWvxXaIHqX1fjL0UhkbIZLC5bg
Oy1xZsbl7enFMfd7I2P+x5B5meXrzr/ZAftPjKUEOrmiN9StW3d63S+ZKvrnQ+TN
TVzyEke4CGtLnrZEZZYgMSCha82h8ArhHwfPxXV2tN3FJvKr4MU7jeqPuz961nJ9
05VD3F6LoHolgZfGf38Cpcgq9tTsMbGHiRMKnAEmPNurufjwK2jhsqOsFgACpXj3
LA5/UfLA7WV2zsZV874lk1nISuXHN/q7VT2s9U7xU+sHh591BbN2bGwW4H48LP9S
ZnJfj4maUGcjQU5Phde2NjfU3KfvO+GCXlZIddPTLErm76kPrqwMrsIICh7q/n3D
FNtDO8Ar9W4nuhixWluJIkXyZa0VEyJaDQUaHxCLCW4uy4JNjTh2+78pwY7aHX9r
V949bokBSA8aO+GG1h67Xv/8pK65b1bw3RvCorxnXCcdsvwzfDMNhsaVMmx0kSq3
qj4i2wjf9UXNQzIh+dNSCMKm6U3KsUqD36Vk+NlPuxX8rCAPl4SQXm2qdAXbraXe
Fp86+gDOLLj0ZwvYtdj7s7Gwc9pDuICeU2w6GTlteGB+71qgfR6eCzUMIVKMysfz
ji9G5DG4LAkkTw+ERKbvNGbdCA8AefBmuA7t1GuJ4CVxuCqwHi5eyucNE11A6vBC
Xwh9sKXoiUwKSQu05i5GSH/urhXUwcr5lPpM/PBu4cjhnpZFkgL6BuwrzN2beCs4
VOhYzRL8V23pfU+hXne9/wZwR9C510862uasY2+W/ZXANZZ8t9zB/U8tjzbtrMOD
gttm7ALeZ+9+vCGiMbgqjXvlyQhgB/uUue0YeSbTLuiKiLiTXVq9k7nJ7HQDL5cn
JMpIbLZnzhawP02ZrNlqA8/DuSZLL46DViR0ARI0VYdS2i0u8jfczd5DCI63LWKt
X+RhaIdNbApL2q4Ka6Abs8irqfNb6949RuLzyrmmRxkvKNp6wjNadI0PA+IUOoqE
Q1cEbm6ErQKPs+7TnhK/UzaVbIA0dIqASDzf4y/Kr7tp3ByxNvckyCoNNnh2O+h5
EKh+IPJ9/renlO1tPQO/rXIx+QnikalaFNJyfZGkF6GiKSOv3WQkjM1F+MI48Rce
H4mcli6d7M0OgRSWQzAzTgYFURnRk5RFyBdFBK3cV2MPsjM7iljwQvwzuU4mMAcp
Uj45xnq+xJZDWdDEfj6dKrApb4x4HNVraAGwKvmjDTIgtLrx+Rg8BD2x2Q0xmxpU
muB+Bx+jnW5zlZ43WDYdluiJUud7Y08owZc4kDiM5pPCHFIhlsirRO27Iyik7dPT
8rGeY4SOcsMXCOpN/Rd3kagc2xR69dL0EkxeOhCM0zGx6bmxsUsAritIY+kqvBPw
VDJa1emHmSeEzry9OT7Akth0PT3FkT/BfFvuE9uE2VHkEYdcEyfWO1MNdsMOItEz
dbkjOjgJSy2ES/lMAONzKWvw6eWmnuXSw0fLorIOlEy/v6Gz+0HTMGZiKk3c7WGi
IvMVGrgAhHShwJO7rSlkOjBzRQKwMrPC4uriNMuNWb13xGpYZWKsniLba8NjL41M
KCDG5XyroB89exCA4TYyCCP4Hnwmyta1bvTrIKS/zbN6mdLhelfKcfV5uY0wMafp
QNngVnfQHNNfDhBkDlo0Y2aJ6JvGPSWE4X8DIAV3JVZy9iISQ8WLEX9z0exHFK1v
a3mo0G15Skn3BLKs1a/2W+7o9x0cTpWcj2jsED3t0vn/O+Z8WfYvG7MOQ/PgDowV
f2ihpuXqQp+MnM5mTRUGpAMhzDl0TEpWvFmwRK4kR3rU2rmJ6fk9iaDAJacSdsw/
VQ1ZLQq6E9r3S7dvklD80cphA/f+Aw0dhn0TvVhcH+UVnBLrL/Zr/59TRzUiiZvf
TPczc6SXLxcVvvFs6HbzBhVwCiBP9HOpN1TFQjX+GjAFX5Nnc54VcAGw4YMC5H/7
bDAmVFp8FZYWX+s6vZ2Au8EP7gwekuRqzgOXZ5zI7JZFfeXi0WTNMZTBS3xfDBxK
bnYbsfw0ZFdveF99W1AlHazhNjToXhcx86cIAt6S85sQS/azZ9bBKV9/mjLmuoFA
CgFSx1GdMk2obVmUI03SV0XzP6fQQ0M1DwXGHUn+Mk5MjmHx6IJ1X+8yu6Hxf/0U
7WAzT4JMTHYtczjXReYx8dZrkVpgMQcQtXvDlRYlGEv8boCJKO9nIhpECutUZLMB
ubUWbGQdIsbxqklGiz8CT/Ubov+k259lpTh1tRYgYYIntfYElTXMmNbAK4H8yroD
cYR+iOzh9GghVm3KSLsWr+6AT/yS/VOXW4atrLXjwcdURktaVklVAGjkycARrODO
9QYHaibsH6UCUVKww+zfkrtSRONuIs2h5nHjUJdCsYpE0f4Ih1F+Kn16rOsDkzh7
d+EqlOmXFTGarB6hk1IG+IRxQGqil/4+lG2hobgpz8zS93Vb3sCp15PTXkUhlZ9L
8iNJDoxW5BfvEFrP4jSzSO1Ru9m3ANBYutUxdG0JSiEWOXXayHUCVhrbwQOBiMxb
pcLwh2NMw0XOHXrZwWGCDv5Up+5sxMeySxrJRaWR3TNDhQwcRH53EXfk3nwuP6af
IowlbSCrNtVWPhnXQG+qwTDfi4BE/w/4osovNooOUk/vb6LX1W/VObueXFmtmsPF
wMd1xuUhj/dMuRAKUGtvXRNCdJd0n/3a7S8FIYJdLUc2fvU1Rr+J6NEHlkb9cxzh
3vE2vYkwMBi5hw8X+6s0X/oGT9ocZeALBhi1jL3YTrDykcdO6oXHKoYsz6ggxiG0
2GoazMbZ6UpCD9Na12KJ2rttzHkxWpX0P1qQ8GLlhnp9gTkUi1hfbIhzgi/O5ZlZ
Q4+lp/Q+Z/DEU3UcENiXdgwDplFbHt/t+bKUxLAnUHRurPgJSieT2ROwrZCsPT08
6D19ol+2oWpiNIkAn7nillRjbohoG734o3+26mmFx7tuEqRZEmy6HpkhGjA0q3eL
5vX2W8FlI65PRNTLo0fkfVHb23ffItLJaR0Z50nvPvwUfI+TM+i5bKmryoHVuX2a
svEQ1LySmuedd81LwjzfaYTItgAOp7hleiTnz/FFh2nCvnHK6Ye03Yxf5p/EKP5g
L6E95g5GtG2iDwBkPrfUdYciW5hHVsyehjzSi+v7/ZiT/E6fQs+H2xArBk9KBXWB
329UAAYyOL75TsFsXiXSCsg7Nn7JXo/7VUkZODRPT5v4/vgH6a79nxu02MrdpkIu
asSrTMB7QkgswIeTW+LEMTV0nLK/ESQ8b9XH0ixy0/JNLf01ORByCLzHh/EenVi8
RRlZfCPqKjZIIw7jiv/vcPlv/L0EXbHRjogM30i4Wc+zjFumO42nP7ruaF/RVnJm
QvnxS+JPd96sYtzXHEqfycXZWUsZoWCleH85+M3wRl4EWuyqYAv2Qf0VQVZfhwPl
Q5tifuO/9DQrrvugopMjmREtawWoBozqJNbe68uDv/t8mBVO/giZzdiMiCVq/ntB
Ad52/IabFuSNLKTQJ0k0dSx0UV3XW/KhfWKBEw2qiJYSpc07LWwAcOUHjmKlrgLT
b7j1UWNr3Z5LomPrP3xiv95qhuPegaYb999zgAjaz8O0ZweMggM39FNHkUhVGqPG
sYrlIxAnHeuuYhrADTHu46ASb+0G1xI4+PzZ77xp2GVESyarl8K+Ua3aU+xwSSz5
PmbBqxNjdML2T4Td3OjRsJzh9GWoZjBzNIyJ/0iU03bRptF37MJQo5ir2j4LGeM1
0FuC5tQYkXeeTfcziHf17gqlzTEv45fIM9i3O9/2eYsKW28v36xGHRn6Yivs7RvW
wNblh/8RK4cBQFJhevxP3I+G9ChYViqsaF3r+mkyYA5PebFGPK0SoC1gj9142MYE
r26gz45KqxcOlRkatnE6dNUVxAeXmpSNKrX/0be7SOrjYqCeU+E1bHDEsYL7bT/q
pFud7pR8XyeGuMn7Ux0Z5aIHGSJoNM4jbPcFM8y84F7W5YNNrZ+y+T3BnpzkG260
6hKJerndp1saSy/KD4rPOQWx9UGU+bcB69SbY5l2JnIQs0s8TqFp7LaaCpiluPsl
JORNhvwxrLIKnl72PVFHN7bpcCgSZX3DpLlmL2pUovZsj2SxOpRWpcYWoQisKPQl
kZypDBiinYu0xZe92D7O4e7fAUv66F5t1CfRhSbijjUZj6bRGwdJZ3yT8Lv0BJW2
s64+FQP0afN0ufwRk3/m9NlTfGNFKN7KDPBBHwhw9V8+KVvA1AMhFJZSLomFTAQc
8mL+eLtLJkYDWTcqgY9KOhZdcAI5XmtF9pIi+gohQomo+OkH72sKJPr9n+YsyuW2
qmhcoNRGvh1hdKrNngQgZgyQxApJBrO4SEQfAphiXYu1UKeMbpAJb6uL2UeXe8b7
ztNdjKwAtAFrQsKGbPdx/CwdNgZz+LlyxLJxa92t9lBEBpvcKOBsoYaMwrhJ/N2Z
susua54TDINezzedSxpaxezEKg9HIpQ5AGKFPuj1zVeuKWADA06pUQKkyUkYSCYI
FEqcdB735Phf/HwTS3Oq/dMA+5o/gfmYh8OxGFWMzCJW7bUBefsf7zhagZhTM6W7
Szg0lLuRYoqd8hsOA9dl1ZBftrMGQfEJrMExxLfCd5UpHyiSMR8zi4J+xz54HeA6
ks2rrwc3LfvWEcDEQgxFMo3JY9gZYnB8LxdsnP/j70vNnEqN/qNCPUJENQCmbG1U
JJRdskQvTmDqZnG1oVR4J74fihTCejjeqjjzeyBFnf76b2MAE7xq2bE9gtDiVo8v
L5MLgh1zRNE3ZXZV79Yay6ybJEi1mUJH4snh+2RprdpmW4BlQobARHcDBpXXQYdy
UqKQ9lpToMuCsfIVBDh9SQifNxv2oM20H3FTZ3lIcf99j/CQnX0I3Bs+5+m3PJPL
K4c10iLL8tcoo88IPTNwReooDMebnKJ9y5f+/43UpKs9E6HFa9x7V+rguTNYAshn
qfqimrXig2jA/DBfFdzV/4or1/EsA/Bfd+4FBrqelv71O9FHnUZkbgQw3j2s47YB
KLmSTOK/RGazG1LpGUXacYguyGvlPQvrcx28oIGy9FlakcdVqA3jJpLkwUSKTrJ1
cgV+0gw1lTRb22Z+aGM/LF8yw5O1t5EjaVAe4oiRO8IYH24KfZFokClCxBtQvhyU
ro6pAA5seEvtVeJ7hV+M3tdPSz6ekFLjZkfCDyWd0h2CMFtTwLCseXTWs/vdD9Cb
+ZcY6BGEsRI0KQ88l/VDCHndmUeSsl5ml/260UeuaCo8myfUP0ViA3IRVqZP8pJz
KXrlPAM58inNqxoiz72EmwddhG/Av/OScNoqMWuh5Cuq7mCUjZC3WAe93likx61P
vcWE7TtozSs7b2t3j6QWaS0HRRHuwSKGNjzRk6PeFodBbNVA4Ux8KlS28RfBLccP
OctL4syH0OKt09XUTviDm8m40tefNxuTVp8jTEq/rLfI0zc7VgDs5mR+3Sac9uIb
kpDKB7JHj02NaUoSObqdGodOT6yWPoDzl8mLYgmvYC9sn0hxOyAZdkJ0YVXXn1bi
zu4tlpspt17zLdeM+HQiINzj/eb/witZS7tIZcPuLABkRgxTNePWuLbVvHs8W/XN
fbRVyOQ/U3LHmGsOuEvCIcahtECMP0oiISEbSN6Hw0dbs7hUelSbjC9t9ZcSDY1t
6WnzsYD/c7xxM+4hszjvmVHiUl7hakiGnCUHOSsQIZGwB0P2b3jQkZzsS4hhFZ9G
D/E0Gwt+NbI8tLCHWhouk0t3M4d823AxpXs+apKpQpEXsXo3u/hP2aCKl6wldxu8
1f+m4AIVXlu7y7DRmj628JZesNobxEVO+5cWhstS2WYkkmPvSqQ5Zl68nFv/lCfR
Z7LcxpDOn7oR1a+OR0L3Bmqxd5LQ2eDc0Ylqq05n2m51NrGgvud7CiXp5cNdTG8X
gZqyt/sNu/Wd0kp5UyGCpojSqXcbkFeYtLJ3asjTo9otFITcWjP4FRTyCCP4CnHb
WjIMD3KQT1Z2fPpN+nSNduIz5QgwLl/2EQLTR4gw0tH3Hy7mo/C0Qn1jqD1YpbZy
iHp0LPwFvASfqPxNomoYEmp4VAGPJ9GhSM8b0N/QNvyjOpob7hb4ebjH4dTY2fI+
sj9OuT/LyeMiDLLOLK0yAudFI7IF3S1GEhD5txcTzyl1RP9qtz37JDm/W28+iD2x
Cvz9++SuxMUBA4ndjOw2VVZ2g4hAQr2Rysy39kw9OGwTb4Fyle7UTb+GyG5XlUkj
COchpjy3CssUUhXl7ORn7b1SFQeLJeq/jX3w0K0g2vysRFT6Mm7tXY2DPkqnvWe1
rZ1Qk3Fj+pJt38UHvMTWnTa0bM+0Sd0ok0/ODkvY1rhACrbEBnHF4XRLfhyuLrVN
LyZQ8ukxsio2cM+gcaLumNgPIJL0aty+1gVtzm6SX8tKTWKJ6F8YHxugFgHWRIhB
iqScHxw0uiivggJKz1liYrGeA9IJSykxTQH8FrR7pXCEz3U9a4WIEo2GGZqYfIbq
NTspoyIK86DTahogv7IV/T+8FFJg/C+0y2J6WNUe50jgf/QfOloKTGXj493IDc6c
KrnGvKtMD1CesM/fJBL7s0FdTKjRjba8n0FklrFvSC9opLxVCnvQpKnBxU8kgc+H
RHQ8x8ZHAv6ergMlG6TECdx4J49lL2L0dPGYMEMrNyJKG9JFmF9p/3/pbg8lrwB4
3VPG8yK7n/zKuACxBRr/6md1FVVQ/QBFekR4bTuDH9bCvPNxF5rqCgvbY8ZhtaCJ
GnwxperfJcPHAWp6ovp5Cxlpf4Xq/SPbwE0ZElnMDrYOsQfWktetSXdTAo/nLFTF
moGR3gsk4Xupvs9xvKrGe635jmcCChI4GXGSD4sGQlnkAjAH+VCMD1EfXO1tp5MD
GbJdW5et1y67qvqRtv38vmiCUDLLLuJKNZVy9k3KL0TLcvZTybRBl1c8iAShh//P
q5FQSvcwvsu73YJ3hvoZq+ZdKbIB627n+S4G1dczGNdBulLZi2BcUBzodFXnb/LZ
4kcPCSPnhPpJmzB8jZNs1PTBYDQd8fQClxk26JOf29Qmib8bAXPq5Yz5PCqHkwyy
CdMFKQaalUuvif/57kfFF8cN78+FELhCgStSZpEal28R4O+Js7M8Ah03DKmUTnFO
RlUpiNr/RJ4e7PJm8ddhz0qZGsIH7wwh4+xIJvubdGA08c0Gfnd/O+77G8062UbD
6TtIYTkkIa1nyyMfqZVhzUPKh3h1+61hzqiXkzalFbvui7kzrZdyCDJh10Gf0SJD
9HRmNR7Mk64YAO82+IYrxLhwmR6wD8IoLBBs8s41mBxMtjCMDvnmKxEaA/1LeMV6
kWq82LpSykfISyl1IFDEvT19b3umyC9AdHtgyzv9APkDen8urv4d2jNwW7Hnlzsl
gGdb3l9hemygz3XXwA1A5P5ClfWWxob89E7SAL9m2xi/lasdwQJh4QDqWVA3U05x
SvwtEGfalh+OBAFfElMJJX2JLiDx6OyPWI15fSYx2J4UtczbDjeWT71UY6znWPVj
f4TrJSpEHiJ8T2pKV+U1ONDi+BCyiAuuttvmje4wEsnU/gPaCEe/AT7g4TLihxUg
LpEKRIP/WK9ucPP0nPR1K6RFcVSLmS9b/rmZjBWshVCGBoL3k7PB84lxAdAIF4H4
p5WFAaeg97fAmv2LPlx+cwMhHbVWgTMm+nz4i/pEmlwpvJ1kqzgOA47Pq+5uhj+i
L8UWaVe0BYc0usr+wEp8WTmiDLj5noHiaNi28JLyq1HR1AxWzGPgPSXZ6Uvv9sul
DEXiD1SGMM4KVQlYvDdXOkBlsfUTCRllu8WlkLkpbPPRdZGSe9p9UmeCAmIpDEpG
I3gn99q9DZzi8wdNUukVepqRTP0ziJxFzRMbiHiigpFzBvSKPNn7g9K0n57JbTvP
LiWbjB5uW8taJ8WD9FHfWh7tfg1roMvHMtn7m58PUcFvyYwn5PlanAWAqkUiWQo7
rqD8QqS3ZvZ2HB12rW0x3klNWkqg0fZpzNhYHipp4fWg/lw5QhXWki0B+flY0GwH
pyo7Kbmng4lOHbu0VRSUmRN37VDBtAbbR/b4hhQC5RRZJwMx+4jrGI5pJHKHTzrw
2/A82eNVpuBMz0lvIFKMDT4WW6DTiin4dj8RwiQecNsrjv8p5Re1jafmuWJefE4i
5VOw+U8okUgwFabuWqsVxgZima3S5Qi5EdqktllpJv65yBsHJQW8NaxcQIEVSxQa
3E1BYr9Nn3PnW0P47KdSUywbEnLce/2DjZDoB/BiYAToQKbI69+rmc4WQUtYoN2i
LnFWrtxmHCcwXHJzIw5HgxJl7srLTNPodByICCL952QwsT+Lwvf+V2QVY0uvQ6uT
Y0qTp283EErNLJNae/H2IwKsxxjvn7sF0oASEHzDMaUmsTGSURxidkqrLV5TwX81
nBIn2tbOyDRKtHwR3yyErg84RrNpn/8xbJ2XXSZxtTz1cNqZmb8HsPOHiCrmSK80
FoTkDhtqbCjT/r+DFt4j7ISQMVPaSks6ekKOMSWU4YUu/ywYRhjrEqdySImdI4Wt
wzzEkPCFP+0QxmH9HV5hNdyMc+RG331sjRq6nNAWJXf867JbAsILlo694/DL7mN/
aKIzysEHQk5h+hbQwHdclG+SYrjjsh87y+ibXG0XyYE5R06ZK6D5kr2Cxr80H5gk
7zwtLyxEH5hg2hK7cEtekvg2eq2xrK3OQT1g7VXCI0K26U3G0dRmaleFFJm3I+Qt
QXXF5vO2Eti72xyi+7uay47fiDSFSThG7t49xLDl7xFjNf0uZVl3UscgeAdhRWpB
YzZ7yWhkl6hTj9NTD11M5hBtf+vWTP+Pv7nGrik3P4vlBDlY9FibVBRWIhFj/L+J
VgrVcIhlC9W40PSuDAG4B4pxdVCxiQl/H6GszTgAedClFmtn+kbAXmXEi6oLpnGW
bsOmHz6K2hNggGIsPCBN/19du/RE20xP/DqBPKd6YLv+F/6yx8djucFbkEpRbLa8
1+i4im8H2/mNONBG5lMfPOSdfBbgvyhm0yJErlUyZHRfbyK75F/dR1EtBIdZd3C5
pE1fEznDJ0VqkFgLfBX+ypEx7BwFS8EP8Bkw0TMYuWrA/DiiTe6AydqV1oKpEtMr
TaeA0vaG4GYygEvZZDyNhdESkLqHwzHblAXKRGfVejaOOgY2CO5vSpVvWUlrYNpw
hvyajLrGy2CPREIzIZAmDiBM9Z1rfUYyPb7jjKjMbJdqCV9acrbwMesOCtnKSWDg
7LJk3EzF0I5GZMzmRIa1A8jXgv6JJHF4HRgBvf2+cZDRxr8gHsBD+5+aCCPdgZgj
tyHwEtraqHNl2YhY63LG9lBhwY8YR602LvA98NqZQI5Jwf///myq0TCHwYY20psk
pXF8+63D9EWfHn/CHU0p/SZRa1clkoAMZb/G5ugEHK3i8iBJYxjZBz7d8qQNvwtc
7iONmHInURkhvQaytrcOl5YRcSjhkbLYGagb2KRtF6pmgJMkozRCFS0BmRQUiuUy
qAgdH6yurbPVrbCC1GbRS5j57wlioICciibutDGKsoFXFYvkYTozvXAn/Nta/HG9
tWdte6UJFdbot4TiUCsx1W+Aty6WfVChEKaVlvQjKS1y+hqt+IKzZ52J4WURGk/Z
gX//iKYxaWVvL0a8Pe2KCGU8AMx1dvW2iTOaJWcM4YFq9BWjplYKNS3k86hQsz2r
CNxCWjY7swlyNwkQwMOecB3SP7h9/mZLrAiD9NXzCZueUv3qRGjHevm7imB7eie6
96jONVPZ8ji0rXrWyWhhUjuh6WCKM5iwlmiezvQUgmtnuCi71rkSyvbmMxyd31Po
6ptWe8K5p3lulQQR0dTOuNieMg1ISNIjLLMIAwP4dKr9QgEbcL/Mfj5VO92s7hYV
7BpYo6AcEkuHes4ZWfq17XRUKnfnBZCKTDiFa22S8EP7J0+oISjCE6nT7WXX0r5Q
SkqjssKpUfyloijGMmivA8cEhtMdazgOCzf9WB621jMym6jdTyFS7nZa1VGjm2QC
>>>>>>> 426889eb8ce467b9c9a9f74dd4af433c5046285c:deps/flexrio_deps/PcieUspG3x8TandemGtyInchwormWrapper.vhd
`protect end_protected