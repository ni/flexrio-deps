`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8672 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
hRRAlfE1xLfeNfywbrz10IjBDB7enrzlaZqn3iPzwO5msIKXDkQK0505fPGwFE6X
3+h1Qn/3/i15h1gyFKBCsy8jvtWER3Vf2oVoRfzcIu+KCywkBxHs1SxzoeKnqLCz
WGsQYZuuKzhEJQIol85QuD/73QJkzmqqJ6G6wkCP6p8J2XLiXCTEe7UnA2nR0fmG
RnuJIrI0HUQXVowT0oxoTf4R8LAVQxrI8uMHSKvSz7gNJB2Ahf77MKCxwKXcM8yc
M4kuDpBQCUScSSPSHszCqvSISzwkMAyJ1gVWGv477izN7ywKNr5BYj6ghHHZoBRo
4p+AfOGMbHeHtv78FPI9SC/6J+zSYYpo8Fmlw8INf07gGlJFvXTR8GTJAbtzpf3H
5XL081sV+dRcY3gZWeaVwQjboUZKsxMtJG/ili5LCQT/LKyImnlrFqmtgXxeg+1N
clmNwWH6owv3ox1lfHItMzAuEmSSsKS8lr6uQzWa5mDJQmVYI81y/JE94RtZX8lR
aq3baA5nJPCr/eG3nStPaPivCn3El1WiBdTdY4fyigQ/M2t4b/cWnIB2m8Ytp2ZC
RQXgkgE4nLeyHl+poDjMIXA87dmFuncj/oDlZN9q26YKqUhN5aNiGFsatU0beJSg
7MfjU/Tvwb6BMRg0GtRLjXiIQgWcFbSknpgr5yPb8NELR2dcMHfTaIzeUo+z/kBG
mR6Vq1je0lYj1PEuQkpKdCiOtORYMvo0DzD1Rm1ieuh7numYL3x15G+Nt5NhnV/P
L1Eco7Ge8bUMIq7MWnw415ojFuukshY7Jftbyou0kWNa5+4LkvbK7yjr4J0XSFdE
fz/3gaINHwwOiRWz39iMmQ1dEQ/kBCZfIihLGOuJ5hf218OC+c3kN8C3G784TbBk
+X6GdWIiFkQ9kU9RuC1yGoziVrFChlLizvUiacjG5XgXcWajVBkoZiaa1WjGr+K+
rYFztdbB4R6/+2XEhr7rHT6VqiiPy54JIMMb5ysTsYti2t2+Ps+hRDW22+WoXWyt
hr+XmsO9RmqHVewj2THsBFLz5deDECiXJHvXZqMKRUD9J//h0zxJwHdRiMTu952K
wus0HqKzr+K11X7TxlJ1cOj+V+53P/P0v+A5SyogQpMcaxaN/6LkErFxwSSo21qC
WQ73wikffc8Zu2qiGUKem+/giUA/YlzTmzuFbXoWf6Qq70rw9dn7iryA21MQZO4X
fZzZrdlhysiiXq7vLEtsV3aJt8B/4+sy7Gh5MUcetb219a03Q4YUfEd1dzfm+Fql
rwZwC8sXTX37k91IAJCaGuiZv6gkkDWI0DqwU0aTyDHkwwR3Plu73YiILBRX0EXT
9J9LraOX0Bpwz3UvljD/VcM0CU4SwTvKwr1IHLPUqTFKwhHLVm0s597l8s7IsFvN
91HFVOEU2JUNpEHw0ZI6z8mHRAE6D96w9/5/7oABEH5x/Tqb5yQjHyHnlPyeN+pF
NVz7lpNussFfDkPG0NjNW3CoXZNaFj+42SNBFoa19ibSV37tKMZnLYglb/vnt6gS
Cvo/jm98XhqjNA2vzveI76fOSV2+2aYhfLA2RW3ZvKsn1wUUav9L1jrK2DnCTMTy
DaQX3E78c7Xv/vu+hPqcwDlQOQ0iGwltEExUPa6T4vidOUJcOzb+mZ4K/strG8tJ
mbCeu12zwHXRufjBFxinlhYZLmQ8C6y2/ZL82Vhc3ZiHqspENJ4Nm0OMryWgfYbd
7qX/mc9iCs75WzwlHLO7PnVjtTvIhwp8Fpwqbh/zfvGfQH7ar7rqp0LtBteUSEDQ
8UJ880DMq3FIglp/2zNCJg+WnMq24zW2Os8Y7lbGzL0MFZWQ18Q14cKuJP3vWHuf
/vjnyvX2p3fn1NFP8bb0B7m9mgo0AVfAFU+Z4qzLQcNPJxsH5HQL9ZxniX8m0YLd
g50QD20WkUmhoHBN8uejTgPB1aVeLuux3dgnnCC0HaUihXZpE44N/Z3rpDynPPxY
/9JDDlz4VzVfKTzg3VCgUYWU/OkcJmwJBBwReU9zZ4sme2PDkSaR5oHbvhm1aZYD
wG7sSBqN+7bOKSFNdSttmF3/o1CX/M+nGmSyPSml3KijnA/OxXLa46DU2a3mYHkB
TmSPjKNO77ZX1WKNFqRl+F7Ftn8DlI/3vlXKLGb32m6kYB9G56SShA8EiDQMVzBl
HmoaJk7JM9qKOKNHR69MPb7kfRdr5dmHE8jxc6rc7zaduGtFeUcKMXzpRzpyP272
mKEdAuD2vJW6VeGSI0a+APSQ/MoBcyRA24mc7+kBNZzb7gZe8ts+dHTEN47xbD12
XDuY6LrGYM8xC2BMtw4xj72GpOJQYFo3D+Of50OAeZYHxzyi+Iy71RCXgFWQZ9Pz
awkd2aPowHP9Wm4AeKMYapXVY5+d2n2CR3Hpx1OuzmniJ9pjDlfGlJfAOFTF0nUS
W2yP1HmbY9UfjWiSmXZ0JnSdwYkXHnACkog6qctINb8RUVBVXGbe8yVSwMDOZRJH
QEHh8LwneEmgNBTkK4uwAYjjql8Dd5NI303zZJFBrWtm76NhbXO9i01dh5VQ1slN
KG6vq2bU1Rff+cBj7AiYJxyBY24WuuWkdGx+GvQPTUIY4dMeimyiNelZzvCQsFo7
5EtNSg/weZRoJVH7Uu3rhX246B6jmz8WAOto3c7nVOT9r+kkOyd7/h2IP/FDbXoe
YnZrA9jRBLXVFSlb0AMCLceFWGqYY0AYvXb4kYs+dMVd+X7fEsW366xWBDl/SGAM
wJPEngSgoiAa/nc/W5BHLIqjVjSm3JkDZzl/jn2tliM5JU7c/NQStFXfHNVWTwI2
fe20V2cZ7HtcbhoNWxpWdtHyHU3FeUpAeamaYsHALwsvlQuz51XAXEyiu0EK6fuF
Ld9B8+ydu5Q3ASY33T3s3OAQDjMjaooDzfetzHEscg9gctHt4zdmtFTaYYMfFw8u
8DGvKhgnDZFqQ9e5P/KCS85KIHLW/82jug0vIGnwTAVbbLr2CRHsEdIxERt5VtDC
TXVCFFGiTq6WQ2PhJAwTb87GP/+e1IEyCk8nOVrb5mQa/ROpLVCJN1kWjKR/C04Y
89qkQllTU7/27ooXDkJkv2Ry/wNF4Pkg51suctfvsgWviRdItLRdLpEsWWvDxvc5
sqLkA26HI7EBCp7k5etSnoVEXEOPU1YfeXm/hdugFg+94qke1LPC+rnV0diafDX6
AZXAQSqM7IBVM+9gc092heFf3PdsswufOtdvpateqWSLXYf2KfXgLKn2DvYnF31U
n7PWqgLs8xtBGiUs25xBaqcVTyPDyiLyHJBDvBoo68rrT1qDVUK1Fn4WBqcSect+
K7yKdQh4Kkyo1ck8eHNvXyn6xOkoY1DmSi3hArl/HWSgdDETkolFwfuxuWjbOBiU
WeADQvQPJO0UIE7YJKz+MMU7CUOuqX8aGcPNh650MqD03C9CGN5121av+i+YQYDX
2gvVIdzuGJrj5PA7q07/4XTnd6BHS1680aH0sPsXdPtMdF83f6NEdkbXbGlGUufR
7FXNuFi0I6IVHhZVhi8BPP3S61HRgxCl19R46HYjeTod1glRVfQeenufG6WjuXB9
DIAZa+TimBUpKTNsYZ8IS8Abc+CTH+uoNoRNLTJb3LRxc7HjsrnYbq0IdWzi6TKK
rvXdP95XUmIYabhCd72QESaFxqeG7P7gQXGgWtxenZc7Z+hyynexijAYKuNjuGCe
U5QwQWaJqIpqJ2uU8MwAyGW45WPEt6xpLDViJ+kQ5YJ80QLHvoUS21SPXXJ7TyQF
AtnX6XaBO9S2kdTnpWxoK/3nE9Y22GJVzicVk4phJoRYbudtIdXH4al3nTqjT59v
4DPMBut6B5yqYteaOWe0a53SxZRrTCnuy5wi+m7XN/QQBPhI/jEYy9HuArNky6bA
apK8smuCvIpYfrC69v0Vve+S9yoJ4anK+zqpNVBhx9mMf3C5sxiVJLOSVPvXrFcZ
1cPNqr3nbQAm9V5D0Bg5yb/A+BOfBuU4jqYRUOnI/5cgDaBUsUSImNB3dEgzrxVm
4jR2CZn3jeNAzEXeA5pCC1MXu26sx2g4eUOz647ShKE6H8SWbp24kFpI5yjLSqhA
+MiGw4WYZCKoMzpUp0SliCfE1g7ttlboBpsaECNo4DvbAvyRUiLFRVOOp5nyXK/A
76eevC0YWG3GoGdRHmcyv07GdCG+adtXLDemsUsT8YCYeZ+VC/uBSq7wMF8asg//
5h8kBaWXA4s/3X2Jrs3qCiobQuyhVBLtprseHp1m7uHn0HLeQN52l+B52ofxt1a4
Uero50cVoe51LVycFnyA++ojywVWjllX97edIbwGf3XWx6gPoCQhM6HNVe0Ulfoe
QuP6NcC9EHEylWNlMH/CcxO97VLfoyrGk/AV8rR/rSKzzFXTbSESXt2AoEC+ma/w
VjhUem6kECNHqRqCm63Maz9iIOFldBGzR72Cdt034t8h5G8D+mDH8W4w++yfqXRx
pWvK0LvdFL1DGtJ9HWrIAaNeRrSnPUMbSd2+TeZB/oAuyi0xBRIHPezkrdMFa0zt
dn+IK91OqEJ2O2HkDvl8JqvN0uqkWs73LdsgHiamyJsDFyUm7gO6mFd4Q8+m95kK
RSH99We8SPOut2O5JVwku9bRKp1iSPmBNLpnS99MD9ApkoUG6WcxUy2HZ7e5YRhV
SlfSmPu+eDbI1QJUHzPueOEsdfrZfwGJgI+TKrQmdRMKEsxJZprajQXDA5s6a5P0
ptDcKHLGDv7fVdvfjDd+RPIrlpiHhxJvk96v79oRylAawMVkEbJso8VXlBiQoe/W
Q+7ERd6mik6ilBOU5DiHIf2OrpUjUhovCGBdUfh5SUzOyDxqUJryrvybNbL4n0cp
AFaeZmUGKIQcOH1lTeAswWHMZVkv0GcHGdUes2M8VrlvlMZrg+cAXc8VotY1G34G
B5WJQh285ics5A6faMM71mJtQqqvYBvgeR6eoLTQso2KmitlgZ0Yo15P9mSipac3
XDUHUJw1IOyaB03T1YFk+1f+xsSbY68oBoiwNcbTTMs7k5QRMHMNUhRje1N2Ftpp
WmNkB30BbSy7JuO/CdaH9fv58OFNcqgqeuzk4+veUgVtGlrlioAdqFpI+m+nfXNp
s6Nc2JRAUhI4F7eBTKPvsXp1xAch4zgLOmfVJ9B/O/ZDyC/RqBtaeDh4SFkTRtmA
OLwHXxhNCEE6jsbyc2ixyqd8Tpq8M9NMiH8Ds+/kYA0H/Kx5V1q8FnARXftVszkD
lYWmK/reW/ZaYtuH5gXzG+dsH35wBXm2W9Vibv/jAN5Zrf1hPKRJdy3fF5WL3vXB
1DG3TDvit5cNNOMBS2UxQIfc7wrHEibL4qyt7JbApWskXvy53Hvx7g2MuiNdWuif
PtLYm+rwAPAMyjksN/iTE32SnOsx0d+BaRhZvO6nsFvtukfkblMNog5+v4W+FL/P
4mt0LHdlKrPhB2hmEX0Gk1d6/isN1C9nuR0mk0hBTws6B2dNyPNoNELU31xwIiTc
Hz9IFD7qaIMwLJHQBVcax2LNTUlxurJiLEdDthjwu4PojAIPZZ+IiMNka8LuJCp4
O+mFqppSkRVEDOW9LXmxboQtwsp02T4PGPgCQqkfNKhYXWOjxx/r8oPckLSZi0pL
yYE/q1RSc90/et+FfwrH1JyVxOe6dpfq38Je4QkRR3V6GI4y+ufSk0iY6RAaa+or
gs3q/dnlC+u9PDynIa03HefRY2sLXk9v4GM9FcZMs/Qo2w7b02RwirmfqfNDPIcl
3tk7hqs0XD86a0CK1rADiB225wo6qCe+K7fK4/RtFLnsNURRpgbxH/c8+hh0wo8R
MMWvkDWmgGu2Cw1dxa+GlvOWmArCMCrWIGKCoChp7QMf+E8R3JeZ5L8QmKN87nnV
lyqmDlQ73Ry5jG4tCQbzW42R7GYSSSYKCkQ9lN0PkIfPGbLMDav3H5K3BZ2FBG9e
rSvvzyvQaL3FiGEkbAYMLrLC9KmX3adUkQh//cCLvaOP5lsSzRRU3q/XZBkZFfOO
1/y4gLd1QMCGg9rLu3ScEG512j/i/GcQ9Tr6VpylzVnbY6VIIQ4+8uMlDrogVutx
/jE65DWsg9bRkmfFL/25PRGbON8HJGwgXv+shLSeWKS5PFEejOisb9LhUNiSA38o
k6aMMnWEzlhOFQiRrN7Kt+GeXpAZ+50SWJWYmOSwIYxx0amUo3yWkJzGys6oxhou
XeSYeJztO2BySsLh3rlRazHW9KeyElSwHT6rn/+0SLKeJYcSUcNe/KiptNe9RyoI
ILhsDk1r07p70eS19DSfyC2B4Wfs5curY5/eDy043vUscmIdUKB2PDWQbj+yhTPJ
y4e4Au7yaNUMVPzxEiBK4F29NbrSZH6InTkRMkb7owckaGc6/rXsK4GDkXAALAho
7OmjWt+smLYZjKyE4XicIOX2G6JaKf3sqIXPLayyZQ2t1q0JoJ3OZ+ZZZFmUsD5w
iWGPbI7skVWtGHr4oM832WbyWPTk0Q043G8VH6aqLT/WPZiwny9V5sCtCegarmSO
JwvHRgzr+Ap1xun5km1GrrjHgHTzcHR0shnGm5uIzh8Wcuczr1/+lj85IQEuPLcN
WQxYUf1EmNZu5Gx2iqpdsas63Rxqn3AtPGrgA1SDt7wkT3Ss0QXtLeNdTy8URCbl
i5wnDHBVGEZw9FkjhNWU9KzmVzp+IetXmku43qYH/ixofmCKD3g/qBJ4gapfw5pQ
6i+V0096KR8/HGo1kAJUdzHIPcnVdhl6PhTfJmS/m6fqS/FoNaS3U2A3N1IyFAif
i4NnpsVkuK99fSJ8ze5ik2IZUvzs7sicFlw9RN97QRMUg+zlPS1e0ydEIro3TSMt
KQda+JX/SribrhYBpBxqIoV+RAhP38mtpz1N24BP+rsgSk7cbyMHzGHZtfjiGJoI
wdkXXqxMH6UX3LglcIi0xZ4GwG1xKC1eFxHt/qINNUbXkisnxJqWrTOqeGerlxa1
oCsG1SZWZAu/nHHkqn31CsQWjIT5cml1nKT53wSPomMmqRvYb/PfQlPuffb5YKWV
3g5E9lXzeABXM+F4T9EjIO3+5PzzgfCKgWR7NxcbGHllP5NTZy8M1KtiWAiW2LBb
tHFFPCJe8cl8wYRTS9XpGSZqzq3gmueT69BlxVGaYshvToc4zSR8a4fneAG/FYhJ
3+g62O6fRJVnqxuL26hXL414P65qUrPov8ynrMT399oy7jXWbYdOJsakoQrg4pyi
HMhCfepFIcWC8o63PuF0sPE7PfV6y7KfYfRQGYAt6uDHHwqFK3Q1VORMrg2tFo2Z
joZ8FsJzTy1wOLDsQqopPrtc9NSCzdwJMRyW9lVbMsqHrVW3/WuUPEoAWxNqG3Ii
MAazsnA/a5waHTnzZMLMukhqCT96cxdB6ynvxD0cZMEYdh8alAWYZQCCZDjX6aqe
WcnVAQ/eaNcQXJKWwbmn+PU0mZsvpnohELxckGRxamRkOhNMml6XOUlenhHL3D7j
BO5O8Bv1y7iyWG2UnISiwKN9okDAiukU/ByW8rOZtKQYHk5bJkVtJy/rSrA74SIx
GpCib9VSkaKscRNnzchYgX8WNm+jwOAwz5rvpDlTdPTaOjeZQdMewzl+i0TOmbyW
UxIo8guL3uwed7PVA14DNYhd1e4/j1cH7tcSmtBj+3n1OnCACwFTqmWcMChUOYr8
Pd3buDN7hDUYfpNYVJ9EwP0P4fsAfleCIqv8reP6BEg9oCxK3L7sUXZjiE8MH/wk
378eWd1R93gxEf1vdE3AsuLEaW3mdwKfV40XsDE6g9hZa1NUsedbZp3msdNJKukV
5K15bTy66mZmc/lONKy0smU16Q9YPNnaMpFv4mFVQPjYxHQ3niy8yQLqpReMg/sb
5IGY1jRtWUAMGm5W6aSI/K4uhj/33QmdjR+quOmZknBcXg83vEPt0cTQbkdE3cwF
giL429Wkn8dfq/fcA99+9CiQezBbZeZagnCeimvW70ELiHIEGiXPD5zEmqzUukb3
U477wLa40Ahi21C4UhXeekhob/ORZ0GyDgE96/P1dxarLvBkiTBaeZqmQB+NmPr2
Oes81ljmynB2O+oKU+Hvdedg6RmXNZBW5rjh5gdNVFvffu8R9KJu9pqnBNJ9oxQ0
RSv6LYxJCSI3f9erV7bS8Jz9gjyzRNXZsXF5aEexCX2B5V03bJhi7qUdlPKQIBjM
cq0LzaqdWTGA8CdeF7xOJYQ6job3sANgkhHwSP84NvReGY1LN4bpxE2ohos1auJV
I8nJKnw3A0hgMejL8sWjvevxdz2z9SFFaJxI8B5rfg9jt/lJF/DgKKFlW4ezIHeb
II2F1ejP/glsMR6nh4Sr6Z+1tl7sjB7mPtFZngXh0XNcajLfLxqvkZzt2FxE8yJ4
x14+gxhnEN4Neby6Ga3hCfBjzAKmUuwtY472oa0m8DOMUTgVq9JBJqkG5HvlVnlk
aKfPsev9duuwSP+AD4wRPUjbDs6D/fEugmEIyi/AXvcZNGRXIRgB/7FJUX9orbgj
s+T/Nf0LiZe1LbeFRH5ddX/OhmmoreABQvn+1rOwPxV2n0FwkhxaWBmvHhfWpJFJ
o0D+VfKAZ3JnoY4/3+QMu2/NPXzRY43LEayr6Izw9YO6psh5wScp6Kknpr40DEML
ia0DLoGtrnG9l4i7uMFw6bp0mlao4Fw6jC7sBRO9pfC4KI614EBqR6YkH7A621TG
+u3jH1IjXhYdtxEl6SftrkJ+8NRCRkIK0agnB5fNU2RDAthtWlvltV/oTFuwE+NL
Ydf/BIEWE2+2A6x895FeK4TD6dtr8Os4uqaumhaBQ87wxJYd7CRVjQdGVLrJj5aQ
OQzBpJXvg/PQu8Kbx5oKY/QdzPYIHl0I2oEMsh1QXCg3pVxoWDYxq6fj6wDPcmK+
SpLydFZqy2ba5JnJqYCYdchYuaR1qENpXPi41Sz9fryu5FXYPaVSLMLEWqwRlZpK
0SiTMa4sjD+CTJKwat1X/7Xx3zzV5S31yZXj3TUJeSraCA9hhVx9KPSkFtHta+T6
sWvutiUMG8d1ZzvqPSzrSKQR71ID7MLfhS8XFZp4e6zewDRLmsX6M39qh3h60BKM
3TEXDx+uFC93gnWrXcpCPvd04TpHVE6xM9DqShRamf3aJuER75yy0Qo6nnSSatY5
gtMUFkIqlbRiKINglGeMjecPxM5hPfacbTDZsPnuloLpJBnLxTVeq2mN1GBPGW5o
pOw3UX1gpS/lTm45ISJ0NW6dcgJoARU1HR8Xkw+cn4lEBJm6Zff0z6gIEzYDo2k2
nZ3MvMna+mELSrLO2e+liTZ/Gkb0WfIi3fXaWBVOoQiD8oVokFAXWrjPyBhV7TRD
sirKIOh7Qv5tIu7d+h1mk9IwZkcoH9YtbdTZBVLIUT+IuQNQfa2eUt43fAG3Xclv
/eUmn1fnm5P2TgwmIatmyG0pgOXAPtjyrcIkTleEvJ1+9cDLIvUUzkJxwwnZnxiF
VR4Rb1LU24hJtOPGR3az5qlsW3ofGvK4qzYw1lzO2J3qxKLrmYVVbpDNlglkwu4p
r9gKm2jtWI3BERM1xJ4VBIyzAWnIuWnDpmVYWjksvGV8zITbDqgEA6X7s6v4rK87
3FrJqfL7sw5naE5KKy9RYaw3szCKs6c5M7aPImkDnxJHKNAucJTCyx3pfrFZCT5I
MwJ1Y17cGuCeuBYd1PtjDeysvos+lxR7UFUL/Jvxp1FHy/jKyr1wA01Q6bN+1Ghn
nW1seoniwEUJ4LwqVl2dAe18GzVubXy7KXrQov4QQjFprg7ZJmHdI5ZNj1nRV5uK
cChI8+L97Rv1aukZnwYw2dHLA5o9uwpkIxuG7YcBJPizP0SskC4bOUTAo0tL2RWx
ur8HSr+XdkkyRhfxXMGcYaZW71BPSTm+CCjX9+RGtU5Ftks9UfhLOD80qOHHIxwV
ztFmrvzjvj04j9NB52lMkXCJEf70oY3PYuUgjJxc2g/x5RVuVNxwD9ad2UR0oiJo
TwpfwvH+yaDIbaiQDWRpP8c7iHzPGI2edXqTWGe6WM2ulVBPR5G8nkKCz7r5L/Gk
2RNXBZDmk8l0UiXkePeuc4CT5vRgsrQc1KqC7jrTYkazFwQ+DfOP42vCVZ+qzQxS
4ofKP6P2gvLHAVcF+HBT4MFWXpPhaYsCyPBMV1bQiTVfCp68rBJ7PSj122karsZf
S+uMaZwzwm5n+d/7gwKq7eVVD94YIjlqDANi7vtWy3ULZkVXshEyjLE+/Ca/cIOD
g3y8BlzIZC8moom3v+wVmseEMi+FoB61vM4tzWIsUiQ24nnnvK2DOYNsNI0toqtQ
0uYAzWdCDySl13jrPLm/n6F8RVkyA9+vk3NJFxM+nu2efIOapn50U2Ahmh02nUma
udR69oc8peyzAkOnJs0Dgm8Nq320V+dj5OnKH3c7ZY8yOfKRf11uFRYItXbE5XqA
j9aTMAYFPwiXkqQW5rApcDSsKjaqui2RJcH6aigexFd4Zwi7l7+mIALeANdSA31v
4ADErX9wpgA6u/QxJag9Z8kxtPNZliXUeFnyUL+jD4wbYc5ZJHRTfEiVCR7r5z/I
ZkFjwOxpsH28JXExPksXzX97OlpWPrNSEXN6/4fhryFb/fWsmyY4nDTy9vLaeak9
uLI0GWiJZNqDnm2rzrMK+QxaiEd4k3a/a4f4RpNgU86d7GEuM8NjRseutQxND+5w
mRm4y3xdC6C/ykYCcdB4v8zGaP+ky6kuI5hH3A5kYV2XwlKNksQmJSVVhaqagsWj
CQrQtTPOqVSotIDLA0ORcggRbMzsGjgeosHY83aXbzvIp7ZfmtuRbiD+c2Z1/srJ
xOXXjmyM+aUzamw/plQpUvb1ErfCUnmsN3PK7mJh1kT1jO90NhK85mXqg7G0p9GN
zN56KRbnwyQlz0Je2q67+Q0lTYX7zBVsAluSJPEq3GP3RwkKtmMBHL1iYr7AKAcT
BsLkRwbi45b3E1Wu2pREaUUbm4ykWG8t+Zwgjd/CENSSnr0P3Toaha5MhWLMTHkT
sogJHikpOw9NtN7Jg2+v6sUyqAf0rEsIQlZ3go6YmXfhr+FtR3crqEzezf15MXId
jwEAfr+geQeCy3pzPRzKAQskoEMf5IEg8oijsVf4membHwbeaQkF67I6ZiRsg7kX
j0ko1zK2Z7vAYjHaOmSmaJl1jl+HSKa7eQngdDxw+lDY6yQQaLCVUMza7KHfP5lY
FX7/KxjH4EnDHqR9jd7T8Pym5sPm2gGQKfKpki5047Xm+x5x2pPL1PLEYyTjJhkY
aaJzRxoPBzv//3VzvBNASNcb4fP5P+k2+rhfR6ToP7jZ69aqB0LlUIws527f3k3q
G1hB8M7BXFAbGsl3aDL03VXQCFb15JRMPPhjTCuXVsc3qE2KKYwqMm9j6fATSI6f
AdDeSKsI0yIQhRTXzcaQDOtjsPe+1XT8NDmJPV+VbfU=
`protect end_protected