`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12160 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRpcw2zQDHRgJxPf7yaQH79KRMqfN1CY396i18KXVzLP3
AtV8fZkBIM0v525LE4mEt9+6ozD0UU/UcBYn4J96vibR6dhDiKcTn4B5o9kpsOxw
ioeMLGB5V05cY59psY7TKXznLqx+u6EDysfzP0FIRSZOcnGWbBlWUXQZWHkFzjc3
xKicfDuj0E0D5mMhWEaHnQ7QCa9cUJIoJzHNiSpb/pL9Y7U048moSa1wkWbFngG3
DijkalfTVCDmSfG1Yp+PGyH1Wd1cUDyOeSJI+ezKkt1QFKAFaQeZLj73vYUCo2Fu
r7lh7DlsWWF4vxlad2nmIMxz1FOjUR2KmuSYJS9pdEnu0UL/qHLv9a4wMvgX5EAX
ScMuR8109K5UBwncVksLhvGJXcnSRJdD/vQbNjnzBXlHIvOcZcyXbkcuAktrYjOe
XWAvYXWVcAJk3qJfyEVlTe/WIs/lgaIT/qXhBeGB8G6acSl9Ixht4H8ImcRN+dgc
EtyDYu9CXwffULcMDNBbEzzdEcktVHSXcOvdHNKGtd8SXlNvd3/c1ZTYAfcIuMaP
YJUv5TYDVJwcTm2hstpzYy/ZlhEMyuRzKmDc2k+K9t32PRYKkaKMHBwwcE8E8vE2
/n6B3+v3rfeHnzwmk3JFdBxO5NHs7ZziV+ivQkU6MMIzcYDC0QZDIjck1YLF/cmm
1+suhQp1E1ivqWrU8IhqI6lVD7NVd5Vv63erdfIjMtqrs3LQyC40aCbdO/iE9DiE
WvQxjoZsipiyh7IPH1ph37Wb7H0dEzYo/O2pA+TF8z84BZc81HNPFSAig5vmWmeq
vmyg7SdN2Tbdlrxt7Kg3sZJP9tvS8gvIa1BQgz9WXun8/1Xu6yeUc6x/TUrd9o87
yIFu8w8XwGs3Y5HfRsCAgQlSfVmRAJRI1xqooGa87hm9wU4VoUA+uu2L5PbZMO0z
/P8E0eTvS3zT7vqsLAoTnX6C18Zn+glyu93UVaEMhDdaUZycv67U26D5CKX+aeVV
NkGqvQJzVwgOcCNpjeTOAnkd3mv+YGkPFKu0RQscC+ZLFkT0Mqk8HV/mwABb4fQE
gAxjBHZqLI/H/jar0kygGmjZVzduwbsxGpTcYN912pO6lKif31fn838RQSLO25Ne
Dty4gFztIeczU2krWfgBhs55pGE93/rfCZqB+URxbQgop901j70t4Ht2hk7eWAjf
a68oTGQe2ysExs7qIn6B/cKE1WIYTPINo3XPedWoL7jxS1Yuph5UEdQDOALRqNQu
ikpK9ZgfdSc7IqajOgHPb+dH01kClcZ0qrUDvL3SZqKNpDIMg8Hup+c+Xj6ri/U9
+1TwekEO03UvZQdo5+9+8kqDVW7nw45vuLnp2LuS71xXJwF5rY6vc/lhT3HPnZh0
8VzGzDDaJQ5PSekCXLZh3PDSPe5rKCq6OhRKryykduPGwo7c62tpQWNqANYGmy64
+phDUea7q67x+jyqQMu9UfKl+q4TSl+3GSaooGulP+SX2KgTlGXdpnNPDm7lTGaH
ohWCrLz6VELy1L07HiRr4ge1eQSlS12pdxqXDEx2/Da/2kl0DwarBZboes4g3RU+
PF3WoSXRdy8quk6mDFwjeideEWBsrF2ULQ2NX+xH2pwMMIHMBYi09p6GGCLJpRZj
ngX6XgP7iIeNB0kUa1gJMYq4mYX2xbhr0cT2lhaICKuhR3Z4DztVBLFAT7xPF/2D
GpsTAMYkg8N3FZ0FxkqlvrKDqGB24/X0U9MOry9+/VBDimHSczFxRVe0p1SGGo87
vjL1S1sI9LEFXzgCrR5YbEaeqjWbi0UnfR+iK6EBL7jCchdKFJDpYqy2/qsl/q+V
rAsKiYQDX6E+eryNoEtB1z73rCwE0vZ2UKelWyGBXYOozov6ux6Eg9zcd2Ha5WwH
3eXJ7ymVmTudzo5X8QX7uDK7BOom7Q8bQRbnh+wRoBaEXl2RKfAADvPdvpULDEj6
tJz20DcoGb+JXVOEjHhZQENYB0ACBVQMXOAKsoJMomNRvMTqyFhcXIFgt7iOd5aE
2N7ImRoJIIlS4ICcXWT1QGyuPRbraxti+faTKtw0gNeMbBrij7ci9Q0DBQWhHXOF
cGB2bZ9qtBCj4NMwAO0VubIytfosWbkU3fidTqvCTOu2ChAfYgOHerRn6rQSGKwg
j7ybROy64gYRJjDYPCCkcCT4GJH8Cn6vI+KmRkgDrW+D80NeTnFh15EimC8ZnqBE
Pt9tY2j3Z/CsoXSxSDVbYNWDMlheUQj4DaWsDDTw90GI28KME8XzkJQKiF4Uyvqh
/Ejue/ktfdgIURHiU1EXQx72poYdpNxf4MRJ1F/F5gWkaLMcAYgJVNO3w34DP92w
n2Xnfr7gZCgrVTMFEjjDM//ULqcoC4ivMlYkdzGr8ofkMOaBlyHyf2gjWkI9/zAi
d0SVPd+rTun+SMGLkqJGtLlCjSbNPjQvfoLd790NQbnheVWCLjvNh41whn5yNIhN
xUZitJZfCXLoz3xrgIdOxU+bapYjoisO+iPxMpwhFF9Ng3kX58wpZ9biTqOc9HWE
Xo43Hkb523bZ+dLzrEJDhKJpvxvbFJ2Sf/Uu0JL6/ULmIVTcH+xNHXJmLDCzVYDC
8J888OwI8Cyl94BrHS/i2FGCMDBl7CPOw4Xk9apByXIhGXLXLjRMsvDcUC0Pxuy7
h4WS68ixoc5xU0mTtw//kgX+cnj+CwS1qUN5C6mp59diiDc2hAVfat7XoIcNxW5L
Tg3nylVTXv8GMlXZsh3fec53UXWQ2YaVg5gtyIwR8GZKOwH1pp6zuJrCf0KR/NFe
+xSeaktPizF7CCDVE+rg3U2j/aJpoD2Giluf6OztVw62QcatSNwa14g+bnBIMG5m
tz/77/yTBGn64xe24jOB+W1TXcuiMeltxai780hfSf1SNUGJttZjB2wMRqprapRf
cBZ0XSX4oRH7rWwn3MEWHDloIHwO+62EPQUmcIOe1ifMLKmR1knihyBpC9opYC8j
ICtMnfaK90y/Hb26b5+Ghpu6W5O3X+5SWFKlFmB0WJIOlzca3rNxTRrq6aEoPNDv
l/xwxipctmQ7J00AsC+MVW5/6F3VjD9bULr0UvLDAoOCqwE9ucB0aIM36KU+oFPr
1Cei0v9f1KdWxQELkHdhbdHr3d/W0TJLk7+s9EonKs73Z0TZ88ZgRsjZfFHVCKoC
JC4ZAyyzqhh2cdmn5Q+Np9eZL1jIg51BzS3k8Sx/ahWjB7K+OHuFtMH66Ngg8X2s
/oMWnpyeX8IFsN9ndceyiFVTTyeh+wmVYJDGpc8zz93bV5TQ9NGYAAneARWvqw/+
Ng+BC2Bohx6X6EvcYarwunTQ7CaAWxQBzpjY5ud7F3WmJN03YU0h1WyDqAtets/Z
e8GjmwmRTW5fI0eEGGkwdrBtJws3HxlwAni0g4zP+ThCxPYXpYJWthZoVMHCrJVk
TBM04kiKUk/zSQpr+u8pGKEPPD08Pt5qYKXKMeoA6DBGyr2cRRsfvH3Tvx+/U6H4
2NGiI5Kp54iAJzGUaqdw4aeuKGeGz/r8rMZcI/faI8+lBJAPW7j2Iijg/A1lp7dg
IILyrpm9/si0aqJvGLMjoDlVIJ6DUY90uOpPaM6dkvSbmPMc/4RYie9x3aLC1zYu
9DIwBSTsXwJTquG8XDkM9NX9R/DawOgJtN/tB7GfawcBiklbIAi9Nh+Isl1wjejp
jYGRKg+CZKnLNKigZBmMojs7LIOdD1xPYHh7q+zf1u7Gr9tl9eikXw6A5AeSq23e
NtUsEtQsLV/zR1S4MZrH/LJOh7ny3tLIcJyxTZnEJCopnqOGRgQ2oAjrGJBa/VA+
KlsEIPwvgIeP12CO1WreEUQQ/5sM+TKLdqwgDYMuUfJL8B/mLBcGIAr1ATA+YYsR
1ZF78QWDPPsKNETxFnYdqx3C1v+fcAfAPWF1JM9ViJ2QTWDAYR/Nu2T3ZTDf3PFk
2mYKnN8RxZVgcymHaFm9Qmeul+rkhX1tdCA6vBD1XF8FHNtFyROKXFnD4zKB048N
wpz6Lcpf0pz5xhMYeupr2GLBIbtoRAJArFwtLa7GDuA9t6KsoNO4hzpbUQZehFjX
yhnP0hwLZioixq5ntREJRAL1DhZb1aMVP6A9im/i1Jp69ODhcrADL0FVPISug7QJ
zuXwzldp2pcIf2drnaQUwpXwsiWLKXDI7eMCXQ4LqP3tOeE77KYqk0FHMxD7iMhm
2pHuohvfsXv67PKcPrqeC3kNSSgFh093kVPqlcni20JzHBXv012oBKVGHiy2/5Xh
unJ6JVabrqWudmzmBmIhmWvo5ilqz1+NLiUgbizj/6muRqDFmPQTv/3eKP8Vh52f
B/g57l6WAvpDsLUgU2MXq0lDsRFl/O3y2ubEXX/qzsw3og5VrxL3IGzBQ/Lol3z9
XwjdvHVQTgZMWRMsD2AkdSmKeDBvlSE235mLR/1nde/RGqBGyB0HW0lysNyjIdD5
QhByEA3PyIc4u6dL1GOLcKE9Sf19w0gv2Xz3Wrn2kvGtxoQMs5dyaGC17UyHBR+t
tTCSKpqP3+dJxdoO7xPCbaUvU5oPi32/5XwYlA7XhjcAHUSPnVrvLtA6+sQVZijg
YccrX8xgGWdOXSzEE7ltXtmNWiCiJsWcOICBJ0p3RPaxpSw2klY10uOYoPBUOOo/
bTbgTZooPnVTBohlo+0mwI16CghY5U9g7eiq5QlP+f9W9IoIeEP096tdMlvAK1G+
uO96PjD2T6cx86uuIRv0BZozN8Y/zg2DKDzrInvpEZ1KHPJVE1UEvmf9YdmabqxR
Jc9Kfz+HJ0iWlPCxqmYh84KF5TGoDJrY97hfuNQ5RmBjiCMViWovpd2rSOjPv4+T
ncm79gcHX9CqTuViCrQbzKmYW4dSVfrvvL8jLMV79VPBipfzY1bn4sIphmDlt8Tu
NQjjfv+QRUDpU5nSAiPTJlEx5/sLaDn8zvnE29+yFaTXbg1Hg7edYyV2xVpJlXHH
l5N+rN1MZ89gcsWHpSjrpizZCtBR8gub/CxwaI2rxTkApT2Hdej/jVK3L3bUtBK2
FFW/N+zH7f/I4ZZKJrT61ZoclbxmVxBxmtsMoSq53hgntY7BF7W1UhaSsmQ1oyEV
TssvZmYxzxYEfy3F1AvgyAqSKsIQpCmEQVDHPqN65onZdKTbQlkcgGqxwRvUhhGD
rxBKb1rT2aQZjbp65sLYelhCTUUKdGne73TdB5lz7jRlrC41QUuv7W133MuRvY+U
7u8R2+B9tnaIh38MmwD/NItRRkTIo0nJ/n+ehDtoZ6Tqq9GVPhfjmp/AOoyatoer
Q+DF0Zl7nUzhlV0sw6PUXgpCMRbxHpwAHRtUozSoxvPiEW6zql7f2r45RnTGBfhL
WmrT4DuKzozyafky5LifeF+VyXpnfzZbRDAbSLuYZyFmaiHVP0tnBNqoSB8vWgMs
Wwhd9fIBnWGBiZpIt20h7Skvra53Psi4qgdKfAAPSnN3im8QRLVwQZUJox8PVnlE
hdPhB6HE7dJLLljYCwMNwWbq2RlLUTtVq0rANuYtzDzdmPIAVYX5KhvmoOPv9yVC
MljWqe9a+7qKfjddMIEu07UMakbcW+qUqs6IPEb3oMh7Id5QEHpwVHYw0hxxjaAc
MWJ/zFTjcHihfmfLWF1VFe5xzsWvUYIbUxR/tMRJQjnJ0YtKrImDKUQxJz48WLKg
XNwloSYJxk1CDVl4pKTyQqSbG6sEwolax5qw3yMAnQCD/SvqVRy1ayCEGoOrH9+K
LesoDWvn2fwoSH03kjMqScRe0i+VWF2rpo56DIFGT9bSEAfZyhavNAlrdrYsz6is
qvByCn3wKYb8fZZQ0tplWisCwildrh4dvIP2+DiTXNII/i/w7uuJ5lDaWcf+igLk
DSqq6sOqIT9rJnMYfVJObkBr1c6LAxzod5SgcruL5MIamKX/YU7URG4tP082p5R1
vOelHjwDvU1OOWz5Jp95AK9cWx1ZR5fwTah1jrbhfsPYHPeWlma8xigp2IEHRwrA
kBI+8bixxm+V+AQ0JauZGnKbH2vH5+6ZNESX4zOSVJg1xqLX5wL8TGvTXgR8D1QQ
FXy8sBOEuWGtjGvaEpSVG3rNPQuyrtd5BTkk3s6jCGCVD1MX4egirJkVb+aUTbDq
MlPIebmvywFgKC0ZSu31SQWyrKlvP0ogezLTaMK9DIXkWuIXyNhn99jtWD7uSkmy
aOWM82eq5DRWWm59i3AOtgNZ6TumGq3h0nUwzSoJQz9q75vbYJj5uo9nyuTkZqDw
vLoaWmUI27CEtvEEaP4TSN1mh2wXTAj+5viYTgtVMrCclstf65wK2Jjh2IOY7Ru/
vR0OHYyxkCy0XosJwopduRUxvJG9AxFTwr++1wSGB8V55tsNfcTiUjPH2QIzLb32
soyQqkzs/YSPzVFLQC1M2SScjAsf5uszemVvPXsGVIheEPPw6IUsNewsvXvnKUeQ
1A1Icqbs6qucjHPJSfyGi1Hb8wAjL0WL+nnA9wp08w7RYeCDw7xh9Lf8lqbINoVz
oLhaXAjGaQBGp4Hsw/5mxJsS/tzk2Hk5epV3T/hlY0TontQFoNeTDZxZWmDNz0RU
Fma1ClOi8GZ/Wl/ZuD5kcyj/XQLfV5cdo2blV3Tba4at5r2LgrQ8YSV/bTCJUmyx
ooo1YyTqzVbW+//wkBQjdUi3KHpDmt0dlsjGDMvdEJuTq1B/AtJE098rkNqLr0ZE
j6qB6j5t0ngsvt7OgT8a+MUIv+nXZmx8lkv9WCuB4ZaNf4xCH3yUBOd4OhIn1TGg
PdLtz6jhtOa9FoVdWYRkF8xK1N0df2Jk/DfmaU1zZq3H2cfY/wLQ4rIkkoJIPpyM
POq0xYNcAjOnRBJajjXKOCAX2IRmWfX8A5W1UUJ5czDdEFv2oZSi+bf/dDswa5ym
llidrx/1w2c58i60xE7H5NHmt1r8ll9LibmcAMzgRpqkmTOuPcJlPyDttAZfZzv9
Vg8RLW6oLgzZPZTAvRkbdNhH56ThjdUl09ZEMGvqLqLZ4DY7y61Y0gB3pWoSRl7D
IxynnXLWw8RWStv2VZL+02CxcJj4tpeeZhwRgaOrKGONTGRQRmeDocj7G7vDsB59
dgHAVztVrXx24UHffG7w+BOiKat/5HBrUw81rkQoVwKO+/4D7rfgJ01m2R1iyBJO
immwkIM7rA3CYhtiE3AZAhYHBZNueONwWLXvFQtDLCt/9QMpV12gdToR9gydfln3
vzC/sW3OAgsBicOcGi4SfvCSvt/n+V+/hAezDoraqUf2hSnFtlHhf5K8eImOSzaI
GKcnBBJw2wJNsZvMwV9D/8D4Nx0hzp0r4lZzCJ38r1FOJm0M8a9RVqSQa5rx5eeV
EhzBTR82MLZBbGCNAzbRC9kxi4haP53UEgbJyjBUqsXk7zYqLH1uO6QGtaxkNa4V
OfuPYud6v7GgrCbRBEjTjM7rwCSC96idxeG7zjFo/cPYsIChs6blnGDjgDooGRpS
qmhypSJBChr/xQnhp7c6pqaXeyh4fXeLuieRZuxzkBY6nTe8mc2kBs84aDPil5Wy
fVg3eRx2HyxjEX6h1cPbfsHFOXFEekgVgjAqhWS4zHEvDQFUdf01EBQ2GkqsFcdw
agtU8OpdkI4+iVxvy0YN/18llLqz01mg248UbNpFFnTA19v5YhTpJ8OvS7O2WoZ6
lOz9EtljL4OAWh/XBv4gKGsK+u0lKIowhw5jy5DcEgSqKMg68M3JtnnlW8NUPmCP
S1TfSdVhNB8V+pdd/ElFvqozyaU/XZjhiSv3uB+2bMPMXwSOaRtM+vjplRMCXFCA
S1+soPlUHyilViCMW1cYzWOPjLVIWA8wn+2fc0NKVIIZv9Jx2JGJ5rsIAoS+HGQH
NHwjdU/WdKXJksZ+/AY/3fBqrfio9Iim5Jzd8X0AJ08kMyQ19N4aNJ3oxt1MLCRJ
vV2/ho2VqBVCYxRqQ7raGq3FksNtYScwRPA413rC2HHA7M50CmTGwcsxf8pj9j5w
NGoD1XbvXVTt8MN3G5NaZDkeFOk2NCrbddBsNoEM50IBOUCIntqp21yx5bh/ppk8
cx+zhnYRfuVkcP9UZaGMGdHhOnV7DjpV/YFT+86ZUyt+exgpaG6vsnkz04XB4aFI
YmirQBITozzhl8HkDcJCztCQL26AbBerMxa9csw9b1lwDFvS1Z2E5lPGt2iiJ4s3
5VxB1mx0RzA4mjV4BAJMVHx0LOWR+0o6RD8evj9AvMBLYwC7Vo59MzbAIDTGH3Pc
exXqAefCTX0YtVDI8GpOyHBf0A4VvXVXQEunzX3W+1uVCyQHnDYLXwIVIs1kn0mX
NxweUq400Ntt40Sj6VLnOWGPrbb3LkLs6H9a5b78r2ZIYz8lc4G1xqi68Z8FHy9j
wwOVYPIqly/PR6mabhVUVdTDrWB+XPG4tqDLs0sxiNjh9RQPoasdKtJq+6BP7Pk2
o3grz7DqA6z4t7NNMlmln7SlDwAgCNXx2p5I8SrIYoyEgg3Cwg8BxuWR+F7QFUjQ
XSy4s5UxzMmTYSkxprVy4hjqWIluQQ7u2ROxvg6RD3YXAvSs4ni5Sm5mrDLhBEx8
87aS+TeGiwSq3bAHiOMyWfNgRFfx+Z3Wp9vs1ljKUogNWUGoaUullbCzNsCgKNBl
iN7T7sl43yA+gIqzsMPWC0lyWggIfl13yadqOTTzSdCV4S4MisVt0C5xgURhDYkd
vH0iM0SJCNtBUFViR8YIcML89HeKUKQ8YFPWGgH/OiLqlmpLCLebp72CRgfiVZi9
9hb3FkJY8h7JByktfunfBRaaWaHcAgXy5PFhHj1BnXTF1hmpxN0khg7z+pP+QyFq
feOtNceQW7tpLLZwP5qV1/2enJ4OSRPBx2FOaTapvKmobmYoDIBhH47EZXooWH/C
tRfcconmzzDKyawfjN8HCxleRD+CReGkP9qt3jslJ+FIbCxnpvSM9sPYUZJPfLmV
C1DoDpLMBmqDTe/SJrowKJCkJRlR/dobZ/jmdV2UPvzOrmBaifxCcZC5TnistzlB
gGi679hcA9oO2tOoTBk134qtV3jlg4AqyqFvwnwioddrUSFohEgVzVJ7DW94/3n8
zRo06V2bHemMKRcRgk05tPSufExBDv1+0cxn7e7HKQES7mWswRqz7zag9FkRK3sb
2jUerTGKWyWM8gGWU9+WERnIBJ7zsnBtbYbI6kmj8m+eJSsNoYYz+P4UQ/dWncnv
vYHE8b+Nny+kDqAaOyzxR+iacVaAKp8yMhNilCU+xZO8gAO5JJjynjHPAua0r1Vz
I1rBROgd1HWWbQVDihxXh635Fwetw+ok8ggaX7n9BAP+UyVLym6/Z2cRm3Y/hXH4
183Ut0MLElxB6Oq54FKgX9PjK6YbzZzIuhgRgKBt09COfzH/e4EaBbffX7Wc0YEz
qJU+XqvOn1+hAZGsMyOK2jIO1jVr5NrFlPw8r1Iap3FMsYj0YU+Ksj4bfKW4vHJ6
hZlO2zYnZYZe6zsN8liMI1bFO2Zj9AfY5sk8phRaRt8KGil5dR5xHTbvpovEi+M4
g/6VRYT4MRswbsAFDRVChzRi6JrbuGJjZGaIWsbejM1zn8CypaYA65hoLTJjncmq
zAC8cUxf1iAT9yTkZktVF+6vaQLiAIcd2Xmd+pK0WzEPByynu/QVIcfci47/h0Fc
Js3sEcKn0TlYSL4fJ3uOPlbuy1it0+i48BurLrDDlqOJH7CJOkAai3yhXxr6YTKv
hIpZ/iCesnZYrjkW3YlMKkqPDkSBOgXfGq50IlUa0w9wG3jrlnr2USEzjTWVQFVW
8rZYRvNOTJnlCxSTPWKq/8uh2Q6SElkWJEAi5YhMvZrOxiHHpYvXQGbWpJblD4RH
duwVwYnuq0hrwCaeZYQNCR+BVKYxq0ZDuBWsB+Mi6i07TCfC3NMSP2yr31mtnZxj
bURrgWQEDVKNi2Q+re9Ixy4g5i0J5/ARJWsvH6S0uUzaC0wHuFTzIsr6GXc8ku9K
h1xA8UwZ+eDIUDV7oRYWVYh4RQimHrvKT0iCqqgAQgTuSxisA3o2v7JSW0y9u0L9
rzVGE3mBCFlsPdgBjBSZzLoaVeQyQrMFmUgs6DWJVzI4/QQkyMZn0055BA88Nz1d
E8OyHl+QeuVdq7HK5DaxNwhgy8dYAuP50dOuJHF7fQ8B6yR7JLh40mH7a2wGo5LZ
H7XD+aZfmsBFJG4iLSL3XU59BXmqvHXqBMJZK8nZ5J798h23ZqQqy5aK1MMImCZc
BWoAHFWuou8/O0NrB6nBtmH5jLMF1kDls90odTfVpUFi3F3mynLj958Mru96+4l3
NE8w7Br4a3NJkYn3+FwroXE2MIEaNiOHr1Y9eMV2YZ4ICcgd1v57e1vXXjfTa6tF
UEAhHO/DnRgXggx1Fp15NMB4AgZE0+G2TuWQe0XBBVNiWh0lT906YATM4CxM+4/H
FWoLQjvSzUPT9A8NFd1JdI+9haTgAnwdHucWKN/o+IMnTQmlErt2qwT35Lb3THat
w5l3YoZse86Z6h+93A+wgllcdr4Fzhec6XpgQOIf9+lDS3FQjal47AgSAZWdakH4
lJrtZeeNthoihgp05CCxGlK0kLTW7V/E3K+5bLDd5V2gzdbKeBnqpRxDumiRf/bX
A31AykxdvUrUZPcHLTnw8Q82sXvaEg+nAw+vYMn4/mL+ega95CeJe+7TpF0lb8ds
0TjdxR89p1ep1Rh/FsqmdOab9R28jHZAjKALGn2CiQb66S5NumvhEJXil47RoK3Q
m8JCdmjKVF0u3tGh6Jkle+lWil9N+5fHlsQf+se+RhzmQ6OkXiwmZcVsS7spS8+R
26xEAw19Ve5w5P/EvuW23DDDpzQqx8sWaBzwAj1tHCo94xAp9KMLbtsPBjgpV4Lw
7FyhLqdTJYxbrRBsNZaSNKixzTLUAsioGuXBGwvUz301m2QrSDsyrjwBnjCDkPS8
GgPn2M3wnv1SmfDe3LG0eiBIal9Tb68OZwAWBcXqH8S73Gy3SC2/7v8vlGVhcWWx
HWXeu2kedsQIjhzzdSkq+U58nAsrv6CwH7daQoE3Wilore+tKijnpmerq181wexb
vpB6IF/AJiLtSsEVuxGlEomqW/HdJ4J5BIjCsV65hw9zQo1qmieqPZtJOF6vqj4f
CRkAMCZG205jWatiYSCu+H4ojbLQ0Jym0GHGKqbOohk475bdBLBdrmzoIj7vLZTh
uDB4hhuPh027fi2BrpZcg9EyfY03Es6Wh2qEbYLgkTabJnaJnmrgnNK2GkgO6NR2
Lb7PyTzAyxVMnSyFj45/1oOBlHDJMFsdnxIdP/bmCd7IFuqwkNnEgnIsTVUXlYf0
rHtRJNRJN9ugludocmmgwUtuqjGajFkoDKR3m677wq6c1Q4wTPtRQ4htjXH8Kx6y
MpqRairpS9R9rksMGDjxjl4bKbbD41rzzCx4hxGghH7fuEafsv0c7IlGHqDIQGbP
4NVXHuPk/FtjZsgcAWzRmlO9dLOwMe9IK4kl4zf/R7kjYmvloZIFGmahN+cToi/V
1VXGupVqRti2+g+S3Goioq8BEpXJiQfSLJmNCoh/W1GRdvhgHWsVu6+HZPvYiSCC
RhbD6TYSwsYtKpVKO+Cwvi7QW0gt43BVebKUkfuaQQUdNNYZX/wX0PMiU7Remb4n
O+Aqng1fzfMTrMiyMEEpuEv7QOYrUeztZRFSLYAgR47k9dHGdyGTlJ57tOysqUBF
jQjMpiUqLOtbHwD8ysDRa2n27iX2QjT3JahUyBlYceKwyzH28URfDJAaDbNgaME/
ZJixYfd28/hveCjeT2baUuH20kwDwTH0g7bWqZ0B3Vr4xjEKPiF+HLnXzPVlKuCA
TAaTZ/VywAOgj/V8aUzVDdjyMwWapiq1T1VIAz3HV3c8i9vYLjTi7byR0ewHSbRk
W3Rx70SqK1+lTAlHmOnfcFEDJ1Oj5HkIYa+8mMuwfi6vjQzkcDh8jef+MZdR2pti
VE5iFaAYZP/LDEOcKjH8dBuVmG9TCyLlvRRacobSY3140rlosaHoLU52OvJNFJfI
aDFQ2PXH8G75ckwd+L4obutdDh2DGW8F6guXFgmO4ZgdX2ejbuFD7Y64IU0Ux/tG
qWtbVXfMOjAL2Swh4hOVzplHxaDJz/+5GyoTbSTyFm4XQAtyvGgAZJtwRT0n41W5
BwfSq0mpw78BWUkPKqi7kTuVi2N9g2dlErYMW/1mHOcPWqi+LEYIkpzaVqyiX22B
CEE+xmw4DcpQhOZ663Xa4WLD2jO2KILwgc7JAnhqhK4jOsvwo/XTIYVBW68fmGXo
IxTO369Et7IyguY4K1IgwC+NYO/BZcg7yw7md8I2e+kC6blq4dpOCqJpTuQmG1Ad
DJYkaDS6zx12NMngWzPLI07x9tXL7LEQXvAqfZqzIqVk8FAAnz+5MDN9eQAHhIoS
QriJbQ/yYuWSteD2Vc6WZbtSvN+zHZbxbbaWjeJ+yadDUcX+TNgpn89vCWxpAN+5
DrB9PtVNxwVmhkswM7BA7mGUv9GgjtFTIvPBmKnk6vBxx+coAWD3z0ETmDpLLNP8
aFjdWXz1oj4hgkz5DIQwfcga/ol+9faRTTcHtRps8nDprK8cHd1/UcVjwfOe1Kss
XwqQ9ibIfOOJyCwaofpSv+ny7NTh0z+S7egi+9jk9dV4zKFo9AGLJGMoQu1GxKLH
mMEXNnfbjAgC3ytfDBy6M0Y9kKk57Qk8wR80n/rZe5sHVDnNToNEvhr2UiaYFcjh
tiMLxfmjMvBH2eE9urgWCr3Wq5mOraW8LoJMhWFLd4PciGEHW3m8n52izIWryPYw
TqQ3oX7SSQ+o47lPq8RWjhC4iYovgeS5MDOYu9pqR/9SD2AXqwjb5Bz0sWxdIVD+
N4pgp0Vanya06UhCGXCneE1uwVi/wzeh+j44B86qT+Pr9h9B5Qs+Xn2YcVRLRehH
83/3cz+cL1TXu9mIldVsTNaxIKzDQit66byohsk36fqEeCdeXXsao8X0RoJdtXmJ
Jev6T3I0q0HGmsP1CC9jT7enlS9P8bJvf989Nlz+FG+aHho1VD0fGgUw0qsAM36Z
+QlkByWMcotLSGB2oeAHtkmd4pF65uO0c+OwZMfYcVo85hDZTTHwrUC4DhJYDkbt
Ie/g8d16aOAPkND2C+UqBqVGgCOIZLzF2CKQ56j55fIAF/CJDvYjnHeCNtASn9Rx
Eq/0yc7ZbVOfIK8LNtNE2+jrFO/tmUKJzxU04AxyMKjk29ZS+g0wNWT5VB70irVQ
VPvf4HaPcNMkAUSR+KvVFVAUNtHtoerlKh32ePaIXP+yVgfhTIGLzNjluKjDD2HO
dihvPSo6+lGvNsY0YinNs1i7WGN/Xgkf90dJ+Cf7qicyfaoXUMBATAgRt13AmA5b
5ogkmUbblbgR5Vc+tURUPBvbpcfJ9NWKEoD9x3kDyq2pO9YBHzooqf3wmnylCIik
fQ8G4gvx//AZl6Nhs4LxZS88YB5IpgMvfYNA180Ru6mfJG61mkqwtMY3l+nobtnb
FApL7zvew/3RvBBlJNhAihjmFoGb/shm7xsRke/VpDiqo0l3BcqfK3CXCQEoen5V
wtSAdIGcyUgC+QYcliBMGGFBY2k8EoL/AMGq6cxkBMrnnDLmxvAwPjgckZfaHaSV
uLyVhKu3mHkug13wdCPltRsqokNuXapi3/wkys/0sHU0h2F21HjZd4hsTzjPrDfM
2o6ij0X7XP/QyjszQyTpVRvmLNvaQBVbDboshqzkP+iVKNpegDRMssuSgbuEap2e
KIz8WAZcreiTgtBhlNKr6HjqefrbW2hD1PVI3WpsQufU2JpvR8dt6mB9OsTcA83v
V2jHCGU2ivw0yXJ2OK9mbhBKAN6807AjDneZrBmHBkFLerlKxlj/1q9z77MAJ0Uy
pIYNgtGO0VniNb3qx03mIvoBwpapGN94/khVX7YxFem1JTU0uxczif5QWFQVsAox
Kro5FmXOCl7DuqgWtPXG1aaaxb8r6XVpdBA4Dr4cc7omheeuXjzOPk0IjmrILkxt
5gIWQBkbEyKo27ePh0bL3tgjBzbmkZ8y3N6Nmammo1KHgAw304Kx9FNsKaXg1fKR
/4DLocerKOX2Nxrmz3CUa3YTFj6wB3kPxfJCwwthGgY5oXyZgsWcdfWocntzyHZM
xOLOIeNz1U9TS+FJM2J/FJsIClylUhP80cGqGpn5Ji9aPZQsoHTswM37CrpRLtFs
Qpu65b9cxm8AWH+BGG9izdYpWXg7EVwA20HgbRe6/B5fDDOl77oxs8P8MvxB6Y5x
iUlniXef1DMy8c1/pKd8NlPciOvQHbDuIqcGWgsGCYAPgUNgI+l/dj54NgKcEleG
d43w3MiUBu1Q0WpvwP1kgHc40bHKBfo3uRYW+9HnIxSsRiFFTyzWU8LNuOwu3e2R
Nfo7nY0KEi3QWqhyO8kOeujQr5MkYXdDJW5kNo/ZdzTerV4Rx8f7cfiiw2exUsPm
baUgyoiZ0nA6QSC5f+5Pj/02AyU3OylDWzOQGxCHTrMmBiNNUUSPixrXa9DeUoJA
eUBGn80KzTctzvDdePWoxVm/lCFILDUoQ4puXSBteW1e86NWA/gJeiuCKV2XvSnT
FaeJGum1NXhk2+izZFot7jMYwT5bRr4fzLV+XacXEXelQIFZbpPRpi38D0Ha8yTB
C23vdoDkiKXCxis9QdYsRM2t533nSy8eLEbBhN91tZ+wgeWgza3H9ZS6YfZdIheX
2wvN5p6D1I4voU5Vku4ukiS9x4bFesBwPUBkc5q/fzljSAPpYrhQE5vBIFmXiGql
eMQxNdwecKNhnV1jl34AJDEeFFN8wEkVBTnOSkCMmXcKErzDOncSZ4V7yPGRxAMO
42wVeoCp9v2u7bGanXgJXC3pfbd4YjR4F+VTzJpTXw3g0K0eunu2jTp+sD4rCiVX
kB5d8z5shOmQyxCQjvu+WIwRD2voBmbQUzrdwwU75PDqLKoJHjJ0j7VMJq3KqwCZ
pFmqMK7F9jMcSy8DaarJXDVjWx1VbankdeK7V3T9qobvcbDffz4rhhqg78Bvuafn
sCfUyaMi99Kyr+Vha/y9a+INZKJ6nW2FxqLEzpC7o0y7v1ONCRtNOG7RnhZjwZeB
YK1gVhjkkhMlmE5qVgJ+s0JGlrMoo3tYNfbguccNKvH4nZMV8RLFYI5ULWjutX0w
rHvBLzLh3wmO8Rfm9U6PbXNQQ6GvEp6dKv6k5gnlbIfb1IjyA+lHyZKRWQciZiJb
Tso3SyQu3ZUb6osDvKq0JhloRR/6JXjkr/DF1uN1RJmVYuZZSZZOWa3m2uZUjcba
+r476guQQzmb/aNY1RHtqSZ8a22TzSOte6vNnGHsoMXUolQ0YoCQQbT8/q0jKTla
8oQAHID5wQCEBwJBi5TQCfFUphOSv2cuXqfmzn88NsQHikV8V/pgCUZGqD6ZCxjp
n4T3U/eEC/P/ieKQO0KnnAFUD3oavBoD8YieX+Ae+5+p1f5zlFojIY4i76oZcluK
kn0dKFcXzkN6RNVjNngaZFo/ErJ/6QHPT7/8TjmQLUSAVvWdWx/muMQavoF95Jlw
a+O+69dhfJHRt5VvXTZksYcIcn5paEqMxkeL8aNEm3iJT2zFxR8u9+oTy9Lw391d
NjcEkfqgt8eymSkkg5uSNSn1Kcy2uO3EUlUGg08xD3Pgf7ryQpZZxUYOlYcnCgop
3jAG6+lEfaGcyofLBEvAovP8HDw2t3LhAcZCTyI6WJCivXNU8czKslToRXHfmCCZ
MQ58jcsHgSvE1eK/bt/IPJcKsB+J8/vwV+iIhjIDg5uH2Aq0QEEpKfG7IpuC9nA3
gMooW6dffExa6gHxrGqYxcgQsR3mml1cWM2AVOq6cCO1UxjT90lwmVzifwDpP2ww
2+tVT4SulxLAfHSv59cGcLWDH4LeGaYjKUPq7TLVfIw/KHoYUXzAWDnX8a7dwuLa
QDsA0wmbRswFm8uQ6tLHdqp1YsrOydXeekcabrPNAVLr82zS6uHg/PlWvexYHJD8
DcFvgZwG50o+bZRVMLMp5hJu6sg63rOcKPZJTZOU8vQ4rMfPLffKIfR6mk5LrYoG
Dbgtt6bEwMzAQVuc6jBKLA==
`protect end_protected