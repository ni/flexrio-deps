`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8496 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRvSzIdqqwO5JLOHm2ufP7ErxMLNy/dY8s/nYNHSIBPNi
jBYFXhYUdNAO0R8/BBV2l3ATp4QF0HTZH1iwbZCSB2z1/VuiJ0k7MHGNN1OnDfLa
IP7R4cxTXoZMs3s2l/EVAwfrZineQL/+ny7cDtaWv4UAJbtBvwXAuSUePaYQqYp3
vL1GGbHe+Bmzo9r0R1F1aa+KtwvvvtX7ovg6AE/aIaJ1eA+gMRvGAGwoehjeAtMZ
Ppfc1U9WUZBIsgbt7aXKa7uZjzc498DKDBOpW3Ysnx9X0aRMWr/fa34Pp6Hhlegy
fZmR5ruPg/sKTBxh/RsaIJ7ePXHdf7/qsD7auhDlMBF87fAUZWRdu1GoMzVTayEa
l/aCdHmgqzeTuSBZdtipbykR4n5y167XdyT7nGGRTRBDfsdPCo0yjCM8Ru3TNo6C
jOi84+DwfoQBQztWjYA5a16PIzYrnOGMK5iiiJ1IDjXgBE3Rj7jNNRCN1dt+LmQV
kVRqsMc6snV5nrpkBk7qbp7l/cz4A7/NKadAuyMg1T4VVnkfVX1He5Abb0fp/iEE
A+N4qWrCeUeXpxNzqd9pSXpLAMwFnSTMMBQrKi6/1bCJCai1kR4/m3vbDanN/jcW
uUhy9tGdO0PvRD5rgQM16pwzEgKK30z3BqbpJGzpW9YN707dogw7uvPF/v7ee7+l
etvGlwJnjRs3oxx/hVtMTI5jQkxzd6Dp/y1dv9zKw56h5Qd3yqab4bObbPh6MwrD
ylttvu9Tvckg/bH4QN2QaENcmTfBFFBl9/pjKRrRkcx04qh7Qv50DCXjOA2ZZDYp
LPPwqgR1i0GZnpflKayPuGIiC2E8MXRxnCUGp9ouMWbuBHWOwkU/5jch1N+yuxi3
AiCN/XZV7bS8EB2fpyVjtQEDuw+y9vmKUow8VMTyv4jvsj2/J0slyC8LG0mIcePJ
50V2ag+DUo+CUhCWuyQy93GN/xrWV4y3fI5EFrX7cc0apTdmILtKf5rSHzek+ur3
gHqHDgX8Q1vXZz9dkJVoY7gnkZpZXImaHX05Nj+wWGOJKoikl17tEUlCkFy757eE
+Y5s5YOwidMDWlH3l+NgJcLF7735McowF9hKLMZ395hvtRsqStSPTU+1BbA76K0a
QdLyUJ154V5Z4cpy6H3juwXpU7bmBxZesf9f+yQ//7c/SB2AXbhfZWBcIhPuf+XL
w4qhwUYr6JMqi/NFKFnHWhq0lZUds6Ov+fmz2oWjO6eYz+gzMBHB9ImYb58qmKGt
E5e8BGi+4Sg+l1f6vVRFx5FFYH/Dfm9gNgzqs4G2rXqgyQ+0Wn/GzL5xMVtbl5eZ
bBy07Dj61ipy2iWvOg+ATdkptH/FHIwHCcc9AgSfAQv+BEKhve/qnhOxXVHaaF0g
oZbJhRWZUeVXji9NhalcPopMlxMjVAKwjw0BfzSoKGy17mK+uZXJPtQ4dCvyG4X1
iFVcDIwYKbn9L0jUSvJloxiLnYrJbm2RAsnNSOUkjdgiSrCAtMLLfZaLm8KDQ/LG
q3/D/kiO5M+1UgZqQ2mfqkS9Pk6satdQZRNCd7BueXmtU96TSdsRNJ5XTJYX2qpv
fo6ddCNIb2Y+7TNbKMSOS3L213+vSNgPFK/JrtDWAXEGiU84bt2z5LaQ3OitR47t
j0iH/Pgt7wp775HzzZsKIe7tEBsHAXhsBnwGhyV51TC5mH799lTYoAuq15WkQ3cE
8CxQn6Rw59TzAdOCt1su+yJhmMXnIH10+yEpp0I4DQgCj/kssf3cVkJ4CzhZtDDG
lzzGKcofPb1cqOcyxBj5gDIGhJoxPdfr+FJTsDanaVXhwBKBwxZZgYReY75hjCNR
ShxrnqwtM0OZCUJcnIcnDCkX9kXzoI9hhRRiHrzU95Pmdkuq0KvcJnuwy1Z43D1z
N2NHwdwOQ5KW302OhT+VXfLEY5PCpjOpDEXbojOB+Hd1lyOnm/qLl24NyIaHcXM5
7xrmpfsvQ8K4RBz3SR0aov7BnphACCzm4CKLUlFNMDwtUeuWNyrZjKQ+yyim/yus
Xx67WqquGB3Is8ZPWs5EdhWNUUubZUzMkS5I6yCPYRcWCoeM5fURyItiP0uu3I9Y
RBm/3at5GmVtLFPKXBZbImOU9xlOjtVeS1n5fO/sNhHrUy8hu13ifA2zrK+GRx9k
ajSt3INL86clZ1BxJY0/DWKIJq0pLNPBAuhrmQbJgKYVYhXLFm1kjh5UhZDGJ/zF
gFThyJrSUNi9+lgWVoh7sIXBs3X4tSOG3k/UL4WPSRqoyo4DWRmb1qo/2nbCTfC6
Ezq24kCgTpYqqjygA9eYpot1furcKfDCFdkTP7wcBd0DEv3VE6oNkoebS8EqtPz/
ksxPre+hFFPfkBxyFSPNAyO+wr3lkdx9c2AffTybdTPeqiiSCT8Ff57r5ctCwNgR
Wh2nArpUc7moxrQcMalkDiADcGfbsivNcOuihwA98YMYi7Yo4aQqN3D/7RYYVWbK
Qe0szd/VvPvigHinGy+bYAxDbC+C4q5ie7IRVgO2YqENTg23N2GJZkYqEqMmR3oR
PKUmBioohP76sQUEvxENyJZSwIHxECp6NVakyalSfTz0/tNflO7ynVwjTd/uUaLa
242Qn+N9KT9C1E1OZ4gFNlcM1VQbZeI59MIq/jcyEzV/pbkv73EgIHHRTCxTGJ/B
mEbxxFxGenKQe0k7dqS/8NYS/ZVtjSCzU1D/Cz28HnCbcHqgDvsVXpjqrEnh+ixR
85Cvgv294rpjjUxX/rsGeTw6HIJuQe0FhHrZk+8WC2/4AhACUBi5xychSpL5CDfa
vHS6VX6ahFEtR8aBhUGp9joMNpKfMyniAHxT31h6wZaCv8s6ppkJTaVkTOpS2aaC
37zUWmir54TP94+uKW+8yP8vk4OKOW71Udnu1zda6ZWleV3L47FX/J7ZeF76YzN8
JleJmwdjbz1m0ht7jrhxf0UhTQiUv0+4+TaCM76tPT5eaU+MYGihtXSCzUWYb8dr
ZBm2lvDiV1q9DrmNp6CmKWw4QWVSTVfp4hApEx9CZwncKAI4g6eLFxfXiwyVgnak
t8aWzWeWAXQL2lV2x/u7zJfKCEHxwgAINOCZcSFlH2cPg+Gzr2gYr2RWHLZQn0v7
85s32JDoh52x1AGYqiI/ghCY4cyAMlvJ8sfACiLVnOmMcULYWzlasAA/Y2ezzYYM
zqfLRtcno2tlDdFS7azuNk4cSmgzmunPfr18B3eHK0Jtdg1Z2W+HMiCHPwj2U8Zj
rDq4fKRJCfRymbnNG1Ydz2xOGxw44NJMn0fzKXXFkxmmP/43INLEgMlvVfRGszwk
SxNwLXE0BJjjWAlLmBhZQrNoq/+CbMLWkUrMU4rkAnRoSpdXZhccrHHBneDaffQ1
ucZw2skQSv6TpSXDQljf/YOb2H56YU4IUjHyBy1pQaKg1g38OsusNP3BHUoAI20n
68seK/cJ85RscHo2Mt0Hipaz8Wf+K892zlaS6C+UnLtXsRur7zG0m0QoSFuxl3FE
Q4QaxBaifYDfwpGuoCY+BEIhd00GZyhl5iXg7sxcyN2nCe6LmHZwt5b6P4sWfAIh
68lTw8H8irnIWMbtWKMatDTd8K2L8m1Z7PT7CtqmEeCv5wqdt2cUAwol8Od7GB7S
DvczOCujhixd5F33+85zLq/q49q2fgnNHzbCL+hm9/6iKVixwRJsmmYPnWbI8uwn
HxWvugV5P0ra1FwjTywS+Kg+WiKD93R7lT4x4SkjRfcLH4FYiTt+57iiY5D90wqg
RIyq0qxqKcW31c0oPn2uqHxFtgKqMyjtm3siU7hVlggF26GprRhM6+l0J+YheKsm
MRLD6T+FW9zAs3ptKG15QLN68dJ7BvRnDyBkXItxEpzo94MplpxafsNbfpSZE5mF
M6L6bMrpBDyAj3GCMppptiIxI5759ojjfLEBKjOH2ywagukwgJKz/pOKRHFVYmLo
++FpwEFJzzSDZVsIxF6e+kNETDuMmuTdkcg84OmdiYds6t2pckyGNfViIFEhWkVu
4TliY7XePEYM8sY0UMJW+oMSbgrwPwgzWkeVICkcpTbV7hhzChs2eiTlGSVn5rv3
sZTpKufXSVQ4BSc43bMep+erSbH8Zlzq1A6Jgxvx0Lz3ytG1HZjmwq45lK8SAxjr
Y5HT4xAX5rCawtD/a8GHMfpdjZCgMADA6C9C4OpCPH+x6weNEURg6hFR7KEGJsgR
/W0Gdi00AiTbUIc2CmLBKRWT7SNPc8/Db6HchUcxqw2nUGMfaCPQIsq89AhC8n5c
UBAD1V2snGjMy64m4cSjim+VTNYOjgGHWK4SUaM35oQVF2uQ0UPeG02iPsKO5B2L
xWKxNgRavF+7+yAG55kUFZ+gh0Qhzh8OmUqyUPgBIDlDwhI+1yj/Ck8K3J2wToKu
MJ0rYWCfQos3318Gnz0jv1HKvVhFvSJ0OyVo5EcvqzqZAb5M27s8lwNknsJTKoHM
sv1cOyzLFvt17wTIPIp8T1Sy6YmAExgHaLvRl+9VpU7B8gkh7hccawndBn5VASYi
nbiJcdyEZbApbUABCVgYr/tpovdLNStK3oASXTsSTfnUjwHVmKqJhbsF5K9DrR3o
VXVwpzONwPrDubfb2hKWgcDxbEcQbAsTYlc5nk40JzWjZBAQmLFfNGdEdD0Kbu3/
/ZjiNGxgApb7C2/DDAvzheyExvssEWfEiv1KsbHVu2iAbP6wrlLTUX4jHjcLVx1d
FcDWLy507z9dR1tDYWKt37E+5hwXr42hAY/Rr9cJWvdi4DnnwdNFd0sY30h7k8LQ
iS3WI4a6h8e+d6ZXEY5FcChdS0kNUuD2wLzMEvTt/U/ov5OBmGx2OmGpp+uVNBoX
CA1gfMEZoXUSjHYAwEL4o0dB2D0Le4etRP2TJnhLc/ZQxroJ7M/wXnR6IAAakSgI
Ts3QRk/V68bWJA7G+9tny3No3zmo2UisDNtK1ZLLQcsoivoaY34qBeWHi6DLIkD7
9DG3/9T8U7EjBKMWKIdFWCCaCPw7ScGHNROf5rj9O5xVW5dKI8jyZWUUIDDcyAWW
C8o1KWx5YhgXrKFUeYxTvkrTDlknB0Xkg1Z+diZ0CZylkleVSxAWvXrgMJ603h+O
51HEX1FNj6BITFT94IEiQcv6CJFVXrO1kxI5liVyu1eRqec63IR6QfhE7Valk39C
+aBosY3HrDILv5yS89arMI+EIY0J0fgDUpBQZP7KmQ2NtblvYPl7lxjz66HseiFq
Am64wo75yOUIJjum8ZLJc0twv5hQ8ugu+Mvz+KKehPTStUqpKJ3D/571KkifOcO1
XINfkEvS9bWVEiMKoifQfCiTzVfcEp1zIWLEWBg82y1QZIR+JcEBnSl7sn/7lmRL
mMc+9yEHzYxUom7Xw5ofc2nm8cemN2m5S8xkWywgHX5e3qW8LOynQaoqwBGT1Go5
P22HScgSHSdBkWnF29vRl1GiYEeJVbvi3LJXPgT4IsyjAqXPgpbhRHl6q8EnGSjQ
rWh3R2S81RGrkpaPZdQW66bOe1M8w7vbUmmyRt8zDJ2wovHX3OR4FS3ywE/K4iPw
DN0ArMXaxfB4TrOfKbjWL+azfBNSa/0XehG6T+was63FidQz2eYHJMP3nTKCua0S
g6DdYmssgaLPLq2LyXGJ0lxW5mtNsADr79lMgS0ZscUxlF26XhzT+Hh9jDCAGQQS
u8joUJvIcFd8nmDTpNWIozqG/G/TtRK22kxcU/CKltpIhg4VcgZBPKPtErtMihxu
yvRMAl+BiHNHkDtBhwtSI1+PE3GWOfI5rvPYnL7wCKoTCgJD/9sQ1tylCrbOl79O
a1FYucHonb9JjXjnYdvvK90FW+ssJr43T+WCjKpsAklLep1MorxZJA+UaAli+5/A
x5fCSGQ/y0+Oc+WKQW+/n+iRTuHAqVtBD9YviPCZFcW74TnIiRgJp6FbnJNbx94Z
UCfQoXM3aIYBxQTuMPWu/3hOZWnvK4XRqCFiHoqOvhWoIxqXEeU6H8PFl6D9SPTu
dioJ1qDN9yHoyA+pVg46Mp5ZvlbgpYADpK0nR6ERDRRY/G1OKG/TZitmiPCyL4cK
BRbVQGjobfMveX1blCQf68HJI60s9sM+ZCUzo9oGKIyXhfd2tvuUp6H+vfGW6LXP
P4qAUx6efjXW0XrBieOp+elRlMjdshhDOUFIJVTI1pLbkaxN+vMcrL2Dk6YubMGQ
+l2GmozO99WIG2C3GOlJdhhnF27qtZYbDVb/DUFeAQk+74txsuKXnILPdN0XM6U2
6snJeYC0WMF8cihIA4nu96IpFaUoIH8w4x6zbGRq6hYLpky6xTcRMPRF5N32BsTz
SWTDno5qaUoGbntrU3pz+YEuYDNMXkmICaInJ//E4NhI6wFEoFduG8omcNIdLZhn
uJDd3zBgYno8lemyV5Zhwv6rGO+Nc9PWu9KBXsTnGUL7BA4/6BXx3Ulqht1oXjDs
HegAkz8Xo7NWN7D6p6B8boGTuZi/fk4PK83dX/9/9f5rzO1SNR6f7L/y57CXlaeS
9jWwEIFmL4TDvxsjYZ/WVivFpPowxjR8ccD2GLWheiqFLsPb28XNpbY7X0cjp8Or
fex2OsFbKSuq3DbX8C0vxpab2EFzprasBLpDZKF3RKPSxhXo+IrUQ6rjo4cqM776
Sdobqp3ppRHsBTBbH5FkbfL3yiNg9te9dhbL2SUiIGgvyHd3Voks9MYgLxVGjRQ/
HWDBFBOFCBhGKmUlH1aIVYr53jAqs1YlSSP7mNKNFKKkhtSBVsJXUkOzhydepq96
Aims6j9N8T8G17wi1O+KCjBgeJ9qLk835RUmDVUG4YXn2/rAoDp4JPTRe2crsuK2
3K5HwMX8spIKMysKcMPKQHWpc95PpE5nKHrymSnoDq3k4B5adZHJFZvT0LcALCq+
zh5BtiCfOwhCdV3SfRlE8YWM6di4E2f9TgAb9b0OUw6hW8xxrZJYaGez3tkkArWt
jAmY7RRPVByQloM86glB2Ut2DM18z44J81NG080oA9AICbTYGQp0CZkOaMHGBF3e
lFVFIw/YFykV1rOYOLl3A4TKZg4BxistUL1+TQBer3JSt7MKEDXr9jufmufGVwb7
+qduobIP9dHCp0qagLgUHpKzrbzhY5C9otEWcNA8xpbvb6GSU88od3k8yEzubyG2
/5MLYTkitgBso05r6eJ6QrWVXaSZQVjTPIJIQZvjuF/0muKdGjaTiQs8STDL1DDx
crrKP9NfTH4ZNbd8GK2oAydWjuKekN1KFZS5uljSwTdPYH6C0FhFbpe0oIpd0ETv
3+4PmswRc3RUgAfymKEFFDe+F6ORukZt7C9q5bbNrBjc5xxfjAwjaFmJrsH/fQ9f
LgVXsiCRQF9Mfqp+y79+pDLIKX3MjCNCrF5NfiW8fYS9AnEYsjYoU8ugdZT5ygVH
wXZkaneaWd+xFqsV3O6HV2Qjpcb7q062QAjGsOt+TibdhAMdTjYHTpfb7LvSkcCC
fse61es5EFT94nZfKK1l9reKSvfxQ/x1F8EpK0fTqvsGoqxyf64U3wjdnPR9aiQz
z6QUyWj66ABLrkBGB/9D28ZeUNxElaayM04H8XeWR6fHNp5p0jCCcqHcSnx+Ur+o
xDUdp3WdwmilPIfOWMuJlmsesP5wQgwjvYbqH0CzcupWg0C0QUe3k9bxWzQWNzWO
2PbZ09QOz+hL7Ts6Sr+urqCmXDfDjf2EUlL19h1f92B1+pPvd7DANOSJMUXjhKsB
PNvK3b6Cn78EfMECRmYP5Fsqlf0tAqoFGJu9O0lqcZfjbR3+XmPeZ6/aUaEr9jwW
cklLTPicRrbTnpnQZJTWlBmmxZcACdGbVnenVmicPCJ8LvturU+0uJNYIy5vtisb
OLnLH6yF+ZzFIX/gs1BxqrYEJFz5THElIY70yxaIEWgY4XFMlRd9hoorJD+HzSo7
CiZWmmhjlJFWUNMuoA4DDKPMQGKJw1GcX/3ZVGQCdRXiOj/5t4tERcXtTu5V7v4R
uwOJmmYbXKbYOv9YZ47AYnskmWbq9jhuBmEhJbT4Ouqv4KZjATqgJyIa3RtzwT2H
EsyMxYmdKuXMay+XyCOc6Sse+FZTokVy4efUqfAgHYLwdTNVs28s/IVTWAF+vBRQ
IyDc6LBNFDJU0jyhSsNw0n6+DUBpOmcwyGD2eKUdTOCBqs3du2mpo3BF3L2XU7Vo
/cOuaENwx5noNyyGSr4Jtq5PnNJ0z1/qBSHD4eLdA+DjGiZkFZxw0SIQsUNEwzv0
67RmYkmBETJzOpl4YeOkMgpNVxqVPqSv+QwM6GXY48fvh6QzcyqlxXKIPGQGwhcw
3qyIBRSSpOoqJp4+Z9wxT3S+Pl4hfSDgxSJo0CI9LU2li2eyP4syl5bFXCQxpSxJ
NiOKO90+Uiv2BZ5+L50SBM/eHPPpTMFqvSTx6P1v06jtwJPwb+bpoloHFasdS0h9
68zI96xgwKAFtQoOyZIeCwyx3MeVEt+Lxw0ubt3o7hjQP3Ed0tx+BTqGsIqaIwVy
Bho1IiDtgUZwA50swZChcnEPJSmcZn5fLOAo1iX7B5CtQDmEuNXbxqV5bNMRG/PM
8FDRH1+Gh0RCVe9nRtTIcEzxPFjiiNagumPotyXnbRqPeXtV1CmFUpguyajn12hH
YgrotxFpoSjVDCgUSJJLwQJRRE1VJq37wyRyABzyOflp8u1manEgT90l8ZKeq1ED
kcoxkLSo2VHHUdyFDIGyJa/dB5BP2PWooNcL/4HtlJ16J5Br8g9N0DjbvAdhgvgS
9LLCa07gzY+vQQ0IrTkCGcr1/8LUE1T4qcnoz0u6kTby4DWxGT+Wqzzjh7IY2IHB
Wh15QvIs/XDtQnzZHVrxDkUrmBFRnDCvw495hUgo+pnvuX5vKhyrdVqk+Jhyafmz
ky3UNa4315gVJs1RaByin5g9jcSeL9jCixwOKGB32GMLC7Cb+RtGeeWv9b7tnM4V
1tU7e3OqCeydIlpfq+hFy6Eq2+foRPQr0EJaYLKruSQIL2vkiloGtz9c2Bq6YQoD
X5CYEE+3F7CI/dJFbwEvr+DBg832ujKzR6lJtvk6ldjOavYj+BhFlrXt+VToXEBg
pf9fkNg8vQxE2e1LEE/psGvP86ZnGOQwJJekeKU7rtH8cFZmHjusnAYhY/5BGHyB
uX4V3jJFkCSsR37e/4CWKpOLbuOZTwRO8Pj4ATIS5TKTdOfELRl4wLjvMEdg+DwW
XbpG37pq2AP9Le0jNtQP9yyjwFwarKyv6e/4lb/6odfqMDZqQXJ7deh2UCZVEBDX
Q3DHzNav0HQZ3yg03P1MZ8tcX4Ji1/jhK0JFVqBc05SyQTWH+19lHxvW59vbAXro
7WcUohX+jOfOaz64ijWCmAyVPaN0IdBKXK/a0EuC+iKMHhHUzcrJ5EWpVr1UEvCv
34uv6pgPw6mD/MmucQ/xfvoetqhZOhTIIAPl4P/nOXfn7qPIB+A5bc8TR25LTd7s
1grfVEwa5coPQjownX1qcvPb1czjK8fsVByhff7YYF6CzNgH5CfleETtNyftB8aK
aQa8k/7idN1KLOkIz9TzB9oe7KfU1KhR0IuoyXpK9sdbbe8huPk2OCzayGKD9BOf
wszzYfPmIhkYZPwwfRHp4tKYpOv1W0z57+6g+OiHULiTFUS9v1PtVd6AtpssJ+Dj
0ruSerVMnhkRJ8V9QjC3PphMZw2hGaIL+nd8+1yWaoT11Tn6Mh3e5hzQTvWPy1f/
17Ujd8AYtRHOt+FJQQLU6OFQAzG5mZQHI/K+lMr42SFJZOuD4snKaUnytG9DfWvw
jeKoCM2DTl8fDlcZg9MMZyKvsAIsoxTY9B4EjWouT4PEo2Irv/fZ6MUo0JAn5HHO
7l/ilBrLvdVTaqMJO/Epm+PoP2WlKK7oams6o9F6kgX7Cy6yDFHmiKSrgxW9uHyG
yGj56a93e82D/b191W0+0l6RGxYqmKqy673ZCFVZDa9GJ8DeKU7wTiP4SQGMNEr/
MYfD2cp7tlzGbboTupzXhXvKtT4MVPhRhv24CPC8vSCITYIpRSZTRI39kY7h1vH2
ir5UpzMaOYR97Q1WjQDrwmeRZQHff2AIePVQNRfecyn4xPzExNXC7MdYK6mLoN34
9fT3LrCt9eFBuqhdWTa1Q/JE7NLI59plIQIBy4tCznKJ58YU1rpbJmroq80YqAy/
D4MeZWcXym6c6rqHBaP8bJv6TQ6f10JiMuNk84AoipM+Hom4IKm8SVkIxFc2oESU
DX3ewOSn/eQZNa/oFI9hGtHYvrnlu4Jeb08+Iu3Uce34Xjy6787KPheA4H5Lf1sq
TgYowVl4GSVaAUdrudv/z70HHPJ/aq2q9xur0Cwl9wD3Ve/qavfozfxT3JfBcGNO
sBMxqk2TQZ7P2md5sLNSbNpIUNoa7Rtiuij3/KfC59N9VNe3Miqy0Lfe7BcT0uiy
wfIVaB1dT+tfiRI3/N6pyO8m4JCfVaLhe7cYE3Dc1pLRcROnQCOv7cEh17C8DYp8
kR/ZAG7dzan8PRkzAsTckpH3vL2f5fTeL8nTSNbJ7/l1mpUMxEdZC+tiU+4N5hJ3
0sXTMfWyb9srzuk5dpquY7jka/U+VGNZHkn8N7BnfyHVXYqOlhczDnFGWgaFXD85
PcPZIX66kwbW1wa/zKNis+MK/xFC4K6qSE+MUnnqFtnnGwuBAdBH6nIl3jmwqUIX
NvwyPgL4LLZMUVvHTKhW9cA7gMZDGzTI+tUBM3uZlQvibRYj3zideUu4TmZpqYct
lPpVWRRSpvk9AuKzna2LuqHpv7p2xLFVPup5JM30jbYdB/AaoRpr664TjB/uCZul
+AfCycF4AaCsEfh2h/oXH2dcE3MUnoW81Q21N7fEls2kNtGX/qIeJOrdJVxMa5mY
bqrzmhCSJNsNMEVGKYSvclz+6Y0aLC7yjR0NZLg3nYuLxa8sGOGkdJ0BA6NbYXT/
cdkUz/B5jUCM4KHJsmlCeWtpPQdRz74oGjEz1C9tJYlVYmKsBBhXkmP1JhxY37d8
gld6gAuHgPQVbADZuFfRWHqsawKXS27VCIM0KgOSKUvjxh9aYzGo0TTHikEubuIZ
4B+zOTTNHWSb+ry/rM2MuL1J9znBN/9SJWdWzTmb3vNPnYmXFXAjN1BVxIF/9NvD
INwoWDdYLGKEhhJGBVc+DcUzwROqxcxZQJQPK4vQfdl5Dt3hGvSDZFSf9S5eqI1d
`protect end_protected