`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2864 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhAUN1Tg6/Lt8rBz7kpeJnZvkqEJUgFMmnPYYnXTaEG19
O+PqujiTadj2z9Vhaz6tMTRD3EZ+d5fYIGtrffEIgXWYOM4oU84pvht4+jnGvMWJ
jtEZofP8VlZhhcRLUZx4FmqcB+V6FV/ShrThkuT6bVQh5QGrpxinweNbSnXryC+H
IQPONPzzcyAd+aX7eYmiY7/2nnDlIvW/heHV3dPvCC22UCL5YPh99mSOwW0WTX+1
JJ6BAFQH3dK9HZXqaUhJgna2qdFG354j65pLhNjICq5uTcO6IvQmOcxW/Mm8Badd
ZrzMNlP+9rpv74AEakupE0Pz69wTzUQ5Q7FybxnQNQzPn3GT266LAkn7xV7MGGCK
FkiZD1M7qskR23YQ5c5oSe1XlsklHnQU4xYvxBWGY6p8Hf7KNrrElvUH1stVKJ4V
nJRh7zUIxgD+HI7ave7Ofpt/jkBm4zHJpmyfBqP/7br8BQSbG/7si/OBG266UbF2
kuOTFX9X4JOV/O8xDfIRzddhwD9zOR9JOHsaP44GP9tr9+f2Ore4ep7ysXO1/UrB
I94IHaJXBL14e1P7vzvl4dmfWA8KrOwF312r8V9k+nub9yWvFmzNwRa83ubPKSL7
+ipNdLQ7Y9J1C/LM8DYiIbtg2MPPbx5I83YhqqgK7yX4Mr1uZOSIdVtyKrZtP8uR
CTBPztPPjRw2l6bpMnB4tKSgC0MwHa2pMONb2H3+42VleXZm8eFpbZp5+hzGUCOS
rhEBS0JwaVMo2GqhuWDebsOmI+HZMDgTLHmu7OAkSXYU/6GWHnDembqhf+leqWWC
RC3BLIaGyc8pY3doWuQSMis/4Ih2eulZFNI6frpsbjizyenL5HsDUAR0Rk8pb9rm
2us7mpd+fzKx5JVOH1HkVae77D0FP4YKGBM4h47jSPyK/sjL1BVrQec2q4tFi45/
G+ffb0ofywMZ5F7jwH03M2hmcCVfdgFNAoVfypgDeC1ogVaTgymTOknO+4U3Ddr3
ISK0gihbgOQJUyeXNjGe1N7I2DsDHIiE7ZBs9i4hgH4+XR5c2Iv6vCmH9CzZDYjb
sA2Yy8T7CKEqx+5NRGjDBvRREOfZlCKBKU7zrSVkgfG/7MeC1vtHkfLxKORmwdNz
4zCLC79nDtUWATbw+o8lHxXecdJDFoE4kIPCd61Llv+sUeTJdH9fgF0Y9nwch1EJ
7L0dYk1oSucx9mV2jFBgLLL2j06dA5QzgfTugN6geTFrUOF3P7dDWj8x4MHHKsOQ
I48psuib+rxV2ZnoS1rMXQUn/RRkNoQYlWlmctYv78L0Q4+JDtxqPK38UN+TOohO
BkI3zhN41VFuP/yrvpmwRqIYkpKuJrLq1wF+NkJMFmep9zZaEQTdQFp1YU1XtwMk
8vED7vDdmgUeTqw+WIFZ/AOk+tDLkN1ptSnhTo2x6fP/x3J3xB8E6YP6dG+E2Otz
KIaegfB4wYGt7XLrNe8ceQASoD8C8qwZbFrigZhq5WC4x6yCiW/fMQprYrW5O55c
ikZ5Q9sUhRUM8WnD53+gLkhlIt8WXC/KivonE61Fq7mEpSlFsTLBPBfqCjDkt24S
FGHPDlV/yq9XDdRrrETKHRVm/vYUukWALJFi0IMzaXzodjDJzq1ZmAOH5smuWTRf
OsYpYtgh3Jkl1nQpumHVtA2ysOzalls14lnFP6Or0L7edMjY6JrEox8xl4XP6Z4k
WcYyTK28yHa32pnHIpULRRUKC7ayCKD1EcfxhRLEIcKQN92J7tVQNbQTaABk5zfd
XSuuzTzf1SJxjnAcsZ4ksQRkrsxLD4XDOIVYgLfudeyWk3nMLvzYZO4g0CilCqvJ
mWfgdZxeEljMMM9uDqmULvmIf9mrIH8mdvSI3Zj4nwwxE0tbTcs0nA83s92s/pXm
Gd8ggm747Z+DM2aDufqD5V27KoGJqBFMF8hLnsQhqW430hM++a9+SANEDMnm3+VV
zyyYmGk+y0vUAHnHcUXsLXw/RwAqLrnnS7S1+H2WFTIP3ZgcYBsf7rq+io4x6HrL
adpctqVoYfxmYFVnqPFmYRxlc2BxzTHeKrNFuf7t1XStZ1EUEOPGCxtyHn1KymEx
61FZH9hCXZIfV9K0xPLF1XUi1ZPWuNs3ZLo8AW/cjX08tajqS+3F4jAcWoJwgTth
GcyPvBd57YMYwYTVV6PB1w4R8LfrxMcYtyPxyme9zO3X5OnUXMyxCcgQijqWFmY0
N/cTyD3T42/eD97dZmELnS3+ckrsJ3yjjY+q5deqEINPJGfn4e0hdlCrrut6kiD9
9j1bpLpqPmwz77r4kWi2TzzDsphhFSVihz1R0p7xQKx8+BlbY9qlAD0mHZUxm20C
GMt0fD56E/V9/cNRHO08VRTNwnfCYbuD82Jj03ciRKFm86mCvOfbtUl7gyICBOxC
neOqthrRQp9eGg2dRHfFCqEsNToWpaJeWqdy81H4jdCugRBdNNxdiv3JfHAHeliN
BAzcU7t9SSVXbnfelu3EJwC7sLy8KEaAyrviIHz1N6M+25FoSCD86n5u0HIPbeWt
2UiygTpuJpCki6car0dz9jYREkuImv8tp4Q6Pr6/WTkbZe/rzWIa6MBhLouQWugm
cVLNhKMUCbpA1jbBAS0JXXXpQszRY+WZknUvbrHOFuECxJoRCnHffKkITceH6yrS
+rw8nbCoydncjwT13fVs3SlzC7KXVs816tLh7KFy4FkxP4qbeO5fGrguYrZ5zeb2
i4W3YAu2scIX9H6z6++GvvTPE6tSu15rviz8NkT+I7GdMPVdtE6p9KmJFob9ZbLl
Gc1Fr2zEzngMHAxndKJcnjPT3pMafgU+Z8+hWu4hkeg7vqsrOvQxjqbo2DeyV4cq
qlLZ8vKP+MwGu2g0oOSuUKtLN8iUiY5nqft4e27I7A2EgTKzhcUflFaDTs+fB4+S
9TTmTDNdtlGYi8gNj+FnXDrwTpsnnrZN/m3ks6VOW/wDBiGls5xKhWa5oAtf4Wo6
GwHSQz4vLGLiMEO6zZ0S2bhyBEiul9B5Kh03RKrFDTIAvkw8Z2S5NBx+lPKU8u2J
NYUhL3VNF9lgYc8rAFtIIIKnI8olrcWcpBUgGEkewTgBHs9RvhRoBKVA1wmkjcKd
eB4PxOgGfxoxs73xAIi8llRs2ngX8UgrHPh/9KHZazp5xw8mP0rWO8tbmbhI6yYC
35Ka6pAS9j1kH8XWgipsKWgQXx6qqXt69f5MMj9TLS28oEWwcG2rQLTirFUQJI6D
xUuQyD88K0tc6dMcfh82UHDubYTPIk8t8t6jGMQgGJ4CPHZDmVwqg+TtriFhYL1w
OTay/G1Bdz0obDMTMCedr/96GpZH7eomiX9vIWmvOBewPPVUvoeB5jh13uq8cvpC
PXux2kub1KggW+RcQAHepgHzFYSYoFQzy2mkR/KWQL9waIcY5hZ5rwEPHsrzQ4Ri
H2/KM5+WAAGnn7yuRwimbCkrpTs5q+fN4yPpnLf0o3Ej2IxGmFw24PoUxzxq4UIh
NkVVmp0PnjF4W6YFU74nW/Vh6FcaXwgsKwx+AAr/0UL9JwfSd567jIfA7/0pEaL8
W1EGttnfEGWwuOcXFUfqogtH2bRA028MDFePM/oqhg9DeFsnrQCpckSPOsysoKza
ZZwam5NIFmRgkIiTULPovfKNZ1IlBFkmF14kPdtnkCM=
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2864 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/T97rZhQva68T7JOm4bkq25
b4BW57ADAHEm2yg/Vzsfl4adqDo61pA6GIOSqgntE/F3zNsb50Cl7UL6VywDEhuH
DzFbOtp3CAjjq4eYHEDr7PWDlrEKjQwcK1Q+HpsEAaHj0frwQ6R07pOZHMT6PqqX
JLT+TyErLJqqbN9TtNyCoI9bbxY1/rngF87dqMRmEdQB0u3Gt1iKJ/oFHeivohh1
gat1R4ydqE2bBpgdp9MBm/LwNiPXQrZHSppF3Ofry3mxfuv8lhEl5ycVm2GjT1TY
LyV46f61V4nn5TXePA93n2MvedlTfh0ih27Q0q8Vp8XNyhtB7ynbt8HDat+atay2
O6GnkdtzV+7fbsNL9gY6NPA3sfw9eeIOGzGK9lA+nJn0WfMDnEVDlyrM2Ws3ipVP
nSFsLKrDq5gtAsrk4sNb6MGxewgP7cqNLmCQnwLX800J/GaARsSXfhIFj5VxO1RP
5PWY7v4wHj6Kvc3yGZK161ibA/A/JmWzniRcweWcQK44IkXq/IU3PKnqGqqIzJrm
FJ919m3lEhzWkmSOAxapiN131MxCWIKLOjI6X++ILfxMl2aNZ4sZS9aSEJMGmd7j
R4Yu0vboU/5tJXLDvDcsrHr5Vuy3EBolSeEcSPZZylJbACNgq0nLyXVv4fz3X5mm
C3UznZgH4773pkB5npta4DClml7mLsSCJaXy/XC0huHo5ooMgmbIMlSnxzzd0nYT
UVhSte40FeCCk+hGGfHxydEG1cfRpl3F/k+WQbdGYXhpD7E8H5Nk0rNkvRMAQgdz
8bo1P2D5HrKyg85x17twbGHhYisSxZ07bPhja7AciBRdJ8HkrgOdDS5b3y026AUs
2lhwnfHM69PoC+2kGxfpheo0tyt3W542fPYZtx25XZnvcZsUq6nXL9iBUN6o7Rwr
82X9+Mz8TlzAqaLv9hd4h0dLbq/yCLFPO3VD02s1CEctqmPLEcHNCbkYzOUK7wlZ
CbUJAY4hUvZmeuc3yQhhcFDdCfyg9umkRslbhfdgNQPAc/QOMCoaDIU7nuoiQMwY
1j28+ZP+cXg3EABI6d5e6zPXlXcPSjSsFHlNna7fSIaGihzcmlAi4Vi0sFesLzbn
G2FPQ6PFWmsZQKg13Pc1E+EPazD/JF9VmqoQXn8zd9010Ck87bHtECeKtuEuwcII
mwVZvUmntkfxBNe00u8t0Cx91Wd4OY5dkhqWCJpf+42LpVLbwvAW1Bkrs0dFeKy/
2Xt5Kg+rkireHW6dHUuf5hhqpeXYTy0bIUhNDLn0sfjLQ8EvS+3FIMxGL+KPk8zJ
gHs988p4w54dPWjrnt5P58Mcfl0w92wGEC6Qq8Z6p6ytHJpogXgD2SyDsPwgdDBP
eHsyrSwxOZ1cg/sYKDuYvzd+3sklJ5dMTZBvzzEYanhu/c6IX9udGhD4RTXKWRoB
kBtXFnyQn0/kIURuiBijkYiuPOKGdeNaE8XXetwEr+lWT6Vcc1qrslf0MgOVZxRM
2nRx2aMzUE6vel/B2aB1uarnI7lRH4g6MJ2uoNtRJ02NUyrRBFkBy+G8n/5AYPNv
xGoi2DJ9f3T36HWYl23tfcim1q2hYcSKwNpif3srChE6inYB8P6TjdYb9yp2uoEj
xcy/U5/ICP2HR474lbS7qTaa6WH80rNm38Tq9SgpgpPJRwuSQ8A8MBEGPgZTcF1H
X1XYFPoaM1SGiq0fSrXjspEmYO+BM77eiuSfxlZ2Yo1knZQwE+F9oF6MarySw6jJ
P/s/setGU+f+V3a9p4kkAUIVj5nafCEy24DIr7FBelh9yTIkmvDJXhxu5ni3zBH9
kmQ5LzKLdmFye8dcM8xz1AnrB+jaTp/7HB6XSkoIw1DQpNcxgLGXpvfYW1QnUKT2
Vz3BLGtUkiZ5qsLJ67QlW+iXD30LTwqTSUafHbtdiKUVRrJLcVn+KQl1FgrrL3As
WaqYDbo/s7eLdLWpEv/KYUCOAbY9g9S9tE1CZAFYPtcR0kwyFzPgFhKnpCquyaGH
hr2T6+wbz93VGW79ru3jPedvvlBiyDBd39e6yTpiYgipmQnKHh9qBo3OSUvZBFym
zOSFwdFt0hdR+thyQF2wPnXd+GlGiVlSMvChMEYJDnLth1MA8+NwY+Cqe8RS2BNN
eSTQDN0J5tlKNhe8zSuw/knn6Zp4jZDgA5M87gIungKIXWwrKZYTr9+WBaGZIHag
64tn3LBswAacnLz2hQBB01Uj8+2dyyCkypfX9maiXiSArQ4yxKcLwyAPgW4TRUZ/
8CJjJVx9fPGvSv9LCEsZ8JiHaDN8k3UlpZndomUVoC7aKgYzlE+4SLq6hw4Mb00V
VHLaKfvGyl2UOZI5uRbLIRj+JivDJvPah6Lk4+5G2bbHz8SbJogTzx+G4+5aTVex
Fr6/AgyMHZBpw2/DoE8FBCl3DW86nAR4B+yzarxqQ0b1T8cLyLgy/ODH3Y7Hts+H
L86fVnfM5nCFcZA7pQT6aJdC2ZmRWp4M3ax0KlN8Wn5RGosVsRe/bapJOm8Zx52H
TBILjJafZRFpsW/U3obQ6J6matIBSFSicso6+SiZRwqFCW5HAYYgMxNxTNbGvQl4
yAltttYvVwUkrwLLNKwoJEp0ewMZ/yOClAq3ki/5yMTZAoLlSF+50xFO9/5JPxYQ
LI91KEMckzbm+tvPKzKSLXTFjyuGpg9ycbjSpgBf7zhot5kSu/TmzJUVHs8IzjdW
VAKeQOM3DwQrGM4BaJeCJoFY3qg6hltuMEAUd0fqDZ/5gsIU4wgCyFrYPecYFOlK
k92pFuvSp+uTfm6T2ckjRgRyMplg7tXv9nWrSdEnNcqHEBMfLA/zDlg4KKEmq+34
RS/xUZ0Jvwuka29z2WyGnnP4vYVmjf8znKm4rQLEn10UWwQGRFjjO0NN0gBDqHdu
Crp++f4A8cXpAcbMSOLczU3SpdRI/12YRZEoViEbaoh0DsWK3Wo+LeG8WIVEcWWB
L/yA+n/Gjal76K5RJUKdX3RKZOlIvVK/dR0JFGShdkRpCEa7REFDJSZ6kEK4qKVl
HNNIambZ560NTEIIgj+LXHgMuQgVGewK3Q794fq5mq9fFBbLCNyfi2aky4kCF+kz
C6u3LuADxso16Q8z6hTqBAW0yBwaQJPt6OZIab06emczl6XI3u0bDWu8OL9COeEE
tAVQ5mCCcHexWTLFV2eSeDFYthlYxgllrldbTuS2wRZYEaLNchiEXxoO7ebgkeH+
qBTGL0wEmugIsZvU/oXPpdEwJJUT1Kp9uBwt//IqRvAUoX8/XQxXrdzNy0tw7AmW
x2r6ChP+m4EBnIi2DbSFWNd3kp9ucDQlAgoPAXWAv/0t843mrZ0jS2GACcF7f9IF
pzyA1ldYZsg+ETMuCgkH/q6i8Kdx8o7jvkT6K9Pfv18lZfwsF4Nxa44getGfPQrH
OUmPAaKE4x6naNqwf3jL1y/4W8uIv/Nv/afVG7gnVoWIdNY4F2SHTtlJ3Z/YFtBf
oQaPNtf7O8FtEpmnQW3McdAdDgozjj3G3zRjJwKgxMJVeAIkoCq+M8LmAI0D0r34
l2XXIF1apXddjCHW3LEh2wtbNtGyYMyVjybuMeFfTh54+T8+cRmhrbH+Sf1S0/3f
ODvB59PnNk/XkBrwRFB5TwiPePXnPMhMw8Sz63afnYG9NfVjGbv96su520BNQ7nx
+Hrn0SGwVNJe/uVVHm0JqXax7Zfcv0dOoxzIuzEGjQ4=
>>>>>>> main
`protect end_protected