`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 27696 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nn7oC/bbltaB6y9f4wbJdgh
0G6WvBg4Flfb54G2gjKn2wSch9mNVw18QwvXVG4GOzYyaKu9QgGJia+vWMMKhirG
5Qqvv1o09hd5lbAOAbt1B8EGN07agjysGENhqHuWjj6uCXLy/bg9BnT/uG8zJKOQ
+4T5V7blZCqgcl8AHjZ2LZ6bnpOkjN4QGdfBf/N1X+w/OXgc/td6ZzMNP/jhwbth
tZ3ERGKUQvIFF4ZysrLNpYQZ8urC0UOWVYYF8a6kSHzyu/4N2OSWkNe3XpVQj38Y
vxkFbstWeVxKuhpaCG4mVSerBwGLvauoCoyKof9ToqpokiNCHEHfSxbb+5VhNe98
dVLYXsgdtsOpYUNhn2JANz5IasB39wC5pThndgYkGj4vgKUh40nxBjYPTG1BHIEy
piMm4oqWzT1Ubv03ZbdQsDfCTE77E0bgdppYvgOHMCxMf3duZi4sR0c8YUZJMUSt
mw0U3Ei0nrpaqUHSIyXaApFFFBrPQqyaO49nsP5BRgpA7sJoG4gYGoYvmERJ2Mg8
0ACV31ZEbAc18oWQVI9P/0aywqxVojolfz1NKvCQfHtwqcyRrkBWVlziCmYnBV0s
5bup4ivg+6im1LtCVJlxPf1tcX8JkyGP4xlHTfZOeawCrOn5N0ox4PvrKGeZMiOp
xuzYxTshJdlwOn9MmAWuOojdP0LHm00WJ7dlnDPNAadqHKYrf1Wnn81PmILU6PDq
g7ZYThtdNcGx/z8DzQ/7L1DFxNSyWAZ4GQf50K+AXo3yyyigBzec8CFGEBZ+51Vo
MAIfE9R0Sj7mi1WLo5DyDA3kYnkAVMl923tCo+MN4jaB2SiHHu1ts2w9U6Nahoj3
3p3eomAJhylcTRSRjUoOfDpQDNUUCl1fWF3Av6V51A+40oc+CaRGjRwu17/z8Q8i
VHq9bx4oBgAarti8gyKcoZWngBvKIPmRxntqjkvrnTNpVMQvV3P83gkJ+bsheJ8v
NvHBpu907BlM5B2amhq36EqGJJD+6eafHNucn0x2hnzEV6CuxyQ8fid/nCYnW4WX
otV4vmyYlsh3+U3qKsIb8JTAmpt1LNkcnZNqS+sJyEZkExh4D9NQvXmttcVq00oO
5icfezcqDByo8lASxOkdX6k46fF5uYMS9Ki4m50/JybPHFi5C3GU4+yzO0379fkE
UZNtar4RRblb7D9hY7UA1gjRkkwd4K7rQEv87EPjtaVxw5/4OO+XRT0COZxFmnZc
GKUsaCx1xNTrNupkmy0QCxmy549exDwpGLGgDCckGQHd6+JcL+i1OTuoJbPlDM3J
uaqpf1TOnqeVDVgdeXsP8oQIVVdzALAy8DJBXBxDfV6ifvg+vGSwmcMV6URMEay4
sfYLcYqwA4Cdkd0fXBI/SjV/j8ABYFt3xnr0ntq3/dISEx1M9JPLXrFEVYA5IV79
yORUWbRuTXnsXHAWRNWOd0HUA1RP5ImtEp2KhitjusqUrx6oLAoUZ468D2T484ke
VZQ3lFtWbvwmYNqOLWiAmjcu9qFyxt9fck7xNIu5TgYSH4fW2QN+vnHdcpUkVwWJ
nAwE0dG0tf9mmJ219PKBHUJU2sac9KP5f+r+FveE/epd5Yc04B+ImshSMrqTnghU
IssuISt8sDVMw5YbephB1o0vs8mn8pRQnd7821wzB48C9zFE2ORzXSCJqTORFN0t
3f/3XkBM7lBEc//NFolNkoB2Zcv3juBQHeagza0zru6Dmh/y7GTz2VEMz0rbNpPe
ttH22ydvfUNkxLfbiMC/Sqe0dK6tS3qxEd5r43DZnIF21+RnyagAsa9tl+pJGl9a
RYKTR1UNV61ryUA5KINhaMUnjMJgAWttw3yf67JIVlUpfyxbRTsSaj2lriMuwo58
qruO9LOg+U5nmELhUeZUZHLsXCSR+zqY0vlHUrm0wX3dKwKf1PcA/jvpNe3A/8Dc
ucSMANHLupOjn7AwxcWC6sRRrl3txL70HJqTIYOJuCaCOjeks/jI+nJnFl47cQBL
muNopBbJvXFotJuJA4GAMGovXRct2FCqKKxRP/lSMtNOZv0Uv+fEI9xl3kh/DndT
pUoutCZXSUZ0ab2xEfZsshFnkYGaSZB77YyHmX/knjapOdUGrCULgopkscKskhlw
AuUwDupsls3mkEYywdcb/aHU7zmMhSVgLoQOc5L4ympETtE8jZ4lqEUh5z6iWxQ9
AKm3/lwsflZWgFWQDGeucp0Heqp/ZO7YWgriJJ4O68CW8TPQyK9wm4keYCjwPqmA
60JhbaQD1yaY+q+TD5G3FXOrQHC2xuSwivZl2IdXxYTEUHOApQ+wLwrVBKP8/5Zm
/RxnGscMCe7rK/j0xUB59xz9+/LWkbAgP8OcCc092U/TqgcXRQ9kQNUPIHzGJ7j0
OPDE6lFd+jDtZcTn49msRXU2MXoq62ZQGjCs3LjGPVY26sI+p4bWj99z1w3G+VEQ
7QJr/aDujeJPWWHCmzUHW1E908576TGIOCJPVGvFon/udN+tnj5S2rvVyDkWkvM2
oBW/ICLPF5ogFz2ecgqLFmZ1Zs2rWuXK5V+Z73y2MTZHhimhAoEsaGCkjGeuOX9a
FVHigz1SVc5XXSrFLhEIKIqbRdTZZby/FYe4dCQTe/ezYvGRhOruMmlkOd+Ztt7j
pNur9pqJxLRVVdV4cQTE6QBizWolqF97SJxeCshpXWC6OJ/YLrqf/0BC/J8bt8Eh
A6iOjos8xfhtXCxK1aM0un6A6xFnzvOazV9XJgjHXVgUSetplC5HE1KouQQZCvlO
kGjQTl9q5Vz6JfPTOOcsa1UmLGrXdhXMrosMpvsJxcuesNaiZ67bGr7fq+bIG5IH
s9n2ruho9G8IzSb4jtU+9RRwsFUlK8tLHZi96JUgIWLAONj7IhpScEaieJM6QqHf
07V7/aJbFiA5ZluBmBrPHwDGNrgecvQku9PSGxWh5BK9encR44XZJwsIoQp1TwNM
1OfceiLV51efoHj1akZ3CoKwpUaL/Hmf8wS3KflZWF4+i9y7ylNnFXjMSYJzrj/E
/FvhGCe1tr9Iz1oTTfm7nJC8ZTGrH+18app625e5sWFhlu5kaaFtCX6AZ5EcHk1F
fEA3ARuvmFIqT6ngSb0dnNobpIaZ04NPsdwXSxVAgkY56yY/f3aTvi3myHp4DeMC
F15rwmqh1QGWONNMkYw2h91rAHn3/JAo+5W9epbkGNumpYiMcSPZvb0HYBwmuOOR
T4Sr7vaZO6XWNwp4VfELOGsBDyqRub90NR2eeQ8IYXjCP4M/a0K0AjoZyvcBL7ru
2khsOTBDM+1ku24CqLmTEeU2TSZrZSGOeYMhpA0s18CbsUUi52QWCVhTjYWq4P6c
1wrNIcIsqLq3fCrT8VH08+yQQyeA4avXdBZncH+11VHaltXDt0G49UvVA5nxyrUL
3gVJQ6UBTS1J/fHY4dnwsJd1qYekr5FfAJbGwWgc8tXtEoyNW0Emsy6Io6chUEe1
S0jX+KC/+BBjMBLX0AZETnSWusOHm9COiLHQFW2KEWJkVBGYB4KDBVq2wyOAJ4ch
9XoMhIh5G+fz4lssnAMhwaP0vv9R6Z1EJKogAzhqzlvhLoAlhGoJ3+fLBbYEUshZ
4jNZmNszVq8d4CpesYDgnGG5SiZ6fLW9ZnPoQGG4EOJH9z4IIzwfBWUrNDX6CodX
Hs/97YY7ozs1Bq5BKROLa3f978D8O41kbVlqYqtNtgz5OslHhCAPnBM6YpizODpa
xPhIez48m9+hTkmF7V6XHz3rjxF/7wd8qXFY9z/yY+SbxQj2p8ckzPSO4PXVq2Cv
vZFxTXq5YITcDRi0qbb5MiSouH8/SqIIzMq+w1vyQJR+2bWPuDw8QVqiHNv1+i2A
oVFEWPmTq45+tfGVO1+4l63gkj6eqKhoAY9/2U+J4Q40/u+1Bc77v9FIMFY48MlF
zFA5d0QP5SKD6QZgkdR270dgJk7Apuu94wiZfw5Ul9PVWh4yus55Q+pWXNExj6Sg
TMZNkAwmKukX6PGZYeL6ZwYpt+QchDMzeKEme1bu2EAv8Fj5uCsgkJv/ody8vpHi
pG+xzavYpe+qV//QcIQtsImzLLfcNA71BLl8/HZFa75DIirTUtu2OJ1hxpGoU63S
DExU/Kfb06LAcrPKyTlgh45W6QawsGDm2NkrbUypfUMqKwm1NqjhcxvBf05RiAO5
Yf+GyVuBOG1lAUBL/PiBGvk9pyEr4D2YkSkRYP38GuvOs+WMFOfOuWeVs6/laJqw
7nMvq+x2QoykQtkUyWGOCSREBf08nFboOUOdEItZfPkAa9KeWYsRDp2DRWIbpkHo
v+FvkJjQw0R/yXBo7viYpj/akyo1NbSBxS5ad5CM11+B3GZ6szMGilZnremxJ8tD
YdaSvsoiAdR3BDbsBOHv31vAkBX25Inx+hZh4hwwD9ysbFzL63hbjEWwFVI0GZLy
MH+4tDhNM2HmMkxfIgTVDkl9fEhY4ujDEtCPjsmJYdfhVKO5pCAF55H+5A/tXg7C
zzHeCPHqhNXRx+PvNzZ5+KKmbY51uaqG8hOTfs0LEvJjRpeQKeF70Sc+0zc3JK/5
LSJzm4IKWBpBnFrEERPSPgWp4Ef7pdi8+g85/vTtBbdOI4eDeMr5Pw696xzpKOlz
SnpbwDpNn3LyGN7vfKn1mu9pSGZyzphawOrbAf7NkPdDbypHbBuDY/sQ2yw73vg1
LBT+yIhGGctmiL9Cn/dtGynp46d2LMLXfRZ4i8MCElmECt0VX+6y3CMfHswwsoUx
vmHuR8A53evBv7my3oIgQIvoYA4E3Od6B3EPHroXYvrYkhkhPeO94/3HcUNkIudH
rJ3UGnUGqx0yRMf5DLeG8oMiQJeMIlfAaPDNY511k5YXKE8MehDJpaX3uUX2U/NQ
bBBzNOhSuWvLUmqozYzk7Uu1yjrzUTiXQG7cO7dehY4kKt+3fNodpYmkihHhyKQf
evUek1pBx9JIt49/QB8dUoTsaEFb0jW9vFZ05Icv3eLWh3RNHycqCehLv4ZUrHok
slFlMpdLAEPcFa0F6C6NrPdS1rRldwOsQL8HldLPs/wkivE4rYSB8jAiATA5tfg1
peKCfjLl8dWB+c7Sd3cTYz5RCU0FE9Bt/+V+lpH/05GDiCIKUGvNWtfIXtvlJBeS
B9BN8s8DLcEIpj5Rqoqset1frV2w4donwuZATWa/VG7XIXYvBAPD7u2//atLyyzg
fd6V3kVitaeqP7+wVtTX6qplNE0tpH9OPenDfITpHvvpyX3wn91IC61v9pCEPMSl
cRWTAez/tluM0YnooJsuZN2eNcpSrrouuUISGDMUiuoAsUnEPjhZkTnovmY4Q/+T
e/RIzFZOcGwNTJdu11sufBTkEzmn1PQY9I/+KRfdrM9srz8Or1/kKNdlEEXYjNAC
jBC8QI6mqwz+14FxrRtukhmMxGb/reSagm7adaclpV857s0qRABE999ry09eKXzq
xTth+agw46hhWd+o6Ud8Md3vzaVYQ6RRoWhdsq7Arm/M/+X8+fy0hFX4/DP73n6l
iSOLjRjyNzedZUi3ECth7z3LDuf+Nie0lDv30dfRICczukOtDS3UjV1BVmHrepb9
f7wC0PB6EKaG0wuZuJ3X5+Xa5LKAOgqXHxiXZXGhYn9SJwwibAGf83gTKAp/shiz
R+449/8YAWVQ12j97I0zO4277sN9onG3LxFvidEksAJIfU5J9gC/Q1WYWbPQ+GS+
C9P1/DmGQ/5XCji9JlrmkfTfOGs8eYA/VT85yxUHnDyNphulxUy/crW7K1E6Ktso
rhv62dGAfHdnJZrqGlVYTuVQSAU49we7bUaCHGyW52C4IHDbeIYuddQGbxv1W5T3
HiIUCj876cAjfJmgT9IybZjk/Ud3l0y6PPNAicSoJYUc5dltPxvpqbEVKRpzDGx/
lBsTqL6sB9UHSRnXYcDsxrayRVyp2qta5ujRbkdlk0NeZP+GZ8dV+K95K7VL0s2r
WISIx4wRZ9aW+CVKSjEGRM7jlKkxsiEEbu3KVNugfegxC5bmRsQUGG85FpVpnXkj
4FZP68Ru+1UOw6k72W435ZnDn36MsfmA4B6lZVjYoSF8QrtyTGnKUt7K/MVOkGIq
3DwhbieDn8vJm+mse379/qwNCoiZ7vmxw+7gspc0VLk3Zv0t5BcpZTOEDyVJiUuA
lXXeZLDdD8wFH8eATU+7OM2cBXz7UlZMnQy3qee0SDX5MqJefijtVHD3FkntJYwp
0PVQoGG2X6bvrly/YH8pG3tsBZo/O6Tt2wrQnMugEqc65gYmOyFUnaYPuNcYeAZs
T/j67efXowR1xCuodpYXO26w5YL+eR2XAgWQTkN8t0VjKQEJsnVzO5GeVSAPqYAl
OyO/KiZOBvF4iKUCQBVhD11fYubshGUtJFD7wBr3mIMStPNxaaQIhdfJ/CIt/Pu2
G1rvjWHvIrsAnXrq+i9BnlGGKIQgoWFApFtxGMfiyrNxJrLF2YAf/r5YwcvCLzSN
hrSf3aslbi/d6YehjPd/MO/WlkoktFVCpWkPdhvZGBXZjROOFZ2y54TFnRihVbv4
E6YsTcRZf7TUjpx9QYTB94kR8k8PSDAIiX9u17vqxt+CpB+i/TJaYy4vHhZnfkAL
5b6aBXPM/N408tVhJwaJjnUUpLpaC939zxCMMRfgPixa4xhdyS7eYH90u3NmhZmq
9bSR4W7erfnFFgYSw+IJr0lsIGfBPRdJZ0I7D52BMye4fSiiz8Fd0VpIC+kCjvyh
N4vcV7RBzZFkZjrSpHJ5ZCUlvBZ29ZNNZIGkuXKgQ/I+9QGaw7E7wu5d+7stRI7u
xOeujSqhRGpB4wPuImf69nVwn0Zo/Q4wc6ItO6gaXCB6hZyZzSS471kqRlzfAaO3
6DVnk19HZiHAoRWtu/FA8c/1eJs7LkEoRR+wyltgU0n/lEP/x4drYMayoELA84Iz
qG0nRGLTnRLlfWjCsX7O+uGq4niMPkOjR4DRCNLt+VBO4zRpSnGOqvzUcbj3MkU9
yx1RrWBdKPKp9g/Zoj/tz0wIyZN/gdT37sNQUgcOQdw6YoidOT2uSaP+4qiz728m
BJ5TgLAS1vXCJvDkXww/CQiul5ykuCQQNo+pfTY4/w9tKgUwBs4IDOrAkIn7X+qw
UMKsiiehRuFAFtWdeUBhW5v8na1ZIKjMYc0EtwuyQWfUFmGkLbO2FTBMV30dqXcc
UbB1hqnxd7aGUETk68YHUiCpG6/k/T9HajWEKHYu8MvzXlA3AW3zOdi1qKg2RqFR
Y53Th+BBTk6fJKjUE+dKBxU3fW0s7H1J3t8vv4j/P3SttJjxmHrb10bnfurPBM+7
W+oWa9BVwoOIgDNBNh91IYt5rd4FxcWZpbJ1NyvRohucAqVLEIULZdnpfJioc47s
Lx6Yfs0yOo51ljtHskbdxaTjlNGUsoM5+AATnaiatFaCizh+Q+OIBBlic1AtTAhY
IGq6OBeQ7zqs1BV36G/U5fmbW4YEVH/DJbvKa22nyhaGsqZJnKj+jygRgHGPGon4
gCmOK+27ae0S9pdnCue0yyQDL6dwZqopZ0YpAsUPskqtAKUUkMa9uWK0TUhiDyCx
OyaL6jwky3xRoICS/nWhDsaongqFMZXrzUQCAXoSjrjWmD+sM2SdJf8nqBj3/U1E
Uuslq0ET/B2htoVaeToOpCVh8UpymsCR9yJFGoE4IBho4CxttMVP5e/0e1VvqAAE
a6s2++hjcAVp6Z6umyJnq0oeXo7zvB60dfZJ+ya7aiKZIvhCcez6Lx2qhpUvOLkd
avPeiZCggfjg7hcVZcXrMYznk3HMhyyIF+2C8E32VGRpnWiA+t9iKHQpVwnNkRNx
A0S9FKr73cLYN9JTDYq+mHptFUQFbXDcVWwB6k+GEieVNKWI4w9kHwQIyCgqRpqD
0r0QLIOO9uGFvSFIpW/4bBwI6xKUzKmaZkZH1UG6BlRhm2qemcfv/YUYMSKwoUHD
omER8qExvr3RvoY1AjlviflaTiee2Z/Az5h7qgrZSEixZ7G/HVv7/jXQHqDge8Ry
AXw3MiDsa7Vq4xoJ+Dr8gJ5rTss1widGXPYzcvcAYnW+4m3qwWaB6391p/hP+p8K
vv/zZOzHL/fl3WN8AXmL4aoGJfvDbaVPHLebd2xoU2SB7r5q6FbjhgWT+H2aeDeI
RNzL5x6RHygDeUfwDP1lSgt6OncJKlzn6cTZl/O8r5pnmc3ZArL8/7msvkEM6sYG
KclmWLzEHyIycusqWeqUqEPekekYRRfElo/OsSaGTX6xq52OcPF1VbQlAXXUa6fu
E5HGPG9luuKFIUYuPTt0yYCQfdKHiFbC75A68pQUDXoMQ5pSxoLIkhBFwZ6UY8xp
Cp+gjYRpB3OXhj2dRcrKTUt5TSfGs62XwpTqRvV/Iq+K2N214whC7tIWFxbGwTjn
9S5vfmFLvQB6foMaWOqky31YsZwIiczprxNCeAZByTi4H1Z4dcQf5UiYHD7krt+k
rQdkIOZxq+S/XYiNT4wAtRf01/paXwXSUEc7wbXJhqb2OMXntN4N2k/k4PFRmCSZ
h01sCkHWAa9eqNW2dIL7pMPlbd7QgpZh48m5UI8bbynah/AFFL3adLFWBEcGs+uv
EhFCp70l5jqdBn80A3Bs/rvC9HQ7LKd6kKc+ZWr9UlgaO5Td4VfFjjV8ZIrn8hCr
pVG3/WJ3dq1w4yHthlil06jIENSXTVatrC/XXdzbr9DPqFUxDwbzsiENuM+Gx0hU
sUhqcOkCORIz2xokVc019OLPwQ2aDgaJs1YxysJPgYcSxizp9/Din7Wj4cNJmOAd
1CWxl5SOMAJMAzsn1lbBbVt/RlUcyI2URcdzR/UeBoKpvw/WjktouPmFZ58G6cG4
zZCHn/UlVIFEkrk/957DqpjdDf4NUMWHGDUAbos1GEg3mtDL5Aex4KrpcQGoiQtM
aKEos7pmN21+n8sPVp0mSwUwNUiOfIIgzRt5v4JmGCvb5esdUrlbHCesA3M7wox7
1xys60xfRyM7J3eeSIQne4BV8YZZymPgUQq3nN5LdcB6xpUONUh6t0vqLF2hbUFw
OWNAsY6Trc8BfPthyin+0F9WaZ811N9whFNVlb4vMjYykyNOn7whYbvNRMyLu318
iu/2WWoY61DEmPRAmbe31CymfoEQf5A+HQr/BC/fsLEWNIRwPKDd0E4O4dUyOEHn
3nZ7+V6S5SHSSX9Kf+yepOmBdPEHvUQ9axpYRAP5OV+yaEs01KCp9xI6P5JQzv+F
UKBnKyf8Wd/GbvUWsRCAGtKaQq0mP/5uUphwvKf/+suwxlp1qrvShcK2WeKr2rFE
1lWWpR+GwIirm1tjfiebklkvBoR9J5DbDh+T7wKzwaOxkBF/IHpDs4+9h6tULKX4
TOXnlSX0dv+OTLrpcF+qLH2IhhFbQAGQmCnZqong2Bk8CG5ZKIh81HFrjzXqP9cQ
CIXfe/nM5XMWLNfiOLQnGzgSiTulSRFZ4sUDcu1fF9AIRKoLnNbx2tUw6K++AKL/
rD1CNVrEWrig2ASN/LyGlN8167nUti4Ei+JoA1MHS1YoX7a5S85LmxIcKOEPDvTy
yVXpRzoQhh0O3cJGv/INaJSn3NXQulmFijElffgRXYq18uO5iEkitWEIanBuaU21
ftRxBx9haegQ+4GmasWK4I0qWL1OO7mFPAHYrdmHd0tfeINeNgc/llia8022ZeIm
x+9XiER27TPwaJCO8X/KGsVQNHZ2iEhJGE54MkjYS4BV2Y8TtSttQ1DIOGe3yXYd
uB7sWaSm2yI3ozljaF2453OT5cyM9sCar8JbRjYHCbbln4YW7x/wYaGLtm2vdBHF
qvG3bPg3pkxqvIbyxdSinW5FPl/j5QQ+/8VUPdmWGTwzAGFD3UHLiOFYGWB15Xso
7MGTMyDk0nP42HVrt2yvucqHN9ukT/UECgMG9rstSHhRYckHhWo8CMVYThQqEHlD
GV8bFpMp62L2iwS6Hs4VKRxYum/QkCQBmmOXsFtL3XduTzb4CJI9/y8x5VblJBmN
sMV23cglKZnZiB/W3DwNXqoeMKQaGUrczNkMVaPMEdWEEX8YEnJNSkNHHhoYvPTR
iotjMg0alqS0cVGwl75SeFuWHsgkLvx/kiNEsZtp3RuhFi+lE6eTv1G0Cj2vp8E/
iRnkP7YN1S8Tq2d3WLLW1Hesm6eYrAQYV1kg8npIdD9dNON/PYx32OW4R+h5Z2tZ
qghv/11OGeCjUnf/lk8JCAfGCmsLd4LgNEdKRHE5+qHnd9vm7epORKeJpz8X9xBp
0ERpXv+d0dd25hpmb/0QUbryG788bHs+BKs8tiK2pAXbSKjlqOurufyCWxOK37da
AzQ9GejeAoXO8EwMeY1G1H6h7to7qag/MWZuS2h6yWx6U5yJWCL/CPOzdVMSIb1O
dXILpQyD3U3R07eTLenY8IRKjHfelf6yqCM+i8orys5ONV0J6HfyyPDr1UrvM0lf
uFX2ZnBzsUB7EJHsHsmBzxAJVEkkf4KWYpRanfNxRpvlz7HYmLh8FWMESvSm/huN
2Vz4yVmAxmnAg5NFS8otWhEYquZIQUtPpPVs3d65NT05MxJbEoAj+lubNKHxKT/r
6EW8j2IaGKzbRvt0B15goBJ8U3fo3nyNd8/aoEkhKasjnK1vHkXsT/QfkLDU1uwz
MVLACo7w0eDXJpkovl0SXVvZpfl6mA/n9kVmOM/cXR3clyk4l+V3t2oA1VfLjSLe
GUbqKBv9xhuCYyeHQpvqIsG4a7Ens8K1KajFsBn+p65AEg46neTl7I16KLM7fV64
Rl/nLIfsL3T7fnj8FCN0dIK4xvGlCGTPjWRdr70GTcNm8WadVPfglIXD7IYxe8JN
nGGEV+nMiXoTU4VI4rn0o0AvZexq7V1qliUp+OwCw6OtYxfpwxYtS70oysjcCW1M
HUnMglUPtquhB0EMJ6BEHqGvD+MBqXswLpavw5d4FK+7BEAcrnj4zFXsACfKPacy
kIr4ofEcHsau4B5nas4dwfSpUV3ISpNMzv6DfteEZv7sZLEiao2LEBSNFFfKdfK7
5+TRIccoD7X8pqwZeO0Oup0er11sjX6qdpxNtyhMvW+1YUUzWPT6hmbKC3E6XR4w
TvhkEYejsTAzUycuZxip9SMlY82QsDG1jyHkq+6SZ5xISnZC13esXY+L/bbn/0D8
QqoP31xaRQCwBfhgqeR+AQq6514co/CQuva06e4Ey9KWFTI9IEI5q9xUisNSK1fx
/4Qf9O8AJ/FUtwckZSqx6gvsgKsifieH2esQQpzk9Q1uJ0GUOQgG5VHbOS/wxQsU
5ToO0hxZNLLOd4pKX/UWxok/niz0i9GXOI9Bvt7zWfCP/IBz7MscjHPfivhibdwW
+Tx/tM4hEx110TRJvAEuD6aLhtgYbn8hHOpkeJLLBATaOyWLREnk/BwNtMZIz3h8
Yc0GVlKhJ7N+zztXUDB/LgaW13BM7VvmSVEOnC+si7oy170Z2AyYrN2x8WIxD3GC
+nENpCH1tABHmY3+2RGYJbS2XESfLQkmpPK2n11AW3O+5OUoy3sR01Qn5sboCEEN
JCbuUnrepuqedG9+VapWRb/+WZQ6jzphIj2Ixw3u/eHKQGLIOJ2qLH+fcxGIEjz1
sZmh3K+9sBY4SCFhYqH2Rh5tgih/wWzpKgiR43xYLSxVal2vtc6tNCqxOoKGUDHo
ewwLgXBEbU62edj5xoi+ve7vPkM1cwhRjVyZjyUCSq7PIVgK/dyQ9+LygQmWuXJU
XlZILGmHt9GwBmps977KyC9BKUwJoT1nRdtAc+sqsrp6coAUvb1axywB4hufPkOo
jvPAJeEMOt3kPcrXdk7AqoyCpFxu5FAkslHW81G1T39lOrukO+CKVmWLbryq0KT4
OedTsZ3xfZmlHi9E4UMJSRv3AIRKAAoD0+lPQqs6XA0JsjaepjGWiFEsRFINwCb1
aPyy1tX+m5JdfwtZVm7S4xlBuCMTYP2MTQyvNOjLoCiGdAXgjDKNhksBJghAv/Ej
vhhuxnCWtJarMOHI2R+gV+s/ap68aeG0WWJM3/GgEnQ8vuP0LphRxR+xUo7hWBSa
fS4M4oebMh8UPWUXQF+5UK/t5235gt75uEIrVffo/F4SKA8YnUPkjqTnG2qD7y3n
4Y4Qa2aqAK/TBnQnvj8q2B/wG8R/2UckmUtYqydt1sGwQP0rkpUtgLw7wHolZSmc
1383UBXK8psVceMTlHmFpmYPccxhapNfyeXiFdln2lb/5az0rNAzucENgJ9lVYo5
sY/PsJuIqpnPqGtsy9Sh1TPXKyQ2vI9rHMukwKDjaezuykoWAWuQsWX5cByV7pbl
KyjbYC7s7TRO/nmva7gWAQQ1e2JySgMYpS7AHl4Jz3Corlhs9g/SveZAJkIvOQip
TyEmEVNL9IprUmoj+rYEP+tKUha5PuyjreluwdPntBU9EuLYMVAjdtrj/IyoA2jF
fhIA22vvRDGIHwMYQp14BFogWqyH55yF9+AtHa0eN5sOcjUtEL5+aXi1DLlk5hF/
UmU/P49uohMXhZgzdTD3ZWY+Ox1jorXsboMBdGxgDveQdihGpB0WXbeg86P0u4u2
31w3HdxenFxKRAlTHWtSUZULKsh5trZumG4pkbob2J9DBYeiYLfS7DYwLJoE+E/p
y8mvorBYTyRzpC6p+di1Jd0UVVPP1/j8Qu6IhYpEboE4MK2TTtQ4HoICKiuCG0tI
ce5AOS6q2EgxoD8M6fEr8NKXhkFV7LoliKqAjjMit5IkMq2zGF3JTQZ0Oj0bSsdA
GOyhTK+TNKLbBAsX1ypFuaVXm78+zZEBd0TcicdkGdVkMb22veUR+HmFxPOGia1P
AfSat8aijYzG/kgAlKoKaZNynm4mpdO1tiy6EJKfGavAtl3J5iAeckzXVlXTrCe4
hvtPrCMN+163enL2dwpU7dJ0cNIGiI44o3UFeeywgvxW3Z2OINmRXmv6KrU1buqN
JZtnBNOpLSndohKNcirpHFx4RTZgiKDm+HFfCGHfHt+HPAAIgWDxD+rYzksxkfuf
BoWcBBT3EqYeRxY9KovgP+0ujoKN5+zrzM7bI3SM7iddpdNrfJXsJMv3BZeuBI8Y
52YIZqd2v38Y2UFbkT8RvjKNVlYtjr3w0A95IwGQp7BY+yZ83wxwtGuU4b3mr3pT
48igLVl6bs1CHe+wy0B0INvAh0RMHLYaxmM7CvdW4d2jbXphMDThaef16gagT4MQ
lssJOP1QEtxDfoMccRkXZ6VUpFFvyyrrTTkQSEQVvqflkggxotY9YigRfmFin13R
98acDikUDsUAx6ehIYljD24KD9WEFXiePzBQptC/6rvMmi2ps63qGVNHdX/+qIy/
WpXTTnZBRh78yErWhrpOEyTiLprsrybFWfTbUe21ki9Zop7LnSOwboVraFmgMvVS
xw1uLr+nSWMqNt+7LzYrE5Y4qfuHqouvNWnUfmxg5HoGzIhrrAJxLfKwoSOrGo14
y6FCWFa8yw1P1Wji79+SRDHHfDaS4AphvFiqFPOGEhCrqxEGXvTcUQa8e2JKfXCZ
eO1QL3iLxSgJg3rC9qo9kOXOAk6qY0m0s155ZEXmdoNKaRDxGCRjap0h07B7c1ix
UiTF5Ec0KTYi67lx+YlevRGMYb6dQ86DuYKccykKUIlOTRahejqYeRIqQK5Q7eqg
FDN/sKtYzywJ6mSRChUMy+KkU5GGDfat0fG7J1ZCchJVwXCJTN139ukm/0HvHxyo
LSabgep8TR3U9psRxMkjHU61GVj95jpTCKdqAoy6zU3rDukLmTNq8SKEYZfvY6Gq
Gya1EGpzZZCMXRvdhLruFfhxFcu3F0FwjUFL0Q8k+kCiGHXkRx6An47Aq2Ij95Zp
klq9aJ/EOV7OeVQjTIlCamBhqfLLCZxK6NqRbXppIw+uolOnzW8pL8j/ILj22XfT
5s/JXvcNHdXCnrYYQWN3a1N0w2eDnk/GOdl+fkd+PzCu3Rp7616YN46zyXlDUEY+
FoJnelWPRuKc+bHJSB0oVBuDe9IWa+GRjmwGlQv3Wbq033IO4Uxgmu7hSfRX5J+5
bz+kf4+E/jzWuLLxdMmPHq7Fk9/uDd+Af0cAdlFMB6o+AC7cw5Lvab2NPrCP/Elc
4KCoy+7krOyTT74fDRj44Eu9F02EK6IerdAosgWsw0ZRgdMWDeFmI02vV3UYXy9/
XDNghvFaH5e1JWCoTyhzQzkv8E91o0tqbMwcNWo/70mdbuQPldtJHn6l4xtDaMAD
lnE+48ku28VMi0hJKYTmTJJDFPAF0qaQSyMXY8Xry3lDyOXBvM5M4adVwZyQzsqO
Ffqs0qilAUDBhHjT6Bix57p800lpP6tujP5OtgdbNGkIdmXj2nCKYN0CYi+uP24s
B9dStFZQAPTlyaZGyLnKxkjZ6Yco0yWsD7DpEgR5uBF1/GFv1YHniMBKcnzVCjkM
QT8957kxOhlEm39V6TzUvZXAidOl8ogL0/oNDj7Je4ARTX/G25oj6A0mkWlbfYdN
ewrlLDsH4jGM6PhntUt04jS5qDLZI/YGRH3NAqHloipfpih7qqS+ix5pNy3GeOfx
ikB/R6BMhqUbHLZ2KOvzYXmOg+BzWcNnF+KivXBYcxUyNT2xjL3dmyxTgqTL/lEz
Xg6xCnWtSmgkiQuSjTDxsu1PKq3dq94fhwiE31k2qiGhFt5OPYgBgDDA+mWUyWzC
VdfW0hQGkf8AN4CJfLMu5e5zsEusUWIIGtBJWoGgucO1D7Wk2HVzMVUd762GlZS4
iJbRDPKCvc2igSL1ZmwBZa+cjAd/oMrKXQucoBv1pbzBcuRXE78TOdockng8dzdb
MXK6dTt+Pwob04hgmlCQn4N15y6fcux9L9RGNG+Cb94aqMJ+ahU3duekTBIkGDol
RGY5lCM3MQhvMjSN0aeCClb7VSiLyUkrrrFV1kdcJ7kbDYVKlSrUPQRIqs5z/Zho
2o5dx0VW4ATmqDXlxhuP5CjhtdfFqxkz2oc96v0id83FsztrB9Fu3Nn/EeO9E8f8
8QAU3bqlLt6HZ46HgzrsU7Jz6Mmc0UBTflW5QKFvn7OWmzL7/OK9lOAXZD1TdMqS
LdNnxwXEcmHO0MDS4WykoLuLGBzslmzHguINySmD0y9/CaKyZodzc65UN/q91q69
RBJz95RnDcj/PF8XmNEVEKccTpxK6zY/H4c3C9LpNJpc3HcMRBZyVafylbF6otAT
71y/L6UcehzoZdWMVAlyASVm686v9+Y1Ndqnb53im1s9l2OSwyCv2Sxt/5tmCAsc
O1SCr0pBZ9nha23SIyyIv+bCSuSWTmBIMTdU6+4F5i2xJQQjlrAxEnJ+tnNTTy3g
VeCWXaVAECQBXyGdVvuV99GV3+QqM6AOPLIikFlH85i9bLnBTMXDIIcmXouD7w8B
SETmSM9XghJn7HvlcLcU0AfWIZQHKfY53xat0uU1jsmr9O6Z963RQc0sWVk3Qcj/
TaJvSlh8OnNMpQpEcZWmA8pBeDYzEGpERSckqFLStN4oT0p6rRbPHhQLt66RJrn1
wvG9bz5NVjsyXd5NsThpJeJyHfvaM/TLZmB3znvVJQwoAcyzMUJu+UkXbCMpF2t3
YCz59ado+xKJIJE0OedLmHHecd71bKxmph1raWA9k0lWuAEsnraLffLit5RzsCJ3
UhCfGibzKVYrNqAzwaAT83/nwTpEqtoPR+Glx6oP8KGIrQETL7eyKl1WTPr34xma
pB/BBVsz0HDJTtVgRkugo+ixSUvmMyRKsMSLd0ioX28VTu9qNtP+0utpjof8R1X0
dJf2GlUPYlBeYjwnFfl/OcP7coNUlemokKG3okYRaZAfjAUCGDY3yPbFahHblT6d
18pmGerj0nvjEO2yb7vgPil+Sfu8FfrMgXESQLwX1xHc5i4ejjIBuJ1MAp3YFV3X
ywr30aRW6sXTae5csRjxOABPQduIY6jP2vULpslLxY3PRnjDD4tWc+cMyDs6Al3Q
4cIHqlsNst1aA8FeW/5JCn4lYFf6CbedmXdyvYRMDsbNLIzfO/tRlsQejeKdjQkG
ANdtYgysPQDbj3PJiPn/ijtJtUBPXt0rI3W+Y3lKzMRQDsFpHSJyjTqVkX0Dsfob
n+lPh7MrvKtZ/dETKT27k1Z41PtpovesbpUsyD2UfSflVbXoQIyy10rbF+5wuej8
d2TdKLbiT4m2b5Plmn3bcAY31foOyg/xZv9Sv3YgnvZafBtsRpFMxUr4ZHxtWeyw
/HipVPnNW4lE6CnaHQjSVmnWbvzXYr3rRwd4Dnqe9B1SE4GRoLVKY7dOJ8dIOYmX
HgGx4s4cOvCa965ukZe3L1pxBkb5l+awiBCYL8AriCZ//oQvGNY1giX0OlGBVr2j
5OyGU79P95r0UAqNiFcPKSKV5HLk+k13RxgJsuehOHL+icmPSbk3coL6O4mBl65W
SIg7bDEofsoPYLtGgEr7C0JCWOXOfquzwqbny95jaZHldSZ/x+qFOwunvG1eETqU
UTdNncPCbvRK5OS2gqmDiouVuQc6exmEmrIeejmeHusVUL4Hd7bMWjTwTvo/0PWx
R8zZLbjhRnTRFatRJEu3siPYI0/W4cdxuW78T3BMsvVDjMjtgjW0f8jBidw9OcKf
oUOo3mYkGVxc0v0UhLbeRvTT0d9k6p2KtC1wQPQe2rXYs2l74GJbZdJCUplg4p03
0eTgm+MSGI+qZ5n8Z593PmIS99orQzpL48wIvD6qrvZWGY1aq44eZTBw1nAKqt+S
MIGTrci8Iu+OfGWrLXqmIA7CBLS+v4wNIiZT+a1FpArPRGXjebkNPLgbL69y8axg
JU/NeoMkyfH+2LE/NqF7I0W/1yRxv9gGrKY81Dxtoa1sNhhwt22ayPPoOIDLb9gV
PFU1R42iqiGshxGeooVIewywONeSs2pqpoPWkT5H07okDFdpIVBzimhQpztkMVG5
yGjo7ZxlcJXqyeOQTfQUK1xA/1jQLLdUxsYHoeyV2TrjtWO50G5ueRiecEA2VgF8
CSeBerWQ81jpgLaJFkLzoCPQO/gzzRDsh2PnvNrCwpTBIiSGTPwuJchHj4YTuQtd
0BLgXGtsEPee0uQO/+REfvTowK5yUt1GvVUdVjLw2BDtZeyvDhcN7YGPLIcibcIu
UmisQG759VmojiNhP0HdmYz8xDlLQpwfaVR5QaFRXxsWldZjdIu+CV1q/tYY5AD8
a+3F6NYa3zaS2tvGqy1cDB1BiqHEIGiI+Zu8OEzNFrudphi65s21XXHNwx7KK4Qz
CqdMqs9fiVeFC3tGRhJ5XC47OBMX1s/Y+h8rIGKKtEqGB97KCmLU0vWxtf2kdgAO
vLcaoBGT36U9NyYV2qlvuL0k8ppHim3k74NdmnrkIl8PdneO+xRWv2qTq8le6GJ7
R9PxaHY4k9qV8GQI216FHT4dcMEEnPTQ8ccjFMfuKa8C7TI25TuY2lwg03/BXSO9
kmWi5PR1AEngpTBs06SyJdwtvYod3AR6M6RfwtaUUKD9J8e3CAAlhGPI5rU7sX5i
2ZtoR5xerHhBrQIdCbBWJ/bcz9+2XXcqh9VQL4pPq4UsufmukFyEYM+198lrXQGv
/ABVi/uZmtI4Rq2kB5+0KoMQBakqTGXeJxhQq3QVN0AMOVhTMrO7gUhafBoRWynM
NOaEa5w8PZI5DdpOHFegIcGSfT50AEM2SmZKbdwNw1GmNj6s9YlGUD7WY1fm+ncI
G0xZGezPIhNqdr+i4OCJDGgD+lUESusYZNIPuCJdWOy2u152gmYbr1I5EbgcLyYC
WRbbom0aVMb7BbcLaLyDWnL0RKKhDhj9C3oDNl3tzS26ttZmGsX1/81f9xPHeEEg
5oRBoyf2c8UkLQD//+CXf4h9ktVe3MycpFtcVITvHM0BGAW72D5J3zNg9buu/8NF
eJIc3RzrRl7OTZxvXF+Ef1DIE3fOlKEZjrMh8KHKsqG1N/vjfW65BQNZa1R88ZIz
grEt1X0xXX6quNYwd7zSrHwRp9vSRTxhv0p7E14SmaU5/SMuSM/yXbRoXlInaK8n
t0LyTzQA66Y6XERkNI9zqdUCzOBZzzNMN4TKOwm7mbS/MT5g7SsVqh3UI3Gds8IV
Bs4jvF9itMgtaUdSP1gfKp+U4AQt87ssjjOuRsI4x5jh9Ua5ZWn0A7299f+KSKYw
bIlpTFMU23cRHw80sGwUHENKiBTGBr+7ZNkRqX57cHp4J9KrZzs4QqYw8nF/rQ85
qL6H4KrPiVwtkLS0lpm0RSQG+uAt6nzgGrr7LDFAZJg6CZvuNJ0jLNKe+791YZgm
1V7uTU/OXClZK89BxYZsQZJwjMEDbrQZEjzZzlRDdBJrkXBqCEReyXwv4amAkhTY
Bc8Pn0/5isiwqfnPg5pM2M+U+H79fXwYYsppYKPrjaFZG1qrYAfwi5ZN6Wx/PFLc
BF6ENXUpN7CXVRnxPNRU+KOuFYoNVuh27+Dp0VIbUBc5MlD1AvOTBN7q7CIgXCiV
nXpyHOKGvEBEzLFxyegZMk0JjseNds7pB9cOM9Ph/dXVnxM9s7Op5223xxcv1yAG
nn8Qj67PyWAu6MCfj0kqIXZMzZmfTBVk+fQ0zRXqd2hgGtOtNhkXnM8+R9FDFX+D
7DINBwcgaUeSJ3IEu/vmNmBqJ89AaOJ69QwlxjD5OGMOArQLqTn482stPrId+p+8
W2VA/IArtkefN7pMCPbhR4wrVF+M8fpu0X+k9D/1UebtLFKi8ObLmbEFhhsuMz9L
FgHWRQ8pcpMAZc5JLfx5eYfSmUoRGlxeAyF16daoVFYqPuwf5XKODM8V2KP5KrnU
PmaHz2JuoxPFGHgMFtytHS58YxwlT/VVEgqoNSVAdf+82021n6nCtAGB1F/Ozb98
8GsYxAcEEN1QZQTN5hqPOwRl+Put6zJxkCg9stUx3PxIIDR7H/7ElJ7OBlVdho8e
WePwAowoqi0Sb2gw7FPLWBNNwW3R0z3s3ZsJ6EYPXmaf2+PRFYphLfLC8VL6Ibnn
ipp8tJfJBzNp2dQYWm3GrOl9GxFsmXu6lSjyo+Cdh2Caj3vryOGbgS19Si9q8cd/
SNyT8vQ08sE466fBgKwhkIBeyjfPnP9MUFxjS4JeUTgMwBTdcJCt6h9E1Y4UVT69
F8k0PwUBEFakJNMriwObNmIGb0xu5JFOscjFC5lS4CzDsH2UkOHg5sPdUAtxuSqj
27P+R3fXlDYn9ay7GlDjVPzu68aPVOjThvBGngOHuweFmgyKlp6Wn0Mp1aV6/DAt
JjIIIGAHEudEy0eVY6UDwKAHU7nO2phQH40EpsPU3vhKNHHn34BvJKUSoPc4lmI7
yLrfqtYDJE7uHdmcNAlp/KBKw0z417jyouqw7WNj+f/ubp/FisyV/RRfYmOTXifu
45aLJOoSN0aLSsBueHm3g/aNj2AWc38RQjT8k89lSiX2fJeKInq6qXA8YoxRmiAL
OeSsn/mF64ZWGugJAk0bE4Iw/dwV2BkJHHhf+hdO0wDfanjpdTv/iWoYt8LbG+Al
fFR3LGGx6LN7ZdNk9RCZ3gWjAc6cw5nKV1K3y+LW5JSCmsiK66oWiE2YZd79XQ8J
0PEWX2lNgnUfpj1cEAwzn2KOzEvPKA1Oyt8O3knCj2I6Royf1uuSOCifz94xSzjk
2DlshmbZ8NwktZW0Ewu6IWud9LVrQ/Mb/AK1OF05Oh0G+BrLGR09+mk7gF9C14Ih
hc37QV22RoCcGEWzo3y3DQCnJT13Ep+6sQQwG9FRhf2x13wAJXyFHA1cajPlkRQy
/J3EoxWGkKlRVg9rjRPZfAIs36paX04FSoqN4UZCna1fzE0eIQ6HOD/GRttdPCOg
uuvbl0RUtk0qZoxP0dhSrY2wpf3j11EKPzDTwJ99tM6bfy+9buk5rghh03O5+YHb
BePkWsbeEi4jgttZ3pytvi4i/3Ypzp8NTAmA6xaD+lSdu1gd+GXTsdE59eAZBIAs
Byvm83+AJGjuKmHvPUuDoOJOK6Uoef8Lu1+A2gbhbPHckMj8sufc5W19ZYa7IJNC
E6k9SHH5y5xPlKyFXbQ25STQm0Y5tLteqhey96Q9sbdw5i5mP/LL+dr7TiwflM0W
ebylwwzM1hR9JBi1YpddhE4tuBcTiqf8SrJpXNrezcp84Rs0nh9yLaLDUF8/xquB
pG2Wgp+yqUf7+HIxRAI+RQehZJFSU3kHT5yQ9ex/hLNI3jtabJRCjpD0NR5sqMAZ
meyU0A6jgkUK288OQDzGbkUMHZQYJxdvhRJuRmhZkwWUonvGRZ8g/jarp16FNesj
2QymUUs2s5+Wb/AcKSmx0FzGS2RwqVD+6SDXld/O6s7+8DYtJCXxIpHhLR/x3EVL
EsBbs6dvQpEsvtHx0JuA5WNMmTMFj+4epNEWP1BVrZjx1uTy+gbS3EBwa07rGaff
nPcglEQwa9D4NSI8rpHF75TktAL8JQGtcy69uC/otH67E26TQTpKn4VpIntyujT/
cCN1g/NH+HPBqR+2iO0j6vBJLm/atk4MX2PYR02KRE3OHaf45RsEAO66G2huwvyX
V7YAfTpxDsZOqqJr4kMqPeeCV6ldxGRVVhfJtNPN+pk7RwGVLDHV/5HQIXlXAdoN
8sgqOA16Vk/Tu0Vz0zYyWQDycSfFSMYv18nvLq4u0ZHmggAXymWt+bot8eQW0/DJ
IvyAxxNdKI7SB0hmXUuGkCMHBONAvmYDNrVuy44tXvnbRTOjRmPMevlADkYW7YhO
ERrbiQBIUivg8m1lRPh0tzP9q5W1XIghkIdhc0bWwNNQp/2w5T2CQUhrKjuaVShD
WN8QyL/FOVSKyEmmF6SIQbziqXiuuPEoNDIKab8kRdH09xAEtuBDo68KmHjP/Fwo
PKLmsXwknVjRyw4lW8T5LALdQm69kkICBQW0nVZbSA4MI0lN8W0vgcYJVDxlAeEK
sGU/iIKRAfbDPmcn0KB2fniEeKtEHuKrytosqxkoPKBt2QTIauJmt92BVq9jPh1v
Kgq+WCsYtercXRifXVgS06a0n/PIGUms+DXKXnHJSsC6OoyA0AY+K3/z5MvS+rxr
Fu4foNbbfn120haIVPzjwFibaqY8UEGgtDBqMSLMAAVs3BhXcgMv0QHEX05kxlM3
qqJRUlk/tA7O3+b8Nrdn0d53VI3pKAxOsvnVPUovh2gyz7rlromTYHIexuS4Wjzx
0tR+9X9awLFCRMBPWNI1iGhX9z0lbD6V6IyTzZOKIyyF3USkilD8JPDnE6mfMLiz
70QosFNQZE4UfCJhdeTxanV56q2y2mXPRaw0BvIZo3txTEPYBzHGUp6V7K5JB1K5
njkyyss9Ze1968YW+JVrNjw9+Ad6aBViSlwTwJF4k0xHCnAtOR3UYk2PQY4JBikE
9Dr4+UWZDtuusrfiWUirTA4GeqDnK079m9jzwXjYa6eAwhlIfV6L44+818/bJlxJ
tzUeOPqV8dUWMNqmb+4Oa8j/17RMAY/thMAUWp6sBgE1+tJhH4cH+JvyQqBcxAEA
O0P0yu1xucZzuqKG25cQ+ZjWvoDlEYYL+E8dOEqIbrfJ3MgSCacd1zVKmSL8PBoe
CL6ReikdzdgP5h2zCBaZhgUPd6V5y27cGc3nGXBAvXs6cU2Pi6Hhm4WBt4wjeLz1
3fJlyx3LfUId9FuoewVcx2yQKZLc62mFjINr7YQjFxN1gpvpIgAFGo5i/BTj9iIx
1Nqj2nP4e7Qtg6Fwfk8I1uOEVyWcf2KKUXaA2ADis3T2hlzqWT7Zf5cnFELjzuWk
AkUrR3FWdCgiT6UGoX20Kz6X7dc+xRbITJelktrL2X1m5IvYw+Jp2k1pZzZaAmMh
q5Q1Ggo0yKTLhvsLmeTkJu2my7Qcmt2WtjmZjyOTtaHUk6Ze4u52x+sBXQ6OfAkU
3Mj4t/fjbpyYGvRc/WkfTVphawcjTsqnlRX/ReO4CjRkwKY/PlBXv/FgmRu1Pb/i
vrVN8QFWWjfqmTbLaoB56gN0sM7mhuNAXCvqxrBeQELPcgbH8uDgBYUJSivqwQYs
Yyy8x9AN9wdHP3rTVha43O1J8MQjz1rcBwfW6qm4EEvCVdHJ3KnnugKx1CgCgDEo
9pSZMXuMzUZ0yki8Wo8IEujCIXJcx8MkgYAsGm8JcLxg6mRyKqHb9m7TeOj59dU+
Vy4MNtGFcYNSaq6O3/+UFmQV6Vy6IKKaS5k3UPoTdcWAzcxPAUbfmaqO2XgcsjjC
x3oD2VohxhwEuT5JoHxp+/TmCSO0pyCggKzU0RGPfQFzWwsK4eDsAeYZBen9Mrpo
3gNFSYqXexOnT9qIAChH4NbqJUad41OwbkzPaq20rSb0O2EVwq06DAlrKYVHtdlt
c6iFajGN0XwUkRb7/WwIXc1zNqy4yyj/5pGHNPdOj7MBUdLAa89rBeGM56lwsQGj
fnH+hRySK7JJ7sQdr5zNB820lAVndi5ScdKJnwRq4fjHtiYrbpQh4lNSRPPHH/YS
E65RZB+EE8l81ssoVOECZhzae/f2bA+jnqJINBBRSc1vznUI8H0DbFlR5i1uuLid
S5O5M7MNKazzy9EnAUCNr3IQtNjCCYtlS5oVVKcHfPquCLVztwDSlWVHkILZ6DjU
+goTPv5KQSA69VilxXwVzfD+pZcCb2R4HnKeJJQugsW+/ecco1n/OE9eIjsrKE3V
OS08MSFWxlKCnX53x/oYPLCOxBRgAptIJtU5faGI72DkpvE6+zttPCtqOQbVGTUf
4UWxML0Ap3Yy1bYYOlcm0lA8q49HY0f1WWA0gn4VEnfnJjS0CoEwzjyyuOwIQ8WC
m6+gKc0SQ31wp8piHTN7bPfW8rdk5q2GdawA/ny4P5bHm8i28dutyqyFQ2SYFHI7
y+GAafdnD2S6jnH0hfvAkE6iNvuJ8Z3i3r9eLSxl5jacnotyM/Ie+koWrFBZSqVa
1IOpVNITi+BsmNIjVqhc9hzAxzEG1tjIRvFo5M92PlmhETDzj/MekDj62AnB6TrQ
rzUEw+drT/O9mMtTQGCKg3l4aMsyPiFxgbS3E7CLKGajy7J1uXggqi/9jU8eBQe3
MUeMepB/QzqQk4EjHpXpovupnmnnRe7Mq/K0eTqw4kStT7w6tPH5vYaPDo6n9XEN
40tffJaxNnWSpR5ayohhOHWW4U9ULgdqWapXRh1ppfvz8GuF4Tb5dieFxAS6CdVG
ockxg/uMB1ArUjQTx6T9B2dHpW6P+W3J/a5ncfuR/rqJUkj6IA4VH2/zilzyGOxN
a1PIbBVPP08awDYthwCc7NyCG+ye9uYtAiOvjjR3RuvjLedCQpnUUrZl4XZUe6La
KH2PdvXa6797A0/JTTnp8zg2nZFjZA5PspUMD//RtL3JrGXV1yAw3xIaNlqLNlW1
InlkO858RYEAnhQINpSSEMmsocBwXYnN2kHg/4oh54vG1UC2cCMe8zRBQ7uF5/Yt
RFkXuSWncCRclYI0wl41eXV6VbZMZouSCRoUjT9ZjgbZaHsbmawaLr4ErbQTNIlq
69sfPjITLdoZ8AL6Xg4Fot8yAf9O0v6oKQvBHazI9POfmIThFEKWC4BT+Zh7K+gA
2uKsxEzib9I5b9kmoSVyaUsGt+cHUr57uT17PSW/UL6M7M1ufWLXyW79Ma0aknFk
pkV/LWuH/7Nssi3qGftVAg6HwgpdpJ0xd21/nSv0tzGYG/9YU9/oJjXi9qQwggK2
WtwFfr6zJDA1IffYpR/Kn0qGs3Q0E5/VyYMFt7RMeV6hHgK+aF/PZVtWmVmhfim5
DUbBOzllDKaUTrotKwI13ty30jMrbqn1bgSuaOruew4nfRaYZcL3MkvmeRTnSXEE
FTE8DNU8hpbOsv1C7fcFz7HWQ6U+ekSYAAe3T9XPLJlESbVD0GoQJLXmbO+t10hv
u0FyQ/eNwfO6FJg2yLwCUj11afoBwTtuj8Z+mdZ9PTHO9hVfj8p3tR/oPmA/qtcC
vD3ALfKPFG/p+8f9mtvFEmA1aTCuxig+QzGvsjpvfC8HrTCV6W8WoZJzs2n2fyOS
TXIrhYPFcVHtQIZHQ0cSodm4togXQk8F1MwD1t8BfxVrOxW8XTj7jBxF6ORTD/62
nj8DevWRQpoSEk1OOp1Bdiy48dmesrKy8DYMIb0Imc5/X4qt5vSe6U+/tccU/VtY
zx/yea2W3BnDETtZZrt0SOUJ7M9Nm/nuN0KNggXksQQ0zOOcDl1YGPcuC3271Ghz
sD7JCYCzm09HxAqQi6H36b1YziAVQdVXazLUYvZf6dFWl+9cqqvEHcfTEeHTvixl
FnBtPSnfMJyWbgHdFikETremeYM+L1XDSJRoqTxqWEyr/RiukuQSB73/tLq5pRGz
tIphhGji3m/tGvfI0JVVUoNHODinVVuuW1Jlf6EZp2y6iyK/rSFA/qXllcw0pn6U
hnqS0RNR3UM8/g9+ouAZ/34iOLBlbgnoFwekKwxdREZA8mTcIo2e5+VWtfohv2k5
x8q/f0n/GjF18+yXbLPWqEY1pplNdmAQxTQmeFDvGcK2GZbh/ofceVfTADhEvKWu
kRJh3ngn0n5OZ6a0zHExvJLRaWfaBYFtY33MwP6gWbVRPLkgpv5NVhnk7sISV9Hz
Uojaf5D/IviuoqPDV8+unNKF0F6yh0yVb4KaaefIj6HQm+7cAGQj38MzTWICZJn9
iV/nuZlkZTPRGlyrsQNcWAPTwqnIeeVd6seeh4bRaYE4v/yq3vF4s/Qamf4yUW3q
m2KP7SSOVd2+YDnRwEX8pqbs7s7IEbfB0qLks/skSC9oS2nuoLbsdNP3ijtBSZaN
In68N9K/wyUolfZkmetpAKUA0WQf5Hw0FDSLraZGsAM/aDQ/G5nB2sPRDTzrbT8y
v6KgunN/VE3TZ3UrOAAIfPzo6xFCo46Tv0iHQw3uyrb14qVES5UMyj+6sDRtVMCD
APyJaVr+CFBsi+QhQw4o8M3Jtge7L1lFUtpkJk2Z5v9XZZxnkMCo6Ld6T9xP2/jh
7mSZLZFsOy2WOG5RcdsM00tsXZmh6ugy/uAbfzA75IFEzCOapr0EIZoG//LKyZcy
DwZlKOqH3J46mIoV1zzqVDgB+wfpTOMwr81/7/8pI8+upAYRBeSC6wzek2Xngyi7
z/dqKsh4K9BnM327ZwK795X05Nyvi4ltOf6HW2pM6w4pzMC9fnJRmc7lZPYpHAtf
KO5HIeLk1cL9SUKGTcmtYL9MrtPYBKtf2+dhN+LRnrFtJ0K/dAxWef+lUicyJm0Z
gf9Tyzz2/EYSSB3t0DS30p5MM+aLbB/MujvNyXBLNiEb3Lbtikv/RFCSmobe8gr1
x261XAMH3uTkFkMnJ6H/ogSO1prjt40F7ibt5keb9UCCjlKYwACiHGqwRCzoxg5k
bJkFh7LFWsI9t0Gu/dPEPqf1BHXC7ETLcBEkE5D++a8wR2dXdvL9oDd08iMCICc4
GJ3H05we7VemX6DKnTeFU365KSW/saKlQIbFMf1vIAR/Q7MDvLk15cSDbdb255QJ
iajqOn502OiI1hqrHjXiropHNftnH2BwUqiVIMLsUGmb4Zp6taYMHApsE6NxBr4C
iC5SoMrfA0NMWjfFI4PgYnmqy8OpUI5gS/Fd954LemsdkAa/SIb6TMwlaoiQ1ef2
XnP+wl7+H66a2HX5QIbZc7LmgQUEOSY2GDG3CMXsm17S6AMjsTawAn16FvhS67lA
tAXxmToxUldWXshj00xJIYu4khHZaLSNwvoAFsWXE/dxrmo8lRRPrUuc/YNUvp6I
sHzGlMF76A71cd69vj2C7g5p+uoigTFxkMIgk06m5TBXQ3BbMeCZmip5Ni1f3fOP
x8R4dS5maKDFc7U5UJFetcfVsOccP2/8uoJpuqemHFbC1+3QftiGyCaaOSapX1Mz
SEzekiB8apeSqIv9MY/r5UuzPlBjj30oDls2Ed+eXylNxLPPW8IewmgcaArNAv1o
FDnPZVDQ22ctu64rgw7rpWx5WFbLHAUV9ip/4HDgzvbYxOHnAu5gfk69dxtXYBxZ
RYDUkr+jwPG6EZWQmKYOhloRgLCAE6wznbCpOgACGNca6Ij3EhrcDWbCRxMWUXdS
GoCFB24VnqSXmofcMRglqzuUnp1dHLNgUP9mOP0hJA5exBiyPTlNP3sN7xKTXYeN
cLWRw4OjJvA9wzraeo2CffvOrYL31PnQBrE6YObOs8Y57lInY1eOgv1w0Q30ys8l
TuXHKWyODAJo1yAKXUSDH3mwpd0KRVXL2dGQxWpf/8pz2CmD5S9R1aXTX0f2ZHVu
x/8nZ+gYd6ng3u/yy90ne7jSWEqQv8Z64YGjOb60AuiLA9hIAy9wTkdG+SL1uckd
1/cJTZDnW5WTsCh4pP5R28wtIoAeTchgsQUWmfZOR4nF/7IsWJ9J/iQfdCjqIBwk
0U0VAyhHdP5JUe9G78C4vUK9hx4EuivAE2uNi0e8p27SYzUBmoTzw4hnOrwEvRPl
DBDEYajzp8YZtM6XG8NcNCvJ0vLObVMKvvqRr6rJtLkCbPgWTjXBQQqmOrHDpuRr
9434uWtvSIjQ7Q6AqnasK/5IQsxU6b51eUriOngmOurDfTmWa5GzcI1w7yD9muSA
X+w9VNQUZGhpSzemIrUSbVd5+ZOebX8J5XFxaGiimU0a9Lut42U2/4RMUbBDMaII
Fs7UC7kzj1M14+UXX90zeioQ6tv3RXX9RZjogvpVwgLlq6o1rEWy8Hx+kNN9wCJC
XjKNnCjs8nu/mpH+iJcgIQs6iGyrSOLb/UvKAPkOow/smkSnu12uaPz39ZSvK4c+
G1aXOJtz9fZs+vFYL4gB/iLQQeVRoPwwsloWUh3fvI0PoqQeHc0c0SNLR5gcbkBP
EhiQ9d3j5SBR7lKu4MaSAH+EobDmREizy0tvrh+ulyoDRqEnvtmbxySWAA376EdY
RendyYLKA6VXY7VA49afhL7PTKPq5Fbf3kdx0FQExgDd5Qa9EFk7gDMbgsYHetux
85Y8zM3dBreCTEKx2WGYZz0sl15VG+oE5xzyyIk36EzSlnYBkGYkiqFh28zqOe6E
kKM36zx1ngcGwJtfDjjyyjsdyG0oebHzxtGUPnfgKy3YHZsrUTC1NEB69fVaJKJL
pp7AvUlisxL0gLjGMjAHfN0C8rvvZq0V/Fpn62fjtZGvB2UBdE7k7Kw2tsSyZ1Ov
ShVE/bRpuT+YOXkemGzp/hbxvknJeFfkTbjoj/aA3AgLBHbZIGZVJz+EaEzuRnVX
fDWgjjow+d1AnLQ4TaZM2ZWxDNVqjN3YPzissOExcLXmrNXv5ZlstUpsYYaelSHv
wF1bmH1E8XhYiN2hoGJf6MZtyyteaQJh8tlo6rKWHVqOuJUQroKXyoBsj5MlK2Mv
HjIc4LrLhswjYBq8TqigfKiYwNoudSeLMZ8+ZGSMIpWEC+Ic6niNnTy7ZZ2ka7b/
T5fdHi1Yh1CB+5U2becbkaMAdNxrCZKqqYHXaTjC4P2XoIpewcjhaFgYfEAqUw6g
K8ZXXLLrPRXKVvou5V36sXSg+/rlbb+URynexTq4p6GGtVNSdJPXm1gghhlxOC4W
75nep0MmpdJ47S6wJMzUmmyBiaQSTJQwbLv8twz3IW3n/NS34nN5vL7MP9KhbaC5
taxnB7KeeAj5Yht2kbq8OMSuhoph7T7n/DQLW5P93OCSG9hvN+xxTzir4Y6FsQz5
npbHqVprQaoJghTXYy1vfWQc6VBMHCJqPyYvMrXaICE06rVmlXntDLdujuSR8oQy
GvX2WyZMvuKb2NNe9QhzGFQbKvm/cVazk7hXo6njhZbkn4Tkcib1Kkp/oZHswY/k
IDToGUnF4nb3Z+k5qPu8yAnSn0PMeAfpMeU/TsG6yCagixZjgYPJWjPUav1IccpB
oRpypMajd3XEweAdIlQLcI+VSAFMGjJv86hjae3mAIiQkxm34rmPZEUkMPx85FyO
HSt30Q7FMOLwuWzPrB2APGc68t6iEaWMHZrnPU0BKqm4GykUxC1z0D3Hxdtf6O13
9W7mIAShBEzjEXAfwilgKRo3YXMQJMM0BfcNH6sI/atRO8VXbWH6DdKbr3UzdPqr
Bj2o0S635RbDn8k2KGIDCRas8TOq38TP70YfR0QFpHzYKyu3/x3LtyFYeACPcPHN
SulwnLHDPnX34GKelZZpn8w8Os4sbcOde6Lj9PjmmeN9T8IWmdnGmptBvercgWRc
e0lCqu+zAH27k2t0tXkOODQgQfJALa7iuBJBcufHLEnX/NOgjYE7d/0WrFIzGvrA
5jLOyOAaCoqESN8T/BLZhZ6XDHo6Fl7ABElCt5fss/Ti+5BmVWJ+8xzGTnsaGW/J
YJ497F/sJG9BvVAe4UXUFqoBTZKAXPuWikwKg+nmU3Y+4O8hFodh+vVz41aR7SQv
lgxlcSYnOnKDj20bcPy0z1dpuwlxecJz+W377VDRch3iJYhG40h5aGZaP7Qz4Slf
dfwt1cD+A2vv7nMAN79j4+DkZaD43g4XPin/kCNRPVV3xp6Z7CLLn/kyBpgO23yZ
dNBKRhTClW26qkB6ccTnew24g8gRzASW/ctmwGOqIoC1KoPHGAzUfmPjQ4RSuOXr
hxAeLZp72LNgiK++RjJvxQGbAac1jJ1oze1mu8Trei1YHVd4tv/o/9pg9GXLFVRU
c8hmZTf08aFkGK88DBnBRDAPyBKvR/PYF81vpvTs6BqiC3uCoVOMdVTg8TmIqged
TNKo8L4Vl8HS5SmzywNnnEV6pEAMndeQA/j/GtWpnNjL6Ld7R8aokAXeYfTJQhLz
+Hsp0x3QAXeQ2sXHd6AEubrbNxCn0yfcyDD5NkJarYb8xCYJV1kV70/cDgWKWJYs
aHUobfdMMTy1MImiolRjNXXyS1y7UFavPFJU6sALiFX1NBQRddfNQYPBgniR2WL2
HcXlD5ppmMok64FWZdPsCa+EEXxiS4kuRkp0oCZM2rf83NJyK2tDbTL+Wzu7dXrn
YsUefOhRioNLQd+c2CaCk4AdDQTrdweq5UV1GS++BeBB65LE2EUE1Wd0wpIzaOfV
HXDZM9/Xm0IIsTg+prIn5c3cKUoVrp7vULIFhQ22mOxP+YBZ1eng2vBrPwY0hH9A
XzScv9c24+ZxrVU1jhxd9Z8djyF3Ze6oq+JL7BflcyvI1/yflFjcoO+zrEpUqD89
V+hgvyMn6Zw30lpt/5q/xva33hb4XzRLp1NYU7aX4PmpyO1R2HscAVjfC7DOb5XU
/CIvTtfpixWmYu7VCO8dQ6U8mHX//K5HsVLZcTYOU6WMT+GjkAFOssg5NW0vs/E2
nYt9vv2Y2/51h9nTOsOApwbzyTQ2XVSm4ABvYXLKflgPZM4y7Y91BTGIP5f1wJHd
TM6k8pAeuW6ZbHiyyY9xEib4w1zqf2Rxz4uII/Me3j+VbQj+5dvpxdQWa8tYF+Ma
sh12YrSPJqINk6wHW25OHVxrtNi77825e9YA/DtHqOP3rJjLWyV7ETOEuLB+1Uvc
NArsvUiAucAri/6YOTL3EAs/BAkD1iVgusvRYXuXD1oQw/2H06M+9kPxJg1kKq4P
IM+VvLZJ5P720pgyYwcTHcndDyQi+uqWpu0LoIO+TO5uWUqt2g8sGQfnQGHNQBe/
krHmlWL38F7DEgnv8G8Rt9IRn+aiOwjyvsygIoYacAm2PfaAlk+pHXMTPd9/a7Iv
RBmNAX3SMp56hZwhXSszhqch+AhG3QA54egzDTiovTR5SWck8uTqsz+K1Vy3wT3w
EIcL5TsibvpXyJ5mS6jOkkgCXd7KUyqmmrPrie2g2zswJzxkPtQv7VlcdSAJ7Ush
nNhxKcVOWLLkrKMATSVvygXd0+9r2ymMZaX7CM8Qt4XmKidJ1j3HVgyJHy8sgOwj
SnCL4nYvskzf1YRPqbbcCzEevk8eLDu+blwNr6SXQha5dVcJpAH97lRk2fIzvpRl
cvlg35gb7GWzdjioiXZl7mVG9jK8KtC1vpvHJsk0zbaT3iiU6vmIjjPuCzmBR8on
BuO21+WMC8jI91k4ZC7iBzmw8O23R7fFK7usZfmFBQ4ENiog5RXcDCSRVhUsVndx
52AU9Vd6euZaEIDiPV+Uqs86OvyHPijZbHSFqlUx9WyIwX7nL1sFwS1Ozx3hVvsl
0n3RUIkDvrtmEs2btqYtmW06xXr7KeCoeX57Yl/s0obLep5fWLGtpfbgW89yDTjH
YrcGVW2JkigxAs4/xGVCo9DOTK9G1Wb1iPrGpesDlAUfx2H4Usgig2VtS90SIiK3
1XVeZ0qLJepf0CyhnriknbaqefLPwKoQOmd/fVtoN+1WCQTT7/Sh8oS5siC7Zzzo
Pwd3nDJOIRnBYbMX6K/ULv4d3AdThzj4GT0vWotT0mp2YbTgPCmqLD3Dgly6AWeT
gPKvxITTwSUr+PrST1FZKgJ6kcaNYva0R98qGl5In4T7owJ5lnrW5m1ZkPBqUSuy
BJQjm0nOqRjvmD8q6JZkncVHJCrEr4st05Wg/4QHMAHrMiU5oKsw/hfNdogpn+ve
/2ua4LJfXZCJF78G6JZ2X2iOroUKVbR5c+kVzYMsQhwf5+A8S20k+orbb3saTD8F
vjnb5Jqogqd4Y7cThY6a8o1MUZpSM9K7gMEdXe0HE5e/6Al+YL3c22dT08cEgiAG
7zY7zupnVz7GF1MhKK762U1yA6+9ztzQR37mk8mwKfJtIWnCf22F8HOBCtDVfRv9
rGLUDrkwHarnpKtjQ7Ck+1PVHDOGCsLqXaAOP+iBKr2ovrjbfGZrEBtgx1RLhcrG
ZqeX1OY+mwb9jZ7wQmFI3/Km1Ry5mwcr3BLZ8ou4gVWZjy1WcuSYEEQutOaa5Bsh
vAAby4mvE/zkq+mWT8TRpECw1/cbMK9GKTBKRfyCYgw9whiiHuJN6Zefd72Q7sCV
OCL8hVgl8swVQv6VAFVbRSZQhRD/bjz8M//egzcyQ8UKMcAUqFO3/TDJwTzO6KIj
2BVr6CCN5+BtgONstWYLA2n8MW2MM5tTnnPMEDkX5QHNqNuFeTALEYEQCxWY1RXv
6zWr5L0s0UbrDsw92xQuhSUENqGorr2aFG1RKiTVHAzyhrl7dJ0zUWNMVBh6QKga
POREFqqsY3uEprCxyR4gKgkMyDI8W8CuGSwM0fPHy3MG0OgmTrGpqhnuHO9rjP4Y
dcMsKcq3F/SKMPR3BIlzQBkR7oT30K2mvv+PHGCEp6UXwSgB+Rz7hnY6EE+yJwLH
1tKlJxPo1w2uqihkDXWtNMaEPhUTxCPEBwBhGIzA5N7L3s3AUiDQ+R6OBLKFv2MC
GuUYQJdrcyoAj9Na2iGCAMGZeIgq+1HfUnsU9JGdGvZ3W3CtCuOeJFoIrSPy1TPh
l9BtylqgiYpWT7Cgl+jsiSjRdUDP6RXEKj8d1D7MB3ENnKldOLwuFyZeju2tkiCX
ClKvh5IJoytJBWI5eyDd+s8td754otNS3Aqy2ajcpFtLIhnjheY6LNmNqYA0LQwB
jOXxsac0Iz3vkoU6jh1QI5pyhwXFFPZipw1RupTE2YrIojmhTahtaZrnUR4x3dUL
AUS1r6mlLMNWzfsylHsVZcpd6EJ1vPr2gqPXS7BsWsKH1lg2po0KI6BkJPU257jF
RIbfg1nUL6UJFb8r6VuERaFg5WcuHbohwZ1pEROWt6udN1aU7lu2DocJH4VAIuGS
DPP36qMav2MKhunuwxK+SbrtbSNmvMqrhwCG+3/v5z6olX3t0pp8wBx0yTvufQ7U
dqBU+p+GykUoFgdFxxk1ZKUSbdbrSeb9e94FdHmJk3A3TGuzHwwmlppSuP3etA9u
ZlIwYPMvLErjq+oTVbueEtggYieEgkV5ddfXXUMXquPu7+8B0PdDCByuztALUk/6
ZFEIcE/YxvKr8kgMUSRtTzMgIsAN4LBsjmK5NaLQekxZ2SkLOzvM5D+ZDlsz99tp
aSnWES6ndK33w8rYMxV0LkQbCmnjZpF2jWiiPcSb369UVD70r1upWPDqnpnaEmvS
8PNMMDegRlnmn9Hd4RSwWyr/oMYU24X9UItX44ibcC0qzvpDigwyacLH+aPm/XjD
rkPxioCh+TIQSDEN2b271qIsJgLKgDwcfXRksGjLBf9b+5x8ru2hnNNRubZxW1If
FmtPbkcd1fmNyTly6m+6/fracCTryiv9wtt0jcefFcbHWyseVhCJqAmX90EZEAh8
WfM9InwrZEw6wKbYYbFRW1LDQ5Po4UvA8OxAwF17ZTWsi2oPj+cgbuuxnuBFccxJ
8tzh73oPx2h1Zd9UnFU43EsP8ll3HN3OJXUFo+0kmWj0RAa36YfQW6dOF31VagyP
o0OjMa2MKGKuod60EV0mUmnyTzaeTllnzYvFPTp+hfc0haMKaVjQxtHdr3mYmg/M
3A52zw8tIpVfypMp+DmCN66Ez8lCganp0MvbX0t30I5pcW23+A60dIVKHEs6XIsu
FhEYDLyNlAMgH8LqebUIIhaZUwWGuRBi9MmRrzUx8n4Jmp3a1fAtT6ilkef80qvZ
ss0dYo5/j6qxGnkAr68nCwpEw5z3IEm6E6RjXETR9aKgz7XJwmVuGN2jYCOkpny3
aHmE5tCkdNuPtHYxsr0I4A/eKbEuh6bJjroaAIWHtZW0nL7Onvr6zEz0vEaBAapi
5H1uvghRgsBQs+9+YhYJJUlyV0PtFQil6BRu+0VRjmcZ/v7+jLJfur1qJVSBwDmD
yw3k7DlgxZ40IKrW5SfuFv9ebR5F4iFJEThtrj6+t2bp0ZMfOzNFMydSMuQvVFwu
Rq2KrGVGLPmOhZz5PnWpc7gnnb9SGk8VMqkmMXp8gLop1h418Ddufi//YSAyYGKk
Z0W0KjWIG7NCFpT+ksQFW+KR62/L/xEZE6tQJ5rY+sFthKgj5GQ2IbX4B/eySAXU
/KM3e5/OfCgcpmpdd2+uNDtnp7/kuSm+M1Snp9HuvF3EiyBFdWY1y7A/c9lwwVHY
gph90RWiEjnk5OxxZz7GMia5SAA4c6mqtAL4SAnLBVUHcXZrEpT+euet5gRnBp+D
lHnLP37SgcbCVbQ5FPbBFLp6AOkcnpMp5BytSac21MmF6DetUojArn/VOKr7MqZo
HTktpMc0DZIAIYwy7hNBxgD8qxUs3cJRV+9LUmKXwz8dLit1N1gJF3tvJNybvOna
LTvoGzkx3mqndrvYk/u4jonMUDQ7mtRzw3BvVWVHv+2mYZSuFJKUEMhzUvxT8kCj
Vc5q5J1NEnU0nPpvOTbN6i6O6PntXaVo0ex6ZZiwS5p8gkFQKgWQEjBGI42plebY
PH5gB3HN1dOhCnpR5F42RSGqh0qudZE4bpENwDrOOOvWF5SIGZ4OQOncI6G9m3HO
SwZEigrwFxKtLTKvFEuwWmM9Bi1Iwfm+xUG+qNDWgIBbgtqq7ktWu5/Z4ujXVFqO
Ku10bBTVRIExVul9xLAweuWMO6o0HmPIMRp3KO34ths0a9cPJoJFw5b2KwCSBTW1
PnarBPFSqyoqTcNzYUEyzdtTXyyAagotkUeObciXPWgL0wTUYaRHW6PnWiGZdtRN
lbr+fKhXXRQpfyeaOFUt++TVGyRLcyImq+gQjYRe62T6sETJ0cjrM/Q/9OaWEvcR
psEIDPTYHk4C6ehmcvuLI0ZerCZJg6PotdBHk5pWhon3b1jcUPIUfB6JGYFDPJVf
3fjwXyP8qPycntCE1fK4R533tLjGtZ1QwBDVwxEb1HXGy3Xm5hFp0jUQC349gh6d
pGFUdgjx8bLBrGNLHiZiYKn93PAHxLFT0yVzYUMUTkRSNfFPq4aTp84TQ0AyBTeG
Xu9Pty662L9/ipGM7NKHF5dHECWTnVe6ZrkK9BLfoiSpp1xucA2vdOPSGSv0LxYL
0Wh2TRb9Rk4Zbd9g9xe82Yhs5Sl8cd0q1w8Lw0CpQhFOp9KLgn7j3yHEXJprLsnX
DRI4FRDlfIEFd3m4ipqDM6uW4GeJz9Ea8iD3AUxC262RXdZ/OoqNZJjw5OazOlU7
/T6WIVxaW5NdjenVRXZg71lnECL91Wzlazg/I5XmUG3ggVfLU3JbzRuUvyrlhDUc
b9tcomvQobPcqivoV9N/olALuvTk9QChdiDhOGH/eECDJs+g6bDfiJL8yEF/ZFNW
Rd4U4OqyipZW8YBanIOLF7W2Uo95LwOKa7uX7SiF+8WcrbgXZwZNbiogZAyjfQGf
wRvHoj5GInO1vevp3rQjrbjhwVFxv0U2WEU/qJgz6rJIWoHyTSYZphdJRqKNfJwT
4veexdQKtc1lfjFuZKCSVH4Fh1YiS6za0kB9jgSawkhKSo04IePFM/W0hbffKpkd
U108r1xegxsVHorSuYj98TwUCEQduVIs0JZwE2Geu/H23BICZTne/PzulCL+E1R0
tbHp+5i3DyMAqzThujiEV4NyHFxe58L8JhDFwWMxuKMzrT1pyESB1GNYjWDpLStY
d8mjgdWiPNLDCJPp05gG+EuC/wOAsLlApIghJbwYOzilkMs6ZiNJ82/85fzOyvpp
aeBZmu3uFuRjax7+wGnBsHzWQy/t1u9FIV3P8ZDyUy1Vz4HY6vM6LyoSBa+KTDQk
gbxpWybqOc2Hn/zI2UjXKKSsmyN0gxUoJYZWhpU5xheWPKsLrOoBVYLRkVNZMbCb
hihnuDt5qKWkcuileAb4T4jLeSocw1zUNDkkjDpfXbJ4tZhpiJlUAVPNUg4T7PfY
rqPtx/4Ovswt6VmnMZ1Xh3DFMFYBTegP3Vioz7eHRR5M2VTdjApw9gXR5D5Hys/V
zA0SmIjzIuYtlNeTYWxOgVuMosrmvGU18Ke+JfE49riyAjzg5twtAwCMPE8cYf5k
FPLvvD+8zeF03klwOHKSkRmxicMqSXkUep0UeLnVEhKc5BjVEJmgqszq7PNGRAqz
qp5QbRLw7oC4rsWHtha3ceSx/Ul+QEjh17xpJEGuHYl76ltOeN3xzZmNZ9gxoaRr
99CFegUX4VnQ/cHd0aVtT0oLmeZO5oVwE5wXACa8iT7R5SETCfdXrxuA/Hl/NK7R
yqD4KlDy7arhj3WC1C0GITNilbpw34aBBT9m5qjBmLEe7DsxS/PXYIHdSwy5vUeR
wJCgwAvWDC5R2s4R3MV645JqEoHzwZBlXKr3a+Q6/WpKa06NKLYZNnlmyA3kO2jp
W+1cOGlvEtHFGQ5mhhdkB2TufN5MfWF2fRZf+YuOgPoH7twdx4c+616gjnNeISBs
ptMgwcuv0zzmBBEs4sL+VYbmogS6gi72gL7GNb6rFEB0z9WaWro71hVvMxqnkkI5
TCAMh9rGGrPvBb+gEABx9vYkSGlkbxUX0oPowpCKhMCFriSOXFyHGPXZY7KpQloX
xoYchbO77zog+9q8AovNMXNi30hNlTRA0bsWGU1pfMLgfoer98ZHHAe0xbMRXVvO
RA8t1B5vukIUF/HU9uF6ww1AZNyP/PF3Osb4ka6TEmhMPkmAzHYOhOkK1NuQnObi
ADaVdegeSkmjdoHSbMrGJlSUEgAEnvlHDooDK3XtjUK3Ub+hmG+7Jo5Pt2UDnhjQ
fIxx2v+EpJ5qRgJTHBZHpargvPWnNkQFeM/b7R83Kx2XEYrdGJp7Fn54XsRMKZv/
6zaOyGmSEDljhYH74QrcqvUO0tDWmmzME1G2T3haXtMiWb/Ct1BiGXJONg6yxnZo
+vYMf+XxqVk0Fs+UDcLINnSIRvg/iYalLmEw69yF//hHDG+IQAdzETAvSgFKaXyZ
i8Wzs6Hked0jUFdnW2iJj/NpE+C6SkuI1exOAlKmyXsZrb7Zh/vJA4P65aS8IG7L
ghfN9cScha9+jkpGFqd5fMEKcV15R6BO3aLVw/uZmO1sHpWpmuek5sCbSXdQsIZo
GnUPizg+mJFfmd0gROlREcSArm0qxjKELMi6z4lmJb6x+UGso2sYyhvOQMvOZ61W
8uMDsXLtGLWQ7ZqMvifU0eDjRndSbdnNHJrkKqgdEUo6VtKSkdSwoiUD0tyx4acy
34cDh5yxelESUyYxhiqENXupD2bTY4m1wpmdXIcx3d57x7LJ/CwBFUQavfDSAfC+
RqYdeGL6/yvhdyYGlMiEQaaUymyoSrWsk1rJexw2bRCaksxkqZ2Tgx+UU91Lc6ME
gYwS/hbeCrSqt1GMpY98nNpxvbt8ie03V91slCsndqNvSRo33k8GP7qitAUc2rjF
IfmgoAwB9j3POhUI9QYt5rrm9L17P51M+KZ/G9Zkb2CATCscdoR3BFH4HRKRVKOr
iV0+RW/3LomxOKU40HTEKKpZtA8PFfw7h7KGksX4qqgvCqiHxZkeHspClqNeaE2L
UqdWiunXc+lGZ1eqwfKe0I+gkKReSCWnGOBJO2P87NH3nCtBzZipxFeFygKb+BX0
go8Ix1I2CjsiVM60steE7cyW9o0LPhrnX4GUkbYJASn86IwqLa9kroAr9SmUuUsA
j6ttnj0YbNGaINa+Bdd1SPUFooKfJfFpPoittN3RFWd1gRIQJwMnOCipqZIo7hWZ
TqGI2qJbWrPy0DXiW3fYsUbVBS00bm/DPT7VPAJmfQsnKcOEiWTk6zviQyP9/I9i
ijlHBoGuOwcTzufQ2AeCeJWFjgU0DYHLBVJbRRu27SPZ88sFup9OY+CdAHaiDWyb
kPJSalpxodyVQeXelJZccL3vSpirHbTWBhNTBh+xfLN80oYq1eWyrNbpsd8wrlkm
MzEu2e1KB6gnBAdUaDTfo4+FnTj3bk9s3Y5uCSKpmZaHESF0K5340mQ78MqlL2lg
x3REPsGkcxfdiMRe5m12lrzp68sOWsecdX9nH62U2ZoWw5W+H1Gej/YP7o36Imx2
ZizeIf1mHneRkN5wR+sUkiQbToRyV5ikgpStDJWlgw2hwBzulqMljagQFwblfjCk
9X3CdPUa0c4v/1oQeoAHhpNMfhff1AJiVAsZB78ME6UWsE5uXoOA8gyb2TuV2+rG
`protect end_protected