`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3328 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
FPPR7ws3fN+RQyk1V5tkgFbkxRGWqYEWfhT461hqKlyY2GcW0/VFFrEOwKWwcSNc
Be+NyYt/XxARXJoa8rAxrcOZljsnRXuExaL4s+v4Qzlv4DkiI/18CIDcS6OGr+7w
GWywo2PujbYY6braR3+eTyApnIBiqonF7Qpzd0MqxlgJ6SV2PHikHUWxZQDTbHKh
F0H9d+E+4NQwjbd2RHuB2kDFTBZ/Y2ywQWFO8oi5n0X8r2QEW0DURNvwa+q8PFFB
zO2T6iXHYJK2SHZWzLCTef/by2M/jx3Wp8Rln4whIwA79/Qqtv2O6FXh7/m415VD
cvwThu/sWT9vm/oPvOwiXoqbOMtzyQCeiRp3lpK/SxdQJD+0HXrGKCzdKVAsxT0Z
JnaIIBrN2iN6kDGTjyd40C193mCQNRrbX2G7zXUL9Y/yCSpbIJbAKjRiviMyEDRd
CuUdmBNv6Z0qbKAI4tTqQdDugbugK2bKyWYX8rycpCW061imqCKmIIKZteSG95JO
c8ItTeskR7QO8P0bA0lkmc/RhRgd2/IxbRhN8I4bwtOLAvCcDvVbCYd9PoUXB9VP
fh4UXZx+sYAp3HsJU3lFPqq/DtgOJDleRU08yP0t+tpkB01E5zW9mGv9qkeAeojk
tt6vXLY2n5U40xEeIGqBZjUaW2cF6vhwM5VVAsNe5jQd/zd/V5pfvt+9/nshMrrP
MC4Jv/xCVY2pgDFO7n15gs0E0Pi/JmQILshSYB8RraNpEEqSn1XEO7RmHsnesNKb
mfbizIO7wxADmiAADs4yaFn1ObsegweFjUItQxdotL2dPoIZ3yMFbqLm/RG/x0eA
wzTFKuA5pI1GOfAcRzxsZZWcVK2+lqEr+RgL8nuA4jdnS6F8mgKQcRCYRG6tO43C
BL305Et6eiYLiP5bkxzqYKK7DsuG50tP+SyvkdKfLKxmEEpyyUWJC9KrPulwcssm
iNGIBfA2i33DdTM3F2pI//dQyb9xqnOWi+tIlZy7VETwZgDsQ4HqUtEOSY4kvI+q
fJmGISzz/oQVcC7IkPHhlyaoASK+uTLYu73K3CDh+YeKtiT9goPaOZ1Kxa+KTSe3
V6fjAAL97Or4/Bd7UuI1V4X+yIuoB58DT7maFxM3uqrFgfnuLL079LWnrsKXmvwa
btvzzKTb1HBSxFIIgvt/BbryLuV/vllApS7uMOHh92cQG8Y8Pj3pEa701uyZ6F5f
k17fBDtlLcUzoB57D7RJ/B48gA4Nxh++tagz5tdtn2qMz3Icg8rvMflCL4kH0YaH
D8LYJcedUjrG0QmrrfrYIFf3RNRasrjtTGklXg9cgXHSZkrzpNuO8lQKKsBUwAhu
aQGI5PyLIOwUe1t1qZchdCTANhLgSasoASPt5KNKJpTYseZzhAMNA8AnIeRduz95
gQGbji5yocksCe5b33Zu2KC2Qi23yEDTLrKDMLB3NgPczNMfqzJQ6A+PTNWZb9sA
nqzsmcBeJxk6/7nP5gP8LZ9SconwlNmbQUEUEIu0hQ8CRssuMjTiYUh52kaFJh3Y
HIIBmO8k9tOpX3G4AuHbMMymVI9LPh2tJSL9p2PAHUQUHzQlm1gGEkeaXfxge9OX
vHnWls9fQntzZUbaIUlqqXF8CAQZ5e0/tWUaM8Pzhu6mipmQi38dDteg7AKWzM35
ow5oGayaD0TQSA3zjtjb7mJDOOaQGftFehxfIGDvev8WkE5D3n2uMWbbuujrOt/O
UHVjEGshPjes7r5rLwC9I8COSTU6SsFkIkF/3ylpUHA/eWd6LOLsx/QsfmqK4vog
VE7kT6G/oGKtSac17mIyqqqD9T2wTBmqhz2ivY3zVrfGkWmTkMR6Kv+ZeZp2KzBT
WjcUncokYx8wsBpk3fcwfvoWn9CT7TudCoUckxKOFsUPc6WW8ylQM/SWbUxbbAPc
OnJEtGYLkO8P7jh36Yze662s0upDrABSCwTg0F2MwjKc/2SwHvA6ZyPcavtThC91
4txSIB51JmxqLeB4szIqTX+jllZkuKYvRUfyGGta3Em1g71gJkM0huv53hiI7Ahe
bOOOiAIWgPutGGHp0hCN5KWR6jsALguCRkptp6yAXiktZlK5rnXtti6OGUZnoCrc
S/62+5hrj3J6tTgigyUwqtBNdV4B6ns3S8AmvskgKcsj/2q3rfsZweFTCbPC4ABW
RntbWgYYj+aGD4DmJ+e0aeRrFy0t7477YjYvn/z8dctUOkhuzYVtwlTnMURH6Yck
mwEilQhWqMUkemzxigzVX3eR6uE+7qjp1zG7b5EynokAHYGDQhHX3Jhh8QdYfeZq
LvB93M3SISpdhxQZG/IW8HRDIe+j/DiN4QyNfDhEuXtjqeQneqbIhaGplDrmJiU+
/v62F9tzByl0pPBnQ6yeVNi7NH2o01J8exV6nFG+7/OJFQCouKjW+BZyKGIEHNyu
CDXRx9zMj+jjBPd1Uhjm3TDggBV1/l7YGQGeQXIip7+wHShJqqNmKgir0GpBDnPV
rl4iIyuhBBpq/lJGWAdHoK6vlDSaZTVDvYSWh8pVCKqrbp3UNT1rgb71fBT0j8DU
BN+h43ER1QAvV+lBE6t93tuBDLrRKxHSKbo4dqsqHbdOhKKxnT2zNx/Gb7VNnY5w
gcrN6+14He+f0aFxaYVQoSDax77m428TOnl0WAcWkJdYl69V/7A3PIc0rmbpRKxd
OUNTuQHx9UkKXXPeCiwwQKdXH4+Emr3T/oWKlIYn9XJGn+YcVsQsv78CJaSqRKZv
9fa8VbsUxllPEWYGiPy34ATNAzn+jgUvKrOdGTPaxFxT0j/SAyIhWUVyGIkgj04U
yIYnVYmxUiCXzMkzBI5ujFD19Z61gMy+3jsQSNUKoPeuhvHByuxC3VszxiYpoR+0
qR+x3VABwVxgzDhdV1yzu70J4MFzMRkLAPuAPUtMcjG+FNj9vOMcrjRcL4ongJNB
ALWIsDxrJHTjCusrbfJRfvwJddLoamqPv6EIcRfJUCVUnjUkMq4vJ+5cNY/gQZg2
AlGO8fWqfSCDoU/IoqMbDmWbYjO21AlpVHJiZGcLtG/dmu6kLCyYU5saqRaiplVw
44NuamhY5jzXLslZdVIdunEtL+z9fws2bcGAZ779/gF4jYD1vxQz6kXsBjhMG+FA
UJtL/sgw2+lGBTVISvo7Sgr0iXJSkB2bUJvWLJEBxRmsanVvTUfV+TP1MHhgceHx
iwr+XznboXxZc1kM90DZikP/N4vxeWUdADn+PEd0z6zP8EzakzXUyMuBWKbWICHE
XgTZKqHeMNvH+NYwi2IzhWyvVNbrI7eSGA+QCi40j9omOskq1/eM8b8FQmbUZwhi
tYnYKCbvWDNpIE4w2azmgPwLk7dVJ6vwqCCH0jONRYFYZuKn1a9dxHDkapMf/qta
yRc1hkx1jBLiQE2tS8iR6lLJo8MYqaU+n3JXC/C89d0iEDH5u9AHnLj79CAw+mIt
F8sLfI3hcuaFYDEu/uXrJeaYHVS7qRYAPNTkU9CED542jEcP0rK2U5AhXZeZjUiR
AVPW2MFqfSrOLZcLX1nFJaGQZUal/p+L06BPa73w0Wp3XUSSxqrHUt7wg74TM+5v
QsNf6Td3191Mk4RXVIzk4g4pgVoQRbCgrvDiwoQvoYfTs8NryUabvFApVJZzzWE8
I2DVMbAv18UohMQfA78sEjoD7lQ0ytmmzqRwtSV/h3EBwuuf6r2SWnpZ36NbTlz0
UqnSqESPyWNUNQtWQlyCE/Nr9HdUprG55J4NWWaZNN4q1+VvEXLEta/+vSBbITKp
MRHkJwcpQlyRUEwGmDyqTFdJ2KaF/IeugYO94U1D4Ts2ZQTejxltXg/NqFnSC7lC
xgnUYeLf6foFvHji0BwhBaUz+GYgf4x4qEZb3hWlrULn7moIU0x1OGDCEI4IE3wa
hg5X7pA9rlQ2M8+xZNpMSg6Ut9yYRv4E4FR0dkPqTbrCMgvVxMW3rvRXltaHdRm0
GW4UDtKw4g0k2+wy05x5GKHfTg2f0/+/+8puuOiSC3VZuSa+mIK4JS1LFewlhc+J
hXyfLtnA892ZeegHkAGVK+UltOulIDVSbaQAO3D1SxmJofA/v/F8LcV0FjGSoiSa
lCLuSfXjjy6SsI/IRzRCQKxUcY7/6iN3puH9moHIn+l0WU3k5dIVT67xLR4lL21v
AeQ7S2jz7UEioYYnZ6Sux6Ml4SCRXZiR3xAZ9R7pjOcFss6HGE83EO3VkqwQ+OgH
9mVQ7m8h3pELgImFEC9ikQl/7AdyIyV58+SEsXlGKj4LnEdP37vBcPAja7NLm2Fw
VKx2rgGCOtz/D1941MyiGw==
`protect end_protected