`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8224 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0gQgIG1mJzulW1XOK5NnZR8
C8XqDUtXW7uOWTnSVqbIblwOHrDC/GFb3kYl7b/cVSRAu+acR+DcVvHNDrJf2vmP
c4Xg6etCN8ItIbctZ8+7byTptpJqCgrSN3iR/dcAU42OcBiv3n6vj1nsM9p/+9KV
FIbguLHvt9V+vPe7X+JY3JBlvLX+3Gs+S28lLf3QW8DZjX47HJSN3aULNGdHfhPb
TicV+xCncONb+oQxipDGQXvpDc0CWRxcN4GzhTL8gsa0cg/DE2tkJ0Zph54lBmHL
GhmgDVjgVYYPTNXkgbDwiA2dh41QPumWSwvJX1m9+xCDCjpccIUGSAEf83LlkLms
GW/y+PILlvr1gOeBl1++1KmQgRxGmO37EjHb8qKTtEqwP+lfolcvA7wz6eSeIBzb
wni10b1dFAYrrGFHjdRUmxKsHBoK6nIVkRpk7jtdaw10K/ur0Kxz/AgIu51oLk99
bG7fPzXYqFzXbgWHBehFqmtknb5sQfnPma04HwCMvpBAZCq+7CKxpHmvlvPNEuAb
7EW/pV+/6S3cT/jFnDeX4nCJxW4J9Cx2ppIddqNDY5BUK9knsGuxZmQP5bzlLaqV
tiqbVwCsA3RAvVKaQ8TiqYIBSlavy8ZGIsSAMfrBF3C0zlqmV2PWKrclvKnaNsau
Mnal4KtZcHFoOgO7tAJ4ZvbSechuBapUNjKWb6mMpEOaZLqJaxkvvyIxyKpyvSO1
yUigs/aK5AtYMA1ed397seSO07kTWE6n3JglJi9QtFuqdjESiuqzgG//9Zi9KSe9
hQb2x2Xp2/WwkZOESC96tKM7duLGIHMNCRRjsl8WAk4j/YV4FpaLBQdqJ53mLM27
YWF9ys6M1+frUeYIGmZAYOQCitClR7zNXq5lMNE5MF0GDlpxJ3UXN1Tu+yWo1FXk
kia5hIBwEBYPbbxRA5dLwuhHn2y6T1/aTtBIGYTW6cQA0oEynuRa3lzkU17yzY+g
hcnbQMxn2wXTlYnAnzyxg7rh1V0Ay8qcxIFt0sr310OrRVjFEoHo60Mgyul1aDtY
+hvqIaAV1KX9IiwktW3uBs+7T2LqGK+hh1+Ql46X1cInue6nlKhHY8ncVu5DNpoB
bWBzOwJ2w1hW30A62pJhnbxak1sLH/UD9QJb6jH1E7hk301Gx/UXxllIjP02Bbua
EtNqGdszVtCQoqtqq4w5MeL1lOTLpCTWI1piBEAzFjwFoGuMidrAHK6UPIFYsTiT
sbp7RT8XW5WI2oAKgoqE/WdL2LXWf+B/ZeEoVPA7UVCi4ohWYJg6EgK+fz4D31Bx
aCf9sBNG8yQXqoAoAl+pEIqu+fJIUdo8mTSBYX4s4OzFcFNlRU7Ir5I9LwWm4+la
DfT0lw6WyvWhBP7yP80kUrOn6vCL3Ylb0zp+ZKpOQM7Mk+0lgkawgYZLNpE48Lc3
DsNyoOgZaxEy7kpmHPke08n0CgCJFsp5MCH6sRh094WD0920k87kemhfz4tFuOMS
jDLH7Ue6e5m8FdRv0Mtbb6UrVPbYuTxH1/LN6GRT8bZ1qlWCCv8avfX0f4/KRAy4
3tz0G/zjM0UkemccMYv5+ydlD8oYakAzc0M81g6L8qxUdHBeffcfPjALohCqI5rz
OdMAZHUdaL5m6kWnVVWqXjRYQRZ75pt0wZ2frd+1Wmf4xQ0HloNPMeVQEoHuvWWo
Tpcbe221f0od3JU71eRMrVOu9ais3r+zKOw0lw0PyzfTvlv1XFxZl0CWk4ey63r2
ZLZWFqtkx1wjTFJrzCCyUBjuTc/jz8yrByatPvvG8x9c9nimt+/jZDgfAeEsGAK5
NsvpjAJCtTkqfFCyWprXYLful6vpARScAc6jRzLnNV0Q4CtugTzsxQu7QcX8bDCh
b9WnnixKeD51+0hNBsj1r4iJjxitR/J39Qzhzxq6UbDALeFH+f6zC/BihqfN11pJ
otqJsteMZSPPqybXlkLqGyFHpceK5LtAr4vftUje1lgL0O+FUBd4NKA3e6lBOOcC
zZh4/n0HL2RcqmTg8MiZftbM7ilnLsBr/luULysMMpeYGYnTOdBB9SgfC/voVqFZ
YYbT2Y1PjhWe4zGT+dzlow55GQl3eC6xWSdbQ8hOZSoapNP8DLK8Ge3eRMSL9m/o
EP3MdQjtBraEQJBDznLqMBm/myEMmWBHDG8QAG9J8o1evVSQ6hVr7Nwbq7fglv7j
VidzlvHlHSQicASW4Xx7XPnvBV3Y+ey/Q0QzCl2k34vMCoCGv3x1whEtCDwATx+w
UcGvD6yD5PtEhpPRWvA02y/8fdYm5LVAEJ4ZiYLjcik1yG9KGJoBooZZpMe4p6DM
oX9wFMhboMoO+3N3Ai1x8oaosTln3UJ9hnS+RdNnttRJTduXaB0+wrVBkItqtnF0
4snkib8kR8OYwR9tj9aXiwvoGIigagfFAwfo6FN47xeE0wn5pY7hin9BtWyp10b5
ODcCH1D9AZ+bOiv4A5Muy7dUusJt2M8BftR07bJ1GEIgs993LKWHoFc4JrvdkaOl
/bZu9/Lfv+82IuIfbuE3dbkCQhYAJlgyj0WOUW5wIgUOWr5rz0rdf6VNxv3YiuJ7
lD6Ci/hXPMqT/o+wtY0QP2o9TUImW0F7gw7BK9Ub4dUuVjVB3BA9k5KZx27zcG/7
Eb8qHdkVohe31uqtIAkz5Lq9wlKYNsKVBJgvKE9EILrE4j6tqX7dp74X2alXscXb
46O+UtPfYRhe8vvh1ZVnt3qsKo1qW9iuTCSWFcemwUu+2LJ/UzNkbrFPuAxynPR+
dMKeFemoF+ioKPLzTQMCPTxSb9GKzde/COlLrWncu0Veid3r1zlKB6vvQOKStvK4
9d4w8dOLF8BY5wfzsJKciauVT3Ywo/kCuf4cgGfSA3MmJaVVLVL9iCYrPQ5gyvKj
6DsPIRCPyxzORIhVWwdEoFYbhTMnnNFQHGyIt7e1pg4H7gQCkwrQNvTQAGvsDg/O
28PnxU7NuwFc7fJspF2pd1ZKGaUKT8XFhc2EcEfBkda0teKR/2Zb97/HJ55kp2SA
FqiaURP9xqHbxpkltA8k/wyZs2XEsJVoZ32Khqt9cGGlWMAUKbqY6oJWdMr148IN
6EtjyyLsXJ49g5QYRh+KtWdNSAwOiGdJC3t1YWHYwWvixLCF+4mlPTUWV8X+FTGr
fMyDL95RLy2zD9390UcByBzwD9AdFSk5oJB8WJ7vRZ1+bX7N/C2//elOsC6yVH7w
7ccPzg6bVoSsLyq4LQ8dLtEOxdBDIGt2pUCoODwXqXEhso8hsmWE505i/8eTlVd0
k0WAwOHIHLnCCQVnx0tKCl1TzDW3390kqBihCM+0Rs/BYTQF5DBLc9+NyvqX195D
iw68QNvE9Q0sFpxX8O76Wbx6TSxgssEcZZRKiRbQQTd5+RKBpEkF/YaJxNTKHhUX
ok45MtE239Vkov+ZqWGhJ5Kfijcx6tflAI4/27txndTCcQkJcKlNenevEhFivZBR
cQZ1Wj+3Ux8gdzdCvbQ0yTnBgSu/z+OuVQhrYoy1pu+w8nG8QHYjB+5SA2baR68l
csn3A7X/Gj/DzRgsMtt+35NT9IgO5AlE8Vv9PZH1ysF7ijAlZHCJHCRWzszIoJbK
FBN7QpA36zieYCj0oY0DZhurOerpMxRlpLPt9rGA57KFuXXjMv6hfX0JTqjSGtY8
bd2YL+7QFbhnBUN0mwYzgM+0e7rZeB//9p+ROpQES8VUUE7lfIenzbJSdbTKyrcv
sN/INYDONPN8+41AyDMsy7S+7KlT5vnT69xmGMQHQkXBMt+xM1RzX5YUBlp04bEc
UaKQQoZb64EidYrtWaGgukLQmQTa1Av8cSQ5LnGukxe4L0f6yweTIsm0VollNWgz
/3akOXg+D7AV6BQUO/zMWMJr1icYQtzPhc/cLL6CW9gwCULXyMMk01W/fNRxXbOR
swfu+nDlvGgrFkRlfFiiwZgxDNxQeikrLB3JLkadYD+dx/ew1Eu+8bFWjVuuIAsa
LGoip/AInF/ZC0TxDkClqH0vifxXYNMYin8DpjBUp+ethNzWjjhVNDKoUYQpG7W4
dGmPpSmEriNsr6MBVTTmVwP/zJH4APLUSxc92IbL6OC9Tg7xG8msN62tCgdhMD9w
ceYpfJL7pzRWzcAACFCYE62DOFP23eLveTvZzAAcu2tP5Wm3jMscMgKiC/dAa/mr
CfSwz+e264XStLaJSRtHTEEsajGHw2MrLJ9zVIPChDlya2dJnA1NzdIAIvQAQB6D
6LS3U1hZ9ZFDGf5Mr855XHYKy6ts7yinlsy5ALpl4o3TKkVsuVw9j5l5ccgbrSYF
Iv+5h319AXrDLad9nH3/ndEXCOWfmYKzyXVZim7pmm0vSNTz3T1dALWYLceaHTlW
qCvZZTxIqtZR9mBw5f7GQ/QkONvsIophFY6Yvz5H2bOr1HNkUhr+8fGS6tUcO5YR
VX2iVYa9MRub+x+u/prrqrxyB4gPZMpWAYnstUyomlBJVwYeds0oEdrAHtwLlhv5
9/7LsvjUCCr3HKfkMSUKh52YgbsGRx0/cK31BvoIQzmDPDE4RaGuvRvDoQpAUnmK
aiyMRl7Amy6A1Rcu1y/Pg0UBS3Wd40Q8/xefYWMyuZaKV9huehipnSuvaLS6Volv
33C+SP51rgh5sMi1/0eXyT4ShRK7v8tMrklAinOTYQk/2rv5TWPjtYbyHLG3uo/J
3FfXUcyGmHBKVKynfcYvBTJ/mvORX9uxucXAyX3Uy1UAZlKeGEN+JQ1pI/NLoEnB
rm16p3ow+mrq0DPlmM5ISM9jGfecwZX7KXtL9oKzoMUHE+lenuXzk2mR2MTLmq5R
msNHxWBQCeuN0/JgNAZWvH46bwqRY5VsoPjwck2AfVt9OVt2ZHGJq8ozKD7GYE8D
3H24BkT8c5QDcgLIOvXzBZNKNbA+JENUHx+GI1OQuTdVusimAecvbcBmN2YxfLg/
6IK4ABo0XD12RB2dyFLvAFo8Ky+ey8Zt3E6uyFUyVJfSGSsuM2Ou19KqygsU+Rrp
W6Sy1KEs+gN5Ir2owqAEgHw3coNXv+XlQxfn6WY+iTh7UZjxQgWiSpm8PA4P5g7C
NGjRZHb188DAF50pF/L7vx98xO0rmhC8wzjLVK5Z0BVDHTfymvvOUiWsRe4OTEQ9
CuLK9d7pRfHGB/a6Q7HjNTomfP3hoMPMcRcRRoEWLu8cuXzmuJhZjxBF+IkyNVf+
9ngVmpRB9lKywgXfgFTKqkE64FG8eaRATgdXZI6DWKrqavMx9Unxl9Z3SJ4THqRb
pqTykeQXNrbyDrpNLzeIKSLrM53BpTkNNjDqBniOyQUZGJSBS6cGUfldftSdauSe
uvPpPiNNpg14NlqHpFqEPX6Ai/2hSgKRjZ6Q7c+R/UbPd3uZsj2hby7Ja07rrPu4
b3LqwRVTZz4sKa9rSsXAPeqTMDdj9O8joaW9gX50pp/tKyMgPppb+f7wgV+A17d2
okFFTfoaYMjl/0NGAM38qJgbMj1YCNsaAEjoDrZNf7Xmc78cn2Zj2ww8UKFIxaAI
cPHQCNwxJE0hV2doRgIPj+2pQk2G9sb9G06W/FcO5Wm/K190RfDZt3ZpSDRXdGQ+
s/dNfPFU0WbBlloqSIyWd4jVdarBUs9+puhM060FxSHJ0MGn7UGy5me7BOKzqrGN
QcnYMhQREu+yTBWJZVMDV0CnHF0Lpmf270HkBzRZyAmFh5AEM4JbPgZuk2E/BaGi
kI9R4t6xBCBhgOSIef+DRpx27FmnGDJcoP63qTEg2uxC4cPuCEheKtdnPZK4jdH3
JYGXH3IsqKnaNQtnGuavM1Wosd8ZqcJYta/UIqNXsHAYJ5WMMQD+sUupNTICPKVh
PJv2Uh596NQj7/xdBzZQ7M341zUH4Pw8OIXTpUSRCyY20uNVRvcPpWXG4gJ47/uq
Q/ZcYxwrxOPbXTwMMiP1H3VeFu6yurR3PAMQ7+e6aEgScWn3AqnHXWdKLftMJXIu
MqzPwHuCf3PXfvzTPxCZJlAhgiLbsxBSFn0t29ESIk65RE6DgawnbN69HXZ2o04C
8aR8GKLRee7CBkZqaEPYGA3O+7nY+nCohjcGbldXVfNSj8xmVabMLNs/WxuoCVJc
khYmI6Vb3I8mnvOoigj8BCle5OuFiAFQ4NjowwEATGewxcOcwfDKrpMeIlwJ/T8m
FFdPiv9wD3hhW3nCeuGr8yYnz3qpreZDzOHoo7NqpM42gXelQXEEDxNX56ym9Wub
dOU+SwxP6kCUzxAX/aunMd+cLX4R6QfItwHrqeKLcqD+uDbh7dV6pClLW2lxbxei
RQBqnvd7XqsODVGMhwT+WTpIdla4nz1w8KKr9X2MPuxk7s111OU8JKMIePmILUFW
kOm/o/zqalRiuOecFo6DF/fITnPhvRY/MecvPhfDSqtil12XL6F96UnaSr6NfOlz
nC6XDYvRTWCuM2akYjcR0js4XgrXCZduFqiVD+Qss6Op9dl9LkNsYmT7oGiQA03q
2UAgXbpS+FaHGLU4vdLtNxyI6RHr13Ivh5/3O+x3XNAjtZW2Uz2wSE4q0g9Y/l7F
JXQF0ADjuX8fyXX1M4Pna97VkLY+7bQR94K2pORSwIpvZMaJkBgYaI9Qqiz3suK2
JEE7bwPN4mwtOjczydwPKsttJZSH702hVZFZibIC/z6Kh/EVdN15RWKQ80qatDso
lESd9QwcASenwRf2jFm4JFOprLdp4h/niVu5jbhT+T5K7ubJN4O28cFa7x4nJkUA
pY4b7sicAQGB0eZtLuFmsmldoPl7IPAAhPxzxm0OsMIABI1B4m7GxSDyvtjaj/ly
5OfRzA70teL5eoffzDn1lbhj6jCFiP5qbVqgZj6rUwb9UcZNWUlS/jGHz9bn6/Ai
s+8FvnGgHX3RWAagqjOMmRpdMnRDtgxC+2DHb1sZuoIU/nSJEIoIPBxC2VtV5TS0
qgZHTlNMWNORS4fC4O64flUVYoGi0w0afla2Ngbz3nV5qPa1eWmdJvaOQngbs6hr
MFtT2EHkqZTXCjfIUjlpOI/qpCj6f7ZRwepwjXXCVek2baOI/uhZTaAgBuZV0NVN
Wis+J59pwpjcTdhCeOWhBWik6ux0p+eovu0kEcQNZbc2F37pzYzWNqbi/pxoyRUB
4oz3xkIOf5BS35aqemqst/Jtc1B2pQShxegQ/a3094kb9tj/baIU1YmJz+sRWRiM
swgb7j8YkKmPv42kplB4K2Cv696rmq5YKl7w07exlPvtnvrcMq6608v+e77o0U2k
iS8/nT0bUqZCHE7Hz+5pBhsff5zQVfOk9XYcgKJGggNwuY1uhEhFpchwieom7qzU
tvfTazrZWRwnamkEuifyPPkWtrD1dRAOPJHSAKSsUaGwTwimZMHKOcZ+OkWRXAwz
Kajbek8rDRjISFKJ+CLY2zGoWm01m7H3lUdk5Q1N1nLTd6Lemy3Sa6cDyMAbLQHt
H2WocJD+evYlhULMHEzEkzMv276Khu33k5but12nUHmerOhf8C3EudXh+cLQSfA4
+kwMdJhS6AxxJAjh2qQZgJPISiUHppPdhhrvS3mXiKV1mPR+ttQc/gnQ4ARijxOi
c9la4M01CO2zFtyBeHy8YeID1RJ6FdrJdOa3gu/M4FqsWRhh5zpTDJhhZuD3fQYK
Ee8/mngEGnecu6O/hRpjqYtMno3AX+dDcD8hNfpaTJtCGpzAomKhoDEOMYybgluT
L5LfFKWkUeen3jd//0v7pv+8VlNYog580mawKbvFOX/fsekZG7aEwAKBz76nuKVz
OcpJ4prHbw65t4qtlKfLicdMeMGqFZ+fcLbs2cBiCyTlVxx/M1g2HXrjGHst/ayT
QobhOtnMZAGIiMxNtPwvgW4zW8ZDc+Lem1bX1N22sU9PN9NXAzbyB1BQKb/H/eF4
JSKt7E5u66+ecYyiS1qG4ecStiV1NXn5SJBrBA7ECT78FYKCVxLlDxJZynwvr39R
z0W3zn70F70jbv7AErn9CmICFqATXl3DqMWVh4gMbdmojI1FkuBusYKfWEpL+BF2
WXEWIAXx8vOrgCTAFTL5LHWFIBeD8n+xX4eUiCLsq4UFAYLG8mirSOUpRc6yCFre
d1Aa4VbLeAgen2HoJWCJ7+vczCkNXyoC4rfbL0LFzgxIL/dPf4AgUyPrv+1L8wFQ
1HPuSBFPhwGbn17C+KR8ZR9qyfPqUgMLf7lI46hZLFruRiUXg+Iqk/N1pRa5Ttrd
T7XHAXeSKGdSlfheYOL2RRxwG+VXrclfyWJk/PftrzDZ6scGHWIU19baKUtWL2GK
6Pxf4o/vuJD4o9bQKn8/rOF2h5A+L8NdisgaSZvpTEI1nFq1NBhSh9Wye4zh3K87
IU1PiL2SB0KWwarfZctDRoeCRtOQa+j4FYJHJ1K08sCFnKxN3gNG1fciDm559du2
CJb5tSm7YT5P5Got6cPX5BdPWJCWdpZNKrxtI6Uj7rRoFVj3lBKAG6Mq9F2KastI
Tr5tmfujKHwuUyHjGvnL9IxNjZ6GVBkqlcy2dYKZ0P7IpbAoTxuGBSkxsPwxgqPb
Rf9wUPEHGbznScK1lI+nj441WeJYBFVjpL+7I3G1mqA99ViV7gl2Wmtwo/AVSDZg
j60PbMbO2kPUQPHUKBuRjlieGx1n277xFE4nXxliEgCH45HnT5lqStTJNKBiiiAe
Mpi+8Uq4gM1hDWiIiO9gtx0Fi9fcuQCoQgZCJsQyZJ+qnuHa7NEt1jEau8ryZ+Lk
ov50dXveZ42L53nXeAzLwR12MEL9qRFPuEGLiWRUvTNQZX4Y2zC0TytMjY1M42ZK
tNAgEAc9w6lcQaZLyPTCNyG7jCA+Bo5PkeT+ICAPnOz9ssZeIZRfeXqqhHbhxxas
5y6VEhoQif0aENzSlLv4gkp0dWqxuzew4+M9H/f/I3/sPnGr2/iSc3dQ7ueIltHv
n1GdvmI+/4U3GoVBVgNEO8tnm42qhtwwtfeoq1Erh/++jwMFI+dhh+F6SX5m+kOs
SvT7cru+DTmI0Iwd3JzIRigZEVhvViWnhmh0KY1wy+aVxSBYGMf0Rl+RQZHjUYqu
JcaXg7tE99z/GHNJ5lBEtlwljvSlyQajIrXugZcMdsQb5O7dnxUOfQz/GDn8OLFj
0gI6wlBlE1lEq2BJQQF2zm5pzxonAo9qmdpfCAvj8TBxyFg4MSBxnzLw5wWGucpH
HK1/PhCsn2T/2jaRiSCqGZT2JM9iAmnO+dp3i42YclhYJwZFSXw5C+4DyU3Qlbv8
JZaoGAIMvjYmGxpOxzqQtNWw8OB7hvBIJfxTZbRROH42pTi3ib6Nau3tNwktbVEe
NPe9hEyfeaQzqmgKq19O3FWuCHRtwOpdQjyFHslJgfVBz0o+LBQGBQfk1pe6zl8L
c7C8SzneVI7aMC3CVkXl4ie4+tXrTnUz18iDVRJDSwj5tm1nQNpJWx86anuFvmUO
2nBcygWPfZq5aSUI6hkow6EAClwv9mIlycjl7Df3pZuGksLnpoZZIjCJBtoXafNw
BbukSovMXul4oZN8PkleRYal3gUqwzuq2JEj5ARj1q++q/nrQ1Xw9/reD85Qr5+W
jPaj+C5IzKJ5KhNNUzbFQ3emCuwQyna7P2Zdchg4gebDhDZbRanCWL2u6HFJ0kf1
MI4WjOzwQJKDHhNsO26/q/eoIqv+74xFci8PsTjfIgLPeMzqGuqmPpGRHcLlDasq
8RNuVTbl/oStnatshrSgm5tCptmfKMw8OWrwPkwaKT8C7gALD9+cR00ON0indebO
XC92zq385xcqPTSXESsQH/MBYTk5FDJdvojR7HfKaQYSzAJAH8i2W8S+iqFt7hDy
YJb5pUBgd8EFWwA2VdRHG7O7/j7y+UVp8EfJE3aPbbq47rZYMFMREHB1MTj88EfA
4VGCohiIixw5mgFcwIyp44skb3Nd50lZHTW2YVAl0xMdsJqkz7DbQhfaE4vC9v9I
vJkeCHDa4Kba5Y3PpevycE1+Nm7LFBaRrSUIrw+fGW7FM8I5q002fGa6Un87kWsW
XG1WyKv9MJS7hOp3AQPPoHeOS2W49l2X/GLs4BcQF+w0Dr41bb4X12mOAvSbhzG6
xjOgrgttmHhIpibFKipaLVdPDoAWLZwqr7Z/UC5TzE3+Cyj6V0yqEORyVTqHShT9
JIO80HFCq79QgmsuNX5zzBX1IVfIbDd4zmvrnbOP8vUmOs0FCrSL9tqEX/negSpN
kM5SykK+WySoDasGCqQbraKyeQbUrHZZQOfDAtV37GyQYtsJmapWmlFfxAuclX6a
jRdX6Kc/gmQiRNM12WnxfqxqTKoFGUSh2NhnbKTsc0fFhglC1saP5tPiq+jGGHYI
HK1HAnTj9YVTQC6IEJCTC+egxuzehZftAWZ5x8O2fbU0xZNOCzrDyuJcegLyJQbW
0RmIKfqUk3ge4+Oz+vw9PduRKcyoV+sKl/GsUP1vTc3Hlf4HS8pEaKhJicCRLokB
ul6Nm0G2eP02oMpQz6ev7MLJlt1L2fsxqUPW0hbjveb4cGp1JsPfNr8S40X7Es7r
AslzxLWeGwZlxc3KXNF0VWlzmFVljaoBVCQg8B25z0eW9w/noOXwXx3H5AoxBHyq
VLsrK4MO+Bnrtim8jXDzseW8bID6o2iLwjNLLzg8g1skzbqS+Ga6leldhKi9JHPy
fdNy1VZqzYhSkeTKwlUR935DIe1zq418aw5KsP1DPAeF/fvu+78lsfSD3sMRrFPn
zXXWl/pu1BMEOY+wJ5ezVaGMN1MGQ7DnZ/LQpBSKb2dHQLAKL005PLjbiD/fYEd4
7lPVRfOe5zuI0DirQ3C82DxTnuNpWxbCr/QCrBMQ85ND1ubW5jjTWX6G9BLWyT8Z
X7LRO1RogiNYuCY+1ElH+A==
`protect end_protected