`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23616 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
lWGnzVBrTm10Z7M15YtSo6rKDpuAW6gYRIrmYyRQ9MgVfX6Jsf9s7dk9zIqylvhD
bVCEsVTKEfpwa1vaVpFLHA/2CGWEwM+iUO4Zz4TwavjN9daZrpmu4i/xpAVP06aq
vV4wODy97GRJpfL0QHOkEnJkmfvej5FPnIA3wq74LdmFF/NMANbOazlUHY8knoIn
slWmDZb4toEb3eUya3W6SLjOt9etlOiUfUOzh763jdWrOxahc6FMXJfXqophKXzT
W9z3Aj0E1CglPgscDS5aWDNAIFL/2hTui+7hjuSE1+5kUHMwY/xofXWzCXXh3fKw
jAvywtg52ARK6ZguwnoLEl4PJ5VgOY+wzI4PJHz7ih67wUkW+cgA3wKUwbeXCk7K
8+3sVCnfo8uLqVVw5SXnSAZRy5oqLm3wErsILrRMMRbMf1eDiGaYciEWeYyYDQzw
fWJUY7ivk10DDQQhMSisNU2Lxa/79ZlWtirzuERrFk36OjMMCiqXClOQEiooDhm0
QQKyPcMF5xg9haRLHAH/5an6hfYfMaM8D9BzMDZpuo6LlgWSPIolq8IrWiQiZMPl
njrT+m3SSlaABAZ8SKQx6NczywlPt8GHoMbUiw6oDoLizGx/85ia3kdMw/SALee/
mtv+QsDKRNrlCs55DUL4IaWIGuOnyw1QISVa6cbP9hJuUHuDTiYTJt8xo6aMRoe2
+CHn2IdPWGT4Svr5xFuG5oPGaomd/8pdCxVF+H63hGf9+Vzx9AJUnYr+rSMUooRD
CVFCUHl4cMUyfHJISOi5P/U/q2tYR0KGh3qo80o+PJ7rz/ZwRQb3HCkRzHy3FUOT
JiRS2CDRlilN2mdnvIqZy55hkirE09yvW5YXXnGOfw5xI16YmTh81W2awuRFPFlu
mNHSAhl/jGFIwKIHp4JkUdVCCJi3svZ1IILNCjMVFVZa+8I7CXo3ZrdEhHZZr84Z
9YlE1zpDyXOv0qXeZLXSi0EHr9bCFsEHpUl0sjM151DLxs96jdkBwdGt08jOkWDW
xDLFLiCJxbcjZJe72kcjFHHt+gVKCqYRWIqKhxHAgiwBNbr1HihcUjRgRjvYssBA
4gSWqcpVrKF/tYXm+AVjv1GBQHoT4e+X92JqUWWBf81+h/VyyLxwPxeR7ygVIOHD
dY+HhvZNwiU6zIfZ9R+BI2EztydRVsENasU86LGxcMJ6m7eZacsIBXtQ0dEIpjOa
eeGKPic1N1SPv5mC0iV32x12JeoFBeNustdUqD1hONA4Z4lHXupwK5fAAnc84zW/
3+6xDKdUNdd49oGSf7gcQA+vuz/rSjhl2Rgvos1GInWzTrt4dhXa7GU/6LLuh8ZJ
Hu+s5TlP7zpVaP2pfGEAV8qev05+OZvt4dW68IubAXMEb+AAoXTsVHQVccmD+Xxv
mQ6AF6q5+TO0jPSFwYaVNc/j/HeFXvAG6L0yR4RwtqxxZ/KX8eA7MwgHUuDVw34X
w/0XhcG07vnRCyoRNXBZZD1gu3AhY46IHVmlWRzvpTptS3tVWH+oCkT9h7XfTxgg
CPTS/7T7A9GywMcVPe3wgjKBI95YIEVwKPWVkHO+vqjVz0WEMsyF/avQO865wKh5
Pf8Svw7Pp6v5RWTRJ0xeBEu4yrL3dH5vt+h8XBVinpX8bEYYnEySP6FAkeeHjKJz
Z/cOvZ+VE+feQfDvCJBr9pb7tXRMNpArOwTi+feAn+0kF/fn40h5N41i/P+wG6XM
bFee1MPTcEiDwsrkLHXGsBxqfAmTiWU8ZYwmJ0pSQP0b3OENoAEnCdw+KSGXSbAG
62NpcZlf7xSOfCOlLzY2OccXYgDZmItx7rJu4GoTvogeo0mz/jd8YfbjclpDXV6n
KrmMC5v37OP+7BMeHnUAus7N9C4QhdpR6ErNaB4nWyPgPjhstydDyVT9DYV8EYZi
5mkYvP03IHMrLmdgjm0c3+WHXAlVj2Zcwx752rbxkU2kdL1y90ySaQz5iGESlS01
5aNwC8qSJO9rI/NYNjKGqKKAOcGtCmogMQGyWi6rdc9jhQZVhGUhs23t5xfbYA+e
dUxUoK+brxuBuy+vtZTIrfgU8ry1lhG8L5bEuNGaNAWYeztIeFoQ6RVAbDXa1DHZ
Z/1NwDxWZO30mz3JMYXiFk04HhZCVrXN196g1D7dGTKp7Kk8Ku86DhKrXO2qaIbP
hizl+247CEnbIIvKzN/X6u1xCX8dF1Pae+N8oJO8DB2GR+8s1lwJFrUYv4fzbVU7
vGS40rxrwp0rh8Ed5Tk4xi3LA+9ofNb5Q412PrcXIZMSNk16+j/7ubXB5T/NKQ0n
xxZ+Qc9OxJPPSBSRtkXSC5eBUDr01F4Z6M55gdlaIYLYEN0ML5uWfUCxTQ2igAzR
FWGLhPdTuef1zobtwaeNwukZfT2Xnn0MbeYsob3j+7pGi2xiHSdMKYQMaxOuzhlR
N3L+wose87hJg3ccyZEhx5QkK1EcDo1bswpa/DJKWTfaRriVs1aJLBEkBYl/z6rM
Zgsjry2gOFvPtJEeUiAEz2IW9PR8XyNUfPSNJwUp+TC0Lcklq5HLqfx8hqawp+OD
haZM4WWeeUBYU9wfnz6+dkPCb9TnN25xY7fDoQ3vYfF8OaSLiwpsDpdgbhHIhkQk
tGMGKrfXvLf1hqo8PWAxmSC36h51389Pjas3MJubBwZfkddVl7UltLWaUCAXznWB
Y4ag3F5LQ3tkZ3x9xSCJl68X4Ld16/+SBi1Hn3bS/K5X4BSOak7LntRCM0dHMF/5
6hz398yJZEkbKG+am24Rb8B79UX1+zrEMyOdbmy0EVubLqP0w/cZbEqmkkz6yPJk
vahzAC+D6p1E7lVbaHtfXmJhZ+oNYL+hZzin41NZEct5te/RawchJfH6qw0NSNK8
mbcCQse7qPOcmmC1A8pcRKaOHZhlx94A4lrw/S6ysVaDVel1Oag+3U6ASpjAALxV
TI6bfEdswK/wwPZ8rGuwfRlFOUiE+6Hg0pb7GUfKdOxne4M7AkTQEQtjOchZcxyn
2eOjB51JDiO13HjaKZGPeIAeHkffQSZ6DgALqRoUtnBEfG8yh/Z862WeEwb6OZh0
bdiD4s0Y+gWrvkre4+rERXoDIuEyVNQtDmW2Zsi64YNG5PYBP+gVQH6n7ePNISbh
EW6wkuy1BtdJ0GvWgQXKdFJsvPxKa4JteJnPp5l1O5VduD1OnNLKZ5s5IB4SVk3m
sRCHEbCoeOdKdR8fSkseRC236ygimNKVlIIikxHnA3W+AQGHok9cH6mOjUg7HsaX
OZN4BUsL87i1h3giFd02xNiaESVT8rRmt4qaHF8x3eesWY8cywP5k3TpGWiW8Ors
u15OxyxrSXbbY5JvzK/jBcydElxj+WG7jzywp8euqE3eEa/FzHfaWu2aGyDdQyI8
rIeLcz6Cp2G/uAWbXCVW+NfSTBy/UcdWlHJWnVTREKlsI6dxCh67eESvhWdqv8KW
4noIfByLiBIQ/gGxOuDFoMwrAuz+9wXWEhYqPNPwJ/VecFcmdF9AS+AIPgewxvXb
Dtg53DqKiw6ZXdicxCZAejZqKnunwmh2tUp4WxtDJvbTz8uwohUK42P7kAODp/hb
JEavLgimaO+UkSuA4LXkyU0oQ6Pfg4+pycAiiK4sCOY8osukEFKgdhw7kRcUIIuC
uN1nv9Yo3NIGlPy4yHS9aq3no+YuNJVmKxf30tf/4eTuqW1OqOXBJtx46gUbi+N/
5w3O1oL7+WH3ydZ0hCJipJ6pmrOuSlJnPjvyfTWlYEw0NE7PrYjWPQH84bBjShju
/O1RiFKAmLpF0qap/tn3GZ1ZveMjw35KoqZgEY8smXx9amPtf37V1VbKGaiIViIv
7HUpChjhGOvdwtk9+Q9IZBahIxsqvy4WnKsmPwvUc+5c02x74vcP9mTINjv8gRas
3h6MZ8/ef3oMo91c7oQ2wdUWCmEU76CHJnHU4iXWuLq7zKPnx4DxB9c7YMjfRWtw
WPuT6sr6nz80BoxOnRYeCUOoFClsd8E+J6Gy1eN2xCdSdJEBY/hRVS+1VtW8gwt2
gPG7zebZb6iEq1I5lnf6KiSz5D8tuYTHXE0FIKr1MoyCwVhrakL5/6vEmkZTG/wc
qHXH8LoHY4vWmU1nqgbYfaMjqxB3rL8y1qkjfDK1kVQFH//bU83lrltBaEV5X7vS
rO6eF/AgXuaU1NZE0Sy9GPJANgykWZWJOcLrdOJI21jNoLKgWcQLKh1PIDCHhnYp
ksuUNDIPYGKpR9Xf9ZU8CEP5SjpuXKkZ6VqDXBGPKtQg9riFUF3AhCXALUC1AulH
Z9DrZjwk+Z98/rwjk7cpzDm2682ziR0KHnMtPF7er3M3EMELXyzuUqHhjUaCd6EX
lnNf0TKGjklx0WxG+nE6F4/tAeQOreh/q60PLeWIc4cF8g/Qfzh1f7zwSuc30aMc
Sfhk7HVL1INW6h8NOegjLUrVXOFli95GHHzdPglu7Ar4+Ue6v8ROqcL8xISak04S
aTmALdmcQax84c0790EN9lLmpvSfDVomu3qDlCTELx6Cb0mZEo8l60wVjjMrgnh+
zj7TUoDBEBVAQEaO9A2J4+yIEyVP+k9aYZHkxoWZkrfYS9KfLbHBrk+lvG3l4Hef
1LtKQnf63Yxdwi+VLVfnQEFmDmiNYUct69MNiOa6yF+mkly/D11WtdDmHIKXvqc7
9JPJJQeCPSJzNApSChvIJ2uJPscndewVWLSTuWs2tjsUleekgX3WZJiaUHnOGZLE
kAupkvg+r0N5mTXQLnBBii2UEi9VKKy7Xm9ZAl+xHOtg108WugHEtR95IlTN07k6
um09Lj2hXqjOFx7HapJeiDrjBJHEBZazVCEcqdugDg6FHX9ltUfYumlhQSnZ8/ia
vU+DOcHnfoGN/H/u3/SpcsaQIszJQLgq4a7Ldne7zfjKGr/IKRfdHAkncV9/r0+/
vKwhdWn1c9WF4cJvXDcFmtbXDG4iEG+BoP+tNzB76A9cW4QD1WYMkhqBCL7IqXNb
aBqBT6SP6GP1DUe1QafccU0Mj8PlL0ZgU2ZCGX+JKonP+BEiVC1XRJgHMOY9TGfS
hz41Pgw9CY4PXsioGLDcuz6UYaqTgozMxcVHlpGyntJBDJdxxTMwwcBbgvsctQeq
3biyzQL9DJaXQfpAIdDFsNbjR+FuS6FHFwuiueN2I380EHTZehqOjbcMW7Zcqm8A
Crf8zMS+eTXDvr3Zca+BimuZVrFTr9FMreJiSpr/zVZY90wzMe89KC0SKj1/m2v7
P6+lCUeDtmEQrm5hHgp6lUHUdjcHYXdzdTPXWWhOAqkShe60priv3oYutlfnsAUu
KsZnC/LIBKgiZwR6bvqgnKHyHKzhFnKTyYP95NjdxlTkb8axCMWfJ9jS0UAJAaRB
JwuTAj5f9VcaGY4QwHVnOWRHg23FEkFuzijrOSz47q6d1TrgZ2fK26yaQxlWLYeF
hynd9YSt41orqICj1PDIkD8JO+Lw1h7nUciYg4vpJnRPMXQhrvw0QpbszQdOtWIQ
YFt/TWO3ySBx8Wr1oY6aPRA46Giv7iqw44fw7Tgb7jB5E3CMJjP9UAbN5sKhsKJD
2DoINq1VXbNcxHNgN5kUFRWjnOMnDrqW6/VGnvnptX+61BHj2useK2ECCfvkqL4x
OHsf/ZXZD9NaNbwWdrhsRtFfdejmUWqqKCydp/Tl7rxoYBmlkgwo54YEpMVOe0WT
HjilYmQMTG5GCRvbzcUpDYX1w+Ii7xrlp2B0K9xUgjoV9CV/3jkg5k1oi3Xvic3g
2vD9jKy5femI4hjO64qpG2N+hscR2t+Ffrg38uZgOFgs01m1HuXo7tsut6UlrftO
zlSsJfvGaYv3VjXI9AApUzoqHL6mmpQFiTf8jaSQI0vgDfA0Qla/45VKoqX/UlQr
LBo8Zc/tBaSzJmTd1Hamzd1QE6KjLwiKsoarfZP/DvvvxKAwwsXU8BaQQwpcNgDt
Rn8eaqWiLPx1IOjTckR2kaZE4AhWrjWWljf7h8JFkJDQwvZxPRQKcq0TwMPgrGy5
L2t0k5kHgb/qcHmgaz8iR0KPQpyoUoWnGKje4IwspE15kTfjCIcoM69T8BAjj3z+
Eo9gKk5LWSBcFDeP44ImNg28yXITwe4LM8wQd+CedpYSA6k7tB9pfmHujPt5EuQU
ttrQYujwic1zJYFXGsOGErqJZq9VpyMrzVCy3rTWhUwZmw/eygDhAKmlByg3afBJ
c9ojJ+1FjIy5MQbJOlV2Xqcj1/gX14bJa9zziTUCbOUoCKZ+HolU9/sgvbnaM0Jm
P6QDdzHZL64jAWnMhgRpNnh+7ndRmoG0dUn9b87Mpwed6liyyiima3+Cyp+iHmaq
n+w34UtGOCWAJnpJLb0/CwWttFMAqBa4J9ly2CM2E+KgIUfoai30ow8kGIGMSn9I
kRy8ScVnZNAnGdxL06wVTbOAp+m+cdXoneDmOQ68QPt2EEjw5Kjoqs/2rGIa5+fv
ectj7zvXSFFI/QHRtCoGsx86kpMx1ABRRNADNTnuJkwB1tsZ8ELk19REsFYoa13Q
mqPF0XSYOwMK00i15mZ1gjI6StYdXtqtso7+0NqufO4RjD29SPzvfT/tyWJzIZJ2
pWVSY0016Ogurtwp6kC1XP50GrOGMBSTfPQPfNuFSuMuheN6qhHGSER+b4HVqKyV
jsYKsjbPTK79dCPLojICOQZ6O3KVe5lXYMSUquiZP2IU9y750MYIEJAFYq2rsp2c
g4F5GRAbbZ0TPj3ssDlnLSGmDku66l//Wt58AYN9sHc5WbkTVxQ9IKKHCrw9ovJ0
nrbXSClaZ25wr5SbAitbrwDVNel2x7doYEahcxb6cMMWiHrqIljeU397ksiPi5Ma
zVpyhpth6YLZH62lAwnjW811Ry5c2v+At2AY1md5g8mFclhJTJuSx0HQ7sGLRx6U
+GTNPCM26ciPYzFo6MuR5RrSUUJOjSlYwKiTlVRdV+UvWjWgzeEtewMGuclq++9f
60qzog/M9wE9ZjTzeFYXIq3la9LmmjW40Y0jfn/VVl1XPpErfrkL6uDki2eC1Hay
1IwYu+kdaP2sWSsQm7A9k4q0wEMQPGM6zdAq7ILRhOS4YK2TPPnk93JY5MhUOcc3
9vYapoWN2mDgaXgWNMVTPl3udO4OU21yqwcmUwL8lkpK/RcI3brf5Bxv73gFHzLI
QIw7pH4UN5WG9JfwqJ/7oPLIvMsMpKP0+UCuC226TP5BRWdzOGnlJesYHhIhIw91
jU6dHB39BNj0P4v+9KlP8OYWAjcpSDFPl1V/5/O2kb1jCRiaJbcq7zT2R+mxzZBN
qMH8mBpuU55haDoBdnsagoe3P0xLxCT12YEnLL0cy11uKJBDiFuYqciLIQ+SGRPC
StqDOFZypwdyLh5rFRJEW56lUQhZ+sJErHaVYqEYE/+l5J3mmh6/VFn6c+0N9Rmw
qQ3ZUurOe9IHdySKv+/ReylMIym/cspBs017VUhKGcMV+qLG9qRhMzb53qJh90Qg
RcyRiCbF6GS0L25XHw/0qWLSWBBE6T+1/qhWFVTm1ZSAFEIv5HdX3BI80naepEmy
fAABXAgXjWr/NbViXNZS1VzPMEdiHd1MgMW6Qxdkf8CNCWcv6A+/BicVuN3sWI9o
0OPZnfzGB8wksTFJIeBXWgbAx8ZJMS0axib3fGT31FuNfXlyyP431CmpNmxEbapl
3ycpSg8XV7AeReWV/X588hOSCQone5IwFFjEyHd4kHEu9tJVwLe6vtaJ6Y4d7QWb
amYLQHLzJEVQETm6YrCotqGiaD5YuOZAIYrd767YmrttfSevtDTp+T6/Pd6GU+7B
22pZQL+A7XnG968dFGVT8tIuoybw4nKvRV4EaCjn6bLL+eCCtZhSVyWQ3itV0rTO
qvn6Z74QQt87I3Rm6X01JNxkEGffPF5tF+xtul8p1zP0/209TVoWM6MLU5ZSBl8r
zDelXKofek1L8QivzzPjVtebuDvf3gxZzvEmEm2cxoJn6wxHnNr5OgCU0GOHP8dz
zeOKUB7XILlbthTtBUy7B6qB5E+L1KZ/sb4ElXbl3QegLSUysqwFSO3KHrt9+ijD
1Wc3vKm9PuP9RKQNKT/6RfZapK0V4se0vC1jJeMWj+k4F7ZiLOiXluH3y6huDs8m
FnIq1+t+Oav5j3l3iBoxNzuM5euD2fUrGjdnBzju05t4SrQuU1CN8GfavMXoYceC
5V7M/15FE/QP0q6akYe2IwfpCFEV5x4qO88USswAQd5Ux8npbhCrC3A7uoITfGXi
f9Yb7/gyaUMa3KodN91ekOlPGrMHZXRMVFW5U2VqrTHHueEHC/DxNWYiR4UetaYZ
Ot13si83wDmgVnI0wkcBwoCS9hy/4yfKSZmceEYe9Do9WCvt7Wjx3y85Y+qfDMKu
dob22AOQmbI1tEuR6A6jGkOHaumuuH5Gu76gH63ybBGCOjHasXXactJiVgRxc0nt
QYsk/i4z6+YCna9+Z2PrUSZQzyzK4bx1e8pWrXteHtn578+JX6uHG83DypWUCaog
B7AwScSN4/3Tmf6gebk4CRMgtN6+ss7UySYqG9ofDpL8XCGfkkhwdwH5PQlSN8ix
00AyOYuHbamSh4db422wqERMo+NFGQKSy1dRWSSYzMn3zVnfjlLWJHdxnACTKVXO
J0tS+BHD+Oamk3KOHgnSeSiTWVl2gAOADVQtUYZB/Gc/qEOjJCV54WDHQLggKz77
yXQ3v0JFx3DfyaGZUTZ9aqAFK4a+3yHGDYlIGd/4WHMUOhVYo89JBucw4Ti/DDdq
JrpvybLup3RFMuRTrOmbPGgiLcTmdopZAFXyAoLQzmjeK4G7D2YBrN/sFyLwMMcT
sq871oY1Ec7aJUanmMEWYs72DoSxPDvBpbw0W7dDUwPgQTMSjUYXovqCTlpDWtAZ
Vts17slzqAzPu9za3goBrlR+czMCGW0iCV3jZr3O56giHPydPqw/Gt3729cqelyG
/XGdGCkDhhRy8vARJ/nXtivBWL2Sr2sl9bQSwOny8QTA5HfT+onBq//BIJof2w9b
gA870IkjnIQY83hnyg9zOmSDLpsgm76nDDeJXsDkuWn8IqoeTfy6xkTpFkIVIzFl
87sExCFo7WkNGyAKUrfbw2t3JYB5nVQPK9eSW+/iuBHO1YIzFo+8ux/d5kmiEJtE
a0YfEA/9iMGfNir3yWkkGJpCvjZIy3qRToo2eKSdPnIE1jUyH66g83GXHcSWvtp6
LlxLxvLDey1lbXw3f9KaMa4pjHQKnh+kxglycjj38DzAGoQHn6abS7oUpVZDhV5f
B6eyAv36RVa9Fy2wES2azv0uN6HryVSfE+IKLhfW5JUz1gNRci+LwTj+S71uEXoS
LmJ6S8Efhae/la3akmbRqQCmgiRdTJIp1wDe9oaOCXnpXH2ervUqU/jjaFOL7Kan
ZwGGJMcbioeYbfbMdp4K6MevPGPbW9hclW9FEMFsGyM9BjmI3/oG7nK1bSTTqwBA
xdn/j4C3nwT1BxhEcY5IRnoeTUcjIkBFtb6BBauBcWhA7KQbNRrErAYFx9RtN1Fi
6HGhAgMXij+g4jg34pe+UUCHGHmfIjuaL06L/dyIsNzu8SDytCfGsOc52jb9G1Ty
EBjyY8h64Cd8HITH+QEIidFsXiWm7P7Z1a2O61tCw9RHxvOAQk2QesZLDDyDy8jG
NUcTlBBYhrOG76O4eYk52B4KPVqqWtvBDWfTwvZ+Y6zd2lcMW8ic11VJu8kjICOl
UtnZLZS1E5mW65PcUycAWNvOihbygDQTjvpQy6xQMR0yX0c66GbnKjjL/OgY5tcn
Q9dcNJN9TwrVtD0if9Tf6DCKscx0Pzf3NYUq8pV2NGDUHCbVJtomX9l0yBcOi04x
vTfieCbQ4lH1MHPX4zSEtLX4XmmIlivi8KOX9r7xGNaVlzwovhbrqXMknRGXnfuW
17HeG9WwdNRgz3GtQDJYC6l3uxyamqEiJUWrOWWjPm9Pa3Yu9Tzl80nWi4En9UoB
Z95JencBKN4A4KD1/Dm1GPjkewp9wPwY/hEc1h+OrwGjjXDeZgS+RJJFFHu4KB90
jhdkC9br4I8FFK7rbV04P661xHhQRrteAgQLTxMzYd7GS7hpSp3OHg54FuMFzkDU
UcPeCrLn7LofA7xVWpMv++gq1qTjR+57wb7VQV6UDzoSEjGocqqqGQZo0s4pC1wi
DnaxYV3wM/NRDTNYF/Z4lCAZpwRtNiN8S0eRMm981Q2gouMkDYm5qbYJOLLe51/9
yCEX58PvjvI7FLyd1XtsRLrujVwLGQE2ff3AeVamIS3a08fxLqM6IUilrgbNoAKy
FqNpq+UcmA11nPpABNV/5IGWIcR6RNEh3if8aI3giS3F7LEWaErJprT8XuLImp0a
KKnV21VGjh0+8naHqmjVelBQRFvsCCbz2NJ0O9K1/GE3GUwbgXyJjfC0ras28Y1I
MNbqFMnQs/X3gLNt4Tckubv7+8K08m1PFHmVG/RmlZm+wBQnNncNhHXBMjRjqRjF
8YrnZGZJrb1PThaWojd2RhzYTi44YaPl7N3yzGic1AK1icC9guW3CeFkUGxS5hy2
IdbLzEZDLqptnde2AdXVLe1WpFoe1VXOr72XvbOINn8N5CAZifkKPabkxqbLj0k1
+r3l2/kuyQ0KjAWQ8sgcLwMnkPkfsx8zxBPkEdxI/HasUPDvLtvLeATXo8OwT37P
2wene6jQhzf3VG9yt3dwhH0Rg8l3+PgLdV1MA4r5ptq1M+GZz/KbyxEf1lK2wyL8
IoOPryMFBNULrOT8BNE3x6mFTiQcOyKqB+mFKkzYyuBwyvy3/rWbBIhlGp+nfzcu
4V3rSabBRhD6G+JSg+rHpi8hcS0SkZnMyoaL5i/hCTWY+Hn5/OieZYOtKzmNo1+/
V2i+wPAG2iKDOoPZBy4UOAwhjsK3TmHkztWMqEnMV3YNMbvczvvw0j77jKlVDl1Z
yx/STrcvvA2f1M44trL3MzHN4+O+s6cRPGCCPLfbx2vwFFAnneXHH8ynesd5IUJK
mLqEoTmm9qZl5wH5QPP2/jdXCEGQ9UsOL4tLVIkca6hnC8HWkzwTOm/oWDADSR98
Qn5mv3CMmIPnwoR/oB5DWugbzy5F3cMyqtPrb+5NyRUo79TKYmn32p9cnhY9kRm3
JCNSJ1DmNvpvsvvil/u4N+x0jjGFTyF4PkMb5bkd9UA/9H0EXibiXM+1VD18eBM0
XZiRpJ6ofr2XC6pFdWUdZgG+T8z/piH0uOJPMnyZi24Js6pvYyGiYeyk5glLHY0q
7mSBBYo5XzAFNqCYVc9SomieZPSpP2puqWu95YzodaRUFx1MFA5NYnHFoe3wrj4B
1gpk6THFP5ip9a8OUEfrEB9RMrjYmsobA3v36Hf2PkrEXVatwDpa8Iw27nEUb0Rg
N/9tQtC9gMO/ev3IBeAh+ksHJmQlxSu1W/c1ZvJxHIP8DF1iSYKzxvI8iBAxDaGL
gr5MIpZWnf+ZqV0Ud2Lb/Vx6/KI0mCMUrjQ9Dw6VrMo9f4OWO2nPnay1MkvPINEJ
ORdLhYcfytInQwPhgE8weY2lNAgJeLsOu1fdcFEjBrD7lZVvIiYLy1zHkzyn7AdN
LiiXJtOU96WmE77bpkX5rDlk+tpVByYge2GZIHr1yf2ppMklUe2zDKLXUKCjRpb5
HabRWqi0g38+yeOVr5qzqMsakQPoJWBZeTBW9sNJSI/vQUyf+zFYkAL54zSSmaad
zGYEa4xovHJ1R8BbbMgVzFtURipsg/MdEtcOCTYmsNE3a7C2tsyAQo1mjqCsjk+g
5wAomFSxkASRrxkR+bknEZoXFFMsT5raNrmVPq/T6oH1iEByfk/MD9/6ELPqNbxz
/DjKGRYIanhzCXCRUTuQfz+AhXu6jZdP2sZjXwBRBveKscybMiLm5vpftM5jFS6j
vkGNtqKCTfEvpkcov0hSDFItn2BEF+n5yN7D+zgaxUUWexCCcc31gntULoQwC7OM
FVjZ/ZgXxGBKlxi4MWv1/WJZlr8HEUXzIEc4AveHpEcbyYeqq5CcIP1z4qorAe5j
tlG65LJnDFP+efo5Jz6tiCsG+/bE0/Oh2JCTZikziRWSYtPKeEhIUNh5242uIeio
5lGwLnpsF03lMqj5QnDc11GPAENwqe1dh4JKq/Q2ROJguczZoPD8KqIKiDW0hUEk
cb17gCbqc2FCiUdyeWTN3ns33F5wHPSjzHvCNi+xo1S6o8X0RAEO8B4vSAel6JYX
o1iTW3FDQjBEI0URCR3A7GvUBGzhq464xAiunnd4Eb7AmqR7oB6i5IEfar5picuU
MAmp1pcJDV9TB+XFsWYDCdl8MRKVVP8JFxJ82vr4tzwU4kuWe60nqsGe4wMEmEsp
MGt51eTWDJkJaT29uuZLuW8zSmdrGBdaS0OKt/Qvkux44Jv6/zpOqm1jzpAroBPW
QSwvrVnoQja/2FEEk7RrzHHGmLIp9Rfkes7zaEcy9rOO5sy+wxF1vOEgzXLtuwBC
rrT2g52yLkd5P/MqXKhE2hwoxVOcE2ZT+QV+8JleLrDO89ubFXDaCBSv+1MKeCkE
h2wANzUexESBorhUEb/GsLVZOkvfON+p30yv/f2MVFjNM3JsVA6eb1Bhp8bxKSyy
BUuJPxE/XWjZeVoLsnVeHxqu9vfUYVoZU3gKq9qc2OY6MUWjhtjCYb8OKWrRyRMg
XKXI+iTfkaYksb3nCYvUF8jPKAJ+mwi0rNLK+J0DppVEYY8voJNPn3ybNvvp5a7+
X5BXexfUpEFrK6Dz0caWudAXqEIJn2Ay00lWerGmLk04p6rKOz6LNxcR1/K9a3MR
/ZGfGoLwj6jzDkuFF7/IsiKfvt9DvBk+EdY8ceKSiF5xx+hTH6ObP+CJ8ZRuMcfA
wxHVZtxVGA04pxHvzkM/rokk9mjOXp/PaNI+625N9zgChV4mh1omwmRcQQPr010T
JpCoK3Q0bS3RqUgnrfpfitm2jSTwYjiCgeSZKWZvrjX4Cs9nM8sfLgEqEj2PPjFW
uIY4wvujCzqku28/DjVyItYZUnb9fgKszShHo5vNZz6M8uSaiidKzrpiSwBJSPMt
ml8Nmt6bw04tqp/5HwBQwfCyVXgr7oD1N1ejC4E9lNLz5sG78fZlYUYxw7Vv+XGI
KlPc3WGR9Qr4o6pFBugxiMvRZSdbzyPhb+UTu/7AUGgKgLfd+f6l77GTpWX52H4F
AjR0KlzldwjC7if/m9140NRKap7a+wYD6R0Wv1EyF9NyrZARouC+xRv5vbJw0XlZ
JTLhXFQ5QvcaksL8UVZAnrzLqL+a9AwROw6eXfLXCapTiytbr3V5A9nUd5NDTzbw
a8HnDC6q20AY/3lcw1YQBg8LsMJKGpTSGkGPXX9SUbTyMPDxWxOfW4poZ8W0Cy/q
n8gDv0DV7SKrS4IV328GnjA6r6A9JbGav60ebJXOwD2F3QxMwd7CdCHWsn26sj8D
oLYJrTJlTLzkJT+TSsgslblZ4aPJ52LrFNWXgx55PXy4QlGb35k7ru0ROoApI8j6
BTlibyOWtwpKQ8RTmMnCpMWnVBf0RbVlDEBBhyRejl+5HBx5KNfC5idHwKWe+wuG
gI6INZPw0XUAjN6VsVIMhwxdpnq4cjXZ1Guv67se1r+NN9xqX7qKXeIZg/166QAP
JYNMytgYt4y/nBzSDwyQkRAO7GIOueBmnkVuMRHPbCvK4r7/kK9hynttK4WR5BoK
fryioa0gPTkDrrW+WOQybl/ZFt9/k6NYmcdKN7MMpDaMnJ9wGYfYMrHZc5VWNSaq
9slIkQaj01W4hWgbPUJoCmGISgqysHGiJUYNnmsEzF1BAMJudOZtOo3sAdR0ynTT
MfsnPVxitN3v/6NJfPyosTsG9aMoqY03DI0kNuZ2OEs6Box7Y9LtAhJ3CcKQPEcT
vZWDPwIv9a/uUgHqcSl2IjNAZFOo2JhQEATJMrWuQRjABnPN7xSB/rvxviIXxkpW
8g56GRdKLljKPq5d76C59lzBarG2SlS/YLB5km1D4DC4lQFx+v7ZopMVZCMjoSB9
TSYv2FAh3Ww4E44D1FTgFothoBfNOwXnY8391CM6wTndiZ6L481ZjIO8MovI0+J2
a6PZ3a9IpNnCg5YbncVM23/aPctcOSM7vlT10JFgAd+b7Yfi0v97nHKTQGDajkgd
Bv7RPSyt2zHmXghAl0JMUTwwRL4iQkCR76GdZXYnxqqQV/FiQQtAJGpyDK/tpoJJ
jrzerwiQXEnvRuFjLhiKPDWbFA2LUMsB/3+wBs/TJLQqTp3rrvX7hLx+hpU4oVk3
Xg3Hlij+fxFi8mLAn5zMz6BxyWgwUGzk0PxB4xA7hPYddS64rQaUgLq/TDXDdqko
uT1oHV+LkI4IqE/KIxH6pPwmB9Upgw6elzP3DV7A+H0PAbRDSba6hZDtf80aPP1W
0PdKTSzWEtoHGZMsAQemgeQk7f0rodlIS7sNCoiIwXonUAx6aVMmhYdYX483N5on
IH0guwFjS8A7AVZsYbY7g7eTrHJ/x3orWoSPOPGdUX1jMrFvOAn1MGOSyd2NCdzY
NywI2ERX8QYzxBKfX7S6X2BTxQEIaUtSR+q1zxV0F8VJoAVcUq2x33UKJ8heb8Z2
spE2jR5YieXKFZKK5YX8k6q5/WMIbW5VMP+JCjFIC6qnWBTzK7z0Y4xo2QWoHld6
pNg5nS5Jf+2hy552L8V7xCLqjMIlIRgdIqfL9pjsKHSP0a7nx6gE8RKu4mbGKv3j
bI+bhK99v1CYb4BsQs3vPFoz/qdGXrrUHfkqbwHe2sBAYnCUqfAWslHLff+8RVbb
m3eI31uw54tnGHcB2ohWA1VPH+9pS52zJn94fVRQKqbAQ7xsUs+V7RbxjKNmr5yr
tOkAGX00oSzTxBZ9PE8EkX916zNGmKZtmfazvE+Zy60K4L5c3zXLbLRK8Vza+hTP
DmkLOM8QybCjgp6XINC2Lp4etAN/SIfrpiZZz4KalFmXlYsLiDCpWcAyIl0f2LW7
M2u9oe6kM+HS+RX/6n16AbtFb/qYjbsyfa1sDDSnRgd4V1VEVTPHE/Sx1PG9TTwP
2wNc59XTYdEdfGUmWysc105PZdiW8famAS4UqGoJgPTz8Ylr6aIjtOpPi/xlQn/6
lb86MvbNL/mKD50qPsN6VDv+8WvwYtB7qV06jAZQjcVkSh/5jIO61T618MiuYIgL
LP5rEniPnEH/eSqLOe8uEnrXL9sDV+iVbkqAEABfqEYm23FSTH9rUYxGrTp0n/8I
VSQWr6b0f12Byw8MyUyE0D3zXuLIEOax7PMLzo1vqFmglyrsHkfsh/3bcNzFcmlh
IecCQyUxnkonbU1qtS7yZI/D9Jp0Sp1EcFJarLImn5xSslq2i9uj/FwNYmKlp9qw
S7bWlLFJND4N5dr0cJiaJyoHcSKzIm/eB+n8S24Jt6PPUr1xylclz0MtsXCnugqd
fLlXZ1ZHhY/3oG8DcpL8ERJN8NSDRQRGlkY8fVchbg5yGYw4M9GkIvwrtMgUi0Ie
1Mrd9EvZeXV2GhB0uXlN9BHmH6I/AWYdBir01KeyiFfZiNgeHvRdr1huVSX7DIG0
fUm5l7aWsyNYsB0T7dm/8VWJdweZ89upYQi122CqJ2wgy/BSAczkkjEsi2x5ME+H
5XSCjaubbK0ZRfKrulYO3E30ClwsVZvb4XsvHo3duVTH1x4oiW4ULq5cEmdw84pA
wuaXQMn2cRXfrXY48svmxINkg9ldrQ5W8o5sUmdWdbUi1PBlv+dVvvKVsrB3KwFI
cPA6hNKg+3KywCODInRoylYp9urrd80nWa9DRzCzQA1Q0cATj1MLJ5tC0HW/TwD2
xMjZEr7Qzr7q/KynsRCjnPBq0lJi3wLPR6PBIvRvF20QfbgUNzLGmZ2SL5HeixKt
IBBUO4B3Bh/xQF1gEgGD1Wk+zZyRLA4g+QrmRL/JZUMmJizTE89Xm/rG0qHLKip1
WAO/v4L4nj+dnp1X5xMqgIEEZDBHx4YK7GeZXKvFLDdpLcgtZtb+xvx07ziT+jkE
x84Z5843DlYLTh+3ZlgvhanXvkWbuVGq3JyhT55x6x7364sh3gk8DvEp4IgUGAxT
1DJcG/VLzceIxmgGKXqMVjx2DU11cVLyq6Qzd3Du7xAjQ1yaYve8DCckiKxchQfF
yM+z8dpp65HKxynBpz3HqzcvUpeZqE5SWBz7/XVRpBZ1YMrgIHX7F/efhv3loJz5
ggD4RgDLJE7J/7nZtn5KuDj4WzIecM+bSrAnXvceIKXkOuPueluPxJJHopJZz/9G
dF8N7r/foryLsTCnq0WCtAjnlpMjxHZ1PPLbYTaJR6becAw6okz9qFJmRNN5MEWu
BCur1lIdDfZbKUS3C/G3P/oFpI1IRdx8k/IAOPMD8+9dp1eu5rgqhwk2/6pw0kKG
OqDqyVWMmNiszQ1ZlQCQW82/Yxj+qfxkzp+WlOzpsvOF92H/1Be1p3+Stjd8Qzkj
H0HKkOGNO+OT04sd/iWCZvGU7RkAw46LVlyDj4wih+nYTd8cS/kcfqA1NayfYWVe
FFgECRfKyAM6o2FBtDs4TBWXpaXGWaxNa2E/GSxD/XF3qqsJmvufRi0j8j1vpOVB
30GRdLmEw+5HjXk7F9qHpcgDZEMW3IayZIPYpstuTWyXk3F2r7ZHtxOiOYaw8Sws
FwposUlVRj0X6U9aKxU0omlFFAwx3ezUL76xAoYpgVI48BxuhDoorMGk3Kee8KpV
tUx9CJnoFyR6wMTbpe/gTg7g57YEdXEiDUc9wO0UXrakcmAfs6qovVj0GzJQYn2a
Xfhg4nhsmqcRsZ9PR08+jXrhgwLh3S9y9N1dUXnFxKfarQrLKACrCjGi9/wW3EjG
xt8BZiqeN1ychUFWe3ZaMnKVitTMoDcK72YJZTEU65+vOMFRXhR7QcJq9+tibHjY
ugD6Y+HlXEkAefH6np0qciQEMB8W5IdriqC5pj2k+SHltlf/jvktCdLvQG2eUrN2
CqfLrqc3gCIi1ywvxDjbvdvSBrhFdvC5vXmmmk5O/4dIt2flM0CnsH4gUdQ3DPbp
yOyaWjpiCTZKaRDuXJe36MtVfsdgWl9B8cFmFEoMJAhYQBDi3FlHCDk3X3jy33Xm
1TQt5RtCNsszE6LRZ4umxfZwTpvj0+TwzidOBRbVi6kaDbVo5umBVXvffnTDlpPB
ev1QU6IangjC3iVSHCkMJjtkxBhPMZV9aUtFlGNRKg8s9boxHyVu2OfFvGJvdgYX
JuIpwcCaF06isG3Pwwvoy/sHt/xh92+4qNWe+FYDBlXchH+iNY97hlvdLv3OXldk
Ht1CL/4DToOechfIGV5Cv2wC1J4OMs2A4w/7tz6PP9r/gcr7rQdePDv6OSTEbdxJ
10/G7W3Xbj9wv1sPW+9UF3EteQoZRXfEGkEaa2G2IMXvNkpg3VhaSu4Phli7zzpf
oF7odkvM24Lewp36kTFUTzdtmyJd52T4ECugD/BR5/JELqFCVEYFdetVRHrt4BcY
M5wPW9d4Nnb8K75ky2PhAL/PHMH7Ai5y+NhHoebJIs5UQtO5vqVG7ONIiGTg+24L
mK+4XgzRs9wzeOk0aU701YbZENqak7OvGGKgUJcA208uyNKB+ByFUMgpr9EDhpLb
fryVZ/aK9RMSlt6d4Wg+qg0J6Eq26l13RZ9lCkSysdhOu7ET6VrYVKZCV2+glsxy
P8z1f4ueDnNLwblHeuU9Jn/JHiuQskO4NXPcM9dKwgjKHsU9idjz5d7ca5aUpdFm
LgXIojt7YFI2pUh16ZEUybiSp7t675uG+oY5GovlHVo0WAEv/gwJ2c4I1Bk4jjdM
+xREttlKe8bPkyySEXQVxYbOU1/+iAV1JjkbRy5ZkA0HNPKTnmEgfkdIW+bU3hq4
MaFH7573Wgc+pAZwnivwc8g6IQBqE/BzNOTFPRnhmFfBGOCiX/RL5QzT+p7Xpwcn
Q1DB2dSNUPirdXuDYAbwqsmlW9R7YwXydIYNJe7qBGCTyK3XGaWtoYetTLmy7F3+
Fo5yl8uUDROu0HcAlogq00twKXQI5sp5Mzkp+f8dNt9dv4PU5o8NWMSEEaSMgaK0
0W9/KdTiK9UbFdmDyCWnlN6+TiFEacvwNlHVZ1a6Kv5s/9zqfulVIfE2Rq7JL6ot
yGX6JwF+zsTazPO0W6msNwyeCFmvJ2vPHPpTyQEDKLqicrQprISu8AFAmTNPeX74
GqWR7CjdUjGhdcSOVgPNrxJatsXmDCy/ICMEkYuXRDVvyu6peh5X3eDcnSwlkNOj
h/n0YXH6KoaDxne9onQWembheqHB2enocUL4eosJLlBrv9D25SbrmN5/Jxd/c3BX
034VNmIwBlCJTEe1vzyd2NjQYQw21jlNgmMKanehgvEB6xWbhLVa5tqoEYodJwaA
j4+tcBIBANAYgnWz5B78dfuHbU5TNirWwZPieWjz5PRWCwyhd/7HlVP/PWeKnMjW
0HWjAzlE/KopU6nzDgWovJJDldokH+pQqQ3di9ubLEjPVnbQDbWk/fkcp9tzgfhf
hVUaKCt9coyIgto7q3O8z23cwkU18lSp8ZFoiATNzqyHtl64XyzAoWEp6KcvgOr3
LkqCN8lIGax5NnOHSIZng9lHoIxvrWud1jZEfmBzBpwl1EJM0VqBfVlefX9oZPul
jv2DbMJ7G91F/+4a6dZEdCEkJ+FVL68ODBcDrqyl4lUVMug34VT6DoC8lCCkIYJ8
8Z1L/T98wJkCgwTSH21ctQlR3/ERSV5sJzH3L3BxkS5AvxXsphcoetFgMfGicazW
nTUxC5b74gohsh2O4NtLu3iwb5zj9hM3swOxC88+sYPa8WmJUB0D3CE6DzNh0zFg
ughsAoIi31nQ1d5fsx4/Ejax/4q4LEF0/Ea4EaKVNXQP2R9sscUnMXCx05pK9+9E
4b9TW0uFh+2kfX0ksEB2IFq/+/p7JP0iUfQwlEheDBE3F9+G36Y/HoeIULeFDm0J
xUw2Eb9M0ETWTIB+GbcOp2yIEDt8wnX95pnH42rn95BbyRmHVmUfdBWD9GTq0b5U
WOZBwM0qSfmnVh+5ShjOnb61d+GF5qlR4xxASXC5ed/rO+7JpJ79PbNhWyjpEB2G
PHdM9mLlAdsI1dZXs7qXfnBSF3liUaSqSQ5co2PmbkoDznK9Ustzt3WR267NHk/N
UjcsCP8tMrcL2CCYEHIZEI7GFNz2EUS+H+Rvkk2G9w5L3RFUfdCN538xohduUB1G
dwSwMLKtXsD3iguQiaY5uw9CnDjQFPUsDcbmKY5umvnaabHAcsIo5T6RlIr6GTcz
/uUQM5ttuIQeEzFi+MSZ5wKKNnFpCDSZSm9fxmOXOTHcJFhtiQ17bSS+IDHZiGds
wlmyNzXLtBERq8Z5huZMUNrTnzIB7mUsXtAU6z2FaVtXPbl2Al0kvLPffv2HwNhh
67AXkITrCUsXzIR0QWyYUtaAFSqdQBsyr53PFtjLefPfdfZDGvqRrc3mwxFf+pnX
wuNP8grjZD3ZcRuMmHsEDRpW2VDMwa919A+P58O7REtDpr0Sip1y/GMSsDweS/mU
lixQRXPCbUwQjAl/MexdnxmLYnl3eofJshqNsLBEQusggsJjjvJruGmGCw2JD7BN
dnUTAig8TI5i/aEie4XbXPY93iXyF/PTTxEhEePyDcsxDhZd6c2E7KLlV4Qow3nx
mdnSDJl4LToxOWajCvpP2VdzUdrec62xCilTynxbuSDKvBcjizXBs1xPtiLOAfiM
mRtHdXgDJz0vxd7+eIXzXMqzudQucDgZ8APEfsW69a8tdYhlvfNa2h+esdtuFST0
eqq7LJb6LTuaPtfeyo5NSuECycwSIn61kmEr3NsW83p+5+bV2uEqT+Uaq0jWN78h
9wAPuibBIxBLcALPCrd2fGVClZiYEN+GqcSu8ruDvf1plCwaHtP2kh6gGuvFTg1a
DStpola3SXEs2zzait2lVvoQyuKtr0CWPAnXOsM9chNa2GZZxbhHtlhn+Xu968Ce
4xEoPuZtwUgrKL/sbMt3JGSht3diRwn5fzMLd32PnB8CXqFWktNa3Pme02OLWfXo
OWdLgd3Su9tkCPHk+5+oqci4Hjrj0vJhUwqPcYyZEaI+n1HATOv70XAo2iQuCSGA
YSL88yQVOBk5emGMVDBvZAVyHHMhWDOvIOcqxvP3QkAmAlSOvS68p5kA2Ves+cmu
e5sgFsAFHn1eSoqA5GiZXRhAap5VpECzThS037zGJsCpZkMNL4dmcWnWbDYI8a0U
rRsTjgE/26FqdA0tPLjCyK3f1LjYLfXMcgwsmsGp2LQuf6/Kg3pXJ+5K5ARpl/Dc
OXo5NQglKbW9OrINGf4/9j47KVH7BnQodH6OHgfFpngjBmPDWZnFRq5UnDTGNB3+
3xQm+6aiDyNnJDHOEaZA43LcSrzis/CtPkrAKTG1tyPAhwh6KnYSymRTV0abZkp6
rr5vuHAFnDM1A6qw0XmVTqTmbA6fahHQ2oU/bK+mCMwrcl3XbyQ4SXHI3vem7oJ4
wd4M2Zf0Tncn5vcFjoJV+r2DLQBMit1JcS9XOuHxaCPbiXj/k0pxJMC5tJ1SHtlP
2knf8z29mKAXlyslFAmKNp9uz6iGsIYypW79voWu40S2mmYQe1oWYD3rIs6Qs+LM
aPqhz98gOkzJ/pcX2jIB2vJHHvBnBbU5kZnsDIrZlE42u53f5AgmZneyIfHz0agI
aU2awoboM/z+UVePdEZCxuh5fvXJ1Zd4sDiw/emndjcgzYgO7izzemRy145rsl1d
olM3kBidFLWtzuxyH4R9vJ3DQ03DLo0sfdSe5v/+XZBWv4Lt7Z+So9DSYnr9jK9z
kPci9Cd3BT4RTZ3Lc+zEIxwxr2mFmUykZvUs4gPVyjisKar+q0eNRaYb0/O8OTNr
Laf60vw7lfGQnPTG+inlJc8gnkkIz3kmjkTQpHh2HKeP1grGRsLyN0bOnc47m5r/
reRiphozJQRn8n0NpvVE36Pt2tjbZ5Koie92cbxflSdKR6W1ahnU82jTzVromvuq
Ubwzz+GMnhs5M3b4+5W0tgpwRRTCCgQ7EzHAQOa4VLD4rTz5r7UAofcE0T9y2bNM
UbTpbkm9cIoRSnxunCr2/aJ0IvZ4MolFQtqkGTjfeidMxrjDUE2ku463CyUL6DsB
gm7SIqsNbGuE+THqmv7hBo3G3IKuBXZOUFs0WKBjjFhJwdNxxwuPybRWgOPwsH7O
7jvWbFyz791wdb9/MG3pHcBSbn4AwOxFgsHmEKjpHB6Pluzcdzn6NO0eZKHwPnUD
XmY1kWz4gEz6jxy1yfIxrOxNDr5ZvBid2sC+tgMCy1SgS+jBjYdOev2cOO5Dgjf2
f7qblyF0qLiG7K7e1ZUvXVoPTj8oNkvvBLocn84RwArUtYXZRpKt+TvQAXpNbY57
L3uURxxVnTvZOvhUsY4NDb9XxTtffMilu/T/hkOHV3sq98mg8+eL7kWKtw54pJiJ
EWmC4r99WicCXpIaI3o0B4NH0oDTIJdgss1Dvw1K+fPfGRPvvDdBqXyCqo11ApdW
+2uyJJx5GzK4ep4hgGDzJg95L7m92bnHiSjunpJWwma2cFAFSHtfazv8TdKR3MC8
OF/tsgWB8IxlZOtmVFOjsY/t1ajEuzLomH1yIfNoGwmeORoE+XtZ8xQTWzY3PRSc
hAVHgkT57wuGyF4Ub4FQwytMPUurwvLvJAOlbQVns/ldujIaTwaAH6aj/u4aYLxc
0ph9e8fXr6izwFhM2mCOi0FITcgUiBw6BIvFGsRXh1EM16/inOE+uy29Lae7WL4r
+FNm5PLsiV2RzYzvPTMSegxVQzH+Tq+VzFhH3qnUiIeQfO2C55w0G50yskpzTS5o
QuhjDibH1y3tM7j8XkBAVpHwDVFV1QkVv1n+NxQJ12whiB4PSgTg6OgSZGJr4DVb
m7azxXB47fYkKcVOrpi+T9VHlTzykDQOqST445IZZ8fstKfiFYd2dBtBUwk0Z2MJ
YZKBW2OdGEmeGgnSAoJD3UQM00saInZHOpZt80gMM8MVQrqVkZbMMP9RVpcFh9uO
ZgpeUQ7CWERo1yd2U6lsTeuNiugrE2LflUYibFIPqUkSLx7rskjnrh2O/iAtmP4l
omezzLOm6xsyRLrDTQpV0E3txOsUY+oCWt/AebKSLKlnSMoC32dzAgZfUuJCgLdS
kvdXRqM02G35mkpqqxOKbx9STkXy5omqdNNc8IRrBq7lPGC45dQ6hADojXkrhWBX
8+no48NTx0WXc7OFbN4qheyW8A3lyNiaBjuMrBp8T27Zp1afTxRItgeIvCYGhzFl
GbU3S66ctKWwHwBEKGdW/hQ8NVdsrDw8UZsPhEhqopmcK0XxYGGvcL05pn/NRBax
hI6CPkDU3A4DM1E8C20ONWKfqtb5u+vUCbaXZcQm1yj8DxVHIC4gr2UFvQNY5q8t
NzXErhuAHGF3ET4QQ2wqg+AJAjRyqB83q1PHoBy9PFpa7WL7nD38LhnpAblSDfm1
11Xw4JvoN6CLsgcJqzfggz5sZdakj/EcW4/2hUZnbdBXxFnzJ6+F/dh6FnTMtqXT
COJ2mOP3cJGGKl35JeoPeVBy6hjOQ5prYidyxPeBF2dFbEOUnjW3ih/SRkCbPOuQ
NURCPZkVA0LcCa9CSscD455cF0vBW4i2hRw9WUzIFyBaEblzijCnUdEZwukOORfT
h1ylKZZwhOSnE5zEZ2l/r3xhZ3bMraJzckLzO2xpAevud1baxRRhH5cQzhdHeTWS
wYmmtrjlHoWUDW1QHJnQWzMSzAoTq9bdoU4Bnsphvhhe3yxyRk1acCVYJqfqtq2n
E0n2cTXdVtizn5TwPBFMX+xuPomazLW0PkXaKJ9ri+Y4ev3qpd7Qn/nvcSqJfsvz
/TvV9JFW+g/kvWtK2dbHJ7MK3sFT4rcCfk/cuKmxeGoSl61ey/Kij/yy4wzWJhSx
1xwe2BNrqmQvR8tEqCVk//MfzBpWm1NLMMWblYw7tJwBwc8kT3YKScdk6eEz6yC5
4396oJQstg7wvdQedKG/nmNDITNcOVGoMpMLspoP9UxmrXNCejhsa+kOIBgelVte
SQKqY/rBFMOIOIredhsILmS4gdr0k0cmXqFtgErOJBxbs8tEXO8d9aasBzcl8WJO
nPRbKH77YIHhcckhLNx0CyHzxTyvzEBQPqrsNdixO2taGvKNgszz07NO6hoAQGvT
we/ubIZInsib6v0ubkdOHCdXftT0DshDvuDsz6dJrFpLLx3pxrcV2T+FEfiybOpJ
9l8wWwULEB4rDZOePJGbrJSoQcT40nK3GSiNoMVO14NmlITsd1vinyCjiOMZeMqg
BtvB3KdIYWZyf8LrtDAfr41I+8RRS5VarzC6lzwn9enyRAebJ/UuUEz4REBiI/2S
8Y8iZ1z5dGzJH7KCTmvjBIAHvf68S5E6o3w+yn67ED1TwW7bX4jLHquAuC+LTIN1
01TwnapNmGJF3A6km++sLH0974VHkBsvot/FvVquEfOG3Dk3ianUE4IaiZX/TVPf
8chRIZzEFXst5Ik2kJHZfVwYqjcGWRxn3g6TFa7+db18nEA3VCQqTMLbRyrI5U5q
N+u9tzln8XziApOrNdIeRpyC1zn5+AypzXaUpSPBOd3M9nacbxe5kn0J7ofrLIVB
MGK2aq62CZQIAQz7xo5/lTZnmHJgRm7AgIVHN8W89ErKER/lt2jw3lHTdyw/oDMf
Lp1nxfjSJasF4Z2zcOqizHYlKYil+u5Ga3JmV7UsAjSQ6AZjSQ+tFuVBx5XysrMx
Rjh8DrlBEd1OVLCHRFnxhV2fVbXyZG+WdkkkWEH2y4AGSEtURT2Y88BE9oA1mIJ3
JU5RcfcHcu8CeywnO8GWOtnCa19UL3P/oSGNo6+r6OzREjmpPObpmTblmoRmjFCz
Gp9cRRKUBy6ZncEu9qaUhWr8TbFr5RI1eQIaQjI9CBy+IjthYmZOsgI+sQeHrfTZ
zWuhy0mJ+r/EHPWE2+FcNCRj93gWBiaAUNGV5gqQ98cAKA39SWbPzzZh9qxwz0vi
CVFo1gau94KeeZJ/Yj8cMW3bq3rRBMijC0uizoVBAIJoLW2v5RoYLk5WB5In5ZGP
YH+nMyEjYxLKeH09D4pS+tKrM9thndi+7Waf9Il7W0cHWPtDnE/IJBbd6ZXaIhlD
esrbn4RH+DBOCsjJYdvbdL0XKZLm5HR6igXmmapxN0cnzBwwZEMiwrCHyQguv9+L
Ib2qKo4U6uvAe5tTh4ZjyhiHjmTc7pr9UsyzkGBd+OpOn0NJYCrOPurZjXBb7S9t
zmeqpqLnAN6i6rzaFy6eGs1Y7Z3qK722IEGEqmmkXKGZpRZav0CtRf3Mg6m1kNdG
OwAg9qNKiaqxJLhhBttEst5q6wzQ06VKY3VsNW1JJNZEW3ANThdDRe0hEbOPrRaK
XP6VGJRaC+MQKBAKzPTk4JJMN8WGLqPZYIddiVHoabT/n1EverkB2rGoa7mki5H5
ZZVx/FuVV85EpLK++uV+0fTGR0bW0R7O2gSNdxmJ9riX6LtYWz47xKGt24Y4cc//
JhrLp6I+oWwd7zj+OUCtTqkiNvlot3Dg6/ubKRgYPz0lRBnCu0hRf3kJ4ida9mG2
BmtsJx0cjYokV/Rb9bu9R6YwW+7CJwC7jluZ56KPizZshG0zPfwR86tSYAH3Col6
GEfPd2svi40WbtP9wd8QgPApfBoWVrc1IDhiS8+v4osOSETdIfWzDQXy5ZBwoWD4
8QKL5LnHILPdyYxQ96sEQjwnI1gOMihEAFM5/BYAVxokvHDdLydbYx0WBkURAoNP
6Eog7KeSDnhd9yoQvGEL83iXNdWxXxo4nTj8ueiKCjsDCHbsNi+JT75fUrNbTzkf
aziRbgfv42rWqqX9C+45obig6n0AiBizNowrv1ZhPXxPTqvuHkxACDuPH9MUPYUe
LZ5ZzHLCbhgDfAVxJzac5fLzpD5A8JAAlyPTDhvPQvvPl7i1Ap5m41MipnciIYg+
R1oM78WrY7kBsurtNDiLRnzVcm+K1y5RSOqJqSew7/WJ7TlwxGbK/kv7zSdPVGFF
yDIqSZwmaUXj1o2s/mPz95wdUfZESHtnonne6YjNyquT332anyJu7D+j9fZfdQR1
YYYIs5nTkEe4WEmyrQ9VZSJ199wOD9wIahahBsmBepNkymLFxSfHWGUIVNlBPc3F
Ju+ig6Sjqi8DT38ZX0JKVX9mv/vXwTwiVxBlj6yNgMoYvHAtQ2E20TX5ratG8VM5
vFb7Iu1FJg3fYpozGktH/6KW5Q85vsT3EqKzk9F//MS/0497nW4lePioINrbjHPg
BB0XoWWkOV2C1OMD179IAf+WDCuDgK30kO/Evk534S8bG6KFpE3A3SGtacnRDMty
dLrI4YtL36BTjqq47ZrDpp7fh23Zi7FBEuj9wasBz4BcMC9aFLxxBF3bA4OZle3k
uBr4vXqDVOA42yBTSECmHKIaRB6PTMZFEIqpFE8DtwQ4iMj7bkHS/jlCle5cE37v
TQ6XZT1j7yXH8bbwSoHFbnVOgy2rMmtIBFeqLswE1IYPKXX0z7eQ7A3GEKrg0ZcI
TBQ7Nj3JqJ2bg9am9yUytQYWWET31kET9EBdX3q0zf7MI+ZZcYEZKwRVtiHlfTe7
bHJ4GiLkSs1UASS7JxsZYEnpAJHRBggeKY5qM4Sp/l6TA6Db3Oeu/gYKoZ1uXL0O
B0KAjuvPsrmIPTI8y9urs0rg04lYOqmFaJwnAq0GQsLvwp5dAdSP6fDaxKJtUInv
o1wDSRBzD/6XMS6vHRjg0nFZcSbelO+gYpN1OfkrzcTTFLHTm44A/0eLhNPvBfL+
rbgHA5cLx4De8Tt2OFPNX5t7luq84FwYl6hcRmKo/ti9Op7TeEMOsI81tZXQpE+1
MOR8pQWH2vfGBb+nSAy7Vnj6cBqGAI4ZoeW6kSxNoGfNPlInLv1OnqkU7TZPaAgR
Pq5JJzI7D/r+CRDRuPH6UuAS4dVUL1fxDDfC85UjmUI+CjFMdWtAcFY5iE8MnmHu
js7uLEL4EWmDaWSR/0eG8UGfHS7/9ikzDLe0Xux4yCnbgiYU8isC8gwlTOOLYFD2
EEcP46/yjc+pdZt9ai19CSfXem42/nyUX+lYk5k+Xysp3kdNzVOkzpOd7TYny69K
TrmAyhekojqRJ8alCxSeLkOPOfXocpFGZqsnjvUPmqKp/J3AEXDtJl7JPnArNXMg
DLxKQHmln+d/uR9F2qd5ZX/qoopwjeIhbFaNusfjqwJsRcYjz5qFAVOSUp9HD2e/
i7PkmUMjDhtlqnLcHzQKesT/8ddZRz+47qXAl8Kj60WlAW6H/cfNrSqNplwmHhGx
rgsqlFAl7PpSUwYsda3p9rZa8dOFIZKoOMzaJ/MBAj7M4IkJAZo/LUsXe0Zgey0P
Q7Ba+IhzNUAICoXzxem2VpOH90+sdNKYqHKf05XVtodlVAQuVG1C3+7JtISxTObx
Oh3hsqpVrvzBMv3PYjSB42gNLPEdJcU1d+iTOGD+7iyeQwuYJp8EHUYSdQ56NEeC
4AKuEyetIEblI6MEqfX3q6YrZs4KlijqlwRHbo8nM4OOM7XfIyFVSYLn9Z+6nRYY
WyMRQ1Q7PQ83r+Qo8unzOqZc8YPLgwIf9dYVvnDtexe1zyZNci5yOa1LFB3pK475
kFSogWxR0PwTKLRZ9lrMWBz37zUiGW3Sh3DlZb9NCbGGW5SxAa09PrPp45Kk3+Pf
Ms3l0meB1frKzkOF5PWB3E01ula3pZs5+jAM+2wGb08mOJY967MNRc0dh5+PyqAU
pGusCCIjKI0QFlQQOSQNnuFH+Rt0K4PGa00KYALQ0wtOIxh75LVdn9bwN9SPYZ4u
Wb+vAqYjxL+FTsIQajzehhbESA7tXIl2bFQ9l/U64eiobiPvRcOVO+8iWFIRTIoQ
aQVVaeGT2v4GovtMajIQSIi4AeqbNIbbjUPUDklei/YSwg5oZ4yp4pZuTqTmdbGo
5pmNBTKXMKhFbUtcClzS2WO7uUpVlgpwhj17+++LoOWH2yXyUW4axpjHdGHdgqGx
HpMnl/q1M8vAACxHgXpmhj3wm6U/RefwaGUUy6esX/67GbBKT5GHQ5Vn+XZmebg8
3eS9Z6O10TEJYOALqHXVcZlto+mjtwLTqqKY+3cpquyBckE6Fipn3JWeNr9vyq8o
lOwyyL+DNHy0yK+nlURUwSq6EkjzyOvRqYt8yf8MeSIbYmNdXUcJF5zbtTZNGoaa
90Ypr4OO+9DdEq673BYPq/f813ogFGWuPZIgETlgjPlz3nACKbi4yjKIr19BBe1R
jZRQ1iDPITaxBH45k16DMA7ZQ6bRCPufJdaMYwe+sGs7TsxSukl7edYB+JxDDI5h
KIqLT7dNJZpMaqbBr7VoXkb1dxl74uDaAWJ9XqEYzHExs/3fSQ32oQEtPrKW+ISQ
I8LOy0YoSCsAHYxIBpf0UD7Svh9s6A0XJX/JbusfC6VrTg7h5qXb1bDxubsS9j8R
gPKYj9N3wlLUQmkFgrX8E46Iudo/2BfVPf/wzfwzkt7LorMEPUTvxuXNEBQ4KMiA
MUgl61WMCc1zoSG5XwBp1c3sSHbpAETUOXc8b0X7vwB9TqeE8GFnBe3eYnq14MGF
34Y4LlSH2L5KVKi2fvsR43bIzRrcQk7g/kEp1swrPY2KnTuPRcclQuiGHapd8o73
+RBPxY6DG4ySRKK70kFsdoy5UKFG2CKnKvXPdln2Ops69NOdT6MMEbOIiSvpkJI1
STyq4UCtZiGU2HRjn0O/IzC5LJ5YXwDWFIclyNAW1ASpFoq3ex1xGdYPKEMPNnaE
m39GAkpugaJzlgS+d8uu4uug5oA6+f4HBT4ZwrevPObgroI/74VtBONPzRFeax/2
9hDlmSAX01gtl2ejt5LZvlFxQnTD1Itw39Mx+HgUYHBQMsKex3zKSHtq1yAlApOB
d5jucIJh9NGRHFXXZWtpaDdRhUC6APMCoUvtspQVIHChsouzP7xoybnKKt6RrCMi
0TQQro1RWOWCVsmX1A5evGpgDQE0hHWmXhOF+25jwwzSfmM14de2NB8R183stCGJ
rOX5GIoI4vBsJiPOnelOKXq9y5g/46ytT0Q0qd8v/HN8QkOW7Me5KqIktxgIxHWV
9Z3wA8d5SYiqdF5iQ9gLeYm80NUcBxMYpZd3tTqygLin+Q/53SLfG0lXcmqYPY/l
cUzxRNWbnl67vS4fAkRkD4e/ft89uvkWHx9bX9MCmIvVIzfFUjyxpz++A3JokM59
XiT/Y85h4ZOSRkjI+RDRHu4pDhy55RkUJhDJ5Qe+Q/oZpw6A5Eas+7I9ix3RW7R9
PNCEA0sP19jnCoBgwjXNmB3WSoN2ZhaOPwNaYn95jFzQtBbVyJCGJJnCl7IHr3If
fVaG0D7zqnBabxJFCuARMe05gBWzPOhzp+Lq/KESxEoLz6f7gUCDAzzAjhNHMIV+
mJFVK3SHC9VN1HFw1dGsANoneHFGsT7V+6po0XDQHD7vA9Z2wufI/HbV8bxc72+M
r7ug1PAODvcPG4+imt8ALTvJoshDAnW4N5EtpGfSsVOs3vJEEFMHaSryYNrvlkgU
tbmqwwmmDphUcblXXSovOlSFGjEgyW2YmHDBeVXGpZhzI00FUEbwvWH9QJ2R5it/
QZj+i84VsXM8HBJ+UfB0vcYcdnIeKueRGoIGOZOGHun8/XDJ65ni6/kYqL0o7etO
GuoVvApjcPMLA7PvGrl6ja+4ZEqW/fPSp9SfJiomJsZwx7hBapNpZycbA/t9b5O/
WnZOl3H6PbfJXOSzbHlTv5yxupM46xSZqrzug17BPRgJa4aBGTgAzQaBZczFrmPp
2UNsXe/Bmudor7Ec7wsJPyW5S7fz7FWwXKfj8gnpNFxzXFTdTfy4nZcL+/zLdz6+
O6r6RyiDV07pr3Es+vgJE70d+LrMR+2t7opzdJwPVatG5Emuy/HU2QnoR94bLvfj
ZfWO5B+XRTZovm3fbEUK4A+4PBlTqK4/4zDBe9cr6cJy7SvCUtjmIzqTL9R3ZbZp
waToIdwwXIzhF55Gq0pXjuSySKIb+FglVG8Bf/6WK0CUsUrM1wtofXZgOC5E8GKv
33sToj3+ebGmKu7FG+eC1BUUt59raNUmLFdNG04XvpMZR8W3C3Q4tCg8e0W0lXKE
ot48JtHu+B0JvmyMQWg3NGL3hw+GWgSv4EZArF7AwfN17utV5aGA7rjHQYI71Z9K
2i48Z1fJL7Xhgj/7Dj8b2gSbtsKHuE/v+OcrOgWJwdP8ZWyXYHlqJjrQ6MCMipb+
phkJvHOruCOdNgOBzwoZQSd0J3vpPIUHXaJkLA8dgQ5yyGvei/TjPRLM72xX61yy
Cp/BfKZGzWSnvx51b87MM/jqz1yA5zfZAOO5nOypctRzWRjplUBnwJm7W6FLOFN/
w3o+DSHolQOumWnDD5IxVGSbzs57Mv7PHSwDT6PktPQLOnkXIIjKX0vZvorpEFnq
p8dkd+uoIZK5yKbS9w8vpBEaNeCXXmH7LXJ5KgTQeXeALrdKZb9spTYtLs/FUgrJ
anwqtmb5OYk7fryn6b9/yGNKd0GtEReEQctXt2vnHXDNZdouF2dCQ6bA+zz8MWdV
H7YNHI3qx9lWymqy00K1L7tfpTe0Iy4Mcn6NmMt14OxVEINcdQ8JS8asFLb1D/tZ
swpU8QY0KuMSTJ8cXjE4U3i06eOfVdeb3CWTZxMkWdSDuSXM3AyBWBXwyW1nBFR0
e3KiNSfwpaO/ISJJGCufZOnvVZtww5QKtLQWHXF5a4Mv3GzSb08SL38GGpo6viZR
xUPs2UCGHx5V04bmGAP78QXODq2k9qBVN2mI7+f+wMACSk9e78afcLChARwQTabe
bZOgtiJlqtLM+D4Zg/aLXNuUHGjHUZn+Epy2jt41Cv/iSyLjiHKgKVmh7S6aoZfe
29p4IupoXlvXCGcAnPjc4X/5GckmdHrDelVkwxhyosHgjKwY9tKf0mCZW7Uzh4vY
CXuqURt3GPOelSxV92We2KDH8aFWKioPJ8lYUCiisMjnmZ/eRFofdB+hEYrb91e7
58LAW65bWVUchkIlOp3fMbO+2gHX8wpNHOnbCvZDs+yebniprqgyaO3ZelC7edU8
ATJ7h4BxGOYZ6Hkecs0xCVd9Aapih5mehzyQW9NSZkIDcqeeK54HLVnZIYIPew0Y
PemyUpQ3q1hYwtQSE1Mx2SyKZeKIce30FDO5QdZhOKAQkG6pp4j+qnHAuzo5bGWi
Ub9GNvJTmoNtWGyv48QTqjrMOGnu1j8+ZagKjROaZ+fqCqGmcq1Qu1PtYcV1nPsO
7YMxteOB3MQOPM0+fyX21Zd+/IUTxZ0WpeFQJgc5EyztAQ/To+oPqnl7nbHZgmyK
xaYutPLWy4lJtlQ6c/bbWNGhQ/UYWN1sfdM7PitNIpRaqZzUN1rwWqMr58pJpr6K
pMD6PPzNaa7gL+I3fnMihOiY7ORz4BZQW/8NRdk2W+mIP9piENai2n3/6nZdfzQr
83ZJStJBId1/9CtIT+18q8a84sEzgpSvrIpkzK3pni0hPYUcF5eNYMVR8F3NsCVY
k5F0SfJD0SLYgyoVAvAx+4uisGumGcVxfPoUeGX5/VJJB/BJXiZb7oA/hFSU73Hk
gVJek8iRt+yc1e7crc8RhoMvEXcpU3l8r5TS/l01Cs1Ab75eENvSC4OnLhRmc6IE
irIXog2B9G+52k806MBRW3dEINjPvYn1ZGztsI4Lc93GpixVZk/Brjz7BbjcngpP
CJ1eLs4LV4Es5w0+ZmcjqbU+yWKOJqd50tWTqbMwIO8YDkBqUWlifsgG6tIdGhUX
Q1Ok3YSY/Nlk+gOQXaTdBtFGS1l5T+STtAc/JOAOg6I86IZrsd1cHkG8kQOMULTN
4BuHnjSIM/qgsUcltiBkLuJSCEo3fEJrwnHVtyLI+y7zkNgcLqUH5IbwMNpigdyw
rxDj2Mk+T/vqTjrJzi/NdPWaASwz04Ytus0ioDvW7MuZ2BtRt+tbjps036NKF5r6
bSgeJLO88eYRUIg2qtI24UCYMfbR8jdmqB/dtxgGYWWZijuJzR+nAok2iBqGtd3/
NL58V+9oDIyiunzk0DATA83r402A0lJ9mmYlwS2wcB146a3BmZAW814Zaejm+mwj
hQW4U2CwQu3pfRo9McV5VvzxoWv+VeV8mZj1Knhy4gZy2iXgJ4sRleQI76sd41PA
pu+Vu24RcARz8jomoymfW9+jlgI/4UqmOfyWf8iUKD/dk5FzNcXyDw52W87Wdwwz
ALsFhnDLwnxsNs8n8H7XkDqsn/5salJt+drj4JpC3s1ouqeLpZslff/8QgIzuSvB
JxjXVtG+ZWZvYXtepFZ4YgGJB+sLQahT/4WyJEfa3stsGKbmrOLR/ZU5FeVHwiD+
`protect end_protected