`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10080 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nnJWG+6JMiXgK77Gh3gyM5U
anW1IIHecJDlzcHq+QPH5/0XPSFHLmf4W2T3zUMDb9U5sV6BzITf6uP6LAm4fb9n
sFUcItTLcJmDdKvrVxr2SAwuwtYQ7tje/bdBvvXAFRE7HqpQAWUUcVeQRuPta35c
2zcxUB/EgjYo2T/a3PtUTchnsJmSrK+GoOfq5jLxALGxdT1xNwXKu8kT2Dcvdc6t
WxptreEirX3ysV9EtBmt+jXrz8E8gq0d/dsFNmDk1HizTUOhMbwVEik/XpZAmGP0
iwDOlB3RIG3O+56vwkTiGazSZL5B9gk6PzKuvQ5U4F14l3W0DwTViA9NzvK9gtSU
iP0q0ZaMj/SAR7YwefV7fp0wwVYb0uLBzM4OFh64mPCUei7siR/zDdHRgWqfrrwA
z3OhxEJW+nmlJCRqZ8OYH+TlU8sNqpOiYwq2XFhX+k1C+N/QTFbmLcpiolc/8Rd1
1RRPX1G8IB95kpKH72oetPdiSe9zpaiK/B7qwJJ6+A9okfE6avcw5jsHBRrXlQNP
9iqpTmWsEUfT9ILOus/aJu0mPb39oY5TtHw+VoYhpDg1xM3LikEWoB/R5jsHROaV
YS5wNXINSYgCeYwE/+9pBAiIT46qKw+OR6hfU0U+71ek2axeHatz9K1QwAME1UZ2
LU6cLqdIpI9gzy86KV5k9eccTdXB3qFvkT9AU0IY4fnwG+7eHK63/BGhOEk61su0
aMVjV9rXsxh30nJ4rtyxrzV2DdiHw2G80rgFExcEx8tg+pGxA0ZpRT3eNOzKZhdj
7VokNSoXVcu84UNu5ke/K7hNUqRmcuQSqzPxhYM/dZYusMs62doJt+ayYiW4vubo
EfGO5Jr5PyTVRyhWEhFlXQqFGK4uzENSrzck4nnJKDPfSlmm+adxpzaKDRSZiuwZ
73ytIg4m3wT+s2Cgvnz9uNRdJg4XSu53yq8cKbCK8nJcJnH4fY8iBUJ/imusWrRJ
CMzyZXKrrfcgjzWQIrxs1o4e8T29SeBNGeNAbOlJcN+/xw4WCOF5iV9V4+7RJOQI
YBeJXM9Ee2VYue6+RMy+wEEKcIkaiUDbM0FBxwHL2ScI4g34hG6B7jqGBwJGi9y5
zVBA+Eb+HfUFCD/bBBXFsglLkqOfo3NJ5DZnKiqw1dra1nWySF4f8SqBdqnidwvV
UW9hFQcQX+tKou1yvHJVa/rSZtS94yTZ4dBjb+F4JfX8D8f40v2RQ4eNCyFnRTR1
6nxgCRIQP7h51mAIsKEQKF79V/g4wriFe7ALhFoywMXMjksrLGQMbzQBR42V1/1q
CS46Aze8f9KE2PigoUTEIkppNHeACNWmm5fqFN1heacSMngxxUhwfo3DiJNEzY34
b8MC91UVVWmiKtQnw9D97Mv9Cg+hq9ex5d+0Pn+wFOAOc4HISKk+SxO6wtMZBikH
grtSTy7V9XV1S3N8mm4ObaoEG/MYmf26mAJPpyjqzKeelV8O7QG0XS4AzNhjwcnm
v2uwSzV4bNrkHJA2mgcg3zKI8Cn4ULqif5yWMZNyJzmUVb0nTxHhMKm/MknCFLAi
P+y5lSHNR1gifDrdpbdgkvXU6E4A3G3oj8BkBNHnMx7IhcMTCi3PmnYfwG7WwqJP
8/Lp7e/2OnYFh7IR2sEk+YvdGL9sAGse7ODCJfYqO2UjWaq8fEdQF6JngXfXz2Hm
7SM0470wSePLFm9/MaDghSLGyp/4kiko0CHIBAty0wUZBI4hLUN2MwZehj9Oq1X2
251QYg1JCIHNI5l5SCyV6wz+gZQQt1FgneXiT4Kw6lRpsje8HNEziv/C74M7u6Cw
8fpFrUQ4+AhzC2uh6jVBRbsz9y5M6eaPy3qRC3tmgN9NqyK4LMzbfLsi08iGyr/1
5RCCYOL4suCRu8E5o17pvgQOAeLJoS058VQmDAjhZvGV9vIxhXWoO2nv3MaQJu8x
3U7MjuRnSQvfl0M6TohHUIqTCB7CuSXHDBvHJS5i9BNNFIBiEMrg3H6a3e/nnxif
ylkkYZGeW/b2eNSwPxKyB21zJSujnUsnm0UESUo3hQAcWDp/N3ZyfS7QJAqqo4Gg
jC3W+D+/sj0Wk0I27+n+yqm0s7fLS6nbg46X/Eqrf2kOpsiV/3L+shV1BqZThzMM
05isKevW5YArhebu0wGGjGqzHY1u+HiV1s5brjl1Vi3kCPiCoAx1Z4tK9nnq9tBB
rRs0HSOHviJbacYgj3k/mjtDlyDTFYke2qXK6Htkv69yG6+pc0dBBFeGZRmeYj0D
o1nCgXP1vJ9bY3/fQJTKPpa9x9/OZj/vbZVNLrTq0xm+av5jRLefUxsZQKlsjb1V
BrQ/WQySl9fUmccuJz15qOECJhaDiKSUC677QQP+cZqWfrV7zJ9g2M/zE5yWvM8F
0woxTjenoWEwJR3hJtM9rd+GW+Tgl8z/E943ED9PoeO4o5UjDllR3RxaCk+s2e1H
H+KdFnh+pO1yYu3fmN9qeweYBbLi9SPgXYNtBdqU9VkgSbzSWW/CG+Q1flNTg78Y
mt8qI+W677DMTOnQs6TbawgOTuyPcPo2+XfEwlF+Zxu5C7gThGeAhvrgK2Pd7fFN
8uNC97Fxj7RaY2NUFXeFOCXxBZaYXWsXJWA+8+cUzkxKmA5VDd0E/UFesjEC/Gjn
mtX3lXHS2k3m9iJE2jpkuksXNPXHO951MkD2yQMq0UH3VRC2L9xAlyujZ+37ugVi
PgOz3UEAMHfkOjmOjaRIDwv/owYdxTJawe37F1Fi1A2ypjn9XJLsslY3uZ+2gmLO
BTbEKMxMjiTOR7GljAgsmv41zZieTSX+w+0oHbkJsXjk7gfbCHDeXYXVZVZiV5Dg
WVhFr0xNc/KTBRLtBENNxpS2EWW9NZNGLjea1AGE9GCyOEAuovCHdp9xSooXQY9q
wzkhzEI+PiBm3K4RdIVHq63+5K4/OAMLWCo+sBetuwl5nhbJfIeJYcSaN/2+QMSh
ZDvCWgN7vsQ6ZVpHppvL1unp/Xm3K1LQ/erw/2rZEtXy01Ie/DB0PUc0DD9/noJp
XXjpHohd4wUDpE7GDWsRBPGhYmFGrRuvas2yunpfWKyjs9/xYrn2Pp1NAluYkPCm
IzozbxONzJMKXrDppEf3a39dYXLB5NNpizWebfPreIc8z8x+87MhF+j+f8QnnEis
dD03f1xsn9+Y63QF447ke/OTSh2gUjEZHuHzJk7dlnamROENHEQgaHd++rmLValb
XohmQUBfObKN566xw0yRvdep0D4REd+mjfU5kRvUEqnsJkoDLY+K7EIOI7DCO383
+Iw1/htAc1GsMsY1k2Qav1cMC8/ezwQTUKr8JdVXieoQ8FfXeNuxeA9P1+IbrpdQ
IKTcBeQLMg1g03CRFZ8uME3cACvyIpLZiZ/EO/PIjs0z7394IXNUZLsmviV5O/Hu
Ea31Y/2z95fHUmEY1pUN7ducTXab3M6nxHhr8ZqRtqMZgN81JtgpNYHuQEmFBS0l
dFL6QV0FYVqy2SVig0wqVxRa2ABtGo7Fz+7EX/mWElnKGKzKqyKCTei8w4f0z+mM
4KIoODi8RXyUpINv4KDE9d31pycn1mJ+vJdWM0L2nZoy1pXTDWIqeEzSiGv1kCiJ
zBVokC+fxrWXTHrj+p2XOe+8WCTbf/6Qe2sF1GjTAzBGXg1V+UZ8HcIO8ca4oBRJ
/b1aIoGUDEhC1yR8xK0dWtoAeAkr3Lrdv79IaXOKkfROX5SbcKMmFFEn70bmxoFR
AWM5fJvFSzmZOvMXKQ2EjJINBeYPIp1lGRw+5fhy97gRmYJ/wlUNLqCYsOyqZwro
ThHu5RvjrBgpsL8N/1uPc1o/pITyeWzI8ViV0cx1PYsBvbkQgMxCUbAjhxX8AB3F
Jb9olNbxt73JN+vpxpIjpMXG7I9UIfV+oxUPgS5pzj9lT65LROaj66nfV0feoWLZ
qrOevneT6NR5cZZLqm0Gmlql3/RnXDpJYfAEHb3549zMV769LesQ7l1FkgZXK1oS
RAkvYD+Qc5r7OdUIWmL1BlNW307ERtIOjASdv2FGMfRAMvar+y9X+ecA7pdlhpxB
l8209bKUjIuAGAL3YFDs9ZeWmR0aHonf24KCUfweUwmswhDFZKco8EMTge60gLfC
2JQvbaXwCJv2INW9X1X6UB7pYGgBgLFbGbMpMWRBR3qycOzezpW5rMqoYYbEEBXD
V3/WSQOHXc/y4dAK6jmtsfSaMLqu5pIlBGx+FjwpwWUox3ZDTJs4USzFKlJhajmC
MUeS+mHg4Zd+Rsqp00KOsgFUEwL3XmTV55drMKWO2s7PlV1Gwa5pPT7ePWwqHzj4
4WAHPTszobH/+hmnvbnwrMhY/XZw86ISqLnVC8kEzBFn6pWae1Z7UjHRAeKujUA7
+yn8EyfKjcLHCQKeWxxS8sRPuO1JVnSSwKGqNQiewOW68F1Ki+E6UWIa0dk4jqzh
hc8sxNtuFoX8YwmOdzlF6q8imGrVWNzbpAbkuYIxMejQSCyrwv0/KM66aDD0kHeC
wupj84Igj2YbNTZAZCt6P540g0u/Ds5AXFeys3FbZN5m+v5GERNrz7fCcYs9bawF
tAAzfJIVS3od5CVShvyNgsTuTkSFFSdSAR6p0aZ/zRuSd0FhxQ8GObJgPrTKjbMf
A/g9I106KDFNLXgpAbEvJDE34IVwMphgzwImN4Yw2oxvJBQVeMVIjfPKvMYwCVU+
RZ6406b1ufln2SzFgzXqsmxsHXiAi18iwnNnB3b0XV2LmD3ZdKQd1LA4TJ+9QJP4
VtGJwDZk7EKG98eU04N7kzhhfHofFLRGhwese00nfKj08/XuNUdMLmM2sXcyEDgE
PGfiV7Ifrq2yJQK1HPQca/cSGXCHkTRSL3sIXEMA80o/WNGDV+8uP1u5BGskh3SS
JIrTb275j1pJgtnhfU2HPZKfEoKkEO9/r/AFenILGVGBUta0z27dKfcF1ClrqOBH
cfzEF2AQL2DXRMFJKwGz/F9oKIHbx0K+Llkg+pmcr6ZrXQGkh5CA5Zytacw8IVEr
fnj+OIf+yrtSc7KQQ6HbanKufPOPz43tp43W06LDFszAWic1SYuWGFwbgJJnSbmf
VpbmWDkNbmdiqN617EkgHfXnCiS8AJ6QxU8F9IqyMv1tMDoQ6ksEQaiq03xcSvOv
f5hcXWp/6l6QtlImR3F6RzRV08W/Hib/BRrw9blDzXXBsrULuwRrId5ZJf5fOTHG
UBsk+slE9MUSWO4vrTHUyJ3lSfeV1cZawM8kCp8ybxf3O3+8PeD8EMBeR1wBnF58
Ux44Go+B2LXfJEkc82s6g7dibb0U000ACTk2dUaxODO+nXrBtayLDrTTnxfpTDXb
3B5SWwOi7u+eUoRAg6D/cE/pfwwyoaZA3JzC3wjsDuemyU88u2aRmg/c/m5yOdys
ZxbX9jud9QbPc/HIrfMluWXdZ/n7gOVZ7bCdm4P+AZ0uUf5y/nb162ShgLHIDc2C
kSE7R+I8ekjY7P5eml8kBquLhKE6fqxpt+H/fbPxZkakEx+hKGFYFz53tqAC/Vq2
9UFBDwjenhctMxABBSpuR9ZecyTUQ20p+IS/HPWY2t0hHjavxUeH+a/sbhgOTnf3
VOHmTKJiO9J14QqUk7EdAhVoRlPhDINjGxUSdDqnD9lU96+WnBl5e/hWXQwz7zmR
7PjuMpSdvkwM1yzINJBVr6JFON2t84wiTAR/uydB57wKJ5BiF8wFEG5q/7Tu0aJ2
sYqW5hH4bElGMZxKpUcJ/9ynSIzhg2aFcjtkwB8HkwWYvMmyunA+olc5PXLlb1Bv
ge2WHuXXz5q1zk2FOPOScZvGQ4X+8j77eHzm8lFKaOqgzb/0IebEJzSdwwwUpniX
WNFeuiVrXUbexGHm5rpGVM8JUBn6TsEHOX9YlB51HeR5RPRVfX9I0rZRU2/ozrpI
IivJ42FNHzNZvlRVtwp+rhq/+XrH346ZQQmbl52c/beT3rHYknhNu8Zb6hYQcMFQ
Xo3nhmcRZsncoYifWF35M9XHAxV0ofmrF1IfIeRGJT92NQ9UOfASACr2j5djTJR8
AFSOCCxtSRvwsVW/9H/Kj1XBAFqLCddQ/dfSDmf70QD5A9MS9DAY32NdSz97vshA
aJXzCmi+RT3LHOLlECdIn1QPeG36ruARoDDzyW7F8mpgDY5fwbTEzvCYpOMPPrYF
enGV3zs6zy+jQuFoH+L3z8v/9aL//6XV2qals4gsFnlqdKmGrNjFP4K0g0lGkDsd
CjG7E5GX5gkahx3VYCt7MnEIuVsq3LHstVitwTDpbR69oJ72XOnqUv1EVbx5UD+x
n1l2+4yoSHG9jXd9JEcA1tgM/hi8m8KPaPnSy6ddEWTZiONxY5NBTfJ5jABQFMaL
OgD3/Urknd4V4mrLrBRdytIUaDAWLol+C6NhbgO0sCtQtd1GsGcVawwO7FgBn0pe
6Osn2f9V1v5GRU+7QoG6i2VS+J6G0f0LGvdJAnDb7Yu7PAwo2dDUcR+K1hztMFUL
XabbAgjrrlSik2zw+1rPkgANR7Vpjvma4kkNgB6pWfe6RzDGf50P/i4q8e6sdy24
VeAGxU2ZkGGXQpeP9+I8w2pl1jEpVnfAUdZp+QDtOAbX66Zl5MGAr2aPxxrySdel
qiikMvYt/QbP3ZYSu/+teLritgWESZEDQyD/mWkKzjyGJk64JNG2V8g2rJdFhQ1a
UyQckG9RX4MkqFZ5+S570I6e4cnOFb265D/BVqvZTacfhuHvitXShCwLzXWvW2tC
kkmCgDSgroWQPNjODOTy1xLpvUDCFEpFpZvhTY9Tcx7KhhGGh9eiQTbJTHcvW504
fe71TWcwcWwMTVWAowR7HMQXLv8A7NvnUXiJduCDGDy3TfQGOqEz+HtmRZhb4D/v
xN4zIwmigCeq8I30PDGIBFwxfnOlO17IGpRq8uzkuRqZkHAg3Sx/mrrEfA7e6wKO
qEOGxMKisikslUI85oMVqiA9AA3xazlBOHfo50w93menXiBiK5jvwL/EnSy1yD+g
q4b58x00Gt6s6q6YqO80of5x86MjmvjcUgarT4SvHi0pwgSFRcOzDWkJBeVa0xtI
TFNoKHy+53xk5GWNFkkGa0wwNgYP13HnkbynCDsU/+1fHtjHiXa0L8373m9pp18Y
3wx0mrL2c3YcjL/m7J6FLEaPT9aEF6SXk78sArBFryEYQ6Y89Dab0ezCXNGyoIOH
OvZMSElos/VOH8c0FTEUHat2XJeERkMp26+DKVZ/XpGqx2H/ysWD9taiVwe5Agwe
Fom583S910Lyoz4EFum/v/jmqyfEqMVRjhZxWKfdH5HGcfBJ61r/+tpy+9ezLWa6
XBtwV66G9ZRAPqUnAEPzODa7uTR/0gPB8C5iNJRaM8vl+leiyuYhtK1HRiabAZ+S
QVLNFKHXudAJv+nTyUB0dJ97VvoWs5uE/Qg578HKlDDMDtiwNqsT6BbE0up+VqpT
FOTHej0A0H4zOMAMFdgzFMBO4frXF/tm5rPbX4f2uRTSK75yKONdE68IxHBSwLF7
/Z+cy8JvJWoP+KFQgHSIbkkBA5l294eh8f1JgBULSb0Viy8sTw4jBFla6k+iVX+o
K2+bTj4skokor5v1KaVQ8TUE8WNtJXcDQtqqzYVBC81yzqBUluLuc4McyfMAF0OG
pGeSNvZVLH/XzsP7raYe2chFgG5kvvrUN7YQ3hTdfU3s405Z+ugy/wOGOGM/IKyg
fZTgkV0ccRTzUtz/wPUbXzw8jBH/2ngMchKbCzwm50YUOx2gZcanHQe94mE0HQuX
DddFIT4Cig4+TXu+OTXZ6c9pxJhA2NBlma8jazNIXf13OSYHWGof1q9WbFI6IOwt
vSUcjmxVDIZnYBCJwP8JUF9rGSs3xhO5mtmvkjjDnPtmCQVF3DBLQMNQOlr7oFbE
/BsfVh1Jmi4n7l7ksGjGQraRJUlQyA2v/VOrVLB9h8RWb/FrpTOP4TpVj0FSX/Hh
1XGkcbTaEV1ROjrLmKySUjYdjWNbASOTB7V8JBgYe7nv4jvzw+ourIq3BRIhP51S
H7bPIR+mYGMttw5oUP1nZme2C41nOtrAuH5zXy0ZFl087mJa6bGDAxZVOth6/gDj
5rSK51KFZkcHSq4Ts9tPls/JKK7x8pomQI7xLOoorxDwBbJCup43GO/sMH1U9+E9
CDxlMnPWbQUQk6QwdYVUwwD3cwMm7pjsbS/qeTypI+iRYlwH+a3oPgdHOx/dZ9cE
VJV58XVamwwcP5auQwqIKK8rotSRM4ejgCjejspEu5TxNfMecXJAVNQASFgOQWgL
b6uRmhRCXb2FjHVg22wge+Kozy6WAwjSPcyhk4up7VrVvjvd4llNfgpWIALmcQXq
oNSa89TcfuL0cu5Bml0hqd6Tn2+NZ5KnK6uAHQGUsTAGZkTK2LlRWYDeMOHi5Vi1
YuPQNo1znqzVsX5FHo6LzfVtuhHF+GwkEkDGT+MzkVUXmeJ4HT1ycrHUmFkg6P3W
Pqn/TO75GbO6jvCumMgVwdUQQCi+JCBbvjde71sjccWaTlCSAzYJbc4nIqJFLpYN
/0yKsVr3rrfkhrM9/MHB8lIvSZ06wqPWRNhZcuJ5NHohyqu8VGUS8AN0+MpGXKC3
rsSymFDu9pcaka8BJvUb+wtrshorjCWLAoQxbvBQ4bxpDIw6Ib7mto0MoUMTt2Jp
jsuXZzDpupLtu2fmSb3f+uVF/Xha1iweaw2HDpn0JnhC4yPHZmc/hfruNinizgOH
AvHGmaUghvMjk0qaW/drczc554Jupwp8FaahV5+qQXBMNST7LI3r9GdNTEQyK3BG
dFIXjku9cSWu8eJQvseFl3odfpyuGFqHB8iRWl5GzFFWtKth8o+1e3nkLf8HcfkZ
ZP0QnTFMQgNoPaJg2E+jzS2M19LxnBvAXr75JepJIjFgPXx4Ji2zMq0iEk54GZ2l
4qbHmogwUHfpZfy6Zm5vyCFRsAFXF84pdokFX4vZye6MtShD9Lv6I/A/FYZsrU5n
BPsg38RIqdol+j8UwP3d6/q6uaXDgY71Gfk+F2J7UcZ1bPxwNDAFCbS7JSSwxP7f
f3mTLjwAS9iozeLb/7oRBqIIfE14Nx/+z2VgSgWHqQMwZK0ZG0UVIhfuGN6c3aiJ
2mt3cjUL9mYXd0W/nf1Hm+3IuwKRycS+RpqCaeoYvN4/p1j+fFJYmNrtvHSY3hQY
W+/r+0TYn7nm2StuEKNmIX3rlXYJ3BKdFFDwCSFZX5KgIHmqrG1V8dP0pZOaesOZ
iDxpZLDgzzGIQ5YBYcguiaqaQqzAfpwKXy20/SSzOzQwqIIBuzHpqlMYOeYCyUUh
tUCHDpKiA5GEhbl/xCdZmYy5IwQ637v/aaKXi5kByUBVbPqNYMIugSSzRYDgOgyJ
679GEylJlhnxqj/sJxZhElQu8qDZ4JXqfPSpisbN+BuVzbOpcH+M7LGep+0f31u4
IwIf9ciQij7GUaHPkPaGAu615W7n7eOlA/Oq37CLnkay3TRcNwrKBy/uiw3rr8t5
aj9MrsO397xA7T3bJLjQcrGiOPpSa6uQM47pxGQ0s0VmAxMt/ALVKKWKb9szOxYB
7jLp7fJjQEm9YzloNbJ0PRKHoubmxU7PbIKoPL8ed50+ZzosuYsQFGeHDSRdO46I
0amEuuhCbhoEBoa2ZcPRCPIPSprJ2GxOMTkRZHc7o89LH6kLAcycNM20JAmHXK+a
vGWSseYZFpvVj+TZ7CfdcTp8ilHlHn28NQs/VR0iZcFGkYiT/R7m09G8bykgkXyj
DRsc0fJZX+KReVAEXp0+VF0u/mpRGdxt5Qxy//9OgkfuIF2E+Fu/vXKGDd54eHEc
JTK2fH3xESTiHtXyonQ3DIDCMfdsAI2r7MrWnUCfqK2aRs+OQEX8y1Hwmy5DSUNm
SRqwnGieL9hscaJHPx3xf107QYo7J5Ze/99ZsgIZs+72f/5pZgEntwZCps77iOtA
cVEijpuJWGkc3pkO1ej6OYorZhAADvA7jF+PL3GjgD+CvYmgnNWqZHU6rQzHM0Ck
JUzlbv4D6mxVdKYEMiqkRQgHZPiLHRkpzsatIU1Q+j2HTeSqjvFKMwv0eIwmcuHv
j2sHec3OKW/441iX9JI5EMXSotW8Mzheu1rQqe8Rs34bz9T7pOH9aDnpc5ffU7nd
Nzej9JpT4aboMN5iiTn/SClhnClEzjWlK9hX3unuvUCDvZE72xWXy3tOo6O4iM4x
VEzpmABkc56azSpp6Utj5VXmlTkGTgRt0jPJ/omWAsn3GU+8o7AxmTXn8MNkEM1z
zXjPSu1tCx77R1lYA+EVscKbz1tZ5R8gTXpZA7f8D4zJVntukbVDbDB4PHYO05Wr
ZXKqpMp+VEBFPDqir1jcfBCDdA9dZ0x1AOFnMr1O2JeN/eGzlaGfpvilUVZr2HlF
tmktrBafmW0wMZ2tEZujmFACMA5rRT3qDeHVTDTLrgXaTtzz2UnmuPsgCu9P2iaE
NADlk2GPcMiqHB8Aj+CWncnLUBBAditkbSAnk/jWV9XwdHucCLbjc7SmOKD4vwaA
GeQk8BbML67pr1hjnccoBlKhh8H140zLZQpYhbGnVj3HlsDoypjekFwTfi3du5JR
lvD4V7PGecb5Q0uR2aSLHgsmkfZr2lOHtm8ixDG6+Hn0qcucuXqaeYu07Fj4h7Eo
SsjjrGvzDwFfYTYLopliPaweUQzQ18JsMJgq3WYv57lvRiq7xMtKtnjiqIuo5IGP
JFTpT6ysVyLUydt7rr0qiROHDAQYLsdjkJBJZVJW0SD4j3bdxhdOFjfz+JicKhIk
mf7P8rGi4mfShPNxurSh6uWYPZcU0uFNIcBYBN58aD8vOa6fzu/2hv8XabYV3Ky8
yYSpBqaw5gYrTWP66KPLYdbiCLL9OSliWX0H/nYI00YD9ea6Wl8fyfK8JMrd0k9p
RSgJ62ktP7ZQBX2nHdVkfosBQMAqp70BGiOjyVgs3/Q9NDH/CmAw6Sz+EXMLnVra
L6xTSJKAaLHrLsuJ2CarHViCfcRhbGUZKOh0wmNWJl+XuZ14tlKZq3q9/plZt6C7
ScIbAdGZe6iqIerXhGyvHxG52qKk3rovGS28f/IzrGVIwLu8RZpDtBjRiEawyZk5
xY+L08QSwHv+bdDMImYOt/v0Ax8oULs6/AreTQQaSYyfv0xUUSodR7ljY00gk2BJ
DS/k+i/7TUvx+0BJfa3Mmzo7zkNMZ2+6LuszeHU0IFPvFacpGVW42dD7v648Ucuo
6rFkluiDM6ACvzbP4IQQGU4TqgcXIOYaiWl3KDM6We5AwFYhvlihskkm955daHHI
p98YmJoShIzLHxfR3dzVThMpK/5MnyQQkJteusZHATqhTUKRsymHFPkexbPLRYdF
2CanJ5Q1el4XCdb+fyjV75cdzws9Epd06GDGlJgFUju3YG8ek6F5tdCIHf6Klnec
Kqp1YgKG7Legq4VddrbcS4cP5QutYAn9UzOl92vl3OqBZ0v+Uqpkj3l+Ew81MKlS
VzWs29VBIVMUIy314vkjB6W2W2uS6kRzDhDfgZdJ1r/sjmgWRAvunCPAu8SUFsDw
V2JtX/4uVz/FDOYHReakCl9KqmL5wp3cVc0T8wZ03sMxnWLgI26b0vatCLtKVOy5
PB0/JntIXHJ9Z60QNzKcJNzeN92BJHauBzeJLpRRQfyGVgL2kTJSmyYPxp2Org0I
7cBqHaR0GrtW6murCya1EN6Vun4aw+FdCu7ew/Ex/N7wy22CXeTLuFCkne05Miif
UhD8mqEXJgymEboNsbYHnuhB3pi7lNFFv88UEr+Sc1VVk8QsrvvIFmCvDqsYrrFF
OXYSVJcdLpMzB5TcTAbhDTVpSG5mEgO88XjCwcWr3TT0zA2Bg6hAfE6eteXrnfNj
tDE3EwLZ5TrnBvwwzGZzz3cgHHzy80K2Ntd9O9w8vKSI01zG6IWp2JLS+qTH7jTI
D8rFl7RmjOt9M79IUbJUu4ylbFcXQrcgEB6gHyFM4vifAzHJBFi5rC9R0+NF8Nhz
M4Pvtqc+Zyi3bvWBab7ArZ/vc619+EivWZQ+cIfIiBkJb0PaKL6nPt1dXCIm1+kV
jUQnh1qjqGgYPIco+2TJtD6koWFmVf0Znco1Wv5kfTcrMl8jMcYqKtKDu9qoq4fz
lF4oz4GdjNmYCLwvwXrIxbJ/3bJEF4jsUlcVTgs5rc3irGK8owBX4lRrQkBzirKL
R4LRWvDENZk19owFK2RMQ0Slcz1OFYjjBmrE+CqkNKnlkAsQo8cPMRLCPOg5iL2G
QbrFLQir24yJ7AZOMNXP9nKPwDVO/d9Cuwdv+LCZW5Waus3w+aL3NiZ2JNP+6E0I
zCeFUx+cYILj/RsTiKwhtD3A8EWOm0jZ+dEXF6iiPwaDi5i9a0039xga6YzGUYH/
szNQ89bxNvpVgrAxoy4u7Jlkqalx5PBimo87HgFApBSboWzYAz47VK71i94DPxHs
Z3DMBTF+Xg5476pIUSOskx5OcKbOC3cSwNhWl08VKk9HlGvgLG3e1S5qJHipjLKV
0Wo8dbGTFhtjv+snpWrxhs/LxtH/ANeyWJiZyMjPx+dx9d0NfkJYdlMfdnlxlsa0
hCMi995epKiBx4LKC99lLjPtjsKSrk2dGMeJuGCXBiCA2lmHr2TcGBntpDyTLr9K
h22tGr6DmhcR9OTN6PgZJ3l3X9hVV6p+fGw0FXqxtvdRRrubvQf498I59FjAJy7S
b3Lm1wm2ybHZuHFFK3+5GNZgqELH20g5igPdJZJM2E3Jkc6azmeHpMuzdGmcEY11
SAV/wgyvbdiITfbw0ODdnlScIvcVQfr9ZUnMiIw+4TqtLaEyjIvTfrLgPc3ZS15U
YT7QfOl/E+DbHOHhNK7rB5gNC6r2XAtH0ny9vzBxjPXRdFxdWLUB7Hcb2t40wNEI
FahUJfoq3Uqq3XVM9F+rDtqFk2UbgwFNCdGNvv+YrU5RRdY0XULCejH9M3XmvbdI
gk0+P3Fps9GePBXTDGUWWXymGhDfSb4IOfVnlvrgFQ8aiWshIQIuzQCNszZeKGMO
2gULTaRD1UfCLirzOURH+a+gZnXjPEVXanDrpzDfZPJFCxGmX5k08zsPKD3qRHLL
bNe3OfLfU9cUXiNAahxC6+r6Rl5qIuTh1tqZ5sdvWDryoopEw/gCcQnl42EtZxlC
wi0H2J8dx/bDPfC0n8TVcmvthPrTceKhLY47RSBuBdBslpwMuNw4mzy5a1633zWz
Vk4cE/viSoSF7A9KTxCDU/9oG7UnLaNsN3N5nOBh/qfqx9VFC43HLztHvtOhfI7X
NqvfSeiectpqqw5SxDcpa0YYNdHFwiRCpQWOwBPHqqZXn4oM5CjJGpeVrF8lfl3M
`protect end_protected