`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5408 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
OyGGrfLtuV/iB6oXYN0vYG1Tpb2FcbJuf9mPuaaFmHkKhAMaX1+ptqw1A6pSdQLq
pdwyHOmG1vsHlXrnmYkrpMSPmd1PU+G+ONt7NAmhk7UCD20NdyLndKbYzaLRaA+K
UvzW0eHRDVXx8u7TYQ5/ggYvX7Za3r08caEp+QD7sxmswF601aNK+D/hiutseC89
i2iEzRm3EjqZY5kCNkTSwIpRs2mkGIr1fBtsiLfbDKI0DRo91BCQEofqxKwihTH0
7uM1QYU9iZHFzKBH3ZwYZf/g0tmy3Qkqxi/13PCEGJAl76PXNlHampfUHlu0hKA5
mzXECwjSRoEEJROJXm39xitcB7UA+O/r0HKJtw/MEMb7oPAiC0tXV62dv7cyoU7E
BN0wUWuk/UKkt2vXjN+w6QLHpJTgLKn/ml/8eKggKw/lRu/cEmIQ7RaXepnOfRYU
rlFI15AkgM6Gh4is2KT/d5o11vi0+9SYqoDyJXw5jb/yeoxagTsda0XNHo/f1s8m
HWlvZfpzLKbFm869a8UGmZaqeh6uIZtXeBI7coYlig1SzoBbtwWtmbYXmQDYqhrC
TONuwvrobY+Ud7cEyg+rZTB0odpQtn8xBcnDEeP0eROiBIa0pI1Z0fMJ+OcvxVIA
9IBJuUa3ysRGNMew8YdDq81qSe7DErsiyNFDZgmqBCYAleFC5MGdHE6qs70j6c3s
8u36Tiv2XV81rnkqaKxKzYbnVLbiMvWBuKSBzQhaDxx7HnmwZjQvge7Q82hF2Rme
DWhyGK9CaiKCOZY1+p5xX9W2NG1PH5mKozhBP2nja5ZSpvNROS99wS9fgt+hYPtg
bkLH77OUIc1Enl2myH5rw5vk2jmADVf1gCgJHefcw+LIh0GaKRvOrJMtxkI4TGbv
S1G1ucDV0CUoM4/dvnKAyRYj/g+t8ceCNNXCjo5KH0hHuQxm4cfr0jHtcryN+Trp
/N5Xf7fYa8fuOdMXj1qaWkl73Q2rpu9ReXMPBWtVv3y/LLEBrTVM///lASC/5d/u
bH16UhghtJNzRsTrZRhLt6RRh7d5oA/xgrFhE1w3Ej721fX5WnAM0SwNzykzA4W0
9TMJ9JY940+06KPIp8+sap24eTtI5l6/+s8gRO4b/uyCVbTRkRT0+G4Mukf+q/F3
rLUkzHRnXB9lYP33QPToPPUamGIZtx6YktZaIDiYjmpBLSiRrtj3zN41FzZcM+kw
V71k+Vz/stvDo4YG28IuNy5fym4HfheHYnM2muflIDxJRegpvkRLaGWuRcUWypDE
6K6kTpp1pav6ST7U9/Bes/ItVYJb88pGNxlMx2AJmP8FAai1SPzhapOTTrIBXTo4
TxZX3T7MA+piraTf4nrL/T1hDJ0r8YAXN7Hlg82BPzU4wWspBjOcngPYX+b4zubr
H9pmC7SXn2vNv/l1Bp8Aahy150i7YOTbgyQkej0EIWf3mGapuJMfvcYGfUZ8j4T0
eQslU88Q/Oe3/knO9/BZTk8TUegXVdFaqg4xr7qDVCoQZpfB41zggC/cOQ0kRpOc
GnFeQfzlu3kXMAtz5deeed0i6+MDugXnK5sTOS7Qwvh11BbKBihVaXNCZOQAYy2n
In8ZK4zuXgeGLXYTEb3aAe3bneLvJerkVFqQpFdeX7NDC4hE3dkGsqoduhxWuyCe
9O6GYN/CLOZuC9sUirSwS406nbBdjpTXo/f+RcqsHpeX/aiKZHbz+5qnBOPD9B//
rCz4WnSPNogg1rl4MGVd818jxLAtgqMcP7FV8cT5GlQ1UGmFTrWwHYw6fF0yrYfw
C8nYpJ/l1ZdwJBdYYjvAj556L5xkPtkU6Cg6JvTeFt2whY8uf997zDrWzTOvb+sf
0A0v7PknmXAHgu0PRZn8xbHvl9Tnzc8qDFGOGnHtnW+j4updTC2l7PdPlMJdKZjI
bdZisbTYAJ7qAX/v28xWnRlomNudb0IbUGhfm2CWJUPgkaJLmYqeyLcYUXL41rAU
uqo6K00N/XZWr9nv9v2uBBVumNRi31qU6FTGzKXZJvsBzFjxeTTS/AtjBZ1Gvf+x
SE2ni4KqJ/NIiPKS/MQvlKQ5RpDZdb7Bl9j+D1ZY/IX9RLQvKI4ddKDlJ1uRtXMG
cgG024xMCbWeydBcZbaBWeg/q/LZ+53Ma/TqAq9FMzvfjTcj4HZ16tUtMRgquTqh
zjvOURFtiOeXwGtfpNBCyG8tz0Lm0YL86XHnAoapFGFc1UTqj3KCRuW9kMrp5QGg
EGaB5iqPhQxE17C8pJZMgH7qyeDMgpTM8yV1N2o1ab2r4W0BKY/Uj9oLFB0aXtiP
p+Qa3yalmxbOdgyXkcFnp3/S5lM1xgL90/dFh11nd6SaRvJKxfVtNju5mx11SWmn
YNDqS2KjlVoGgtlCvM/KkfZzfK0wmiVMH90hCXlBmFULIW94QpZaqkRIBByXxcXq
vmSXiWiYZc+lD0s5X18kAaIhEIFug6VTDqPyYLFasUf7ySw5yZKmuIHyf+C0q39Z
mu5HUVa409G6ffqPaqHkKxrmvS9a85xnvojl2MQbGoVCABvyoySKYZv5E2w2xoCt
UB7IRvuV3xEuYYielgELfeGnCPjIFv/4xBtJjew0uB3gw2BFVkjXtMs5eigCYemf
z4b+9O9ZvJ2HMLgtXlYPB2YXlXAOl0W70GTwZZyhO90ApTIJd0i3+wQ/+u8bUfCO
K4Wur/c3JHjCPpY1GngmDsRxoM8lMkk37T0Hafp9ZrnUUu5VDRGqU9kOUVTn9HOv
7hCLeozK0GaYLKlrlICalqrN7PamWuCQiGuBqmSWX1sXEXbo+S2oWRMdUNkpOrYg
VQ4es2lW+pA6eXD7Ww8XIq/f5t18bQgJOk7B/r1OsqieqNiznY3dlMq4Pt5czvzg
6aLxa2lhNj1rh8CaTdTH8a8zqNMgWxb92+rsQLcd9fdaIOQ/qd72eiNqEAzve+P5
WdZco/zjK8SRkqeY1OrAnd9KGsTdfUiIAPbviRx0fRTOEOcU7cd3FUknHmeNSMd/
UOLBGQ3SuI/gsGE7T5M5y/u1vf6nuDtAvrP/dm7BCXZcJKwMJUBzSJ8qLJNkmhG6
AllfgoH9IlSL4SUJQKsJhFPbStYVPaODlW0i3SuNpB8uXKMhE9I8sQgJF7/VzsxF
O5enNwAuv0hRDk4vOW0RudsJDawLu8iXXuqLlbrlUP+ofjFG7LUXdeQjH8IAoEKg
xnXObb5ogVoaGBr0LQsJ8ysoqLW8589H6kOOQ6dzvvi06DbdiHZlO0Fh8XhalzIR
CYmgA96OZpwGoTVZJcP7n/rm6xjX4z9+pQ3sDm7AZhyzg12TZ1467ICCR1Br+Uhy
d5LCNeLOe0MIKBfuViuTQ0j1BTqDu5ahOzq4OO1peZJjgKCa5tnryjAufDWW0jO2
/gyV/JqlBj69tqYnBftMurVBm7nPS+bOK22L5WvEnFiVNz4M+CA6nZOihgj4jm/c
SHz76puGPWPNmwSB/IbBzG2gjtf8Zie0SD6xf3JXZUISOC6uZHCIjPUGnf77efoD
zPrVrXMnHReWkTBK+qTe1MjiKIpZj4vMbJTfHGV2hEXjPKgnNnbqJu/RqJJgTObX
WD7pwTB3Pr1rvMk0mRlnwBytsdjyoZAkmQJpEWRwE53jQ19u4S01rWgOdqveajch
8+yonPQ9/vtq6vDcPqhhQ+Pdzjd/NzszEn7NxTIsUamORExHpG+BrQ/kAt/+1+jl
Rcff9TsiBezgvmxUpxis35+47Pmb3LH5jLHdSEAqd/WiWnDIkWbwIBJMYRVzduOI
w8xwNNYU3iU+a0gdSd+ja+j0uHQcHKjJEwU24yT8Lj8r+Gz/uQsFKgsQ0ki+Bjmx
cTzS9M96bMyUD3KNq85useZpF+6QbIhoipCcyPMflZCHlryyHbLbprI+IrAIy+7i
SGMXiukCE89N9LUiWqPUukFHtJZvDEFz0CHjjNyvvTUvKtbUaAw1a4hEhd8dyyGR
cJ8z5dNI0gF1HxldiOr49+0uy+0BHQr9xh0sSNXt8HwAgVscUPS6aQx0wWUhQJSu
SQCHPJkhnZH43KjoWWPvmX+CKCyLwiopc2XOU/aIYZGJB/Y3BUU/W3F1lJXZfcNX
cid5BbTlZ7MIIzmdQy2mmX1YKX9cXJyLJv6npxvn5K5qCCgJ5UHQX3x6dvm9IP3t
zzD/6ehhR6OhQcP5/n25Oc1aDX4KLIW3il+Qx8+BSSGEOndxtArXxhiWCS858WUw
8dXTgnZXfRe6pxhGUtEx8qOfXZ56Gj7nUWUTj2lr4dZ0AaGgKOs6Q1eA6boNXypf
GAkRzfkhBRjXRVIi/EXBdblHvrJdaPksaZkBZuJ4cdnCCFIfJ0UOkZ5f1wr38VOB
MAVGv+9qz4R36v3Fy2LNX2IkoeBbw1A0v2tZaU/bqwWRtbHk7RGgwPYKFK7W19Ap
ZBBMVdf6/Wc3IlMalc0tRbrubS9H8za4+GEMgzXrV3Peyn1uY1S32y6zZTZDWBV5
vv9MhaIR6OtrFnRK/k+xb4G1/84b7LazNYSQfewJFg7moSM8oNxIsRPkP8DMbTXv
9mnx0kYCLJ4XKKgAHScW5UDcFlK/FcpHNYF1PU6J+BuX7jdVmLbB8mwnzG2rpXZ4
zkmGwRyaGaP+3BEI1N3YyPpjtRP1sJ9c9+BRynZugG8/EXUW7pLTSCc1VV13+EFg
vVi7fOkdf/ro4p7KA6UpICOY5Y+PiiGXGvUkxO3JoIihw3hk1pnglNcyEyyg/kI2
5ZJYcu2qdQs2kjsVF3jnn7vI7KX9wjb3QEK7YG7x3vWSp3Ar+mV0mF+Q5M2g27c/
mY2s1PD0oROJxg7hYTkYUq3azBPzckombPp//jTF/AVgquB8jEvub/bcNn1JmJHX
gMvht9Ah/YXxH7oAE/R8eGaH6RVGEn44gaWitwwonC8vkfV/fdq8nYnTyh3ul8vm
ybuW7/KDMAQX+bO5UIgSlcrC0pKpt7PW0sxpwH6vaBIS6hbQuo2LBwSdzrJeqz1e
6wYfg5fT5tDul7CExWhhCcYwifgdse6LBe37fcaPlESt/PLH86LSyhtpmKvfPkPL
lh3//L/PlERZCOxnliNKW/bOJEdWZCB7terjXQSwwAfijcZg1vA44x3IXgW0dQnF
R9oqBiaPGrUKcoLj1OQnbB2BbnX5LtZ5QhTiKbh6Qhgoq6hH7I8qcCD/xD5MoY8I
H2qg2f2BVuof5t/40bvArC715iCtIAnPnFHfUuMZwGf1M9fS/ZS368Ra85/FAO9q
emvBy2QJBOYHSmcVSzlAiw5SdaChliXsOwQIv0UcQhbkesrsMahumRdgQAajDXW5
hh3awOC/Vpw692K7brOpnlfC8z3wdV/lco6tIams1qgnpqTRTFnE4vTH2b9AKhUZ
OucqLLbGNisAHsqHKbxdc+S59oGSWkORa0qkCFE79ndUUGRlbXt8sxyBH6a9q1jU
rekSgSwgb4uiKH6hYwTabI0THz/paitg3S7MZvLVMxQPtxKwTuODS7B0Kbhazb8v
rHMI3sU2GQTkCFT1ZzWv1DFOOK2bDxtmLgJGRPYxg4FMIogXoKBI4Dmam0nnNxBt
Bq5FrYKX0tBa9OWIDkIcZI0DdCMI4L7KgxpsEBlTRBKP51MJjpcc9UlrSn3jDFfu
l6uszDt59ecSANxdWj0X53oZuzKullXGSwAObcy2uUxILYZoyPBQnJ1ANcoZKmzK
9BrMWOBoPba8Wg1lS9Ls3aXulynXPhXGbib8ohrzpUWZqOJsj52R0KZvkZhaHMTK
P+G19hEwOhYorEYJ6LRI/0tnbBBdcpkS5qmDCIVgM6aOBbqdeVyjQU2k84guz8u3
tz8XigYGXpsNnnmda+dLiW1YC6FJtUcCfxKGcEzQeHQL82S07nQr+4mCi8oFzYAJ
XY9c60Y7ZcD41IkkNPCYbFOzlvZ99Hlo8o6C3xiBjuM4glRZZdT18+8Pf3hdnm8I
86IALs+nMiB6GZ9PXbMPKzrwR99McwW6RMeUtZXs9gBUt0f8Bkbu/hQ85E8G4iL3
A8JBxfs+1yssJXnZY8jH1SxaX06YMfr9b6YxQbeDP5clKi+EcW5zg+LoJeHjf3tW
mApYJS9oaKxmDDfiT3aqDZajWJwwCZ6RozmVTVgG9PZAcoX4XpdMA3wedYgi7Y64
w8yzIAiQ2Vza0N9ofGjgW2E/m11d8hT/foHY1Mx0BwV59/bzIJwuHk9edai3sPJE
7kOuR5Urw8nDlADyusAQboFC3E+fY+G+ijQ6R89D//Q80FaqQeYwfwfgtifP9JCF
ADWZiPbLxjAB1wrry0p2JW9y8T4jaUP2cevsO3jIGINrGOAqB40u6pmPEqp/utYf
rTx7Q9Cd8n4NetMKNyzodccrUz0KuFFljG96DMaren2ZkvqpDpTM9/KXv3SirtPt
SOBZgiViTWAiWIpsN017Hu6jFpWDL7VcMzTipXwT9c7vuHQYSpQHTGLLl9RlT/Wd
SBpcAWPLLpSPHfugPoj2tLuuY1JJM7/r6BvYsZSpalsHqsMnImjwfGElj5E/2Hq2
Xu63wLOVwdihKd9aVV0ibldAH9t89/lwrL4+ucDMttel108+Fvh8pNqV+Ka7ipUX
6BvOoNFlmAFXJ0+CDkQH8kkIIa2fHOJP5iolMYrDqpUrNjDASEOmiap/aPeSzLKv
7dwCP865qjtz5ryzPXpAHpq3D6V2+DWAdJ1s6rsP1WwEEUjCtEKKxnD8ZO0a1+Yf
0F2VwAnh0Mw7OHoPntviLH4SMGcapJWTKsytVDGD5od6O2Pdn9DbjEaZkSXhcBGw
Z5ZH63AMxqYrtOrNyTVlkto/vhZ/AdFbAz+qTlU/mo6SjLVrhbJnpxTfe2rb7C1M
hZ4Vgx5QZ8CRDZwJBHkaDG5pIKMo5XfugYVH2J1PTUY2C4YL5jDfcqeJ0TvR33lT
ebuKKTZlO6hi0Fz1Flae8JqQU5zQ/nPoKa20DcCxHMzJ6kGzCCdmN3CzdSg6Dw6d
A/OBBUPIQW2IiFZekgFblgkdG6jTyFneaqxJ3ZuXfG42IZmqgLBx0kERSvFS4rSL
s2zF4sehGYZgLnxKpVoTNlPFycpRzdwGmR1+M66wZ30=
`protect end_protected