`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10128 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
ZIICkMu+S2rq/yOQyqhpukXuDUJ3ozoHBU3zo44aVFEZvI8EnK6I6DtLeXG7z/gf
OD74d+8HoG9U6+f/TCHuvSIsAvfiKokNXHGLkC3VInuIz4eZgamGL4P5yuwGXuE1
pSWSOtU6v84OJ7e+udMSU1h3KfuxeWQCOPEw5JCrTuO3+I18gnQzjsEzzeCmVnhx
mj9JCh/wdF95Jxel80kT/u81L01DwZUE1TA6MSeGRedv6f0kTZmOUuA4bDWBFWa/
I+bgvTPSwp+DhcIOJ4tPgzWqIAPIgKVlqEZIEiL4jELbjoa1v/QDLn4Rypdjyott
CouOgzNcnRfb+bX8vIeYNNtMiXCF15445bfMLXUOxVpoFoqenzaTFEn2xI8gdo5N
kVrZ+KeEK2ARGuLguAAXjFm1cpTcjkSOefuQQHsfIaxx6S0/K0qtO5WtZNdZ0I8O
LAbrmGQZbZZ43xxpqppdtsAPdNsyiTtaWzIabKhoCLhQV5pSIg2aUH9LVWwqomUq
bwvBGNATzliUG0Txi1gjxrGEKBRND8Y4rTxi63W/iklKRhsqRelgYfRPCEPFw2KK
N8Yuncnqy1PiG2ZBmO3VvGBr3IhH/7EKtf2yLx2NBDT/pQJsaVoTH6AxQ6ar6Ubw
APWbty4+PtaDhhRxfC+JqNaRCIPuHfyYXbDOZq6K8B52NDeurk2Lx6xjfExc6HSK
IOUIXNQ1nsL5ag89DrMeBybBzGQiakYhpAXGLntaXuADveYTV4ZwI11pcQlU5rEF
JsbSoI+8OvGSBqzFxnghnolGnVmOEiRTAs8emrQu5elGn7Kt9K3D3K33kewSAA1Z
JfA/7kAArNsV0g53WeQsfzZcMcPmziGKw/GwbACPL9i6U8Bvwndwem3Y8u0sJiiF
Fzib67UzZB/EA8z/eDjlLJKicApwXb124O0OS0zNY2+jX1rQ/PuZJpwrc2CXCutc
nzJLM/rijYIqdGewLQudZ5zt/Gnlo8jmaBTOh9SDV/V3zM0csuhQ46pKQhvhUL/4
ZdC4jmonc0tiL4Y3kx6NcduLR6/4EwL7puveQ9Y+AsdVivI2WLwivoFSByAJu+6H
pbWYw33gZxbVKI+uc6mzVwJDE9Zh31xun+GJiGs2D0ehIYdiyP0H9sPWQZCHZWq7
rRN0Cr9x3StUi+lKfohD8IKlHoM9e78Zj0QyWaNExCEMlYCPDuUBg2faATYrQ/tQ
xNB+7A70sR9TGG98syt8nkVdouFt1czG38j69QzH6satVZ+69cw5OIRxkOkWqMLW
5LckeSKcsBgtnzwWuUR1E5IxWxI0/6AODBWXpYdMyminjp4DwAn9lQG9emRwlH5I
6oICflZv3LvEYjMBx80B2+h1ZGpjNgVF9aBxegbCGAoRIXbE74Q7+Kr1mWYziNTS
t3W0jJP7JA9jjO3wO6e/6wjTMu96Dzq0UEiQe+g0f3MFW82r+siYDzOPkoUy0MtZ
z7G0griWhFkIL4GXMJtvvpoMBvTfSREZCeDF59VODCAhSKi28cQq4QYV8I9UYPgv
LC3hApNlT+MYj5A3BQWqtjKHZ4jG1IlqCP1uIGPxut4xzI7sichYea00hoTIPn8k
yxaHVe+kYGxuAICKzHglCczB1tLdhBCINJOQlh+sAjbAz9RnUEP57TKgni+FXg1U
gIMgryWUcNAJzWNk69xAAkvAauqyDh7gzztKSvIH2Lfx+Rz0VONCPtFFBxbslr3S
Zy0Vn/jNGwb7995AFDHPU8N2mLnLBvW9XG87jfMmRqZtVX4OjVXw+tFLTHeEokVg
XPtwTs+2srPxHGhYL7Ju3U5t160dSjRI1WTSxv4m/7D5jOLQK6tUUC2GQIgrX3JF
ZFN8Wdv8qe4orrByR5arbeFBCW01QRMMYAUsj1v0UP6owQ3Gt5PUTea7OWLOubJC
jDAwtGto2zZPPOzxhqlZTgRK4v3pCEp7gmPH+2k3c6wrlhHNLMpbdD1sXyBfL/9T
Y9w8oDnSJHvKaTNHN7fVnJCzLBoCnq97Pa1hRLBxVnltfW0dCaTd9JImReaZfNk6
5qrsAuhEPPstukBNXBRjJSNVMLOW1UKn+fqS6KzdokAfMMdCd9xakWT90ERl25Gj
ORC4mE2iw215lpSLNjxRbSKppYptS7coLEbqz1npgRFo03MBeV3L8f2EmcrpAWe6
qfvW8XJC03Jii0pegXrPKdmye0JIsV5SrLXSoOtWxSCzN5aT4vxNBEQbjWZ0BVNC
Wig2CBS929/PDrna8/q2hJVGKwjPUil6S0mMDQcLeAL+nQO8usZQvSLy15mG6R/V
bDkFje9/bkk53sP9GXmyFwEdySylz4vwmmGSCadzNBTsTwI9jVqZD54hJy1mow5e
5ZVsDLxXwAmeQ5Axscd1qmV0N2LBDqkLDygATlOR/ebCIAVevZ0H0CRo6yXk/k+1
mnPbI8C1BnuBgX+EWcrItmebJirkTvGhR2o6ngLIpLHEI22D2CvVDVV1GoMv52/Q
OMjNcXirAvoEVfVp4fzjFdGsJCDw6WZ1WajoUC3t0k0QlCHV3eWwLtbjvUS7/Tvl
MbCPHACb+8ecxhqSkYVz4Hrtcsq/8CPDJJ/Bl14P/FuANj8AbxhXCBjxPrt0L55I
WpPOZwXf7bgovCekAv4Fmmzi1oZjKodtJt+q19MK87ea2mT3Q7LJ/OXVLsBp4zpQ
PrVU9L+fr0Y6Fk8PqX7WPiUTnfJI4SRdx18FhuZz5n9x+Jpb8LSJNRHEgXYFEL/B
nxRdF3hjK9zoOXY32t8UkiDQzD2GCmY8w+Gh2P41Fezpoga/Lduvf2H6cM+bE57y
YiV6QWuF6pmT0BYLz7S9pJSv5+73gSdgZ7jg2gEMzqcMd7/ZefRIhl+fLGdITlqq
rinmo4QFSLWVwMDR45Tq6sAv5PGj/tG/yJ9v9odJxtIwrhM+rmKCxy7P6kqzuDge
+f44iT9pPaW4N5xbTEz1Pb7a8aGT5JBx0RPucNOIBG8SBSTkOzJhZAFudEd9fUXn
7UaUtiwvRhcD3eu88DE+E7ixYLK+XFHcB6jVt3jZ/MammhBHJbZu6jnO+v4ad2xf
HuFBQr8QAW4PV0yCevocx+mqKiT/qUXrFCOFGkWtKaG1Nl+Q3O9lMN7C8mbAVJBg
0Q3F6t7rRNZoCHGuQNcOCbe94AD5vJp+8bJtwp32xEARDl3pscA3WlUqILowv1/w
X8gCoIyItl0wPsKPODfJ2xtU+WCLiWufG8P04jq2BYdIGYhElyC+OtIW4ygJeJNZ
gKtEvw1bF/lmbFZuW8kHv2AuLRD1ycfgivhFjCQAlJYOjg8fcq6gCc6omxF2QeDB
Bq9wIcJCc5hPHCXuoeePRuzc65yEyZikJE6FidsOO1jHIcthWFC1kBq/E12G2rYb
D4yLv3ddnM0od/3jFOKk0YLzbH+PbUr2i6bbsM7dz9gg8oL29WBGx8VfVRBXajRw
w4AoBnCtSDR5hRUaTMaLHKIphsDKvfTRlDzmjDghzHRUKrCkujqFEJjhNO7+U/N9
3tYvpu0s04VStRM1BNaOdFll2TjR1gOSlF0hB/WEAMbrWZz6E19mrVr/Jp0g2L3N
vZPiG7bVjaz7LVHCYJPs0TB5E0emtRx8A0sPbK5tI5zAimdgFY8kXJDWlKIK3Tsg
ZQjBDpkl+BkhyRMiC8SiHomMv8QGHjgHcGC8XF96zyhSNfZHmF/oFNXdV8D9QI6q
B5OX/6/YkfU+DaZG3+XDCWDHZNcM8k23S6Z/cRSwqwk98no7PIEJQrVnFFVergps
s/GEOMICquVQ+8co4Ebu3OIDfRyEyEUbynAuC0kuZIf8NcQ8LWstZhYPErP+qEw2
TqgC+9RSf9Sybs7I7YSWBAr5RV3V0g3g9gpBxf7jXjR5Mf8Isu+cVmNxzWX+rxt0
BFV7yqFTfhrQiTjUPVfi9xO28lLhISEnnb3As+i2+JorWQ45LhBdvFze5g5zIead
DvhHDXjdsiVxie/eqp8GSTaNq1cVrB8NxHe2q2QFf+kch6eHs5VKMzGgJ5I3wYA4
lV9lVWmpZI7NG1IOglzGFDFLrJRetKeqvPFnuD8sxtZYcZ6S2O2MEOPaj0BXTfeD
XezOMte/crOgoxkHWfvxAG/KvlW72rFZECxEXqS1RfARFdAJQKsoMNADVh/W8fx4
hDzgqHEe3dVN/JHm0k4eMjX2aXdRMGasOggo0BE69ggveAn24OtDHB5zuXoDtOqe
5OgJAl0TY03SX2v1TJIHKYmMknd8BOcWQ/niYkANw+wBf5X2533BdBYOiiwGb0AI
CsP+Q+VvkmcAAqafAhF6lzZc5qpnyAA5hg2tU9b/1tC5CuCEUqJCJbkKFRF0NiNR
pNP/glGwjg5p65QPCvHC9tTW2UwBjwrtim0+3n1TZRFNCWZG9HQ6LL8ZkO2lAwXD
fJZN/qVuP84k4PdN38bbo5rNkgj7qZVRXMLcTvV2PRNZLQRFP8Xfs77NKQFwl5ub
cILU5PAO16EmlNdXMscuCyjCNalDUuBi8Up/abqMbvytvojYy0XIC4cO1/KhH0Pk
nPBa8/FDxrR1KVxm01kt3uRimb4xAbrDyxZz8x10v5N7shaH07pHDDtHFyfokQXc
zqpa6iFyXUhgi9DDAjHiyh0FxmKYUVcGSltbQ4RazF0JS51uXOp17XEmQGcD8X8s
shYUOMnbOUI5Zx0CJ1zdeEHTwnw1L8ijNp1JAbziMVOEGNrC7gvuuakY9p2KArse
QY+DJEh0GgcmOdRRcOMQ7KwTDes/VRHL8rrNVBWFI6+o6Z0Y6ZDc1tyO7ZhjrXV8
A/S1hc5lFH+Gs1NDlXcIOCebUhBi01eVG1KNfKbyjkJSlylXrw0P8LU0xyPVfejQ
Wr/xv05J/82TFfKL/LLWOPHp4Br9CtItrowVidDHwW/5R1ipcjx5PFo3yOiW/1GV
Mr7iivi652tp2OfPg8yw44WDR7/E7nn6NTpoYhOtJibmiM/k9URDJ1tGHsLeZ3We
ia63NzVCFYrxvDeURoniEYkaRGdr8g9zgAWwYZoUh0jAnkgGOlAnnz7phEX76yAk
jEyh25fJuBVZdlX4fDvA0NisWBvQb2mgUQ5Md+I2qfJjgTTkEM7DWxzMf10RPzmM
une4uy3nhuu5c2wWG9VcFmJTB44MmjwNjvl1Sm9ZxbX8mZKv4TimKXKItNrBHazW
M63fApA8x/f+jt9GVziV3LhohAQwf/qb3sIX3B2FXYFnS6T1eyL/s2OtT6/UNsSr
3fmWvtbw/uSESZJjRns7mIxWb+4ZNYtmNsutd1i6Kn8OXNEL10TcWJesWgf4PBwv
iD5VmwfrmqgiD5+9siGpRu1UvbgZQaQ3ul5uoO4gARLDrrjnuy8603BQko2Ghsn2
mPcGHp1QTDwsMK5Kmgn2QAugnmb65/DM/YTs8q4gSRvIdAseKbv+Y8CfKHijOAW1
jrQFJI4YljwBhNoQs1QIfrUZb2/OpeBzFhY3lDrMlWKYdbxblntdekRYHCQ3A60B
Sxk0UabEtUjKplF4b4bxCmwquJs24qy50QLf0IcYjtLUfKB9gQAVzs+mHhgDiMmZ
mhg52Rz6iZhP9LVdFNzF76lA+O9Bi5irtGiSDd4QBCqjKlfF3MpdD4pUdykxXJwj
OP29dNGkam5b6H4gqRJTr3CsL0M1cDwxMPmAscunPPYsP6FyUHkofx0nRCKX9Qys
RAdQHGhlQiogMX54mDsTthZ/IpjDihQv8p7og9LzMAKR42JjTYnxZrnwAhCS2zbT
vvsWlSALfyzSHT8WpJ4HJofDX0Rdthzg8C29NzgPaLcZzirS6jk3nTqjD8YwsGqc
VCh9zi5iZslHdtoFLnYDyUb3RYFPHXw7JV2RguT/p4QI4seALukrc1WDO/asBnMv
LawU7vu+r4R5p4E+EgtM4T8PDZwFncy8YDhkFbMaXc2cGar0nMJnIZHj8AWLM0+t
vONi8xJ0ocVWsPRzvgZS/VRTbgFBOouQHKwGt1f5Pe6aRSpMJQpaMBEyQCJXEwkn
Zb8TMffBqBWPQMxzO0L3gK9NWeyAeHR06tweg2a48oVSBkvpzhkJfUV8IzKBrsUL
cMmst4dCPcWSqFQyW0uSJhKPNDT/HRJduY2F+EV5mUXO1Sl9+bAnrgS2iWyuN5o+
Qg8osanWFlv3MoXcnXlhn5adfIb/jmyjhExwVQZt5v/cVILXQm8CsjZhzA6ULyft
R1J1BhYq7Vxpnae9uauEDck5nco73dRcHDVF1yCk1pEKiPTHfYuQ83FjI36sBSd2
2sucJHiM0BGLPxv+mpw6+3+R6BkSeGttpdnuU+fXbUnoRfRxs1vWyG6kY1BaODbs
0TqMi4f1nUe+atLBPcW17/njft2oR9Fnyj0h2nyGMBV4J5yo4lx/AYgSZSZDZEXQ
qV0a8qiBSZtcS6EzK6E9wW0d0vu+ueO0EnmIRBV4v24tibs5nQJNWv1ecCnv0rM8
jkIgsUleI4cK0CcMvVC/oZ0veubVXUxRjHoWFVdwwx8y0ZWDnypKlxL3I9qDxc4o
f4jfUAI85np3l4zaopUNuIhwexx2zafsSt5Q5JrFHCRnK6wPRAttIIxvVOXPJwTm
a3T6YoQDLlNaxQRxZ5IH9enuzppiZLW80PUE9WgLKQ5AyT0KMvl03iYsWyYpsP45
I7VYHYClvcddbXxKGeOANGxmGa0pOGJjTE5hBzG9xY6Kas6zFP0ZSLC5t9KNHiHL
rBS6j58Q4p2lI8PyGOIEq/Taa69E2+T9v9T9AQFvm0cK+d7b7WLopVYnpQg6AcpG
A8vYRbFIj/pZqvxItgJYCjGCN8YU5mk/Mj8vMbLLQJp21RDb3ON+2QEGrHheFQjl
23kT2fH51Ksq2OhQw7NJvXqKI1rdY/LA0YBW/U/a7iNrvIvQKHQt4XxmMZv/233M
aB+5XeHn8Ld3U7RzZhF29x+Zxxg55CpYc4n2jdj0Y8fWL6Ftr/aWXcJisbif5huB
2ccApvXYQDoq1hGEWAqeRPGtV4rnAy0wq05FAcJ4cRx1txcAU6RuL176FeNVzbk5
gU6CEy7e+CmDUb1ve1yBjK5bi9LdPWgirdw8wPSnXE7kU1QSXLa8gTJkkETCRrJS
hQsw2qWbobP2VAy66avgrFVK/oJMbQGojfOozH5WR20eZ7tqBAbByj1hWAsAbuOC
Gh77b1Y5o3futL9vM4uEd9WL38rX655qcf9NL3C7E9Wr6kIUY2ZyeaG8PJP8mmm8
n/bQzkMA8Ln8a9NOYH7i+lO4K48UExXIbO+MyMNRygJx9ZnwiQQEXbu0L8ikDG2J
kkGlgcaGscEqwLH0Dlz92dxrlmFeDHN3rc0vezsnLePFG+aqxYO7oWfRSXw1kiaj
6yJC3L4SKQ2iDbnd6miCRyvcFwfLjkngvejemntQJYzYojVC4vQPwtB6g0NGavaq
PuZjY77YT278KuZ0ea20OXCQIAtHr9jhBBfixx/+ribGbyIW0J6kJq59EPUvPJaJ
8890iZfmDQWBi92gSNrWYE7rZNzWru0qMFKugDSXDt0UEQGHeWip2w/PSWU9l7bt
m1HEaVkwnQe6BuVZ3ABUOGq9y0qDQ/z3YtuWC9A8lGhdrYLaam8CECAaoSdHuCrE
fWciR0yfU/GMQxbg+x1M6vIOZ5GEeasRYn6bw7jUnR3Z4NmM5wW+5B4X7l39p1+8
4lTC06+m8PNpfr87A5qi9Ihfs2b/H4c+UXkSF4Fp0V0q4UvniZfg7bbHGv+8/Gtc
oHIXhC+udwpObP4zuRIvmt5VsUEkhN0HPnwYdfDC+Rs8VuvcllCpvbYm9k6ZE9gp
wCZBuvJk91pgcxijO3BtglJsmtpt+gpkHt1pqJnK7M9WFt3zwykLe4Mt6IbLgfay
OpZo0EgMwx7mhN1FJMw0HhN72RleIkKlo3fTvInzPITpVqnCVoONQQaPoNLpVdFY
1jRPOkfRkSJH9/1ZGFUYnLP+NUI4K8imkmS4Pgs2FzT4rHWMYM4h/u6QW/FroKAQ
LDN5miowg90XWQRXDA6Hd6V1bJVG5j376CT2IPGEFupyK7TAcBrEp+dTluipSv/N
iAwiDInS3I10IJjjqmL1WtbGcBOzRdVB8eBGEsdUMO70F0AgAtO879RgEDmIx6NS
CjO+8kpPjwZIZRIJUhRS0aJ3dw2zwc8lg8CwCWOuHP3hwNpsaFHtud6gIFEILFFH
lrShYS/8Pu5kieBMNrU4v3dXTlrG9brLTl8ccflIdUezBB3nL4+zUYKwN5YLviz7
KI4sYth4xh6tvEdgqNiKJKSZOPSzaah6sQ2mkvebO0rA0lYCG9A0d9jkgQ6OhzBG
F3xQEtcvUPSp/LyUVpL0G7v1KUXNnkx1Cr3Zj9YFwtHNo+1CDdfjzAx/9JBBIYvw
J2WPe0CuiFNcxREPT4ux5FPgRwRYwnQxBtIGp/CO1wZu+n60jemZ2B84er6/MjAE
JKnQX0sMFPrpIe3kqMe7dE5en9m180Ida//YJuN88GfAvXtsdaXMXkoT5ceMl7xs
7HCQk5aDQgVV3hP/G66SEbG/UtphHD8y0E13vi7G2EUAw8VJG7fbewmP97rNJMQP
0o6nDmBbLhDfEQY0CjNYiqxjld5fTjAikJhKkVAWYVTfSq6JvXv+eJX+E2jSAokk
oyQ5fZEbruv2CnLI72FEX28q9cIhMzDwZGYMazweNB+W1xJjmXaap78Z2dU5I5K7
hiaHe23MQw/xSkZqQDV7SnHvEh4I50FfpZHW9Cp5qLgQR7yzeWngkzOtUOsqy8Sw
t5X6WuHk2S02ipyxTLoOlfpTLNEuBFi3gUSgKc9itWJf8nShjFUac71U5NLsKAzQ
wL1xOzEkeIyx2wsZBY3gmJsGCxQlBeRhyVhHuqLFB+o8e5MsL/U7kjsrjw8zLrqI
Hsml5+j8M712ciEXp67d2BC1hnjUwIPPh9SHM+n+pjTFeo7NYLbM0u8+8XpA5Jq9
j4a5einSFeuQNo8H8O+hXeRZaCJObTzhZ1OD3UYZ+0KV0dWH+5PewZjC1j6CTTOH
hlIBAvbJwCwd1W795dTO6UYMJHhnMrp16kZNI64Hzjd5X/sqC78fqHeq/VQNVrcZ
sR7EY7RyqjPeTIFh7xmDvuMzLi3aQ3V0XouJh/Xi3+dJYN5zipF62KnUwvXb/6HX
Am5sqX1H7Rwn+W8z7arO+OeICBBlYR5c4mOLYdK9Ez6B+Cn8xziZGYh08GAkNJDR
lWJfcLsd0DNpwcySu8lUyl1D3HgFKfNdxVpTggl30G5kdP5ZKeWNEtVuzIHQlj1a
G2/KMtfEJMn0eBoHg0sPsPRaNmkVP9MBTxmySz7mcTc1ZM5RB3EZsIda8oOTSRsk
bWYgQorSjc5K4C7IaREAKK+HmjVAlQTGdqfrqHVPiC/HvImTAIlXuxEu5iSh2eoo
LnNBPa5TK0DT/OTRPJBYvXyLmQ79//akphlXKfJwpt00SWfCAw5ZGPQ/DxpNERqz
AR9QSecaj9XaZj7szQ7tS4Pfur05iv8kxlqPsGU54niwD9+cIQFYsdn5mK4C3Zo3
U9eetR973CqytVsr4DLfU0d3GkKSjERXkZfLbLCyRbMEnUJR34X02/S/u38b3Fao
67tvgjCewE5a8bEp52aeaodzqjwNfHRDxRu0BzogR8mbikKX/GZiiDoWWIaMeE7l
5aWkPBmhUYlo7EOGp3TVDD9wQE7LQNqbUa2SOKw2uIQP+y0mtDsLUb2Gg98zxSpX
0nOpHaTXVEVsU3kA9ot0CMU/luogBnqIB5JythkdDxL6aFFwsZhPeU5R2k/0wnen
cllN9y3EP4BCuVft9GVVo3bs1MTEfQYii7K8oQcsLvvhl7jwn9BpmyyzJqhA1wtH
t2TJylJ26i/nwdkaMpkZ/c75c5XNQyDjs226XWs8lqdd7n5p2915jzm8sqyfHXOl
8TY95mf0zAVrWTHCwKBsUWFPwXOmKHdprZqWdYn/ydZt6nm8Ygph26sfGPJwirfu
fr73mA8VbgBaLS7p8aZvRpjoNATvR+xdN2rHfbG59e7uLyunnRqE11PXPLuJLQ/0
HhZLhS7Wa2m0UAEeJ48DAB6R3TnbwTU5ZRNWWi5a36FF7dtsTOCZpQNyZ0qSyoPm
ZGPAhP7g9xmJfrXLHqFSuIv4DyzFpsnxxs0vh0eMoe6+MuwaHGmpmbqSucbk27Vw
mwtqcSw4k7o65hc6cdX0mGtpCjZYRkRdR57w54qSXQOv73rwHmD7nwkWCL/raol4
sB9ZN2bcvgB/iIFmO8tKv8f5UKfXzTf/YmuCvLPKo5AAW8XqN+Uua2WuoaLyD23e
XPZeHVZq89qHYgsF+gypVM3c/cWqKqz8quJg8rr4FUfTLbJP8BDdPuopFd0KYjYK
JY3wGFsowCEw/Os7JSQxX7d5EWMyj5pCt0/bkrPpZFhfqcbN3Hl96279cu/U8Igh
JmeFdS+Rc9RxGCYJvzDNdMtIYpjrEce48CCKizi3FQ+efdoeAHm6XZmIjZQUUvL1
WTqkvb+yYfIwRd33dmcaGrW7XSy/HBIOA0s8NNKYtfZIWEBqVI4YohDJCBqRJ+v7
A8hCzMiTdWG2g2jyVV9ckoyR4FsoHwVxfUGlcgTFB1YK/bqBqXZXhNkZps7Bb6eC
MaHJbRi75t+W3AO5p2sQoDBAJscy9j0pJy4XjXkjni3qNXLtj7YRDrb7HOqYbG+m
gcNx+MeDKwe7gKRr0cIQ2eKue11SR6m3gJqRG87hcdoiqKXF18EaKNzJsmbiKKBN
7lNKGzwVQmidtot0Ug34cdCUqsIfxKBHAkegO94HJtspXecOZ8BJB2LzrgyJynNi
da9eGlwM43z04JBrKKXHXSt3DojYLKHaI5ennfBJTY0ZEEXFJwcakKxBWA5iGZTl
6qZbb0NIY4XLb1UQz7Q313sGMnGor06YsSKwNCMnK/cjBwHO4SQD5Rd8F/Wx4gDI
5EJ4r1bd2zV9nNt84ftfC50YP476n3neQyv/5cTmznDmlvS6wtDEOjtm/ZabWzzF
x+dgLspVRmsm6m0YBEVAYVl+NUyK0/9ohRqFZwTbfIUAvcH+qdP8eIrJy4J5Z67b
QroKsOYwkCZOt+dAsypZOhLAgBuBxK7scA3HkP3TsiD1i4CSuo639FR3ztC15Mui
MYeOT2mw5pQvv68eQjUaZYWr7Lgsf2eW0kv6stM52EsMXxTxCq7NzxRfxAZyZSy1
keIFLy8ojP51NEQ81VWgeyPZnplK/gTWcfFmJe8P+3n081WrLhnFQiUF9/yPlBpQ
77nYzmdNXW9LwfwtYZMR9dP77aaPcX1jd8U3ZJrhilDFnA2RLb42ypIQsSUJ9Px5
dMISJp3R6zliR4jlSLzi9cN/NSZ5dnmttDJMDLY8B89TSqSC/lfPSgXOeIRV+Rd+
mNLTojjk35NVdU0MTejwM7zc0vCZTbrU3OG3ghTk0KKp5lmfYiJJf8xwLhvejZfb
mqzE65gdAqtK2NSj7YNE1GvmgFTFszOdSDmK2I+mxvEKtQqMxaOJmaH81I8pAbo+
6JB0AqLKTgmHSBSvwzDE/3Tpncwlt1pGbD5esn1b+OXwqrU32GLaSIRKW+9ICE1h
hXwP6GNzF9nzFrYBACXvobHXWw18Zn4k6isR+UvOZOt6Aez2A9VeEYbToDsbTbFh
v7CrvtR2uY7DSiL2TzOygaQrGB+UVzuSlJUxWZzV0UvPu/jQw8QmwLoS3Hi5xJtI
wArUYLdA7CKpPTz5YFwwSgoVyWpoYkeSd61hcivRKadvM6MOpeHVjgxZiZz/+x26
lpdn3qXW4OMApUDboAFXUZOeuJp+ihpro0Q/kO7mp8WvaHZVKG2nuAtdQUcPtL+7
87kfkoxqCvrMUM0kDEzOg/XssL6Wy1hmTh2EaAXwlUfzCOdfnfajMQ7Ud+oUEIIA
BOaaLI1rvUKnlDrCixzgv9K/3fHz17lDp4qTrisaK5fNKxW0JZPQMNxZN5QH8OAG
vmED6BjNVRdYDhFoLjN+YQgB7eGWsltSxKJdCxWK1ICdL5hjp2yNgefCV9LpulW+
pZaHX8P62LyK8redylXhU4+5DcqdsTDL/PT7anDI/SpxqSX13ylPsXEpKe+m+joS
l9PPbCISQqJP//2+pXMiex4rzi8NXYVsGhlaJQR4iGDvzVnFDd/57kWIegJNFT23
RM1hnidPsDOseD9XIKvXzegkArOtZtXdZb7FmhpgbxV84/ucKUOGNNbpCRjjLzxm
1KTHXImJyOtGFOXMqaYEseyhGkcR31bizn6skqQ2+MDJtDU8qTShdDgLXaLf2hbK
HaENbbl4Paj+x27LIHJc4F6Az7YJtkmU0HMwvAw/rAbAgDlXi2P29DYMLcMij/HT
shbZY3np/tiZhU79aooTLJ+D4vlz6qqCkLv1BPOO65dfEA/KNas8sYiPdgVc6J2J
AoLZLL7pxRWRT2Ghz9AXStoThZrzban/t9+3BVFORc3FcT5Np+oTDS2u4NnBlnnv
Rp0GjNZAZGPLJStAD3Ed6lTp0imVe53b3WPsnG+7BNYPNbGa8L+p/qCVav6hmLn6
nATJKMI9kckQSSH6SBXOirDJJhZBzSV//76mfymK2T+aqmlJkXMtVq86mzBdTNqp
Ute8lnPnAcLtMaCYW2l3vK1f0hkiKVxVPoQuQJVtX9M71yNJu4xiKkQ4pahrahBZ
PlvwtPFXS9+LgaRNfql1N860wVbbwm5phVlL8J4pY52B4f5W7dbv9ozAI+UsIV/z
B3P8vlZfHnlJ0aK2IeygtNfyv0xGQSEliv5kyt3e+TWDcT1qaUrBk8lz30Wd5iOf
OoD/SfWuSEI14nZFvC+qMA3P7VG2ZCMMFNi+0VvYfX9OCIvw3EmtbCIvD3fpkmKl
4cSLGJVC9ZKRGnVZOFoq48dRCtqOB9fDKkGM4A3wTH+tahCz6p5GZlzdXRFdmJWv
P4/G17zwhbz8Ba97tsCe7CA5GaYvQKYZNPL/ZPXqPzpVcoLMYG+8e65IzxgT6s1A
2veTfovh5G/Ms5d5QrP8VVO+Wyo1f73Iqkrf8dDXIH7ykdgSgbg+OMt/oU1KdFgj
2BKQJda8ScYuOj5YqYxpyxgKaujAnVM1Yts1mgqtDw12vaQchrlfONxYYNDazbsU
ukLBUY8JCPHArg+3m89n4+TqkGk0rqR6Ce8zjrWOKCzAHt8jppQtF/Q8PzamQrIw
pxJHrZ3WMaNBMRPIH7rUo1VdvyRo+Bvvni5F/mbmYR5EDlKJtidvlRp66wzybMLS
LFxI5IEBXQJu1Zgzj/eZQjMrqV0sIUBFDUhyLT5d/DznkIQ0cbSYFzFspQr4XLBJ
Tdm33BK18MFM/zn9JE6ybSOd78bI5mKnXFa7TFLmC4Gp/JEiUIwPWvPVqNUti9Gw
`protect end_protected