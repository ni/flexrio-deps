`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5744 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
FTGcP7VlpSOhasofAJvqcFdPmmCzpJH0pPSlg4bqDJjaFpICHlApvOnh6lJaRAlm
IWmtfVIjrykrihgo79y2lJdoP/voQsAua/juTm+fnesGXMObPk64OZ3iRheKAll6
y8C0dGynFoIn/k+/11HU5AQ3Sr7BTbTCqFpbkwZSRipSYreDcvlTpF2xNMP5OtOO
CK3VTnSse+Y/YzMuXRZIztifkMbi6Jprlx4hvFvw+1R0LEMdsUaKslWkOBdUzEtj
ETRNKaMdMtVOrNiUAE/X4BUKUhG46lQhchzPoGpfRx1xF8D410Lacz/aNXQiw2NL
6+ZkYfvQLBbeHATJik+oteSCnJ7RynzgB3BLB1QwXIfkl/SsyvxjuagRUrQpzbfS
eoZz1CG2Qf7NaT1r2aWhnNcZBux01PoSo6GmggTTnxS9KmLJakLTGLSczp0jkbJf
PrfcxuOFjtuyiJU6cf2ThOyy4yqLu+NWx84pLvi/Maeb+GFUUql3g1Ggk9DLlU/C
7WdbIdBJ7Se9Qy5aca/a0ygb3GLUett7FlArNET2tRfi0vWscTj6x2hSl5APJJIo
HcVcLhS4k7hwfBHM73skkV9w8ivV5EjL11p+SgxadOlGymg9F02nznKLvUElAnNc
QUPSExfDOk0vv1GpODeJFYS/EPU7YfUtR4Krove60Rv106WRmn/Ygnqo3iMYAd5s
ODqt3eGG2sfppKVgImOuiYyKQKsDuKglZluAIThoBdUTZZk5T0h53lqt0+gQFROV
tbfDhMOGgKgy7tP6zWiwTtEtLWq6svbKEVXOmNxPVb+ALOKiKSsRPv6kmRnq63qY
WTkdZ+uVtoFTWiXFUxi4sQH2JfMnRt9prlB31WBjb9JgEYC6IdwU9wgaUO6f01F4
ZqOOwPUep6EcdF7ZDDh9Ep25gQqIYju6L24JCRJEY6KLuhJ8hkZQDt2BZSu1h7JU
HBKCO+r9bQ52/VFTSvcaB5y4PT11kSF8TDSB6JmFQ+TkqACjScwCLofoKAC+9Ivk
FAR8kA5b5GBOdIMLoblR1V8xGXYANxzQGyM+erhRfgUe9ehGym1GS29ALtqwOMZN
qtITdi+K4z6PGUQ8BksF1+wuRLZ9UxvMfUDBg1fLEA+dKtImRRyYMr6I9xkb4WBt
a38ywD9uSvTa+cqgwz5gxoy9BG+xXeeCPDcjwuCKnLXfXCY0ZhqpJOZmiLFAMh33
ALN9GYqhXezfTyuuMKofLyU1H8/Oi+mBOhkWjmHkIxJQXpxgVRRC/IRi0T9XE1jY
1OAS/rhX1oct0BX8Jod6uJDxbR/7ubHoTVSAqW+ZaZKnFYu2UUQ9TgLyXv3WpKtH
WBshfPZ0Lyom5742QP5Xma69aSVs2OWl257RgK5cqt9jEOzm61Y8tf9bcSByzhgC
41GH/3Zw5fbzs9GArt1cwm7QWNGtTMGlfPtCGDjV1AWFxo0SFevnayfvGlb723Sh
LnEvVcHa7clcYygoIC4M3nEjqKiWy2BYU6C89xpwTUt1Rlj6n4j2Pz5AZAXgteYV
aD9A6cRzWI5OIY05gj7cCO6Iek0bAeA9tyZzShBW7RjII335dHWm2HHLjYU9U7MP
9PeSX9OqdFmNGO9u/5zcTnhwECLqzwJpqOYp23feKLobb8zVj3cSLIdRgXjZGv+G
LpWlKF9cFXGXvisBJb1M41L8DyGXR1F0dZP8c/nLbG6MGEVaFEbLOXOGOiExap5k
o0PbD1COne7lp9oV5eiUooNtBTECTMkRK6gyfazpyvwIiOCB/E6KDZADClit9L70
7AYrdwZuInUEa/ZPi2elaYfd8+lBZBjWNpF/gFkLr17NvhFnLI2qC4U0iJ5cevUd
29Qomcp7A+EexS9lS9qR0xTDY5/VMIMe39ECjcqTAdG0fQassFJclMmi67C5nz8b
x1fd8bh/gURC9oX00fu8vMrYCRHjyHczmSTCxlj7rFjL7cL3WipJ/dAxn5UaVutj
GSS43Pbel3YmbgAZxx1/nrDUm4KmLVt8pgP8uCzupjNIGlgqkwLv3ba0lhyW7802
ueZFLn61aMi6USdN9M7dQMtE54MbwQ1voRCEVIR3BhIWjqIaJ7ZUniwq5CgcO0T7
E+/LWxjJctMXlfhLS9gVC70QgSE8W5E5SgxojT5n4UNvtypqk1Gn2dTyDQDpxITl
Dku+PkI6YrwKt+h/2jGN48/58O+CPuHx8Omsdh/AN4J+WrDPTj6IbPCfLXL92V8C
gfMdFepOazqvay9F9SeABfmDcDHeHbFLCNvV4pQiTfN8Neo1m2+ZZvZKBCTQDpmD
vtMqiReF/WIXOVGEmyxOC2Xi46DPAFp5+uA4GbLzoNKEu89M/CHT2878kL809BMM
MPMNlH3PxZ2Xo2ADNiQpYRAbvrEGCkS19AAbJEsHnXn7RscOr76rp+IXFvLLpqeX
jwZswwIG/bGGfT1mMzd1uWvlHF/fwaZXjEVhs6fE8YJfjO9rev5VRbuyI9xo5Hx/
ajHfUDPkzvngwHKgqm128/OCtMPuuenf1U8hqAAkZMF7mgrcYAJRLyjOvG50Acdh
nCb7xIJPmdgZMre8IV0T4EbkOO0D80Y9sqdrXYzZJSmpgykKf3dTCUv1NVmFXHPQ
X74RozYaNalFC906LO7fkiOcOe4VBz/3ZgYzld39boZEGTUQhmlq565ZPHe/IQAt
zI1EQb5hqPd988Ul5gqH7V0Koxa6ZBRUn98Oh7vny6DD/TQLI7H/aLUo6suYQtEy
jEUWszMJGZ5k4nJ5a1eUnssN4abnGT0wq4sm8OV3tJya0rPtMjohxzKdkfmcfT4Z
RQL6KE+pSJ3ZvNN+8kcgWJuldR9CqjpHtZkngMFLF8pkXn6L/BlAV6hMMlpQ/rFH
jasHtu0+Hz0rXYH7RDQHI8oI+GA1xo4UezSAX4TeLE/iUvikJRiC52Xmvk6dFS3V
1N2tVWHmfZiQcKKjtAyzh1TNtlRs9QCnWGMN1bDAyPzJIyzE0oCT8PevvD1TQOf3
PjmwUZUgdVoF7Bpx8/woir2Nc/S9BKvuuj+/UXx/j/+z1QKNzR84ImnahEECBovM
2sgrYNcUQVaGD+zSn5zKbQMhVSTxaIK89Ujy/Xr77XXckdDI/wSxGCazi2PsxORU
gm8eAEYNeei3j1ACO9QqFZrdcwmvMIISbcPRywgetoKT5AtorbRsyGx7lzKMnYbs
lJmnBDqifz3v0uxMFGHLHYUlhNWBJv14rWqSlKB26q22K9QNHrRocJC8NcyLnVWi
mo8MuY6zJq2V+Qm9tp1nGRBP5WGI4bW6WPBnOWhgtF1+RtgZ1Idnx5lJkYPT2tFk
DfMfYp54bBsC7qiyuaeKI2yDJMVHlPsNRnVjAuuOUoh/8iaJWXhncmdSjFWNZhO+
iRQmyPl3jjWICdmgOw0WOFAoWHYNoyE/WOQtCBzTBuqI/7AUMT2DNbT25k4gAADd
svVTYtHwwFVuioFHrHQ/hs9alvHuHlV2nU3DrdadVZPStngNqpUIVeVWC4416/R8
pan6vc/ExlBd3G/BNsdxf97LLrCKffmBws/RMbAYvF6IJQainapqy5mombSIBsMZ
KpYfD6SfxAl74RQ7p5Q0fvwDh4HnUXJmtbLZq80Hn+PhzdHeoO5ULuT3e8UC532D
xuaT+mor8Xjaqtzcpz5lMmgWaevo+F2WDjFAJkcBcvu5Y6PyBs9ygXwy6i/+iT+0
p/RP9+QM5jt6WzPT0ril2CDN79LGxhYf3/KKJmqfYVeE544IKfPQTs33Rf0off0Q
/ySyRu8ZLIkO0AzHrBZ5YtZ6TZ4NpQnlHsq6xmO3nm0ReAHkIViyxtGna6/vCpjA
eJZGOUFSKsVRIz7YzctMRfHtrm8k5Jko294Q/9F3AAfcy4f9MBpK1WyHZPFrA1EI
smVZkdmeG/e3jU7ZwE3yi1EUtBM5NydWSEimfUMe8jIOFCpCwak8M6ZBzIkv+mmC
zlZAi9h+hBh3qQ+kzIbT5khPtE7IyOH3eA9x8BBSy+v2/rhnMPr1W2Ajqr3NYoIP
4CQRElV/mKu69tFJI+jQCaUFvjNGn3Blpru2CvvwODS7wrkkFCNq0NGk43ShnYer
mxOm4L4iLEanWluSVVxYt2IHSf/IN6oxZGTvTgWWC6nwcvs7Xi0uwv+uyYSGLBUz
zIa1qNtPJSoVNwVYTmuI2kKNgMjzKFfNNsVor0vEjUoZp/vSaPiXgccB2tZmnnuk
mu1W2P9QVDK6jYKGRwttLy3HfXO/J7YdIw04M6hWWO73rZzXX7NlR/HdgeQ5siiu
Ci4SpAmgpKUY5q8BITeZwJhOcRUPZhycPW7W/DP7uJkTWUyyjGLdzSgSpu+Q6VZD
2WCTXR3YOtAcChLWLZRzJh7Nq7cXXymVoLNihZg0cgLqpIAhaD+9Gfu84+OSLttu
J0vySxGoKjnz+clkiPjayUDfErUOUz6ygByQgMUgbHGJPOTIlLRzByudopjulkL8
4jdi7Q4Lk7LSbmiBmkzDftIte+QzODdjm8RTeYS5Xf+PuF891c08w6caVEG2jP8M
0dmEOAuKLauvCSpLcd+7VueyzVwbVKxYCNlLUoxKoaCTKnbkqveV5b0c1W/Dj926
OAUu2RnUdBtn3f2y/JJ933pbEUC14a3jdAN99zDRe+3ajhe6dptZhY3Pf26eZfoi
quT8gGtI6fG1OE8YyyRQLp4B4NcIfK2/OCuHXmJxaAtq2hI3rk50eU2m2DdPe3ok
CwMICcz1abu0njWAjXp9ASTIi84bFggUdpVodSKE1KRmJdLSlygaYDrXhYeRZAkm
rHTLznfqQazR9UjYJmWaPjFW6XxkqUDReWXHr1c51tjA2UOya+Y/7RMVYzFr/Xg3
xrfkPHyWLOynX7d2cM+FpmUTA/0l/MWCnJsgVH0AUSzkn7DO8TIjGF08Y/4XNhXv
5dcBwSJCM+kQveQPVmNerDb0omqdo01X+HPe3GpX2VI2VqHbFqncEwDK4WCZubYc
I3er7XgJE7D9iMEKcgfwyW0k5dcVxAor0hJCEsOupsktEgriwl+vIQC6sJUXrZa5
YReKSTyYxtUGtXo6rbg8wSReBwWvK3zytsEjVoGuz7Po6E6Mq4QUn0kfB4EBoVqY
Ipgie+nIU9jdfw2k/9zZPSd9EJ7NZdlmeFJrcea5WIgas/jWizkvPmIkFWkxibCv
0mf6n7vAHS4DfUPwGgeNFMONJURLwJPNgu4ZncykVxDp4zKLKXvkcqnjdH8NlO5z
LeRV37mSw8cMbtHO+rlSLiGEaroYo9bIH8/Dsw1juzGxDEjtY7yu3xXvTHWzEzdw
HxXJYpTzyG/PQ6KT0ZJsyDPfxpysVLVr2IjnSI8E6GdUu8fISDzllia+rPBdgL3/
3O2vN9PbMuoLnv3SatldDeAJxQFnp3i20anc8UoqfRUselicLDgfwMIynmXAZ2bK
R0tS1CXioffxHjDmgYzWb1hRvC3AvIIp4A7V7rIsGEOGmlnK1mHzDupDb4qLWfvI
tfwsdoIMvqNOcM3rC+MWUwzPcudtfUkjCNT/8lGC63UolRzKYZ4GC5Z5pDbb1Z9F
eNVNCixVshoVxAynNxvn959R0kKC2UafjJq6ie0RyHooVl/lHIkJKHmZSgISA1W8
b5GwLNjFHjxkbhFCzbAZPkR7GecNae/FLwZAKTXMYsY8D2YI8SZXpEx3B4Me/97R
BzkO9sFQfCJwdjYc/6xzkWTvwhtNARaxi2AnQjE/yok3+Gtn7VyHHTMApGUf3OQl
9BVUjf203rVyAShZjaVH9FI3SaQ8zsTq9VvzF9bI2CYgXARqkxubu/aneb9F1/0C
n0EIasBI4WSAO+fiJDOqlPA83v2HdLqxUYBiy6G/4wqXfmuBfc/8dEr2ORpoHQt5
U6nW8JWP6JsAN4bsdMdD7wEPGbQchvpxPlrpAkALqa02qz7Vditl8RtbosGoVz2p
TA3z3rvYRW5sekHnZ6N6qouRwWb/zNmmQpLJ88TudDWyniuF6kVUvcNR1efJ1m82
CtBNu4jFRSrela0PqoZ2mfOPienQ9MFIN7kyDBnHscS5+5/3jg4pPiwbdILw8vfp
ywsI0Np7A1ykAkQmKsTTi+KgkvAVyhSys9YNwbLIeDaW8yGmIBwy/9PgnvLTTOY+
wFIxTzPbEn+9wXznXW40aGUiqzBJL67YXDhBFGZ+40upMb5oIbXL/zcGJjY6KLmP
07kkx1KlbibAyzPlFE7ZM30KVOdHm34cE/qKalRDLdd108IhR3hzgcx1KRghFgV8
c31fQzNCUH3Y2EsPYCFBO5JxErRNJc/EYrF4UCy7T7pykISqpwkMssKnJbjGosPJ
G8PP1Meka/sa4fxsDeknpP1S3ft/cuDQ6qqtzdFlSZ7HFc9ghmBg0nrBio7sHjPa
2ffQVjyKHyopTYfuZR0AQOM5E2V7EH6AiiD4Y7jJNxRpa4JbQLu6vd6+nTGrVNx3
BJvT+7atSD+XMbuBM8zy8QqbR0mdvT7P7GpjA3q/J/+1PnDasLKbzzrAGSN1ESkb
uuFDTolUZ78U8Yv5GzHHTrvDMSfoiGWGMfJMuZKf3pOw3g0EJ/aQdVjEzq83/0bz
HtVA60UCcgaVgLz058RSQ+nLiHXMfbCVsn55m7su0oF0rpLa6+YwyBujITpwHjGS
zwZXB8CsS7IOWHPfSD4RIC7uLnYVv9epvkg3wE3vZ0vQWQlD/LEBlWyxZwdoXd4n
Kbc4lA2yoze/E+e+qPPJetHZPLg/7ktUgzmAw4lWxrs+pJwttGmoGNm+COIN8SVl
wU8doStgN7NewGEqfgem443abk9bUEi9rh30MZg441YERbktPtCZsMdSClLVSSMg
FiMtml/Fpz40PgzZzl5jlnJuPD9qYVPYOckK1Np0gm3FxfABbv7lVVMOz3Ufboef
TJ8euDjn7g1SgGoUeGjfllK/X/Yl/JjEjwvr+Phh3XIEecgRfUkHEn9X4hWGpLGc
MmksOf1E5qWPKKi+c8PvtvAMr0PtSLdRnZ5d+7slRWvJqHswMuFJTCaM8jxelGcq
fNAVIEJetDQK+XR0yjBfnKFiOr0HXvask2Q7R+J92h57dsH2n4/+GcKdq0YABVI2
ucWgmWFpXwIDB4Kpqe8OdT4VU51cDoF3J6SDYreJa/ndnUpe7XOkXIDUN+rXYYf+
4FEDPllriAmIryZwcU3F7ZaAokwG23xAXyuf7n+9FG1P4HH2nMGxE6vDhWs/0QiJ
7UB0Br/iwaH4zA5xbKITxrogpcdLjNQS41J5suZ758JUaGvEyhIuKM9Zti9XR6IM
N91ZTmfftRxn26uxLAYuad5nPwAxpu0f9cNIAfTqKRKLAxWJ1hHGkuvT6AMUSGVw
XrocEb5u4bWhMcFDmf9pbBq6dbNhuVBINx2ariR8QfzNISp0SQKT2hkDizXXHL1e
EZVUsaw8z6HA+f4wePFb6m2NLUOosGiOetm1bkhSOq5zA7kaSPiWSDleKEo4qyWT
idhYGFIe1YcJxAGOMyKdRt0MnPVUUVfsMBHL7Hsm80M=
`protect end_protected