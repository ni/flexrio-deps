`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 16560 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRpcw2zQDHRgJxPf7yaQH79KEtnTCle2MtJU8K/kQpZKH
fI8TvDYlaRaoZ14z44xXz6ci2rrSUqmvS/467lGm4zRRVvlA7F7l9itNQXGa+vO6
mnO/oSbTbTCAXI3avEwDaVujOhOY/CC2MYEG4axSht7g0qfL6Xr8KZvik21YzDAG
pqh3g2yidzfwN0PXAcBv05ROYHlNqP1iH8ju5RR0tc9BOJsESgvGS9H5H7tU9aLZ
KHf2t3OSH6hGhZDwtnFEh2v2zlQwlajfbUGIyfOlQJe6s3AuZPEBNF1WFFLloRKe
+Eb29jPuC3SiEgaPaW2mEiPjv6LmN5DtyF9x8s9263eMC0US2bHRwtFEX2GWiVEx
SQpxMeIaRVYXPQIf67ay1vOez2QrpVg88/0xOYQ8pRyvDFDONE71aPgt0mSjk9lB
2mQzmUXGZ96kRRlnuxrsPOtO9IMX0OVupUWWavHSUlXVMvflyLXWx6GVJl2sqgg0
dNqaUccimsLnazlYwgIYXbDBw+gwLMZ6+AAfPL2hKmiFrl9OkKMH+4V1CaqI4Ydh
0sTB6G9rm0cIxmJN2fL6NRypX2mAXZCLoHoUKNHPfQpbabVsmGc7pEquPUTV2+kb
VhPAfiLuAKmMLzTHDcoy35d71duj+8IYQmZx9wzcCmXhOtrsRlsIhZiisgyP08wS
zjbnXhPFqmVuu+/HM69357FFucUOXFcUsHGh79vJYwMqGvdOCVMRR4T9tfbgj/OG
xwudlkMJBkJ1FvsUTfoMHBp46ZR//WGyBUTh92qZdAomIY1CZ0/r9HUO5AJg0Wiv
kIo9qeHMGWvYVYol8kAY+FRZi0rb6lqLsbIHhDTlYpg42XnklvRvNZOi74ePgCKJ
GP0XKCXW7COhBryLHfpEzxPlhHcv/wyy5cKyz3LLEPDQz/+TMFjSsjHd0U4q6UOr
DoU91AXJ9Hq0YLGjDX9/GTnlWFeJYSXOgLhLSrElE+7tftkwT77pqoBmWJpgHPiL
mbr8lv08boXnNuF83uoJPfTamoUmZzM4RgcNwBkNSVtkXwqJGzf0xTt4gk0PaGyO
lbIaVV0B4/h1qsH9e3rvbbrjdhapDhnw3LaWqzugFTcLk5kzc1z4NVaRTWD9e64j
8MA1wJtdPET4UzTxGGultmYa3/qRj6GI5FhY44ZHFzi0I0FA32j0E7Wp1F5gB/RW
cV4j5tiYfj8FNq4mjrOzoVmRkP3BErZp6MoqzJ64Xd9pvGd0qgDP48N/xbJXSOuY
4oyrB06WtNnv/P9lbOWxJkq4G8wkDwXmvITlbvwSLFi2QX1lrTftkOjoShjBDI8k
HdPV3oDhsE2BBGQhvFL2HjCgRuuZ9NozGhjNhJnw2vhE9R5tdet8jz2O38R2ILEm
gSFwlbQliCrym6I1RRjV59OglB4Cj/OyCE7Sux/18hl9Rw2eohCvb9ZsaWpfs8py
lgn8KzySwwakvIMhVZovwzdIAovexiMOPJHDrfy/LYF0SFpa1fem+mK9gRX5qssu
AX2tHx/JgdtICHaKK7ndBiLp+FjiUuYahW4Yd6+BK5BNj58WdQROK/IRaWGyha9a
oSzcoULgdptsAOTtdzfNvGNpIjyyaRirNFhrpK4y5CG4x6AFLQvB7/RPWAuCKONW
WRCtV5CAZ9rukPmlzC+T2b5CiJ044jz0CEzSyo66n9FqML7t3t7OeTjwLoiu9Qbk
D/QobQWSYqK9OeEc65g9LHipzSIdnPVy7TAGykMqfFuFQ0F8wo8o/LvQShrqZm2f
H4jpYEuod0wJWSGK2etxf+flr6LLAoSLeBGu3cqzMU+wuYF3Z/f9bdTBmcnobvQa
6uXXrakCn4rxGc+sMqx8xr+MGBaaOlvciBVQNhvIxtceNNEctHuXtMuDtvpIxJ1M
K8KyakURu4wC/JmUFjNpY2E4KBLxomsF7q2/tstIu066DKdJpoF84yqTWX92wQ3p
S8NkZDNJhk2DGUSNL1/JgFQGGT+iz18FeFMfPLqUUaACOSbzNqB0Y3miaqtMdJiV
gPj1VGKt0iMapsI6KGvpaO73QdYUaqPpBalw5ZWdaohjHEQgOt1QyN3rENpY+y8v
Qj3CiOEHNAAUrhLWcQgIzGxDYs60b95BkcwPdYzSDUR4lzF398FLC20zs2tIJH7l
io70WlHjXUmeZb3L5tWwBpLCZT+i+VStlG3xDR8ZLB1ynJrbv2WXXwYii4NmfYth
btQbpVg9okjco63VSjcLsWGZQu9StBcXP0uiKNShu6pmxJxZFojd5ioOkFwo17qt
J9pppvcZ5CGNoLs3/ZCzA/0BXzUBsdmsZNAB8ovqwjRwYcqm/JhqUHbbxnF9D3hn
L7MBer/FiuwMuXVdNl8SFZYIKV2YCBMOguitpyZMU15RAdYpDmpFKcUWwGmOvBJl
C8y39EMVRhuNu4meeqI3y+nLxOccFSWuZPIcdukrVllhXb0HAXJ3ekAp5kAGSuJe
xn7YOZKOdevWo8ZXsOduwAh4nvT6DxUEvV0wRunjPAitfrfY+Rlp+IT/mRHIEm/6
2sFIOph6Rd2gK9QrvOZt7g8h0f7pQJkpDnDuvcHxTnfHysrIs1Gqd9k/zz1iOZGY
PHPQOEwicNu1Nm6y8wFk3mLni0HHHTBuHQiR+xTa6gmrt32fl26wZ69tqRhj8bbL
Av2d8wvz+JJRiiaJKpyQv4e1GEXi9HM+6QH1p03cMe+N+7fL4oRWr8juQXP1cRcU
a0A/I4+Jqbg7G+N17l6JqZE/y+ntGhlHXnicJyvY9J4W1dMsWl0G4M4eNlTS35b0
b3kFyXk1kZrMAiS3/i7GaU0+L8hKwlvt6ioZ0n/jGWBEeh1PFxYfsUkt5fTaXN3I
zUL8jjYljDkjMucLNfTlCGDx0S8Na2QPhYQE1YvG2anUqUkQdDNkhW3KyftboJkZ
6MmL9AoWqLgnOtqZAyRQon9cBf5uNlWOeu2ZeQ+HaPOVkV06l6eR/tAOsnH1O1Gq
EQ+iiFFbFBjCiwueIBlRO33JJw//u/8ZaES1FjXWkSWkDYKxURdMxzNLrl6Phv9B
fY4V+BSRwl1ptV2ak/sXNhaRHMxRRPt3x+v3roRJuIqlItVoBUJ/jbItkJAsDugx
hnOP1J7VGafjna1fXngTD0gVHMNA9kGf8ysLPngPobCJnGVQEVc21ATX3/AepqrC
R/fhQ73OGwSr+95d+S/bsazwPP2HCbjoN54YlByJS8+IPLZsYCOoETLSMoJt0yQy
s3M4MXBUsmps8zbcAC9Q8GK1rgUFOE9Tsdz9XVOirVMh6VyqCzsGKLPygCoBah7k
i9kYd2hM6ut4ldxEnwl0Seb8r2esLs8ocmLeVADQBuLJKX2GgvrmWGJzkCLYNHjb
o9yU9rDkrSs5VNAVQLE5C5he8Be3fuPlNPpqFB9lYwr1rTrtDU8wSdCBCaMumedW
tP5MBTY7NhsKs677NzQGGE7qXAZfV89NLAnVQX4LUPEyF+DtN7W8OZ15urprARVl
aJYYZeCGt/gjuQJ1H+9jLn7q1bSOLPWKYZbHFjCTZYsRvEd0VfXQ3vYZIEUAu253
q50gmEadNnh+IG8uHPuUj5+ka0XG3gMO6S+U6EakF6FgHw3XVojK5Vz6cm0pLTpS
orRxTkHbHZ2zBIC+2UmbVsgMhmo1i1tgEXlwMXBrdFde9UOLsvo92CdTOj8Gvs4E
le/bI+x1NRsNdlZoFsZzrYpIixtu+FHPXd0t14+zbEB24yAsx3/SukbrO1fWujD+
yOGPt1igjBMkxlH6U+kF6WMqp+qeYtQ1u/00Wdy0g3mVNR0Y9T3Irj13NuaIRstF
HmZ3xRvtXmcPz5HWc80GOE64xftHJ2aJ3Forx26rn98ehtowFrGwKtS33nSYioSz
oXj0RI59DD6rwa9iOVHnn1tTntbu0iN8agsakGS++0xr6GansS+V8BN7qInxXDac
TDdQRUqKPqpbjKdUHXd9T33LjTq12iis5Mp6r6Wu9r6tNBORpMCU4Bk02SrniZga
Ygd8YrbCyZSHMYOzYJUtlKk5FT0WqmsYazhmFImrrn/Co/9bZaRa0THKtnTUlRnK
wNDTGhLcPeSSlwln23eHBayYut+bPEwCuki2pbF9EeEFOdZCtHzmPaztEm2k4p8h
xw9/+IKJBZjEM2fbEEdDMK5jsIoTwNokdKj7b+RJPn8ZRfkksc3UHD9jkzWSGk7j
4dwjXYUBB4Q7kyn/COwuBske9gTdyiTj8Iq8mahuo8xtCw3BW4J3qGlldBH7ONIC
2v9j80wLewayygeCk+CdIJDPbRspKBrsczMSpH6r8fmIO9MgX0XvL6iYzaGkIg2R
H7e7G5xJ++W9o3bMnV/vrYmBL4flxLCd+llf6EhRXADfs8F9kkgLqebA4sAIDtUb
NnRaZj6RQs52ye9VRGVayX4Tk80swrWuoh8GI1YlTrxf8vm7a3gFHjJ5ZxjRUBnc
TkvCWSSA+ZTHeaCNMpvnmhP+TcDQtyOWodIUe8hAk6wRBdXd2totTXpQzz+fSzH9
g0CTZ/Lg5mkyhfhkrfM3CYId+mTdjuMRtCFRgWqsgERvboWo+7H/N6o//tiCQhGS
uFy93IPlEJLPHUBYRsMr5WUFaUZrzSUXN3PSDHFvleoPVwo1L8kCPtDrV8LoRIg5
FX5t3kNeCuwkW27GPS1304P5m6buwzitVqcPLekOhHlwojU1/IFeNofErtya3gD0
x0o/+J8n3ia9h07BZM4UBPWWZ7m6nN+ydeNXQXiK6zXLelSYg+e+Bs6bP+/Mw2FK
i1FG0AmHp5XTDI5uOVVGIH1UKVjAWq+jylxBgTez/0UTnAq4KNAjzYXVkvo6VXDK
qp5lPI3WH7UUudkNs1RrJIyVCfOvN5Z/qoRcP50/FhpoXlx/E1cQIFLY3Jhs4V+p
lGOuo0tlFOetnB4YwVlLobwD1W39abHqm2PVuV1+ZcJh/YWIQoDa97PeXzgnBEWj
59maR0UI9ThYvG1njI1Wd/sib+scvG9IEu6v9AxvP+uIXkxYgAe/u2Em1tOPxlK4
lrScp+bwnl2teVDjhbkGXrdL2UR20gCIQp6sBeP0VjTTrgUUBLGVLTBVk86ddSTA
JfZWrTT4Yr81XIZejE9repGKwrRlQobqJHqjE5XNmIz29xTaozegfjjnYkpK7LKf
UvHB4/H/4qMFnaFtg8MItlFQCrgr5PZzayJjXzV6NzGPJzEvHen7m3XiUJL/An8j
mZGgwKplNmWnpBvRfjOxsttuxGS+VlwfZ9jX1ZU0qJbgYmHPBTbCavlBL9WHJnf0
sBtPD/eqMrO8lhX4D8Di5QnvGf991CpShlBtagHWPF5wvaNXbsE1tVZ5t9yH1V69
k8SRh2gFQpM5bDxyuN9U/fLB3CQ1FBRKAK8+9hbGOYIfcMbJ5xoUY2ottj/L/UIc
1OHoMAlvRmnl+Lv028gzbvevxXwygijG5HGu3eHk06d8S2olKe0K7VFhUwOpLvcE
89zW70aGUeWsSJpPr7b3QvU6GZ2tUu18hjjzJ/zL4NRDyqDtYCOW7wx6oWKLGqJE
uERNqjUSxDzjlxhNP4yQX/0aVsQ1+yTjg9NPV0hAk/k8RS3nNfRWi0Jui/iLbW9W
AjMQBn+CFOu2RfoNbe0NTOt11l6OkwYs+Q+5/oWDwlT1i8G37jTuPjNKRDK3mIAH
fNWAPAGotHVc6KTj7w+ePkYxmnfXf2ERekzwd4pVJd1NWZ+f9shC/DlVlg0P49lW
AtdQcfbSKjhrDfnV/dtmiyj8qKBvKnt68r6zJpJAY9UfaJv425kcA8QzXkIYkaPu
8s/EvRNIvUTchOeXJfdX0/znpON0PM/fhEYVr3Kjfn+JBdx/i8K+6YOp4W3Jce94
mdX3FzTS2zZqe90II3yJVEhb2SyMaSou2Af6dzLtZkzKUGbWs/gNCHlmfXa6RSha
Mcf4I3t7aaXmaT1jgy5Ow0ZpkyjlotMbU7DkbzdUMhOZjNc+6XUNP43LUQbIewRS
svb6xblihOgOHiEXdZU9u1G14G0ikcHO9gQUuXddFuqrWHuUL/bb+L5JYK0Sr1W9
rIz5RGbG35fzsLExn9EHp7mDP6PBpNMe03VjD3EBT1ql2Q4ri69DNyskoQdS0kDB
7Tm8ic0/U8hY/qrLEQKUtyI05+RSHyJqCDvVeaDEkjyAkITQQc6qF90fyDRH7QIe
jglKhGgt3FflWL8reXfBXtWaSWi2nE6bkyuwutDIgGgj7Hix1OuZ4353sneKTRgp
mA4WhJu7aIfVro2FD6YXnvY1S5yVtKVqigyB85z4mo7qDP2klW+/b3cvSQX7Ob7D
f6gd42BXhKfcEu08A+2j6t9ehm8w9rcxNFPrfsga0rvawhB8+HamS/EOKuKxeL3P
6lRjWQc3ZZTBIFsiN4rf+BBII73qiDAy9hpuJA++cxkIDUuUovlxOvKO+NvUMSRW
ZHd7K2GJRmMV2r4fN1wj7B0VUp77gKHU4h3bwXl0lui/IDwu1GDinkGO3amP1qh8
NnNBCBeDhZ3Pfbjv/KNcwtksIziRq0BCZ/QUpm7z1ERHjVAGk/e7PgN/q0Nk2j8F
G1jsbm332jY94jkJG3FIY1mUW8huQIjDInNMKQWGJK6pBDfTlW7rjBSS+7tNxLXZ
2FfWN22erIoKxBvZpkQE03/VY4z7GNfoDoyx7vCWNiHs58WIVTYBB5A1QZ/OGWQS
BqLV2cDng675VP1n0PIXuFoa5IODv9qiyGifmzV78aDXoSQd1RYDvSpMlISmVYwq
SI8odsgFSQkcdjsK9USpz6UsWOGe0X06BLz3tqmMcDr0uI21jBfYHz7cmQtXwAxg
+ZDPO093/Wt/T+El6XEXGW7EpKDIuCg0ZwsCG1i8JrEMioEeqfwOlo+iMkyARlfn
WciEvS1AnjfcIGN7Ve/pE79dlhesDcmIjy74Oy0pV3XnzI6T/NKa6ehSUgFDr4lP
noVRAptkvU1MQSrN5P7J0QPfC0UiCq8k8+qEg15g3LH+1yM6ud+JMC5w6AAhmec1
hYny9PUnrGAr+QMxPAONkBKuTJCVYpdjdlOjao/k49ZcTya/JSclqn7i1b8IFOcA
dMCLqeb8BftNx4j1UKoJJ2l9X76K4VfeGwD8xmCgiYDP2k3EhEuPf/Gvv9Cj+kn5
cj5vSVij6kgWTQlHqvFjaeXSrKt1WhyO+W4rNn0QeclGbKd5nRsE6uwHrLzFgyQR
6tjPszBPpM1JbqBEMVTDeZBqXVYR7t2X4RLT2YfGwjBPIXVfQJt4xH1A19V44cKs
kmEK0R70lCFV8g6FSd6AuJ7vueENnmFJ+HxeVpNkHzYgvMPzl33lJcJI8HGXFY2X
Z23JakLo7/GV/mofjqeniIAAk4dyzE5X6qTkuh9rOA7pPecyL/PjyFZantJL2Q0O
bqPr6pDZFSRFp2JzYp30W5dd5IFdWSJeBeIS1fQ9WIsOi914WqKnmc2t29HjhMj0
UtPdtfznxWANfBpbYoxeBJ9K1nHNL5QeWF3luiIKfp8Wpk0Cczaw1ktP0efRNgDG
titRUMmtr0fIJsnJWV52jKPhDKRNJdr/tr4qK8S8/hAkRzpHy9uC8cxF3IZttc7F
orKHxPIjAjry8fQN83ML5S7xxN3qcNCk1dsGKHNyehG+GyQeC4Oxluu6MEIbtkzk
guvZAo59tKKbvAbZjf8tNLdROLwR5gbcJPk7S3TW35hPcJAaF7wSO0I64q5w7nEx
Jz5eaDsAuPd3QFkEJ7dKEVeeD1ubs6GsFo2vTJHLHbVrEQQ/Nn6p5Wuz45XpwBOI
Pef+QplGf/NKu3mQyQhF/ejzHpiUtmEVmqfAHUdMXZGVpnsHuEPPvGIZyDXh3q5i
K9AkDFCc3b6SsQy9nvGPNs3AdvfTWYttc2Sz/M2AZYJTJ+zsWtFrYq4gMPvL3DDU
p/zdgOpv3rsEsBUeQchlA/R9s+yLflakcK8gFmfIS23srCAcbvauzg+tv9ziFIY0
8b7GN9o/afNImm92/xyAAjbMfIs7O+SW9JJ/EzrezW6FnI8F+1nHaJkWcFqZk7Uh
yVsak3RvxKh+jd3TFhPzLimP51Z8Kfvzn/gJa8RMfBVmAd/BVpXndfKoD4cLok8A
Irk7X7EKcWrHEfqnLF30+dfyk3WgoyTRkd0wMOn1Iskeoi6Nt+eRKC3BenNrBA4I
iaYUJ4DxNHR8NfBM8ChmlOcO3vCe9AAZ47Uj+LJdoRPkRvZquooSjIaLChZLkaBU
wSd+/Mh5hwstZFXjqOd9tggZ2njogfPDg78l3fysgHb2Wh/qt0ESD+To0gOpFnBC
ZMEru3Xxn9eNkCZkYpkSdw82K0K0hbu5O8aWn4tFxG6W0aWDM/jWUdp74mG6btmD
zl+N0KVvwCVoPfDYL9alL83e7v5TVDB30d2U3V3XTvtH9eQ5TS4nveheUhB8RKnc
TiAo08tW9VoVUGdJvw4pKOTiCPDM9KQByvf0kzAj3P7hFgy4GAjH38bFJZoZejv8
P6TlLzPxNhzXDeqQKkpEjcm0CJ458Vc1qRCAA2C9/2L7FshqZI+DZMFAsDXUUuQr
2qtiGbthvpVaDYhFof+IyCaHpHxDJhZwxCcpk3MIP86WHEVu7ZVVAQSk26vGS72w
C0DpaVuW5RDBqoJL7aia/0GlscztnAbAHqB5DD+WtNjOY9c+sLOCKmTtJt8c/B9o
ZFQizVrDIhIvxTjKDTp/JZiopJNsgoXRjsGg+NlMZX2Sq5fXnWXOoZA+PJLc7hWz
ZmiSk5hUZWz0IebjiIfODoX7Chv13bBE4hwazIayh45IHBlHSJ6OGe+oTDd4meE1
ta3cTV6AGvZNwjRUEpZQRidEcexeqWzb0ZPyZCEhbWCFrU2lb9i+C3azMsZ1Nk3m
xwxhIL+kHUXB5iGZiUQeuPPNdsarJtI0lHSwyUrJ3WTY3P4nufXrkO1bVbufgL9g
BIQ7RgMfIZoZSRs6sqKJeJXRS64D37ioPdnYSfCyi3gZoK93PAiRrIOr47ko2YjH
3oqLKiRM3v+tizMri3fcFQp9i8jEBGecOxAyQ05F6ol652uW88AvnvhoaPzxAz6d
1OGwX/iyCqOhSaXwgbtkymYLc/PMVedJiYL8FBCSKve1Kz4za0AOTaYxfEjyMUJ5
WjAqqi0RafslHs/1/TSZC0wAWHlz8IiTusVjMA5dFTodL0qDS4D1hAyp9XAYUmbE
cvr3G6ogwyfb42NyHQHtqenuA/YJ2R7dRculNInB49DRmGjNuoP8ooqLVfGhU0e2
smTap17nUaBpiuhDehRFvKex1svmXmUsnZfoEmxz7xbzPsy7T4/+THLQ39AwIWIs
iQHat1MXZM9y+gLU+tzCn5Diw8jLa70ZZtgb+++2i9cY0e5A9mRlQ1jsEIdJhgd6
lDbJvkx6XY6G57Msc30eyIaqY3J/qF5BZBgH6uFHzLpvFaltf/XpSASSJFMv7yYz
02wr1K9bPnterDXqgVquZpWiyZdysoLSqpJrdEe8oNv4XJJNIOJkQhwNVBahk/Pa
KE8nNlcWmU+BQij1SakrFTQUrjS2eV0CPWEMirtHl+Il5D/mrNHXyI+vzCSa+0zf
I0BOYD/4AABEiYGpAvRaSHU3fKVn3T39M5EDVyVUWqInuChoCkRrhsMRs9SIczah
exBxCF0CaHYr8e3i+C6FejueNJXz1aE+p91ovRLY02oHONY04okp7Ke0mqGyjktb
PgYHYsUWjHNGLiWHT5vf5B+mtVCKfhxOacWTQvml6F8kkj2yP7JAZYQycGUTPH6w
BILs7CE8X+4jHzfMuZMzFq7avTu9UKQJzKaDiFx2uNjC7wnZ5/goX4Rj29n/kT7K
rcBiG7kWX3wdVuxgWvFt6FCcLItBA2Zb8so9Oabm5D5fY59SJpm2oLorY4h4ckeb
uY0pDJuQhJy1btLANzRElllLQsDsSkVDu11n+PJoWu0crxd8ElBcx6W7a3fo8NHO
/LHgahGmMqjWNZGpe5jYuV0OhIDUsPfdkmXkEgx0LJjWi5EbALeHexniwHJa+szR
lCi44PUEoRRppa+BHKokOCpHpoiIdv7EPF9JI+FFg9OYooSGPPPSn9IGqkS9Bufc
uM/nbhjtQDgtl5fid+IjXhVd5M/go60yuk4cKLhmlZA381073YbJ60xHbXhZ+qJd
v4hHIjoypQ+mhMmZSc2w38kPqwdc9BaZeqH/B0CRlOi/cdvHI4i9PYrzN/J1wpHl
LeielR5ew3iHDmzv0mlrbs/3DTr8lsl4KCIEBEuErR0BTqMxOyffAjnVFzKnkuWe
ZPBHRr3b50SMyZWpZjwRmW3u++gcqpFn6k+IbC4YJEKjp1iEVWfl8TqUkk6tAfLr
6zAd2N98R4a8qSwVEcpFzQZgXESSP10J02DKAyS5wCMsUfJ7cF/Q+u4LxDMSKZK4
TFCaZ9LcXISZsRDcmLo3U+58KPHhXkwzvrX4P3UKfAmc2wh8jHj7yeXPec2DZfXv
ejBjfoJASqlte5xB8HXUYlwoc3Xjpdk0LrKGy6LNBFAc+AnDjtWXnn16V+cVe/10
cDitw8MEBlx40vtuPLcvZEFYkUB7N2/xvakvOea7lWEBllpW19w79k9VTMF9qAVA
RefzUdcnKjLRGY71zn7Ilu3hgmMFOPlHHGCnncgwIr5CwsSHaxpbXbEw3RFNyN5I
AGAHGaS0wl7p3juOUV+eZE6UkpkDxFnPirwei/XdLXAjTgtWvpJSMD7v6HY95Nh9
mH4/eD1SJbHDeDHScvAWPRSrTFSmV1456i+T/d8odI0/MFGZP74s4rqdO77DCWNz
0ys6WlylrowKcHfn0mcV+ehhBogpSQf1K98tPw9yA97UteOG78bdVBwGwwnh9ALa
3Fsuk9wUpP0FGkOUyReNGG4tX16m65TJ/huGkjFNklgnWwNqp/caKiy99OPKX4k3
/krY5FbD47OPUhSyDQxiDj2+t6FmlsmCgenAJY960texgf0Y48oXp27ETUzY9RAV
LAARGwHrFhet6TSZu3GCRYIPBxuqsWakFK86ophGH25lkO5g+wc9f7P32anPEtfk
bVPRUqZ794d4WGzN554Ow67G3pcTg3LjzwXhSJoAvhNETuObtJSpq1w4cxvAxKiA
WI10ee5zx+wSv9h7H26/E7Xnab96yJE3vvnYZIAGd8r1kZ3o8CervGoCZKYg5TJD
DGIv4AHuxrVNMKx9aSqQyjfKs/LMuyj3RyVyflvPTOb2kNy5kHKHX+KqxIqOAwkK
Qc7vqMMIa8btN67BHUcZVaMeVQX7Jq1d4Y+SE6DZHF3xOI4czJlBNdvuKDtbznXp
Nlhh3IPRnoGRr+r7KBS5B4V6Zy2B7l8Y+La5ncVUEkJwrPLprGJJmw4BfY+xRB5v
YNDd+Z4RY0NSV/G4O3K9IQK1TD7MwBdaZzamP7vKk5gjsHW/jZEvq7fsRFwFV8lN
4GxepxKqay8OLSY9YRGmB+vZVbxE5obyb7aAd+2saO4QutNJB2ciCJRMuYymgFEY
GGP+yByh8Z3uBEr+YySGWatbf5HnQi9YRHiYyxuZpZFn36PuwKELFE3gu7mnMF8N
chLAnnJX0hlSdQFI9zRZ9gQoUptzFDyoMONN9KBdq3xQusAaTNCHIjn94uHjTlyT
sUII7wzUuJTc1mFFso+czpP49tRfMdRUWL45yKckqrkIzEMr4wIAprr16kjFxei7
21/dU4yRd5ypnJ+FBLfWIwWpKj8SbyepAb+rJ7FbUUn0WJaHeAwh4iirtA9p7e3N
Igenw1NtQY/Nxi5qmJ5GXbpBeSWjzhUf7Y0QqPlGdhSTOaFCrTEwvv9Efdc2qoZa
ifghypkIYi6NA891MDc7LTOjxsajWWj32hRa1VMcKq+eCzHo8qfpZVfDBmWkwqJj
RhKMNu63iwQt9exYQm6kzWHU/OrvOeVz/gq68eVk/R+yOjl936qvuTjcQh2rNYgN
Pdt5CrScgGn7VuUp666uTDASPZ8Y6PG/An5TiA2H6v4fd4DfVx5jh0nwoe5fHLar
Pcwf0Tc+EVXDiYv80BzrUXFREC9VpFDMM6u1UY4Zaz4SsfiZP7T4kMLR0VR0mxJd
G4KnPfjC42RAkb3uxFWX2HnPApXFUNg5wJIGdD+mf0EhNlDbh+URaygas4phDWFc
DzuTm5uDP7/IxmJTLZ63Tnj9Ts793pzNqeUHixFn9OqgIrBdVJMuX8Q9xAO7cZ+3
0WnIkU53LBQX4f7TTi5/jt24ZZ4eYsHsuUwMs1MstGmpDBFKNiQr3zTP7vRRnnhj
d6HQUhbFq+jES8SHgm7hrRQ/ru/LGLXnjWL5lIC905W8RRh66KXS+MGxXzNLwbGr
zAOw9e/7fKEJqqdQoBUNcQeH6tEmSeAIGuqiJ96aPv/qBvZDcj+cfktoVl6kcLBt
ByYhmTL0XmawLlp1FAxeVelUccTG8BEwbxtcBswfLEjYkQkCJQ/uoLye9Ds3bYEK
ikhg0Be64U0qIX63bViOUpzieotPuD1kgxNDdZjfZnQZpZ48HzMY2GOzsPcBboCz
97Iy1Lff3P0uSVAddrA5QzrvfIFXDvxNhxHU+GFvNtu6Kgnu3L8q38toezl0qwaU
+r69X+W830KCoVNBP0fvnRqONUFGkCK9r1LVzLZW+kpVWiHyXe6FMVTY3C1d/63o
JJTavjcEKgco5IUHs6zeGWXY15/e9Fx67R3K7aETeTkbcWLKLuhBISp+cxyYwP7B
ocZmyqnr7+ixwU42RxK75PKxZZCaN1lL62SC94w13UqnW6ECWTN4EFluDijUTSzK
w260c+GskKcC+SIIo4reZumJ0saxLXImVQqDopU4jpSiE41/It0Ig4Qv1wDJb8lR
gKRlYw0/1v4zikJFWAgRhlST9/rO2bsO6e4QLNSx+WY7QHYVe6zag5C9KwXSBNZB
4OpHJkwARGtMG4wZSsLUkqj2HNFyjRLplhMfPlpW3ybDe8HbA10xv3BTP9P5e1h0
+AtOKPbZrf1Ascs5b8/s1mxW/AnYNy6uCj3NsdgZb0i87hZbMLnxrA86bPk/62kO
R2hpYhumUrvXkkCkFqoJ6p9SgqgUtxH0mKTcDth/JYLF2ixPnKrYpIdF+ulJu/AW
A40baXrgxanpDglXOAMvQ0KuvKoNw5LFTyhftectRHkoGHBSzASLBNzJSeu9mYVl
dgtaqMge694wg3Mbo8PIFLzkEdIBQ571PhxmsNgjp9EDtk5/LXXWoG+UQzGuLPxL
80ydR6djxoi7zmcG5rv6k7zNWQIO+cbojPAewDGpdetKDJWgVxUDQ4VasxcLnVyV
vzIBQj/KiKX5P7n7cdGYHio5PBOcx0D9WcJ3kIyZgmNTjezKxKUW3/t0VnEfNEBJ
JVC9cbHH9CbauDOlO9UAdPzvIq70ITuQhyxFHgwAygxe3FZj04rO+iRpQg7XUkb/
c1MrQacCpVKtLhj4BBm6eujPx1fjaU0UG2ahkbOWyaE2sSBMFb9YRe6d2wPwE1Cl
bbxLH6XrT0m2sEgiT6lePQ72QgFVEFjj3+hxVQw6UJ8o3dVIKAc51eYh2r9h8c1q
JZPg7st8x8zLmbALm8V+OKVx+P+4+fu3n+qDbRYT3qvpDXJ43KPVeOkaY+kI1IuD
73N70mzKbMZ4akX6wlbmclptU2SlDe8ow1C4H/F2DPi5lxI2Lvr/vb0mJonWf0cl
nAiv9jzb0bchC923EwBqJm3AGmm+jgGZhjH6Jo+t1oj9x7jD/EVvxVBQ/K0ho7QB
92dHV8/5BHN/qbp9UU9ETe8CJfQAxiavcUI9JAeuFjtCmkSL/b96ne8KqQJmpyqk
J9H9KsjfCJNrVsMP3PDwfEMxo4YAZQ9RfawryvRe+4IqnBoP5RqBOUPwc5EHLHic
azr+aqlz/6QXCev4ti+uN6s0wtOPBkvt3TZhUxVJojn1kjguc3eDxbtqLBvCG6OU
ePYjf6JJl6JkiSGL8uLmNZ3yYJrZIQ4Cv2+WkgrRXXbvTL+MBI8WmuuXBhP4ab4D
pNzbXC46HTSdHFqymoJihHm3Zx5S2alIVFmguNs2WlX1THdhw/PDlxbxslcpWkvL
h/34yL34AeLQcuiPgN+gGEoaX+BdNII9buxm/UkjyZpr8tzkB+vD9/gCBymIHRKj
O5OA60lXOLVgi0752czLzrWJJ+ZMKKrOw8E4BlvlGSb9gUt33FVtst9e/FCnPKc7
JMrItBdrtlVF4sGy9TyJ798Rh9dB7oRj4dPMT03in9QNC5RTxkkvJkANGH4KF/M3
pTFSem3NEF3F7w0LM2WY6/0xEReaIFzj4L0RguXGbXoAFGhIAueDvlF1T5OC04q3
zgHtSXshArZeN1wromPcohqo90wqKDr3L1wBCCKExTsxnuuj0Vb8IK5sXooKTdaA
5LDEahcaXaMhBwg4InmWEnT7oj5J5rfoXwXEo8ZKmbiiAHeEyykhiEQkq1jFyWcV
9535MPgtCllhm1aRMu+jTfe0Z2YRAtUtA74UrQjNkPBdlHhUv7qKR6FVj60lpb87
U50uN8iih6yTT+ZVQ14i1pkAoluocAHIHFAx+N4ePCJnRGOA+riVJsoiwmGUQs83
1MhR8ZKx3njLx//TdwrbBzLb+AiYtGokz0Lfo+0Y6yyDtQFt4kBlIHbZONqqJ3YP
y0iJS16qXARi6SBdp5TkI2mcputad1Ofo3IfGJ/Fy+PCo+pGqlIr0hFpXM5XO79l
GaypnXHp/c+WSG8/i8MRtv+P1Bz3LEh4e47DR/JBoK935WUgfNzh1kbaqJj/flBd
BpRPkjO9W8frUdgUIpt2uiKPaZLHQGlCEt72q+v8F1emLQd58WhWYKBUtxjxSrr5
JKEaQDZy+y4LHHnS3kH4r26MkpLTFe0BXUYZmAf31HA2BFYdPSj93/zYCDAXEaD5
nNc7dTpilEiKY876G6AQ9LtbRmMsm8ZeQzhO8MwQ/y0WXLPXzqjJR3NvQhU+F8Er
dUF4RDAxOCNqby3pkM/NR1tanr1H4FZJfziC14EJRkU9uvEi3ZJpsg1TohV8zU/y
LdXjVnkuwmpliUC3YBZArZrH92pK7K7aQ8g0fEihbKy40KBNGqW7avdTNWYuFOyZ
I2N57SlJNDD+gsS4j9dNCGpWYnCN/OUVa8ba4diy/ZwHjaBgUxTq/ZmsOCdms0Hn
whg1ZAiiR0YkcilMdwPlClQD+b01K79w3qFoRJ2wEOGEIOVQti0Yx/a32DM0qt80
m7m8+tBmauQOjCo/BxgwdN6bG4aACDatdyzi5KABeTUTyL1G3oYsVlxFaV13pgxR
P9l+s2IZaJE7MToKYZkmnlkC000uL6XsPf6XWZS/Qw1SSWTKgGIb//y1ksAqWsHF
hK4K0+Cw8loomnjAK9Sf+cN0i95k7JVTMIHdIuVBI/nfo7DS1N7LKdY4RoGUCJ6W
+K6RUaeEM6FPcKFAShlWF6K1of9xW3NYnZE/zDl45zm9iurUOqfr5U2o0nKuT6bK
+LQsoqsIIL43JappqoYHy91pP9xq2FU2ICVB12UwtvyfyHUAbYZVGqzaWuSWvFkU
LeRbirYdEqRkmRfqAI+UYcYk83L6kkLDRi0CkN21IeBuqKj1dFXY8fNeELFwJGLA
VlgiIXk32MtA44Nfk6LfV8PNysZ+6rpwUYV47EisJ+t7aqsLsbJrL4JBVBum7FTv
75h1UgIxcp3R7ndMkg1C9ToDyqCMiDTmBw7QLaclGhqX+whO4zHI/bEK8q0+TjTa
xeZEeEvC2WWVnl8F5VGh6Uv+E+e1dgtKeKJxduDz0NH2NV9jIPAo0LpcjF0icUXR
RmJ3tY2IbOoCmgjDXi7L2h4vyW87Khft5L6mSDnGxqQIt4PjDB71bPHKHst5aKxy
8N4278nBWskxr1GtDGEFnr1K09pFLIFaxFBh6AGLgPKnHRxvtpF/Z7pK/0wwYgIc
KpxHiI5OHRlq0xKxtHvaxkq49ie7m9htJXqWqTIHLGDq4nwE3K8HJhpP+UkuySGm
RjyJRopdb0gKam/hFHrrhbvFZK/J+s+/SEx1sYEzOrsKxKu2eNJa8tWL9ynwPBL3
iHjvh3iV0OlGzdE/ZUErr56ftMBUlQoCN/R6Nh/RDZbkpUV/6nXzrUavmFVoYI3P
RA1knrKs168zqg0/JuI7FuYqBq5dlXNPx0x0W/9jjrKKuF4TvfBU9pwK+mPYy6l1
6uVD7EGQIFm42La8d8jZGBEQVzgZ4sp0VnDbwkJghfPHSfAYLL/Sx/skV32gpRRK
jZcGYgY6seEyBLhxBawUIMLZX2JzQlUvS5FZbC8IOnJS5tuaCsyNi8LK63trWPkt
EXOLu33kHQ8c0IluExWd2F7i6oOJIO2jVrQkZ3k1uA61vdtZ5hYXKxp1dG0q1NZ6
CYh+Tmm/4iRADkzo7S46vv/p8DxH5nacWh0heH0uOsxMhNH131LrXiJcCkTogmen
96f8HaF8/uhts7FuxJJXLgJFCj1NeNIdCPah95BW04XC0x6oUmMVvxruS9osCVJX
QrzE8yzN5nLAgpUlPdyEnfcVnOkuqIHo/HHbUHj24TJ3RJVZX9xSqMqN/3MfyIfM
R0G/QIo7kXseucdl+hFNeeQ77I9mbwh4uLn9aPPjNCCnL6FMi5TkcqNrufY+5XDp
PHpw7nQ0iUhZrsQMknTvWoXxnU76V2z6mPtDqaBib9mFJTzmCaVbY0hN5ZwVv4ZW
/SrbWjuiBYH3oLwk4HwNZD3bKSapHM5fisHBbsB0gebyWBPWJt/+PkL6PB0WnUjo
VS+AZSN3uMiZJh6ItrHWiQbIn38LZFLVsx5nCJpz/a9S/0uek4AdyEv6OAGVm5rx
Us7f+7V06E4E3/OZdfMQx7RJcEb1PzyrVsqK02gT0RBTaXMv4eXxiiTlnTSpNMzW
S/Ls5i6+9bDvrq49FlctwC3HsYG1g0lCkSgvNRKe1EL9qIPR3zuX1Z4l+PxqYaF+
mXVZrzJDCwP0eZeCdjGRlLKeiZ5q4socCqsgcdFNp13BMYAAlcGaGb/TuOAbQWe7
V+CNTW+RxlyoUqM7jvJLIKUy2NkJcp326P1ltw9lG6nDjn2LA3HNJF9DXwcLinFU
I5RlebWFkJbrx9NK9t66SqZKkBWI8jNEXp7oMVc6z+dlgO3QYtf9aUDQu8+/9AuC
v0O5fgCiVYPINlGsAJ8fa19vz7bQcBRxLYZMu10tiNHJ7Vdh8etfZRiautXtPG0j
01JrlD56wBDM+3KlEBrx1i/UqRI8vtTCrFzeYbIBHgzS8J2uGUJN7ObO+7KwXV5s
GcGMFTIAcXnqxLC/yJGirdDb4V47Ky3eE7NP0FszgFmQ3beMLK2huMspb8iC4LmE
Fz5/MZMcrrsWPZGhL8ZIQuCdIdJEWm9CAEkT1yvgmYq1YgZns4zDlMCoK7oYzmDd
H9m9Hyz2SRyu4RDHL7eyNKZG1XLSK124NgqnagDNpC7r6rj3Q5a+puZzmqZ1e9FU
NVHVAOLofMSvtXk5Bljb/IXIW0TtG7H9Lmy0p/fiMpzr0zzfQNg3DEOXt8umI01C
kv6kE0BZnAKCJOAvzupLCoCIRIyXSMzr2i9Fn2OWoJyh+4fUG7PoqZPYh/SWJ4yf
SCMYlrvbc+14gdBgLzRuUSUhz5/0XineJnH9TNw5D5Ph6SB3azuHNetmxWuQl0VU
fB7oNFdXlPjQRxgjxyyLp9MRvUe05tkddvkcdMc026T6yXsGB59o7GfYOWjgyeUy
yl7tEvwn/Ebuj/1MNTM2uDsEB6R6eR7eZb/kNDZ52x4GgTO+SSyR/PXpqmLIzH46
93ANAaPEu8fL30o6m1BjA4H65gDwDdBTzJ8tjSlS0RzN9+wjVB0X8yqYrNXk2HgG
AQu65Jje/4vLdzST6LqwLPrLZluPQxZgTB5vU9K3g9AbPwXNxcN83YTt91Ndn4L1
zZY+i9tvRFoA79afuktgmUeVIHe9Bc3sj/BnK7JBUexiDLP+nQS9m5zf3IT70jal
yQ03bvz9+twIi0pu3+3xGhhBjkD4RUkBKcyF72PW26kL4l0MnxVECXehXu2CvpDp
x2Jpy+fEEA2r+EcH7wMoMnFMqvRHM4BkgnUOJwwDYmp+SemS7YxT7CgepUoGtIbs
Wv8xIeoJ81F5oOUfRjtUJD6wUT6DrEOxl2CSRrIVbwDs2Go2CYyXgSuR7nAV1Jrx
IH6ZDPEQgixrV9hl7eRj4fRE4qPpeDbYkymMP2l09YgWAxaTMw0vCP/bSMdCKwvY
DgKZbKKvxkjFSkC3eY8ZCAE11Aw2suyNVILmg8DtXPHfNKDhxSGn2Z8f8g3lDKrD
2ZQLpRiSvPsrkVgzvfH3goTZKynu4MPsytJE0/AHVxU9fxYahQMAA/WK9EPceiGs
riLC6V2YYQ87pTKhw12acoDiltnl9/0R60+vItXVAoA/9hxhtiScfMX8uwiGvVEi
zU4Oe+JdSbUHxlkqIpJAylLuAk+S4eNh54p9c4yTey8dRcZLhxeMVAHFh0NkCHI8
CY7FBj/2TzbmGiiGgIepshgILGQ5+qBIUfxbWsiPU0yTgfCZtnT78r45QXmG4MZq
T82rbfaP4HWSFVP4EHkgwaYxf6M5E/flUYIfsBAUptAFoZ7VCSKnYZMPNBZkyhJA
9LtGPZWbEHHtuiSVm/6zP5XTsEECzBEcWEYZ0Q8VODw2YvdKcjvQmd79qciI+nyg
0GT9Lr/Tqd/wXb4t0AZLje2BbwmJMUCTRnMc/Zg3dqzhEhYG5025BGL5o1YHtUzF
lzKemyO9CGMe6fEi3eb8sBAj9dEYXt4gj4NMeMZmrJwsOWUP76bBBbeEuN27+kqc
4SNduBpFcqblAlrt4TqU63+O/F72YvlYbp7fzmDUnBJvQL54u5iRxt0knHwJShvV
QQTPuuUPH1AV0Rj8pQ4Qxm9Aqq4AWdnnpmnJND8/t7HMkvuBAzOtVzFmvo+62/pT
WulyZgQ0pyBSvXc7dPHKqRScZZ5m1flZTy8Dp+Jp6VTk9my0G3eFMpwIB/qKeHZR
H63SuQLO6kj6m0qP8/+u/B+W2h+2+tpibS7M9Ju5xAqAn/PnVYqe8IusVI4W6U3V
4CyFubNeAxihY7iRiwxwx7yqZiUHUx6QT3txSmtsHFhFuypGOA/XSlslI5q0cO0Z
hVNjOic2T9X9Pr5RBm8trkVo/oLgnFSxPxwQRjiJdMYw+yBcGX2EvtKk4Q5J08PK
jn3Y1fVeX4IWtNMMDBb2qknvkLHRdpPq9djWENWGKW6bE4XlyHScL+yTRKm9pyQE
45SpeRsGIRCw244SZ0vapwsGuxylgDVKGX2shpAZD4En8ZaFpGT2tetzGNAj/69N
bpD62S0UEgdizQpnGCYAsrnR+XpiMnibyk+JyN7cVJeHlFpzVBRFiW/YnK9nnSBf
lqivHbjZLhtb3pS226cFYhWfjPcWhXQJ7G3illfL1gSoanAJJEsXf0GW7KyY2inU
4fKgAmXyMRlYuW+Rz4p1oJDMIW5oMEYZCBBkPoYLxAEOnhhAN7DFM5AV/tfnGcno
3/dnsatvKHqGQiyIOJTBAxyQwhios7B8IIgnv4Xxpu97p6ZO2X+7yXhMuAWwEoD5
x8mfHRgnrhuCDAruykhiTPTd0EtfAim6UQGOajlIf98umgjzivPZ5RHLEn3A+zNf
KFdmOfUAqJzUeTKHtSz4U3o5itFhp17IEuO80y1KEdoEnbE0dZsFcLoMyB8ajl14
/2X1+B2Md6tBwsVSJVAgjI6+i5SA3YqlaSYC2MUCGqdrWkirN8X1LgpwQJq612dl
uNL1xUYfo19KsxubQK1Pcpvy36V0Y4CisW+yMD06qYx0B+siWq2cZz6QKc4FLTHK
JuEBoAN7zDOHLJypbBQWrnRy4BFGQlTxLWRwjoFljm2zycJckwGZ5vow6NHHp/+I
PUEYPRUOp32heHp2kQjb4kYafOe+2cQGVA8LFHG5itJq+lVrt1VXUkbAf9tfCqL7
lS+gnuUQg7uOFeR195MSkh+MAW3u5vNATGB850KnEB3zyQ/+kFUQV6NY4H6C2AUk
1f2ORbfoJPP6UuYMQbH0NAVPT7YI5WMR90OXoq5XKs9cBboC2cHanMPMVULjYiUG
OIag9Em1dqZdS2WFPLJWnsjZobPIoa8m0wF7yKbRUs4CwPz7ypZWRas+erK5oPsV
erM6V9TplYRu3p+QYN2e5R5dcYdh5uJjFIKH09THrOQ4L9i9RIDm+OD7730z0k3a
kXwZHmLyv3dmhv26SOmnmZEyPz2ePCXP9DAs8X2nkdf/u7sIJc7YiPsLvV9MBeuw
CD5fBl+QZ+jGjBzW8xiM03ZOGNr3m+ly0sRER9USq1MsPuSlHh6mD5SsO2PDP7fJ
GrwvxmRBC+VfZXWNPxd5dBUSYcf2quFZa/1tTvnoK0wMy3ve2Fxejl5UA8ZKYZ6p
je7ZNr08AC34pBKwwB7BV1Zcchc/3/xTgZFRAQ1UXvjAcVkGSp/jM40jKDzGKuwi
LwbUK5SMd/2VysOIBm8CtNQq8xyDsVqMQOOIu3X9sTs7tBqUSIeTyLQK35R4gdaz
sUwGDccBtpy3zyox2DYEXiXzzXrmzDHJUfVOYjkF2F7vh7anT40NBGyI2XhHOeI3
mW8VlmYnc+hkhQX+CYz/TbQptMHbfHZiFG5WZ6g4opbyEwDn6p1GvYEiYREfhkHi
+XDVOaDvH1SrmVz9SBW9W94IkuhVrO8lAzTGdRwyBHQ8IT2hjS5tyUcKxGp3MYlN
weqZhfIsLco9riQM1PIe8+hi+sHG351w1QVGcNBQndu9tfKi5gcqXIItw+LSqscu
04BBgzPtES8lgfzfzXwDk8vjsdfAfRgpxAKlzf34cgkHEY9O9N9j6bp/S+pHv4IW
vKeORx8Tm5o6dZ/dug3s05b4GwMghelc/QA9Ej5dvwTkSPv7zQNOXt0cMkKEpojR
gG9fyPUXszloPkLG2OiDbjaZlNTbm9/+RiH7CzijgnWSe/U6xjp64qrJ+ScV0R+A
Xr0ZRSFym6CjYLDUm7K9IRfzZCD2L6+fiDU4Umq8xaIkDKe9zUT/GkSbldiIi7ig
ACBu8CaON5yUkDyAIfwJ5pBnBN9CUou5yfrYY+VrAsng9xwBOl8Dxh6xUBx4aFBx
lTSKA6oI0QhS+NxbVKx+Nu7ZaXtUZURuFyycNydiAghengvegortcKr00xmZygu9
xhxewb2p1D0oQfkjg/iRtbgo5UO+Ya2wVk7i7zej9OZ8lUvoFgYgWpfBKgoPvx3R
2rKKNu5RJqZn2J1emE0AfPfDkgSdr/9DwTT/rJB7lLGRi5sgG/G1+/xmkVSNIwy+
WGfk/8ghGRWxhq7azAs0wbLLo8CRSAg4n0S2EahsyuKET7joYX4Nh1ziGZYX/Koa
Is2CM6UK4oc2a8MpDqw4IILJNmW16Udch1VKshU6XD7TWkfiscTShFjqbrmU/MOS
e43O+Zs3qoqlRx3w6Nq9u8MALDlErDwYQGzoJe0mCmZhe1x22osWjqeE7PWkiuyF
pwGXLDAghxesgietVR2tY8nHIql0KqvZHVgg6uv8NQCnvZpNBh08glZBbin4V8t6
iR93+J49nqkMco79S8NWDJHtJDBe6elXVAXZ07FAkQijJDu759as0bZsvgJUcTab
ncxxIP5GMb3DUq7NqUBtvp40YLOCt+vJZcqteXG4VCIk41OyCsTdAVaDYyqXkcfM
F/INE8yKYRRuruQ/c4O1UDm2AQsehIpkX8RSlGgFsBXdZBBaZI7SYsKXnqftaO17
QhdJqr9s6pCVo8KoXgZv0Q25kZgWmvVW5nERVj+m+uVafDgEnGlnxpHz7AbE3Jy+
P/Z0aV5uebNpqaiAh7LMqW9V+L42ZsxiIuTmqctQ3cg36osT/PpHLz2PTnvMtAHU
1gdUet1sEVjZRis23PWPSM1NGwhuIHcnDtwSSHC+fpGqd2yOnZlUuVWly95+LeKV
`protect end_protected