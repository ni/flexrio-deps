`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Jm2uGAVYfY7w9Y5qKstopObZuZAEY3b/Io3MSEcWLhjjnKulVhCBBYAEQrAzzGsT
vMbffkdZgjdXQUg8jOLJXSHZ0Dgbnob2vlppjZs3bgyHCF7MoJ35E+LOsaLimUA7
hlqStcK49hR1hdeBPr/OwfT3UeVrRtQyq0eJXQ1UksinX1G9Pz3/CmcGfTZ/C72x
p9icpt0bkY4/1I4GBvNCsA6FFKH947JqH27OPACiQQRW/K7JToQn+1uhWr3LA1od
lbVrWu8PdZi7zW9gK3jiW5GaPjwbYQGqeGFs3bTKBILjb7sYHxfxw7eDLVMAIu5D
W+OTIN4JiHiE1gCnNEvkSQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="pm+c2fYA/4JT1uhlJGVUubML8hZi8lME4xPobg/m8uM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
nBaXksR//iZ9fraC7WMJWWSrjqRXHxmM1Y0+KKN3b10NElDzVNMlR76DLrcnamFd
2n7uzsxWqhhJR5LBl98SXO3Y90J6BMbw+OBG/MFM/zUulxh2Si5YK5G9GCrG9gvZ
5JomxuZFDu9CzlWGTuRUt6FsE4Lr6sOL1P+hraQDpMk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="M8TXDiNa0BVMX1P60yIvW2WA9jKGGy8GtbuPknDnC9I="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 61520 )
`protect data_block
/5TNZvs8Nu0G+mfp7M8H+iVAGG3Mh5DYZ0Gn3rRNhV8b5CcJKgjQajrRoGl/gSxp
rBAhtT8Vd5eelHgtvBjpvFBA/EBUrRH6CG6pqRt9r2qUDt4UernbZbxC3BC14KYF
uTWOLC/d5Ruad8g2qo0MpI/ZkAWoYg4P/ey+916L3bXUAi6iuy6Ku/HHIlaPt7SK
cPafULQBNY45ZQh45XgULfk5wIB4ti2W0xTz8IpBdskCIbqHREF7S1WXPpGHX0VJ
Ovx9K/NI0PJ05y3pByLZWThUT76abZwyT4fbQgOf1cSYZCM72EJo1ivwxs5oCvj9
nb4wty6hTW3ajAn9XuXPWOcg2a0hCI8NUvVkTh8w3qCgB5MjpPpS8VJpH1Cineew
CEAAHsHrQ6W1kEZROI69uVV10mHaKMJGR2tGwieAZcyDFdVLstn0MtRRQhXguXxJ
vaywObkI/2ucWCLSir+QU53NeJN3l3jKMUJ+ZCN1ThHG8q5bmzqR5//43nhUUmFS
Sicizv3IZM1yDbLyL/1bboSvON/QKQoRRM2HfYIHRES6If+NGFTQky9qcMIjYJiz
/VWOtHTh9at/jsyAv7KXMc+b3m4UonuxWvIbFqr97j+sME2/XcJ/6YYyPfsjRBf7
38zSFaCan0Okx09BbBehfddDgXAkzbERVpvoLrQ/97dTjCMEmAVVJL0BrwGqofYI
SyzEYZhRkPGvd7X5rOvvm7qkiSu1GgdsJJKVR/JRvOYjm+BBnAUpRr7XZtLbh2M8
dZBId8o/x5ixSmD8mhUFUrqrkmMjqYAl0lF8Q6oBudfQMQ8I9Z9Ezpy+f3kHMSC/
nwMuNlCulT7CD8bIAaPz5XaaI4tptrOSVpOm0a+7SYEYAbb4gzGKSRIREn5CA+7m
sDa1/WLAWSXnactNSHikVsommTuvnP4GoHz2IiOD3D78gpZKPuLnGXszpbQJTZx3
c7otvCZZkrZR6e8IzrZSxg9crqVeWpMO7HNjVTg6FNg5Xiu47oAq+7p6ZEBCPsEo
Fz3zyrzAAPeg/XYTVZTcko64Vus3gLukBB0DjBFGUoDlcrO2OVzrswQJMdqNqdnb
i28MTLoVwJ+iS36PnXi+LQ57Ey8XAtIhry9MlQs92GVkSHugJsid2/2xJq8f9fuQ
4Gpjt7gru/GYn86i1iwQFsPBoSNFwqHFTVdPht9NCHhAuHjLytyP2BOgCx/GVLwD
nKmA2cUKY0/nTyJP0sJjb+OJe2L7JT7oFoXuLAHhFMS7E8pRUvag38/co5TB8qW/
wdTtVY6LpnWNPFKYc0h/8FE83HuO++h01fyLmKoJ5SqtJ/gdTa4QvBorczadjqc8
vT58PYX24ECrmCakx941pJpxC9Jss60NGANnyEd/pPjSYvDu5wto2sPzD37J4RA1
Fo+vhne/RMINWgyaxrX/tZe+8AOdYLFlboxkcpYF01raWRyKI34vGNR2d8avJPL1
UzHgNhIkxLZwrjyBJGGLUMa/40Xo2YRvyKXXQswnNW6vx7uCTtQBDfZs7bFz9EhO
aXYSXQfraZq4GOMOKTueD90gEomKaVEqhc1cQolMcikHveiqnaZOjx24czmIitWd
N+oIpGPQsZiUVPYGgTpIjOA6JokHUPTYTqbOcny/5x5v71evaIjEfKQarKU7wViD
0u9RsmBuiV/INDOYTyzecBmUtrhlB19ucrRlcR/7JKmwaIKH7Q/zPjeTlfD7o/9X
kQleRilWLOLEIx2Wirkykc+uicUx0932wngdlKbIEhE/keEN67Vy9BdW2C95EUPI
LhDi52cNUoohYV+LeXHagky9A28QJdtpTxTL+1EwdbmBUeid0y5TDR2NEo7YtbYE
X1SEmddO5PElymcHuCxWe6OSuCCDBAzIbwwzVvAEgYQVSGQ/bB5z5T6X827oygDw
dSgm0rXXqVnUNCxs9DxBWnWNL+N0uEVXkKITzuEqp4Tv1iCY0lGldkuPjAQgP3Pe
SFXAGgULp8R6+pBGFjuZgpM/07/uUic9oEQKflHg02RdgS2qwwbX2P76qyp2HVZx
wHjyvzTLr4nZbGNS+iuuhuNiJtsHIN+vbopz7JRwGRMNilVAyTPmGPmls1vkSRBt
1TkGvHPE9vycnIABD4TgYM33HcPxukU4T5os+DggXs2H3AGDG1J02kppZl24zw29
3ead19I4r6t9n6A2ZoIRhTmSQJeFhPz7yMlAxujSu8Av/AJJ+n6vD2zDlHmV/kEV
ZlVFHyXCDhe2iBd0oqxIcT2T+aG45NuBnk9tFetQrUDez1j9HD+/pa4uRfrXGHRi
SMuvlgIdKoMbqE9YTgGrdFNmEtQKvNAth/RtTF0WTlBwhHrrGIGTclIJpPu8ej/k
3byxC6rxQFKwSy2r2gbXAc7OBwL1A1ep0biyMRwUyJpn42XgW9E9uSr9QkQvO/ta
bqvhreuXyZnEz6+FQEbaybT3S0nIQHfin61wTYUOjKiqk8hRGoR6P5zsnerLDqIr
X/SFM1Lo8XSxrXfw5KEgfmR1hxR2M06LkdPax3ULamOZhSdBgdLBS85yoi2kgjMa
W0j/WNMUS6LhfNUA41inLV1SnKB6R7hSflMjmF/2XpEZjcZnLY/kTQNuIinxkrTn
TXATQndVdKZp2SVMVfOqCMno0ZhKRry7f/q84RmkXLD/jPPHIQRgvz6YfiUGYTfX
dV8CbDSDa7Yc275Iyj98SKEtSuBKvYzhibj8GUuBmyZODd9+8sPj8Nch+LpPrFfO
EhK3SPNRDgi+0eXsNBFpA+JNGq8Eb8JHUBbjonXGsTh1ccSnQs6nUEJcAZU+Zn2N
MZ2FX2cHvJ5CefGiMmPFnAPBqxo0lmg5W8YaVuObcQLkc+AMdrFp/iDA8px1W0XD
AtoShUkItTv4OWg7YZ+Ppydk0mJvWBNCcXnRNivveDJz543yc+m61DXfJQ4GtLz/
s1jzhNqhHnc70Ms8D4errRJlVQ2Lb3bnagxiLW0pcCSURbaYn+wNeT57fg4JG4eg
h3ZPV6eQd2vGKPz1oHDr9DrRARPsRmSq8hq13yE1ppUemJiRXc5U/uNBtfpSvR/1
xCsmSweQ9mjIGANwaKsY3KVwQIJicN3gGqRZXqceXeGj/BTT0IQ+nEBHcaJeiRBt
75XEGgRJr9smI0YS2mvwKoeOTwHJd8ZfbTqMwrSh6ZB4ek3yeMnBvsin7OZzM/VD
LKthoK9Nkgb8ucQ9rvtte+jovkrHJaxYG0hZE8GHvZGk8lLj3T6XDBo5wsFhSpr5
DqGNVn83Yv5a6G/x/fimBAoewLEqVTUTuhSlDtmrtcMeTQFFma1THRhTCIXQnMyX
ACO9ypcRv2JTzw7tYxL9ax11jUEoK1TMpuzXKIOALBlbjx2wn8L2D4RXfxHgl4dV
g8xwJMZovod6lQc8lQpjjgLO3S6/gJ+LHlNe8Qt0oM+DsA2EOBzrxvUJXedAujnX
PaPXPSAgSJevgcBr0SgBXsnpFFVLf3/Q7UNdXFR3/MDuFefD1HZzNyNRGQcxbVvq
vSdlaJuPN5uzsdfo46VOwG9rdssGHEAOEQr8K3fPv3Rht4kbYoNXzNt6uook3M5y
io0/tyTUobPH3DYJMeKgKvK7fYf0WwDYYoptJOAdA3vH7mwNRRZxmwPYsakNf0mf
v5aEVNaRlSgGAwHcv9NFgiqMZ/AAoupbjFiVKGt5R4NLkhunO8lMigkPIsYwjNth
6eYzMiAam4MeabjzA+uBHsb1C4z2h/st6Diz86QlH4bVnkfjKCdXduVzyKWX6U/7
RRtFZQyFEXa2K9w4SV6AQHZuZdHana8nYzmvN5xGX1UqEgOgw/MHh5qodc20PE61
uBUToTcRfrx7VC0mY6XfcNGgKA2XRkQxYcASsx1gsWxCxzVx09dA5g0Ng+5yzc3X
qfkos1ll2dBy/05ZAg1CQIXvAte+pymReSggpVH2UxS6xOCSRqgKPYiQPkvstN0s
4KPWK97qeGWv5h8zQjYT85CyOHgjhi7Es8TA9B+5K9jnxnDUwJY0MK9uUDY3hT9C
nTXnFMvRLSQxSSKQz9YYqBBl2dpbyt1Wz8yu71IosYf4JKcuPOuOSo1A3NCH0uVD
4GgvGpm2uG96K4hAsb+hEQQcwGEVMB6U358dR6LwiQkJFvnOSZPxZGdrHbv/itCD
lY9QqVAKkwRwEE+UCI+AEA5N2LEmqHkd2PjWfn810ec8X1D88kKFo2JsFouyzirK
5ogSkXm/qPXV/Ym3OhqYbzo9ZWPmobVn7s7GLxoIMnxYK8f7p+FXq/ddfWbntle3
p3pJ8jIR3jJ4WI7ekv2ZraKiOZvGpJPmxSNVx5kh/Me8YFya4EltCw3pLIXW0nXl
NJ1kgngcAy18zp2eNRnGsUv6O08tuODngcfIJvg7jv2T0DOkjXOwUWnslp2XZPqh
kX8EC8VULE+cg/zc8qNx1y0upeWujPV9SQkNZITef8TjN9ebtI280KtS2r3WLjhK
E9j+8Gw1DIjCWxoIBAvh6LArP2zrC7ejjP5fUwoomTlEI3edXyjMnKfKyhk2eF/w
f9rB8B51zbS7XAB/LDaHtMgKv1iLZxoqObuYiRoq0DPYeMILPp65RNdoiZdhIjl1
xlq94l9rruxSnUALa05STddNGDOVhLRZJFpldwAPylYV7zAUz/fDda+eVG2qe46D
EtqgwVWp1AAhdZCS7ltaBf39GURAcDSbTVq+5ju+B9CZMZr+vxsjbmxDM7jNE5Sc
PtnUgm7Xs4cBlhMG2GTlAanVQ9Qt6jZkiD/UJ3rn3QuaIlE/i5/Z46W4ln7B+3eG
fJdRxd0GYU90SICU3ZnZc5uavC+z76p8cQk4RlpJk/o5h7yiFvQ1nbUAyL0WwcdE
EmQW9NUttfOrdVUzkZaxIfWz8yBX3GjCMhS7CsKwMWYhY5MH9oTvB3Q6wZlIyOt2
i2Hq1GoW7d6gqpVeSAeVG9zICBuO31/dEukQARhbdTidj2QEzNGXmUh3Rz3SFTMc
8KvqXTJyQgvGCv00AXqoBSMETWHE9liEqO02ZguB2bdU9rn8ilIqGubk3ZusXwyK
U5ZUq2P+fWscZzQxTZHJHEahaokar1sCBvwHO4d6tiSQE8WER+T0jHHA8MMRpjU2
ytm3XeDZUSSd3jMtxkGlFWprsjSsyv5UraGXE9yyX0j7n/v3yBLn+bNbvUoFeuG/
0uawdLdYUqtXqKRfKJIu7XhppZprbqxwpueDRQvZls1v0opxrZrInyw7WZvBPRpJ
8yIF+CHAiUqnlIaFzWrg5eEl1MUe3JXz9um7yi59SOyXlEb/KqinKvN+Y5PGDIF7
7DVhTYjjavXMzfTL3D0K9OLTPjVUzM8l5ol3qyt3sPelKukdbqURLo1D+2ng5J/D
MBfgn36TvzcJ8Yu6x+uGusA71aqbt6W1MaJNeS66mcTu0OxLAK7QeYiqexB7zSRo
L+RKQSDDBzTvoedhD3zD1LrXJAMAsSzZU8Fp/7P+TenNfTuHblVhsVan9c4mU+BQ
Dzqtv68a3iHj/TLk+lwCaFggWHSG77b4GoZC0DuEVSUe73YkICYua9OpStEumu6T
VEVGBX/Ef57zl2yQmScsJznattCmrJm8YeUVW7SPV15jJ6Oiihp5zI7SjUcU1n2w
R/lh2p8uN3LGCmBUgc22IDzrNQcK9GkzrOWnIYODOQ0B6JxpyrAd4eUBq9miAIZh
ifgt9+dVeGpKpv3WCOyrttTCBS9akN2mKnu9rneSYZx3s5suOzkUxcRodCbUAN9v
9U018GcxntNnaUTKNa9v/RrUm/0BW/8RJONIL+u4iyUhf/K/bEtjz2IWg4nHBN5V
Jez8wUulLg0TV4opNWhYvkVnmTqzvq/jSik86bE2M1RfirK+xAt8P6Z1Xr0b599M
uoL52USFglXnBDjFfZnYD5StOcKliX1r3F9CjCXffD+K3q8yGLM4fQs2V8Rm0iz0
U2dRB8XIMrN+f9HH2rJJHB7Oja3LxV017VSErsmjJUMv5MiU10bv+tmQLVJAZM6F
BS0JA19KnV/oXaDUAtkNvENrJIdTwHK5ur++aNbsAGcyoyCFrdNb4TJykCCd0V3d
pCJE+xUq1XpsgjX4qtvGJHg98DTePbWcYDUnHaYDVXIy+R6k3ng88LpQM6awscHx
4J+xxVooNwUbJD5ztR45W9nKPagTGyYgWdbcakaSXi3oV/If7PVxh6D7uN1qjA4r
JiXwM1r1Vl/XsnINVkepTb8MJ5lPouGhouWxtaTe7tghZFNeOYE6OZx/JklnAB2a
vGFrr/mxgOEsELwCiapFqLEMDAHqU1c5JCc91iMutPyySrkDhayjXm8CRdFdZvYS
ac6YZiAJYEyjdz84b9DmwzEa+yYqOvGAgJKDtbtz6D6z8B/Op5Q6fUUdkrZkB74s
Rc6J0JU5yXEjAZpXgrOfrjhKUty6CVlnKqAQn9g9gn8Skx9JOloitkYH00wWGC9d
Ab9j9C/moqSaAvUxhnjt9mH5KQNQwYonxO/J2QijTIrCr0/t4V8zvLJ+BmIrHiJI
Z92dNRCk1iC1BO18AVK+vqj1AJ8QNgCyUZ/iziZQjE7yhUaK7uAdh78z5SOBXcyS
4uwJO0BG9O9YuDnPATgqHVPycPmJNZaCpe/xrps+wCdtikcZNXLhLILQkMTLrjbX
6IYfHpHB2Lb1N2QRHHJ+K2DqzSjgeQ001usiRRtiGVDCRZUjxENwtqOpAxWl/Kj3
flqhihBACrTZi0+6hqSODxjagzoYMef94Nj5ATN5+ecwrkxcZsQyvnXwN3I7JINJ
SBpxrEs358iSFck5GIfb8ltvekn0GWe9EoG8cRhhzuyc7VINoP4fmkBD6VEyxWDa
EFoKr0AO3LSIkh6wLZdIK+RHPuhX8fJ1JwUCni8qoafzT9F9lg3ughKS/KpC2L7p
7soG8jGOxKwpY3BUjvqDBwyvyQ7pPrEKJQMQWD7EVg+aF5DhL+mKloi33FKjZDgv
7zN29TQyS2sSC7zvf+7uk029s3KEqqLl4zdFRijOxhAmN3EjfsteUHgL2B5ZGU8g
pL+CBKhfll48c66WdsqFRxvWRbbrnx2msiRbkQzXPSpQHRSf4xtInL0Vuc3q4BZx
EIpnDIdBB6aeqdmzRc2aCCi/VOpgmUlTEnlyATZXf0QT6FXzqx53UawHLfkEk16e
UuN1Yv3kbhVVRL9g5XtY4XxorSdnU1yeZyqU5zZ4K3Z+UUnFyXqIQLg18rjSwNhc
1fyCweuw0cQyevPTjYuNt47XidPqJhBTol1LfohXfXpNnNSdUXrdPqGZIGAJ+5Nc
gIFwU9gIT6lQQOUzLAdFbEO9SMBlybTLoi9GjxmkTMX9T/P96pYDE6zPMjw6ji0u
TnVhvNLSYaApRmJEwklOJ+GFQplNGIRFfn2vELNQ2Y6f6BGuCG/NN/FAnXP7DdSx
8g/atqdnuTBhkiuGlBbhrCP81VMZnym96cPeFF3nV+8Hw+wSv5oOJxcI5K0FJrHZ
E1nMIg8wKVcuqzGhLiuJY8nhGt2l3TwmPOKmKK2Lz4IYRRJkLUA9ZopzAunHR5td
uIpnFy48sbsCQsQa+GChRmdHTCgeOsvOSMuP5a+mECNNFwS0V+LtgUd7YJcv/AY1
ERuxZVa3wkr3RqL6q2ODK8c6kpQm2f05xWHSEuOwEgcmf8n06rA/ReZocfFPq8g5
JgA3Z46zjXItu23HyDOawtbnEAjiE+gHhQDajA+obsjQ06/Kr8yKl9pRYwQnRrxG
j/YvGFusavMtqZlrw8YjmQYF1BBz4aZwGoi7pGsysFTmRxE7jfXTjADEXFakubcz
3Ot6O9JX0Me3TV1NCa/KI8n18PMLDqd1ehLH7QgT1UGLdVdFSwqeT/BivQaN9b5D
+2lKUlsPHGNnFFgb4EgOZevvc5ze/u2sk8UQOhtIl/551Wp6QUjonPlFWbyuPDoz
VB3BfeR+LrSqmB7Nxy+BLNitJoQOtuIT4ghqXjK4hU83nvsjxqdsVyHC2YyGIqtY
xAxGTTTJ/LjyXN0kdUB19cmCY6RUX0FUWlgoUYUrJ0L1MI3FgztOhME/DnRXhb7w
hHB/gxg3W1bL2DyWO5mhvpwpNuSyYJ9BY3XoEkMexlpGqlIjFtvThNGeAY7ZHhy6
aIdl52rCHZ0EOzNP/uq+bahBznB7jUnWYrO3X5K5QcLqZon7vZBiDNo0O5dAzFyy
e4K1vY7NnfL8hulZYnBxp+BVB7ORUjKtBY8W5mLZ3Kjvt1NgMlo6eJjtKLUcr7ld
ZSLD50Mo9A5bYp0lqM2dcFjO0rQzLnN5Nv+ZHhQke6FGB9AXXN68cPAeVWStVs9r
I4PwoGlSIeM4ZMJuJUsZZszduyZicp3iMsjEBp131Qijj8AvQjPl3EuvFsV43biv
hxtX+xa9/Op+YfPkED1KFDeiZ7W6MPJe8EPc1bcZrMkvY7El+9J+lho5mUTnKfsX
S+unkGsGnoRkj/oejeoSvcnxq21NQmeY3d+agal2CytvOKE6H8xPrO8PcufnfEoI
1ksvwULEmAxCdFfGmqkkZqFxUoMXxG2JnQbSEkQ2Q3OSL5bTJ2pmlXMtoY2nua8k
QhOeranf/bMChcQ8NEG1kwIxTZV6U6b3CvhBkxl+MU6bZweq4y4IVuCIZC77rLG/
QLv4yzZHHMqLKMD5wQOpeuIl99JMbThQb/XJjpEyZ7dOr5RXYFyhwr3qAnjJZQyo
l0nTqBCsigdYejixOdlH1XFn5wJ2/ojclOxw6E6Rfpt29Y3EtNHBJxLV9sw/kyGH
it/Kd2SgzKOfWmAc8s1AasigsHVikA7fX8+VOiz8CBjyyjkLYbTYH2y0MNcqg4xF
4iwksLOFFIEAXQ0+oFWPl/tQ+WH31O4PI4HU3PJow1wtbYWLS4egcSIjwK7PJntw
ngIX7XtF1KNoDlsTJu4gLxem2VB9xHiTz5mnpGs1+n3m1zB+kSYPz0KJtx9rHEQU
2VKOXGjAu0Y1EfzUgfzrImjfjSC7Em0PxQ6u5ArD9KtPpr8neI/DpC1wXx267Oga
4mslPlMZRa+H+AI/tgN/BUVdD+JM2heBqDpkLPIooLDpJPTs8eYAyF7qzUEDyJnA
6+hoEgn3rLx7+yxYGuF4sFCdaZJCOCwVt+gWbltZn/TIc93PX/HQJOTfJsBJGJ/Q
C/T/OQIggUSxUYpkWqv8swpRXU3ZxM6XqdXRukf/4mvnA0KTPjn4Mrv/ATrbseGI
cq6rujpCxDmWg8Z3NCoolO6epxYtrZzVTWDHVoOPRsZJ7/L0b+2ld8LG0P+j1JYf
K0irfIoPlCGuEafIeSVmqhR0sgUciFcOUzQllx88ZFMhQUnihQHF0eAy9dLJ2K+w
UFTtCHbrYs4pUoYM6MBak4DFiGv9UOc7QOx13yZqINomNWioYA9KGEjQII+VYwQ7
2f17N0rJTv131u48PJPBGi1Mfgosk2AoKn26lzqEBcuYNuuLG4S4mtnWT6HwprFE
EW6zfJu7gjZByRDAlUFj8K49O9KwVcyDYmd8XCe3o4gSiJGNZoQwTSzDrdR6ErGP
m9vu2jEPPb12mcHEGUBawcq+ebtcg7v8PH5a/5xxTApEeBqlFf50ZVL98c9KP3gG
Omjb4wpqlKOr2jpc83dqAmB/hZApC9SyXdD9XjL4Hukt+vXSsUkAjIr+xPIUs7Nk
TMTBRUDwCkxXWo9xv/717my6dJiq6M7B9aMrbSpwwyxKGqJTcb6MA0XapwjKspBB
l8z7Di5RL7YJQ22uGhwagotnjGKlPgbc+G2A9Qcrwu3QrOYzFJNsXJXQr2e9tzcG
Wp34slnCap5Kx0sqKBpKJ9LKFVFej3No7kkP9dg5wiv2TzUnDiHRQ7RocL/hp4dc
50n+7/r5DQt7/ioJqBHXXhuwp17AgGsztkLU2zEwGTAbOTqHeup2EFZM8/Zba0lM
/5TQYwQs/Dc9u/Ua3gSaQUh2oOqz0zGuzzkk6EV+dWUUIgWhDtqfiX+LHdigbjbR
BA+JoSl6MsgQOYa17qStCXAEizVn8dCTeyerbjrKHgwY+oWKG00l6xjS9980lhkm
qg3Je8gTEB0mIZYvQk7IjQeWgmlDR6p6wmUpXJUtHMZ6gI7yiWDxicSPTUj9TfZS
Rl09pG7yB+a2bRxkNLePohcAdlTzXGNsAz+APVjpq0QHsC8TYCDeIAWyNH+WjJxb
Bm6EM4Bpp7Z4CN0mREfGr7ZEQKuYGt//F8V7y7xIllMRPXny5SYtxbA+YbWLCGWI
og4EvpdP3aLihDlH0doxOLOMQrLhjwDXFYtc5kpgT7sg3Bz/NKqywz59WXj03IvJ
UiyzQ5kk6QGKAHSF8uV1ZqZSheC6WcVDCh+MPkMBhhBfXrNXaBhWSXCjpsi672sA
61kRpn3RzYSJc9QtJl4923MUeehSe8PEBCzI06SGd2PR3OvrzVFB/xALQ6KmYKRD
4G4G7YKrBa/EEkEftarEji+GZnGa2DuDSozDoMAP6K3Z5wqlbcPaS6u38v94U2yN
UAg0/TY8Z4ei12iLBeA9fx3M16LuTyzVAMkhsvO006mcimUqf0ECMCosThRwSxTg
Kbd104HiPEG4ezhdVECLH5mqBZ7aeudnvx+/usohSpn/C/zbmSI4vlhdDFOTIdJq
QkvBtIXe2yGeQ9c7j8VM2YCgr8YU83c5WSoITMzKRJzud7mwgASgLash6nsgKEMd
JiyofhBRDtuhlrF0eqT2x1ea8esTiYy0l5yMpSESPk+FQGvldqPSJVxKSHC6U2zg
r9Su2risGwx4daAyvjhI1Aqxn9eMSUF1ratH8uJcxg5psFIdGoenvPiAtcJrHEBr
yvaLijexXGLxzyn7Ab3V5J5TqziLTCVwAg4/iNgnk0n/ATyy4f2de63gec89Y+ld
9ATmq8GNx5i1wyVXOcHXb2wBuen7RB7vUgKo0TRJL9kG6fVcQ3GWKCwywGTdBrTc
MZth2gBgLLOBiWH1PwCn2/2ie2ORi6jIMeQiYEwnh+R159AtBO6jAsfhtSvY8t3T
yAyBRLakG2RSE+8jrPzkWmnlY2HiJNFtNerN3xtsu3H7bDrTFCqYhAQTn4lFrSaP
vyy9QGKc4hCD5Y0qTMY7UWC2u0M6RD8Z0PRcQkpOUg9ihU7HOXlwCoGAIV1qQ4kP
/Y1tDUKdfSdVI+HTK3T4Yq9T8lKr/vqZ/Fb8S6SYf5uVhj3s+dqDq4nizV/o8TFX
FgqMBuyiF2lY0t9BrKtQ1DshXLVktgIqU4SN9jK5/mvumRMS75eZElYHwwbhWtZD
NZAVaHlnVy3UT8QWVdNGb5LKuQlq6JJtgnZyscuN1uMnSTMV1UKab8W44v5v9iVi
vZ0TYqBvMf8wZWSA8tz/5DPhfMNpw1f2uS8EMYQODVIaFvIjMM6vL0yE2OU+EEK5
ntVcwpzOcScvX/fv1Eze7lXnhGTvoDDdREHvxUyUxvRpeldTzdQJM54Cn5zjeDib
DpQtBe4k0t6xu9iCtgBvf1wqFgqJRVdKDSd3rgLoyZXi/KRw1dSgH9qGWuWP5Qmo
kXBK2NWiSpSTAcoCkEqseTk4P7txDdkpC/X8N4gl6HrQjr6S3XSma7QnvLGwIS3l
Wi/mzYNaWXYz+l19chs7g/gOp8E6qR+n+I78ftk3xEX26mk+jXbUtq+bKULtifOL
4vzHUfXFISxzU11rEtPr3ZI+YlIKknPmf2xSMT9ES5qaor3THw4JVdAwY39J0Fam
5LVXzi1l5fw4Sis26JpLKqE1hpTB+QqLfVcsBrRBKmLzBD+gykC2OYgpyBHFdwYR
igqlUa/5HXeV007RBkxxIw1jzrmO8G3u6wumlp9FAAGRa9njHvdSQ+eQXBAwOilR
2er36s3L5ridwmZv1O+WMsfekDd5rxYgJdpbcZkPo4wV/Ortd57kTReMgGqA79i/
xsfByR1mHLvJ45Hlve01ipAylmGkmyWBBn7gWfIDSrevDLNpqq1DYKG9F9XQLdwe
Xp1Xcxsb1xmYXmMR2PVY1eEF3KMZsXlj5UkJ44QUSpvulv4DUssEaT+enm7lSPwd
MJaJ8SdFra+97T1LKPdniij/vThGEoGm9zlEjsNlZuGLmlHUu7rKKEgvjNE9+9Xk
5yRk/4QEb9ltXegaCAxzRp1ZTBajEscb0sFEfG6ENilxdp7TOh4K6n8IOCpiPAdK
7kuwKE2VEtBq58fq1z20YQd2cJLnf4H/gMHXiR/01MGoXrEVay2CzFRvnlpQT2hF
XBxpaBCxI9Hpj7WvY0WJyo3e7IK5auTzzTYc92A7O9mBR6okb+WtrI4LzplB6xu+
EO9dtOhgKBhuG3dCbCY9X6UsLGfvugzDq575gq58b7jS+8wlCyrwrScQTJNzunV7
Me2e1jOKbN1VtmEbHQ4i6+zP/NMlbZerCcJTaBzLMm1DFMQNo5XXYjp5AIN7i5i7
hRB00bLu4w3HLRf9nas/6u9xO3vf4sCH933RQ6eDD2Z5FdOhhxo05qV6MPoGZARM
0JrHzkxAnhgypG7crdz7cIsrr0R4o51Dn8k7adscpZKPDBk2YUj8Yy8zB+9QgXqo
uiUBoIdmW+lsrn3Uc2OjcAAcoiW22N98vtJ/a2s35KOmuDMKzLNvU8TVRTb8zfT5
8C/e8PpQ5j47GfzmfXOY9xXnI75QFdD/8fDxLo39ZKqTi/EY1S2n7LcWZ54ryJ5L
VlAI4Zzrb8XAGnjQF8Vdj/O7REQCUNu7CEizRHpbBa5t5PGC+rdIbYlUeC/eInCC
LrOl7d5jw8+6GOP0PYs5TS6sjUjukPXMUpoGsS7Mu/+m8SHNbnFcDLdQFjMZ1O3D
2yKm0RhVyA106QnsqByB7VqYsJ+nAMPTP7aIK2bxyGL7O/9OGtM8JSzvC+w6ffhh
9ehm3l0ElqppHkm7S3q7x4/csECx1zUBxDzaz7bwb9SGCNXKY+5ePJ57T4WEZhnO
Rh6d3nG81fZakRzL/p/Nstf2f4WoS0VB/en4WOJfDzEwY1rqUAnxsqeOSfec77Mz
ZI1DraseChCwABGlwtI8eo/fvQqb+S1NWdUdNzcruX9F9h1NBbiVaYd/sgoaBdWt
NaaE14GUTZeaaVE2I1lMzcQpcvwvY1yo9YeR/mfy12Ok+VdFF4qT8o4C21JVE9qf
TCP3yuq7aohWegJLOhqT9XBdMsDYY0TcxN5EEg3rLRjPcgdcJ1vegGuLpBT4yXTK
4C9YM17sBV3evMF6hSxnzUEmWABSM+tl7NG5Yy+22hdVt7tS9tma/wrxRxo2Fzey
EdOAWzgrvlq4q1Gfu9WwnoWnpolCjDda+jbNvf/KbrMwWI1RkfBBd8loo+ZUgI9H
GSOT8+JxHqWLI5a67zNkavSEZw7qOssm/bEdU2ApZMyRjvMnDR/SJiI+N3sSlwXb
VXY24HS51h+AjUqdP2bF3p6LOesh67+oSMa9iolbvcPAYZ4sp0l4fI6x5Cgxyo3a
39ZUVR2ldwhBx9jFCzD3UoXbhCbbynYGbBAxax961EIrRFJJDbyOhc8L5e2uxW+P
W7tX/P/OaxoI4K0k+YYF4hzTBUZxL8PmQbTgLtz5mvb0lBWiZHPVp2jPoyymWOoB
ookCBEmCfFf5K7RqP6VL059j2o3zmZzKQNKxeUNiuTXEu4pL19hJQELqQHMzmaKZ
9o/y+nixr8/8SamuWaT/V2kmjnUxZTrMNOPv04HcfKXqdIK7ZtiWfYJ6JaIFMJLG
p/oA/XSUAMJKJL0dyl+JmGVTVu4TO5J7yv2CfYlp0E8Y9U4u6gYMiJmjEqqPuIli
tSPUFIe/E18J7wL8YIMo7xMKqLkDpwx6BkVjxqcqRWzNJkaLCrJpZA6UH0g7ZH+j
N4Wz45mb6YBcLEQldfymjMU0DcJsiU5j09hYNSkkvKMvNCGCxDc2cw4dDsBFDxJZ
sD3HAWO+17EJw8pF2gnAW3jWrldjnl89uyErFSwB+bZVjPHHVw8hvE31Y5hzFAfE
hMzFwOTyCZ4u9N1DvAnf+LhXjislVwYzqAgwO5+LrxhBqkc4DhKdV/DZY9s3wRVY
+YMbbqM2ZKctDBsNvnHQBUGtgrvSwDPrTe7stDwbkDbYZvc/fix1Jwu2bFrZsQku
BZETw9BoAvfCUh6uOpSyIr1AjWnVX/Ajcc8b/SLV5io2337cOtwz6jCDCYIr3xsk
BVGoGWrSJ/wQsFI4omh0L9PMMxRAooJbq/ZPCXBWHpA/1Id2VweYws7yuGS8J/MN
c88z9+2daZc7LhjtO7FYfumjQASVsXvm5y4Q1knJg3lFhSAN5UMQUz5nTQc11Ghg
yyjGC87jXqIVUYiGOxsTuM1NbpwGbzsH5ouaeS90HCKhYHtt7KCewhJhaSfsYYIr
a2ArUPlEUqRoMIHoxbNs8tTtOxW4dy/tFzWmUAFlqgw4KntGtdqNAMrN4cR7+CTV
ixo1sq98OmntnItGZhJpsj0/4tslrUex1jKkeCVy+0hPlmm8pKgXSrtJ8pGOPXNZ
1N55unHXfgpVOZtv+Y4OKkzDm5Vu41FBRrFUlM+QwPg9VdZ9jKC/Kp/yZZojst3j
yyGv6qiA/y99sAh/QthYh9kW99Bv7kuVzN2IRQtxMhiPLtWx+VqsWidcyJOhFpjf
br5+PracMIVRr839TWg32xKRZ9SHB92z1Kbj8bCrkOotJvbzgL5l2bp2fMhWfwmu
3Z17W8ifPJySX7Lh7oOI7N1IFWYCzVboOpkfDeGISoQuAD+Qic7wGe3eqKRni76s
MSAMttNmskGULIPiS88UMYBg6uiZxhj7bQ9W1raEZ3BmjpCX7/fPf47b2rERQY8H
kqp2xpfkOeG2MXG/wKYBLnBc1wiVp9tRgWnt4nzgJtrvXI9cHxbz0GxmIABlSKe2
ajBEXnoGceS5U916eH7KdeETFRNK25xY3jMi4RolKBtuE2fB+OJ+k3i1ayMBMpew
Wy7Es+2rquCKJqHzjq3XyjNZ95Qq/7Pf/EI2JzK8PiwvHHX1FhaDydo0Hygja/S/
OQcKsOQSzNzxSqbSuh+oHsnt82ew3LlOQUP7Cbl/eWOFd9Pf2puIvyNrbjJZuGk9
OlruEYSDkyph1+cFa7qNY5lFN05EHgvOKTBfvTVcvbgidRBtAar5bIsKYZ6l75St
nImQAP6VotKaSw7XQbhzRZcoW4JnhELryGasKzfytnrUpXE+mJW+cLROa7F17Psh
SX4T291zbVG4lv7+TA5NBp3JZRMPOKQ65GPx8FaXdEX6NnzK8uHZXVvVqeHx7KX6
IQV9nVU3A4SMfcCBHjYl11ctvYUOIj2kK01dXkHNq+mVbipvA/NaYX0DBLk9QCKn
YMpdurqwArS2tYcZrBrDUq+kX5wDnHNr8BpqXE4USg/HReKUhNLxN1wQNjCaoZvt
FAQ9uFndGnjLcMUusyNToealfDLA+FX5KRV9f1Lm5uGOl9QGP4qPTwq9esxLh/H6
XAOxorjCjpuKzj7f2A80XZFkWd27MpA8MPhF7ynYBxV2IipQT9mzY8R82tJTimpd
RHb4npTyro7zxkzYomUZb2A5lCOQlEtirPkrkMgfvFolbpObGcvWEQuZMUqO82Zd
aHp30YaEihSjdvZ5O+yfNkzkeYZyBanIRXgGBp/DQxhxzh5NO2EI6p0W+cfzs77H
lS6GMI0DEmRPRAqfSMh5u1FLP36GuYkPGU6cA6/Y4r41C0l1g0/Hy9I5CZ8G4gbK
dZmbP72Eg5HN5fwwOLL99UpvpelxrUg9WDRkDkufztEDFNr5xikVkdVBMft62RJ5
A8f9iqZD930LgQu59Zh64OvUmFPRusOfIFE1sVb+Nm/EfJMDwINMyaGB6qbh1Z3W
wP5sWE81S50Tsc5Uh/nkZnavlz4+cp8jtSjBVKmoVVkClwbu0QwiRTq8mzzDrjx9
jfN0GuL0ayx4gC5/o5tXFRGy3wdpy4RIM7/LB5bwSgJqNCmCZCI1JRD9iZLl7Xn7
hgxfOTXucNMsJCn/GTEfW779TKJax8pnA/qusY34bA3JJByaE0UF3glRQweUl9wg
2t0b3ZLYcKjA6gGvshzg/vvSZ0GTD5GfH6aBisoY6CtcPyGchMGke1o+pFC2l8wi
wbStJmNF8jcQRrITHtF7jymEvQCS84/VLTXwTVJ42Ek5e3qTb6aLkZ+Ri8OX7L4M
EBFkvnpfT9C1Da+to9IO1BuSfOmbYiQzAUEMJom0URmYW/Nu/oLfL4RICadVtkfz
PrQR4rgQA5HX0knsiUaThLN+2LB2JAg6y7pC6cSCTwPCLpCXMhN3ZBEeQsDucgGp
cy61aSTbq+yUKXdMq4gij6znp0pasflllYTi++ywyord+gg97280SlAatebS3Q+3
yTIrL6irptGaDB4ihZhOprrFD6l2QeEBs1ofDz1s3jHAD6PlnFItQndrdDTcjb8b
lQEptyF3/oC6jHPG5wXuhac68ohSlVJe/hXOdPDIdvpiQqraSgsCX5nZm1eQQBtZ
fKgHXDpfoWtfwos4jNnPmon0+8GljRxnlIigXpWXlysZAIaHNPWxlC/TYNB/qdGj
8P0CkRvDf8k8+DJNYHqRTfVb7G1RIdhrjf37jq5OSPnA0mroQlh2EyBYyTatBgHe
86HtlyhkRwwJs9jei9koTAJRgVz4/dxH1JbeABl6fNoEth4hQBhUdL+wAK5RDCJe
em7JWR/E6UpJV8psKqFEuDjHuH7QYw6KVxYgWfRiyMBx2na5Tg6bBlMLVVsmKtfH
ghofGok9dKCg8Gq5Y9FZ26TopebhjNDubrHQcvhEsm5/iT/iABZwIUeCrC2tpm3v
GC/oUdMQZDJpVSQxtkdRoUvdOX16VVk5IItwWznXAu/fIhohdoKsQk+LrnC1Uui1
1Io6iID7TjM9vM5MEZlmQCVNBj2va4QHXzj6e8OKLBDerRjum6RueN9Gkm5NFlbS
ddIxFwqzGShMuubxKJLJMHNTgnaHSc9vdd+gL6YoKOZaIxw77Q3B11JY5SPwm7Hu
ubViY3GhNK4HI0f3Y14VUuy8Ofthuj00/Rer/pr4BhsmlZcjjkiYajKeER5eAhrN
w6FF2Jz7RmB/jgq89w2rPX12k5pnPssiu3mvp2oCK+cvZt0aumr3aX0hN7pHkcaU
hGHtRWLZZewDoUTSorbtzj940pPTF/VexiHh/KUCgEB8t7jMnZJCppsTa3EA4/K5
GJS9nlh3YAM6rIfGYTUuv/MLfgrGEdkBnO0J7ZCCE9VNR7Q9P7YYdfIVrZEDaQUP
kCwfu0wJ+ZQIaF4loIlf5UEDQM4tOquSzZQEQEa/iQQWAGAI3B64/U0YdvFSgGt5
XX3nXZv+1TiUfPPpFpbAzuLYXWG/oTGwaPTIBAArNoHkip12DjHeDBqw+sXoG0QW
XdVpQDa3I06P4lbxY8/sc8Pyq8BQUAABWHh6RYKv/ml2OrJVhS4Ua3g8sCKxiB+a
lxyIKehpLxFQyv+dWO5L/t0oBL0i/4jElFRBQBnIZisUSN+QFQGFrpWgAg7HgP5u
B1Ep33Lb9wKakBEDnBiO2XEYwQcQbnzqxX6qhtVSlX+ZS5TaqO71k3RepYBF4GmQ
8L8MsOEJfeKYi9Ic4B0XfwMQPh8wIMkSTJTS1yg8TOXI8sqYiB41RBrdiBxva3M/
h+MHO+aoe7eRdLa8dLHTFnJnbZ9fHz/FhQbzwhZt6HQLHdrvXAwn2+phKNi5UPvz
Zfr5bgv1+0kQUZan7NK9aGfxQZr6EH87bBwEcYpK1KWrwQJnI18Y+IaPCoz/LNyj
bzT0ZpUmpd2jGWREOTSyRySig7VyaR5QPVcAL7IwdTAxxRmIsM+em1FaiJY+cLGR
Y0dwHW867Bt/iXbc4akfIxzGcomrDkywkpjhCZW22L1YsYZnlhXSsF+WZcilIDTn
WqqjMX1Kiu3qUt9yp8assjHlOZXfVKIEaTyPl468b4qgBNPnJyqc/Eqmda9utWrw
OJH5O3h2ZMs9u5OZ9idZKByM+vMYoEJZ3T9W+JisL9HdOVPxPFJGd/upbyRYgmnf
Fbuc0ZJKzNqi2YCxlIxBlIhopkNBtCRa026KvRnEhiKZrtcm4C+vCCvoY+Cm+ER4
/1toLBtZw7yHCcfXk8tXMxEAZYFXN5ooeW67XqItqhSZWfxfYG82TjP2BhBUhqVl
Uo5aptSwTeteZk96y3L4S4tG6M4vGHgiqSXexDvtuVVwraSi6AFBb2UM77bopGLu
xzcP2tja8M0h2HH+ePdGLg1SgTiYMAtGBJiIXhCQeFZKcFe+KR4EeyisFFMo6mur
PUq7KcuKUIruFxWTtirURhScOdFYoxWP7jQOrDCy0B2hbWQ+xzos2cOqnm32Cd2D
FmYxCloggJ2UXuQbIDSa4gZQCyDUa8yi0pV7wHX5uwGIaNYY5jMC/UofFW2vk5g8
WC+ywnS0ZMZ+nBaKhnvrJoNb8T5HjhY73A6UbhQVGspcDXCsfjL9stYL50+A6vCX
/WCLFGYurVHQ+V6cpZJ6GDQwX6ys9uJhYoRQvb6nmED9ERHu3hYrRLhFMK/jXGVA
dQ0r2B5CJ7c2slUpUTDStryM7rMYO4GrgMW2jgtAwjnri+7U48qXiooLtH6OXOtu
YQnhsap3KVmYjix3hKn4uC4CdJFkzEdsXJCMh+s3pe1yuJOffxPH8oVH0bnjHua7
xuCNhjkxtUlDCXH+6gDm71VQ4yi7Rujk4+wIjUqOaspr+LB+3G9Au+Ycj5F9zePW
o8/5qg3VYO1xiBjPHQeBLbg2vt13f72DIeclbzD5BZiwnBYBgiVKidb/uagqQ/cY
XM7SLJZ5XOFRDsgVekaaaEAAdKC5NpmtNg9xRByFUdb10WHLnBFQfD8PYXgVyxrI
ocamZ54exHlqvY6Hksc4Z/xCetrk13+UcS4HveaC8/7bQpapa4WMnlJmcQGF1nll
qAeUsmtFcYRyAte3v+xsPZDFwP0LbPn0Ks4FzTIJRSUmFBNmKhVqUxz88UNebUNi
DZ6nBx7JK4yVulR2t/cX4ptdp7vG9yEglRxEMv+ovtKpPhkHm34wZt23VYIFo2cs
40kz10KT0/v+1WfrP9x3mr7tBp26VVmrh9FBKs3dvJoO7mBKpiyPfhA2Z8yk9ybZ
rFltz6kELSxK4MiFl6VJ4L8w18kAQNdjetxtBUNQxaA8txj3fmupd0yubZkM2Gv/
A9ssm9ZeAv4CmQ0c78RBLfyBz6Y8rUm8jg6rriL/22S714ZnlWAgkg7c45Y1Fa9C
DPwpmWgCsiGL0wKJxpDf1YS6Vpt6ZxF4zHIdmbEyyuEBAAoVdHCGyoQZ4i76gaM8
og6XWepttOXd5AYiEsfhhQPf2MelKX4JwSOoOmOLyXm94kAvkJeYifwpkPDMPpsv
8ZXdJ66x5szHGgXADZKq0KQrf2qk/VRGZhl0QV+kt2TziykSiyzNAHYlT+fzRVF5
SYFk2oqmbSDPwYiN6KsvzRekq2FJdjTqmB/IUh3cwNNWPmg6EIeqofV7vB5NVgKh
lziNX1ZFbykKSlCWVcwRIAJs5RvSEKdsbR5+5TdlRCDXawuB0nyeq5cp7UvBJlys
LROUGTdIFizCG/r0uLiRx38HZeg2m9SYSbHPHPGo84M282TFlXHTUyN11FLmGcd7
4yppXxfKTVLYM5ZMt97g/Ci2eytuWGwQNsTlYlbTvH0IXTGhpq5/xXLpRWv4pvze
dhbvMiK62ramapon6c2yjOIAsExVE6A4INklYstvpinJY1Fqz92NTdktlMIdkJ3B
3nVn3UqW0y9nurk951SN/j3iGdv0D+z/96qG8Kt8czi8DOtoiYMV8zd+9lf6eK9l
ijC7Z40YF/qCK7IjKVQg963QNOnQOKn88QQV60UdHND0/iThWs2Dx+j2GfQFi5tC
uVF+O0ZxqMHT3ckKYnmD+6WJzfTFJZiceA+eiw0MrpeulGtNPJ5YK1VnLqK0eAd0
I6Rm8EpX+uJ+uMCHB7w2KBjjBdu8RA3dq6z1jxFjBViey9mr5bL0LPjNVFCaNs/4
gNG34bPaodZ5OamoFSGhcs7QUfvLSWz685jDuu8NaUwt6vBowGXdUo9GrC2OPYX0
eR7KnwnCww4ueyeqarn7WVfYmsX9CjMcOn8aqaEuTIlrdI7NdchWhmSbmeQlhHj1
llrxC/xIXWsw2fybB96E+4FrAcAmXLJ98d9Mat1Cn4xEUcA8B1fpFVK6NZlZt1MJ
Ce+voY2iLTCE6HnSXV6VKOdvqWl8SlD+NJPX8TUkkJXeEtUBz/huUXqaPF2/ZmZb
pZe/Oxe/nxgl2x2pkGyro6kmtEFkgWfuL/r521G8OuFBwuUwvUr8HYSGw/eVMbEs
wRUyu+g9x5LB0FvTSu5muOynd571jrfSqaEbhW0XK1ejb2tuIVrYACO6bg8CbMrd
cz61xEtfD5CQ75O7OEKcr6J89Z1RZa6a25LKPuh2b+SQUDcsIFhL5z1w9R9s4Mlg
wLnYDuXFUbyflcVasUqGBq0t+lu9s8iCENlT0zOmOENhpYBDXCjgMFR7cJu0awWf
UbRYrHFXcN44warXw48NIKVS6ni9UuL7QHKU8oPmFvpDpfD5Xi9XChH9BJjYQy+R
WkhD8yc5qdZ6zGuRIh4inT7/0CcNoGB9ajbxp0nPKJ8JBnLmILVSHBRBx8hgkPSL
AxuksyLiPal+QrIoaFykvcU7dE8oB1e8waOhJ3yz+zq3t/+pESM8jcLBMn1z4c9u
C/90cerBrwh3ohE91KjsVNyws8L4QBMoK6neHPkHBUIoGlFaJ8rPrxXLr6wJQEfp
DbqxEdQMh5jN3o0/JhTadQ6nA0HOIuSk9ckjWqyD8KSz8EQKKVBOcdG4HshGM3Q3
ZsMBHm+OL7Bf/hypyYclcF1Uaba3eW64PXqzvGvZvVLwBd5yz1XrDiQlVM9dAqEe
/PoY4tofWl31m2u+YwCq/BYmclajkKiYhww2gQ6Y9+Dm6JJlttDj/eI07nlS2PAU
eabd4syigVV67OpvfZG4i0Samda9wStDM7/FcDF1qrn50rkvMnIKpRG1bKYPr/oh
64Ilq/ld3BU7IieIGRU/7v5tWBq0xfzQZ927bc9cl/pAK8/HCEF9xBkCCQUp878N
P4c+sFI2+CrHHHqRQxvZDwgFkh3dCGYP0xjczmHGfIQ+VvEPhCrMZPJLdBUOSmTi
h8/nLy9MVL62sfNHhlnSF4Nkw0wZBUTaWTkNftRDKY9aQAZfilcXQGLR84/CbROc
AHItklxxZ5tKtnOI1PrDokZfSKP9NDvJH5A3C+qLVXULYrAIto3679Pq44E556Wa
jVCsQKt+eG76tgHzhLgIws7Tc+iVg6omEvSqNYmmBQ71cZFa/a0ZYno9tT8n4RdC
rXAPn8Eqflp2mI//X0GbJTPOtJZ5giJLT7dhbg+IWTWw1udvBIFaURGxKjIn7s9o
9AQJwsTQMMDuomOMIeajo2f2PDTGlD90SHeFA3ZuO99+17b3JqkQmzyufy4NfvKj
ETcbB0KON/ZTC0p0/j+CRib1kdhDhafLbjeiNH4wp7xT3Jg1sC9p0DtCHIOZr7Qa
VwCbzFK73+OsNq2/qiV2r6TFWwcU2ZJEK01lTTBAEnyA6BCBeQbFzGtuzFposYnQ
PdY7uTqE5XWr5IiueSQg8CZIGyc7tPnmSuk7Sn6kGLD6io1KDc6sIr9R3zFo0Twn
RXswxZ9yZf0jmDYManRk/ZKDE49R4QdpTt3QOW5gFW/ATK+9g2dgljAZqHx9gXdz
rK2v0e+uPZ7l2brT/tBeN3H/hja1MdSm+4Xn8s5LoHHxPYOBBBCtjCvI3jEfQzyH
Py1r4a+LtWCDpJlkNfdDijoliV5ZJ2+P7YcNewp2NmYwWVmCMEGsLmDa3YFegIln
UlH3y/ALP4KcQOiDGeVs+JYSi3kqhegy4479ciqDFfVnCIk710W/l7zyIMxxWdll
pSYZxEdyAZMT5LvEdVBcI30tiCMm1ZrKfI5fD4ol+fPvgbK2RAcvFnM7oycLjuWO
cTV/yUF0mK7je6WXwDhDLsZ3gDOZvyCvV4uKyUc+FJD0IdJ9ShaWqN44cEMuDnbu
aRiRauzK8THBtEpzG0Ju9hLHREGkiUs3gqF43pUDMv0N+8Tv2EpFFEOJB0+XSV7M
4E/Tv7NcKZRhacoEivRU38ZoAaAcSJskmkkWLBQofZ6urhuIuyDKOYfHrkJIxRXr
Yjt83vbQU4QPhI9pM4f4sR0W+OFvHgan1wKQMQY3dd3nhl9V+S6sxi99IL/4W+K7
8ll0v28xLBVqE8cHC52vemzMzAaq6j7YGuH8C3ke+GAmSUWMuZbjyjDowp9pldZG
yIYRN8oCFomuShiyJV+iVcisUAvc3KkvkOQ97LT9eZ5DCYststEOQOEYeIdtK73y
q6DwJIs7qOyOp9iWFP2wt8ThF+mgH7bJbhYyLPE6VY/dbz+zQSPOSARMzkU/gZ7v
wlZ89MAFrJ8gOgY+BwaMP9RVOXTnCybAd+NRsMYjUuFFh+miJCZkXjZQUGMTOStY
7bKILRB+XN2QR/tVsDcEVZASEEBNqJbKXttApTTopxGnWWR0hrEBGXgsTbg8OhRY
iie1GMA3xHK5qkF4yBCNDVaiUibbudgRXGoHvo88xrzv2H/bxsofTdRbz3MoD/6x
XgPOmaoJD7irM4EevY6T03pABeiWLzEaF4CpyaCq9/Pxddxh3n1g6BhAOhqmrtcx
5QE0CF4o9jJxvyMgdY4JXH92gn4vkEJ7zwBiuNnrOPoLE5eZT5vj6Jm9dSTVzqB6
pJGHkMgV5dCWo8slQWfpMu/0Lzjgq9N3/izVJTnkkC9TiQ/fNZW6/j52P7BPY08m
fQEAAcuMMX/eBwR0niGHs7iYS+NJav/k1n8fEEcKkYX0vzouihAjRTTOTE8M6VBc
8lM6jxChFyExdkmnuA212RktG34uhR2uY9kcHKm3CDOrqqCcebpuCPgrslSIl8EX
B4nIZqnK1N7hfkZbV05fSeZNjSEXBRiAuQmq7ykV+8H087F4WCk3nhMRnxWgEdgT
HY+L/GNqsDdqOf5p7LhRRk0B8MsLhhJiU7feQ6SpKXwYgEcC6fVrIGpI++smFjsb
5R6G7jp2xic3Q54KcXOxFIV8lWvenVsdNJ08G9bxUWUGE2x1XGu/N9dmTEiYy0nJ
imQiUiQ36oLITVG/AXQym0X5hKbQzvYX4hfLtoaUXezaPtWVrmTBrJdWHtcXpRfs
gCvJALcETnfyoUL0KFA/JOOwjsI/Mqnd22hDFa4o/qP5niwml98CdCKtK4lwWGUm
mB6CxnKJYtDznE524cy08TEojMK7OHiST7wmUL/HRUcDx1V8A4XVqbHN6LSqM+it
cll5pijnxhiwLJfvSU0LP81UILjy8WgvgsuySdtY+5L34OktPQcIXxKVjYdwBkJ+
myCEP0boWwPpydNJkAOS4UMfq/J7jLOt7khA4MoT8Of1VMFmkdUDph+ZOeVaxacm
f+YAm94Y7/UweOqXoCgQDrVw33XJq5+CavEkGuhCkYKGlxW1Q4df1nPd3pQj2e5X
eStXtHnQnYWr4QZZv12mCEXw+0Z7kdFw4x31tAmEb5AcePXLArqB+7iKGxF353Qv
DQTM55LuuNBk/tkpmxvOFFgV9AlE37DRB2Lie/rnVi4tf1vWuf783bycJ5uSKJwP
+sGfXPXLEYvoJBVDkKhL2xjpsFeaSk0GV76WJA75IpJuQpvlyjHMpIh31hKSQUcC
rxLcjYr/AMY4EfAQX4xJXs4ESa6fScefMm2sd3bz+X8Nl7HaFX2QIYk/9w6Doz5f
tNb7+GM+nDo2flzu/He2NB62UPYxuqeRKs01/8wV8UJzPNHEA0ClYbEsCogW3svK
bzKIQjXex2siPEVMaapoIQgJpp9fM7L/E8oUkZZ6aSWu834mgRfs3k0AyiBpEcD2
8lHTEAyNE+5CxHVF7ou+hNL3YvqK80BTtk39ahcwwO56vaRDOMXBFVeD8GqPpfvs
vyWXFlVjWVCs4cUG/iE2/a4wW9tOKyDRwBerDXQfmKAhnpQhjo5wxZMOz8tiH0Ls
D/9s7w7omt83sYxAXrZt/vB7jJy22cF8gcnUPwBm7qTbIjvOb6CjPLEC/cnFS4UW
pXThUvVeZBzhyFYYByTbuQZdWrPHXaPpm0d1c3Sg5OCNcXEeZ/JsgJpfq/d7EHV4
1T96msToBrfxrLU42gh3CBBtrc4vVRzq8pSTNe0lCM0ZTfogivGs/viaOBcGwUhf
DZKSjolaRXiAzTkwDZb9mPYyklgWFNpVtsHNtCviA+k7fuLi0JRyIy35oX9DjgUF
dins5q2+TjoWsE8v79+2s2xypaBuSA3db4bYKgw6152RvQ2+vw3nr/dLvPaMNkkU
9OGIdQM9UJDBprIJ0g1+5ZRrv4fgF5UTivn10Z9GkS/bCoiUoiwvajyfzW3bSwAf
zKgzxYfPcVWcnkR2PSo/yDPerIEfjyBR9DqkSAoy2wplWCzqJGrCkLG0tXnVItoe
ZeMRClSLfEvadl5aR2qKEQNhY+rqWRHOdfrtSqMdbIYyioYzCfDKfMjy2W92l3O2
MiN1DDdz6g2nIYjGBOyY05UmezkiWX8tGsBwuyNl6jsHO83k3PafrCrg81jyUTPF
3jnVPTHt2j9ry6YAZo6bOZt7W9g3wNPZn/S0/3X32tgXfT3QbkpTyyYYfiRYRNlk
sIWT5Y8diOXp53S4FVi/UMXv/SRZ3dYKCJEgxB6vSHP79Vach6Qy+zba094b83p8
XJVd9IqEJ1JSJqw1XEigiVRc7okBvRCSrI/hdHRQBlruSjvK9Rg3sM+aQra9tpTd
kpFHG8Hc9yj+21n+2UMhBlsCV9TMvkOshzSqHQ4QVEhl8jc3L5VGFo3XbXEeMJ2/
ZVGbCEHdPbZeQw7r/GFi5mTnvMAmNX1q3CXO3rwV01hFqS1qhG0HdO+ctC74GelU
ASoLZQF8hF9pqEtAZpPx2FzVd6LHWpa6yf+pFDLYGf5eVSNDISOLnySOj11Gq4WN
ekF/Hw8Wdby+Vdoww14vwE8+9zMvI5qvbH41u+Rx4JmTtWNs3GnQe+8pJJqX3Xfi
9/zGYX85UOxIw4bMEHtFEVkh01AMpzB5B/vCBdKbKYq0Qs9WU/plPJ5G96QulXFL
rNIXW59OChBJsV1OEjd+n7UWfoXcHk/1JHdF+dTCK7RoyTlNlEVdnayhF2BjZQHI
7l44ioQGIwxAbT3UEk8W8dfqUFlrWTZIimwlW5JvEwSdrCrZuQMjkKV9tAuPIaVY
xrtHfU+kasXL+xSU845/a+jYC2aVcRY822wPQtsSgrh8YzamyM3DJPYYAJFx+0QR
6ryIZp7QW27u0HGW5dFB+/vQboUoI4jI85KXGEmxD4nRyW2NHh9pSrmt9oXclt7S
yAsKzgL3CXsx5yVBA+bitsWgIaDLqsicskf7wGu5dw+bxL+iWgPoVU8IrvO/iZVw
xdn8tDVfhdVaJyTOinEWEHVMySxvsGnkwD8PekHEqrXgbRrOGFyiGk829hatXfAE
SvSawjvZl3XCc5BQaULiSpWa/ejfAff66fsHVlPMLZMYmqhSGsHBh3aaavb4UEH5
QGMHEFkvQs2iWwaIihKUOzr43qgZVTmrp3qG2JE4M2sgXhb2twOENKiBgjNHAVe7
wUQm5vN4uJWedeyzPJtWrOMIzntQBTDLnyUh7eHrSNmpCYyPL2srcR8pzN9tBCBP
pdaKWKewhCtKiiRHNrxArtiseXT0masK6CIwdmIViWrWZMLUNrDkbMJgssETNJhO
h9vh9XiNysYAVoj+2K/iu876oCd7SUhk7SVy+tjoN5VQQbqTY02E50fUAREGp5Pq
9IV8bGijj219FPuiRk61qhDOU4GDc0AJsJxGYxQLKbX27C72zCW1ZEXbSwBoeXRM
ELRzpEm1r34+fusPDPXFaUNGc+4eSvbpRzMpmyU9JmDVja0Wi/y/TLbSBTPazZ+2
bhaYyz4psD19c7Ca48IB7tzSoUd6fEZ+3XBJOk3rL7KWhIg8f+J+sor7iaFBNspd
a12lAZpItXeiTUX1fbTKzmTVLb/KRQdu3MfyP5xd+CjIcfmKjZ8eQpPmdUFEFs+a
+wr/iYDaPIeXcKGeowXGeRxWBGYpApHn+dG5rxLgYTn3zn0ocs2I9w0gtB4juGgh
Mto4DZLcb6lY8RfnK7uU4MJIL/lho19Xg+idn1jbRk7PjTlqPyOWv0QglMnSE+bW
FvAvt9AKrceXEooe0B379A1CkL0BgD2dUme2yJcF4MwiWfraPB2NUMjZNSKQUp9+
Rm+GBsBKN1BEbcssmwEo22lJBbmnJPQ8XTdJ7VmV0sdECWR0Ll4hnEGu7mLpuz1P
/dKAQwlpbZyhxr9+sCDlW3bsYYkRKDIfvLU9qMWOOkHaoqsiIf2GfSRRt/RPnNyE
G5rchiaiGH9VRmn1q5b6/3jCbci6Av4a7HMsoZyJ3tFTh+5Pie1MZ5PxyHUKpuHH
Uhn396pqih//C6cIZhdGaHVOnln/SULBOvYiUB/ZQ5g7tSgLeWrXKQwzupEkpx4h
izJPydzJarQ/M/8zT0jN52h9si3j/O+5ekFJ037V5dZL3QtkbBkcz2pile7BUw2L
miYH+TGKdxdr68KtBy0tUnq9dH4XBmerlpsyggHA3YGvLuMXL1S786mou8F/fjea
gdeI7Q3sYwJVd40L63A/712UuCNQYWglbSGlvSTG31IBQaHbgjISIVwFTyrGVUI4
4WOBJX6oa1TUMm+iv5B8xMlIFE3MRXaICgUBQmLfyfWLs8wU/E1qZH96S4J09La7
LpECS9d1bIFbeaG1rwoCZuhRt3VltlyMG6jnxI7Idc5m+dPnBQ1o4zHtZ/FujvEX
D7mXCm6ATTsohocoUHw3CkLoAjZfO60DxrZUiblxGvrM2u3P/drTpOfUyUastYxF
rqDLW2/btE+5Y1En3zpaPfzVxnl0UHqnJqMiQ4Uovdhy79hzjfWBzOSc5Ii0Ac4z
k52XQAsAIkHZMOcdiK+UqV8cj8qwv8LX4z8iYjMVfYu7cgaHm6Nvgf0M4Vr2lFZx
r0bou9F72Kytnm2oK/xgIXZSMvdhMUEn88t0+FWV9nfTP0iRXQsFJzrtNhi8IYta
TAVnSQ6D3FT3UAJkMkTqE+boPjabtlpG1zrJD/OKyEYlpYDnEWYv5c461Zz8ORac
K3wUJkSfaJhGDaSjB60fzr4ca8uP2+h9djDaqgMc7ykrROqSKICRuD82p7dELs71
ohrC5/+UXazTzY0v46R1URxBBs11qP4EROCQnd5NmnUzrokaTwBnRtcnqKFsafTE
hhslzAwHbvMrv6fBybs198pclLUIHS9aYpEg/U9pdXGbfTcJBJiJJtwUSP7protz
WPJFN22efRpmctbeQYW6kXs9g2unqVYFpLOE96kf4bdomGyPuIvLezezrQTDBtR1
esf3c4foue8bgdjbGsgHoeuKqouqGyGCKv8u9RxkY5mOKXkOUl3HPp0T6vhQ/wE2
lxSYS0OO/7/YhQffCZ3WOlKoY6ttnrSnc9VyADBMJe/Ix7winFbWdv3mwdBJS7Pn
9kOtbP/M5BSUL2Sd8X1wmG0FkcfUohXUhioAiiSWx5iKeWOpWs8yOI4NmRdlSojQ
z8fdDLbrPk5JLFx3Gk4f5oyCsflxjbJt48n6h5MirMtx8DlvOD1JCcY9WKiBPajL
U7VEeD3iLUX2PpJe5S0ZbZJ0G0BT4vvGR6iEzcCW4oGegm4HXdjp5HJ7XwYmrOlR
vSB2P2+h4fpzTvUi+0OAkxJru83PhEKXiDfjPZf9SOx+cFvqten5UEhi0rQbPdx+
/iVn1uTpGsu0//eU3v1TpNaXCmi/WSfoEwjAiW/o+l8UUZhktjzoM4vqSzPuUV2o
1lFKKvSo1754NWFDnn+QagWySX6nozOu5CQRyaof5wHbsv8QlFYV2X11BfD13Bja
lwmY3+jfmYJJN67ujAGP0sxot4vtzrpn1nIboYanXJL5XbjekGi5YtjRKvCtNlCA
vU/6M+FS9DvqgfmSHVXqapM0RcVMjX1x+iWZvRu63h15fQ7PtV8v88h7FjcYwUfW
GvXJZb2NF/HVwx1YkcSBwthUpOMbEYrWswPfzugo/ikA2QvuSs92gynuAZP8sKZb
BVG/5LPACFKdT1vtsn8tp3mm/nza5XInnoc6YhuDihhvSEV78KfUjhcteJ75gB5d
9IBlLv37qUoB7NOveGqW/ri20q9OUmysRXJf0nJ3isCRaBk1ztA32t5gDe1RmUbp
PQdxz947A8l2QQcy5kPfzx2+SzOu80YTD9fmGGGdUozhFE4l3V5uvXi9zmV6Lcy3
/7+ac6NrB5wSehsnXAEMLhH7gC99Xb74Mz8jgzf1G7O4ED2ESWr2S7NAzuGEeZOJ
Tr2wwiQlbuR+taABmONkVykwz7dnGKrGjZlhuiQs6/KB67mK3byXs6Z695YhYOOI
08u/GqgngWhzpgu7nhpqpOT+cewYUTsqQ4hxvDkgB8nMbrB9GRVUykL0x/KNaM7c
IsxUiagXQeTqmO54+mnhnxxTklYYllGYbRMP5uLgHZfoFnEExzHZga32eMvNrclV
WS0XHg+vWZWVduaH70RNGxJW4jaWRkH3j/FDbePr0RTRTi1dhHFvwI/dqSPlVds0
+4eKcZohBaNtFAzLXmY3QxfA4jcIxg9AgZqpjfaSC1gPoQTbx8UTZIECa44nfyol
7iezQBHeINBVYwwJDMU4CEZhSnzoEnvO7qa3T3lSQEFf9AW7E96dwRo7j3ckINSV
beAvkQiaPqE9ojD5fnQlpFrrsf3WYZJ0lmoexCCXFW+eEKtRqoCxIXe6O2EirSsq
SdQlOhwSHkfpH8XEfVPB0y7EuZC3wYjxsBiEcU8Xf6I+8jp/WWlmUegVLa7oU7u+
w9fbGmDBUPvw9gVYlPhH7sLCON8MX0ugIg5fHruVw4dHS6NMPVDcxjEKT2lK+Csd
9Z9HnSDB2YOT9wLZoDfamoIIYQHeOH+303DUgCl2yOZA5W+pUBhf7kySL3jhBEcM
2yuMaDGfKObNBgCyUtVsisWmsfX6nXjhgaz1/6MAEi1lur0F8I5qQ8gFMV4g8FP7
X6cEPFk1ItjL1gSAxIDmehnHmv0CehO+iv3zKCw1w013dR6/MF1ftWjjjFq2FPXq
TftOzrWKKpKFc6Bmcyl2pfNrPcpFL9ksGgE2rLVuNnGsPuy9ZbE325fhJ6i8j7Ah
QxMEkmOCzMRneVJRncbBWaGVOXsUmcrKZWbdrMjCKiwYc2jJHMC4cmyHY4T6lMRD
I2H5Wl5zVekm4fmcgDwfyKro0l/CYLZsEbCOm//EYsTLaP0lS2BrXHN4CGS/ksH4
AsQXQUrSyXPokPvTPYIWyRVvR1754AouN5ZAHhk4WHO1RJqaaqX+R9QgXrCe+/Xr
zgsXEP83Z5mURUKF9VG5rwsY4fkeBFzgGa/ERB5PmYabpr790TaT0nMex/t/gOZe
8c+JPfMrBjq/UpOlrFLMLzK/7Y6zOxj+/WMp9gBhSe9TDW4Rfg9HSbYeOPekbjLB
eMP0NyukZTg3gpOT8wWFJw1fLrJDOoaEmCRY/Ra2pR81VQrxFPfY8uP2RyqPxJja
om8NKTB1PYJS05M218J1wT5yqzpxE81KKIG6nwX6D1kIgcoOcSkoE5vQLokEr1PQ
p8QRCU/1Vlh4Y+oywD5HwN5wU4xp4N9A44ALRqE7oUy9RZe2EIpTCycLl6VX7sdC
gOjyTUP59iWHyJfuWqJRT7qGdHeQgfrfKFGBsqGPQ2UDW8ra4r/Q78DkYmutOjQD
1OXs4oAxj0h8u+AaoYoW20QTxMP808EdnE2XnCfaL2BtXjcWEXZzbmOlGp2N2x4j
0QsLzj6e7Ab5htPOpCuoH5lpTYjZCkOBhDqpViITmChT+CQhOfFeba5rbP1m6poX
zb14fx5cST4nvWuOgs8T3HygSywU/3E57qDTcyZOwzTOnfKLhzCpVG8FJfOTnb93
JgUuEC2+6WfpVdwSIQdXwjDIYDCiQ6vvzoC5lIXm0cEbLzrxQOkVJSguf+awTXFG
lelFFU8p29Khh43aUDubDbCcQDgBh/TWescP87VfPVuRL2ufeDEXIilc2u/iOyda
kWVnc+XPyx6Amuom6mdMBOLaWm/zxoi9w3Ge9YM+Xk2bs9Q1Cy41uvpWanPkk4Ms
je5G5Dck34U8vK29ax//8yMJvj072w78BnuXTxzMOTpeWq6WhbRoAQHo2Z8xL5R2
XRcNCEa+YJXPrrX0PpXA7wjdE7h874jNToEzqSofT/gc+ZLSSyNjNSxjJNBv/EKX
W/Ee8VukyD7R86rQxJ1+Z+xCjbWFOEB5NE/pS80FXEnx83otKiSYtM6hkLQJ3/Cl
C13qNQQFwWpMW83QNpBAmvMHHfbwQf3k8JDt8518I6MShy1zAnm44HFnnWXN0Z/d
+zLsQY2Apra1IWA1OpAJ5GBMDEfPX1TyQKoh9MQZpKqESwBwJJZ3FkufXK1hDo5Z
aD9S2TZvpu1potXM+pLJAd2/ZAH16pwkr0PCDaK7yX9I0VaQpw3fzV0/frsNoUSZ
BPhmLhtZMNyGwgpYfgEivvpcDRPJhLUK/uBytly3Osw9ZKzcmSwL5ecSpGS/US1s
dqkhpAW9iPIoT+4OBjjNEtcsUxTVFFONFd/Q9N9ikie5PXJ5Ch8S+6PkXMtRvxB0
AjrbnTzbg/l2iEe17gAexI2+Jcgdaia2KWSlGxWjMymjpmFpkLSBesUaRQaxmRoN
4maJ/rBsUkWVcJ/0kliH2oZXIt3nCrLfH46OrC/886a6GZihhwZBThkam1chXdko
4MH0omWG4/UdIVULFNszakgqwoJ4kX3WT6EvPhAfCPL4TW5pSocjfxpzc8t6m1rP
IN/98dywXdm4z/Mp3z9NeuQSsrXmqsmNt7wPNzmyurtEsJwqrC12FOvdPsz7t047
q9NTUeyzlvDOpyHjOhluePcMSthg6ifUMSzczASWXA6TuCZh6ZTNq3EIjZOk12jG
W2SKq5GhSgUyHia6ACdavT+iyLLB8gXG8BbF5bjsIP784o0M/4K1VNILdANahKdn
vEfxlUvfYH7HlqZ9z73qwqtx1ydaHZzeDtfUEHLtqMqPrxsJ7RJEGVWicaBlCwNw
grFJgBwCLOPGlnycaGnC3gc1WHOMag7/3aAdi2gyvr8roaDsKTKdZudfela1E0cC
BSf3ahN9KnegsZzRKOA+D4Rz2mJssW3NxuBmV7vbODaOmn1jk6yzRJrT5gnjRShi
WA9ywQtS0D99Tut4Z2ol1Rm1SyIC/BL7jfSEiy2wXePO4A6UVmSSwZLXDAPsHlad
LnRzZ9Hwpb3oacx8acTrbCW7TKHmQ539IMggx5dJOa92ZFfkoc8GdftWgb0geWZU
mWXxwbI5Q8wRhJB4LXDZ4nl730l629qmJD+kYgSsEigjsntDxvLUB04l6tcDW/ZI
goOn852s+78iE7+MYNRj6jpCMht3uQJa/eetFX6KDXgOh8IacJD7IwcY7GTy6aPJ
eRfOY5oZr3lLetBuG+9XQM0uW9Ga38fYlM5+359RDyxR2nP+XmPMwRutlyJmwuSh
j9hW1YSSVT9XWEmDHFzsBkYEuc3eSw8BxyUxYKLpJyFRCoErrGhwUH+ZulnRVpEL
yY/1CmQ/O912fjmhglFWOJPWwlZm5FGGiWQ+vCesbqc6wnQxA8xPaN0MohaCRC0p
SUe/JbGuGhuO67PZ6UWcbVbuDEfyPyqZo+znBK3SaZO3ZGeCcHK0BuXFVJYwaJjy
eB/f0Ao39mr4HRwbacCfa6vR0XEl1GE1kkdg2sUtvsesakVCR5I2fb6AzUKnz/pc
gOyhhC+QfgPzUnW0A0cA8Xo8ISyGExy++eCPskYcscNYGyc0d2tAWvXRMg8L4JCw
YK8GdX20jfiYGejBmVOMH5s5tuSp+092RyVVmR7pAQhyt/u34lEqnmBh6LKj/C2Z
URxlya2leBBz14nGCcmszbpPXNNrQKt+2QgMg3x/GuBEIS5vJhOjNLywdwPbBUqK
Mc+TTTy/E17UrB8//QeceacBHangZCJsiAhNGsx8B38oP+FmOsVLyynbfCf79VHU
EGV86qjLqFlNwXg8pXGiLIvvFJqLMVrFLHw0qva1ZOQ2elJHvuc5TEU/s6O+CiWD
f9YCAPJNMWtvpCnPUqjkRIdCOIRA3Vb5FDVsuOv7Wk7PqPPTHokaC1iZlGVKa2+5
wR1uN1fMGpZF9NQRjMZeTjv794+O1TCX05sx6Rj9OxDLeh8uB90zSM0ZoZR0+hNI
65shdcfxCxBFixQoeZ/JZc9KDzTR8F7TaEPioeZnAOq6w8D1ZbBkrIuiLjp22zjW
SVU5bM/Mkw7UWmW+z95UPV4IsY9wxdcu0hfZTq9n+jdszLzwm2kQ+R3k/KNk0wLF
WtnShDBLZhaKW+dgbtiKFa0itO7BvWSZK9xDKvhxrGJlGkgZg413FdrOeyNViIda
YXr4h5KaShOqf/khn2G5cD+Ppci/HNJ9Sf1i/IQQI+v4kh3qSa2pHuex3LWV+MiV
H8YICxAfXHEUe0MsCXvCg2h2D3qa+gEwoUnpquHA8Aw2PIg8VNiK0e+iRdS786Vs
jADySlxFXe4a7lXm9Fa7ioxZ2bHiNwI/rpaXXn9yw6ohA7upRKAkGLW+hJ/nWKOU
xV1JlPMQ/4X+Rs0HwZuC9vL/P4wrEUzBaL2IEQoqav4wULfIEpL1+tJeHvhIPxLg
jfbPHth8nZmIJIRBT9Q2kDe24R97/9/00IY6WlXWjV6uk8JtW2RpWnxpvoPKPasJ
cccsVQ+gmBIQxAzcgFTYzCWeV2IwJ2ar6fpGpVvxMGKtWdu2+hcBvBcCwekptVFT
HYYdEyBD6GeR7VfNL3R2p/BvFcEZ+GOKgd9wzO2WbxhCkGvFzzMHjSft8IGH2zIS
V2VtcNeAmy7avNwxz1h7ItbwsFJYyepvM51HIa+aBdZEKS4Guca6EL/xcuUkP3Ne
NDtAcsk2D+g6DYbQjr/73VVHqQXlGfb3/zqAlBFUxoHKxQ2vTBHudY0DRwWc2mjp
w2bcaIwUjiMz0/EEOkeoSalJZbP/fAw4C4D28bTkMEDiHoV4zUTzOjjB0LbieSKV
+QrYng2r6R1umz7QMNslNnuWKOTt9ZMUA6MtXTz+69x02ESi6E1ar7lCKQwMyVLn
qBokUGSNC8YiUo+yzNKNOeDrMD1ZqV0/KLaqTVwZCFsC0gjtEF7v0xz0t8HQi5Pg
C8k7g2yP1WhLguzWFVMZwXhsg8r9DGxCC0NyPueJP3FxMimvaiBzCHODMf4xMabX
lcgqsNgyw2zqcv+2p1R3/aIk853FA45L4MYHa63TnMuYVICeJOh2K4qfdulNWi+O
o1yf9deVXl3qmBDIeWwG2BYXAvbNFHS+elcn2VyIYs5FRHB1EWv9kpwC67TD+q2G
5BrB/0scp4GMavrkSczcMiGoG0URG8gKZoncPuPugWb3vZlbVno+xCE3n6DGNtOa
fj/XJij2/mB7PD57J3eEPRyNG9XhnRKbtXyH4NA8kc7R8JqR0lEqQWgrejRDcY7E
baCH2c0oEyexMasOk3iDapXvXLnxBUWLClDyLjLNmqC4sSNXYOKxSyZ+1nYI8JvK
PaS0jdREiK+3bmHmaaKQiSKH887sMkvA10Nx+BBPLCarOy5dsELKXHfJFWecRy/X
cfUKSsTWrruhVGKxoA5kINCvLnmq+jZsHOEG7TaQMJqrFv4zrzl1eXtY1R8nsYTt
1QZmqcuOMRMr+a3+6ql2tBxOTmEaNWVV03JJL6owBQeyUO0kP1SxJFAT0T55Akzz
XosAL5+ocFDDdJfXB4fkxQeVrV03G8VPbbC71A0c0a1JQZxBgeCEMj/A/7KDljM2
XjAJmHleOvFQwXvGykIUo+WRHgKQ2xvfK35ByMh0aqZXll/vYx1exfAHjfGjWg05
u79ACGv+J91I4tHM5lkgUhS5Fk90/pPxV46DzNVWBLaPC6OpJTOIIwtuolenUzg/
Q0uLugEe7aZoCAeqs4yW/EG6u7n2pqxSrUw+bAYXskFtQw/hAYEIJd5GpNpD1vsM
vvK0Rocxlba7JbYH1EIBwTZvFZrWtWCZXPNRJWNCkF5M3gnA2rrxubiMl7Z6vedc
LmuW0wLDsF2rqm/p5mR/BhLRLqVu4WbhE7tg5j14/Fng02vbmiD6lThOcwsvA6VB
gjKjyQxb3hgU/mHWmVqVM7VKggHjopyZhB2tkR6Tlzsy87b/XMUUv39EiyhR/JEY
TpSO7RonLj8E1nKao68Ej9RJj/Z3UPQWjYqxne0y9tPUnPmSHvrPhXuKLoU0mnJS
dSBUQQduKRggAd7WIvNuxIFeqif4nb0QIx+zZSxUuMGljVY5NK+lHKnbDWSljYIF
X9z9pV7R22VcycVjAP1RLCMzBudBh3KSv34vX1k6azqeLVsos7dj9v3YeVtePc1u
Pk1cr7Z+HzWIOGM+LLW7TJdsBuGwn0kzqZth41hSzTH0FeOcUAbRJkp0s16PcijK
efc6dEIDhYhP7Umwp7/Ij5QBX6NQlJMzfNE0K5wbXhQDDg+NdxNxHPhHIM8i0n4b
5RRIu1bYGc6NyOHu/hAqjd3eDcULQYbwmr8CFSQbcHRXrXwvqisNhK8xR7GzU0HJ
SZ/9N+HB2iUtVoEkBVz4QHPZ+sVCaHk8VAuiH1jQSeDhPL3II73rtXY/7YY1W8h6
muqCNCEUEJv4L5WiOhykj7YnNBGuHnE8PUG9brYGuEEWW7UbtYVP+QbXDGragiER
M6mKWatVArrTN58F6iPoLYkr0M15bDQYKzMiBF9vNwAjQkVOIS83DkDdC6EqG6+c
Wdbx6lLSHz1o3oVKSocErLvzruSGSVNtFiTvBqewjLyRTJuDvIpV0i+OtO1QpVah
z/qeZ42QneSls0jcSfVPLEP7LmsFaoxCpUu0DtnC/gV3WRUBuv4AzKpLglWG3FaY
/j2VO9FPl1eFAEr7JXRn4oKtlWmH1VdImOvNUIchmB7V8aAGGXjvkcTUIFOp0dvW
klMuKxeO1biMoenDQ6egbhFlPBHP99sz38J2ugN8sDoPcTlcg/WEA792AOF4CCpi
Ld3gL68eUcGAcxEqe7hmDJkiyavRJUZnt58vCCkvw9xHAw9w2QEKATbmD0IA2l6S
D9z/APM1Wsf9XCbqFZSA1JARYGdMf2bcwZFFnadwNmkjetezJ+1A0xduWrRJVxST
Oa6m9C5BqmrWOWLXXp5JHxNQikgSHufVtF3DiFDT4h7v8CDikOPARzn0pWZ8sTL3
4CoeK8PQdRJYdi9/YtKni0/3q8jLEYZjgFHNE+g6W5WEog7c51D5fqDw8UX0eCho
G07pxyFy3A9IBKCr/VQyfbYfNsVsKlQAWO4Tu0y4whfWTXrrpDX+Ff2mhS/D9nmW
UZ+CoO7gZm0JGl7bdcuIkGmnImcEtFGpHAle2chRERF86jUblqGPDbs6IvRWuFEK
7dzMndpsYFy/YOT6sSZUiodUgG7Bji8JT/i97BGSRWb620gzZcCXmdqPILU+00yT
1BDTi3HFSeya8pGxNy5s2Wewa2cIkkXrEpRdTd/JouTN2nlcFA+SzYrd7LMb4wYT
QyGEDquxSz6wsJMEmdv04dojsow2VklOKD4FligVaZS3HZv7S3Y4wPxFYJKUQoM1
L8DU4H4u3k1FmUgsgLg7UyU6Fm7DseemPk2SBrHsLLVSieLghUmhMe8nUJK0Q/PD
SUnI+5E57KrLvFC7w/mUkcemWpkahJhPxy4lfjFEYBZ3pxJGPZv246lfxBmAfAdS
YEZeGXLbeaxzmhiRkqod8aa0dSjPqOHCjUnAPQU4yPoWWD/tPEqXbWaseWMeXz3O
RO0JCwkgbuklOh1OcSmXEp7dpnL21Op6CGJzKUpT0/k87z7kKm/vaeqvxMSL3VAW
h0VjSWmaZRWXllktb2VW5xqOD7e0DtthbCmmhHffr6pbmxSlmmfKr7XvBypsOuPi
0ThMvasNSxf9UPupchMwp0ce4PSzbyw4Sbsdk0FiH6n0hdVob/fOUDD5APsGoPaf
p91axhR3k+qt+b2OFxqqktzrS64QOlAys2F3jreg7nMkQGnQ88m2lNZYooLBaxF/
lHC964Q3aZMgrgMp9YB4732L/mhKm0PwDmnFZJJlkel6YfFLVD/5FMoLen12IOEk
L/Ihmoeuk2mClByXRgEDgTZ05ZFyurd3AnPGg1KIFfWjI6R2A95aTDi7Hw0kVSBl
dnOloj0fZQB3YzWKaTXs58s/1p1qR9TXqeCy6gh4QUNEIZv/V+HTtR6c+ETX6VPJ
D/RCpHv5m6q3oxxJWb6UTRyH/iqbucAIDTcT3D2MrMF0/qlWXPVWboMWaSg0eB3x
9FU7YRKUSNh8OJPaTM85J7bw6pRvQ/crDG9BPUTRgkUzJzzU+rnY7c0Um76ZOMD9
SKi/YMqN2PAWvtjOHTubEE7jOYni6rbFcO/6K0UJP/c1aNRrhcUopbpmaqrcTZKS
1oS5Jt8Z3cBIqUi9NQsuezBOfuHyZV7Nr3XggkRgcH4W2NhLLnscMoZr42r9lQn/
h6tLqE34984dl94GbpdrB1LVTNDQkE1i7bcp1eMzIPCdqb+dtnq/aHVgicoAcSjP
HZYfkzcUr/JHpubA7+OrtQLttroHMMWebXZXtRenMeHuCAON/6nTkJmAk6zUtTJA
XyB1+tcvs72nVy39r1keHsQAdsL2smKDGJbTdwbRX4yikmHcfWeQdJBrpFnatR7d
PpOXLfLs4LCN7DOrjuqUmrqwg3NVirx2jiQUcVyLhigULZ4lKXyc72dnbYusliuf
vjMMDi+y6COB65HES3HOxFYdtxXK90KWrGWq+8S9tx8KxZB+ejjNg0gcyNSNWsFz
dDE/vL2cSmuy6QOFYz9nZzCSCidhX6ghwlZGVI3XY1W4r9z5Zl+R9a/H3Eymvu4I
PcmH/ilaK2z2DE7DbM5gtsLThT7RDM5eN66QWNzhI97xUmn3y0nOKlRJ0vWP+Zo3
pNMhBRKbeTZJT44fv1wRy1UPXLvXJEUvWVTXeilpGX4f8OXnUa7r03TQby97Qi/I
UwQfgSXguHn+oftmIINbveGG6rw8GmV2viCvskiEnWyzRAIrHAfX0C9vBGToAYRM
mEKKWumBWTCFKyB4iX3vfX8DdV07kWqaGqrU4iyRstNIMQQV7HQ4/wKGCjcZvu3z
ASSReKCBhhzXjQzXh4iXq0JuJlDzas2LhoxOHKTXkEWegU1yc4ojnAVBX9mwURhw
JGNApHbYctN2vRnS1jr7kRiFz8TxeiS/AzlXp7Ie7tezTSqYKW8zsAz4QYqxunTN
8/6WvQJdOkRmEtUknO07H6TL1N1XbQonQR+x7NzZ9JfMNste1BnbeyLHkDfXpOfr
/SJ15fJOq9IuNGl1lURRcbjkw7Zuc4aVeUlqgnFhpNt0ldGuiiO2SAbzYFT9OLnP
FPX7TfYs3gTYVplsewffL4a3tD7q6DWKiq6HOUWJgrigiJHKL+qg/3DKQUuWpUQR
SoHGeeuWa7wzbBag330JhsLeTb9x4tkJOmndlmvfaf5uwQOOMEhtXUpNrK01AKAz
pIC67GtHTuAF5toCwXjnLWqmaTBkUz8SYL2lQ4tu07ZzzcB2tkG4km/ZI0RuRkUn
DsY5TyIU5v1G4bFJc3WJqBhwGKVDIaJDrZ7DoQG0SxNEcmzMmSXYxLp1Tj1WGu0F
Z3omkJt9RlAMGYwpuMb0x8iq4eZJtqqwU6ID0Cd8moGuGenEbWBcRcKx4ni3O0gf
HpPvR7U7SopQk/NlwOoC3Y6TwX6mLft88UfPt6aAR/H7V3QsAWT0tEgL8XPCGp24
pkm4YHAfwb3N+kjlsGAaCh+O7hSCgJ1ShM5zOyJ7fZ554YtGZWhAx8VDjo4Vag7t
4mQkt5PS8mdqfTsyka6fOmUA47wuM8Z/qZhVcrYYyVK63iZ2cqYE7ayzvVgE9HKr
05hXWXc8AB5Qr9pXo4v2gJLKdvuH0QBN1mU6owaJsJ2fOIa89vxs7AwN8BzaeuIF
+9dKpISZv1DFGGJ2HGYcBa1PfO/H/4vblgQGhXB/NSluUSN3CZyA+7QSWNZqould
E0u+TMiUWmzQoljQ0CbIs8/S4iyclCwNv0HvChRDGuj15l09wKB0STVLxlOJiITJ
1BL/66bfcItEbIdG0VQ0xf0PU/1O0AKQl9lp3zRnWQEEWXfCazZN1T5iNYhhhUbz
TE64AOU2Ad8bLCpG4lkAAXp1wa0xsL/zlE5UfdPrxdwJ9N6c5r+/Zvd2g++QR3WA
V47GeUmNfjJBidNtTDzRcoMtR27/t+qlXkFeLOTMPyvEjAvSdmz0kAaZHcYJEmb0
nNkOd6kFIYPxCF56nwZnK0qm4wWpMbnQstQAzgN2TFGxa/S5tCa8GUv19jotm6Xz
O2jXVn4ne6vgOKlt5twc5JLavZ4u3JmoqTj3rXkycYyg6mw+6XUPrIwqT/+/7f8s
ff31OB1EPm4keayV7P47DNZ84p9GXm5GfogOkjJD/WDZjuKDNUPbUTNjAj/jijtp
5xwuW30Ag0A3T0z4R2fucnlFS1t4c/g/sdi7z3AyGYc0kf+QQklwR93urK9vQ4A8
IAP6p4ySZsvnz7jHr9xlv9LfHs4nRkADaLN60i0f86zn4Q9dPwNCsJk3GZH9Nc4K
Zcz1+hQgxBFwSKYRBj0oXQpEaZ103pLlSrBOo9249rhX520B4O2EBYwABe6itw6U
lTGiNMvcz8CmexNgH4TJ6ZKnR5KuKTS0uDgYC04Jhy9fYmk1nqjjrxXu74lT3G5I
UdMogwfz0NEDldArxMLB4fMjSSobaIKJ9wcgmN3vkFzUHYvJW9OHr8k7Y1TL7/72
0hfZ+sQUnSZdeklgWyiPEwKWO0Tak8J7MonTcdQQ03Dm+66qf2u8EthLcAf5DnrP
pRvAOpsnPYOwexIRNT13wa0j3iYDgRO8uXUkPdYZ3OxXT5wOSpd5v++436erj5Lp
pWrZCvccpaklLiE43uhndQfZAHoMf9+hISvNz4tpO5O7Z9Of8JhjrNO70Mh0BwDi
zMULlNdu6UJbIaQMwLpre2g0uAF18TA0GbzJtpJhC14mJWBP78+1qOCWJX4dQaqv
AWLqKnz/CyqLpywmDiwWxvBYSReCrB26BhKM5dIWpQm/v69+stQ6YX8D94CNnfAC
smalyzu7IocBy1cCLRn5dIKa2G5jmjZ/jvSUq4MlTFM6ufLPod8CYmMW9dHjN/JV
D/XLaNhT3kXhU2CJfuzxPotbmdjbvTlUtGJAEOHdM6JDv6Oy34JLlk+mFvupP1iY
jAx8m/GxBjiAxnzd/xDJ3EKHghYRhFVkPp01qGWfINJ3YxrzNIIDtIE+XXRM00gv
mh7M9AuOZrQcR1ZV9P6RD7rL68UxBfQe2+oN/OkBCOKeDw2UIsvvH1T+TQM5AEHq
REey1wV+V9+pmimifnUDpkxg1Ud2RMEvYMKh2t2+e1UHmv71M2wFIGFTAdFa4NAy
C7fmyE96ybENKw30nx6ezqqCZJsuah+tIPT47KdVcRfz5IIKKqKH3mWVjROWkk0T
4lPxd/IDkpe7PZvOvn+FKzlBv/LJ9BZ8Pya6xW4J1HmkR4sTNr2HXkUMmSySLgHK
DrDDYTbGzmyVUiFT59iuwOQCv20VNyUB+eBB9zlHGXtmKwyVTqA87YZ1HwZBYWRQ
pQuZyFFhqZfib21XjDQmeUlJA39uU3lThotrKF45V8Fkoa0iY5Lg/aRLTNfXn08h
G7MtZO2SnYwivKIhgsNeIbaw/9ok30fjKxCPaAksRxdsAxKGXC9h29Ujla0XEStB
5V7cPdVFXgicAYaUf39vpCazMA4EMHuaC8e12XjXmjKuVKhcPBkHED8Mi4aj5MHw
iAIkSP9Y1a9y8hZNiEs1xttz5oRVgCv2oM+4DypkRiktBQlAjwHWjs8KKaVCKiak
fqVrcprG0VWVod5Uk3SXuJVyBtThGrj4e/n3TRGr83XtitzKE6ik3uXI6IK6mgr+
m5Jiu1NgECaMOx9gvfN3u0JOdPAsL+iPPmPvrus1hUkQFu4jRUqMUMXpOdilmlty
UnTgX16Gfug3Gn45KMhxekP91rmd7KV1Ag8+ixp2mLzQ0rbdcTyV3dKIPE2ZGHBh
UzLA/PizcGSdW39ICj9NE+mdZuqyAE94mt9hUUC7DR0MSDYtasLriOYzEmTEmsyJ
82Eu3CZXTQBMwH4XrvAPmt9xIAf1npJohI8NLDihIBgxdaejKY6I0T4DyYkFxxzk
it7Xn8/7igCYC8L4ARjRXND/pLa5WvLNzfGP26+8AZovyUfsKOPiLIBKF1EkLqhe
oOEVHFlDR9dLq9h2Z44I/8FnkhET9HaGhEHiiF2HIlJ7n+uGdRF5W+frMzee0+3q
LOk0Lv/J/WbIUJbs1w7W5E14OWGntqKBeFzcAv9dr2+I1WlfHrsTlAihmNr+BzLH
HplfIWnxiQrtmF51JDmxG73b4c+UG1RTQVvs2BzS+jF7AL2WpkOvSiG670IwzGNJ
+OBna9tU75pmN/a3e5HnTL9JU8qeBZ9lnhivoDrsyC6RzPCs69fxqsh+K+M1GQ4Z
NoTry5wRzm1uZ02FYjQfMS6ZkEDoQw+yTvNaTOFzCa42L8lTGptgdy04I7J2cq9v
FLASH2f9TxPYXW4bZ/S1Nkm+M5IriSAY0B7zpRzy1orq1RJOjz3ljTc8JRkI6Z1L
LnLjJbuAXm64YFpkJd9chHl27O2FV5MC1hcSMCYa7GSDisoeFPnkhHLj7C8wcLtG
IalbypJHzG7RbGhtoUjoVRx9IadSdovR+JuXdaPWLj4F//8Y9V6u1/+IMgnwwYBi
HwOqXNjIrxUn/HwOj/ij5LyrwEW6fA6A056oIWyr+5/Pznq0e4pi6lzSbDWX2Kb5
lh9ctP5lPOyqlLZA/dzyoR3PsJaG0YZnxWNOsmGa3WHvL43TL/0Dr2dsiBl40LuT
M7+JZ5ZuZR3/gSP79MSxM0gZvzzyBWqJwDke6HuVkXciiKjdcIO7MnHUXiuTI873
UFewTOJJuSV7F10DHK1ydbuNEYIah/3hGq/YG9a+d9pQG1M4HKAh4sXTsOnikoVR
IptR+Duk58I6w1LpdOtwrazDxD0089tjTuaimeaTw7QNCRQ8tuLqyZcA/+NqurLP
iOpe9G8KfzIAnpa49K3PkUrO9oLHrsdzYyUo6ow/4RVt36diGhK8qaU7KnfJmLWq
A9hOCDZKjf6wLvd+2gomoJ8yldf/wq2F0Vji9UaDCJ5pADWX0Cf+IVyorBB5NeJw
bXLcIfqMbzb3m6K7Oi419eIICohHrgbot+HEX3WHUy5inqad7JFasmsOhJEWhvt3
WnhmU90EKZP+POubZNewXAXZvDnkn2jsXgROydxDE/LLioVUSufLkhifsjjnOibV
1/09yHwrMmCmIFoLA/MRQ73pik1fF0tk+AwHdvyIxTAHU45skTif1kqO7mcIz3Tp
BudmvTnmBD/QjDudfmGBZPVQFXa+MSw5dJXdVwPOGRm6OC9OA9z1DU0Xt4uFEdzp
FSEj8xYIEr43XRVDTeLeG/B2Od+CjUcJBwVGfsjyX4qrduIE4U1xt0mRByvyu1CT
Amn+5BCgpO6iH2QpReA64q3RgFY2ySvjv9N9c44VNCZsEPmYziLdw6OrtmSsmdv8
s37idr7nCFc4Ijzz/JNiHT1Qye99uAET0pYwkgrKHRFkZYlUqWE0tDqLDCU33zGb
ERpT55cj8rESAsSjjW1tGHKxgCbB8Fx+fWrt12xDczv9T4t59EcMLnrB5QU8ybaL
/drs87lA/PXl30C5ghZUXk8iHb4PfCQTZK/7ibjraDsc6GVfEOxjxe7DI06h2TOX
XQNX97s5tWpAJ9EG5WysweaxkoD4+aPmlEb/2XyMrS6i74g4XUXgPirx96whbmro
nRCHzIg34yIXIaXEE94TA2+HBk50kPVo8xESNJNLb/IKK0UPBYHNJ5vGNWFTHllN
8sqSnUI+1IO5qW/c7kSNTDQ2AuctZZdxbP+a9Y8iF+71OqwdS1Mf4d882/VRF4hR
reOowIFBck3Fon60c2QOq3vf+dwmVFhL1e2fXzhPQmcaJslOqqqXXJ4ntI+xN22Y
HWqgkhBu9vMcOO8+Jp8kNb+n/x43OfUFhrBne0q5eNAxQBW5gM9KGiHEKTZaAw/x
ytBLZzR+AaWPRmoeUcOvJuU7EiMII4UF5XTpcrwNAnUkU3wofuGPKU2uymtqCAkQ
mV81WSD62Qz4SklMCsD7D4haULvLgSVvfd9vcfiH3bPyYDTIdbLzgbiotcJSN1zU
u7OYiRY+vY9ZjNGIuwosvaMPhJqzpG3lTh0L/62gXb+JGKZVj/0vNSz/IIHhDzCw
zBZMVsWJ/IDGu6W9UMu6+ao+7YoUNnvSVTlm6B5HjbcP+xmtgPLWxGwwuOHta98E
4gzbSErVFTLHcimK9QtgWBruEvB1M+VEgXJxn9P6eU53WJyNxswt9M5/r+1jpVtW
Geyct0OdmuFmplw9TAxWZSspO+RbU7sD8RDReqb/PkZIKTuKqliYm1CJr3GZ4cB4
2aBtV/Z6mS7Nw8YUpCESyOnzAy/2XiiE4tjiNXu7aQlZqStCZmYYQho4NI6OsUF0
lS9NtKAABNaN3oeQKwDAi4hQ+as9Hel5QkRs7hlz0U6iFDd5g+8EIqFga6IvzxRw
fTSGACJKsKDpz+BsGjGETB6GLloO/mJtoF01ZBVSxBJrkcheh5zYfvmYZIOQjV62
Skcj6qN/1DFHp0CHKuO6ua6LFr9huxdkJ8W6MGj9yMYkA/b2OYnzxfnyO/q3K4wJ
qNtzSvAjWLyYf1IfJKwmBzM9G/twXJ1pIF1VK3uan4G8sngFYGTh+Y7KgN0MjZ+a
OPfS563vctrQzbeY23Hy+E+29HResJ2OQHZhNuZCFoYoVDAKM0ekWXx6T/LZ5CeY
mXDzhh3XuyWTvpb34bLPfnL7L8xMXa+O+4Dx8gNdyDGYg8cA/VkLSfe01pSnamdZ
BX3+LZFMVrvCyHoi6YBMRwKfh1dZvwyGFVWXfKD944Yj1kZ5480VcIcU0eCiQqMM
YavMVtkqpD8g4ze3+jfBbEo0W2fN8a4R4coSKEOIsMG3ThsYnZ9yht5Lc1WAQ3yF
q/R0qm4syUHq8nf9w7hK4HUuZXNzV4pszXkjH/tU1gd7JDAQlcWf1WWDiFsBwQoh
lb4Y1Z4UPqx3Vxa5I2GkEMHfrtqyc8XAI9cDSjl5oCy5cCnLkNzbejFgR87Z6/qW
0FK1TXkt38nTI5IqS17fH/wD0nVQ/9bWAeSyzBmtvU1uIRXc2Q+XF013vQQLqehC
4lwDgy6/8tK5cBGoekTF0VT3GNsx/e8/NeQ/CUSiF9cvJ3OjQ5J07BrF4v5AIR9e
Lqg2yMUWLaFUC5+1g5LcTsh/UHQfYgBb18c+C/UszyhiV/5aynY37ZGCjva26FJi
FhEQKoATwoUptiv87vUzRBJjJxPB7P6d6jFcG9X8DDZ5p7kAGfs+4N0fG8E2HK3+
cVWSnuXKbfxD8UaiH+V8EpDDPsCZ48cxjEqkc4vDrh1Hq+CUwtW0N7Rb3xNOwPFo
EeKdtrG4YFqxfUPOi/eW2n0GBbWyzYsRK4Ojc0o96F0llux3rGIQTwX7LUMEWw17
YZJyqInWl+BEBRZk0QWgckBOioQMYwIKr+RNdDY3oZwtnA3PGIN4K9h6aYadRUp+
9wmYRuHsAZIotGdA0r4+vQdkS+9t6zSHOJ+rj2PQSyTwPvUJMtR6duEf8NZ9NjRq
2VmEdottDscNg0w5a00LCFEbSexH6jFAOF1nwH4P3p3sElUUBuomazwYRa2zTalV
gAvZ1qPOr2G4bIk28MrasKw/ajgNCZcHmNlKw7IhjfqmMWK2Dr3sDYlXsJjI5kAL
NdI5RU15UxZQYb88mo+z1a+y9EHMLs6YlejPGAtbt1OPjsDkmaej7bFzvtlwKW9c
gok0fvL3D2i8BMqA5naSTp39CUzZ+uYZP0rm/d2kvWWrNa92y9/RUCb843IchjjP
vN4qeQwUkNy81B1c4bvLe52oIzEa2VCSbLKJW2DfQyGlhVI1GX+JCR3fCuJxzmma
haz48WdYr/tOxy5s1Wa9zkeNPBSDyXjTnhgum/oMnQ5gly10bd1Vz0cM8Wh54jFe
FzyIczpbQRGR0jSY+9pNBeMXxiOg0YkfadMn+ERJMgk2zh/d/OBkJakTaWSJfjQd
9hPiqY8zk7wua3X2LIH06eE7goJpIg8dZir+lJyCccbpiB+F64K+DT+zDjQ6glZK
CN9BOkx5FqDxey4OHsBsM46c3bFfsBjJXecAsJamHNLp05e5qtAWHPO+MDOtr2gX
zXSKDNRnhudoS9jcatGSYkB9QyEKlV1cIVmw75hi66iF8cI1cK+72ozcnlt3DxfL
099wd84B2hcJO6RGUNFsuRhABF+FmPNvArOEa/KlIQ9MgjZJ9HonQj3tk2Jd2XJs
us/qnEDu5miDytbNpKp2mrZ3xL4W4Agvr0KT0lCvucJiRKTofMkJP+JA6UjR3Rya
J4SGQhYhnIyr51ZPEJcghwlQBsn3s+3AEAt0yMsiA7zNJNXc4IpJGJ3d0brFum8f
LWZyDIAS5Z7xlax9Uyq+e4OhAT9nPuVpBci9S8XEGRtTHugUixZEev7S/mP6/N3G
mYFH6stKFWeHVTKLghvAg/Esmc4+aIwAb7GAdbgzHa7o/m6Du6a8fkDinkIpAb4+
qK1XLO1fnh2rBfaeadwjwB0CTxsKgBLK0TEh40+4iTbdftCDWSrDr/q3zNEp38Pf
RtwZxFZ7cixvxezHh3iHOTJ/52TPhEvKBMbtxpf17Zzims5018VVQz7aV/XoM/2C
SzwoAslRiCFP83vMYQn5mU5YwDY1pIJeXU1CUqKQDg0MDgO805aonNkTtMsdlo1j
xxS5CMaW1IrEicJ0BD9E+zf9Tuobwu525P/w29NGqi/npvi/d/f/vvaRDaMHFWyK
owZDgS4ThbrQ474PEQi40izT+e8Fi29Ll6dy6IWO9+4T8rADM7VlTqiqAPslgpeX
U4SOF3WUrcJFkqUe+gdNTIyT7qz0yHpPZ8tzgjp96FnXhLrMg3rozenDXlSehcXI
7AG2GM6t/xdmGgqqGsWJrOxtIEsDnEpTnvtUsz350g4vpERT9MkANWf+rQ5987xn
PqLuNh2YSo0yUD87+czNhMETrAdZH5Vij3dnt0E5rf8ddiPuHzoybPAdunN1NkgA
JYp+eOtCM9j7kk68niUU9p/SVhpW9pCjfTaPVilohLcMawgRGTtpqnil3Qvpa4EH
t3frLALb00vsedokCjDRDGC24tgDskSzc2ghK5mxfA3pqo+m1i0X44fp4Jp5z9j0
L/pf+La6bqLVePa1sBg1PCwxtgPOCQq2Ah9ykOWrZ2pMcEQgeMbM8wm7xJjD9laA
DLo0JMPEXfG8WDkReh9qxJL57Uz0tvzfdy17AO1yRMucABlQsKKFRd2pwsZOpb96
BGfpKN2iJK8T3QKFIYlrXGcjdfk5x4gvoPACVGQ4Ezz80Rnmhdhs07nMd9NQj36w
alBOB7ihMmkf0zvd5j9vX/sUlQHVGjB6nkJGkOeSrz5S5STLCVuHixi6KObH5/dN
vppaTUBTe2MBONVzQ3uiat7OhtjR/AXQ0unSst/KyjVOHtK6s5ow/a7AmmThiJ5Q
vD07ThogDo3XZXe5NjJIB55YWKtqOTVumbMIz+WVWsK1X/fEAlxXmHdbTnntdUfD
K4A1lcbT7rcASfWravf/goRQU1Ma2qNeQeMkFJZmfxg4s7znsQifxtkmY8Zor5P/
Tph1E/bLu4qQAXYYNg5Mn+9RFRrYUFlok9495IQxK+H2344s+fN1sH7AdNOKZZkj
9LqEW8EMClB5Lah7Jp33ODx56E8wLvuP/XlnLq/fJAyk8nrVV6CQsQbHg5A05Iz7
acJnqEs2bCrKrhlBmEvW64jbxAbFrKKdJgA2T0vlagZDbHmuPoYuc+zIhYjYTQ8j
GzNsrF321ZagtY6B149IfbthVAsM2+6VQxy5KbR4b3FbP9h78V9dgwWx70zYHDkJ
9O+VZ38TxCTqh1ZM775JXdXpbZHkZHWRlnv6eEsipWyLbFjftLuD50/ifLokAm38
DJMk9gKTUljj39vS+NjyaAilIe/NkmYRRNCwezcQYW7Tv9JXlK5aUfUwyeUg5VXN
i8jb5pIwi/KZPAbzKrmBIeup1o79n9Fw897JqX05AEfyOVJkKvGSXOO/u9Ze+i/Q
HcHMINZ49Le7s8OF0RBRFYmOd8Xugdy37CEktC9a8Tb9fgKYHpg0qrdIkizQZY+R
B1GQX5ojFFiNMpuAeE/WcArCbv4y1aa8PzNoVnSA2iEJRcRb7clNUGeOA2X1gAOW
Uh5d2/Hu1MlUKl1veFw5OgD3vVQ0yOA4e4qeLVuLuXYe3ILxOaIXm5cCCpoQMcRZ
FCRGyPSb6CCJaoOtzOkAN6KVYnnr4HMvU3Ih+1K7IVOz3AeUGN3nGDGlZGC48zFG
K0qKtyLBl2bmkxqbBXB42BpkrbCUYM4cQdKC0qjt0IMpGSaOvyMlDonV1IO7xVF6
327sJPFlhvCaSBpue1asB9X0+ajkZpeKNgH1VE6ulLVx3I+BZDrWRYKgpxPrYMZx
kAV1G5Cvl6nTAHxPznIbtUwM/x9uGx7L19fLJ55zShSymE7oBS4V8L5T3uvHHb2O
9CtO0xB0aTqle6kYBawBW3CxDKK/B0TXBvmtPplCL9Js9VlNZ/O2vylbU0IaPesx
D7qtnBhSubQnCtQCHeLdAvsusHNYq601Jo06FTfsh4XhC6wAP/kxSFyMOh3I0yL7
Ac+y2tMwz3vidfgsICrypDZmb3duyWESqOUvsw3gX5+zftivBA982I+hKp/SnJLl
TIeU368zRq7MopKSDEgizmvIMSkzAQdI/TtDrNqLeyfT9YlGdbmyymL9d4heT+lc
vFv+udvJctD+fu1XeAeR+NarubhH2FlXycRyXAXTGddeG+z74lG25ZVTk2GnAJw/
lTlx0QzGwl0CTcZGYwSQz6Brxq8bh1IWqv8bldtOn0MUPn2ojzJryx6pLUGjDS9f
WaFSPhIxaCf7nBKLmDhOXSb3FOx+4oWAjJ/9cdyY7Qj8/rHeXg++qTuCVOjOkOVJ
FwjuT4JgSq3sG+yqal/Pwx49npFpLnOTKXAZKzqSBWg6O1VORcySrQbSDl5Ny1MT
WUci7hQf5eL9eJjiwxjPvuVSFQfRlEpg6UbGqkn8H0pRvTWta5OcQYVuxp9GBBxm
YSrpPpEyXt1UFG7eSsIH94rzTgfFGIef4dAF+9MTirIY+DKJNzNEEXDTXEniIYhe
5nQ+l3hJFJxzQaO9XVzJoNTQPZ8zyKi8odFjza/LMCtnHz+Vqm1DaCgZH+leAjze
6uYYB1W9VyPnKRWglrqDiPu+sqRbxjPx5EtVpIISxLkvcnZ3RKme7FRAFVQXdnRA
Dow1ElAsksep61eM/xnif0EcMdaAP3LSDd7X6Z3ZYPWBcJXik+Dmto8ir50a1EXK
ishg89Ez4VAY7emPft97LGNU4QsUbx6QaHMX43RNT9kxEGWOaMJMZzWMfGoO0Loz
kMI79ftAxABdVKO5C4sr0vguIlz2Q31KCnJdiyNw/T+v0ia9EI/4dAcVjxgLP/tA
iSGPKCp3DMUEU54zyXLPU/HM2p0D7vptirXm3c4W7/n9lGTk288zk4DWetRr6A3v
XotWKCy/JWC2DbIScMVz+1qXCitgSy66AsEokF0XZ9thY8LZmHbJsKAjzNBmHhgq
BRD+IP3LPPUQ1zSpZLeMOMQNALRWXeHv4nIrK0Le4XsIn03+rkuD/1Ik5OECK1YF
0IxJ+F2TzgMbYum40KmMysn8JPHB6W6Y15ibenSDH26a5PcezApvugmknjGzPoI4
NQgnkGmY0PyIUBo/o21qMLdxMURAfmPC4693xsL1PYvRBwX/vnPAjaoSJmyZkAWX
F7qpGzHLg151okUCkt92+MyR8zk+59IQZF2wwbaF6f73rR3shdd9O/U1Dw/DSKRV
AoCWoY5Iz3gBRl9NnjojxvE4SV83wJBiDlDZ2svbKq4moSoxW4QIBq9CdRlbAl7w
xQPDHRovV0hLNUw6BT2eR/ERiD42rgVj3Wwk0Bz9yMYJU0QZRBJs9AubIugyhzp9
WKxLu6aMA079hg54wvPm1UguLtqotYt/d0XlOSFMzyaVrQmh5tMI+U4ViuxU6h0w
4si6N6py2Eo5E/ehmkbys7wbLnUGei1TWHaqMdv/SHYkQ8y5INJXdVchYbfAYWGp
CO6SYIPT4rw7W3wj6I7+n39hEr3mw65Y9P5rIiOI9Of1N+OhTAgf78MugOAjlwxx
v9i2itzR6RzNbUdiFW/1i/C29zDClH8b5miasWR8RXnAdWNfeRmatzfhQvvQSHdu
dc/FHcgRm1hBOoebL+sKYKI19ck4d+C7GK/HmW4eUaXwUVABLp7vSef3GQDbNI3l
+9XzE2obbNks0GW21V1tF/SuLJ0xjKUtsuYmtE0+Y2Gb6nNIofzzlXdAOnwQ4J3w
4lriWpauWJ14hNZEp/BabBlVhn4PC8DHXctM4Z9zg130iigniEtWurrRtUCfqFSV
f8rPZeY5v33cCQxx54rP1E/oIUMNp+MzC9QMpMwZq1jT+0QKgyyZdbOcGATCDJHN
H4+XPYObpL57mGI3TnCKyOKNKT70V5xqV8Qe41xCcBKY3mx2ph0wr2vTsuD3fzHd
qwd4dHT4wVI7FEa0UkmpOP//4+uq2vfMMy/sm5UU9yMBFuP8X2PzV8Nze/IyvaFK
dkwoTPdGiuZjJDOndEnTMuZ5U7cel/+oTtCF0Znb1qBiBbNILL9fAx2RiTjTGkt3
eOKEJ3kGnBVDso5jiALMNNHnz3n0g6E0Vkd/9BzIZlGoJYh/bKq2P7+0qcOXFi7+
RT5LnxZWyM9V6TLmS/H4iQgX4sCfhWtDcR/rajH3K2sgNOedjHDI8JQr/co5R6hl
FaysjgmM5j7rdZ+uW1e13f53Pc4I23tHBTo7mwYiqHZQYUEQHObravvfYGxHR9tX
OicF7NAHSn1SaIx9KlSvZvNHXeyzTeJIBgQPf+0263ncvj5oR6Tu21OnwMvrFXuP
0rjmtDQ9QudcnRrVo37SOUppVyXZLqml7A8H+Oo4J1HWiCGYR2yC7J+pSyjkTe6d
Wz9RnykrkdezWkWE6qvHCY7aaOBQjkEQth3hQelljclk2Z10PsGSWJTnDwLzL9e3
n2w4pFRYZQOFCouMMgDCC0fSUhivn9x9yPccbp1Zlp9s27s/bene0767V7EbEWyf
k7Wji2arxvZI7u3irN0zeH6gl0rPmOVi67q+8ruI3QD62O6Nh/YVogtSG7b5Q3AH
noqFIwVaOEQO4YzSapWroaQn8ZC3Dl0sqN/omoUgQiW0k2+mJ6S0Xiot+lEDVEsF
9TEPu75GaLKvdQ+nv3GBkMdmQfltNHWHFuEdkr5NhGeWHnPdq3yAAPALscdWIcwj
8Yn2DEPbRUdEL2yNDoEWwdrm65PaLVx3bvQ9R6CRTP4uYrkc3/opfFoma0eQ/FTT
GHP2hvk3QZQKd3PBwXCg4kT7EIQ3kholDu4CUAKaCH/FDvq05/WxyxYbblUoxVvb
Zy9+RTNsEBKaczUovDxx/5BrrywGoBws5In962gMKhOAx617/UB8OZd6wSIqkof0
mgUYA8e3c2tr0PjhqIV5AXYIurGXgUD8pWZri6QGdRhdkkl9z7DXCiCYvRBRYTGL
zMYON3GfEpc/x45TBYQHCUtzR8ot1QOLK7ea2VhnAUi0fApxJIJqkdSA/xeX+0Y/
3C8pX3AQO8r6OKBu+qjC/JqpLPwp1zIacVOfT2vRL9HvHVNYXQ1NXHwNxFIQ6YcH
csk8K8cnB/a6xYpLpmvA9zsudZvo030bHHJ6/MRmkuAmEv0EgQriqXjmr0kLKqX6
GUuWP3VdlQiUaUNlI1tgQyKaMzp1Y2rzWycDeM2KRz+aS+Ixaq93ePGmKcSz3/M1
Yf1SkDADMs3DW6NCDutpazQqM9ivqytY9oBSxB79Cr1Yewm7Xlm6ho/GXp+xSv4P
f8OjiQ8Ai0/peZomp2MeqdPEsHgqdmCFDUUDBSltk8ZARW4Xx5GTF6hWd6YzW8Md
3Qg4D0iGdPTEWq8iXy58L8Ot0eSnGGgSqCRl21OWk8KevZklWgH1IiXc+x2F7Vet
ekHdEDsM8vkDSUWnSp2zpNkfz9YxkPHLUqCFxciGQejpTgzvHx1z8ZwlaO82l37d
cm+sUeMFZQuJ6pH3XUCMzUVZmDBQtabHoleYkEc147WXFoyfV0xPdigWkGulbuCw
WGIdZI2yXMTtjcbvVCiLvjqI9lBkgHySpH0eR5RUuJ4EWG01SLh2pxmvEeoSNhba
8mxb000JyXx7+g6O0QLdgaae8O8yNpnL5nq5k1Hiu9gIXY0M7JkHQ+av1czuMTp/
GCVGr92h4X3i6JrVOiEXUwwB6YCY041IPMG8QqEurCbOehFkKZXeb+JkD+R7cV2U
V+nOZ5xlTkcfe50J0zwyPKMjAG/SjvXNNBlB8efFc5ov1Czzy30+mM047+MH93C0
9E9g1SWFFNnEe1Opfi2r4gp1nGK4Rwo9OyXOlTtAPZ+KYwjb8pEYMHDjPAgHFbea
NgC41DBIKYuNAee6yTrj6MNc8JS9f1ljJCvEn6dIXlgBsdhxHtLLCxmJ+9249hkN
6Y3uZ59HC4p9gB6girxVRQJNmpSjXECwE8H4nsm2GNdxXfxmwMhduTb7O6HqFNkK
l6lbIx3qAWQ58dx15GexKbIssTP/+HeUHgegjHITlpD4y7Sh27mAu7rmUQpmW2fT
6KKz+DC/6nd0sJEe/MVk7eDB+1EeTnh7bbLhjX0lidMXc43VcYZs0xTtX/rvQ86U
NrJZejBXUfYgByy9kaKkQY7iirmhuhJcgWWV9OiLrvnzm6MISAUnXDdU9AvEykw/
ICgT6oW5rbKyvqw8l/xU/aOHBPFXPtU+qo6rGMRDykIJf2vZPCrn/83W+SlK+yLC
TN2bAsqzjeuqK0nzNHZD3x4wqzNFuL9t2CCGHBpTPEDrdu9zGmD0dneJGcJInn59
JGZZePBBs9gM0EHJeB5feUBIO533c6WL8LL819TxkWoVwA2+1GZln+owtaYXsiLp
vURUniXj1wq5jpSr+6riY7hPm9v/+cdkhass9E5euoX92Vrj1Cl1BSkVFMV8a26c
ziFJdbAb1iWqBurKHK03pyT9EFi1cwO+dqKxAAn2QNKPM1cQ4BtmKMjHwwanugqY
EQpu0bttFc/KhwNizIASge5EsStm075ZC9qSr7dtbquEl5IMhUECU3owrcegMKzq
Wzb6zO9PjQIWEBOg5orpXoRGmDGmk8xND1j0EevLLA8WETQe+Y1sibUcvVOfv+MD
k/8Z76XvbQ8rfAKpoYEf/hqMBlu53/gW0jh80iE43b7UVWAFYi9zWtR60wFSXfqm
PKcw1BfR43M9ZgpC5hFodUD6DrzYpTVta4vxYsPjvPIDDTY9Wtfs2D2a+dfDdkko
W5gMLLd/WAK1ViYZmkQhu8WiAdH7/k7d+/vSh1m20El//5XDNA6s+ld2OXcaEXjB
OZBy+U9OKO9DsWg5jVPun97z8WvgPPfMbwbcmeV+n75X5uhJWakJeX/7uqyPlv5c
bk2kYzjRbPErQBwUEJvmstIWsgMWQkK6FnNFSq7zbFPYJf+s/khZwN78wKeqgnM/
rEyjjP2DN7rxZvb7RYxthHCPgF1MAp0cMMc0daNDg36WJ5i5fevtJvkgwjPXNBcj
mGSBUix7HZG0lNA75Pi0CQii0c95BJAMdvjRMl45bT/PCOCV9SrIRp1+476Ignja
vnM1rtLJq/xF4yRE5nLLBpgBIrBjGz5U9DdXvf2Zg7BerNwPsih0ZgOuw6uztDi/
Qo2IZFAq1bDv2RUSq5m1p0PaIlN52pT9Ai3DImnEdEVPYqf/zKdCuEsyFd+A+cMW
1YAhLylMrgMUvbRi63+FcJl5lcQ2b5J1YMM1lxUjMbArMW6PbCSwzS60B0nYrxuU
Wp9aMBnT6a1WihyTuuAtpYJGUoDSzmc/9qlQmYo3s4EPEqLydSPvuJ7dzyZiRAj5
TsWYPLeiR9WG+6jGVfuv//Dby3kufwifb2Y1uQoUwj6jbpE6adq0cp8x1lBdRk9i
ysgeF53WlpN6TWvoCBsonfmrpoGqCC0NRQicsgTPLqbZzPRmYyjBPA/b8sXghIOv
+H2vQapcwQQhD55K1LIoEKB6ukSGP5dEOtDqnahwl8A1pD8SllgnR/SbBX64HIuw
AlPQMDJUWy8OCi2T8bXWaE4u9JsQNl2r+HB1vF4935cm3KJVyBvPsMrhm3XZOLmj
JKdzQiCNUgNYMhLdlVqgIbdvLnUQOf7YnMC/nvufgvRM1O7nb19z/9iccB7fzH6a
ci/rSyg/f513zGNtmG/VBcdwtZyfEYSAFe81Pk0Wf/2e8jY3FqAR8Ao+tsyLtpjH
fzUEotP3sBQUY6adv/zAkQ+Iuyd4n/mFdVsu8rkLCvfleeG5kPhlpY9Zc9rQjjnC
BvOMXiFJpooyrRGktz5SwyuN9hMDDBFizQNEcbWtaHNgKJt0pFByPKcVdU8txJtV
lfXX2I4rdYsrYpRUeEph3uE+fN9/zeeC+zysUR1KBYFDiDFJ3Njcx+L5qgoZeyOT
v96D1Hlt30fmhPy59UPuG/JQqFdNCX89yzkc0wBXGE18onhSlgYV+GtEYKXZeIJD
g69o1vBD+UKIpf5zv1fikOoG9npBOrFGQVlSulwd2s8+QB13cnQVY9VSWKgk7A/S
bQTSMz+wM18qXyXevMRi+Mxw1WeP4Xy0lDjpMf8+Jqz8OL1+IVQhSaU7dVOqQRjc
k5uonInfuCxRg1vqUbZbHbaAkJ/nWh0cHsbXB79++zmGxoN65WdTRcOiPzMofjkN
+8mqUekKVDevKjNHSASxD8sdztCotCDTZmU/2zhOTGq5iozhJPJaH8pOoB7gN3J2
CyGA2mUt6u/q2rlMrA/GTwj77EhXfyz6JXzM9ot6Ut8hpQFUzfhxsGYsQp+/BZZx
Wsw450bAq2KrwcWqdjxmEv+rYw1u4LPai9fENapxLkqMFVixu6owiMuCKTU7kITF
6hDHv8/H2CeaH/mTpZCBxzCHM+y4+etAjqz8AgsCZZDfWRrAlVKHg0091Bdi9HWr
8c1OR6hdXJJ11Enw9sNmXu7RcNzJle+PfDCx+2iMhtf4wlE5lA0c6H2JDpBCo9LB
2SvCIeMzqTLeHSWUJu1S5SuUF9N2q7AL3s9sOjq0Nz100JvAJbSMfFm4wUA2yYuv
0oL2TZwSgHrrobWewsXnx5/uF4kccG4cl9ObTVkgsg3ay/0u/u6in06kEkhZnUqg
ESDKLf0zMpA46xznTkx+a2uuAcw2iozO7w37fL+6br5RetcWBHV3sZQg/KXm6gZT
C7SoSnQOG1txmjaHUtJEeC+QBbCul2b6FNFWc+G6yQahq7C5u5eH21dL/e3AkXav
deQe0U9i7/MjgSDTxcKMUcCup2PsCmKoCx1EmWf+Ox1RyJpGlVGlw3BuEOB+SrP/
vZ8mE08zs3KaTTx2OWK71nPofHcwoGSM1bUIdV5RWSIq1vYsf0f18u59MpHzqxNS
e/gE+dYC51K0SxS2LkfrEft8kzDK1mZSlXOKQ+DgWITla6/lYoIi2x4ENSuDYJqJ
ununuSCAybc+qGomIsaSLJTmBffatzc3yVNrCBSy5Esh0ThbHhhPXHBlE83cnSgU
InbLEkwG8KkvAD4tYCQJun/+veQL4tg+pSS8YAW7WBIhBaWyQ3MTL7rOmoUQufuM
xeMOtbSmO7MzUP95VkEa+5Maq1Vmjt/OGUTcOPIBXdBa+g6BUXVEb6SQ07gkh1Xu
OK5m7b4Ekgyrpx47GndQw098GsnyPKWiAVJfFdHeBmhqZ8d+mmQBKkvrq+bfMDDy
DW/bZJmT4NEfLxcrnVL6YnhuWEhhW2jPupZ41tozvN3IWcKdhWPLB5jE/JP9uq0C
0lN3G2AMwoq+THIbFWVe8+Bpa/x8puIWtrtDwt2okzECptwJfcBzYdCNL6xxgzVd
oFUPPBRCAeRN+F0wu9dhJiq1MAli5UbkNfp6ki4JWFGbjD4WdyxDsh4a7I6Nt3Rz
25tdrNnEKNS1Ab6J1Bf5G0UhbE2lJmNm3bR9XOnxS/6TPoUGXVE8GrTlJeRlcSQI
rZxDbsdT+dDNLDVQruuDkrT0AXArSbTU8Frmn95ScVYTcCtL4xEp0ml8h9H5zczk
QOKS3tXFUIJXH8g5Dj6co0JhFRlYqVW1J6Pk1H0lyk9EjolrJINvwIwCeWa3n4Ds
3P8IN/2uBoLs3JUM3WmrA6BJPN+ufYNDWGRNRbXFM0+Ba4RNG+RscASZ/Z4X8xk+
NoEK+cjwG5s+7RkOYmsfh8xSy6v16dwEUQcBnSyQzuOR0lHrUooGDZKgqpqhOSXd
NoNtQil6c2zGjDF11N3bIlS69PqNVylhDcrk9ssVCybFcU1VQFiG+C6jBx1eS+gq
oRc2chIZiO63UhjxXzLD9b8lJWb8bjwg7nDBapiPFc0qSU5cILKJ66Xuoktt1laZ
7iOb3ZXpdNTuvz5EFvIB6yPM8UowofTQbOjlOrRDyG1y8bY6l2J/3dsC9EWipoJb
2FGpHe8y6gmvqP9AGYvdN23bz/zwLWuMN5+9duIctqjVnXEnpGjaqpdL2yw2PVNE
UtS6NUe6W/qJsSBld7ghQjsxtQa88hUWJAQfQ9N4+/Ge5NJc6UsVac8alF6/qJ91
EC0E35YjFoV+D7HK11Zj93tw8OMFJQ8BBvVzWM38zXNL+DwtR/CeEkchkM7CPXCs
mEVwMIsaAPB2XCkN0gqyC01kwZvS59v7cy2w4dESrq4MZD3Z/R/QeVoRIA4at3i/
oCWG9jGhUXfDl0eoAPiz/q/K1ecKZaBzNh9V7B6KzAn6OX3JJOgSWn/MFreHjWyO
FSp0yJhpVj6LDRMkzSs65xoNALeC67A1e7zUyWBd8mvI8VP1dn8HQE07EUD+RPjC
tUOTlOa/KVaqFc7Q+2wd9zk8fYB7MriyK2gCQr/c3TcsXkWyiG+w5rHwlkzogHSo
xLwTpjk0S4GJUE8lPdrIHckrgTF8+4OX2mK4gv5/hNAzGiRXABaFZ28BgkX0WE27
ZA94hDh/KfQHlpxEi+pip+70w7Pseyz10C8GtfINRF8sqmsTrYpPdndmPq8J0o3k
gfbiHVPUDpss+f5PCElsjitSqXypVgr7RU38Nde7HM696lxFHbMKuEjYasidc87i
5ZJ5725lU2A0wXsp6J9Q7UZvBHDGoBnoyJn/U/OqWS3HhZvUXsHZQVrss++FToBr
qG2kLoYzP5JYPN7LF3qVQzWy7B9iNi3tX5ouaDSK7QOd/2CvKYZZySUBvoGYl5+W
ifWUvJwgYZmNhSHX79atYOME1T0O8GN5O3AhKl8n/v92xXtM9sGiVh7M9dKMNXhl
BcRks3j33Jk1WHT8lPdQe0ae/LqPTIuOLEQG2t1HzHa2oV+WwP6TH+qAcCi81I17
2JCNqXT0UDsfBmE50XSls+AfrX3t/2s3CIrFa7f2NIlv5CBjUPvDTpEii/1EUSVH
PM4ZmTBm+A+H1mj0Sra181JpgQHQVebiLcDOwFv7WXxh8ArDWEzpWTxefaNozi7k
7HzSEG3nOK3uJyEMSkhjQLGICvQwkRM502w2aqnIhvKTUyOM9MBiwVNPvzhm43h1
UWo0r+MHqBNcQ8Um+7g+pUMLHsjrHtPxsKJcnAO/HmTTAK4TiyR0ELpnkweJKOsH
DeScddRziHlAiRYbhH6jbcAmmrpGm/GZ/BIa+oeORjjcmFBMklDkczcDYFHGzEW8
dCJec+4uVdKCkXKYVrXIoUdmXowxnVoznd59mLdh1njZoLqr0ZqVobtVgRAFJuvR
nH0TRUoXQiAdfGV5d+GC26h6AFBznx5BxMRp/eYyrLC2B0zQZLA1H47zHqEPSHYR
mLj3GUNcGTD9YhqAlzMIoc8T/x8ykpRJaIabkzISMhrIPZmIPFb0TtsZvkOfMn13
MbTh4RVS8FHRws/d0k+E7NlYiX1xP4egXctezXTh+Mhjr4GQyOECUqkCaPtB08VA
2n7aeMz/C9M4tW2QclKsU0ufoGc9QPkefE6C3A+wQk+wybkpd+18X7o18uIeqR2U
zxfTnQUwf8d4nJo7qqCAShcZCNks2hq2NM0fEDtR/5XHAZoTaJj5BWC9WReYd0Ic
gQSqJ8VJZEDWq1elE0KxjtBLUh9Vlxu6agOtJTsmtYjVrejXhjilLCbqsNlTRf6F
98f1+QhzlM/dbmvhOyQvUojEWPV9+zmvr/UcSAgQjUAQwTZKr6rdB9SxzGq4eROm
RT671fYj7xarJ0mi7CzppOlGnIKYz0xIwQ6XGT68TjoNNzqNPHIpVSN5qBqfYqCR
l6gNiAaHszlqEY/yCAt4i6AFj9Vi6p0/1C66jyZiT2nS/eBwPRojMYG6g6lMbYBv
kMoN1ptDuOpfJvZZ0a+t9P1C1lqibwENRr22nr4uUxtM0FBQFl3EMkyDjIlbDYho
3V7C2QcJm037TCx9IQo3NIAkDaG89kJxpS9NTJ2nkhLCqBe0G1+68zdjzHs7bXbj
KT8dT5Bdy/FhgvhIZGmG6HzVVtPCNym4d7Py2f5cTwhHKy8VEGf42WdngvRAifu3
JaH2FTEca1gvaSjpqKOIc4kS7RM4tqXgInSpE2pixVqzcgkF2KF/HKQ6wk4h+agD
27R0cYWjYXuIOB59f7sC0CJlX6303pThSalyo+aA7Exsp3eKJFAOqapsgKvYdcPz
JLp8OA55FGyvy5kE3TsgAHozSpMGad3L8leGvArHy6cOfAbc7XjAzRxmNjVMQEAE
2guQyWDw3jA6oiKqSw5d9rTA1DUhzA2B7oqGFZPBfIdjm8CI2e1gLhrt7jRB6rAa
JX8mrCwEyoG89uQirOADOt0z7J6JHWVIiGIVKvl8h3QcfSIm5KQwV8iNEwXHOpge
AqVcjQNzt6M+g8yr+WRy7CfUDo6fxWJIwnffR6SMD+CM1k9WSFvAoiIgM4OlVU3y
4wxTCCJG1L+1wMnomNCC1iAmaBxrhdNLKqBLkbOaiUFA+jcz2BUxWuC71d5ga5CY
OkkfyMdSw7m1hpN6lZywnc9IXFe2C2iAtFPtRTftv/zHgPbvGSznM8q3mhmXbHOA
+uVPs8xA70gR5TGMCTdcrlcJqIYqvm6whKAhZ5rAqXwc9IhioFEoZfPqaAwNLUKz
ur6YN7Xg/wUZF+TruvedjkEO1mfRdOn3osVEVziW5GxAb+5lRJJdhu0v/CxRwhKg
XGyaSjvQ0qiis5x6ffVtM84wnosQzqU8C6EQ/zhV/k2yByTXp2M9vLf8SKolKG4X
oNPJbWWCMFiPeHb6GaRyAz1Q8a6EQg/oL8JLBmooVt3F1vHfDrOBhFl3slEe/ezz
kRU+mco/552wIyEKr1SkgWAlQjn+K5bpGs8h7AMwVsTA6yL/OEqaamJZKfh/mKXm
A1JYQ9NnbVnpUozTSEZYXnsVXgmMOOGhbSeW9tMSGz8E4GAfU3FvE1hF5LM102aB
T/v3RvXuefB6qSIO0SV3K+rweooG4vzqEcBv8ttP2Ro+rzTYpaKK3D5X7cEIHJ0q
aHu8Nzazk5kkWSfzCrseJ2E3nGbuLpEiDBA26AerOS9kMQiZfXYZRBMv7hdyXn/7
UOcIoJppMOdaeSHtPJsSKhEhsGJtqpwsGByQHdSHmZ/VDski5Rx7O2q5yTFO1Ykd
4XRAeMQlPXcyCOeorMlPRPEets4Tqt25T1jB+bAnOOmjGIdbXKcJjl4RNCFNMO6f
WQhb4BGWOqH5tu4P5X/fgWvBnba6bywzi9o/fsRt+1rSu07fwRzudsTQUWTZst1a
W+osNn3EnetF7NKmJL0V+KI7yvaTGuFtIcr2hYmyIGcrlYjjpmOf2E5UcwrzCkd9
QBgWAKYOWQINLY6JEV9IAryMJBMeUV5QBDDaPDNExFQzZSeOWLB8TmKj3sKvptzk
CSKmcHXI7402UKz1Wa80fbCYjbTTReKdCZ2Bm8whsOPZba6buqjsmjkq2jOkdtjy
pmsW9508ytbQ/WJz8dRkPfnkYG880jYyeWY37fXJoA88rNG0PcsZyi3Llp8zfd8h
fdVDBq+y/skuyIXDvowqi2PSox8n5a9TKFnsgn+8VTSE4C4Qo+esLAtVHpWHBoSU
efyBMfQ9S8JXjazaDSSe1zw2lWOtcju2wilsGD/wsWudoM8UK8YzlQGeOn67Ux59
fVP36rSzRGZG7ACDoPspJB4EobkCxKhrrUakl7zxqoxfWl3wn1uR3SUq+P1IIQ9w
6vF/bJu+Ngk+Chg9VDhEPihWkJfR3PmAMPaa2fLd0H81NF4wg1rqBFwAAWLHp/iU
A6V5VC2WuSI9j/DTRne8c7Rqdo8NkOBEo7mLdiyglzIgc+7DPwYL+aXpo0W/gBp2
rAr/PFdUCeJ76lsGeRfKGoA4zIGSPl7lUaChUAFbwMreGVgLCe4qYBnkESdbE6tw
aGqU3lp1Iet6+pbCV1XVIA8pgUykjiySv68KRUL9wsNyyYKsNDcseYCKCPshoo3+
TSpFpoKvgn3CPV1SLZKUFKDNN0faY/LyGyGPXKA2Mo+RpPXOjT4WtWk7iN7QEwMB
iYeRNgqYPvJWXA3S0Pll7pLrKTlXRgVp2p0Tu0xSPoCprzNVNEbFzsBYc0o/Wvx9
smlB6J5nQBECmF+z9/k2xSHYd6m6aEWGkbb7bPTSuRM+McvN24BveT8Qhk5JrCPn
OPSJ1nSU8wVpQ5+7lRBWJOEahJfLZoHnyfNYzWjYRdfJ6ndqUh/fNFi98SbSF5Fa
Q2Lgw7j/5whgO+wfwv3ko/x08xol3fIIPVqX87RaCzrK0/5WPuTJBrOTGG8fDKmp
li9zw5Wl/ytjYvZq8qmWwxjfoBwIT4OCuJj3MJ0mbcR/Z6HqsmC1F5OoHw3zJGvT
kp9iHXOzaxjwkS1AuCVUzgshbaKF+/Kv94sOmLqPrtw5fStVhHeRYmPFxLcOFmF+
jAMHjNlp201/ld2MuplYzT4I2KiO+tjBe4QvnLbmDa/uyxCm1YixesZV0pP+4cAb
uTGiNm+En6aklCAWIcrksobxFoMtO1g2rsZLjK0Kb668fOvnugEiIDve9deDGI/V
7BNbfKAnTEhd0KxINqvhPM56kPKqzM01faL/iW1t4RUagf7HlrvcZNVRyb0mUI1G
HQWH3ol6riDtw3BawGWTQUlSTc6A8cUu9sG+CWkljkcPAnOxfRxoydkQvAETJjJP
/7Rhl5Hja/vX9epRetZz0Qs2NyMO6Wk2vW1BcxbW0v7reMJCqoU9yBC1iiND+etL
OU7+U54ggW97nkqDO+geX9/f/JcSAdb779PjB0K83GNWImHw6H9LEVYmuw2sNFMG
8xrK8xygyRPQyGSICozLBLNu/yn2zI9Pa+Eix2nTATxe9XTply4Pk1jrkXmSPZzs
Z9gvPrO8OgTV2J6ZAmApRkEvinyQqZLGUyzkARXprWhCrBFs4RDR5y5JYZOG8OGk
I9U70HzrSBE+SfpAOOdRKBV0MJLHbQRe5u6IlysOd2lYZTsJowXpww2qlYlemK1/
9DlMFTSqcQxnjeQSpSVjdBXSLaGDL62g7ThfPZ8/Nu1xj5o6ScwFE0RUBqo9Q+eo
lNXiybPBXtoLzqGY0jYkxeJx7T+8LKFzSIr/3lYgAW6CPcCThVBSTi5v9DFGhd+K
FOicOInF5SJbDKkb4ljnqulQ/wzW4MicPxEbW5TL03M2hAu1I+ip7jGKWVKHjqvg
PMSb69aFKYOU1OcpPuVypbu4Xpn28YPKIKr9bWg1rOxFXNHmBnjYUTSVpvcsQRuA
cHq1Qhf6tYtB6badjJIT2Ur1W93DSIlbXXMav2Vqjp1k/ll2VLGvD2euXVu5T0Sz
ju64+kyaVh5C+ksMKcYbanvC7gXkoXsJbu0I6Gq9TzaYcd1yIPd2s+1uFo/NnC5W
I9t7YDpgKJbHuWtrNXakr+0nLl7vyBmq8YEFodkBtL9zWjGJ4Gig8jefuvVaKgrC
KKMKfYZMFjb4QBgR0omE7H10mjj70tI+ha0Vk3gPPnEgGtnGzd/dY0zUjnzM4rCB
0YPgoXD6vEz5XliLwWM15m3zV0dvmn63EFmJuSU9sdeQreow5KQy12NWOQHvg2Yv
VdnlwZtVJC0hUXVWeuRswWRfNdIlLrMw7HsUmKnAj1fr6/IpqhH4rqXURbmG9u+s
sA81RFiqxs8/eQSjCaMQR7AOL+auYzoJRzAt3ytsaja01M83t+2vzTMjmb2M+iA6
qv7LY2JjyL/8xRK+0H8vgYSbh+wAHuZzqHKttSsDm1DFVcx7dhZ1Ph02DdrKJpPB
52eArQsfuXQsWafyBPl1OJT6BsAxb8j8uPKECYVgVtHjwvd8sQ5B5FrkI5INGxSI
y4p/RFk/LqHtD4RRECeA7LHB3Z5RcSUtNBy5xycHpyUNz105fO5d9h/PUNK7sGzi
gGj8b2GaZKDPrkDOxhuHySQqBCVETLRaESkMKTYYRFB0usWFmI42Z0Oq6YmzHegC
7/4z+OJ7jEFiE2aQoTjGPXizF2z59wjysclyb4/NZIs05Y/VhxglS2mq735bKLzy
kYV2EaWKYPVwFVXgU8B9G2FhmV8wg5xBbIyvfUswYGZiM2vbBS67QrvzTD69Zxjx
SYwMbiHmXR1M+a53kZyUJDxjmW1aSriHfE7qpBMZlBzpm9OnIhK8OJmdKnFecl1b
zU0UmmE6PIHR2Rclt1YwcaXkGsbj/6M3KpKUsHhOksk6Re22u3Xn7gnYd0/V6TUg
vYiBHWter9NQzSDH4EtPO0gtVlNmERqVsmoZQtrnamLV5FL609KuZ55OTRZEcO/7
qqUI98x/fGGGhY73U2SNZ7SLRv4OuCZNq+sHEvDBZbViRwQIrPG0yeavvm4SA8Yr
hSe8h/71TS/f9nDvyN1Jsy7S+YhCG8s0ZnK4DWqCj+qxgDU+Ep+IGSavi1uusYYn
1j7f8qqnmoCHAA1PD7Ehf/2VBUpdH0H+fNqCaJcYTr0w8fDet34X3EPeX06QSi01
IcwJq4nJvltn75qFODNyihVZBP+gQA7AAl15Rrieqw0xbAHTpK4mfAPLfx5UfdzK
QmA9czv9PAvfePSoqMjAzJz+tNZKkFAopbJrVApxnKjKy3OXmmMWiqqQryABTGUu
544noMLXkR+v8U87LgKR33Uyy8lhgKrtsgFgBNqTVq5V3ahxvbxxUja9tOUdloYc
0iGRljqbag/GvvupXFe8KMA/LkcD/P9eVR19aaaW1cKnU1oijlJ1u4Zy410YyBa5
o6DeVDpIgPV+zihJvdq+hWXEpR6t7egeDWdzlvTWwMHwT+clT/r5UiP50Obxwuzr
ceUoSAmxh/kKs2BwhIars1oM+RzJfWbwHQim6bW5HVCN4iNPRGdZPVJDoidraJIJ
29EagEI6Ely3zcfABbJLsNvk2JbvRuwPfxYycOH2rIrcO2M/c2+5ABxc6gDGjm0Y
Ro/0LX7Jq8eRckNZUnAwtV8k8RSVeQL3sPKU8XM4qnlRGKBezAxi+3g91UlsMGfJ
cEYaG3jcdbxjdWFB6EHMZNczlArydsAIKUJUZ0uwWcSIGFRdeWP+L8yQ9H4h5m5w
hzcR/alyYop/YkL8wtyszAjH1Tyjzjm9jdFMfTdRaiGgnOjRh/taictcnNxVVWs8
BTsF4ZW8fzeYMrFRONEw7kZChaJmEjHwWrOCSOp+DDFhDKVT2Hcy7DDNZm5OcAhz
StZ76nz7is+SRRfAEvnW4X0JvOCtNyD79GZjB/JiKOVSey1bbuzhAssT5mBJWm22
8mqvy/YHvU1Hzr59ZiQ6X95rELJ0CU5FUAQNlzKMCCIfcgFka49D73Xzki69BPcC
Takhpbgzscef8KBnu8O/rtvvH/rVSzYL64XSRwRePdluyXbmALMXPPyRDTFrDaoD
iqhpUJc5FXd+y58cZVN3EfA+3KsQTM2ZAzT6tcDbYuAas5NgIMi5O1hU1xD/Y1Rx
HsLYdzTz2bxrrGY1KZeZhm3uk/YGGjt3ntIMCpG02jrF/Axcb4impwLiQctqCmNe
rOU5ANES3p4PwxjfVbefoYsARzZZbhs6OX+ak0s840seQT3OsqCeBDG2Y55cA1YL
O1mVMRPGWE0XqrNchFwSsO0DYFerzIUl4EK2WyffGrzE6qN4YeyLl1Kse67zwolS
wFHEaLHABLTqcNEGHl+crkmb+8McRifSJ+HfGMEadcwmT5LvNBgzzPgklEYVWGhu
ToCYL4SISJ4osw/0/c5RMn7V6WHyVj5JkzUWFW+nLgdjwgjPbXsBrdUPv0jNKDuV
mQ0ncw8L+AeXQkBL+KLOqAtfBsErx7gF1U+jretDD7MPoelty+Aehx4ZsEJbblDE
yc1/HJJ8O4woqGHsji5Kh22bnsRuhduzR1BOlSwM57HAeYcLb8IjelGWS3X1kBEB
tGO4gS3uQAmNThTDRfpBmgFKPY3tKPtgQDdHogY0Kcve/J82EpHCAQE0l1Hxf5lE
G68FVx9FivIjZuaW4cbvKBnhYmXs1MAu/uqbrC7lpsVV9/m12Ir04kd2sBz8/pRr
cmYraFvDwGzIYMkc3ZgBAEjQssIRgcfCgZ3faUAmYzrxLjlCBQ4YmhRGs/Z0YuEi
ro02HDSvNoyMAEFF7bUeDYN+vZExrPs7l42liLGz/S2rLYevkrk4zB/iIDd5W4Q5
kbwaAHQgfoPm6Of2vEWno78p3eelUAfyT9YPlO5HoxfwhAZcgkHnUBh/+DgRvXgn
UkHYxBuCKldlfJVESVqwpPp9H2E1haeJImVdpGR8VEDPw679F+ta9UnMA+wrL2Am
8Ff2Xa5Ef5xoaja6rzCeYTcKHWc/VsnS4DmDC/fvLyXoUdCDv7J9ml7rtxT0OG7a
29ufz6U6TbAB7Ghr1QmuJpGdbYyA+edty/glLRWYQ2Cru+IoDel0+zG4SVrT3voC
1YfcolQ3p1wz7EOisb01ojBUL8UvA/HkCI1ik7tycLkBCtXOnAtHl0adhNtWU1oo
k0ZTCM1xzRhRyQIrlhrZeB2ahdgHe9AJuBR4vSEUMx0CMVUb2UJogYMDDoPIGmTo
TKPJz2IlXXKZXKo6k0fwKKiQ6bB2QWnduZ9chQ78N5A0P2rwUz4UUWkEpXPPQxP6
yWN4xhbbCraQBazJ+/Y2ZzZA7KQxW0WdRVcJ+OIaS4myEC9IrkCp5zU0/8Gk1Bnv
PM35opQ2VrHa/rPJYlS/AWXRS1BjH/kmtbDMMYVt+V6z7q2t4TJdtCOVuF731e24
sq+TTYmr8tcwGYwZSv+5XJm7kH0MDbVH59T7fKae+zmoACjHVRxuZn4EK95tz+jo
gDYvS6VpFDit4MG0blZDcrMHX5V4DBD/mpvnKhuESPraO0xZwwkOEqJxxY/q0YJ2
l/eXIIUi5sGFnXSDebgKH9an4AhFLgKGeW/bSURn8cXYoWJgnd907dHw0Cbi1weR
qi4pHpEnB9V8iLCDMn2e3KVZzzxYf5VNpjrw8V2Urs6ORoSjR1gm6xildPzJVrtN
quZGvImh560kguRyB094cos7+K7Qn/8vccpye6PHXlW2E+m/Y6ek7ymOuz7FFTbX
Xb8txCZ83w30Gx7Qj5nNMbQSsj0UTugUB4BT6SrmcfFj124Nomzb65kJyaTjQzTf
l6w0N4L1fu2tWa0lTXyMPTeFNAf1kt4ev7mMJBlGcFAoTjrdwi3wsPB9GSfPkC/f
+UB24+r/+UeGCOTcUL86wF/p/f6NBqOErefxg9DP6cJgsl2ClWcaQiwJXlh1eYPs
plDPkPlpYrKAaJGQ5prtnSwnp5HMxpSGoYeQaIoIn8GgtxiUB/6AV7n4C7NA6RZt
jCOhuRJKdKtpaSyxbMKSH/aMCgS2IMXJt2dbmmhoPVMIXFCgz+707tBejj1CHtGK
4DPiGOStf/w19hMltjuLoWGcUDrs9VZJWeCsyJULLkFQ6Qf9mLylk4M8DYW3aGPc
0jNjTNRrCmrRgFWekBdPL+8oqbsdyGDyBDPKDZ7gQtpfkPW0cHL1osO+a1oGyt8O
AUa9Ga8vuqEKMXOWwy3YCaAYxo3ic2u6oqa/XFMeN2qOwHS3D9dao5esnCiRYoZY
N7EfOa3Hg4HbwzRfVU8o0DZDDZ4ex5yE7hbAHiGuDdT7Y8OkxoD75xgrRSQi5DF2
5R58DToH8VHzS3qXSmvVJuzjJ5/PC6vNv5TfZ1IOTKOLMKMBBi3hqFI2rQwSxNjv
nfIPlsNV7eARdr6Gm4w0+Gz0x549XU3zSzUuf5OKYmZ4/5ChGFsrk5gShwR3ciCG
iUUz5wxBOllE/4c/Em8OeBsUwQeMzizf/rXxt2AkG5muer3W8QDTPTr01KNC6whJ
LflW4TbJ+5M/+xalx4H6N/qcIQ/o32CxaAW1CGiDBSxe5qdhDqSlr/dBMloseiUP
mkLVrk3aPvP9i8Qw+3EBexBWUzsLOZcKDnOgIQ/C8smTpITVPCjbCsOn4/2NmG9L
aqe3Y52ulxc+j++epO4jwdOFPFB6WrejMr45yU+PUngJ5dJXrVCGb8ufgiNdMcSs
RK4bMDEdAiGUpfjzhX+Mfs3nernB44FTqZjavGhT41QbogNtZjo6Vsw4O3gcX8zd
832MyqrYk68DgSBeKi98wgZxRwSJJOWMgIe7OBjk3itzE9jziVuHsGzLhVTUYnjn
3K4SYFOeDEVwD40fG7Nal73pMK/J6lHzPHjLWxQ5nf/atDMVObsoKXJ6hKCu+hu1
ZS3HED5SXwsEWegzz9rAWKO5BKXxNvHK5lSobrZAkGvW3j430AX3iBrq8dJ/mTZa
rkrgbO4xiiMlsnGU9sdO5K3CWSPOhaCo6sNrpuRe6lJTbN7GBzKJh2yQ+q01BWjU
bjcS0nxt/AoL4Lyicw+/Ko5810jDAnQWhXclqbZ8R03pOGLD2C7PHRpBAYV0BX11
p1Kj4liqSAX/iEZdUKmUjdKXL7EV/mC1phfGh6s6vDgKU+ziMN3XtEX2wS04Zg/L
DMq1l2rrcmweA9zLtB7nO5mTb8CNSBIKp8j7ieBz20KHQ6GkC2+xgU3ne+nJinEZ
hrkG+dHOS8gSKrjvYeG7SzcshT1tsQlOs/7coAQJK9MCrJTqKzbZODx/Brt35Zgg
uM0Ladh+qV6mY6Y5cCq3srjrDqoWriJpsCec3nXdS+fL0u3M+TLm1WDsTDCxj7Uw
VUfWO9oCF2xPd3f9Sh+BEuj0ntwurNcJrq0n95cerrKq0yB3L9JBd2n6RnNFs781
tyYWfUu6Hm6qJTlOb7d+HoYx2xNGsyr5w4FtpyJElyqbq98BfP0JOfV4peQeq/v7
UUI6Z4D/k6LSwf1/kFWNjBqXzhsxvAPpvGHoap2sMfb1HkijmQWrdQMzD0yIl/hN
nhdwDpHzFLRF47EyX6Fkbhd3Y2iAaJqwk2XQuAoTcjLb14889qnrT/1aH7S0CE5W
Z4M1OoPExp625FJwrXZTI5YWfct/3UfWMmlRoxixHA4uJZuQGo29DYbg9fcSLY9y
DF5PL8MgeLfwl6KpU2yeZjE5uzZ+uIoR95bQRnWDpbuxtyNdVfm+b0HAdoFVT7oJ
iHujg41946IC7v8ywnn+NGZn9QkSPOD6mzpVvhyqiLvG4rbeeR31H0+Sz3Jj1iQq
QoJzq1FaWxmvH171iy2atvv2c9345zuW0Wl0toPkgwn8BE01+2cGNMKQ4smvyIN4
Jj8p9Qx7N89uIGBMglLPlpzPBRVtg1m+GQB4YNqF8sEXhiSQppVZ98g+/6UGvAA7
3fLXtPIUp6G48z8peyzdENRBp0dIGwWIHJ+hqfubKPmvrrky9s8ZB6RDAIdSKCye
9b0vccWhvnUO2ZDbeU8J4eYmV+N1fmJKEW4ITl7StbftKPiSm+QLeT3UzHqggLo7
Uhw+ao6EA2bna5ohjocoKl3c6O4JJZ35THDYwp6wmreTNPW/3w7B/HGW+9Q3WadT
K6jM+B4Kv5QgHBEqMNYbv6bSgur5gj+ty1ZEjqYC2yrUOS2ZH7qoY5Fm2357+jXL
bsfvEZobV4/nx0ifbGUWqUlpsxPcNfgg2aLHMOgKELBEtNu7j8UYHMvoJiR8G5fV
gbrujKHAm5S2bU/xuO1PE26qmOorsSvWLM5sisiPyjmQe6Lf/ImdjLYpB5zAro9/
2WbXYmezLIZE5tpf040Kh/5mplCbf99sb+Lsm+/2YH3jBKAk1LOndpnPyVvNCr8a
O/9U6gxQSh02/9ItAmr9VmbcHt8X9uLFpQeXXeuCVJI3KADb71ANP5NWDETzcN2o
43bAfDZ+84YohjR2vOV+rskvt36x0Tml2DrydDiQa3rDRq1K+UIzcOLr28Gf+peo
Qr1eczCVpogPElFS8Ub2ZLToXYOcw3hJAfASRgznP2sfvhwTriPK2llSJMAMTuqW
T40ufMnllDaW8vnRHMJVejKpMAFlO/LabHjr453bA2K4pX5mR4pYN90KKmOCMCUl
JaK6mtTqOsELL5gmy41vOAJ/trP77iJiyDdghLmt5Kbvt8xIldl3rmsFlY1r5tDn
Qflzyr6Cj0Y2Yy4QyCMFHs/JiqqjMdhK3O4oupM+6DmiSSWiTLZQLVE/xSovPh0o
L1bVyHnUR8MroS8dWXdgVvNoOlhDkaYZGAhPqbg/764Mbjm5lRVR2JdkQ3qrNVqm
iA/O4gx2WPWDkPSqKtPf2rB530gqvgXacmXx0ISQgGWlbDwmw+ND5UlOi1aBKwa0
MJupuWeRpCbrRBaFy1CxtnjMMwAi0rtdHpMSH1K8+FBcjnyV5yvEmySxmufFehMs
UuMRBu5ZvbUa+ut4bqZe+S1Jx4b3EpucgNmirFM8rsD2SUwvpyvR8sUKFXnTSImv
htyne3x+Jo6b2/844exeC9o7Eg/fLPBlRw7W7UcttUc8JxbhYcGzjzmb0/UGfJuV
OOINn93RYXMYR3tbzeRqCfwwcYWYafOLqyiiX0PDc733OeQWroOcsLK5nu9cSzXD
/Io/0FBYsZ9tK50MLn47TovlKAxeMN4Cf+9y6Lb3pJho6BZMvXXo/8X4Dtsx5cNJ
Kkj1l72H+hM5g40rnVWOMnKdCS5WpbmmQXyohsLp5kwkheqAGRIWKn4d+ZhRo4xM
OpXYJ3U/6M2KpoQ3FHz9JdUvycTTxyeq8AsIzdusVY0dvktQFQaZn7t5ZgO45S41
ufSmMshGl0sh6Fyyb/qIdXiV90KcnAmb7zYvM6R+e6p7nlPOVJH6bJZY32+UgBvH
DUtUYssES7c0uQzFxbYYeJkN5PIAWZcxFDzuCENfe2io+sjyxULNOG8ujp3H7b3j
l6OOMt9vjQDR0Mqy2A7Vm/e3YA2LlWarFntRQrg+DvwBsaapEkbJ/6VW5C/oi87h
4BkPMzhr0ahM/dhBKvE4mOdt7CBz/PWP+o5zoH8rTrNwWX+jnd5uaTXlpAM5i7df
o+GXGLpHFCVEI86Jzj9RHBU9lbty/fFxuiLxHh1JStW5pDHZcObkDqbMSnIQe1C7
X35/BZ0P9l4ZgPXKNVC1HfhkahSdGAwA3RA8ULnf7exBCQjmvPSwgZecRlqCOe7P
6sMT0wqfuRkszj4TW2Uf8e6mO27x6nL3+lgu6VKzHwBvqvwusa02IZBGsRoUlC/p
8Hr4iWZMABrGw8iMEFTczhprZ2otgSxgmIZ076B/dimc3wFOfnEnt3OB582D5YGR
/GqGQAJQne/bTkFcbfnr+1z0Hay9w48B+r1cOjE34QUW0KT1wPSlMSBVcQ89TbYd
Z24UtG/nj9PnbAJX6b6WUxzNzdLTgHZ8vLfvr+FCy1S0WjqpuGqVQsxDu9YdUATg
gW3mkUYySrY/S8ZP4Dm8piOFBxM+ddhghWhSRyWnnScoaqw8fokzvSh7gLjfAdu1
t/ON8Pd4eTe6hTDzPXS8SgkQsMDRiWmmE5VEeNf7NnXuv/dpLQcSEVBn/aeTFVeJ
YS0IIHk+E85GdOtgj778nNB8V71nF+KFu9VhliNXtZRfPJgRYjepovXo2tCArXyJ
cbMoVy7nCIGvFhdDtx9coNS/HBXU4XeE+q8OY4WtV4ZMMgVBS0iItL3JrcRDr96U
EuEu/8d4L0oqH6KwVomdi+KVdlvpqn6HIpc4/ErDWMphpaN0Rt9IMK5PdPap6seb
qbwlrGQIzuxZFy69geicwTW9zbAvBUcl5obsBzFpdrzE41amKJgJ6Qwsob5xwtYM
tx3GfMz3UEFMj89lZjN2zgtNyIQBV5cfSiblCaFH9wnhlrhWAygr4bA0fLJSgMnY
+LyGQvwb9VK3iZpsEV3prtghHWIzWkL7EaVlg52C3R56OT025mpq5MwqINh0IIzG
hsxkP+VzwW2oZ0t39pyPr9EDt11G72+JZByQUBHPAGgnNncZH3tyxJN36XK9BIvg
uxg3id1vugvPplQIQsv0GhpflQfZYGMqj12Q4DYUd5uEBfalU8zUmJdiM32q8hsi
QxsTIa6x0ltc/nwZdgGYMr4EnOB/TWs+8VVvVyA9HdmzLzjBHnx55SwGmyBJu3sU
7tXxg0B+xMXYROWF4CZ5ZpLr+bEQO5Tc1XNFc4x8PJrHrksNBY6uTkrhfse5hVtY
fP85rkrHBtwWPJhRd3Jt6JnFmxYoZbFG2fAwOsmYmoikLvm1vrIRmFM0/44QJdT2
WrVbPykJOkRtCNa00I0O1+Lzo5V7AUVpjHFj70FKVcaybCshapd7YiVVpmksfIZc
kseUEbJjqI7ZtjXYPQQBPn/eClZPKjMBeOwyTiVhfsDqhhXyM+bse0xDqJcvU7oE
4bHo9E3KRM/tYpp0vmcg7ZmvpAHNr/y583ow3ESaaIVpZdAHvqQDpsw1dCtq52DL
BAKHA24Kl8op56JLdHRN1s3FTnMl3fv7QoWH2KAUmDkHc5Jbx0/IgNWEYFmKjyjp
dhH5XNgnzGC83tROzO9fmtwcMwDGIVrWTyt8jcHh1TqEuUOsQJfw29jOC+Wh0N6k
qGAO91rw7bp0E6rek9VcX4XITT8gkHfR9McQxbixP6SEcl9NxrpbfO7D5oGgeb7i
jHLRUafkJIg6A0wtEUKfTYRsPZN/LnF1pk4E2V7OjdGKDHT1x/xWr/lYQfPSX/JV
gDINqKGyjXxZjgFfAnyMMDJ/gvPoQ+PPg1XWR8IHGMsdgWwr8tECnMNJgHvpFbc3
9NXCc7NZrzBeOKDhXT2z+SlSocOrl/K/mDbwl4Om9cymaAB5s82F82+FwkpVZF/X
sdkD6vfk36g8tR7jwwHkE9oDnr0otTbsaTQE75KgZPUuZFZMSpF4Ir009hWrKnK3
zhzyFugF97hClxMzD4PL5s3Zsl5XqCB2Gi03RdIW8NGtTAMiqap7rTUP3MynGdf/
Ec3dYql/Op8yGLOl3VrkmS/UH1fs5Ht3xijzxYTHPDBGc+kVoT/1XdEToTVqm/4B
NCKBcOVBeio0Ye86wiYVycD2MAgNp6YkhVx3+0nysoVkM8GlqqLdtiZvbKlp5qrN
0/7KcbWeqD34cwGZKVHyfEw0ZJmG9M8TkK5bi3KlsXBhYTNn7jgMjRTe6MXTHPxm
mvpUmrKEayOLXtb/WTLk3evBsrFdbdw1oKpeMWSv8DbRbHXC3gmJ/P5NGTEEPvTf
CAu/469HiVFduODvKz7TzbwXKW4y2QJCOJoSeFiU+N/4k48qKrv1yMYdhRmJE7HY
RKAaQIfNwJDImzZ+Lv8sIOD/4To56cVoED0vLXnp6mZj8ibkpziiuuoXmrfYzgk+
bUYtRXRWEu1irQ1DBZrC1jQL20P6f80QgoO3TmmfJQpLVm/NkESJFLDIPRTzePU7
hh8rsrKgdo1NwrEZuTSIHpo8zbuAWojcYClWrOat8cC/ZtMck91TKSpBs2Hvz1ZP
SCwiwlg3roEREHByDEgx1u/ZTJCy2AirAWklNlr/PpxTOyELTkclNH3RHthAi5ms
WOp24jNIyjCmMmhaE4RzafFvRgqgDFOLN0ygRCyshWJyPFV3OUjY7eVjC7yfw+qA
ThRKRWhMg3wYEc1beUrVJ18FTQTALTjtkMIw0B7ojFhdH70bImjlYdTS0As6iSip
Urx8vITCBLUCed4sOHIdP6I5FlpCCi2/4x2UTy7pYWDyGm1PXuvIYxSKB/+so6GC
17JSAcymHdYx08N4sB3Y4PsIJXHhjqWMvqe8PQ5CjE6r1jBdJ1xJ8TAhPzMjum1Q
xQNDwlIeW7fAhotGG+yB4Wu2oLRhLTsQvbC+UARW72iQDOnPgFTRnbBprVvcpA6W
QUGt+DrZS/Dmo1G9zAVkBlKDso7t4kVVapcGuwyqKIVFM605TRr8AjqcfZGVr8QH
gwCW5dBKQb3M8Gc4b6C2kDxZVI1Xw9RspZJM4OdRz8vAS1ESSJTA/n/Hjbgt8ge/
UyGmt38qkZUegcF+1u/vJyxC0UFsLtXzEPB10hECvVBIHmpG/IO85caCKwjn+RWL
qsavt7iDbrNDBP6sBHglKh8B8lHoVhv4IAR8mudnsGQ5gxI6kij8NUnPV/pujeB8
Ll7NE7U6hfo3k5ef/8h2oeLdULdioYZ/jM+0xvxdbn0oWKufUy88rziqWhgN85FC
H0S7/uzO+6qqGcW6MovnLptW6koTfz6SrHGp5E45nC9P+AhJivP75Zb3iVBwAG7x
YyLwqEI/7EGn2/3OYFJgu5kUW4VxL5xmxCBAFAyuq9ddzOJ3Rcw/tvm36chJdnbz
I6xSQie3T9UnMjN3VXyBUy9nLO30asxxD2yj/AnvikDHxNWeV4jO2c57bq+75yxh
yWCN/8lCJVu3TCalzAqzrzDO/lNshAM3kE/WyXyU9nxHe3rbkO4DfjiuEtiGyCqe
hSvJb0a7g+/wjka2x+Crp1zQfKLP+HMK7deynbXybkyNr8coP6uw5V4Dhxc78Jv0
CYWVwcVT3QdgBistLIV/ZENc5QNFweZJcglZ08jP2Lm0gkz3pmm9mC1+61w+1alR
Ta+gHVGBRU2oPKltTzHaaXaKw2XKMiDRIXfJ1SfW6c/pBu7F0bfWcjxZ/IZhgWGK
os6qVW4pnG1iDN1wdMRAIcI0bP1/wOsqbXsJX3oh2SSLNB8bMSk8gQEy9/dDu0WK
1Ggon+4OMXjuXwOBHxrwmnPgMrYtK9rthfaOf78CMTdskvJ3wSQRU7lAJk41w699
AJpJqytvKbmMVcc5POsTLp9/V2MJ3C08VBXUj8yZggJg6/LH+3DBAr7cVgtJ2fye
qekWgzuBkP0aV/f6ZAyHmoGBgWLv/m5MLJph4dTLGOX0IQf98KTKMkdxZ0+eOblp
YVy0mW4W8ApZJ83rmWxowWnYrYZaJjVJrfdN32G0rqVq4NkbgyyedhuSUilkL01B
u8VxSuZggLGgKN+ffr429Rc8wwesOcTfhvRtuUZ+eUrETWNMOiIMIzQff97fs0sM
3+939skGxUmQD/VIyTQxoiSmUcNSG8XDqbtF1Z8dejUpVMYJliDOrPT0tUvaK/Zm
nZDfJMVsEWWB5faHKLl/PJrxLx27UiChQMJJYiaRuWoqpSLS4zcQ9GTzp8xh+hMx
IiKrch60pni/S5xhZhYNqaziy77cXfr8I11lnwZf0NqD9jtnk3/WrTq52OARL2c+
ARFKuykeDVJhBgs3PZD1wDG9vqwnyVVmSmhzyAnQ6xTMa7jsvhUmsAOXhaYIIAji
aiMmP2ZrYjh4/FVKxTS1wHIZmoDdpfqQgb7n+fPKoZIKWLRMekOmCkkQ/b/1aDlW
zRggxvIpfdlhfX8Iksk1oxRasqRlIvSCAvjR0cKTS5vAMVI5U9Ku09z3U4mY60zR
b1GF+IjqYJlAr7aq5ukVv0SV6gTBtKJrldrAPe3AxhLeF09dVZNcHxDlrVSssXSP
Ro85FwiM6d8WiUm7IaNRE9qone3Nyt5LRUfsgqVJ8LJIN9P1099MHO01eBs0cTIj
SOdDWl3EU2PIhaEJB5RLtIJTGB8o+KfVBWRyotmN87ylncP2HvWQKIMhp0ETsLvO
Bcv+D01WLWM+6tdojW73W/htctB1Vkuq1CjeQkZKa43OsGYXF5b3aGZi72syxi7v
YsN4pwNA9zIOTTrBA1mZB7gTcwDBflF+LzD7XZEP70hGwgEAP892jf9cwsKw43go
r67dMJ0ucj1IPxs94e60W4pseRa0eP3xfDASnIO2boYujS2CQOQPN2q9OfXqvuF0
0gJFrlVWzf+N1CV9K6y9Ro0RITuh1P9vILX/XLIL9XNkuQ1mVUXOMy26P4d1FC9d
kGMrBTX/FbgHs6+LZqMl7/YRzfJhJyGBm0GpSctCPscsKfGhA6WKTy2vev7To911
2qdwtGdlOfKZ+kCaYKbCBl0nNrySKG8KaMvQh0McIqpYRct27UAepdrviAtFwEqY
JjIdRpBR5w/Nl3bWTEk0IQP7SCZVRVvRKkfSXBfKun4oeQMiAPd1BWDiZbjUHbQ/
BbTYy+r09EsYNVMsrTxj6704n9ctL0sp+Ri7ZGhIs0rF6ZnMHN5OzijEy7f2W2Oz
sNNjJ4/2dejtCWTn3gLcRR21ZldRIRLMuoVbhyPZHsyy9whU+ALhqzP+k5wOLHzt
RJYJwWOlHsejqjPzyfrtjAWC76MCByMJuzthRDhNk2NSnSa65Qm0w9dCut9mDgtQ
efCVmrPgLR1vppPhzvSNuNdmxBv3dumAVnygueF0A1dSrQEwOmM8/YKuOrXpk2tk
ES8+ns4zr7I8kMn3Ri6MGOanhGJjY4G2kfMQb0EnVklWvgV38D/r4vKnKlhzw7j8
bYqyb0uHLUqVQV4lX2Hf27CzacCaPYCdgYSQg21ghe1g1LaZ0CmaK6isGCZ4ipDo
qM645YsLfxWHBVpxs6UYr+QOnsYsYp6eAdpsdUGXgnlj93ESsPZQoIwsheH0eHIq
0fYPiVbSm3yftYx155p6IoXdhHm1ttWATmLNyHPO9VO/gNPFMdVtQCVLEU+HJRMf
VSSOP4dp3+li87fOxCJBoDtbjDXFjv68dTg2WKlDycgEHz7+4E5Sn6FXm/mfGjyB
MlmpGaX2z+LO4P8xh/QYLFmlW4KU5B8+oB7gc2dfKBlgIrZJgC+dvTXD1xn8tn+7
pKYUUHFNFVRCutixVq3N2h57VKmcS+VI88nGNNosLua8JLfDn3A+4CBR5WcECYUq
sp6p8ulWcjsZw+EH7Agoz22iDezc9rcZid7d4f3U+juNQJy1b6UOWp+UdCVu0Hql
Z7ZGbphsiuWB3gi6KtYqfoW1XNZ2BiVGXI1T5KOgWCZWy9YyTqMkuQKmzkJ38Z1L
j+qra5u4HEjVSvlnGWbx9QfZz8ZnXW4Vs355uTfDJqI2EgkAsPCL00PYBxbF60ot
8oX4+yWvZ+9q8CN3HF+LkQKfGNDKtTooKJuNAsGlM1unlFfFeLLU7fDcZbB4aPx3
xib69YCFvxGm1Ms1q0RdhdaiNFe9DlC1Zr6qpxAye5HY7+JW1EqCTu+IXmEMHm9L
nlkjOnOqhIFDupNT7NQLuKddu4GLaOLWw7Vbaw+NhFiRC4LAi5jXjz86LG/C4Bzl
S01aqZY6ufCkSd7FBZI5OpSJEC4KbszurREMplJIoOUn8iWeuPH7tovZmQGAT8Fh
btVPxCBIe5eEcIXJk4jlbboE1T23HPgO8saNn7cBvvR82OKIEaDe+z1yKm4RRKwx
nt/2l3s4YoEEx0wUwHFZmH1diCcu/BXJNN/QiVMjsmgE6tsctV1Wvi+uyPyqSL7n
C3xOcqPBuCOmqFQI9aMeWwFNzDkfgdfLQAzrmc0nBf2M9SwW7Jkc/y6MT2s/6Y43
6xUd2JRxyeVfuzpnVOYmdFg7MHx/7pr4DZ4Mfiem6um4CBfGo7+VCXLTezrQBJ0t
kxLTUWHYmkPSPL+QTozMKzzS412Ypx5xY+bKnV1h/6gR+r/Gx/UmGXtRNa7RtpUI
8qHkWnMEk5GBu0jU5REBJ3jRHRcS0kYWWAbXSz7TidGHzb6t0RBDuSA73isqVnEs
YTipu5Gc34nqszlGj8Q3JTXIttXKlmPPGXOujvDQ3KJ+Y50SRBYsGdVcdNdgks20
ulhgEZh4kbuXMyJgid+FstTm2c6gnINdPMlOl2qMou+ezESk7yt6Jon5RYACX49I
TWsLmScc6y4OzJyBjw+LM6rflJS7sbF1omKraIL7JC4g0FMvCMoDyUOoZtDPQqj3
ngiMK92mftBGRC3ACQp5TRcSkRuIIHHpM98bGC6mDEq26mC4k46/JXhXTvX+PD8b
8viQuV+OYRtYfLDpSeuTPfZwbhtFsMmrwpUxF24Nr1oSr+ELeUrCdhj/GXYNTN/5
CA1ejyQqSQ9Ek775Ksy3/7ji3F8cskA+lrFKSMOsHlGdNg1AIFORcYLrdOXBXHEq
UqgVpNTkA180FLRAjfllwqbnBf9dICGYHYipDd8wq/F8W3g5ZWtsdM80rsICHNMm
GlumYx1V+o9c/1HiumkJ+dMP+v1TJnqfYjbllIctIfR2hMJWjLE1hFu6y+IBNPvd
fAhWaO0dMWB1AW2knbsBrCLFFMHnoG7Mwdvp1rL8QCce9U1XA0e5z20rbreJW/WH
ssqgF6Wgfd96a6cZZkT6oVhv93pR50iZpCVNofrM+NDn0GthwiYB8igL6xGtJmqP
oIwUrAT6aNLuZBY8azJQy2HerhpGqWMVaFsivqYYxReWaxcx74T50Ybsv67J/j0U
1pznK/miowrvcgZ3qzNFHLgmWk6tPQMcEueKlGBTuq2fKHWRHG5/kFP5/vRYyexC
6Z1+CO2WqVGGjM+a3nygOSL8B9pZEUesNSMvCoTWRk4pppykGtZlQ34M3FlbBEuN
67nA/RaQvfzziCs30h52Jqpfc77EYs7o6HyGRypyyAjKELx6i364pnAXERD1z7eH
y+t8rKrji5He/b57+tCRh4q++m5pM90iiFHQxaadhbfScoo86Eef0Wv0cts0MiiC
nHQVT3zF0MqaNNi5w7VwrLAC1eXe7fS1Rd2aHs3KBfwyOkZ2Wt44eMQ+FDJUIsd2
+qGBRQ5xXRwPb2VvkuE1mVdnj4t5bLrdfnv/ro8q+oHZmjQ3zPi/dCWOKrE2ftUl
8tY+bvchGIXLhuFpCfgaDpKnyymQDFKzRM0WAomixiRGR3tPCrqhuanryznuEQfb
KayhBDVqwCZe4p2+F6Sh1YvbNcC04lufKPvrX21+BofQ4jfnCvsyMryIrvGPH8LJ
K4kwvw3kJvgYJH12my6NcPVY0N9YcRhYRL0j+IP/xzegx/vLqQKR7wvNg1doBHV4
oX0NcqhmjJrgqOCGiuu0uJvpCniNJElSlBiYUw/gLyKhkKJrspUtIWjA/mDWbw5B
0xIHjhLs90acb3Iz2GuHr1tBEojFHRvEvKYM6pwOy5nVMzuZptCydmAz05bzDSNN
Rsm9RrohM2UJwWnXxeD3KnIBhvF58lOOEgX0wZgC7ClFGChY6yKpNEDEYCN8mLyH
l/dxu7Wem5Hc6iSx+/xNGaWN9M3ye3R5/jJvZ/UX2l5DIQjmBPkiqLDBvKCDAvBo
YF21XYBfJ33D/cjplcNaPkTTfStSTEka7+qWEU45v7cER5rYDYCFxQQk6oxRvZiJ
b299/tNPGuQIt0VRKv78oS3h07trU4WPVJj7QJP/sLQHuzq1t4+SFHc+dILtN0gJ
mTu5U0Ms/ZaDDofSeg/eH1JArAytY2+Ciotafl2WGRq7fXx2TH+lUpdhIUJ3Ej9S
1+L0pA2e2xe80dcoTGPlSIpvRRFgcII6gs/fGgbXdt8dvaxFDVJIb9Lu0xShxbTd
shfaJUHbXfTjPg8FxE2LYqysfi6I89HOh2hQKAk7L7TN76ybHX/RrhR1soruZbQO
JKsy/EI5pLi46tgaUXW9u1vCWdIyeu/kuhYNy24KWG+4ghn8QAA3B7o/4+mBWrCW
qzHJCKcF6QfSIvBpfVFQVaFJArr55B34nXm31VAiaJU7ebajTjhDPNFVCEhNMmf2
pIGxp3SNrpSlxYluVYO/vqafvar9VGs3RGRMcxGyPvxLofTXubxoQmSOfe6YkZVf
Q7tA4sUA4IS/9C9Dv4VOFF80UYVBUQwsz/vzg+0ffbyfp3y6Boalcin5npRnizNu
NbOjgYd+eXA986OJlaVE7nAf0gvXq2VZZ/Eq0KzU1B/tgysa7cxzxPHOrpRCmYXj
j5kGaLU5E1/IeUTlJ6MbtRxwLdRy6xvQ0fAIJp1f8nb+7bqAGzaTSWbv5Qc0qrIs
8moGVyBnVG8Kiwko78Da9pA1LyXFuSjM0Yw7NmUYW3vDGyztn14GWKEFo0kyDkkB
0WkFBpruWS7EShuGG8mWIRQ5D7IdaO9TrlIy4fm3werurj00FzcqxdShYN7NCS7C
tXdAeLRjKaQr6xqjh9eIp7eAHo3zTtaXu3rzncvYkFMi66u/OGVOgiBaC24KwpBE
ka8k3nthafXrS3ziwmJGs0s/V/c4NM3AbIvQVbKCnn8dbC01BUiHgxnU2hTZciXd
gYPZbx0ZvMsS+dScNmkdCDzmlUgWwZ+AxTGHk6QaQG5o9BpR9A2Nx07iN3A7xd5+
OdTBQyNpCrAbDxLb5tAXlgU3Ewtrp3wPd9bk3Zah9LeknUSOBk2B5fLhahj0wqrO
8UFRNTVC0mO+Xky9bI09bRDYb3jVWhGc9DFr2PZkWl4rJPW2z6Nn5n//g2sV0rsc
PJGRL6IZ+GT4YJmBYr3B9wT5/OWPI3Pu7CPFK9J2MA+SmD3Rj2HCl4tA5OXezSPZ
EWM5mn3IvMjPFi2bcnbxJK3wRPLlks/xKqWcL/vVK7L2d+A8qhBYdQ7CP8o2z6cQ
6EyaI1cBrpy8qwcjjAnQBNLx4IFrgmI9PxcE/6OYJ5y2S/ujJvXmKGcjhuAsbpIo
Yq6U+H7rSlxzBcDzE5vVJ/zZ3+hHXBS+hJYEcSONe/RlHVBHxmhsm6p3+8omE0Iw
EqttJ0bfxCu33H/Im3PS0jyjOiPeINDAd1bD9WWxYOUaoQLuyRGF+abEER7p+C6P
P4JmIN6ReaAJ6NIapkYQH7cDqsawrcs4aVmBtM/RMTx4LImJG6Irg/MLF8QxM/yb
wOyJl8pMbtFBRcUStO4p/jzHGtDdNDfiwiJlB6YtWU1ao5sqetYAoWjXtIvh8FdZ
QGvqULWemorjuFJfT65keNDBG59cA9OOXdZUvvldfhU8Gh6G6JYjPrh89/uIIKSZ
ZBOGb39nyz8aI9l7q00selyGqz+9b/Z2/FL4Pzim1YPQI3Z/LJW/CSYpywc7pZsa
HrJAY1xW7Rm5HUkpxQlhIFbGUOAtejmRQTVsPF5GrgAZXRICnSmgMM95LWw1fHn9
pn539uAqFazsvEKD14pKX852OrDUBYhyPaZY/BA8rxVg4yeHDVyHiBNsIAFA3kyr
czqGzc7MHLT2KcxOU5KhftgmcxehrBLm++sEbV6OEM7zSNtpDjQoKwIWtZrs1ytF
kGl5dsMVDbYCwf564iRDEnPJP+BXOa1NutBHptnTt5nVMsXkIKi5UXANXYpG5AXZ
53VPDx4n5HOw3CEoHAIrlzLdtslvJX/HEG6W2uMgsESefupuLNJlMauaoLvk74u9
Ki95kQ73+u2n8UcHTnDemEeO5129EE1UXhbNgzLDWvOGPxqlr6/DQefHmuRcGWAI
iSc/9mMnwOuSpJUF4KBHzBa6gMz1SpjXyNQ3YF9dXTt1cVmwnz3ypqWb9ofgvZaZ
GsJMcIxyY84XdQme4Md/qhDlJs88At2lW1lQHRExixJ9OTF2wD/DDXQGsnLqlvRZ
j/pFY6YiE6Bv5ZQzhDZcB3Jx8AytOcs/EtUdaTHQEkgazoJw1VcmNwD+SbAWlsni
YEyRZQTbzfWJS5XwidANdZJwmNvtaRkqmnQYElRcwjpYy72clKFzofBwRucfCGM+
xnyGJt63ifdQegzGpjdbZvWxWcqMntclz2dsYSSlwzV5naXq4UNoJm2J8n9f1fBQ
cdy5rcxHmdzxMrOCmqoQdx8KlcnJAAdfcdE5u02lVMenM8L5jiz3ChRObNZgnGle
rNQ0gqFnrMxgq4CwX2UUIwPLPTbmf4F0JGCR9IDKHnvK6yX5uhJ+nsQBAMICzftV
/dopv9ryxAL3vfkbF0RrGe+TSCEX+6+cl+a/eC4pNrNzzBL3iCvE1No/HUWiOVEr
FMMdUJb9I1Ze6tFpOJvwspK53Tan2EZjq2sBsj8z7TK8wSQTyusnPpIDUEB/37XW
Zen7toto36e2A0PeW3GFhD5oAqphbFZeP9qi1Gw/0H7cuSRBXlkVQu2ec4xA7Xgv
tktlPAMz+/4uNrgr3xgvMmkR2v8Wu2zkxp/cUyA35z5WJGTP73i/G0MgLrj9O8+t
WFzFUNby/VxvevPjiEAieXZewDPEcXdPeA3OwY3nP+bn1rrYpKgSJ4XjoTACY7Lk
1c0etEfYDdzzI//DL75rYlATivLLibQhAJv2SQMaLo+Y2Ui0oYVMeI9+1TkyE5ml
I2GMlT13N8Vj5QRSXPwsSw+97O2mr+Vp10eAb4anbIOWwsBwVxeOFwSz+asPwY95
4mdFDgd33sHwQc7Sm7PB/xYY5wDrtEITvEsx3a8cCRKDMIwDzYwF5KIrIlVATRlC
Ja4I+e0RyhWoophh/joRQIwSoo6i7D6IAgZjdaaW0anZhBdmtDYrmx2Yg7/jH/mD
F6ifwsg7NLS9eP384K5KFUi1Nh4O3JUNZ11PvUInm+tVYbZhffjZGXHYsMU6tf5f
/LCRR/72v4L3FDXZTAjrnbIAW0CWmgKXhlFne962iTr8ymqgjV8IR8X2qiSxbwRM
kwA+S89ydlnFtRRfFoiAop3i8ZcU8uf+9hGw/Fg3daX78ivRN2uxK1En2khmBB8q
hRauSuIJfCTWl650k+grg+g8Zxu8vckLwwbPyWJxHgNzoFmC3lF/m7h6zrCCF6Dr
07Jw74LbQ4vmWI/EkHg/JzEsxNvuS5oaxQa036KjNO094IM297TETov2YWy29O60
Pye8xHNjpQypuSCkfKKo4eHrarep17MEzLLnDQlNNsFUpcVdsbZr/+eDRFC2sX7Z
NaQKZ5sW1PK/AMy2apDd6ifMSsYt6nZ8G95/FQzqz2x3QsbvZSSW24B9yCteq2sR
rs/mjVw+Fi+A4F9INn156yxW3WuGINWUr140pBrCT44VRW8gKOF2dlWRbzpN85j4
1HLLuVLot05PJ/aaO8q287IwCJ41hvvX4i/Eca+hu2D8V3JKb6Tx5P8Zdw9bPKr8
7wMxsyvmMANcKBSnnwy7xWtfuHPbHPwdSTs9QL2YtzIdRC2wtPzTJvYfcXpP0qSH
U8IPmOAERqMA66dijyAR2IiimOQgMfmwx0TEZFuHfs5uT6ao5EDq5Yx7QBuXKgTG
hQVYTlCGBFgpZcfTLe1nbl1D2LYDinealr8GCBBle6TJn0iUQba2fYSH0VeLVJ2e
x/WmP7XIINuq4A4oNt3Th5Cw2Q2yT7BkqlnyzAZiD7k/tKN1ZVJHkzEHdyc0Z8Hm
YMbBpyf5o/s7OB799cTrvb99ztnbVeSWK7PZxxG/6EyLC0YqgvWG7NvYaoaCrUKy
Hn+PmodArXr0VX2V+ulqiaMksFWTHgMbuury2ahElrINwwLW9T+cbUzavz7Zh2kA
nMVaQlzart9tPwfj8338IG3oOGLPJpw//o4qxfG1ro7h5w6m0Eto9F/9hLzAK3Tm
58O4Jdsg1wJvL26sAd47Dtw1b8psTNJESaP2sevLHePkVH3ELOY/pRH6y54xeCo+
+AdrG6QrAh3cB/nFoXFe3Egun+yb98oMsrYJqTB5TucGvcICprzN8/TRX28gfuOA
yr7Bwn2apIYJGMqMhv3tJKkGCs9GElVHEycu1xq4RSmWA2w+b+Rb+2DFOHcbbTiH
kZfrsoie+FhpZ0xgyzJET0w6OJZRtIwQ1pRMEv90/eVXqYeGohem7fdLNArzu50p
482Zo60PCvHErnzEBGhsDU9pZCsqpG0LnoqAmrdHF4vlrCbkyAQ4xhP6T4EUYT2m
CWQQAHFatstvPx5kZHep5X72bUc+hzpbieKVN07nr0MRY5fv2qPHpKq3WcqspJ4v
3Q3CpnCWtlrt7HZ2GU8rTh491Sqe3RgtX8AYyU3G3tPxi6sZR9Moaoo9CS5/h+hY
jpCLKllomJXq8KkKEoD3uim7kH6QjD1xr/LH6jNpePDvlC+GRKforEcr9FODuDUz
P3lOod+T47bo8902+8D4l4itHbtZ6ZM8NmXOJNmpR1RNVKVJ430eblBkIxpTAO4r
sKgSF8mG2wr0rpxXapoD/qA/i4S4iLpG43T/B+7oWSA1Bxr7BPiaIc+slBfo4k71
vpz4qeFeaGmZAh06mwdTqYcltaP6J7Fcmr6337pgfPfSGsqKyQxYP44uBXF0CNpj
PstyW2geVuxFEvmAlmLPx7Ynh6G3zDhAH93pqiYxomV2Q3l8zFBrwKPiza1CgA8f
WEYcISESGbV3Uf+BGDUwEpWIr8HwwIh9QdpOrJIXeSM8v4koKC3gVkfwYyVmmYZL
owMDPibOARnRZt9qIZEwPZUfjYH70n7rZmrXFnoCkjIvzYGzYIqeEewS1DPV+QmB
w3xboTnE/HFdRFA59vtkWfrRaTAdm/QCGgAp58+kiD+PAu2l0IhXa2opUvEtIK+H
KZZB4JHwCsXcoQBF37Z306waI1UVUU3VIxmvTdvnJ27Bh9GeQmuK3nPQopMtpX/i
DXro0TxHYvvciC1IcV85FWq+Pab7Ils9iDo+D+9tgA1tyfzzWXfs0ili/w8LyHFj
FdOh6fGXnp2iNFVcWVHOVJdQJEkc8bgsx25VR4YwLqTd082pWEHdp35/UxDV70jc
MLB9l5nsabmH271HVNjixNt1IxLN7tdIWKEw3e1SZ7t4LtE1fi+gzvy29ajQ104V
negxvXhV7fu+hJzh5dxFIlBRTZ0KR+GgmVwwgokQ4Xl46ClbTLPSlanLBiqmaiYd
B3vvrLCWMleVoZXMu6CXLBxTVfY1WiUk8XzlIKl6/wSfY/OO0AQ39BabFKbn85Pc
x8VNxRZvFFGdBQx6T06QGuwM5kZVUxGCYBcJ+m/zMReARr1K9jr48Yc0iL7YNiXD
kj0CZtAgPJXlncPy9MLfI6LBI3XPqtkNJtjYyRf767//bA7lsd/u/ez+9vrsnNc8
l4I5jb0mSAlXVBdvQpVCPXc0zp2ykqz2iAnblbZcMAReDGvgv8s2PUBshbldkupU
TdA6wehfNQc4AFyFmstu6rLHk0FJApzx8a8FgRhdAdG12pgsbmbx+9F/bhpygi3z
hdLO/3gmFAx5l9Me74iQP5/86jZdwY2lQ2w6FnvS/Yo336ZYl6rPdjq2XDTNS2Y3
mmXkq+N8F5CfM8OpRyKtfeQe2WAt7/FMM4hFgu9ug8c5uzvozO/hRQp7dQxh0ll7
rQGrjQuUJ7Ijr59NCtNiTJZDO3YoruBdrlbqoCU5RE9r8Kxle9VpBMJGTNjTlwox
WAMDaf9sE0BH3dFMH+Sao0E6Gt6F61WmOz2mbPMZKOZl+0zvKkcfUx0l0gvS1eQ9
+7KuYpZIqP8//WVjX0DYed2XR8wLK/S6L0L7LVDXrHQDOhj36sZu0r2llOeWI8Ay
LTworCnDQcvarlhPIk2pvezcltIzBnIl3OWgyOeoUMArvT0i5W/6siCELkwKHWo5
iANYKfaI/7ZkyGXeFT7GgcLItfMs8HcMMa7lj8N/ZlcPPgTn1aw2Byzm3CLgnSJt
u9KDAKGt6FNmJHVhdfWnSZcPjGuB8TZD0C7/7iFQQynuc1ji//kVnU6IUvvaMF28
rQQqNLWJwXWCA3R3qfygKLMtx/pk6Bbq6dCZyHPHCe9EYaP7lojcEef08cKoCE6H
W2K8FxOxAi9WxXo9YtPDRwO5uDwZxZhhjY8ItXRQ3Nc=
`protect end_protected