`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 13312 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
mvOv0qUqD+6HYGQ6UGdqrf9oeDe49grobbVyNR9DlJ/ozJpU+IuOSkM+3DkpvWkO
0tWB6EsbCwShPAXdmX1WX2GHDts7iM23drZUDYA0el846BLZJoJudFZOIFcqGPOg
HCFADEY0ucpjzaFMMTCMiTRYbbnvSRe7JeZAKWv7dE3FWqpTqi0ME5A7ftn6SYYw
89BCYE25oeDk1i10gMuMeZ5r/SMCsiij5vcUJhNKWTkBg1t8v5wVHQ/3DlWccjCe
ox5mbqWl05vstYFSYuRMV8WSwOS57Nv5VQ5iSo23CtRhnnX4j5FrUhfgH7BuctUs
djK2knn1IHMVlSEacAN6yEUviKaK21kknvJyos6lDNyN9upd7KrkDVSiRV8nUGON
BkuhLNzy3O9zv9gRorhcTyONoH2PhlSSKX9t+DuEowkpnsoZjx9+9ryGknIq+YS5
ofSApUMLwCHvxjs5Gt3mItLA/1K0PhlftdXqzPhVb84QQfiMYLwT55FqoFqCYuwz
7a5THJvXA1/4qMkRUap1qFqKxd9kbQLVV2pbPDAG5EnxeEFVTDDX3nzU3oa49D91
rTCvMyiDnVVowd6tdFpCfhhzh9ubM2LwdWyPNC3Oy2sGKZqt3JuZ07elndaHb0Dw
lNWkgUnZWY2YknXcKG8gn1ciOoGiUauzZsaJ2U/e5/fhV9gadt1gu+hLVQ6x8anJ
a4OHkQ2VaSIuJ1/VUulmUwpAjXVvGGBqe1070AU6jv9OJaL4YpWNUKW69pIOGeP7
5eYlibfLNDWeEDEPT4c4hVgxie3yXaxEUd5CHnypq35xp2GTE2/CZAfkYo1jYlcN
clcDdus5qLW7wrEGLTH/WqFRMr0h4oeOE3fCGLuqBOxOHLy6FObpwWA8Itk/3xy3
19VlHKGWYSFZUqzHi9gNVN8HKR31K7w9SMP8NYNI3qwPapZPJY4Z9wHnk1/o7J6i
QCGH9hX0AGmGWc4++2fvL6AhHUDyUcOS7QH8P+7BXhD0NQAzmf1oUlYqZsnJIdZV
QT1svjZSIR+7292O7Hhfk2CDQFr6IItiyYESfuTWHssQg8h9kyueUo74uVrXu/y/
usQPe3bpDpboEF5Dvq+2IgvjPGRBj1RmxEYYQ4gbMZAqZPqVJ3iGJ3utBTxRcuIi
P11OM6RdNARaoSQsYRqoqZtaSac8o1Pj21C2oVzTk2Kw8ZDzRfWP2GDhc72K7T1d
pvi7RYkev2tfTZ6W+Lr70uE9zECMQg05b+I4h6e6OkGlvM/qbmIYwhjIPseCKatv
/906tuC/TMu/99qoiw4nW6r+EM1Jkx0of3H+tBjUZXYEHJF0jYI0ITNI+HWzNvzu
TrXa7JRywj832+tPwXSvuAo7/YYq1O0WkESLodOzL9SXGFVk1ulsex8CH7Wll2v+
dQYz2egC2tGzcZXbDz0FuPnSFNZq7VrA/ZbbTn6LqoKe9UgEL2mUhvXPBbsh+oi9
o94oHkn02A83InoHcnaopcvQ/lslwRuN4L3BC/ZWIkqnuRVG1qt/LsipAbFXvy/X
Z17Ga5mTKWLqOQgfKtMDmqlbfkAlErj8dXZMRyxGMw10rPiZp4frGNc4UDFtBmAG
rpci+XwYrOdtMPyQ6jJHGENu1K6hK+hw1Puaa5dz4optjW23LDZPhF4rMLbzzJoW
ZelXVbXyso8yNzqSdlUP0qxtWmtBK1sDml01E7M2R7Ho9ne12AgJbPb7qyKfXmKB
cm3aOjK6b4uGZ+eRppNd9lhARFe+McOkHbXPQDmz9+XLszCZ4BRkKJifS+zSwQrh
70GOerEs4FcY/Ks+kzZJld250bfEkvsp8WWe+4WwxLIkh+L/O2tEegiSTHEFv6EK
NeaQ7Frunfv72pdZBEVHXsiK4FSWD6pHqo3yWY4Ey70pu01DD8ezk+788b/vbS0G
yBGeTcY7OLdCiNKYz+eHRSQjuya894WMgIabo39O+lGcF/h8RVZueteS0r7TcHzL
tLe2Tg3Zamv/C7HvSqmqUABD/CoguyAFqJ/zSoHfgVEpde3dZLzPA8EKoVszzLHT
6QESmh11i4eUByEQHs+9gcYNnCh+3CCgFB5K7YCflIc6ZaSWPJDGo051sazLJCUI
IG46JvwjMiFIQz1vdIoAc2gMki4BAEVZYgwBr2gV8NRgyE8vz7b7sUZrEgwtCUy1
4VPZGktgj0+6ziY48+z9EWgRpOjj5octNPHLrVEKVWO/QxiUd+rIoicTfcCEqk6F
+hptZ3k+q13vHfJskneWx65qt/bS05/GnC7PWI80yanKbC8/kquI/omEqWySCOXp
mVOk/FRZbzOSDGFOdTSV9h4jXbeieiVqRU2doSNAUx5pJ+Py8g3pqX/VZAHAfpnC
UYkwdwrc4CflX7mMGNvVQSWGRtT4TmWQIFxNaaKiC9wDkDkj76JEsZxgXsXgKuGo
2TsHsvEkqOL5HJ2+mt+8DSk2YBVWwPVC2yXT+2XACthFvliksZPQ6yqt9xQBjKRG
RNKhRQbrQ6k6M4yWBJdvPKerVudhCzmkCPyuKh6eFpUYyvZu7Rogx/p2Id7y2MF/
EwDVj58XE3tZdHi4+tSCyB94Z2/J3moU8QyN9EJCDkbY5i9iyYb3Bm4OEMI+oGP5
K9g2qBr/NDc14jUMLSh2NWyync66EfjPUh9EZOgjrMP5UPgmxQa+WC+pw1Nko1gN
nh61TZvoK0uZqhaIl1jnUCvRIHnnfbj2H1OnTcIrX6B/ORSX0s6ZV0I9RskryILj
Dr2nTD2SGPxlJ39ndd6IbccCiuTO4LD4fGLScTylr/yueDZTewCA94O5hg9OvpFs
XkZLeVFQDjsBFuXcY4D7j2OHNRtuC2AgzJ4+Ql/eC+x879pMwTVXvfQKuOb5KFpa
Z8EYJDRkr7oxAhqDvR62n++uJxoveJGaf629KkViBSwSeBo/3qNUUylD+DeKVYXX
ujsonv5KNwTE6XJhHrPyNJWSF4aKHPntTKVqguOOBriQIWLSQcbymW9fJnzzbXSX
9Ljdf3bwesfAsFeCneQdFCKDzloe1mK83/6aqUNWJwqSIyBvydgjefySilJoPjSC
6IbrRmvO3N4NVE0JnWIl62/HSq81umkZGhanAOe30EmMewoF4G/XrC37GkIDztHt
0yEmox4IiGN8BJRBEJoW7pJAupvPVOlH2Ie+bzFmrYXadX5JPintDSjUSoNHPgKD
2o15F6BbUGCefiBHqfwxYhg2Xr8tKl6tq9sdB2QJQGlRJ9JMFpHc5ONE5kGF5xwG
ugxLHDtHKq4flDEnYZBbkEWS1b8FSE6fLfL5rH1xvadXW5vsmhz8rlcACxKJdrbc
L7Qk3IvVNcualxA1H87WHbljNxT/EYbNsPoovT5GT1BuIUSpzyQoE+6xqt6ixw+N
oWwKtOFd2LaxpHRs+pnigl+EN5o6yEpfXsjakZxGPoWEp2+mCIAVq4GmUvWC+5GG
UQ8F65Hts0QdfkLB5NnyJ9hKj+S3YJ2xRGEuVwYCrn3rdz8RbGiBVCIXAV9O0Gxj
hL5Sl94NRFKkRpN4bRlt1tI2JBawfT8UXXW9dxJTtL0aRQ51CqTzuIqkrc0l97eK
Z5q3BEoV6VIDnF7lHZnh5II1f1LkVeL9KbY1LMPxCv+2h/ZSGFemzc15xAR1Uu1U
QanjHevSROOuPJmf8uDtF7SbL+71JKel6Q7qw/tbfD4ulmuUz41x26y6ujTppZ/e
f3KNB2WX7KSAQiwJNdq8VXg3v9wiJgARRWt9VNTaQzIpYYZL3/c8RaYjXPGpp65+
OXK1GpKA+AxcjSNnKziZgHRSW1HxT7uQ3HfPVxXuzWJBKLF6tZTMIcdVDTBBGc+m
dFhmPUbnbvWw1sw5SsgeEqblbrZTUyJBA9MLQbaCbYVNBChzgNfAkafxhdi4oQOG
e6nfT1CTCs9IbehEj/FozsWc64/Pd1fjw/Hx9QhFGbCefjFwPpaNhDJ6HrAy4S/N
XLn0ECUpDTYwU1eW9QXJ+bvCE3KEwMBq/8kID7Bmx2R9Th3sYrZkFTAa2wNCQYqJ
R0Ir3AtoDYXgoXyA/F+bxyXcXkFY62hpq6pahV1218ObksONohedlAP8vmLDbLTp
dNX8Sc0Fzc1LbdwMDYifziWXP/2g6iibFiMjF4KzPnArRQKav0lpXjzlOvhORaA7
XXfh3mmQIW9iclRpmObuz4Abtp/zpMop3t7rxCHFn2z5AZGMzJCSgXh/hI1NTNGk
6vmk6fU5xjdw6pc3rUjGBU7LXt6szoyR2o5C18pGqhu02cDNlxID6og7Y+j6Bu3q
fx1e36bF3Kutzggrn/b434p69/jfQe4w/CxgpR81iO50ClVuoztcBNXGqD1q2dW4
4SuL3MjoKcpjSdGtvzyfoq1rrMvJcO0un4TYx2RdeAJOgIydr95o04HTcxeQH849
fZ+Ijsvv20L0DdU7lAMFOZfAwLxmeIMeh4cDT60L9Y8prfxNuMykMe5aMnzFXRtv
eQ8W8lpBB4NeyhH5XmRSM8twuXouQOCovhmXjVXct0WoAEPs2FCmyubSrsnGiOsK
oBSEnuAzTrZgrr26Y8edgbBysL4s0nmcd0smbIO9d8ajQhgi8e/JNXoKki/Zq5kD
2s1yE5XeEGQMku7sgY+2IqBr3WqWAtzKVzCx9Zo6y7jUnfMvVQ/M3GQVIVU1T0Dw
jSY4y3NpBa97kl/TXVJWoXvjpN1wZzB6mJjndlHqQq4Rq3zUfhr3SOAMVosYJgKV
LwXsICa0K47SrQz0h01rgJLFg6tHrYyP4UCct0gth97ZrfUtYOgvR6uc4a4luTdB
EV7gnmmu1VrXinYiVZulZnq9ATGrTvtCKyO13MBcjxQJRWq+ZeHIKxRmYTiM7iIl
jengUtlWlio/oJMiQUDp5H3lpTJ1BDrUcmePTYN3enmiHeVoNlbSJGsrM3DLFEd7
FTMy2XWLqxzUG9pGayk+WxFYWITtTi5003AkVgw/PmS9Ez15hEjM/tsLWgPYvw9X
vB6oGuUptKr1d9JLt7NGWYEBu/uDankoHGsCRM4vYdmJ8ZpJz012Bq8chWjuzOr2
VBVTnv8jM5J2TDCzcLfEqg1SPta6J0N9EXZ/4BpVejRCsmxRYM6YC/rZfbxNgzqf
xjiUQBzZLHJMPV9m5fCYVXFQR+wkMg8wBFFjGAL7IFo3iI+/qHC1k4+JmXiAPNGp
cED4sHeFX/W2OljIYRf0WYoZEt7TC7hTUSeLvzhun6vTplfc6Kh7HygxK4e+smuC
KVazOwmClcApNox/laN7tpwtk8uYngxhD4W9NDeTWOqbCsSJw/WKRn3s2ZdszhNz
EJbLarIYyT0sswI+Mjq2y0NNQ8juMXtLryxI1a/AM8D91NJkOFVirqxYSG1OleUC
iFZjpXwm4kIysLKOkOQtfVif+bU/i5V0Th+SssUAcA5L0LfwEO4iCrKclAaHx7jX
vtyFSLd6l5RCLhTbDkv2sKdb+9lplwXv3m0sk8RmXqKUW8MBFMnp9ARWmURMaic3
F5FH593+b2bGzS6shqETLzV/2D22bVFxRuV9ZW+7LQ0lGVSsKKWKcrTUv3e5qe9/
nQxrb700zvXl1xDX7A/JJk3Gujc1tqwfA+rjYiuYrnzIS5VbEC4xB32Jo8Zgb9d7
KyoDzWNuRhJ58QzRRhy8LJWqUgbnh0fJW1bXMDRh8YywSd29sl4MzysvSZ7T7u7M
g5ZQoYaCHb4poE2rEvW1nfM4pKe1+U9ca14XFkph7AdwTHWUKj/KdF3QliVAuJ4q
rs/ntdXjaxIp8+rCFSd2HMWiN+/DVP6IczHotypQiaPz4E5IrMhQokngJ4RW1j0l
8ns1AYkcxLf7tUUSCFaJcQUmOUr0mMiQudD8kaJtdsE74WVah/XTVgZHoGezfBCq
2uzlUf1uDWzq83mPJWqq6HxxcG12f0SdrhOfO1kAi51/V2CmjZ867pUIP0/ATA+L
1Snlx76E8OJJRW4G5W3QF5/vF5TYQucF3Q5Oe2D3WAuQAftsNHooXl6odAIn3+H8
NH+ZLG0bPWBYEQwaa2PccMnqKRr3z8+u0IBE3c2NC85rBgVvHslpfsZTqSKU2d2v
sdheZjrHw0BbhKFgNEucSjiv98iBy4cj9HE4g3nWB6cfMVPVCFbVIO95cCZhmqTJ
VDRXnwzGOfrNibKRrR8UTmUgg6RwsdZLefPmKIDiguVUKmGzPVLpynZmmoh0nhwU
qV14R/0RQnqGlBNa5RbedXHZ16CEu7mBnZcGl3ssRcehUxSXlCQhZQmrnCy87hco
Y3LGU1OhEgDLrKWFmwr3vTWW8octZx4xJ2ZftMJyDj4W+UoEr+IjExvBZf2Ld+IP
KENpTje1BjV3Jpe5VIrRthSRML69s4NQ4tat19wFqBIvatGFWXPVkS7z9BKF92B1
3OPgjnI6Hv+BpSE/7oAUxGv9RBP65o5Scji5FwsJjAVYwRhi5pnejVeGxJJngQhH
rgrPTxpm7stHmRRtCFTFFUz1l0ng2VPnaGefp+98JVGZLiTEh6N3OPCunfFXTlQp
UsvDbtXx8ncN0NII8/hCed/DSKCk14ubiI+bqSKevh4OtOimgLQRHf00ka/qIq+I
y9erd2kBW5ai6+Ies51RTCgemc17TSCtysL3SACubeVjYTqYl9gXhk3Jzs4xWixI
bwSSKFO5a7Fd5JijQdlypkcBI+nH7kGyapJXCcJvWTZyzLvseMOXpfqQBvpaWUJJ
PlGa6awRDFnQVFXP5fI+a+rTggMNYm60lhRpt6yB6J9BWMzMjjomhoC0mXr4VxBJ
FXF+yE3L3N3iouEvbdb25v0LZSMXGCE5xRoQlOBGrsKotOTt6XUWIdR+P04wzxVs
c4D6Y2QPKtSGDUxmUTKRcsgwes10jpFDEYuGI+yTlsQnBJLE+hd2sc/Gfy7DTJ83
hRhk82D6omBoGs0s6wBC09cjH1oYhhTumqPQTGNVUXDHNHY5HahIvWHQeQi/Ds2L
QIcjJhBHuvu4nUbHu7inC1oEjoVvhlWg9a53FhonKPfM/JOLKUcmxXLRxxDVTMpK
d5XmGSz4d5bsigzzmPlWILba7YOebaAo0rCuPW3ipCIxiY4LjFirJWbQWjJRFQEn
MIdVoeiPKjndm489ulH9rpI5aSH04FggmoZKleBqYDK4pSOuw6yZR/Otm3jrCYhh
NMvbT0QYWMlFLjgm8cuR0UMm2DAXf3JLgeKrWgmHQmYfLyhl/Rb/WM5MnPCEM5P3
D/Z3G6a7F3AJOng2m4JBy0VQNU7bTdYOx07AduEYMbd63thLkK8hzX6ASZkNqJ2B
YderjiidEbg106XGVZ5FF+1+LNWqEnvXC9Q+QpIi5sTjl9xvGP55IqwiTIQWxwW5
B5+uQnsXXFxQWBNV3q7N8zolMuLFrLEffW7PztrQfKZIeyVj0wsLXl7ALMBmBEMO
0jDlKvamZi9WeQHjmW67Bgg9m2FzGpPxDLxOwvqsJqQ7BNHCxDF2ZGU7Jn/nPEni
Cmpc4rOrjTGqyYD44HeUqPIm/Vsk+QzsyHjqIyrOgnmXQ4oXDVaj/d5yswS33urp
yKXMHUV1AjPL8GOLTfIYRaE2047A3OfZWtF0CXOukHL+pktBtQ3M0ywBRcd67Rxw
/eOxD8z6E8pEH9trjE84sV9lx4X4RiOtAE8uiEQ/XSwyulGzFuL4MekT00ln5I3k
H37KPY++KpBYioOKbqwJqJeRs3lvQZhnvJ02oV22aRs7JUWbNNpxgbhPYohzF4Dc
4y2s68A8mUvZdZgp5uvaWyvE2mPk3gLIGmmrVX/QhX9Gna0GXuDeFxybhfnS8OBl
rB3uG8m4X0+6Qi8iQ1T3P/dI7/DECZir7yFZ3+x4ApYYfbZTGzippu6tl9Ap/02T
cTJnJObI0Ih+knDB+A2gQczw+hMZZejmTwg2hfn8auJ+DQmssmGWSOhZ21fIYipp
e193+1QGaUgrKcQ0yp4e3BuTr7XuLfj124lSZCK+mKABMsGoq7lmQIiYja2EFQQH
THOCGJrh1UrItQ66hmUdYrvWxxOp3puqqQJFaWmH8fmNL5rjdzbgczOXVl6E/0Dp
sAGsSmMAYQh3Ucgc9re/MI4dgzIH4JvrKXJBB65ZgN0r9AXV161ARN0jF1b+XMgW
8SPO1xsZap80JUGb3t8wB2TNVIa9Q6mJ8x8JfSQKPVexVRrkqL3CVO4SfOjCum8A
DN+teU4RXyeWVv2ivX/feErhH3VBpp7sL/ELf/4mZXsbUi2he/HRoHkKK2CRiCjx
iozpSRLreNos0bLSTvcJgLssQvvnhjq19Fbkpg8RZWuQBLdjoli2tQP4fYx8Ga4g
O+AI/wUn2Yed+GbLSv6SVyXjawmsilamm76ciO8M97ZuwhCl01OriWE0XUi3apH1
9fEwd8z+bPhg71QnJUvKA2+JIPzV3j/WQbEs5tYuR95AOjPeXlzdXF9BjUxfze3O
YgBaw7EVUa407W27A8NSdHHONqhn5dSORBtjGHhLY2q0QSPujdKhs8A4Qy/pIAy8
O/NnsUnpc9TvbcFm4fkIcGqzhaQL/bWMRHVBm9jk7OP6Ij9/ksHMrxydtBRZLPXW
fzfU8UMbbVSn2jne/hdnU8RA/I+Wk5qY/Ecjp+Ch1Lwc/N0zvmKgIeEr8rumSrom
aT1hqCfgMDJtbgDBirdEKyn+5a4H006TvziKlrm+iCrka7GKTSV4jz1+ejSwZhEe
I3ZTpRSO+1yknGWYr7HwcYv685rDLRv68lUYHRHF+qMz8zFnf4xTg9yaP7zfvIu5
o/MyZN4QSEUtWFaBuxIutOKw6vT+kb+cFieJUccaTX2QUrj8quUQsDPm1cfmKGvm
zQ5l2Pd6hXF/WhkeTxgn0mquZSGHS99eJOekrN/Fqa2iAv+g72hBfnFnd53ySRPu
SLlR7q6/w3CVd5cU0tbFDgkygSYyv1O3wMAvWyGOmuhozSYxkggI8DjvmRpe851/
SmEIuR0Jh/I18cFIcfuiSLb8/IVVdCzhQCadj96YpHdTSN8n/0cL8xBnD/Q25j4T
SfFYj2Lswxr87e5Qm2JhwpWQaNSw9lQhW7noJC8HL3U3Oamumei1ieBWkKrJZIHN
IpCpt6dn0E+HXHiHjHtFu4qsRcn/TvmfRj1bxwiQk5s9IL3USbGFiuKn5MGqllED
xtY0a9uIcSELB+QY7SzVNvBNpXsFr0tFgohyk0cuU9PU5tcZoNB4DCefKMgYXTKH
lL+y5n48BICUwYJNcfiDNCiHxdB3Qs387bhPPnH5kEUbYJiewoPPKNHlxI4hySyL
cRJHecfrA1S4Q7HCmOQBrgYUuO3Hrz1KtwMvFm+siwgcm7lX/x965pOyjaGrTorL
NtXPJXrCPqdiYkmlqLEXRp6n6bNcgqnI6HvChvXDCwfqQnJCf4Nnh+h5lB+No8hZ
sR+0IZbt+0q0TPEXoyN3LYP5UEKMHST6g0grmiSVihlj2eGny6nlU56k7RCvtywr
d55PtkAuzCkHSx7leYBaTpaA1nlV2T0XksNEz5MnaKHsAGcOUXlxl/FpnNzRnS9E
CUEa5fyHt6/eLG2f72n4PZNMUBE1gfxrXioXa2kdgbGPXTlGQqMqgAlb+LlAG95u
RmVjUPEJF4LfE58s+U+ZRL+egdRngjPfO6dFU2SW51MUE0AaJRczD+dqJl8syJLC
LWYWHk3lY5QD/on7Xr1+0gNmG0AhL4znn2F3e1OE9GPYVK3QjYfF80hDDeSRb9vk
t4Ky3uwzh5rZBfymFahTUZXmwPfv10/iGBvtJXZ+eB4XxVL9SPPBY83WOpkrrCK3
B+xOMSZJpYm2uMc77rVaT6V7FXTYpwQNCpxoLITqnjttE8nL/W3ClkKayDQYdQWN
5Gt82CJtF/6EmVTpAtLdbgT76Gj2KU12V6Z759OobesbDJCp89LkjW1idpRSCEtG
nWqGZ0/Dz77l+C25UlMzMVRJ7//QPY11efZrhBMKCvYeU2e51urs8I9b4rcu/qJm
7N4ACTvheCUqQ+WLHQAKVDJ6MwBsoC9bZOlNsK95OOlh+NoTu5zVhqgQZaWapOBZ
B8i3MJ9XwmKZCrzXoIQEuRweyG4gWYAjmBeykA7CrNPM1lnrdcPBIGiKXDYYQOka
/2lydJtWQKcpvcfbcLnypqSNBRnzDfNaOzpanfKS1xJxokbR+ZCDKkDHFRFW9pIl
3jjhz8Oa0vWlc7g2ALJ87xUhY7b/grRRa8OV0LsPHVTVxHd0DgDKHW2katN2rOn1
VLzsAeDpuXbZ/Q8uiACMrHz1kCUu0x7EoDTz7GdtfcGSKAzEOeWj4D53w50ZBu+/
HjOKb+KPW36mDoKJtRuvsplV8C2Lz/MlD4Zk1p6BM+0gOjWbcOO7FCpfpxnMphT1
14L+OHz+lfkm4Vriekibgfx1CoFRGzdYMtTeXJhiQIC5+tIPQWiwWk2sy781eo5v
GhIgVA2bwRuemorj7/Ozi1wS0/cZCyYAVn7skbBOIM0GyPpcIGjzQ2pBdcak1aIt
DjV+AcXzVkSE2Xs97L4rxkO/7COZh0pWqDcrx40jgPjFhL+Z1QWSfXfsOcoJpNUr
q3RIdsQfjqwLFlB/2VJV9Xwzd9tSW3Vk0YdFP6zdnitJ8zIlxinmpaSfzhka/njB
h/rVzReH+lAnUCpVYzNXLxWqiPzIlmBexWt9auRRf+stcNGpd607YRAsUCzI9kKa
ipIII/VyVoopajPWyMijTNdnb73+o9XAnVA7F5FeWgtzaGdV05y/5gCXymETZqYe
Peh2CbHwv0xGpqPdLPpAjVlw3Mzelr+dsYG0Wix8GlYVIwE4OfVsQyETH9gw2TBT
SqX0/6LRiujaHhpVzUAWW6ztx6HYIouvzUULU52btvdYwU/gkTYu0vWaIvPX8WzL
fCf4vTD+SexVHs59Wz/vW/pT33Nb/Ldd5j6WpP/CtNtLOCAp4dAYxU7zmIXS/2eR
7WLtPoghnc6+QMcyJhY+S6b3+XUUBY7N6rNuew6G8oZ1SINOIISaQ09insaRyPNa
IzeycvXWrfgPg23f9cNT6toq6aLARIC8F3JbIqc2YxDGVW4uPfJAYWraKFsrElx+
GK+mn+oQsi/aXuAJ8HFfnPS6la2jPxxM3a8fQwXpMXGQzyJnpvphifJPg3LA4qOJ
icBu3UZ8PeXettEWR138eN4G/Ap7R9fg7nBrUwpM4afuHvDWJn1IL+PPopYqF4Vj
ZGao8bSuym9TbimFWi1x97YwwzwKzVzRY5rkH7POk3AJDqmGxU/2c7mEW9oJBJ+W
9m7w12xDC3ezW3dz0fejmY/rz3hWvDpG+3voDd4RxeqgaRXwA6Gys7tfhoQ2ONXz
mu67jLQVM1U389tIkMuu/i5Oe/zZJhZeEecvZ2fUnIG8vlKHb42u/ysq+mRoHrfy
LlnRodl6539sv0MBS5EsdNdY2+gPpuOjqIaxtsgzai99MCJdYNtW2UXlkoUV9mDs
I617arg+L5t4OPhCWetEguT94AU6LH+YXe8iTd3ZJ0p/Gn7BrLqQitQK2FTZRfm0
7lLR9+DeYUA6soYe0/hHv6jMk2rXyHQQ5KCOv0MxopkKVe2Jl4FarnjuH3nW+JEr
MOqOv/WvaYgLrPHEkdrZTj5cverJooEIJYsGPiu4f2gYaTCVqYv8ZwOfXWG4f8Nc
eWSU0G1EK+t8Dev8r0MhiCtmtyFNEucGGNjj7BhFI6l5BW56QmtoOwRdvBSrQDsf
mz2ehfsvnKRPahh4kAGz8w4iOezMko+X0y2foebvkzuj37F+/e4MCmGyHrciEyLR
cBL9X2RVB+1RlcP6aHoG4VxOxR2fu7vQWczWyzN5g4RgtxMB7yCYT7hUXj3kWMQK
cCWe2huB/7fEQCy2ykcUAYpHUIh9rXQ+OX8IpSm7b4aIi/0PpHVO5LGYKt75p80T
cOiMgTNwxLNoe5RxBGyJ1e4Ii6IhWA6C4JjBnPduVsmvoh7L4ReF85pceIsgwhhq
ThqP7KMyV4Qssp26qmzd78i6isdusFjChlDrhcGjTORazZycqWhruLT9+JbPSfoK
7phsHBEPJ2oC/PV3V3d3yiavqnQIoDEQF0n1NKMn0LglL2xZxSFLlRiyz3CzuNUS
i53NqelOfI4Hdpj3yD94o7e+Nzjkvr4/CBRv3qqiSFuQFv0U1KHGaQVUh4dTHe2j
VXdPCJXm29I9kc70kiZdNfHoqjFm5wNfKWblFpQPHsYyx01kUq9VZTUOYofCNVoE
EwfBsb1XkNoQ5xMmPjVws+RYHQ/1f+8txpWwx7rZIBqkor9hV1qJdYTy7WIf2guV
9+QL6MiHEYnCItE3jX4TJjsTwxL0kyvHwsSGlmt8rgVdXj6InjUSU5Z5ZXbjAArn
LUACbV+s4nRc0Yy6aLMEPhwkiEwpchNn4D1ufw0tAUsT8e7Is+sGgxLt4/EvkLrs
TbBjqeEUVZ08Vsc3ClaPvY7/D6On7qh4lp1eP/CBH5y+RTHushkuXbXCyf7+sH9A
tH9Q7Jr7q955rsBkyMjy9UuOLogjFF6hnzzFgUwD9xX9I14a4kpcvyl0hZD9ATHA
XkhIQEpCbSALJS7j8u8M4za11fAAoFcxD+X7BxU+LfrsG/mtpTZ7m6xfo7RWCyJ1
JYu5Ifhhfj7DtwjzCgQsGkSX8DwU60cRKDbphIJBoVtOrohia4XGXnBHR6EdmT7M
FBHCSPodCm5WPObjtw/D9+7lpjD+cpDMPv4SoPD6wvpo1S8DnSyxTqr8AZ3KZwjk
D2s2hZXcrSEdkitZT99IxykA1AQzwjrCUF0Jsgo1MM0P05kRscya+nz72447oyjF
HthYvAWI5maYekPB7e81tJV/B4dykMR+0c/eBgxr96l62La3MOLrSc53HoO1HX3h
jaBIfwISZvte5s2bj+4rgS2NLYawEjMb2zCNVmR12FLs83TPvyMKa7BSGrUDI2J1
vbmxILiq0bR77Kk0oDn+BTlQFLHglXcIw/lxsHtN2pDmos/CtAPM3MGSqJpv2y8x
xJh9r7FG8LSLIvEkbAScgFOeHXiPL+GtnejY4mbu4K7cm8g4I0KuKp2mBYVw0pOD
Jy/7JQmpUQHbpwF+0sJUzHf1bmeZwvBw0ZzU4dUkwu+LsYBjvQaMHJy3IrsnZpne
HzWn63uI2qXvH0/9LTDB9+08CyccNS3UuQXjakPpyL30E7ARihr02WXL01pfiaMn
q2ZNzArm64fZdItJpLhy2EowpGuBv0DsyiRriKCdzV7PMufPUxXdZfGeKoq8a3Qc
0NAUiSd984vDtSA5IgiwonoqSEK6TSdoINFkMUWq4k+o6geg+2tWgr3kiflhhOxR
Bd0/kCVCHnej/egb8ePd47aIi34p4G8Wq0jGaOu0PEimaQhEkMiRQMvhgYheyAzz
2EEglgGpiX/AyRK9pwZdwwUYQ4RAcYBBDvyXdrSRn9IhWTG/pDQuLBaffGbOX5kc
Qvjkh1XNaIqJnvvidMw9tDLlH43CN0zS21qlYdJXLJW9oKtYXWLqyRZ8py9q0QV/
iqv7igiY9xsiapyau5qL9mBop2QURhuVJMVFEtgZR3pK7WXXw0ZFO9omgBaUyxtF
QYH1IqxHbMhvitT+RbGkG2Zn11YbaW6pP+oWYoI1+7J15sw0xJQk94AypKR/7ZQy
wmjqhOyG7vYanWhfsoi6JO2PA7Cxaui4KWm3QseIrW0w8iCtz7KsZBKYo0n8bK7k
W+4GqWt2wuWovrwf0iDnEzuh0vBrPpDiMmzWK1oFciilOL/4N/D6c8IZZCnPfsxL
V3GLo1QZVK+OKxgG5UMo1KZrNf5nyYlfv5cLmIO+39aeHLChomZFuFdgtVANup76
/jBrFCbYRI+lKJVIS/8Tor+4j8Yygr7t98hXk20etu5vvAmwFl3teZrF1NY+UUDh
J3Vvbi/efVwGxlNKIhFD3cYigpUYwHj+XYleMs9Mftt0G0ekjsJ22YBjIVT7huXs
gR6TFMQDQ4ju580m0PffK2Eh9EbSr3GFZts60ujzamtXUK3vKmLHYB/8ZJorMBfn
WFtCNBSJfZFOr1pQy1g1Qi/a72aMZTYq4xRCEWs9CncB52v+5A17sopblYRHTz4c
62BtaXO5vPY+LXVDRt0K9+xjTQyEIOwe2R4XyZeKn2WkKy31vmHAryWA8PldNEJP
pVQh0jQ4bwJifELDVz4LqOPM0//F+N9s9FFqsNvBQz6rYxRLsvR6aKo1wdtzXIvP
dO5IszvXXM0yhFSPLQNeO5UDLMtPaZrQAXR0FSxJQMyzb713phbVgyDtoGZBGAmk
03rBT92IWnKUHx2bV8Q/ugqokQxfb+B3iERYerEhbj+johrRVzh1eqj/wmeqZ28L
pIAwzUmRqiguQ2aSuCi8ZvnaVLfYUy9yjH6E5bLZqqgXGJbC7uo/q/oW6/zWRibU
lUZaJYv5hb5kdLVCVjBrULNLN/FkmJwsRTsEDybrRt0+4oQvnpzGTbMFuZYh+BEz
6TvW/iY78b4IrnPKDv07OXDNj1NCas0vAt1dKS6iIaK/YtDjjsvBkeK5BdlW6FQV
J+sG1gPLW7g9DMFZQ2m+bx7zQMcyw5qoDZdxXxZ1Ye9ayC4iAXhsT07jdzM7PJkh
KL0qktRUj2NRX3GsRWoOoWN0Y2lGZQFhV7SkPAy2p0z3EmPoZYp9mha8e9HBe6+9
Zp8Tt1aqgF5gzkCeXhBxZcvKDW9JaRComSNpZ6eWmtpK/X4nsvNc7qMCMtIPyuo9
GE2ODWktK3z6md0I+JDrM6CMMpqaZLyPG/pzlnv4sD4dt0RSHaZa2K9DIA3LLyFe
kzgNybbW69+fCrcT/NdfI/zvLD+OjrowRvLWNb8s39LlffFLHgRvh2Z+2r5v+6x8
ct/yV0rQYVEvFJELXZ6vue7QwmDvbKJbh4TaHVh+tBOnHvZtNOBVNCNVcfwo+mtb
O41COSqRvoWbLkSV5najxOMisrxancv5Z9UQvb2WigzBnTKfCRro7OmmgNkCGg2K
nWMcPH1aSmOVaFxEmWayF0um66DfYXkc3+5zjchIdzZ7OjKJOW9ekbI+zLrnf/Y1
MgTDG/2TaYeL8aUF1NXwgSVFww0vqjPGtUDSbDfUVLKrJVNaBaNPEwVQfpWK6+aH
ZNwjL+RWE07dok1dbPP9It99Xyyh8/vT49fGzzIDDOEPsvhoSYDKEZXW3Q7QVReo
KJr7AITRuXXBhfxlRZkoN6jWzl4TH55myf8kkvmDCqAP3/UhDySnk8n72PbRy5/6
C9vdSa4/hIKlVZgZqkoQkeILtLynvVQJ9ONUt7c/uzZiSLYvq1DS6RqXE7CLc5tN
ggJpYdSfSIzlvlFdM8GPYjk/tYd8mLZf9iXTlK9zhZwgCxypGK4IAObVgMk+I4a0
JKtNEBHazL4sWPWryuX7rSAKOqV60wgweTXi5WqyxMmbXSfDMo5zOwmbbgIN6ZiC
cxSlsiXTjc/MJH+2kswXtQvCJvOeedtXuwTK9vDQ64SAFv1BZhqwzwW1bzIrIzL2
gqz5IUDLmZgj36PayoL8Vm59vd0Btjjxi1w9t2A9x9s2tFfGAEhz7kmrmSmqD/R/
NDn7jcn1NMLgPCenXdBIIr9VbtN9HYru5LbSa0iLryt/HjlInWsWiElINVGAdUll
SUYBNBuHhrByZw/pKG5hhFhzUcWm2UmqmY/Vo8ciGCS1AYOqLl/dzrkrAzDBuC9R
vSfyqKlvV2tuvlUW63yllXtGUSrEeqdVKSO74KO8R6MBlJuTceUa+x6gWnD3n04N
/+4EiVvl3zFxoqxfkSUgym8oTofZB+RPPTU6W4xZ3HU9hoU5OD/nWa3yzhZiQbAD
lw9gr90a1V4MxELcwnANLMxq3hnXCW+W/+Cq6fctn+OysYawEqsjE3CarPPmadrd
Wg/Ou8tCX06j8UIGrlHWYyNx16Ap0968Babe5EYYXf5IR2EiPSNZlv01lqtsexdr
ElgkebLxPSahxxpopudfWxuZ4uxp5PacOA3xUAlaRmO8OGIjCAPKvLGtgWB4uP69
LJE2AT9ozPlUGqEr+PWz1y3EKI9Kcs5OqgAPg4jQj1iht81qIN/VI/vlybAXTTel
LEqljbMBWkMf75tA1e2Yudu06zi2Gjk1WiMfxpUJz8WcSA0ew6RzzwvuamqMxT6E
Aceky+kYRYO/xTCprSvoUOEBK1FKm0dsCo9BRRbbp8f6Ry4nQFtqoZXqbwoJqMUB
Gw2ji0xmgc202px5U/O0CYK99tU+LmWFMLzTOO9JDnJS0DKDfF110p37fxuM6BSF
+FMx05qqMbqYYp1GOzzsh+KCeG3dl0FyyaADOFL1P0YzGFMq3crCwgHSIUFgyTM0
u6U58/0fq+Tadj8hl7V982xheeRvL6ns9Qmab2cKKMohOpRzJ7iz2HQ+jL/7DROs
IaD0qCPODvFf80p1qGq+eUuSQsiD5jjeJhMsaNFNnLdqKBrp470LKKpaLz9S3rjE
BNjqh+ne/GcVa21/hpiapoMBn1kD4Enu0r4uWCeb12gkndGu5DugMXZ7LCDEA4et
dRMWHTqDZJJBk4K+XnyOQ6Zl4gTF7Oc3X9FjUALTtl49A+XaGEuLrvN+MR6mgo+t
0mme+r5GgPjPvO4gqf/dgK3+jZ3zYjLfEJprRGmJHmLlK24OAVt0LVY0xgyp36yR
1aj9Cv1EEcgwSK/1zY59kWBGT1iX+srAjejzkzxbMBCKhimQjTpBvGmRc1zs5vJs
+h7WQAOgyKQyL3SaTplA3DdT4Q8U8gDask8oZkVjOSYMWWf/cUIWFAdufCvVtalC
20d+QUWdcxLTeImpRzq3Y/NkeIzhd6hGWl2XXRAdwYRJVYF6GLRqGUewDaZJZ+Xg
oYw6DUXJqxon5Rsb6Ki6SZfvqTTWh/x4gcYRUhRl4BNtWkLJpKYBOE+j0BRMaNw/
mvIhuHUkl+KRkKrl70nMkvrwtoUxwAYSHWZc0YY1AZAKOnNLfuHZ3tgcG3gkymrf
miTaqVKeRcyG6aMkMvetHocN/g8n65ynm2PJCfYcQkugnEB86GWxDuWFos2XZH4F
rVwp6SqrxmEY0Y24HAB73/XI6XUSoR+VDF8aQDyZzMfs+cHRbgs/+BTQnRuz0PA6
y3wDaC972jTNZmiCqGGvMnT4kP7Uzvrr3LIEekhH8NEmO8a4bp1IsiNt4qAUTihC
Iip8n1XRv7Lyv/ikewaOr/CrXF6d1EVDBE4+JKXzpAtgjvDbcS4H7avUeoLjzZxz
wqtfvoEs9Zp3rKG/hY91QLZhIP3QaoqlxyaBvm8WIUQVgmBYFklHFSSCu7y4p4uU
lNB6UDqIwhquaSChJTTvOC/1kxIz8rLAAKoDPsBSgzXxjWDVZ1WmybOXzmQ94ffK
OHTVllsrjvnS34nJOrvpeKYmYshKi+WUq6setxN7zVnXa73XNeuZn0h9cI3JDLMX
CB0crSFBnEJGmAQXTTF3aPbhlon9yeWdsCeN7Td1vpweEC9SQ0uT4JPNr0mg2YOZ
XB/wqRv+a7DuUPDkB/b/TssmogFNyuPs642LfjBwyRJYrO18bnu6sR8wCquX7iAf
Qsox4HPAtd8JPqqGypAY+Y4a7FNt5TvS/VVFoc2YScHJuQNP+AawwjEdxBlaeQz0
cIvFeXvj/XQRagMOlcrcTA==
`protect end_protected