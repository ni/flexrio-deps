`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 50560 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
lmOQgIOM5jiJrGbWpsW/8m6AI0QamD6tHhrixTgFXzdqVckbYoid2UcGpEmuL2kl
vu5boyY0/2xKM4IdoecrpUNlRAKxI4ys0z6wrU33o025gnWtxoT2300pN0LOZs51
+znxeQBN1iiccitPD3mVkTob5fpKN6/RvVjSqK3cPo7Lnog6L18SBaDgk21SJp0x
9mJ3YkC0MkI4L8EQNdkRg+M7cw6oHJI0Xmzgehkbq/rM8C37nN4zjeEPBNWN88WJ
mJ66hrWW/HSyvdveV24pc4QN+M1cR17Z29dZCTpvcIEdNj6CO6V4DqgrMcFBGxCo
EW9iCrQngtuJP1VZoEC8xs7Hjq0Zu9rJv7r8TzeF7/hfmysTo4K3uuA6WKCfBQQd
AedQMt0CJ0GOuDivdm5vq+CMFW2vVM2oM5/3puoo/8UV4qRw6KrWE9gMsCL8wYmB
OtoKC2Jl+0ha+703p/ply71Mr0qN+EvuW3r1hqcnIVFzmfsC+46qv0vRKm6xs9is
xjgCT7UBbJnR+5vdvfRkys0ELlKWrS4fw8BXLV465U1CXX6Kan/IlVULZnfRk81I
vYt7qJgBRGbQiE7FfzMIl3evlxvZbDC6YUDCLdCyDPA/ohJF/BYdxeGf4HGVNJ0g
09xPwQ+OepEeyyESZP9Yw5kIbN03qzD19qziC1TIReLfOYE1owVlg6tS2b561BRZ
9AQrcUXWWe/wkhuH+Fw6ukYX16H81IkhngQeWKA8unDHx+5Of7hvWlJ/XCX06Xwk
LsdtQQR9lo0JlHp2s/M120XMCLUXR52vuX87iNyOcZ6G0BCKc/jhNeTuR9DC2tQl
JJzaytxCIIMnPN7wf0PmQHtg2K3Da29sNF2k+NqltFQ4d0v72rHtBACUaHvVeTz8
LIOzWkM5+Qj1dCbX7l5wZNI0CQrzLpgmLkuU5wNT6Szko0dj+BefX0uGapOwBg2X
ijQZcAdpw2IKMH/+DjKeES0d16IH0+R1UKXHyM/P4Rb485DHJreGj40GRJy1MgON
JveaNKmU4WbbaqbP2PJLhVcM2iboBo3BAoB59RQ00Fgy/0/WQkXjm7R/rfWmEnYA
zJYMOsyPYsleqHBVfY+qiMudojr0q077od/pJA/pKHEfWzvsTpySNf5Kii1Cqle9
cOnPHwFCUybC4NyZsKJRjUH310jWiednastNAh0oQQBHDJEscXB3E+/d3ojyKRut
VOyuCUaQwnzvFUGixP2B1R2qpzRHHZuAvgAxRieMfV0KX4NXR2rLOCIP09IplU0U
U2Cx0lsoWPhlW3SRbhmIBRsAHADcj1tXDxZ16Zy9coj0ehxQzCx+lrWL2MTY4PIc
7rdJlUblGJ/BZBuneg2srK5ezqCinOlEOo3wr6cm4vMeBbM2ekmIzBEJ/Rrke9Az
19v62tZ1Ehu6WhAPQUKEsAROSfB0au8ObMAKxIOoS2DL9mbVGEbQdoheJhzD2zj5
2T66uEk4PNeByQwS3auq/jbxCCJ7tvb54X420NVS5jaKVXhagNt0JJBp9qA7PakU
hFGt8zYW8pYIuB9bke3EJ9IvLUOq/5QF2AHtJAdp18FHgqFpPBsVj01FG+9+6rmI
mD+4hvJRiJ0De4L64zVC4yrhpE90djY8FmWWje+aE/eWRHGwXYRIH5rKDRPMHXKj
kB4pV7lNLHu7Q2r5t0P4RQsnO4NxGYkH0Of0DGsCiRBJlrZHpW31L47zh0muwBO6
ITWGURv8gm4OkA/gQORMlAG2DbcxJlVK5PWcrV9ZiZg+d/OTXdQzwC2dmpDVgVSO
cLIluXX2sljbDP3oNi1a6klss0yjqorxRCwi5j8BfJqobGZ0evoAsY+CUUkABbM8
fvxMc2LxiidMfwGKwhgMOc6FiddaVI39KgdA1SlTfbeb3CbtiGLnM/RrBRZgM+vQ
/TzE3n0ICrrY6G8i9TSCrAApklTEV9iOA1NvLzi0lyI91WLbLq/tp01vxCszHozd
EvIDQSZx87l0czWX83ozc+LeLpknI2Myjkgvi7GNkJEDtfTtD1Hs8w4+pU/FFz1E
aRfH2v3RuBugyH0APYbRLfFzTNX74aRerJBPF2R5yAFRpVxqLMejLpCtiRgOpZA9
xA3SCnMiXloTq8YEbfJ0aToJvFDXfyiwzc89r03AMzCOJjf40HfIiu1xp+571c05
tuTTAPkDe8FkX52VfNuM9JVGNfIlo75vwvZfGoV71DakoiD2nIHgyUQD6UzbQ3e3
YTVFGfSBsqvm1Q4vneruQUxUkxScRPZwhAGANkbmWtWfsoW/8QaXP8ZtUB/r85n7
mdwItCFJeYZ9V4i9IWchKQW2W7z1RT0GgySThrM18fxAwM4WUFZPmYra0JC0YZDz
6371uI4hgyP48iR6xyMFSA3C/63LI2lGoW0jXTF42gmmRAoYiOLEpJsmC++Zn9pL
/0+5K8GTY4HVbLp8PpPjMK4Z9X6NDFJuKH1iCKfdtMSvzIK8o08Li5w7fHMAshbB
Noso1YmM6X8cKb8GfL9rCbL1PnJi2sxMdyrQXECd/JyKIV+KsLYSws6kHtCZp3it
nH/ynOT23lYmXALxPEtE+BpS1A9WOYkxBEVory2U5NAfLwCZ6mpsPp1T8QZijeIy
JY2PMhuo+q1XPrgFHaRelxEc1wT/zWZHIQMMG2bpVo4F1fohhRy4tBatBjsyONTY
LaAmg3cBhqAEqbL8BFCWMEkc5d1FI2Wt02jpXZatweh/5LCdLbkkoib4p7B5W46v
eXYINRvxY81ck5nlbV2QCAGiLqw/UOGWz+yDbOdw4TOl0RgJvWIJvpPCFAh/0chq
rurKhePBZP53YBMGGeqedEEniFTEftBHszQKGs4In5pUqubVy0gbDzu7XuH5enCG
97RAs04WZLGbfW0q1Qaw3gzLBjRhhsjF6ZND7JwxNwL/tRx8vow/hrl/BG5tej+V
8dzwgQLQVCu1du5jXG5WinuQyrI+ECiY4SrQx4rZfsNOm58pq882kYbQBP/CHScH
r3XlAQmpl/qU9xUk0EoAaeag158uxH1CRvnQEexpJ3Z0zuNOiGd0+Z1MFzGjt+4i
xiM2L1MvLmmeoXW/TkEQdyotn/7i4wQjyBf5pbetPF0+SolG877UGMqbV74QCrtj
Q221mmR8KdmHBfX9B3dkqnux+BcacK9BY2aezbSPoRLUNoIMky2p7tnte11rPdll
12WltFC+OCsw5L5TiTPuQo62Z5EkVVYDA9hrcD24DWzlyrqwF7gR0UgakCTW4wPO
imOpc9CbGa9ZS0xpUB/BRfpqMJc6uvIzPJoI5xjgmmEu/T2hy7b3wlp+GcT+TOpj
TPiTaFBlYXW+qKPuMTBcDeYTarVQHWxaQmvZJP4A6UFKDVn7sXDY2FjogCL8HdKs
VDpzqYC/LH4JYWYny8rl8wnnT/9xzZVnaEp+U3grc5WLz0cnvph94DONkw9O/hpS
nY6zE1xA6xSyoxmg6DpC7k4PctCSz+nXEd+8XlCuYJTiFPY8e0k7k3lM/LoUW5iH
rCRVUtKuZ5TP7vvwiqNNnLky7WBaCZ6nzazf7cZT8o43Q5DM7I/AWIcfYxk0dz56
qbEcUVtgcm/3enHvc7p8t3uFlTUCR76oLbqs+YC6vCaAJOBhZdd0Wz6Xiqsz1tMm
+UrtzKnial5W5aGern0C31TYj65oHfSr8TYhDb8eB2jDrhfRAf2nZENY/lqWXquO
1Tcc9Q2/3nZUsOSvfUgdz1jVFWC9BmSRDx6rM7uYBHwemOqOwb3QYGsqiP3ujnUp
uPXupr0cyWRHAbiyces1TcTcXtgZkK9fXeVuVKraNEFxYzVgct5oYIYdoI3X+fsu
0OLjrOCJaFiL4HJF36Af49UTIJKYS3lTVTUFDKpCAlkwn5cpfo8kKYp2ckhVM76l
W7aMsjgWUqSyCDoEoQwRYDqF+RjZov8Tnoa/myRufOJD2WLJ6cEXMfeRNTS+24dJ
0nAaIJoP+RTDg0+f850ktj8BSRes3wv+THewEN43ts4Lie7tjjw7w8fEuwt+aRtc
zPqqb3r4nfKgg18MGLIX9J6lqpKW0fC4e//PfoyDCEA2nDHU3k54BDl2Is+Ouoql
xgH9R4j1L18AYcTFIH21qBfu9EI1UTQaqrYmyJfgkeeFnycTFEfia16rVer1E8Me
4negx4WlH7t9VV4LypIZ8q1AtE2iQe5xDlMjl/qjvqVxO/hE2YxUtyp1uICb5Lw9
ymFITBqMdxrr2fQXLSOvcAwW8Zyin8+U+s3RG1FoD7XDFKmHpvDGQASjimAVPP74
iAF09Csa8MHTEGtHuKNDH4tERB9v+IEmK08BhVD7SVBi3BAS3lOdmA82WjLDZaJh
hp+xsF9OvdDDcz7VIkkyKA3Hyd4Nhb1SoxmLlzPp42nFqtEjcTEx9puZWGE2iU+9
XniZGO5du536RgB6Zah2ooX/EpFY0RQBmuKBJNrnbeFPK7RAqDE/RC5KX2opozCM
rcx6UhZnAyIzOHK3fMtlvWowx0zCvqOIt6SwgkHlUY3/f6H1cZsoaVf2MxDJC7/w
SeLAs/yd1gucUqogPNmBXUcc6VNeiYkNHW0kDpNj5aPjQfcg9kd2cui6fW3Jwu5+
yGb/QZaAlpmnyntE86MUQfwarqfdxIEZ1RjWqbqzdPEJCXfvE9CyqrVt5jZhLUN/
JeliFfphGc1fvvAfYNnQIIbKAOOXzrccAvcvSNFo7TiQSyIK95Z+4QC9UAgPUm0y
bouCg5DBQ8FQgpAklSo8a8bpBAnuAnvTR1DAM96qqtRmHADdeXtW14m7C6d7p6pO
mpkqE0Jn+yydmTSWy0kasF+B4bhQrzuH2lVwgjTpf+LFQLku6buu9n9xm55tNzP+
MtPuVfQa1odU4VnRa46Ye8FDG5anEi8vU7yu8xEwHz51lIkIAWZG/AEUJscdJmU8
miVHNFT8nTBZ29SlEHyZJerxy1ywHWONgqKijTqN2GGaSH8IM78ssck5GyFq29Oo
c4l6frHAnpxcovn3ru9yEnbZNwYvLG4bBRsEqjAejTAeZYKOE683o019pEkh+R2x
BtzQFNzheDS1R+cgPtGAQNmtiCX/HRL7bn/jcow3QiyfQPBLGadQHLKQS9F8Up9N
ubwUZrYShIJ0kbckMOy+F3nLaRfCkaI/8Hopb7m9/vSZRjVVt37F1UDRm+TXigPZ
t7o/Mw3bDoN2pfBLgvhGbsaV9IN+GQdP5yW1DfUmQPjMGwc8p2FV6XtI2jMflt33
fFkZCKJtF9laxPnW2lQNDb86Bdvxzfkrdzc/ehvLrlcVJ9OfvJiKm7KIYMaMl6m5
kYT8UV2R6eG8SUxeQfqd1m5wYxnD5nzjfRmuG4BfmAJJGiiyNxYSy6gLhFYuHuGw
m7KDpZqTAXBXeggmLWShFYFXuAOfvdZGdiUPY03qk3U9ET7GmcMmbtNJtI2HLrqe
eTjzcJtUHF0uRSKyNnlGtq1/r7Ga5B328Yt2wMYATjYJ9GPsAldtnS9N9pIAV1HH
qd1cR1FL01DPtJSj59XaP6mm3vkbcOlc74KltntVL6MbNk4G4DEUKRZvjGuYGRzS
fzImDnq4oqh4ZYpWWaOfI5fqkqSriBRTP5rrq3yQxcZI0J3Pp0nDn+tgs/5tNWCd
5yhkfQo4vUIaSTS08PKuy1SRLsOsHM643CUeOOMd/xqOedqeqQSle3qC4dPWBXKa
RNCeUngSQjPhMAWi4+p/OgsXVEWB74D/G2JNR/GeFxocg6exH5Zd0INqEv23UW2w
Mo6YU45Atbh/VL7JZMpyuNrWUTEwMZsDqRYssjcwSHOmvABem5maUERSi0pYal0s
p6ypz2HA6/w47NFdUN6r29tnXefJakfCPCIkReHkIVBCwDQUt+NyS4oNrdnJWVA0
uWSFLVtyP3f/bd5YrPxTbtuf+NjoL4gLfnadFSKlaAnjbNmrgekfnLPJscGv3P6z
m9AHjOi9KZSJYLBRCeyBk2KpG1SsOreVkqoCJzvxToDEfYqenE9wzzLjls7uVb17
5W8w/yqATI6Sy90zbVR0ZkYM/C3ZZZ1HCwxTkMUHh0vqnkkB6fALfaADx/hLPkuR
Jub3cIH6Ou+y2X0fJRVuPeKxf+rLXs11+v/W5MgtVONK0K1WYhPKmN8g7RrzpSAl
2c4OEAicCc7RN37e7PsEXoXJSB8dAU1Drkcu9IpK85oh4nkVEV6DXY0S80pvIpYV
fp+m7hxCPwHW9VNbQh3h3AjbGQZcc++7O4cR4XMrz+69LWAujU7bXOYIAteK3MFs
r2mYiI81KpEWTC6Ste1DJh6159rn/IaWBy1vAh41UAhauApSKPRlrgouJODYHQ63
CVwZBD4kbwh15hwOGwzZcUcsHYlq6tvD1FBcreTprjiIa6AaZ3uy235Z3zUjW7NG
c36B8wAcZ9KzwLUOb5obiwBfIaUoKtTfI+dP3i1ryYVWTEHHlN5eacEv0fV7cchw
7oMhdS4s+sdOTYO2BtY9ud/odO/2h9fbzODLqhoWJ+ITl2W0zDx9vktYKdSuz5Wu
rw5Xhldy1QD+CktwCXarQpxU7+Bc0hpiKuq94qqf8QLQtzty7rwJ5Z33AF8kAWI2
Pt1Jt/hlGAqVnpiGv63Yxrw1/2Zx2yCbYzeFCVzf8jG0G6tC4yeURUOkDPHKQ6qa
7FCkZ3BLuoZpIa29skiJ2yAiHYOtQHL72BTiylbA7y4/jPRhnd9K3D/V69bcek9U
bPChu56+I8EFkrw8epPxo3Sk/q94nKkMIiaKxebqcAesRKjipM/KU5NyAXcuwOVJ
sAba1Rx+vUA4UiJ4wEhLrk/wJhUWAg4H1LR2yzaBqdyp4zGur5/+9ETTdwGnX0s5
wpT/64i8UQxaNvE/udQDU6yPiGTAVG/zgg0623osWPxg8Jnu76Rq29Di6lBB+Z5p
uR606XDf6Q4Xzkdt1zr2B7+6Mu0P0uBY6EznzUwDFPhH1pmeifKwqoykwRL9aDzQ
1Seh3sCDFT4vGCPlBUSpN6QW2WZdv7PKumDPlVlyGgKqYrIoJFXMEpnSTdlsfm0F
iC9MJpUoTsswlA9TiLVIYJd/8njVfsDELJID17U8Hgc+mLZ4kC2ILKjbA2tyuSsM
pIRyX4dIJpJVB1zsIEf6TAejLbWOU2vbAM+Im0ZgJtI2GWFGs/v0iSHFz9xKVuka
VQoX2y4ykTEYX1faSoD2bb626dgTDsu8LALBHwdWnlZfP4l7K1WBL/qLTw5+80QM
9LPl8zhUdNiBulW4+7FDuYVjRBBi2I/A+xpMWA4/AZUCMvmruJyoeDpWa9Da9LRr
XF/M1eTbXTt3fjoTaPbmUdwNlQTg9rVVBzHGALDqb6XYQIO7sgYdA5aAQXQTmoDu
XRFml6YHnbgGx5VVETXWUgBDYqv2bNmU2UqyGTSdfgz0LthxhFRdHvxBF5bsJdne
Qz+6T/39wkKXUuteR7lQ/2qt5p5zXjLEAc+ubrP7G8JyJswn7Wmdx7O6erNN1Ti9
sH/XuX8KC2CNPSg98xqlpxD+ZjmoZsORiuSVVSL0qmXREcACuWCBHBM4RN/LUxtL
uBmJeU+Qi/Gub7lMqnTZFl5GFxcRBAriaBHQDoqqzhr3D3yzvwmWviT4bykBgnc6
Q4yW7Cfis5eQZ926MnW6ISJ8LHgqFiYFYhYr+YQjtriHnF4x7jq+t8EqeZ3Y/Qj/
zbvUpn+brZ4Yag3j9PowTTs+oY5a7eeUZjtS0ZRkpnzRKPqq8YXjAs90jhUzfKq2
Ef3csskh6hvPOsny12qXBn5gS/L5lHkQtVtXv/FwrJNV3IEb2+eZlNcyQ/ZjIEMc
3q44V0E3yxaUYFpBNyhHBPB3OuP0fr8DS6tWqejpGadUzj3PYeHH3gkMgDWHlCXG
BQwUQL2j6t96WCbd16mUjZebDYqBQrOY51V5+ozKKW6XXo2fkcwrxEMJeisvd/mp
8TD6FJVogsyN81PM92OuDx0a7ruq1am95m96P/sBVU3IS7SEnALYy+DxoMtt7Gfx
KLe5yYITjjN75VggD/Sw7LYCK37yYZxNYtkmUrvzPUvYFV+MdF48+qwwlrH+Kncy
F7NbWpHyVzvJWYRNCyDx7I/mjoK/WGQBAiWGX6RXGmo+plqCJbp94gZG93cmlmLK
YrEKjOEwKq1goyVWXEtq5ImwycwbUWSUGQcygRIdgKe68dn7COJ1FHJTuL1FFC3P
nDCp7/oI7piSz3g09HEUvW2vPceEC7dhWuBHokeoBy3jmLv4tGi+5Nan7vmn3oiM
SM5UV2LzKIMRcRPDZApFLEqGyYaFz8e5bJKBnBodUigzHcKVizivXnyo5530pTfJ
Vc/PO1Oj81Kh0E+907aZU9Bce7nYBM1ZF4LuiPutKMyTyg9VbaHmbK3yfQE5Bkgq
M0qZMpaOBYxabu3sYKR1Jm+KWE8HcU26R4buheAmqMVFTgdtF2XihdRfX2NLFmfD
9CpR1wUdLjpgTy7FH0RlRE2Bq9xdei1t37GPNTh1woKZe1XNZsygvDLwrdOiOhtW
QXUiJctP3x6ekKcToxE7SC/Kcp/3pFb15M4lP4Nlx2TD2Bckpj+bB1X3joezE0pg
KV0+NIpp2jSBeEefNwNakei4vl5r97lTY3gEtWaNRUOGDpP1+ALWGoOUwDBVkgQD
WUkLEoNCRZJOVi/idN4xjHRLbOxm+fGQspyfbR+7OnDFAuxwyFFbAfDPywaE2t9k
bAMSsOc9L74ONLtM6aLVrXp7BzZ5iXNs3TbZoxKJMHKkoQbT9ulcUSzwGe41rvOw
GH9ROKV0gQRItS6wqNtoyEibdUjeDxeJA4a9pCpBzulRknDZTgEu/7vgt9OMGCbO
t4ctRp3Ur9oOoQolHz3H2sr/ugZiqDZruPRVpTL0kjrd9WP7+FxDMXGwsMqIDRB3
0+fYGUuPqsV4whD71yCPxRSYIBhbBaTKNbNC36cmlwDL3hhggquwDAq27TobiI5Q
IqFOittTVUwA9YA04Gvkoe3Rghi0Y5/mnFpXa/i7uhUsgzfTbaWX2O1FkfSM9LeT
+0FRARWvyiyWSp5BaixaXkExzXEHj+pEhNe/QrU3rVD/Bn2GcLarzjr7k5s4+pXd
qGsHs496pAicrUZ+jS1wa3gOEF0IgsN36N6nqDoffXPQlqhLst06Co3IYgoVTIwB
orXE8WwopB9DZtr0jR1V0WxsVhuxAo+ea7V1XZZntbIpyRUUiht/yLRcsdHewyRP
Yn0T3s+mRIf67+4qbeoOZBGY6SXAggI1DGVgPaKmAUQ1A1EFar8ZcJXsdQuhgd7+
bETboVLyYdsuFv3hk2ydKsHly9inP6YzL56cz6JdeF1hnoiXu5iTeT8KrEU9dUKd
Bj6pAYOCWtPSaJ5wKetoF8uqoYzz/pue79rM3PTjHQ9oxGtPGrUpZtbDrxYwim6C
f89Cp6lGtiS2QdeOEveR8hEwASuVQbpVlt4j8wFgxvBTO0sytlzvob0dwxjBi928
D7mFTIDATqh4ansFum2eQD9K7kgibklN6pziThLyHjc5OgD2uHZylfxcw4xtbDBt
sHudL8xANlhQGjU5kOU97H3HB0E5q4OYfe2bdUz5cfMtR6TwTDKz9+zACfnNl7Zn
5RaNreXVy+Q68GIl2y/8Atu6j1vulR7a+KkJ/lBAwRbWvlKK2b8xVrrd8mdOpzxs
+o/HykAC6obP9Pj8+Jb8A6LhXOAzeQ0q+KWgdiW/DSD6/Pf/fXd7xI0Fn7cYyQmN
WEpPf7HaWlSIBCsWN0crCDNvnnt1bC7+IZkiI4HKvRalUkjXksikpqWkqRepLc7U
KIiJt6+DgrHvDfTO/HpttEO5VBV/w5ZZHE3elV1phkpnLJFBi8XdlFnjsL2xoGvi
fzZYSU9WzqjIb0l2ovByuu8JGzRyrH0slfXuIvOKTqcsoGa+LIMAReEKBiEvDrXc
NyfLUTDLI1TVTjl9RZWgPkXHG6NwmgqAhTqLSdaLcmy3ontUx+PfCfJnIYtcHgLZ
yEklyq8retBxW1tLUNnPFa6tac8CCBfQRp3QsBV0StPNKzWM5D+7DjnYzt62uV+2
3LLDk8JJPj3vdWZWtr4VJQezdodKzrHmroNB8HCJz/T+UVRbeIXbopdDO3w3W9BN
6jr10/ZKa3kIS3jXfJ9UaA58uxNB32olyl+8/X/Ls/BmIdWukjlMQu0POeRg4y1A
f+6LWQblSI1/9Fm4LRiukf3lTLZjC2X+R5ks6ewb3p3GajeFX6RXtj/S0qqa2WMY
PPD6NaT6HSrGUNmzgU7EuxeRoEVXcICg0rbwpJNCJCkFQFsfEm0YFAIIEt6+8nUT
hxwUVZz3TtZfX1QmJQu4ebhkaV5WD/fAqMj/yWoOlxkfDeJf119uhLd+81bvJFdb
E8v1NkX9clPUG+0briw7NpAKuGmPYwpNaktw1xnRYf/mtpQO7Qvmu9Ewuu7Qnsjv
32aNGTdIFFuu1Ha8pLjha7eUoOtyn57mELOxPSwwnJR9I5nvhv7/bikb+PXtdOLE
GrChZwhLTTDy9Ulz4sPoETH2LDaU6fOx4oHbhVu+frxYe54/nGhs8xP16xgAS3Yf
1qNSdjLx7jW64gjbVCEth/KAdSQMUCIJ7+QD0hWvrieoiOx2BtDlMXFXE6QZXA2C
PQFVRFPcCS+rmM56i5AGGcoGelzNWJ3wDGO0jtaijwDjDbjNlH+7dRlNdrU9O51t
vgSlpzZYgLjJI8bLlvUpJHTsb91BwQmQcTFT/cEk6ym6v3yK/WgfRkwcqjlAj+LF
IrFwmp1c4mop48nb2PDOHyMHywRtJKUxtquH77U5GxmHi2OXbFsP2gWEFdcYFsW4
obUwXeSkLbko7+5ZCTET0j/qvzTfPB6Vs7JAGNRiDSou8b1BA24aOZj0qdpoPdX1
8a1iIrpjgbt3U2m1pz+2tZfYvdQJwb6+jbzDOvTI+yIgUExCe+D1OYqOi2AlLxH9
kJ7csb95+QdAmANnnx2iXKIqfHwQauBWCwPsuQZJU8ZEsotS7VM6nTb73dDiVsap
vq9VRygCmV7/tyVow/F3kcob0Q8Ujdv0QRQV3vYeZsB9Kv3uPUWot0U0owQ8S7Uw
kLd3qdcxooJFCT9aOQdSOIUFOvjtTLPQvRrpgoSOoxjNYrEqoNK4dCRzQSbCE5Ni
iS0yh3KBepo7FJXItHac6YDYYtmcfp5AAIvjdQxmNWuLKMRL6BymPLm9jr9bN0vw
aSi/VbD6LAN0lKCrIIykrgIcCnkW3y8g+qxs5Nw4vqf3PT3QFl8g5hrUUhH5g22G
jsWnSpvzAGI0pZ8QKIua2TVkAbBcoBlzC+Fsp4v0vwgXYgwdPV42sgP4dUSIWQZU
FiV2ph223F1/6Xa8TvfiB4NkS1GUsF2toEc0i3ZDHJ1vExrR6Q/ckJlbeNI7gKal
mR8svhhjtf/oD4On0b6mi9PvgVYiCYWtvxznaLSIE7gYAiL5Ju6UbbHpOoW5u1j0
oXfxKbGG8TilDlbXDAeuT7Ogy/qNCdEl/EmPBHX+qXBKUuL2vchHlElOR+CfBf6L
7rZBHlbOYZl7lZps+IQlTPGuSIDYvhz3stPKoNr9t+ZGOjivGoIMSWCz6spH4QIH
ju285469m9PFC98ug1sT7WT9Umd0QRu9RgZJ46qToyL5fin0TZiHqPROR8UU053+
FqQjSfB4wYtshMHzIWB3IkXsSf5nS3J+iIbM1j1KJUP782wONvhHFX1uGFx5q7gP
HFID4MTz1YcjuBfZ8JBrHTBECxM5fSVdgeJvXqvLFhqFuekberZR3jNWTOZ/KrTD
lFj32eyKilDYGWdE12se8woD2n2fRlP0Lzd2jYsc/+NieaiChKETbXLmH5CUJKRk
ebQR60iRzWG7PpIQ+eo1fAxIEgWuzU4e5TouhlETxxEupAbcu2FgTjgsF1sWkgth
y55lseYJMq+fMD7EUCkNwu8MF6mx5ksU6zL2/pqOcj/gvDWPrZK6e36YnQHCzZmU
vAgPARfdbdqXKNaOrt0Bg9KNH9sQChIA8/n+x4o4exeQ8ESmuSufybpwdkg93aXt
4uEmJUxHzq8rxOIQ3WVLLIK/l2VIkiHAJYZ8P21YkOcmWVXyUwL1tX0zYm6MDbqB
CvE4RIoqGOpkVdJWOuqpmLXroOLiW6jqq7umHO9XxbwOLS3oYDsvnosqL8NFIs5z
UEeg+86G3ySNyIRQziCF5qw6Mc6NJdnoBTce1m/TDDYFIjoA1o84zQCVhe3vZEXb
9WVjLJgPgBxNSpepuhVcyEJ1Ya8kSnyzz7QAihw7MUfQwN1uoITuaPtap0xJHMhu
uMz13fdW7uI553Wumh54THgTsHuE/exJMVQiznSwbMmp/TT3TXqPvKcUdYy6JX/L
pEj5+kOt47ZjDNBUUMtCqdnFYhCLuHhaSetIiZneYNaEMHpIJOhK/Hk1sDIhhMfw
r4Ite5zyZFITBK+ilQXEoeHuOtD5QTlNTSwnAMYsOvtKYDBrcl1gbxXrvVumNvpG
fHd74K9xutRI+ui+Qg04uLv1EOZgOn5g3c8FfF01FXeHdtTr5yFq7wWXLGl4xtQd
YZsYcK0AgNQW21ghI8yGoOM7LmcU53ns3QxUKsLmz9IRw6ATqiDcInUnIbn8dQGQ
e1EWLevAigys69xuxGxQh0nH23WAxBqq9/SVEWey4GXYZQ2dPLn5utdra3DqeoKo
9nAXSx+iPAPG/7urz1EfpGpCdiRuevpsQ0ZvvEXEZr6DRbLS/QFAm1deGq2OK9+X
iRhIZQORzYsYrsUOHoVsukp8pGgQLwLmI3znS7p3ReK+GM8fqHwCRI5W7w6wZlOp
H0UmBx5AxTTz2O71jjddfEk4PA2kQK33UdKZLfJU4dfU3Bju7RjjeUpXnVI4xhcT
+hCA+OqUeg3EqPeqHPBAJlHgSozjz9kJ8/1mRo4csz/a2DBGFGi8CF1KjYG/Kixc
EeEOf0Qr18wuVHoJ1kQePJqnU2M7iQCI6zftT4hEB2lJzszYYxuYjcToG0zBHTFL
f/8OUYh4ZAgm2Ct7tIagEe2NOEW64WTqb+tFbZGxxLFXwY/WcD0+7dPIGkskhVk/
J7BnuhH+5dpkEXHBu9D+NILnIjc76N7YOyHry9lN7kXWTlZW7exnO8O398kQf6DR
Ht+a2IHYyqbCL+RYZ41W5J/u099m85n6OBbHj7M1uauSjRzQkXKnn+/wh2xsm35T
foYy3ck+rThZ5F2ZkIBOEvpgEoTNki3kOjB724Zb10dHeD0Uc8GFv013eJ2d432S
hjCTje1AmTVciKmQ2c/VMeUutrIv71H3L/cYjOu303az8ZuxP7h/l4eIGhahhS2Q
4kXZ6RQU5LlchA17igxS/FXeEDm6q2On2AadpNS3A/34+fnSGMYRmaEnTuYRUCpx
w1PqHY9XLTSaK3JEzmk4cBSwBIX2Q6Dpmzh/5z35WGBCRPxBnlgf2rtOIRMIAPAI
g3Go9p1JFtQjDlqHlZpcmtjvjIua69dhWBielS9zQSw+q2eLdAcXxgTHSyhRWgT7
/xiS0724YHpaR789A5G2RFJwGljtOGxwTe4mfRJtHR6i3U3itlvuCWSHyNJMXDQ1
1p7iabeWH1/2+xd/yuFDrdyl5a3QlMBw6hEVx554YunxA5ef33kqKnIYJS7Vg+Te
k8FfocRXM4i7GbzZTN66ksQ6NQv1Le9pnNi3pcvvhw2c7qAl0Bpk6/deyy6AN4my
Sb4QuXh9/AlysmmQ/G1o7xvyCNtWhQsyjv0XpxfXYS6rvmQfrE0/mEprL5/3wTxa
SLsNBW9g87hCr8WbETFuVjBN6hCFHXxLW+OqNgZn3511AFwnIu9YRxtsrrOLKRVj
qiclb5W1MQyF4XHUcxRngEugX2K9C6aTjCBfymrH5i6itObOyqnZOZJLjjJmuFKf
+/H/IDk6OwCI6qYoJ1P3prK3wGIoeI84c0a2ubvCBSWH6F4v/5iyOOagOTJ8WOxr
rcYX6AyOuTDqeLl28vikLjnVcjsNue+XWGFD1ySB3TxHXjK0oUIeghVpxtuPNmR8
bo47mFoLHhv3MvrEbPkQlPQ9resRAuc2iJoHx7qIGMdXwJorFjjubxBDPz7lzso7
sVY3GUC4Ml/ENIokbFNf7Zd94AXEA80T2pA2oPGGzZMfYqfakQ6TktvLrJci2xOH
zBQhc3aLp13PpmxoP2B9ZCnOBcd3/IShJhoqJACo9zATb1Q4VuATAC8gYMqUc/3/
ezQpe/RvZnbKK5tcVdHIOlr+rzkeOypSrBDOvsRTvW9MtOqTjVtrG7bb4bI4KsFi
YZqO4tgVeU6E5uUjPZuJ9hNdr0pr55w5LMMhLsPae9Lm/Y+JXfUc/wXXTPRgceO0
DNXDmUbs3IxgMXGWV8MyNJ7vcXMXo0IsqWM1pgFQ0pfQjER4hX2NqfZnuspyOEuw
q9i4yS+ttO2+RTtYe5/dt6K6kW6YDQdWD9FBx/yJ4oV0iu6FTSF4n0oha8Nbb6p6
7GCdkkkNPpSbeR5IzhveMQlGyKZA44LXMHpDGziXQrJha8buZKR4ns/FEJXbb1Jp
BTQMSafTJ1irJbq/iUv4KFxclaVT//GOf1YNrZIJ4BXfp3jaCRu2Wdi7thwHUsmv
2klpME6q61oBxO2B/0omp3OlYuB1pgbzr863JGyDhWPpgfApkY0GojwMsOc7qs88
fpz53bYfAUARjis3tSAXyLf0czi2lL6c6M+LyjevwTxdMGXt6xhgcSKPyeHwVaaM
PovkddENI86MR9uG8qwCCszxiGRV0MAEvj72ZwrqNZXQzOgIYQyMtKMDxKMeZtzt
dn4CeevCBiC41/NDJ+nWWjQ43H7L1S/5+6VuYr4DWfnXi0NYPfFxUldcUQ6Go6E+
lzB0RtA4BVRanaaqUSr5Fh3b9e8XAlyDuHMBB2XwNu74YHvCpEAk6JGN0g4fawHx
LLMm9jl/joK/8WdIaSVcR7IrtuxJhMV7k3EaL2N9My9sPTMpZb/h5lMSiNyZN97K
1Gidj5nIOJc0vCZdFQpgy2jK3Ske4+s2InrogMw5xVlrN21OhtSXySz974E6v3PP
3E+H14KerAXcwqGk1aku765qOAieFX1cQ5pTBAoxvJT0IvnuYWTmUY1kLLMQMI2R
uJwb4g8PEAsuric4Ojn2TgiZH60CX/1qCol9oBDNVyDJqEY/sC0vZ+RyQblpvBrE
q0IjXAMmqmUyYiUV/F8B2L8mP6q7PwW6F0PzMniLXq8VG04K0XEMpcQ0ejInOboh
pPeYKVYD5x63gZRLO/s2fN7+F/IIFQ5k/JxXIw1aUaDGr7u4OZQQKE/AOmCAiSZC
3Ap+gtDi0HRkkN4CPTcAOwjrwXsQx0FrNUiAqz2Aq5LijLKDvmvNdjpPCq1JJHPD
a1CspdUbrjBYBYGYCNczirAQo5bu6CKEeLW5P+M8UyWEBq+McCCr4mFcc25MKPXq
piEN0lw/zZ6Er7ZU3oT7BFPFkfgESFiH0WxUhl5ZkJK/V6RSdpFOcEl18BXL2I2t
iqQreBWGMwzYd1Kk6aBp2ObAQSv1k12VBj0T3WQxLZiy4f+gf9M0/NkNEa5jut4l
FiHyVuMrvIXY18PKdZfSPQvDhmgVeA4MJsft5amRXbKJ0MgjCyQLfb+whet01epb
w/W+TFm/whvt2RSXD/jqTl0PHUipmYRHSix/exx3u41LbTKIuKQ/7l8RCRzomRpq
lB93wdSI4oGOwYnmIrRUBZeicsmHNMy0/1eJPrG2BVQOH67n+6dedBpRVUx4ykqp
jr5fM4Lp2hQyHfwheLwZUkZ72bTz86Yhrkbztd27rr2EIN/cDlvzNMRzc5OAiovq
fzYGDhjUqsJGqpE7VJVNkgH2QvWhNqX1QFRqksaMaSdPNmQyLpHEEuWM22t4uZCl
glSBHaN7aF4VammHloSZsLtLz0Pq62acSakKsScT8aaCpEbjnzBFfKF8hl7OQS+S
53GWTqffOawWLWyaTtU58yrw6sEfIH+r+0UeS8ZvM1lqMfP+lI3jAPiHjhbrSQ0B
rrLXB/+5r/z06z/QviwGm0C++OuNzCM5bOatefb1KwG7NtS+vKNULgLwlekyva4e
0lJyVaaRxpSiXaFocafJHHOGRJViqDOvzzS0+KjkrWUfTHudqn5cKSIPLAopyeqO
IePW2StvxLvlGscu55VuYxLn8mLP1IfrV2r+qOJrHg58K3tJLm7ZuWQeN+jg5Kip
HSrPl57Lfg/u/Q3+BweGBjgXeYY1nEgrir5iAJv3Exp4e8CSvTaWVZ8pWoIOqs6+
cJyI+S/o0DYztSnerEBvYRMnHW9iZ6QoTd9P+UX4DJ5xPlFvm7tPOkYSil7akDrd
nvLDyNkXft2QT4QTzhjXo40UXMRW6tXBLy6ffLW6jS4m3pMx1nznijClpF4RD6xV
VJkPqbBHNUBaLqXKUn2e+2SJD3IasM1EWXZC1EE9rzXZ2secZenVpQ/+2lgj8YLr
GZrzDQtLSk0A2A48wjpQhV7iwPD3NONh037ZfUTx0FLR+/jVYfMZ4NmipHsNe+7l
DOs8wLyqCcvErpWHSYmTgIsN8JNYabRnYY0ZFDrPUN788TIM9+wYm1kjNfcFTqJR
cN8w/i6VESn3y1BlQ5lcOHgiOC4sUnWq+2QKUAJiD5/NHxHi8K1Z+MNAicPmkpXb
weR8tjjVvPISM0pxYLjUo2ZVK+Es3S8KVbHZOFMbUaIjXGWfPRUtv+7EjsT4gbkF
6+hmrj5eZE/RdvRFFqYu8738Rt8YAPr833RVZj/dvjUVjBXR5/cczRCPMMt39P0V
FvD+6jkzpttEwirm58JKRCV2XBoQjlBBSK9r2HkRjyRCxCXAfqZEV5g2RVq84iSn
2JUnTvwjiKo+nWCbwbiZJfHzqdn+G/O5+e80B1Cuqoejxvuq7p9Wee70KNRhEqVx
b0sA5cSlMNYNOrlU7RbTlEz8dAnvBi/JX28xM+H2R971guuNa2OcId9YMR/VaxR1
sXfP90bOqnQndyYd59sg4PsI3W9vLZhaR3+QBOQMWvhVrIFEY0xKiu8t0CU7s7yx
B8tnmZ/X7JPScY85pTg1WNAh6d2oV3vJyqxktRtK7GjRxZbtijGq6brsT53VvVZS
T/r8xuJCOtZ7IfKlGBbKDssM8MewOUCulvul9b3wnyet8KTyszElEP4Jy2ixGk/1
Sza5zVr2UH6C22urDqswwvrhiJYFRrnrBiiCXFT9suNvRO90iSivgU63v3dH/dXk
S5IdK95e+PwkcdUak50pjEfSnUdge+CUWfRevibtO0YyDg/NKD0ecKhTNkUCW2Fb
Si5h4sS2lm3PCm6/MFf3hULNbg2nJKpF92M9l0ZFGkeVx9RHnCuR1q1sk6UhaacS
tg3VTEHeKWKSjSQLx8B/+XKcLiZr37cudnMq5rns7iVT3HSXYjgPFR6/AUmv7trn
hjSJrZwUYxPPf3KQ2Q2jou6gEaHk01d2nUV/QD4TXGKw/YYoEyNAH9PirJsR/BUt
ayjCUWGGP44RoKMx5Iv1E5HoBnqDCwIBxh19bKINvKpFlyZNCqfQm6hVSaVYnahm
8UHzD23uP11wcmCsBNf7NTqXuiVQzDVCL7xTRVLciKZpuyoEQlD3qPpBtHwfCE8E
xklztbrE2VH0oXoTfI7z4FAjSpU+YfkJl35v4EwkUV1Q/q1PZZZZSr7uZweRUY+N
QyFBHMUfOhGrYni6KpI8eK1dFI4q+u9KaSiaugEBGwq+NKmvU7WEQztXOrmgolj+
FxVKNoXIaF90IGaMklHNobb9A5+ZpNEuHLfJjKaf3JAPQOSWcyVvKw4yjYA8Y6+B
APGxHYg1ul8l+UaWzAJ/eGPTxDYlV0afJ5Es40l853qJe2kxUOB4TouJTMN05fcf
o9rnyfGh1dp3AXj36QilCj8EtqJji10EkkfSvstnWmNbWkWuckLRiEPiiodPuAZo
jnUB7qevYW4erZVuRNfeiltNBLmsKrEEOu7WclsPOdNAPGD45RldwueAv6kI/QA8
RDppEBF3Z/FRLvSXQI+LMvDJoWxJBd+pqOrPdMyJHvpM9r8EHzZh4dhZoGt2bnmY
TnRBWEEByAIr77K/hlUmQRbG0y+qZ7fZy1Pm0MaPIOUGqA7SSzgskgpONAMJDO5H
F831WgDhECIUgj8ZRdfDMzcpPR6dHVAsZUIEXTb2Y9uaCrEICzukaoAOOGONXZ12
nh0gsEZBjQqeE6DuFleZ3PeH2KerISpxOSMbzFK93bVu5OaYX9QSgMqtlbD7AWv9
4bdkMRyO+a6blRjGJwI6LqeOhMIODO+tSkaXUhAARdan4QfE8l46+q84+vHQE7ne
PVZ5Ph60+Dv3uJR82kxvbCCVGmOoKMTuhvJvV6lll5L/QawFmWbHoJiWudTZZ3Fn
+B4qj2rioPWNLMZDCZLEeW8Ck8n3qHHDrU8Zdy8SIzrsxB1v3zpQ8WH6ZFYfKaSQ
ZeKbD1zKKrrWAxEz+qikXN/s+G0dXc+beu695ppdvy8/ISKqzDNHJhGxXa18yCMA
XY3kdPh90Y6KHL2Ue4grkEtWef2kBn9dFjO3vJAjEwFZDJh4AxpD/sh2V20QHxo5
otOBcPGkWAY9KgB4l9qXW1p7nDVB0YxkrdevrjBQilEkMzMH0KHw/gzmcJyPkpX4
dME4v7wEmDR5EN7vG3/OAudrsSZsedKy79OeBN1d/U37KahIP2XZCTS3m4UaG274
fHyLCxo7V+VJgTfoTLnUDSWAcjpaokwd/w4A6HPjojKdFy0LMTlbWtp9DbPb1lok
ZrwcU7y1ZVPOl1nfImrjBN7y4Q5xsZ50W67C3XTwm6/Iyiz5x3DR73NoxfbIqo10
fA/7LDXET1sb80VoPZIFMO/L9DJfWdEWzBq2w1PqVNmz3CL2Iw+CYZ9c1NkGo3cQ
ZPrWXqN0mxpNCSh8ATl2A4RQUcXGpRyjSKxQdh7Jdu2h5ntg5rQL9AiJA15f+qHi
81FD2XTaZ3c9n9+ZepH+k/4GiK8er97P9ljc8QO/8OwmCieKP+QaLY9Jkwi+7QU1
R5UVocmVMnuXTKFtCGYBcann12ed/rK8FndrrvJzAhfIgiwpUJ4BKA5hgDJKORVr
xl6vxzbOYNDcXTVBZQHI6phGwjlRUSqCQvdeftQWFxTIumyqb7KS8sS50exxN/iC
HUpjoIdhfW9kfN4ByVqk/GIr33SnryqcTdXRgK2L8LGnPI6l7NFdulpRELSkdy8m
cSWLVJauQUPFMD0uYdiEyd+YTqGKV4VWQ8vKqPd13a9qMxTdGOdNM26JYDJvy3cH
Uz7eWzJpYFnrqsSPkT4/7UVte1elvW4BhzyLox8nBUNP8+Da1i/L6IapaUS6cxvC
voCNLLhwQi1XKqBK+cjFEt5IlodhluAvstwAx2ccW3fw+M4OP/HDPZmJXGIykxlY
vdgAywRVrlYG2XDxFtEW4ILQf/QCcGk+BbqcirNJ/0IHJtlHG/4fMmBR6fp5pgaU
3qDksi1CXdGRo585HbzyAlIqzzYHe/90jZw4Pn0WKamnv7PdtpiDxsXti9NW6iQh
R35/BbFG85VVjee8awn5PC59bDyz7nUQZ59nf23oqUpHD064YtwCs/i32XiLWkF/
Nx3rNID3vkltk2FWY3i9+O7070pST5KjUvuHX2A4ZGdvx8uJ0GkWv40PVO2+Ut0W
CODJhokGBy5uzzWzmlPhYw0RfJUm/Cbw4bpa0dvxVxNVme8+5ENU1j8ehjDDPHw4
lhr7iBfj9pOFzYvxBu6MAdE9uBseb2n09i1yZMyBLNIUZ1n2FrtL2jnoAq4aAQsr
iGZdC3S8uXqAUY74OlILWZIBagKeOpkn14HkKp/h4MXyrWbHtdslcw2GJsk95C7+
HbtUvPW7N8D4iUhm0jMJNeW1dCV/9RTPyL76PaTaTQAPudcqEUFRfFivpdC4b1FD
QcElVSFfW766Yt98Ymhzny+EWPrXTCNb9NcqejJLPp3p4lXSvpf4MafSrA2bxUau
47g84yXxVlpRpWI9++qc2i0rshepLLr2m2CMm/KvvQ/av5nNjgtz0ADLpIOfMAOn
hwZ33L4V2hgk2n0l+XtmoqXZlAsrZIBFs/7KJmI1Mx1iHLq/Um0QrZrvCCxCTzVk
XIVH6UKFJdutSL9GEcVG6cXmPJ1ULnTRWnoAMLFIfzHVadwaZ5pImVGF+Xn/vDRB
hw1PJ/ivEv1TZmQFeAFiX1Up9KyL2lOZO4Y2taTIWR/mzzfvDgfJ4wHRMFrVZsku
Dx/Rb3OZIrjaLAjWZf31emp6/yXrvC19TP3/B8KMZBwxTORNHzZNvcFa+DBDGQyp
5nAjIExkCw1JMFAVbVkQW7zEmAzOo3PdTpN4Ox9Aj2+H4gasmlyZa8zZG0s3Ys+o
JqzHYhfVi/rKrkCPdpVMgm9y/crNIVm5O5IJh9+Q43sIgO/aLke3Kzb7A3XRcDhx
cgI0gWEOIMMhXFQdfwBX+UwzCeLkMQ7J0CYTyyOFnYIfXaGRp+pUcI5B74+lEgcA
wZ9Gs4qy+V+2C0yoVQh/Oxa7bpMU8tylN5N+Htg1GWmIFF2NXE8MLFOPle4Pp8/L
jNV5d4O7opv+3GYLuqyEGHrMPSqPwZ26uvQU/IhnBzXUEIHVH1JZQTCwYTmOSDTY
LnIb244p8z/LnSv6657KsrUyCH1XAgxf3Nmnj6pxres2VLdkc0fh9+1AokZxbDfy
D356sWabqNhqWMXmxXbB/ESf3TO+y6EGwNKoOAMjRXQ0j+0NhvXUojWgWB24w+yo
MhvCOVV08RT8PTMcXjFd/pDKgcbBA7BiJ5FWvH9eQKmZDsC29y+GE1cVKD9VGD3W
9CvcvuoqeqUhlVR276iHY3lxTUZrFL5SPFxwy5Gh8aZ4PAFrrGoexWg1BYgVNo1o
I1spFMAQMeX93e0Ud6IAhmHs0w7+hYvQ16ehE/sU8rHRPBWi765nBqRIr+9744kp
aFlrRUK50TkaaOKxdgbj83/ZLvBaQjp7+mv/xP0CSYH5niSRWalzKT0OGoKuKOtZ
GHQsrVMZL/ZtD29J1iLeBE0df09j/4eVRSqEGVXFgrEzKJG5hSrQ8iK2ZFhT5We3
bD5SW4IPF6Jxk/rocejoMkRmTmEoxcIr7/bn4hejs3A387mi7g++ChTeySols4gq
cYFsxOv3ZOXQCSicz4vqI+ugO47ZU/mnGI1kU/ZPBvw7SHIqTqGOqg9QvsOD+40h
a6/jj0HP6n288GpEIc3Ozbf3WuoNQwSo8Wmwvf5uhzACDupohC+/KYDgH0lz/YnY
p4n8qa8l8LjKFykTU0HzkfghKcpkmNh1xgz8cGOrr5hi9SKeHQC7o3Ick5GDmqLT
8BXyv6DR3AovHjbPwYuSHuvTfHJ5MuNFx1Xuv5NnP656AfZwobBq/InZnkCyFPXp
E0zynRcXjrapOYfGuoUMM9HkPubSD3OSCji6ekvuwion6YaCBdQGE6byazFSvOs6
NCHSc8Q3N05eBzOxP3Qif25ebXtffD6E2us4OmA5zY5gfmjFxmPTPXNuwYVLWZ3C
JUGofpdK9yiAHaYXn0FJcCz+HzunwBBz02PyhtCFG6pDDp2gQzr+Xfg20tipcdQ4
/sC1pkl0jmNAhrEG4ykRW4PG5uDazYVH66CsbRUWB/4IYUlmqSsjLcr56LfIjfCx
DJW0bo8tBqcq4mhGjXLg1eLvg+35lvc4r/RCYPY4q1seOLF51NNIan8hUhsJ1+fG
umKNgjow/t3Y4fNWY9Oo+4MW2WOrugl3oI87jVcd1jC74h2ChNhPrHaoBWfEcP/a
iwgmuDW2c4H7SFDlEUf28WJrzGJZE82VCXi32J1k93SklgOl8abI7UKtXNGl1ww2
hNBcAh6fEmuKdm+wV4NUz6OneZEXNwlocEKAw9fv3puI+SW2ZmPAvXYZ60hVBDM1
Nfe1D/lEqumKEPQRI5ALn/AhrV1nBv1a2Dd8yXDht1WCql3zfPCQIUYCdoxEESce
YgS8UbQLt+JUC6+BG63tIAARovQ9asppgHwgluxWLle8vuLMOe40p2qfj2rsVWds
Fmly15FbVJ/WnjCTIYV/MeQI/UoNmOjw1xtfDXZGwRT2KexUnjp6kVtH5A/ZMZJg
u5gczgr/ogNYTWz6bbo75uftNP7w5Ilr2Md/P9Bx0Ucf5KgOLtQqVgEh0S0swWuW
zJRUqNot0FC7gCQ9Mar0LFYYw6+A23XMmaWwpzdHDPvgoC8fSEcQS5IYuCe7nFli
JliZeCHn/ZkXUSX2UFIMQGPShM6DMhWCW6YHVS83lepinJJu19WzEfROr2uDxb48
TG7V7EYG7YP+WeGacGHMxO4LqFyRGmr69FvrSwcEdnp1C9dkU7d2lRrpVCV9Zidq
SzCrfj8oXG4PQbuAqU8YLctll2gpqkZyOpd+nMKU4JuVgBWFdTwu7yAAMQj6VNW6
89mefvl4Lu2BkyA6Fa5G6C2+4OWMPLYlplHLU/6M6U/qZRtSj+P+BU5rAQVRol2O
ZSj54XvuXldioRB4oDDyP4II3NeMSJooQWOkQ/p2C96FdLEJJIcMmnG5z5bLajPt
JhtiuRu7CCQglsiu7+wvdRuGVC37NTiU78/ETsJRnzirXIM1oE1sq00uTTaScYXU
v5hBNkxrUSw+r8y3OXieyf1T270rwVFumqBElGIZ7slXBNISug4n8iWI8AMyoV7Q
eLqWHXpR8a7NXQdB04bTxVlUn+1sHJD+he1lCQAhluuKW8GZt893AUgyUG28RE2s
0N7R5vkfJPgehqOB+s8q14jQhZ7ZGB6NJYZGHhgzY/GQB66HxCJ2m/xZqiMVpGCa
CBNrTUc0/dsefPKO+r3jj0tt4F28u9CdGpU953kUzVrPKtF+MRoGc1eTHrXDSW3b
94Wl7h1AlKHoJ+SQiUus7xFXo4d10TbmMRMW2ded7/aY9/xJaJFEoTQX1lrDN4g9
XUMbNJ5CO3HKz84Bw/NCcPoKFuxEMu0bn/9wcbg2fS8/IvZOUjVce2hEippWa99A
5RdFnrO1OaCk3NwGt1DpU5fW957lrQ0L6u+XzATkw/Y00BEKeivOeatZrhzuvlPI
1CVa1JSwlrylFRDwYBs8VL2yZuORJiXpmm99GxHhDJoloXYj+Bh7a8XAPfRxTaP2
8PzTISruRPqu1fZH42ssa/02eDG3pWR+xyFLwdkfjQshCvIbucMJesSVJEru5ndz
0suScz58F9+HCJeBCSH9lX9W/WUlSVOVXzAa4n2fM1YAPsgUxfFmBCwurN+hMv+D
99JqU3uUqQglCgROh3oqx60K4m/G4JrtJSz8C5t1yzKGdZvvoVjouYj9efXr1mAQ
2Elmk22iqLy0LDti/Qec5Xne0sxzuMD989D9xnBiWrhzITqXlZKMyYlMqK5mZoei
8S6WoQEH6zqS5SJaUus32UYgyYkgWr3oYWedJ/BbLQ5iqWQ2AyvyrJ9MxqiZUaMW
iKYI0lwxqJs4ktnb98Y9DFl4qbaovgZtC2Q6yBXmqGMlL6vXtez3sPaKQYO1I73h
UfBkNyDTampiaSiM1vSvUymR9c8UzqYllVK9igIkY+OyKF9g1nlufv50aTrgG2GK
WMbW0EkoCqzJdr2U82rSni717T1v4hYxXvm92Gy6K5WfRHxG2NDzqIHxoUBeegpL
/+4Unb27sq0LmBATaLyJ65ov0YyDtDTEy5OYVdzzx3Pp5a3jLChfX0yI/sghSs/x
reIGSOsHgByjWOfiJeYM6XdUmozbMgpP7eUcN98xZePPJRdZtmhtpjDWV0kipKch
OFnSSBfUjqcqR5vkBbu8dvYg2ueI+ZDeSDXwOv81F+3HMEpWAZpv8Rjlt+NS3hP0
rOil6yNen54Loy8uRQ6vYKSy911gfQH1SAE9Xp1mvHG65i1G3SfoasMybdPCBgsI
1eNeahxRnVWUGF+fD1lkpymABHIf82a/tAh3/GxqBxLor7XIDlEJpQqRHFfCzh+8
n8FK1yQdGkUp2WWj8iybpaLwX88tRCNaq6xj7otf+n0UUlP7GoQlSPEwt+MZ6mUi
Aj0Ww54eSS4nOghwkPAu7JtEojVH51wZ7MkosX2dflUC03AuRKrQuBhmE9xcr1cX
NgZYGEnfi3KJ8hCDhjQaXcrgC74s8d0QOhiaDnBTbVTPDMFGjVrLQK/pjBN87hhE
x51h2khCJSmXOoP38nMNSwdBl1VvwyiRpoOMCSDcihEpvEg34qO/MUzD2QVTXk0F
IQioOMWrEFoD7oUv+x5qj/SP+Uf7sHBUa5SOsjSKnQyfCwZywm3IU93wYzad8CKu
1xcY27FaBTKah/TxVng+rJKoLYXyxW85DQ+uzk4rTUN0tYm0c3+V/xapJgqPdjjC
wlKav1Btwceczw0UlgwFQfWmqezF6cX+twSbAxyRyjLqaSWdNrlhwHE6tuc2FXwx
I0fce2+TKYMrOiscNLN48jj86Nw/r0enA86LWZ6R99pvmOZa/W4gs3UUWPCwQCEO
mDGaHYNFBqH08ep4OuICsmMi1Wg0taz0QkV5CIafIGQj5mUcRcU5uEhED/cu4hWg
xT+IfLwMNspOJCKCXqBVlxyauZ2OSaoMNTRMU0P2e5Dni0WBD4DhMjJCz052JFJl
Zu1ajrUwX7n/IwsW6G8hPISbw17sgW2ZC4HI0xKNRs4+Q1KeHKS1Q9N0ibm7QeRj
tPJlpiploMJsC4siuuPNXX0y8+VKnSTZiTUSWisZX2rYdFNXAQoqy3xSy1mJqMxb
ZNKNsZw7YCh2QansGnhBO7XawmP1WWDf/bR83s+BkSGi9TTHFiXLDTVTKXOWXIQ5
G36PZdwiKqyaJN0pk0Iu+uxWSI1ch5/hFs/vOlmYoyMsaNfkyxaLkAi5SMXO3V6A
bb26heRekRzESEasxiYcWIMpQTIgayF0hi3rseeKx876WdJlfgWR1Z44BYTFiIT8
PDyd8Lssc8rAeDreJWoNLURgSnKY7dwGczQiRhGOtxnv1Ef3kQVvbjMzlubx7pFm
rk9792DU95NCW3fPPKpkBFJEiRRtdaBfgYuOq7hh+D1HPNHZY54MJW5EuPJP4wR6
xO5hSn687ZsGIpTw2fLyQ+bchz5jNQEumrH3z52i32VvRiAHyh7nLu1tzbCF1nOl
b/p2MCcGnCkWXMP3v2Q/QectzB9usOKXVovGzyK0ELOCA0mNJu8hYlVUIuKcPliW
JXaJ9XRBG/Z2O86zsMaBh7nlnlmg3UZJHsqzFHZBKnviJN2btN+vz+P8jIGRaban
Zf/J3+0PReHB2JzfD8McvBIIt4HLi2bzHoyZOzgn5PJpGqSZsACQZPo/C3FuuRBe
e+UneqmyFIbbxJjaoOzet4PqmBlJuZHTxAE7o4i62uJlq8fZhPZ3+wXUBW6pPbcc
cXh0YpXV7CwLnIbWFPTWiGbWjheV9mQ9i3ZFMuR/ElmBj3am4wAqu+uP6ldr5hD4
mpVpY+8E4Rz+/Rk2SP6hcjXVeVa9cMo9r+WhFcUTDboLer2FJTcENlkhWNEm2Ji7
ft06jFuV83pJP49mYYFcu1NPwwZLXUzUOZtvWFseaoA3pxLPAg5RidGCA1mLJ4aM
aZ1w7Irsp7Uf1olcobc5NYS5UT7X0L+gTrFtnxUcBImpfcySV1DLEyOdOO3nefwn
UP1HDxyQjog0ChURGZ0jlPiWgiGzJjbE9U6z9qJsURjUtxRK6F4+B3uikpQS/Wkz
qlU+cUcXYlIrEhYZZvHZTGhsZKeUpsLSxLK4C5reO4RwtmtuSt7XBGsI8CYhhCEp
cqe2MPR0gOldloFqA6t4RXU855R9meTTC11JNYTN2qJeFtIo8NjgKOArDcESnoKY
EwzuKNgFtfzBX0D2OVP18Wc1yHKLemeu7H3whEf/3HPX35VoS7c9Hwlzzs3Mw3FX
9gUQjf0wUmiJck+QfSUDMKdskUKRhh+uI0l+HSbQSnWk/OcpjKEKbqhMcl84H2/Z
9BeTHwJ9ResrM9kFzDgrLKnsb3zh21/zXDjlsFbZxwklghqbfeN8Q50eNqWTvYf0
Magcn8uPCFLqZ7r7E6SjUZdMtgcQQamIjWjXwbmRhryknJckKxpbXTUCeCj4Rwa5
vUKYLMfa7Kksxqs7ooTlmf5dvfxvXAUSrymsaZAm4PCRrO3kILwJ+qBZPIyQFsA3
PmIo75AmBCORAw/fl7cICO9HOOkcXdOO0fvwFHUtxjjeCJJCYzG1bXI3JBPbDMzt
de064XhKxY8h+f8jURDhHdhgVBju1QnWkFXVpAnBPMBaujYAtjGeFb+hsCv+knLY
YBSPSMRLKeimw95MBIgspGCsTHKRsznrSIQYrpNjmVWQzGgagiJuA8kUqLVkQmtS
f5fKo9wOEO8AKSdXFxHZgFBty+A4aGW6/FXb6pK+84aqe0dqso2dOdtQq0yFrfHf
1EwOHSfjViUocXphafz+wnFwi3XWKks7a4lcjXPf+nSMQcub2H9i/Uk0IfrzsB3b
YJAd00TW3yNzkiVDayuEl1daBsi0/jxtWolUXJNbKq33v+eU2Wk/k0uLp1vywVx6
fRROAXcyr1u7L8Na3nSzmz/5G+0FtJKHLHXEaiJ7wxaE13du42kgbeRR6wnQvhWp
UY8boLLgl0fSdo/A58eC7NwqkCbF3e18NmOPxy6cXhTy6sxiS+bY9OWMBC4cov52
QYDVwdVP9ZrlgjtX+UBO0LxIbvErKQHFdi97f03gmCJtNq0oOCA/8Qjm6RCDux4C
FxPHqSBoci9BBt575u0LHgsdc08QdmzU0xtNyMKRhHH42b6VmOIqGLY+JmRLqnVI
dHQaeQDPu5EVyxLa+GbEGGgYmVYfi3E0t5NBbB0JlJ0adDARSh26nP0mUzobzsbv
bS0SolTdGLs2qexzo+bWKZBj0l8c6asMmCLHmNCHGfuX38YbOr/thZECcaP/jaIX
qYxsw/kkCtrWL1g/XEXQHR08mt61dJby5ElJUReiyepg6OVAZUjxx/2Gnmd+Y2US
dwkRKf8FXjDnvng9R/Ao7pOiDNFcdsBQ6vgMm7js15qzYPSA7mKJZC7idftHd9oz
gfbd24c4Henqd431bYHvnGg2y1HfD0wASZhOPbvHqrJv19RoCSP3PhUlZRmC0zeD
AfwvojrzU8cOxB+/awUUQmch7EhdwMeEw/hhxdS5nGWWE0gBzAHb/kHxzBs9QYyf
y3gYMAnD03h6C/ir/2f7tAhBP7JulER8c9f2IL3JYF6+aWS75Dwrv0HSpGyCaMvh
Sehcedh+nSdylG3RX6oqXLuaG5o0NhMwwwg7xhsN4NaoG8WOwFkfaupqfjD9e/E7
bGBY4VOU7dvKpseKHzvp4JtzFHLsa6UDVuAylZ86tDtknA/LxFz8jZILcZ44JsKc
UvoMLpnM0IwPF+LnSd8cd/5hsbtqxSLL6p6mSi0XkL0ee2GGcYXSOMJC0rVyDe4X
Lpd/ufIn7WLoVcKpezpBc5e6w8CYYZUQvzTw0ZjaJCI9GJKimK23YFMnzI0ovdam
HmZGDtGfIVoPEdvHleNKR4wtbrN+l7vf4r71X3YlgT4GFLoja2z4JFFR1aKu2sQB
CLN11hLmjHKDmZ6Z9jc3oHfsos45IoMyiPMz1FpayAOIfQcQ4LgHMnhpvOT6oCnV
Jd4X66D42FP/P+gWdj3EH1jtpg++nrHckO1JakNMdc2TM216D9W/pyBmqrp1XKU6
FZD9+mVcC0HCPXU5eXv8GUSSZrRB0HkYE38FX9b5v36/19YX81il/rh2DUB3Gn3s
m8h4qY9Kb7FenyJX0YQpA/4yMVRdXxm+Lo+8kOZ1nDjJAdx1JORqh7O7UmnchWT2
BHQKY1BGNxNaVj9cnt6rSEAqBnpC0tC9b2dQxdL6DEdkZ9uy+FZjOvyNsgHkT6qL
bduL5Jkb2kAQZ7zcZJmxjNm57RS0ZbDe1/L2lY5smwavpyuh6++CKgKlZc35qP5F
I58TEq6QRtJDJ/HeRNg3QSuUU3rbcViqCIWwvaGGePsNpcu55XsEn+4nrRuhpvY8
ZcULRe3yHWgRzFZwsE+4T/mz90OPz/HwUBrKf54FlUHh0v4GUpXoR2C5oRfQ2WaX
BorcWESqC3z2YZg9B7U7lJnVAEhRyTSdihfI+mRHUlKzYzZWUuTI5mKf6YAoXqLD
E5m82ZFeWOWt3cuk1sQDV7byKT2oA0xj6yibVJSOpwwskaWQyIAkV1BNZ9ZmDxh/
zcwP3VTqLf7j8uB5Fm8M1GJzET9H02VymQWt7iR9NFPiLdCqXkrQSbW8y0r/nJYa
4bmt/U9mn9ioYVmJyz+DgHCHFL8neINJU16pr85jpXVvTQt38pcMNRy+vDuZL8SI
W/wjb3ExdCXC7oaKMaAJeIde+jrWTJDV28Rz3BqJ08SHCgoWPIAQDxLFL3fvHtf0
x7VwVybuyveFl/SkUpyJsw/Wh2lxVL2kpR2C6rfMlpEf2u+7wRj0NxC2E8g1pELs
uSJpNkTqx1N/2OpPsZ2fk8jDTN3+ZjG8JZdS/K4Y/UhWrCnDZS9TxelMx3mRfKOC
LSnoTYJxP0FIgSPTyT7EXxP/5MuAdKnp5QEFpxniEoDKLZbYnejNGw5WucGAzNRX
Hg+JPCkyblrPt6Fc0ZHk7lPwiEpl9EwVNU1T8H7uMKJFc2S2m6DILz/BLxnd1jvl
qlDJvgPrP1w7lmeHEhB/iCIzz6MT/c0B8mwY+V9KVdgDcBCDubhOkHPYMjFLFduD
vzXo7ZADdaD2wDesdPRlCwcBAiNZTkuZ348xylwHQufBFZ69jxkRccuaHuVs4+GF
cGe1iGAW1Qbmig5TV1v6HWVkED52b6OFG2ikmCJHGz1UzVgVLjPOCAstJDaOQ8Cp
UjhfLFz1jcXmgPWPAwRyZYqc6SIbtjhhfr/hRfAHes6JFZ30X3DI6aBvznPRKCNN
DTZH4S4NsRntwLCnpaDAs2B8sp2LLpq7fDEiqBGAlXy5CEciiKNAqX1wqmQdPRyZ
mFaPYenUkqu/V9skxO4rD/Nm3zWXv59IQfCSABmw129NxWwM2BL0H9yfKdZ0R1ae
A/oA9w2My01ciUG+zVfiuqiXeufM7cBGxdrPfvNOY1uXb+yZHOnqONlsXw3eypLq
J9yXjMjhdOVl2FSNtaNI2vKKlZ9S4IWVMuAYEaWy8RZgVjbhFAPHuA7GpkkgTvqn
zym3DoO4W08C8PmJny7/bcZCovVKPQYWFvgvFlEqNvKiSh0zBBacxpReBS20KGSa
+K+SEmntCEk1NgvW9HZqyMWBsgtZU9z989yTO0po6QUC3PuMhS2phBFlc5xjbbLb
ZSrvN7Ch7kWesOfWh5tKcVTC3kI+wu8SPF7OGbtLMXYnFKEj/ppOqDGNd4jE42Ra
M/5LQGtlbBo4hFjH+L7MOgupP4q4l0F6ylh2YD7+nIclLwwJH9zApyFN6HitUUeM
eLIRUOzjRqs/2RLrlM2tRJWZGfLdNhHoPhqG4AOUkCxYHFaLK8o88jC4EHRBLS7w
AgvOlbCeidBZAjEtyGmX/vrx5a2QRRB96OgPgleYeCtC3QTE+R/liugT/Y5/Xl2J
x0KHnBexbzs/rEM7no7pvWeYjmdUKo/aqAK2RZG56OQ7dEQE8E4BBzUxuAvKzFCf
8UHKJmRr5YbtqlFZtFMEMuU6VZjuOx8ih5YtDJlDEDfaXq6hlhBa2BtlFDOseLh8
POqlnQL7cYMiMlNn5aBy0S6aO4fn+yMmK3vmD+PhNakdMrAb74A8X5bBDN6daj+v
cv313JPeORlWnckENIq3vc5DZ2ERWkkAORNIcGVTeMWrZ76H4W1+Pt+cPDtaaGOs
HT8ocAZ6Q2ssgOu562kJ6N6+kDdIzelc4Gpef8qSf15PaM8pnbdgVeRfXAznafaX
m5haUqHo8RkbvQFiE5r8xI9HdNQ8amErMBmaGg0jIFsSriEh54to5u5vG8kJ+YK+
JFWa2YwFY5y0gmvCSpbIGGPMGaKWO++3nNeFMBwL4mP5Rfyb3bvNg6Gz647KXl4H
Wuh4D/Fq13lugVBMcFt/SSf4R9W3jO152LJqWH2SE/CjTuzwmhPdAZt2zcGMHLKl
pxVdvZUgkXcf4riloneUSTkTRkDyESWw1AvV0G7DhKhHdt9pTMlZge6pOS+Nh2ml
kqCdXzgYtDHnzKLzgcgOrJdAzykwlJr2O3Uj1kO2pFGKbxoBBKLXDo7ipwEnFCgE
i8sIfYjDSlG7ASP6qmf69Oa/tw9j4yy4dBVz6Lk1yBj5JZ2id9zdJ/YRAfyEBWhr
vCSxsRd5WFwd4h82yacds+uPGWCATev3V6OFiFN2kV0vSArB1PgmvXOA9N46mL0h
q1sfGChe2cMgbXK4kPpeUkUhDJjmBmfcMi3EC2ZqslrFVy/ZHen7cG6jTioCn5jU
7z/vyD7KXBrk/N5NoyzXddmlqvtY+dq6Up4nMBcbtt43XSyQgI0T7KZ7E/y757QG
d9O0QJsVbjcuXTPWz3D+/zFqhNB1E7+9KoyRCKnCYDFM3LlUn/aGdygpnyn5jnm7
kSepYOzW3dvzQWJxig4EXpk1NcTmaCUFHvQlFDIYmWLnGOn5lugZ47ekQTAhZf68
spiSmWFtgoiCtCBivuXYopgOKZwOTrKQ1sajPcjZKcBVON8BV0KCh3B7zsMq+B1T
JNJ14YEIQxkNhpMCaQUafTHY7tP89RnkYLkYShtXzFJtXMutZNZ4ZMZgHYEMYui/
hAcyAf0cKQBovS8CJmcb6k42Vz3C8afZPfDBtsiH5XJUfR7TqEw1C4C0CPPj6iQ/
kcvJPSy9vgzRwiDs5QWM5FtMngSRrWpxp3FI+a9gwRU0otoRZmELpaalXtKIHamC
/zIMfvcf4f0KI3+rF0lwjO825z2DM3KOQDXURMqXeO0i7CXak5oynMoTLJQOE0Bd
RQ+lHIefOAMfTNxhxY4f6Bu1phC5fB8hKuOb1HsZ0mN/OyjOEp3kt60JgRuQz3Rl
XuZ+LpTKoIlF5iLqnyUYfN4JApcuFxpcvKgkpYoo6CUqHWURpLbDgKA7dD6G0CWW
CZwIJtiBabe3g01I72BxQ4M5k7SccBwsz3N5Vbvye9Ol1pNmsyw4MAMY3ToVSntO
BhP2FGkWW7LiW9jUj6EhwHvIRxYc2RGtS4jlwzDhr3GCVA+lkrd+m977MX5TUME6
VMlTyc/QFG+rk+/1KLrrM9gKMVqJTxwwNTTUJKW5b1JtVtDdHb8ieS2M4aEc+SF7
wH5HpmxiVIWKAgjO7dhsWgrRqHhqUYzS7/1l16wuKUWQejpTgwFmKPHfVHhTLQ8x
HUN+YuFkTbblh6h2TKjqdMkKPMJvWv7a7/YkTHEc9yJVmg00tgBvMoRA2ZR09cUW
yUW+xhZshfjVHTHaFdQO0FScIQOEeLWFoAphyOYzTI+rywHDh4pGteJUxlshEiCp
yEqWNAk9Lj/6zn9dkZLfSDTtI+cAqveVyNNZcwi6TOZ2K/DxTAjk+7qrtbUVICSK
bXjBGOWPuCikjoRfVMk1jTPlt/Ejm8f9cKwbGi4+1Y5i3bRHq4GOMTr7rmZ9BCfs
mky8bEtyF7/IPHiWGRx2rUUj0/rjtuaD3Z5UTNU28X7zfc6hjq+1KYbOerRigJas
H0d21sDXzzO79q4DkAYWNGYuAkiqeNViKw1yT5GI6svknjyqmEE+WiBcRmp9tMLh
jL4bl41S7DU70YXdAjqzuAuRIBc2Va+vaWv3QaxlgASe1jMjiauLiaTkP8G/cZ0p
/5BodMbYBOBiGhc7vaIn8kSg1s+Bi0V9Ne/WQx8J9aNTFU4+/s58glmuPVLOOBAu
anLTsMnQJdSjGGP1eVxcHSV2VHIzDD9dkpEJWhDLS5rth0UPRqvaPh4Gew7vwyu6
whcMsSf930X+sU6ZHFh7327QEteoG9NPr4LYQ1zSdwHJRgdHOtsAeHzKjumZoNtM
Z8BvxSnb6heb5eRKq6ltVJ52z24e4mxu33SBVipEvMSnVd3PtQr0qBDhjg3vqx2Q
OI/UzCaAJh2jhwqc+uw+Jwu0df7piBGfko49rbWiaiXYC3u8G/7znjFIKYQBuXKF
u6TA/zXG4DfnFUB4GPteE1Mb/NxdV4VAG/J5JV8vZ3VI5riBYoxKyPo6hRj6xQmr
f18Ex3xClIBSaCK5PBFYRV2vcITC0yU+AX2Bf2HqgpWaWzQwU5WoTEPg8/CQxWQJ
UzBa4m/94Cc0CholCUZsghLa4dad7jfoUTDJTDfTk4UmTC22SplMrnJWwIRDQuuD
MpcqB+3k3211DRDtkywfvLFU3kzpnqfXU+AAVVeB83FdZspXtfcN2iy/hft68aPr
ExpBN8w631SAIBA5dsqGnTCvd5DzDxnWH+pL7FLjKEOsXQpvDwk8ztv9JSaDkEK3
sC0PLNT2gRM4DkXMsgW9dnRGt/NgeYrqcxyD1tVMSfGQi78EqkvQqc4Q77owISnZ
QYHSMrfubfaEStz4csAHhBS77UvleV798oYVcHkh0oK9NQItf7jDDs1N2jr4SxQ6
oApGCzzlhf25BXwSXgtlX0c9LVapxFkWQ8lZm/S2rw25Xh1osIZ6yk2QDKOLss3z
hO2sTA3Jp0REAwB2l4f94QHPb73JmmmXB2Gxf0KD+PolpvDVzU6IlBTwmYuz+2np
rj2kECzxb+3B7irH1I17BpOUOnu83dOoQphfiP1zzxeWOxP9Uzrtl9JAVExJ6ICN
dAJ0kINS9cgVfmpUEhyHzItNRL4F6PqcVcnImQP7a6KLZpsndFqtA8o9Y6/5nRcW
mnvFdCQVnDhUdw6PkULkSgo9Mdvve5Fnc4mzRdzOhCj8rgZuZZvcrBG9E6iKHmRh
VvCsyBzlOagFnobfUfukgRa81G3ncSDbTTy5HYs3/dGnJ527GpywvLSXFJslml1p
B3sx6DaSjneqbcs+zEweKWYk7/Em6rvCNaMtZ0nT0IAExhjV6h2NItDIpIRgAKqq
3wWQthicY1Gk5ltzVSleChv3hZL71CtSoKh2m8SOy7+Cs+Oww7edZPrg0HFTgl7a
sAJLJkM73LZPENw97ihiM9A94UtfYdBc5hCimZQZLCiH7GVcR3ULpyCDqfLxQmwF
YoBtnEzntHX2zjKgItM3X2eSyyA5UkEfsVAXLt5FlaJeA2DbJiGQwGmIRVFcpPPT
zPcFjqd8I7iKDtnzt9TvKMI240evSki9m3BDmQGPF7z6KWtbD5sp58OIK5FUll4B
ue+GDsjAH5mnINQOfYUNmC1y14kYgpHWSJTmwW6x05i7RV4cfx8VNm6wuM8cqr33
skd0P2CS00ZcZk15A9OiOK4IDXri59myWIK2m9Yui04khKxhwWs1WYwLI4DskBKs
6c2uCtF5qjYl7jRz4s5yYbjbwzAmvTiBvrugqp7GJ5Ga9EhWex4HIGPAWu/V802U
l9KFLSYMviXugDGq4i8te1dUnZ27hVwb7615bxlfe+LjAt2dXu7lR2rlPntuX1ZT
OtQ7qcLhrjLou0ky5GnHt1C8hI86V3u1wocJueMNeHJeFYITbp+J6A3KpG3GNgfc
1XOUACXp+CWs0QwbYZCUUj2C82rlGNQKRIBDWNmbDpc7sK7pMg5fXmvbTLaPKQWP
ZED9xwjJYxCJCZRxr/HgYKqYttKbmjZuQND7KJLQLnwphS/X2pDe3xJAcUBRyrbY
P4TzOiFRIu32qFzn17w/HJKTUcGgJgUvWFFgSaI8Oh2p3OJfTkSdYDsPh7v4NA/2
5T+940u9Sj18goORxGzCDw9Y2E3Oo6i47Zvu5jkEpG71XMVKSoy6IEdrlBacmuuT
QddR7+PfEFuDy6UNgs8S3MS0OXyURUhxH6nJ5+xKGJfhMCLVgJm316odb9Swi9PI
ct2ABaIZFzCx3pTKRu1beh9mljgW00Zl6gHYFXT3dw+gRLnE8n9jThBUzF1Cc763
0jMUCbkpuVIhhAp2kCjXWtXOFZPE4dfjIP9PpYcQ1a/I60brOzsWEtkeYcXkBN98
RKGHwMCvpEY4TYiB4VOwfMFRfNaVYlYZSbh7FgnBn1S6tHmOcbsAE6hiUMLH8+vw
aNom7mmma3DXdn7+k+zlX0wFYJxEHnHWWcW3TKikACeGuMhJTE7guAHT0fXSZTOI
0WsYvDKTucpVa38kL8XzkWalJI+l/m853iXcHa1rbRdN9wlZ9FrGxxx5rwd393IE
OCvWgUChc6ZBCpW3BVBYYwEnBM4Ojt9hv/EG1oumPssiJxxpOGZCD6yPZpP2NgWu
kSXkgOwmO9zlPFjIzd/HcU8Osog39DfXUo55VkALFbSHYTZCOL4Cfnay3KYEMyrC
ddOYtmjPjMGCNj8CYa/TRU22qe1pH0+hAIChk9OyURQ+Cc8qyaRolstnojzSIVcR
CDVbuCSgH/lCXJBwPZuwFwqSP7KNrSQC1AxwvsV7XbDKX0rCCH3tP10AJZRZQSra
evGJmdMMkuB64akeCaccujwpd6JfsSMl0nOl1BttSxRMXHfWfLGiR0t8SAgZR9LV
GTBpfT1P1dgCI462f2lpNHVyr+mIcW6SzxpABGMUw2sGuvgfOIGj7QoC5dMT70BK
AfNT/8+33COgRewLn12lxjKPxg/F0S5Mh3MxWkGr22bRXxCSo6sIT9kthZculwgK
xvXh+itKnr+YyczLmYX28CQ2pydQQ8rNU5ltlujfYGBCranVg8zKA6qMRkgihyrd
OmgTPotNH+sp7OlL5UyiJiE2JDgrCEHBybEgHZRqBgqaF9m3KPGVrUCYyYCyMxWZ
rms48xyBcvMoQpdRf0SQDJsiYBe3itMBAN7yfSAAPhrllA4dQUYDaqsWv51HDH/E
K/wvxbBw7ZGWET3Uvr3ymnWOpVfl/544KhGd6tmCBK00cgsrA/lxXo7GqfFvVabq
1MEBqvdSHC9xlGgzXxSOEYvZPaBd0ZBkhZjy2gXGSGEKr7+nUK0tkj4xeVA8Sr1k
5v+74gZVSAifeO0YwjfZQ9zycCbOBHVHVuVg5BCeRZxmZDiZMUpvJJ2TP8HDQauW
vYMrBS6hLd0uenhIbVjtrV9KjmsGiWwLmDXxMuGe2MsYbg8FamFvRpC9ULHBK5LX
KKmk+QvyyIKpYDyUuKyyP84f2RaweQ0dyMhQYKAX5luEVbD0g+M3yqvP29vbp4aM
wEAP/SFfHzse2qT3m/msRubx1W0oACFYch2SivVLPv/quPqnUg8J7/PCybbFez1n
YOENn2P5gxPw+LpdxLMhO0aAedb2lwcWiQ8x/LA5tOBizfLIhcEoDBMHS+xrkdLN
7Fc4DhfP0XGp30qmBx6tlS5nsYj3Wd9kTl1g0yX7WidG39O2aas2cBO3BPDKf5bs
3XRc2qwl57c8samTzMCXBoCio1XDKmuhnULp0ItQi3siPaIJ8dQZtwv9TUvl0In3
PP2P2J80p//Yssac7ZXhQ3z+6mgKpLvjcSP57+ftqGX8umf9REBAjjG30l50KASx
49fVE/JM8Qc5vdn6Bx6H2FqBrEzW/4jtksEbGNT/PNQjXVvETF6DPsBRfFpjwGtk
vzhlrGu5E8U3EVzYKvI3EfaQsadhA5Ttgldfn3OK6bZTrAmwYqnyv/znglg28JgG
Pbut/vNBo78v5HHdp7S4eCTMRjCFK5u/3J85H5LWjAEgxpuevbTIVNceVLUR7Kqj
TrBpcInlj9RSGKc2qlI0waqd7W9meh1/uh07AK6WkZu+Y2F/0JXTKSDDicGMyAJ7
PokemAxc1LiT8WELpJDD2tHpurFjyFAWlRKIcTEg1wcMsyn5+MXwuoiVakpynRb7
hiPP3TOId5yCuyIa94fo/svdkYWkSEReAqfkgm3v/5As5csxawGwBf01DYtI0hdu
dz5sFPZ1y3TkPM9tOWvqi+OWY4LgnOww640qO+GPwUypaBSgIMyqrqER+3uVcQGX
hC4QN++P3cs2Sd03IMz+0/TYCymabmmMRzqdmZCTubaTili8w3iq1ohY4se2l+sv
m5ZaHWb2qdrjqt8ihxfMtuHpfTx5JDAtiwdYb+BGEQj6N+CNIipl1rVkgVb2Qwnw
JA9uyZy6+0CE1EJStw9SoldjNhUv+VSjhn/8C4sWIf+4LpYZbsduGoPFPwutDRWr
aMk4HlE3/W91fXW3I4ADSR6LPRSGdplEqoVdwIWrOXRZIYLgaw0R26AJgoPSgSjk
4XB+1RbaikqdjZ88tgdqVBVk+B50DaofDCbwZZ/JpaNkjORe+TqBx5dMh6uUtWEc
Igp2goyd4J27o3BxKVDlYgC6TR7mmZ7F50N0urayEdJFm2jiCtso2PwoS+SAUUBB
PEjikDRhNuLKKH/OvE4SCHDo6o4hBQcHX88WfmdZKtSSJCjjnVoKynB8IuQI+4Go
+mv7lYcSfveqz+rbSaPy19xx6sohRdZ/haGuy74IGOEUINeM6QqrAv3wZH/dWH93
i2MNn6po498M2GpWTM+E+mFlNzt51nLaLMPnpgME/1mndA1AexnpNSYCDRFwCF+7
SiQpvf9YRfTjkopIye7/VTjIGuGriN/kIxvekeeC2AmXhx36HHbLkPOZIUwjwyEg
+oicA/lSBwKPdchln41qZbZoSJd7BupuhTzgStsZtRAWXEzE6hkhPTu6mmtW82A2
hREsLw+M3q1Nv3zhou/mTMNVfqNv/WjETbLMiXvH4E0I6TbLI6FWF7gRQtwycgx1
GIcV0r2JMU1DsJvG/uwURswxYWlJYKPLG1w+gu8Hmkg9y+UCcMNDxceJ7CJEI307
eQfj5kH5ClQNF8YCitDNxQyKHRgBeG0/KhWh3tvfUuM3cW3OfBOwsVEO/Hkq8OtF
3Jkl7skWf5NtFNfxQseQaoheYnvePON3HQ4UyZLe2kqZFefHXRShWTguqZxTPS0A
wK+cfYJOBJV3bRyq60nSdF0EpZLiDCW8yq1lN/JcDLyMu/+gYRhTZaXkorPsh57I
FnHivnlTzpQNzxh7hzWnTq/sAc1yqG2fV3SfkA1+GI0afwHMcTt/XQQbeTqAaAZC
VaJhqv8+7fK/WnUd7kdNoT0CWTjKyAG/OK8EzOSyI/JPnNdX94tYeDhvlfGdImci
DRErEWObB0C8oQ1pFkI+61t9aGYPSiV+twCOvjEOv43UzwLvemshGuTLqFSxXmIG
iwESLntXwB/ug0zNchDty1vv+RA41KvsQxjBd+PpGB240ofxV6viPgqMoYzecVRj
fmCnyon8MJ4f4Eg552feKmjlxVm516l5G+nk9hTRJgwNudQr2usGx4cKNYD6YXW+
XHexkkPpFUPTNCIrwhGcbGjfy6bfMi4Krldh5s6FcczI9lH1QVvoBmMXGpKPmhKn
H44JMtTn8N4Ywe4Q2LRCZKNw0EapY6be/aq99BPTfNjyqRO64WUUzq3XhzcK4MZB
L8SWN/2NIVN9mMoDrM/87fA0mvlvXH+jwk0fX6GZXhLzLQuduBxKXGghpPgBE5FC
IKQGRPHEoKtVMD2NHrpe970J29feyd96MYWtTNFZFil+YMbmHjUX/S25rTyGzw7m
vpYeKaO/URhV+cZFgthnNCBa1cSbdGAzR3+zrcBBOIStp5Onnj6B1r23X9AD49MK
2/A2K3yyV4JGXh7DZ+I69DSS5BYuZaMTaslx1uBsX+YqiHNtAT+xH9flHG7UBq3i
EY7T3TTrRWNRKTtSIf9rvY8POKT2DW+CRkMZLg8r9DeWw0+/xJe5IOpjo4iuUrD+
8OjBdDCCUfdN86Aj1tC27N2DRy9imebxRKxOdY/24zKnOPkFUvmvcz3XabhaZDDp
/Bb2Fqcrv7vTDQ3EWNeuOIYzcJILM+MRiD76Rck2QtZeLpPQPnCukZMvcB8ZyZVV
azPNXKYVVKJG0KQ7BZfmZL32Ph32T+vrfJ6A6wpvQDSH4yfs7HNJDQkt8I65oimK
xFB9JeL9Eh7dJozGLr/jsTCeCRGVVf2HrbGu6bL8zPuVKjNY9QCnV295ARzMPeJG
nAtPEz8rYO1XvUcB9RpRG+r4CHudYgAK1HWYpcXqvMb8VZt0MF5Eqhn5NE4tG9pn
UG7QlrExfatMucMBdYGJK+Eu8MDneRheewjrO6eS9r/gU3WI2PdtRPC04qxoHpoX
NFDm0t4zHqnyEKnSBTH+sE+SZa1Mp3q51YTAdT+6FTLF6sjB6AFkkcUjL4fXOJU9
n+HhaFOKnNpHwmNSCeAoBIUmSRAC1kAPCMO3DUqoNMfL+MseKSQfH5WqfMDDBB0r
Bgtyk7oDRFDU2NdqUzGrX1kSiOlL93E4c44gH1Zgl28wNRRSBxnlHTf9prc2XUrk
sPHGR8JjU27cNNR8FuGwTYp52J8VIg/iWDiUgVL641M/IZTTdJT1OLeebwxL+sAY
ZLtskrF13Qsz4nHyFN4BKLPydiCxnBMdxX12SfLeCHWPaOUlDz+WWaw1MM8Lpq9u
I4s2yNZbzlh4k689Sq/oKxuUCevY6NMc682RP32fGq4HBwptM1Gozted80cgHRbT
2wXrAOVd+icK50+TJzlb23f3XOu6CCX7jAI1ZvuHDJ28uHIOVMZisco2HoEdl77j
qmsTX+cfpJxaGV9a2Bc2nmRS9aMzj1LqWCaaPYjp95K3e0FPAMKwRj+smSKVEmn7
Zp3TMvWg3TiVsngm/XadHt1Xckki6wL+17esDvLOgLoobtHK8zBh4JavRPIaqXzC
ANjU8p9xl4jjrHZtzix6jWLHMuXgQ7nQK9hJUHGDtU3nqna82uFhJg/hBVlqt8Ut
qn0JOSPIrnKMs89VUIRpn6gqXIrE1qQpBp33Ih1cG1C5GzQHYHXrbToD6uBVAjuf
76s1bPd//rHlDdzD+aj9TBlRgmV8N+4FMZxibetHFADn+jHBQ39r8rSbHwOL+cm+
YGyI83zULYA+xEw33MIh35pIU1AJAZrDmxzfZh1PJwdl/ZCE4z8sUK+s0bSLUM4k
GXsKx3GxelaqBmGhCL+6dJL5Mv3zuYfy/+ZmOGFRBzJ+fIceRwdq9sBzKvs6nUvJ
YQIBci2mAMOy36izAniyTWGTe7vyMVsxAVw+9gvOykVyLiROUQ0am6mZALLR54KX
2SPj6jmDseinuwZjHnJll+FwpY8Muu0y6QHWy8iVnnhdS4Tx+xtIDC34cfDRY7rT
CGeti5hOeyb89/PqHLO6N2bbvqDw0X0tMUy8E1zwPXY9CFMUxDgQH/53X8+vlAn3
GGnzUux6Xo1LPagx6ZbbCyCvi4nd0NM8BCWnBQV3RnSjjtBh+Hz0DiV+A/V55N63
FHuFb+fVfaGZjjBJnCvHLelGf+h0vbTItOXvk/nONAS3IkD7hWFpY4NdHyC8p/vg
/cOQD8aBkisEnLA4C9rT5IYBcRkjbCxf6wGoYaMIbrppFBkld4sv4joD+lB5j56l
J7lrgQCaTOStJb32T7pyTKtbA8on/h7qOhOC0uC4JJr8aTHwgMth9TL7fHOo3pjv
0FJhCQAzdNmkJagAOGA2uPlDTeVCH2eKF8XSceqP178pRY8xDhaiYMqSpL5RqueN
HNo1FQtYqzf7Y2QLXJu1VZQEkjD7oiFoBiIGoHPXl0keXmpa3eL+4II2ZebtsQsC
nNkOj594bptScADQLp21x34QSzr2zgJlKVf8CQ71XhWY9hk0VwqRHbUSNikelyjC
0Q/8IB8VHBJZDr0v2wTmYuK0iDaK3nYYUshMR4cXuOUyYqR1Sx4CHOASPGLk1XDm
iztXmDrkJYw04JAEYFeBmOJu7yFrXcqe4FBtCsZMZ0HWPFR86Mbm97gaIM9iJA7E
KbdX1Lg7lKUGWGBNbUwy/cHSTevDYmwhNDlH2Yt700C6yYHa0IoQWiHNkO4NkIAW
MBabl+bZmQFhbTk6Delh9o27Z+Ynl8MXLmlyObzwSRkKH8jvhoxniZCwStvB8JeZ
xGH9v4fbNrwKiOVJg2fhE0HGcLpGHFpsIbA7duOYKoOcsBYlS9vyoW9yETG6LZbF
vWLEG+dy1njzJypgLf506dsxQA7p46oKj7mSlyL4Ay5pLSolIhL6/dixosDZyvjY
GQctJW4IXFuJIkKl1331GLKfUNDmwElM3E7gBrNFNS3Kr6kWkic/yUkL26Z7YgRp
5DxoOIVu7e7MYLMGXMOntzOJUEZMWcuZYxFZiKK+NMu6jtlQ+aJIP4bUXB2giADx
5JVkW6REgjed3VA/UZ3+imLAIbUbgMGVOt73y2igmLDGxKzsQdINuE9we4ttPiVp
jDMoptuQC6sJ3shkNNn23CVbT/WlO3hmFd7k78rX2vFXbZfAvoBsPBZ/ldtkv5xu
H9Kz/G51X0nHuYzatFbMeUE8en+EJdREnY3uGjKoI8K6SLOioB1Kr3PdYnYmXwe8
eDrhFiEcz7hHvJIOV64I14e322Roi9RcPFx7rmktdcuF6WWfWlOQyNVe90ErB2q5
m1j1YYUb+m+66VqTnetyOq++phaivjMKj3Z/KCsMkOvX7NKuOJx7aICVPAooaSNP
GPGpdf4sHXwTt7YnWVc0rAMd5iYU7ZUNBSjwkzlmnD+JpGlOUZ01AXa+zTJ5uvk1
voOr/N5PebSEWT+EJo3pvJ0KT0Ej2Yy6bEHElPSTVPYnfcUajr4lZW2UZtTw9/Wg
AJ4pCzvXDSV12sa34teKV1C0Vd2YXZFY7/zbezx++m5WKo07NzG9BCSRHuDX06hK
G8e11QqCpoFFKsi8rlYsl3aKUp7gms3KgwEPi7Rvcg6uXDgsXYLEkgzXGT7xGLct
0RD1QOB/+E0sLMnDXMISJI922DFDaCHbKvtmGs5eh+lgoJsiIKJwzGNyP2mPVRWz
/1/SG7R+xVfGv+vaGqfOCaJ2eT81tBHwgxrqjRZpzqkMbsm7TPSf+E2uzsJVUjXs
gVuIr9YmUpG+HrGlkWN0KkMEXgQw/qhQlhF4mLi03KDe5nAF7o0HnNo+HPG/Nhpo
z8amrYej3oG/qFB7k1bzCtduaevBet1Q4qBEJNtv/hF2V+6wTOq3nIBWoqRUrMJV
FqmHtbnlLNC1OiXmne5Wo3GqISjSyGuH1RcoT5u9iTVtpKW4mKUhFmGP1wm52Kv9
F56hIkovIH+jdTX198ocs0OQuZC6CZVy75Uo3Bov1l1AlJatRXWA24yKdkuV58Iv
Xe9kPAaWj1mO+JzCx3dFQlxm7YUuphmDknRZRGvm/z/Jmnw/rizM/jo34+d5oVdT
m/GVSzUzgvQl5Q9YVM3eWxkr+JbPfmf1k55RN2ofs1j38DFHxL8YauSyc4NrFdaW
1w/dv1mXYVLpJPYaaXjPxlvMmh1e0M6SR6qsSt7yltCbeHYYSEI60QwqJvw+kufk
Atrs6MQhowzF38K57qjcacCCMPKEd7c6tsUF6NsUj05UC0bZ0+1kbVwJCXqHG181
f5a5eHjH6Wr4PS+bOSdYgq2vHLC3bUXFJHfGFY9Rfymp2246hfS53UDvuZBOhcsu
pcnsHIRAae/XKE/+ML551/BVtn9+L6eeLQitrOficaKQ2l2n0cS7ho7ptE51uymZ
PCyaa5poRFquGROUI6gPUWVJp/XxHVW5cjEe4eE79CRXldsGmJJWYm3wtFNd3v3y
fXlK3GzH9CXfi1NqES7Zpfh59q1+06/ceTt+aznkiZnPMjPsSh3FDluZXuH3Xdp4
bCVwbd2aifINTEMxEhlBxzi5nUfXScS9d5vllwLZDjOgTM7ET/3QXnjhitwJibBp
CB71mR9sxzZ8QCanPWYx7GKoigo934SSK1IVuzpDwkYnmfnAR1C4xvRReCZsSpf1
k5xj9Y36nemVvhQ95JKgsYtAsYFvg1fqyL4CD5RlZNiije7fU6SPP9Y5llxJx+CS
Z/4Z7deisIlFkCXYll9flbx3YBczWyniSpsP0dkPyc5RQ59/yxlndHFWSwDPN0Wr
pCp6AVwtbmnjmroyrR5zatKUf0Og7KJi3eVuJbxz+hBkeH/s8uB8+SWyA/n9mgnq
yXqliu8SQjn6zd3CgOxjOw8q+oXNlvh7QilNoBj4JfKxE2xR5AzxCsNvq0aPBKVw
TquAzOVdUPASi7O2bbGl8SVytsF+kp/CfzWpe6rPJstG9JQCwCsgsBjToSsGrr0/
GFT63SN15xYjyiO9PdSi3IxLoK+XSzOpVepFL+y9K0feZrJOS/ysKJCJD7mY2lR2
k8t+9fW/4zvBi+y0o87yc3BOEMwAYk5bMeeO+2F0KJwGcoC5muchNBlQjLBAj0+d
l+Xt1TccpFllsEV07BNlgTP36AW1uD/wGR4r1u6pKvxFDSj5wnzISqZrcWSF/r9T
G7IuLuNoqhAgh5SBsyV9FyJODit9tGnH6+9eF3Nw/bTcYZVJWiagk4Q3i8QVTR2J
z9Wg9A+8idDenNDjeI12GYaNSetRpnFP6x5owC51BoGeEs8oVo/Bz6Cs9rWdABDb
t+p+2J/L+ilDTapqXc1ale/8aXRvuDlYM2IsOZexD1Zjd6nlL4H4vamEW4Z4uDy/
7NSbtFKxHMK/4T6qXzKHXVIbeq04d6tEj57udVXJqmtbnwwgDYUrzrkL4y6/4uCe
Dp3BXr73ijJ4+r/Pgxvpciu0lwNrxr/a5MOiNJpuR19KaBh5x/ehgKF0NG0vtaZN
FchbD3u3A726XuEdTpgKnhYbyzVnBglDHu8H7hiXG3ZIi0pKbtIX/EDJDwgzujqR
xtP12LzTGyZkob8hAgdc7XTtfP+pnBgLdgZ+83AYjcGFIStaUxt7Njyfr3ct02JW
zEDHw2GFR7Fj0/J9MNo3yNd6XfEdJmgoBgrqKN+EhKli8MfT3CwVMmYMD1LdUI/T
HgQB6n/9WaAP1b/UThxpe5v3JNCf1pHJnZQBwM5dKvD/VC6IldFSMHHWUSg6EaM1
Cmt2bPV9qHYg151+AVQ1Kj+x9kEFMcrQN+Y55xSYfVI9mBFT2te/IAYJ6JOWpxR9
Xhe8pKUaYtWeKBdWiWQ8x29YoT8UpOpXysTiqkE7Sp0VbLKrzyN4ez54eRNxNtdX
+gfCvdgTyTY5fk28gqG/+JZk2FJVdm1SMSDxeMi+uPYWLYKgz3ohbHq/p4Hbed/J
cYcj94JaBzf28T6kBXe7tnHpnMOgnHILMdK5/zsYE2XYnbC3kgvEkJaYHn0Sru0o
xyAvXlfC3tKM0J+r6K5EQJF7Nd7xBgt9mFvqgGEYIrl9L7A9/4jahT8L6/NnzpOe
4m+Ga2uNDLida5MG+YZLgwFbvjb0MBqwVUSBEP4RmCfVuZW61vG/GKYq7VRzaTbi
o5KPB8HckUhy3kCJt43wGrbNhubhaAFENqP2+ivn6ifuOUjEJPHA967/LV+UzF2v
2/ICJUIaqHh7MeHsWs6LvGPrP+mkO32TWdclNdjNlDpKYpyqciJYWTaYa59yR3tG
75HSpZaKLY6C4sOjZPsKo58bWXj53PRAFn60HdLbyrUdL7pWjk7wdQGUFLNgJ8ML
F86Oj88XrwsiTGsK/nHN/OGzI6iabXwbMWmkNq7xda/a7MQoPHFhaSpYJQ3JJ/Jo
TRqPtq0XLsEUVq875cVAofwoKe2u9+7bna7cu8099byDRtbNHEZ7xc0OCYnVBorf
UAWufNt4MqSm9pmw7exur1z8y7pWWXlCwxxK3pezv42I2Tyly7id9yX1ccbb/hDR
U+ylQml7CgcyPqUUkQ6G0pb0mvCcqOAYaZanL3mQJ58+DZycYAYor0fjpUOyrdV8
954cbBXx6eXEgEQ9+DD3OhbPoWWwv+bbGe3/TeWu8LbnQ0obNIWQbT+wFr+/WJSK
nam4Z9da93HKjQppc4nfelpQMogeukR1RLp+H2zKdPJkwgvwFUeo0nm4bQlKqXN0
uYou3TmONKvG6+Vt/hg0fP/ZoFt+jXxeLlkZKWATL1615iVlWvRL4ugPLjhwkebd
i27wnY9AxmFUiEVFPPSpWQlJD3SDAAssNUDHIuyTFwEDIWHZX3/u2+H9r37aK+kC
ST6BLieJKX/1IINjd7ZF/TBnDHUQCrkEfcIPvXYHxQN2xJXWqgutEguQ4xL4TeCx
RDMZAeiapKPT/RSwiJlQtgUSO1L/RTypvdzgbED0CSQKjN3RrQ3ndt7wx8HHFJlM
XKo300uhTeGPZm5kz7J+gqdo5xxQ3e6M+NDVEwkoQBWaeA/zzpZpiveJul4yCHUc
/PQE5hqHl17oVFfdABdV+Uizqm9jD1qEjlaGXZxuvy+cxnHOUFVvszj/daTnpmQD
2ZSriJbxizQ8LnnV1AzRXbF3wD6+7OHd1H70fuSmDjGHGFIVSzq1qLYLL/X2CQuC
oW3hA9Vr7uOUnUbI4/cnSSw+w45GucQU5e3S1eg8nHUleWAK/jJ9lzI3Dz0nazhy
MsmZGs9p46Sq4RYhE34mVPR4ocPJqT4dJ10OQAcBS4nQAGsS+AaHl4VKi0WCuXlK
SXDObTOiW9tITkGxDSWTRv0MrD5hCUT9W54FX23G0qCNe7VA9gX8hpuF/auBZqE0
v80zC5z/UaSqOa6HqzCU5VaP+vd4IFCJzj2Eyzd0RXUpiXAiPAfRDS5B8yGFXcg4
YoHK0Vi1dMKXnGQ0m1UCMnLELk9y6G+NuvKgPX5lyfRwezr9VCQ73VBDAm482azZ
us6lrVxUlM2ALnX/um9FE+7mrQkN5+V98VlB6wargPdNdvC72n8QoI+nQ42JyWBF
5j6C14gKLvoftBt92hqRGgJSCWfuUUQ3uYGGxWBxI+IUlJaGNUEkvpxIFZGYWVwp
7bSC1gSsxWn9Wab9g/NnE9UHxdKJW7uI2jCxNHW3FZX5H8AW2iZYFYuHj50OYT+z
3pgXp6+L/VrI31YkyjCestO8f5cvogFCbKEQhDZrw4PE7A5i/7Ju8w6yoKtxKkOQ
Vx/fOQjLh1NrptTFpr0/Rb0UjQbhwQy52DfOC55exiPoAEgpsx3OwUCEAGxiD/S0
oi9U9HkaXgqTsm430nD/40Oyn2pFpvGGvLcDGtUojMEeDRo+rC1nudsGK4w0vnyu
taRi0dvSmgkpri1g0fugvvpJ0D419qGt7uJeE6IoZUU8DSHr3lXRnau1xNjdGrQu
cwZaQMIx3qQd+YuXlk2MxK8EL8docJiTbwo6KCzpatZ9CCtP60a4YxaM6dFBo1wW
iZN78d2xh1Z2ClFcCrGBGOOxpYzrx/xndTmwCY9NwqWbpQeKu5N2Dtv5bPR2BHMM
NYaQ5me+zXTwR0+Q4PonvBKSyUJkHedxvj06XpJTbtW3GdBT7Vgdw34XGP+7yju1
uP3W1OFRTj4FuC3QMahbl9mzVyMY933FSO/guG1ge25GtLHYpQ926QxP3SKFfz7v
Fo3cwQaLij8p4VP+/Bx+aU32h2DcA5UhhPLCt9n7QFTKLQeXnk07UJ9LpOTxyUEO
xqTLk7X3wOaXrAU3nrlyEUOv/YDzPqeIDW7M6itC8+Q7mUi17ft35kX9ZSqGpEBh
Qce7DoHpkwF7jFGn64q8ry+lT2L2txMvZy6rHG27ukOgr1bK45CPzr/kAUns6n5E
9MKqBv7p9TSNvIW64M9QjuS5talVAGSz59Qu9R3HguCEKAOkf+xe37ViB/VqYBtE
auu9rd9IgbnZ0a508SA5yXZNeYoUfE7wahSSiKALp2HFsOeyc0H4sSReI4X3UfXF
0ylZZx6pSXUeB50RgXuJOgBf/o/enhJKn1vcqpvo7RfWcAaK9YNDpMlQGwLipMZ4
OfjH1tl2BiQuvyCzEvm/iqvWEWeh495rU9yu1SlM1FLvavYFWeUvdOULCi+FBgNv
sfyyvoBuS6+XmfD3TFMxk7daP7XObHLqLneKcVJF1B7E0DdJXt3dNvbH2PchcEMW
jJeu55bWvPRQa4HBClbLU04UZDmgWBv05D8EolqVSb00xkFkf6aLvlZhB2Pk40xl
DNwN17yd0Nf/jrz6FHqMRXE7Z+WGOOxvH93EmjhTqgmiR67s0+982dcBhyJ3xVQJ
pJfDF7XQ3fSocBXb9nkn17IiojQJFpnHcWQTFfsDHT1H6l2jgLQ7LtIG6YWGP34V
FufdQGSAGgodWcb3+e/GkOhf9EmZXCHjrgpQqnKcuoC8eCgE5nxOcTdSo0Poys6I
ad31Z4Jt8u8oXjDIJHtxdIr93jOwy60dX/nA2UXqBd+KkvSU/en90sSP9ZU+rfyT
UyaWyseLfL6PijYPmCgD5hHORzaijEOvPoCOMiEEWC7BHeCAZZ44Dz6Fvjir6UUz
8adrwKtN7ESH8lNlw3lPoAAbjwsH9dxJ/SB5Ys4okcit3rQuMP+DWKYX5LJ9KZXd
pXVxpe6NOyk3iSQFgH3Vb4ztnfpyDS2pYXOHbKbz9ff9HVLr+2TNPViH3pTM+T93
hSiQfYjiTZYvuoycUhi5dOuPtG1sVJh5LdSCHqjLrnRQaHcQBTeZKi1boub6mcxW
VFGSWHKDzAHlydM0gQfPNPccCyI5fLZKeGCfdT3oGS4mNeKdyhopFkQInFLIuyGz
RbFNZzH1iED1VKyxod7LbPePzzc+mclRYR3YPwD+FVPqkPufN8pIonW4eufzD4V/
04Jordz6gypJjctuGeYEtOpQblBEZz5gpq/z+joHYbG5YkNyX5iPLgTXHjFyqNvO
r+fbeQAHZUIfkne3+sAvz2pwcUQ7RG8nQl4+ek2IgxpbF2ThlCEkvoqHD9puyBmF
3E6Bqylw6qZxqcQQkNfS1qQtl9ouZ+UBBzsC8eS1gLNtbuG9ujkQgQwiSASDHlfb
CGMkq7Dis1Q7Wx6Jra6R3nkA5Omq3qa/aoGzzls+OoYaFzyiUH5Xpnb6fPNEPQXt
7WrxftChv1P6V7zg/MHxpYMifsOzzGn4YUl2iXlQ5ejzjYgrdWyqmUiR+4MGb8g3
0toQeQUmGE9B+nabFppfVFzlDy+iF6OiRILae/RHwA42efr720ZlBMOorjtpvq6S
X4QavZWG5imy4R8Vbs50cLkdegK5uURQbZpaC01LUcnOBW6spoyPFEI4/Kvc0yYc
yvp/sJoq3DpRrxXqV8xfy1NGKzyt3LpIfhYjlQcm6XapfZtKxoh1B/oyd08R468Q
qntN4Lg3xeMcW5iohZNj67ybuxIy/g/ddS3lt5D7j0IRMU+G1IRHt+xsX29K+2sp
AQzxK0l68Hikrs8WUyDGG58agF9NzbOWaFkB9OaP3NSoIv6HuuHkbjEQH2EPE4ui
X9XP9J3ukkW/hua9qkQa2iyOaYsD8eqNSgHNYRRFFBqueBxPdGdwhVYPkNuxwyry
oJlJPFIw1i3tf8Q5HfCI8yZf0l43MQj9RgaWeGswcFEq36+1URDm2i9PkGIh1ymA
qyK+wkdR507EAJ/fBpIyS/YYKOQpeuBXDlu1VwKtSf0yKRuNwlmkCMtlrjCC7fG9
rUZE58g8vv4HbCFaCCW1xSaNIRma9wr9Hkef9tVLOIerq3o1xaJK8d1zzfIdQ67l
KskiibkRKP89J73EUcARUlMNmD/3iVOyChkx/VCgl1ykzUPn9KiwY0P0DTbKgRUN
vsrZ79OW1DZFD3Rf6uILyLeS5nOPc+llAjObBacvCzxpoS1cpoF9LX3+5q5aZpoa
MmrKWfpSYotQ1pL1k7IUG2JfqPSEcFOKpdueT9DZBz66OmB1sE2E5bUoZwEWcf3d
6recmtnXHHUGeR0LfCFVpH3ewD1rA7OpI/FSBBOZ3+E1i7bDX6gob/yZdWr+a8FZ
hIrHC2qVQVozkykFgPCu6W1WEaZjGhFdwHSLrsY/hv5XYQ6o0ZTYxlsGkhP+s+RH
IfeUakJqUHCIMYD+JDeGqFS6v9TmBMzMA90nvFLM3f4AEh2a45Ih2jFV6dz330P+
Ra92q1OC+KL4pxtA7y1OVGCTFfC7lOtEYjQZWB88rzTpFF93pYyht044jLUQIoUa
iGpWJIGvMPn5Qe/IZ9RUDjxJkdCwpEWuhTopw244taAMyvprUvv4YToAtUKVHtXR
bD+rWRhcxHeJp0AtzX8zzuY57n7rNAWI7GsOZfrZ+jm3NHKH+g9qfP8dTcjjlkYj
o49skJMzxdnkSXEhQbKQnFWAs0vbeYLCI+QPVr2AKdHrX87yF111r2fdOCQrb+6h
lFtOUht0qK9gsvlvyeOOfwTMZ9Tr8RrfsR9UMwohpn5b3MQwL8BbLjDeuRSp5gpT
U1Gcjmx+Agxcjlnm3E+rgwYl+6ly7r5jhoYMOSdqqMXpkbKQ7KZiDuBzmJt0ZsEd
oILfd67ae9JYykZxkvQ9pkm4VHz1WMDUwuPeVr90x9L3ytD4uiPu/uXi5Ox90aFU
ur5dEn5GbZZ6nX0sEnTfAiUdioZae0zbmtweA2rjOyskuN4jVGbXUOyJycNPYrLP
YgJcq184cRtoLmqbst6L+Nwn1s2hdkHb/uxYHReErLQJkjUT85gm56rdM3Uez0dR
w+CcYtkiyAxgqdm2wfTdAGcQBXzJrurGn72nU9Uit2VpHkTY+SB1ANNDvy4aidcm
PR9AdEGWCckp5GHDuP4w7FVOdtahksD9nu2TMkxuYxzKIp4HLvDvqWBFMEv/rFuu
BX7xndjWwN4tfSUDifJ+0y95/Cw8zWlfqsQdSoRj56B7bRfOmWBzH95DxHTR3STx
VOF0uv3glJXzgIOIn1VD05G1QtkPIKlneqNmDXC5XfWBmoT2kqUsuAbLQ9yFYl8y
N3SJI7MpA4OnaDyg1F1Vb5bPiintpg0L4DgCfiD65NlKEK5jJh++fTaCwRrg2Q/C
syM+T6TdaSzfo98zpSKzYiVux08bXLATCABjOP0NDehfTJ/NeYGsL4J1QijUDYgx
a2MavBjchUbj2BXXv5wy5vuiyRDGhPOI6U5uKize34yt8YWj+Y6QtesCzlLEKuZB
JFmN26nyoEpHdzaN0dIhOoEy66qUi03dbBNsNqiawFCQWrZKxfuafFBdCTGHpVyO
+PtPA/DNpoF+CjzHenkz9PLXjhHdbM5tZpN+fcFIruu+k8VhCO0vDfKjMtS5612w
TEaUzTPjEkKFL08j2h/U9ePhnDAaH5x48sNyygOO/2BkAR1D/8Uy6yrhZBdOGoEH
k5MlE2dwRCpqdNb3sJc47ZNyGQzbhQv/P8UsdV9zro137XO1QHoVRRsLKz3HRNQk
STeuoyqU72aicm4f+Qsn/WOB1afSspZ4uIIq+T6911DAsDRG6C1JjzhV/0VZIRng
EIecTx+VevgbsfDRvSPgNA0MCQTT2WIH3yd/TNYn6mrvcq+ZKsFef0x48cyR9Eek
povGoyko9/Du50ev7zLtdAJbqwe4e8qZz9naM6t6erh5IZgeS1IJrzKmjKd3GktE
mQamWOmabYIR02Bs97t5bZPm0juIFsqIixrZovVnxhKu3gLm0TxP+dT5ec6D3cHX
2xI4q2wC+wB/rb2S24KjUTEai47bYGvyCqjHFW9DYTpUIUqqHLHWh6yj6LhvelHn
ZE7s9OO8aj8mi4QJfOTT1p2BaVX6PRPQ3lRoVhbWxr8j2f8mg2WO1YlJjanfDCwD
A6N+/Dq8Pqu2ZGk5UR6vNeZH2gPBgfkw70B0rIot67U4QcdJXwWdBruK9ABmdPUj
38aCuU/4bq94sp8JeP9bWXoh5BIF4cHhtn8CV62S/dS/gaiAHLpKFUfO/c4t+fkq
gyfVOTa8WqmIeVPmlQUWqXh1G6RpCf0FY6H18sBhcGB6OvZ9BGcF05JDafUb4Q1A
6sV3x///yNckYOWClfUDsasnD8bRjSE3+Jl9EjVja9HL6wa73578vrlDQK6ET0PX
jUHqO90W5qnWWxYeURNbdvht3FDYnfDkHvEq+BbuGMumkj/L73wZAWTr2Uw3eHDI
slCZ0V1cOCNVUeIrOTLbJkNNgcxNssThnaP7Y0uahrXNVDamtzL3GTM6KubF9g4W
Wsasy//PsZgsYcqdh9SliR2uDc/btHetaSQ7Th0vE/n5ub+NsTDifZwqCF/q2iei
fyjv7UgbChW1HU3K3YJh4W2mDbhUdUMc0/xS/bKd46Gnv0Mtc4Akm+XyfYX3RgYN
JKCgU0PcB1183XjUIo37ATZc213TQWUzdbOumyCtGH1tr+Grse+/9Bym+IszbeMH
NqWSZdjTR6iaxdl3WbZo+BzOTU0oPMyn7hEM021x36PFV/f33BHgSrrpqcgLrXKn
S9Ji13ZCXgvO4e4Ano4bHTObWzlAuIvY0Qc2iuYqEymxx/FOXOZE9ZkAAmrRFcjG
+4OX+SgEEqSYwH22DAIjhPhxABou6AzS2hE3bOrm0YrJyMuVOlkk5JhuZxtamiGL
9jUJW/sIDBcDII+H5uyF+XoaBo8uszCZ+CyUh8SWPIARp0YZmGYtXBzSwz41OnKj
swvhFWMhCQpew8UAEDdAimWsWJz4d2CkqdibAljzHpvJI7ejOggR+hS560bgFNyH
O4IYMWbphhca1a1sFT5rAAp+pXBOU/k/wbowVBq9nANo/rrtXY43rjR7nNTKxRnN
WeFrN/nYqdRiLquaBNt316A/F3O941esEvhO1vLw6d9oyRBIldM3zebi907f6gEm
k4LC5IdGDCKQ7mCOGCbPEs7INCK7/vWAwTjhQuGoqZw1Aw8C8uMrcCR2d+790YWh
JXNu+euulWTKfAgsvwGLP3r5xtkQWPzP/bC8oRx66m6fbIhA8BW2DQ9pT5XkSyak
oCtHhDIkstgrxbEn8zf/F/m+rA4CX1TDam1WKE6S9q7SoEyuve0s4FhvxwsUEb0J
JbsN6uArLrGtkGkKlYUSlKzRtCitSjRFnthbAmcrEr/Dgpu4iEQyAPPfWPgT88sg
W12VXrmtPEs9jaIP00+iOqllp/L/fAyg4mPpXS4ph+mnvZznvI1H/O1hjbL6uRqs
dJ49LHnpyAtHG2FNHQNx0HIUt3vhcAFiDme4KULdLGnIUYAECzRIuuIiW9CAc+R4
fQsv7Uyje9S2ZWQ1AvMLlhwcomiFsGR7HeBd6r2J1jAYzeuRWqHOlE6tQEaJ0Qtw
Tj0qIOs73LfuPlwJGlMlAbIfiN03WDIzxBxhk34x2CDxIb+oxMrB7hp0Eu3I2QlD
AdqY7IGHLgsHCeP4k2WLoSuRD17c61ZtcwQAUoXNsmwGI8jYTWYCzOn41FezchXt
GuFAEaQwjbMKh6eC+xcgbr8Zz8aQ7mq6dtreugpKOP8fIt6P8RZhQaiKl5VblOXO
GiNw350CqDnPqReaosHyVT5IOKLU3u3js5PWZMf0aiii19hk+A7fuKpkPfdTIDBM
jJP1ujq4GiqRTR31O8EKalLbiIEcqXYgt+BKa+N7R6y42OG3qbhBSAmHEIJG+H+d
ATrw9RWid9w5I3ax90h8MAAduakNjNEhywkZirM3ydDKKx8jjswGv/eAdX4aL8KN
hWrdamAH6s9nyVfpMnkO3QX50svhuIPll4sl85vSElTFKC6rJLwY6qs6QG0+PKFu
sLQGNlglUhq/qF8aZfEQ8ufDKfL9oSEyw8uxOHt8bDZ2NycBokD41YV6xxUL1tVE
5nCyk6RyBcoR1sAhUVbPswMoQs4MaoEChkLGfmMn3siwBWM9D0biiTI4WK5vZtnD
Tktw61EcRh7ZqTmJpDFjXQ5wSe27Dp2q6gcXkOLc+AdkND4hyWR+zsGDgJPUloo0
zo8KUxK2HIly44sAdNG6tJ5pwYiFMKWr6yPEr3gYPJv85LRJbh+Di1/0+157ewaL
lZyHDG6JIhhM4tDhNA+P7iCipg944EIMKPGnvazTZCiYExOaQP4oGiJfyApQ2x0m
cKqEbpLBitKDUKquHSQ5J3Z7aFZfi6JaHgEGYdAJ66BQa1yGsXRUEZRxqgEz+CVo
19MIC30QSn2kZkabzUnlBTb8gRP80rOrymvkUmtgr+nk72BESHuprTcANmit993p
nxUlEKDatsVJRxArvRXQQX2BeOKzs5xQRi50+CiigiRJsqKlMaJVlZGbkmPM8jfK
KTQLrgOFgGYstyvsSJAThLOsNH8MTyMU4OZSIa7fwnI2IxVe1wXLcLCZM+mokXVI
K6lQSdvkvV9LiwtCXecq7pYExqspz/qhYsNKesnVFVAZSSV056leVAUT145eor01
yZYbaJ5kfPWhERWuEWaCn6iyYx0b4ocCWL7CJdc0eAaE2CAbPzm+jSOrWose+7FL
hpyZv+PfnbYSFwMjaqQf4FaPOjhJsKOr9WMx+rVGXEWr+YlQUCq/Kq2AOq2DVAQ/
wWi3IphktbFUp1Ah5ipVG2amM/PBouQRCSLidpsd2h/gcZ2gVn6TfUn8VaIQn5hT
0I2yeQ9N38KALcwNngxvsJyvuvBWKu/RmdbNKFmKiSXjllMmwrS41WK2ch1U2BdT
i8SGklSEy0F1wQdF0qlm6d6ItkZfx7r88fpRzxtpdOZREPgcitf4q1+EB9PomdiQ
DG8yyKVYc8ZChCM7oWGMcXMC6qfFdtQ7qpST1UYyvlDGl2iqs4046PtLNqXOja36
+gYbjkpGwWEXxNBIEp8/9qxEdiINoWCogVz36mH8bpMlWmYI4Xlq00jgm3OBVXrp
YbG40U4VVZCVSX3gtj7f+avT13Bu5uLjpt/ASR6SQrFbC2PUZcjAiO0jzKcSpWc/
UToXC5FlVMGxnaG4UTlC1zcnDPii9n0wUteKU2wlcGcJaAzo2AdNFRlErAwZ68Bn
HSHiUKhSEzFyGmWlj4QTYjG0rMS/AaiOfgwmgRuqCovHhha9JYC3ueYGAZF6qU2y
tmYZJR4Omfk471/IFwIuX8owt1z5VBLVfIq5Exloces4YmTaoebAkhc+YVQ35t2p
Vey9pibH9eEmLzpNE6KO/3M9tEhvP+lbY2oHhz38uGNdHo9H5h9VJJwgciZ4k0fN
pYsn3UgNnr8hypinTQ2a0ClTHlSDAGXS26k9/tjxO4rGYti3D9eS+ma7j+l7NPsz
+l8fiF3JlotCscUZwLGgaK/mYuy55JkFiHqUqSZ2dKnhXvHprICcbOACEJRmjJvI
yaQe6P9qn2A2zIdNKYRwISqPlfpQoDOenSmS17I9YXLhi21BUDnHlyB2cuI3BIdY
0cUFY9xJRtHJvWszEK5sO4OHWycbOnNCRIOMUZk558UF8f/5kKhWyo5yhUdJLrSk
r6T2iPfWASuPsNrGV4Y8Bg1q+ltas3T6MmeUHJykdNIHrcwsKuaX9gm09lKYzocy
0vpwqBwide/ASXxPEkzezickM3HmxLgxCKHyaP/XAe1sMCr1og2inbIq0FHgO7jj
+v6/OEaETv/Ny8AjtRCDS0wbOupoIXsy4SofVxV0vGk3BK7GQtVjZAz4JGJPqho9
TI6RxBqBDn/TlnIDk3ANSlNoxpRHPH5W8x8h2PXvAW5sYWuq62CB3tHLSi53SpCj
1Ebxmbw03VBDkGFS/kh3iMtyAW/ya5Jt0lz1ZiMKuldg98cXchEmNnyzfu5pNt27
ptUSNGeG4gzJGxCZkVpwujsnjwqIIHAt0eyRUDSz3+GDHgBpjiGtKnC9yXdXONPo
10Jmw+X1eJA0/3Pe9djq8OZg2CYPL/RiiWsLWN4DQMaTsuGFboSWHqxW+071OjDw
tKOYhL859JjGB5SNXP/7Yh8tTmFupuqC658MiXnRgXbn7ym8CT/HwjDd4Yi6clld
w+4BWHYUSsTxfLVWt5sqbEPt96A06O7CBct5hs9ZxF6xB07nLu2UlZXksMjcpt2/
NgwwdU++HCvHqF5AFHZoShz/nbie13DOBDa6DEruCSwPLJyFANN7k11Ijm5zKJDy
cWIHPMKln4aH8T5ubNMOlharuGwcaoEZZgtVAeF0PAawborQkfOweAg69UIbl2Df
9c60+juCjsTxEEJFIUqRVsiEcS69UTr7efaMLKfvL0lJsHpg6IW1ZBdDWXwBE1Oh
78tzN9y/aXUuHXH38i5eYAgVgOA/Xl8R5wV8kv65mmZCESTafuJm0GF1CwEvlmGT
wGI0bVtESTFRUeuYWk9Kdn6x0P7OHMONISf5tKbcBQXs9JqVUge4MCSAO/X8zu9t
j/ghd5B8vIC/3yjCBCxQMuvOBNZyLeNexXwmMOi+N/Ewsv6cT5Cot91kGeKQ4D3W
70Px3+Gn5gUN+7BlhJJl1RvIynubONDsCumg8u+0OkwFKdGcYJ4A0W5bV5TK0BrT
CEqVQO5ZgWiMmF10RGkHKD3QfNOeqIXwvfdf0ywEvvpJGLyqi5RA5l/1Gz30hV/T
26h3VZMe+RPPI/rZrZFJCZctkcWsw7srxfdA82an9LSgHkIPPR+MtphKKuCmH3yO
tWNZweihh9CuTWiQYXChJLcgrtXhCRaSCw2EiubOuVqepK7JNOa/GEv5T981V8xH
J3nDRs4pvn+xt2GYCMBRP2PKLajyv3ALt22qB3i9T05wgqhzvamf4pxYp8dF6en8
Id212vxb1/9vSSF0Kug03/bSGr3UvOaXPZpKCJ+rOEBz1Aex7DUHWL/ilsF7fXv2
jvcOeoM4R5ijEY5HMFVZGYXhWR73lAa28NQaxI6+pU5IgJovifwijlTHRt6qFkC1
Rdj5yrbgqii9wFL6zgwU1ne5Gflx3Xc81GbHjdo2+MQdvVmnSZQCytQHUIZy5JyK
cNre8EA2degJrrFxwo1z5T0yWDux4wvlVTptkHngl/1QnCzvMszmmmo6D7S6h1Zg
ldxnwHqIjj5tveoI45Ankcih3BlXfd6QSZYOxYsyiqwrkJpr7lxfaeOZInSQOX0S
lhN83EpjFbaWwbU6To7ZwDsw68OQG6ML/1JzmK29ALhmCNpiWtdWaQG8N+k4bexc
mYuqQqTG5lGwCsDc2/Tp4L+NkvjU51NF9kbVJ+5n7wlfDeYheWfgFqH/kNlX9KfS
dqPGz8zXcsxtBEnJKVqHYSn6aJjsfmS0XnMbwOneGBUmOK5IsevpuQEUea9htAyb
P5M1a6GBJTcoe1BCbNQ3v0EJlZSTMX7iMs5fvn6ijxH7+16gitIBVTwFVK8gHXvh
ldnCWQMzIIlHW5+/20rQkYTRALh9qe5OHkGUiCN8LsqIx64CL2Q8YmJdOQUIpxSP
nOuAZHPl0z4SbxioARpJvLN04GuOiw3YgcYo18nMcPPeVBYHMv6UEFuCIXv9i7n5
a6k6bbA8/45eHh+4CdEyyDstp3IiS0Ub+LyT8A+Np+6XRYxMDJfHpBpZrjeKonki
khFgyG9SyMstUVVOylmD9w1m8KjQwiY33i6eon87awM3NjbkN5yphr9iYuziQzGh
DErNQPeRH44ZzTp6dAiFyu1hfcjFDKvoW5L7UiDmwaMMVlp7XYUBp6WE4a6adoDx
tZnYjjptbRmV8FkVeDgq1ugGVFF84N5/vXAuUePsN+0BrZtRLG1+xbQzs4BouIsN
R011LYlEu1tePj5X7G9ob9uXInoEusgF8BbBDJMGgp7UVSno7LZTsX+LCX2EB0uN
XPDDvkgLkS9kDnsPXw69h3mhZ9QJOwDiowYmtRofRZyECzCyq/Y6x0tLEABgs9dx
WGPG289lACmYTYVbZ1Ga8u2efudZPJJJ4bWfsRXc3ToWo3MXW3XZnmRkOLGSXD9d
9nCzojxTII2jk8+oq2r99mgqLnOJKkNSeJw7KDNcQ73muNJredMsPHZFVrIoVikM
5wHdxjQRuGbZuY3qUSRPSYFibWABgBoIOcAPi8cShdzxm10CEzYk6EYsOB3EF6Sp
x1cbhbekDGM0bnOCZpDHZgDnz7bm+EbvakaYK7ScAXYJe6t0zTHrgLM5Vuvkuo7d
ATLlqJapXpQfYOxEE65n0opDYQwkbwOQ9IpV6Ta05xvqkeGmADrWSqK7pAFh4sOF
j+Yg4ayhq5RRD3vjUHZqpbViGrR6zTCB7AaI8ZNAyDAWHn70vO6RX4h8bK2upCU4
EvwNeX0gqjdbhTmY3dRrIqhYgaoGeLcYO9J+BH+10lBhOguDskLY6lQWFG0p6pqK
sZBI/Q1wMMe1LLx9qneRefEQnfTyN7Yg4u8hKU54GDa2Uqje0DZlxK9hC3GaZZVE
Ieat3or979gsW3/C47G1g9ssEaW5G9/+Rn7xZPyq5SPq8hwwk2rYHDY9638gWGsu
Y23yCMUE6OWtKLkZzoVpF8IBLsueupdYTKYh98qUp0Y7fc3qXOsV9sySAGFJVzU5
aO3rnr/LCxQvAA/Efyq7uDJaUvT2JzMIILYT+tMT9FiCMADns0itCcPdS3g9kq7q
U4DAqenrOZl/XBRjVPWOqb8V6WDw1qhOgB05rltWNPWtGbPSj6KlA+G5osgpII7t
EDgflrn2tUfqUXVzOqkJjUP99JYtMJL4397uYp1bNZuTqFED/Z1rvA/0St/UQDyH
m6c9s5AEVEy1ArJdVMh9kNmMsxxutEeUhTqGARsABsmJYR+PRUZmoCgCdYzZZ35p
puNMSx91vlvVeRSaj8T4bY3wH7ikN+I3sb7CkmceQDlNYYrfj2AjghcidkMsZ1FJ
0kL09yG/pQnXuE023fed053HYFnT2fC3ZO9UlS8h+Snv0stpSvfK+erscLDHZSDo
V2fwG7SPlz9D0TGHQwhJtMEprfL0x4UCFgc0HECiihbA4026Uzon1qNNJdLGdyZ3
u7iLjK0ggN4pOwawtO9pGBGkGfqS51lVgoUAOH+wN7GB/5rOX2nwavwrRWXFzVgs
UPzeE0UVpdD9vcn70kNrciOkeQHZ4dJmFR5/s/WOmyolOB+vmdE51OFcKoVTF6Fc
Wttmdtrg++a+jPjlIQQRNQgksgADJVJaD8pAVNKAsp4+6pfVc8cGiwUeMg2Jo99l
5MCgypg1R59HwHrm+BRuql2GCjud93VDWG3Io1dsoryQDgXLQl99nTnF0XSIBoGt
/prNtEkc3OCLPQEzO4HkIjb5LeHfkXTMO1qhIcQMmvEQavWSRTrilF7VCLdFNq4m
1daBaMMhpgLKF+s/VQ4PZMEFGwXQ5GyLy7Ev4Wq2IV0ZC64BUMPfO12GklBBHH0X
F0jMQ8aW0n+NIXdRLWzEI16yZ/bTzZhP3VuhfIo8zgQMXalTLp+/ljlIL9/+j7mY
ikx8yTby4tS9zOaq3wsw31IYX/5lbrbRs6vgur0daCu9Zg1O/7kM8jyDqMLGprhH
SeQmF/S/4N44CDhf4iGFpWDCGyCiehygQNpe7MrHRimDfRJL34iIal/nMeVD9oQs
npYdYBvWOvatAMjFmk/qLVyvcTchdsmW9ddGP1P8NtQVh6HA3TxtH78whh9t10Y/
PLWfjs1ATiwFcbRJ7Y601RNtBA8mRQ7WZHCnvreWJ0tqlIzVelIXqgmh6YglX6Gn
KAY9bBjvgNcuP04UlKRKMauRXlzrOcOLivajRq/zCZa2knwggkN7U92wGHZ7aVKd
K0uM//uwKP6YaPRvxDl9XowtW57LNi4Rc3dGM1Kh1ZsWHtezNE+Q4iGS+ud8felX
CbRkF43cpVDbEw+F6oedoF1jvcg++maUfaAl3wEzlTcCONnJZN8HowHxkEECQzcn
X7dx6WABL7a8j7kq6nmVSPY+9cGtY3q2A8G3TM/gguYVEK9gBGYdV1s4Yef/TQPT
zj0Sw6mKda2tHB9XX22u1Kf8UWVOh4WbG3c7Z2xG0M7c0R+PM/aUR4See7nGYCKF
lKiHZCvRwn/Bmt+YGjTHHV+pX8ek8GZiIFCY4ZovuTDLwExCy+Aq5s48jhR0qrBC
KR5B6gyYAj0bhh4IOqBlHydWt7OeJ9BqbFFvdulXk/TpTYS+zRtC1qZlhNhYU1TT
Ts966/ZRSIZV1sfVjAyxAp2/xH/wEiNaxfIKGE1vDJjw34Qnw6iU+y2C8DNhKBH+
uh3r/qYMiCO7HB/BOzgdRRsqgZGMf6IEWXy1p1OW4QsJJcN3SMW3aSadCNSUgiG0
cSGXH3acFtSHFXlzekI/6zJlJYbIhx+t+yL3XLMf65YJ/lRGWwBPGNxsVdKdEkjw
KZEAiNxIHzFuCvXhLqNm0c98qPdPHitRI7GqTfZYDVvcMMs6cIKB977iTUSW+C67
Unn964l02gis/Pf65R8MjdrrZ6JmOJxcVq42cNGcQsB6pOUgYr8Qy5cCzdmwqqCa
AxZ/yL6099o3odnfsaOXcbHaSXIsS2Fnkc8d8Ce4MJiBGSXYoQroCEzsOaR3aac1
HD3UUDotQCvwtDRvQKTt/QdaR7QeIQJ5+zNKfawCpMxShDmKto9I7jo9vSTJV5cT
jFGFgBY5s9dZ3fXGx2KdlYD/SolXt3qPlNJC+gWOJeJ8UiqFWX4OUlIadFQJ8R5y
eHNtuA67A3T9RzCDW/u6KVkVAyfMZuZVdtmhofdvNP8QPU6TmlMzpz5cYaVCv1b0
8y1P3NeQk5XZ2NQqOeMzvx5xPvi1CvVVuWtbrWkiz8MlTGSp4xbLGlScDs7t5vxS
25FTytZ59KILm4WWtAWLMxp7R8tQR1s7gwu3CFwVubJwYk7mhwmDrXSitYrWD0FM
AtbL5slPcty0ZorhWgdQ/T6gNhQER4x+MV9Bh7ZatRVZd1152OUdip0Qq7lv40aO
Aed5WwkIS/iktDi0Mb6r0QIon8/tQD3uoPyEUvCI28VoCfd9qmv5AmNCo99/qCn+
QeH8/OZr0nPN/Zx9+Xp2MDyvs1GYMuM+uadyZV+FWOf9Tz2H/cP9bcJHnIeEcqn5
ugtwLFYT9JfQI3zcpB1/9vjw0SJElnMZr4mjwtGHlvPaiY12ErhVQpJ42UvfHWWp
01/9hmqP57cRfe9XjFf11PKLcGSrWQhENNrh3Rjw3U7nVCEG/OBby/D8N5qqSu9I
A5aRnRh8g/UHm16+JCgBxu0N0B0CF9EJAr6VMwTynyCGCWYWyB+4DdeBUPkRGnUn
Do5fA/T5dMdsHoYaOaCScmed8rdaQ4OJhq2PQcAZyXp/r0wm7y1PJKxKm7Tt7RzR
bTDehEMPCQgCFMNZXe54L5hqpQG9+Bs35AMRii+VnsfHRwtJ5s8YobHj/iLi44cr
Y4yGO3mGU6MItyvJq0PSNH/GM9yGUF3AFhcsOr3aiX89l58+/wvQRWobSzMEZkwi
UX0JZz08QUqWT84Bm4o6DKSBQ/H8UXyWj8ayeSPQ5YMWAWGhJKMN5ujyRy/XnYmG
lJ5sb/k+sh7nMaZEFP7FfPEsuC402EwzH/kP7G8MTXL2KLUu8BEnLTfk7vfCfOFh
RpEwbBu8bd/NcTFGh51pWNdyYkJ6GbL1Kw5JeuiBp3mqUHsZLLLccWSxBUchC4E3
LhXIrD1J9WbWQuQw9l/rArBubSC10FSlo3qTvW0JyNuP8mi5Pzw1Nk15ykz4i0mZ
b8maqJKX9I+vO/PFr+q9IHq8qeAoeJ7c50YGHGpPwVwqadWOk80/4Xt8ipaHzhCV
u73gzPyFBM6Z1tmlZhYk8acwLGSmV37sCS7jOLdiYfxiywMria9dVuSQIeLVzDUR
GWJ96o8jrJb8DNbJ3/yMrYCT0k3AtYXFf+5Kp2nSnRlInRCKTMsSgF5y1o6Jam28
eXMkPmZQBdi+ZSj2PZzE2219DeXD4h8VqXughV4XCM33Dk7XETXWfBhJcLs2RqA8
XUu34OnvnHo+wL4mZ8RBufnSYwdZQ3O6RRFY6JWLDGiGdZnjGI8GohnwlNp1WHS3
t34Kn1C49B42mMgXrB6/LW9LkmuREWGkYh9YFvltj2R2eugIVJLdHI3r6OQEz/ih
N7DiyKFaM+cPaUl4/VfOVgAoqJrezoTxZ6adFVLXNENLrQsd1+ufH1rp+jd83x45
HkKGOSNESCJ+k7MJ0QOrMuONGKIyyN3zW//zkDLPS0w0rkoerDqlPfNmvqVUaaVz
pwgtXSTDyOnyljTRGuzgsdzA3WA4sF0irZ1nn5qh5UB6/baCdXVLOKI6pAE4N3I6
7b224CKjxPlY/+OTO1F6GdwJ7koRqY/k0o8VWefMhE8Yp752WOd4h0U9GC6k0KDH
gy4n4YR1CfIpNcgkq18sEmOLtWLQSYdxLiYfVaofE5v9QigZXGSkDqu5oR9MJXa6
jIzHxvI43VPng8Jxj+/PTwP0GhC5ae01DsuHmkAWwIpfe6iZt3oFx3lrTOp0EAG7
ItiIaViWbqDMG0KTtb1DUW7oA5fukeFdOWQHpTBHKLNSwhXSG2VtbHfIve/HB/No
p0nw6Bob4ZBlsF77pdCL5JFuTkNljv1N54wt+MYOewL/DOSNazXv0RP//4c89Dtf
ZZ8ohjbv01OJjN20NZSq6L46SayhlfEBG8j7s71AHqOqbeOGiRBaw+nRFuusvwCu
yE6uWdXBasFmaxnSu9dHYo/tHzVUXKgRJIMgi2N1ubFDRjB56kEsd8mv+OQnXGw0
LmYjk62zhFjuS9YggcwLN5VrLcSWEaKjoNaeS2E4aCpRa1TP84ElQJ+m2MWqk2tz
w2nHa9DshI8l4Cy5eIVHetkWFqfdsXVIYZzFasSfrV4ej1gHNL1PK9xPDv8HbG0s
dyCOLW0pDggBSWjhn/5lDAT1S5xTHASQUegErtRP+Jy4DCg57Vluu2q24pEp/q5J
QZ1NS8fRVWSMOD3JnWgD6w0MwXjqzptwl147Tm31mGr1ELE072hd16is1ygQWNGO
4VaFpYRRdZCi47ix5hVpM13p+50CFdQfdAqe2FcmPBuBT7sju6PVcBoIOtMISPw7
dkb7J5fOTWLiAjFWRKePBSMBS5PUfikpgE/kWrn9C3wmx8mIEgG4EpZ0I3g9ubE3
DT5zMCG6LojjQshUD/hZv4JW8xP66xM6NN/cHQAMgxuU2daEAd6UcuH4HFma7UgV
Zw3u/cy2JXI3RW3WlCqrUO0YHlhFXkMyJ3sMorZhosQdjUGF5yApUaS6AftwccnT
AnsYYqPFoHAv/XSsLktrWOHh0DNlpMlK05VROpPfSZoaDsfCh2A4FPmO02Mz+EUL
DnRfCyqGT0kPDp9fA+eO+wb+0k1GQwJB7T8Q9+UAVb60f99I3fI5ryKyrjFAEyki
CZmQDRwcgIddT6KIJY1LsBeoqeWOYMYUXGh5OTBohy+THJpdxZ6Qpr2LYVVSOnt3
4oSAWOBA/enbzd94KlRoDu+fu7pBjbsX871hI6flkor0RwSVIdFpG7oD/sHHkYtI
s9h8Jx4gMxxoiLRbHr6+2WWBIo+jzjowW/AugmyGdeQj5EttRABNLs68EkVVk1Cb
Kx4kq4Zzv09/iPM8ZMyGlKXKCd2+iwhZQvwdZ5CAh5lJ5TRbcC8UAG2fqRH0GWLM
Mpp/7h9sCJct1nybx0yTcxdQudKPsonsiWHhEFgdCcN00f9+5qRdxHMzi5DAXZpr
z+sCgV9DCXvfp9X7+UG4KHJLIcmR52thTJLUAwyQ4VV3p+UpAAXKAfy3V7+vBqV4
oT5KbgToKNHeaDwH8KpeAkfXPbB32DzQ+37buc7/3XQlsr9gpaIhm1yxfugO0q2G
VA5CBn5HHmUL/Q6Hh76ug0MK1OBQJnrjopmjQo7YGf0Tf4pEcmzdSsOB8EcJRjcj
mCmoLgJpGEO+6HRtkv0FC2yjK5MHLWMcNj8dVUIcAYPMwIBzE/EJfF88z/20PzY+
pd99lVdR0b9yz9rhCfnamfqqi4ARkvjYG6mK7O2GZ0Mt+mFcnrTCjBWhbpWErWGs
BU5U1Mo98K8tOtpEtGHXR70Lbx52VnEWbmPTSV+cAKT0Lrue30cWuWbr78iVQYM0
xxyGzcbkm0BP4zygTCLrdEughNqdSNoEAI2d9zQuxmCb3wmdncQqz0TaeVb7j5y/
rHOuLX7RnfOeyTxUhiJZhnZIHDVWcjLD+PeZLQA96QVtxMJJ+T87X5GpZK7YW1DQ
KfJvhOBQ7n3dbAYCf9v0NzQc4BGf0oTY5CwwedvV+IpJ0daBNrmUYXXVaB3uQ6Ea
ymPDNybckZHkEmGCQJO+InRW3NwLaeeapn8H//8krXrjKaOndWFJV/xCjmeTnOam
lA8eqApgiDn1nifwr3YGw4hRE8tja4vBvIAg9ejYGwZJ6eFQ6DT1Z57JPoqMunSa
WZLlHhMEux22Z3UmW4EPS8w+PMiJ5JRp54lmqWUh+Y269F8JfzAVLdBwQgd1pES6
BQbx8PytIOc4E+5TFNWLZfntOsw8y6vBPtz/ZE3FxctNjR6wvV4X3enlrvWTwA0e
fhgrbJYGDrSux0lEajEcuc70LsE6slksdbljGiffl4NuMufDGIMy+bIggF80fEhz
WL5u60ccUQT+MHm5BWZRrJUpNGJyRhqKUn5EX+Pb5ev1fCOwUPTTcDyUjUsHPdea
m8gkjd4sDJyJPMG2ZyrIHFgDz4/nryyy1h+rnm4lC3SDaZnReNFjR2KSfSnDp/JF
V6LWbEpcVdY7l90SjRVkWL69lpSxN/b2Su8AzwLiRmwgvKYIWdTOOzay1qnhpE7W
rbfDv3+sYQRTbhLrgcylARZcBfJz5DSMSmyzvXiDzJZewB8u4lLQ/CvljAO6nH/v
UOLHKyzoWdeYT6uX3ytl15s51CjEtDiXleUaas19X/a/CzsFEUBw6jMztF40A7Rz
DAj00l239aO2E4EK1sQsa8dMNEAWsJXpHHj3qWdAAFlwJFJNdvKub9rNvJotpKJK
Df1Jf1gWkD+G4oqBEcd6jUPmblT5ij5reZ0gj0po+1gAX8SMqWE2b5avg9fmEtVh
2rsQNTeoi2SusxS0+RLS1x3YPC0fQeN2hkuPUkkCbDKg+DPs+GhY4QFxsm+8uFim
4ADlSJNCfEP+RJcn/h5EDpZmJwA0zWJc+cNJKCbKNbnmCijtLBJVn1huR8ZisV5q
KTzqAL4FcKEdJGGJgj2ojyRx9nUhJfZp680QmwoFT83zfroSPCzuSWqm8T6IcdIx
+IuPWPw5zpKu4QNizbbLN+eqaXZv0E8rzzzXwjxG4ySwrdMY6K+PyS+P/29tZj5Z
Co9ByBvYvACDNsZAcJBOUevs2SjHJjERcAc05teose6zda/8Rm/TCRLYvSQ4gN8T
sbuoA9IPMQAEB8+a27ttOsRtPPRP4fxTIyoKTEPHNxcf85meE+aVzc/BVeK5alYk
2S0lTP8a/Gw5A45AqQtDH4RgaJdOc1Us97WF+VIUpkYcFoJsHSGcQ1TtVL5YMcSV
84rUSKnRDC6hbPJ4rTU8APAU3vL80f/uhEAYdQFytHFqtHsMj+I8VSDP5YP/7L00
wkndaEz7ErrQENs0bQ7O+iSKzt5jI/K2/yEEYkR6rOt8fpP7EtRiryM3UATaiahS
2aLxZfxKz0miKow3A3owsOB0AEupuWd25Q5AbqedQ6uQEeAeIIxB8BMfFi+1pX8w
W318v0uP9wlnwqPGBLsE2udMNIHzzRhgU0U/4qUgkpjxmiL4k7v1IIt4G532Gbe+
6M8NGhP/208XimKUyPv+dJkDI4Ka2fLnytbn9U7xZeg4nNqWNyrLCDNxdCPWyGDb
kgTnsgSMw+5VYG1MpS1iQf5gMdgYImrlh2NKWhntOoYNsAHU7eh6+txgCDRHUqDa
YeVmRw8xiaMQw6R+CrXWJ1UugPPoXVtjgPjDF/DZGv3c1sQxz8w7jHlmrhAyZVsj
hUhWyWaXhV3SZXHwxc2yi9Mm/58IxUXFKHW8TpEgB4z74JIB+1I16n4wQOOy8Qqw
L3rsqn/xK7HOyQQbPee/r1lp2qyGHtTkEGETQxg6lBP0MYFwe7cewsXjh2cN0z0Q
aTl/R8kB+HpkMzEpGB3+/HYJ7lV0h7jh5yVV1x4Tg2QjZuHYylcQ++MwoHUdtIKF
hkWh+u3z6QX4/ovYVCKtPKP9TFiTxaROLoNVZsKEYVt/m1h5ufkmBgPSjP91RhJI
mhfmZB8EIIBRCGiYPZeQEAuQK9+/uxmPybXCdD6INJZGXXFDlPpX3Ay8hSnsBpk3
0dhKP/XmWNxuGEOWsTOY2jUNTRRiuNUP7ECPVOraKbMy+Zfpfbpn3yUWcns8KCAK
uE34Q2eTZeGynUCGXVfcYQ5PGy+peTZZwELwz6b96wPiK2lPdJuqtNdx0NvI+1Sh
3R+ovQ8pGg3SBj+p8dXQRcCt2Rnv26Sbvt6U1C7xO6H+S0a/O+iY/ycmRqMLLVMh
CookkNXfs6gPxYBR2fVQ+aFESARB00tKeDCSXABWX9+h0T8ZUy82f8OeGgS+So2z
3q0evU/LPFXrenn2Ffga0xOC+yNZtOzKKZkucbMG0nTlJ+nJ4fMTxsWT69WZb9dq
nRnKVGg+O7QFItKuGPnFeIy0YL3m4pD3zz4ejWRSify4nEhcNRdMW7VZYrpYdH/1
TCxXuqYjSphpmptlaoTmqYFvDO9Qu1MJqZje+2IKmkYBBP2CuFeiKDN4/T4ieEcy
8QaHyK8H362KWzZYijKB+sy71q93xX6Sl8VPp15EsFNRPa0kIoXlUZY93SFIZZtG
jm7dILwTpyQiIHiNz0B0uxa23stzuqI2ZjFz00Uzhom9BlO28blX4bSG3cXR/1hB
QI+Tc5atgD49UOQox8XqxDjELHvCr+28FgSbUv+s1GJuhvqgDaFNWYwgmHNyn3tc
fGm5tQOQj37h0bwd5uuVHehPGimSwFbIDgDQul0FD5hWxctYV4mD1H1w/jIY9Hz/
cwn+AmoicTIUFNhkxj0WmKtk5NO1cQgVTV1mYhustcTG2ErclNuA7e9p9i8oIV00
XemKL3f74iwNxAdKTgR60MziJGJksftOKaZCKzZXXPVUlg690lqc71qrtNyS2465
29l7igdwW6RI/DElC+/RtrmPZ61AWLCvloSDroWRMIKUvWEjJIiHitZMpMymRU8E
4RnLjn+uaIMDFklkQ/oQPJI9a6IAo6wKFpw3KZogqLcxLaT8WeCYZIkxD7z/OsvM
x8R+110HPVxvXlGLkG9hqmYoBsL/aXkAkj0Ugv3e3GawfKfb0vtZ/jwuy2KZS0an
0/+6nAx6PLZgnIF/FRwBc60EzajYDboEmMBEUHyT8qzfoADbsXdsxX2+1x8VdGjl
NbywUn+PRvTIZDGg3P1aOWun4ws5oYsnFDVbrX50v/yB8NBoSaBHaLlLc4NlYF9Y
KlnA0oJMzmo6/5fYhGNHJcWZTz21Ex9flIL8AtkeO5o3dlxCaG13kSkcHs8vsdEa
AVnYABSVDNaSBsIfLt1nBCqsPgIOi6fynDb98aeuEpZLo22IJRGSAxOPGDKymbVW
Ztb3Sk0kfH00raB1Z3J/Tq48gNj9DNqyx8mbJFm/Bz8rbtd0p8wUu4gkfZx9abA3
S2HRyUMjq7vN08aiRwCMUNBLw9hG0f42W9FxqKXWzqYSfrE/q7dT4oh82a60hoAj
Q6b4lzc+SfRm9gR7LdUc1IiYus6PgnuF9PBS4y/sTI1JvaOb6SirAy78LffPhBWH
A7GPa7Q7Nb/fTtT/BgQpEJ7SHJcXk1t0xtrO/rbYprgGalsFiH1G1DIW42yFxljk
CvfAi7McigAf8JUleOIUw+0a189zwP3NE7tyhrPrE50Vp/zM6e8Uao3mqimrvTP9
uKvoYqMzr5odV8A5+dFknBjuzHfTDNnBvEgwxW7e8+wW8P/BuI9tn79OSmMOyZpa
RqqMc6MKt9mQtAVgsgAMRz0X52OBmdyUHJV6yuvmRx9zzseK49kGv76rLVaAJwj3
ZSbxWx3/6X/kbpD8QaHJVz82gHs6uVrv4PwNVz6wBv/6P6s14M8uMPlTJFQ6Arc5
VS6l3CzFcrxEfFzqm2qgSlvlorXO1+cOFvFD1gC3XgxnRAhRLXtkP/ZwYPl9IYjZ
9uDiIBxRYqXuD1VT9cMaFiPgzA72om4++92XmCxE+E+3c7nNpAwJZUw4WgVzt5C4
smWW9Oc4PQeErvjfeCPPjDQRUJOvxsKEntBWY0cNnqisuYFhDsN7b5L8P+k2dbGp
LEQJPFlbbe9vwH7tD52PPWy8yHJNIDM7YHcNTjGrErlNAMfHTj0vYEOjDr0t80l7
cpHE46UQMgMwpGOhvryy5NtFiv+vN0JX6Jcs9uvCK5yAB204nCw0/gvCO2XpgVLG
3Yk8u0LpeId80ZTLTBybeV+ti6Pamob7xvsy2Nqsjryas+ROUVuaybcIAsY8cfum
7chwgzCU8qOa5EiewlZgO9CYiwJP2NHieJur4TGbTuw1F8o5ZaP9mxgf1Z49RmbU
StwscGZ2AlNuxKL4PrVmD+fU+oEhDoS427jEnqw6ix1KeEpo+fdlkNZrfjIawVwy
eE6C9NakLvVUpqaDIkoO32X/v+ekgFQJ4z3QvXuYzbNxl7YOzmXGA3UUYxQauZno
l6Y83XKkcFUhZt8U/N4d2ux13+9+5XuPBAVkaZvjLY9Yt49YVgv6s7wnOx3K+YfX
Z1MjmLH/+V15p+ZuSMlvLZn2xGZD8h6teo+rsjwgRSG58OU3DTHRe93WeZirjTFa
vtOjS/mM3MDLoX7a69olcWLcXtIi2ZZZgmznY/Duy3C7UASkOG3wzFQAsfveUogn
ZSbrrtf9VY2x240UIaIMUWmS5d+p+HuqhFHMqSOGJk9CwPfhbF6waXeejMHNTBYw
2AENsRFdqT8LzsmUr6LkMl2iS6Z/tKyfP0VIXF2+ELXoq9YpdGMVXrSEnnzav70m
r2x1qGBTmu7qg7kE7A8mGQ/HXdgyDBOZaTLstS3ALy/E0TSJ5ga5JZOkuznmFoBe
sOO1Af3cjPFf0FmqCEmkMXzULIP2npojq5BqidRa/Jg+XzsC73KF597tBeOJKMMa
a992N7pTJ/JaqWkbl7rNx48OUQRiuUt5Z9CVAVnHc8QTDjGgIIzhVKdMfst4aGuy
kyLMBYkwkiKpXzaNRIv27ArHeVfsfRGTIjxs2Cu5r5ex5DkY9RP3FCe/jtnu9k/2
hDdnyFgJSDvmp2FdbG7tr6zGf2xK5oBuZVZjdj0hz2KEhN8oSC7To/7sDcV8TPBW
c9r/Qs8vik6aVzWR1wV+6tZXb38D+cnICqbQMeiPp1DcBaawPHJdcm4uEQP20B5v
r1IMPAC/Sl0SsNd6I7YKQKROc+vQxrgMuDxjN8/cG2aDyCOyiFEez3qYENkTlJLa
nxU7Q7nDt7D+Ia+gHNVYWcavcFMBXQ+VNnkf37gIVuAvKV4l7pPy/ciEn3mUE9MK
9FhLbFqyTnAw0BGPoFPj4eDPD0lc1WAw6wzfIzj+z7w/zrWLQzDwHbbOOymK04HE
CDAP8cRFplAZRefWh9RN2gsR20LNUKZ3fLIvrVYMKsxQ+aEMh5q+nVh+jr1ep3MQ
WxEhDQeGq0hgeMyfHJhBod2BaWz8A7eGQGN0eV/ONON3LERQ2VH5i8QATz6h9B/a
j26LhF2IKvn3jLGYKmjxyPyFETL+UaJw74Ehxa//Q25z8BpMs5QzA39fh0WfcFc5
7EPUyxvGIaWIm6SRgAktESHY34XA7rGOA8tMsBd5c3u3ptNAjh+r5ri7v4KLOXyf
UYgSHqPgKCFh75psLrGFqfGVn+nl2njzzoyLTC+zIXILCib5qerqdZKc3MILSU9p
uZMDAT0svag0Ew2jEtcL+HnqxJDW9llLmKN0nDVlsuJkBrDSfwTEV1ohMXhr2KaT
fu6HfLh+URgfIaXcIafEtw==
`protect end_protected