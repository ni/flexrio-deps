`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6048 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
4NnOUJJFV2nnKBrlZQj+t7RfsjMc4346FJTtvmQANmbaD0tjj34J5kvASPk9bfc+
AIoDyn3WYDjYtr/y6BCdU43G116mamzWPgAY7mVDMyf7cOMRpRtpNW+tPZapv1MD
nwBGmBbJ86w4LlNKBphJa4pyO+pV0NhnsBuGWDPM8CGDC7nNBFie9FDXICsgCgI4
TYt6oSqM8j0YzwJUdcTbmABhi5RSqBCav7y6Bng/g2D5sJpDHV1p+8j/q1G/AWYA
bS0UCNqq2WvGl6F5A1V0StUgRaNRwNi6DA+ml4myLzgZUi+rWuLm0C6W+MFyP42u
I+xa2ynEOmzNvpwmYbFDrYZOFlMvG1I5JWdZfnfYatTxQbimDbYBzlkQj/+Gjh0x
cfMtZJj9x/U8KO7UIEhCxUl/ktpQQ0TD8Nma/7LJAqUmX2mNyx6E8irCHW9sINWO
wSASnkfwgAIsEhJZ8wMGPkqufz5F8tWyP559Kjjw8ljOa1kT9DleCq1M95YzST9V
4Xv6byfIFGloAXKDQraPRRAKU5oaca6PsMUJNXayAIWaM2rHSTZG3UKCZ632W+xk
XFyC1RgSj6CMMM6NwCsiKsshRTVMfMXAL0NjRNP1V/P88OsFhecHJuJjK0jCgb0b
V0fB/13vLhFimUbWXigJpmTpp1B5sJoDofFb7cfcDRi2CMudD4RmO81alfvW0JqL
oqc5oAzyf+6V45US92VamA5qd3fsOUiNegGZFAMpmC3Ps6txPOEiuMvouup9abXo
GcLzRuTWGCBO2E+PMncRlb+dNff0u/wwQHahIzPTLORITXr7/A29vFxdiHc9I7lU
1aV2/5L/axRhA8JGpW7bEnkVXEJk9/ynHd8ivNkEG2eFdJeiJ0SSCk519uEZcIz+
LSBLtPTqypZEIjbVcjT7jETmM+UPPsaASBydRmXVV9Y+4G14gA14uXJtC9ZK1mdS
if/BIxxmY34Ogv8llAJ1EgO0280vXEITBdaQrQWSSVt9l9B98/ZzhXGTysHmkPyA
hhM/UAyNxVVUyDnBYpO5IUX26H6jGSOfDePPMHdzMu0j0yc/L7KiQKJybReGQ5bV
l8/AROr0UxF3bdA+zoviDl/XKAfJ1uEUClFS24E8aM03od5lX4K1Eo40HfChKFhc
/ULYDTluS0YB0bvRI3jgwmgvLwUtuXt48Inlcd6i40OeRoP9b1ulKZw1+zUFAOuV
7bXNzz9HR0/74+yyOoW1dPTYCXyl21nNpWcED7I0201Zxpf0kpE2SnWQDAFnh6Yp
ILzs6HRVSQFeBUMRp3PDQz9mju823tJIP8Ud4T1TImyZYPyvLJCtO6TWZS36j6IQ
LXiO3t1dtvBN/9WABFpNbnceCZLEBHYgXRFXl47oJuV96thySBg6d6OYWcR2kCVM
Zxi8D7nZ6NM56Sl8i+wzYdgXNr1mXx8GMb4XPx0WaJtaJ49pDvsNj2RBzK7ocg11
GW1L22dd9YjgIIEJkXWewWkyHD2n+eVnvvdAfGsi3eYWRoFmKn62wl/GVE+IrEHZ
0QScjeTQQ9kUjJGP+gxKkeiiOmx3eNCx0rukvgw7nh1ixYiYSB4iga47VQLnvH7W
RoxVm4oD+w5Jo0y3OFFwc3oXG5N/Ie0VZ2tUG9VoY+5LEeYo4B64SdwRH65XvtvX
TaHKIniVNVhbp3gvLNYCdGCbU86RAaFNo6k0zZnDLyZq79vJSa+0epiWlLO3Em4G
mqxgPmmDh/X0ONTFji7i95i/8gOssXWvDZZvFjZyCsg+VyuBm0ZooqJrI9NQP9nX
RcgwbLiPa+M+TMwFQNyhxl7I7GrXz7CmbJh3NkeITHWgo5uCT/ZWjREaUqN+btr9
d5H/iftM+T0KZNM/7ayiBwmDOFTnd+EG3VYLjdubyGspfzXKOKEoYv2zAEzpdc0s
yxMmfSDKUHNRa1T4JS0kmpUn1N4s0msJ+d4AjJjNp4uVt0Bt/SW0qeQpgzCgq8AQ
OqGtUE5zQ1gSSQVLpGpP+eIPfG+hhd9EnjsHVaSvakIIlVt74BbM/38UoApXdw9P
P804tCrfDELSPT69IGtJ6IkaW2nC6qgYFiBmtsryS7B3soijrqdirc3UgsTk4n5v
gTyTY6dgOMv0jQUQBcSdGG7LC+NxPOV6UvEpI8L7VXpZUFb1qdUZeiw5/rJbyYEJ
dtpVf5WmSMQ/dsoIMJhg8Zl9ZZG5zWoJTpH+ALKtVbavPxLOVgC6sFGlyKKvqmsT
E3Mjbvq0+BDiHZe81lAQYILosF8gG5MnrhdXVolznJ9M5iXxRzuOPjsdOtcRYVdN
bPGUJpQ5sWztNIiv6h6ex4uahQQ26vPTNJ+fAwlUg+wGWRVMVhqGSArpBOx+qJRM
75M6Ckh71ecBX+2yOMHqM+jgJB+lf5Jjhoi9Q/DRTzChjigWBYZLov0v72dV/mdr
TsXy7Lm3x7pIW8u1YLtD+dgA+XPw+9HnqxaTbBpBvaNNex7c0itENbF4ND20E+aS
233Gw8KPl75FukYDPBbU1Cro+kAxP2ih1LpAxnWRq6yMraaWK13vN9tbBfSpMr3b
j1BRTHXP4oXAlodtpXH/Yt9SfoXPcOj6FrZuUC+klY27Q6lYW2WiLxVGobAdJF+o
Ek4a5dUaToES8JPjHk0sMYUKp2ner8xy2fyATyoiYcjZmN6MpTRKoZ0bBLj5HEpz
25ehdgk4iWcOxNh4oO5GdbhYvIjIwYgdzgotKHt8q6y0uOQ3myIJva+sk/riKoem
3WCckdyF4dhVZrUtrHPWdjrAiCQYTqdq6jBrsX3EtMoMGrH3KRbJZ46j1FPPbJHZ
gQXIFckLHXB9hDoRo1iVL4voIoKtvWmU6RaKjuWRjM3mgBapq1eVgoOiwkvWX+/4
jxicnJbgb3WK7ktks/P0FHFM4pHhVPOLS934MAaw4HFB/fKZTO3C+KJt2ZnZO4pT
LDaReHJuE8B4Z64DtS+ggbE6BNLRCzWxicTQd5JJ/kSpjF8JtG9NhpR09IrdIcnn
ZgYVYaz1K3xWn/Xdg7UcwtxAukUv44n3m+tITliiJ0hFNtbETP8DzAGBdpfE+kax
KzkPujJyR0QVmtOZBJCV30nSQNSDzog5Vo55FYM+jY2Mbt8BqHk2mPGz4i9XC82j
VWmSJXJBbaWGynilQCei0s6T9RqhtjX7l64a6pyJURmJiANUdRuvNq9eDEGc9s50
Qez0rSI5Z7ozZpC8oElYnGbstzS1tgkfhGkzQywOaM273Z5sReWdj+mceStXM8Xx
vOEO2AKatrekvxxDjtujaHL3QfA19qfDNgs3nIg2qFZXpFTuNoac17ppR1UnDm5P
qW0BJyGiYrOHUAUJwcDG1bB1XDpydGgp43i2rQLDgn/RixW6ZmpU2x0fUTTdE6Op
Zm6bKR1CSCrSXaMsFbd99LUHPVR863/bgyN9QzrTGd7nygunzzBerCcAQBCYI4j8
JNqMaTNq+q4ZHS9XSuOnICUSyWJg1VThMhBYHW40hmtlFDmhWALYott53M1m47te
QFtPGXwuLevCv/VfgQwU15+/JLu13RL/cLFqPf51IUth+IyLVMootGN6Bcoq7K9p
horEmq7SNe4QxU9h69YGw2havR1PfbND3IU7XoU/PzE6xbVwanNTfWnVlT70vs3V
/0aCheusnY/ceH7fYZe8ZSIKlGST4dXanl44r8l06dsfsX0FyypH9cNkT9zzU0fA
6y5mpLpiIrNZ9V0BsKlF/oMtVfb/z14pOraKPRVasIE1i8I651I+V7x9N6u6Jlxq
Ier26ex9Min5yKdm+IBcLIO3Re5+wlN7BopfdxZh0EjidxHoPOwShK7pFgadnH+9
FqW0rP4JJCEQtvEc+hZgo+uJ5VQRwBUH7ZGyzl3UmESsLgZYcpBW2+6/mV+WOSOU
8HJiIrTYxlZu4EZHfktujYTAeB+zUxNH6rcFZrY2WYCaGNmzOke+e+BtuY0z+pO7
tndJhn9BLFdjA92M6RIMgzbZ9qpGJbCmnnEgkHKWOMRaQh59z5zSRoDr8xsZ0V50
QWWtNuz0p7U6QuFQ/uZdL4GbuIvVfIX8YkY1UkHVyeNqo2HJi+f9VTZnPIHz/NhX
qgDE0YOZUHLEc/o56Mcwtt6ceEfHH21+CqIl0C7UmQJuOWWbbDdc2MfhGzDuv4E5
+1V3lmPcmW6aTPBGM1wZpAz4eZffkhsfANWaTrpUiIRhwGRf3p1glgQjz3zOnbdD
xohW+sDkaFuWFl/xoezWfRrCBKE4wLs+ElTvzx2ZF5Xhdef3p6HHimltMH4qmsho
iAv1Zzt9MtOvzGvn7+jiQBiYKWH2uX2rB7CNnyurUbg76RdxO2WVczAWd+1N5s8T
7iJOVTQwoTZnDCUt1BecXVqR1QhkM/RsfO3fiogzTLaYxmdX6KcAso9KGqUwY8lB
gxlT5myFJEvT3R8LAu5Z+uuOj9rNwq6EyJ3a2YpalKkBroI8nUnlwETlcvVmRBJQ
ylD8A4xgda6Gl7hLqHpKFFh18qDpsZNAf8ca1y9QOb7lZU/pXcGC54bgdCKpV/Q0
qlX9nHqqfTdNAgtNfh9jDoYDzjv4mpJMr8gBXaURGih9oPYLqaKEV4UgncbcLkWE
1BlWJnq+gONPIg7KxHYoDCDJl2e4SDBDsaRlh6o/ZEZbG6R9bHf0Ju9tMCpD597i
uZot8rHr1IGtgHF5V5ioM63Dqth7nu1b6qdOn/avUHo1OFii2BMaD6P09wnUpz3u
L2m/NEdMA5kDu0kRDVKqX/AKRv3NL3DbAlxrfZJK34WFArsvAeN5obaCoSBplGob
I6RzV87BfAdUPTRg/1LQaikwpU3+b2CqiVFbQi2hc2gmnXbiXT+zw5lIoykitNA7
jn++6WHwkYCGB+8l0uqnYMIWhrUL0/ttxqJ6s5jena5Cn6tQRU5otOfr3u4UGWsW
G5eBJPzflEBg//5FYi+4NEkLgpOxbMUky44Tg9A1Qy5oVevKYvsvio165gqcuMX3
hZBUZErRSsSELz06aY+F1Zx1RLDQIATOLKdQbpb5C2do0orRpJ330ZqVbCld4FH/
jiPZAdYz6RnZVaBw5Gr192HuzjXiHjNnlqcRpV/+sP0qF5/KEMUGpDvJNigQu+HS
oc9o4CXU9KsX9C9W9Z6u2vuyJJLLynjrYVgzVpMxLwo7/n7c/uP/ot4dfyyPhW/x
C4W+4DzPRjWtwxjvk5fqac3Uo0Dvg7QYwxtTGWPSCWSMgTXYgSkHOypX1T52ZDvz
kGgwKZvO9R0WmezsLhc3mqkNAKk3Zcap5wQRZManjsRbTX1h00GevxwA1koxqg7a
cXyHjxRURj08YD86gWJBw6833N8wppEqVu5WMrryN7RWO/0T97CBhZL9119fLRvH
aSiu2Lua1kz/lmNkQWGugw9Lxnj0yr0gaDr9yJPdxj2bv1OkkP5qY9slHy1s3Tdi
PIaGo8PEvPpjoeDex3gUpEoN4fIPpwjc55n9d1IhCUlQ4cPIt3hY9PUCV8PUBKyj
b+hdU7siAm+d8Nlx2AcLSH0XnwqjnOWsSeekOWaI2Q49OGz0Xel6H5pk7z1z0hOj
QSC5o4k0txz4n0kH+pqvVBFJGRrp850vvhymLNAAYiDhP3TnRxZJHY5WMClSm6rN
UkzFolIhAmPbXQVltp3IaAZ2IoHdd0iEQ2eA7L9u0zXVuiMBxDd+YQPQCinjDYkI
76R31ol7Yw4uGks6DA5nNy7PpnM0t9qU4ixdvceqKAVeQv8QkFklHbdSedeBAMpF
mnpTs3OvAvqP9UGlSqshQvoi7kDL87MRu5oN9gePefgBmaJfIiZSm6PP4g58NEfA
J1tiP4OyJvwPqh+0qRoSl/UvaESEeYioXeb2ugljhPs4qpHdZ9IjhLVl3/PsRBbw
9GGui7HU79OIXycz9qzFOmMd1m6VuQks9bp1qUUZWe5MWJgTypuctqu5n9KNjjAJ
mEvnug/SdxlffVC+VIrTDK2r1tuNDEnXZkW+wrG272pKZspR5WcHjNuUuPFHjsDC
z+y6xtgrkW9bWmxeat8xXaCTx8t/ZeuUnCctWjll85tI2oW/txrStYO8Gz7b4ubm
oN/qxJfbuyJbNzKox22HlR9O3Zv78nPXoTHSXZds/T3d7kuhnK6dIgji2vjJZD9/
tJaHnJnsSrCrhzhjpuHuB8PmeFTnzZ+bHmzZKk/tTikV8TVBQLidktbKahk7IFba
tOsXA7oV6qo5jK8+i0uGppKROK4+MH5uVMov5FmGJXfWco91JeyvDxlTETiFAFxD
1MCj8itmLyfEF+sx5O0ZhoIvaVqjKrOhaGNTB+mos4ude0MGvtIsqoea/uQtsZGf
L7/tjN1PoV0KD/+hu5QMd2MT4IBV3rXPUVZBSfhN+YL+b4JzhN/cO9h9s3kWn193
wGKfYzR/YCs/9DCZmKNcDGRf72esU8CHrtGK5/wMgQoMfFqd2JjNkDOEcu07d89v
AQ8yp2/uOzrOzQ22frp0rHoJJR/RAvoPWqWkhIsE6/NRJ9QfmHW5qRteasEc6qUm
uDKJ09cQwq4VhKVj7Go0Osz5SuzcQT1X/jZyndXMTtL14/Ov2HLJgQdW6xFGY23W
zsN9QtXMQEYQF8/n+gpaDtymTuknzNZwMZS9GOsfxmGwrN6mM7ckRypKWIoMLBsi
aq5yCVIejkTy0ZTxOO5E5kZTnAI1P16V0iYGN8soXG6d5xZquPZWZyn2yoEiHPIm
e0vhDJpydOHmamf9PZ6Rkrm3KSAS86arwaZBFI6u+9LHdQjObedBr4kFN4CVf9St
9dgXw0QuH5xxYeaHWI1XB3jhGN8lMy2qVYsGvhFBHRd6G3pLgD662axACJgmUqTz
cjzu2/UJscMPq+bqSKIydYNxNdXHYWIVIJAkUnWLG/Ezj97Ajx17ADwLEDXBbhl/
LPZB6MRkZhv2Z1uW3olEifhWNfftczdHAvhygqXyqgtMvL/Jk1nbj/nK0gSdr61Y
wRDDFnuYR2bzF8lpJqSvcNvE3I9IVhDEJajgbtnmJiirP3tXrZkWVf81oLx+Fs5w
SdZ/I6yD4xD0HD4JlEnmyXl/VX91EqPE7PztWs2/aYyUOkB4g95GQhF2M3X55xVF
iMGzslrDb9c3GMofhDxvyEPWUXwYcEW4aetQdiltBGQoTEMI49IRPzIADv9WsLeq
kDWCakLaQAot5mMOVlq21SGlb/ddBj12clzi4e7dwkT5Gc5GkxB52B5QH1VycMRd
Y53zWLDJUiCgT9WFG2h5jEHpBCJyll/0+Dg0+yzNm2SZYyWDstFyz6iPejX8g5pB
lfFtNZqL0YRMZpblP97d1rp+zSkU00YlPVxszkAyp3Nk64sf8QcSTdC0z04YXMpv
SYrL4OLFMlAv4lwo/tCcvfdSUvIVISvMmLKvWLZhBJ9IrXtXtFvfzkv3d/YZMveb
7ZE2diCn0weSZdS74jsQxXsfx445ZmWHM946h7XqIV5mlR5fCev+MZUFqqWnFxff
BQVSx3C13dYqwQqsgiGTH56tAV//Zxbe9aZtmXKvgXy/Gf1x+SFuMPMhn8IoPpdK
JuEgVaR9tY7WrPcY5JtdBRwPvLlV+vGDWXomcrKpwvLLuj6pVLlUCI5k7xPbLh5I
BUz8gYqip1yWBBqCHDT+/3dwxn6SoZq328VRYEWbqzYq3K0brQ7cziwarN8IGk2P
3SJmFWwCLfabi+MX2LnDL2aiQ2ihr/NNjn4wzBy9+JwcO7PmbBqVsVXlt9G5AbQW
0E8eQZYAmA/u45Pjmef5RABsGpWeQmTpqESF2ttWOs6rCPlBJ7zCYW0vEmZAozSV
/Z6zF4b09IBLZfpYYZzzPa1cocfopHq4tcnTsRsgQG5kzmWbAtL9IIRoy9tGrmC4
SaWS9IWmvLxP8JoZepWr34jNJ/pY98pLQQpse0bJMlJX59wNEpdKUwnrzS3wdNkO
`protect end_protected