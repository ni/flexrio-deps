`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2864 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhAUN1Tg6/Lt8rBz7kpeJnZvkqEJUgFMmnPYYnXTaEG19
O+PqujiTadj2z9Vhaz6tMTRD3EZ+d5fYIGtrffEIgXWYOM4oU84pvht4+jnGvMWJ
jtEZofP8VlZhhcRLUZx4FmqcB+V6FV/ShrThkuT6bVQh5QGrpxinweNbSnXryC+H
IQPONPzzcyAd+aX7eYmiY7/2nnDlIvW/heHV3dPvCC22UCL5YPh99mSOwW0WTX+1
JJ6BAFQH3dK9HZXqaUhJgna2qdFG354j65pLhNjICq5uTcO6IvQmOcxW/Mm8Badd
ZrzMNlP+9rpv74AEakupE0Pz69wTzUQ5Q7FybxnQNQzPn3GT266LAkn7xV7MGGCK
FkiZD1M7qskR23YQ5c5oSe1XlsklHnQU4xYvxBWGY6p8Hf7KNrrElvUH1stVKJ4V
nJRh7zUIxgD+HI7ave7Ofpt/jkBm4zHJpmyfBqP/7br8BQSbG/7si/OBG266UbF2
kuOTFX9X4JOV/O8xDfIRzddhwD9zOR9JOHsaP44GP9tr9+f2Ore4ep7ysXO1/UrB
I94IHaJXBL14e1P7vzvl4dmfWA8KrOwF312r8V9k+nub9yWvFmzNwRa83ubPKSL7
+ipNdLQ7Y9J1C/LM8DYiIbtg2MPPbx5I83YhqqgK7yX4Mr1uZOSIdVtyKrZtP8uR
CTBPztPPjRw2l6bpMnB4tKSgC0MwHa2pMONb2H3+42VleXZm8eFpbZp5+hzGUCOS
rhEBS0JwaVMo2GqhuWDebsOmI+HZMDgTLHmu7OAkSXYU/6GWHnDembqhf+leqWWC
RC3BLIaGyc8pY3doWuQSMis/4Ih2eulZFNI6frpsbjizyenL5HsDUAR0Rk8pb9rm
2us7mpd+fzKx5JVOH1HkVae77D0FP4YKGBM4h47jSPyK/sjL1BVrQec2q4tFi45/
G+ffb0ofywMZ5F7jwH03M2hmcCVfdgFNAoVfypgDeC1ogVaTgymTOknO+4U3Ddr3
ISK0gihbgOQJUyeXNjGe1N7I2DsDHIiE7ZBs9i4hgH4+XR5c2Iv6vCmH9CzZDYjb
sA2Yy8T7CKEqx+5NRGjDBvRREOfZlCKBKU7zrSVkgfG/7MeC1vtHkfLxKORmwdNz
4zCLC79nDtUWATbw+o8lHxXecdJDFoE4kIPCd61Llv+sUeTJdH9fgF0Y9nwch1EJ
7L0dYk1oSucx9mV2jFBgLLL2j06dA5QzgfTugN6geTFrUOF3P7dDWj8x4MHHKsOQ
I48psuib+rxV2ZnoS1rMXQUn/RRkNoQYlWlmctYv78L0Q4+JDtxqPK38UN+TOohO
BkI3zhN41VFuP/yrvpmwRqIYkpKuJrLq1wF+NkJMFmep9zZaEQTdQFp1YU1XtwMk
8vED7vDdmgUeTqw+WIFZ/AOk+tDLkN1ptSnhTo2x6fP/x3J3xB8E6YP6dG+E2Otz
KIaegfB4wYGt7XLrNe8ceQASoD8C8qwZbFrigZhq5WC4x6yCiW/fMQprYrW5O55c
ikZ5Q9sUhRUM8WnD53+gLkhlIt8WXC/KivonE61Fq7mEpSlFsTLBPBfqCjDkt24S
FGHPDlV/yq9XDdRrrETKHRVm/vYUukWALJFi0IMzaXzodjDJzq1ZmAOH5smuWTRf
OsYpYtgh3Jkl1nQpumHVtA2ysOzalls14lnFP6Or0L7edMjY6JrEox8xl4XP6Z4k
WcYyTK28yHa32pnHIpULRRUKC7ayCKD1EcfxhRLEIcKQN92J7tVQNbQTaABk5zfd
XSuuzTzf1SJxjnAcsZ4ksQRkrsxLD4XDOIVYgLfudeyWk3nMLvzYZO4g0CilCqvJ
mWfgdZxeEljMMM9uDqmULvmIf9mrIH8mdvSI3Zj4nwwxE0tbTcs0nA83s92s/pXm
Gd8ggm747Z+DM2aDufqD5V27KoGJqBFMF8hLnsQhqW430hM++a9+SANEDMnm3+VV
zyyYmGk+y0vUAHnHcUXsLXw/RwAqLrnnS7S1+H2WFTIP3ZgcYBsf7rq+io4x6HrL
adpctqVoYfxmYFVnqPFmYRxlc2BxzTHeKrNFuf7t1XStZ1EUEOPGCxtyHn1KymEx
61FZH9hCXZIfV9K0xPLF1XUi1ZPWuNs3ZLo8AW/cjX08tajqS+3F4jAcWoJwgTth
GcyPvBd57YMYwYTVV6PB1w4R8LfrxMcYtyPxyme9zO3X5OnUXMyxCcgQijqWFmY0
N/cTyD3T42/eD97dZmELnS3+ckrsJ3yjjY+q5deqEINPJGfn4e0hdlCrrut6kiD9
9j1bpLpqPmwz77r4kWi2TzzDsphhFSVihz1R0p7xQKx8+BlbY9qlAD0mHZUxm20C
GMt0fD56E/V9/cNRHO08VRTNwnfCYbuD82Jj03ciRKFm86mCvOfbtUl7gyICBOxC
neOqthrRQp9eGg2dRHfFCqEsNToWpaJeWqdy81H4jdCugRBdNNxdiv3JfHAHeliN
BAzcU7t9SSVXbnfelu3EJwC7sLy8KEaAyrviIHz1N6M+25FoSCD86n5u0HIPbeWt
2UiygTpuJpCki6car0dz9jYREkuImv8tp4Q6Pr6/WTkbZe/rzWIa6MBhLouQWugm
cVLNhKMUCbpA1jbBAS0JXXXpQszRY+WZknUvbrHOFuECxJoRCnHffKkITceH6yrS
+rw8nbCoydncjwT13fVs3SlzC7KXVs816tLh7KFy4FkxP4qbeO5fGrguYrZ5zeb2
i4W3YAu2scIX9H6z6++GvvTPE6tSu15rviz8NkT+I7GdMPVdtE6p9KmJFob9ZbLl
Gc1Fr2zEzngMHAxndKJcnjPT3pMafgU+Z8+hWu4hkeg7vqsrOvQxjqbo2DeyV4cq
qlLZ8vKP+MwGu2g0oOSuUKtLN8iUiY5nqft4e27I7A2EgTKzhcUflFaDTs+fB4+S
9TTmTDNdtlGYi8gNj+FnXDrwTpsnnrZN/m3ks6VOW/wDBiGls5xKhWa5oAtf4Wo6
GwHSQz4vLGLiMEO6zZ0S2bhyBEiul9B5Kh03RKrFDTIAvkw8Z2S5NBx+lPKU8u2J
NYUhL3VNF9lgYc8rAFtIIIKnI8olrcWcpBUgGEkewTgBHs9RvhRoBKVA1wmkjcKd
eB4PxOgGfxoxs73xAIi8llRs2ngX8UgrHPh/9KHZazp5xw8mP0rWO8tbmbhI6yYC
35Ka6pAS9j1kH8XWgipsKWgQXx6qqXt69f5MMj9TLS28oEWwcG2rQLTirFUQJI6D
xUuQyD88K0tc6dMcfh82UHDubYTPIk8t8t6jGMQgGJ4CPHZDmVwqg+TtriFhYL1w
OTay/G1Bdz0obDMTMCedr/96GpZH7eomiX9vIWmvOBewPPVUvoeB5jh13uq8cvpC
PXux2kub1KggW+RcQAHepgHzFYSYoFQzy2mkR/KWQL9waIcY5hZ5rwEPHsrzQ4Ri
H2/KM5+WAAGnn7yuRwimbCkrpTs5q+fN4yPpnLf0o3Ej2IxGmFw24PoUxzxq4UIh
NkVVmp0PnjF4W6YFU74nW/Vh6FcaXwgsKwx+AAr/0UL9JwfSd567jIfA7/0pEaL8
W1EGttnfEGWwuOcXFUfqogtH2bRA028MDFePM/oqhg9DeFsnrQCpckSPOsysoKza
ZZwam5NIFmRgkIiTULPovfKNZ1IlBFkmF14kPdtnkCM=
`protect end_protected