`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1712 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
LlZn1WiQnJx96B0dQWSsquxHKWOA3beP1pGwRkQvF3Z6tfHfjf5al2v/7zCrQFRY
rTqHlC9txmupYs8sTRIG4ndW5yo5u8BhR+KzFTB0hZIJGHsP22pcCCYu2KA2L3Al
oriytYln/tA5kxIwEkSQNnyF7+JlIiK7RHb79/myQGE0wEC8R/Y/brFfQDYbF3Io
rJ1+79K+sF+REYlWVdlCOpv7qhgZ4AHmbQyjcKghNmHI+azGzUzAFo1q0xIvw9v6
ZCBkQXYKtuLaXpQCWfgHA2JqdOM3pWbIiPrW22SSKexqEbmvVP54jrambcb/kqBH
/gQcyeN6fsMbtKz0VLWY0gbTTwGblBJNuMb5qd0W/cL8fLmTMoV/eFS6zvvx8slZ
iR5HuH5FxYvNkBJY9yXYjUCnQvtSOoOR9rn5de2499X1oUccymyLC/4YBjduuVgI
quwLA8UkLJD3NMkaO8icSp2w63yZqHfM6p/QHiDSq3gYFu2nAGl2oogDEONoHLZ9
pN5yXAs10CwUqL65mu4w5rFcxFRm7IChLvSb9kypz4Q38Zj1XoYt3ES9qHWa+Vzk
9+8C773hHw/arxBg+hqRY3EBrs/JfN5NUFh3EStKHpXuY+l+WKXvg4BnU75xDoqG
MtYjf8P3H4jMi5qm8IB3+iKJsggid0BdUcaZFzG5tMCC0IgtTi9CxMXEoyHFCsYw
0XCYl7wB7DfUpTAdWsphDeLg0qJ2umn3VJaZm7/UXD5EKzcrZL5FUukb8k/okBqS
oTMvPn1M9Q7KYclr2Fikb6LB3fq8IqJuy4iNBBLlBJBEg5UTKXTa1qGVfiiQL2at
HdsnU5whzD6S0M3QMYFBZV2K4hVY4/GQrrTJKVeXfPj198faVubwz8WAUq19l4o7
pEQItBXLNs5Iwn2l7tdTlg7+1tkQTsFTFaM/k59BLD5YDn2ttfWP2YY/Rl8nvkWj
7YACLOwGzzQwb3YEQ6iyWRBUMm1us6kS9/Gp35Aazv+H+/YxIBZMtJMnlXoqE2zl
7/F4CNNll4vucrWIvXVaDj6JuGpEZfV4Q6zQJjSHM/NXkexahamPwILmeTPf/4fu
K973Z35lGb46DBYifJDd68UDI7I/AYnepjE6lcU1CFRZVVgpu6U6vMISFlCFI3Pc
ltSvDyP6Soq9GTEkWWb6PpINRwMLNWj2CduJVyjTyTlpvci03w2V359nj5rE93Gf
7Olqc6hx0ISx5QYYdxoHPpy3ySMWCtUyFsrZSToOaqqWXJrKzWLV6jAiK8o1tpin
M1zuIMqBZYiVK4mKCygjj/2qxw8bxfnmIG+WG6m/rc+zi+3/3ZHJPulPRWxWMfOt
IBPdzIjcErOxUef//x1RdUi2haoeUtyApGRqM+pWxtaxSnu5uDXotmNzRUl60z1p
jI8r8ZcDDr4ZaaEc5brU6W2hCOUAtD8O/lPBzM1vtDahhcXt+pCKmh3sEVTkzey8
apJ7Aj1VpP6Wz5GYdxCHZzViORwBRqVUFtvN0SyiNBVcHyQrPA9cLEh0urEDpMnB
wg+EOHKVi3FCXS025DFCrPC65OR/GtXXus4Tc/jQCfxjkEHk4lblnwORO6wBlTeu
o3LQaSjCcRahZg9nxX41rgLIeait+ZKthdV+sCK/WV5+SvIe9y+aOBmCodog8Jbl
iEQfk9iS4zooYNpTh6lQoR5S7njOpAPWqat/YPSbD5Tx3O7Q1SWbaCTU7vu8exDQ
iU9CiwAM+mnAcBIQ5+xgEwzy8pO2z0p8lN0vqRNP0cx5g8urJ8koAj2Uir36qRZC
2/POnVgsOtobyFe0wrJtg5WVcObSeM74y559Rdy0eMN9q59LGTCDgYayCVTHdUx3
K+z2DXN3J+/iQPFEeFEWJGlehRP1MNTGmS9Yuvgk7ZFzDGBz1M0RwuRkUVEDnrrc
ODs1xeDsEFYQ4WwoE/kVT8u7Iqmj3NfSMzmTcoE2Smnmv6sGAw0KmkudE4cAvkN8
nKMmysWiKhemWE7oPYStSUBvw92GVgKjgUDAzb7uAvVywnEoE3IigrZnP+e9Y5Fq
zFWHb8RUuPRaqWtYA1vNkqlS0J+CrVsSyiDdxgkQGZmbl+9qcFMxfYr+Rj04UES3
A07YKdniaAE8AaE1Na13A0NS5bnaiUb/0fwDQNRjOAI=
`protect end_protected