`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7824 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhFhUxZEeYOohtnnSQTgbE18xmbQA8229HTO9+k+PWoPG
8L4gN35bC6dbkfsizDLM3S9LcoQeq0AGPI2+Lzq7jEKvhMTPIlF1lPWh/58s9gbq
ncaPVWhHp/JM/MvpMhhFHzISq3Nj7PIfFGx0IcTdzLiHOzErShuTJ+ekjPw3saQO
Zas040K/CEb384xPzCD68QIKdu516NpAxMqxE3EyzoPaUlmTusCm9NvNMLxIdFbT
3FHo8rtzyfli87I7+FWpbULrrH1LlQQ2I9gWsfxM4ualtpLaR44sXOLYm4v1/Zzv
rJGmdY+DRtttI6+grFHVb9GMfkda7Zh382L1FYwh1F1hlWTvVgv3Ii+3yCn2A95Q
OCrUqastrksl11S8v5RjHVRRWJeDTsB0Uh1AYqiW+m92KnQmREPja0rSI6SAY0wW
nknzCliYB04G6l1ubKOALPfMVUtXtuYHxmxCV5NareMDyLCJbaz9OzgbFh0wXhgW
sIhYYL7OxizSF4oF9IB00VyW2GMOV4HWXDaOi6O30g2sgYs1M2jh2xfXdd+Dm3EV
/YPuYdu+kXAs+gwV4EYFZDVan4IifC2YHodMU/ELvYu8yasnukhrqt+nBEfuovZd
EHC5f2lWm5/9zFf7BBl7VYa37wXEzeo00pB+mIPXKOL/14AjU9Lh1uBFTrDQM4DW
qsMdLL/x/XAq+iK8RVHzFOyVWj5B/ZXGgTvWX4c0nrOGHRUOgswhjhuiW8Yi1QIe
vSLPdY8yfqoPim/QqJZvJunsLBnlVYENc5mlzV4YK//jZTgTeRExI4tbVmAG+kFM
Pw9FXJKZyqZj62pAQiESxioCUIuddKtGfnQbO/69LnK0qJP4JaVbflIgM6VXaJJH
ExxC1fErhIAf9cb7CEe/IzmAXYfzR726SQUHfavKV0Mpl3bSGvUy/PHRPl0guVZF
zj0if759zYOWDfhgHVqiNPTwn2v5JlwRbFf8m+gz+t4Bn1asY+ARMxigxYebxzw5
zD9BCk6hONZcO6vMhOddj0jzyNz1I6QNXYUdgw1ccbYbkLmjlfs4vyio3W5Tn9mF
QlWV2nKjhcoFh9e3tuJkUPK0yAIbLHnt/xo7p1+YySrw34nAJNqxu7sV8SyWVyKN
P/+hTTXgdx491mNcqEEahAvhwB/3SiRQHCoCGJMilpx2nfZx/4t8qIXyDpy+PLxf
XBVoT3ez+4aoV5YZLQFK0q9VneH/GpJPs425Ibsq/t5/a2gLaLst91s+pUZYVyXF
/NEnbBS/a56WZ9lb/OFAqdLIvA+ZJtIdAsuIYtYzrZ7M/Htryl5W2lnkozOqvZRz
bMRJtnOmKsMCSvNPSbT8IPW1Fz94RhuOy3Au77NSZ3lhdRd4s7RQIQ4NFh2zXMB0
6QwqGS+gJM/Qw08O7ykqWBMEfsBtYEVmGOiLzzsYvC4b2Q+quLW+CKEUKQ+Dth0n
vb8dO+ZEltEC5l7mpWsP1U+SfUrwsEm9Ii+2bke5J8LVZTyyDQ6jgSzmmDdKrWHh
6fUD8mF+At2trLEUYdEkKfh9ussHwG6HBgsgIWP7lrRLOk8pIPy4cXJijJ+kQQ+I
zO+A5N8yYnZZtSSKxPgIsV1eCAdhRevoLOCXkEpIYy4KkPRK1JPvoITYuBnRgW4+
CTyE3a2Q86Inafw+WXzkaGr24O17jxY4S3LANO8LGHMH3ov4KaOI5V5XrcINQqB1
4xzoIEu1A6JWRFujEhjhL6IgAMHNCwkzanHiZ4rAgrWvdJ29yG0yRWKa2ise4Uqc
BAWqeX38F0hNmpc9hZ1HoDy/YJDjcxpt/Neu/FTdKuAyihOcMjPQ1NCiWnFll/EL
Undzts5pAbI77bhRlrqr2wL8unDfeHBg5cGhFc9viNw0S3NMqeyRqkVixkEJ6GTK
GysVAQ564djDAmp3ihak0DeNr/6YvFL45zJps5P9YeEIOAAI/ZDfBv7IDUrfD9RB
igCibTdgwlc35gUIcXoIuwlBHaRHbXteClmMViYpW2rpU/vE/f9vCNhLAwk+bJY6
oL5OALKhz+yXjgQq3MqCxONEITkaICQCSxgGHPeoBVwZ8oMqPz83+8CWgHVxjkN1
LeHZshQCr7CFDshZ5NPDEUY2WuSzXG1LYrRYg/NUCdqWwPukUtwLn5ilM+O2dPI/
MMsUv3Ed1WDoqtQTAdI9AFm7OcWTFhFhnx9DggDpfkdi6Ez1/BMOAjaaVlGdmUeK
PeCUN0CWLSlP1hJXnptbi3dOAELAETKDjYaN2bSfoqYa9gFE2ZBro2rRlAlPHSdL
TEEIviS9f1LRgodAC+gjPejvkKHYiI2ensD0MTgR9NYcILLrWlgTS5jirV73ut+5
Zdg8gApP27Gp2uj5jl0/x034CM4i77/PWCOnWYJXhpKo5JjCNJHf83DZGzndEOe9
Bka+Th5L1/l6TVB4pof7FkOTQ+3ZBELyaEZ/fTlIBPO925LXLveMQEP8HoeWqdy6
DXzb6ARhvUD35/PF9e7ayPpjhpZGEmxk0bYeuyZzsBUph/2kB3HivMBd6wd4p6Dj
TKJZbwCF6x7FiASC9lX8hN5CcbMU8Qistf6trTmavCzgbw44jJAWevPX6zWdfhi7
4k8tPFC6dvFzHejzD2LlZdKYzkwiBk7UhGEdNF6CsYnPL912ntsg3po8Qlc54+o7
9JMmPzqyetUAOg2PtUyEq0N18Ee20m2r9w67riNB5dZtB7xzFEydZnUd/WD6SGKv
mjOPePGFi5h1vh2vU8jjWoHKZvfuvOlbHimyBcSC9ny/K/Xk5heXpj9wayxpAQ0X
kuaWaaAwue2911/R4Burr39TfHMsg7cUgdAAiByEbTBXjEnY6Y2RhJu0qAWd4WDn
DAXJgamX4v6+FPnuSr8Q7Y+IJf0uVNrg5fWbe5J2auqF16c6baUfEJfeSzitAgp3
sKkHSmsxWGBsEoeXwMvRFyf5JUfDb3jxYRw9RY+4rYVQ9VMBToH8yoLbLTvDOHAK
32/x2N9uWTtakWBnsY6Z5xKOCxKIzg0O2u17B/ZbqINKTUGwwr39FLlaEIOg1BbF
qSQOk5XgSWxBIz4PT1NteLLljVcvJLe0ZQpPd4+uY9hoxUEAUpKR2k/7HeheYkI7
inoOe3PCT3OWbpWS35huUz/+H3gb5yAScHGMT2hm8aOAdH/DN0XMcOHIEvazC151
HpN9kweQ+sC3m8dOmabgyyoP++RZGRH8cctCJ2nBjRG5+AwEtdFrS6LBA+kd1qqe
nUt4QFbNSGLkLZOgmwJkj0NGE4ffycNP/wWD87h2sbVyEY/+t/3LZK2MI1321oEF
U3ZlRYtmNFunQ6IAAGPXNhJ8dsqU/vvw9HXaFvfPTIVCn/Xl0V5Ttv3s1dXBUvAh
/Q1QyAtaJbu04csIhLiTlSsN1PpTFz1iFA3vcwunS3IFLOKCpKca8mYXlntRBub0
NIgbfp7bZVU/SkqeOtjk+K50Phx1C11FuDgyjhYZWT+WoqIZWudjnLNvkv/LW7A+
QAteOl1amUmkhi7rtN7pxgFrpzYhSgrmyVsmHg7vcxd/Tx8zCZ1kF9yw+GUAzizr
+NgfCXhVxDgT5zhPVNI/8IPC2R4fhvjsol6YjNTUDoTCEoPwR17x8NXLsXPaXYPd
z6asOEgMNLIIg0EEXu0iB+SCU3qRxZ9MSv0ZNLKzJsWeAMHWXZ4NrFqC9xNFPgKG
vzYWwXkDEvCxOzAhIVN8lkHcJDRXPmTdpRWmr6ayfmroAi2sQdlvOGlWk3HT/HWE
A/Fa45Z2Fz/XsdDXU05AhU1taok3UFx76PO3bqEJGstJHnJNBfU0p4sLlMsnXoR+
QW9LSX9FiQAhBvBsTSjNjZq4iK3FzO/gsoh8C9bx7ZZGiDjsSRgLW+a1yUuM4q1E
QxOO73KR4r7yO4lrthe3Kx96AB5xFDgyywRVAvpccRkdIbKQOUtHbmcxdcXXPRKO
VXBxz+QQcfRUm8P2XP+MdQl3eNL109fvzKtuZWshooErqrK8nXZeKuQAKji4AeQX
w2qMv24wBBVtPom1kVjPLOpLp1ctkKftgqya2tcrj78Skbo9bjprrtp0kjwvU+hV
9O/HMcvB7j7To21rvCALgkWbFZMON+0xcigjq3xL1tDpL/y5xY8P+OMz2LTqWPP9
jH23V+5jIzCAuY0BKOlfCXFxiSbg/O0XN2ebphsxCStVEaDWvqzds1eqHsbEKygz
OTkkhf8Kz4L9RdSegRuVois5027MQ16wycO9ynfLiO471NTWZ9tyI/GSPRf3caCj
HrbDBDx+0TQNUIBmzlIJiLwOENO/bK27AjL3WXS9kYx2fr4YaGI1zEork0Y9pXRc
XKzrF/FTOphjziqi0C0OZpNHicudXA5g0wzTfzN3SeXUIGz3xGeQ00OsqZxE+5di
1BUaRH+TiLyIrv1F/DakMMY5YvJNLvLWwdoYLrF6EvIBGoKkHevW1LWdAJVKxqxY
4ab1kXbqc13mZMfP+ab5JI84y7Bl6vsWIj/D0n3jPrVS5ACxNjmr4cKK0XXGZOBD
0GOVIMY+SM96Xeaj0RA6R52BVV6NBFlf3ZBeXiHESuXjtqKmbowlWtwudL1RAsWu
Ir9q7D+S0RQHxr886Ij9ODzsjlot0IfzrGhG26LYJUpOPWGtWOgeZEBSPAUX9Ip6
wzDp0f4JrFdWT6nMGhYyBU1E3rx7gDzNTOPirNimVGlyvHQB9LemgIJEjVP/eIcP
VO1rrNmQGjBQqJIx+FJwaX/+W/7SK326XOFB78VwUz9rCOarIGsN9OMxfWA98MjI
sQtG8ehiC5FCT3dcPsU435sM3i5l9UG7ixkq0T8/co+Md/wN6mCvSW5X0sEEdIbD
2X29GKVpQ+5TlxP2bLMuA9JBGawaYmfATuoosoe2S222N88tUPFoWMtNcE80JxuQ
iah2b8EF6SBMIQCTHwpEALETZ+FCH8ltYwq4txmHdwUyYn/q6i6Zi3M7PQipoUYt
LqLIiBtN7Ldnt+9TyPjlkAfpFAmHCKcYpLBxhIsx5noVHcIXpw2jIYRxWydXUzI3
LQRrA7PRMu9Y31L7DeTj/3ktXsSDqZyNQ0m3G0EkDNkoXcAqsGGPX4B966tqO5u2
cMau1fiOrjxH597HiB+G1sq9qfc9CyntnPpm0CPMeCvAkf6baRxocAwCC9KBZT73
ho8jdpkhnRmm65Q++N12XkWeflCy1ynOeeq6ZV+NJIHBcFj3CjDwPhkIfNkm48/C
IuMm+Zu81/M+lAO1iycR6K5xlUm5r7lFutM1v8i7xJw/KkbC0KnjtCdhCRCvPGRj
JGiQwiHeiA4WmYqjb3+ihAJ4Hs246H06gVoF+W7MMKsa/AyXk3GLt1hSKnHGuGlG
S3SFQTxZgv8tPGhrZ+PBuj5S0AsUa4Pg3PkbqG5xKnC1zggVhMJb5tIn+LPy6aF/
FiIDpfDM8rXvCE7ZGBVSpth4bMcqFwOIuVBBh+TmfkIkqetGyv10JznTbSPEovp3
fsZS+i+dmJZmkEl0vEo23dQOiWqn1yBPUK272wZLW1bL5QAvOK+SuiAtYjCV+9mj
wbpfOr8ln1M3o7UBb77VFZJEpBRzzvDbuXbyRAD6UJhsKDYfu9AkmSW0OL5e8z2h
E/9jwStutKe8do6QqV5Kow29NqrpauIVerivCnG5+Sn1cnCoDHG+vGHuI5WzOFOR
+wP6zvFjzVeDKXSAU6UUNTnFJ+tf3qcJ8tEqJigngCctRxsWEPeBUBQufv7tFXJh
KAb44Tk1wCuo3pQ9SIplK4UnShd5gBTKv8xLhA3foPnQXjLXetGrtby6EDuwU1BC
1a5hqBn9Ig0Hku525Sr2HZrGHnpEeKQyrHR9kxe5AALIiZ+asplG1FRFNL3ajIKj
qZCSAPA3Gfios9QxqhIQ2tTbuPqsFhjjxy2UMmiZFX3q+awFbL0d/lf+8GPwR2hr
0f/u95cnVqEXZgr0gmzKLGkvvzH7zQgQh3/UGjjKQqkGP3Mrm+Q8/5yhao0eYfVq
IBXwzEbMTL4vgewQMqW6lIUlZbAdCkVbDy6onPoaTxsPk5JZKF3uu2JxJoOAQOtO
jXwKn6V847PCl5nlM0PgYiyF4hVv1ipHnok9gyFa0iy+sKXJVA0TXWPmCJ5dNp2d
9dQbNS+GZwSFehYe/oAk/7MLf3bj9Uma5PghtaSphxxzmEl41x1xYo+DF7J8BHQ4
ztY2ftRFnfw/zRhcE+3lh9sYKG+lGW5pan1UiuhLCKwTJaryDdC3vKHuiUMUI3oK
VWlUbAF408raXGwUkqwXEIUx7ex+qATVzv5FbrV0O7jw3HHWfMFL4ufAQd3VOJPk
ahdGPwC8OY+omrJOoOdJfo5NDmaxXM7VbTwu8cfkkytkOeYocpF1llxTx+VQsIm6
fYa73JQ4d/NQV2Qa5iiiIV2eO5zA5x+g3OooXXqD+TGqN0V5t6ItkZZhpHgSvatG
GbcSnWfEWQm0vNJLYJEF+kQv+JQXoZyXTD77Fk5ydTPUqzrN6ojGKg1B4yq4cxbr
Cx5+GOCwisMaMcIbe8k8iXUOlcFSsH0sX3320hNF3OyIpJsnch7fyIXlbptqBlYe
Ctppc0A5Qawzxa3l7r10RwYQKUtARFl+e8iY5hQh4N5D+bPPKOe7pR4fB4vTk3aJ
l2a9tP32ZoqL2WTN2wJgPWQfstncQKZZ4CnPHXBUBkX+S+eGRhC4V/AXT2OR3RzF
5DbLFlN78FRMzTWqHMwpmBfrTGE4TPI44th8VeMJQ8WlSq/YUBbmv9j9TcapOteG
4BEiWjcD/hfz0EGdTO9x76HHo6rM3G+aaFpokLPqzz9DB6tKDnx+cLM5H9apG+Wj
7l5oqUlCw29eXhPDh55MnN1jEAvl6C6VRZay652NrNF0uCH5xqiEulcC8MZqcOIV
+Ufeob+sek134XfWTddtvqpQD8XBTzCyTylU1g1VNGdYSJBNz9hbEoqxC4vCXBia
j8ta6zElpxGQO3tDyKbkw87Sjvp7PZNmuMGJzpsNUuFIotQxvuJwF4e7/OClI/Uh
YMvPFO2NX/h8zvaQpWH6JjofMxr8gz5knC69U/+mmLfic9goTJvyAMxH5rhzoY8E
E3Ikulce79c4A//7fFWjxx9SUUEMN8StY/2iVMDaRDhzYxqDCIFNCl2R5ikIsdtn
R+29Sc8unicYq8iImhrKbDRyK0gyL0uqmptf0mF6kXYKzdP2dgnjEj9WvKNdaIAf
3bTKTZcVkpaph9+aHA1PoCLXTfV69Ol+/hCn8kJp11ZcS3tV449hndzm4IlauMx3
W4uy5zd4VPqSOdGOBDaX+mKMj888YCwhQR0p1YbnCjzIvdz1eFWI3kk3gjPpViab
oucT9gB/uRuNlE0LxwKbu0A9MA2Kt1ERjTb6gkEo2olk50MGMuXPkpxckxp60pyZ
SDugHEk0FAhL570/LSkUMBHmwA7JUWVEA4hJeKOXzyTczuF3cbRFs8tbxZ+HlowN
+ui/BGdUHJK1Kd9YMKPGaUV1zZB4bKwaAFTKSNsZhkvPonMmIi7IND+duexcVo+W
8xhUJrqD/plgRqwCp97A1r/xumLSO2BRC6GLa3LYmJZRwDDYagfsD0mm5tmaT1nW
teMnV/zRP8dvt8GBAm7+yESAZ6jiF6Zoa+8GZutmlrmwEd1jZkFF7BqOlB1l0kIW
hbpCUPupporqzUx1Nx038tp9L+VfYvPkePUXbGV4ILPGoBAD8rFnRpREzWYIMRZ5
VqsrmQQqaeJ4jaQld9t8gYscGDIC/eZ7o9eto0uqY0pggMPaZU8VJdLlX0SXHix9
Hp0f/Co23YuQHz8u0SJ0UO9+VEEqFyjPlNvpXMNA+vO6p7a30Asd/5prfu/RHjv1
H3it5IN6Wx0eEaGL5bbjVT3eDsqLGdrD728BDFNU3uk4ShfkbtVVfCMS+Hvv1aah
IRcFTRm3k3H1orUd0Hy8IJd05lWYI7uRU8a54G5Cdf9E14zg8t77GgbZ4Yt2HAGW
UNwsmvEUdxcVooZKjMqWIrUnJthrYa1W67WGzdf0FJvn1QIMdCC/GDUuwe+FfgQ7
L20oU/GcmLmw5mEqphQIUtlANWu/kNf2yncx+yQh5O8d0SHNtGkmVsLLxpS5mJ8f
5CKOa72p8dBdnSn5Qw3oTnFz5K7iJH5VmRYtKI/O3A0dvkBveqycpHRWrdp53r04
Wfo9Sq97tx6lB5igoY5w3OZjR43WvIJuTQF+LAApx/ITjeGIoNz4hjk3/MLgtg7Q
YISr4X7fV8ZTlgdPNYxK1L3JqLlxtsAMuVeZiIh1Do8E0Yv/l875UgyIeQbCKa2k
2KjCnAvjhwzNl+jLUMZ8cOj0EjfWoxg5KtNdTdmVHxgPeAsXKiPukOSyTA2nOnyl
Sk6vb6EdMxJg6T9b+G8Vl1xsW8WCdCwSOr7SxeMbGGyA29MDJRmAd1BD7Ek8L0le
lACJfX/qUF1M4bw+H5pPIMzy0AlA4bO3tpnw9VlZtOe23Fik7r+crtdQY1Vk48aV
afIkdcOlSNuHzmUVjKJ8ka66z7aDz9C848hiwTLGEKgSca+/MIaAn9NhVEcPerPY
fn8I6rqFztRxp/nCwai8MMwNrWZvZ9M/WTgG/fiz4apbGVaV5o3jPKHBtSnw/hk+
op+L4IbtsfAV787dUxSr6qWOIcQa8wjpyH6GCu7n7bq7d2HHpkflzwNVn2ao9SGQ
MmL4saggMTYqRwwL6Fo/ZecfVTON776b3z5vh6J7BElJkINrqoYVZyIW9T3JWtoX
IhTTVmxwkmwPvp2W6NKj2YjlVr0Cg8omf9jKrn3CPb5CifHUPqoKQ88NhaKJ2fas
1HFtR2lN7XNOuwb/Nk/34LiYnO4HVEDKl7CsAiJ+Dx4R9z471WU8/86th7F0mjZZ
tM/vZRk7qoCvReYszk7bSelEQFHQkYWEScDjXdtOj3nfGQfqnAyoWz7djai5WXXC
BjCp5CVYJfu1GRNaEYFkfAr1fPh9K00+HFi/Mtk/oZfaMzn76STl/H8/O91samxi
AoMvD+7zJU31R6I5ze7ej4Xb/F694GivTrg/BHmDWOPClFRjUIU+Nt+Iqu0AwBW6
3CMyYAbzKWFP4cqEwsx2C8+nQCMyj96w5CdmJZqlyz3NgcCkulWzatLlvW+yzQ0X
KhqlVn+YPmW7CSc18HSeeudARrhIwSBAjOfCrPxwZsIbldYYvo6mrmBYKIn7yXPQ
YJC+TyIxUbqNYZ+KAIPrf/DOCnNGx0FEowJcjFCgaB1J7iX1OhebZbri9sPt+tMY
gdLzx1Ymcz8g/qdJIs79Ydy85pNR4K6uj8YV2m5FDwM34s/nQW08kH+iZk7MqLYe
l8KTVxNtLmhjtJcId1QgME/NIn7hUwwoda6ZNP3G3ORZ+1+5KfQKdJJ4cChs6Urz
Thgx+N9je8IvG+CqCScQqw5s30BgyowIumsaWUNTvdT+ujqzrt6hjwhJ38dFxM90
tdP75G3bT6l7hINwnrz5hRp4puxt0sRuxVlPMcHK9XLdP/a1aHT3HVawsLuCfzgv
q9BbL99Hin8M5pPQsOCuWN2cekYPDd0lv8YOHKfiRr/9wygNZLgxAs1IKI2ArQl0
K9z9uDN/mmWtWSDpEuH57eHLTrJwt8c2OwSvyfqHoNjgkFPcEl1zyHZS1ouDxJaf
Frqqyjddtqpdt6/roqx+O9Zf+6SfcOvLbwLifrp4RFCS1hRl81fPcEhR+KY7d/wE
SvDjgQPVzzXWgtHpyv3Dp0sGkxb2zYePOHIYGpJkPOqhd9bhzarggdO5CfvvE1vs
L0c6FVXECwQHYsxvKqfdFHo8K+W5EaGGAYXUNv8foeQDjwHSJtkcnJ6eklS0XOVZ
GJ/4q8v0Ag3gIslZ+BTiMF65nQ1L4L+hLCfj1teWxLcFhcfJfZhcAKRkh1RarYD8
LFqy50VT86HrKzDAkR1BZYZqh+fFPab6/3itsRvDfVKNuTAiq+4GUUuG7Zbd33eU
Zfxi8Gl+B6IFcnqQlvk4B+g9QZaITXAQrfprcsyGtHwllD2RGy1ZCMErXwIC+TVm
fGae9B+fVVBfuJ1dmgB49sGnfAxJdgZN1GKoU0NTv0bBA+XmY0kiSWqtxJwZIGZg
p4fociPP24sPpeDdootjcnXQn+wbH/1x1jMAYpQ559zskALQRmQJ8JJSQVZdS9t+
PdOCzTTTq6orcnin39Go99hMwOpUQVVRhvpMVglsM5ZBpy1iBA13bcW8g6+5HOoc
ETfgWxZ+D0ErkSSU2Y47r3QqfANK1sh5YubIVwhwzMpx7T+5Gq1jg8AUbHu9Hh/U
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7824 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/T97rZhQva68T7JOm4bkq25
b4BW57ADAHEm2yg/Vzsfl9sAL1gPJW4UBYWsaJqdUHW4GN0oJEvOLjRyct40Hcqe
j1qvcABB2LR5KJfYQvTB2gz2NScV0mDulz8kGZSPWLwBX9EK3L38xLWOrK8cXeH8
H95LQZ8LOa6uJTXD3aOkuoD752T8+LeizeXvTfKMZQjHNk9m0ak7/uPT0yldhp/h
yevSHb0mD+v13+ym+CIhiAZSKy6KqJJDFIwDtowQvStDlIgUT9tJ0suX4e6gpSGz
XtW4EBo19qVSthkA0qB2XIMSLYtZxBWvgGm2WAiHW8tTZqdzYVdBToNb9f5bPp6/
H20YU5hckB1BGwkCUb+ZVwY/cEgtlUoYW7nBzTQNh0omUv9ryY4JOJzOEUpOJwl6
R6Rn0bb9n+fjxU+7lkBdS/J3f1D19wlfUOUuTC+jJNbJHNj/0/DZVcpzTCeEQtoW
LZ8Tmd0Tvklm9/Edfuio4DbnBoNrealRlmiQbpRqLOb4iV8u/mzIJ8vlAA4iFC3e
5RjGw4zWSqlCss84pWhhu4mkqwGsQsxI5f+ok6GtULZmQzSehauaWRSFXtaD4d+l
8zvImD8rnLdFdn5OViocoefRt/UqAAjB9JPDi1QVZqnL7BFQRY5CMzOBotbDTWEO
U8tn4kuAkR6p4vDuXYp0KlWF3qTVzovedq0o0e9usEhe9Ix3KKdaJrrZsSh/5J2q
O/x8HiQGOnC+Vy+ql0iQleWNc9XE7/Mfz35VrEm9d2SyV/EwIcBv7Dtp3pAbXZiQ
T0e16lkINQZpgqiTBszUjrKtnyR+rXsYPc7yEq3tXMD3dw+KvXYkERWBE96T1k6J
RGb2JGGzOndRxaYSjUHSmruZ8ByVS7toIF3BkvbblckgpDSGOGxk3bOqm86glyxx
dj+IA/a5HUgBMiyvRcBdbG6J4mJ/RN+s5WORPV8lOJ3vUfylheKrULRvSsxQBrRm
NbP5BMLtbAgJxclp5ovpmXluiXqDLDms5YFHCbvmJ5WLdDjC1r2V2/apUeCqQoI+
hbDKvj1RUhd8rf488wYP+gy4KOsb4SQ10g+PqHXmdHkx2NkBk9UQANG0WiCWQ+A5
39hWAFYYqH/RVosv2iETIK+sBG68jbOb59Sun6ixFtXE+P1cLqloWAzE0o6xkyNy
RAzaIQW2DeSDST4n66nzIfpp8OIrVfKF02h0gciSRmW4DgXgC/9x6zKM0eF/i0T2
xM1ra3kED+Zhg47ixFvDNCPMFXNjVMYins8H9kyC/dLyeaBmRZrhMzxhYBt5rSZO
Ye4CDdaBDRk3lpHMWFchg2OB6RrVVWtxy1xzxkJsHjap7433ncuXAlWJg31v8KNX
0XIGmYJ+j9070Ye3dP6i5m05sEVKFs98/ubcMztinBf3R8GO2mvoGGc4348J5s08
7u/x7eVqrQrQUgzj+J83p2xngwx4BL+rWOHqGFYpd0bqeBKCK0TsPCsjSRdiF8no
d5JFhdbuafhJZ2EbQUqkXdEG6N5AUolBPWqwE7l9bbkJCpMf3Y/5ulk5mxmCR85x
eF2Z6fFRAM2cnQM5gs+3n4v6Gj9zreUu2H/Ah85BmDJH8t8wINTk/4Yuz8o0uaRN
vIj8joxpfFOC0bhi3x+ef6QI1hqjTz077JRQPvkGjEUySrJg12M/jgJa0hSaNXGT
6OIcqVsH6mtE46PBI3obVdBdpzBvfsSKK/TMvMBluYGEQVFXWK71pzcaGJMKAxXm
IgqGdzDbvPY8yKtdbs+ZVGXAJGIG/lARbIxjtgjhNvrsABp30Fb9RMdRh6ntVXD/
MoByeb+xi4VKRWAwrFK5Kd0EXZAXFGavrawl5sK7wT23yPnGBttMh4XfiTVD5P8r
FVMy33sgb6Ss9uisXSziYNmX9XnXq4Fo2PisZ2CfpV3qSR/PoBH2cvZwIJZ8i7sc
BYXwVterpNueGf/i9/+RQC+cB6OLfqfMAl4NIKxGFsxttWmTN6X0k1/+0CCvu6+4
kwiF5oFuYmluCvL85K9T13SPsB7F289YFSgNOWUjPO4DQZ/7Fwf0iQcQ1iSwSIEx
6mL5Z0Ky1/KU88/e2jpYGvl/+/5tX4tuXpwjoixQ7VPtLawjo1uIQAi59S2fH1nd
N21SoV2s8YLYfWNyuOhTQnyXVIbjsGIOt8CP0FDKv336WlJ/57K6yURvE4H3YPYN
RWW60wz1gZ8boAR9KubOpnWCV8eUuGFm/1VZpK7fLHq511aC12Dmlw0qGLCFiWGn
i/7ynQs/asfME4EW97sMmdRcp+5KuV1S0vkqBIlufY8yTw2wAi+KSTxxgQsJOn83
dw2i0yGy9KLuHu2zxnTfSQ9Ss0QZR8Ff/NlVtQ7df+YxGAhJEoXJxh0DeyUJdlTF
zJx/OFRc+8WxaD0Z+Olq3/S/VuR3Fxhf0ZaWnHyuVT4+agosFVf5eTCuU3C+a+p/
nzgDNHaIIui6u8bLoqf0tiyADl9pUiKz8xzRDRGuV1JS3ixBrc1RCsvXHRrPZgl8
NF2Z8sXnLy8I50MSFPDtZSWbu+SZGfoIp8LQPRD6U4iGB+FMbBgW9rS6x72eUFgs
ZIzfkJlsnJ2Q8ENZWPmHRYKW9ciC0P/Vz4wMR+D+WsAbfjTHv2FYv6rcya/dtZjk
nGTolvK+jecC+xfWlDl/grAzMHr0xq/pI8qy2JjhCFKUxD42t0FJ7Gd47HtNG8ZH
GEQpbVGKsJqWNPQ2KU2kwQigWGGAe50zYErPS3E9SAYRK5IMV7PWjKT7W/Y4hyjd
kn5PVumEJp3ToKhGHLQqgRjk0KlraHcplAY1+tReGRqviB8tkT69ad6XFSBAPuar
cNn/CWUu4vTuGxZ8oPBcXjvCM07aejcEl0YEi55fsdfG4BVldpzSJwfWyPRqiUGz
oB2yMDswf7dF2gN+Zz+ASy2LKFJfJCIazjvhiF8whN6NF4kKYLW9zA9s+Q8puWgZ
EjmA6a4OTSfI2lFkEMvtMjl/BgUnUvLlrvzZYvh26wN8WPxVKcVt9kw+twUNWC/0
jj+hOP06nLaarr9FFQmT2RH3tD8ASHSYF96Gy5OEDqlWUsN4XDYITteA4YrIsgqN
THFw/wrg78EwxatorFU7kw6y02Iqw6G3dsObEclJ01xtDnsMmPjmMeQzaPxXhIE1
YfPPl35y5UMZTSAEptlK0d1nB7Ljj5PAIQtaiX/nimGgX8lp1DsqzAbUOVyMlhdQ
M28uBLkrlCYoOByGobhMhvl+VaFOq4Og9yjsO4uFHQ0nGWoLURIAroMvR6LgfPz1
luFsWQB9shn9lvsxMXyZQDvtXJpjFFZjou0VcPq9fQzRQif2ra5/TkM/SrLLPMXT
bcfYwDDfueWor73dYLVpsBBVU9TbMco6jxu2MbSJI2hSVtlr3sbEGrXCEQYxEh4v
FPpaP6Qot3CzhQnp0qZNerA/WscaBN6Blo8Y0knJlNwAFw6+Rm0IU6m2Rd0P/u0S
Ya20gt87JbLhvPQn0s+8v+/Asodx784zaS7GSzZeptcFqJMx3BPj1hfCjBcciC27
nUP8cD5Ptj7g2dZ+ABJiH0ugG8QH4H7f3O4mcCcEIra+pAFjv365p3m5XMkGcOXe
fGbQ22BF5bAsxv2tVZkxD378jkPbI43tJKSyLqptOPH2TFQ3mPi/rLAKjMsAzHA/
cWgAKFmcJfcsz2suMGqupDTOUuKs7Y3ojvfYfS7U58LME6Na54d8jqmq8yIaINZm
thQab+TagAYhFmw5YEfX4V89SCk/hOa6mDzWi/vOALHsaNfROVfqqa8gC+MTutMn
C250E+KtWg+w6HygIdbS4o/pJiVEn/Jf1XwQ8Kqoa9BJoFPGDRJz/KvVLMXuqRM7
J+a/uVooG3U/gOuSkn5RQBvCBaYMT4gi+6ITKsKpq1GTq1w13dMc2/dx7ixyLWi7
dlImvtWfPrTsl2zDTf77uvL+oCozD0ThLV7m2vghn4E1RQ9QtLopciAqPPRbcEY6
5sIZrFY09Fo7bIWg0T7zbbegQBj2T+gudAzedzTrIRonxFcZgjQJmaOJzBohbbVA
XswNOY+QIrrO0Vcvv2Y7wiukfXta2JN7IUgsyTEy+uZjFsuTd4+FdEasFJknNfMp
bdxUqqudpWOIWehw8W496vGxn3taPKx+YONpXLVuTUfG0fzuWesIrjN7L86Gb6nL
JRPdn2BaIUX9sJ4RQHWl3gr/KljfB8o7KBiv14YJIDYBN2CZ58+WndIGqAVVpxwn
XWyCWwJbepLrc0vZEgDUeMa6+uHjnCcESmBcDB8IoUV/Bz9k/4P9J4XCtidcr93l
Xd4WNhiduUQlGO8TpVSd2xam2n9MYRDbjkeHmgAyqEJKo+XeTtttSFyMhH18le0n
KRhdcokWS7glcpqD886G09R7exkRmmgzflPdoKA9CdBPKQs5ltOW0elPZnLyKn2X
A1pEZPUUmdcWLSY/hZYVulqUMQJ5dk7yXtUqTervKVla9FYYKnEQRH+h/xDj42IE
HFbdvkZMDeMh4K2qwORmbeviW06hxkIa+dwbS5R+U9SaQEjdAbhccJGrlfDRJtCJ
DRgl0b541D6jLiVjlaPMEWZ+n2uDh0Zq1eg/cK3AestsvzcCMmVgkBE8YxsL5Mbg
6JzlzrLX6ftFZPv9XeOpG6MSrMAxJ3bAIThgyRpQFlzYyRdO8IozMGFE+6U3wKtZ
kBSWKUn6FChBT3jdcsfX9Q66+7IPZazlTi94NXwUJxcWj6OdE9yoTP5dDYv1Y/9C
4WPIEeGQIQ9WgmfxpaJr4ZsOLAdVRwA34zlI5yaCd8QDNjbqMRC4Tzh7X3S3L/4b
9lIiTGzme4fXpGo9BJ9yNOA4B/WagUR5WLIbrkK0qH1ZXzNXQqofS6tbyzFGCQAb
uV2SQK3mAFpQdeGo+maut0OV0IRapUndV5j6J5MkGwa6D7QxaDK+zdjrmIzIQOVD
fDgtZ5tLPkl9I4ncOZ2y33NydpIgwSHF7SmuFmelKqqa/EarDvjVn/0JLaktM8+c
GboRLarYhYyMijO6o6qA8J+A0I5WmkNrJOGMUY0verkbcxSwT+D/0HzA3PDK1hHO
mu9jqPRBHCPlQQZOHMrI0sBEScI7oR3kJmlJpz/LnzJBmf4BgW/yvasYa5zBM3k8
z5cgfL8I6WbIbG3FyOaqVa72v1e7BdLYmxvuSSoobzclNS7zXup/vgj+yD+pcNMd
nQCPWJ/hOjvGLgnZjamAArTxMKeYgeN9a0gOgGQeHKgcj6OOxwEdZwy7UqUihPG1
GrmVZDO0u5lA8zyAv90Djgt8x3e700yzk67vlQyXshANXVz1Ez+J51NGZBPbuyz7
kjlZH7TETFvd3YD0NhxHCeFZy9G77GN2zKFl38nInF79Q6ca6liPasKCoIfPisSo
pscIuKI+ntjKYky1lpnoL1nJgSjSIkOpQdxQ5EDNOJyPY/SXu423DiCnVxNEpXdh
0b4s8BpqRO0wdmysu+V22ZhcDz5FYIESmEwpgFwGcdBwPDke/qHRd54pQEdpcjxS
KZcQCnRMZTz1OiZtyts2Q55ca2w8P0ViuiZqocuLVcxi/JdduovVYaveVNRJ6KEh
9LhKUPHF52EuCpp8o7W2NB9EoZr3p0uSut5W9z10I1EU16rgAFn0kG5NSHKDRGvz
6Y3Kp4bNY0W1DGp3gnvLIybxyNIniakcDHhLPASthCPfx78ZmveE/r2UOJLasMoH
74bQ3JzeyObNOGlkkbxcp8N1Eu7QOB99PDOsv1aUPkIVsxzFa6Nhi6aLvK4NMoyD
hAQd8ne4r3ClyI6W0TTlDo6dnZGvvyzbJF83A6jd/eShb93V3hxODeMipBwIDanw
wOfU8CFgaRXhQv/PZ8E3O/XPqOwdEnbs+3vCXI9ZQJNBbtJ863q6hGkPMFkFb2Vi
J1t8BLsu3vGKYFP0zNKQ35WNMZhwMeHh7XUDbAvEUPcDbH2BrURmAfObiHw97d7O
yf8aQfq9nmb2UPuF5d11hHtvCPn7iCVMyPmJXvEMR2uEre506a9Rd86eiKWDw+GA
PcOOyZbq/cPLadrYbLXakyEPw7nf6EiAZAri6wiH/PHJfKBjyxsASfLyRvfFUvZD
xmjGMgtndc2tnMHZvQRtKe6jAwoyz0womzmy4bDQGU+9sbeMcSb5LMqR4C30Y/oj
w6xwGv7YmRFYoEH61hpeWTED7dO61Q243EpXuMvTIkTXstXvfSeNvjbKKXZJ0cfn
s15J1fMujWJk5YtjA8Uc4i3jbt+H7WUgKyIiUxcK7oLlekx9tggY0U+SLPE/htAq
vIoiUEYs4iD7f7J4RKtsyog+b71CTKOUsRWffEDZnqSfsNWqBpCepkUtY4/7LPSe
3JJT8YrHjqHSQH/miPlsQQll2B1e9/5+HODxtJZm3i5PQxAwU1XbXNIdCwAosrgF
VtTLJIxWRKyjNK4j12V+9XmhG4x8ZYVPoG5OsLpn7r0VU/g61kDygqJKxFj1kc4a
kBAVBu77gh3edJWQL26P+wTgkTBkLpHs+75qgLiKHUEuKL/eoeW/oEf8GFv+Q4Ei
MHEOlS2a9FwSIBKYg30io46JngIExL/Qnag7oHgFBOLVePZN5Air36n6YQ2nNLWE
zuBxaCzo4n6xepSktIPoz2ISmV4wdGR4d1OBB9AnKFOERoxhojRbtoI0BM4wCPt2
eW3kP/EwzaQYTGbyVvvYbJGrbI5U0MAJaRDlWCLc4ErF3U9Lv2p57/qK+1VveYZs
TBRmwMEt0VfPYodNhPI0ThCur7gn7k6o+NERe0F+miSFHquU4ResIjJXJnT1/bqi
YTGs1k3WtXAOlgWbHvVMOUN+wT3KkCl0BB8c+BWSc3rMCZiplPe59n3FxqOexsue
wtbOaGKQdJgsPj+YnVLBhifH36MmU8P9slwixH006xAO8W3bFh7invDED69THe1L
L1zrAQQiUKs4AMGZ3CpJcx+PYnYrwlZd7feKDYVFwXiydWGzhf/QotqqHQpOMON3
IjF/noFKhKaBkpkjXK59OqnyHW3jbkpcL4HiUJIVrtzCNhqn9VF5ALx67kYrPfqB
/iE//ounMbiuUhiWEo+7/cwhk/lASsXC3YrRpyG+nAZooxoOMUUeGzt10ywEg+sG
NYq/pH0f6nkXfDiVMn/2TFr2evUjGFLjYf1wKsUBnEwY608OKO9ZJSx3rTtvXqbm
cWIRcN2xrNguDUnqbIRO49OoIl3jWW1aqhllw40P0ou6eykAxzoMssnpxzi2DqEd
N30XJyi1HW8sjnbgTU0eqG4ogMlSghnbY646qalH2bn0kxNJUZq8GwOpArjJ5Rsw
nsSCJBpzRtm4f2u2614PLm6fk++RwtXS7C+/igLE934lDNPvmwbDTO3XV6Ug7OVy
rfc6JXa5YkasD7rXmrOFG5hbBM7bOj7wdjEacH33df+VTBdpWATUVKGVSCU8A4tM
GB2iO91rhJhSqtxD2idZdTxu3mpzgexJqj0RPpJICimxxvXv6eO79MADg++l8jPW
BECcz1POtheJHZPS++SP1RWPYeQ/OM8XNM3xOO5cnWs5IWYUJMJdYr4Yd/Vu5cBA
vsvoZGICi2NlgQwgJBdomgKn/+pgOdYzKDAA9ou8jHR26dV5JW9FZrzknixla177
FW0P772hDC0X6EI+/Qs4FeWRVpAThwZ6/Tc+21BNvVAFr8uep1iKsA7F++dDYg64
vQ1acqTgBrdLolbFmS9XElNrLFpLacmo5RmQ54Pwbg9ADTkvyPk7Y9Hnwg87+JIk
sn5bQXkkgseODAAWuvyZvRTqAX87waZnZxja2xxG85ZYwF6aRqqRmZhuibijvon5
KrMYO5BmmyOTrl0nkWijy3RoN2mmXE0tSIA0P9IZxMVUvOaL9EibPdWMC6JO7WXJ
FO9KE234BtFLvDdExbp9zA+MzbejxjOdS2ICaxxwSQQ1SYLma5P4cDdd8VgXSVRw
yDc/4ddiAwkIKovqNCwpx1MaQF5wQIJX4ycsCa2w3G/Rp9ruxd9SyrRz73yUV2Vs
Eqy6/QueAE8z4C2ipnwznZXvw88JWfGtPc1u0ugnJ+lrG7adBbszbJTDuurW6g2D
3PO53AbisEBkIJdedXJ+ppjqKArSNnX+nB4ebFm4Ons0XvYPmMcD7QbLFy2nCT3c
tNH70aI0qJnGPkjg8nfWYT70PmlCFJGNsg9gEhRRUFIuqr+hbc0V+Tlp9eQY8XSo
ct1YyKewODIyu8IaCZG/vcHQs2ejicz3yG4NaaILbsP9Nc8ltRJTgWE/0DfAfEi9
GXA5x+f0tRojJj2GhPEGvcLoiX+D4ee3hJdAmv4Kd0puDq6J9n4JbCUfR/IYWQvj
rS3hTeWKY2pdtVOFMMt9hAMtNmAcwB8sFbmSJ8SedPEuh2qILZfqSdpE+UgEt0a2
jwB42YE5XV1gFGeNfSNbRZpWpFWtnrymoUchNrIYVmWbG5S/rHIWl/16KFVA8eM8
zk/Tfx165q2ZhKhROevQUL19nRCbVqPLwand7UDCc+gV1966NhJNhdDCbzA4AP65
nYCxlOaDTZ9pa5H+JTfIKmlqsjVp+mhjw6/Sgf9Rdu6gNLVjk87KV3R34upW115N
LdHZ1lYGEu+d1mF1HDJw+lX9+JVOzt6BXk7eecmNCQS6INCHU91Hxpvsr1I6BVSW
a3T2adOnWmnIf4R5DXt70kCggpIcSWOjO8H03qGCIfltUUhVmdWfPk5LYXzIppVa
fU2GQPnG3BXTI3+AlHvdzF69UT/qV8U/jKqmWZUkHOGOrQj1CToHhT4ZiZI0Rllj
Ju3ncq8Reb/WiLszsekznL/DoFM+lf53isQw05N+h/N4IhXUkQt/KV+0hjSE6ohw
JItGwPUU9N1/I8xVV7AXFn8Y3uYJ+4CDzxwG/B6NQ40BGyUE+mhLwCURUd6np2PZ
sCwdNzWPqEXIAaqnINuZ+bwuXrterbJcAF714d8wgkZ0YgNqizR2V51xVIua/EA/
ePktrtwzbR4HhbDp5NQ7E10XRMAsfjj7N1DHUK5kT5OF4jxOAvcOdro4hEtPaVa0
ehm91y1JkltpQ1v3HpMPM6QHZFzwCxXbYwK+3503Kgt6wDJ8JkfSXj+bT9dH3IOa
3pCABIFRGtn9rIRyiRcJrIY0NRv4SrXVrS92/4UcHeQh1jCEMIz/CW/VGxJS2qqG
2fH1b1LBeO3hQuSZZZotRPvLMohW3lKWWR2oqkAssQVBHsGQB1HzRzPOxAtGASQ+
xkwp7Os+dhdRRY5f+QBKrCSGjLTgLElwkchZW0z7r0XOGZ2ygp19m9TMTmzTP+mq
f8giE1DohW8EY4uBEvuqfEMHmaSKvTM3AsCEbS0+d375nhiqHstDUsytoe6wc5/a
zl6UXCXczY/hp/iBH6JIS8X+lY7EtqTJLfBK2w+HCVFnBXq+/2UKxGYJiwGO6sPM
t52q4FQcRtQNfwBDxl3/KPwb9MrTwJr551dXsUjJQ0UljWXEYLQFex5gJ6bG/fkp
dbQqsoewuRJft7Dkl+gyMQNWWRk4TOWfOvlNGAl2sZnF5O2gQ5eht0t0tB8YNXJW
QnynQQ0iIx3NjQl+5AmJwXiE0OhGsqgpSZd6SCjtQNQKaNET9WEjpiHskQfS1ANa
bAtiZKa9k2d6dQJBD5uxyFCJ0rghfEtsEPWei4PX6jADMrnRK5CkjRq7LMRT4tf1
l1IGvDwJ62fdeZ5vU3GbFBl4lGFBOR9BfiLJz+WJdAaU9Z4luEUDopGkZMfTXpbK
cQRJdiHyrwNGPKMH+uQgTmRP+7+XhU7VE+4KFKvaw9HUJbhGezotcpRpXeqdYNME
WHG/ZvTFleF2y3Lzlz5AxMN77ibxdN/5D6Yeh8EnN+W1/K1napZ53MQsZuGPMLwu
0oC8nYskm/Y5qRxhz3vt589vpMnXWnVvvfi1u8cHk7Y/x75XN7JX4k9wsaAxCGmw
gk9YMhaveajAVfdEW72uCbch6UL6zwTXOtZ0HFaqdg3jTkbCHXkOOtK+J1bv/9LJ
f7JwTIvwCrI7WZhisx483Q9n7N1YG+Ptez0UV8304oH+fqp7Qe7P5gcJx8SnboVS
w6HiWzvMtbn/PFMQ0tORDosRISK7YYOD2BxLhk2YxsAExsvbmhyoO948AKz7sCD+
tLb65MbtTgCr9Uc0WT2SefqH1mkZJaJVvAyomUVN4qTxvRT9PhvuNH3OIQ/HKTgQ
HCEh89O9sTVX1cnAdlIuLAJUNydJO2nriVi9CABBxWhPEc+zXv2/qMan0XrhMOtA
14IXkm55tuZj68QDmVwD8guxgqyIzyuwo8lQ72gdMX83NwnQJAZukY85vNjzEJeI
>>>>>>> main
`protect end_protected