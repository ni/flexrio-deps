`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36768 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
yB5UT5oQgw999PzwDg9vEoKepf2TPySHYDB2dakMAbkHbKVLlbau/xbQTdPquu8w
npOYJGYk8RBD2wez6cwFcKcRi86ughQp1L+s4uaoYdR+2+22lBh0h3oM36naLYAb
/ZxyGMBhOi3lGHP0a4gXIhx0KJHDxb63PvLHemgNYr52TDzkVyWYNfNd+TTgNV54
b2JNa9FEnDbbH6jFLtti+oQU90B/fpTTF+G0J5RFU+Lxijhs6MaIRoDd91EsgWAh
7gfMZGWussJqEP35ikb2kf+HYdse0L2ZI2Mcx2vhwdTZ+cD/uBf4msFKl0Hyj/mh
8JiSvJlcM4oaPrbaeY938aSFw86aH0fGhINlW0JluH86HjWUi8ixUYgPa5PU5I8w
zjjNXD+/+ITM/TFKiuWlCFyoExqjOPR8coMt0dIck4f/yivoDXSBQ9FZN3CMwT9+
g5/gH2ghELB17k2eKAWOyTHEevtQj4vCOGwQ955mD2cppxo6PxTG+El89ArqoDez
W2+U5S5pmgH1+LS5fFh65sqvZ7SkwVxme09GGa0Fi6ViuAAP6V4D4JXm0vA1fHcQ
QgGTTMkfQ7k5+Bbld+HqSkLsAAXsxpZlAYlbLUZMaCox9vn4y7894n3plFIy/m43
PzFRRxwS1dlqul+PQKl1Z6QxrNsLRM1Fvu6KD7X0CoHHjSOPzBvrLgK1d6UZaHpM
1OUnt39WCOpvUGq+eHWruqFbRbATjGjcVACmTQhB03nQPkYCEitWYUzVrwBvSiik
sfQPjuIYPKtEBtYb1NK6Hbpd+TBjKdPisQoJVAo7CALIHrA4TCCzTuCs5ntaxamr
Hjmile3UjpCUaZlMY69x53RWsd+fbs6lKzd0OwFHFvhmxtUZ+ze+oklZxxEBnpsU
QNiedgP5kijPm8gujxn/7UNXuXi5+la2fC5FYb7pr8fXNoZEaGNJV6dHmZO78pFs
LMlcswa9pF2TGInmoLXZNUOJyZ5v7nh0CQOmphB7Cw2q/CX5qpA6f+0Pqfih/ADJ
9BUYN1L1at5WZXhIIZTUyxQykY/dxjmXdpBWIBi6PV+ggdIzh+Sl0i7pMAuM9Dye
VgqyzCoQchGQRLt4e2WBJTkRY10QHf3ZHdHoACjH4EAOK4wwmKnGDme3rE/oPcpl
murCa3MHiyVJ3uGocC0FAy0XLKjtJC3vGEGEVvccrY1Veu8uQaFNRDJualttQdmX
Y0wGgrK95eQkvhwffWQcnBaMBGy0SyuYj9Sx2q+1Cxo8GGcypaTCHAX/rXtmZfgc
A8+GMGjV/LBYQgSrQgvs/YJ6h8gBjU6QzfFcaqQXJYjtBeCg6OtVV9J0tGhkT/md
HBZ0AZOTeiXLhsz5FS5yqn7X9m2UxKgcnsv4T8lszSfImTj3rii58dbtKsTal+Lc
Q/aush4wWzypV0hFAGKuCAYsEZEtZ4le68BhGskBse/b1AwMzOW1Ro3sF8zaMXzv
AkAhM2S1Wf04Yb2NW3vBgr1f7yVkNd6b4wqO192H18tVKoiso1dfUrfXgt/zMc7z
FoRmOfryPjvIF7vQR11469YCpd81sbISTNl4aWR4n/g2awzqVLlmqMDlkeg4z+b3
brYBh5xbmI7ddWMCkieD2rOpQL6lGX21yb/DP1uFzlgkb1/IdNOd2ktd6BrXA4GH
RqTxMpXima8PWVjTgkBsLEH3Or/s29hhteqSST6MS+J6Xw7a+2Jx/9IvtRhXHuqT
StFcDNUBcJTB8Ytnwc6usmBDJbKarG1CB89rSM6C7Ahx/D+inBvqWhv0T0sROiav
/pJfENfEz22QI+TWMLxNK+YSZ1n7CY6VremHXvBrFoHLqiCqmDpd9FsFt/L0Pa0z
sOaJ/FEAlqJU3Rw2tu9QQXEXDQHq6p5rOj++7n8kekcKDeSPVdjfSTWCJ/4KnqlT
TG+WdPyfA+0+qCn1ivorvFiSRRMTx4487fvTKBzp2bufLtNHnlq6hFcPLsYegTwF
k+KvnGkEgL3tLSMUafjV7nPhR43cduvBH1O64dOg8YFugkyvrXkipz9HsM51gFI8
485RL82T9np0ttt/yztx/u0IflC5i/4K3LifpGbr5ZFvOmePBwV7JgJ+U/fWLV8X
oUiNg8IA0rkS2qt2eG1zeBkIfc+4VNVDENkfWl/3H11kI929WPJmZlxCpktoKlfy
bOztfxoj7xQ2hx7HnSMmRsJjEdHAJ3nuG1Ok+e1YnEUQVre4PB9tkAocR3t4eM3Q
iRLb8me8C3654UpaG3Hi+EjVDrMNGs07CgZcaLtLdkIkOheqD/nyCLg5PzL8Bjee
JXLBX9VDaMQ+MNVHXheAoWHTADwQBo5IUDWwVttcciW9ttZy2oXbsImCskOerd6A
/lncJSYEGSt4kCyNy3ZbRsUeRW+aneZYbdUi0TKRIBLN5zqoQKO6ZKCg0j80tL8H
02/FgUhb+h9D35YEcbTjJsuifbMga+GXN/jF01lrG4CbYrL3yg+xset0Idu9s76R
QyUwz9VTpTmT7hwalXHEmHJxPXq+KpNbA7a28/gQGiGPLRqnySbNOuKeiJqhSPHq
UIY6Mkjajpy2a+qBzLXyQvmFlIDKC9q4nsi3zwKIUjh8X1WmofmX4kxPaETUwhs1
hltQFmGXDnsCKwbOKsV7++vAUM8ch8bGEyBJYOiQfK81utg4eeceLZkeC3rq51AJ
LKhE52evVyrV+lyAoPirPFBdCjVaXUudrPGht25xYPAwXeIUWzcbq2h50haAo0Ic
9z4zyYiHfo9FW7zP8nBznJC3d0z1oW5ZDQDraOZIpp/J2kmFtBIa4PVJykQa04Bf
sh6FEDXNajInz0Yueq0/lehQcnHAQrUf476CluGDbJCGwPOjT6KwU7HVSTSqgDQx
HGPrdhGPEsp3g6cRo82l+qcM4tPv7cOc7aWoDGygJ7gmrHGEonkHPjWnFRjWZwR/
UKyzWHbV5+Xpu7NAOUDQoYXMWwEtRaH7hjpvqT4IS0R8KDGQYiGKeBJANfJvkiYA
vhPRUJUERvVoFP6ZsqanIoIPYOvd8ukSg9KlxVqZgw5RADDtP66NajOWv5QwDCAm
0ftKjWfKAz/+c3dcQZKjAE9qOc5xR3P8DOttE45fXs9YsgiQvjkINRThZN98QKZR
6jNeB55JLPgUcfhEupyVkOZHbQyK+yde7vLx+onAVj4OwQHNMknt8R6SRZeqRQph
I5hjwjbOUNkAB0UFzxuy6hx+KTCVxPHWiShGAHrCdKfD7XEtsuIJ9pVrQXQw0ViM
gug0NGf1QUbrgdD/+HkXHVLHVNK2BSRASznDnbI/9O1QdqwidNfNiRtBnXC4U0BV
GvIaEqLgCMGYXIjUKwgUtod7G90n/Qg89fT+jQSSvY4ChazSc2If0/VO/HEoloav
NezMIuoEZsL2gm+gcOZUXEWYGmyLWu5DbfxiORNtSi/jEcoRoJl7v1ZNpr2nkmOk
Xc5u3mC9JYYfOqUxUwhixI4X97Lb98m673eWKLv1hsWav7FnK51plbHYw0T+wZ77
QLgrtrEL5rKD9eSDny8xeQcY/hK+/JIr3jTkPL47VbK0dB8QVJImygQIG8XHj92k
7lZ1xbUtnSgFu1/JzalLK8fMTYf++s5uTb+lOm9DHhAnzzzho1mTVAg3xCvJabmM
y87wIkOTc41ZniYbPDndSgAMPvGFo0QuV3ukT1Di94/YfjY1KDqxCoS2O+oCD8Cu
/VJoz7lZX+Jdz/ZB53IojxGw12NyE4ZKNLMT6WV+yIk6cGvpKzjkA0kd3S3Sj7Sj
jdkIbf908eZO4U/3NEuxjYdZ0hJb5CexH9z05/raIZC9rwqba3ks9Wk3/fouNfvg
XT4KRr7HvGECSJAmXQDhCg/+CHxuojLaYKjj0QFEeO656D/La81DdQ4urQi89KE0
xnnHrjtrOdtly2mVFuCqQyRlT4qaN+W3kZyOaN0KG49UQsJ8003X6Wjs+7xIZxWr
vs0sPg9V2rB5gYt8DDdPZSV2pVM8+C5Uzbdo1phcvyRcUKmrnE0Vn7l4VCxXanQf
wOjyf1yoDObhqlE4M3g2kbI0eX/mwNSYTeov7q2++vL2GjgheGsa6he1Uptvbp/i
SWIIW+86StJ5wrcPuCo4sTNJJP1tmipAhMsjxSPWLsEwaaMgKTeGdPcHNxFd8j71
B8Ids1u0dWPC97ImZPm03szRh5vPzagSwtSBd4phGvReUjPmq4Wi77nt8/scADtS
moh++UCdurlcx3NKJtFkfYGsYH5vtbB6A9LKqHypmgHti7cqM2wafmXM2wHgacfZ
G4KsW5vA0HdTdwnDMhFfwnKxtk1aWvUD0cATvtmPV1rfw4cN7ujWXCH067Ch8LnT
p36wmG9tdN6ei7DFiIJm6ADCEfo4xmmAPyZPb5U07wD4/4XTuSb8sj5jwQO5NfFe
AunUFacLutEceXg3YihetlOeZl1oZ8IHUF6sM8v/CVhx3yWg3/rsCvWh65XzPWCo
tSyXnhZiWa07ErCeWTD+9gY+9Rit1cN4WkHfL2JwIFdkNrc3O1Y/NEs9uqTIDrkA
LfSHWqAmsZExq1WfPiEupd+IJxxwUZGiqGKFb1WgOCrcO85pzFHihuzEuqMSN3m2
+CjhsakZTe5PtX/19NuJcWzInhSNVbwp5O0T5uqSEGlEa2GzCkdRBpwFrY4quomK
xGNGUFsADfn44JcSZxP3+Oi3xNJPAz+4oFmKruFV+1DsHv1NmtZj4dJPsB4pAVyr
BuHeQiITnovVbaK+SyGxQm+pf9yTPiPIJKaDlLRV2ZNgUxHPFWsK/RYYR47BNZJU
JRzA2HDbGapvQmuZyBwbojExGg6GpMgdVPwbdK7Tp5gUge3L2o4p8tRW6omA5NHD
L48cI7IOay2F+EitVF0h5Mw7mKuQAejKuATk1FY5cMYE5SeazgFrZ2HDPiTbAY/J
ahAOk7212n0tT9nV0LGYrOL78Nf23KoI68IP4by4ZlxxScVc02rL+5q+xi0Ly3X3
FSOiCvtyfLeVzKTf8Do+TNs+JI+ndXT+5NCLYcuFnYryMF9Z/TmtmHAr0XxNc68x
W9adrWWekC1pvKNT9PkehMmtWm/A3jQtg/dw4RXRgH02ydJ+0HiXNyBDnxpyvkh7
Q7YRbw2OIkyYlorc/Pmsv9boq0UMsBwh+cyBPcKJUeE3ljzx0t7GQyfThDa6q8eh
H2tYtZQLxSR58th2ewASkVmpfJlb9/AEzzRJdTBvDiYYp67Pxv8PuEWy5zpj8yGs
tTaHvBPrxOzbY1lEmB2egmbV86Vt7XcIMpgmyTe6JD3WvSveW8YwUx4gO1uZRCER
4J+MFIjq6w8whOzsdWyboZzJZxc+sTR2lKVFawJjlUVxqASjZy8huS6cxW29XcP6
MjluICJ1yh2KS5St70lLaVNiyoOJhVgagi+4mNkVyPRFa8pml2UAIdIEHKxBcyS4
l6qSYi6QJfq2gePFveSXH08oCdPXpdOSgi6eKINSX9q98+GKhfSHE7YUgoHs/M2+
zOA55X5KkAUqtv3/jHS7INbASzFos7gM96u2ovcMn+VDswCnMICZDMp2BGZV2Dsm
VxHpKtxSF0xPHV60XZIJWp68MhXOUKY5J8BMm0cASdw0TylpoInVOUSSAkURvg70
hLmZGKPyi35BmgZy6vk1A20WjeVttQyMF4DEa8UXShVROao9OddicWujbhr0acL1
kJNu9Al8wJZdYPy5lzmQuoxUyNDfAHYL0+LU23tdMcNJ3TevLNWyTLNykB3oDaGm
D/5T5tBzb6k8m9n4l5Ge/5c8bU3fJaFlNwQYVBcSpDvp8cZWF+5M9N1+qJoUmR7a
vy9wfD95kB6TnwJCkwCNcmvU8+uyyfAhq5mNa6V47IHCwaGK2bDkwAR2YMRO6rQD
HOz3hETxUBaz2xwHIErS4OHTX9VITURYJdEDaJ/66aVSpw/iP0MfV1iZZFRrCxYg
sZOg39xf6jrvTuBdecfb6gpRjInAYeT/IYRu7c4A/VEaHiX0BlWHa9v8FTzgx5hq
ie+ny2E9NyzvPzAsVfhi0vdLsL6A7+wel4nBvRCqJDLfEBtgvOw7+1ogrn6R5ONJ
ISVx1mgiw9k4+qr3shaJWeAmV438S/WWnfhunTEmezb6wpbPK1iXjhLuz4IeRlD+
H6pjxxAEgtk0RtD1TH7uE/unS7f0FL7+pw1VkIYe2Zu+vXlK+ZgTWRVbDyon53bk
3ZADqBu/JDC6WNRJt8iPWhLHpm+5qku9e0UdMaR/Z7DfkGyM55FHLgvtAlpVAcxA
FfnLS6/eUimSqYHbogbbDxxV/25O6ydx9xtQxTmNqljkN/985uYUQXAo0uLvXfyI
Cc7Gf7+TBy6lSdPiMwzdASaBGR/buWtUrBHqhZLoFnp8nmfyPeIWSyXIK8zjzBXa
M6G3FLdAjEZboCS/seKH01QZRFTdPwCze7DZVyaD1VopiQeKs3kViLwzXrq3JbJI
hc90BJfo7LYgcdEc0KuvLYju/VhdXJ5TT7/bGdCidLNR3HCCaoVluppCAZedE5W8
nwTRIUO0/lh/4U2fbk4eNCW22Cpch7kbyfLaxIhOqVEzI7thndIFss/EV+i6kAh1
/IJRV1w4XuR5TrW8TDI4k8C5ESgQ6ZiAKdFYjbinSwRMElLNNYoZ4l4npuzhoCER
XQciqVUeLr3FL5aFKmCaWvW8kfn8KOoOX10skHkNVUf7PRJn7xvFF/uTOhLyX4Kj
TS3FjoMnY+gPujoXJ0IkSQdvt1Ith/KztNYprDaI4aM2PMMDyRLg3Jyb3N66fUPc
GcOnsfFXf6bhyiFnYNqDyqufyiUgY+kHb12wzc3yAvZezr8X3PHYbQMNhvz9C4l6
2sb8oqxohx0bxg2I4MztgKBGe5TVmCVsg7dINIfnjWbCtlSFw5C5WaM1aaoDnJiU
bEKBM/Po1kUggEb4Hs+MGlK7prOPkPlziEC48laYmptNR5DSIvfzcNnFPQYOiVBf
Rq5hS7DG1VoDFczq68pPfds7JXzIirQcj39gSCX/DmXVr+BP+O/0GKh/VUpYYq44
8r7zT/YWlH23FeVYyEjVAyeOlY2YdoIZYbGwXCpTXaTHxNq/d9AdjAgMVhXGJ7Et
NGzRvhPkHxhJEfCi8Fxi4s+//F+ci42GFY97gkQwvZm59GarzHNYgCDlVKuMGYMB
Q1CLj3eN8Zqe0HqKm8Gi8B/Kr/BSUMrL3VkLSTgy4l1joSYqyaCExdcCiYVG6zhG
L8UiKj3TXwlYtxr2A0D2rJMVeXA2hZ+eDwLle2U0AfHqIwta+PhB6s2FO+Ti04L4
khySeSj/RZ8BbfbRVRbZWFdRV09jHceNa65E3M1RjdKKVHWeiTFhkQ9PE0GbiY12
erM7h6P8nBGXnwP3dlOEDuXPJZtwkaktIgvNwy09o9sxMlQTOTuVSAF+U6Q0WS5p
v9wJ0lJHm/G63dUOq0tu345eSrV/5DLrxWEecfkJTUuN+H/Jl2vXB8Oc0X25gwaJ
P1JKDxnhaqWuIi0q9wwTixkq2UYuF73IbWDa8NMNxU2uByVSJFQ98iLmazehQmYK
YcnCviA648Csjk+5RvzSLgNYw1u8pgUnevqHv34iWWzniUpLxEjUpje2FomBkPJT
IzijZjR57c2JVSXQZm/8WTvXzvqAS0NTWrlQhGRtaO0ZrqWPTl+RCCJgv8bvs21D
6vqJSmhOBi0UpePthsfQQAsXY53mtJ9rXaa1lRa34RDvRR3ApWnlGr4p0SGegnNT
kA9z2jFseL7S+5O7WDP7wodKC7MWDHy3Zho/1kwxbx/TZ2+HJ6kaWyi8E8tFLxtG
M7mwNBH99YJxxf0LdU+2goX45DKM04Bg+Pbkc1HFiyPbMnzctAPw8uzeO1fmERuy
9WyhjdxeEvYrNh+TJIMxPyZA96mdPrCr8PlBL2r6ilSWLO+xXr9jQpsrYSvMUUeT
66YrFL389FnVM8/qPKFKlqszM1CfvRmG8H4ZEofiPGiZNst6R153jf22PTrs9tv3
+Tz6tYLvEki6SkclEZHVSxgIWld7ij2a9agilpxKKb79L5PGLA2PZm/mRtt0btK8
NDJMSWlOpW1SaqejREJmSyPsalIdQ4O29pG3JuPF2YqkTXEpyUuOmuwIk970E9hy
Bo8WQzOLsQ0+ZheqFqzjQQeWLpnHibEMFpJ35yuIN9p/L+a+Q6PTte1rreKgfKj5
qJV0icqfTAbA8UVh0m3rSFm9AM+wj5UyHOCGyKaFBL8S8vBIOniarruyGzTbwuyw
gOzfprt4lpLOEkTg/ElQu/sH0SUepp4VGACcNp78ReZ2pXbtYzQifVMJDBz5Qhde
xOOsXPtXnywRcWnRkJ24xHQMMP0pdTAz+SIrlZUNzSQFAsARWxR7YTtgEK35TSXy
T2DoD6hh0euioyE9P5KcO2yrK71FTNydJScSn+NfOPeM55Q4D9tt09Ba6SrsLuDR
L0VQCrYeuACQkxiWIlCdRoB+4F9OB7tDWeKkKvRYKnULhvHl2zuiVaf+OUL5Y3CH
po3nrS69x1ReQhWUSgrusj8vosQsMrTKn+VCfqcUInMIkl4HFJGaNH8i5sxfgJaz
l2bAPPNZM8rAcVov7kwHv2aWaeDnyYPzEEUoDHK8ocDyvpTeTYJ1An/8XfUINajt
VK4EnWqXQhQfTwCkjrikCxYGbIAIEmAPIN9OLci3SyvmI7hZUsBUlt/Swj+nzq+g
wG3pf8e71x/fd2Nuf8kEHYi+ytjMOGkLRKvA2zkR1MZJymqnBnV7ckfjOQJwXw/d
1/VQklud9pWpcR4MH/DS8Kb98wVPlQTT8IGbc/QLtoTQQvEd1ERHQeJ1srulZimX
yRoBIoQl12KfLVZ1o8abmuWcgK55rG/N/80rv343QtDHiRJik3dVAr9nePFTuTrg
ku+h3W6bKzx8jO9cFgGEr9MDTqmOnwiXbrU+hMNg+WRwCHdD6MVWUa1VFpnX9Kxy
imw+AsjW6BrRNsnxH6+JU+QmllQ6gmoPxf/wjr0aFVDP/BkhBFpdDKj+CG03gSn2
Q4+ZJ+pt7JJ9ZoR/JPtVeYyIRWrJ1CUAEscOrvFWL/RJMtw6iFKGHBWKmVoY4hbo
0P1F1Xco0UJ64Kmt+gQAAYAfM6jI7aP7QFybt44ooT10E1Y4SGchIwPFJtvAe7PN
hLyh7SSqzXR8++pxNZ9EGYx2ENNT2/886pAPQwUDG1jGmV/0t5CqUBAkT4Xi7tu2
lgQBbl+Vsk4/3gSBpKZ++o5MK40vOb0cgblPzepofv/7G2mtcYA+40lFi/6kFIfI
+2+nmPBhE0JFL4XKKYuMHezTzH7Z/ijkzH30dNSsaJ3vK+GEY0Z6d7NVdWp6kk4Q
vlW2qqxyoyKqMpbzp29H262PMNW5qZZaiRTTjOqTL3VcylvTHJVJt6lOYvtTlJ+Y
7HT063lSq4vwNqyxxqP1+KDUaj3AOHG8jbki2CvAh8OKBQy4PbtIwaI8xRFJBATe
N19ooWLQ2djvL7PkArHzNVFIGBkVCyCtuuJ8vZEz/PYBerRvGHIpdOT/SFzZNuUv
afTzJQ5k/anvgpb5/qV4OHALe61ALzSSPAJwGpfWqzA5B9BbieafgV6Eg/X8SYmA
PrB0WT4BdeTyoNhuuDvSKF/+LqrwWuQ04b8nUxttapB+YsnvHKpmqUvZZ+1CP0xg
iepdKvCGyc2nFMf6AtwgWA9f7G0Vut6OX1o3//+xIuL564wpypQGRZqcYwtq0cu7
I8jt5D2DVy37RU1AZJ5Lvf1hG7rHKEQzU0JqKl5h7eexh3te5iGY9pcNrJm9yl7m
g2wypGzqm5/YwWbZyfpJIzRQxxOn/Ep4J6aXBanGIZV1IINzjivIy5RrpZXUAPt3
USC+iO6/Sd1neCHk52MDeKSN+MO/r40FU7hvJ3Ms1gjecdRELMcRWyftediI5xy8
lUz3U6BuUBLVKG6m0jh6Jzz94q6RbFgFDoJL7w86E2CPdfSdKh0Ea6GsQPpudICo
gnJ0fUXkpxVEsxaixefMn7x1rNCYUQkihTlbIb5IQ+NQk4UPEJBfnEoG8hNnF6km
5Z9LAAVxoWTl50hIMF/O0lHqL4EEdPlvnyYlECLoJ+pchTazfe++ijEA9k3gqLEu
IAfqD7ZAHJAWbppAhLfpFmlbcJdqBvcdUZ5XadBEcHReFDRKjkC/kNqXJMCjqrxB
H3TwkACCUM/SNpeTPfwP8rY0Y+vv1PAfLOqRG4xsUaBCOa0RJtaM0kI/MpnI7YrJ
h9NiccEO0BgzwSOcKGcFpmcZT3XIejDgpiecXHT/VJwp3aIaFyBlBKw7ytt29fwQ
pPeJO9G0NIo4jFBNH2myb+Wn3SduAh6CEpOVQIJgBr9CNEhevodGNo33txE+R3/z
L7YxYHf2G9l0G6ngCgd66G31tCizDcBYIXXJ9Iif8Akss5yxt82/RUadgfwEehgv
rDBuGcVQGhgcAfks1eP9txnizB3vhNe7v85UE7IMGWsFXdD3xor4f0uUgKlEkU/5
mS/0ScZu/KJ0I52fmBuVvLzX5YVWo2ukhEK1bJjHKKkvj7QzlOH7s6FTN0tD7Umr
V2vH+nz2i8eVwiSBmQb6PpmWn7N9kCA4hIzvsaEk5Th6Us1Tmg4zMxV1Ky5/Y3nN
d+QNRCb1fVrFOSUHYCueSb+HxI1A0Ht3a7pVjv1LIv2XDSryoxAN960gbk0O2NJz
ZW/MsHUMrfT7R7glkNQ5tDTCoaYVD/AF4mPsPw87SWSd0KQk1mI5oqOmv/uGnwqc
HKhw4FUmsQISjRuStKzi9Jqfzk2gARe4NoHJBLYgTH3Cqu+0MbcYI4Mq9HRBW5sx
dm+nGpLztSSVbtjK/6EA/nn+b/bhEdW5bQOAJwY/1elPOS+QL4QVv06cjq0yO5Rf
Fl8PLg/y0ia7kX/pjBlWkf0cCZ22KXgi4T8WbiabDGTmxwqsB0M3tUbeYbIaMqbj
0cqb+70mk71DsbTtYs2bcRBLcWNScbI0TZkin+Isrl72dqZ5UH0/oe0EvUCqEWWK
K4lJ5V70z3ELDDXtmRWWX446IZoWupnuWo303RoPCiuoOgzwi4FvCzHZPTVrX09J
209zjsDmU52RMs++S/Uxpi+Q0D8qUtNU8p4AXkGE4p2OC/RskYw6QnWbRXgznoip
vPf+oaKP8J5nF+Zh6i2LgrPAmVGg7MZ+QdSSV7/kfEhfy+O3WTgBpkrowQcDoqzC
VJglJ+QeVKo5KbHaX89DFzS7RNjMcx8CeT/mizMqcwOOs2RBXsJcFGg4wDWVUkwn
VR9pJyWayP4mwmai9JEuX1v/gIZs7crCxtg8e59xVFdagFGUFKrCO65a6LhEdKLu
2ZPaBeliK5RxRSYQlLV5ZctObbXZ7TPDAgtRhGll8Raoa8nq2k/TlxUhYyJSZRpx
bjqJjBHCzK9M6mcSNbpF0GRLz6YrDrByQjo4jq8s1rXDpSpOztZ3/4++qvPsg942
FETgAWknSaH0khNZ0wDiVoCfBAgjO8vwSxDX5tCWK+CqoNmnmMUXUPEPkWUbW4rw
+xW/GXMARw4O+P9DtTGb5QNyPhk/WPqdrVAijUYK0vzGheoO6RZjpy7JiWfKqAZO
myil/X9y+QgdmGCug7P9N4+mBlZ47sIAhCBP1OQryLBB741EvpgoUtkU6im3d5Gy
1J8N9dl3sLdJn/VxcZc1vfnZ1eLIeUoRYKntulo8AykX9Redyk8rDLmg8Mq9Pq0Z
CP3SaxvCWzyzTLnHa0DVHge4htLTYN0TXrcS5bYfrLqTO5w/VCXOAqC6viJ2QtQm
WPvTH2FWUHtXQ6o2hyUz22IwnW5iArk/7aqJRune3tVY9QORXpngs3TebS+MCl0A
KXweFxY34XYb15r5HgNEuJwxnPO5WVWWbWdBax/uvpasA+9cNnfo76aE6mOdH+WO
wCFBEBSqS76gw71IPND3Zb2vusEC1o5kPAeJU8SDb2bVcITtyHPtu9BMUjQ8xMfR
TIUcgWpbX+P8/DvB+gYYWNCZV/t7IvjIp+iB5yEyayrjNgBea3Ak54it0OyUDIev
RCJ1gvrPoOE05xXn/zLa89JCDrxmxJiwoPwOLMQhJTgQR3ts30DFN43T2vmYQ1vs
UKGW+tSprxtVROVvsHORwcroPyVwclPWAmyuI/+Gv5vMBIJedO8VxU5z5h+Q2PQV
xh9yS6Z2eGh5vEIWl8afa7zOoMubOFGFvmWfRwwhUU0EQc9MeJVyLXQfZLAEpzvc
UP9ySkN0JnZJvsrH8agRhPvXxP/Y4H3tlagqNkVRx9DPQppINR2D1PA9fOzZAkpo
qVvAbz+rWpP9ZmEH6fCEqui8A2uisYkTMRIK5D0VdKZNLVKQjTJELsF7ClxU4WXL
DdrcD1xke5ogNK0hx7j0lHD89k0N2PxqJIbzIWgXoyk/Nv4BQgKUFUrE8kR0z+AK
LztIRwW4z/SVMKSVZKp31jFWZQmUHCxZ4VYHtls/z8QG1zWV4/XZCu7YZFQSPmV5
RhXwmUfUBtmnZb5FDmvpwN2mNBQzIaE2SwDu8d5954HIaHyrIB9gFBUSFA/P61dj
1kxJqvJ2pScUEXJVd2eQBhFGx/FL/MqwWnlY4KflnG+IrI4zjPunND8LBoJ8TBc/
nqxu8UBjahF3LZgAs8oEML3pCbsrLYCF+/bKevz464i7k6yrgQ0jq6eur1fEzjU8
l8lowySFABK2rYwBxByX+WcvuXb/ZQud9zdOajvcb7idc4eDR2GkSf8INU40Z8wb
ugm/GL2l2udBqUlaE66suHRmDnwY72d6ZNJEPcIfpgEze83IKyuoFhNXmcxymw0g
ONLAnIV/NH4ykyVVfOxnY0wWtPT/RlspBsTMX4C4fXIZ3i1qocdoPB26w4pSHmxj
MORPHfFxJ0uIiJr5LD9Vmp/sgH0MiiAS8GxxPPtgbrs0OaAEEqyRwtjm4Kqhjc4R
zliOHoZB1/4qXIwkAJqUnT09v+yvfUNXEV0CK/7c3+92sWn8+2DEP4mQIP7goMMt
59D0SnSRoyadA/yKOmvVsiaXMxgbh2OQO/bNGnwEzZQSB9fuFtDJdr1gbYcecUjG
oZzGOQeMzTT39RL9Hjd5bCiNBXNficxONDhJ+SQcYl1PGrVH8OGcrQE1zeAhyJtk
pm1WqVvNai46kcqaIk7DNXuswn6r+ODNMLgZP3AyPYMwjgPCeN8cVHFdfr49jtAr
SRc++pbdZO6rYIiaB4rPRpg/At5KSNCSC8vWJAIXErkGgu9iBQQHX17xEbsssinH
H25hvV9S+mRA2kMW2nrqX7ZRR7O/re/ZTHaT4Pq4y6zp0HLvuRujGi6/roKoeaWc
m87UhbUvA7RCWNpVrg0kh93ADnzgZbkX+meEEfAGGI6Qwv7VE2DQRIeYeOQ3SAPS
F1qVzoH/84fPYMNyZAlrFNZXr6WjQT+4unODq0Wol68/ldutSPEKwIdkN/rjD3tP
5I65eD7on2e2HdFl4DcDoLAV9BdkyRpn2NYr7RwcKcmZZPoSGUNYbp5bu9f5BrcM
KrIen8uNWMETvpp21mBig+LgbtR5eUrt1R+TWokSPmrhxyNf3Uiqlvli2spZSpOs
FnY05hpnYlJL3pwdj5wdatXpbadM1NnNhMZa5zWO7dcbujsyyHsoC9wdWT+vt+Db
/w6pSfFUqz13ViQ+onadq66p9OlzffyTkbp3iDWVAd5KoVHE07eS64ze/co6g+yD
yFMsHYjO480AA0iFXVpqpvoBvUCfGhRew8qzml5XpVhBLAf5CE5Bca9zG20ru9YI
HTfmgdN1zR49SLtgJLzUmamDvoT5pxmKI+P68Vhb0FhW5mPE2N8ZftAc5tzfId+e
R9tTYQrb5B6BLRlEEx6nWytpFLPat16P4y+0ofWTumtC4y4eeddDFs552+q1Ia4b
ZYCTgzQjMS6j1DM6THX7G7ukEdKYTlrNn8M7EnORzFFrrprxb8KWVZTe9OI39cDX
XzWbpBfKmsoNu5RaCICgqxQqFT/v9zj0QNotgCWshownanXQ6/5rVGxvFUCTTvw/
FVK9h55zp9BUPf21awPTTCAcL1Ex4oRu74PwRL+vAo8oRxluEH3gHXiA/sqGFtVQ
5/SulzumBPkZWOBnnxSKE6VfnvuF0QrM9S8RXGHGrFJi9rDA0mdLY7CYf/d6c3AC
zMbRJVHCOXVdq5Gpm6wPm7B4k66Uy5tCWdARfLyG3zG3Lul307bzvuPOkS3tX/2L
tJSvlig+Nf9Xu2fcqlrN9VxlmBRFdTkIWIk4FlZc1MGeBO599YvZfNsBfubuXsZP
CDtXeQzkdnMAkxmi0X2XWs5L7+nEnQRj0/lrhpqOIHhNDzr4ru9RUFr4aZQDM3lW
OTJ3Hz9YtY73/CBLg6ot4hWflMiS0PrJmR0Va9BTEnRNXLeKAgfYGzeUi7+kCikn
xEOMQVga9GWiHNAcDf1lkBEJ/YKdyHM1qsWIK3wVnP+ds0cTYqHIPv+8kEYAoBSL
TYiEYlSAzV89iJv19Aan6YGP+oeFZGjhtSIEoxOXnw2ZfQjSV018YgzqHk4Nto2P
QqWVsO0AqTifiCeoFBoAtu3bjwi0QeDj09ruZeC70uR7guNwqOk/8IXtu9MZCvmg
QhG8l8u+mWAayPy0K3FUrwmx5+bu0jQS9SpmbBJBJIRNM9tXEA2yKEvrQ5bi0GpZ
X3Fh+kRJnrOL3FrLC85RNTzCY4B0u+qdQmprN250TgX5wmgHLtXtPxJZyEii8hvM
bdEQbm70iwsjyjlRVtmZy+WSBx5Unom2bLV1cbMPvBONk0u4mLasPgWCNfd8S2LT
J6m1sh/bBY1SFf+oX6L61AzfK62hSpKct15V5Oyat2yvJP+1ovObjo15zZ/lNqfN
o3sKVW/kwlcYeZUbhj4ND0prHG2piEJ3x/suD/qVa4kfzxqlozm1lCEzxMMJ7LVF
5ValcQ765ZqYYLVWKGEmp+NKj28xPMNg64w1PmTSrCkpBHQpojCp2VN1O55MANT6
XqpLsCOfMM79KBC8jB3BUwK14btRFFktBPH7CsA9DRAonJnU4CDiPvpjGYzsmHpu
JqNX4xULx3A05e/Mvx12MdTGKPD5rudPp+GoCuPcb8U31rGCfE04EDMXtBYgHLow
hVvVxunGaurhi1HxS6T5iqzcsSpulaBLqbLSUCsmXPbLPbYeMPTsEa069XiSaDmU
cn0ovB1DjD0Ab/HHMbKKfifohG0OEjx1iNOef3gGirKWnR3pRHgDUfYd68NW+yy6
PycdPRJc/UoP0JmexQMmwCF8O1+2SjtAEeX39AvQMAFE1zYHtR0McHGEx1AzcdIy
Uf2Bqo51MQDGVYSyvjtpad2WhJAOVcOAHJQ0eHC/I6lOC6kPGoq8nYQQnGih23h0
4wwzcsgFhuDQrrN2byjkTYm3r7JH0xhmRM951aXWl8sn5VAL0kwgjDBOuDRGaGCX
LkLbLrsGtyUtIuh6DIzHfPAkfCGgkwFVK3ADM3aukt8S3mShuMijEHnfLCTzTdLZ
TcT0YcIbppVFkL3kndogcemyhRHDFKpkN0+4jTZw0sN+rwtwi4nII1iOyfAc0Pgc
ItBf1K/dEgnFZFC24QbDUGWwCDRP9ojVuD0kr0MwYaVvRnnEMLiWL+52Q0QElM1G
IZLegPNYnWArQlJkyn+NTI1GHoBbupSwM94v5GDX7W93qEfsubMUw+LRIEle21Cd
aiwglrwYUCHkIVqurhx0J6uO85LX76XPclwvuMbRXq4sXkdnRFUA8JBqOwlklOeJ
iUpB7zIw2dbV/vccN7M5a1VFcUrAt6g7TANcXxfFzi3PhnrWTAINfCVNrfTvyrjv
KJ8vVBe1ijEYf2Sk/JxkXzMb97tFeCgvhTvkN702QDPo0cLG4H/h3NqfiMaY8xNu
LO/pdQR6J9XVzaTocST0iX1wMPdU0opaHzN7n5u6cq+H7llHX0aPVu2DyhP7ejbM
YzIrcjb5HPtDNbdgyShWpj0b8D2ZBNoCgGvdv/n/7NY/FR4dWSTaXJF6zuqEpLlm
fKnT+hNtBs1lQyw07NSpuLFu99rpwPQheXA/0fnVVz6bPFxVjZRchTFRNv0WwYho
gLYyOTronDY8IKf5bDFFKvSMQxjr1ZuOIhx+7UBdUrhoo4ZPA1BPgPDscu0KbZjH
EJ3sh4Cyh/q679ME5gcS/Bbtcd4wImILw7VY5cPFeu5QhDr8lCyFjKx3qzL/CNJn
lJyy/86YUXiFemTuWIQEp6K59aj9Cccn/+/J1qwI4txEEo0ZqGsdLvSlTq72Aiz1
gW6R+pHLinv6vYOGOX0T7GdGqqO75g7DmsR4kokPQLeHmah+KiPSFb8wX7sUE0H9
QePrF/qSu1NqqvJmEnIum6nL5DaQB+lWPmMqNqtlxgmA/YeWUgT3XUNRr4Xffqe1
7hqtrTdzkU8R+nmKkRGClKbv40wSKbnp2ZWBcgJsREwzmMnhS355fozBaODCowRQ
1GeC3GGIRHEJXfuexvgBuXkt8sjB+BqTUgkLnXywA8e+7lhfygQtM9yE1+XZqFLW
VlA4PXXohFII70Gl20H7GCoVzwGoo0rb3TaNASwNq43H3wfl1e/PZKNB8aDCMpUN
yaqA+bwUdskRBtGodj8hT9ASM3M/Yh+ps+XDpIgPuFJ2jnWLgyn+9thQcHrtIQoY
aV4zCsfvFRj9VO1FvAdarNPC5Ay2RARrjSFTKimPX8TIuQckK1lIXpXf9oCPKzyF
RtVcZS9QXgCvuxjUuPKUj3BsXjTRiVVZhsu2y4HBKR7KVYYCBbGn8COqQhuEDrkx
87BFBORmJ+sdTAoqyf7FaE7L5GSQFPh4/ni1cXBrxayT4Hau9Rn2r1+sR4K2HuMv
QJCMBMJKu/Adra6y8cU4KKWCAsFQip63/8cHLXZ2UEQr99UZCatcce8OeOZr2i7Y
0FnZIMeWctFmVM5MXq+hW0MV8sT8rjfZWSd5v3Y/WR8XOkz7rwfjwgQKump4yjme
LSbNXaYjcVdrnny6aurFOqfKzVz1XGw+TowYmJBVLRryFKN0oYQtBIOV9lgVFY/X
Q1yfZjinOM8kq0c0yFFSBnGkamFswK+Hf7JXMzU+P9zuLi3/xLLlxnMPm90vTwuz
cBqhtTiOnqGrCBUBAAlU/N1BTE7asjLBRI4wgDQkPlMLacERHRQN9bwYBTlhEuDi
HNoPgjTbGcU/aDJu0bqi4U2fIebL1Rj0RbtjuEEPWbt30eCtWYaceZfjR+LS+k0E
lU9SdcJvuv+4j+evgSn/ZkRCnxolCJd5UEONx9DKGR0IaWporYX6zr47XHqwrJda
Qm0dm6NoXHntgodnseY3vwU1Y90cydfMP+1T8dsqWDHMeUjfegRN/g4LNw1B+Cs1
qR9bDGFEZVYN8Ftb6TodtoZiUxOrGA/+srXIhlFQTQasjP8/qkEuA8Qj0X1f8Fjc
PbNzL2cEtALDiq9UB4ayLXjY2LFfu6W28ZpMMwlE9LUfa9GxRSxiN3WRaOQN4wMW
mb6Dh5HDBN4NKRFcxdetXho2lUflIJHzX3c8mxCNjnbbTaHaOf4Z93Iiy6qv6+Xl
av7nXhg7sZU4nQwCiG0lHgmsApcrL9h+/y1Cc6DU3DLWDgD1OjgSvPWxX5tE/mvC
IyhUmST3xV8/QaEBHJVvHS5gZt//zyP0AjuGueqjKhAXtClHMqpitONjR0VS7ChF
ubYC06MbyyI74v7Dq/zKfcfSy8WfKgU/nr8QbH15pP7Ky5y0Ud59frEdvN2ZPjtp
aNfzTAfQJpT4AwDsth7UBP7xggOjQiAUaGnovZtykCi2CQP/duG99oF3tXccznrt
Z6XzKdes2v6tLPPzaZDfF/rN5gebw0Aik0mor/zI5xZcJ4WW/IR3wP4msUrr7+K5
ODZMS+I/GsLac38SVhu2V7YhXx78IsM2mORYzEo3oVwyFxLnjln+L79Ac6lRjAuC
ej/ag1GZmU/249YbPKst0Tt6Q9Rb6yoluSss9P8QlFBjf7sfSAC4OWrCPwMMZe3z
CBOdDoepB+YLzn8Vh5rKduL+d0/VFYX2yiWF59Nt6y4nn2pk4s5PIL+EtsWZqVs4
SZlGbQLfOWeRbyq9O8egHKOoGZX5UIgk+6wA/dWq0vV23GUPg5ytiGUW+7Dy+WaJ
WYF40uUHOINmgAVdDSs9V3bXBqWUwPbs+Uj+ep7X/AK1E0/rjdUbm21P46aCZFy9
g7vMSepGSDibbNxyWSA5w1mb6mMvxiKg7BsyfBMeyIof7QWbKRBa81n1lD/IQXBW
2QEpfgy8jYrWE8jMUAsfr6sZDMhXBJIV6yvW8cKqdH+45QcJ8nct0l/X6P1xp+C9
Nkga/uRV7ZZh6i9g7WVr41LgwPSHAjCYKON/ABgVISlnnU7pcy4zbZcsXHWPuBkP
s22GLR0J5oyzt6yuPK+K19bwh/WUP2cokMeA/tuJDHMKlXrE3W0pnBctjb/VTWFO
v9ScambkoUf4CFsWj2bWjRUuY5dRc/4QZaZmqUjoLA1tlse/OXpDJKobSeWq1fZP
hjRkCqESYniyy6OgnhyWVyulo9ValbV+the25NsJlxcKk84M/WKk3vb9dR5PohhH
8gJYLViod2VbEHuOya8E08gAPZ5PlYzI/SKjFyb83Otp8+TE5MO9FUxCMjHhL1T2
lfCjuROQKoIg+zQaVyoWnKtOGGC0R1nWywrQ4vvhwamcCFQTKOxgx6hXMvkUEDwD
u+pHsiZdpPIzjEeOAim0L6NpkvDh9lJdT2ilYNPD40KpNcsh9N/smdbjsl9JXIto
W9CemMN3nhKQSmZPruP4WAIIFTGaAC6IvZgNt/NDPRnz6eS/vEd4AGydOruKwS6y
HDFlxjpN4fcmPRprsm+QvjescvWAld7RxIM2uzbmkAYr2bt6XKlQWMdHkdufW5oh
l9vun5d5ob6O2A3nIg5hn4ORJHbHLjGxdt+WndHE1czIOsnAm1CDEXwHr9jaG7ud
PmoqEOMncvxERxsyCAc6ZEDOhWbQPDMS1ezX0UoLY/dPhdPhG/xnEdGEcZeHTlIR
wLt4UmzK6H9jRpkwa/Ow8LhK+9Pa6WVXaM/5oSPOv94pzg6ydopZayvxnumnuEdB
vXav2ZQ4jn9+byEaGa7h/+wifpwvgNBMMHXO88koWIXRVYA8CO/hgG/sOnLVNuiW
uS9xT10fl5WJzhIzxYoXgXP5yhrfX+xFsAbeXOYLkbB0wZdTNq1qhNkmKWXVnYcP
h/o7JKvEJAoCm0SavhcN3ynF7OnF3il+YkYgwBLmQqvj7QAJ6MCg/8jGnydiZyp9
gu5efRfAwEDdDB1dLia/Gb4i8Nboft6J5IyJoymdm/LKVDALEQLV5U+eyUAu6d1i
WMjlH3NLrXJ5uzPBNV6zWpIrzwCoN5+5xsSNQ8hDMHuFwE/7FGXANJImB9OytMu7
wCZExNnLhdkG9g9sWikOr7PxXCTWCDwEThHFz/cj/nMc1TOtSrBgFPXYMfV8UU+u
J8dyzDb0cRL5Zeh28wwSh/jWVgmTix2ed4YzApO+7bcFIR/Oo0KXtc6XWgIMHewH
sM2uRiulpUHG69kka055iQ2aJ8eo9l+opwJob1QptMUkj7cq68CPCLDPznEctuPa
VltW6ahIUBqkE/4kkywOWNk78ALasM31kgr+KWj7S1CTowsk73SICa6gFa7PUZmd
yGox98j9ElDK7Fm9+2bsumt7OthuoJJJ4L8VCjdNTh+ne3H+X4KQYLjsmJ/aq4Mk
3wPjTpJxyv/8UrdrGMMG0EcMO+HyhTsfzU2w1vI605KHSAF9q1Lf7XMG3lqtChRR
07FNo0BMznS8vCxisEM/Ne5ZrgDSaV4INYJUlcZyKna66lS+AFUju5vlWZgGE3d1
030ywmqeNykFe370/AclxUpQ+tEUVa0y5zxJUH9kaLwICaczXymWYiMxk5Kv00Vn
Vecy58Oxm2M18XHowDruuxRBIvPickEjzBU5ADIavOWRWT2ftBwaFftXVRXJdAue
kpfxtNqrkFcIc3n5XA/HfylAPmLfMglFm9xNX4FV7ymylC+vyFaYUqwOcjyaB4hd
OEE1hGFuel2tZE88HmFEeFb0Sj4imxJSyG1pmppNxzS/Hh+M3zRyMqnu1s2yx8wd
4gbxt9cTf2f1kJIz7rcxE4zRd1nPP7mAV1UgKOH1dAPVeWRlNxIQV9Wid95MmB/N
V63x6SPQTuP8NNiVRW+bKSnrTKgUZTgrHF15XXLnBZb30aGK5cleCe6lGfWZ95Zy
1TpR+QYE34t38IJtf78mlcDY/zn2caaRvLD2rsEvtMVpieGRFKNr4vSvAjznQRVt
Wi7jpxQ3+sOE/3LAeLeXwefO/myczci2NpoPGqGwQz1ecEGItQzAfglhzjGCYUnV
YLYUHZnTlT4BgOToITKusrTZApmzJSBWQ+mB/qJd0TWzxCQwSDwdL0IFij/RgnrG
xe8JtguqgriJ9LuxKrCPHcOeYw2/48jQs2ZyIbhQ/DXjEnFHzCPPDMwPwOADPyT5
W5OQ96rn/aGpXPv5OiokB5OrAYkYQvapF+awp6ScZiYxYfsC3THtuIdQRL1AVHWQ
IUFCzMzURBqb27BYqTc/80CqvssRfN+AT4kKuV+Y2Shmd6wyS4cV8+1tltNH3+Al
z9Br/aWxP1xnyZ39zhOJ7o1Gq45hDYVA/ORmDtv7p+72+DufSCnykvZkN3QlEpkJ
XsZOcgBMYbazQ+Gdg7Zny6NbfUXU3oG9qae7sp4u6A4+WTPuPlnxi6aG1ULC3Jv5
TB+sKIuBQsf+EtdMNFlAV9L10QDBsMGDM1TYmCjG6/s4vi5HhcWVob1bzsAjE8bC
MhmV5mmyK3VtMBNIEtcIdxMKpfYDNp4Kwq15ecSuHLY6o7svUwASGxGa9o6Qmibq
sFc+0HME7gbfOEleAEzsyuFoEw3EVydwCRx0QX632y9l0KKQA4oBo8f0Pcei28mK
IEoOtmeQxqLPFLpqHOMIjauWYG+GZOiwD2sALC7Z5E/+xZUJVUeH9X+pZErRo4i9
9JYOBrX1EYXq7wDhQeHK5QT9Cgi+055M9cZ6uQfy0Rnz0LgLQbA1Ljk8ztSq5oqH
2dxidEEOaIW+HEPiRvIK4sTHaz3yyf/1ss5vItINIBX+6+quiQ/iBDXI2iU3ws0J
8vqeBxDwwqf3tgUZEMzwUko928zjXyquwwFYLeoxud+2hB5/4WyMXzKaKmze9JLa
21CHExsgv5icIJRz3N/4Y21UlGBRg3DubzvRVzAd+/hCSGmoKgrn3op68rAMqZcq
4YXW4jJ0Aij4kGfEPcXazBpqqfjfZpZuNeJ3/ilL9D19JyDG8OAXhp1ncACmgKge
m+/G+KzIjXWEj7ppHfOzW02e86747kxBAxE/aLqTV/lk8hUTwUTGTzhdeQXTfNbE
HbN8BFz+O9sKiVs9DVqEBmeWKanmfEpXTosEmG15K2G++aQx1pH21KogW+bbi4LM
4wWrJ087aWrRWPvbbDyHsNk+9YbagPXVsbo1FwyO+n+A5By46zJEEy3JXKNcC2sw
U0IN0VaE5PZ2xswgJZl07BtgYxwvMg/6W5IeyP+KzSZkLeOOUXEyZ9IOW5cOazKd
kIZwX8YE3yhR83d9lfvS46hodL+ndFJ2rDa/4k5u8G0aATmOl4IRAUn2nxzBxYm9
OG9WPV9zQHMljg5lteVn/jUE8FDzsbq1ZatkDxvx2HnWfW4FYgEwS2PYQhoGeN9R
ipb/FAdAIpvezluGE4/9DaiNCjJsNuIklVC6vYAH9DIBmxWRxTQcYDAOSpYeYvc7
eO6TUp/A7hfXWpzNohL/ADAcfioiJ0j7QFFG5vHb3N2hf4Sg30sH01UnCReDeTkt
3I4eVSkDjkkG7rAWhozbxS796h4HAB5Y8TxgjVYpGTd7VwNX+2+i3EoBLzU7vsOO
9zCu0DPVv/i//GmYvHMQk4HuKxq/MXXcc50DR+atFTiOcq/QjzpwbJMn6+4eazBF
tnskWQQiLKR//UgjnA7x1o2DUfijwxgLtEELW43MlGMXhyfVZ6X3SxV6toBOkyU1
dxiW3xyeZtcwRmQH8KoD3+eDge4jpvRmW/xPAGAYhhs2SseQ05T0LlUUVmxTX9/U
U5zKpq7edQZOUDUXCi14hmHvUMKj0gK1SqOIrWiHcpe2J7rFVGaH2E8nYmHM4UxO
rflFrUC9KBorcfuFkAchut9GXV8oTntjXfmaZlmSrFQ3FdrkDrS+205v4jJ2MVBn
b6ef/TEbZcdGg+Jmg9b8M8Ou+RuDQjjqNWEmqN+6MIG2UCGfGqBzld+d4JHwDuu3
i+Ebpl9Axeww86UgQ4o5/gjXuDb9ywRgOYdV4IPFv7E/3+BpzXMYlQN0PfXjqYU+
2VNZ2eMUANu7gwwPm5VIuWm8ux/JduoaGlMarcnp4594lytV9x3bdHYY5BNv+ZMB
DEtF6zwanltATLBOi7RPnf7yE09LXoc7e+Bcxatj7CWTCJhPCRhXBi4B/eQcg/v8
n1MJ0dYinxZhZ7HGvT86BaRP/oOmnQHC54kK8Yuxs/N5HqjpfxIZVi6fKIIBiu9A
rrxt34RDhw4nVYBASkgJc6eIJ5qI48zMJ6GJLL1d684ESJzx/nT7p8zTNlZ9AQYp
DeU3jjACWgriY3zFfk7ag0HE9A/3Q54t7IVhdIWIonu8bMJPfiL9wPZZ4QFNFr80
NmmnZXEJqFn53kAgmP1l2rxeiU4U5SeJvQbE344D1gXM1MSS3+tXlxCiyo+c0yMC
LriELHPi0bWIgTCO3IZVvDPbnsfdNqHpjLwnYzkMPuWRcE5Z2Apf2nvpsGDIttu7
Ui8UbrAf1qbAiZlfHEo70j0bdwlnq+DUFIiuzY4UQrdcFL6X4vXwoUQm8Zc4CVwa
eX0juZttLnksV02vM7UAhfBtzn/NQGXS+V9KLT5JA1wrAVERFbBTeWDCQD+Lodii
fRVrG0/u2q7UDzicMGqvSPhXeNB4MHGedPn1L2P32BvQKoxQ+PnCdcZQqqp3Yqxm
1cuLc3MQnIEnytSilwo2CRtIv1SEWhy1pk9k8d81+YaGy1yOxhNK3WFe9Lex4B8p
C/S1D3OdPEFxsyA9cOfTLF/e4AFXCgJNF91sZ7/EDMYWyFNWg69MRRshwDN77W/Z
Fhb7XIsLCQg1q6lR8E4Z8xi1RKL8ITkMiTvUzjVf2/hF5bqk/sr/3EktFVwmyFF1
nrIkbD8zXMKJT/b2UxENB11zM2ej5xkrLf5/+UMCFLbjZGHEfW2onN+ZeacRDE/E
ga6Aqy4gI7ZHFmVbFE9eDLraax9ehUP5mCNLWug5qAmwLjBnf78+1qsuCzXf44aL
lkqrG7J8n0K5sHfL8PMBt4yAPDSjVzaczMUduQAtFQ01I/Go2AiESRu/SSMB+5KV
wW0TJIc4jgeURUB+oa1DeSuF3+M/A3ItMOOIYa+1zASUGyJd3/XPjR2obFQ/gkIY
yF/V+vJe2V4cY5wwwUu0wCK1UB/R8n6cxx0mKk5DSsUcz3qPWxyEZDwofqKxcEWs
jigevg4HPMcGFQdSN9MiS4IJgvjClFgefSyxRieVFLimqn37rBpijBEoRkM+KtGQ
fZsYwjdVKqDVJQORslKr1QFt1MISxPZo8PjY7KICIx2HFIbVlzZVTJXiNn5j7yML
kcEsAe+qXwswMN5JnPR5Nmn2Vta+VT+I8HIxIFPwUGMr+lIafVqneesS3KDoQXpR
71vuX4jdjlmJU6RF2InafWWyIHUwBqJ6m5Q3cN+i6PKH5fQ74WnCUGSLkdzGqNmP
hwYHhoq2dxCYws670FaGas7q1bR9agNbJd7ngVusbDcnO9RumrdhKJUkZI4D/M7A
Wb7iFDTnBVW8Y7SbM4IYAZJ0BJ5gJ2WCgJCVlq7UzZQjoJsfXXM5bT0/hpQ+OfT6
O1xwSPUtCfDdr1ncBj0oN7rlK8Ebq6G7Td8Qt9jIE7zDSd/uAWEWf3wcsHwW+C49
bFulpBCOBnXPrxcHgeHZPYEy9nu94dI6tAYkNcpVmUUqbFspxCn3VXmGZ2lZ2VBE
/tB7d+qA55zw7F5asqFqkrVUDa8J5Vl52NR0ytRtVq+IwigeA2XFIwTSf/q9LhNe
vLjGJzgd/ixP7A3FYSwXUBB7NH8X2CkTxcn2GMw3bu79m1By2yooqkm3pNHz90Fa
Qes8X9RJKdjakvlAzF1DGnvkgbIXDDNXCRCly8up2fzaUeAwRRdg1WxNV2EUTBZI
/uYoWzif5WywZ1G25sT8lLDcskhJmOrGN/wY+ES8XN2LCpjo33rllCZppFvfgeW1
b9TfkmHaugcr0bODSqi2hpPXRsgfA+omQVIiNZIlg1qeMMFgUg5l3ex4CqS2dloA
pXOUKJ4XHIsT73y6Hfnb0HSxQyQf/yc6nsJUzLyxUYvW419A0FxtIQHoc3mPxWJj
MI2VhEuMe9hCLEwJSLDVKpyy8CLGoETe3trlw2UVVeH9YJTk4CKWYluZJILesH0V
0YDjxgs8PcHcUYyNEmxLux1S6trdH54nAX2CukBZ8LODfEIvmXpqBKI7MJ/csKoj
MMka0D89CUZnCyoNz9LrO0QsPoYI+66MIzuLt6heyyuQ0TPTpTAswCmRjfHZw4CM
+LpZc5OSReaqTT5NR2zJ/F9zbGPIfe0ra2k9qXK8oAom2XYcnY+NoaZ1l4FkSVU9
Eo3t4n/a6BByfKQjPWX2nNeN1o/Hri0XvdfltSyYSMR2Uo/uW8qFzlyfwlhevcMY
2iIUb0nhTaaZFRk3jNCbygGRylh/db+298eeAumbDKhAie7BVd3h1LOYBDwrfQ7o
Vh9Yg+Nwtb+OSy8J+50BDPaYKW1/R0P2TsefLv980tHD+xom+bWOMSApuPpkUlsc
Ho5x4uOLNUkXblE/y+ZaVHcxzHkjXcf7eRU1Jypz5oCKRsAqOKfT8ojWiWKNiyKj
VQ7dCXgZkjV7bQBo8HqUOvhIhuf9Lh9WwhPVYGoGnxkicbbY8my315sG1UMMPspf
QumslYKQk0GHQN3FjolyOjtLEzGl9Ivs5IUB0gRGQ5bISn52lPBHKsBU+9QgOCPV
buplnpl6gNoKRgFuTsl7Lh2mkXN4wxrfV2xbjabGb7Vnh19a9LuAUZyjwLDshtDg
d8GJXpDI0rxzhnTZcoVmvZiTX35DtvOaDfcq35MaL81IOhK/j9UHAkFwB0WT88zj
EOS0ASSvKYYaVUILPVfBgEQ08+dzhIX1S3gZDgK85EvwiLcZoPVNnOpvLhD2o9/7
E+K6HRZIF1czrZcjHCJ00ZpJT2Ury6UdJCQVa/BgCNqPrTtdrS2FJxhyixB+aeAA
TqvP0UM0QlNzL0bOp0hioAthNT9H+gNgm1Xr3l2nSfF4Jp1yZrr1UtOUmiVRK0Ak
1AXEAw2BxrZiE47b/5PK1BApzyknDqMBhg7ewNzprAsDIs6B/oxBlM9rr+A1L6Gu
dq0D7ihtErePTTRIhHVnhxxXIzgrGdVP9s0ODqrhDQyDGknsj3gM/eyx1TRcv0p/
BS0Bzd2qe/RuBhaclHYX73ToRawsfdZ10wk+KzDvd76qW2K2y5yPj4zFvMaTaVhC
+obgBEaDpCxoSXIJ0jngkUZbB/XkqmP7k7xmMJrOz58cj9R00n84ocQgP+wxIwE/
8TVAXPQ4ncgRmY7nNbgZULj0ugRbJ/FDYzMTN0N3WVHjNN8CfJLEBuxYG0W1xKnp
ZMRDzmNuoxzuHnPPtNuNgFuoyn6/vNXQp3qygOfEqXTscryO2Zlv63PjZwoB8nsP
wOcarqAwBkvYZUWlbh+EWC2XJQAb7BLcqWWtb3jziDSo3XQmzZ84IGwk7Acxji9o
50UI0FNrV3Z2WaJNgfmkvb8APFAsKsQ8jclLFAn+pID+lK45jtoPyhKKvtFLdDo7
6rmp7OAz8ze+6tnaqGOr4OTH3wp0+e9SE40X2LFC3kEzOtk95+pZXZlnDnrTp9Cu
vrUQGsgn4SS1HyCnrEqWltGSSqYNfIMq7rSMwT4t7vNWYdHtxU9su2eTAH1mPQdk
H3Lj29S8VYHICttAg1Ubmn5vVwixsEXA5igx/PVJsG+pfDZdsKPNqy4Mi5TQ01YW
cwHRHtFsh7NV40zARw8gvJG8KBLrPVR6EYq8oL3/HcuS1GOHUOyXHVjY1lK/TgTy
mTB3FZMEknnATyCONseJ0Idm+jAnXljHANXCedBNw502jZhrVMTIKlkoFjCUXa2n
348GNhkDVEIDvRqHNinaOBwwC0gQrBvzOw81xvloPv1yjEsbBOt9+bjW02w9WgpP
63RV0Kxv/6qBup15xEcCc9e5tTfTAA5XTxP2DYqr6vvHzKa/yUj0cWf0+V1G+nRu
l1QjlxVCFxzvfJldXgWfpDzzgbiXyqV8HdBxCH+dwtgN4+/e95ZktfEG/CJ9NNCq
gJVi3gx5QXB6IsPOk2JRfRGvIi6cEaY61Y4qIxoE/mhqjOdg6Knu3+81rMs5CIIN
6JBxXgPOg9gnjZpPMjx16vrlr+2Rv+Ft3cgeoBPl4u8hFf8cn0fUebZNQm+flK5z
Y890divUuUFFROHe0ifQ7HPr05Cf5LJrQoMmlK+oG+jV+Ofzu1syGkGTt7KucZKz
X5DdbYrNT44T4PEugMW/ZgWA0cPF6+s36AFqRlQgchxrVAYKmheLkdfG0y/axDWE
uO0ozASvhnTvPS9fjUHAeIayOKrQFsKmbxXJ14Td5dKheBeAraV7/T2bxpNmt2DJ
hxzdJAtv304jVAeZAoAtp/Mfc3Zm6Hk6zYPH7A8Gg9qqCO0SAxGNvn38CMEBOXjU
wujCIdSw+9qMb8Xp4K8Q0WKSMvrOLj3oxYLAj4TJQm0X7SJR0hJn9EL7sR+TZLLL
QnxJoUa/g6t9Zk7NCy4s9jM1Lrd1gG+CqAn/KjkEF5aXkJ05F+jMd+PtWNJRATvw
Khlxtx0ecTUVz2PE3xyzXl2xlG1XIxarna5OyZw9x8r6oqwU94WebigaPbUOYmda
pDNk3bwAZs0d5mmSITlnQOQ8E0LKwMCttwZzQuVUDd6kv5MThuuaFBEBJTZOtWtL
3fUw2C/7GQdV+StHyeylwFOffM2bHrQC/JptO8l9eSke8NL9GvaXOUMTj2nryBXg
TeZ0woHMidVjgnX5Jtdr6VckKd+fBmIJbik6mwu5G0iLnyX6mD3NY4pkbbxMl+e8
jBo6PZMzzhmYBP9YR8aLdxBw8QuGb5eZN7zkGlDOMR1GAKAYQFASbYaP806VBnLE
blVAcFEhSSH2EK1+OWscsr2Rc7QtOjq2UfFW0HHwfySZRQnhzTsxMqWcZPc3b4UT
5/cQlQ1uW/tA9J75eJDLx7jkklfnwHHcxUeojIG9QOiyh2t0zZCsErOUo2SUYYQB
wxl/cMmvfvt8RQZMAqi/Niw8rh8HxX5iT5J2y/+K76vizcj8UNEns7g2YzdHBMTj
UeYjUQW+fde2//cwMBk9YNq1NKarqhQgdvp6gkOASaDw1pCGh6Ac29i/tfe58WrJ
5Os6fZwGgOkUXoRBGjQxDYaQxfVg8Mk/+IIoubMtiL5nVTBBkAKH0drvzZ+ZuHW4
LbxvsLtsGFy2JRavMTZkOzFa4JFxRdT105R63nMv4ZlVGfDHhxPmClCj1s/NmzDs
7NIrx7B2JKuzI+DBqNQDvO1qdjOJw8L1RUmgz8R8/qJkOF4FdSodKyD0dqAxsEvT
A0Jotmodo+irZbk6b81UKuvTZtiRMsUBTazrQa4YQG/lBW2U6xebC7A5xfSCuzT1
8c+E/U3/1alC+uToGApqEoOmFHV8FRihAMjw+W4Q+GaYbR8PmMWpuy9ImNKiQ7ow
Xmx/f8qzYA7V7wr4DtvjzYJNlcORK3c67tQfW2U8oi9cogPRYrO28pCvubwQeiTO
jnbezzijTHkeMDi057BYKZBDSIrlWaLC9f4O+Ni+GJzD6bhTfftf/7tNaL+SOu91
zYgixwWv9oKQogLT3XJNwigevRhdrlwynwr4T2MTYIs4Vz85iQm0arMmqpOd4naL
30v7afP2nSK8l9O7gJ/LGjFBuR92Q4c7BhhxeTtRIbaBStQDerooQh9dV5TUi+/3
/UcksyBjFKz5vqDHu5qiu7s0eDd+lLWVWQuqFxZxC8LWuonZHGexlD0a7dATKBML
EYQbJC8Dd95rtOYybkKsQ803j9pjT0f5jEpQFHRL1raq4K2GrDCt+a7DQKb5sf+v
Db0l9MzapWnTZ7TG8X6y9eYZdzXAV+cGt6qu9MqiHFXl42xJXc+yF0s1WLY8yjDf
8/PYInpTzL+nrdqArbx0NlcmCh87SwOCn8smGSiRCOgp+g8A29OV5j7+O4RrPlxX
+pVVOElb7iddwTVBGX7tP4tkNmdwdthsRbkr4pYozCO8vOUvIU28xjW5ZRyEaQ6n
bYIbmtUA4tTX4CZ9LHI3kQK6G+JlkFVsoRsxp5hqDrlkqWGfk3+zUWAPn2PKxZu4
FV1nFi/dxNcTOsMsZSGX5Ve9Q8qfnSH6oHUtxR6DU5i/zf8rhZOd5jzhKAfNuS3s
IxJzNCwEQo8GtBpNVaPXJx7S1LrQIqjcZ30OxsiW4knUBfG9Qa3J4dQUnYvOxVzY
ameIApEONqfEOwiU+uuvjH9KDOqlZcPegbH3fmOuRKmF89RbdToGqZHDNGPCqtke
jCzLlIz9NxgSdUmJG+QVLUAwvV5mmevBlFWMDDq5zwIjBkb5jVl3lD4IAmwg6q3N
U3WVTiApE+B3JfXcT4px4QsXqxT+94tgSFxiNXY+7u/5lCApGWosdxfKEbg03Y9W
20LmCKvuwmhTH3lWPBZ1/azjDySa91IEjkXKX+jOU0S0AwnuVzvDpF08zL2SAHe6
4VcehtRIKzM0mWzj90px7BC9iRmQVxwCvPilgFl1aRfpEM+HLQFP/IPnZSigNJu9
b+zdjqBcyOpNPBoZsKJ3M5ItOPcZcwD0tkEh9nEHKdEC8vI2eculG2Jc7paNp/zj
7j8leB1CY3/BZGjAn68cZHN4cBYFHvJJFMKlk/i6FRYpWVdtHzCOF7qefflxnsV7
GGA7dknVxoyIQFqOQblZg0FcXZdMieb1vW3dm+U4zICoHPZBSf7u3/LkiF/58CP4
fqOl4E1wTlGo7k6mXmo8124d6SENMMj79VMXsBNFWNbM1pbt/gtbZh4sgh3BlQP7
Ca6ueFTCo9Xk0AL+yHcwSA4DBVXAr2duEqpXWbcdla3fsc3TIV8nLsMDBFGPMHIO
PHyGDrp2E54MqF310R6zyNBnvesfhQMmiSFGEIwxGzemui1GId69vN93WnKbxOJ9
q/TzIkzAl5lPOcxEkmLDW9hldlL1Tl+kzrUSDfbqIVfqN+VhheMl6lT9OTTXD+X8
tNBL8TQnUtouGjk68ycJvOvn2YJC4cLifOxIytCuw5EbLoq1lKxZfP5Jj289pz7S
/eTWvlUSLpBomIlzHbkalEQo2oWpH4JiyOO/sM7slDiw+x5vRxQebX7JPYHRFSoA
RnLqENTNxivboTaGQ6VEiO6Yv85kBwAPbnQVvV4wCOeEnWJmPG27NBg+VbefTx0w
IE7Vveikoi4fzrXiyZeK8yEpR9Kb508tANEdJxPGjU/baU8zV9OCP2/7ZDq4pxJI
om9VA4AH3fWJ4iZG28OZXSVD9T9lN131JiQ8btwknayz9iQwrpwyLoDyRgEopJsR
AFPdGYTAj2GCfADCOg+HI6BQCS/pr5bmlzdXym6WmHIDJZp8SGB3o/Za65zFTAKx
hvqYdiaNLCFBBc6wC/0HYWI88kUw6VaA0hDtquHuR1EO1W3lfMQ69oo3p3Dn9gGT
auAepTd9nQarYKybeZqIuj6xap/2zKuYIncOyeZ/DXn9U0wTeiuXHXYIIUFBBAt4
8kGONUWU0uY3Rly4hwEB5YN1TmAcAqC5yfryKXuqKZ1LzyVlFdaf95ceS2QsDEdU
T7eRp+xw4cP0ZEoLX9FGb7U621B9Va0lkdkaLPPd+Wzg7zXphjV1Zou2ZEkm3iBH
JzlzThHVJPA1zVDfYC/VWg27Vo9kfVMG9YCpTekz1+rHw/HIQ5zryePx67iI7HEV
Z6CJ3HWFyfgDoA3QGo/xPh7I65drBDQS2Fz7iNWWqDXbf4kB8S2Oy7HVJlJ9DSzg
E1LLriTaG5F1TUiuzE9mJt+/FyxKzxNFkScfyFP6zbxtZQQWiNPc2KjXulpwUaj6
7fCrnpOh8DWOpmA6BxC8DNBpgxHzfgLofyXAu1+nd5ZX16qzomiTQMjiRq0M2kJk
Xu7ZcJM4tDRGItAD1KglNEnocUMV6NQjDl+HfaZe/FgDCEfyy4VeOaMLpiAom9Jd
HAOtE90cd/oZ2YQnv/sHzFtWmlDry9+0CoHBX1qopcECIJ+fToAFQaFfQQVUASU/
GeCLWG80w1G4LzROK3DhhBZ1CfjOZuHOWGdIx1owm42HkGbHeYRdlG7toA3I4iSW
HmsgXb46nR+8wH4I7EN9PTTAT69Nm7Dkh56DyLisZCJToz7b/lhoQZLXf4ytw1oX
eBWodzYdrcOzbFZniPwhZu00Ttyng6iG118Bp16uShTDTWQnFkLX0F+k1gnYlzSa
EEyXpIth7VLQ2cyJJqRwbgSJ0y1hPi+WNi327UKbQ5TLgR0GSABa7uPs09i72UYy
qBsMt6l5WB14H9Z2ZO/tX6ZEz6J+qzhUDhq87FpyxZ8BM/ygCdSC9Y4GajvSGM9S
hWW1ELihVTepQA27+rxfORmHhibk2DNlB34ussgyWN/L/0TT9DUUpd29WzYqt70K
oofsqSkoMNKfsnAOxFPUowKs3As/UCKAzbHUdF8/RzPO3N3DOH//qL2U7Vzy456m
xVk9M6vYPIGM++2x4oP30yf9/u4t9nmUvoti8CzcM32/dOD54gkYH6MOwwelICOX
7jQt4B92xsqj1oT+yb2qEv1sA7X6pI4wb2iraH8PbjcnLWquavLEAFE70SUHYqic
B0IAl7ewFIieOtpGylpDVukJGLbshrQUNVyhhKDkaDVFoK2OhsfZKO50WxI48hqX
ODEVV9oWwX0TQZ5JgbaRqLVEMDngicO9J716Hb91elimjZDMDMgKoXzic0fQSpro
f974i8wyzDGOau8DH/RaV/4mwZVYHrIbBGl3v58kZT1t1zhsej1+9TXRX3Hi71je
QkzApIu3fqkF7dWjLQfti7wvmMbKF1hBVzOU5f/X0LHq0spcxxsUiUXVK+IkhV5+
c9lg/qrpfTiK0qL3lTYSodAuXsw27FktcbTMwZD7eEPoX5vk+r8NgQ1BBH00aNbD
ng2DUYr46ocQ3kUekLsE+TEErFLKxjOtevMoEmeA7BTN9vofBmBezzQSM3mWvbxw
UMSp4PgA9cdfwUiWFnBnhN1WGfI2HnrPeXbNekomBqXmef2Yf2iF06gGS5z4E3+l
VmwLXpqMlDOCY+hssffKHSsrf3fAS0OOTs/XdgbmxBF8LHCkIYpTMuwcdoPcQr2y
4DRNTnPrT4JtBBL25RklYPM2QNftbcHnRn/G82PSeVCrX5sd4vIPph+N6soYdUER
A0JxVxGiQ6ZcMd27xdKSAWx6ZVVnwbWZJ/aNWlSbZzDugMqy24Nac0CWoYbxyxzw
RFgr8H828wbL/aFFjub6s4YshNP2Vz6XsG+bHfeJKy+iS2luWdSghMLl4NAvdrxw
gak0wieph9+unQUo6hC+sRZj6RyTSmn/OR+nSNK0q2Z8rLnWalWiqYszLgfI/xDD
/PGFuqCrJIxqdWZ+PhuiD91PuAXwi8jCGFB1kUouJI/46IygvEpXVS0DZfJtHuQd
EXfGzkyfob/D2/p1ad5fIcy8EoSF4NEUGrv8afsgIlsyZk5m6Gq4dh/nByCU0PfR
7OyKdBzLvNGRoP3h8/HZU5iMXkBjXD8E7F/xGXNX01U446Hn8UPPcL/iBZ1CCvf3
2eEeBD8n9b/To1GeIB1QXRPBEoqkA1dzgBUoDRO3EE3CLUGqWfFcWYUZ79M6V+5A
XBx5fCsAdHSojsf8Z7lWBxfDWUzfdPDyenG00xejMOXllodpDgwPdBiywYN/Cc/n
ha6h9clT0nq0WMMaA1DIHJsWV7ebnscHx/v9wBmUMGPPULq4W8KQyrMPI+bIHKZJ
stcuSpN7tMimWpIZXrh8vj8Bva004GBbqsE/kYlfN1JzASa6nQNXQNTeQKZqoHjc
aPwWU6lClHde2D9uu2fxTnpCnTVAISZ13uzJWuqb547a4rESebVdYNt7bCsSbslw
DyBzxyl0kkmXA70ixr2sEuD3cSs2EQ3NlFiO130X8QdueYZQz7vQqk8SxJmIUbOO
4r37EZBh6GAj5SsVe3zLTdxYleZ56JrltoaP4hykjVpCDkZmkzbZ49qJW40TOMTa
RxNrN86fVnTYGpPn0H+UcZM23p8K+DAbV1gQdi9V327/voHoDusxpDqfdqyPX6aI
JF9elvTX0O9zo1d/NydGVY/cV3D5jMm6/jZtR3OCJeZcoRJWPNR4G/SuAy1VAJEw
q3pb3tGWO4RTZpAixfy2eUw9OIBxnhBLZTWrmvamU9R4NxXHEXpV8iXrpeCAJ/PB
1e0WgUCnf7Gk6C3tuRxlDyPDiBfHZER+WlsQ4Bbzd5TTRVPFhDxqVVkH5jYw3lHh
Kpjd+sgfuaYyKM8oNiX2lcIZEVgZWS7YEGWGrDmdhjhOaeTx3CSfjKktpXNhcJz+
ArJZOB5zgIssxRV+r0XkZn63eW94OdFf8qtS/DjXj8CIbyS9ydWgrHoK2C19VW/3
0308Un5aNk2GeVVLaVxZamC+han8t45xGoyafb9zrZR6jkKvftp1Jj86Zl2j9Aua
IbZP0G6ucLoZez34282MqLHK8hGKPbXlKgrHsRB/4XyeV5pLx3n1GlmzppmlSiNB
pu8m2WDT8ECqP6mWnxR6mS03TrtKnmCzwtiiO6RcRkwq5Q3RsY63uvZFPbtJeprk
yylP67Vzk7gRMTuQCH0R08wM9Ua35LThCUjE1jdMhoGgZFrP8Juf5bhhUv6p/7eo
DRUexxOghU6hn/kzm3qftunO0QYAYA4X4vvVmPsqJWXMpU/KLmMqsi4WYfbRyH0Q
QsGz3fHQ2PRJEI2SYNyOyfNr8IjiaPTPHeLnuNLryFxjD+tzxB7/hb5XDesW3Iv8
qTCJCDl+x63sNWsTHZb5nS2HWOYs9C4I3fn2/REpDM/Vzjs6ZTIWqrxspkeZmXeA
h6yyL5/vaTJpdMRQcuUIgIRVmzA+PqGO6w2pWBWgI8YKnKYePpwEvsWbsCY4yKkb
4d7gqGGqGXjzxLoa94lJn7sqaPDhDml2XkX0QJ+H8gIuIxkztKj04vOhLOJErBG4
E4GbKSAQg9px4vR0F9lnvGBDRrxra1XiyAAhGTTnEBkU6NP2Df/EgRGyB0b1kDEP
DuOiGgDT+Sw6ATnRjRVup/PnxVOmH3qk6+wZzO7OFPW2I8Za3LyT2Pi2duDnMPdJ
whUyf8CcjEa/5l7dHIvUWoK9fs9qYRLL2tWZ0wjeQY/e7QFHuIDaPajJrszCdL1j
t2jhQSyPeOZDwOFtoZ0F75n26VXLajNSUgsjW0fA2C2t/BeFhJo3JilHLKSRgFC2
vvizdR3lGMsmTkCHssudAlJEWlc87JnBm+WsMsDPDzV8NeeawhJ0pDYcgG80UwoE
z39J9rSA/PQdAl2yRd4GBec1y5Y/B3lwijV1GQDeftvpUHLvLp7JEQpp4YTgzl5r
vcuNNjyRL8DvndhHIr8wfOFghAvTLKhN+3WPaFCOYjRlU5Q172JAH/kPNCYqMmJz
SMu+yRUQFsrZKnFwR0AdpRKcj+BsDUR/Zh/4fwSDNLI98/S3vQD8awTju4VNd0O0
2xog8QkTLfGa+jvY0Id0pVKcffF0pK1Fr/NyhhGw0DMFmEUVk/+MsOmrhWiOzBTe
DtuUq4mMdDBfWCDeVqIcA1thClCiu/IgtRmwVNQeAqIopGWZomuQP7oz5sKQduHb
T8lqKO9i2RVIijnOLjxEUl8FUuTljWuF9D0M+3N6SJAwbNs14dP0VHCqp5CkcJ2u
KTajArst0QufKJOzHkP94j7ylnlRwwLGK/P6j4Dahk3w91ttC6qAC/T12Vc15mpN
Q6w9CdeDqa7hvVkPmgl7Y0ETFxeFlERoSwXIxa5fpcBTVlOtNLmjjy7EhhC1tp/F
2Lwo5WBU4aGbjUACQnFQs1uL+P6ecICZ6Mzyp0RxTz/FiVj1RB+ssN9CCEkto0YL
207STp0ORT1hQM/j1i4uHJs+ZpT1orRWt8i7dst7nDW7g7/Q5IUmgED+aRSr2TvI
lc1x9J/TTvsRLiv6V9Y6mUV74krYwWmSb1+/BIVI+/pEypVxj2SWaCGfwj6M/nV/
1yAbe1+8ijTe8WmbTIF0YFdbqBzJTIjHRU1s4PYgTYmUbTyHSos46KsueMUX7FgI
nbu1Vp5eykAWgPT4838uftlxMLV8UnYA9d3t3/+yGlWlzJURVqLoony7CHUwm6SS
3I7H19KLd1UeAJCzAkGuT1s36ChZ5vfs/phzSjAUiImeeUClIk/b8ezjfm4f+wl/
MX9IIARAiY6RsyEXvWSniDGe2etC8JhOq1JbG+Vi9yGGP+nzJT6YxXHhAKnRVEvK
GwMrcp6yafTpMpg1mq3Y0n+Ub0ZAkY5wZ7LQYDIYKR7x1iXrmAZ1a2B5tP770Fgi
QQnLxwRCdZkmbbSzrVOpoEF2wJTVOO3LBjMMrFmYo1g4X9g+3xwQd/ZbcJCSChsA
p4zadXKrI3b+RBU56mpWy7w7IyucwZldaUVBwt6KU8nf0akMitAFyGX+cxDBGt2F
+Qg0X6rvAGxifk6w7RggUdUz2Qip+xyq6wCR8JqBozGlc7mFWXg52MIuN/oZBxfk
jJi7sYlh3ubAwyu/okVfVQjrXUJAwQ/8kGgNeqkSXJylp4dJ4k4yCjwxGDow66My
hjPbVybukF+mNadTYXTkgQPJX42KtdErqkUJtFfkzu1j3KlWXwUNKLUmcvUm3FZQ
srJ1xP66s0wiIxpLRdMho//PeT/L1MgYSPdLbJWCVHO1chttJRUgLBx5VIbPAO1G
YhLIETNz0esfit9QD63Fa2jR2I5uapBiZrcMwU8m8ubHrrKgVPXMV4JBQI5cKRmw
xRlk/Tq6QCQGbCPdDKw2Vuyrr2AN0M3DXbqzTW4QVcCe7gBVp8SGAXfHJqWwuHSp
Urn/sXHJtGLZSl+hz9ETnibHWGVcYeqRSlI4VxI/GbtduVOahAV9QZf2gKRj3REK
ZvzLH7JPynwEdVr2AIrLBCdOJ2AGhkUJdKkctOnc7ayxj3I0mSVKe0AwNMRahqfq
MZT7DNCCKk1Whw1RqilnrVyK5t25qtmzmXtbJQihocrOShKLRxIlM6I4s8vfSLTs
K8cPW6g2Guj+HCsIAjEKBy2vn1CP5N1egLr5X9K6axqPMXdLRCcmrW91pArQWXx1
dLZbe6IwmkD2EDvf/cc++9xSOokf+qAfljN7jVVpC6R0W70k/BKBF2G9T/pP/c6J
OquugH3c9RKOSZ0L3QqFvu4X6k7ZENgse7eCuub+l/nvw6dsJlsD2khFBK+mV/uF
uYhVL/cvnb296/ZZxLXkzPbwCm9A7Ctp+/4VYC6sjFvx9r/lfaoEZDxvy4+Czgpl
TravJwUCJoWOyDGynaVpRp0MA/F3lGQnlphxtz4hiP6Fj1wnvFejFSETkNgjgDNm
wbPinkypzf7YvMtO+ZOZspRpctBcqjyDDuC6Uoc8nj54nqOoggpKDZCr1Ck8jctA
P+AHgSNcN/lKoVUZpwheApnhlKWzRgWAe8EJDkUGdESjoD11Y802OILuxzvrZ5jS
L5uMiQe1xk5Eql6UKezPnAmIYUFemIhTaqA4rlIHr4zdPeh8lBkC1s0Tr7BBmanK
eyKC7torlMQnibRB3gy3l4rdsGjCHuAuKttNwtuvgi5G4PK8OBsFJgKq4tZSDr1P
ySDo8xT6K4V+eD+m5VldvQNO7Jkbbmpfg/+exCdzrc7mK3/Qg1iAtvXqDzeMF7kF
4FPG+ygeBBCTI8w7gBOZEyZX5Qb33zfW7arPm8hUT7oulKhzUjS3x4JVqQxlHzQ5
81HeuE95e24Q+RzalE/SOiCoLQIBpRfk+2sIoxxkT7Wt9XgKPRqlTUOySS2OdX8Y
l//HkQUWY4DqGVhmRQ+392ON+bHgfPxMJs+H6+iZeCJE7gUUj6dnZ7TilA73JV3k
2FGx7CmZL1IpSP6Ni5EPUHhdgbuNr2N0e6DUs0oUlOQRLkKtPkhxhQP0waJ+wfCa
ZBnsaBLuprAOkbLKmKfj7Ga9rLic3lqJ4/h3J0LNOHHTFLDtVdx39Kr58DgDxVKS
dEf1Lcan9rU8vk+gX+mFbgpqV4Ob/sPwOixhpdUBO4/4iQmt/TSSpX7iZXOq2wEr
onIHyj6ua/9TDmpblHm7C8lZB2VOeWnp5fXLuaXA2wWuDuJBzeTSnpfpwJVqXLYH
lsujL/xL3tdrL1SvuYKa+t/e5u6f26pnewsDCGdvKocKLpN7fmR4sH9wnz25Nhgp
F+XkiNoEcxzk2lm2ofuSEKnxU8V+TgAZO2g6e6FDaMTE2plJxDTAugi5k+sHv02Z
BanPzVE//g335HUt5ds47VOczKArhSs+CfXxE4UHny5ryWU2OC4E16civyDWGUT4
RC/vR01BD/vMEi4oETXuQ9cETD0BRl6xHNihVt3DrcqfCj9mGtfm5qST0qm2wE2T
XcG34bYF5FsdwqejL4f0Jw9SagUs//+N6Ja9rVMC/kNtzG0a4v2oMqUL/24wE37/
UdwhqVPQaRSty1tQTj7WgrLtB0mEEzMOoDjs1HsUBzulbgIpk9UND/6bwDK3x+54
yLqAxWvKt4+jNCK9sryYkKqwGJcDcQxFk/ioCa5VtpxUwtq3QGMIkb13XUjDtwy+
VNqJpI4QjUqqMAvJa7zS3TSnOr6MlwwCgb9AMqpEzQw0KtyWVcL9JeWHco04UMgl
VStTI6YhXatRkVnSEBx/Ip7hbrjtfoxshmh9KoESZRs3swODiEZc4LB+T8DgKPCC
6ngNShklT6fHBrkqBMh94uGbpWZl7CEAzn0Mz8CLyfI8u8bXlxgKbx/BRjn18dY3
LJubXrkjQMTIyjTmkkiqgvnGL3K2VP/2p7sNOAQCsLNt8ZaToPpMuf4cvD9EHR87
hEgV5FJJvPwmrt1WfSNTM6Rja/Lb7z2AcejZ88lmY+AiKlIAHoLIDBaCr//NeI4U
n7jeAK/K4TcteinPugIP12oYUCBoWKnko3Sfy/6VxgzViTzBFtXKuwB/F8ADu4JG
PPgD9Cy4NZlYTzKivAUM8HvTe0aVElBtdm9CfI6I8GXrfHm2dAH62/U4LR9zDAuc
5pRScZayNKRWfxGsZ+4JYJs4jktmke2abR4afB5ll7ar9e1Nlj3EZgjWFRnjP/HR
vTBPg6E/a+gpU0hrU5n8bHzGzbi1Zj+eH1ukH6EYwzPXan3QHz2J0eUxLXi6AobE
RztY5Ke8GFBZOpfvhFstEL+XiIZ5qTKsrRjNb2GFiTm9mMmgxODUAM5sxpj14RXo
AjTabqaWp0sSNiafivTJ1+f05uvWe9926s5xqYSmEqsPUuQwJUegx21l980SPnyx
WMvo/DrWHUvU+VpcWYIJ3/ZuIiI0FtF+Z9YnHWQlOCopKiRIyX1X2RADCWSQXw1J
1xwy7ZPlQHV/UgxU2WQFVlr99QO/POqjhZfh9jzLU+fB5r9YG6xmr450mngDPkxS
Lc1itj0E4ngBFoXwLeTUEDYOjyKHLJ3YhFtbXzJY2bEU+joGWF3jmZ9ICs3/6iHn
sBtaRvRK+r+N+z42pRuzcUeHsmBlgKE2sy+ezH3frilr0zSDVnjgEsxNZ5njzAYW
uXNdvU+eJI7nh+LfMYltm45I1oDVxzTUfJS2mQvm2qo+7vjtFEeshPQFFeA5deOM
xOt+MCvt5ZpMk3YwK3WG8mClkqQc710RPiUF2n+jK7iZ7LfOWkucYRIKQMK7vPjc
OOuvW3JcVb26XJEh7cJKexCrT5U6QBqVw8HF/beiCz+jx6xnzSuR6U82ptH5MC2x
ybwMwCrgWIuC0a0rD/9WHdLiM1vJsfSe6hR33hMPNOSUoDzMMjc/EHeHd0xdc8LW
xU4FOj/MVGbNH4luxEdMySxxy6pmrTizDlcYIpx4HvyLfdxDW9Cf2B9qblH0dxSY
yboMB8I5AaebKJg9zZxtEETnvDdK+Ml822c+mZIuoyER2GnvjaZDNqmjeJXZEzXL
yKDenWR/lZZ9xVP0w0n6UgbwladAy7rQpiQPGmcevf93U66VRoaZwTGamlhWgWrj
Ht+ARMg167k1Otk1ti2oUnSeb55Lt3wE3Hyp0zIUvOinCWctMGC9uKynfLRPl1AQ
XVIU74iUI4OjZT2jd/i7fZOzmrGBZJ6ZX6AlOxMv/KX22aNAQa2k6CDf64ToF1iL
8nLhh9HHHqOEtWPOPXILzeEeDp/+RYf3LZe0Ls85ySuPJ7hYqFuECrNoNd3s8zTU
KFrpULne1xn0kQF19LSHn/Jkcq/qiFoKHmtkJ7h0l29k68WgwYcgt0I4s1C7h80I
0fZB0bqx7ACLX5n32cMZh7zyZ/EMeEk53LK0wetD++BOJpu816Ro/2UAkpkVgQ67
BAMatInSG0LPvzo17PDO+mgFiUvTJ0N4t7mZNik65eh1AbsddBgdBQ8AMLZuF7B7
l9YVjEp3k6z+ogUaPPS7eqKMIVSjMhqcSxUkLdlrRrzD7TUhiieq3m8sWhdS6B0y
W7Wi79RXu5ctyfRtLJOv2xyQYRpAFU8if+asRunED+3luwNbHYk3jV6BIZUnOb9C
zIh2M7kXUNfyFqwCy45j2t/7R1Fn+euJHfrirHMT5ERPO1jN2gDp4zzAAmPavchR
5X1hEck/9cp2mkZyR2uTX6wzrrT7bf1CQAAMt1DbjRhmI6xOtmohI9IHeiezl5YH
SEnWChWOklW3seSc1ykFcCs5uv/jym3ODyWSJjSy9FpmRCTRrujhmA5K0np9THTn
ej67e3uOsan5psKd6XeA9Z+TjTaJ9Nsdjmjp2wYPEdS8WOIa52WfTz22PWqrnd14
n1zjXATBQNXl+wf96lUB87EoKmh/grkKc0TKxDRAJ0WRaqZF7jfSJwilObB3i0gP
vvCkygtXSr6d3S2UUDplvCZjlhQ7CiCkYg6pmqmsRQYDFArpEs0mqHwbAizDneig
1PQrSUQfaRV7eCPHTt2RSKYGLrsHUaPsIGjbOIaRhqk9ouwnxqUwU+/PEaRZ57b6
0jvvksezYmCBjZwxwMIPD94RFhmF4j3vvz7vY+8EYNG8FqKvRAEhP1d9BJCraUtF
kJ7vj+MN3s/oLo8+bozqyif68HEhPyO6rttcyRI4zfjZkWnkGEcqcMcBKOc0Mho4
irw3lEDMoy4LK01rqPESy93UVQWhgS2X/A1Z1uAi/ccpDGAZXD8kabl5EP5TfOuV
McxRCYuhIMZ66I1DYaqME4r646mf9vKXnObybLcxHKiNqhBDq/pzP5zRQEqXFDzz
ztUdNzKnogJM3KbJl1HeJ6wSmXL2e86TsC3UJNQc3rLWXT2VRaoj6lUohrSAUuZd
UQgCfaWx9Ra1ExBiFi4Dtng/NxpDwU8axfH/FtLbT2Wb447+wotgGkFucoSqPXDe
6hbKQLpB8pQMM69SHMh3aYsokwoim8IFGkklBYWGWvk1VwlgWsmna+pB9WhmitLE
JhZo0ruHdx0quOnwx4U7QuC1Jawtx7cOG6Ag/2gaoyg/yvv7HRNzwd6X+Iz40BPX
pbKgSJF9hkpasfedXb3v9WzFHZeg70gcNvl5A3xQQCGXIof/oO8ZwgWgWx6OsdkC
YQeZw9TH9OQ8EMxn77SmeaRPXCFqCXyeUyJDpD8h5zz2S7PYeDMoiCRwx4G7RUsC
2j7QTkE9FcxU9MNwxCuCAt9hR8LeHpd6VpWtaH55HxzaxpA06GMM8gxUgDbyH5BK
yKE5/BfHFgWYS/YvpR8gItnrqDLlobN3Y4cifJ85fD+0wDfZB82QeqWZfsywYX31
AHVFw7ZLEoMl+HuqoBeHYAwIMY8e6JHfxWbfgBUW5bN69/Oq7IpaZ8EoC3bwIh1b
lwTbVb9Wc0ChB/OnDkeFD0gYSTYO8GzFnAzN2Hsl6K9Uj+qMa8OanDiKRUwrSFhi
WRWpHMmKcAFFjt2B8tjDL2z7rVkq1wmLmku2DjyI9cAFhqJyCxZ8bKxHNUC7gyz7
ue77pBk9BLaqe9qv1oemeVCw+o+YXTEc/BQW9j1UNsQLDPxhPm57b9RsWSu/GSy9
x7pCqZMHphM5EUs1vnK/T/2rt+mt6gLce3vT7VjRz+luauxUiBL5gNeJPxACSXMp
cGZJCb+55aH7todPveNGzgh5HYlzRx7wSwlGJDyFEntv9Uwgo/ykkjNu9wBMdnHY
GYGaEl3Se1YbuUlibEvGgz55tHqv7/PV9TKvixWdmPx03DxXxuN9hY0eaSZh6BXa
djNwtS+FXjB3zHh92UbTbtli6MrD4NUjv4C8Fi+Qf3qf5VxRAxQKJmJsZuMbOskt
tcspeeSB8KH/6pUl3BARNebw8SNVsoyY/1Q1Wy3No3FUqkmO3PlXcCvdaenM6fpk
TqV1noCZkk7UFIn2UsViVyJCxv1xASCx8JcZdeReYr2NIOPkMm9hSNX/175zk4cC
I/ymV4jTs5REnVACDk/jZaaIxOK3cKU180aJLhSpVWML6iqvIqtDaQl2S5hhqinE
PShkD9616Kg19zAP6AFc4V+zfaW61DfzHH4pDtxNbtnsnVWt0K+Rfgbyo+Gyr/cY
mNLnTwq5X+dUqWHQavEqX6jVIBY775s+2kRdfgNm8L7dGtQb3xd5CEIbenG8JfHK
WL15+MLprKVcvyL6MWjwfjO7mK5yGMLiGxr27kPkXbHlGlzsb7kbBQSRm02lP7ed
z312GKFaKf73JIgSso/O53q4iYumIK0x61Gm2XkstwyIJxPQHkqfPPcM5RzbbdwZ
gRMDYI2dMzhMaEBiSrNjdasgXmjgS8li9TjE++PmZKyuHtrSybi0pKDWKKsTUWr+
op1PADGHF96YFIB94BXwDzRxE0R6evCpUxM7HV8x/jX/jASeRp83iRZuf7V8cnuL
ObHkmrqNsJE+XoD1Q1mE6xiQZ3InryGHrTndnSgxPNlNrQan6t1yeHQCRVfoFH/h
x/EKRkdtqhgk8Pwn6kSCX+H+32F9ECk0lxkFKFhDJYRAXVEA4wPzbqdXPqAU7N1K
Q3bJgLbfCXzifQRbxXBGgJUE9OxpoRJINSoFdfekTm4x0+NdXo9FQYi48rKqYLJ7
4cBZBmhAMhaw+n4qaSdWrdIrswyjzlPybrlMeBg9kCWijPfTQpr8uCJ/lb0JcuyC
7w5QugLBLjRegOvPTkaZozoegmrBM5kZvcohWucacewqdmjQKQYflpqtvT0JVsLe
exdzGMBlh2PuczwaTm7i7cpB8AIhBONBmafa1IuIYf4nzwIpfzYIVCJjNwsavms+
kTvWSIeY5YUqD/s+GLBlGSPioSp18CQHtacGSiHWvY5a3FGOCicDcN9SVHHumnqP
/ZroobiOnluTa2giPY+QyMPqDG5raAl5CfhiWNl7KnQ8yN0ufvkasi+qQCokXgsv
OIPgyrXloyZJD69MgNv7H+sGoC/gChF+KnhH+yJTTlOeBtfO2boMc58Mw6VjoMqX
UiE8UZV/gpyiTyurIzq6sHL3kebl1cUMBxxA+chCfTE5KfQ5gFrKdsVaJ49sve5K
TG0BDKv2B/J3t4FXLM7ljeX584VWY+qmvMgP+pIEWC5EUdeAj84y0fC7vLKuntck
3DwXwL6y+EAXnK6Po0hkTlA5GTma1o0Xx36fbN3g5/Eg3aUXDSD56bxnycV2pmTX
63qrxAmsnfDF+3TPEUVfsGoJtVaHnee4bxBdYS3x3gz2A6IfGHRx9Iis2IHTuH5F
uyTOH27LAuzQqxEd3/2rgsoZFJWI5hURi6OsdE/qPu7YsTIYF+YCuDdcE5LBHkeG
S7MQY0Py/CZjukkv8K3W690WF4YY24hHtoEpBih5Eci+T/3onLtFOm36rKJX6uAK
MsssLjAbGZdS+rrfu6KAjGJpT5P49CHLu8wwtFOIVJzHtPBb6VRy/QV4g9S7r6PU
eaqicOrtOb1KKvHOEIRi09uNfMEZVFYav82+xugSHPwGd8MzQe446M/hsfyD0/tC
fsxGyZi92Haecg1cyQ1vsZM23EzJqFfN0NasPICjrbnn1PGrhafcFBNA+TLkgKMB
42omI7NhoLhFg6FY5azSciLqLn8hyo3vm6r9mGv1P2f20cm+OBVYKZq9VuZh6h4R
Xd0RCPycfDP46b75E6zzg2PZNlvS4vh9WJ/ubNXacVr/aH3fWze2NLFqafrO4She
+SbP33qX+qjvFbSlI74t3+WXYebmYCIVxaoAJkHH19WTi4dPRcYjuAP+xA5tEzQ4
N/q3nPBjAc4xqvFx/ct9EoUAJjza+bBsghDRZxwlSIyySDQh2lUCUE+/EiKLakxF
l+8M1fqlCncN7ptGClISOOvc1fWsTZVcEAfPe5dsnRZ3ma/99IcTkR08vO8k7QDK
RwJkKnpAak1dtl+bz6F8DEEbjRgGIefoSP+v5LY0XH8Ha3hD0aujbFtwiF8swVg8
SG+nb6uvSpG3IDjhIbOKo+y8wDB0sxO/VyfQcQ+xAm9o+Fwe6d6vWs3/TSooFUwK
Ut1rWnX4yqtsqKhVSoC2YzByhscQ3/e1dgj7jHTnJzFZxYngZ4KJ8SjqkWPUQGvP
QTVAZ++1lMhO45r2wYmSjGrv/2Oz/4hkIi8gD4OAX9UJsFXO1+dv6kC2u5eXhEki
jXJFxW96BCBB/DsWBXtKv9sO5KP6sgL4EiLbmYF6P7sFoc/4Tu+1hCK7xSipR/ZA
Uy38qqdFZRZR302gU5azSywyKGfu+PDy24c7ADW/q7h886HLQn+qKa1ieez4O25b
o38SRMriikD8n9d/H3cVsWOC5cVorXslZuFUxoAPR7oF1xU9x9cBnVPb/EdFNEY4
6tfUldjuR9iIQFqK6clfUxEM5nPqrRWK9dMvKPfZICH4vcFpumI25MUIVbJj7aEJ
qLFArhImotUY87XcMWVXTkM0pg2dwuybZhPFHZlRB4OxXGvvtokNIlTunw3nuBOw
ymZCOyfvWgiAvYI2sYjw6H5GH/yLiL5xIJfd6uVKgZB/TFR9v+NF83q5jBdlKw5w
bxF659kqSJ121o7Zp9juraAJ/zBQZnLy55ZsFoDGqsIrh8WRixA4G8nxHnfJ75pL
L7FUg6bDLiVcUlzJAN++7awOkNddDkAlKPDNLmQxHgBXW9jp4utvq5uF4aQ912en
L/mOXhUMU2I3nbIBGKEncD8est463WUow6NeMXFvN/CndGP8KGl98f9iVYBCiOIZ
3Gzd2nix4Vy+5LSaNRxx3tbcCOEKGuHtH5ckO8mIZNf2FrWwgubeTnx1dRVeO+s9
1pd4tK2CJzX4leF62YZ1apgNSBA3ZkeCZiTdxIApNgjo6h9o8Rl+7jj0EVYeLSbN
+h6sFwbiwYXWUl1FK++8uah5h+0OT0YMt2hGXt8kFvmrwXcYOaAI0G0LZTbXZ2DK
ZQ+bgfmxy0x2JrVlRNfohXCbA64LwxniXydIZmk4PwT8EKYs/QU3PCT3zlL7Kxk6
yaonUuuZcd1ylXR/3QPAFIut92SEbTHJx/MtnDhzUunQ4EZ46c7yKoKfUmEaj2dK
GpYTj2iCT71Xm2F7hfVV0qZnxi2riSILOT743iboJ8HfTSXMy8rk9pXfJ+pRnYv5
JSdg+342Txyq+PaCYyspCHeN5KT8TBgN4JKPB8DObfFwpzi0z+KB6oDTalYiCeEZ
DuhrFU8Hv5XgXC+jcG59BGa8ybY5cY3WdAgi0K5ljcLb3HUPAA7OLXjdqjcFZZHd
9FE493XGQj3ulJjE/5z7LMKYhX7ql9GX2KRWVFtzeN+sl4EAJkXA7bCc4gw85uMJ
ejOf3ZZ8XSuMxf6hfXslHWRXTvvJ+8D5I5abTFIqK4HbzxrXJDyylxq2UItRonVS
U7pTXAf6NdgViHed4P97rrDjqklIfEUarJFomeV6A0sd6PSPBFPEegiwh1Uesssq
NnJb80wLVTN3XEK1aSu5zCuJDE0+HReHHCS3SOSIEeLt4BHliCFrsB5FOiE5pinn
jmaoysyJN7RcBdpkMqT+6KOOmMFAx7AhBFRl9yf+npDF1kekdI/F5Yt9yLEWBu4h
sAV1Qa9SQg84EVJaLErqLh3fxzodkUUDgBHYRa8KDBXngdcBra29WDz737tONDhv
yuCgcLskR+epMHVHbbqhjv7NA3cKHoxt2KMnd7kZ7ybyrAb6fed4ikPpAungpl8L
wA/+Rym4YRym+UXYVmrs8IDaxznByJhLz+TiCM5hLy7GMGS3rA3VB/h77i9ZX7eg
WHWFq3GEm/myh0kwEPPfW5R2HPblKj4UFa04lrCy232OM/nDvOjbpMTOvuI3WV5n
z9OMc2Emu2GlQqxZPaMUsbP5g1TgNkaWBYhPS8SJCeFXYsK6A0uH/pcjFyh7aaWG
nXggZ83BXZqRQFGUGlRQ7mc6lA45VyHkcEba9602cZjpdNR+jEA839FmmqusKW6y
HtwSQauITAK43Lubl75l+DZhhB3uFl7qKR/Nbpxn7usXQZVh6i+NBk3dmcUxu65T
BjtCLwvZ8umneg07KZbRacFoKiEHo/KcZgckSo6ug+TlLF/RNWc2zqx2gnvqHK15
lj/1BzW79U6kvSKMq1dcuAKuUavGX0/WZnWqsDPjzJfXe0N1Zd+MkGdaK7Y4iYqG
gh3EOynLiA0ncPbXPf6lq/2leQjTkEY1XMOtuSenYNObFUY2QxXKiHgGpZaHe/TI
iggySJ3G49rkYJ+Ow+C8+I7h5+BYgX29yoBoGYwCruOMXagNnwTesY/ks6NOrA+r
rqfIXXAMKa9l5bdbe6wgpbuVQdMe1neDfCyayLJbBhqxKpdW+/IuPUCPKPsdPChP
lJkWc9/rCTDKMdyhaUAqo9giVPfJufFBngpa509YwX4fkYnM2fgxH2dCchTK2efV
og13rgmzJWivHseYFxOyb2PoAg3MQGzu5h23sZM5LUS91FCKWA6rHYZZIOY4iDDy
RJLCZK4sOXyRH/VsJLNl40Niap1W64S/1wC9zPGT5d0Kd4dsTvut9gpu9plMKcBX
Si2poMeqP6C5qB5u3nXQoOPXqIYnEirgnZA7Paok3vXwHCWlu2dbsWLbXfnIuLiG
9mRHpC11G2KmKJJPnaZ9wM98LYq1K+AVj8c0U8VvEEqRYEOMM0dPtNRqccYBid1k
8ZcFdoLSUqgJkoaMq6UqxmPxu+vRLqzNUm2J5HmNaMSAVrbA2FaTFsjKV0i4tMFR
Wsrbv80bUb9eqhh1RsOYfkJrYUsB+JqtND7tGR72G2yoF86a19qN9GdCnVBlBnmy
JBwq0nadSX7AasgZAibxyYgB/qk1O3J2rKqeNaVsCEuOZ2WP4nC4nBy09NetsSSp
XPErwC6RhxU8OFBAMPh/9JePPY1q2+OlPLxm2/XOh6TP9ikAyygdYDS8gRrda7u9
EdGP1vm79Drs19xNdJlqGSgEPCc40DrU2qxr5qr6dZB+aH+ljQKmb3WAd7rxi0vk
/6AQwHOdQn4iowkKLsgoXkC5XZ/RPT0Cf7H/shfuFjTPhCowslI+/97DERnj6f8n
EadnRMe97AMV3Gp0xS64tr6NRqGUK/vBsp0hbWcA/0zqIcjOf5rvjxL9byHAGap1
i43Rr6oKu3BYZr2i+rbtIvic3o6VbIkEFrm+s6K6F3XCfmBvajvKvrXRAuHuhVAV
7RnmS9pTngad1UNumV5qX3BaaJJwTdK7RXixp9Of6EcEti0b9hQbZPrc9jRCBFGP
tgzyd/Uey/wjVrpgKXBXZHdpi2FIJ6GtwlMpRk2GGdSWZF5hXWECJbtvJvmTBrkn
147DqpmdjE9+2oDGK8+JWDv30EN9HQTpOBni+qWRW+zq4vpfzaFLIP4aSdMCVQ5A
LYrrr698yJ1Zsr6YBczwvf1P7JtLbMjW1fesRvaHGneL2hu/T1GEvDmunzqwYdXC
mG3tKWHQKjBa2Vf5xd5+QInTLiIWJJQTGgVE7LkuKDP4hPbSopJdhsrcew9xv+Qg
Lln3GJ2TWLPL9Q+bYPzLlYFiqpjhv7UdOE3Lyc1Qe9ftbM7v4YQo2Do88bG98PGj
iZOBarOADvpzThUtjdt1DCQ2zc2DMluSrAvD3letyUGhk1DKL4slEKQ7yKiJ/U5l
6hjECFIUxICco0v9Bst8d0M0owGc0eMyxk6FH8phV+r/L0MRpLnjbPlLDwNfva2M
Zmxn+TQCzzBTfUq1Y1r0kWXjW2sA94Qawco9Pjc/V3g7vZDp+/L+NVOifLZ0VOcz
F/jLa/QFkliJZqO2DCuFv7wqulWXdJu+x8XquWwYCMBxZ0cdJCHW21AufmYarbJY
Dpw2JO9zqIDo5sIfrxkmAHfra7KQXSEYq/aM8yRZfx5BikYEMXGwdlTHAF4pgFGn
wk3UqMPmR7la3xqpAQMpxW0GzYusj3HnE80UgChtQK7f1wGSBbBkgjnFUvURV+ff
7h7FC6CdchJmCY/r8njHP783gl5SQmOqdC3z4QG8l+W243tEHQgIEDHJfSxirRY8
fp+ex5SHKCcRMxSCdf+mTVpmGEVY2V00XpZKa6f28VSdj+x0fQbJEtzOaehKk83r
ZDj4iXKdqs7RXmvKm4S//YdF2MnYdUAMRePHCjbgxzgM9g5v5Tp4XSesrzCOpmiC
IHqx6WlLCvUrwjcArjJNSgJKrmk1US82IP5mkZUptzllF4Pun+VFwseEJ7AkdvrF
Ngu2N618pUf0ufbsLMn9FzEgad3bcpaXdYhL/aI4+8LMmR3S1sjnmpz046n3mVwp
t6yISqWnJOASHXwto2E3AetgFCqq1Wc3G4Vr6yMJBZb7+Oe0M7QZiAa9TzI1aiRV
gvL8wMNsBaCbt4dyh0UBT2Ys4ixjfqXcDO7YHkM5u0dguuQzSq8csCtg2Qc8VxCK
K0l5MElsTGccpPd8zDuyLe3EGv89h0/zY1D2teszhd6gu6g0ZbyZ4pdk8vITLo8X
jc2vUYD+xUw86P3z4Hdd6SjTI8zXGTxA2xv/RZ3adaOsSReEA+K0OxW/gqyOEEcb
lr1+jNnMRZhlvP4nIYCkF5hs6NEmnIIa5OrS7ojWgDMjQwPttjm4p7IFPsGLjpF1
c9dOSlVZUsyBhpER9/MiRSKRb1o+0GjPevkBrte5prMeM25ie+YNQNmY4BqiT7p2
UEWeOdN+lCkJcM4od/cHDuQSMd1oJCkD7IwK//QQKTXToTuEVfSsP+Vj4gJ4diwd
1/7A9V3woialmMtopAw9xbXlanWhQZr6f6qcaxlyCzNmN1nEVSX9nEYpGvAYU+ug
0FXcv4iziEO2lWIzbJ8KElMOWqCKmasRHDjBQWSOlWG5qrCi33sS/1v7V3n7sbbD
j8q4NqLzuPRd3b/0QospL8W8LRm0JVy9acYkGqW6xckHcwXGO+dDXeYGCAbYOyOo
xuMbDNJOB8yr7cTxySSpBTzY7B/pEmFL2bXIqVGWEWFDTL68VKYhCh0ldxbftPRK
q6z2RE11f4ogu3zNQ7TgIQfgZxBbNXbJM9EpRREYOSRX2B9WFDVotKQThmkK7Nxb
xP/Q0JYCXbxGaE00fTxJOUYN+e73m1Fe6myBBxD9VXG8DbZodP6qvfDmnyvJVuBO
eSKNZRvQCYZYBmw2Rd/7kXCUl703akvPgQONwzAFh1DBc3gWWJ+l3uu6Grr3KqeQ
l8iBfHG0y0BikCsVwn3v7CXMv3SLB/KBlHVMPYMYNNqoMj4YgNusQ4TWRDfUXJdL
mGuXY6f1qAskeJJ7ZV+xSzWORmjULSQD4WjCbTF4DNl3LR/8sT3z7suOd6sEIhZN
NrTQCw3MhwGJ59ZjXn937PGTJcheIlDNV3ecMm9P8ig79Gyz6E6rwJJrRRUN6xCK
hvRs+AvmBUP1fWhkbG4Ue5iqTk4zahVb1ElfcCpGweMeT60eGRlJRXuSVQHZKQM5
tUn+cvFCqpvaWSqyA5TfQ42znurct9cUBVgSeR8d5GgiLn31MlKxYI4aShyF6ba7
QcMR5MAStCeBK1nrFUAided/IemN/0jXagJTXYnoHFf1bhe2JAAR6/gBGK7/lFuP
cgm8G2Jp5qO9yiFuP9V4XMSPTi+oUQa0HuUMLrEJ1VJoYaciHIXflZJXDqOcpWnG
pLSx/TFMBGSpwaamBzakRUUCQnSGdWD37wHl7rE20W/e3eFinAXj3qSr3SBVQO7P
sq6WStBoLWADivMERZ/Ff9YqR3XnJ5/71He4+QvDq4rpUlPGvnRvRkMB/8gkLmci
1gVG+rw//gTixFyYvcTXxzUsKz5SA3zMN8MF0Zna+hIJFlp4RXUr2jaN6HmyA9Iz
s8pGWaA/Dg9nJp0G8BLg1CA1ATjMaKPecHgDqjju5Fed06L1J4/hkYD+LV9VIRc3
TLJtFHC7L8F6N+Nvg0QybHchsq9n3wTNe+RvMnjcQNI3KyE9qKMBW8Us+3UfI0zw
Yi0TbUjxRPX2eBsu+1Z/16EWOlfNvGz+lJUxYP64EFc494hyyzMf1shAiugW/PdV
MGEiCm2qsbKfuUyPfwhS8iUlb0pux5OiHj42PVAXfXmDyQX2VEPlydEVIT8K1nHg
i9ssNrv8tDx5wpcvlwxAlOkj47P4p/NvCuUDnROUXXCrpK09Gc/mvMtU+IAFg+7E
5Mpn5YeAhmMud9fy1kdJx7A/RwToAX/lIOe8DI1aex2ndEfFsKek7berMDwuHn9N
6eg4rTt8MR6oMdhH0lqIEZtnmWSPQ1vmToVsvD4eoUZMib3i7UMf6QZiGj/maLwe
`protect end_protected