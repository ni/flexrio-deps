`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23616 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
pmYWbcAdKoKjCg70FScAOlDcxgpDo8xp+DafdVM2qQtReLE2HwiBiD8eRMQF1bAJ
/HMNKtJN/1RbsMoQ/CHPrSgc2NgTa+ybtT2LBcnvsj+EnCcKztqpw37ZHyA9oSRm
PWT1b6OW6JOHoOupGI1xsZ1ZqIAjBOr+KZAZddQWMUjTHmAHb9Vr6l4YR3yEr1Mo
/DgSWLfMTAT5TEe7HgriMw2cmyOOISU1qQQ0BhlhcpMBhvd8G8dIOA7KmZENt/N9
nKqFPuXPCEIm/R/Tij3KoSdcfoppbQ6XRbrloall/vdsd7cw5p+X9SVsNRyJBQUB
7Ii2E1sLyXWdYDK4vrwn433nOtoEnhqP2CBzGoCQ6sUG/6gKn70Ua7Du3t4jXsFx
72yFG6tEG6nL8t1N4TmpMb8PwzYu28JRJ/7oVQIxT9NZwZjLqQz6l6/CmsB9M2d5
e0Ygp7vwxDo9a6vT2b2lzy8/TCnvB7IiJqNyMOcGZo7FSLDFiMibcLs3u614azp4
rfu5WwIXmaUYrEYz+0TLzSxQZGvRg7FEH5WjOL4hdGTSTy3cavq1c1nW5KXf4y4i
6ZGixDvXwLJ5TDgEiWR9U6hKIsrLy8wSgc2RRG38wCN4JND8EYb0T1U6tTQ7TOPr
LTYLLHQ3fnkYfjsX4tMSCs2abaIxCfXZ9SIIZcqZk18HZDYRunZR60Yz5PBCRnAd
baJOUPZ8Q+/uauBdryKKFq69ycs8PRHMKHRYlLfZlVlTYrXOzZcnHNCdkb9u9woc
Qhp6vvdd8MjqWYab2xy6a/ICgiaz0vcF4M9eMqiq5boaMgEwVioYIDBnO1pJb56R
Xmva9cJQ7v/K1OnRklKZvHHXmD2GqTxzBMG3uiK+biRQRXPgS15MU7tvPJIljdYD
qYYMRYCOj4hR06kVVOsVEuHlNx/pK+v8I7bfdpRiuPfPxt8DBP5HWjzMpw/qAxaw
uc8tBuWa5TomhxvaXvrzhVac0dSVofqUxnblAwdEHruI8kp10ioGhLOkWvtSbCfS
oy+aXBWoTrokcsmQNRwFQ6WhIUdFw2KswQPPJE6JzxygzOqnHywX4W69+cPmh5Ck
YhtPC35oLYZ2uMSicQUS9QmKBPXXAI3QvBybY+98S7LkwHR7AzkZ/KQBonQf/knE
PZloR5GXRzZU3iSWVUHE1JRILFqqreGQWRi0a7nIfr2+4wdMaPXg10mtNvEpR+cE
sj2MFIK1hPDz/mRVUqDZgCZgAZE0pd/4jDnoDjO1gAMmTIjFUam36fPpICDxJl2P
JkJY0iky13af9sX/2aAf07ty1NdX/9/cgvEECAaK9ZGsMwvRO02b2jTD6aOP1e3k
Yfd453ZDKrUBz56w4BgBuWF798KrO43pdRPAjBVXBdJ/hiJp969k0TwKp/KkieXu
IxZWjDeqtK7AzmsWwse5iRJg4u2qqfdjr/eI6hedt1kQBsX2HAdrRAglUb9wIkmw
VbJcLAnIDsCYelGBrAahQjPfe01NrKCXctqzXkxziD3OUp9xYpOjX07odmuLhmm/
eQgyDizxFBs+zTklQUPTNl5DLsROYhnZNQXsUJHTfyxqV4VHXRwfEbst0Eg9orar
+hzaBQ3Qih3tzJqzupH6d5MNWd71niPZAUVGyKN/jxHJzMaX9oxlUsNDxCrCpX+z
rwRrB0AKOseJvI4zYDaEEn3vBbp+H4KI7C8ghw1UxZeoQMoDX4pvkuJvLQI+RrTY
xGD3wU+FPdzSlOX2ZPwh09hXnWfb4IgylNEiCcuH+Zvv3yhQZA0q6kS1cprFrWTc
+jrc9GzT3ebzHsDE7WZRpiutAZtmYrmXJNrew/CtElhXnKkpvSi47IEr+245mhU9
vtynjUhoxvN/2QFih3bJLCRCixuJmMxArLMOq68En/tdGCr9z4ZCLK1BwpptJOQ5
ek006Iz52edyJr1RLjmh9j6lQHv5HWn6RWfyN70Y/uutyJKoFtq/U9mi3bQ8xl0S
WmmlQPeQtA5aLamQYtx5V+jcHfv6jxrtCerJoRIcNkiR4ECwdR/YwGRyOpSUQJqq
n4oMKnwrhDCIJAnBP+p71H4f1y4XtTm/aXyAHPFh58XOZ//+LEyZnsPAoKdTskJF
qoojT00GMskAduJbiIFVRDQuwZWS7FHQiKL4JzBg8nV1M/w4twkWhnuhplSNayyw
L5g4siDVMZe0HL/RpTXJ2L5XPTkHGqjChGI+05j20TPcH8bYnPbKURLfI3EzD0sZ
5eYUfhBARrpGXBQ6MaDiG6JTMrm0hrYTCdJX3jssHZVjJgl3a4aJQ6jDQst8nSgu
0/pzoVhUdLZnsTCXzF/bm3Pv6eCpTGsico1MxVafUrqqYXAIgD7wGNiEXpuB1kae
6EPF4HagTSPVoiF15hZVhI6UfXPJVd6HZtVSQZUwTnBubglxmvo5uUgznykw+sHr
EtFYmyMF6O1TuuI13HG9Ot0b+emnBIlBqeoSv+ql0uubOg/4YqJRqhsO9X1md3Yx
bb7GmqVjdErVepJt1hJq8MC9VmqBJ+VSoPLA3R/Q4Xtit++NnsIJL2nxClDtgti4
oH24PpzxuNvhySGJ8f0GJsZVW3SNPHxe8fGehTmgFFby5wZVnJSJF/94SRmamkih
jNnh/mfLkEb043rveXIb2wxeWcGWA5dr9jDBKat1sMmRmZwgJdlfLafJEpveYUey
Tzua2wAA3n8m14YP1dZgx9yUKtMeWBiLeWqVwPzcWU/ujZkU53K6oR3CABjWCdFC
RjBS/InqylQFyUXMojtu54v43oFD76VpQKlZRartECCT14O1diZ14KYqyg/6cMQC
UpEkKoLOZbKACpsdH7uV2Gy8b2KCs+PUSwUdrrVB8U03D5r5BTO5z33itRNWDL08
rotV0QGxjyrYYCMOf9bmW7sqlw42p66KgqaeyRCBiT/15Q923zXDa1Ri/r3V+wts
ksbKhSwf6KPYn89RtOioxW+sRbDx3PYem4fby+m6IbXUGc2IAUvkNKo5sRxu/Q/x
mGgqJ1H7Sw1wLL5jO2EuYvHe/ytRyd3VhkXdda1/rZgnzwAQPqzFt1YiSS+JtS08
SIgc2nnMv+oZvCmOLL/ROGjxCKLtL3z9vcMSxKK8kFbzYi/YUoVufNJLi9UgmaXP
aDD3bfjfZCJlDYDXS/iqH7ou9y/6Ex06ANaGH9ADMEHrmuY/hVBR0FthaT3mfAtR
X12+PRvdkByIEerdpw8pv2XFTK7VuTOPY/4ow53WmWt4jtFRROQ6y6dXFoFFajsG
CR4kNO4+4oXNNoaZCUQI2en1lbnByfjKouGuzD6U5JQc2T3k8+XjrIAjmD42hBo8
1zeODVp1z6aamNTvcKonW/sbGJdvn2TMlJS30HP5mtNpdO3u/H4PwBp7inY9f8Oh
ZAi1L0KAZNw5w6WRci5Tv/jbvqermE9teWQeC2CQoT45uJtPJ3gtD4T8UAQEpwbT
StqPvI2A7+5PC8t/wjVpvqglYcSVDlybK+RGEfVplu3RIGYLJ/G2kEgJr8wKg/f/
sfYHt/1Jq8Egc4S1eApbITj51qFCYoaxqUpK74wWpVrbg/ZMX9P2HhA2IVeImhWL
J68pmTRCMxjUIMIcbM4divVCnhN+oFjtPaKkM2z3fWnff5Z4mOxJhACtx14Dy+uI
G1fz4xWIZBX4lFxGoDGskX+U3sg1AjXnHakLeEikfRS7sP3Tuvjxer8Q0m0gAHvJ
DOwVojQi0y5EjBwNjB5cW/8PKywF7raBcb1hjExhesunEVrJQlql7PIEhv0kWXdi
of05fjKpAwdhqqP0CicOo3+2Kp3pzFd6Jnjx+aUNQ4ZOOFON/w1gQ/UV+1rlGviY
YRXl7FTZETCbMypGTqOm/Fdw4QrEycEb4NrquWm5sXI3p03v0Zptz1otgz24S9+P
4zz65EvhPA6AGxyyDuRpBZpbjcMNo7ox4HPrLFX71WGyG5pHTooeRQtn+ECJzUix
Qb8LKklBnOHllPTcK4YBqaCcg7hJxblCHnRAen66ch/X4nusma6Md2JuuLupx6+K
rLc1HgS/dgSVrE57P/ecxHy+GUUg8UG/ydhXs4LGI8nOUlZbDPFZMXXwj5VKyTp4
up1e/YcuMZndGIYZmPrkEIWYyXc9WVYLPnLemkqrgM77+9h/Ju8k+Ww4t/Hw5CSX
0qOIplB3pLV0ahxpbthJYHpdKZvF8ehy5kqkQqJX2ezQo0YdfJgVn77aUqxYzyzZ
ZWHCZVOnzzzoFA24pjTN9RXcyyoFNfeRHBza1IBi2RWNKCQhZYSjgEAo6d8GgFMO
5ClnBLtY1836DP2rNFCU+P0QARLAFKdv6irUba9AVAMR7WIE/IVK4ObdFLxISOoy
6mDvOBm5FgWo7p546HU8u9Yq1WdsdILuYIYt3hUCIRa5AjlGMI+OSH+dm1NTCdHY
k08KZlAHHFsierbM6/suAMVcSqPRSwoh0zpqhO6evCCDLyzDig13kZU0bC1Aj7Up
9url2P+dJ09O04njHJYOcXVXyYaol3+vyuLEglqri0bOwUK7hCOYKfPGT/r2nmM1
98COKNPt9r03N2xP2+jbpb6EDzz1p4rVwZsKSbOCGk3q8VlfBkGSSbatMyt09mTW
tyaQnsIqeYOtqGsqGUpVyLxi2FiDMa071l0KJKNnb+bydf19ywP2/3fOtvk7X2aa
AdJOo+3feWlCdN2wcwpQ/Akvo8pEPknQsDlF3bXLVLzHGpRtZyPgWBPT8dsniM81
OspegYdFIOzTrr0FjZeOXTKRDMHUsa8hAIhzMPAkByOrUAmHFhOKqXW3utueYvw0
SIKbTI9+vmpNpDEm6cFY9sJ3dxAV7TIOyniAlm10K39wQcVc7ZUUZSqeR0Mqz21u
0AvbDp28Esb9Il++ol0O1RncBlPoR4OKKaffW7af4RpWJbDNKIHHj3kTOw7GW0pp
b6Xu/mPEZNWoiykxx00IAtG6rVQmORxIX8vuKqVoXqDfKkPMiqJjvGekd1X/GWWT
LxihwDy0n1FY7usdTCz+qPzXVrLJ17IzkmTNp/wSCinM3aOH7wJmg4dXjPABcgQw
ld3ZT9V+/jdoy5p3ra779Fwtuf6xIQOh5RGoCZs9uTI77QnBOLZjVKt/ffKTj+JT
h0LZvDrkiuPOmOLbm/vFp9Fhg2xxij3Tn5mgY+4NV8MeaBzMKDSvtL566JM5pn7d
6bkOG8YSdKc/nXRGMmM9HgLztoj4vKTAfKCvBRwksATZaUhOBLcapfr1iU3if+mX
iRdZdVLI6a+yHv9OzprXlTtgLurvTffhOIxk7Zdq9tX9SAF+WYB/9u14g5CVEnot
QfRRMlD8FawMk9mbBzXuUOkbe6LOT7q7QreY/SGBKzNfNt7R50n63TkUVZISHFId
e9NrBzvHIHWtaiIzuQmTVjGUkQ9+CEgZlAtDK65iTiqvmYzEoyKGJnxmUK29KxSw
tLK7cPh9xnEWcxEu/Xa4neAD/Be72mWQcSuUC1BFMrP6ksiFMk1muCmGr/S+RibM
mHa452Ui5tpKMUsmIZVmb4RF7l4P9N+jmqTuw655XzBUrEw+b0AdgMhdCeJUbfR8
+E/5XUPx0Q9N2D8p2x3GzCBDlomPE0saupr/ScJlG4Q5yPH9AygFHJeJ7uvyN++4
5ivlzVeREGoF4qLU++esNXldzWvld1Ei5ME7jdS2H/IkgaejTE1ZPdwWvIca0Lj2
LgxzRqmYTI8wAL0gSJk2Sr35E/8ogbvkZPaFclShBLlL3aMw0F2fdCQd/OvMYP1D
/nqZvWhEyHeShy5gh1nwon1rpCTIX1MsZaQ4/JAWUC9qSfBGzVuPN+hSnx++ZqCo
5wdRKv2+jVAE0txaa4JQKmzaQRyKOc4BYxe6amHPJrPiUNmATi4KkbaUEc1rI4/B
T0NR0SQBKsVIA/eEp5+IsdCUfVKmCeYC33no8qVMsrlDGIDPvqh7AdnNXDt57AEz
r+MQTiBcVnRaE3EEZMZFCpxE3C0fBZE8MjdkoIWO7GbTs0QpRUj9CsU8p48v//0s
VuapuNHGFT1KYBIepOT+KmkmVi/Ru1nYv4u6jbuQZegnO8DE6UnjGEnt9NdY06ZV
nQdJgKsJ5UAsK4ZQOZsOVRGk7QQI1vWmiOgikjuuPusFEaAz1d1dUad02xJvodgk
04To4zQ3zB9SmcKWiYW3hpHuDsj80QEvIlNPMfgpzbn7qJwPjnmGXDrFiBljaCA4
omdPRLHzFqxkj1u93LGrYn2noV+G2j54dl0aA5fZU9G4tnclpNhEZxWRGyqwPi7P
dmd9uCa2Hobupnmnnz+/iNnxXPUgNXeH+tixqUBsi4/+Zwqhx/0TKU4oSVVQlyZ9
y9ZK4oQvH0WeZkiZcHfksiP6KEi1gVAYNfty0xyG6AVMu/YCa7WpSvIdch0LPg9a
+tcPd8tL/0OIu+S6sXQSQ0I3moNjDSedusJxvYihtYVk2yP4RwZ2bJ7lVMGMsjZQ
RX7OAArvRqIpZJrWehM8v7Fj/kTbOjT68SHw10YlhYMvfkm10cW22hsxQjsICKlJ
9VObSpamaIz5oenkHicbruAaCpaIzAPEjOiD5lhuzY+zr4bfS9MBX0Ul6NbBbs7c
HnPEcvbUtQiYnQufmCk10FlIahC9S1FjpuCB1t29yHxYIny7OWyk2JL6RQkEupLE
LZKjPCjAr5Cmhb4iX3DXVb033v3Jn7Z6VCKi4wZEquROT7ltu0YbAuHC5M0HuAzL
OVMFGj46nzVzAkM61FsnI9a7wDY/xeQ+8btcZ25f2Vm1TA8N9YjJEE5AbnWNBfos
oW33IYjk2i2G0vQMUADI6uoEfq1XAzd6vIyTXi4AO8mk+3h5VknrPvZjtA8R61CD
KT8euavutoaDP6VnKD76+j5Dbr0S4HgN6yokKG3fNLt1yDhEKANs77igmEjAZfOD
K8jKBaT5qCxnAy9ykHCGmiMzKhSacvyM77EqBYJHlcimxKsQGQ6gGI14Xpc0Y3G6
8w2RivCZJkhVTcKFWXkFEABBt08W5dowX+tACjX2i85AipW8ZxhOKjLJTkzZjPDc
euBMp2DDzGXPcgf3XRzXpg7ac9s85YQ55XcmzsL6vwNEPDq0TqezVerGv4n7haBe
K77QxXAfgcq/5DmqWvRnrEA0o4VP0n2V3iN6qWd9OmjbCcjMUX18anZW3dBUwUfi
1SsuiMK7UAqZdFRBsJv5IX6vZlDykH790pN9VDlD8iZ6gPSsN15BQ7STHPJxNhKN
DsqW1pW094aIrwApIfR1glz+vWbTsejKxzW48KFzaYP4CmWpJ2xg6djqLHXkfxUj
nWv6sEpou8E8T/xh5gVmwvuPVJFvNtKqfpJwOWCthPAkNR4ouY6qUYmwzmBrYcmQ
BxSbKHHAXm30E/E4oL+MIbtiYjhb8MeXAii/NLZ7cnsqKx5Mn9XiKRZyy95BLwFZ
iE3oIMcdtGQzvRcd09orhe6OmOmdSGCAfsjo7iu7jpnisbegKclBy1MrADSgF6sK
IGJTOGt1L9VNvfTNQuO7NwsyZ6S64TD8ttaiyM7x1sQoyNE9YXR5pe2i1ArFh+zq
3mq8bqnAkWvWCbVRZaPnSoYM5ztt5NXdOR50n7PDrOtaknyq8O/Siidz9MCAO3hu
PkmZOpz5C2+RGHh6TrzcgROvgEKBZjvozxKJUEoGZgUq1NIXAPiCbeOM5l4TG52u
sQAEE/b4F9myveCLiKDVFKOwG+xLK3MjIpFfFhsWgktjxH+d8qiGstaRknWPAPFl
xnHaVtXm4K3izrjhdm/K5367B/AIqyy+59ZLS/k+9jgfs2s314zawTRcRWg3KCU6
+6QYVCNfhEK9W/DTgMSvve/G07h9+cjeqTIyDicO2lrcG+xpJRuDvv2rR4U5ePCH
cDoE2j1FUsc+oSlZ6KlN+Pj09HyheGi/KGWc29PbbHagwVoXIXHDSV3s9YJyt1Oy
Iedf1geNgKTmE84idYkWZfs3hT3TeAoMNbFI0egYhS5IfFkDftkS76Do7xcGTfwE
UFHMjeFqmZUouACJTbT/BTq6s/PhE/wjTyG85AKU09FkO1T9KhOQ602Ivkq1v842
TPbjboy4RMPKol9F7YAEMh3oflIj7GeXxlN1bJ+WpJdQPMmNhSOrnXsaQRD9gQFg
Y4NmxNI9SYJoZIAXVdzu2AcFQyQ5HMC4QmOGnaTJAykI3DKcZtCHjqnBXU1Kgq4i
O6VsQ/OjBrQEqYgCrr033VOV1k5Dqdnsn5vI4UXySmEKTs6iOGO+hsqwmAQ1O0Nt
Q9MWqx5cKeDzViIqbz4+zQUgDrcz94jqmDTWCiyMxLAL/zjiXkH7eOSmGs72LiGZ
/Gm4HBVdrtALaDnUW1VSkvFltdylyz3ftuO2EtzalP/dgzgjnFxMppbv8IQYB1TY
rwKSvfRa7RRW29JVAiRMv2vXY2qWkU/PqKYRQCXVA7+Rc5XqKmP1Wm5j3EZuiCEu
6X3KvCqZNy/G9FIB4LQwJ3JERFmoQJ5KrKLH/xKWoup3AC0r6ztDaPa/sC7i0eb0
EseeFnHZneaOTW7JbBvz03MIpZ1QvUNoIAi+7U6jlbyQ5pxxYWhpJEvPelbY3peU
niwZArXXj4c9o/32t6X0aYgJc9ibTA3B2bcWwQ6Qle9Uz+R0hH4JPBmUTc/lmjnP
Ix8hi6Myu/Fco+gL/oLOQQE2nMWZKZ6zbPUnPVKImBG6CPE3ICoZq7iJIYk6squb
l7t/wc0Sn4OLur5lMJbN2Tr36Ly1neXl0d/xqqfmaA7qrtqSYefP8no+6MPWeAJB
/mVMlMrvfcN2pnKkCXCfAA3IF3BJxfw6fMrwI2MBcB7Wu73cvbE4A7DYUCDbVZwn
wTM1QsFvEa5nFzk1j476taWXY6CQqk45+2OzlwIzaReZt3GWFmiWwmFvFwEDo7NO
KsyYkKSYsMc9un7qznAGx5gt5lmDzInBtUUuOt0evJw9FnGRvFntXlrgIoc725Eh
QeYAUnbYCBg+k/hX6aYl4ry0epYgtUls+n5BgPivzaNXb/Ou/tHYp8svsI74z5H3
6TzUwct8kSG5+1eW2f2A0FdpbrzOfjXiOLV54LqynAuRNzSz+8aPLsN5jc+wgWjp
mcf2xuywqUy3c2X8ypEiR8h2oTko1Xw+1tg4BAY+ztu2KXazO9I6pqtxBzlNDGqW
njPZFa+MfDQH75ekzrWUl+hEzH0kZrpybEbak1MK+91rl39XB6fjf1AxEzlmXNpp
z+L6HX0jVOK4bN/5NvpSCEp2sgQCu42orJWmMkTSJyHB+7VtPCjCx3pv5FhBWQc7
+Me11CeX5KAlf45oxbqcwbpg0tZUSg4qOizmPtswiQU5UezS+7RB0Ojk4TUtSRiY
AD4zwfBcrcnxC4Uy1nlfp/XpustWPx8Phxv3Dye8/km88UZXUBfEMqvr0IQ4m+xp
+GGCJAJmnzrfaD4wqpB66kCeplbjLVwwYv8z1AOFK2ZZXNI9OoBZyLjYd2HNZmUA
xE8RbnPbg3LElqnLQ8T6QLZfEjvxnOiXKTdQ2Luj4JpyY0ZFhlI4+Y9r5eaavVYC
B5seEVK16CwGaF3WH+uMjZxsdcuf32VpI6OfhlD5zgpZy833TC84Woi4aImwICUJ
ijTYGHtTbCymm/6dI0oqBJ1xyMXebbNV74llEQvr3PmtFeYZpK9VDirZ/yMDbJOP
BuDaInW/QpJ5al7zlprTQR0EhOlUZkISkLsw2KBEMzrqDW4X723t2rKN/jPk1BtM
2v7sguGODsI3eerovFrvvn3QUwIAuC6ygs+zygWAxeOclVle6yt6nIoDmUaoSAIc
7COa76qKStgxTsPaSAYTnNY/pOd/EaQTatUl/D43WZ34Mh/DBVjUTR+BWeHxcXNp
NcihOJuKwBHijNhaOhPRwU3G59xeISuPtZmHNwB3WvK7CzbsPo+0F6KiUJIEvxHi
coK4VlAyDa5NzfFDIejskOq1dijlO4nQ2FfvfCdUxsrb8ehfgRCVu98jlOvMPrz2
FrmIQ6279b00kMdr9WSM6N7CxiRVs7QDaDcknLu0MPrZJRJZsjllEFAhU1IpnqWr
ZXsLlXMkj/kJY7bO6JF70+nmvxambRAW2D4chY0xsp8wyCDs+fZ0SehKYg7NQvZD
De7hjD3JLDq+3UTWsBE0WYH5SwvHi9knjqwTkLvEbsZFhvl1n4VOTdIvSaPzyhQL
vL1V/xRKdhytVZxTKdWyNF9DrBnSoOQzki4jChGn6Cbnr5gITE5A8BzpyBHqOLZS
wlJCpl8KWI2yGuzM5bgcii2cyEK1ooHfh7X3yzpHcfsRDQhd6vJhVpwmTfg+X+3K
Vi7Qq4UD8FvoKq07zAzQeAHbfhEJmnaNV6Hro2xNjjU6L4TgFz1PWQ+6V1KjmKin
lGSUgVYu8T2lF9rLpTBSxv1euFuwkH0ynwQSa2HhHOWzghUlkiYtVWO50CRy1sac
cUnnvS3eXypkIbDUduTVA3pDbW6AcAleXUchx5mSzXX9oRSd2MGMhtZPvfy/KTry
fAqXKKTMLpduwIo3hM+kl+Agsn4xmJVqYOw8qsk9rZrre479YLarWLenCvQmxk+9
ZSIEB/IDsdZSUz5S7e+IDhPhB3ITVPndvYEHmEH5nkc6q3VE5YSOj6JBVC5l0aFN
f8uIhxggm1HtE6ehqpCDpMD/sMZfeZrDyid8ytjGkbvPPD/rv+4VqQMMU4XEPqGE
S82/9LRjPkq1jc2Su6DR/UA+E9eQ1W+TPMVB8XE4mhOruX9sUEvmLCtMi3rd1DvB
1ca18Dqs98bzGH9TUP9TOmsEb0zswObGNX9fACaJOyNh/6Af2us9NAJ3CoESH4Ka
CRW29meraLHTuMkQFI5ad4VBDMofz0OJrIqmaWhKET9X2HUEi2OQdePmjVAvutFl
pmZma1zqp+OTG4FKg37sC7F64ZyirRgqVTp3+YfBrJZehiXuy1IL35DNj3EVqM2q
cxnAN4oGORMdRW9w8C1DFOKV/UPkA4P0kM61Ucvv46zK6z1BUV9GoWkW4dMTL2Q0
9oZwxSsc4QdonNW3TBWIg2JoUBNQ+iXBo1wECs+bA0YU72wp2N1nl4PuisgLpPLa
2Dbxn1xz2vINa3Qibi6GrLtEH6mrwz69PZQGhXGsRw+YjIlwVJjn2sVfiBydFehN
ehl/jafXjSf7zyE9ReHbvTZmwSL0Kq2zxmDgqPXX+mX+d43nBANgB/C0Yp0S/H23
D3jcC3jpQadebEBqXDUFY6ySgt0LG2Uum7bvks7uJAQAcJ/s/HzEKIzkshbyiTRB
oZfl0en2pKDG0Y/uBKX/QtM3OW2KupH9Fiw3YKZuVKVpuHk+YxILXJCzUejnrOpH
w+PFRmHFKf81LylnLWSb/Q+7PP5ko/erCmbg9BcKXdHoijBiuxcL59LMogsFb2wb
gd/XDVFn8XzqAzrzCTMLVczXg99n4Trk/UqSwO/xLt8Q2F1xa2bQFPxv+7cFe9tC
8UZJvSFACL0EHIV3oMgLmxI7CKA2+xsWqIcH+qiHuz3siXgrK9jEGAXEpcT5F+cr
1twEIZH8kRjhcl7tN/CCX9PWY1gaAJ12M1Up1oOMXYkO5DtZb3Vave35TDGEY9vR
ncVFD7pemGGCQX1wCTEf1WegMAqd5OLg5avN3rp3DnpPUba7txFg4vc4aC4YZ+GK
4ljxeZe0H4s3BK9+H2EgaAYkz9CAQddxV1KN+YeI9z9p8ulcAOsbjNLySCoWyilb
sw+XV/WeCDSlkL5EZ1JNLq/C3Og+S/Lpzrma9s7eLN7CiCZynT4DpYBeswgjkgth
mgYzyubk1dYieoxtQ50JZZF+asvOxCyfSlP7OgXGr9JIKjgzJCgrwZBguPA1BUUM
3AMQqPajYUZMb3gTCnHuwqhO5+EYz1cjMYnpgFU16sD6bmNf0OBkwZhFFJRRiGXt
Ywl5l/1IfyUmoT+3HV1IPWZ6nI3viHwMFKc5zbF5iTLisowHk7Biw6Jfvl1KKkEN
mKeKDretGiXOUljf0PqywPQlp+WGGva6BrZOupgrZHOLyhVWl49LQzfLz4/6i3x6
x1Tqhn6rew6EIZIinF8X59McfFEPta53caKrPDllnC8+UPYZlUC5k5yQlBvbW9iX
avRtmvMKHFAU+rZJfrN8awuRiRhGz3xbxcy/7vjeTN80o20KFeEC6SJ+J+niLfOA
YExfruVJnfv2r8QQMf4iIxWRR0TwKWQgDlbyva+/kMQWIIf8BtWWCfcy0jXEHvtP
6eSmv/BLBX8a9EdX0xVGT7nP8tnLL5zddSCcU1TNil6vI0GziAjfh2XUZgrTkVms
pfOAXxlLnHVAF5O8jXPWb1VWfiWK5kFDyDR1jHZazHJLCPHE70CYWbygVk3fZSit
fcD4s8Buu/cEfui2k+YC7g/GZevzikgtnwleSfC0kOsdikrohLFwJ9GbQvCDfA/u
PjTdZheWk1nC6OKoiinNSw6uQPiZHqZf3W1WUZuxWpeKaw2MJGaJ/+zszTJijs+c
RdbVFokpR+t5+T3AHwtp1yESCBkuMc/OzWiW9AvJ61V2HVXfkaFyLuqSSidLbd14
fH4bv71pyuMFAQGvuO4B/IPksJAA7LXYFGy/7NsJAMmEh842ZFvXFQyjkPVp2zc3
+2JmSAUeRAMLP+kzj4SHSoVlXyVD7gLTbhQYDDK/T0YU8nJ+1tbdCtVaS+zhe5fK
F1cK4YJyr2xhAUeARxcOHpQ8kV2Zz5ZOp59SOZ2lQ3ykVqYa8MZ1fkeiHjQIzSsP
sLoE2soY5N4FGWpV5KoZHnGjjOXUZrLOUpIonr7etyDyJ6gsduDRreP/PjWAF+lV
lNT0RXHkGgC6KceR+I88YP2FPxA+rEmD0OEh3RYPy1D5DCpv8gBrh0xc8ievDkrY
Ss5LiwlpbaljMgI3dVFf3noTxlczCryy+390cD1CW5sdWE43Jv73jFlY3hSMfjYZ
pBQLxysjQQSFhxNrAJt6fE4GtxkJe5dvxddO+vHWQFYvc26V7o6zQXPK3PLv/Z0r
rkpbej2/Z2QWMn54mwzMDbbMJIh2z0PK3Cabvhw6gsFZcdsJAJN1ZzGKwULzXSi2
yWzcszHGbfCulWYPcVrKDkupvURID3wPEU1kezioOTQR0IdlQaYJ9R7i/G+TMGVj
OnEG17vOain8Sx+mZazyWvq4yzE5y3XZCHDXW+MnJOpf3bFIRKqazh3D+6RS+r7t
KO21mLky3RCbKSqrrepHpbStSm/QjMqbAOONwEc8ftYDUgOm+UofFZuWrVkBdqyz
hS7uojAqkfYw4/k5Jwxa4TN9fQAj88HcybTrZtX7TkDP9s5oOgW7vYcUQs5FyFfa
Ml39xUy8dQu96FaaArJ1mOmPUPXntT9ogCKPEKNMyrXRoh6ZHVYAGBy6cz8gxUnQ
XgvajiyOlSJHZPmyMhAVR8EZNahMWPO3+HhUYGD9bD04Ydr/s6CCrOazZk1BH1Fs
Qd81qLGxuKOlfSVt/MmDiVYNHpD/ubEmderUbbiRJmtrUSpqO15si3O/XvxR7CIQ
SA3vKGUwdRj6Ii+evJ+MgYMbM1XZdFRv2sJCfhdk6SFh+v6gZWNiG3e7Nr1oTZKi
oBAtXBlnMV6V/VMC7JnCRWCEPiQTJ5T2pYrEpRRMT5aKri23Xehll+qzCMPnoYCS
JnKceLRsCLSnT6VcYv+eu/QTfKnxX/DaVGdRMOPKaH5HdVkTE9irnMWe0rBNSUB0
UOGQx4VTRjCS8ERK7HhZhxqftk2t4VA6fcFndfVmg95/BAHd5t4lreo47dspDmMv
7Lx9cY1LeIYAbfuIvkMMlomq2o7Zv0tinR0GKo2127rcczbPQkpWWgmoTD1xsSRD
c3X5zThhoqwJ7DvqkrW/rKPWweqXEMirQzYEL9Bg8IFop3fBs38EMDRX/k2eXZbd
QWZQ7h72eRxZsvNOpfRcl2SHCF0O5D0ID091w6dxFmBJOpY1xFRbWiNAyoJhYTXk
/VpauhnMMBaTQtczdot/f2InZXiYlnPAFgsVm3+XrMG/1HR7GQHT4Of3uYJmMUKI
hUN7cSkr1RdhsPLnoEkLmTGsehAUlLh+x1kP/JTZlQxY8OAhFbUQkJub/tLt/KcD
eX79dxC+knBivXWlePzqEddzSGPCKreMlkOvC2OFvHPHm3qg7w0VYo6ytoQT3e2s
zLyB+1CjBDMkmIxODdJGPc7CaImm6xTFUvAv4XWwGPgYOiQmjRr/W1yoDUs/myY8
7pIDv/fGyqVEE92P/nrbOEepEJP5Ft3vmH1bfiVKKD0shBshkBy4RMe/geQkEyFv
gQ+X64+SunpVrQGfuflRuRu81+sZUju3XTCKuAswJdDZcmC2SoxLKLE7b758iwL3
mtf3Jtz7yA0oqp4JqyFgt5k2Ot7NKhUg6QrzZF9ZQJfB+KDIjRNNtdxPs2smA6j3
bK1GF5ZVZPrngP95TUi7dzKkeCpcE3ZFJUIjed6iJuTIITpkbQFpJzrLHqhE35Np
kLxSzJwz5Uu9YWuDodYv8tf2t4MGLtjb7098UEpXyuLpaYGVVDeC8oPmyST1YKzD
u2MAR24K/BxApkSBBcmYxt/jLcwkCXkpz+NPSGhHlvPAeOk/20Q0dLAeId6CnaTY
XsXIP2v0N6Z1u0+bNfaM8Q9I6mZAKzsCqR/oac5xdUZUfuXWt5F+NgLf+nnezmUv
b9pxYeVYQb7Ta9zQHUylIdEg5pL8vQlvDdGGRH+e9u6BGTHg+JeOMc6yXUJZILKq
9pb0rrcO6lulD8l2zQIKZacNoGKkSh/sJ+EPAzLI/rmnr5uDl2ByiGrUvBSwcGmD
dDb9rQsK3+0y/tqnxg3J/pu6C/ybdIvrhgAz6uiwCP1iChyOU2gwio5xu87c0ErO
0MRLyff/O0jMxidswyXd7tPbjUHu+fqk56k2rzSgcQGkpG/pltD/KC9/lwhCJ3T2
efLY4zsjLoQzQzNGIf/wLLRt1cbOtshExBcg4MUuUEVqNZqQ/wNaqB54Qu24qZyj
eZGMmtioqE2mQX7t1b3QINy0pF+YhiewkJQfi9n+kUacwThTCu+x9XTTsszglBaq
2y0V0O5uvzRzvKQjjDCjkpBUD85MEIt+cz/JokolkVLW6POElyyoSWZnDpe89VQV
ksgUh87Ip/Uft9EiVQ28xr8gHl/DTHcHAfy99RODTmbo5jk6TejAkVg9NHe0jCqx
mWHfizIuRMHhWEZv6utK33xttyq2OTwdNiuIWZh8j1JUYsnzPRvrJPtOetkZEY2w
69gWij7WITH0328cGcuEfmf0AdMMY5SmiO0Jj6deVfcY7gLXhSV9O6tsj5VwwkGk
pFdj7wTYxxjLRT+z8Vkyea6EMKLS3Pwnc9gfrJjQ/IwoFVMAUOh5SxgynT6e2czs
DFrjZvLbDJwFfiuUiAbY+S3X5wurCJr0++18V2h7xK8lxgaXfg1nRrkILfG9ucIg
89Ay7FqxBqX2i2wPja68auFNIWPLBDGa9lwRK0pJwByQOILAvgzbUV+wIKrYu9PO
MpVPfTh+OAAI3ow1P5ZRLGM7W/+NMUwfx3gAHRjTSMUwhBGi7afHy0iI8Lwc5Do3
l+M7z3TxKhzMgEfQN+koDKH65/WKZizqIECzq5YrQ12BkcjkXGZDNtUhKnD2vicD
kwjMH2C6+uFKyRuhgnsmDlgpeRB4G9Q9HgsqUI18wYro+WigRzhjVy6UzZBH794r
OrZbcrD8qUEScuNfHCZi6mKQ0akyVQnUWo9/BzofHt/gmaJ5ywIrfD46o/aqkQta
ahF0yV4TrxOCjd2mDDmAUtQDal1lxPO7U4T2FXH1TBlmEuBG+C8fHrQHLkJdg2Sp
U3VMP0tFRnVJ8xhbFWr+FGPS3udQL8w9KTrSvukda4EmW+oBN+6c3TfbDrYtuMFe
8VIHeWSa9M5ypwLz3f7KazXfGnYyV+PEH9MZz+yGnDgc2+cgV4Nruv4JtSOjQlgi
3e1t2WcOOXnjqI5ZOes+cWWEARVMlu2Vqjl/TmELAVoXbiTw2El48UBLF77yFhvU
Uc86G+1uNkoolvxdEkaEFPLCZfKYeTGCOXLVV58BfG3H5xnKGGexxc5EIb0jZOqN
1SVi8nsKBh68Rvo7aXj7WfkuO0FkKhexEkwB66vFOteYTUzsJH6BAF21Fr3OeTxE
ZRQx9nFm0wQH7LjOWlOObzp9xzlKyyo+7jynvDhOVjCZHlq0OPPJTmsAOAGSDwsp
ENkG4/JwoJ3RWiqgmo1bClRP7Ytc+9+u144+Pn7QriGLxc+vDoIGWB/CXYdnuged
g1aa3leT3XQxkPUtcFjk3SP7pLOVVnldZFK3m7itiGTs7Ov7/O7GLhtrOoLNlBCm
kezi4MplJgm1to5fbJL+TVsDVtamY+J0VoNB65KC9cqCxBx8jMKPZLEZ8k5kZMuS
FTMSqPjRcHInvSlHEN9+iH0smNZAqUK6Gg9MNdD7aMAwrMcU+DQiiiyQZ7iRDLK7
De/Fh+q3lQBjgzm2j9dPbWS8xNBfeojZeE2fd6MhIKeQkwXU2lKvzkaOewF9Gh6P
JJFiHas0O29Hws1z1nj3wA2u5f0zkKqr7BEKlPgxoNxslO5yeLpAKvShb+5eOAWj
zg08+c2J5LyfiB42LY2Wuh+Ropml5Dg2e6QW7KH5V+DO0JZvVogcZOa1WVr3Kq0y
FsAb6AXJW9yhE+OlMtNZ8G8US0Gc1IdcFnAWPkX8ay4Hj6WS1aBnsJ2HXHpweqQn
zdad+ZSA9AxZgUDTM3ROXU2yZCOZy3x1bk7F4ygvQR7SfToSfBfTet7rGYmFRSZL
04tm5YfR2OJwjAcfuZK5frbJFXta0LV/ZZcMv7U5FI5y00VDCy3CysLsdnuxoEIg
i8BGMJRHqd3dS3E4ree2U92SaAqzDhverTr4KIaPkcQwpxXQIPxGXQ4RPezA/m/R
M7Eg1j+j5bMZF6NOcOpbEEEocHmN9OUXpcfoY/YJMDquJZAlnvxaYnOH/GNgZIIJ
3oXAmEKqRA38kjiiCFs7twRYZr/raX0MB7xZ7hVDYKcx9/sG1mt6T2CLsUpnE/vI
8vMKOEiTKTkAmCVfxr465LJQObLdLZrvlP3OumoeyoocaOSntYDZpIwsALGeXEGk
jfoJOwBxe6MO/+i0Rov9FPPLxXXHbwVp+C8tRyrHTTvNxxnfCt+faH7UHs0kiUgx
coJy77UkYaHqnZY087gkQgW+3pVl6gwI+mxWcEoJ9aA+jOXwQ270YdjIL57RH7XX
WcY5rs32Te+LWLP/6YV5agXVcWk/JbEIoZKl0jGLg5mUFoZBBv/IN/yOugL6JDSi
eZnFhEJdscpFfDhwKSKjQ6RAh2pecBpOgTiOQLgYXO1nu+g0wYUMIBgqX2fgDgSr
r2JzupsbxWmBM2augYlB++urtSxqQu1Q0HuKLh6Yf3lL1FT1aplYoNdBehn8g8y7
1aJOIN7ApufZ3l77MuM/1jIXKrlFAsmfqn2j8+3fMy+DAyb51YunRaCZeIqTJdh/
5K1MxNSrQldUrXXLZEhwc3RX8BZUXhAIfZd4e1jia2mm1JEpAnsAqxsY64wc7rch
VbcSYvklsSz7zXqCiAXh53cqgop3xRTjrCo8xT1Qq/O2zToxlGbCEZmWoGIpzqlW
DFOEB00pvrRF/SFGZf5gyL0jsxVtU9ahMeHGgOY9j2UeoayExLnx/SqBfBKaEYnT
aB45PYvT1rTkuFeZVsUguGHvcSyrUIRkl2Jay33ojT2C9mFZvL4sq1sThljHW6nl
eS5CY7Cqdt2t5QpDBK6ZqO4yXjvFn237y/rHl9WG16eYuGNLfpuYfRHmNd+CzVI8
UrlsGrzoNgFZB6kOHFX0OLwg6fVZvCDn/Znu0GhKDDssldoD66FCa35PfhAxc5TU
j9/RuAcU/easKbBQTIYbedVyF5qGB0MhaGiGXjs4gsbr4f70IBgxH7gfoHxJ/G+M
1GOrULzs1qomDyJP1t7XgIfHaWoZQoAXJ5fM8yS6mAKGpsI81D70Ubqisv1YOOau
yvT6wdNPv6MuOH4BaOxKDQRTm85L0Vy+XkDGZJFTRjDLwxiGBJvVKXhGCi/6NGa4
KS0+G0AT05z41qnMe/X7ZY20uglpLs++XRcPBZ8dCJLz96OAOSuT4Q5UdlT93dZF
6NPzzeLFx2mCTQfKsNGkY1eBWFiDMhYoJy/RgFGz3vHp0nQLVq/vUVSEcTqiZdP3
8XzZqwsXfQkHNkn21m8mf02S2YGfDy2i50WVKodwgSzOngT3J1c+k1olJgDcfqqB
tndNjZJ8bSP2RHkF2rREKwGXanXqRBZ0H2iZx0JSkY4Kr71Okc0xzUKOmV/L2Khc
iHFtGntKt1vKgnPIc9No/m9TJz3UrLJUAEqJlvjmOPEGSquoCBXXeDtR6F1GK3o/
Jzbas+XlIyEHRmOIDwO8ozcKvL1uksWRCMefSOq0rWE4irmfCmPjXhIweAFNnUKT
07GQ1zR0xvc5oRMICwGgF15KyLuVNS30FRY9UWkWzf328V0iUKz6s5LKNKBhH6iH
kw1nLS2TEuVUTAlbiMSSz2PIT+RcBt2/ie7/6k6LWTjbANdBvpJzDQ0JZ4sl5MmS
Djx41q8vEyXi+Hh4aE505fkH+jpjox2N9Esiycxkw/EgNT88acvykVjWqTjnpgfO
xd/hzX0YAHJwpuEGY4BaOIDrMsx4OjhD5A57N9LmUe/doBiFc8UB8rhf/TC6Zuq/
3UN7p0tr0yMz5CNJ4Z+t0z3jrM7Bn55CybXF74y1tcBTTKAiJ5bTYQGFEN3DnIPm
iY9k1jzED/+U9BHhSIAtG+HFnP705He2xkjpXWm2TlZO00Yl9ToMDBtfrJQxsamB
6jt+TUVYemX+DIzBUezALUZFqi5uVtne66FGlmuNl9uW5brXJgxluOsDWpN/p1Xd
IfsAMP/LaSYPc4bbLoQxdxY4yUVerbeknrI34pIncf1YziHPwmVJ9bKWob+OGceY
99ux68BsucsAQromgtHpprb8ZctGYbIcEId0BEQF4evWVmsX0cNO/D8kDT7wIITf
by8oq3BnT1CDZOGzSlauOUmrXh/FmhcjipARU9Yxh9EyKh1pKxaoIuK1fG/3Ve2I
QTu5phKxMrMNWXEdXjJHfNA2QXXbLotNulZwvDedWt/ElzOoP+GgQ/4NefZtXxK7
tY+eQJCs/vLEGqqp8w7t1wZwXBKe7znIAcJl0ROiYdO11vzj0/ww8+UxC32du2uy
VDmkyNU0nCrnAVBmDC/o2cF2mP2odAr2WlgHGFC/dGT9i89PHf75qXOfGwWgZk3O
357IdNBP7tvxzt+EE6jzAMf+7DrVX/E6cY1bzom4ysv1ITBMIsZhbeffDnXvb5XQ
rY1MGbRQVPFbipOJmE6g4cq01DdOqq8olNxAPT5k//IbE4F+/KrRRtjesIyO8whs
vcphWWxS3D5HFPu4IjixbOcH/zpJNco//xA2uhJn9PYkp+EILD37qjiaj/93pd7w
xQchzpx8SOGO6usDWf0peU51Kd9loFN98PDFCAWygPvy0eL4FXwtmgSRck5guiUM
7wAxsiRgoJCZrFIzQgxRSREGW3U9oFDJpAO6o6kGAmi45h3WPkRNqqzDs9qghYuq
NrPwYPDHTZ2xjTwCijw+mg1GZTv7zDgYkxlvojTAierTbduur3+z+uubznbNSeOf
djc5EULbh0Q8zJ74XEDY29bzxl4JwzOy+lwiHrrIlk8CaFzc7M8p6ORcy5QfTG2z
jnI5OXmXmQeDIVecbWSRWUBoKMJYKgz13hRivwYgvbJFPMzUwgpXg/LfHo8jEaAq
YCAYkDsGs45x5LfFDquvlG1s+c+mKg/8TGSp1MHGBkzwKG3umldwcbbZ3wfjmReP
3d1gFQ4Y6xt9LsUWzpwyzQD1rEH0huONhqpty40+FsVzsMOQzIbSDmjaM4bly50K
MszpQqLxxrY3m7Galm9VU++Wr5RwcUlSepufOdTdV+KHE7Ohm570wePynsgTJ6gs
lhGML1pdB4wB4y4nS1yOvG+xDPl3wFxdcMbW3GKOc7LtxydbWqr/NllGi/sMkUyO
HeKFmALRJfYicX6KwlfqirSBMchMA2U6n534Hd2lnyjT6HVWRtvdDawC8xl1FCjb
OEw+QSsTgSS0YyjYKKjig8S7xPXr0gXrmMynguWQhyyKbfEgOAw5nF5PyVOiib4E
V8ePUVl8MzfyZssCiZs4IUDVTAr0zXGQQxAQ+GNIH2DDfVNkohYe8l3TvQM+qigX
bZE8FgXaZ+8WLJUduUSwo0wj4ypOtwZGW2Vv0faD7q16Zc3HjLmZeZPxHSs8Vh5+
QjY1xIYV2gvDqcrrGX3hX5y3qbsIsOvdsOiSzrkLhh4Xc619C2044uZRrfOcZEp7
dzn/wsn3ykTsR5BX4UFvXMBAUxLnOlfkFzkPjOSegjQAChMy395KlN82HUZhN9tg
hTsaSRoDTAFY8CvZWrxE0nwHNNIyk9Qax3tJkyDZLL4uYgReXQ+l5cxw/3I0REtU
5A8NbmaVBpNph7MeIYM4LjsP7o8BjIITV9I3PJpcotAUfxcabJkIu3Ue1wwA4oGz
ZpBkRrk+bpA0GDQe3dPVY4mEOrS9jsjfZOkYo7NrPSxTCcipGrFzx1ExzQOZvNqa
dSfEXq2I+5Dtb0DSDaF1il6u0+2O4ZWP07laZtFZuzsklevyD4fW3D3VnzEU6ja8
wXHj/cepJYuJindhCFo+CQ4pY0NP7HL8E9EDJngAHaxn3uVwFK/eoVr1zWSD9GEg
fuQJqqhWlFijAWDaDAbOQtxdEurLP7zyXvY5BN9xsM+ZTzioH3cbxcMlst2E3vTn
pQZnVbSDMR/t1GuxUIpmxaZsDMg33WEpSYoMvjAgh6VhzyZEJ5FDjDcJO33fD2uA
srMPs4BAueqkeO3sdAbp/A8E6tiFTQEQdpJ0ygDQ3pNT9rQQ7fCkqCNytEqZpQOv
EcMRNPkSE4NgQABwPH/h4Jsn3XW8XZ+UZoMY3/uR7wvtS/tYN1oxUZq6I+aJprGf
BimlXQ1A2b1dI0j3UYJZjg+ZlELtUGwAABPNA0/Ettj6h7ZxiVE2WLi+MMJBOkLW
Lrs1Zw4zycIZUJFSXG7BsDlp9frNPl8ntny9fTNDsv59KMexM/FHybEDgj+jUWsY
L+JmSZVG7BCN6zfq8hTlQoW/zoBz57IvN9K2DefmJTa1t9yaqv7lzbAXsYE9g5Ls
GZRoYbSZgtZf3IRx6iytn4Q9x2ltFjjDQsAzBcFl8qXbGKqtsL4QXjgY8BHpZjds
mBvRurgayXFJP1vFEmzCEs2H/eklmjIPaYdsREQCgAgq77V5eCsny2Rr1wJ3IQn5
pKBFKCvjKFk5eAzYMSAP8RA5OXgGYK8zKu4sb+46s9WvWV3JQiU4k5xQHtudIzO/
JsCLsPTZ8KIQCkmjo3mL3ybszgWOdl1X6Vkv7B2zbXSpD7k6kMGN/uMWcFWCSs2x
sG1eM4Y8/thL0v9PUmoRV/aoo6B5hSxERjbKI6J7yiqcmtEDvriFSeJAiNui0fxY
iO/DuDVGkxYk232UHsc/EglSaEOfL++TcHpW/8nSwozeqz6QHkgg1ktSkyD5XZQ/
1jEy0ihFrcA7fiI4GSf8gq34bGMNWERCm2ekJoTaTKSkutjogxVVH7InOc5shnR2
e8DR4IyOMuIweamcSlw3MgoWIkNpEehuvtwFOqFzVnwT+GpDiMSEia4j9YoMnlc6
PBxYSDBvVA0wUgcH68+oIIfVXCOos6Sb702Xu7eiQDWS6GBHfpd9WSKRvG7G3wax
avysdUPC4CGk10vddQQUVf36q6+jEVYgFb3kpnQSMreoOHv+EN5FNRLHLzm+fwAF
jy8r33kQysExbZsVTJFL7iwX8WVK77PVvMwCe+JtL6cY2JYt8pRejVqm952I+1Vw
+/tw7AJTh0XhhLd9jWSvuVsCCNm/DrgNRsJ4vOTKStKLk1CblqiVV8dBdjoI7g/k
O+HIG6xGWTj6VnCMsMACe8abziWeMoJoi8fv3d7WxcJChbJSDj2hurviNI2+igYY
n8udrvZuqk7Wr8NOCNODv4SdhFZr/GYveMH/k3+1V6HrQdAwJ7yIYCoifRzbcUJr
fsbbobi+GMYLXNA4Vrt+225jGek9tEH31w2UCVbqIZnHhSFmp/7rv3JOe9L6XndL
44Nq7YdJvlrMxhbCuK4nXcOlQB40lWgK0oF4eIEB9Z3FSyGQdUHLxgPa0y+E5jEH
VSCFXGjTlYHy++Q0Xy8n5g+Jf+MitzbrdJCGhKxzCNKgyClTB7Yhz6fIEcBMefSj
j1CyDJhv187wvHH9gz01qVf9uwnQ+Y1KRjZpzau4WaZUtY+6VGpiIjCG9PS6Zpem
vRSRzxnurMW5vGikd5GrT1nnocGgPjmTJPdwGFv5DJEZl8i1fpjY/B98Wb3JGsjF
7BE5GLppEWS2RnxAHzrPJRNvUFA3Gs7opMIBTn0gFxlCL9FOMriTZ7OEgKUc5DBq
FmteOgNwYBXTCIsVy4jIl8SsmnNatO4jkypzgtuxlY6TCW2SYl2TcvfpJKfHT1gV
J/4WgYGJxpErMcXpx0pYMSMQ+othnQvmK3gYQ5SAyRWq1lKm/R2T4IPP2wufSuWo
GdDPfiyZZ5pxJ4TgYjwbcqC9x5UI0Mp6vwwNv1DegcZL5Xu9XIFLlRYbOquX5ry9
iahWdv+W6Mgvwis1bH8/jqUNL2dm9d/ret9m7vs/Mtpos6cvaqjYXn/sY0mKF289
FRrt0F5lvFSbUbeO2wH1jKjG6lAo2AG1zJzq5knrwbTUNHWtZxF8apLBruBhP4fq
5ykZrOeOWuDRhCo3CoxPlBRWBDTlFLKyAR1R5PnRJoncnX48XMwy5yBeFvfPmDt3
Mi3GfwbhwaVHpFaOJAegIlwK2bRJwulV+RbCg/ULBz6P4cPPwEZb7rhUBxIeq7SJ
SruO43m1w7utw/o+l1vYvWi02GM7ejEi1oGO0wf2GUHd7wxVctrSGlQvXfOpSF0J
sk5HlFedhGKjVRhvHQnvlXFFowVAVrHJAfNHmd1by73IGZpPtV/Hi66hXIkOnnaS
acIeTT+VIFQzvD8U6gTPC0dBzvluAomll+QWzSh9kkjX/fH3sdzSr4jmx8Qa4eLf
BPHWyj8wkp1OLYJ20iVNufZlqBWMS8DxSJvHmXV5QE0DU2k3nStzoQXTzK/nzUvg
zTKc4NjduKTo0Pd/hIzGeWB0W58wGoQ6MW/npMWEye+lSJ9FIW+e7HP42hJy5w+1
+OP4UzRqXGUI7N5mrgvcATsRbbEJ7VYemXY0tmkw2U1sQ1w7aKP73IP0kTNykhnF
jbNWPfvNn60npEpr+cCG9uhErlsdSAPMuIG6xlSM5RbfCQYs3iR7p1EhKEFLHSLV
PYUUEc79p2PHBRb793kVCrCVJlkbgYB2rCqJUGK67GzlurLuJFDNOSB/bCP5GxHK
qQZyrQF1R3MJUNydABxm7YlUoh4QiTpUIKUktmlLvvzmeNGlZ4BkL459HXOBxS2l
V8krpYW/LavqawOemwM6IV1q79UWxln/ziiMWIK3ROOPDwS/pWC/QU+2saOkAPkl
X4fLGxiyIsO8GuoEPqtjE8kG07bQuSQGPpnux9IdW1NFAf1jAu5ZHJBDFwb+igtV
xBATaa2dPjAwZksFWejIz43JNTBbj6QPq55wLfo6WhJm0dX4Kz6Ez8Wl+7Nxhp1q
VU7UikQ62T2nLi9SXFhl64jJqdLGJenS4s4cI6XTRp+tchDSX1K7Aufv9By6pzy6
Rq0tRhL57PRnBbsfaNOP0MVVxizAoTi4j9FzhZqgJY2/b9vC4RxJem5xlE0aaWJl
U50T9IrJ4qYCADfXxA8jJoBcScVp70r8WdufR0ipjGAFM2p+hyostoGb/WqBVGW2
2JGz9gMBbBMQ9hnWcCBEF9CW2tEiv41PD2f5ij37zaPbdvO/coOS7B+hyLGjoxup
2AI/iA+eKtfoN1iE/c7cvxrELlGreoV5pOeo3qSfyB8BtxsA5xJ8HSw81xbo8oib
uJ/JQR5wvoOaKh0oiDBZSbm6FaCDKlxtqK1wtodzig7TZ8bTejQZkoruPHMqKTAu
vN76FZS6Whai9YXP5KPDPLylztflEQfrFEQc+uZav1+5+4pfiKQpFx1iPWx9NnhB
oNT95G1BPNMOQ00o5d1VbAhxZT1Vt0KR5qX8bdNGHnmkeFa0WZx/11U+0vE0EDg8
qV/BsTbTyDekihdVU+IB1H+lo9StvCp6PeHGnZn8xZZylAcdXjL92Si5lTZCSOUb
/YC+8i/lOzhvGE1KUWirXR15NOWRnGVawNDfmtI4LW1shXz/7BJQNIVDkGxW7mI9
5LDCTIi45CPdrxBw066Ig5Y75fje+bX60FeFhTVLOh9S+MXowwV0rQkiV5FXEqIJ
/UlyhFoGrqf9ggjBsP2xvowdrxYd/RGuEl9wYHqLkR7B78JG2hdRgftK3wC6sAk/
tl66EkFnM1TkVDdWEnnH+GNW6rTCsEYrNgyv8X4/vo0MeVyFrOp7uPcm4bRycLfp
BjWD3/TShR2IBava8V0STOv/3HrMSfAN5z/kGLzBxzNVb01O6/RENS0PoPhlTnwX
i/BOOfEwupmGYeUxG6Ohm8LoQkD18MiNcZufvLR2Qgpfkty7qdFJqG6JNJDkIxmB
Eyn0w4LZCSGqGMmIO4GheDX8RAAJBZkaTMfkYcRNiDAXLzkYPArMC2B3lvVpaakv
yXiNWXqQn03qZGA6nKNjA1AN8StYHsja9YwZyn3EABagpuY3UVJrVC8OJkUUP/th
mZNK2ZggFSkDRPkW5RJ5xRxAB0LKt7wlRdAQ19oj2Wkj2hOZc+eFcXr2Lr1B4gZo
Pu6wB/4aG+AWSHwWk/EjjueNwrEuQzOuBhO29iaEb8xRn6gBztSsZ2wzFiYi3QlR
mwH/t0MN2SybFgIiaVnQ1q6Y70vnXyJp0lXTvF7Zn3hvvhDWG/cxn1n67TBPTE4O
W7zpwRO8IgfXVEGAbUzQrtCeW4ZqfILpfHu532gkvKuRwCrAIl+prz/6GZGyRNWC
38VNzJuxM968svBppOZyebjhn5riQSqKw1r1EUv+1rQ5Q/RDynfMwq6WowbYGOCm
ZskJLOf8k+X8Vo27TEKYObnHlNTH+uC6sj2fpgMJMV6UY2Zh4FfVURyymVnVDB6w
d60Ye+DwaLqjUYKtHBAQdg2LfKuZcOVe9qP6X0ANP/Bf4LHddLHGtwGRqsRCi//t
+nKjdvi/Qi6ZsEq8iog+PZTlTNkyM4OyW8h+x6/mGtYpJ0N54/jwWSWFItcNZY4x
NovfA42rHvIKk20SI8Dea9G2Lce6FKLjNBNg+kXXGkczulwgnQAZbLNiF+3iB4wy
BwxXG0f/Yu8TtUu1xpieflrDDdCRKNGJf51ipZMMXXGpKSERR/NNsj0X4GbiMplx
QvKY631v4+JOZxqqjIrC18IEtcLQdz21BsGcSrQXiycuTifReFxVQd9oxxGmeIeH
RkbWWTeeggPs1BuS3mNr4tpeJ0Mia+CUHWliZ9RjyIJiLmRAge+XrdrGgkXC0HO5
OQdySJQ5R5PShVJk3IdHlNhmaMk9+Lvl6I8PAofi4BH0g5s04MSOp6dRvY9MnjUh
xCwB8UoRCrpWHqkQsHLB/hxolQhB6TponwqGgIlFL/RlHKQeA/XaOg351HHsvE6v
p81g0MJvpp1JdT1q5/x2fjv04X8tGO4IeM66bemWtrBPANLHkOJ1/JDj2qo2g1w4
ZyWcfH+8oRh4aiyATiIGG5oudYqwDNZu+yKWtrh91jb9PZYbkl3RYzmnVOc8/yqd
0WWSgnNI8dESO0nYG+YYchWZy4yOjgbMGRUSgkslXxlFWxyF3IAfPaOxTPXK9PIb
KKKmloHAqozmDU+Pmf5OOhJImb3nlOl0akHHdY9bzW15Ho7Wbd10ukgJxIs/8+GD
sFl6hJFliTpwuI+BNJxG7ddV4A4VJXYttR9LsvuJpTqCiy8PyQWKZw0fFeabX2a8
V1QmxXVKV9JSMbs0oDSrLXQrEYmRL20YnKV8ZJ8gGzxP8JuANbgQVl9tVuouIwZS
jFgfF+GvEvkmCGtevGhOx7lMjKjqb3UNdLTTvyHN/b+dh+1aJPlqxPllquvXCMdw
i/ucrtLwSrx5abii8CS440gqfqWMERaaWEpcbYwy3NEKTIHmymE9fAJZ8yyalBTY
6+FuGeEKDy1OXXW33TUnImOWt3/Zdk3DbFTEGK+giLNlAOUqVGSyokPTjR2SRKBG
xoxboR1BTqJbh4dUYR0ZphcvnOANE/2LKEsKfvrDrsyFA9sYNG27uEfApQqbCwpP
spUYdGMCP/M2i7zO4YC/Oig6wmyEJ5q9wn1pBgUHmbGdQrDBQ6cZafE/GAVgrfmz
da/0FW0ZrsCrrFVtzgdG0OtaAb23RdhQDxWJAMp66jyxyxe72UT3VVRyTQG1yBy6
mSowyf09mrYt63k8WtLplhEX5sQ3l3d3weYvMvwLJpSojniPxvTbDr5CrIc2CJP7
iO95izMFmABddAHvLWTkSRG8fawnl5lfDW9EqmYX6bj8nBizRVu9vzWu6qcDpODC
ZPA5u7eC2/8UoB+i5NQny5CrtTB2Sn1ylcEL0fx38VS8PV2YNP9Dxcun5yrXfSAs
gbV2sMJOyB0uyqlhxqP0UUwRELlpudKk/DHXSYN4G9SvXg6b+rz+bVZX9JJj5u8b
uGo2sT9P+yijilVTMtbjuh4RYcacoiYsLoY+1mIIgoyZB26txabiNxUSs2FaQEFt
aufb8Y09yhgERABqAaPKCTJ18F+8qmEYHTSonYPQa5muz6PJRrq6RwhsK7+3T7kh
QanVtJnTuenayGjLDU2cS5SB/Fg2kQyRA+dN0lMp2dLOT8K1h07F4WL3bSVZYeA9
XgAFuQ7pmJPKjRCdFimVtqePkhX6FtOK/pjeOv7Uhkd6Jou2cgP7FXbmWmoTLCWF
s9QUikWqzXDnm7D2hRmk1p3B2+0ZTVaG8YPEUuxkhxOhQjek4wZ4Y9061/jii088
vT31Rglo8ee6iGKwLKS58PnqViweknSkFfh1MlW0iept+k4cqcSvuVGvP4MpBigX
CgKfelr+Q+N3WF53gwCQCt7Sa1CCdBZcNH44Jd5OycQ665G2NxNazcfC0K1/rDbA
dSt1Az4WJobCqTdjPEaOk294f7Lulc5q4MO5sY99x7SHQCjg/ioBNSfV8mCJ3+7r
YdwSS22YK3LpeJGjCRyJLi7OeuYyYin4LadlIONRg18wWCRowrvTTIBmQn0mW0Vq
uSenVpDSJsRQRGjaSebt5VEpfwH60lTrpXL3/0pCGRVSdO7CJV8MPuzlV4tsGegE
fy9noI1GXOpQfG7P7Ee/jhh1AazjtUR15ky41yFrCn3isqnFNxaGU4RwnW3BmNEJ
tK62iSRqaK5NP0HAffrV1reCntAx7P7dozzGIosP/HUWSYGHfE839icg7d2SBvvw
vwQg19Cbv6GW8rle5KyskDHUucKecn9t0fE3ohWwPjrCfcl9H1I45gWtyhhVRFZ5
MP1TKmm5bpNcPFgMP378G9GvGkACDUU82wxmk2yTa4Qf5s5h81P1IA4O+syUfJ9U
C2QOYT0lyU3oPFd+kB0yFiwmYaekEtGBW/53eoWrkZPIPMccIT6C6LSIOSwq0gFc
AkOofEq8JyKtCmGhYjFOIce6KvxwXEehBAhPf/8PnKXBEWAlyThN9awjBBHmNISG
j2mVALue7SJuuRN7n8dOxm6PA3kNEuG8lTMGVGQ1vMvzOi5BA18qwJOu3rEZM9Vj
cdfnQCoIkhEA0SFwEbfjFcoCpnePcHdihT7pfj1gqcQAhqP3j/jhXCkkCXbpspT8
/hCCiLTwpN6KSBgfrWPtPijZAWroDjhD8QRdUswFba+kvxGNX4e5D5KjCC8ZP3yA
bwwdulL/WxbwwBHZmsXLp0idCqZRNwmYNHLYEqqZUctTsRoDtoPkgXSKGY8/D8gl
IR8aga9FzAWLVs++LkXb1nv5U53KMlVSNi8RdV5cdxGZ4qUA3Ab9OM1BHIgK3zou
63i5Y73ZzWD0FfIOIqY9W0q7fL0It5tt322UCMiCBzBDZYYtSVumRL08qy+kKbnL
3wlsUW+6SRT/MkQHtnbw5wzRGOaA/ftdTMsw6Dylck6tu8nlYldO4wZe7DIWrpzP
7da01oJN9EpxjHUSj5Q7QQrc7QFMbtKcbadFFwcC4XKidWwKG0bW3hOnUHoF222x
KZ2lS4Db+W1lBvB7SIchgUmn0NJB4r/YopmjQhDZdngWqqsENg4CHFeXI370GlTq
yu354pnermVvh9FbtdFTNZ4tgBmDuizIaaH8ENWN65dJGOFXxo3chXrjbC4GiH5P
8Gkh7nz+EL3uMnaw9s+P07NM4sEjf2Nct0Pih+xtRPfagbM7ZAVM8Jy1jwAR1BpJ
LgAceSKoJ6O0nIoNss1KuokGoNfWi5XeIrKVnx0bhaWXPgc8GPUfbu5CGiRjkQ13
0jOHiEDi/WZttzQWCdFpO0KEPZzHmE0RiPU1Ws3wyX2ENcMw2szg2MAcoYjz/HqN
gKFOyliK/C5Nwm4NT/T2F8gCEsfuu4aWbpJ7rgwO6L1Q+sJy6/LeXiDHuToqeD/z
komxuK5XgRVVaAD1v60czyGVebRQzhPnwG0Cbf/7LpLuZTUct2c8FA+3Z1elfmpJ
7TKEwWld23sb8fILzaDNsESpH2eEQsoSjp6n/pRn6I5GZXF7sKljAcLl2gpYSUrc
+m5Hi+glvyqKyHyM4hNWQ2C6FeX6A986lcSDOdxy6FIy1oD2ZRC//iE8fjLY+bjJ
TXJBI1bGxE+KAK/t+l/kj5BLMza8i/9/dbKLtbk19bWsZ3QDPBVKzJfCl1iFy/Gl
VTrIzoCTzU5wJ/Nr1iibE3kd9HMoGHfQxRof9zpIVaUAdblc4pfqlLVveqWwiRhD
WzPmTM6lmVT2iigzYkKRtl5sH/pjlQ2Zh4g+9PETtmbiRYUuuqBIE/QrxjxuLOMZ
W2pGToI6ony9erqWVRSvWTyzd5LxXYyl2xYOq7Dj8MAlmqGKTBCp/TsyVrMuN/ue
vas1OuJGo7oC/saaLCyN1SwlPWRqeIp/o84KUXITudals27WGUt93rgTgyQpbjQb
wi7el28GAO2o/msE3E1Cnc1sUhPhyWKBOo/DsUqmxfT2rrlr19L1owVusbmVPjcY
iz9PjxA/HioX3Kt23WhGMvtd+M/QQqB9/W5r0TjMwVh7sGI0ahK7ftVQui0g7e8C
/IgVLakc7kyaGFMaGwP3T4tq3tL7sEdxRGReYKbzP6hBOa2n/Un9EEy+hr8aKczn
b60q7Y2Sn4U8yNrnZsdM9EYQTb9VlFHo0AaotpaO71q2vegnjubxBg0sQ8w1/ls/
4/hN0A+pCN6AlXh8bFozutX7c6CSWzuHhRGqntcxEnkznVYUUDbhMdCvVgw5M5bx
5DXksiLweryinYgC6qHIi6a1Y5cNsMg8Xw0QORzjjX74beVarLau/fYBJf5l27TX
y3mSrwtL0fOaQbjO/TlCTegdoAoUAu9/ivnNgcI/KllU8zqvxK/6xeJEByscDxqc
Ildlev1eCjyKQ6fY2oOX6srYCX1RFaeuR1t7CYd6G4oHVki/gl08C7ihWBsJaRKz
9yDcFpDjN7iknwZr4Y93CjDUYjDtnXgqDIBBiu65dmOQArFh5kYp7TIIkIGJjtrx
nqmRXtQ6JbpLNnr5UBQSV6ed3AwKBz7mDhzfVjHf3Aw+kO9A/b2GYhMWgULFHP8c
jWkIrC62jsRjvhCGLGCgmNmyRF9elpp8p2DoAksxFTT36UXemNK/HtggcvBFGaXs
bQk59Gv7M9V2vnvmGsif5AEQX6Bots8hLxqb2CgGyumSJiOPksyZeLyLVxF8xxyp
XH0qhZmYuQBDrTt4W5shbiU7dsJWQs4nO1ODm6SD9qomRKqLLfNarnNoZFMGp9KT
mPViGAXVRJwjMpKoX2a6E0g006ZMkoFo8LJ9BGej14/2tjEs6Qa2Y/W2ItWVwZQF
hf1CZGKSPXMQoHBUVNb3oq+WN1+SAyMq8OmsPfU+INvZhtAusHGU5YizpvszIunN
443ljLWEpz4Qv98zvnsGHaExMoT4Iesm4q2sGfGA2/h9QKW1B6EXblKATEOOJsvO
LqHNJ/13POWB/hU90kyVH1V+3eUbM+CWwst1MjVZ95uDclUFGuVYBbOr0X5xkL4I
LDlJtdCAYrKi+4Llz8BDxkqpluhMMy2ISY3xTYOa4JGXTq2Kddzx8667NmcN0xSJ
RbxuOzuHIMXBqeHWktPskyuoysi9uY9Lx8fl4rpP0ZfK/r3AH+7EYKwO2et0QROR
CT8I7OE6N2zFKbRqcCkO11+yipDjWVDcG93AHiXhsurYWCacwvs73gb3ZId9dy0O
N/mYCV2ep2G4Gt5ucJEG4XGENg+8QnA3jj5aB9fM873u77fyO90ZruYuNe8UwIte
yDB8/rA98MPlTj+PMSFZKc/mirfLZpe3Hk3duPhRW2PXGN2kPfDerBrfS9PSgRe1
Dz+2SmXwNLNO72NAkqLVmktgx74YSbEWvc/xUSlhDMKmlQew3YJ5AbDpFqkeWVEr
IkjqcLiU2IQk/vyGXfxSFRl3gW2Fiaxu+g5WU/lA3BQCkd5W5V/717JMoipDbGQ6
rL4qB3QS2beC8pRWhWr0+B/Vzp56ZqWD9HlNpD5hbqyEusA2t8ZGhQoC4XjQWcPS
AYdJ+1TFkBYG+TASi/zABNbzQYwJyeCgZXSlDu3SA8LjboaD2xgzU5ut98BKCN8+
nt4XZfSI/PaM1UES5BLC5rxeIE5W4Ot9hU/7a/RHR+ogvktInNaHNylszRtTJE4N
6IjpV8oAOYJSAj5wQalxJVME7W5/PDM65jeUhPAtLwe/Mbvp/M3M8TNy3D42arQQ
TqBeEKHGq5dyIw85DAjAWnB1WScaftXzvTxLzCt6MxIf2DzvxdKFepdIcjAuCZDC
EkApsL5MRT8JVCtCgRV4fxSYf7jLOHQHN9Imrx5IygCfHhABtjo/Oj5vjxCUcFyp
IPJ4PmTuvwHRe6wMxslV3UVjMhnvTQUCoxxe8vcaStbhvYEXXH9gY2viPnDx6hzr
oH8pfCswtW843dBxEtKzH/uXm03bD5IaTwrUqQvxsAxTJQXKKv+ty9E/AjiK2PGN
1ouT/yT0ivlVp2kudSoBOLAaOmpp3nKkj0JGGP3xL60vqvxT7XQajYF8uiHlg7KN
PkKgvfoS0L17bMWrkDK3CgqWgIaqnIGXHXA2lU+93jp9oYrI/qJTcVYeSDEKYYeM
TymOlJczNWrvk10c7mIO/CFU0Gat7E6x0vMGNKgm6WjGCQfUgYbQPyxfg4y2mQWc
`protect end_protected