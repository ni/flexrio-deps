`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 45040 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
Oc4fq76CzL4QYVrEyjSlCNlYxeYY5ZlvWbKLL/krBMWo1pbO6liVN9QjZ/8+WT/x
Qn3c+RuJDJ4LXEAs6/ebg1nGMMRtxDPbhptGtSxp+uYOlSzREatarHXbLb1vTh8N
RaNN2+ccax3Y6xDibu8S64ZjgSJr80yRzmcrVEL1UnyExAhqlH6cA2zGNc00LHP6
KHaKqVCbMoQ4M340hqhT/uGNWWKx79mPk1PAh+iG3SwG/GwB69k5rC/yroOsUO3D
bsgiEQmnvppVpTzKSKOInNlRouONbGYzckEKZvH9XZHJHndhTZ3QZE7OB3nINC7L
xOsUovfLaRbdW1+L+kpJdzR2dCfW2pPg1J+Re9M1DXDgINUHxTSWVv12PyCSFzIw
YwVr2CeswBG9VFVkqPmRBv/G7HM1aWs7hS9246apwdeYYn9MBU9IIoB2buLaDhPG
drfnokoWgUpARqavlxuG1uuZqTYbJ0dUfulBIpl3C4qmQYIoOmOjewtXYaBxi39A
AifqtwwQSBrGJ5Xa5jGFi4agbFPd1DZgLkSuJqQRsciF0BqKv0rBUznYv1cVEbH4
dZ1DYqiTgEpYYTr1jrId23YT9lHq7wFjVq76D0H/hYwHL5WkTRzeXAkOmPdkGctD
3pCYBHypDMqzDAM/a7xUIwRYqLfr1WaImIwn/d9Zf3evMPJGcqyQOWRJFu9lfsyo
FaCHiznh4AvJzGjlwAxv8aKJhWGa9YX8C4AQNXXyAxE1F5Df3uGNF57jUsfFEMix
8O6VOgKV11bKZATpfaqt5PZ5cvlxjo217K2F9vLAFgwKxKFkM2YgF+aeDXrAzqaN
ZFBWuvAxHe5T3sw4sJEZ9D8CWXCIYR25I642uO5TfEUF5pIBbGUBj7vNEkco8Rns
XinqLH6uxxk5tEpi6tS5kEd/o0gLntxYRO5VZD4fTtchhYFY83Z2nMASsqqNVRHE
RYGmB8Wu89LhaOQaTzCrZ15qWw8pe+3MN5yul/+bGQO4Q2ORezBL3Zn+OhvSMgPr
SmrJrRI4bkkMlpbAcvSsDWxf/btVVdYASI4D6sJ1HaktOjuMDCJYbxsIeFpwjaaX
eC2Eae0h/U1V+Q4bAQFRfuchU4NUt7ogixBXo9klGGEI8z/CWk2NzCa+7FYlU0r+
AEFbVQmOzd9O3xj+JlR3mrqorIK5Ip7etVkFIm8O//lGRB1WiwufCxLk7BmHfEc6
EM4wdw6t5/qATsrG3ICjeojnkTzm5BOxNU5O8zqVZPl6iKzXUTI9a8TPypZp6333
H1OMUfX4c/KAGkMye9IsEE8/0FljpU08UISlZ/0h/mhVCbZpkIycT03HHOyTc8Wz
0ZNWdHXMFw8tCIeIuaT7TcOPHo+9fRuN5wJ/txDK14FJp2LOn3knF3efcq8sMr2m
SK9cwa3/3eNAwv3/p7J5+hvGaTjaWupSWH4ToQcgFQMWWVDhAylRZZv3+Dl5wAuT
fb7oE6niJoMLlEhw8ofayfe52H5phr92yrCWwJzKMIAAjYiHN7kNg5RDxQpIAetg
PPlG8kK/HKsT4ZJkQm5Lbsrv3xzKl/wpf4ELwZdwMj/jB9Y0Rr07t1XcZy3E56V/
xtnZCV8b1jwc8v4TITlpzrjZjSItxClOl7MnUfDNWZc53J27AL3cFxrcOa+QRIDb
d20uTAHT1BsC2DLq9OS6TxXFT5PqH2aV90rfR5U8bDhX0DXzLr7IRyEGZKKmCIzt
PctvMaRW4VP0NP7N76YG1o+jhxYpu8qcesi1HTH58rnuGTiUk8I0gLIvI+23snZf
ZWXGkRqsyNxxz0BiIehRKUDYyItVCA14iT9YGsqVgO0+fp3ndwIW+W4MpgSP4UeU
diYD33bwht2f10zC7Cq4LkKzqPkZArN1jUMbVHnXHULwKsQSndW8B4+YzHlQKuOx
cAPlZvSqUms1gp16VTLMk+LJVGJOFFugyAxnJE3+w1k1dKgV3ni6MckoddLF9eHM
g438VX1IaEdawbl7PCJb8b7cdQiUKxaRK5/Bvtg+vRANeHajj0ZhIT8to8BF0n1m
nSdvmDJ1HDKLw7ReRIdlurRi+SPxr7EiF2cvtjNNaiL0jVMAHugd6ihxZGiEjJmW
Ceg4kozTwYsTdVOss+aU97I/B9Z+2xYbV3znOpsYcrmEfbrBBWdmCiGKmtcouhjI
TtTJCOvcb7H/GKwQmiFzBbv9Pn7wiEdls66riZh3lPL/33mp9fYFIC7X+40h3p5O
duIDt81kHoxS0UyG8miaIRn5uw56geolFOigKZDXDDeMag002So2pGaENKrx5ZOo
ydg777/+Da2EdodmWWV8DbqTWxO8Q5NcvfbWwR1YL46D1leeGOuGeQm9i7nwvlOP
oKAzflkkCaowlgppF7GqovHbIzBrvDCYKfkFhIHf6X2IXTzONIQ8ZjZlc6Jb5Ofh
FLZVSSuUSnBqDDS/Z9d0nmFQxkUhUHVKTCjWk+qWVEDs/OXMb3cc1t3+HXqYXfdq
SzfhXM3eafIxzmYYbTwuGXaaOXc/3IP3tPPWuHzClYSSi9JYGVPFeid14bpbmvYr
skRvo9ZrUrd6NtBVb/CAi3tuAtTxQ5N4gYSkG+FZNM50L58LivVHgjT9CvndyPjc
60cMmXfnYturJ3D29WfwjCzpQZJyFCUHKImWd4ec9rguvAY6B59YPq1tXR++xMd7
pdKOI2IzMZEXytcxmOVKHxC28fH7i/uz1NGo7HcQ5Czpm5q3Scl0hDpKl1pd6PMi
UZE7hV4ThZrVF+ZtON1NN8F/yBXcCZp+xQqlD/clqDqNX0mr1FPlfc0HInvSUBXf
D0wzJ+DktSxZOrzHyQkMO2uwXoChbwQ+Wp5crkA2TBb8YS2FiLapDYhP2PN0IuOF
okofB7wL9jlrq6+9IhshWC88YjqRf24N7aWj3A5UQVWZhh1VW/EcLSkVGgFrBNPy
mSZSkKwSSGqq6ayTopHJ1v/8FNch/LforH9nTDVu1jE8VgmBir3nQP5x3awHE7gC
ggQITGytOlDMJwdA26GuNB19JC/4fN2folQ1gqX9t2YLiYBPG8rvrKEZAYMN+bId
FeAD8Mj0L/mh50awTpxkWah515f9x8F1fedja1k1lRHGAvVYRdFZwRuJ7uCw30zS
RQ61DYGJiPI5jxw6kyfo8VGqWhPkV59+FmrZ0zCZIzPq6vppYNNUzCuiLE5pXrsK
wGnpsU9bSzNpvqLo1NvO65UQ7kcIXpOO+3xUVnul5zrTTwqJGPsnWe/iW0oJZOQr
HIkaaE4qx3NfTofiY7QqhfksdsGvpfd0alc/VP9Ox2Iw8NZhrX4enFINlbLZBPPq
b9TMXGVUROjWkxrTyeqgKkeXYtYcwvaaS+B+DjKCbe4Uy/t0mojJl3cHH1vKydqI
hTkBlwaDPEDQEOMf76G2whg8wl9heFFidukVO159hO3WF5tjZtV7wB9/MOxCR7oe
/AGozNhqFMTneWhB4PXsNLRE7KeOJcAnXgBHoy16EkVknbvbDU7kKsAY++XvRMpO
6YHt+VlgmaulnpubfNg7r+0wECpLjTYE8KMcx0RUFqncH/nSGlKw1tqRwZiSKCzm
ummyejb2l15SgdK2ZhdDgoNCn5hd3YEsy8tgcIwFBNUgsY4AWprC0llI3pBeF+Vo
8lvFCcELM7Dy1BAPdoqcDZzsnQYz3SSGL9XGLSNf50U0CT+eaToi2s7tgp3auOXw
3517bJWJaAIAYfHfd+Lbu/D+z6Ewe8mFZFXwg28vk14ghMlsEuK/P5C2imb3dxzY
SfUEuBoTX/OrxgmRffnmD+tI07IaI8O8Ckc9sgo6dUimKACaqCPkJF+lptQG6BWV
FuxQ6v+t4y9MUsjlstZqXP+ZSpbbSp8NowGIviQS7ilLaV8P+5JQ2YLsL15hPHXN
5574+V2wFWG947Rxy9BplNGf3TxdNKnR+grZUitzqQzchJH4ce4nhdOSi/pnQFSy
KkuOMCF7FKrtXHOfeCYYUlIY7T7tRQbtfGGtCW+qdVMAnp9UHFXaMs4l9vaUN2m0
we+qciElEpuaSKInGJc2IbWJ4lPdcqJF4bBVOeVisWRq3p0mYccdiZFljyYFulx7
n7uTQ+CA/Bd2/NAjPYucLf3MVc8gEAOJI/A1uSeOELzDE1BX9X8+dOY+PRw9g/mU
cQWGtwzYbam5ICFg6lilE+vx1nSksuLd5usDlRWI2V73TEhPZbjfKzydMPEoeChC
UDsz1Ny9dJGjfcS5w4Zf/Hk4ehDVb80h7fWRxsQ5RDlDqqc0oZkYLXQcTPJd7ZpY
YPqUDwXBC3QHX95BedwiSjELPZ4Mr/xvrjCHyi7sSiVYTunU9kkwOWVpUTjRUk5n
C71IX6qbG2ZZxTXfRI3/2mIgAGI3MhBjJxjCX+UBeU12djNuaaFN+1bqKg1Y6Adu
5Wew1bXtSeeR0hN4nVtEICC0ReWMtEckhz9rSllF/L1h2sCvdsMSacyB1ITeLpaC
1PuKFtS4gIEu6ILZo7xe9L3K03qgtu7ALKvwMBEPtdpvgUhQQBeUXL9YwFvIFIRD
z8DKXovLcH0y8qFy2EtT2GLKnW8BoSMjiAu+qKA7yAGXWguuE503zuQ/x7QIplvZ
OJUfSBim+gitZ1x8wfcWJTkQnGs72NFbyugVWWbW/25ZHgaQXPakFhPo39TkVw7K
LLt3MHGj+Iz6CSCLc9RthYYWbdpOWEklzlMg9DFArv1iHIuBml6LWBkts26D0q/4
U1hEYzWPUcjYbNvczH/9LXhi3UJ0G1BZGsQ/tqn8HgpU9SPpi9+LvXdSBzQF7TLm
FjZRTf6dZdW0GSgBbtHJlrW6RiFGGC4DhgXg76dIzVka2TZJIwjEM/MdeH6M3wAG
Z9nkmr9K/MExNwT8B0wa6Locq5ih+EO/OW6pb+e5NhHQPZ93XDHuW7yD14733JMG
c2pPneKlRn4B+7qv4Tt8EcHSrF6gq88UB+rm9N/Kv2EUSIH5HFyR9L68ODUAQDQ6
PKGXXherMZN2y9sHff2ApXw8FEhE9ZnUPMwnYQarmlt0L9/DKqw1Y7tqxX8XpxoX
DVZ5nxKu858X8wyrxhbFiq8jFBCVHno25we6NWIC/z41PqTKGC8JxY4l2dgPLaL7
LpyOCckqmeSvrskOTPxDG5kvb0+nZBXTPAtQpH9p7+aMyCU79zqvATNU9Yb+XRJq
UGNNNK36DXrA05RfVTbxrR4wAwUTK0ITA4odTKu8lPTjlNbQwVMYQOBBlwoIO9qO
c3PsxkYwIY1m3/OQgq5s5ovGxaU5ZaCxZUugap7EokK1LioAWofwbKPJedqU8wy/
J6AIELFPcEqcnQSAwKrhmL95gL+siITRuKBQNGDvGXezyAfYyTubaVXSsv7Y+V8F
cSqxU8eq1GuNd4VxS5aXRxs7QubxdrLZ2gvQyKu8HphqRX+ZrsDLvO/DlsHv75ss
WzSU65WxrYlGuFG/6zgKSPIqMp+3Jd7S97OO4GT2XkNkLcu/CwmyJ9SnAOqS3LYD
03mADOcRgB9ZACnMn5x0E0Ghgady3zksL2oCZsROylC1cTsECC4ok1PLb91+RGKn
rQiX1pCc4ZUI+wHUUZLTnkxwxy6Ua5ZBokJFiS6uQ0pXoLjBmT/WVt0zEwjN0mDc
JUZ5l2w4PTWEvPnbqokD3IXmQUa0OF4IjgypRtndoAMf7br5v6gHcMDhoHdzQcl4
jkFm69sq+RRNrWBicizALdMlHuQ8nKTVE7IJ99um/RWTnPYntg+QwNn5+lfnUCRD
AC9RdhEGezB8u8AD7N6rSYyw176KGBw482KogiUETSbc3kDjBjcVfKZLA483M7e8
Fbmqrmx2CStX7oYqAgNHUT0XpjLC0Rkx5gCFRrQgucAv9Cj+zFnBPJudhExbkaXj
sXoAwOvB6bVd9p1FoN6OT/cvKpy1wnh554+AWSWdDWZO3pV0QA88GKGnU+BQyAOt
YbgPFAwpNDh3kml+gosiYthNRvHbnbz+lQiGqhNHR3IE+Uf2kzZ9dK5nJEOTHwc7
er6/B6XYqSVIqGVZUCGnqL/c4/osAta4oJiO4cHx3JxH9sZi0Vv755bxLuM55Lv3
hHkhwZ/seQnnVxb8dsyyniT9b/2KVIcb5h2ZixlwFPgjNHvBTPQG+zv1jchan5f2
Gut1QnJpB/z4F6GoCrtZqrH/RRHwvCsyH6RjHsospSH4G4AwxnnSxNTq7ngd6N94
aLg7xwRMPsizmQiwd/t6tw8xCN/RzFeLLoLPd1hVaXE10xrmtLFJjvabtmujp3HK
hW79pVVwPkKVHt6cpbU8wzjauaGRSSmrygxxP1vsd7mH0nrsYFMEBh6cVkylNzo+
LhuJwB+ak/gzoKImfXWLA03Pb44AmXeRit2+MHdU9yI9G7PyMP65SQwpDv48U/93
e9MMFWB3dk+vCNwhWUekFcvs1GEtKiA4tmyQwdyyyxOibtMY6wPbGh1NqYfTQKQY
B5BPdCVOCXPhp/ZDzZfxDnV6zypAcYJ0hcriC0hkfCJx3YZiAITZco+wu1qjqB01
mh/l4gQu035BGhv9gSWwVfebQmbFCRKwNNMOIYPtkyxwOcrkghOFHgnIjBrldcwg
Vg9AG7S6olV9WSXqVPhA2dbB3NHz+lB25dRwP7zyQb0YivEXqmokYGc9kP5H6Zkk
ry+vYd7UuJxlpTTBpcF40lVtXRRD1VeROhSCRvnRA5JIDYpLGRxct4jnppeoAixn
+soG5h6pQYxmj886wdLVls2U8wgSPjwxYPYTsdcv7AC+pnWySXbjQO0AcYpNs3bf
yVJEoWv7S0bzc4ZiFKTa0mgzQ6hTdRDGPyLjEFIXgxtbmeTl452pllsdI9QEQMDI
bamGdqr+QTC05huAk6XdcPSBQSuTF+nu+DFK5FNV6aeI5pQdi7EzNHVikCB19KNa
vD3Vh5EeewC+4cmkIKWyXAkimzrBnIb6x0LpGNgi+Gc6XOmvBz3N43vR7gM0xbks
izJzDEU30KzToIOZis6HooJo717EfGUnD0Wua7eordqGaFIVlWb9OdxAoYWJGKu+
qS69rLhEM5wNG0SzA6FH9cD1TMj9L17cL3CDOqwgSZxH1eMbS6U4CI3dK2oMAv2Q
L3pIx+BfO/Sb0GAJkTLJr2EVfyhjNofCpjHCp4DD4rzHDTLz+HRn4wyVRtt1uOpj
8Ye2eDMPhEdSlc1ToX83BpUJYnfwiDbiwPNoyj3R+KDKU0Brt2q1V61wBTG8CV7K
grivbRNBc1BjFs80X3yhwrmVEsHFhxf8A/QCQVZT+TZuAYI6ELdsCXjTPjT13/ke
kGRkK+k7BGsHWF13VqcMByRkt9ZOwbh9jSITZqYMbFtP/QozJY30ECasRLUlVkcU
L/S3gtbaL3wEd2WCs/H4t7KZqxnAeOS3qv9fyiCl6dcOgha8UHvXIjZeJceLnepF
JkrhybfEWoQwWt6o+UlBEF3sOzIxAJQIbdeteGnxQryDY/cZxpue2Sod5FwJYoxk
qsRG+BSPmYR7miXRXbuJLuVS2Y93oe7sJ/S6IMJSYwOhJd8q6hG7i4bXNqPkqRyS
6DEdwopiwvoB6HQo2bRJJms7Yd+piMlxycaaSuVd5qLjxNYYJxXQqzyGDxaIhJ1Z
Em3PsFLUTO3N5TCTdTXWa1L24L91/oISQakbAhRRKeVA95s/a1jdrIshVq6xI4fw
WniNjuOWfdjXxImy3OCyyytVW51JPDfwEDf9cb/eDrLOOenH2c1OmMhBENtAYotp
DMxD9R2ySrAhn4d0qestwgJSRPbGyNJdxyPSIVh/8G923XGw1zPTq+C8Wd5E9rz6
mN2mNQgGXn+iDF3qnzWOzFV3JSL6F9ul5+daIirfmWcMiqnVNQZMZj2QM8XrIqKA
omZBAZO8A3TBSdcOiQjzPNiLT4yT44uwsVuZRIQu6Z+z6GW/I2CJBcz1a9dXiCt5
1VaK8oLH3kNfctf8yzkOZtBw6AJNgqYufwvw4CrqjyQSqeTKR42ssNxtHauQXuGS
CGvMNxVKYnVwn9bzocd6F4F/dbMfnGc0uxUdpeI+BKNTmxXc9S1VhRorWY0Qy7Aj
DYesoWKsep0FPw544oF66h+lEhyhxJz2kH4liez+EdmZOT5OpZvA1qbl+KJi0S/b
i/zg0QtC/OceuY6d5AmzuNkKehMeZYBfQiaeAAClSvhXYmLWxOekXeHUiG9JrXY1
YQbRJevMkHE5DUD5ow5aWLMwFe9B1F9o4kLPjpEFCqWcF+SfgdcG+NuuK6Fi7Q3D
l+zSyFYKRUEKXRKv4RkqIGnt953+il9zF0H31L1Ion+DPrluC8rLq+FT647FBtrq
ZfEi2FpJB5hAbns37UmEMoLJuoZ/C4ejiFRDy9goz7uLqy0HiAqSCTkAmbaACMVX
kfHHgXJxxJZ++uvM2l8CJwUD2rA1uHSOnRj9Yr9o7kcGujlXeHPVaA5IoxAcAsR1
jIuI1KNC5rZuldG+qtvvdnXTRuSHvTWMGLNFyINee5U9L8l9cxO8MjJxPYzoqpGf
KyFegV2KDjX0EnHKURqzOxBONis8Qb1rpadjWNpkNy8CmxtWCwsPyRXxdFa85Jsv
oqI+2kuuOX5Mf4dG//beK2iXvBDHR7aNqWDzyh0MVr3mWfgA9BelnmGNiITSpl3Q
QGMkLiFzKTc5iblbYQYyJgRWr1SaRe0l4tGlwiLJS31MAUZK9rcRC8kmMuqiwqRY
bfcO+9lC1hErvJkkmP2b2KiVgVqPwXBZ4xaArnKgGUyypbKMHrs3xUO9G989ZGTg
H1mk8MzsmN/FFMhPh1znH32Dg2uKSrTT00EyWa4/yapK25z1LGx4/DyVZbOY/AP/
SbSxSH/8fKDAMNYTB9sA2dqOQuOSrhBqlBCDUgmJ07x226aOI6eQMlTlgtdIxtQS
2Ubd5P6PRXz9TFJwY1qxnhahJIJvcK1HV1DuNd5Q0+ATJAuSHges4iGM1/iu/IWY
QCtOn2hpHjujWIfmZKlC8ougmkb2uoVqvKqLYcLAhWFS3awulZFQlhgNvPU9EDEP
R1OZj5WrEk2/X20CT8UaTOmS6l2JrUOOv6yNVH8IRjjw8h7aXQdAC6Tp/tL+0s9P
7vxW8SyYBncZs9vKELZbgVX2NXJWYn7glz0bSGpTkyifHVjyGyGXQmc3Z9Hp4yaK
dEtGZoaK3eAxSWDsl37D6VZlA0qE/1orQPyL8p0kLNGQAnBjbBjH4JslC1fgM9hT
cPlfdMZs0VbAp4YvvQSWAi67xNJUW0bVKEwhRnJOiZSKqiO21MbDjrt+ISW7FGjH
RuT51zTNfrmMelBTFw41Nm1WItogtO73uCGiVx/4HTgQjPpT/SqUbGSSgy5qpnwj
7OsfO08DamDmZHjpDqYHzqw7+MXsAfoySk2OZCFpIdDgFQuFhS0CnScEJ8d04UF1
vPGTqm8bjOzv9SJENl1BhfKCr21jOtulCDcNgqltNGG5xgR+wkr7dbxYZmhdfqKf
EHAg9Rbaq9j6bdroKxX5cq52y5UoMCfhyuvdF/BP7XV74gtKm6986I0bJnvdX5Zv
SIXWa/v1BtsUqqaGCwX+NScF2igFuInHlI8S41zu/yxuAD+AlbF+ee7wBFzKu0Bk
XyYpGAqTg3wwYK2WUeAo+jgsfXbw/ofFMUrgNivh0A17+FuQsK3B9T8AQ8O7pW/S
Apfc/3CMYOCM+l4j6Mwn1YbxG5Vucvi5jixZCDYfhuVevzuPhcIoJBJAXYqbtb+q
MuPPa4B1IiAXIOBMLv1Yi68mbvSqd/qlEIw2OSnaoe6A3jMmAwwwb54du5JjMpu7
sPXeIzmICO1gnTJ4mPiy3xTXkObTyxDNpao2mW+IrjvlU3MPto7r+NOEq0F3d2rE
Z5j7RJgNYWMJPfPO4mmYTQ3cbIjVWGkI1AN/WU31CdxmnyOD3XrzLANCxmJ5ITdu
ZNNQSy2lwcDyRIn09jM/ii/0BE3m8cRBwnMkkbuhOrgefLTYN+qHWO7AQ/RoQ0oq
K7VVaVZczb9PghWNN41Pjt6rVOVftmBd6w8CovTjagbJEPMXM2GIgpyChqfrnguh
mkjB8R7L0xN9fmPvNeIG/dfvbz/5xDtMYfS5PCsy+iBQVlhri4xmJ99V9WU+Pxt5
HiIYrUfiER5eSIpJ3JiEjL87EPwPf0jlHX09zITMR3sgk9kTBvvQuVNuydpfXrJK
J6f8uBLaTKFGb4AXbnsqNgRUlkRQwcz//hQCzMgWBKWmK0RBYdwIPOmcyZEnvqO7
5EOGWOClIBUKGzsCFVw7AbyiEXm2+tRvqxYQgEj9O9EkFo+jyX9QCksGJHbBr9/c
ZI498CUB0vUYCjo//0NMZdGGHGaxFK7d9A/wdWn/RTEF0NYLC4nZP8eFUhD4FzVf
VswTG2SMbrFlSPRJRNTIYU6YGTwvzxfIWJrcauQeIGMz5uUup2sAYzHDQP7LqzWD
csbzBvoMeUkp2BNEUqghMXeGb0YKMukvbQztHJu5vVbWxCRAoa2Pnk7hb0/7vZfr
V8rHMR3h0YZu+2Xt9VYWWjLyhBg6u+FuBu1CEt8z539jXDXD20ukiGZgEyjKgdtr
IS1G/CcHKmn98cp/Mca8rhnOgemqMEp4FEkthybLMoymCuE31o6+RU3yeqFXq8f3
MhT/DC0oF1QIDUEbOU2uEIwakBujRYcwZMAacz/srvRSu/MhJaEEDa0KOSwOgB9V
wDbmtXgXKTYkVSjZkbYN7B556mDHcpwqyTeyclkJzjGTGnE6MD0Q40R1zaO1z0LW
Nzrhu+6DswSRKbJGD95P9EqEDDsAzZxuypL9hQbqI69XPd+zU/m/QmJ6rKHImcgF
5WfusuuCTTfLdXYoPWuTckboGRMwZY6t43N0x/9+HWRJLY+i4spf/sV2AyE9V5Kz
pq2MBhWIrIRfaAJP76Z/64/xzzr0EB7rDYLeHdGslHhL5TtiX855MyhMTDaPWqeb
Cx/KmDhBErr/CF2CHYu70OG02A/g/IsCYWLJbSJRxqH8QSXBEK08HO8RpNrpe1kp
wWAPuG9Kz5KrOu/YheTmF2IYNo8KcuYagIyAvW6+XG0OSEBYoDHUcr+9W+kEib94
JvekSCY1NBChuDq88nAfvqC2tY+Vs4t89A2u1JAw5gluF6RNnQU296Wp97HkSqBz
fQcTSshrtLMBXTIa83QGF0fTVFsIcbShdD6ZkMJFR3nibkrfzUIgo/N7WNu26A0M
WwA5bCRvkt3nqkA1zEJxTwnjPWvSG+X8VGmma+Jd37Ka61/4wKCgSwoXG+KmUaFg
K6PKwWui8rvMDEavY/mTdC6p1dmZxjkOTxQPTnyUTmjri/BeTYFk+BFxjzhELVzc
e+IyEBT0AimtFJ++fzSWK/5Vh/gMtuRxbjxVgsKCt9r93+s++FkIRzbbS+N7DjW9
5ndYGL/rEXRQYZIvSSZ1pkTXql63+ASDhPkQbo5sftTEXCytA4/WB/yrRglMVZ+5
LqrjsNz7V9Q+V76ff2H23CDz+Fx/w9uEQFB9+K6wL2U1zbDBJPVMEPF15W6qGGD4
Vuci9nwDfuYbfu2OkSuLawwSn5nvyVta+J5JoyZGXiw83FjkT9Q/qGgTeLUQIePw
8TZSeR3N+9zvj7J3JIT3pr0bGoCT+63r/iALD22I5S0Yc012k09l/HSs2AOW4oJu
qF/QGL71UJx4FvlSqWoXdl98Y60lmsmWPdlpBuN6Cno9j/Vy14PHt/ISraodqlPM
QV1EVIw3ITaT5x1nUZ7EnMHWfLXJvGsVOJnioclILqVKNCM5Ljd3D7pxo4PskwAo
IzzeaTjEq5GKq+x1HcQwHQogTEjk8Iu4axq3slEPfD85ev5eAAk3j4gdExCHYLYT
TaNmCKAn92QTsW8r1RDJwXa+gLee2y2ywno1DiBTMyOE6l2iSi8dMKzL3HWu5N8J
WMcku8aCYOZf1DQaD9yjzTGLcXW3kQZoNqsXcU+UU4SLH69nDOwzVLod8W30Xhu1
vADK8UAk2pheCTc+UT7SN3/MYqR7Aktb65tQXn5Ra5MBDTyPcD1x5CEPXlWVzgrR
GZedY3pmEDIhbFwuSfEotQHaUscW6tGPNH2gnlqdAeac2LIIP+uNPA64JuP8gfA5
fbviDfEZGsfSzKK874OpQJZSHzD2uGfCf4vJ4suXdMP5jOb6WiPQOwjqftsZ804l
NYKCVlyql33CEkFvrgP+IHuQ4ZEAJUDNXLNk0cHR/stioJ9ukniWcdZkUf5EvC3S
NDXZAs8j/8jYZaB4SbZ+I2/n2VkcKKszUR1i2J7pagJjf4d1zzjL1LZDS6Fr2QGH
2vJOjzSu1c+ba2JTrHeM6Upy2ubz4mQTEffJb+LyLMusRf0hN4UKM5fqTAb6/ftT
X2q8QY81rKZ8fpWYF3+CVa4DJKvMXsDaddHXfdK2mCV6vmZWL2eD2JMS9/PaDCfw
K+ecwg6O2rrvoEQJK9aJfNeLkj1Jgho7x7qH7tKuD8zCX5JYOnrCKBHPyo0n3i+/
anSrO85IIIcer89b69CXutbr34GKQnw//baFDk1OKJEr3x3zD6oaDln5GlniFDYa
M7ZCZd+/cTTMnnGnW64LTEJsZAG8GKr93ed6n8VJqhrGjnQfJZWuGmhUemBMUZZL
GuUgQJEnYWyBceY+DZdcaUJttPDoQTf5hvxcfQqdaHElA7UDxYT1h1WjLB3FKz3g
kzS4MLylFGnSH4VYhHzXRIs7O0lnDQ4vn1ngK4gaNKQSE6X4PBKdD3DzQ3HV6jiX
r0TvP5fgDOAu3mxzI/XdbvG4e0Zi/K6+rLK+ElUgJzzet+XYNtrtSdZydMMuOpM+
tp8JBKh6dnaIDMNfJRhS4MnqTpTxpJ9HIh+u2wFtzl9Q72AAzSQ9SkEt1l5S1w4V
ZVVnlkLws6aWC7o015qnlz4SNI0RtuVcUYTOFqlwRrCfvc7gxtxhnOwBQF5lC09V
TTJa+8X4ASiOqgcUrmTGLI5XoBdcvzFo0ekQYdBNter/JwiK3+r6v1xjtHYsut44
dfYArOsM++sNATMhy8xf8tvsihaoWCjnzs6Zptvl9w/s6Vur562mnuBKOdV6ZeMb
6mXq3ZZBMm/pIGXEde8ivX099XCgBfixvc7eI7OWjv0rrpiEmekrcu8RGaLI/ITR
7jTuDkHAzq5Q9DzC9oAvXS8kR/MDkQUDCcBl6oRl5+TIbhlypJdZ05YHU562ZVdr
fXhUq/no9RPLlZOHrdB2tjlJ2z/HuUm9dp4WXi+uPIifmeaSOAHijPZtpwHr/H+K
h+GqNV+O0fHJRVIt3TYeHUiRs76tqxEbQEoNOdgGdtsTqXL2UMS6f4E40Bhlmzj8
b2UxUBzOtVd+FBf/yGekY5hzaxjmhF/uGSR/5s3PxktAWzzwQHXYrf9EGGEFR+oC
s70KzcO797hj3IV+wQ9LAXSPjEtp10bfTiOiG+BQOWmzv3he3j8csLckJfj/bdWW
9OM62Yxyg/nIBrHKj6hQrymF6WRSyvD1vp6GsaBRnbMD5edi+YHEKMtroqFcXi4G
9SGbfKBh5YOERYVr8jgjqlcCoW9P6PYJIOb4wvSYJ2HsWeYRZ9CvOZGaQvLOSt0b
bw8098k+4SM2GtGuJe1QGqVeVFoysbZA0ufm2kni4lJf9JnwnRdv5PvqpWE4abux
qr3wsqFNj1CJ8TORkkqVN/lsFNC4AKCQNA4sM8tHEjeAbC5D8FCz421aiIUq20IQ
4zrvWdP0fJd1s4MCtA4ppZSQ0OkxRE36jyiHSMykBUqJiG+YrMW7FYOXg636Jco2
PBP0JvSSa9L4MQlVIq24YKCqW2NaDtkoHC2YqEjqA4K4DED8CvH11FBbIzXe3G/V
Zn/0NujPQg/mbVFkDFL9HdOXd6KzMq13U5KGoFsMKPbf8PBTz/05SDVBF5LeA2ez
C8TC4a0PeH/zfZmDQVTpysHRBur6b6W5d63SaSkj24hwTrFgusaHk39FDCKJNNPn
JMV03YKdbHJJSIdJBjbPI2Xap9n9ZOAbgvpm9Ew8I5UcL1LtnerfCxsjD095fhpZ
PrgRz1CP8+bWUMKISt2axw0VYAELFWrdyhAlyS2sC4Er48Xqoz+eF7Gl559l+ov1
toLwRmrl4j6rb4y5XqHBgx/PAg222+x3w7TCCILP0gDKozXYGk0hHFp3RPNsGfsI
jOaAAb6mt2hJpkXdraTMPzrTvi0OYGUbsEZiKbbwRNI/R7nxV0CtQTBWM/R8VsOc
N7PzgfXMc+Te6e2EnMv4GkRgBuIB6ZCS1Wy1SVwb1hIOMLNKE8CSDuSuisVkSfGU
qFm4/vq3yR372JW/5YSWqFZd7wGQ9YCQ8P57DsZ/Jv0yoVgcYFSpDrKvVweYnx20
Vl6HvBK1j6HBzAB8bulABPJt2srfvlQuxmJTr/u1Ci+DgPlVdUzmj3auL/H4WJ4O
erB7aQndSIn4W/MrRsYZc3wuygBt8FOy2x10fg0HpHcTxKvzOXLGnLUhTm3+HDUu
icYqZZHz+1XGHEki665P941RFcPTBXROplvRVqaxbjNlk4eS/vaan52Bfl0A3cgr
JTSiXWtdVJWK3kx2kGES4KTTMYnjS9pfurb76zjZ2eOAK95FwWoLJH56Nq9WKMoh
WE2wKG4g/W1scXW3QteK094Apdcm0MDywmv+GEABDsYVy7ljCpafxwUonuRw8L8a
dDvVcS6mdqppjoWl7JH0FG1AJRrO+VrdZ2XTumjw5HF3e5edhBMfs8vfn8eiQaFQ
Ot1lOHQSdpxrPpW/bAWmubiwIvkCkTj9USK2l9pvLhWHTbt7QjWvSrBj03IMDnlC
7mkERprAP0EA3VKEFeGaaw7BGk1qF7eC2wIZtqTJwrrYb69Qjz4IjjMJRV8QwwAR
rRijHXfLtPRmGEbYLQSlQDEJobjrbigM23cgclsQfDXRczcEvFC1CpdlW+bMOefv
tf1BX9JEO3eC1RDFdwTqzR46RMQ6Ii1GuyfND795L5QFZYtxLUd0IXyYekztn3uo
1SksvWheIBAM7iD/DDhDXgi9tNzlVN3UMcioVU86qjBINHw6cT9PK7PKHxhv4Kvs
FaXKJarDdbSzpfurDMeLQpgsX/hLS0z4AcoDAXg0J8o4RyZRNyndZ9sRUTr+Znqo
vixyTjxQb75rmvxqqIcA4ld4n8rcjAU0zGg758xuhIF3ms7mMRIb33Dp+NIDmaIH
erhZYQapyH9Y3mPjZSMpLYDCy1dZJHFIpKYti75rsb9tLK2iYLf1TGfCbQolpr1I
k8A48Bco5sC54U6WWc11fp/zWFyR6oO4E9uhMlFDEGwWJa5eYU88aWGTXO2ML67U
uGcICFZmB/7N2AIqmZxcUZZYwZZjiF2kTBD4FqnVB4XOcuTdDgCPHALgV2iQFa/V
PUMY2qSi+MLiTFmxehJCih6qgUPGo5cz66MENS1XGF9XE3u73jhu9Bl1u/sEUnOC
6rzB5lzn/F3pe64YWBIwhzSHWa4Zgqec9tvaKXE9xZQXdVsA489OVHuroMICCSGz
A1ZuhAAXwFIOTYiTHtMy0GPLtyZQRzuSCNnWoCP7zyzvJChl6kBfmfs/YwouVKOM
bhmqu2lO9wTHtkklpPqxuiRBIxpXhV062IgLtc/ieWU+ISqGOFzfvK8ZbQVX2/TQ
6iofY3qONQ7DT9/WolY5vBd1aT9wKnn2k7pQO9z0Edv3v/t6pP7CjqL+5/0l4Azs
bfxHOHe8nMq0IH7t/utAMbiJWQQNPF1tKQhfmA5IiBv+PjaLIhhvnI7PyS1Fg0NR
HQK/BylIiL6tcb/8R0Y9wAMizrSzyWA/zVJNAqUqp8yC65EhJqXItOoIJmfPrHlq
HCWHVciLpUoU3Fel6KVCMptIIpIDZYdqhxB+MGTbmjihLc8KlDbw8+cDa7szVxFA
+bGudYw386vJj3Is4xREJylbBOtz33N9de0ZWJQsLBM0q4uvqZ3qWmG1KtQwGNsz
V0ikwWfzl9p5ajrAnzIuQP+vu2P8AN+JNYvKeR9pO/tHUy8Xxb+NW7IeoT7oGOfz
mK9KQpd28ssKuwdRmoCNNKj2hgn/aLvwIdH6qnBMthPG9NsZrKyMy/rYRTM9NgTb
nV7r45kpxgwqkP4gi+VHgKAtfo6aMt9JmVGm0wAk5sBzpEL1RIOUiJpsNTaYbI0o
QdIzH8ujN8fsPeHpAk11fiRLHr7e18Snnl2LmOuQpkxGOzzZjMAaRp4o6R6bX90z
UlkvS6U26TunK0aOVxjB4Ib6Hiv46yFZ8F9GgwbtjM91b1/J3nAIhf60xAZ2URku
4lay9kqHFGcdQ67wl5S4dOd8SucSZ+SSz9ebnACGM9fiFN9EVEmxEgV29oMZZfE/
jsnBciTvtZ33uDDR0fYIMqZU3m8tu+QngIgmIlvQChtn43xnYw4hLHmIywExPR3t
Y3rTOJYIY0GNNa8vzdadjeCkjOTO7llnDZq4iE3ohEk+3JiNZSp1wMe9xrr9peJO
auPIGzn8DNaj7l0Wa1ehb76hZ+owRv6d2MVXcpxGPxjF1lXZ7vgkZoiKrJ0zoMvE
q6NVOSzLztpsHURgDTRr5ZCa9X2PTBfAD4HjRVt6plz1yng0YCuHWcNXin3L/Tw+
ae6oFljlAAi5fHxnuGRymDQ0buc3mU8R68edfiYdBK/VEeqIuS/VK0ZvvysyBWNb
hY5gTmQ+1+XSFGPS+BcN86XgFO5Itn87Rta+Mwr9X/zpfDk7DOxL3D9JAeWvYQyb
LY8AJ/YpWpMA27DXkWMv5EW9gd68nrjbciIbMk6y3u8YjLNg3YblLJ/hOW+BSB0Y
YqEnXRGFLS529J7z9lSX/I8uHomptc6/TZlbll3G/SuTQpjxqgStiaheXQdHKLxR
hN0+IfGta3xjE1BzqcpE0zFD0EYKXpI06fryo6CwF4N2tAbHdMMivcOaHH/faqQC
vWdvKpu0U7F8C2zMo16JzIq4m2vOfSkUCv4VvlcYk0V+uzLW3TAJ9SZh73AmPFZE
MJUVj5Yx0BoFz9d7W+5v9IUj8/Zt6u6O61wVnfYnwC/CRhcOBlMEBF93DI5i6iGo
wlv0vbjUE6Befu0KYJzGylzp8bLffCbc63JLPXpeks6Tig2TuiBzQQVhZKr5FFQM
T8bSMucmS+mEWy66jKXTTVl/E3YtqZIbWlZuc1vUGKYxUycW/+ex835jK6TaxZBp
8bMhP5hZFfbCASLDbWVOhXkmbBx7ylehgWVicncQ9xE+mu3ODBpKAG6qBJJx5urz
18wYwyIinTsErwkrhNQg+bhndh5D9AebGo3g4VNxvcV/K+5aAsI3WBnMCK6vwiy4
pWcI+pgTP/RDzrdIgfpMBSPu4fcYbxGZxj/4mWEBuzY7CmYzA6TzZWZNUQi1JEsn
82RL5gwFHwqATs4/8UHEf0BD3EUa6uUmXSo3JbzwzvCmO8T0FHHfgKur6pRqkeXa
axrkGkhBan7s1CuLb+/4UlYT9nvJXUBTQx67k0k7Kz3fMgCMG89hSBEl51NzlBF8
1WSyGEMMFCov6pmcnOjfj2RrLs3VT02Cu1JVipL1V/QikypQqJO3hLgWpJBa32jc
pyQWT7RTgAv8GGVja4j9CtOJMSXyEBaxhCRzH5QYic118zsrRd71SkIlj9Xj5aQn
4Xqfb9e7qQb/9+JvOef1cbpUqTzCbkemf9PkoSQ+ImucWgG4/MwNhr+aRnS41pT1
YyFSZtsA7V5An7CBYax5aelQPp3ylffQ5QNfTnQP1NGy0mjyxHAxU0K0sztXGwcn
gXDIVypkGujEGVav7PcS+4J+c4m3zbTGSAeM3qwEIqPS7JPY2TFEJCDYw0yaTPqG
tjLN0n98h8/lX2BHE5saeok8wuzl5npTQPF6iI6aXDUcnSvlq1Uj1b9iWB+7Dp2j
WM0Y2/N3x8NU9xO4skv1bF7nwTZllekaRuzvf9cw7yCNuzqveV8lXBMaZIX6DQ96
uz3ZL8ezCJrlFlI161dJjD4hw8NRHozRmPWhQuOrSNitwVfkFLxJGN8X+QTOjstR
9AyEftmWavBGo5RPMtEzM77UynVwpw7pJ5roD1k6aWwwbQFbIvVPfFdP2WKHvtoR
dtn79iz0+z/uM4tJCRvz8CrLYs1W+kgDX8/vEfPbAOjjqJ+A0u/jXIeMITESuisn
yWjLkj0WyZUynA5neuRD6vullQZ+456uV26DsfdbOq8xlVsYA22LJQfapDUKpxBz
Xrc8DAW6pd1G3D6jSTbHW1uAMv7JPI9rRABtkfpNx5j+M9T5p7OE5Su55BI9G/2O
69Sd4f60GRKcz9aarCVdpKcHB7ojyJ2lQHtSMfRxcUlz3K8nJ0beEcNb0vpQpl6g
dRWYmCk2M+HVpEEtwc9NZk7FbbpLc3MiXxkeeleEzbHxhvJ/8FL946lAz/KILWMh
yzN9jPb7EgJP6rOlPn2qpMORhjA2BPLYhvNzp6w0SPwcuzY1Vo/v+YHS2sXR5BdP
fmoj/tv+7WwRdWCsdjJ4jp4Rqty4RUKP8uFdwyQIuvIaxaIIJ/q2w8VwNLftCkuR
gX97fpB4kLU8kz+69uaWp6u7Wq32sdPE4h2sSOc7+N86I5uQOcQKWb6PJGuF6+LU
7QyCDxwRgPKAOWYhSo8yfM2AATJ/ZdjNNGNt7xMTQAaweyiwb/hYO8Zkvu4FbH8z
IhHVOc5Fsep6TGAAFwok7pAmQIe75eIZ9N0AzW649giU5w8gdpio+tDSc53a7dtg
0bvatW6oL3a+hqo/Yk52tpuWXBiTz05JmtV5qHe3+FYcDRU31cUypipREkeC9cAV
SyT7wTlJEHbnbywUVNa8xIwVVO/qQKWw/hwUF8+jCGlYtrFbqlexyz7uEgDkSjSy
Vb0Z3SYocdadXL/BMRHYI2VMQgOq1Yxt/T2HPcjAooaKXCwwjkLkvg8u4HQGPFzU
JLGTV7Izd0wHd+Ri1s/hpUq5qyFUgPb/Cdun3hRDm6xs9aaaKoyKST9YRgKIrZPn
O6wi6VmmWlHCjLM5F81dYeMT3uu6v9EoMh84OVXAyXSROWKlGogKuqRdDW/fTmFE
xDZbao8t4GlFfWAnjyEPGtZJpulJ0TWIXTcjqDtn3N5L+8+KHKKA6CtbzgxE/pGr
xHO3nTz7O3hWHHTUnyPAJ7xX0qMQueJWG1hTM5B2XDrge3RbwI6KOwoBlFS9t1QM
1edHtaZuDA910WhX6f8Jkbu31ZAsyNuHAfJ3rKLMWNQdJA+17zSMcbn3ZC/EzfPI
qn/O//CKRD+NKxUOGVyujE7GZHolIoClgUtPQuhmAs0I8w2DyQRAVO3Rm/xhDlo9
MSOgrS7/dxIH8eosAU5wbd/CAfukGMi5zNueMMebNYhrhfiLDDADZzhA2/8nm9Q3
/R1cWDFpEv7sn0RB+D8Fvw+BqQ0LvoTdE1i309oc3biPN2P1h8IHui54l2YuL8sk
c9XGPwVOVIRqwBRM7x2+MEkE/RIbbU0DopPC9c6C1aEzreEsF4VFC2RfhXpFh1N1
4E4Hu7//W0Azn729OUbieJvqRbCJvH43T0z7WC2ZXITMNMMXvEMLS6QKEhwgbyBS
Pi+n1pA7H+w7hvxeVPe5klzPlk/3k3NNvcB3/kb5Q+2TqrlOaAbmLTkKG3mF3lZk
x1OEwiUNMBGLp31YHqfr6B+ozpGtuesNsuQMizJKAoDYbD1+G4GW+vxnr5zEw6uk
2NnyCDx+WLD4N3ntD/sCcKk+SRkE6yqvTc8Y8G5GQSyiv0XoPC3+Fru4hoDPFQd4
QYaPFc/JZE/9IgyTT6JmCdNYtY2Q5UiJpEIDJ/lw42zyjGHJqreTPGP24hv1h1MF
jW9qX03QryG8O2yAfpMGppWOkBW1QtNIceddQyaVEAyhEwBrokv2gcYM4vrqZ6XE
J66QPndWAHDeP+lRCWIYWuGtJ7ROBOJflk5fSx5Gvqi//dIEW9wNewaYIgIfemS+
ir56RDH5ysRvyD/T9dimp1RFr5j8gp9GTkpy88hcL6kOWpu2du1Dhp/djhjniQe0
mocat0Y1QscuPh/njLAqr1XTpImA0gl3xNR6dJD7vh8GCKqa6/OX/NTas5ttphhA
r7cAQqUGJuCJQ8RL3NejLMVZbGsI+PgTjbW3WA9loKDYIKR6YHCoPQXuPZYozEIy
hyRTCfPbsYx6EALfsytdOHkPpU52ADODIDqrAMoqAVAA+17pG5piXcLMU7FqF2lu
kW2fQUOPQ06Zvp1lOoF7KzcAeQCKLDHNuFvEQiPKQZZDjc79wCnR0uDdmv1Br9t3
XJeRW8bnw7BubImSNtk29vCftHfxg8XSl0IbiN65/Gi+ozsfXQczFj0KfCcMR1Mn
IduU4in+AFYLddpF8fRDnmwpOTb6mLldXJCW6HmJNazQK+NYjGD89FvPjVV3+IS7
PC526tr7phpTXEbcG1FnMkoHxYKWSdscV7ZJ9rmCoGdxwl8T4Fr+kabzhb+VaXQb
t9+UdVtdtJlHtaii7jmTJ9jdOxX+WsypCtuBiMuQV6xMxeCb/GBCxGGQdvfWaPep
ElJEpf0gKlopsJdbb+ANugH4pMK9EevqRS55Esr145andVasvjHsM/7Qrih6R/Up
p2qw5Kbj26TEmQuC69F6HwwYkUEIEu2QRL77p22Tih0zXFIicf4S2Qcatu7zKlOV
YhD1TjS1OyBHsbegW5iB6OUeSOSEDhtDDl5LlEPSkQu67h5j+n3T95NiIoVwU4JM
BGiq1C2u+Dwt/aeGH4Pgk/MBQmpoFtCi0yjWWKzhmPggr6UMq/tBNaxF08UjgRzP
S+dbtkHGkmEl/Kf5V6WmHf8aeZQ8gcXn5inSasPo5AMlrkMSE6P0mU138r681ABD
gEEpnfK+W6U8XzWwtnwhB1R8U4nPypPN+Snse4XOiBOuiML6ufhOLUG8VsCgLViG
bCKSkE+AqZUCE93NXwlaDQdB2ChG/VK0/jBmnEHOKcBCTdhv8jZ79HHf4PpGNg+E
care4dqGWiw0VEY44lSuXsDQ6bel2DsdKyuPAXCw1KJdaXk0TFBJTO3GfVPdOqxx
m14E4bbl4Qt8yg1xX7Clb8BS7d8vr0nQZRWHR1s8dfO7V6ZlLE6d1LmTN1e8I4Dy
CfXJkZzPgva5najZPecaAJiK4UbaPwEwr45qt4NbXY1etvZtb9yuHWVagp4Cyv6y
PYrzkrN6zbWXB5Y3vY8pGv6m9To8j92JqSCphAunbwRQrS6u7/OcY99WLHooQIeJ
Gh7CTomcp0d+5S0Zgn4Dtkw1LLAJ2UgcBIjwMWOkB90oDR2eVYUpaDiysqvzyitW
rOjO74EoB0Dy8qKr+gD6hRgyIbCJgZEfigXPP+IT7Di8LmJNRPxltfVJsuVA12HM
YJqtakv+kKRjp+ilGoyUlseCZH0I/PSeyvQR9wSBFCyqOGl49QDOIQ90Uq0yFgvk
zkDmgXfoHIhI4cfsuYeDzvwlUMymu5rhVMQux1YPsooEnVYs2qcLSdwAFO+C0f64
mEGJ2I+sc5/v5U+/ECuUQKsdz4ronqnnr1Q2Lt2E42e7wr31OERsfqvF+kikO7lC
uqr4Minxha/+pWL78cIHefRsz6xjvMI6/7XgP/aFQOEpRAag16sXpK8bMm+6uMA2
ZhwK9pM1qNL/6kmf77jae3LVjutFHtzzLSsKf/pb+XzyjakGx5ZWtOtohAGbfVc/
+WbAbWish09h772J7Tls5x7yl8DHC+KdkrcBJqkFaKNRds8h8y8tr5bKkkMr15aS
StcMW3usirGbcHx50IKTrHI/klYtHIvvXqW2H3ykp+xx5DkDG3hDV2dJ88RoJ8z9
4ADHXPxLc0noNcNG5UAfGdcmdsgEbNcul36jr7DiyZdmaCFo9FXASAtRqyWhA8WA
27bY0h+tVkWvPLaUE5quh0+DnPzRYqxbVCizMI2/UVqdWRXiQYhN1pWRcwDDevcd
tLSL0F3Q1BfmNrFrSIghJG0kyLK1zkrhh6kWRQ+XrriTANEnt1M3dIZIVvx2y9oS
lAbKNPrtZex44lGzu8LoMVKTrt1amecTZ0i8Xw2F0LcnwtZ1g5nKxHr2+vYgvCCh
5zns1DqQ7IULfBSE5RJq3a7CCj5fdz7tu2PFtogRIyNq+ozc9ic+YNQkWsGtWFrw
sFeMCMIHLGL6+ZV/hHxQb2OhQuSjVuVIzyv5S38zmZOpMPXbAd11jrQR1KQ0/xEN
4Zt3YLMEawi5BE4NTvjdQ3nfTxZzA5NlRMCfjBY71JHa5hFIArko7WB3Oh3Vt0RJ
u4ALNSdgKEokde9AZ7eNjcLQo/4DrN0ZYueIGY++BDDiHZfOb2FRuc9zOSJ9VHBX
szOpjsCnj4KP58Cc15dL9mvqT3wDogF/jpwnW6wN9NBg5gcXlc3aCZsH0mKaPjyb
3j+3lFeIw3s2sS5LLL51oKfzSKIxYX1cBRRsraA7ah/AB69lTqI53pyz23NfNMQa
n6tazp+BmHLYWflOoqxX41ZKFzOFjBHuHGhkX/UNak+eT55GOT+pDdoiQ1TJlCvO
ar1AHfOfECVMNCyzZL3TMJUP9VWkRhkIfJILbJ5l+CxSz84PeLQwOOq8v/CM9Zdb
sswXewrPbDv8+K/dk3VuArma2hs7jJfyv7v+4lHjMUWO0mUx1f3RVGy4UahGEbA8
YKNQQHk5pnNTMP2FMhhrzcxdY7dis8rEUAV57U9+psCpV6UajP/yUQc3l7aJ4hZJ
bbdhGVruBOjdM6uZEUQJ8ZMLvX6E/Ng/A34pVIuYNeQWm0EfLBOxDT8VbgiX+5P2
gV14+tWOsmPhqJNT37hDwsnFAQ5jmuG6X8cCvBVPoh/prCgho19eroVolj6Ys1fZ
pT21zWePuaMK4B0DnYGPSDb3F8ABUhoUe8PurAEN/qx7jAR4sVMN7Dz47BpGNoEA
/eqi4+Eu5dHpKYfsunVM4c5eUu+W9U/JTYBzrnRkY+U2W6e6CRM+ZMWlCRayKRLC
GpippC78qp2JNyUCWS9+tTMqBtUAS3ipb6+SZwEv9jZnFkFzCIhViZzRlp7u9459
bKaeIfsNmDD6A1qtAilRMsihUjR/75vYGydGECajBlxQ4qTiB7OPmhfkuEjPY0kZ
hNZmQIg3kavh7SAl7W084J/HZo0za1M/dAq8g2gLVrVmo0EWcVFNjjtbj2HnVtTG
dWoBpQXpkPHMlR051V9hKJWotsXZZUvWuGnzveGhmCYnFZ39VpdRC3QFGj9ZtBWQ
TRdgptnWTMP5gwyNSWrxU1YnMd584A1MHkKmR7s1kd1icoErn0VhDn6sRgM4jjDC
6JwvxNHKhkTLcnCQQr9jZbtorb/wqNCfG7FA46ijcdFKdiqPrqkfWqaA0gjp2JDY
y3b+m+GeYA8MDG4GZijejZBTNa3gg/a04wl93Ge8/IxTl/H6lwfb612bKGs8EnI0
tOPTxFWn4luXfXgpWRIu3nk0lowMVIAVktsI7Op4NFgj6Id9GuP5wx+4uHSvqrOu
/vD7kW4aCzqGKENuccImgjY+HE3NRPJrB0JHyhKS8O+P0hCS6AY7g0tkyeiyRzo8
pjvlJP+Ftk/pQKy2SwENBsI4mXGobwGCEVQ4ShwGc3RfgGu0tNpFqal/IRTNvgNA
l0oKjxdCgjU+tqLNkWY4bO2Lp5bAT9mn1YF+Igj1ZCoylYWx39GQTXlk4b3KxlOZ
pxLlB3QXSl5NLb2D8j0yhsmVUoKuVpaKDy18kANnk7s68xze4NVrYUo5qdmY+uDN
FBy1NRCEAldNCGat5pjq8HefWChRZVOXGI6jD0lMFsvTpobHIu+qGhoLZ2gam0WI
dC2Ghc8kBL2UtcSQ98RUEzsCagaEjlFcoUw0gfjDuxStfXeV4KfaQomXbwar5ub8
5eimxUvuI8l2RLhrF1NWOGh05uLUTm5+J/oTQVi5YEw/iy1H4CLYE6A4Ablk3M3J
XpQao8TRbhepGn6EBHptoLRLZyosRrcI0HBRsCQcPdRBdIB5xlLEWG+Rx2d9131i
t4Bv1l8favpeoPjGYUE2Oh2Er98w6EazL/OVKmnM0k35Xodc3RLJbQ3I41aAar87
jk2oIcmtqcrKRhlZHgd4AlHTVTeG4na5FbfhUG60bH6jX6oxU0fF/2Sx1G5/vt76
Fr08JoXhB/xHymgbXHdau706wnjboL5rejonami/p6dCZ7dVh3O8DIsM4LVKVNLr
q3tCfXKmtHggqCD1kCalwxeCBxKUAfiePErNHvt+Kf4+LGMSihHt5LKH5mQZOR8Q
LUtcTI8xjvTgJSVZnItueXfezAtAjTSP3dot52LgCOcHL3sUETsNBo8IK0M4C6AY
fGn2oErvZ/zFzYaLwzMuXwjzRLCGwH6s443eu1eO84aY0PTrRX9Ap7DggyqM6pBv
KWmw2Ogj3J7CptrSNlI+Y/xPtOoFACffDHZlT/cvJ3EVNYyZkeRlhevyU1VXOosN
d5wXgXVhILd8LEHJXEznaAioKxp8Xa6ayp0lx9rOLkpqvho0Jw3sm03kkbEiPURX
EbNrBmuPWrerdpoxsppQgJ4T/c1bNLRp1nSR8tkwM+cPXYWMtasq3cY10KVVKnMv
CUDpclsSeopxRvXeHlBGTb0N9FZtGvNw03PLK90uM1ul01F1jfc5giSK77fk4I4s
JqFECLdUAlkRaWxnozvwfihua6ikjuNYkR9QRZiT322mpMBhLyFe623RYh9YUTgE
W5cwaQ8i2S4WG8IxlbnsDMlHJqh3Ub+05LMzWc2JjFBtYBKX8lx+f4LiL+ArHN2J
KndDeKprjtcv4rVwrwxHHuNiT5h6VbZe35UFx8iVq6K6QSsJAq9L5wtWmLMIKhXN
IfYArfqfDV8oJu+EDgCfMbTOldXP2KNdcyr4lnYOxpFTyj36gSdco4dmzEYianJF
tAfXphFt1Wnoywq7E8dkLxiYzgA602YNjJSCGZOAyZ0NKLBx2RDEDYhcakZkS7mJ
097U+Hp8IXXjrDRJGugKVZiGuIPoX/I7VQKJpglrhCluuOQq7b/n11X9wY+S87Dn
FrNXAWfgRzE6FRwn8+aBxo8dx+ziGmVGk9XUzSMn6hNS+42JsAczD5eYKEBeZBG+
P25FsDEuwj5c4NEIrD1rxTV/8yAPzFv5iVRtyyDhj/2zopnBjqSWnYBeftdaP1yp
ykrhV7ZKX9CxCEGfu+OgJ/2HTUEP4tmta/kL+uWVZ0SYmiXmSt+wtiZZTOoQfRgM
c56H4xAlY519Nimv/pkhz7Kv2sUD5JlMfb29k+a+cUQxvlk0cTeSir9MLhYE6si1
NYmFswLXxdPFor3+zqm1igtYPSJDiTg407kHqgPSB+cG8SBnmoNzY1VVtpzrcmqw
lxrAwBNzMuNFOIy7lkbRBk6e1FZIlC4LXJjMMl/cstwkbxgaht2zASDYxYNhKSwz
QT+Ouy/1FvmFw5LIJjwbg8dQVXmPoTYiGdW3wnnIxJfmAHbquwGXptJ4Oi91SolM
PUW7AIPdthq6q/M1+oNAFRbmNMr7u7f2Y9HcLFAp7YRunLvpBAgoG7Q+/Etd7bk9
wGBKlCqpluY4luH04eedA2PyBpT/pl7fGVnvOTwjr/9QupNi0qfNfXTPnzm76r5G
H+r/t/lnmAGez4FPdfvhy3pYCxMQB65DLVUeM8Rgz+d2towo3g3RINIPrrU/VRa4
XrLlCtmyv0Jo/dGAeeeraX80dp68LfBRXxkOPL/c4WHB+QwvvmA+NGNdh1Fi7M8J
kjssmPF/Yw3b+CGovy2e/35StovzQp5sCuPSFsP8e/jWX0RbUj7/J0OsrqfouzFj
tXc4eM3i8BZXNcSb5xCZJW+EUIIcKz7XStq6FnQzYrFtDf7BRC+C/skMdo7J4Dr9
ab+EtxpdWaXaD5zgQmdmviqahnBcPCXKZCDbYZITzjr8a8gvLtFlZy3CHeqPheH2
ibUbMcMbiyj9y+1rONGHGD7PfRDOloa6LY4LJ1ei6VkbQDQHjS3y/uJkDio7TyAt
b1Bo36GQNKJS4jw51ZzCQZb87ifv1E4GwgB2OCzUY+96n5XmtQfebBoRXIUPs01/
pvNkU2ZGie4r2vwTzbAmnnuI69m7fP/XVp8r0cEEV0WAAbvvePkze1Y0UNsmHk+c
YR4K3o9+R+Vr5pjhq7D4Ckj3Ipxseq7Q5IvebbcYz4aeLh64KTnHFK98+7XSrn8v
a4jujQPN4nEky0Y5RyJ78WDSGhK8/nZd7MzFOGoWpnunF5lCM5ibm3YOntovEfJ3
tOoR2p9L7Du9+/pQn5TCSeckeDjfAh+LhP8jTO7AE7uog+ArXF66gDF1JvrTpww+
mVphzH9phO2NhaHrD4oqrpRWgeerjsC9+z0sCVMrXIML0eKU+57nNqowYL34YcMj
SSttYVjfVSMv7pmhyFlzqpCrhHE9qLgMawt88NTdeiNWfoQCcCDbPLn2ePmHP4S2
KBGGiQIAexansZ+8+TdnmI2fkkaDMDVwsvLd2ksELM6newbPdZy20eceoGfwa8pv
g1h1VfAz4OXOsquHWG6LndV+kOQKLtxP/Vt9d/+vHqdx2BUMXmpRWPKjWApSbww5
W9g/SHaNBCe0FqIM5M5pA6+K4H9VE13B1VXmlnIpN27dAdczCPz3ogTT0Au9y8HR
AiekfRxmEJrLqaAkx3MzVZO/wSKBXHveOwYEXNZs7T1w7w/5U5kC7m2+x35+HmsR
bGjiAquOlPs51shu7Udfe7+6vciJ0XcEltIE7NLn0q8UVx8E93ZgONRZGuODL7Pt
rGFIqiwfeoOvIHV1nBzcwcGG2pwQycCeBzpc5gcndBUT3wiQFqKTXgXiIojhS/3N
b+IFHLOIdcuML1Cgc9COX2S3uC81NAv3KRuneWe2M5itMYSaQgg2jLDcOMfT+uqk
mAVPTbCetrMVOU1+FLJDJY+sfy1TQJZjUyMJx78JlSmX1BffLu7+sLVWI9c/MLmv
sgP37gfuGHg1jV/KCOw3uhRksaAZ59XiRSb9UeQyHgrzeYfoWCXyQGxyH/TXF4VW
tVDcjX0px1j7r/5/J05vc9yC6p3nxc1pGH1A90CA9tjYSgp78JYwCdtU4XRAlQBu
jB4Q00T4kGs7aOo0oXSFOrkBINoEpWyQU7j+Pcfm99vMlmj15PUdXNQ6MRsISxU/
7espS37yFSYh5s1UVzfyP48eIrrZCJXryBu7cFkN5eJWUQHeyCwDHCoSZ4dLEE2S
efzFlFbGjoSPBGJtbL3xx9hrsNczZJcYvnEd9qnPcjlHK2eBFVc6/9x/quaB5EUc
NraWkdAl2LxBzz8pGr1tvRwm/s77Xaiaanky9FYhJmqb0sA3VLI2oR0Mhc3c4CsB
IURDOECR+93IsmlA4yjnYvbSfqo4m5lB2Py2HUqr14VilfXW12ZYRd9FHQlh4Cg8
8F3c32zTrkwNr21mcxmlhbotGoMAjuId50s9Aew64ljhEuWNcHUaKt9JXFbmV1YT
5WCDXaMluZlrkJs09EWUiXCl9UGhk51bFCFR3tpnMm4cCQN5K5o0lL86LxCXXwBK
lgj6NQB3+s0noFOWsaBQWyMwkWx/aN4GLFRv6CkNUi08xQ7+KuiwL3LnO6EFvCrJ
BX4lbJzYBehuifqzO8JD9aRJ9237YmqimiLMLs30Vu3N16MWJgqXr3hflIZ1Mq2y
vVXocLqcQ0+m88GUGtfpUMF3oixuvLD8DQuFewx2fRStknJXiw4e1KxzkDhCzCPN
iVYqdyZGksfahGsWv1+OzMY/9X0n7rdZskosUb74DmrA/qc+sRYkq2c19MdgbeRy
UU2IRH+BFMUMp6/KcKwsYv1g5JJEAFc/UTEVL4TS93T75hVvHomiz0h+OuxIr6qM
nRzZXGj/kTmcyIEbQXvMMpHo7sUolVPVXKvxKdyeWBvtVw6Hj7T8GJ8vcOfKh3Jf
5NIexE0sae07hHGjhOL6SsLa/oH9uv5tX+u+R89Vz2YdseRVduNvIQP0/FJFNSde
MS1sx2qSdQWnwPjDx88N5WgJdYV8UpXKI8g8sO8XLDD2zcl9sX7jtjl+MQi/LmrF
KmRjhpx4S7BF4M6pXek1nRTB39DZQ93hYkF3myYHFwCvDfhxiSMH7uhOJbW+ZcsO
v0wto99FDYxmor0a9iDunWqhjvcDnE7r0Z0PqwTpsoLOaY39IxQZ2VGzZ4xy13N+
LcsICln7b2i0eMUviw0MrlcDhA+BSmD1QptP3w8xe3HrlFZHds9kG8LlrW6tJloU
DvORP+lBKGLosPqKoEpgOksFEubO1nENvL1QFSTsE21fZDwFncwNyrpDxcMQJeJ6
B7v5FfpNYBXwTLvp4Lsta1lyM/YvM6jHQJqyOPTIkBwtFFXrvJSohClYluOVQ/+k
LM1w2co4byvuM3yd84ksm/ENjZc4qDfkjANLSY7UmRLyCYFk6s+4LDecrJmG3vLi
d6C2wpfpRB/Bqf6zNQtLIU4qrAU3eSer8Mo0RTq66hda0GmfVUh1wi83TjOBmETi
1cqL4kvaeIAJzH8SfUZvCNjmf6ryTgQGk43qzCdBI1h9lMcAzKlVjcl+BkJwEVsV
z+GIf7CAc6g+fq2dm8SDxIIdd/qE8Cqd0nmNxxZb5irxPwBhVVLpx6VXTbDsvjBj
RNCc7jBQlsSvo9wf1S05ayWDuuYvPyDKFSsh7Cm7FJlb6gXZO6igE8KprmgJau0X
5HvT5mvp6CLQOnVDjJVlZfviYJBkUDzAjm5qUQD/XNEge0jEph6KJxYwbDQsHEht
8D///gOWLAMtNqsmZ/zwIykBX7T0jcney4kZaLRZ0DAhjCUqkgMhfefb+TRN/Xkg
vzvJI6idX7BcsYokqVE+Ff1xR5P54Y7rfkceL8F1NvSMUCvAOCbLVXjP1kXI7xpJ
xK5GCN+4yZ+oDjIVgElLYbMNIQ9k3SwItJKqfJcrE6kPZvi6ICuF/7ZyduUKTbht
09xJ2LSNrXL8PUYie/GgR6XeXT1X6i1NfzzB8cXMAv91FRrvJFCgXw9ybNXX49PH
1OvgnqBTbrYkjdgMQKWeddA8RT6vsr6wiYrthsmkLI3VEvr+imukPqt4/0tdXmzb
o4mUYntJsMtK5KXESX3VXdicf4c6MeG+uyzHsCsgUvHieEyhLY0LSBIL1hzEXHrI
FV1e402J7OgvN1PC4BP8e9kzQ2RHK4aMqNqiMoVOzw6cpSMfOF+V1CyDmfdebx7q
CaKtr99UpTMRjwot5nhJXci8dXz7jYCvyAJQu0q28o6jz541DAH9rL3FrQwm1yMT
LMjMJmqrFffeAw/jHjLZrfDhEhEqqIPM9gvQgyfjYbfCd13zGFQ/w+onH3R3tOBu
sGJjoPzmeC4tGYHqYE/iytwCpftWVemjnPqhxLiebb+GY/mSn6MCIkrd4mYhdj0p
Ee2vtCVNcs56WkdQi0Lv1HnMUbN3aMxMx4l/ML1cFJtqgTD6zrN+ImrFjwtVE5tV
lbyOIZAVZGKm+wITRyywZ/t7iDu5ptiaIVRvLvGQ9TKM55TnqDqARv84kFWueLHu
9efSedHkOc5FzxWuS81Am+CC1JEoCpRvsErSNM062Tj6I299Jx6Axs/vWqbDZuF0
+gEUcQzUKepWVYl+TTS+AUabDGDt2s6m65YMEIWS5yDhy8wz7y5Iw/DmTojPz1kn
AjaQqIfxZvrAyh3aHBtLOwySUQ9fZpLQAVrvMHMXsYX0M1q/ZWLSZqj00P9VUSY/
YhHy9Z/Zhwj4vXuDJ6WINP7Zqq/KgeoOxQ3LNrbTGjjnEfrK96BbVRDsyDhfr3d2
lqyCNvDWHgEGAxU4q4iDLthV9avP7LzuKP+hvASaIoEo7n3NRoR7g8vFg6pr/WFM
EIyndYDXajEU4inS/hO67Z1yTXVk+l3t+PmmX25aipqr1dVVVUaGT1kWq+HDhHKL
yjnhDSftDEdUyE2yXcAZ6fNLczepAYIeIIW/KYDLm0MiOQSadXOFGzh3II07v0Kd
Oy60m03W8FoRkbt7OXZJov9KoORPdAJgKJKc0T0eogmFUQemLjIKaXXR7tn+zl2X
rJfcpW6aPwBi1yGAzmdLeii5TjufvyhmmSefszwduIeemRXZEBB48AOB6X9CXJZ+
HZ7by2jAom29UN5tw04pQgCK7xu+Nre1sG/nEdci1YVFJi0d1y1H2eV2mD6cc6Xy
NxX/EjDwrQ5nsmh9jj74VXzsL8980nMu/7xPOUTvkaTs109QWrTgIxLAcDIMZ5C+
LcNqwnbbRdsKHMJE/kiYkqgN27aa8C8ALr+Q9SIlny73M/zdbpcStJQoVogNZXDJ
UIQ5ItDjDa3hvAbwwydjgEdFw9TGQiA41kUqS6UucYniz4/c3cWcTfhbYg1Ch7Ba
bqxJtnYV7o/IFRFO7TXV/Snig1NtECD+YWiV6Gliid5Wiwm2ZJL4AZZVkahj+rXj
oMtA3lwmp7nJU38vuLWswUlxLr/o6PlNRrBh4yeyy9FKOlWQNwm2EWhdd4HLP3gl
DeqBhp6SzYcTsjhk2Qhaqs8dq5Sp59ETJDVrZpLnfNJki2Me0zrZuLnJyljFEPkK
rkfYaY8S/Rg0HYztSsDFZ8uyQYPbi1oyLDz2szsSUUMos8Jxv0/zlRpR6eewCGUQ
BRsbEmeReZrCu5DofqCcG984koTLNQl7pMcYlCozPz3y6i1eeoz47N/RR2kYB0uE
hdJPToGSPLT/XlEisQ+IYPy8qKGvuvTgl16zPYktiei6o6HY+e1yK8xWw+IvSOZj
rtM3pa7TOT3coBC3N0AQRVM+9NAzvpZ1J6PXKPhIQiZCrdFlrtWZLz2fDiIHmboJ
z+59KOQe6LZhLh/muAu/tltI1M5/BqfFP92AnxQ6boF9bSgP9VUefj8yGwsj/n8w
k5QmPixgRXKZOqhPFAXQ/DrRhQxaotcSntm4+Z/DAgKu9hjTkyd6Wmzm43q8Toz6
Ubk6PYrrVGKy1fAgl+5DReYSzjU1JlWFRKun2QMUdjP0bwFKe/XyZAIFXplFInOP
Vk97ScvD3jl3lL2s0wLGQLiLJWUTEx1Z/oIa5QCqkY61g5c+Wc85pN6Iz0uTNnvB
ZEx3vv1x0uzGSk20Z9rdDAh0QqX7wBluggVysD4s64z89ozQt3M/ZfEX+FG1zpHY
frIPieEdg89OkOhuyIJQNAZYnmccmGHe5EsLufPI1G8y+8ZQrZzn1DJYaK0jWqr9
zTevI0MOYMtRPqvCDdkN1iX8JKn+NsbkrsKF66kQc5JRG4vzN5oM4HJHZQ4y8UFe
tQbmrz1NTG0GpGnWfb0oeydiDjHrtmVFMee6I2CoFqdRD7+vybeXXgsWizP5vynV
Xu538RYQ6zf/OYHlHQ82tmfJRiAIXauo78bRSJfMoek3kLhJ1T2WWsaW31eDxbfZ
STGC5YwMHT4T+rvVDaGyT5P9F7yuJeuMPNC/oAUiBcjHw17j42OnJgdxkkCStTUQ
RH78LQTJWzDz93DxjYk6cLcdhhbwDe/LD3eVPQ8bFvJGbM796mePRVeTYWLJaoCI
dQ/I6k+D+z8xyxbmlXITYRJwi/AhKoq4FpV/puSaUXU/lhU8+rZCnTrHgSTYlXzy
eCMUdWvxWF8BNPSYyYCvsuZzkAyta0QJ97YT5ehJGXPYh9KtEidIn8CW60LJsYEh
3NCQaP7BllGBGKQVIl3KIuSZrMogRZitcq+J9bcVc5I0n8gdxm1wuvin5FYf9aur
9a2v0Qspc4yT3TJclF1DQMuqfCRBcIusFQ5eCRHt+t+EHCRdHh/EkAD77mg2C25D
BXVJKlmAc9K4b+QPrLKROY2TzLX+TWxNYkO387L6z1yPr0bFbN5vWErUttU+0GIe
Tcp+7lP2Xrg6oWZ4juwHupH1yqqmTMeHjSI/ipn3CzL0SQYOhnY/IzYzRZPJvD2S
WtLCE3TyKZzSt7559Zg8K3NWLctnh7E+Bpk+NeGvf69X+Xkc12PqrqmxcqySUy7H
0y2nnsuP5zkU4WQdwVwl99dwQYRdu6iYz3GnGPPKolexovSxC1B292QFchAvdzbn
ZEBKQGUxhwu8MUD/+IMxb4Dhj1OrAJiztXA0DH6XOKAIZS9Nowtyw9htcjQ9+SE4
btRwhfSCRzqAw2/hehGmr0aYZ9XoNyhK7XbX8NrEKwQSNeaFPK5xlj6/zvKQerkA
UxuXenXBqZtG4cRSj+ERVQr8exldQ4SVfV9V4BdhySwOBkRhAfXLSIhwRa7HBUea
l/laXoPvKTNSrQlCDdsLh9GTWEIqnssGlJ/IfPPUUL59Cg+G2jmAT2a3gNvmsN7U
xNdMZ0PIYGiyBeo51UkhPyj0VsDrc5iORLa0oBAj5CmDx2mrFI5fK4LPxsWabrio
ldF9ORdx4uxGUcUjkTivn8L2wEr72QJqHtKCpL9h9ZK90diBoE/gdFyNI1R6ixsZ
dxglfZCdINnWtsot4FQYA1qMoXPAk8t5tD8ln5hDqpHq2nf8MLJ6mQMv1dWRk2Ph
shnmqRyWMrCNKlhZWcGqgvFeHfKb8mYLRTz3PFZ110txihJAYR2x/C3Fcph/74e/
TVTsXlMAHrUipKfDtXXudzqnRU9vHDnlXdJ0Cumu1xnSxAENeTTDHteC9yEsVU8k
CFg1lWg3H62XnnYqvA4KETGl3wp3qIemgV4TWijntNdSzx6mMDEucGPx4ifABW2b
xH5kJgan/OcG/vZv0SIvh1WY/GsaZQrnHfF5Y46Zoa8CdKv0sDx/7NnI+f+QGM1g
IAhW95JqFpb30LYLMbAsmmwTY2c1GgUMAWmrJj7UAlmOFtWTqUhzWSH7RdcA+y7p
xSe2RmQRXNWxd/u/agUexruvZkG+j+QGmfx4vNyo0J+ElihxhDZdSR8S66wKMoBM
6eCQhxv2/buira/AEqVZw9kCkfTQ6kxPqj11qhki7pYZY2yZ5xS9Cl5ZUBx8VI6C
tOtdZA0oP1M0qoj20wJRaMrhhbR9CogIDQXg8raSmJSv8Mz+Jqfc5r4BNoBLC/jx
KwMI7ju4bFore2aVl2h2YohYipLFJhaFasfpg4A2ZE+cYmHN7GGYVBzKhVjmPIpp
Xn7iqT9fnwfl1nWZZMBygyCQQCT5EWT7Y72BFLowJRTzk3wkFylco9SiX1we8OdX
cKl/atImxBa8rbQz1zuoeZw9+BHyNgqJfgQw8vb+E+V1v90AsWVdcepGLyHHq9FA
OLmiFsqKkFtngOOxLlaz9XQyz3WwIYDe8CPeBlzzCEzLBAOlnMI7dHpcCOJs2OI5
dPyUwhCWPEB7p5g6FIlFoIr9XaLl5qXWlJqiR+OM52cLf92g8XWA5MOo4QnS4rkM
EGNTFrf40thlR8hL3v3nh8kadqqVNK684+AUEtHTH4YSFpekAcPPlyF+v5iN5Hgb
eCMoPZRPXoY3NfB+1BAAMSHHBA4GPOevCvBXljyCzuV5y2W4B1dImPtbfQjKLqL7
1A2yPyToz0RMwfhcbqtzjjVnZm17sJjtIJnLHAzviHNCIwQiqqcL/OtPpN0QcEOU
sw4JhZi2i4Rm7JwkzAusOd/Nmw7F5wFTMjlQQ/Z9JdqOw9V7sWeLknQ4Qj4GNL6L
u5SoSSg+t1CFRTRAqi2ic90INAaL/RzJwcOeq2k3XV9kHyUQvMavTd5W4DXnKiZQ
SptHrkcsyEc7sLYi9p+04HAa6zMCTN0FPR5O/96QqQBVd2POYeqSN0jDAHg9h1IP
rgHRswzRzQ/fHhbPZEEvzmWbicBHnUgdkFCzpzkzczQYYL7bPnxupM65Wj7PoW2F
l+mApJpsqlfi1cRSVcgmoFMIfWishPjVmxAGdfK/O/GLyn2kp+1Dkhl99fb8E9TR
9KsDSuCkW2iS29qgZYnGSp/OjmfTCOFD/ZiydVg4buJOeamFEe7XxWN9I50g/SlZ
BqI8ifM2Lj1/knNbTb8tMxHxnz6MjUOg2Fnk1f7qI7zB6hJ1cRjzLZL+A2ShYOHJ
tn7ebjxPDTar7LdsSj5DKAFWuWB+jVGXciRlhsvz7z7mchjRHXkqxAApzYH3Y+4y
nlVezjFJoc+QZZNiD7sYEUlzBBIkzFFj0cwG5sftcsBKax4oBPxwdBIOTjSthcN7
AuQZhUy/kdxpfa0xe2k9uNrwfcnTfXcxX6Ia6mXgJ58FlT5lKcKxZAs013Hf3FjX
XZpjAfmk/QBL3PQMqcaPtfT24U1PF0RJyoosAly7mD11rve1gAdbvqA8kb5qj8S1
yiERJY/v8ADCZ0jg7ZyXkiZBLqvXR0Iyw4d+brviTCc9plo6m8lAgiiPXHNS4fjo
sAaFcGgpzxqKIEA85D4wgA5mRRc/n7flcNoPmkkY1RXi7U+d7Hex18d6GE6HaAe3
q20KQSP0nf2eWgRUpOAed4Th6muBGkgKAKPBGwFYE0nHW70oXp7BLt2Jlaj4Zboc
dDUJny2rltzj66JXQqMmfcKZC+vh4Hy2FKlXxgP4Sul5o7v3CCAQyf3mZaa4jUIy
31xYB3sKHNQkiKi15v9nVjxgAL1BBWxhAISI8ASIB6W2TLOmceYMUvNqqPNJ4x6x
OnJBCcEnWx5hwnqCoPcJO0mxq4VMXal4YSfOzZbbIE4HTb0zjndJiqmuAxF+/otH
ngvqAaCck/1YjQdj2v/V99p/kiNY4BXAqy0jQVfDqK1vzl7kEWPsX2JL9vztnl8p
bmB5BdV7DtgUi9vTs1kA3xCH+xGP67HU03d1S8CcgOtPMoOE4jB4nOwkPNSKHIoe
LcVqHS1tBOKk9B006G03UZU8BjZBdu7gIEOZ+U/AipLq+D92zRAUufGLWr1nSKWR
vMoFI7/sCc8sp9RM3k8KAz7R9mgtkGvQeNBBONI+nProk1pof+PWtDimwqsvur8B
TYWQHl/E/KD6Q+AuNKa+ykFY6l3XR8NpvGP5l18MY7CLUAGQDs9+QnbMH1PqWjMD
E/f+HwBS6nOs4OgWHWcq99CXIM2pHI3oUeCuTU8IH64hnagoGts5/+UUMStg0kQ9
WGsPhjvujwFMSKNBzrjowhV2PFrAmb5Zgm5dGgTCnmqUv4vNgiBl+xpyUjyrpt2R
735lVvUqyCWmRehA0RjZlVvfF17l64p/7ofaVxkJZymRKh1uyQncbcBaOngUGmtA
D3Q8qnW9dF1Wszs8Tc1O86mbdFILf1xZW0yTudPYyyEyZNp764NCYLPbDWoeC3sg
YHeEl++WVvqYIaoinx3Yuz9RlvDONxp7GDbqQVcdWawc5UoOf9WBip/0vQIpt0to
MvGxQpE3joD/3kYQEZcBmSsdv+70yxUGv1OGFaZrAX2LZhj/q5Mw/H1h1ArVtyv6
Tx6i6879PkNjq0grMTihPlCqKP4cxATyNvoTnY9gns0jvt0GvwVbm3Xs7c2gRcpV
qozrv62EgUxketaAK7oBYrWzhqWrwvX4ibj5cxiq+xYxGX+bbfCTseE+YsO099aF
9vhBiZXEywR0lCpUjKUXCIwOT15ZocH/pfh+TJOs/9UA9vwDL/PCtmgav5JQWCcS
a12HyYjoXeR56cwi4A8urKZuLnqsGxBmDfFDViVE2i/7384mUAV+vlJs5KoVrYAR
Q5Syg2hGmrcVLeF8eoDALAbm5YfX2iXk/hJcZcMpkhMyPWIp5IOBcVPDEmC0mUvp
26UWuwzOv4ZnXImeVR8CSQZKFc2ggE1ZE2KGZhstEI6GR/VrW6GF/2sR59n4nFrL
nyoC8AsPEWx2d6UCnb1ooefrK4vjb1P/fMl8cjGc41ukl+26iOrO5RXLMHb3eqvw
IbwWybQtTlKTawLcLLqo2s3cyhVIOWomzVpMIkHcizp0ValIW2i4yqiJm35pTPUP
KlNrEzovNqh5IOaosyLyq262apJvFfWN4EjyPuwAh2fGHGnY+2Rcc13a5IJtesuB
LGaXFS87nRtS8lX+dV9WGoy6mjCiEHxs8kYWKcxKyyuVskvR5gyVedWv75VRjk69
aUMnWffOvxsaIGWQLaMKuLq2LPTpjJhLEPogKiY28ya/U9ARO37D9RRw9qcMSC4k
Hw4K8b6cP+LJRTiWiuZgKAbgPPZ6nI/P7zOOMOad2HjAY5Hsty1zMMOaVUytPrtp
zMMAdF4YMCYgfL4W/FZWPK4awHGK1/7oUUMbTO8tFOk3yMJM8uq4ggOxZnCu1xp4
wfUXXyxL8z+U8BLzvXrPEdR32+l+MePVoV3MnvGoIY9Gb5CA/vAn2aGhNRFBoKo3
HGg/+fVmIB0tQyDLazDxghZuf/jh+qDPLDmchw3f6qjyn3TowU/1FAahbcmsmAD4
qJEmVHkiUu+JsG2MGsN/s6Qk2mQqlvyVANXSuuXvukgRiBIVGzeHkv8yTXGRf7dj
BGEVC1HtpedBRiql2Np2F2tijtPIa3hMOAuTQuX8TvfCHWAp0muY1mkjkL0DCepJ
zKXvNc6bp7du4iUo4jLuVy/KG1bhWaETxhtaJ9preyEHCOXCCNLZ7bXERsjNe0w4
RfVd8rFN6Dk185HGzqXj20YBIavkT8/NTOiePEF6Lwi5CJbm2l8z8+WhtuE7+baq
qc2eMIDFKuFD1ZNkCxwoB+zC64roivxbX3gwBjvsLVF+sQvifgi2/6WKOlzHG02z
kKa6vq2xrmgpi0sJPM3UpQTQ7UNiVEzXKH0UTYlqzvACLvzFs+ZRkq2yIeG0p813
eM9JztM8Wq5wogyTlUgeXVVNcuXd5ZnSoG61rowpv0QkKVWg5xaGRDe9sQYSRODU
O2xvGbuwuigADa00JQ4mm9VrBywqQ3u5JzJ0P7tq5AYBqL5gwXN20a0H57TJEgEs
Te6iLoEMGMj/k67HZsyURdzMNQ/N7lvhnuA24pQOrQ+Xt/w8Z2xNJsT2Ps23eZaQ
gb4M3vLT9phikQlLbQM8kP1wcdN4kAs0RNLS102XY56ZOOQLqVW/+B1TuxBQr67f
02M/kP0wiBhZvPdvOt+vRAU1Hcf48Jp9r3UYZ6xfrERbcC+qQJTTdvwWFb7cx9lJ
XAg5ARTJ4KyCtaK7TJD123FsYdNmeAHTbmo3WU5BRJJA78wJ3EvzT5lTPdZ80K4E
BMtjbLwTVfv+1fvD+iIYshZtZ6UH93IwwFRlnPjcECAek5ceC0JByOOMwANAGxR0
BtJy9FYzk3yCkOPZVq+MGtIwvehXuIo7IijQNz4ts8eo4UmbRw51C5APUTus+W/9
OHy6nCiNz/TZXZSBDnmOhjx2A9t7lik3goAqIXTR+97LbYqwjfyfAwNg5LOB4fzO
CArY9GieqELAJr/6QJN5FjbIctp2QTOwhQ86NKbsayL5SK8F0MiteCzZLk6h4gw7
ilhcidDQ8yJnFWyKi3+NjgGvkguwXovz6OytB2BtWy7iGOL8lC4+auartBuz1BPF
74HBSWWgick3ajMZDthczhZxkN79dUVbbK9nnH9rMXPT79t6vEObffZj07c9X8A3
xwskygsG83Pjr67VC98Y5jvoeCbTWLTQ0c2A+sCRFN77OnwL2mtN/pjri9ENVZaX
iaVqAwROFPQgC848yj2w7Jrq1I/z56UyJvCCSmmw9Gp0OI3/e6YKT6TxeKlXplNc
HjilfNVibDHHgEiwTQPoyvs0iV7PsSKLHRYl50WCknPt1jymkJ2Nz/RW39iijTxk
dsexyh4S+Xy61XpPKVIKAPexwz9K/mUR9Qh9chwQv2NzZloEDtuqAVO2WpFUitP2
iUbseTaKLh4YsUs78Uh7ZbujzMJzldU+yE417G3hnJs7Mr2MhofXjbX7gO6963AC
N0WZ5P8QCakAk4SM3RxodeVZjUIfvrRJhp632JiHH1E5NHlMXaXrEGD7m3EuSxnZ
W3l1TKTRg//kA52RUApDskM5ZqxX+/DW0g7dy2+00Foz+QC+9U4zz5yZw8N6qj30
MAmhVSsvfNskNtyUn4mSraBR4mU2szB62InPxq3AsDBKlP7P2+wbw1fiPVlvVfT4
RfEYRnlYw0ubTCQYiI+PDELLXJYEb2Gu5i7YjeWs2rfYSNUBWYXJsKYFiRadNREz
efuu6UUCrZHyxmwHRWN/SGPb0HdyHNCecncnJZKwlMuDnkDupuWoeS3vPkis2a/r
WPR41piW+7CPwMhHhc9/GkzWOn5eKS7X+tzg542zpkG2CdyJPxb0ToayvQZM1WgS
bxqgQRZZ1mBQRwOukW9kH0dXSuqZyN4aeFC8ap0NI6HUtT9JZGmILif52fjWPFpU
jMfEQdqrXL4/xJ4rrnHvk9D2sQZC40Ofin+GqgtJohLLbbFzBj2j6ALPcIAC0qXq
vrviERm3toyhTQ0P6YYniakgu56OaOBZ1Kd7d2MgsaAZzkCsalmouo1COXLkGBC7
AmraQxx7e5ivxS1HXBBxpf3eN+rSW8wcqbHO5SlHyEaVDdoudZSFehNKY/YjwhCx
8QWoLEA1cu3Bi4fAojIlssFerCf6COfSOH2KUTvzj5vvALOprbAaob9TbSaJ40ft
7NFr4+82gdN+kzHZ0Ek5UtwWRVBkGlz6iKKvd7NmoQCh8FrksH8xDa5wVSZMvGDr
OloI7ULYpgbLPscrN0jahJYwOpc+i8bQ971E03ilZ1eRTT2kGK9qQcOrz8JZ9DCM
/j83WUSreg/Uhj51hSpqwC1rnNzEDobo2hAINWWsYRZngW7BGKqTjA8xGvb1G1Gc
419ITFlBM5MeW2m+7o4//RYYXbkcQxU7SNjtxyH2hhrTJDQYoGfU8icY7h+qs4SW
a5FGmgjMaK/63DgDs05rWeQsjSrWBLd4XCCMkUoD0545h8mZaPODCdhH91Gw4hEB
enqSEDXmOwezbBq2+VlTFiLRyg2vSaGu2z2OtGfG7Xp8c3TmRNpqwbNS7chKhh6b
wm3DNeL/K77xNJvtmNALZel0z5wcZf89At2H8yVjiPZzEb/Y5U2OydMAlZuMWtB8
wQVdXfPBYNO9acWQk9LiRqXzl5LwAyMzyFDzDKzAJuzTEbF+Gb9RxSwl0x3qy2hO
XsazlMBIhPpN+gNTywg/SawqbpZmxszTPHpCGsQvQS4vAH/RqenMCW5HMagPoF/D
aRazkssHUC3hwGPJja0BlTqbGbriqn2injHTO/MAuw178lQxHh0j+c/4YqfMjd9N
emD6GfpNMtGEAnPmbdDBVv7DKQrl0gjab1r6kHu4JSceJqLqVgz2dtfNiAmWqzTj
qM67I4gwO0/OksQfFEXsCOFolNxOqHJVFmmEYAg9WurymVIXnIrP1StWTSRQjh1F
SNgJN+02ZXXtRcyZzJKhjdh2FoxgTdUXhPVPw+ZLiw8LDN3jCvjWeuEV+SkmyiQX
+W7ifx0ROoWm95Oso+525nHuJlm7LDyB/cGWfU8965Gqwkf/SKVNHLcZZ0zjZ0iJ
1y8oIwi1Yfa2TjVFSI9cQW/OhBiYu66TIj0R3FWt6Kqm3ZxD2kc10O+28JiChsEw
aNrv9MtsZnOUzzH4LRE2w94oP4bl0m0IUGI4dirpx2/sUC3lPBszpFh+ynZZbzYM
jJNi/SHuQCoE7HEMLDyZwkcAU5TREC/uLbEVDCLTIt5MfM9vxvthLV2AQ54pU7Ev
vl5oijdxJY2cxD6RgPGMxmYYteSrkBhFyHFd8XmH1iQsBwUfJuEzVDERZtvbZj1G
SZJ76zhgR/23uqnnFQTquGs5J8Zpp8uXN50K4UkDa5zf0DKSO9j4hoHg2q5c3Sf0
qHPw6TNhw0B+w6MdPriV7yft/xJjr50TODpI6jKZBqyvI1zVXTe0bh5z4AOsn9lI
qERU/uOEx8iczPmzlhwOtYR0dcbgAP5yy9cSYgstoKcg5sBf1PILtZ244QVC2SPq
190P5o87OIlTvjF/apWAeZHywQQ/uU/vp2bywDno4y5zNeEhytB+vGo1dK7BusAb
TN6BCK9xJN166IHi+StnUiNRU+tes80NPEVhibNgnpWjEcrfoCmMROF8TRiIpbgy
hEzgvQnfAJ0D2MTbaXKgEtIrDqHccKU5o4SMbsqZWQMInGeVI3lDT1XHDPgzt4z+
xzwg3U7FeH+SMeBp68KT1LvnzDzjJ83oW16aNNGrrmOwLjtQLpxY5uhb4d9Wvcm3
H3zYCrQ/cxqeXDw+aVX6ui9cjS5xituT59sPj7exRKb1LjnsGZ6nkdRJa/EhN0i8
mxE9LvTHY2VHaHxfzDU8Oqx3E7GZBuqWTXnMqwp1GCQxiLhKkdOmGK7b9ApvYv83
5kU6vRbOdLr1/nndhXAKFPw2RXhXEPN+60hGjO7tIsVxuwmLa2rqBp9g05jNg0JY
QA7eHHgy9jpajO8DBqElgtVeAqdfF7MxC5ShpZVUiTW7Tp+XSq2Nxjiqnx83wq9u
Iu549ap61sE+z/MDlm5HzHOI8/i4UeLaZGn9ufSh5MolrGpX/rXL3nl3p1Z2q5a9
b8zYg5MO5wWPoTEOblBbWCDH2Fff1FRSciaek31pDJuvnGGQ5fPxc0S8vIyHr3q8
S4oJvtdoA+fduzWljk3ejNLGMOuF4XRVz8t2DVgar6edZ1sybdRGtt0AXq1fVz4B
fJrf577Ge6zxdzr4tOcLEhCnFtQWgkuRXJ3ffDfUMyOjmB3Pdrm8biAbm6YvFyrR
oFdwsHyDOZzxpsdnVw6DSSlTOwKOSwzIJJ2a0Wq/FzruCI8egoDNwn62AisuhNls
Sb3Qs32jmb3moAFcELdypo7WZWKouEaIdsQtOgJRnS1X311EgXLr/SrmMb2zdmfk
Xo7YkKxUpbJoeyCtysV66Rc27RManhyE6okPv4qQtvCqKCVk12wDPSHdfh/jwkpG
2qx6dwo5l2LuZHWdOk/VHyGgBX3dJV3plERrf5FMsjk0W1NtIfjTo4IABj5b1xP2
fe1OnRWc1lhydX6CtBQZqEDJhAZLFJQn0pkvaA9UsKIeJHL5gAO4ibUeLGid302r
VWSpKoXR0mC/R2G3H8GDubmGD51m+rc04OsM0ryiNb7AqHq7sNUnWiRCitODXcYN
G8oE03uC9SBZ8HHguW/XCUSd9mTq6zpc0xfzXf9RShbgHQ2Id6EA1aPZh+vlMe5R
tLjgenSKWG+rg8dpZnfiuyUm1jJUKZjQ1IiEikApH3YGspF8qERQacpbEUKLfI0Z
7UGB6tUk+kvU77Le/6YAhR39u0fng4wsPWNv7mvqfk9PEgHo0FpsJJUxUM0yNpjf
qkOzgqijvBwlIhBMKtolmjuXQKDr9LY5Os0cmw0ocJsCHSzhwSMfOW50Dt7Tfm89
tX8Dxy+zIFWrI9Iq4F8A2pSzVZe1iBnvhORcgNZXhxrIx0K4XlyJvRCF0DJFbDNY
euKdbFosjsWb1DA4RNGrB6yXa7Vm399jC8WKfg+uZ5mvuciW+3jvJsPVIuXbIKms
+IwIQ5BzddKlp1QIcN+vVjZwCqaUe2S3e/hKGowGU+eSUyQqn57dMxtX6RM3W5WI
6YE0NDBXDgtUS93IDArcOounR3qI/Eml9hFXMxv4PESbPjtgNgJ/rbqZmGPDOOg+
JEvqJm/2BKKwaoqkB7daYYqEMIfZQbxk3odw0ftUlF6gCbTcck/SPGKxEEVefc7e
TtOPQylpeIQmNFaTHbc61hsYX+Prmi8EA+tVHyZUNAJzI+N8ZaS7fgELCL0c55oL
nbVzze6JU74fj4z6nn0TbdMchLUEFn9pcyoJ37ygb1TNv8/G6Qm0fTr05o0vofWA
ybVy+h+OGYudlg3sKmmDlqz6ssPabAQrFWXZptd+Zsayr+NBaCltvorollAnWhMb
Z9IVVEFgQl8QCBB4Pg3mCmL5k1o7G+eXGg41TXaYT3eUeXBj4rlf7xarApt35XfJ
yRyBaoZWqDND6WzQpz4LdYaV/6ONS+6qc6fINEjVI1DOvbFtySI343gh/OOPd/rh
baP+vhPIERNi4lV4VBRhgCFy8RWHWdw/xU9SpHM38bKU7uDL/2wYPeRNb9+rA4cg
DmoH4c59phivaXr41C/pjaPT6pXK+8z7ktiRlu1PdAJyiX8SFElU7+gqH2Oe162f
5ehiE79XlUyiIgjHMph+ACYOKDyjMGYIf/Lw+AKSXVAXCuN9B1qSldgLqxeCMYpp
bXJ8hrJ5rsmgVpO3nRY+VSF6/ocLBLEFW4pvPrmpa5FcRpeVzj6d8I9QMI6KX7+g
xb/VyBzgNoViKP7jaOHjw8CN0O8+J3JkBmSzRGhcK3RJzi1uZr7vGkHMvUdJKc5Q
mqEtMU0CepOpjKp0hDkAWFpGdpZYD3JfWOIi0PvZtvU/sXWuJSlkei0OPWcq4NpY
fj1ee4hTZMUySLMElnOehyWg/kwfLNprGyZXyYfEDivoeYvE9HqhrGR+7IUHdeb0
ONUkNNcTsjS7Yu9SCVuyPktsyBD3R16zH5Wqqun/Gn5IhwV/0wCGzXi6dPsi9sg+
th5QwU898shbZgGw3MacT2YdVlk169esn32GfEPxMq1joNL/9A0hqsL03n7+XRxS
ZnTtpR1ZRyseH0x4GUmvDBgldX+0DbdgpXJDAcuv645WMXCkcLzU0I/ZYer9TZuO
jO6WhvrZLJmncVBMpMW/DmLaDVc38PHzI1RRNSCtXE/IwQu0NNyyI2i0Z2+TUeJ+
KBru19v3aWbPQnQFZ7Gwy7A6N5ajzdahcXtYqQOI4lqDzLQxEhLqvH2nwXSY/g2f
vuHjEs8yPXmMGS/TcXFmAKIH2K08OvLwS3+/b71kKJO61voRvKnKl4GOViI9z0EK
fmKE0Bsa3IOct8fB2yPOUt0BOynUPhFaSq7TILU2lkF24TDBpq7G7WDswB6D4RzG
qIOt7zoJFBSKaliYSoPLtZ16iCAju5dfV/X3fjO9v3UulGd4r/9Fsr0SSWTp3izB
qKRWKpaWOeHhfnHoPJjf89Cj1HcmHNXviwGJYapCmtIA+D+/eOgczTH0rRmgFH+p
BTA/39xCCMgZZgrGeq/qhwLDg8uI4xl/JfUztUkAzp/U7xgQT93UzSZGVT5wmMX1
6Flg8Z+dgU2Dx6+vZrqYxZbrUaxV2YkElk8LOqjAweHjJfW8T89w1uGRthi/WCQb
Ef4U4dgmVANO3YA0aU6G3Mdiy6yuovcA00ygxQt7VycqZ1w3QChZQXNilsV6h4eW
bm8sDfFCUli9K+FetRi/fswfOulAMkYFRgEn9YlyIrQXBeHICG5iX8E0vnbNesd9
5gNziTiprzSmTTORjsCdV6sQATpBHHNg+v2QtdnRpUsTwvVJvYJv94gWDOdz/W7E
hXbl3zrdh7/KtBtpK4J2z6QdogeoDzmpQiK415MvTvYjJkBCVtL3LanrkoGMMnHX
uG9gNZwQW2/I/XWAu2uHFyFNZVrwnABO5hfZdZmc42WpJuKwBtJ0svQYADPDequ6
SIPydUnYBoMNzZEdfpa7/8duU5iWzjGDberUfHQzjoLBGvcj/JBqzcC5qhy/SgM1
5RHDco18QFEkxXKL3Xfu7W35zpOBAGTFJ/y9hWsnUBvSHCsAEQ+nJ3Bq8S9M6Lwl
qhTdnRuQR4g11sQDTFPkHEylXULqVi2MYJxga9gaWTa3KE89Ss6d3rGvJ5b8osyx
1Q7rKUS00AW6eD0bUZVa/yzsAD2FXV0hX0+BzHBLNSy1A6dW8p3r1SqkjNIgUVNf
h43xL/76uaew/HN/S9oPRfGSGhKXFXv/kM+ZmKzHhnWo7aOhuLLa/vVtnhBHFP+u
YddGcFxPkYUtwcAwhnRLNdY7rHAmS+TOc/6NI5CMPzSKv17BAeXvRpOQlVE87v/E
yTNqemAHSuyg4AnGA2vvjXa71Ciaou/UuFcMgXGV3G2Gna+xATOChX7fy9LCnmrH
Ijz14rj1T3cFilpdBZXwC9S/KA9XiJWZmt8q4Hje7GEPTyozV++j1MrnD3Jmil5h
tH5dNPCCfDelB23duX4UVuuhiAP3wU+xuNxpL1am/fubBIhZVSrs+dXim30Dj6sb
qgNI3FhMigicewJ+4xEYdL4TDDaArS0dcmwHLiSjnADygYIIKSYiGIOPRjwklr1+
L1ipwQD0aTztDol1IF71eb6kJnrZddY35jKIK7/AXqm4DEaZT8dvvxkM8Gqo8DgG
NblKcckThn7Y7E9ZbRl7lUz5PNJ9s2yJifLLM95ZgNYpCbz77DLfxRyJAZWcKadx
TmNq+idXlu8kCmg7DHO6znr4jrCVeMY9DYmfTHPQCiva9IhJoLHEck6+T5DPlCuS
MxNv70zYoGDeHnM547gOQZDEEgSRgfAXhitwpRPZUDlHDFQUi5ZK8aqBiHdCg2p6
QU7IDVM9HVou5HF5irAFANiysJIVBZ2GbXG2ynCOJduwwYCka8HLHtj81tpCTG1e
y4P5uNhsMrwaW+OfDnoth76vDA2xJ6ZFu/90HRYsaORI+uPujzSP5c0F2AiPEUVU
rKyW+dpyePC7Z67rAWFNZ94HBA7qVLbQIZGZpRBMZx0MMM7uKben5/P+9j3Iyyge
RsEQwzAwGhSZY6+OsAxPg7Q8AF1taojjTLlmHk85Iuw6ch21tkYBbBndaL/VX+pu
m2kzsRiXY95fw3wkM97iw/FdJQheKkZQwfZAPKFuiyzEl7qW+k4rbTTc6Wko77pM
AZfV+AlqGi0yCew/naH1t9WAYOieFqN4FVfSft2D2Mwegd0uLLlvbeOZ+0tjhvJd
nXeUb6FSbqVSkB8Jq41YIbc0GpL+i91TJRLOQuZQlJ7JNlLaT+KsECbUoZVhcyMU
pRLdWVK5OBA6OvAsTir1QIlYcoazKLESCLdpJ5lPX49WvAGboV12pX7Gz3b/xh4T
IKmuHbycBkKm96Hv5oVt8+HQxXKqiZjFMegXdw0mW9RFQE+LQHPPc9G5sKloPNJW
6aPp95MS2zAv3GqmNfxbZHGNZFg3IWWdaMak+aOH5/O+eLUe85USlbzTqF3J2ahV
T5mil/o1i/MdfJmn5+iYXzLaa1zVIbhsSB4oKflomOiJhYgJGH1u3o/AFUP+P1RK
v7d3XGy59KbQLqIThtmaRiL6KPhYe4TtS5xz18J5rsaBJ6SBZtJnzf2EpXBJjzle
sRQYFhv5cH+6zj/JCc0fwkSMK+qCTMD7YI5ulzsE3OlSm0ixllSNZrZ0drIUf1Sp
UFMTLpaMglSzRgFsyfu1sFpvHaANJujtPgcc/6dXoa/Ajwn3HVLqaB2P7QEFsWH4
xrJPsN0vNpAv0qqGddry1VTkMWGuP3WLFj5A3uleAGn+WbAbOg1MHw9pU0QP/Gfs
1TopKOcMhGP9YH2ZAkzofpxMXI4dIJah0om9NMO2tEGShXBIZy85tvF/sRpVqNsn
7+wCJ4z3klVK/fiUUmDKys6ZpIkgHNGbZUoCQdf9eMd4BJ97TctHPMCGSAPDsuIK
OeohNkB68Y2jfya8Josy291PU7dJo6hDI91RLy1mdA4HoValekL4kLWZ1ojl/4id
aLbtb2NWnEZNDx3ehru04XhMEj4XzhbOL6BMlT3IHPNqrm8I5/FNbjYZyZVaXZNB
rFf7ykyrKfU1J3maeviwdyj/hixF63c4wZUjhvb8ZF0etaeL4zxzo/lbSaxpwUO+
+8Oj2KXQ5XyzJ3ELl7eH+BWmto1d5Hn2Pz76bPniGb6ULwRzsvhrYebAo4nYGLKG
H/CovewWTtb9Se1OSLGujsn0arq1KswuPpmiKJ3pam0feIooOyxB6GJKsVsrABv0
vJEoUYrk104o7ny0fG/SwZRknUwP81r7xzmWIOeGkTNMiNYojmWNuy7Q6yWWYlV2
IqS1KuXjCPsgaQktZcITma9NM9YULM3pzWO2YXyVbWSu5OIdTZYHE3RolsDspFCS
dk6KzIjJD81HCKP91qXNYfd5OeJW2Pp+0W2WAoDTnHW5kQkK3Zxn92rCJjpnsMQ+
nA6JN7WWKtcwb/rZhvSKW4zz2o6ExngT1laggCqQCDywI64JFgJm20g4p4+Nlmjm
m1gJdHWuk1YLKWK3XVPEUPDJkTGJfIlM+jOOdoTvcXrU07V1Aepbu1Q21rnKEsX3
BUdA0visOOiiJmL9dqboUOjPlMAVJFLPwdY/DyyDN49uiBePU/y2WH/dlKBQq9Bo
boV7BVTm7J9FmyPxKEtNSWFZUdz+FDc2xkUKnD1SHXRg9K1lpo8E+u//kvMpQwvU
7oYPUo7SdV2wDPb5WvQTjZEgO1VGibJznCNT9V12CjLDKFt6kbDMr9iTsLVbYbiy
wwIdtjFARpXxo4nhV5Rrizy0G0I8K/JhXSKaT5V05PjaAsWkcxX0c4ihVRstAl5O
7v5C/w8ctvyusi7VcL8EpDXQrf/C5o08Lrg8E6Xn+oARIdUKv84j3j/ILUUZHddZ
n0cu5N9+o1QSZziMPXJs0snk+/ggxgaK6sCah9ujIzQIJqpXR5zmV2MoBmdneUPS
Vu3EQONyhIFLj9H2pAONJkTBRPWuuD4ZyWmGDNZYUTcljdBOSfMWPQ2hNSJJ89Ds
aGS2WsOP1k0ECM7OOSl+htud2pt1srWMCMkIT4io0pNqrQ0G5zDIzS8fiwhF0BJG
S+qCiFLhJX4II6O33NctiXcHQfSOUr2XAHQyR+2cvE43m9IVZA+39duAw1jcOJWn
uoNevThpotPgud4ocgK2WAn7oIe0CoYWQT+6ChKMMBDu6LumtSEJ0lHU3eBlvV2d
MtVGbRABjJsSx9Ar4sI8Kr/yc1LTq/3FoPURJLqMsRuPRlCJHnQdOso+F044M9si
QgqioUjTSdY4L57UsZuf0Tp2g5XVHVe2FbvluV5G/lmGxlc27CLiE+OEk1OVm1uA
0+l5LyoaBiKD4yUMIZ3zvsSmEJVM8n5PPE5u4PeF01a5E3EI+UDKu93P1wEly9WR
49/V779zBTpt0xb52BtONf5w81E/GqMVaoaoCThOJPfIJ0O7BKdlEC9OoiSyWyZj
MvGDQVtZACL3ZtnpgouZJnafo9+Rwq0PNQwv8xZ9wl91dlUUtprASbyO9DaO7hlE
qOU6bHShsxNsz5b5VuLHl2GC8yD/Ec97cc66PQscPCWazXbh4ia55e3fWxMLMlB8
dI/+d+/he8492WM25JQJTB8jSfx50WFikPNIAuZLSSrMci/KXPOkejj1Vddbwi2r
w027tW31mpv7tpoZB5EZDcJxmNNKprj+yr/wIJjsI4U3z9emS0Y9ZRGIjpmfnogi
AkFbAXFhjgo6PUuE5fRwhM+OghhsblPF8YJQRABiqwOZnXnb7pRjDSs0CXd8hRok
qbLW3JlLEhdma9ffSFt5WuqFLacd3Z8vJ771RD0ZZtEFh9RFgUbmW/foFEzgbjm7
TNGpDwod0IG+R6+YgGzYmIWJ7uTQOwZ44R7cWASY7rKEegs4DGCofstfg3PeyvWB
yxXbqHrFOAQVC1GZ/RlE/yZAFFTqCPlLwwa2a2XNtDdgdj4RcbIUfKu5xqLzfMWl
RSg1D6OzYBU8HgcSow0XeAdzXj+DzUuzSMo0HM3/uWlAoSEouaLm6215pqPQkFln
ovBUB3RPaSjspxdQa8TUCTShsO8Nus3tRoVDsIhfhLdkCAIJKiSQVAwBWrT20Yzf
sIgxQj0FrawcNsBge6nITlK74g0gr82AVjffDJ+RKtTVyJvYzP0MUP7PvUGnk2qX
D7bA4GH+bUDIhyr3vr6URpaFxnEY9LX/s80WWXvJIViikqnrYokfzuqtRngxmaxX
jSFXFggFwAYfahZH32LM0RXfDHEY9BBcaJr+cNGEVIEy35Ka/Rje33pSS+L6VcvD
1WXPrfPSmDw8/R5biKjfGpjlnHMjj83Ifv1tOIPw3lu4OzSUlkTGCnQ3ajDIccjk
x4Nln6un7e26CRvKqtwVOnqrztvRlN72GfZBMUsmOMPRxsfcgQM5ee2MygRqoK+q
lQOh20E/ngHaY2ZtHFbLH+TXic/ZziW1ikB6g+YcThDQTic+UNNjWjYvbQZCf1QZ
0ZRkdmQzY9qMNdvWFgRb6S2uLl+j+66aCRc+SPnSiBbSh9IIleP3bjN1YHEhvoX2
7b9/gvVTCgUybjjEzN5zUENB1Xm7BL9/3tWVnUyr7MtqqB9DngzHkqEl69099FTo
fvBr2dxvGZw87YbOuHXlQ0SuBCJ99YruTfVHVNwtCaQGFZrCexDgwjQ2T+HP2Eg5
rsTKNmXjN/8okWhG/rn7xVW2tBV2N/eA/UcgUY3vtJ07Tr9T54/ie5GKLKwnMe/B
f+h746fWU4ci2i/NHfNnBxHC10NB9lHY+BMIiQVREmCMgEaa1+mbNK0IeovhODye
ZCr8Bn7i1RI0EN1nx4iSVrripFdl+Mc3OuWmVvLfZVVNGnRuCwUK5IavqQIC4V8+
2jHyJktHmr1ZbPb1QgreSekk5mnUkYtpTJWBp3Hfv+9JQ3SKjrTMk7MLG/U+B02Q
5YSveGPgZNqhPy4sHK7dMfgsDEE35Vi5IvaTSiQvC/SUT6XmUQdGjXi/rD7+bl4t
3K1Fpi/Nn0z1jqa1fHQC6LPeSvmgu5TJ8b/1Rfggqhj2I8olY57I99mxgBRizQuI
S0+OECCdjcXT/P7VPH3ONpY8VPxr6iYxOGM+ViDGRIxFBKxFXQAYthEriyTV+HlZ
qU0AW/drjgrz8jN/5lVkqiYGc0AfQR6xfHKw+J1wSkvuSUPTiVunZHgvsBuPTy9r
eger5V2NsGnFVLlpjJ2Owly2ncln8ySJQSfq9gAyb7G1Sn4PY52vFuqwUUMyy1DP
0QteL9T5RlyJo42AEwUq940kaKaGnfJcJkDKZRLBS+kG17LoeKp/QEGj0m7J2hwR
FG/UUKfnHLqae+mWcn2q85xYYz48lGkMuyWVkjCmqzn0XtdrlMqcAw2TRDt8YZ/P
M4WyMMGx4KInLgFvcMaY1r1C4yqNzpfKf7H7wCDjUu6baQNtB3O5cN/BMZ9+jTsg
tFwhHp4C+0qHlmFvAjbgBuwD3l95ROIDq+hZFodk7+ZDPnbymnwSzBogV6ls+xrh
bDaK5GR/7xSqgWye0m3/GgPv7pNl2edY4T9u2V8UnIkD8mH3QuwmGz/jEx8ZUm7m
0EGT+Nm9xewRW9LKWBjPaV5DNDt7iyn+OOd4OE4LolMemx2Uj9dcl53TEnq15Ndp
bvqpa2GCQ5xv9mzGo3H6iI5RlBfAshIuRReXobt1B0YOkpMCAcDjFeIol+XwjMR6
CpRRuF2qOAtuD5Gy1Es3vxQebifV/6CclMqQUjvU8zE1qASTekiu/02zASuMbMGn
fO0yUron/Hf8LKtIu4Ml1VnS5m/gfOaiBqNLdl5AWHHcAZqPf4Fo09ZntwWfYFZl
LnvtVekUoTMIU/4xuhf4tdbAz7/YnjRIQdslntIRtICnwwMN1tZCrc4CZIUlK3ZF
r/zlY9iu+kda1LuVRpGCrdxF797d+1Hj7Gog10hwjdcpVGmNi3tr2CeH6ADbqjcX
kcYogCInMj2HwW8uYYtZhAaDYfbhs4Gqr7KafzNKdHp+fmu6x18iy4+vM5OwYUXO
c74WC20mobIX88oAgTWQzloi7FIYEH8oYViSkXto/Em2NJTrg4AebmAD0G21zw5p
9g3pdWVlTCKTyeowvLL6LITti4kg1Y2L4uF1AqkdweGPI29HhfJomTu+poORJWvV
kO7P9mOZ2/Oci3e4pr+A2dW6ltnDlNZJ36fnaYq2sS1lCQFffNbAcxir8cQ9IeVB
sOJwi27y1qRZTN0AHvEQPMHcXGrygBYwbybBsCGZjkm4mvjJ/WNEHMHmtO0SHpy9
eDprz7UWX0StiBFEVIGd7xqvYU7of/BAbt+BQ8VrtGZ204WRQZ//Y3oN6RPOUcET
gJiLzMW7eMsP9LWaVUJovNFJ7G/1AMzUwydUwyL5fc7Q5NaqayRo5Aaq4bNEu8fa
lDw7P1m7scPiIdluM9Sep2VG2F4ioxtKtHhHh0aY5NQ5GGGlmavlf7ArmhPibbuP
3iiTZHxR3ai5e86OBXAb3rXox3YBo8cxEfj/n2zn293gvvPgnH09KDSN7620wxYp
lEJiKC7lUnUfHcceLuvRm22OZAbxVT9oOO8sEKIPKdzmHgj2b23nhyhvjdzf/xG+
FmWqNUYbgSKltSF+ffbRRaxklmgfCDnmtH4rjlGw5idz2j9kNPxPHCqHHq3Mi9TF
smQtroKaquejyEv0qpW9aBeI4XdUP9YsGf90Rq7Qr9p1lpyoVbItIE5Z6VeFDedR
HAm85WgmAdwGugKoXVgyuH3JnJsvrcVNi5K7xOsX1TbegOt4w+chUjWCHm7O26xi
UyYKEf5db3ZzL2mYpyVD1+cr/BA/KAM2dv0X4XeAHiioy3pD2AQcmpOU/9kGstJ4
quYiEnQFV8lc9n3fRB8MP4vfh+8L7cqXF82PGxpeLtHf2JpyswVSiv+yFxf/aJxF
VCH/4SoASlz0WkGk1wRtHsk7nvQj/tUMtug3ryteN88LjhdmsRIISSS0eSFlkyvn
fFeNiTItBWHTCev4VzrdirO3MU3Ejfz5Vh6xAD/fy2J3UvMemTzWgZ7iVJOAMGel
ybWwUvLpJupYG3jueZE58ZXBQ4ffUAQafI1fxim5jvDe1XlLfLNQki8q+xEAB978
WJueHSQ7t5N5wdPQAPXj+MPA1eg59bC55jOIY80UkQpCQO0dtBg9HedxHB2/wOUL
4CH1T4KWYjkKa/2J/L9jxo5t+3wS9ECE8EhvZWA5Y2n3REEn6nCb8N7Q3hw3ZUkZ
n0Ny/7e6QEFi8nqXjsytWAEoYyJX6IMXA7ngi8Wln1wHYkQZwmdL0SgHGcsO2LU2
+I6wYNnCHHfvFKDigJY0DdCm8vahQPb5RUFikIXIOgPR1FxODYTFcDF8uKEIGqWf
XEIVaGF2STjLeRbkydKO0imon443xdIMY6Ch94jHC+ISGjg0AAGKaEklSkFM3php
/VcITaJg0k4bCK5Qvcsw0lpLGS3DiRW7Ajx8QZ64359Tr6BB4ARnIKow0vDONYiv
qhDYCMBTrf2JtyihQt7QsA5PBWwSIEKv2bklx4hgdkM3PU0dH2O+u+KsdPS3buKF
14hZ5FeLzNBcjzPyHRwIFJ6v0esEGlMyOkd8F2NtdxBpqZphV8KvIcfzC4JrE1Dv
FjDgUqJaHzXC/oWv8Vud+S7XoSCeR8IYfgNzh424s7y9xCwDLLVBFK5St7LgsGOA
8ktXa1ZWj74yGNbgw+i4GfsB6X6jklrLi5Ng0f1CkfbDxufmAr73Ls2Ck6qn5QTR
ojQUZy9cU1+9Y0wm6W1ne2jzxAyvT6/IFc+qyy4WnKYdVdxCIQvI8b3drw+NxCjS
NYICSF+MLhEEsOILkgF/KgJLOzSlQh+SgYhy87X5LhKNeXE+hWcWxFabRo36HKGR
SbpCq86b0I0Cg7CBvoSEcUZj4p5A4/QSV9cTce8JuHjmY0Xdb929uo/FRrMZAeRC
6ifXqpTL4Yj0a42xm6SZ2BVeiZc+kmVg2l+usKet8vEBUflp+lPy8l4ITolsTvyH
iSHvXLtSj3zvf+h3h54rhrmH3nUE9kcNyXbBXHwPRukT0ZTD8EfF8AfGrrfxMpCW
POVMYWv8Jl6h0kJRwwFR/Eab0WUKEMAcZCORemeAd7lt6DKVKUCWx6duDrodRDm8
Ft8MnTnZHXnWmCFbhEDi+f0cBQ9/zM2LNv0+B1kGfPYnZNMl8xi8wbssU8DzpGDL
1V5jkIiV0BRjWb/xXtvZnVCi3aNk0wsMEzTVtnUVtrMeq0dLGJLSZ6yVeYUUOwSd
XjODykS6Doc7BBVKexRYY/1zfRcZ9C53DtBT1C9HCBMmyfLqhW3fJmAdzeKI4egm
21HhiEdcCNnsyGOpFocPEMuUW+9luZ/RrOVyko6i7pPHprub2Kfe3wygBTZ8eE0p
KtCrAw48bdqoSS04QLTfiR/m/B3l44sI0ENW3e8qoDw95dy/++truqNnWUVoGQZo
WtKnMC2w9uuIt+3q1mekj51NWhp58BiiR+TbrZ0gSS003QYGBMzUQjRXzvbvpf9B
+AAIG0Ty2niGew3q+6dmsSkxSZbZ2mbGsfxXvb0tdtBzFsDwrLjhXZIbiYcIYlu9
CAsyUzxibqzxqVXrmxQphIqFDFZx7lHQ1At6rJFRQbPI9j/4Cm40artMPz/J0hxS
HEGRJbwgHVHkRk2l5o1VebONMJtFQ0jYILlr5qpsuSnedBzRMLfiy06Y0Pe7lndt
Z43laRHsgS0MkjBQPxQmtJLbLgwirabl+CwYlkTega+J/ZaiSvzeT1QO25mu1UBz
zkBerwIHJXn/kF3K0zsKo7WHJ414E0VSzD/RY4SnWbm0fg5rwiXXgVO2uP0zCgdb
1tv3r7pllW1uObxUT7CgVfLFn5TWncqV7Il9QPcpfJvnuZ0KHKf81e5WfKUiH81j
yGgDWTmpQZZkpGG7F41nFMt9IWqxomE+kHXTgcWSJNgWOdHmfq4u7CBXTrvwrl3e
mcyju/UqwfDS3fDBKqJsPDSbqAWYIPiXauwBKTlrAKFOh8WRXwlmQ08RcEbzO8b2
QkVPvGst8vxRwuV0PlwZbdlMfzBrC1OcsvOwi+XY1dKwiYln0FkEwOeuyuyYqC3z
koEPUbTTAVj7ckD3iqzBoXWiYeAo1aLUoxebV7ikZ4KF0ZZx/52hbE0eP18DIlan
3GWPvnl3aUX+bYGEImkEEGKitbHfd70K4cdfS55d/fzEkV2dHQQY10Okd9P5bgJG
QnbzIPA/VVLrC+nPnrFZ4k1SjgQLCEwjQKXjAtZVt3MCJbeaG9oXBjd4sWfDyEqb
2YcCDubAGcA2Q0/HoiVo8GdwLOHoJb6OhxT8TKFUoTb++hNbCX13cWLXt4J6XKc3
S4Q4nurjZUUkaOh6A7itZolOK5TcH0jDd8DnrDdlTCaRzDWt0Um+npoHICMIrGFh
X88Ja1v4afKP++Bm6Iyv/Iivp4bKRePevN4OZyCg2AETFDy4Yz0B9Yy0XlRAw4is
hOLUXV1w0YfDO0Es0ZMsuFKo6K52PduTurMB8K2sNzQ9I1gDHQsiOMNHyBaKoaTQ
xo1CZxwIoAtLUdxbtr5BHlFvAiB+fCJ562NPbgVBShDII/FpSOwSy/r6RwREoARa
FD3HNQN11fdZQbXpexlb6VXfETH9iI6IE7IgHWQzgiEkdDpCNiFqOtOVgPaiwMHM
v878IU/n0e9C9R2HgPbT/Q4/EDHRQVeCJStsAflxdjlwq7Mhhzr9e9oULXQlj40v
n3lHuY7BctMljlrGnud/j01zpL9a3j8Uo9F8pBh2YZtYzHztpR8z47qK/ZQgQdSU
1U6/ppK3Ahioi0fmOj79pO4yLhsVRfqUW4P2lX8XtiCsLl2VjnKzJoqSr8H6No2N
FCds1PLHpvTG0yMtCBdv+HRG5+SK+0S8/SL3NqNq3O7LIH4erlnLXU40jjzq96N6
dxl7sReOUpWW72vXH9Ffot2s0ra6t1ijtC01EgRi7HkHHZaem9Ht2srFefqT5so7
LMZY2IcJdqtH4bDeYj/ncqqJhHavXVH/78XTiJPVAdoKimittBd5/xe6mIUDj6Ir
O1LOHw58XOgrn5ZYG4/PO6NDThIQQ9HI4VP7dfebeFKggLoRqhFBztHYYJtIKgBu
fe783sh4hL1xJFovqXJZHUQ5da+9BK+rwY9nrIJezFgWWWWxVdJa9eaT7RWU4Mjo
Dk2dZsg+FemxZCWeUV0Oxzno+X0t8mhbzCF75FYrn6ee+eJaxOgYSndRPM3coMuh
nbDtK1S03FrRwPDTq21KK0bo3ezQKbOM9aLZakujA+pOTFMSffyg8ADFkGGMCdiJ
rrsFDVKzsgUU/v4oDEbBczXjlaCawxDw9QBfORIE634Bkk8cLXVehDVUKhHHIG5o
Djxgrxr2iYoT/JZLYp1a6CpiBG+TtaMDjKBsu/+rB/vE77oH8N9s4PRbQJqBXbuH
KT5TSrODY8MexxVAC8ndSaYl+zhvWGpCeu8RLxRoasWO+Eihk+9oY+H/kWN7LkcU
WKmLEDaix/SC0UbqZMgt2zXmQKuuTwH6x6b/ylA5X4kI8qJDYbC/PJrlof0GTJOA
HFp5g30gJiMfTRSxcPJJ8E1xV2h//T5LpHk1TqS0kz4izpWCI6zv7tVNjjYRdyA9
U83yz5pSm0iktTCdQlpGxlOh047qSdIRj8MGkc6xGoXLPlO0j2/KYr8grugq6+tR
cauqPx2+ngRtzE74QUHLePMO2GSjFTBO5Ipw4Uc0oC7REOZ/k+ShubgOtstKsQPE
d4rFcRcunQeX61LzmZIT5MHV8/uwL0mCKbvHkxk6zEVaYqJOtf8CRceiSTOzvFX+
llk4CsKRj+sIpXR1Ddu77M4MpUHP7M9Nu/jop1I3325bmJhrb6a8MjIC7Y0garFx
G2LpUOCl2e7EQGENayqcBYoeb61ra0r+tRfOz2kmP9D5YrOyIR1Macla6vcDXzqe
FPvRbSh+brto7HiQzOxcL8r0DZb3zhlfL9ez6mPhLdfldC2JIsKUSMFmTBAWtk9l
2m856waF9ObALiFSZHZvDajiJvBlFbwjCKYmE+dY1Aaq45ZcVNj96MHzAprugrCL
Tjbjdf44/mIDJgBmAqsEVHoNKX2J//LPa//CXKPMd/7Y80uYfPKZGYZxLiwDpHMR
u4kvCXly8zcqEzRP/4Ocl8RRyRxWpC0PNYT2ivPQx6YF2+5fRo5Xzz4liSxGkjc0
8+QXrHoFcE4ZrgUxgrGXvE0gmbqDTdrHSGBKLuxGQfLWx7kv5rL3KJsbGiOe2g6C
S3JKOTQ5fnRC9S8O4wzGGGGUMrjTnwlL8uvGLzo5JCNnobpMS04ihDCQ2zm0RLYE
Bc8KBSk5lOSuFwZODNkgLLW0jCjzMrtLr+fEUYr5VbAp4Njfp3abHVOINuMDTIe9
IiTM3cvjhPyU75gMgKBZR13zRiYryLpVuqbhSzY749hL8Ir9VQxADNoiydQ+OLyY
NUfqB9dSwEiNuH/2oWpI04cIQklESODoPeX41zHdLAUQutFN2PWRI604wngxagt5
jbNhMP1otKSUq211oWgE08BNBj2M4vgxN83id1ri/jbE/rApNAXU82qq7jwevTQD
iIQwqm+qMYoPvwD4AG5y2cCxVffNghZq/Lpib6i+/laJ+tinXUDYt0Cj83LJELEf
/DU5mecYZOHOqS3AfSMdJkTXsBzsKLsTexNSFzDf6CI8sBfa3kTsMW69onk673QD
DkqTKrOXwmrrUplNyF66qxJmk+GaLpBJoODNtwNYl2HkftMUfINprnCcFgJsrHrb
9fJlgi5rPThjT6NL56/TTAdUcyNIBoFvdNiqbeLq0LDxa6+zWZOZIJTUUIpvxE6P
6Rv7fMx/b/0BysypawmFHtPh02dhNLJGdb7lOO57wy/a5/kZVsx8mtHrJgF3Rmog
2s3k6hLGSEPTf5fFSXopEiMQRL0WqAHB3u2PVVlM+Pu7QkEqTVCfF73imExw9Ob0
vVYfkr2W96p1BzGlHzgeffizjAjBo4mbb5SIEJDLE/ATa2sasFbCcmDSAzGtMa8t
fi41kXDgitU/T7MiXtzN5CdA0+LbVU0gKvOKVcur+gdYj5resZZIXI+1CPSRyjb2
sbO2cakRZJbBbe1dSw2Hy8Ud2TYgPDiI/art/ATXHPeF/0D44f0S71uf/BaqvcbF
+yPUQEUKEUs/SaT0gZQEe9px7hRxoNO7dpOorLvKd4ohd4mZuddZRPyHE7YE2Yk1
e5WPPTUkt+mq+tbzvpvZXGPxyEG0Itbe0NlJ9S9v2xDbQRnElrjCAwm7Ls+SetIB
32DqXHTROdvpxwxwcesWPTRv70I5ST6BHyPFaz/YRduz0oka0M5EupEa1IDNgunS
3Rc1QBdtMYpIe8RbBZnSol57FDX2WNsmSUSnh3cpBpyPZMImMbcpLtA1ExDOA8Jv
nL4UOTVXUa5uXUDF9nmHKWHliElSLwDpaBETxknL0XwxeO7nxEjJLhHlzLXH3WVy
M6OUI6J66yNrxM83Rkq3JN4tRlFPaXUjW+pNPa7NkJWmS41W4nNOYvPpt+utOAQr
9vfn1/JftFuGFiZaEJ1WKNN2XbMtqBrEOy7gJrtqQW5Fvpri2Ilj9r2G2AlGELui
HR9zdX0r+Sk3yKqYhMTU/Q7WBjthX2LyTnm+XbhX/h1tXUcBYFaiwlvtgGA/v6Iw
SFBG3kC7Wwk6Qzxq9HZZPY/Reu/OI0jaLo7py5elhxA6EQWroYg3wkXlWfQjJuSZ
sgPmvpa8rqSwq2fzJsQyMeFQUxtwV/4Kyy285OqDkX7b8O8teXmouIJ+Z0Z42Yq3
OGaXxG4FbdNTD2pokGkhRIQZbdhxpbPQz0ROaYC3Ui3ZWEXC6D5fn7tszIKI0Vug
buwJmXEvaPrsPNxDzgnhqonTJ9hiHS1CQCIqnw458UIGj12QFI5SDUnORSfjnOW3
81srG/sWJntlWi577PtY5dxlDq63qkjSsuaku9CV5V4nxrHeOJ+tryEu14S9n2y3
NsyZw7xSq4Mt3AJAPVegiApxVWP0icYyYJOxogFL30upZIFzPVV32JXs06oES/l2
t1UOHG++rB6vMLkUJCcoL4sP8rACYuNlwnb9rA3aTU/pFezLfgSSdpE5eR5ypP2t
bqVCHF1/rdSIOUtMNgT1ronI/ooVgfq6WKX8e5id9gApFX8nlM7m/osUzIySBTMB
AzWxHsyUxcAI3yQfqBH00TCqbYWa6aNbGNF9oJhq4FpIrDjNJtq+p5aCKYf9ooXx
WM4oW7MM0/tUjtFV0fU7GZlfyeoqF3mQh/+NbWM6uADtTZbOPaefHgTv9eYXGUa7
bzfV13bDk0Ii5iAqChlcxXybQUfWj/zZMsbHCRwrs1WctcvhwLWhyvKE1KTKJXUZ
2DeTaD7WS0loMXZXeT7BaZvnxw7RRqKUVUuIcuM576NUfvpn06Yy0t8NnDICnAUT
cgdGGT7mmribAXyYMrVoTOawahUDzxq7UU54U+XtBUKydHOkv37M2oEMHSI/C0Kt
c0Z54s8lZg4sumL0b2Sok479eIU3hQHdhjR7/xPM9LTA4PVMm2Xd/0RyKkDfx81b
8i/SwoQHUnI6oEJbeXuup6j7a5z8toV0UYPabtVTkKu8vnqO5hpgiTDYfYawRv2W
bYX7nTSavnOiKt5fKqJOAPegjPwPOBtfuFu4HFcov1J/3QG4DC1CBZu0BL86/5Az
4X5rmngoWONk5YXoHvXVmYMz+bLLeh/MB4HZUfzgknemWvx2YJudlqAO0u6X1WB4
gjnnA5t/BiVYSdGZgBzPVTuyQh2BW5rd+E7zhRKexbAY3bVhvHtQcHiTh/dnw1rQ
e/0Ktf5IJb13Tby/kLJbatf8pNfKAuRYIaeoQFHiDnT9Vum+l9EtY6FO010/Q1c4
i1j0mxDi1MmwZ7mOk2G8vJk855xZrUNGEWey5W3Fp0WNgRIgYynt6ZLojdXVjuBB
9G5cXXbXyrkYKuXRGlv4QpmVncMFBnCZOqxy9jnOTJ/MOLu34VNmxZ8xIQaoBmDF
l1W2eE971QTwD5sDskP28iM5YwHNxO6yeRyAnOR6plEhS4L10A/3HZMMBQFEMFS9
oeZqmiWQZBvtszzjdMl4aFiW43lNBS6qjnJZ9n3SNGGbFe/O0g9Z9My9+dfia6kp
V3WgMqjSCYx4C763H2rVcFU6nKTnXxda7EZtpFqhyb7LZLMn+UWqObUxCT/TT5j/
jCSH2LQM7r6LXV8ffuNoTIhrIZbSi+eIhGZX74VJl4yxCzSCB+0tWMjA1/SBPN5l
JqH5wODjDlGHK+hz5ahY102ouenLzjr+281jr0lHXhyCCeJH+U7paHjaTF145N14
v9WxJj0NwpYfRVx1w6OjrNN9C7m6aZuqzNoTWjnvsAWIvQWLHGb+rOJdHPVBQb7a
DVuvEihcmgqAED5S8Pt69icW1sPOuIW/P2fgAJxaWkVG7DGvij4NvGPKwbJ0Pvl1
59oErdquG+oohYgwJMe7Ed7NrWKoq4TjUfYV4mY1LzI9GJGWQnDTLcwPRaQnsefl
o5pHV1uWKjbci7zIzF1+qyBD1D1Q8Jl3uykebZ19FLsDL+N8el46lzH7WjPqWfzM
eCgCJCiePLzJ965AkiSXBmNp9LakI93uNHHmWtE3vpqNarZX472SiXGrR9DNUl1G
iKrarStjRPakmU2RkkQ8wdm1Kl+lmZ4gd25kOEy7J+/Jqp4SYr7vdmbeTl3+rKRD
0jEoa9DQotVViqpzcaduXBOc6WbrGbz7Do+eGXOlKRgnHyrymDZLnvCZP9cvhL1e
lfD/MZHGwLX/6DyXZNZRtjBxogNZuJEo74oVdfmndwAEQki/xwux/yxhhOcc2qPv
WB3DDpV/8aGqBS6EndhehaZwojHbdz15M1Zcp6v50ziLG8p9lS5+4olCjH7xZ7+B
V7L22cCi4gC1sqpQXQk699uCIN+LGXrvZtA5rrEnfdf6x+2mwgA78dGkw+wXu3kz
3GKK0rR+VDpDt6KMEVFK9jaojJ3H+0vgFy+CEBqtD9VJjCMQtjXqW0jdgmYrov8r
k5TLa7bGeB92Tg9iNuABHfx5JYHfKeE4AEu85yB9J9zLCz2W565oFBWEngzRquCg
N7nPEUPx/o4GLlbXik1PH+ng4ilzLHiC0t45vm8fUzVIuOEDenO22nAhugw1MW8B
6ZrAcRE36aGxFe/HRG1qMwdfHMoh3j9zVX8IfxpBmMd+Vb0IYNIrXLuX1OKYhuc+
p+R716MXrCOKd2uKkqtk27+mJkm3bBN3qIvU7Umy6BPPqyLb5sp99Yvqq8bEWLaj
nXFJfUWUrGyNjC9b5STt1prhUsC+OUyLgfpPw+cEOzyUU0zGsg0+VDbcMenQ3REq
7i/I2Cn1o9UkLQ+0qnAQee1I0QhZhGH5JIZrFNWQXFXKLOl/yMp2ePMynQnTAosO
1ngMJmoZLusWpAZdbpZD1TvXrKDuXJ1JCVF0mslJEoIwSbyVz6uV5WqgWqkJGHTx
nGVAuRZ+ANbtzr5TFRZ1EfNlQoUh31c5A9FLE7N6+C0EfDEIke7TaXl3YwArrojy
HkTEl54SmvZ81lA2rzF5L7YOtcDRp3/X2sJH8G830GnkNcz1oe73A2s35zR6vfxg
7atJ5V1ESaWhA48r44zgRPIcjMInrXuIreZZNfy6njGfhSt+8FK1B/R9JkC1ecOT
8fl5d+JjG0jxkgZT3n4k+dy9D065VQEJXj7hY9waLNf+at4iiNwjJhQ+InwTNQTY
7ka+4S7fDcGFxBZsh2PR8Cs7KkKBUYbDGciSpqSw+1KGSmSdzbaMuXLg6Ld/Tx55
6gNB96OpJcp9lnvNGlkeybTh2CNs8Tmtk45r+O726fanuZBsIp1uhePmepcXYRjx
kDYB6i4idwkXfKBd9+lUpXfx/Et5/JzixvNknoeua8YZLmNaA2T3aeF9evCllaX6
3izcENGXee1+LxRoO3mDNX6mjJVLWkc6VDe82FRjLJJMCMG6ZXwTYC5giBx4HvMR
AzYsvA01GnyQAIPJ9ikllC5Fb/IFo62XsfcGrS5VJ4qYOfZBpuKdTQAtt8TsDFry
s5ZWHmHWGMUY3jZn30WSV9nDoQHTjuaraP5vPLH8RrCcr2dMriMGE8vY32OPXg7N
2/IOQKbhnlsqpInfH6kN686f1gnfFXJPDrn/IdOJGO4Cw1/iZjdvEVAK8HNneXux
sS1K70HtokV070SPGCct+/6Mcilx/bRFCRffYNEgbzy7AXae5wIs6CRsZYIi41JF
PkpBobvIH+TlrQmdYNxezjTulSrzQUVSmmfCwerH7OE1EEzagHs8IOJd9T+9ucDg
3RnF2Pq9VQlSb5LhC3HLd5QtSwPf/3Lycg5YHcjgIFCOtQXFDFPgH6h9jTKLFIN2
X/sJTQedmKhpE8vNk3h1IcMCC0nQgaazzvbG+UBgQPaOksTueNfsoETap6ThCaCB
vSL5VC2lzrVWsgFma7Qs7gxpopwPREE1tzdLyAAzeFdho+SRBvuxCPAZTMDJLiKn
S2EZbAfiGfp+eUNuvfd6lWy80r4gUODbwi8OpZgTcgHvQSFFwJ6aRGIImD1x5ZIP
1RA+aWEaN6fLZ81Zru7RkZCCIsoVE80gAiV0D6skWa1TsCszGPdmra/1XFbXf9W5
bqNFF/DT8PlFb+qquMRtgw==
`protect end_protected