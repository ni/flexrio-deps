`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14608 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmWdo24EC1SLhDeUV9o12ewQ
ulXp2xSZ5P2RSggIKJUy/anaBVTumwtXp6e/AWaEducb/8FQ0ZrUn+5N+LXp7t8O
LmuhF8Fni2/94kc/UZwTeEbBwen9S5qZJ2aZ5HOAGlo46RaS8abaBfkBQdawT4GT
vgjMErR+L3owar6Cw9c5g7Mb8lgNMYHovt6l5EmBldQrGgdkV/h30GVsRaArfbVz
rJDEZ841WGkfYGUYH9lgIuSOXV8oMfg4a1cvUWC02S372V4jTKH3kdSlZzOpgW6Y
Pz/PdtsIxpUxpQJ+nQuEWWpD/Adio8+SVFiYOhLu8BIWjZP3/ZqWx3v2dfgZsTgR
Zscck7baOUNgHwLA72Xldi7uaISRWFt3yLoL9Hqoo8LatWKqmQ7Z8wH6APzxlScn
kETKKWkk+zLWRD9+8+zW0psB8L3msdTLwHzUHH/ZFJHt/QcA6YF75CI+hSYFMkXz
QsxATLkB+aYVMrChCZZUApuPo1D55phBGUHI+xxwN+/G2D6FBzvX3/c0qUSSwakB
r4tdCRrjInvo0XgjHI5xKmT8lbhYaKKtiBq2XVLiz8DD/0DdbM6gGX8so+XkH9xC
LrXSoTWQXvAdllZNH4JA0afa62zEo3k1NyRqW9IsbuZfujWcGxixL91HjCWczrf1
DzSovw0yF64+8QlCdDLU3FLqECmZ1+OwSAz1ZWS6v20KN56JiTq150EqoPIhp6JN
nw/8u+y3NCWTuvBFpSRA2Dcfxodkyis0W+kGxKI+O4arQRGtly1sQIRq5mo5G+TY
jGYkZECFwlDdEMEK56zEncK9bgf9yryfVFeCcDTU6eNdsgxZc8qCxBCIJGxwn0lH
KuB+eTdsImg3zS95GWbL9tyVH+wHd4U9YEPkhQ1u73vFM/GGIEz+gwjbO3IAd76o
Enr8v9VlBoTHSdZoMzfb7q6PlHMOLsLA0p+ZJdsZNsZjvB2mh8UIDxtUAkMTcjIG
I5hD5oIRCk3UzYN8SuJjawyv82KQK7rPAtHyY4MVTRp2Q19mmhCyjGFuLvAYrOpi
+MJzBC1rGv4EyjN7lHT6fHXKeu7c8RFSffpNOoOAI+ZO7PyxPlAqEhF/KFm1fGti
HdkG+NZ6lGM81fQpPWinI4nHHDLAH7hErSNM7xmtPnvAeKnVGgLEpctCgpsW/FK1
LkLR0rHOW3bCpg6vpOtg2rB8IjG9nBDsBoTNsZ9xp3qQIs6PVvUX76vnqpX6P0Rk
BzgN51RwExs71952ZHOphsNBsP8SSY9YD4W+PHshv6HreBs3SEawUqXohhVOJq/U
PcghiSQ62MRseDfuXfq/50eEjsizTMNwUid+nV+Y7+wdq9ZuTBEa1Z14kKdBmCfM
OVDR5RRCUUXdsRBLXrDBtiq7NFDNsnRoOmYjH5kwjusdteaS/2XiZ9hKnVjwu7jw
Tq3aSs+edqu3yAZu5t4G0dj8IEFYojWpAqfB339+Ohxuhc0vHhDNOCifskslQNun
Wj01EgpFf0QtrT67S8rruZ02m7i6F7ytVdX/GmqrzlfxvZRL7wiNHcBcyYz0R1ET
xUGVvyfjvlXfmMH7Zi656BXvnh0HuE1WBFxgZVquaBcZ2lrODCeUzuOUKfgzorch
j6vYZRi2OV4K4Et84Lw8YoVdnspw2Z8X4Psttljoa7sSQyRBeugzxw/5D2PQPQBB
xvc3McmPWBhDxRqGuipUeoRw3aawwHsI70RqnifIsZ6Lf7Gdtf329CoOX/7UeuX6
ikWN0/2x1dTvEqzZzMFcVs3mCyVQWVl44YTDAFj13Dnlo2AzEgFGKMH/u3+c0tAc
NppjVX+VvNWejf3pwCcho4ps6ql82FUILR9HXy1yRWUQOSrtLhtU7oekbZArXG0p
dX4RqYsZ/YVTyOVGJneWqJIgN8VBvQaL1r6JkGOpBFUDErPyHduK0BJLQ85eVDt8
VhvVzfGYYKBUklZ4YD9wsObthEn2+KWHAVTV9xtN/rMSjA1SD56ebDIdJ9G3IZSp
tH0C4TMo9t6MgQ2kCpO2N8tLvazP7rWbIHCLhMTUewIqxQTOqX+VnuedzIwup/8d
SF5nQyyIa77I0M1pycLhva9eBNk4j5fZ+wXQdIKXOBqrKmUhcvXoHHGpgH5+If4X
lX+TAwfxHJmxnvTaq+cYclj++bWWZTU3ZPUUywTL7nj0Jn/lCkYmD/HGmcRKWQ5t
v4lmdIQwqEV6A1BGw/9WZjJRt1ZbcZ0dLYpcwHqJSKKE7Lj25B8rUXiS0bsNrOS9
v48rQieV9NMnWTYdwAFlSBXWoNXAd4M3jE/MO1leROq7aXC48TJOWvwM6xOBfyzJ
GvEQBG+RCIyvjCUMh+jmKMeW6cadDxpArBbyXuGM6KIFDhjm5LxabptWxo9NMoCq
mUlsg52SE09uv9JH/2fCQmqsgU1COy02KRFjwRkM8nYTIzuxTwGXlSXkClt53MN1
qSm5sk7xcADgPGbEwZALZjawlrJQzolAF8qHdwa47Vnhpnvu7xl3btd+KFoLBfBj
mI+ZAxXkYfEHF8c3mGFPtWZS0PH0pJBJmWewkuF7laUi7njwDZwESpsh+U4po55D
yV9lxB2RuFt5RNV3rjGR8g821HYbFzdHPb9ygWhBhuCDEkFmSZOxktHSwMYaVes2
VsUMx+6PAqg5He0+uJO2nUOZtexgsznS3YkIV3Qj5dBa5l5oZ6OAbeVxyu7fMF2a
/l/I9sOUHiLBeTxSbZbitDkxuKn11DtVts49mTiFYp0F/asKgqlhX+Ek0mvBqLYj
NO49s+yh7maFg9V5joyTXOwxsmG0yPD5Zv2xMng3doVEYYXdlpL+HcM0TIU0U/FD
pcbqnBtjUiksGSkFSPtzhgo6kJrdQeT0MKc8TNbogEDGdAnwxUGZIZxKo9eOUfII
0wlAn7Iu8qwpTnJl2p22279Yj6IpPKwCZ6PPZcWAtDbk2UfjfkjV9rbJIktmID6i
ApEdqJ8JgM+bvF21ysm9QraQhhMM3FsQcv7oPTjIAnzBcJ9ygU74A2fSNQU5aMd6
IJqkIhWoNxFQc0QH3+1VKVNHLqxmIWKEVUIC/L2uQQFGHFOD2utDNCJ4NQ0mdC7p
lCNszxn+5wEF1MQnxe5q3l5urVzxzcj/MvFTh8HevrQC4K2xOmndKm9Tzl+iW2mj
1zXOy6KrUYc+JQVQSZ4lM1m53C1RhmoJkBbfxyrSI0Jft1GqOl3kKSsOtafOu2lU
OMxeGDyxKAkWfd83IvGf6ksk8lzz1m2no7OkNc+q87fDiZr8jFbPej8CSHCahFSW
AOsPyDrRvKko1VuaaX/P8hmPUqXCti+PpA45oLWAZtxVE4r2/H/8efdhN+oM6KeY
3Vb/Q2zkFn1nsH1IohoDJ8yJFwqpUGSjC+lR/woXxZ2iHQowpEx4ytzntHgG+5+k
qFON3M0Bv7KvhEqtxAfLxVEO9uSbKN1/T/dDWj8kfIpd4/OLuIvD3JUugzhMFhcf
MTIw3bQB/ceGhUhJrHWMy9jr8HX5qO293eV8OPaMQnyP6Muf2Y3/SD795Xrl3z+e
xmp3T9/rrvG2AwK/EpqeCiZilZL+vk4t8K93LO0zIRh5Hzn3l3jrdvXfCEyxLV8T
HAcDXXaZZbNhaYLxxWbrMeMNGqAEeukfjuYZJRZ7dC0BvcO4XUaaJnU3Z9TYcbS/
PBc11qTWRQhoSWCrcIWQWwiRofNtmZEiGXbfV74GrvIMyeL/INa+SN1EMVOOnE8p
G9yjuFljivqUyLDwOxu4zRY6oIfknPSkDP1E/yZzrFj9Ozkh+ys+HYN9u5hcJI8S
ykEdmpHxTZwHTz0tklCsOwdiguIL/05WldgOQyi+lqJqBKxisCEE13rCVzqeR1wM
IVSrkTsihHTkhrHL9st9Oo6LY74g7NKEz34S/qaj+F3dLKPRjt625gs9OjK8kRXU
XyzU2zCZ5sc+ZPNlwUi+YZ6frcj+yHqmHXku4dyk6pN8x1M55t/FPjCmlImxWqKY
nEa7etN5PxmJr/d5MShDDuatpKLXAxr+ybmVw7tNwRPk5BUOMAsIuyrLmp0a21IN
K97ZaIACbUJicHb4+QVkbXd/z9uJGJXL+BbTlXOyolWv42zjVP1o4RLTNfKs3ifL
E73+5IMOAwE2MBrQFssk4LkdN8o07r36L4HQ05ZJzXGI2PBIsoYd5pxz0yGiMZgX
JFptAXy1WZji7r38RsNwdKVsbJw+7pwqBUTRuJZqIrMt19KW6z1uNfCEws9C0ovf
Dwq3qpu4pb8aadH4+RyALcfq8+ZLAWnlIDpdR0znXUTWoi099AIeFHnf4hHOyiTW
VEQvg7i3rTlKq0B1K4cZLYHIgCpHXUH4IukBCJ544dpOXfBJAJLNfnTQYvFabJRV
wOW3QVr5c44wrxDjJYetVHxrs8HzIVjOix5smi2/veKWtzU2zgKARtDHKB584w0g
vcu8ywMTek3dzaijuQy75paLUJx04/HBv2x6JokmD3qEREbCbaXYPCtuKeLcr4q9
RqzScO+DQdM9MV2j68c1hIOkkbgvsDWrtl/0G3Zjq+Y9toPwF556wb1SGd42zJSL
rxxNqiRRk906+XvLylpIImJ2f1/uWM/Ux7JclDIe70lTK+IR1KySt7ZibE5xu+Ko
QtDcw5Hm1Z3JXU3XtZgLHCZ3/Gacmgv7zbY4lqJ1S5okAhnXY39TuYp7bsjOAK6Z
pAbgepuTPnxXLaKJziTOPnjTeT3CT6Sflnmu4hCP9KlmC84cxoQK2n6nvjhMiVvC
aWPb3pXx0sQ7eciqVi5+YBAuoo8bSWN4n4EO0OturnpYHoVVg5qu16j8oMvyu8HM
WUxrc6oXuwJUdjMkYh8MkSEjgPgSDBa0C+mLb71wWy++Tl5x6iXkS1vb7nEdTdcO
ezXBr0ub8JWpLVWjV7HwylHNE0obeRM0KAf6JF/OjxRn900nazPj5eEdId8Il+OT
MViSdUpMuOf5/cLQUIuhiaOkA5ayb5jUQf/mVt4gQnXdgazgpHFBHT5cYh5nN2iL
6VO8Pn/sSxabAINXc1k080UClQUzmX57THWwKK3V+Pfru11qQmiiHRWP92zZ4B6C
jGSxr4pR/nG7q1CvdAMJU+amC/uxh26KHN6EN+lzmEUB9wm4kFGrrb2W/vMphhy8
/JOIYwn89jlNUEIHn176/3G2rhLTvQptwQ63t1urP+HmUXZHK8jS3c9WLqld9jof
TiEjpKKxYZO2iIkhJ/p62UIiNZ8SyM4QRL2m9+vsAJm8xwvT/5Z3Wu4G5tR4+MiK
lIuMhQivvlgX3rgPLyycCOSMsqzalBFrM6+vHcTubT3hJv6J47diUjA0uCZh8uG6
VakiSpjPEDkAIwB6/H0VLpw/m7OtKkMrPEpbTJamxvL7r1jOG0Mr6OFadzuDp+sk
j5A/37I7H3ueY6f1er/IWXp4UooEjUOXnN08+E9DchyjlsjO9iCqb8GMqTzCfU01
j96q77MP+D5DJoxT4EXFmu06i/0EpsoFzEPuTOHPLr/nRYU+J1liMNEZ54JNksfY
q+Z5gj/U2UTYILKs6/rTG9/5r3liRIN8Hk3lFCcqQ0QaMtxA2JYuasoWSHCAbyp2
0n5FiNyg9VdHgQ8yJZKY8evry5vEn8YpXa8pusXcHZGuZCenrcEorjR5sbB+EGpV
aTpoda2ghRK/uSrOc+kyR7F7kTlIlbCX8Ig0+zN4TMhe2RfIcuP5Uk4g/7MgNM8S
X0qabXXPO0OLeUTwsEdntgkSJ4fuPoS7u/70H3Zt+Tg4p/iAUhX7jJvV/Wehb6PA
4HKGImVhTcvb9ouHdWMr+L3bW1+2FMq5HuKxBE13bW1LFPJs2WR6J3mUL9MU/p4m
WYqLSTulfL6ecxKk/c2pJxVTCKaocX+nG75aobcauEFzn8xJfR2Z2bCsBk009Haa
ng2QgRv7D3tk7Kd3wEY0wF8wWhJXBO41GyxakhamJc/ILXdSKGh78c4m+5A5EtsQ
IXpKWjjBrfibQwa0bdAU4Oh21OTT5Z1WaR9EFxEt6dtzvSMnfhJ/1BRB6mE+drNv
btOCYlrh2BiJPNaRNIKGLAXDYyoC25JuWKrbH9YEoLksPEFg7jc6wfsz4x+SpG33
ijuVVb1L2cR/q014hI52p1kDRpKTXDqSMm3E2wBXauOiIUGFUqW8BjVUyn3IZtMt
8ZOvgeZ+NopDJ6/fQNTGQ745Wdt/gIt8zCP6C6EzmFoB+VoN77WLkHSovr1D6KO4
pbEU7PuWzrABqG1Qqc8PB1d80EHKi/Zfe4MUVT7fN1+ioFKTnjXixQO7C/HFJY+b
a6wSuO1UgfU5+YN+bZWJ7eIo6KrfGc4UWOAbTPduFVWTmvzQlP2YWVVQaAEWz2s/
3NwMMlBUiQHotTR51+tPShdAMJ0bFfmu/RPQ5IeDUu0PZDOzUHmW7Kp3wZQ0Rot5
l71vqE/pBDVFua4Lzmm/wr25+o3ZkuYpJ525oxemhWyAwmeKo9p1wDiRXvMAiR/n
6vSD4nuuuUVZ5o2F7+eaWKWjTk2ojRcYtS7LaC8dNBkRq/hyK9QXCpuvPsDbFFfl
2pLFNUU+po7VMkRXbyGyaMg+XtQJ4mDQm5GDCVNP9VUZ9OgK8bfmFKGtqS0/nwls
aso6nNoXFJgNA5qVr004wWw2I8OV8PtM64v6YY97CVhJyd+kMJJGP78rMtp9Exma
hjSSeb/YWGibl5mLwRkk/wdv+/hWvFAgO8XbQ+cBwoa/pw2UHGqgq0/ctspvpxhg
bXrHIT1xqfpdCV8Z8ljYlbubjvfcARrvWAt9gk6ijLjgZbdEDP03eN9243CxLGmT
1qlf7iq/ukzRWrIbA4VM4r0lbXeZ5zH5uBAMTGM5QSw2C9uFaPXJihVPV39NGtjq
rPDm4bgNcZer+7aO2t9vUn/QCBLulfE09YEPlPgnj8W1tfKUFyVc5rTrXJ5y6A4z
pNlFst/ooJLpeGh81uytkvaDJKaMP7bJgrv+CKcipFX+kBT7ZNdAnmsII1mZR7uN
1cf57UwmEcsTyrwGuyoIs7QPVjIYkFC95IqBwPzQ5NS5Mv7E33sDKCywaGE8/NZi
fsOBoQRsQ0imPGH/iMRpDuqgqppy+fF4hJY1MPw1cHBA+Kx695U0S420CcZhdnyi
l5ubjOYh1fpNpN4ZXEjeUEgYd/qkWmUqn4EeBqNgW8oo+Q610tTk7tWIwc5qYzlf
3osVr3Mi+PCnU7nQbP/YecQkxT2Xpa8TYinRSrFVcx53724b3Fr8ek/YVmUYmup7
EJDbqR8T544Of61HQc0ZbWv019J1RoplxO2zA2RFWdGrEt1mkWpbmYEZU3h8xNue
cfWXSs1QTznIopRqD/lQgzuAkZp5vu2JtSbKPS6JNaQi0n3Ke0K/eQctxNRK1WmL
P04SN5YL2ibDE1hKeS9rnKY1ZKFeqm0GNiI5f4nZPz50UABqpp8txeIvvz6uQ4Vo
tYifM2PXqQCouWTGnsl8Lv4k/SNFc6bX4m9eIIrD1kk3Fb/pyopbE5Ca8bM7tohA
+CvidB3IRCSZ5gJ8lAtoj4Sli7IoPznLK7T7qcOqT8TmWO+COCkxkZpYLjWIO2sl
iMW+KMQ7bwwTpx5xcocFTkn/nC3JjHQVgVOwFfh5CxneHHyX/Y+0iY2nEYF3s4dx
VDGExqmTHMVJ3rATsFN66lRR3GoOrP94ZRbcg1WhVB7E2pMNqum8bFHRCdsgrNfD
9fKjH2LJpb9CLk1CZY1MeXBoWNyzjT6inmjYcYVF7+ghEJBEC4+tS6UQZEDiK8MN
GoD4MFcTXaQY4gpBPFSzFXG/SVrFf/NIFjrM0NjSat41sGITaDu3jw6x1b+5j65q
VYJe+VD83rdVlyWnSAebjpTYXwP5ga6xOSaIjk03K/CkcqHi8Tf1G9h9+IOxMMlV
GxaZIWw3eoV7MJRbAAHJDJMYgXIvY3aeIQsj10PEhtjxOvpo50I+2a60wt0Nrrei
W4/3aW+EKwU0QufJX5mnDoeRjhoIff+3mWTzkOeTyhMW6Xz2W/CWIlEyfDnGLXwR
EH8ivZ+9v8tUAMFVsA/jRIKGyxZ90S3Zc5yVs7TbqLoBfv1Ti36MIOgzAMAxaUgT
cZ5E0FHTHPaUeROdcXCbSlZEGBsHHVGWwui1/jmLY0SjGntOTGIq/Ozw4ZVZUSXg
87UPyyanB0jyObdbexZmAlE7kj7ENB109mPm2biAq0tQlaTUOakNx9+iqTMiNYEX
L3+hSY+aztKdgPs39+/tG9tUUpQEq4hWxMt0hIg9ZS7HDN+sv9mv+FCiZeMZzUUR
FcesriAF96wdgmXKAKheMVeL4yzf2F1SwjTcH8Kb5c9gdVK7urVt8+q5kStKCYYi
uOQVhJOQU7uUtfPm7czGwpPF8Udg9EIQFF5s+ILG8DrtYZ9x5b1gYTWvqpEhkHt+
0WgR1UysdlP4bEA/+mZ/xbJMlWj40dps8Xx55I8/8FBwU70/7lvrmV34shFhESxn
AUAnYVk6RMLR1lZKxew1uuHVMEXTHehT46WvtaUJ5sYpopbiknJdWwY3gWZdcvK6
1C+5nEY/PT+jdNAQE4v6TibQ29goXlmsS+n6SmrRWQcxs1u3LvxnFK5ybRR01wMo
8w1AqN4FlsNyZztYi50tO51CUKH79drQ9xWtSD5k5mxOgU4ittJmHOfnCp9kjoeK
cOuITADLlOPjTp1jc+eowK698O3alhvWcXFc5w4OLvOzc08HEutaBuibKgI0bqdw
Ff3W+WIrjk+YuNuIK/32pR4w4eK4Q9G8g3E+IJxaULfVafEcJi9cSOxtlO5Z7ict
93Q6+CEW2/vNq+VQiX9uwy2sEg+lC7GZ2Ffa8tnQ/4tfnHkdmwvMQU+17hW0+Ien
9pjgJiipd5Hj+mBhzXcZNVDXGIZF+tf910uNAKKtDCggSct+1SgaYlTctyuYd3+a
5QbZKfLgVfjLWb3NwHHVP1frY9m0IYYgNCYTKTcdKdwvIcilMjfJ3H5LlojoDVSW
LtzlKm804Xo12s/ank3KoupsBe5jyub25p7fudkdd3mFYX2FP/TDpeFJFmRM6Z5Y
aOH7KVLLtCqknv0AHyDLuqYxR/SJHwzz36MLGF2mST11hvZG1ae5RSl3dm6ASeWJ
jE/Y8gSN2mxbPh+Bc2OBtvnjfRHZ8/qkwKFxvf+xVaPRR8pa7awixBYBKlles0la
wDgomFrGpM5tWN7aYtdXt1RvBqV/6Pmy9lQKSM/mgCeszu84rKLPSjDBWqG4DQw/
NZW1fbaWob0fj9g9mvkHLdKbkKT3tXtyz4XTNMo+bL3VTuEXB95iMJ7pLibwmIX9
eQSSHu2r6TjjIQ/f/5bsJunKLGouzgVn3nmMSndIFuRIwwu9za/HBBnD1pauaOaS
tpRCKwpH99BagHlg4uJIeQW9S/gjXkS3teqxNuOaD+XjG1r0K1eDSfvuneT48dvy
i1Ua63SMZWA03ZbvB8IxEZUelQ5RUF0UvEOaxR2WdRa3nxyuoMEOtH8QA4mpFr+e
rXgIGMpy1noJvxJ4ptb8JTtho1XRcK7vGBgaOuxCJj6t9GuwBlz687YIuHS92B76
NzbeMvL090qbX7FKf+sD0TVl1nIPhe3ZIL0ooGuzJL54NVBfBWWEmllPSlOVogVw
ePgdADq5yhrGR9otXoRdYdX4RadwvIVmx6GX4EPIOBS+H+xeX+z9X3cD+ANeuxVQ
aulbZzeXd4em4M7PqVXjatiRS5Ohvtahkht0m7WM69ieBdWNzI0p0uIEPYYxnfpe
gVH5DDmZI8W0npFwKr3OjfN+lnv0HGofrc2NUF1CQ7N9ThscEnLYWcwdfKPbBRcL
WJDA/n+p7MCnMwZ9fYeHJtRXKcPVueOhQ2RThwVSZiMYlOzlHbBaPrN/hlo05Vaa
3RqWRHOLXxtZakiQE3INyEE2TZM0wL6Wb07OcvMtTYZQUHF8yy/wLIeJr697q4IT
527LEjZiIkJVn5HONdrv/dxqBmxKm0y3SIM5DJu8LhPBHkGW2o3LwwBBXRJmuE4x
NdQDrh2DUT1O4My9IgcCWUk/uZmH8PRJTldrAeWhSV/g07in1yCKcCzgP67kIGgb
+FjnB5qU/LJKcv9AkvAJsKv3zFMh3oeinusXwiYR9YSfJzPTDh8+ZZ8zNrP6D8Cp
lcYhV7e1eTxjRlVHxN/5VccISuiH5oHpwEt2gKcxb5Rn6vdGUd8T7ABu2Oklzsh8
GuPON2K4IZ6cM6+/JrYyRMSBYIL43ccF+1OziBS2YM90MgSgz1uy0FKBKhnsPrMT
1EdRJ79uEB2zo3MBOgGTQH12Mfj6/iazalv45TP1jcdAJEHVia9PeYqpzuh/8Y5R
pgKAXy98PdF3EixjsuPbgvFLUmx5o7nRmxsXQfhgkNtC2dwohfFwWCIp2CL4bunX
9qhSHyM/fRxa3p6/3ddyoMzuiKXfeptWOdOUW30oYyTZMJL9pmkt75wap6QSraDv
FhK43oJ2BaC2yBfkTtDa4FzKWRCb2kYAikufWO3RhY6LLTP3BbAZiBG/8Ip0USD/
BjLPDkImFnKasVp2DANBgAyDLXwCUwHv1lVfugw+oyqNbMNKJJRTCZuqTYRJArCe
JebyEruYs4FIn10a5eDXF02XEKV72hTGZDgs88OcNRksG7p0gXa8B3Z3lAcWJyIW
Lb1asPGA/c7AfKaT7yN7CkkJHwAZM9Nu/gjeUPlI1VRGRe+DFEAjDo0GNnFsqR2c
sIfJIbcSHmGiwxnIpCz10CNahFKVxXKXxD0UuNHCjMvFOGMnoTGqbh0iKL51I7D/
kwWwFU3a1o08agBNuem3UHdEJ/jwrunhxkxY15/knPW5AILDJFdV2jf6yl187Vgk
8a7Q7jwB+KI3WOHzThaqJTBgvCnt6+DYh+1OJqu5w7TcmtLz778KNeA4LM1tYgYd
AijPrVRKQMfmhi4k06QBkhy/604+A1wR3c0FsH3DDO048hqg+KxACkj/0I/mPazZ
HI7IpjLoBPF5DQ1wZrlGlFmY8/CGgAqVbbc8IBlF4PxGcmz780u61JfO+30SDgVr
mxpzMx4cmcbItFVd5T3laA/mCHUv4maopejbo1XcInerH7F3cNw7wNXJfdCHyvSe
UHnts01I9XWa5qXVEf9862la1Ro7wUajf5qEBUtLFX2lHZ3fV78ObmqRWQm7CQoU
3rCMTW80wy3xiVaXWJhv/xaJP0bPhUy/pS/tMZ78mpq6PfdmlEywZ7BY/EngWObJ
8BVGZnev5gAZqjc43MlwgPl+wEdABiGtHrzDBWfjMLAU8XtgB74YtfSdgojfQ9E0
KuMTtoRT1uHyq5eXeCtEE2HAd8kFSB7sAq/54T7GqERNAqm1Lz1txNgBkRqZBtO+
fqM07mUw+PtCuCE0/4fGEoDcEZS8rx+AWDW9Da3Mz8ErpOLdsXxbDp7hIbmuQGlZ
nQT69Jewv9HXpArtSRyPMneRdMeEIZTAnXTk/KFCiSGeSbeuFzfjHo0sBqk3u69L
v05tSiaxBC/dbVqD+lgU7baU6PislhCtTuHM5HN7Izm+oagj0LVzctvJh+c2tzsc
4l7Np4gP0LDboqPeqL08uTOIA2yOnQ6yIh1Ma8cKhWXHP35e82haJ0B33qTtbWfd
q4iQRDAY+YdmXW/VZ1v6mFVdJeeh/jFMbDzwhsH0oJdTAUSvk4pTWENmbY++3+ny
FJLc18ZBclBwe1s2Roa1pYcclAEUkEE8ZRLJDj5MfIfBWVtYnIWJ7PiwswL28yQW
iuUE8E2L2L3YlW+qsdM3j4xOR1e5SXp3UoyPQB7F9vJEvgaxJh2xbqUkvGSAdrSB
R5lxr8dPuhM2mmTj4vggK0o3QJBs/medYk/k18vLQQ/5FF2DmgJXbmTI3ErDIGtP
fIEW4nnCniqA4F4/Gjb7C5MmG3YV1oPcU3/C9AxQxx34f3GE7g3kNOxaw/1dfVtr
OXr2WF86UEPsiD6ubU1bypOz7mU3ASXvTFqLzaRwdmJ1hqSmiO3Y64Fh2/9LODg2
oP6437BGG/7fWG3mMcuJ4dQspiCkvCs03kHFP5ykGB0qyljmg1F2iSxYwE92QTWu
t3WVSV6Qb5LKzIV0hJsa9bLWWjjfbz1KfOgO3ivVvdcxQ7Q7heXp81DADnIxg7Cf
1tNJuTwHWy+8bfwKUc6cK94pFDU5Tv1l9Cqd8ifFTKj6nJRNyOS9+bRtfJQ5WMCZ
RfwG+iXuRjRBVfpqQje4+yONyjSleX2M/M86pr4Ec5rx/4AXxYK8v5SEkLGQpCyx
MvStdNoYzZg31V7DaYzlrwLgylvVRb603FXkw5GuiV2EvjiHrN4g0/Hekz/wW0Yi
oDY6o38I10h8jrZfFCdNua++we3XVw+V0V30cSI7314LCHhltx1/gl82K7WApYKU
/YzLAlDhgP288ZrYZgrvVnDKm+RD4o3xf0M0vrWphwag9wcI9inL2WopyN9bpOSa
XwOcFqtNBqjmTibjoS1WfsL/zfyu+NC7+zlRSri+2Z6ZtNYqnH2bXh5aVSB5yS+x
UGvEr99tqQhuRdcf61RuGNvEi9HAqsb/dCLl+UmCyH2mT7Er8xku1V7a0AGW+N5z
S9rJly+svuWcdSzfUhpkizEKeDZqfRHOiKvZtfSximnClYG/BDWfvAVa566rVIqD
80BZ2Tzl1aDgl+Sw7SCBiYoXAcvN8Omwg1sxuxDEaO1xgMacp7SfAtTCTDpwnTMz
BDPh1wnjyslMyu1GVrW8lDDhEGTN/tQs461qm93VoobOLJXAPdMKb7hx3sPE5rtN
6u7xh4wVcyCg7qcgjT/ow17WRh1wSi14KVgaGsun1DpnwLsTII+F5Bih6GPTWYuM
y9DuSWRXbix2TqLueOVHgI5hPQdi4hOnMePTapCkoRrG1WfDm692B/mZB554GnZI
QZSzy8kh+dpRj60s1fOwLSLiQIyfwVX3mWrinDn9+HOOz92JYu2V8b2mgXqbLxrI
WJpTsV2hlVsPD1Rg/B46KPuPpGaWEGjkL/K4LdadZOSLpRRIH+t+KRqoYPN2p0Qu
0un6s1cXi6T1dsUe+3LF8sluh2co6ysR9i1C/EvBFscaWzbSp/jZtAlXJ8AEPwB7
4d8UCcvDom8EUysJ8ZnlqQQMTLQckPBIO7gx+rLAweKUdCVf2LFHxfH48UNGzToH
Yn4VqedHsychH5zznljJPfgFsSdhCQyW8mvCjg+vh7+94k2hDHWbeOVz8lBPSVqp
e0Z1m9j3GEZMNVEBhSRFArVvVfB+sWPOYMVCDJaIDFMsllcWEEgQcd3XIDvGf+e8
ILJCVxA8NHi9kjV0SFVNROnlCdWGiGchPOBqqih0uSQpi6BQaAhevCEZGg22ZOYj
9yWLZlc+tTcUSZzSqmteZgrIWWVdJmdNOQksxVnWcKx7CDNcYFygOc1kk/algc4X
0SmHHx+BMirBIJDR/nS0/qjLpIjibNGdFTeRFWEQd+J/lditC2NUeg+ZieUJXGW1
FhN8MclW2PEBtUcs2Mxei5xs/U6MOuH0EZ6DamPGZWj6o0bS3kal0sczjKF/kwV1
m9S0LKZU/1sYXPonhUAYvODowAj5tK7CH7UWGeeLjNapekRr1AhdOAScyI29BCFi
u/hzDQuc0s5n7Yr2ehOF4uBhh2L+IonELmCXahPnrxxoC93YMi4ggtAOOiLhNJ3U
r5SHn0TvXB6dtBdLpqy5AJMNzv0ef6aiMGk9qxIfuIkSwXW3VA8MdEuCkWOABykh
Pv/a78F7ORBkojhFydqH8V7xys4ADSLIH7O6gzV4JqbwRNQmlI5cmYNbcI8pyt4x
xL9xevIxbR/KIqivQehMYVtkyxQSG9IKygRdGbDreBu6+uclUT6vddgwzVNHj+N6
XG44865LDLhZvzF1saz7/Bc35OLp1wK79FIk/z9GI92786YW1lFknNAH5c4Nfcmb
aOPLk66bcua6sECNcp85ZTT/sfFPkDgkBowIpGTyUgDXQY7eQCPVeH9yx/V27Atw
IPeeN7BCGBazg4Q9tw0c7w2n35oOvQhW/sv3kVYSthLzzMVePN6dXqxXsmKFkEas
bHIRuRqR4Qrn9IOyS1IMgl1+zetrF33/RrvWj5EQPb7CGkybVkwwLgeKLcxGKxdd
KGOxTMYPugxZxp1jiLisA1BQkmRTRCx/e5XLCdMCTBMLP++rl0mxlsreL9k6m+bf
NGsoQXAKYizCpDUySzEWZ0+8fDp2p5PNYJl18mJa++c3wuDkOZRplRFRlqSOxMsU
kmpsRjnSBztmGbC4ePvmj+Z73AzYNy+8JD4WB6MKOIKwlne1r8MmaSRXVL43x+m3
AIeuPAi73ppLgBQip74gKKFRtlNmj8cldFJhtwlBWyGx0POlOsPHFcI55ZEwbQSD
RYS/tDMMSz8RMYcw4M0KkEke/dHdhmZaPJ9mvLKUiITbDgDSHbdkYAgg926tPVpE
y5K8xKH+BQN2Gy17M37Yq0Xj00wY3vWkuypyMA+G3urPffm9RHI5TYrEJUyXje2T
OZGpgxZn2Q30itVQRsCifaIY49jj4N8EchNjLB6QpJl2LFo2CiPDcxxhVq/NKf04
DGCb3Nf0mm+noRnYfQKGTDRbVM5b4wT5PL2aAtZSJUvwk457/JCXlCenV6rke6Uv
N6PCn19VjntEAiZjj2a1ABFd2uWgC1VZLDj8TC76mUlAHJhkrvtE4ydV7qpYQQPf
9UPliwQCg0LzLyvAdIRvSSgfVmTb5S6ZZ2paRyp4H+Zzd5wc8eZtQj6hes3FaELV
vmXREQo/Sc1Ud4uLlLLaBuohTKtxvPYSd0oQKdrs8rm1eYWvgaQ41RjUT9/xO8Rh
i7+72ta2SECB7WEGBT8/JyPWjzEAG78uUXiHFwC2Z6Kc32U73zfKoV4+l+Mu0Ri2
n9ku0em9j92EtvVlcYpafgiGxmO/90ScuDIozbpNAgf8eEQVreK0F5qEMvt0SKNj
qJcrP2feR8troHl44SJWP83n6BakLX5pbwJ4971N+5C7DxRssJ3w05Pb3j8o7aKe
EOaNc5a4T9z9bSQS1bIYbHu0P5FD1fun/i6sDNxA6skGJSOJoKIxePNotcPfg/QL
vd7X1IaUS+HNCuUcQx8IurjwLe8YUcRq7YkiihVhwFsXX4vL0u8ThyCUmnUydxmz
uYCUtsCwHzXIyNFRymu9SFkXpcmq2w/zOp0p3vXhDQVUVloDJ/dvs2eQ1nG0TOpL
8TwBYqLJQB9Q5hXqtWIt+GLAZTilklXlLprP/mmAPfKTgYlmuQN8GnhMkJE7H6Ea
6d3RvXkSFmvl3QjbJRUskL0WI08O1O8CUWDNnbmxzR0heALJSd4O/1p+CLzcs5Qo
AQh2zAaKul2Df3QnRmeNhmj9XfViXnpr4pFMAlUnWT33W/gX+S4YQRfWjU+k5ral
ZhCshbs120a7YdbopGzeWyLx+5rprFM6JLFTvja7QPm/AhubqvVLnNUSR+UUpUNV
gxJJ18Trvv83nC0TzwuZ/70z5S1FlEJIOo1CaXUK6vhy0PSJUovkXpDjt4EfNkaW
VJYQU98ykVsicf0x9kkxLyZdfYLLtgk3Y8OwvhUyPj9BKRwb6+9CFwUrhAoptoZT
n0be2UwKvhQIiioOzDy9rmI5nT/CmHxyaUC2H6zNlDlO8c8VM8rkMdhXBUu3vcH3
yDKHLSkCdYwlTm9aqo0ULi+jIEqTZG7CexnGJMMEbiLSRcJ8zVlMR/hUf1C7omFK
UP+zradkeF7PFKnU1YmfJsl+C2jN/HHcFXebvFWbYOawCIM/Mvgcw3ie7t6zszT0
ol3p5FBEFZEakB/48j9xx80BH6a+t8c2420uTsIRTgRItjpC6xgE2jDiQdXvAxrv
AFJcJmkTuwmetJH19hucI9vxUpS7CsKHvZ2m6MrCbdsv0wqguadK4iQPaSOrTfRg
yUlnr4sodT1LtEDA84BRwCEWSEG+SrCuAmihrmVvDBgw51ZTz5xDGEqaVoj+gltJ
CnNAodSaNiNyOqEVAd4DZyDdVG6vXUQLBjPH2W7hLJNL4bbQuKjBLqyv9eHVdDCG
UpgRdzBhRPEBP8kDrAF80zJLWk+Jak4St0uqoYV3SnW+unn/0OKrFV7D/cn84taI
x5gwD1WhUS/MuCvkP8LnNZbSX5x+Ae4jlbIrplWUDeXWoG2jaQayU1l63Nwa7NER
fZQcQDZFwHRhGIH6tY0/vHZAyK3FEkKg7jq9kcO63I2T5QFw2blPuy7Toh7PD+UA
WBhYV+C1HXrJl7n3pLj34NJk6VDXh6kws3jzcl1dD2hGKzMI0ZW2yG1OIeiyre4N
zmE2Yw4j7UrHuH+E7FOwfEsELTf3cr59v9poByGhxS5FekOFkxB+q8dlqEpF71Ki
7AytJthX5Z2h2O7X8UTS4iMdKDme66haFmyo2i6asCYparmOmeDoN6eLw4KcN04R
dUyNS+6Cx2XEMbJ+ZOqoOCc7tYDsCP/Ta0rY50+0vmfj+qPqamU8RTLaNcyfVqK9
jrhXufOxKNZqeejOokQLYYEab+k+xDrdX/fYsaGFEr5FMxtemVxLMpReY3mU1mnA
byQNGnqn1FORd19DoOBDZoXCHgA/WYm/QxSwexTz8a4ondQqu+taP9mfj2/cS8ZA
5qXDOuCMpBghrKerxve2tn80HQZevqypARfgBBJKT5GzIJI4Pf2UPdlOoDfxqB+T
gKvwir8GFxDChoqWabfvDoSSMBCqsi6oyLVxcZJVW5fu0gbHKIfTdoxW5fxZPwjB
K3dcQgH+VYwC+ICaoLuqrU/DnyvFuea5QeSfvmbyoVii0v+iMHPVSxQT5Y/DmT2s
hGfTI1sbIReQt14lMos66hSLVoA11PneWms04r1siHWbc3DNTKuGG5AKSHN330QS
0SGFVLII11/4m+JX1iOseWYmccOslUVtohLlxpHWFWwlsizl3n7jva+UEc0yHU5Y
DjJdXmcJQmtGfWWCFGl/Ieof1V0X7eag/qsJlHQJbul//vNGNB40ahxSwv4uZaQc
ryG2ImKL4bXyY4L0wCCt1OeCnXPpYDHpQhfT7BSzdGxUcqNrTNElbTLq9adEkOlj
Pjnsx8c1UCYAzLBFDYKeotLnOTXuAPJ6CZcqeUta9F99j5T42Mieg74vIGCfYhvF
RqWj+i2awwuT4R6nI7Xr5lYf93y8d//sC+oJ5X5ype2CB+1KdbvjDSauXGPS2wVd
iOFii+PWfLCjB5SdZMjIFi3xZs5mpzLfrL8uuswjPAyZitzh0KN8EWurt3PjyP7b
bMqeOlxAXGLcLbWUnqGF7OwPf2LZofr41W30g1RXw+jFYa5XHIccqV181W0nw52x
X9gKCKr8zwh5MAspN/26oBgzf6EpdoTK1q4/gPTm53wVb+U2SeufD6jUvVxfC4at
DfKuXlQoZRedOQTwGK6lj4h0pZpNX1qk3Xe3tr79+9FbKwvWNlGUuxHoaxU4GGBt
CzPZs1IW8nb7CaJuZmNhbM5gWw37QB1xlizzKRUmneNQ7VvZkYwLsXWfR+67/KhA
o0ZkA34ZESC4bv781UR2rj07IwSeQq7FbWCXsbYvc3Yyf9pGABFOxrAJ/eGM+LDQ
eaCq8N9ukOseaWcWDOezmUqPs55PfHWDVR/rDTp306H+C7TgYwZw7L4+tZ93X/Hw
G5Wj9Iq6OrokbUVnZ1L3KvNJKiIKo0RXazU4BA55rFacyuuD962PXm+5QnsBoj5K
6NjyEdbgyRp79vmSzsIZo90rA9g/mAMLblPvVTJs8B4M9ZHee5N4YDYkEDe+0jZo
WEH2AwbPckGq+XmUWBjK4RvZIHWizDNwOTKuHLeJXM0663IY10jmkm1jIcPnkjRP
LPiMxp9yWVmDMBn7x3g9uLizjHdYE7ql32SMwQeDbJizgF59GbRWFJMDj48j973X
TlDQNou70kO+CMvv8eeiWr1DJn24s4dzffepTtNZiCi5L0MNhkhgKAm5pn1uCU/X
YLb+FqD5H0yCWM4u6ZKW4IJaTnwqBwWKzjRjLyKFmvbwidS8OCV1+aL8k1VK5CHS
HIJTlLNhbgCU4idTYVuxBu3QijlwcIgzElg3qhiKSsknNep50lh9k7ZMJ3JGvpY2
D9OKbn6cFlIYUKf2JTkzO3Bds+P1b48c28KCjGvbheu4gKz5rkh/IsD79gb5+9MC
/Lvt7fH2aKnxUuisZyR0gv9tPd93VfkUs4whSUO2w0a77U8PmzFg8Ld/k2AuxkjI
a9GoaBG1im+Hy5V9HEScYNXLPGxeZ5j5KLaZX2YE7JL9I8ExNuICPYyYjyXQIV58
XiNWyJx8QvJ5zdjdMs8zda+mijM+60L5s/rvHPv/mSOF/H7duPZChjZFHXiCSBCi
hOcV3216PD0VlZoXYGGTtKtHT1zfMckGCJURUy8thzXxT6Iw1wtP2RqWe1NqRyiv
5S8dvyvT84ViGsdnRpXN8fzM3LMZaNBtIn+QzATAndr+5g++C1mK0eOx0hIxTpKU
mlQ96ikUTKZXvRkOs+cG57BbZx/g6RQ1baYTL28pWCwuwj63p3HprmW4UUu7lsHX
GNFxZ3aqy7FTYgYlhp8/qzOlNrT6o7sksdGOn1rUU+X+Kwk1rnrAp/wKsvHsH6Hj
la7JFrVyV/IOGO6yW68QBsVV5Z0MSNXGCDvR6b8pEvrEu4UIrzT0wueiIy58likU
yJm3KidtNa7W7hdlQ6TP+dl9nrh3S6dKFromgKYQH6jp+A9S74Gw8Z91DmZAPVtP
L+ZlfX9lMbVzYIBzGNTZQSw7ISmgREvswFrN0RZDfyrsPzZmYWTCjW8b+WbGQCPc
Jsoou1+XXO2212bQlfRypoUyp51TAl5sKP9hBE/zDNyB6uD146cvde/jz/THnEpO
KR1aYWMzycStI5p57e9kmaaBYyoY9w6kOvyR5G8EGWNtyInNd8+Wq98vXjB1o9m5
UF7oXWYtVz4brShRSKzHRBDU97zsIOAblojj0EYZIqoDQIqCpuA9ze5FM2x2b5Cd
X2V9qTznso0TvO+9J4EsUyafbRuWTswx/8nKSpEdkmpTh35pZThxqEW5KJneAgRP
UKXvh7+Y9UzxdBKU+nk1O4zgrHw/tZSqFpCZXQPa+MQm9lO4oAdOUq2bJeNNdrmC
A8PFb5KdNhFNarZ3S3THxUooRtxVE/+pCA1X2+mDQQ+MZp/KiaSIZtriYTetv3j5
LDAc72gYbf8eriA7oIK6YEHVlo94So1tlc1qJHObfSyOAgJzDkc5QAmW7tA5EL4D
nzEvl9TqmURVQ5CRxXmbj/L80eB9ghMwOF6nUTrAwjK5XTlvGwnQFKYPCByKmiLn
wZXDRY3jyOMgTaM/gjBcbc+AcspCdUQdKtcylUrrWMdemEsHFPHT4MJJgtZwPqqY
CzCt5ysnXDDimGsW9Aj4kw==
`protect end_protected