`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24224 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
LfLaKOw3utJqtz02pVdKf4GU+gQRae2CP5skAzFs9BAjcoxYWOFxdnDO159qgpCn
IRaENpO2gYmmkGuXGP8J3dWE2g2eS2F/qJp/dvimDvYMS4ZmRsR2GInLlijY+EsP
1sIRzjpEFHTrp5ZJ38Jy9WmBNNffl5zxK++7z35XET9/ClyB6XqXVPpmQEFS3RRC
aYLlvLAZwOG8yXv/fbT9xMkDjK3UWDxptfKjp5FJw6F89HSg7HXFZL7l+LoZ93AR
MjjmHEMYdAXVUoXBR9/4n/SymI1ZePQZThDVramJDDWqkGTRzjbLKAXxlHYHe+KL
0hw+dkVk6RiK7+tBeNvngVGYVALbiL6G0GNeCV+7rlPssHQ5lTLLWEDNp2a3aVlq
AYx81mFJkiIOfB5k5pwjOJGp+h/OhpfguJprOZkzAUxZfwh/E8vszK4JbIr83MQS
18PSFcFy+tHiKRdvppZbx+vYvbxLLYnlwbkW1TdkiXGMhy9Sy1ZxpL/kdi+xIp0B
sRkxopTpguP03EZ4pLKjtMJJrpVJ9N3j1izn8KJzcMbxHHao4NECC5J8ZvRwPMqu
jf73ygCILmls+J79FCrMmNxHu6j48e1xkw3kFkfYis7H6CmWT8msvsKUWgge0Cmq
+B1HWLtzdMqMse4YGMXiggOibVWs+lS9Jym2V81w2yZao9IP7RC4+ri/MPuZeJlk
hoHFZfJnOpnlJI6NHOIsbA0q11L4CDHuhCWJRIzllsGKvOgNMT/vzXUeMf0TwYYg
LrgK9MuZS8BUz0HgnrxgkiBLLlyyuGS8qvr9/4/NFA+jmjQ+DIfZcZY2QeEsQUdx
xJQPUnuxjhwswrYCJIog0QJpqRliRmLGMVelnCpCH6Ui0tyS/TsA1vmQz+KW/QoO
GkmuaWsbrHpWhvc5PSo9U83f9XJl1N+px0n49HZZdAAyKh6Vo4XN7etQNMEpTPGp
FYv4HVH4VT2mCd0G+Td/9armY3tyfCzLjhWsjnTkj3nGLSPnonR7Q5OMyF1S4jZ6
k13ee0u/QsxHD2/OByb2qgUHsnqFDrBDGoNgm/mFvA0AjWris+SN4o8Ylb78U0Ae
yuB09O6qUYNqazolH89v066nm/6jPQfJR3inQb/ZoEKYSHrExKCDfB5hIKE77srL
U7xhkFwMThg6aYyXpjUv75NsUPav86ZfjOoviczqhpfRSM71gZ6d956wnbMZCxgI
4KNjLUqylDj0WSqLzzQY5LtrSQfSdG9i3Qlrsldljl4pI+c43nt8neCbG0VoUOdM
JrBM2BzDqPrhLkQHiIL45y/DVIYr49O/hkzUXtG7dw82ocA3SAdG085YhD+dxLjr
XfOd4Nan1mopaXFWcuBrTlIO69oSb86LsljZHrKzMuMwXD0dtTC1zRh7y4DbGVbc
EZ7JTj3nmXyMXSg+iHS6j/TpivfTBs49J43rIDoHWacTxDWuHoYae7I8UtODizHg
OiDIQsr4OYnctWgKbwDoJqvgeF0joG+uCkxYGUSoa+bNxIGoaTn31lEKwUV3cN35
qjaelAo6WHieteNNd3P0XKnEFgWqKMpZBeXsD6bvBrXC3R4JM9KTkatOExPlr+uM
OaBSuC0WV30bndyD8kp/CpL6eZpayHHafsgdu8qcnOcSN6nlWrss9nWSeiciXGTW
IbfLIH2OcH93PnDTSpraL6SYz+o2zX43ilVzo92MgAXnXhopONDZ3NvK6JO+/nSt
6T+YGPazRHkP2kNXisvFohk4p3+n/kXPm7p8lbWGHiz5jbPx9cEsB1DPF5ZLDXm8
RQsnTHk5rr0zWyWDDKo78CQGwPdH7tx5KoQldY9Ybkuxb+5Us2KagQvwDHL4Z9Ob
DzpsTaZt1fMMhYGXAQaeF0Jhg7GYs0U+mbtdYufJHLCmUTABzYG1kOd6mZlc/LA9
qrJCJkJb0oQMlxXMWHvlEyyzBIKxj5Sfo/9eG/ApLVqVT/HGSJZI2VoZdrq634Wf
8+2FAPBB6tYG+4RnvCO8+mM3W4UOaCLFhYZVaWyWnampFhOcZE8Ld8KATS7Pv7zU
YxzOnmkSNczZBRvO49hoyWpnmhzbgLWR9FRMBeks/AVQa3RXYOIqGYHpf5U7oejO
A3HjKN3zPzNOFNT02GQlclfo7JDyXS9rrP5RLP2X+/X1SOkqpPW+ZIwHfQW8QvDI
cZWfp4bd8swCRBjSKU2yEiKWbL2AHsFUj+zT3pgN+3ZXG76mop64jWux8Tncp2zO
RsfhlSmhSgYzlY3BGGhf8lKiEr7brJzfP2LZEsUxTXFeWRH5Yl01ipOEoPdw4NFw
NWY2iCClsLPc9eRcjBvY6plF41FCyH2Wd5+ieN66muKiReP1ly2hJ7B66laAd5Zm
eW8R3amBF/Ux68xnI5RTNbAirA4WDNh2shXMa4x7DU6Gi4E0Tm/CytRoI39akD/6
h38Xs99a0ekSVLm/OAuve+ai8j9GpOH/riv+SsfZn34+JIzCR+PfUTY7JyEbz2/C
bnUTuXnfT2T7FFXwt4jvDd9EIKYcqSBK++7Mp5A6o6oMXR67vt0DLxYc2OMmY0Ux
Vxfui4dZRFX2f/ziKA+2fkoYOamJwQDUlNFgJdR+IvPf499FLIxFyGGd0JzY8zzi
nbFMtzAaaOmIxpg37Q+Rrg3RARzxZpySql7FXfUm2pwca5+oKoGdlVAkySaEWN08
uGdPO493PlcT6IpXQYxKNOTWoQItlSyoESW2Ni35DsO+gRHjRNfi1+SQQgEKtmcW
ggYzkozLEel6P7QiuJdmyy5NNflZSVpgkaMkhNnNxxr/zFBZo7TpkZZT2j+7YfhM
Y7wBuUWRl9Yn25UiV5hhnszXsaMBFCfVBBFBh+hdHB2z23cE4F8n4tUXCviKlYW8
apsSw1b9Xg4jYyVzbCfRDI6zZ/XTkuhdEfQcYI7Evn06IHj0MLJEUJqRCqCqVAek
D+0NEOC26uPi5lqY/yHldZs/W9g3Nv/mHGa3bp8iCmqXBaGT3lh0xx0Jz4rLq5+2
DA9tm88vt8ptNrec7I+5Gn69u+93+SLW0CzhiV+CW6ue4MI0O35XWs7ESViFAYP9
uBo8xh7bRDnZfAFf9+K5dXHy5AgKOtpDVBSsoXvdoBWYjjpwCh4lR/bCcHppCx5Y
kOqJj2XYydaOrYIZRQY9ITEAM6aDFBgg3mTYhVIm29z5ZZmxtmg7G+9lXsxbkfQ+
kY1A/lVfhf+BnHJp/VB3zvctLgK3fUPpR7tPfVFCHAr+9f4YkilwhXPlSCbZpkL5
rxmJshQvGi73apr0veuXZdV5TyvMZ+OYiDal7xTVtgKO0wjZgAyFR8F+RIBBbIS7
Jg+idBGKsAFHC4B46Lse5uCu0alKefKIs2ZxAo4bt2aRwdI1bMMYsOPo+k3Fc9fr
sNwBgVe1yDHed8pNAwH36B7GtdVc8MIE4E4DpqGX3HIVnJLOoxAAnFMYelyecDY5
2gyZjYeAM9PropYct7zC78PlU5iodV/HaYqeNLIOwV4ngj65SfG0/NZiYUdBsy1n
hvzoBGiXfswSIGoic2mFvX38cEhEFI5M8n/uYB6LCMxUfVlytkgGHh8xEopVu3Cz
ou63HDcJAYIabd8UCjxVez6BEBF6bbStscvxCkpRG7WhYvkH/Nf1KDooZaChc05k
cVFJqFYqGpY3qeTel7dalqUG2E5OWDBIWOqsSn2Oi3KV5WcWpxTan6VjcwHn1/QR
EQPAA5mYfYKXOf1+3j/o3TO0fkfVVlUMumN30AXP7fQRVBVrunthOrHAWcG2qFDT
hBNhaTVf61dd/M6eaG9eai8WueEb5UePTGR7jk7UXfkumBb2Ubm69fc/hMjE+ZkG
+ri2JleGbc1iXdPMFYFZ46U2j9QUS72abDZs5K+RX27cnjIGVph5oh4pMNDVY56W
ioLcoGJYWwCR1fwBvxTIz01Z0kvEFrhdXRsU9DQgORKKwlEZOKqYRRyOfkC8P44V
KKbgNMng47tu8SxoBw9nMf2UYrJ0ORpZMpg69Q6rBUSyY/2mHSXteHqsWNqIlXWd
7fZhpoLXgICTp95FGoofmDjEQdVTGmU/wR3CxAGl1OpY4I82HXXkvlj+xzYLQ/rJ
pOZc0GnuCZTm3TOzHBbMf9lzNL4WstkGHG/ZPtb5/3tUIkpc8wvetQvkApPwbSRm
vVEFka8EyCIoV5ci4whoi6aLyMmPFZihrM3IHJyziUEovXqY8aClhKFo5k23WTsu
WL0EyELGelKqToNLPJOf4S2KAtAW3Us4AWvb2VLxFNR1qlAEjgEBv/DEPT4yl+Kf
4YP6R7SFUa+Qo7DQ1Cf2c2SKdlDoy8UZcuTuST5g3DojN5WLxeJAeFCLzKoaZo0o
lv48BejX2KeW7oaFHrbvyt13WJ8IaYnd12Gs65mxGSrAnZey1yZbCVefXAY+us5J
uGlVayepyWBrZJuS7ad1JE2y0EzYB/6dY+RbTgt55VkmhB92WPHMtaqSPD8V6tUE
XpoQhXoAQINjCrsUT3dtGKPxUdPmoXJu3KQNXuKOCtXxmy+nLVHWpRf4/QdiZEA6
7GdIYivrKPGD0Vb9f2s3wAF3a5p75e5RnFBI1Iz278EVxG/e/0M6nXyiju+HxwTA
Q1Tnx4YSg9H4HAXavNZx2ZmH1mC3an3PcwD0qndIrHoMzSToZLB7y90iFJd+uP4V
z3RlCb8vzwGKIPfl/uAaqyDGdf1Tkuf7ZEp+s3mslUXaNiN0iUD4OHnH9g+dKNPb
vPvOYgtKbs+7vb0BA/KMjpDNo+OMInZ7tZOTevAe9h4DI6CC+85XJhc9Qdfp8FF5
0t1/ZNUsZISqwKBFDxMQDCMtCSxtQ7OB6+BqffESoNo/xD2KkPmDDwrtK2gw1M87
+ZLAbZ3HBrVYOTVK5IC1m2SZoQvu38RSzGHqa+2Nb8yC6aW9isyWyYoCIHN2839U
qyeCm5OppNmqPi+I8Au+qJ+WzCNPQ0v6ouseC4Kxu4wXbKVClyodcfw3yzLAuj89
uXVygFtIKpZvQtxjaIsLAPtpzaPW8Pxuv5TRiqz0tRQETda1wf8KZ5m6PvPh73IP
KOT7zd8txSTwz+ITqRFKZO/1t5DsTwjMkfuxRU5q6BSFHKWBEs0mfnkmulgLTi/s
VO3M9de6TYHk7qd/IlfnEc11T5aiXOvrNalXXz6SoUJbqhED1YVEuN8Kc4tsJBZZ
Vg8s/fvq7NEDeBfBMaDD2DuSeOp/s39DOZc+vYUEaAHJW1OWUIHWD/TRlF+K9Jrt
eFYIaIdMrAVKv5qUv09hvjFAIZ6FjZxSXaKN3+PEZ8gVZiOw6l5JhxV4E17b5t6c
WjxNgAZ5z9q9vJ0xJk4GQOGYkT3OfKYyWciKC1CgzzzpqsT8+dW7u0kuEusHz5D/
CUlIutZFF2YFFHuM0qs4zZXFSOZg+/MSCrCmoM9eF+Or9mhriwI/y42yTQaGXG8d
RPlLsGe430m0sSf+5QmPCdLxyeQjetufgVGUj9H85jVBheu8Yus7bZmuqUcGuGHr
4vgZYoBHVj+6WUPCADHLsXyoMvczIj4JVtKMGXszFVLIqeD7hUaT3SNBlabmwmah
N22fEPj2PeM8OZ34Im+2gw3ot3a4rs51015dCVs/U3RzHcuoyrkRXWlz9uzex8mU
rIhhgmyfUMzsYoOtxqtya/9BwrkIHdH93xcvSOuoMs1at6FZXI+ZaGwc1HlBW9Ai
XFCp424ML7eNIwK7rz2uFlbShro0DQM3HaoFzCFFGtBd230nbvteMIOHTSWhjRd8
JKQE440NC+viV/fhTJYVvECV/W5He1KOABPtzO57MGHgvH7KrJgtwG5GmTEZLvVA
uT3+C/CRivjg8gE6mFx8rx3W/dv8lBHrENen/Ly8VEHQOSJlDHBxBzdbqiKS1Ma2
JK5EUP8+yp6bOsr2JAmiTMUiMRmp+PLvO+bA6UDdcfnIps63mfoUvC26eD98zSyP
0QzGDzg+YvHsMLeTkGp6CEy0oyPGMTUJJVmOelkUPVmG94qejXKc52L9PgnHgEba
pwyMV/71dd/Yieyqot2BNKStmyu9oFTIb9GVVKv4CZBJ3ROQlKMe2L8EI73LLasE
t6yyh8FdQ/dfT3r+AlEr8Vi+5EYJDpNubNYbnAE4fFazXeip4/HhSEIsTvicZSWq
BZr1pM7Dd9pwGpD37BZ4deYgARFcdR6LSGLWOY/OlAiD1OWBpSe/9zmX4kYxZLfH
Jse6Qt226oexlnhaUsqhSgbELZSNQOQy4ahoUDkk/yvGHgm7EPpEXtcZ8JKImvVI
7BI1SnstiQra/t2RoNjIpnjBSZJEFVUbEYl2c3Mbb8JPbfEPoK1XsxJQK3Rv24vs
lzS/1sxycSkpgcMzArA/yUu3EzY3i/JuTGQlnlSWUWOypELpJx/u2RCBI6mDLAbW
njYsXiGNkTk06nJSkwmuWjt/lgs374cBN7v06m0e3/HQvhxSeCe4f0yl0pAqvVbO
sfeYuypB4P4u0DwOOWw7piyJjC+RZrQuXGBwUqNvsvPoZYNHD65OJFGOOjbe0m7f
cDZZQuwy8hZLyaY50QaegaOB9jvwvGiTqCxNYCawAxKIg2WVtZ5I5mbqQazKm4Q2
/nVQHQBzVUEB2GzfOq4SRCYI49GLUvNcZodGhwinQpvbKRSFjyNR9y44WDxBdcf5
x/BdM/nU5DevxOZXjDvl1ansXGtKtGANdpo1c7PZL8ZrWSwew82ZeK4YWzjOd7Ny
cTDI47HoSInAzcJptKgVxUnlBk+2pm42zqSuo8xMt5MePV6iveqUy461u7qXSKYC
cxG5RgXQ3wllEHR88Vimx5KrIY0OhC1sPAhxPDu/X/ZUwyq8/ZJ93ra+bXyfjspW
azJEQhUMZghhxc/kMXKLKpz1EgpqWrBNQbRDQeuNffH6XTkgjPuJvdVe/K22jPnp
3Aw/hYLbb02hK1COdXq0VSdg9VOb3oZx90tr49QrQba0ZCQmUT+QyHeYJ12jEt0Q
fBDjGKgUIZBSt2IjioRu8mSnUDaXcndpbCdEARVrOAWvX1zVjaDYfbo8zxtwW9qt
O3Gb999g10kHm6CaJecvz2den/ru/ATjLO4C1L1mJELrwvx282nkNWq4ays+Yqa9
6vXXw42Vy/KogX97rbfw7+uelf3BOSd11VhECRKD5utzbPBi0x6nJdV3Uij+ElEU
2ybiqk7GoavdylvtByilDRUxFp2f31ITN+847b2dz+7B0xvQ8UnBhG8oUnfCbO2A
XvEVVUNRyVWTdQCmcXwwSl1z0aDZB7bzm2wniyzDY9wwI8VY/ZOsxfqw/7JcbJgi
USCUTH1ZzuSgIhFcp8UvI4yNaNv9lM20KEuYeGGNknKMMkZOLniTJo9pTxcEMFwV
G3EL04O+zx/Dxw3fTeYVa2QEnjlc6oEa3M4bo9dkeYKkQmOMapkTTNbedRpPEi1h
TUXkNNK3o97wEByPDc7r0mEcXq+eWcYP7PZwyBGNPDoRvwe7w52rk4AyP7jwYsiP
CNSWY7v/fvJmO31vHIXvQJPFBn7Fc9vqJeXbzLIvdIuy+CCcUqVBWiLEKnIyTVs3
lhrs4Q5VitejfkM+iKsXxcCyUYuXjUVe7luyHDjjRvgcEjMGZezwg1tLtAlM/An5
0euL69oXfqU9+cBkKP40xZ716YtyyOv2jqIQg1H+dLRPffkLBAKcCmDxkrUIGlQ5
xpq53b4mfqBmXfh3GWSdMRhtgsjKsBIVeFAcSl4GJtTb/MGUogsESscGy2+RclSk
QhpodtqFi2tP1kd3KtwbITqLdL0nCJSsrPvKdIIW4dAmkIR6fKalZE59g5eSIZaP
4y5W+Qur9FEd7cIa595qIAiBA7f6/8Pv3/12nadW5cyGhxC3Fl2hYsnYGG81k7Na
2rwQnVFvHuw4X1aNPlQSZn/G7T8wadFYTER3XgeShkDNEVIYx41VOOB0/KVPMVof
ul0UVLu4P7wzL+pA7mIgcm4jGgtiib9TlU0MmwnqCW1Wld1/MgKR3uywxnXtRl2Q
jctgvoEeURCqGfMgKGleLyhTq5iHii1enZnYv6l/9h6k1N7OOtIrM7KxxmWbDAiG
Hd2w4v0ieBXSvcR0KHQFCgXjEpzUuMSqv7Bu9dPuE1rX+39q35ee1YB+J//FelJ4
JcbPG2Dv2GRqiyGAobk4IuvkUzPNshMkhPDjV66TaXlblOp8J7PGHn3N9D6NiR8U
XFSx5B7lLSOcAq81ROpQtnomygKkQwV+JeiyfZ+/yFXFcqMQ+Sp5x3/cf/whNJvC
sHUGv/cXpJ4cXc3eFXbDdHuulJFJQQd3a0og9R5jFkm0FP343Md2oMQWAxlQwQf6
RB6P4CnjCNsAH+V4O/Hc48wZjdIHmRmxb31nKzxR8/DBLxTC/0Di0zlxmOF6hpth
nEMMele6Tyo+OrP6uqpbmnX703RAVHv3jXpVfT6i1mrXhMfvcOa49nsm5faILXAq
qNU0+1U4meFB0PFJ+hEiTeY8bEXJKzEFkW8xiyszI6jPfLLGYyWfjIngIWEfkD4u
xnyvc+FfLN3IRR4qzYSprbg4RzBIxl68X6KAbgJVUBXidConlrNizKp19/o10P/W
80HjjPphgJet+08eBzl9bC/rp1/JTwR061ksJ035n58ZZ9dy+Pt3O7GTrCEsvbwr
B8vZzaZw4L8iWhozeYTIR7cWv41YaDb6KGP5GP0m9qFJ3TP6+GFOl4we+y95JtgU
A2HQu/s7Idcw6Iyu+ZiGdCO2i9mI3b6337OGwCmMJ64O/VPCvhVhNR17V5vw1LiW
eY9nITv6bfAsuEo7+NTyf+cgE3DicXas9cVCVRZ2cNMr6zMjce2QTu5qxauN7VtX
ONwKdi3R/u7X75a7Def7NxhaMcdxjh+psdbHMAQvxmGCVqIdo0A/DUo73Rx4zQ3d
kDY+Ec94K97lrpN0EIswAQa8Z3xqmGQUqxLTyHU+XrwgidZpd0bR4BscfAhOE99m
+mDKo4LFGQufnKTLJjdZIc/n3OaVcHe4gymkGO0ZspzhkCOhyoI/ifokqZlmWlr+
WBWK32SrcbVA/GQyaoOif1b3gTm+yvhHHAyqpUdbRynAZCsP+XcexbdhB/elsT0w
dKipnWRxUVQQPq0VKsBoyEuQg3MNgBsVtGjW6DVEjQR5ZD04PoK5NSXkiv2l2h7I
2lzn7uE/3VVAbNQyChcJThOnRxi+lG6Hjf//0sMdAQwsz6IF/8LjOY/U1xeblgRq
jAcNvtB+gTn5Kj4HPIi23mbRgXDPwP6mHQow6C6Jo+Igkpzps/t46vl5Zid/a6ah
jiS1QkippVNk43ilnKyh7bKC7BU/GkV7Vlux8lv4vqmz9LpNhjtLJUwFCEs+Gph6
p9+8pBIYSqYj4Zjyd4hQNt84E1LCdZoYKzhTm95wEl0jcYa5B9MgVqKvCgWrac++
e323PLaq3xMsZBN5yHFxNMTYpSBxUYnscuUVSHjyiL0GavMEhnjWMmksIz8k8cDO
30OsJKG0lixkRd9L0tfvDcUrp7YvpzmuLBIoqaEaheR93z6Ch4hOivzx1qIkj+YL
PyjCSw0oKYhgkqcBT0S+wBCCFvSVqjUWg7sc7DXEP8KFldu97UqDrRyAWb+5SMZW
zT3ckshnxQYfhhJm/NeAyMc5e5NSwbQmWkkx7Kq2YzNliFarbaYcxUkM030Y9Ydi
JIrph+XwV3pxLrYyrSuQOHSogCbmqv5fYG2R3PISH4ICXEO0GRpWVRANOwcjett6
CBjpMbFD8wcqO4msachf3OguSIoMpvIScxqbP0clahLUdgn30pHGsFEWLfN5uGXi
dncihvB3yVLF22YpNzd6hpbo7X40EjaDKSugtajAKf6+NbKrC1TX30EgJPZ52VMn
RS9JLofIv3h/CQqSkidPfqkB/UkgQUMPAndS46tGJPu0U0ETnjOclR8WvEBWZZ/i
Gd8G1GnWNCDXWWpkIlf4V+4tal3O9TPTab9dfXlkksWbpj+AL6EFDgMB4tN1l+YI
jWdtq9lbWlCqV11aL/BVR0j9ud0iHUW90dUKckUW2f7ZTQQx2vyAcCkS+JQgQy3B
OfwUlScWkT5R8rhzY07KmrkO9IK5d77XlSGQEv4X32v1fh8ARrqRyUYvpfJerYQo
LpnPZICDQPLthp+2lsI8XftFpbuVUtrWadHVZ7wonm4/Uz3o/qsVddqC/cpMygV2
g/qWsX/XQeDRxTEhZAamPs5kmPmezamuqKD3GmEKyN9CihxP4HCzYvKhtBEW/4zI
Q3NT90GjpheN79dAklk6LBT5q5bdsFfhagIq1PP37rW+rTKzT1YeRJXkW6W2m0PD
d3vqmcwSou5GqEi4ppGnofKeX59IdtNcLgeDxrUOZlQf/rbDOnNkdWWJXiVsztTb
5kJnbTJuIopWWbNQc9Q2gRCuLhYYYOxR2CCSXbIOr/KBPlGE5WHYuVRJOsv0P0h/
BKcRykJ5q15S8WeYOlUKjxhr9itBk2iUO3lmyqitiBVFDD4d3V/3106DppJNGrsi
LVP13DVFslh7m3Q6j2shAkQ2ANJrS2LiCFg24u7xqHFHwxc71+WoslTJcAAlghnm
bTOkNkhjHwIalgOgcwsY1hM8ku104nW1NOj6hZrQiMGUa4FkTt9KpC4oAyglirgn
9X+pInxxBjRUfrDvdajso/wEhSKg+4C7/9oIohj5j3pnc2oSiHwEAelY1Jwy99/8
pmIJRnmsnYFWPGCKbxLu/y3IlfQof1ryZYC8GFZsBya9wTyVdwdCaue1tH2U4Lvf
yLkcamXo074WJz5ShJWmZFc6H9/SdhN3kU04ytalsh19tbVqn/P241htKK2OZjx+
aN34lIExXVljiXSQWYL75wkvh9UwkrBgbbQNZ7/5SgB+K9LxFzxCixwvlN52nNk1
Cm4RPO6Kj6JsLPO7YKURMSo8d4MLRGO/4suECgFM0SBlQ+ZkIXRI15XQUrqURS8T
22uf9DgAAGIDsxtedrS/YAVMuD7t/jbdsNUhOo/DL6sPUTwLxxTCHHbU2NzvrkaP
/2wBOINY6XFTo9u/E/B8yIuYH0z3/tXDOBeqol1h7ORSR8GZ1jz7/HPYCU1I7Fbh
6JCaVJJ1LdqsKyw5fNH1hM9BJJXKyPreDNUBGGQyymeh7KpaGZBy84pOxDje5SXr
XQLOCluwcHhvdy6stmb+cNe7hHiCQlRoFlZO38+3HlZQM5pJObQ44HlDCFoKn2YE
uauQpZhZUJVwlGEqTIohbgy1/CJGOr/UW24/plSzSGmPunin8qpeRSbAq/UwBLoj
6ZmILHlpMWoCko3lnJkaBbE9P/0Mpk84UqJScyP1QhdapCKaOlzghE2qzS9Vx9VB
RRfQnrUnWdK6UT8RdjSD3As7nV4hkN+1iJw+abp1iIg6UrPF7dYX1pWAUq/Xpnr1
GXHX0qH5aDFqkvSjYmJ61rc6q5UO/Fw+J6rU/FLF2uKHtnQzKEQ/n3rQcDfWBNxw
ScAY2w8QfRQvb7FtB5JMBTcwgzg1T6066qJulY3VjugdhdjZCEf2q/gMbM/+641t
dZTdEuO8AmOknULX+zcsH2bgT8AKX/sb2Y0nywQFYnDvIuNFeCki7nesgZYpf97j
a+AXZ5oYuKl0Ia5LAmmEwopuyE9VZu3ouaTXlcG3oEcvEXNC7qT7QbLml8ajCM8f
2gWpLoaAC0683hFEYNAAIlZ9twU0C8z+VJvGykaCD52HwjEmZesM6JuXfcq7W1ix
sJEDkKqIQ9SRPyVou1liE4qiJmnxF+chNr3uThaww7pNJH7GFoL0q0El1hu+QhuE
RuvnWHSqP0kkV9JIlGBOLr3LOo+oRG88W52XCDI7Bf0cyrleBS/9CCqttPKCkcaD
fUyFc8VjlscLimBGcPCGqXyAk203YqCDBRRSYvr9X4KCNp07TBxJC9Zy4MJ8H69+
gPMgPZsEolbtEWRgS4qPfKvFOn97lVxZKqYnS7ZSyyo9HDZqgmuQOX2TU0vBZ1XX
g3YVgxNdO+o2QT5ojMqibwqi2/Mas6Pf/MGyhwHixnxrp0qcsaTSU7+Z+GHZXeed
vgkQwEwWOz4G6e/eBYGXJAOnv3hYe+o7trwUdhMCJH4bdlnFW7/26RFW6cHsbbgt
dcY4E8ks4kE2lme+s3PQk0ClP9s4YAkyIyGRvPgTx+voB6mwUf58tk63nPnwIvbZ
CFHOqaeofxHOb6itAjWU9WHu2vOUyGswYkJkFfp+ywh822moyBM/ZSULwz7IWpHC
EU0N92JSHy2eOuZeXNdericcV3HtWerGTER8EMjTSzubedIYVoWH/VB2Uf+QJCQW
oe+iS6YsIdqIFyvaIB8VgGVqcj1sKVp33zHhj7SwRH9FsW9m+3S6CQY4ufRnQdPf
k1OrRcV/vP/de9jrhbX7D6IQEhNMn+y/DnycFQIhTNBHX+ZkMne6GJ7CIR5hN77R
hbssTDwRBr2KeHOPoPNmWLoywTf+vF7nzf1COHNagnt8neJ3MoOLPI5KC1LKwYm6
U34Im58lnaVId0ozb10vcfJGG5B/ZoCVpLWmfyPPW4WRQpaiXjaMGtcJKWL89Jqq
mepRRtyd3pQHooDc2aHB8xTe8vkvxIhzJDYTU37r5Nj/u2VGS5xEOsi5x1FqfSmI
Vks1NBZFIPlmMTE+F55k3tqx5chiXEuIBPy7LFdfdqMCPy1wGzQNvyfy0ukfSiSY
gfoQhAWkiD4R9SCTYkwFDkHj3xfYPrkGZg4ABHVa9p867Dl6rSp/TGuwVsy6qQxw
eku6K2VIAfGkk7JBxpFqHY0Lw7CIAOqzUdpDlhjS8rVLIoz0F53IOhXfGN7cIkX+
euSQGdxSRQMfT3X5nh1kR9iXRu80JUvGVjlzkM250pM9/CiV2SC00CLlNwZpRFit
SfqxNK30xSkFXOtBxsQ0Sn1sQiPFKDGxuIUHbgI+OO0ooZUJfzR8RrPidaqPZn1h
Kll/gMjiqyu9mzjGvxd9vj3f88q0xTf3k1QthIuU+4dmvkZyS4zv2Zp7KPQ8+cSP
nplV51DwWJGgDrnkF1nDAI4zJGYK1Y18ZIYm8SZbEbWGiL0ZGxG0OrVUQuOMx4s4
fZd4sguNNcZOO8iZeJ58KBgFwgurYZPWGgleg+efhvEEwgApEuxUAlhwvj1D6K28
llWD2gP3e8zXwKpTbWcmaa33R/6u2AKpHDGI9/HPnNi1sb3Cn6E1xUbRdt+6hZ1h
V1VcPQd82W037uWhgjDOL8MYGBV/xa3VMfm9U3hMI1YMotzr1398vzLQddeXUjI8
NMa4eVPNgZtL650V0kTyqWH1ebXZwXkIG6Iw96XMRKqlsPSxYB7FiKhJiiBDigRa
AoMF0N2gb4vfdRAM7yM7Nco93FlnxMJpoqrlvHJ2zuoWKuE/8g3jTITgfWftPA99
LGejXGAR7NJQ88U2RcnfQCCzaOXMOu/0AZ143b8ihet0wgEMhAJAxwc+mwuL+L7i
qYI0KdSosNmGZUJCFZZxb4+6adlLzCUeNQLvMoUtdMNl7n2hinnDfbqQjdj2nSbK
/u2gWS4sb3tmrI7/DpdaJGq6pTOVbjn42pINIdeWQJWWhYtyKgiF0GF2emTo/L7X
BBOtZfhDpXv2m/xtxHuRVjY17swsqrH8gsVKRic4qLvTOI31TfuhL7xS/vbOQMbw
V5oj+qT+uLzfrnfWxtpvV05TNUZtyHLIg1tPJak+oHQWiVc7Nf2KnFIsKRJfBSEK
aSGla5aI4r26ANevu9YI6g2iADF5SnV10k9Kr6tfEEFVlVss8pO6taCn4e00VQJK
q8OTSeRC0qg2SsV6SM75ibo3nchBhhtYBLOtWnGhmBUx2C2HVC/qi7pfv3qiQr2P
+pPGWiHWjMp/4i8njoYLMvtMyigy+Zc9ZZ9Xz7SlSJezrjCA9VKuK970zdrzrtyU
ltpCZlqpGxs+XJF3ZcJv2IIM1Moh/3mN6m9a8BHIAsiUliH9/XQSrJyNQZAB2PMk
1oSucSzXwrmHOS10Cvs/eCXEIsJixHL+cBTvwfZqULsFSuFYewZ7UmkbFRhKksyK
YFmlllI9g+3Qrd0GefXXOjArFnFlMbsIwF/r30ZWD8MsKCl0BKqGFkaBNHw/4uxc
k6z6FJipF4nWyywa0gRpNSu3fc2Y+muX/VbSwfMtA/vOGSbOglIBCM5i7V5UjZJq
QobBqCrE2xiAISfBSpgj+yAMHFp1kvP1lG9xhO+4QEqFqr1p+PZQX6LMRQQkWZsk
Irge8w/XJanZUoCW5F7ypksqwxC/aJSK9xHGVQ61jNgKpAZghB0kHtDvO2nNyno/
KmH14nPzdUsiy20QAM+3GpOKO+vWSL3pf8HcItj8x9xpLarisK8TJQuVsYOGaJmT
StltjqIexT+SbK5jhpGKLONBjgn7wtzEADGw1wKn0DOGl0RqafYzOiTFDCYjL0Qk
yADuqd4AENaCx6rbWUbXNpiokpkXXGMwSI2xtAPS8KXfmxC1hD7OYE+zcCn8f8CF
WYB9ole6JOoXSS0oDvhYhFp4jaW6YHYd7MyKu/NrMnZBF7/7cjBxuuGnwP2HPAhj
KxMLGgnwpqykBmVyzCFPYI9QCcuuQglPDRSHdwlGAAsSxKR1ykp53zh+bxVWYKzz
HiulWTQBqgnzhaXi1WPNC6fMJNlYX57pG0vw0ZDzWqGEVPnwENPR4eDOcZLiqHCY
/j9uy76ajh1CMr09VwIZXkQrj1K7Kpr8gU9pgJJzFKtU+gF+zN+e0Ef0toDl1N+y
YC5vKNU00ApSkPFfUDTMR0JmF4k/d3HxxHjSdnnnVD4tHYsSs96qNODUFzRESZhi
cadfbTjAObuyUYQ5nltF3HA9WXLfUlO7ogfpzf2Cur409TnTwnVrmJC9Eq+IwFIT
S54iKsLmipJU5e1Zn7WtiHys3s00eB28a4C3DJvgtF/BDxOC4sjKVQPDvGbLt0A+
9DteXbWJaR8AYaiZvoRrEPIjZ7sY/nozipXtRPlvRKCX7o+hE2CelpVLhoMxWRt7
1dOhFzvYk4p9+qiQeXv4oDqVemTPW49H49vB9LLIub8y2Ql7ec376tKe2tKr5CYn
yYV58XTMPvXdikYFffYW3xFTH2kuX33BniVo6U5Dd7DwMohMNIAcBOZq7+/THmnP
Hd9tMxyNE8Gk+kYzNNySSDhseYBhQe6fZdyEuDgYnMQ2GfW0xAmI4vvepdVkn3TM
+Q4N2dmjVtw+4aWOC97cn/d/qz0s5cKActcN5R0U7E5xS1Y+YpEUIY/5/uTUUaXB
C5eAIOK/oDB2ke6u6jl84DmXPG4GQQMHN1xelVr6mSJ0KhMiHi5yMArc59aApnoG
MubXHQomBg3bcLqYi2IZq5ZoodVqhIRm80ZZitM6+HdYSRYOQrhld9KRTEiROEzA
OaPPkKEs9I5ZkkKsQ8oAFQ1kd/hQgl6gNYzMFUHJOX7c7t6OhwiJfyKtWd/hEs4k
AUvO400chRdzNa9q1xhV+Nh92qi7ulcQAZvrq5Ka11z9YwjU2mwFNXbigRLCBHUp
yeqHrXFw5TCJ9K1gX7ZcZfunKu4BYUtW4FPHH5PbycMdh5Grb+bAtafxhh1W+rQs
teCkkyLrGiXwNlVPqj+o4tavFecBjXi6YnTsbv3x9Lntm/hiztj4Wa2ovQS3vjKK
1M//QXXJTRC5mLmUER9oqDF7DyvK5s3cTZpX5BggcZwyho8UORwMR4ivHpkQuKzS
9yShkGr3zvUiaWLxNEjssayKKIaAbEB2l2VV+YsBTtefDSDkTwsGuM+jlpgKejAH
/AqvkR9UxWOw4sJMgrNnzFTp/7nrUsKXqPp0/ACAYAQP7w9Vw72Bd4FW2VEAi4QJ
Zta6QN/o70nJ6T2Qm89YlUgGVQnepI97JF0SKh19dbpvfuWFJYCdE96uREK5GU0X
z5JBy9f7zMDo3vK+gzpZ1NBits7s4faTINLn8qrfwZJKvfFx8Dn8lDxlA5oi4s95
U9QqYty7ly3J+DKdKTwVAM9CmKnZpSzU6RIakNCrFe6IsHYNVxatva3g9F6ld5+B
N1bInxyOVDSvDelhji5bo7DpY40BR2mjy4G2UsQj69RyU/ZDsn6ZzqojJY/Ay9i+
c9RQQpz4pzj3DmRnMR9LxumOZrQCZ0B7ar/qnVSIeamMYfTOFtWhW3zzCIeH/nDv
4ZnhG51twEWoYf3Bebf8tnEmUiIDBsBiS6MGz7TsREcPLAdxG+/B4z1Kyf9iOC8f
OLUX4s+zfudVCamaBlFJzJ3Nb8SCxk4/e+dexD45mWij5aACX7xxByM2VHN+0UPC
S51F4UtKiKQ8njIJcwuSxWvIP/X4FAI/vn6npMZujcC0yDn4uARVYBRgHB4UlR+X
IzjLpDKt7JdBSOQ9d1VrNsz4fmsFuhYJgrsf2NVdre4QlDHQxufwZMnj3zcqJrBt
mKjSXL/dNwbgqru/eRPDwF7vcRXmJcp1vbds++GncK+SjWtp6Up7lACY8SJd8fq5
/YaQ1et8goAlA8EDC2W687johnRU+3q4BbPqdb3SSF+M11Md3BkBYXrwYb2vtc/C
bAudVPNFIyEqAJeBfNU0rXigpMk554yOMLprc25JPl7uDkTweY/npvDkyNF9Zthq
H3sCQ2tRr63bBqK9XWAAJ8sYfw9a9yzq5UEeYsOfTK/Qz4DaTkmBtfAgW5rfFrzo
JaeKLVow4bB+LeLwxokni5esiL4rqdwZpp86p7oI3yniQTvbVF9XW20WNbYLzPhf
hBpx+V0AOU1lOjz41rqYmmwmzpWT5FtiWIbw7FpWz0ClAeQWt0icw2qSs3vh0W+B
mL2xuYCprV1XUy/uyqAGRLHiBV9GUS6cSZeTJGlDdaelaEGe/mVCcJwUxidzPi3r
kOtUGwMzduhKiPm50mEvlYhA/hyUDVEDkH/BELRCVUy6JVF2WfcVu+eMAtofx2nF
AGjisYz+zkw1CR+XEtnIBJhon5qtnRAMC3YIHtrXkEqk36+iPa7DuTKRNgwUcEbs
G1Nll1/fvhdPGdL05BTEhGYzTPQECq/m+pnqbMGomLcmN/VhFYJFbzv8gwXzzX7I
BDVzF4HoJiqJDu3AoyHzTzbvFCLaBVxvYE5bCJNwEz5qBjZ/HEzXZft7EZdwsnPy
4yMyBxOuarbCuUeS2WXzMGi++u/X1PwvCxdtUUyUBWNPc/g7O02p/Tc7gGetKcFg
A5ufsGjUKfnCSWb4TwlH5a5OPnPc1JCbwoC2LrVehdE7LAviSJJYiNnNJUgEptwE
2DKUSGgMBXKQ3UwPK7WJjGohud39iEC9XSX2go2jmEoxCuBnU2rNJ1F416vKmNj4
RJDKvUhZq49UT3XXUNkJ0S85wicEAzddCEykCdkkKQqBOzFfXS3mqlMC6DyFhzFh
Cj2e9qJ6WQpvUTgqkIhXTA9rxIC2yBmHCYILqVifVQxP+v58pZ6U7UvMn4O02j+f
nOrjadH6/q2kC0kWlO5gquLm9+2jumFuG6xxwlx/Ie1gVrSAfOf9D+Gj+MfDDMDy
i2piIuPuXt4Oq+Xdt7JGr4XSyTI/ybKy3ePNBoQBgaZUZILCUb366lGMtMOB1kjS
3nzwa6WtKrVvrMu8HqHYN+cDdpcE5+KnmBlX573h3ACMAoHwPnvav1CdfcYGS62N
6MCD+0rnFcy12mY0++LLcwEpFvNsGmlQAGVpZYRU/C41WR0SBkdPqAR1JgP2ZEy/
scHQEjShD0IOguHrD/1UQxn4WErnktzH2pN25qcnAEBwmdouy6tfFQgTQTjHFzDh
uvmPm1gMSyBlFx42rAozNENcLJ77alhTLCo6aMITt10o3edWZszRN9O2SlA3MoJY
UPo/wyeOQoxwEzL/F/DtITr5I+dMEjTZrwQ+YMp6/IhfqzK/B1xL9g1J8LswtEZb
RqCE17v+MOpmFXr2DnkOnmZFZtV1839/SgQv/15OPv69/8mtrMzeT8aIu8Lcl5Gi
RTPFPRgUAX8GgMjaHbM0MIKW5QrpLjF65IYZe5D54Hy1a4svVzd3sYHppqCp23qo
J9kWGG6nOSQO7nQmuv+31puV2l9P9UVFQ/dz9DmfMvmjhf1iIvNPsx7ov0oLOuEs
dOGA65uim6KPnzb8mXeoRx31DLLJJV3eBGs6a5McVs3NYOq2ky7WoQQbI1TL29Vr
BwQ0LIWaaZ6mEoAnUzCq/XR8mmrBkbeUQpfIFhtdFOQh09gCAVvA0l59y+rDiNoM
XE9v3PG0euQCABk/tMfuTHYjPuacd2WtLaynnmSZ4BuohGc8hl1WYbY9I+krQPVJ
Ua5XYEeohBpFzSezwMgcaszlcoSr9DpMI8VsW59ng0lGLiQLgN+yyeOghaMHPIsq
+64GHMjwGUBGXJdmAXMrp/4CVxJu4BlJwwJHgvRXWhee0UHY1m7HlGr1khzZnzEC
WWISYN/hmTMT8BH3QhDBfdI/ZRcDnF6UFa/0sCJE0J2NA6Y1ZRPxMZ8ezgdTHBuq
/y5GQjAuy8y2fzQAuNmGA4YuiMvagQQ0YuUluGdkNnjag81be5JASCSkQYb/ikZA
Tpjw/L7v1g2/2pxCuyhjVqOXicvO8e1TwJ1h7ztBOQndb7TZ7Ea69xoxFvcEZhNc
YIWc3+sr6+PuN/uI4hIvAB05MM19vJY9f9ZSiAhajnmQoFrFQroJggL7N74oOKxI
smAOIQuFsb+1xY9PKXC+NKAwxXKAvCrfQWz0x++XMPkonEUfGqtncDQ1B6+oPTU9
CHhySKm+QPzNZ1DxOREs3DMYwzHfurjbQHAF8CFAcfXPK+nd3qnq5lg4fzzS23jF
UkhuKFbgVRMrowHz6utiKtRRafgSJcrBQZj4r177PfmTx1h2RMVwvalUAVPR6V1N
pkvF02C7GHIYDjAkCS56FGAMyWCLZhIY84bCCXIKvLV1KIaXNi2YDz+yrb4SfHC2
+hhBlifDaFYHO2vmCjzob7vHGlmQIhywemHI0/BZOY9wX7xOWQF4Q6KBtNGsp2SM
Sq8l4NcHRSKq7E9kCmEr5Hatyi4TWk7bgvj6UiI8myw4J17Yd31HtALLZAnIabCQ
/5GjrmTpnovN41Pd2/snuOabAEB+SqXVfX3JgEbdLs849tVKxYjbDIKebW1ATGWB
s+jjgGI5D33c9cqmYuuhZrd95NGsIb5ATL1C0hj0kRn8km4qwpW/puNPLmfBDezh
S+2BfW0MV/Z5QQPo/AHAB0P9OJbfcBlMRgWhAhGAKBtnIhUwSczRleCcnuQNTwCX
vaAfzCGhZHwqH3MQMv7tlII5nGU4tQMvryAvj/SYp78iKbNrROeCkn7h8zfuTeNT
omUSzFVK5eRtq1Ke7xpg1n3gb9uKvvL1yVWE6RYo1QyPgyxhMlo+F+MLoMGkd0vs
GNIvhp1oM5X28AHzlcj0dzKZ7IK2O4k9nOL953k+m+GBm1dLyXU3owhOSHakrj2/
LuIrcEA1SNrydxS7wpixWVnf8nLRPEEi8byonh4IT0aQGjWHmoYaQWX2d9bAMsrV
5d3RF26PSkGDMSusDCr4mw8tJxkDCJBI3s4Kwu962V/DXcMus7GxXTkd+VbtGp8G
qoLq7tvhiuoi5rldvxyZ3chWW2Hm2TYmN1J83Y/VOFghaqD6lU6Pd70ZMOy1mbOL
u83xgjBdHOKG2GQcBix2FRoATU2H9uNFHzVPMzTBjZPn8/N4vVYkjPn7WQZ7PlNC
bbf6sOuYDQ4elgghYlZGsizuF9MHS93rXwVW432kpNxsZ4h44ecE5dEAXpGiSjUc
5zeBFFVjUy9Luer678NxprLfuWk5y9u+JppMavTjSxX+pfOvqYrz0PcQCfxo+rje
T/50HmZWKfcikAbTgnPLV67fLUtxsGU4AYqR37/hIIUBVYHIpbG9NdhKOGZ2sqm/
/Gz9O03sWKh7UGGuZzwjmyJfetHpl235/7Sm7c+xyA5yOtEOMjn96bv4SW5smoYV
yU46leJdBZpLIoVXVUQILN7eQO6z2t6yPeiLQA4Odhd2X1AlTDQojMeZ+Uzm7/9R
pK+cv8FOlFCrlxnJ9dwo+f++CkOGOMkaueV9nx+X2cn7FSpDgOwe4nA+YvzRadSH
Fj5s9U60EJJwBqwbc3Z723MzN+fvbLEo/J/lWN1p2r+hapnH0Ai4gey3ROttm082
8iOc7KgCGj5P5Z7J5BdO9rNCyctxDqrZ/zeoBuBfO1pj52KQkl5jMEE7iUBWyxjX
U++uU0+l48O04MQIQk1e7xGwjvGf3DETKLjZ/q/k+yye0Ryz/t+6KR14RfHvkoXA
KcCZzZfszIfMYNBSEcl5ZPKCR4Xi9Pzh20PzdQYmrPloU0vJ+3PVcBuK5Vihmzak
75aWqoLSjDfhfrCoc26JY3mzycYlA1Ck2waSZWQl3Hapbg6hV/wd6ilYcEeCfYDl
YAUwgLjPOoeWfZrvswjyKFwRus09iqkrmHdiK/wAQ9NJZicnw4FRXeOHXmlmlzCA
qO+rfeltPYF1M0U7eBoJktPzkt/yTy8YJ85ZlkHxPLgSinCZmT5PsjaZcsprRn6G
sv5kNwBvSwVK0epHL8XhkXYe+18tAnw1eTA4kfcmaG4uITmH+V2nbk9CW4kzRmwC
HhoG038u6Ov/Mi5bTT8ueDcZvFLSgPnfw04JXrQES4gMH3UJjN4gyXHuSucKwjj4
MLJnB6cGnsZ/ij5MrxJsD21qsBQ+3AV50kqskKDa5Sczfw20ShcS6f2Tet8aQZsh
6o1dAaWpo+gz+dqH/Fw2KMh+ZG6UHguRdF1PIQ7JD7oPIaZVVpX/KCJw5KA5FsN5
QNcVQT7juB1sDQQSLf2PN0zWf+E7QnEkH75SIOfWLHk/wsdOw7WEpwIi8wlokkAf
4SrS1RdylOThl/MuUH5blnVKMApd+ws0/Hjm/CxVqWTWG3zMJAM6srUjlhXdrsn4
/MgrrIidn3oICG1PTNiZrg9QGVQaSvYtUoG8teHj0i8b7ag/If+x4GrwIafM1Wtf
lvu9ArYpchqk8ah/5NeXJ7s/VIxyYpsVXBNSSAxaiiDdVvl8fCoRpPolyx4hhQLK
n3FQ1jhljlUbKIfT8y6bkJNb8jCqQmkFakhD5ey8Oc9zEVVY3hU7eoEEDrESFxRE
1KZ673L6F6/sEOPTTDJj/RlDSFDBu85Dh7wZukaL6beNfe7djFsIW1uvKcPUynSG
Uhp311YfjPl0l5E8w4/IAcQ+g1e7erioulV0Daa7AhfIPmNxY0AEBEex7VEILiIB
rI+eFUgp+1+nMpYzxTmZqxyan5To04FIYolL+nib56o0hp2/PJy//MhNylzWe3aB
D/4actjEZ7Cg2k1OvcHH+hcMcfFvJXZL5zTiQTKJhaDeh0qzPfXCRB+3YNXFb+L1
8eusdU2m1VDAF/W/GqI+nm5UevAipRR1ysgPBqtpAHwXsk7MTwLTHdQdjTYx1oG/
zJ4tDdXvWZITM/15ATUg17EsMBzkq9eR9u47S0p3zQ7/nkq931q9n9gXOaAW+ngv
+tHFZgynOeV4R5EoxGHZyMLB2aNJ76cZB0fcVhXvnUQfy9+qD5dnFuq+9IZWu4+P
FwzcxIxgQgTuKTWorjSReYMJt9bDa2UHrYSg+oR8Ht4NLozh4pK4+OBpf3SltEBg
39lyo5LylFg1QIO52RIdUFPihxWwrcWnhwNAteY1bTRUjYWoacZn2k5mGPkW7K0q
xHFy+IeIyjRnuy3jYAb+ZM6yR5Wv/ceMq1dAmBfwBXUlm83uCJ1/8r1VfmXw3oyE
ehNnXVLH1SLcBN3iE3ByK3RV0AID9LqIr8/fJ4AAAergDic3vjKUdN1AhzUJ6jku
e81Jc/HSXm0OVeQ6XTYPdGNdOPnThJfFaRDcwMhY+VGaNYMkHPMKnAbiUkQSE3Jh
jMQzrLiH9UJpGPeVGlUMIfdqYbR5GOaYhbzNkGTEUQPGX83nDdL1Osoi7/0n//Vv
BFhb5iDAHR9T2CFnU82w8Ydyh9ezg7CSEiFslYajazcHgDHIjj3qPM+d+XAj0OQt
6x6t4Giz47VdkCx5wwoF11EGR3QN7lRFPKkaJMLrNr7I3FKxWZ9pValZAVkLV4XK
cRBfYHtXORxlUoGvaYi1/wnJtPHUkoBSWwoixdCwgyuViftdgLv2shvttJjMJTfX
KYI/8FbwdJI76OsN248BrJ5OR5EKko3ckLi0HE82QRQzc1nnThC0ejtPjBR6BPBI
poaLZa0XgPemjPSryd0F1ppsKfXy+StwB25/cCHJOe/zxqKA9xIYTFLGg1jmdQPK
EYiY+kAivbVnQ1QHcOEYreGQspU90Ae0tbxynMu2GklgS3gVaYrx5GTF1+UNW04A
9iWb5boAJ0Iqs2lCTxw/xLexpLCVHV3EWFaq2b3DRFpkwWJpz+GlNCKwhf2uViMA
hlwVfetOLpSzb5RLl5RdsSL8XNHd0z+kHw13iN3n4R9PyE0ohiU/GErI3oj2kqGU
Z4mvVfgmdx+XzCsEdqlExvKm5Nh/NmUiGyIYZ3t5d8RaK7lOGwsG+kIKXTeIChIA
16z+oESTAlXYDNb+dEVPJ55uCBL8TWDEatoFBFQ9TClXUmj2jmKA0nexgH/EXo3g
c5DNxAmXsdp5g1qWh0hXxz147SRidTdnywhcKDneO0w5W4/HjoYtYB6tlsp/wuvV
fgBty2uw6z0HmG8TIsdPlOV8mV3b0AilQDMAyeAx31P2WO5C7iERw08V/G9hWoZ6
be4TmquSSSC08IMrsRskBSocMQhSRsEl2fcw4OYMACx653VZmhNuL+3w6Y7FNvCb
Bps099NJcFsgG9Xu7s8cKw7xVx189NMxoRIF0PVJhlTA+t8RLJkwQVRR9pQjjtaU
qKZiH2t4S5TQw4MJWv+oZ10xiKFL8KJgrmZDkTGDJiXYy6Lne7a0obJh7XNjQRO4
Ru+glwrKcw3vTikNUluW8uWOQ6iAbPWAG56FxFqXT0y1Q8MeTjxJC8NrDO3L9rHJ
VuZsOnJAdxfCXjgntY5yKkME6SOI+10LjhP6IVVfqqxwz08Wbazn+tA+JcM0jXhd
tgP/CaEk56BB54PSvNz0Lwse5Jl53hPNT6uWFzt1/HNzuViAiFepzYFibdMDNSlH
Ivv69p7/rZYYTMLfyaYOKkILo2gor9Mb0WgTIZdFgDIBnPNUo/uIhc+s+HOOVfEq
c8VZufLaxoOwY+pMxAQWFXWXxMIyx4imnBxzToY+NXlOwCc4Jj44y8rFhz/sh6UM
0+hSOzCLTDiPpLQtWi5+nyJ231zGK6qPfpVdmwfz6Vz4PTpQ2GtjYv2QXw71yC9y
2PENVN3I3VZ+G5YYAmt3+6/KfbddiQtsGL9WsYR/Aze4TcJ9JHfZCebL9dm9Yl7y
st2QsKOwy8uGSYj819pkUAZdmIq7kRvnYDpAmmle8EYkYecEJAvlCrVphvXVm6mW
bkF2p4WrTxE0SBgwdZkhzdu/NcBZvtvtPPTB4hVF5h/U39NflEEiMCLY5MQl0m/b
2uiUDL4x0PMHMB63R0IW/nektT3ElQX0xe9E9R5CW552zVy8eyKj8h2aqP6S/O4z
LuGi1o3hXdShSbC/o0CnhteghiEQ8Gv1pP0ZW2NeZUz3xU9RKgpp+DddmP9tKqVM
SCTbzLY1ZbxFdPBE3k7EDvPBFAAqCGI/oES/4aJfD2PhoJTjyTGRIO+shAocC1ih
HvflozS45q8/TAdYL8GKKA9D2sEs4kCo+YkWy5m0CXZ+ThdSVhbBpk0adLsbqLn2
VKm61Ta+skEMNgTQ/aDFkiJ7is9Ns6cIBJJys71Du7DDWGIupXxCpk0BWnBPi8Ut
FL2PitQcpxc3hzAWvch8PdmkgwKeyDeqWrOLauGOqdAF4dQAvlu2cl2r98UDqCey
IaEHWbVVEh87Icutt7T4KeQvfbUCpj9aayX3rzZOLgrHTweoK3AN7qc6R4fDOiqA
79rXRIJHiRU2jvYVSg68E1p6iBuD7kO32lR3rezlfYmtrjRJVr4WHsZv2BeL4DC1
k5uE+Lvua2SulIt2xSqqbFVsbddCoS8KJl9M1Vm7vmK6XcKRNFWAkSBBwLpTXrtL
aDmrcDQEFQaadIQWThMCXsvUlNxqa2zB7mmmjGW2JWMW0jpnyHEy4PRX5OvbdWQt
39IHZZuRIgPU+apzwXUMRWxa9EXBwx9ZJ1zHFPyQ9IhkXQhlEf0fg2PW2/QeEGfD
ydMM+kRW6FmaISIZ1Y4VBckwthaRLPnI1XuqKCbbAuvy+LPCFQ3+nkiksH0owjTw
eWylcGakgyhQ6BcGvq0p6ZQ693AZoBRuuc1seLStDD6cN1Tdf+Wg+J/GS0SBpVrC
CPyBQ+m7/i9TvA1jeWuFlPH/ufXhgQFzOPQLueHSIpR1uAzL+5wekTC1uqDo7pdQ
pV2t517bAIrIllrDxbDxcb3ZK6OD4Ilg0gWk23Kk7qBMVLVgDousie+YuwTcQYoY
w1c08O40MMTLblCg1mYqwrkeHoxZVVbM8NEAqyQuOdehRUyKpjttlLTIBSAks7R0
PTq8mbCmlXHnodSaYpr9dcxu7dtQgB46yuoeVex9xlpwgdKSSrifKGptNqIdaCq3
1N/yzsTrYudaNhujg/z3LrXC7C5E/CZ0R/FGbmjj4gASmCaN7mh2VQv1yIYGOI1d
kjgpzrQHx3rJFOaYM6RFdRCXXueX0+5CwtVWxxlyRI7LCB6+JKp2wPiNJHl1Bw3L
TkAhKkSYQwxFf/mGkflyPNTAz5uJgzw3i9kBHkHfN/N2DUJJh8CVu3354ziU1XNB
fQlenbSL/o+VIiADQF3XUzEuPUbhzDWLPPG0p6gavt++qG4As3mNofoT5EhaiyVG
KzIc2EdlVCXGYn/XqCWfpWtHyDAV3ixAvGHqNKJTyVXyIn63tB0pwJ61v5WsBKvo
Xqcss3UUqNy+ezdFlJlmiyKwQegtHAR70rfBHOrCZb1Mo1hknofSncpFTa10A4aX
BtyWpzT5G5TQXa2c+bygNcTL6G+vLCx+P/zUcI5cMVI+B24xrP5yW14ydEp4/nwh
2QkP922nCXBJK3aea8h/9RgPpD/5Eu+W9WNgas38DImIEr8ebO5zav6m4q2E2J9W
IKJFOtOXthhFs2Ewpg71AqgHmge/+OeMSUvKCDko/O5PjxFmABgi5dzqCmUe2gJM
8ApjDyks/MDG2NiODwzFjg39Yxijz2dh5ZigvwJSO0WR6p9+xb9hpMKnGv+5K1Ef
w6d6y3JJP4Drf0GClbjG08eoEMy87kNn9DXLiSOl2NSzx4p+4L2V0iteIHG1m8pg
ojLCnreahh9RrzZuzfCi0QeBlrRTfsUaxPD2qcAdApeU+VtUZTBJsPs5b1Ypuihs
UUPsQHbKtehkfvhFiRxY6ffhnLVI5om12Nhz8DxPibRAoShiRhvUE0gEsHVz+ihH
Q5ECZFrJJL+aKmDB8HRMOtXPdc25jro0HZ4FMO8FJOwz5i8qvhV2AdxxbtzXBkIl
tRTNcGtka5y071YYGsuLmH4RwRghuWKVcnCabg7LgF3HbQntv0fNDk798JewAyJr
fBIyvvesuPO7hwSqArpwg1/RipLDHZlqhb1XylsmkbTv0QK/W2pvnG7/8rIhic9R
XgGFMRaPMy2KP5eUBNlHyw3uuq60Ku4Pq3T1xKT/qIhfuSJshLqc0I0Ko5rRcjIK
T7EqB+tDDQvk9bKSdVE4ZamujBwhEk6rXAWFkBwvZW7wmuJZcC2EeP/53ZMbPBsX
7w8D6d3HVyiwz7x2420oETBrAmJMIxLTWJ64hYVWNYphYI4QepRNN3JczIh/Ee2r
SfUF4/+Y/DKYpFerCnXTgkUa4QiaJxgMydaFS4YCDwiWxYuaLdRkumSUJCgx/Plq
6vCtUOzXcJqQ3tt4EE+LzyP7I81X8L2mDK3/cNUVvWCUlDiEOvYEVFhMj+bqCZpD
PGQjhvcL9dFjqeOLI3AokKls4yIJLO1vgSerhurdvpb43qsJl2lhfMKVbLDGmFKg
JgEafhZlyG99QheOIFgXEoSntHNypK5d5uGaRHeNRL/avlq/AfIuBr5MMYK9ZVWK
K8D03tklI5hlf29YMTGQ9XM3lgzYkOKlR7MdtzTz564rUIICHL4OvYxfzzKesrWM
8Qax8uSv8LXwvHzgxdriKrs8Nk5Ar2YbRPJWNP801evwwEe7Mw2kZuQHFICyqO2v
7DR+SsAtQsTI98QOjV52Q4Fu1dIqA3EAllyaq9jCa7usukjU1xSofma84hlAKQ4v
arEdc+DCo5Lr9F9JWCRvXqySIoQ5omlBICObpQxbmDURTKKE+IUU/j5xyRQDGTST
poIQbepyH4D/G8aNmVEJPARuYLzog8OJ8cMAF3pQlKqNC1bPbO/KvJTOBwVP77iQ
3wxJjhfCZ3zAT00QTa9ZfBqIKnDtGvP25bbYH8eDg+uCMlukpjVl/wg0TfpD+iYf
o9dSRPfMdVMAkA7mQd7fsH/uzNNtAkai3jdzpm/gemRTKdrWzw9La6d4iAsXsBqB
9C2p6SMpTkDXMIOuBHP+nHjNVgkLClAZ5yQAKpi2isoYzL90RUVKj4OYkocdNwko
He37LOAqu6qcfLRro+qEKDj7iII/BI+AtUsQk8YdGcuEjt/5WZ7dUnJayLFiPblX
jiRYX++otcvqVFnCmZeOxRL7YNLmPfzWGX9DAJkSkhDDnBQgsYdyrZxOwNF4mzc6
7CuYGtI5G9xIjuTrNB/9v3mxX9wFEkpPMO9W/qX0FgtAbDcQCG5QdF8zZs7UigZH
+86sVelU1DrKxVEssFxVDrD5YA0Nv7RA2hVM9r+05x1qrFb0CKxrq28cSkLBcFbP
R4qvhA+BS1SbaPOcD/V6Z3so768QqVE1VTWuNFT5k2XfZdPCU5d6DL32JT3ltxA/
3hqSF7Z7Mbp3zNTwyOD70WA6TNVAG5W6tXSHMeHegN6jqKkIgcbQn+EYw3ZPJQ1k
+MnSgs7vJ/kR3O8gEl8FJCm/X1GzTc7ldXffIBO1Iin2mmRqBP+4O2WTMMiDWsf4
vdPXJWit8nu9VpSR7zB7Soj+ttu7v5zD9buxGUCqcMuvyLJItQZqNNnpjdFFIuma
r88pj9EhPsxgENZhoMMd2EyIbytdahqBK9DMeNlZdtZgc4zwFqBMbPNbZDY7lKTQ
Fb11VnY7QkZBckX5Hk+pEH4bEh2d/XCchXB0nEqBYdHtD7Wv+k2JKAMhEfdxkK89
8504tt163ooSKSpVsJ+5jckAocEB8DO1sac/H+mlS8lj+tqQCyaMvQAyETUOGYtf
KzuVsaJyEVnCz/eSdVX4asTlkze9Sfm4LFOyH0+hT9TcGobSDqJUs+5Hh7K0mL8k
fhDlNiz55aLZnXyT+ZunrC8nJYaXRBHeoF84EuP6Yu0B9nZ2qXgiP3FORd9FRAWw
OvgttF40uWweRF90Rl8YSYwj9uhaR9L+0Zgr16RE6+JuBxFox6JmA+RrTDBkDYfo
sJumptuLX3Fi/CYyC3HUO95qyAhb4D36PYFLwJjLmmneMMMwyK1mOiOKl8exC6DT
xYAU/8DpnWAXh18OOHeYu317zKgcyja3hnPrANl4LXY99MtmB2uNLGdIxxAoiR4i
/QB1Qu7KJAiAbFJ57W4l3ZqWqvksdir7e5mBg7S1Otx8d8oX8siyxLNFKHgjKq6F
mkGKb7ceR50iTmddLfXSjATRX8NIiKHQpLofbVfRFWdoiDSYBEjsSa+PcfBplbFN
UbIuY7E1Df5OcoKUU992PBVnqF/ndabeoagizEz1ReNy30h4idYscZ26st6CGvaK
UgY8y1hNnAzcmgQrkznZSlGaUPaHr2l9sZqccDn0mJJO4Wy/3A0iCkbSELX9n38U
JpIAM5BV1+R319KAI0Ld0utnupwwfMoltmsNxjEGuVebHU3NXSZ3a4ynxSsr1BaP
32VkT09cfuETOv/TQY5EyqL5oz547rxbSxnvQ3Yn8GM3NpHyOqldyFrAx0bPtD0u
AbpnZF7R3gQJYRN2o2zL6MPsPm21ZPuoy4QaTi6OP7zdUxTxpmWspzB0/XCUxAKm
05FcH+a3iehVL6YpHGuMcz3z8RJxfxIxu2FJiOZYoPKK5e+jBEg+mM/8XO2gSUjI
n6HdnNMQviy9fdkABrgrfphgeiZ9t+NfukzUgLL91aKvwFq20BEOs13oBK5T05ID
exnDUpMcuQjrtMNzqKTGKMOC24ziskmdQzsL3J1Tm6+wRE1ZgXySegbdvE21Y2IC
ZfxQq6huxrVN2YHti8i1VS3EVfbowKsWZnzT49FOsIHN7KKK2zOEe8FUb813UcvW
WGeUmBqkXva0PBWUMnWiz8UJ9EkjX1Yy+STtTCp/suSh/nkqBga3Aki2Mgc7USHm
Z+tkQqiCuyjiwFOzb/MnN/Z8Iq9pVZZXTI8gfw7U+P39ox0+eMASRfgS4z1MGk2Q
OmwGyKaDJuEAKq83CUe0fSHVAWbMY1bdsV7IIXzXy8LTlMFhgEOsWPAeVG7Ac/gn
AItz6JkU3DBCiTK/Ny7LVldyXWnMSSGDX3miZUC9tkJzeRMC/qNV6Su7fOifNYbB
T3rZMZPJ23hntHeKHHnEJCx6pCq8uQiI+leyYRjECCfUIm84xoXltdogZJYGEIWx
qGJBxgWYFGfEio2oLfP13CAEdwncBCChVE+/zGbjSLrvWs+65oLL2o+I2f+OxQeP
/ckEjjjEnXLa6125ywh9KSn4MPGud8hNejtHVAuuYe6vsPamMs1Ipue0516s7psZ
zlOuaCCkWRg/5u/q+zuBbSN7esDinmLlmKZ1nfvxYYKCdDioEA0woWuFdZjc2OCY
s2ZOr5oNEMIuX/cbOHkpImg4aAvzMycHavsJTrn/1M4KohzWQrjRB9HmPQFMw/pQ
XrVhZp6sVRLzLg//tC1XD2LlcRmmwvPHWxcBdpWXOFqlzmpBdzax+CmkxPx5iAur
ND0No75B6++RqaAjVI7ytvgISKN9olkFWMSZvGKB19gCCM0Yw2o5f4cD1JN+T0kp
kYGr/YfLVAGtsp64dx6M6sn7RPT3ASQ+7sPHakGJo9vf+HoXJLnZC/BOfdSYUy/z
afuLY1s+WChJQ1S//nzasF1b+Iq0BIwX0qLELEIfA3qEVjsCumuaRBNQj0zGalzU
KwuTDMPtJgsgyV/Z4SKYTdsgsQgMnnHSjSdWWdH6BI57cWUbqyRKu32y8I4IZicX
FAWxImNGj63jlEgtnJH9uCylAfRqPYWer9E8vhnXnfN3JSnzfFWd9PQpKYIMP1vs
QcTPe7UzY/js7vRFKE4YTrGxYUQjZXdC0Y3FrkY3R5/AqO/tiZQejgvR6854ADor
Hfu7YlaQt36zKy9YQUvgiB+95N5eLijolsbYTtpsi7+cH0pVeZVSt9EZex9IKkpq
xVdekNhsnlpmdFbbsMvnEZ8kNHen4wLMuChMDpWv7iImoh1If4BveVBFcdhFfA1m
6q8w07K7nah80+HmQXBn8kYwseZCq8XEtZ/CvW+rq2AtFRm9njYjwPGK4+qpGWPd
tvg3PXwOg4fsR+spG21K3ogiXthzZg/nio5nSwegymJj/PWr6c2jOeKAtoT2oyZ5
9/GeRqHjTwfvtOaI7w7LZNG7duYcFUBs39oxYzvbA5C+uqJ0AKMaKLJ71EyiCoxo
o2U+1HSDV9mU8QynrfNfrsyQojtKLiIQhFVsJuZAIxSxIPm+AD2J7fwVvIe1dGcw
6KeWjDUzaq6vhz3QHHD2OoRGOj9Nzd5dL0m/XOGAVtOmOylhKINt1WHxktANGpyB
UEIGxQIF+z6tvPJ7CS3bUvb1AVXvBOSEAJxN/5a/zHzAOcevofmsGCfHoEjg7Cjo
2Qn1i+Pap3xgNO7zmymB4j00jysA+ifzW+q0HsPi+tzVa+UqDQHvNkWC6Cy4LgE6
zpsaGUmoRj8lZUYIbcBNEo3wCDPeCwIIR/0TipX2Bc5gJP0pdjXoy1sttE42NH6n
JD38DwP1c/cGDtOgcKplA6n014OjR+7eQ0zB4l+6FNOJ03ViUjrhpvwUV5BCqlDb
bmhlD/KF0nBKtzT1rBZWnuOTMjecl8NuBffrAlRMSiSCezSDsK3V3LzbRtXUMEjY
TB5B3W9Ktrmz9y2w4yZgZVMFzulPoybWSrY2OustLzMsISHIzgdai5Bc2gCGUAUO
H+yVRr/8aMxhav8RZxdtpYVLB957cji90UukD6y8GP1yITKopZEDYTdSeWL1jJkA
9r0LECZUhFRt8hnaW9m4CT195KdcPlufuTGMetNYoBuBdNtPZELoSQ2sHrMJS9eB
Fij4yia5MHqrjlC0fzW/5DQzKv+dmJbXlGvCbC2iFs3tj1SLIGCrsun2rnjn/FEc
y/GsyKHT+2hrIkgkn695L34G3E86rbjIAI5dMH4OUI/sEpsWEc57xdVwiv3b+pWI
HW+2dlFpCytbEAhzssMAe20fln5yWEm9RYcG/5KqwcS7g9MJ5fjiFoCfsPI8PO1y
uWqlDKuhJuKzoEzpOeBGRxbWGOL5rEAigd8OWeDMdbvgv6NbVNgAirPLa7hGRt+m
Fz4RgMfym4UgF6xyZxa4xYu4+4DYYBGp1QtCwwHCun2R9VWQDOuz4WBcSHL3d1q/
WXT4jK6bY/Ib+/HHQBxckn+wia410G9xAB6SWI5UdU97neFpNYhy0qijIXP1IY4A
g91KHKUXafSjnWwqUm4hVSDkUsNpZsD9G4ZUBAtOioov1oyurZFaGypOXAI25fXa
X2CopXmL19erh/SEcXWwnh1Pasa+5IQQ5Gwolp+1t5qAzO9aEhnXRw+POkbjIqli
uBxoGorJCYIGzgWiYleaTGZVeF/LbGz4an142T8RlKKcPxjotXOViaPbzFHZh7nB
0xDCTnh4a3ncOUSdFWfqWuuldmrT+QygIIzxSkq6x8w3VzKRkyzO/Am1Bcenvqn4
l5NRFOZD+gsVNrE3IHcQght9ypEtmDrRkb3dOKWWBkWU3vCbAdhQwdb0GSiEpCGC
Ii1PVcOd+AWQtWDVIkS3/jUEUDkPUFCso2Pj6a6fMoyBjJbL8uvoykdlOip8Qg/0
Pv3bwLxYprzmJeKkjKpgqTAIfH9HKtph1RalIwWVjJTRJu9yeEyqBPQEnOC2HlDO
CYy21paey+tpNgCCGYfkKsJB2iyQZp+IALFftO3uYCqT12V7TWjfkH/vazZQZY14
GbqShgZKAJQfXH5dyPWAxUkD8vhRfse9K4idBpLJB29TU8eUoWAECOb0f8HldutP
6Fh44PJ3AaiqGKVJqikxs39Zlz5d8Vecg2bPac3mn4uQXz84kahlIfCDPzCEBdTT
XrRp0j3VDYvh8Sh9oefO17hcOxle6zq4abP+mnebZSMKAAp5sO32S2LFaJUSozNw
lhxZtiCJU4yVeA75UMCtPP8O711OEJH7upD1s8yZciPIPXBGAFnggO08D6QU8zGj
BOlaMOy+xMY8H8LONy1EM5pJS3d9W+kx2rDudgRmI4Fe6ulNXXXuwx9Urals4YCm
zS/TzrpcUpK0SZkqZbavUYfQhMwOGDDwOChcRB4MSgycEHRNOCtqss4+Z6r6KQxK
jDXJ+x1xFqVfvbGpqauFIE8wcynCmMuvO2ENviGGmFJLJmgYnX8lWXA1ARrETI/j
ymE5JjJUtoTfUuTd0rtUeRSr0KzBThIZHwKwCFoUbRMTTZKclvSWU7eGYiykbGV0
QcaedH6C3SEiKTce6d56NzMjwnud+w/LqCx9JtIS/fNFjLLMmwx+mOVwx0wR7r+T
xAmwuJgpAiqJIU0jV/P+OZZ3ELqMgdkUbO6M5uD6XfuptKIcAdTXJBHC/DNqz49+
1ov8wlVvN7NXuE1jkIHQ8FWnw5z/vd+Tk61dL21HZNwiEZiOp141N0av7Tj+Aqxh
pSY+8612Plrg/Ypy8ROlMXbg5cHeyJHabWZwBSfUgvpitRPmnYb3gBjrFAIl8Cm8
NemwBY/MZsQYeFUdyFRIvsmG4KYk3T2N8pBYYixRCb2vIuoZk3uhG6SiXBFL7E6J
G5Jzz0MLeFQ3OOEaghMNgCEEC2yzyyNSngH2h9/ttd6g4Zj0ufJ3I4gOLyPmG7JY
YAh1uc075HLpvCaRolWNgVmhCOPstIOuZXflEBYeRYzsDBzan4aoVfHMSAMjnrsC
Vitprui5iVqBaiq8/XeCcvvVjjEpSgY+ZKMmOarEuh4WJep/zT68NYQyW4VdgnZC
7v2l0HqFsHrH7n9owQOspaDNBPdo+1mecOCNSTb5DtE=
`protect end_protected