`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14608 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhBNVMbsl6PTB5/ApNH6uD+DV5N7cjkYfz/wpcmHBtutG
aGMTCOe8GY2IPU/Fh8AdItvayopufmQh+ov0cOirMkw3XqKzts4RGspwhBwWGN7N
4mSLBb/EgU7rUjh92HIIa2JpapWY52bGLNzghiT2QPwtn8HtmgZ/ddgeMc1W5xb0
Fttu2CyPkAi3a4UVMb3osVZlj5LlYe0kfYxaIFYziQLaLRWYfcV+czxd3ncO5ZM0
FAMWpLixdfpZfelwrHKTP2g+zG4kiOGjN79ueFHgFpZz4XZM3HeVaj/ON1IOVlj3
j8oqjdGp2gyLAABdKQJGqadHuOK57z6zyQ3Z4ZAUOumkMyHeQkdJtYXGKF9Y4fS6
ia9OY4e2DDmHjYbeOs8/uWzR3bqTPDg6w/7p3anYgbE8nd1QQiJThS/4IlQsAcpu
q6aJHY3ejFflQXPvPNpS7yQ/gkz1785i3oNE+Ky9sTPskcrjSearWnRsGY51/QCe
lqACo8tua1mQ1GLBBCGtt6DtYZ1cz0Ao6NyXB3/9KjpsVznmQk28SWU6WqmHeSjp
ikkfbNT2YixvUgZMS5NARRkxn7bo64oz5TfRnEGk9MIBlzFcy6iWXP9Td1UrybfO
SvtYS4ej3mVzZPL5K0VXLWjgMpSa6/Q1riXfu+YxtdtQ+xIGe7A5cdGowps7GwZr
KvgnHbJ3BOHgPj6KjV5uWF26cVF04ChggmAR63BGx5ywiFSvrNOT0bIAcwM3J8DR
mcCEO5+2vPPTnBc83/0Z/tt3Q7zAZHSpNh2MOGa4ce2fmwQ/v9LPIGtRgaIha3Zl
DN3REmR3idg+bz3fPTtdbJ/DArof+B2q5lWkupLt1GjQPvk6fItj2riBY36scdcA
5YjksVveh3FR+nP3j7X2mRrChukbcHM1pLejKcsYnBi7HY8wAmDLrrgebCyTAVq/
nkJfWgcRDQ1Jc+6QerGmzB+/5mLjl9DUWUS4x+ob5Eol0Ic3yNPXjrD8FPltOcFs
h0moMEK/iu1Esz2Oz0BWUrR05cYgKb2QUCXTi2wPWsapZ187WEA3zw9Lf3onuW0K
QQ/QLiHZO2RiRT8+0ulA+RvKiDkyulodsYBoVkWgwk2Q0Wct8uvpPwzAfd9oEWsE
H8AeCVgJ+fRGut7JEMGNX3uaz/3Pc+pBCld0P4tV+ofnngio7xBiEv4oZ9v5Nf6j
GGuAD3kU4t9xLkx9bWdNQFnz1hqXTYRy3s4Jqi2deU+CNjmL2AK9aeTTsjb5l3ts
p6eXr7gytCQbJMaNln1L7sFs9MdipLfCdoIHLzrNAVV9bRV98OsbqiOPwBab4coD
+ZwYHCgl+yBt6Vr0HXRgcPKb1N9Hjn+CLFKXPnjUswZtW3UaH3DT/413yTtp7Q+C
OMqiwHSNzdbcVfc0+yw1NRNyRyorIltXoG8fUdOO6sGv/8630i79Ci/FhvdE1l35
yHmDuDZFl2xAmL4ZZfAA5AjEauFWLGk6Mxzt+3IQPJRp2wyBaJtZHEG2yA6s+ZXa
dk/EX219lYJVq0R3+Uwmv27+Wsmq5Osp9Dv2IMJs2F3PAcqdmNsQmm3Kbpo93QY0
8JxADe/pH7dpqEbKYfBGAtlSaZtwEBP6JDqj/BU5AcYxzrJiQALZ94G40tfn3wM2
y+1YaYPuOfKqvkM7uCjUk/CRHgpErIEAYvXx9vdzy3IDMdS1Bf03ixne8zrp2gOo
yklhX2NAvYMyr5S9Ndb1jSf2FVBKm5Sq+cHGLCNl9SwwUZSTl6CBDxKkv/f2sgbz
fuQZlpYtoN0JV/nf0JViT6Z8S8+5EL1mNW/j+W5CKn+jdZtFTbew9BWWr/5xMt+h
CPRx8+26XtvWBYw2wv58YJaarZ7T0MQF54Pc5pKfAFH0jff6A1L924fPjICJ1wY6
2m393/IRKIsWR76+klCN9+d7engTDdefE/Nl/daxspUfeEpw3KT/00vmXcPuKQH7
qaL8D8dAe8e7W3XQ9460jl8BqzpYBZg66IIu9FgRl/VweHwgAlFmpf4+iKAFyz9J
9MFGVNT3MALFrrYKKKdmrPBIuu0wpWANmem1yWk4+sAsiqEzIQJCRnXtnKaxpdu/
DrhmZlxyIWac/a1bV5YX1vbghT4xykxLMd0XJNnr7+1gcZj2opouKBZd1yohGjVQ
R1XHdNUlwA2F4a5GSgBnVL3nTWbsd3dpP7w2m0pzA2IkKE0RmzIhGYPjlc6zXf6a
F3v7lCJ3+gSo2L2VvqTnXzd6yIbvuDt3n6TiUUaVi32SAyP3ad7h2AE//fi2niq3
rpOUwlkiCbfvwMVkb8qBgax++G5XHkz5MEPbTvOzyTH02rt6NNJqlEW6+yAbl2+I
lG30ckg7xWp7saBzBKcZSzs9VEOKvEiOid60XGNqsESj+TFC8iTQmvRVvToWCc70
1J+V3MrG3osmXrHlJhu9OQc71OcQ7OSqNKqwuMk7XqkLTg0Y7W42P0CxiY4LB88i
WbeyeIDBh76qM2uhjnM+J78Ft0G75SMkC11iLBciiU5qmnBYTmIecKHQpz88dcyG
AqghQRttZX95LFsJLkOYmlaWJzovrNaFV2kAtHtakzllKY3BEJZ1zJcJzjoG/RnW
j8Kqy83qxVzgBVWm/eoZ/8ebjE5PLfvCk6xMLSRJltJKv7igNv9h1ILdpH+GiB2e
0VO2ZOmdUawpNwsz1SDQYpfi0i4D3Ww3hojwEgo/tejzXOXwKk+4qdcsZWvvVCw9
c8yryhQh7yjU3TlUr9kYvOLBeaXcuzXv+h2f3py5gGMeyVda5bP94PTSdjSHroqZ
bhCzcsYNHdHFBkwKQnHfO4fCqv/j5caNTrpfLSwHLoU7HycIgfZUl5z8w3dPWwiF
z7ytaBLMjh0pjfzeuX15lTsFJrCW5i3JxyOwCIQ/awALOwKfPcgjYHarc3koI7qI
Fw0grmZr/0osZg0NU6LGkBCtMfL1uEVLMrIlfHoyML5Gbj/WF+wqHRz6uWwmpghi
RNLYjBZcY5oBwJNZcjD5QMClytG15r9gN1BLIwUIThy2U9/3Ggj2AqkjdzFRjwkD
TRkW4OgcQxb+WSbDf0+E7qUZViEy08wjDg0GJC4fSod6yvilk1VYe1z4AFoK7Yy4
g/BuIVplPWNBqGp4kvfPhe6w3xzZQSblRLxCJanGD4gh/f7Obyd544ME6linCrLT
3g6ZT2jH7Q0h6DTy91pcGqtSZCfzX02xgIUguwak2jLoUe9sJheaipi2WkkDYXK8
g6d7BGBxFg7GIdCOCeK8oHfDTr/si2WXlUYsxZD448fNNdB+YWCfwnXL91TPylNg
n/cZVoaDhNPhO/W0CqZRJqa5VTvB7EF8vrfXC1n2o8KpwtTKsXr5VmbcrD/3ipLX
iYGCCW6vUi7YFvAUgLXQquIKYGVtMtdk2kWa65zNOdyaW3SpSmc3z715uxqfJ9sT
hVgUecKALn9hkDrIVNi2d2yZ7Yq5TXn+GKhDv6+l0oTcTA/H4qI99bboo9Bm+vKL
7T+cXXU9hxOTyzqJyBwNeztR70GpC6Rr0ds1k7WgxkOv/mVl0NlXsbzvDtMoW+Bz
jI+QzMuF49hrOt/Bf1hrNFus0+aTsA5shqcuSxS0IMeFqccdDBDBktvqIZ6JJLP5
Nr4Mj7Hc/2wm65+WBSmeAKdXNSycAsaouoPFJuGlxYrLSUY9sNqKtJ1taI8p9rLx
+Nk5/I1rjN4HUdDxtaw2BP3AdtQoqBFj4e1Og8jE8m2/hVhczCvL+7fWDWFBkmM3
q8MgJBWninXir29sJR2KdYW1pOvvJKPcj4ZE/HGcjIyWEyFFVLvDaQdJUuEaXfDz
fWusyIL6c3f7qJm+M4u2nYpByfrnNN5CIjAFYM8q3zoESTh36hoZSiyAUcYwtd/H
BmY3qdOrEHiqtab4EhYSuftoVQfRiVfLoeYI6MD7hzvFB5d5p3mEfA4kCb+jwV0H
3xBtoSkEyTYAqpRMAzFeMNDcI84jJ7pTpwEPTTiEIC+GgSPad+Df03X1WoPWES4e
92ckTDcZiMgRIFJwfeJLlN+gpDx0faWZnjwEMgXUscdJXactxfL0b3xCA+QOI7El
V2Paza7NdQKL1RL0D9ZdhGtTCSSBq1jw5nRepVJ3xdqGHUHZvRiopYTw0AK45AL5
I94RgMoe/niIlrJKYcyArh6iA7bDtg3JKlfuOs7K0QYQzWmrnITJAeWJTkTnfyfr
bMrSp0t2X8Jk9aoKp2Dz0sWHSNShvHtaQNh3mc0/TilnwwQgWFqGq13VrFKf/D2f
gR3NWoJ2GCkxxM9qY8C8f8PjAWvgRAX8p2QuD0Is3d3zfccTOzAyVh4X6jI3ZKz3
XR1Dhp45IpOJ3T9tUgcsHasZ4PZoH/PF/qdZxiFWtIQw4L8pYUXAx+9N/imCKGTq
w1Ka/7/CCoFwfsms2yvNp3EUplHz8Nhmh8Xvdt5WZbRtbeBzKmlhyEhLDNWTWpWR
J1o/muH4HLDub0mFGohWr4/oVbE++giqxG8Kt9slqzpMfWa8S25YC4ISGg7hJ4tK
yCvzzM5F9R59zkPo+tQAdy17jAppVfWZcI16kWjSkQ2hMxO2MIQLF0hHhIsp6o+Y
Mh2KUBaWDvM/eK0VtxEBTPsKdNbYJCdxjY4Y6rLnPWctXWTWB7Gb+Y+EhvSL3VfI
jwcOISO5pyesnylPOBnURejuegipA5jgl4hnhThdQf+T25tHAU++sPmy7ak3uBBM
+OXh7qBOhuyezc1FohnLxmeTV1nTz1tCDS6YzwGwavuvYyKm8goioE2HtkR5I6tu
7T9+EW0ehYfDA+upxyg9FMMf/bCc5MspS+9ez4DNkdMDHSCZPRFMeCYBKJq8c156
tHLovU9d4iPB8ywTubyBvKCTnBxoEdY9E/Z4HlPHAnmkjQdCZevCe/7no5y04uM+
URyFc/DfKTpBmsRqNpLIbnfAS6I5IrMJlyhTu636fe8UqHRPi0f0xFxELvpTskt4
rbYOAJJ6yEvEsMkmHTunv95Ayo6qO/5lGxj02XOF3di23eY5ywXWFy0Ax+O7HV+U
QBnIAYqViPY3njkAK5sfGc/H2D9gZ8375x6mibvhQ+sURB4qWq4lYzMZ2nGe9u+e
9TtzhgbC01WKyQ/pBFahoG6AAwGNGi6TXQjg8/mdcdT+EAyPIlUFeBzBEbzseKVu
wNd7OjqC9H675faTwXOp0IQwHPEfTmgNKTDoZ+2odm2bEmzWfZwL9SkUuQQQZfSS
X9s2gDERpxUEiE453NmmSMuTlppGvFBV6tl7R4IIZDRO98BBXYnV2TYzayFtRRAd
+/1kjsT+F7SnDV6Lv20Obh3lkbjJDyn8d9COy6iapJegsa4SVPK40UOVI5STdGxp
acFXVqwJP4c7DmzNhPxqNS8jd2CNKzXBiJJ+y8EqaISs8LnsHHbTKrBnyG0sRG17
5atzGuqZAONV88Na/UPzbr5k5NBc19SY0M4tu5QYqcwz/3l6is3TCFL1kKyM3mqx
X+8/4Zp/caVu9mliYn+h7ZZHkZwBdRtW8T5XauctiUUyMJl/3TjgBaRx+npPuKwp
FydK5Vs+7DdPzb1/n6Pjb6KymWjhyzYIRnJZu5l5qnTV4kWYCFCow5V/WTbXaziP
OsBPJ7YTxqPA/sVqJxqlijAnT1XaBpzZoxdNTnIx1v9XMtgniz6sP8ejhi9VaNKb
54YI8UB1NztDg+Y4sYsx8JgUY2mFNsyp5AuAtjI6h4N+Npkey3v005vWDC/kCtUj
GGDT8fP7J+/VHA2OYuzdw0+551szsJYW5ULBkV1WBWkCOkXTlO0kP13rAzApBlsv
NXBCLipzTCJ1OOmGfVLOg3XTdlnt30EsNHDdKiEKOr3cojWevl2Pa7I/mELk17w+
1u58IwjM8vO2TTULCO7meWiajEo6vvJXcfWc4zrFPOrbU7919s2M+1xquZfeIO/0
qaFScV4QSdPMDODkTij1GvOWyDnWubQOBFbKPbvlvazsrA23sqxV26GK+K6MVgoY
QpBdVsd70fTEkf3O3aHfah7Ad0VuxL7gElZlEVuOf0qLPx1aKqPqQg8m4MFHjsO4
PHtcwG77ILQdKuPFtQgSyZM1/KIF6WM1GK9WnN3VUHAQjYMadG69XnBEbBKzgfwk
XWyhBZJ0VGcH2bObNwMfvM1yJ48veIXSywW5ZaQ0SCafNUdHPN5My/lkZHJikfUG
KCAA6OxF9M9DeBMxzh3oSDl5DUmomOkdvhOqXssGPBFrt58ZrWlKHyCbY8hu/r2D
HdZ3npUZpYvru/jacYlQzEg1T6lV8IwCE2tuaBJkxdT2+x0CNw//QssJTbrDZsFe
dGbgyy5KSMGi7BXrShYHhY3VzSgsUxjMAAKwWtejQ75FeDTwxwMxtEjV8opQw1f6
qmguBgjPqi0ELKYcQN7izZh1c1crnrvVRXgJDKosBsyaO2aD5Q8g8wthThsxjsln
iBPQ3sr2HMfoDFAvg5yIT5OT4QFkEwWTQ02/nbQxjsJnspugBDX0wrpI5VET+VDL
xEgU0IkrbwvxhOu++JKzfVL+ciXLvUt04zLcwbM0JccmbHIEgyIWWaxoNkW6tE/3
sj1y7AaRyO4FWJJLDZubxZM8Pmr3ifHmjUxn+eo3HUK8fE6K0ni8yVQvGHdX3Pew
D1zGNkb9zfFjDtfO4Vfj2J1JeTSMEUTVFOGc5lKtopodVrUJbpsMAUScaX/bbm9U
1GSm06fGZ2/9a8qblBgRtQI/XySCpcTFg3QfDF979e+QFcSEEmmowSFfGhckasse
1cPFgmVszz77H7tWZMKp3ggAO/swkymDGFVlh8K32Fkg2BKCJHNzWNX2k5aJ3BtU
kj2I/G7qWWt6wP2E7E2SJ6TmYee5az1gx9RaWrJis/rlGTEjFfmsFqiqtyvyPgiY
Iix/HXi87iuhx2d97ZDT7OIzc9pfB/p6LoARnE8dRIJraw0NrwPOosegYPodNm4X
xsFYZ+Lmlwb5vQfLMm57qA5u+T1gf1Cu+wWzzMrpW490sq7O40WAr4gcKt3oJp6s
qmUoxF3GALZW1hPE3Z+pVQcX0F8ScvRoQEr9qqUYww3ITT8Rh0ae5WDrbcSEd4qi
Cbbe9li+hQXE9k5iMV1Uhba2JNnqtGcoMTqiSaNjP6ZZ/8Fm77EJXcPk/VpdzZfj
/1V8gCtBuGYbBeWvV2LDaAXv+w9KFM0sN1Tpfl/TEjZQQPKNqVbws0vd6r+zo1kq
kp9ZXujbHMLTnBSh2e9MKbjs8oaavQJ/RpbtTHkv5Q43NUl+1H8Z8Hg247gxkZPV
cHgNixAaD2TxChWD5Mn05pxS8DPapnAgwPE9zMU+0rhCfZpqCrz+SCN7CVEPQi40
f4XGMBSOZZGp9rtkW8xavPBvJfD7qu8Qxk0PuWgSvFZoejHjbtbnGLR6d2z8WTyl
z7My9PH4I5I6VkPQJCt4+DyhhbUdzk+gComr+QCpH5Ep1WhzmR/5OljeHguLJBAq
jh1OzU6Jw1J3OUogOcB4WI70c4W63EeXeZDhqETXugPi2R2itnQ4njvyBKMunnko
ey1BLo1RwRMctIH323q+43RkBeaQb6a1q0WTM1wGD72rdnNV93cGHa3o2wXBmVBz
nb6PxjPjEmtHQF3ZUC6/s5KobgexbilGkjEB8KZ94wJoFDTKgLjiC4xoPMotV428
pH4+tEdDq8r2XO8onLKEV8RhBn/zonDQmXGp+NfU0gSgJPZOijiRzbbK79b1kmlN
Is++bxH7sRO+S5oREtyITiDxmQYJZEYEly31g6iRmyBhaPCY8SZnVijnCN2rFQU9
imGAtBDTr7KEtJQmp3NnUDI1Kspwzd8lsCq1VgCjUmUv7GIiJ5MkHaBH3yBkMosx
imQvT8K/zmR51tveIOtJEz1yoq7cPpp2yAZ6I56mW8dwrEWr7qKaIQhg3hQR0YV6
njX5DPW0kBboQxBNnp9vTSM+2WVZ9EtB9hIQ8MBDKpquwHt0Ec4Ck222r4rv/24j
16+oJ6VTWAcsHts8mtSmxFUtztVp3w5dYKCQdjhrPezgs/3fg2MsWHy4FG4nNGE+
7/n02vn97/GPCkX3ir+LgcEaW+EVUJ1L5Er8vGj5YxflIayktbHMJZWzpoGPIA3L
1WGa8Olk2RBV56odacolEUAsebe2goDzUm/VkdzuNkNlaWQnaWE+9McYow0Jz4jI
g+wdgDWUgt47Id6WjzCPw0qmiN3HOf7C0z0L37Bo0O8sz2ffdwwwdk01ojjhcLdj
EpAI1C2vw+Yi7DK5G7Z53+in7fy/BVB6YJj6MX22+WZ4M2fsGHWPXD4R+gy+UMRH
oDoJHwUWUT8OT8mmXAlyElHKJKmBV1uW6fAZ3EHlomjaaTsLSECSWxBMn82GYtk0
BaQD5QUr8y0cR6V+rwFye1qqeBb/SocqLc1esF71TglAPhSsE2EfFTLQ+W3BSEkx
OPP767lxH9QNio7Qswhv+PvpMY+VqshfuYFY/pxXGP7w7ppI+zDw5Ans2YSTHYa2
NDvrXwu/m4plZPvDziqS/WyCsLV8CgzzXSgmDTU4S2H+lL8sTT18x8Mq3qapWGDO
9GKQxlP3K7ZFMcWnI1DIRv0j02zkbM0Of+Y0tL6VUFcTbEtvbupQgW1CIQcJI1yM
K2oJc8j35AK7bOqwyIQKwWD63CofQEdgJsXt6LzrtS5bJ9Cfz0O42Ru9/NBiNsi1
MSdsEos96+nGzogJ+RouLgb+ixTXeTMzCJPROD7GrVoEOfVDgm2FMktHMZTTr9Yj
sZjbXoS/PPH5kJfXVAqUXsqMhW7Z7xml9LGqREgj5/CSlg4kp1Oxb6mBCaEhyPPa
VeZvAoqCdCLj4MHYw2MqAOX9sg4tgOFCtOaRk+AmJ3PU3o8TV2f8EeIHWu7sf+eg
PSHntz9c84OZ++QdteKP+50vehigJ8/tp7wNzDBBstJWKVTLYYbph3bfmfKkI7/y
Gld9fBxPZUWIP48cbz3aZ+83q83rgwtOpXL7IEFH2sArYWZ4+0Ly5LK7L6TenZRG
76Z1IiDSMyzyMRrO6RBpafAfoizmp5F0LnRDiGMjs1YjwHtTh8olu3kf+NwsWhYY
aFn/Rf3AsNm5MxBa74MYi2tW2aBM8onxwqJ5PgjgyeEJFC+hqe4xwWXDVNwL9wtX
DMzZ2Z4Xsnpi+IzjMl54yPFkKVZgyFfCAQx5SAvjQ+kvz30ru6Eou984+t7v3TnD
sF+s/81kdj2K4Ysi/o8rQpyWjGHKDSWVB9Mc0edCw74y5aZ/Zv06OAfDp62cn07F
kFswvAvqBxa3Bk726bl9KZw7tLSirAEJlTux8i0N8XG4JW03aHV/41a2eC1XE5Ym
GGuZnaKh1BFdpikz+0z5/DvxX3vB2wVCP8nTzqa4+KYkBAfWW+j8fpIdd5agSIEx
4wJR3esh+PJtDN2G2lO8W0NaD5hdZWhl5yXbCs4ZM/CWulApULjYvqq9HbabTqXs
/8219GGPT7TWI1wW34juc0uMQYWzvldhH0yVNahAMq21dqO9ULtZTaD7a7bizshh
OOFHTVxWgMfpQz7mVJp9morRrfP0MfDrRg2x3BjkIUQXzOCjINNrrVRZ5Uwuj2B6
0m8oPoPu9cJoXPdai9OUxDtcYLnsHhbfISPiwHTxUnesDOgLlKxpHxkZ7OwmdFH6
kk4yz9TeyaMsPU/UaJcaJVyU5fLyKSEvVWYdkTZUE5aM7FDw3DgUPAy32C7VMJdr
PwcJmOKA6i0TcVlhRV8VCYaud8XET7rsYtrCC3I+Sh5xdyXo1Gn1fqqp04wFI3Ca
odZtjKWgpjPEW/GisOgX1NzOubxy+Ay7WKqWEsPQqea1PK0DsuJqQ/51zAjbQVvf
0W8ZLY8cBsKoQShx54o+sSP5LCBb3odvGECMguSU4lmTDiz/Wtkj48qSMMBy0sWb
4+lY7Kr4qT8WorwAd4eiHL1Kx7WJzJMEDQMm34nAxhu3m2btfd6FEFPv8J4jPKzp
IMaaOZYpzCDktd4j2SmEDyqLZzegbTC1tPnAsetq3ceFq0qtx1xNOQQdl/kzNh4T
UPoQiBQQQACCRUM6TGag16Ljv6Evn8S00yXxVqh7vnvL3HaDE43VKZIN81GFxcAz
YpRZ9uWpcjagOuuoRWOBcsFJexiXRfJM9ToWhDjeu/wZcKcslCTbcm1pkqYuqUDa
4dgo8b6LYayDIaxJoniTxs1CTe0XeRepWeYVrBBqdo1Rc9swOJY7pGbux5LVAFUg
UqSy6rqP8Crcio+BcMAsPdi4NM1406KN2xX334uNdNK1WBwaITSo/HyqFQM71NUf
SjdLPS2T8lqYfvvxtsPkj9D0kV8a4rAf8Id3DrkBKRl+Vz/fizfNHimXse5LDTIy
Y9LSgOEKhY39OWHNCsp0MpD20DX85EWocbxfIEMknd3QC6z97S0R/VnKKonVikfP
OOU86ktNxPNURj66z/t1qNPpCSHgWu/iweiAodG0e4mHtbkqkz2gGr8kzkcpmCbz
Jb70f7GnPUZ7N0bqXEco4JQqxESFqwuy5aghmOuyI+RQSF3/wRvOHN3ai+q2a3wv
Z/eyyzFzQPISjXYpCO34eHocnCWgSCBT/16f8OLFp2h0ugqZafoqEleK+APsnOJz
ErnIv9U+76P3EXdiT34VJnU6o4pKg4hStLA8zuEavRakCI3uJSj7XnI74C73Mlev
Hvdr+a2Im3dJ0xItpKh8Ka23+PxWwynI4Fgxg429HNGze3Gg1fAGRW29AkPEcNRp
83CB7HJVb5k24lkbZnn7C0BBtwrLKWAOkObIAjgUx10hzvRx9K72zKjn8hx6cF+T
KzpRxKdEbdQ4S48Dm16P0NpVeuMDgdze5xKPnoK1TNm2mc64Xp2hfmVysD5Qgh4Z
uHPjsmmXAx58DXpGCJV/lSa/3ZcA8V/B6Q5FsTwgLEyzpn+g8L3T21WMizFYf1qE
dcl80crMPFRa6OFts7CYOXp0eNEJa4BVw7Y4TsG7wfmj3spICOuHhc6T7MCS9dcm
LMmLRXX+zONFGj4S8R8H8nWiVfys0iLP6mjwh01B63SAYuvUjlr8b1vzpseXfefV
aZsl8LLFOtdaiPUCZJJfAyyRE7xeFM/+9OMaTkNBlWhhkPCTVixy3EbwrCKrWROs
3GNy0o8uScnWUTwOGy+GzARF57R9OmtYoeqKIF3VX2bLjfhl3y6V34iwd9tkYaXN
olEsFJNY1s7SfjXEjCQGUPhYY6FeisQ+DpervbnPEFrzC3WiQTILGqFi0HfrBa1H
BZaDzvyH8QKzlL8R7PvxGbmPyI0+79KJA1IprmGlQKGLkd1Fs1wz+5b157T+aqmX
TZOJxsJy5a1FGuYbamQqp1XdDSN3EZ/+IcPvH9+hbdo/O6j6su1zw5uxCvpnEu7e
HW/jQuQjqOMuoNU4cRb1/gpKUwJ8w5HjN+aOGsBd4c2ma0b190w1cE47Wva8/j18
Z+nW5AlgvnpacfMxuYCPgakIhpynvBCFvz6FumTVFTOB8XqhigMs0pNquliazghT
5JkfBkZQ1qmm+O/63fZCWj9jpT68/mgoh0QQXmINqKR0/OogSjm01AWE7wRzImW3
uAoLC+2ttuclOk73HNikjP1348Dlpd7OamlPeHg8/awKYMPRlDPcO0itKQH3DzKx
B8ag3lAScFEXvZpc4kOSV0mYEc576qkIHi+mpwyxwGi+MDsyldYu/NEHo1506L5n
6LLutAroBaROUAf7Tj3Ue6G3bSyaNPLKHUENm4WX2slh9Vx7OhpxWSEsTv/T3fNW
sUculd9BwcQPUY8hoec7OigM5L3c6+8kskPIpahqaugrBiY1nPQbhI91cOSmtCPl
UKYb8ClqWYnYHjel1rdsqrFPdfo29kJIEqVbCGXHhlDZ335SgH7rRm/UkBKyp/qf
qkdVwRLyp+plTgikt1PkHF4+mzpzlNnWHdgTzlmDX/IegEOOFbvRf/7QKdFM0lNz
eToAuKikiMMFuyLZxVaELz1ztZfWS1aHP2Wt4q/ArxSpL74GVocllSzYMP4GK14a
oGQ96WMwaZ9ieJOTmSzKUBXZh95a4VpVfE7n6J32GBCVUjXfbgYmMOaeZ/R3nXbu
GKazhJOCJJmGGftPnF9nJs113kFC+mx725IqdERW8X3l2k64l9njduXTCOqr8oRy
b8qt7rg4G0/INcv1ynf5P0vzsnzD6c8RrXsT3+N9zPOWKmO5ltTrmJTxCnuUfxMj
w9Mdswgr7foyNuYo5pRXpiaJgyosvpEq365ngNISp8Xpm9kb7n15cpX4axiDTs0g
SvmptJNtpwjx32O7JlQBZZYhlIk+c3Gn6DzTa4j4YjFHVQboHOdM7tGnlYBa5y7P
yN2pwW+uNh/jemPIYOdNs0LvmiBP7nGIq3HRYoh318duIxqlua8BB2/BfcOWbu7l
7bADHsi+evYzSdYt98xn6BF63qgpdCa/Frl1EwqETuhz0FvnGGzDK94+TQ0ccZ8V
kTvlVHQiEffiMwZKJQqTWychwjLOXSXw57Ot54Z2nMppW51rpyUW5JsdPeMgIR9O
Ywg9Ux3Mt7IK2I5JGYEatNVD+sbLqb0easmb9OA9yybA7OC/sFxQKfr/2ZWIWY+V
neIKi+XsbaziPD1hJqq1Me9wMcZr+rOAprYiiVA7uc8uJnysQzGHybUv0cJR50j6
2lJkhgt3Zy3TA8S7+yy3rAZB/XQa25hE11SAlUV84pvIyKbbQfym47Xpza0h1Oih
k9scWXOexjboCJDQZip4ZugFA2ClpzUCAxnIrxz10eouxacbJueEAp6H2DeC8Be9
6YV6W/pHJq2+jgMBAUc20NtRldC1Ldbnc5+qMUzmbmiUxnF5rGqS70Lra+wdt2l0
npUVRBzqo+N10j0qI+L/ud4Qoq1nAZjOFEbI9Nxo8jP5LKHtp+P87TEeI9ipe3BF
e7hIyXlDUO8GUHmykBPzuYKO0C9pRzfATV+65N8sxBXZwDj8HYyI1ihJJOmFGwcZ
eA1wnIsXZsmIlToonuhAUqAUpSdfdyVoGNCzJtz1hyUwuSQzmx1TVljURwwLx65e
1yBSMooQ1I6Rm1TJaWVntNzyhUGqXGJuh/n6S1KTe5Edncoqh8HcRfPkGJuR6QJG
KCkaV2PMayLFZTZqXgACOjAKHgbOe8DZIWicuhLAbKeHGlgZ94NOETm+Cs6O9FBA
GYe0UdXWcvoWSGezZvG5/qMSGBdW+kzEihS922wnInHUsDC7AkmpyhV5XLdR53zk
/o/RgukTB7hqmADnGVBMLeBMLCUxIjnan0DkVBVdxpmGx/n81XRtueH5leVhGpkQ
3cygTQo4mqcAp8hy7S/a1pc10tfltE9nGIu8sbwaXtj1Dt2HoqT8F+5mK0CsFy8w
p2+a2ljBB6Jskuox3dxHyVjYXOgtBdfuop7CSeKgL1vp0b4gemBQFCBfqJEq5x5/
fAM5gvgQuMxNshiVAccmf7VCXDK8q/nMzQuLLFg68eSHP9HKWuQEn4GZIlSNvVw5
Yg6ybz1iP4/zwVmlJ92BnFICHkTcFrARsqMrIDhNzZJXrbgB42dIhAVlZMwb4V4+
xSnwxJCZ5WV12i4r5GroqTNel0N5HpRxwgYSG7K/QbOzC5JDLbY9bRzTz2vuczKd
qVop1+LSTgm7TzBpg/bD2TmhTMj7fkVe8Ibqk1iCWrMDxlQD8POtBe1tLBvQVhk5
a2E5iEMEvBQCRe8Mo9DU1lHc3g6fghXHsU6w1f6jWi75R8YqXBKcPbM3TahpZxaw
PbSbd09sSckMoL7e2waN6qzBnRahdqwFXGooT+LKdBROsYMMTCN5ZkwayUlsht/m
SqHaIpLMBnH1ZW0JPGvqQJN0vgHwYrmt4cz/ErCN6It3AMUhRboEc+pHQnWcDHeP
F64Qj6ckKTUK4+LnmqBQNo4rlcqM9Clh0OOrBohUnR8Bgng/7TTGTY/vb2EUccSb
AUUo8NTSDtuqWKuqjETOY8U8xS+yLS33kYF8D3YRwyjmciLXjrmTLx2bm9tzReBY
lqS/jb2I3QAJJtXxuRxUZGxuzBvZgwDMAFoocnauS/buH9OAVp0lVIYU/umUO2Dw
CqHHG8R8jrKRpaTcE3ew+HEXP55yEP9RQS4W1ZMRzYp2FzL1BHmTJyxNqIpBp31a
/nkqu267Z+NTbokkBI6KVeY0Wop8Ix4Y4G/SHVb/p34PqDRpbrIBJ/eU4LWPcaVO
qWFDxL44L2i9qcukFtoWfv2VpNe6NFoezBcxXCjna2ZOiGSJtqTXmjXErIZI7IQX
ok3KDNarHBIo+CcjywBA5thcRI9FZ/yEcz/OwpxXivTHj78z/apP0F4inPNpw3nb
fNxhfoafSsKqc+TEaDh43VhMSdA78xAZymbLK5mXTHvFkg3KXOgb7FM7JEng++nx
PlxLORy+3lnIWQLEt3MXBrI3Vde0qCd10AtN5O6mBWbvfXlRR9ukD7bmu1AEuj7N
uqGbvmGTjydHw8mKAzl46rA/jkjlPMVdr8S49IL84J7uaRvuceC+vNpmOWZAvoiK
6Dkz6zsbyy7C2w84de7crRdYk4Sr5p/ND57Je2ucc8cMihjSXPJgLU5CSR+zVZK8
hBiCiuU35th5a4mrzuaCfTx+WGCeCLrKtMF24E0Gm9tkuci8d/9qh9gKOoWchibp
GbCMLWcZnk/Y7h23nUYrBn0vrjXzOaZ6rY+7yqmd/9XKbFwkJkY4wOoumkGO+YbB
/VJpsxb2618FMgB3/DKhUyZb+oXI5OV880pXt3gRxwgU+kdNpP53UR0aQkE5Z7N4
Q023G4DXrHPPK3C+D8P/ih9MXmFZ24bDd1SoHJBbdwGqaNogjsV36dl6KOssy7g7
6ZkEtr2cOoepSS5DTUwBXDNOySt2kzOBxyyuuwiuyaCQj/7WNCfltpDMFTqd1SiO
mjF+YFYT/ZWNVL0sciKLJFHeZMgYWq0Aqa+zopQm+Nl5/DlNtzyAkMyDSL2hCEPi
WV7hHFO4jlqJxZZzmSd7yw4uE6e0+x2Bn/2RufGmZDZe4huzQLSCeD07ylbUb2yR
Jd9swgaHlXQfgbKzldv6UsyJdvY6kjCalDC3SYmTDZyHByLh0ZmTOik79gc4I+kG
WftNktq435AwyxKsRAU+3GHlpTeJlv+6+jjhC3vWmd21v6yzCHNqQfSSYIKVIOP3
tF6FKLH5nsgTXAW88Y0Ia6V8moceEG51WPC7HE0olk6XUDFxlxpTOZhCFC0kMmkz
3gk8n17FKZ8H5H4JMnErh3iUrnoy6J7YE/Cj9yCmbqR5wET3ANorhpQCcuKMHUwE
BzQ+DyeNe7w59s+l5ZA+FDnzabF5zIkO3qnKtIRXdtoAe11aTvIMwUKzftUhgaxX
UTxpDmsrJVt3UiZSFJGlGlBklLAgnLJqmvYxM+Fm3KrNIK4s2KHIYor18iH29o98
7rOi9zAYAouR0ofNVNIoj1jhcXTKKaU/c/ajzvNAbP826Dd6RAMoas3TCy6QyWTR
W8bWOFqbpiunTmO77RN7e3x33MoWvotRSzIvCUui8y2YrFivODq2caOe+3nAURNr
hlKLuhZ/VpRWAiR1zU/y6F6gucwfFWk0eR9kZDDk0PsN9Sei5wSiII9G3OwdvpMF
Dg3TL63M/GMF5Ombq7JSzdV1yZHTNNHNRNuiMMRxvcTU0pb/EdkysCbeZXyW4sxL
ZTPXG6zTSlb9kwA25D2npQkBYVCEOkDpmdoMSGb/Ca7C92GFDyiC3H+ZKsaznrkv
7u5Lu4ymB4XCeIAOrVo/iJCmvdH/uDjppPKbWQKSMPq9A4Q50ARzXujdKibHeMPj
2DzUmoF+IO6zkLu84FaUpYTY8+E3S6a+oWE1SkPgHfUofE0dGhfX/E1j2jjzpoUN
GDe0P3IoFpAiTQVabDueJGoPnTCy6pk5vE7mr1T0GWu2rWrnu3Y4CqO/1YN1Fchm
pJQN3mOAGJOXPJE1YSOvBbe8lALagfgE4ds3KKSMpagycf5XWEGO11A4KAuapNAy
dzagkkK4rGUTUiEMex6ajM+Vqyv9TX+kml5wW3lGFZ+OtrPKgubzYZKts2YORHaZ
0ucr6nwfUPp7XGVVYyEv2U5TY5BuagwxAe+QNeLGCslbzsXfVz1GYhBuCDx/a62i
5jGWhHcZDsZugdHlfs6YwPB3Z5mH4nDIzz8r5oo5JFA2ChrG3UONTxMEKZD20S9r
i1zsUNEkOt9WKnegU0tv/tgdfbvQDBrNyUUlWONyshx3VVsNhgD+BnDsS6zLLMfL
5OBIHc+fnq4KAtzgnmnvRwyaO1LoVavqW9dyx3GZit7esGicntJs+ru+r5awJFjl
GcTqrA4Wmq0+id+qSZSBnn3yTtC7ucsh8Zne2MabQzFnxUel2xV6dmjEeSJ0sDsH
XyMjk1qHnnpjmD5xInqxDRPVy5MQKfo8NA99x+owWgEOOxQiIDlaSbMK8WXZ1CLw
/OfSyTPMkmPEDTyuFxXaYhXqQzTk7OApxfUiLdt1pd6drRNLT/BnroCSSCH+ba7T
aPxuPZcI9AnUOqslkGOQRXCf+TZF2gBbIQl9bXsTuTOWp8oki2d6Dn49/gazAU/I
8pg5ZUidyi6YYlmg7spwtHWJuDHW+MHgZFsaaHsy4b+2SUxe6pSAlLzyAo2h+r84
RmFNsxzVXu4vdjYPYdgnYmdMUYiXu+CksOdvxZRyihNoQqYH7zxCBptoNa7A+pws
i3piSXx/l4ZcXfAw8wCCxjCj9TvR06HQMpGgGKs79Z6/tpfLf3Sc3PouiAhLiMQs
RXiEDDM5TbI0QHk0gh77w3RNLj+iUJ6WJbQqYjjM5oxlAU0G1AID+aSji9ZdYXeU
uu97uwB7Pp7S5KYZNVJXrZ25vlH6wCA9erC7L3XEaQaPWAk3xouQRl+n8DZJbml2
4VGs12W2h/PSOP77xC8+bA36/esMbMmzdga1DNjinEbDEVzhlplyWVSWa/klJLKH
FCpHPbFMirUL3JVwrZMgK9SsP+gdcnkKH1EfnObOhKJaDX2PR36COB9scNSXc37J
PDMAjJ4Cn2NyYgCzBUgjWSaNBM4v7RE7V/wFskow2EFIbEk4Z8UBcmlUzfNw9XoR
JloZjW0DfcvVTDOAD/FZ+54QJuGw7Wqe2KkyXoUfruCH1HR3MDa1eDS8BWxanV1W
tC+xADKMRgMbgAreb908VXYjGUY8N0v/IiEI7iRPzL+9eQg6GyVdpScziVD7O+aK
jkvlh7a3B9r7nVbDgMLsBwkIbbCTC0zogGJ/2QEh59s1lRmRLjh9RCKLoThohoOa
0bJioB8zJhxyN0XwLF3GqoyEXfuhk1+qL8xcY3U+tvuTcfQeXRINl4kke694oJL3
+wkOw0P2Zvg4G5y4/L0D+uHlNolwyrpiPtQD0l435oos0Sj681gxpZ9rP7uyqSTR
YXAL19qys7CKwAaFlIHfjCpG1N/vElT5QnUbjM4YJJekxNx4ZWo/NZ0Hq1QxeyYh
5wT6nui9gQIa5oDBTytSUCGLhsrZujd/9RF6jBhKA34OQCMMuR97v4sw6qcSoaod
mMlnMm/nU8TkqSp531WOuCJzm0hQTUKyri8ODJFZhywBLGsiFCnj1/o0ZYlwNm51
KZC3wlw+fipOJu2pJXlnQSI8W0C4ZRJZCaob+gx+cKFJtzUIBoGCPbNyqRFUrGXX
EcIv3TDatcYGNjhnmWa8aMrEdKUHOXyXwEUp0F5ytQx3p8CoVdoDkq3KMZs2Kg9W
++8Rl9tGp/2AxdViKmgqIFKyqQLp7Wakok+odpvUV5tBFvqLIe2WSDmts8qAm4kd
txPhEyAbIXiF1VtyXWcpODRaxqBWqwxPhrWLQKagnvH+ZNfWx8giKjG7Knb9niv/
oQw2Jt9T+h/0Lvll2uCU9BdZgsojwYO8ljEN9I2vKedk+kyn4EGfnSGi+s16wYKP
KgIQR8bckxqGR3+5KWn8fvzYr/uoBWJReSOokTIu8nJTP764n6q3CRiFPVNVoRth
U33NGUhnOwTWVN6Lx9J9quNcyHJuQv1XppmN43V+5zGa6vEoDr7R4UXpjWhszalr
lFzLDiQWHcmBHBHO+ylDYhw3dsIbHdKLooUuGmLr5Zv+/ze/QSvrOBRjttPvdb7P
T6w/jKoL03zxszNaPsEp10X0RGUs9+ifWoe1Eomu8M0sHh3dbHYOvtvxcgeD6I1O
RVsZTEx2//jheQEotoYaHl9LCk7ox+UWk4Nm0QVx6GV4HvJXAv0U/UW4PN6OaiCo
bGDaWBRzYfR74NxGhXyo6Hdqa3cjnich1shuy9YKM8QmLEE29ig/jVX/WH/X8kLq
lF6aD7mQHFu8w9w+OZrHObGOcklgmyT/yhL02dD7cTVJ9EgqhOaP/GKEJt8+5lLZ
ORHmh02ggOglSZPopdBveqkAlQ31uq2Csawi61DFrzzgHzLvPrgMLxX/E7djs4C5
tRiAMqCIWdqeAoH4Q92sIvXYYKK9r6SezGT60E3APAZnVoBHRma1Pf1KEsR8nUK5
hSB5vf0jYR+U/rO111rHxNlXYgevGW6g9vh5pSyEPnGOsrMU7qVqo8l1TQRjSJOe
KfohlionJOpkPVsLMGX7P6hdCWyrZV38KUAFusLhn/rlhzZ3z+AjzlhdkYN+TuA2
qokx9XJ1BwYq9u559ASvWAdnDzwd5fZ9yWJQt59dw5FQ/+mvjSJ+lzXvqC6K4MrY
oBt7N/v7WITqp6zbA4ees7T+XzaFoRFZVdv44wwmT/SdqMhD83aQCFIh4OssXtzb
OdH8+oa4flHGIANo1GQlB6mG2labLGn8Cb/ukD07BRYB4h8Egpo59DSYqvkdoJPq
6yJR8s1qNrhZwmYzvAkzbn+UYRRkEl++q7935l7XAgC2fPS2QVHN4F0cECCAXElr
yAnJYd/0I6Q9lJf3ciNL3/yxwF4fQM4rPdvjScG+CiOQXpwkKIciDqvfiztbFhiE
T3bOY2figPOGfL/4r1PVmglHMwzYKXigLhcZsS24DQy/ezT7DGPe25Bbfevs51+T
ivu9VoSbtLd4wzi7s2hzZhZw1e0dOydR9+Ed45C+ZzSOJeKav/+jUDUC+npg3a63
IzhKyjpkTqpOiWYpa8Oh0g80tFOozklWskj3MzmEaHbih75Ugb7fNWn9jsavfBIN
8QPz5vqXenZ1OfFiVuimZTGEj5yMlNZ4ZqNvVFw2QJZplxa9mNAb+7c3fGAjioD+
U5DtbMImCTY8DMjckZ0vp+YiKZjDWtzvRPlvyQu+Bg7Fxgj++UMWhWh53D2gue6f
05zBOU+xTmMCmfjL2oUJpq2HeTWgXHIt1Y/5XLcOK+idO+/YtQY8AroEudsr3uen
5UC7kWorIlJaSzXH4d/+cw==
`protect end_protected