`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4816 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0gQgIG1mJzulW1XOK5NnZR8
C8XqDUtXW7uOWTnSVqbIblwOHrDC/GFb3kYl7b/cVSQC9gqjWEqYWI/tJjtbw12V
xUJjibHCtm91BnTYcetncSrOUOEm49l+0aQFUibL2i6yUVUGJh1ItU9i3cXtZ3No
SrAkGWP0MEQ3TTKPz8KFFNyg4XBKs4kGyAWm8w93v2c/HM4gkKoy1vXANqNwODOV
jixwmBMuYVzjSsy2hlE+KqPBcR/Ji0roZr6LSHopjS3dbwD28eWIVFBvdUQ7j5rk
fHojexkkIc/sYMK0+PSKs3Z0zbEBfFXnbAfOoZ7kqYj0zvrbBycdRZVY/K7Dqupy
86ju0vovflRy5TfbFfEHJ/ItoapdM2EwKfD9Yd3AOnVLco2RPeuIdBrR8JLAV9Bt
iSHXE2a+/2jSWV5ElulJNY2U/vp+ZRrOis/H5M3D2qU19dOov53CnppU8pAuUGn5
L3vZdbUwQA1qDfrtJyOVuBOlrCxHmLHOfFRMgYUmitwuM72i2t/bmTLsQQAQbxtq
OGifjMQo+N5cPi2K1d4M0QuV0LjyhMU7HqxA4F44Ff/PkKehDQPZ9LQopkyYjomJ
s9Nj09lqPHu6kh2qPcB5eAvR2q1oE9x2gXiCYYeWorFWzPglptLjYsUhpbSVd2JR
9LU+GPpyoryTvT9785YgqlISVzXWkeqfnnthPL/Dw/sW44+EZN4JaLvpDloefL9N
sLvKRt4QeK0J1YvfsxLPyDR1/qGNUEhBvRBFys7d5YjvGYnbRbyuG0RxpOAW55PU
jfiCRuzndiVPADTENU4qkUmLHvz7I1NrEs/S0BibxfZn23+onN5tQcbXWagrwrVz
nrWoP3K96cRmSm2qW4RGj5OLQnT427fYg2IowsRt0euAyuqyhnQFopZIEySL6Wlb
8+ckfcNGEt3jaAKw/QlWMNKQ22c4DbQLeRKcis4wuFwuBF/Oiqum940GT6NF+iPo
nE18+4zmCFVEC1txbfmdLkakugXn3PrMJQNbVm0KPz8O6cehUJHX/iiAGDnCPSFk
nTypc/WrnALWslW6wRXYT+tO1MviZ92YtaEAfHT78XYm3ZVCnevKnzUQUGNkX1HM
i+gmuLhKR2vA4j5sl5SsJv58NhSjeFCa1lcd9f4VE/7jEW9/94FhW4WFJ5co6+TH
urT+YJdreRWbefrXWX2tgnEgT3p7GpVtYEf0MWyKKt1tZ95tuitROf1BjR33f/Nl
rUDm16uXhMu8UKmqZaxq8YywqmWsUqO2TzK15KPgmoKX6u79vWQozWBgN2hNvFob
pbm5cUAmscinMHxylej034rm9C4s/oqVjSj964l8xMHOXWfDHqiE7ayImLe8aj3d
SdBIT4wI28RrjGExfe6UdLevJJCgtVx6ZAlqIPEERmuYSBQphc+58+TO8mX0+g8w
mbLhpOdnzobhbIY92ygVvejyGJFS3BRif7f2JklxomuwBJ+kTs4EtlDqfbSUY6ba
aMbNN+3hAQ4k9ldBcsGw9+fq8d478a7WvW3jo7nta4DedwICk6ULQoADEtDjwtNL
2QXT15ftfMC37RqufcqvbHwhJicGSfPy07AubVtrm3/tFZ5j1v7x6pv4tlk6Bvn7
25difaor0Gd/BX9KgetNFcDKKtnkCp8z+qg5kB9TECvS7qDewuN9GVU+DfuEjooW
pHBD6KVEGq9Z+6ai5jhu+2xA/mP9ck8onhqbehW0co3Cj5ycq16T7ajrZYSrTKB+
9v1ksPzjG1KaKUOhY5zYCJ7KC7qEyDmIheKnUwMisYu5ebcI8LDLgHcUwnlAybcm
/AuCjGG6Et1ma88QpuqsSkw9tXYJ95l10p5lsKWvJj0RMwvoIVV+kaJXRMCJxd8h
c1Mqim1tzfZhJkFgVSxvcE3JgEPbHNeL+SS1Gc5Qcy9VCpp1X0iM87iLihyZyOIu
+QahgybG/P6eZ/wtMID3wiQZ5Vnnt7kUhovwj1r+nAPORoYMXwvAAFl80rQSs2I7
Vmnx1KCYnLGFJemucBpN1hIpgBLb3dwNWCTm7A4a9MOq/dAbkyuhQV7aGUmk792M
LeHwXpHWVnGEtrNu5+dtrV8b5QnNC4uF3G1EbJs+FJJYLvuRCM/KEJvhZ4iHWuGo
odU7qtB/RZR6bVn0xxYGIQ8oUqjeLVZpDggOW8xd1iPUiVgerSJvSthhJ1wI23Di
rTLYN0hZOiOY53g5VCUj0ZYCplRXu1RdEu2egq+8ZoZ4wP3GWy+SVOLbc7O/b88Q
COk5vA6+E8FRio5WbmUIfWIuirgwQzcXcZ29TKTzFygcz+unK3xDtkhzrWE84UB/
Jzliqu7Gfwh1HFrxsryxxrLZ7HLIIOM94T6ROJxuosNsq7KYjzaTl2Xs8t9xQR5P
+75qfdKaNP8aJVcME5gYm9piuD8toa63Rx0QmlG5sGGGBWJUsNK/LbvVVF66j1Ke
ORazQW0IJoYjkNlvmE3s00IjcDFDpTqYDqopwPiw2kuxnC/hV7AXJPZlYXxGPLXO
uabs+06EwXq/2IstS6kK9xknWxKau7g1uykihRbu9hbaOaEOeBmuM3t9sa9VB7LR
zdsH0v2A56OP2IIcm/aQU90qUcstIdTTxig2O55mrwDuAwDFNIxyRVNRu4GcLEjq
ZzdMAgUqxwyDPFaQ1CNPVRHuE09AjfdjwCmkg/loj80Fp+hruEFkwufqI1QEk8ZI
f9AIqieY2qyOrgfk0BHIJttJftbegnbUQNndWLFUHE6k3y0aplOT5P18yiRKL+rz
WAlIAHCS7GT1PAsQwn+JlWAhBCFWU+z0OLOEuEH//rd+3wPNQKrMFAkIfcVTpGWj
ZStjkdjEKL/8Ho8SWS4FqootNDRPgi97nrz3dh0beNl1hO0vTEEuX+PEd1b5ZqKo
aVgkBt95zoA/lXDp2frWfGwUmtujbEl8Y78fV3ZKuZzmIZfgBDkowW37vnbFYNp9
A/F5RXcSV6w0A1sS7I6arFITLQ2aPD+cD17WzSrdPIA4IfUdd3jbzKmm9Iz913Zx
ryIGmG5uBvPrivPmy6cfXGtbP55LKwpGlpKnk6MaikK5WO+YQXieQ17FKDhjtb7T
2xdsxZbaDgsEgs/Nf0HdX+Tp4Pi0ID9RfEORprYwA26Be3ALstARRtet5BhfJvx7
JejGMtE6/NqsnwzGX9neY/WUbtu/SvZwMUMXsBWJ0iu9E9oqNv+VBny3pTgyi1AM
/W42nFJ6NLAc9Dc6kmKukwDzcOnuMJNoRsj9vdTy7yQz1+Z3LOleRcgHAcKIcoxZ
cQwLb9jxAaqfMQEwg/lbnbwPLo6M38MG6NXOq24k0WodySHGcHNBTZsTKGAc+WvL
wtXSXHY2PwZPMW37RbfDujph3/AHCzpeVFDpYtLSOqMdXxIOiUVhkJwX4lQKIJJC
X/yJ5BQcWox3nwJLUClollHMQ9V9un6xQ6WSs7BAp/aOBeaO2X182OXyjc1Ets/2
VDkgU6vaNaxRTmblfhJ8tVPh7y2z9YhILFqBp7AJz+rPKpvEmRtnMmCHL2jqO/BL
837l+r7drxxupPW4BxHMNkWgGarL67QXZ8lyvVpjlAp07saOfotSO0X/2PXNxztG
6UC+qpgnKtdGBVW2amEtFNiE4IP9bb1glz0/wjZ7wy1Y0eVMAGAY+iwEHfsYKRj3
EA+POqOUnMK4vvx6g+a3/uuc6tcmgeuNt9O+lU6P2uYrgpTJEb0GKT0eQDkSZE7p
+TMTg8ZRt6i9KGCAirqxqSXWA8JwYQI94zwPoLRFBsnGfPRCNuROyGdehKhBL9pb
1Mi5LGAsBbKFociIAonc0Cqe6ZIC59sDrNAzEAir3mvm4JnLanrow0NyA116R/W3
RAsdpqrvyQSIZDTxC8X72AEnEr333CsYzWFrJ849XDwmG6/4WrAzJoGF16p/78wG
QT/KivBbXGqWbFl3Yq66P46/Cdj9/bzDxMxq5W07dGG3UYbxUWyohS/SkO/K4RVC
4ey2c2CkBwUw9pZbJAA8ddfHybE9ayOTkEa4ws9QQZctpra5V9nyzSwusf61E7aF
sHFcphUO4JDf5jgyeK0RdJgdaLseRAwMbxWpnzr+lc3kdMnIi14jERZA+/yBeYCN
XWIsLv79KzNbFOyLtBdyMRtCLLsXXuxxDSJyltafCz6T/gB7bELNf1vTheJmY9EY
Qa0NuhpyIOW2FzvJhER7h3MIM4STnheHU9VaMURXSjmKO00XECix5lcKVZcxmyzC
Xv+ly3DOX5pQ1Vgxv+uDQkpB1fKbiG79uIo3e8wf2k3BkSm14yjyTCcc0ElXfaWm
SuCTH2YkiUXv4B7ZLKcMUg31380VXY1Kh+DcJWaMZmfwe1ZOpKM2XpMgsSWWaO8d
A1pDco4YwSw2V/bfa9+rTwBKXPJ40lOz8zfHgOrE2VQnK/bbYsZN4tAzvvoBZf+W
trIUTaCWdDJY4YJ+r0sqVLgZk920JCEx6n69p7Eg8URPJ71TJSM6AVQfNutbEN9q
ty6LYQ3vTEZRp5N/9vG4m5xgmX5zH3e9q110HW4JdP/aFugKnb9ZgVNqUAVs8W7M
fLkKwLQlz8IlhjveX3+Z5/vwU2MmoTCb+QP2h0ANG45QxH+S9vgD0WnAw+nv2rml
x7204jZgNFl2voGN7iGeLPPe31h/c6jKjgczfpqHvVNXiDwmX7XrCy57lwWIj3ss
m4tn3lzDCyliDZcQJOVLY26B/U4v8A9kiETyIXGg4jxyf7PYGs17tY5mB9GjBbAS
bgfSS8RfawgeKB4cat95Rgsl7sXYT2JXK7H287MsTfPquUI09VBqKpwh4L13BI7f
E6JlaJ/OrHzrfQwxNq+NzEU+3LeBtitP+nRH0bFn78Lh3z8W4r7GgteeIHgP3XVM
scVGNGbon9qn1HOM6ZSJVbwL9VVEqaqAIgL8zdJfTMvy0xp3dwbzaeY5sTFx0sxs
R5HOsEPRjWVpn+tKUSGD8i/x675/Ep6HO6Mm0v7wrU7PEKFP1ODbx94cCc8nQ5TI
U1Bx1ieQFrgZFl91r89WzjxKFn/Ctqp3OkY+hZOMbPOb+BNuNB1nWHpleogCEGO2
sUe2ajOkGTkAGod6JXnVJ5x8f8Tsm558NW1CmBhyHCaS3dmCNkJfGhCih9d62ZJV
CoY9LhMx3H5n6dsrtTTACkD+5f5UcVOOfwDeZc+XKY4vEEyuSPscCYGyRSWPPREn
amFZEc4jrOF+MF4y4al6xzJobUWRqe9isXodHkdzQmudVI8yN7J8eV+LhNorVF6b
8rAeXP7JGNAumHaq9TLCtmzhjuRxIJCAawIIxmPfEnySupoq3oouBETNAzjl0Txt
RJRht/FyLLMhqLb7pxy9lcrT9k1iMkXOPSb6Sjsjgzkvd3di88NFhmRWrxfivgJE
Ekt6xq8UpdeZEex3bk5U8dBaOr8+tBOMxYyH04yQgm2iT667Bi/jaNhIVLdeUzEY
X7IV47QObUZYyqgYL7KrLSgsSHFW+/DuT08OFu9ciHJt/S7Xl8gxfcTJlAbgnpxF
MB/vdXUchfmmNh1vO6466e78mBi2u+Za6obDDkG7xrD7nMduxtDYYRen4xZnzmV3
4RMur93zz4zSXM2q1DoYnTrWkYNaIXCMy863jYdqW3MeIjaugNraagp/nqiRJBI7
czq0nVFyWPBGz/J+uo4Vuj6qHZVn9YXVdlm7yxtZvolm66srlMdZ4CdhFG/g/9h1
ctUhImDkmprtYKdcyXyYihpfgjtbeZtr9KN+sIcKFqBqPdUepRzRuk26yuqZJzX4
eJ2vu8F4IXNb1N4uUyeEd9dEHmd7As9LeqaAfLhWK2IpHB3r5pz9vLiqq7kZHlPt
P2fE1273hd9wM/LDn7ybesm1WmlntbIEYUcWjUY1Ru6LqJko5t2AhNJJXYUO+a8C
2+IR3cznvJjAHSukwPDchzs9UCm7rF1iu0XKfhjj/O0N70tkxyrYeki5VB+LUE+i
5Sf3fGTb9UKCiXVpxLNEHO8L1yqzs5QMkpzUwsWeIxAUDf5ZjnvgcPpwkqx+sd9j
jq08NVCoGO6SSk8JB+Y1m20s88c9vkzOUvp6efK5Xz9O62sijX/GEay3YomFzpa3
8PKZ3Xw5LjBrqOiXSP1jPmf7MfyVK9D8sGXWLT4yRcPJg2LgpuQyH0gwFPClBGxn
OSMinTJ6oOmMR7dEWRj4C8QYU5p32Rd2pA2eBDBW/gq3RmicCoJ1m0hasvOupkHu
FdsJE6DIwBd0LjepPALACDWcTUdwH9klTWXzEZSBqspWmF53yv9xV9mO/HGkZyNh
dXgb2qkJ9c8gpRhu/WU/qA==
`protect end_protected