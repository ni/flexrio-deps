`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36768 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
EQKoDAcJ/8QYHXxJAKTmMGsAEUNjlla4HvfOonvoLfIIl4LuruOoe3Tcx/8SZDE3
aKvWK7EbMTKkA5r/rE2KC2Wz/B1WK4Toe/a5DzDi6EhBtAz8O+2BMo33lY7Ie+F/
FtWM1iedczOLOiMTU7r7DqH3idnh4J3HL78c0Z+/23XboUOftSkbhUQeCDzcQsti
UaerGaruYJ3vivRHbmX45PM2tWH/UFs+VvHot0dIJ74njca2KFEUWeKIMPs6DfHo
tOjIxSIli4NOq8KR6dBClR5S48uYZdvRXj0RVsNcsRCOWS9hXHM13sd89TiZ5pra
I7yDebXykIVmlP2qlYzG+ArpO+iwGDVxsseewS1jL1Mi3AJGBF6VOKa8r/dSyxvJ
XHl4bqNz/Nd8fmxshHDp1e6fMRDP21JXkFPWAGCfs9SLQxFgNfF28xBPPIdSyPXt
S/50IR6/feBczo9oJlJ2YY4bB6yxaFMhaVZR9awVivEikn1bZfA+4yDUX/sLk5Oi
y+4amjuEP4GPTsIGBCyPqNvGMhTAhOcCP6a6XT2COdzugD+ExIlXTdv/d1/Da4B5
o2MEPOMxxWHlX2oPhSd6/1p4V/Xxvo8H8KfES6BXxC6gwHYz/DX0apOgG+NKYA07
DGFcItzVLBWL5CUb9tgyid/hQwtsbkK4kdH8IO5U9ExGooFK7Txv+QWODZMWwRB/
dZjrsMEA7kAh72mKgZOCkc/wig7K7nD/iC2BNcFCG8YIX754eGKPiZFRRtwgQqn1
HVjWSsOW3J4w7IR1MZYWnoswvhAQeAH9V+qxHqTeiTXrd5D5HzRyw9+1WNTNWQB+
FBpaOpuIV9q1zj+UDDvtDOPEusId8v9WGr21D3YLJUzZJzMPGZe4ql8B3BW0+Eqf
1yNVZiPrVD8mtHIRgphtx+rsM9+VGOAceCMd+AZnAs/cjKvmAPq/05P/aJbPVT+/
YL3QB/+yPdGdiaLOeILa6CdSViUb6y+zomp0bbh7RdMP3JRVLfseuzOKGPFM1WiZ
SUWCmyh6vgzQWOkuiNd849XZ1sH3nKW0yrMdxaa74OhVqIXS7VykC0FfGyvqP0Ak
DlVtkBlLyBtuNfHrF5f1mcxtGWRT7bm6m9VoqPmJi/uI6sH4j9LoGYiIvNTREou1
1R5gI8geHvudGyhXsuSReI/RE74o7TPIt1jwIkv1Mu6sKyFgsLUD5NXXyr5dBOeX
qOON6+jdaPHzdCzU9BoZjByN1yOp7KHjv8tDhai3gXGKK3NU7I02Yn9fxyWPbiFz
dB+YYtCxB7jfyGr86ITPtHmDOnMPfPOmCwF9kKubkiObI0WhN0D4mJTKEpR/44Ty
JhWY+9aRBqcIJJoDjFygcwItxpdKDLiTwl/U/grO02pzcEGU1lAuPVmwQQbeMB20
I9eGP2iwkVomGPjRhwqaCGYahe0m6cT9pI/GAiJN8wmQSsuuETcoBU+K20AIrdXe
7DSCIEdRq8FmXxH5GT2OkhIBFMfDhWoZEidxh6dKiADlPRxSSFVdq2auQ16lwft9
fyuC8GfANc67C2iTuaF7bP7v+har23POnCYKlRs5siUP10+JlWBjrSDCJ59QeQEB
0pxyy95aDhtdV1gDn8qgC2UCIFRgHxYL6CFbQ3LdzH78BaYTJeSxrxIiSViO/M/r
JtbF9VYDAFOIzzuvWxkcHH3X8/3mXkIDTTGvH4asu8z5L/WMD+d7teR6t3jrX3e4
/F4vNxGFJqr7uS+r8KWwK9Tb68okXYaDBhKrFAT9Pi+exI+4uQmZjc7Y42r85OuB
o9UUq9ppke2TkgISqFzydUFUZk5+zTfYO3+m+WXMd1rgNFbzoM5U+uckfidE520f
ksLTOd9LIcMYxVtC9Y764GndpcDFUb05fSKH+zOTJ0Ib7TgQp+Bp1f2DitT8smxc
kU3BYeTlIF0PPdBXn64WTSNv+ce8aDihd2GiNVGE+SIEbPlnpg0x5Fnxc0RoaZxt
K1Pp0Adi06V4vMrZMzF90fGlpsruq3XGEx6uyz6B8RJdg8L9n2Q5beSZRpffBA8G
kZDoDze0aTDefqRpGlbZV2pDXNdHtv25MnZOtanC5rK1IUrussn/DJRc+uziCLGs
Kq7Ix1ItpFu8CNKXrBAt9TWk3M7TF8hfc+hGldEVhCF9/dyQIIo3ofPXgvdT101V
ATO+V11XWeFSv9j5SgfeVfuRoFOjhV7Kgs2paMoF2wOTSZnI7MCW1gmVSGafX2Of
hWWi70gKlensr9HYOqupj8QfYQLqIQUvFlmhqZ+uixO3iqWL87KvLwe2uJUdQIRC
1O3zmboyOUTTTM6ayC/YUyDukVNCh2Z9UlkZMIafYPcQkVm13AGT/PPxWSeoIQ/y
O+nNNkfDZoQJMJlh+cRij9w95NGle9S7VVjRIVNpVTtxVyK4/4A+mGaSbj4eT0/h
rCIsn8db3+pc8ShsH5yuhYX33WhyN5M3hizohD/5D3nZD4uLBORXsKU3ZI21TEDG
PcZ8s25mcDj6WRT085exXshXIpEij32aenCJe++puq/oTDlErOAG3H0azOM0ptq6
H3Aav+f+S5+6h1efOdkDrEC6A/pfyb8b2Tkn9gq4l8DNQOix0RDYoxPhlHH0SomU
Tad31KWs5ofx0Bnvxo+YC8UokaC2uk4dnD2h+BKMMggqGndZ1kOu7JsYYrZu/K1V
ou6BgAZwERPjUoB7KTm/BzbLCNd+9qVWAahDHz15h0F7scKvbEkA/B0fKyVRmMZ9
xnsyBGEEmHRa3jsDjCdLuXEGT2hpP93PWtmEh2v82iYRIhTQKISo3kPZhZwOur2d
EMZRd447BU5xxnlZ/iasqEMppojv3gYdQdpZ1U+IlkB3y31X8vsl/FgXtnyoR4fB
gkSCA+oIaDosj2U/hVpEss6Hxc6mWbxiZGfuRJYcVhnVodwUHrITtTj7AmLB+fXj
uqpT9V0aHVnFEKnOL9rgfood+Mh1N9wQckT/l97hII44Wl/dgcY09xIvN9gLctl7
hbW/xEV+CT94T49hCx0RLXAX2vRVKuTTlp/Wj5eM+FdaWKvigsbP14MRvWnvHwUZ
8wvIR6CMO89NvxCj9nxQHCJc/2aHxltnOUwLPvYXHOAlRB7z/8W7enTrRkFg6nQs
SSHZXEQPqeu3au8WSC35atEege03MnaiwLw1mfaEhYtPsYrpQxIxNCyDD2xr85C9
ioaYqIc+7CHWD+mbAiUteFd9ZUBMP1k6ITLf6MiS4G6OylaO2yufVb8sitFg2CgZ
9ZuARDW4XkP3djnPqRRVCnC7FO/VVmHpJ92OCadGh6xzh0s2BkhBpFIQ7+ucI4/8
b354dxqX7d4yR/MRvMz5F9cVSQhnQduJDKu9w40IkP8f4XZmEibi0HsvYy+TDr9f
Pnon1FeM3DigWjDaryrGdQBhg24HrRvP8vzTMal9pk/6dIy8IJSIoeFg7Mxp8EfL
HjB2/5bO/DMg/S+xOPEiW3Qy9r8YaNqJnKABkkynbp0lFuQaP/Bze4T2tr46lCpg
6ezhIHHRpjCy6rPhkHw8aG50rqMK7XYJ1XGzU0LjosRoaHMDE7A5U9AGgdB8DwmZ
oKYxIV9EyJqYEv80syAktTfsAkw/xjZ7bpo3C6Nwx2dA9TV5Y/kk9nT6nOQzsdFQ
DhABlxUyAYprq0xCs/guxDvpyt8O1yjsqlp6HzBluG4rWL1qvavkAyxh58/1YT1r
ZF17nqeskJiVG87i8LwEicdA1Jk4gA2sMzQ22etUglRgbkCb/LsK8TA52BnZ2OiK
jDLZVo5/gJHBNzDN8HlCC1H8e9uepzfX36GR6xQDJX/bsUFhuc1NsAMze1HKMnBh
jrEECcA1l4KKMc47VTvtE4DzqEQ6R0XAarFKfyHzQdAgFTlXT7AtpY7H+LRK+veN
Bz5Sx4mf95XVcB4K3y8xWm5K+XHIFERX2RXiyRzQ8+iQzfPAjGp5tCaRjdhCq5tx
u2/wjrJOIY3xZOLOpMvd+NIFMGUbx82MIq2PGr74svH2ACCcB7nerkrAMiVnsael
U8a1fmdVfUHxHKbdR/folJ3K57GMrptSGm6UD7uZbjGQXiV5+Q9YrGVOCsDxgQQ5
mg97zJLOyIUHhI4E03QldK9U40/433mBs6WeWgcc8RFyFgoJtraYVSea/0JyBeBg
7+GhlXX66fNLb7soSg8XcikKZXpHDwJtkU3Yk7B/E74lbVvJlRUhNsDkTLgdsgUH
DJyjblK4SdLPqjJVkf+z5r9e+66UoeHXp8FitgJiTmx2Zab+RwAYewK0hDBq7eEd
0fcWqtx6LjFfp/hMfrisNEAqerW8N1VB18bgwaQAQi9TYLpe+Q1I5YwXOm5GCj3H
hJ1TLnR5Ovef9HOC4QGycmRG45DEx1jOUzHdZ37SvseVjR2yVJ0+15R5yvsbgmPl
iM939/vN4IzU+CYPWa/OBmRJt3UMVxpp3v0LL2cDjmKY6ZBTyp7rWfHjPyBFfDKV
QZFVnjeNpYUeBBgI3y32nhbcfsVuAXuioqaSj3ES2/9obT6YN//pR7wtCN0Dkozx
BGfoxhYE5jb/WXos24v1vzG3srIMwmWeI25igu4PWIBXJUS2iJJNbOqeHPWgQOSu
bnbBAGwW2G9vzNhgbrJPLt0yhKIR1/F7q74CBio9782ZZXM8vUocDoPTH+Zx/XzO
A3Q+6W3qlQI+Ec1WZkYn4KhQLz9eYhD/IORsshQpTj02feaHmEV4RGJJLCgD/L3n
6AoAMzPbZmsca1rc0Ii0vdRc1yDeqM8Pfkq2wI5xV4b2eulbvKvTy2Ke3fpK5t+L
NL11DMArqSZ6akndeXggij+zU7FRx6Omd39gDSm+zOVMYIn7VVK+VtbL+GlQfAwS
KmhwL6sTN1k2aUK5TV91uQ2YDN6cIPN4A7xlfhxlT1ayIK+FK+AL5/OnGv3rDE2B
uFWKWtlB0kLdU78phqiuurxboFGrtmzaRmwes9TFDQBo5GWDbwdPtQ9Tgu4GuiAV
5qlUyQCUBqje20pFQSx1LQiX9vbaShjY9btAcVpPJU5bSOXT7ij6NEZ7euSMv31L
q0CEBUaoTRZ47c9s6MbtLSKqH8jvD7WPv1EJ56TXubdU0ATvtC5YgN2998RAMEV3
ZxJb4OJcw0vJGrbiZ0jeEJicvnqPcxvtxPYrPTxY4Grbv0mU9Tu6/z1/VQbP2GmO
/RfIeKxlB9orLCGp6z1OgNS2q3sVs5jj3CpgF8spocHAmPB8BLKd7UFvZjASgS98
zP4SBRsCwhw6/D5iEpP6KAWxpUflUYHhpCuiHhuQK7YF2TTXCq7C6KBEi60cpzJK
okYlqZe8jO7oRDo0h3C3VyFP/skWC5yW5wskT2tJJh3O+GkoEyyDi/9SOcdM6I/g
p+WvwiTGd2Wl5i+KaiIdJN0LxyCaMsPSEyJWclfBdFOddOARwGhGJDgLwgGaQbJ/
E3BOml5jJ+WL/Mxfdkch+4paclxceTpTP1TJBkRFARPnPYoc67EX4NC/JTfR6zTO
XL0fHDic2p66iLKfSixgELbikW0RfmN2L1eweyzi6aFaTFAfyVmMqpUKrj/IQHZ7
MJ79C1gl4/nb8jsGxOkKxNb/RXdp3XUFDrSHdlH5IZ7BvLwIJkOccNSTFXyTRR32
fMVaa0B7Yt0HYUz0CXBeHo0FJq6BX+LYTeXlDVXRVzTkMFCMckZiE+zKVCCE29yc
BZmv4Q4i6DcK4sXi+oyfZRQ81SnFSvcDWoCI8gopcLlLvUJ3uRfe5jqwy20NDx01
23YbvI41Hz1E+H3tClis2SgZrSWY9AlZLjWzU9DxpW+Mx443YwIHiN+r9D9z2kCl
x9anfxl7MiKPfalQMXobJep6fzx5AiVci4/qLOSooJEuT9j2aaTOwLcvygDo0ARD
KgS4aIb623Uzmka7Bxh+OqX2+6n0r7hfwuM1mwwBlWH7JmCR6DWNsaQcx/sQu3xw
m0tvp2EbTG7Eq7ia5ZE7azh5wnRxn7JxwJZQHO88g0nurLhKr+QvP14I38msY3hn
a4JSbLq8Xc+ZHot6nityJv6WSnJzVM6ROctUn3fvXJc3m5Ka0tX1WgeBI48KeJFf
OHkIbNwwoiSxEGNtymtk5SHydW0yYwj6ge/3MJ2yyCv3AVGQIJHw1inoMja1MqYw
TBYA9vyKfXkcBKp/M1AnH8E1UV4JgmS97g1U8Gjnk3zqVnHpQ4hIBckAAbvsQbke
wK0d+6MzY3g/6bcSXMWZvWbh5AeXDXdLjme8oE+u2YKpLGNilBhoNP7PFlkAcpMe
67XlG2OP36KsJPmylJvzGt8lZDIbx2ix+3Nf9jFo/f6ZtPzm1Ik5kaa8BjH6VSa+
Bus9JVR64hXNxqbPOncmfzGl0+ViTW2LJ4ShvgwBEIb+mwmCiXPguNORyjTi13CN
kbd8jfNILp7kw6dDaQc64EZuGt2Z9LdM2qLP2qkKnwqN/UbHjbmREl97Rz7UhEH1
aDmU0t+aXcfFrwpwSDH+YrLbQhe45qTLVmwB8tEVHDcvopbeuoFL2wctFgw2jHsL
o87wMm4an+6QP4OZaGEaj2Fh5ubHmJ15aSCww62SAn7gPTjKEEeiUSactrkkwdZ0
Dz81MGszPyipCnzow9n+AXYHKRvqYhdZecEAY9xkeym6jVuuvniY2eqcaj4Heu7x
rw5V69QE/7exm7EU3b4LJg5JOIaZSPavQLR1+zaoE427Mx0UwuU7wNCw8YGsSsmy
biH3WBi+BJ5j6vwM0N7Afat3rjXWGvomghtkz6q61Ao2w5WWkr6zluOBSyyCSWCp
flEm+IXQKEBUcndHFYAVGdL+YvSH+GAEJLTWDNb6juM4ZIhRohzWZlc1/mABK8B/
4yQTGbAM5VuqCksdrCAWF6C2m8Epm+mBeHmEEBLltFGiGAVJH6aQY61LPkxyDSy/
7R+PFCdSaYWDyUZBMJon6Yp2JDc3JKYx96mcV2MDYvm1BUmh7VA3b0Qc86iJQk6/
0OB1fCcYTVL+fVgQHGFKMNu1WGWdc50bpgzQ6uKcM0eN3B+lGfMDb1bhxbAYRCAm
U62uFokFxnreWeZCCjrpU8jYhBgiYsBgdxJjJX+jJH5EAFwJvy+Fa5m9nrmKyFE5
QHojwxQJSfRYfULYiTsWvuPAmxlD/tHazLg9XyC2hkD5h24MwHmaaFFkbWr08p/P
BpN+17s3qTiYSXomg/s1a2ozm95EeUi3oHpBaH8ME1ZY2QkEBVL0W1JoE2qoOh8q
T4w2yI9T6/u+i2KPrp9GE7boeYY/Osdgtk0n3n+NdezeC8cmkJDsf2gPTpel2Oo5
UDDwMTjmp00qKnVuqClQvuKKGkk1uNt24HukYLLNkkxxhpchUfGPbYnuzfuT7593
OR71z5iNaTjnuJW8e6O7/Y1XFgzp/UGkbFlWkqJf9ZEvK2QwVXlcn/YAuaBUkRnz
Ur1tqvlQbykX6HKy/6jTAC3cp7IB1l7pZ6isE/grjjUpsOsZZaXbqwgte/5zD+kH
EVeuJ/oiBJYxiGSgmfDUCAztFbULkvBB6WiBNHr/nexuVcCKFZeOoI3Kd8w5Fe89
BywQjkR8s0vuOlD8EC2oue2qck/YAoPzIJaUl9lpvujYJ5nuW8qdpmuX6EZkOU5h
xoFCLdW8hoRAwqb76BezGJfcoHsJ8PeFNt0n6Dj93NiJ/8GoqcJgh/i4Eh4etVnf
dqWFa0Yiy9XFLEugqyJNjRCYqy2quG5S4Yb80u/4LiWIRp3xWCKE8XbgDfnclMQH
tGhnlCjQrueP9h2X9JZInG+mEdWlD71vQsz9U7WPxMfwdjkH7q22L8XZH+6EU1UO
4HhFu2mLmn0iT96zNUqE9A6FSoRvo2q929Jucu9JuybRhwG7ZnAjBr4GIsovan5Z
nbgkKzg8fqKiXUsBjfZ4f975ZOZ/NI+K8+EHfBp60JtvGkkkXhaqUb6Az5E1w4rN
HKKV4+iRbFYfCmDNiGoFwpqboqu7dmJIZkC1250GcLQbzKEiSlmKSEzJ3RghXHk4
l4DdXUXBILymL/RSdBoIGFC7M0jhF0dOdx2Tga8bZpYpg1hIeCfahwmutXTu6QH3
nU54Tc/DgRRG+LCXSRPiNXUv15Nzl/cMXVDc8T0/Awv+CCIQDoV38ZDH3jgf076E
ohx243ts9+upBf+GEOq59XE8EbnYaP+ZgRN5VM7wag7kNtooA/LD9oMhr1Gqqfri
1+fwIAIrCxCIcZGwkJU0463/uVcZZ7Qua6vLsVtiLtV6ILa9/gH+vGyxeyLTtYGH
1YY46kXZQfU57Jkb5HoQVl+35xirJ61cD9AASahkAkIhpQov7c0ypbuOJwSOWxoa
p6qoGd9w/lHRyd2Xwq1suHAQ40Ve0tXYmAa6aIgM4VYAUOVGfzcJwQi41WF/xwP6
OEPkLQNQoHNJp5HvlDhrIhHX7Pm6m4mvYPlVGkCMj9MpWumN2v8yovYmkSh8jLbe
Crex3C/v2RIkb0LDDjX+iTh3NTigfs/2n/OwGs7Nhs3BPuiYGOhEtWYXyMIwTwVi
DTF5+UvdVGPsW/J36kMvU+x6pYNaE8+Zj7+HOznIIAYfgUDpRH2yvLMJktXgpeOo
hqtS6sKhpJkzCa6/H1bB80PIRGOLo3V0+ttdmEUPrpW/mpJjyhCW0Xlta7BZhueh
xkD0rqxmMwg2Sq77ViMRYueKimy3UKiMcp8RaEJUbwyc01vn5xmC5GAyhE1Qqvek
d7ROqZjOX6yH4QeFakWTwVRZ3Nh0/2nXzvLjIaBYlWqki5dAh0zo8Eb05UJ/qAQp
79IIaPyinJDy3wRsCsoAJ+hc0IDzTva0RRlfXFekUk2UeSDlxyTTJK8UycMq4poU
j4cz5hYQH3JgwAJDFiTwxjk2jeo+i6MsJlp44lGRI/NKApmssRG6lA0ApxD8eyTt
g2u9Vf9I4U1OH1VKjfLRvx2j0qB6aCzI6B6OZnBDbohXr9vd4HPn9vP4EaYK90dP
408lBBP8VN0mocSzVGNBv2Npg4rcjN09fS0jDUvSSY1Ks67HYO/wp+ZLBQtIWD6E
Q1aPNlhV38TXS92quxdLcF1ewUYgu/UpwN57RLmSGwdE40H5hbuOe/TzkrBI+zxv
fLJwOVHu3V6U4ZAq8tLLFbio1TngngzAhbW0mEmaDcugfwQjRw6wHeUZqhhu+VW7
eFaBxsDZVdmZHJUd96rAcFzDezsqFHESGzfN0PDts36P9CMo8z6RiRN3181M/b0M
xAb7btCvVLv7twkL1DWzobshmvVNCLZrZjdKqPqCQWa+FN7buX64z9FJURgzzzwr
3Ql237/iWHowDnDeeBUxe0HRqZBf9MDiDD+2K3Q8kJ3mg2wkE9ITAS99wYUcsmFZ
ObeUstNuwXLS5vTdPjQVXBbKlow5j4JPKgV3Orck2aTZfdzeqaaOhkCNXi9FtnlY
1I3LLBtjVOIN0rm0MOwHa9RWyR+b7VGOhcdu486N9kT4knOCt2sWZi8vpnWKN0wl
G21mWlHRSsz94Wd1QmiQ4nSyCEuRpm08VXvkt0IyQ7VM2NfcOFsL/TSGvHTyyfJX
B0iFTBozCu6g7eofCtzEhOEFoZpsyblKPWCukT4lCuAIzDZYT33/eO9pFKh3kGZk
dP3Rns2E+DUMA/E7T3KIrwOD1UFGs2fNfpQJnIOeBRVDpmGaHe2heQURTLquKNsY
3Ey7St1BM9LrU0h3OYTR8BX5EnCQfwQic9bi+mU5CnvV51cOdWR28LP7/v+tLLzk
yTgmLzqc68tIU7Yd03fbBBesyS0+jqOAtVNV21h+fMstvQDzPqv8jZ7KKbNRKtMX
Cu2s2VDpXN15L7wfQRotpupKSToaJUiEAIg0imNSsNSq3ZWZ8YA2/BcR6nSeMH6V
a8RB9EVFp0L+qQIwWPv9X6XIQllzTcUUy9kbRZX3JLl8KzKDdtFuisns2TlVd+S7
1q7Qy3BJH/Detw5QBdUuRMYtYCAX7VAHNllvsubqYuAdSv0R63EztMMu4VtxpQzP
gT0+V36tE04ZpjQCUE7ZE5AFoOqF/g/alAx2gZY1E9Bgn/hOXk3589h2tbBmygWE
mWqi5Rh4GFRQpiWgxAdEoZJkuZQFVW/4goEg6TyEuagjmQlDfAfGT098h7IQF2UV
lstQGwBgA6Cu5R53oDz1bElv9RNhezFOZS9iQlGlfEAZHxQ/X8gkaOdYJvPCiVgt
njFipFuNGIXzL4M8xqF+TDxId/5X3IzL01QMoGN7+qEJzGzQyucrfSM9vlFvm8ZV
RDldGDYEmBYToVP0l9C/syDg6ZCFqE416513xjsnXA3KcmtL22BwzhEHE9fooQY/
NF8Cegla+1iQkQv5VQ7s4nzfh4H60epyrCRpHGMf1J1i4X72fPOl8lNkE6i18YD2
k3llZ9dl4dcdJxZjih0wL9Ra1jrf5qq+3sbpfAIeQBcFMsj8X/oUWUuJ+IaAP6lu
9GiNrTVarPsB1BAsdtHlNe4tOYB7qpL/8UHgvmKM8+4Keo24BwT+fHbfEQUlHTZV
GXy4nVhT8Y4ruC1EI7QG9/ozjptTYz7b1OdNvrL5ZFuqltp+czkTclMhO3xNlf7A
Os+hVU3FnCok28cKB4tQVuW6cJXcFpbIDhZFCWe8aUG3+IdiI/vCqJhAAtFcjXZ0
etoIVg1LuLQeAzRNjfnV05bT0779GO9GtHWT0YPbezeQOq+SKC4bC6DWaBE519j8
TY/gihtYqVIIJwe2eU+5TicJuhy0qy2oMzViNKgGYQ3pYr/dJbvcZt1Sfm/ysuCZ
BBkBE/waIaA97gY0wi7qC/mgoF2vcizTwTYop5hKtk8qPIKHX3l1KmOPPYpkSLC1
u1nP6Q22rrqSxfZB84RZSfZHje8b5Dv7CZZKDBmobxEflwuVcdN7WJJpS3RHYEVq
dcII7UrMOJ9ooiNzH7/H0YRlgvsRUf+YOPMrQubMz2o7zBfhnFZpvgfMLKCFmXCg
u8+KTcS1FitNvno2i9/UOkjN15CCQpI7t3isZtbrfeJtHRS52jRD3ONDDoe2cUlt
rAXxoDRhASZubWf1NVBI+KKnCXo4CNI4so/8mIxLejIv+HJVnRmdvIG4IE8Ux//J
GFS7uEMKE6ehAtAY4zmpeYUU7yEKJbMHgxIeI+7+y28H28OxKhSoZO/lkLxFf9fJ
7bmhB2LLT2rPAgMH+AwJL5LQHnd/0hJL1+qkYSZa8xMs3Mtpe7nONzJqNZS3WhrH
0X4mMOuNzOuhFpS5zepkwU0nO91ej2YmtEHrDKn93awVu2bUdizjzbunHYKeJiYY
vCcQNX+nFBgyHsD/xDECdQPqGOaSXi7FGFOuOVkQj6SYf1t0PFJK5ebqGcTv/OQs
rtqmwpv2Bv1UXYI82Xavq1UVka0En9K5j7Xjv2bWrb3tTcAEnAcTFa/905eWvGCo
MiXLR3qT9BN8HkpS0TJxRFqHDHFudk0FcmW1bmVmLgaFoGI7OlLihwZRikTQJrFg
iKqNWzI6RmvGz05DGBVMiRh8IG5EiHC8M2yXRlcEsheXcNaJJkTbjohK523RWxeV
0NSVBh8VxG0jLNvapUGqaD3/zt3+y9bYZSwF8MJFxMrRxVrHtmh3Ia9PVktyRfyc
cHYPXNa3WrekT6C9W8G22x2u+lO/UldLrV6kNlYCBf+V/661bbA+GURZ3BfSp4Iu
aRI6gTJ5MwWJS0W/eoBtmRatpN/kOtaicHmx70YKYCoDLGXT2J72B4nstUDDLkES
bmwX77VoEm5fbF8VIO4YpE2+qhu9uMRXsBu9wSuqK0AHZFGDN6vBzQrrygS19gYh
yYWpi5xJyDE5XNDpwiksfBiVKgAbDyaGnxZkq0IJ4iaoAQuHDHgKL0lC+cBWOvnY
xgAPI5d/kbxziPJifu17iPb6uHDPJJH9VhWG99U3eQeJ/pE3NxG5fTG2z0uSiLB6
oe4kXpxLkCIVAfRrJCHZvWHSRrqtP3HmzrBK0PoVhmqMXPlQfyiGJHCq4tMjRhO2
FkAmOTSCslTxP5GOsHvP28+nkMrM+Je22JQy/CDmhYfz2+wCzZDzE9V+41TxLVWy
Q2VY3RikArSmWSm1B1CmrIl+QxR1JoAvORZRygViQTn53UpCTLS7OCtgFnPDN47Q
I+8Y3EuvC4vk5kk4LanrGoZAYtjy3ISlxD1IRlXzlu6WFfgiyL52+DjVddySejEy
mMMU0ky0bS5P3p5/QiWhaebGKLCgQTaQX9jqw1jDueIqtBraTzU1tJZTpYtOwOEv
RGyJzcA9/6fuUNaXzr+XLHGHh2VaxZ7b2tvYgXFd8hVU22/VaBet8FWUzLN6GSFY
rq/VrCL4a8QjO7V0Q45SqHRyFqYXSkDpkHyMIROgYznQ5jq3CkBZzdg9Fd36o4ZF
eidGmOQkdZ4IVeD/cbY5euDxXO42QB2s8mkHMTB1xTWbv1zxprTk3q2h1rnI1cdl
XndlW9qHa/ionxJSnxU4w2/zFzs9n4qTSKz48h/aPrvFv+MqaS4a3NHHkLdUEQ6z
pwLg6SZ6N+8ObAAH3Z00aCmDAHaPqpPQ9mCdLB88BPm8SXb2NSLSgurQrNWwuYj6
8cxtv2nzDYg+2ly4xsr8soob7qrHHc9bpoy/dD02Dv4TqPQ66n2sjp4v85eSIJkz
GQfoXhJBbIi+S8RGmVTlZA0t+dJnWabMivLt2czi+1n7h/mniClwjnba1qEH8/ZI
B85lc4mcvs84EkbZ2/J1MCdqO8LdNuLmbtt5Ngvc8irVVvLIBkatkaf1nhomUx1z
rM4mX4nERxUjb9IpW+09O9+iSeEodjfYz7bP25l7sR6uB41lTe8Y8CFLYJkDfJXF
vkS0g4vDjkXtLVZk7yUEf7TlINYDdMxstAa+3vGxVZJeinmXXTUjrkej495vfPra
+K+/5/x+Lw95r6ghtHWRTvwZrFCLjX5W1cH9yz1lBaUIR9zi7xCTmlBcnlsgenpU
eI26uOnzHj97LdAgxcL2kKLLXuwP9uGc+0hpN12LK8XpQHlLQF6kf+fY7yPv83CK
2kUP+dj+c8DRejOLrOW7Sja2m5coSw+qgFGsMailxPGX8NuP/B95yBLbmsPKcUyI
VeRdujXgq4DFVBKyttrQ+dzouvNFCZTFaCTk7Eap72Fqx1Iv+9JPug8iCjn1PBuJ
7Ag3tP8pCDosaw6EDymkkeHBQeXzjooFmd2Q/UlJi0lCc0ky9zJ7eUqG03sXx1c7
ruF3JyyDR0hxr1A2gDBdUNyQvtRESuDN3zX7uNaHS9VnwQ20MuNTEbItgj4An1+H
r47J3rr/ZKpirlRrDWyVFU9Vc+RadnTUGtPx1Wae2JIoJOGHSD9+acwKmLeyXIDT
z7OdJ53iWl/g7p1AxIWFPsu6E5kohQ82vBUnBinkmmd4n54mzI7YO7iFfcDssTxZ
0XJH1rJf+GHbiBVuNMkihRhhjByLmmU64w2rybqSl7/M8h4CIZSIvCvPXERLsBEn
mhMifZusIChnLJ5ByntY5kXuPNHpwYWrSp+JxRC1BCegTahZr7qHIbepKEjoy9IY
NV4UiNgRkjkTE90Q0/gFZcRXDTXBJAZWOZi7UhlSje8f+6VIgIvHH0bNrV2DqgWU
Ed/HSA9xOFH+WG9yss22SOEiQ5mDjgdsdqKRMYXPdECZvZXr23KbhF/q9FeQRzaQ
fLDkWmSkhefqm51AW+2aecaPLe4XNIUqcOw8xrLtBU5ya98OubW9OEi5+0EgqWee
tQsoXET5zYYGV2Sqj5bBb3K+voJovKZJWSxN71g/X8uDpoBI34G1ZwRdVSI2YfSd
jfCNtNFEaOXIxIUFjySRkXE5W8XpQmXv9Ae6v68QZXsJVOaRqEEzmPTy7Rzb4AzT
vST/HU6BqHDjJTP9Lh+WrhzL4V6F0Wc4pcCVrOWEObpJU8pVxb+AzksFnT+/jxkF
kMxdfih5x40yksBGzAniFXhOXgYqR7yo1B7RHNQ0VRTPb6lL7BpWNvaRYq0dLnR4
FERMI1nKOxhW1BZvJwU385QNgqWfUCmw0vYZw6dIXbBrYAeuRw/ZOf1QBAOFqmXf
Cs32wcSrgaJyLvTwZgUeiV2QnthZQ9TeFHiZQjJPSnVuGkmcqG1xnoZ6oAnyHzR7
dYgjb62tY1NPBW3CAsKUEPC1cIuPMWgSBOBEmJqjVrkzmgu2CgYR5+feUW8Pe7ST
/X82oBQ1DclyZ7Ys3dQD50d28m21tZZZagSF9yBIQ++CVyCZhiBo1RvxPKxQIlHf
ap+0xa2KKgizfeBvcu9Jg7zhgG5ifFC1KBmRvYGYqP8DpkDSXXocfnVWIolKWbY2
QtnWKxDQ16pQojGXR9RgDV1z58efrxb53xTD2Pg59pHG7LekaLLadFNZ74K+sYpQ
xNaLnDV7MeRT3twyhGhlEzB8Gqoq608HW39DtDuioNJTzGGD6+35xOPhNMX7EKLC
vIUI2cSvY0DEP1++XyoNMh4W+0EBI3GVho9tNB129hSf16E7Svi/Mp+69pz3+Zkp
rDs+yUoLDWwuXQ0mqkZUGN+cgDbQM6LKyOuJ2mdXS5ymgsqwGVXZsZIalXxTagT6
RsBzunSoTnZ90vd57YwYuyY41QqFVSm9ibWcRJCVIWGaoRIHnLkeoSEHPPWKKh5B
0p/LsCoCnoUajLX5DrjCMYu3PFoibLBOr/GVjyVSUbNVV7nXZsctefGV1gbr8+Zu
mPJIxps8oV4TfpJPY75WnJJlMAwMZjyzrkTi+3O41NSJHBnXFKWuBe2TJuNNItQc
IYbsSSoLt9Dr0yjqcw0ZtcYD5TbFfbn+UXNXpKam2AyiAm8Jk2ai+lD5dJxeu5He
P21Bs4TqWfyobwgT7LEF1bc8j+XxX90aOVJHSlp2v1/lBcHwxF/DVubExvglRb3u
8TuUDA1/Pc4NgyIPd+ykFm9I78gEUavdMBfO0LqzaFh5rUyoh+fOLokXoRpTL6P3
B2kXFrK/ZxISk4tRLqTCkUIZeHZA85MHcfiuUPJDJypopoZmE9ROEONTAbe1Cs5V
Hu9NJpJCz0TouNQSUlNXOVL+cplwYu0QReHEh8xhRMtdXDk2uDkvT2vstuFzdAgs
xXBtvK2P9L/tVX/ONAZf7OcK4ZgOD6YHfoETrS4YMh/sweB1wEcF765xxH2URfnC
hzr4p0gk2Nc3G2FfatonwxqcEULMRqkFk9reqZlH/i+fXzlZadwTWoBDw0HXU5bn
gJ+rC94SjMNoVlUKUDXgv74BWDMbs2dNXjeXCiOIS4VXvPA2oOHonXmpwxyoacx5
7ashhGUkAZJytdQKsUzUWEEX989lWjdAgw9oJetfQyOQRHD43OfhHJr1Dc3FEhFV
oIpr+5+JxVw7e+tBSnAN6s5pUANHLaYJ8HZO9iABQC3Mv4ApFwHroere7ZQhtGFa
Qf0aOX4Z5i2OtRBxQzXkXAKZy29TQR6xiSdbEWMA4ZRX6D/NXOha6KF9BnIdL3pO
jrCaCCLYeMjxBZ39EX3ler1XkOf/VUkeGTsRDn+0TJB2HWyyP+utswC1EcOxaM7a
uQVsKX4ce9ixqHUxv2tZIfqMPLL3wEsHxoWVtJ5HthdULBQeUGLvicGnbDuCDNlf
QKKIkon32JJEJG8Teg7h8VlQoHvKJnhNNcy9ynjtU2EtcNt3GJoci+Mit837O7fm
n2S1g8uKT3c9JEnVMgp7lzs015C+mBG1uZZ695/7J0vTfKb53AnvAUpQJEQEy3zQ
8WpQhDle9uuIwXfNLJDQdJEam2n0UwYnsXhJg92b6T8gpJO/NCxruU+5E7TvG+4f
jxcybmQ7Zaqq+pXtfnz61ARdkRt/wPpFoCqRcjEXmyKXCOryoUOn+W/QNIGTpcWy
O9KKzWRYWj+RrMp2DvUvqzdFIhr/jAwWKe+XqFMAjXyCJT7txXdXljkaZZtknQu+
gsAKdR1Aorg00wTHeaw7NBKyMfyWLlT1w81NsDtZADvF/akA7pVj2GugSLd/nBLc
M5T1YhCL/5L4AYam4+TbZtC+lx0F4WiZEsD1W8f1Logl6C5sXqLkBj8MSUUFQSIw
drH9b8qg/2ysx68kwvz+YVOygifqHwE+cbG1zEZDS/eZiRNxsSbWKkm9ZaWaWGon
UVDFm0UVF2WDhZvHaYKM1hesi+ilzrWwO69y9GCqqki2LvvqA6QCEcpS6nIZo3PD
3WEp17OUwQUYRw/g6bCpCC/pi5Dwt+Nn/aw92tS7+y4tkWoHTyYcWsjLeb2UQvPJ
DYQhwSmdpnOEDNWOyVgC1E2eUD8+UCQ8Z0gdTDeYEzm///+bJCth4g5zlLYla/PF
PdLXQcLLdFPWhTeOMPkJjfFqy1S7WRwFKya8nzeaZc58X6zqQAgqZb/ar98ouisI
GFxdlTUmUt3367xCEtYshWyUhQrJTyjqkoJWoYO5NJ693pkgwolghe2wTQQ33ILE
9Go7r0zATHTraIFNmlxcubvaAzFFtMlX3v4memwYLNmMiHdbInVatduoG8AchLPU
qqeJnZSj668GUDACLzUMt9Ds4DGkeuXMzVL/wbkUqII4lMPkcfTLWX4A8UY7YrXY
ny9Irt1Yjj9GUG+Y08lo4BhjL5oZ8BbiWeC+cA5XziVF0IHQMW7QjAaA4hGCETC8
njsZpU8pNrGDvwOodW3weE4J+xoLptdUco5mqAF0PKtncXm589cH8vZ52AVpx3LP
aFeFCfCKPD1QDa7URj0b/VHwl5JLeEIhvMsEEXM5rfjkkJRP/58xvudBok3kmViX
cZwaW6SnubcQgL9F5RCNh+1UNFewD3La2H3JRJ6gMuKfG/oCKke8ZL5wCCxJaI35
TpU8pFi8wgZCpDmHfJMrtNmPulm9O/a4EXfndiYDiyNMPt87p0vjVcyYIjC9sDet
xKNzeLdL2gwv0fevT62C7MnJ3v+UPdK8AJ+IFpLlJy0C49EEHPgCWvhX3frMjD2z
y3xg/49mxbv7NW4ceYySU6S/LHAakztypcudarY+FWIJYUEKfaozlGpyhgmz1GvH
U5EnEupOXdQQEQsZ+1tRIOu+Otea+Bj5mmUwgq0ZYcVNadqLx+dHWzKmKUnp1Uk6
iMoD2C7/BSCsIsUToeyu6SxqCGy9+ZNE+yW3AyFp1y+81y2H9iodSgpxw23ETa6O
U4Uesw3sCSBVC0dnqo+Y9bU9OwytmmZPZwSxHxwTYnm9p9h0oNvHFwQglDWD7YLa
YGSMqPzrtWgPi+/dcEFpIV7hOx3ScYrd3ct40T1oA03Vg6AzDwAmNwzQKNQsvfi3
61KxJC2ZWhoJF8Epf26RyFUmobmJW1G0qT+WsmgEc6bw2IE2AjaVS26BLZx4UFT+
nKQNRxH+0BLUtLKm/gfkWJgnej21o5mztcV+zobQ9YtrSpXOorL6s55gVnSt4nc0
rZCtwEqbc9RUsh3CNrth5tOKpgLyx73EVuy9ybzck/wxe/+lh8qpMO1xgf+Q1TeE
f0MRYImkyMUYTKDZAb7BrzYsYVrLox5ZA/PtBZZdSm13pmMqDTtdEcnRk0E56JbI
sZYy8akAHV1vFgYQpUDOa8UJU83uXiJC8Uxodsuj9thFZxi2XZea2fzKrzxjJokJ
efi5crBqREzmdid9+ESFncqLtAyKLBZ6MUFvtqKNm8hUhfNjH+RnjJmS+WUmvlMK
hA06OLABV/QwRN/5sMID4hl+l4F05DzVc4ELa/vthFxCEuy1I7pzFrWZ7zePBKsk
PNO0DIJCuVl9EHpTWZGogr7DP5qJ5bzBw5VRflEHv05xd4gvSHMTUpePiSLT57zp
5DxhwZ9cpoa9TXGWRwo+HnTtrIVr7zHJKK1XyECm/lvscdxmVkaWX4f8Ck7EOklw
HlTwG23YqJ+1wbBqP3ws2dOKko6crepzu+d5TYx0MWblWkomDD8Y0a/MlaU5lxIl
RGpOtt7pT5pND+vIGVE2UhSLb5glX2WCoxA3lzwHkCyMYxlntFm53uotgC7rxPDx
tyMgL+5W8NeX/solC+knbJrNKgWpbDzZaikfoItuweJ7mU86vadytbd3oW/Sp2Qa
7yee5hx8+UgQFzHvuQs5iqRKJ0OqlSEHZwqrxJnWMh0XTw6oF6XBc6uRNZsqLHwz
MX3PYkpZLHQAkSh3n5sGhRQ8tYA4OCQSrrUyVUB7En+L68SnnWmyvOicKOe6y+sd
t+bcx1fPMQ4UCySXyvzwhtc88HsC0boR0ZRYPWqn6uIfYaL5P8mHaMLg/mVoZmf4
7zIAfc0RQND6Y6u/sJpxn19huV/HxL2bH2f0+nRLezNuy7OLwSl1+9PwB56TIv3J
9DyRQUwbdHmP9ejpZr0Ped93e0Lcw4s6XOVKsx3L1jUs1fFB7YGyrkjZ3CYsC1HE
pki8SPcfeKoUeDaM6tRneh87eCkvhVWa2FDMSTd0Wnio+ukFCWxGufG0prbYuTE9
WMqlYM7if6OpedO0Vf+0p2/Yx0mO1DXhImku8HY5IYro5SoyxMdsgbnmuiNiJ58H
uSeQffjuph40hswnmfVKhdX/xpZcs+NAhPIbhGb7G1JBf8Y2vR2+TGW2DrS2oyTB
X8m6ufUO8Dx5UxKF/e1FugdF6jE0GpTPuHD6+W7n9g46bRQ5CjKWmBaVsB5nEDZk
7/MHUcROI3Ou+Vu9s9a4sn6YikghZZC41nuYe9N+l10d3tx93TdBP3UDgDkQqh69
SM+MUVMo0Uh5winFUQ2XS6l8tM7MGvtRDc+i9Su1IljHZ65Q9UEkFR4D5ET5Rt1O
Lp1Ui44F1FZr/yPrb9zSllgH9kThJ17yeK6bGmygkd9F2BprmIQVua4qmdznVszy
Iug/eutqLbA0NOFmu+GdGu7YzZhSRTfOCcsQheW7j6UngTnWY0KHtAgUGxDU9AYi
rOJrP50NAoUPWNdARu6KR+z75vb0SHHswJjAQMACd6HZ7RJpzSJmRbGgsZfmdzTg
4XpI2sEky8C+3njzI5Liz0wnxaQx0tqZbdgd8cc3VFWK16KaY57Hq6KyQDvK3sQ7
gPXwEb/07ZSE0locw2iWDjE14zQSOAnovlASIJ7qidj1NhsbQlGqB9yxyn/AJ1Sb
/dHPDtdJ60EPPxbd9kBO9bSbRLc89/sz05gu3HI6eesFhukCui3+Xbd2XwraHuo9
QyS5zcKLiuh+dlG5RkzVVWwLxfPo3UkUc+YskYYvpFdcuS0KA3ZD4627qSPIDOWh
uioIWdtdLrcs4DTAQcL9gOA9vnKZL4Mi+qcKRf0yOR+8Rb6khfbMvDt3AevznVyh
MRmNNi3fEzosV/5ttLJrUwxjq0C7GnjAiGYxtkgRAAs+Bg4YcN3PMoGlQS5tLW3U
omO6KYbIGCKYtEFweadqCXJpq2GXcfDPt02ofslmwXWq0DabUvTtVYMBvSwQ5nSN
NOIww5V5afHwBiaEUKB3/NrIyjMeZWQNkAnWWLkFFENDpfBH7dkT+WlwrKfcorZZ
FRe9Ipv30wHVnuZrFRftVQJmw7bkMRsQmXHwN72LiO9JUhltyglYxYtYatjSl8JQ
oflhzQlyB0JqOSriKB24sY7GIe0NUfSWv151kOceHs/Od1LSLHziGvn5qVcm4UP7
eppMsP1g+JU49eU6zH5fBL/oDlcxZSbpuyciCsg/WgO4eVsMJu+wJdFmzkchrRIu
VkBUc8cFm4wEDJVlr6uEOVffkETg/O6WAwqOQrsUQ7FLpZIpLMlUQXfflqktHI7z
lr6+IOstmkd0J+IcPGB2o3rGddgP2g7SbYGEGuEnJSG7ueVTDfG+ZqPjIjktVh4X
1yHcL3GumQZTjy9NKzj0xUK+az5jjprtttCze8om1RcDnm22ybNdr+jisHPEst8V
B2xAIjJiTJOplr+P+b2iBBCWK0HflFC9I+VyK3tXyhm+SFe7MzmXbs2nfszLsOx/
burlai0GYs5JdlViv9GQHSuE8kd/a0Zy53QYCvL+yUS8Xatkp4+HYUWfZ0vOcUf9
plt0MHP0dvPKKPh4US9iOofKwYQYd38rkCtJsqZsYLF95nDEQ7bXQMegxpJc7ZCu
/7ecN0ZPRsw5z1QVV3yUs7SA+x7qYKvhZsdnaoryKq4xF6JhhSXvSsIMTDAMkusx
q3WyI4BWtAb26czQf8Vv0aaXid+Wm2HYnx2nuLLlValjgKGbK3LFELbMrzfNCZHm
SX46silagdtneSjmIe8AB3CbIEF7WOwggRrAJeb992e8jc90MTuAvnP/B6VV2VbP
1pluG5EWMLe9qlbVjl+EvRCsoldHbNzmsVHPc4EFAm+tQs8MRLXcLzqF7McYC+eN
usMTrd9YvEUt63e2q3Y0S2dGi0GjiUytG2FQ/7Yid/lttWg2UweDk7s2XPvUhCXp
a4hYvmeXFgUByQhhdHBV2lT461tUp80HOBDIgtxGATxefYvBZqpR5Z1JK8A+Wmja
3Kw9sCS1TD+ua0qxn/ki8UckuwfAVnZzpx340ThCEptvcF+La72sXbDaHRMry5BR
FSvs6/PDUi+FUtbhZ6dDpGsYQRo9J/rM4X3cF/ur0EOEhCuASS65/AsE5YPz3J/F
aKjQEMGXkJii4FJ49Zrq6bupE+zxJLX6bfQNeumfynWHH9OZXCuGmoU+Mn+7+nGC
Mpq5tMBLF01mV430PgtWzTnYrPrEojdWXpOgI0a+v7bCEErvdGFPulLYyD+90yv2
qn3Utg+hYj7xrMpfxsnF+kPnlhd+l5DHmIx161p05VYJOMtVbVBWX0pUGpPJntcV
fMG44qGSdQM9kiadezVHtl42h8MM7ldvyQdgTPfZYMbIz23CKYc+7nI2AJneLoQo
aQ1DC7Ld5Ou9PyBW3h71jqaTXMgzlnpnIHVrIR1aZMnnVEl68PrSicTXuCMISPud
aZRI/VnOGuZ5oBRshVdE2fz2IXD/oktlzbQSCSgNV4BCuxjmGfHhzHXCOr3Th9bM
oc+p8iSWvOQEHJ6MkfYOntbUqW/XuDwsUH61fNSxcaonn/c0feXLPLCVXAU+JJkn
8sdKITYLfLNL1vh404npetiZQjuvHrxrMXt+dCCUk1g/kI6UDNay7vHLWU9+VGOu
OlAVw5+7q/CkvS80p5TnG/1Ymf5K/dXr7MWyYxKmOiJ7JNCPTbYSZYr8e12u9cUW
5uDBGlbUidr6/FoSofWoseKt8JNm2s2qO28gQDmQEpo4wTDHcB+SnNgYn8MaBB0U
NtQ0thKXZPERlsp7LWGLK3t+/ChQ/NDO90/6QgPZ5ngXy9vAAMUTTv2NoDSsEsni
PtQNRVK8prpcD79Z338uTnxDSckN5kwOsnqOMS5OUawMuThsj6pWTG1GGI/8KNeX
xzffU2jsKDsNjx9SHrQxrYlrud8LpxZOmahnN/ptESP2Ur4xQ/MUZMnGD98qp3UJ
7aSU7fp5+CtJsMhKN++Q06GdiCl18U+q3ErDr4XTqtcUUsGfIOPYhsa1WDdaUPfL
foxBsoYNHYjqIJCFt4KCwLKaoPvZVYztYo4N5H2FyGT5S3Y8nlmZ7B3yjOVRVln4
r90QGy3Jxg/XdsKQH/nlpY7EZ6vFbgmHkFpVsNW9IOu203MpKVTzL8zMfmvhXrJg
ZwS1Mg0t3b75/PYKxo3sypTjLRzTrIxtuQejU8N0ZP8OQQKrKcKswnKSQpk3IorG
gbTxT41FSWXFMulQ1qC+aJmIBM0A1qb9Q80hagsCkbhvwNv2rNLr+oWoAhdPI4+8
5dQPZ/GWKKdMdms1nxXIKuy/aXLutBN9XGXmQWNoHmjB7y6oXTbFJpSRM4/VNmVN
5DOK81FafBzDIIr/tXhWHrLjXwMbvQXWIXB+z759Tc6E+HK8/jp2ObNyd5ykZO12
o0prPnzJA+3YLTC+JsS2DN9NXtUJhshsAqFKv75BOLe+p264FynOjw2sjuc5+zJz
cLCFUOwqh4p8zomtU3Uh5FIO3lbeBIFKrnvQz9DgrKxH8V4SK8RgdHOZ+/J4MGFO
BYQLpYMK6BhLQ8P7zT8vnSQXZMad1tkBImPJo6YUu9DH9ypboKkJuPZLpAFWbvfB
Unw/WpiVaLJf5/tdNzPc5OROq0SJ+TyYiWfQeWmDfFICO6EEumyYvIVuy81dlGYN
H8qIj4vWm/5d3FtZ76IhaGR6ruFagv0l4ZtTKj/4j+849jTDgEIrEyD4Vkjgo6Et
ag8J65DvENrnMsOlq80K/iuGTlUwKr5sdneIuLYHKhdtjNp1jhy9DgH3IkV0NMeq
vHlZIujrHz8ihoPZRq5Atm0lydZ07BuiL/ic0YOk4FMlCxVU/C4TYeuzj/CVQl+K
fhO80p3t+mKUg/hjnfPIvn1Pra0NDAu3mpni+0Osz8MYKvS0E13dxjHItKyoJLOG
Toq3kEJgOFSe1jSJfJsrWBdXtSueGYa+NGCZ08dA4iqRAhaLrHpFyTvrvh7RdDhC
bX7JcOp7V4n0a9eopNhHgZpYpDpLmTZOZRT1zXNzI/GTwaGTBul+C7pqk1I323jp
qBMxwqL8PWXqZBsccpxnUX6FbuIvhNbwmjTic+J/goKsjVvs93EXTME2sbjCkd3Y
BDlWULTRg8F1jWxLLjBYk9UvHJs/yUTMsCWgHz1T/UW24DRwpCEXXKn3glmPDqav
uBDcl912JVx+sZuD3eLphkPQVTsHimgchQEsex3JDtJzOXUkDxJVX+iw8x+Cqp/v
rRN762OWNRB8LE80rHjgaPYvAiWmLxvgn6evM5+ymBYG/gcP/vN7JArdjfdqa6TW
T5G+2YOimVpnGLiLAkxruNMBzqjdsBjw5cmYsyQbtbBN2MKoAv/zrnEdBA0i9nTg
7upMTWuPq+VBIRqA0Z7aUZu0vlOeW8BEyij/ecGur+Orl0VMmGxsq3LKTdEoZkIW
Hf3huaXIK05acimlZhYv7L3UEEnvS9tFijn1iy61oFCfif1+1+V6uA+xFHx04lbh
g0y098Wlj30ei6NXc3ax4lE1v5AgNu1A6T+GpSvjBrZ540ksDSWhdu1dCOuFYqAg
Qci6pcm3HrG0n5MlJFQ6Exze109HAHpRYsN4eHUG95NfJHctu2+RV9PoUYgVZp0N
dUlf9srtgLUjKUz98J9dOgKYXgEk36tMCoueyuZVGBPo1vlViktnj2uHDS/XZX8m
zL+mrMX8cqs4OUUs/WHemVWVm81DzuM+5NLWWtGD77YdykVSk6HjzP1r8Nyax5jp
Pynp6BbJ+cNMcHf+I/xT2XeBNxOsbEoivOjGKub7TlzTcJUdYtdX62ADT2x/Tru0
zZo6w/7sKM9SoL5u51pTktPRlqCDggZWcLv1f/lPjKVQDb6M6hvQaHMTUNoq5hZF
ViHLLVom+WdyiIc33Mj9AOHm3UGsQlHSg3ejJwLccxHEDWl27nxS1xt82CjBPC/M
oVKgO7py5W/Cppli8J+WO0abQTYkjfjwugneAl1on990ZSZO8M6CB7wHOVnfJHeW
wBLvVOXle5bV3UnpzUbtXUPoJpLFRgPCX6IXIqp3pYNpwUJ2/mAa4qtPFaCwlN4S
Wt5GkNaBkgWOGIPFwvfPrItYbqyYOMGxdvf37GfZ6uoZwczum5stezrMdLN+rUUz
HkJ4FFwwwH7agTlAeoyMBGYplxLKeHBJzxWVVu0fAQB/H6I/AZC6fv8jStNberKs
/dvZdnwWXWbTNy8dt9KynBeUvyq+JTeZep++KNsFTQITXNrfUXixDYSNriMZ4F2f
0HKMHvdpluc4dnCvcWtr07IQd4y68E0IvdLkiDvvNFtLxi5zVgZj7J2MRWDGMCTx
Q83IfDL0wVTXSI22iXysU1VE8zZ5ztMsRKuQ8aWqTfWepr8yH0v1b1tXU1vZjwVd
FATf0ulIqZB8d/hkjVHmTYjWQUonW8FqHg/BIfYPV0MfIPiqT3K19KQqn5nyK7eK
GjNqetwrLjjRM6soKVXCs+kopF7Bj/Okst8kOQfpn+WfhuxBGRZDZx0GhQdtDsjS
CEU4LcviPx/jqzVUzaIFrSy8oo4av3sbKFo8N1zihr9SB5dnJskw3Byte9CyZNDq
p93004hlDXJVk+JMwSppkNG61Q0a571XSaNy8JXZ/0z3/HFlwyaprpuvDW3QCoKa
iEvidkW/sDO3bAh+hJsCw3NbCpC0zOTeCXxYYrNTvq+Y6QChMopKhgqTxmGOHCr2
0dV/guwRziEzSTn4IluWnrbFhJSLlh7Ztt+j7Tqc/at9sWjGkJYFRhTy0gOKPtWS
4l64i+xWHwYxTIQk+9izcufP5OdFvjMZCA0vIqPbrwmWSpWWhhF8m+OUIolJBXZ5
8oAkZQ5tCWkUXJF8SN6cQRG0aCjj2Vt5RXVu8j/HUCnxCjbXvRr+4JPrYSX2HWMo
8eXHW+sy0PRxpIIbJIoW6yRdqeaKSTrd1kOLF4be1VbisopFCLxvVYVDCzZ3kD9w
CHLQW4ipMAVBp1GjuPJoATFDdZsxILlNooaqUkc+crN45kHeubu9BkesAUAH6QYP
E7sj8SZdnTf19b1hVKNB8v56MnzxK2ra8aarqqPbAe22qVaE6Tj7Yaoy5sdrOIhG
a48TeVubEca/7NyCf8O6R0y0qQm6Tmw5sh7LT7Hn1LZgw+ocG6zv+SaMACSEWcvm
AXl7GNwMG6zicF/ei0+hE7Cgtq86+MzfvGvUpL4fsMaLRbvnRFmIyxUFOeJdHA8p
06GJPAgVkZi/kOfPzp2yXJtpHudtAz61Rr/2DM9Q5HxqzUgmpGxNXmqHcBuggnEt
kbXgKbEc0d6XYhwe7JGDhEH9OuPgZ6C9l17GcR+aNnwuB0tjZWBGNEEvZPREM2mC
9JiK4oIq3gapoBZqFojUNSaqTz3SuHh4nPTmLXI01fmnxcbyhtkqOAEmmoRUirJ3
IML/G3CZq8B4J5wP3TtM4Nl2zu/AM84ekz9dHiMrCK6L4EQKk3f+4ZE9oVD/4eCB
nMk57WsrAJh/mkz7mr62Tlm4melBOuFnMVH1G6+oQEEYBl36rk5d9Z1EC4xyXzjq
o0luwAhdBf3gJ5er2GCv0z93FukW2u8Dh4YxkFmaekx/AiKXRLixcnoH44p8IWdY
zYASAhvBQAfJ8LM+DpQP/oyNummdjhHj2BSpbreiE1+oH67ILH+CPrRr3eSACFMX
robSmmwFj0Xxo77pYYmYG4SOkFQJbAWo9+7/JMAW0Ql5/L8NJ8FNi58ayGXP0WR2
NCnCDSRDua5HdZBapMKLwi/G+XQA7s/Wv1NGxmBcx3FkFad9eIG+X6FyehtnCfba
o4vCUeZGh63q1x04VNMtizmO4Vd5Yv5ukbyVBq8DZCjXsqWwU5zM/RFNZsIUovuN
Pbd4asl/FQGUXe9jEfDnpXURtkWmMvoaIPEqaRE0C1Ugnzd/PESeuNNkRcH0TcBD
yga5pjY2/ASSZ25hQsNhqihXXDShU6aO1PuvYe2tGZ6Xsq1vtegLa6x6Ii0/wFJl
MQ15fibGYkYf9UdZo/Yed28zRjLM1jBYH49X32tOjOUq3fxoA3a+A+x3Q555Tr30
l5JIoWAdQZxfZ8LqhRM3sKydOfy0bDBPRnsOd1Ty+9Dd6aUtjF3YsFeqTUoXjEny
oUOTdSQ+1stb0aGmegEdvOy/NITAJeLx47zh+GJhPF7JblWG+719/DeOkhVM1bWs
9VkWbclCQx255tXIKizX8x/Bg6D+sEpBFow2HycSV1MfUr2OqKls+E1tclZtVV27
KGrfld2ppjlPB3QJunwJhdw1OekJnWdjptxzC0biXgOVpm1Labva2a3FGYIihi/P
CdQB/yhYj9CYT+bfIrF93nyydcrNtJKgGZnABg5D1AeX+K9V0Plr1g5dmCLNxjna
tX+wcw85MNsozV16dDYkXw69Z1JxlOqrTAIqtZSXqnpirnl33x0A/f9PyeUgKmzz
WxVonhkXEIQ6sZbn29jPULLOl5H3i+MWCWZplm4ouPeV2YSdbqkapZkq1NZaAoYj
Hza0+/ZNxFXviuLGLiju8JPIHPWYYYWgD/9pQvEqz4up4EtfJ7TquuVzXg7e+yDA
jvCS4njaRms9PCi0vHSHVb+qjiEftdSmiPhmJiproa0UpLWBw1N4/hLs6BSMlB1S
StfTNZKfJI6ZeGoC7BmkdtIWknNn/AZsp+uOXWlwSNei0XOOY4cBU3N1g3uiwbeS
nggc8E/P+LZjQ7Jgxke34IUnAO0F/RCu3eNBfk+wQnR8YvQzhRE2WBT7DfV8/buE
DJYRxJVqwgdI7HKW5KePTVsUJA7Eahue0wuh+nkdFT8QVpfNDX3RpCVQaf+kiTNT
xC5ap1B0gVtC/sUdid9Har0gdrdA3I/fQLPE0hIWmboH4PZiRQyySKXOO3Qyhyrj
zMPMZon0PNcsNF/VTrIANCbgGoBmb6oUrO03VrFMae9j7WQZD6NlRkDv/+Pt98Ak
mWzWaYCQ0cjwOWfak+vlAqria4g7DHpUxqPSs02tkh26fTscxDfmb3ZGTojE/hue
PzzaSYwpIYRiPMD7Izrgg/jZNTEw/axYmDps+lIUfB1p3puJJml3zxYuPr7kGjCm
007ZQye6o7ybvUa0sVqxl6ZfT1HPRPkHLKFNfnpT/Hrj3m0RAJmLlx8DYEPNoNJa
tGgyU1JmysW88R0sv/aXkKo/j9cpej0LvRt0SpeObuK1MIeAt48rJqudZuIexMbB
aG5yWVeSoUmCy/84T6oy4ptGNEwWU8zZgmrytO4gbtWMqkxdj23fci2EdHflBzAS
qQ2jRsjVIdgHGAfPKMoy3XAGKeD37jmgT9aT6RXSCSMyZs6hWVD7MWh48IxbBkXz
ZlcYic6zfEYShKRPLawTf0gkjXqYYGalPX7cSZIq36HS63pIs7FgRgkHY0w7OY7Z
e6RFTqHDo7MxW4awWGKwC/Vlnd+7CwER/luWtCaUPORQ9e/lgqj4Z48emLxmQEtW
3P/W3O2uNDhrKjv+0JB+6fUstJVsbF5RL3WziAi56paer1+VLN3FoYqOwNrV/1sF
v9WYEWHE6P2NZQPU2QkFoliBv60GSpW4blst93weVQC2lqtDaY5GRJsX0+FAMGL0
86ngbHE0x21pr8JGY2oczrjFwUpTKz81WTAd0evoxKAdCQWq09SaAhx1cGDD2v6Q
RqM1QaEQ1NusSVl9Wy2lKtknqcfDbEedrctVF04Y/OToiP98I2KToPC2PI5B5XmE
9Cpv2sC85DW+Df8vfrbtBlaoFSAvpA6UCbgOmbuuralnkY4itros/yOloz8jEg/T
VjnVM1LfFdGBcPRKSVkqNAA7oisNZeqwUpVtml1sBWEG2ktv3kU9PlLOXjbhVVEq
v3hQZTNrWQJHz48x+pk5HWyIUnHjSfdHIwoj9PIuFUkn+Tdc0oWjEG0uyeWp6C2/
1pqyIrK1F7C97EVdriPCY608dJwLPy/t+XrxgFaunYtk+2hyJZs+guERuTcbCj9I
s2X0MLT4IWLedKIKB9mrqDQ4/9L5Bu/FbmF3OyZh2VxT9R1480SjLruNB9tQr2Yf
U68YPzaRaf0sed+R+0UuZl0m3bYULPwDd2rFjc8tQGwYPGxoTq9ypnBrAhYxB1aW
OXBx2Pg4Ogy08VMBmcf7TCKnERBKZyH5JRX025/xTXD+V+iWwR/7OukyA5JH9kQ/
uQCEQ/UUzys4IKJiJLTIlT3rhADp+fPNgkp8mK4dWf1NR0OWdGrUZ+NUDxO57P4Y
QnFzGJSA2EZF/msCBIJuNT3INMxqRvp+OWw64g9HXwKxiw7kNmApos8a/lNaHE+i
k9Wec94fDW7ld+ACLaE+QPtDAbNCOCrHiH5IU+8JO5l170FKKjBev5JR1ZhVDh7Q
Cl1pG1Za3/OoUT3d3m2saPyyurT5qThfCkaE1ACl6+PYiwa88xiwvHbNUaW9iMAH
Qqnij/ALNmsTji+hvIMn8m/9UZ10r4wkSjrJdk7NbHOnVEX2sbuEMkibU2w/GVow
93BQKo/Wg1s7VzDBKvZ7vPJNNukPq9RRnRxHo8Umd6tsQqNDIkjdzIZlyPQSAmZ2
cuO7JszL/PuXe5/3AZkxeXhV/uQW/QWBKQkHa7eGXM16fu1YoGISn895NfEK/96F
EptcdXg2c34+AK6DPgojLngxs/xSc7EdxhuVoQ0l+V19m2iqlWksnE2km6AstwZh
r+HxwMuxesYeC9maJP84zcRLe21pJynEMEEVohQUmLTW9REKCjcEo2+TOC+4QtRs
zgH6eXTwinbX6d6qofVfY+TXslUN3bN7n26T1FvqfwdZ7nnUTgrrjHgm05ghFkCJ
pfDseomZavcyB82FGCJMLx3ZTthGyEXWEMSnRi1c2fSR9iv+An81oRdK5hiu06cL
mqiUiQHyRtQt/hlL8zs2h/+Wxxe74CjoaayRCSD432qz7I7xUjHMJ4MY2sP7XmUG
QZfuu+FiCwsXpf/eJIF8cI2YralYKCfCRabykZ4uQGGtBwdZKQzLi1op7YJ5vgDd
GfPGFxNCn6zUe3NWthceeavmAx0pQUFgCKaxxYraccXQEvYFdDq4WFEb6L9rQA50
tpqxy0rqgn68SN7zVt5WcOiqS0ioGptzrSLVt35mVsrr2ZsbFJ8E47cTFybkfGRj
iK3JtP/tMld8aZkeUnKkv88EZaGxYXjkoFJn1SDovhzGhZIP19O3xpHNQvGqIXCM
YD8er/JXhwUZeOpn9ag2oeukrUj7VsjVRldHyUw7lq/tm/0nekySA6hwHFOdQssX
jPveLllKVl6n2kSgRc0DsDb4Ef14wJp0lksRet7YaNvkCB+sZl3eLDg0skQ4MpJ2
VmVMQCu4fnXGyO7QveoWPl7WnH1h0PPbvq6+hlOvy4m/sc+0pxjDpFNTQkT5rC0B
lzVqnl95xHpWn+qq9EKEEMPNOCoNAaY3cLU/DqpMutdCJfoDgg2MIVU4YkcGCHSI
kXj/9osQlLNp03VJci2lX+xYkKXi4ljvBXYO7Is2UFA+DUQNy381wK4N12oD2OwU
xqqh8Bgh7T67h2L7HAP9ZsXW1ipAOZzuiEr18P7AP7xnKyUivCxE/ctONfKNH7Cg
I+nJ1z4spUR4ze5wBvWohSxDWITPmppR7bURxezXJdvpxqwJD8/PsJ8ztjv/sQne
jEHlJojqEneitOS84SdtqmBoizG6NTVcXZE4M4mGYSLWAOIyLbJZCRcLnFJnmqqv
WZ7BDS21zdtb1Df4i+klYSYZKtl4QYcD6sM5k/um+guIIWVR9eNyjKh+PHN4qRcb
E0KR63UrL2Ud5vvq9I8CrrSjrVOart1P2RyvB3Y+33XdoefGFPckhGjlbxeM4SEZ
TMLVx6KBNPVYan5Cg69TUGjDPH/s0jNA3NunHazQl31FqXBccebpRI94IwyHyZov
idBKEIUJK06LabMbrS9mmSwyJfbhm+PF6v5mZvyWkwtiDD43aIknxlf5kmQ+6uNK
Ct7njfINQPRPFMZGBrrrQ+Ab6E+cGStO3FONQXmWqnN0eP89RmwNd3M3CmqDQE92
jIesP1B0dAJrxuiVDFWuRmwbSs2SLxO6Q+A6QAC2add6J8Uer3uDEP5KmpeDPd60
rCmrUFZxvCcbpXeDXMFSKtkIUWSh0WiUNUuwmHAyAR1VhaIm3GbEk8NpgXE6bcOo
TyRVQGO5kt2HKEcR27gw98OSx7/M5uztggFjjsAXjvgWunkAQxiuipeQrFMkewdP
pJNtSCafzZGi4FDQvmYJBbEjp/VmKm0ylJyRjQ+xX4fHO4QiqS8927/8qMGCS/qM
BwM4ceH2qsBC/a+YfHjkF2gwRIcKT3kYOMNJOq1kLB6XP38PiW4VyvXWz4ZGuUHl
IA1JKS5uE9yK4VZySyRUWcTYFTIKeErtyJnsTXJKaJDbr5mSX+GhrWnq5KzX38Kk
aMDcVzqI7Km3rF1W5dxBRf2exVFYmc8gcQQqp1hgI4TuOBNBV3CWZpBkjd8JBtTF
icwt++RI6KD7z0n9EI+ogXbfsiwf6GKY1vUIE9bi0afOMCKOflMzQSCiAKTsbJU3
qujv/ZtZ3ZWCv2eNyzz2mem8YQvWA3tFwx3ACV7N9Q5aeGUrP9+2CwNGtnEpTjZN
NmxQ9F6GzhG0C8HlL8sMkUEp1SS24xqLPFH9IbMvogseTOabyJ1Cc653Gkq9urku
ygAY3sdT90NRixiFCHc0vtbnQ1QXodipmqC/FfSHUlMVdHvQDAJgkWcdjFTvEeCg
7YvJmsxYTewPwCIaDosWQa5wEKkiIDK5QBUftXn7CKJZztFvxG5Bp6kW4YwhltcQ
+cBUB03jfsHP1FhBlf8sfVT1jLjpWoe/aUlOoxY36++ZuRaIYgDh9HPsJHWe2kFR
7kFycsT6oMFgEiu1aTIyWyJ345Bf1tiL0Le8YiQGHjFfTNABLxBSSlwNXzTJAIrW
Rq6VWNCu7pCwdoSr235c8oCDrzA3suvg6kdnUl/qhN2P7h+QMKCRxHe9xkMlOfgt
SNpS8xgtRK4aCJ2LUhH1YC4IYQNWq7FjecwgjSuou5oqahV8gnAdLWpGCyu4aIbB
0ftLUQ5/D8wtsYN0TObIdNDFh/xflJWhvqJgPisLFPrt3qj9k8aR3Qj3JOQuPs+c
9bnQHeCRpgZiwySOpmCOTUBX1CkQKR1LcSOh9bMAiq02oiz79hHvODDxZwxE1pW/
z2ZF3CYflTC9JWve/v97YlRGp5QrIzlkik6m4Bbj2WPVqRrsLFGA2IPG+15gE5mU
02KVk/sF2aDpYNPO+VAdblhgJCrtjGftZqB9BJPpN6Po66T+lXwElZBxF0Nv/BL0
TyF/UEFt5XrocesMBHu5ixcTdzerRrMItqzZ7eFYUZqcjhPKivxUMbH/233eoLhL
QMUyrziBEe7gn0rUq0pbzl/S6d7EctiBRL6ScO3EqxWMPur69/b1gQnTEPn4pyDA
OkFdPFgmujoQXefXPaza35O6EbfiBoLB5sI8iFGV6JINAi5H9X67O5E0B75iUnFf
yGeO3rJZP2ZmaMRLeii4VA2la4+nbW0F4yBGjNb0nLmEskWl5Sqndf8lq+bwj53q
YKSbGu7a8SYtxM6Ad+TES0A7j5oIRPNakpmjFNhcOda9s3/V9U+ADwBdgvR1WPcd
+krEnLEY57K5tfB9YDT+mVdPmQ3TvfaTpS0D2sajSp+dhtaheywUDI5URzNBjb6I
2Q7bjmwBo1K1ECZjMfjnvvdmNEZPttAsW+Fn9xHTcwue6daD1SAhRjq1qJ8rIPz5
U7OgVU7Qyju4n2LUbeTSQlSbPj5N6uulrxL1VBTOOJF4AN2X+z9glCPS+aJjlmhV
+kSsquugDlf3cN7hJZk5ITVJV9qqXoRTawxAe4wby9H1gxxChBD+X4Ha5B1AmxuH
XUCS/emVzpLI9lbM9Rgzn1hyzYfyKanNM5IMaiAd+hBZW5jcNjxKK+G99XNPNk/7
wfkCie91YBpjfLQhgzSslq9XXRUAFoeNc3Zwx5Daq1QLhZswtn22RNgpjehpff6y
osHf4aXllFRH5nw+eCQoyF9wKna0F53YLD5Q55ZCDGMpz5P8uyNDf3VGjPKctzm/
okkhM7UiyrFQGBwx7BMybfc2ji2sMVVdkpfKb5a4l7oL3cVk/HoMM77NoRrK6B8L
/31pmZs4Qj+LL5gGtmaZQ5JtDXT/5HNtGwBRL+c4CoVDFpxxb9shsD7iI/sjxWVg
JZmATPNJc9ZyOTDG+wAHD7r3a/NhF5Kop7sBSqGVB5hJDujLLgb/qlWsytWf/EGM
nS9vmtTp9JdF/G52zWD+IOcj5LEu/FPBH/mOf/JleP86GEnyJ78kqIXU6WMhQnJ/
/kbB+3uJX5govCV+B4nbT7WHsc+YNeHB6QHs2cDfewjRnNWDANtIG7EisSOOOCIk
zyIIfEKigiXspfOwU/T87kkWDmaSAYpBf85U3fAZOAs6UmV0DyvtEmVfy+a2eLpv
SZWEEZubxXHNYoP2s8rn0O5T3fQk094o9cvJ+DG2UdDqCZVAnpxJptw40P+KCxHX
f2wMITMqN4q4XaLc02RF9CtYIHSAGFCh9ipm0BY/KEh+P27uHoQrmo21Eyyuu0mq
6jQWoRnpJyiv656wujDNhnTkm+aVShKo+Ytvg/Xx0ouV0XagL/r7hAycTxj21Wzz
gEIdORM1ZW7IZ7FHHSNJqPU5TwXJRitNcWUbk48WeSArrn192VDLJVOWo91RmVTE
Mo3DCfRfvyyjjV6nLEFU9LzVHzPSzkqTbwMzT/wea3mOATYnldEtZPqFqs0NOKox
I6lgozW98h2/+avW6Gg3PImMCZjbubIo1hF3NvoSqlJeAQLmh2DEJHQuCZtr/zKN
0e57ZPoQVDIPxzGpwCP44Z6tEIhqAfL1ECjaPffSHp9XmAa4U0wY4+9ToQgU0KVY
GTOTOscCu9tv1d9U2zLyw1f5xnamJTF2RDeK7/OJofm2TyNvBdhvicExrPHWAPOM
yDNt4ZDaQ2Ialrbo4v2obBlyZ2rkI5svLmAKVr441FL/HsOa82H+T/X9Ikky9ZcY
UgY1/gQhcnwkTrhzCr2zmg2PyFcbCdI5tDneVzeNhGtsIFwhGzKPsmwxssJQAEz+
wKx2gOd58Jbee5gjteTD3/Q6+anDOMzuwhnNofhEUlUTZiLbAIBX6t4ZWMlC/BFM
Ld8jALl8dVCTjHsIRzGrsI8ziEbxth80/tsTzKI9IATZ34G+eP0vqoYo6t08yrKU
uWr/K0nDTJiYMIooHRYwOjMf4Upu+P1E0mpi6BUXUHEcsDUxvWkCMAIzUagf6RCE
Ik1+bE7juRrEqG2knhr/WLVJk9Nw6OrPA/zeDOJzygUfcLhEMEsAVwL/JnizgykN
L5m3MUwHO1jLcMyX6quy04r2et+hiG7nHmXAnIftPtefdR+olK/HzijHxpVJ9j2m
N5i3zQPH/4DY8mMqpSlUkDxaEP/RLmqs8507GG2e5t9fZW+3YHbVSF/9LLgyZO3Z
UwHMHBzYDBbGl6AMGns8AAIH3nciMJ759LCIKJS8O+HlluzMeGO6kmbV1pzr0vzo
q+WNp9UwZ7t5WrjO1zbvvQZl81Ii9fxefF0Wm/WZWvz12krxbYaska6VwqI3ScZw
5QEolC9xcIzs/8Me6vQzZtG9Wj/j8IGdyKXgBc89noac9DiU/uBCVnt0sEBGjOi7
it8nUHFiiKXkLZlcyZlldCf3eAi7OQg0GmqOsoxb5evphFsiFJc5KFqZ8A5Gmctr
RCKdZEec1HrVwYQ9r6bDjrD72R4J3X1tALy9VPSmrz5XsgjyLzkyvW6UUtV9BJlz
Afmtn8UwEt/IGY30hggUFPBoqlykC3CMHeuVlSYhHRc+aYIsGMxYWgrq4niI+Mdl
iCMF5USjKgE9QLpM/QmGwco9kxNTEZARAQdWctYj2T2bDtLbtvk3Rhkm6M4yJ4B8
xXvFMfI5Sm4dGKiBSSAoh9vX0w8+9mWwu9X+9z2tj5DcjscqIcE/Pj0cCMqbu5mh
ejqf+HZt0DNkP3nunMADC+Jbnc6kJsRlKCE9fgJ2VEaQ3bl1UT6tVAQGTkBQrRRg
mMl8bK8Px/koM7hxY9unmR1XyFbgNoTtHq1o8Igkp+rh6PGEyZscCUL2wROCjTCG
f8yz5YqMWx+0Yqb2rEmUDMqN7q9saOuaWd4fmuIW7CDkuW6ggZA9MvYswQGYg/ZJ
mnRannPEiNt95afr2B/BCtc8DrmOmENPiz34JbTlvzt4eisruWKl7AHFmwmTNgqA
/3jH1LXe3/FIt+Fv1MMKWLJioEr6p+RLuy6NXkJTCMKCbB5mryo5+1uywwf07b/Z
NTZsxfV3urShniZJ9lp9Mniq3/XzVSI8b9DlQJdIEh+S+bm1MCXRu3Sern6cZ2aR
7mZuaaB9rWujbSIReHtpjOGQ+IeSLYxLUL7Zxc5sxVnkQsuSmUD6l7rfdXHIzxlA
6ozHLBafiG6msFsWSbWRIvT25zRhn9CDjM5wdJvZ5JInqH3FMLbkyfxPX6N6KhQc
EUTc1s908aLQ+2Ijpke8Jy5LkMRCdNHvvWPxSVhM5NutEdV/6hyqgi6dp/Qkle6B
o52NicuRzRDwJtA+89MnTIW1xepo47r2WRx+g2ktpxtpZr7jNwkhl03b6JgVFctR
+DHHT6sluruNenAVosTBt/r7QPVG95/m9dZ6fGjNYItnk290eEkaXJKxL1wTZDfX
FGEffzTbyVTB7C3LaOo6zMveOkGWuFxocVg0/+/boTQVYJau5kGuZavpva7kBwJ7
9bj/Wuslf2hQwqZMJSliAImrA7+InDjbNN+cUJW7oUfTihvn9hM7oxpoxGlDKBQF
EsJdxeFrwuLcuqBlnkddxKJdq3QIPq/C5kr4L2dw7Mq+ij4UnLtgHtS0K7BLMZVQ
BM846AjbTG+ZngdGF8umjxl+HoLk7oZ6hbJd1GnH0D6RhtbKUryOf+P9MdnB7P10
hw91Ut6hcJXDYe4BCwSBkMDNAT9oQrCsLeZRZuV0l00HgiMBDfMBdl98FQ6gNMu5
LLHCCQXUyPYMtm5RcjwylJ5V4HwrKGHtT3yqF+iNIZgVGjSSbIlRJhgaL34+A6+l
ulfivr/YgKkV/nWdJ5H7vwIzPH128bK0QRm4AEt5aVlXe8J/3Nd7kuQBDHG3n9SI
IOODVJ3PKtUT+OIuRZh+Q+FRYtXsPslhpPqGOY7JQYHlEcT2RzmlTEFvCv4mWtBK
fOiYVNQgD9J7b0Op865E+O0t6WsxEACWg3J+ZFT6SVI29VdMpHhaIjGn41j1fYMp
tSUh2Rm7eKZin1KdXgleTVbijEVob1pJ0mxUkEurkEhIAJLktGA1V061mqkVFjss
ehtrqFRo3rZL/Eivu9yfEIkyffpP6n9wB8KR0aqrMpgqOXKX+11M8vK6jNgzle7p
7LqzWNxZ/7NTK+HSSPaCKZk7gxQ8S26RBYn3qjxX9sgSRfZAGYXpjUjVXHGJC+W9
6IyM/HByZHmshzBe6u1M6HNulR9nNxRS3mR4qZ1OONBR5p/UYAcT2RE+c2btrlPk
CsoH0OeMNRu2cwUdxoYAJBLaVPg4HxeFKB/YSqBfJd1zH1vTrLaOydCIe+HGFHTA
hgFTOSBunaFBACYiGVi7q+6BDKvH29NF5rEHXbR+0Cu1mtxFx5IqVca7R7h0pYCa
KTNZXhV+XhHyXAOJsV9Uw5PNF+vUESU4USXBYj6D7wc0IlAlMq1AFTahANO42Qp5
pEzU0NgV1F4A/NoZcKDnASMzmJmCDocYC9smPBqHvDRghvwFFqNsYuLjmGPN0l/D
yOKDR/c0yq8FifWHRYTrIGAXSBi5tsHgiMS8xrXAEMIzlb3lEXbmJvHd3JLWPMBw
QDwHocNhuAvLFaj36ss3L7KGDV0zAZRZ/EYUeQF1YRduGdbR5CM2AWRqLFqlLmcE
IoNNFaOK5YXx45+9luJvKqNAjTM+YAe9+IYU3GBxU3E0lwu4xkRLePu0ZHYkjOWN
wO8vTrlx0sxIo5yBvK1iuILpPzeu/wuFW2d1F7FGrowQ0fDK6QKcOrsAb7g3FUlG
OE8QYaGmyoEsL52xVziaw6ZS39a4K7FsH/BlvlWQfdAGCEElpVXBjDwJM8KLqLt5
KUebI68hAGMoL36GHSkirnCcgAHMaVkktmk+gatAH6PMicroCGj/SDqjKf4y/JtF
yMQkR/ZH9hj8L3IPet2TF+nh79iH2eoHBM26Z1bFeA+xHhnfuTQV/CaSUBOL/ZYS
4OW/9JXOZ6IU0fJoR6MyBHbpBU4UE0tSfaLCRkxuO7+La706btBVC/J7WWA24CMV
QK6gsg9gh7sLL0n7JUm8UrvMRQYVoMbBw8u02kcZ6HP6gcSadXJA+abMIMhKD4Rz
aaBZ7hxlwe/00HvjApUvwYoEFHS98/rFB4YLxFP8FpKQw0TvGbjn6x6NM5Jr9gVU
PdXjCAfpNiJ7sVDCkAAiqUOTaWrgPEanjd6wqySackdSUqSkcLyv7fNTLXwLHrMS
PfIdhGl73tjYFHb0r2Wnmp5ssrg5Gh3pwBGHoWUdpQKcXuLfcKpK0GRkiqr5A1VL
vhg6FzlYy3Feqkl4SnTlWlS48tWO4u6MMIQ7K3VTKIES4971Ax5rixiiOd9yF/qd
MOwI1YmUaQjDu8HUNSgUdu4slVHanHYHK2G5W3hPYV606Y75S0yhiOISw6NEp4PB
XKLNr92tdgoHIrkcuWpcVslwAyJhNmKBXqC6fFTkCuaj7lYpLW7e1CW90gR9Q9pB
ZqNQSzEjIJwYIaTDkM+t1HMUPAEHZAhqvdLxNPkyK1phP3pugqIRQIQWh1DxPmSy
p8uACPxduJER7OnJEJ4suFKcK3tUOIhy4eY4dFEcpxSJ3UxonsDFQReijZ4BXBaS
xn9KscYjOJbnT7LltBmuYs2EwMtsM+YqJxPH8REC8bpF4yQVhyLzbIGeLcjafh0E
iowu159A+AajLetCtrv/UjV9EobqHJCIfJthsXMohP/OR8JZC/rxgSMDKIsh7yvd
+uvlWGbMAIU0yqf8mwpUFiao54GMKq9pdZXxB63dp+0FwFxxrlTknd3y8Q3Jm6pj
TqUDIGT0gDO/akG+uuSaRnh0qvQD9HHvyJVN9xNNNtIej96ahpI3PUqhr5Y1mpyn
If/lhexbsG19eqGLuVkYFFffjrE1FvuoMPHqtW5kr6G4rBbHhCZ+UDnmvvzknLzI
dwwhrMdbUX3Uvi9hA3Slbdb1qzN2w63RJ+38sMC4j8Pn7ogHwHzV7SknzHcj5sbZ
0MIObb4nGFShZaIN8ED5Nnuchh779+UKjQDumHucSwsWlN8lGV5ts9wPA9dv5E+8
eFGXVLT/cyfjABWKw8PMRcKTIg+xYowgvB6SkUFb9F6CaJ5PzgTI1zFgH3ikPOBB
aJCKw7j5fhJ+ELvLnxY4k7NXEiQdsgLPpHghl387SOb0fsDo8UGPnx6/b9FVVFy5
im99Mf+zwrsi9XbYWGL8lee06AswfnRTVLfR/v06jlZ0DHWq448M+d7hucUIH6jx
FauO1CPHvAc+8ZoP2V+uRJuZy9ZK8kYgoJR44GOdYAOo/YDlwZZlWIusd5zHmz8X
2BMbgwtOPgkttCvWQdloyG2EYNko9LPTRnZpPeTJNW/BLxS+kgezLk6CH8ATbZgP
Vo0l5Jkcdnwnle9OnTLpg28lMrelJK71aWJTDedd+oRXT93lo7uK1cO5CIMwhVpH
wjYe6uiGEg7JY9cw0xHzdCmuwzKUzegfvPrVpMZWkfivv4utaCLXO+zaWGMOy3R9
JXZN3OjBmxr8yfP1woEX7Uh51otKMhuI6AHovHFUfDPcDAblfVsqb1hWqNIiBJF0
RLtUG+9uAwKZMv/UTgxf9Z26uW7KBuR8ILPEetroc1ZQmRDIsr8lfP1eoH3un9vj
x2dSNxbPqtThGXQZFkFVO39N9qvwj1cEdsNGkDs4NX2HWR2Ry5KApwHOlW9sqj/C
/FvJtHYwz/X5nTChsQ0xENopVfJZ4u6xArksv5BYfT42ppL6CfzQqJiF316svlNP
ful2jVqkI7AmtPNh00+ZKjXtxZue0t57cUhtxIV+zu7hhwpd4JkJDINDRjKjqfkT
/Bvz8sHwAjX7ZhBeB0Ajr3MJrgSv44cgOHBdDeR330HGgrkvYwYOYby6xxblMyrk
IOKMbclUqysTiRetos1+ERf93b1SVdqgwglQbV9+Zj3MnDwhsRUFvyvpZ7i/V6pG
gUfebraSoMuPfOc/JWgbXPbYxk2nvSlZHW/pPiUz8onKgrYDcjp4UNDf/BAVO70a
39udFIE9Su+o6W5gVzqLRZT3lVaYyO7fWyOCWdQynYfTR9jnKW0ABOjPsMzz0ndX
CnpVONPpNDhxKSbeJefePEezagFaHpBT9AXiQS5e1toPsbJoJLYQ3mNAbVy+8tF8
qjobS4X/W8QCZF5rXE5nZ6dO5eVQcWY5PFTRjupNaa0eDDXbbX/Lep9ViP59Ryry
gEt2U65u3Cxpp62GUHQddXm5qWXUccdkN1YmPsPdpcttNrIrwac2DqXPLDKb1+8a
0g80L8yn/iQiTwpmgxtI3gnTsiWjr2ihY+3EsY1iHTWuc4uNavPVW3qI+DzNr5BT
cbhIUKd+pjrf6o2YlDW+aeYcVu1E3JdoZYIKDlHloagCYghe9VHhR+RpruWhZmxD
P0R+2tEHG4mi24p010i9/UPRqQstZWllRnfpqpbOcECa0C6NwKRv0feLD8vY0+y5
FUa7PzLGJzT1pCW5CZP1vdJx5i5r55niyzXu6wTjqSvuYoeBBnhGz5IT4NT/S8Zw
uRPnUNi4hvI4vLaDSwHO60pqyxH7cT8eGNsjlL54Fu2kljW+CK/LN5z0aU9Wrot4
PPUvXl7ZbM8RxNG/emlfBdQ8K9izP3qywPUwPorJAYIH0+epdYlovs8XowK/1Sc2
FEagRzejItvF6agxivxGi1O67yocbtf8mOt+7c1LkJY7Ryh0nAaIJlDL9/6ri3tW
6frVACVlP3oYurX0e9cJeUZj4CcrravkwtgfVsmrYw9QpGHt6xshdsi6h4NaNxz/
67s5SkViHovujerwENXrqoTQ/eZ+fG3zciq1nH0Pyqv0gv33ryE3q53kyoYiVomu
D7BLnMbJYqLuZSp9WX5IDEw9iN1WVTmVU1US1UIHWJnrLLfuuX5y3jzgawaU5GIG
vGO8+/AaXP67pKG0e7nW4Ntl5RGh6k9YNjkpauUthUeSpfiEm1WwrBwkhGd0TSkf
S+2Ds+N25b9cgvzfPuDWv34+3L1L238KlfvTCT0XtSC/lRblEmYn1PLpYInVUmgF
7N4gjcxDpItPmvdfXNRyQvzXXZWTaTSAZsTuMFhrES8ucPmuHFO5U+KbkWzqENxT
rC42Gc0zJqiQZ+dulKf05L8xaIkzCkmFB+9Ksg+gsYE8R06qlK9qJAU/WQQZTSMg
DT2t6CcjvBn+vV/DZq7FN5QA6ZV4M7IZL4vzV4JhnrmpKGUCQujFKnYDRWk/jwYH
kgth4R5Sk6BhNJ+8wbvo5ZxAgUxoaKGV32i2PqSm828HbZA1F3fRjnKBggn4PZ59
jHwM+ntccqbLQXG003Z+jbjPbb6+G13tP6h2OCJjWn4ORD1qsTWvWeCVz1qJmHIh
hiJrBnFoViGfOMjasBC3Lm4E+3PsHTFlnyEcJLFs9Wy3w+p2fNlzLsu0mgdgwSLo
gawnXwMt3bChohgC2w3bJNPspy81Ydmm8FmF02/uTB9CAx9zW+cXKTN3ueH2pm1b
ZbaalrrfzhvUbHwV/0FHucC9flUTrUYZNbGJbFyqzTVYTeO0P1oAirLuZOtdrlxx
H2ST1Dcr9NiKlPJyweW6UacgamEkjhxYmxg3yzr/PadhV9l53LqhAc6cUkli0duE
XNPvBMx98s9X5VlQPswk/qhAvyc/JnhYvi34i66jKTm1hjufgL5jAkI8ZrDTd5Sy
06JyJ/+6q/uVY4wMZ8USEGfp9ut6+LFhW5HdvGqxphDwu6hg2mhLWl8pla2forUn
aBBNQcqTGrZxJWs9jCTaFYi3Adm8Pn7isr8zKx05XifLwBV+IBCupveZdOKN06vn
tpOuDk/UXToDzXMMQX510jhvGMK7OKwAjaZxeUeBDp0zNWMYF174siUmcNDtCuSh
srUZ5jQ43H2eY2X4BTbXiFKjjj6SdVkIBOt6ysEwswGFiUdJy+VNmZzoXpWVlVzs
1T6GK5cokG3Kc4wgGdteLDRIpv8v5b1mSmeVr+/3HhMJ1ia1SJtP+shr5K3GvBRv
m8oFic8+VrVtEBDa2enYIHbkyAZhf+Xj26PavKKtd3pyzn38mwlEvjlE2CcI0fTx
gI/bxLEjI3/r0lvICNZvE2Qx0RH+K/cxNugQOeHbOBGI2t1GhVWl95Cuo5NGxwY5
Y7MJsMIDFXoNoNMCKPve66TuwaneeBXBOZ37eSy/ndcQiMxiwjxdBy6VE9mISPVD
R1VRCtv4wDnB8dlmTRsSFSSBEoEWiwADLgExD1Kf/UVnXMiBWHPXqDAlbmK/L9p3
y8GANsEvI1BSR8LTnS+2ybP/XQduWkwiths/h/Par32WiD6ZRxeSNa8EYDxxH7uX
R+mWt5ZPt1YjTipSVyurd9BOrSZ4/ukCoZsG+rNiGhSZQ39wJ8c5c2bZNqv4vmHZ
UZAkkHByz7nkpWfA1zV4qwHbe8dPGDzIIVdOnsSUPZOPKrc+UPQJ8FHcNJ2K83UY
gStcfaSDmBq62O9/t2nRq6f40rSTBnt//JxQ8P/qPGaT2eTmFoBTiWoKD8UpUV16
vPxBgKHt/2DVS/0oJfA2Zrqmzrh833qVP20hQUayr3FL/RfDoNp09dBZ4FDhgV9c
orkHiVkDZ0T8CYu4mpyvzBwt1UddZ1TdvfKifHLHta075b4+vszOlToQ+wq94vRo
oAosW7WFd5flM1QmOde6RH94lShKzj+A7w7nBQ6pbWRGFA+TjE235MOI6BaIcrRH
y07BM+v8hIDi39XA/G5YaNFq9e9WVLjt53EDGENF3gXei+QJWQu9yIrtd//275n7
8QeNjBq4v2A/0SrS4q9DRDLheRInC+CXSc0KkEOqKlOZ22j30oq8RGUnFREJnObC
OjbhZxGDKrXXpfCv0P7vL2XXB7bKTRsR/XDh9DokMbXcvb9Efq8F4BwESjqJHuwj
O3E6YMI/GMgLhQnLMkKz3i440r25bQSHmPK5QFFsJUaNr0MI+b2YsXidH6h5pVTt
OHhCAo1hlh8iPAG9d0tdSOnQ1Km7BsPziu4iB4k8OwFMPT5EpRc0stWIsI+rcKAB
JcSinAy2/xkR7y5zmwTQfysJpS6HUWkLnSy8eEJ9G9YETDWrHh9P9b0QuSSaC9qM
zvTzPSg5b8MAi2zsYgpNKKAikrAg9+hhDHse8Ep13BtV1bEA/flFZh55D9D/05gF
v8rVzzLVog7sqwoxZgA+TJ5zCk0ivMfUspZxCSbAISGCvcYrUguo/z3gaQ2soAAd
Y7Zd/Pnc/pN1NzPE7enGzL5X7v0tNHk8kk1tqvWo6xpuCe+Tur26iiOdSR+rPgZl
Yc4nKtkqQMBoUd5VeoklnAFDOFbYA5A7yrFzC3lWASKTSzu7qHEGcpTuwhg57yWM
iTw1279cWKFu/TMV6WGX0lThN7PtoeffGOfSJKrZZuQVdLjsr5/yh/9s8mZfeAyl
KeFnqSn62vUpylYzC8bYw2A2Jkcm8kqiEqDG8hAJz/MserquOA1s0Rbdv3HM9f8q
byLB1aI5+kGCbI/1jzdZuyi1gFOOkgNtU/HiJqkybDjm2AE1vSWWrsdyt+cG+5s1
gIMEg6InzGCuiH8Xqrc2CrryteOMKzemEIp5CGuzSYfvdevIBrajQFuk5IqfBUsh
90+mpEuc/nUcyWdhRN0rL4/5IOEZnBWqYVbrLijgrCJB/cYi74uxqXu3+MvvlhZ+
LyrrSAuOsLiYCouqYpePSb2sa0DdSnbFUHAZGvIn1+XsZA1C+XV9dZaOEDiJQ0KS
6c+UVM8u0wco578rxfKjOOBxVCKVnIf7Z8Wnt/ew27FZuH/ynE7FvXBkVaW0HN2o
ATeIMFyEv+yg1UGQifmyzniPTPaUmqmMaGJVcxinLB3XwYLFwR4FofLsMNPugbY4
1bmSdLYAdsmqRKe1mzksPP2BQTVlYH84z/2DahdQk+LTzd5fpwG9mGnaLOJmEv2b
Lzy88WELW/nBEb6xuFroU/VVrb0j99eL4gXKDHVYUXXRc7FMFAqxVyxZMKQxvPPl
a549ugqEmeeLK4OsSg4i0FoRo2CjmodxvDn5e4qCTFU3skqZnOexNd4AoPXC/CJD
ZvvlVrdvor079AD5b/1vttOH2ugNmuo5V45CfNSSTKgnr2dxfPgfEQZQWYxGZRLu
uCtGn0NWZccdg99TuRjwBArYt//PPx5T5P/6zj+6nU/x83JDUW3xzacZBXU0gUJe
WSGA7t/KDNHv79JBPhb5RRFQEJPGbYugujrSit4MnQU8h7TpBAKRdEXfaVVRjVPA
fnHpiFbCd4HBgU9MLvrOfsrZmYNtUUVT/dWaTaz4nJ5fQ3GwzBn8/57/f+Oqbn9F
u5KvoZi5bG1cDmVbfskproBgvjgZrrHD7yW5Ixqivqt7IexGGcUptuSDbT5p2u9b
3POcDXmQWDx6I68UCXaaJQxiVFyvIvIp1NZZo6xbPfQmWwyWhLZS4pUKDwTyHV3B
Szg0VIU+EzwpQX8Ooq50K58FRXms+esa6+ON6LzVMvEPGgAFz4nYthJ8vBqqh3kF
VIR1NP9W02y26E/6gUGPKRi1Xax4UHO4a2Xi7HUxsT5m2YwtDC40LMrOqixfzc02
9PeSTlttmSRFTNvf+IA7lveJOvG7/Erm9zFwuwQLXvb3+OSz1aCdzVY8yQvmbMnJ
xfPlAuqLFPiBOxfa69lBeord9ZvGR4I+d+U1bRfuO2S0I7Ekc1KXi8ydTCU+ur6b
p6VZsLjJ1dAAiCd4VRybFSjeleyWiXbkywfCM45rxHnHFpNHgjPlOis3bl0lotCq
6Dnl0AwnUUyQEdHsTuTxY6RiToC2YR/pd1aGd++Vhc5yS2BvjTl1tbIh4eDEDNBT
DIas6yvTMbW+PzKR106TK6YQxW1GWIg3uJrnPxfv3H+PXQ6sBoTPZWLEBlnyEBNl
eMGEzjDlVXdfMJlrs8kL1N8uGLKZ2oQqXrmh4wscwT6AUvac3Wh62+fkpm0Wg6Ms
DQiwr4mYTPIs9MHk/26X85dmXGy9LEEYPVo6x8ivAcwfn3B3JjvMKNAmVjWOflR9
YkOzn/i745kumcdO61lfQhF4YoHHuW53T9IOKiPf1a2RDyfvBCDNEZ4BpaV82QVZ
jLdHm+fLcYYSu0Asp7+qo+bx2d1XjQ/gcCOC6juObj5zAUID0xIY5urpmk1pyp69
IwkOQxQvtfTMTqTjRFxe0EpMGLBbvrtpwzVGsmYI5FP3BTcpx8yuWInv1s+kDnjN
LgGLmef2GBWWqNjwgPRtvM8pgErsJcYHQ7qsq0XCtj6R+EmkapiBhauyXsAb84oS
ARBZvYYJiirRro4RIaF8i0jG1HtjAod2nHB40m0RUfxwDL6cywzzJIIIlW7+8gYX
la8ljTRwJetVG9tzi104oLUxlwaMFpReSU9A88KLNaPYlpFeX1LbsdsupWV+iTlt
EpcT1UAXDFwZCYdyNZgHs5ATXMKkxQrKpKNcIR41fCt7IpqxkEH1jdkdsQavbN+E
pH0e6+C3JaxB7FrZO7LQbY/KNaUfooxC8X2Lwav5OoKPMCxD/prEBQDE4oWK5nzH
X1l/5pDXLgFVV8/DgxV857eXl2GpIXHFXvOmz5Oqc+yy4+wCjLyXOlchD5IztZVz
in6xVHKDfT0aLjhuu7gxacQ89k0vrRyVo71KkoxzkLnViixfySLnIroznuFucMNY
EcOEQN7yqbipobTPkJm5X48nvF+bB+PXuWznwBpNRx0A3bhRp162oiURz21PF135
0fXfaw6UUlhl6i5sWB2mJV533Cx3RvQkufwQya3ACPg0HeFLQ7edhEVNVuOD31wO
kP0ljdflHdDXZucnY9G6l/iAcy0jQrGD5i41LMMyapgWDvp9OFGS2S2xe5o9La47
XPuUtFj4sXRaVvePEzZ6Z8qpoOL50N8gGmXlnwT+wdYn2Bj+v/oPrcb2g7n5gptC
a5NmpBWeZItsQ1m2qEFXNdWFvLD9KP5tzIh4mQGhGA1jJwwktpzfPGlqqYxoRWhj
zzZ84oCbpOZ3dpZvM4CdMYRoU7N0fqqg97dBomc2Ot7wulcRgUq8wrBCcdLuOCrx
QcECFXXsKAPwIt2Bkb8VrvpCCRoXGLGcJwOcSc9lAIoJBsRB2KDSpzs9qaTaLi/n
poWFY2m9SM9O8p6AsGO6TqPKG/+d8ZIdhP3ZVaxMoaNl08F0Xi4dZkCNXzdy93Fd
sOG9kPYGxMy/eSeAVq3k68xIMCGVWWR3BWbdzKOqV/UIiGnBXnKCRbD3JUJb5A+y
8WOw0o9j4nT8HRb1WcdvWEwNiX0Odqgp6+cuSTy8zylgLX+SKUQbO70s3owk4b0H
7J0eK6XfXVRYrBC2CUlQPf7yHYDNiBFK//11EMEDcLOm5KfgP3bsLUxc2STJfbJz
P54UDgtQpW7W7gocGQM7DcircN1mMv0KFQ3kAIwVycKkmFCD6fqaNbZ5tQLVRFiq
uVPyL2dOFs7okvLv6Uhz3BphOOyywYBfJjk3sdheH/Tv/xtLWf4nf3Rl8TO5v1zH
Kc2ffm/BEsUYsvAdxuzw5aFe+UQJw2AkspAOFX3L5CQMH9+tUylnHRDbuB9ND9rh
bKkAD3kKPMa0PUd5orlQMMR2g7EHcQzOiv58jZ84nVVfnFDY1H+QuZg/izbyyp/b
T6IqqCpZKW5OmDNpY76PiMCaZgSP0nhNpxqPUEhP0TMEGUIAcq59HFL0/kB5zAkO
WeKwvSn3enHRYZenrc9niq5/P/TkQS6McfQ9BrJQUJil5LCUJnqiOEFmYx1Tdf0P
6SHnBZb3nz6JG4MSMZ4lFnnmBvzPiCZufD5C/uH8YsqApPHTbKNwmGrgGmiApt/8
I98+vI8/L2xnd0VRLnmPseZQcerATPrrSN5qeTAPMPCcav1UTZtr+vQmgNk4hdJV
byRCnNgwFpt1f67Cez+5I8cSJjnj5zda+IE2jJCJ3q+7GVpFuDu6FOP1D9J+jzXp
beUsMHYQJ2KKaK6KcWjkCeSvHSBueGsHQfbYPSUMykldNlA/tBRWdhOQzLi3yhIW
ETuUmgWEDDjHgoTFfD8GwDbczcDT54UPRhfwswmNIooHbV1Mxq0FCjr/BUA7X4RO
M2y5cZgM9HAWtHRVg0jm6Jn4s/tmL2uYvaZPKJjrHaUN+wBg+u8hWGMbj9q3J5BE
8gxk07YBBSOcz2nq1pd9mnaxYHznFflgDL91GO3ZUqTNRfIoIZH9XGQfcw8NPZvJ
VCXH9lenGObbU5JDS6p0bfx5EuZR6h/Sl41zbI7mS7MwslxbXIvaLpJpwb4VTBCX
6paSlweWX3UtJ3WRQgNwNamalsBOdZCfYISYzSPQCZrdgiD8mqDrRh8qnbWdxB0R
fG4xjVAC5yNxrhzVASAMdZVrYBoBol7PJ5k49SbsgA9CVzK2EKOep/IWG4c09L0s
lVAzES74aVvdbqQqd2rcNVH+tfBfOe9N7lLcCPerhiodAuJDUeQd3SmC4Ramopvw
nbrKSRm+Fe85jNt/j9FA0L5vsFJ5BvHAHF2cNizaC7FZrH1PKLZBwU0t0c3M6Vgm
ZIgEjut8qoEhZYhBC23Y5N1TRDNd3biletqDqmsI6pQ337pv2IFNhDmuPCuvjrSV
AVZsSG1ceo+7GBxaXvnD2evEA6ILpbuKCrupaXi3rbCwD1HnOj7CKKiyxQvEhIfa
bPzPWn3XFes7XAoZJZ4fHLT1ZNqn4AFBORKzSEuf1bRs5HwIOa8g9uJiANqQ2syF
cNIYJmIcMjwaNWgj3JWdnuR7yHWPC/AT5lCmPeEHvCstEkZ5JZ4AcBt+46GHdA0m
IBJsQgEStiGNG3u6X/LiCx2z4OdXTC73MTIAinNxI1OE1l58qnfjWqoFFMHQqnv3
ngSmp9fOiPpgA14an/jlnMHp+E06eVrz2Ax+t27wNg9z7WSvzJtfvT4KkCljlhX6
SHGx9TgQYSwcQ1tk2oqatAsjXB6SUOmQG+aVhZwsjPr6HMBxd0O+qTl1hvsENjCe
Gb90HMITRxcto91BCaHSaG0L9tyUupelZa5zYAOd/kwYy5IEEZnnfAPO07nHHzXR
NEcS+RM2WkMWlbyfTd8W3PxwEXiuXjGpOpG7ZPcre/AOb+SIYninjO178/LO9CsK
evsb9wc+Z8BpRKyjrqXOWPMk+VK74mwDV3kp15GTbnxcmPt/Nc8koPAKC15Fwt8F
opeCdoA83AG/tM7St8sO/zD0L9b6DokrjvhVw3neIlDl2WvUa7luT6hXGNqj6PL9
vxv+g1j4B3XSUjt9fdM4DVe7VbrMYTQkvfbZSUfzuZLUuBT2WhYUoqFkyRdRQbxr
2Cez2TV2y36bKeJ9zTEZLrut6xeBicaDdIcNyUrpEz2EbeicECwCweyfYwsJqg9P
DYwnrdI91ZNnlZEXQ4yrEfmfuOLA7qwVpQms0xoTzUfa1+VzNIB43MzBQY9c3kmp
s4bIfoAfAtQzW1BKny0KqbrXKddvem5uFY12KyY06EQ705FzSZrVnJC4H8/bIm2B
6SLcuOGJbvr5i0D5Z4v8tR3GuLpL1GozGTVbdqjY3m6RSJQn/sqbNWWcdQ6FE7nB
r72D31E2SgT8lznGp/cDCGhFs/HIUGjRd+nFGMuO28QbZIzLhHZxP1kGuesUZDAS
o7AFhCiMTtKrNbot8g7QCIcdn71AsbXz/v0gLIlUFNHucvq+ABJpLtYf2v01mz5G
2zI9kh5TTE+q7Q/qo2cnbbZudJU64mpkDg7n9XzzWFxglT/QQdScXftS50dEBQYp
9f16+M/X8fvH4TCIsUI+KfSKIkGt6GLmTU2cRoOJNvuXCYhi/GgtPEuo+knFkxS9
6sUX2Ctx+8EEU6jg318fHNLuC8XaEd76iHQRNg/GTMavASjOi/Iw4Mpt1p66hSVe
PzjKNPwNaoN9wT9cgZeoQInSBakwV8/1yTIFXdV21Ig/OHFqXVrNN1TZZ1Ke7iL+
gg+lLbOzNSYBoKK+d3DXza7DaqWfvepiNM+7eG+qzgbbFIVKJbDuAmS0FGpPhuP/
OUWNYOg4avLuVFvVVSD1dCnAumTB/rJPJ99CnNa11r3fJKIq52VT4hnrYBlHjV8c
KGOl+VuxuOLIgVWpVf/ANkfceCmNxJ7ybNDvwGsGdO6da90WrAjModzhzK45H4Qj
aMbBhyXW+TYhdMEPKPfANvxgW4PPZ5/944iH196fkPhWdk16JBbCQOjjDx+m4Lmd
wKM2VWS8qf/MSDZWKT0JqbA5yaDjTPHAxGs7Q1UN4NS3bulG82qdUy6SleQdyac8
VDkdmPWuqX0F+vavt4UL4B0xLw7Zer0R41I1I20ZIEocgX+wHXacCOIKCKVQFW1L
x91yAvwx/1llAIIu5FKCEQTFfGyXJv02jvCCzkYsQVHpU67YXY+RNlEHKvPwvzRm
6+fC+GXLefa3KQWNnwSTyT2n1wwTRfl8pwMQ5IK9W8LGWThD7m/eosG9JUGPESyM
bGsrKj5xrYHd7y77PbmNV0SwPzuCd1wrS2X88eEPilkaYTOgp79S/WzSTmCVCgAC
89NVz9h6PFcl32a/y2vXV0Y3LzRVUVvTBieDeXqXrfDlymJILX5PG5Hd+Tkm/RBq
XJ8VWmiox2jmjkWBeVVLGhZRrdpBySbZAKPP3myosMxZeuYFxIEEDQKZ+4I1D/GU
5TxPgP+lwyIajr2XXX0qAzdcDmk8rnU1atTCiYbsfl2NLAQfET0dvkpipt3uV902
0wc9o1muHdbTKb9fyGKXtJ60PZHRk6M4Fe8yDPt8A1nFfO5cQTG9xLbbAjLJXBAt
G0KtIs3aEhyfoQAur/kqm0YrKH3Xis3xGOa8N+d5XCJ6XeO4JckH2v1+Ca6uTa7E
tH6rBy/MBHsO8NamZPZ0PblzBj+hY7304bVnwZIBdZfV3tIUZRrFKIkNBbYOJTnS
vWfZDUKCAlyq991RdbX3IzL0iSxV7duFLhgJnWe7M7mVamtXuSfi6kE6hdvYVDDj
Fy53JHVR6GnciOfYA9lRfk7Igzvgok5hiDCBYm96vqt0cmoAhuB0uPBM2sUxrIoP
RpOLml8HjOr7qFJmkiD3jxo3PP4+IZy8Rat6LdrgpOaKeeilptKz062zqyX3edFX
ILfpanjD9xBldYC/mhY4hiLMtGlaCnM9vGY1TdmVL89ZCdjFSkxx/MVpLe1ODWcK
zEXqQfnXk+yNj2UsS25jpmiuUg8T21sASxwLm162CiKZkcERDSgACjfyOfxcQw6K
8x4cNg0/58vuvGLOMT3P4nFtVCUjuyMIjuMNpcboMO+ippRofioTTGLwJ3RdukPB
5kZ6vXWFUHbNND8VjJNaNi9wEU3Z5Af/PKm64NwnaDQ6xvwY8EwegqP7C5JGxPMc
KaMvqizkecJJZrMDtUx9lNG2s3Wgp4V/q483C2JfyzH5ZDCxLTggH8HOJxhNKz43
sS2zVZQq7D4vPkOXmKYbpguV7VaJTMm6RS0+JuGPI55xXUy49IjBEaAyPitOHRaw
Vz0vTKRnwaaAOZXkZ7iF0+rL6IXMb7I5vQ+BTlyvpgHkvMwY6qN6lla0Jg3or9Rk
ykIDgriBJQvhVLb6fbuJV3UyrlR8cR5houNQMoTZja0AHXZ3eZ8WrgmqnqsZLC8e
XCQe0MvPtnsaRqyX0hGHp2JcZsY/mmnJ10l7ZwJj9QYYjgQBbZyPuCh75ME3K6S0
YQtFtmAB6wmPBqBwndyzX5vfKpRJW1PL8FeVPvBYx5/rRegQdo6WeXlsCjrihnsW
Sf6IRs+OMJ0L5S3YXZ4cCcA1zOhIuSRyroKN1zcIyDflXbNhvOvGfH8MLP9PbVdR
c1yG+0M/pt/nInk4bt8jEY5P3Z1EFCxMO6xuDlGQxMYxHfhc4uMDs2sAiRYSBco9
HWfpe4YJoCnYwbZPeLSw2dhAxEdbrC/H4XTNoFMXo5K3tAoUDGImlSb2u+RhnQ2f
5yeYCXT9EiJv1CToW3qAeaurT7tcC+LIfPjAyyIFhyA50U74uOy5HDXS94B++PNg
MqV2WACmk64auJ4qmwKTHHobrsb0d6XzL/wGgoy6mq5FNufAR0JK6qUXqFhoRHvs
zyeYmLIJMBXn8EiVdzfneLfN0f16dEt0T1kvCb/ua3ESK58kliECcU1e2tgTo6pg
9GDA2JuD6Ap/vrQMyfBo8XuPZKhpAdnniCTwVUAHf+5jWrUcf8wOTXdWD9b5fWRW
C5CVf3Boarr5WCxOQparSdyn+fnfbvOz4r+6WpNSZC6qUQ00WdT1MYNg/RApRf9B
wMIrjC+vy+S/2rkTSICAfJAv6VDqHmzqt7TH9XYeUgAbYF8kg5Yu7yKbQDl6jEd9
`protect end_protected