`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6272 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmWdo24EC1SLhDeUV9o12ewQ
ulXp2xSZ5P2RSggIKJUy/fb5NMnNt7XXpoSdQ33FnbLzkSJ+E0Yhh9EbsPBePL44
K+Za7YHZlGRiqJnSFTxcObwoiFMrri7BdYu4u9E6b423kevV3agtdvYmDIkejuY+
1eTKbpoF+/kgOlJqsqKLNDkMWbefsEZURXKgsoIexa1gdDJArewFBEW/y8dTcUeA
o9MfUVncSUmBj88Tb0vbO6vFCyklXskJ0ifO2bZ6A3FF/FBgwSGxjg2cLMSGEHfk
bVGOgACk9Ow4z99ADal28kqqiyoCjkrNqrfs5YKGcKGlgHJWwPGdv/U4mHYOxhsc
05GhC3jS8LExiGP6EiBBZRHwW2LY6kkoyoUZtG5HFkuxPpd9WdDwCPA2OKrnEC1q
qGtq7/qryKI6oYy/HjMm9iKYe1U/udVv0GT3caTdpBHd8OZ2JXkc4iTEB/qPOqrY
LCNFXrp/FIJ9djcyK7cDQDIurXy1kihmGrcGdIsIpJ8z9k8XxSMbf0pbQJydZ9U4
FLI7iX90ttbhTscjG27gCZJpHPGRCliFhpf4mbfVBaONC/LGW3TwLe4hizusRedQ
zWlThh8rlH4B81g7d7tz8pon2f94u2DkdgXeH1Z06AWJ8G7jDf7OYTRrn0plKtyC
LjSrfLtLkrumnTbOofGNI6EelsI7/6eTAaI0PH83pTkQMiDBWaYUz083c8INcyuX
E0s7YiR/AGYB8Sx8mLvDyiwKZM6BqRgMD2ZslKSYFn/glFJOIOtYSzg5HDMrMZT/
Ie6fqQSVxEvi0zhUxnvLTYQmylSK7nqp7b45P24YYnaSqSc58RBhN3lv8hRl5wDn
IX2VyQW+5BL2mNqLM+2mMzqm9qzaI0t/1ikjqNmVIygOBjRfvVz+IAMnS/Ya4jyh
LGnDhdYul3kTjcJW+ESxC1IzStUgiTyWiz2EJMy36dsFkmm2H0nORog48zJyGojS
k/4FcqLRtJFovEiSwoLwiUyNfrk6q25VIORjds/TzA8MbyckVXFh4O2KV3lPI/Ym
xADVVvMSkBc+197TRn94PVCOs6k1zBAnI4zyO2Ft3X154Bb+i4lwYjYsxyY4/HJh
U4+1wpeW3VwsZ7/QONCUviu5znLpDP4wWjK1oXTnnAN714RjwmHJ0nmvX0rITtRI
+K6U9F2ED8vbs09xW9cfFig1d2uLqX8eo3m5ySVfh1ALeyxaDeDmJnKetnzDfW6/
MLslnrLC60rZlGHEwB5nb6B1Bz3yVwvfYCTmgUsw5+C/FtrhP4DtZjO5ALEcHbyo
nXja5T0cdQ0TTwO+XG542kJEK36C7t7elJIszePW//tcu1E569Zo3qZ+oUHDwf23
8E9B8oxYZd/KP93S8vGauDjmwlF9XyM4pzTRG9J67Eep/9r2rrmmWTyUVJWi8AlJ
qrUrQyjz1SG2AhIFStIRLE0NHbhEEJSXTOYxUWjWYOsv83FZNhrHFaVRwnC0q/ky
luilMvSI0DzZNrl/5wtGsZsDjzXbfz254sGCBcvKcXhClSSs+g6/fIUW0Rj+4Iyo
Rm1LFSUZNXMoQqzmHkiL3Q0Brv2jseyP5u0uf5aGuhHBXNmzyLmHOQNkeZbz/g8o
bNwZvXLYhr6VulgHvTufh5YAUfrxrclAWIyJh3yzfJ4rCVMjtFBeqn+a/BxjjBB1
hCB1herTqLL9n7m+1oDG0dgs/Iv182EJifYqxt9xLqM9bKSRw0O2Pok6ZkU/l83b
hk7wYKyYsO9WcF+KIvv203Zrzr+o5A9GXYSM0wtNIDhTauhvZjxsaUz5/3q0o5X1
1WDjWr254fmf1UIKkCWrZx8GJ0YrsVgLwLB+dT7IEpez/vs3F9Zc4gZJRd8+W6lu
FIBtpj6iZWSF+4LDTV2B7jaXtvTiTYUWfgI9EguRWHSREJdUeS1sZetrqBHxPOkC
XtsGu4KqM9UQOzZhh7QPdmTAGgHqu/RloClFUpG+7YUvfDvSUboVFMEe3puMaoPz
ogTdYRAb8Vxbw+KzNF12A2zkVznlsmHAjo0s3dK77R3PUSTSDjuhufAOO9kMNegi
tOSTQhkapXtxo1pp+aD+BTeXk2uR5Qask9VDm7SG+mx+7GtM4lu95XtQ2uxERy9V
hW/TIIkRASGPq0sAQy4Rb2fDDGOMDoW8PdoSOftWU9KvI0O/z31ztcjRUZgordIe
g+sCyIFUnKs5IbQVbNzBRCV+BEwJOYihoZxy3OfY0j8h5BXE/L7s9batCLIDR+AZ
g2toyHzhBicQ6N8mohpGpyMLCaFGKhdTcGDsJa+lCFckjTbHJpv+HU0Cvx8iHMy6
6QNvBMseKOsxtooEKvoXOVmXh8uLvWpCnZjl0dQ/Tqw1nHt8uSfj5RS3mJ2l2JG2
soXt9oJtxTCmrwITOdHHz9uMAnc3fpob+S2ndqDRoBL1e+ASdr2mEgDvV+8MJ+FB
8vqgcTBdvvKTC6Qg5HuEvfvCEvSEjZtvtai00LOGGHG+uOq1NbMAfIugQwHlrmEl
pb0cMhvbAphS+A23f3dAVxoPj7Dvwz2s5HQFSDswv6dWsg6ETx1TGTFepEQF/434
88UH3IKUa5Z+CclBVBGLTmcdzVvXv2BCGm/V3iQjIRM5SxLIKz1YgLKzGGJhJ1oS
7rUmXs1/wninDGQtteXaUAMhJ5h1jMQGT8dWx/9WBF8tnPth/PROWilsK6GUa6qq
VRAPabHcdFS9QDcm8EvZg1OQjFDewFvNdteL7mbx9XyHMDnZ/fcOWTQZhcTA71G6
TwNu+TZthAUZMUTJ+Hbxry3Do+OMAYev6wIQO6HVn26i8QF6L2zgakMdaXnh227Y
Am571o9wRNlnRuCOFFisVS/RP1u5VgzWFKWmlghpkfiKo3FneawYTaXoFqLoCWix
/aeNfH0sc9r4qr/5XsgOmgUmhmpTN+sszacH0ffECHrcaz4Weish3kz3M3uMn7ga
tWztGMX3HfZdVHXa8SWi2vAWoFXUB0x3rLp8W7dn5LTvcOz9RCUge6PfLyCoq3p8
agd7sk7RlEb+sHso8KtPOxgYg8D6TNafrTPP4EyKwQiiefbSbTCxQUpzh75t2kHO
wUzS7irMelLDbdBxhPPDWDEKSY9WrQnf53ZTDZRAQPw/7Ub5IXaokEmR4XgxEH0m
54rUMKVa1HWLkRR9N0WQHgF4MHdyf90nMIoKHE1XGX8eixaWdQQc/q1xyDxKUTzi
SI9iBtKo1WNW8N9ptc++p2ZNFAyTQS89xiSYIFXtfuvHb4Dbtff2FXbeCJ7shqlu
xcrCEUxvRQlDf0455QP7qhLG6crTf2j/JMKXHtyVuIXalvrJSy0Ykz/PBz91uSph
cPrgp6KlFyabUwtiScI2nDMtJMhhTz2d6AtYSHXMeJXIVJ8rWUknA893CC4Dse6m
lYztWyi8n+y3Y2WNHEe+aF19ku7SBvD+88kmKH3XomPRFk3w+zLhPOqZCoVZrpKC
NQizu/hw1cIHDL+RVLIMcuRbXiJLgcNYqUDoa166+1wNI1EHtxz0RMBvT0jaasr6
En25Ey/GK2e2eVfdjIPVCfkPXyqz8xTlIYpPZR3u9H0humboxxQmML2O2RKEKdX0
Ws2EOwcU0YWfGAa32ymwxHzIjSLSGjsvL/u1ujTtEU390FM7E4jRYGusjgEO7OTy
jY/VAwtBmK1Nt4WWAwN1YGg6kyjejVZopipksqlTsThiwlwoD6nZ6gxFCLMRxrWq
k55LkZ9HNwqLdf97RJfSsD5j2vnc5ccXDHrYQAvQzxAZFBv/2zY1089QZbbzmkxk
KUMG5++LaMHjtp/0mzFQR3GVTQ8Bjcceghzc4D8ygCEdEwkOMBE9xibrQUvWDVJ0
9zeCp2VDxig7TOJdCOEfp0jjy0rNi0GasULH9Cv4RIwBvEAc7ksyZYUwljgqvV+X
flW2Osg0QKNqyZQN6OzFpWoCxZuWT15d09V7JSJArPX/rqSqt4eB5r+dJhvtRa7f
vszc0EfnKlOUYiiPIwoDFj9suWR2M/d8uTuEBVp6DtCDe70TmZf5ML8BtuJk9QRO
hpC/Lrtj8c8XPIQ5PwOB754KhOz33gbTybn+HIbgbb0Na1qaAbW5qTD0/Hrsnd65
dU4u26DHGqUk9YDpWUNVWXWClSgdb2OY49rgdmFlyUr/Ti7+si2gTLJ9EdG0HoYC
Gh1uUKBtEasMsh1tQMpuokZxsi/Jw6tCh/Kegr21qW8IuDxFAVd6xzb+yl2eB2KW
RqxHxxrGbpYGrW7N5TqKRr+3nN3UZhh+oeMoT2eh1TtQXcZRGm09Gp6jUKCEH+UC
jAtbFYHinnkz74JYjFnNlYiJdzXm/SliDpaMfGShxkVbAPNrSUt++8p5r3eRT+Cc
XUQK4TfSygcvewDVkkq4qlE6GkTZYGhaVRH1xnCuc3H3HdTuXqI06o46Yt15qe01
GLyvHLvz4KJtWDQC8Y64DnznHczFXsTbz7UpudjlWTnSeE+qIrCkqkxqKyahZYBy
vpeBsFAqv5d76TfeZHOedSdQu6LvDp8b43DFlJnvVJhDx5vHOL7dHYCai3bIcV31
VhQeHuDxSkEtI6MHGN9tK0IxJOgf6JJrt1f2HgXOT6ptMGKS0edm+I84w4Kn8JK4
HKW8/8EQSMelW+TqRPLvYMXat4e2sK7X1kMBC47C0oEtg7Ce7WPVis5gDRQmJ37D
glQss7ak+grJ6Xib9VUNcyxL0gOXSre/MWLGqIMgPpDuWyK+eDg4+TurVAQzW8Gh
v23FhaibxzAeBx3ZwBOQUPnF55R3yOikKIu3i+p4u5jky+ihGF9hmx2LSpz+ah9G
DeXXLAO1/SkA2NB8lmEG8aJOQ2AaNLN1PoOrj8tXAFU9WlajgN5qqIc4PF6b3FEK
+k2jDTM+GtUeOl68spskfsrPDe8xutJl1bw6YcwPkW5LmvoY0x41LkDVNi6jkjSJ
G5cfzrXTYmsDkBbH9TN4urfzOapPv/XpL642kASAidf/gPnSc+1i29GFYfJaEE5p
92hN1xZkrvXHMAj43Z9Ov0i0/Fw/6IWiCJkzSH/A1xsnPKoCsViaKZJF2abh5G0H
YXiI5anLgoqBxYxgHbTuXKMaG3CV/tNELIQS2WNefCoCEpaRWQpLDzvR9XBHBVRV
788bSb2+1UCugt6YLaImiV9ngHfhnmuQ/l/1HJeMC0+FXFY0t9U1t5OYocJYVdyU
K5P2LVy9CXz3Ro36bDFzpTGrajVgJZqjfNrrBMFsGakPTnJ1252uCWz1NE0FKxKX
HOizKwQWMHKXVJ6JYC8weQcf5ckCALHSUt/9UoaLOVJUMcTWw3PIFmSmiSpozIZU
acg1tM0cSl3ynMURcJpPkgaL7HksmRCb9xRh6/fOrgAlWPiX/BQa7hOotQ85VzGL
VOuEW7bQcHjQ/S8xM9+QnC4H7I1nEYio9sINs6fmjl7SO4/uIVam0Rn1NkbJshiY
zChlWPjhTB0YzgUfzNjTevH388mSPk1iBxVz0jO5ZTYqWNFajqAwBXgO6YHOTpmb
MrGoWMswhCd7eEOfByQt5+Vnv1dcQBwwvWn6Jec/Au/Sd1kcotMm+qXN1BzzOnKu
SZH9EfPwxkJ75lFc0Ss6FXohI7w/O50pvDhAvMyxwNcw8DoLcR21rSgFy1HhgQUg
3GLBvaiNJtAleEghegWrfU7rlpUir1yZIzCjihZsIqvSNNjNwZ34369tu1gBeEo6
54M5fLayHHAEf37/paQEQLT6SQGrF97z8sHyvmeCZAZSrqSNJeajLvyb8RRg4Sjy
JFe7cvDRWjTFP9AurX+e+N38OvIZwqMVY+ppY2UnBfoQu3vkwoyJrFAJAY90xifb
bZRzxV8iBIe/eD2jK0JGGYIFgNnWk6O8hB8BgFwkQbXp5xmPJo4BY3DUxPPD+bMi
L9zqCaTyUFR7UYGRDd2xf1nh5vU7iqzDNjan1WTbKioMYepxueVzVzX7EJU87y6p
4HQ0RLaulBzs4xqOQ19wE4cYgqQpdAtaxGonKz6VgVAQwrTIhPDsQVh25rGva7gq
iAI3KI6+64zS82LeQTNpscJk6F2WDHQAJvCNfur7yKCI68/I99UkEhnOneMrskbK
0H2oJM9qbiqzCDRuRLv0dQzVvLdOOX7ef9DC66ADmUdFXK9oriszPfQIaeWP8yE4
mz/aO2j43iOr8nuyUoNly3gcY2+TgL4vQCrGxFr7G6Swb9ZANDoE7XW3r2y2CSZo
1fUQY478IjMXBCj/Xtukx943f62pkGKpbxUmx4GUzNb2xQGuOdNbQngI+F3Pxh9r
yWLEJ5s2yjkkQZF7Fph8vmfvt/5bvUnymFByvSRg1WAQ+KatUZ+0sZgTUKcCs2ZY
El9R6ypbW2haZAyU4vteRw7n5Ia5Kjix8swtDP2mVHUiXg/p/FMnGST1XvzAt+xo
M80WKpA3+6oNBbPo5YfA7Wm3PjclueDtdH2Hg1fO4ZcfyknpBqeJDw1B0J0bey/R
KflScyK7bDaj8+WNgManrHLWF4f9Du0tzb4Yid0VcLod5Ps/E6zJ5tXuiaP6u3RD
aw0Y3lAMockrJJfrNWoCbKVZzGSEiuzznTmwJDh2s/m7hiidPdkqqtCBMlGEVAS2
VPF+E6KLU10uzAIkPOsLSKyoi7gGKnkZWxz35tJN280JbMivdjENU5cEDU1kqfD2
BUHdX8U+pnkqr0WdA5P39KBkgJ7qwy8TRTV315mxzmDO6ekUb3kKv1JYQhOUKcos
/g6eeB31ZvBBz0LpDCxfNSGAg+PKAi+rD9a2xG+gE0yFCk/kF24OCNP2myBDe9qt
QpDbrngXe6TTzCeSpEUfShks0GfJeHyyKKyCj2Vj60Z26t5R98I4bcncGAbsU+Iy
V0xwB/TjlRh3F/j+QEROrZijjNRmPz7+tjhGm89hAAAoefkd3WDSPxoZ/RhSp4/k
XQGQQPRQQbOkwbqoxNhAfqb/lu1FW0nw/gSjR4X5XngZthcLm2OfFiLIPTcqCZV9
580vcil4c/4HK9WV/WybKr0w4pS6fKyLaXKL82SAOm0Sp4Mn63FtzMAxF/nBZHyc
BH61NChfwPv+Wa85PIdJvKC5DidMyOBtydJQMWBE+DNRsqEE6PaTCvs6vhvb3CHm
yPAzcwzDbxikuzRDNZ1/rfhKIg5gSogmvI+3Foiq8rOIneFNyRBIbXK/bhTzcIFO
Xnc4UtnYaUm1nwayIO5LdaCx50wZ6Xtk28tdxx9H7WvbVj1M5t2LgvHoOt1n9ghH
IkCiKO3o49SweHJaaUwjJH7KRGoxt8Tv324cPcnGuI5htEWuwbB71w6aU9zDy5Bg
8Q+cbjNMpwT7h1ORcXzKsAWLshk27Yo5hQg3lDY5iw4M4lgNgv2ZufuHbzt9NN/R
RZLAR9le6DwCndXuhQhWIadsCeKi/Id403RJzDHRaGiY95exdHBpEpYK0Bj8g7hn
VSYblMMFKwM3xv7rhRYu1mYJ/a4/3qslEYsPIamve4sq1bppeBFqGNl9MoSg3GlF
onwvWCehCkQ9nQj90w1yKVhzMr+LBzRB+tjsVTTlHwcMaW+A1md7DFEZPHgzQODF
4fPyIpy1DLQtvd/F05Cc9LZ55ggDQxSMAlyNG+F9Od8Yd9YMX3Ft/Cbo4F5N64AD
y+NZ6aJF1p9b8nXUuHJpn/0HQwhx0rb7Hu1nwgsVQAOzcUdjrNO5myU6ryY4iTnc
XCXtQ1ZMrL3ne5nqpQjK5kTdbRS2SxdwVlT2POzuWO50KtH9JZhPWKiJiOzIBp71
XCqcUFmBZoxbIFHJO771bcRMDndUTto0YPyyFRKeDQjlTaHG/B55OfPBy1QsmTnS
0HatFnxPXKGYrqVE1F/KxonSEvJnJgbfV8+R5TtIw+F7xa83UQPWp+7soiWOIh/R
gAL4LPVshEldt8u1NeBGnJo1AOo47o6X1ftDkkZ+hS/bQT8xaYyuVwnVHZU9fgmn
VBTgH+LSo1JQNOM+vw1NsGqjM2EdXQ1VemGAVjun51FhaGpJqStoGSu2dDspmJhU
gCSqA1XhJEMnm6UluXvtGl3wRu7Mn4V/dp2m7W+89e7Nrl3gr84sp/1IVen0T7v2
etUaW3p6cnDBSOk6ZDfXdt9IHi9OwkdQitidKCdSyyh8W1cX3SNltUNZPGsT6He6
kuEUgl4svw0lCnXIKH5Y4tkYow8SU3V6hrmGYWt69ScwN93/RDqWNp05ge88b9ek
61rgTAGmENpcuKBwuOAYilZWam8zTJTOb2CTwHk2AoY=
`protect end_protected