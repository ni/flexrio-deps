`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2048 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
K21MooLiMCXVPibvGUiGAZYWqqRtfKjPj37SgMdgGfmCFJtiMYOCGEJAPc9xJ/p+
uf9aao9P+By4yu9wcHju7RBxymtRF4xuFhlKGYFJjWnn0avml0oT0GhSu2o5h12u
W1d8YyKKE3g4U3iLzdHIYR5j7GTGpx88CiVx926Obwh0HjxO0gtzuA+fFEyry/da
VuA0h1Rn2Dk65NWdHBQwjrpWLk7R1ozsaXTzxTIN3ZNWmiQ4Xo99q1/uH3sB2Cur
RWcKNKQxlyeGQ2IMc7LBYnVWVdQJJjIsqwMQQGzXu1BJ1ufpEpP6TRFuHGqaP9j1
q84p4mwjl483IKrBiJIE75U3o+d5kg3cRr6/77ly5tgjiqVJcSb68axbe3YkikgG
wInwxDUy8qUSwJ6H9FAkFHFT1VlpjH5XM40a2cTAaKARz0CH1Jdrp0yrwpH0/mcY
XyDW9/0JypnFDmvyTMQV+QrN843e0FuHcDZ/5lafcmxqORxbSswU781NdTh1nWed
i6mgrU99hfxI0qN0to8AzrCfFg66WDOAKe7t225VDMLqViB21mpahgKfvgZDMNHt
vtPVxuAqMIovDSJmHBbJ4TVlZLlorWmdH0sWHdE/iT2degKnYNzBXmW2tawcmiKP
T9/1FtVq+EgGtbQ3W9xEl9KFD7yTSsip2fVsHBrT5McxiKUD9zXvG/sdAz7gQMHj
KCnlh6VfGp4C4ho443WsbSBsbrSRlFzhZIKQWmIwXLFWVMxlbir8ckgiVR+2N8ne
hyXRosNMnsMA32rX5YDyPQvASs7yyFy3v5riL4AemZorXKyNMbaqK/EzT0VQrs6M
pa7nDDtejiGxBOvEWWFiNcmEbTGoopG0FNIHymc+B8HQt7HQFwpHPIiJBaadoj23
VNd3xqcUFj2QKlRY0hq6vUcKF17KohMnuD7+Ec8b+q4VT3mmiBAEFbh8FTRUMeIO
orcnA+/OVYPjbScceOMYi//cwanhYVF109mGtKaWsiGbijQSU0IzWKudt1DHc5Js
v3SEOdHXgiStJ4Bm/0UJpS95E2zyLD/XaZu07J6FBC/RpxbNTb6P1TU5uPZkpxzC
0oS7yCuv74u0ECmrwrFzCokmPMYrd8Tsfwr7VCZS0tomgPMSOIWCrgOYaGz1Djai
upqJW8hkOTOKldzTLHn0cK2nEUXb6HhU8gmoDJpYq044f3480sDJ4iEr+DiuceON
T1kntjW4nOPVMcJVSmw50JBpM/mp6b6dt6pQTwYje6O64qsCLABMuBgZmHE/J36I
+ca+Myp7M+aFKreTJMpjkGTiPQyxMvCS2vEUN/XkiYHcjPE13UXAC7wMyLjx6Tkn
qISNpWgIjwTqi1yMy0gYG4ArzHNK/lZTbv55lY38na2cPK/0emixP0OgAAhV3T3v
5wuzj9Vwnc/xQ6fhzoA7q6qnZcR8JAUKYQUYcvU8x52buCKmI6akb/wm+hyzEUhf
DZjCrIr0Xi+xhNcPmOPzaEZMj1aFuG1X8FSIgp639irDBmaaVG5nkkwvbKN8XIzi
nZKcZRZYT1ptlW97tDMcE/Vv4qegN3S+9T0jXFlHaca+A1c4SD54LtiN+y9JBsBr
A7P6eROdWRSYU+LlLVHLvNwWoKmV3lGfqsPO84m8uO4zBAeAQUHSzM6TbwxH4/L6
92cBNUZXnmF+INGmA0kUPWhK1V2v8va43YB5g/uJIJL6F9+a6QABYuJ0phBfSqxz
xLx3G8dAi6i096KMSXFSzMvYYA5TpCde6WjtXpdDeMlAl7O6Uw77qmjexSawfAWf
MZVsTQ+dcvaZjg4VTQQZvJmIckxKQD4Ci0ka5N8KlID2h4XZxhWC+vKFF9lnVs6S
tt9yzwd5PK/MqdS9RRB3UHXDUarmp/xcWmb4fX6pLDpQc3CfeEfRiRmasQfTzXwp
0ysowStrFD1WnBLPxZBZp8lG366yH2G4wiHBc8X7Ff8luzMLbzOFGjcLnP5/axx8
uBWpyIHsnzhMfXdQ+E5qQ/XEkTw+sDQNZ+SOE9ikfWatAEzNiuDiXVf256KaYu1o
Nw4hvKRqbtU+NugxieFMJ0FwY39KT4zxnVeUkznZJ2yzb6B3HHxrVFSKVS6WGn0/
UoswPPH90ZqncDK3WzF91AjEi7ij6kT1OTfr46OEhrDjVYq8QJRBUc8+dMtLn8Oa
zjTLI2Gh01aQ/xY1JCh7C+cd6pmN64j2OsaNbSMaKcwuZJWP+HfLfG00oCA3p9MY
Rgsg6mlB4OKx/DLxyOhDBrzVg7iberR9hIbc4Xbsd7wgNP0cZVczOw7zy/iMoAJb
o7cxjRTvhZb8q6IOXKq5fdfuYF2HrLCPQ5DP65EIXiwCXQMpsW8f0zyYBMlFaaDL
BB3kGJuLxxU9GwWS03i0nUImgbbbPAC3XVovJFnfUduwUnjOR+Bo7RUMCxi1cdRA
qw2UKLwo4TIHSLZKn+vIbgKQ5riSaSYOUJpv05d87/+oj6EQ82qwI6UxH2mrcDS+
ouIjDWNh1VV35XIc4vQNQ5EYH0zkYXhySR+dXGocbgyEQeTxHQ4Ux3yMRk2wDJHW
EtzF7uKLLrWq9Tz0u+0B7/FqZ/uRn3HqldivCeAPKZM=
`protect end_protected