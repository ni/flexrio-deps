`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11328 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nn7oC/bbltaB6y9f4wbJdgh
0G6WvBg4Flfb54G2gjKn2yCDQNQwxZwi/Rt8/TbFUO7/UmwdvMAQdzyqbiXDYS4a
JHDZ/1E3CPRHjWSjdotJCPBSco1UbApC4cgI292qfHR/R+yC2nbXJjQKZ/DOHqSX
iHj15iEU+YPVkf2q0ZgMsWnJb6wGxYXhbqDdKtyEwV+mLg06j8OlwoxvPoyq7Aeo
dmrE8adGMzx1xKIoS9VJIaOIhe8w29b/qra/scVd1q45mTCEG/wk6qvWVaXHnOXB
stbLO8+HCv4XH1qZERcozMRlcYqE29ubtCfoeKLDq2E/OFRUJXT9dnasAlcXD+iE
BxVsgWmjEyGGePjPPF7mD0X+atiw9vXKJygVeeRyPj0s6ojtAYSrYuNqmSwEijL0
xSZFMZsEjROI0zeaCPnyNr1Dkcc2OZnvhEKOh1EVzqwQyi1C5MWzwDFwsL7lCKYA
0lF4Gq7qJ2H69GfutRQBZX+pk1Odpaufpn8d3fKyxs8ONkaHNTLjYpt78mouVp6L
JAnNeshwY/Ucj7opM49Zc3kOyPw9pMCMGA1MohQ3xkuLz/PL7X2lUWRrUgsOUFRO
ZKbXIJygxkVFNguREmOLAOvAnYCgNZ3ibxiYeLLRY8Ed6+rBW4GQ7vP6h5z0JJm2
cJYD3DNbms4XH0qfRUY014EkuGAcrUD+92R1DvBCaTnRnwUKWa8MOC/McNyAcbOs
5qmfWpn7DEmMBZYsDeueKkTNTGRBdjtJ2iIZreIzpB//LzSYnTR9KnmYntkHJeNb
9TJxI5LKzsu2CkZtAdhsSt2r/JVkjRnhTL31rhBSai5aF0Xw1guHe9c9exThYuhd
dvkLRhgd+1j41qwj7rNs7DgOxBTzZaXU+8qiq8riRe/Uo8dNJShfI0NWyJ7H4qiI
GRNgFN6Sq1QZne2loUZKcsRc/3RBD/1cf30Vo5EmrcKu309Czq1le2bY2Iqtfe2r
cdmNl90Sq3y3M+/zsIO/h9MImOR7VJP0DhAsL3ZMU9aXNSIhv+elHh+NcYHBnDE3
j/LxImZbi6xyytwoLsmQAL0WCA6sOVVBCHPZVUurZzR7+QA2lkbGYtUspsAMsKtl
14KI2Nu4OpB2fEcmUW4xbEZaWiJ5WkPYaMTJGbDzrPyXx/PfIB4FCfqz1vg4WSCs
ePlyh0TWvu1LzRMu2hDpC0ux5h14FJMsNOo/klXOAg2qBfaLMSvlZhX6CZPGIrmi
Vn/8igXb8zIoVceiprW2hOUhO5ce2DwlQ4A6jCcYeGjwHIKL3wfdMD491fkLXLbY
TG1BK51Fc5a5pQ8CwNm8POotdbtxR7nvMYK8Edo08Yt7X8U4YNLhds1dZAU0JjXZ
l/JxeldauvzNuou312X9aryUNrGdzaV3q7Bj04vEGkMy6gerJKV3KhO2fT+T2K7m
WcFMAIJofeXLHIXk9iwwPEq2BdymCn8tDl9Qi/ihNqdmlGqYWLBQEESDD6kiGOen
g26RnBa23Wd29iLwz5ikgJ7frCGZ0xYpx/rtSS9GN2Um/Sh5yHuvJJioSGvZyS13
5y0kjUhayDEfDbxczPW74o5KqJ36Wr3s0selAw+Rwu26T+UUwM14ZWWO3+teK1YS
4UPM1vDcJoIAYjAZ17SX7RZj0Ru+RuYFUqIw3IU7Hl5eUrQP0JyPk9HaujQSQP3L
snLeubeaJPSOeBP977dWmvlEsw/HxB5VARpFyz7etVu3bhjQKc57goQostHeKuQ4
A+cLOMv3rdw2OqO0x7syknuuIGA+HbusYPfqUXK1PHn1sWjrHiiOU/hqUOEjkkb2
WsGrdqTRqc5W7y84URLSla0PExaoeMoz6URTy3C5ZpykMULOiu/aqFwrVDIyzdYI
hWEGl9xao1CoqGRhzcnF4I7QXFHsV4YJERlZ5XC4HvlEL+H9anPdBGVuFAiTm6bQ
xYYZzEwlt7QtOrjeeQVB4z7598jDyJY4e0pbiVHYWSbC1gl9H7si2OR0EC/Af9FZ
KwSbOjtYYq3uKTqNYOlOnWyk0GFyUS8WfnWfFCbeZW5GDgAYOFxjlo8OZ7hzfNFG
vdkmQhYq85kXKRBudu0XExoAbzgttIPjpgb/V1uUO0Zy6uWUU+DX5Uq2VAc81q5w
zxyUVEIAfNGhdnL+mezdlsHUEUe7M7OxX9+F7NsKzjPUamEmqFGDza6kIDzhQEV/
6AyiRw716/u0bD9XVbOYGlGvTqfl1Oth+S36zJUrEkh1p6diWz8jMo6g7bVQz9LM
KxNpHx5EI42fNboiumU2WNKvDNBpxT1ZovpH9bQKio9CBms6MayML3yKAdZiEZvI
9vQ1rOIQPhpMdR0Wqt7O5pWaX/4DI/M1/BYRGwlepJSfeKy5VL0mg1VPm19sXrM1
3o5cQQXh7r4E8OMuexzhzeThJvng4q0MiyDMfY+QTJ4ZjAN30FyRWi4wiM8XC96Z
9QXTVVXNUALyrsX4YkzTrASmFHW5G4Pd2CoXMEgU7zQi86yN+14+s4BSxrjXLv53
6ZWslXFkG69hy1pXNXwM/ep6PtvW8hKxF8vx+gvtusfSbOPqnrpL7isHvQRheU//
WfRqHOZWe8lfXIT0WP+7SWT0t45csvJId9JHdMRnM2XLLdnLAhFYWz1HUw1+Xt+y
lNedG8MqtbjuhsVE9I0v0PdzBin20500wm6yVl4oS+MgWy9pt9zFcs0gu9xD+0iM
cFd+Q07idPxA5jnOtZsYjWM0oqw5pOygkCtlKdAs64AvDGQHz5yHEaY+j00e7+ng
tBRUb2GVN/iOJlwtD8lQz9BURp53YlwY6pKMd9x+4y7kkwCd824AhMbyh5y/GZqs
O73D2+OlokfgxRg5JnEOYCs2UV42HM7CHWHPxr2UeZ7C5jSvTgtRKH/NDo3rsmoe
jAbI788o1PDOZR+uQ4Vw6oIiQ0u8t3W0HgZSO0hpTJBhf8gjjN5uj8PYauadr/sd
PrYHzDKZ0rAQ+q+6+ejGP9xoCzfOr51MOeFuEqAcnre5e460REP0j4c3+wV2qndp
xchMJrsUFThf4B8B5Dv1uFKnTU0l1JfxYnMTn0lGOyBHoujy0VJeeLEzz/G5ogB0
RK/565UJiqqoZPWbiNjSDFB10tN1dLHciAQy2XZjg3h5RrDrWnoX5/WkDkJ0sqHj
VDFj+JadmtJPpZyIWC17FTI5r72MMj+v1yjN/lEx0ABFeRjnJz4cZbAeKV7+gBzV
FnRnUZzwNAKssYClPd9BBbsBhTGKD5wfZG/v6hjYNNlWVS90jHm61p0YbG9iUz3i
gIWgVNyHeQv63Ad0ahJLnG4NatcMrhq99Nt4PrUUqAI6VRjCT+Oa7LysrJENGtcw
Pue8egc/67aBF3nP7GERIJxuJOe/j1wv1rm4zXgDyqLoGYIBZ3twcsf6lFJ+IjCA
1Z/NZM6V4fqETp4HNYViKiI3OYM02WAnhNDeMrEmQSV2gSc/anYcn8OcUyZboLlX
MbawukpOkf8BcaMN0f59p70R/MjSU/P5+N+O0GKa7GMk7ucYFVx5Nl3AlVGEg1kx
/Ajj5lDofisOXoWm2IjAc7/D2oEcotqMSVTGU/3/o6a+6J8IghRuDjRahQmOlJus
B5J9PJNBmPpYoIrDgvYndnYDf6PC7dQCRrk9NXwJK4lbyTx+NRLdT6w1WrfzPM2k
8L7RcTsFxShx2atDPuqktOR696UUvIFpjEqbavWCaWuZp0+zv/B9Bz1HxcNOgznz
AYi0vE5M/Yh36hOrsFcg0/Qm2hZkuRrikxWZGJKcCbkVectF1xaGYrC09HgcFem1
zLrmGEKI3zzJF6MAa2gK3L++101qO10nRaR5ryyFaFc9M9oli50Bxa7umZhxOkrg
H3Bx8CRXU1LeN29ecsH0zNHRCugALpJv8dRLRV5zzww08iybdJ6Rg4NoNOz1SdG2
0fDKdXMG33HNZeOYP1eW9+hKUX9JEv8K0STE58K7ppuGM4PdLg9WVKR3YwhPycpu
TYdt+8uVIibeW+h+0vl/FIf6aG0kdlmJhF5sCYY+WInWbYCzQCAXdZ/jN/zBmYCC
NgKKO10aT8p2Itvw0ET7pDyiLMNqT1uLq/OH2bc7pOa1wjbWG0kqlxICJMK99ult
UiE3CRI5P81TF1uuAjQmPnF21JYbds3Vu3YwZf/mW7sHvNvha0cBM20FNRZWIWSV
ByjMF2TU1R6Fv9TaUoUYTACXGx0AaS432F3jkrlpo5ffrcUPLTUHwNI6yA+PK/IW
PKDxeKq7+b9S2HJPLXVkm9Mbik96gq+5GaSIChmvZXaXeakVMCZwWuOfdDf9o0wY
4qTDf65l9HY6nPJeSDW+xgFZ04ZnaauPqvgIdAxBbqrIOZi/nxJ+YOxPFAXfp4+u
38naixtDnrEukT3b3iSz2QViqd/2HFREppC3NY6L59ks3SJFKjJsds69a3lu8Vsc
wNjRI6kSjS5YlVJWCpHjH50r5YDnkOCq+uUnAhkm5IW3I5po/Rrk+xjHbxkxHR/V
z95x4ROzQ32zrqAB4ikwu7JlPId2Egejdaqw7iHLLMLe2vLbsDzal4lBuJK7JvgP
ggp4d3wWj6xqMlNP6AeJllJoWDl8jzmsEl4eE3WNdvBqzz8x7q3sML8hgV8VL0EC
JFmiacmgjqUaW8w7J7ZfkQW7/PrhVmoHxSiADBcza7MxC9PebNbzJ9pAoyJu30T8
ylNKE2jQuJSxj+1CyxHqjpiQbTARbdTWlIvrRn1lZCl4reka0AwyQUpEpI2z9guV
OFH6Jf0mAUjGyGlxwiKYcfb+BvmPZyKl1ogbA3VikjmdanjQ7wzcYJDZOJUOCJNP
JSANYfyVVptBMF3YlIX6bpzl43nqsRsU3Fahjflv1XYFWYBCD7vdSmdAU3hQoO3u
FnA61pInrwy4MHRwC3qOG/DhHyYD76Zn9yKD/WeSHJh+xcH2YN2xGDkjMhtUpofY
Mih9SP/R+QtnIJGqVRQkJuF2mVADJae2+HUuPqJuKEK61wGexyJtuFTkcXF0ic6j
pPx2OpV9wW9YnItLThOyqCeTvztCl4ooEvgpBjjA65MCD+z2/ayHe1v69WMY8GI4
MGTM50UuYz2n5uNzH6/M7P+9OeWlcS6Yar1KrzeGo4Z1234xffamWGLPjcONTCPF
IPlAF7SOLXxVq6YZkbKOL11HGyosNWE28SkOrbh8dJ/U0Wb90FaYcROTLxhCk592
5tFnEhnFxIlXYKsdCvwFrpUc4ozk2OyEaMxLaNUMEBUvdGcG+1tJXSX9FOC4pZ+H
/IhC5JVSOCns9dduqYJBtR+lzSQR4xSQSpR6WiR0oY6ymSlmQa6e2ekGNNgvRHdT
DxQSUE4c5VwRaWYyWH4GODqSUdgyL6PLu3JT+IRHko7+H3WEp7rGRZ1bPVNIX7lH
VPbWANGkjAgbf1P1LP5Yj8DKF1FWXMuGLKe5Y6Y2thvZQPTSiG3wBVvEfB5h50/7
Map+tBZfQqntmJKINXP7t3zJPyqe67++nbjXLMLxGyFno/JGS3t6z4Y3MO1M4mVK
ejEwBgbSsq5uMe97Z3LWDzGphV7SZJrvXBg51sJbLXA97Ag9RPfNqG9TgJPfbbG2
n1P5vd2AU3T7srbb6vU+8I4m0Pm9s5X95JGTPEjcr61uqQ4LIvrwFBoBQPono0C9
OWoGflasXbsTfxmmUSe9xFD+2mnZzp9/znVyxPNSWnI6ijhWDG5+rhm35KuLKP3W
tJXN7DiOTRlISBRNj0oKbwdgLJ+7KdDTZQPaye/pApMGIm03R1EQJghu5TYuRS4W
oV6sHSphWfW4uDXBXU9gnRnI92QjEnqnFiyIUQ/B/nnIsBVzFqJoSc9qJDKUv6Of
AFKpSAnQqFk4T8k/7RwuF50CJ6yt2aR5kFQjrVe1vaxQWjq1rt7Ep7a5GzdB/xfD
sMhTRUvYNB8UisOz6rNaJYh94hSS0vw+18aq988nCS3o7T9kNK62MNrWXry44kyG
NeMl3/po+9xSVOk5cgYlJk1DmYEnNk/0aHZ3AE5UN4aOizuVGf6WBin3UwmfnHSQ
2D8Tdb5VogmHHUnOQck39MhFy1nsGTIOLLtIz18G1HIllp/BKmgJzlG9Yz/Fo9LU
KSdLO1ynMQ3muz1dKJeAnbNJr9q2UdSURRk0CrbEJ/LQv8xW6bQSmsi1rMVgrZ1w
9USl4VSlfU2EoLwBvb2VFm3catIRM2B01J26B1ppAe9g/mtN+8NEbEJorKY/kzdf
m0FjwIshevBw0i8abnVtBokbEd35SV2GJG8HP7ywwBGtfL8R2bERSNJWqlcsGxR8
FkhoNFmjutCEfwBhjkVpN37aaW2jlheljy95mGgB0z40B3nC50WI+KVFnQXozGzA
7TrMb9DqaIYAYmu9Hz9AA9QA+8SC/NX/tMVmYN+IqFtD/+DGwNvBoCZIlb83PwM5
FRhBbR50H1lBpUT9fP84lLJBkGSFxtvOwZbrOeyc5rcZIfjiJvmxm7uCTjSRoeUI
VLpGIYDESy2w86mNqk8vAyzWKbsN6DDsyuc9r6cLT755XRPoYODVnfRrhrH+wE4Q
BEDOSrAGSsy4YZsE/g5zWmMu/4JCLcY+SMrdVYOamTOJuXzJRTFuVG5VIQdnLDcy
jUPD4CZuPNuhgEpHwA6n/GSwvynj1Mj2Abs+/ZQx1Mj2sOCXZBv4VsHRAtZZwcwd
TpPgo1kEl6uqAqb2oXWEBz4Pf63ItpoJK/t9c7g59YxLeh3tY6aL59/V2ru80dGS
hix81kgTv92mNcp/lpvshTIspKK7odCa+2Z0LJE6mbGJYz7UOjcQoEZhl592gj+9
/md670FxZJCZkcspn/nvqpiN5a9OraUYANCdN8mzUKObeOVwFuL88wVhGV/OITDC
nmsVdf22Yq4L0s4YhpIB5OHC79qbx6KTroysI+aKRQHLKI2ixYh1yRbIM1cMW5v4
TglpHNT8H2QuHpGmBUuBS1KQksWt5U7vxFCih++dBJintX1n0nxjrLKCdDCcdS6y
Mlz60ZH/hXG4m1jHKCmNTH5p+1xjiow1aCdEzGs5B0UDC91XMfZQ0sx7gNunG+e8
TQSsq7IxxgCnsmLsKHaGV5v7KaGj5SHUvrz3UsPt9b8VngJcpFqHPxyHFBBFfLt4
SdV0vsVqhwbesNpcZvP0tpAeA9xweHi6RK7oy4Ar9l+/APqfn8MDAi89a7zqkw3I
IdKCR5xVhukvMczRPtFCccRCFzsVKPOd+mN1AMaVxkrzdblW5iOsGcBQkeApwSsA
ejKdngLglD05ggpzwhY/0d1YTRxo4PW6l+y4As8XolbBxO44n2mJP7eUSmFyo/PQ
KpRYSUdipIvaB322pL9yUAeDHKW3viEBZfXP2iFrS7lVk0zDOJ/5ZykSesK2hacf
GUAChzKB/+BFI7v4KL0hAkUV0vogLEpjV5qOc4EorLLpjd/+Q5H4A/4evAxl1F3a
Rl8cNbFpbmTcAZY4TcGq4PpJXnLXkyXeARXUUy5AwlG1ZwDCwsBxbA/otLOMqalX
gGxbc4eyGszftb+BpJCkHBLPLdiSBuK0q/kzMJy0XaT9/147FrBEXYEaAshzZDfN
ij7DOAkbroRXhSdOEpN5/AycFYUtNb3b3dPGilgIO3aNqnundIkHZBJoeC9S1icH
ixPuGWdzEf3P7F6JzAHFPb26Q9bxEOpz3R7jIiz5659ksV9Q5D8uqcFfu3fnHsh/
RjBrRBlZVEKRncs8Mc9mCcAvw1WMiAr8eRjN824mQTmvXivt+66DMzjFEP+Uacw2
tQiXPx9Bc36L0Q8pWEvc07qMy75zvcp5t3Gmuooqbkz52XabvBLm3hI4L9NyNcxE
8kOvzHNhUBFpQH3QE2uuxhy3Qe/yiloHdMd/aXb2eMh5iPID6oOguCdmBrofShw0
r39mWTkNlQRJXidRY4tZhmlPp3R5a+hZlt+RHv06ErYxrpWxKakjcOihudHfLMmQ
1qMxoYkqzj0KHgMRKV+QoZttX542ySu7QLHfwZ61Vnq3zU5j4yogqkVonjOP0TOG
BhF/1bNdUKT+ZPNabvZNcJSnUClibGznKrXpkjloQYNvJowwt2tEOBDo6qyBtr8Z
M0Y1KH+uwGjaWzogG5Qbl/HUtyJk5RBuGutHT3yZ9TWKMKFU2LurGXqA9V0T8v6V
ZMn0k3M5cmHgjBysaNJtbreE7WuvHgurj83LOHh7KrgdrLu4NIDOy2dber4L7yej
yD1cr7OCQp9EHFc7TBywGxbot6wCovYzMuu8ngrknDEJ+JiKIORCJhXGMxdj3RgQ
rcUNVKxqBQ0HNjzAuRTTgP/7gLDAN+jtpHo4mDiY9+fIibIaCVnFK3lBRhAXWWne
boQFBc01wmsmia+FCT+SXI2Iw0BGmhT6A0L/h1sWacIJqmFsQoi+IgNcX3UW4vV4
d+8YogBLdx6VZIuapuNNVJCqF0CTjwDEbq0zH9I413Q5OkEFE1bdasuroCPod2eh
G5TaonFWmzplOOQ1KzzS/LDujp75BN4MG3PzzIqqM7/mME6az7y3mtfEnSjquxQo
Uwo1mQyNdMy/PADW/j1VxV11ehjizQa6X2wSbPgRG+Ge+t7NqmMbTC5/qR3S1/Sn
sqjQY3fqPbN7THt4owaG3Ws1Z9AT/y7dbVfWB2vLcozW9+c4kTRrM2DR4a4T/V7V
aMTfTSJjKrMslntkfI2FH/JhNGGnnaBxshMaVCXETaCSZ6WKj/FfdHGcWGymYUXt
h0mJQgUYvJBQZLpwZxqs1nVFsF4UnwMnIQXTCFRW7MHJ5cc1ZEFKV1Q26wxVRAy8
drAtvn6ZE7r0ndSOHKtwOXdXa9F3cpkqZKSSVGVD4VzihWrITdxtJtYzz0j3PYSX
qq9Aa3VUuA+9pKklLKhX2u+PPfqh9A7uo22oTl8Tg9x4hS+S1jq5QT2yZRNIA2vd
tAnhkJQ05DlXCqnhYaJRZmblMiGr0lF23Rdce1WdZNlUlQgERKg8YxqcLJjaw9nq
dkBA2mn05YaNK1COH/ACfLnNeZHF3VXS5Gv5oEWeuvpiHRqLBUKkCCFKBdNHowrf
EKrsLT+3Q7pFzhCrfmgPlhDef+avEWWt7VtC6S7Lp3yNkSzIvTkgabu1KUpTibAd
jyyL/H4nQLH9twnMhwvuSyGMxZSeze6iy10CiAsBVHcj/w2wnYGxbx8aJVsChnY5
OGZkfnrowB6eWmlWOzp6l/PeDbzbVGgsXKEz6mU8tt2ZCb9wWzW3uRtNccY9nFuH
8hV8HfhqW9k3gPp6AbHfkKySfECW5H4M6Qd0RIKPKQL4pmdllLQ0rDcbaw5k0jl7
yA4WoWNF36o28hfrnRFaC1+y7moHZgwNrV5Qdni/a400de59N/FpBuKLg9hn0tDa
4djEHA9jD5lRomRoUXp8S718nBlDqi/EhyUxZTTUdhcLYohf8AQuveIhwyvF99V4
Ddr1DGO9SYxGHUCrDf0eUvmUvIuGFRfrg5HtoXl9iomYYa9xYrTHxVEs+ki1BJcK
R/D8l8N8PDhfT7ni3BWgPEKUiABTwqJJtXmq9TJc3EgDKIBrOH0B1Unn5Ds0k/6X
7dxy2LavywVvB+cBYfRxI54wXocfyQOdhVKEMxSW0wfqbbX48BWPJm3OSRVwYlAj
IRLpc5rrInFaaBF+eQbYy5Dpoi6lUzDJ14tvIefTQILW6UA8Jj7CRR62fM6Smah8
l3tmI6i8GEwYElWReiZqZWR7Ygu+k5VGZCMJVpneVl5IXiDVM/L6Q7kmkNOKFu/P
Vyg6/qfG38wkiuGC2FVws59v1Sr39RhT/ZMckq0nRXTxjlRAniHhQA/ds4clr/LM
63PiR2h5KAJdzKHr3/WBnBNQ+0tedB5KHcHhhPIMfIzrhNTNMPppWIO7II/uW/Js
Gq5zeWLoOfOMl6RyQTlSXerO0PHTKiErS1TpuKQ0thBfmJnBd/5R+05B9Pk4R/sV
CotsmqpdOv3OJ2GoNcARSxz8LMbCwtsPJ+sy/t54mL9NuR1ZDhomRWlwYJR7H64l
0k2bbjexFn7eSJ2oiLhcPG9KApe3ciEdTijpp3cTHLt4uGtUXMHyERlP+ixsaBgn
58umLPoLcLmy1aNh4zk3pxNABNJfzAZRr2hFZD+vXERXr0xLHJ4mTI+qRcFNpmOc
ijk2Sy74s1f9oAmpR3mYto4uoD30EpEKHiL7EAneB/bGJV9lcVdhIoDYz6p5LYbZ
u/uAp0lJF+e8qw3ToUjxWf2VMz9YcQY9UQ4amEEnXJjYVovH9TW7X2oXNlDSmC1e
aqEgtP/qT5/6R1gtdQub+hZBYyjEU8MFkQjizQsh02i4SMVEjhoKPyV1Ai5V+atM
jnoFvPm+yMTrZFw+ABPZHw8cF4KQrBUSlQnwTiYKmcyopgTqPzkYzcMgorYzGswK
FJSxnncxyDQloLLetrRbdulQLCstWARxreJ/3vNG57UBkClC1Y5K5xKo0hFCdF6d
gDdSi8a00K1gSPgTlsEqQ5V3iOuAW5RPZOwgk0dMSlsblxc5grY0x5VsG/G0tguq
vxIvEc5f1IlN3pCQvTYrziO/k1eshaOsQHXHDfXfYHnK867g2m126hj3SIxMI2eU
pDEX1lcfWtAfSXT0T75Yh/3ml7LMrHEusNAcwfEiD8qHcuSKJudImt79ItkV7Uz5
xtJIvFxa6ch3XQurv6qi/ZNGjF8EvCmllJk1wOIjCwcudVeaz0yb8UDNql4y20G2
Yx83Bf2wkqqTPbd/NBc8y/KPrgEifOwa45V1Sk/Z7K54T9fQ5H8FMfyv6aauIXh5
5Cr+dZ9fK7gOq1o+3l1hPogeY1U4P0UXCs8LtFw4Hu92XjufT7B3kg2P6eIzGKrC
fnkUJJwvmYGwKY16NiJP3agvH35v0BemMz8bUbSmxrzD/6XIFTZoVklqZjKSYqbm
VTjUHcX89hkxA9bXeBmo8CIS0LJrO11ocC9TQ6UYTGm5iSHM94xoasX8S8qC9lAp
hZw+MB0zAbkdga1ZE34SA+6lPvB+GQ0UuQE80KPr/fK5RGzBEPAHQ+MZ5OryCMVQ
znVXnfEHH3smXje0Lga8CiN7DIkaYuuR5wN8AwCGHxw+qMUIG4wFpXwTRUQtaOLk
eMigcJyJ+/5ub2sJLVwQt17Rcfn9q4kJOuJ9pjG9Vc9RfM0nGx8SiZSMm+rk4mWl
d7D9myZHTGvdBipN9ond9BUzJUSRq9JDtW09WjUDk9jbQAPIK2wHqS2eKMZVj3HY
zT5BZHu77g5xiMX1+tpql37s7oHtFRwpnNhKCvKceUQO7iE1gOf8UtnsoJA6Qvqo
qZ97dierzIo//J/3uHWNldjcAckUcuzosErlNbTe4VJ2TWY0ttkc1yb9/tDQtD8c
eiQnPFYhHHpBtM6d7MeTU7KUv1MsouzYXqlr7VLWzQO7owcTp04w4ftAzYGeEV7m
KGitg0Vcym9TYGpRSXhN2u+WlsCQcWKATcfJqOPpR3/V/wMrRn7k/u2n+ckGnQO8
qG7ZwmFC9hOQTK2SAxCChVNTM6ILvLGJGr9uEx0F4Zlv5hmU39PgW6CkQ0LuIx/D
gEPfzy73FDly/w+dsOyItnSyJF6CchjxXgETYzazyBa1T2ZqV8bJTFqY8nxhVU6A
ea7L/Kd7zTxwpgnVV9bQXRPJ0snj/cFNpAdJrzPkW1SIG9tyg3nM/sBWJ6F5QCqd
ntUtQ+rsPUr8GLCuIu6NzMXon3dYs/OkV8FflikHsQnyXCGcd68rlUhoti1tiA6s
G7cnLlFjFS6hlow/OupRPGy58Yl39aHa0ypGhq1fZplQ4d3OjqDOgIXznDQthbN4
TI45j6EeNa6e1yS1D6sxDakJWulqedYdSP9/QXth/C+vgQ0VmQcyEwFqnXSNSq51
TL0H9gbPE6NHBsTCOz/TjOjj8uIDWIIMnvg5prn0WjUnh5vSGn0xsBGFk6EBFde3
ueXxdFWEVUD3N8LfC2O2wpbBL9cGDmKfu1Dzf8YoakdZyc6mmc5pTfYRlFfZgSKC
H537JfdassQFdJCpRLGblI/PV18vR/L4PbwZ1tz2O4PzRLhiHYHFX1rHBEeFU0Wk
TCMlmMm3qn25J18kkJ0CEJXm80YD4ilwD801aYN8ps1UL8nnIYvckGgUT585ahW0
bq9RQJjz0sit4jBNP938tNVAtwKFkTV/uaceVr9FdtxAOOXV1HSi+2Op9/ReLopb
l3nnWXoXwRejKdY59VoHQLnWATxuLb5VRBEbkY1SQkRmQSPSo1qUFoNL1T5H/MEo
QVpW41nR39sd3kjd0/xS+fvFgKbgWqRV610KU2Xot2klS2m2FD8A8iwjEBBfNiKw
8U3vY5qjosXusUma+Gdwpv8fN02p3H7srGcZal0DyAP4ulgoPzqlc2gl24kvS+ir
voaby5+lNsNZ+QPWnlJPAJweNS3PjPL33Bp1uTjS2dflq2m0VrltflNY66UIb9sx
0i8dVZ2E2KYeTxy4lY2+Bs4bCsMZwpY4bQNJAjCwTfxGQ7FtDEQ5JU6yz9mOiNec
kUUrB7wjKEqtzSGyP/Qh4X3lzvzu3PJlEyhQpE9YQRy+9OuQ1fWHCyZAgD5e1czB
fyj+Q1cUfJwvmeAPqj2B5CqCc+04jvtcihSga8j2gtDt1X4Tr8cizqD/tyXsbEyy
/gA6PGwYhMMIIo08kx0IYOe6CHigOngDG4ZtF/40dwUO8MALOfzwX4+U270YVHZl
0aqTv6K4SmIU2p1cJ4DFRWZ8VgL3nt8t/Nshcg6gpjoFZYoFD3PkyXcj4qZDIapV
uw0NhjAcI3o6FVFJ9UZvZo60UE3QnjRzp13a2n2FLaeIx0Dl2qiPttyyccgEyA7O
NTaJ8jm1nsIWOGuZ2uI2edOuIEBr2Mwtf/NQPNhUbmL/Evp0O0eLB2Q+QiJhT+j5
dXpRJG9+wadqEO0XHzZ6NZEmtGk6L91T2LLobwKV9SMl/Di3L6WeyG2HhrG2tOmS
GLyR9ytDT1jN+95qExSdSe+wJQ5ba/VLAj5g/VLasTQI9Hu8olmkEVv0h50G0nEN
CgF00XJ6RF0d8JSm5imI2avSEsidrV1G6+aq4lG7l4ksXGIN3Fo4JL6gpcCy7yF6
+lKKJF83rCl5bXUEZaEq5AMXoWw/xEi4Yplk/Qhyx88GanIOaHiyGabJU3FkeT3u
hPpVZZiVGANq6pWwa9iYtF8U+nEZjGlf4HwNy5hYLCJ4PtJACP2oesOx+Y7K2pbC
qprbPkszHInqzQUkbrG/C8QMXGpRiy4J8RY9bOS+k7Orcrff/gPywns2JpL3Qozb
Qh0/jJ5cADWpnRxZSdedPMxWFDUCTbmoNWWWuC621oioJKjGS/0k8mSyMNihAL2C
vEgimgjNxN8CRTBMwG1dQthvcBlgp8opx/3TUtcMS+4MDLnMARoMXEQUsJqFRYLb
Hrd6T1zAZf+NaAnS13ac3CEJFp5m26Djrmrgg63cqDoQo+LaM0ztD2SLRcAE/B8V
oJXAVZxld30POCM9KDx9VLr4HHNBq1KgMI65tEyrr1atGj2JdUQn9ASMVpYOCuBv
STlPf7wj9tuGalK02yTtVGYsiSEKV2VToD0kvkyCpmE8bEGD2Ph+syzbxT0Y8B9L
5ct1NUO8/22b3k+CFeDp5+PjOGOdZnpcSmTF9Ns3XnLRHzOch99u0GJjPMr7rT0s
rV9VeWaIrXySc6Y4tKVj0OKzvHbub23ehzrxtVzZSWdhJtI9krVbMrfNJ9DWATHl
rXWiQ1S9j1pc/T8UWS6JPC5V2BoitDzSo9W8NLPn3CBl3Je3HtmhtYTVf5WspYf+
DOQ2UWF9zYFMORTomisy+RM7i8SoGcUiUjEUW5YVZlmUf8MWWKHC6KsETrHn4/X6
PvRjUMR1Bsrp/rrGQhXzi3jZAFlqZQAY5U6K9lz5kv7PrNgQC3ptOMirbz0jqIUF
8fdhCVMW6vRoMBcCcDOvBDItElYOhn2WIPxbBf66NkPF5BxaqmJmnzV+jvdFBy50
OE9FFEkZA46L34CZb91PBhButPfvlNg2Hb0IDIHDwmEEGzN11JFlLq0ePSmqRlTX
A6CzyDPEiEdXSLpk5PlnMwSkxgShGJtnqA3dd6NwjPBuIZ0Q49H/trLKsGIDxS+U
5QoA7Eok8Jr9b0i01MlxLjYLY7FIM7QZlZ10FcpnlSt2e6fTxLmmz5PJw3hTlpoX
MvFnx50RqKFL0HYHvG6zM2Lp95BXcRzEhoY1mPbHqfdtmZ7rG3Pmzjp23yRetIht
Rc2FSlKYwMl76g8NuNZnEz4mwbN1ezEpjMoaVySbcL7HFfxnfyAz4F6CKY9bZy3R
ETTSH7Yf27acrmTlIJVvuNfk5rVn3pbN11xsCg5237t5ZqsDGsh1nJu5ODZ5UqHZ
6b8YtyvZHjhE9BQsEMzFBJSUF8e77l7M9dEwUsaE3Lsf9IqYIRPcQJrCXTlwXBx/
nryzrq+ifn+p6w5ZxzX+n9qNj5MMKhLXWCIkEub1CBNZRH9lyT+33w261Td/aGBh
TOZVSqVtdvcrEz61NZ5xhOtSu6oUnn6/6LbDERuiNWdSYBLzaiignaEYnwFzUWgi
UWyaSZEUfh4L7dfHrQv3BBIZeS5IzE4KI5X4Cj6HI3j3XTY+pwqyekeog1J01/oL
DBLxdB0SONvnfmbQ5sQy+lIqDMiGa9/1iowPJIafSLPVELx+y1wiIWGvszBDswdr
+oivrHKpeyBiKdp4TbzdYRSSQiVS8qtZSm5hKjiiQ1GeInHDl7C5O6EQDeS1lOdV
nGRzXMAGZ2OE15b2/K5YtDBsxgUrN2JydichOSlZU4pcYCMYARaYalf44pEFgwct
ZrWtdhjVcHGmJVSnDrjWPBga935xDP/Fdf6E9RMyQpG63uZr5FNrqFGPYhsHiY1j
l5mGqKdHUfbhnrQLiQ4iKDR6qrrGVV6q2+t+rshXgu4qtnORVUmfE3XEs5TbhtG8
M4EnmiePhAcrVCrOkfE54wBtJNn4ZsgRTHFlRVxnYpGa0hrOwUVxXMck2pdNeQ5c
`protect end_protected