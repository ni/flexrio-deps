`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23616 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
laSUciT835LU3jKjm48TUBNExw+LyfGj6IKL565zkpfKS1u6CGDoOYY2p5lnMH2l
qViFU7v4NYqLq9Il1HhjKmzyQAANqYxjrt1zJgsjMe9hkP/NsSV/dCxEvHRciMml
H0r7FLP8GZPy1dp+SkKjdbltJaevokG5/9ubC/XBHHf+Nqg/s2fz82Ryqg/kKTP9
2FHApvenlLCckNvA+ulYhnTowXvhifACv/HBXzRXUgf5QlBfm7jhREkDrlcXU5eL
Bic8OwCakXKc1U4RW3fsc3cPt9UhChk+AUcCO01+g9fIH5DXf5cWHFwCAob83Ewi
d41ULyIh1Alf88swLGGQsHQwu27eoXDYYBQsAxPDxdg18DT8Z8d2/00XXBZU8nLO
pO8PhJsIiFk/Z8/GDmuIEuZs0BlChyvEgInHKvXQ0a/JQomNkA1+0MWxY+xunOXf
VwMjBLsnBr+3BCrKagZ083tTQeKckALwCCn2Ka73rt2W7qsUdMHlQnUaJs4V59KU
VFp22y0nvS2/V5FprQs97EdXsC38e+wEyzYKBr+hJwFBskEDI9H9IuupVDGRBWUb
Az0JhdIooxDsngwAMHuUSbiJiThHw1/gLhb6g+y7zx7Dk2cZCRK/K3NUoxya0FVW
j09+ZPt/n5++Bg55NmwTH4Tw9mtfTa2tsV5HgR7XKW5o2rg0sZpqUYf90adqygBS
HxA1rlE9RvtuIXR6b+zhjkhgT8b0pTM54BxAtB+wEEW8lILHVMPtrwpdEAYE2xtv
XIbsOKWv4DF1HGHzZMYrlgAXAArbDcuQoiIkg1xoVytY6t7Uh784mRCDJAxWCbOw
h2rnLxaJny/3ZysG60hlYWFja7sdZyFF5PaDlO24299zJJBB+UuGJ6S3CQHQxoJs
a0QjTSM82ca7qz/PdLKHKgOVs8CoPg4hhYqiLmi3mi/YCtbXC9kmPvyofKgswrUJ
0d/xRX1dZ7sEkYydL+hgFlLWWjn/DY3zEIlzjp59/0w/jy/6LmrKDzEG4Gil5ckg
dRAPq2U+2hFUxXkHU/j/Up/ouqQSlcn5xQIMLHUS1BManPbRMjNRaRCM8USmgrdo
tRuHTdrkOg/tVIaae7cEum5LHDmovoyt/ZK3pYKsCbH6xvP52CF/xb3JaJfA4kV2
yf6GB0xBh8jUNJx5rzhOz7fEEq+mfj7GdLuKra3rrWx/f2jcsnFbY9bwVwVm3289
c6Ajgp8Udzu/AiyNyo74FeAONDRCa3WWe9sVu/CUBwqclC4EgDd3kcGmSls9o+yr
cCB/neVT0y7Q3fBiFqthvxXk7JB7h5bsplOGWDRrT2vk8rWztGrf1aeLt+xCsbok
XFs9pFEbnaS8Qr3VE1+SxGurm67+N0k5kXLNGaOuw6hC2wOZkEKC33LsZasAA3Ep
HoSSnyG8+ETbrQFtpJmwQEHoU6DbBTBh4s0ek/PkYzWQtqzj6BALSwpV9/EQFvth
6R7Dlg2qdmVAXanBteipgT0Hmiz1uA7oCITs9i/DWkqwLaBI9guhCq0Ou6WpFEop
/qyE/u45Lh4S5t3/iKiR4Tv32VIC/xAs3OnSoGt8CxAiEfHtBzV/F2kHmOuhO0tf
Afkr1Ee6mm2PF91ecLUHcWbnr4wEGS8jlfPyjBu+qb7dnlPbl+93C2JAbTxRN4nZ
ssABEICuXWmRX1Zi9wGdy0LPETuYOdR1ByUFpsw+IczxKhOr+WKxvKV30bIw44xn
35yXJyEVL5FTOXjqkQZiqYe9F843KKl+m2LZsgElc37K0e4b2ABQgCdxmbBD6s/7
NrVhHMg0lUJYihmmOkTuDPWFqrz8Xj8jGxeQtJHNkku3xNeytObZSxqTS8OI1ffR
aFkUL+rOzz39bchP/M5TT61gRCr9gqJsUWCmIgN3wcOjkhqn7aWxd3JtnAJANtYK
pYvLaNUKjoqR/f6am8zPJd2aq9MwJ2WYylOloZznBF5uaE1YMHZKXw7UlAeaGhop
lW7Ks1V1vSYvkM0ytoV97nY6wkILZb3E1qqTzpffjWdhUT8XFxkioUO2OufnuxLy
ZLswhR0QqiAxe0NoeGzZHmd5QndWceg3IDg1tFITS88BXLtKuI3adx/nQBJf6KS0
7d0xRC9hi7qgdXwIH4ag498ecFKe09j1xZKo+nSyVl4rP6zlNCESJnRxpqVRnCPn
H0ff9x8iM+oOsnoHk8+tOTAkGJQqbb4DmUTcMvLWDdJVh78+0ymlCOtT1nVa+kGm
yrwh4eB5JpzTz5YFdNx7uayX+tztouOptGIyhAxzphtES0J7dWhy/WF3TGqpvAUQ
AFqMXs42HP1oIqgOcXOidWnD8dGNvJOi5zRqkg5Y5V7h69+IaENqBG9RuD6ajW//
g3RIzwmdneqHS2lyusFOLPxN92Ff32Ek2Z7++YdmNJV2qysk+fjrrssrpIYg50f1
RymL5KtR8kwvAQgifMgpV5qVfnywDJtZsED6dll0L0LfUp6osI9bi8rG691q079+
1PKf2EnGRHx4bQXUDJZkHUiPx0UEqTvw9vgQVagTt1qU8Oh6t22gkbe4VycMlNz4
uBYXRpkc5jEA9dBwwG2tcVBVlZxlhzEWHFbgGB/mTTTk9ZiaWTdvASuzhe3Xieip
1B6rVR6c2PBaarENb2AQeKX4OGrFAwH+CmGNN9ExjBQKIgeRYlbI1t0suZsN5l6t
7MHJHnWtnf16W5BoF+KXyWjJBUh2eaP33k6XqubjIykSfm6HMcLD3Y/672BU4Fyh
Fm4bnPz++BCf2OreAdHknjRohHuLBz5uURy88awenNtLvsY9Nbccsv2++M7uviGW
1wYyP5kbMBBSF0qRIIVpkqTR9B8IGpR4ty2F98SqimnaR2H4nXZ1yhuIvHUV3J+K
33kNySrsBPLhnntpKemfw5DX36t/AyfXWqc5ngX3x3t2sD35YapbgoWt+hvkMW57
RPx8Na9Iua4EF/EZk7zvCONfaC158GckMyLvlvJHGhbJ0zNxbH/avZLRrjv9VSb/
28OpNn6yG6Nir4OuEc2lh0dQrtEt4ij/jyRq0pJKNQq8juW717/xH8K8CLRgeOhr
kh0rDSyoOEOAujUQPtCJpRsK/Sp3NXsjN7kE0+ETDRWEU4LOdL/dD+LwSOZ+sBKN
bKs+PR6gYMlFIk8B1tw3j57sXXdpA56o+G05gjMDaQUjAMhGAzRz/AjmOIcJzUd9
FCKt61gg/GRrlxVQ8zsY1vtjv7h2LQx15bPXigJmhMvoMq84yraQjRhXeKKBTPF6
+qrC4LJs4G0GNKXG05+JA7IW/jr3LB2hNIhynh2MzAVam6ezrBIUT5qkiuh+MevO
hN6ZyfYdrpL3WHcY69rApurBH8VAIEVX8xQBTfJECpvmIgpdH5pViHW2Dioseh2S
Wi+jsue75fruaDG2C8XrKcgqyzUhL8g/SqsQtGXCFe18xowFl3WtMwcKWhNMArEI
VmJ0QHRhUwr0AZr7Y1gcQb60q1JWdSmMg/No2AdaSSzmC/Umz8yV0t4SBK+ZGskm
aUPvhlCiSQRtF6gNpqYxaTaj5AmbCbsgFR6+DcRehYqwzg83DS439HvCMaL076oh
3w6kWcw2wuaLQL5qD9b8f7GHbB4L9q4g6iz6LeVajTWzRMJJMprG0XXFPpKhyLAG
CEiwpQdPfMsSxGMuxfUwcwDwQgwGljzq6DUb2cf8lg/IflrTLqe7ClTWRJzzncdo
BroyfboIWg/UGpg31RLIr3MfJ9TNmovajklEH2HS1T6qJD81SSndJzgkuteTnVeN
W1JLPS+mUNcK56hUl9cWTsPJTGLiKv7aPAmThybtS65FS+kApuT9pIIrBRCESxQV
KlvY2uvqF24fxULN/ZPT/vVa+qcpRBQ+H+O79GX6LmR7Bd1pR8pBqoBpeE7+8pWB
0ZBdBU3e8tfBP8RIx2wTlVpyoo+80HGGF/HanzScLFlChIEMKajoXc69ElEOi70Q
QRTTbC55wDtZNXPo0CEtSiDWC8gg9lxXnqSyf4loqCxMyEWC7yQI5pUzEgRPNpzH
9o3TjXdKVoMgn1LQy1Flx4UdZos9lGPRLwP2QhJJrzie7qCC8eEtwNnyTG/icZk4
9RHWmkY03Sw8vyXtFeirZzqQvWOLvdknOPOzmvTPdPmg26Dp0sTrr1H3vkd3iiT8
bOsv7U5IiF3f9S89/IbDSCehh57lwJlJpJMIomflZMr8UuuKdDEcV6OvKrfdpaRV
uqSKRjq33njl8RMQyGeGGGAbJFAp9j7ySPhmOYilPyErBUJghq1gvjztehCLPK3f
0ZWJMsnj0JBJD4mq0zGiLQFt7Ei0kYl5c2+OOemrS5J2/LP/y7XSmwytDor+AIVt
p4GsqvKQOt2wAg26SkTUbZ6hHiZo8RPI5oYVHktAeyQLN85GJeKl/fGKQUnoYlO2
Q4O5jpKhDuDqbPiqDDmdKVovXXd5dzvQ/1VSQ7ZcE9Oskz4W9/bQai8QDayYsyQq
Ym1ZFoA1qUbHh3Sc478M7dUi6LoPgoECEopbyn2xIjY6u004BoiTON4iM1pg3M/O
PArg9u1DY9EvkyPDEL53Jj5NdfM0169lsoy2eolL0cx5nGuehQh24Ct92TTznUKH
WbwfN1Ub5Zk6RCWnpcIIQzInfAY6i0BTNlthah/OIczxo9/e0evQmAqSvmpjKunu
9B67Wvb2yiAtr/VgAWz8hecMgWgPQ6VTSlr3NXWCVFnbLrGF9AR/CajjhpLKUOrB
QP8ieJrYHK22/7M28db0W5QFGJbnaPnhQcuPTKMVwxUvgpNszHNN4yD2Y6dUUYqb
XzdOGi35H+QNnuKPAiuhOfgsuy005Wu8KEfYYkghNA1FHX0VjXF5AckcU4n4ZGl9
XlbcCRPLNVsjxQ+jZQsdSSB3Mk/VX0buR6yf7BoHAJwECaoEfnLet/bhygYiUPiZ
3fQio9P3QrphS5NPsgwHwdBkLiNTzVYBpna5q7LBDjYuv86Naf+QEW79aMuLK/j8
hXgvjGIM28u061xr1+YqdAL/iz4hK1LHZb4NnyPr7alpNeHjgi2LA8jGCZ3Yd34I
1fWRSnH12LLj8CH361ku4krgSTq99zAWZPNh+iaOhBVOCkKxHLl2lzQl+a4Oo92x
+/1Rzbzl/c9Zw74Ue9oPGqcHFjmfu0gTjoW9CsZmcNX2RDavA14sftnmug0GSFoU
/lAWxTSPWFctdXpCpRykZ5k+5CIr8LGjX3KaXetrBcC4FDECZS9STL2soqqrlWn6
kMm6Uj+j5IjHKBw6SnrRS4Y52ClX5++9YwU8xZeAFsCm3ljzEOmPNClODoCpL4tT
7V4l6A5IXxd1pqXmd7ubxdoaUrSMTZ+4f+Fd4LRO82/0Ctp5Q9x7NfNQyHp6/ktw
0V8mjiwby6+8il+ZwzyvvRtdSE1I5FADEH6+wZAy2KwjARPEoU5a+FYC8El3BhVU
iKRMucGNhnLAlB9Vc1zZ0WozO3PG/vAU7Ly3NoTwV/sdumiHHiixBRR94AX0fOtU
tY6q9KbCyCl4yZELidW6gFwxbFy+tagiF8nJlfaTrDvTdEhfeTciB+fQuQBib9eH
/XKsTG/wGSuwVEOoyC6r1y4pkHdr/GqaKOD0vOu1m94EW5aJhp8fjsSRfkvPQX3U
ovX9T4T4irG4ecVyBegQeTGG1RPeSYYBMHaGD0AJQlOQnly9bloF1m/ELV23MHRN
7Z42wApAtB4Ut/O3OhR8YE3PCx20IsYevgRP8ldz5vO6civBqlfCYpKQSqhENlZ0
tAhbXtIQ+eHt2hCmdtoWksTxBCoHmX/8NNIfGrb1hHxhklg+fsUickAlqwcwe+TB
n8adsKz1X2flcubFYyHokIdq9WD8JzEcMm3Tc9laxoh/Gc1yRyrVvLbkDyREZIIr
DGcHM0LGJ8Iiufn35hWMx4Snc9dHbzTFN9tImicOKgI5+IgGoqyTvBHov9FmyWIl
h/HI5VQodGinE/uyRSYM3C0v1ROEV5l5hotSaxtNO8OygZ+G2rLu/RYTApFMCIWz
EkVJDwg5gahhHzqXn04UL0QOHRT8qYagwyHzUKW0eE6k6HivW6FdFXS9YtxblR0K
ztykf6JETAoSalbnuvFTFNnF/e+CNRzMVcdwcunBKx+uTZs6HClizIZ1NfE7Fncp
lb0uGes2OvRDKhINYwgy6rWVwt8QnMJ9Br54Tjb8uYNhlp0I0dsrYYdjU1s2PBEZ
fW0aNu9jCpOstOpHe/TOj9vnm8Mvyngz+JJTFQSyizxlvj/SY4fZeZpo2tjOxtta
5VzKE4qAt5D52KiwH9niKYqMn6jSfoKKs+uwGdCc7+CIU2hK8j9AxJlbQSIs5Tfy
eKUizq5gSYbH6cUsNgvKQjrOI3f9r9tG8QDs+AOBxuDbIR75PXBoNVmji4fE7wch
XhoWl7d9QDU7tseROF3vcSyAKMDPJ4ydxLi6K71+U/5mJOSxwymSEfnvPcTgqCXI
9gr+2s4fWr4QHPSJdkUD7trIjKaPGVs0DyL7MuyxmBIUxRpBKyoEl2htNguKGdrz
xYob2odf8dfABqyHbLQEeo0VmUpDSqJr/kfygrJ3/9xN6ZNsfRXeWYl7WF8ADuW6
3z7lLyqh3uE1xW2WdLB2DvxwuL4ruZ26GFQKV/aPxk0hm3BLABZmPn8Yr68ypG/B
lRf1si4KllfCUkXmRVyDjPd6qx7xX+xQKDlSzxh8EhLRQ9HmWjySNGMJjOF+JE1I
sHwfN4ZNR0Moamx6wFpQ5vmiUlScYtu2xiY9FgKxX43TVe03e32FMZILUFJy3i/x
K3ETldNBZBg5fgOMNdizLaomWHls8a2B6Q5fDNrMqtkuBwJ2mc1wqc8w9O17VXpR
uAz6lR3/5kttUIqv1MlQ40q5d+7Nshd9VtpLMlLsOqgbC1s8rJhmsyHgLeMTH9K8
8g7qiCUAhZAAcIzMQqwam4Ji5cpYXRpOq3KneAumPKVFt9p3W3X6wTyyC1SGc0zz
1eJab3iqhHJdJOU98xaTDD3m+9kjLkdteU/vVlbP+vB0mYGpi8t5cKAdYxo8er9v
henztM7+auaFlAVS6KA1Bm1Z01f2NJlfBYym7rLv14tgha8AQD5gIgx76Kg2MOdg
gcEHxt/v4ag0oL94bacD3cfIaE0rjiqe6JGrlxX6XysW13vXZH++IeFrfAPxeIZq
isGvqtvv1tLf6NjqELJXLruYEwxyihVRn6f27ZTlcU5syp2f6QYihFvFEm0GoLV2
1upJOydXSZN/fFXp7Tibgk9bJjqaIf38JPu+tpuIGqf77J/j2XkbB0YXzTbQzQcq
kDa6VLngoftrIKGlQXir8zhuv6tecsrkjzB+38pRdj/sGORCtSFsRroHjm5CYpK6
rHy9Eihl19ALuf+/tKeqewH/I3QICFeaTPfU6/n5zoi7jh/BRn2GJxgF8hOQv7sS
8GuWMhk+e487LuwAUs7IeIDSSoD8CgJovuedSOuPGpz9Lxiv1VGnV7DsqmFAHOmB
MgImkUb2klGoxJU+jn9jBVgI7ZUdaJN9LIcVyfoMClFvnOvpLQckAuiOVnuGNdSy
2xngWOA6A39RLQLgQ+LHyCHTsY5stv0Noq17ZuyWWydcJZXSPACBnchAHf3xhwGD
6zHojDQoj0FyuS4srvpfNJ9Tt1B7K9U3EwD3HdjbuWSE49e/9+FgKKh6SwQ6Ng8N
0ThRIPyrXVSxR9UE2LlVk9QsBR3pLiMty6LkXjeQx6jWrerfJzUeylAfQpgJT5jt
DVa0U68MJGzDY7OJi2O0Iuw6Uha6VgKQDsdso9/gaUaTfHgkEuBGm/nybQt/qgeC
7nPOzQqwRR6kQUQ6g7Id8l+hE5OLDl2XEAQ9uM+CBFqrtF+ndaViu9eGKq/DgTDY
RZgoGUIEfxPM1Wqt9NOCXublsNS18nf2zbhZemskOGwwBAKjzDzQ5eqdJ/aALOQP
x4KR5AHbGOQMM9Qr8rC1jP2IQ0KZF+kyd2xlDn92zcFlhFXH8dVtqgxLzByHNSzB
LZDnDrdcYgQsQBNSXngDPA/KW7ZZK0JCNwWfTSdf/Tw7kFxULfHtTLr4BF2+f+LJ
bu6DsKCnPZ3Ei9YPispvtCrzd7EpzJDNfEEiLg5jalMuUATD1i/Wsv7wQ4rIPieI
84cBF8IuovW4O50QBpbguvW/c5oFhPRs4vY+tyMagLccRvn2sPiak1s8J44+Zmwu
8KmUSjMah8Ihzis3homK46QfgqSxk9NYO53Qh6Y7y+Wfw/xgXwbGpclZz76lxVkq
Jlt3F5l+GHCQNQX9p4d+bBhwbZ2McQyprk4BFnN7FRWFsaF9+UpqQsxbHmvlxKf4
Fj6f274VeitdzZdehhI5XihxlV3kxet08TrUjn5JTyLrjPxqvNm5S43eNXXFzUl0
iuc3M7gQ/eDc7hjyVt4E8xclUBQ2H3whtv+o6v/SQUHsLxtzZMlna23mFMUEYCr2
IAZjbHKm0N5gN/g3Dut6ftUzdoECEc8aLyziizesUnkm7YZLQ6EB+aKT8zv3AvQg
23ySmNN3fi9CLE/Pwi3L+3/T6UnkrFdrKm0+AWFtJw8gYOdPmiuc6LbCJ26CF7IV
RaW9y28IOLnaK0sLtzpRzbtDBlnLMlZCS0EUW4IUPx/uHSzrWw3HrRv74dUniAz0
7Ni5FUUJ87UgL/57416G3QIy1a5LT2rUlSF9NuErTV2GLEZ59kPh0LZw+f5xGi7I
OlJB3ub6E8y7Frb0VJcLcBri4cmsqC2f2F4dSoyy8p9xh/5ZZ+rOlEJYFGmCCJae
hl1SWWLa8ReKfsIBUBQK2+OB7l16lv7KZaP9D1bkX087WZ2fjPLmu6M5+S73WXGK
NPntoWy7k3L8dbpVjSHjaaBhA9spjJ2keNTysQ7u/h21/3S51oJ+hzLUSZ+2vCdO
XvVl88opr851bxXMmshia4xpZ48nL9Q2mGd28Hmc5CN3yGva6yS/SoCEJNks0pol
dbPKvJXi/AJipJOuxZMHFWq1LNWE/F5hLkPdrlN4XpU+uXX6KGXHBIp3FfBnql8T
Jzmozkwstf6RrR6VRND/pPtYlQQPx/c1jur8Ulo4H5AFbhzgwChelLImDPnCM52f
yZqh0Nb9wkIUq36je4z7ZNSB98S2N3eJC5RkZHSxafcGOMJ22NpAFwgcTW9Y/CsE
ufV/LVRm3YvXiJweqzEkgS5HU8moWgfSrDqlAU6H7/0zaM5l7wh5MDUUD9IhpoMP
JPz9S7lxlhg2GGG0EMwAZW5qWUe2dlF7uGQVGF3A+Tc8nP6Fc4ge1Sjv9qgupOLx
M2HRJVrrO8/BzS/DleP6MzwfOJetqQ+RL9VwT0rTmLO2BQPgBIechLIfezS60YiX
14lr1NU01KC7KCyOq8yobcs0WvzqeLo+Wv0jSpYHgo2XU6L6JEO+0I1xM2VC2jL9
GwbpfXgt9chJwe+LjOtGBLg0nQrNhlbyBgvq9JTld2tyZE6Pmdb4PiTf2vemxLfI
4ZFYhuxQ0WTbPO4rXeKcJb5FViwa8gYDY/FvXvoAXVeqPvKogVNMYiZNB7REnZYu
QguGbuNLBq7qegl0LP59hcRv4et38ZjCByltDCl6vYKddYkH606OGVEtJEint2Ey
+OZPAN87rlw7CII/zQGq4JGw8Qsr+neXMeUzLDbJsa/xVUoI3tSRCSRV4lZuj3w3
fvRhMsaTxsIeJZaUtl7DSVQ3nlIen3RELNvnW3JY3lh6ktJN4NpM150IQxDZhQnR
8Yp/MpHwGj3t3hPgdmt+2LXisTS+Q9C7B9DhV/uFz7tK3D9CbxLFBBt5K6HeHe91
DXQDPDXogWylrO/WMuFHB6LY6TcFoIgqf7Q4AGfAXE/x9rU2bVG3V6e0HKUnBinP
iSxzZkdqKa17vfnSFGSf+wb4mxjed1UIxNeNsoONPqgW66ELVLhzowi90TnTPUnb
GYxVDNOBIqG+n6tnbYgMGl1D2MHN9R51xe4nClZi10Q5uW0mjaj7wW/E+W0HaRAa
cHH/elUrkmAryeBxuDukTGzo/dqErw03yCjsy59W9mYuQVXQcTs5NZ0KLTkYUHLu
jdjisg8Xm+ymvuWm7DMyn03tJQXE84RljmHc9o3sYq02qdczk2pOsZHrnK30H516
NBA94J2HPSaX4GqUJbMv+YghJgUwK6hlOAbb+qa3FDSSv5Iar6KuPxzzHRjD5o5e
/B+KFoQSPjivyQGsg250zCB51Wrskw7kXJ/WwfoWVqAHPG6kwBJA/D/Xt9THQD+p
aIg3xi5dpmzBB+um3aSWWFZvsD9r+f3dITOd9HTPFlQnXqkZYJ+ZBiZ5jyufkMqP
6hO40Cb5iR+cA4CBWWe8WdiuxUnLjZfx5PXBHSsV14lu57rjIvuFWzpFxNzluYcw
6xqov5WobRAXjDECwZdW7HkB0R5SIVBg01Fr6U7FKZ2kh2ROXUCwLZ92kr5wHk4x
lvmKF+vKS+VjWeaW+xojMV4dtaHbPB0NK9daGAemz9Xg/BF14BD0aKAqCoGpz2XQ
Q7cE6N/5AVe3MSjs0LX29Jha3TJ07osmaT3vm/IWLuQrNGgg6/NuFwvg+Vxs8VeV
cbYiontveY24smfcvTGWug9XgtfsWmt52GCyrhBh5bJUznR2nBGk0FjUpgaRQLd0
XOKEBUcFJYOi5PdSaO+H/CkioSNgWmY4hDlMl0wRMVoeiv6LSH1z8CFKB8PvMq8J
UI2wjB9c8XtKEGfkCiMm1Eml7TXMKdI8MS7ZiDrM5e4Y54fRXqvwssF3uNcW5oJL
UzNSjGX1zoHTJUZcLjsOOV3FnbhGsn/UQmrShEBXEvKwConSU2JFUeEB466Z3XoN
/8jBOHgp+F7iPExbzTOENFNBmNMjQzF6ePgYLY4YfgfXzmGqSuNYg0a796yivUGR
rQq+S68bNho5qMMVEhU4jMr5w/LiP03p3G/sxZIRcD/dbfyZRU+1jrixkU7gVsao
f3NsIjhVrqhVRzggDgjMSprTyN8w1n9M6z4NoxDAnufg+8dLTzDcwYlgwPt74co3
q2qkS+oLVxZn0why/Uv0i9WFhsr7efjqSVzxrQ+GVLUNf2g0vb/j6tVADM0Jx4Jw
cWL/r9bPsZ9K0N40+vVNDeFdqQfGTHoTFj9wMSmi9bumvpEuQGkluxcjPlIDS+L9
LDeKMUs4MbEKIx0pBnfUQVpqjVfEdPq00Rfc50yANYtiW/tHGQZwNoABXnm6gZFb
/NzwZn/d3vO3cEqtRjTjuYjz+QJ20qvmrdHcxz2+xKaprdDvTzpTF0+/dCDDDV2b
tUFC62gfV9XuPPp+HUlQtKeo/rU0GfzE2S23CxpyER9TiTa4hPQ6E2LAYY8dqOOD
d/Htc2lgFgRSDbKr1DHcWWcAoaGPCYA4w0hLgHXA3e63Xe7if3+m3lEZsBGxHaXV
KVAasKdvuFF66v7dGu9QJMxCjcB11V0fVxMXKer8x7afQ6rIuMhsiIQhIIpIv9rq
vR1ZjiBoK/MVNKZkY+FcdP1CZD97yyKijPVQ6ob1glxDYDvMfP0iZXX8Cqx+ha9P
j2WpILJqkfcNxJx8wA8EWO5l0QbFn3xnfqfBK3XDT36p2NdA3rKseCAkaDj/amTu
AHXxHGv1H+Rv3NdtALrOfzZcZhTADP/U3U81nxu/Do/VCvQt5czUdQhdDnAN+sYh
u9VDgg2sME6qKmm2iqdADWCcu72buNUaNpYimEr9BmTEMBv4AUkqm/mCylcU3xb9
KQc7KTYNydvfQTrLXG5BVwoUhVIgue1X44ErPm24/U9OKV2v52PZ1BktE6BarT6t
ifUIvJX31DB36sni5QnGiAw1Q2mP4QNr42ek1qipPy0jYeeyebeGnVrjHlWCUXvU
m/rcWyyRTy07max/ApYU4+edUsJ7b0rohBQltP/K6BwZt+ei35WTP0Sz9ZBzcOMx
F8Ie3tvRh4kbb2jVUNvX+Gv0bWEg2Dg1sqkBHli1wnPEtAfiRQwjhp3CFsTgS4P8
K2YzN0cXvkW1hVr9e0ER4TTbIBqmg6HQNC2v3rHlagiUqJpPIFa/0UtPUzs96gZH
6x8MFZ0PMyV+OfLGz+ygPmWYatENpU+n1CYTQDHen+KtA6TmZvfyeMU0ycdHfnyD
9lU9K3aslc+r9awiI25vJiYVITDq0arKK0OgDT/pclAiHWdevAgljxLMRSq4VrPd
PeAn7nYn4fYeSq6U/oLud5YkvThPimPBtycp0N7Sgr02K5V8erDffJBOczYJOQIO
Xgk5q40JoIIivx63PyGN8vLYWibXd+PUc09zrIoIDMc4O0pW7Xq9raZsUSXkN55B
mcDScXXuv0aEcAwOwkuWKCxT8dFBerMOJ+Fdan/ImqTZdk8HUCpxLIDAz60hDZjl
9YG8eDkmEae4paNCtN8bbhA1blIXu54FctC75tP/4LNsAtJZoS27oNHkvt0qaQ4i
PQXndnRrUkKdieyxyFh+NVVkiDfmGzTBN9lDGRGr1lk/YxL3Q/7fM3HEWSnp4xNn
VlJcLZqVn+nS/nbqRFzbCoCFok5znL5HuslM0bGgekNF05VSnGnzRtX7tOVYR7bZ
f8E9Mmkzt4xfxBHfo/4xtCwbfQg1BVv7SZcIibIXyIHEhIPzouyG+c9U1dDGl5EG
CYbdPtGwUL5GlgifVHaOT/JWEBqwq/mGeXkIrKR+9IMgqwXRI0XnHWV37eGMWftF
OMIH8vTHlj+AIEoZjBqe+wC6sRIGn2S1uqDdsJD7KVEqoCMGtSbgRNQz86+BNXsX
7wfNF7u70TAjonkJRPQqvu/bgMT5jyVWRNkgXogBfrWMLLuNMPQYYUN5Gj2Unt3P
NIN1jydOB37f/xTkamn71F4ERR/GEWYEG4iRgaawCFdfQErQOqP0wa1lEpXLai1J
NJ49t0n6MkyXmcPLMWMrKvOAkIUYq8TruXlS6s5P9NmCZC6QPfFQgeDlelRyD9C6
14g4VIWtXIN9TD5ZiuhPYyTj+6Oq5uiQ9Cbi//1i+R/e7IkOo6IX3lA384i/otb1
ulEXJUJNzNjS6VOFMYkn9Owf6MmkL9p1g3LQDgDG44SpX61HW82LK83DFSpXt/aq
89coEDZixBSbYz7iKf2w/poLQPx6xSOaksizrDCXRjbhE3SK50UdUy2qSXWwrWYl
kU/7TK6ok9WJNNYUR0BIp2oq9XEM4ecaq5BvogsJzFYInleUFdrLpcm20Oilckqx
UhB8oMRROSrcxCau4km7Ugjx+CsT/F+jtQv0k6i59kGyr8XSmcDqAF5Pmc9wyog9
YKCT4qe5y7RYOcvV6cpDUDg21JKP1yVBs09hpIu1fO/vu3EZaGonRX1KbGR54KYl
QLiZGLZd9eeyEMa2wgUmQp2YIEe/4Fl9gHg6+ZKqX6lDW+BI6kYIBDI4HwFxZ91v
g0TxBlaXt8Kk3CB7LXuwae+Sg5vX51aVU+89rIMFW1ZSnHTxFmY+kAIleBFVolQD
uTbFMWF+RJNDyhITmjcWzNzzREP+/3LFXwyrCdB92b+8Utdt9NPX02wQFllypXEo
PDaVPF25p8pKHO2i59FPqwmv1bbq4AfnN9f3j4dblPNeOsDYh4FmRS0Z2thv3iKg
qYx6LuGU2KNL6HKdphpEZ2yUbWFeYg9rWXlW5awcLVu2Yq2i8u4Uff1XPPqUkclD
y3hW7HIP5GC2ca/8U3HqXq03kGaelonKmKb3ZZRr9XgYeF4bVukR4jTx0+ls16wI
QvHb668Brvb8GgiptAtqOuQr5pMplNpyVwp1T8eFBGtX3Yeye99jLYksfHBy8sEq
dWdC1cdvjZuQXI4/lhLzetGW17aDTu81kSwauMT7iuexyk5KWIXRCIKB2tzPIq1M
NhSdl0feBTEJ1nNKib3B3nidBEAjRoX0D44LB8An1XyNaMEty4CzfZSneSTTpbSL
EA/8gGelcXXpprkC1IP1T5E/Po0fnLf9byqZj/EIYURD6ZF27N90I9fJ3MkxHWn5
TQODpeff6CAPPHY2ihMGKSw8LpsrQIxJk6JnzceZAqvlIHBq55z9fg+IcAAHSb/f
682dKWQa2UMJrD2KPOHq6g1qpZy/pR5DFc8Vp3EjEtZNFwhFBfGHk3nLVCz4ujwY
HPGyHN0xIqC9UPlWhRkoC7YuscbOtssZqeepTTclNSVq+XthLaA8P1aDakGN5vzy
98DMtOzGAXTE126VR/oH2VAsWH5eToM/zHHw/x3Uyxa+iOD4JhGCL08H9aFXGPPx
5z0HzF51+o6DbgTbLiy90rS0QCvcSPQ7FNyfbN5B75GBUcUvYhyM3/jKviVhSk62
W3KDxCEx8Z4UJFZZEYhEAsUC1+UFrqFrn8lHw+Ptg5fWoP4fOd4FXZUcHOHLgpwv
iMZzPpTT4pmlHBMQyfijamG/zUJ0fpvTuhIoEgB93UxacwTTYK5iANxIXfa1dTYd
Opg3d3/fDEMDX4YPXF4skIa6Low4oCDq2LqBK/Ea3HUjlZfBkascjbNj1yqrc92N
/Hq8t9WF/6tqs1BB/5KdZF5Fk5LbuuJtN3P3xQ8gzzIaz+6cR8lLZeIFtO0nYFiF
e3k+qSiNaH4HBPQ+zimi7GBNxYJeLSROIq5nm2zWPRIdCr+B3aEuZTpiMRO9m06W
ZA4JVAlC3USqzdVeK6fS9LueXMV6ioghT7W49EiaQ4Zku++mISNN4Bsi1j9he7bH
C411OXWpIxRxK65x/Mt5PeMtdwdh9rZaF9lRUA4MNgxshN5VpqQ6eHDiUNgCG6pQ
JfND6mNT3F221kXnnO4stv4EZW10o3zhk2E7AvXPT2Sf5KnNdC+GuyLEh6tETUMg
qPfdOhoQSCV57+O2AF/ZzNuNaJeCrLYericapA2tydmo7h7VQinJUSjLAiIodjOU
/9lrKhsq6V/HzUWFK3kVmIIdr8axO2fH3ufBOcoX0S7U7Gbd68/PO625xYL9AhiZ
x+B81eOREu7q4Q5+1Ydg99mkpUWeYTDUx/pO0vGYJwknxrT/fsn6Xbit7tuwC174
1gf0Efda+94/PhFhmi2D+XLvYtp25HrqF8WUCQiD9jqePFknffCIHJkfZlyZRfQw
+ThuYmCYXNQr2tYeqGg/9/5YKtpvlyBgw8I9j1f8ZthZ6SkiETtq/z/euJxDSoFt
7zi1s+RwtcQRKZg+yNA9emBexugqAqEt/5yjIIwod7hmslsSzBlyEQUwudPzpwqH
km1enOk/VBK/xQdydnT2CHc5gQySSTf+fIEAFZKx3T6U85y5FuW/Jw/rFUVfXyN7
MYsdmmbsPR9zX4ImlU3UdhjiVPBIsb6WQFz34B+3JkXtRafzXJIxvB8qDt3CrBP5
/P4VCTGm1Lt2smugc4o25bxhC6zzQpwkmYGKxMAiB2wNsZS471D+caoKug3ZA7uX
ey5nkxl0sKFs9QuuYPJ9FP/Gkx112PObr2L1d586qR9SOrhEEOBVU6h1dzeNh82v
FHNpjlonyuMRzyIqlaEw0TptHcYd1n6cMR189wOXA8l5jsEvTFgwNvbzGWrhLOJG
zgTQd+ICrSfhinTwE9F1L40qxIZ3h2mnbejkIMPFeUmF8XM/U4HQYlSA/Y/U2Xl3
L7T6uIJ42TKPZnsZKU2Z3As+miEl29xsWixifhCsNX1pxGnTwSKUQKenPmO2y6wd
hz8rQ3ZPVIfLzPBlJlopTjTX7KwBRR2lP+eKp7wkVA2LQNaCItsafhyRScHYSBGM
QuqfwSYcUi5FPs/OYmieNgaAB5i8F0SMoDvM5cxQHaBWSrf3hTVfV6pJx0WsW8YV
aU3EoXH2lIRz5NXY0m11zYuX/jlkzfbJ3IRYyrWzJ7/qShodb1Ys+nVK4pF6LIx1
QWCwYShARNBT2X8c4weElzKsGzISgUbX1lZ1AWLzvMk3f18V5RWcsKly0M/7qmTb
wLZTRw0QCtQtxooFCc0aMRx0CfkVVDX9MdPlCxNk4sE9QnPkWhGDlyLbFli4jlNS
09gTXMZB50HKMpTLxYq771n7GoS/P/ZnJiljbKiKpY6rEHgTsQn8fiDeWLvQ+Y04
VeZqBS2ztR11eBLfO+v4ar9vI3Th5GPQnPCboHkowtUQjK7e+hf3F/Z94ndiGr1j
zjpTxq+5whEegvlvFtBnYrQJ1dcrM5m0u5sRWOH5CHN0apbP6D94tMZ65jA881fa
nd7AysKVD0q+uGCer/JRWg2R1Wi5J70K9I4dXZkaP8gyQQ7jKMui/oL8PulZfIyS
v55v57VqTjgEwqd3JBPZ1vVKMcNui6CA0iu4WX0OLyZ19IXN8uBNydPGP10WeUzS
xe7DfNPkuN/vhg0NMbRxXuBh9av29UO+jL6BJwwbTl/od/ulwND9f2NA0JYhChn6
9HKOxpBVQ4+vRXWcLftPID1LG4mGARenAsihavmgSuwobn5eJJZWpGEAWqjdDufd
CqjEmIc6TxswTcWe7/NdWtPH9PDmnh2NtJVYfNPqSooN6szbaxJi27crtDCwo6XS
GMWdeeoZKbKZgYAH71V7Fi5nLSMaM4ox8YuSz02CoI+hO8fKrnX4PVhGymW6bc5x
8JlnYXPtTpyWenM13vYlcDJhBtJaa+6xPdV9g15tD+VeTrK2TgnETyFPRIB5dPnj
UvefkUSBO6M2IUB7mqedaWoAcHxUerUwFkff4/YyxZLQD3rCKThKR+bfQItcICzP
W/ylUwdPL5X0j+xGqzFSDsmMX/lQcapCxlKJgNi5DCwAgh0NJVcEHo1DjObUau5G
BrgvWxjbnDx5a3YYldej8Slc8HOIeG6ic3r7qflIO4J9FvayIYVOtA6AIqDyEYNf
4UHKGvSvqEBQTJ+HrHjxySuZEtUd4KEbVeMeu/IAqXnLRrFLbT1T1HCqhsni8U0u
MJ/m4I3bGQCDZ/Hsurl0GHarZgown3rPeQXLxxvjrvaDCjYXquOn5UZBelvkv/w3
naHLPnB4nnipdt+GW6xW6j+lTxfo2TpJecStstMqwj4oZztZ5EEjRmTBDGoux7Ol
YYRAQtSpqejL2JXZDG7mhpbv9KMlePw0J0foFvf9H55jqlIMGWexwgcOV+zZxN4T
5LWG1nQxGOU5D5kgDAW56kYRQI6dugZ7BBzrhNkclR2NDUupKiZnOA65qV4LoM6W
ICKbSSB8c/VFe99hLC0wm13i1ej6oephaCTEdXB4HE1Vy7Cmj+m0gibUb171WFbp
QaYrLYZpw7+1uEok4pH1aZXrhyzUgKznyvyIjifhOQMqBaebg0nVfz7wmlD1HSnO
1tAVhzw8VYs6MGStFSrv3hd53p6kjpIzWbFe+zVvn8RgxgY6qWCDYKpB/i3jNahI
rtL4njFbx1MBLEORfDnk0vahZYnhABEbEV4u1Gyvjhm6fs5zFnCgp30dksrF1JGg
5pDc64b64fbnAv0SRNg/cPEfsqcBv83cWt6GwP2QJDQlfzZjsKqsXHrjPHk/igS2
LOpiA5ER0H3kQXCJzPHsSAGb6eMlIXQWPJ2Z6jHsjYqndMIyiVV/vTejy4JYF58H
JdS10f8MVbnVNKMi34iz9PpICjJ+2ADP3u3sVIKGrpJ4ok5NhDqke0SxKlbHECcW
aEJFp5t+2eps6wDu6/WRKP6Gd9JEmydjl9Iq1T19z+ggPJqZFtivByRUMJ8h0O7h
tMH66i9cSv7kBzddWZNXEOBKxBTGQi9ipIVIy4LIV2rksY7LKl84pTutniIIxy2A
cnpwMLxyn8YE4s2+cwEWWSmeuiNd+e5kfq1IpMJzBm6XoCY/oXzFxIglbGGZR5y9
145iLAHcbK0TMEqaS75aGn6f4FNZvl2ChdR9Y/GpL89ZiZiOwSrbeUsoEmKggk5y
c+XZa7q+RE3hGPx3Clmblu9i4TI3RsHKLRJRrKHYmkSAD4QgxstHCbPMJ+RPvg6C
hYB4TYRV/PvZE9CqXgKw8kabEHzKIDs0xdmCJUCQxKOPK6bcOWo8k7Z7wX/1KaHF
so6Y7zExEhqnmp/1N477A6FaRY9rIEZ3PcU1f36Uz2nCChkICIrNSrgsABPz8ezy
RNhM3/e81mA8Ym7j6vByFekiaqRiGOWJ2tBsydj08QZX72WC9mmkXqTwHsdPPs/T
PqerzyR9nGfFS5vldBzh9PBjFnTgs+R43VLi0b7Le0pWkRsj3bKdc5gJRfQJPcgP
g4HaYGF54sBEaAFyr8Oj8PeqfmmHumjw8mPxkZ2ee7SzDRUtQ2z9ycSnmjsVyOnz
wfIcZCuxyn2vOx7zHvB933fFNYXLhcfHZpcr3AffOBoKiN+pknVPDOlbIIgA3soz
cqXVblIwAY+LGqfJCy9isxPS9zRBISewIdVucLdFuvkc7egBMpUd2Y8HJ5uBjIzX
5Pvej2Su+Ejtb3LTdN0t3zEoFp1MlzaDzybnQmn5iF78tlnGRYvM0rXRbqPPfvK8
ssc2jg+oLJRYUgXcb1SZTQHsLW9VDJunpYOFT9lVW4iXUejJZzEROXXm2ER2ruZn
Y4OZoE/ZymyszRqwTs82G1PBXJwHmaKOdZYUSaeY4/gzHDfgFhc1z+hSDpPa+71A
b8uDjR6cyh1rVS5L2ncDTynTfKC0Nk1TBk9zIDe/TTAKN0e3e1rDUFWvFXbYKr8G
ZJ/fMQzd0txkM3GHhpZMrfpawmIKvNU/gIhTJIc8yGmS0PSV5J/WFLTbUtX0jjca
e/qvtY7opEYTn3e3d2fI/2JE6v/kqDQXh52Tj5yU8kXI/8dStvZUGYekRrdaxgfe
UgjXB5C22FBNHrs1MgY3v4UFEFZVW+ejSoGzIdu7qzrPjE2O3L/MlGLHBNjUfzlj
ep51yrLmC3npx4U7ReSk5dcJp0rUGQCfedPVezfie5I6uJbdLt3DMcO/XqP8geC5
qItnNKudGKJiwahoMS3iD66ZT7QHUT47iB7m4rxA7BZ3Xg5hbACVyvfb2n+I1BFx
AH+DBOq8A7dKbY9NOzmqUVA7c5qBgA9R87wfg9b7gkjPHGeZAg9RmlsZLyV1/O8b
JLs/+Fk6Tq2HAcIEmQfMdygUBHPFCoq14Sw0afTXlRxZk5i+9mk4CBJwC34M2oyI
EWoj/1n6KsWBRbLPcrxQpnL+jarv/xcsnLjHgJevtJkni68wTSw2wynCux+OTGJv
b2kSW7WFFsyCOFm8Uz9DhZmxl2FtDGQYHfgkn03BsoyYL5To7jU8RpGx84yjKyGT
VkRhSIHGi3saTOvBmG2MLnTRJJWFrEofEeYNSYw//FSxZpApUhTroMsQd2L404Ra
zqPmz3mrYhwyYDV/h7h1O9m8ogtQaFKWa4l8eO2CrRWuH4ZTLl/dezG41VP9DI2m
zgL0/6xMTYvZijK78YBkNXGr9C8JkUc8+ZPxlVe1k72tQgCbx+xx8GDqDRkzzSvw
vlHle523lrzCNaSjrBJGDBMRLETI+YHME2OH4qWxus1/pAntE/lWO7kEV/K9dqj9
eCMXeIJvB7bmdaCkpJEo715GOFt5TeG0CwN91NYnOw1La1nPJJgom0QoZgiZ8usx
opGGxi+WzzJlp6hLPRgYwbLi/Vy7cZeS68LWEtbPFwrXWR7cAuBNVhkFqirz0SKl
sN1bcU1OMxjqcRdPGz161PUrPHkn/DQ44epP5KaMb5sUHuW8iKGJTq3EmiqR+Kgf
z1AdfiZDSqmQKe0HvqUsX0QEOvHSj/6q+nw0jJ2VdauMcgpwTELlRAijo78oPYpw
0Z2da7cd9H9Mq1twPPb4uwFf96xz6gUWSozFEypZ+8yhucbCzID5tnHflzEmwF2x
W/DHYWu+JYxPFJo3M+9iqvyIo/Vy5QQcGPGTqxdNOdBwJoXfb9AY5RsBzeOeejtr
B23xoGRCyvbzvxOmvaZS/G4h5kxwz3/XQU4/RqMqvXfboy1V3BoNsty2Xt57laeS
5w6qXueOEhuW2U9FwwLezx3LO1iozjXV7ebXI5Ez9VbMWZm3XOZiKO6qFakE2a7/
SQUvP9RmMj/dEzpJbNYlVt4inpN63zdY7weJ0dkWqtsZXLr44GrUP+dXP+Xj+/Lj
V4J9fj9EwWNL3g+qxJNYnZCSFGFN0jiJmourHVej4dZMIqPbsZrq8PhrPsFeOdQP
zumPdnxZt0xHmi3MpplucPVZiUk0P71V0ctSLDoZLhV8iXLJ6m5agXD+sMdbZpJp
s4lvyMgCarZDpP7rKs7EsxdMn0u/9Nn9+EU3krmPuT1W0sMoMTBF+3uYF+OOfvvr
KOzZSEo112cw411QeqZswqL2pFGSINDfLbvVTPrm8rIrefYzn3iOOR/wwX78QLx9
bJYNhKqFXaVT/zL44LNuhoPhZPTg1M018PryjuNRaBj/eh+xa0IpXzq56TQpCnvL
JxgYiskvyrKhmCUnilFp03K1sUGNZFo7XfOFjgfEPTg/q69cnw+Au1Uc6zRo+Lym
xDKM5zpr++MTWUWoFqZVPU0T0GCi7uJlEsNjEbavk0vbBpIDGB7s4ubX9or+RskH
xtuc+45BzSXeKMn+QSppNNPWa/nEPOQEjd2x/dNmTrYo67aktBHvsd60VqAQOh1m
WcajFrepk46dCjaP1kpFyVgTtBuq7/R4gaSpzjbRrAksLz1N7z4mbphrLQY8dCzt
94voObSAw2A8Mvj6ludzihaaCxs3tgIHZGfgVAYr2j2aiwDTfPi6zHqeuMGZRGig
/Ps0G7RAA8aw0W854++fQ1typZFPclxKuKSorrkYbn80FBSWq+F+Xu0gUNExY4km
KRiePVXBG1cFfpdsHBZBEDOua0tm+Sgm994gAPTLN9AtmiruK1OH3QRiuMtdG/O2
FDvEkG3fOi+cc2Glb9Wk0MA8tPXtRSvlvttS92XuXXagHrJjWjrR0ZhmBxy/G1MW
os58m6I5l0nja6zNZ80k1lNuyr+HnAYGv9FDZLS+hBFQlNxlo3PF5UwynZKXKm3V
QruzV8OJuhkpNBh4hlLHkeBlVOxm0Nc05VwQe2wI9oZJW4TsEiiJRxJhISvu+L1E
/a0HGIdes0L5C8DXu5UXfwlcrpCpxBW13ANVTPpzXj7frtuJLaHrZOb2zyGZVJdN
gdzd8alb1Jrkm0/PxIbBl7AFyqQv3CsrB7dKxOStP9VbAHgD1jGGOd8E/vr4UVkp
/pJMbJ3q/vTPablIvyFlH3wEJOu0YAG72YLm4xmkfxqFdBI6SpOP90Ljv0WOzRbb
PNLiKNabhAmM6AqsREJSs6d2OmDL13NoNUG2/XhOAtE0i4i6XlJ1YQ8dO4mgSI5V
DVMKYR55UN9JTK5+zVp0oUd+4y1SXi/qmQHcqwHax/rIoqsbUEZprbeCxC5i/qZI
neb2MGJuDEDurqBZXQwUUIpt65fXZE7xnQLrc3SQdqXNwLiYk3VnrHcn6qDMkhAr
hMZ+yNckDLyfrGxo3YPAR3r6Aa95Y5/eek3Mbyl7ZfWpAtFy/bzssz8zBiuapq7C
ZavntoPLL8Ev5ECV5bbGY4BtS60WKoRiaxSuTP2B4v+aRAjIfwwYFYHAotXAIbHx
2PFUrM24/6wBDIDchNELowEdlB21XOrzREWoWV5TkdTc2MfTddbfeYkWncvfEkbp
G8+1sVfGCbGI38d0OEl8vyGpEJedA8PCmUkpVOIaxh24l6jkL4/2y5dV+fP+4TWi
LK7M8ks/Fo4fLi6Uqy86JED2TePOKmc+tpX0KL7kor6r8IxLhR4QCehGkjuuFIOo
EuXdMVV0j3Clif5yqCyRROj5UCoaF0Vk1e8f/3NyONzS/pYAknPppDPfUtMbhtEM
GyNcjrTLEA0rr5CdPwXpAFdN8V7LAWJVhCSWAAV3EYdxccyKelzx7ZdpCLlTWekY
7wsVTAs9MOGDVt6y5O4/4H5Rm7IGmrZsLPUlXChLrZ60kfNZecwPUpj0UVal1iQE
4FXSjnjmDpmvkLxiFd4C9Ps+clbezJcI66PC5Qaq2H82991T7H09ZXuZPbS33yTb
S3oJ15wpyIqzovmj9krLJjZWylBqtIfqKVGiOc3budF4knO6TvkWNXTuzzg/mCU8
yAfRK29sAVTe5R3o/npsqWgVlsZpjBJyi+a1/Wf9QRQGHUXbkGYtgpEM4ie45eOy
x2oo9hlAzuu79sUV1m7vf6gkZ3n1gjI5/FxKtVfEbSVYWLsQGXGPS1layIEblSa6
130jOysr7LklP82ehXmyrM7LuBcmDwcfKdBRa6YK+CVrhjiR0Nw8od4N2u1m+oyn
GnaIo/bJA+qUrtdQV0Y8Ff3rMwjJz3KvWM0ElpmQoViol2vtWivfxYMigXOASlls
jN9Bci0jDTUte7glBC9H4wdteQrG+9AEXLwG97ipETX35tMBS2TstBH3ohZsdWx1
Q+w6nRaJbYwpCkXcyZWm5zaqGPiWYfSPz8+/zadhgzrbyg3G2bDJlCYl3t/HUTOC
19THtbMrcxMXJ8wFn0A1rttefSO43dcVgeLSCNE/LQ1oNeHlHuLBGnUReHUHwOl5
jXEKm3zdGpuDTAEFbyv1eXH589LlNz+00Ih0tnoAMruZWu+oBfnqvcNkCf9Fn/7t
bjrBE+/u/kOXI4yS9zOuUov8yJnhnJintIwzMq/knES5IhIAsydJW3W8Qoe8dA2W
W9AnvIdRQ+cAruHiiUElvHtH9fx1WPRWX8Vid0Aa+1Wfv1PPCH4oN6OjLu/yBjLn
31ZI+SFI9vxlLYwvkh95PzHjr1xpPL542NWxjtqdhyPVndooTZiNJCT/DdXrUi3M
DaHQ73a8GSeetQI/a1GiYpFGyLtOvovjNV/K8NRsL4D7ycVjsqdc1cNlM+wAPtE9
dJ8kRBh6T9Az8LMHU12iQJiRvuh2Vg5EbYfmFLaiNXJBhkei2zE0bVXkJZJeIeSN
sOGRHn5JO970958K/lyOgwgY/zl8fZp8bzLE4tAbCLF86sDnJM9S9t3FvIKeBaHX
NIO+kEVQrXkkWGoZMZNXmKheA5396jhHp2J1CtzPaZSBSnd/cSOb0XJ/O8Z5VmCR
oulFULlYpqpWN0pqOlW/eD+sYvd12pp/qDqoWLq6D5aB/GTWDSbDXlMfDCmFlTLL
+9eDvuDqG3/Ro8iepHCUkESxeZHEE1vil+hBE8+E/mAOReAvdDS5W4s2u+oaqEQ1
aSoVhPkpERlnFRUJAIHRdfOhniUZu8GVa9bIIFUYEFq32o8QFiWG2vn2hEo143UV
9BeAv1yRHTyu9LMF1Pmxv3fnwz8Jd7EaudDFwYP+twCQ/8RJPq7gf9TsRVInnLSQ
h7/E36Dy3uF4ihS73vaVSaJ8eVeYleEzWiQgcZ76cEpCm8kB6Apbo315aOgvua9+
VRGYudu6NcG+DITKJhXG+fRhGau1aE1HnNcQviF1Fn1RXEZ0Ip/5U/52ya6L2sEI
gjKMuLxFITAsvCmVIBNdFSjeDzqLg9QqaI3Hr20wjZDYGclBbasY+uP2rEJHDmrC
ctv+OMA+0Sfy4mDGiA84hn/51QW3E3ujZGxAwQkIYJAWs9iyxJzjcKGJ3ozNHDN2
ThUN9afGCXgi/zPJGhrmEpgpY+nx+bMpCVW43Pb5xmZIgpWRGhE5rqs8H0kG53Qw
AOOfpXofjztHPsbZXZCprgf65i/tS00bCSXPMQWXsKdyT5j+1VYoeDqhUbqpJvEh
3DZtGvj1xzxhCb+uV+kucS9zdln0AJFiLTYN7CM/e/Rah0Gpg8PJgKZkRwTWsPQf
yboQAYaqA28KHEkp6xE16eWiK1aaSbn3KEJv11ukSz1WSGgu5UtCITBat/wU/+uy
0AlChtZU7od+WJiLKzsWkk0xVkEjbtOuiAmMzHGSERqKZYzqsPL4MIcs5if1iidA
+KpxssIvpDDF8AjeJh9eO22kyyfQ4GYD0o+1f367ZZkHwibL366pfpSY/jfYozDa
wABC38YHjbr5Q7tz5u6IHYfX3V0r4EkwIqIB7IH2RYPYPraJ8ElgSOKGtd9QzVtR
NUzrnYctwiYOEK45j09UcFXuPuxK+0jJ2eSn8vW4nvUerGcppChL/X592tFSyrkA
mIZgvkfndK+n3VsSEIa8F5vY5B4DRUsmASL/tXl3EF3fgkjoRUIbwxGE+8zDK+uG
Pxia8sUlkRY0ISVseHSRk3YEuzqFkQZkrDltW6KWRisTSqgz+Nm7TO6Vqbu+0nrX
pao+lFVm5Ueiv2d4DJqn21zbAU13QJwI+PPQqyuFNiTXVN0dC7KG3m7Lg1NdnT6M
livRmwiGyj/09cMU+TsHii7S1uBVWT7tiBgOzZztKl33ZsNTs2iD2P273K0b+kHm
qxEG8DPQexuui3gksdRmBKxQM6FgcGnhwG0CYgDvKn99uRp2SBQu5iYYGjOPSS0x
/UiJaM5W5fGFyxktOZLIrVPYMYYxZ2w82THPRnifmGTlk+46Rg42y/0pFlEi90C/
8V+BYR5gRXhRGzmd8bVNRTP+Ac6mMsM4soruOOuNLZsBdANN+gXX2yW4H+BMlWs7
LiTK6teUC512mAVOKwMzQ3uy8Z3OHxAHqCJfVZE334iG3EGDIHOxroyDiWnjAeKx
w+Gbgchj6OvT0lC6divAnjcOOdy6bZgLsuCAyVmZjcy3m6fvIv2zP1yT6NHp45Z+
QLR2w/XPkylNvNLMwYJki6DskBcehwCqtvXLp1nrm8Dsj8fVJL4JQjwJf5S0Ne2T
ENZkNbxIrOfmrZKjLsfaQXRNF2BufnCfxnf452RtJQdUoAKYapU1ZkWLqqWbZlC0
gvOVekbi5tAKlGRy81uNLJARF8Q72PtdSqeZA6xjJiKChGEC2om9hkfG6MXkhzk5
BptBu16R2wX20FulNRrScPRME6JnaCTLUgd1n3Vw6Vx3XJExwpbPLJYusrbXPLDl
THH0z4HFcpQL7DrkdCPwLbEZ5rk0LymIOb5sZsCfnwkjyV9WZk0qfVnyqBzc5dOi
or8rrcrSl4n9y8y1wEfTn/P7xX3zO78wryjZgXbIyIcubZhW740qGgdQ/au+opLV
cPmlc/YzBgvhWlz4MA6RFAnQ6/JZz5wUD1ZEu1BWC1Q4g7kxnIOWkjerDyTILbID
0CApQ56oOJSwwhFP9HjBzUJOS5ZnE+Jx6M2ACTkWvPLLtlrKSTSYZZ4gT+GhUuDN
lAB5pTj0p1MnkwPa32tvPb5h3k425et1zehvII5LHB5ZYTegNOtSn/2PAsiyBDDp
KLxSCPpMiH4eHte5oLMiNTb/TOO8cpqVicf9wwDVWGoNnrP+pe/h17poAqIdRqk1
WlIREj6VldZUcURUSU+M8drZdjZ9a/zUzJxq74Whnl1JT6DrhYf4vWtO34YT6qH+
M7dEZAxQBTK7Nhxgv5kB8kMsOYgbJ2zu5kiXmo472FDEFs1F9S8aqnTQYAw/GG0V
kCuacP860bh277S7G7t7uy3oUfYbmRce421baexmzYtQVGG2sMJxLUP36b+eUNhp
15OZLwSmke1M4/RuaPJsuDEUMByDs4auJ8ATJhyYE6UrsGWV4zFVW/232M7QWt9D
gcSBt4NmfkzgcmSXgvf7EBctoCoqcuCuGDl3NJPuaOVrZ2JvaKSS0yhFen6T8MeS
53I2vdjAT/QOe76Avwqavl0P2iIL0Zw2u9psPAkFyvrUc4aWV1qFwHhUXW8XAFfZ
lf5kbhmlJ2BGCtT4oBlBQkNVITUbMKP7rF4tTRKmZXOv14IqXE/y7qEEmGE0w1Y0
T6AGEm62vJOzbSQwAOgoNynOhoEf5jpbXjCIadq7KVLrb1JwpmXH/hSRzkYIEiLq
w2vFlGvipRJ84HJma4Pz00CoByGh/WQER/zH+JthRGK6A28GQAj34Z7b6jayJcVs
dGaxjeW5EXRmZefCSFDFHkVVfCibJDWC6GCkDpCglgPyVYunfKy3Ah0ucE6phgBJ
mdat/vrjUGZ1ZhCn7KtzgANFlFTp76ZID5e2QBN2+ZeqJknSPH07d2V3fpPhvC33
v7KjXc6Y0LE05MNy1f794DRI9f9Pzs2hzFfWtnpWka1kC7doKNQKAsTLxyx9OtSs
Bu9dUr3X+7jPlpS0RXY2IdEuXQaunCCXDcjSMbcS/f8oA8YHPkjZN65p4hjFGkDb
gcGpljHkerwlkzsrSsk/7Tzouu4MU18woKk8M4jypf8IjN6yi0Aw4Luv2X6RcRng
60MUFcj9uhy7V/QLfkpIWwCF9jXudeL1Lx4T+E4TeTaJKiYZd97QA3EetjDBI8uJ
joRkZuI2AHh1YrODQPo8AOrFW2n1ktBM9QuN79fex0m6dHLezPAaNciPClDbnyrY
jfMZSzYSkPIvMoOndT3H2xhKgK6u7dzhSU9D/IVx6g+bDIQNe6+XoTy68INIOJJ7
lLWKJ9iS+gRUmSRHavOT/mhHhn4SuToAyDgCkEvvZ904zaK0QalRyO2bzLYEzYzi
AVzNsWlsxJv6B/T9X1ulJ6FdeoaAYk20V+TXCfjwUyFAo1VAwsm0rp59smzGPBmE
gyAHazj4MKrfw4IOcilayhxrRz+6tP4vazSroudmwFm2m9QYaXLLr1B1EZvJRe72
j0x67ZXp+0teVwCk/0LK77IekTN1jrci9HMjQPwDZyISDmAeru2gQsbVl4Ut5tzY
F7AV0M7RMT1G5wcOL5cbTjMFItGiKq+32aVME5tcvEIl6ux3X5qChmnBZI7+i5zY
5RV+anQuJY4Oaw+pUBGAGU5gvUVx22mUmEtBiHmYhAoZFd1abW77LmihFK2OrXva
Vl4+sABQJmYyq8OanHRRDl1EmAVHEQsB7JHzUk8JPzquHKgzbWlbFajGC2FeMmeG
W1zCPMBmeSDNVLeBdcMH+NjEyJ8ggjEvqHlMGuIg7ngNh3tbvYeJB6TTnGTjci3b
diIur7u7X35ETg4JOGdEK5OiDPkMeYEwmMSl8425ptUFQYHCI9Jw1Dp2l5MGopYw
L0Lv4y8Ags+ImCaa6DhKed3QtzObuJD5Qn5nTaEWj0TqR28DpEywXO73Fv2RttUc
Op01rHfbfoM0UOW0xInQYKKlfGIAy8kQaImFwAgGN9sF5dGnoSIp0ltYL6++G8pb
Suv3SRGkL1awNEUxXzs15fX0MqkeedrNZG8EsXupwee3Wco31Q9d+0uDDRIWGF6L
99Y3HyA7Q7MXnv1iL26F2jYuW9Hl8kEYVEbOjYxONwH17buiHqlyNDeXuZlk1GBR
pRiK00w/aJ2W6gUz5sOTgPXhB/Xj59RoQRjnBpo8DNZJkAALd0jOTpP8b4PoOP1c
os0qPv5PD1nj4/w/qgUgYmLwHZbEnVeUfuPGWsj5EEnWCNo+7FTZwLpy+JzO+ZOj
l5JbIcFctsfCe4K4uAk/xSTo2iyFWxEDWftLhMNWwTEShsOOULBzz/QX7kNmXMrF
jIfsfxxfauZA1WhSpX4ATdtkKxKnlp7B0vCOVQ0l/j8Jfgo6BlsXb4pIGCj9H1ow
h97PN9TF8K6t4CuKj8ghimxwbaSOVMsPBIonJpyME101U1mXdqtV2rZ4RSimo6H+
hSBdwqhSKjfpJwT4YyneFWjsF6/lu4/cH0SnrhqcZKmp8cqQLy2F6xa9AMRexg/J
Dm1NAAW4PG/Hx+MWCarNgzVgYOO52r1X/6T5hHFYLXi+K8kE/VX1wDG8UXNco/gd
66mxZWRfJ3ZxpwJjcFHxBXPDzFzlKjcMc3cATmx9A73gmTqK0iDeW1tkgKfD/wEK
WMFk0qoZor8LozC4QcgJ+LxTBsvWsBB7zdPkeIV46SUbnqmmlCjnLfGC65QJAYIl
e7tWwrEOEkkHsHksyWI9OoeeVZPd7QNPwEqlbgu3Ckr3NePCcGW7f08+SxEr5qdT
ExsoGjZF/c8JZk7CYWKfDGxN6CBzpHY7j8w7fo15M+/S3uA+CEZIZfmQCP7A+Yc+
A+esHP/gZ6LHtRPmATRqIi1zj5qKZ/Zi1/82jiba4ZFr5O0KqSwvLqLHYyM4loFu
u0AigjZruhvllLfvqzsHz+DL1ozf3gyyrNbdrZu1EnrDDwSfbCC0I6HhvVbQRZaI
zpimqWixnBKjgS3GNzDE3iVwXT73f2D1AiVbzGvg79qk1RphuslQs/LOM2+dty9w
wrEXRSyDEa1pFFohZBiu1U94hUu/CxHZrmfQ8Wugc+YpJqMEkfaZIku2R1oFrNmI
viYCJiLUlK77mNGBdx8DkujdWSLF+4MSAZtxTnS5PQXU3VTgMqx2KY46m41iQhRK
EuDEDTSONE/W7tweePjIy6pVGwlOobnWA54HRO2AclkMqRCUTJ/V5DlsLZVMhb/9
kKOjR/lSNOLIVUNFzI0HNvrixWXiE/RM4XlzxhQH//jTsB7tEmcifNjCy6muHbj9
WLlAjCntpK9vQ1S2aiDAvt/HCwQ4uoAZ9/8A4dYJ3Gudd00pUrv1h3NmW3hpMrBr
5AdXRO+mexxEgrmhQJoRVPl1IKtgUHaJmvBUv54eYFJwkUHN9J2ZoQeoivC54PkW
v2AvYpwZMo0mGfysCneXybdSCl1eaxmMjz0+dkjt+coROTWrM5m2U5h/x+sEVAQ8
qrixQV0PxY8LdE0xFabLKbTkcjxioTtxwDDmDmWTYAkBEaasRzULQ2ELq9dZMOtx
1oXeKgwnRtvhgm8i61ly+EcPiJL//pHuRqaVp7ujv8u7dSw7hWUp3tIoRyIgGNdi
9V51S1oWFO926WZC+PWGMWhFwwKeThDKsGzwcLDElOPCQusN2TGD/SfeTLNnnCoZ
Elkzw1n0QfYkiE4G53utFMQ+N51rgtvAmyBb96JeR1nGZkOW8+eH+PXd0sUXMPuw
Hl2ADT1uA2hrt3B5zL4EgVknhn2VilZ9YollFEF6iFGCnN/yDf2PaG9CXkb1/G1o
/ljr6It54Hu2OQrDiie9YL+Qj2av1rN18Qt3R6VQOEMqmoBk9rW5vG6qqzFtdoN0
ayL4PkNtk10iGuVq/Nelhpkl4HMWYyQa6Fuo4yyCs5DCEQBfzSdaI6cROwFvosgB
Bf8GY88M+9mdTzGMv2SgvTJYf3TSyu1yM6JLh265rJ5BKy+JoClYW+fotBEARqHa
rtlfs0ouPVKaZWWyevzcplB9Vng7XbR0TquEBAMiOOYjpmbN2q5i2TWH5c9hrqqe
VRfaZEd/lmYnBFMQb4/wMd/I3gHxjoW951lIU1Hk4/bOnAPwt2TdEaYxyFrME1sN
zkGVe8J+KGF6ymfnYwZu+rZufjfyI++bS5P9BIGymMUp9y9MmRQghgHNep6Qupm3
VjYOisNCt+tgAI/tT9TSbkkpgp+DedT8BHxCQuSGcyMo/8RSbkWMgrYXX5/WR6ut
xJVr8eE/PmHE6aVIvKygrqPOYFszpe1Tt2iTqt/APKFNgoygOjmtii3AnG9DpFvm
yaBuLa2OFl7aIdsSBwOGora7QNgvzI2H8SdxDOzOHHZFNs6+HEEef6S06jubc8cv
zr8worPaA60P/MsQ2hD/sdXW1RgXthkzbi+ubEi+Nr0H41TSfH5IyByJI14j6V64
y2aXzWnsqcSlzvIE4MiZJP5Gis42MrGBO4WenoL8Og5Sc1AbGCXcnR1aQm6d9BnX
SVYSglRI01TtVq5GbxEfItEj70NDYdaivpsLdHjb+Q/KJjOLggZMQEpfmwA1vRHv
aOn5HCKx9dIHmtmTBRB3edGO+vwoVDpVFO3LmXMoZYCw9lw2vvyFjFN7uPBIRdUd
qRvxtDHPsJE5fnwxjrP8igvwlH2FWFhLP/XExQ9UxAbl7s0CnY3AczKWXypjIBgG
Yy7sEYFVn/KKV3S8mVL/FsBzOo1aEhRBiYSJttGCy0axyahmoqLT9gPJdcG2Shiw
tgFbjJ9KBxmqseCXi7Ny5WWdGjNo6tfSgywFJenOqT05e5SOGByQM7E/4+QwJXTB
eDgHOtXz59yLyHA2q6zBlcxzklgQ+Rb5u6y1oak2vsYy0X9bBfTM4FBYZ2isGRU+
uc+q4OYlyjfrilt9DpLY0FG1AfBYDV1Hqi7tnAcI2Pd0kdcpLbvPo1ZAlPl4Nrl4
FcKv4IyIa+AoYwqe59bUEXxAbbjL81xoEIL4gK0wdmP2Yefj6DFFPEw2D63ol6Ts
iKXpL3L1kbB/rDXfvHZLupt0Y1YFyuB8si7sAOLxrhuGQ1kNtdVFakQ4f21VRf/J
wn03Ql/l/M28mibqCp4KxDJPVg3+zlgIEBUdweczFJP29xKBNE86oKolz9aLmDN6
T4TmGGxUBYQWAvtvLGFYMjzJSA++i0JzaY/ir/sLzb+HdH+FSTtpAhhuhmnw+/79
48vo10jrrJmdJHB7gtGszXB01bDSQuBzIiu6w+O+n3SNAruz0LmXEGRJA2H8d3u8
J9Y7MlBv+PChHf6pjROIV7YyRzSG3/coIwLo/4AHDTnWO5xKJLgPZuk4+1BgtYZp
e4yqfLUe/eGyeLMu1xs4PfUxkhSv8DKL6KkuJXokHfDpVdAdV+sNaPXD78u/uGpq
5rIQim6GQ0OE+xC0hwr5ZTfmKoIDsnPE/e2r5OuzhlN8VtsmRDQN9CHAU3yFYMut
CXKJKkBH9Z97jU3gnDH54iM3BYMf9aeCrk3VXrBlcZy0GqVQ+2SCf3QUvhiNjJ2A
CyFf9/h2OGR8ilLHl87PR+b2YZW/H15PThJxV4DwgIR+ooMJ0yVdqoklrG/I8TfK
fajz4NNM+inReLFbkwwuUuwrlY1oq0OencfG98mn6YCxSSoJpQjQqQGn5HjWYig5
KY4nnEpKFlVD0KO+on2ijx/fHeE1a7uuN1bnGkWAcmzX0toWQIjG3Rlkn9CH56VC
qAh+hDPekgtsR6f43oSSpP1LagGm2HXUL0fvRJ5B2cg6qan8AQT8hb9yqG47esPM
rJudfuOgpT1Z60Q1mBKfmP/2mffvUyj49zuMHtupGUaSF9H4KZpLOrtmSDDbDv22
CwclCUa4+Aw2J680CBydeSZvWFCW1kwm2JY9uSfqYaVqVjC0QC6Q79m2ICT5Qo6R
4jwxet+VgDt9VFl1MLkIRlsKMM7imcPrEk9bvq5n0hPu+wjxM4ifJCxbUzjb95ST
t2NJiyBiO+Y82wRFPSgXl9h7kq0iooGdqaXfFKp7OUJRpHkC7KBoESmH+2WUbkNB
aB+KJMnic/p3jlTw+/0zcBSy46vGoxRhYlxnAAr1ud902nz02mAi5Q+u5MaXUSKI
+FZpu6uK3EZq6tQ2cb6DocJ3b3a9ELWdHwFzTE2ymuybXcJzU6PlWhdegTCsL7vr
IerT/YE2YQxNPInonumHEHHOM/ozQTokU3/w/u9m4oLW+2T9jcPUT2COAvlZOhkc
b1oC+0VP8CWDXpNartmHg+fXGLRbnOwkT1F11O92btKuRCBN5Z272f2n1+wXcU2i
s00Z/Xuyl6UhQ5NKHs3G1313pjAv18Y89NUGBZbsI4H4mtKXLEIz1sE1V2D9h5Rw
dA8CAkR+rb3UlM0JL9nkIJLdBXC+yUiBPtkREtC8btR5pkC0W8RHZYhJ/0pH3zio
`protect end_protected