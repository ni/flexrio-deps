`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5408 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
e7odJ6CQvoTnAodZnpyuDJNV6PMjKoaz5XVnou4CiCtRaI0S5FntwioAUOPSMkFV
4ACXEUrjiirl7mX2oQNZpPWVDv7YbBOD8S0Axpf/RFTTrWSv1fDSnCwlB6MkLo5A
O5RLbDUBEaqwCsK1ZeINruS/3XxEmeP6zLQgnOtxMab/5TTAkH3/et+qf0KWb1H6
5sY6t5Ygx5G7fdjMWS4ymq6Ndn5t4BPsUSNThfK7TWz1dB2oYEv8U776E1pz/LM5
lFAPhDPXxDMqY7/Ge+5UPRw58pox35txCWubm99hZGRiPdYQ9tvUSh3J+bHy63rd
6P9cNIFX4f4w4rhzSwUOj+A8nz1qeKKsnLyxzQUxD4JWL+fiFQ+kP/LiB6NkaFef
5BNALGluuBVrFfxqK9SyMATvyukAg7s59pfdbMpsMK7S1o3L2qYOLkpZ873TjO+b
s4gHJGXgoBAVgRbci1PKgwg2mFn1Jn+zBEwXMujIRyyi3QuZfy/6sAkuTdvWiWf0
732fFPB1yW5LoGHqXHRrRyxz5HGvIN0QXQgvGYLkynJ0d6PsCloCyuTmtDt0gZal
ZE06PBx3REQklNFKwno86Jkrm63slTiuNpAT9HvG2JwCG49wNn4KWc3wV3aWGbn4
zU/ZIck4EnjaEYhhCnDwNNhaO2DcUAK1iOLlus8DIYKRWbQZ3ngu9H6oU0JH2zmx
bNg19T5JewTSiiuMwcWZ7NmhklUfTCx+dmixVkYXs1A1pR1wkRizldi1jtpJxcR6
Ku4yRIzh+c41HSXI7GPBYWY13ryI3w4GAV2IW2hYkL8eA0Zixjh1dSn9hlFJ1xT9
YCmJdwXqokbZfzJ3pfwQL/KFxEDhXrJQTAm1+3y/KVotGI3EIzmqwsRmHFiK8XTR
l42Mltyj6PM5qWI7R1FGFu4ZSGd0jm07gpfIenVrfbHjKa1x89yqePWPS6sR2Vh8
un4I0Kyac5mCN1kJVaTEFIangU1WYpo+xuPh2PdH+7FyWwqn3Gj3p7j6jxND/xur
x1NH7B1tkWcRYFyZzdoAmC3C6khEKg92alsrIioHqFgw6GJ2N+ZWq6frAxNrVmWY
Dl5riZ3Heb3i+mY+96Z0S5AwGFfL3WgjsbVhtCPKdBQ2uHbJ70E45sDXN9rjbgf/
iPzxeLo/GYWco2J6N5o2SVSx54unifpNVa3LNzXPT1V44SdBuW4T23UXM7y8w/s2
QdhSkLkM4Ln8uNx4lqQOxY5GeyzgyW+IPvfyL8GOG8P5tDujmGxZkx4Qcl79/BOq
lcysGod9EBHSa4yLuj7VKorSf2ftXr37IGzJ+J76MXXz/sc/JgJaUcKOotq74Igk
HdIUF4OucBgUCZr6v1HzeQoadcmv/NhkqmoCaN1ks3dGrTYmBhVCEqIkB0WEy0sO
fGLLaXffMJ4c8liZF4jUrifWgGujp11i8cgV4fKPiQlHVDEXM/KY30Lz9ZEfF7OZ
5q6XnnUStfqog1ml5xn/bBxRaO4gCXoa9GxvqYdLAK1B+uW4U6zaPRRcqYGu3zi/
0ReoE8F6cWtkITtoFHA5fzmQp+Xxw88ZdrAcn8hPENDh2DFm8PJwh90BQQ/tt/At
S08vLzA9ls5V+T0U+efrbL4xy/bCKfsQlM65KVib4vT3sY+zwvj39NEZkMELmTAy
82u7/yd4hd+goyBcCfPAV931xxLtGUEN7rlA66ecO+GTS12ghYiBQwjKtBCeyVbh
ztWiik2ypf99tdqs/t+9kssy/bx4HJLB8I7srQVE7sL0S0L2zyvUcnP1pYOsM+Dc
S11v4hcOQlA3uQlJ5TGyulM98k2T9YQVx9BJ0ikGgnN7KVp0xdpGb3d4BhMw1Wp7
n7Swv311nUMEXwAIAZgy88Xi3plkOw2llJm5ywV1NvcQp00BusE+N1Mc7PtXeZwE
2/Fth5RN/QFLDw+yi59TEpG/h3/e07/QK4spKDuOYntt/kdj1ZdSshpJZuerOEcl
tswZXMfDKlN/uUdo+zURXUP0nSxoMBgKvajYT/GvPvYbX9P/L4TVGAZnnSGGJeA3
htk0V49+qOkrHY8SGgoXAvHb0mseBlS6lksgqOK1KpvY39bcbzMR0P8o1XG0Vo/q
zYMreATFqW/YG9z9bTzaNCTrZW922Nl5Bv+PAuVi08NK0x8xuCtjLml0Zms3N9A7
r0DpEFrmBaF++foFmziogHnBlHRBqgjSqQB+KlozqBNXX1lZfLHRdVIF+8vRicN+
HpdC8CA2o6QdSBMoaSD304l5qERbyt4RZG/WBcfFyNVHlBYD1Bl74JTD2105uXK1
+k7+NrSTYQMMiMjg/Pa/5xcyCV2y9HUOVh7IuQUkhxAdBpf7ag6EVQYMNr0d9qVA
DKqPFkM/0Qe8ZgN1SDr1N50W7XDauiSq9pyoBIax82E73RNKA7nsUKwv9F+lWlP9
qKXsQOsUSOaPwHimSbcEezGcdKyy0yf3QA5oAWqibDRxslqGuaw/7B27S+LhoGjX
p1lcZEtc17MKmu/qrSijq7RD3jc/KPnenXdGtoBHmNeJVewnMG+hc2EoKhUkoRvV
7i5TbvhqEOiy/kx4yXfz/3/RMObtyn3lFGMnH69IZgaW/EtGx/mGqntuaVU1ciry
bzFXgZwxsclaBuJL3N1Wlzk4YJEDBuq2KTXvqc/IlKMzJPOiGYRdezuht502gHIV
RLLfkIc6T2AtGN2EuUKq8xBjmNxA8Z8BmY12SO5V006hax02plSX9zYiKmh4yzYq
zGhAWWS+K+YHz2d2XehK5thTzJg2IxYxepyji298y2Q2tlxrQBkHR788hebQz6Or
eBtdPN3BZkxQlC9VcGLELiO6GHuLgX5ex/RayVUyueiez1M9TEVGb8+ciexjc76s
GHN6rrvx3wQDpjsHAmS/zO9YVLRfL6PCmJKPgmrXdGG2r/KuqXwjSWmffXyFmiZK
V8eUj71577OpkVtihinnzayN9PR1KA25iXz3GWN3YY3xPB3jx8gycEHmeFk9hkUj
IbhromAYdGWLyJmw1Etcsj3AAm03UIy0ejAu5Cf3cI2DP8AKj7t9jzZZvbKookx+
eAt+aLJxeO5l0O+meuUV+v1CI6cYxpdyb+DR0tsM2d+As94DqTq0Fn2cOE/VO4XD
ciIX3hbvWXCAwBFwlHSV6V/EGPUZldGIYIt0IhSPgH62PoS6Up3Z2DPTcxvg/Ia4
zTrlQrlr0QsbLI+YdUOShJlhR/RL05DD8OxMDfRNH2c6XY6OMHTu0ykMxMZZY9zz
J/b83lovnx+KwC3fbAkn87WUC/qvjjaAdiV3ziE43WUOAFFe52Gay7vFU1TBDzP8
6eytzfU1CYKi5s+zqPTxo2eyIgc7JBiFB/VH2Yxyn8rOmQpGscAXawHbKP+HT1vH
eTC2AOc9PkM+xV/OzSAd0Mxa3KPyUNTq74aoEX9V6ECAzFq6YIXhKCNxqZTAWkcA
yjpIGDOlmX5P/DIlF4yIzgNDmpbMdawAYFJ280aME31s4ey2aeo83ZBz9mTY3g2t
cvrncyqcHT6lThG4hTV1W39MElfNjp7gLBWq9ntS8q8J6MKexTT9uXucKajCUSxC
aFgGVgTx5EJ4ncQqvGaZg75y3W/39TN1k40wpKhwo4KtpiExVRma90xNsnA4NAVI
uDld97GTEEyZ+nOpUuQSNAdJpz/fO5XscWM8+KORXfh9bdHIgGYKN911rDh6fjUv
qsoamPU9/ZvbVhsR7qrAk4iJVEvUrya2tEZJQ+08NNXgBBp2HLmreRXLsj1FCneU
a+os0z/8bo/0Hn7W56R2lmPA6i2PJhKJqNBwpB4MOlaGNs+gZPpjfjhH8bcFAnTA
/6d4vvBiL+5rcj01a5aEONvb4pBNgoBbKXvgUwWsg4oH5ojl2TTvDT1X/LfhG8oz
C/iGXYqKMtHJEGQfMmNWXKcT5etRauzfi31JKEE+7vVbSHN6JstZcpah/MB45cqR
qV3g60bJwoUAu2qMtjg9EWJn9gcgq/gBckPtHylvMnBh2DprSVZUz9oLRtNnoiSR
AWg8Zxa8PYLlTZ98mF6GHYmbYqyD63kkGqR7JLDlJsT+akgG7bBByfxzCpL4h4ur
by7pXk+GdOz90jz3Glko9gTwHurmR8worUNcznsZ/0SOHrFJqO/LoCQtnz/lfmps
9R4HFzCl7zWUamTjUYtk38z35LhdxxicHsOjfDCuY5d6t2+H7h6oNY3PW/u+1frp
1JIinb+aEe8MHhncsn2u7WECcgH/UyxNJ4I54a2QHr1G5Fm+Sx3nRhtKVotiMIYf
XZpDKQpLp+y5IwW417JDxqDFA0VedUDTaarRbMLuvHy4Xk+rGxot1DxmTWYle0VJ
hZbm+CaLnrN2w1iqLelZtv41VKNgiK7bzq2icz0rckLbl4k/2Zhi5DWWuM1JKutx
IriQ29dzPDqCBpAgGVTD6PJck6YqsFgZuxUhagLg+iUL0diGNR7QzUX8MZCBAoXJ
GWG9Dlj8tHXpG2MmB01AVUJ/IpW2Je50se6xfWjVQxAeXtyH7T9qg3GUuS1OVE2g
ltqTzb6R/t8GkYBxWI/xURi8+TqIUSz0+lDbsTMEfh8DiwpiUyTsoiH+uSL6D8f1
/o8l9q4UKf+zrh/ZlRKVVJISFHzC8fyIOlM62OEKeJoESu5lHTa9J4wkDDVAK4up
SAjF5Kkkd8P3qDu9ypJHhy0WbsuGEAWtonIJcyFyJN0HFMcMk54fOiBJzgyFxx1V
aQ2b83xHuQUV31BnBIZeif0geojXvrU5i2CF8ohDfelyxiSX4Ika04LfXYx6OqPL
hGNtHZw4pvcnyp8RL057/L28lsC2fWY5P5vnNI4sqvsjfkqCMlocicsyHxNLbtSQ
iLLZ/nTIkKH+B17bbsbH7x4/kWM3wEi1YxvVLMoSRPaNU7xBp8ref/hnRqbKBbIo
EvQeKCk456Gm9+0F7+bcEXi/SNZMf0UrlypNBTGt7BDVioR6SYFjxRTU9aFJ1Q4n
kR8wbrH727/hP1KqCZd4C02x19znvchKPXOGdV6KzgtyKE5QvluvUojYpU3EFFuL
YQyGM/SithOA9FUgj8axqvY5deDfhI6mSp5NbKYWkcFcAqh+SHjvreTV/0Bo8kSI
O5NZVziUGqtxdZKNR/GUsbEV8U5CY5l56gBhEkAkzMuQL94NuyeiXdCQvj0ilotm
W7KOACehIJqKrBXBhwa5DuJzOJ72sRKl80pLpHagMGermleWVsQZhyljaBEUwZb+
UxvYZfnQvcew2xszfblWkH03UK3OVZU2jxlxRVLakEdZUUohFnzuh4m24kChqK8T
uURxBnN57oOvhAEYzbqifKAxuFamZ1STaz29CP/tug72y5RMFWCfXDcooM2r+Jmn
dCls1pxK2XUJwCptBouoYOTDO+NoBWsDJzHin068h2/5cdvFGfDwWRcnGeqCB/sp
zAO5NASMPbUnTH/0CCscRyvgFn1N9jPrDUo0Ht1KhMmPBej7RNy/T9/6TX9nxORc
QjmIEbO2qL/y3WRp83rKlK9ZmLGI0oZIejfR37m/IKZFkTQPE0Zx78tuZGVdMFNS
9/wNmDVVGP4hJiKUQWJkAWsM1koWP0dBzTZl2Az7QidBZvuCHlapcXkX97IpbRbd
7bebFPfZA3QkmNPeS5dZ7Ng5s5B+b/TlrTNhuVl09NsQe+YLWBtIpFn8FThkkqnN
GdcSEgrGKat7hixHuu2kq3Eug8IjE9JzLciEN5hpuZ5B5kqNShnDYKl8DpnFbeQD
aO1YOHaF/2NWJ06J3SYd+6eyDFS7t7dwGWhHrqtG7aIG3eBiEkZ9LzQ8XELGTawu
5fmKrGsinq1lhc+GQmxv8gRmPbEo1zx0qx4R+YsEVCWVWHoKK2pjk5klI0zC3Wm7
KIFNfaV4LyXGgMI0ZOUj1gLohzWYRQ4Ce3liLnky6IJ2HbIfjUjX1Ij9CgOubQsA
In0gF38UWdXPCaHFyphJLvI5OdFKREVa19FTwWepDnwPwVedi0SVnuOD7/1qQPSQ
vsJZbGwoSxWet0F+Fm2h+uD4DNORVY+UM9HxffrovVcMZ8hAJyylR2n2qb6s2TCA
qZUO+M3TwHAlclZI8+EDTm7d9PeXJtwPzeEaZXrtTElcgUx6aAsfLO74gQKkAWwo
q6A7aahIvN1Ll3P8caQ/EUZbCgeviFY2yPE45y/D2CpAPGiVYG34SbWHR7oNCGyI
3oITTgFK+yFSeuTcuvas/oCBpXNaqRRLHWwig8TyLNsCNm4jz+vQHua7Qv/lKNk2
4yD+3tq3WWvBnFGEXBpAojv6tfyDKQuRzbEbnh3qhM5JSo4isx8MfmRlcugLoA4y
xC5Rg94LxqSj0OO1g466WhwMYw6hVWWNhCdOvQAPM8T0fbYKYdJ7qBQyBcIrxUyH
44nHUP3SqKaoeOgIgOAh/aFRS/0XaOGxoj1GbhDMbUilgNk6I34Cx8B8Vn4nnPYS
3WbFj7aKEboeT8CdO+Qsf3KDalNjJq81UeItpT+SaDiQ/863IORjCH/UhH4a3/N2
NQwg7DX989LbdQT1oKNsvKSxdCGIB81/S6mrrgF+OgUHSTBBF0LLalFiLwyJM8DK
2lxGACcyEpPdvtfUy1yhNSY0d/CfRV9GEMSItcZ2k1hUk24pAXjuPu1GxOodZQcG
K5AVno/hf/ShkstJz209TspPlNeyWkOz9qtQvDKUpMOrMKQokukfXOL21X5gMcmS
vkJwCvSTnrF5ziOIlDfCnGkeftzbk+9XqpsUR58HJ57r/Y7edZRpoYWpTO/PFO72
3UaAdELfw6vNmQ58oQSK6qngUFcl1m5ZNxfqp894K4lmc96dnzjBuVHiBHmRuH8z
hMpJlCMm7FZdS9ZTl/dYtNJlYIKew0YmQ5B+PjqSTY9S42Q04HsyoC2Tb96v3VyM
D5oEKF3JVrsxKj2rOisvQeqBeWJaPVzlvp/1VLokQOVLtwoaCTtSleQQQavjvNT0
IJL/gqZPHHf6bdAh3NhvqoeVS48N3XC8d5LQMMoZUTEMEaGbXROu+6dZJ0MUiZSf
FT4wuyP4+J5MpQuJpXwr2xy9hbV+VUxf26Ckdrk8qk4=
`protect end_protected