`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 35344 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
Ju3IpcJpVj/VshHyynUPTDdvL0SF9CTSCyUiktMH3efn68qLyRYhNbpK+WXFC+Fs
bsO+GtFEqyOLmceDxuMlVixrLKssIQi/kgBs+eTVY4w+kQsc0tz7mxbnVvsBnNJ2
c+31TkxJQxnyfsKvu7DdCgd8ykvYWXDxaPJCEJrh4f5WMgZEi08LXnOP2GPxj1tW
g4irNIXmVRU+9l5NhklcxvYpTHOdglcB5pgaUt4RabviI4ayvkJRwKt/mgsWk/u8
91E70STkBpMqOrYfefip8qPORJEvNYdQrpHWzJ+7Y+7737n4urV+TpKYVgIE+0Va
iS9fMzxo5rR9fTuksPmaNq5uXkjHv1agJ3JIt6+Yl2RSHVo6zFGltaFrrx+lkE3n
WgDjAkghROA+2YMDFqDKOVE0WKclXMTFO5yIEXwEEazWxcSyCsCfFKi1jN06r3GJ
a1DR/ulDHizTk9clHN21N6Hp4cEoHRTwraVkFsbJE1GETWtwze1xTj8Jwb0lUTsx
SmSnj0ZX6bs5cFDKm4WQeucnS+vJeq4PhewlEP2KQa613C9SU+YkDs+0Nbh0pu1H
DpOFoL77kthDztpBP5px9x/Z3j8iHqeOes61UdJQeunuErR65hGGPU2QHkFR482O
/c8cUuJdATpkfo5GKrzFbxMOfeJwRe5bOl4xiSd4ODwd+eB6HVc9T0PnE4wPPG/N
PIE3Mdbbws8M0ogttgda9iYLnhxnJ4yPmF0co43jdj9U0oq14m8N3nf0oGHD6kpr
HvjPyPA2WjRoPcBgt5/36xbdeh1KD6LB6wiwT0Z1OXVdcPlSt7QY4N5YtIXAmWGy
dZ0Nb1QHmk65p6L8ckpa0SpXfjj2igs54+VzFHIRfFuJGLmhFFl2lTl14VEsX94p
Hmvu6nNEJ4gRo7lIiJknPIkzqTxIOxkqpGxG9N7MbEjHh+2uiCAufAOJgKzN/HLt
G6Bmw/IwZooFTC0KxZMG/Blgyy46djmhBjTz6l3NrbdSoOlDK0d4mgM8DqGHRE+3
j9TRxOYAPup9YDlT1cvaPi4KsGdPNwBzA9cZ3dYQLhUT6aSIlFVA+ueR3lW29OrO
DR7Z25fSk3T/CpLL5QYvYu5sNDOvD6clUR/sqpXvlecvg5tHUQJv6kiTMejOsxxl
Lhd7kFEqsqVhcGdZVQFSfqT9mUvkxvQzCb/zzdvgboRW3OUgsCQy7N2N7IqreqzH
CKvoVZ2B15/H4DcaYFBQdY+2L5Pq737fNr1ItCbtkmRqfFJFVdpmD2DaZF+bRrjf
PEjLaSupstCJx7ANnkodpkFzMwMxJXwJi1NVohhyYzJtANXVhORDuGuu7e0ArhUA
GIUavnj6p9xS8AIDS9dSUCuu+0daEd0hU8fn0ldqMIBFrIoTddwNfvBzdkU3SAHL
NvYBs2FOIW4QkSfpeNROAvXbbCG7k1PTvoR6MVrq7sXvz2uxTGoG0r/X2mODZp7j
OHcrNNJiq4dynkHPauY3wlUMTHALlsMNE1xO6bDn3SQkON+O6+/RxqTG0SZgTtxi
4xGbfYUSmeBELnbnLYq3cLgOQjCToB5BQZBMuBPNbjeeKUHo7GBYZp8DdVSJG8pr
CfZMzBGIQ9+G4eaZv5Jy1if+VcgoCO3N6dO4NfmTk0Fh/XEZyUH3G/MWqxKc8zJ5
2pdHNwXc8njkWzJ+i0ppcUSXS/40UIBJwnf4aEwSw2CFzfFvkmjBpM5jSy4h55e6
T3t0dH32QH7XjPu9riYoiFBAKFYQJTGOmu145QQshSsGAxjyGyiCIKA33BOpULc+
uRxOrTuvMjdFnXxefXJIJOSTlzF4RXyKGyx/6tFt+KGeOHp99iXpd2cspVQi5/O8
NV97sZt/xUvduucIHMzbNuEGbmEfCtkQbxEE5QJiR0Zm0WBj9HbTG4/0zTVFbkb4
teDfjmkpeMRj8DnnLduRtfy8JJDtAD5HWAYphqObJ5E4CThxduyq3orwuI/I6cV1
VX8WCLT50gTcbpGuxZCYu+xAjED0L1fdCfziQmRntgwfFjUvkwvQqIyNtnQ0Argp
IJM++isbfZqaIAEXLsx7t6RD9U9CwfCACH5npUKb8l+66zVvozQoIT1F+oJw6+C2
1TFEq0+Yt9aSt343c1k3ip9gWW4Slw0ECMtuMA5hzfRbhj90OMeRDP8AtX8Rypug
edrpOujjgEFu6aiAoyr0hC2J9gF8beUuVojOjiJcZHJNd07MSfpV+/kHGguyRUCe
37GSKYy+TZmqQUmKBxr9MepXEdYRNhXml4HEVdko4b4Zbgns9k7Ge6+FtzJ5Pmvg
YzmSdfSWKYzBQPEdVr1JnfnEMGHzKsa9meETE3OxjjabeTSNBjo77of13yh65W5f
0ftsRVgWLeFW7cBNMk57lygo1iHJ84hflrtaOBm3wpC3q6m/ZhbJTeQqHP0w1yBp
CLMEcGsGOI3CgW4TOBT+dNdZwoKCukAiTYpKA1e3c1bh6N5KvBKLTj0ykl4gGiy0
90cUQu1dzVNp96Auk3ANfqw0VjQTHw0/6nmSrja+wElC1uBpIfEKO/anwP2yAGAE
EVqYjEoFVXz+3C8YQYu2M0LEOgr4JkmC0yrPWC+iyXz9kVsG7uJG52gUv0pGrKo1
HlZn1bWAw23HttQyJM5Fp8NplNdxZHLCtX7SlvKDNDBxr5vyzbjkYtxIbv8WYPFR
p9erofsXSmm9BvNOiEp1ik7c34zAVgn3s3HmtVDcZfc/ZXmMmljvevawVUySW6Bn
noeTzj5vT2GANncjc0GBY87LrPS2X9PAtAcPSC546uja3PNbeHey6MTfCCM+BKR0
uVQxoRLlCdFG8PechoYLf4kVJ+1zu7PVB9+Fjv4yFrBOH5fg/u+Q1N3txnC91Pnx
6dsXn2GfmeYAFIb1Do+O0aKiENLNyfdakdra5Km1IIrhq3vC4jxRy40bgVaSUfJn
i/bzpOXh5lk8cANBHKTu58ndz69YuKnI/AgyL/Qf0CbJxJWTzSZvqwQdNbkOu62O
czyKZsCA4zU7cqAspx0P2EHFK0FexzmPMkEmryzBAmHGL5HU9GQKU8R7axPXacZR
56NBlhb4S6m3v5zLRjL/jXPgi+YrGU4se4ozMznn9k5jY3bwTlRuL7LTKOPq+jOf
NuYTNph9glCwNfunMREZsGHmJpCfHbtL4ae3Kwan37ZZEPm0NobmMv4KJd/Z9aUk
7pNkEnEtKsNb25uuQIcIQeNzmR/yD7zM91Kbnk/gArVMDmdUtO5lWxW8mvqQCHE8
VtRrnozw8QVzrlmpzo+TgUpNOlLVmpfRS8nTEezt/M8t2Fcm33xgF17zkkCYzjih
q62TRHfctX9LQWUFtDxBUX0ABPyk64731ZR8gW7y9/BpScRbZ+syUIH8LhZ59L8a
smRF14Ya0WAy1imncdNYrKOKafroevdAlXafg9jnIOxYeWq6lF+3mRA3+pgruLr6
523Fr/UAmrYXBT932gFuZJDz2ZXaOP11wJQvs+PDEtYNF0Ps1OfpkKhjs8jy6pbA
ml6ZaLUC+QDCCl9x7MPSMByBNaQ4AsBZ4XkHzRZolgtCDYvs5Wf7oqHRkFXDioY6
bJUC11uvHvNQ51s2mx8yJFbEoJ8G4nVogrtdAZIQjcpn5dFHsHJv+6rCd+4xBy2E
we41UFoouumi9+I5MoOzQdfla+Q5mmvRJGQOc5OHL9Ce2j9XCQDwDmTin+6KUSQB
wvwBXJL2hGWWdn6MzcVrUqhEqNpsNhKrplEctRNA908zULhSkZcmqZS4TDN2Ogp3
V3Z6NRFCemAF44qDxbGFUaJMAaKxo9UDFq5A2S5EIhZWxdX1bhzou3QUaJrArxl8
musUFvvH/X1qSIP35W90uJ9VmAI3mkotcrCig8PhOTGxKieazf08QrCY52LmQtQf
xAqf7gZ6+38EFd9sovhl/wQj+xlVcTELVAld0DUChfWwtOpLHfMgh7BzEb0spPjQ
x+XD4jvmeuyNxwE71saPdm7Kli/s/ubLMX6L42IdHUw3ovf1FKbfQgscW77KT5DB
Aptdjwuad0IY66qynjBVz0zFabttT1AP3Z190wrw7uu02yQSWW20kjF+YkhA22P0
b1LQEkyLi1zit5OXW2H+Uvc+ghLVUJVWgp80anQcFoqAdPt4YMVoAIYOQToJ2yvw
1sLOsO/Ags6+9t3XJ2p7xX9MuKAfgYDBCOUWJTx8pex8YpBCk8JhUFFXQsmh7oHL
GHAIPpYDO5Xvi0Ya4L442Oi+kpV0a8vyOYt8ZtmxHx4fqvKUEzfzTpYzIHXyJuYk
Q+FEkiru6sObxOUZdPyudUu2E3ra5WoQcXZdNXbtQDGIMqxryh7mGd95zg9ddWol
EdZVUpzI7snra3CT0mt9Z0qDX0fISDjIICiiNC+JFA9JLAiZ6ZPcde3p5TI64g2j
L2FF6h2I99X7IMwx3/cI+OlgU/4l6TmnKQO0oF8v0C61gils+Fk3uSbTNwDWEIu7
sgHnJWQM/+Yx52y6ZzA0rvg9jXshHqR1w3Vk9X+9xBWXgWDLn6MPktlPtAA69F8T
CNqzk+kWzx1onwX/mvwfbRcjDWqZUpT6iFZI4w6WkKs8DvzwYmN8CzbDcnMmijpP
0YgjX9awNbhXuirfBoAEOOth/twTzZCBHZVMQW8F2z9AMXmZBdvudVp0TJw3wk2Z
NyYnDgmTzWTMMGx95r/QzkvZptpQeacrTXPqNSqPwJxozOTbEi2aZ9ZWJq8u97H9
C6zo7hGm2syOZYj9SpeagYK8LZ6xG6zgA6/qJ4jFUlu1usvMrvIjopsh5U/mWEVz
Q5/oiMwfD6dPDt0PX9uu3P2JxKQIwxj9v1FAk2szUN+4J0B8Qel/rQ5UbrsrLAil
CvlokgokWza1gwARwMKfsgSAAFnRUPfyVZ0ySdQ6A1X+FWmkNhFPOFqfXJDtDrbY
hctE4PKWlLcYTYLaA3GOs0zBUCZ3BstvHxeJMT2tfhQZ09Y0BpyqUH0+Tj0bP17A
VSOUOa6qOgmANqrYyWTIRdffLzEPxiJwYW+viODrUfa7GVEHoddURRpN8V7VQ7wM
YIlBqxPc1BrBZV/Df7LOF3XQltXhgavaKNErHk9gBxN8tCViAp83Lv80+/5Ei1dO
zWNQVkSTDd+lCmL2qySbcsXHIazUPAau+lHlUDKA4uvmZKpWdOqM5X4na64YkG79
U4VYp/FnzI0fKHeGnQqglxd280FQ5nUk6EcawEoUjDrfWZbcYSLV9Lad43eF/eS1
s5SC53UOHXotmYddLE/W6zmeBQYGmZ05FBJLPRwfvAN+ebqLpWy8Fe7lnJ2gIdJ6
j6W3ezH5fZzCrf+QyULas5HjnNd4WUbTV2XOk22qeu1oBbVJQzZRoXmVA5A6NRBm
aguamhAyjs/40ECSc75LnO7oqd5xkbQGv2MEJm/mPEilrkD+kiV7SLdc45oljd7I
fn9RRXe9uj9LLRwAF9ZHkPNbepSzHcvGlD8sKCgGRDao05lEHbxbiKQDVJ8D9IHx
K0kYklqDuHyKwwJI3VJLeovXs7zmZp677BmhVCbe7jYo/5KSgnFvGFo1unztHtD+
QaEgS7YxG1VgJTeiup7kheHRz3V4t9X7nTrNi2yQd/gFmkLcQKWSAtsWzwLX5CWF
NpDOjd6QTy5uEL3r9pMijkHtnrJLbTgMWj+7m/au5+9DYrjhmDRirUqpjNciHFkJ
ZApLjmPzbYcuBlO5nOVN03BwkAVB+R0qhx87hJj3PFBwsfWYVgBHsT3nvwIF5hLe
RoRk52SqUjTMoCb7aPoJZZZVLKc53hV3ZaS1xTOTkb1RguZIEThilRw140x0j113
ICN5VlvB89c6RNxLA3vT4e5LF1zCMomWVitJp4S3hBo/socNDRXWowK40fHOU09h
xKYgc1rjuRzridyjuRQwta//bC5H036rEL+DiRlsS6eBBXriZ59T1U2qK5PCWQRw
gZfhV+jA35xL/yMbrQ3XCbS+qsnxBUrdmM5pldLy+rbaq4/cv4T+r56P1wOL8SCk
eJMKbtn2ZAoMgNFG8fp936FxtmGxxjoiQ75UYKwX93TDxFviDk0vWpzD9CYr+kFm
OFADQc+0JOjUra2Fevz/jrhnrcUC6GiewPuL1gnsRFdNPgTDlcDKzwB66e4gTggh
7nzliapHIy1Efr8Iimc9v9tgf8iEv3y/lbs+91PFGWg2tU89DfR5CckoQSCawL5Y
lB8v7sfPYErgChvZEzb3eCik6eQNjpn1JNo3kHduZFfrh9Vb1wevB1ueaUJ1YhcY
+a2iCE4y1aYPd1OdJazXaw/2t6ybXgIxV3WK+pL5Qk/VkgA5c8xKlVk/mVhhhv9S
UoGmyYwbqoJk2Werg33mJUlz0pCPgKAnMt8ED0NQruu1Y19iWVbGhPJurnyfuXXa
7jZvmQSzU39V5N0x2sciqcrugQYdVl5/t2Jt+bGkWQbwb3pAwCDD+zYIULbj7TiJ
5AbXSE6gfvhc8Iy/zbXh5gh4BC8VHIDYhM1qzn0cvC7nLM4XYq8XlNtN1srWUj8M
GUHRqZvgMFsA0qg6vDFdherc7euOodE9Z6clK9/GHSR96gyGi82KBd6ZYDtiWIIh
MlSjA+PlYFUW7u0AywqFxcVkX6p909Tvm5Yi/U1LSW45/APCuQpSPC69NPgqFU3T
ct6UaBIML51r9ZvYNYK5ROSghZKxq0Z/qYj0s2Vipepn4ky8vLOSconRJ1R9pKWg
D8Zp59ATVfRTTXh43/9LPEAohnHDwOTBd5OE0dmzFX1ZK6MLB/NSHrDHrf0w/YHH
x389sKQdYAxN09eEGXDTrFOuuquVQrnUf05vTKre9noxIct8MRgpOHb91lGjICR9
9wEDe5WyNIj0xdtGX3UCxXx3YPabPtcrF7mXL1IntUtMu+tqjWIbpaJk/2PX/rtZ
mRCzcOt0gKkdruqL+PQqoPbWNBbwVH4OcMXoxTv+W4kP1ZhWxnpbMvIE3aAZXMi4
Y1a8/u79dmcWRlRa5vArTc+B4saaEDxFmNtFi4zc2k8a0VvouRpbO2ZMQk3zRVRw
VPfRrJnliJhaHP6lWNZXTerCkPlVVlurMvfvhd6XoAuWgYsp5NyGoZ4HVnrbUZEp
zRJ9WbNEmV586lqdxE2b9UVoUVKLwpIKF9u2KRrdKBvCn/NtpfkT+8U+y9cfPI2C
Gd0ws25Zkdhm30xw3uKD0vFabL4k2+UZ+xokutGETafmBYg0so4fC54WXty682C1
jHELn/jKTdtv+LNOwGDdBhNWZHQJCBp8vdUQ1NcCZP/Y3iWpPuxwi+sVhh2fy76w
M/i10hf34OcKzfmsHScVEMLM3N63xLKr2whqcoEYtpBfpCpEuNkvEyy1IeYoCayV
1SLMHFwOCdVgImfXlySoC6L1+x6fbDPIqSecFkcr3Tf23UGtZfv5l0baPVEqfOBd
7w3ZRX+SiwLPx/KPSlK4zSyTJWyo/JfwiicpfDp4vy0i3CW/M1Rh6YawtQoHkzlB
NiTVGeGQynGxRbQnxY9nmGX31uImqjLKc5Hj3SH9zXrobeqGfQ5/hao8izSf13Ef
TS7L2dxN3Shkj7RjUrNtiQMM6PDvWcpBLynZ0VkwMmo90qKmHpzm0nyzhwqg6EHH
T/MyZss+FJ9gjlaPDOC1PGxxt1xEpI1jWmZn8/wa0m0taSdsFj95hQLO1+Vrzy+h
9T9tgtkIePmJlLjedqxH7wvTs1Dh39Ij4187lzEceAGhs3GqBdmyRH3eCGTKBpPz
pULNFh3E6QGBhUqFX9UgjkCusa/PwfWlqL9mGH6tFdKXJhWNPhr1k8BIWaHknbTY
/gwt/4Bv0nZGgbigLR3awAYCxWFHZtiiU1CXVrGVTT/q90uYDBTS4p9hglS8ChVe
1cLJbTjYjq0s0tOleGtZ9xtl19i+Jz5XNLj2Fix+rHnb3nDK0zdKzD8J1vI34rWg
94LU3ctzUfjm+h6Zd5zzfEkFtjAvnW/CTqPLdpwroMXD2tRdeD/Y1Sb3qaPE1HN/
b29fsHjeWSVbYz83jmnl6fkiazeycLiYcUdtNFJ5lCekfXLRb8Zoan+E7dyKoEtA
XZPfFqGeXxHQ+Aq72uxVsmvaHZ5tcuu21hkgYZ7Aj7uPlCL/4222l8h0BL5yfIyB
I39oBEb2eWGsTojot8SFW8Bl8K96Oy5qDo/YuxxwLupW5QzENu1rsU429uMj9viZ
M5jiuBhAqaxwgxYhcwEjsms1CjNwfhKK6lHDZKwAsJoC6J5adr+JMOMVNSbQotIs
U4FQqXdPZr565P3cwSd8ZSyeNUzBIkGfkHeHruT6tBx/fRFdFkZo3Toxntip6Hxq
QZWC8HwMy/gNbqKHxUKrLkp2Mn7eA08OrgpXh06fHqtI/WMLwrbE4o6KgoXOtyDE
7SORoA2kSDURHauhd0XA4X3aDXThXh7gdUXkPJSKAxWbjqXpzXh8MvZd4NoCDZHI
wRHMWwgDe3BQVjksgzjo5fxwxSvGRcgYskEAWHqP/S8ATo09eyzJHW1y8drgeaB1
IsN7u7/Ra6REGc1QFz2+2L66WlfAKoznSfVUZAZbEnleeLb0bRhVbHsq2e2WuOUt
h9RKhrqESnhNJhgvTcH9r8gRLvAz7a/Mp/PS2YB8GEkK/06he/nl2RsVpDwo6Ysv
tUKR1BIsi/5tO02jwzsUAvdOt0XQk0mEFX/EdYWWOwP7Tgsz7WMszu1PuSqktuHw
3vHopT42WAHac6BX+OJh8Urjg5RsQyBeN5UYcVtoF4DRW9UQXF/guuyoT76a9yCN
2EeBbtId9fEfHI3qQE92t8ElPl5viHUUk+LUfFfy+6uORcWEgajEY3hn2MQSgeI2
uCcVaXloe54z9k8+MlRM6Ekt1su3ur3TpdFnE7kex/Zf4ijMsW5yiRiFgcbSCETj
k6iPTKBDlEuwuzDAF4CqjQog/+9dtu2NOFpJ/Ky4SV/5W8pVJ5Rj4nzlu9CHmUTx
kN0U/NYsLIk3f6/V6p/eN5ywm2AS8lYy4awBvED5VqYp1L602mQKf8L0DJBhKFVl
GMs8JLiOyGRcXj4zd3V1C/hk72hMzGSv+6tsL1pNyBfvPCJzrJuxC2Zss1xiMcFd
GV9La2Pwlbxamvk2tio5nu+HtFj1nfwc2JhfPh5QmClBArmx+D5s+eIolI3WgUTC
Cpj8XbJZHmtmQBr/je2OlPQD40jgpSwGSNBw892yfb8YuMgZEkaVnQUy+zNhuxJa
+NK5O2WPljaLh65mp7JVMsVjQAXX766Z/HTeRKqxk/nLSqxihyI0v/425EXRaabc
SVdUav8FqoP0YaUEAqIs80M83P61XRkm4ODWOTKLxOFb8hyaQtS30OLo52Xwc/zm
JXbgIfw/jrFc2kHDCDUinamezdubC6rTNKhTH5dWWq+KGi7x9vqzNffNLvdFzh9l
rtGhPbSDBgK8LiSIQdzYz47H4p6CkYltL+KJPQ8cOf9G4OUwVXLMgxwhztazMPXZ
g8obZI3tAdLIPvXz2MznCAKDSZzDtrVJ7/Ndd327jDJgc3CcOwRL3hhmoYZbex2u
PHrWI4bBaynj7ou0VxqKXesDx5DI+GiJHNqmCHaap2bHtSEpdnsrvzgfLoK6wk94
KhypsxlywRipmUr8zJOAG2Ooe6JB1NNhCg/DjkIUfCW9NJd4l8Ubl42BknNggBy6
Qq7cCbswRDPzo/gMaifcczqXF+MPi8p5u+xguWB7/t1NvIw9IJVRMGb+xMr1jhb4
zEjvfXGu/o0kf2hL4hG6E5D+bu4XWgP4iWu550jubl6rHm8QSBfIx2bIHsa0tUJ3
DSoCq6r8PUotoFAAMK93VUPbiYHK6hdphc0004/JxPtUYSiMZqCf1gQo6Nxo+dwg
XvoG2wq5p6I+KEZtMNGQ+Kz0DvGTphKVBhhb7SlJ4Ddbg6FCbB6ISEchCbr10r5T
K6xxC+1un+ZXnD1sx+I2/jWRO0g/H/d/tSH3n26yRJuBY9e45yhFF8KDvkv5grGN
K10ni3ISCIKY4SwkFEKpvlsuTZH0HMW7kmUtE2Wi0v+d+7Uj/ohPewsiMiYGeFmN
32YVlpTafWfi/+1mrPG5IUzuda14yFpFen5/oq0Eafwhx8ZTa48dCtpW5vB+x1tu
CLGliiciJ2El/uaNYM9KZY92yBHY7FS9Lnqq+3Jhf40Rb2RFgczLbdNNi7rtTjDK
QLnjK+YtIuN1t8qEBxYAOqv3FBau/uyiqdRsXCvy+e4lOcr67cQi/hzIq7W/ff9Z
9gTIRzijHBIE/OT9DRPVCx/fTSmNIvmrNYTAWsHiFWFolOuisYF5rzQ9zKbxwyz8
cqgEAH/lWCflG0NuXxob8c59fH6SD0dlDqKijK3bUzyX/eTbvJXmdu/dituQ+vsR
nulJLWQE6L+iVNzsO+rP0ScE3jpubOBCgYJ9V0Om/8wo8YFqa8DiesouLzb8SuIh
5RWMxVrUrkYeEtUM+pyju+6xLFHI9vOZzORXIdcVdBNZYZcSFqSMaQl6OGXUWxjL
7vwQOA6T2deqKzRvuredEHnJ1wvCxAqeg+pR9eY0B1s6oMvOxdxTdhkK92kzk+0J
1bMoatMwmDHmnyXJ2su8sI7dUAFhsCGeTT3YNwn1mduYU+nD0JKqX2bTQMk/VqWm
spc2xt30wEIYlvV3b74Rz1AOmzVgBJVvHIubr879nuv13T4Zde1Hg/lltqVt7zgK
VvhMxNmDHOltpg558FoUEhvzDCJGoxlwngFtrCg5kl91HYYxErs8Xd7zq/W+mtSj
xlNqgoqmonQeKOkYa5OJRN7AJF7tWd/8HN7cUth+3DVFMmHob4g1ibIuiUfymzUR
POHTKtSs44xUkQCEUBRlBiGzGEtNx5gs3trkxwE/+BV1FDdPpg1BvWHLo5tKbVDK
yhA9GulLc51UcEUiGAzQIYkXnzfseAI+zCzTnXKAZuADp/NRj/qWjn0CkhK1m1Ex
ruyrHorxHSn6YAiEPXWLCG0Gd/0xk/JsOSPeTFimple9Z+t93jvNT5mCVcIkUGU3
e+vRxKTutT5Tz3uokNAyPS9tnYJJgK66Ns8cSFNoJ5Ap45hpJS4y3XIxuu+hQsLx
HfJ1hYJprz/H1HIAcchOB1W2Tlc/LsSo+VE+2eQxfqWOWnL635XOTt30J8Qs5m35
b7ytTl3BbvQaNYfZgR7vRSdGR92tdnsFyOhwnnlg2GcOiArQ6nw288m9jY47+1Lg
G5twqL/crU8Q844xv99C4oE+thxHVxJiSicxN8FteEf5pfhIQUG2khLorueZxVry
UhePpm5Ydxr+wuNKG2MrzvXRiPmc9+Q5stNZVw7nL8PYU7wqzGg7L5E4ODZZuUXZ
TekTuVB7tfDn+X+s2BqFAhowcxMlpNDtwfq7O1DGqnjsAFqlsWOnlii5H92BQTBS
BlyHp2MvTzaEBtTmYUIuT4qiB6AHrRmxjqblQlGuZ85ZgUF+0bw9umWkE90W9ctU
pjDjS3vlhIDHoiR8Vc/Yd+G+KM0aoNnooMYByLr70KKCLU64rj5b7EFrFd0PUtLh
aqvgykfrLXCIXXwRJd5/EVWanSxNbdreIetXM66Fl4Y8ddWpouHqi+YTGPMHc18v
ku5Gbg4EckuckUmAiCPjHaeWyJMBUWGOpYymAvbzZkZY0Pb5CmgIQD+FnnTK7dpU
m6lS+RGHnzXdNwe/X/mr2hOFozQdXB3505V8H25fmgVmNo8WXyAmKfKPVxSE+TIw
coBJeoqkY2Xqa815iwN8vFT5KvXXEtWGqY4q8BPEdYCSICz31OM0NoO5/WWgHvv+
AlsVyt+GBcNwBnOcK4mELZ5Y+YDm/eTEy/lzSQcE/DB5SUn/OuCNb8+6R7S/wyKm
fdPu2Lte9u9x18jxH/eU8gZrwMnEMr2iiOGVKWDgRvNnooQ0MMN9Hjd0Slc/nJ8T
+lVM1C5k92A2UBn3dGl2QU/yQKyiOhdpmVYTcd4B02QRRwZcI7cVpy/RM3THKBmM
zjitps1TKidviiIacvT+JMekJkwRZeIU82XJGRDUuuEyhPpB5AMlhBIDl5oWqDsf
1pDy9Jq9qde230o1cmOMYnVYjRrqtSCe/Re+D+2zstOh3i8fAajok8wKv3TjW/Qw
HXAf6HVr9aXeGG1lMQAbmrI/8AjFtBMQB3s4GFL8SZMvKRhMoQp9AhZq3KYkTwRM
Jgqjxvh/ubRctsHHB/6+0tX/rLMqUX82d2OBaTrnzcQcQdJZM58VQgiHihCqROtB
DLtWKJs6YCGjFsb0C0R9EoV9u0zhf7dedZP9heAgtfWOXdVhuZOGHTbObm1FLtyp
BZZPCHNPfoerrc7mC5Jue3NKx+JXaK+TnYM/MVMeqCWGLVesFgSlG4QsJg4GiJDi
qcrfrMYaE2a8EZSSRwxjWyS5m11usCNZiFYEJXR2hMVgA8M0++8MJ4wnKA4aSYt9
vtxSz5wOXkgzFvp4MnqTLK62W/4CAD9RFNfLtQrN0ekx7ScI1R5b+51inFUSFzg0
IIiOTyIqJN3X+VzUTpWVTPsljGRyLDQjlNw4/KOTmT3q0llx3PYgorjhlVqtdmxw
SRbWhbjfCY/dC6G7sn8I0Vqyc+VnucbUew5YDI7OpvuDD0sXmcytI334sABD+mMQ
WkPQZu52Cqy6egjRgn6dXltV6oMaU0e5khP5Ok1o84unq5AE4noAembufT3sKHyF
YEz/NfS2GPhkaMdUlfLBUacjOHfjvh2CA//UAenXJPw8RcWnwQWyrX6/siP743JL
BAA4XttL8VjCkLCvuUgQ1TM3daLQ1IK4qEnJSRoJYOBc6PUE3PyyNS4VNW27Dstp
xdz1jbfs2Aw/eJqVXLhYBfhazBc1KDjvTZbD6WuRWz/E/x/nW90Uk8+igfp2Vn+b
SdAHRY2jAWtySMnZh0fjvGQSy9+Ovj73hpdAe8Z3clxBookPwY3ACO6c2+PDskSh
05I84hxZbtVJa+VnOvyy8dAJ8KX8Ke18wRJgmFz4mSTQ2AKP5ve6A5W2/RlWIuY3
rIWaw6AM+OPVA8HKuhQb5L1f/51urfnRA3DMK87huUiWvzlyh7LPpNFJ3By9Tosy
PK1+DRFP+MtzAlad8GX8/ZDwV4luDxZj74xkGF1FbKaPxiLgMEo/7gc3ULSG4eBh
7vLWvu6HtNnyefDWZ+tHmaYgHXjkP5GcFp7FdYD2EJiwNOUeq2uhw9GjtuTCTmyz
rHReJB+bAZKqmG1zBXBtOmhCnJ+fXCoXQuxVq7vlopZAY98cKtWdfmOa0bjtStC6
NWhItjuu6anxCn/LE1tGgXOfJZYVjvIkFZbN7AvG9kuj5km3iq0lOXLKl7aDZYKk
sMGAmKrU7QRTGRn9h87SnrzMziNppr3PXIuotniP1/Teo1J1KDR/aZxRoc38PqR/
3AZkQh/kj0Y2Xe0i3VzD8DUUoS7H6ArlMLChRsC51xmSE1JUMMrMuvuLfUihDooE
gzAfNaqKGPN9+E4V8BKbHkLB6ONlG084Zp94LJvtrClJTv9BnubpPwwoYLayFXVq
FQyrQlTYS3YfvrQ3P/TRFyXk34rpbBjQHlWamGY6bqS3hQgffC/h4TC2Hy1xC+89
eIjWj+GXIjD4blZhm/Yg+cKrJ0UlqVUZslPhjtCVLBbt5Bowz/vgo01Fx8/MYGQw
erHIUN77Nl9Ly171Kgcr1Q1JpJxAXJ/bC0PEC0aE1SB4cIvaJp2H31GOWr4wabNm
z29TXE9vmO2y+9RjzaTDUbevFUnSZESkd4bI5Vv32vMlJ5/CtmzvJ2EDekTHYva1
XAMqjL3W8VtZHO9a7oHnsOODnySXkk0j4Q3aqtlm3hAs/bSTR/fQmFQ6PHNutMPI
3cZ7h1vzyNKdDgFN2HJ0OWsnKRurWkYRqACMsnZOBFXvXr/e3LEk4wOvuc7jMsoY
ptU8MGSKOmKTt7qOGGIDq8CKihxVgtojNZ6+KngyLRfMVipVwLc1dlYDZRe6Jyy5
v/ffHWk9aW3ZQInwIKWyowUXWi7pgSHE2cgdFaK9otBv/HhcUYTbFpoSA0PGvwuS
HNx7YqxP8++bOqaYMb+eEvHbW/fiHIeZhrxf9DiYs6ixXu5H2xOtU/nhuVRk5BgS
uKK4rI39jsjM//3mKkG0GFll7vuaHE+xhLqukrstj9xui8OEmtruyPH/vXqvrn+a
2U6hJFkCm9Z4GZa6kzsKmdhoB39dFSh91vflmqawWcdWhkzOfOYVkFNXVOpzrnBs
hNVwbB2xFmAP7pnY76sqesE0NAyvIi0x1XORUAct7dg6OwB2dI9z3dt2MprOgETf
skfWFD6zvVpVhsAQPoXdUhMv8r2vxDjzV5HAhrZ8MWnz1iMdqrmMx3J6XSkr2Fm7
sECA/to7QCqXDhX8HvhuRueV6yuq5PRJYcyqNXDHCtZLxebFnDT/8YAFp66dpmXG
MtJJJmPpBuSI6jfQjJeEkiTehFZpYZeNyZBcqL8VySv3Ujw15upqWq5cYnMT7pE7
CsNMaqvFJNtVWrlUNZ5QcQyCAUFFrsPqYVCLtnLJY21h1stdMVqc4UzRpFkV75el
jZgdpr/+chKVNAhVao+P5ajaudKA7JZk2aHCug4nNSEBq7xkol8l6/qNiEGcSP6x
K6kl8HZyhNEZVfxncUvLotuTa4FLTeLvYBXitnirRnDPNqYyECZNqWhfEwNaNsrw
TjG+q359uGKNXiQQDizOGp72cxZ84Pmi8s05id61jCrS5V9TBu6ybxADK+kftlYM
20DRvm5o6fW2A9lxQlOb7GM1xsqDwUEBMvMe1BjQcwjNWbbDOdtBa8oCZNAQ0l3Q
M2JkYU8Ead88g6oZ0O/neV17iPjaDDN/OaZMl2g8IioalwQ3YjLauzQUQGzFzV0B
KBx1R+PZk9cQuEolbQLiQnDIbkWUa/1+6Iy4RKskAE/B9Q4r2O27FwNwX45HOP8+
uie/JsHzU/FY7e0fHS8+yUmsaVq9Zhc4AdLq+qxQ08h/kYugXRCwaJS4PD0TC/CC
b+L/ZF7aaYwgZSQ914HTBk0Hm0Cyb5zJT5+AoZGhUGTvk9QgSPQZSmSyMYxzuX9R
Afx/KguITmEgIk/H3y6wlH4W6buXtVhhogEV1ycLWQO/PPt8/1bW66IL6ipvRykE
8v34iRauTk3g43aIhQ6yf14eNqBeZS+Frc6cqW9kPsJvwKvo3EdyLr/Ee4WIqSba
qN2FAFCODLRkzBzOolk53bGkCn8CWKLnaj9LpMa1ju79nXFeS10bMm0fwocTbMk+
k6t1CCBIwrfCnioqGKfpOBDZ9hCCS+XL07LmM0PzDhUwz+ti9099iQuCJxIRcYPu
Z1oMuPP9CPtvEG1+BODKcTVJIP273iZ7CxxEHgfNMj8N/x+kDcbtnh/G8JJyWf/Q
dZ0g3Rc+ktCj/pvus7CINWP1/mfEoab2+NoAwcn34HCgcNH6KZNn/2eMHBN2x+zt
pMgdy5YQUmoHl7A4LeSEI24rxvBTyXqqDUqDcl1/nnWKhdVUNDdqKTLKaw3uKAZI
B5RosGLJGB/YsghhM71Geu+XTQK2mPab556S39RaDAqfFeMwvigri6R1RiCinbMU
X35qLuTIo9jCefANWqnQ8ptQiKzrHfJwGRDZIixKt3QPWuKyuanbbI6DScn9M7pr
lgNE7aOYZudEDOceqUarmyr0ECAauQ7yHhZ+pT7LLtO+RzQxB8z5/bOylK90cchv
Wmh1vFSmPe6895mnsKcLpmPGzwHM730iRWtAqZAI473ycYyRnjQ0iCnkKzmELZYj
EtcgZeX1+wyP0SplENiK0yVGPzDxL+ROsOrGse0XZOEgpsRIYG9hQun0OY+tMCrP
QFPv63O6Q71vgjfrf9yEwACxdhkxWT6EyC2YR/GYMCBy8asNJMzJpQ+0DpHSURNa
vY3iNG3SEp9WpBeZlPRZpywlLCWvjbS3i36OfMAyTSt0x3uPH1hjSmsu8oXID1X2
aznsC820J5nzXtpxIg0BcjcZwHGG8Yp3pJjQ+0QfqYqfhZ47TFMvvLMxd4y+HRA/
76qi4l6JsUTPE5kcpS/ASvTfT2IdO+yaTs9UjMkg5psncwu0WVn5F+9m3NsKiZT5
35CCjMtVVjhucWM36Lj0+ChkN3SKjd5k/5lgjGYmB2RNEZoRfp+sdjFgbf217GWO
HKkiZhmhRHgHuG3eIOwddoJ/vYsVS0bWa+54op1Ys7+h03p36KLAzu/WyUhv0lJO
sTFz0kAJ9FxyraiKa0ElptwNO03rfnOnTI8r14osATn3xSzrvULhOcm/Pqia/nt0
QXMy81PYbdTSZW6d0+3VVTh1wr3evm4xqE4HM7RJuinYkYwO9BzwAVvybSEkBImn
R1uhnE4yOADo1eK+lgs5oGBZzoC80lGzTgEScNgX0OOahfEE/cHYFwkhz6cJTI22
Kt+3TJi2un6JnHQB5+l66BqfDz2y7drgFG8cT2AKELnoJiCOHhhKnYWqEu9zPVsK
AZGSQQudua+LoUh7zydlP4FtYwc9JiElRTyfBmdZ37t341vQfhsev7bHmBF127RL
CFHnqFaZVjK6PBKSxW3vkAkqgwH9ILodAoGWBbEnw2EgxU1PpH4Mzp1olIwkNs/1
pCouVwrj8V9WkHuWOACWCOSjZ/v+fFU+AjZLUvojTu52FVoIrHjK+t/rXR+VLsts
pvSx7HLBhdu/5ddssPbKL1k9U3LMqyOI4KbrfORNqNyeSuuHrylfY2L3sf2fYzii
2Qz0KuP/E4y0ekrEnYUP0XSqheLknUqFe3MHw0x22jKXYYa1dC1NzHRWprYI04f/
znhmYYfOwGw/PqhoLQ5MjHyYfsQZTvbD2EOZClLhUWCQUh4++TEALp3qUUqt1dN+
ogRX2WYtofz5Q82BtYLr7uOJiE+sbRqgE8OWW1IfDPNsZp4qBYDykuDr+umW+yrd
P6jfpACgXS5mVbO+tqMT63UwEMUUBQ/+Qfx+RmjJWfyTLBhl6MxBlKc4jCsOqSxt
vX7e+GRBUql5ozQo+MD2Drnx5CmpSzkJCWEOMXie+OAbOppAfdrtHYsaZun9oRau
jVMz5dnGQRiMfN5hDZjp4Zjhkb/cxCGjE/rGalU9STlz7Ywn0N76JPmaPtC3ZnR1
5fTu1uT4rPXZnwLeHK/Af7qaN5Rb+p1oTK60RS1SxN/NrZbqTErLyQduPe9vTDB0
1HGdmcMDlxQdUN9jYGnr7TRDBdHb63letiVIGaINxmxfZnu9GoOBROZ7918l1KPx
ej7ic8xrp07t0qTLd7vReOh4k2Y594KAqdylzib71X4VfeRAacpDifHCr8jPWq5+
8XWdLZuCTrA0HuOzC8cJWZAm9r3ueotkpu+kv37zCecyLwPesvYRXvUXFtiq9ok5
qEYU40hxNydcaCaDETtCwIv5OBt1nZLhqIdQkUfnjvZPy+9XqQTOiioI0ooWeIgl
wlor/vNOdPWfrFKMlPs8pRBB5uoG/CBxOIStIjNJf8zY2C4wlen+qUGhOQF65Hpw
HwsPI5gGG59OTnqFbeb2+3aFCM3UpQr6i8cb8sCivhTN8kqFGvxKTfWRwAeI4Up4
eaKP+fgQ+sHaJgae00o2TMNun/eBVeZNfAiv04xGKPISBQ05kOEoDhYtVDvKo4b0
O4VsGsbnx/lo8T3ShegeNWOqnTQ2ELnb5cjyB6ATwWFPyv89ANyGpjEdW93opiLV
OpCrC7T/W6DWx98KdZEtTlePLaOn7q90kiVLpuicEUdzMKAV8/5LKbVYotR4HE+t
sqvaipIUJPW0ziRzlhjaGfDWz2AKEUtoSm6SQ5zAJl7mfpo5ic4GNu9VIL6s2XVb
7bPT32rGs0G6Cj4TqFX8+w7TD9yp2ObJDuCUgQMy6XvyatX2z5FCSbMhMKYUMdtT
o78IbWSP8ej7W+P+FnTuV7G57qQqJP981JL9Spk470wcXR3ETy1YY+jhsEziiRr2
a83acxp0tZIIv/XwIjZxwqObgruNuWMZ4YNeKJEVOg5CQkDKq45uPMpD6otvC37y
5CkORUhV288HLcLjiaZ4aX1E4dGlXHDYxYzW8Bt1yORHTcOp31QiiWYiehBBJpAd
dZQQvKevPcrAJTV4gcgfSZYUdGiWYS1Uw8YaVAriWj9jv4+oo3BFLB/9acWozv2R
D+mP143+XHkMWXuayUKnnIi6qX5xJS0UPGsg/5GCvujEMuXAiQ1SSTLaK3uDH/t+
bj+FXbAcodq9+dJ8jL8oBD74NoPJOZJ8aLGhs65/5nn5qO6dl4VDiIZFA00BqL4n
69zkF+Oe+mateI2JnDErjfzNiUFPy2q9clXsmTY/bCcQrqc3NAiAWfNVTrkXeBPb
u8SsbnEpa98zEndZyDERhV9i/XP+EQX9RXelNhsI1WiF8scB9dGcclRoUSf1BA0B
ajUqMjDsInLhtWC0ATCYBjW6auUL9hD4V0wybt+n3XgP0ft7398AsIrs+71Oh90G
VYbTC6jbz0tKfVXvH8nxf9pAXi/+qNwpe07nVToCzausJzDY/1+n3m1O/nbM14u5
RWe+hiMIoxDNSykskroe6rogQW2QP0r22eNJgX2Bk12cOrffyJCLQWXvdDkmHndd
Se2+/Rg698tMlglfYtHuGwqNcrIkVXVvsAEfb3u5FZsW/4wiZlShtm84SPF+DHrT
Z5Iu87f9opy6SxXylkYx2/eIUUjKgUTubPeXJNE6MfUzqIBGRL1TclgJiCiF81Jr
1wS9vAv34MsQHhdXAQv68UMdA/80WzfSKaR4JBhto0dSx1cKH6KnQ6Xcsd7EgUo5
vouAZ/ukPsXM/e6nEXeUj5aKLe1De7yOjW3CwSSvk+TGi94uZs4rfe0nBkg3U8AP
DLenwocodipMSQMNT21W76L5i1+OruDm8qSEWOOUnGMs9fR+btyjkLMBhFk2dL6z
wd5dTtBap6OiXm2PqUB9H/t9IzWONJhB2iuQE0H8yJPcrNMkC1T+p0jHl7gHcZGx
kL13TdxqHxEiLI4ZN3Z2E1aRU7sqsaDg9830oJFLv+D078Dcrbhln8sBQ/oBID4K
iXEWK4CeQ22T7dYgCIDXecsRrNNJGVbqMNX9hNNZl+awhjBxDV3msncII0TgKoQb
6nOM0z1PxFpiUnSZ43WOVn/xer7/gIOoCgDJMjWP1S5ZzTeMHfffNvoDpX+J76IC
wYx6VefRRRXf94kGT6sB4niKeM3Mv3T+/pAtXjgp5sJyTWpVSVKdynkjCFSKxKIN
bV7hd8haTB5y20ipMyXxHq7bO9Dm1y+wLnpWoUdyGA/L72/ueC/qHDW1qnM7QZm4
By49t0NcZXfDpWEARr204L5+uFt1xzcE0j/FQFVY6POI7TZmGt7o/qKQtRGRsz2d
QSmfWhfXFMjBmgb1INFaqHTcjB8hCD9n9mL+J+nmrnaVg5uqDFFGBnoSC3rGQh2V
zaNYeGWDgnNqdJerwLOPrXgb2EC1u6+8zQwQgRQCdw/0GuWuCQI9qs0oIhh1xlt7
hqCdDd3PU3phEEn1/LtFi6HpfENxuaWpj2nfOXhGVloyXizsFIMVU0B64Sj0enMX
0Ado3HFuia2+Bqj9M8fkiZQJQ2ZIUZV/zPhHSkxGHUCVHI2t7n15DGc9d57jBA6p
mDYwtN0qf4z9XYIGUbTMdC2s871Hw4Ry3U+t24LfJIYIAQ9xghoj5Uxdx3A9aDfX
ZnbbwZvJ1Wsldh+fIOIL8JsG/qnR5WYUAhIp88KLAgHdm5dSmk++kxuPXsd+g6Ar
qh147esq2LzL6kGk3jrX51g8eYR4Ei3mdJL4XJ/zZMOYrdQQ50oqTsM7TnO5KQNl
5iB2Mba6cgTYmokAfwO1IJt1pqkPO2nDigTWAO11B+bTpFs68OII6AxUVz0MVCoO
crqTPO/VAQ2gx4XC9L6hPmswEYNJ+Mk+OCoVcAbcMqY8AJi2MrnLHmXuPiyfaK2T
+oJ6LwQuwufSINCGqhsLWZFoz76zhM3F1aiNhfaabnuU13T8SgvYXi0k7LbvlX2q
vPGlPP3Sg0AaCZI8jlHmq9H7iXYptn4fMZDHzMgdzN+bALTRavkbwDGrRJ9NmrJY
YSnpYwSsc2KV0d/Ng8Z6RClf/44IzUPx+LMilQ+cG98IjM5EKZdao7kCijGYnNcB
ByamkbkJlhuaN4OvaCynI5RQaZqf2VGi7LF90m8AlO6+zTSDcSEERA3mpt6/xR8e
/2TWbuxZXfiJHi9q80XGjOSB0n3vQb2NRQTiUbaxqa0rDVYamM8+aOZ5mxirRaO2
qs/qWt5Umid1YIYQn5Jc0ldLSmBAQyPFiJciHzKlcNI3mtDegoO8WjF0bFDk37V1
Xv9u30CrPaEChQHDzFfnR50ztnti5qEoNs535houJUjpA+uWbTXJ6wdfZWA9N2j1
3kqzqHtrl/R/ORiQVueYNUx/T8IzEyvbeAiFGYF0sn4DyLeVK0dmhBLFfYbhyCBM
XLWNOlZfzc+cqHUEC3U62xRdDtw4/TAYEuA+/ZLfR7Wa2Qoap/VNQ+bIaX9D9WCC
8l+ejtermQD6jf5ReH17u+XX10u/8j/tEUqf6UwkwPVVViQXqeLHERSbqp34pBIR
kfX0wofZ/4wN45qlF1vYSHjmT26ChBm1na28FcZnmV3YNo/yYMAmmG4uKxnOlDNV
iI+2QAJKzxhp+GHwTAoUXAlj1VL43uEPEygEE8ADbM9I/dzqAMfJrfbz5gQOlruF
i2F2pRnUFfDN1Hc9lOgf2LqYI4huSmnrBo/byWhaRpApotPqTkcuF5q+FlxNN9wR
nx5hxkumMNOU2oneemrkLhBWwXnudikpYrbR/ZTuiECFLNZ+7p9oi1FurvULHdxm
767S8FmoMAQUaU1y52lXHY9G20vSt5K8P4Lhlwe3C8v90vloIcosFlzZjWoiQa/3
YKhU7P1r58E120FOjFkM9pEfXvgFlZEf9E9RbWJOkRurGn8s7IcI5TePS1+Uvxv0
8+5FYiAlpfaX0mtaAuxTybYBqBDkYVcdFAu84Z2Z5Wg6aGh2ub3sO0VvyxIrt49H
4la95fskYM5/S8pqvmB6jHPB11IXHdegGdhf+d8qofauwtzrVsDcn/pYi+xBfvX1
K+dG4bnN79JH5LPH/3EHMb2hBpLQDLFHNzBOOaIxlmEH/gdyI+IuROIAx1C/47z3
6bGgCjvfHFXavBfaNKhG5KaKiz1effob9NRamOUtTx5BR7dJ7+mjwcpm9fL4mjmb
8GObzi+KBV2lrAmAktx2OAyoJrUyo8V9mbYOFXyArsjOsufgyXeibPvwmRSbHltz
wjimKrYAYmtzF0x6Pod9RyD7ZJCiaSvtR6TaVExLByUrCbUXDJaLd9K99oZY+PL6
v2BidMMdvXxhIf5KdudrlkDQQgkgPcmKgJWF1OQX2JC7HXggDWviIxFUHbMJzdcX
TpTna8tv5GOQhfGvPBBUOcVsmgs7MkHsiafaNerDpiTRgi7BtWjrd2XbOSmtOvyc
t3B0bPW+h7g3bDNiom/qsHXRZAvUMiqeDaZ4GaZOqL057kRkEgalA3V3nL0QA8q7
PtChqf0Gaqt3JJUjFl9QvZnDlzsrkuPxgbXVUZPlSwPiFZa+3yx8XoS70KV3d0pX
Mlny1EFfmJP7Wcb8Hhz95zakC2x6+ncOwc/ObagOoEwodbo0JACpOJNvkFKLOsoc
tHUMUQ+EtHW6wqOKv42jvFRYAxtLuueJlh5zgU+1sxjZqDyM08y1kf40dmoY3/hb
41XVgYAbna85i3ZlbGhxWdugnKSj47b/aDZdAzogP/j3Dt19cwFN3890Vk8w1Xye
+a2rp1X9YJ8MfaUFQiXjp4j04pHA7+Mj1iqrAqw2vZG696XYUv1n5E+8YaYh8h2W
ZSsVGPGtQXjV1yj30tte0wLaxMCXvIo1olfS0h1g12BkhILDJ0jf/87uQ7z3aPSM
tuU769fEOiGgHbNmWQ564Z7UoVMcmJqVPQeNRJMsxdxEiWFDGO9JsiDdoSBSvF4H
9fla09sfmW5s7RefhKFRSf7Gm/yBHTEeA350l/bva9+6PmSGqnLVnjB91y6J7VV0
AbmJ2FWMFzhtWiQuhd+8lsc3/avdB64Sp0dFMmOaMT18C1qlxV7ACwm2CzB7y9gc
EyhgKSFzgph1GBIq2ZdAKp3eSSrHAY7mI+4R4F2V3zxHPaEvI79sHgXDuglDDIgY
+6dY/qRYDwCzIoewS+31byXWq//JqFCtuKQ7O8QblUjeLbHGUXtEiV80mlj8F6j1
WztyJu9AkBgBhpUDcq3JyB16qLS3ZTrhgOO2sTYlW1d/q1eDjIPJ+DtpXj9YQj5K
2aqj2GqjqG89wVrHEtZBbssEkLaywIMhtGCIhb8eoXMJmO8DislxXhp4yirr6+PZ
YUhc1l8ohwYcn0lFGn+Om4fS5ahqcBbqmQ6Xv+cFKgp9SjQj9+/6QbzmW2IFtxiU
0DaHHuhCZKKNKpR8GSYg6Tf9Ryz5geE4YOMgQnORSgyQEBZXyejEhLP4VcvzowoY
wXKIEzlA5RqTNTNqxVoSG1BozgAYBCZuMH8oG0FWX2eLEHQf9jYwwTZpRloCogzw
Pn4TCaEyfedSz9JH0sif652jP/vxNrhvjLal4GAPZVO7U/h+qbhHTIUqzug4h8zn
Xs0RSD+fBUQHQ7vGjPgtMrD0Sp7dDA3NIWbLYPv1uQycI5pI7BK2lolvcpDqiPq+
sWy1sjLofbCZg42sX6M3daz20ho0BBKWeDoW6FXArh7RyIGnL59KLKP9LQAvITZ8
GHeepM3ebYRLha8LyQEP05GflI6nnk0/Q7PCJXNuMECGDA2OlihBBbNKQZoORFJo
2KMKSnZH/1JbgNXxklhw9c/DEbWT7RFH0CbzgnUJjDv5f9+mteVgCMv11zUbHiaH
HgNTkmVAQ1Dk0L/o5byFUyVbj0YuCWuBh17+t20RDdwyLTOlS8/6p4ckiTQPNBHI
f3FdkwClsGMkObS869hhlWDp+yJC++GI3tWnS6LeW42QaxZAQ31bkOOwF11+hVjF
G5ZQfBh5Q7dhQhjIoCC7BQWr/3itzm06KxAkVQvwzsnC5zvJ4wLJcJeopENtcjxn
Hx+EP+9yhVEaAwYK08T0OSBXiN4UDqpOSkNo4Yty7HQHCWk028fbBZnBVf0yDRl3
ORqT5Q5WD/G7723v1x2ODop49ELgK92eZxLzyxkzSON7Lf+uYCWkF2WO3Z5bvnTi
BrkYORyjJAVlqCdzQCmP4liSYht9GFWNRrTyBTnonvUFnAoazTzjQLCw+NCJ2mk1
iGWveHa1AK5xrgKWW+UNTpxQoSXJEqeN6ywxv3JAzBDyHapERkYDor1cXwh+rwZX
ViWOlwNBHDB4zNLklFXDSTz1iFmPJf8nKrG6KDU9m92AFodcWYGuic4AsLk/S7f6
uXYVLtAHLDFV5Af1zgEXrtbm1XCQPYiKtd+Epz4N/UVQ36lCsLmdX176QS2U1Jx+
NrGa5iZcrl52SOi+KafeJHr36SHUUUufwrkx9jXyLe2NtZgEg/iPzpCrIYBco1OK
5kBF9xYhCLmZgNy3z1JZjNRaieNI4Mk+3V35J12u/k9skzkvUeX20CCQYlDuyNQ/
lfdUrSyG5TokKu05lmDpecLeTTkPQMITnJyQ0FAKa5SrzI0ayCemWrJLrmdqbxTq
0MPvYNxS/3Q2T6BselZtI4+0WBNgVLFavvNKDWXGWdH+aFcC4nk94yDz5kGS269N
y9fj8W4eEYIr1i7hooJZ311jmOc3n0NZ1psrBrw6mGSrLXLzMGrFhdIJSHtV5/eK
yBvtRAhdjqpc3xlSkGaSPSPNJ9v+0hyLd4k1JhRq9dCJ5RJX4NNv2lj58x8FLFkv
EgdQ+OT6XXv545uuwN+AXgyI0QtrSP1gMENedr4H3aMHNqQNirhSb3bWHPGxw3PQ
TLPr2GIDSrGlAgkxQEiKT/4Ylx9dVZzrBSEgGq6DHYwBYIGW3pjMBONAcF6NdUES
7pNKtnFVlauXnYcLWZMHr6SdR2vMVxoW6VcqSAwvizmgmKeBIMnFZ4y6swkGDhnY
IfYhat47aX5L5LwKwiOY/M1HiRjBUhVuhAL72arCn7tF5EDY/vhKyoAxdJF+Q6Ev
gRBga3od5BHIubSWbptbMKyqjEGbMq9mN3ZM+nYn/Ambc69N0clMtFtSm3G1pl+S
ooloqSp6eASK0Ho+iaWv+yt7vPyy5vgy+cRuXAZfCwa+PHkrV3vb3vfKQ7lT6v1W
3EYWTZ5FspCMmli2zRTb9gJGrxcnX6Jhy9OnWTx+Tqoze7U2Pj54ja59oyFVDj2u
e/LDCnk8eRLzcQJ+MVYO5hKtHI1GLPzsWh+3Q777bUiTkuaz4lY5bOeW0gahNDkp
6lb6c0HYjU2YqYr8CcR64hpPnTk0BeVORF3SBr+CnyGxEUEYEAWIOdVaOT+iWEtG
Stam8LyxCAsZ2XaWct6sF/cD50foEyGGmj25InQYJ20x7+ghm3MPkvPv4NGzlCcm
Ms5O3ckXv9RbaBZgJWbrnd1iNuT+NSIvAAPFGSsE9v2ZTQ2whVGegL7aRnMZc7CB
0vC/7O9Cr39Gwy3Vzd5y4WLR3p5ps21TRUe8bunXGUgqFonVAPZAXbgaU/lUuQgE
mrk36Scl2x+a6srzapXOptZ3KpfTdeTYu5mnVTbmAjQHbr9Vnnn1FZYRok5d7bpy
VIJRmZuPDo2CISDqGHR9Lo7wRsE+YJc5FtuUn6QmgW6leQm+D+U8Yl5lVjBimm8q
w8jSZb6S+FsDXMD+4GlIpofg+p6IGnZUNUfo8S23J16l9Y4TY/12LbaTrqhyDZr8
uO/1uAwQP9WOBGWCbXBN2/diz8FJPYnYrNikxxyGORK0XLEKuDgZzQ4ckJFgkFGn
oOhGNDEjPjAscq69BpjY9LHcoZun48XysRvVR9YnE+8yAJA1VP1bpm6QGVnmcSB0
DHSNZppnGooiOp4TFqcfX4weNEoREI4eYRVQaoqtjXMw1zZ4GLuQAJZb/2jUV099
ytMmlrxt8b6Kb+LDJ8Y0p854PfElU25FIeLrewndBFxd+RtnKYhYHOsawJNzkeda
F/fO9J09bdaQxLbvI0Ghcs6FZSY27c8hyc9URsZDdiPLhU47N4c4GmN31NzMEpB1
i5myVwZg5uWHiD9gLvJiPWZO0IRsy1J/nh+bsEmWdy+4rCaLXB9fyEFYrU05wtr4
xdA1AUvv4Rn7hnyeadgYxTKxvet7HJhW9AhmMB25O9S6KJz1kZy+iy9SAdN/yV3V
z0EeTRqnZR65TO9PsgEULEGj0/1g2TpsS5SUk2gx1C4pTGdFsbcKlartUMgongQl
JB2xZ3Pgtg9wqYWgHZpFPuhL0z1aNQ+Rmth2Abs2RsIsa7smiwN1a7zWTqlHoC/A
YwpwvLb0INypNNkeI4IpI8kbV9XTGQjz63pJm+LRS7Kb24DHEzc7oeHJKVufTihr
HUhwemp5LRv3xub4e48ycjj2Sajcm/B4QXl1fFkeNdWz61Rk7bYAVkKACigMsGrF
Ju9SpSq2hJ1hJg+bd+xy6LQhDIVvRbkGrj8brliPQA8UFW6rv0hVnHnGSD/vNXXb
xpU5KOvarQGZjtflet0rC9VY1MituMPxdyVqOMix7Ylt1SDRwiSoYDXn2mrmPYnJ
9ii0qxG6bchW4zA1oGdWEucJdd5ku7qOG61yrRYbXd67GX/gHb4KOn70N64LKvaI
BJdPlmf5E9LpCRiU0i4h93oR8JkoJxHYBx1Y1PTlywQtUYjtHHUBIx8au/f4xkkP
hWxot8C0Efi2uLK0Be9/8jkDhB3pINczJ+sCy4Si3pcV3TTMAMpqtW94BvoQww98
PsHl50SchonjsImDkqHbfSvF252uNUYganpUTojQyKEc1MaeLT+NvMMeQnCgH3W5
lSYMhFSCpXtJr1waF+lC2eRlmP44wkAJchaNvWpd0Ixu9Y2704OvMFE9nAU/fN0y
pAfUvBFG2wXTSCt94kBqFkrBmBAngbriehqSJRUCaDibszwWS7jcHhkkixsduPfr
dtRT4SHmGF7tS3/tK/lwV72cvTZlBTBziVPAOz+Xf+25Yz+xGDtH7EJoHXab10yY
7gLypuE8j4dltMO0GqJxZtM21PHuguHZM/UDVBL/BCfMJKQAk4qe/ORXDRbQHjbe
dH1ZQUgIG+zWxab+AGNR86+e3v6cG9W6tAfZELW9Wv9ZTu2cgLCyxlq6rEQ4KtK+
yTk8Owzak4RQ5G5EdutSt5Z97GvvQA4vh70UF3XYKCJhyRL6aFYvj/VWckbK/6XF
7XpwtPaHtPPP55h0ToLfkigBlesSJ7hFngkMKKd+3Mg7Y7RtELwry0ZzLaov9tS4
aqr4boXN/VxmEyozhAfuxF6yZ7wSbLXl1aFNbVJ2mB0mZsUGgK9AgeIhE5GYm35R
UShKAtKHdl9Mmw2LXow4qiiQlfGQGGC03DzNDtlqwLII+v+A5vDad9WmuT/vcSl1
brfHR9u2qH3trkqh19ik31/PJqKS2GCjraJPwXauJ4dEg8bG9ljIgHu3IFZekEBu
7iiG9cgppFgNNmnKdLMbamPI8Yf1tU0Wyh3jWmL1XiRNaimxarr6YrLbwH4u4b4I
XgQNb0PgND88ViUVouvOboIym8wch0cx0mxUXpzMZcWj7dDXJ1V+ssmP/5zNIleX
ZnN55S5Tg/bIZR6t72sz4y+jiDflm+ESp9DWpTlbsYduETf8440S3ry0wG2Bx0C9
vj1QcoW4hQFcYPKcK1H/4K9JyrGwcjhgzXYGx4l9BHeGkmIal4t4+a/z+SSw+5Ws
YhaFkObLb3QMhdufD9jBeh2a7//zq2zj9bpeJzekwpyqR5URvxFXnl/cQkEwA8jI
eJGftVB9MMputaA8DL+oUWaPdB99V29g+TcHe9Ld3oxcck1dtn7QjzAi8HVRQYZ/
6FUnRgVGeFbNho1ZlVlzIt4rQUFfpDCUCkTzSHjqNZcmSLO0ihNovhYWUExnLLoK
9+4cfRd95H63ULrQTYDs1sgDJqalXpxRd+ndtY1EO6uW2H9pp2MFPt6asRrb7Y2Y
B/TIu7wFbMESLsqtl7G/sr5Jft+dBEGTl4XmPMJBKaJ0/VtV0/WiZdIl/BwGCM1h
oJRQMt0o52khUM9NfI9O2pGI1MbnzW+vU88JyvtT338wSXx7xRg8m4Prw9Zj1XD8
m3UsjyQAUtN0N4LU9imxhICUoukdT/Q4QsT7+4UlKsHOxXA2ydCSQt19scpm3DOI
pfzg3ee7EU9pFkzUn7NPV+OhKpbzCM9LmGXiuSva7kdlEr1KqpQ4JnUXoGa9vyLE
FccFc4HJraP7NtNHeAKWOpz3SUE61OfM7dYIB5QD2Pn9S0sFowFVWtsYbDLKmVY2
PTfvoTSkLcEgCDfMJXY+AIh1IrMu/Kyl0/osZ8YjXhDQCbjXtPR5ObrsKqHqxthq
uLp5VQ+XLEyH6h0lYVGGMQG7DaccdFcr72NyaRgbII/p0NBN9L0D1ydpzkPFkFGi
Azg3h/hr5uLa2bcTf/acHYDIWI89jluNqLLbwsz1cKmuOkteobwl3W5v/9nFzrDK
SjDn2YPx5GDpakeulQ0u3vTYMIuT5/jVIx0V9DOQscBPKSTyzhNDglGqCZlTuG7L
l73N3n7J2bRwU46B058PyFoXEl8tFbxhwYlGujcT5ac53JPDf8uocQDNdtHwG2kT
TDQnxtdASAYYJb9wOYSWrMIXWvlwFrWT40ueeDjFGuPb5sA4NNAJ6OBglDe8VRc5
fsi4RHkyH655x07pCRDuBPUdlDqustcEIhmoWo3qjZ9Ok0eArvOUjIRGKtdCKObH
Likhxzgu6PDVw8TcsGoD4e11CGnEiwKF66H8k9FElM/bY3f7Ll0zU6ahxXlq3B8W
7IopLRd04vuoCeeVGUe4NAuhSsvNJajrPT7R+Ax6Jpd58rwPU1klXTauJip5NdDy
AMjZlwnYUttpd8IlQVsfR37IXVA92zpkpL8dCLskOkrKUqnakf5/EP1wj9DzIAsJ
8hLFhxbwetY3wztSjn/y+OPtcWjVsNiUHFb+0afiVBLHrEAh2DgGhaCpudosScZt
KUbLY0pyvPKzp4eQ4W1l8D3HgecpBbkAzZxJjNYjXcmgHZyYX4pP5lEYUzIb6098
VpM/RPSIQLUxXNVN/I2FxF9ot4RPkavoQ3hjIaIGD3NMc6tyI2YYdiI3KM/0hsbp
Cco0F3CEw5rhINtII5GzxqLdbYOnUuhPLBf3V/kuXu7dhJwn4X2KL3bMYBPYorqh
MQCcBLUuwCYE1IvuaA1M2lUL/B3Jp2YIQur5/HF58wK+gWb/aol3xWNztgMYnrVY
cP5L1ner8f+aFMX2KWMyxTPovNSfNdSEemJZ4OwV/jODe96a/ZAw/1sqGt08Mla/
0wFZHi/H6O4UZPgvX3AW/6sq+AYUKQ8itkEJqzMuRi8R/p8kyleegNArNACGiTjJ
1qAZsLDeNLR2T0zq6iyfa5O3WXE0qoBC2rAg73PLFuwAwd8/IBvebbvfSfBhFDJY
Uai/eTK8rkLRPc9VNIl1TmQBpkW14m+RVE8UQarcQWZ71h1GuejfW2CVMg5sn6OK
eZKfPtfS9Yhzwnsmn6W/krAuW44Nok59KhxYOlBzOWjuR2YIxzSDCc7zwncvvltG
HGC/Z9mFBu7do3XH3qXWHzrlHKqPHxH6K/kWAd7+PIzGCXOiYWjzOzSTeWSxKCHr
OM7PXhrzNwQ4YfGeQ7iqFkUkS1V2RtMXQc+11YERnu3lPSWF0/TGj74ILjs50uLw
CdPzLOeOHqCm2rjCZFuMI+iTgPvX76yqLM/r8RyuDBLd+0sD07MDAlm4L0EyFPWF
7XrhQ/8ViqdQnZJKzEF8/x9uW87C5dLwAWkBaFD7yUFfQfYwrYdHHpTtZ/u2OnzD
v/BIdtCgj6rYblH/BnJobxCLlBn4BgMeA5zdlPz0dPhzwbCOPSWbIYVS7stov7ZP
XO4XQM7Cw8ksQlKBWOs8g5amF8SH8gYl/QUhMG04ohcKYxvy8y8MY7iRedkYK+ep
WGdDMnxHDAN8GItqqmkNvVcnf11R5tNNElnBE9IRlFRAIOuV+PakTPjhsmqaAjpN
l3yQAc2/uTzzvsPGbmQPvECvCjlZpPnkPtZ9Z6gqkCWHPTtNyZn4ypQRbQZa5VvG
ZnMvU/cTEqTJKiBC6KZKYa83nlEnC1VDa2OZ35GGx/k36x11SiUzyCBZk/UlojAe
9ugeIHiW0a7VxA/yr9nO+hiCwYgN2QsvfcyE3rLjv1G3kMvA0GCla5Qlon3gLOTt
tgqYMBBJYHz1GXOpRseicN09elhn7PvgFHhab29vmhh/7hpKSLCKaRG4IKBdgnU3
J/6Cvp8S+lRuqgeUJx5vaQ9EVhiug1XYloziy4wic/68H1+zfdua8RWSHIyADdQK
6mLvP+TcOmb13ETrYaUSjaWbLZdYB9noE9Lgo+xn2vC4L/n7sGYUD0dTsk4je1ZE
dLHVTsm52Zgye8kc9m08aZqddtQYca5OuHOv7JF1XwOBhtxXF0nkDHqzDM4gUfMp
pkTm0ueQAdQDPQoMqisjOlHQmCUIzGXVHxbXuslSdFiJ3a1xtAk2zTChYfdFu0kl
TgvHm8HqjweJVGP2n6UJsLOG7OgLY97r37DLjGDimi1D/ckPrk26RoeOdvvyAkcu
/dWF+2V2IG7aIwDpKC+AmqeNhNm42B3QdjZF8rPEQ7VdNRy6hEjToQ39VZDpfapv
O1MWwIH9Wvmy34PK2+W8MXBx40N56tz0OyYbbc/OPm5sizndUfhIPBAc1QXUNOzw
+3MySLYHLY3jwEfVqKGFtdtH3w6+gS6Unhi4CO+j2Ah0SwqGEj25cZ2Wb5d2Uluy
WjLzQ4p1nBAco/MGZygWyejsVLXrl65UYKdiH+pf0NGyDV5uBi4h73wZlxxDghDW
vadn5AAGNtC/nJIWOMjnB630+BjVQwSOdHzx3JeSZElgpg1bQiGZxGr0AQroVuWk
Gk7Lc2wXFPOjaK71uO7YpzaCnDpzJIRcqwy+HimYQF8vDV++EPzQT4chtE3cvfJw
2Y/3wBwng1+aIfxNX90+qjb6ltakNAtjZKb3anuAVgfT+CKvaZjKe8rNntDD9Qwd
yQ2X3WfOHxeU6wu5/0di4B7XTnuCZtc6uZQVmgPBXE1lAF8yDqniQowAhcl1gcqv
zvwzFUCk2hWb9hFzDkU4Ih9FWToiqxGIhnXw4O6STmljkLoTYEMO/FkYTJSpT1My
zwNgmjBrgvcV7WUMS7BS0PqLYl4+mc43WTSBJQIjYdY4DwxWvw0EWncDR4MG/cej
pGoyEmK7LCQXA4pCPIejakyl9yRaLk/yJaP6Akrx3PhJZla008juW6dS1pBUw0QF
PWkTmtof1rKgPwOPwGxpl00W6gM/C2SedY4rcxSACX7GYT/VAbRs8O2ccE6wjXYW
7Qv1xR/MerQ5xQGFBziejCF+MBEVyB9a5gnIvsZAAH8Lt1gyNza9x3l6fTRqQogQ
w4AEaixS7Wq+i9tBzkJuPh0q/PO9k+QCuBgFLW1Cr7nPQR40A6dnl+PmjLND5Z/u
GaiCxEPqGX2GfKG9qmQq4oefSq8i8d7G93ygcZsow/HSw4RbcXlHiqr4ab/fzns9
ayk9KLRMKwWf5Kgin0paPWErNqM+Z1HeHvCkbZG6SmYb3MYYmdbNO4+V8oNYUIft
+KxxUji4aWFWYE3vHLXsKgI3GgRrk55ClX1l+BrMPp6pbi235BIPKbT8i3Q40/E3
iSEI7yHH7rH7DnU78rQUFvrB3raE3I6yPdXckhcRwVfFoRQ9g2cyD72oe3cEO4Ds
gwx2DHlDUNKqc52D+0IRdvENc6YR6l/WljJpg/J7oMuIjxBDHleaoLlAB06kO9Nw
PfRV2FXKgQzSS3oUJGvslGMdEFLjZVHdfwc60X5Z1xn5ToGkd7ifcgX4KZOYXUYK
tJV22BLKfaOrytKMw2v1EnMViU8t2/Qa5wVgeW3SbzJb/meOkubWQXTnHc/gS1rQ
+7x3zjnp1ichgNPahXw/7qs4+1GSur3jTA6l7aaa1VyA5hHacrdyWGqFJTi5LONh
Jtbqkq4Z4R7i75ip7Q/FdwS5HLTjSGCTHVc2N/GgsbvkP47zllgg0sTpKI9PL4lB
OPO/QVXfa+PidewVqMkkaOM+yvQzCWxhUWi8ymL9kYZgm7oR1MLVAKQiQ84cDToA
1WrKrg44ojmdM9/k55Dwa9XE7CAJzCt3J2jzc7ZJfad4pTIax/dbDKAP3W1Pl3RD
ljehgCxFnq+AftH80Vt5ExF3ztcshnbEchAWqr323VvaU5kE6DOFhiR7/UJhq7tp
bHpYd4EpZWgCnTVbciQ8dWhHqI7l3PYsCVEvG9VYM5QvrWaEyCXzwkMILYeHd2E8
eUBH5T5h2UkZBLUwI9cNSZs0ohztdXN38oTXIku8YLqLifGuOBWAdjtPWW35KTfI
31dxlLRfvF/pVJg987NLyAMv/0lkTDop5S0OLBfsc4xPTPF1jiI9RUgbZcwufX7E
IK5XD8jtV+/cdlDoUOJFZlXLyw/L1g/4YOp+JdM4URlUeqPNlq+DmRvf/tLHI+my
iKUXksmUhUdPA5rWOIXkZPmUxA4ySo8KhUkfImlnAgluWgml04Dah5IT9XjwnWM7
82zPWHs5XdFmWFbEWKJi8qSwfV5473SIS89Orp9299ypz0+xI7+NwXKCaxF/yThp
WnbhXBlR2Kmk6vwQsu/nPcbjX7nsJcFdDFlVvJr+CcXBjuuu1AkpEB16lfLRp5wO
YwDZmE/6BbCszYEFhaS33WDduaRtTw8niEqPQ2gHi4A5ol3uhYh+fbZ4s5uaYYgA
QkPzZ7lAKrPLdy6reoa8YO0zy4JxRDeBm+mHTUGGnxryFtqMoe7oalNIcJbv94vG
Ofo0nzuSPJ93sjw0jONz36VhxSQLnv9gb5zFwPHqWHp7VbnwG2WMgPw2EEafQTBj
O+0Oab7kswMG13j8V6LbH3P0GZ8nw6UV8w78bgiAeuThmFfj5ffz4jUQUovpLsqI
Ohgc9gwjfj7tI4la6KxB+MhCrfKxFRzsGWZ/VJEfWK+mDKMhXaMKW18k5ItmKX9m
EUXxzb1ze4p3N7kB/zWpq8RRQbDXqZHKUaH0dCpLFnnvcKw9txYCZaw0F7OQX9uL
pIzGcalBfmh8eYJ2NotMoZlKhqpg9CkiUzTHxcDQDpwXaeNr2TfzGjEs3Y0pc7UY
2lCSec+wYE3WTwdgk7NscEaCEL/SAxxk3x6tEjvG/LVosjfAtVr+9ucMXa5XzNvZ
29sKV9KWqyRdYrdTpCWhOxleJT74un4BfbanadcDnfoS7E41NmUthj50301TtjaZ
lNzqZBXhPZ97dLMPMZ1hs04kiJVK+bhyUNeZ/l8gZ24noyhZCuKgFRRkIsDZ+GwK
qyjkpu74vRgQNLAmGkAjSxcuvVJImQc1u8lIenX4PDx4zZ4zjgmiJBYe5yOf1UUW
z5BW6FtHLxi/fgxEWjJCna2GOTTf5dX/Ms24RYp2CHfadhuzvCzrsw6rPamKUH5Z
tp4iv7pVwnQ4PEH2Yh2MRH8gFBdleyxFp/NLE0VbSpbBZE/m2j88+hRK2heusmpB
C0xUBiL6S0gfy6UmZtg8z74g73iB2W9vbMDGiOnN8JwR4D3jeqqLJCqXrugh/f9L
906hHhL5dDiI0rpm1m+DcKO7gY+KdLBXowttjEMtQ3NQL2DPadRpYeK0v3RY0Mjp
iq9LNzedlug4pXqCVrqgbpBlhg4SWS41QuLk1nnAZZ6JN+d8dyg6Gf9Fv5mHmCkU
B1diblfdKd/yD7fS8sZxR32DYKe0JoeLQ3mo3wBi+OTZYRjc1ow56QyXxnP6/5EN
YoTlw8xQnavnRuZpFY/yk3CytOJM22ypASGCjtKAOgEaarxptWO3RopSJLdbRgiX
AzLOB1vLTg/ntKxjuAlc47v19iak9LoLAI8JKVJNn9f8Ju77dUShXgFW/djOZRfe
9p8tt2wfmVdLkZDYHeDVD02xbc3AX+hFkOnNKHIUvE5QnPt6TbKWOef/cZnrGZbp
dNtaKSOQ/TNKayTigGJJ0nPGdTHaDduvGaBtVkB0DxBcp0WIzYIlL0XzlCWorjln
Svw28VeokXy43AhLiope2eoZSicHe5T0qBpEkmceDOG1Th1eENCpujfDIalwNXJs
cprXj2/kutLaWLK26XEmCcc2FCPaqQamIc8vaR264rapKUIO31gTGhK9yPiLmzKp
ClqgJ+1urlallrpl12s5l0Y9NvI1sxbXbV3etxOmVUGWdVrO5hxNY74CB9syCoWl
N/cJekwq+MeSM+F+Q1y4x4giRl3+J4fEuLRBIKRYdgw7rQa2VzoENyHsd9fF4Hl6
yWPMBc7Mij/dpysrRA3j3F8h+X3fwP18KuB/HN+eX/x5L9dMi6K7UmQGRs7Hbq8p
yyBwK9OgKEbTyfZZDJaag5UBZSHyRjLr8x6unify6nBN25az4tv3Y5r1/V4XhMGy
Cewv3gleFZ6sjSKlf3a/E4X/GmrG6TWrNWv1DN8+sLiNcRcAnMMLHh18Dxvh5zTP
3STOePuE+v7KkjOX2MIXGoY1He/7iqXA60sw52SAaWdXpCw2DYvqinzuevOdotbG
DIN+Gu0XxzZLpKLNU7DOu4sDREkO+LVz/BFPnlCJdSAI9CgnPAJAWVlgGa0aEh8V
7RYI2+UbPCCn86c5iV4wyevxCSly6W7TZrhc6Kt2BLfuz0WzA+mNdNqKXT8tmFJZ
u1fKrfqwaweweiTq6jGMMfrfOSg/YkuW8aaKZS+WnYAx1iYcO5As8RKzFGBkHJEY
0p61pMU0+OTjv3bC2ZDa4X5IimpVG4eae0ViZZ3oBs+N1WQn1dQNoa+LDaC3S9dZ
A1L8m13Ze/2q/OQMrk2ajMTDzQ9xOvThxDCIxlYPbmNC0GPHtoTzP7qzk00Sktxk
vor9mqXvaO4eBuuxMbAKO0nbxIezRNBiDNtHTC8JtFFlcMl9ChpwV9KQVhFfJyBj
zbnNC379K+vMfhO4HZu5crEYzg9+yw60OovcCQiteEh4tfSQwf/MKfpvQR6ZuXOu
9jIy8h3xudfU7RrvSurGpLu4tJVO5zrmS8sebt18ScRiOQrAZWZd/AQDPzXkRhZ5
2cC06gBQVDd/mIovRGCjDgy2+3klSBtq+GOQTWLR8N/q4GqMnbW+RZdBstN5iDJe
M0F2p6rwucS20IHUpgUosiuFjDC3tiRAb4aNQY52D4bkt+gicloEXxlyKIspYAv5
pPrm30V0q9QEzFBzSzZdtmj3v2piTIkX7f5RDINqOFo+qUfsXrB4+v0fil2Uk5HL
KlWep41kL7jtFV/yQ3TZG6FJ8E5evXPGgF63ogANNNOUYrBrzcFQjTBO9Tyq9HS5
fbPLp+MVK77A5fNNyyQy1smHcm6iGA/eIdL24O7CrSPWzkJ+aqDCQJnpR73AYSkz
Y/h3ARpr6ZWcm9uHbGAhXh27D0cYmP7FlIwykBP3FRKaNxSD2ch8BliQob0ncbi3
BtiNNlCQZPiKaD8JTtlHupEIOah4Uz5HIPpGvJYegDA00/RyXxwdNIoATCe7AjaP
bPa1A3Lg1qm82dttTeDWmjcVH8zg4nxmfJKyJB3vB7XDDagk937bXzwhszQS9vxK
zmAaUqqPQTUf2kl39D0AApXYXBTKLtyvQEFlPffD9/hqyAPQc9L+O2piXKQ4Ps8l
+CBXXpln/iXNnHP6jNUKUK2eKsJ3M4YQuC0gN3dr8aa3sajYZ2fB4mzbcvRt+pt/
RJLhyk53RVE6HHYRvVfIS7kA6p3y49vWQVIdaeGWcBKmA3e5VpPWIVTe6C2dxTiY
/4kF9gmZQVfnE6DpaFg2r4+KY60gY1Xp6/H0WjNrezF9WEuZXszgLcS6r0D2VdBo
Ssbf104gQn00ag6dIhXKLQt0KElvKyaGZxmptrteXNNwaYznHZcJxvD2uXcVi1lv
0xzwlD4Vqq8CXHcOu/6jRbR0t9Ep98Px28ZIBIDmdmshKOIyKkQLK2gh6Rqb/dkE
a5C/8as2qaAsTo7HOXsMmG21SClXfXL0OUUcvK2Ta6C/Oj/GQm0kQ8QZlc4YtNBU
bznsEjnWs6Nz8jH4dQfj5Hx8bfgK3pFtTS2k2nEFe66ihAKr5XPOocMK/QjH+h60
0uPtHI7b4hDNsnSVOYp1X+zYkHF+bRKH4k+HBGtNZo76ckGY+aeLANze4nx6LQ+R
eIKijCHLjoP6XIiR6Ws9Cfe7BfhNGtdZZgo4yHUNUbDfrh6GBDHV+VrEsuWFuYAf
KCDeo//nAbu7BvC/9Yeu31uINpb3HmWbnkjtD+g4eUb/a9YPOrn6to8iWk4PCYv6
KPfA9dC85dyw87BJR2zOlWpNWh60QROoQsFSg0aWCfH2QBNpItwUOV4yRRQKbyTl
CnISiQO/C2fwjag0VQEQhZQ+0IJbSEkHmYcQFUeyR9/Ev2TknUUrdBmw4jB4OJJX
kEEnZrSvNiy+/oNCag1/GJwpcGRcYqrp5epXnXZ9oI5vjCKQTST7GcayAS7U3Zkd
IXW2mKA87U3/Ot4+XnY3aYKrkKpznzK0BL5rFz2oOTG6emP6o1yUooEUD1eRzxpG
EV7o40rFnAEtSWEv8yYO7raWR1106pLDZEMA/ff+DdFPB5MazTEj8+cYhE8m07bI
3mX/S53qLfBiMNKTUAOz6leY433/cFPqb7aL5WeU3PUjCwdw+iY10a0e0UJj2Zqb
csQDSZCoURyrI1AJiai3p7ptfc386LEKx4frqRgDN0qZtfyd8rjIicZwcY0BOOW5
i7AVEDDtkr9g0r6Q1WH7XSN7Z/cLaEJTuq8p6IVpyqnxLwH4udYcifSw2ew0BSvr
qzEur5VH9v1+EmtqePcicRiYvCxgLU3W6DdcBUA7uzRFuSQXH5WryP1IJxcsECwa
Iztkbqe34bgHCg6RWnl1NMV0Eh6+O6AcboKex8xUwo4G3PKG26Nr2FvfxJOpdxea
vIn31EjyhmWewXbH2xcGxhd3CmMzKCgW1OQXUMubYYaSiqQirxkwjIHCNiA2hRqr
3ozQk6sBMjUtsEoWwfn4bcxMETkR1Xkcxoq7zOIwEGcEJ8MUDa/oKPBvjhKZeT+F
9g6hcK6ded1vl5GLPwOkQkVsmq/nS5Xs+D5QhW1ZCDat3iaRY979f/UCOdwJ0feM
Kx8PsIqzSN2CRLx660j20dKegW3nebhgzXfYE0BrdyjDQWPDZ4+tkuHj2nX1ws9k
RsitE+QxmRw9ovTHPvnn+5def4QWABSV5/JLpHQ13ha0yO4jjsnQjzAuORY1MA+E
0xQ8V2n+JzoYb3UJfBWEE/AEcI//QAaXU8f8QtrZlkW7LIqHbFsfOYYpgGIhOp/7
LMrywZX88z2CpjeoVOj9I4TI7ADiFVnNv/Oa2LVTV5/32fdZRbI23UcfQPWqPrGu
nRDFUm3WnhALuyS3aoSRcdt3O06Z6L8bgk1lOYPy6gLdB6MR2c/MhV4yp89YVsCb
70fOrbRgUcawBmDgFDIjoHmfl0s2Ife9EaS+WR87nHAoa/pGbj+3LPKgTHwwmm+/
B4FNJUwzzfRe3QrNxxkwEEB2VaM3BMylLu5JueNwquuZkJ3SdEFjFPUXQnPYidVs
Ixj8MIylxDYUpq7da3rVHUISj7bePundZmbPhZhnBUHpTrsB8G1HS8lYRhj7vUZK
aCl8/L4fk+ETA9eDw7HhjoAAFFN230fnpVbsf1RqSW1SlXYdrMFTSY+ZLCVXRplO
Rpk3NIcE4Ys3uUlIIvpoCYFb1wRKPynNpOZIifT0JOho5PYqbPGzdPnOGH0iPLY2
uaM1vXiiF5iKVTVi9CdsLyuu6Fh3So9zkY4XAhVHzv9gYSGmf1DQnWgADf4fYlNY
pcjGq+FrTHoao62m3HlS2qyv7AhkMIf3ukh3S6BY1r7X+3DGJAW+crxfTrzbLV1H
8+uncRU3OQTygowDNnhg62NXaZ0svZqposo0VUEt0bRs3lmFC9pLV7Ze0yfiCdLe
lQxiuFcK163I665o9LvR9KZUAQqwq2aEeOyCfaOEMsMUjZTPReQbB5NlLRC864uQ
aEmqGZ+R3zXs8tLR7B9MGTthtT1yq0zm/QaMNRutW03X6ZH2dUpOaVHuck4B5sPL
rEpnoAkCkORU6nAM1kchHuojsnRWsFtD6Z2KdsrJiFCdjqoBfRxiLlqYx9scj5CP
FvTQQe57tJUZ2eAZy3Xg095AQy2Iy6hTB7lcM2auq9/dResXTjXBBpUp8ufH7sZH
RRImjDK4+7rToorlUuRT8LI3SSHHsrmG4yuhcvLfMmYyOiorlW3QLLmHaCWN+LvR
InENR/4divPNS9iaR6dqdIR8sCn91sOB+rkOvH7qHkMaH5dAg0zaJxfnTjM6w4ry
mceh+pOGAJrE3Rvb64fN0hW3KUIiNSY+Umx9lOnPefMLu6YNhrB5wAM4eFWbkZdw
POndNvWpdLf6tc8kl+Qw+PwnsMrUBZGIeQhvFOgolIbLf3+rahJJbA1dp78N+Dew
7AbEfXZ4z6rppqFkAqBveme9SGhzoWH6q+3j1OhAGAIcQzOrCEzXu10K+yzusiS0
8pIRP7sqZuEB/E5MUXe5fu2cVuO6mzGJwynS8v6Aq/Mmi2PxMyDT4wg8ogXWYxIe
WeKKtqxFluWX+Gg/jZy4MBZAXHsnqZZ1IwAcuQN9dJbf+6jC8hA2i2kIhh989z1S
JQOySzfi8hK/dZoI+BegQEtte5RaapaVrW7iZvgCSASeMLE8K0HEiuGKClRWYJR7
xIP94uLjxtXPVmCm2UpqSph39N+SSsz7Vyr/FfwUAX5q3/LBp99a+sLKe5BJLUYY
AjoHbYSCKQ6v3tw0dWsaRSYN8X3BqGHdk6Dq1fubHQ5N3SGYX/+dbb37GPBlv5UQ
heVT4WqOIqXbz3ZfyCoABjQ1qL635mr379/FL3IqrrNtMms8oevcrxG4xPzrMOTV
W2KUUbQO225IhjRpfErE9TTMUC5pb4Ow8L64KR6N8K0pWr/eMHaowJDQQ2CTAIJf
76YUWzwZzgMcHsPzJpEdR9k+VL4XAsWSijuzqm54LLewdiKg8eA7pqLZLeBoiaKU
GBrcl7hsCNhPUh/2APJ2IEBRIPTq5onQpZ8vItYJG4OYisRks6s073KxM6A2uwSg
MXmVBthzTMlX/2mXazlicFIHduhOFJQGWQ7J5pMcL0520yHv6lGoD+gEwIn71h1Z
Y0jgXpGvEV8nz2h8V3Oh6341QHmzdd3ZApF5Qa86HoLcUWruOGKo06UDdsAag4/7
b1V/KkXa2DpPu66OIIuckeLDgy71Z1JpKFdzne47mujDmTbwTwM7D9AUjHPeH6Pc
Jmr6MI06StTFkF52PsSfj6ApxPHRTiA5roOFJaTPIkYHJ2TYSFh1207d1z90csw9
1TqB8fUpLl0m2rhsL7qP+mjdHCGRUrI9r7cqGJ97lr8GPtYn0t2x7I11Um1qw5HG
a3M+r/yaqW8tJb2FNJWims7v8W+eaKFH+DJUj12ogWxVz/T3h3kWt35TghqrB/z3
PVh1PpGO79pVqNadKVvpV4qxRECCSryx6uC5B4EhQPtA2w++QxoMLT5gCl2G/J03
tvN7smdwL+P7+/6wOgNT8CZWIECE7w9TVM0+AKr+G6Mi7p7o2RVEH/16+ZN1M/QT
rq6f0TmEKluhyATK17CmsdWn2lBD4jSTB4JDDzx1dazz4iL3Hv5YMO2zfEEHyEPL
t7ss/NEm9/YH4PAzSYREz5xCMBZ2M+JoPDU493W8+GOITfPhxboWKlKZhgHvtbo8
B58lrZvOTWg2p4BGiYke9oDPWcX9xrH1ImNhdaR0Yq14jY2skn0QIqZJgNRfbxCF
y+6/38zJPRSQWQoka6vYMkJCQ+RXPWapY0N3JfB91zab2PZoYlyuwysQO6Hmxll5
04SYdRDYeu4VXW3n8jacNjpaFm1+ii6Xr7yXHaSR3jxPGAD3lU2s5ZXp1mm1ycS0
hA1ZTmbppk4g8nTgWGoA7oG+faMU0Q1/bL8zoTsf96Ne5v4RTAGByT+5vpJmVSTP
PV15NTg83E/gpHuviDVxohcTvN/2KJY87RVrlR5M4KbaeYj7J3HI7GHSii9UO9mj
KKdIH5zuPImhLy3NyBmpXJFcjAaPYj2r+2De12g95HBWhPOFtLNALpUHzLi2rGru
+2TcYqGzYEJ1lNRcMwl7BrI751iY5A69i12z+PvdiCNjHc/Rf1KdNqofDoDCQL+D
z+VKesZNma5M9rJl2fZptFGi101cfY07whVsoZZx/nHNz1GtWuGO1iiEbjYlfQgZ
WZp8F1xTigs/XHGTnpeHAOHiaO6hU1aCoie5ZV16fLvksqZmYihMQKexUy5vUtRL
DGG3Wq9A9b+eCAQRzJKGFgfx/YOflCHHmdWP44FKbiA6ilrEL+8Z98bTDTDExpii
XupbY1VNtTZpPiOHBiT1IpyAq3c9fvhrChKcwgiFvj1FrHL3ccimtrelEqPglYVo
nT6WhF1nYh7Jbyb0QH/hdS/o0f+GgzmQXvsIzGzolP3xlk6llucr3kLM6GJ0u2nf
LgroDwt9AA0BrqPLs9WXLAY3CVudD70lTxbmT8+H/HzZ6oF0iRU5vijmJVl8P3kh
iMFZ9slUIgq6DqFrNIInOEOXdaYDr4ltIAp0nKqZ9PGuEKf/DxozWe5DVtx4fqoW
MLYz7AeApchVPSbT18C4Hw2sXetg6WsXHWuOkf0HKnKuezFQof2E5Q7dLiyBCdPf
Zqb+QyilJri0eW4i8ITTP2c2pAllV8QFwNW8t1e3PkhAnIzlxjuM3XiRMRgBUZZH
9P/vLtu5MnRLWx2f6PzMDcZuzRahPdYIj5Lnc41Fi069OwoM/Eimf6BrUVqNrdav
cyTIOfEmoU8evizuxMW2ShpotKSiq84rpxmKKDTOH3eLy7yn//vuNSvQQvOxHTco
5kZCTVWrHavslCgH2dL4KnCLcLOSFySl9lL5ewSx+dJfDIw8bwiOdPZPk2J/6ZEj
ViqE2URapFWlkwLDiS33iQiC53IZLSKJMoTB5RkEHB6uyvhFmH2JFdTj8GcIfof2
pFGuYP4gOFFZfZ/jNL4oWxXQ769aBOMBxUO215qs3RSZ/jgHfvPksNQBWESOQ1/f
7ZNgB7VpG9v3YZ6WvzWCIoIOtXhfh7VAkbyHAu1J7plirEhg1g03VAR54BihsXAF
mHbPZddRRZNTwTgJtjffwtzuwzZpFaZl377oN3WXddWm3dQ8LiIm2nEAuZjokuzW
qzNDf/OZ4kTf7W59LlI+o55VoZJUHWC7/NjF9b0AkdrdUzYz6JViLln8osOblg3i
NXHBLZgZHCflmGG74ysSz4jiAzO4IKK6gsjY+c/NA+aJ99mfcIiUpb3901W5J8v6
+1cJamkdvvnPgs9LrLYRCj3BS530qEQbc974+/+cMIYR1o8hagS6RCZEgD6PFS0N
UeWnS0HxtqsrcdEocP1d03ZvcT/21N9HYiVc4ki2MxeHXikXCKoTtehqeQ2Kso+b
wcPKM2Bgt8sIXTttt2L9pB9Qkx4i4Ax//ptRNXfORoj2Gk/961cWbKegzNZLfbBJ
j6UintgnAsU+SHjufyqomVQf24BhbyK9/MRoBM9TuHQPNugI/dbm8LX3RG1TVpeU
LfLSfOFr5aDEb2alUiTD36PRPhCEAUdvcHoKtp6rwoMZ9CPVd9Kf83r87vnMkfiY
0D7o1lAW17lKw3twNgJa/05jFVIzUfQCNPjefZsSCkRUGOt/lBhufsCPGJqY20Rn
pmGxWVTFFtSe5dw2y0Wt9eSnIRFgRUgwz9dF7Wm9p9qMAR6lSqTcuQ6iwlXwoP+C
bJxkyfhswd8zy3vbybuUgnl9Vmh4PlC3GmYW9lFeL9GAHVwHmN983kWw++3vpFEj
R5Rk6ydRlfDNiidbnQiPwpkVXTlY72k4ZHibZOPIYt/kw95nKhj84hbh+1gl5/zP
QttNBWlXpV2P9jXVsemIK6ttE9cRSZB8IPrVA5F26N0bnP5ji+aDTwV/eifgweAQ
/oOl5v1+fpJcmhhURgn2lsCng/tzQ7irQgzhTB8vHYNBgTXckO8zaSS1vCo+NlAk
srDLgBdkIrGE2Hyxtsvn5Sz6FldvOFEDN4wWvIq9Y/3hgbnn1/iggUQ75qZx1SDq
8GCm4DL/gqBgNy7AAyZW6aRncPpJ3/SrpSSG3hy/jxT2cKzzMmEtyiauO/JFyAry
OojtBniIdtGefNoExRUeQgo4ObNdAgOqWbeG3oN1CZuO+zP0TiIyOfXmQL/3Z0fE
ybm0ui8VIfX2KBZiRpufs/RV79DCEUeCczeYL5YaY4zCP3rlCxaehmORheZnsa/M
y952Bz1AI84+DNHTJgbjgX/M44KDBvYCPc046f1N3fTJKFkWxu6GPWeO8yKS0ckg
61+K8Q1rThAlCgANHK+4AdxIycvWSGDx21aoSA39NLZrc0HyI+BtiO7lIEw/KQZm
ZMrN90Ws3l7H3wSjbfn2pJ0klGrbCMf85gXpRz8AJfuzor0X51qCXWqMCTpYmt8B
EBFi0AANqC4C66LII7v5KDzxypj13j8E69CMmLpCfLku28kgfAdhB/9wsT3E58gX
SgHhsY9Ykr2CvKLJCjcCpiAVENjaguqKokFZYK7cr0rAuai5BKi26Oejf1pagFbL
7bGQ80pgpMEfcPGpysIvhFYlBsPXFfnqZpGPRKlCK2hYpHvpPVBaZDJ/4tXtiJWl
UUisrycoNi+LUDMzzqKNChrQ0JBHWUf+uZQX5Bygm2unnfNWCLRVNe+H0r5Qr28h
KvzSauZrt2paUaKbyMxKxlARYHGuenDMj7HTfFTOAZ/kxW4JBtCYfp7cDnV7tu7h
g2mFo9Q5qxeXVoxlClM16NH0p1tKBi4wazzjHKYprsolILthFwo8VsT7N0ZZurZ8
REK/MFr4snOLqnRKmOJm5W4Gn7cG1dCbKyCsoODwrcG6EpBizVXhns3MFQJIHyzI
kj611WrYkHQerfTaTDh3qpelyD0huDmiZBsTeBthdh2DTmifEPB+GmVRNK9aOj9A
v1XF3vBcGRRxe/xI7rexGQP6CSFWbv5vpuLyY3uNlkOOkoplVmrWoJyXJUBUdrqG
XpZhH9ITzmIeA0nzbnOg2hDwceIz8W8Pu3jRzpnf6g03R5dOaYcao/K3YUjphMUb
CSqdpcb4KLh8cKGspfnzoJ9fnEkqPgunKCD+kDaprzXEUno4Rpckx9bh2r+SlIY2
6Hy5Gp5glaDJMHFfiiyHMaABWzJvyK5PHUKMlGRUZz80tFgjZl+JJNFAvoPbdCei
2yHDkTT9EIcbdaGxT4WAQd+6v7RhCqVtLH6ZstizuJEfUUfY3m6eBWoRqrRnioz+
FsxXGaNC1sdU47afs0jmieq8S4Hjvk8+nUWaMAz95inuPMXJ707dVyZbQqNm0xpB
N60cm+U9XsBlIZMqrtZDFgd9cwzka4Y4DZfq8N/vbAONmoorsxiPVxAQvmlIjm/f
k1f10sE1JuCSFoLvervEBrQFwHqbFciFbVa/fMjI3m2iasEhwLmneyt6dBHNTbCn
24/SlLFNVSRN4Yf3vY8KqNfAJZk6t3RgT49qz8dS8mPRkW1K/X8SGO5y/R7CnloT
PH2XX0R4bmV/2duyCeeHA/pT87DcBRi7IX51RQlNufM9fn58Oeyk5uGn8/9W4Fbb
1rvuoGzh+6+oGsXoxKQVIr3PwRpg1SHHLmkuti+6J8xSVofglAHUFl2EzBo+36pN
hVuapUElctx7Dpik89H85sAdd0VtT2g2CDXXbzg0jK2P4zlt448Q+IfAku7uNuy1
RpYYKVqTWchbqir+eq62CrIuGIMfdj9fWHpO3f7AZCh/+tv3Qh6+yEMs0o6djeDP
sXEQCAZ1hDzd0tgOzvnCNtPOLPdvHlD54OWFholkbhyN0Yd36l2kScSDUUbceXzy
6AZK4Mfj4/ppscC8Dv7G58DGbTnqKIwuvN5vPXLGJqNc+NSlAV8/jslQ2WeQPajW
IkcpU4kbsgYESDLYcgmRpZNFAQRSwem9bn55y/pDe53RWC+It5lM9zwBjPZkyiB2
ofI1rTySEr08/6r+zEPssk9bNyr8iFnXW8DMWQeOoqQQLB3pTv9W83Ywru5bP7y0
l8DMQYc6fjeGFGerR88LQiXeb11jhxsSt46MQUOf+6eCFTWHg9VcpkniXUTtDICU
9aGPyAF1CCuflOAnVkTkdYjLXfZPNOOz7PAf/I8WIac5Ufd9zW8qY6YDmj2G+LfZ
4ZONAgO5OpjjDEL3YI7PIpHk1Al289Yc6aTxGToO/rIFbiQMHJL8t8uBmQTPnFPm
VNSRrG4L5YuMLQ46pQJ8nkmDeDyhpc0v+hjTfjVoTd+bZZYIPPxIj/iDbEtx5Z0i
4S3B0kegwe93pxnnnfrK7mKyjQSWcMRUzQi8lxo15m531eM7b6wesY3ye/6iCRCk
UWz4wVUGQFF3fIMXEQlOoKscPlfdznR+81ORkQmZzRR0wpQ/Fo0AfV1Aam2rm1au
fuj5PTvWQ37vaLjAHHevgbACFM3vKHf4qqLwrpFR4Sb2+AZ+kk17HPevHtCEK5c5
k3yG/CjjuGnq+Yj8VLMO8xbSa33Pl6sFPQA293PzhMFjlvyTt6ZnIS8g7iu4OoBN
GBbVIpAB9lhc0S9m4sqQSEvITZLebsfx2HpYtfTkECMM8lFyf1JRnIrS/7uVSm/W
5eK2nnhlV0maUPam418bbPlc3oLouZHjjSW7L2phXvDIi8qmDaqgsHM4Di7Wc0G3
iOJ1trDtAHCaOvhqH55WVu7qmauv/ajcbi16YQbbvKpxLAEEjtVG0gvNa7Fa5Lcu
lJTn7lSryJxqWjmsulZRUHc9EIfpoXtP0cvbC5iGPGVPOPUR6JOJdV+LGr2HVDUE
5pfHsfFsg6kH9WQhGY/nkjv/cYkCIyjuHWfRxP3MniZKT5oIcxGVZV/P1sR7gVWy
Yq2y0UlIyVZo/TylYV9SAB57RMAvH+79bDuifC4EZdVdsFq6RH+iOvBSdxNgo4+R
U2brj22URFXK8eTAudiZaHUtjhiVz9bkqQrewFEQ6FszbndwYt5Qk8r4r3Ly43Cn
hKFNsShxV66wSxzOo4kSRtEXLsmodCa+IAe/ltBPrKZy5kFMXtyvRRdIpqCoYYB4
sy6jkFELAzntzOdCLHfGiRBPLi7gDMue7pvOWZSDM/8lcOpKIAUXTnIqNKjHhjVq
6joKVzujRFpfCJI6t6CciODGEjXvcIDjnK+ndHBdllreM5TYV2VNe3tPR83VcX0j
ZdJNscnun9eAGFqQ8BE76/LjmZcljTjqotYm59L9irXEMPHYUArOrxwTPOmotLEs
rNAAkpJ9Q9+KA5Pfr1imV88ecgCq1Pu5FSpmxWsQ53Otf5A2G67dObaNF+CZya/1
4Vjdp00pYV7JDSLZ20ayGrm3G85Gw1mnSEmlObGq53IKgoVtI9HlqAZvke8UfqtC
ElmQU2sktYQIrnlrhp2vsV/zwaSk87NA7Z6xvyx6BGIHQgSvqogtLBq9uCN0Y8Na
BLtkJsD2A3QmA86B96OkurXANCgcke+k1k4tfW5o+x4En7Be9+e9A83sxOuA0uO8
uyhqqA0ievLsDqUx8Ua9SGPuQxWOs0BXUDTlSVYcx6EJyDRSE/25VmIJkWxctib2
iPEEMoYnBaEQGOjCVg8duE2ZZRx7b397LnKRwtmq731F3aaPESlLZ/RqWlq0Fl6d
CUlh9P4SJ9cSmdaF3vkT0d6BLbOYnpnFBnRMIkqkA6qSx0XiYkJH/6bIuGxzLUMA
PuftaY0wMdIbFFstzDvK/mrVPxBJv5usdwy+WEY9fofk5oRGYunM+t9j7EVm714q
5h8bUpCoPF3Bf5csXXhqCGeNUIdFZ4zYMIVV+ddH8XkWzk7SVmASuDA1T/3oFdhk
vBb0ICpFlBuMVuW5EgRB0WAecYEO5Z6ijyYXFAdy2nfx+/yV3bTS4gtT3LHxWTzf
dbTU4IWUY9YMo/Wrlyje3mDl7tkFQPfQK0U9d9EjE77e+XSt1lL9kFgYxHAeaIw8
XYQzFvAz/qVUf+a9Se38oJ+J0g8UoQP4XcfntFfo92J/PAsdMIEk7zDDVSP+iu0a
BvpldEMwbtcWMz0HKcYUsnYB2Ubnj62P8dGCZTb2evIQf8uB+JCIXpL5Yw9uBzJF
4SfGvdNbCmmfxWgM/Cao9Bf7KD0caaIi87eH6hP0RkxhL8a+PCRK40c/3WNLckmE
ISd3OxqYzvPrjmIkrvVeC53Ts/f0w+pRialgKjdJZxQp3S0hFzpEG2yBjbmdV4aJ
L/VgZXYphtI43W+8wneCEJ5h3n76hAd+6vypuHBCZErEmXu4owQM6KIwR0Fw6n+p
GCs5MrBeondRTfpFXuYhcjJ1FLsUItVXQB4rrERmOUxHqP74vzkpPhhNJRjkh3a/
P20R9utCRht/HzHr43sOKzOkKT+drW7qkPWvGYw29Bbud6N2USUpduT0T+ebe0BD
1tIbiH2ru3PS/OVCOPY30nP5wEfQXAxEq+JphQOu4/A1fkSbMScEh+/+c68+xqeY
YuLKI3HmU+SGvjWeTXxF7PpmkXe9d5ko+MO567odYqSlLQGF5UVAmCwjOr/0TvbR
QQpueopjpk+5wQ3OMHyddr82UtOGTp5xiRmhnYk+KYj2CW/bTx9khoJXHZEsh6Ty
8J7VWpD04HjnFdpHgVzT7VafcNltxGKOHFGAMFkLRvcJ6CfYzLz8ignn6fMP1tH3
lXt54em/Yxz6wCH24lFNTmoTvrB4oRKjfJSG1wpw+zoNgIqpSIyVEIG7qv23Nf8r
nJUB0uFvejMu2LoI0zQgSpRWHMPpD8ef9KLH4tVVBotRA6sDsxKgo16stBkIyP8u
nrJNNz6dBpDZ8FqeAhTjZ4fkFeVw8KQPUvzL7Q9o+DUZARdoK/Aiwd+i47b+oP41
11/JCFzXOB4uyIW3+IvDitXS6X9iH52LuO2XwWXf0B1KcbnTQ6txTXXdgEmiFEYS
uUbbSJGZeDXvIwJ1f4ILyEsOWY+J0QY5AYgV4ri0HwpJjvxUN9KPbPflHEnnApOZ
P2S0S48BZwasSimF9V+nb+VGTAL5CwiuMC3e6mfEBqbUFs5HGSlvAYadJkWH34El
ft2w09yvs4YfeB6FTzHjB4VyHy+xb2iecuZUaCry72mSwz6/c7xZ35dgxEjwXX4W
dPRP+YjAH1e6RdgfvkU9Rg7H4YRp8Vf80vqnowqhSO8DmKxVF82cBpDdzcPz0GLu
snwJN7nOtYiEWMyxqIbiOGfhkA8UNei+jHngYFtuXCYA8azeo1vNLkOFsokgbT1V
tsWgzSQII8cD1bpvesEUhs6ktZ9I1FFjB2xS2LIElYZBWvBrD0FQtHwP03XQsRPy
i9hU9812bwC5ID45lSijgsYSgaCGkhU55HiF3xdEpV114lxoAalJqyeOK0H8EEa9
3lcFLzOV8TxlsQA5RkOYl4wGW1aNPGb1rmHAZqQEYUHnKH7MAv3BU6v8TZvUSI9x
RUbZ2Nlia1JyC6yw2hlbwmTpXOUfOCgjX0LGwc4tihiM+mUi1OKzPmoMRPFv/2Wc
3XBdrEgLyZgKtnjiDmVEnPxtpPOQF8Ovjwel3SA3rFbpJ7h/+zkWU76+PCZMhi7w
aW/phlRVP+d1NQefOTBHkhUOnuJXfLtPk+f5Udpr0e3q5GZ9sNGA4nTutz4BjWDO
H43rdq4VGsxNjtcXKohfRoQoNaYKL+5YdTtxmi9bSwvrkVS0wMEN3cm2zU5Y7Xo7
lHFwNZZMjWEzbGn3ISu0VXjoQfGTA+6N8laSPv/V6aa8AgXNYeHboDrZAy3U9GPl
t8qtoO1D4WQnjwZgWJRTrb0UrVq+NYd0zTSePDVtmDXYpayAL+uEgPTwTYPFQMv8
pxbRy1TetzD4hgtP9UN/Ye5Kzw2q9t1uldLFlnQZBufMszkxmVu5/q2srzzFQ/pR
VkSJeSOxaVXAAgKnEl0/Eg==
`protect end_protected