`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 21376 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhBNVMbsl6PTB5/ApNH6uD+D0J7Nd1ZGkjioM/q0trIs5
E/ZunsOVESFcQuX7N6g7zhp+QpEbTj8tAvEaMvDcdfe8WEDAt5sXLI4O0eXeih4p
tOFk9u6Qv7GqDWuMYMtXdoDBhYPIA7bUj1JKsJBlvoqCxwjpWKBFqKZ+NaN7bEwE
tQumPl8+12CRHA3JoOyxpz48K85sFzeQh8aOt5/3Mq0OSycFrfGTtYgPWuYHaFBU
G1qYL8gpxN8D/n/v7RCGhSFBlD7YLMl73ic7BylF0TLYk7Qr9GFf7znezLZEEb4b
PzuTjr5xnpQqc1/obfRZm+ewBJMvNCL9nqhefQYXcQtgHZNgWENDLzaeRF5lS1ka
mdgm1kqBHwSvb9IiL4W982Q8QNZf9qQ3h5yDaxPcDbsH5mfWCvgx+8WmrZR6OaQM
Hf1ZVzZLlbUZO7OI9dbtnZLZ30mlGnuYIg/p6PInSMYd//pWPcyHLcjBqdyDHnHD
ZqPIqxNGgRmAC0W1XhlEeE1Q1afv0AsI8nbMS+64PkPRI2lDmIqxUqncOmmQEsA0
HIkZnOzuNKRtg6wWf0jJ9/+4CCm/jQpMFYdwRbEC4oVfgYeyfsuHQuYhgoTOW7L5
J9RfquF/porkb8PzwxCwAK8aDO9F0+aPalnfjx+BjQqfLhOnjdQZBe7IAkbV1c+3
MSFi0Huzc/AmEWLFuF/0BCxERKlFeFWBhhS66s7bovWV9J/8ASGsTCmD3TZ7HtOO
fBczjbXN8t7bQEjJZQnhHSGpAcbCsajpnugHgwk381rlc/2ebwJ3HEia7uchvG9k
9MBxLB9TepG1m7S4tPbMdpEXJLNUH3HU5+dtfLJl2P8+QKihZFP9ssJbOrh++wUN
Wzwdw3mjzP4r62m7c/aPJlqlhXcomnbPHiHZDcZyeoTI6Xa1a0AK098CsAioye7G
5I6qeikWUkG6mGl2mTObkwyKSxVAT4sNDsxPA4e+UYjohipij4/zkWpnBr+5ODLF
QeVCHrydGd8ApJm9f19V8y+UT6Qq+IGtz5VtN4G9pv/rFo56F01BfBU9clWCK4o7
zXMn48osoCR+Ch8erghDNVmLmG0cgM+DqmiTwuc4ysFMOq8CIb9UhpBHC//7LpY6
R+kx0F/JSwW/7O77w/dZ4UCmZzWL/Xb1zH3b+Dccu05jIBZxiFtnyfVjJpDRorYC
o5dKGLMWXXSTEinbEIuEGFEqMHVHZv35oNig0r+DwNZUN+3RpP7ZVR5fn0JIzppL
wv2LJHdzl3AXriGnaVi+jqMU0Ds3kEEHLhG27QCHEpndkr3kOmtBiAkiuyr1/iZV
yU2bjnwBEIIil0XCvtnrcX9MaMwjsB3kVqHy1Cbe7ktnDOixGojzXuT7dL2y1fBV
plOSEmCl8b9/m35OPOmmFLks/i01OD+QuRHW1JbUp2WXgscThIGLagzU5ZgAKE6y
1zlM0l6rpCVZ8N9vFKZH4ANFsn3yfq01/TrwrCGwlKgC6AOsO730ReUT8JHUQVZd
iEMAwFBreruu7LYPARMtsfDJDt3rZymIjJlOJUVrN7ixuvO3NKuy1zDDO7wxoXsE
u05xz0VR4kCMBA4yb20UAOs6ahKLsgjV1EaU5v1qozIzUSvw5KH/Yzb/k63Sij9Q
Ki1pvfuMvQroMMr+ZjTRuFeLoDZH3RW8akmcIYTXsM0c3SRdP+tcRrXGI4GvBb8s
9YI2QKxGW5dObcios+iq60tirUvar55Ia4shvWofGWaa5RcA1HsMQpZ8vlaK5CmE
zh8MfvJhT6X4N6vOamvUZpfc+v8AEg3Q94I5IgYcz6FEMwebLMmIx+aepkfXTral
aKqWXzr8XqAfQohImUwdd+MD+VcqKZaqOjibxEXFAgnZc7DpjHbr+Z3iSBlrORsh
tjLk9MP0vmTfM0svhRZ1S8G7Zi8z49wSpVVHJFVHett0cEy2p6VgS/MmNoJFG6ye
g8RMmJzfWqKoV+xShSwJJPyanO367tfrwsRUbdpcG2h0Pkg/+3Cp5ClpOxp1wkT0
/hrier5bfL4TxV2688wTr+SRl/8KxcUjug0YUNejzEz8yEObGSckzw7EAIcQ42ih
S9Kx9l1XwCLk5jgKljWnTH/BdzrsuCOFRRmVYJRwnIo+DuVerAlZzc9Yl1bfZqCu
KBXGa/8du/mEIpQqjuJUBN/hkL4pUJ1M+IvnK0P/GbNOBf77vEcQfpgAnJAsKKoV
Rx36U0muzKvZVD1u80H0lA9M9uIes4TuZWC2WYcpj+IOMEQpKLuVe2YQwVSzpceR
bDaw65HSUH9KJjl3vlB8d4UL9dZdxDz28cLXhzpq7D8LwoQGoPHw1/SSR0/mgA+C
p1SjgXrSrxnkL6gYN8+lHKReIM8kCJkz+XkeChCZY2cCAEJb/j1NYCUC8zoDPN3p
xKD00NYhkoBGGKJm++kuzwVc7HJdWHZiz80mjIioOAqaLyY78aYXD9mTY2zbqnl+
RaufsDJcV/O/D7676kL337bwrigKW2nNxrvVxbGfbPdYfU2I6t21zsT/bUZP91tC
6ZYzDsQF3HCHoqWjhZ8as49RKVafFm3ffGKq2dE4ZgD631GINWCGKRLV6xEDDOqz
GCjUusuQOj9BfPJoGvBXBOzP9uWXw2wQietzwliKqmGb1wXVipx0uKONDgrIq1aE
GeYMD0Lo+2QoB1KYR0XuBt+oMD6ZRm1ltHlkWvYI1jyn9wP36d5JnO78LbEzn/E3
/RqJkDAwxld756WlLLbjD7Hx1nx5EpLvC2q3Vc/OSP2hZnkngPeJD2L75zZb9+9X
hbu/YWTx/S1Wtg0tWW+FhnVSWmMQOXPxKgN1dYu2iLquO2JgtTxgi845CLdKaR5O
47K1ysVjXBKlygmI0gFxiVqzR7OsqUFlN9Zy/QMtyMVyFRrc4ORkQZm38LsQPUR0
+q5WFmx0yKsdew85OL2LrHb367GewUiwCcXEGzHsWQZwQxbKIYjRbMBCVv5iJiUB
2fkEMsDfRbkI+QfDm1lkk02chkAjxrVlRQHXSjsORmv1pj6S4DX02nMAs8RID3qB
165NElQKW4AewedcoT2IU/tZaTMIdDffVso7DIcbjzGgYqp/vWqkB9Ztrr/Ok4ES
FePforZKngsWpAZCCUMQJMVxGPsAFsETKuRkP83llXYlcKBU26ysmwoYpc//4St6
CENgezczYE708tNTBHadpZ1lrjBqNCUp2hS7dqVwXbpRIjHew/i9TkzwnquBHnNU
+YAHZ9FnQjJMi0kIaMWHjw/oD+BJJHyB/UvjAqcoAQ0SyusARfozD6yukdnPIOaI
+omkyfk+t/WxVgQZhi6J/ahPhTI2drT2YhzYzQOYuJYb022eBUDlfl+0F4JQkwLO
A5hPKoGDb6OOIECoMqA5hoMe+hSjYuI+wGlInzWSBf+DPKnad3tENcmvYNQujll6
9sFQLkKA4SUTnNi7f7vs+u2aHUDNNNTyXkT2vJgDDgx7p+KFocUEQBiosK9ekR2d
jjOZyAjjkiVatLAuvRCu7VE+Szxvq2MklL7v6PUwRMT1+cKiSOampZ/Y2oHctO8y
fRSeIlbAUMAoljMg8rSxU9xM6/Xr0fbKBAGSQZ7lbBP8S2L9RheCFMhLw6jsJ4Y5
2lEJ92TzxJANrduFBOElVCmmPXIFFbNc4rN5n48UW4Qlz1DNbeT65Lq8bdTdnsVc
5Y1TInwU2OaVe8+vtLrUPr0AHdj2by0CvNosBrLXM9fam2Z/lRsUxyaOoJqkBSnR
Vv1qpgPfJmzdgBLmh1yOQy/kHOBYPa7y1QNRB155+n6lmUrhT9U+wpwtgAquYq4g
0FLYPuvHmCn2gE90L7oJXv2ySEIH//sZwUwMntZCw/8Mi1RjTpmDWIX808GwkWv2
A2IsBbqFFmqq0n33OALCBH3Ci/nzWBioC7ZAPyw5X7q+NI8UCwCFCI6Q8iNkRFTH
vS5gC4uf929GnJGaf2EaFKYt7P2/6gOh8zGxbsemzv9kGGMXq9nKlOuA+Z6oDY8H
Ih9CZ7M+hZQyGsm/YGuQAYg4xh0H1m6ggF2IUtERNbqKxvFrI2ndJhtyOZcAK21z
jBnNht4xXHwRuENPmp3sRgBWo3zB9lrIWvR0HcSrRCjJ/ufq5qnzcI1L9cdoIcia
eOpPQ5udp84yzyBvkMiADdLOOz79E+PS0PDKZ1t/AJsRURTi9S3lPFpHgpHVjsu7
F5ILitIkr2CxidtL+Lc4820KCMnXu5EdKSVN24tWCcwA765r+L5jRDLDICLBUX4J
MWYXPgkVGIJlKnh6ZJ18kxr/HcxKMBw6rctM+Czwdckc9sN/4loAk7ecj4BgE3ev
lXqIsYPU7rjF4kxWos1Qwngyc9ZOSAA0qMW74bitITj2u6U7EJUItNqJxwID/plM
49eXQCX5CoIJFU8bFjd0YdpC7/Xt/lGXPmAqfb8wdVNKO8OI1ew9tP6o222SAPex
Rp2CcRcLUyRBqGXe5wDIOG/BqhEVRdZkY6AsLXr8B4wpP1IKfooin39IX4W024GF
8Lk+aAZlTa5l09e8yuhmzdbuP6AB6tbnzmY6OZc2Ff8ZVc+z48PFQqWyrTXV3fNE
m6mu7iO8TDIQI7V2RHSDEcIj8Ybho/o6BRSk2lqID51tZ7/PCtEZLhMtbt+feWMi
wKWlMZi6WWqZI5eUpuiByW7lMun/y2m/RUe4jSkxNw3NtQ/LZclADS+z2RSHTJWJ
md6hjlmDtDA+U30KGjpKYj7VCIzbAsq2q+g+FgA8yVUxwfyoHi5RMvKb+0hf20Qs
U61Oldhj5kwFx/KJA/5cYyKZXV0i4xO8GtvMhGhgJjpKhhY4P4xFqOuuRyO5BJmB
FsN/2YLCjhWSUyGTtnH3F+lknzZxlGbCH5fQXbwo03bAlTjGzLGrWQuVzh/z+0Jx
AkBPeCecGVe6Scv/Qs9PSTnLDjS65rxd3NIxOawx8y79VKIykwYBwlCnAopFgXW7
UYI2/2idYE+1CG/Yax3Yu+aMf9u5azGRJJfMcV19ASlz7iZBXLTW7kOjxptWxcZB
NXo5HHEXrH/JNrclTsHfoaIJZaNfdTTENqDSwSA5dU2sg19oSYTmL6vyUPkdOx57
GXjATIxfwZ4i69MAAg+HQhBDkLJdXjaEpCaf+nxqBrBCwkoF/QRPNpS9G/kKnInE
JOaEnFGSg5cWYiUF912UaicjHMWeFdCcv9JdjNVpzeJEgzcmFo8DzfR2AjY7E4ab
dSfyYJ/M+lPYj/eHEU05jIrAZKeSAKGg2+xUKXr8a0cFa8iX1U8Ub5zrbU7XCP+w
Ags7r0RqtHTiH7180IMktC7jEnc1VsiDffyD7npoO2f6OYx++mwRT8oUhwr4BUYs
kIHzNTs1IFw7Gf+RcZSBcpHo0uvdIz9Cxp5wWzs713wF/YsGuQ7b4C+g5dXUVUej
jnXbyDByz1yywcy5xHZ12ur+xZEVYfHDz2l59+QBCBc0J1HHNULfVwDClIF39j5r
1/Ml/dC81GEjYtmpeNoDHHlW4arOgP0BBqaKY/UrbdreyrB5J9Yjh8VW7+pfTsQf
82jtYYWhHHWR93/GcUwHucRuuuHZi71XSGi7XOBoCP/wtYQusWeE7qZ94NvEBGSr
WcH881WlD74ROklXg0X8zrpGSHCtBwrRUMw9+Ar8NzICgFjb0xL+/MZKmZj1wQ9h
+/C9PfX5lcnWqs1PRzEM7s8FqoeYhUjAX4l0Gh1tsaqtQTUUwr7vz/WSqn+ejdaA
jrU5w8GV3zJaXcrJem33WoMABvRVOknauBh7VuL7wphI9UXxp7xhHb3dDMtBEMZU
BrGVIFrGyyMPTQo/vPVseyOzMfoVJaicGlYEa+lfQ5TpJAADXcOrEkALp7/UlspN
IgKbcFyIxN6JgvEL2SEGXXTCaPfmG3GXmP/ylw6pH1w4lVVNm7J9RDBq8eFXPrVD
yVNz+1zSaF9UE6SMN3gkl5PNRGquaAhJeJ97QO3CPrWq/nXpP+218w3yDGBmcEQs
izkmtsP0IJ+3JTq/H/mkDZXEWhfc40OH3PrGHyOgJXgW61BF+9RRsHxZn47RaARk
Q/rVLnj06Mo2TjOtt0ZTKgYPgjFFY8lFUtQn2ECYPIZ+QRZZITUZrDnySOyOMTOU
v4Q1LLdIo0KENr49IwFsIf0Ydrnk9ioYfCSXkAshnf/RPvEWReuxbDKTiryZZ8D8
yg+ZDV6OqfDOgUZOqL+BpRW6CvrHuCFUeF4L7MLGdHFptZ32Z4wpxHWWTfS9JeEC
+WFUH+zFSnJIrHiXRuXAf4gl3HrcHl1NiIaJzhAYGEp1qS1Ym9NM91JG8K3Qz2M8
w0Zq2S76v4V553ATjb8PCz/SCMtt5pvmvPu2g5jdgZocslnAl0P9qJ/BxSTck6br
VmZwuaUFGFi3dj9LcCH05zZJ3pjGC2vdr+0Aeb3ts4TqPGtgQaTCCGxVFrN17AEZ
F45J3g47Db8ug9KkfMvvxNkI4V7iDUNcXhFYTAcPdMTnKDjNjJDUjX4/g26gpWo4
EVeerv+aclGvJ+MnBewg6FnDYOr/I68rB/S71vYhm+wKobTPL84VfjFy8ixFh7Rx
yuWmonC7VgF8tNxjrxYdLkSlVH+xIckdrLlMV7AYpDdRe3e1eU0nR+6fk695PzM0
x8kcRvvIarx5zENUPY9o1af6hlTdXJ/jvKtL5VGzlC47rJ+tK36k9ipN2jg2/lEJ
0Ep0bEZ2yGX8v6SfWgldjKEirpP5ghpSwavuq4DRQHMGVDHKiy2MK9eUchH6XOOz
koNWFEOo1/hbriv5XIEtxLxfcx0MytHIhyauEqrGCpNh/NOhFIoTYSPpjCWyqj69
bLODagBNIndpUgdvGzuoqx1F6S48g4VePvnLYkdFTv9fso7hg9LURut5YbisPb4k
YWgh9Iue0dHhi3DjGYTcSiVkZjla/VXUce7zihyavtt0WK2qSvnRDT3tf+2Qq+rI
Wolr5IdLcQCioSYgYw/h1xV7BXZYr+1HKzNucXaHAoVcVRgR1CZl0v4K0znR3EEA
CnB7zv9rletgnkLRAVbrGjb7ofiCD3HnuDYZFzz4d9MDvcH9vd0/P94js3dMK8aA
nmp8CuQKHCj29LSGc861KZ8ancoSQkrxWA4qeQuloLq1Mn6oHcTXVpX78KL1VPCy
giD36Uyk2+1uOOxOgLQnELYqOIvT9z2zSSw9Wd3Y2vqFe4ttWsWPXqdufwtaWTE9
sGubcOV08wX9WGeq2bUWBNhQsu1HO6sE4iHR3Bbyj9+PQ4VdZ3Am6OfN9ZVC/YEG
NapOIV9VsB4QdhPSxYU8OwoAhNeBUiQ0Bmmm56Ud9IhvI2Fh+8yUVzwc3l/r0TPQ
5VX61PfWIAZ0yM+zgRL8/2I8PRHTNfhstlWXTdNTQpWmyfvNIqUfD4Q7qMhV6GUU
zeu2prShgVhQzjUo1IbKnPvug9pG8aIqoxBYpbl8AVv4Gy5cdP3dWrDXosIlvz4n
rqvy3rcJAXCu9uuB5kwqqtEC9JC20xWsgYbvEKhwaRsNW4LfuuPXFtEG3meveo78
6eCSMo/GOTUjNAwDUs5EJ6h1UfrqOLRbM9soX2FrIlT59IDPuRuy2pd+5j0Pr6/r
2STpVa9AQjRaDaIVZ/mKtOZJaqRCqa9wUHT4CrbeeRxr+k5UKQPUjssh7PHxDzWt
R/22wWMbcbR+IpgbEMhzfJGLX5C1HS/5JWuMFitW7B/gOGziGYZvPkNnsTCLfjVu
kOWmnylNxxE2iPycCf0objOwPD1ffP04Yr50PaMHFkgEUJxQnYoHTZFK836qcyYK
mutYc7nFlFgIsufzZda8arpXMOMKL6cEWKEgAbkWzITUwHuv9Rxf7NY54qYGeWm7
y39bYu1pYUC4bDVm8+aeG5npoRbFbBsJ/04bD/QaJkKdVJN5zjfhFb3fy7BQFof3
gWFdrpXI69SSoDbqEDaGN/g3qofyoTQoQsbT30QGv1sUaW8wCWbC05fxBqr1j3Lj
LhJgL55gUNTsrxb1kduHQcb5wHiPQvhrjkfFPMJXL07r6Fks/emU1n0fuQOHbmJM
9PUV88optwCYmww1QJMaoYdmnfQAc+1rII/Tzezk0O5JiYWMUlTYHsivS5LsQNIl
kyyCLMRjY5mhduHKOIcaEZoWQFNziA7BFPTjyvVYMfAtfWELqnwqYIxObbdIC7Kq
za+cH0HMArjhErk6rKkAMScKBIielR1mgN/lCN/MH1+urWW9rV1ms1rx7DqZOzKY
0aq9L1Br4MieF71DhiIJPQbtb3+CggONJAIvquyNqoFq3KbhJfO453G+gLuLqfMB
aPN2lSDuhk8uwxd8TeI0Tvuaat4+doluCd1GgH03vaMwX0aVpm9trthxFZ3c+v3a
Ac6A9aQQLa98ffWKdGiVH+82WVqU5u0gO+GPvIuLT/9fKC6spotFrtBC0sv2ilVm
Nc2OMbS4anp04TQuTJ+LRH3CquBqL4rNdhtg2an+WwJU604pWOFaHduQeHP2G4vO
ZLxQHm2ymKVa+VwzX/2FkzohlaR4u01RdS/NVV4tdUrJsQo97o6th+A2HNE4AMd2
ohOd/zd7ii3gmm4cA7FjNtDpum3HaVNzpmt0C/C3J7g5bfu8DehJw1Z/+mJWaSmN
gMGpuuUPchUTt5tTO512aniduT4zyZItI2/5zqCgScKpOwsvADRNYcYkEQ9gwYTX
SfynAfDA8ka/RMEAGNS38TRAK+g52OTtVcF8fuSbAtuBc21G30Eug/uOl+Xcwcpj
yWLsuY9Fqg3EHP24mP2LtdX32919ViLEkoLKS1gfNsOysIP53fZdCvsB42RrvuOQ
jN10Z12OIU9jPARj8jexb8x7UysDZbQSthi2mw//vg6Q3IZoiTrVO9IWJbBUx8NC
tezUNLxAAOTa/nXL9lqeG/zKJyUQb0XKxR2envIEEVSqNGvtr2H6eJPT9kLQvHK6
87wynRLvguXTkbVB9VOUVcdm4h1xc7eWJE39kYekAKY+JdgX87YDnppC9vYGxPGQ
eXYviUkYNoo0xSsMGtctjySGe0mbzmLwuLIsyFzm6kky+bzs+IC4agDiqrwI+pKr
m4hACXGFP7W4l8D3KAafnHi0QRX5KCbiTyF02xuWwxyEp91Y6cIC/zkBuWeIwXi3
rzp5lvGUsChjKygSOxIVH3RpLMvrDZWu5UsxfbyJnlTd7Y/s1zmQ3ZMotUkGbtKe
f/SDJbsGK9MAyv68GlhyAD0J0fI6EV335H+q14phmPpkp67FT8/PGHCGeyEpbO/0
Eaa6kRSEQ8FdUCtS3Tw2gOgDnTQ/eBtlqA3tyV3R7UfkxAOsRBcQn69G7VWJ3BDc
9SyqYKTTV30BhpKwSouB15CYX214yZOUVE2nFRxoOSTFxH6N0UQZ0rV3oMg0p8Gx
kbo0wjQOBtRqjr/RCCnG4vrWsexGPvFno7Bg+EdXTYJ996ZH20JdcSUnXfkL/gzx
hb2GvkCHq9yjeaUFrs5sLTcF6bFR8W5Ujw2aFZzS12qdOpQrsveW2kZKLXXwy8Io
d5vdKnHGK2WGm6zTZgBYIMARAtSAj/XknFRv0uzS/BGsMPdDPJA7KSRxckQ7BkET
ktemw9J9DkxoX1suh4lAyoT+Z+d/k34Ueq3xkPfMa8yGv8YdGQsoGDl+PDfk/onX
rwBfEgwzU+KpOeyNjpj/4+zw5aHyTigNX6SlWcSQEggb2kRTPomL673YyOCFLOxY
PLTF2c3jwJcJZaiNYBvXhYuILbZOZxLlJL903MDSpUhMiuvj/bOfcQUZAXLQVjhc
ffhhUlcsgSR3WOEcE+/ABdrGr3ZnPprFzmxzbN4DtHGtUwlQb037dMVhsLW/q/aj
co4T1bgeeACWXf+xC8ALj9h313Lm+mHkn87AzMRLjlkgbomzoWH7h2ONd+UPFOrg
wTCv3uGBpL92ZPvcPqscKYcUVnMBgQUfj6ApzvLLKLIJxvf5Mn6N0yNolOMGVIVc
3f3N99wQRbjTKahTsGrM1I1N0tP7tMVwqnlU+pu05rmdbknWPfgNtyGT+vnF3wC+
9U7/KiQv1hS+/8mwFuYPZKRMx2NBSqppeQLhuHm7Xy7P9+e+DiO/de6b2sGPQ8yS
Mw+8zNn5LK7TALatWdkLoeBAaofu+MrDWV0OoINfVkoDP7UG7d/czafq3v5l0kVg
Siq3xS3wlGcoJNHQ3Wp9d3iKvzQaSUUORTFWPgjROo3EvUZadS/fimTZjvgMHotg
cyJ3zAgdksZPt8essptTvpxTT5eikqVxuhv7izyNSKEaY24ygGLXpnpPLXe6GE28
qcOQ72kMqnpjtlv2flSi7TWvg6khtlS5arWVrVgvLO6aIACS4BGssGbNcJRDZ6xe
ZvgFJXUoOvo0X27pjHQdz456SP20Mc9ojfjTEt8UwylUItyKxl4dNX21wyDiQ4rU
Pg3nxQwCjzFXfvaQMzfty8q2EvlMk6rcFKXKqDlHosIl+omL6IS1/Pbx2tSOaLO/
1tuxkKR1x/sn72ROEjaGFruhDQzjm5NOYe9Rk2Y6Q/bpyQ2NEtSEQp4VEdhMcdWz
Orda4E7EsEYu38o2wGlXzGZUkF/6skFHt06MqNEjrlzguImNSB9KpwjPu9qjcKgc
hsTdDAwlbDf6La3UfwKl5ZkDynGVsskT/s61p0h74JU3pU4N6GNR4NosEEdV8BCb
VppiBwW32m+EHKDYwags9ZEILkcp7XZM/yvKwZPtVpt2cEEHrCM8iScXPy5qqdhL
gyAFsTWX7NLiFA+mT+zUrj/m/Zbd1YElHXQrKqIQBohuaBhOmF6sRDWRzYAY0sLq
T3hfwU127pqOO1O+aL7FZcSxYR7VhKaE0IFwCxJDog2kqSj9wJ5RU4QueytjXdJl
k0MoIe0amtDD0caPVRPIxDmk4VTYYyq9KrQVWoWdUp/qO9jORkMOfaGWpp+CNlTC
MZrfe8r/IaUDnmvEQXLFhHNC0kMVCL+frXx+qwHnEG2xfvv6CeSsFRZNX+KTknUm
eIdZ2cY8Wbi5lldEJ9ShVdO3Su5fDFBWoOpfGK0fJf4QbHJF063AsCm4OmUV/J5a
4Edgxp/+kVR+WFzoFwGW2AsNB7arnBrAwVMNWjBfvpzRYsym5ONJpDALrBc7Ih+S
T/e2lSBhlvc6/nl7gM2fITcnxJVxuI9hdnW+Q5RMj+LUfLBc30d+kT3pJjyjhmK5
sPxEuiVUYj8FuzcKpupDs7yAqLMuaJUfBrq613WO1O4RA59Qe+HVWyI3r8qkU/Um
twkZzCdIjNFCgwULcAjohFMqCmdQMzM37lhr7dAk3LQJVw94FBmcL4wYVhEizhre
boAvm2lDkyDC2SXrLvK56De7wZDJ9nAsEUyppKVnVvi80XerALQ+RERYAMt9l7LG
1mHutoIQuM37N5VAXTIx0x9dyE4x6E/31sYBVYIgnsx/65o7gisButcovUPBhouE
V7gNJMCVbieNFz5Gv8WUiI/HyfIraJVHEq8Ny9Y6PzVxfO51EW9EB3tafBG9guF5
HjHPJMArZmFF8z3dxv43/g6jhuA9JCgzTWSme3CptsOWNLZ2URvzjsQicG3vYaHt
ao/slDmO+CTlP5Hm7iXavxqzhimCNs0+UmmfEGtzavhAxVycbb2yx9pPu4L1WuEh
Ozf8x9ZgQzptI0Eq0N6Ugr7NOAk1CGgA6Aza7dfWdojBvo56wj8RrI4xCiWbe1/I
TqsPzdp+DZdHkBPTDGWcHn3kMWqYWZ5m5sh8fDIrml/YtwcfWEszfy54LpfUH7ZY
7CVwXaB9TzNqihVSxdVOOdHiUZBtr2PVeohgDYwZGNmyaJJ1LSlsuho1AxaXTVmL
uJQjwRc4YQ4kMjsriwBA72vvHA3yYgxUFqgwMgxhffKJVnpQGGktljWwISrihie7
jXL5CgIk3ed/YlQf03DRjU9MzsvCzK8XyiOWX6rjcvw5JTgMV9uzoRk4mZf7FSUW
8W09v2L12meRBjNq0y9jYigDfTZ/lg798rEsujkyJl6mgilyCd/JvIaczqF2BqLm
SvLhcrGlpcz5PVOLVbNKlr5SKq6/hpP+XDrxS38IqMKfsDiUgBggKa66GNqwh/UC
yhbVsJzA4/1KEugF11lC5W9VewV2avLUkJ/QaRbDmJa1/bKbqNNVThJneB36LJR7
M0pt7xMjPhyryyZw0litu2GquSSQKZs//iNUdS2OpsITJhUdJnMacJm6Vgc6HXMo
Fv+Q999uBTPZobASlboIH3SnwNLAgQXsZDIkPs80DRvryxCl34+UiyQmIkv+1PSz
XogrbIxQmzOH0h9xk9J6EIyXIJn4WXi7rBMfOw+btn6ng/K4z9eC43L96mP37Tis
d+iBMPK5++iAuQ0ohcIHFSuIBLZOoewuK/GdGWsHgHw5JzKgpGYKBiSqKpBRf2QN
I0L5hGVXFLiT7a/UtA7ySnBH28M08tf9XtRMRQRoNP0iRol84etS746XJZagv0Tm
aDBsYTBTzoCzXWXvjny1oPITUJvW52NdUcE2QhauAVaQsyfGeLLKrXLUZpTVCgRj
m4J9J1N8jZqayMUXo2DN4TJJIqQyVfdEGYpCWX9FJTxP2/tQ6EAMdLjGjMrXQj05
U+aWR9wsbDLRFfoGC3Oc0DmoUG5hafGoIPy9LSEgREmZds2bPGk79GTrhF4ZJMHC
4716D6/1w3BtMIh7iqGbFczAiQpo17bh8qT8AH9c4y5e/NhEk3WIzOmFKfK8KRGg
ZCRtG/69AE+y08kG8BCyGFihCQTGIDXOEmlFbCOG8oBD2fDUQiqFeFYToQ/4SDv2
IA3NmT4d27UAQ/u5aQdTAsZxuHyVl4nr8ZDpAn1v93X+lhZfRybFT4w6i9H+DCO0
idT4/mrEisXfGMY422qArcVUwufprvpJsp4LAXSAKGLUN7Di3kbeuPJITcVHGnhy
uKjq12yKiS83teh6qeig+mQDxJ1ZTmIzsR8tWNHfdQ8LtHW9wMibcUVHEL5oMAJn
SDnWgUgTdF0tCSdf7oHNk8tmmOpMm1IcLJOBzSUKVkquFHm4H5o9evGkoKlVoC66
/mOmdkh9HFf/3KYxSyFPAwKgYwETEpS4xyRMqWPoLHeC1QKY0CZTlVIuVFSBgJ2k
llBvCoog7lz7igdWxnfV0TmJyFKi4mDgPJhSJqE7kCT3UIc84p/2YtGM21EgjZEK
UgAKXeanIMRIHAdTlMrIawF7rjxavHctzvOKttEXrqVFekRivilLFyu3VubS8zvE
iEgVaftXPC/+O28mwwuOwxOPLsLYHnoKsC0NCIkXevX2XFkr8CQZvaKG20j0ErI4
oQSMMWW/Ne3iqdsaLgXOsZNK3I4TwXSSGikbvtdrZbwXbh0gS9q2sOLQLDHCFlQQ
uBmpzy23i4eBLGkzAwyeKNYBSUsNFV0BTcG9kROSYT252BWA7nMmXuMTL/mIaxmq
yEEbk5O0YRIAWHgG5H9pBoJ/E3nUaAzKlKItxvMgywJR3dmq35PB/hru6JHSHkRW
fIaK3LTn283fpxwW96Hu3usLYt+ROyZTo/Vra8khK0wIGzSSR6s2VBOR/1qfA0gO
rMnlR6ZgoXsmaSCQzQUXpzYcpStYLOYOUBQs078YLrEZzkp6qdZNba0sMHwsDRQQ
9NfxXMBTnAaIi/zbXDkDLrjiJGtPXkFz1hbpScCAw2M2BXiVZ5bAxV2mpbcMzfx4
B8fxLOSyeYTPLUdB0Q/3xDQJIuqkGUO/8FTJRRCvCPhVb0Dbym27ht9XSMrXBe99
7k/FEyyN4hi60k21WrtVV+3d9+b5htMtBqqXuvf5LCMkkhu8s9euzSUcMcxGkI/7
gTwsqs5zHYmLLBXriFviqKwxw2ezoU2HIUov3Hb9DF1snM61qyVpeKAJqcx9ZiwK
15wtwsV2r2brzpLAqI/xcDCkOkpFZKAifA3M7dtVZux6rn7iACb3UDhauGmqJR36
wNRf7aWLXWBfWn/ra7mSvBKhHLEa5IFxfLINOjikK6CnNzOX9nE09GjpOwVbUKiN
n9mqGxKd6VhpK9kO05vplcriJ+eJhu+eoC4alANPk0jQwKKCQ9XwBWJcMtSHpOhs
dcRF3l4cY4tLPW0yo1v52BRlK1biKtngYMkOY28rGK26+dBoJNr3yosy7WZXXlwL
k4AxiP1nj6n3mK7e8Nltd0gyV0HpLUaHzrXSncP3N8bL45jyXfSfsUgd+lDykjS2
B5LEWAElegPDtSIuawQ/gHhILtE9Sibd+1Ex5liweCD6oi0dAFr/w0MNWT8EVg40
7qov1M6bMaRJZEoKubq76caGWf0negLyTgsmxka4en50R9CnLA41aCQy3VWj1848
8i1nRJqwaA/IUVh0g1d0NrXyjDu6iAVQ5pwEh9J1D/vzOOKW+Z7qpAlsEgf7qLii
T2wnass6jGP6PsYsZlymKRwiabd69hF+V0gj3SBmsOmBxc7EcljMCEP2BHJkqKC/
vztGsNPpcrwaZqN9QZ5hUrHCcwbrYHkshQN3efoq7ppjj48KBrg6wYMyOeFW45EK
ShOwvhaIdQt1pmSL3kXm/uMosoYBi7KEve5GrNGDFm7isoz1t8wHVpfGqZtdPpkf
WhNQEcKtsv8w1tIF6vKm6Yi6QjYMzEwyh4YZR8DZYgm+BTY4OQIyyLOphPeWoTZL
dqaUI+vbHneGSu4P5ifagbZGCEo25MN+NKrT0KxBLEWO6GSo1KNSkiXytXAIdEY/
a3GoplzwggByfjcRWzABzuoeMVHoMrkQcsVMaFnGmI8kmLE5vlPJKWqw0AFAHSQk
E4Qw8zpcYsEeH0sREoQuq7QbILsYadd//TZm1DtN7/9YCgr3e90WXu6Pk8knc+Q0
VNMRVt5oghlzUym+bMGCnP/vtALUIBTV2OCTpDNMxHHTbG4Nr83mnaspzEtNYWT9
pxqw0qQhhniWLs4/cCMLOqOe8DbYZksk1hZNqqgEfA4SOo54KQ7yNXJW7pbco+7u
692KgN8/clWbdv60hb69w7EkjA5FyMKCOovBz04gJB3Ad7R4fXZTNmu36r860z5+
NkPDk9epEUp2IYO2xfPXsmSo5PlLqVi38JrZh5FnXV/yrhisX6Avgr7GKmw+WKVr
0acPET7l/IUOgsDvCaORuH6Adt0wOlgwbVbdlLrW6pbUVU6TVVx1aT22VOPes7Bw
Xfqs8liDUVpQqTfCXqp/iTlR2KqoGqOA/pSDciZBToLTBkoLj7Zpfm8UkGoycAvp
hXoFypYMAt71C1m54diQhAPI0dW0X7EcKz3gUBOuSU646Pkex0+kf6RK35SRp90o
1Nlgb18XJk17i5LHtZXVXtbyBU860UJuxulCSxRADFvwvsBs+VxPcjXcrF+6T0d+
D3fhH7Uyu2x7JvW1wNFoYS/VmeQmOOB8+L7jjGuOo1jgnga8+lRKig6MnyaaKUT0
OXP4hFwlyA0ProY4bw1RIIxJ9X/jtqoBg4JPChfrvAAhDOF+fzvYHIjNwGINxAQa
sdFFUPN/83iXX6QjMGyd2Y/Z/TvZIdfNSo+CKBEvR6EY5fTO9xXqbUqFHeotqxan
03wN8TXJUP8760DjsASbvCOuez4B4+KWb7MWzAk0diyWfgyZn9J/MHus1sv2nuxV
Zl/rAmWNrgMfXexhCZ9Xcbrnc8d27abHZZDydCiJWKuohtkPSRFCdc4ivMa0meMv
CsRE3W/FnfuL07yxUrwtlHP7cZ+uxYKqzMZPToYXIKSVq/FhiCFVRveWE9/7oLJH
q2uJQpAv1bxfftZRSEFr3+JQEkM4UismWMAHXVJ9JXPvXpS1VvnS6r5o16u+bR1D
ZmX5MC2pY8BU5+nql47sX7IrJdF6otG1clIJIeWuA2bqNpSs1lJFHTCq8vw3d7+o
j4NuhIlSk9CrgZ9pi6h9pX43Ph9cFpJcV9XLr1ol5sdescZ47aKpsDw+lpWYQeuZ
jlNjdjsyAxtXUjpjcpK78yfnSsa78kRc8qmWHGuWJPf6npF3ppb6dJtsWUn6AmY2
H2z0aQMUy/gNf1hAtXsWZ2QW31XxGIWWsC4zYV1wKEY70JGjqS07GIdRoP2Hcnaz
vJiy913E5lKaTIRXDYiWB9ZTh8Oje6feIcCSVfi/ixCLMIDCT/41jPz+DDHbpftJ
r7P6mun0esIdJ8nM4xIaGBCqnRjCQl0heR+EAC0Dh9LA0zqOav69uA5PeHqTippJ
M/8dUaeQcEL0U3+kWemZzMXNQWxc1qbmtsb6Cp9U9v1InlkXTfaNMJx2MGJ/sNFu
f3tKgcd3CqWjorSIxO1GP85RHbsPqYJg9ALN/dCtIXsxgwEVuRljDeOsGx+MHvQK
AtsxxR+RGn6wkUfBsN/9P9TCRG6q+kgfW0mhs1eELpzQtHy+PiNq+P5lOTL6ITix
PT9ccMIISOIgJDP3KtCYuprBzShGJ/FmnaS03LsRd+J74LqaXbGgBy8KKCNFdPjI
rz0ICQJD3crzfDzA0wbPsSzhnQeSH4zcrYMyq8/2gWBMsyy6ITBSj9wYkxbqRcQl
CrahTj0/zql+R5z8tVMmwvY7cNC7QNAyCoRKzVz+V5znmOQHuYJz855hn17i4NHO
h2mfJmbC+pSKdqOD/yEtVNPSh8y5ddgAdafUAFSA8SkY1hC9jeqbeIp/JfgO/NPr
SAcPxKiDIEYatpfnHIt/NRzK2UKw30252fyYitPb92hR3Ss8WmoSdZw5rDeZs/PI
4YwpP2oQrtyaocoEUN6HfGEIie1AqSGBAst32WBYIB+HBdrAcVCR5yuAD7v06G6K
Ct+7k24+YlFKZSdj+yuxXYmi00GVDJ6EoCntV6kOdrRXvuioBSDTiEDJ1uDmWhQ/
juCYH6Pw14ClXbb+z59sGB01hDbF+WVOMYjoxboi8zCcar1XPf8bYIyGtsy3FJlU
udsZVikFM95PuU+FTYNezadon8N/hv8ExPgPKOpYlptSUaqxcD5dHzhol+siqDMi
GermIlM7rCS6W14TspMUIf8JAlEGbIYJ7aop3fwXoKzVATb7icKgBlH1ARRkB5MQ
d8pm/BCADoZonfKNRvyJmzaWTkOkK2iylbqKrOY0EeLeh3FZX9uia1NxgsCBXwY6
ty0bLpHJXbLKufH8QQbU6lVcUlwFdw4t5o4qbQh7Zuv7aHAJtGqQpuZOI6df/jLG
bELDq+r+fvB7I2epOGnZcdFbyZLlWsCslTmduvTQ1cEHMFKD0HWsbjd5eO+E192v
q6Y6APkCcN4XayZvxoN7wGHuc8VsCJExLIbXxgzOkt8ytOeKYJi8zDRP4htJfRct
qJi1hektL9UWvy9xl0BkgVjqdsSsUn2N+dNOcWYW0Ql90NlEE5hFJ5W96AdjX9Ij
v7GQpIaVN9EnNglln0K3yUnie/j736lldDbPLdtyMf5VBvtIlUQTP0Z1dmnQqn4d
292AQXknwbz+Q6m/jQxFPmB9bvv+YhdA2DtkAiDeDmG10tDeVTgBtMmb2ktRwP6h
1+YCM56jPlRbX6p5VWIt244ZALtRq1ORa3/u563IXTVsgQm4KElmSDMK8/twjDyZ
SQMBsgJuBHC1Fonn/B2xOs4Ynk3lF/QeMZB0OTsm3rCHN/e8c0VKZs66CukOGxeg
q9ziXnjKrDO23gUZccdVnQbJYy1jrwgvU+yHVDDOUEEaZf5TUiHKmMjZvazeUjpf
9LWm716d0uATA2OGxjJEFZI01YFL/r2U6wtpOyX1haksZ9Jm32DtwLUUesXS6Qfv
5+cU8OpfFZoNCOY227P/Lhp7rzrsLIpF5rVpCmyzQP+Ra91Li0KqYzFybg6DqKNM
xMUmnKvgkFHvqpe8/MqQZxect80YKAQx2BERfILw+TNg4Cb9KSYO333YIoxXM70H
ld6x3pSAFzPBmppj5QWxR5fVHBdQ2Ykm7UH5WaKUrDuVAnNuvXN3XekFfjkm8N4V
hWYOGg0TwVE4XgiYOlTbSzSSSdUSyE5Zl4nUveSSVtR2clhPtK6MiOstlZe4ADN7
m/+/P4uZTIXY8ZukfQ3QR0FQnygtf0/axJHZcyH1R33a8EnuvU4MotgYiOswfwr1
LjWGuIU0VXGtkNOI06Kw7XLdVUWPqntfTlkO34NsXBzVloDBtc7TRfuCc/rwBdcz
roSq5RNpF8vH1PbAKQ5ZjUUnPuNQetIUFfR7xZncWwRJz1yyL7Ri2NdaOoxpTPmI
icf65WHqGFEaokFLzRQQcUl5hFWFjXVO85khaLXp4lwyyEuMOJIL4a0vNdb9Et20
MR+MWn51pYk5XTG7CLr9mZybRFLYvPc5cy/lzR2iGolpTMtAVGn/lUK1b1dr8SSg
ea8zBJ+USqWYMcB9njrxSUlBk98YPiAfLCPNLnfyeWji+PI0WKKb769xTv5YQsxP
s4lU4xZhwtiDu//J+A/r4e3HKvRkWVfOycwAFwm+cur+uK0A1ocE94ceEejqZ5is
vejEnOg10Yl/flgt4J3seAG9AbMA4ydr/u1dMiFC7hjrZpE2Z/HgoVFwaY9av86c
Dxnbxi1pWZ5cIKPklITRcQegBUgfJQ1OQWHxHMXlndN2izauzyJ1rNaXOsriRx2P
h8nXbxopWupGp5Q3WuFtdUxt3Ag6JOs5OQ5yj+KcnZfnNNtKy2RLq79+i1x6k6fg
8rvzY7RhOCBcgvhXjIrhldp2/PnO7Vz+MmGZq3T860TWM+1BXhzzINVdCvQZC0va
WNMDZiKO/z7chemXvKS3BF0SUEGl64XRxzsm/p+NXMyDUh/dmqSloGuah0mVnTwA
afhAx05cj90YChHGuWUSYNMkqVwB7WE4JBfjEuU4Ugmo822VyYRe0DXazoSVfiF5
93GRs9/3TSHRJDIAHytirZ6yVgE6/Iv2iWLUobPTXQoNPu0B4+gkCDOaiXm3EwdF
nzHOMllx7+g6y40N4w10yoU0jMr2n/lJQEn1U/+TZqmrDOIx/Rr9+NjoUwQGARts
O5ZTUQro7e7x946kDlK8X2u4PoeTR2DtZC8SIXhHBQEwZi+bV2p5HX1x5Ihch33s
OFOeB/rNlTNnSa4hmFgOTjlP2P1xACsHSsc8gBmRVR1fwYRy5iRDE+HLcNpVJVGS
iLUUT5/C9Njvb+L4/Iyl4AkajGMLlWBm7Wf1iO6qVJnoCFMOgzfKdpOZa6roq7QY
7n35C1svyiqCQ8GC55j4UWrti+c9OJuOkElqy77iJ36iyv+nwjSkXwmxionnsl7+
KZhXeDldyOP/zsR2NeK35e+HIEQ+lVspJDrIYod4Er+oMK9XQY4USXhDe74rQ3WN
Vlmb8dR7U4+bHr3h7qs3l5xoVLPE9MdA0P31SYiduPhcYQXcBF26HHrzd3VWmGtY
dHxLjFyctwJ+GGfs35S/9zwAXHS752f1HbZWI+ThfHsozMrKqMI+YZo8g711lVjC
20Nyb66qLuelo3DEKqowD4AeaEwAeySeah7wmb2r6aTBYRIl7lalCvLRCQ57OuLh
nIVLigO3j9HcLxt0DlHy0RuSOPM0cQBic71H8BpgwAqneCVjxj9BEpvcM4hgH0Fd
8+yzSlS0YoOeQmlkc0gLu7WykgB6EkHaa7PahI+ngTmG84zgqES/6Aqkpas/bQEI
cIdc4BT9KDzswK/Dhg8G2oHX0mC1dSis2TLG9fzhTIgdJRPAR6xtzIqFFbLTtxYt
f0/Jyy7qC3BCWiic4URWyUOS8/mXGbrREBAC3FE82JJVJZezPKPa9GrGE0NSVp7+
c+LA0IqVrlfr5FPQLKcmtjcZ51+0UNgjouRsAnDBRWBmLd3z5p7Vg3yphaWR/YQn
NZ128T1HoExrHRojlWWbLUm405AE6RcxDtYkSsc9tCsndzBEYm6x/mi0JEnnGisd
dje1Ov42kBnZQDfdWehr4vR7vMCj9RdpejW3/OX8lAZruwxdu6pJC1l8Cg0uCoiO
w+HP3zA2hKcpHvJxzKX346Kg4lYJLjXwwUUQgBjqvSiUNqgS8cOvM40mloP52Ua0
sZg47E5sWmDryWWdjsl5rg4jLVrjwZkLLVWfEX5CKDb5f9+Z4DmkETOluHI7l0h0
K/jdmBujAHyzBBfH3u8i9AIKLwiDx0vIgtmrKywG0zMkYKeY2AlJyX4a4vFvJ+Gb
1gg58tzSATC3rQhDpSBmUO/9grRKpO1Gy12FlQYWuCUVE+pID6h4rzX6EJgx90xt
u7cfv8xUnf2x+v6J2H50rDicofZWg3emiWNEkvO9tX5R85+M5P//Nluc8b/TA+g9
anUM8WJt9YjWK17KpZTtwD6hHyFbfgRjl6l6H6wetzcySuhauDHmrE4MaL+IEpN+
o1DRO7LWLGWqKHdPutl4c3iyZPC5DHM/jeOI5yX5r7JWdrk7dHib4Jho2dXX+crP
xbt1QUd438hAovKfW5uOaiCA8dvT5HJYFfE7Mzd5WcZkQQCQeb5X4HwpGprlFji+
eCygHJKUTBBu4ntPno1w9UtrpSK3mKG1M6jNg31afup0S8jgKKKH9raemf/kLv1z
ing4YfXg7hwC3Y82TTRg+oEE4O48luJH2gzbmodbKju16dDOh7JoKENI/Bf19Y0d
Sn97ig5Femr4xdx9VqxVzD8eEGaYvHdUauI70cZzzwmtB/+/97IieK+NNPthEeqX
nNTuiK4YU0JTBj5NhYFrE8PGvxpmmTQHQb5q8/XR0bD8sVp2AZDCw5j+VR+PK35L
BFnArlDU+LxqOitWhTQHeJLiSOS0EW2IzGmgRJxKj9LiYrhB+e6Zek+84nhBZti3
Bst7gq7CBUCEs+0wRt1GpAvTbA3Lxw9Crp17efuNyOyeewR5mcu8x3IrtrSjubyF
ldy+pr/yfvkOfffevMmS6/w7lvWZcG3wKYZ9tpkoXU+42X1/URzz0mQsRLoH9TO3
t9UxedYeB0UEqJpWj6cCto6AnO54zjyvrbBz/LcbMpS8IEIQG8CXkw22LcI4Niyx
/JP+UiPdyui1q8I3BFM8oGEYa80wb9jcS+bepcsFLwNb7uezGfZYe/9KLA9hlz7m
ysNI9TVuhLJVBSJP9gsOrB3HYByJYESyBo2HyTwjMHCkxHBW5toYAiUkcbvbgevC
qVUbPq8gaxR7xnXcPUspDwfehBufmJImrHMm7xRB5DU2qgfulCJH0f8NwP40iya4
f5KHlaYhvMQRVEVsDmW+L4MY/4q9LHb8Jmns7fx79GfEBQ16V7+2sIsCVadzSVVc
tQMuhlUqcOmzKltmD9dw9ZTCpHTDcnGoBXONLREZIHl4wbcoCK3OVctl88u1mec+
IhVMADJ85Io3cEh7Z8nPOTxOKmZYem1idgPGTLHo8S+1fT3iWTvlBsF7Om83S4rL
pA+Ajl4Chyhry/8+aNRpyN6jiW3FOfoBPVliZvwVfQ7vVkkpL44OxyjZk11fV/5w
+KxW2XE8AW433QWAQKWUpOYCvgAml2eWEv70Zle03HlWC3+eL66tu2604y5l8ZIv
AObmMpHW2uzoRx/Si0g6Tw1Q7cVrLqUdx9MQ/9vQ/DVwpXje+5RflTMJdpRC3PNX
8Ax/5W0umTWi5D8V9cC4ARlmYHzpZtn+i3JbwvB/Nwdz6aCf19arSNYmOFAPqrMW
Hx7J7KPbZCfagF7hNw3P8BAAU8JbeGzwXHGGcbRSP+s4R2jzYN25ZV9St76lWqsL
W5a/YeC+FWlO6cI7aK2iInWR02UbWLo6S5TiYJWV567Ictr6nGeZtGoUgilL7xkN
3EyLrbR5y7T04l6NjCyQ4BS6OmLy5Kg3MtAf1pol4cq8dIMBeu/rg137Gzul8eEQ
v4UC/HIec6HzkfBsKSG8pFCbOuwn+OToEi7l3mzOqcz/PGnE4B9V+1Jf9uq2l+PI
2QxlUh4ZMtatQ0dpuCSGW8a6AiWEvlUCViUXyVININvSSGn2J9VQC5tdz1e8R1i+
MEsjz7mGNZvnPpqyUN6qPGKheI6Wi438FRqB+dqFzX3/SC7SiaJfLmY97vEIXXzl
+KjXbxA5iWGOtaFoSd5rJBUG/cu+39QETIk1k19y5nmMO0eDPar48wu1CcMHIvCM
eY5a1soskLRTkzljpTPy8fAjR4/+3/a9aDWnMb06J03ePS+8uU80gK6ceCrrjAHB
S+F/tFSsgowtFosvQuADuWBsx1A24TADemw+v6GGfObfmnjeO0LbmJ5boSC+tWpy
CCqEigi6SAla9E1A5/WaOrWZBNBcKemPkhFhKnun98eMdJQMSt0bT+cvSjb6v/bj
qa7bkM+vy2Y9+Q/7oWH4Un80LG/c7/PUDOIX5b9pAGuawHZYEgmqDDmRzCBvlvfA
8zsqnY0o3x3q1KTyTFnJ4k2gux+wrYa8MPA3q48tsjs8Cy7gI+dadxtd9YpMAbi1
EBfleAu1ZztlA1jIqsWlt15Jjnb9Q9gL+l4DPl/3erMwOHXcP8STNlak3qTSkjEv
sXMOJB9FSJYnaAf3vsNwm5hWp8UoE53pmff5XtIn4htrY4h3SrJC5JCEmEmuNCyq
d2NnpQAWWpOrJWEDkSU3/BOqNeXsFpAOr+CeM1gHoXtAJ/+fk4lRo5l2VSnIkrjE
DPw3BQk4gJa9FvLbR/31WqUTZVmIwSyy7j4yFwb0KM5+gNCsL+SU+62L2fsnqc4d
SW8KAjwWksCccCb7AcXfbbf6Cz0dLQpu8dBLvhBh2uJaUEfjHgIrtJm/KBndpLlW
CV5ZKOEIPTbUmAMJLNLhJN/FTQc+/SPjDiusEMPf9YSt44UJ3adT0Z56hbEAhS/5
ol+hnDOtnQ0Sjo2946qG3YfdM92JG03KFc+pDoM/kVc0f2ccbHYnl1j8/geCnUjy
pZChoBBQUhiYizaX82dTqcOQgV+cjNVJOGfsIdwJc8u5HVePWe7gev2sGzE3imky
WBJDPnDkOLOWnlFkcYaJGtYVMDvmTxEpgC/wd1ZBg7gbz9n+EmCabuvHd6+seN9H
adHfXym/zD737TDvxQpgzRwYelUsja0ECV0U/Ar8cqUsEsYCXFBYixiEqnwiHNaG
xwanpsJMUgs53Vhx6xlxYGgDamVyH/zMBxiesS9EUFfWevqOwzvho/Pmjrc6Cymj
eCQidGdpVpY//jSvA6P+mT3h0knWIoNmtOFfHesXDEd+40VJAKQ2aEWUAx+54wEx
+0psloS+KibeOf2lyCRkI92hJPKBLUH/mrDuhpylK/dG82eXHSP7de7cYOMznMu7
RuSL/Qyn70dmTTHIRhtjz0G5q5CxAqMjHfEsMNSuv1s42sWnjbLLVp+kpMEmH6Hm
PPKHorDH6o5lJbJXOaN0bmMqX8b3mfKnWSEh8jz55Z+vwfwY0Ntq6Xjha4KdFRTT
oMJlLn4SlecYpnxu4m9Lw/tIUIqLhza2pa9zW2mxQ5RKgiJeorc/ZZ8obLqWgnjf
TfDdzjsU7Phyl0rkxwNP0zCPMC3QSJ8l65B07LYOT9+pNZ0zVtswMbyiz8ILMV52
+WhI5C6pRSMXiDjFsRABwOo0gLtUV/BOyDyRVQVRmiG0rO1Vesw4siI1Cek5jvKd
Xh/31uj0KxEviwaGEVufd6PZVlPuhP3FM8nn7lER4w6nKEOS2yF98jQIlDKmNWjv
5iWy+V9n/pPxyTKjQIFEIjxGRy/WUxZYYtoK1B7g4z0mQIZzDjH8N12L27EEiKSI
iU8k16uvdhRJwuhTOJonK9ndf1kSeWe7LasWLiKotLCkYZYe3EbvhPX71W/Qq+9p
VPjX5295sqtTIuARoVg0IuQNNhq/6cW+4A6I9/NNioVrIz/K61gAgTEPKZeY0mU9
nkQMCFurRAoy1CxVDevxwFukdGncb1Hts2b+O6z4nUu+X/gYzxzM9Bz0o6TL8ZXl
kOal9M4Exj33gRs8TOEE/rdsDG4Y8MUiGp3ni8pXyBMqOds5VsuChfxvaG8BCbZm
mlSKz7oIj8Re4/uNOI1ssnM5hYv2qqk1jYWbU1mLy0HjEzY6EzP3SEjOhWL92S+Q
EKCrrFI6f2JxL3Z+G/WzkZhIP50YIVsEhO401VCMKzPxZN9yUGVyhhVUU3YlZsIm
ltAP05X3QoID/74QSEvA/K1jKsv/xuIwN5TEu7ULBPcbM/JPlnlehCiiSrU5fYrp
BRsuHvAlsqzE7jRAbZBkaQcdsmmZUF21/gvU/p+KuLwAkzHRYdrDAo9FtIiVFw0w
/7Y7WKwmttxplca4ifxHU7iXFwOY/CH+N4YZL5TzLk6RycMiqxPyfg7Cz8E3Ka9T
m9IM2hq/H9FLscfbO9xhiwVtOXgRQMdoT7OS2fuo/vYlcIFnTwfmQA0CXKbwauzy
oViJ9Sr3puauDG2jBBXy/dOdsgAKtKCUyCbIK2wtHjMZR6E5lGGZNxJms+6ov2LL
QUwn4nqOrDyW0XJTboWBeUydNHvnRlweOa2Her/FeigCIkdweJOlTVy3FOeGIpvF
2qjMIx3nxACb/PiCpIU9NUXRek91NGo2V5v375CvvdMtsPMN6/uzrkuWkgrBlNQc
8r7EojAINNff683pnWXgOLhKGd+tg7SydP+Zxs/AQj4oHY5Xd5o/+wyxidtCpx0s
X2sQxBoaUWeK/TM2le3pEPmCe95mh1ivqBMrsgW3qml28VUVIPBG0UOD0zfRPp03
Br5NSvag62FH63SunjUs0tFHOtjqB4BMdMKWHKzeu+8aBiKlwL4fQDlBngoBnWnl
v+RpChNQ740fh5+nZshcFWlAZnj3cHXpnF8wwTS7G8LPKTuNzQiwgHiExnoVSBV6
GaZoFo1tSDaYXlaZ3b9vL/ySjl2xiztfqBkCQvkg23ycE9eUcgExx+OH8D4yZeF7
zo8JO4ZYZg2hbG0COgK0GjTQBIvJuICCFLQW/mPnwQQUfjM5s5SClTljfM/A9Ft2
X9TCnSJfj9rb+1txftE2cUid9fnNVE/IFsvE29KSFPmbF9rfe3uiLMS3w0f92p5v
nI3vJfNO1zC6/1vNHjVRu/fYvYuUepOmCBiRU66Zyh+zLNZOKYovoGAdWYqeR5wW
Pjm7PIhudF6foggUdgTtT0ZA2ElocuEwiuwdEbuzDvaUAhtwxpcqgeJyIYxiKyIj
pnUZgJHuQ9pG9POEi62Nt7mexEHMON2YHoHQTRqRXZLIeQ1gpy5AejF+N0oT7pDr
H1N9m0B+NsBmAsJ7pGe43jY9E0S7OensY07ND189cxiTLjWBI/73/qHqDnTcoqDJ
k2s/i6ysQGwPhwxeaE5PxXEGy9RHC9md3/O6N8E4qonTlyEqMGmTvr6Q3KBwZtTP
0dY4MGsFO5a62CsmD8Aq8sH2uj4NvhYGW8gAQ+2VJ+VKsoI2GZNYbgUTJZ5odCqF
VYqbIkqq2UnMqBw28Uz/yKF6sAxQrUbG7OGemmwNLjUz10rfomNOIFjbVXiLlcFM
rfuEslIHjylqP0HtvbrrT9fe4ekNqQMug0d9s0MaO8gi0umFJD8npgL5hN8dNP9A
bsvRfUbTKofqfdm6zgbKRtJQVZXOAQeoGXTJgGXjUIAq0TnpJPG2D65SCzrEgEPR
LrS/KAhmZxrmlIwiht2IH34tJimOkbJSzaSv9DXfmod8Xgpo0WiZPr+LpjHo8KM/
qNtFilsW9WBfeyH7bwjTC66oR1278y+LUQqkfNmwGRQAfrUc/uVn2jRkYlpibkAw
ae7UFaRpMWL/+/NiOR7t1v7ZVFO3bjo3bjYgxTtaQH86XAPf1bm9F84fwj3Px77S
t9FxDvEOpN+tAou7KVaASaZvCakz5A5blofLxMFUwAzaX2WQaXg/nW9pCpS3hJap
LILgmfnjwNh1JbIGA5lfvWAsEHclRLp9mBfGCCP1bKI+NpoSEEuxlFlAxxypTSFa
L//ey9K0LGAjPVyQClytkAO4urW/v7xfZh/t17Wv/UQ7Ff3arOAwa3/nXdDFuy1u
FqDzaZA9Vr4IijyhyLs6BMK/zvb3kAwTsXikJIc3g/8yQjdH+/bX6X6UpATcILOA
UwTqBKF3R5NfNPN5zR5+siaXDPL2ekhMZaNI3LHsAjau4JFMlkUz4jBEUe6Ds2m8
KpDv/ibY2wqHTj9/JGCrVLOLbQkqbs1DsILDUlIjJcCKE6aApzz31A+vKD+lPnfp
b3QecN9u8jEvFExGqTkDy9fe9oWmOFOMgmmbin4ocdVizMVoUd6LAcI4uC7GtHdW
m66tT0hOHLm9p6EQWIEZuXBPtKxLnnhWVxMrErmxieGrY0cUi6oTpe3zY8ycTLrt
8Fx3BSBsLJqCKNC08I2mPapA12awsvC7QTqsztqIJ+jBlWtYlXjICDuPnTjj7Ysx
Mq5P0x5NXEs7X/cYukYdReKXqljnDhOmfPeS2wUMfcB/OuDf51NbMmpGwXuEWRF7
4FeAzIIjthLXyAm1PWIAhYcQOfvXcXOmJmgzc8kjvVo2eUeQ1DgYbLN5yIlsxiQv
pez9dmvgu71GZcJ//eQtyAj7lSUR8+ttnRf1D0axrarpIcT+Zup9ICdMZtVhdXBn
hAh6XOB2KemEGng5okwrG3EVWpxt8/RVS3RiPs1J9EQRxNcYMGCC1JNAaaHxK9uc
BMk1w2YjBK1Xhi3hXAseadP0jsrSvnbXUKyN8iCTnNGqMuiCPpALzuf/cC0BK+xN
NKeNJegEz2FGnF5iIoyaKwmxzh4Q/MfkcOhtnyrkxTnxuMtLRSVz2zIxSZDK7uBl
N49KQQPRUzYKr+auRUGZKpJZ7kH0ZDu50mz9zs+6an8FR8Qwa367AGzQD/AQjlJV
nUtnmSfv++1zTMY5Sm6RkP0y0IMVJ/y7LXrQyEoQkuviSelbxCdO8p02cQ2OpKGK
uaCbKrKM9tPDahQkRWpNDPLTrBGXkqk5haGI5hkVs6XV4flaLXai0Ta7btmKwRLA
YyDJKJwqXzGARcE0pcSIhoEqDZSkU1n8w32TZiqtjxrdZcGduvDpXJGuW0RskSKC
7hx2Irjme6a0vL1tRu435NqpX2CkLtKmCHFpkOeubx584eSfQ6oRB16oB2zkg9lP
B2oHV40yCEwcPdi5Q6xq1ZivD27fV1PKLNUYYp/bhpesuJ/k8VNiDZDdPJwqDWUn
zxfhKZKBYrp1ow1uKd9Me3o8AuDbglNUmgluaTnuGLpLWB4qY6IPwSKvp9EviCYT
uKOYyOMKrA7woQbqzxuSpZAzl4nAvArSLks6W8wCQEjORKi2Px1/1Zkmg+GySd2l
z2uRc/5+r/xZHnOElVhupa/YWqgHrYEjbWXGKc1LaEqV3RQe7tSUTDV8cV19so2D
0P0Z9WAQ8uYYpRbx96yrWyDSBsZKhR+wHVjjj3j8ZGKw9Ascg1h12kY8/HajnIVM
Xwd8b7IVO+vikpArC03Ae//cvARn3u6zVysuMOjxhDJgHOnNwNRYnG/cEnrAYhcM
anwh9SzaUXgydnM+T5XmFJAAGIvbr/z/HEkRZIbspCJCQOAufesscJXfgpWoVR5e
qkV87ebqEso4sowzBAMOI3hj6A+PP/+lRf1ApR23YeeNYossLX46yIXi3d+5z7RH
jQZUYSpgpfNCyn27odQQTfcAClxPMgPPc2rmGtPvkxERY/C8iGAz/lSsj4Tve9Jl
REvPcD1Q14GU654CTI7g9AXv0LFQAuMzyDjKR+ESmK5u4axTnWRV4YgI9q8GssYe
789VvkWOAzlYQrJdmC3IKgY/FTfAhCmnzXScWFzbfzW4QrOvFRpTYFrggblQPuDE
BXY5F/IAp65BfCbfLIvimaEvnFxHNLdLkDnVUs94CLfYai9Vs/uxeRHtEyAgthhj
ypVBQfEOPQRcwue78dv4oaw4FC3bN/cyVrVPx603NsD4u1zyU2K02EclnjSUBwj5
ju7FKELWwDT8mwuYW0AoDjMUqQoFLzhgCtA2Yn9COk1pp9QuChSqmBWyMFbRzq7s
3csupmt56nrI7BJ4v+EFkJ2TGbqIS9Gp1UjD3reQ10qVoi6RDcncpZUG+OiqnbPq
YJrsbFO6haP00XicWEp3/1g9lGCRn9797EgI1JYi0RUVcv9DdguQo07Cqd69Wx7B
QaH8G19TQgXHwaFeoGhwBgLHkg2p+2CC2oxkCtQojhnwrLvm2NH6L6pNCIc+O0Ji
mWTINi4JvZKuwTH7Bd5u7gEi+NYqzJ2CKi9MiZM3WIcIkJTnDFN/N8ua0x6fyGEE
LzuPfsfBf5Vn++7rpZsBxRPRZLpxEdPjTSTH2xg5yNSCc8V+wSXRWTZp2j+JdsDF
j8X3sgw+JxgR8xM3SwPfY0hLeJR2Y8WiM2zQOH4hT6551tAwZqe4XLeE8VIkpTJr
Wq+k3koY7Yr5i5osLg0VBeugwfMJM3Xzxg9/gcnx/X6UDwe4EBNIInZhto10OlAr
n4u+XMvaF1xunjcb84TvZK7MSzH3Lbqv1t8KxyU6NYd35KDwdMP1WKL4wYLjW57l
XGov8WEQw9NU8IlXvZPZNg==
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 21376 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/T97rZhQva68T7JOm4bkq25
b4BW57ADAHEm2yg/Vzsfl7TOuMe4xzV7rdHsSWg325sjWpFWZVqfqawtQjhOV9Ti
xjsylaiqHnTulnIowKyUkoyU6J/E3BHocHBw1HLmpZELKO/XkVV5+qC/Okl0Nt6p
sL55m5vHl5G8JtbNpJDh8GdyLods05RwSew7j8ZFq64fppRjMO3gR7FsxFi6hnn/
I/mFXhYsAl1s9wogsqF1aYh/k5NnqL9W/WGqhPwr/uxfwmJhTX4jOrVP5skEQ27N
HaDmAKO/FZzaXVTFwXxWiOxBvdYGyXtJgWs+PK8adaiu2vV3bmWQJ3Psz+p1Y51/
fLLqkTWISKW1B2KmT6Yfyd9NTQiFbHQwoCd5F1gDAg07Ogz/HSwPor5rWNCZV+Kd
SMNNFLwWpWWwTmw0DSjIOrL0BufotBm8QGh0I6cT2v1U6B5RNvxL3An0J239TpLM
nE+okX1072T2ZQiYpFTk5a7YLJEPNyv+ESd5xwyyv7voWqmWFsulXsGC50kaG2f0
Y4zWBHIK3fuh0sLplWu0J+ZVgvtXCWfCSclCHIIKAXX/i5eSlSFc6JBzJkA4zgOp
mQwWB/rY0O4R7ECJea+TbGMcXkDdhBxmfnMOUbElsvg+9fv1oJAQc6gws9jp4+Pn
LnzI0pJZ24GDCNHMDLHl7fhjy3uxHwcbf4LWLsfrv2k4wRThpVF8GlRj1g/YsH9u
Vr4SEyiWopm1A6BEqlb8b8ZyciCotk3WgZA1hFMZXXkJdUOS5H/kQQgHAsihEWs0
WUutRlvyU1DOP5nAGaxBzR6qo5El0kDuOphfhp27VF40ye+0cwKNzbz1MOTuGkNo
o0pdJ8bcSJ9B2Fosjll2v505go7Ks7XFbxN3V4J0eNW9e8kpPgCGuLcFdITF3cwi
oT5/o+vMc8uPRBRb4rsCInhzfq/XSPK/JivBvSu2qTmGh55qw2u60Ir8rDewBXGE
c1Watk+6L3an+FgPqKQyfCyDYHlj+JxkrD1Mu8rVwK0TX/5VyWijZYOmeSEBEAUk
QaRdUfLCaiFR9L1wEt69Lv9oTt3mzUwYkwABIvls2b8rT2p0MiI1JEw6lKCTWT4b
5Y0H57Jm81EBmvLl8OnjRwnF3016Jc/XHEEa68PrrrwtipRZEkKAm1KdmWqHjKhe
Vm4uq0BSnipTn1qU1ZPC4/f8NKt5MdfJLKWHRku2CFTTH1OV5DrbN6bXt/zAGdpa
uflIiLj4vSJocIzVPqe0gIJFOJlccnMfPD3+lnJXQRWwml1t/0Y88jMZYR8lksSi
rFkmKO0Jks3OGqKgBFSQMdifjT9FSPIjCLneFJd7Oxjd8E27FeIqUUZObK7FMOTR
PfrUDxvgYC3tNJYPRJYoQ6qi3MKWi7f5SxaN5b5lpTkyA+TXinV9W9QYrInIgree
RnMBd16epnUyssYyhos+cy6yFlB90Fzm8anE412i4K46OjOQo0Nf+NEtXXjo7Vn5
QBCdvUV4olE7A7JvR+tv7lxw/lftqI74+Cccm17RneO9YM4gF6rcPHYDEd/0qNuU
NYKAaV+kx6ZNmM9Rk8YOjsssjgsGzctoORiJSnA09VS0yNraYKYIL9bg2whKP6i+
KHgxtv7BJtq6v/RGJfdpPqvN8Ca9fftTCpzpCUtf9TdCzJ7i9RVwt6nrXI3s2hLc
xjZP1HksJJZzNY95Smvf3LAn75sgWWICs7fESF6DiBotLcmhoNFu6IHn8whK+f6z
8mDVj4E+FOsfdPAhZGFOwNmf9GCzd1Dk550uZPyM2hGRnNl6gRMNUZiOiw1PdKPb
r9oM94iy500dLOtlQ/eCBfng77UmjZ59VnPdY3AHMNPWTCQPmVxFnOHYn9ayGVSI
kKUrLPOXytMut5ZaghJi2ikIl37L2PhFo+JpKmzKKBPL8JMJpRwW8SoMEHaO1SHJ
QPJl/B5yn8xtVpS1rflOsFkg0+6wEateuG6gZ/MGXdkYFkL/9/eG1Ft/Q8xEbDfc
MfBIXGZK44i7FZqvFMkD3cC2MLSPbKYHBouhxnhf71p+C4JBOb76pM7KXUjOZYss
t3aAa0OBtNEcyXdsjUMmQ9AW4w5N4LekjySIAkjE8m+Eo+0TvwAETbQ0JH1IidRm
rYfyUptJAMNhNbVfy0OaT8OCq6KxlXY4IRHDW14tL2k2/2kctnwl7MXOLpSwZKOi
lXjfcDTlMCR/rgWrsDL4vR2NMgNzWuh3Wyay7IhGtuhkk7HOW5W00PJdHE1boMM9
ffobYnX9pqOvbDwyq56s2+cm4cz4frCE+Lp561Es0886jxWkSp4f4oGB755ls6/c
nslfAEL+pnyOxj88HVMtf/RYweCSFNqiPfspONwiqA8x31so751fza58S3+aAVdq
E1DHJVRAv4HVPRFWO+N+WWYQ3lmJXrtLmWlIaIr5EEtY/c4ivztMaqm1gGreM6DS
HMoS/IQi8dq3QaI5LPFzxWV/B31OgG/A+Jpxa1gty4COGCWnmW9Egqqe5P6LqwWe
giOOyzsV3D09AWYP3fSXB8XANfW2trzdSSuEXXE6Z2oq551ZHYIDsZKQH92f5eib
3Ep+whI+/abpar2UZTFUFhKPX1X6ATdOOSCsNCo2qkvjuxPuFqRw3TiMdYrYkTdJ
Kj/QOXC4bytMj7lS7JunzKv9Rljpeqfq2O2/sH94Hu+uLz7Qwu7uCyIkWJTen2EX
sWuHWdbMAicYnrkjzZ5eS3O2kWlqaqJQqcAMF94CjNdI9d3eylT/gUtl6gdOBBUM
4EQdmXEh6U/sJh2xbc+G4+ktRDpzE3o3VARPoX96sjJutqarhSW3X1ZgEyzsGExM
DJfDtFQq6fnlglmCSkcEciN8N+mOsFNrYaD3WFEZek21n15McwHWivjtZodBWtFE
C0uXWGHr8YYItZABGljwhyWuvDwQvWvjej/FybTcTbSL+Obu0x3KGVUP97RDedxG
eF3cXO/TNANBwcFueHqzPQKk0+CfGLpeu0NU64AD4+hqMpLjbiGaQlW37+jkjolc
qRvEaLd9GHa3sjIR49GGnDtVoYI58PlKw6x9fV3HBurzqyISAPX0n4dH/1wMxygu
6DfoUOUGkt8h7tsPjLO9oI0jlRr59YPPdLoE/oHZIF0OnxijFmDlgsJ0juzdohoV
Ggj2DclYNQj9BOtQt1s22lVkohAGHHadIO41JongR5cBofamc6tik7eWeSgzr42x
0ztPj5gzNUIGL5vacrglhSQ6GkGzsnw9rlhnPtYdEMHYEfKQaOiIQ5uTsGOLQZYJ
v/PKFw9JmhWVaNToXm+1n/wUagoSoeMq4Azr9CiBWTChiuyevEbA6rnnTl/3M5V6
wZe6V/uijN9DafTaxzqxoC1B4nwVIN3zCvKHdVNUfjLWL+qO7rXG6L9yfkEuXuco
6CHX5rptcmH+LPT9WuceINzUGVwHGsEM8abf0Uc2mugodZD2r7oSHPFLR4xOR2Lr
4dEWbMbMj/5tMUVKnK50XEhvqHXFavMCc1JDwxKfqBsmLlShlNgYJznn9irgCuEd
/CRbgTklX7DYnaCft4TtLgGvXdd0HzENhabL8sSEIEMyL+MQ0yhitRhIEqVSwkzK
ky+j1+zm9yiQdHJjGmwQva6Fxt+jG4GyGVBevZa6VVO7NyQ+/jzNqgIXVg7awbFx
2ANkdPa+3zFnB6/rL6Lh4r+A/8D9QKZSR9SdT6czafWoLRZ2oeVAlztdzzGPSLKv
f+jb3qz5BNbcanakoKULnCz7C4z6aoMOsn9fu44We/H6iUvcEFqhBYHLys3f93wD
e9K7tGczLuNsk2gOBjRVvXpulrFKnhycW6cr8vLTmQ0+WjtJY0i63dIsVNt4Dc9G
lvAnQz/c2PAwsbE4Qg5oEYutbVHvwcu+lRnWblZVC5oWWhFoSJzojVryTJmLsK65
z9FgomVz7foCpsUj8ISUxOfnx/MmdxR5SMYU2KAX7AtucBldxrqgucbrUjOjZD1T
xT+meG0l6y9UKovM5fgbMkaAUaDcsclx2oJD+/E27cOHiYxxOxwhCbMArGz+ia00
sfrXS5yueThVMb6M9VSjpmGBEyac9/BtOrFI7dDFykm4bkFOGfsH7YtEeoOlpfuy
sH9TpiFeMEdOzvrDxZOYXNvxDvb5aWRLK9Ik91R656LcsIQ+KjfJD0tMakMQH+xL
BhuAV2Jx3bhrkuhsveP7jwl3UFaYVf9tGZ5EPj49LoV+GNhjszu20Edf9G6f0XFj
mWTsY8AT8izE49YXqI78w6kz2bPXfQFqM++GfqgGnLg1D5tFqk6PMNq4UDIOkJfF
UgA/Nj2YOPQWVspUBwW/1oLaUMpvg3naTPdalAlPcBtIEtGEupB+ugoxcI3jdCpG
BTyEvzTFYZPaj5PbUkPTRisRccoCX52U0ws/oCeyfUjKuLiuCRLs6oo5U5v8VrJo
lOL5DZE7GEq1M//IRFMOO+bt98qDYoqFm3QSi0mfEYDIQa/Xxv/PrzHxUwIINojy
U2jYY4SjCsLEi8gB5dCNVPLSZmpQkfwpfnPkoaaqeVg0rryTprzX8bFiHSXaAb13
IL4DxB0cleJq93FsnfDv31C6v9kT3AYFMdEsjkQkNBIRbhb0rLqG6qn2h+p7p9e/
z+dDX/9lMLbILl9VDZWekF0QRrYPFZHwp9X6Xc0KmatUPw7GU5IEjKqwDCWfwLpI
7yYfGFJEFliFONPAxcrF8I6Lvomu/wm03z43RDOjP/pGK4yXv3fJA4XsRUy0dCcR
4BEkjyNWOpHijhlqpLR6bYkaA/v/wSJHieGFg4U334ithGN3nXEyNSugTwDURPKD
ZvzFA5YCC0L4MHjj5TeRN++y4bkmDHJgYtqI8LPwZeVC8ywos6btD4RITYqkhQPn
jf0+9/EMu9qPGj3qDmH+7p0+lWutrgK3x32SIegXw5jeqH3G/+tZ+qa9mgKdUsXn
Ug6R/LkABXG8XUwwE+9zD/vcPGr3QWjQAcBiRg5x52K56luOUFMtJs63kFhSlkLm
dX18iCp6LOaiGWJXkEi7EWewR0+8AdKgShBqBs7K9apXHB2A4Yd15ii7oPRGKl3z
C9vXZrSV3u/R5fUjhBw7UBo39/V3fvCvXU81Bn6dgbVbkmZFBHG4BkyIbuyCeIrP
9nQ/b11rTOnx8QYoxuCoZoISSrBMVmr8pm5Jr5vCfv5l/DyEjJ/5o+730Zdi8zSC
U3SlXpvgEMXakq0uLGDMmd/PY2g77lZ0uMeMrOY6xSprWtb/twWKZL3Afa1BOQ6C
K4gKOfcNGrX8RSUQC/CRxtP4FhDqIMp/drwj1r72/sk9gyI8CEU1m1g+MjdQw85V
quNDwtediBg4Cc5trJrxhEJPMq2ck1LfAHZdnf8rUUgAAtCI4GD/khLpTS+8AKr3
mZ7tXijs64Yh++RT+hsuY3ZZQyjYhqrf2q6FE77I3LClIzoWFuIP7uQ6H9boewiI
C1BEKH7l8f33kn2JspnOMUbLNxh9PN4YKs7wZO2UmQLP57t29XcJ2lHCkDXyfsH4
k0TP0Hf6prjSwn/Upx+XD5gLuU52m74Todfk1UQzS5II8Uag01Z2IJbbk76/fLvZ
XY7lVUVVgn1EzcuX91hodUA2mWdsVC5TkC9JcGcMdkS8QeCPZ0XDt3U5K1XfizEI
NhBz4O03nnyjFe4Q0g2rvTSgEQpdqI/WuxGlrbdfx0mF+t/+MPVOLCh40Hll06a+
ZWKtwi98iF4VpMb+xvR/gNv9bwxpqfgwjq5xoL38dP5yehCcvLJyh/SluCjYOBJj
w/biVfpYNvFfTUJRbFxVRJ291FC1nIBVb/zk2q9/00NbY9QcbvDVlB6JjUZizwtg
LrNQmQBRYA08MKI0ajbHoYsvz5R8Pu0V/4/7ywuzn5jrQlYOGBoee7J+wLka8JHH
urF6rRKoFpasH+TOluI69WC3Ot8fz/HIaFOgR5yDkXAcjncpVrpAW1GDKinVVY+p
uR8PJ4r/Q2pzT5cWD/SKPiHeYui0MkRON7oY7aFY0n/7vwbmrn7DlAzZU+9lN/Ml
yf8YS90V8kdW4jreHrM3/FV9ZTghKN1waREgHLTxrgJURp1/hXyb8IpPBa+GW5N7
rf+ogaGWvJjYkTQhEuSxkf58Tr9fSSs8H4ucYsYTjPIe30+6lkgoH15aNUpMLCFm
xzyD1kkHetSNtdN0MrvuvXIgd3yI1DIh8eLZv6OqYWzNSbsKFphc09FytaUhydxH
uwAQkzqh0kwJohIi7F4so/WjFSziEfnA6E7v8FKYgHWy6qivYQp72bcp10sjJGNP
ZU+nUK76BIjBCMvXtNDY2HcNLX4VQvscDv99BfgXJi3RsivAfU5jg7cCYqr6mXFz
q8c7E2QRfI8ITsIkBT0bW3y8MZmT6GsGgSGZtQNDLT0zjcvm3xbFXoW0q4GZ0D3E
s08T9rno/K2tYkY1kiU4/3KKH9tfJ+Lih4LppqJTKOdOSTHmGIHnR3GoSolStXMs
cJWJ6lb8Fy+gUm0USV9KZOLXrPdOrX6UuCtJ4ECSOghRXsqHcpjKQFYx17RPNOaO
PE28fO6pft3VCiNmAwoY8H3+HdWlMqL0Zj1P0XSC/cQ4VPiJw4UWwXSGMCpHIj4d
0cJFKdWvTqSmqewIGOnjPgW3Gll5/GKw5FdiSH2lEKN+VDCQ5LSRGoLj7oke0IUi
299PJWG/2hyZaD+IWU5qxmQY0pT8yS5/+CcOXTd2aXLsU5068Mc2v/pS9onildXp
rgsZMeyNDjiBuv2LCvvLIgW2WyIPiAn4t+VAo9tOgQ69Rvb0mNRwjYAOddfAyPtx
w9nRnhrTpKMvdzdz/GO6TCxS9LRjfNbdo0sS9Q+tDeDUrxSx9iGas7ZDj8+einBO
i8w1mxM2/2DBYrqvjxg/SL9mvokzPIx6YBEU6sS4by5WpR735x/46p8WqNtmW2WW
bUzc4ugWXCsjtY68PIZ/RZnCedE30RFwIv08TzmuRpN6wU8h4hOIDgpP/sf5tdU+
Yy+icdkUjxt5bw2HINo54g312mgcchm0qhDXWqVKs3IGTZDbf/Zh8FAF5CAwCdKE
snpQ2vUfIIUGvl0Ip7VgJagHORd9j3tuEqWh2VYyIDIkTImkl9few7H2CtJ7Rf1G
3FhpT0chD0+cBNY8vcGRAhPXoGofYv5LZuWDpCaVqYQrE+LC8W7C1GyL2yh0YwKA
IvtlLj+6495+/j07F6FvzVcHm/8UgcUReWv9RSlKmohlUvaPJEtfz+eTn8ANKmMa
7NB183oa/1xpJSJ1/PQCxRTf6oWNXjPq6H5P7bLnPa1bZNDuhHs02jGuU6u1FCCM
9r2QArHyhGM5Awoc/3W4t4kq34RisvcFsHw91jzGjj0CuctWKy+u1fsgnWgMCic/
JEt+4D0gWj368PXEpf1oNPIzsGJrvkrwS6IGmOCZX4iOr6GHxr2QiUROfzPyTNHR
HRfq0o+zJe+fj3Z17XTN+O43cy40reqcyXkvsQ4Fc2FxTLw5/En5JFwBtEv0eG6n
MWA4qnrb/VCyhUcvWIX6I3TgTF6qeKllAeCeaQSnkOqc1/EIDTfZb+Yv96EYD2PA
OhIvzZni82ggWaM2oh+8jTdFNfTpcjWiCZ2O802QTEFiCnWWlNRxk9D5N++47gxV
nDM/ztqC79fCEWYW/jwvlD2Bt+OQi2VKpwXW11OhDNBJ7k1hLxMiaH2ILjL02lSE
ceXpwHgBazCZlOJefeB0g7lOjMgco4ntq1/s2Zr8T+V8wNryP6wYFSsUOe+zlglM
aEerPJ/gYSkX3R2341sAxmlSRctL6YQaKLx/ZAX7dEugbDeXiW7xZDT7+MPUsSH0
YN2uY9+1aytB4DVWNVsvIpexcO0BV7dFp99V/wNCtmXmoJFr2eJJkj3IWmqCXyuA
2EwLiGcQTxQZ6RyoWJ4FrVKKjDLETZFECRlZgTRV+yEm7AB2goDVkxSkj+ipP6Iq
CRS3sZBWhaDJ0ADoclloRrQYR00xDbv5Gu+/2prZO1FWyngydmPTayfEb3dUyg0U
yLWRbuYoS3isereIItQaYc8Ms11OWMhQS4JxVRxYtMl3X3LdamWlXWTnHqHzs/gI
wzmxKCPV9wn00hxbTvUeIhzWgO11AV+ByLytu8+iOppc4f3sNHw49VK0Y1V/wANp
khRW6e8hqagiKadVmLUN6T2cNKg/v8V9ao03TqIY3kVMJ0nme5YHJhyOkmgELyFP
vbJdcbuOtixEPih7ec7NjHgcNBRMAHGmjmp3sbJDD2/P6jkYJTT5TPmaGqvOvX1u
/B+f2yl/vm3KOy8KcZCvL8ORTwDr+qBUfvAhiloR+Ur8IenovG5zvLQT8yMQF6XN
HS6HQHabZdJ4oGSPvmNFi7Yr4TPb9U5wMW9eVHBHBZZkWicT964GCTcBaRnF2vKJ
R7gaPeywXlgEOoLYPNjQJRn+x+AZRlIEYYxRT5C9FGHWf5LWOb7W0eEk3klleRoM
ciSKkZHLNiHco6Xj9AFJNdiZw/4uDRa51dKj12qS2qPFI6MB3rJnD8ywbFVAh6a+
+M1DGukb2nzu9aU5Om9y7I34UBADI6d6NxSAMRXLeKUXGT0JX0kTgXKZ4aY0OO5r
TbhVBS2QI/CPLIg8Ti+x6w64OqIMO1igWMW0SZdsnNZkzdRE2FXxWLqFhOOXaLYi
kEOiHL3P6VpEhtbmSryMsrRSzwJ5lgHNlnd3pdZJHq9PnGX2jLhGUglzj20Gvl3K
Wsu6K7TyaCtihhEfaGjnXPSH6FKaO3z6oAMw1W7/S+LFRenWIjrT9JeXHX0wcRIR
j1Xq8nu2nlkA/X1Bg6McK0+vltj5GR42iyZYOX+BXuEKI9loMLcThaaxD7PFMiAc
vvHTixzXG0LcIdDJNV0FcCuDGqBFoQdtX1VD4sFcEKLhd9qA4FFyOG09WA9W+5Pr
cV4IrI/39obIAX9ktoPrCbcYY20KsUkt3ZNAbepfIQNqsb+QCT3G9uUD94QEBKTO
CjKF0xaF8pX1lABXdKyDtHFhCw6qnrd0hXAQ7uK59LILZpesAv5grKsV4Q2nWEWh
xLBP4HdGf3gZGjhY4SwuVUebHlET93r3JSsB8Am457J8XezMjPFBcIv6O7SC1/wj
+LFFqZoHwBQoqSTIWaLNMOya+0yocef2rgAr0jQmMHlpLrXkYudqTTvOA2rVc1tR
03d5fOqnew6JJfqsGkEEdT6w5jGQQVSEm1xcms/OmUD8AGmVK9tPCAKkR9H8Twwn
UPNC6uNJ+JaHL/NvXpUHfqPukyrBNs592dA6KlzXyNCsNgqyasUUzHzZPIZ+gU9c
ICwFAB0EXP6BH687e0kYdD91oQvuWkdzhFf83k+ppN/7n/I/9m8AMjtDvfzzOflD
vI+XewwBCz5kuxVDsp/ReJPDr0BB73kfa5vPNCMLPI+3rD4sqhgArMglJ5nrQPJx
sJ72nWAV+GHYR97uvEfIA7Q9eautWE5kTOJAiwz+I0EfbcjOKsGSQlr/3pbLL778
0ABSFgUqQMPApr9L3Q2mNWYN8EA9f/Xmpnb6GqOiigpC1Yq8nh3ANtUNkoC8v7Zr
fU7FYugoxy9xGiexK1zqM3pKcAVHcMZh78D7Tsirjlfz2NcsZtg08FMcMbkDjaEn
VWhfUvpmkiz0WeLZrlnnA/o8DeXJOzdOdQK5xpc+aW/Ke9Syfz8fNKzpae4DOWgl
Dte1W1zoU7WZVuHL4Ni0tsngB/cv69VyZ7Qd7p5Y+eoK9II33Qv5J/rARbFKCxDq
eGCLKLgIc/osSTcBlBakfdcdpSqIricVJsolh+EDQC5IKDX6tYxPgqPuIBLMZDWO
QZwl+9GPLXAcvaDyfWjeXNMpeBGSvB5bx2ertYbSiuxXjObVLp/FY/DYy7Ln/woe
rIRlByI36Bja0M6hW+18Ma6Iqw02LAwFHymeiiHXp2v3xtrHUYnAlYKs4JRvs5B5
ukr8wliBShNscnB0VsfEsReY8oPAB2jVn2d0ziEScrqeEwss7JMzCxHh4w5/l4jq
aStcbeTkZ5RxNO+xBKWIPV6z+FxIJ/J+GeaUfzIgkXoF5r1LawN6430ZdH+o9/yT
PiOU/yd0uGorvsRKWTKENkVjMAI8Sc50H+QN8kQKbfdu9ycUi8YAMZzGjm33lGrl
Bxb9LqHxALfzIcXXaA1pC0o4SIYgA+tnDPsy1WB0SvCVwbCz5FGVmVnMSxFj7XG9
zKtpK300DnC+OsMGF3EhnnXdjUe5Yi5OnVNt0YSPxSqhG5SrZ6Rkafqvqeh4tbfX
lJJXMMu00gjcheiYpFaa3g/NcoNbHp30f1m33LsMKkQCtyruVpJeoz7yKuRuE7/Q
Z2CjjG/oiUc/OkR/nzLvtjEXsUEaozTr9cNJAkV4ZGUHhDj3XbNjetcVtOZL7feb
a2DM2lGz+04kQavufO2EQB1WhQWqZe1VZMncPGY2LJV0hSY+s2pEIKlH/5iBiQfF
4816KVF3R6SuIWePE79tXeFcgwWCXJdWwDoXp7yJ5TCiVOWXU1GPkoGide19uVea
rh5oSYYXKSth/uLopLmHerNSaZ4uu9XX7nA5BR/dEyr7J9eybuQYPZrLy2rZ0pFw
F5TZGvH4yjGQ8vevFbUfvhN2SKBeuIQCpMFTdmcmadNQEQtXE1hulMZoUR4/HxZI
j+f6OWm75SbEpaJDmJBL3P1zR8ijJchauHfozTrchqx6syHDtZvhd9uEwp4GXNIc
yKFVeC7fIKk6HIxmT8jTS51MK+DP5YtLT++TBvGQq3yGM3d4fPqeqimBCpcmJmu/
qwLZkXwJRRfQRYRrZSRgIkcD0DoWXodoTrq2vRtfWLLYh01fm3iKbwWtwXgR8/rh
yHwa2q3sjJtYEsi2F78pC4NiwjTat4I5lIYj96ogTS1QHeyWwUceASvjawLveDSU
q20t4Xwb34EK6vfXF4Y385mbgrFIXlx3LmZ/fwdjIZPlemDTRDLHDMJyEmhhFxke
ChD/l/nN2qAwfQjCiiTSCcmw2nouLKXRIekBwRdd110vHkePfV70i08g6D5v7PKp
2hn3rZyQIUB02aTgLQk5DyTI3i94m00uNtplRQNUqSIkXi+E3tN/pWVhOUu+7JDK
DrV3DLxrdxTUzXwXwlc/JacaIfazk123WEgWU+FCv/QKv9X5GbHWAqPyYtYU1yqF
vy1G3R/AbGVGcmOad9hCbM3p2tzkdbz9Y3sqCuN4rBYRJx0XQsYIfH5bvz6y1PSf
UmYz9ajTWxLLh4JFbh5PhUN/PclubOAoEyzPTUZttjCzICDcrNsPYmwfdYQBawqc
ot/zqUTzeCdHkL44YSUr9tcX+EXcD3qF7p0vy330z/PHWu8YRH+YPQ2Xf3T5ROYd
fmlF8mNSTfGh20OjoRiacFSjVxwmIvhWXo88wTU03sBkFIdHuEJj8OdcUcU3Zl3B
7NBJ6+sawU2hrEZ9fQmMAPpD5ti67qWgbcu7EpO8n1yI5QzjHwjWEKyP6EZl7xMj
e3i78YeO3wkL1jZg1EtZy+7kpaJONQwI1+Hick2iIx6yVkm18m1SqJbidk7+CvV9
0oDeiF4g1gaarpQljdLtkVtgGIbIf1i8Fd/bP1AYImUZ4sMs9zM6WGy6UIL5hqOW
L/ZJS5Pb8kv2rdi5kn5Cv2ZkT4WlQpPmox8DJEhsyq3bz+T3yPH2OG4Zm2d+bU5/
n5J6vAu9N6BzuQQqUL3fz6uYQQc274C50qQffhxocz8vZ3wa3aP3iDsrqsKzd9+c
Q56zbZD8flE/a+OJtWYahcvpvrh1oDfi/CPlDF5GlTOyzbxCeYWH5zutabvNppOM
/16+I0nQHUhH3l/Yep/LlstbCPwZtY3O3NpZRpNjCfuS1upEfsGkoK+PwfcE6Ojb
WMxkV4Ocd1vUBEm5oC89Qvvx8By2vAv3LtfvyqJ4mvMV2pDZ5+RoqSyjHpQ4smHR
kAI0Tn1xJm/8D07O03JhxgkxEvWRk4a8YOkTWklKUuvRVcGlUKfdHLi6Yy33xEi6
+gp/IJca9TjrL+x65Dn7ErupgcJNmCJPwf8iWtanEoQr7XRX6FCskQd+t/ydra3m
thcbaCAc6YKQetEAmivEgma8zQj3zmascblBrRgvI1XlUPkycJaZEqvToFWDnXgp
Xs8AYFFSMmO7DQhbN7eYm8TS/T3hGNxDYuagEGj15kw26Epn1gCWDjOeKxWPAP7f
5iifkmTcZve7IGznXsBNFJejFy/ODTs3SE1+5/SB6cUGhiJJI53bpDAkRpr+gdrl
1kGRIVV3m/GPWHeObkO4QZJpFfKC3Ff9wwzOv51om6m4Sw4mXwAECq0llDpvN7e8
Wjv6gUqk/mKi/ouPs5LoMOSCSjX63ReXzm9TLsTZbj2Hpqqu3JoYeQaCnC5OhgrJ
aOWKOg+Hql8oK6zqhThWMFhu+cRC4WiQUwSUZDfGpJy8Xfp8wyEEt2y6UszO7+UI
iyXGP8mEWQ/EWujz9iXwfTV1yZ2z1YepySWzGqA4lfjdr+HQ5Hr4cooS3Nvp+3GF
d8VPPOerXCf0vtTxIYE/i1zIBf/XYPBCaVmM5TS9tbqWnQCnizoO44/zKQogb3fv
INvfZdKh/OI4n+uUnOImtRFYgSj62pU4LdszErL8LaLzwwoNuNKoCOloIG/JFVHH
jQOS/TKMz200r3e15zkhwoFAnTi4y0lOrJ+jhb2wOZLFaiuEoM165NQWs/AiuW0T
0eudBMwcJ58XWE/Zmya1UUrlK2HipoCOsqtr85OANEzM46+X4x257yISLFH3zeQy
gYfh4rqPnZHU72uxuECNMjhdas4MMCtjICq6ebCb+ZHkozH495W9OWELVDa04+iq
UE0ykiC5UgcP0BzQPGGhWzeyF1/JTkT4/gjwpZXpXcxo3tkhvun4xkuvyeb3dbUM
d5yO4m7JVZoFeCWCtNmUlUGveYXs/+XJ5fAQOfn2F3J8jb1YCOfOPwpE1brbSW/M
nTNtOLMmc9hxEKvp/yt1/nWNQMoS3cEOnBb6fP/Cl2iHkZ1yFWbCTAmXcJk4MhVF
V2BYwRYEgeflTudq/QPvlCjeJvNSxmmaMJUp0f64KEFVwZdL8sewbHhtw3sDZxpk
6E96YGFRFPhi0DlVOj8Oq7GG0Jg/ulx+h1y2ofwzwp7iGj5E3YdnnXxcLHR9ciLc
YVXU7RQ7ogvvO0azpoQyeggMfrg8Qummh5Hvq8jQmkAj1ans/qFWudjSe/ZGO5ql
Rasm/dJrhyW5brdzcdTA1b7gyOaH6vBCSuQa+AtKoMg12sBONUNvOH5LiQl3xfI8
sy2mPC/U3z6e0N2Iv8/mFoO7p0PCr+amLZxCPDq45eUVfKRMo6Mvqvw19e8JaiEP
zdMjzO+5YBjpMIbPXWsmcDlaONkkIr5Ic0N0lqp0qZEMlcKOdn+3TkRsUGJ2ln1c
WuFqoIONQNriALKaB7ikWF2eqXMdd+mYa8CDL4+ylDvyblK4YXjyVdw5O/P5Yria
88p54OhmsVgaCpIEn3fyVKj4Ie1OThCwv/9uHaa0/fpq/eLP2kucomLJpLVKAyEK
/NLQDuSXQ4PhxtzCyov9BSj4M2alF6co820LrEK6Jo59qfrY1iEi8HvT1PEeztnJ
RNH8QnacuYVgPvpvuBsWgeoPbOI02o+YKDVDvvR2NN7oToyy2DiatQQtgljRtvi/
y8V/SULch9VFJRBFepCeBCOt+5wy4zhbvLG2l3Eb3pzBIair8GBITMpg2J7hsBDa
+nEkzWvEg7ZqIOvK5dU3mg2mmvCB7wq+KgUsKSI33htCs/NUMFzYoIF1a+tPoMuA
wcTGVAfYoVKbjSKoZpBqC1uStryoiwGoT67rjVcJ+u+2MYrAqpQ9nNGXKTt6z7cq
A+Fv2edpWRcPRYr7fvTCahkCCmN5hMKwMIgmRrOeukodbs4mHvNnpxTNE3pzhh3L
wtoIZWO1CMVIIHyADpCdHJmbrrsCMwqn3XJlViHbUVOK6rir7K1/YQ39BtscHOTI
I1R8Zh51rZypGs2ntPRunYconGFZmx3rL7tvi1iLH9p5fNWuAxBUItMWby27cX7N
rkp2wU48UmII/RQ1Taw/evoL9BeruPz8/Xqkf5iPYXeCnqXLGN7GqD6KhKul+fCN
AqpBHO5xWWg3kaYiDkWj3m/NsAVIQ1610B8mBqFYmoZrlf0NhG8izi3sVE/L6dJW
TvoZ+8jXD22J0aPmBSpG2ACflHaWDmXmqDtDh/HEZxtjJtdH7OTAfIqiQWD3pOi6
uLmjNtDDL4BoD14IOZKjHuB7fG7N586PGfnxDmghCDiLn0ff4XKpMlX9nUeIdm6p
1pnEhKDeDyxkBRfpxlNRFSjebxXyr+0nbc3xItNeTKY9dGaUKRIhuqpix78faWyo
ukYR7XQHNA8aEuXOUb2eLagHPEax4muGQmex7NPv1c2JrxPX32M/B1RyLPsfcpfz
ewDG/UUUAJoIEucj76qyvka7hYdXvbowPSfzDC6UsX2UaVX/R68XqFhNQnp+e/gS
jQg9VgwnG7TdHcZQfB+Rn545OFq39EuN0UHDQ9pMQgk7I4qX/GemdIS13S00Nh/K
ZnPahd6uoqVZ9DFZ1HZh/nhsuX+YwrUSYmjmlYxsjNuqfL8BW54QuYI1ARZG3Ytn
zid7bJPn+XQhyQB2GPPneybgUwiuxmfuh7ehatbFUlxoJiuelq24Dn+rxcFsJbc2
GELJQUbSuHU87XPP5O6mhi/GAQRhZ/BP9oW7B6dx+uXomY5MPQB7jQU3hC9Gptq/
fdb3e2ZMXrbxVCfbfbgzj2PRq8TSmXH/e7c8uwvCaHcmUtupagYh1CEyENxVEC4b
e9VMxaceE0G57xLWnAWXQZCgBuUUYWXFSiwbVZuiQKiJUD+d+COrr5was4uFJ1Ns
OC05jeQAfU4c4WlbC6QBE8pNLYgzC0dKnGEjNf1eQykdrJwYFQB5bIoxjpV6lnNx
jTKMIhyMg7GhLNy3ZdhWVz/AGHsBy6vZgC/M9z6xYK3kxpnOVZfpauwEW61ZtbsY
JkGM23zGQmPRns2706DO1+Y8/c3RhU8GscsolbA+r/CWnGQ0+9d3Js22Uq3AAXPS
eam6h7Zv2ENNL/Ro7+B5YGG60/XiLpteFMUsTs8crzycrAMMZ1cfa3JR9GAfk7HD
YqMXdhDor6pCqKOzbKhqMCckMj7oOp0RYjuV1HyA84uus2XBTUKlWKA2T4Lr3pcZ
yX9ogH38koBQYgkfJBU5arP5NZthOSZL1j9aiGGNR80i7Jkr3bpUvfBd78LC/dfO
oAciLMdr60oasVxwqcs5uUgjz2aDzBHyIPlyTlQnpGbCalikriI7pnuxhQo2hgtg
z7URPvTt2HEkYbsjBKsHLPuE32ZIA5ZXCsrpSMG/wiaMbVY5CSkAFzS9+IeePHjH
FKmrmU6O6HE4w4qzF6lXJ3TvpSHyc4hA1u1kTdVfJDrcpMMQO98o9IqEIlx7HhUq
leIpScc3poAEhCjE2EPY9IcPT5awPWFaEahba9Ft+yb/G+SbUccl1yHK56o/nJ4f
lvTCD7PyNuONT67KO/9bySEe4EZilQXTfyUSckujBxZE7thqABhJeRPraUeJZpbN
xE5B1ehWJSEssGskG3pnD3MbBrnTAcX3RYca8lD0EjWs2Gt1tGBxwtbGmenDdVqg
ucYa/oX+WgtEIbGW0do30ERTbz37amqtWjiS08zT45Bm9lFZXSJE7Yg4uFiLzLiF
NnqBA5lDjQI1847+5ydXkkuRrG+7uop3f9p/G8fmLShb8/ZdKWIXQ7AzYZeouI91
oxAApOb9VEv5SZ6Wz2C/1vTwpnzDVe/hsIizUTSIhcbmqxMsjkPgO92p8VQOx7+K
ZdVpN0OEDl7J9huVtanebYVgw1Mm2BBj6hbD+PHJUA4fvym/XgIBjQRL4rnKzyP+
e71wirmdvZbmec7HiqMDJLD36gcW0I4CtL3XoHJ/ZfPlM61hcTpUhLnLk/k+bvoX
sEsM8ZVxNra/g4zs2vwKm+X3PSCqloy6dcWurlb4w8TD+UJmsSRSOOdJbG8A7hFW
4PBOqS1Oj2zlet+yj4BY3P8+v/kaM7KPBUvmGSOdZ1L209z8lF8ZcpQjQngCzuto
eUQVA1kooiYsrlI74lYHERDOKb0xytTdhledww+ENJceM9wurhmom+FuELDGL37l
sHTFV2lZBet4qU/JeygD/K2jxSb5Oi95rAqdvwio+mlUhSco8mmwuXATCzQ+Qdwe
FW7lDcE9fF/stwTCgOZA+nEI7bzEAKp0dEepxK0GILBSzFY/bHcQuXkrvHSMaDeV
JlF4aKS2UMsKHrtZYm+5/v8UymOmCStL0HKigGxSlJX/wJrPQkBZjTJ0LIC3w5Oc
OTd8LhQZqwIpWdlhEFQcBfvfBgJJvNPym2t4SbhAud7+iSFgQH7+hvcRDIeUAWWn
QBMfpgWcFPYBf/3JexOJkn+TifU/xJsuF8IGkwJhvMkFwEHVr8wGGuEezCQ1dBMk
kmjEhNx9tVkgtj9W0AGn4ghZZLbClbwRXXofUU+pk2Mo3rQRElKJLwiGJ278taov
I4M6EAfpVWVEyIbUUa1htgqospPy0qnUJnzsi61Qg8UYYXu/UbvGtkotWDAloGpc
z01p/fEemfbjlyzlwmKfCGBi4kXK4WaFwmeRWGmaS4Z5f5BJAX7e8LAXt1JKNhsT
Z/RA60Hy5y02HGw7Y6HCW1UsY3ywMG2K/nGqQFM6DGCCRhzbAgiufbHC9fTUhJaS
84txPcP/Qhdk209zRO6boIlPrNKRYNegU4RiIOqH1Om/WHhUwTxp5tqaaJvopGNN
cZdW4Vf1wVIsjiyNUjaGh3pAnUwKVcSULImG3VOEDoaPk+XWSCgi7YTvIkqVvQnc
UCccBmDGRItzYzeU4kz3ARAaMfRsweGazVyo1VYPj4rAVC8yYsAnDHflmfXmRgj1
EFLwpZP7MeHTC2ZD6YDA4NTrAmpWgkADZAd/rQbf6Aw47w8sFjj7pvXV31ibIz9J
OiKT9qhLPS79cAJPr1+oxKc182vHV1h7ZmDqVolOmHSy24ITUXj+kzcb0I+P1piQ
vax2mC9DX9RQPwa3gpuo4RCtmTjIc97D1ihwqW8/cfSDs13+FzKhTQabofU7xB8h
/t0J6pPKHye/KPWo28li0LYdoiu7cA+vMN+iII2W5hCvw1ahcJryF8vnaQr4RXv1
w0/eHsM6DqdIG/D4qbtefGVGcoAMTTcUhf0VVMvLa4vMV8HxO883eywYHEz3AaIF
uAmelGdOjbvIYB0ESfVbP0iQVMsj3AZ2O/xgu391/44d8lYBRVKCIyJvIg3xqo97
fanQAtS+5wairvk+uZVjRX5G6Tl3GQtbtMkE5Ota3inxMnOocddpdOG0jROlsfrl
g4nMQ2kRTGuWqngdI7gOMkkd+kXWPQz5hYRvd8X7cCRXh8CBentQk+yVzKRwCtWx
rXUDowMr5q1/0+SdGJ9FaVKKdBUAizD0YUyFEYRRnGVJKth+Sz2o5HefBcDldDKl
RE/EDrSLd5E2vb30AoI6KAItNFGaCGDshTqXoxKeMypPgjEp3RAtQRt1JTcGeH7u
fqoIyHhJU1PEVdLJqaVK6GKlsHqt6XmWFHszSSfHnmGt87ZjJLCmETUzDYWavpJi
CiLQEKZy5q7xcGojqvjNpl4j5CBYaTqYRvYRxRtUnRvfeWv6fOdxeNGT9SNedUBn
wjcgzlJCSZZMBRmu0VN7S9OB1an5hA0IZOlLZmYxW5wr3xZq3Qwkna+YT9tim4ra
S4+9yuVKaHaSjMRhAQrqcH6r6nmQxkIv4/HKHe4uGgoeqVX64K1TkRQUFypFst4s
qUAjdzjX6lQ5xuHdb7U2dQPQhUVLhAm9VUFFAtY44dQ9ChUNgRsa0QWS6l2TB/vL
vHbMmO9+F91kzTKXCCc+/YHb+U7Rg/qCs4JpaG2VVjSWhG9N7x/H2vyjVis++osc
sXz6fBd8x6y8UrymVEDGbGInMXMzu9ruichDnEaZoYsHR9zPjIdFaRiOEg6mO79e
B7KwqMdFdvINSidfk2cKCGDKYPexk8zyc+23pjDwUt5kcu3A3hZTLwk2g74dAI8p
96oiQbaS5Dl1ZFi7Bxu7GQOqH8YXeQ3jVlQtoYNEcTJjSLQ/C8WGN1E+oK+KfVuB
XDdo0q5oKWDYzNKlpvMWHwkxzBDewSGL+MYqTkLtZV8CreRCzuS6rq7pDRcc0AW7
yVqPceKRk+bvkkwaKexVipT2YGg7JvmDXtyG4zwxaDUJlWdJgNF185RG+dHfmE2R
rgBuXCjOZXb7WkmoWY75Y1IeAVDBeFP8HnULQ8xgVfyM3YWsbeIozq4oaT1Cscio
VtxilCggI6OZIrB9Ufbm4X+XtFZOP2oivWc8Q06+pfH2Fa681Ii1sCXTGFK1GPhO
94qfixwGOTOI5Bh1SjzA09Lq01rczdrQhDZ7cxmx7GpFTp5DSoxseznXHNI4vCWg
XDzvY1XvxXOaqwpTp76zKE7X8jDZgweSzVb2edMFTTOwmQdYsNGEHnU6soJU8on+
Ygfp+lIl97ZGdhVEBpLTVvFE05J62XDghPnYMC9dqmNs1N+ncsp84ZNJd8CU0IEi
RKM0VqLjfWMd++2FAwh5r3AgwgtywIig9lf/wPxy7BLCwJxOtf/OdkL7SjFNzN3b
S6lrs9hHW2h0XhEQFlHS+AdyWZIstY01lEnNDWAW/L+Li5xz4zY663T8Plqph4wY
0i7w7uQupXTzQMP3tbWliuFGYBIynquTWfVgCIjzFP5/nt9VZAag537ckn9Lfcpb
47fsyoL/HYjYIF9PhnxWXg33GkN2uvWBgiHQU00keaNFDdlIs+f5r84/3O76px2f
Mk/znfkV/yGp6/0y/HaaTuiAZSc17XyiZyuVkXur0ENEWUQtnfYfA3Rmn0Dz4dZI
bw7768KNaWf1U0xfAW+4srhWdXp5y4R2OoY0GOzCiAxXyv5G1AfdyRBub30b1WOr
mhXo7I6oG+q3Y7jQWPPSSW7vqeo+LwRHl5SGNZjgtP6DNNGCJ5neFvzlzofbGm7i
giyJ3f17ChsSmewW/IpgWTB5XBYQ/raknQklsDnXpxiMCujhX8oGE0LArQZbOc5J
+0xtbZq7g/S/4/7V1tZgJa9YvKY7BNUS6B5p+PCjorkI6SprQC39RtIYicZNu6qF
ObrMmU6FGAOUXvdc5MvssMfTWTp0X9L4G13THp2Uo3Clm31KgSxH89wE5FDTLhOV
dm15hImzg4e6pdKsNWF+xec4LIeWvTUzshRYlkgkg20hvwJfuRbFY0kxOD4f7Rrc
C0PqjknlkduzDPNXfs+CUH2H9z3IuxfQZjjw9qlIJrexQELtumj1I2V8V8sN9F9e
YP8rbshk5h++tMnbsA8wBfihKa73gureLCbcBMfLvrKzi5uLTE8Yw1sD6VawTd/2
qqdX4TpsSzprtzGQqp1rzr35sLzBXzPTlxcltR6Gp2e4R7Nl009gcq+3gKilk2XK
V0ULCCULx8Jc9gK8voVZl+d7zLe1ZtN5ch1DLAtUlDVnv8nypIvYWUg7UYrWdM47
ABp2xacxOBAFveZyUdfNKe8ucfyT7McgxEWYd58v71EbuEOCN2X1Og4iAIJ3a0ju
XCemtRBP2OeT72+YHZ+kLP0DW1Pbo9AjJTdkkjiW+wrov5AKEyN5qk4mCGIXfN84
3vMTXAxCLGNsXYrPnpQIKBYl4kVW4+AsAKnkr10ybj3xg2mhInjvfjPArVHZ3FhU
eoUSGm19U2mzNAAfgPAsXiNUtAndUymN4KshQK1axK9wg0fKFxNWibnALrwOCgCB
rpG0q61moyLYMamtNmcwCzvTjDKtTxXsbkOG9+gonn0zrGlt/SHrlVtnxXiw/rCz
xYYNrfHMq7k/cUTohbX7BOThEUh3Bf8symgFATOMIrEnlJo9Rw6SDyhc3DswQYB/
K3I4syEkSxMK4zg/1iNnRJQ0l/cL2665TMim6r31d5sfCXxkedTs2juzgNFeCOZ/
wuGjQK9X6P4UWhFPsn7O63KZ+xkwhQ4bEd0gVcMERqKdt1+QpYPKGIQSmoe6qNrx
i3JGx6qFd+oHxxMFpjYNj3FLn2J1PB3TVsb814WTVbJ8CbJN0BQFoe839Uz3fX6n
PqdRqQoaqvT5mdtCtZsbHluZ5720K4Yy0sDHAPZrbq9HqAfZsb/0BpKO5ucuSx9I
9U7nNXgLHlZOpiReca+zWreMtDGFFgw3JXoIag1DV9zv8bK3ChnL69NL5aNWRreF
D1sF1SwGUObNrOaJx26URf3++BztllQWuqULnDWDUhA63QSguFPPTOxSW+mjiRhc
J/3BbduB4W7mdICYVb1qiNkmKk4oqBw9OW3HK/PO900Ei5FYulbm7FCm5C9hKQ5k
DK1r9SXdj6is+7wVoxp9AIN4CfnjCBYm5q6oKjxuxehaekHU5aXet4oOFbfDW/bg
HK/fMBaYrnNY9SA+5zYW5TGI45SA9lgTQbqJrOWxA1JuM/egwwGHAEtiD0hd8ytw
x376js8kUPd3MJMYUhu/AMFvDFsBkL8OBYhRkA41I/L7hRLfg2zDNXMC1n4Z/g0k
/OGkxegm/+aTdBkDcWV7bB0oqsHRxdDZG7kzIWdr6WhRrCKnItwkrPgvTczKMaGX
vSgZklnbVwTdsUfvAG7ietf5KR18YWyusQ/pN3+uzhIvQ2bIMewRnn0Yq3XzeSQ8
wry6kO4iT6lQOfI3mAwC66YZ0XLjmtQ1BiEzKVAqmUFZ08A90frDWKpoVDZQwVQj
jRlQJak97QjH48twUnkXOSvn++LS3vBA6sM+BL6fhcHZ6GxqmpnNI6AsllkeJNRp
pTS7BpEWWOpSEQEBPl7+dT51JfB7IIp6Q2uOM0xoDLH1kj/YY2R8gQIKRPs9zVfu
XtluE03U/+/8aYfMopDIuxaIsuM1a998LwdWCJT1yHjZzWVqssue7g4XT1iHzQtG
7t5jtnpBnd4fLIURlFnwR7iiyvCo18L0y/jCJ+OCFT47IfaUoo1h0bn7BmMJ4d9A
vwFmT9j5boB32YBbL01WtSob9J/nE/46zNwfPLicFKMfFXui1V5/kS10A+pOKyV6
X3hTCVuZw9VEJR3CrqsXQkFY/GT+izzbiRn11wkBku3zzewoRc9uWuQMhjEm0IJZ
ijWM9ToLbchvOwSEcgxEdYPiFCrcXwCeBjx/XA7KTnKPg54Zjgm3FXrLf8+SAtTa
GNjEu+N5iCUmC/UQIt5kkGdl/5+eAWSYn7GIucGw2F5hOGLiI6yUukTj6qZ/wuIp
Pvme45m0lgBunASIaogjkAo6phPdjXPxUjM0sC+aRj4YER2Kf2krEu5TJ5HQLs0d
X5Urud4OCCd737KgOccjkkBI1FfYImy3i7BJFjmVIhjipqU+y9OHK9832gSO71nO
8FqiaX86DdyFxo9gBORCiULA/3DinthHstJbXOXYQzhnd97AVBL8yuNkZA+mdDZc
okd6BybDUnWCHfRCrtg6ObJELljTTPx35JbXe7S8kU66gYjTIEVa3yLp4RAowGSh
2uy3W2j9JUNyoJpqHWlAalRNmhjck2dntKPQ0FHP5tqeJ9qysIlNGgBFX+jqXczj
ULGnq1/zX+Zb2KEVz2MFpoeXv0yAMJwI0fJM4j9uJcNkpF/0pwMMfqI9IZKsgLZQ
Q90/eNpjtTrkJUIGccUJ+mCLcMfgHWaHbSf8cLv4u6QwMsDoztJEW1Rx9a2/PNCr
PmtPPXIKtTQbtRyfDtXpV2jg5I09bXAWjovNZxfl/iG35rMyJQuF1HHY83oAiNXo
U9HbK0ji7FecQkRgPSMW4H/A17Rivwe0hqvV6egoabHA8nZaKvR70R8W0bLOk12B
w0lwYwTlw3SPJ1XC16ad1kbamQAJtpfZ4hNVg6LIa8ZLf7vbR5GgU2mRCGsyJIot
/CSGD4E2b/3l6sEfJEo1GABTalx0UOcWhgJ+b9tzdJs8hcexfyYdTvxzg8La9mu6
d2iouKiYLMH6krykFrbwk0AXBqkLdY1VOnuGtlbgUDazjIJjavU6jCc9VoPwbh9o
4H6FhXd9f88UYYHdODjlfg8J+7+Mk+qKCpJHcYOK1tPBuekqq8DU9YJt1Ci7t/xT
bFJrJ/E9VLEwF8uTvR0rPwrMlyQJv5MEcTkK4ecmxosX+KBn5fvCXv4Bbg4nhNBW
ZGSYMpw9RZNwUxJfyogkayzOWwIQVCfdZ/ZbrYVwBbfdHi84+yEiMpd47l5quatV
wLvxHWSNsQQ+/szK4AJsopJ1qnjqfpiY09T623fhRHlU2iNjGTrN3U37RQRGMxls
MLz47Fks0qOmc2BbH6tGtpue731I+zNLMtYdvuonrJtRKYJR6Su76qMlL8rPDoPN
AXt7CSMzLJNnaIXor7UexpQLHFtHH6ZeXMXmQGzYnrQpSxK2Bv9Ko3xAqMzJ5ZJ3
u+tlRfqoX4PKuncOsvMiFsM7oXWTshBlgKMAi/2Mi9Rxgxs1PArZkGhNUBQWJWEf
q2GxdxZbFSPlM2Y4tjtRP5DrsM6mqbimyQV9XXe5tkXomVgl72i24gJHY1P96EDb
oAuuTsGf5lop6F8dn9GEKEnntClqICki42WD97vQOlZ15iqNLVC26m8xE58eEhwl
oi0Upty90Q/gYLbfdHzGaX4KTuG44iDT5vbsVSceY98AjjndKfe6xaCmvKLRkyzY
iHm085JFx9HsUDXiD2C0VBkK02pCL7R+IGTEcF6XIVBDXPd/mJB0tC/mlOsB6zH7
kQxpRe2fOtGk0Ek5T0VuUf6KOo0TdQJYHuzNI87ek1FP8vGdSpemMWszn09b+bD4
7lKz3lalR3DaEVKC9+DFJ7Pck8gTGI1jgUy96ncZKmDG0mXRs/KOil/zeIfRZbk3
ObjXiSKyT2i6H4LuCplxCaj3vDMWPE6reD6ZqGtejsdUBhwK9O3vJRwFSHPRIbnz
0S9k1qUstqF4YCGswJBeOvvBnvNLRzKC3yh9YPkRprMjYuC+cwfr/R+GG7Gf7mI/
YM0Zq9k4NcC+17oTZ9DZE81bykVtVEMaLbwJ2Mmz//p0TnawwW7lFZFWCLNDuuVw
WYxuP1KOLPpNhyWwSLnLh0zKvOfVogGU1eQug6HO9YhFUxUgavxx+GwdiddQ8UQf
Bt5FdvxEegTqrdn1dEfGMvFc9/OblFhzmyt0o0+wAh+jTooaddAKAoyP0GH65rVo
VdG2Wj3akWLVNNlcKusZUYv0mgPAna+Y5In+8oB6ojsMOTUU9tBCvRlqj3BWrVil
WkWe1XCK+aI7Gj2ARhp0YLJxvwBzFRFyNgcA13LcVrbHN2sycmqPTWq7xswclzAo
Lr3/lc2qHtxdxZNkXbrCxyD7JGG9hXUM5Nlkk/IA5tHnNidCdmvH5cX0T0ef0TQO
0KA+cc5zeBfkfpi7GvJwXBCzo6Q6zzWW6/BkergFB7oRLXjw0VZPoGTEYr6mavwM
+jstHZbsmSn7f9akrA4IgHiGZFj/B21KPy8nFS0kicqNa9OSuRUsRHQEa8KK0V6L
oIitf7RbXO+ITae42cSRvMlm/Rt6/v0qY0/48gWKT3wK6bxHzrYhqM5cOJN9N4iV
O9ODNdpvBDwVsOVGhN9Ygk0i2vbVlihfpLymSOBOyF3vAhGF+5u6WC6iaxnuoKuZ
OwM1Xifo5CUkHEgRtrKW43VYUL7/HJTXJ2iskQ+3PX8EAdu8r9scMBjyycWTdnED
7OBvBPHL8cfRHmPZstDPhEHzgwSDi0bKggCBD4kw/1Wgy+tPsucwc4vBanJzeQIk
XzryU+4i+6LtI4jUjicwTsyHn7RhOMbeMuL9NXR/ZFk18ev5QJDCDZVSmS4VNqya
SMOpAB9HhNzijLXUD6EWTPHlPsIRn5/J/fp7OVr0Xt7lpp3iiYtTUJG8k62eLc9L
2GPTFRHs03MUlLUJT/KFDfi1siX3i+VNhO2xpJn+cqmqg4PSVw3RFjb8xckoFwyZ
vUjVR3UVKLuDwyLtXGj0j14e4FQ39zuqMX82zgOxb0bXvpAcA6cSLwZdSCRElQXa
XVeIEqAjafRQtfrRvrPAs3TktO8Re3u3dy8p1NwYg8Uk5oC5v3pLpNrnHMQuM4D9
8QpXSfOWcV1yMOnFIlI7cWS8tP4y9MR9EeQOKEcHOkefN8yf9ainZn0+tzqgsXRu
2iAtWjVjpyERvFhDss6hoaegl6R01bnFQ/qefSp2J5eOCi597elj/j3MRkj/SLlL
asOjYJJ/YDcZujPWdI5OKxCC0Am8Xir/pqeftH9b62NVdI7iEFSinbCmPwqEk07m
/X0o90zIpHAuEVNUccXnG3CQjHRNbLbj5gJAFAwvWFHypyD+ObM3CbtuiA89G2St
HNJ6dCL3zuZUGLZapHZOXt1E/E0aIUoSuh+8OYDtzS/z9AId1OXP1CM8lYpb3Cde
178JPdOd513yTGym43KRxaboqCC545RqAz4bC5l/YhBxLyV4/zqL3bnD7YpY0+dz
UIWG3JZnAA9KFLJJg6dysC9KW0bIN7quX0nmiqoHIpUUr5q71ZIvjKA84ZPnL3l+
NULtyxNtEAuz5G7ITSMpVJjap0qeCLgIa4zHUN32N5oboEbV3q914it2DgnoLQd6
fzj2pmax7UeItXffAE9m8gVpaaFJRC34Uf21IRB+mhv3ZGyjepQtip0x8FXRmvYb
LapilMKjLXgJ8pND29tevNja/+ezkiohiD4QIRUbBrHHa9PKTLHYoZY7faiOOQq4
M6s0Va+CcjB8ldrzlVu/i4n8pFi86Lo5pIuNLFDTG8J0mbpoFHmoqN4+dkdVNZGn
ae2O/B6ES0XqoOu5K+AshAuBVHVcpBuBVknFqCyDaLByRXURdWV/zKqD19FknSCm
DG442ScUWUKzp+kGsH3YZu7Z7T00AQYtlazlzomm83edZmAVpYtXO9FOne5dIIbs
CVMlKWb3xA5qROP5jM5Lv91jJGP2uOoVBHz80liK9fjrohyNi8TZz99PwoZKkUNu
nAGNue3JAHWcnpc7wWVEgjDQTzJ7ImEvJU2pAffcNC+yT6OvOR4GzfnvlE0MoLnm
lZ5A2nLuaZ7cd0PFHgOmnx6blJZGRG8x+J3Vy/5SXlLqsPV/xxfrvDUMqTyiVzjm
gj2xxs73rAym3v0gdCyFO/niwJ8TSctaFLoLUYJQmFsF5IQtGZBiksrmhUM7t/+W
iK7n8aS3lUgC/zFR5Cl3AbEvBiEKhkbua56R+rM+BWzEIKXJ9ENK1VQiHFKvVGKq
LNXGpU3XoV/5QgpVsZIQS7bxAOqd9RAnJ96mycuO9ZsU7pNPCrACZW1C1AxXO0Aq
bLxCh34x6u/WCZOUpj8tTAAENzG35Kt+4+GmdTP0ERowY1BNNdrt8ogFae3YZA1u
PxBbSdea701y/baDVJHBMUMOiBzGDF66OHAsLZ4WdGjm64mmjqt2vtWfEe8p9pPx
5jSpLUOEo0RSFJP0lzKiUW8EhtBIFTaPJoEVU3woBQZK0Bzfo9BTqka+aFU/OfOE
mapVXbv24vWQA5v3sZ7Lh8IZVNJVv3K4V6O384Mxdi4rohkFSlHgU6Oa6SVUBWzi
erL41Zj+fXaio2tTPTJCIoI8SuMKK5qz8ogNIx9e7PhrguHGpOnhOOu1kZl4Lng1
zP5wNInrMupaQf1KRRHELtJ+9LA16TgkJ0QP/ff2u6Ntf4OOzUoBp4QkEAomq3Qr
RYNldtW1o3KCKRDeDEJNQLJNyFcqKo23K2aa2Eba+d14j2SU9L3X6yAyzG4j5VYT
gCQW3+nFyliQRqqYqjwF8v3wBw4UV3aSvrSUckRE4VOGf5GHT3dITkBLQPCUSwnv
0ljW+WXvYbmdXQjrG9ig2cMh4+roZSkJ685sJtpNsbwdKLIZCnuOt8g825LMe/a9
UZO0l+vM51RwNQKIHdGF0IOhzvpwsPull4Yx1V8jc0R+1xw3aqj7vPBFiVsgd2OY
/p2awzVgCX6ri+gFSStCln5FNABQgIDikQtd0GWQ3CL45MJpxooBRkKjXm7VrAPE
pWIjB8N6I48MN3/Syh4FFgAa8AMZz3m/sTrmfCf9YLTLvN9audfObCyx5h7jF3jl
nIH0/urt23qwhbv1+Za3yxN8TQbNK41lxmBbA3TjxwINZ80BEv+1DO+7ZStPKwsM
QwcCECP8hhwJvZyOS+TKzKapmSTdStZOsxKy0ntzhTOCAQu4xquanc7Pe30CfoMR
3e0LRqe0CNasefLt7LDl6ctbxRwkJJZz7xJRusCLk5Q4cuCNtc055s4bQmsXj6mb
NLxJH6b12SKj3NaDL5WoglzbkZNCgii7AlYs7pEDiQy4IwHdFfFqV+eiiinxgEnq
sQZYC6WVO+o9hI6kpe84xRr2fykVaIDGMEzNE8xq1QgD0KBGLVSa7HhsbwNCb5o6
jqOumjWCr/eB0T952kop5xS0nrZ5mv5Hunp5tWRm+ip66dcYnL4WAvuPVV/7xOyw
uDsxplrxp7UQV3Olx9UOiMHnJCe5rxwTPIDpFORb8S8Aig58CZ8PFhgjREVnBHQb
pU9NjxJtTzNcn54+hllJ3ASZpDmk4Y54ko7ImH4oztDl8zDdNiDC2bu1QgstbAQ8
IUWF2Gh9SHjHpuVJl20cQ8y080iPUsnCoPPkaQVCLuI+o66qT4Y1lNznSlajlgES
Pn2IjRrE6L02pdviNxxUXnCLmfI6pM0ML6C5KvLNtM4yQUzTaJvPF7TLu82pBwdc
qX/pOOzuQ/VNPSVu/Ft9VCBxqg0MWlfa60kX0Yvsg2kCKJPiF003qaJToJ270obs
E6xF/t4oLb08K1SExE4+JFluaa9733waf41XbQ/Em6siNmqQ176sNYh2Je1y7OrS
Yab7AJG5g74vPB2dVktp7wO4IkZqx4DpERV5MDEZQPg7zFNVT8in7MXYUBDPdaXw
oQpQ3j/QYg3cqnn7xbX6OZTg1HfWASqw78ytOwnVoEFtTIwCj/vBgrrJSvOMJ/hz
wf1fHlhbDpsXAcsAhZTsTsfyAXvVmAEzFVybLjtDHYROOIzwHwTiuHhVaorO/oYK
FKfwLwyY5f5R2fpAj+K6yhoD+3TotAOG2t7hbISJ7ngZQL1/sulE8r6/TB2xQQeO
QtCbgSvUfhZbMwz7kCRzIfWaW78lmvVgAeKRgGqxP3+0O8QE09O9/IZvH/w7eSnH
a8xbKBZLpQf4E5uzmawLTV3icMZocjRHvB2v7+AMwviFDoSHTDhf3PJADT57iIdN
rjP226m7OsisSd5eHZF+WL3Hfzubs3JeI/SIpwzRfOfYv5wtgy//BmJzkNpWxuKl
ubTJPhOFqZiaYFDB/U48KC8lLPZkaQWsJ5qprBf0I2u4qHLrkjwqeo0LsXA2OV1s
H8sIUKVLzplHmwxtBXXtDgZjrlYkJy4X79+ImxEfXrMPr82f0KBjg2P4MwKRSedO
pVHRi2+r50ctUa0Cy3HCB5efc9uTbekkH7rgcuGy+GUO1KqQHaVi8EeKq3AJAbcI
LQF6bxst35OdIHyltgWovEOQvkny2iRtzu70mm9dvgG84Cz/G/v2QQbxaHWHrRNB
Cu0y8WlmMlARWvrscPHO0TOghY1TnOjZBh/RsKekAjLle90uDu2V4QxzL6NxIkv/
3OVrJi4UtyNQj5uoqZCSu7fnC4wC8t2jkxekxhrmuzWftXzHZampt8LHHFwDuar8
Gq4x2svXiCgZN6/vS1KZEx5eSCxPaGtkj8dwmmPW7zk5fE2lHs1lLDVfrOatFM0M
O4w+phSM8+TUyTXP7LEZs75Is0t74c1u8iqGKlcUvuaKsvrHyNyTyErDRGKaQ68F
9Xs/fhztEJe9PXuo81zOCBL3ETqzvGljrai6kurbnAXT1gsKDDA/nwiIbL2acAVs
wgZdhsZ5tiH4fFLtt2JDe9kfZkxDdLoP1aPA3THIBYcMwYGEr0cX9EwGwvhFpewE
Z+IH5wb6NMrZviVHpgT29hE/kO/7N/uZfGEyX0xnubrBGqIn9nwapUPy5TUcIwXN
mS+Ioqx4NFLzYQs522f7f2XplfTecBLGBXd9RqGJ/kEVTwLMxZDAHCzRTkXvbwg4
sBXfkx6fP+JrtUvUsdIUNt/r7UCnnh9cSl1ku5kv1TG5AtavV2JsKByh9h6eh2lT
CWCBsJHSus9sddVLM2plYg4qVSt24VfCDsVqFbdKupHQZ7eQgxUB4axFGVGdMhEf
4z4RNMSjmS+2V/UtzmOO7tPe/GeMo3wTSHd9YeqELi3no+AYX5NEihbAkPEghrvR
mYXO4BpI2QWHm+5u/QdU0z1VpgZjiBYsKMRToDF4rA+C/39WrPgk6kIax2h/Qfb1
975TkK3uMP4lD7d3z/eQW0QRwM2dK+dZwJUDXsyDgM/1r7UAwdZiCM2yhSY/nCj3
lIAU9w66SYuYPACTkOVPfA==
>>>>>>> main
`protect end_protected