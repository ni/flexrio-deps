<<<<<<< HEAD:flexrio_deps/PkgInstructionFifo.vhd
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11040 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3b6eMZvf+eQ8z14wALfTJHs
q3E8aWgVMNpEXpVH8GIRPzD5NQ/qPB94fcGqRTdnakwbdkO0gJ+pS10OJPPz0Nxw
/LCTk1hHkMKhE/EfDGT66XyIg+cyVOGir9iJ89/Z7Uv+mXu1IF06ZtSNnsEGT5Pp
cj3ZXXGXHSI8kuU7laNol5TKcuvxEbPWi5tcq6ROJOgxffIDUUkPTczMDGNN4RJT
5PurWnCUNjXFuJntJob8FCbkQt2voChMbYQA9yxLgPge+Q8CsVbesdQMxt785StF
I/maLEfW+sqGszMa512zDV+rUHg3tDTMPOebp76GnRVZA3/tq4TXcGwwEJyibpi3
T9YgLsVjLNbrCZMgW9vIgFAf7C+VH7lKvTmqlR1ZZG8Oapk4MIzY2r5CkUoVbZIY
WbbtxiA+eejTZP01SPuZepclWsGVTrMpogMH0VN7OlKYzK7mNnRbFio31IRegRKq
OtsmoB8EiwcBlQrU1pM1i5SQ4GvWDGpZxjzf71ZWUvRzcYwGK/elo9IhGca/+6UI
BFR+UIyBXyye6+7/wUjt89B5n5Em/njKsZEgAwqMer9GkMhHLJgvNVcQiUCkg1Po
Kw2MWNFGC3M2lr4ZpIvSCq/cocbkaFLcD+36+gA2BgvAmXwdR47rlODD3IQDL0eg
1eDhcDBA5U7BP4Hzld/k/xS43/VkzLjxyOVJGrYIY2SELERbSaHRd1vCHyA0iUJl
GQzPoHLii/SXqCB90cDEYdUj+Px7l9YwgTKZscHeSP6qpGWF1ulDAh0v4j81Hi0F
idS+0fg5QSrhU9zQEKadmnMLFtmrFJtFsnmP2uD4JbCKPl53rVQi8usrDl3ZwQ9m
KbU4UBbI9Dqb4IH7vIA15R0ExWt+SP2KOIYpGutCxjr4zkR0hddkcDZ8e8s55F74
3y6gQHroD0IIw0vVMyUa3psgELVRDFgBs5d1LCwMmOvsuIg3cnmvMt8QKZ0qW3wr
/evAg6e5EnfsB+IvWcx2Nlax4auoPvIB1z4zwUVoYy2Pg592u95Zc6QXHw37ucn/
L4ij5O5RNNTp/all9BwQCqy4Z3u9Te0IJfyk76xx5iAo5a+V14ohOYLIk1MbYayH
Ngp3LwEUIMKv05B0mJ9eXqsRHGCTiZg+ayWhoV00IxxqNlxHWIf7R4/HrCGj4cXp
FySuxBnCMXNmZkZIZMrcagJsg+CNBwdYLNCzWwP4JVvpUsHmrEEUYDRwm72ICcRp
CAuv6Z5gEOMYgpzw+KJ1UCupXN84lnvP3AYWCWOXY0GwD6Sz9AHFuedN0AfxFzh9
FHGKicz7LKJFyBv2acbue0I7H6danyk2obmNrGtmfq4YNh2YGXdVNf9vCwrR3X+H
JGfjc0g1le1WWoxRoI2ybJfMeFZjwAZIa4CMyil2YNDTM1RY/lr9bbQ0IoJ/azWz
qC5NM7oTMzvtKL1/FbT0Eaxe0e6yz7FJMioKVy4kGd6fazCnkBjPiEQVlo5PG7gI
N+opoGYziQ5+lkySUmh7khpJg4thlcLOFwaa++iN2GaNrHpKqDcX7wNeApasg3C2
vW+qvRMUkyyKh76pK0TLgdrxgvJecs/h9AvOyshH8/2v0SChsMRkyRsu6Q5U3G0q
uyEhX58hvdtyqgg85/ydt99CMdVxREySbJYmkvpwg0QjuV3aI6yDKG9AsPy/nSd3
YsJDbLuIc0TXJIVgQHDAfS52X2OMGumAGO2vOQUGYSzoj2Sc4RS20GWFTShrDyFo
2FdE/1BZ08Fo95+YccPoQJraRBu/0jzC9MmgGWfdo5Ljql6k+syhPsrmJjeh6vYX
9Jw3t9Suvqex3RzGjCeW0PjTccyVlQCKbm5omDb+W8pmyeG0eF/bxkkK5b3zo7c9
cP4omWjuOyfU8mqLcy1e9OytytR6szqf1BlCtc5Fbmk3WQ5nRBY1DzONgMn0Lb5L
0JCLfkKTn3uLz/fpf0pdkuuERSo+/baPbS7SCpObkdoOmn8RqMQWqldr9Ywk5+H1
H77vkI2iNgCJQoJVWKTjyKLw6q/PZXYI9jtNt16zpWnib8GVyS9pCXe2H9YcX9gL
c7KUWwtPlAqZ1oHl+LDMsG3zC+q9gyjvp++0YbbDRER5vE9jSqfkYcOglG3AjkZ9
y1EWjlYmWwqDosLbPstKyjqFK5yTr5jEsWdQ51Natcq6MOBr2ht3dlaHqO4Gj6YL
RS/gwa7pvZnKDQ777/AKo/++Pre+HzLQutIQMCwSIsydBUomdFy7XbJ53rMs+sZP
Yn4JPXn37jIVSpUFfUS71MqCgFHAAUj67CeXfVqMEnYRweQmVrAjoQx4b7QuZuwp
o8LvPiCK3n9XbcO/uaLs1qBhwGRKvzmcNzFdEjK+y6PW/hvZU7vR0MV8uKL4Q23c
5WLBLq2mA5MzmTBPaeL/RM0jhHl/Tu2KNNfdISVYDVkyjBbUoslHtqlfmLEU6f56
NBPnxbB6IePolAREcSReL859RjvjS3ajb0fE0qWI6YP5oKZW9QHqtiIGkKSfFdKp
J/M58IvfOjQ4wGJuqLbNlQQ1Rw+WPlmwoR6Gkf4NKt6vnJQiKlcjP3ITiydd24tH
ztfSc3e0s08mEKaRG/o6l5gD2NJktRgX4Wce+MmG+4hvrcViFOmIUXlfDvo/u+OH
r7CXC2QJYzxL+rQ4/CTjSsWJuMM5RZa1mIQewzqEPGYCTt2MniqGGjaJ5YtJ0tV6
QZgv4whlYUO+H5evQVtJWSyC5X8308ue5sLvNaSZ19GjW5jp4vAcOpZFz5JdYh4+
ZT1sK4NYbNyQx5Du8d8FovTOaghU5t0+tDs3E4AJidhWitEEQMmrmPdc32TcYKfr
XP9MUXZa9BaYs4lE416kOu33zfUiYBnO7tJZsutULF5SWhR46x/KIbmqPGPInWmX
fzTfNs2tDzezANJWaYDVp14H2SdNF4cX7zXGMEPbbAUw/UqgD9+N6LUZtn7feVQh
26u1crA5soEUxYMKEcUrHAH8utPikEDXA7Z2oCNzdrSB4IMtAviFweEuQm2CdFzu
r7oyl86han7v1c2mzb+nQ9vX5t5t4loOcW3M7B2B5vRUp4xTPTp5g3kdUio+jaPf
x4PBLOOiO4/18T/C5fHUS6LX3Vj98EqcXaGzu/2/46wL1WcZV40iFzptmZ8WzipQ
xFosqWBJCfAihv19+xsUqttOJVTyGTmFJSk6/WkejgrRR/2/rIH7eiCp0FXBA6v5
ruUFuBythwFiKKUQy/17ZjCbRwQ024TaBLP69U+mC/iUBJfmys2ZQjZdF7qc6feS
XCMMEHkOfAdnEya59vZK26txJw5TCth7VQfMvM41craNicsEyzArhGj204GsqCE0
kxPIEVp3f6IlGEB5Q/afLno+fUNGsOPeivv5+oFT6psUMa7pJ4YExtt33cfascSu
GVSgIUXg6iLGHykq0xtkSuAaoMFQE9t8w/TKUhB/o2bLphD8DQjJxtsvRrktxTwJ
d3/HgsCwGgLrdSfqnuaIjpzh9k6vZN5PobO1V9T5L/mzkAogWKRVTrq1x4kHghy/
LpExCj8pfJrIbDX5yA8NA19Ml3GA0AWxEGx6Rv5Kmson9VW1kSQoFdrnG6/IpauN
SUEHDI2VBfbvMU/77FCDJzWcoZjzKnBvZpzW+SRAugyLfEixwQk6khfW6bLpx+Vv
hzkeQS4MdaGdqs2Qzu0TGzTmPCCtS8xYhsnBbtgIjXyKA9qwVj0/hIOKTwFJPRTk
jV6LZN/IcOrTjQxzpqDa6U/l7PNZE92qRLOa+vLczT4bZArsPVxcBDhnKJIkJeOD
1AOpSb5NYeHLiji7h9/yZ+EEgEtR+JsIwVtOlrwu8Dmv00csWc2I9J6uhT05+FRj
WaDmehWqm0IbcT17XRqfVsrOxoyGrrPam1r9zC+lnh0IF+/6n4d/v9yFW9jhs+Wn
tIbRIAF2b1jv2gfr/fQGxuFkpdKBAFC6G8B2u0cDP1gf2f1ktkXFF8jADI/7kQsk
a2aPVRKmphn4FUfRAG3hVwQdtCnSDePmy8Df+owSOfNLgXdFoBC2fHUYwQAh4NbD
AmsDE9J7jcfdhX696ra5RCVSBFiI8kk7w7IXlDZdPDpnKaAIAuUfFupVcqEQCP0S
dGg8+FczYPmKJ8/uBv51ukbKtsjtV570u60uoqtTrYcMwbBFFY9a3fUGw43oxisy
nUsfXbp85TMxWUXuL2dHe500bmxLEwyLVTzspYcFlVA/zrDS9UAb9bvmlBa+s7aQ
Wq0Ru7WCTfDXyztRTGjmAr1g16aps2FwDBV7uUftXzkirkanI8JZdXIDn51rphJc
kr+jaUK34Jc3iJ/3+Qykboh5RNXspfH+PZb0g5lzm+J1d1phxH9McxVSmBvs27iL
+8VA1evVDcK730GFNSTYA+mgiD6M+GWuK4pwhTFsCIurkyci/XZ45Ajcdgh506NS
SR9QZt4Za6iHgXd+RysGh9eMNkiUvOAhw5FgB9Y4Inty8vM8MRx+TYzZjv9mL8E5
5+ilKq7KHYTRBGIN10XRIbZFDJrlSPtN0kRitqK66k7C5vEy1t+7rrgJJI3IuXUG
NINYhf+cJjsJ4looni/mg0viW1M1LOUWPpe5MaFxcEktx42MNja/wzwF/WnqPcP3
rPKEG2mwD9mk/QRPvQD1xok6c49iUz1sn2/eoHVY02owOoErl8+QEWnyBIa9JPRY
R1F3rD2KsQnT/u+fBNvfxzQj/xBbzqVmV7AJIzv/aWt/y1oJQnF48wRp0yEzNHx0
EE4OYAbTj/JjttB5bcRq/0YcyIqDAkC6fLkYb/fu4UByoGD/4FDAR9Q4xBaxmHX/
frvmvfMootc4OnR2+jjyIzpheaYhMJxHNlOz2GnE2psgFNH5cxkUWb2iYNYaqKxJ
KCyiicjwfk0lO53VU53HEQBWAKcCKmbpZPzvWNPtI5TAxZ1oyXzL9LQErpJo42fE
2XsEjCo93DwEuQpcow8h6S9zcbOky7gdJGAeHi/FAkja7mmLCsVijkZzDPoP3jVT
68zuu5zH4aXTczBzzLKIHMsBA9hLoKKHwbvn5PRz51ua8vgo6Sop2iSUr6BaePue
nnafnmCpy53oVSKW+WV2hRZT4BT7KTH14Cr8QaloSbs4VvwfJrmW3abrmHor7YBF
EDYFxNHJUc27S4UEBxDz3IGsg0TrGjla8K+0ylxZnSCtkdqAIH+F3mnGnbyMr/uO
IS0upHPYfgMjHgrUGM8ig5+5DyDu9TCUewVMyLaaRVzF+sTcy5/UBVCRqqZlCeng
1TtmeAqcPk3biS8HVVoeazLgCFLgwzvttogm7J6wIWnRfQ6ugGbVH+VZtr/qCuhQ
0aj/Esy5YJOvOhl2TDxWKDWMdQhayizl1/0wQhVj4WW7qdcSXVmHkvYtbBZTLa2H
9zEjLkgRRn7187y9AT5LKtzvkQEXXq6DqSQiKWSuI4rS9VBXp4qjSQy468GH+g1K
q6GJYTohOyOiKAQJXHcaldbOj00WUUGfuWRHqrv0O+EaLXm3d2TwspsEndYa/VDb
ElePjQBDBWKY+eoboTIRw6q98GoOl/0l5GKF+VeJDNe+zM68hy2X6zl7OWXBF9UZ
40eK18CEO0NrAcwPqGp9CStIYna6zkOb+ReCwwkPnp4RUIffRSurdCOds09Ah0gJ
d08vuc/QrpR0r5Cs8zL/QYQcC/fyqs+Q0pqFyksOY6afIXvUqvJJQPgA1chkmLpN
FZSZRXA7E585GxC7W936t4TFn6Kz8zgfqri1BgBCinx2SOf3D2vFteoGJ+ST9hdb
y4moJFdoBexnVEPeyT94vkKpphZ4mXT9PELxxzZs3Onk3Mzm9S2fbLhNlR2ElzUg
nI960EWxkjP0V2PVqagm41r29roi6SGrqt+kPVFjyzsv3L/H26AAqJI9RpuzGP1X
MKuFWXpS9WTl3MSW1YKxguo18g66nZVbvoEz49zFfAImlOjXbnbtncdsnAOv9Vft
V8eP40Le9pOW3Sg0eaKXWC+VXqfLrC7JQ3CWjsCk6ir4bfgzV2g1RyXzZfBF0UBJ
6kCNfpKPQ0ZJumbkdAD+pwYDX+4p6EPVuybrHd2k7cQVBuAhkHnCoNZc53NJpmv8
VBn+jLKPF9eWgd473I8aqRinnI25oqiEe2U6qeA/p2wjmolNLnap69jBlRiC5fEA
JZWZfFmW+hJRTWJtmOWzw2VlIOCDepAXByra/PlQrVRFyht6D79BCrgn9hhgnl1u
Sjp1o3wUF+w1Ha+MLqgpFkytbZXlfGtuDSoUQndXTki10M55sUn6rwuJtmmwT1wF
Lc3jocu8xPcir/EeeBkCpWMgw5g/t+SNs3RyGodH8dX8EgSWNJO3p7zw03VMwwH1
3wzBHgBp5/OzCi2gSTHWItclV1+gGcnwSqiZq1pvTqLam9z4gokdsBYQ2+B8WD1i
GZRcOnFIS3VltuMqnGgD+biedwrt4NTZSsPVEJoqr26tXabUhOviSInpE1h2oi/h
LAra2urTlI45T2QfedngVXqDqG9TkaGQVeTorZoJx85Rh5CpNV8PJRO/iesRSEwZ
ddrvsFZMOvqdmu2slfFyn1kR4lNBBz7ANhDyPP4/fsPxaUjO08hMaZ/ta9ZLcH9B
gy6VCEv18icFTkmsbBdJEz7/Oq36dqVBT/LJHZZCO0FaBSqhjMwukb9XsrLPgnnw
T43gpEq76b7zDQqyl5uYUrEU6150U4hz5xr4PzfkiWYv10cebqRvTY5i6E6XHroK
W74Z91oG7RerZ67GjF0WN6rHVsTRzWLHl+4WU+ATsehIIuFvPa+xReo4TJBtoA7T
XxJekVZpLlmkp1fTwlimcmww3KQnuKFux5c0Px9uHO8jjTWM4q7EKgh8BTRFlCPV
nu0nBcd4dYQ5vf/T4DyuAo03hIz7238ui1lNeOSn2HlPqRqT4qkAUlSD64I1Zka7
8svpR8ZUIjY1wjfwYODj1jY1N+DNdFk5EngdmWg4/kmMgOE6HwD8ddFnaE6qcNCd
MEOiKzqGyE3HFD0lBiegZfTs2AbIToBxYtiNWAG2O2QeM8DHXCklTnMOeAI/eY2a
sEb+mwoFWex5t6z3AtAn/Dy/3fDztAS9WoSwoj8UIN4Ndvu4NvNApDw7uJUjN9NJ
fu1VAZE7P+Q6ddghFIgu4qGJV3LFnh465ulpeDa81sm9EJjdGTc5ofh+nwEsFxg6
zCBtCTmhcKyCoSxfvT2tU2BvYybYGJE0WvnRm4M676OfAPlS0xOPXmCj0qaxsfqH
yzbHySZK8fII4sD/R9oLwyztj1/cexFBMSTkIzqGrcHDf+HjPbyM817dr58TIexy
Pgd01X0hn7HUXM0nKG9Cj+EPcJ9sj1uTZ+tr8gMKBdu8J6PhlXcVmkuWAeBuJ8TS
cyqAWV/zkSpIGD4eZ+LPOBucrpMZdgWQkyu6p1hsD2mHFgaq35OGQ7i1c1t6HoRG
GlylBpkHxu5MMkWCje/RqjBs5cTL7KbVYehzn6VBJVEPsEW7spO/9EHWdg3+9JM6
8L/MKa4EAHXrmS2OjLA4VPpMV5usua2UiBfU0GalGUUsc28jHoF42d2Ja6gvT0Oq
aENO8tFkm6WD47ZUoUkEbOMwRbYEwgh591GmQJfoc55PHJSWc8UJrNZAzq5lZY8h
aLhJMukIUE1VSUGKtlv60sOOLsCD6sbq3UivgVhDqt1PJiKWsfBPIeTEXpKErW6s
jmYsTRC+rTcS6+JIytHCRxE3LzzvlwhBXKjDlXxiXGATxFNa2hvcC03ZRODH81tA
f8M1tAEWozeelnkaOVzYmPfdwUQl2AGXUuqYJofPeOWlRu/7xvQtdTJ1P21r5wjk
NCsB+474NSEYLq/70zO/dBOOCxIQow+H07dJCjhveQ7BBVTISDFbYtyopO7a75Y6
xAzErVsxduSxyjTffPjuIRdyO/KSxohggpjN40Sd5DPxSsH2MnPW0ZibvCwCs6MF
69CW3BckJYAT22r8+8r9bAHgV1ehBnv8MfDJibLhvRlQoo3SiQzXYM0PJkheS4ez
iBumyyV06AkmhF+4uzlkyZN/S453WO48K0xX1cZOanU+jq2jvonPIzaOgOrlInem
h70vvj16f9d2VGZOwXwnXtIKYAgKsfC0P2DJ8foCITPyYCXs4Qdk6u7/E6s7BoD6
68FE6Mzc6qB5p0ICTIk+UTUUah+lRJ0OW1UwJCQAWHSutMT2/HlRHHWxBa5a+0AC
zCh+c/xkexkysMxXALFdVbBKBpSTwUjkE9m1n6VqFhi3PjHBjXaav5kaA8oAbLmJ
VytBHkCbEa1dTMmFpe1f0Wx1pobKFRd7PcrzsH4TgFyrdSB651KTuKXMAP8A1AuV
zlDAO22Z+RRfkwf268ZmW23nue8D1FFzJtVj3008fKg4b+dpEp6JVoyyWitnFW7S
ihTv53oGML//xjVEVVCTBHPvOquHBjS0Wmsg0VKcwAnTUFaoD94nQfh7A6jgtEQ4
dA7ncff9hYyxnH+f8wrAVipz58QQl8D0dbEK39d3amNDE7BKF9FX0zgDK1fSEttn
bq4J+W1xBCPnH7tdY9NdBFCtkLr1T/9rnPvsGc6D06Tz+3ok+ag3vH05gWyEPFNC
QSCffydyATLG4kDVFUIfuB0zLtxROebTKnVgNFmjgufcEcK7j/Lw4OGmrXGLBY3r
jvP2SF3f0rKWVQAtsBRebXix4ohOp3tUL89Z4nsR7KueeaCtyOnXH2/CMeLhPkOB
wVNJrnuiW03tw/y8DxA3/NmUqCiqJs5OuFfGm7OxmgMRDC8nnzRal8pFw0NTVw2A
Y1adQo0xJbKC6+/N4hdetfRbwzLj/NeIgUhoFOeyIajGHFIfsveq9sgUAi9OlI8l
XEWfiMycegR8JNLgd1xTu1LEwq3LeKcgN7tom+5fghQc/bBtOlXHSfDpnIcWa1ex
qz+XANAzTWToi6SyNlmnpn4VF0hfkGBkKsKvaeUUANGOyhzXjqGLxzUpQKfTd7cM
kzXjw/PHcF+PNP3A7VgmHF6rUtTDrrL5X9OpMoUIdP315RkoiuN9f2BQ1or+J2Ms
Xi1fScgdp1I+KTYLpzxn+7Mrbquu3JepRIkYbVnLd4wU+Z8l1VHOATDxOjyYnBIz
50fl9zs4EH8Jp4xHCxTswLN3RB3+k7Nz9NdtG7bALC9s+74wgbhWCdXg7tmB+ixu
5YScXupQyGoSlKCY9+RLArMiHh+73M7+PZzH45L1XvUqpbOhZuE5Jn+U4/hPFByd
Nvv/U6OsazTlgJgpCT6asAwGJwFDxNn6Qx+8Jy8hqetNQgxUQgqTRgreCBuyxzgm
B5u0+NqWJ7wMQ0EoO9dITTQ+tzYz1W8StTYNMmUX7mHpoGYgWW74t41K4StF3hPX
OpRwW7BO7oydBjnpDOSBLih4es43pnNDKRHiOFptdn8SfQiVlx5c1fw39rpCSRhE
DcMo3k0bVnGjfIrCQCBZ7BXI9OIvzIrKO4//T2tJxX4/k88Yif3Bqq/kmaW2UPxy
t2vZqLy17x3KGp5GONMKXwuiMZMayGGX88LzB016PqONyXeSKOoujvOIC/NhG9RY
uKnz0/Z5GpH6bb0a0ss54HpO56hfC3NJrRQ2KmqbALUlzE3lR45i6i3vxK6Rr4fx
ZvL3//f+KOM+C7Je2Gv9Odt2cBAUEsYr44po2L73bH9PJ5NGICNDiA6uWARIkMpU
27bQAqk7W8E6pDVbX8ci0oYWOHwKiFVzZnyVVU1bqXPhK7ooiACLMbqFT4JKLL/p
cmJGjpxUCtplJ4cT0o1leSVhhfkFy+vwlQLj8Q0yvegtIz56ZceKaCL/UTsnqrmt
OKzz4TjRdcbNaWq3noceWVcesGWWg99ZKlCZpGeMrCM2p3CoMLjRoq5f5e0yADE1
HN9n22fYRghiHazsvRGRARpL+oQ9TXABBWIETWdeKGi669kcHfpjtosoVYKeHHXl
9IsPOb0mQtmkJsTMSKzJFuUNHRArr9XLfxmwt49+IBhCawh3AL55wpEVn6T38bYJ
IVzEo9AywUBiel0RJPiLFpPWB2EvNUBPaDwfmnvVBLAWiezGiYWE+WAybMuiVgNe
ECnRS8XvlA/ehFwreX6WXp5quAKUnLU/gWoDlhZ5v047pKw/smAVfda0vCUFTtSz
V01k+t3dIj4uLJfbnWNNBs1NlYJWl04oEz8iDhxVhMOHJEWnVl2jFH4PKid9CGgH
IsuNQ+S+ObK+quAEH9a8EH2jv+4APYOe8RJRW07SpWXFlqR76q7C+Lj8s1zHKR36
fykG9BB4S1XVsA9yiXfQSsKBwfCZLBdUfDCRV8kgfgquybNFzzB4dK9T7Y+Ayzp9
ovOk087FKpUprmyB68fYb+ZrcK/luDKTY7BAm9ZoKzwBx3kLNZwSzgmui97zmOpo
Le06IO0vkkFDKzs8K41BxAqWtestjSLT2h1vtAbcY24K2DlqCsV3qWupNUZ8GHUd
5oJbPf4q1oQ/sgBTLkaWu5KP9eQEY+7RBHcnMOypJFsJ3zBv/Th/miSXcchXViD5
waiM1AEYI4Y6mFm5gBI1OE3KQ/Az7tx1W2kogpFtYpug167nzB95t/Xe5ZqE4BoG
ItjWQdCwMj+5+uR407Mn8FW4HGWYLnyx0KBjAxTb0bOi16ldUJzJ6scs0B8mCA7x
V72dpxpD/lYfXMl9p2A+q+9Yak4IWthTAN986hhA3zR7BjlVMiiSEOgRSpiA7kqU
HTPQpMmZg9MJzBd0f7I6sDVjVtgR7eBbQUOItct7EmMxVftFZihrfVPFExw2+bVW
o7TP6vGhiW6zxM1ik//PTqjvMxTJj1FtlBR1ChaPsWpLil9nDYaPUvx10qn7qEyC
mpLIWNz4fKiei3lFS/tdkSpgVkmbR072AqkKhEYi5nnKMnHSlUkqrq7IemAz3302
2k7Y3SkBXtB3cihNcWqVHFrusWi6P3TSRQzBB6sEcPH1yhF4nGF1ixh1votR1yIr
4rxZNNoSm3vPvlZC1IZQdLbmVqtVps87Kz8yMs9hrD60fZTq5/SoRmfD+ZIhsb+R
nz2c6uEaShGYinY7eUxLoxqQbpF/ghtfaXf2RPHx1s5zbyHWGLgGWWK4avOBgelm
f3iWGO6ZSzgnh+nEcPS/bsVAOndzHOrgBLJE0hV6RvHR7mcIns9jOPDbxs2TrCxQ
6Aqqeaa5M+uO6Lfipg2FpOj50b/+opeG8fuMo6By41HoWTmUYpg1/kisFkXA9xYs
SgyZBaJu9qErijOClOds3NnBOnnsLId+45G6u2PS0ABeMG3hMbD3kGt3YV7xW6co
mtFbcla3Eislm1lYeXIlTwTBwyUbr5R5rpg2Lx1r8oJy7+hswrlVZ0ANlbr6X8l+
62y5QmQeBI4iSWJeiHQSkcUb5TQPO9jPSsROTJvBqetGEUoicMsjWQOjUWFX8214
bVNmFLr9yGC5r17AEt1MLXExxxxY99QWyvwiRlNjxfXuUAVN8pVJMFH2SYddR+R5
76u+Czws20PAkAjMtgSWCL+PWelJlz4NQRRDQfA5qYbM2bNLXo+WSjcEflZWGNCc
0gyYmyU2vbsyX6qbpdCsMHbHWayrDRcLkppKGXPLRGiATBs+bYdOPrLeFm/tcJQ6
gvVBlnRWyqqOLur/HiQzZY70tfm3O6EIAMDV/VBr2wbXWg6ms7uyFJRlOaZU7BE/
F7ng6RhxHTHMA/zYuaXM6g2LW7jg/srLS0yz1H6JfdoTPJiOfNmv1Fm/bIZMvRdO
9VG13BeozxsGC1Z8yu64lNlGJanxnT30T6SEZg61cHjNULbzbZ7ybLhXDRByKJ7z
dlpemTS/niCth1qzZW7jVRdaPP2umtfZtdRXKSap93r1f9rZCWLXWaVGn4W+LPhe
DH7Fs7KzcVhWlDeyXd/qM0FXbq8d6MnQoaIzALSer7WDkOHRHtwD+FLptgcOad+E
gq7mvqX5bPacaezInLL1vYjoP/kxxORUnKPIlNJhXmVJECd1tHCwXf121fa6q9un
8mdWJfEmuSAG8Dq4tImVK+yP50zM/PrGpo0amrb2VCvLEt5zxAWj4mefFTB/d5FM
ZEFFHVo6O5MANOAddp2sfCWQIND67YkwEINLskOKmX//jCRSxOfRWcg5jPyVajmi
U5iEnrW4inmkyZUysSQkSg4cHzlvbGzbJwjh4fsvlpKTUKVIcqzvwDdGGpnhpSeE
0igee4lF0BsQ4+3I8ThdrPZAMyEL1Wif+YggNPVkq1rjg7NqXIk6k63aw+RPr92w
um167g0JpaJgqKEevjbqRd/dvyA2Od3HmDbxC6F2/+2VPxJoXBPb/Wg5Hlt2J5ly
T+CHbtserjvax5MR6W/viqBKQj+BAUMtQSgTUwY5lE1KujuIjjRpgY82wa66DBRh
GabcvrJTpr+cVXLSvTsvijJWPQ5u7Y0JtJaHoCOBqaK0a8sFuqMICFHwAPDt+OlF
YWlWjzlPALeCbHFyq3daC/7hedXBqlD8pIxjCvSGdy70ik4QLm3IXzlSxTTalxoG
7fjgR+VRtuAWNcwJCDEm+2+2kiJsmjlABCUhUZhaCCWNCesNTCFIyLCTDMCqdhe8
+JgGwH/GhGhhHx2KKl+Pg38eKxcm32GA625pjeRdkuqgGkJsrVbeyB5IGkhRyv3m
kCcE0mFcIk5TsGLxoEKw9/csZhJPCpW2JidSB3e29nftLs7aRymbB9tJ0WSEJpBK
G0ftwSToFple9GYcWJ2+Ddmiff7GSW6PhuR+xEpZI9d3ytcV6bZDm8nRiWeCDqjH
BbibrMF32HpQArTVGqiQOZWB70oCVMPZmt5jTY2fAFRpBUMOY+XowSviOm+RM5X4
wks4LWYO4MDK8uQJ07IvMVwz451XkeGuVzhHR3q7B+6avKlaTLEylXSHOLxSCYlu
Sipbwtq023bUCTBKKEoZxDiYfpaaw7tJhmSVTgn8j5KdXH6Zw+NMJyiDyrwrrOJu
ywQwhIGgQ+uKbQvS5ZfRM50a2MtRp3fZxfohAGa0v5HkZANlD90FoLgHz3P712bh
cUc2PoWiMQHYKoLxjTTN8qxJwWwnxjuc1bu+4C+GX/PUVQSTLpThXBqcpAku+0AX
gWROlTudqBzMZTSUAL/jfeW8IWd32iSxWYtwg9V0RvjWBWQR+LJompNTpGyE9J6N
2elIz/dLLQ3P6+dU4KOAqWknSSav2VSeTE/MhFvDTo/v+TCXczTX+k11xhVpONtL
ESdpcOA14BARMlTYcW4gozHzlZcOtgkUpDc9qYpiwid9sym9kl0VF4OoE4mW3fpq
62orVj6jV7u3Q+iKVs2BsFePE2UHd0tpdkOIqqdhsYcC7YQ7lWsgJNKwyhzFaOPf
tj4/S203HFAxILCGc999ZBsA5PtdCE5y68aIWDlVQ0p9Ens7aeJhQGiVBJNfuIvO
0nf7laSXHb2e6arJqieZ2P8CtFu3dn9FxdiPej6x9Cu9OstPmfVcZSW2UgrjTL0Y
cqxq3Se25si0mdFbXWu+npT6O0Ezh+tK4+ssY4dGNLCJWP1Rru3H4ijzU6ikHWRF
Krpwymsn4skB8mPpAtMJiayTbLQOa/ZOX7InANadHYBZYyg6EjSvpz8QYpXCoPQq
7n2bmTFw9g98kTTGzYCq4bif8Vho6qg+sL5LjIPLauh/sU2Ic04+v9lIJ92EpM7L
r8iqlc1SjQtRm+v4/P0Vc8frN+eoFDOkpHZI5+FMY8FuweYrzGoRFwiYtFEg8cKA
nGauU0H4jXzTi3SoN/S1pIc0D1z5Kb1rfLVIvojKVstPNbT8JUgDhL4riGvaLhbh
5oJNkoVfn1wnVyw0MVW5nEoEPKaIZC6RpWLK6X7nxU5OAFhonvUPhLX1qCxW8r7n
5BW7/lS8nw3Ij6M5lpIdFe9PYZSw8VtYaP7hyjwe62EyjLzX1u7Y8p7oRVXYHeSq
VmXQ0qCtKVGphVSZQCi4FStvA0EbJZqarxwbtehKoJZqTLeqVe3FMBTz4/6mH++r
S4iYEp28ubInYv+pgad2MquPZrUMAmLpEnUhDpe5O/Oyhk4iBeR1v8UxJD1uK/Om
2X5uVzFgkYJw2oet4szdOBQBHx26RK7VDo93+MCirjrBtGElx/cr5cDMGxpT/FVk
W1Zs+3Fe8FeclXRqw1COxo3XqxP0xRjzRHdbRx5R2PhdNi8FCEsWHD/jJkH9166d
1txhgGAcbkKolJ8SFxHPOBVn3H1Enbx6YASRQ0u9W+YxZMzcnywI9Y61gq37ncaU
GysVq9zF7hx5KN1E0Qr/J7s/5RKoZlk9epVpbpS5ddwnZrCkI2u8ssuRR8Gty29I
hM3NuLti6Y2HiIw5fidOzbH8Kn193yW9FYCkm9wGJ7VE04PWjyXBluo4XXk7Ai6X
ttbk4XxuVHtIgIKHcMA82tNqtY31S1UpLecRdsWTtGguWMrSvwnuCEpj8Frc6Tsx
SyrIUhrPXCGFXnnNgGGH0pfP07pCVPVmgYRQJ2zWk+of8BzEEL5cjJ9LluxaNaFA
Tr5Rho9hhaPkwzMytEg6wZrfUUHogX8cpI9bKGL3pzIRfg7piI/LoR8xADzZp/ox
suNf++TIMr3O3HrKflsassdeO6vDFHwW/T5dfwt6AvW7I6aSFpLRhMNwL3maHMJY
=======
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11040 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JXz1+zHgF4n2s6TEZD4KtuQ
ATkS0e5WlIVeyjNZ91Ns34mGmqHu6EGvs4XJ/VDUJsWW69tZddn/e5K+z4bIHCK3
HzrIiflk9Ike0DA9KOusgAhjZJq8D/qpUOTPkoiCr4r7ZnLr+Y9Wq3GmvYmapi2+
AdoSdOniOYAhJKaaSftqEuykMH/cCJDqJO72+r/7it9LPOIXlrPGEMoJtsMsBNur
/NVWHM75ZLcMLCNJq+Fh7GFhc4PFud35I9/ST5fJinlvpDNOecjbSXd3HtD+4ocC
3l5TaMmz1qKkVgb5Sa2EHWsLqDTyiPzAcvKgiPetVMr7jxwZ3hG92P1ceY1RSR1m
I8C0wgBders8kRcpL4JxyxBg99jh6BilHereIGtymyS2s2p0AhvD8t/hQ+GlKGyt
mqe3k7h4ww3nZ0FcRf7GLNUPvLdbsZQvyYP5/R2hOuB/4dcr6Jszs9ezBr+1x34B
Tvsghm8hT5Qy8JNH2EsF/wjzhskxqvq0zgjEVVng7swk1v+Buf5ow2HZ8ymwYvlN
npHkHHokpt6K65Fs0FqJZxZhZ5kOHa9ezH4LXGtn/1wwfQqmcILZuwR2VtS1pazV
u4Ah3NWT+RZ4OMODpB8ylkxuw2BU0N6GNsh1cs4N3ud/0kJjqnNuF4LigSP3Jef7
zF/xsdWa0K41NNf48rm7QI10HbR7yWP5iPeSEnS2wJcTxqPoqZrfbfl3BLGqA7TG
ToVexN7kv5MJqA/YETpCbQlsZgcinl/6erRlAf2ziitCmPp9qyDfdPBmvgvV3ySH
jySeBIOISLbQBn/UKrwLbOBtpKpUUaVPvMVVKE7QQnjT1EEnEfWgv4tCnGbIDHNG
jJAitq9fcX4jSz0WMSbViiSg6eWwrhrMX1nsMlYhIOT78czYlG2z4Z3yuKn906Ex
3tkgasPxsx24x5jinHvNqCsMVR81UuVtSDPme59BVi6A5XJ7PkVVRko2/wOnw4Lg
03PZBgx9359EVK2hke0QLyvl25Lahp6ih+CyP7EcDQm5BIDLK0wrZ6hwJq5iytPG
08LXE9wez3ImvcopehMSxjmmq6iIghHpths25L5ueUIw5L4qcHv5SWBhoMUaSBg/
YiePdyAyGkDXZbPUZClt95T9jJiSjKrJKdCTINgAabI/a2648vKO5HXASUFcs1yl
6PCRgf8AIQJ5paVKFvrFMJRKc5vzL7i9vIKpqvd9GRBJ56Gdl7dFTfkh00uzR1hY
DvB3eDOLlnLvKse0D+yIBQfi7BfWX/gkDlsy4VfqJvJjYJi4Vog+SYvHntCOxYWD
FmCIInKuKLie9YHyRWw5KhPlBScclbJqXd1u/IGJlp7KDP7+HXvXcFSOSMU8R1l0
pjUiP+3WsJhYdbqqKHJfcppnb7P8F6I84MAKK8T5sb7jKt266rpxXg+Arw0ZGNy5
osVA1I3L5NIqjPPTKfEYqGfm5i4OOAT+ZhEbc2b18SmNJ/Gj4qS/kkNoGCrNGbs/
s1Dqcnd5qKbXi9QhlzFtvw9y67tRPX66kMC9mBe7/8cJk0pDozAsRejHZveIgux9
3IUxw7Z084D6PuSaUpWjK8P8yQ+EpBYoYS2yhOHHavf8jc29yZzwlsVwfkb3LOb5
b+p1PU6s2UWVo77D/nl3tTCoT7ByEaHkASMVnP3Qtk5ghU7adei4BGyRMD+LPeJe
OTeE85QIuBAXOT3oKpqrW+lwjsfVRPHX4Zs+ZOoaKaG0e3szX8jPrTItwG/n+XgZ
RtbTA+jvvsuHj1pTRszYkTE0brOkbsnSiLte3KtrpXjNPqTyPqZ+avyAHil7b2a3
gVuZMZk5Q2PfLETdFQMRHwjgV9U9vQAYRwXqskj5xLsP/LlgtAywpdM/s9EQsjLE
VUYl6PTCIB+cbITgSrrXRNnfkYYBjaWYgxHCKYEl6DuVV2O/Y/vhSBxq8p3DTZ/y
2vdc2GwC+z3CKnLiwTkHmCmiQtbc5jyzWmFk5Y+uEIYF9bLUwgXmeyrqOYg1yDrT
ZKdLFp2aGEkQHQ+rWG6QqQMJfgKxfZD/B6hWDsmZAzpSiZ3cvu5ADFMADsDlu3XM
KDUdOh7FDveEyJt58aCnwi13Pj9vPErVDyVoshaAkfcbcHbe3R+4iI9QBMCIuNpG
UP4lJI4d3157NpjBNhpLELaZ9GJoTRIHbtuThaYXk+dzDv0XActclaaAH1FvvBpB
4eK17YvHKX1TXAMd+jWZJFvqYAfauSN0WmS4ukRCeKMwPwx1xxMVYnb1LOZM9TT/
CdmhBKxLlSw2TmJfEUwOsnKQxS6oiGRCHQCHbvwezRGfVy5uRDVZNrXgyxtmdAdk
KGBPKRfN8crq5eJCvTd5SylwemCpWji6oXAz/SBj2bxz3vcZoZFD4IbUnhtlFcbB
4ZmFWAqe3hq46m8XO9YiGmBV8i3gnzYOcqGMMtfU2UQyEMovNA1hW7Yb7eIlrJv7
3K8H6+1c5i6gkfUnNPNVTdTZbfPiKLqB2NrhT4vRVZF3eT3fjux1Or4oCuQhfXGR
eYWYYiVZLTLNXz2BQi/6sWiPHitEWdTMP43vHRg9AR8++3TC+AWNvejGkH/PCyw/
GZrBqaOYpcezT5RDIEVwWJIzofLsi+ivf/AvWE1JdLhlR97ziEn5QPyK0jezl1zA
3yn/6MfnjNrrwOesMZejRYG/z27EN/3PjR5TaO7VzWx1x/kCHQf7lOA8iQr79Him
kmO0aVPCFD/ViYvxUJ//3UfzBzSZrtnvBJJQKH38gF/pDOTmKuOaPaD1Zpi+BVpe
88bflSY8rIQBxKbgnNEZzpZFaD/EYdVbynHNiHJB5YVeb9ZJsqkQ6Xjj5Qqj9ih0
tGa/YDiIprLgs/tKzB2WL9BvOKp73CUw+6/rGI/JqDqS2zaPkPRFW2Zv95g5uBU8
XAueJum4j+J5BRpA3BeraOo+AjowvPMzya9iCTPEss72AFZE97E73kvRxhXFWEtj
XM1u8YRjuqMbhUVWE+htZThWdhqw4ZG/IvFciR0DIIR2dpeDEP9pWTsDy+rWEzd3
UgtypH7DrH3gGKqgJjcOta9ohu9rdV0OvoFI0F+BDL2/2gOI1P+nvhOQaiunpX8w
O7+vHGAN4XVwYbZO7TWTIezw9WwxIqs9d/swub2qw61PfAzxFW8T12PEBEoN/Kb+
Nuvuo1gXUeeUDjaIoXhu4GvnkhMI5avEQa7+SRcMV4AxXMiHgnCMN99U3jXjiai+
KbqKCnctSf5Me/lejb4TkE9MC6pLPc+iktySS4/xy/P9av7zo83M8hOpJMxIFAwC
hJRYG5FZy/us+eNghUWldj8YUepR4kRraR/CIiHfRF2Wy81JiqbJNUYQH0tN0iut
iTP72C7S+vxrsTiaS+ZzleXzvjqnR8vhUkF4yU3zWYsyNzajePT81KEXs6OLZ4fF
3VBRJC15eS/K7i8KGDJiGWTBSwXZ/5JOhbeCJ/7fLYou3RJo9FQ+/7/g4zycnI+2
yjRupsfYSka2R00ioJgEtzydUrRs3Urn5vBSo4M65ajihDL+BTlwO3fO2fODd6q6
CPDYDPs18YVoDVncrgomXsz3jjziBPZ/ACfY1JEN4hqIK02FSLgA8CWFdlsNfjcL
jOYFTa7n8vQVkJD0hixx1jTqTeEcdna6uEKRONQ4j+xYa9OJQZYMpfsDs7rd3HJ1
t2Mhu1/VV5r0Pwjfarhd6EX2N+5GLT2vrkl1zkmXNkplL16+34rEh6e8gcQvBb2L
M6nSQwp9YDqayA13bE+TkGb3E6W5blzuwQKnWmCZUruPYdCegQVPlcLZqI1okymL
HZUPpz5fsBYNQEX4iN2+3mj7hDqO+kkCu9cTf0oKqsxI3bzBR9kwsNSd0bGY8B9k
utP53zYRCUwYVOVphOMN5jgR/xEqsKlFbTazlAgsy9HZ1//F82mi9R1+GodufzP4
q23wLkQhVez4p05c1yM/gnjy/Y00DcBgUNwQ6DHgDNGxg7s7ib+F3qec4Q8Nf60c
nlH4MgKqxVvKuYMTs+tknDWO7RLe45t/Wabef6X5o55i3tId3SDt2AWhk2OVJcDz
ScosTJxsw7awkBhCZ+0FhaVZPF0AMcn+GMw3tcVl3aVosUy6rxLWD2ZmO94AqPW7
UejGaXRlRCSpWJVjYiihvZyz40IHmZ9q86NWUKdmKuVjfn24p2z/mxdOu5vVUNwA
vq7L11Fi7VZq8KKSeTu1nA88r9Zi+nkgUSzye8tpuAeHMXBuQl8qyYTVyTkBYDqi
kNhvuzVPnOvyhM9XYaK7yXQ+n/n+BJChfy0S1CJlZJURtqPwPsc1pBUBw+8fAROE
+epM43SPC3UCo5qKzoev4C7UnvqoXskbDsuU3VDKX/XkY8CuXihIqntdSjlZTxqQ
njG9EwJsyYx/Ks68FqE3PEcAlPi5SqhtFTawroRODxuGrY5VsmQ6KbixinXjuNGC
6wTZ3V89Lnt0X22gnG+Qx8FZ/vVGZ6bzD7hrOFpxdPXTZvlh/dpYS/aRRt8T+6yd
rCbEZNU+uvWS/sk7eoo6ACyBMnTL+/OJpO8df32Wrn1mzCe9QxTteddTyR8cVDXb
6zdUSuEhee8bSZOu0jET6ovdrV6tp7vkCitE8g5dwxeFylZk4gMvYUlAgpXiRjrx
hV0XCTRh6tkzagPT2kcsK/NoC/4TlWSAaCY5rYVbKwmKQ/hiKYhtudbhErx42B2Z
jA7IqsKGjcxl6aTjVwN0Hp9cQZ+lHw6Zxokumvj7Aq+5tTEZk1bTh/U7h4bWHVgi
fLNBx792VSD8SCoCk+x+7CNhodESypMT/Pl9eabshAsF3/9WUQsNLkqp7ZiRXgMB
MadxB+zqYgVapxTFECTDj4nH0IviQW16To6uEjmsrp72AYsTvp0tvkzZSIffRhES
xrzkS4MeN7nOfPABAlvND9FQQz8zEKx12/5exxujDFOFuPA0193LWkaN8hvpm7fq
WTRJDt45NnTWmSeHziph4jbJk1NiMZoDAzCM3ATPUsQk4CvVUdackZxDOUVLLNfe
LD9XdLfucpUIZ0rSHNsQvqU4s4Kz48hnlVjy8hbcf2dm0zA4euVxRPXEu/Dmfsn7
9w5Y3jWxtRHm2JdYRqPDtpkm7sofUVEc2g0lM+RL0LcFkLuKOA2CJp+rCdLKBgz5
pyAOF168xptYXOuKHvT8S5Xhs9O6ZioBMsATqMDTawmSkhpT+aSiQwMHvfpz7Mm6
T8Ps998fpEp8R8DS0ycREBb9c4RldbB2CawML2AG6EBGjsBwT8/UDoxSp7nJDGVR
4121CLLeDo7ZVMPjNuCrkddczihFvjwNWclgQc/HeL7C7IBulKII/ny/PuWyjzrc
pxk3vJD33HdSqb1ItEEE2ik0GQzs2Y8hE4CjCbQz9BoS+Tw/w9L5Jvc23HoC6IuX
LoIvRubDPqOxf7e2QGAgrTh4m6CuI962pt7Nbp3F1lgf7ZfUBv+yRV+LxX9kBk4w
3xQ1+jC3aq2Wq/co0btx/x8dBjiFNrj9TY6+IwGAjIrcDhdwkbg1Qi1RHWGTLXVn
L4X2vmSwZlaHH6DQmhnpf3mM2PoOC3QwrAXdid19Tb0KQ0DM2SYkxLhMUM+NoOZv
U1TQpP4/iXerrBny8Cg0/4WdCjm9kMact+uLuO8493GDtni2etEAXwZih43cJiiw
P/m+GjvH8sG3dAMjwvrJd/shQcDafEwdDcZdEstLkL+sKx2v4XrytSxw4OMJZs4J
OVGr/fQFB/DAq227JtlKjvNUrz/GLBH2SpZVq0gAmk0qhMu+X28yLj4ykpPCpM5l
xQZ3xqQrsONllgUbdkwp1cXfpn9YeJV0b6vOxAwR21W5lCOGQ/6Zwotlelqo/KTU
6BYXDp/W9zA0J6VeAczDrBziz77tT0wDHn8GHnMW+r0QNIZTMUjejeLCzW4UtFiE
35T4P9QPgF1ihRpSLR2n7922JYNDw9orfoNETMMlHedCp82qYXizP/eksNoWAmuY
FA3nxhgMz2HRWHssWDX/oa1uJ8fg7O0Mg1Pyh8xcjicXaXuNuYkfXBT5Csv8ZZQt
R3FJwg0uy8zKHU7ixd6z/OwJZrMRKpjVXwYgvOnGBO6eN9SRqDRjK1wyffYM4IIi
TKfv8k6SfmX6ABqvilTWDbCmpA7dXGdUT+j7oK7xnAtqqvU7kSRn0oRAqJ5BGkVk
pfbxGmp4y+n8i+XrPRWW+XhfRbwvmLGu63DuVtRvilgRdlQf6jnLnPfHnWWoKRCg
e60AEgPtsmrxay/5kuLiBpwuetO0yV1Doz4dEcvSeq6omcM/hHyOauwS5hagiu9p
RSDOwo/RhvBoV4wjFnbVTzI7WmqIiC/uph7I1iTmWT+jX/0gdrRDsJtTFupFp82h
jM5/5A6DK5FexNIqSuwMhPps9wkgTp8plM81tWq3UHjZm2bwCoZCkfwOfUn6DtoX
F/a86wmpY9FMT9OBVXJt0B/z5zXwHybI6gS8/8dF0MTimXVOFyeSsopefK8eUEtu
6VCwxcppdI49DQmXb4NuRdhlQ9GnmYAagPmNG2I5MYNBLbprM11eqHuJbj8KVfia
U3RovdkUgsq8FbIYjfIh1MchCNNIHZYdnUSnFbH15fiyIr63FXReJdt+pEZETBXz
JsXi/VKmemNH8/hpwjzwJuG0V2SsYRU+ChJJmAElU2zNlqP7RDvHegUr3maG3PpC
/k6vO8ZPGnLu7SqFSw0vwhnhsiX+HLtRXVisk7Ejv9rY/EDBd5628LW2gk04zTCW
Xq6Bj4Jav4o041VYfICz+nqWIYBDNL4fwH1BuwByI+dGwgBDcMbxF0MDzSQCT0tV
k9Ew+dpG694/Y2PTXz+BFr50Kp+gaF2fQ8tgfTqBKTUUAZaCgSFX6Muig+kx33dM
pWdGjoyYMzSSkffNsjko0kNasyYimLk4dyUOnWEtQREkRcI5rdJkufGnpiLGDAVJ
Lx5EgUSGyNl5mBVxhyS27g2u57K7iotDecMLggTr7QfXLNiS5yOyelScP3Jeg2UR
KJWakYqhirAHAFT2EslvsamfiXDVXuLqDiCa8Bspvo+XNK4Yxofl4Nq5Pn46KBPI
lxqTxZgnLoqdRMAZHlrPNOXSsb+zXcN5TcRu/5fAFgAaOugToxUYtVAOHb9KdGt2
Yo0VfZ5BhzwuLNcUtSmOVfWpzROgfE31Pf2xakk2K9q2D2xmCus0UeWy/hQNAjh9
S+L27YRXamUdchQ+nqQHiLMAKlLNudTi4DOAzKMgAHIMsvZ7xN4rXChEZceb+pPy
7fxicL/rKC3kUoddsTfA6lQa9WsEFasoWujTSyFqhofn2/EuDN9t2xQPmJ1I0l79
uZ1JnjbwY9gGIu5x0U9ESFUsu/FXCsxKst83Kd0JYyOLQumgFOoq8XeuiNpj1ZcW
amHHpA9RKODZGiHDhYIris0xi0MjPQOQwHlVW6tVYIdf8BiepMCU697vHeWHXzvE
V0zWP1eNKtbSKsOpu9nNKU21q49ENc9eN7FBi/jRHzpI7taceSNkkqzhh5ZFUvKr
679GIhSATbZUUbwLXEPZOaZZSOlc8YtHIgok4Qh8UaWbInWUfHyDuCABlHz5FqT1
ISR6zoao5qPJ/A2uHg6ht9kygR8kucMnJ3Q6vPwirVXQt73q7QV/MY7gK6Q1UAyk
CzfSry0OK+U83IrquOch5f5x3KVoNLXxFci/5zyu6YesMPMsiB16hy4EGkRHTNUq
M+PmCoakB9UztMIZRvx5mrXwQrJf2g2+7qTKfWFykx1PfCywfzVPfYR6DEdpzAnl
N8hZtupSvtj01Po/2l/kHWk4o7+KpjPOcU/rYC/fR2TMZfuBI1UAl1WkjWHb+z99
GmdvXYytIxQtGJh/fAhiygxrwFuAel8dlWVlvkCjNkTHq0fVdrpkbNAZG9csa0uI
qFryaaskKXXQaFV9BRKvGeWYdve0sU9gylfS/Ux2c8p9zBqpceFPqvg217kUBSFk
MwcQhsSyrEgMe71GplAuqx5Z0Mwfw2naB3xjzAnSt336c8dvs5DfakiUKFAvhQy4
He9JfrlN1My/W73muywLe34caUcXH/mLrtX+P5kkVgGp87jW7H5GbYtW7HrhTubn
/h+ECbkHN7Slncy0ciLYooJ+J+LZSopu90bHFyFtcOAwS7gznMKfsLgNCuI1iWVP
bRzPXGjsi3k5Tc/c6tESFZKi41lTCCnDpFIWRWtctCkYKRIHnEUuriZxxc5Q06iX
XUNIaUKBGENVgum+3ivxQsNIyDeiiwSs76Yddu5Oy2TCTvDTxVdaAiDcAuA0NycW
lsTFXtiXDdxnpjJvaB75aPDk9rvQTMHVDt3jtmbU43ELpS3vWnI796BCFILxAh0+
snTK6pIvwymtuC1rR9JQcJ2zpiGVMfgCrnJtOKNHJc30OzxB4HjLLlg4LTYy4aBW
8pnnMBpi9rn8NUMkIF7vmmJrBZ2K+RwPrspuP3Ok0aVmD/DqRic7TAFqJOwB8rpi
1YaQuxwnaNizKM9j+iIzVJyH7CITtYIdtv7MUsco4GLDh1Z200VgxSIY0YeMe2eS
jye2ZsLQzBz2WjFpAC/kCQ4QqhK9glsIjokQaSCuml7koiJxL1wKiVevBvIqernR
ale4DjY2MsMiRxASDJsjOdb33QC6f/V4A1+EsTl+sbLHJPPHGV6C86/0ZiXRw983
OjYDe7Vp3IsPyPbBlg0q22G7rTj1cuKjs/whqNY2fwACiZfDwNuQWxK1Xpku5fvf
jn0i0uXreSIctU5cxSLh7VnBMWdjGqnz1IQ5AzjPURA1RyXg+OiFxghS/AWdT/33
1UcqETnUF5x96mPedd7icV9mHs4reo+50gkWkly/5Z8VxCtfrklgChkzawOHFAKh
5+wTv+aTskq6guBveLOXuV9TT9rd9PEMQd4u9pU0pJhkPpyKJu4juwQgL5V0rezB
Chf9MWmCPYcqV4/AH7WLRrTzXJEZTItgTPd+alBeS3EaqIgQjQwXxoxr/gGctvxL
TVph8sPkkmn4vitdbb0ujs9wp5MvQny5HsLQPTBs1McMPcLshWxQmSnCKtrp9TYP
5Fz6qeI6pi9m9EHmJ3obvRBGUEgjB11TlpPWnz3ut9HU5jMTH8KOc2WwRVlAbVTl
EVZBMthJK8Hn6b58Mfo7HPun5KDwdE7vUixrVGowHtJnxOlNBLLmsAtJCoj6UcyG
/2o1KPjGAegY5gCZgVVOjXx0OphSXbWGMBx6GwAPde6iEDBVAw+gb/j9i1PhSRVI
3d3xm3emVDotCuWPDv3qXI8c5QaFHEWwKbAub27KjX5cuUNOIQymR8FYGeiLhjC1
t08xteL6qq7aDnU7XiRWROUtVlpbT3wlid2h0N5i/1yLvS5kjxLTxchwHBGmqZmG
9H+kcDi1M9FUj6nVegdrVDQY1ETtDHVEqo/ii9CHiwBNQisIfK71PJqYpK5s9INm
1UKF8mVJKEmKU1/pzZ2hmcgEIVEvzt3LE9LeukE61WB411g4zGcjEf/PHADhy1Y5
mYtoHZDg6L06PfI5mFmKuwHWr1PcF26Eo8a3/IEe0V5etZpRvUyBVZnscqhTm6Gd
Swj9qMFIHEDLsSty8l0hiMHedF3dx6Ay4isOTucXUr4Sn15x1sOGtjRPEONFG3U6
xzgAFgQ43UOYDRLXnXsRydsam7KbBT8/n2RxlegxYh2wkpTDun/OYq9SSfBEQIJI
VOGfY5mU4upT0AbRwWz9OkqUofwdRYS/LEBk2lDlz1vfOtPe29POFIWbtC9EIxIQ
OS1+73uDsnhVRsHPzorDi8zs/BXSr4UjdhB4bT0PFjlW+/I3ehkU9JjfNhKK5Msb
JkaAF+M/ol8LuwsrvBUMo44JeE+1RQgWpEgKxfAw/AGeDClWf5Mdb1Rhk5E1QiU2
vtzUCTxWdIs6g2PNhRqfCa7JCpNFnxbbXHTOpCjRuDO89o2y3Y0xSSj1sCwTP+Nq
NKZb95juBLKrIFXoi5iKcTK6hDx18q1YNR8CZDN3pyo/x3YHTvWvfST10XNWhOuJ
B7E1YeKhJODu90FmOyn/mX7tGe7BCUnJ39nyXfZsWEArG3cR6FlR4uOj+ERPa2mj
gVC2pBWu+xD+IJ9AuFbskBxaa8/3+dCmYavdAlGWOCxmZTV35aZmVviqMkSVGJzL
YysHb/T1bj9EtK0BgyBUAT5xNtyyFVewJ95K35+5KVmfSv4n74Iu4BLSbLz5te2G
GQ2+3mNrzJ/Bgcqqor4TZrkH0yvQNvSt7fi/teiltD8AXg6P7lGrN5aOYtjYhwYO
pA3Wi+k+LMITzetEl0zqXCCMDMBkgGaFqIKncafvGF0PlbbuMDsTtO+H/V+QH3Yq
vgDM9fWW9enFQ/21AD7GW5HFV0SJZxY2Zr3YJxSvVlc7t6zZ6JGn4A31M+xlJ7X+
RoQxDa7vpfqSB9bPBCC+qIsrnu75a2+DA4mamHB9WiZNFUuN9VQBIKLvgSGHCJ0m
c4DDy/S6LIhD/KiRWT3JOCZ0TBHLz11pBfETD6lMciWkwXWw5+UPrEGUFe9yghh8
WsY/ZEEotITBbFq4jxqB0lppTp4ars0ZhC1Rv/vEspRyCVj32wnZG9Rnocs0G6AX
gsXnI5cdY5vuckf85phu6Yl431eWhWpEiRTkNJnH1YkHDpHCWKLHnwLlM0V8BU/Z
/pC6PGnk3BTmJM+YFvVbLOmYQk9qR9OzGoFsh+bG6Gn+SNkGKf5g8ItTxJteJYMw
vrTobvrXhjKmSI7+eIKtPLTvuQYOWdPjO835eLi3UbkfVjedZxMicCmmIBMCeI5v
UoRVtSjwozP1bA/GFvhSnlNdx5FuFj6RaDQT94qIeaDETa5Dn3MzSTOmyzGxHuvl
K/ATG77IRViXUm6foO1R44vIJV8g59Zrc73uWHr7wlTL1kNka2ptoJciLzOPomYD
dErkv0zOPNopp0NhdtQ596o7kmRsNJJc/DKVukmnOs6JAOkNLqCTS5xx27GE9YTk
WI2fuVr7V08UYEyUD3MqXUMquwHilvYM4WZKOBPfLnp3Tl5ttN0YtUrMDINYndue
C0QPeH4OM2UEo6fWfTxkl6zmlQM0vewIJIh5yoOSvS6iF6gGG0u4UcZqn6zuwCvB
3awofttjtju8Lu2vtjIU7qJJi2GGKtcuZD+5AFf8mRlhVgr89Wlpu74SRyW/rB1E
yGVSRpvbqemTiFNvaERxePX7eK/p0nHxZLZRrw/0ji1PA0lI7Wgu4tfE101x0Jk2
BD4mw4gFCYzFJgomRWzEjZydwgBfD3Pq/2Tvdiotbm0MwRBtbi3vns7+JE+tk+Q5
+K2+fvGEvyEz7m3CiX6I0CN/SU/Fl2OofnL7ETZ8D6TDqoR2PQ8FUYAM+BNlSoX/
SR52CsyHB6nkW6KW9eLVqcBA4BQyyN87CdWk7q/VmtA1XRJ6z2PpYi9zMPFXgGSL
ojelLNZHXDpySqdP154Af5ng66TVPqmXU8pNMPA7KXcBC5OPW6dTri5bUTX4MtFV
6YzPDLqhKkRCki3BhzAneaSVBIrNMsVglbjwQ3c77RMIHayPqc+Enz4n5YODMweV
pmaewZZs7k2psrThmjBkjBP74OxaCZhBcDWux4CZTn3DhO9LqdhCFjFzKB2eMGx0
8MaEh4phUjPgWM93SxNokd2Y/+JmrNHPqUC/dGIEW8CZTORlxk9EFmCysH/3s8Jd
11EC42jlYwzRGvh1sGNLLyfnvEALOGdj1PykgEWQl7xTlr8UFtfl+gxWdn4Z1Uq4
QhhgYI8uq4OM7MNRu8Rtl0H2H1k6MjU/MIyn/3AQAPKKCVRaNGB1VSwk3b/tgUm4
7B5tR5/cKDGmBTaa3X/rfCJS9InA9VHG9BfLqKR3+PEKg477eALPYoICrJEODKl7
BM6C56Ob9BiOI47XwfqEh7EzAllDUwgpToDEy1ZPi3svfZuSYbftFOCPmFqXcEP/
2lXJtzyR2b2Q6NhgdeY27Aukdk+KHoZSaPsj9UAXOjKp5W8NnQBpnBR9QzFC3FUW
TmYOHr2qLOalH9QiaExfKYfnNXaNZpolfsVenJ/1isvKihqDM8ooHocqlnXd/IOx
zAfFkQZoaLr5Bu8qhvxuSdzuUkWMmvWkX9QzGVjYQYK4aLGym/kP7tAL7j7RnN7U
n5ZabN++csFhSO5X3B37WzNorQHrrhWkzK9ZVbAlzXOnXYBoV9i0Et9oCCAMoloY
dmlLx2g366/Mf/mWGPEfD3OvW1kC5KODaDyz+PQdJYM3JPONoMUwLlJT0M1A8VFo
Iv2XAdEfeB6F+gvsYPsWwnKLzFL7eKbHij/KSBbJVn+D5+w/daxuafNGmTzL2wFQ
/hhn8fRy0fdFICz+rGOAMXut3CbazWk7kIvBEVuldfXRpdGZFzYz2iYlf/8KXKgi
ESjDo0U5hBylm7wZZQ4gVFN0AoFIKHac9peXM6VqlGmcZ4XnEdKli0HTuI+gCwP3
5BXgzgjChbjgax5iXURbzQjjrSY6eiS9JztO4J+4/9kbz3tnaybqY3lc30EWZMPe
zu6qYbH0aX+rkNMD69jz/lJjLVR8moYsvl0SShQ2n9L1h0+2XYBeKI/64IU9vjb1
Bt5uoTIKsAaJHsBj5J8AuL8fcLsbo5IEkzCts9ofOM7R4VSnES9EwFnPJiYTO/zl
YC3gS2QarVGMBUF34P4D6gOPlANZUxDVHmnVoF2VCx3GteT5rgmMCjvG5JON6+WD
mr1qK53yn9P1z9bQwKXl0USoZzMmwr2fjbHscYEOFXFcMYf7FXASDxsMg4P4aGIu
FKnoRAWhDeOm/AsWF4grkroVWpT6EOdLXV75eiN4xP/tZjEA66KEa4kuHNzlnmlU
PmRs4za3w0Tvt/6Zy0zC1VFfIipgU45wDhV4dFsEvdhrmbS/KaRrsjA9Hc1n1/F+
fNm/YQ+zzvWPMfAP5xw2KBTJYAm02L3LSzzEZqIIqiVhns6pXiO+B+qIs0HB1bGT
D1fp9/AV6M2rNbBtUt1yaIKbUw0jfO+NBwsB6pjBsmHFTyKqR4feIU1qNM07qxok
Wxt2hWOdblTAr6coRsYQpbIgbKg9GyqcEDNOHiZ9MQXo1QMPgxqQqNPjQoM60ex5
Frh78Ca3Ukgb7pRMzcKeadYwml7NF0wOqXk1JyGomD7rpJTF47RWKZ1xpUbKv88x
0J9p/xlzGrQf9gVPaoKNX7WYSZOsv7pz2WXoNAHL8jT+FCG2H/0EKoo9UZv7vgco
vbbLYr26eymTplkx8WjW8Q3SrAcCi0z+SK9IBnPIu0VGm1xMsb1PK8yHAPESdBVE
6Yl89GHSTCXtIrciqze2JtzYeH8cceFXzGy+fn8jzkFsP9ZoFwnHF3sko77rrJPv
2pwn56MROe2kFGkWNFPCsSHC4v+eFKyorYy5Z4Uy12wxRyF2/FpDovLHOrJp+kcr
kSBszskt7zrFWJxyf5oEYizHRAH54wZV2WuMQ0pSiP2RbOpms1Y7ARiYc0Iz4/eD
UFpdnwzqAEHx9UJ5bnckvg8LkepYLxGmzEXH7+Nt8QGcFMpbDs/D7ltiFRbvodeW
XJjTMM+oPpMcIBYB2rHUWN0VBLSHhs1scFH9fKLHoI5IRjvonxeVo1a48sg+W9at
mROTc3emWmKY74DLUxo/CoFpWTfDXHr58/+HJl7RODIWXMNnaSceeb+FxGaOd35r
UVRxE/9wyvGZeN6nOVwr5IXhiHuTkEciYDMKfn3AqqO9UZGQC+uZ/HUnLizfzi7K
yhDxduCp//jo7i8EJS6owJCFvd6nRX1++CkjhTkHcQ7EAKIB17+yYV/6w2ykBSfx
6x30BZNfKwcjup5asowxPWbEfvp3huiZTMJ5IXZL/5j6v1b6PkTkMDQ63oX9U4Xw
umYCglGOq+W1Xii3A486K7cEoPj94KBgq1MGJgVfo+zpXa9rEVALT8UqPXvHTaGq
tOZOkyu0rrRUiiPsz2/FinCU9RdASTNZJEBf0MjT0wmoSqJ408+M77E052pNW7q4
5tGUMOBLC1vKqlrxWFS0C3hog/gPgvQnb/MXcKJFIqbir0e5kJrAisuS0/CcLdz4
Kun6WM8rDDr43fIX7B9CJMoLF4IKLUkKyHXgNsgKqAb93+CjOrmr/pWSjyyPqAP0
h1IZLPio0X2026YhLaBGV+pAMdtAnJzWiDiVx5qIWuof532Vr45AQ3LKcXYPkpEH
+p0+6plKg9GUtdWKP1gQ9iYZ+e+0umTuopvp29G2RjpIzvz1eGdiVY0WyMmkJJ33
XUgqvb38qYk1zaEhFIRqO5EiRswH++CD8Z3jGKGLCv0xrrmr92qqstH56VD7It1t
HCtiI1RqPlAzHUDNVMq/TA7Wv95TjVAMEjXXarPQ5pR1k1BBf/ppz0G4B2SebYz5
ILKw5zApRCbhJXyecLaJV2PF8yjh7mXrN9618y98YiqSZFnqdeFXe2FrXFiaZ/SJ
yRldNf9KK9o3qw1KjYPDU/rYdvVETD75ZLsXV7JG92gUnAweW1G+tL/8MZyCV8ol
uz6boxUyj3z3+U8DnPfhjRdfwLLy7sJcG7M/NJvBk9e0/mqEmY93yLh63wxI4t9X
1qz9mX9HnpDlMtgDvqw7Yu+zArafdRZpej3EfS/k+iGwgUT8NExSgamtTRJ8EWmO
>>>>>>> 426889eb8ce467b9c9a9f74dd4af433c5046285c:deps/flexrio_deps/PkgInstructionFifo.vhd
`protect end_protected