`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36368 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
CZ/1hjxIYH4XUI6J5JyuXWYC6+in3UYJTphjGjr0OUqcrvrKlYeacSOfuXy7eELs
f+X9EseDy7pNWCxWhqDJWdYYue3unZ1pW2EZHogdrnhOXngpKSsMM8omDgKkU/Yb
MVBI/Wkw1uUAmR1Am75qYdD8goKBXVTjK3P2ucH/ZS0mHU5v/0QtSETUR436gRvN
LHwx3TYzYy4Lwz45OScUT+n9NP9GuOUgDti7yvtoGTbjFqXgNJmmOC8TJREQsxjQ
G9WHT+PlLRZNDCWb2Z4STNyFdHaRqFVR22VWxpDpCU7eXws+KV4lL6trgZrmeqkr
tIfZWlKlkOgyW01pcxhPc8uV/X1sKU2M3ha85xxmIQ5qzu3VH6AqFNh3WzUezBVP
KXCC9VxpI0IZKclEkvglae1HH5SK1pq1uYf8DGxgVq8sAJaK7CNIIHOW7ujoubRe
hTe+SZz3pQxM3NhPjKB9chLudSFeQFoHjns/9FPBHgKr81Ww7F7mDBlArPyw/Jsd
w1JUzR8bCDy3mEX4IkrANkXIzm837zF1+xX8cm7za0Mp20nZLWUdM0/1yEV4kViL
JdbqONn71Eoiwdwgjuyx025h6MOvqnP1uELU3ERWfwmKkSnv8PAzTa0cyqTX3BGJ
Op2jlNI8+0HNO5PmBkIz8O6ITHssqq85X6PI0A0H+h7FQ/95/4SN8OVDwT7slEFd
abacy34I3rwWzDlniUEUDd8h/Wx6CUBVHiPZMgVOTpmpOqYmKfK+9SLZ4xDeieIO
Y+KXkY/dtp0Ai080JwHcxBytZ1mSsa+17kTLAPNRwACIfQxAKuyi4VikaOdTGbyh
0mvUkT2pt69kDN6+62VZb+orXBzSSNUeNhfn+8lO7DGyQ7CxNs9nVxfPEkOQLKw9
RvRnC3EFAH26Pickw/BX14avWJ6JsZxzp7b2jikpZTbdkmGwWX7mzkb6iTTjuxNu
sq2GnsbXX1Fj3/HFVvg/LiPR1HviK4PYFJOr63u/y8ITmXJ9Gc3Wd1hBmYtbbanH
bPP00t+KCfsz0X58DCXvHbJO3O2ufoKR9qy6DZT53GThDVR2Tw8mEBAjxGVe+yEQ
313PRrhEEGiaEAAWP6qjrtogVGEOcLcZ08knVjfAY3Uju9N5wzft1x13lf5QzQ+b
fJPg3KrgVC1aHvfJCyaORQeOLCMmEgAqAXDW7kiVpAXp1hFuVAcqMJ3oJZ5Hfj9D
pq4FNawvhB9E5362STf8JGW2rbVoH2ll+NJYcS+D+1uMU5ol7UK/fPBHZmVeFOYv
gTCY614r+XztjFyI5fqxCSGTsusUTeFPhkA3Fgb0AqLN66iCJ88XsKhAW0Iav8GQ
niAX512nZsq2ScJ2TDhY4Qb1O742Lp36iiVpz3F8hO2t0/kfEjSHBBA/hL1rfCvJ
iXmLOifLrr1n2xy0cdfkr2NbjAS9ZlpSxXhMajPze70OeNm+WZntmFth1BN7LTCO
QaPg6P25YSkXGWeXeLhatpF82ibvR7MG7/ucLsh29iUIggWxd2+ZZ6IQxXk25g6r
K4eyB3f4J9FG1BAVyiKPnMPuHtNab31ddcq6OjJXd/BmHiK5hrJRZi8Jl6kdfTCI
ZiiwlX2HQodGnn+1Da6VYKKfdKzQOuobi5wqEuYWZIGF5Q33ZXOq5Qoiff3q0FNy
nYqGg3wf9EqtjzRHvzw42x0ZawiaE9iR9AQlEKSKsXvsBQHlH4M5qTd/v+xxcyT5
2ZuXPqRCSNIUPGycbrO3ltlnVCe5sU3ai/gvze+t/7zAKGvj7aAxpvXmIC0ZMoKX
/1puR3oLAFu4WQcxZGZrlKBrB8haC7dPcPa33L2WzM0n/Oy55NcvJ/831HuvyLvD
wE0ESlt3Ll5JC63qnnMkNnvoYRT7N3U9wJvUHLqlSvNBU/kmNMj19LTVeqEo5gvP
UOenB8Z1VT19MZYfv+/g2XjSXPuQAetEENdoiiGfnWi3vJ5qGDIbbvcM0qbOXI1L
VrG9EK0HV9CfJPVkPi9F1Zal6NOIKVmrQ3Sfq6+BNcBRzxlWTAdiVWWSYWoLxOBh
V6IEsAddXSfXp/bIAMyOh3suA+ZazjbAR9H+JGNNK7WQUit+pD6I8jkTQEA7o4HJ
c2ywsrizcunozs6evGLDVQer+4taNEFQyU7UjlKF6MLMwkdNlKppZDgaihLDy1k/
abU/JfDJIf6QIePRqygW6/1j7SOkXdT85E1/YKcQr5B4FFbkceKu+mE04sHCI7dP
E3szxdVwksWKejzvsW6fbg0TO/BYx9L6k0l2XDb3i9XGluduGjD1hJwUuqsW48Sp
xYjRlsjftts5XBvHGtayHjTTWHNefMdmFFcab5pZCgynho3Mi5H4NlAFmdJVApMy
U+2RnhGAP4UUd/5V9cL1S3jGg5ekPThjUPJY87DtYjD2PU0Yr89i1t7R0VdhKPtA
khosEKnDj/kaiRxyNasHG3U28Lf1u6SWhMrzM0kqNR8C9vr2EzFJKxKL2VKOE7r8
xb2PemGiol9Icv2PpA2UFbvo2TMl5xfi4d/O7Esrg7eWZn6q0cfhluxQdGT6ign+
7/QSeGDk9wmDMbUAqSOKmHciin0scPtKgOAjo2sbnnqQNi/vyKi1vhSjDx+z8KjZ
Ca8NIE3nmL6zjj5VZKG6MbU5NkiGmvIFHYhaQeTQvlncxzylMRRUH9bdogrCS859
f0l5ohEMX/Ki4aVZ/djiAhhfScJC2XWGoMppPfJusGYjg8nmxi+Bu3BFCpgIoeOv
G6fh8wTSSLJtVZZhAfNkLP5Ee+voBoeu3JjOCnckC9Pk1behxXqu9mu0RDqgn5F5
21uXXTRIMUVwX20C58LiGqPhiF/0kUGFsmp6Xh7a5DCe4X4YLlXgC2jB+dAbedrv
6hY7gaDeL/p+VKBNHJSUfGWEf6JFeIcJQjaqe81sxmlRK92IpmD2iaQFL+lN9Puv
E2JlhChxxQh/8+trxxQVVOqIjavauLJWsuUDwRGYJU4Z7DzsJ4ZnJbv+/q/HuWaP
Sis+RbiA6Ibdiv6/8U75gE2sMJE2zfcbagCEIKWXk4x3A4aHVkBMh7SgnI9QwfXQ
1sE05me1o0hEAyqtD54BLmdg5ILBvyf5r824Y9G2XoOBoB8mY6qHov4O6GTyWfHD
62NhL6hoQCgQqNc8dk2UhN+UKhEc9K/ncPz42upNmjjsmmfjh5FCjQf7IAuFV2EP
0jydpEKaSctC5IragbBwtz5pp1exZBX2KLbsWqJcGTRaWiWFzZnQsJY+DiGblI7x
VylBsddtm0bSM9IDxLFj4THz3Dn1Xtp37Up3gZOdnUNs94HDZ6ZY3gMgrx2WbpSK
WirAJPi/TQHvkhx0NIU+bo9SBy706xO9G7AijQOWo+1C5M4G0qgqKe94U+vKBKYm
3pqBJxQEj7MF1dfdmcd+5n+X1LLDn4WojIYuHWzPliaYEPfOsEQlU53UQzd/+4N6
tr0AMh9SFe5DqzSSRgfOVWmTx9sD3GrOqLH0q5LfMuKP6iaZi+LO0RupUtn18DPm
ITazTICjKs6Z88eK/0EuTLnRVI4LAHUCG156b9CcIsM36LD1Inmagw6JAdQedI02
cI78FZD5s7l7RL1o47ER4LdQHIqmQ9d/CupgYwZWB8SJ3d/SdEv6UiXgjtRPIUtz
2raaLzaPMHMs5g0YmeqWI8ROmNeBAhhJzrDgogQ9/as0WbYl31y26uz0l5As9x1h
CT1+NZX7ELn3ctTgAK6sRS1kvTh/ufs2a8AVHUjjdBHWZzMnlJw9a4vXAwJQ7vBf
6Z5aQnYQvt3xK4AjeBiaTrPlMS7VVKGCgaUAMZpF2cog0fzJVsF866qkt2fX2YZd
IeGnL2ZTzoD68doDraK85OH+OTyjJyu+7L/CWDTZC1ZbPKfmLNEUsrg9OAwNnosz
guL3rL+jITqDqiytWRvcwwjC1Sq58/fCdT2EvUWmD0KXcol1+qV83NZ3ZtAXBBbG
c9hxZmZyPYBxf1ito22xrl2iC9tMMorXyQl8whYf+4/gnye8wKFnDkTmTR9JQjBr
kFiNjKJNlmcsibE6cVK9/vQnJcHN036R3Qik5xjGOu08JPbTC243yJMS3ASjqnCf
sM3UCP7DIt53yHVqZDdwqrM4ML+3qqrnkrd9oiJq7TsX70HzrjRTLeK7sBWG/rnO
jnjfP2dY6Us+rWMiLe7wUUnosMrnsC8tDeNhzzixBPehGNtFLHkGtaD/hjoQmeC0
RJFVlHJgnPAjZbZe+GDkqjr8uqbH4dsAkX1hIfuj7HfCW2EkUTbqbEjBYwR93ky1
C13hgb3J4/IHI415aiwcunlGcRPpQBzgpNJYYYwYN0DXDR3R4VFa+6gXyy/J4IVR
+MQmGewcMVynr+EYD1Kkt/OSE0MDUSAGvDSDLZaGLyRBBdxX58MtgajHrRJGcQXM
34PBNtpoeAKS9bc6Frcwe+v79+bG5E9jPeQXumjnYY9BaOPRE1dC6xpjV9NA7q6+
aXl7Cq61T2/TOjGJLcE6+YlJasS8YRwlaTUysohBxAJ34OmG9q7gwJJweB+kU0zf
W4JbaR2/tviDFfoXosE/ylcxrZvTWl9c+bn2bPEnp5r0sQIkvgEc2OjmxAMMHQT8
OlkLsGr6XCBCAb+wnfKzFDfQIWf5UxaESHN7dKuvorezKO4i9FR7XfLKXj+YClV3
CmuxrK10Zeuzh7l4qROwVEuB7K9flvov55F7DYyygGH2A7fGLRvvby73oA+E4w8a
AeQ0TPk1ACvH5EEWuHcbq1xBiJ/4i1jGFqj0tRKICf7/oDafgW1Xi1RA5mjIFfWB
cav81ILjkb+Jh/XU/6Nx0eSkhMk4/2llulVoofbytpLQGGQWQ8y080XLgxVxgHyh
nAm7/IGH3xLLWosIWR6ZK7oWuc9jZoBWzqPr1Xe/u1b1MiTfP1wYEuwEp2YnNvcz
cvvjbPunzI6AVwk4/QOXabtBCB5RpPkY1aOUE3AtN5U+Qsf4lJkkaehnFcOUODJM
aUF7tOro+bGSEPwaxv1CFU3VSi509vqOLDfyDmUaXxmHE0Hbr9vGQatht4GJ6fDL
urVyKhBg7OeFlRFxRPrERepT3vVZS/HWIwMRe7cblGwViL/eofuCL4x6lKndMx7D
FscJ5zNmJ9EBOcub2K3dYNf9cdoYrYoZ428fbdWTiws7C0fFZAX9ZP7mDIjj95Iq
GwSQrFHRM+jxs5omfIB68pfCAbD6ZFtAzM5AVh+q3fZw4hdiwWX+ocoB224+TNAJ
WZ9dTCPQ/UgxYNmmXHV/RaNdmtaIKda83VGI08CRf9wz1qsF8yrd9T8+yOu4uENF
59oVIud8riZ09y4cD7O3osvh6TnranEIbvc+7+8ECOb7raoMdFReQZ6u83tw7zcu
vRYz7/iJt7cz/p1FY6KfEgQYACJxKFyjjL+/2OksOBZEnRISeI4xPe916fdezmuM
WIU3WLbX2irhiC4Y04KLfKdT0gCLMlH5PhMus7jyycAECkBs1zMxQcpnWIJ2HtRi
ieMdAk6dY3lmNU1e1zp1jzdJ8C7BfTtjKnSiGODr6+7/hxrizfB+1yC8fxkTJm5u
WlJj6+3G9jLxj1Xt5Bzt7/4WlYRSqpY37Y5lzJPx3Yo+ivCsv7mfoyV2zaGU3nbr
QsnzoHMRVj5F7fmDkHrOHrvOjy8XkqIM9g5hk+9AvEpSbYnXDCJ8s1FEqF7RatR/
bWQXbRPnzRPoYeRK7KW4kNQQegm3a3cBGnQghS75ZJU5d9f5xifj6zr9cV9xTvEa
/7MhgMDf1PlZ+GnDmVq/d2/scyggu9tTxvxnRr4imYRgP5EFqteGiObHUffyjAaA
VUCsrMF+aTyRLAeH65TssaHBm3yOYrlXSw7do8OEzRhmn0JPH04kad3R8lswPGB5
vRavCSX4Fe1AvsZw09CpH2XXNN6c8GHhxv1llW3LfR8fQAlPnwJ0ngw1w3IUk2ZM
JvgxsyxV6w1tj9R5zb6Dkn/D3Zg55snLJOSaXhWgweBpI7mDr9XgvkRmm41o1GOJ
fzPkkP2OCBexwnNJQbt6HsaG87laiMZTYdl1AjiRW3jlCWNk/6E48SwPTNGdvhmA
OeEe3ldhijw4oNkYs0SxfJNuGAmbIe2LGRH3hBUcJZwBcSHOQhecKdDgF8AyHBbX
aMhwZVHO4oaTbVAwTiqYNlPEFuCZboRL6ztjqfvAyIEkuMccL76tXwiFVOmR82QO
yqGI/7JdjdEGo10d5VptwHm2u3dAfFZv3ZQPbvIgH0WogiHaVHLLQK1gA7fylFtw
Ejsk6BXeQ7r5XLG915ue/abFtyvV0ymYr7FY2/NlBlBiyA+6RhX+4UOZ10CTjbcc
vyDPUFareXkz9BLfT1MWQY1hW+MimolX8nbvCe65d4PkNrIUecbuAgNg0TDF9BWk
nOK2+VdgIh3lg3P/sPmbi5bThmnQkeNGg6v83upIbQBNIRPjSgp7lS/zw/I9F3Nu
P9dB/wMrnwq4GdspwcD4mm/Za3UNr440OodUshWOS765YjwYA1O97puq9JBL3qhO
Vkvd9UWzBN1cWV6ZAHCFYb4Sa9vW7fo4qFykzPETRAHJPd/N6e1XdDh2DJ5sbw0B
8u4thGD70SI5BsPmZPn8OPM5quIeaYN9CrY29zC+aSudKzioyn7OvDDdk2q99+VT
OqThkrnlRaAGOz+xBzQSmXh5qu0wQiklw3L2PNaCHo0FWzZLxR1B6QSBVMdiLkd8
fzB+LFWzzmybwtwdcqDRu6l7lZ9qjr/3et6b9FpFuoDGVbrPzV7ZHFXp49KD71WY
aF5Ocm+TljY1pNDi4KBRgsHl/fC92cjmMBvkrg7kao2Kgg5pPAEK5OJZdzLLdz6E
dcE1heC7Ocrj7MgDFVdFWMd51H/faGj5oMjal14pae8o4fIouqHUsOlm+T8e4KYg
vCU3pOauW1t914MQT94kfgCXNntAj0/vpjLKqqU+YuPeD8mzqdqkAL24u/qjDFXI
unjdgJm9SbSf7/d0IZSKWWw8ppdhALqJjDtVJzcUyuaK1TElB54KA9GRje0KBa6d
HWV834lhitV7OlEufYpQSN89w/pBcLfntGUIDhekhoHMK3Wd+Cl4N+t/zNRGeLNP
lqc0hTngnZaKe02EXGPg1cESH1yFV4XbbH/xfnIogzjzDWelQ3+CFGtMt+Yknxo7
dMXTMFp36kDqFRSS/gqOz/2utjE78p7HAUHEk3xzDtHjzx6aa+k94RieHS6UKlh6
FH5/t9Azqvs4zD6I1r9tyhOlQuGXSp21SbGhiCWZN9nmxxj4vLHmedyoCWgwxFkb
0+ZevbAzo2ZE8crUxUn2Cp0cGb6xW0wuLhebUJFBxEtTFVLgLCCoYeHhVfzutLC9
uVlZAIDkgfWHDoIysMcLej3BRnF04+iazA0ZrdLIWWNvUbLI7x8pEJY6Ga3h0m5h
zaQOEYU6PlR2rdXuFiU51ap5oSTO45rBAfplcQg/UlhBifGGj7QN0UMHtnQQUF77
qWl7j4y11jRAkQWQtJ1PLVQHNdWNYE39EcHW05Bk/4PSjdqcr9DXXHmzmbnAKsNT
f1pkb6ER5nwgoICHuQ8LRt7K19+LK6bJyH/ilnzvyjJ+ENDxoOfPECAZwj7xa0hu
hBxQELwNU59LjP1assTk+rPqOhYIjNeR+IWoPED/mbwYLIQNiutYSZ3Ter31ibVl
kHMzHzQW+EQvw7HMUYXYbZ64kR1GJmCPZpbTeA676n7q1BnA6f4q5et1lAd1u6Qe
03OhH7v2QltseuhViwRu1qw3Vn00aXJlVAFxRF9ZfRna+UWUhg1WopZAc6DPbPzC
fnGQSGJUE/snUtRtFxKlxI0PDSsWOVWK8YpDL8UUdNedOLhVrJ2mw8SBht7DL5zP
QJNO4p6ypcSBs6uSpywiLNWlEwHhUD/TCWXAGDLUDgtEJCIgw9SPm668efeyerul
iAw8Zef3V9u/wFmu4dCC+5je4v4YXn8lTRQnZYcnqstBgf28ZrvZGg0snHnNf6le
J1rrXcv4e/vXFYwG3ZaqfAAfnLUZGYY8EJvHmE3fVzTQiXAOJdqRPFsvELTe5/6T
NIpAhrAnZE1+mw20k4YvbCnDH5fmG2Rz2V3t1gXU3HW5VKnoycMl0dLN6/jlefoe
FzFdwktHxyV/Qf+H9eVmD4los2XCLjU4X3JVtheo1TcDk6PNH6P/e6FDHx2UxcAS
cKX8JJxGs6IN7PzfVrUj4qAhESAzaan4L6lND9zEum+osMAusXEyOIKSPgHmidRA
OR7s77d273UML7aoz7h0pDlYcYi4EmRTYCj6N1CTPlWmPzeTOKjWhjWUFSxd005w
evpjpSNMKjE7MBeRZuddNladJMwzb3+E+geTxM453pl4d7xo0dc+jXXX1wgeOl1r
7RH9bVSZ00escTt2yFfHm/622xTegT3VaDC3da7rIaHCGDQ6xKTBcsmcczQN6a9k
yWQxFhNu0Z9DwfSuVjL75dZZieh1RyxcfFLL8ZlarNdbt2jBZhRw76gBHnsKo8Dc
RN8vzLtJ5250/f/LWDspLfUATx6u9IeeT2/G/R7iMj8UgU08ktyRPqH8EVIfFE/C
fIh+0QDQFFRJudnNDXa2JANgseMMymXHQ/D0SrnXkrPlON/17rF9JLFr9Meapst9
q7AtWGidLIh0o1okJcjFbjzWb8gxXBZIP1Ys8BSVvGts3mWzvgiSeI1P+PvW8Eu8
X0aaTn/pSIR63qFTEcarkHd+OBM/5AaZZnhlwPNXhPGfOBh4KuaTHijM/vMNesTp
g12IpwaZ48Pfocs3zuBfUX3Y2j5tMshnI9bit39hczxFIVJhswcT3rnchiUH3cc0
Fm0az+qE96+vvyKku72y2pWtrzcezKS6oC9inDLTHibuvixzX5wF5ol64k9xUXXt
RmjYJlUC6hrJoeBE2s00HdIwCphL2dqojmXix5OyJTgCVPaBIkHIlM1RtcFmQ41v
NKbHb4nItq0OPn0Q8k0u2QFnM1B9/EKSpf3hCn3I6QZkkDhg3wQwqoGw9l/584Ss
gJCpx7scUVuFmfIyJzX0eJJY0bM0evBDJOixVtFu54NYbD5sMBJvadEvVq/T6uTV
1CMDavB1xjOWS+68KmnkjjPeaX2gDJje8FnL4fKTht++rriJyt/o8Rrd6YkdZQBM
BNdMll2gFYyYQR98kXzszifzXtK9d1HXTmkfUMOXItgV9+LNQUzRyxIEu5Tc5jvB
mVVuuNX/p+gUj1qxFOnL5sc4wORzY+9AutcOD+wrhFIen1GDiJIAmuakXAbBrq3C
kpEvRXfuA+APKXcD4ttZS6gjZ0L7DnH9tGQLgmuP6MRd9aGj5G8D9KhKTiOR+Vik
MEn+w8KYefdFEOipJySgjB7DdxfljEXJGKo/neozAm34v9+VIXUoPVcf5N1JtQuG
S9YqOyEI5NcuVJe0NPCVJ4rVdM0iAv4FmmkHtXxpVytFy2cV9uSknkI5+zqeqs2J
ZavATvX74pwUBAD274Tw1zJmj66+Exdo7zRrcHtAFyVKBO7x+jXqkEnO7A5qZ6yr
cdCQaIjU8hOcWg8y9gt5+KV7tQJ2Y5s1bSbTJ4tNXtZbF83q8ChnirZ/ZCdKfshT
69mG0k+JxhJfAPS+04wwMI5oV7cc+6tPjAk9tth0eOC1lSqRgoPlKAgzaxqtap04
p3E1p7Yy/F1bmft3metJQOXi9teqe6rwdL1FMn2LvkruAFcPk3d3NMv7msmaLpvm
Lh3f2nzjrp1WQpLXZ16s5gmo6jLqCY8tVsY3PZoxs3G1nnO4BH+OgPq9sRiCUarM
afiIOY1fagz2mIAYA1kcfmjbDfeO8VMYrUyx6TyjdMBQro3BQNVdTbOiG9f4Kqil
Ihd34B91p2Pp9h4Y6X6K+Cpgg/TBSq050xo9nkW7MCL7JgH4Otj1VYNTk1MWZORA
guGDg3YDWiYeJ5WklQYlUSSswRzbvHSNTdEZyEZPrU+KXLaSCGHasC0+x+Y0lqaz
RDyUj1JtPVuM9j0eTMFfG0Y5OFjccu5a0oGfznzgAWx0qefxfD+9CWpRp6qTqFLE
H3WtGRdc3AGjyQ8GPCvgaKgVo4NLC+erdTVqBXc/WF0J5aUCuGn0uAbjLcNDUJdm
Lxn7xK37bQr56N0qElfvxZxUNfE4VrRd2TFGD005s88xHs2o0Z5Oj/FHtuvikyQ0
GVb8qqYddvmZeWCa2NnI7FK03+2ScfqMpdcCyIpnHj/lAYSPtl8+S+A37jiWvksm
iwwi+zqEiUts/uKuckNm32M1x8a7zsiO25PpxWomPF3UY+TC37kAA/EyZatUBanY
JTmwj1afmurVica76fv8S7Q/nmoSRrruLGj85mRPxIrEChHI5BMlwC2nvC8DcojT
LRNmlvrhURn+B0T85HblbsEvnO17ok23NJz/EKeiPjmtI5UJOaPli56xJESHnyV6
8hRGDVDpzkOGb6k+ZMykD3pdV/wfDfvKtyUWiWKQZfXw24IfNIo45ISele5RJdK6
zf/BecRmT1X5xyGHTYPVbyPspE+SxR6Fu0UE0/Yioedi2+nVLj0jU4AEBYwfFdyl
vzJFVdVp319+57uWIOQqTTOXsajLZOkTCceyH+Tgmwhlhg94ERQMqchLjKjnT55E
xFleNuRTMb0SzCgxGpM+XdcxVlcMTTdyXuDkbN146AsWxDS9JAUBPkpkvZ9VJVGN
m3DYhYc/lDZlcwIm7rJFi2oTL5Sbs1N59Vn8RehGLW1kwxWFW/lqHjCkfxBpyboL
GEgEosmJ6fmMKlX3pTKjSRQ46QGxIAN+bnKw5wfVVRWsNjv4nsif/nT03v3MVK8x
x7Q7wUpK+C5K+J5nDF1e7t5DZA67KHeim/X4Wd/AZL4vN5YTscAPF5sYWxnCYRiJ
8oBCP2VLskfBh52eUduQGDXDFm6aYpDwfPGCe3Nwjc1vI9Y+njYrcECNj7UvgwL7
ob0+26cDt8iqoHmORSrLixUt5R/j1vNbpJIcFoCPyWrxsQqn7IC6e8TGjWSYJsNX
d9gHTth4/C10gOhlNgKqubaazfAeEkIXaEQ4/adwEjin22TnnLfXlwd4P9sN4ndM
3XCxFl9kOPbCSqu92FOiRmGHAg9EiJ6ElSUK6k6WCMESSTCT5V9kc6kTg/RR67sk
8UOh68FfK0/RLg7W1tqGWJR7VI9fx5m99V0bu/d7JDDzHqbCUmBtVxDNzZrmsOfO
OYmLk9N2Qo/GFRzNWR8PceVyHUM1H9ruENJ1DpE+A7DAYtfNz0JlTXC7YsrSLM/b
6jM0jkX6nXaqqSMOdlFt83Z7ktsDh3BJl3+s+bZinkoR42Uwz6anzrOlQPlp0+Ok
sDJlbIgBC0C+xZsg0anBq8G3aeWe7YA8X1dL9Sg8WqctdaK5Khfzz5Jv8snHyAPi
EnNtbNFqqEAqrtNt5ekeZhtKdJYX0H36tkRvbVIpPG/EBosfuAu8TWabm5C6mmNI
xi52tpPWEJgCgagB4ofewz+6tUKQVpENVRM/i14wjVJYJn/+oRdo2BRcNL68Zj1K
tBKlDuY2hfUpveAMC7PfPEWRHsWBs4/vUif50LZX/YLOdknHYLUSN6xFpXHoSrma
Q7ZzCtkU9qxnXGPWEIX0RMIRH93fpcLDQzyXnF6LSPzhhJB37etpYLhSDvYSn7Kf
wym7wreDO59+xG/1fAsNhR23iP9V3GFtcIY2n89zw6cfeEaM1QcVuOBi4dOGbg7r
sQ+4JkUQelFQxHSD/VwFQBkO/tLA6L57ZvBv178p66SR0bzbi9nnMQiZYDYztGAL
UDhORB1Aj8SlXemarKh5/ESoA1HEWKMB9XBps3EZbwvGfhJR/Lmf6515IzT6CjFT
pNmFTChWhdFUnMz3ARSnTy0XW/v0AdTgfi2UwUfz/6B6gltNe4YZlZEh/x2U2A7L
3PhwGIx2Z81bkDFKgIi4YWF8WLtmtcbKKSp0SUfoXOcIhVZSO93p8gpxHhc3zxuE
fh7WljXrT7GnKIKDqsdz5csmBsnD582NxHIcLFYX4MNB+asTmTp4ryVnKY7/6/nL
ADB1VsnGIgpuInLMXIDpgfPvNHfCGxH/7ZuI1tXmz68cWI3PQJHoM96dH0VQvg0G
Rs87SZtR2DW35kolJDxKv0H5tLGmG1xgiYlRVt0OvgAXObia90R+F4AxhIPlf8tP
s8RVHCeS/WbWvhyqYuDY5dsHbUJl+WqQ/FnX9fNOBetUcaPVqBu9568Dc158NA6r
DtF8ev/Eq22Iri6aQu3JjcvvnkPudGorXJ7/EPlxKZ5A23jSf3lOUjVHy1BmAmLr
Pce1ooarOntVFybqWw2ng7td2ybKrL1vXjFpxhO1eoBAevO1lPmaCdiZHwHbfr0x
v7ZOpn6R3GMz6faMoDmnyQivwydGpiOxcEuGsPRIcEWZ05PKeo3NiFYKhwHO0NHE
5A2714C3te6emvXOqcb0HPww0MnmbBMmY9fXYAg4ybfRKNXi25D1jG40zaGegmvi
roD1nTV5dE7OP6WrolXk/quo5GC4YNDs5uBwSo2TQbPVT2nIHGLGFceFhF/EDGLq
X/M6A3ZOdYArI9wa4AVsXiij4563fAJrGF2Z3pUJFA8EQPhonf0mNOdHyNa7ZgwX
I1UxvNLJWKc8xrDyevr2xeIXC3T5MFpOHoi3/eOkUjjU4nKYdLI8UI7qzctmWHW5
8+jIs2SobZg0VQ9Dw3qlLU6yHzKFeWZ3DsQ+aH6eqc9iPd9pazSUY1XDAxazGyya
Al17gNX5kHf6N0aLHtMs9Zy5oXTC1ji+aHxi8HY7q4UoUWhfR3RBvpI2LU0ekPm2
ReRkRgW2f+ttPG1ANPvcVlDzBeEKH6nKzAYlmz3GsxoUejKWcRtM96LokV7k1+qJ
bbdgNam1+6Vm+JMh9Kwk4ArUlA1hC1fqMIqTJPj9D7dA6hIehQFehMmodwMbEweb
tFa3o+Q2rxs74A2SkyQGJSJfz84H5uHW+3boH2ggePtqRek2WBTgp1sC0z1njLmJ
aCwRIyhYPcfbb3BV/+Jl5cHjnJlKmhaYes9L7dVaYxZU0IJuZDuFx/44HD+GsXTX
2qfLVDfZBj0I3lfe5LduTMD5KYDICiOIJ561uwFGXoa/WeLRbWQubn9/b9AmmHR0
VvHOFApvLteIlZDZa46Fb1i57z5GVxLeSbl8H32wieXmMucLc6NzcStB1sHVQC6l
Q7pdfrNitBUkIVXe/g8jEEhRjyYfC6k/O1/dPSkskcIRG96OTeYkoqQ07oNw6lyq
cXJXcF2Zz4bb3jejqOsFjVPhZZ5sEBrvoWfrINy/jJmSDoh3bi0KAB/VKI+wNk6N
MYRCD0Xe/Ui/TikFMXDwnkSw9OVSdCqkda9GZ2xgXvZp44GFr7CUeRJeRyY4JkTf
/dpeiXNyKTDswjxBUwO92q5xEDeV72N+fNUKNP1zg2BTRfCcI4i4JTfY95mO7N4b
WvhTatxcVyFgTeWpf4mx3/N4HFnNbiOBw3DbQ7mW3MUjLcHej4IshYgx6HDqjcM0
iBe24afhX127H2JywiWhZZ10Lm0loX3V5jY+WiR/ZnPzl8DwFefc/sxaEWGuPgqS
ZA8CWOCZfqAwkrhhZ3Oem1bFSvlrODvXZ5XpF1nBZpE4BoluLbzm9nIUHxyNzK4K
160nwvolwbp/qnpRKT7BDxBf5CiyY3KoJx2InWLzW3BXXhjsPjpsJA1ky6Y7pp4x
ljqm47A3XbIjOXbiotMyNV6dfs5UUiv3CDzPTePouBxORrmslcQGCLhY0pIEaBX+
K8FcD8fhheLfOo/qPMGVEA01oCxwBfNXyqTwv5MLbV7Nx8qjFdlfnQjYsuTht+At
76CsGyWpDJ+e2CxGjnkjtn7GVZkZpUUtcn0xD8w/cb9gwidiMeVnSzybcnwwGbnd
o20HBichcG8Vq7pGl8+gf6oq1VZvXGPbqoDS40dTuN7xdSEzt1VKIGK1TUN03Lkh
TwkSvhnhIAiIYG+1Qt8FlJFgy1csCmWDabism8Uiti6eDNQvPwtstjOX/3IaCaEB
C3SBEMMyHcbP5ET0euZ7TSWksEmfLBviT0z50MIcuwiUII/EnP5pR9s50ZxqFNlQ
UPvwHbO6kpSYRV+ACffhqHrVbAZt3K2n/dCCH+rtjqtZIzKKjYWBAg0pJtkeR1rF
/ckNvdJx5t8K+JKwNKDv1Yk2Cv6Kv7Q6g+QjivUngvdf8ufZTcyKJW7xzbcs7h3I
16LPNVyjAFGXPs4FHTRc1rYm9lw18XjOqAIXsa9Hht6yPEXpJRUmNhXBy3QtMISa
gwtLKDcjXxMx/4LycJKwL77MF7duibvkqkuGZlkIpO6WSCbxJGvndx04mO61WQC/
op+CNhlgTVyOH4SUyoQLZo0VScMdqxNKWSt38/qfAJdf/+UtTLYxFSiOn8HAZbmr
lmp35qD8n2LLkd9mgpyF+YBA+LpqYitC8DzavBrgD6sd9UNMuI4VXUfPHG/mpmEh
KrzbxhSLZ+AkYaH07GA4CXho5Us2NK2tRKedTXgT4I91K1w9Xyj009X3/Wp8Tqyo
s8sOHjUYFtVxsbE+u85CSH4opCVdH61lS1dfjPV4miC7i90QATR5j8JMswzeVp4r
LIRXDGXgocO93tcVCtX6P3uED3wguk3nkJ4pFiX2rVcVaJ/kB4YMjc616TCkJcWh
E61ZNSnEgw78vwZ6tGwcmRD5nvqzJyOwNZ28vkYdoderxMWadQuT2S+WPiOx29jf
25dhyvYqZqGcXZUERoEiiKpTkjkorUeXpAxELVRPxw7hwi6aaBv0KVS7Dn1SuF97
awL0W/lN3VViQtOXVWab2xiTWRi3zPenuVK/UNH0t2tKbXMjKYTOjX0XR644v1W9
TFhvn6LC4P5TDrzGYZGTM9NHtp7gmf8j2vA5qzNnOadyOUiwwcHRepC/3iqR/Gm3
+i4kU5OiCGO8z1MlJgVLHTdySP6CV+QRW5MHNb1cf90sW3NGPv2g2CVtoK167STW
DbDMfOajBuROhBcBA2bareDK484JPzfPKHsljP4twg5QAg4Itxg40TIQn+X+SmZm
RTop5Q21e74vswg+vTE79hHYEyJVZJHbi5QfcmuCchPFyO2rXv6NBuiKaeg+c+L2
lpyNeNPBwxKDgbqghxMdQhLOwkQ/UqrS0Dj5zZDZwKM/iaew1SPVDt7V8WhKI6RJ
4URlUw+1SvYwCkulgniq/teXScXh/uKCRXqZLW5w98yNf4vwFeEhN+Iv94pqrT+N
c1IOb/kZYipXZOltSHHs9jFU1eKR4hR8DIyUoW1aExmfcSia2gtnD6aZ+2feTjft
I/5wJW7mdykeI0odytT1tKjAh65tooc5Zs30MCAi7pv+CAaDkzRjkX/CKYdggwZ3
OW1ASuWd+cKHhqafE9cwn7J+5sPre5xb4FcQCHb29vTC+pxVN/c2gNCIxWb6nSt0
GX1PAnIvudo8Wl81FDjJwLdYns8BSs4dHdLdIORoPNLeTItvLEALC38cJ0Bwt9Mq
z3bTR+AEPmMT1PVxplliIm4dNKaNaqP1DVprYXimKH4q/rgtLtBKiUwyW/EFESnb
/mb8CywFag23Qwtp9jhhnw7/ioTvBRTYQVDYrdtbeCdIREdKBROipNBaqoc3J41y
HQi54RMsJ21QtqskpeAmqaXFzOkyLMpgqxIsMMaKU+SitcW6ZMy4FA7iMoqQcmcf
WLv8kEIM+1Ce4n3jf91lfTTFDo2lH/g2uL0OWKrNxuchX4eSGM0+D9jLdXkzmYeP
tolmZHedTfL0bV/igO8+7w9Y3AVoJhjUYWiy2y6M2SQ1Isu1fYwn0m/E6kw2z3Ed
CdzBUP0OyfrT/lUooxYuZeyHTQXnAAJo4ZCEZxnC89Lswccbq5ynNHD24xzQSth1
1y5dJ41mKrbO3GoSUIPNzmVudT/O9TVkod9W45q3Q8+s/Cpet/Dy1uwUTd4k7RWs
o5UJ2spVPQdKygrLel0oTRErNdWSike+LrAjMgEkDxllTonIJv6s70w6sPJKch4k
PXyCSP4OA52pKiXhSUgNuGzkWrz4sYY//4kN04S1XnuXfvaRRU8FswaSJVzDUHTA
gKRfrg+C+VNsQbhXsGC4rF3mK5LLK8rJ5yyJGrPO1RfeCCcHOR3cI4WD1tIw4g1/
HaEs9cIYux+6ICUlDtEAmZ5CdMO0nzQQLRbIoI4pcA4JGDILPjTpxb6xpERTz/Ai
f0o+XR8AFelhjj75HmlrzNIE3huGBnDGOYrW94QNDQvEyk6Orz7ObyBdpeCEjVRw
9D60wUt2Gtgb+bbcr4s0YkpnmVve6bKoCB9aCARIqnduhQoJoGPGXY4KEQ3Z/W0l
CvH1y9XemLOi2iSzUP+rk9cxXpj8OkML/WEEPgCo0Z8/yFLG/Ff2xDWKPKejQhZl
SpP3EQAuieZtvSeFTmrvs5ymUQQD+emFDJIyP2b9yUT/x8Xa8XlrGRjxjy0yX0Kb
K9Pm+E0j4vrIlNorRJC+EksI82k/vFrIETeYeb6Y5jVnoKoqPGNB4PF7fHmOd64F
tz5U8cev+v3Mj+SUwiqaivJbTkxeYYeAEi3zbZTg4RH3+7JSHCtaqGYlSqKTVecw
WDMk4fQGN0Ahv5ZvM37dHD2uDUYMOMT3aPTPFBOCVnKPeqniNd0PTOH8ogu5+uAy
WprdIe0yH7gT/86m0TT7v6Py3gwzacDNX4BKBgF9XmPO4JpR2GK4/saXB/wENlwK
hZ07BLh6XgdojPppNzqIPh9BlkBvyA8+mmg+P1/XkZAsksGaoh1WKrdRp+3ahsZX
VfBWSfGpWqiTqO2DsYMH7vohF7JL06wZaXubaxxQk5rzEaHdoG//4zVccFJk6kLy
emp0RyCjQ7tAczgBn5wXSvq4iFcp0kHVpcJJuXBM1PVGHyy/ZR6+HP48C0O255rP
hkDGiJ2iZeLLrGfdMzQP5RfRWH1TzK4PhoPVHgS4GOXZVX9Tr9Mk422NVTNTfGhO
7hT1AbaHh79BJr1YBprFLkdOx+f+WCdJ5uZp6GF8r4la0ncRL5xFuXA62QQXG2NC
v+SrFfC6ryUgSCGvrE06xONRZC4xGHE6SbEcf86kpzxuAumxAmmaEDt1c3jrUB3h
uHeeP+I+f+2HJhqEQNPV9Bo7GotUBAKQdwe8RCY6XUDhKbom0VWd433wa1/dbLNQ
GtkmCx9oKzlItq4ka4GC6a/+FY8J3MaGUNXhqmkvhuGMQ+aQw0HIdwU/WVU4IGtw
wTefScb2/rUFET3pZ2NvMyHcfOZFkn7KVGHl4/7qqD08R4x9UORcfOVT+V4QTTd2
HUggho65CGyLgiw05ShW8DEw2uW2m5Guru6wj5kQZ38Jr0yjIi4AbGfFJalzlPxS
NagBcEsjxO0oktK/kPdTewo3dD6pKywgNTYFZwRSmrqodlg9wDlXSrnZvqz1pEiz
6OI4L58LNZVtqMMqwlOonumc4mZP8+JfWrqJXcHLa4bePErg3kDMk4yXOjbdu8Pw
ezOMMqS0W+Hd2FTrW9FUlskn7MRcXCxtLiZ/CFcHooq/VqTu+dbiWkPLLDQXD5va
A5tvyoPt09eDPwaeZPmCcY2v4Jb4goDNEmeUQfEO9K6QPE3oHovLOzCeAumZyZOH
cn4X0A62apVmXdPUmfnNJxu93MFPaCM1O2DtvSqsPLrRclIyL28BvSJO9keL8ntT
tA9AAkck1D33zVva/pMaVX8X4cOQ2IKebaBZD06levSUO+e4aiAkLQ+CM2v3WeqD
Ccjc8s1iz+9UR8UTM+0VkT4amaqe/rU9OwnKDHRqgGNkDPbutJ6zTUU/ygzCJrtu
3UY7DCaGiURvD2iakkzKyBpCNdUZnKpdiiMXX01me2a4zKRgPy9vy4fUW5x2PSUo
csE0VWbqCNlBP5i2CDMXbolqS1lua82DYe+S/u6Ti0ARy4psgeqziamSJUsI8MZh
UfvsfYqqf+TSYmey1uqnG0Im5ZW6oBN/Iy5auEzNayBo4Q1ITV/oCM/rhaxZKIde
mA93BKiykOoL7UhABLN0cO9QBXQn8foRN837154aO6kpk2bIrb9q5II4kSwJ1DqF
0+RP9UsM5DCdhSZgKu1UZZJkAoDrVzagoCZ8zU81GDXcV57hWpMPaqSLrER91AjT
w85p246dXQ4BlsMHMyGsc7kNH5UnE6W3dVpDcikA4LVYpejErFP3NrPvBy8QK6Ef
r2unk77F20fp9UkLIJi8LO70yR1HqrOcmwjgKqb56h/VkteJL2FW4kpqZNBpbqHJ
V686geF47I2w1xwdgzISw4H6klt1uSVGfvzYr041pi0yBbdfUkJ+gAQXD6mQurPu
XDIwM2y6RSeEcE0y+XkaNPHymNkAUtemoR6fVikWBtDmqKvZ2HId4jGN8GUNE+hF
lIZXFySwPRmMlwYCfVj6i6FqsjxbFRJDieRHh20L5ZiC7jbLQ0LGV8mDGTg/Wzfe
xHXAl1stFvNHiSRRi79YdipsD37exE265/7nkxg2jRIs2OQIu8LquE51vn6FXEnt
OuDY0ic7bpvtVJDz75FDfN26/SYdb3BL+u5J34jFyI05oS/v85MA6VNW8mjGbWDY
KrMMelFhLdWMpBd4FOGoMHkzLdiCbRFmTaB0EDRy+VDjivA+vu7MINwuE7+PfLiY
PyV3darWpoEz2SpFOOBx6UO3lhPT9ESoyc439MOf+KRcE+WKoF8H1FdlatA9bWfR
XNlnHxNmgerhaNi5EWhVUicJcnjfy1fKknUrGJys7XndMkRcjMshGTbtHBUvtlUl
n6lOkvPktYMudUWrwQarjQo4sMRkseJaE/Th791poc86ytNLoE64QfJNuQCtZ1s0
keLe4AlqgVWpufPU+ujpZ+YFQYq4QBhEGrbV9zwR79ElW7ztZnkyNxBaFoQcLS0m
l9vSEnvOP5VrJ/jaoQsT6JqOIanpRNxikbIHRm2JmpS8l5vp3As4II2C9PU5idzU
McROfsZMz1JBZFA+KiTX3MCjXj4yhYDimu7gR92W6ooGz4pZMWPBXJE70dgTiFAT
PU/TJFrJ3olR7KFGA5DSbLgqeUu0drME1w4gJoN7aLZkV982QGGNhNgqKV5cUhzc
8crJnVMlle+4SuYpYqc5vR/A8SF1QVzmpOLZHo+eRq7AFHTIGIqp+5qVe5OYrffu
c2Z/731LPFW1iiUjVL9ySsZsUNDgGrnua9BxDK+n6qLPixLEZ6w9c1gZVsPIbaR8
ftoJBhzzf4e192yaZBUeUVWGpfsDS2WThvSik8FmBZNHbdNY4M1VAmXbVzsJgzTU
eZP1ibYU+TmIbKWnbK0hep/PFqZTkpJ8LvPfBrr/6ra2G2HSGInRHHkmMlxS4g/k
4Ivg+WA/zzQcvVpq+Rs+rPDUHrtaym9EFZZiRhiG9f2X+CvYdZHVnxf5oW0Vhnhg
I2iYyBu6fCuKm2sm6taXy+SjXnlAtSUk6pvdn3kJWFBHIg4CGrVAcPTIFhHexRwB
DfRX/LT0q7JlBzTnbzA/WFF7TqYLpl8d13kSU0pUMeBcRkOq0WQTjc/PJyU1qsCA
x8awyaGyr09gDEDVhw9dc+k9hrlhwgkN3MW2qrudUeV63xe0m/2XPrpDg7V9Gao6
6ttVHqVMEPtnp02LeA6mUZkFNvhtVh8QshGScIQ/zJSjx9nheq9z3m2DDFeer9mL
XeG7DSJYdsJx5Vydmewq25Sn9dGRiUjIf7uaRvxArWh2h/BsHoa8IUNLRkaM0j2I
522zyUwcg9H0wK/RPlf3xH9zG2EG2TozR/sWJhWvkgflkTEmVNXh+WPWs+1yKL33
gTbvriyODCWYAHtJRDGqjLnBHUS8DYAR+QHWeD1no9FZs/Hn4S0qfJ55kVRt8YSR
rp+uUY7HC2dX4lbm9LtnGzv6ixNX8XqbJqkLPCpcS7vqJHpq4DSPutLG49AOQNbR
78AtwLf8eNZKWQkdW4mMEPjnI4PkUKY8PG9avLzK+nYYeVCpyjy3/pG5S2ykZvgj
jhRM768RKaj0SWWFcinbq6qhPSTROqjSMn/ebpIdFrgHic1X62fidUQJAQJDLFFV
D0eICVQK53B/itFud1vOoiLvmEezWGHsu2pHcgHDbn2gKBag8eTA8MBRcfMX1Yr3
j0zTjNq9DPGQ7+XoGTclwRtS6AVwJ93Sq06NMxGSXuBAi1VprJvhMhE1NdtVVzgi
KpnJlRPyizcTjYDbRaQ02fjtrc+JAUoIjdU6E6M2soglcwFo9KZ12iP7cJOAGXvn
EZWMdDV8FtEhkMatc7RNj0MiAPMLS6j36ciSebN2MssDnD6fFerNVkPahfi3mgZu
PvJJn75LxqwCB1unXmJiee7Lw5glUEoy7VnkkF87voElXHc1WKuOX6SBa+1nBOXB
JcEvv3aPPkrYjqQ3lzjhdKHU7EgmbX1ceHNtWLfbp/NkuYZqebdhRWZt6S/ITH7/
nPlgfzapS9Jl9yqKI+j/3aOEw1/HtaRLAA2rFilAjr7xj42mkt4425S+UiiozwfP
y9usAZ3Xz4m2zDRzjjC47LYxvO7L0ggsZ3srTxn/Bkez1s54fhZc50BqCqqqS59z
sHtx7GHj2UgJu/O3oklj/HzCr1ljTtEC85giZWwAfjM4yiOBpb/FlX/h0A0zGr7h
kilH34aiN/QGcHg3avCpxTiFfwFv2fkkLHaeF60U/IH8vnok3UAEeFeJThrMyIWz
bWt7+62KE6I+ZRd0QkXsTkY0LwN/2SJvTF7NDYebVeKeX7d2CPU5OWdoyAw7nhUg
dj1MZI2MFQEb8+qISC9x2g9eriTKF4MfFFwIvZ/R9/RLaAVLW44JNQUcm1COb0D5
Pr6uvufqeykkjgAadYBGuKw7mCS3MYNT5ss5tskzvUdjB8fcXun0pn8WvHe3lBcn
algxvxM2wSfEguPn+yiIQ2XkQnAPL8dmHGSF7yW2d/8L/6QhoC4jfkABmtFWFNVn
0S1n2g9W/HFOGKfKY+h/kfZiibDLGiME/WoLkFGdKj5nSrW5cqWx3VhxUDfoW7xi
HTNdW90Q6EdavMCtLe6D/xlK7DzBOMnekkx+Rl863mQsIB/cs0yd7AtaQj5zgEEb
0b3qzSV+OovCjwXNQXsKZW+TDQqBG0JAoF9eKZpNEyoZTCcH6lStRyajCdqnButT
5cJdsONrmno+4ayI7+9DCR4dOpIbEdWsQ4NQP4FLkVVP8NJQQzjE61BvJdamXDZX
obItYm/S0gtnLkRvgtWPlPq6gjuQi5Bf+cZW+h+iBgEHl0VtqOJR48o4y2idIHsp
9m5cFYV6wkWpP1Azc5BES0Bt9Tjr5Mkc5EmUzaaYhEmXC2QivVYmz/Q3fQ+SE0Rd
G7XpKLXhYI20NOJF4HPUoN0NhZpdWJ+VNyrgT1vZG+tibfZWgUzdoZy0gSG92YiW
EKShEDD2V+jGQVFgkDqFbOmKwHAMTjmA9NV/m2J2/tvhoIHL9Eg0RbBUHXZbK992
+ffqlY3V6Z3l4xIDZDZPtLxakG2UPARLQJVMW8pPMcdU3i03skOse4sZeJKIItKW
Q06YEkKs4SXkdF75Rc0lYXhUPUjqFo8sTSza5E84dFt6S5PIROGyZX2xQiHRial4
1VybTwExBzSGFJ2IBbC+JdrNDf5Spk0TJ39rZCSTi6jpWGL+iMmBavn8bpB+sAIL
dYDe9VXWDytgo5ZK0jpZrDF+e7jJyfFLbz62Rw/u5zpesGg3QsBOvGDng9brTtK3
GoKPlU/zUVt9GmQmw1NLvtO1U6RtnXuB2+PwhHiEHKR35pYz27SiF7+odXjMAwLH
4Q5bRaGSMBcjZArRbVIC1cXyVJ0FnJNO9XFSYk7qtzX4U0/b01/KD54rN4QimX+c
DgK2Ixe2v0AcPRW+UoGjzf8f088jXqHJxa+7azzlZ7HPYjp5ZsVERrs6+n9fd1cL
rGyD8MzvBd0nAnnWRG8bMqLhxhGukO4aIQ+VO8UBH9HsshTOiYuAzzr5pTPWcueb
VfulRG5Vt8jdNL+LkEZYmg1etLdF2wlOVKsMO2S0MEFmMXwPGJihc618/Wv8ttW2
vGFyoP8rP+cp24FBFPLNQi72673KTIX+7YtqOCnEaaV2vv+GhepAhvPPl3yvoMnq
y3MJdkQzP1QMvdZX0wh5JAM8udgtakBmyO2aKKekFBu+nP9zp/oRdQTp6zzt4nSe
zTKlo7l0XU6fIncJzgaff8HnMlAkbtZujmKv4vWlIkt/pRDjF8F4jYf9AC/TIviK
GYc8epMN4BPZpWA/lM/N9+BLDDm36rEHjqEUeBXQVuDORHL7cTdYmnWJPVZdbeT+
a9oo2CUAOt/R3AiyfnsQ6UJDFHd52byRmm3q7SbMWYbm5BJXlWRJDu2Ga75XgCGm
RqNeMT3HkJu3bNpBAgLpwjy8scwYr5gpOjuvnanCvYUdUQvfM9zaYCNkK2FNmiXR
nLe2jnZiwEuHHLOShps4FiSb0o/DGJRoc7YNrYvfg3pKoz/vs0dhORC/XA3g4h1D
KUCKU7SBq417Wr3O6CAAUiJOrIH/oWr/4JOfms/yrScw/J6PCOAKdO5bfI0u9aGY
rdmPKg1Lb38sECeqd9COjvvhrS8iuDkfoovHWQMKE+JSxXRL4Ujdrsk4FNUtDDzg
y07BZq2U3nGJgu+O58ArnB7zj/T4Hdq0pG9kY6TIre9kS/RWifBqayu0u4gsbDif
aPVB3wR+IBBhcAp0JzZdwe478mXHpitaA5gtBAb6EJadBRE3VCTwAs9uhhQwKXlG
2i4QPOlFr+fCVVyig70LodgJVofrnIhaHvp66BM5eoxRuXTnJnqGRdb478XWkrBa
Yt0Rp2TuizW4sM/B7WCU1HdXWW5XZkXyqSW/zPXr+PPkVybhkPQo+bPAIihJvAdD
HemxDQyawxoLqcn6L+c93qtxz5OqnaTRceAtrd0ZYFD/vTf6dv/6rlMecGX6nekD
5g/dbJth/iWK4KszQ5zQcjVW/IUBcSVQR5m5IaaOEo+DESKFXf7FQlBC7E4zKcNe
ZO5r9ZZ6CId1ayGbBjsthByezB9EADEK61b98TBprDA/F1gXpQ34Q1cm3xujyeku
PqhWc//J2cre6N4kCgAPKiLhVh7Xfx9qUTLQH5MssBymRs9vr5N6IiBaOyRi6x9Q
EcuWrIuvVkz8ln6I6X/myjeGv2IrLOE4kRmKID2o0R0wfzw+EWF2MRKodwr8RrnP
KAuZusL0WeaSK5Vgnqw4a1rqPgP26vtsw341AKeQ7H1AqQ1+v46DVHC5OjAnf9u9
44jNwvrJBncLzo6I9Iha5rApTENqMgH2trwBQ6TnDD3+uevfZNiayATm0tAO/d8m
MAgAIMoZT8wSDzG0vH3wkUwqAk+X+CQh2GgOZR9LE+cWjq7ATZuvHk3sVmEsGKR7
lYfgTDer77+zGmJa290CV4R2CWoUNYMSrZe5QvzuB1v5z5KSTNwf8VO8UKEW0HbJ
gIp6+tsU8BG0N7t/vtd65WQDIUB1W1t67AuTvSQJLvzYeOsFWbGDMNDbLdv9PvEY
EKxFr5Q1p1TApgm/vkoCrTBZ/5fs7FA4FpljkSUtMkOmF7snXdwvORHsw2ilXwfG
pIHnB/1eUYMNj6WyqPQCWLMHkgixYn8+u2yEFA6wuARW6+4credaG6HrKSiPB7IA
qAZX6xsawt0hnvOqO3SrolXHlLNaQiSqCUKoUyYCnIEqscNAo1KtUALUZyjjE2I7
JD8BqijbO5vzB3VH6mXJraXxB3J8gdtKL3g0jP/N5v/jW1fJyVIxazbr3MSEaii5
B8HlMFslRByvRA7hEIVGr3Z0lPoNJo5L5sP0RmGW+SIuFs3XKcjYe+l3W0B9h9BH
pYVhP08wiy0xisY/og6QbmBkTE+F4s3OMtO9mxgmSaIcsypRwFCL/nCVVKb3npy9
Qd7OhVzJ6C2SH71Q50x3q1OTVEcNbBgQKYAhWtch4I9rj1tX3q/gHdvwW1B+BtmM
0EVhwkbJFhFCCm7xRr0DFF0M2NLrLsn1UpCrqUUDmdieBw115v4NG0/vBajyJ7wY
F6MYGtsfKpwiW8G03qZXRrCBDfgp8YUjV3Q8pps1Dya4aBh8zhEJyb+r9QKerJsV
efbBWfCHITkFDurSRgA3h95q73VpTfm35B3UBwkkaIz6SxjyPEDWeTfB1sleX/7b
0uK7eTA1E4kn7hwKz+Ikw0VglJiY0hF1ybmRmxhIk5uv7g3NUIkhu3XYVbL6t9a9
h7FULJ6Owk+iFGV1Tj2Y4dhZNZzlaT23D4xdIF76fZPHE9Zhi7YYkTIjt8hF129g
IfvHHNbe+AUeJITutKMrxwFCHFowFQxAaa1vFxIHmzShv1vwLR22pbFPeCmN25Wn
G962oWeyNlRoj18uTTm1Jvvbpm7GWEOZ7mVMWtWyvEeGCv5WgxWjGfiL1Ztb4QHc
kIqZmhYKc4v6y5NYjGk25W0GY8hW36VGTG184CtjSn4fdn5SY9lKyFFGS+4Pqx7u
+Z8x5Fa5AyYsCiuxM9cUe8ejkOyxtl1BK0qfiI4KIbRPoQCU/XaTy1T4bRH3QPjP
X99dR9PBlBC7nr5Ogd3L/+kcqjS0kHx39IOHVroI6OdEHzHrqbVH9j4sxMcyrDtZ
k1ZYXnst3WcuTawWdAbw8qUkwAQHg3m+yu43WhyyWsOdZHmcLDHI8EreOwum4aG2
T/dQDLVcPi24wO4fdDd43LyeEV5lfRAytY/QsAThiiM6fJleXNXdbPWKnktv28dn
HaEXf+IsRCbuYv9wcYsa45OiU5oECVWYmYDbuZD461NerNCoH4ompBAexisHmQGf
n3CZLVJ6EGc1TL2YKHh8c3p8aOrRKu6qcCI135RDbWeqUs8DF8XwNITPDiLHZ3Yh
kOzUp4PQ/yvuj54OUF8S5iqpHyzpLClIcJP1a/kJQrKKiqFTHVTENygOYDZYV+Lh
TIyWjyTYtUr34RQjYHbVWoFBCOeaQEGYCNMKztDGtWbog2RLAP72T2R0UtW7KK9e
UjL3Dy3QRIVSObJChfgjaaxEOHdMzyy6KRErDBvyGNtVgT/+8zOKZh3hUEDeLLmf
g1xX7LAPiyM44FVwMp00JNE6tuYtavJIF6zbXEywZ7gZeXfZB4Q1auXYVRS18HEF
ewEnmq8dM3XKKPN6urkjWrb0RvyKeq4mG6IiW5uOPdDDve0Hv4QuvoW5zveH2OfI
gDMzs1U79yzP88su3eTQ9IfW/+XE1kpAeOgVDEKVrP6jTcm9N1cfyUv5N6RbeP1m
65i5unVt7NuVmLEojcwQcEG1Katn/SGJctPAV8HP/BSrZnJOSRHS/vySyCPNODN7
F+acegXpKn2gmZlBjgCZNSsD+odL/2buZ+uc7FX4gStUNqCfnnbyhaxPwLHs/HGS
rW54PReWLiRM6xAvYvzpWlp78oR0T8LvSZS6RtCGKy9nMtM9MiJOoHEmzK21piXY
Utr8CqKmQIDzxWC5D/QwSsDP5isodtHnSDd4Or/XOjwWA0u+0HQFwe0czI+NI696
8GeqI0UOIAtaqjcQFpkDgAx1euW4KcxwOQhBzp8hBvXyE0M7ZlznXfYCVfeBrbTL
9ypqWHCWErF9zphEvU1Xh0wtCFp3tW27XUdsDR/mD8vD5kNJ5ua6vER0ip/r1f4o
qerobdg51XhQvfkPzKdih5maT6rtgufZGhBbBCJUgLcW7kO3cEm9l/1nPEEwwtef
Roa+MH6OsB1ZFSasBUTmv2goCByTetXktfjsgKwXvTnO6ltVI48rN6ALsVn/AgMX
Khh/0pkUn3s1b2LKzOKWRUtAyMAB2bClZcEq3dS4dDKB1lkhsmSXevCmC8poFUdV
fyeqgLA8dD812ki0pzNihDVRMliVzujpPehZ6hUzCPcFayJJRds0nqRbPxKS5IHc
kklIjC3kwKIDrwh7F5O6sgxw7aUPjsRGyxaJ5oGO5Y22iv17HIDhM8QFsEXTPz3P
24pCAW2n4Od7zFcjwjTY++zR6XwLk5r+FtCRJyZVoxvKjeCP0c8NWmPQa5gOFzFv
ju7tm6GEvbCZtZn92hTWZYuNgKJtGIBwujDr4M+JVLZRBRlbXHcG+/rOzzzzSqdR
tL8llYPEn2gf5/5UU5pMP8HJqfXdQVjbOu2n3XKtkpzBSq3C/qBv8tiipggx/Onh
ivKGs4gDtzT55qybHHuGMUwGczpqKPxP4dNOOvFJ5k9RrGxsx4PKLVjPKNlqPecB
gG7nV8UlZQbh9Gkb4DGkTAdXp+t6lTw6AxOmFIMQnBiif8bRr+TCEqB0qzyBlE1z
X2YsrcFIqzn+q7f/fxo01ZP8PznbA35+UB/7aG/+r6w3Esm9aeew4hOrriuTXEqg
kMaBdNZcxoWzHveZmhR+nAW3q9zYLZ9c1fAvBz0bQFexlWU6Dmcfojgw90f2QD6r
OJfcgKvxOasefBVsvxED0ueOjYltrKDkdtKOfCIhjbJN0yYewBN/ahXVSLquXz2D
E47JpAFLo4WlDxf2yQz7qKdn2DxqG01e8CfIOItlmBW/g58fiAmCD7PSTrQHKD3q
0PlpAt5N90B/uM1UZ8Pb1PFOuo+sQSVIAyX6GiOatJ1SwfNi0T7RXh2OE4n1P+GN
sE3KzCQpU71CugIKCbu0uPLmX9jPfQDp/l9AR/V5fa2fB1C7hyQiC0ag6U8lkXRC
8dmPCAW5S/jE2LXmdHsZyDKVtblE/SLOIZBHRSB2c4HJK4R+t2kCses/ivpORx/3
A60N8BWZwgxd666q9U6LAHt/9mVB8TZanDe0fkghI3gvtQzFkpsPiNloGSCTtT5/
MjDXJLqIt6ekFMEdwF3ImQJ2eTGs3BsdPSqK+yZjGq/B21/yXnUTsGjk9imDwQ7z
DBxhdllm9YYFqoUO02fFyfSEHjVciTvBGDbbOPeQhdb092bKvMg6njXh18KmoTrQ
ZLHSB+NmNngECttEA+xs4+QLIP8iZ31THi4x7JcUDtaOwNrlgYPIzMdNUyq31Nbe
3eIMvNp+IC9adQq3qx3U1U1YgFvqc+9MRGdbbXK4jOiKa5bfFABx8CDCkjiat6lj
z3iWaU0A4z9fp0IG0KamoTVNEd6w8sstpG75SIKkswmmJY1yVCPK1IyKUStHiDrY
y/vt5E+JWBvk+GxJ5EVEs7XtYPcmpxfUQOf+4xobhAqaUg5buOgx9V72hyBs+EG2
ekAA0mhOlTR3Zz1uYDUUU7NfZ0bE84LWhyUsW//f9B7pcS3ONxAjFRFEq4o+ibr9
gg4GnxEHB0o+diSzzcxhLoHtBg9UVkr9B6gCiPaGrKPFkKojhTCPm3I8pvV05SKa
UwLZfBMXH4xyo0BEQ0wj9ivi3q0fH67anYyeez+DJO3o0+PEo45CIYgIVIVmIiUr
ZOLRlwIBQiNPTUcjLWyeJduOizqRXRbm6SzzTh7dXe+Jco4l498N1/cjf+2A+xcM
zeassKVYbbtXZUgmgBvl9TJxG+vHQqNwvDCDSHLgYLMR+8KL7WtAGWrVHUsL0w4S
eQ6aFEX/wFPbvNBRKDSYp3u9MaqXrCWAiqIgZQRRQNQw/PK9Lu4Atfs+Rm1tm3FM
tHPet58gZwv26Za9UcSWri8I8N/uJzKCcRVqgZjlctDo2sd6mbKf+es13doM2MBC
d0C5VjdBOzWUQlSzDglGmoL5bIQKBXi5dqg2YepuWzC5vhTcjv79CKpjWlGio79R
JBl1KZe5dABpnNfDqPtBke9m7tDSSlwZaq/1R0VAFLecJxoJYDHB+52VjEwbwLUx
Oe6pZbVbXBwT6QN3y7b0A+DBZzDxQfhPxVHD708Je+LJFjqS+mxC8jIslE4wHh3i
8KiJvhOsiqfjVkK0vjbA3PforOqXCsl3gCvnsvdQtca2oipOptrtkmkN0BlKTYRh
/CONClPoeYUe8izzSeiJpMJkjvFketQl2om7AJdyykPNuJYxRrxocs2Ufg36Hm4a
nvwNNZf62pCuk0ZMMgu8ZyPbrD90Z1pjKtpc4eUgrUWAB1WbyzpGODt9rjR/J2pP
mvkiBr0bDjVQtjxhs+e06jEFlnaVUXwBgJWu2CEDCtrYfK3Nz8+jHEFr4mBmhl5K
RhLV2+GuimdMX401PGQK6OV8rooK4QIEw/Y68Y+eob1x9zbL6Eq4ip+l55p4vJmf
bhCFIvTYaF5dh8W33zrKRHaj7Bjo7OkedJSNp0zYd4R6In/kc50PpzgXXhdbRJHz
EnVO5UbAcui0XRYOvh194pfBbMyvCM9c6qNyFDmQfvRU5o/AGKr9LakwWhnja/eW
36vFLCiPMzRsSTmMxSxc64k0pzH5rtRsYX2I1z15c234MSM7XQhr4HpWzteyuQur
J39ZzynZsIKB06N36jExgui1ilvAMsHF9rEOmb1lktQTt5uXnGFginZX82kWJZun
9GJflAZlaB6eItKdjm4U/sdiGcDV5VcMv5/aera6ONVu4r+iB5VibScZF2HYNCDf
Z3LAWsfjz1zLLkQnK0pHyYgwbcR/ARt4dUjdGI5A5QUlMWsjf6fwrM7Gfj0FLZwt
UxrT7ffMoR/d//WXo1a9p2JJfMdbqAMVMAfHWgAQ6RyA6myxORb+qG6RzhTFrvUO
6419MsjcdttjhGpBR/F4MCLiF0Rp87BmYjlMGvYOGIZd4p+ymSd1gxv/TibtILlh
LieCtdJjTYZV3u7GoIwHKjErS+A9bGqA7Kq2XHKHbH+ljEQQ+90eJkyAsX9jTc+J
LjKNJTrdjwJbNuC+1GiqFaKcgMcUjoPAtdN+JzvkZ+qMG9Eu7Ry5xkVVmTYkqMDs
Hs3y4/q/7/xOg80FE2u/2hXNaYQ8s+GBwY1H/TcHRtF6HT6ibXmZza330bzULC3L
ZJwnuD3u4WpBosqQrOQygj0tHpZEKAhcDJg1bEwlGDP3/tnGdEzmTnK/A7oc0606
FxdlHwTUc5TBZPjqsbnRBlBawC48tkcWlJ0RNRNRZY+62KPc3dxAiOhbpdLnKICK
sHqSYpvzlwlfnpql3iGrj5AsfY0fr7v64Utl/d1MKwK1KSk/+1MhsisILWOwmHiG
WS/U1+vTNyqD31obKHBZd64TBmfSLZ5hqBsAo6DKvYSxTtr+LVN3LXfQj2BJ8P/L
0BNnfgHpgt+xuSneLzaNDYjECNgu4zJZ+BMB/GvUC9VxW3ZCOrBxGjJEK6jv6wP/
FU194RHJB7BxNSkY3uCRJFAxSCV0+3nOZYroSb+6jr1m+HUKGAIubjtm78W1C2y0
kNQRX1SiMYdnFuZ2pCcgrdFVVKLD+q5d0ZJ3lifEugMlrC9GiBa0Ms7cq3YG+Xzb
a2XnPR54H3bVK9LdQmpDq2o7cfWG9LTY0lJDkpC9LFKjuVR58gkUTxxsQuzIKDpX
LKkZNUAZwc1+W375htjKQs7mGeZKbPDvm5zWPKrjN8HDwhXlKKCtc4R/k8OBGm5V
TENN2xsXm8W5/OVRIEYoMFRYIb5CWouvtGCMbbHXCnrtncLs4XIPVFe9Wg/p7L0B
voxb4m4QJPaH8mN+Qu7k3OdNqLHC9x8K/BD5ECS+M5H6c3F9MO3wMfm5UKLEoRwh
SfuifMIwfvxspyGnW9QOCMur09l/r99u21C04QIGLegQgvK3wDLzekAowMwnav1O
zMZ/rC8OH46JxGHjLAQdLKd3kiWqXKvLTKcobdUkU705ZED1+He49kPiTPsGu0DD
/DC/NvfOHb8FsRcjCkIczQMyI/nF7jctrfJ2kiSV7AGIzdHyqJ6EQAigSLxqo7Bq
h2E2E6WxBwwhKf5dEfnsxRbKZd0P/a/mAiA59G/RJy4ToHL2W1Ugqsi8AtFWJzRe
8UqFGBjkQYrhBKJScpVjziE8WkjAhJtcYuN2gSxqoBiin/MEW3EpIP4pFD34L4f3
/5jToAvWixM0M0Mh08U7hvly5jsPQpFybt98kYcnujJRjV+AeRoQM6X72mKd4iZU
rVVmP4RPj8fvxzeoc931KQbVc94Urpf8AjUTl2MLpWeWNWwOIxdNNlnmzkIeOPz3
jSH7u/hlgITfzOQiGiAefmJCbqAfHrwWxxCYS6AxhsAVl8xxp9uNoZLcrKFdRvaC
OvDFigy14IQA5TYOfR/cRrznavky7Mjf8mbWnnt7Xgu3KZtdx5sgXKeqxog9sqDF
6O6mOiY26NxxpYcBZhAqKHl7SNfzjHySh0zq6HL8FS1oR2kxhNWe3aGQI3W2qOoR
1i6E8HKH+CWlSROKoZIqqdjII8laAd0r1QsHTHDLAptD140Ew+/QturIWlpA84iU
HpdxcN3tnw+a2H3qzbac3iVXGB6789XZq4XhPudXlaCyX5qHOaB7j4qlhT89rlyF
seKeHwp1u9iNcUj8kR7a5ifY1V2jzxPLTx/4YTdqhTOv62ZCOHIB4j3iApuX+92t
jUkaJPiEY6pg4hb1yzH/lSE8d7AG2w/tUJ/ULwUhCFn9tJAIS0+L4DpZWnZe/d7U
1SlbmejlAbarTu1TRqGGLRoak5ER0iTM+5rt0EfEl01eSQVE/P9EMR27pcdYu8+1
kxbkU+Vm3qC0pWBZf/Ho8LHXXEFsHLh1gjyQbF9LuO81vYgrLvp0hUvvCY5rh4m7
8VT12ytTamVQQYf01rr1Gftp4zJAeG0mqwOpGtukMl9k6qJpifMo16/AE8Nej2Eq
Sbi+Gei2fHGzAtBrADYOTP85KgQtl0toitWXZ1/XpQCvpCYvXylUxE6mF4HWR1tk
pLxeJkjTt/72s2r6aFaHWV91KmEKWdZji6nvxfn1yaIc4sutIVoCeodyJnZZeCAM
eVq3kse75Qf2qhs3UAgJP1GcPzPsBM9JyKgKvRCi0sc7eAfbFqFTN69qr+3nl/Xn
S/Sp0p1P395R9x5eomPiW/Hog5BG4UVgNSSyxEj59eCfAuhWudCLLaATxpFHsMGs
Oibw1Gll8EWaDzIGF9wi8E6FrqbsruF4EP60DItqzWKBkzPbggHjbl0FILBHTcGR
6yxa9yDbI0fFClJj6AMhP5a5OlEpMqtkiXxCZAMqQC643T5f2Y1/b5eMoJ7cdcbK
5tbvCwwZEyVNBDzxmm57ZfN1RCGMIjFpM8bnkaWPEZzuFqf0asyore2NG3gpQW+l
05liUJgmIgBe7wArjuOXbXB57Tjfz2v93ORvLVf7YPszeFUnukTCnFMqubOR6KdZ
xuSCKpMuKrRcBSEYS8fK6Z6yqlmo8Rj4iqdKWr+7o+FKz2ge9JZKd3/4lNYGrNq9
AEeCBzSsC04cu7OBHdPvESAA3bhO2O5UIfo5UOQyW/VqGlltj/Zfm5WthZS06FaF
bGQOWYQ9nyPEGX//qX22U00xHG/dJ+EwktYO3xsfqrzg4ms05oNz4PegwZDxOwLg
AYyTLy/nHUOH/NaPRa7W2eAWMxzRmaQ2GeBVMuOITr0ObP6CulwR4ylX9ywbUhY/
DYrMplHuwyC/TgBTxbfcKsJYILV+QdybYLmtvthfOjsmoUG1Ni1W9kNEJSOFpeJg
93xsAGcC91uk097NyZPFbKsOwc3jDcUURel8cD1rXZum+7obNsWjxlcBt6qzEg6U
rmkb08I6THYbdWwoXZnDO67A7i/W5GKgeV6yI5r7Cxr0JmvXINALMrn384F06Fj8
KhFeo7rKGL7ui0SXPsBVH1y1MrEZoC1pIkC3UBat9YtsLVHz5uhfYKkz9y/X3sJs
HktuKloV7m3PxhwMcowqu/iBD6iRCdJTs/naFplcmDASyeyb5H0MlTUX/BEIg8eQ
MlHm8nIJPfFajXvkNvG4aSrp7qDEhKYSU9QHBylY3rnNPUN9GACCRJ6lXcdb5Xcl
BOtSUG0KLklk9YLffhluXk5pz6l10WxcrgOtGKMlIS+nXrj+0Lq1RBrm6ZZKc5w3
/QOzquy/pLb07X7lzJHOXwafYJCYEEGLoP87ukqZf7gedNCdS0PPp8fRWuo4p16i
s4AWHD5hqXGzITn2FAsgeguPss4C/n+yZLCEhpZZs84iv9Fn+JRkaP3CicFnDQUO
/vUWfg71w58c9u8DheUHCVnQ1SL7z1guuFxeNWWWPSMaFDRkZAh0v2PrJNNbRdxp
v+VZFNPLSnikyfZHZZxm1vRNVB94K1DrIBOaeXN+zUXemjQeU7jvnvhHcdbrTqqg
Dfv1oPjaU5Sft11uH8Koc4qgNn2avfVxziR4BryqH09hSDtceTZ/O4UZf82kr8F5
tkdoNEGrDqma/9j7K9Pkg69aWLwkpVhVomv5qcKEqNaMoWsYwN0zWPWlQRprXFlS
wYJwtanXV0kU1ZtVp7hrTmeWdLJCWDmdCu6v3p/N1D8yAQ3hFy0222BwZCkecd+z
lvgr2YDhT2L2K5d3h7Iovwb3nELoUiZ5nt0i09sxl4FerMRP42sGcROQR86Xe+J7
6re6dfaiQWXEMOL1PoaXy3eF/cnSs0D3CgqoFNmhk9qzIQkGbSTmhxTiZRHihz+l
BDbA0liHFmSkCWTkD+J4MK7JCJfURMc037lZ/Ar8WjAA92zjRx3lpV6l+3Wm0OXK
JQX7hFN3ztHy/6iVxwmfL2gKXO+llh+CPqeKCnpXDLktfETke/tan3IpI0fblEZo
/WI5MkUrH4ZdXmKi0ei+IkRgobYiNp4hQr+ZT1ZaxymPl9zA2MyRCSXMfdUHu1kH
8lxCp7ynL1vAm53lnpEF6xr7j1H3Ih9qTQ2XIsg5r5xxcoaA+tfo5/+CMAKBCpCI
VwdugH8Q3rWtzlMVMJKpbw3j/tYtD8T1ZR+eS0HxWH3TbOqWWiKirAdMPA63PDrH
U/LbsvUsyc+c28ZVIsxrEgOdZtsnBxMfkBEoytp9+7rjbMjZRY7FhjX+vNDMiSqJ
jJz3psD46shEXr5b71eGlQsu5LeYbAMb+vhYmVd0izFLNhAZ2ib7KOaNff0E0WGK
poDWYvOR2n4Pw9U9R6Q2OJQe4vpnQmcw3ggRfQKRcctJbYxMePhGYRaZ0ivbUFuC
xw41TaXAU1DcsIVAUNPOl5h94rB/MghrLgbZgqi/x1yiOvhh0ouaPK4ugLjH2NKh
T54WdydEx+Woe/zIYNHg880u6MI9LaKzvCYUgVoCer6SE+AaCOtq/jF89lk83wk8
YiHF1UHnG7mC3W1Z6kkCf3VzHH2Qnt30/DYMgTrDZWNu/V7rlJ91UXVZjta+bRET
k56rjrO4tAFXoUswi+SZE3Ic4mR8Xa6J86QlqvrEGdELf7xtZRYvquDCLa4rWc+N
8ISN1g5O9BJFoOmbpK0RHpTHdgMSjUha+RXhRFCqKlSM3cK2LoV114iHHM9wTXV0
Ox08XXmlm0k49G12J8qXBCkpZlrabX8xbNusuP9susBdPYdQBLHdxL0Dh0fEZu+p
5dLO5CzcblcO4zw68r66yJA9zH7doiJ/HASC1Gq7SFluaz1u7cAh+BnjP9bPUzsy
3vDw76Vl88xTvuUyJq5tuoHvpjwo9WSXUGab0GgIUPmvkAiSEuK9F3HpDV7MNxc9
gBedfNM+r76ju5LVUeO4oSLUA9gKokiFCTGXVAJAWdk6WIq7sSa8AqSrO9vSMuw9
dZROKHsQQNPd85MuAkfUO8jhRxNtNdLFU9xzDKcYof+qHRnaT6usTwDL4utftFnx
iRnPDdgOuUchchSHDvLet2F6OzposWi4dqNMDNcF04DtcCF0pHB5jwLayA3kZVzU
JAb6y6iTFObgxKf+i2UT+nGOxq0+mnmEUYgvZibGVUqmQEDDuN0TZj2G6efQOrHH
dLz/sBY3/YfmeYLWvvAhSR29XogyR5sC0NDfEpmjJEmXAQLTv0Y+YYYcvcXQy0Ru
Ri4Tw9KVKEwGIVspqPxPgRMq1Y1hAXYzXy2eKzcjEkmSqfwsjWUe8KBZX3NF50y7
DxEkBUGwetTBsumYZePwkR280WHLHfVmf4OZhKq7c5Bvuw16P/D8VB3N9e7WymK4
P324812zxXvZHbbdO1l3KJHU6kFzoROtaGcEZ5yFXQisQ7sF37szI9E2RJYewWTf
X5S06apoDGoN4v4W7YfFO7MjwMrP+0UyKkP10JPHzBuutyLWRQGtlCF8x6PsTL6m
taHgBcsbwAbxsLMWdQ7MiaDyu/q8EWpi4nSmgD5KwCgTWrFPiyfci/0qBWCcAQpl
hyLcTT0/JYh+kn02H4NYjoxWFRfN84XT+wno8HU9hEW/CMwMon1GVP7UXbrBhi4q
68c95hGo4hSDilvVpnRfoLoSfYEo0BLay8Ld4pMGPLH88icgJYmi9sA3xUA9dfiC
tyvuyyyvo7N8jY3B+A97nisyNtBVEqhDpDuMeymd0x+JgIwrtVlV0LScO7Hr5yiu
iVxjQcP0BIkBSPC632h14BZvyGNGnaNk+AZZcoQJAfNW1ijBabl89NGoWQDFIt20
AOLuovZ/gWrloJJV37gDxCYbuQFOuOC87qBGR78dv8YDWWCVwaHvqpGkF89S2LSn
JFDt5do1OcW+9khJjwVGbemTH/AnXKsJWtHLdAC0RsU9B75SIPAJgY97Xu/si/3p
coqSXzu2J63qTTbK7DZ15QWMnKxUoQYEyZKrDE5+3u+pQCHBm2olus8SUuekxUQZ
G4JqQvLgt1Av+9xSSOqYSgZoHEx6oP4VGA4KUAxb1D7a3P+eYlafUuG3CAyCYrfX
+wraf9/wDnKqr1GsvUJdrUizL8Ixq8jh3BP8WETsvO5XPEPQdznEiXq5VK86pbCG
hzTHFX5dHdl3f6g+OG5zAX7FJTu/kXHgyL4jFLpg6KeFcY2BRyf9DqCdU43RXh1G
Ul4LBcB7/Hk+qi+FYE3p3TA9Cl+5UPEZpqd+9US/b/sUzUaPlUFwZIPTncjaTHJP
5s4C2sRLENWsEYspLNT7onThHSSgnVmIKbBwAng5tIN9z+RF1WnOCKYVEQlap/m+
WlBWIXFLK+brM6larorjzw6l7CYzJTzIFFvzFJMj1EClEqF5W2Nudsj9Wd/LBW9E
2nxmELxPOOK8PKD/zfnszAxVqMrVjxFYnWZNKvvevftARriWP/d8C1F69HYr+IEi
+f4SLAZh39FlIt0SLoUZuqlWMPQDL+6uXaL5q3siv1UjI6ouX+mWOweGGuweUJ0j
/Gn+9BQN5Icde8G8oPhL2wu+PVmMyhEzPL8BUwuWZUO88Cg1iI8MBc6XhHQCs3rZ
hhuj+AUBNsPMYe18TWU1yTKPsqebb6qbeS8N42QcF1nHuOQj/bAZaRNk/P/kpN26
piSTHO6r3Qg3N6h/H1GXvssmLKIlkqCOt+xJmgAH/tMfQgbFZIea8nUi0ujgSTg9
uSuAe+JBWJuy0yPRh110PkyU2IFax94OG/pSDuBHFKszfDhnaoLEZ/AYNpXHX1bc
gJeIuMS/x/zYzKvLh9qnfkuYGqWDFoftK5pdX2qFXBQGkkWVU1YPmyFN7UvcTOxV
efROmWBDc3eJiZrcRQqvrxZnJSPM3Wd95O42Z+5N0GWQbOwcH1Gfw9Sm7Oo/P7gy
hIrF0T9YRh2DQb/4KspU0IcdRrC7KNZxaQ8xHDiBk5Ab9hWu/1hW4Q+hoSxJXgiW
PsgJyq7Zcy626nrVvWRuH7QsupmTKuaGxxrgjFUkNueOWDIUTKMMBcVwUlQzKMix
9CacFb+7o4JH33rZP8hTGuiCC/KT8vjT16jrQPsn5DVIGMtTyujjxDD5bge3lwNT
4TbP71CzldhlMul91Fl4aauWH5xTox93cfCkJJoVqWXbUVjusXjR00pilr5irGHd
7fklsGEEjA+MOtNskgiJua8NLosrP+UCUDS3K7eTMO/hw+aIqE1rOeuo05hJaeIK
6xRgVChH5ov+0rtIaWJIvl7ohcN/wr6UEVrNh5EAyoHCZv9bjR4vzHhIt8gG6+D3
hoybVGAiDAGqnqxVlkcchrfXfmFgRl2rrqQw/9w7kveDKSZVjcZlH2+Oa76bJzAS
jHbLxNWM2xYAEeDbuq1kk7Fl7ae9F0+UvaWGh+DT9FnNh/U54Ca/0w6BOxKXtNxH
lNA/XCfVC/e16KrUHasUHblhNVfAkISx+ODuwyeL93z8yVXtMZzi0GVHlsCLIwx7
vQ2C1E5ffjCVhnlZVRXkValKyD/BwW+6uJIpAk3QHAzEjd96mQSulX0KLkVsGFCm
LNCeHoxCwnF8MHNzwi0eJJnoQZqfUmroEEe973vhYTTKZV8WgPLf+BX4ZyLCfxR5
mS27mzllpIzN5ihzPki24WyJdWTTC8gY5N3J9Gu9EVu6TUDudRXEDx4bfL8pmkZF
ddCXRs1jsFZYceL3PtBY5FqYYbaGA7IWQnWdk5NRwWoYIbE/yBNBcQx8pgZMqnxL
sNh/yfboYI+yki13YSIEAm+2reL4OWSi/QRowAVYgqXOsfE3s368JxSrNNC7k20j
RcM7FqlF2ngTo5cqFOaiU+ZnehEO7azlT8eWcO5A/AL6gfWPzMNjmeCUJ+dgzyhm
UoYg4Ex55v8pykDlbruaDz7atHime21elT01nAUVsAyuTMf4Z6+PuEOXS3ozAvoc
XOua5IhxZvqR8/gfzkN3oMCMNo4dGyn4dFeETfXeYM8Sj4tZ0Q9qJcrg5vm49kC/
vnM8JLdVDu0Fj3EgTAbsdP1/WgsFApoJCXuclMGxM5pWL/gNvZooX4hcObBCVchG
UyXnmY/O0hRprCZorSSIbN4HVrGGuMIu++SD/6y1Eraji7aF1sGYNNL31EzhtJVG
wVdZ+eSzmMAjZulS+hWXwuRG2ylLcg6QYqsRrIUtv9QcaEkW7QcJCeeBH3sv46q+
XBRVG416pMztkXU0+Yd6DcW4ZrOQcHiKl7RIW1xl6SVqCSOa9xbHKTV5/z3mjM3L
i7zs5wH4DetNXfejpnSKNMWk/0xSq3YcHiJ3rOFIe2JFbZE4Hbc1J/cz0ZAlS74r
PfwlZa6HaNcINcD5OGJ23KNNuKbKcVBSYTW4Wf7Rb+WeTxm+eSh5nnCzGu7I2Isk
7E+4ZG2UFwxsDayjzNe9kw8WvlXaSBidBAyiMGT7GXHbmu/H8BMELq1lrOjwMw1i
kG8hewhRQtBnOh7dafPyRZp49Yi+des1WL5hl6xC8lm02xETTZWqFNRvVpXAmOg5
I4yfFXq/xt/xUBUsiOZrUsRNGBQcgqIRvxU5KPITQ1Rq1dHiG79G358BnyaZDi7G
Y3gEL0Gx4ag7p+ICiMsq1Uea/MQnBCmEaHQN2zV+cBl3ml1W5qFYkcYNHEyWsLle
GJAEtciXPt896yCJ/pcInPRe3UO2J8IwcXDlAj28jiVrIDNwNPT9lFDk55kcDxYF
SjDK+f189EQ6EaxmPF+QyKQKXXBEvEMo0qumaAU++EXDECGIYtsIvzG+JEDQSS1N
/lp7T8XL4rv/xUyyLcnhScddr5+3++x0ck0cgKBTv1hVFuH+DZ3fKmd/tuLRkKUq
3lA+K9WlUHT9w5JuMkpqxpUW7FHgUzrE0kni0lP7zrse4qN9ztbHiF18iGVCxlqo
dUdMoh6K+63SIsiEbkL1L28DI36byBD/PyUhvxUtwNj3HKdl3ksKvbEvq9WmlaCe
onqjyTEje6riaLWYUfXJ9lwCDhLHWaMDDXehCFV0mv5a1VTKP3C/HNv4SVmPh3m5
pUfJX/0f8wLl7i4dglLeAaYmEOZQPq4XGkQndSmiPL4QDvL/jW+vnEJNPW8OFihx
0385WmyCCiQ8BT/5EbsfFoNgQ1bS4CiePtOeJympflBsB3b4siPjKiwULmUgdBeq
oGqmE6Uu38Q8pV3CEMx8cjMSWz0QfW9x8kUvw6Y6JbdIQJ31AHvwmiqhoIBY4a37
FkrovpftMNhBb1MKQVeS7IsQcrz/8o+jKa5fYTkihR9Eedea32HMdM2gOvRvwurk
HpTj4sJ3yLegc5bLUZJ//h1+L8d6wYEhh7K7F9r+CdNqPyuYFwfJQdadlbuCv5/9
EsGs3PLPRD6n3tTT9N15Op+NzgzeZpY6uCaAm+hMvEYsOCUQT3r8c5h0AJ87Hl5r
G3FHZcYSME8g6k8WfA7HseBLq+7B5nIvrqvGY6UqruAp9zPxKpAgGD/dQgoCqFOo
ufaH9kdpk7rZ7/p+M7A/59qxdLA17fLDe9POp9WknbckPWh+3OMAmjebp5urUk2H
Ylw7oYpwyOmYIrTV3oGybfJvrU3nb2JLyDqyau29WxNJQms2W7Uh0XIQXqW3Y9hg
z3OOqUQJlWMe96OUg6OC9pHWTFAKgWD/WSorcb/DNDlq+eCFtRke2v1DB6tAMjQZ
e8c0LbPUMM/iy5t3T0B6Kbx4qVqbyLkTD7muNBHJvya7qrEJ4TJn8tdwSpRi1y05
rKcSELdJKA7ioBmJn2dIl6PEZOw6I290l8ttuvxybF1436xz5ikwHxBa7tMgjVae
uHJIMTef5w4jO6GBU2sTRHYCH1AzgxWfk8vmgJPiOaM8sQUWHCi23pkWGe0QMtL6
itIBHG8l+TMjgOLNeU0EITpijw7eNrO5/DIro37qNEh/MTG0m4JxAgLO0soFc8do
OGw5FnoPgH3ycH2NhWi9QfDSlclbCmNgebkUg+5oln1i5rN7iWcmjpoHgpznIxvM
TqC191XqHab+qc8Twx74x9JP4XbzFxfPK358jlwjL/hyCo5MGfd+qyPbwlPaU+mL
HDaV55wWzyvurSZRpPkNKjoEg+dxp/uIHV+BsyzlyYRUCsnuJRauaI/SEabH7VyI
M5F899EL+h8CbYVYCsbPbMV1JW+Xy28zw3bs/k+JMUuPADOWYrNW0duATZfhwOeo
tWk5BoKlKkErob2H/XQhO4wmshDrsnbBonx0D5uJ0ppZDvieZQ0belmUkWsstSz+
nj2VWu4a6UB2r/cdAn2DglACKPqssavi3AFrjFEDmwAmQy+sM2NrFFrHEWBfnQ5T
mM0/axUilG8jM/e3X6APX5JzHlSWJ3d8d40/qFxuB9aFaVIq7F/4ilRp3+lcAK/e
/CtfQHYEfjcwTtD30qsmVSBA5MXNiHdUovomQ4xmEeinBVApZgJVB5IT4CvcqVmc
CUYj4QPgk0WOCIVDRTGA8KEKWg7Z24wDuAQqdnBgHemO7Bavy4p4S2u9zN8+Hqwv
IYy/Frt/JZuFL+2fnWiUvlg+qaQefYGRjPmk/gjluPAVePj1gjbnDnOAOTiaeaCd
fhkhSzZeL+g90t6rEIkTcMXa4MIAHCBUZ89hyFcj4Fu41NDoq1UaUydq16zNMDQY
LutZ/5KEbpOzlRmQiAxMnJnJTI8fLIXkmbJ8JG9feeAWIL09fkxzotdT9CifMEog
+mb3V1bS5OO6Hmx4wiD0qS3dJPOwwqNmNu8liyMC2jYmdpclf6q6ktfkJ28LP0+S
1x8eg/kXhRWg5e/oksjBgi0w8wnqxTFFDdCKaQzY0Xf6shUBv3o6t0kG4TSAQyX+
hpQyB85EhBjVdn7Xe1oPWleWrjlXmK9ItpRIQyuh9qDwELcE4R8+VySEUrbJhoKH
NzUwZqHYu/HJTSORJDIR458xnGFgMjilAKwNxpCcuTd8dS9mOrGhzzB8ySaPqJXI
XRFKsnmdiqQ+Ld5V6Fse0usu4+MeFe9T7CzkG7yg2Mu6ExrTJdj815lYArSOIh3R
xqElzw1aygB9gQzB8fqoi9GHoioTOlXgbT4M6/650urygNAyS5DiHafi0cKjup+z
dVD8Iz9UjqmZWzIq9o2wJKENaoDWjsmx9cAeHbP6xFEfEtA3v5H+TURSGbqZ86j0
D5AnLR4akTcRdz+YkmEJRX+QJ2lWt5lTxDocAq3LhbzY5uZ5JnJBljf3seEmg+Hq
cS0biPVpoxe9VLetS69Def/HXaoR+tewywvEYYYrE5y05mpumaAzo4Fgn+rTYG+P
wCv8Vg60Krt1xqrJm1Grlzzhxwh9AmcRvERYkmrQMI51Iu6OrPw2q8/ayvoBF0jO
i/vXI0WpWd66MjOzjkZ8KEXyNwhNPZx99zbxK1pcKJUtoDDhVSqdbmA671OzT+eZ
36eu7YXK6bQMoOaLhUlcMSBJpJ+Jv+fHCO/SI+Wz/YgnWdg2Bpvt5A5Gy+7RBX9D
3SBI9KCfeJwB35SSkrVba3rTXDj3EPdlJPOQ1dNxvHolkI1LSRk5aG0NgBx2jaEb
Zbh0rm+puOhh2NKkYbceAWUXsV5I+7Lt40oneZuB5s5TW/lzmBf1wCZ7JkB5BkAQ
Kzrxzr3XsdsTwXB8x/g9MVj3iN+f+Vb5AcXzy+Ov2BP1dEgkkBL7iQI8Zmz7bQWB
MWB0XdSVi6hhjq8eP7UZtERc7JnvGexcXNszAomLh/zKA5/7NoB+V5zobmazUvEm
76lrtQiW+NxtOeL16IpdJ8EZvU6frr/2BbioSyymLPcVGp82dbhO8dCAv5SijU50
kTpwEN8Fl3UzzDhw+uiS/ePBi+ZGkUk/MvaEEiF9AMF9GHJbDj/xrlMLm/ZniPAu
TVbhu+nnHC5vUkmY4NUgVAS9EGuZyvFnpZdc+PYwz7TYL+7EXR1+2Py7PoCFcsiK
zeXr4snhIAuzvyQPF5pq1Yc4gf/nyONqOG0qHE49h8lJh94va8csD57B4rfw3tey
jByh5DXoDpMpn91Zq1KBy2cpi3EHmuosO1psxM/jMVXuv55LlS/5y39y8ec1Kai1
4YGKqwFIPWT0dV/CeYvgXuPwbacyBSsVXoj4m/z9/QRXDGXjfR997C1igmSQ6mF1
hsTX9CuMju//U+L/LfH2HRpRdSa+itSwYO20uJ4PffcZ/6QdjjyofvpCk2s5QtjG
uyLuO1MuOnOSKlFZXFE9isH8uChLbK0UUiEgTHQV2bodGXFdaBgEXVh/zZP41H1W
Ggs0h6zX3AcPqq7N7OrAQupWC5QtFh8ZXVfCAAUB2yUIgnzxu65SEk7Nj8fQD3Hm
N9Nz6UEkLJaQhcvX0AiEz3Vp1XfX9QhQbVdrqx5ZaKb9Uo3EvAKhQwr3pdF1pJ/z
nR7x73GNacM4G4XMZP1SVHdK1/vqeT2cpjFI9WVFPfQ/xZRYQm8nCwFC091z22Kx
XOVzDoQ+JXv4s4dRPKVr3v68JCRd6L9O7aqQNCnL5GPBXoggZcDYlC6HIvLlJkPR
pwSwPaLrvzrCnwuqdHnnZNv/Zq75b+M1HXK+JOsZ27iXSutwZEHxQHvBcWgv/V/b
vzjqXsqQBu5RkTAlRfa0aUDa0fZLXG5EI8INZUm1wFY8qaRAby7+NdsJ7QghFbpn
9u6Av6z7hpQHDFxFW5qTrh9hMUEnUxTqjr+BFt7hwrc7X98pSyd722klUy96WQ+B
qCyCL4Pz9OblkPneNjz4Zko5nnQyhFEZPfuePVv1glb7fsr+5LtFEx4/Q1V7BA9j
P5ijOBuLQXNcTAt04h5X2KGcU7muQsJoY0PH4lCWaVCYUgaFaQvmbH6mg54IxqFQ
x0RXogLdAWkJOcnQ6bCM2djjWbHT5YQ3Vbojym1SO4ng8E8taouMG2n4RZMTfAO+
+vUsfd1C2vt9Udk9VHvxw6cI+9MVlFWdBil5sQP2kfIxOe1MAcgCU0J0aDhh+OBe
2jwpSw8Na+Jl+qSQ/GDQDbs15K+kgRqhS4wQmf2wV1E+DHR8yqi/4MkKefiGqTGU
oViZdlkNE4M6RrWv3IYHTbuzMuioeszWEXqr8oBaP6YG0xvSv9IxDyJMuqa1bobg
IJlDI8zES+V7VxqQHBc9TrPnFi1vks6H2l4XKDu1hHLCcTP9No+OlYTGNKqRSZXL
8kO3uGrWWUc2RCVzx4fudArYWcVIvl/8IYwAmMmtiy53NrwOjwMrmgITr4NXaAH/
LEjtvE1Rx2ln9FmpKlnxOnUpae2gsIixHMc5PB9/GreffyEjD7zpHJRxAzHH2kq3
dvgU5eR2g4NcBzhnim1h69aGWrsZt7Jthm3V+kOcDa5LKQqLQeap1TGo1IEl8JwZ
RmFwzoBCguNaS8/RQE3lW4PK80e6ZELhj/eoiKc9QC7G/E9sxN7DN1cgQ2vB6f+S
cITvfEwZk99ijnCsdWjBmIuxY368TNTJQHKC88Gh628tSt/GcqkqG7Wk13iQJ4nD
2iZ18G79/gPEtsCju5EZ1y40szpDY5HctacdqA00eCGW0Wy8F5y8OLYySd2e1DzF
nxqpBpULS5rENhaFoqlAKA6xyo0AwpAg8hetfiJQUDnJFilGsmmCEGnyIihxmbgs
e/WboXE0RTg73GTiHPI4SZ154ueHk62AvlnZJ7M/h60IbG9QUroaS8HN8Dmpf6Of
Ibt2i04p2HaI5TNSqVmd4NsvPGRhwqoosIUxl34TlwAeXz9egF2K6Xeh9nTnFh4e
uExeJ1fYP+D5jAhEMkb95hROSB+ptbCcVRWQN/IciPDcSrO7vYScKw8cGUFRCSz5
FIaom1BdtqyCx0X4hVXt68IQ8OCSxm4+BRYvMaz2zgy/21wF4+9yX18detQY3vtC
ayo3KM7boI42LLpCr82g6CVtH2uz1m8oqp7vtywjDP2P0GFiqwuVCCQ8mQUJHEM9
mEB1sERS5OW0Bz4s9JE2buerXQxUTOg5Ep7OGGOdN0oWGugAEIb61ACWEa2KBK6K
m0jQcf9ogivbvR35MNTMHtXe05Ct+0eA8nGvGjXKE/oDSeJGjYsqsOW2gdiLtmMO
tRpS+Osk0x+DwBQ/XUZT3PE4viTu2Y80clWDzgguC6QPFWaS8JjqwiqasZq9XmvX
AZZaukQi/3lJBklPYgfDfdwUjMn1gZlLJsZch1HoL0ydKHZYeYdHWa8HctFt3Y19
WYnZo8b0GVDR0Eo/YACimw1881S2ETP1TiRBJ/GChyo+UVoS0C836P/oK8eHFwi/
0en+jsJ5oL4FO2Q3ofsfcstJlHGGnEeOGpk43sGdqHr0kKLjt2FJNcAZ7NuEX852
G9Q2W4Vdx1Hh7k7pjgnRAiMjBCDC31c5pRGJpqsZV3eUuyVEbgsVyZCZ2gmEWF2J
BAiJ/vMt9g/CuNIgvIMBJZYPr49CwZW1VAazlhW91T1RMvdhRAgv8H/bnC5RT3+7
p6M104D3wKFklZB9ecuHU51Ou5vqMD1hMBnlH6517zwFZrc7qXZEZ1QoG5UhdJPh
mzQXq1oSs2FbA0pxd0noYYlWYcq9Shg3BFZf29pDkk/MD26rmlDpH8oFHOegZAvm
n5stp9Cy5FozgtLIrw4kauUfGVet16pmZymclG/HddaT0eUuRclIeaAE2+NRjv4R
/UlOZ58fmU+Y4R+XlOgSGACyweqPoAE4mcNeUQVVPYhykOtwYpuxZEFp9cQaJc7D
757/1t3OrrKWa/ntfd7ZIWU0kxF2+ZudbsSK9BjnvXHAHztRtS0akzvswB3v+64C
7fPMG1gy0u4ZcP0dw04YUjkvw/ilmT+ow4yrZnfMXRIbO/LneJZzwcJ3nJf1kctN
b8jup11Ai1VI5HARMvMhlSRurGJ9j0aBuOK9MOkHRmArR+N0d0doVW4JN1ia1YI+
ssN1SG4V82SsOLXykpYsOKqgxCLPqVpNwbGNX+gIJ90lY+mge4ifLiSxJ2/PNSzq
+RTrC1QHJ4LVhSEVdZdilbixc+ziNwYas24XdlKNDhpFLV5+YWMl3UvT0DIkaPPS
fMRXv+qd0kais/2h3v8bPIl4GnAaUWYAbXRXso2L/idQ7JDAFlbxNNUUf62hXDZA
JoUwRuQKW7kI+dOSYZ+6f1Cqyefh3fy8/6qSjz/mc5d00/W4QvMvM655stOQC7zh
ZotkSvdyWlnmMqM7F7hzE/jQkshCj175RE76Og4OHtHXyuntV3XHS9OovMn17Xi4
bYBubMuI4iV097M8X2r2vDAn/yqnvuvOMO5EiT+awEIoo6H09WdZTTKWXQI10465
FNloY+vq8BrNzEjpL+Sd8Hm4iEcKV/EV6gTPD5V5VFD47r35wjsmr+SCFhzU2Bjw
S15s6lY8zWRFoFf9EnbPay6gE7Xu1ltzIz0KuAI29qWi8WDtPNckOS/EEJBOgpld
S96bNeqYIxRMOsBqYEmL5ChLX2+3J4yvqapxUgc41P1dBL3BcuJncQlhQYj+l+gB
81owLWeYrxjwgJDvEXQOkEqUbyIAtwVJj4e4seFeJmGEVOiOSoZjSvhVvDp4tcLi
LkwBa23uHp8E+nkG1JL617XNqRHVz1ubUBo4Q0ZR/j8v5zPfhBLGjh5bI1TjQ9/j
Kkh0T7D85AifmZb8FybwwxCrcCVypj2DzidiVIyQwIsIw3yiUADwudkc2Wf0TQg1
qtk802OjDaeGok7FN0nsOckL00AF5dcJlrpKw0vuoIsSAIerI5FaID+IUldZAnAK
8pL92syDIew02jXOnS7ueJcyR5L0OjH/f2nc3Fn+aNK8/fQJ3Nvi6OJ7IFWtDVSw
QVThCwX4g3NgWblsF/aCgwJq3AzXO6OZXGYbZkFb5uZRVd03MOzTFqr+nvxLdGcd
BDsCs7YnViATDbXZcXyGQcLjlByfdjV4iTcEtl2ViGXsQabfuYJp93KozmH+8k8r
d2HLmm3Fknm+ZFeRyEiWx6wIaHJ/2MEr08j+EVJ/Tp1OfWPDE1nRGw5w2jbBqbw8
v+9Xk5NUqHfdu6LGsWfXdvnHbBEM541Jlu+mvXE7Au+G0AxmgwbQNJ2BUTXF3jDX
82HpPKzNhUNiVVrUOM1a8UZLvLmt/R3Vn/TKBIcPPx/cGksY2TJUVUVxGW/t0f6d
PoN6QHyQvXD42WIHeNFOIHjsHAs9E42BK560Hkpz06OMgH0+SflArQ9gYxllRSbf
BY50Kgg8NNxNswomaWkU8zvuC/dXa//zAaJo+VL6WwuiitADYW89kpA2kvjX4KEJ
csId3UZke+Ml/s6UX4Djen86q4NofYTe4MqmDO3pgbDPc6Xz8mvQ4+Ms9drP6LBn
eFOUr2uY0p9XmjBrZbc3LAWU+TU3rVSqGVkGVk4QHXi9qPBZ6s0PFMR9VG3pMyOM
KgdiaVBrQyNEGke/qB1xZCgjXc9dq3xIfNLtjWxwlgakyklpUOTL/PveIW/NJB+u
POyDpfPnq3xa88LPTbDQtA2GffEyrEfbht/ooEU//doDScjVCd7ZuaiEcVu0CqYm
iXfgRmgUVzYuwjnzGv9gIBlpRfVZIbhrcJBLqf9FQz3FKl3a1Q0+gOdYLdDFvl6p
3n4TMT7QfQ4uSeV2hFmlKw4M5yB4/uAfYRvyeUOLaTI5j8q3AD3qFTOHxz7euGPw
CPV9R8WBr6PUZOQNuF1zKySNsq531CAXS20wmVYOn9/3VRrv3gb8IDlZ0QVOTnqH
c/oukYEw87N5YQwm48xhgQj4PbCAb08gPHrypShprHF4Juih4BNaIffHUg3GSJYH
+x5GweriXdC+E3WMzFrjMLxxZR+3Ui9Vh/Z32QuNxM/6XgmfQlnwBIcmvtC9Watm
92ZuKV/Lq5xSYG744pDP54WrB7O/9Hq9gJypqf6sUva0YsXXg5WXJuBdCNFT0ezy
jHxh7gn6Bj/hMANnM2MboFpPy0CW66d7Bz9UCJwoZeP8ljZB9qtbFs+4FeXKISu3
zCjyFEtNg7lDHB6BRfa1X64QkXBWrGJF2VRAM6DiaNZXj42S0gxEVUYzBmOUzKDB
wbygyi6v1SB3xGfuXim7vDBr6TctKw8GDjjH/LBeTThHY1mk0vhecqiLVBOoIalz
LM7MXi2K+gUqbh+7zuO1dAU/6t8jC+8lWyXdl8dMfibpU98nFDoFgwnDA1QW7MuZ
V8L4b3cRNO7wXrzPjIM6BVU/992YOIlc6+pHjDCH0NcUj3oHqFg6C63NfOBn6bvv
PBPceqHBF4zz4VdqNxDEmxOFkLA698rattxhDHRC7IyWBlcPQkwpI8kLQVhg8O9m
QS7C4Sh3x+kLNUw2p4ytc5qfCENYvrkxvqlKkI1ox5Huu0j0yabBVZ3VK0z+FJSr
nik5PcG2cS/nC4T3ZEJAGjEYWXIFOIFL7xXAC7asopkJXrSZARaWyqnePzq/O9o0
w5qlGFuninlq9AJOVIewhVWMsBVvY+00meo9xAZwXj+vuerzNAFgcUUnQy/ZDhdr
+B6/YDTlQQ/5Bj5rViNkkyFlwTOZzjQHAPeBvMuaLaTXPPtHAoI2KVd7GU4loanr
IpHB5Ah3DcZIOwsNGseg/8h1WWtM0EN45zJb/OfRW78DoSbHj0728jOYHxsu5EbG
quuX8GpgT7U9xH5b6I22QafwhvzDFWFVuzpq6hh2gvTVIbOHtIk5EMmmT6vIrlZ1
DEgUSDmSMV7RbX/vsjs9KY7cq7KMELeZzA8gzxHwRDkOt+nMJfQQYG1uo+neB1x7
RCtPdtFupOTDZYgw60+laE3S1bczVyhiTq9mKWqd92QfSQLT3nionlISRQqSj/FP
k4+zbVHLBv2ziWIsXtpFlw03kzmlGQa6DJOEZB2HV4wPD7+guGeLM8Icq4N53H8+
BoyNa8ETOZ7LcT3vzzFhhyxAGfECLu5/yWt+8AxnwsPG9Gm0BB+Hl3I0lmY4JEoF
qBq3zV/jM/1qm5hI8rbzPw4nMn/meJB/99oyoXFhoyVDv3u9dkpOLxamXlX0efrh
DNYWcowxj4fIdt+rD3l5j4BAwJAasG79mdcFV2wT7NMJGbdfc9cHWAH+YJuOoN1s
zr7sVBEl+RCJjn3HkgfstJlhnJr1bw0efGfBHd/7MnaunTKqHRLaTmmu84KxH6dl
nEMkaT9m47mn26fsR2fqOzEO9Bkn4Cb8qUZJ9ZvaDqDgEyzKnb4gpd8Nf+PY0G5e
CrXeiRenZyek8anKS2LgwxRmaPPNtJnAKB8KNLll0/uk9sJIa127phGoUwMTUwMx
R4GuhFZZd//cl+mgXKq6AfVWe1StNjAlbYNuPrd5ZfsbOmROir43bUXpbTpQKxEZ
JzHnUsKq7npQrRkxQuALEXSI6XA1iOPigBiOUPxZhYNuk4jSgqkas9UIaxfQ2NEo
JEEBoWzrvgLiONlsTJ5Xx0ViS3yVQpvRhZr3aGmgo16hRBAuI30ZTLu0jcRx0pW/
vHlmyyj6BYu4oW07hqQm7avPxYxjcrieySY8yxM90y/lVTH9eEW14yLv7VPi5FoP
WvanhYJ8VFUkDyy87EzOWTEr73Rh4RgW+uqyTk+KYrj5lLgA2T+doGIGgMWzr0Tg
Wr7PSqj2PEjSeEZePIqKUrLEF6+RdnKp3K+axzqPMU9RBbtfY4e1DO3mRGIwIydv
SUFLT+oN/iq+YaRPC5anGPAhj/Beqxg2q21Q/w7dY/A6SW8hZSc4BIMWjnWabxCw
CD5uihbCncxYlZWVW51HdULX4qKkJqcwiN5Lw6pw9KeNZTGw+jI4wb4mPQX1V8wM
HLKoTrV7KqbK69b1zTQIiJ0JyyJ0D8Mss+kyYAapFfMSgBP/4gKlZvw+QsVqeJ4J
EKK84nUu/Xpq06LMkL9DXUwWL1inNzO+JDyVu0/gkOHq9xSM7aj5oWbv0zBcObHw
VBe5nrxjNmNC9QaW5F94HGPkRFuHRnYnst9CyEqz+jwacYtM5b0DJBnudNrObsNj
NShOZKAOyLF3x47xXCfQdUNgwPXyYQuIsdWDmp8jzVOzDeflBn4PbR5O0f+slJvJ
vSfXV5bs8SCiqKEeHGtfff4rivUEnUftkmxZQP5jkWaQBFERb1cBFAEqRtbLkpGE
96xfevRFIjIHJAWZwhZD0FfIVGnQrTgS8qdg2lSSs0H/ckOFPTKJh5zj3+SvAIDe
m+FR2z1IZEE04sbL9OV+gjP7qvl0ap7kZFCoaMLAgv42rF+ZH22pIjSW7hFIbcPV
JSnPSGZzDO80UZ3Z/MzMvSEkNFlXVVDfqh7SRbtWH3aq2b3BxSdw1b0/hrpSAtlB
xNzIWXIZM/6VqHcuZyuRGDb8jwnuTYCz8DLF99E1S97Tiv9OXBN1xaGL5RsLplgm
RLdwoBQ5L9pGQH4iL/JhKW3tejcACo0qXDZxD5jMRplqLHKQSphtfudBbVQ1Vn9B
WZ77IPW1gla2re1X0XfTTNWWBII+v//KB3n0rbT8mi3TCJY+c1kW1dPVHCQwey0u
XmooIhzYYacpKnRcYtr0YLAVyRIoamgSwz9bDosuJw232OvlLwzvMIKXs3OVYE4a
r/qQEhSfiGsHVZILl2lxe98uM3iauVYlavtFxN9UKepptxF+gLYxUgiZel4A2HZc
m/4zr5rWXDnO+pCukFQdRWjDpNWoedDs8BkL90sdCYY+hYgbf8UBJaiQJa+2vDD5
SQEYAZKh1FSbtWWLAOLs2H21jcQhyz6kj1KQralAXIWTlwYFLyBVzw3Y4oHaPWHN
tmHl9pnHCBiVNDEnbXUaMQpIbBI6/ynVcYZ0Ad0hOE5HQuL3jRr59P2Gnn0PyeTX
BimIi6i8vmk+D6lLKE3pefyP9qElDrimgMlsIg9Fc1ctOSXtGZ+/8LjLo8Sc55dY
pYm699xegMB4FG/OFQw3ospzbLSXTPUuQG6TeL1J1DR92Rp6L6c5N1P13MTwOO2K
OZXHi9k8lYK6CdoG+MAQhhvGP3imqjWqVRyJVSPXzmA=
`protect end_protected