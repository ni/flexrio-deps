`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 38064 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhKhfkQ1RWny5iJ5zpOL+J6n22O/UCwa3pitUyyRK2+2O
+nk3oq7qNLyVXq5jOjGxRMFyhObnOO0yxDYfjVnz87mQica17ynm/Eo8Vzxkya4P
pm5lIyt+yveaFj645+qHCjXi8KQggXJySK/qOT5+FVm6MLMA6jGyi3dHhs9857cb
8BilGYT6pWZFohWPutpbhJfFBg6xuDiA0pDGrMtcugOj4y+5zAA51o1jpGhYnk3E
U1GJqqL4d2HZWc4yVmvFEC4ve2HFyqAczqzXM4xCp4v6b/As1cl51kjJDpZiFY0I
OTnJL4MjcDW43OzkLImSV7m0hLOka1gufI3O1ZIVlX9EyE/yZWiR2SFgHVIFohfQ
nBxFrkA+crRsg92A7UXFuxb7EAJqD+OIZ0RZZ5gpAC8gMXakn3NoO93gs2rVqLxY
hg3Fnd8NxHEVtRS2IuQqGMPzztuGuuqrVKkV1sC1LKk+UlmPzoI43TIY+jxMTJAw
uSiKn9Qmxq2MokGsR6J+J5ve3LoNlfSlLg9Kvpu2JpxHFALBkHWbyWjIWsN7JwNJ
bc39zdYHpEqfgZtCvQcL5jKHPlZVTvirXA/wZEx7Y7w05zkqsN1ZG7wbPDZqzGxc
zf8IRct88ShLEvYGtPX9EV0XGF0T3Ei5I6gVV7JM4H6dZcFfF76hrSognYXSzhTf
QPWN1nROcR/+Z684MNtPkSySWfymlXrZAoCG7UIgfv5XenmztGgYfnj5VZ4tTqNF
FppDWuqZMWdtCNNUFXK1nU6ZpywGdS//5QYL0gLUiInvI9kNquZIyq8Xw34r4VEx
6U2Ck0ev5Vj4J2zopwQ0fGhRON5pH/B48qWXO+tmLVHIQ9pwQSmqN0JKi8NDyr01
GpVNe0jnLAhQ80dAE6PDj/1irKedn1PmZc5Xw2v6c9aNysV+WqXLDYKAF9V8Bq4N
csOip6Dz8UzNTO2shqvB0mz/6RGnr/ETM1xsW7eZ7Q81a/gvVpAeEE6s4NWY3nA8
OlCiMYs8gl088Su1WUrKnGXdDAZ7SRxpOKw4vkjxJvjfWaj5cTHqj+pBDUb7MrLK
HuvRz6Rtby66I7S+bn5UZEiMEbSC3eEcBFlzjQBIjkCaIT3Pa1Xpjy3juncv5oz+
Y2EHNrjgb3ikOzG0on1XrJ+9nOW24XDi8ar4wTIWRiouhUK+rX8pier/BeGJvKxL
yl5pa2s6KDywZ3pL5MCfzPirCShin+YC/T69qkWuXRjnhWhUsWc/cw7okgSsivaZ
yPD1MCjEBDUIO21U8nI2YIcZryndBQgXQKBZOMLdeVUzxi0BU+cO/cqMtA/NC0N9
vUn47OJ1fAoDpplxSUuhrzw2gfcGGBqRNim/IV3GbcOIFPnBUSK4MUJyXzyVZmfx
ZmGfz35ALbeAE20ZtbAI9o+yQ8r/2ZHjE4oEBtWBKs4B1nwpGyAlMvB9DY766r2s
+REJlfFVBGCbI0Q7GQpzFIRrOVBQv/EDkgy2NKQRwPQCYwWOfq2lOwg4xEvbyZ3m
t598ReNYO6yKgwNrccc7qhuB/vJ6Aw2TekWI24JF/339RloRwX+EioFm+bz7TBt6
LYcgVqfkvbYE3M3KDSq/zddABIUVdHMFpBoOo4qDWiNG+cu5F3vVclke+B+MTXhv
LhUFUTXabSGp61EC8RjSDeivRNEfAiVF9InYVzZAKrFtZ7w+kRrpEIDI27aMOt4O
yYeNYMFABMSv3iKtWjJmAyp9eMOqBVtVd7Zc78Iyb5aCqe/XuzpkBEcJJM7xYsJV
J7d51LpTeqguhkEzlPQHrDAi6mToJgoGpTiUNWPPTIO1/jMr6oV7ox/Y0MkH6Cjv
9x7NTaG4zpNvkdlhuL0p/UVsPgdiXm9YPJ2ha2i5dyYbM6eJ/hL9xayWac12GRoN
oW6+Kpw1aUFWccjmpGYzRqhiUT5vN4ypqWCiRfEFnYZqMXUhTP2qbhHIeWB6RIZ4
h/sSSKDM9ozicRjRN3++2NDb97GiZVqpxZOOtDO66Vr98p1oKGtrAimKkwvvtuLo
fObe9zwDF7xe+91aGV6lIfenqjxMbXwLA+B1JyEc5cN75NiHDcnCA+BUX1CGwwNQ
staPP9Rg3T8LmVChq9hCp4qvTOFPzENPTjp4cATnC2SeKUkYdnzI/TOicPxiNCdD
cMWl0ncGrOpIvb1PFNEpn0qujidyFBwLWYIfpD3kk5ddi4Ty4/sRKMoiEjTvAD0e
ay4GMtaP2h8GVhzmAky7gqPxQ6tyGWWpFPIj3sIlKxU1nxyfcrSr7StVgCpesuw1
GKrWasljcivRgvR0ivJNy+UE3SV8R7Afc90aN90TYkNH0jZjV38w0wXekJexjnPf
UYgHntFQxef4QXqzzjFAP/5ZlI1s2E8Fj7RacFzVJaYBR6FoYzMJ/qF0zZp1Non2
gnVZkP+/F9sI+h/yI0bo0tROsvePhzpBkwCA4VbcR3rfCYIKeVgv8ne9SDwqIwO/
EJsTBIuX+r4kQ30MslhZ4E0kb4DGRG+ugFBDe71aTZYWESWkCQnWfomhx1Msod0V
Ik18H58iWQv/8vw7StlwL+TaNds5OW5LES3lS7PehEKbV8xE6gCV+V3i+Fc8oWuE
x9nwqyOcbvBvtWURIpJv2e5tHyxUjJYI6HDdZEHq60oBSiIgg9z4WsA4IPnpwkfz
5LdsOgKambmHtqAy7YVe89L5ewtEc9epZMdu//iusjYSor2tpHwxZ6miLBxNEby0
X6xsnP9733A7C61qjyvi0vmYQF+bJJpM2SAY61RzcKLjtU6wjhH/crAUaNmFszZg
d74D8gi4/HPXiGZM/AM6/e6GZO9cSyAQAUv4rGtdii77iB5k6uX3WWcYemPE1/Po
hcUAzaNPV7godZus6cqcehAlouSBa6+0UrcxVmay9sVn7ASW1bvWeA6z6ovdV8tn
Tp8GaMT3uZvv9SZ19sXtzNebzLX19wXxc7Tvon7cbWLRKHECKJtfkdqeVBlZs0IA
lKmFbY3CYccSM3/E2gHJtyohDoJcBwyZx+f2T7uDUszg7vrYDBqPj6qLikdyn5I2
vNU/Q7/dygQbdBptxqmy89R8mCBiomXsBiBJoUOi1E4mlNrFDjzeb+vcYSwYkkEB
EAxYP7B1tFYXLw5IzzekLBONPfV62ha7JpgEsaZ6BIuWJ1PVEBYegETIdT5FqC4V
CytPkpbZnovE1qnlN6t9cXrh4XgQR5LWxDM5uMMvxVb0QwyX7IRq5mcL6RuM9Trb
qGTSHL/AF6bvWlt5kvsiXQUdWlqw++Axpa6K7zFrqPlajmc3U3isuQ8G86+AbaUW
lFBp8WBdxcnpFUp6njxssZfByDfdEirxXobZBDjEBjpKfqmkWt4YWKFsMYAP6qID
i/IvalqDg5WVxWUIKGx4A2wOiXqXb1QgPYcam+bTtwdDrPPd8oM7YiRsjj5D40Ro
Hv20SfKLNixXolv9PI4yR7euWiTaAOpQgj8RvJqiKXwWamwhKfAPfzJENLYXkzFf
F9X/9VozjuRP3cojryWS3Gi7znXgf5IVzDjuR4IKpVVIljhIWi1msV1tj9DgCX1a
AjuMe5RyAKQ0phK8Y9eH5Wf+bxicSUrZQtgpQk/vvEFIpiNK2nWLAAAmEX1Bxaf/
hvwWh5bCdcovHHzpE/zoqqxnM/gnHs93UC3ssrEqgW14x3czi6J3lYdknAMUuCRZ
Q1xUty9OG5GYQ3KnPnU37Jo7GcnYlzctwbVXiehhJ907mFnwImAMcAM3n9l7zDf5
PSdM6w0z4M4FsxOSuIJrbv5G5YwLIjEXy9f+7Rn+xT/omdu2TgUja4MQC0xxTmBs
X2maS7HPhA9LZp7hsehbFvLnDTclHqzJOynbIwK+qswpKQX+O2iQtvb2Ok17OCS9
dorhyeKP4pgG6n8I3QR49SNSTAMUSYpa8Qae+DdxAJH6NX9MX8D9Kr0yjrxf4P+s
3fp0XzGuXdtzYQ4bpP26Ve10y0ih7wDDrx2ExKV732/VMQ45L7y9eCMLg+ch5vpe
Cskv7OF+R/+NRZCzQyYcw8Pi7gVdDXJOEwCoQ3JfpDHLXgmw5VXqlZ1XWQGffwh7
H8g9y0XKEDQJHIDO0uq0+qdb7YuHmLD4FPV768Y0fNNKA2uQG6TbBM2XDi3ShrNz
iDTdyFGHQWMNcm4k/6QwNUGbWv6i7Qp5lcecP7L36VRY/0rK2fB30YdyXWFfPCVn
qBCBVT00dYeHtfHXgQXRotRGzQCd536WfZ2+6SmfGA/IiEW1XThOg+ZT7DFZLWZu
dCcdEU6VrAX49Y78xAx71neO1AGBmIustuRZSVSUnD8voeNPKHEFxPYERpumleou
mNslwzeTwVyq3Jlz4eWPyUU0Ajw3GsGpUQsAWaW+6rqrYkhVcfZYPiwMaGxzHLsC
J39tpOGWYzfCIaNZyrmrIDhUrhuYbTzwVuVLctf9R6jRQwrjV+i+InwkBm0Nh0K1
PbzG5vt+y1T8PqaScLanqAW5nq5HQvR9v2vzyFVEMXU5Mmg0H0xDcSBklkODwhm/
SE11XUvltH+lHK3La3iYBrnaEnZKua9EVGVc4NnKpuw2ao87pq+TTLDumzNm6L9/
CpZb3Z+7O3HC/r6+im6dpz6ZgwAjdHq61M3d10VHDw+VcdLDyzbRDlJ/c7vg0196
LXBcYK1TYd1QBaqioUT+LQnZ1bou3akc5SwGAKrHGuA1DcQTBf1e1ILq2nOGPs9T
k49U8EYuZn4SZiAWG4drK54Py8q/nFV6nRj5BdyN81kSu9zSnAUC8eB2Ku514GFe
mAdJmCgiSqBrcIW3Fwj0BFqwXwgepnVH26Yy20qBEHXMF/tcBiA0AmJ2x2RO9r7C
NurfaSJajBAWweDkWnLby7hnwZNg84y0VowELgUdYF2JrRtWeLgjuKYhD/3RYVyK
zm0Emc+0AO2yZeWRE6AM4BVpflZiU0jaY4Zg5mbA6rerZxfnWlHMdUb0xfQipSCu
IsoR84iF5u/4GwB/g8qjTAcbxmdlDNIyUuQZ3+NUUfEqqwI+AbyqlRp7QU9bSBqx
dfp28p3dgvJDfy65DXLG22V535k0PKayhftlm8A3GCNs8ekGRfDR8TuqFKptk2Qt
0cdyKRr7xCIJ2l3v9oLvLbudYkYbp6HH47ZcGIlaEtjIuhueZ9dSq5+11rVtyaaf
I4dBI4idAUpBjMk0L4pFQKFedRRuqwcO+JDFUnZGxSSQsMR+oi6DUHFOI55TuJ36
l6bDZ+xWQHMmMe4TwbbjJ8RYUERjtCXmtJgIol16yFoXdQvTDGxChhS9j0OHZnP8
RIn+RJDQQ4fw2AtwWIG73WkBR7uqi+Pu37h4U/Q2nmpvh9/rlzJ2ujb+aVZ0IFFc
DJBfkU8joR4/IMyt6YWRHQXHAGFNxR6MFL/2WyYxq51uDe15zQ8fanQl6+UJyi34
TmQ60quM3fi1Uq44LN8hDMsnx68w+nN1ArbGSujzQCLpRjGwuEwpJyblQcIKtRfo
pzt/v4BhlGK6FQaqS13kprdg9idhfntodetM/AWHSb0tnDjWT3+7thR3Cg0N6JRU
ztdMPYDw73br578J98XtCqlSH+mdhVe8sUkNS5uhtKeAjQzNhARTFQEwIdAi+Npb
VXEtEff84Qgtl7o61azmdHkxZM9pZno2vROnGVRLrhysz7qIs3BFaNuAn73CdCrq
2iGFSkXciCwHelLm8vGCX7f96jDyfjZpThDKMJNe477ZYMKql8l3ycyjkk/OD5AS
1mAVtF/r2zKXEMW+AyPnvSYjEVdnS0M0WtK2nzWJtmI/cMEzlJcbdLzITFvasjVR
9FqyRHARww/J+PUSRrOJJK5RcqQmVoG2JleOVFZLVuqVI+LC2SD1gaHj6y2uUovV
ydJctZiwmjjjGoFqcPLvbbODja8Gf/U2eb9E5ufpk+sl9HCjExXiJxkT1Uf3HQrT
h6Mbr53KwHo5JzAEY/TSZJy7Piht1stj2ow6OlyNBVNrLOjhMfbz23pvEIADC3Iq
+XqPF1x4oTxv3JBimSAjYA/vCipuudseIzNh/M7OWZGS+OqRI79P5FPnA8tILvQw
l0DrzpmGsZpmqY3Uoky3JEayEJt18BC4J7hE8ftIcpiXMWXanqreSDSWDZjki3x4
n14WTQ3GNO3QneoKwrTjXpDFYuYVQ0TxCFHNkuxZbIaFTRIDy3TCjgTOzyKDuSJR
F+M9LY66ao4fvnLAZiM772qQhcDnk/Bq8Rsr2aoTfrqnkH68mJs+fOFq4CwvF5ll
DnviupkBcYTWnAMfbnqWov5EmGSKvd7671z4y/XxR5b53+K6Xm8qYRhjhM27B3JT
LlwsUtLfErLf4KQExFd4+Z7xtA1tPaz2NH5XEoHk3kJBZU49nLjrNrX4luAl9nTS
v70yzFz6WQ7l0QPREYQMR9es37REBle7uMlWrfOv7DnvygX0aHDLmnYsboNww03u
0ebj3oCtbLcGsthjWdWgrNFbB0xlBsNLSXLh+kfJsz2E7zPu+yRl8sYN/dUqNEAb
2rPRomF6lv/+CVfSlqgDI+Gdxb7TuAJ0cmtgD3qB4rJTKcy2PP42YtrAY6Ti1pzz
JE7SWJS8Njer64sUyJVkX0j2dU94p+gJsF1T9DA9x8vukJASqPlbrQxJwDoJsYk+
qaUwxHvPYNx2kheVtAXVOTEyU3dN9bIkwW/MOCDG6e11zQhVNDf9o0aMF+fYgPS1
atEQI+rdQDrYYq3U3rzufbtfsm4owuLAlj3uERVhNxvmgjYCrj0595525tlkIMZG
nnyvoP3AWmWDylQikZkxFYYMNaLMWoAFmu7lQwySu9jjzlKMrWOvlA4oEbLPcZbS
6FcRiU2N/6V9JblZ2JUHXPn+zQ84rT3hqZUAi+tZ8Xts83ldpDffjr0MRCZ9hVPd
hdGImBjxztlDItIQo9k5n2GO5oTq0vQS8tNyqfp1LnBX42Pf6rmh/Sg8PHNYFsrX
R4MgtrbN81Bz4EaeMN9PIuAxFyIN3rls1X42jiKWi+VGh9LBvHWOOCkU3Oaj+MEu
IpCg1Wb/r3ELX+b4VDtEsPOxj1Em14tHX128mW8Lvvh2qiBha/XT64fDuRNqeVch
1PsRJzpgmIpsNG3uAm9J+pQNdgQWqPnzRvWROaPczkcjLF1/XaqlkVwWYuZLAUrR
gdn0ZLChINuxkCVC4ILg3dPirgvXhiN3S2GkNT1X/tHnPyaMrfbec7jAvsPTUzGx
12HH8Th/X1WV5yAwXFVO15r00oGA0i9OFqP0eIm5gY65DIhbVdyCsgCy8qZzJjD2
npvBBVPsNye64MuOGu1KPpdFG5g9pTtIlMF1e+qZLsm5zUHE1sNEM2PQLG+nQ9Pm
T5ULirz68C3Kp5bHSqgCG84f5OJtmUVsmAYvu4sB4/eWmtUuySDvrH7qLiC6281V
QEOcR1isDeQmYDh10gwFi46PREKVuXtAoEUGtw/1wKxYEl6iVqKs3AgsNDpwHpAc
9ioWLfZirs8em1qXaXsG/yW0tve0G9j4Ib039tvCca39bGX8XhgEkqsZiYTHL1x4
I+NKMThKjrVb5OqYcZ93Yg7qJdmkwYGo+Cty6k6Znh9FePc6p5MmSgiQPN4YY7Ak
GWLqLZSBQci+fhldWPtnY+bvxTKhrkXNK5e05j4hPciHYxIjpuQR739yu08Wmot2
yZkZxQgp8HmgRYq+bcUwRxewUFP9IYSYC2NDt021T9TKUcfIRTswh6uQoEcrvnc2
unsL4LTgw7vKnrIx28MRq8iV6eVV+okG1BIyyQYZTYISUZ4/VGGVwZjXo929IML0
35sriq0wglyop405ktKtnq3aCXvanqTngfSRXAV92kweIk79RlKAJ3zlEJUEcfnI
mLGlrZuJ8iKvjbzycyh7rk7pa6hVpOBdTgYGgsxBmZtfPd06xQdrzZQoYtIFnycn
KSzM8ikm5r4AlvK1O/Gvd2EmIgP9/uiwxeA/hDmdlr0pdMHz6Dij8Ps9kVEvQiKt
Kj28/pO760MsUOWwJ1urL9J7Jj9cJCGw60TuJRMlv26NOUAVKGBLSOVSNkoNWutY
nukTbt6YDbhmQ0tIr97J0EWxiosMdw/R90G6VfOsEr1tSmNtr3dlkIzWjkbm+OJA
oISvcx9OxBvl/xc5gndJ1xgRccJYuF0Mo9D3GfA+qysyCfbPWF/P7WbmU3LV7vHi
8YJU93CwwdIGpjIZBlTSZDUB3eqfy7xnOE2uULGJvy7Ra9ScVS++FkqnmkZQvdtX
/8u+ffycZIfj3LPEViC9vAfz+nGBPtspwKC2P4/LDycTDdLByGX+dIh/GvYLIuLG
epb1ujqJfL/pcY+BHetUhv4vYKQuGABavMWnoVnuB7345Vhzgc5QTO3/OTH9W9+R
gsdJeVjNfzzTg4Y+IvRzQpR421KTStgQdML3BDYwgMz7+Ce7lx6aD7NAjD4R7X/A
DGzEWfeoKbosQP+OZ7TFtoF8ubSuzTtp60dx5pnFxWuAM8L7Bj+6Hw+WsMjLgBh3
i1uAXh0DjW+tq9uZCcR+qwcL9U0eBFsV43MNLwxVa/HHicNZEXCMKeNHLLy//iO3
fjL+nxZWKLXYYxAf7MLVpyjuGh5ck3tqTm3Lm5h4xqHLov5K8TbF76TrFq7rO6oS
5LILOcObwaOQi646Anouq03OmLqpdxdPH81wRqIlYEjdBc9ku+q4qlZVszsBoe8Z
Eit5b6UC0Zq68H0kPczHuTfU1F9V0sbvBppPlMuhVqZksktYbtCIceD4SkbjXF2K
iaY+JWjHw7lJ25havN5cW+RCUnjslSAZublRHX+04JW3Nj5Z/uORzo7NK/3T46YU
NEt/XQ+ldbeJrgH5mJotaRcsFgdAt4PmaF0WIfXKI9p6OKWyVX8g4deKNDBvXzaL
4NeooJnx3il+BfT3us6MC/QjlYrsJLXi4c1Qr9zj7zbObkgSAiQbtTvIzevwIXPF
SQWfL353mQEDUPDVRdSEJg7kQHu+N92zyy+SWm5ntdoffEpQD6eiV+BD7C/4Cboo
RGgqBP7v5WokNKDLEz9ZF4ZkG2d7j8DUKJMrHcJcpn75ahTKeev+SNMQTi+1lwL4
HoOP2YEe+Y3Y2OyIeMKfQ4Ixos16zKSoRYCVM1x31Kk9XAazBXkQ+vHi32WcS1Oy
XdWtcpVTLVwXQo0BcH/dBio6UDsPnCjrwyGMSw0YHfwR/gzW67K4qShm2KkXxnB4
58M235eTvNnd/ikepYoAFFP0mu+hCHI0BBnwoSIMRvVrkdojJTB+aJQ9FTTLvUBh
j5AQ+4osXQbsQNSxSQIUHeFgoBjI83xeEQvBRu7XPL/qJCVYBnne7KT4CNeKjZ1F
txEWkK4zlvSiazDNYYZcsi8rHY4RQo7nZ22v1Uo0Q+Y8PbdU+kFHE9l5lEx0VgUW
PpfC9kjt0BcPC4Vo+hH8xiq/eQz9EP0FBJDcu57x998keUE9qqpTd78dOarEtlTV
SLnKxC7CpiQMs5joEiRZZDRc6mHRRayDuXUp9JriB3BhU4U3CTAJgoFOP0vNziuS
agQx6a9Z+TJMgdScIxOZpUeBwg7HIiEuGBVGwLe2X+QSkYSfiYUFCXhJWBHZZRph
MJFAI3Z9RoonQYLQVap308Sz+wOld+1iZNgD8GD5+wYO+dOhOeKruQQzR8OFYOu6
rsejmVElzTZjKsItBzgEdzWXM4ILeekWjPyi0uUJ3JaPRsIq7pYkxZ2gYsXDhMLp
SCTO5GPUiy+VfVaOLWJ0p3zU1HVFf0ZvBlaKTAI83AaVw5t6SgKit15AebtHaSK2
9ZTjV5+IEWbfb4x8kSA630XPbOQkJcpbdsdpz4Q+pjT+uY/6MctbpMTqhmGiS7Uu
KFpSkSWpgwTkP0UbGyPZVZRVfOK6pbj+MXFMny1nn3mDSElqyW3/y7ZDxey0dg3+
kd/QBcQjp5WCCHGQ2K2Y1s7yXyDAlQdneMOwKDP78pQAkszGraK0/CuPG0rhcP+N
FVmWtX5ctxQIEVlNv2m0oIsc9wxJLqylria1qnG21WOlweq9P7BM0z1bNDMTMhnJ
qYeVNQxyl88sn+NkIeCCJd0ZhZQ50e8DSkz9W5LMf6pDziPAVHPjdXZYVEiquTlC
+/DSKszC66sZN2wWGFowc/jqG11xRp39fnK516PhRog1Z3M/XRo+U39fxIZMp4+S
vWAWTVLy4rDGqPXGJpoKjRMzI1uOEzmWef7XCH8Xry19BMulY7xTSp7sY8tJM5lz
X2XarWgS2b13+KOxTM7fRHgchLanHBpTil3R0kOkC6Wadq0rLySXXzNw3E3F8zPS
7cPKlw2XMhT/Ak8Q+Ys5uofFz5A2D4xhQNn0Q63BlRUSn8IfKmczAeR8mx6J9hKt
GeE6mVTYoUs3BRtFSG7x+No2zz/sXivPY3AoACHiKWH32Two+fVTKZPGdjGzoBKT
AwCykX8Syf1Ig7SmqUXwAoDYVqMhFVXyboqh4io9MMo4XI7FZP6ur4kjoULfTuY3
1+rQnhDQYpD17F+D5kNSkm73LfzO4V+daQ/ICWjtymblzCNuqoyjOCfq2oUqVTuv
RTbBEjdBsb0RDonc4o3SisbC7Bs/ijgpmes6XGFHQ8F2uec373iOgm89dfTkmrsH
SnEJc+/kfoEV6wkSUJ5AiI5j6xD0K6c0PefykqR9eKrmSYNZnFSuHGRqLbk4zME5
4ofiqx0xv1InkxFX86LYCTzalmYjzUAe9FqFcla2dQSRWUHkYP0VE2ZM3hqATSMA
mkNIULiesbFHoUAG0FJgST5jh5pvLSkJtIfawhp2aqD+1RneLbWgOqyevquVeKPx
AT/9+XtB+b4H2obTTMKboFjsR/sNVPZf+WAqDVWbkRks/hrrZmqJZ9Dse3yl81bh
Ed68MnkM510FkUkV2G5PfjRivyKLTMUO7RtqUvy+FmgUZmZBs77k4j/EPBO/XZBs
FnLx1VY4iYcVjSqRLLx+jJvD9QDee+D6N7JozYPBSvSjltlrPN7a8Y9vWcLRdNjM
foBPqW8kpO+cIwOaQ/JsztowZnfSK2+zEouctFveetka4e9pq1qYS06waXd8pdxf
SlT0giPslXkD2aEI4hK6RANFD9xaW7I2PvZxFHZV0XdAQUucWvTtaRhg6eSZkEzq
0JPUKEozZxMArSe+SpPyWMjhpHSGB4NufNDd7fm/dp31wJxkNUIuI+RVOxUcl2T4
t6cpPN3FmCvDbWB5uOk1t2bkrFGW5RWbeCtr3QHnnekYCRpL3I3Y9a+WS9fsPdJ0
Ib+Ha5L/dxkL/vIIDI57L4hvXaZSOmTAh4AUDcvzQa/taKd2icj1I6j/LxqNQ+cK
MYVZ1csq6wP2X/tdgs/eOXC86UNHz3rzZm6pDCwhQnVBfc+lL1SdyJu9Hrbz8+3l
eqTZZ/i/nuDGAeKKDZO8fbrqJBhEbIc6Av9bS+5NB71jvARTNN3H84Wm1wHJW2s8
9b8bj89cd1YJj3WzZGsYwH2tgO3uo1/58MqYNPPfJmMmRwZutrJJjziW2hGz/qfI
8vXeb9mH4qW1VxIkYtx/suGbq3mnoXCo4J9QW6fQ+6DfEvlHUcWBpa9LRTe+0REG
QCDXFPT0ZI/Y/J96zJCzpNLTqGOzwvAPnlrI3c03T5B4778DYZ3FGFJ+mxWHS0T6
hWGbb+Ik3KPHzDh4GuNWFxpvQVFrfzYoPWz2bFS1DSWpoQHjDgz0CaqYLxr4FjZ+
PntaCjrzABi1YmsPfqTCHb+wsj2sEUyDSjKYpwwTXqjX/vTMpkUo/2OH4EocZpJe
aecou39fUGPbrqTGuUYKqSsYZQs2jNj1y1O8r4pULWowQpNqAyHUAmQ95/OZYZ+9
R2l7k0zsfdAm/ncBkVje957F0FyQsYlij4mMHARsYIUPEkx3T0jvptNPSMKW4Z4n
fid6SB+55NTneinpdO8kA3Bk4h9OPEE9UgwQHkVLnphy0fGFj2axoe6d4102iJvK
Hme+cfdtUl4+yVC6ec7vC0RWnpT8/ePt3fN0YX27dDpZLqe1J0XmtTzfgIbXWtTC
9mOGPSIjZNStO9xQLR6k3uA/R63BEx+FPCudj7Il+kbVgWzsgfLoa1l0jZwD+2B+
p9CI6efHMClfrcstC6rLkfxB/sgviyQT5NmR0UNLtfQeabE8EPhsOp1YfDZi1WcC
1sP4GMS9a0qBwp6BbCvya7bapZruJ0tMIimk+ZxO2zLTZWGZhO1TCupl+sCFoxU6
3SvbxVoArzNh6pBvx/CptSwDBKumdwDErVdis30Tzt4C1LacTTCNwfbvUdj8kvc3
NFoKmSqgH18HrCxaGLR+/c2s8HOS48wthfn6Levlvn2YZEG5omdamQMPqgWvdKxq
wNS/AsnJvwQrrqXE/saIt05npOZo80e05MdX3OFvSITStJP4UK5KhHLqss1sgMef
MJDM8FZyVi3ejsI1yeoYwLWqhEV6jA1iquv2gzj6Svj8h3fVyOALZ+suzR0Gx/tk
tIUlgSBHFR8xtjuVIrtgJiRv5T0Po/K5xuC5MEBwb7CJAlqynlZPjFvQIbD+Pvql
Jr4BBxysF8Cj/Z5HX9oUC7rhc7VB5i8uR7KHhWo7/QIbfmFHfc0/KzFpK5rbO+r0
NcQlfV7p6QxtHcBHCJqrWd1RfaILojIbRWYCX4Kx0oYhnBAwD1Av62amMuXheDd+
5yqVtAUynABRHoov11aq4WF005oAKfUYa3vLd4Q+1XmKJhNN4gRHX8BcpzqoZbzA
KcCPyz6roelzv/Ok0CZTu9IQYPDEmOwn/p8FPpFwEfVEz8v5UFMbwJlswfL9UnAZ
M6hZnYp3wrqWNEw8ybmvkvQO+mpe0AyWashGfDdOG37Jac7sR/ERFKAscfHimPxd
KhyT3JhQ7HWLiHH0b1iq0hOkIRG7chCRgVuNTGqZh3W5toa0/QDry0NlpKXfzcHj
CUui9b0tn5muh5oZkOWlsioqAWT/Ar37PVaLRoQbm+3Mio3cY4BDewJvECROxlma
jOqD0xDp1EiGq9PSFiTy0uzQqwDTq91j66ebHxngjTN/Q6eXnaL1r+6l2aS7wqse
73v3IpzhYL3i6e26QV9PRL0mOvvfnRRRi/Pj5b5kHsD91B/cSANqjdSJd2p3Hw8/
wH3RYJFDT6XYlsIKXVHUQsWEINzdDwyIaHpVtggyqY9rRUFQKgYr5ex4oqt7JSmf
0d4Ins5ZOPcPU2LuINgLbi+kdmhV9Of2T50UMUzu4cOjEnBzeUEjYjYS558gwZkT
FtDYUKyjZYjnlxxmM+m0ZklXkkZvTxmi6HT9evVzYWjV1XKrEzBDRS+tpaHbyK/p
09ib00rm526PDQAd/QGQoGETpu8gmAckjtL/vzOFAeD15jQ5S/ZgOssVVCcDmnxg
FgklVqMW/mePhyWYyuhKLXBdgTf9uPl78Dp1H942BEI5BXxY/5IFQ2E5IKRR7/ID
V3al2tCOwgef6/th/9yl8Oetdn96kK+UoSbFfOfGUfHrqTWYvKFlsnG8UMK0csmW
O55mdSthYEoEGoB2h7YkhyWjn1kkVZHevRciU4BIv8D0TOCmWT1/Tq0gFBF95dFo
kLfq1HPAbbimEed0lCXnzSr5/T56QtJxXKf+Ua/4t2ZaMJ32pHY+WZRjhZDLCCK5
pFJAC34B5RxlKTeYAE/rM05DmeNAUIv5TXhUyoJz0dn2wtmONOX1oeG74VE1HeE8
sKt7or+eZcTrV9WUQ+wQb07apzZf7RDsUYtPHfSFsspecmOvD/Rg0n5RDBjlhRPk
QyyEiM7vnBekqdXD9P7Xo4iNPyoYsOUzahJjgqbL6jgb3gCA0pOt79yVRl9gHA0Y
hMn3MapSf1SldkTOraVfTpQ40dvQtAuNXJUTCmbTNekcnAGKKfUmNAmxIor07PxD
qRsVCXKbgplm1DWgsQjFPEhpxBw6WwNRgAyH6M1ex4TX2A/Xrkd4arQNIWkDhalw
UM+kQGRjILO4ogpb1s8v4M1y4tXJ39x0Gg6C3Ra7IQ7o8W2ZjJVFweKmMLnNjqcz
T2m5IJ7AIF2Iy9VYOtfXKFTUoYx3dKd0N59QkUrz+4TqO2dmFRGJMn1FObMPBcSq
e5h483jvHU7GDIuJUg46uqY42YomUv8VbP9J6oCTxkQoryxoybSReqLjRIZBY8lU
WdkuwcMkic83M1ifK4uL6fFj7dRi0LY70KBAlKUsFAkFkU5b0qO18HYBUnviUWg+
BHR7z1OyHRcyQyA2Ol+FpvGIp0aW1JWqNaX2AszhNmbfAwTyrGNmpdqhHDcSOFbG
K3E8+76p38zcH78m7QmZSSVx1g2Oj4VpAHRxvDTp44/KBVTzsk8XRQsJL9t/5PFd
LzXCU00Md4K2+fB2Ud7TrFABpOq/1OyLDmKo2ulpqLR5y8MEZ+BgUZQqWqzUqtcS
ds7y0hqoXacG9bfnuV8J13k2K3Er0jC24oe4lnHJtMMS6Yb8qNb//+2HCnvyM7yO
v1yWIqne8cGUTNBEvabVZMImtGylJPlzONAR3c63y2xpmzSPjJk2ujrHAzK0VnL3
C0ztNIN0ll16ltkouhZUp+PT16P9CYXmLOFh8ziViPaG3uo8vcESoEd7n9UNQccy
O7xg6EYAM0wGOZ8zrMIh7fBmMkxUd013dfFFlGNoH5+loTm3rCjuwAp0yNYi3IoI
cyGIwAFFJC4faP1dL59yvgRFgaen+tswrdGa7Jksq1XAL+htEn/iVGK43KHOs1oe
oQ3GTl4waNy1sik6qaY3lTSqUJZRx2G/ZHPk0s7O4V7wvriIy2QSt9jp8q3VEkqM
m4md+jr8pdL59qHHvnz3vEc55sgxbVegyrNZBjRr1nbQQglS0b2irUa5HzgDQ5KO
J5ZngBOF8kIw1SJNMCeIolcrP1T0Z+gNiOcY/G5OlclvEEskBj2uycN2M14eKhWl
LD6ZxAH+9n2QCGL82FQfYtrHmXHtmQI/Us9fbliZ2P0GHPr6OCExcHMcnLYaD0ZN
eF3hiSYNFOJqfBfA+RgEnUwXagL0ktU/jK6zmaar1R43j3OHD+nrM4xGc0GTVYr2
D3c6flGLy0puy78ddYm8nQl9YB2617Q8cZQ6wfWxPz9dinpb6Ib+yfOkF1gY2rBA
1yXBwqF19wr45bXFVWneu9nCqQsB7cYVJthLP0sblcedB/GYq7QTuwsQv+0u+f5Z
tQZwoA2WKURK28AH8fzwcGkqmQTRBr3ix0CM/Fdxxrw7Y6Tw84hg0wdQtxKPB0Wm
KNRvNn0ZmlyjNikzIb30/rQsBXnJX/NzAvItU+2tgE2fkdE8HLnEMfxWTJjbXQlc
RFD8jgFbieafK9AZ6Wuyg72n/POulf84DgDAhk2Py4oOF38ByAWsf7R3lQbjdg2S
TQuhrPqwxEsGr6DLiYU7q4vR1DrqY69n2/eIULs50qgy7APBLax+t9ZfKoe+Cr3D
61Jpe7YvJYQVmpWozhRKCmigrhH1DEUlK+swLqHpff5tBEyEnLwf88Fnx1myhXVg
qElQYzf1d/+9BSiOyh5xn7+YB9qMgILDv9HLrtOq7EQ5UHSliuzVKfC+wu28Zg4e
2UTxfnvr4yYANEejTpiBoLEJ7h/Kmtsh+kecCIId4eW1TPxHKZkm9PxMacW4wFiq
TG7C0asJv1xD0dfF5qbh0tgYHYgOc8MSedbMRx2QMzIt4rO/GT2mmLYtncxvUV8B
imxwwxVZM9EeqkyvdcDbOPXiuekpbztTcL95ZlYIYdRegm1uF25zmoowBqBM+FSh
Oic+yo5UwIvmE6MZeNwRJJ3Pfw0z0UDtljDVlZUoD31JxbyroTQ6fCrmY/K0h3Om
VOA6lE9q1Z3pjAO+XV2NACVWeMSNPlWxG67ogRRlZ+dk9ePnPrzJJ/Ruo+ueWUKO
FMF4iB4EuAwe1lCSFvy95YR68EshDNDGtigcjJafT/vZzQ/XpcSh0ze5klFUiIPH
sOSVA+NmG48J9Kh1umWjQmNfex/+05ym80NHO8zGsvy12/FsViku3jgATCrFC1W0
IbP3wz9UTgvMc/Z/HvGaYzjabtOHwIlKlM5hSRItZI+IP+LZnReYqHl5+LKzLgPR
9ZU+fXbf+RY/JS7f7GMYVVh1RVCQMDDRAbCh+9ZSN+Y+EcwNZ8Ma1q8zqNYDIEHg
A6yzux48T5C9JDUmmMGPXJaXuToyrFkVEDZ7FgAJB5pt6jW05AICHey1OacwDKwp
pGe3puZVwT8M64sh4Ug12P2rP/wL2Ax1b5oRvLKjsWrQuLgqJcw94UTgaCVQ79Cl
TaJ2t9Sx6u57UOiujv1mxuAOSxA0bC9MgBE8AYmtzPo5fpXRNSAm7lr9PQfhtpoo
eI7dB8eSMpyokNiFiAaEbVk1GW8H95M9hmdNdUy/xIt0YbTFtyFMtCnoQPpbCzTj
3kgQGIXI8OeHsA5aXWxBoDvHqx3jju6H8CAxr1tDRFYgtvuTQ5428S7M0EZmXEwM
MznB5yUDXwBN/VCBz9cnAt5huFIYhKbhCDDoSUPmglIVT+peXMcHwi2GU6eRLZOa
xePLzurMQuxdXcopgDRx6lgNtGfMcMyK74Qn3/Ql6cXNFkjD59Y8CAHvmGOVaUfJ
dXIlNK0QktILiOkM99LdTyfRrfyNZ6IARYPfdb7OgWgvHmN432k7q477W9OpQSqi
tDSTnwlAKU7GJmT2uscl/j0u3GsugWHb8lkqaqk8egOX04Us1PVXtGfZXZNE47Vf
YTD9HBLREO3fVDRSVP+TnWmpvlUOksDpwyb3LjiovUKPKE3OnaeDT0U9NrhXcS9i
91jp8ZBJO9QBGy2n7+bZzJqCPK3Dk8cSW4cDilEZHG6rK1tHWqKoITK2aDvYMiEa
+rDo4Tv8ITgx0s8b7/DNrov+WaYhrmO4mWLiAHPY7KLgcKoKmLQxMakhs9DftB5K
0u/rRu1RvPRETxfKHOgcdBXnsRZKUa4sPR25MEv7ZgOObcFBPqCk/ZvTvX/gtxyx
MX8jafo3ttz1wmnOGGIHViRHu5OYRyP2/zznWh4MjoImqkail5oZjsswjrAI9bLw
BtG+AhhP6BKBNgyrv1nStBn8/WuKXt4HUiLqO+SNdSJxu3GCdMlwihgFNFlqTBpk
KPIddzqudKu+PzDvJEKXmt2sSx1o/QtJxOd+ZBqo2R6VKVPC39UCqN3P6f2oIDqu
p/iWnDFztKMAOLuHFdAlJg8ppwbPv8pwlQGYYaaB5+36gY3JWdS4pel0+F8lKkY0
WcvjuMf36SOLSqCLW5nnY3gOtgJ6o4lqcxk088mUSsEHajF7CP0Wy3fpBQWav/M7
7RLU0yzkZ9rDXGrUbwZXkQSJxghpjkWF00e7RXRSoXV1A2NWJ5TcE8q55obwRXnK
LQYdTyKY89qJx3fx2uIk2kb2NMsIGzMckTAaTseNBEUC6wXKIaXL86hMKxlZk7DF
YrTurfDXsqzdPGiBW48+BnuEsBByGJsnZprgyRE4aqlproDJIESPXu9f91w0zJ64
j72PPM1vJwbIzz1ldBXfHqg9YJp1mdjCh7Hd15vvmvqtwzdcKqZQNADF75YUbaOB
kyZ7eOqtryTPzknkFWeuSTwzTCHzzsJ1rsVgIqIdwY77RewtiDWDfYS3gtUZ2rhK
tIqgyOX5ejwwpC2jkUDensNKJ1C2h2KUKAevxydprR7oBz3KqYHMA9FtI1dXpRdE
0thiVscijhh9TfQ2GLognWnDdKSEnO/Tv0hpr+hwRWGCIvi6XZ8oGOiOCtL4uxVG
bGJSb0R06ZPuvIezmf/dnwOn895Q7AaPPgZTuGFif9EL4yax/EGFi81+mYxTW+zZ
iNQLGY08MG+Vgj123odfCvNusBVw9WBWlj5uS+qetU0w4DiM31qO43Je7QmsWlHo
nb/Ij+7javkkvcN1QxLdtFYvnUTgGuMMf1stAmKHCHt4OySSBHdRaoXybzhJpPoq
T0sdR5sZ2mdsz23BBUF3RaNreDUdDZT2aO+QpASuT9YUJCt8WaVb7LHvH3HyRXE0
CYHbWJ1FypXPdW8NoNjqSmPL42Giq+VlTXgHJ67CrEd9sfoN+qBAUHxrjkmC1ZKm
eXKC1SNPNWeTyvvCEhqxY9QPkYMDkQSXr6Es2waPQMCxXfBhKTgjHoQIErDDptIJ
zrojN+3WmbwtkfIp9dKLHZVVSJ3eFKEbnc8f8kfWPFc9sh82GHmtarxINoKyZT9d
eG+yzG05lWeAU90JLhVSX0cV/l01EkkC6izvAMTHb45lbAwmqWGIR7+5SkngIBjo
UeXzgL/K4iI9dk3WYvFjRweHW22Vj02WVx9Eln/T1Ys81zr2BSoukgbUX1VswdIt
TC7AAcn9qVx0r+UyReY5QeGuNfdrBWzAqvOEqBmOvNhqpKGtZSWicHDlHDHIlmVA
8dC8KFwPUgk3NHE3RK+3RiAHfYqHs/1t/tJfyxJQYxplk+wtfe5n5dcJDeNa29MH
8UJEsdAsN7mss3sO5SedMLy+rSOkxChLlQq5JxVcUWOWInZA6CpnPQBYvwNrJvWT
zC6t+uAyKHvcrpjV4YwmAoDQTI+qboPlRzj4BerxekBbHlMg9bpp9K/NCjez6wLq
h5TfUtXDHM4iyUvc4MYHXWeoXd9iEJ5YgoM4WV12RhGj6+UPXLO1k2e5VSFRl8Xn
Qk32lhmQffqdm0NKvYY6ek3BFj/sxiYRONyONrJkmbnZXjzvdBEBN6zXumHXAhKZ
JBct39bQCxiGuCWzSi2WJfHKlg1oTuhTBfYHNzXSFfi0n7S5QyrzAqOt62DENDVL
MuLJk764GKJfR8ZkBWtCzR0eT95tj1Z8PqKPvypIfurupW6hzqpAFr/iADe95JqB
xMagVkOoBmghNMjjRn5m9MsohSNOgfnCuvspKv4KROnkXf241ji6/lqpoAOaPdrq
353QbYf81y2eD/JvVhlwD00zapGpBT7RSxDQZLpt2M0GeLrq46LRg8QXYq44RzdK
8SJQT+8ahQF4sK7lo+UG9Nkrv1FbzH/k0lz0y9skeG95Akzl3cnvQAkY96NTDPkv
ZrgeL3RqiAtxowXj9jNJ0gO3SMMBP6b/ZjpPjGex1tZ4JtrlrFHpQZGUo7ygh5si
pFim2SKHL2I3CR4YvcJlU82ZfhzEJ7rcYbjocQT2w3cmcr82rxR83zepu+44CvzF
tFtbQS1ALAJyazQnmFsmUwpFzyyxBchEIwDHsA+7HRCXvR5MFehotPZtABEnCD6M
pZlq107Bd69KyrTbsmj1dPdcQNJrxwwAgJnDCcAgHJP+FSMGbACkRehhqH6donCa
EMSUml0EawFRVr8Xna/jxZFw7F92xR8h09+Yi/EjckzI4qHcMBjtpHTKjH4fQEnh
RMxDEFwwiakGctel/t6WrBiTjqTVHf4Z2AX8eQH+3GJmT8NzJixvEDiKL5v//65U
JznzJPvXIeN+UIVqRX8mjkuELT2Dp9vZhWdB6ACr0pSYK0a60accOCuXWx84Hy9f
VWCYU/fwMQ6Ox7WifjXkIEi+M1dZxJVRYO4IaDjORBQYxYtHbvsSzqNBuSk4vaSo
3UCb3wzpV4w96QX737zfu1G0GLD9ur/B+IgglWwsENSljlMMv8zWcSxY05Se7btk
aI5khFrtN5DDe48+Be+qgWmF4yoePmOj7nsKyytD6m4Xw5+5NYDIAtnNtccUBSpE
IdTdL+aLWzTLSUenO9Z0kdus3ZghuUVy+clbU4DJQ8apMY1U3If1640366cfFj5q
9z+rKxRdEs/maY8xbMIbc5FaB6Y/fTxQ1D/LkRTdQpJUmmrgagOdxqot4sA9QZSz
kX4wKYdtgSVHnSuLWDgbZPT8mQXL5tFmbqCHcK7v6AokB7SgZjkV99As1wuiTUhJ
JGHD0sMBuMWxhCSoXsaOmeOb8wFzvdFHU9N9kDQc9PLf1tB7+S3Bwn+U0zG2V7lA
ucezuv4iwSwuOhcnKStOYox3YdcqgXgoU9ze6PRrzphAyb3Y8YUWdX/K4Y5xCqfd
CJZz2sbgxcRCCrqa3fBcWVXBcaVW9SP11SLUPUeNPyTWUFv4thv7NmTlV5y4PteI
zJXHrQzfkfYazK8CS59LvgY7bcRAr4zMV2m80fhmeamkQCb1wemI6qyEGD6C0c3f
PJtxzq+4l7kRSIx495eyrRDAzGeNVTZRSc6F5F6cJEFqsTW0OOEa4LuNUn2sd7Kn
fsNCfpJqXSX57ewO5dUFDC4LHpH1QKyIv2GQqeaLpGDQ2KnZGGuXi3hPhoSGb9lh
bsV5CYlOStFgIws03EAN6zSvr0JMsDcsS/tmYfFH10QJFh3YNwPaH9IYFlJPqp6c
TBeJo7wWCd4PLzQKij4w1AmvNHLiWH8PjcSBvzh+meR8vevH1gwEfOTDovd9GQJ+
ETUDxb7pupZcGZCnXba8croyAhlsx5Vj07fNhYD8MkVnnRYUs0PoFt9jrQh1aYNn
hSd/aACbGam4Qj4Rp4TOb1ntqEMLrjjo/d3bjwWjpwk1/4WgOqNIxcFFLnHaf3ID
JrVO8mQn5B42mHOVnHrqR2zcSwGLSF6VySQi4fdz+6HS+kYwU2+CyidjutIDTS5F
0CnB7Lj31qMufv9cZqXfjge4ESX46DtFVmjnilPoSI5sKQjJTZOkTE6Z6pCXtFO0
46D5+2wo146CURRjhHtqLTQnMo1AJ0heacwAlO2bQO6eL+EiOhosU0iu+A/3NIDB
Idh73yaJbispgd158915QX2ntG9Gyarseynq6sJznnel64gWngQfNWv6kaG6e3Mp
oiSTi1/FZA3tGzOImm9nF9zh7qsY58f/dnj/tOQENA2q2mV4OaQYjDQ++8LOSHeM
FsPGwOO8mGFjMCxwRIELNFuVLImY8ZpQdOZVvehSXXTubV+dDXIa2I3SGKEEkeRF
+WquRx2kGqS1FZlwKMNsQ+i/AogpSP5iOGMyPhaW7sf0JKhnu/b3cZIW4+ehLiE6
fnRLheb37hTnSJugv85aq2Caxrqa6Qk+n2B6NVyD+HFRMf23CABR9gNHcNnoEaSQ
v+BvdW327Sw9v87NUjiPXmDFIVhDKYOKdminJRKaePZmGDd0zUpj55SWCUkUhD+V
xhwlpBhDLwwXvzbXwTGpVydDW5/cExFzmZaGfsonxtjpimFHNadR/+sQxlfib4XD
bVODfBA12/3zS/pfeyrANZI3MZ1reX6+kGZj0CdPZJYYZCC2WhAVergdh+BqoUmq
2JUJGsDhRZAhTkZ+4ihDPO/vMSIgPomed4gB/j2eFKatRTi/ylprzRIo5RPY7s+Z
ykIg2DhX2C0u/wOLO3eX1siiF/U/n339Jm2E9Tb4IxqkmPCMSkbVRfT42dyARNrl
I9KH9WV8hBONnoWndhsqCb0tWv2AMDSZO2Y6SSqLn7wFEKPHCNljKv+SPQSWJE2q
576JYzL8LRPnk+FzEq6xPJ0kQ9wSBCbteur8kx/b2zc8ZH/9xrjO5v5wy/f8eJcE
ErGQX6SPIewYyg5FxRJh9rxqAWZD2uPL9UgPzrPfIboa0N5o7QVQt0OhnS0clk3T
X5iabBEt0peHNPvvkjs68WXtr3bxq9k46gkUmb0c6q17Ll4sJQ8A2q3f7MXmek2p
tMtkJXJWqcvMSOhToNRr35TW+jssdSHtCc5bcTgCrE2dBHEjqaLnqe1BkgNq/8FZ
RXnG20mrILjWELKhuxeBsQBjQM2v0aIfmhWP1bdb2mA7vzZGh3hAsR+mTM1Kmncr
Kws9BDjltPuKM/sp+NWKxhvc4gySHU+DAtmgtBmgRE75N6Ume3XkNbgbxRJszQIv
hpEpl4u1gOZfIBTrWe58MdbYs6tHls6MB9BLn6X5CKd5wl0pRFbuCD/f+fAzltfM
URwLiJPoGiPhn4F8wlgwfUBPbkabw2QdejKtLH4oXsF6EQBInB8OsQJdmcj04BFT
m5t8FxCug3/UOCqnruEXhuhvfSf2HVh+1Jt85b4VrEWDiPPKIcSqw+otkC7IR4iE
Lx64l20nPdC3ZjU6hWlgd5n4v8jtG7la2gO9a4tEPWMojgO71nzz1gd4pQYTWHh2
3Nr7DZVmieXWPCITjkfhdP06DR9UPSx8CQRTZzYzoKps/YIkf9c9EOqTq7AGgzkQ
2EBlK6sJU7kwLsMQfXwP/MjzivG9cqee2e/ha8T2rEJGcG0AE10vuc8188iEiCMq
BZ9EXvkw/fO8JjHUvwKCSahvx7vwocJ2m9VBDGak5A+ykO2Bsa5f0hXyLjSzvcrb
dN/VTtm1VxiEwc+BpNWSda6MOCKAWtLvKCEhwfRS/ee77blqNfICPkF8PJ7DJADw
uiWHWl6NrD+6wc+sgc/osHklvb0uv/ENJeJajQyipAgD7z/T1Z4jhWrtaSXnDZGZ
XYMHif4Q6M/UBqBepfBtyA6TSWiiT6k3sGU3so0AL9Vso3Z9BAPETIwe4umyBIj0
v1BN47p1Y4T7rMhQNSGPxhVNEDz2L2g+5R9BWcMDsR0fKTu9KomrBNKlkGgwf784
AN4Yj08dEUaTk0LmGJmNcjATz/jwfwSKodRu8uy2L59sf4B9HVgHGe7arjUZFOqs
3scl5pcx4vBnEV4V+N5dqxaOFuGWdS4YwcbtWsut+i+nhmA6xR83rvZZrfIVD5DN
v8an+S9c7mwexbxbeNuWSePRqEAoeR/WFn4o071RYEbcosKLZ+6VWZ3XoiIyKm0z
slRWQuaxs4oHYX7WlDk99tHEUkR+b//1F+RYL3ES2FQBZUgKYN0bOGEHdiliDbpW
d/lpKGNiJnfaaZ5QDma799GQDnJwawGJNl4avyhOE/OFyYrV6gQAQ5xFdvxXIqTb
DEDqheai46tZ9LD7T3heL24q1ohqUchbRepBS/tmHGa0Nzc4CRfxVdfMCPJhzF9A
j+MdGhBEIXnXYk9dYAXZFlPvpuurPHo+FMjbLnIhbxEgQ4cBO+b59Hb/DkRuVi99
r8m8ycypVza4MYbF1okgF8sHqkAYa6u6Vu6XCq5TgmRntaltX+BLwgmSW8B1cwNN
Pde0+uJmDPQ9zrplYjbAaftGuwFyaJUBSIS77l0QjYCtIetTL62y4T9X7VZHYce/
wsRfCGknCBLoU4eSe2KrPZK3k49JYPml2IYl9/SBhytQXX/E6LVjBaKnWUVj6lJ+
VmoNPOayyn2HpgLAEtmPhCR5fHwxTexVcdtnObVTqOvr26OIe3C+zjNv4nwnKqQW
9dzkIem0zEWDdmarbh0puT8X07Ok9tnbDsFy4agIuX6Xmh/Ziy8NZXPucvl2Cpqa
kpDRZxHZxT6EX69P5JmDrCIvW9miIAhVKqqO3ac+UW4tpwU6IXJahuYlqB59drW2
SCyEePiQWXMOf2pdMK4UQF37LCBQY7PMJx5bSVRHhO6J4ePwYfMcfIWyUvM2mlj8
21s3w8q6brx2syVY0pQiL05fab3L3+vNS0GGTKmHtYpyk0pnjbWmuQpC+rdLwXEU
R/JfWfXuG/NPku+Jmka6t4bwi1ut6+5tx+6a5tdDo8wuwRGnCFDkD79GPJCNPZoo
dDjQ92wpNhklpFZVUqHhX7sdQf5dvw7TuLnVJVhlzPKIHbDeXwnmcytiszsNxUZ8
GPslN4VW3jcCeWQKciFAO1nklnL0WbD62ivil54Q2st4cqEEhv0rf0wqsutlnXMf
hnoEaLCNwBx83O2BuS5bOcN1AqETNk+cCo4QS9qvcNy8KyDMhoXfBOfRy+L0o25b
3gYAK/0gwxNBUxUOfO+TN8RNaPl3WJ/9Ak0w5ecmju9+XQ+h5e8ea4xMWNK7C8Rr
tBpx8yIcOpO6WSVx/klbkXWaZ5sDqdzFH0VDKJXdnurW2GC5lydjBUbv26Wezfg0
0wBXEN41E56rhh04iOMa1hYFFhHroiUoW7mFskdSBoZNNOnVuSVemJH1+4NknEM+
MiNtFhAsuDO20FyjfrLqeNKkcAtzFpUeyuhSRWFRVDKSUb4TwwEptgkjF7GCN+1i
CpljoDkKKgqjmoaHeUxuu2CtMHYcY4f5ecBTtBbEkVsadpaapHcQFbn9yLIztq6U
IZZzVAXRKXIbN6mYieIljTrN+jPAAwFHl7A9x+YO2XI9ftBg2OFCSIUp85QVk8a+
dKaK7UWYhxl/gdjyZn9aLBOQ2VTLinvLdrOIlh9jvP/klzfbsOj6OX7RS2cqhozz
4AyDCCHVciCoTdGJj59242tPs6oCZsVo2mFmlSrxG6gIfNqt+U0u/QdGEU2dS8H0
UvdL4kp3dowMdRknTlCNAq9BSIjJRyTfFAl4aoktxoPQYpittGGeM9FkCjdkIA9F
D3vNti6hdn7kQLa3IJMexhKHLH5XCWZLJFZfaGY6F36yHY6DcYqHtEs4ECKwNyJw
nBaN1z7jlBqfH3cQl7noTw1uF/9451FYalFermUwRXhUtQnLgRKaih3zfDDyn9Pa
KKQoYDn6U8j1yqlPXcRm0Oa3bpKBzjUo/0kPEd3DmxJlIyoJRVaQbxQHLVFhFMTj
FBLhFlK8a2msXIz2KedG4mXVFlXSqkUQyPvDa4jiWEN3zavLVUvZ/QzxB75PRUX+
KUENoVtipSuOHT20HIHcJV2tvSXmmARFNjpaDabQEAdBUfC+U3vWUeaQzYWH2k2K
cDDvPV4r6JWoLSoszOxz5xzIH4JdHgWNaSIoSNptDtbFW1heOVWdfQSwNgAapGco
KAi46IrIMciedco2I0X2oyvTvpNCTjclnD8puKu/EEFD2F/MhpeOXxn/6SGFVnvk
p1m5PvvbR6Ll52ss9h9k9qCel9HL11DSJnPv5Csjzenq1IvsJplSSrIcjAzO3U/L
FuIIXSvR6328x6XbWSHRalkKiTDF09GzCtZVxMM1mBAwwPrXrOOzy0bszRL2MttO
/Sw6tOgR2d3ZB8/LSdlC+W9RRzkQua4hQzmufTGaESjAqvDKt+kS0kSAwQ3aZfdN
tavn+2ihaAQ9X+VGPV2XmsHlK4myHnqUAva3leRLsNyE62TL5W9o+wWhLtVtYAlT
GvG4g40yvJhHz0aUPsb2IYc16SfFeTMWkTiQ8rqeqceDuqBp3ImYFyLEhvLv0LAZ
erNf8BYfABBsVr2tlzPEDF8QneXmb85Be4dHyZAv75/SPOe2bhb60MqFIUxIrGHQ
F6isGjEDXsGXhNhOwNcFvbpawZTs4HGkIGl6GXMif0bgOIFrRD5rLLlp2pRlbmci
RHlhnBxoK2W8GjBDK/14tVIyaz8uz/tSVNM1NASnS473z8WxqwGB1mvntiIq7cQ4
CdV5Jq+omzvxyZJgE/jTfXoI2LQwLmiviDTGaDgbydYmrtG9ycdT9ElMfnqwWBbL
WJ7hggdyMpCSQ83x1aEEfBzs8CZ6OFLyMBUd6NqkltR9wQLryLo9jUyZekwkfGLC
tuC9IKOs/DToTB4ves5kj2uYpAaGX5Bu4Ljn/E3RCwmip7jT8lD0ozpWvO4QvgaU
zQc3adr4pfqNxcURVeu8AsVdys9xNSsFUc9Lb09oHlKYjRoNsSfrBhFcPRtSGjUK
rV8Ul4GK698aiP/OgFJhwqyDVElRZdPaa+jkwx0Fo26KiwJ3P0MQU0QeKlc/MlL0
a1BKR8TVpYRUWP4FTBVkwW+HyS1euoyW34RtZ/9sB6nRGbTKgzdayyywNpnMs5JK
/cetJsyUW45N9p9f841R/LC29J9Q2Rn897P+jQ4sOJlGSSrZnNkfxDjV/EPhEBZ8
2hxux2zHsmGnrv7Pajkq3BFnv+qN3Vjnlb332/hzDRD/7xUqd+uaJ7ufKziLg+8h
yxuVRkO0XBjEwYv0sRQexx7uFhL2xTuRRgXv/zuK/qO3RZ1QM6r3z8+fjbu09Vni
RS1ywEo7nRh21tAr7+gdWKxzAjERNpvTioTSC4NtbQLQor7XzzBuTiwoLrn9tLIz
qg9ZWbyUYm+z1xz/yxgJw6MpSLApEPGRDEJ7Z8KIYBOPuEg7Cppq1TvsGv52R4yi
LtSE1uSV/16TJGfQqWRNCuQEOwNFXZq5/V+2JSpkRSPgm9EQJfAEbyL5hPVzpO2M
jWi6VYZo1RYKdSMEOpNLHO2kNkoLopjKgMNfUbxutUAs17DZmRZm34x9HTcIrais
yJ9tffrOaZfnfWMtYvLuX1uxFwzHuOF5eGiuo8sAu465WhD2sHc7lQIDWRDWJZS6
iUWxojOIDDXjVLVNrIo+rjEGl8ZplE9cqTQ8u9qV2C3ukx6AqqDL1/Nh+7nErAU+
F3md5l5STu9PWj5vSYg984jh+6LhAbqkAtHE/DBtkpTR5VwBZwwJmI61DjBLV+3t
/diVPdcEY5F+jxEP2frkxik/Oqj6IJsrJjOX+nPjAXAQlpW1uDgFOBNqBz21fzf6
AtjFidQ+HbyKEaV7Xex5AH0hSnfnTFPm+vOrufd5cr8c1BBXaXnMEeAD5MU/288K
T1nZ5UpuzdOslJZzWhvqFLR663mklZTOx0Of85dEExmvV76qipoLUxTSLc9zfPMb
SgT7w4Vi6laaiDzQ0F/kC6lp+yoW3w9F61HjGUeDDLmcM0uPEP7Qn+g3PeO5wJLG
M0/yqz8nydDotH5n3qm25nPi0NZw/vUODP1IN1FJKHrCVxSYGALgbjvrVF/2oV6V
Iwl90Jr40ko0qfaBapf/JxV0pDhg9lh/j7zgj5XUSTM6kJMrdpYYXxP3xP6ZicX6
XWbJwQha1QgBsa+89MHm7cwbGHGx/D3A2xL2j73rbzLMXUdo+HTJ8gc77FkscTC5
puB8in944hDFn/3AZ8mQCgABSvbXmLOUVv/YyAK9LLK+BLJYT77as447n+XAdCgJ
UnBM6bOe6yGlxNA+p//X910sdh7RGBOWYHsSnmyJYbfshDFKLtYPyaCBwvfHOG5x
Xj27sSIfH1oFF1BMW8vXDbLpZJeLCyvv8R+eeYGh0chzTFHCfp4OSWdNzgqmrUQ5
bI1jbqlfxCX7DmlwW+YPvar1qzMfJhUAG1Yzn60wAcpPQpEobgsGEGl/QgPz8kdh
B6LQ6RwLAFKcWRM5DrdHNJV7/kwLRgvfPsIbfnQPfty+1iHdZbua9eKLD1SWsC1F
TL0J6g46RNQVblXkZACiujkLqK0i/D8r8ZjLdQhRatVb+E8GeePd8lE+7/KrvxV1
WYSpZrQlVhNXL8aFkNFAD9jAsl7HWIjZ5vgx6WDMzgaIr5mdSdsvOaDf3a+CAyy/
E66zYeYfDhWzTLD3hH9YeAcsoJxggoH7payRwukSYNyl5opTq+jrXJNvif3/U+Ou
GKin79VkEVxGAeFHx4lMwLnsoD/UudeElazlFh211sbikWuUetS5erEsA34iMOFf
pHVYW7PKtAZnJmz8hkRiTT9xzmDtPE9bcl5NCkxqjtfoHdhlCQ6jHPJjX1ihgNiN
trRBU545wsQTQXQb4QwgxZqGS3kqMdkdj6thRpINYZqz5KU/Nw9CVdwKgdLx9/98
BYY8yE+PoZQiDYL6R5mALrF9SAqcv0ezskMfYYBexdO9Ztqmh3v7T9yv50U3kKG9
pUNAvp0wlX+h/kpCGx/Lggg0/OWYRxPar6jYPvcnRuqHVp6zCQyiQjFiZLsyfqBb
OWMKgYpD5BdUmZ+1Xhw5WcWOpFKr6s00TCBOxZUTSfB+69zzLyF9laOWrLG8fI5u
rGKr9lUTWLZ5wcksJezW8qPwVmHud3KcvqhzCm4AkATOQYMTzZjI+sJv1mIhNWmO
vrGtLC35cpwnd4gN62WN9fYOju19rjrrH33LQ0yPFptV5OznyN+EnxcVeB+C1d6k
TAaOP6XoBxOBqj76AS9glD0m4abojB5VNJjgWcS7oJ/gLqhrQRkU0V/HQ9V3wSfO
N0Yt+yImgF1SpEGZF3YmpO8/NxSbAd8hVJJep74psjzD1hw9u9PaxzMVYWPjdBmx
OHWcstFVCUkeusQtra3l9HvLZwoOSwz66kwkIofkJ3Z8vuHmgivzqB0etT7ebFtC
DG+/9dSEwxEMwUPCNRVMC+IpmiXvfqFm9OyGGtk1cJKjFpwdHHS7Dv6afl/1sov9
U4XA0Tjzgx3fT43GjGekAN39d9Zx/KJbAP9Jsk+NuIP2H/83Kfwnkms3fXMKdMjZ
KIggFz7qsSrky04+A9UgkWEQFS8JkuT/tn34Oz+ks+s33ab/Uk41ekGHmxpotGGz
VMQl0zWkQss9nvMK65R/BMbWyzl0uOKOpoeDj+BTbQ0lDg8ry6xxiKqOXCFJRrfP
HFbaF5/kk5QSgw24fNTo8leQe/AS3NpbEPTLO0B6yx+NtWKW2VoYEu2TDzpm5ra3
s2uLQ4irQlpQqnrW1SP1bu7x4fVlH7uAIjUgGL5h5+N5n7mhGjB44O6eZo4/FGH7
tIpdkPzenSKGJ+99N2MRgbkjo8SAbI2u4JPRIWiLWM4bCY0sd1zmCBQ0IqidqrEm
CLnMUFum+WJ4FvJxv2S1FE/a/YtgqwYQd3o3Ok3ysEupp5RnNluwJgZoyhQV+odq
faJRPlaMPEcfsYj+8x0jhp62YjzrQuvo6tKoaCvEUItKLForRMhUVcB2CVdSrr8t
cmKWfvRLRckGwsuJf8HyNVo99c3TYibE5cOeT6MzrmpifYqNpXUj7ajDptYjCb3/
XOYyFgRrXXf6GWE29qp3Q5MKfRhRwYmi/OUv8Id2onMZ10cCNYyipdSfwkPwPgrf
PIWs2jpbRcpl8Q9kPScpQ1IYwyiuAGBJqlN4uzzvt+1XA5AyfxAmp/VxwIdYrXE6
nwucLGkwETG/BgROgjgG+PMGHSs01VqgIoAJUhrWIAwjKCMckKiVHywvFHAy+q+j
Nfojp+/hdcjg1poW58p8GbIAeGyWXAzsSWrokW9009022MWVPFk3OQ2lAl/Pn14K
2FPcSOOEp2ZeLgX2mg1NE6zrAFIySwLCJyjA3pY2henAYEX2XQ01GfboRoKq45U/
PGu8EZBY8svo6QyS+tkhbBtUbAoroRSD2fmXoyefpvXr9Q50S+tbydNv16dm+LJK
bNqLnluh+TkJVlaqH7CoBDjI/e6i0UGoJAw/ez4EulNcDN649NwM/Qw4Ix5he3vA
nXQMa2YlJV9ikUJ7y195tqBYwA9XVXBOEjjhfuN2sIv+B0YCGbccomLBy4Il84Ho
OYn92HAALM3DWhAArBAsYvdK8aWJiE4ma+fI7xhIb1pOqs2f5PaFTPJjcTYakV90
eGePhjl6mY7e84qOyTUc/pdon4bOfrUi453+YLIyvsDrYgFYbx9dXED2jTpBxr98
wV5en6JcrDycC8ThnwETNt0d3Gmi3ym8HnfRBaIZ7d/Q/bsEzEBbM55n+1jDsN49
CrhZA+7+0Uuj3NmvU+i4rgypECt2PzFp+HaCfRUFqBG2NZFqNFi+j83jIpFhf+dp
k6IywH8cFSvMG8mEftILMGciGsGkq+7mJY41SGhJZnfqYfgDdGSl+ud2bWNI4Wvr
WCZ5+FPsyr0viBjRz4R4CH9rntj8yf9LHo3oWIfB9aI60uIlpgaz0ugRmRTp1hDE
X7cM1k8sg+xAkxs1PZhOzJuPG+uwmqHfvPgTv44Xu+tu2GhdLzHVfQz4oiNBZMh7
mDmOgx3kFOzmhHxJc1/QA9NzECdvhG5R4Vuy8ixrbqnh4L9zE94JkhIvefWW1dOE
AARFwBe9yv3+Dpg9V4f4hnQgNPbe+j81TmnBpkHRpTJx8xV6DwTdtSMLOWoOnCuB
1/cBVoMbPeKeom/YmyG9wWWVlvvFN3SOZJolmJYkaYzvpaBb7z5neLSfwEBzsuWo
Z184yHIg1eoOYKNvPo01kuTLn+GPutE4rFZS5tst+eTC54r3ph1djPVMMV11AuQJ
P+Kv7U38hSDeQykwKOQ5rTDt4vL0NbJoIPIXPQYPpj7E3glCQhvbpSkplGOfiKPs
9coazBpK66aPCeJX4HV6CjTsxXgiGUZVXvhnqIyzE5T2k+UFctKRe/TlVxq5q8g5
RQdVRY6xiSH5FNyrdc63fbTfYp15EAYz2wRGSBUYwgPNvJ4cXvpN3xIW4mC5dh0W
1Yxy77IwnqJAJKTn/7Phs9s4hoVLmkpYJjoA/RnmMxHXvlyYRamLPkWxKIVFvBg1
COp75GEPXJvCF+hB2VSGfCjgWh66yfNEVF35Om6sP9CgS6X3VOYhhyZdslJJEutW
NBvKRtcNtRRcPNzaFkuakbTHQmXCQ+6klGnSJF8jDWCXdVVVFYVQ9XumuzxmK115
Zgck5KK2DlH2nzhAIC+ZI8fNMiA42XR641r7+1IU9iTKF4W26HmYqzQw6vs2kSkB
UGtB08G7Nkm6d92AjE79Ogq0gY4jEDJkztHDTj46MF7BsWj9sB9BGKN3bKYOiujE
Z7x6eGzYOGIagPxzH6mJHvp/AgOHT0YsJIYvBCCIRbmpxevss4ltC/mJBGv5d9BZ
Fa79lH9Q58DyjLpT/Q+Hw8/687z5wqVzJuFfHnLisi8W2BT25qseoA7A+fez+Gms
GwAu5ytTwObsz7IjFK9G5b9X/RK5SCkHHMUpDWDo/qgkx/3c34k+8V4ybY/ZguAz
xb7hIjt0+i9gqbrH0U4zHkrtkX5e1Y2xAMfFp6HiwaMOX2TZObk+Cyg1+htwDDSN
bMkJ02eX+sPDq1Q7C35fFz9EAwkA9ts01iIZYtdOeq9yRsboEo4ixCLv3Tr1GDYV
6XkZfZo5O4mOqbvvSn52X9BidT6C8yT/oIcX2rPsFXCfBSed5fc1BzAsOYpJiMIZ
vN+i/U6h5cTOXo+HNaglq8iYL/BrHDwzYY+JJh8mcnIoKU6ZV+HvGA830jw6C4fI
5btR6uR+Mz6RfWj5uBxCe07ejqmewHrl3zngU05nPGOCjqIdk+2YYFp00wYAMP5g
4ehuXRcBgQFHgilW70BgvtD2q6V/HkovFwWAPOIgdR4+wzW3fTOxePOmkAM0/+en
sywEkOHdIBHRKH7Vmc05F71EBwI+jtDo8tAnT4JRy/VYbtxpaCCEB6OCnbFhQw1S
sDn18vbS4ng+94AmFQHh4N4dxCby+xcSoMKAOGFL/jnd3uyd0b7POX61wNEg4hU2
L/dWmIoAlc4cPhmiKL83kOilFxSXsGlXijG5BKL8V8CdFuM2vUcrCKOEqV5USATn
ES8y3ot9DV7kwRYHrX3OetYwG4NSsS/1joq0hHt1/5dheYI28WrW03w8wkIMSK8g
TO+N6uq0c9Rss92124tRoiyLjoc798J8QzhBCDAvixA9T8m6j4pgThJ5XWJOJqpA
ZNLvaECk9JOHG2UQpyOn7Grc0QEP5/m+h30nj+wIu2LQ5FskWski6E5p0Y3FPeWS
D0p/aLP8cRTnZrbF8T0pGmGUOqyODYQihg3OiccDkdGHk58cJ7/akUbe34gLln5N
4mqObqBPcl8IR7zXI+A0zCiT/swWiincK95Qns7T/+1EasaeHJtP4XP58kYDrB6Q
jlWILksXJ/y3x5omkVQLMzApPzdUG8eUzPA66PxtwZbABUVkbAv9XT2bt2F21H5J
6AVUSfc9RozlLG82nsdco3gPMuxhoBwPNZei2NTP4glz5CWmB0k26XdVKKB0yLKN
uQZhFyWAk+NwxWt6cThztwznlUDS15X8fh2iW/xQcN0JZzczCRl91xBX+dd1Sh9F
m/Gc2wdoBEPZzNuG4/4lmeFS7SnnYbPBGeSPJC8cpyZns+4npCNT6XZaR+6o5By3
Yp5b4buf2xlWC95kKCyXPStT0UwiofbuA+8mnxlodbF8EVKnIn8CvSldxmNxT8zx
Ao6NWa/dNqw1Out+HMQuwNKjHZSM/sQGJdhrPOgT55Hj5c2yp521xNKfhjLfxpVL
f8DH9CC2qN+mCQ/ShHzm9oHkLOBHFrusEGv6/VBLB2gu0TvQVEgqMcDxvp5TbUlA
CF/QB+AmPv8PDfYNEUFIKhv9lsMIPo5JsKe3+oNDplaR2slJLVRD3eeADPi4orxA
3oyphhzkqqMxX22Uej3HRL4qKzZInJjD3IRsK1kR/VcpGWNEZu8CI9frCOoz/i+j
8/3QonFaDDtAYpdCzXNu4zCnCUJc9iJa/brdQq63bMWuVj9ONaH8x3+11uNBT09U
AUkIOPMsLmKifhntF2g3dl1FOr8kCNHuhwfBc66PJqWwLb1yo7OhulvTJdEXM0iM
nmYKxMhoclU4ievHH8m/2AUjxDMTlN9TO6gu3olnMKzlUlGaBmM34qngz5eMvW9u
uK262rL/gNIFsRmmOlnECe+a9XqP96lG7cAH7P6ewwQ+Qc3k/+TC6IQV+iVHmues
kflEqrOjGL60wZpaEQb9vZ2zhqDMfITOVdgKhaTMWWMZnv8AQ7DFlItEoiEPIbs+
uqr5Rfi7L/gEes4Gq8VIyd8IIcPu8XH687tnY9pb4HclllgYGAaLPBBkUC7ZwkTW
4sR5jzK6L37qcd3QhzHneZHom2iA8GjhwxxNjNuTFR9iPgCF2ZQDn4QleGYQEO5i
YHNDEbo6GqIFoG58HU6z/j2EMnW4UtETUEVj82AMrD2aQCIAxnCQ/pAdQacAAk2X
XSuWDdrkz7jPFYITaaLAqzw92KejtCJXwPKKlh2V1EDYrV9JtCeGq/TIFDAmJfIr
Itro7p6gT3xSQ8xgZ0NJbGAMofdq5JkKqUY752tCvexE07vBnkswwdlgBR2FrB4o
gV9AtYzE8lTRwR0H/FC7oNq3O02boRmipE8mj3vFpUhKz7V1oaCYTDXHLEiUFR6P
iuMDzDg34b0AogJLnLK+9LTN0sLkNU7tt9V+MHWSP0rSLCTWnkQ28m5m1uwRI3d9
8lCiVfnUNnXSyXnokFj6fmah0MckaqwludHZcZ3uSl4Fp7a546Onut9nKOBdO9Fb
+pvjghXwOCuMZvdJFpQxzcRSAVRNHi3a0ktRPeFUrauicaUni12xyjQ/gtM0TAB/
yddUgMfRJhAHSYeaiJJnqaoQpUrmFmbHtLX6CWr6+hW5dj9DxGaKzOH9n/OGHiiY
uWbxeEd6lCh04+XnASw7zSfXztJvoFbDFPVa/b0Wpkqu4TF5OG/1HFyNNWfl1hDU
u5/dSyhXjaD0r3D8y19XU3dJoga5aJQ+QHqI4zHO9a+fl6siJtjHx6sfplXAj2pg
YAr6VuHMsNM2S8zhsKVTKuXnQghyRvzadwpC+jfAECdLt6ghRp8WxN3sr4mhdQ5Q
FT43J8eJ2ZbcguekV2b0IQG9zDkhWkIAlkpTum04yUumSS41LgaHPP/YJFp8uYB2
p/J16KqqJdUQQWoYpBHTAsXzwxV2o9l6jZktsbF5boygY+ERwdBJ5PaZDNOunbch
/Dd/reWTLP2cSIdtEC5ootsItKKKi1sMb8/v1kvYJeLDQG9NHenew1gmMbtmzsXj
Mi8S9zYtgnBBIWME21BfjyLkQBnzwn+iW0gwZyNuZfCC1VaRfqWxAp5scyRXAcDq
WqYByLoI7NepYZtF8RbO8U1dfwzZ3pHgB9qH7Rb9U5keysvSblKzRw9OrMCuy89t
2t74fqIxb0BbUh1Ee6UwLAjpUDo130MmH4jcpWeTfsL7TwjpgaqFgBbHPx3jW5EV
zIce4D+QFW4LZ0N5B2PnD6pWw5EYW62tOmhfPDjm380ozpQhE+3MhZ7sMjNpdruJ
O8N3lr5zFEvLPN6/N6o8ci2o1E7NZdfd5SpSsEKkH5T6l4DACQKFl8qmSaChwW1/
CbNEB6dUE+fI+FIz5CA+9/1nkUetp9S34+DWF32XVfVO3oE88/UfwInPsDs6FSFQ
VJ0xUfmlk7F/0lTTxrwrKHW3TjTtsMN0nBVvgWIZZdCfi3wXoDvKzGsI+fkZSxei
1fR7VYJx0INREXfl1ikgDJv+Fk8EUpLAqZxmMX6Hhx03BTPfFXZCkTxgCKxoyzNC
knHuu69kkohSLEWMlOieSTPr/B1kaa1+PoWeHHkOHAjt4t4m8CXm84QWAnyFl31i
oUemrIJVw1C/C1Dgrvx7k9yZTHLDBxif+cwsM9rLL6x1bKPjyXDs6aW5dCdLxEb/
yyyG2/ZrhO94/hEATD3UHmkqmTtq9V9+/+jllDr9mL1Tnu6ADiaB0kZs50JgX5Yd
uFSFtItxD3OjnQgsT1YyPUzPoYL5HoDxcw72goon5tDUqfMJ0RGtU78J2GuSUBWh
4MWzz4o6SWlUtEVFIru3WP8rTROjFIsKCtuEk+8RaaxgJ1LI0yA5LEcKNDBw261T
OZeHNDvfalDzIHFrPr/x8Rr5PxVvlu3DsoSj7+gDfrUypDG6xHbW+8GSwzgFinbI
1Mp68qM6BrRXSCTbymXvWKhs89m3XUNkvrg5zFNNeBIhH/mb8GP7EltN8kGsDQkC
uwhIDJeDbf1y+DXKYiX5/pDJOw+doGkpENTWiND3jnYozVmLL60a0eyDq9QoTqEx
FBqIBGyI0xMPKGZzF+KXRqPjl+wn8t6397XWolQ+uihce8mGTazDepqcxyQOhRec
dCIY1yd4kElV5q0bheKUNhW6ShZafWGdqk8KDNTniERkTS56PFCzBAMZ9qznGA7L
Xrw0sixaIQh/e+cqus2YCReyS+wHoqnlMAaenJqD6HxOLJ/0hwTKhzrxckdFtePE
J3zQXYS8tK2qTGLSoQ5BJnENOSCfDBNXv06soxGnRFTVGm2lTCtjx8bW1tedqaUv
ZryRM8c297jJIido8VEPzttGSxNsdpREpuyinGYeCFNowxSEttlYUBvnYrY4xzAg
9aeCG88wE1nuKlx7jQvdrCokLAB3Q6OTPlHjSQPW6/mXgHeLB4GYfgwfa1QzeNBp
HmnOOFCVaC4tagYQpsHcccluyM+YaaZJjncLX/PmsHbFIoUaZg3tTRI5aI6pkm/6
CEIRGQ4bZOzlk6C3j/qJgurhCBZRDosBWRcSYNStj48dcMKqYVivVcAeVRBVjwfn
6e9TjrwYTTDhY5jA9mLVEZCRrlOHHvQtqiIdxIZosVPE60/0esAPO+wRXF/w6JWH
kl5qGbaXAGZdy3sKi+hm+i+gO2Eshw1zf9UPapmOboeNwpB25LOIwqABCmUPI7TN
oD/XyEBgkLF/8qmbMMsgxStgp+WkG+dTsRMsjhjLupAWWSjSlZJDG7UpJTjXgw4s
ASTIh2b9zbIrV+RuE2VCG0ibqsxyPU3HmpBeEa670guPyZIYgAxQw8JrvBgEuQGj
teHyHhMBL99KoOt7amt0cmcujWrdpYX+ZMzr2bx5hdry3kwuF4P0UHGL2e77zqGO
ctI2yRujVkHQzeyHAst7XAR+t8vPwMPL9QFXDBG47yPcDMOKhu5B/2k6clklXaxA
R3l4qF2erU8VQlKgBDMJH9Cof1qSVZT9mGvQwB0wBghjWb+kJLNuHLHgEWEUtMls
m/G37zOG0MdTm77hjqrImhi0Ps02jS0FRZdkO3GS2GzCPn6zIWcDgM/MnUQudiNW
m96XyI7NF/U3wXfNd7Nw6BAVBFPU0pFrQAZV3KRZo6Z7m/cjF1DbPQ7Qa2jc2HT3
H3iYgj8PY1DacAG5wd2YQtUpaVNbhNN4CecVhwXi31Pwspffk00w0D0pdAMvav6o
nN4sFjEYWVxR155UffM77x5FE0DFtlNEFSg3iPvYfBkOR/akyofVClmTJ0Q/NiEv
PDMAI+ZpLJ/cVtz5V65vfDrHLYp28YOkXM+VOOyQWZju1JG3r5mf4aLpxppsTAl8
vIA3V0cOWM2kupd+qA+udTso8+O4HaLgSBOCDRYYWmvy7GO97CWXbVMtpiWE1QVi
mx1pefZdZpg1X+e46sAw1Qf30Cqc4xxeN6rXz+Oq6KsLDWS+ft/txSojMLIU9Thp
pWYcrKVtIT0rthIW0zy4jQUrRZB+LGTaAubGt87dqykGEvMdt0Z5xGH0yvURuXLg
HWR7lmjgjzT0s6N/5ETafTgOhfsubpz8M+G9WypLMoXC7RqDlLXlrSRd6qx9qB7n
Y4Lq6MXRV2EqU1FE5N8LnHki1PVnfFDKUMBCRC2ayy3orU5fD+FYzP/jf7xNgtH0
n+8SGT5TpNN9jVso+IKZcdZB7AAH74LNOGMYCNvcOxymw6INqvo1CLxFKB8A/Ga3
QtvHNOioa10nN0z882gxuprw1g4ED/wyTtLL55QAsOnh8Y+T7ri2XLXGzOPs/qVq
cClN5ectT98jt4YUesyR5bLAyxCyDrhheS2fo1uBT1TkrkjciqLzX/YmghXXfJT2
U0jBTUwIoX7lIjleBZoMmk7AO6wcMUZEbZzEgnk9zjLaaTRvARpb+ylf+9iXA4LN
D7JJv1C/Ak5bJDEu/Pkvjr3FVawutpmKIzqUqxKdMKcVOWjC3IaPjQIynqDQSjUX
n1Q9nZPGm8Tdjv3OWHIHr4Is/wFgkNAX8WeuN8lEfRtfhBdIyUeUpK10IENqfFF5
IsHZ8Jm182qgsRZVi43n7QkuP8jsF5PcfKnt4UrHBSQuwRCwtsI9C0bO+IY1DjpS
VKJ2aLGmDa9A4lU5OLaaxCWGg1v194IaAZ3Of/YHEBIj1z55eNR93Yq0W7PHBBz/
bHpN0DDi8vJoDE+acaVMNmyjybhFqsYMzvsqZ7O+G1U2qFNP2RXC06GKb2vRIaLT
sas45iiZxkEeRgFmvaWEgOE90W/v1lkHrZ0SbM8eoN4WG7Qy2Rbqg8q2EkTBKCb5
TalcMQx6M/hNRSQ3Z2Yw3kyU6GraiXeuBY4hqvkoNjdzL7pGsUI7C0GWB/KsbCmM
yFVjzPO5SMPCxaecGHWKH4jsCvCCBUwXdTKcJKdkpu8xZBk7yVxx7p6bS1vzBbO7
R0enSLByNWCkPX+Zv9tqRkEga9a6iBvK1X3KLKo7/ILoKdXvmeDpHCIpgToji0t0
eep5zQ6VdJFCW1Bo30pQf6SL/WVclDCM7SJcQcnNv0Fe9/8NzgM3jLcDpZMtUvfW
/NgUjfWtBrQiBqc5oKBfi9FSoJQjMHr9hi5ggU2OHQ6t3YbjN+lj0zUS9pvEC291
AmKzD3+uQ4k1bdJUK5nr1Kk2XSjYYzVtkXtMtEXz8Jqun1O5t/jFf+5JQ1oKe0Rs
Fi5LcSJmwWy8I1wlDZfazSKTpsR8w8wK29PnhNJyuugk//KBIOff8QCMxql97YIb
GXksJrMGowRcXSOFKOGLP/CjDfNUXf2NJKnsYtoVxWvFuHSmNQJkm6IbL1rH2ri4
zBMO90ufzIaj5hu7ySeK8z2ClHQ4r05trX4Wl8iu7AwGVD59YxzFIvSKMCDxGE7u
xcPa94H3hbbrJ1dHY9OaCWiSQXEgAsFL1honkvhbw7dmik7cLmAkrSLTVIWpWCAk
/jyGt0wzIgAb8Gq8/Y7rdrz2RQYPcgC012BxOPBAVblNdZU7DL4F2m00Ij8nFpKT
Yc2XSEFBXkPYfiy9pq3Sv5nZ6r/1cjECbF1pjzs5hMu4cAE4KVAVPsqaHd/ho0iI
x4ay5ANa1gIX5UoPLTHmuHXtJPcYJmBh8bZEPemonJ6TvAIHRyOG6oEOPCE9/foP
1ezv6iTzP/9/PE9LWSZd++Xzs/8jvgcEcEDWhBxMV5WyZu3s1WGJbBU+mPxOD2Qa
Ja2Lf26alNgaYvINxVGlAfF2QJc5byxd0nbHsf3YZ7McWJq0jpd8hFz04qEib6d4
w6r/5S07QTjJ7NWX652LPvOeHJ5JmGgYKOiNsvW2To4w2olDa39WHBDWeUp3h5uf
DNG0juIePTvzftcHtLsEHeBJhb5sJpMnY2SRKVLSAeBGLb4Ey961JqFJRwuAYs7H
BJ7r/IOiJEJptLOJrNNWmPRKQbL13C190aY1fz5MLjSffBM7a3CCuFAwNb0YnY4m
szKygfE4au++HQ1N5nYBe2B8euh4u8iYiesgKCHQyzFlaJ1vrfnNE0EGTBzLEbp5
k0zhHQTNdYzMNAsVAWQ02oJsgzYkJWgu2rn+Q0FYFZMTXvmv+56HZMa6QSZARY+J
dMyDMqVPzUvqtZrQsBQDLaO/wsWm6utjg5mkYuPstheJwuhHSTZMUr3c35/us1Ti
u9KS79JidW0qHdhpYxHciWQVXCAclxLnt71vm0OYx5PIVtHbQkqiZoNO14gFleKg
FySwgHr8m+l9H0YRpHcEN6SwMTBEEfeQ2+v9FnQV/MMQCyvjdbBBKnYgmo0WgD5M
dk50ThpNz3FfrVuUiRGg2Cej5bKlyOXmXtJ71tWRTJAwlE/vLtt75G4M5WKV1lfk
Qrs3mteMeuGXmoeE1g/MxTzy3xiMeeMkJZ7/3Kt7RBqVU1Bc1LA9/mwNr1KIIcVv
Ee60WHTBfaoYQza8cgxwrZ3642xEjgRSXazV66Jq3llzrD2OGr2Jv0nHgZBqZkRT
B5NCdIetkVVWIv0B8wsYUQPuqNCrgcThwYuqYyHauWHhvmkllEzrkuSbZYmWPYrG
O1/xrooxWcHnJ4cHLzvCpwW5ZKwGjoyrv5T+vWWowF3miCNu4O0TlyDuPtoIkSwI
nKTeLDE/JmpezNNv+LwqBo2LxKNkiPpUnKOxftQSnOx3bwoVcclOBdAy9GSjywzZ
Seo49gA4dM2srQQCtJfDqT2sWvfXj9W+t1Or6OP3L+O3LDZLf0Hl2tLNRw4Ncba4
dqWkkuXF4HhvptW3oR/2es2SlpxP99Gmg5MDX8J1TUIqhIL254NSu5ERanqrg4F+
B+Kg7sn/GehP8xucpYR5gSaacOyOvhnNlDlnXx+FAS0//xexcBrwW0eX3AJ8SykC
nWYZ93MFAgNbEnlYvKt8ZtnLGd8gGF8MoFS2sDf9Cl76YNEUzOeiBQNOOLsbagp8
r3wz8xJbCV3n7cyObTtjM5WxxpLozKhW1huuczcJJBUUB7Qn/m8ajl4tkzXMll+N
0CKE9UCZyURAA8i155Pwb4AQxbYfk/czjef4DwS9xJinrYLHkZq76+ReqZHMd/Ls
yTv4dhMJKVj2Y7x27dxWFdLNbvh3/nu1C+o7HYhZsOrThwRkOiz3l+J8Z54duuoO
4GTDxqzCHNntGEO3jasv7L1O4qq1VqV1hKLM4A+erbMXVtIo1tbOIUWm5N8N9dee
quVpbRYBUlL7thuXPE8GqVSIiJ27gHkj4o+X1LqQ6Q3rnl5PQpUT7wK2G2KZ7FxZ
MDaMeSdXIb4V7sQ8XpszInWWunz6kO2A/VPLQ4jj1yI8fPO3BkP1ElatzdC0QlIU
pGo3MBgg3ZqDOtmkZ0xbJi1XmEL225DzPtodsXOqku0bd7lbvocqzmK1+AMwx2Yh
w4UOMzt8P5YrT+Oag3KHo0xpa9cBF0KmAJ0Uh9fS+EqK0pzV5I50B2iiv6IvUP4/
9ndqceCkvURFIGM4YZLtaA2BJKLzkgWuSkmtP4LedMadWKqH0FeVvviyIUagaTQJ
Z70MUrUNd8AucJFkrzRM7NNV5i0/8yFS52A5mH7WdtT9H6TwTyu17M4dlLAZj/hN
MvdxaSYTWmL6XG/puh7B3zl4IMnzxZxwCJpHF6rqSLu/hYJ70neuVESLjrfVSuOR
C99N4txe2i6qNCN5VtaL8QTAjIDDDq4Mt7kdg1Jp4zsQNjAurEtoQSR5oG50IpmX
jdmpKAMdUeQJ7pAIp4/VrYT5cBkkUBm65pTr23Wm9MS4XXdAVW1nXW86R/8skQOH
nKBa1pEYihYglUT2WV7uMgBtFJFZlIyaYaoSnSiQANOOy8ckAiTf8zJb0YoOpR3v
wwgG+EWFWatTrACI09JCt4A5wOlN4TWBuojrqt7gUIWu86xkaZPy5fzlcDIdq61z
GedAEbGUfj1vxEAesJ8XooLIl/eZfBblb6auLXbmDf/M81NmOGTtzK7EWbRtARJO
D6j60UZmVd5lzQcTqX9KlS+yx8doWCHFgOZzmOZQS8qc2skSaojSLGutqwNT3hPq
HaQTZO/eW5H6tGrOfEhhkl8OmrJc5uThJWzy9m2lcOFOcJU3v6FcOH1vj4F5Zqcc
w1BaNeRauyGK/H+IjAyfVmY8r0WHkWCl5fZUdFWfGPzs7OAYn8TqrigEj+ybtOw6
PrANE2F6Ann8gPoLIsPg8zVAHA+TZylzQq1qRKuNLxByMLgTGRT4TbpePQ/GyhLO
WZKkKLwSL9iS9488RV7zD4KLVXBickYLlStYlflSwER62o6fej54HgmmjkZw3c28
Vawx+cmcFhLZ5rUiDdXc3AFYO53gaGsZoMEGx0zXko7eQN0xV3iXvHHE8NkgV2lY
xMYlchiD8AvURY0fsR9SuCe7N/9gHePwi4ftld0H/DElEJSCA+21a+hm5Ojt03Tl
I+eiajQ740Q2ftuQIaHVwN6ZzqkLUAJgT0S8cXKw9cqRYCa2pr42LS8RTbhOPsTE
Vkb9jBIceuG6TlCRTHDOKk/oEyPBxEaYE8UPF3MXqrZFyZutxWmmmDxWagLwKyHP
gMkaCMLphHam2tG6adW9fxl8eD/7b9NTNXuOQ/rWNACRkWkgW0Y4bYj8PbUY3gRj
WMo7fES7oQn80WwzI0DZKweC1ryVJ7CMA3u8V2Nh+HFVxr4BpJDgv5n8eNThxHR3
lizojITftDAOR5BrtS0xITiqZsUxuVrIbL5PXJSljTLrNrAzjQRxuW9kmVWEtvm4
YLwcsLNxe21FVEkoRL+Lsbm25VpmFGxbtl068gP9mvc0CljXQnlIJOh0vFtFNNk2
OY75UKmFEHEl1iN7m3yp+u1wrsJiWKw8rMY8MvdHsKabvBW3NwomzyZH3dz/I5Jx
RlHz7XcQyJSwH2Sw08IjWyQIo9l5DSe05n0lCztEf3B74WVrC4qY0NSXBMrNCyGp
dUAX3RMc7yM0Wo/NMc1fqxcc4Ys3bw0Dew6rHWiQYJoXAKtGmUC4tAH8FPv1ORP6
kwiwdBxyr7ApOZVtiXaa/nrLQet9orLwxnfEgL1nq7sqVcpxJ7FUkqy7TNmW83sX
2htMGNTUcGl0I7GaTCxYZw2IVO9M2z9XgfyH59hmY3FtJw9qrbiKmUed9AQ4QWWE
WbGktXKeazslBEzvMBLTZ4TGgTVnnlHRW77iNBBRIv3mArTAKEFt54QJLhkpSl3W
RxLU7+gZR8QIXWdXBi0forMYdSaC8CQaSCuwNFtLey3Ch0teHSBBxkue0Zaek5oO
CIKJeYlcnbYlaRQ00CrWbp0B2PqLvSjL1K6n+HXGwMsda8YWz6ex57WhDkM6tEHp
Vur2LQybLjoUIu42GkbpK+npj3/YFZvg/nJsGyzLXk651TGyyKmpK/aKxCLTqZlx
M4l11CgbpuITaYk35HTCXrMQRNF//aVwSdYPd5T9AeuUKbYxkWCwHrD9n//xIAGM
MDtp3o0o3bk3WELmpcxfqL83JBKiMVZY+jRfIBGaMGqNkqtXVu80VQFZu8beg6c3
gmuTn6EZWeTauewWQnzUqaKm2crlmxCSZP6yoFKhDuewmcH0fseGKd1v4NtNzuPt
oD2bWYa3nHPQMTqWVEkXs7eOETBsD2zHEbnNzsk9GtCrv0NhQhJsqMu92zBD9Hsl
o6GshEx10RwzY1c2kFDwODm11tagOMgBoJkZJvxTIKG7KZdOCJmDQJuxEjyNa54K
++Dbg+aIxnx/IwflqJwCv7XsgL97t0qicvYuSm2Vn1YAzBu/dehQdRmSeMRrzvaP
Kxvkj/Umujh5ctHfJ/XwoeQP0IhR8B2N7TQ6dFWSUqMcEEm4TbUb4o+37n5Empsi
B+JjPPstuP+n0k44mOELU65l9qZJ7nVFtlQaIhE6hokqOQ7ZGy1665/8YlWIiysP
MBf1eka5MWXPj1A4zb+YLwXPVpU43Nz5f0QxwL+7frwWet5bH/+kLSR8vCdx8FwC
g2Vr6ZwghAuPj5iSba9zenm5xqRY/PnP66t/K827wm7kmLpG401o3mE7iIe7dbG0
6AooeyXCpyo72+56H+qNMD/Ed53rDfiXW54GETWgCxQug/PyNoGNlz5gKdEwg0rG
UnSXwrDVnfkluRbJL52f8T023saRfrCVtOfCcM2KOvaIcxHovfyFHPgxyfhOKA+D
GGQjhhf4f6elnqbO6laXzcSCZ4/SkG2VeYr8LVj+iiHT3LwbfQoxvQ4eJ+ieIbAj
zJYYp3aWti16eWgymfsB3aSuBbkL/+s80M1lHBmvzt10p8godNlm8ScFLm2XS06B
RAbjXkSRgUnbRFdln+S3Qyxa3olYUWPOP5gryCYTQwIoDYsfMiMTgovLKEpEyKDH
PVLwq8geEg1ybJvxpcqWg4yk+6f9Rbn2/5Lekunq6m7Zd9qHVzGnhN0E+BfRYZ7t
n2opSmhQEoA4wm/o/JBx1HccZDnNP+aCmLpXB7Fpbj5SB30+BkEptA6LouaDBgbH
j5MchLprqFk9tUtF5dTpVipKbK/NFMhIJnly2Ah+Wsxd+MmP3miEDxd+Ppi/DLMp
Yx7xsCPI0sqS3OBk/EBfs2fae/odwFcpzWsgiRM7z9JdLFh1Zdn9+rcYJekgs8au
abv7iq5kL1Ou6BSE8UGAR8lAbkPlB/x2hlxQ+8NXrLTxEGvSfGiKkPe1hW9QQxNh
l6vYB9mF/r+Y31Z2gRjEzIutrr2Sb4VVMG10SdXPlMG4BnOsFHcmghYOQxja7CNK
VMNz8s9vKtE+ASipTzpK/tP+Mb2TdAWJSL6ferQ/vlz8+fMsjk6kh6RlVA3ZTYL6
EBnYdQeICmqvFGTD8rBzKt13mUa1C62hse1HR+sU6XfRZbNgZWvxn+sBgid4eEUS
GGFtD96pXrTrMWIf/1URmBXzozOGNkDEsQjg2jQU1jt0Wpz67pCXnc4xdmyDaZNi
FP7ycb+9mcK8lFL1IZMwC8k0+T2wAxcb1hW7vUyZxLhN9NwKH2goiykT06lFF6P0
8kpvobV11pcYO9L2eNqSd8vIeBiG7DSMGFjJEaSZDzxPrbQ+BpW1Ubmdcp3oRqF3
nnrOOniJMsBGji4iyLWGOoLAyX2aRJ0R0cOJkUwsvOBuyPBtW6/O+Ly851lczuMb
3+AB1h+iDqGtqb2YbxwF8OdKV6eL7OBXB9fZg3sv5LvzxokTxLS/gBlSgucp7CO3
ST0l5OGPDLy5zXvLSfyNs+cMzWUhhnLI19++ks0TOhN1K0mPYQfxTCL5C9aGMR5Z
D9b+HPxg8QUK6sR+6+EEGDkqlThtY1Tyh29iDJx665CIGzyJaxcV69rsoMQiw47U
gIsE8bOis0dg8wysXMnYCdQPNblrxK9MpxAD/3/iAI/d228c5UtjpBAjXIp0pt+e
80av4C8C2iOjgchLMK6FnQV2oHb4zhtOOD1dcqEbXOnD5sxczKIUfCMwzMX85S8y
kQJUZyOcCxeeGbkgSj0u3JHlQoE4g9mOLHeOL/fxgZdsvjW68SXDu3clNjd0w0Xw
uhtERyiiKxtP7ApUgj/0hNb5CPuZ4Uv56KKN54+TBkNFbBCoZGupbc9gosGIOJ5b
X6WihirWW8DfrOGku5l00fA54xIPvEmebscsuSBZPH91B5PExCQ8NKAxseRQhnlu
x4SucH8K0kvnf8GrEVGwv6RUSlg1XZKS0UY021ynXYorZffSpJFyYABjRCT50D6I
3gbORpu1EigD3uM/ZlbsAYAVreW5qgdI7WmRRSeQviAIXcdA89CYEt8UzTAwkT6x
3H/aHupkJRWZVwgGMRn3/KIiw0N3CVts22SwiRzm+4n23tY3p0CWPzkY2/3jWeaz
RGp3A7m/rbLrXOt0r3k2uRJqIfL++ze5v4gkJjlQfIUT2dhPe6To6wBbKDK5/oGx
V2JBvvqZZ8A5jVtEtxRtvetOJ0C79daGwJdwgpPVHNNEad/2k0VEL2KG0ei6cxDF
4dD7Lx9quJvzngPoYBOe8sS07jtSPxX/NvxHwWRJkxSQ6i3vYZmsme3K+iJq41do
yqieDu7gOJD48RltaGEWH9nTreoa7xiqHKX6Zdy7rz19McsO2ToqyEztkSfVs1Qu
URpLc/Vq6IxAep+InxtE3iOOXpn7AnIm6ywNw64dujk6l52Bb/MsyuZ76qqU6KO1
Y02l7qnl4vsoj/+X2bppdjkrIq2P9MfmdPqWyO1WhowQJj5YkelLTzxtiq3LaRsp
OvSu6bgB/E/aEgewE03qlKyz4/iqBuXQ+dfCbpp48MeOoed1lHIcjuWSRO4hfPLk
wbyF2TS3OS4qvAJb/7BlSOm0Z8m5hbOXqlfDSIOeFo6wEwEbtpAv75SarvVnYnAi
oXCiilex93Ez2jLeGNWS7ViBxoO8HKT+Hmnfs4HupX1pD15QPnurMQU3JMoa+rLF
/SYU0NcBRL35HxnPMEHFWaqlMnm7tgqqgrtnldgfv/Vvw5X9Tny9AVPSARCNSbSi
aRPZXmzt4uCRADORx/8d7zxxejdPSAp2A3KA8CRpbvd/b/LvCHF5ht9pbTctbUkL
8T39bZcwAQkI0HhlzT2ry1X7Ja3CXMb4ZgD3th2S1vgWyTAxC06VVUoD6nsuHZoW
z/6+anaQtBGCtJ4hZErxRgnf3NGxn5CEbZNbLwDpC0ubVPmE0DxoDE2xCLEDOePf
D3NXMrqJIOdGQbd1rQdQ5LMgtoc1iaVxlQb2aIROhZSnIdAG2is4ipfrnIT8lA0d
Je3loeNVrgGxTc00tCiQK4e8LpEOOfrUxS2RgS/WF+QnpPiUtsO81q3ri+ORMA08
iqq6D5sFs+2vFbzcEnHqVDa5CfEARw7B6FSx7Jo1KMC01tTTO/4NUN6+hD9SVyPh
CsefwuBbaSXWpeyit7UxcS3kxp3rD+fwR1AzLGF8hnMliuKNnKpljJM8Jf80rbZf
4xeJzGduLzKjUe05/LXptKf41JnXYMSKSGq7Nd1Hm769TeKchfjsOOfXQQv722Lk
HKN2MosPh0ooW02XafxdkkArtSb09mTKfToAD2bDDRAHNm3x39oQVXfujbqLoBFB
uaZHueAJanHdGY4TIFVeXc90j4rZkpCECxgmee3jsfDMniPVNgNTiIzQHKnYV6AD
OBCx8rmsjzx+WGdNP6UBxiVEeu+/0XgtVwBgKWkofdL8+DIkvHvhfOwWhiNaMpg3
lPB2VF9cVyb0B9eb3E54KrpFNH+sgq11vNeaWL90JR+KhEng9fydZL0/XUh0ZQYX
qWZybWFS5Bd3uIkLH2aDd3NgEJgmGAUEfWaCWj7/Dr2UwjJd7vo9dEmLnefOgT3S
CoTUPzvwLOj1LaSrMBUaAVTjk5it30m/2Sv21c5apIoQU7Vw4qEOJoxZebZozCU4
HTsqobqfDIAVcfLzqpkB+T3fo2UgiWdUM6WJkTpWaoXwxO5VTNWtBEwmCiruGKpk
Bx6/JIIgvQNiDZYwTWK0dI0WO2EyJUjM6FEpiAvCP3P+B4GQoBeEYnjY443CPm3e
2MdQyLSr9bdgSQvD71sKoF2gydRYnpUNgmSimITd5ZdQytqhDmmA6kmffb3EErVY
NESuBEgPvFdY6ezUtEUMAFmwiWVGAXqfILruhq/LYhYCKicmuzP+zVFATthxoy+X
fkRq/5e4cSrKMkN9tDDwNxIp9PoTY81qDPNrx6FWerKgVMeLb+F7bKy/5zQ99z9v
ikeSEfoXeS63hvoHPuzqtLuczLHLMA6GP8toKJk/J7+4tXmAqxLmySxb6u47jJNc
bREe2OTInxnqkTW+EA4302lIMVG3N7FLcFyWfM3dnDYC4DnahSftzzUc3BEvFaiy
h34cm/NX7xBQNGiaME6H4dTLu/L66rqm0HH1bl9OgQr6Qkh4MTNhkVztkI3Zx69N
5lujRKWMtJknIRxh6qnWt6kzh7QHS5xEmj70OiMHdeuw7xM0Iir/dL720bMuQGh0
4RN5QPBclrPmY/hQ1zeNDrssJqR44IZ9z72sV0u4+hAI0AFyQB8SouAtq/Yfh5ub
VMDYw+EsCWbpWleM04mD3wWdLZs1rLCC3sLgFDOOmW/I92GaTGQ7rRz5KDhFnqdh
+ezL7vJzJOwW+1RWMI98xTrNdUPHqMxAJx4M5asNsHEVzmM6rF7Z0ndFeee46LJB
OCDHcrUNkcn281eo9fokxBicCny6giE7ErFii0y0WKvIADLSOtOD3VmpTr6Kvn0y
DOpqQB4ovY97gsFoVp5yGJS/9LHV4wZZX5XDUGU1xrJGXfh2X51fWKE/9xnSDO4Z
djuyDJEZffEEwOfpIceiRoiPhtnPwEEFfskzA3fh/jCbj9JR/LrN+iost3cW3ofQ
XLPs/z5BetZ0gohkTnThEu6kLZgMzEsdvJhrhdSY1eSmJNIdFhfZ+GqNoAwRcVkp
SLibbBQSvVwsTmH0qHfJPFAJjyAJFXVkYIlOe0ZhNu/KzlLb+mQgykbPAYxgUOBP
Bj+RovXgHM43Pljb8o0TifQVrM5bX3aV03c2puICbVJRnn1Q7ID9avPYNlxI1ns1
vzw3v59mwIiRfhBO0Pt6MqVnER35RVx0de3OF9RmIeqZySzyR9h3cOlj0rujt8ng
7O/rb2Yq1bSl2PaqpLIjDa4vXMz00jQjD2r1mRiCNIncFGlWaUFl4oyEjn+pd5Pa
hxBX0O8xKC7e3gp9DZE3Hl75B6kjVNJ2fHgbzg+DybC7H1ds9uRTJYiapu1KXxSs
q3gwgJRSgXrC4paDeJ/5ZEo16ix3Hr7i38Vmnruai4T/L9zw6Hl4Z81vJ7KLKUYA
7NB0+CZNMs/pXtsXRWV5rKfy8ildp8xSlENngFkxxz6VGk05l3WnD1xtP7crAmmO
egFTgQlUKGxP9ZbB9DBukebr7jgKaFG4oMjbr2ygaEsXU0c+YUe4X7chjjUPmO7G
DTAv83HTXybSDu1QWS4N26SlaVfELMD1C3ZcGRJzvg5022GM4y8QlDnwGqHnqEd6
l/JT+tQ6SieBGj/qZKIbbkApY3jjkNlZVexyczyOGH/48/2p86JntpgFXcpKDIyQ
uD5pfNvdELiufr0VcUaU5LNWqTe6GdxSpMKgvts0HO8QSTJwA6jVQOWd9wmqEhS6
lDhOu3VFgNItCYPM4OrtvA2v1r9obetsZceJBzha2CKXXxI6joJKPTx/Pou5xigd
zU+iyHQTW1Nvqw9FZcRptpuVakcHumke7bJxqfvcEBtzs+J21yj78Y59hUqX9DHI
dwKzk1GXfrhVjr8VLv2kJkGyAaq/LSC4iDdlAAdyNNQ1q8NDCJMUhOzML3PbxYmX
Jqj6WYrd0okNuDceHxVeMOmriBVEA36HxKh98V5RuJlrt0AHu5otF1XkeKlmLPSG
X+k+eZnsLrnPr0WFce3cC6RDkhNZqRYhPTHZ22ofIflL44EQu7v6PwZsLt9EujhV
iSGbD1LtACxUdmxuOLWmkdNzpBufHzOJ59q15fLXXILz+Yigo0BVq7n3BxOw344Q
14JybXe7ggWeMGNOTeThtOW5XxRfw+59nvID9QoNvscOEWIY/v1brAPeRzg5pp4y
f/nZ29uKQ3QkdWQH8lfztbp32HBLAPddgl80tVuW9XWUB82HNsK6ebFTOKzQn0EE
15ZAj48qp4ads3ekC0bnKej57D2Wx4R0Cmyk1czfeGTs9EuPgGyqB0KuXQ1Ne4Af
p6H4BcdRJTc2OziBqIqvKeoDdgCY+3xYI5xIT+sohxinMXG8xh/aCES00Gs6ISgm
/wquJjor0o095R9xTbq5CU7OeF5WiP5gz70B1hjEH7sXpqaLR6BcbrULMnYIvUGk
2wzt4dmevgX/f77zwKScfaXQAYQ1uHNRCFV4y/uXpkjmUlH+x6p6ICKJO0frpoUy
SBr3u8eIR4x1u3AET8cED/DqLjMZjfncSZsPWZ5lklYVGmgrFznIwUNxwcOhLDHF
UCFDnbxa7lBoRqfQYGzMK9jO/5R1eSVAqJNTfPSRfrsEMLJJjwF3JcMXLfp4B5PV
LJyH2rYs3C3WSneyh/RuaFDqZzLyLqLR1daErMOMFRtl7YVMv5NIuUXMGrdvsIol
FdRtkOjZj+oCHftBKPm9rZ08i1wpvlqMSBBpTvWioK8x6bPQc96L7zfVfADL9EfI
/AYcbM9F2Gzho8oeMqa4Y8SdToigQoIhG1/W1oFRRgYfoI1K+oI7pKK6Vx0wYdBH
XBxBGmb+8Zc7/3wwJM9HgNioUS+BcpTVtS4G6d9Fr6jAGq70L4lRXMKbPJpVPRq1
XmOD2lxiRw1QHrJJxqqacKJeu3Xm6ECMNe0DHNET7O52LvqYICuiZyXo7Ib4GBtv
82SXAbC7Sozxm25g6bI1ryHnWE4npVqygVEZOEuSo8KMHIUCUNMV5DsMn5RYDFmW
DuG4QRnM2CXsSCRx8CRhbvQgqIX+qHPW2MQvwOblW5SfOrkBNSKXOEQcQ4BZs3pD
6mCBFCKwOVLNClayWNrqaMkL4tkUohytjbSCn/Xl3Pmg6gwmoluhF5KE7ILsERF9
sthWSY/TfkNIdbpEyNzoHybz2J509PJix2Dac8vUApkHyOtaa9JZs9UO/pVMP1TX
/thw7JOj7fQLcwPCZyCmpEsV75yE23qAb1lzrtiR2HDdoaucGIYCyY4KyvjqV6iE
tOz0flQ01qwdOdx3XHzpuOL0FfT6+h9TbwxKekWfL1LCrlfmaCB5G1vHv9XpGN05
HZl+6wNOUP8Ia5ZuRqGmgf/DxuCWuVJmTDQDnDV7x8aHcwJA65OiEw69ndNq71OH
+iSuqfqafEb8Wjpc2XIrdx3gGF1rLStuk4fxZ8RmyRMNiyY5/Kk1Mc2QohO0u7ud
rvamVF8mbgTY2chs0c81BOIqlA4tj6xmR/EnZnQifP+Ba0lWID8F1Z4eG1q+6CHt
q/ADYX2yIn9jz3lL53x6kk90frIdYfLhzaYHp61BQHHkq2IdJN6TfGQ1IY5YWYMu
CQcdz/fX58pB22aiduTP+JmJjyu9dM3XpX9iZuGr1tsxyLv1YisYtJK4LWKfkPeY
NaNj7vxd+Sqn900Jk4yyXSSrdrkI7wA+Rx8B7UEspCTmNQ5H86WZYIWCVWTy62Um
NV/0TlptFf+29UDFxoYQE9Qby199nxCkozAXpA8w+U8F6bnWecjNagqdeHLvlQ0K
TsB07vgjW2eorqu2jADV220CSKXMx3IRC50Mru/idXBkvkZeBA+I+wvQedBARBNF
COBPjYeLO+kWB4OhuQB+LdSpOtu3WstZekKtGh/NTx+nzXTGosKE1aHc8lEE0gvu
5lGG4bSakeWmumaJ43CiuSa5WnmC80OnfvzJIoGiqezC4rhVnzK+zJ6oOl8FZgtI
mUkejS2sfq1wleTn8r3RfdWycYHU/2hRBP4eg5MuPMJLHKDM4GUDNWMw9tTIlncv
qESU3qm5VZjvbCFflTekRerTY7ampmrTR+Knx162rz2+ho9q9u9Z1nqKK5QdfGzb
cWjqf1mezQHyxb8fRANqTYoNlIE+9l4Ubta0rwC5ESSvayCpg96ODeaCnJwYLgwD
tFo1seP8XA+pmbGGIWt/0C1t/qHj9UmStH7znIFIh0KCqi0batvo03xnRIWP4vVk
I0LpMpVE8txhUAv7Rw7mfGw1fFlRBaTIW0Ac/Qdd53O/fB66DUvzSz7FwB0BUP+W
ZrVI7TB1mO5Yh0lSkSNapLDuQIZBVnCZGV7z6JhzPjCBqORWlLcaJxv7+F4y0Qyy
A9L4ntefGtxfe8ArV274WQb8cjNFGQeII1eDLX77+WyqkTMkpV7XH1PzOdN5ftjj
b7BJv8aEp/afJGeiUwysxG2f5Zt5TINvTmpNBQyizqTqlf/gAI1l5fEjc6JxCkZS
xPHB/lWBKGllUnguh3DoqgLW9jJSRO/hjRFYgaDOcxR9l97l7jFoawgoNKjkExSe
cbrCBgCfWexS2RnIjPL0ej27iHZiXi+rvqqMEUxr8J8i6rPbmyGnPVu7fL45vHrg
9JBw02lUemhQIXgbXx0bMiCHOITFDY0vbub1iOkHKQ/qXejhzwLJPJdM40AFatoG
OYbIvW4/6oj2NemcPkCV46Psf3w1WsbLQNNclgXKPZ7WjQ8g+MJFK4y4njjp0v9z
WajuNUVz4gmJOb2EHXS7y5Y5/9cnKhT7zj5Tj+fqLLQNms7X6P+tjM8jl92vKKsn
1va4/Vk7fQFNNVU2+NYzHdmKfCNKwKtmFj528AbAsbhkKiCmqnhAeK95xPqF9o0U
XujyF5zzqATYZBlYhM6KCOMguB8gIAneD/HErX/qlk7WQ1q2YEzBCqIqiBVucbg6
2DN7mNuCJLyHmaAD4pjGzB9eCCRsgy/bVuf8ApFIFQVAj/dFaBq33gUrAffJdiaV
xQVVqkILe84icJDlo9h/WnLd2suDqzmMJrynLi2YfeXgMD31Mo+4QXqHE/GA0xhy
z8/pU/yISiO26Gc2zSAxPC7xwuDPKjwHLXhQTp8F9qm3TpODz690/BqvSYvuYZOU
oKtJ1vP92dLqJJpdNGx98SFKjg7BYqR6Ka+F200gFXmZhMFiJK9l/+1lITcUi4me
tHDA2LroOXYSPvbdeJmaAS4MQaxu1nBmwdsTP8L4EWP7uGnn1ZbWOuAYIgkRb2EM
lELW7Th1pvQgtH/tKvV5Kqx8yVPwxL6gWD200NVxNuVA4/8pG0A0dhs+puRomHfC
OT/eM/qTlNpT8RS3D8DhEOjNMnaFuFwVFFLR1Cx1uwVnDeCDM+OINb1ci3ulkm85
QYwlSi5LDdCmh6gjvG2r1v51/DMImcra13jrMrpgNBxdA+Johmp8pTAE7dgkhi3y
gZQ3gXzzYyqxZUDXTKp5V8wTf+HVmGYGs7ON+nhLrH32Yc31s6jqaRmdBaZOuHC9
Cr74S8NnY4TYdNzmkQ3ioHz8x5tmcR8MzG1DJW8RuybiL+0QttHETJMv6Ipk14MW
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 38064 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/T97rZhQva68T7JOm4bkq25
b4BW57ADAHEm2yg/Vzsfl+TP9hfO7L54Tt/n030B3RbHVj//PaP2/0tOkykM1X8r
EC4GwIaHORukYtaNo1F9qjM/8go/MvWETRpNrIaH8lD1Ddx6xPb4e9/QOG+nLICc
0rkNyjTJDeScavgyhDQek04pzOok0QS+YL/NvSzKRzJTXnCxVF9QhSoe2Z1DmvAt
X2PEJOWQ/5+SPCJqPjXDaJFYYrvb1hP0eC724hDD6XRUt61djauSftbf1EJQr+uK
feBMGa40XRQBZ4tDFi6AdAPoLvzhSXql6W68f9Bvvrc9eRGWqsH203OAzYvnKmOV
RWdlUGmV0nI5Ag0/wFRDMoIzhmhI3m9HsoCTrf8ofedcK5BSu5JwKlKFjOKOgMgs
knUHAQ+d9ievPvPWg8bR/DIYGBSV+9nJPAjOFqkC9tOqYMHNtcrrHM79ykjWC3u1
DvFOyfxuFDPuD0ErHyL9f77hH87G+SvjZtLda3RAbyCWXznBwg6wQyf5odi+UBk8
C/Pg9zxwj5bEEy1+DGgnrz1VG6Xp9J9KB74UzOPjJ8e6LUKkPeqEDjO+T/Er8GFl
U4DvieOKSMSbFa+F4qJKrM93WV56CmBiMgxlqvxj76iHF0SXl+piSQJ3djT/y1mW
qBKtRQ7oXPE21tvk/Amle3h6kXUlmLSotd8tE0h1Jcr19O+7v+8UIhUgM4gt1UL3
7uluSNAC7Kcu8ZHpQ9Od2IZzJN/Ng63TdvqYSaSGnDwHd+Z9EtPyIT0zRdex75iH
xU4OZNLeuyYMvqwxAdw8C+6wR/F0Zt+fN0q3LStH3hrLU0QPQLLr1Ho32GeIIIPL
X7kYF01cip/lx2fsQIMrgmj8VWTt1XFQ9xeV9lv27WxyJH5e7/uGMhBfLGsQ6juM
vQJnN+qVEGxkynyMv3Evw/KGqYWwm8K4JhzWzBtVvQVzxYIb+IXS5+Rc4RrMWgFE
EXavXmO2OQVSAsjCv18tfa0ILWfuDbMErnTLbRwuNPLm3bUI2m9X1r9tnpNDOk1U
Qn0AOZ/x8vwhh3UF3xobXe8bE2sTtEbxHDoBoRg9jFg4jZkWcoNLG/0zB3GTY7Uv
WNleOTYhHkMm5Yd8zGW6qCgI0xDhqYbRuksgrIGGzHZgkVmoi0CBbKgQ1thVKChr
ADRM4Xy72hQwzsSUSZ1NCqe5IeFKAijo8/aaAP+NFHI0q5ZB03yf3Yju4Hhlrdio
6yT9JApvxrdfzNIcnaJdsWeScx3xLE8PNLQBmqhKmVIiY5yWCEK7p/i5DzBjkmTv
D1quBkTF2o0iOgPeEsy0UU07UrlP4kwdQLajksYSks5u88qEUdIvQeTrWmAT/0Pr
AoLB1l0jcNQZkDUi42rfVbZKX7h67OQvIyeLos3d0XNPEhIpjoqtEkaQUtHvTtt6
ZTwC5CooXHUZtArVu9jqlRRum4utc6tZFFQBxmfzEXfxpod78XqtiY4hW79n4O4S
t66OF/GPhRok/1I6/aYdKeXjO4m5R/PVd5Gypjv+JjPgozNSzJM0DDBsUhrWIcxx
peddOiFKunBmHLObDxDqCC19CRghLszEVU6dfnP/CEehEJSwQttwDkNCNwHf/52o
fewKEKCObyqlyq38cx4nno2cO8B2GJGnAzVV5aJ9sZwpljCEskfyaH3dUlVNhIQg
PGTSptUbniesKZUB5yR/jSzxyERft5NraENG+d0e35TePl6WR5/OI2J7ssvGLRvf
+2rclEXnNEwarCJY0VjMb/i7xM9N17z9GNjYLQpTDZfbL5kI43TE60CgxJwAIIvu
BXrIiEnNP5sDBXA2ePy0KW3loIf9P8u04iNZ3VwcBHt2db76EpXbxi9kLVSqrn7A
+uZYUSnqW7sq6UnpsWma0y+1VFN+Z+wjMlu/fmSme3psFrJjJYhLrgvJ4pqpr+no
Iv0SAPcOoevJ4WwPeZal9r7aV83aCUEYvQBeZaAxdgIwXWWZ2FpLtY/vcz1QGg6F
DhTUDY8rW51BLYj8tYxdgzR5OmPfWj62jyvYeBqEXbECp2ogzBnUGQaWCm5cz87I
rsjLUjFZ5AVCfSfyc/QZFbk+nyHM8RBMeygh4EsNvUdyh0ef9TbJCi/A2Hqu3n71
IAFyAMlVa0bt6W6knStf+UdAXpRH3oUrzma4jBWhJ1P6wNgipJLb0uheiEP/P5sf
4n2xcwu3zD43876EaS2h9q3lNcFwghpNOFTwL+vdttHUVQ7FD7YL6lhNr1y7bDD9
EyJfeDOWoj6wku7dn9zpMa1/kDTR38QU4Rke34ZKymqzzI3MIUHNhJP1SHIl0aMk
ti2s18LMqEv0kZSAcwCKAR8KAMkPwYTGoonvMSOsS/O43scN1j58avAYykeuTwPH
6E0Dy6EWT8zjUL3qvQSrlosUuB1CVNAhyiKBqNsc+dkmtLlR6/4bsxP5cdkW6QMN
so+w2ilMDOJSeBGa5BE36Y3mcXwVCdf4/RJCNdFY9535jPqWKpzc1MZU3koVbis1
63wXpdW/e7ndgX4TWLija5JnftSPS/feS0nUudDm7vkvUqIIfrpUQ1OKsKYD1TvU
Ohk9GeFqcj0eDPmc1GyZ1NTSxVTo8NOaN7QVWurcx+7PI5fVSgOZReEEjn9BdjOF
ul69FVPOTxMHtAsOApRQlCNcWCJxer54aFHnNWmMMt65GwFK8S3xPATFoSXEiFT+
IcefNPNoHOY6KvrT88mRlWkG77x0CE/Zi0FnjCAYjyI8x/2zt02t4tHgp7AmOUXj
MIzUUFa37fSbQ+1pbPr5M7Ikxum4HZwBDjFLx2BFXVhvtIc4f5q3+EbsPBQx48TO
yTV0iZcuehOILUUJ4t6iNacQml8398mK54ha8lAQgnu3zhnVkRn6/Z1eza6XLT6c
v/kfpFdehHbBqVJJQ9suFA1LCofsegwa+gwYmlX6SIQLvTH16+r8L0SnSiV8q5yb
En+n8Obuu5ZeK5zcf5cua8zo5HBrjpnrjU0nUSnrIzPgxYlJzShubk4k+t+aJxx4
sBUgG+DMWf3qWJv6Kh5MxmTkGGkp4L8nzVvdevxOJzd3rwRMltwk1Ato1bXGuy9v
CEQ2nWarSnJmZywNKl5+lMugEL3F2U6R9u+mgblg18AbEXBS4l5oeJtKVTyXAsX8
HT88Vxn1PCozKP+O8/HsXfyfdQPftYPdJGb9TJLBKQVe1StukvpwcKLIWVxv9g8i
jjRztEPjFyo7FneTOUvowU29ySXwUh3g2DsahJs3VKe4FtqXSu1rDcLBSF3mLe/3
GnFOMNp9SaB8jPOvk2NY2TmNWzDNKO/JM/Wua/i6P84ow5nHeA+CLkjKEbMyulG7
aBfe9MNEVDLF2+aaJwube+SM0qz3GZd37FyZtD1FM1hK9H/2Mln7fZd+4Fs+mktO
AmLfJKbGXyOvHtOs/ZcmsdcpnUfuFZFSNAInvO3TcZbBXTaljUoJuU+LaMM0I31H
s9w48OY1V6Bho6JLaywxs1bCjrYsxfSgpqOSKPFlVJwhzM1f6bWuxLPbAGdEvmwz
jc4Zu6U0kC/BlO6ZB6NEc+jOj6nsk6j6zU6b43+is7AO6eNdku3ostSCVIxVyJzB
1cFisLTsgIM/WvAXUf0LaIUx4m+hF+w94GBPw9qr1lxkMaszHzc1C/BC6zNjyVe0
2ChESEsbENAH97p7ToJQEZAtj2cLumyc89V6fH9UJlX7K2Mg/6Whn40MAym7PWo4
HR+OWXQnbw0UWgwtbK5WoMqZqg2BdvEASKRwnM/R3SKxoHO3BtKx4juFLK1SWSDF
iphL87KbmAWOF1ufyUd6bPy6RZQ84Q2jZYq4uueZApIce9ayhcnB9mAdTxuJebXO
pKWWqYHn7nTPfpgJ3vildJ3hUvobWdKjpp8lUoefRo8fKEIpmQm/VrjI4GzVk+zE
ula+LY3QMPnuPkK3lx66FqtM5uiMOYgd/EuipQAMtL3pvDo1ptK8fxCZL+mw2fAd
wV6Oigs6GuZyXq5WlH/1YALgFRnZm8i+tlMQgcPGHBxN0vItVNHEie3JDnBQKJaL
cdTl/geGMU84PMYGSHElcOhsX3dAdfzNjxJwpUn6cCG9j6mLl6/np5Uwhi56jxOW
j8sZY1pyIefoCteHYJF5bjOPK1K63AXy6Kf5DR3yxHQ0qz+VDX63/FD01Xeoz1oy
895V3UpmG2KeHxX8qJzsd1t2MYZMnzDwNDTBxR9/2d83Y4x7No43gz2ednEMdxxT
ZSDCkBDAGFjUXZpX5v+l2h6ROC8KdPT7kFBCajazpBjs7/TkpD+giw6SmlCb/Aot
RcN7UlC+yfSttwtVMp/29KSwQeO9DQrvbxOAW8bw3Jwv9xLhXrDpCSj+PBvwadEA
TrlTfpHix1GoBBq7+5O/9H5Gy1N3EEt8t4+SuQgWC3yF/SbIiqTPw5AqcumTMh7h
pDDjGweaiLwsUu/muaifBim7jbiMCv7cJB62CYCLt8xQOlZ0r6ZXz60J8zCIYfLC
uM4pqJmWJ8uA9Q1bkv2mGVcJnwIFeqRHkmm1FDR7nx+pPXirYsqvGwoayaUpFw6R
lqjQC05YNxwBnN/0YbvRFqF+vh/1q+mJNklx+uxO/CoY/t1vBLA3ppi5Kah2zNxO
t1xGLwDEUPbNYcA2U3HUAC4bctSDTemX0qhdJ9Tqsfg/7fD/hCYzgFIeuKIVcFOD
1ac2N8RKUla5PAUs1UN/TWu6J/3qQGDeeF3NPaMkqHaCk+YB0rxwUmFxj0z+zvro
izC6aEqcsAyrKCZ7VXbdW2PLPPrG1DjxFyd/n9YzJzUjRdJKVkZvvUS7xvodg/yA
B0RWIZ6OWGyrEXebo7w3QSoxLlQQ/COKehgJWVshy+nd8cr/jBh69pY/s0QRHzmd
rBkLgB1KilJX1+guKXj652zjOCqsLs8BybjyFoCcy8nB9vWpd3fcOujYky7N1Pbj
AFkKiSIk7QBzVCQAivcz6nfee59I5+JWT5Ly1nmi+DLs8NP+N7IlViP4MXHDhu0t
N9fSlWhLtq6xTIKj/mU8P4D3aFvaYES7Hzo1GDGPDYLxld3mlFBrHEYtL3vR6G3x
FrfBvGF+SunTaQ/TM8qr2YG/kVTtfxHfZ4ABxiyCGr8SRMdi6tT/TXn8MPClNhwN
ioNCg27OtjfdAXHci7u4+ihjLOLRdSgccsv7FxdvtWt0cr3/6nqy1NUWKTC6JjzI
hly/3SoTyTdWpCEBs38qgx1IQQrHiizxC559lzJE9w7gObLe2cRKRK+3zOlMGKBN
YgxjySdqz2yci4TTuslXLoO1YDr0+xHVH7E1phbJ19T1sPOo1Z1zu1DlImDymwlv
yZRsoiMMi8JHK9xCv8Ht0434ZpUPQNXfKsKcL72gJY7hDT3jlkJtDL1owzXT4McE
rTerukcwszJJeTA458Qv1iWv5yq9aF4fzgo/zNjz9U7tp7kcW/yTVKSToGqX1Obd
KSvUH9qaa3tmSQs/u102mc+3F7fU1NPUydgPQPbYTd3Xkvpjfk7yoq1gw8FSuM0g
o5zBnVmfaJUmX6O/i16uLJXjTZfX4NWXi6AWdikjmAAD3IWT/AkNy03+U1ZVO6CP
e/PTI4iHm96V+ZIHqu+ElapD8FMxkaPgvoSaFvcnNEHGXi6pt2/vsI/PZ/3birB7
p2AUUdL0s7xi4m0fnSpek3I92Qjde+iUnQTus7rQbHNdonbiywvKCqYrtftiw3UD
Rh60JP3hQFmdKeCniPTGtvRnIpL2p/xGW4Pr7PRirX4iCKsL6amSSi2ncimpRSCv
kL+IYzrR0wHBNzSNwJX6rMXch36biJxqcJ08bFc3n1a5PTaWOOR+D8VcOmXjQ1SX
HY2hQ8lRuyV9sULhd02phPGHa+F55IIGVTTuTd7ixmNqEINPRwIolPK9cKrjfD6c
uwSzrMi+Q1C3Wid7bHoxSUDVj9g2bHjTTkeIEGeg0ZgpBaZWtg1caKyehhZOKE4+
ljQ5Wazn0cFAz4vfMGLCLFBbqOsj0VjRoxYl4MwAR8o6yAoXoaYiFpikj8dtpWyM
G5g2c5dsqnofpmYvTJWu+/uYLSeKvJ/LUcnQo5JRV9LLL25BfOKsGckgjsGmtD0B
Kd4C78jPd7OSGRUKE/sLVAXKvejKl3U+uVqzShQi0hBXS5WPUpL6lZ/9XtHhuMSB
QJeeWQUbio6c7HS0WWtxtZRZIhBopeSUevJ4w4tGwk2misAUWjoJmRhz8Mpf3yJ6
cHW4PQuacYJa8FRF4QNqSRUKOIXSlaGzG44Jk4lp/vVMlQR38jUE4TS0yEX95FDw
eIUBLUxjCaSn0mt2v35da2gj5Bypa6c/LUuVSYfq6isuwZw447C4ps7JjP6ib6AN
GGk1MkD1knqbhXohraxoDXnQgTOVmjU8+ySvS1zAJWJqLj1yHNbvy6snxzgOWuvs
TXJD0ikoxaool5nxFNJZNsxaCpk+jyskV+raodNxO/0mqiNuKSxe+Vv/p2heWSwc
+VBXFD3rqKu0H+hLVwLH7/QWr0HCcBfRhBf1hncP3/6+qvIO2J7xzVZh2SCMbdZO
6/8pHFy5eFwAW5p7BaPX0Ojtu4+jm5wpkpo2nKEGhVbwXYJnA3o0dwki7AhyPs2S
/JcbWV3YOeRJfEPvRAeT0dziG7W+Y2gIYDVrkHKIwUyNDWp+UfbWeVy/K5QF4+sN
MoRYA/bxKDElX3EPh7rtAu0TJGO/hY680Exrs4nem7lGKBwpR8Oplj5df1QqpMqZ
a8p39swZM+KtHh4RjxEUeR/IO8ckD8IkUkudFj02F5m+oaWE6vJcSskPzkans4Kw
ZeaIumOruWB+tVU0SdK9KcjtnLQmmMDYvWhgMUwO3oqsIoTAdbb2F1UfAC7uNqPp
OWQgyyAJDSzNu11j6rZaCWG4RV6Z5GNssgTY6tSqsGOmaKTEgyi1j55YegjG8Vbo
ctbsW2lX78uyFwj4Gq8sBoCNP7urMCCfF5fnNZHxmjB92sTFcsfKwzC4Sxnx7n4k
G/plt9GEQlu63HJMeM0nLnn3KdmjS2zPfYNy5semwINLJcGH5r6MPFtOEsgcArWd
0Bc7b6zT/c6TTj5yIShVZKBsmtdfYP9DKAM3Ei0Ac6yRlz6oIfgamS8KfWsVAnl9
rrCmCXQWpA1i2dHrjDwjGEm1ov4DIcq0nzORjVmFDBcPKIhVABBJdEAUoTSLsBhR
KwmsUOvUw1Sf8Rsm/ZCg7WYnRuOU1uxvz12GkrvXjueR8207VGUdS6K0+LBapOe4
SO58+uJjDFhOKi7W4kXJKSGQJxCI/08DkW00lBY8fMyh+m0HoHwSgBvcpZzW9ArJ
evIL9aVNw7ZyUIshCXZeNT9e3+XmTkOqQgWXWdnpbRzsJgsQDPVVcGJtcg93fdV8
idJGoujJkOBoEAxx1UHVVujc3XoWQso3msa1oW+p+cYCNwSzeRFrMMAB58KtoZcH
Wb240N3hCoqBRyuHLMvDd517lPemWzI2cttkUONGwkhmCMhrO3KLo5BO7dS7/eaF
KecBAllUjcyyhgozEEOYpbhb2XN5DlbBqX6VCdJvRnYEyVkbpJj5djmOt9QFeYHz
V0KS0qN7S0rr6A/Tlg6iriivAC8Ykkg6/VUeMUziCTtChzfTVuJOkvC/+8iObmBf
+LWezsY8ndpdQP1IyMDuwF9UltY0sAzPMThvwFfhVSloFsJ0Zc07187nHmawo5Us
nPDLNse2vn3jPhtcQhXmtc4fwTz3ZUkT30KHqNxSihdliH55FH+mdcj6vUm4NWZg
KE04UIR1uzwRTZ05eSJykwIj3uDsna7o60rACAYCXhvHMusiebd258lPt5O8IEEO
kgbHgkanoalqsKoLaQaX3XzSlSsPGFAczK5pAVNc2mvqQ9G2BZIXRbIoz2g1NZNC
Swu6yCNqqTaZ8/CB7oa1ZqZWaUKDrXjfXMwJ8C5ZwT5fNFyX9M4sYUfWMDf3IuDw
lcaA7Q0pdi4njkXHnKBgqk4dsoZe0COU2Y49PoVFtEuCNiaQnybCCb4JaH/s8IVn
HJVttLUJ6inKT7qNdeAeWRalqMmEx4/6BN87cJTZsFYzrFbzY/mokG7E5mAe7B0+
GatH2DMuDCVfFwdvNzxI5UXHAzUyk5OPQUbv3CJLPGxwXDLoaxuJKzKi4NmpBLuO
fkQSb9uM9pwYOZU5hc91Siz1y3giggy8x2/2dMYMakWWv/d65g+BWd+udA+dp/Zv
l+Lb5tMOoYKb0g3zmEEqHh3S1mRtsXFU8nX+x0W3CWj4i2daeDbhpk/elAe9O5Kz
tOmwbz1HCc8aIaMjMMohZ63WJonRTqPuxJv+EZcL8iijOy6o5A7bofqzNLcdCHsM
LXT1l2tOa6BPN4FzFMr6JCcr+7K/+hqQGhxLHg7aEK5riiH9JeL9yfVrOhYGMd84
NkBHJjGB/kqEJ9O2eTI6wTfyhGRn+MPWz5vLTjnpSk1iQOfeCrPFihoxITYvndEw
8TMA+N65/atUbEDS6JNWY4DK3EJ/YQ0zL/jJjU+XmtVYhX/4iifYpnVz+jDG8Zhx
Y0Lsj+3Rwy7JfuWqSfkseU5o0HTbjWJe7evK7/dFtCFbl7FiorJU55iUsA9eRJj2
UHAF3n4LmFVjF2MFXJVHyczx8pOsgqPZXSmBUU3NHSks1I5Un5gRgXIc5yjez5Q4
uPeqS2E3Sgletrw8xQuSYmhdbl0RiuMDxVDSdNWxq8FUj8z4j4odnF7evQ7W8nbC
xdoDZ5vs/tZKNHIpHRn3yd3gOshx9v/hWWFk1/KDBBdteKvH2k0FWKuxzhPPYefz
bkFTopXdiArC/3fgtkPy2YErW9auSu6skIwHtJnBY/mR4FimuzKoHunlGFhdxenY
FDC5iF19N+nvI6raJoHD7iveaFxxKsu7qdsu1E9q6yIRVmHhFECYfIoqOp2LgXeT
1paHqVpr6asTa3Kz/bGMzzKXOGjMBnXCUlP6UBJhJgjK4FvS4hJ66RAG4QjT4kh6
2Iy+3WoKeFZW1ngCDPq3rbHfv0vzQ3LDKlHWMFu/kIGDKgiVWG9M+2QMSZ6Zh+d+
agaLym67UyueyyEvLOWzHSODY3LBqZpEFEW/G3iY5jiVEjiTNXpQYmauQk6jAqYo
ms/XRmWQiOAB/MghANnfX3XzXXgrkrKF9o3IJwoYm7pLbUTBEWVrynrE7QlpNPma
+5XZbPm0opdLSpFYsIRRdWR65VhghS/Hivc/sCSFqC+z7cCoqV7hfejxVYSgh0ZB
wt5N68+UJwEDeWF8O6QpR6LMuFvPwukW0GaLJKfIPB5I6UalSsAp2RknZjzFdJNk
k+bWlaByFt0amnHoYRMmJro+XK9uX8I3qlZW0DfJ7HEkRlBxV/O7nfKfJi8idYts
n+VLdXPMg8AkbyYAgdhmdndIM+sM4h8RYSw1VH+kLG2qWAUbivY6s7Ef7Bua+gOj
w1sw59PDZQ/DhWJkEfRjR9rFlMoWz3zPz4URV+cyDo4Q1T90ZXs8RTVwhL2FXJmO
jO9t7zDfEjSLg4Xyus3tbuawTQfIMbG97c1S9MwV8+8DgavMpNF3ZWxtFK200sqq
UEurpz93EdAhIL8jVQwOVXGOBlaXt05wCoowml5PkCiEDbw22Tur8RWInfJXIrY2
hDN+irI6pgNuxdDEFcPSEbYuJCGExcWtGJCDl/eHYqdwANWQcFLM10d+1ZhLcIg7
8qkywHw9CAXO6Kee40hTBvGmOuvaeyYfrCTWrNrcxRElLu1gulCLTKk1pP+Frknq
3u73cPAJj+Rq35BGfjtExKkjsuvpGesRPSYGPsFnbiy/kEDhTfKwxeJyNqLANoj3
k+8axwuykHk6DMfcM4G+Fd4Y86WaqlvL1KH2Ea2Sm3gMyumvQuLZys5SkHIei9wk
ELiVcNLPVE4LlZPq8GPqovNztAEChRAycliKycrRZb3sAUCOElerA6+h95BHZ4De
8wDJVtvRa5sv3OKUwh0DPSuz4BDmJy/K61zmXkbQSZFTGBzJcBheetzoQYmGJeOz
MW8Rtlgxn145EVpFX5QNBDR5yjsq1z1R14EiS2rzmwa2ULRQ5ETEQRpRx9gpK+ZZ
IX6r+jdgwKGhlNsfP0J53jiXyYVwv1CsRr8wVYPQpJ3kfTr5JKIeBTQo1rYkoba+
3qK/HQ1E2liKKoQGlBYS12E7RcD4kgC4/3BK2U1sMj+jUsKC2LVyvEZerfkRyxET
MmU7K3YPG8Aca01A6n3A/fxQkPY+hO+TQy8JnveBcIgq7EXTLn14U269l/85/UbG
kynd/kUj2pcsNS3NYsjmaQoDwBlU9F/CkbnuKc505Q3pdvGjsQNqZm3QL4x1N94+
Kuf7RbrXiTWXpAYIERGYiKMtqTObBRtuRivWk5CFOdGmSNlvvN7Ilc2+2sg6O3MF
Dqv/fe6es9szToB76WZC3FFLwvpKuGiZrAGl+ywhJ+eKwClkHlpXLiQks6aqCUpg
FhEFigQd6UrgnBJNSHwB0wZGbrj73/QYM3plnw1yprSYrrJlliLpSUWQtfPkUk5w
79p8jQ0LpeJt5Rz2FkgcI/RLpLkE3HItfTVc3m6ckvceDKZ7Y7b4rpI1B3X3Kqy4
J/lk3PMbCH/pPX8c2BIjV5DXwPTs2ytaqGU9DCajoVrhd1BTjgMk/4ac75SUyMUL
nLLtZX0PhOGTTALbEuy+pSBwqfeQ3xTEbALzWpsotTzQH21qYNwCtskdvKXENAyW
a12892fbzqP+gNBRVn2tMv7E3jtzbF8dnlKnbzaR0Gy7sQVwiTVGgFELK2ukq5u4
kU2FojvFNNpGQu0kRyFgTTQKnfdoVnWE7QrBfY19tjkK2Qxv42l57bbx679AwANJ
CnGAxGG+Ks05ARrBtHaAt58vq6xWCYnZppazErbmpS9+N6RDvy7+5LvznpBBFCRW
uLsH8ySjnR37KdOA6rJrW8cZczgIUgvcFtkpz2PT9MvIvEZzGHpz6BxQTkiglEez
CXVZMEC5H7QvdepRG0h2ZR9XEwbg7EKrvejJXj66gbT/dQVStPVSNpWerZ/42gWt
rilR0V6VU6Cdy5UqW1ppTPeTsNgQY1vCUjtmiAysLayisIrq/9w2ctNAVZrzNZdI
xe28cmtEaPGvSTbhGjJQOzqF0j699ETafgdhg/Sv3Q26QpGeAF7mK7IZdsssQCzk
rFaWcj4GJ1TEImmFqcPtHxsWcph0xTBNMjxHplOPptk7bc3buAv0GuYvM0qrlWX0
WPFyzHWlJr4ly2H+fHOkAIRAYUEhiEHUUmoQpOa1PzI846sjygTZEZc50E32YtqY
dY8olGIR3q6JQDMRawZuyR8EK63iQWL3SfVen1/HycEE1H64F/CBX8nbab74FXTE
E+Pwgl7NRCxKc6Mr+ye7SXUSseIivojFe0f3EyXijXfScbdRpvgwP4DqvyN0b64A
b/6Ro3pOvfvIqKe/W2an6WBDR6tJwrfTcyGkwZIxp4iLmDkY4UnNYcG/WdPdgvnI
/MXr3HB8OYSsijOOn1DZW9vhCsInx3xoJanRJQqL2b1lQx/i2Kq6nfYezy6gOUZG
1d07j+uPoJfX14UphKsNgUwKeFkAX9Bh/HfbMEQL0t/0rcpySzHqQ5/eUma3QXfX
pxE+w3ZAkzqCu8pEJvilXq75L72A2OJrzwvvR46aY9JXbIO8qZQJITphbZvbuN8d
w3kf+nGEIxK8mFyj8f1qmRUSZH8iZ6CPyinzVbjQcADD7P0JlyulwYyCThWyYPD0
f0wynyUX3vrPgEK1GSUwog7hvnytWmFVRDn/qtF5EJYQAP+qMuf2Blh6udAy8gC2
mXXHzAeK4VL4zWv5m92RWZ//meENFHvSvJ1Xd9d+uw/QJYjBUS1bkHqAlY5snAbB
+STrk9yRZ7vHFVGFYfLWZ/zyhh1lMelyax4S0FjC3zGUAV7GSZbPj/wTwu7rJLvG
Fkcp1g4rORfFv8vGQaSC/QU4dKAiwRE/60EGWG7VSAR0MLF3nlDAOehwHGyW9cvv
PW6ipP3+LIeGJi04ky4GTNoRSCDfAoegTqHkJxi8MVdRpewsxkLgNREbxDRE22fc
L+A60TKjV1ytnp3CpV9BCXGc5GCE/3P3RSjLu6TcT048LyfEu+zRpr6gmQi8Xg7R
8LWqQy7EnOJNDItwZ7MWdaVgkbnLQoqnwYV6cahHYVsoBVYyVBzvn9Quwp5sUZYh
qwI1+vFpp0lnCs+tREvEOIl4RuIREfKITvI9mmM4FTWmVJnMVSp92iDYyufP5dXI
H90hfCDNXX2ZKVLpZlQa5cNXwpj03e6JxY/WELvKTVZ04IEyZmXsw8pYtlWUoEXE
yG+y0XAEWYkY8aSDSgqmZVDkQOa8dOEgTD/1Og51G0C3ua/6E82TcLX/1gDEFQ3V
SPlCHwcyPIG5r8dS0jklF8HJcFYFJSb+fiq8CRJhC8hCP6DFBjBLF7U+UL7gWMsI
YeJUtop2NIf9ng/lbyWFcjNqpMM+K2quNQVJEVHOAVvn+xNRw5pWkMwDG8dLsErF
gOsB5r6NvgXQlUjALEkjcDfnQWvd4SgaPH9WaABLIIsKf0DAp69Kd8LUqY9mAc5t
kFlNt/x5M3uzsRmYrxagnQ6OOR2VQtUzAsQYHaKeBJYLSaoJcoaKTZ2Wa1xQeQoB
BpDdKMSNMG2fNi5uFKz+LTRQWn80LzRhJ1dmPOTA9uKwZs0BTW50Myw0/Pe28FmQ
xVvMO5KiVV81zj6ymnzCcFUz9OvMxyuqnaOoFByFOvnyvjc4QXENTcqrNB0jWRqI
eI6X44P5GeIkeqxSOcQWuuVXkkNDnLQt8Tu5RZAHRl8fgma+2nGLKnAMRwahjCKk
VCkadpB1aaRjXrAguTcvAPpOp+Bb/qaD5b60Co9BimgM6rpjEdA0UrLKfdgFz3eb
iHO9fU3cRBULzNt5PqjU6MlvH69Sdp9IWK1Qg8dt6KOCjETS6K+epLDtEmuw/XE1
oLZwxITrroD/P2a7HqspCEkem6zm0ARjIXQIgkfV1utbPXmZcSuJBRZXtQ9YrIZO
GLYahzT1xLhdnFitAHfj18YWghzJQDPvdsZTDtLYDEwtVfNALqF4Oqh+Ike0yA+W
F4fatb+diH7+mpyItPN7OlAsPboVKI3aH3NR+uMMMdjxA8ldum17Jbb+SFh2rRJA
7yGbOMjEDeMGxd4LjsP1E8AMeCsozAyfK2MMWt2rgCgCKM4IoNfNgjXZgvo1fcfC
yauetEr73l4cduDPhrEs8Oy8kMYkaKIBG/ATPeXMVhl7osaaPHTe8Dz9WnTo8NQx
OsDy4yN1i123ApKBYyP62zBWNwbxwH5J9tixAnjoq3qthMq5OuNtiROVV+WC3xiG
bfTlc3qXPcWUH+e/JvZZYWMwf6JuQ3aRS/w40+6dDAIPHPJmckjl48Lm14HD2Men
A4VkcOOerpPTQ88r7cvl8pN2URghcyofYoS5zj3irvgwXI3LCYa7pNoUJ3/O67xg
kqvt/ImFTwrwoEThgUDqfEbNS4v4Osc03MCRJhO/N4aSvJ+m4yBoR8TAtkJX5Mdr
S6RA6pM0LHAr+7VCaupIDxkUzQognbJrLj7hlrjtIqOMph6+g3Yx+pS7t73GrDZu
MSZgUtE2nAxqn3/XJYSEi4K+PbDPfzEh3poyM0QTGHcdQLXAtNAwAdHBX2+qpxkc
bHVpI43f1fUKyq4BwN6EbnzAqboM5hQ91zNlGnBAy+1zcnhK3MzUN23dyI8/4jGw
ITIVUWjLarvfZk9Uoq+m7stjvlssMum6QhNeS5qf7412dnBtJeas/TQUiK/9lCib
3P2R1cpqBXvaSKTMdZQVCeFCZaYHTKsLCd1o07Ox00uheBbLEzPUSm4VF8eN5Psz
dwiakTvlFpm6Ay/dSLxP91OURfeVNm0OXEKru3OvaQnmA86Uw5EbtKb6wBm7P8T5
ipeHAnGGPWCeZbq4K4IFF4y0C9AcEW/mKZ9ulLya7T/9Z02/rIVlSTuKMDmjgNct
uWD7jBgQK62EjZDy2rgcR2EyD3Dat9OlRPQL0cy0Ng0F5rKnXEzqMqoDVwSB/br6
Neazm4FU6Ul5dEpQScEKCueq9gfppHBGbLB1hNJIZx1LjDLRsLEe/pSlip8FAFbl
WaWHRcxdj/W9Nnrz+nr6gAnVh1bk0p/xR1aKYbT1afVzfiVyNKE8uy3cXgJbWXU5
dGUKXSHXUH06zPV0IvM1o9N8nzXutiaIzRjCZFwi+s/W28ETd17aD40VF7Mb7zMM
p9CuYrP0I9XpWsDQEINtbvtT3koidyWDbydo9tlU4u/AXEDsGF+gSjJF80+ZUEew
5z1/FXY/I9xt1mqSBplhKSx6BxJJi/IL/89FGcYLpxtDKWNpxxjNJ9pQmRPknq7k
naFCqmNS5cxMX2MFuhIpz6hy50KZDIzD3aUYQw0FyHw4P1AkE2gvQjEISgQ2n6cS
WHmydLb5GaNkgtu2dvYEH93deml3RZ4DMiHG34AQLboKoIHEqvasjleKW3RoAJkO
Ky4srmzozONLg9BLDsu3hwyLui63kLsb0yr8KzUpX/MxCDtrv5yBDTX1TwMCzGuV
y3O27CRdN4MMLbs8qFM7J4zzpqmKrkLSQFyW99xzXmygNRVP8SVNxBbTDjRLf8pA
UvZiUEDz0HK+XSTrh2Bir39t1n6ciIxU8qVswYiv3joTvTZCs3DYMNT/IMMHRDZS
p06WrtNHWdYJ4+9xTqMnMir4eGtL8BYjvihtUZr2ifaa6sdUbpqCAPTJnRapMaEa
lRHA+gJCGnIIidSM119HZAKrkEQdyNxcwnIHv2zmKpmrdxl5b+fCN+vnmZ1fH3sh
d6tr23aRiX2cGRsKfrFhbMP6gjB8z7hs8kMU288fx11zpsE0hTyiH+X/m/s73id1
+awmzMvxGaC7t1js3lt+NmqlNKgQqDzHWg400KahG9iqkqclHCWKtrVrsQaymjrS
r7tvfjaXm+PzrXBMj8ctn5zcGU1mRs4qhKUKoLzYnF/e1aW04T4nsrJOrHjffLe+
Cjvdbc2KVI3J5G3zfyYFHNc29OZfX0oaLSONi93RPg9Il4qHSwwnUMBrvg7y7XvI
mD0ndCzWj3Qb0GJmYx569kxFkEw2zv0eCDr5njlVBSGe2w7uYGqScmai29GEf7j9
9YS89QitGzYRfqGkm1m3GCeFU00H6oddNPCP9u0m4cHd/TGV+zg1yUV9YOvE6SaY
P2ObV/656Y+yxBpaQ1mOYc7d8Vy8AY2MCpZUaXfOlWFTFQFmmPq9torKA5m2ylfC
scrpUgyW0IupUmxV0wMM0eA/MpwyrqpnKhmGyjl2UQKQhy1dwxxt1Mt2HlfK6xgB
zAsgap1ERHGP7Hv/Enzrd173DP4Bn5/TtOm5xCjBA7Z/QWnTh8DOuOOnFkCxdHv3
7FLrkN+PFnJcfukSgOUdw1iyD7FYJhzi6ZM3KBzmmKHRg2yf9Q/t7x4gpeVALDpR
zAAOgR4cpAnQQnShXAVmu0F3FwTR8MpuC+Y2oi9vFk/0qUsyB+pZGwWP5mUu/4el
o5YQ0364QxrqqMRGOxbRE7YF7ynbnG+q8Afc6lD0YGmTPTnq2H9EQer1ylESEt82
YuMxqUWkHvbzeqhiWQY+slzNqMntU1PpBcCDTczooEFCUUhuuX5C5pPRQE3NNwkz
lXovAPX3ncTOF8pCluTMiMqb5/1Qxek7BMpLKoo7dkfecThTU8FoqAli0c6oVO/L
k9N/UbAV2gJ5FhMBoCNzTvFOkvDsj9c1yQ+GHoE9Z5bMur4EsUMZWAggRI14BYhm
nL3O9CzmhTQpqPe/59jN9WXkw1iclsZd2x7aUnXHz6fe/owZ7J6TytJmwgPTJJwy
EbUHG/J6LhGxVyM8ywiyjG2atXwJJZBpCCu5qvdTSY+2q1rrPouAF0hJL6gYItcX
QRJhRncTzSCUilwStecEG6Lz5Y0FG0cKvbRJkK18FW4LBVGCl+W/X2OtXGitsb1B
xFnB46bOwHYsEstO9/I3Db3mtlBYA5CtYbM8/aVmjv0MDj8jVeZ1y/K9nP3XzVIw
JKXl50bmUinlWGNNbcQci9qzAAOQth+4pvihToxx1EmclXuXqKflxgFW5AvG/QZf
Ru5JzYTxPjJqYeloVIcj39MUSNJZDUdsMWpA9+wuRoSK2GlLkvGPtWds4GLj5ATx
XLM+NEKQjOvxIXgb/ZFYz9cmQLTDnWKtjU30bX/UQkROseHLD10dZ4Mr6H/j2duc
5ON6DvKNmtRf6uR/9wBiF5AMSGIzc/0IT/mk7RqgOENf0+BUHzMkkGDMVTf7xss5
dkUSJAV69xaGsiekeGtCFA5uYOHL+JJ2roXCrNc5UUOZfcZZKpZXshZxmn0utFI4
VuT5KEIB+iP8Si0CUXHEw9pmy2FlG66KXFWaQpBSBHrr9boMzye9Bt2PxklxjJtO
oWxwRpkarD93NP6HTIBL5nV6oMjkh1uWxml05AcIh1QOSuVjwKVCC/ZzqpRiRoUK
AaSEMoCMeXtgvQtZ+ZIj+hQ7czkjFY5jML/yCbRGpYZtBN/Oy6+gD/bLf/GWQGPz
Vem/c74Izzyd8gwIiKPCfPX8k3uBQxRqQ7kI8v5KsYKolP/eVDYgl88gZwJQWV+k
mxli6BXyBOBVsw8RsW61b3EZBLI39WnDIf33aSqqoh6ve0RaLlrLcbnZN3raFC3S
HJebFsxePnJJlqQ3/yQ4T9kNB/9c0ku721CUhEZa6aX7Kt/FuAlaNvYRVuYNW0n7
LjPVX24mMAi0NKoc+vLtVcRpuacYvuN+Y/vHXPSNyzDnEFObRhAQD6nk7PYNlDvO
jW5qXKTiZas8qjFYFsnG3q7Xu7DcRzoPM8XDof3ub+uAAp9fWSCoUgOYLJc+l5v8
JjiIOCVHSNwRVFf7KGhTtbbAkP4JErMQEiSrocKx49yDwGLiJ4G1U0X7Ln8Ipzi8
HuL5SCjjnKwhRd356ZhzJx6pEeJAp+mX8sV0DkI7Epq72s7YVK6jqLCOTehwI9SK
i+2IagAPE3eDS60HwSv+EEy2XpEG0gM80XQHXlegJDJn23CUIrgRgrGQZscZUo9e
IexnN9i2K6XEFXwHVzSt0Vn5NHhfRslwaWUuUxh0g5TGqRHymxcfplKd0AdTYBx4
rrpibP6tJ7kG0twcxjKeGYXoTHtuZO1/Yjstg2PaYc73NY6BMVJqmJzFBJVuOAOQ
KmaHsRc4N+Y0iB/VvMEDIGliYNDOwCYIipV+9lJeOvabWWwEYiLLAnY0+cl+JJbY
khK4nuwumv2FyxnmgsYuh6lKFqmV4tHRPeX7tH6ME6Boy2mFJ/FJSekXp33Chxjf
9UCd1Y9kWLXs1hv2IWliK0XU71V+5tjd8RVhWKSEQGOlpzAeSzs/yKAC1qUMEMbb
phQ0j6j9G2EiPS4xARr1TdxA/L/bpu+EbIiiLrwVYMtfFqhyVt0TZb6Bx0sv3gJV
LYQ//K0PWYD6B1sBV4deJO4IO0NaTOdtyHuPk7UMxX0p8b4MdG/Fe5wuUw7rxZ7a
P0lxDDA2hPLmFFNfEj7qLHhfXUD8TCSyIhUlxWglfpiXpWxkVyL/4Jc5OKk2rKex
x9bKpuOWGAhRvwks9hXGZZ2q/r17EhLpm32I0Wm9Oc75IqCoXR7lGCechZAmxCY8
2kGe64pTf+IKEAE1yPqxySqoFwLz8sP8PF69oN3mK08ecjloQ2zKUXYCTIyu8mYc
G5PoDDjiaZUFIxd9buOoBzz2AM8vfLvswJpvImuac1KkiCSLMSmy4H1ztgVGtqOB
J0iKCMcEneaJEpORrnYeL8cePf50xao4m1MNvdZxDvrTajpq3pjDRPJJ990jCH5v
Pqdm17wAG5pveu0/pHmjZlsPbhLDnoeZ6bzZe0bZk4y0749XFUcH7k8P9hNCzWei
xbS/FxIdQOPxAIB9GfSF22Wjo4HaPkSsPsZG6mq9KBo6cC0a5rAghPI9kQTtxo/M
tgPwMRXsfor/YkjrIDa9p+QJiDkQLhdlJxK8XvB3GJ9IPPx9hr0LttbaB1+p/100
gzwwUMI+NGiJdwhTjT9WY8ipGWdC3P4FeoIPAxu5jn3XX89DOrGK9OtvfKoVceqR
NWmGGRYehon5nVM3vFC+whQrrYz8Hc2GYkE6v9YOF7QcKBhG5VLaNd3VcocycIdU
bW8JGYYELpGkldBvZkAgi5aw1ba7G37ItgZeJ4aR6obt3DsV03uqEEAMzzB8o661
e2AYwwsjcCko8JzQIGfk9cWSHk38IDcQNAhouuFiiVVgG6jvVKmVJLO4OYK+NZ0I
JT8fUpJOXdu0u5r1o5OEZL3ZhSSh+bfkRBTYDQBaWTEEKkUudi3N60Qf/poo0mYY
RYXQwZUrqQQnfmViDmsbtmVOpWm5F9QDbocGRqSjotTUpFZc/dAVh7Q7IsNwLVV0
g3smQi6GRT/P5GVYH20seqNDvfIlcLjB9s1rCLe8n3FxxpdYLqJOkc1kJzWg5+PH
1oMWtVtkb5uNi47+eKQVCfRAiHW505J0rpDpKb1vANrctmf+K+nlvAFkOAfxq5Dn
9KZKnCjXHHTtzfOgPUo7auDBFXwOIcg65O7SfBffOLmc5q146xBPeq8+68RwRuBM
VXkBqorMhfaGIaRP4FZZdAQZ5wIAkcO0Ri1Jb3NrfYi+E0oC6Ts9EjXflh8tZSGF
ojzCN2Fwucy90/Jg/A8xjGm7NorlSGCaX8swU5KUrKJJJqbrcgZDRp/n4WEhcDKl
3iuECDKXjVv+nYtTwmA1r6A+Aq15lz/1JhL0VlN4oGkSmN92lQTGj7vHtgnT0rMj
ul+hMGUH1STLwwNHrjbrErLAVjDM6grJ50HHTyvozjnlUjs4X3e4YC/smdOpOnyu
poDDDgCJxjadfLzLMKJhV1W+uved/UM2c//umDRnvPR91XN+Ah6Ufa4jTtMxCV24
bY6LIjrL6MdfxTUfGnX+i+5oHlZvdsypLfX0CTEwg7wlGvxOgmtzWXT3cFlLmFtP
F6PL7upVj+s5JMF58uyLJvWm5SpS3HXV3EZAnaO+mQgxA6+gsjAYGZxKhek0IE4O
JDG4ICqDP5SLeXeO1Mcmlg7qNamU6Z6Rxlzhr/mCyxYUOy/VkM0/oC/0EKI9nFba
L4USLh///jgjksZBns8GsnWc70fVCECoAVkmOump2Pu3aKgdSaD2e30QENp0r0WH
5JpBUuIzjHzu7E3ru6TN2W9CNMiQjWfFGnMXywJrbJ3KCvDFFEDGpKKEsDdE+ExM
sCPPwxZWJKkMHHr8U0CSb7t1Lm38G8/S+9IS0PBr7bU+Xviveh4mu8R6Wbg3mGSr
RKAUCkArziNR8xKzeVU8Hnrs1pNuu+5qctWkVyFKA5D1T3QB8U1NWwxuWyXgnR4q
7UI7lgF2lyXmpxdw80ietj7AQamrHBphemRc02yO7NTOczR5BrX11EdtCOE7NOYW
AxHK3VOMO+YLwORRNF2MszjduRMyMtrxHCFeTYAe/gBvwOiRXCvuGHoqjZ8zozw3
AcM85uLUitIoMtVcvAHcv4Vv7dWcJWPyIvX0wKaZZxVvQ2s58vPoFaGOz/zthdi8
dERhJdLVN+HPmqtYsyu+KIwdkEuYXo3ha/5HXnBerIrWB4v3EGDOQtoDaFD81qch
rWFD1TWuOSV8/1/nKY6ByC33yZxMg0t+dkD77Dor4R4Y5oRFBpvZY9DmRDpBjk8z
2acOgDJuwpQYBtTYfM8h5SSPMtF1NLYoZsWxAgdImdtPDvvMWrTpexFrWpwQHmbO
MuwzsFTCkb+IEo95IUR2S2rV3VqU6aJHcJzc0fEAFNE9EQxLvqxh3HpgkOlyajVY
8M0rzE7jTAcR3fHa3zR1eJZROu7t7s3gXiqSPB9/wcyjf3eWk79hY32snaQyC3jz
ASKxJSWr/utliX5hk2bBQ1buKJiMTtR2rtAioBKNS6SjVRdheSoFTR6A4g3gs42S
ePyINsAjB9cb3x9hDrtcgo9KB2/TNbxpgoW1QC4cL/pKKuWmMcFFF/u97cWUQIZc
NsW2n+3bgckESQTZToXCeCc68vk2H+lEcoOsaue9/cfux0w36Ds/iSFQwJycIq3K
jR+rQUCajd6zwqNCsjjuqxt+AYOC7B4/Re5p1fHEC6c3Ow66W/84FzZ06ZjGuoYA
CFcIGZMoSWAQxzoA4t+q8dqbgJw4hh4qDU59xdp0oSnUXZ2b29kLHS83MDmxdt/K
d6ntaL96HPesRez3zrCcW9MmVLfMNoy9AiDkeHL6sVkEpn9RrZ6cfPG8i/Eg457V
Lh2ZmuBQ6P7UUiPP+aS8cs83LOCA4JVkekTOfp9ElB6BnHqGB9uqalKVtiLCqCi3
RvqT1JgrTXVmtJ2gXNYCi5OadvD7rPtJ0fd3KAXlDXmx9Y+BFu72YOp/BevTkZ5h
+zH82zQdRf0LLPfMx9/D9qOYGQAnNJPujk8rQEmQGPBccPx4hgOrmI01oFgBD3lO
iWZwOusEewApxt4NYQ3fNZbxTnYZHkHpOidzs9YDTVHTvDpt2oKw9qzlAX+2ZIG6
C0HbU6Mt2+YyKKWgPWEJ1czSyPciHLWhhfb6kefursmLrDuoQ0RAAD/NDaf3BwG0
/J3pRLeZmL0Ap2D97/QVhZzcdivKFq7p+cwhKwFbqoLeruj2IT2y7MqdkKNcf8l9
6RYkw1ie51ONjM9FyugxEQiIuanwDeoum6oDfb1xrEoVXhZvEOeoBhIWLNFDEUuy
v6WQvi/5slvGrm+wzpFufcHINjxomkxuuWYy5JqdTla2BNwcescpjXE2h0r87ak3
RPPKeJZzE08WqTIG043kfWpKUB2a5DNGj6cFUpgyQk6gPh8IEQ5i9DoXqNzMwsrY
sNIjTSv4szEfGof5ZvZtnnLv9clDFbR84htEufTpcBa0FC8bx6hDzo/7QNlU4Glp
FyypXUaEzyIDAQh/XNeZ0Q4sJ4j89EaFYGlbKGj7rTqqpWy//+9X1NrqMoS6ryix
kRU1QdRhZMnKbc/8QpQwFutuqOq8MQ/ptt+DjHH8tot3LRoslNHGLRV1m0cWnQsF
ygUfMSbRHaxWpuEq5JX1tML9vlSfBl3zYLc8vwkC8HDBmbIFQDIQlokAeRJeif09
T9K9C71Wza0ALHQKrnVqDe9Qmd264aveVghn7H4NOiS1D9XIE5JiymuNu31+43WP
+lt+Q71RDaChu6q06D7kObmVqgAWuIrP2ZLXtDSG2Sf4Ck/lfpkyY4BdBYii2mHJ
blxWgLYMp16w3YwycE4oEYfTWj9abLQl+gzewyxTt6esk43nOkFIEgDc081UMtH8
rQqi3rPog+YPQDIYyLjrvXBx4+/ZSoV/Kec306eTKdvsqwzzCtFzmeIh77t1mCz4
ix+fjZG6S7qQvmh1xaX4buNQmOhvtOy+ug48LdSaHyrL83GGfsuPRgZtEfFcI/2M
N6uUWuZCRX2CcSX+AEjm5X5FIlY6R99Fe+McS0ECXZGJ/+ICJ+e7y32MlY5VabW4
G8ZOJDwfUj15nh0agqA/X1oXJ7GvZbGe4ZxBy+EhKGhGSBZF79Q/RPGYjNRB/9RJ
vYvx/vBs6lYKuLhTWaH/HeXnftVy9/+FJ3gST+QQ8ZAlFC3eY2oQ7yS8KHsrYVN/
eQjmYvCIdFOxEHp+lXcg7sjDOd9pDDEqGzgPnqKanW/EvfiYuShXZFXOIcWR0Nqc
XDj18usNzNXnQJlDhRZzJCSavUHsKUtd7GkhPKoOXsnWox0Sjhk87CNYwdMHuHqG
Ngc3L4za+4ceGwBsZxYtz2MyveBRRc1Tb72hjptiPmErr49ZVzOPb2eFhyVC+VpD
nGvLDE0y/258iEhT7AMdctEHjIQv7tYCaKX9AlvFaaLh9iI2NJG/svM3h9+03uqC
6bwrSoXNxEFmXB7ZDMObtul2iXtnVQV916GxKKhOGrALtQNSQO4rQ0ITZfR9UuIP
35elY80f+UNHY7c/tGgP9tMJDcCgSKpj7NiYDvFbThRTSxLpsCn3tuGW2VmYDKgU
P9RVS55LyAffPPgl2shMPSXOL8aOlN3BT5e31g48R9LdDGJYyNB+3t5jOgxUJ6RC
5hWkXR6olyBX+o6bgnkulTtilykb6yTJyZ+Rg9/eCyqY8DYuSqqQMtDn/crnLB+j
wmM1Mrh20wZQCg45cROa7MFzMEeoOU5JAM92dBBcLBIkCPkZnC4Vq81BOrXJPN6I
TbSmG3R/gF/TlcWXY15OJYT4scuy8Ul0E4eb3IdBjjAXmvJItFn2iCXTNcRjDpBJ
3Pbindp2xXbbajHahdIKI47yjMImzmoT09m7pWMj5Xs/GWPpZfhWN6XATek4u3v7
i2viW/QgmbxOEsoskuudZ9zc5OQpJFJ3DdHqjMUjqlnaz5aI2eEsDe/dqmJ25tqq
b6+vxkc3braD7EtY8t2spG6CTR5SETzoX1Ytc51gJqRzAAwYbzDY0Rt7vQ28Zp1+
U4SomMFYBDAzycag11aDqt3Vw++7YMm31WejNiDXVuI+CeY4tIJdf7YcuutkywYg
nDvnfWaFsjTA8CYJ+BU3rrEIrb/4pVoQNO1KwnNhFNBxSY9fbU1bwDD9o7HqIFqd
3dAe1h+E60Y7IcVNnlXrU9iaa2u9AJ8bFksY4uOPYig58aeJJJEwHpVM6ax7zykd
VWozvy7oRjvZ/GOahXEOkksfx0JDQAwRmBtWF6zvICgHnuhAPeRDEsKjf1kq+vOm
0u1446/dL155a2xZaBHfPQqTj7tcUyz5YckNGoYK9a2FBumwyykhx+po2KPL6aNQ
s6sU4v40PfeaBdbB043AztLP5iVGCqEHjJIUlyj0mlOsY++s9zKH6yYuYPfOelA/
1tb1nv+zZXSoPYwRm+e/CKmjIBZFt0XKPQhmnY1I0lP1A57J7x1c3TZCNCCszj93
iFcPvrUJcnkmZcXKnvKIHozfFUciPG5vabNtcQp11vBg8s1m+VltoLGAkQ9EDjjE
yszs55mD7QALTUFnZ1nx/Qhuy8IdxNN1xaZPdTGwtbDO1wacQjhKZJEzWF/8uB3F
wRKFjVuoeN/mbJ4YKvo7P4kaLNFAlTTDXRlpgSjrqTIEYn9Ppw2nEJ6rX73ic45K
aJofxvB23d+F4b7b4Ek8Y15cYsOGSBFOrS3K0e1F6ZkfRQ7Gt+ErS34ps1gu1aOR
gwSkmyOx2ohVwjzl1/ypsJapAYlPLoDzVJKen9XS3y753Sf3iRvwvHrqxBo6m5Dj
z1ytPhD/VWZLNTYLSblXSQGY6RVfrVCDcf/pVzz88+nRpeMrVWgBIjfenIEyrij6
mUVfLlrC9TsBc7UhoDLpnVfUgyl8j5X62hg+UEgMIDyBpjjCK8chKYRMDBE+ILen
F7u966Yt9ws0f+/Iw4ETnSXEPrIuPGrtgvSoTmUgy3efd7EljhaXLI+aHn8qRd7I
d//zvwOYux3lelZ4xF5ELr7nkZyxBcuChRb1EhPlfpiRpH1R4PQ28JpyRFclj1W2
hrY84+OE6M6iclUKjnU8X97pCradZj98l0jOI43T/buQRb/k81sb330fJ00+ItPX
s6EA2uEUbK+wIamV3DGe/ocEg89jDrrXyY6mnwGg/7rCqHowcp+bu6BtJv0xCsqY
ntQaETLFLJAAeSPj+jasnAaLmr/W+ZHMNXlMITuByu1VqOlC55L6jXwOuULgrtsS
GZod+6koiBjLuDpmCU14AQkOQQk0mm3aRhjst50ux5YKUzLF+QCbjUqtDx2UwXFb
oQP3aw3wO2210GwGkb/v4RRWs754ykpRLdMl80cshrvXnyzwIIBqNSuHuc0YdvW+
Po0tvdYIV0iy8DwJyJCU45V6IqI83LOAKgj8qhuYKUVUmXER2jFPc3w88+6CNuCA
8QSmM8UCXo3VIZJZZCdcEgfWbIEQkfCZlX1/9tXx5BW8MDtOgBz+DnvXaPpX5md6
SY+2KlUm/el7vzMJ/8bhFT8Qfes6NgNeqs36v5Vto6xJvTQ4tPDmm2RcopGDJsQ7
DvBm1IaSpBsf3Hwh00+o8bUkS4v1YeCWR1JjnopowvHc/OcOlaCvQwhyeS5oLMZf
J2tjIyeyYsiDIUJy90fBS7XFz/Rl1lKTFEwnmyWnoG+exP4cDkufL0pUTes2Gy+F
bWSIUOFzfVa6wgUyT5T4gJJQeJywWussv9puml5vc5x6Tueq7+CpkwHSUuP5bJiE
9YA6KXSWBCWM+AY5aUufo31XfnB5sq9abFmOQY6E7SLlx6EVQJkeGFsXsP1kHPmR
mlVfVQwH9nMTqX6drBpRvQIZ3fvC5eZMX8UoC/SVYZhKFHF63GrUEaCo2jIWt+J1
DsCWkm6rF0EYHs7kMCygmaCotFyf5E+5Dm9xnEfJywLLtNXqL9oaCmX8osH/yil7
BL/x7Zuj3WQE8Nd2EstdG7NOVIQIPJC7tu4DUgCGX5S4qE02gnVHuUfEc9uqlwjX
tYoyG/4hO9z6x9zAWGlNjOCbzWxHiQKVx21j+Wr1lFDp3gaHIDLy4oMwDDolsm08
tM3S5z0ExVZzPtvOLD0uG+aaRyC9SuJt+N7Fg8p5b86sXkdxJzQqHfuocdWtVYkb
/BHwKobwYxkkNNdl7Q55Q94jinJ3TETAGtesxiI79KSllGGl/S+YkuhsOm/xIAJP
ho4Z2Dqp7p//v/mn0LFLuj33817p6fAtkn3oN5u/V7b2OVuS58pCPQYHdrpW117M
itmI7cvk93iQI/29VOuEgyy6Yp/Bk9IZtDg2XyZNnyF+BN7pLnOyKVLYlWSYKO3F
rclrV4BXLHhDEhhPaqaBhiRLVg4dEbNlR2ZKnRmfaExnOfGWuuHrpj9tGXjsodvX
m8z6bnexX/4mk6AGOPQ6yYlS3cIHU1bIq5vcuF0rYD8NZEm3aafrgABJnTA7Od4p
aLsURgj5r3gVRDSmyQtsbbwu88w9SyOhNQo7JC97FStgcVDbZh6uZ8Kq2Zkqfpm4
RxeNra9g5XaZzhQHVdY1tGXdm4EvH0fdWBW+wbCxwj1MFfBHArVCJzYHwJqiBaOs
Qe299IveGjOhSwYrpEvzznpBxVrAEL5uxxfT6e9qFaLm21XIh23OGjsrq1KQanur
i0sOSlu9R8PXKYs10f7IEIIcu5j7w+E1bDeCwqO3zLvag/zrwL9ckBiW6RjQKWpj
Nt8nVRaf0/lxMsn94z0BgcOtZZyRg+mQA6YSVOF70n5TyQPUziCLmOuqWDo0jn8/
8xQBNDKUTI2/5cqrAw81E1NfpRiN7J5mML5KYLnSRds2GWKx9FnMHoRhKGTBDYkL
DwJUFDThyP4KWq2ek+BOwanzq72GuO1pIZx2wBZjO8jOWjvVgNXTSoK/Oz+XRzwi
CcUwHD6PMpfoiUo9hbxJZ9rueZLJA7dA4UilNhyYQFMW/IJ+y10xH5dRjDVHnQ3I
6ptvVBoco5aKsed4MJNzPu9SsN96pL+K9Ii0Hsh71bmDZjZLhQYI+mqrwmC7xtDE
/CgSn1IhrHPH333Qgl44ZRkoLBCdxLB3+KUaDk/YXPFLBV1yYuybs5TbBMgDUddF
krsEz0U+2EexpAMkBB35b9zwP+CqAFvHc50TiN2yvFeIyl91m9iouLkmPN/u2wi0
XORDBKdedwPfvPDLWEWbo504vllGuSkn1ozCWL/FbEZzGhp8rGsTg4rqmu1HRwLA
cWA1zqyn2wYI1e1ypqxjYaKwa6qeXsBmqu7fev9tgJjC+Ef7htS0Gyl4iMO+pQsy
me/HuDX2IGYTqiDlJzRaBuHmMZEN1egQp6w1tpTQwTssOD/CEHtMYZ0ArMUmhzUL
v9is1UgNs3/sePn4UnJ6ckVGXCXpGH7MHi4gO5W+zR06HJkImmUFXanYiil8nyPc
b6Eki9CcH3t1Wiyy9Xd2k2CI9TfY0LTJlZBx6j3+3nWPh3p18F05OFsx0goESuQA
afujQlyRLyjoo1K+UYtrvrrboYCc7kW/Ptc6XG06dVAQoEPyW3Ens/tJ51tT8w7t
Wij6/Sand51QRFKGvKqEIdjMb9qYs8U+K6W3h7+sbYWezPoxAPtr1xR+9lKN3Eqt
tLaeBZF4mfUsmQyqFThQKnpEZgFO0obFXRre6YbZZTh8rk1FAkP9zNOIFEqa4wxH
hDHbIan4HAn26RaSbbt7D194GU8v7u4QCiOT320wBH4p8WNrRqJZ70SQFZdxi/B6
vJG3LNYG145jxjI3V1MiAjCKLbYmKJV6Qaf1xQLfMFfBTlaipxngl4ZJKgix5rbi
zp/ZGBFu3DR2+xa2a0Jjp5cORLAWwhPoB0bQ/wyn40KnBEZS26XqStN02nlYyJwF
lvG7MjDnFc2gp4ezd0wkBJSdvzMGGwdZ61M5zfqxU2xgEfZsHvBd44wKQrtZMDoS
nJeluz2h5CRa5pyA0uBqaJ2fPVf4cHzQBzQETyCMW1b9s1sYfglSqnJaOagzQGDl
xcHYipW3qpYHGjfUpURtkud5e9dmpvJo/bgOVW6V1dtx4/v5prdLUI6oTzvBgFXW
sVGsLUJcGhlH6wOsMhlOm44krKsVBIHJP9dNWRUeNKNPe0zDPjdw8ibZggb7/3dm
EDGPkDtCSGWg/ybZR0UUTwydSJDZV5AD0NHI8twc92/spVC2Rz5Zu9vE19OI0uOk
/joEyOnIfM67p0kNW9t1ohlPkp9SytHGUgYtQ5cWM3mEu8P0Lvg8RErIP6DaRohh
8D0DbfKxtigQ2ML3vTpITYkbG16xCOQ56vZqacI98nxbEsQPj5tZZWMfjXbEWvNj
OMCQMv0+HqALwg7vL4P9HyfS8lpbnoK42bcXR2XMzRPHpIJQ9EsK3ChEBeknTlW0
/hYBZ1pUGndX7kdSYwt0PiKx/Px1rm3rhPvdH8cykgVOPvMud1bjhQsIvvjN9Dvp
JuKMgXEImPvFzz6Wih9mdrLg0gU+a/nUhVDLl0p2TnJrQjQbEp+7Y9Qt3peW4F2a
sHMC5NJj0/JmkrD6zl+206JFAB/yrYZQaZZvGxJ3FahLkvaQpy/Rd7wbKDGCKfLW
cywKZ3zjtFWuYNI9LiLJVf9RlthrDIkRJKWtqxS0bwbRkJYtpbcJdhW8EV3Vup10
HTM+t3gveV8h6gzmaA69SUfAlxK/s1Xt+fCSQUUgOsbh1i16XRKs4nbzgcsmBunp
KI3eMK0RUPJNlolkdWhMYH4Z3t6CXxCoG3PjKgVaClYI4LAg+PA9rNGRPKvAo9ar
32UeVyO1wGbxT7zAec4ak/p7WQQnGCVkOU8hhQAmLSS9QWCKmN34Lz/7aqzTCVlW
aUHkMugnSDBw2wKXyGkhT6jsu1nmJSvOCO1RQCMGtZ59ile+EV5xCA6qBZcBgkv/
v1j4+lrybHnGv8xBz172rEGSyktjRFJdDpAHZJY5tacMfbUjIr9g26pQrMsCxLLO
Y/8nUhoPSxTmlbd9kFI2+EofgRrvTmG20Rx4+ISTIW3kfxVSTn5aIEDuVdWLLGnL
u7eic+innCt5hBZHIZS16zYeqxM+T1YHAjKZVHZW/6gI1JKp67oADamGQMwtm2n8
JQZGHIJqUGNe3MoYe6sklrZPFxEXgvce9wXncPUnXsmIgzy3i3Azv+4tCcmU2r63
bHkaRvmL0BvZl50xXmGLLHR0McGeYyoxedgEIhv+Y/E9AZbQAsLc2MMGeJd7WfaJ
eqRQZFgok5UGyQrDuTwQkA+LOZKa3Q3LBsb755GJh4z1h55kCNsxZ4mmJqnx3OPj
Z9Qu1vggpVuo/HpzLoSeqju9HcWLrLgJ/CeFrowLnJXFCwjsgRU7IZDRmAZBCWom
VTFqqv5g0BZhJbBjjF8ArfA4CPDwU3RRf2alrkPL6lCqQBghEb0Z1n+GK2KgpKDL
jK/7ckJ7YzOdZ8xbckoJp296ZDFxFcsafABGqw5IV9DsIr8aofRLnSs7pa5rhEQ1
134odDpVUouYC7s98Mdq9a6Wu/wVnGmOF2ijW1aNAKU0l9i8FZ96FI+XgjANb86m
1LYcpPN/xcvaVvTDdSKMVGVClUz0mhZkqaWk7CxhrKOrmtnvJ7dbF6+4mvC3LeJg
o3+NFck1Xm31iryXBE6z1hiy0Fhuh682XCE8uHEOiy+N6LUTXnwlV32LUWVvvAfZ
LpbnDW0WUSIRh1qrotN0E+5Zkcq92Z8XdULdl1hhtV7JYgYCtA9d6qlZno79X+v6
edID67RQGUoHbmtzUuVc9JGoD44pZ6uBjHbCD+3JsmyARv68/sIWofrGQDPZtaEJ
Ttnvmc+PS0HXtYofqf3lN5ZhwL2r0dH72wkncp+/XqUIiGrukEXHN8oen0J0MMMS
0ulfEek4dFxB0R6fIUjb3eLFTQC9OphWoDeQ3uaMTp9pvwVsT/whG3mexToZlKgL
iTO9ASbdAcggzKpeYJ5CUCP7DjHit6Jx8Yhxca6vAMzheyuot07Ii3wkeZKb0TvE
2fb0i8G4/ujONqWssDaBdWScGyaFwhJwe2WFHdJThmXyT8/crZSZbKMA7uk9zmPI
sl2C77zBz68B6/sZqqXscklm/SMWe+4xfeRQoNbw0IzDApgT0NfY5fDm7kEF50HD
CD1aANk4L+SW0AkudQ6GcFXRH7PFWMt915kr9KrUDE/Du6TlftUFqIcGjmKl17V3
YS+wkw8tvvYr2yRuzFjn7RrDDcFsL71utMiVM1m5Gk50qYrzRylnMjdR9xnI86RQ
b2TEkiO7lci4H2iyLGlvsCdVAPNAJetTSrU5G5euOAgkeC8Q7HdfQepR98axoNJB
5TOO8yoVIDzflvGNhJtTyEIt+VJSIIrvrZuq/TrD9sEGXpO+HZFEgoYtS+pE4Ns4
NqigOMZ77VKGXsNSnvA1ZUuaU3i930fonpqDiwYcgt3n/KRTzbGglpDy/aGAQNik
eEihDsSzrKDRnOe3980qhXLcMnbda1eaCwhM+kkbtw9z9WpyVmUzo6m0KGZaoG6K
fqox5Em8rABi5l9d9OcZsS/48WfyNgI65QQuU4rAE8AN5fRrQ5NtgGSWnY/rGKmQ
4olaxF9hNyE4eCqrf9kzuKqIHzN4RsACwAA8b2sUuRhn/ijR1KNQOjC7KxyqEqBV
C4utJi0fvwq91H4TMTefqg40y8Jt3fNcsY4ZbGN/UgNZjJwB7n+Wd07OgaUGZbPZ
D0bk4SO1NWVYZMtywzQFTlqTfnJ0ZRbCEt8s7AXur1eul9erc90YqAOuocEXYp5F
8odOa2cmsyFlQVrbXTU35E2An1uIzNa3o46sL0eUs72YYp1P6M44d4zrillIo16Q
WOBH81hLSEmJKF1x8tkIapZT5x/r5AuNRB2gpNfoqBHi25LaX/DsTsP6pGxH3vae
7uZp4N6KjjG3PCiufMO7LPt2k03gNuQ1ggrrnm/6hrqVWCZeBEkaEjRDS/c9ojUP
ueAPfPKJ5axrF79s/Zw3Oj6hWsr72Sb5xjyKaVNg41JH59MwXpqwS3cz+rmI9o1b
p1V3XFOfxMQVrfAn/yEjVGsS4hfib8vItlImeMBVBhirLwU6OmHUbLs023eneSrj
Dp4vEq59TfeNLY11m+uhOFmXx3GH6ypcLZRgb+2TKmBy7GgndH9J/AVvmeTDjftz
nYsL8BK1bSGBGDnZSWNtRX699xHcIiFGYWjomGj53ciTg6nCWZAhD6+mXOg2MqsV
bjMPPCgflJjGG3tdCN8w19IoIQIUDJCmCS24QYcRPM0HEIvWOuHuMS39ivKhiH7K
sOnqhKGWIUTA44ZVYodKcjBYrQ47W5ohF19Wrm0qExdfMq5I6Jp/IAKHLVokpgFd
S4HyURDEyKFjZGuKNpmqBtbAixvP7iUTNlX5T0YFHw+J0VkncBz9MQIf6Qt6f5uX
7AhzrSm4UGpCYqTY7FMxykIm9Ha0iTgoKzN6QzaRZx+AVkwxQxpobNFxG0Q2EG3x
zSU8AY21YGe5r0L60WKASuR8TrdWyhooTv6VDTVCrciIMrmLFOMADmTHYqizAfxw
bS2JATMxVFGQqN9pvgTPFbi5OX2sUgMf0vhhc5OZWOGoji+na7IltkHA2SdkhmNJ
xEnq+OoSaU2NzdyZdrzKxwZArtDNmro1EPN4sF/JL1wpJmpUYfhOZEHoFwqMzMTl
IeW2HSqu0op3W7/AH9ybbQ0ls83ar7nqDKivW0H8Mg2qTN1Ug2D9jSz+nuJyBd3F
pkjp2bB87kQUUsj+hyWmEIje7T+J+7HLmcqw0XxXt27aIHNC7ktraLcWETAlWzft
VY5cQLAqW6p1LjDe43EeKH6zNZezzqFVaFu7dFvm/8knX7YF/tgypmhPXq0mjA+v
fUgHfNIqn9B2GfAkNyp2QqERb8ZjW4hw2Bsi/4KkP+fkrWOlWCqSZc+fZ5dXnY1l
BWYhZCmUwMAJJoitydVDUJ7aZRA2fZcy/j7uh9jGm97bDpLNBYcZORACqQLz0gvA
b2xnP/NK+IWr+LffOfKz8e00s8R++BZlL+XXYHWrQN5ymYIOu77V+eaLFwrxor9M
HEQbqzlEz7oOY75Mlkn0CXLMCz96dPLySdeS0rl6a867nHtY1aedS5aSC22l7oKJ
2vCLGmQ0enWkUErFSfSTYr622fcRxIWfkH2/WxwW6D7n3MuW8TA9yIVubpQvCDLm
07x7ZlfdqdWHi0u30/wkOeouHYJwEC7C2SVoZxKEqkI/4/rUdpDxzOvBmLpRFKLH
OUnvNashaXDtcTsstiUyr5j0adHIuEs7dDZ2leUVhswT6HX2DhbeTmaWLDdNGJoz
ju6gYNlROOavAVanIYsn1WrkY/SQc+MM0B/u+FL2SmLrbvLKeUaJgm5bW9LdQRyU
YoogiRlgFhAiaRRlI9AGy4eUEJnpgrsjrjSKNaZzvmjnwmS5Ke9Sz8HBlakIWwYe
ZIfgSNllWWYsnT+suICyB7BcfpNS1b7fJM66g5ewvudijRfmobaGLgkX++QIPTUN
Tct+nhC/jbRJlsAJJcS1rK5r2gst3RF9EiZSPld90kNLV+NK1e2RfclsLQ9jQK+i
9vfaP+rklJWIirGxntQDLVA6MdV07aXheETL9EtXiDkEx6w+dYL0NxLy690RHsXu
dH8NXfD+8OagQMSUXkrrAVt6QP23MSg9iIvm3gPYubT7LkS+ImoHFiwt2z0dsEhY
/cADF8KJdRXreRgfkI+e446E06LdntiOH3r0WFjHgTru94t9hUiVI+gLW4We83HZ
8bNlJFks6kOErFPXFZjKZqm+Z5cJIN8lsU+AHISaXHmC0hm4oz4tND4rrF+4vfrC
iwE3B9vY9955lnONNDZRYOpMBH5l/fb8cpAfnDNxPnjDtx2cRhagOpBgcbn9V0Tk
Cg9dOVIKx1cGGxRwADr6kqgOGuFc/PIZLw1TTqjHRFfHUwWfl6RK6nluHrorwP5t
UeWeII/vAMZ1KI0IaxmzWz9hNWzVWpzEz6bl+olBFppjOXbuiqiPipe0RKxXyizL
w+tuUGsOfHfRxIS5X+C4HpztDx2Lnt3urBxP03ocT2BP+0bYv6gjMzEKozARVaN7
Budwae1/Qr2iDRuII0GEAICT9pt/ZBkQ4leABBgynAVclyFz32xLahNpcyNrvXtX
LmOAvBuLyonnhu78gOFn4401KVaar+2IHK6nyWyN7OqRCeAdIYBTuH5xCdMiSyM0
nHJz8rp2V4yYDFtmq8vfMaJH4SLir9AZ4Qw7krx5A/ekGnaBymId/dRBDIUMzAJn
VydPz25c70q49AD11LOleKOM05Ljk0ZYeLZ4YPTRkbnSGTDzJBQRSPGKMEhzCfsD
aT8thyEItdfsVgv6LF3qI7brrxx05b9+ZlI445lTLhZYOgVK5eNrTPZtmR/MRlQW
iv6o/6PJHcwV9ayfOsgULJzEd1n+Jl8sKug5yu5IM8IG2NJY40GYBtzihU9hwrh/
nxOsFRAZk3KRoapDHSSp/DEGHJyGpbl3zrHDeRLZFEf6D8OnQhYYaDg6Q/b+EJi/
YkV7YMstGKmfEBXZExuVQTLJ/3mmjwEZ3bv9htQmuAGcC1XowFc0Mb7JOfcDPYlM
npRteYThA0s5xop0jGqHfsVSF0jkzq3hJG7Vbtw1s/XUnfPcMOjLlT0A2x3ug8co
6zMKvvp78g6YrtlSgh/6tFrVgzjB+s3xlIIGo2bDi/26LFGEz/k3EKy3I3KaYBDW
npvUJ8SX8YY32nGYPl/MR/wWLFkwmLg5mOCUoWEO8mq6Sjafs2ZiKOZ3Xpo8gCxo
Jw3KsB3qLYv4qro4wTs19oaclJOVBUUJGIXO7gOv4nMjnEv/3ME99uIlWO/u1e4z
IspkvSbdQPTiIJCjjTLPqQdjnJ44KwU3Ng7X8xFB2IggxZMX0qOYAQUry2eaR2PI
atPrrUXwF669Fz1gmMWJMaPfWcKlQ2nKKWW0UUdY/ntNVd0IRMWcgTPxT8b0aoxI
Yqwi0tlELxBZL3IRcNsyQeDw03qquqrN4ZnXnegPpbqa6CsWCyBwON+f1d5Xn9li
zmYAlBxGhJt2nxgutfmhaJKEyR8+1doFfyRI/LqS0AtbZZ7l8pbFqYLjDlTZ3d9b
ENTCJzkl87N2oVrs8FqdNKlBSOtR0H0LZocsivn5jo8/zyC0hhyiuJSFFu+zjN/b
0MtdLR+kQ6S1fka2U6YXS5q5eOmT18aWA5e7lGmZKc0wZv5xkyHi9F1b6JXwQeO5
ItTJ6SQFg0cTaS2oZgMsMreoVnFpu9VVgVsTps+fijnjzZZLwtzEoO6TH/XNnPKO
TQ2BQqXaX7bGZWk/yhuWFo1kLBYTGkM+w/E6rCc/fE+R12aDmrfuqSBB4p78KdnP
p3E6Cw5NE3EGMtQjnEivDSzjDZE1ocdTEZ9ki1Ysn6pU38hc5nrvuVTSlff6uQXY
+ZTOAPzZvr8X1G3wO4BCfPK98wNcbNDw4wss3rUIIbav7Hw6PbHjkkdfjr3fX2YI
3mngWTsLEIePyEPkHDM8cNOIuS/O4GwDRpu+GlmQ1N/ZZIpHJSX8oNJ5Cpo4mSa9
Gb+tXBeg+GJ0JufTMmarzFJFcaokDbFGPnA74kc8kRqKPYMn+L1olqgMTzMbexmF
t2EpIro7ZjMUAi0xHpZtKD5oYn/rLsc4ZU0UZJneAlkXKxDD9r4zYUYHk3+w/sUr
uEgYSDv3vejAHIbmwaKvDBs4iM5eMeqIHDfLiZ4ecIBLki95K6X7ZhXc683LIAQ1
JzPdsySWxX/X3wL7H0+xXHq882iIFx5rydCWEMEaLYQm2HVPByjqFL4r5CQOXUWH
hseniIcqNlVa+cKLkcRy+MaCbgnFkN0gU88Exybe7b2LQXK/b82TWW/NFFB6aeQw
DYD4xv89CYIeunz/j4L5GO88PLB7LsV3jgzpvyubnvB2eOP5oufFfaVssrqiIJ7g
vvo8Hfh/9u+mEs/oXrQQ4DJe2Z1XMYugqzjbFGPRNWli5cXylOXzK18zNU9bSbJv
sBsavl6KdJIya/jwLhkD2fdkhsBlAvitLL4xAihZW3yBx17AqoFmhAilMbVeUPWi
WySg63zGEbwyaw7R7zyeuj5BFrFFu4RSBME7qS2+Q3J7hOa0+Cf7QZg/35egpfm/
02+hH+soDZd/OHV5S3+/uAlIikX0oOdJARozUoYzY3q51l8+mjfbkAWdWdyXSmVa
VfGL+JzX1tPnoLRm5LCW+O47C0d+mvzgDi5cicuzXvzFDYbPWxDaOVOjRQ2/gkYE
pj/FshfjjZylsYZIF63rUKIly9sZkOvDpACGQY2RPEDvTl/fMU7RTUeQIbs7owKY
eZSPa58Pnfj8vkEdZfIjP26zcOHeLKETc34h9uDYZF/3o0vhiTToiz/YbS5pumWD
Ll2+gNcEoO30yIspj65UnZ0rqQEaL/VkLcI+peBDWnkuNRptm+WFtGwmAu9Mtjbx
K8lHIHZLToWz3kFpoRk92lSzEVbfVXFYQBiaLQCthUV/iBVismojGDoS66qX8kwy
y0LN58LgQrQgDGcOixKgtEBCqwztJD3pAX+HrhTDYRGn4FyLvg0M+BgmivDJblQ+
nwFPe/pUkUjn828XTPeC4RV5cEB86EiZ5OWt7Yurz8HF9srFRgBp2+cD/pBK323Z
c6l5osARhIZ3HrtHv9wa5AUH4SbUP3kCnQxme7xvegePJTA+Lztx6V8tnJTQAVt/
KxRbb99nMISArvZBOdT2vfg363Re8QWVb784heCLiN8UaEzU4rnkT7VfBk3wcg1C
V/ABl7E8ix6yeK1a0VlXKIGYualqNbJYHSyPZAsTSS0dVr6C+gXHOGZNKbmm7OJV
5CnBFae46azRz7ESj/qgo6GgyjJvFGQVwYnif8gJGUVIVB6/TiWtOZNfdZ1qGgwJ
fohGFHfQuaLmj0MngccOZa7ABWRp/m3T/CbRqTcKo3REFZiCkO6FgI7sQsvWQOaT
3v11YAa+WmgDwJbfFL6zXIRWiPmbspr1SWdXysduaftajEulBZezHNBkexsRpZph
aFsTJwtN7mcFyemgF5sayiQ5X26g4LarB2oNMY2hrCFWqu2ot8NcSy3h6i9HDgdk
jyU0EtNLAwfneuLE/PJCnUE5ObKaE6+E1tMZ5jzN49NJLOD1h25gSyatv2itRaLF
GYig5rdDK0a1ZlDSPdrsP217io4TL5EruBQIOCPVqttsvCNfxtLcCrH2nq6L7YS8
m3uUvJkONL1LWFWL/GIOIBcQ5QUqPtczHtu3gPjQLxh3FYdsKSfJdhyNNfUSzuKA
3RpdSW/q7RitkJ3lX1SXSp+NrzCX6SauAzFTTeOu2spyaYz4/mEbfIvj1UQJYxBt
HSDc2dvUFuLMGV8+SJymT6MUj465NB3aOHKhk0QcLtdLMvEFDK4U8wjxSMrlUCf8
K94lL6psrQTQ3/LvxqtOH58H7STlSht/5PqSvTkhukD5BNYwBBHVIb+Du7O9LL3x
JB12hsrjUTueRBjfs2UgBJWCeWoZ9TYPT+eIe94kazSyDQIlVc060B+CHyL3NxRU
g8iKKovw36VNabN02HSSh7NAUHmQiz72BBTY/2SxjE/hPlewOviZQ+9fUnmDOj6K
QWUkpCObfkxXZePCXfEqanhNBOkp1eovofuJ3a2yJFSsF2LUocvWqB67EI6rJDBp
sk5rvTHE3B4elxpdbdFTm1xbixnMMjs6uUvGA9NZwhBLxL9XLIYUCLT+xNNFfBQi
/owrBFqpWMYB5fE+F10teNg03I+YkspiPf6LZ9MnpuBaOOzGtqIhA/XPZ6rJ/YO4
GYQIk2GF5B6lECA5aZlzxAGGwt08tNYvQ+tR17xShJDudvRUWX/bqSqpjyEgfcgF
eJiUVSiZ9Pb2e2FrFvwr6r7DVBA04OM62vjz6SItFVDnaBRqWP87dmRKqcKW6Ftf
l82IkdPkbYHqljGycdH5xCpgCFK/Wg/AJ7FAOpY0XxcbRaq1Bwu8T1GzTdAqZhxe
MZmXsXMHBxBpmgmAnUxhsiFvFfuFTXribpugn0u6cilIzWPj8LgmPui5pLxLVKZp
ItadKmMIVzsCU3pDCeZCSnJPm0/cq2LYWzCxxyuw8zsHCGLIHlxjCHaerXuHdj/g
dV/sJthwyCIViF7SrKPaEFJQ93GJwljFKa7H2E/e005FEIsMoeWfg3TvY3UDa8NF
UMbi3lYm0eYw8zv/NtOk1oJoUhVVE1LZ6rXpWgbE46XNYHbvtB77TYL7dAwO7bAb
qntuTJKfD7H+SBg0qyRqOWRt/d/sN0G7GucTTvm7yjoHRVh8WVvY/9FiGYTgHqUQ
PWIATMvUnpYzX7Xoayqq+ljTSEENeS6BUUnpxAXswxXDSTMf9O6va0JQny9Rlvg+
jsF5DuzSthuENaXn/OAcQz1xuZ0qTogh6jsrg3nQ7QI5c1KXlfx+xan9fYrZIrXC
77P78I2V4IrelJddPouAaw/bAz1nXMTuqPUAUsjD6s4JBrrLYrKD2alCUltP07TX
xd9Mgz4omhxogS42IAimyB4kd8GEopQq+vb1zeoaSYLh4uhwEkCfZP1QwYSAVQeP
ONCi8/ejlEWq3lhbSaL1/eFYagV9DDEd7uTywHUa6mm03TfC2BB90YzaG6ecEUn7
xF6jsy41M7pOvnNdOlmuGCpbA+xF8t3oTNfGQohfANpSNga+rD/72D/oJrUgvM0a
T/OtMTAt5fXOL3FL/zIImPNbyxXwx7G3+Bhumm9gqkizW+eRwMZd3EC8h6eEjzS2
8ltuttwJtRkP6/xFNMgNtsicpFxC7kJiG2Ilfcm0WL+yPdwxD8OjtiZw9UU2a9zL
ABelzHK3vWBSx5l2vcQD2LLTvbZlOyF1t0EwjCPhKaO39LlpJvOiydHX3nD5VKSx
OBB+c6dpnMJbYK/dIMGt2hFr2Dtj7KKhJzXc5RO6AUpuo311oqMGtz1Lg82xkdx4
1Mp3BTYiicpj0/sLAM7zbPEI7qk1aWArJvomqFxxxUNfecya2f2xkeG05tx0Yr/n
FnE3x00qTtUWHJde7EltU/B/ETVot28IAmlhUZHBD2C+O7UDH+/9YDT6oRLs7xj9
KLoprNnoas//yLIO1DeLsh3HJcoC1wR5JCt6iXkfi3SMQXPO+p1XQ00ne/emDKBu
EbaGoUyg/QsTddolpnce8HeETGPAqWNTLc3HGM8abBf6ECt59Xfe00/rK2a150dl
PbMd5Y+bFTxbu4dRzn2GKGZf3pToaeieMxAw7YFDGFKUfYINV0FN5qzbnNKj0cP9
btfmswMV5ufXPzd5+jGSMWu/4vDbGwoRVEe5N04x3Rkh8ZkhfGEr5yLvVFRWrZG5
emAW87gtw9+GDhPeOJidloMpQBE9gBIrvROD7sqtDI9M+tystzPf0/q5+E8i+hI8
QzOsfb56pGMEbH6nnexEBsfm4VxV1HLSh7gYaT1oYFnDv87eqb894xt6aKcHyhkl
4HIYNgHlrkSP9uBTM50PIeDE/7vCQmm0I4bJ2nsEI+IeKWvEdhxHMmdip2WqLfuF
HiXxLa/EuJIZcI0DMBt56eQ7qIT2A0Rgb43SehrnYTCliTwKd9NyA0VFNDJ2s2Sn
PNjbx+Gj1P+Tpm8ktqnkVhliMh/C9ceZ54n4d/ahI+DYFGB0Xxqj1Czazd2UM4df
ilw2zUSw7eD0dJg8cvd+KkWFHxV4kkWFf+CrzIHElo07rUkGEsj8fUbc7tBCLuf1
Jrl7SPlRtQQj+VPW6IUySQVyoeaEp48oAl+O4irlHNIwB8b18NnrXA4i4Y1gHVdL
c/AJVP593Sw9SPxpQSQ8DCausyNbJgweOitjVwbrH9eBBTgTYHL7PpBwh1StyyWa
zdFj/EZWPwYXm0eHY7eC/QNbViCOGaziS7TnucIvC7m77eGLB4AGDYc16mdP49Ou
v8rmOWnp1lDSZUkHLOiCD+DoOhK4FhdpiCS5DCYxyUPQOVw7pfaSSSZdCtAxko+W
X0iXe0tIf3obGKwuJzS9yg1eEa0PaQgBbSLEnYhl0XVExyK9IYoxNo+evMWGryLD
OXczsZn0RdIaziP1hstaJqenwWh65tLKF5BMqcBmFli2YJHzUJEdd99/tvbb6ipn
wlWB+JqefYhr23ySYKQAZQmg6j90BoiFkbarf6t/kKoNJu6VifLHf8xnfO+ye0UP
frBcfVviAUnL/YLgjZsXkn4b1gO1mRbT8zgagFuJLAPELCi8S6cQFfksl2gN4gMC
phN+xH10p4Trk9wqBtAH2k0oh4Mf4CNuGmG6lAnj2XHwOfVkqEtFP4wu58GMOrLi
vxd7taonTi3lb2qEMFyRcBXBbwLzUwZWDwlA5jM0we3VJnmTlgZAQQukQ5zVK6Nw
Znuv4L73+JEbSNivA79xBV9JJvnQUEcchXwSxtYBWrMA8YYYsewWaG0IrGSUEcDV
zQHem8aIepTMcikXJnQlBJMpTa28xIwgpWXLKxbDXT3pcuubwvQLDcoP4BCxk6+Z
Qzg6x1Ob8K1O6rk56rw0QX8ka5U1aZo97JKkMSe/DnZaQFSoSxVOU4PQs2WHxE9i
D+8wtVU9+/9xf54vt+lN8Wt2gOTFD/CwMp63GrTuGOv1tej8xgzUtnxpqQjvOskd
E3kvuZ6mSZ7uPsgXBcUCu3bP9t64xg2MFWwC2kGihCTfUzTumOsyb+TBn+RmlxHu
EuZ7BKifVQeo+YGmRatVI9M+6oju5V/8ebKDX7KNqbjhqsc+yNWNkICETp/9UwEq
QOfONyjeZ3ZPKX5k/Kp7OWywREwYvosPoLQwLglwY2MlgidVuvlUsi9xiOVuYU3q
15QEA0IQVbGxEWVsASLcIwNg8FRbsTj5FynTqx6mqEei2eudOJCtSavthNxH2oxE
JtxMa3CSj+eJKN7DOw3Lbaz+TJexjmzGe7JcmeBLh9ynvn18mfmW6g961tf4cjUz
bAlbiRvubR+tsJMc8UZt96UXaIl5wf15dXM+i5q3yo94hNqyiioLY6Z8U+PUDwxP
W1FayvdzDiCtlSzD92x+5TRP0RBZhBKxvZgPwHanPJs/+mSurpptGdWcHMLO8QyO
prlp8HgbNnl6Jr7U9lZnLOlbouMoNBeHsANXw/0UobNsgxmgq69yo61WTxljiVS8
XAoegawEFz2b5gpoJEhqOIm55UzLRtnm16GHmxTT990y4aeKWAJUHHVQOx6XCrPj
eOcGFqG38ffd8x2MuLafTzdH+QOCtJSXPhIxJSuIseuf7JGirZUTZ7xrPZB6dUtd
US8hCHA5HqLzp83eWCrQzHO47jZS8b/5XuHhTZ9Popeu9CLgecMq1ynGQ2+nrMHM
rAJX4lLvE6fDgvX1Xgu8GdMw3DNtiQ49l4SMlQt8J9HklZAiEa/wFgddhv46+jt1
rhGTkcDsRTqJBX4Wyw/4pEPDPiT9K6J6SX6UIb5DuL/7wXdAqFnPvjFRk5O+S80V
SGF0xeY0fMp70gpcMurmdXRHWLBOJny5typbXq8s9dFVD3LUbEmlNFz6taKGlLT4
oyHY58CUIaJu6E2Su/Ei06C1YbgyHsFist2aMsiLht+Cm+rPk29lLPJ67ShTq2bf
BW7SYD+e7omhUepwbmKN1qN0hkRTzkP43LDEHf+TNPkdbwW6RsBCA5eM4pSZIgk2
Att+1GwQz8cPYghqGoKMP8NBGQHIp0T+K79hfE2cpI6e9HY+SPjVbXWogtQcryAn
C1dQUxn8j1j16DrFTvHFFmhOkQkgykBikRb703tXEIaEb0cscY4GpAo+rYceAOca
TfSdKqVmkLTVi+vrt3FfVCNevljYeQagunrkRs3ZQmniLq9c2vlxEVUR/FilWzLJ
S9TO0AiZ00L/Qb8ZqkA4hZF2+sMuJt8f2iDaikrREBkyOIozgNff3pa3Tiu78Xp7
merNjKZDqhTQLkCA5L51BMW6xp0TRmUmLK2lufVjvXxTKaKYr4ARS2bNJApfu+PD
ny0c5kKO0j8e8yPUo1wHVidFc9dU9IsmdL0Gn3qvehkXJ0pXM6MDgCKdyP376Mlg
EciwWxErxDfbuub4bbj5z85GFCKCejKXzNLBpb9b+PAHyZt0G81OKsQ90i8Glxoy
LNRyZsR2tguDJKSq0TgIBElUVMmfV4oEWboSVVrHZ9sOs4Zt5SQxVthDxtwadId6
uoH/25HwnHP5S5A3brsFBNY9J8kmtc4XXoh7tPozXlSJY++Z5IChN4gJqCsuwbwz
/kkfE/FlDYXjpS1nPCrGBRDw/6syz8xiEqbK0KdUa83sZb23oKIm1OcC36BeDv5T
YGo4MeYZCD38ggpGGzvRkH5eLDtzqo5eM/AG9waDosIBt6M222/pYcF8MZ7q7ONo
ps2S77BHrS+leaxtmuShgkIDLQW8zyZ9QZTCZkDQwkUQIfnA3XF0HQMmTLdr6Pg4
zgKoO6soYBdI3gVedClcGIGOsSkWTCyVdD1c9AK1CUITXeaeDQkKQgFVZitEnv2J
zDECvWYxnljYEhJB5Nj0yHeEcPgdcw+Iiw6GlZKgO18qXDdnCjcz/ge+iOvHbD3j
u05JlwskvloBHWPPIoMy3FupvzlfOxTtF4PJ14Dta7rOXPwwY3IwXk0dpdhSjfFg
2/rLaYUM1rtcp3Z0HniUfbLzeQmWQj2j5kMci8dspBt5GbUM72/bf+qOGpC9MEW2
SZpe/RndfJc09JZYeMqY975m576U5GfsTBPWZ6H1MxMoYKR7H2KpKPSk65G9dKUw
xruQc+TVNq2koPudGj83w5cFD5n+DKL0XjcLrAvkR1Rlbrj3VuufMSXZShaiXRD5
Io7iej+L6uG0L2sY2mwAjCEm1Tq1Zhn2YfbMt0uJruYgBmoAttURRcu6UC/kO63T
0gUTUsd9RHMqunCSutnd1Ot4zicAioAo87ktvNdkKV5m+SbgBcltGOb/EtiH3Qph
rpsgVOvMv7k2REzA//SisFHELcOoFsQfKiCFvlVmgIq/EyEVh9Djb7/LwoXWerKf
XjSaAXOFqMbQSPXA7UAwPDYRURZxJNIMuO3gU1mJJUEnjsJj8XqwZbRnktpMuDVx
AXtQRfB61T/38z4MakH7/LHttt8wj+46QI0SVTykBBHWv81hR9KXS09yM/RSzC9a
tX/vxtK6zpc/NZRgN74E2PKdL7wst4RIUzzkDhu3qJnWFPIqGDv0+FeUmKA7m644
HCzQ15/BP6sUl5yNWfs9v3+p5iSUCcWKfLMuXrkCmujol+lu3wAE18CgbFVdQKEr
9fbup9c7oSA89EopTOYdTODWBFIjoAA+4yXPEwilHjJ0TY48/9rsf5GhXW608M0Y
L2rGmWUdD8eRWd+4fKni9TUXLEXY99EaULo8too1lb+rPWU+rYNtNgC6yP4AwiXi
RZIS7YaS+7FMlvgZ2ybuYQF88TI8lLefWffKmYyaRjxNJQRD70PgFD1RFaJZKUok
wkWcY8wRbxROLuPBLxjCN2jRpnWrllwlKGizawiuJawatf9wulf1IbYV7To7MGXA
whEMwBx3fDNgRTip9dW6hClon7dcUUJ6vtWnk8V9yld4PVLHAiQZd7YIurATp2b+
Jf8QG+cfpbAK9TxQyVLYDaD+pcp7SzH6ECA0Vp1VQJDukKewf/sQixmFLqWSh8b0
nqZKAlpNR87rdfgeqAbLihXngs9f7+uTZaryn/wSQXHOOiD54tw46hEkWr6tZpjZ
SO9GHWxBpZUQlbLcSfzosIXhC7jU+QKqXahc8VNThwaNgYhWVrGVaD7srRvqHmzV
UqT7FJACqOvLJsoxJhI8YIGYzUw0Tt8dqRSJgo/DUF6vVfCTvY2EwgjhFGk2tiHM
xS00JjLI8Nd/t0Jtf3sZ+kkowYnP6ecM43fIISddiGX0GjdHuCPYE5FZIJ9vLh8D
a+nnbZxJr80Ayc7PQOrlKXXFPKORjHpaz6jw98y0xPT+ZIDLtkPbv/e51/g06BEg
rdqWMGGR/vtewHlHKtMYsH+z7kXu0peexlzjG93kekADRonTc7rVHxNNhMnMO6lk
QoTTpBKuWkTG+4Jt6/9D5MOkb2YB4mPfxBWHmk/7tMYHse6nugTrNZPXewSCBPBw
FXgrxoBa0zfGVRVDQx+xcreYOPQbRovt5kzdyZuskXRJfPXLGtKRmrQrk/s6oLXE
8IeuHjwSYntqNa1Iq469sJhYfzDC32+2LFRXR4WeEZu2EVmhSVguXqw4s4qCQ0XX
7Pxp/bztMQry/MuvHLFjEEt1SJBUgdF0A12BtA8dWTKyi8YJo8BFgpBRT8PTGJ4n
vQBZElVnslpsdh1HOBCAbV0UzhX4OSPOX69q0xGeIyAULpyhrpA8lzD+FAotJ1d/
o0OTE46SiJ8grFFOS/YMcXJLWFMmrnFLiGVE2H20Xzi5GE3ztPtp4px+dFOEMc+3
8DQ10zpbRTYCTZUf10EP2kO2u54g2bve5K5rVWWWmAst3V1Y6uxZRdgnS8ttbs9C
PSsy115KNfo2KNwvu9AlUtsUUhKyyujmOGyOFlpNsMhOEDi66Q2gdkdkCtD74Z/f
7tnstiTOGE0I1zhWwM8BK7GQgn9M7m4lCEXjc/fK2HDRM8cVIhDjnOrRj31jyCQi
FTwkn47uRmGM7DqtZVVMnO2iTb/EwLBqGAWMOMbqBchu19t4b0pmd4u/+3cMHCrk
+a5XnEecwhyyuw9nQ4usIkEiRQk4NZMapMfeiNHj9ZCHvMnhHMT3SO0OQgIVh5a1
sj+GN4v6mIIo0SGwRLfJzIs11SX6bcgO6Um3vhdjlH1yiaXZSVITMy8tv62fMJLk
KpmREWJYzY1h7xP7dlwaXm7cBnZL64hvSCU9v8E1fpQD6D6OVhfIHoG1Cfixq5UN
xt4MvwE2HQX2GfcLNoQsP3TV94CQ7VeTRyko6nsqsWvVyNgtnliOaz6l90TsqzUw
q7F26WMCTRd67bXA+jEnHfhBPG1yCqM/Or+3oIMuqmaOerAfeDRnTZsuh06lgdua
1UYdtwkjyESPEyTRuMThjsicrOXYTHRDObnTXNxsZXLRfNikWeJIEYWS9iSl9cwm
HxqgSGPSPpAPKmId7u6sxGKKIJ6anYYjL+R/j0JAyj7gDJrK2EwuaunSI6afOcdi
4TKuPQb7jwHT4LmvOiJJ1a9Z8VdOojrVGz/Lfkg4NplsRdCtSSJSIKAtUPo4M2jD
9SI4UajtxygdYsMXw8ZNOuqjEI7v3gkZbqYhoP1pIKaZv1T64tTj1S0GHJ0jRBBV
qMEjyeL9l2hfJut55PZeWVFup9bEP5ORmJ+42UZxOFkVNMYF44tyN3jsOhP8DRrA
avUwAQxnaH5Pfzb5t+u7spKif71TvF3JTlnaEt+kjl0ZSVSMfnI0uP5PPdzOZ9YI
HJsys2u46BT19oj5OGItgyq3tPOuyPh/u88etAKptan+b32O4xaigN3rBWAlLYa/
EMjADV9Q+T4t0Kljr0sFnJ/XBYOpSFXuhqvf+EdGnqMaeQ0OQSEzimLczTWA7Fkl
H40MxBKTkZxo3t3TFenkaHHdIeRpT83UbkbuvhOJHwGzDzB70w8WpCy8juEj8ySx
wlcQb8HAu/5k8IdM9/JPlqQx7s59KMYK28xsPK+mEVfnJwa6MNVabNi6tbNtFBhp
rxVJ/3YOjgg4kKaMzmA83pViH5WUMr5qnFm/OafSX26tgYGL15IufgmJH+na1EDy
vtsmBOAqvdKhT9XnZcU9B2X6TfOiGkLFXrJuRhuLPvH7rdYpkOEg+rCXHWpKfLdB
FQQKP0EhkdzlEBVxmq/HFzgU9kxgZbvjc26CyH7kNhPvifWg/t45K+e9UmljlCWF
YUjRmzswm2zM5vsL5Leu+/HQIsBck2ZJ0p9FH+Zj967zZ2m7bpucYLnNH3kRpORL
aE+kWPS/sIfuRRU8h5xJsfyrHyMpXvprkaMEIAmK8dyZlQpwie/9eCtkez4eDxt+
YKAWyXntZnnrm07HRSBGZUFyVRm5E0jyDBmqCAOrHdJX/UaYmTkeAy+LAHeFNf+s
7gTweGQY44CJhExmH5j3IBdcPsmKBEdwSFDEj4ilimclvdo99TryJuXkhUIP5TfG
rYiIu6YES68GcgGdUoi8lqi6atk3vMgwNRdMfCoxwrx+hWIIy05YBZUfVG6rMzNQ
gctKkqQdI94a9v9HB6SEnj+W1GJRkPrb1gnFU+wjOSvQLS/aMkWZA0Ll3orkwP0n
WzzjhWByvvhN9jiU04yW3Lc1x4arVyGtgePg3T2MzeIVU2vz2PF2bSF5+R7QbuRS
8lMAkO3ODJt3PCijmS6nJzfIrX2hMvWphi6jxfmx2cVWV+EF1079O7ZlRHUqLKkj
F96rVYBjXp3XC1O1ir4X/0mujZJ/ZTH3DcmQhNaJyw2YBVtjynh9OwNMO4JkBox7
XGt/Kx/8m/J9ZLLxi9p6snLFRrENrJwXYSotUBoHGc2dGs1ewGjxX9IQMOuGXEi9
oS1gIMBtiRrSA01CkZdxl33w4fMpCHbBmXcodmMlEP3tBMLNrcwbDTuYKSxkP3GO
SWIZOc0P39a9e9YDCFdChN9yXnqetzxMZdwVkIwm2DKX8K9DJaVSKutnBcDSXDGZ
sZcE7d4oeIuAZlcQ2DHLC4wizRJNU7HGt0KbxHJyhgnGDOATS4e1xROXtNkEA+Wp
oQqp58BlKio8v9CF4mkOdixDxGDXW+yr1gjj0yHtTaNr4FCXLUVb0ar1mrtkuL9o
D6/7QW7R8yJaIyxTHppKFOrhk1r+6naroNrevSPqYGtj6vbe7w1VzI/9s5MiGrTI
JseQBTaU46DjN0wxtAcMf2RivgwlwSSDAqOo7ti9oKkccMIK9504OcyaEyvRFsT/
sLdM4XweKAUkmzDlnn392uPy+KM4g5puu2U5AUdEiVP/DBwKvHW4ugTDq21uYT6H
+BdAvCb9nlwfhediXGQScegku11V/C6fbjEWupNir2mxDfobYQfQUEXSJvr2Teg8
XMVGZDFtN1pVQXc9HVJ8Js0X/pWe0nQhW/S8Zukyx6P5dZ2n13VqeM0ZpLWeJxaC
KPAGnctYnpuVCaF7gaWte6UslcSuShzMzj4ce4Dmd1GU2pkaWBZRYtO/TbhGerEU
t1o6+MMTCK+zWaEzW3EXlhXmxRX1QRS7egF1XxEmWJ3yKh8v8cNq6MKocOmSZn8S
ECtzBoEZgPN/lI7gaEEMJ5m2ev9QmdLdQT+EPnfWkEskMzwcjojAL9cg5jSdn4Ax
pM0ra2dySxYxEMSLrvKjkNkWSTuUtjpxJv0yfd7OOaO4sCFcjkiBTy0pb+S6a0GV
DXnqiCpnDBaQm49oYiWHSvYVlXMr9WHqIkIIHZfC2MVbHKnc9CxD4vpj+dZznaMl
H+yoQt4LHnPobFhEEiwRpMoy3IYMh9tjFNf+U0n+LicqRB46VLNMfCumUKVRQ1jP
McEwcr4hA+lm4qHxaYTgc7VgamGxp+x/24nWf5MRKK/R2rCSOxwKQ6EL0leLzC7z
xBpE3igtiO3gaBKTmJr6JhxHk74Rkc1PUEqUyvLal7iGKwMOyt6Kek+l6g8D2rw7
9zqOhMdVBLUISPGO7IcH5YZF+R4c/djuYZ24OTiIcOTlkrcsjpl23ZJSJTfbvEM1
QYJYMS3cA9ylvY+wxHl4XZA1bq3cbe8SQx6ogkcdLe2Dujp0gGYO9vj7vZj54esm
JY58ozKaegl9Z5k3Lr9nRYNiHOWN0nHIgvIonSdqZ5dk8ywUkQJ37KRDLRrWPggI
42KZFnRvClZSl/Tlo7T5qgfZZbEdYfOGZETXNMSJtVS07zwbZPr1jD/HCmELPX1t
04Sgp5nYxN/e781RXj4DXfF1SRRGNQkLjmNxFVFM8HZPDeywZF7OPfVsnJ/x5VDD
LD33jug9+evtJ5vKV5nU5fmyXnf42KwiNinldXJ/3lbaRZXf9ZZ4mio1Otis7lVO
8QoTrqozF2IH02M7yvhLKyaujYA3pRt+4jb5EBGY4EiQm/b0bPuHe+o5+NWMyH9H
8ESksg5hjkR4Umxa2wS25gpS1hVQeo5ACH4DcgkDq3Cv1M98QxPiqqs3ZmNXxWm4
kYV8vhgvophTIqMH4CZpZeGHdbYPny3P+zR836b2e4+VG8nBKzsWyTievCSxwKcU
0QUP1WHSWRBQ1nx7oyXap19/Oz1VDpF8PRCbyR+8dGCuLqmFpvkhvZQEg5oVa7Tu
NKnwgtg+Kepaliy0LWeuuUKTgTYPWIv5WE7IVcxfyNZBSHN4z4G6rVK/bhjXLBEd
seZuDrSSKcKI4dGFGRyOdn5vQA+oUcviPxNq5VUTZPI71WBKU8JYzsn/n9NzMHGB
d6d3hJVeeHt+uXMKsAdHACrLJIum+F0nX1FrH8FpGTKNvr8tHyPdDboaYQI0Fpwg
3AtcVlpEF97kMmy/NpuujRSC+mTqsynwBOITPqGJIxyOWKjX2g1unqpxLtnmYnRo
mTQE8hv2DHxK/d08LelsNc8xwzE2G8sGVO8O7GeEhBjChWCRrUrS7RfkfkHdzXD7
wKqXc2dJtnNAFFR56NDatBjTZNU8ISMmxGTPA+CPz49zw1uiDu4wQi1iKlmkkzmm
vFEXhUHeeZbJzuliKPgy87VrHhQEmBlsZbgf8yb7j97Qh7833ymJonF6d9CJUdP8
xBETcdyxjs1V4mbHjHoI7zTNc15cm7Qq0poHspY9VLv/Ydxywg0JKepfpIPeDSnd
DyK5rKGDYzSG8wLHDu0ozY0wpPR5PPP7rmXivMjL3ceuKI1t30Gx8Nyv1L4kWWZ6
gUMZtKGi13xZzZUuCG+12rGePrji1rlh0YzwRRe89VLdtXjOmlr6eKE9adMUYb2Q
YoS5XGDONHK80nNEqS5noODIWVVUkWM6UQNBfOMp2ROh2LRm77nl33mGl1lS91oj
+pWcb1JmnKyQ6DNWb1NF7QBLJ8SSo1bs8NkRVjsuh+xzL1rzAUqqvRSV7sIZza2P
Cq3qGEMeU0XYSYO1M6QKAu7EkVcr/QV1cD8bLWh5EeU26Crw8etqCByESltWD+GO
N+mtGGD9zkuCmv+QmtPuVACZbhN68Kkydph9SUX19wj1Qkx1eIQ+YAHZFJIARgMs
vrM6dCI1kGYCvPDsM7X+UORI2tWQ8mVEX6TD5gTinhckQmDX5foyeGmBGeYVrW4j
2YgCndOZGK2xkmCxVErqKxM7l8BtS/a1Mw3TtFIchwWonMEHoi7bECs5joDaI7vH
DaDMUYMIHfmzxkBDsCtaToei5AOf/XZMungI0hCzzipO3jDAbeJ6qgJ6aCat1UF1
ie2Ei7FQTr7hpNMrdRQZK+TzeJaxHr1DYE7hjHHAjby3TUsBWBXkWByfudwlyCB/
jJyoxtht9hnswhgoYIpoi/qvKxfPD1l4gcU3a5x2dSdweAg5sS0NxsDLd+sFcUH1
0Bd7e2ZOZgd5oR49qOZ0SNnVQCj3Z4oYlr4PofItiBCnlXVm8ncDg+Xrf4hjE/1T
4pHead50cgFiJrrMgFvG+VvSuFDczJmz8nRJVORo3IzbmRSvUGOd+hWr22eyMJvq
ZunH8Qd+H1cUeNGvgvPvrQzAb7vWPwliOyHP6kw8YQzh/coc9NJWfGX92+UMhsrj
YlmbdfpHyNemz8GCh8BcFIxeZs5Uo0OyWsiK4DFCCeff3pnaqZsjHR3fBDV/3D6q
sVEcqUmxYPuXv+Z+aY0vIaxCcylKsAvtFHtkO44uTkGZv0tpoXm1XkG03ayHeqG4
VrUmCfTOR3g6zNikm6T+qGXmFI7CW50cDycADDgVUFFg+5QkPdQNjLSxzhNsVf3r
y326har8xdxu/oQI8BJCfFhEW6mSVIbf4E+UdtGDlPLb9UnAFQL3EfGE68Ht5IZq
infSzYL/qo4EMqOPu82QjMKmM28qDdTw9/EyUwYt0vKTHcW7jtQ9vH0mOtCmQ0iT
72nFiABBFnKVeAuc1wWViZIqCdBkaUXFEMT7SzhzENUju7Gfi6L2lK/gdU0BB2n6
aVMSQlPfawvnPatS+Keej6kzMTBtulECiwblde9vNYgn/3n2JqVljkYWwnTPwODj
/hAZiiq8Veij29kSHYuaV0+1utliKmdLntn8kgT4hrtEdJ2cwqNRzGXnhtU4OlLU
hFRJxH8B7ckxPaMtmjXPCkwYC16UR5WtF4h0B9Tx5b3KfqDLjBMMsK2v9QHGWS1u
eIAFoeAH9vdk3VzCnM0THMRo27ccKhHMajyyEeKxXUR8ib0VMtWznEYftEeQXxzO
i7uDS8KxcdqPNxFxA9XeKxKlIRpITgva0LNIoVLuREeYCu74nyKPbJO/+eS6sEmy
VTkCYeKx6wbc66C4OVpv+gv13z+NtGamOqPJFJ+Ahp97YwMvkJBdv4T9L1+cAOK/
wDSaI1uxSjM2J9nveEslLcacnQpWXG1URiIcaYnjrJtyaZ+tPC1Y1y2A3y3Lm0t0
Br1OFV3if6SVydqSP95oD70VJbfdgkT6w3cMVlrGM7PiVx+UAdzm7+Ln5QIohZIO
NeDIiuVzpxfBnHM6MkOUhBKBnqJm9MfLeOFQ6C3tGgwkbPymfk1h22nDQBe6t60+
oTjpBrRBYNRaqN5ic94KO58vEuujCo9q9pYdIt2JcgRGf2cMdi7hKkPJCmbW+PDG
4HN5e31ViDo6OD6oPAQNqIq+6JqJv11T50MBfk6P5RuXdyQPyVfCY2QX+STolaTn
BwNzvHU/n8RuE9K7RZu3Uav1X0RqD3Zb0LtfpIhDrcGCa+QLoSKWkNO/u4SDjHq3
ET0h5nYeHTd1bUkI4KlMf1J1BXbz2oTb5WeSpXytigPY3qbEnHxY3WnMU9dgsDFc
ijbPRlzSW9bW1pTj2TCPmBdEyfab3X97hpcuV3wGeSRbO8RltmaV4HgwCUq4+UnQ
SyZRRm09mSextEZn583QxZsry3M3l5nalP+yjlKTmWLytJFcSfh0mza4ZhnXrx2d
3QWsT7WzCOTtxGKLAvl4EbCySPWpGz7zDlt88Uq4i2tS4nIp5h5wwcXRuRtGHZV2
/2d4jL5/Pb2h50FG0ymZhDKjPuPbp58MsDwEtE4B3OaeWSAZBU51SFZiT0RLfgXN
Nms5ZwlgvQCMc/spz6LGVX32shbZrfN7Rt78+3ZzRhWJVlsfTphO8d7K1sfKARfk
v9hIDbytPgY/Wrnek9CnGHNQwZcWPLAVhH69MkPW1drLvDZE7SVC2IlArpfYwyc5
ppAafCE7y/Wz0tRhUPDb9uirDKqBYF1zWY3cfPTfT9H07W/7HtWVq8rqGbtUxcyA
yRKI0fMKh/y0inHR2SFmHwL2qIZT4J11rkiSP73ruw/rTqXhdA6jufrgBYqnAbuu
duzWUdXIeq/oFPusQytZlkmfr/aZC6G3EPyq1CgS1mzIDXM3RJTmpE3tRP42h0hn
CPyFOHzE1gEIaWCXeuNmSvnh+XyKmxeWkQ0dzSw5E2MU8OXW1aKpV+QudrtVSpMF
aCghUf7Q8Mhu1RKEBXtd5gSTp7CSlBaxBDG4FKIl89wkgnFl3KDGm58ETCXpQucg
gnW+0DaAEDkpc0qqfjn38waqyyOAUJEylPXoNpxJei8ymd2Nu6PirZdOYL2b97Qf
NElqjuZJLOSZC25Vr4K0wbTdOaiylQT4UuIEmoLTE3dEAhB9qCbyH2LPnEbTXSVZ
EfFLjUUIsnFjdxn0McdTFm4kmudMbrFn+8YSMe/I/l2Iaac1qe1t8h7Y+tQZM1jJ
6wkSRawVM70KX2yEjVaLX0QhlOAVm+nM8N5PY5sUnDolF4J/7RaP2PU9WEoJWEGn
Z8/Qwlm0fcZcdI7lTOQZPAZinZv26fC11OJVNjIKh61rfKspBjSlyFApxmlHfg/5
oLQor85qqdKndEyFv0TViuHt9D/7qXnKUc+yYYo918a3MSeLVaqzTR3YMdHi+G6g
lxQA1UkOUL2K+/m1gFKs9DcZGMQtpfU5MphbvjQgW+/3vGbG9TqCT3i3T21Wbzlv
59iD7ZwLJdKCi2JVKVtViaXMrh1ayM+CZ6+718W747xud7Hr4N4AawrbtnghTWM6
2v1CkNOFBUE/VP6+DE0x0qncqSDsfV2MFhDive9ZKJdbGTgmeOxcd66BerjD76od
LqKkzbNzhs271MN7VEG/CiOuQSb4Uftc2+Hrb62Mq7arnZ9ZnmTDZI26cfTbG2Xm
xjc2125q8MdVkZiBNvnrozjqY2k4sqYH5G+LCiUX4WYztFOyVZRHUgqir6Qg2AuX
cXd699mqhkn+QFiTBLiNkT46+anyBObnSl5TLYw7mTdOcHAxRwLACD4KrmsE+eij
yR3vozHt7AvbMONDyCqkp1OhRLjyvrjeNWIxpxb4fW7yxSIhbE+9MqQoHREXlvUs
qIKNJ06I6tXknblm4F7QBrv05yDG+e2r3bxxfHzvC1GURO7vsP9HR1W++4XtQNhf
Lj2336MnZCgOBiJWdkwrtTxf20VWDAcOzFTvn6Mmlbem/4AgaUwU6M7y13IsmZY1
hxS3JguWRAUopFtxh8Hbq3gUb+TZFpCOEMCX8GF8NNf9N/NOf8/O4/c5WYrIv/NW
/9zHb5l2Qk5qcKIKmZt3xGxfybW1+IbSg3blnR+5NK74nW36uKXVf08oGCHIX4H8
XfGQWmmH6nx5xmEPu3guHNnCQOexWdq9cq38nYle8cB4/ND1OaxOlXWvgjKQ+QO9
sdne4avyT99e/TxPO1b49HeAh0VmNydqhh91wUX18HCVtWWIJ8L2qzKPmprWORFV
UsZ5ou0OP+i4htZ1n7DMzn2uq4gjOo8kXfHO/H5uBS3cNnOS1Cj2kjwaQheLg/LJ
9rW0o2EBpfuTUJlQXF+nDVptmyFYbh0lU4x4QiKy0i+0l5XYb/pmxaX9WB1Zt5sJ
HeyxZ3LrndXC7GghY/hyO8StyDSTiigtz3jo3dGfpCnETG+BQXHn3NHWrzvFFbWP
YuzjVglaFVXINoS0ZaTQ22V60nmA53NLCKvumqcZj1Mjkjoondx9mnqpFkJ7O7+n
WPb7nlhDE/o4uZsVUai0bX22P0AXwps9QeiQ29ijMhnbEUwWqs2POqb0VTcMI6DC
ysF8zjxe6RaDLL4jfNE+Y+rasrdVN1qoAh7x7T7d1ugyeB7yZVc+/Hf7TT54obex
uO7fXNBBGEx46LpS2n0GmpV8q84AXt0gKuDmWCsXiW1jiddwW868x9q2XqgnWwEh
ojz3/G/C7rIpztgf1SZzWR49wJBrL3VhWNjqAgLyLma14XCwGbQnpWHdoMWkBDoO
DN514mjvXa+4kgq06/fRgO6qa84UMmNCJ/zhpXh6YxPBj/4ojnkE5PkcS7RPwn1w
>>>>>>> main
`protect end_protected