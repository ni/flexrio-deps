`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 41760 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRmObns8czsvRiDtLMy5tgPqPJJUfbqxHLHroaSda7mK9
qS2YERM0dNRPt5o7iFWWN9VTn2MFCBH6BQgZJQ7GCNvM8AOb+gUiDbr1uk+GeFH7
qTERxzRPOgTZRc63tu5+m0+jqjZUmrybHTTaK2p8MCXGFj5rHjuJKSoPWDGhEIA2
sOBYFqufK74HmtkNYOTve0dWypexw7fm96KfzX748W5P73Y/GHRSncU7NAYkRchL
Kh3HdZu3bgwCUH8PbE6ljN8V2BlkgDKWNc2HWqEls/CbEl/J2LxrfVMDmOQNyaEp
+RlEt46qU4Xj7+kozGfXK6J8b4gKitKkgumh7XSxrx1n9+JHSESL0y5Wfic+9cYR
UzvSIUo1/zgp4C0swCVg57DtEVzcKMQQKcyPAJ5jue/8O0M/zjTbcA9VFi4cfAoP
fJsKqewchl6zAuB2HlAszEXDYxLtXOrrCapo0f7y8Uad321dE38TklTqJQjZzH28
4WOOkRMBtQgBHpOXilsjqFKb9NnQwYNuBm7WipiwiMBQh4w6ZZpZbnZgBRQuO8Ed
UXsbA5dvafX4AwPqyN4E1Cu8QjFrygHsoOireVRDx+2+IULXNnYOZ0hM8ZBJW4vI
I83t0RDJOgNMaaJqupEqApfhAE7uVMggbe3/hYC7ZV9i6uf6Wl3H+EJumvtLF4Lv
jA60qP71Mo69CR7PUFp7xJCmRkSR/WhRYK6VpwEBkTgbtdOu4N2sXpkemjB3gTdl
3JpIn6ZuU7sJXYRM/Mbt+HxgVusy8+5jegoxXT4Twb8ySBGBjEJUDLcY13/tr4ka
xQvVuId9YBURDqfA+u0E5toMucvaFAmv3aD0W7PMnwM8U3im+KSw5novGWWxH8aR
MphecSgYSQZHCBkW6mIDmCvR0tZ35UMy1R2yQbO+CCZEr9Kf+qolQhSSOYrZ6URw
oDo4nW3Xnc8nl7gtw7MwoYOicN+bte30uDiBvCxq+S09OenQLJ627JRiEnzz8A5i
JjeQfZVVrZQa6MJYOHa4Sx9hpdPRZ17/u+SF0ZSLyZsKwh07H9MMpPEyj9sbX/on
Ybb01uVn3UbVwbP3wIax8pYCjxLOps0XVlTgBr63loLiBwYk3vQ7taYcaux9Mwmp
Hv3V2MYiExsB1Qh4luYvFFBIW9Ks8Zcq/6fnld9lkKYeGkYmOedY/L1l1ZUO+TEo
I53dE7eGQn/JpskIUgtyW7ugjd3yO8EAd/9F9RYXaKsnNOphCNQjz0hEfm+HDaux
bcEjyvrcSVE16a3RHnL6D2LDECK9JV4fnPXgl3T+XOuNNwSCcUA9Ja1Zff08QhbW
sx0kIwINaKdlJyVe+P80PSxX3Q7D4x64pb9ngBR4wWIrW1uWbrk6+PpGkujQ0E7r
n3BAYomEonTy/2MQjSqyFpzLS838/Zm/Of1XZEd+5gXj1QrqKDfgBpaQbUbC1GDu
alXVGEGPNhqsuBHyED6425ZDRrdI3yQXt6B8GPCdCvFW//GEERRSNGyDR8YQUpeK
ZCEwcsqa0SLXytU2BWbFUHBSzyNEQQChyRyuSngKZePvxLjvOT6xka1heEKcGM4Z
pXk6tJ2czBINJSDO5Qg+20r52FnMHSHrBVbq89raXvNHcrHoD46NEUvBl0OMgEzQ
olu6jpiZX/JqX9FzLOPhdVGJ2aHH0hSLEUZ7vYBDTEA18w2DOAoCbK+1OZCJ0Nj/
M9ktIjgaVaAvSjbySexuOSv1jnDljJzjOkm0vdSWDL+96NwMIelZH3j+wA2vktxD
wzDJfK/xKzJR5oHLauwCJ2jrnZrN5Sd0XmAYplJLjCk2QvmK4Y9h+IIHMhaxg0n6
w96oMpmvuGsJm3/k+lEuLY5+m1j8cElyaJokL16PldLjatGUc3auvmMIgB9CCrat
y6Xpudp2nHnJANWLxapZsA8+/h/jQbM2KjaSPBwN4dwcCruToKSag4MblTKLaSVZ
PRhERoN2+MLWEPrAf32qm4eZi70PWhJfC+jJp4oTsVaoaXlaaTbq/eEpzqPd6YzU
FmNO6VW6WnlBlbWBEbHdN20r0CdaNHiOIxNr/mDPmT5QYq3Vz4apHh1ffIYBOkkl
2hCxTPqcogMi2gY/1Rgg7ymwU276FveigyH1oCzcuz4U5Gjvn3qTPogelhiQWQxD
Acj4KeUZaI5aOADVZzQoSyAEW98iniH29EPikwLUDFPIeOpFOayjltFGhCW2M1nH
Jg/UnnIXPjs6ELI++C2FevJx8EJRkdNaFl73nIyFVKbXlSAWRWzdlKXS+0tUO8wl
pCGpnWa8crSrIEM1RjZVqBP+WSqoI4gHimt1PTLJPV1MuwZUyX68CmtLB5rttvzZ
cT4uyTThJtWu1SuEdi0bbFUzzvrUInSnd+8OUZ6xYl2cBHb1Z6o8K7v22Zp9srZq
FvFTIyu6s5hftoCUxDINFFtP+whD63ru98eqS8QnaXB5BJ1t0u9nTgw/JIQDeXLE
LDTvjLna+A2RsVntxptvGhUvKan9MVZlK3KfxOLsdDWyGpgIAiZgMal5qC29Ms5K
q4R2X5Q9WlvU3fua+LT4jyLDNyu5xCZ6EqkmCXXHTn3gq1iH9fc8lX5e0nZuho1h
yLMxxEGoX6Q0Capzo2VE9FPWZEH9zurnTSG0Y6wGEJpF7CHkbrdpqXKGEnOMzW7+
VPID/8cnFGOGffEqtbU8YY5d3SH18YCxOIv5QK2cstwHQKXbG2VovJNbPfPyol2G
3l5cvI/ZBU8Mf9SPMb6K7LwFjp60MpChAERYHu2dxrCVgDb46fUsastoaxe+ZhkU
XC6txDZ31G3/9t5+h3UV4tSdXEtsIybSImS7zTw6b7FZxWdq7FUZj6S2cJMZJzlH
n4URp0jd2OXrYlr0RQujwLKSw16RN7C3vR2sRYsTcdw8WsV7LfRiWdP6QjGSbUJj
AJu2KEZVHUL81bIFftzSWq0Sey+v1DoEvv3sJ8O3IwPkZjW1I7VSB06KaJW5s7EB
aYkMnooEuujYw3uGqNwnH1Xpsq7O6N8czPherNgWZCr0oo7J9h28yY+pQVBImDPf
fRvRfPktzgmypRQ65HLN1XVrgIxrsFbfLLuPqfmqboyUJ5Etq/c5CPhAeqDssKth
eW3sdhvZJmkSXqQ3yZAgz+gfEKbRPTWSanYckmXb8X44nDmBxT8zxhlWndpF8RzD
MHsGO8tTTklsAvHkqAJ6LQcvBV349xuuvDoH24/cnqnbdsgM7GM8nYuDoJrZ2/TZ
4MrzQORV9FbLcc+YBSCMW9m917bCWrCVqAbXANgv+/aoP6JU/nahgdo7HnidFFi9
yO0+PFNJEOXlmOXMpt10oxl8FbzjuBM7oq6L4y3wFzrCrPou15vP3vW0G0BYmtir
b+2LhQ+y2GkWmzGjlZi3J992tvlS8bSszkFZaG2jRl7qQtTvqlZ3EL5jx92O/1xK
87Jrqb/AB0bG04eWiHWTjUUKXTb3+4TJxactOtuidPfzZKC1sljShqTL6X2F7+/e
RkNkTs3BLf9RnsqHI84V7UbttO3lq4uarPAAqQqKb6gs6PGpr3/Usj5O2TWxOMEE
mDNd+2M/oFf49y8jwHHvrYQKucyiaVgudqrqa6tS4Hihk+2oFQE5hp6XNKRcwOt3
GlSIsiJ0yCbo+trbBLXh7k9nwy3nKJX1It/9GagNqbnFifq2bpjxct5xEcWiEBiR
xn3AMae6fwWRrh3PmnlCGOdQWWQFh3vpAphUddq4jy9Yy5kSxslSZsyL4arq2VAV
cCiSzOW9hJtLFWZjtOk3YCaLr5rWlBsuD+6ImmIQKjN1IKyBQLH3Uj7VPoaYO9qo
Uv3nENvk2B1aqT/xYmCQJ5j9eJfXm3q3jgWMFpn4tGVIxA1bwGCdZZ2yQHWO8Qb7
uuHUrajGU/O6aiF2VmOOAp0zwtRagPzq/JyQAFAsROteC0cVAaf069l+sT093EHF
pqN4/JyS7xrQQ7HAb1htpc5raqR/Z0WPuuqxJOQeV/ZqhULAYE4fKTFaFmCk97CJ
w2CeFp1bWMWcMmPp8G2tpTrf1tzk4baIkWCZlFk4U0iHllqCZhcA2CoMl1YQmx45
WEVVWQ6aCmPDke2545EsPWZLW8l82fsphG51IRSYjQFfmmIHRQyImVI0UaUCBb3x
i3chA/l0rVqfdUKJAcAVaG1bI6jPKIU54w8Hi21DfuViDIwJyupsq0LlyG/K6+AQ
dz7j4UtzG8CjcuexsghyuezAKXeBNDMVmDFTDqTIlY0XixG0YucBNjMki3MJni0Z
cJn9rtdlDqOY4heHGfMYnnNBeqS6wR6dC8Gd7y8hgyaKW7EO7/853nI7DRV44FlC
oXSQCYAfsMV4PryECmR7Xh/Ae4jOOCy5b7UnOrnv7WeYfkXKNbgfIlIhegKfDa9R
hRHTnE7XznRgnHT3i8iVpic7xrM67sfxIGoCkFu0fTA2+PaTl3WLQBH1t60ah5bJ
sb2JiLFUpWwoebWQRB3VkXr861hOeZy77moD6VH4hBA7ly5AcRmTtLHeb52WmA0d
7f8ZV2uNeYlmSe6dmGmPi6z8aag6bEwbOZ8gGgOtv2GlohUzUfXM8QZgGZ4OYTKE
K5zAdEKjaIlBUol8DGc6n7+84thGwCJ1z4cAhdYOvpI6BKRbTB1ZIlB0bVzy3Iq2
t+JWDvI3kfCwXR7PatD6f7MQoyJOfftVD6k2g0Oj3cxeu9wQ9bPzZFh7CrnSXMNI
5tk2C9/WPoYMotamVtEL4oosqt3ntaxw8BJGiPMUOxPLTs6fEeS1p85aCsabm2vn
T4s/HDRmTsNnwOO3O4eYE9zRNfodGTm/wsPtG54f02Mvmx72Rn90uZjNA4p0lwKj
MZrtnBLAXLb8LYCKzD2qnS4uDHnkvKKYb7X0K8XdLD7OMBJ1HhGbm7aWEwAarFzQ
7tIbz150SoMwfR6hPLGW074JmYTkKdTJle+xbJrAQs2wpHzbTCMjU9N3HJPHA33y
TACxWFGqwH3D0fvuJErCe7bGNafqu5V9NWdwY+YcDGViMhgMMyP6rvGclYtmJCjs
Gee0PztgkolBk0Xt/WXoFSN2v5e2h3O7+GurgZJw0Eqe3P6TSilkoB13NUvrPVbo
uzrQGTQMXb7LYoCuGiRRRRR8YNSKK7oUCI4RfUSJQsqwkI3/fm1mLmBxAzq6H+mI
y9WU2K14SBenn/3/Z+hEhDhGxxY37/Xa2b/1uhnFuUPFwfqCRxjOloaFsf70QmUl
pIhpUFPx+yxLi1KQjA7yA2W60RPJ7Pmy4swmOhEeUMd7n3HFNsN9ZgHALvjS5fo8
WKeXF4PXiM0iccOPJabpdZJau3lTcn9pziiv70zL3uX5iPbrAI6BuFASZfzsSqXg
6bQ1XDlZqCszVz85kLoq16PGfftyXkscZf6/C6xaGLVGMTLt4r0Nph8o76RJ6r4J
xpxoSl+/uMAOMIXy7+DwiOLStWGPz2JdsYcULND+uz8kOmHM74RormCZUXRkQ0ML
KG8WsQVpjH2Z8tyxeszECeDKMJyGV1Q7Nc/DyATHu7oWwZ2NCl7DZvRZnPUdXtar
O3tk5WdUuBMs5KUtaEmU5mKn312NJDj3ZsAmTzvKc8J8VRxpm7MNAiUV7yGQf3zW
w67k8Vt5LISed9Ydvx8LFzvClFtGC6d+qaQ52hCfd2OAxAwmfUe6qCnXbgV7blyn
83bU3sycWfdkK2XiWc9lc8hCsjTmipuMurNfCwClYyFxfl27xh3N8T+9dcUDcmP/
xjWNXraVFKEbQr6xEqfcbYMwHq3LeR7uZwcYhJbjX+KOU//Lx9MhZsmA++Y6ZC4u
mLBTopyQYFBsAQntJ40Vg1llsfEeZB3kIZravms7KHPjLK2nxA/TFzQ8cZmW1/4s
w6hYvWdfBHjLVGnEg/RVJTqBxx8Wuu5BNo+o37qMUNW7ndmeN6n4iFL9AtNcVHZ2
vEIYOGpULCjfqK6+OWXP3pyaG4hmi1eJqHeSwnKs6AaMQO2TcipyJPNGJH994BAu
fQK0tbystIRzMkN2+3sO38wJkYDo2/oxoy6Dy3Jwa/8Inmyd72ymxdv50/cHPP2F
Dle7Qxo9p7pnSzjSA4R1IRMlsREZ5HlGSjOCjOTFX/linqd75IaMy5Dk8f7i+asG
iZo8StydlhWB0nCtoqvkGYzaNblYW8khlzs0wZTHHhnaoNcS3tVvmEH+8dGMy3NN
6Xh7qJ/U7moSdWD6WTov280wQC5bTtpbnBA+OTb6O8xh81bg574yxqYwCd+BCwo7
abI3tqS9I6waETJMBp5w4yqSPKATQNKouVr85ujCRhtvWGN4pBZYPNd7JPrtRgzc
9Idb0j22Wrvmid7Q8m16KDF4N8cEnxorhCrceq0FHsBS+o2HRzj8lYo4mSQdYp70
y3B1llB9TtU0WZp3K7gnyIoahwCGAPJozcuW5WDN6WdNpDXXcr9Q1PsFM00pDECZ
ojY8XtDIgPjyqMeYz3brghJb9cy2fl1PWzbS0Q9V2Hn9Jvyktz6WmBkO9LBQWueu
uwcQlXDmaqKXEtGwYH7Q9Cb3Dl0rWppdQgXRtQZBe96qeenFs7xeF3wupKZa9XFT
NBAJxg2O1BAvkR9q1pjX6VHs+Dq1sp5uW2FRfgHkJkxI6BO0XA6PIvMVLLVVi/lS
w00ULcg/Y8KTzxVi5MniRPGpzWR6jlGYMcIkuEP1aPWgxDkNxFTozPg+E7k/Fw10
gxR9EeaWJm8mz6lkCFkIMx/n+MhVmMhr9iMUHrlscX0uFpTwakuoEOWzQ3o4dY9t
jDnM0WZ+6O8ICXrbzMlpARXu0L5gSrcsDTbghPw8kCDeQgPh3wtX8t7wvPAby+8F
Tt1AJjvEmArVCc1m7MK9bX7+U7sOzYezIOYXAsWjl4WQCMcFqbJH4qyrmSUN+8Dw
ClaSgcoFItTf2KLm1MPysZRBdFbZ7IbVIRdZ9iZ7+PyKqQe/J+1eH2bcJjGWCZ/O
OSd2gHKTaaNJm4TbGhoucwsyYCfYmBiq4rHOEFxlkx6FyELiqPu0JcgQlbVWjUOj
oy55VJxsq+RvWHhLfnuHBIWqOyEXp37tSJsgq/8NEoPmQCZhm8Vm3tBbQi1eBf0u
Zc7Odim4KKf2TGBWbwynvRHbk7WDVQMxEJljHP5jDhI6wwtDUK/8bGo3K34E+FAT
lqLM8H1kJ/frkyCBdKXpXFrbS7xpl17QkKBufoAM5mtYhAemJbb1h9kfCUtfBGwO
hMdFiwpLcO+GONiXMR/F2Ac4SCHpPE6pDpYrDAIa+8so3iLLTgLlEpzWjf21NDlq
EMaRySiCztVEGwcyklVSimTSRqPDx/ZwNkhJ034EjE/+nwE0GBKNcCLa/ZY8BhJj
P4v3mnsMO0fEjXhZLe1+ByJLRJBbIdHS4eoSEWMQ9v55HV/H/DhscCClrWuiEBko
KEp22meVqKLqU75EclNIPwtQ0RVe3RThYyzzcv7cz2tyQzY4OFJwwCQYBLD6eoRr
m2UIXoFamWWUIDoojPQ/vodoBVS/wNeukyP9SsNNaa/CJxl9rvO1qFrUrFSAkQGE
b2O1P2BoKRZlvPVohe9XxqEr3fzJOMx5oowJg1QKlIxa35Ymv1sT8WLTDhJmm6s6
qszRiNR17e3gIOOpKaPIGGUwKeu2zKhoT+tiTDMK2HXET4tAkucQGS4z6304P5Qm
sMsfiwjucjao3+3PDo6YfwCN2K6a7ugNv70SALBSyr9wv2PSqk//gsUewnr4hUbW
99VaajHBwxhzWurnY9bxLT1tUuQr7Rfk8e0QkgNYw1/uEziJsyR77NOYi+G2BHth
2fxuUlJSl7S1K+NDcZWRbmvm+wXcLT+UOf/TO3OmMBoq5MzNYHM3J1T0c/xB32Un
MRhPWA+5cIiqf4UHw8bjLe1UUVNGAvy3uYqr7MA7dH7+6pmBuBs+RpL6dlAgkUdd
kH8kNYd2n5A51XeDNa7SRkjZbOj4Gt2xE15Fpnf9A+e80x3Fdnwo4bNPDUHSzKxJ
4e9NxSIvKX5DJsnjU8ug1ZGfUvCIrRYu4WPFYJx+Rgpyf5GGeUJ0344EmSzDjVsi
lBgRD1OkgfTzSQ4MZRnsysRBlwnLVLsUGLHP2IB0uOzx3dvBECjpHGg5SEU6tuTX
Ugxa0y9ZN/40lThipn/aWfCQyyIRMpDhHu6aDHjGDK9gY5O/QcxX3ZeL9MDYp1ug
XDfQdaXVFGAEOHMxsG1CDBvUi/MM421HFYVD9RgduvUeH3lb99vdq/QghZkfo+Ut
I9WBF6Rd7Sa+jyn870S/1FHz7PRTynnTLrVwkFJrYL5w9Ca/+9ZV5YSnrkJ2UNA4
bCIt9tWSXFL92kbRXCweT5C6n+YBq+3x+Pe/0PZTZjctJb8NZDANGF7UsM3MJWvu
ito/FZ6yXkSXdwMr+QPvXLo68M2T9OPveZ3Ybbad+dp+c7x5XfoG2xnclFHCxsm4
OeSOQAu4hj8zu9n2JakltrCAkqbMrpOs8QL5naWxqIjrT8w8BItEr7eldbgfxWtP
6+oZ0UfscxfbeIs1tTXSpXmgIypWwfqGHpJXOWseYDRfZV+xxXJ0Pw2PnNGJ2f+6
FHSW8DpClja/qUM9N6rQChQZoR1EMi2oz570Wf2gk6dqwm8Q2OuKBAF+tW7MyfJM
JEayrXRbkcAlIslo3LoMu3okJQKP6bcB9Mg30NtKN04TYiVQe9nvGN48aYlOOlyQ
+sVN3Uu6edHIgKnP46mFlGmYBzX1UZR5K2UWyFulGH0O12RvWLbGrKnZR5oeUAlw
1oC7CUTBmvMK4UkC/nYfEZzB/Xx/M28ibinsDQXfTaoyrzXAYOtIrOp9lzFoRxty
oKGfwBvTmTaHhTgI4w3G/Mq32+/6T0FHkX6N046cTSmVKhWVMumLrilT9tiIQRk3
kGQVFp7p6qvfFm+Wn6B2fLywghTJ2YPqTdZjFn1q1W0QxKOFtZHmQXrmEgSdcWA0
NFgfixA9crhCmZg09VjZzoXgVjCRcq3OXr6Gv2x5cPBiRcEPpGiO4RUHASXOYGi2
T7VaRMjMffbsE1QhtNxLn2Fgv83UnoTCEJNrtSrjuUcQtvVhySnped8YDe0x3rSa
Pd1zBChGnb8Z9LeVngtjWrqWK5dAMdtITqHvWbfVkr7+ez6PU6qfKDpSW+uNOKPn
UQbDbdzmjEK9C9dbTWmMRF5aKE0Y/DzNYQBOb/SzdHlaO7m2m5AgJzMmpFOIiJev
Eq4/YTvfmzJCfDpvI9B1gQtjTmylodRh7PVjaRnTY4c9D+vyKKOSlXWtA8hJvByt
PnbPXZ5MtlJKVz87furRtruFD0zpbLR1Ft258v0hj2uCVmup21LgdRdMuyA+DVkX
BRHAjm5BX4YN3gy22xCm1NCoepOU31WMUh7U61kP/kvIij40zo4Zx2X96bcE/uK3
MIdQrZtMQX5RHgVEXaHQmTas30Pkg3dd2utIAotd7IkSOLUcLDUnx/Sq5nkbYD0M
ytqE/gpsgfXFVzF4DbdlaagUsrOrCrbyMgTDAKQqO46ipK6kGbksbL2GHOozNTqK
gYBHGfowqO34V5UUtrcMT60614zoqxxrEobzykllRw8/GV2f8hOxQWLy2y5sdP49
1WFpItvA0QEIIk7dr1NdPutg0wjY++5+2RS4OG2S/pbzZzBkI9hEUZtu8XVmLH83
M1ah9hWVHuCbYoinfVbt5O9JowcXz2y0JAvDeWtZSWZlNTPeki6yssPdpJs2NkuP
9Bz+Sarw/EmIb/7tBJjUA9jBeZrBLdGUaR1BRzcZBR1AAdSBdTsX7w5f71kgBJoK
HNlVfPMT7fG+IFTdZe79KkGwpQmitpnttxrfYI/HLBK4/y5tittrVR1kwn4H/Vey
VNBKF6sPYDeSteH/gXaEx5ryip7gTtFwwB+F1jQkQm8NZKAIZKXuH84Pn972MlUw
LkJAhK20Qj4uJ+3J46Uz0KUtvHiLVbPL+0kktEvFzo+7oCOVUMt5UvPjt6+r+Yde
hGWbKUpBRQPqQ4rx9C4b8sSFTuMEpa1XkK8GpW5FDE00gsizbGRtJYMcsbWoCLmB
5V17y390B1H/IO4XydFa8MS7nhkPMd410Cq0v5Y0Sek073dlWnpiAPyxe2tfwP81
ttqehRiihD+xzUACq+Ki8DET1Wk7CwrWibT8zkR9Pe9/xeAt935l38xRtwiR6k2K
tv1C4ywxKO6gUpJYH0FSt6ECC8qNYNVGSSdAJAvB7mnrKl85Khib9ZEWYuJyMTe/
1yCUmsAoIBF0fEPHLEcjWgsp7ZFO5wc4bnodXf1/nRkYne/FiiuBRde0GBzm26pe
vboR9h9iPR6iKSRB/kKQP8TT3uOX/wJ2XATfEQCkqTNgovqKpZGZbgJay0Guq5oX
S/5XS2Xfgxi3Gp2ko2MadADC8w/e7fZC8WLs6GbbldZaYvGM9LFQKr2VurEhO4LO
eQ/mTWu0QGwO8MFTW26Xcorj5e5LeRL2krHnZwpEnD0R0dCv7SxR5nVbxIJUeasT
wmjYYhU+3TSNWczWmJ+ZXELCxeMHFrylzXuMT/N65sinpDX/SU0NIRcCtnU5e5xC
1ZEFfBeRToSlVGl3uH4zXf5jmhTd9PpYh0GLpwVoWYHCefzZmp9boavczZ8MpTSE
oKR20V4i2AlDFC58/PV8KRNxhSa55/nVN5KIZMjNNA3bGRdL0P5IyMLA0KnAkxcH
uu8KjBfc6KhqqzR5adUcdFFLpEmJ6EhOMWSXzGfF/+1FZPs8liKLVyaXx7pzH2Xs
m7xlTxTU9Khn+xL21VGTD45RO6E16JCgaJVpIOjHLAZp4ElOg7c3LdRekX8aIo1e
V1ABN3hbxvpxWReY8rH4IjfEf68uSKIdhH03gA0EH4TfQQBf/vtnIbFgS2w40xZQ
+PTcPlx72qyRm5IfuVdNqBjQe9uhXRSymNwxl0mgdMs9kSHmCbMWzxEFhaPAMh+s
RmhURLJWCPh7UQWt6lIhJWGfoc+llHVE3i9Z0WGQzA15x0urguLlE1u8tsr0xdJd
+3573aOohI5w9P1PomLiYh010AONJ/pmkSeauW23ApyGWZ3ATBIL8uwb3jzasrux
DiwqMcQfewH3wkoo5QG2cUwVZivOXeUwPCy2kXzaFDagrZW1beXWBzH9lmM54n3t
XLxTkNxz8aiWbXw4SqG5OZ54ukaEQ+r0vn5CzcAV18GthkqsH99rstp0cVnVpIAx
SWSvs/I92GCzRnA+l5ct72pC2+xzpgdQvuJQo7kJnFidueX3n5xx0lPn8h2OhHya
5iAPr+EcaCzAK3WkQO4Z7vtPjQz+38iFWNTHQiz75pciXgCAmSuCyxkh9vRSmHIt
Np9neTm77S8QhKcBiZdBLqBytpTZbfSMDeJFSV7eqz8hjtPKBi0nk/bAjb0tKFcs
1hKEzzIGuKkdGpGcDxL41tCglE+82MKmLVkCzgocFo/QVH1Zo73pQFQGVlBX+XMA
4YM3UCKDPZDrCA8GQ8Razis+LcVzH+mKI2Vz4Rc39gViADzD2W5OhY8b3nhCnlIi
PTSOBcmFsRF1LtYVm/ETCBssH5Xck3BQhNgFtZYX77fm6HXhRorsdM00wj5mutRQ
5+lDQw6bxAED7MuDLZ+4fDQlRkRYjDLYR94aYBJ+x4jeOlAxfQPnS4+0Ap7C0SVX
ivmMP9XiwssKMceLshyRJgegg8Wwdtk/Dw6X/oZEdqSH7VZCUisdng3QRxFornB5
3YmJ5egNQeT5hwbbNAFoB0fHYLPpfH7M6yFZxG0TgTUfIfmzzQTJBzw7zuyNrwEX
dzbjTSYm9+AZpdtU/o0ifoB4WDJi9SQWZ7DvUCcMT3OIl5218RKgH5uoIRoxy0pa
h8kUTyuo5pl/4oq59jD8AIzYc6Qc4fUWKQRnj2EpwkdV8hNHRwhdal4veSsncRxX
VaIQJ5CODE8HRVs6OLMRkjEjV9QWYc89IFx9WBxpgnrGRaZeN7O8GI3hAvookc4b
vpp5X6eT3G/zPt8IEAh8V4WaK4UBQ2sUPWunNOQp916TPOlTI0UjOuOiEzPwwwY7
hsvRvVPV92vUuVIi2yEs+OEBKhN6uWMEtLvRS/anfGsMkQB6m6mA7yCAI38zEcip
ek25iH5jq7zH7sVRExbTaogWxmeWP8scAiAomNNs2XKE/7tVDpEmTPcGuealMi92
/ppfmd/coU0XjKZ58eHRWqq8+w3Ua+FLQB4zSEWNmV+G6GGz07tZHH+cOZMWfASP
tSoDqEGHL2W05oxadZSNSzlQjD5oZA1iJaxbxthWaZJk8/vcW2Rl2g6J8pkdxOJz
PxXOO6ZHwu74Nhbb4ncPJQ9BjiBRKMB7Xd/ppKowHUSAB9grg4U/BvEpjItEx1Rm
tD/jJiO+/GsAmWqYfjRstqS+27JsZdyeZ5FZDCV+6QOoU5OG+mcI3OP2y1Jh1b3H
ghGYdYhZqpW0tqyPZt6WlhtJLm82Q0XyQ0008rBjC1+snk/cDXeh26mZFG9svDXA
eM6Qz+8Q/MEJSG+EGAJT5VgsLCEmwWOFB4gCTeWV19lsRIkzTqPjUgFgdHmw1WTs
nTTUiIbmjUrwKl50pdvVprk17a6pSu4TK9A8p6jnv9TyrKg8b2+WIL4uGg27lsCa
nrv28K4MsRSrxwzRpmKPmun9GAdKYokJqCpGDzFJ0H0zvc9YHzvURCwMSeOki1ji
/8mOjKmkkW5CL7+iKOwbIW26BhwBOagIYSnybU+G92R0QCRwz9IYPbbT0CgPzB7D
rrFWtPH2A2NcLeoSbS6Hagrgen5VJznUCtQ7LjvFlXKMjGY6kLBtABJQJqh58Hev
WEbXODOADKuMnE70NhduA0ZyWXGhV/eVLrO/58yJ9LDykqunf4b47uBRAyC/S1B5
Zar0myiny0Z+ucChNEPE1TMShGvu7bSf4Mo/Zi2kt/6FHtxHh45Zk9rFvhGfTGuR
6Vv5+xvetRCd3dlUmbuh1Cjd9bBVS9yoilohEHOcfSXN3j6DScFZ5NNSFRq06w4K
cvQA/9o2YLQQ5dbUfdwkoUbhK3AusJur2m21JkpFNXEpJDr0gH7H79NkEHOgGq9N
isLKnPX3V+4FWkrqbRPkZCqE8rl7mbnD0G0eGx/0ekKHcxwyFThmADCSieVO05GI
UNaZBq7hc75hQH5n1wwikxbMe50dkidHQqNf7tzjBeez4p1rlrC5paeAt1VNWGNH
wKV0fbZ1JqOo39tfHnyW1WX9RerV9oVgPukVZqjF3rmDp9DgkeqjKWVH7zm20sq3
W0uG3veaXmpxMwKUHSfnT2ZgNsYWqd1W0L5Ogzbfel//Q3eNR8Kt8GnI5WUADwhB
JNWn8qI739mVGGFApp3Iiw+nUv5MT9c4JYVfHjrfAXGBDi9BGLeP1u5ctJgAl3XU
zWdiq4WXOuuqIcGnd2ebrYQovhY4QoaA5y21W7cWe+FcCNL8lVzY6unmSRMC8qQP
OEdG+/kcIimDVVhjhqX6owqht3EpalsQtX4AwnSL74NKFuAxrjN/pctaARY8hxco
2i69A38suP534nTsNSaJVwIDTo3bi7yPcKmyo0m8mycoDtxeGsFtfspaXfUpHw5n
cIv8BH/xVwrZOdSOSFc8C6sVNv1DJvwJvPaLHCtG2vyssDBLnapESybf0QOG6Lio
FkDXvl2+c9X6K+tQPA5Km4lRONzXpSVCHhwRLmi6hNywQPl+FjJclvdOXnSyCVzc
4eA2u6VcmpDHrAbUrK9pnJDNWrmhguEsXsKSutqhrvI1JnsnACK+JXJtKJCfEAiY
x0Am1eNPC9R3TrINHvPkkR1yEVQxsCDcqqzsd1ibcrgNqkY6zGGi5NDGZQzHgHZ8
LfIxvhELS175g+LGTQZAQ5Q1sfnuzGAjLEDQlBXGBr3NW6sCR35+3CkDWSUIUUFa
da2qZuIUvj1Nj+LXsQhR/XNQEWGekAsrts1jMEnb/0ezmWU89B0p68/oBdQnJIwK
gBHN9HbPCNdbenadl6tIMbS6a2cYW2cKd+nSmGs1T+3KZHvi+2CyDbjBHhv8/Jt1
9Ks6/T6qHvIjKAEMiYqDK9Vy8U1jWIFgKN7iJ44OuwB0/xj6ktH3ODpKoqLJUb85
qyiwVl1i31H7DAwXQdeJSx9Wx8a3fptWE+GWBvzGshbXbm7hHXqrp7PWpSm6SK8U
9eOCDXaFROIIUwMPL+fDEMrnF5nzEw1LO9sfALd3fLqFhMGNXW5fiv8iQHzNRenE
fsLg+wQyAR68MtCZqCD6C+xUwEgYIRYkiN4sHChJuwzg82qCQtBJJ5Y27jng5BlG
lhg8b52s6Nc+/7pGY3eNnS6cD0/Or9dCfhzayyQ+TPlTHouJWNJbc1eQJejBpwxX
lpDNpQJaNRc44hgctM1Ro4yfPCJV3y0/sK2ahkbmk/tx+Xsrxy+1OuXyUjtZCe3o
8XVZNLAvK/92CjScWhUixuDE9XZuEbR/zPG4RmLPx11d7ODBOEvKYFLIhiRhyDeB
lsVpbih7vIUwIgR02t6UPL46rmXjfoQ1S6FJQrNQBCzJLcZpNuBEtlPxViOX7VXj
IaP+vOn+SqxCbvbgeSnsocvn9sO9GcblEqmaVSfASiawmFswLF255mBHJqZ2YM3T
wE3Ty+ZZW+udblTphSJagwMoLt0ORuCmTyKsTiHHKuwTS+/Zxxgonqvz4GxLIDn2
q6qn5IF31TrhIUhNM7JMOBHTcFuXW9UxfGuWmCFykt7zp6BlkJvnpAhRW+rhPj/Y
DlnoiApA+QuVWE8HXXC8TWi3SpgRK76rKe/gJPYbnCVkjs7Z3E7EB+eH66yyMpKC
mefoDWFRQh9s9jCIuvr9MOHADcNKUv2rANpaBk9K/lAdJX7/58YKLxvxXAD9+zPl
Ikpt1431IdwMoAJMKfIseBg5ZuWIWc16O1T3d+hgOPVzST27P1AUHUvsMK4t0k5/
BnW3IzPxPjhLxkNTObZ1B9E4mNMvzsMa+gb3uLjy62LFRtuQWPPOoppl8zaebOGj
Ir1Q+Tlyau+XAL4O1Ae6LrhFynLfl90//yUXIRNf4CyXTbKO1U/sBY6DKAxrUolk
IgYAKZVshUJkVwcH1ZyEi+crVP/nPMqtIb2f+41vjxbWxE+Mp2r0Eb0MTs5nh/5O
tX+NCP2OlFbGJrBEG5E7BFjo9UvPH4OlW9Qv0JcoD6GcQlWiFQwsed3YpSHr8NGT
EVeY16V2gsc1D5WW9it2VE7Ng9r450VpLGD+/d8JSN2GMp6j0A0dHGKISyVLvKAN
c8iG0Ujb8WmdFa4HFoOt8s4XdXuatdEIQiiobX1/6PosEAy3Hxkmp91/VSpcq/vv
xSw9IDlH78uhTHZTGwFHZVeMdrDn2ZFBARl/gxylSFOBgdu8E4Eh/inSGqsyXW80
RlPzbKjl5YrjXPttiaTWKAYq0cP9oIj3pvN6WuLN3c2zbbgSXy7ObTw2fRcuKPR6
SdbhNXAIrB2bKI6wqAhBNbQD4FLW17pp9I4kBg8lAYFjfHfj5bvitILbtoBPRvw4
gOPuoxpBkY6hnBSSrliF9lzEgTMW+X0gte1d/51eswfGO4/PnvwGoRV2PVKrerdd
in2UmMUbO0BhtA3V6WeeDRMwGsoqYHT7eYKpU8x5CtOTXw1rwbN8zx4Icfe5XZwE
f2RwYzQUu1zz86K2ZIbTErX6azhEMc4rAo6FEc70bo/dhCV/utXhuCNG85+FYeVS
UDNBZNREMvDii684BGS5XYRjCxusiqX4mv+3X7nvd5bqXsi18dpPH1XavBw7UTch
jNVRkmZX9hGjXNwoLtFIePKbAihzsZFCmcKYU02BXWYce3kZgYba6pMWudnzOrNs
Sad370uf+gwVymD6zKdTE2nYMPfJBqNrnUwr1z7Af/CsM4IeiNukT3ZcnLpR66RQ
3FiQ8h1pWv48JOKy+QrylzjRUAcW69jtzwREOLCVIRUOXM4XMAk3J5bRmrSIC2yp
f/9k1oOQIPaAIqH/8Ib4iP0yW1GGyoPBNReOoylaPKBhfD0Dk3AFaO56OT9cJpwQ
4nJdWcLZnbF+1998ZG7Eh2S9mQmrYmypg3UbPr+ePtpfZSytvqRHNWZ7vmmsocko
AV2tXGBMmAqI4sbKcNhLUOQlZWoxqarkehoN4EBCMhFAU2zEhOBXZjHNYPwu04OT
Pd1fqbvShHp3Ce8AlkntaNMAs8Ok1vBbnSbBAUOuz+LcIiZrUzeIPaG/n572bGrz
DcW6gGK1wvlqFvWmKJyqR/0Q4PDnNGjjb5kOi9ukBgkuNSgQT9uX0CCk3LMMzHU3
SPN8doWjXp+8gY8IZooirkY4/MiDK6HkRJGYMQQwkWw9Iby0NI++CsCwTjg4lrz7
srtf9Blh4lNNRg0pHNrE692raFoX9QP9af6FOhocMn56VTBhfX5ykMkWwSmqNIUZ
Hmauqp0h544bZuDo/oWJGsM2W4tEU/Y7r7Pb/KHdfTr9q9zxFo+p8oKCW5mP0bZi
el2SwU/SVnWxImogJHLmAJGSzRYgOoLQv2IQPoxEFwgD1zx7VLpt4ylRtLLeuqJx
ru9DajewQw9av1r9utAG3i5IZVITpBFBl7wEMzXjfPz7MWqZPYlGz7Glnc5/D9pp
w/wPJZKsNOKJwnJtJXvkSYnQx6yjc0x5i0UP0fu/j39Y20CbNabe6mfVU49CvwhG
HcB6S8PoMoE7rOR8WxYFiiiRh1miLBAPhVtNkw6dQOqxIIHfPUXVGGhuigeJ78wv
MbClytx0OzrgSiJWeIxDtjtIPLQTLeFNFZDFmKtWowyzXwPiY7OmixX/f5Fxct/H
QZv0znSKlmPbaxa9fh/opWaRMrWdbRVAq+s2ChU101NrfnhIeeGnwWIdFWkup148
Imn8vYTp4N1FVL/xaIlQMqrjG2BVwvBfR7qmsieDI5r10Sf00+uMkyEdGyHETe7w
bGqLodRUJiK3zMU66kF0rkdxWY2HEB9NJRXWBmNo4VSgV6SPGrYlRIY3ZcxdcWhY
7/lM+8rzTYhFIw/kHJt5F4h+lihkTzrC98Mxrfm0nu8phfq5PijgdS72BW12+l1z
rcqVcXrW8vFlBnQkniIs9nhpzjvq6UUJBOO7VkKonT9khvEwg1OLXqct9+m/i64y
OrZ14A7JqZvhJ2m6MlRPVLx8XkgaaVzv5+BRPqEJMLNxDO+4Da9TchHJqNjSqaUg
KsiKt3Dnpd6nm5vA28Vq4zY6V//uJQGbJbZ1c2LHAtCqhwS6rpzlajWSStZZ6h2I
ifRdmTmNfg7BYb2R1Tr/9tw1xUj69yvoEj/K/fwxVh5Z6W3a7Yl2pSOV6uDMfO53
aYHMVM7+hL3qcFYNpZxrLNF/QK7OtGbOSbjuT0Wb5XoX/eJsYX9xRj3gI84mZGXd
Aev8BSLCqCDsBCTi74f37rZcCxrMFK5mhHNwWEeHV7pJ8iMt61Tx6fOK2lImkGB3
EIqvQ5M1jffn2R6st+2rLjIjrL3Tv7D3MO2PPn5s94DLknG2CCw0hlnUfeUnHn+o
a22JuAZIghE1v6ofmFHg2gvzLbMvrxI3SWoLoyincQnle/SwmPdOWo6ejTiJKyLa
fNwHMsdZ6G9MD6WrbhVMrcQXokPLdNTwescJ21SwNbNPOuZu886bkHWNiQskHJiV
kanRNZ1E6kJBvD+viBp6cQgK9fV5BJ7e4D/mDIiPEk/hnRifTaPf4wXtV+JTXb0P
oCT8N7NofWvzbmOJxo3jXASmd4RdnHv8ORbYL5kDuP0p6m23si1hEEziLxi6TItG
kWQTAafdQa+spBjlB2BJePvFTR1jPban9OnRbEGWDDkSl733uOOzJisADouEfDWF
5F8Vc4WQ7Dqr5/HWZe8EKrleod+2hWcwEViS2VUb/u/7mQHSgUpQbfyUNGEGj7a0
lqpsPBcJpqAc9Tu2aHHXL12QVQmwgPLO2kF3uPOeWZuBGL/Op6lbMY1DWK4BIRK2
9ujVpIxc2ZWsuHJUmzbdKNTrIh9jxtY5GW7M2T6BDcwoOF0sGnb+/WOIs2uMUdWD
2OFH10t5Qvfa2mL7sKkqIPPcGZoQMWYiyp6npv6EzPEvJr36IJiUFwDjPziYmags
DEoDa2QGUUT1ZTMXCK5MaGB8VEQ+9VyL4rtoKlDcs4fFus/p0BQqin72V2sk4KQ+
yAbkZu37uGxrmDuQQc/ClgTK3i4tPEvWzLJxu0gEnpSNp8vKo7PQV0Uhh/QJQ83/
l3kJVnqzzJAZHw4SmvPGkxl4putRrQ3HSK1p+uD6emsDGqvPql7VPclWI695RNBD
PdsteO/5mC59NJm1L6AUIpWfUuFMxiOS9w9aIXb7cpb4MfLLaacjjTtMNV6dwm70
oXU84OG7XbQA5PS9762a0zZiI3f9MvjAb4ZBNOSDFr9kYUc7gvRTI9zH6wO8kmSo
LmQIYygeVO2Hf9mEozI25cbgmdPNsam3SqN/zwryot5MvJBsqzq0EKf4tMSpRVd8
TXxx0vjCWsR0gbb4iBbzRELMIxulXnBDeN0OsAWGyMlgGcOC7VigiJfszMesIae4
FGSgaXSU85arVX866G3R0AxMd9XGqWBt282qtQXLAVIXvXTF6n/W5L7JZs8Xec3l
X6tjR5qdvkCAoxp/LSDcpgan0SDDjv1eYCk+K/uxhiU6Cfxx8hw8ouYZV3oxsAAU
bl/zkynDOOD+2Sb6sjdrPGOjqFU6qyUO75/0El5PbvybgaI5JDB8DrUoO/4WHOaP
N+ibGzUAn2OjcvG64Gf9GBSJ3qCjgFN/X3Yh4fG+l1pjZDAvf4q5oPb7AsDzX69e
eR8tA6Gj1l82FuJntYZCizNtZ2dq3H5/h1bYXooJBbpeijfpCX4JromTSdr664FF
L1PRe7w41uj6AH3kYCRy6rvM1p9lw7LBNOC0rCQiBh/wL0RgwWNPmf37dGsokQJm
aUGreu6GlBgZS8XXmW5CyXKfQMZWjvm3ntW/26F65dqftI3CQFxiiENphadodb9b
OFS+ATRxLPTZn3VcavrJAUMvqGqtyBPYPhDVQhMYenlLdVlenyS1krbMkDDKpcu2
QWzcOIGGJgi/+0JpwoRANoAi5FRIuj/36bKoRJSyB6rCvjSxMtOd4h7vtyxSQOgA
wrhapcbhahEBfO0BNgsGx/k+XNPIzcx36xU+SaIN/Cybttie+sZqKPh1jXGjCT4o
31Aova8n9X4VPq1AVZL1GjSyZ18D78UHhDT9gJ2CS1kPHH8jYvpsiA1/moyruRDI
qQPSMN/FbqZTMCkZoYza56pKpqQSGXlp0EvTfE6pzPHfUqOLknNRFBW4oQa2zdP/
RdgdeMZKjfs2LkkZWp4xTEhzZg4eXTaIdQjb3XOvMTEg8JVU0zaAcCqpIioemskd
NwJ/u1Sgl+tIavxT9rOOToQkKBnyGMn6Cl2N6/uq2V1L879IKb5piMqcKJegteQn
LkvWcQLBvQtnS6j+9dFl0c+P1d9AwU3crtNEQZQOBJudcdIB0VZEmHwaAwxd+qe0
4XBoph7GxWhc/ZrSuPvIuJHxPwkJBPrZinqmfiHhPOVeVTcynaDmzqxoldfnBSte
LuhNFaPSe0kJO7+/vVMsFjukZkeTLfzOWVHok08uFv2Tj8nh31NdrzLhwDKumDwq
dO3GaWUwJhj/mDsBRdeV70mukVt8Eal6s7Vin05X/eWFxaR1l8vASqD6FXKyHBoX
Zxkxdxh1wMDPPqtZYxQ19woRvS2D3lKKlsTuhsznXQbFRi7uB13WfQX8+v/VaQ0K
61tg1XDj3BW/VgDN+nldZiB7TlirHJ7jjgymM54uSVapen7yZaoh8GT73TCbLe4Z
6s8RPW6LpPkQWVkLqZj17UpT3mpY1fShsBGNElBfBKsd/1cfzFdK2xpxu47Snc/z
jATs0JcmK7oFbd3dkcvnXukx0FSlD+bIsKpew1f5L6BtWyxtyk1fWYyaeu/owIAZ
IYtM9V2MjM240ufY8tLfd96rqFtwvnQCb3lFD1MkyiEd3y3Xx/reQLtM9J5fMwxN
AgyQDDdy2jzPt7ZScdBPQ5s+qtsLzH/MLPzav/LCIpItsPjeiD6wMbmKfuMQdXaJ
z+Q1xU+rH85ue9ryQoJrc9tLYfy31CfrLFTBe5l8tdvNbNg/eCd+Y+0/HCmHfaxP
04Riyihmy6aweLvQ8DcSHbIvrBJFBGfckifHxh7QeywQy8ZfN5Q0shGgJijDsYzl
oqecWpPTl9A0CZE01E+3l6c8RvOV9KV+j7pAt73R9hkNX5qbJ3xbLpeZ4UsETdq+
Oy90kEyQy2aifr2mjBHZoXm1I12J5HBzV8D+3Buj3/FLqUO86Jlkj5iACM5AHMKA
swwzTyyFBgSaniFQDQYmq6a03s/t+wmS8Z6gaAwbA9oEe/roKfmj3tujWNxgGhSZ
gGTGzlNmHcSFsfEghivqyGTqS0eM7zKU9VpM71cIBdn0kTPMYo96TzG/TlRwqf4c
SMYgSQ2+CWnX/SvMaDxyrkzgWMyP3NGXAzbrVQ6eWt8ks/Makjf8V/7Kls0wN8Lb
nBRiX7TFFelqFgSELZzFq7DLKhWd4z+Wg5wwrd+F0aSdzonIS+DF528JGW8qpyA/
ceALFil2AG4Y9M79wc/5f3o0w/DOo4c/tSAIPhZgXT0fYDf5FxEhJLCZgl0yiqyQ
hu1ZVys8qNZQU+7GFzYCkrsNqJ6C0KLjXfDIdhWqOoomzdnVjjGLcf9HUUKdwgm8
glUsA6dpJ8GcgvUN1nWRlCpll9Axbbh3Y05qTMCiRLxNOCVLRnb61YSxKS19IPl3
2MDRHXadLY4w3mIOPI9zB7CKR3haY05SvMOtRULXj0tD5U/m9TDbmHHjBgas1Ltl
SygrHBYeCnsjkdVr2VnLbS3w5tn5Izw9BwtwLdzg5jOWA+/Z7eAvJgsNs8JORbPy
WRKpNeuSvaZPCPfX76CjjNZaorCXvP7Q7whYdoSFQN1UCpLbZgcuJ3rcx6AdExc7
dMjquU7Q9+1Hi8RedfOXtl51gnrqKeB2Feum5AFb85NOstsk962TW0Yu8++LgSd9
kfuMWOftijV89CvMcCEGMiSm04CznsbqGt1y3ZeqYiDgDfoG2N5ruvycsRQcv/bf
SG5IW9AZE8i45/TAAiGN+OyFMGRlFzG2SPLtMBwYzUWS4QBx6OJpNC1CynG4wIUh
w9tipLASB2myx1FUNE0z5Tn0OYJvdDvyrXROQJwQvrwUoOdv04giHf/XFKDmdmpA
fsuq3cVhuuQCXn6rE/8uJfIMuK/tQTw6ETTNkBGzrQie31rkChCNZmNITAD5M8z4
A4TCZfy/LIjYJ4UwhLnImEY3cpC4x1/PJIvSZS8QH0NWuA9TPB/+A9mRWEcA0zJ8
QoRvlHlb+Ma/gMuF89UDnI/amVpPKIKvW0BeTVsVjJ4m8Gms3oKevngTUaUpf6qD
yFnwxB+BiUq0Yi63/bNYhn7Nt63REgV1ATvUhxOHMDWCG7GdVnB6lrsqkjEF/SJW
TqgzA4yYfoOGI8UXV5rPcmd6g9bXgNc1+zOBD43Um+FRvVblWaaz2gZAEudhktPE
T32UyLMAIGk0PihWP8ByVTpiUuvIcqyXGJB0G9bNXYyzlMWv02iNXsVXSAtCMdIF
huhjqgrnmrGGZnqyReR538T3wzsGRYSFjUTH/7j5hG0RYN2lBJp3ghJT9QPw2yjK
16CDRVhLgSXQ888W+uwygAUcIUmADoor02Qt63XdEUGZl+OcW40zuY+vJYKNm5Up
QAG9Id3/LYra2R5u5wMom6rlwfC6K0wk+L2KbhAlV3crZC3S8ORPkYSFMnf9yRN8
IWBu2qxFK1p6VLP+F9jgUcSl4lyylJycyWsLEE6cxdFZTeYv1E8U/w8HliXVQuZe
DlvHssrqofXT3jCmPHwBr1upUIjxVytE5kAVE8oAH/xY1pN2PjU0gNIHQgjDefhs
lty1JLhUBbSiNiuA+AQ1tkZ+dFR0xNJbOdMF3rZkgyAwhnaxZ2W4yj+5zKTF8JGt
R7swens2v8wmcLa8meE9K/COWStq6PMi8En66QXmsX2YBH2kL+JiPdzlF14jn8MB
V+v7h8TsXIio6+DiLVvLs2rsJ0kCxtk9YV6IYZH6l1oJ3lOjkWoxxWKkvNSEj/W+
Q35XS+5uNMbeDJ/fOBQJblFDW1V/C/J6f26+4KGGzujOE14wLgAMWNvaZnhmw1Nn
sfaDnNZmWtOPGXeuIUnphLjxIYXkXivvoEw1lI1CV3fDxaIA5UnmQedf8KsqA4Lb
7LQsoqwwOgv0Fml/XblYGR9ZPvs+VZOiO7WYZOzN/I/d8tsDXgZ6P89DLf9EYq5p
YFJcInQnPeM7Z/+l8208PtnDN7BwXQ/EMJ2duNaiZN/l3OT9IMZqf4QMJFxJcOWV
Geo7Rnwi4mgMIQ1lmAt7ldeqPAFkcEeAbYzwA9LUY0nAxC719bh8/pibTMUoFdH3
S6F4nySczBn2FG8/I1KPPvrkeZvXkWEmFZrcTgDwDU6jNBIqcrONhi1KhBdmlNHp
66YUvPXPkNPnQsZ9QtOGWH4GWr1ITIIN897seeenkxoOIRYP0IMg0NnUf6Drg5yQ
F5hwVrzE8ZVs602XE+k+hPmbz6GCm00YP+msD+y6cBvQdRbYfBd7WSMt5oo0sJaa
F7FMrOT4UGMKp+ug/VxVWlov8PXVrA2MVGBkGoJ0sA5/8DCcE0skqqQtNBGSOogh
uYG3LxZJU9yw53IIc/m4Tjwol26fTrBvte0gOal2Qb6l/bTyD00/VLa1edJtrZ1E
fNsXbmSrer88G0Av/UzDgjIweurhmWR3vyoPKqw0KZhWJW9ZSirafQNhq2Cy5xja
94cN4HjJL49NEPF5XDZtJRa9Lp52cwBQ59fZ3GMmFP48uC1NTJ0yzJkhXi0tyfGU
TPHz6OafwT2aC7YKYVe1HDBsbPCY5R+2U8RiXDh0/mNRo8KZD/MT24XF4Oz0rjo4
RXjtMJcMduaA83qKhqgW84+NuMEsnXmIsEClgtkxr1T/9YdOrNL3EzQFPHDq0Tyw
Nkg09rZtZnCw5zsMiKFFggMT3h8l1IZpPeXM5O0YpvssjOJEokTdNj70gCyO6IVh
SibGuvkvC6kvC0LlCTeaEPXOPrPELdMIBgHDm7L496dkWNZbgd7A60Zm3Ds3LcZ2
Psgbs0dX1eqAKtlEvrUOD9KMCL7CTQIiAZ54yg2Ft9VwoZE1h2r1EqOGNrvKAlhT
4+Ypo9WsXQi6oGSP7x9ITQV/BMr/3fCwpJle7e7wiv3c8Hz5p9AX1jmAjx3rfn0h
DvM/rTdaXsPcwXye7jGlgxydHuLLSii2MDDBt2MQyt2hqrdeZWAfUoO6KymRZ7js
fXE/WWWnLMvSiQNXFbTktx2NWTG3NJgXiv0A8Yb5Q4vulUxIgrWK1paxsVGrzXbN
Bu9nioT5W+tUqNlOHGA0+AAQ0ZGmJPslht3P10Zyr86u8oyZJubyCNmKV9+7EbFJ
CxivmIBFdI6P88VfMidvfyN5AOZMCm2egul6AJX9/oaItL6DRZDInpLHKG12PKMA
LiaJReMJA+eWTMajw1EUzJJYH2ciy6lj9VzdeA0Ch6ELqOEcTmm4SA23gQhLD+C2
MHAcqgNscYtr1cfc0A9PoMZtex+SG70w52A1maXwD/uoIFZR+91gMkm/qdRv6jI4
JKXlmOGBu4sTAf2qKZ09h7EGKlnoZ3FAhnUBOSdagHYr6cl3FJfCVSt+LxvGnLvN
XK4o+dKF+7dTRQbC3Nr9tON217hPIcFbDH16UGxXNGP0Yzr79kHc5YNNxeRy7TbE
cV4jyvSvkVr1a51vQI/GVjHaU8oY62vi4j6uLrSrg9wcxozxbxeWtGK5cSFeTQMU
l76rPO/TLf0/AywvfOPFxHy88vcxjVPunz2GJvbdGyrzxAsPSv0pj5JV/96GeuTh
lmDfurU1szgaTy9nilrZOpwiLhLWBK96U9bSAQoB+3YwqjUus6YyW++WW2wpb+93
pRfnwKrFys1Lwac+Xgls1ukcFPhQU6Kd3+68YwsP/A8nHv0g3mWFW84w7GfQHp+A
M956JPxciwUQL8Kyh10QZa8XY5dn8lkyNGsaVMeLSeRbjib8dBCcI05Y73aQ3+uU
a51CbKqr+Z6XyhroeG6POUIZYFfyWLhJchKGYgxFazICPBZr9n6cAbJtNpXCFKmJ
kuh6uQGe7PzI3OJnqm9i4Uhy1sZDi6YYBzxjgYbLKYp2z1SO60M+CuoXy38bSvl5
NeK8lEFSZIKrmpgCfbiK7qawH7apBestQMcYIrC1ReT6Xpkc4Fg7nUjxExMS30hP
gwRRvak6d5MGa3d4vidHpy2cgKJImkLSEHc6vw5f87shRvU/LW155CNz/vfHuytq
I/KlTbBUiYumYk25j9by2Bww87nXDSqu79NkK6eEidZggEcrBM74jUEdx6Zno+YB
UmkXBF/QYKeYlrlbDyX8CH7Om4xSD8CMCjMF9G79edIeNVGWPRdaBxMO5Vfv+VBV
+Kwdp9eu9am7P4nfbgbyfqRvQ34X2FiluDRUaLjEPMmfqrs96rv3HsJZvolzk7dH
EzpoJr41xgfBkCS8cE4Mksj/CDwXgc8lBSkUZZjvuMLwskuFPlbPVsJjP3kdf1R2
+kJGXCMLozw2FT2oxq4YhxOPNEFJ2B5RISPBXk+BCnw/KDR+BYMVCM/tRPbIMs1G
D5dkUbKG6jWuvG6YDjm8KE2LbhWzQyF07drCOhv53hnku5X3SNaZlzzTku1yVWVX
RZDCiWCCTvi39ajk72FxyAQHQnGYQH/CVnV8IowSL9ERt80NcjtzL+KmM0ul6Ett
4Ni2jVPLuBbsulv7b3QD2s0Ik41U0S8PNUKcuphcDOOCM6SJ8xc8rV8Nnt+2l+xE
GtTIRfC9tIkL6qos1uvkSi9rhzgL03ebq61tPhqYrExz2/QQq9PHvAXI7WiTSZo4
EXf5G441hQXjGqLhlmKsdMbPVQGE4V3ZP4OltBzO9Vxgr4ZE/yqHCvVp/4SMicmo
2RiTwQHTJfn2tA9qeuUKaeJCucEi7GwERYp8mfPvruAV7AQP5A+Vyfsws2yahWJI
g4E89hUMhvfe5GTtymDtvusAFxGMv+6tAnMMCCgLGKADRJzTecMFPKqP3ch/Nhot
XNRvswZy0EmCEK+wrcp1KO6ol1Hy1Zp3/mkDOAE1liJ41Jq+lhX3RE3tzDrIAHf0
sWBn9WsJLXQT2On0QLKB9rBr0YrWg9xtb30sHMdetQiXk7eTtr+zUH4h3jYa0fB9
+vvKRC2x0pv8NsIR6DJRNCZ22nL9b+iOyx9ZtOzw7HmRydvy2mcBhac3yUTNmLj0
XjR3iSSEKxgMY0xDPHq/5aTKU1pGF09lCPso3Y6meZ3vjNtgv1Om+uF3WMeXZewk
PQ79JyTsBQDrlgQo1NJBJpX+1d3W5GWCVUJdcc5U6MCkGd6ZitF9x7TXrvDxa96m
J0P/5rkAyu4Vt65F6woyNMH1NkuxRIc7nvkQo7EMqgOvd7wOyifoCbqtrjImtiKv
5smovs3GyyvjAzT/C31cZb2VNusYLqKdKx1I3hcFRSyMr80hChZU5UNlLyQVS/ig
xgAw0h+KOTLqIkUNhtrQheIo7zGsvFtW4g4uZw9gwPWfzw1JrAImBFTN31gP2fm+
ZduueQuLa/xr6L4oDiUC+UUKo732HLJdsfTzMPK9q40TZjoRC5Fle5z5w6SxbU7/
555L4gnG/qJaBl5G5NnXs7QK1TNYrbqZl+fNF6hW36kjgAeQ7JnhzeXGV8jOL7cl
K9tqChLtkTIytOwlwu2VZsjGAuke5/SL8sZw+pBrE1wNdW2VPqnQ3FbfGlsHXmln
lBqfeajmbhiDz9Y0u3InPwKFoFPGv35ANX4W09iExKYaQLSZdg8X2lg1gc+cXxwL
0vxeB9CBx3m0Iyu/VbiAxIM/oD3lF+tWjXWFFnqgTk6gEuUREyEscdVsPjFOfolQ
ogAQQHh7NC80bzyb+Np6IJZ4bYzTdBUe69xXti6iD/wWfe/DIRFBy79poeDzcAoy
cGYIzTKjKLWuu94ujsnuE8tfx9nmZnem1IqAnEqvcVaCLIkNSfBHt7TxdBzgKfDC
Po9K52zqMvTNw9lDKdbffUO53gEu1mDthDHydeyfsviMyoTbD23znoS2dUgjfkZH
fS5y0v1E4lLRdTofgaGZswmptVQn8DAZv7/uC9iGzu1rhywgtzMLRjFV6E0TWHWw
xIhya1cfM0GZLgKDfNVcjkuepdNzF1Y/iESZlYXok2g7euvMOqbAvMgg2R54/ZLx
wB7JecsnEs+teSfa1ls/m8N4z6NuSPF9SZnw7lItKWYNRFlf9yYDHTvilwvPvRim
P8qqN09GxZe0Gwoji+wZpmP8utUVfULgIkA5LMTodzafp3xBCMWzJnqevYQ2unTm
g493NWzTOB66ch+NGN25opUFPn6F1obrRwAHgoHqQ/9q6czjfSrSZvtZ59AUHeiw
qOO+A8nlAFKqVKAyJAmxz1y0IRb4hqVOOUztlW0sZlCI3y0+yXzOnyS7V5+ijrXI
Bs4uS254MGroB7Ft3nJ0WClpY0va/Tn2VB3vHQmx3wb5TbkaIZ9O7KYxd3olgsQ/
L8izTzjiGdXDs/AAYBlW3YfdKKETgqDhFHN4+1IS7oC70uFBIWYuGEEDzsreNDgY
18CDs1WLzVOIWVqTBbO8ZdMpq2hj3KFRhK5x/iyhOoVtZND1wtpXjescTBBWhiZB
oef8zuKraCmZJLatu+JnpczpOS3JhDgDVC50qTSaPSuv8UJL9rtGi/Zd++gq3EzL
CKIUW2NuGz58uvIcU5SbJjlj8JIC3X+dfCJY1kmFrGq75M1lCqynrcocnn480Ov0
dVkJvEifhUP5brvsOpnKEPYImUemWPgmM8Ank2V1KbDnhNF/VsasNptBXqej07L9
RWzP1V3vs5Txyo0nv/PBEM6flqIkX+C3vd2gm3B/FduQwa1hc6KejPlBEq5/dNIc
dpfUpjR8X+dYs7CU46/P3mIUzFKBCl/yC46afRuoFASquuC4uEvGPHnpGRE21VNo
cMtBQ9Y6AO6HTT+44A6qnr1uzouIF6IR0FtT6jufsO0RyUUqVRFbDWFdoVXNqyD3
V9sb2WdEW19HUUci1wLCrT4/tVLQysusTY+JgrinuQ3lO06b5QTeCPyzNKBgf2ry
H+aJuTkuEISc+PqpsFPKWNTaID/M+N9GcPQchl4RlkWwYxs9pBL4N/jU4B44uqlq
mQpJB8HSaYw2MXJnZJF9SSimPplpBfAZr/G3JrCN9ipdB8TmLpbWdrQcmAW8PGCz
4GtZbYcswnePzaANkCJbxTmwyJN/q97BmtVH/8SvuARZNJb6jz8bSz7TJKQgst+y
RTG20w+X6FbpRB4LH6tXTQkjOH93iXW5YXajmvGR9KOeY1/DVUuWDNr62Ay1GfAj
jk8dxDdab6q4NHcGE/TLFmu4yVTirPFuIHCLQXTjgiw20aygK8Dn3RVcbcfyM4Wg
5bfUbMvbRDbYJRqXqf2T41nn7axEUmhAcGGX3sIleMP9tJ3LWhXnXz9PV+Hyz6jp
+eQm3OIz+PKgt0NUtkaZXcXx86kszW/QNdyd7vwy+t0p9CztwfeehElVxPtT5QWs
9ClCwigPcS8WpdgMdsL4GtQCB/7P6oFWM5WMI9jeoZd1J6KaMcUtYS7Uzyz4CGCx
o/X12tw1jSbYiPtUFrLVwG9kK/Du22HjBHa2l+2XJRZDhAg2o9sFpflXvGwTmf5M
hFP6Y6Ujq0Pq44f8YSs7lgrAnZQLrzVZqZnoagQ+9Ba9t8yk+chONOUXd8WLKo/8
z1S6jiT7btPe0vIy5OjWIb7XHv80iUN5nP8FTbWI0VapzumZ0X8plKGj+HoMUn8U
e38eqCiQcybkcYAB+gwpUI4QJhoumYJjABxM5WqHArE9adKP2oKL2Dyu1LXF3BU/
+GKf9tNL2EWlu9LNYZW0A3orsBKZ0ltkgFFeGNuOC969MEXV2tsptwkPH6TLnZ3s
oaM4bIX+SmsSV/pI4fo7Cc8iloXKf94uGDHn8dLzuo1/mrdecskGdD850LqRvT/B
GSoyKe3uFdITVhEQMwEy9erN9tGx92w94Gxbb75NYHeSlv7C6tgBHvdq4gLMykhT
hIBzdJChEV6inP0AXsgSSu6JlWaLxb3AGiuiKauUOLIkSDzbdYnaWk1475j9vtkM
dxhJISioj4L/hlM+zfFW+QmME6Ld6RMRH+Vh8jdGmaW+tzt637V37cFoTmrfoLVY
44qrNoLPMA59rhbsdd8GEyFW6LCNUd8sbt/uj79cyjN8oH7fDMOfkv5ruefs+FpO
N6sQPOmzvMRF06IvxJRt/aAXosNCrtEyBKMTkY3ohQSQnyzs4Bd6d4TRgfQdTJC1
z28IrCopVzK1g2vFoT5DauD5OqMGdj/qouZ6V2buWCrZaw5df8inrQWEUFXGRjcs
ejlXkmpif/53srYqLm3hOA2OR3eCahPkVFdrgVdwphsuK/5orDyEkH7MMuwiDN5m
e9f2aV1qfww39OldH31WOVxblYmzKedPAD0syWopJhA+rJNw53Tb66Y47Wa+oxYh
AFghPE5m6sf0smMd/t0fKzDj8SxNOt26MYLVhxxZhMtR9AV/Q35SdTWydOKUjWQx
o9E878t5MZVSGo8bFYgu46OHsZSzgLT3qDQvqQC0mcZcnf70pheT1YO1Kw7eLlvN
4ptH5+yC+gVVDumVr/SUl/tpCtC2Sulbj4R3qO+OFSYYrt8Bbi9vyFfJjiIgYG+U
LlYyol7253VwT/3iaaH4+oWtI18BWXSqLu7BVTbU9HankpdrOeRWadg6jxp2c+r0
O5abs5l1SpT1CDa1B+JBMUo2maOahTkVnlepckPqg5kOYhO9wSbS/tnGCZPyAbsS
gw6H3+fJzfJ1HUfei0NRf1lYj3XvVnDVCAGfc/3CmxKbimTPlznRzKbOO1yS10uq
c1nAv7qX0FYjj1WDGL3mIlNrKhWqGdEtfluJ1A5FuyLY0VrkoXJF/hz8g6DFldrt
mFXDlKEnifZj/fFTjQ8lr+c2+9uEbMl1oLbiJ9FbqJwpdqv/2QPyWmljuc2KDX5m
SvXombR3IjF4V329GoKfEfdH+sshqj4+ZBN5/ZhKv1YFVP9BnRe6ngcdq5vDqnIK
gtr9oUDJUXVa8KYJE9wHn2JGRdo3wc9lK4CVQIf5iuRmUZJ3kYzNCjxymWwc0mE/
c78uP4PBli97Jq/GiylOYFv6m1pGQdwCv94wAs8idyRmEHxZObtetIGH/2WBbxy6
atE3DmQ9mFpY6pa26ZGJItxrUvU0JmJeq8Z/Y7voHS4rmv2aXjl1tWgRP3pyip2P
rPhTx+dYqZXVQl+11anFcnOsbhv3YKX5HhUqX+OKZ75dw7p0WauF/TxL6E4iuTjG
7eXcuR9c4k0LU2+JEgYCeLA7Bc7RIBAMnMnwa3zf8KtFzBotCzhObtoYrO2qp3iB
QkBixf9Osm6BgOZTAh9Mh6anRD1/ggYL2NmsXIPn0TGKExW1NzpE14b124fCM21w
rX5vz3l3peRyZGx4weBQ6UjHuWyqZRUaUuNSWUUvrnqwu85eaPia054dRTMjEae7
7fnPycLprPoYqgdqs4fobhF9T/Ft6a4HSNsiMi4ODmmBQXYSc/kuoYiGlZyaVnEA
hZUGNp2mEe7rF2SoBxpdnQIWtAIC6DS+l1c+B4f5xpXooOevcpJ8w9xOYSslncMk
YMSlEdoWBpfbO7d5/qt/veWrPBsTsQ0LHSu81GuXJhc5jgeW0Pw6Idy7U4qbMhnf
dEW0/1/yZIqGZodgJAJYAR2pB1ymjNtPXIZ5JLBKmD+2hvlg24CMdJvU6V9pjFVu
LkRxu3hsNOoMic0XEbi1wniU9Acs+nvL/DnOilirG2FChoDAv0ICRikV+A0CbvKk
2FDz9oGYbsp9BAp6wRa5bd9LaFfqJHYtoI11cmZvQYUSKul7tn667UPUVgNV9+nu
lw3bYyAXj3PznmifKuFPF66blBA5FpCda+7VdhmWvrAfk39KTyCvftSkndsYrhVG
yJLPeaSMLB3fmfCznCjSWi9PeaetFP4uMVl1X7hBpy1i2ZDD9WbIbfo83O4lzbpI
M84v4jGOdK6NJ0kEm/3KimAKJFQdLIBPgX8enBlJXXxlg/5mev3cYR2upU8tonJv
A+fTWT6Ty+jLgi0Rqbt2u1GyAJrf5fAd28tjN2b4sMwxQMysMOQEnevIwzvq0X/A
ISIQC1d5Fk8KFpLJJsItuBpGiCCJT2MBB8a5oSCuIyuJhP+iMYed7njlaE2dAo4X
2Ub0jk4Zw8EvHm84Z4EWxnAOGOtUdolMIFrGGyiXG8CvLO1NMFbUFqwTZlm7Bz1D
u9kGXh6mHCA2IRm38WpqI/RVxJnF6uuG0FthzADqgOxT6rFyKh3Yo+fl4+MU87s8
nDcbOiFaFNlOT3lf1eRswT0SSpKVWxgG/OHMVgcdblHngYkbA11Wsfe9gxBRHShx
6Y+yPgcSy+AuZXlA0pcyKOg21npa1U6PEhhRG4XPOUgVWgjORQHNjvT8S1JFvsFN
H+C5/sGJaL29UKyK5TUy/hXQcoh6xkDirTbOD1bVDQlM3rbilLQhyhDaqlNY+LuO
EnfFrqn1fGKHTmvDEn2yQ7iV962C6Skw+oZC9ST2zzGHI2v1suRjOb34YRTggzUc
/s8DYrVqKEaqgT/wXuorR+CO71Anm//aWLNuYRPcdMHVmbr8Hwq0K57Gaet3+1xg
+i7/QIBWLR0w50fvDedMtwu53/sE7cKjg+gpkSBBvy6Hzjr5L1mvYEBRnddkYAvg
KGLnG7tLRZLG8Ef8UezfoXGVslHwEC5wrTaakjmkBVhZ41n/ybPuBOgz8NvRBv/2
0wFxGob198feObtO0KhADjseLlRZFULZvtK/FImjpEsa0+9RHe/9M2lzXUhkoPEC
02KE/Mf8a/iaKPSdJdplORs1V4Sv4DxgJj9bRX1fsoldT184Q8XnOL3VN8+GadWU
NJTiFTMeClB8YZZoXwNsoM2Lhi7c3JT479aeGjUT8EVFwti+30pcIugWWhNrqDxO
6RzUA4hUNC5VFq0XSD3sSkKiBpHroPLTMQ20USXHQFcmhNN0jFDOoP6akCYq2rrV
UQADhA4adqHhG48Ozv3bNXYmlhawHVTUN95oNdsAVvK5kB+jZFcv+WF6JTNgtpPb
fE5S0clxggyU86zBmS4qfda4K6W2QPWV2wF43YITafkJOQEqSMx7TOQpDfj5BGXO
vh5/ai9Xdgx5S3FdjCs01dIdnq480snvTfgqxpQ1IR9uzrl0ocr8LD942LX0sNgo
bef2x1qNpsXlfmQpDr/uQht+wXRvymdmLOWYBnVPBWaCjMsHYP8Demi+xZPfA0RL
/yZWtK4tfrFaQe3x0AajJeVqH1yut2YLd7viVCa2ov/n9wXOjCmUHB8xprzqYxST
kXFtBuvtqIZjF18Rnp8qkpyopmuQuxLbrIIzcJpSHAtQHbAeW3aRNVY4IEd1z6QD
lhv9M9gJ5x4hXZdqyWV/ZvKckJ5SvAwxX1RL5eeZKXq0jnvFFgU0Ym82yhLaQVXc
9HYeA+7QCEyM2FVwHQwoViZBxjByooDTqH5P7SDXLBoSGhvFB7NRNdnzVHMliMgy
HG98fWfx3s1LUdpgjyoKXcgfR9QRveJ86ziJl0hAIibaJl7EH/QEBrC4IWKsOpvi
h3JJpK+pKBNxBWDMPuA9cW+L2RLCBdF8XDcPGSJxXytK196i2uk7k3YJXEqz3/QI
Ae8kuBC/4MeNJj1arvWJe/lHbW0sFPIxPUn4CuBJqKbCISIyssXA6tVKu3ye9wL6
9MEZtGAJ7BM1uq0MAHsfZ3E/9/HZpnkTWsKUoYyubUHdh490YTxy+dzNIeT2BTTp
CvemB3yJuDmCTr84gBhLDqco3upduiofAeQyXnPdvOXmUb8s6sHZ2PdBlRw7rbfX
ET8DotNlMUi3nhl50uwromWygvkYiJqJWBAVeUeWaNb1OSQJrubgtH0WCNVPk7MG
8MEHOdZ8mDmqB/+wATEs0YWmH9+6Ayyqh7mUzp2OZCAb0e3FZ1oKE64OytZPxi5y
ozxKhJIlwIe2hcvAohoE3d/UA7L6jbkY6W6Z1CKF3gX1C6XKlP+DDSttHdcZveb6
z/O483tNCBS+o8daBeBdHSek2Agk1JqZO0pIK4/t1xeOb5UQPKQuiOkBTHVzTDhJ
xiN0sHdIEgycPgn/N8xpn0B7DhT9bvem3xtvb6035eMmOUACJT5vQhdmYbD8aJsF
QkGP5fBY3zerNdWq3lpwKuJ88NXTTONLiPu9+oNK1xS8p9/T13ZGnPwzt7beicwD
YBlAI7oHBzBB55ISYup65WSVDtwPZWF3B63RqiR3JSAluCHKlNws61I6u4JXFPmQ
8J+ik9LAlVgnscIaGfhnCMxRheOq2KyE/tPQC3Xu57o/8wRZw5dQm1i4Rxd5XT/o
VllxPPCDsIxcbr4cEYm5c5g7QoL1U8mKu8nWEg136Q1g93OgqJnFAm4HqGmtiPdW
+7uxUYnCmrs1uDT3dIOqXGfLy+0UpO3R/BdzsUTKhgyzL/DpUs7G6ALprrBJ9/fP
MSLxfP/NLq3hdMrLLvuQFO9OqvwZBYx8pg9BvCAOZUk+1dEk1uT2PLxnqtrOP1bc
GPObX/sR6Q6GArTmn/cactuv6Nl2uaPcEklngc/Rigsv9+aza10HZtR2TVws2TRD
VtcK8VLm8ZidZgNwON1BX4ZIOe4H2kAYistBR9s/ErIIu6NjzqE15KB03Xvuu2eL
Lrhb82iS3TDcQHczLPVSM26iQTKLKfol7n1jORjjZRVujgJ5iKb0HOMpJze9I/xT
UYykjpWs+T9Eu3OFBdYwBcKGZrV5ksvzjBislyh8tFkkS3B/66ISYZKxoW/gQsEs
1dtfotKmUyT7uQYRZF6uw6BNnqcFO7IxoZxwvxjQ+t5hPq1dttWkcmmiXK9WtVbg
4gDItBxMJKqvhcVQAzpnbsaFPPSdlnDLt7FyxiSNuT/t7FomJwRwWUxBB8vbLcZw
XMXm9yOqR/eLDac9j/CDKFiVwbi46OGSlezvbgvOS9bBbimNAr/giOA9amBFt6Mz
sSBbwlF8SW/74WvkcURfFlzkmVBMeZK5JJQECHOIL1EhS+UZxlSmArBevh1xxsBr
UCH/CVVNbh75KjUkfQobBD0zOCym5hzHhFTG89cooN+OCMAPoY44c3+O3Cn9h4rC
JYM+bmO6xJJ1Y9mixv9SdovMJdjv7a41ZC8EcbuMsDGUpIh8RgmBoGPjtHWgp12R
TYo1rvBsf9a2/grCiZzcsv9Vb+qdsFoY6CWoEdPyA1X14Ohf2hrLNKS6BRCIi6oY
oTTB+/meNJPcYnp3wpLktwzc0qL5T3rBFJMrgADLsHchs/6O28T2tS7T9Z7h6pNj
WVt2Jq2HlI6DtxsIMkmM8oFPoHGKQ6SZcsdZ+Nhz4Q/UZn4gP+rQvj1K5+z++b7l
jSzcUibRgEDYTAD1A3iqu0/ofU72JlcOcSc9G1vmBOtSghJ5Fmn0Q4TLXjnf1fdM
dsI06e7kT6QnCmrDWhZss5lPHakviz2zarnKIKerUtC63VchD+QlEy7Q/8pggtI6
H5H9lkHVjV6n+k42/5AdZoZW3NlvzqSv3JlrofGOZhQCCknNgaY9auYhCpnUwvy3
ltOLcEi20I7DljUjbIBm6zYdpigkjQu1HHRQDeOOuxIAYNZREg3UPArfsrt0mNVy
jNmDO4xysj+pGv2aYqaJlrep7sehv3TlUjoC6aoKJqDBkBKttuBAmfpImhO4S6ub
ybdNN5VCOQ4d3liFw4CB6J/g6m8xCeR7idJ2kLgTJLkv/G4y8FmXQGGGjARrZxzb
RnpWRjx0pbXYrtqU8vOdQm5Aa4leRLJXeNGFnNbwrl2by1CtCejThJQdWNaEAl76
mkD3S+JyYQztjxgeT/yh8hEkl+Jmk54+GSaEvTYJ3SR+KVuVp+3HWtnoHVulqqeJ
7OCxVC0uN/p9mqA5tIJdlZbhqnA4gSC1nd2kFa3E78eLQJNTNdOyxyODIFX2uRKM
wjMsvRuQZFxLz5Pwo3ImFRHYe+fG/BjAz0JO91/j2Kh8y6J/aHUrTNtk8F9wY9F0
1iTOik5+Oq7IUobfOYAqar6f+2rZxIc2OkqOhWY8KofgWnZJlnioEVc/7wbwfwWh
wpL8SgpK8Yn7fuKGXzrm28VZZ2m36ELg58zPFO/I2O0dkOHhywhXhowuKQT6QhLr
jAX5LzR9LqqNggwoESb3lJI8LaKBqZB4udT8km4M0el6NhtDDoxk8OdphK1h5z6N
3ldKGx2T5YtWj0JFJN9ll1Wy2ar7EGTDO7/YL4uCVICX7iLFMssebe40lngWa/KA
2xg83OQie8ehfL+WZIP4CoSnps5bbh3cokxZeVMW4/G13mcI+xc2R6iQk/9tFV6D
favNZ76KONCB0GHu0iYS0TbyjOhGBd3L/Jy4gypLQMCg8WpA34HIIAZ+BZyOYrO5
xr9kWtSHoML/FQNm3U5KLgcs4reUNaCSTqGMahRnqoGNBb7CnOPao69xZ6GDBL4/
aW0abTtd7DNECZb0WY7/87zX403rZtrrhN3BfE5UcSKcJhSos7xH1LNOtd3sVgQz
HMdtxCSKmR3mE3fv3s/A7fQHGAloSq4BfUSNaOgFqy605u4hwbKFLhXEBJz17Fvp
LNMk3VPR0rZehpauX0M5DAxIYnNRXBlfQVyuKF6Tugpm5bg4tCDa3w7vBc8sO9uR
gaYx3WSn8fuLDTNtUlOAWOsEcviMPrdNgIavJGtQqehzJwOacg+3PvcHUkbbwrIx
ynoDjpwfWElIStxlt2tFW+6CtffdfejCw6v+MY4Sc82/M97NsUdgqgA/K0q3heV1
l1baDI/RUe5BSqBh2pVfRfQo0joLPxjpNheD8902euCkJbE1vccp6gJOX+GqKqGz
Ihw1xx5fbsVjC2B9Jcmnki5VRU50abpVhln5LQS/aiGcJchlCJyOdZ9yFEpipC7B
WCEViEH5iMTuvZJUtrBXbd2t/2O8lPYz1PLZi60cHmqnESW/P/JAGYM2v37UQ2eX
DBcAh8i3cZICzCuNTLWImwouC819/tkB+VsqF+tF/fg6FEcY7WKN6ZIj5iEioa/v
YbOdmPTj6Gv21ryiK/1HyrnIi4DIM9OpqVPsqxpHHmKe1klP52mLpIHib/PijERX
ecIWKRB+afqwQlxjxWC1sbTbngugT6lspFhI/hREMmAQp2fx7/6ZWauzOGusYD1z
NyWuoxpj6hadRaDfl08/6UyMlVYyi5X4GIJOLDCzQt0OHOnEtOfBYWxPPKLXxbJm
dF7wek2ui0KqgjRwPC36uDw+iTvMlagTjdAiqN5i6vZPsrlh27lvzCdlehAGMlzS
yzmnsy3huB2nqf4UETOIQEjp/29z2OFGBkb6mw8Bdd2vSRrvKmWAk7gpMyhplSTT
UscibbgmzuLYWAdnemX4kxfG8yKPa96jWnKHKWBt4tMP0fDcpIAdAuKx7YkxzmS1
YKqrsDfv/KQVdTks8SJP6mhwU6sMf852npK5cZwIfq9k05zMjDiu787yOY4G+oEB
MThEuWlbwjGuZdWJZRKIdqAGoWz5gdO0JaERgyhs5Xm5B6WY7+oqaRSjXFPR5W2y
JDyNbQfKkZPpx++fGyekRx9AExrtcYVxUNl+tCtaCxjFmaYg7Ob9sEn3/zpaFZ/m
Q+cA67++Woe8kQcmu1TOovm1cCLliyKUdqs709zq6cdiRy5vT95W0dHXGZ8hHPTW
Ld+hrb1pq+0560RR5Uqb/G6racVC/Z/U0oGvDl9ClNJJs44wnwWHgh9ZY0onEPe1
jVvUOi9d/VFAR2vYjLpkdKbdyqO/ZPFd3xdISQR++a0e4OtMzBMQdEKCOybXYe/L
Tibzb/Ysqjs2S9ZlVMKVlUNCF620gToGrUijBZ9mWu4ez0R7BffxpFjg2/fjew9+
mSLBqsW5cmzcwbf4wysQ11YETPiSQeAFikQdB7ZruwVPx8FcNVRdPr0BwKGQogQw
u7WBPXEh8Gb3BZxCdWTpiCVIZmZvmqOLkCMP9enioUjhwUyjC39k5WnRLauV2bTb
lTAllRP87l46TKEOkkcLV2Cj9upJIZF66Dh1i8zqiONYOvfU1ntGRrgzyQ6BzQVR
y95b8aDzrwTy1ENcIPUF+Kaq+RyT64eW0w4nFkUXkoXMUkxJaTXflW4sa0/n8M7t
hrJ+dUSJjrI8mEpqHJYNKwMMtaEvv8tX6uV7Wr8CgAOkS/p+5soFfEagbrPMq+Ci
iL06qCD/a5jP+FuzKD0UV+Nc65L5Rn2Z71AiyMczJfUFhMUxOsl4Zk1/a6K33A91
oSMKIcdcWcwE9NRWcZdFI3c8kc7xzcahiQkm1HzbEgFf9USspiafKfwsKC5nbPH0
8A131D5IvzJ4EALZRuZKOCEezIcDZ85uwzUOL/LbvT7WR+vrsWxU0nRDezcbKnBa
zRdbZsjN8Av+cUmeBTktBfkttl0vRm/NFqj3lqBLlUffS+Wy6GFCKEtZDlWwdt9q
WxZatj0QWWfbdt+pbGO2z4K2CF+vndfWYUcYOVxLz1owHiQGbTLG25qZagCfCwCf
qBeHwQa4Rr9+1ZJS1/2rtz0rc2GYWIyI31y8Zn1qwrWo+Qxhkm+9ItjXNwnrluxX
0ky68gtV4ez6y/nFXf2A7LHBHvBIXAw05Pnad7E2YxJawgmh8LJMQF4GlJhiP0uX
bArgzOm3AoMIndwx9qr6o9CmuImj6mk63ODC39jy2oc3WUS5fL+Y+xUPk16RJhMd
EOGwCjz/HmOs3ig/VnE8oCLxCi5GcY0yYn5QGDLXyqQJh+E/smoptkCpfGDcrTj7
T3OG3D/6ob6gBCkYc0ZNnajG3dMpXy05tosJ+Y2W6ayYmgAV1iav/xJLOZS89wAL
5ifAe4Ovd9nnivAcx/fWi+44ErT+n2sY2CxcOOqIeQXbsExWm4qIV/9TaeLofXNe
NVnZxqP22Z6Tj+MeCctMjFIB4MK8AscuvWbgYa2xCFP0volGM8CKMtrhZMx2uZOm
DZHhZatvp16HtqIev6ofZjoEfT8rXeGMXFlpnZKqptStXwRK4ZGMMgVWhHYTLAap
nTSZ0cgq8mIDSD8mJrJAgb0UiynoN/4bA5JoMvFGKq+uDn4ANo5+Z4VxvqWfRZIs
3skgEZeXbTGHDk9oPP0t1nIwZDAMmhg/q3EuVh8qSe9pLO3nKl7YV38E3h5rzNaz
9F7b4+FnGlhArAkVJrCV/8DDGPRvAP4EA1CZHvn5ViGdAZJ5y5KjUcHJTPhbwKAp
rzT+scMAYYQPDXyqLQm2bZNo9GGomhspIy91Pw3VV/r60a5v6zRPxHeckz4Ux7dC
kDG8cTxHy7H5JAGIu5TR/l0XJMze5DH7I1bve17ulEwK6OGzTNCDGMP6W8kOy2BI
N4CYbTt7f+0RhPcD1T7xFz/C2o0FI8mI+lRlb8eRahREaUjJ9IGofL9Un2Jo2CQT
3TPuhIC9BOZmpS6uOLWXjmnPLslHuGqLil+arBlC7P3F82vAbELJ/ubp9MJaltLK
WHZ4u4nQIg4H2hSZDK4vbT7Hbn72ABC5sfoGiGZ8lVUm5gfzyKujkVmFhO8ZcPHG
j4JhNRIXhurm4g4ZqBYHRFdxQXlPN2L2fW/q4SkX2qKd3m+h+sl/DKf019s71rY7
UscMrAI05Gj/RW9mneQQxahwgpRWCMwu48BiykURRSo2ARgeI0x21bBdqgMHKE8x
0uaHKmbR+JLCwH4ORnI7mRSyLSpKGXNwGqtrrvX7UKB5hWIPUYG1/HxJqQd96+Yp
+gs58uszTywDik2i/SU0c1+WJjVVIAn+IK9a/IpnRs6+jmpjjd9SA4AGSUqvHd/+
BJek5osEmjPmQeioF10rnIqCd+A7z+V6fDGf+oEUrtXohmQ3Ekcmczjy+fRZt7rf
F/c5ZtpQD3G9HUlj1bpRomU0brga8AIjDJ4HlBy20SRQnCqx8hN7B931CuxdLSGA
3ZTLNeBlN1M9OiTLX64SZia7AC24NGuUxWCCKXp7HGHM/YX0CgwLJEHGlCdfSszF
V6dZxtpk7FEDvbvsQDxtkeNUG8SBD0WNS+ut4ATIP+C0SG55awItrrRZ2624QILj
mKU1UvUXBOdsV7IiwyRU9aBW+NiGJoah+z1eqi3MgibBFIOElFg9lgKRwS6kLORw
LvO5WRqL979ovIID1rRMlakBtaQmGM0czieDeLKY9RrrlabWCQc/U5MTNpRG/hF4
VqbRdwEhVe8XhiUSqL75j9gKf6oZFFNJqtqARMHAgiN5+hnphYwlSU6sH6nlomBG
VbEnQBHlXOB2VoO3mYrbHknwxQqsKjBD8Oa886+kxCFX0yYQbpd1zTfbJA9+cjkx
aP9rxDgd/fGcNKA8Nb9BlhzlitYbVoqQ5cxKNq1UxQfrB/ESllj6OSt4AAMPoXN5
srEMOOGUELliflyIXwqoiSCqMqId5t0Zhu+ayqkx9ziOlxw2b+epRJzsWNgbZ4L+
s8FiJtqCrIeUjNAVHw2IR6PiynRQu9zKft3ZvacIEgI1oZmzeqmcbUuHkLkYO5jk
OieHNekuEzemImFkYZPkUq+x1nsUhH8LGAB8Y7wbhFYEfLG38PX29YoEDsdbWBDC
jpruJ4XjIwVHIjLNAglapiP5/dDD1GVZozBJBSf5VuBEDlbXJb8eiXjM+Adju54l
rRRlLRGnKvkrSFJi96UO7+NII+/+Ni3fpl+v6htgtiMKpFdbHskV1Tv0FPsBUZfW
7o+dADUZ9PIpAacTK3dcguCRAqCbfQg8aaTTZHkuD3hp1jcWOK1b6aKrpK+ordbV
2zrZ2un8AJ99YpCZGfGC4f5E10hezlxEOt0Gm4NMKrCOIqJvnKUHy3yyhUEq6FGj
f/CrQCsl1Fznu+M6gTBuyHhqs8Y4DeTfhp0QYTRV3ni27Yoyuf5Ewe6ofOPESFYC
t+kRxMb1VY24m9DKHAttgT0tuqvjNnPBsEbeYPAAmkf6XSAZAInGusbWKFdULd/P
m6hIO5AZZ/zx3eEi3CmLDyWq1IwMmpsbGmVhi1EjdZKXobiHCEGMCymoOlLt7dFo
kEoT7Jz37Uqom6RSd0mDFLYivyPtu31+5v6oVVqR6eZsCuDGEVsaMyiFW9ViLkXw
bbHVXohPs/+9cuXEBheSOnYOVR+WN0jn5aPvx8F/Cs+E4GRKSdeBNwl1ZtShhwID
SCXtapugmjYEcY6Br8EAUTl+9CdMu9gF4uRnSwTXVZzlTcSSSpmiDm/t2dzk9B//
gV5B3f18V2cuMsiQU2236G38YjkNq7O3I5EVhkLgPRNE4slnurkYrZcCZp+FxawP
8yFiwlh5VoKiiDTs8vOMhuUYbYaBVqeOHlh9Rowpuon3zDYdSWY9dhgfJJL8POFA
pLoqJXjPiIhpLYqO6A/cBmlSAF4j3cWKrhxSeXWpYZthgvlrsrczWowBRoZaTEzo
Px20rfgBtCzKUSe+cigd8PwOzy72M5BcjzDSB3C1tESq9XpHe6md0Z1ELRaVDv+H
fAnUkco+HQBiB0UT3US1AIDB3Fe6aaH79wClCxVeUJqKHgNM/AMIKUBv9ir2Lnyb
tcceAl9vWj5FPi3XTQEwJxxF37attdajTKPqr/BRIyy87z/N/rdVAz0KZ8n0P/EB
Cvaun7Qx4gsazp29NiRyefM+wT8OhUu1quNSE5ct9cAuWayvDts4p/xkNhFh9r0Z
/W61njX3N8l7B5WnUL1EtETsWDp1NS1VINVzM9wlEDbGACMCWhi4wN8F+Q5kMqDy
sRh1ZdfLcTblRYkUB1nNAWZryO8+p0e/QKg84LBma7lp447RzdSIAjvIIasGYckf
J3QSFrZMGZc3T3pajKIvy+IE/z1uYTud4uytRsLGt//QzebN/M7lvCQKfQmkcYLw
tkDhWxYZ/F33ndTSFHEK6Ggeua/qVE5W/SGmn0eT73GvadMmp10re2Oe1zIq/juh
T93BxBQuopNbSvFeK7OxxbqHHZARtg0ttYn10l/CaA6aMh4Ss0ss9XexVWuWxDOc
R7xfj0HFQLWkmauRPNnI6AdVIUBmtujjZBVraaLAqdokmZSODKGfvubCXwbz7Nds
kyxPJGx1qC0++vwVKpsOSsj50130tb+Kt2I6aIhKUFBRr0Q6mfxfosRdmFWeliPd
LYf1NWlQZfLNs06/h1pwd11yx9J6j578ZsyzfDqaPOK6cNUaE16sLtu75KvS8G5W
YBSjgK/QFbhCh4WK3l2UFujLeq7/SdO/xUkcRIbYkX4MumHuGGqeFXSjWvtWRGwr
lHKYJcmJAKPNAHW6tUM1nhbcwl9SMWiWRAbBSEt3Z1KGj/7bnewqQssDxh49YnO1
cu/WoYY7e9wDtaUWe0D4Pds7H7sgksu59nshxi9RnWa4HIxVzOtdR6dOXZmaC/J7
F9v37/AGXj1WuqKBnBoqJuyFE4fa9qlgsdwjgOGmPna53VOwZtANRdCKOX2tTFYL
bibNoPiEfCV8Bt7S5eWN/kGJTUYl51ig04QSDHvs+u8BlreSgixlc9EgQe41gMmy
PvDq9YRVzI/qetSDlbTyOgYIRr/TD2hanyPYEjwwiSYRAkkMntguInaW6AcJGqJ4
M5s0WfYxWas/ISZUgEyQIGgzAQbwqAN38+2YhUI1fdMzzPQafOwcrHuzqjW5+aof
l7C55HRPlY2QueMdMn0m1sw9W+U9LA7Skhai3MWuaB+QxT3UkCnbLJrmsCjAgyYk
OT4jaE/rK46/sfs+vwoOesysn5nTpnyGd3oR0lPh2ddnAqr4ZVOu8hrMtHIelHuF
CGjcvvIbg9fy4YhEpwn5w05mc/Lm7ptE778NguchnhrBoKRzDvyT4OnDWR4zCrAG
9u2TSO50zx50UY+f/Tbq+thxyqi1CVYkvYarryFIk6DfP6KIC7uICOb4vSgEs5Lv
5A7psC8HkciBKHvp2psTcZD6XMvvjPRuEWVA2b2fTzi2HGzstC/uAbdpl2Fw4en1
daw45XbbgY/Fd/tnFBRY4D8KHI2CoB3mJWrUueVwucnQJuhl5jL/8IvGNmUzFtli
om6tNieEVLbnI4+/LWCLrlXNHIZqvn/lppZ+kqkVjJKx0miaveCiVvtScwizfyot
GJoq8YFSrLzY+r7NTGN61ALDrhOzCugr8nZ2KomvKcmHWDayD6MGnK7ZV4G46t0a
DXG9JP3h0QwCS6p28wblDm6ePR1b7VK6yfd7cI7PSYgRy2HHv6EzVWPTwfnbVAnG
QTGd5Xl4ZrLLuDJ/dZNXbqiBmPQpNx1udjIJMux4T1aAL2fynF9ukO3vCkT+7vcs
k2+3h+6pe85CncryEXFGTBSNeKeWvmZVyCiE9uupJiCR86+m1/wDLSb3Ji5ATE3x
i3YjJC7SSZrGF1haNScU0VdzzU1gi6tjBd857e2flRBlHF/77OjR9aPFa2Yorqsi
uBHXt7YFITtOKRg73DeG51cf8cz4Kob2LtoND6NdBEyvLm1eP9BcCv9TW2JKWB3D
uJOOjfM1f6YBQHnB+oW5FZxTXucDIyUNMCJj30K3nnx9sg5voL5J6ckE+uWThitt
m3rQfin/OLPBiC2jB11hgT73VDQqU3oIEef/s0Bvk/2AH3xY1oMzJ33R2yRrlD1I
R3FfP8uzgkfIYEVcQ4Rp0a3HRhkAHD+vmZBpR/OyM55eFyCW7MuCGAF/fqapRMn0
em8dLsWPt6LafKwFADeVFogDBoHdmrbj7xGv+8ZGvTqtyNPjT/0DRD3hEwcdufby
6PZKvN7CxOqbuwVVT4ljmplY9UsnlnL5pZEB12zHmBDrZDd6M4VDdb4ixXdhwu/I
QESoO9A++xW62oL+vkQCCoo9m7W2G+5bmpbpqjBNutCBa91mlvS4OeTrORXfVP83
xbXgQuMxhCUl0g9ZLAd1H2xVOXr5eFRw997ysL4CyAavcVm28GogyNZEQmmF8oVQ
gawToeopQSVHheArfHLlfF+yOEBrBJoIBVqftztK4/1bBLLpY085cpz0YnAnfkIq
gQEDcKDPssUSvg1lawFZzgj7HgEL34QTqnQIg2znoPt06yrddn2MXitJ0J5fc8oq
496fQGnOHeQ9w8Ms7OHV3av4onkRcfpqmZiP5IbfYkj68OhswG1B2w6oD6w5oQkN
nV7H01lKT1cTvnJZUIzz7946LRU3qzqCEW+7afvt1hGn1AyEQzGSuqUAbMGan3VM
OWCouGVtvmLbp39znqvSxweXhxhAIbfbpx8UrPWFR0UTYQkTPZDzLavs+RqGwnZU
BWpjneFGoVzNSECC6cgw/EjbZNp4BGqBZQZkQ3HjntrRldKJSeN3DOnxA+uWXVLe
j/2fza0uWsq5DG7Kh/anKKMofnlomWQZSHatHJNfSj5P+1qxOjgM3/rcePvYPcKe
oPPtZP4gU/PONXgZPtKVNBQErQ6YD4Q78aFo0PSh8u1DYpHFC+oq9IsrdMt/Gdzt
6lqW3JvZbx++ZGTwXrizLKIlkLiESIHy05jW5f8dY/SKsxtK5jw37ZsKwjJwTeN+
TKHRIEWVyw+o7h+Y2RPBhIR0nwRP/5A0nrMcWkhnaT0m+n5FLNtor3dFPib3+a3N
W7oK1kOGLhPXs5Z28xSvBaDTv6cr7kbQmf7kCGyotbgItsat7ehBJdzgl65hiX3U
lVumgo4+jSEEtpypJFl1mYb5P/4kR7shXXOO8+u93Un+6XsEYPrJy1YnD2fxDwK4
cI99KgcOkVAcAVuVF+Ej/METcG7pRDp658PqKV+6BGG7dGoodUZLDXBYenL4pANz
rVru2rpXlSv++wNwV34/x0MCjkLbFMiv/Kuhd7eCBf6GvEZ4gXKBXkqqF+aLr/Pf
DvE91k/mte+QTG8YDJVMTX8CqjJAle7l2wR8PZMpOTsFQZPPiWUauSTDbQqXeo3P
4rV5rOdpsPHwZtnm0GU8WusRRH6OIPOOCC5twDUOjxEEm1K06tx+94DDOehN/Ywk
+aoiVIaJ3XtMF8kxoJ1WXTU/vN7SY3d7ic/qbUvn0a875I4K4ezMX288diIuukty
+epe+VWoL0eZkJdBhQTYdpOhRK1DN4NO8e47lqNzlKWLXptqpGasJfuGljCl6pu1
BgPxViJR5oBsJqlBktzYxZuLhYYmmBHj+N5391LZZdiuJOrfwBWQpvwowDeRdY9k
9us5i5X0kbMNZy4EfWDZGy0T8GekJ3A/etX5sT5g/j4XQ7z4bx3eRlplSjnnlkuZ
141dWdgSfvUEKq+U701eMUv9dxx7IQbomiDZ8SbQhBLWWImMbU99+Et4pVMuz7Vg
wwowaiG/72a0gBBffCHcUPb1JciQMXfOdEAOSnbsM1Q/lp8KHgO7WIettOx+u0E4
AXzKe4sAgYKDkQz4b9myqHCO7QN7EiLbLxlv/1TdJeg/AHyxzFfFbhmSNjLsx1Cz
OPv5Vze7lCG19vWbVSe+YAVT4SEiu3M++R3SCZgLaTToK1cS5yO8peLWThVsxHIS
jPG2+mQV+9DAOkjSek5OLeId+vDqoeu3imSR8Lor5nF/V5ArjWJb58VCc/4Va5Iy
BXOFBPJ0RyG8wyqdjWf7dnQkgr6S9z/Zix1qyrVD25+C7hTH0ZHovdshzUgMlT4W
4cmbx5+q0WzVVJC3hGPPhwIawN3Jq0k244xBgbXAa+80yB6/U5sSX8VY3nhGMDfw
7cx+tBwMrpRKShfcjM7T040GiGfSYfn/pJa48/bXZYJVvNfF4qigigc2Y/yAX+eZ
WJGf3ZM2gL7heypceu3Za5XQTklaKHK586K/IdtYGCEE52TwsY173LVn19Pnfrrt
wXhJRBT0QZRXSzrFqYzh2Y/R5LA6RNxZfz09FJVknyN5fDYV/Rlh2CUsLI9kexIq
tmkhR92CRK8rmwvZXnpeJszkWhtDfpeGkoTHEmCYng/mlZTrag4+nUlQ93+zbXUb
JafFOvTLSCmbj/7+dYPMMz8ekqNyGRyQVDw3sYOAfQtctxTI89yVr7j4aImOV5YC
YzquvzjZ7fNr9k7GGJmTbpHOJYr196QOqbWT+xrvCgy3aKjAlk8ApfjP1MEnTXjB
Jkw4iJFGxDGuvhuD7mIR3vsVhnjUuB/6crtMk/Z68Cw6OBI+tGHzYikaWknlx7p9
ljCClfSLtXPftDcIcwYRU5xKynVD9dQgBy9FH0tee1A0Y7FJJ/RHvswELyIGBwCl
wOa34zfR3nzWXhoFvKaixTzDXXJIUI2NiE/WZkB6ehc27KvgcNLusnUMr8ei9RBn
JvMkyX25SP4Gd+IHQNupv1I+OWcrSyuYO4NnJx3HYsYwSS8wmWkO2eJRmk329GC0
GWhDBnvVpZf9+vLGOvWdJlcU2nE92zPYYr0W3hU28QNJWy8TlsTA4Qote+GK+xZo
na+vUocfJEMSZIGYd9vaI+pJwYNB4DAGFjZnqR7n+T/Ss3mec0r1Xs982QcnM+4O
wp+9HJtbrSL8Z84FPj5m9Y6XUoZ17JDKby+Sc7c9mNRanUkPtRjY/pZl8+HDQ4/+
Uv2JXkig6ILlTRXua7Hi+nrrNDwET3GI7uALSmhUExSf5+OiO2JqzUa76CXtx9et
w7J1+bElQbbGZZND3FykUVgSdr2qfUQ/fb8ni/aEF9+SkOpHoW1n2L2AJEcVTz2q
oBrKK9FeCQb2zd5RlrUVfmRYJzWOs0dOTEMm1VcxdhLjHDK0QsbWvrryknjvUE1c
xmE7x1eDcKzdPGXk3XtqfsL2acFCt8dRksqttZ+4gW7X+GnGc//gNtaY0O1hlp5E
E/06yYZM0fihYTHdOuzzFwBDZZziHzq6NqLLBY+enoAbgCzXtdJC8Va+uel5RJnR
xub6x+er9F7XKNUDKK86TfYRPeYyrRTnb2WrXijr8EFmNLDSROpG937pPFUtN5Yi
qEtGQriKLxLgwwwQK/fb+9EZaIk8u+TlT0/cf9KL+r5VwVpNVOIhCoQ20t1SYlDC
jV5+93SiKrSbSRW5SKxb0/I8YTHhS6oMPuyIJCmDK4esv9cDOG50DIKMQwdqtlpt
XFS0A9ev/c1e1hKwmcWrg6xY2elAlKsEYusu0KuoCMIp3p8WfTEGW0AJvArCtC2H
9BtgdtYHb5nz1UzA3Iw8Y8hShcjV6ooDiPIUNtzZk1RK5x9WtSPBJ75JbzHz8skR
QBaFRtn9gyDeXhkG4Qja6J7/2hvFVods/LGHB7y3TTm2EMMpkqvpgOkd2YiYhlaC
oh8IpyXa7aE+a+UToXydxvejFNr7o8aL0C8bTG4D9jM8AqFtIYU4xg/P32CxtH82
GLH/L2LTrP+nh3d8su9YTcIGdrK26EPYKQDeFZY5EQG4aoM1o9uLnqJQZzpWfOSa
+52lwmRCsyqAl+g0kEseGtYVMr/y7J+wSvagSMC/IkvkBWATWCd6lK7TKYay+mgW
7nl2SiiUV9sBmASyCpxzKqlj1VqPO8WdYxi9xoNc2dt3mPT2D71kOnBeOpHuF2ak
WZHPrWJZxIZ/Xbz34VSO8aJjB56DBy+RPNzjgc2sbP8V9lZ2pYniSqIzFBxBgGUw
rgDductEe3T8IogsJwaxw4apF35v5925nAB12MEKXSR2ax59RP1sj+yfZtpugTd3
zg+kBLXZ9q48BdPy33nEtbIHK50V43cZQ6k80Z4BUED4oLpX5c/Uf9ttZ6NgT5Hu
KKEj0XN8Vs/EZu164FdawVAvHbh289BksOiOTFKRmNSHBNce1jtaTJm1nnJAnw+R
Fxe4Rvk2Z2YxTYJv+TQM6R+TVPgvS5jD7z9xBKs0RQwmd3bDLcaw3jcRbDB08dMJ
WVlbnuSUcqEEbyfn+70FhwxGwTMJrSq2KIlZTLpHkHiMF1dcKpySJJOS83tCtr2m
voB8L7JiYQuQ5FExWOg2zOvZFnKzDVsACCWd8VqLnM2x9mLhnSLqOoNO9RfSxZvi
ZDZtd/DgrvLZqVqsIDA9ZpnUeG94qWjgHkN5uxOA/kBt0CZcllc3R3XGzSLhZ2HG
qx+9JBIISHnlIojLFO66UW5skIqKQ/Ue6BszA0OeOa3AZ9lBbbfdknSFEHUCHIqv
I3Yj6btqlbdzBEJjlEgaBlVCGusUnJfTnsouc+ojxU5QBQ9f1cQAMv7M0VB9pslB
lIhAul95P0Loyo19vM4iYrhtFt1CRKgD4mULJRWzW/okYs2tB8SD9HJ6GNP9NTH7
0fiRKi/0EZIuCzmBZLHwqI7Qi2HBwo0Cwndou7NbDzNAMSl6IwIkHdIGc8UDUVU3
EI51tFjL1TtHsvTTNQU6vK3DezJkg19qO+MeRSUwDtHJZ+NPJNzoS+bwawupG/k/
Iq6U8LkYID7ngi6H7Yuoilorhse3Gjh0A6uaZ8DS7NTaqsR8kWrp/5JzaoZgNBVR
DmytenrYVdxd2pdh3MRyCJ9VYbz7HoMmzYagY+CywF7pJoDzkhBChEIIk7CezXIz
+0NvTD1L2MjU91HR8tROEpfKNX/wKuDRfjD0IdWuiPxMe3sjK8F/xfNe7uwjUU8D
V6qF91FG1/k88Szh0p3ka09u/FwbrDBbsTYEn1/Wn/z1TOoHAJRQsglTk4/j4T/D
avYUe0MqD49geLA9fz1Y53Bv4pYCI/UEN8PyxISsTardhIByIP4XH46X9J1bvzet
A4mJzJe7gcMeF6FzJGPU0joVzaMR+irKd4dj3p/eXn2MqScQ4c7RREmsMt3Qv3H1
ax+P5z/UrvnEoEtdkfbxTQFvjA83nOM8i4SqcIH04EWNXduoz6KQ+lKQ/5tuzfV9
kTOd4rgyMmCNwGlcHq2cG0wbfbS/4JIdL1YQZIqbKLAngjUay3j7uOsaWiVdY5sy
B8Pj1of4PCS/emcLhuAC9ytjIj2a9uc/UxHgz/jo+jxM0ou8Qgd6pfz1udCF4UiI
5Q3SpDxwBFTrSW9jJd7llOOGmb4RoWKXGoL1ir/F0slAE4O8k8bQsVyf0YrmPffL
Av3UehofZbJ4MnCIhiQ8TX67CNb2gCVdAablnMAdU1REPFFeTwddJ9wdFaumUAyK
WFofusQ9hodh2dJm8xJGa9lrWBhne+wZ+PCUbHfh3+d5V/vTk2qnGjWMLH4tPIiS
RKr+Mc88OzX4Jn5FDpCWbfottpWgqBcSDSO06ZuOoZLOD5eCthqRLa1AdzPDudkw
l1Fn3yHWIrAt/bQmMV+kUnQ5TxIUaFSX6DqufGz1rDynMh+OA/RraJ7iYXqhKto8
GFPocS2Hf/5xo8dVxT/Qe++xAGh5loMPFVDr/CqGVTz3JESjp98CW9jr1b4HASRx
3NFRfNWLn+ftaCaw436UEDG32bjRJamaTt3ItRbzRQbve5IZSv6GhjHYiY8qRlpq
vAhDqI05Eags8aGhrfWaXP7fiiud23zA/yoPkl6uBqWiBs3uqaNTGD8WEG2c3p6h
yY4GWJOEibnLinA2QS3+Wet/DhUNYCbZLOqW4ndLLypnxMv4RBTVkIat11k07GRa
sSN4C4a38k4oVgtYEvwrqgzO2HF7SWMOsPAEeYdcFYptB517yGhtzpnR4obcJNRc
T/taqi8aNOJLCkAEzEuZ8ANnG4YHR8Z8fXczTAMGErfH6HY886ysQ3cg0A2NtCVP
Ye3+cK932RXN4Sk9l9LJB4qt5Vq86Vd3Ei706YvAdi+vQFdIw5HD6ehd/VuCh7Bu
HB/x7Q7szdp1mGHOtrTxVaxR77+caS/RuXz7/7uv+LwaEw90a0R3+2th5bEnvxLc
OfCKtoPjzWHdKBuv4Lb7r7CikAzGLQe0PghVLYiM2HcBmIlbbV/RdRAjo7X7umga
+olTDjWmQXs78xFH37xy9OOANn8qrC7A1M9ZbvuFnfW18BKYUUST1IS5VFCujFqf
nfRVXiFMbM4DL+qbU2FKS5O6LyO63cUyGmG2E2+zEqI2kOH+nj5lUKs7/pDXSWHl
osQm3MYEMdU0Xtq6ZkJHC7vNdLdDOD1LjBwcPTFAdY2jWCkrrEecnpN3wnI91NE9
HY2gFVhH9XgdsKx97p0AIZ33lChTcULTLFnHVMgSzakwGmEkJEyRw6oO425j4cHH
YL0K861YgM/VzrwGhOdi/gGzu6L8YeQY4m12nEcCtY5maWnYOudjFUB3rv3HOTbo
sYVMRw3h4gGt/Q4tQOn1dw3IRu42oo9Q44loHsYglQGTEGiq/UXcoEzRFAneCGxA
cTnkGWOZ0hSiGWIFS92t+nRh7O692C/beLpYibRAPhXRfWKha7v3ICAP4PxVjPn/
0BJamkFTy6xvBzF86Rpy9TYWqfacU4vula9RC1Tmx8gmKEB9nRaMWRenHuryjah0
qBlLVFpuLHUPHipGAVj+LJ9h8wsR6A1lj7z2Jrsq+yvM0qmeTul/NQXRtXOB2FRe
cSoEjnKRudMvxjMR3IEFn8jgyJM46ZsuONLO86yY9EpTVPnMqWpuBjTVhOGC4pks
DUEPOp0pYjLV65HdbIAGsM4L6J8ygFomcPSPhJ3Mm9TLC4Izs/v4I9XIYwj0xJ4V
ThXjXG+9l/zXpgPJC5v4Unccj5IRexfwDd7lEDh9O1YpBRGomRyC32Qll2jT5WPG
jcnu6InzubR4flioMallx9dZ59F52u2RgvRak/nLavOnO6ekG6FQPy1zVkXgJzKy
9Cfu/306oAj2KBGcnMl2Eq34rsceYmclZFucM57IYSfuysROfGWyhb91nn5p/Va8
vvIP1JVDXxImyk12nGp+DnG0cveZHB9+b+QVQm66Oif8J0Tfwt+rUjn8zNBwCJch
RBzDuu0LAVsnqCoDdgeAzOXa/h0zn4HW7lKrwfjD+J1dTc5pI02PZApQ31TSJYzr
B6R8BRhvXFDjJLGMx1lQ12GmN2mC9LfepZUMzYFkFvkM6ikNmgOnNxmdTAiJmN/+
OMxIjjcAXY3t8mhxc8/fbV8s0qHOvNq+kmVIB/Nft2IFeCA9qbW9kb2SkMeytUcX
9eB3aFLV77CyrwEkFfMsMnjzk7qftBjGGkT4InFHsA9yA96/CvzdWtLfyuF+KhjD
y3Ci9Dmk1lewa+VQi3sNzCVhygVhkBZZuz67Bgr5pElVpIBVQbj0BlmYxztQuOu9
b8YZ9YjXVMIsKiOneQLe91X+5aSPkcFX/oukLYqJK/77b+N7q74j7FZpMGTWTb7g
Y4uo2Ir3rnUi8jtrFEDd3mfKvaC8ArewMFu7w7g1flyyCBRSx4cgVDbmnQTbv09R
l5ARzQDFArHctgCtYJFzga4vcWVrkmuhzHP3uX6KNLpJFHXrozuwk6/4zvfHGB65
sU6m1qMf7k8RxDLtdZA+lt7Ea72dtzRv3bPLfYlVn8vNyldMLZ07z3G90JWxMZXP
6P7c1tEg3Rzr8WVUfLpt74udQ1vxE9BGboyjDSy6xuUTgh2if+UZ5jvldXAc6wpT
36g2O7pJrWONDHgkvZZVsj/gkJ2Htsk2d/o2DhSQbvVBlNzsCqFyb35pc6aOBB3E
5f+wzv3VAQsHETnFAwTvpk2mRMOzPCJgZHcLYGfY2M/FyeEmUHyCS/MgmsU7oi5+
Ot0n5C2Lg/Sqqs82cLNmrBm3mJXYaLWBxsBDmDNY/r5Tt/yZtuNz4ORN3lhBUSic
CaORdFQRYIHkopUQS1cV8SfaXsHEIxLWgtsxCgCmGjQubvoPnlBIeNuBxg4+j9tn
SkyZeYdi6HTDmYi08nCLtXLnBw9Lp6EtqePrt3jHeiXpKiUsWYblm3TFmmAszV+c
+HTkZLJVyGHRbWQCqRk+6Grf6pkA6/ygc0oTsXSp3oZUDXwsMAjUCQX9tNeVjmFG
o6VP71Osj9yyTSHu46Rbuk3v6OeT8/Cf+jB0SAw0kDyBNw5CN9/VWknY5AZTHLSd
NDfyFyKlDhnYmQYqh0ZbTWk3XaeK7lQQzLqhImgwN4uwy/zWpis2WY8IGganifd2
CXxZk6WfAcRQDPGLUSIRo02UxIm3AX+lZ9yGQ9d7Y2afXGkav8CcnlRTkZdqYHxs
EUsz/4et6a+Pkq2Xfk61Jl102fVRYKtzIvA+wBU3F+0V/pSq6RfQ+7TmWRh+rULW
ZN5avs/v27AWv4dALFwwudIhNsu+Snkdxd4Tj7izOq7sKvfrQhOnmxuwZ7KnfPKQ
aZ5VMMqjlZm3rje1inXBglOmufOyDXovPW+l0a949ReeLDz3jDpm0R+yYTD3jnTl
RdF2WUXeKB1g0sjgB2IksFiS4OGeEo1M0ATgoYxrtGzlemgqbDOACoa9fr5whhLr
QdTntcB0Brc15w1s9lBFiSuAcZMgbKs7eQ/C0KBQZXcUdjJMYVkf19wBFVB3czmQ
04HBjagXe2Atftr925BQENRuPOHx51mL9z33Vfm2bxS5NwknVvxXFR5k9Fg9ZJC2
TDAt9ym78DeH+L9m0h9fcsGBnu513+4IenFtc4HmuYRp4b19PgGHG8U74pq36Y1H
7J4Y8WqfStqlDjeRpkpN+CnPXo4oy21A2rvDcwbZ8OyKj+W8jguzMrtD68XD9CJp
2HJJxHLRoz9f4de+F1tQ6g8DmWNRCbB18gFQD/ffhrHfeU5P3YgwtvFyKFtCE5wx
/TnghblMhNGMEEjdMBIg/xGdNnawIa40cLDbyuTYXeUwkOvHrZBF0m7D4POynuFv
8zAxO4q1BDz9yl7PDm/yQ5LIl/sRvZUIJGs2aOrW/vum4GuAlUr1vtHe76eiKKsE
IBf+VcVpXx+NT5XpM4ugZqiBkTNTZDAnSYvoBcAOXcArWtxjz6oCopMadLGZA02j
JC4ZIcgGrApwMrErovQfr4TG301Zg4YfVtLrihMn0zkEPUDc3TSk5K6VXxivP+6U
9zqhTcfOM+sTdpIRLM56E4VRpKY0a1kglTmvARBCJ9AFzTgtmLBxr85Y+cEUd5B4
yrVebEJOdgc8PE4VTsQdWRsrY8cyPs3+tAFyo6CLRSJOLoTO6PscAOmuwf/QlGmE
PrZv3IVwzBMxlq81uZVuQP3B5YljIxBROikdeTt4C4nPcqMReKQ8BgEwScvnOFE+
kkTAQVGInLBJ+7o8BND9mnX6tA5q1dFHsbopwpMD3PaJEQWCuSckOo0QEXjs2xxD
/ZKPP8yNO3c980PqhSDphfG0FLm//q1pThFR0xslOhitBAu1NkoVJvA77dZgKFtD
EoA90nX36Xtia827L1TAL5U+6qUnjV9Vx4me2CFxWxyQVxixiPTA+VGh7s+j88Mb
Kf/tuvmLzcXdFoCg/djaVD48pjTRBRz/a8NZ8G9Pr+iY/PkMoHGr8+Y4qjoTf0aE
jkLEkU9YxINE9e7V+fHRazMPJnxDqViXg7tnk67r3rCUnHe1IKolUU0qyU77XPmn
YAZqB39JgpxFoh9PdnweeoMjBYKjwBvO6oxnm8yqNs/qwRo7ujhTSQKQESxKyMX1
plA6dyte1qLUQ9iju7mxtjVIujhKYzX43kMbRDCyIl8Zv3AinUnBXuFJL5Sy2Enm
apTZokJpZ+b9/S49ZgpAcrENgVBu+AHklbK3Z0bRzqn0eSANe/6Ll6Wmi3lr79yN
SAs0SiXBj0AsSdrLjCIOIGg6Scpx61wRZLofiLXZI5CG9tNxoczkFdV1gN4rG5IJ
2V3F98qT4idc4sK/tRf0ddZxK3ALosBBtubkV5y45XlSUanUBS2D7YKsDofGNwrt
qXoX4wj1lhPJo+9gslnNsTTQBVDjqF0+/0bJS09MaId1vwpPJ1rk2KfwRcGxAKlh
byWpDusuKPsZBbP6yYtUkHjvd9YQ2+SbPujFBbaUSFXf1SdbIyyKoTkE/+i7K0K0
hKUthOHSABlgAtzGOsj6YTxaSyaNMvVekTZ8w/tGE1HvKyDY46Rcbu6kHv/QNgHW
sFXrVP0M9vEZGnx1A48WXN1GrSaJ5r6cMV8KAHAv5mt2fIflE6GrmxhP1Zpg7xo6
YGo53hPKCFeqSJGp8TPj6mABVGV8p437XplV81jQX/0fGjCXgBWC+fTTLrNoj2gK
CCgzISHydYjPF8KRP8/Nfud4yRcmS+QkkgkymUdBDty8BhvNy3fm5EE4KmbmaIyL
qEQRfBd+Kc8R/F6fnGGexG8RX323R4rEzStUncwHTxNQ9q/d1POzskfzYmvbK8T9
wiWsAF3tc/k9GxZJIrReZvIA1jVSAvDSmKFK4qPTQKLo7bVpyG9sCRJVGFecr1u6
T3ClpK52zf2f864FWY8PJtBw48wCIUw7r8f6C0UEhrldGjr9Joib+W2nJ7vaP3+Y
lY2RViOpkxJOixw003GhMbukctXNi0Her7CmkWZlIxAMBiFG96DDfGLYSPgJGm1k
b32yHOnEgLgoTdgTScV/hTJY2O3e/pZH00ylpqQ90uNxo6CSOgVJI4RbSilN9OZg
PtWE9R/q2cEy5X0vOm619cOxtfrxYlV13ek/cZa6zZ6o9uoBKC0aBfFe8OOG/RNw
cv9C867CRfL/X1uZiKzxn37e8Gjya/VKgQue8Nuv7X6xUeY8H7cOZj4HbLRi1Bk+
bBsO3yE+JssJuR6euQwt9zIZOmFK3PH905uoy+rupKwXkZM3xO7IDgicUjoaSnD6
BOCnXRvez7pB5yYglCSM71RwAgS1MjStQxPER2wTAGx8zxZ9ofp+stxdJTazRiBc
+LfqxItE0kMO1kbuk2dTwiks3qolSKjEsCmZqQc9XNcpiRKdInyDu722wgWUHzYq
jzII7NgHrn9qY3CQ+mBvkoFqiMDY3iBFNonDa1LRmC+b01syyOEy2/mFKgMxVHh/
LE5DY+dk6l1VHRBOw8N9TG4BKfFAdG955P8Cte4GZ1N8HtPgp4ZXiwqVkolBOUNH
kmnq9HAcn5/2Cv1EhXfefByBBpzMVf9t54H/RjGzRPmvnAg0hqIURY9Ih10/z7yb
KYHTlPBJzgiX1+NOPaEbwi2GbTdeKjqezKD0TWEkxwCy9Q0NwrCEmsRn8asHtaTO
HMeVCzDRsMPwM8b/Xa5qVtvHfUINbF6958alDz8fff5KdjERw7hxipjfm63JF0+G
7XyB3sbJWk9zXBxy7GxQqLqF+zZu7Ye1vHn6TSgN+orooRJ9YbHb8Z8/q0Z7vASE
m8gp83SnI9wsgf4WyW2pRwVBEKRaELIQPzNerlpYQI9qo5SmGVkbcQl1gUYIakgH
/XO7MAwbA77u0sSUsTzlgnHrgIZdmbpzkymnaaV03N00uKEQezDHwOCWVq40KYGO
sa+bf6NE0PXzyFKg2b0iHzX2JUPp25xvTmUlBXWAsI7UV1ak02JXeH2gezFYlSW2
mqw8kcMhzSqhPwS4ylV/50wIdr+7oG30hk9u8vAYM+0OE1/oYrikKJL4GET/GdiZ
C6J6/Lzi5i9J4nIAStR38IrP1LPol1bviwGgofOFB9fwcec4QRy/5tqJ4HFI/x22
Zjt/3mhByF8e16S/clU2oDWmxM4Kb6bQeuAq5138ka70xTS6M366Qr/v1J/UdwOQ
eIwZHBNDpZT+HVuI7v60vw9dWpSs6L6FqdMK9guTNliDSfo7FBRGHCiMNSVH2Iup
5nhVxkaCH26VGvAYYMsMa+SPDmaNWDDQoPXLbYXOAewK14M+EZpRZ5L1b1OUYBav
lxzSX/3Mec743dXDWhORRp+mrCVNaf8b3YbnWX/LJruz1zDlMt50q/jnlxRiGHCq
FNxOWrav0K3bj+tn9sJWSymbk/6Sz1hm4183HiUuZhJlMSiF2WGpb0bPt81u+Dca
Bb6bUJmtVVnWHq1t5gZa9RgAIoAhDIEj3Ss41vI8S/PsTJEzk2XRHWmsaMuhKnPb
w58r52F6C6XkvqQpG3VvZ5KhpGFnxLatoa4lqzXztyFBENr5RVJThNLqjReSamUU
Odbp1FZpV+AXspdl1tFFT35zgzHkov9umFWp4eSPwnbENRJMo4BDnu9jVkzYTwox
fuJGc90I9bg9CafY0dK8sOjv3mXk6nKw5iecDfbEpMtzjT2go9heCZRpZPkXfvlJ
JKuw1hKdOzOPg+YUyo4VD2uYHA4z1E0uCFdTFHLCaHd61ITLxQSIvqMDFL38a1Ti
rOp38ZSdOcm3tOWajB3Zxax1Ut86UgewI5zF1dN1pwpM3ltg0iy4xdM7lMvLwUGY
LFAj6PkfRm8XqNhOu7SxJaQr3UxQk+GipV3yRRXLFCaTzvZgt/N4Z3lyDKw5Il3A
esiFEnwI5DjUgR9bALy82V4lrJx7lwfhzemZAIaKwV22mgzkkhCHliOWCvEc62d0
IWbF1rllstxHirIiX9UggGbJb8xGkodcxN+h9IpnE51YqCXk9CkJgogMq0CGYqly
YC/Y4IPZr4ScW7jxPHlNA2LfIMcQ7/azYeaL/UwGyRUIQ+Qph4lkf/XDFi8pnTDi
kt4LRIa22lhnvAT1CXCQ5PE3KkQLTaLq4Dix6WBnvA/B8nrcFbuXsb9BjWW73P7g
7am+jpT68HmEcO9LsD9kDMz1p9YU8GMotBiU/ORUrUjpZgJOB/G2Fid8kJoEICYs
YaQuIP9O/iaaWxvA837B7erPADnTW9fsW4qT5IXbUDu5zb9TEnyGTEsfUIr8gB2o
PIKTg2v9TaCHbJRvVCcLy14wMvwTcye4dmjqyyF7eJFwdl4FMW7x2QTOneb7pMwQ
LveZzKI+juh0KCUjoc2xEs3pK87POmAXc8ZRk/r/9sg4dRz4VI09bCiiKGSICiz4
TtzX9Y8IxHrFymj5vDLFGGq8VNe6U/AyyLNPH211TH4yc/fQR4n0F+B3J6+qeBiB
GlzcglZf2pxKCXnETf2utsMVUlzxiFBEpJSBIEtz944iwjYFvz1DLPF55QyPV63+
N73qqEFU/KfbwDzt84tdAvA2LE6svN3nALQxdDea5T1k3vV8xQCH3eR2m9KaCMwa
ewOlfWLafmQoyR2MRIXjZBMzTYLzHouHj9+bpcRlau6Fn/AoWa7Eh5UecvG2z+Dy
ajEbtM4W4fPHz9TmGfzAMo+5T7JQX5SxrLMyK+/fSCDwzH0gLF4WcgJt9pd0Lklt
M/1otJzvl3Bg6igsCEK9URtoxnOpRF80B07wC/P72Nu4fGhFRHw1vi9jBJriauY1
y2Ok60Kh/gCDT5/AeZgVT7j3jIrG46ahMPld783eIrgC+DNsA8JabgHgCfkbk2uQ
13T+72FumaxXm57hmbwjuwyO35ySUJHuGCYPddOXAtkw3RtwHP57VEzdU3ew3frN
tEal02tKPeO0Hp6B/Io49PybC45zEIJFJgjz46B+nOh0FTb06YuR4FjdCEwG+RG8
iM8HLMkHYbz0JYY0FLAkbhlukkkEoM7pPNY3t3h16eQJjylDcStihWp8vxVbPqvh
YSLi9DA4rd3oO70SRcM/Pg9Ls0uVBbQaXDWbQeldjjbmwb2iNG1rq5p4Nt7CtIwQ
+epqUtcDAngU6oPayC6sU0lewnGHKUp7yThXGufWBFtz2zQl/bER9eOGgZUOy8pT
6f1bxdOWE/ezH1i1OH5ZX3KkIYAMwWYGCb/+EHyudUvMXplFEsvS2pvWV8wD6uHp
ZxRsNCpb9gn7q3w7S3AMWwyg0y13G/GPM0UCAdwq/+rBwYeZP8TNagJpIycq7WaB
`protect end_protected