`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6912 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
XVHVS6SW8Hb+XzH/poMIoEPHiOErKkZy5ZA8/8T242nx9tQTGnir1xsFqxBE8FzY
ZscnA4RGw9c4xwMZmD6vQH2oDraipapv0rGCca2zAdG5LB3ql5M3zff/gaqbKRpo
iUNhSZgBo0yA7WijKLJS0Od9ZsdlGg1Clkifbujloh4M1M9uNGy6XPkGNRn1Pj6r
uER7kiZgwZHByaBzybE5kJQE3ug38tZFT+PmtTNW4m5+j4fwfcO/eiHKsRRNPmOZ
AlZjV7lC9PIOliQO2p4a4K55b2zPQ15Ml2drIOj3sGnpEhYIAezfQbsfavbeRInE
uMZOlBipOcwHzf15gjPYy8+DXwU0gQzGyOFFfmCoQu7/cPCF0SmEY3vh3sVHDghh
r5xGO2E73Bil86VcROt+n+eu0TNku+6wUhsJpi1eeafC6FvRqWQJCvgNayoYwsGw
2JW3EUqtsyuROhhaHY2FHwa/K/Slcy0GglOGTe+4Ypc6DBFulu2yI24Y1R648Amo
YspxOtTDh4EmR6EL8ZqIeuZdvqQNYcD1kGvR9WpBio4IlYuA+efLA7CN+J7V0LCO
qOOsF3ElPOCYCxpm1dQYirRzXDS7pG52tvYwgMWgy6IzmyI3Kzz0rT2khrEfiNSJ
uhn77QLMtF5ocziMtgZtp+Fmjy8uiXvmgomwu4mKAHZejOZEWOUsH4VCVxBkM08b
S0w+0QFhJ0ll3i3wdNUX7+94bc7neAdx7oC41DscYqqxTr6gbEkNYQHZe1N5xriO
NHc/fLW32XT98GDiwmf251HtCGN16pNmSIh83C0FlQ6bZfq/ZmfPKUGSgBYgcUlk
YoVzJNY1FScb00C/yPnK4hj6aVa5Mj7BEZaI7RWQvvO9ghplUzyZmKx1Et7nIHO0
OTHqzuUAYyQgPTmmw2VVXZUXZYWOVoU0zMMSxZZozoGqej2qDa/duTduxcPAFQGv
7UZdzgMwP4Eql+0OvE/ZBBy8p3g8GC9YgLPVe3mksQxGRPvickvqgvQMPUUBRds3
I2+wNOqSaBEtkZQht2kGdbC5MmAtFzq7Yh97c8tfq/wglXiE+G8HpzGKHiZMJ9xL
cEZnTW1TKrjJykUisoBNHROLHUcI1LFTe0ukd9nQWhJfXsMK7i9nqwS92FF/SMNX
gPpf/D48KSV7CaATDuzcyrESznXG9kz8YYP3umYVonFetL9oYhKZYpzD7yDVEv0M
ybgPA8xmiyLMvaf6yvsVK1mK5zcC+ad3zpWimIgKtRebeRJghX91KusbA/UkmFN4
q/jyGU9DELUij7W5sEf18ACSLV7TXXtWPV+nKXsNu7ZTPW8EFwtCxMXEdopPEKsV
+SWWzFGhVd3BArd3WVOCBZpSh6ZwdZEGbx+eSGMn9y25p9HWamMCm8wjfxHpfNTJ
XehzkTaWDHvX/btLulVOxPz9ALGL5QqRMVDokl+6BI40aerq9E6NN4zcgHii1Awi
5k5yo0tasePhriVTHWBbDg08iHY6lPngR8zvmnc8JWQzuXwGHxE69mSR8lwxtkmL
V6DTucx+liMnKEqdzs9GvIwWmG9MZzOLhnXAtAGeyrVGxvhw0lJEzhUl4aoDcv2s
i3iR+6Mhg++2jsfA9oUkaNWFNs8BSAbUQxC/3ragyQUK3v+7eNh5rZ11VuWC2OHf
+aHHXLr8tkcdlNXMQlqf+W0vKCDFvQNayxKidIw4BF/qy2smYow93D2e7gTkPM32
jK8oMXaI2WgtYqaeG9T1yX+3Go3KAGv02aONlSl0L2GlGRKj6/eCJqQ6O7qZsEIy
bABEJoBUYhhDBHSlOCX7G6CJHsFeVJ3AzguDzJejjIYCV5BCvGCEMAiGN4vq7qtM
236FuLHogMDwcce4Qp0f2UsqoZ+YZGbU841CkXbuudgOgPUmS/mEA2cNiPmOseLq
D44Rq+WG/m3yqQdk7n5vmDF6zuIshOkcH0+DPTT74jJJoCcpk/HiXFYLyPWHlk+i
XybQ+qPz3CLorRvltxjSx5oSFxJhviK9GQWs3xQU5HpUx7OJ60eREbK2NgbqQ2J8
WFYONjkNZPZlhXB0u7acfGznRVSlBtGu7rAwm5sZkmzFhbgDRkEhwhqi5qBOrNTh
Y19lIhmfVtVhZDqGaslufg1X3MM8H8pYz+0FoICa/x/O+Z9pWUw+PThOmniMKF96
MeQi79Y6gn+yUoPMA+T0aaTw/qjo8iNrv3fykOowIBMbY79TqC/CAsWxMU4oRB8/
AM7wEH+MEQEYD1+dDSOz192w6BrZ+uIu16qvE4dmjhK1r2u0Enm5rwlmbWTqBIPE
qJIUgceoon6AqlFUqO/zLODUf/VQeVpJPIUVBT6xvQAAlw/6rPdfdqObW0nJA4Mo
ew2u8kXMamR8FtsFSqQBP/Cez0ziqeluVBES90QzyAUzFCTY/PhT816s5ZSRo0/p
dX6hpDEf+GpVSTcUdNMOzqc06uygIeJW8bOWoKVqg0JZ5XtCd6Adplh+YTt5+x6I
nV72P2NPiHcB/DlKRbMD17ewLYgDemh1VVTBvUMFvGixCRvjwJoikxAb8vrxdz+M
NpSI24RJfnZa7pXnnt4tZ/QhIW5UUamCoVnfCJ1dF7f4R5oA/RMn+jBZJIMvmShG
Ff8GIld0Ph3LwQ+Fzgy0Z3/Q1szv2L9l+qezAfulWCyWkgmDRATDRcg8bWXL9pfY
LkW4Txoh6BHgMhfTbPKxKz29OMA1teUUqTw9CUUslAsZGPKLXCIz6PH84cw6uAXR
mWUFHjpUvBuBU38UBSqCXFzKRlN8FBvofkVB3hKVQQ8v6qIzyeg39DGIr2tBWJZJ
GPCajxU5GOrLb3PY3K/nqfEPrUurlO3i/E/2K4EVO9A2pG1fjKEFY96lC4/ZHsn6
S3xhxHMapYY+Zwd26vOMMdSXFtIJi/oQmEQpPypkfWfsq/Xw0sxPrSMsi8SZSd4N
QWaeOSV1vn0dTWlPjwERa/8vDSNpn8NVYDmHHqasuBf8Tg8Ky10akx+S4PaVDilE
L7wa8qDob5FmMfX3Nq/3r6tTBASpMNr8FgnmWhqkIp+0RMwcC5S7VapT2l0VOa+F
+As8I7kInIliKF4Xnc0LVWj8nUIxzBalyD217OWurZdA/pm/Vbb5h5j2w/SWOzCb
b6c1cfVNNiWcABY/cLuxyAaoIUV0f82vGdEqrIh0eQXK0SN9n7EpL4fd0HeWv7x3
bK1PZAi7dajfjYp/pzEV2P77QXdwmX4VdDRR81UgFaA63pzMnP6nxeiRSW20m/9R
HzYEt6LVx2/9clr+ayD96XKiLohglQY0zv8PVk1T6BhMzGkZ2tZYmxFhdVR0wO0g
Tb3YdsM7nxLvXLR61iBI75cfVrupaaTL4OENq3tUhDEA1rWj3R26E3+bY8laj26H
kFVZvTEbUlA5zEfryIn0fROg+W3UTgEwhTgCsEdgjTN0M1VqEXTFtv8yK/aePdPw
3AWUekOu2lhYxiR97fPfBTYM43JS/xTLrFKf8SIlQbaZRchUJ8PXlsnxd1+pBr77
fZqaQIkBZCvjIcBR7X/gq5xEwx3JiJpWFZbP9eWitIU5qhwqm+Qx1RSl8jNLokCn
lvLoNELImLN45iwyksM2peVqyiW6gEb8GDsGX9fx68teywz/2LDt7bDpb2pqySZh
9i7FOpO3/5d5VW8S19Q5ZioOg3XM+yPj4efDF7dAhLOdBTX3ZJdJ/QLEyvDeTqtR
SO/qR6EWRxkpQOuL+kuXg4G41VwaqhYEpfVBA340jHDm3X570wihLvfKOyk0wqOy
Edjclpal2jhzOer17CzXIIwJUOt1NnNLVtANalhxPyK6pp39w/FHSt49WuFTZi12
gZtc6YcqLzzvrT6R59OJtRDqoX0RVd+/mSP3h9o1h6RFP61wnHDPi0FiebIKusI5
e8O+sCPY2/78fnNDbO8q0cFoCu2RyV6G3vOm+AT+fPbTTupJNhSXKIq820hR7KA9
xNAPAEnI+BnEAEpp+Bi+iQ8m1L+ISNDQFPSlzSVCaKURFixWK1wRnM7rMJIcWqTz
xX/zlfarb+euOOWxz7TIR1H7P9pZoRXJoaNXalslbjRrrPjLwkUSYsqq5g5W8Vun
ZGFsBAu9EZJ4Bepb16xv6cf+VWWVe21pkftYDLIerqmPbpjhGxjNCPrUeJMOA7Mt
hvnyZ/GABqVd15fG4K/cnKdvch/2uSQMiaoyJr17HcE+3RJWRTvFEuKTSN31LIv7
wI7AlWPwzeBq9Wjl1Z6K6w7o24dIjwtKw0DTKI9OLEgZIQvaa0E3XWvU4DYdn5IE
eMwIEQXW+STW9TsrFXcT84V6FlL4glrodZ9SAS6/rYjK33RTm2hlpf+eUXXHB5hy
gPgBx90AzavapvZ7bKyfr1WioT1cezjjWYkNcLzvgEltgzO/N/CCEjn3RXY5ZwxV
8NfqcGYVW7uMXEtZw51vN5GmWVLm/LtofPzsVkS7UhKspHa3TjzLFQzx06D+l6GQ
ru7PIgcA7H4irS+5T9PZxfWqbxhF5D6YfDbSfEzGTRtJx2kq9xrvb6QO/FXU9OXd
iuMcvrVWFIbbK898Hr1mJ0eBkrbMKLiW6sFME+88bmWUlYxcXeAaw0I6eqvKOQVL
jEzFiW+lC71ERnsSIpH9u80ApkJPVnWFWo8wkrls76dMoZ9Zkw+FA1chkoO1AGzM
vqwJVq/4UtC3Gq+uP3utV3F69iFAA2egKSracOH0KkqHfR7NrgCQTmmuwcf6FgSA
E9T0Q8BSsBur8pl8ycgOR+1Vtc+XMnqcIHTUj7czNfdrqTcCT+PNV+tp191MSJeF
6xjHkb60ZmBREdkHRKBHU+LP7+zTTROOv6MnvfEQW90ASr3rv9o3GFd/rCJGzMhU
y/PkPJaJ5+WNRNZs4/UPxh4eUgg6MNPCO1eZ508f6JvCTAg9OeQlk1513Zut9yS6
pyBzMeRtqvAxSqst+VArzf4T5l4dEwrP4EvZ4jv2rDloJVKn1LjQvZSgC5e/yWxu
Vm54MuqZMJq0CJ4niyZXjfmR8Qbgvjgt4EOJF987efwllPrRrCVcPZ9eg2oORlRM
mVq48+cQL6o3x/GiSp7Mfi5hlvuCHR4/sQbxLue+VzTSb737DT8T06Rfs83ymvqA
h017r6/OzRCez7qI2LNHnuJgSrXg1s5N4K0R7zkJwuQ3RzMdQLACmOMGgvBa5iOM
u2MwzhsfveooSpwVnSWjS2PXqy1fkjn+NtdtfeyhjqhXEPVjQ8Uh+77gcsO79uAt
bBHQpOY0TG9BjYn1b8Lppk9BZpSlzQfusNtQIDc2ga1AIekIWd/bmNdQ6CKzCWtf
kDSm1s4K8FS9l5dcshUDuJKav2E+GKpgi6GXxIPlF4mLWKizVgSM2OnLwruAw35Y
pXVRCXyDXyCz0rZM3sNGeTTxcjhYt3trpzG9TtKCPH50dBnZDSgZRLeFAuhtIsMS
cFC7ivbhCmif0Y6p3T1dGNVIMFaid2gK84ogShSRiLD/FKlK/RHCDf3D3e+69h5y
IyeVjiKRPRNt7dX6cPe5/99BLhzN+v8n5CD1EciLfOIyPzQxUPKs3yineZp0B6bj
v7wdb3reeGGZAQ/oMjUEUES4+2jbAqAWjXJdWt6iocTTkqOOWgD/0bPmiLeeI6OM
FeMkCtNG4hna46GED2KVWu86Nc6OSIPy49soqCWGyqltmiqIyczG2dLc0rP/tBjW
0/pb4HOK4ivI962YapN94TRz0Aj7o/RsQldJGLh+CUItWzi34Xv6DdN3z8VODfkE
TP1GWyLALEPOaYlL6I5T9hnFHmCk62nbWw84sCGTKOoQ1D3H0pDmmGV9YBu6BinN
4yNAXfnqyV4QjyS8OerQK+vvaaGV3r/+Zyr23Ey9mbs5b4u9Umjk9z6k4BnkomOI
qCAJH5edo86U7rC6hbj9XiMHE3zRl/FJWGyHUnhRNximSwRRe86TqWL5qbQ3/mla
73kY7QWTY7Gq2XbUTti1CuiIYgKfaNtGAphlJR7GGPPTmQ6f+1yVNxxU4DxqUgpi
Ty0mfwEBMYr66X+tk9PhxQaq4mO9ms0kXRxGoZMhfWABhXypaGti6UDgK3wbag4G
HxBTmxaCq79hsNeLXY8kL3P6PWL2HoCJPw+cMeiElzefo0OqwmrydOgeKZPOlXaP
KRGbX5wo2bEeBrjtoTSCi5ql+TdGQKFcwp1eIPCRGNuAGcbQjzV7k3tuKDV3+cVQ
GBt69XBWoXrmslAkozM1a5Y4qyzWQLfSG0puGaWBw421n0RJxHloVVs4enEZRLCA
qu2f46z7yINtqTCWIrnz33l7Kp8qogsxovblIqeshspDwMrBaBwwlphcVZR66e11
fNUH+W1uNed1oV0nLk/O8yRKAcTGBbUZh6fovUbSDQYMQywBQTTJ373DVFu+T6Mj
7TKpbEc9zOst6SfedB8bG9f4maT5ZsMLyjJHZuZmBvfag/X0WaYq6lZeAcAXjYn6
cUqjRoVJU5wZgloLSWizNaEg1BSGUlL38pajym+LHhlrLQjAXtz+dBatUbDqpo6p
AAqITjWlBVBSktv7YQ5eZUGvsZJrGrB0Usy5Y8rFKDkk3HbCzYSDTmfNW0kGeGWI
/mlZrKDVgpW1CtANF1qAP2ijpbQdAwaUIJ13QIHYrtA7b01bQcEcBqVsl3vYCj/j
N0rvTuK6WTV4V5kBWUHUTCud/ejAd83a+XjTb90Ljys4W71TsQ7l7st3YhP3A1oj
oXMoK39GSEDn2r6TG2oxniRdEOjO8aDYQI6BJw79NeQqqcnlbfQTwdXOpAGvBYVq
zb6tgi+LhWksDOFJS1AWksbqVVvwof5pn1bLVoBR+05Z4ThUSXPWUECIm7Aiy6uN
IsN1Mx1UML14976g9rMrm9OP6Mv80zSiFaWm6aJaOYfHWoPKT078pcyhW4WiBCYB
fC6LqQdKd8PcEQFxhnd2xNhdZhTZii1kB64dSITLbQNm1XpDfrj35cPk9gPw0mhF
r9Cbi9r4BQqSj/nL6e6pJKCPJ3C8/7/wrETYfaRvSGRMg7g8KyHsZcZ3yZQ5dHZU
9qk8KesVJF6skUdC7/tWIDZxO34g5AmsQg/KMWzFNA/cznqC+nIPujt3+i31BjPJ
sHqMKP233hrRM9YdMGZOFKt6FmbzdZP9vhVj2x9+TnTPOsaXa8V6E2TyKS4QnWso
KWsVRhXqEvUaHeaN26h61kDStevYPAvAN6hGy0D26sR6ClhoE4Q8a+eKg4lcb4jP
y2hUFIwdI1PyR8ky6xyYNm6844NbNodE2MtUtOb9uAOMb9G8lImIp6OgJb/XW/Bo
WGib8YtvP/LfzzswdElvaFF2QTVPP8/tz5dZ4lyw+/ybyWnDYq83lCKOyXgJigUx
3sfu4RbZl6BbP5stwifEuHdEF7PpNTvAeBl/ZPIXc2YD6Hckat/AFCPe+6M3F1fd
5a+HEr2jcr8BhrOCEmbW2vAkkzEjWXMgFF0HlNiHXoZ7Ie1yWL88ttkpJqyKybGM
eRfgYcIM0pS/1FUIiPFAPXPtTsE82SW8lOKcGOdP7FLy9ExEEsLajwuVq1qrytWJ
ceOnGA/3TnukjLRkgef3B3uAm5mnar2w0LYzKkECMqUsjA7urjA0wNu1zve9Ej9E
FiWDbpVqbx8Hkmo0JQZeRH4TUZkYMTrxEuBZWApghg9Lc2F8NO1UuZ8PupUDuY7C
uMrBdz0pv5Eq5V9XJVniW/XOCv9sBiGeRt9whjeN/Xt7J/6frYxYdhgtDg6CnuNe
wM+A5EdyDR/0bDVNZcFPS/8hkt2iiTmEwKJJmelep1HUMnDZgZeP8hHM6pgKCmj8
pPf5uxzHiIwpuGlypgH03nEaEJxS00LYsjo8AGF5PHdkEW5oA+3ds9GzY6r/GHKR
JF4APqk7d/DWkLEoE8skWRcfexW/FFFyAJSV8H3fwjzYSMsYLD8A8WZMU/XiT9OX
1JppPJlL2vCEXjmmjDjWS+mYKyIw1P/GNryI0VugXfv+bZPpCpLikVp0glVGVBbQ
CLTu2w76oaojCCxQGWAFIFQyw+xbcMtDBqwRGqSMUFb6zF5iXM4XOaxGSirdsaJm
Xx62Ix+USG1gYihEbQvX/L9r3gfsmExMqenQGwAS6bYFQyq5Cz9vQpuMs2Awbeyy
NTRTGr6jn9gMusbGUI8RgyHexGaYtfFDRrYWmY3ItXBAgjZ9vRXoGkA1flwavKYY
Do+Y+AJjJ9wv9kBr6q9HWJUO666qV9hBAovTY4xK7KQW4Y+Qg29LP5EGJmfhPX68
BFtYnF57Umhrss82htw6EcYd8nvIyR6OUaow+8y3a1j2//jp4whU27c5JgHzWaCo
TDS8gr7IT475WobLxrGUbLVIF4CZxGAy+uOXFqIZxIp00tYhB7Lr6syS2gFsLdiL
lVD1dwDlQ0WFFpfKg15TxszZaxun3sNp3AZ8AOscnMjOGNICU19eECX5DMoKp2en
yYpwMnOGDWv+LWSntqbG3MdS3AxTUSizNfYJh9gFpKMm+NoOJR99OJCYvwWEh711
1CA3JIVKcXLjrgTGVMmBROAfB+sGOglPjdOxF5nqDgjxkurojl4aC96Ycq9GRh15
LfFd1LDI9lj3huY5gsl1T4WC3aJ1VejgveK/GrjQQjhsI5XbLZjVWlyIxqVPUywm
+adfVG2A+mZsgc+NHdhKRI5aesWQdXUh1yFKaGViYLz7ZHLEN2pZblWkH8WUumP6
meIu+czk2HWk6gXcKEtWBTqheZ9FzCaxJpm++1LgCUJ+eP+6lB/8kzj+iz23853i
Uetqai3vwdR+vzsuF0aQw+flEl2DSJClk2ejltCt04yIo01InLZnrU6QVJ6WnKzY
Nso/tuQRTY/fsgRXM8BLP9nwCe1/a+0z45OfIi4wRiUPSuDIz4yVGvIJpypVHMpR
9SLlPbyAOcyuHcqRhmGKJ0wPT1vl8/UuANNW58mHtk6qYGS/iEsqMOuwLoqym+SZ
VTGBcxo/+55oAGS/q4CpH7eHul4wG3zbfBSZPRZppAZP6s2NmM8PmAb758acXwEC
LJoMrdnKGTlBFGw1Ay8FgX6SoAe4bqiQta1f6fubHDXPMp8zRLwDtHx+N3GGZrJ3
`protect end_protected