`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 21376 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0gQgIG1mJzulW1XOK5NnZR8
C8XqDUtXW7uOWTnSVqbIblwOHrDC/GFb3kYl7b/cVSRF+w81Th0ZOVRGVCrlYzDv
lB/0AU8lZ0GB1kTTilxo8KhEB8HKVtgGTX+fS+A8JqH2vDLYLSJ5C7a4EAY/1xZW
/yQHESfMDZ2ZUUNge6GtwMPfDU5YjP0n0EbetX70UoDP9OydkDjWviG9dejwasc3
J2WcmDD+51fnHVf5EmGAmLv2yVYc1LLcKsiONrMO8deXNxCn7ao1Fq+jqi97uA8W
cnuKZEiJ9Nvhr6L3S7xtZ0ehXUxBKdxG4B5OeCUIcMPNEs1g4vhonLEXCdM0wW9A
Jrk/14qTUH5y6lKOWztU8lnSmZw4laq7j/KU6NnA7XegUvRygNHsg8KCpqynA8L+
KtSSXjZ2jIAJCatCPhTCPOG9bEUnMvyI1MF2pRGw/bU1UtE8P4mar3Y7Bh1b0OCp
l1F9s2+BjOAEiMjG3gLiWBsoJbdALdhBmoX2mNeQftVLqACx6JrwXT6CsFjLxbkK
EuGWLC0W42hRIhm8XbEdCyfRSIXFsjxEu7UVOLUMKCDbFHKUujQdHHozowEYzm23
1Yx83/fIkD8PkPBrgCZDw0X9DkFKcC9kq7DVEFXh6VLH9XvQzuy1IMyFS3q1tQ4n
CHnFP6nbmnO5fYgiIDUjLYsUjKIZJ0ClSyF5Edi1UZsQ3VNQkeVdlksxRJuu4/6z
IV8RaJrycJdOrAA3vvL1JuuEkDc9BJ5dqLNhwBTP3E0jeoOGDI30f63MozGKUzi4
gL77+nOr0cZPVWU9oKT4obxedJWqwVYFVEP8RIa7A88Qgwr8+qbpTom5NboDCEJT
BQwF98ZPQizvQzQiTjWXsGWp/wV7v62BaQ9GMSTDlkreB0zYXBnxhGNReTbansf7
eVJdb6/aBu/1hMRHsiyY8kRacPoyTiWS33EePZNbnH87YWJS/WBe/qNX+Rktpila
yOAcpAUWuwYUD72gmyuk8tqCY/+OeZdZ5BYb+4bce0oZnp5lkSHRdqTPfFZHCq9x
Si4T6BhId2v2mSVADT7IBm7oen5aLsfMb7RDObLALFp7BOcDytdftHQ8V1gie4k2
f/iL/yBB/K8Lq6kEC9OMUeXAR9++oun/if8gszbCicD1UNJacX3hDzGcF6YQo05v
c1NzVvb7ksHxID6fADj4osM8hh96vRj6Nkbhg8+RzTFg/an3hjKHxeEvjx35n2HK
taWGkoUbQYnksIJF9Qg6Rt95B01GqQi3spWGJCLxViFwuvQC4XQYwHYpb9maLXw1
cAp43w5zSMEc7Qy4wrTEeGBjCuG8HH+9XYa9wgTiOuSGdy8gyZOubfK2s/nqEa0q
zrXmCkY++uGNIFSGiRh5H5B6Qfm+uDn9Urj0GIFQg20Z8os+OTPaBgWK+M6lE8Rq
8w7ofpYUzkteWXqZNcp74XnBDcM0t/cuVK3TB2EpM0x++rWUONqOiNJV/CGomZEQ
2LwRkQlBmEZu9OZBtFFgy/OH7Tvhy/SAg6yKc5lUuHoHygSN9oVzT13q0J/WZccG
FZoZOLWwqu7uVxU9+JTLziD2cPgDeL1BOv7hyAtqneY0qSTtv+sgbUO931Ov87fM
cvigKLEFhougKz3bD62yLnMktB/GK+Q98zX3bpwQrVnoOV03Wkh9o4/0g4WJcJni
DmBftwX/ZCPZdTVRSmoDJh6tAmboVXLhqcLdbh3H22VuH/xqK6bo/IaKBDrjbG6w
8ZATguJ8s6uhFfSc4DMyx4yZWpfPgOLTeKiMVgHuN1d07KTdPpCtPrA/2J75zMOU
IW1SdlOflkbp3tjnfyURn9X10Buf8zM6qeSF2XJb/6WAO/yvsyF0WnnmdmN56TBG
yY82FmLaewTAvKbVg6oonQvbe19gap1hAqrXQqxihOd19X15oS8Hb39aJk+xkrTB
+Q5gbz837a88f0LcBBm1fJ9QcY0qJs620aUctNL4eb8GYo0HYzCYhiEyQSAHPUS6
Lp7G809bXN3k9yUziFwvZvWDIG5n6DW4M196lJVaY9DMUIKiT/538h+D9QMvHRYH
tqOtpg8utNRJIhhjKkxAB763lmxZPgLIFIy3XQq/KhnWalOpI+d4Py+9i4YKuLZe
92A5s3Yqk76ucjpGb7rfCQwtYed6rMJAXbxphtwhmca3Ri69PGT+G/AEvItsd0VP
1bH0slZqFU7KPLeBr+nF5k1ss6IXZbd9R+ydnbp/UWpyGHbRi16mixS7g+49lyQN
BrDfaL635LwMZjMOom5+qTZZ3UGb5ZD8jjdF/oCSP5ETgh1YtN6ykmJxHzNHn5e8
ydqgeBAYbIAKIZjX641e8yb41w08l/EplZ+y0UeB9uKz1CLh0gsRq6SR8Pr2F7AA
FVIj8t/rw/jTyl7ynv6tkDKBkUuIDjWFUibdJekvL74+ARi9TOxxfRqPk8JO2tPL
XnoivWeqoMBtoTgP6FsFielYc+SljgRAXeHaO3TH6AklbM0NNmCgrf2xs0j1Mld8
XJuMfeF1aRlH+3NecrRBvKlscpNZSwoMQ4QIGv3kB1SdhM2yhCbaT9yRCoRzZW+a
BfC998zhSiFWOrYZCkNx6C4ULMGQXGAyCE9ipj7rgi/oK9u7jUD+4+My9x2tFQ1l
DNUGA8nHoASa8g83BQZczfv85GP4kfaw2F5B18wE0H6+cJQpYvxT7RQQlF7nzmvK
yPGkitYV4bhDqaAsCzSOGeYlCPbL2Ifgjg0vGYpKwmPvn/KBGrtYtKvAfbGa1vdl
opNuSRzNO4QWV5YjyaeZAlDbf8GLZupMKH+XI9mFmFThPqpLfKH1zKtNi+rlZNDc
aBa2HD2q3pyeJGvdE2b5PWaw22hheErt6xU7uOGaO3HPyCX54m7WDyQL6Xm/oc2I
SuO19W5dOIcsKc3tZD1mbh7PrjgPzpKj0i+y/JMrxe/ggGHochi67SGkGXnS6Y5t
yzG9cTdRLhSzSo5cvX2omigBL10seJ5elhG4bZtqFPW0qNxdmb6dIMv7OJEdzASP
gZzGtFx8GEZErjjOkz2TxQqkHNLUIlx+HyPuHUqkH44r72uXt6c6Tyfv9uiyO5Ys
787PKDq7SMusVx9H4g5ziBiUOh0s4Yrsd2t0XLHvI4fJ3aatahVVU6ACFk6cP2Ls
nsVlZygX9jAE6yBPvpCSJjMvDZxZmPr4DCbCzxoBMmLKLKZCqWFUQFJaJifm5ySX
x54GSW/I2HijBEqdqU9wok/lKm66o1sKDbx/uaMlfa8avkk3OfGHfejETeMyRsds
E/+/PzPkfwKa8DqyW7BpzoZ2dZEjSf+s3AFZEqLQ3WLYwglnTFbRYFx+gGLgakN1
bzpZikFGd1ipMVcCb4LMC36Q2bOQmMAhiObaaLgdUw/4Y0bzH4rWA1NNVWCcwYAe
PGPLhjV8/arrLdAdBqOcv1hN1gXGedkL2VyXLvj8tmH07R0UYEV8wAe83f87i5Cz
adNcgux/utHnrU+8P5ByUijMZtGyCRIZbTQ75VpqVLrqFpsG8gPuJednNQsHYXYN
viUQWLyG26C482tDIpYVaO61qX0WSKlfo8AVbCdI5DxKCHAtV0kP9aYmieIc5kq4
3JID88fHZZUdgbEabvu5KmJzE3k6yI5+BcptxZnAqEn27zVxM02bHe7yFVj/posJ
srkYJf4UTmdwXssGNL8MEu2LAFFe775OF6dpRG76vCvDUoG8hvmD5l/QdoEZ2HvM
dt9ofGQ6hKZSFhv+he8zfhMbumis+ByCKF8W6p3Gofbb+2C1e+I3l4JGqtziGKPV
nJQGzF0+GlpBAtA5gcEkXchlt4ZjzWpgz1aCT+osFT9dgPZX9AS5sK+MfBq2o40Q
QUGltQ4UGeqMhORwk07jf9awDeVqFDrpMAQpeCHJn/MnJfcIRAQs023VkAwrJcpC
ef5YxRMCke9bopUNhP77bypRhH0BN08eI2Chj5aDnbo+ZUbgJU8TPJ4E/UfPRmHk
KmTk5NIn9NQi+g1JdnXUW5QW1WC+eN3/kdQOKH2178HHVuHmU0S2vYYTJP+pgBhw
HPmfBCgjxGq1OeZWAkwYNojqKrKDMClBPwm4TUT3OLH1x0XpAObtMuj5A2t3jPcb
UJJnzjmqvgggRRZNxLY28an2diY7mHKJ33w1ezkH/Qy0B1j4ZxbYg8gut/lYJLxr
cIJAfYGDpoxAWhuZCzCb/j7rYjFzrJ735w/N6zI5e5wwDML+4BID2pjdaQ5RTW0n
7FS/dlcGH1VNCETK7XuDlLnIs5nFRFMJub+wjaxeKN2iF4hF1zmripk9v1UjAiPp
fWDUorYDTr1nOBtnXTeFMBjyAT7IBHmoPt59ZJecR5OUWsHjogpKrpMHmj5iNXgY
NCN2lGNRPv9mgg4wmxD75/S+N3nS4AhoWvuTc8wvnRW0efogJ0MEDjf47d4MiYdE
r4dodII/kNx6W3NripH4NOeDu2uwrWNGoEEMHx5R+1N9p0/vo+FcFPmMnliY4OTZ
Y04e6wxJWy1O2RNO0J+OzPXN1CcJNpYgeueVqR79iC6t5KUKYsiDWMUya7I44bCC
033Mc3rE8dy9SFauoNNdPw2C92FJKPKMNid1sMSWAtZVORvFBYe1CFkaiIk1ex0t
FhaHpCb00+ukPdPIW6H8I27U9pmb5Wnr6Oi/+uKZdMTVMOAUpjJuft53ESmTbuZT
OKYfaxrcpEcjtywh0QMi8bNrkuZYADskAG8tTtpnDbC9tMHN69r86Fm0Lklst8RI
Ppxp5uMD1OjFZD/b1AnqdQ7NuwoRMRS/7izBFaoaNdVXFOK0r0JLtcDTh2c8CrW/
GVvHzirZgNGjXae65SzesJVvP+YR5sa5X2dVlE+wvIh1oglLW769hNy4op8xpYTb
lsdtmOqm3ldo3LZEV+yVpDrBGuI2DlpgdKevdqbs2DzQfCiBSn7akdBQYb37wdFF
i8INHXVjWvtaKDcJrOXu67MmCDG6AB9vcBgeLYP0kF+GHB/UdnZkReS0BpAJ/z6D
xJnWp5FiNCtjqxenTaRBnRHMoFNKNVevxWRDytZP/jj8qL+qMrCSGcGe33ibFX2v
siIE2j3Hv3S/HRY2hOYqSuYuqawqYQvAoA89xrxXJS8MJCE0/xgB03B/PQKO9Hv9
C6iK85HQIfCM3S6ZeGLBqwrsScCvsd745Whd1Za5OYoAbbYePyQ08VdLJ4mdxWdK
jxgPZlqZo0OjlwjvORIu/IhyrK8KUQNYsy8k3Qzpk2Ou3+hwmKUfLKHbP75lhIzk
sm3N4ASUYfAJlRfsJ9SEB+UWhIqLZCECxgt8oTVjvJ63aqjGA/EoXHkck0kHG6Zd
U4nR4aIjfI7+Kz1CLrJbkVpjHSe6n7xQm+TQHUGp7rYBZtpOl1EKMU9YRtdPZesP
YEJMj7yJn4ywwZ1QVg9lXLBRuKn1fi/vQuACXbGOMOCsXXvt2puBJmLXxWA/P/8/
hCCgASqTXI/MZlC8MspkpT89KRU9g3vZy6LPCFKs9AGflRd0lgBQzOt5/TT7b6R+
rZuwrKh5zeF+GRXiKX/3XE6SQBECaed9Il1ytYohIRRWRBeYwOvip7LIHRmOeWhR
EyYHsgXmvic8yvg8t4gum8hjFLNOpzpCERnuE2HIlssvPrGETs+yH+5kLrrNvwKe
0OIVqJlqOHkcmP6FpZB5KQMroaTXacXbOJfAvWslQFXgUidpgziT6e3fVYJsE+bZ
+74jcPYE8eNpi187Mb+Yk9EBxnIe8lFBxce+sDFK9yIxgciVE2ZxDVoYiX606MFP
qC77RMVoxnwacZEPr6x8pkPgCL+3caqXUDYxhlsR/TkpCqRErtwpP2RGuDEaszzG
tZ0K99YJUOwEjsZrSOokwimxKBVrOo5jVB6zDEkJoBCijgFNiGs9xO/HMxe90FCq
lyndgHl4fLyly2g70u3/7NzNeLbIKLR0qQhGciQMecY7VxI13BBZLxMPJ58hL8On
LHoCy12Jm4DUV/8t9C0kACA3/NmKQAyu3+C8Vwu+luBqCf1f8Y+XTKWj3mRdhKcw
2BnPuFgKj4i3VCSU5HDLkcbV+nnLj/i0tgAxO1Z4wSDilc/V+iV3W2v5rtp6y5Ox
Bm0mTUHkN2zJY0hNoo2y4cMm9MTCDbUWig4YAYlyNfMuIClrqexQplSU3s+aWbEY
4Di+D0ODe6CoS7WQ0anJyBZZj3QA2L5UsktGeO+jduNzPG99Hr16QhLMQ4GvrIlg
rRvN01z75QUk7CFhLBI45xOLwgylkq2z7duhrOEyPtGRy7brg6xUnRM6iblKJx+9
IkYrSCcCSadLjcVg19wfx/f1T7XokM4EMnr0Kf5+i8oluyIwUWf9E5v9oU9vBK6Z
mcbuw/iIICeMSigj2b9Mx+FbsBdDlco2hyPzG/d/h1+VbPBecIFC27UlM5d8dwr/
XrPKfHpD2wlLpIPA0IJiW+E8b2KLbwkKoHIA13qSTnj2h8lE7M2gN6xDcpRriKNR
irv+QE9fGsEaZGl+us872QGAmf13lyTSc5xZ3KSUK7ysrD5MIWWW8VbFJPgrttA6
RR3lBmM246LSSROxjh30N1yitdM/zE7cW8gH4f+rePSLPUeoL1T73KVQwV6KnXyX
nBgJTapZl+DgrkFKM1R/dUl6VMGpuZyJd/k5CW75ud1tu59qHjMqppRoRRw7XlmC
f2Mg8noXND/+LTroj1yQFGgdQ3qu0pwEiKcr9PTeCE1JkrPUfzNsq+zuFepiMO8C
9LKJVKO3glwHRVvG5i9r2HS2Z2Pwm0gSklRSFExrKSgeesxWTkyeYSLaXbr2j+Fy
GK/cp3ibD6fzEii6ahlAgoO5ZQ+cnh0mPggiTY+y+wB7S/DEOANwHkyYzXLNGaxH
zZB4pgszIEiwBjkEiAi6Z8TYjdvRYH4DE1ZBQ58uDwpBbxs1qpDIWxx39a4x1INg
9f/U3v7E5r24EBqm9OUiKmVc8VchnJUtyvwwHzAN5KrJTLKNG5Efphm+jaIfKaeF
OWov63CDh5S8KsE7Z8BOsbIclheuLRctKi43xRvMs3zmJC9SixBHo9Bxd/eM+1L/
082zafb4nUAABlL+SI5nig0fvH2Pr7Q5Zxy2dcL6Pz6nX4TsEvOTAp0sWpVt5Qdo
dSz0cf56FbpFdEtPd/kxT/jMmhBOO0OU4g/NMEw+kNmRly+F0O0U6sGKytsevdBN
SopI1Ppi9EsL/OhFJrU3p79DqLzluPHETJy7kr/J57SL94/U0XTMqr9yHLfHk+4D
pqUcHrv4MvWpyOCvAJQcCihL35TU6M4u3Wh4hbmlovA6Qh4F734SeOq4FTmTDKp2
VDrkh4QetfOcle+39MUweud8B9Bv+EIfziW0UVJ2FcBChqUcJ776IJcwfa+VO70J
HoFSPB7GRnZWy/KYstq3QJXR13qrOgMjxHFiSphkiKqcW0ONvIQfpdlX2/uNfzKm
qpyyOS3flTyXEw7C8fyPLsxy19mRxGPo4q/UZQQzrdf6bXwIHHHFUPCvhUwDaRhY
51aH1MTlSLSVeaVDOrFxRMgL1GEPv/gvdnYiOBvz7nGYkyytwI//FQtkfApLd+HS
feqWoyjDifNrHzV6WFNl2VEwCeQGV8EV9sRTWDZpvqBSAyAtC/WWt5Kr5vCcD9+b
zqG+le0ogG9L3xG16cd3E3qSx/LAkTnmOxmSxqUTLNRCJDlwK3aEwePQeLIMxQK+
mvR3xYTdgXvGtkhvFv6+eXMUuyXm56J944moYTwFUcAn3+ZISy8tGNDufz1V+H1+
v9D/PRWaddb/RrfPb2/vtZdFDOXUAPySuc0FBGAE2kC/6mvPKzP7S0B9dc6Fo1iL
ceuF4xl1oZWRHkisFXBlJT+zHbz+yOgSgW/9zf72n1odrLGcWcemH+TKgh7etQCi
04ygB0kDl3CEHByA9zG+vSi0DqrAF79P4NXwlNBvJfKeHDCriVDvaur4af8j2mEz
ZLorNIYvstPxt3+d8y4gSZgXuQ6ohslDRQE3wyAfb03MfXxjQBGzdFDcNnm518Cl
VgKbGCJHRDgf3fP3brsr5HlQ82DTGoEy/3GYcCNZ4F4Jq3tIAOMqsSCltzHTb29k
3XMzL0+qZ4pZ0bdP9cUTnzlEjsAPLM4muYiyys31N5GOgpF2y5ySTsj+tr350iV7
wo8FTQk0GjsSxTFFETrQFmMMQnbyY+OmAq6zDHwbLKkiU9+l1WbufnFEs9OzUtJI
d+GqnJaEV6Hgf8ubmp4EfXH/l9xpY4sNNXAazSfSSbiQc33f5L6rO2U5c7RvTnJz
ARctWZfvkR1OfnGEUkHDhQ4AVlyNfb3c73xCZ+mjJjEPeYRG0WagUWX9tFHqMpqX
9xhYzwxbbstOXPOHLRIn1lCt6XtI2Zgt6wbmK1TZP65e/rjAL6UFWbZwHPottlUw
gjJM60+hXNbO/u839GfVP02DOBGvZY1M0C/6zkRLTyufzhvbz9e5wYLEGipQP5+t
uC9I2LhsHiSNHq47eb9fwKmgU8AAbeouqHYHXDb36alnyArg3/+w6eib1NXqTi8k
sHii6KMHvPAY/cTzSecl2G+r3mt4Uq0A8enyHREb8CALYWVPakWHl53hS2ds7/8i
60AjJTGhJ+N7uXq6J10sB+pnzNy3OupkonCzQ51lbRaadmhDeT4v+fg50AjhW0Ph
Ve1CDTJGiSxST9ln4Fqz+ut/CiHpsU4PLOZFVsXFc6pJQ103LFMf6L2/ZXB08wKv
B75rYGToehf04wMnnEsuV04psjHFMzAb+dikm+tXZFE0RVWjybdmTs52H5j1phGO
SsgYMMmk8oMaC3Vx+hLnxkf9AsoiVk7wLFa0/ifRl63A1n0Qe3a14/4fMuv3e0M4
/sslwV3rVPBiyOgp0kuZozw5/xSFDVI9Ef3b7D1/3iaoCqwfh6pJeuxcrSP4ERC1
9KWWoU+/PxSMKjXFFnhk4cpP7DDKI81kBR3RhWOe3eY1odOJJRtPyWLcYgL+GKxk
Gm04CO/lctCRqDc1+9ztL16KAtXSlI8EXyvq1Hl3+4HCwYfQEcOAf0AOD390bEds
sj+E+aBlnLIEnouCVeo2kACLCdQ378+g8prBlnVjE714+3CrW52GlTzfCowXAhUV
EofPw+IrDH7on+H3DErldxCorEqyEKSclpnikVK7qmlQkUwskSKTy2PixbqWqntL
cNrIEuGucjpUUhoBMMCtMxCHiC6bb7PGlgiBXG2P61t5W1NwhyLz0LVaJ7sQLsyD
N4nNVzJp3w4cg48H0L/gVcmXls7RTAof2cwvs5jxFXUeG3JUfLKUL0nDKbEuwWYl
yrdN/x4GBj8j+pId82gIx1arFVIf1UhpgxKt/x4aZNSm0zYN1tJyJo0jgYOnc447
YzMdEh8kPWiXjD9B4LwQ4TEFR5NKrqtvKkYdUTE6YBqT3c2LjRloyI1LiuzE4Bq/
CxeoV2n/yLDcMcHUkr6yc+lUiIU4swcrgjXYcF7K5LZo8W1Lp5I1VTd/gDO/w/5u
won+UnekXFNaaoQ5er4W1CRYaQzdpmNIdbyMj2dFN8ADSzUGjJyCblcLR+Qh51B5
4uGT/BH3mf5BNigSc29nLmr3b8bNrQbNJjyloULsxlDahMAw2IZ0/y1fDghDkjrb
Q81VPuAxM02gXtt+E4b0L3avebwyUrwoY5GXbHFN/H/kKPDN6ZN3HmuQvoEVI3X/
oqpuvSnWfdCOjV0GN6KJDZHqCMNbJxALIouHU4993U+K+iU9vFpXA3asokysLB+i
8ntsfhz/3gOIb7TswF2Kj9H6thzYYRIfq9R6dHi/vHCmzRAOHMoAD/PFXtDPk4Dk
pGVeBg/NdzHXR8872lk5XLXHKJgCsU0bEy8+XFcazPz4i3/1h3IN8drewT+d7crg
nIeSKeurXjvIJkMzD7hSBrXvFZq1SzSB59wKas5v3wu9VcE5d6Mip3suXAkI2YP+
rlPx2OZfYoewQiPcSwMwCXOf8hMT0b4KbEMxbG0eq9+RjSKqLubmcFnHd89A9krg
v5MTNm4l1KWF+hKWeJkpGKjhC53zZ6C7xo0LKKzx4o65fvSx/C/cABvt5Og9Le0P
pz07dMwTHtiE0XbI5FcAlGedEGrR7Tuhagi3CDRYF3ZAE5rC95PO/u4eFFweRE1Q
efsM/0hl22WKLtWeBP60+cPZYGCwnpJYrnmmmp5cJwmk7E9BHdR304uK3/+hdJ6y
6liUisRKdPYrlPsqDKr+NUP1IBQLyIy113YYCpnwpuqOEaXrbrkRa5kONP8FReOM
KwrXegdr8dyr6GJe1TeWnmxeGrjBqRHChSZk1+Cw3xJ2uuNzXjA8viABCbO54gGa
0P0BuvZxUrTDjjYmvmU97EdRcpEM3EUGwj2wxhsXZMNgV7h3zCwg5LW4ebL2VDnP
mPMtjP3OAcMaWMXeHNFnAUKPaC8PWc1WIUtUlmTEiZMTA7If1/M3hzBvMMVAwCMX
z5Nxo4iTrhGF93B9cS5RUypdt4/G53eRIZL7vfygyFOu1611bO2p/M192l2JG5PM
PXZt4uqeSwffWpCKq4m5f2IemtoS7eBOjioZE96HBXJy+BxcZ4+2UfB5mYJ+udIn
ruAHdkRlQZbqdn2tfBEvlgrdHvuUOjqJHNR8wy6CDY+1hsnnNrDN0UvOIVeFIu9j
0Ab1riZ8lauN1Ianr9zrnJwX6xn3ChQcQDmUH0wkcw2qYoCtkR0tR/VGRigovC6m
1p6J5LHcuXpMezk+rWPbD6ElqtmiPkdVNKHVnTL/YEJqCoxUip5Xk1hzRORP3WDX
b5LMZ6xMxan+Jw3yI/eBsTvLIcUm2o58SCPdeJ9GS3yjZczPVtn2GgTj3dVGtiHd
Qx8DUaLjoaCMfKLVu89eFzciQ2hclOF1VZwZpJWp5lCALPHs2jc8etmfrjN9cBZt
6A1tEIDlY2n2gwFNfoqUtbh/BLM1ZfZlWG6N4E25ePncCnBNjCSBSYZVY5NLyoei
7jZ7L3SSXT8J8Y2G/H+5MS5Enbifoe1pPLQOAakZmH/iRJ4oXFycC/7FHWItZf2z
B+zttag3vp339PWz1HabvSvD5GMGzB9/9BTilZyTRRWuoSnV4rFdzVETeypRndvF
tSnGqLINBCPyHpwiKidwHG3w3N39JJp2O5RU1/yKFPZIcPyf+hLidYcx9KwQOqAN
1vBqnDwJfM7U0CJy/qbJCxS341nnxAxaWQtxmPNi4OMskvNHwkwKtEYc24tkNwfH
5ddpzA5rSexZYwj/YN+bTQo9fb26xlaVi5mvEluxij5II8zOOkcTZ2sWWUAssF+V
3HCpXorrttZus0l2KRu+y6Cq0kMBLB8EqSWVFhJAzqO7IhIvgNS3SrC3roq+NKut
jVHY+p/bn5xbYFGscOO0dJ0S6pcmMyuXy2EieBZ3wsBhbCPjRzgZoaQeh59Vzsjn
XEMoJtE3TazihzmnPhxONbvihwynFMZVoz5qThCogwxc7EuYVnIC+pCfAsZtwU+n
aiEbE2fHvyRiSY212FOHjfz3dMKG607jGnklWD3xiAHImeUOo5zF+MrbZ2GYAJEP
McsS/s1/E/RQ/bILXjhHpoiVlejdpagTf+TsCMLVzsWY276GjbiRxyT9lwfLHBrg
/8bheVkBOGa8OBfCsrcst5nR8eFxYchIkMktSWO0zMjeKUOVpup0upBm9JNm1isq
YCh6E+3NFlhONoaq+sG8EDFZPbWIq58dcHNNwsexR1zrG0WAfvbHYnEcXfw3q50h
dLlNqPnYLgw40jjjjx4PiGetdHgsINBq4noaw3eXWpghbWikXZtpvsHrfB97HUth
pgDoKcd4lpxD9sbHW2JZsA2tvEb84JDjIarg+zyL6eOjZm9XbwJMWDLS+wrUYaBd
x2Zr8D//yr/wMEY8CRDumCmTYfDX2W10jasUC4mU0z3AcGRA/7FBSmP7S7Esz25t
iWZYc/lGtbLvrRxL3+eiZBwA3VzXSkJ4UI55/aEpLXAJjSL2Lt2zo9K42s4a4TNq
mK1B9VpEwIjN0VumFvfqisD9PickJjDSvA40Wtj2g0hoAsZnNwl5miHwpfSo2yxz
VnhgrESe+nlQ5ZLI3W7qSA8hpjhGmAc7szXTKKFCzF2kfMUyBR88AXHtqDtneV5p
+eKfw9Cmo821sLZCmfHim5KMV4WC8AMSrpMvUaj8NtIRa/RqySW4GIm23kKx6VFB
Ph8zVZc6koTBkMefwL7P6XE0a++1C/4P+rUX+DaGlF+0g/1+/YtAhQn0wISUxiZH
t2e8xW1uC/tCAccLvvNaHeur+qvncqfHhvE9YHBJk08XkosLPTq73ZQuGDbTyTUB
ODU1DaRl6AEfRiuCw18zygHFb0qZuzdVSY777rY+frZUBJFffbPxbn5tlMUsRmKz
WdbXpn/XSN+CH4nLPI+giVN3rBmY8tdMxkDqSfrXUOs9jiBXjNHP5svg9JEFrlEz
3FSLJ2xaUpf0Mp5rn6UsulsjX/OQ3KVgQBVn5r+KfvbNcFEqlOW69wtR+Dy+iLQO
kK+hbi8yg6rfemZs0MpCLznk5zHkpVQwScOLJ2xST5LJYqyvrvQOTuZC7qa6fVYH
1jdU+z5aPeZYHaZNLkY+Xdl6yalYetCBRjY50ylFIXra3RsMMzHTvIvVJYSTDox6
Z2hWasYNhsIOmqN4xqgOpKouAUk2X8IWM+c4TljMop+Pq3uQbeaS0KxcSpjAgKYN
MRAVdCiC4zhE7UPtQLI5kam8OFobKiBGMdnw4q7EmWA43fkX5dzKRDsYWrvcyHNj
Aah5MXCpCbAIsPMaiIcVnhMrDP0IuyAE1rGeF+1DFb3HZEcKltXy3fcRrzZs7B6e
T4kW2nAjSrTj7c+gPSavEVvLWm4Ug+dQuCWS7sQV7D5yvNRr30Eky4GOBRtDbcRj
F2FutJpNyfw/26y4NdAaTC8BqQB1U/vRJCHuKMwr4BeL76ResWNDZQcROWpXLvRQ
MAA9/v1d9QcOSI9GtIiceRXZpbEbybJw+UcY95Olt6gdpVP70TVLmioZOPda9Plu
9d6HPAWEsxY/WGZ+NzEkZWzSW7xKCYTvhFehM/dghugeK0z6Rcugwy4EJcmXQoWi
TpsbNvn2z3Naqf0Cdr5HmXfHyjbMxTPyUHJZkvK2c5Mlh/oKSW0N1RXSrS1vD93A
yeAY3MEp+tqe8qjyDk1fgAe0LFEQM9SNpf8s4GztZze6HNCSOck5PzDcQUW+4TKP
SEjVuDBf3dyvNHX6g1Vr5RRBlrzfScmaoxmhLoVmwdIAjGsrSB1J57lsgIkSfd5n
JFSDjNIFhgyyde60yTE0gVA/f1En5YMVpuUDhMG4eqAz9E70+b2eJTV7CLMeEITq
Ef5WxHTNZiFHfzZicxHzTNdhm/B0W/bigpWRdlF1cHKoaxj28ZVS5ZTvc85LowUD
eKHTMjnn9g6nAmFLJfJg3utLGHU/rvdZB82FInzRcTD3e3Qj9JIM2S5MmsyesRWU
lG1HEs23JsjIEfc0BDa9S27tp4H2eDfLy2xJzXuvxkYrTIxAUObEWlml8xC7MpP3
agB0zSpY+8uFydiSBszxl41YjbNeZHC8oCUGojp79KBvjoKaz/Qyv/ThFH2mUwhN
GJKpsnqDAa5OEbTWNXUeHn3iuHrzO6H3IAzngBnwoCfAjs+neEjh4w1CwLdDaGjb
CnGhidsgxt049WUgEMAp8hqkm+eZRaizQjQlrUComlyz4DkAF8FWczxWRwloJTqy
zUwGteJ31hEn8yYBbVllzLGPDQM6Hem96slR5SOX4NcpnkQApIs8UyMwNgBZgQqT
WloDrYfgNG/PH9XpEB5hTch1u6wyakbCAJtkj1KrUqbyLiFR2p1aSx2AvIzM0me2
QjPaGQuuGGwD9BF/KJEiTPNMstSN+2+uSDlP2KKmJ6MsX986AP/creHB5F520KXL
0+zTpfFLpYOlL383rSojwdoEI6g6npMfIuAoqOhIwVuni8r7usgJtBdSi/H4PQ+H
Wdp+nLADJvAOOmO4LlL6a5qw1mRvPpRx8nQ2i8xIv/lNfZP+JUdj4u2Sm8fMlqI3
88myWrtT9v45LJdhK3NhW7zKmCSIqf6GDgM9IUCZReogo65PCrQt5SeRc9QkSPi5
BeomobosQVVZQF2eYKzTbg3HphNGhqyN8SOrKHnA44R4injghcELnve9l/2yvdQs
lFUye0tFX4RSmOA7gqKmSM5OdHXobK8+0uJIJEbXMIrO5eNwOLXJMV1qBkm8ZIxq
w34M+leivFB9nR+j1jDm2OTXVbmep2QzFQrSMlmuCvNw9FGMquMuTFdcNVzNo8lE
pH437MwLAgqQeEFwJjCmwkLUQoQ7LAvxeeDN8HRwYj2CL3NJIQ7NSx+MrKfxAkMu
4f7lCrIBN4Krano5o3JBTi5EoY7is/IFc2iMP3GKX7HP+dizphDqa0i+nvcA9nym
Bk/MV83h92E3VV7IXQtN6eGScnQkqNgGLkPHTpUQ7hBX9EEuPD6KvAEclJJCEkZc
lszSponx07Xe6h+IvSI5P4DnBkbF9ThSG0lbZXBmIP/KWBRWrYcIi/zxoXI3VVml
/3MfCFZkv2uCxfc4FAP/nWMLOShw/5+0UxxFq/QqEsqJOiBgBFSIK9cVMRUwqjlF
tRyU/T78nb/Q71oMG9hZVFk3SbAGr2Xo7Eg0cDaXAB3TfrTtCBs91RDtKeST1biN
KkRw43kGfLWwyRJHmLooFh3c2GenY3SnMpAdryIva5vGvJY/om/4JRrqR9Eeort2
56dfqdxwNLTkI3VVWGsKBi+2MA0qNRQu3xxfUy8PrY1PyERcnfd+i1gPlcHj+Bvm
KcgTtOdQsYOeGcZLoOGDDhkWHl5bh54s4fLDWY0xnzNbuVIeLXePuYisS1cL7c8v
Z8DSTy9zdIXy+XRtTdlOvY8Sb5z5Kaea5gyTOBma150/X80uXVgTLirJM3nw337P
dg8lQx6Pt0CUVbWKJDWb86kA8x2Idnja+DLDohKzSpCN76r3bxHAQlzimxWbojvk
JFTPw+spR2/oMiu8PneRo2ZKKAcL8QGgPPUtd/AX8VzaIFsxj1n89JXc2XozzHp1
DvE1NvDKipq3pfUtS8NIevSHTgS1p9Szi97exmukqz+H8MNx/peXsEnuShweNokf
oY/qnU1nbrEPMxSyd3vlfuwwfsPWjlqCBkEOY37PR+ta1WHWHKaLB161PUnl1iOk
3iAo9GbNZFwyFLndn6/t6wcK3z1ZQDjD5TNrNMB1rKubuLphqmf4RbFPelhbobat
Fp1uxRdVqI1A79P1LTNOKyJHqg5Aec7mfanEO3N0Y6sN5FaItY6w3kJTWo6ulmrU
r1dyca885ZT315LonN/EHtGABCcmghpWrkM0exLcmHU2Kbu055lqOLxAZZa/Sarf
Ll6cu0Ne1uZf5t1DQRftwg/Q1/KPC+Ner8vun+GcFGrVPq6YBsRtQOgRRlvCCxid
IsBAfMA1gYwstw+SsG6LQLtEQUbjLZSeLxyeW3F5iq2ABmF5/tk9cV5jcn4NlMox
L8hvUrdIv9/YRTH5/rNQEJmLsHc+L2iJ2xrgqpbDFtxjDZOqu7dxpp91yDPa88Eh
KU36Dsw7C4QewRxbBhXL0Wp75UpMFv0OmZ/0mrmq0T/e3H6i7a7vcUqQFWG/qlia
7Uh8bg/xPJghggXWSXjdita+ByAa+bUrM2P2e8FMQ/8WceJwYx+66IIb5a1dcATv
wDMhpwIYT3x44WCIjiMNl0ciHXp2pe8axYA18xcunBJ4dzKg7p+6LBkfdDdS1aTv
Qq1J/HY2MrkkQn6jGhAZaaPJG4Kk7nGpi4uc9jWUhH5AljzWuAXScnJHbVJzM2Nm
Yg821QVcea2kA8MKj9rJLRQCV668C3wx+73jUxgNhPforhmIMMXJDSbxI/ww2ELM
W35HtQVQDer+CRVKbTKUeR/644o1GybD6Xxwtz17eMgBcCbkAKXKh8lalhoof8kI
sh7YgJx3IrR/ryMYit0pcWqIQU3vAzSXtYBGVLcOvW8ray+KJ7NCgmGakU2p4kId
Fa3MfyIfODX2zW+G41aAa4EyGLQRU1DIWcBlBxlW2u1pnzAx4N0kokyNDq8aLbDB
2X7eVttWp7T4DLYjk04Xl9cE3rwZZrjzyGYfl+YzyfFLW1hTFheW1uHv2w7vWSEv
leW6QlpT/Jj44iAUMJbY+PkKyiSHreoHkkaAB4vDjgWAGA4YwDP/FKT38ILQo0dP
io5gnCydq2x2LchjmTo11omcidYRRvR3DPi42HR2Zx3ddTYWqR/4SMC/o61Fe/Eg
AGIxBGunFm0L2ur6rJM3SdXBZSmNGdVwxXd4Z3eU7v2zeq4gDN+zwt2Clqc6ftMg
ZulpfBkHHow7ldVVhGb6wXLUyz7AxITtQ862qmo5OYx4O/+DsR/m7kArtUOyh+EW
Vrci/9nvPsNvGgY7SG+OvnWLKpXlI6vpRaQf9jVPzNIEhiLaqXuK9QoNthggGRLL
ZdMkekvd6YYJyVqEodemo2t8LCRD/PxvDe151X1PYm5tCpuK96INhHHa257L3fGg
oFsMwmdAZuk4DRdIU6Iv6FKLfZAboWnM0Kkk+bWjj6tctRhFnfLTNmzphG5EJkpI
l4T/7GF6Vm9T/bJediYa9F4+6nADh8I+yHW+sOR0P4y2v44davi4mc0pJ0+X75f+
J8wCBi/f5epQ0FaMgqMOT21XyVyIV/0dmah+G5iIjax5Vz9hIGVvFx9qHhZC/V/U
gU6apeIWyM2ODyUJxEryeLNFM5j5YbIBZpfFXDgIHPqamPS8hXpJLQTKK0MHSbRk
ZvjXwt3Uay5Z5dvf7wE0z2OeSL8WcLUf5OunX51w/kM6ilw2vNKwTyJ/TXocbHNo
rOwYqkDgYRDCLHlk6UucYzJceHu6HpB1CV3yBEmz/H799lY6R2f9Em4qfvHeXzK/
yCQK4F7IRrPJurTDv9wx21AlnoFlkqqNMJVXyfqVn56+JqV7DJboXmygSs3AKgss
radh33XKQ3d5tXmL9AwtaLjnqqKejPxZraDX1cXxvBVpNBPHd4bqX3+pEDsMBarR
VRyydyWxlLDZRe1BLhLramPCIu8OvqwkHE5dDUM8iVYRaMlkqSeUBRN4J5ibgCsP
IhDtgmFyW85jlIGHW5OH6NGn1aUinvC6l+X0oQXvv5Fp0VR5aJAhFI0s/JK7NU4B
MNmZAwHbKAbneBDChdd1/9ryPtCEnWqVWi95YMky+OPQp9nz5rhyOt1AjFqDffCm
4chAuYlnX4qM5d6vS/amewfGauGo5k6OvifOG4qKSOrVxx2RRJHfPmg0uONU1VZo
BoLOvvEvxL5Kdgosp1JHWD6u5xgYSKpJUKieVI6DMInVp+FjUi651joBASrV5rxk
fxsRVXUQbDdCYPb8kVDm33JPm+bs09jYZsZmyStI1hO2Rp70a8jLIjoxSpwVSKSm
TdYmly7ZUdUChsudNiyd0xoF9GUMB9ZWaW3MjK7GgoBqDHx/7lIAri5BuxchueUU
0pM4RmI/w2nEJG+TakpQHAhh0fFMylpbCdJV60uEmFeAFUAnS2i5g5nP9YdxPUF6
lr6KAjGMC6zYhCQVW3V0n8iiqSdUg4sihOz3ElL8lN9rHlGS2lAwRoVc5HO/E48l
AgFU8iCmGLj5Bq2FNHPFnyG4jc+fwF7U4UnbVRXp2oHtfQGhQDyzB1Vzjpb29YCg
8FA6A+sug05EtRnaDmskB11iqwuhI+Yqtkvf9kAl+ZJdEVkcLYvAVBxO5g8vd3rX
eLQ9h627znhSpljZItDdIllanH1DO+wjTlsvh6UV9QyTAFv+OJIqEUbX+dTr5B0d
9gDhCDPpzyPODQ7BiC7j6KQmPkxLpDz5JeWm6bNbqE+9nlVu5z2703En++bl75lP
iqhNgi8kCeNebhPD1f3drL62Uu7fuNGDo8HV61E+/qfvHx0sVl5BGZQnRRPnDqiM
0hAHlY/DHtzv2htZN8jacEbWNRJuxluZsvk6g6T7Jh2oHYl47ImYXIDRRRCS+fnt
I0257Ae9vYaT02eFqGb8JMtS81TkUZUtHYxeOX0vb9j5zcryhtdVt+MS73wjayKq
gYkiKk9aQzm19t0Xlks7bwr6ZzVcIFVEurkhU8vbeH2QpLwe65ME6F6QVlC7KKjJ
6xqwnT8/GWOnLbB+PPCntHtWKr4qKj69oKIpReHFTFz5O36xfESlDEmOO7VyX8U5
g+jADy3nbv07ZY2WL6mwYpGVqJNPc8HnF1Y9T4n1PrppJOVgESyJ4xy5kIk7MPcy
WPhMQd73KG/fBgRN+SIVmxwQFgvrHr0JkAPQlFtGXznB1U3Nd+nz/XUWJLjtyuZc
KRa0tWEqpXojZFsom2QsAeNQSLX7S02uVAqBFG5ThVknQ9v8EGoM1iATd5KzE+k/
M6Trx2S/km1sA/aNCXs7EbtE46CD+EQP88rdIPSqhMRLT+udtlUtKuTluAU9GAYM
QiBX3NvX9mtrxLDXd3Jzpz/exi+hC85RhzV8Vz1VrJIW3rjnBDhpiENeuvd5kf+K
Aab5LE9HrhAgAWWsUW/QTdgsLywFwUgcdFd9wUVznibPuesmY9UNNYR1eWemdyxg
2Id/9K99OZHrkx6Ek1dwjpIlXz76nOY22a1DBxmSAwnz0Thq8GGH/U/VO8xPwCzR
spLXjSYUjU9l5+jO8iC0wxqpt3MvyyJ/OOdTDdTzYQfqdWgtrQxcQN5TUqgyPR8u
S/CZ/IIPf70UGIA3ulj4zYV9DCnoqK9GCoZJOW4P7PpmXa3IRWz5lyexs/CZ0S5M
1GrQXDBL5e1wcKTHHvbCZ0ZbEBnGWQCOuMo05o/cHo0/glOs6kNit1QJ6oFbzSSb
T6O6ZEmYJb4rZ0BXBpyNDJFo3aOg22GYjd/ApOmctH77fDx42ibKMdpvCuZXJgf2
lrASjxbUtkqOzQJLePmB/5QbQlkOkQAbB12oa5peNZsJplLORhmnrn3iWgxGllhO
2BEup+UtwhmXTayqh/JBUZJM5orcEZtc5FN9QoijYQ03a8L/3BSaQ+7gxxLwB28E
1qbwmLaYqSuWs2VEjOlMXgncR7mKpz008SDZAh3IJVBZl8TPK/voRC5UILd8ozHK
cvy0ePe+AiFoUl8cWacQByBXPMdsHc8ECwKYKHu93ypaoW9+mzzyoAyEeZ15Krvf
XUirEGnWM9SZyc2OexDz2QASqwCI1zARwPQy0jpgYBAZ9HaJ3B/P8c7Oby2lhu/m
eZkVVRU10OBblDLepHX2R5WxrCh70qDah3/2OvI9oZKfqQoCjaLdOlCkQFjB0Boz
cetwWAAAPCshZ/PqqdpM5+vYlFc8Qaj2Evk+LE1bIedyqKLBgWb8RP0p4N9YQuUg
4fX3kDrIddM4QaXoMOQsw8uJAM9qQDIsN0KqfDQnBrC7SgsxYonZkJQna0PdKJOS
ogKeecjnuyMxmRv6C/73EutFl4n0nRAKYqgqSwZIIGPTj8/PHjF55fBBD/1rwmd7
cHglEeXZdVQZa5DVXSzr35LoJKKQTFloyrrEcAw4neGhhsRzxffPIfOJFNh8g+cR
x9QHbMvpcV+IJlWwz06XR/oaDZj80xSfhiF9fjn5Bk2tSG0I8H+RJWWcyUJmSlWD
Ic+wkme2xcouRVetXkVP72UOwIiOCPtnDq6wy82XUh8DrR+gf2thOxiTIfPcUsTh
cLd9R4TT9VvLscFqkM+P/96S15+kokcVu0oGwvcJpjFoB+uVmMSEzRVxTsBMX0Ad
SN1C0fvCxgJEmcp16h5413yn6lA82sm6SOxc2+p9NlItHyaMrIgkM1LSyHPjGtXR
WKi2/rg4cp3DDWN05AURtUVfjcw9Z9PU4ON4d4qO4mfhjVduRULhfJZGWFWAQ42U
k2ExKl20Yw9Ix/i6eih8R+ZudPKafUnlZUg94DmoZ2KhOYY+g+F/V4Hwu5B2MYFN
kjKBcTMM4QLUUEHJHIjzO3MqUUGG24NCd18ASsBOYKfxlBaVPZuMjwyztzXRMNw/
f/WyMsSqmxAbNn0JN4pwzjgfOtUMvfgMeMite6p6L22kkhNKmsZs6wkHRaXjdbTU
o6fxh9d2/Tr7EFSHKvDOE1mBwW1gGo2IXMgk4dWlkIcQ9xjbiwEGCbYg0hkKvnt0
M6rudzh0nECM5IRXpv8Vwh+5bvVkXy2AxnRKSXsVIqL0rVGB9Gc2S0qdpUBr9wxr
cWUqzh+2ALA/WH/WiFeZaZ9gqPk+gJVhmyHQsRyDJjf/REr4yt9iFQ4yehX8xBiv
UxIc2TCVH9P2lpj2/bIYguw+fLf2d7LfpgOEpvQbLCxMKLyj4wPrO3SKpWLK34sQ
abAynQ+uhyV+qR7Aj+Sq/4iFflpq4U0SMyCsLlfBwKh68f3JERTNVpzW4N6p5nGb
FDHzNX89huvzBj67B7eE1lFx/0rVzZSyP63rTfKijH91qxXOGIufIx83YNqyCodX
NpoFWKPw+2L5P9eaubmkbQgpisq/qan5DGxzYTwXY/2rpx9YT6MkuyQVFsNUwVBw
drtuF3CTZXvuLka4AI4rYJz9wBXn8mDi9R5o1sXD0fmi52RbgaYQsFeyvJEeI1b5
0aDIcFox9UfenuGfKHeEtX5AJfSmvj85dXU/8ye9Zb6ZCtiyOJoyx1Zt4BbIvfHW
Z26wix2+m4rSkhdI1A6iOuZBt+mVsdN5q5b2V5DK/goyInyi4CKsenChbInWkIru
A6vpz1nX3kiLg4uSM8pjiugUP0h23Qz2sVUSbHKUEOeLJ/18NHazNY7slfHqBhVR
diEyNMPp6Zd3mxYA5ZRnyXxJiRI+sNFXtCZEYzADO5hjMEUlLYsmfNoajjAzb8uP
/ibkKGcFmA+8SnMz2E55+UPzpXd72SgL/IjrTVE+HaeqILhzwUYaPYkV2HMX06w9
7ChDUO6x4V+5rpAEvKOsVhoOWtGU/YAPfP5GOV+pYtfwKZlYcGLdiO6bmxmFkkEm
IS6oNrI/th/NeJx+9nvwRmVz4kkOOaHUlN8ecPG8xaiM7c/8CFoRfWKy6Q8WUy03
9LkUg7Akl2CEwc+1l0SKhU1rjjSrLniydd07igy4fJOdPoQ0qz5fB9mfPJKs8ny5
TaqaJW7MCB0fe80/0AS+g25IaL74ubSTsNPuOa2C6tNrySuxRJGHpe1T+YVQAIP1
BmqtTJwCjTw7DXSIuZKI3GaA3EXubzjJMNeAXlQPDuMi+wRETcTizvU8yd8mNoO/
QMIellHpqpyWLbS8V8m8DsPFaxsGWWY4hfuVOBKopyvhCdbEV50OvdADUUGlHDEg
q7eL4G8KnI25mSrbXbo8m9ezU1mbf4a4Zi80Wzuy2ibCCtQ9foJZmnmy77oQ4C1o
7E1/j1XuLaJ1ISkvHTXRyumYWupmYL/28fqrNd16GXLLE7btD8jllXo/EF4TOuzN
0mSXy3hro0LJ/oWq9dLzrsocONRU1Dd2xv6bZLcSgfRZJMq9aFmnkwPVPDBcONCe
4SOHE20tmSMFhLRkZcJMBV/adXkaV+rvPH8Nyhq08kcx+DqiGWZC3NMuFmLXoJPB
bgYIxBWvFdG+BM1TDY7d/q2H8OsbK0aCrdcRBULVMoskRwif86kkRlecVKqS/XD2
q2nWPHdsZmr3NoWwhHdzY9rBe8awe3x+POK5v5o7Y5ajqWrF8A0O8iqPJgBRgh9E
bDduz2ynYoEmxZLxdrmDHSLqMnzaB8ckhyyxuV9wcenqdo9cah0+HeATrG5+6Qmh
NBPq8wj7OT0A9N2Xq+JqiM7+elsWO2I9o6CPYOB/KAtO1Fswy2VgmnmK16qu7Y+B
BOrCskaAQRFNzLEQayFp1Sjyk84d5rms/VriUVCCKK1idMXvC289WiUFnFwptZkV
E1a6PCpojf/hh2z7IkMyu2ZFi+d4/34uh9bvixpCzKSLIHzVqlxe01On6tZCAGen
zmf1gx2IMe0EppCUz+ydHwq5HnM14OgMLzjI2O1QEUCsdwXIZoxY40K1qltPXjy0
J8M6yR/F0ptwenxkfkeyazyN7tTJu1H+DsNIO7AVmrnpatoT8agFXJX/OBxHWjy5
AAUf7jA5dnAeL6Vkk5uraTVJmYxQPbUa7UwAulNNmFtZpJxIoOJt35rQ/ReOfyo8
3R7RsnGjlzhsP/Subnbub+P+kdbvek6b9vzK/uolOhJFk6am8wOoeHViJPvLbB75
JuozgB4y+ZKKj/WSkj9kvRhPRbOSzqEg6L6MvdWgpllSy6MHGJVRXj5doPe9gv7i
CU/ZZ+cZEHEwcggtQQR10jTZ1HvJXatq3cQilVhl/BOdB/bmmEm1cVnioVRc4QoO
7JQu1BNrInVjlcMXDSoiy1VqlKZHzsfj+uZh3DAzgFuzW9r8MKlj1YVVfAP5SSug
xtaY6xlVESEkul3lJxMF3uXA5M7+zY0/RKnHRCl5IbSBmoyDoVr0S15DaXLf7U5q
JYEGivmB5kSUUSgEwCY9XLY8u7fJIJnuKDLPqK8nAp0xyAwu8voaiynJyx4V0m8u
PBp4cHOv+KIGeQYlmk1HOyXb+zHb/2860jQncmPSgSA9U/Pq6jqgoXTYEv+KkrxO
S+6udijbIqdtrmRq1cAo8wRsVXF18xCJu51j1gQvdECdEpcy2GHeNXgn0nKRPlKF
3QTpGh+bNZLD3HSbDHR57MNqAa9rjPYqtcwYvcUv+TyCoNgTCVZj+UR9H+7oh33E
Sq0ncgHN0dU8tSzkTXug/SpkguMMIbFQKEel6oXaHQ63oOt0JjFAMuy/XHcakGa/
27K+2ki8te4Klej6vJXbDTULJMNzFsgFsbPBUkV1f6NycZ609rUdIsRnqc8BaUhD
GN0s8hu3mcaaJllKVqXmxDKEuRaiJQuib7lpreQj8dM1fIrZL6yy+bG1VQ1jASS/
DxIpDt+YWUtDxDVLWqBBIROJYk4L4hnuycDA+CqF1G/ye2zflBSedrl0g2yBZWKq
K4qAa8ynMbn3zzZf9aSST61rdmYzrv/MINvSKDnmQsTgnc14U6QptdwqoxUCGzzC
8of3hCXOUTUZJtX3FPJBgkLjpUdSFtyqeV0Rv0HMit0P3NkQRFWi2hvJHNqSUend
FZf2rh9Ib8LL0VQvHKQxMqYsMt1Zzxa/IephIqx3+PYq75FMlB/0qmPjuHw+2npV
fGflX55nAJryj78723l3E8o7UGMJmeBxJy3ryDGqO5arg+fChNTrDkHfLNodg8qK
QuyUaCxaE48FOvXiOSe284iMe88eipFsPapgR0r1mBsxNs4+eCD1EU//9/X0Zfdl
0TxP8tmtThkYutpztNfWBpS3R6gioEs5IFrerIiiBgf8TLlibOHeD672t8xKFiwZ
OzlTQ71EqsZ1aN1D2Xo70QcSPRHxlXo/EPerI4CPci5Ahfqn5Zp9EXTSTX7r+/bt
LcXZVnwNzfnSKe1ETgZ5IzCLa7xCcahm9dFlrF3YGrNWCBSYLRKwmL60suDItzM/
jAAIlF+8oAbvKc/6VMfAEWwXWAntDZpqfs99SWIWdW2LtFATsB/zj4CU88eTn/eG
DZ37mHn/U/Uyqc+a6lHqf1Gu8/A9BXgZprcq1wlMKWkaNWVK9EhMKeih4eFT8AyV
r7kyEc6v/5CKjLjhMvVWa1x0vZWK+JcwsNiWrTK+cU91+v17x2iRgu2YKWM/jjho
hi0JCT7Ufyox9p798BSPmDE7YFqiRylbsHa9M6XdXfGiMY0CLjkArvw4iXtNjZnZ
ni7oZCBYWcNSN2yWKzZH+jgRhz/UavKsPEWXcH+04CXojoHLRMlqPaSSTNF6SaP9
reu3/NapsrUy1REiyTTAFU7l64WfswpX51B9mmiOcGzPwLexyo02EdobST3ooaTp
ryIY5KL8YhV8qMtsTLcms9LRPhOcM5OEnaf7vtmFMROjeeKzb032wYa8YW7bGLRy
n7MSVcuxxduxBwZw6TwJIb/yESiGF+8pJUytlzZ/zdVYKLIPqSI5jKFTdujD0x2c
yyU7okzg/jS5IBav+b5Kf2SryH2ju4q3HUxm05jS5yMG6qBLj4MPYhH7Msw6+kSH
t6nbAu5KQyWdgag3074hOUTgQQMmCQGAaxdlvxsgGT3DpybJ7FPuxUzel7ChrY1j
8+LMpmZTA8Jd0OGGAjKedJEAxjEvyIIPMFrPZIWtnEBU1uuZZoLoZ3qoYIAXKBIR
K7aHRaIQKTtPQUVXiyQ+Pvsym71rONiF78h/pe2+VFxq4shAhC3vx5rfas2DbzSu
mX3qYUooLQJsDcdGWY756f1+0IjEESmLNuEIb0X6nFyWyGzU9NIhAbPAWK+vuGFb
p/I3hNc+vf7qZxBkANNzjLkkpgJsXLgxDyAz4Dzy7i2+O3J6vuSuPfrhqe5ZbBxl
+hfxcLZGYm0ITteEdc6hqNeUGjuBBqVW4z4kZpNbe2Ks1UuzjWpwDoz2PxLLgwpp
j6touuLjRPKobd3L1+1MJPRL6wlEsO7ZaSgQO8rNZPLDkaqLANA+JbFdopYYuiiS
UYsBvVWGRTh4+XeV7xWg/eaS1vOwYcrLao0vKMXQs7rjY0qeG7r42VPqlrKzUZ4O
p2vqgrBCVyw43PurDi7Hq2UHyvnHlHlsrLWM5eu/Ecye9oaXkWoAhrTVfIFBbABH
cS9eF9miGliq1VWH6UyIBk4H9d+OPPRDsYSVHrM8+L7MTTOQM25K3SLE2qJGteiA
CfGu73Eob6c32o15M+4BjgLNvxSXio3zNpyXgxSU1SI88FxCx7/AbrUbYx7SVs+D
tiiebsko1VQAGYtBr68uNNhGBTYpmY63APN4FcYniirODFmpWTZXun7LfCm6/M31
Tz9EXUh0h6uYqBRsMPWxPvsIzA1G5R2CDy3SOIvpZMreaj5IdU1+csSXGtK3ma0C
bOaboNcYLi7JVN1aAdfqV4PGAI2xH76xJ2phEsOLtm5dkfDq2bNBV5PpjQ8fNM1n
SnVXibn3yqSH/wAZ6N1EcKYWO/kgVDukfh4RsvkFwgLwfRJ5mr5XVVYGyJ9qTTzB
tE/h9lTpLERXCpPxafxgqQje/eE4hzNeD2Fc9qXZW6nCb+fjOw+JGLtynfGVdmas
vOOcNtO4M144+ZRbur/OqtmyH4p6R7c6+pjtw0qnKNY77vElqAUcqCI12qOW5eS1
nvO0n5u6EzdkMbjDxfXHKiGBc4Q52HKX7OkyEyltLhFvrzuG/xRB3NETo4/lR9Rq
OmAKj3g474x1yWLYxmRMh1ClYF4rhk0GHRELPnwTJwZ5CLs+qjW4mpD0GC4CN90A
9YhnSA4DcsdFZB7PQ6UsSYLAPJlLr3cyzUpy+u4Ms6SdZ4EKlSM71fJBjASw7/QK
+K4eaZ7dMKYiAPAsa6vhiAsR3nv+XFWygDGhdM7u9Xlu0SkIqC1ZoD8vaM30+bab
nxHrRshoCGrWaIgb3EcKay3x2FwvwRC3foCa56V4bpP01fx0Oe+K5Vvu76Lij9TK
EsF2/9crIA/Qib1gjwzFIEP5iwqbtYrdcbTwNxbR6suj2wFhN1hcpK5RCc7YTu7N
S+w/1oLUV9nqC9jLcvGMSYoViKnohhBgRQWw2CrqMk/rHQfGof+y61HMu3w71ZZ/
BWaSFOjYPVcQYTadwdsHCSWOxIApb+eqit2KWbwt04zADemT+QblHoy3cmOciF/M
QwQ8x+X1O7WuRL60qUnJu5b0xcb8nYwA8S88rtW5ZnV69Bs9fDrLW4DWvbG10gn5
T0x+smTe1gam5XCfgsW6Ze0DBeUJOmAtEh+nM1jKKo4x0klFAS3jqES/OudMWRMJ
VzMkXl11TmN0NcGFc6rx01Cyq6Dlab1vHxmbGe+gnixqm4m80hHBcjaLm1mPhhfw
eA2lidhuLEukQXFPLmlsph1ju/ZWtgC1I+7adDa0Bzu3bV0a/EehI47ozJHuEqc/
xo4Tx1adRj2hAbmdvcqZ2qmUuPjCJoF4rylaL+VLo+e4mKvNIhWL0ovfIjN3UXsB
8W/3c/IBNLSBpi30C5M2QXy38bXV0HFm7ROsEctMpZqW7MaBtWOZGlVbvHmthzDv
HC0M2mNxxmouZyN0JuY5IL9xH/DpWCsKB0wfKd+hT6eafc+WPe87CQ8Ka2dgy4Yg
uf8DGi/6+E2LzroQJLEdLVm2IAY7CH3fcTUg38qe7F/Ye9HBOpW78kaitUzJqQ39
Eh8EKxfGuK6UvdDOZqhUCje8OAKv8y265zE+tyshPkMPqNxknSHWeLsciXOu/rsL
DtDoy7lNkoRc6JL1+kUxpUnwSf1EzFbJUkM5ISgAW//83I4kN4nuKZdkk2tfGrfa
Zb8EK1WCgKta7Ykk7WO2QoXg/iz65ssGoFjKWDHhvtUGk4b6std1NaEzhYZ/2dMO
H2Npph+j4t3Ui3K7B/1fenHAGU1T1wc7RD8pUz0+oViEkyhGrmJbJLc6VDS2nPxa
vABJlkFRb0JVlt3eM5fVupvaxhpCrmsM3Dqts4cdy4uvddO6UgL4+WNy1G5gYyko
gjPXTBY2AhmZCZ2P9uTCeEYX44tRjsTBASunCHoS8UJaUuQQx1IzH+YKMGzNopDr
6yvDlQQClYZShdtOl+coN0gKNQJV9y//fowCLW1hhbMgzsEc69XS6k87Y3h2AiCl
JYqygHMuQZEGxRzXAyDUglhgQLeDJODwPeOZM1x/VLCqWSlLmyP08OxvDNX+vBuK
3V4nzRL4Db+lJElJrnfV1tL6M3sHuUbWM+YMnM2ciP2qoiNs189lkVU9oHkn9GOd
mpkYSa3B0X1hahfwKrB9y7rN9nb4x67zfnXKaY5jNAlGJnwT+ccWdkGTu5nSR7wd
iv2UG8fsb7i3Xw1FAI+QTCeecOBbCbxWVI4ai48hurxgV4+bKJoXte5C+CLQd4Kj
Sok7BO56oEZp8CK2SneJODAUZjLnLtJ+Nw4fJiHwR32GTn5vfTUHOKDS3f8UtJKw
CSWQhDnvZ37HddcEKc6nhsjOmisVm0VlCED01W3oPfBxSlKqw987x2+GwGMWpbJy
QQ2U16phjnFCxieKzOlFuD4P8qzulz5PdzpniMS38KT+zTgrNOlV8Svykllxskpt
cE2doSuvhppRnOXu55pYTF1EKIIAxTEZbfdry8Ze0AVIss6LzwEOvKpG3sDaDd0g
6izyFXrlwBMEiteeOoSeLK68AXDxWZebcATeMDpNftMP3DBstG9pj7YiSfn/YAvh
B59+LcrbpxA9uwLJmVECoEMLoPaNJczulAUxuMMH5XWHsxr6fj7+o1DoZB5Xnw0a
mClF1JxG58HCHJw9DLf5KkMEe7DBWqV/H8OPIg2MgjneeS7HkLF2BR54ci761187
Y34QJqg7BmLzyL/8Pp2vuhTqGKjmFojM90cgMtVKOtuogxPZBu2tr1dnTTb8HQad
IHq1+dhRizuzjL8ypBu2ZZZMFCjy3VGWYM+zYblDCLcbPtH3EGZsu+/OymnI4ioY
u9Q43Jeo5ScXyo3L8+ZmdEDUGy1elyTVYm437IJ2k25GQ05yMXaxJr8KTepzhW6q
EuYTGU3VuGHUT7AWzIQJcPPsNLY9SQHHzQv0PALqwXPe0WbHT1diUIZOAxOMAPr3
W4mwqz0Fda4xKkxQR4JVFXSoYLg5wsf71MruolMglW45+EV2qBYhEs+Uuem9B5z7
lvTG+aYk9QyQ78vvUD1Yn+36Fk7wPyeuBllH93niCeGRH7ci5JyTRE7FqMdSn4ps
ZfRwlkmFanzkgB2V0VovmbTiAr64Gk1yNkD3Sig4NYZdWWayR9xtJ0RWxxv5zC7u
qrYpp8iRDthd+Sya2sJni0mtVkIVq8sMlu008x1IVG0xcw0jdimmHJf5OI97RBre
HtDARE1XSMfnOHfTosO8nSLyCY5mAerj2fBJsGfeZhXhdSHcXHaVlneCPUyO39LI
qjNuUdpJrGHXhxxHifXy5ZhFkkVYcyw6e5MkJcNF9Q6NzrMsyhEYqc5CCbjuFNrZ
cnmFVhyorihFCkyq10ov437x8hwX7lhHMH61bE5FtUPBEE5aUdGjJ2e63gK654Fw
llg7rceGwwd6hnsasAA5M26BRC6oItIJBoZBiS1DRe6NdxAKxC5F1PH6pfNgpE1n
hd5QsRlC84tT1PZsj3IwJ2AkFdHF4j7VJXr+jilwMaVyg0cRcvy0UilflvqG+vtV
JXur5RiN1B+hlehmzugVJtajW/t4DY/HDW2bXgg1mSB8mTILhRBImipe33WCzmwK
eupmRpd3PwUF0Z6uj6+ShQOVpXbOZFn0nQspOt/oGKOgJeTDoU3s6Qj6+ppHPXLY
ARUMhRTTC/iyNINJEsAKavHHotXnNfjNvshc+nS3iELJcazgzaJ/6Y3AwDjtMlId
uG10F5I1S8QBJL9lcXH9cmilcA2hGAsZa53bQUCZN4WixPThmm25JEPAg8Qa+YDR
YnDsD0i86KmNUkmKYNAIfQ==
`protect end_protected