`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
gMcHP74wBZczB0bB0IzoP2xg5wC5NPjD/GsvSQ6VQgzYAsanETMwwsWi4yhFtJwv
5kY07u0WerSDf8woJ0stqW5xF501W3JLIS8KMiCOd55RHBOnavjYiaaLeu7oUCmB
TtTS1R4sO325rP2zOn9YwRbyyS5Ljn+PzFZZUmkt5xMca3p5NGqKtZW2dV6Babni
5HlLuF20Au601B75m2nv+ZRoGSrpkNElxoTibONmX8gBflpIVE7BehhHwaKSucEF
pp4QQ5zZAZjEC6aplZepouGVggAulz5AahlX5bf4opOVlB1J7IrgyjENtw6ysQ/q
DzybQ+ipztSXBGhmcCVU3A==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="jAI3OJE9Sh00Sic4PtM/KZ4WjwT98XM8AMZrZsQkxWQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hyw9IrFLPQsjvXplweG8O0lkaSLBN9Ijv4B5VdTRt6ipKJT9Kzsb5LxCKvkQyF9n
sGPOd5i74hRHnkHfYISGkfxGJCa55ieOyFShOsqTKRLxclm4oja9vTIey6yFm1BZ
54IDCG9h3PqfDiTD847UCSMRvFssyycwv+BRHQMQlFs=
`protect rights_digest_method = "sha256"
`protect end_toolblock="BnLuc3jxknmZOyxfJK70E5kp9u9O8IQ8cgkXv26kHA8="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23616 )
`protect data_block
xABArkLxBOK6xG+7CdOOiGu0zbCbHMrEntFfAZEE/xRFxZaAZl1QLkuFI77OC2KL
XxG/mrHJzO3taVHgwRXNLDdc8ePbxbAiQfzV3NJLBO+gsBjmIymaCa480cPNpHLx
12Ds7rEEcc/qpJdlPXorQ4D8ZKys0CNzHN/wuOT+N9FDgss7pdLEpirbgYX4Uptw
o1oXKNxMXgDn+qoEkUzTmllBANOvISer21z6Y+sadw7IGVt4j7D2IysKiXjfkqAI
HUIhjDmxUZzS/U5SBquqNrJe2uy+8+Xf4WlqWQ4iFKJvKqOIlZR25KiJOzzltQv0
WsKxbXB2v1+6cxBdcWpy/wbe+2zcp3DaRL05xLBayNPO5IqdDCDp+4KhbpH59hfY
6TfXZIAgdWo3Cag3fERe6cHxEFB8mnmHTeU8gjg7/9brkCfd8sZeJ5eGYfoQ8UEV
l+UD4Qa42N7bL1J0ZhjqX4rptWjAp96Qitq0Xzq/nHnKDQAgrhXrUYOl+MyMwRqt
3QENo14QhlIqQNwMz77QKvCt2ijcXC/inpBPlnFNZyIYdlNRHhiRc5+NcbEayiDM
xUcwP9hPD2dnrp+01K0ohOIsx6o2DKn4prFlYALblzibCvB501l+QWsisrsE3s2q
em644J492chnPcunaEEENR92Z3w4aFS7tz2egG41ELrKV+tNO5xBnji83tOUdnZU
CleuH/KdAI6anS6JjESvBHsIA7OLG4utHGnGABjSwGvxoz0w6Tu7WYB+pBH8SNyr
2fmND5r/hp3MQOefHxTTILEJfyKDzD1D9m/zwgMutUcafnhdBlUrfQzI8Lisrz+f
3LDO9rqt4+p8ehvt2Z4GOSARc0J7EDmEvwxTVm8cXRdcya+8fUY2+uDTXxC1yx6M
q04nKqvzc5xTNHgy8nE1+Mg/pXw70mNjhtXV7VjXkyfqa17EhOdOTqVUNyxwfS8Q
mLXecCJKQ/N65+avMXvu0+UH2JL4P9yYEBwvcEx31ZdXHsnanlbffmtRre9HbMYu
krLEwe1UbvUrYxJvlbJP9s1/O1JtpZbrWHtzsYBg3Z3vxu0hW7DpkwhaXfvVw4wk
j6xtR/JFNxzLsQ3PsOVNZIh0a7MT2t7PEL56hDI91s8s2iPZHrfeb1km91KnKUI1
zPa5i7u1kgfTKpJhoWzqiXLM3XdosY/cbSyDNsC9sw31W2iCccXcX2C9Y/XcEDiz
YiKC2jUZHIQLE/g99o+ro9wtUKLjDn2dTNjF0mUBl6zAL9b9bvGO1f6APUGcFJdO
VZlwHwZl6SybHxcBmiSONaP7BRU0+DA3dZKmuWnfDC/1sgmk04+qDXags9kjdJ8N
fGzK/hpznfGY//Om6+c7LN6WcjvUoHTyxa2bpYwjKdmRgeNFYPg4tfByGhZNAKxW
D/3g47hzQS6bT0Djn8CVSuBJ2QeAD+CFxlJqzdlAj22DryQz4f4mlVeOeNHhhrmz
2b0RUNPiy07ZD1WDVoga0TXIXdqwe8HopZnASVtod5OP40jBg79jaFIvgvuuNkJr
qS337EdvBxqmlHjYmQPsoL/UYl9Mng/TZweOD1UmnhjoES+vvCq8G85KvoW0MFc3
0d+gqRTU/FgKSguiPt6JchET2MTI3NOFc+Ytd5QFtmVQyTfq5XyHDDB5Wm748oLX
eJRFUj8qjuXblW8aZJLRRweNTKG5RZR2UVQ/6jd1OY9HUN2OxzsjXrBBMNEUxolJ
DgeSgnMomDhz1cLS43hSxNMIWpNh1yhWkhRaIoTIKXwlR8Jisa62gw0EcPmaU+y+
5SBUHiuhr8z/oJqImaJ8C7DWSR/LLO9B/MDjtI/mhF6nGm8wiqacn42nZxOGv7jr
X39rJMSosmipv+Muq8aPZfMrujwhJvErNLA1GdMt0hYN6jnAEdrhxhYxZYJR+INS
MbadVKpnCVpa6Cz56RN8N/iqdLBk6kuhfBMt0G0mQIodgxcKsB/i7XnOz+4hiKJK
Iaanht2TsOzhgnj+3tVnq10nAght7d1jL3ZS/XVEPtPnugiXNE9tfIABqEj6v1vi
LuJnGe36BJIbD3EbKLnFK7ka99DsN4g//Zqny7q/9H+zLpY+tvBWmsJ2sAhCOBbB
POO28iLODpBt0W62Uy7KPokIGipNaRS+SVSTzCZI1Q1uxFhqPJxkFfgxH+qBzsJU
Ea+72RCkEghsB8w5NIXM0QJBSqXu89C8TF8wLU0vt9iC93K45vhayjFweRiOt8UQ
+I+k/1FAuN+6aRtFbCHgabVfDRlVIlB6KuA7+X6+4nqcyeZiMnFLAIuPLSQ+hW/H
BhwESRQqgqg3H6OLw+FL38aw4/2Ro/QIIHXyAjUII9r272efmzD8TNNHrXIylRPg
iPDVFYq2d4XyPQpgSNl6dpIsCdMSWe2Su3WcZw5q7eXtXFsPXBhofSxdSOEXCRnt
xuQSJqgDIqT2LgG+bpLQClFaIQKLlRCGxwkR9uOSfVmIQvCZb5KP1UD6ShSlXy21
0fzLRJZIBjADD5uctA6eBaTdbE7Z2HIbGbchOJgs1LNebfesNEI9WzmPZMgvTSrE
18bworlCpTlZSKbbL5kJ4qfCC/UN1EEf7Adiv3BiqNkuaXrTxcGeTw1XgNl7gqP2
G/BdD5UfYvxhi94DHV+Uc9jMIngnh+5yPLUkPyV9iHXab/WVPlqvfoyMgu+mF5Go
nI0qo9AVSY1Id6erJl008Q98gtwZ+DszQ8Q7s3hO7QxWAo6RffU2qnkJzMhQm6kZ
41Qg7ty5fvNYsJJp7LpdDt13JM2n5rj6R+tYpMEBOk3uLKvn6Edj2Zq1cZTC4WcL
jPgVeyaQ5gf/GOFunflGhwI2DmtKRex0cuyqFQKvU66e+4HqLUkCPQyPHv2n0n+M
XMOJgrdz2w+mrQi6T9eT2RIpCxSXtz8OfGoYc52VRks9cf25QjIlEVSHGU8qz89X
fT/2QUK5uBHoIb74JP0D2E1MxxUzyr0kAkK1r3QU46HD6W42yxk5R78+nPK8ZyCR
ZZ5xPHd6jN+FuwI3fZP/dvGP/F2I+oiwpoLieBljk3KWUuJfuJaXqvwdk9HEa82+
uMrPRQdxktVLnMV/C7Cn57ufRAZ2jp97rTX701xktZ2CvheacCqhwCuaZlCYR8Po
rTp7lA5LsWbl1CzsRmhMUlGy106zr1qjARqWtJR544IyS+9fBI/x6kIjS005JbT0
BRAgL+Qlx0EX1vyszoGFtgXXu8ZcHv4Zc19/1cIy6BiLrh0nn2J4PpyE26fi2Fvz
xBuiNVEgHtf10apo6F6mgz1M6Q/ZDbJQ+gEVCtZ8rrxTJHaKi06yKtFgVQbEvOLn
wCeTf1QT5jUOtkMr5nVY5sdbpspIHgVY8mopzdS3dLp4Vr642Aaxq15utO3BhjST
hYn5OilGgqmXjb2BdE99eRv56cDG4OwD20tHzMcq3GH4IdE/tGtoMlJeaBKEIThH
G+2jquuDzGF4TB1K+bCktDVfXHI69NPLh7kyv8KNPbKAfCIPEe2UHQOxreuUTTLD
VLFw+JwLxsxbrTtJKTJO4PrL34spLcN3WDieH40XLCentBLWREh6i24YwzFpVv60
MbbieUp5c+MkxnM/7Wl8LcZ/EkI68tZ0lQn5VLurh7VTpGs41Nmi0GCa8EeyMTPw
mt04qg+EQ0/M7nISDAOXsZnmh9VnfmcqHvWyQ8CwVudhdILp5QB+VRM9YlVjV9vn
vo5OJtUwvETwVtBpwgs7ud8b2KSf7rtktvcuIQIgRWNMd6kXv3cTYoWwK2zVFkk9
WhjMDFw2M7tiHYXL2G34nEKiuxH4L+4rk9SN91xjglkLh6mKCXZSaSwtCP+RLekH
TtCTYhxkxJm/C4o+J/zqJWHtJnEwGt93qiEF/pIYp8bPSTBpa08x/Mwpis069yDX
7bnHVaGuYsOge2l6wx6Xp/kPeFaJGpi7AXJLQj0KX6VjZsPKeOgqpwIs7E3iEGYU
TFSY2iFi8Upld1a3+iKm+qcz2ghfcPGdaxRJLTpInzDRYkw9rhUk6iDemLlR5BYq
3vQEd+t6qIXENInicc/QNB4H7iinlpeq3ZB8YFCnLs7Sids4njcl/M416D7Si0Jc
YEECyaS0xiz2jjr2y9FS6+MieHFG6i/z7GDS/hBz+rQ43J0rmWYspmnEalAZzJYb
F/JuhV4EbBdQM/kGYAxIkbHq3Bl/+DvpUcX6TNTNGk/a6DcisckhpPL3dccW9aXA
4Ublix1dj6k2vuSzZgQdGZnLrmX7h1+T7bxCkBaFVG0yZ6bXZMJJh7o4wITyc3Bz
C67p/238GuTMLMxH7iM7wg6txs/YjUoya15OR3kFfQ/s/BPqtRQmL/hwbtM5cNA5
wZFLmtfUrMoCcGxiu0QSIWb+6m0pqs4DpwItozODzyhGcKzGIlEjg5ThXz5H6IVi
+B7PUMLUWVTxH99vc1XMc5wYSXeW4SY7mveA7YGJgZ8f3KnbEy1+B4oUkpM6970T
xEW+Q2qiRgxvurd3x7F7cRTkYyEAnQI8XaCBVYIjhi1zG8bb4/1/zYOQC1RzNs5j
ycXcDyKmHeKWQqZBr/WEhxqAMB1SP/TIuF37TErsK1UDJFpot2tcww+Lv/pnZ8uD
uK2gLDOyNVnnf6QHoUlBYon6uWbLQLxJpqn3DlApD0Bkrk3pXmKvVBnbR7YIENfu
FODaCLBJdDDmE9/waG5nL9oDF6DVDr/E9UUPAG9udW4Wx65gDIbiUDP07MIsvRUc
1SNzkW4QPW9NvUXzwlgmlTMkZJSlYzEpWaVo5qSTUUA1TXI2iVk0U/5l9WprvyQz
IENEknZ/mZUKUegsf2dXW7ufg8TK248dZMM94JUm0AANh4x0u4hkVXG/hZ58WIy7
JFOt2PcVdSL56NTfwktJCY2P7mBKDVU55flDZO19sME7yerRxUzYxF4nOeLud/9L
6eBYTY4N7IaLb/vUFqStR4HiVG02BEHVpyyt9Io+QcMdOklPKMoapGlk2m580vtl
XWhcxyP5WL2hXUk8vLQYpdIvaiOsw0ZcH2jpQFfn2z0DLsCvqs7Z98kUDjWV1REt
ARex5XK+8WEFjYmHv9p2F6OXEqe9RrDSnZMDfUh85NY8reBGVuxIfFYM2JB0DAuc
pEL0AvH0Jec6QeV3e9GLm1ALqiwvwQV9c5abG097lzKYkf7CWNict8Fz1OGq/cV+
b2jrp+2DjazqUpYJCV7MJ1po+RYkY/0PTKtTivexIFiTCyNuXTl8CtCNAid7UgP4
QTOAtZRNZ0KLU9Nx6os8pbG0EMgWE6LJzYhiA2zacxmTQMd9wVN6cFVfsKnASYs9
AEpIvf+I+WdTLmbNlb+JndGsZXUbttkG+NEaBwD9zHDUybg5dqvjJgM2CQShrKL3
lOfF8u+TT+wkM4VDFl42O3dB0Qj+WP15m0wc67QDgyVoHGi0b1t04H56cNVpC3d5
Ep/J+Bdf3nVQkmRaSvDsP92ubxevSSVEEnFNqStS7eImzTOIgekueoCp6+8vHuhy
jC1a9Bg2LwULuM0tdCYk4PYlfBNabve8pqb3IVEkvOenpTY1zKpl+vTdxKHJ+S5R
9HlJUVj23AVuvuwiVtra2wnLGrIweWO2xhyGedTJP6Shgh7jSWVSivtU2Fx5pCD4
27ZUKEiDeYuM+NN6m5wQLmtL85KPUJ+XXS4dVxKEhDagwqV638POKGd6XxmrfZBg
YR2HM/Dlw+YBqkaW0jsHBY9BaY50CV3g78xJuTE262mZf/gMizQ/TsaSEpeKpWqR
fcEPyuelB78snmehavDpSGADIXn7c4FXMV4/HElt6y+uoY0tTMpXGw714NqRJ5ig
IWj6FDk9yEolXeJBcjoseek7WP6KzMXhAt4wN/F4Q1rUIN8x1JNJKP+DlaHGs02r
pzfifehQWjAgjXEhu4sT7+jcV5RpDzUUoD5/UyaEk9rIGj/sEIz5mSSZGXcC08ES
8WoI22pz6rfq7eJ8hkz0Dqw1p5C2xDLQPVMnw3etACRlh2pwvplyPNcoPwcYxfwT
LIzYvnzwclBiFXgxLwrFbQVcSwOaD8hgRTukg+6Pr7BAe0W1M6pkpiE11wSY9b5O
wyAStJC96h8f9050Fqqzua3DiBKJlqVy+vnmIcURNPtT1Wxj7ybvxGNjxQf0+Y9/
67SPDsozytGrsbQh64p3G+QQNpTtTyDLiOrvHhUoNwRboz5eGm4WBORwB1Hu4sJy
2HPdEdCFD6yOLnJgFTy4ZR6Amm77iFwfIoF6Gb9M2ExuKdXcv3hVz7Yyb5lHHIht
aZ/dFAkNcyU+A3pwmslHcHKM6lXJDTrQet/e4a5fqntZHXv3Fqo5Hgncn3HrnVNR
uIROo24EJDHbV7oTWdNqOAC4BPeYLGzHUrnhvQOjoDyfRMrFjTAceaqaTSvrwrUo
4WUVhbuXTh1/JUKALPfRREpw956nsnH9OFUUDpBhh0o8OzIY2f6lcYhx48sbfxA5
U/kH+pTJvfX1SI3LLFz9byGPbb9VFLq/bbm4jWPhjx8BDrMjC3NQ/sqm2DDEKZ4D
WgCaLyOAYXYNwsBMCZMpYCY5Q9UHTolFnSttW9FD7m0q9d7yFfnAnRC5riUlpt6b
xHxvD4HImVdYndyutC++fgZkJu1WNbiafwUbFcwUjJ2MGN8s//0zsS+cLbZ12Tln
AxeBMbOw98Fl9iI71J/0qsudEez5LxfE0QSeGN/CkwuI/5jHD2aC24z5Gr5giXcN
QsnjgYzcMn+nQ2ujDwCSEReOxK9mfUlUdUfrCQTAoJhHsRa7zavWe7vXinUIjkbX
0V0Si569FbK2Nq0nI2TwHb500tnR8fvtWGCgi2n7Wz6CqiJCLOX248HTOjDEw7vb
3FF7LNFLZXTjU7GerPPW+cITVXSmIgQL6taW5mUkG4b0ydnW+owjbiFy6qpfNLPB
DYS43tqoE4QIQVC92rAhWt1ICllII73t2Hf4urAn6xtcmmXFC1wgCo9GUQrxGh3s
v0tFZWWO345iUFTciI4BGdtRqqFHV0g9FSZSTVAKhHY/GrHSROnUjtDO9CvDo9Ed
/UMuuqrZEe0KYc2tBB9FnAnoC7eyz0d+xJ0gHqEn7NZn0dR21XWIifC7YFOvPht3
Ub669smlDKBpdvdg0pay/LFXIXCeTjmNltvH38PlxLQ/jdArBLexe/uj/Iw05+oV
g7vGxP/oVBO1yU/NDVj8YblZmlFpx4E1iHCEETaJjrVZ//Li64ATz07wqZ0x9GU6
LoIjM0i1Gw72Xxh257PR1/8odNifai79xrjR0rpbnp1H3QHliUqhjHiM7jo0jXWu
EtE6txigZPttQhIvIQLq8t8ArHtLiJ9lNZaaHmVdfgBtqLznTiSxQ4C6IJbPy7c2
FikgnYIn8i1XNtFm9Mdk9PnEKwoTN7DR1GaHHASesP2ctQkvqegALHj6sq38zvh3
bXT1+h6iFfDPJBD1a6fxI8eEZxB7IRJLOmqndsgyCfGsAN/vxkBx+cztetPszfPi
2u3i6CFK6N94agzqj+1b23KZ2nwdU/c8H3LPqdJtmB2bFXUA8dZiGaEkrTVhRvoS
WHDW0W2/VOE70q8i+uH5teS/dZVKYgkFKVBacmL3W4I0HI6dCfrUJAEJAJHh3tkO
CwuWwPrCszuVYJp/w9i+Kg3cH7tUfR0OrTeM7HGSZGHY7LlGzCL8SAVj61kC4rQt
kdZs8fcCgXA87Yq76/Ba1GgqqCQhVVzKn+72BZWl8KlFjez92f7X7OkjB5B1He7b
qStHRIfMLRb0QVY8nP+5e7HtkYcDkvqL9niCVOxNHJfGrJpJ3zwhoqk1MrB7hdsW
2Ga4DzjkV5Vq1m+z3lvDxFARZuMAQREoZo8JghufcM4GFmMAK99vpyLroET68WRa
pDs0RL5DkqVDpywOdmOW639xQEHQSaIPL3+GvRM7tt02lLeVG9mfvPh8+RfevM1J
XQ4t03zgYrmHgwIw0ewdfCvJqpPFb4c/TVjzcf8ZzXxNVWW8uQMzbm7T/Oks3lVX
ooonQSotKowHtzrEoWvLMCycxmPee+bcUoIpfByBcGhTNuaW5fAhGCZnFU6C4d1B
qLOhTEl0LcV5ft61buKf78bmYcT4dMGaIft2fFIDOY9bh+EIzqPiDYkuAz3AdIr3
IBXZ1dpPjzGhbFDg7Sndp46svMNiArfc5EaFJr9Au00CEWpss13JaJEajMkpujpT
g0VixSz6SAE614fMlKORI1cQ4do9AxJ9PjV2bhvBeznyYorTuswa9bV2pEjKlHtG
dGZzmyUmvPazhZxLZfi1jdJWtXvvc/FWnIAn5oxuk0QGyBJeB8K+zFUqLvQLVx7k
wVghH2QyFaIpSo46sVLHpPOZbPEoHg0W7cwrnm4mld75imWYxBDD1HQ31x3Bl8s9
IU2KGzSnTJ5Roo5s9mOUK0XDAWIDlx4LsSzs+F/qjUyZSjp6wDTkeIoo0A36lh/5
D74ICG9b3fcUFkiy804FrgEhwhMANXRfpZ9W8YH4UPE58dj9fB13bICx9gO8e7WU
p30iIhvZr4jihR39xN3LFvxQB5KPTwciAqo6zo92mr5Ah3CM9c1XPL1p61/CodHg
DuCUjhB8eCkoS5LOnITOY/2j8yGCkWquj5AbjkBOHqNTT/3PsspY7sx4MVSOxAZJ
1eXyPa5B843/sylLJYN2iUXjgr4+PEeTSssxEZ0yPuGmWMTTaFTyAEyfEy2/X4Pu
/mfhB9KCd0nq9Ho0JCbrcxqCxAa+i9h/BnBh4d4i0GuUubJcyEixCOyyw8202Xwe
WAL6z4+9BCXjen3xR6OTi0QjN0p2hpAxoUMa3VgYE3a7MegDcHXpQO3gxv7oC6L9
hNkQ2DMAER0B06VrN/U6ZPT7nvPGgn/H64C4Cr2pSDI4Gm14v3bHnm0fNImrV5HA
uFq9nkoYl6DJoShtBSNP/oGiQEzrQa5uGcSsGRSBtDFp+G5fdocMLPamZ2sz3mtg
+TrldGVSAIrXG0NFdho7uqsZGc1ypto4M3eDabfK9VZ9rJeaDCTk0aioURmqo8p/
CoNsGjiks/pbpNDZpJ36qHYZ/4IQylWUbW/7sV5bnJSAUv3NcygT2JafjKY2TVBi
1EsMJYWe151VpweSV9KEZLwwoqhynli/vfH/WVBrEp0WA3e8SW+jEnqyxT20nOmx
Pwb6QWRl251jqfXZrFYFKZSbMFsfATl7V7B2n95LS1FtHAH/Ql1GFxa/NQ9AXxGU
0VTy/lt/vMxjNP/dHgvUJgZ0hreL+nonYWFxJeCdcdQKl/SWbcERq27kyTCL7CAN
Wxd0XVHPuJHc+s4hKkUDys0+gWFgAAX0yHFSywP2Xn2e6pL8WCq33zllzMdEffbo
EQqp/DbKyJhzTnaWSyiEhthbDSGA82U72Sq46mD4/Hmjfupc4U/a/wVwXe+fNutE
MsXL/rewZz1ZrRuxQyjAYlpR8MdeKYdkZbezTAYcyGKOwbdYz9CQ+PHZUQZ7KMLj
XF1Z/an54FJPJIXWWrNixKaO8n0SCeiaItCevOJWjfnbP/Pfw4vAPNL+bJxmqhM8
ugQz4Q8YC0gDnAagTfhtpJcHWK9qDD+xtmKWaxH0deBtafBx2H7zKVkoYstM6Gqt
WIqDfyTHnGxrNizML7q9poTeWGlp1TcCV8HTUIqiwzlwlP+KcIELrz1wGBuVbif4
oRGMwfKLdFF3hwNSXt3L16PT+ooPHrwRyh2YvncJGl6iIhs2zmCdLvaCqMLF3wf3
MPXkor5H7ib7gq48uJLZYFr1nJy4BzhVO+HS+/IdxkNw5OLI4krFUYF4O91qM8Dk
vO5GS5OdCV2fYjJIPQ8pL+BuU6TSbhHj2N5+xKQfjphF/xO87rBwc5R4SCVdJbSt
Bs8V6jtIBqmD764QfwkssWXAz+pQuuvmRP/9B8pixpzx15lFQ4dc8lc51N6vWMCt
Q4yAZKK0oONVytkx3ozqcaONkQjh1YjC9H3xVTNgZ5zrMPiRts9/h86If43cH9G3
vu9QwRUOzaPyji0v8t/fKMr/Mn0q+LuELJNUAuLG0Nmvn6uN0MwJDUiigdt5/T1e
n3f0AtoiTShO6XBZQxfGXapEf5eYu6wakdn9P1F+w2ZxBis/IQFy8umeVSuJTcHf
8BcSf4wQOSe6GHkIy/bz3hE29fRMkqFsZv5+N3HdMIt6lqFa0eHoQVkV1qQG9qXD
mKMkE39nExGoCgzol9aYJTse9+iex9lFSdjnTWlmtwKheibeZJrLzYoTU9dSAP6v
5g0Hf49KIcRYW5PE6gU//ytsdHdJzj8oDQZrgonRFQ1XV6VmMQahVagYqzpjOnJd
XlP5wwwJu1F11pPZWGwsp66q3mSvCVW6z1Yr9eRrsLdn67I+4UeN5F5lfsdxniCt
sPbMxjJxmhJOGCa3GAKIN8loP6mLj3XypQNH088CWSxUxrZfPT0WW0sdyoQRcMy1
I9PD0QKfckuYx5QnuNW34yRkbCglrA9wCW8xJLgURHMw+K8uCg0dzL8NPlp5Unmd
Yc/eLdMhgnphhBbF9ttMQOcIhtDLSBETF1a4BDO50bbabzUkztZXEp2PKrSq5hp/
N+zadSwPf5J5nenPG0IL85aIaoZS80apZnZ//eoLedemPbV5iU/QQJA/oHMQ2mHe
Yay2/Pg2lvuOcXLT2SKOHfuf6buuLgM2Vq6QYU4i+h+NKv/S287I0JFLHgFUxf38
udEyKlfAyiVa+lGQV9RY+AokG4zIkuzcQrhksLOmJ52aY+thAU6Bj/mYplo23EC9
R/RZFR1Qjd5q2Ho6t/kD0IfWcUTKqTTLI1wJmFPmNPen+6vKbyc606Jklk7xFhBF
dYzDBpBxgNh0M5TmkcieU+iMesPsRsstNCiqWxdLRIyGDmdaCB6NA84u0Wnmp3Uj
aB4Mq8b39ohKkJD1gQLkR9P+1jNwcTINZ/d6nZyLdMo9BYj17Xdg/4p4FS0LHx1n
yVuuWsHnN+2tvYJREHC2y1rqVg56Xn+GpXc+PdfpN2+QMxn8Dn06q78HXhbHeIDp
UuKZgZtgHkw4xwN8qENtP5xhu+0qmUsxA8kEXTG54l4lK+NnpTsoGoR9N39aINRO
VmvfNQ7PQM2ke5HaP2z7XxEXayScB+5go01YvemnOFYpNxhfcckNLJqCFV2kgta7
p4P+fSNfIt0COtVxrWw6XNbPUIudR0bQIH7MMVsi9awz9DYxCS/ZZ6VlDlAC1ew9
2WoJGbrfA9mgpwCxKAzJ06Ab2rkbHeC979nW0bqfYVr0ohjMJmByt0UPnVJhouG3
n/DR/D18eNVFMGgzg8KQPxwrKlM8pdObVfZYfUH5zgINmBmZtxEK4G+GWkpMd7wo
wG8hWpPhrCIsyG4QkYG1bVoOvhvzHhIaopdTfBvb7KBySsGbLluFLXJkHoKBl+35
kPfDtMIW3yzZjDiFDJqQJgwT99wpqtS6Wof5fnGrgLLt72ZibexNIGnTocHhAUim
8kG8ck+fuIj9dnbowX6PgPbcKX5dH+92Prcf3k5wEqTJwPJsPNJwdZWrlt2GtRng
iJTBkutqyAx5fWEw6+0AeCI/Pwz8WqU/aLn+VyRBoGkeZYR534WkyUMeTdIuztr/
r1+40szbB5AqtnhUlDv5TGrZmnw8fcXJIpOeoTPYHvyer4YQuyk3PiEcIrae9lFo
Sc8KkfI33r5X3LEdXATpCJORdSEqX/ZeCtw0hB5k+LyAmaWkqOR5mlEXOa6iAKkS
POzlTQaYdFwwUPCItXfXypLYKltZ3NNyRpeIe9AqvFPgz6A4fBPzUzRxQjA2EEqE
bZ7upltt78s1U1idr/13T7gprHUzUKTWm9n0J6fmQsDhCdxM8bdlf3MKQjWKVlqb
uExL2vdCfsz9bC1Lw9Hfg0Vz1x1rTgYQhCIoDaRcUiKuLIw4wGyTasoETKalYCMj
nKkz0rAnYWWG1w1AH9QAQYNr5w7IqLVanZ2kY9Qe4b1XtMuperviduS98ofOAwdM
FA1h+SJFI0ltasKQNvg/4151SjJWWrMZJrDYL2iTNlwkkrSmDiNzu2F2re6B0lrE
OuM/OEsUG9LEJbHTp9Q2deJ6NtfMrwF+7OIqSIeuqh0GIjF+tlwmiUg7Bxy7/Bl0
wuJLW6ODL6dl9CbvJjelQ1r91EGYJbZMuvxS+wsqKVzrlbgwdFte79x4EtKF+HBb
4ZAzp19OKSYDcjUUTc8KQNpGNNjLnttdPVkay+CsLeNntoNZikTpJL6tCHehyqEK
oYCvOnd1kYgSShPKQgDh2rjUFy+ZNZTDIkyZQWiIFyL2YrYRkQxv7lTtVjl6LrsQ
Gpj0ZkCPDUwZsGs2wUdep+T9FMFUf0N0xghtxYOZ2ZRKm5vtSMijtD0SltXKwT2P
a2oprtVFyXmBXON+sgUhAdipN8qF7jtMYYA4L/5D4Sts35uK/k52/w+WZ96BDvot
E9U35SauwR/jHIaiAs5fDQ7FBd+5rUqnl7eAoS1GiB4yAWQHB4e2VnDK0LakO7PG
95DVLqiwTXBrTNovIZyMlbA4utyPLzczB8km+W/LG0/FhbcQXLTQEi1QSjTJKRsS
PMVp78uTPFPHoSvseokSAArUQslAsLvPrUadKKBCDhFgs5JDLYomy4VEqf5rW7RY
ClppR6jsoVt+DXi83lsDt2mBw6UgiNTUzDec5Wpw6fBT+2mFCzRSxKYL2Dgiw41d
xXT04rH9zN9MdIMAXiYo94szd539Me6iy62Elq1UsKBVAhUf+30bK64MvNA0Z7nO
XH+GpRqWC+PKuWD6pvhuhskacXysBa4Td0oTQmUHogGvIJKH+SLcj2p4oUa/E7xR
ENu5TReEqQbqBuBAFB7Fi9bxsbCx2eg3NjdDM1nTBgcd8Rz4nXdSgBegjgf3rQ/x
Jw9yK0QoAhFXhCq+MgMQQdHHYrcJuB3LObLywuADqLAmymgrHBEAMMrmLB8T8jvj
397oBQON9I3lgtx4J3j2cjeSHIHRCa/SKJjUCzkCdz+pE4ZWfNXkEOYVHHIib+Vv
C/fvHB3Cbi4xYs8oxzgBI0bJuflnmiykZcdasvGJpGx42RZ+ddojx4z83NpOpPty
eC364mxil4pUPcQzMuDCnXiIMOeP38KJrUCllq923Dq3yYSCGZrQ+0B9VyMxDc9H
4KhTVQJMqUNUrCpOJrVk7fdG5LdraCWTewELDNvbO7omymTfYv0AxEL6hJFXfSZo
PsxDBgAYOOhT3emJEL326K+5kGcX9RNb1Zly9/Ac9dLkjUY53Ve40Et8uFFHiQJa
RLmYPIV3kxsMXC4x0gWH/jgmsOtimTOwNs7cYnQEV2zXU2MLKIBOIMm8w4EnZz/j
D91f6/jMNyVlFm4kTMwXrG/qiT8xkA/oRdk9iyBakOdpsPKt2cGzvB0W1WCor/Ss
T5Eq5oYdTeh7Wlh4q6tYayX2Sq7Dx3s7poe5ct8E/O+C8PhpBjq4Iv3WotzjUszu
xI0Q9drc30ZLG81HTk2NTCx5XsZvPJy3eSHSl66DhBqbjghgykqh9ojhC1NAQd7I
0S4YfQTPQkWFDWs3nQ/diO/3JLIiV9e6c6IKwGySxZMrH+90fZXakdV7q0OSecnr
qgxjMRpz88hBT/+lj/XZFqAHooGXF0G5pFV1guTcp9MNT/neLU/7xWhTSIEw7c5L
X3XcANsyigyz6+w94LHv2oDJX6ydNRDSSWHpTqw3Bq5UM8fAYgwmShOGpT94KoXI
cTEUxuP8ey4soqurbK5Axd4Fe8HhLfnSDa4lcKP55smJrDKdaxY3hjE6tXiUr7e2
HKTn1pr9J1LA72Cpdx/UaYyijm8pMwdR+NBaIykjRutCY0BAB3SGDve7Td5aIYKF
QHn0NkMNSZqEaSj+60LbojoS7yZGD5KPLLPol8/GPzdAER8EHlwgnPVCE8pD5rA+
LMFM3cNVqPbPbcKz5L0C+qrsffn3VzgWphfIxL+vRCD8oxfc3pCiu5qTLjhKtPMw
NDowbML2DQnmG4jozgD06jFzpUi1lNMHwUjMJ+LzS7HmdFi3YMYr18oCrCIWVC7s
DAyjO8v975j46UWgR7LILB4zp5IzBWoaepdJ9YLLIubODFSRmLQFqa7Q2vS3poIY
tSqpplkDkz4FkOpKBx8MWgqjeHHRRTvVMsteA58WclgLBVoZWkjdcfjNcUg0NLaK
0wpmxgepD0KZKQRd3uXh6bhRlaGfS+nRdJD9eI5Q43eqXQvJEvfptgWq9hnsRpWg
Zv7aF025zbMRVIEF9DmIekUPmnWEvVKOBkIF1UiMPZqxhHJfbKG00HUrehUClnzs
IwN8N3Z+n7yQLt8D4L5t7hQPKnFeYaq2kSIR2tU9PEdHBeIUMHaZHGx4dI1ySbIt
JaG12At8kUL4F2u1kdQOEabbtSgfD5z0yj2OG51PD15IAQ52Nr0W6c9DLgqNeh47
0MTEiU9QtfPU5YvBzpD7xf/L4ZL3Qo3v1doXmZSGkqMYtz+pwdJuetHh5sYfMaia
nA7qI9sQOhcrKBt7lMLuqGoSJCXkQVqVMDgyJq4Q/NnQ8jMSjJI40Z9IZ+2Kt0ZD
oeUgm/YipR84pm4Jgfsd3/3dikCBSJZmuLoutHKqP0StaRyLSyRAEBpzppZunR/m
0EjOGaYlHckjG/4hM3O+PuVyy9sJR34MPKBroFEspbXYFzL1sNRgngXuhcUNhfu0
CS4Pks4X7dvwJxIsk28YuepGQwdrfqtI9F6IWy1tdwJVR5PVHtYJzxqe94O7iH8e
r6S6jaul6xFy+3NyeF17le1SLf4rISMLCKiWI4VmYvVnKnAOIJiv1vWuBerane68
xgbeXOuSYdKAonZ9nvlgxT3XcMv5Zp4d9iB2Cyau5PWmeYcV+rWkGlGQJHOuty+q
zCJZz9eE8ititusnyz+zGfCxnDrtUWlWCrM8q2OiOgVBuinXsJoInND9dC0NTwia
DzcGqf3xrpyOJ+v//U8hV9tUeRLYizp5ZDyH/QNPkxj3UpDGJWBrZwMEjgXVs8pN
xYwWzHfM3mb/NN2iWX+tRyBFfyDjx/rvGrQCABh3YhhgN6hPj4cQlXuY3mpVk7c2
xQ4gOYPYYVTio1DVBZAGqFRI/lXP9Da5emuwhaUnyRZwtgpNK5cePFcxwgQKrAi5
UzZNPqsYHufF92QUYoV8jwLfG1QPoiaF3Vmq+AiIedH5JK3H/Bj1E2UIAwuP5BPc
7LhbiqJKP88PVLcE5DVtv6xrKttyV/QuXkvwQ5lCXGtk3V/xAjBBGOTqctVtbkrd
Wi/sYY6Zha7s+yHUJ02BZQvl2NficodCm9R+xabzz7FWGRwcMpZq1+O+a90Zyh4+
wloPQXWd+1Jr361RFMNgWCCC3rqIrehMvjKUKt9OnYBUnJwhEDVqZ4tyBGwRc6Gy
I7P7BUELiPm0kur/irMASAJH7B0qnmrRoRKAu0MRz+Lqrcc35Mj907ieW5OkqKWf
R1LY2XIJ0bs70cH1dIehTaJ+L2Ll6GmpFER2t/PPPkdUSkdH5zJwXKx8of8JpZ3V
+oOra0qlvN6JSQ9FQXhaemNxboTCQjg91/wr/tRlsC3tPRs4q3udTlir6qUX3z/Z
yWhVyui1KkJPVK7vDUnq5VGN/PKhX+QMC4+xe7lQSTluL1VcYTGr5cI3Oa+grvA5
rzCs8wnaJejxVZqwUcQkVEkGNQ/o3KFCc588j5J9lPfaU2EA0wNc8Y7AqsEWySMH
72/a0vHQSb43lfCbJr1DLDdfuoCfdGviPwOId+sdYMXntiTuZ3BK31MH50F0yDKX
jEAxVzVI0MLdLM712+WtaWl/lvLW6TeArdymmPLzW2yQAba2h4ATXXBzJgs3tTvM
wH0vIsrqhkskvNNK8X3VAT+KK/sSsy8bHHlGQDWyaeOFeejnOqqqwL7H3htslj9A
lBeqPmjGbMcEXiOezxIm4ZUEZQJ8O/07iTj0svK6dDN1Pe3mNAMg28K6PhkV1J2c
nPJOzuSZN+49obLe8uE5kqcFdj3ldrw/lHlZhWTXDFnIjn2HM3aSm8e3gY+C2MW3
6PD8xNYZoGQmDxNT2uA2yHTOoRyApxuDkdA270DPZhRou5VgY2JPqW76DzN3k03m
qpuDM6ffniGlNcHrPLfURc4W6ElSYZUbZzgy5/sm78QF0Ya7RDBew3l1IAihH/gk
BSRGH2QiRvNS0+wq9kr69XnX5p5luW0vJRXJ8DzIec8KnYbAhrBbasTZj+OiPqL2
Pmu+82qBQADpBso01rCCVJzk2L7ZyxEDl43Onzc0PlvAzLi/JA2uWkLBXp0grfdi
PMyfFVlIanDS5REzDw9PnhND2kqm6q7FhtSwfk6E+1q6hQkrda525KmO0zxybkQi
bdjBf2LSGPNSmClrvYV4Ec9wvzue6DogLJ5bgewR7bXy3yBE8ifUuPGdFYH97kLa
uKIQev1O5YsmxN0XQTdK0l5fGiFHXt0xZzQRjTf1Z9lFwtJIz5Z5Pex9g+yEr7Ht
y/8tOyR05+Q+dhqUfiz4Fn7UGMZ0CYi6nI7rWdfk0WdoNTq6MO+wFQWdJK9WbPg2
jmPe1DjMfv3D5SeXyFBdRSCpt5yKqZYKh6+ukOYNKkU0Rjti+8+mydV6XQH28GX8
7O45XxRl/G26fs9qSglfGlCWi9A2fk7e16bkH2EkskDZfkLXZdVhre1ckmQjjnh/
lBkChbCyrJzDbKUMyUyq482L5G82eFM/TTgCEPvsXoufR7g3PPhHjUSzRKP06T1i
NfOOdDCiKA7CeYi5P8zpFo3ShTtAHQUpy7MhV5DyV1DTA46F6/fQU7od6Kl6Sh/Z
Z032kFLrosq125JjKBpdNq+znlvsba6B+Jgpud/LPd2CcyOQuQ+EZPAqTpohxNlZ
pRYVd5c/xqD7jG0B7C5gwGX8jnxN/Dnu1O1Vlpnnn2YoE3uz9p3fFdgBdo5sfH30
020W1oJR0j2+gUJXSLPKiodUNJgow2rR81OpdXbgSaRe3n4tNuyijToDDZGpsYBs
5FD9CStaKo/h0rqTSn4bXRrqNdnJ0/72ciczlQ6thDk7layU7DS1KpPamTgH5177
JJU+NNHAPfmgYC85PQTo5NoraCu46YsSJ/Kt/nm3687xtEVxna6ju+csFSvnFkik
EnazNJU5xdhthFtAnoR6tD2qhka+xDy9Z+zBYmyZ3vLKZ3FhAUp22hSD51aoE882
mbXyEzOKwqgWc3ZTkCPuh43dv0/uAxbDafGXQJeCCd6Tp/AHOR+2AbDJkeNILpo3
nPEsiIJhxcQPGrJtq0qhKpukROj3DUUCvRgXKi6ywOlN30BheEAf/Ly3UU0BI4Qx
HZbjITHvgr9tR9oANLR6LJEFMG1lBni/z8KnGf0CzctVmMXjKn4Lpn145AzuHEux
QD63AaMg+vFgGfBvzHIRNhNqXrSyViHvHU5prSO9m/UQqnCiqFHS+donC89hHkAC
ugkDWPl517ZKnJCPWHzquSjMeYJecI5N6aNWrshRZCMfzBIlFv0MosfLu8fsBJBi
ocRfStWBmN9w74qftd36U/j3iGde5lo0d9RFwry2CXUiwBRi/dhvLdNFOcFHv2fO
Lv5BwoeTaBvpRk331lEmKB93AZOD1NiBAxgaUV2aqjJ9nOZYaSrVQbVbQt+Uk04Q
jSTwcQKoOaBzcitgmdfIccLtE/B3BPuR4T7pnZt345Gmt0umi0gWP5Me2wVSFq1n
L+IRy3Bvj8RR8wEqDM8XjcJszaT2QAD6opHFjAVQfXowiOzVRv9UcGrab0D40tfe
Dh4xG7JmRYngemvXgX5Nd+kuF2knDSzC4j/2gZwVkErcRmkxxBc1gXYUnEcIcmvS
cQFzDZMMOdP6rpfL2dJr1DW4R6co+IYaor5AA2Rp/POthwEz+JTnFyaHU9bHRUXI
isDjZwxWdUHgl+9nkTHupC6WRS3LxIqldXO+7icuMJdPt5nu8BViGCz590u4yaVA
1y18ycuupzDYwj1yuvEX8Dc2gju+SZmj2ib2Xm0ebz6Bcmxo2v2yekn7iTPYV9k9
AhFi29rb8/H3jzkLfAdc+Mh0BSR6gG39NuGMI9W3LOd6HyizlMah2GcxY+XUhjGp
dgrG+4B/hkqw68/KNucJ2nQgzlFnHyPVpHH/tMtPkXYraYiM3X7rVoScUHi93xF5
bkhwqkRadS8GMzzZKrdN/7/Hiq7e77cJN6q9nbE6CAfUU3PeaSvushtRPoG4K77S
lQQwoGk2xNFk3tmTmVg+Cd+upO4m8Cf5iw9hHGWjM1FvY+kK3e1dOSgbR3dv9cdQ
t38dgVMhT6LBQpGuIkSt0ekQNy5JzIew5wg07sE7QTzzsBfPIJtWTZ7JLBAyhOJT
ViE79klzSvobVEbD5xEA8evH1ABvxmk85dRG2HO+OxmlDffIsN8Q3CMZbR+C/U2G
vxBzzGLTzn6R0hNdvJXVqFKDD8bbWCPH/d+88Ckez7+N1jryYQ4xz3dhgrElK+ED
DcLi0d0aWdkz7R/IWRhhXudSWYcQOLt6ns/zg4OBlAItyN3pEQd6rdAbFF3SwF6T
juTs2KvpXUWROLd0vshvF0opOF2F+wq87bWL55AB+i35sC4acoIOsIQlzopeQ6JM
sHJJK9US1LkYaFmg0W2MiOfGc9tnx4jsGUWTIFvz2zazHpLf43Ed5ZwoYvEaUVAQ
qs5fqSPDOGFEtgGuCYwsWwkbLRLbTrnqJqc3l7QHD6xD4QWRELsiqxUGT/TeG0U1
TZ3cpIemxCodcHKvE9NuR5Uy+faRT1cdHjqfJYhyhKLlU9MAzS1DnmLFXyF8pgcs
oPIHY269vWyafWs38g6qybvbKBCAd3Llk/y0Jb4P7oRJN/X8IOw2A2QjRO1743J2
75CkA/dizpGLIByP5BO+q1uyMu2fCPp7mJN1pLRyUynWHra3IsPv+pT4OJnLiqqz
EgqnnmoGMUtQkn2oVwsS4BS+SP8BolbRL+jByGlxM+RUI35nGKSn7eXpc41CWeJt
fjHiy2WFQWuWijfWL1YwvDwOHQDjfbalR4+mGKfylkYnRaf3+iKotkaqxM+uvPxl
FmpXacnwS68Be4oBd3kzJknigmdhG7M5YohQ5YNQXhMyorkopkERE2VCG9BL3BqB
w0D4rLB8xdqfuyBD4W9BmFDuc6jhHYRgkrKqGxNh8NVMiO78v7mHtGOrk1Dparcs
CXvw8apuQJ4wtH3ZYZ17CfrKk6KyPmb3XQlaWto/36RUxR5pRop9/PZuz3rIhaAZ
ReL/mYaxfsaIs8DPzysuKnxxDhZ65KfoMy8H684M1kx7nJW69grANux1AfR1s7GN
mActEzOqFoJF+jAy9fGodCPXaTaph8V057GgjTddF07RG+kU8XrIYNTdLd4ZHfLt
x9M9x9gIBzLQdL3C2RU7z7TmgniQziOjusX+R83tfGF2yepPghEJzvbujiga5kae
itFsZ4K209QutZl1EhOPThxjBFNdO55a3ZBJOfsCXcyF/4jox+sWm3M+cXEm+qIK
yFTuySv5l5ybSPzv2JkVY4qhz+PevSz6fvZTzbIfN2F1cdqgwEm51arBB4t0moCp
SC2GStrvIbisBACZ2I7JpePqDjofz/t91BhuvAZ683k1SSJVwycqB2nWnB+U5zHX
4/RopwuoOa8XjAtNh6KF6gOvFWkxeoqPDkQ2gNehJJIiSsQ/o5N8q/AEv2kysAs3
GlsS3TVPgSMWmxDbM8THlJ8w2bR+mnTqf8RQ6hrCyyFUOWWi1aTb96Rmebe3fhdn
656bRvRA9F07L6swgOxgNAw18HHIj96mcwwS+gYCmM+RslYihYN3FvaHxOP/X2Qc
NHMF2D8sdFE9EyhZVlxqx/MnFxDpgNiN5+XdID8V3KYbn457ZA+s+lAle+OUL8wd
+SO2/68pe7q4sG8H4q9vPAaKIarVlyMLIGkeZlWrAZZ8GY1hCP4NSb/RNM1397Nw
gvElbX4UmMY23sIYCz7ySZcfE1tm1YxNWAqdWDkJF1KwgaqxZlmw/h8Z43EudKkt
yzyNw5upTzYfePwQkPqUC/sp+JMwVeVDULZtZ5Z3QPa8w5veBv1y+dexDLm02xGs
AwDTtiR0TAiwqHDusRj6TI/pXzmMKH/4VqaD3EUFyGnuSWocWo3WJSDo03NIwlrX
EOetpGrJ46csi2EIT7GJeav5jhV8BSXj9pDUi0EeYbU+xcQ0SAezYBwXD3Ub2wD6
kTnOV53GvnQ1iFiNDaPZ+1Gb3Jtwm8p5Sm9duiU671AQHTNyrdaAU/mgXyPm3l1s
dFmUMQhpL2DsMW3b+qwufvZJBwVt8EwtVPQwbU8yoSZne7EHVtFef0+mKNODjokv
gygjeZqm4HQdcnlQg+Nav7L4zSYS9R186ZqE6vbqnkbXhYP4JxPan5o6JsKDQ6Ip
N6ECWPanMxE9MpZtgqpyF01oq1Yai0n+L83Re+KjQczanIy7xmtSfE6PXW5bxabW
DkckWuQSIbLN95q2EByMFUVlnOQwMvp+a2irMdFIhpuFYTylQGLOkTqOkT5qVGjB
OgTFUtepTqSnAD4cuc4BZzcUyn9pitdVP4v8hrp/a3QEPCL3hBmkoqDkOM1B8UAL
qx0aIYp1TlTiBhz8H4FAHNmAeIM1yj+ZOXWWCzR/RX0rlSSyONahFw9xiCBvkFeI
OW8dB1S5Jujekx6/PZJDBUFOJ/DGIBEywvfVlp+Tx8abTHO9BQY6pXk0HVdR6Ee8
iSld9Jxxfdb7uftMW9cBDdCo1eEy4Gspbuxg9PWevNL7Lb23KkTqokptnJitutHK
GDHX3c6YnGAvv605Ptw9wP4sXlTNnatpMXOku+wxUzJDX4R4iPgjUGesDFBbPlln
4e0parsBh56sYu/uh4vvDlXHx6IDdzo2wCfRTz1++22DyHAwwSp3y6EvmYbwJNbC
Cd8ZXyJb8cnMgnUNGE3WiowK/CxEVTtppEBX8gHaUM+I3Z8jkQ/UMHMZ2L+MB9Fb
RTgGYFgkWf9Qt5DqbLGME02RZ4cWJ1HSvCGHoIt3GeqHAE4hLDV4gUeMdjbYuZrI
i539vSpZtxONhK1V9smdHRrAzV9WI2MXlFzx50aihNf751KhggnySaw5MnJcKgvd
KK9YHiJ+akT7yWMdRp0VCFHI1ox5T/zpTPpRYaXklbbApCz0nFj38ZlN4BOqKH6K
YwQdKdNw68T/njT629WmkrWLiz0sRruVE10Y2v7lKGiNAGmpj14IPD3h6HnJ1OQA
SfxMBtUjwe0/LC2Zbqp0rxWr0zclaxxeKF6hYw0VXHIsV77wB8r+diSFaPTDzez/
7uG+lNywf6Fw6D88zJ0lbDsGBjPVA8r0eimvUlNpLVKmH7Q3gyk3krHFdUpiV83W
o97ShR4g6ifDPt7J661j+LPec0LKM4fr7jytel2smHXhpXdT2S1ujJ/jySQQEShD
3h7sCsUlfNxDnma8Tb+/wMR7gnyvU7CaOAHs4C5cu7jIpSIC0XdsmT3K++ayTiXD
RDnIX1TnzM5V+lX64/hO3/r4UjE7IbHYqJNbKzRN7BqF8P3p9V+lhu+OEXguPQiF
eKktt0BLL42nO2j3mjB6GHLTKQrE2U9hUFwZNJpIURdMQWLNX6SL+VgNcrm8agYW
Z90YywkKZLOQIMUfsbjpNp2LQPZIF8IpmUWvk46y1bmk68L7m/16/Kr1Y9q/GJ5m
GvekEIHgkOpCF9BV2dGewLTtFXVpPXyuoY1glcIJ8cAGum2ot8Ad1cxNyThzD6jY
VnpeKgiz05wvcREKTcmL9l3X3zbkH4jWOBbmqDihgiApWAfJM/u9DKYue/dfbgeJ
8VlYYpoF6iBFMhKCQ4U5JX9MGDJZe+A0XWGejOIs+K7I/o8OSi0cfxfug4PdkQhr
ZRYrNpfUZXOVKNTQVScQ1qzv3e8wiNKifYlyi3stpm1dDoyVeKqbfBPmi8IOwXEZ
awWlSuvnCMBMCAeZh1dY59YMlKvYj3K27pjL5HE3/A50kRWgps3aw68idYaRJvZ2
Bn0WkIyBStkmF47evAMn09yhiNg6ETC7xcZIALmj4PntCgmiKXtO82Oksf5SOvxK
l2Dc5HHGbfrrisjjrU/755h2ImiCLoq/r1SgGRPof4Wo8Tkvsutxj5bv9ItRVsAA
DGW4N5YXL/2yAAcuqoY0lTtF4bWgdthnKemfUotskVAfHPYOQxnuha7RCOFCgSA+
hQb2i8dXWtdcIG5DNxz6QqT3Fb2y72HulkNk+sxko6K4r1Rqb6I35Ta7Un1tFnjw
6mxbU4Y5T7NEqDZgk+gjszTwuEo4Y5ueBucD9NRFk/gZ0/fvPZ0F7N6wvSRykTI4
E//c1hrVr6qbfIPXrBORl272X8mhqwDhVl2RkFtRq75R4LNbtOh0rHCKRabkG+Sg
xZTzpwd+lRLdF4XQVHTqGA49JKBeKF3OifKcvDc44gPxFC9Wvo1rFxgkhlcuLjjT
cW4TRLDmdESZDpYdTaowattlXPTvlvo/3v9xg2r47+b+DuE01+qw5VqXhBW1jrDC
GttQlreVF52h/suIQE3t666oG//8uCebCzByGIvtm/1FXcCEQP61iiYGHcljM1PW
dRgHn2RkOm9Ao5jJQZxXyLvEaQeSe36rdqqnYQbx2jq74Hn0OlGt7GWTRiiO07vf
NSRGEdXRqQg/v3cPU9S0NajAVLJ8ZM/DSmvxx+gsWWREBp5mk6/eq9qhW+w8RjWv
1lCIA9F6f852gnPA6jqAe8OldtbmH3544WatZVZdQ6VEcAz5HJR1rZ/npQopHuEJ
nZt6Oi7JrqO01spK50ui8oIrLLTJZlcv/PP40YuR+8cOquYP6RxiI6vSblCcktVi
fF1qSmxkFXmjzShb/BPTl/dAQ9/ylaZGbXmWuExpylFIsRPLQtX3LOvEelTX9Kly
G4zGCiG+7/Cd+lLDqu79uV+YX/w4wlKaShdfXdz3/6Z7AXgHcTTl2IEp4HFCavHO
tMfxzhINceHxa0GWa0+NFrmU4L5vyHiZDUD3cJt9ebYHNJc58CQEbWRMxL1r2j9Y
nT+xRVZiEPZYqWDLhT6/qnNhaw/ApoPngTO7t+fBT1GB1KiMXXcAAudpekXslVta
ikU1FKG1f4jQzIux25na4LtqcYiZbWl5Qx5fAgvS2lTtLbDwS04XrEf/NjRLX+YB
1x5vDOx8THDXaB/WsU28I4dZG+ADAuw15YGi013NCdC2e47tR0oxkD+KRFReQqkX
zk6F+Uj99Cycwk6okFo48aZ44inTiNmba0JjW7rYIE2R3tbVBhFswD099kLvx5WH
AQcxfd4eJEefPdND+trhJ7pQDYu4CIfoB6aFtU57aTmBDZ8ciyOe8V6uDPeqc24R
wAuKbLzQ21qfX7e8jytOf7kimsnq4xt6aQZ+pWqw+DcKTw8jHEc+CjJjaKfoj/jw
P2loDC73oHZr2OmMWXDgIqBeWWzj/6RT+mTgYWt1KxPB+DwdjJfANOpp+3lvXuj6
FwyWcoltaP08V5cn0LbR9DA/4GmSVzIAcS3+LaUCvpgjetzs3T/ajGyC7A05c7cR
//4r6Bh8rvAxtCwvQOuj4KiFZAWZMzjsQodGQrYzo/n7NsF6CfSzBem+sJXIX3vj
jOjL+uEz0A5irkDanXV2XU/7vCuQcqMfzFbMBPJpyyQ9UqQeXHk6QIFcQK8zq9xt
Hz+162MRfQ1CAL8USzOmPnNIrgdnjz+mHwL5UiQ5nIQWIz6/nc9pg/bl2lkRs8iV
bu7mVvxkB/o2K/v7YW8+osuFHoyaKqW8eeNFnIe6p+P7Utr2fCccDqg+/L1VJxlF
3t3M6+EfeVNdodeT/Oo4vztzGR96UoJFnvNMIbx/Dws6w7nDGUGelOGic7L9ONax
R7WdSSg2vtVoPO+Z2I9ZeTNu1qRWXZVsLoXrTIoTgKgri8DQdjgxVT/A9BVva95c
FYnYTJpj1mNuiSJpuoMW7ZBEEeR8usSQQCmBWEt8zqKMedp/2Fkzpzpyx71g/chg
KL8zFADOUFpVyHz1wvzoElvQULGMjnVYfdQa15ev6E/Rpr8xnVIXO2ZC0e/1YuBV
WvbPUnNzu7IQknYSVqWwGIGda04xmQDtvrM6GJ2Ohm51lo5bqpXMTg9W1opocjQh
BT5YmcuGAkNwLEPaiVZjEVa4BwAPnk2iWGN1B14c4oQP3o9tY51dQg2mG2sFV2CU
nJlLEM75935l+YLAgEKM4pun2KOkQ5wO3+jr6na5iFWghD+Us7v6R0f431Kvb+ZG
MgF4J+pZN+7F4uC6sRj2u04aD0SYOjCTig8+WCdowyzNVYut6ObUFk1PNnZBmR4g
qJR5EHIyaQHvTdQe2p6Hjfv5cj129LVjbt8sjNuRV5O/k/hg/62CLl6zTuYNzowG
a4QCIU5IE+yTC5Gl1EkTHNyadRgrSRNXGGTBSqWIxzaWka1GwRhWTk/gSBi62Hqw
u4YRU+9k9XL3ElRr16V+VBYRqT9COR6NIFPmELNyZTVW4aTLHXDu+yy0wb9F6Jqd
l1Jz1yXpQoufCw/BIFE9DMx3gvmEj1jr+ueFI9lum+YONv/AMqQdDyn3pIba4/Ae
1Dr2NF+Cgy5D3Ntgg+6US9up/+YT7JduzPh22PIaoy1jmhnLzMP7b/zER1q3PFmf
0kXdldMr8Q/uTagMKiYGJ0xErQNP3u8i/QwGRzM/2S2I8D6N05/DdHbQ5WOthXH3
qduwFY730WXNrhJ2cs4dWmQC1TWpqvrhcPXsRH7JWUKfgc8BY1JNHAvjxnhzPtOR
GISEWk6HHEEWgntkL8mieiI72pb/FaYAgbVKQw/MQsFv2XXiqZbXUC1Tw5LPPjim
vmvx60Puck5T7FacJN1eHP8ST2973PbmSLItuKLNqjrRotZwGjeSSEU2EpV5xCaU
lSa+C8n6QfQ3JYjCuq3POHm+6QEeUaQxFPh8XW1dODPWWdE5EALwy8RvVCKrdhLZ
3HcFuCZjU3/j9UkOgIBlcdo94LUizdWrDFQh8Nk9Xn3B3b967tjk16jxB0uUR/oq
KghZhwubjWiJT7YXO7yGYZhhuTWy0rYsja6Q2ETUWBi5sFK6bUfKmIQUGk83rlYz
6rUKZlNN898kqM/MLaFz9RtSDr5F3eH5HvApC/n0ukhAVTwj/DkeLO+1M0CnZ6mS
KwO10BdDo+x4eBmOEwjeK+qvPGdSDFkONdAUQZNhfHqzr/CJiaNB5Kj7XJ4mzIyL
i/Cpn4idB3/eIRdq6BQEXnJrySyAbhreSUGZutjbLfHwJaNn+hZqNAkmo1L0j+rt
jVO228RpBLIEaE/sArpszG20cw/pqHQRCMtP51ikS8AFrdNWGAMfWTimdBq4kT4l
hSTgfCGo/nv3TEov1j1WxTw2p4RZDGzvRMK12vwhAoG+3O1qXnWZ/ipZDp/NLJUK
4q9c5c7BB4D2va4QpsN0B8KbAnPdWw9wb+gWzsqrUW48u/0rjG1pnynfBklVUbbf
uLfSRYCFxCiu25v3hFZGTflrtuZfKm1FY8JdWxBJOcssLvVYi202SFhhEPTnYpPN
dHUuwLa0zF0ugSE0EyOrunOwqZzKWwDuAmEtbDzoQncH8D4RTDVUgPxM51wnztGP
pZgloc5iTgXwa1Cl1vCNBmJtlYW2+ahkZVwLa3e4ZmumfpvaFTF1BnmQ8H7AuTpu
b302y8e7IESd3zjDeDLSmUR8LU3h8SOu++B1SKQb+rAIbD9Kum6A2ON6utfeB05D
9hzZibN9noj2EirwNokxPuUzAQlGAazRLVXYtZHuWrTA8B9E+plAWAV9jAhv8O3V
r1v7PnII9+RF2ZKKD+p4Qkb+shVgWUAeO/t19Pd/DUWh10NA64rjmKw8NZ9q917L
A9nSzuwlMaLAwKUIAOHwEvZbNRmD+BLiZ2D6WJ9joUIrC4cUzZ9ai6DR6AkRDG6x
0GrrVWV6ukImdjPfqDNH0Acxk5IgsJCd4Cz4yF3UH6OtAdMMcF0LP7HyAgPVV1OC
r/i3aEaG8qhjZ9mfTlwB541Du4o0pr68ldqwnaMjaxnUSNONclG6tArw8GGbAQvS
8gLaoGeJyagyqkYbKxkuYARsmLtFJBd0yG1/6yEena/r4dLFRKJCsvkLxavZcYUF
zmKW0FQxNQJLpSaIpLf7Lt7d1HpB8isysfKVcGSUdJxts0S8n4UNSyo4hzo7Z8lu
M5eljkZUhExw+wNqnU0ZYODg1zSVxFkwsgQ6COwg3xPZ/vgbCZ4nXPrGJPgC5ugB
NZj7aT52VSj8xmy5j1d+wHbLDXTQS2mS3NHeA/rCSMSZThNis7rmnG12QA4Ppn5B
ISIiFA5k7skb1Req/1nxP566/JVCFAboJSXNRcp3GODFCezUmFAa7ofUyG0u5foE
e1L4FQ0nXKrdK2CBCVG3XCp6AslDL5xmrx+ezVF4blwL3EVTygxCsfgozMQLd1NN
2O5zU1wgzAzGdSB9o7ILgxlXXVOayBBDHbR2rbICv4fsqBUXvxGSTJBjOQ4dJJxW
tbg2RuAt6R+EzHZgv52zMPhfGSI+n/R2zLvF2JbHkHkrsgF0z4ZWcl5QJnxUfVSX
eYjojvXfb/9fKpL7sjn7prkA1ZCuDmv1DJj1toHuYvOw2Mz39LGXvUHeZMELfk0y
5tf+rgeQ/WxDd6gKnGwQUVs8djG0gm77lAf8DUlGFS4RsFxTf+DIMa5dGIR7JY4O
C19f1nsC8tyIDghbTjj0UudMdjSgY1T+Wk8tB14FoVaobJWinaKOx5cumQZdI9JL
TggcbnXL+nYEwBovD6D4inUV7xSvot9J/W+AipSlJL0xPtX0FCW44S8aIY/lWl69
fnB3LriVDL3XoCCBFe/WJsKFUoPMx2S/xVqL/tzOkNV2sURZEW2AuAnrKjjZ7LR3
ug4bUQ63M9gRbQxA2tEFmJPKLl6B6olfaM9rl1w7/NFI0ocopZJznkQKTiHzqymo
Ajxlrt5HjjHEuS8cCPpSrRXcuQhYtfVPgj5aBxvN2mdVC9YcfkPv0duxjtI4+FMV
EWKo0pOP+ifGlFpktz/0Yp84dvN1w1C0faXejIHvokI1vlMdyFfRW6PCHI33DD/1
M9GhPXBvcEbxi2HO0epfASR6zRprI5Kpbf+dE9A07nGILZ+pFgsb8XnKv/2PJml2
0mO3VfNprM2izc7t/y70nbmKEsJb0ume4PuJlw+sMpE99OwoWfFwq3yKzmdsMyoQ
fMWFcJkN5xZFLhHSuLTU5VUGp/B5pQ4AnW+DxqaYOD3iyQQt+M5yxwn2nWmaFab/
NMA2qHIOP9EYEQWRkpFP/BBfCwntkE7Ljml6ibX0ks4lvyAkRvDQHSy0M+MRq8RW
lkbDfuNuvEHOT3DCF79Lfdf0fCzFbnfV07RvMQqXTgMvA7BzCSnphEJT4sbAnmgU
XP78/K8uzgeavMVNnVx9kN83W6rBPEYtpwQe4wvIDq1D4df9s3vueWbA9US6mXe4
IGQnWFkwPfeVFfzfxIUG88XDs9y4fHygsoJan8Z/Zk6x5Fuv0v7gMp8jBgCgQtgf
B/6s4KzJkhTG5B4KNLgGCpXhKFIqF7QrbgKCGJ3ThEkQCop1U67ShknduNzctUqH
V93E3zLFQg79KK/0IM90AkM5ManjnDoSItbXHmZvFN8YOFuo+h18NCDiVrxxFOEM
rtOAPMFeWW81kAKi719Kw3zmiRm9F4bKQgOK4mRSvobIJ577le0CyZ6TeRuzKrfY
wc+4LHca6vZChZbUj0bTrus7Sb4iCX8EVwtrbMvqSJ6se2PBfcUe0gOtDi2Tik58
03pl+Oy9+HtT09ELYh7iXkH+TIiGOUrISjefmY0DaVc9v3oIlAt6uCM9MSGOhQx8
CCu5INbyNQ/VXX3NWaRn3InJiUAAjZxXApkgNqsToeohceKq0RvEYSECfHEaxKBC
N5eARg8XyMlBOslMPWzxjL9P2sSzLSudzEOWMMIg2k9xITXYUQPv3czPBfTl2jQ0
wWrrsttlybyAU/4zuuyyqxgMEu9DoqC+Ef/TdsP3/wURMyleE7dBWcdkjjwnz9DT
M0XF5/ImfGZBqcFuF5LBRKbhafo1IL6mrMmxjThCHyKBL6ziYE4Eo7yQ0+5dYgwk
k1aJalIt0YpFjvmxLN9WxWcdITtItRlm/UdHpjbDj75j5OFyN5NuAAzQBDYFmQDZ
DmNx0l4exopY6pdz/6/O/nPG4d2cWAobfTsw5bAqQMxvWT9FDPREvEeDowp9EkJh
yWmYJlEFLRCIqOygMH7Pe+DZWmhqopzBzpFO4BOAa81UmAUdzHKeHH7qoBnxkVti
UkZnN2t2IU459T44sMj775VXyq6qUDyp4CwqUtGJYj5Grk4dYpZNOcZpR9xzUW8y
/JF7JMuILutF4Gu8Wz6jnr5idszC0wkN27M7ZXhvN0z+guXGZjM+t6yLzFvh+ivj
YlujHLlswiCOQltA2Pr+UG9KrhOCRY4U777V0Qj7ZKd4h55AWuSO9OcW2Y/nFeq4
Z+uTn6tHSzlWT91FBAtN8VVXZZ8T9SfnFvrsbSTS4hN6FHyrCAjjJjHRpvFUEBBh
qmtIoNRFTiSv+sEu862KtfNK/kK85kSHwSeFLxXh1Hs7ekwuba/eXVlgUvXxxRRk
db9rGs7HaBrik6X+gmS2aYHTWgXu70WWbtK21JD5hdNPh9gfRQ26YZLpFnrrVLoZ
PUPO1ya5JtY8SbIBJkecNgn5AneMtXBdL52BtGwjQ0UxcsBGW9LwmSUloMFs1dv6
yREYOlLp/k3+9eJXf7sXD0PH62OEmVbyEAaTcGwd5Qf3PS0SqaIKoAd+7aWOBnFf
+ZQV8YEIxKVpiXNkeo2fOHYfknkBQ9dcZn/i5BGWjRRLo4gqRszmCracktrZ8A+I
muUVqDVYK/V2gCa6+lwFqAr043oJwcEAH95LMUXA+TqMOeKn+GrDsvqwvEW07RAa
pNt9rMIjWfox7vy7yioXjSKcjU7AMiTsbkkWe1ojpuh9S1zvrhBpx9raQr9p1gSo
ePb+DOCjFFFc284oMr79ijdSmYU6d7MQ7yFa4ZtguKVQcQZ1heCcerP+Fw44zfEk
FAAgkaBpC880MQeIcEKZytGIZrjxeAPW/FboBxPTZZEyuEkSX/+9ipEF/xqkyOP/
4iit0NCn8N42majMtxnac8zUr8RrJY3uIHjtWCjJveVEo1P2YSEI0Uoloh+G6hBR
0o76y3p9mxMHZNUi9q06vVhu9zHMl6oupxdor0A2mqRgnEGbA4sha5t2dmp8XpA2
H0bRMQqnBSXfiQ3s7uc63tY4zx2gnTPppCd/xOd68zPEa2YKrJYQzcV3ASUIalBG
HZkiSQnQIMwSmQ123juwB0iAdrDMOdnQwgYeSBXK1qPkayivmU8a6z727w0cRAra
hWxuyJYJRarlBgKa8s74h86M7tVOfXj/huptf9Uf6gxwc5iM0rgRl6fQkbgijVdL
uKKxRwOf4Yz/q96E+Gu9o7UESFFlFYTnsBSjO0oJ1hEsV0arsD7MrAD1D72REsE7
0vcmRob0GS98joNQusbx3eb1niSXC4LGd0CjeOkl6z3b3VgTzKR9sVAdHpouXm5p
TR1GFzDZaET2p4A9EpUhyyaP3GlWb84SaPyiQF2aOPnW04Dgs4RnQnDeWm8lP1HV
oL+ULjcQ6wSMxR3Lq3dsMSv6aoyME0R8NTn/LUWKRQ1Smw+YVeZv0+BVdRk26v4f
vWRUU1s7BeYqqKsPIyBWYh3vR5FK7FGWJ5GF211xebnz0IJO1cN/LHNuctT37Rt3
qQY9DftQe9YhuODibgNS9ikXdw6pvt40Oi2yP1O6zJscgeP1d+fBny7cda9Y5ObR
/yykFeT+0P4NtPNRlTim6h5xDd27C5+DBAf24SykuJQ+4g/kt4N0wFw/OPbxhk6/
uamnp3sfG8py1zacCn4AX2VPuX/unHF732t6ZvHZgMwakFOHWbhSYZj0pWZYUJ44
hXAtc5KYPYV8pj8ZmiQPZhj3tmvpRnYU5H9Fs/5JR7ZzV9hiHDDxWpp3Z6gfs3Fn
2KJeu72Xdhv3NdDh7aRJGFZgQn4W3RkfUj6vFDkV9AsjegLXURWllW8ewufczyPc
B+8JNi5jzCKOqEahQPniM31T/xIwL2kOFb5zup8utG5dIyR8lrErmDItjZz8Wjm2
8NwhqLwAtm3c4VUawTbLzZR0ywRcpF+SNRReyIEfG6nPCGsX3HgB1zixhOOmXAwN
oJm6K4KwL/ggwB6RM55Dw1qJKWPpGsP/A2qKshMKjY0lDXOFWCwMNCuAI5nw0COz
V84UHqPNBpYaj5u3TbrGcsCO87n2BVCk7dgn82fgEB72YY6MYWrlT4MQsNhgYzB4
4igdvxsZk+VTM1wLcvJXG7sT5APKv4QBuGIJsKDjZoZiShobnYtUnpYqZT8blr6k
jOc8zdb1IHkFKSLE2N9xhOQyKfwzh9gJzscah8f5cv9+lATPl1z5pz1OVARGcTt8
U1xR8rp3FgOwfow0qe/XZbNSeiDMrunuYOOeFyUz/Wy4/gOsU3AJGG005pnczuI+
aJqHn5oRjjg6vYTfIX1adIDarcBgV7pPP5qKA3pFrKt5mHKOkiQ4sQ4LQM4P6wzI
pTOIVeggobjwnAscz/9JKtPnfLZhlqIqC7asraURk2Qcyqr59RDrhWBPtMApR/G1
JBC2DkhMNMtEM7G2wlTbjBVML+qCDlD+5BEGue6Ylp3h291WNwljnxwyqlo8mMiO
hU4dVLUexth60zTVSuBGUdNXK/Et0VvPtUqrkX7EdW28/1jDfOpf3s+WbgkiZwm2
6t3WGHDzrqAKQEReNW+Xyog09bPJD4TxYFpxY3f5nqVPDnprqPWAZCqpY+XI6uO8
QHNgkBzobLQHzzJ+YL5jZetThW2k8ixkMlxMz6Knh0x7iYsgBs63qsqhBMX7upil
iqoqZ2ZkXb8nM7WcR/HTmvY8p9Fjw7NihJUaEzQsDzZFz/jUt9W+RBG52jwGY//S
CPYgCHKnNNrIeqmDIE3GqtHOpnoh80H9O41RlXQG9Wm7xgLWtiFNs3rrgZTShSpa
HMXOFlVTUpT683V1g1k8LTqUW3CpVnvmexeggKO4Zeu/87VbKdX9PRPYJe+EiRlm
UN0U+vhaDhPBdfSwyqX5L6LI7IfGhPw5vHmAO/7ReTLz001HjaM6btkfHP421KPK
ejn4rTMEvhy4TPl45gkZ0FHHyCwOHPo9ZaoYb9pILIyFKXPA75Yo7ygdqeH+UHB4
+jCDHrrUhSIsrA/wUDh7hiUDDnjTwMx8qGvJ9ZDnj1PVJHaibbHsreBJJRsrBPns
1W05M2ux04Dwpt6lyzFS7kLWgeMdsbbuC1ZMw4ApxD4x+si0F/JtGi3oxbSI0BGi
Fsnp6oKlllVtJOuW4nJs3iV/gFD7cWeWfXwxkU67a2o6kYVQT+o9MTwmLIRvwQan
3wJmJ+PkvQnBf8iyVxL5LsZ+tq9fFb85AyyCjcSFXa72g1ncCrH+P1d+bacXTR6m
4eAQNXNz/i2kJOxMmz/na03vJznm4Jg/orl82TBoiO+97eqgG1wDObWiLjYabJoH
`protect end_protected