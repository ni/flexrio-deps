`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3952 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1wB2ShNYedzmkmBWjqK4Mg3
8iDfXbv5M0vDNkp8sRs0MHDxPZFWLbNZbNrPVcQn/RYqC8GpKkaLz+06nJOZtPWi
jr8qK5QNjskGItvTk9Ufdc0w0HIswlMU1SWf2/6NbZ4Q0ZtZjNG0i9kMfn7c3+5b
lea7g/bqYA3xXjsI1jO/aRKX/fm3s49TNxbvR4bD1zRKHnGASYh70OjvH9xJe5vN
FRkijuhyR4NjWeuTu/Nv21Nc7+Jd9LrYHUiyvexH1DnqKbPUyB5d+RrG/ouQaVz8
XBfQKoo6cQ9n1gxL7fB6B1OPnOhxESoPTAIkL2ZfO+DQPp3vKiug6Nj5aymOMQob
gSFzyf30zsUeeoF9JIOGDQT11JayKCFBZYMHCdSIocbR649TWKNKnJ5YXnbHmqmX
iQv9TQrpgpWM8AXp5cOeTndvJiBVwQAn+V/WWGgcVK2HZCxUUQK+noO3zrC9s1sr
LT6QwO4LfWSXLYQj+K11WrKGLdvh9mlZwDZwE3xyYTCGKZte9/lx8/rP892E051X
Hh3UbdpPl6bw2mQh+wT+SX5zie0dv6eG3uqISIVo6sskp/FDuGGcKqcze/Dg6Wdz
La6sh2eZCz/N/y3rUv0ud25SqhuqwcLDKQG2e0/akfIxHLiMsNQkEs8YeAbfBCl0
6xr0JchuyTANOAK7H/j4lZEHk0ghBhFpc7lSELavnEI8h7wxhbggLkJODzlrkzht
X2fu/RFeNXqCZcaMSULvQi7Zfz2dHgjqD1Fc4FaEASlNY+ruPoseYgC6RRi9ccAj
Zts6m8WjInSgcoZohjY3NJS5HiTzu7e+Hn2nh/8xp7SdwK3SjbiRWcxBpn2GJUjt
zSMbMGREKIBlEAYHdgPq3llHPDMakJtTOJL81UKVSDw2kNfVITyZFB0mXTCbHHP8
YmU3934Oh6O+HrT4oKFytyH6H7g6y1LCmXsnxpwLbO54Bje1G0IgIFN6MzMtJcEO
SEvE3VKw32nNAi1lOTiFupaAHcVbv0YILCS0hV9PCw6Jghkhn+QcD1O6KOwZfuw3
Mgvb79U1wOutsam6oPx1lvi97dUmHhg6t/S/MsTeJUi3DxCSV2WO5kPlZGFCehYL
EdOiJwhPCJKFH6VNMISfNkDZgDyMIlqBGiYNyGPTSOpJLEA2cLfwVPtGHKM95kwI
A62ykElwXlksOUMVNDiBqk8WsxSpycSfvHNx8sBqYJAViZ8vJ2vP2iFVJfsjDuUW
GXGckwT6xT3mKroMHkioAF5MH0itgtKAaZ/NmpxoWhuFxDhMlZy4fmWSFpncCxDs
g0leDZpFTPfXjMjFOvhWIVx+omO867NrHaWBJHM0Qj+le2z+WQzLUc7nWDx56dO5
6DyRhf56IHdcX1ImLqZaiiI6DJrN9mFrWi7gS4Na7YzbS29a5icKxasy4D/B/QtD
TmHk/sxNov1aIM8Au/xtUKRoCdAa5RMqt/4b/0XfBk9Lw8/ruRAhy54gaVjozXLW
p8h4F6sGfyv+RcDUFr319xToQUt190n+qfm7dzPWz+WCEO2YTZUOBlC+SmEiuFa1
sv+ArpDPICNzQo0BEPAAHw5uD+sThi+OOswnbSt01GvvlNyiu4+cV1JtEr9sKO3x
F31GvAub37LtGriCRqp1dqFqYFV6G9DjhUHYDOOhis4ilp7xzgdppyOwADFJzXJ3
fFFgVCpiO5uNAvuCBm6aVegK6DXYOrqdzhnViInFt28KMITzsewGikNrbObLI0CT
6b5s21rbhYMhEHro2PeQWBtY/64IIe37HdNuVBGDSIZxHaPBSoWfLiYV3SKG9xdN
YxGVduBjRcMqiQJuPvlDMH7yOLjXestMZRyAf7cjSAqH20md5Ke1D9wU2eqICGka
hQLxJFemWgtBygC7VqvJ/SGm5fyT0RA0FDA+tU4QDxwhz3JljPSoiFjpeJC4n804
vrZyx54wLBVWKb73U9rAU2cHZuKKsz28pH6rohy5JUAJy74qld8+nXWTQSuKLUO0
2g+6aWYRdZHutqd9RlgTlm9epGJqON4rMDIfQGwkCQ1CXkGgsz62TtXv2KavA0f3
kNPDNyaKXe4xPe97UL+FTrO+D4dohvePosrCflOckWPEZ2LJyZzmogj806a8Lr84
0BbTrPNChgAv/Y9XZsGLQt1knv1Nn1BZacYEdwWFSnOp6QVtD5Vk6Y4kKllU+put
GRFHWXrpQZW36Kpb0Z4tY7PXVDqhjaGK0XlkU8cBbl5BZFFHxxvGoPL7ltrAXVU1
eD+mNHXzIXA5rXWvzCBSr03won2edxqtbDBMFHeGW2dHVIuWSwUqEFqg2l7JtbpI
rc/+uddYzv3bAwrF9j3R9ZBtY0ted+Bu19KRmM6D1IhWXZp8yDl0KRLiAiEwn7AX
yW+R9ksWS2D+23f2wP0923x3V/OWttWoaZwZoYg8gocSMYOO20QKME2U8xA2sPDf
begp2SZcLPRMUi3XlC8UdBBmZhXxNkwNmD3h1dez+m2GSABsUT497pP+dlWULqjJ
Jq3cl1B+zB0A7CZ9wSJWJBo1bnh42wbmfakKgNsWW22p7XYRC+YVmfCn1w+nTGgP
T5QuLdlHODQOjjxL8X8zTLe5kEofv9IuFqL2QX1+RNXkDcv2B8f/8hFKDteQBQ2E
eex/QQl9guEX5lzpQ0y6kiSSiLykd2aTsCsssSamVlZNDcmftbM8zIpsMtBLf56Z
Z/EUI8INr05Nxz/kNsX7mcTeIV96GaeXpfnm+4dj7XLZEBKFqrdqU87vdFJvZ9Aj
KQnkK45Zu5RAKlnLFryTBydLaa2Rt9253BvZW2LDyOF8Xecvy+Os//TuEmqYFvZ8
zIuEHAra3gyG2tcQeddRZ9yWCuJy7r52W0KQUXh5EftSnMZbDDfyvolEkKmhXy1a
5x/56A8uaJtYO4pUrYFRoOTFE+l1YCfXaa4jINGKkMaWZXBSXI4qzUrzTKMpPZaE
kfTk0eG/SGmkcCE/lvvjC+wnWZlCOLqIdmv9jG0Vp+Gn0q5u8Ds1ta9bBkhdB3dv
cXcOG1hlGpCWoEuKBzA4gjVqP4OBEez80X6LArRVvPU2Ej8RPpDS+xuZ/9I9xcpJ
p4Wf2pUEUNogk1pyrLYgVP7bKLmCuHGh47oSzyzw/XBX7alUrI8wtV7lnW7osAmL
FzBJguljtIWFa07SLSqlBZgY0GEKJTp58Fz3KqVNI6a6R4yY5BhPvN1mYrdz5gYC
We1WjpT7vOsj4YeGLq8mp5bRzbkYTTHN66SFT8mMl8BTGPRQlMNWm7FIoipIcZTP
Vnq1acaCrSy8yhCa5bLzvX7sYbvPcllTQfVbvMRhZUnsui0VFQaKLcdbUnvRqMKK
LuL44kAu78JVnUG9l5vuMpsxlPZw9VV74OFHZ2ikOc+O0NXBhatjyLLJTYLqZRnd
hFKkDwxhg99m7llsKgzjBWmLxQcQKp7xdjFIwGu1yPl/hKVr5CmBz1f4YPI0ejo5
tWzAAp+e+O0P899bqQEKbLvSdWPb1GwesXoX7a1qu6v1tsSAz3Xsg6+09nhryChd
LcfwajASVPFTmSG3zjnClClpv81UYv78Danzu8oK+8WpOiedG0EnYK61YQ96Oh+Y
zcQMo43lPLWatuLacFsv33LA0gSY8/QPSBmSSAxEGuedy++NO7wP2vsQ+01fQBI2
VVZqcqnRhs5o1M3kBN1waFwDVKEfjaflHX/aHDuix75XJtIwFqqTIc9C2s6MBQ7/
SXNmRvi+/6swx3UioyoHIUsxBS5ZIQqet5A5wJ7Iv6TnyOMrps01qCxpYz6MqwNW
w2AlgbuyuXrJxK7lnwCfnyfYLzj11I05j3vTPjISZO1u4GO4XTP/0wkqvbH+cPnN
ZnUfqBb8lqOwOAvsgsUoK4Zdu8eY1Qak+5JDe6JdeJowVkLneHOI181CUSMZtNeR
pHDU7SHEwv1ye7l051l2r/e28tqiJIpPQV6HaCElztrqyzavzNj5NrdLjL/SMkVG
mZCuvt0p9/AxtIgB4gqTo74g0E+IWHbdXrldwYGbr9RNhV+t3uDizpxcrPDOikmZ
Y1ZFTbwOI7ck5EP+fxq2ceAOgJJDoI4crMnwIlkViuMsY+60PP9V5tMRWiyVOgdi
I8kBZZii6CZM2qF2qT0aG4N5QwoaEp1T0WBUGYCF4dkuEsOMEb5g1aDEyZdhJbQK
NUTMjrKMwsohm2Ony99khosZ4Gx7UK6Uzg2RwTNTkTaaWO7OLl2C5xuGbFF8vJJI
5iN38pBzFuMyPCmxlzTj4aIOdGMIWwUw7RsdZG2DgfX8b2z72fCwWrlaPoh9S+bv
w7U1WnHhet9CjTCJn8OLJqg5gKMfREwgRh9vqNrC2ukMfM5zyv2qTHSNG2aP+JK/
MMOZG9/rUK8Z56X5uK7ROGgiy4MaG4u3LQ9vHdmW+eeR3afQv4pTk7j4OGXdRx62
B831XbZSQiWdnO3KEgjL34YhrHu258UjbDt6Oc0NFcEvfxJxEYi3JC0Jy4fxRkRd
77NLLtLVs5l1YOSS8F/+KiTJ7C4Jy/4EbSqC+U4Jk1wbhRvg0/n6cWLfcWtnrT6D
IhW5jWq1+K+7GwuTL/BsM1WDZ1C9/5etraKirvBbaS6VnJlzmlndIoiXmA34+sru
83V3qQ46ArvytyByqSD/7lFbRT4/mQ1B3pJey+uAH1OjsYZAwzkjPIPWVqmsuGlR
bPKVxtlY+wtIbljldCJgPbMpjh0ffui1dNBdN29RVT2qiBYrLrD/yDhWZvex1014
MVQTzDN5YQ6rhc/YHiNcFjL9orgrD3t65uGyzQqDqBlfzzm9dLpNUMTpV2AvBSx9
1PxnMjgPQxQwTOQajBgs0Ty2E86sF1QqlzT9Qp11KOmocTQbhBeQNcw93bZylwOJ
KHrn9sFDDrZpKQIvtjjbZKiuSBIF8VpYoulkuRl5G669RCkDbV8tJvW5kY2WE5Rz
kBXIGd41phM48LJJaWSaSxOigl8WVDczlevMu7ER8B8dpSq56RkZlGdKuDJxbX3s
KJ1phSKZbb6c66tfPiemTBIMMF1LsZ9jKiZmyL9rzXC7RL80pvq0TBeqjU7cQuV7
EISMdEl1tPxx89+Xlpdo61QHzAHSJ9OnAtOIyjnWjjD9ZPm091gtUlGzMqFSWbvd
96TlBQ0B2Ys/ZiRwC1VNMQ==
`protect end_protected