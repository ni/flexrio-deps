<<<<<<< HEAD:flexrio_deps/PkgLinkStorageRamConfig.vhd
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1712 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
5ebVVNMyfxIGIoeonR7K2xe5BAnQh0GQpMvAifjrCMJgg/6tZ45E6cb1qCBdghoy
4RyfAFfaOJZpgqFv7bdAIOFs6C84ubikROIbkByj6FkJh5j6ZGaBF7v38FnlHCTl
iuidkz03oBePjoUEAMXAyh3XZUlH98C9YJfUgW6K1Fcvis+VQJbwO1VkWIi8viPA
/4YUP0A6qKJgo6WBxddz+PLii3jQshRWexluLSy+y6mHKqNhQKHwO10EdyQvSwkQ
mRW2I7+dHkCezUNAGF7WUTAqU0IO7IqNj+w3ZovOF6+JtXFhVjhB+r+UY6FlS1FB
5DyyqXpWnuIOFoPC8mjasXhsZdrgRr8lJC3lg1su39p97bohQqAel+io4z6PDWtJ
FVVV8sYyPlar7Jy9l2BQVNSCtnjon0EZJ+5UfEU2efTWb7dNPIAEajkrtclBnKa9
T5KWewpro2z2VvvxKrsrcO8mL7aG/30TQhPfYMCAc69nqGoaeyPillLuBRd56GOv
YQqH3sqdGaP1AAI3ELmNNAgAlrfbH6kI9kA1G9ZwLM91hY7iSYkPd35A8hCogEqe
9b1GF7EeiNqJKlIey0DvvFHSW3rIRA4mme9XR69B8k+dtdDKgRUNv/U/S4QnnevF
fLk6YMYxAKxVX7JYXRR2v5Th5DRaCY75EzKO4u62ao+IEeEfeYHfRnf86YInhckc
6VjdTNS5v5VmaTIt+IIWVhsW4/Ndztam8vXZ6uyjzoivHpIw+2jAY9Tbo/ZTM1tg
zAzCjurNpAOHSiiWNbWA20+DNqBSOFLY1eIIDyq2ARrrPpnt9llWxqit5+KzNnpA
OQijCVJpCYKYrepFXOOZA2WYpWCsA459ZH1/YK3KMZiF2jrIogKZcvrH2WaTcy5J
eZvlgtTPAvCdQTcEkbawFLEjCp1eeUTn8RIKLcn/bJeyw/nfW7ALC9A3EN3iNMTf
Ql68Cb5uffHd3Vx7nMPzQd3vMs8tezTReF+HFHXLRdIVEk6aL0DiMTXIEpzxYed8
lAaFgHUMrkd3DDd93AWt5Z9b3/A2oQHmrIipQqdMDSU3uMWlQUBJP2tmG7RGfip0
pOuiPMPJbZ0zMiT3crY7LULll+Xosd6HuAYzKre+91Du97qyovAMeajBXCODoopq
OVWugtXZmuV1hnMjqOM7zZ6/yAENXYvve/om9Ybp2KEh/AhrmqAiYY9jhR+bJJx/
g4jucijzsG5FTsozdgIhcjbCk9te3PrjO+UHmrdpRUj2Zi2zcdb8QS9bzMdBfaqn
5g+KvlbKZsD7pX4w41xRcunBI/APlfgnGrusOnbs8qEU+LUhs62JeFGMwp+DXRUw
7GqFZM5BrnDz5BRPtrrwm3kbL1N8njGrs2y/nAo8t7cPC1Mh/4kNQ6S4PEICmDZk
3KFz9fRvk3qNE0EzM128H/4LRX9FD35bCuQFg5nQY6vbnc2zMCHdLJ+1XT5hFgzx
u/j8eyv3XsjzJhm0PbyeicEn4OEMBi2turzTG5dx6h1QvxRzfZM33pMTa8flwfQ2
N4rMiCwkiR1NjzqiBgDYlF8XRXk5hSkKAtki0K03ooGe2XlIQYVs8QgJpNu0vEGc
MQMmd2k3N8Q0Kld2+lGvTfFyKqrTVQOfalWmvmrNPDKk6DhZX28EnQVXn5/POsLr
/ntTnvdAgqaFBU3MAV1VpLcjuwOtSDU/PaSuZqdnmVU0aTy6KH07aPPVx9bjFSTG
wmifliPSQi4zyJ6+Vi8OUhvcbqRYWIIcpxfeNKrb9HWidyFtTRkXvfaD5rVOWSqx
ATxLMgTS4bAIIOwjYzvMladbVWjDbTR7XLsD8BQ94e+tJitr04vY3UkbZY+bFJgu
vDo9Ir8s1+L5d1LwV+i1klJPbu8Cwi3FiW3Hu8WDcwGT3Y4kkjUO/XKdiRnlqIb/
MJU18v7zu+47KoJPj4QutSDjsTTVaCfYt9UqsJUc7ryv5LLtzAGSGFq7wpF5fQDX
5zep+V6A9hIwhs35lKFO0FBX09mp3nIvuFiTFCMTvbvuV6Eb0phhBNYyP/GYflUm
RYIY5Zayp37cAxU4Vknrk/D7zqQmmMflEoSWRX2acFJ4HktyXskx41IfeBbzuuTy
AxTNQCbFCk3m+GGexi3QtfWVC/lEDJgpSWThSLJpKSU=
=======
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1712 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
C+Ri7jmn92TKTC1Pq3whknqcbygOs7hQVjpx9gEuS1SmKdtndqVQr8U5htAdxYTb
CCyyYtoFTPdccgCmoFpyxQUKIJqIyB8QP0jSOiT+U3eGgwrms9pM0vVs38S2QtiC
fUUEeTXq/WH/W96206Am3KjjBgNR2BWNqF4GAoJ6yoSrwtFrm+RZKZrQfUoGc4YK
NdcV4qXrQ88wUCGwzw8b45sHbKhbkfyQc3zMEieN4qvh2kQbBmZCij9ZEEc5sv4n
w8xl7tJBwzaJnLavTzhFRwWckRSqB69XKNZ2ELI1hzcnHCDPaTsVumZFePbjOV8Q
nJbw4TZJGR9A6tLFeTX2DHAQlgcJK3+fwane/06bTKn81cv1OuHky2BMjmUAYBKR
mJAnEmyg7o6oXAPhj1IMj85o8sqFqrrOutibJeJ7gJ0GryJqQ6uqzbbVjXGfeht4
7layStL7Bhp0by5N0bl9mLPdJDv06xViiA4Hzjo+JhQaaPND4unLgC3OIq1N1fkH
wCmxowO9tDjDBo4OrQ2l1ml+YLdkc8FXl+qpmGEPubi13omCtu921aEhC8rD/JZJ
hDnhbU4PhYsWsRVj02IrEC2aJPUkEmbmWMCR7GWJhhOZNlJRVmJ0YtI+c4H9yCQ6
D8r0+TUN7zLM0Dw+xXEK1M5a7JSnAyEn2dE+uVAiRZGWxkfrhiPKfUzvIhRD8PKT
a7xB3Pr3sg17O1V9Xqji1gdWVqINKNdJWoh/Dy8Egn4iJ0YE0Yzmj/0ZoJNHmhbQ
yVDPdbv8eDhPcTXOg9Yqb9n9GJX8UCCs+qW+ZVg4woqEAe0kkJrAtdTRdmvYsoeR
4998piNiott0dBX0vLCPmfiriEaXmTzK8xOonR4kRlkTPDVdgtQhXnv38hidr8dq
uMc6XOI+xrCGqhyUFV0lq96WVQ4HfPPU+CNmm8wv3Qp4xlHJmkVUlC3/0IsKTOOZ
pFxtqGyWmPiJXYLhtLnl5iqqPaPxqmeuuLDYv6bXpNFu9kGD3N/pdSEe/TgE2Xak
XQyEWC5Wyk9Pn9a4lsQK76Xd9lkFE1MD30J/DAKsY/gUJ8gz2EE7hm/X0hHpD94l
KQ8/sfrVw0S1A8a/w06jaXvqUK7b5JcwvFTJcPnSsXcFiWqh7GjsNAXIzE/bEd6T
Ri9Hhpe+yYmOru4aPoPlJKrtk0zXyJjZTcdamDPMUGaps0xhKU9N0WxwkxbTUwdt
EWlfwrSAPu61SW8GEhTRvXJimvqKud+v6iM5AwqOm+jh+SJ9ruTQh279j0Jigcya
uctW98Fp2qgD6J4NaIbeOSdMsI9qWIvNxQXBzhbAEll4weMlxZv7RuwKCboR/hS9
jfaW8ia9QNcA8xYR/LM1qb/BbN/+rSpNm0Kjc/kGO6EojbcJpt64t5NFbwx9Kx4b
9xiS5+e++g1vuijhAOY3RL6cg+Ck2Ge/eVg1Dc8sItM4sDzu5GeaQn72FNwDA825
pDe5qnJ5w3cKdSfKJqqVcQWeOYEqCZmk3w94/wikEmEZEIpcziEudS2q4DKsEI5X
Wh86AUpf59m+1I62hgRyIEuUaC+P6riiedAVt30YqdMiWvbpTMYVvfxMXGaYUJPL
MgRpr86J3QOR9Bs9udUCueB5RpRoP8E7G4lSN2xMV+XcMEbW2t+IP8r5L7mj5fOJ
pSgt5Bzh3Xulh9amfc3biDrov2b2Eas/F5rKBHQL2pWBzUZ0lTjsQNdd+2LtTks/
CSEGE52DHc+rreWuuy1VuZFnOr2FZ19Ybwllqbfe/iLljipW0TAiWphyhWwbvESd
SJQKVNkEjCaXOEi4SwEg81mtdOp+uLR3XAVkRTToPakAc6D/lE/7WqYX2frqYU9H
Q8sBAhIpRzzMZSPMR6VNwiE74z/XHslKeXBA7Vch9UpJYTWAivNAQhQEfAK5KRBC
Ze/Xe0YTuBCpYSM8L+QFphfQHOjNk2ZwRqxp4i2mZlrwixx9jOjnWQrG1Gp60VDF
ZnctcJQKkggdGPLiUwjUnJYXbF7Q8xEWVMEcChZAmBrcMj2c+zLKdslSFwZ6mz2H
N3XXRbDQ+hyILS9pZLSI/D4N+mJp6Vq4YcDAZvLQVDLyASEZRWTy1yNi2+7yukwg
eaOi7qaivXouHjCGEP7KmToZYlL0Tt+mLe8jhSVt3HE=
>>>>>>> 426889eb8ce467b9c9a9f74dd4af433c5046285c:deps/flexrio_deps/PkgLinkStorageRamConfig.vhd
`protect end_protected