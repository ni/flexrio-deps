`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 22016 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
ZIICkMu+S2rq/yOQyqhpumClsy0g10k4V+OkI+G7LQ/PVGpaW5GPfSiBz4MLbrTS
JTHVanGLtWGvLuR54pOxiB6NgeyQO9xSOky9/p5tJTDK9+i2WAJXxnZF0ZofTeZv
AWi7lblEiCGu0agH3XD/hQssfHBIImU3ZP1TxennRgLF+J0kDT8S5xl9eV+fSTkm
AeWo/JFsJdAm3+DLjbTMLLzKM37PKxSSQ3lGsyJJgN/Vh/p00TdOKg5hDNQPa5rL
YPBx/lPioh98NpIS1Rrd0/3JIl2zP6T8R9AN6xO55kYyki7FjnA971YyjCywh5Xo
JO3PIieX9u6lWkHJb/Ub1jsjP2MsqPmWjTMEikOQdhVmdY87kX55SuxJ8tY38Avx
FhOjLHZuIvJIsnoezg4HMG8W9yHAJLKhEySYw3kog0fqYbOI5AgGnj72kuz8GURx
8y2OOHpIzj6wmVWpoYRGxJTlV/mBRMWWTJjG28ByV5mPxTAGxZGiT5Po19pG6OZq
G48V1rFHRfd0/vaqxCUmV8gCuGlypsBSLE1T3um6Ook7utJScDdcHzk9pHb4lsBw
dS+8YwRrhzzdbb90J9cCNsJfwT4hTt6hN1sqpCvG8jqi1hPDbPNyv4jFFXNOghIp
hPe8qM2xfQ/Ra6hsWiABkl8Fb1epi5+phA3FEx1vcNqcZ3ELsT+tNwqb59BhVFyx
2awkofJZ2ixY4TYwR7cy+1vMtPJPmVNpuY/mUVEGpB9BH36JHvqqFZqg2Hk7oNMX
Cfl4ZYghtkaY1DXA0d6LDsvGmOnLTXmVL5vlq3BUWWv93Lo3al3bJNquNv4LgmRO
Fh0Oizx0MJMEc045Orb+A6rsb32Ioy02xVLawhXvDDs8EgPhvEwxgjiHws3lo7/m
W5T9dEXDUtG/RZdsvuLzNvmxGXSQ+6F8atBUoNK3fYY//Xy9PosbPk0e7BKO1bvT
rIrVSAevzCUOosPe38xMJrATeL8onuEABVewKIDUFE1tMcNfEzfauBjT4ScAU9Wh
TTlddl5iGl7CmWgxIIKZyg4ims1kH2dsq9QKOLsqlvs7d0/9B4EqIE7BZylRBxBV
QBwYWAkBtjxihq48poB+sTst4GjR3lN+139moqdnMHXhdHLmvkS9E0RcMLLnqmM/
1BvDbGxzm8ffrsxuTxs+gDap6rvPGsDImvRvNxyCesRg2c/MyCgXHT3NQphEbMlX
P4k6u/MGlAz+0O6PqDVMO4vby6w/4KsSVzxFkZCrnMbF0OsiSkWoi4ER7KDMomvh
ZpMsYLj4WCxPDrl6kcQW1sKO++zhzkjGNM0uSdGpmQUvPogp5yBOu4YD1jjmpVKK
rhG2GDNmEjL+IMrKYau1ZG2mIenVSijEHoRTiRsOv/3vBb72y/F3JoyA0ctOOLbs
iHVKKlMB60LFYuNFThUNfN2JKDKsmGZNKEZUZUsexLzcNuio8e92w86YQ/64xvkJ
EHtaq4a0B4VJFSBauYQn93h2V3OI2ilCg06pTOZH9VjI5g/5ZyHTYv8mZx6qhWwd
UAwHL/qgajCIngLXKX4hIzGlwRYR8ieOJtZkc0qIBTzNgGl9ukgEpkNqyWBPDlWl
BuplTyYswaSnqWdV6NtKymgvRTxK3wfNIhjeNm9zVn8oyjcdu2ARPz5soAo44/XF
Er4CzZkBqIEJPLjMuK3PU2mUlM4y3RT0TBzGAXJHncJ9+tMWN6Usm2a9eXBGSslt
WHYjNjgWtwKNwVXMFjL/X0ybbtk92yAzseGNIBSsh/0Pu+u04pJ9HLQARerQH/Ut
jV65rm8F/1Uc7aYIJZT10fN9npcyyHMjM5TA90+YzR5vQ+ElKL6SDATVvPqPUpLC
HHwBET9SazBtRB/HV3WhCqbT6tI6FZSL9bzOhOhZ1Q8xSaFT/MNWxTy2QjdOryZW
rUjdvxqOKucNITuwxT693Jg98kr61qKmVhno7P/AM6ikal1EriPLw5R039v3zwUi
+S6f9YuApjrnejjNRSjPpze5WhhIh6vA/gQe94zQ/w519XgqcMDMqx38wUcBRd2Z
VbZxk0uqAquF0ywnEJkKFa2ptdttcu7SIH6z0OG7gYjwIIHKTGXuASZXhnHA+MfZ
jOZN/+/TCjuPbBQqYTHlM1NVx4kkR+kV3OzrIfm5rSfnywWftabg+d560OMfEDLM
OoTVjb2a5kkAHDU+mVBXat3RMtE/g4H/7mGsiS2nvYDVgzZi91VNpIpR+xJYKvJ5
5Ad46Md2GBDsvQpa4mRSR4e+fmFC1WpJ/lNfNhiVDfl1c9GFWDDf9zTTUkeynDyJ
SKYU9JiaT+UnvsEHrlj6zwr+FhveFMbjlkoAOkEB+2aAmqXKxfQ1edYr7rEYXLwr
in6EqW/qUR/tWgwLlUxJaua0wfKrabMtfqaE9xU6FA34+xGKxCrh5OBXbo9PsYB4
muZOTQiHGZb97g0Xf31o6TCqUyacfWOe+IgmLVegFbHS7n+3b4g7RdmU2ys0nz2x
2+QERFw8ntUO8HCaSWs9sWXqVjbS0eaM7z8xMG3LaTgTidXmdR775xLgTvp2OWVQ
nJyGWSkH7KwS2zBDphbZI0h/WokStRJjs5+K4JM7aSvk0zaoBbmcTjOgOCWyJily
EeI3gbMKEQFB4ZFggKhahPlQ6pfN+jz85C2pX1cYIfK9KOa4xUGspKz4QDsaUZmQ
dZPerl7sh9mcraPAJhTs8VW85DNNBnpaB5hsJi4BtJnmrlFKClg5MrN+OJK1HkQn
MtQvClGXNLdoYwSBgw7RsuK4KI3f9oEB8zYWG8rZ9hqzuceAqNzYy9uxTy2GyoJ+
s5bDURbStCaxTorbPBrJs+NCw0i7ucJafftnbDsG89jAGk9p3fyGchnm5rnPhAgN
d1hKrJMO6V+OjoheXfKUq5JEQmfniC6SwbpdFvrWiyVcLDijxEzxADiqo33sGlda
ONJHIwBVuBZdSiwA9IyNGjOZ4P2jJNPG6P6nvRbVc9Dxh+YEuaIACtVwp3Qu1cNI
6QF+Plpx5yDARUGQ9tlY8gbbMTl9Kwq5BoGKWMJ38XhHXz2D8ouPQZXx0QiML3PE
NLRNhlIkVgwD9Mj6+sYzhthG0iCIkx5OtGnLNcTkLQ7dwpxoS7duPOH6+zbbj4x0
UefX+Dc7l0mgrJOh+InBZW5TJHtcTs39s/wiENYXET6m+nc2V68wNjG3gEfFrs4a
3QJomPBpwJOt72/kt3atbceonm2KWQAbZ+y+PZaYfchPqalSuEEg0GdJoetuZDLs
F3aRhiFZ7IffA8RLIBOrpdOH9MAwFtPnhy0j6kF1RwrBFYO6qiHySV83FUTRNg7X
iu0in4MdZXJhnmqsOlOlR3E+2vNtu2Pc+iTZBZ6Cfoka9n8334f8XSUa0sJATYcW
qD+LvwTe2GKbX+ylkjutpXpCXZM7oRZ9p1L2YKxHUBZpuVkoiDC2GgkIswCHCtmT
KQfATAc7MClxqdaTAqqcXgnLqOAjEMHFHCB8cBGY/JeB3n2pwE+uCL9/0hAK6tVQ
pRKzByCJtCzCK0KKc3QDGT6FDBPlqgqwymnRNUpNsRsOJW7qdkRmVwaBGr++bloH
9Jb4B5ZIBDBmruV4AlOy0FUExFCNPr+EW7zTbybsjWM2u2ZVny7VjMqsjkybNGWn
d54blCqSkZU2zcKgnuLy+s738ZZYZYyoGRPNGkRyz8Lg7vAVh5m835fsNKBARYec
9a6DzXha8qb7RD+f5ERCBk5+eSt+ZvQncN7/z45859brw+Eh2saZtj2IXEI1Ye1x
4vDatNH6CXE2YKbGYEV8qpxtPP4x2sGyQlLnOcyuyMq+SfQrKO8EmwQyADhQYiD7
sEgaDH9Ypbn+wvya3g8ovHtt2qJQJJhcw0zW3oqS6ecF6KQx+ZWDCPNBUEhbvW40
jo9OZLEkDJdE4tN1VLOrNC/bLf5iMBz4KcJhKIEtLCluOdaxZxsSTptL9doG3zGr
tSX5vJB3jOhjHrZQbpgbX+ozRLP56/S8PNb0MwF+r7sMKiEsOF5+QDX2rnBZxlmR
XejROb95HbQlr5fT5ukK1I3HMBNdyRGuUwlIe8Hx7vZRQOWbsj0IiWKaQ1RdY0PP
80pbXG2s+pMlbAdwWchkHYO4X8JzpcNaL5iEX4d0cCkkDPlJgZsph0/R1xqpA0hu
MATwH5UfJcfYxy4Zb50KTe1kayNijzkiJ3kBURNtF+xmLg4JafGxDINLR2Pw4Ktt
tWaF1EURuntCsf/s5lnnuzZyODdgGJRN0Oncm9zgQNRQBP83iR7XCZpwjmU9tLJn
LxYp2f9Y6KMazS6g+3JbsuTNUmJj26db70FquZ/ygGbZW5Vfj+d84zsYVNzXF3a3
7Lvn5w83WkHHnmxkd+vZb5EHDK6kacrfM7zBsJmOJ1I7kOBmWInUwAQVx5B6yEGs
3/A663LvAZPEvXvMRNQ5NGd87ox/DwA2U7vhy+UCUXdgrgHs8RQl3Su0u2LLf+kA
w4iCXGK5ac202FlSjnUuILY/v3LGX3UVcLuY9RMuKjP31sAA2etFVhAIV3YHyShp
MFP3btQZXGsVRqLZN7JvQTqqJbbdfR+sEgMl9Qh3jed2TqcJMueaVCulKmn1CI64
K925+gsSB7mfVly30OcCJb0BQCA/zfJuDepm4IXuDUDLYHQlECtcEzj5tMvijZEk
Ks490Hb0iJv16Ou0gN+UvDIJb5uKjD2CI08IWkwb7PwaSu79xfSJjdez8snVHkMd
syD6l+Klds6By7j+m1TQx9tlVmcQOtXl2xQnmQhMR1W6NMtllmKMX0ezJ/LVr0cB
zZwXqrrpHpcXwVQ52/ogX3CBVC98bcu4L9V11G0PayBFMz4sWUVzeg6VK3u1HcrS
miIwmUfOPkLyCBVQfJI2rC2WJYRVKlIqUazy9ntZ7KFzsxnszWPdUkdMoW8qmsQR
9cIZYed88IWU4IDSYFQWiG2j+19QiHZNc0wRmOJqHr6VXkcNI0SH1s+jqqowQVbu
f/mYMrsV9bnomV7f0dApDypDab5sVl7cOcPrNlvWCbqPZZzk7VH/yEhV1qcNIJY+
zokpxKK4K0Df+XqeOS5t2Q0kf6tiwK0tyNfWxWd+O6bFfiIs6xBn1nd7KGllnIWJ
cdtFQplPwiSXV+92tkqDggT9q1n3TV/xri449A6K74xEnklqKSNya5VJbpxYTEec
+xxKPsYWGEHlZgDSv+wOaF9IqcItiv64fctd3cQK1w8M6BPmhGuZ3Zvbn/LfeXqm
JqKQDeGXjIQqt64wpULm8p7Yw4fiX9hg+5FubX2bgDZu+7UvYZ5QEUIpqkmH4SIn
nU8pg/zEQO62uXK02z1NhynPajq74FVWV2iQKkBqakSvy7Yn9JmdQIAti/AGz4Ai
zElSx9kg2AfNmv9peGzmKfg6+QGfX2syIXTzWiS8rMyUG3ewOCsPYj65XjcvGGfy
HloMcdMJuqjLIHDHZYBP/zol8wMlyLuMJD/3Q0Z2dBIItBxSyC1MF7zq2xvbWZI+
9tOQXSy2IGx0j+8cKhk9SbO0oD9ntaZ+79YwZhR/TUNTrXRhVdeV0NdhYNCycYnY
Y3PsLQ1KEAjNySC9872nSgmZt72OycOevdKHEBdP/9xo6BgvEztDE5VrIgKLfCdh
rNfZrHr7+wxEGoTJySxk+Hu6rpqq+p+uXTaT8/fFOq61yXqhWLsnvLuKnZ8qamAh
rRs26Nu4wvnETp7qMB9XAxhxRjOQ6eS4zuaTjUGH890WKOn7GMi6XfL+NRKmjYIS
+GLFdGfo1icboyg3++HZwcKZQfXCzOI8Xw12KdHYXW0t+DtxAsJEex8KWreivhus
lHzfr6R7R40UeN3ZbnnFo+SrXKkCt3y4uqilXtj9Ws0SuQZxpPgj220y8DoZkC23
FK6FqxiqnS93CXwcUkViM+rlfBe3Y2GDF/3axeYx9Y+u3Fa83vllYA2Nz81TJNjj
xtB88bnIwE0EokSF1XGCR9f3c9fkajANG9waMGJCHMsyk7tt0i9SvWGVJFWnrBiK
sN3FAVBAPagDkcHM2yNAgkhLgtYBMSeonl7uwfJR7Pb3YUuWn9Wwqh/Jcp6Flk3C
2nUcZbQoW/Y/2J56DK5tK0SHQ+r2kOD2XWjz5MeRzLt0BLiMu+rKJnciHo+rN9ay
9iEqmBrAHqM3rAtyANWvme3xmELtnPv/b6qObrhaCD+Md5D4Xau/3RQPsVQJxO7t
HuuogPMOhPO+rgSDviY+6xrBvNkvvIulqGADEKtRN5W9WmNRTNnk2B3BwUxlUgT9
17isgrYx/VS509cEe7IbmA4keotTs2yov8WhvCLahIfpab7gVPq6kogo0JSEzEJK
Wk4nS+VeVyTMTC5peRovZAa3zc12qlCoJHWQyWBVPQ6F/Zs0CHmaa5EZEvpHOvsb
cphPnf/XDwua7A8v3uycWSWdWyBCvwKS+iHV+FldVpfhO+8De9CEhA69COFK1JG5
jLP51JoKnO19Jg9mnHNWh6g/oTShq6VEmPQEXY3oa/I6z/BqVKgWUKLqY2p8fT/I
ZgTpm1meAmOFafL+qW3szNql8odP3o7/tho/H+ITuddk7WJ3QhPv1pXZ2AIR3AjN
EhBn8B+y7DLAB9rK7fyJymtxaEixeYKYnEmYxT9F/S4tDTdu6QwhAI+9wC0eNbUm
98q5PGL9izJf0PV4z7/hFjlfuglPLgTJF5mQcct7cZZ8QPklYKYB1YveagCGd4Ae
JsoyKAauQU6q/7XI0JYYqpg6aDXi9k3It0b7fazCYiSbtT/6cDynOBgfNMxBYgam
T8Chao3YPdBNGyfHSTxE2bzgKpW1yFJbRFqWYp74BhNptP7T4ChMHcOPXs8iXT/i
qiVljK54s0tT2E52KVuCg91ipd6r+O0G6O3iBEeN6kSwAKSzKwQf6Z0KAx1d+kPS
DDpWcKJg5f1cLjKzzvrfOA/nFPrU+8ziXjDcJkvsTIQ2+SmzvcMzpxa3q4whCByW
hDhOG09O4fMb7etQ4J7FXimXaq8DCkvzVYdHGshsgubV0N3RZKABB3lIhqPpEgAC
OqgDoXC6xgqHvFZ1FUDIEnEpz63mlNjAsn70e+PS9iy5sbQX7s5tJhMsdXONdIvm
vf0v93u7f/tAGFaEUOhypGb3LB2r4FUgYK+mMW8cNl2kwQs9sPj9fxFUAofi3M+3
CIOx94lEVRr7oD/ehYjWv4TpAVUqw9KtaoJfq8JwjH0oa2AmoEwVyDGMwFCDDjDe
+2J3LRA6vWbnIfuEdzoI129CtnWtMj6W0Y/s3INs1NIvEmHom9eaumo1Wzx08MF8
mojSwHBCkmKFmcmG2mVxkJi66TdkoKOC7UJtcyKBP/DEq/rYi4xvVjApGBMIlHdl
+md9MLzkeDupOCyR6cj9zPLMmieiiT2KE+RjMw7a55KFTiM3UNzuja9IRvNXJb2L
QErZemdt6VkM7xxHIdzp7bKKuD8dLhqjiUL7zTRvIZ/v10Y+LFfS1niJ/uwyyEHD
0mIyX/nJ+ZqsGu70gZw0XjDEEGgY59gUKbYMT4IpAu7oQhRdplBnD/8xI16XBfhE
5YuxAFA5vzY/lVbE8N15hpSnwdBPAOspakmCyjfanE/gfOuD1XZHQNVW2kK3qjqa
kWc/85LibTaNAp3zEQnb57MvmKwSv7Es0ET+g39oB7lND1CV+Tfoc0Cwe5/ERf4B
0BHdylybRf4yynKYf1ubFeAj71GFKaFPTcMCmZk9uxYei9UYJ4zCPlAeaxGlUPLs
AYcBFp054ho6uEPZL75D1j8r+xsPpJ6OYFC4BxLqBWluVs5VBN9Yq5WigGLfroqN
X954fDe79RePJZePxbQIldhpQKH0Hhg/6EqJgwsxHpV+OnEcWXikSStLVzNrJore
WRtAfGh4cTk+/dmY+ixGJxsimHFdRoH7ezssBHruZ//rdyHb5yZXybYjV64UpInc
dv0PKbm8yF/2Pod+hrOsAkgrDCNvTRIX4ts0ZPAA53jIzGYve+64ZisEhZygjolG
FSznfoCtvlngQcVXv1olPnTSdADd2PXMn8DyZUAVEoOtt2HkURlBzKT3oKMJSsv8
8A+spKi+0y+9IZZeEemMi/JF8OnNIcBv0YT9gSFvusRTikp/H6RD4PnIhjDL655D
rWC8nV/sEa6TEqyFUYo2Pjm1gJXeObzDGC7P+Xn3SuSJsmlbH+5Wz5zebVI9xlc/
0FnxIPex6JqtpiaVO4K7gJUoU7vb9pUQZDc0xjZGJIuUCBYoeH/E0Izjpwvgd+sz
jNU9fJ0qA5nNciGW/mWlTg/tA9H+wCatqkcGZtdQLjnPEm2g+0ekWgWDwknuTBeI
7DCyatZvLf//Xe4WHtlQosmQrgMNobKEAZh7jM00eb8nQmyomDvCzPmKFncgCBCM
3iNrhZXNfo2C7csjILCw7Gr7Q+brBD7VlkK0zVcPUcHLMljCLDRRo7Lju7pvnVvy
rpJo3Y4KOahXoIR24AJObte0kCgmimgHG3VBp/SDGwNYrsjDHZsFTrbX4TLlOXw5
+zlIEhe/8h6kLxnMFQ4l9EWR4ra2uFhwFlK+xTfEciL1NvItwuzNZtJcfIFSw3iO
5v+xQfs7kU7CvhWs2UNJ+dfT/IGAt5atNtEXAjcHl54kX55FJi0gnqmC66S/7RWE
Z0nmRDHeBJ0/sGOQrFMKM4vPHArfXBRwSsptyJ09A+JSYEmbhb3PXsWoCQdt86uq
f1uaAmrAB/WTESBzSNPdKccv3E/JyTSin118YZsLSOAJsaNMJ/bAaYIf3bsHVM4p
ZZg/NmHwyZXRHhKBjrU+0HMjk1VBn7LGv5eHAWgAdJYVSQ0+ZEiu5GIkLMegt1P9
n0mrn7Gf/+wjJO6p82X6ma+mlxm3JcVSso0fX+GbouQ9Go8PXG99kVeMTDsHcG9B
YxMs7mjPidX7hFPkzDnXdFKUtkKktxExjA/4CObyoFCqpDmKzWUXCNY1PpmQIZ4f
SHqgljGmvBaCwOpT+eQ2sccDUk5yyXBT0vSXzsnzzJwLMN3q8Ycqw+NuoWFmL5/u
zi2HCygpnYwD/6+SgbCGNJY3EViJcaEy8E+dzVqeTJSh/PWCk3KB2NO2tVNkghBs
tFTQ3VWCrqtE09y0AwJEgvlOHzQ1BbmGXws29UESRGtT4Z3WSOdtkPJ7kweVWWF7
vibmjPFYxxmx63K6ThIQN15Vcv68+ERfQt3IArCWNT6cKLlq/VQ+GMflHPW3s9wu
J+tCSx+vMGYop8aEaswIt3zFDIfKhBJcaNJvgXMEQD13eoZFIF7HEl9kWg0I5pKy
8ixlFGZv50Ko3DiLioI3LKth2qT94/In/fY5hMfo0Fp3t4g++OqviE+pbok9Hcob
aK3R6QHYUGWdnzfLDHNuIBPKe/Rt6pn7lZhJcGMSo1UHIh4H88Dm9nzDIr2mW3Pu
WpiKZSRnsLoUou66PdiMJl6owbRasYz4DDsMrbKSuW6Ou71tbwADqPs9xMkBovef
J0uyL/tIagXupZgCT461i2SdXjwAu0vZOUyiASejq3aFYrw0XPnZ58lEgvut+Ero
fG+E5RvcmTKUyQ1jj6sBFQEPYGj01O/sON+337LwgO01YI6KwDFP3DHCfKZb/DuV
Agfi/cudVKJOAembLwMlpHj6MSiohFtyRu61Y3uupNKcpO1vgpPVsLttAXftCBmu
cNPxg28LAhS3g5oBD8GlNUiy3HkqO83WrRnAvxoOUaCVgjQadj02+clbUGPjnzPx
43TBcxSrnusm7CcypAiRShLKgMiyM8OdCT5g/4Vj46LUJLEcoEwGV0kFiakNDQ9/
XXp13viNTBzaPn7fWRt3IhtGBcORTz+OhCYGlVJOGMIWEFFmRdLoRSINLCDL3BIG
K6LfTcsUrR1d2XHH6X3V66o43/aqEHW0uQPzM+kvwXGBhNpssbmTPXDaLTlBA+HV
iy/IEDFJwaBnLLGR7o87erGeKs1kCAcBobl47TKhl3Qoe3rwSHPcsoUiRV1nhYhC
D3NoVRmBBLAWurBjM+u0OEFzIwhvryI9TWjyPzqxJTJ3fK4xZgF4ruEap3i+TmrK
vC/O/hDsDyUaVz77qe53pHQkOL6g+XZWSDU11u6Bh1XGzoY85osB87NJVL73mcpc
/eiFVv/RBnJRwIjQZBqRfWtDjhBeQ3rmwLK8ZAFzD+h9pw8gc3xRtHzQE05lfYjF
Pxc20O05i6DMHCcfPH9n8wu4TjegFXYpcTNvvYlCBR0f3Jqp6sdS/w50LX71NvwM
yf63cagkrVuwBPwCLltbBlzHolE8b3FDmWbI+w/V8rFbaPDSRFA+gKWeA52q43hz
QYxuqVGTOY26b+/PtJyUNBpGjVtQHa3vUej0OE4fKSNYU3URhvq6GDOQbDBZLhj9
Vo1qB9nk7FJ/RTRY329FJ4k7/NxZes27GlBpDAmskCzkyeB8zIm7oF7n9IbFrDOe
wbBlURWCx/bsg6iMwL/zdZQasD46r/j58krwemNrdJ7DC6j2Vvt8GFCEEZ+ui18K
bW+k3ACrNEu6RqJ3nSb8RTPYKKPzs3pZd1oLL1E2zqX5K7HycELwO17+Ndn3Qp37
ArpTSoXglOucse4S0dyrPwjPhD6rL6rBiGKQ+CaMpdBPWUIur4HMCAu6WcJgZHoH
ElD0x7Q81B5N7Eo+F/u7W7zBYa4Ahhb94rZlFG+llj/2poZBZQALO9ymPt4KsxxA
wkGcq9E/wZCv8zpup2BUs4DhNOikdhHpota4VSfJ+K+IfAneHRDqGRGLeQWh6FZN
FI/ePTkQrip9TaAXNunrcRL/AQ/OzcWdkbQTLIWo7ccZrXepyP43JLUfnRMHNdwU
yuvjXE22bQPIQ6BRPRkhzgOUC/AdSLcAK+IZeDPnIuhqulBar3haTVvnNSV6AB7+
nsWidSJD+gdkAUaGeCrDWykZzk0idrFCNOb3HNbtp1+vRJ740Wsrmk0H27RrVRy0
2so/d33K+0xPM+elNJ0DjiurDQjhuvFZRa+PZRICIr8y0LV8+XkZYclYvLdiIcsd
rtQtoyY3ygoJcW6fejerX00DgIa/qGvU5XWcwRc1PbAmryl3rQenTefT9GQxnJBj
0CAT1ckcXggQ32ePP2oawaVrmcuXB8WyBKsfcFTX2gLIOzp27NPD6X+lr2L1BidT
+QrDZP/sv7Cuc3SFVpPFxH7Vtw+hJtzVHNGEq2Y3ErzfSoijDyAKfW8BpJ/2qcSB
Pb3qJDc06tIWZoQVWj2Tq21GaVpslG1dVATju2CbDfXJHnhLy9qT9uZ+CCDmI3lH
4FNRPfu8JUh9XCsohY9YCIlU20r+amezC4anT9y8rQzVqMPVgndaeUn5F0cGnt4y
Z+pw8gbjQOvvgf9tWeGB65tCcMsFAZIS5jNUTXGahuI12HJFYFoYUYMIQHHCX06h
k3wJwuFGT+Fm+Zh1mQ0CMSolRAwN6iZu/KGJyajl3qZQp7L8+/JULpoq2Eo2sW5e
xTlXxHg1jxgeRA7LvxEod6KDq9WvNHH/dDuqHoM1PoXg59njcDMB6uKUaLRqdBYC
NoCEZfO7z4g0CTCn5dnZew5FSP7lHJz05V5xkJu/y3Q5z+vmKt48njGlLD4XG7sR
8r0wfk3IWFzuhm2pwy446DQpZNwVUeKkB0MPQmatSWj/31yyMgHrUp/zRmw3m7WW
00UwuJf1ARtvmZ5bQStxlTyWkyjSzlse9WsmNnOgoJXqYb/JaZgSMQ6NiOAeonke
ZCWiBWmcMRhoV2uWmBRnKgIzEdfwAHToos7yt46dJmRP37LllMqqbW2VQCnDMCVm
BsqGNKgmhtfLMS4FknDwlKor1PtLP4DERCvmnOYQ569NPmIKmhY3lZLalsWXi+t1
hcsl5sbFDtiGX3NmEIyvfXd/gTX0HDT/74vsy+naWKdKC9kgb0FOkmN7b8jjWUTz
ZK7v5qWwXMS9yjAjcUc5G+LGbaXmwos8G3hK/JBmmVsOAdRY+F8bCGeSwRkLGyKc
CCTIu1YAwRzmrKYg0yIu+vvr8MmM/uGEgYfu5anZWiOpLuVYZ3CvGTWX6TksYT4l
qlfMGH3tolSfk7HiTqfm9BthCz1FvMX/bC010vwHUqorGj2UlkkdHOJo9L5y7iz/
rXnOL/ZoIbZ8uP0xV9ImHLLr5W8+Eap0ihkTh2wfdBT40wOk02tp37VTqAVXVChu
pvXUqe0wK/NAhDU+OHrdw9A0Iv7RlOrvJd2uGKpfimUAmysZj97jP7X/RyZo/5In
ftUiwnFqrfoIuwa0HLelT+uefNKMpzXW8BdG1OrznqLzA4ra9Bve1jkbwpoifkYk
bCGSAzSqUCn0L+/nD5pjb/mtKudWX6QO0+8wHO6whUnLIDf6XAKGy84ftUSb+ynA
S4HjyysQhsPg2nlmgqE5T5rt5k4TbwxQKhPnJlToh3Z7+rePT/7gPh24kqcPdmlq
hPMX4CziCjOkUzQ/X8HICVy84S3vAOsX6uu+zeHha9GQt/Fj2apa93p6a2clbwOb
RQY/GQs0P7wJ3pH6ifbca0lsVa64RRMPJTgBCiCyGBB8HOfDlAADqhS+d2dii6LQ
xry7hzJ8+7+zFPvJyaj8W4VHjse4XbxkAP+1PjKE0yUP1SiAKDWYz5i9P3ui5mzs
T7HzQSbzNXsOy2erWjwBVn8INuwi0QsyQpCVFV/7ChMWm0X7bQcAuVjbaLatzzOK
xb+lsgdTU3fPjripp9OyzceZHFfwYRJt1bdBNLESXHS9+GdqqTQ8e0DPhkmyAWuA
But+AzdKLPIUCxuh8TmQQ3fFcdVArh+W4v3j48615BbQ2OktcQnUidKA7rwhdyki
KYHTe9nBNIXXYaisTPRtvMNvbtLg309TZ/x1yQx06ytqXnauF4Oy6KN5ntmojRf/
gQx4btXC3gbe1p3nnakSHwdpXboNR+dGAwhRm1KZXNI89QUBAZ+XFxVnmA5217/S
lUWTcmCXLUcVadShKEUP8U8PTEWFDZWwWB6Rux6mWQScW7YCzbK60hP72vWbpbGU
oLX9oMr1HYQ+47iA18KvUBBug0MV8okotLLkMNBA/qR4UCT6VGW9fDAOxGuXpbRg
+HwgaooWg766EVu2Im8HeWe8/1EtCtEYOZmGVEFYKT1Unj/HgfwJ8+CA+R5s6U/U
Pbo1ZxGqLtKGssW9qjwnrx6QoIYzhxs0/42a0FgtgVFb8Q96Y7NZP5OQDYTH8Mj6
CVvJsLY/UsaZotQ2dl2gOTtjlq7dHp0oO6JHl/yNfU7pKHTb48OhmEfTtOqNk3Wq
5YxvGirSYhlb2Mg3lCj2JpPfEbqs4ZdLHhgU3FQm/Urp8XenGJmHDU0oSD22Zdbi
PJaANtV/6s4ChadHP5jh2qjhdlz/v5leGospYLXpzwWMqHmAk0VggAlrI1bAn1kP
C8BHikY1G9ycRTtWdoH6WhkH868qmbT+LMgi9tB3rsrDN50azK4tVXLO52/gQTQu
fHiCt2aOHxvMVZoMElWFqJEh6rXT3YjSyvfe4W35B001TPSm2XHZd1OYzY07+7d0
BMkx0XCtw0EhSocaQFOMTzBNrFzzKzp4tKYfTkvA5oma/+270OMuoRPnkpCQef4Q
m0J4XnCVez5ucI/QiETbXmQHDPuf9feY3nBx+GhWSILqQR2bX0NgO8cAxcsigEfs
gMrx+mFPnpdcKtb8AtHAPUC1JRIfXaAILkaR+FxzIAcBiPz1YNusP1ef/j0M/PA4
WbRJqA56CWR/xM/9Hnerxx2lLlpluu85qtl/B2VUDhBQAENfPt3fCB9zCc+nyW5T
Aje/l99DqnaQucfljw46tqVH3UkOMt2HT3WbAS7D2peEmhZnKEUaoLZstnphhohY
lLepVpTxZfXiAsuw6D5SvdaYedEQlQMvwASPTu75Ew9yODGYk+nNmTka54nwHF3V
dWzsDw37keYvU2rf2/WHjpK+BtW5w3MOg2GEknVI42jeTgsgAx1PAoHcbC9wTk39
jsYkZsXaagD8hW8mSzQY+omjld/EVqLttrYgNKnH9VLeJMKLMycobfcydAVKcjvL
mPqV4VYuap8rlQDI6XPPUBt5zhkp5tW94YyAvdbtuh+yK1gHny2MJqdFstw5u2K0
YsS29LnE8epnmvEfWfuUUudbRCj131WCB9TfZL5P7hhyo0Q0ug3nlWiCnnZM2+XH
z8gnVSh2BzViNTYF8qEUPUK/GYMWAcXUOtbU3NwU3QdAGWwg/ZAKiD/xQD8QOsvK
fdudoaOzYGbqVoAVMcXBlJztLUGvib+naZlY7QirBSoO/Ys13G9kqRyZ1gVZc3Lf
RIE0quBXy8qBaeMJZLG6IUwWk02QVEWj/yylp5wCBKEGTMXMYCKXmR9I/1REN5MH
LJlGZmzJXOrwQvGsqNJeDTsKoBmS02QNdtBdz46rnGxI0qi0A+V81DOoKbhJLmSI
R3jAo+n44rhUWdZNV0iTDveaJTintA7ae/oYlmlrME8LluIOTOq6fpI4Prwda1X4
9N7ji906E3B6k7FBVtoIkiCn05LxqgPg2SlxiT0XwrcsGDZ7dPjj75bqvdiY47o/
Yqc15F3ZTa4ofp+fQe7FGMroOVgoMNolFzr+v8i91cgYU7p9ysaWNn8/acKXAGKR
0cqznuxnD6a/CrpPXP0yBdq0q8oyWunK3DrLateF8IzP1OVeujsq4HMbxKUwznJR
PrR4rXkkMZ4S4vjVVi8T0PzwkG0cVto91LGJLfHh3BTdiy5VSe6/qitdkDtScf92
LfA6CEcGdPnGpWQmKlZbGkQjjEoA41xj5WEcTlC03bTK1gHgPZdJ8ztzPZD18rdb
d8L/zwR9fnjVbWT/CiCcIRvKbhyfttzVw9Z24xchMNptI1Qx9ouZ07K/6PqIxaDY
joTT1PHXSAfmo3McwOe7qH0tPqJu5p7E/6BzxirIogIXRiL8P4+UwDzh3wabms3j
fLTHM78zdVa+JQONR/UiQvaMh366PGgtma6YzghC7iHwQ1GPDFcTxMFqDF++Q7e7
kz/4nn4dwVj/szdz6V4Lu9rlxoIj5ohuXYqwC9YkFYW/UVYU6lGQstJJqcsNwPgs
lBrsxMshzCUNBWDRLLGtu9XJ6OJlFW8ED682CboNFdJwZcIi+OZLypxxqfb+lElk
IXQhtq1DkaN6dYaPbz1V/bkLwXykX8FuUVgShOYVIHzMc9PvZFSe+QnoKgRJHUlM
f0k1Y/rlbxsV+PgMW/vtxBYzI+ufyIZt04Y3GB2shUdqzCxtN+V2wWEp8M6rDdXN
NZoGaTdrzygGiGWqI3Qa/rXCNBkU4SILmyuTGS5LabCOQCKaeHIVUL9Jpw3b4eoM
LLNK1WKfEGpxpOyC/NZnp+cPp9VZzdHx5TeUzT3IWgzOcrP0NHDziyKN1cLDYSJQ
NqxbgRDZGpsqqOQzogelMNrT4h9xGCQ5ZyrlSAv+Pw8eXEsEbLJrIify6gAWcT3u
jF00AcB7e7/P2IDAe48/bvm/GyFTgSrEkn2Jc5FJookvBMBwjM/OlGaEJxbn6KFl
KjoyCHTsyDAqkOjhiyKFCoHbA3BaNLnzwQVEN8lbpyqaqqV9k+VYCM8ocsHW2bUg
LVSfm7GVnGfRjZqi29n8WWcUspkv5MKTlK/UfgGqpGAlv0UIBLJ5Ki5Wm9bEQG30
Q0RmGyn+CRPAhQJcigxB7qX9kKXipEp0thBOgKHWkfHWpuyvszvzBp8I7xkkcKKO
mWnZ7CfdDW5CyuZr9mzODqE8gxEEROPBpyccZvapCS7WFqaWnQbxI57Ahn/jCZ2I
BCl6K90MD8ZJWVRPbIf9kvTBWCus+KGnahJBtm1FGk6pec8SYGA2g2SaBGXK0ddn
rB/eLgeCnZAuiXpqNjDlC3y0HbMDN9IN1EExVvxJKA+HmmCOaMBVzPn66qTRYm47
plzyr74AwQl9oA6FwhXiAJD7oZO5vAlBdr8XOQqFJY8uez3GeBFOq2+w5dHOumGB
DBO2SBLFjZhGL16FCEUwAfrvNMnEJOryLs3FqHdMn4RflVRhXpJKN0AOxMAZAurW
IfqLa1jtHKT8Pju4TP+75aULu+T41Jq7GLHP2ZkTxHkyW/NgL6NsMhy1l6k7o/Fd
u/wyMoUBC6gYDvewmst8mlC9miCaIwC3eALrUTb6BwQRz4iO6yX5NzkfVsqnWQKC
SfgSeKsN1vuto8wYQ2IDAgCMgwD3p6iz1woEOrKPm3VYaX6vncEspORe93Xej4rN
sq0OuvAgwFnuEBeYz7Yy3mk/tcya67tgLoptkY9yEM5TxmvhlTqE6J4lck1fWwJL
vez8SIxjGrbsLyRbQQPcdtJZQbMAOMk2ZBH+HVcqbTzEoikBofG/r4dP4vNXCI5B
A36dbFDZoWBdJJ95MFcOux4KbYwdhf46CUDAkTRtw9x3ODyFRE36QrZSOOJthLoD
hDELMiMr1aAm5HD8TflEj4vFGDFZniyhRWdUt/dmzvFjYFj4VzwDLBA6dNaHZ8Iw
BiGUBZrX3Fhl5p2YNc7WPfp6jNCgv/l2kYNL/PxkxmOQ60LUaA8/CngD281RA8M9
wd3k40q5X2GVUfrgmdTFAI29e2t++8Ez9pJd1g7VKQ5k90gyYZgVbcfDP8EkaUCi
BKt9mjCsbPrTYOyDFiSVMDleNQLRPolNBEozf2Q9j8MeDF1S6HJQjNWJxgnzgTRx
yNAmmU5C1i6D6yJDdK3jVvlUrh3CUkr6m5QKaStGr9HZ2XZJ6jCu52ozNIJuMpzE
u9gEYSuilJsEkyu0xtDknT3AG9cBazuJlQ73qBjsmFyMrTstIzIV/SsXIC2u1Rbv
0n/J+TNggdH4fuUqwSL/hBovNMAGJpUTs0ds4TTgAjevgCn3AKVMd0/zT5QrpyuE
votJMr/gpm+fehpCAfV/jZ7cZaFB6Qp/fWJy9X213blevEdYFhug6IxDG+AoRD5a
6eyVPK+r7QUBHQq85nlRBdlvfjMCrz2EWy04l2loCZ7VW0skdCA7t1tHzGbmbZXI
WSwnXSRmqsVaFzdpJoT7Aw9bhJkuJrfMbbgxxWIzxsM29H7ziF6zf8Tz9YGA/fpv
kC3CJkJuY8Ns25QGMyMsIMzzhcfHFLG+Wuk1/5Z5MTGn4q3spgasqWEv0wR/oLR8
abKrS/L3gAHEAYW90Tyx4LhML1GA+fjIE+R3yPnmHGkQYAaCh1BAG8sj8CSrgFwl
1IBtSlAorS1+dWzkd0qrUprciEhaBidWBMbP7J9J7PQxof96NGvgpNZ/XaPncf5o
VHFIV97V30/jrHm/MtaYk53I9VPZG/m2DfsilikRVSrkyQlvwLTSLa2VTOot4ESI
7uXedXvtFLjo+NgH3IMalV6PxL1w5Gh6MiLGZIDqMVih3Dy/Y6mGpg3WuRz5IXDG
FKVw75UD5sKQ/hHFjbX0OMNGfmrHmYliBZjepuBh5WyiDfckBOMm+Tr40yLJucO8
1SJGUhliLWy36cIy/SS/HUt3WNvwNVnRYc9X328bdAiBFnfHf8SHfovtgiDmtaGF
BgSDFtuse2o4rFS30z6vGkTWAEtufyz/WYqvK4GvVoUP3r42lvLcWy2YeutbMqWx
meCmhiPaMC5OX0YxkAYnDfK43mxLV0TPWtBQvV8KFJuACLxn+gIqMDO53uWRlExm
mOIaMSZ1AXluZLKJbrNhr+ElSk9usZRvu9btO+kgmJqR/mrDiZyaf+n+p3+IwVeh
tGP9y4qCiPfGcGBDQyZGcB0BV9LVO4TQBwIZp+IO4k/RuheXMBgA5jrKS9G2mVbq
CylB0uLYzdJ9GweIdHXTUxIi+olQrosc340HZb/yHx1B+FN/+LNkXcA+ix7Ag5f5
6ooW7GlXmI+cE4thd584WvIIxs1fapI8om3TXzqipimez3tQ3ZQ68wfDgikJwHuX
Q5VbU/gUfv1lO5/yaCex6lpBZJi0I3yqmAlTZmVJ76ekAk0GnldWNgR46hRYyTEY
uB7Ws0OlwyfdIWYVaNgN/v4/9jIXvGK7YzBTy1P7nCTidcIUD85iCZj7FM5awwEd
Fe4+la9MQfirbyktr9SnoW9jCfL9lf+iyT8QfAc9dQvl/y71s3Zj8bJ3nfIMT/AA
adkUetHCa0yl51cotCMeVDjL4qsSqeLabRXQaqsAWQSZX8UQUV6J2hRfSj4X6ed1
NKPz/7CBImQQ0mNgtBrWt0+YNnqGe4na3MYVT4IbdFgDj60fjQCjqPJ+7dtCe2EM
XUTgGOfJY4VtSNcyS5hCl7pCtsneGy8kipvqrrnH1ArizyGUIwnrbGV2noG1GXg+
gakLn9TPhFiEcOAXfrL4Cii1xCvi1Qh/woYsTj0ZjNpxZutCiuds9DoGxl0WyLXp
zHhyf7VwjkmZLNPPwvMXqFTve8dfP4iRUN+BnfQGnqTR8JADCxb7ECTLUVmBvr4k
J+jRsiz42nnti3EKHSmhU3Ytyn6rsntR/botBasVG0eWwC48AZp2+QMrtwnbIf6e
EJKO5cp2RMgkraTU7BzY83rndjEtdnFl0HhShNLaCRH/clSgLrsBs8kGr4/TVVA/
Cnp/YvjOz7M9yhqsE1SoD4E6gLVZ9l9qsjbB7cmgKdiQHHao5fBbgaRq7/Yik60o
QfQa1KHIpJtnHrvybz2XO1Gu35um0tPQ7EyKlJIuHnATyaH4BqmioYrkZwrbW/Di
jzddf6LsXcKT9w4Web9JDl+O5J95lgCr9KKszNY1Re3RS0j9bGX1iULNjSYkTOhf
ZZLBXsgzEagtTCAWf51DGObv4/rSxwm+HffvACLAnGdgoEv4CXojWiY0QcsjvfMw
OY54GfQ97jIYqNPddLFvoUIGwa7ymDPTusymKaNMMBCbJIV3P82SnTCP+LWCyT7F
wXETam64Lxx74es15LSI3Z6+MSLPqn6TPueV51naKfx6ZAwLM/4OsI2EtNJskS9W
SYXMVU8eRgXt8kLc/AdpU2ZM1lae0RNYN1d21aKVhCcKweW25gd8zKMXQY4SxYTd
19h+xiusRCN9shfiPgQodMmjf2y79XXyqRN/dC057iaZ8VsiwNNsBbHd+HEggNbr
VNOdwaEzaVDlxNcYR0M9hhTcXRJ9sU0zMwGW6VdCtsOn785AHIwO90Rzmo+Nr85e
O8/dTN2PaCoNoarTYJcOYIPDFkjF+Jhiy1Xjpb6V5EoNqUIiAhU7ozOTXZlJRvqq
fS7RMyaBF3JgXiB01tIyRa3nTjMCmiIo++jFfKlgJRls8DLQzimvyRTPr6ei4J1a
tJwddfeoCAV/jEhjlrivjNif2MXi8L3m3IvmXysTy1XNhoKX3UvThG7XQqqLDAPH
mJ4cxojlpmelORyD9NsHLzKVIFGHXrDZEzZWD7TL1Dlr9gfiiP2sgkIQqkm+/okj
hsIsajZiIM3rqRGVzD8iQy//Tn3n6GEI5CY5sesyWtBN1fTZo3wi71eu9TiwTWwx
IztSknX4zavwH/xXh1sE5EDIZxh3VQzTxu+ROCm3VvRxpikmwIl4urouVCusNbP0
Ms/bPSP2AtIFlF3A3UUIh5mj+PasEpGTT5K7rgGhxVgQvC5YrcexBBWZ1vZcEJjW
n5mCv2WQ5Zbjd09Q4uxJrNNmsslxXUzn4CzV0lOprXKgkXt/mpxsX1hw4quAT94E
HlZO2a0/DHQU8NgxvSEgvz6ek7/RHU4zVjpzdX9dw/zgfZDLP5kquGqVI0GA61Fn
QM5o5DS0oGt3PLbhqt3b14bJnHhTcRU3vXkPw4lUkovji4Avd6+74AmkgHzcqoOi
XftICL8RNJDF4ek/E/f/7ESRZjGTBv4/Fwjoo8ugZCW1LY3xdGRq9QRCWWs0xM8n
77c6C/6cCD8WJ9EtC2SKSdiHzXyJHqq+T8GcnkRZJrHSHHLnC+t6NbvHM6IZi9Ri
k5HQ1LexHL/si+dxYMKeG7gE0qpMokAU0e6/EgC7kCeB8fpXyln4bwBl6Hal9S/n
G6WfqjyarHAEMDXCp65ZWUp3vlikjrI6270MG0YkrogCc+DxgKAlPZSGUJTMJmi4
fPlJm2bDA/Q4pVHLflVPUnffMsO4vb5IJLRjK7d2YiGUxS6j+nXRuJ8n9FtVcaql
tmqPqREOf5rsOJZxjQJzlY06EsEQNJJeSzJubJIywyEV1xGdLrw7J80Ay7ZMqHWk
RBGqPAgLX8lRwOhHEq17M9PhVa5C9tMy+cw+gB6gS2a0nwHvrPYvkJmGg3EY3lB2
tLfEE2DxL7qyMRKWBlKXO8WMpBdGq3AXeRjV407GME31ED6lIZhFEcyMWA+w53kK
lCG4hUfcWxIvyHjoYbMUF2ev8HqKVrK2WwNCpX7gxyR5ERWrK1EJntjH/V4tvfFH
X/QagrfYnv7ztGsfql1AMMXZMjZw0QDKmxGrgUGS5gWt2pNxZhiunphdQTTs9Ids
2M9dM6w7aDIu3LeRtLoffEikMy/zemWp0nR1Buu9GpM6m2OcooVjPPPzMGgSATrM
Iz8dwQLVlM8Z/+BSBmPDEJF8WA4e3zPLpsALUO+Xn5uEHAXZMWmhY3PVq0McdC9y
8rdSsAGAqST7ZoXp46/PtWIa2ap+Nlkz9XITnxdXJi/wl9RfYcdwib+yOiGmztfI
QAGhCXeqSv3r6XM3f8Qd1PhD4iHH8FRWlDvuymPiDzKF39WknJ5WxffXLidXPkr+
bK/vfdvqAKq9iY8IvmoQFlQ0nQzUqUc0l1NhflAHHqBVgaZCGk7NtKxUvp22cu+4
/Umv6jZ91nrcl6Wg+9EzvC1WdOSXWI3ct+sn31euZf30soxgZCciHtODDg0UsS5t
ok1/zVuV65bFU8BJyNqwyoX30h7uWqopUP0iQq/BAL8nWXBKmkhKiORfOgWO+dE2
V2O9+vKJhIxG4w3UVpbG1F+B3qk0NW2l1G1mpdczz8gPMyR8bCb6vP5WgysOmjFd
sKyVRpU40+SUy6UI1qBjZeamndkW2YH1lrbF7EaiWejVAqpYvaadQD1lDE/UzV6h
tnPrVKBk+7DNgJlfQsCsE64ohOu7eN9bItM/VHd9rJaYIZsNr2BkPDLdXKYzEVTB
O5YsNcR9uHnLay+uP+6l8dxy/tUBtd9DkwsTBSo3h5rFv4JTi2ed3lOqp5tyxQOD
TBQHkwLEGwsmkWDkN5gsjhf9dS/AU0kufrP2IfmWkLC3Cw0aHENO1C71H3Y3pr+c
QRMbCkt+2jk9G2AI/1PflaGR3DKKhojhjXrRpQOzznUkjGc8VUvZ1SX+6CGNUsX+
JcSQ1h9N9rXNELFP/2a8Qd+iU4bX8NaAdGrMFeEI4j1FmnAmDCpV3pxt4senStje
0n8YySnvp7bRJcXxajO50+HIdgL4uATG+KNR/aoEIqua7SdpsBrhtDGV8KZL4vg0
4Bqf1JDjZ2nlDtz2M5KvOLxfBZFTGq3HNB4GUNQtMlIrYZvLQFMgsKE4iR/mmuK9
c+q9JV84sRwCAGSCg0QhuyyT5RlkU28ZpPX7/SY2sCccoXLdo3TqSo7Y633mLBs2
MBeVjvAHw4A60ki3auEyOVMkYGhoEg5J0H1rF352p0AUpvyQzFonRoF23rftS5Kh
/ixID9BMDZ3wpE/XvuW3dMKL+PyymR1XOife5Zxk6ngq4TRKf6L5t7i7jbWUM6Bk
aiEoC9yMEm2nvroZV+f1shacIE8b0v1A9LMAPg2XvbaxULNbkPlCplHTNJsGi1MK
I4hHQHnm1C5bUi5n54Ccq5x/oyqC7KgV0K2xuiIfO/4QMQGImVe13LGLtaR+yLtg
yb4TVYPm6W2+aG2MM4mrvvhP0hrrWeRggAknaepe9+34VE4XH89BOg+yvVyHqGMn
zxwnfZ4+e4wmdsMyaUZmrPF/iRYrjSpMruu3lsCduSMUQ34EFjsZ5tQ0dzLpmff3
Q9CH6g9HtIV4gKvl+ZVjH6e1fajjW5hf2sMSPsqxgEQdtT3JipjBPSnv8FUg3cVF
NSDhP7rsbCMMcbEwvEnIptKaUyp5IFZpiaJwy5GWIK5xfZwtbhG7QObFCAmuUiul
boRN3UK59hI8j67YN4s6fkzFw+D0GCAaUu+z5LaNrpqj0c0eEg32vfJ7qbNnZM69
GckdkufR0OvoQ9kqbJUn0kOOxRKuaZn9oHvDqBVcJjfR7TfKP1v0Y/FwGnRMCXbO
ldQW5HdTIm8nGfMeLetLo+RcnvC9Zq7EYbMfT8dJ+RMUo/U/uzpGEMGK3xRsnCCk
fQWbd451aVxZV5VEmKXbnhLIfZNtjWdHw+QIyF793G3go/kDWtyMYliTJXlmu7Y3
kXOddUZ+SpmQ7BB0ZiRFWJ+CVsf3PvQBmndeUp0y8DvX+NtRR2UcrRzv0p3E4ZyL
8p3BzxQVep0wguSAvnV/4gGrTmfUIRQVzSIpibD1Gju6KDadG5mmb+1QLB4j7CR7
P8UfKzVj4Gn+D/e1zRda7wOxgI97YNRQ+2jqgBeSezIgEjU6BKPgiQ1aulIaHgEc
YWg88DnZWJiGvut6ZXqLVu13LzQLh/B51k3Cde4NT7z3g1UJhOgV1cIIaRIiQtB2
WCBu2XecHVjoCUms7yQWqO/YAEdv48z+9dQAFphlbt0A+EugCyzQbKqaRG7cGFfI
v1Cg5a9rR/9Y8dGmE3Z1qjuZVFCUTGdyu1IcHXdomvdZ1b3/MiguQuZZ7b459OqC
9d5YCeAZFy9SNkVKb8z8SckkW17ogZ5iPyL1hQCEi0wjeOIGKGRAd85RaEUcRtCn
snEeAQBOpx2UJYLCz9YnFfcXD5/KBMQxvoRF74NMD5VY6XenRUdxLt2shAb42plh
ocWVfpw/+Vy59BnGuorpMils5921IlL6f6IRzvbIgy4sV5MctX5Nh4G+YBXBRPLG
Zxi0/Yar2qHkV0R8pCmeyPcBVNC/pvC+UgFISsG+Z1MaucCf3h0KT2O3gj21IA8A
qkfG8/dJBUfTohepzrTbl3iCiUmvMQew0aCeepg5lJxUq3r6UgMAKsn2Kie80WhJ
y3ac/g/jlGZcDvupiAXc92tfM0ieeGB20COxBFlSfBJL9apbcIYSxMK0d9zVS/M9
BrypXJSumwDtFqtrVp8IqW9Vk3ljmU7lPclkMgtdipR3KYKCAjqOywQ8r9cHYFKJ
OMd5Vg5Mc3QunZMdiGHWcE44d8GGHd5GBuYaw34HgGa2bLvg/ox/eIlO7qkr2ygo
YXknPetEeC7WLUfdbMcyEyakG8QyXjURq6C33qeUK5DozKX+kcqtU2kiDoLftQt4
7UurUJa/QgOnTpHiIv1CJVFab0RhzcRseiZ9/qdWYr951XVRqnnAi1GvZOVVtakG
/cb5oM3CNkZJQPn8tllrqRXjjzfyQnLFOj1wgOmIse+WYDW2DWOR9H4HZx1PHYFz
ObLeWE+2QCYc7c0DHqEJbpwQ+OQLu1w5UOAquoSFBFiSYFzY3b9FrpM4DjcWCA0C
YkWeFAWw9GajaSEklzGVFShu1lrEZDiDJY/VNHdpeqQE0K51GCLRQRjYA18AHXNM
arXcvcR+aCUhBzDGCeK5Qha0Lie2FY3slljURTHebBN+45c0KPoNF5ViXGAJXMQz
s1Obb+opy8xfX3HUKs1mbL1jd4asTyz+5CFngS9T4Q/hYDHrFrvk0sNCl4TSYj2i
bbAcaCdd83nuN3kLXsP3cy76WlQS81SJv7YVQQDCFBK6C9Kf/808fiqtdRa7h+XW
MBUps4DcIMZMIfxByoDo7Q5zUd6nlQ/uVFCblP0witIg6N0joBeMJmwV1aT0VNNr
A2p5x/aEmiHNMvd9AJV3AKvOwGGuzjTeejE0uTqVfFybxtHqk3Q8CtVr7YX03HIk
wEVx1qC83dEYZ0tOh6/Oq2CLmblggvKxyNZF/JMidwp/z4lrPfmRscqXw22UcLqT
WCa0aviN9T066+frvlSmF7oJvBD2TMR2pmpVyON3iUnc+BDfdcZmgLAQWLpApu97
NB4Ghr+z+pOOQ+QoMrAcJzzqs01oLWYWecyqyULpdbh9KEmt4k7ZLc4NxY3IKSNh
GrReodJb+PTU4eF0srA63aluHILSKJ2nmH3S2E34+/wGs39PpOw6/ryS3A+cksWQ
HILX50sLC5As63O9AX6dzaHT94PCsL97GGrHrdj2MvVlli5UgNIPbpbJexIWZ0P8
/KrY5CM3AQxL3iSNs9fB1YT59+9yG8l+Fo+8A8A0U8JIerkzUZeM3FOVFaiaK4CF
Hv4/B97ZGh7U0/RfPrYcGxnQ6wfM8WnbCyY6V/Bp/mWkpcwvn0qeN97Zf3zk3TFo
YXCqoFqnvM0MRgQtS3ifQ7GXTCp2YuCTvj05bq5JgD46/CqDUn4fdN2WCMaA9iWs
WruaEvCEC4m0NX4IH+Yp3sX6IJfrc2gLpc6KQ7NNSvkKW8Gf+GScavHsmER2CVPw
CVWqMcfj9XPeBIbBrJXOgKbRwCIoD9PmzW+nq/QoGeeCvPB3vdlnVfVmsOz/1g2x
wwbmdHCcOCIeD14O0XrJBJer6xQA52oXNXmtuyPYcs8MftFI++UVKX4Jq9gGPrwx
Az6RTIgSFPGjP2mAQoJzO0YumUpVHgKBk31QA4gk7JMgxHBKNlRXlkRwkLvpgFqY
pwXNS0xwJbtvWjoQ/URmKTj+SlvdduGZaCffaSWP044A2rbLykXHcgvxbMmVcxx3
yXuUZKx+pvihYfECb5Oj78dOoysTO71nt2dAGRE/lZrSU3Wkpxh1W3A1hYaz7ukK
7dHRE7kOMHtMoNTOPujZlLzDlOAbmfICJSi1czNeSpOnBaFOJrMw+tg0NLlwKJ2e
AJ/pCA/Lv5AL4T1vmYFB9hrwj6i+zW5PMDuPGOOeehIXutfc2JPjmB5VA2n+L58j
4Ak006Q8gmeFBZ6OWjHb4qqYCcbG3F53H2HBTirnep4CNDjyA89m2+6Sh3LbWIb9
DgOyJYAvNid086OrkOcii/J+kGjhSSEi9dSUCrzZIFsvupZW4MAozPBrI5nV6Nul
sJjV9nBNT82XuM6sfZOV8hybPH2BvurzzZ3N+EAJ8z/19sKCurDTR4oNnp7pz9nX
jrTpJuHMS45ghjoZnzSsSRmPvrf//qR/oOP1TDZgb3rAW/6jqKt+vFBwziFU96NP
Q7BlDf7+PvzYTYwoJ6iOj6UbnZcmndcmTcaIZMMp/AcyWhgPaZ5IVQ6/EKhZeJIk
QooFCtR8SRXoUZPM7N8RwOst0NRKT7oD8KjFqs64h4UCS2eZ9zFtGGma0glgyFMZ
r9PBSXetNQx5RXiUVl5GI36t8B9OX2eeow1qWCcP2j526N7yYUxJQ8T680f3MOGs
8kDYFjqRbeFcI1wbXZ10oPeodMzXrnA3oaMDjH6NQwA6cl8Jiecn83OQUYomvZ94
McU450B5SiDUJ+1L+cK/b31W9Euk9KMe8h4BHfFlBjCIHqQ7JJ/wpTu0YOuoGAL3
An14CL4SSlgpebLqYol/27/hRaLLS/Wm1PVTuImO9mpZfDQpDLoBJbx1rOvvkvmW
v8IjSloi0rghOSNTMmMHJKFHToRdU1QB3g5pMx+HxK4l20bN6Ulrk3l1UghSoIg7
ROFCYBX8wxDRW8NK+3ZNY1JCEk1CsAv/FGGfGNSB2CL02Ml8g+TVnnKIBlPH7DcV
J2RKf8P4ZzQFJTpxcnv2lHl9+VmRy409LJYpsFx00uW1diuyiRxJtIk0laC/Rwv5
+y69PHFowkpzgVUaEDyr7773K8B8fFa8roj9QqJ+EEoo0Ng9ySJ/qw2Kt4QDTsnm
joDq3aO5N9QkskdA0QEXYPB7OTvx3vDBezP1LlHM7esgPhrVa38zkTycb5Wwpg0W
yYtAKTDswRzO0rgRejsJnAGS9yl5sEsId8FHuR9y+Ba4ZaIKcaacJu+pRT4IJQkC
2NvB9bA2W5IWPp55x+eYZHJMunmiQO8gZoQmQPKZV1DqLa85A4TmG7aKMUT5sEdk
EGHJZdYAcPttXDzZbwnkleNODgpppwp1Ab90H0N/Cwl/eKs368AgRdvShrwfDXIk
Xfu/gHMsY0h3HqXkmwl+qBuGsIrc+hw8SquJoY/u+chedXQeHYbvguMetUIVD80h
Dou2fEzgCRIAuufjavuMTxGLNm1JysJoX562CQ5OoYi1WwWJUI0mNZU11IdWI6Y6
E8eScpGSp/8us85lv9djv5+nTSWR8IRFIkIKyTSVccX0eqJlwbpyueHkkMhIA7cS
oWEY/+U63RPFm5BpSrXLJrfwt4X/ZQLx0J6t0c0e2coAAoai+HV0dF8be7dKDutS
7gdmOkM2oc7dhzmrUANhKLkJlMBy5AQua1kvO13qI9VdYBVAnKReqrH/aYCPnVEf
3y94DQEzK/i5WmlRdezQd6XFOfn/drgX0rJMYlXdINTrzelmxmWRyIa3ciSF67U7
E7iluNjS4God88xMMHruKEKEiJ/hoUCPWpZWu16AqhG6ecrrPJZEgaPs2ANRQbIx
VTDTB6vACf13hLd13UKveEB7cax5Yh86PRK6Oty8CNF9zy52SXpJS2wPJRMFm5Yb
FZiViWBk9Rv6NbX9n5Iv3J162D2kUZZA1qAjtX6XD1xyIqNbucp4UbU9gNdG6gAm
erg09xMdi89wgGSH3ZOpYtJI0hoKBWsLBmsOcdCX8IyXWtQ5zd7LygamHTYxvu9o
9IFGXq5zUrsqiq7Y5nB3/iXTBN8GKBcGVyb3ttbyXWa4iDVUVPAIIZFivA7+3/JK
t0yY6HaO2McegYErMKf8yetuKj2V+bUNiKYAjdevhzYJTPD0g/zX7P2aEyLyyrwW
CQYOAlxk6MgTUAh+lSQ4v9uxbFVjolgw5LjTRdrGXQOYLP2RTA9hRheCgEY49JwI
skRwO95jh+uNJMqbjio901LDmN9o2Tn+HS2gDsio4p+LyUlnvPdtJqxEBOr6Egiw
y7j7xLtQ0jkWzHqQ3MbJ6u0hixbCHsp7j7O2xVSwYwdhoB7cpwBmsRJdqelTh0gE
8O3PsxgiZ7d4wrH8mcKC9k7P78zhFuwbCW5WIRyoBJYyq5d+QpodXagscCoSbXog
pbyeJgVdswByG8R3SdMY5GWEcdwETkMy7lPsnqLLThVLNlZ1w/NaQAAxkvGWvw9t
Vc1za1ffA+2GYZNOGDHmOWwrBVps450Lhgk5oXBTTFTa3GgTkE64tTQoPJeLrYwt
caNlPB5pkor+ReeEATDd5mgywmdDID5YCB+bzjSSi57ps93TdYmzcq8oAl7e9kE0
99HCAiki467HecS6I7/ZTP3La6ZroF+1fjWO4Gkv9AWF2glBQvHV+QQyeG8zL1VV
nRxmSFbiJlW+PId+hiBdo8w6oU9255XVVOR1tQgXKNmMFyL8N1Oqx+OTwG89QL+u
MbeYgXclbYQcE+VlL/Xq38pF81LjrZDq0LZT1E6+qCB8jP91ypt4sa1FynmEBpN4
yPPEwbxPRBWRjAZPXiVKLyPBZn/SQHfMST7JzmV8CJACj9ChEwULA+zUEuHNu+yS
AzQO+QLcY9cTtxXOZZAlmsNSIdOEkOMRm4DHFtFAe9rPMmA6xsV5taixzZ7jVUiD
RXoN7kkE2JpjmjeJUZ4ibUIU939sxfIj1cQOm0EIcdc8qH10zCDDZRVMqzrdqCOK
jLqwXtxVvZrRhrYsxmQLAhGlvk90masfnIrN7xJrBDP6leHapOKl5UG1dkUEXpku
magkWtanc8uPCHJs8xLQCs3+ST92mrweWjakvBHjaCDTj5T2+AJ7vzgMr5uaJr0M
dM4Q08XiXS+QUyCEaMClUbbRDhD9bGw7N1fbvBrPYyB8/HDKrUjzCQdrsiprnaBn
Swoyv56HSd4dFXS1Yhy621JSDv7DGFmmf/P6DPxcRqK2Nr1EMVZY3R1ggRMs95Va
fkmnig66UuvTOA60LPYhOWU2rqckldbE5OFsjXjDoh0y2pS8yZGaGTOG6pc6BD30
6lqtbgBNA1DghwpyKPmW4toJ+Lgjch1ITb8PSk+eGbPj/QJAbESS1FgGe7Se0aup
1ObjdCzLsEyGPiblZIh2zmP+FmhJ/qdc1uNtEl1WBm52Bk6MsGXRFsAC32Wmd4yG
HgNulIs4s8IA/TwGDQZ4alQISF7M28+HD0mtkjgE2re+YtVYJL1rf+QH7HSXkjkB
gnd/WwWQMdJAVHdXh0Uu74zQRqqa+U8ZFLZKtzSMrO63bKrLlsOKpaHt2s0gCrpm
eePL76hV0VhUegk2Cw+VN1VviWdD1jCXgTqcsB4C5OCnqo74ioEEOrim0odwbI7p
c2tX2akbVXIP0UPr1tarBK7nS4q195l5bYpXHnyeaZ9F8rQZ+0iFQdaUP4wNv1Sz
wIu0IeBXH4P4smLow72B9QBOnZQpfgvo8mIDq/00BYBoui4BJhjHUyZjG2erOAwr
HAnHyPtA9778toBYdJdl1dA8ZxRq3ENA5tfqhn8gQxNlyghk0XTFXgJCu6Io9Z2H
XB5AmjW+LN9W/tU7xLogc8//UQH3iMAOFZxpIMHXml1J8AG5ErcZWZC6ru72xgel
zN90r7e1IJE349sYyqA9ApJv0bIufpgAsHMgRa/Nvf3hDTxjSpTmSW2PE8dlY09t
9c5TmxmJluJWi6wSiJpSdRTBjfTIWQis4fzyajrOGKVwL1D+qCl2CS4uGwjNctLG
Tz4H7yv7QD8ulhefkqAtfXUmUe5p1Dz3Rer+fznmU6j4JAeozuR4gtFvzUaK8TG/
FMbz3yVHTczF9UJwLRLisTMCEfPBfyhRbLN3A5xRmnENRhYPzxdic2Nv54Hk8I8l
w/XP+1bV8QIXQkwZQrECe/GrdiTjbP4G1h7Bz2jPzExPIemRVFiwRbxlzzeIym4o
Fh/qq070137mPg62wGYf7X++Rbj8VCuT+EWY5FVtQg/SLDWONbrrAtwRSld7EAt3
ayI8PfAVndDsdioow7R9ouXBSQHL7XoqXtupdXxWzDX3/yYG+5yAMg2b5olsXIvl
MU/rz9UHXeLFrykunAgyntZIYfoNhBNTba+HgrtK5bITn5ZCHS1JHj5W4aOfIzeT
uk7b8KF67UtaYTrho38zvvuQjg4HN7bF2Ocqg+PGyqCaaFDbakW3lI7aABHX1LiZ
w+ExWbPGGMJenCXsnfabroL7pr6Bqc23alNfYdldsIAa7OV64ovDbDMqcAFZM6nm
zPs61+sF1EtO3miusm/dZRPvtAbzAG3XoJxJFlCAr1QFJgEJnolDH+zr5LHbqLy/
mZ4+lS1TkCx3cB5X+g85c4iSVbxpEjGrxb2ceNkd3SUY+Pd48fn2ckac9YJMoDkF
v+JC9ta4sDHp86RCHPCjV/JGMQzJWiSpvos40qZan5I=
`protect end_protected