`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15664 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
akBpHK9XojjdOyFTP3pOwt8EsNLFsJTOkvPGprz4M+GOt1MB0ImTOfr/6a70bVsx
+fqmOMnfY+E9uYR96fxzaIoPprozPw9nTInf+L0YwXdXf2vRl/vh1i63U3PRRJl0
2X7nlI+msaPMx4b3Kn2M+/Wyu1zhVCOZvQ8/PNow6k23VabMlsV5eZewh8ET4E7e
n09vnUs9OvAZ7xwEW1FO+FBBozOhCzt+MPLUcsNeuDYx07P9CqUzkApA3hV6iIEl
eB7xT1BhRKHBva453ycfDgGy5yDugN36t5wVWIq1zSJlj7l41K311pT8E+AujOYe
N9T+w2xlwrvew7W11qnrhCuyKUtAFzknNJsKm1LXlYIlCdSaSHGB6Oa5I36Zvb0n
RiYXNcUTP+OoDhEn3Q9bI0mTVIHOtRrmP48pavbhW0wGJmJdwfFEX6TvDZ6Hmkb2
j1JB8rpGf1h1d5uI8A7llo0LZnwencweoll/y3WyIClGdaif6CRB0ZwW7PZNVsK5
IQ9rnYox8ENVEdyqRsB36C4El9qKGz7qPRunVd95vvBYfFuhGo88Ng3ShkVZrhNt
Twr5mBvoKEc/WhvJp/rNTtxNA66e3WeDPH2RxvxiKghsBesLl8Ua/IiGkSvHZiab
5L1E2kbPldIo7UNEi0oirYXqZMBwrD3k7Q++VMD1g95BwzIJNRFqC5cw7es5Cs7o
tIh9YlMbYLitd2IFWc/n5mseUPW1TUF/RruA//QiFswhoU4z9tg2xuttcCIcI3bA
l2BYgrwtxaB7KYgIkhaJhUJjSV6pe3/pT3CVgBJqY/ky5/M/ASstbBFLXUYa5GXE
Bk7E1ON1rCyVLieB1EdLPYVH25x4I+pM3O61RO6EDh7DhMt4C85qu9rFnsmEGRKw
T4sKezr+gfukeuKJ0uH7MpXlOd9N0nA9+RV6/cTDBpTVqLAgAvzA4CLDZd1PHaNf
qrM9fQZq2pXqHRmkb9zxsFGKynKv+t2I0FRCBWVi9T6KhkamaZ6adwvr8znCOVZ2
5RxG5Je6WW381+8oydL5DD52AXUyICJ8Q3roUmbVUyw5tGAkpzdlCDtpUNBlyR7E
SgGboxZDerGydX6KI/FQyHaLEjsrgtf3jjgPudaKdfVXf5mOhM+5+EM9zlkGX6BO
HzG6wN2HdodU59dYz9AHJIrxOHZu7PzQZPNSoKaLa28uCCyID0ZtXKygNr4WPAgW
ISqvEsoRQpkwgfZ8xXjJk7Ay08y+myhXsvivW7jtloNXNJA5sONwV9hg97EYNCc4
seAhw6Gxpp5iw8ZLetuPOjU5GwMTbjOk7sKNxQ/9355hpKm4LQY+RGw2gZTQhUX+
xpD6qZlj9spI2rF6uCIoWm2vf4E9e1UH0Rn9tSMRHnZuCnkeC5z8XgGsdapAePdw
jC9Ytf0dsU9UaEug6QhghdWBxWUxqziHrMiZWwH77LA2ctNO2rPBlTJw2pngtDHx
Oc9yd109buKZwuENGlGGzdX0tJ3doGigcSyz+wrb/1tyovG6xpulHpejWL8VNTxE
/zBcvGWlxnk1WZkLnJbuvG6yhZgkxL+xygHOglDYSV8RTmzMR8vUwm6CQQffekfA
o0+pXfi+T6f4XmZHBvwgAuKAB1Bw9yqBMwtK2cHWYdZrKee6/UpqxPVN4VKkeMTB
vIFLGdj/xGMaNOEE6O2tDaM8Axi1SDF04COCBeHO4deE5YBE7UZL49uce+XqOxcN
3wwTbO+6WUfq0Zqkx34CFMStH7ASDkLbM15MvqdN7WBuVILTmGYWCNHtJsLOmzNu
PCMsgIlHFUpCxtNIttpLf4oVTdg8S926r2DBKPDzBa3IcHzsYRLMpjXdK13d97n0
yHsOnTpCHiOxZvjE9E9C1kGVOxJYn3CaBQxWcfwkHA7Wqcu9il0qDqbf+MTVi085
x3sF8XezGS9Z8e27MmjAd3sgEAUbNxaRz1klCRSpkjTElK79dKj+GjxEuwtrSQYp
HGtBlM9yBLHwuw0cP6FBpbnhMxJ70tskrrlHmbuQGx2qT3Vn+HV4l/B8orefzDqL
faieGqo7Yo8mMIKprZQWYty2Pp+iltqgNyNCyGExqoIPlwezcLGY6Axuz1koce1E
ZMKfmPHeDxFplGh2LL/jhZIzpSMgg00F/7LSLHPhPuuwpT6m5Xn9OTcZ0J4xeFr0
mWIDvvQvUZfrSZ9PS0aQcP70zudJq332tBgGSaGAAeuPnOrJb9X23H02p++mWa8w
3+bERAZ9It8Fv4rG0HZicakZUP5LFaUY1OoVlKzW9C+FMs2Rxwbbqa1c19d84rhd
3m4DolNTgU5iz0AJp9z9A3vIfBmAYLnLhoWR2X7nJoieqfKi9H387qcL4Sdq5Wqp
/XESiaAnDZN7hRHAhx51nNPN2dtW7SUGvY9lpe2Rt/yisCFOwCo/I54lyiAb66hC
A45L44+JbVNL+Ws8OiTxJJdX5LoS4p2+EThtwDx8ubAyuY/iPzwkJb/P9ncqRZ4a
3+Ooe8MQsYKWJY+nrt0hwddtTPsdI8OJgjA9XiXMkrTwRq+sXLWDfPRG2RhyA74I
EAE5KFoY9pUETTrAVzoLFrrZmHxBjmVrguMqhCxtm6qbQl14SedhYjsRW/5FjBhR
lKTua/oyiXD5ZltIog7EKT85qYOSLPCzq5F3Y8OL9t20Sl5uHmDOzf5Ri+9xqeQu
JdU1NgYPgBpI5zL3kzk0biQBgypg77o94w7WYvWuBocmqHiN6ApbAOHhmA7M63rT
GzgFXy2IotMC1pKk8LR7NDAqrfYa9nG/M+vVSJlohE+Sf4FHxvgPrI3WnJfXeako
EpMxxMvlwBNUrmnfcTOkLgzsWbpbsRvbQt1RpzxYXEamIALtaVcqhe+rMbkue6vS
cqynOMVi0h0TtA+MxmfZHjgWFYz/fbtELgLP6Jj0G7xQIAdV9Eveyd9cgzf48/3O
lUjRh5p96CdOvTK/7pjmqYEOJONb1kqEGcwWZrLJBSiXCVnnPmwCE0OgDkX/R6wM
YXnCShqdOMrb0VIfxO4BFQ616U2LphOXMXPQMFeqVAlZ+NO+oR0m9jcD6mUklg6C
TXCRGkJ30Td8rHGokxc9JYVBSw/CqEb11ea/caP4ia5QKG//Btz9yVrg6SXjYjnp
PuE3USHN0C+wX4tfLA9IY8aILm3O0b/HMTaW5qJ9Jwu+Zb844pfSNMlwXZB5I36r
80miQsUa+jfwQOd8300FbaydGlOUnXtLVDGXbqA+RbJ48Qd4A1It9EwUu4WSTgov
HPSIbAdR6559l+CBvFyHP8/qqs4LbWklhbhR21vd6pDO4cBeFs/GMQi5B8HXPAJS
yDHRbd0NoAicdPcS/kVWUjkdFQ40eXusB0HleLvBO+6C5nIgYXZy76ylxPRQmgQm
/ET1j8P5oMFs8uJGs6UWnTQlsJwPIcA4jrSq7DgzGv5e51zzOZyGr2CYUfVjbXGW
PTotlf2X9hJLOfLgs+SvuJwISYiJRlAcA5mcC4OcxbWFVGg4DhuTVaRY6isjsUW7
vhBuZb7PeOyODdJg6dk4Qmd3JQn0YamYWxm0emEshnDzO33V0vGRMbBd3Jn9L/nq
+C/eSWi+GFQ5COkPRJOQJIZ3S9AriwfXzCOzM+dCxnkDlQed6kDAeYg1vLlx7Nko
/UDAfecsG0RkLEEMi2dvT02FqNdroe4wTxAYh3oC5Dx9QGgeIbWhFPyFouu66Ffx
XToc6Xg2MyRCBZsWhHangzYm3++yiK7w62uDrCkKVCNK5RWswp+PbYLzkqfBHK4I
6nWVObohJTICSqxNxJvJ/gmZfXNo3mr49Y7cSRsVlUFoefCkTHZSpaKFbHWAuyIw
KCbXWQjH+BG5ZzKnv/pcoResGfs+SGPFypXXxInCzqfbwr05GXL9mnU2bCpGCBi3
Ozfo7T0I4cBdD29CntCgaEpXkbzG1bQIxYAewjtGQ8TxyfEQTFuq+Xluzaz+Mc8U
+wGpQPk/iFx1QXG1l9gZFMbVd/OlvFxXOTjgSDJOKSRCf+xGJclPnZr0Vmj7iIuT
66jp1DPr7TOwmsI+lm4we7Amd49HXx5QpKMazLS4u4rcigqA2grSQVejFhCZN580
o8Pb+rua19RAywEa6p8dH4cka2QOS7WXcfzh0HvMgu/96JidAbmuNDgaBeG5+Lx1
B6QvweMKUp+mbzI55SQwZ8osTgZxewh30NYPUkACw+Yv0rmvM70ji3IC30ZlfSSz
bD4SA5e9bN7DAJL3Rr05EaAGUU/lk4tJv2XxwDNz4yQIM6wkOdM1bFnO8HxwNfnf
lWsbT2iOHMXL5cICSRFc501L86nBUDFbKXRlzrFAAZykGWUOaw5LPzCRW5VXA+Md
GpKOqxfDKQErpgCEgDamxzKRleQW3soqfoLPIxb8AdhQDvJZnHkNc00SACjBTXTp
AEEq9nYfwG3+PLsQkI6Oup49R7MaojricH53Vgbwre9WMCwJssJEmCjr9cbmbXIj
w+cbNKJXCMIcyw8n3a67w5fvOsy6s0zuhZ2ua9IPKqcLxwjjA/HmRlb7yqi5O+0B
8icUDV628li3aAUU03GqR/FYgvd6jpRNmpCB5cFfDMfZ3wxHNi5mdoZmIxBf1i6q
nh94ao7fYTB30/rgJUWqBHP/5eUY/v31cqzPZX0C4BV0zGGtl3c5MbjNJmVxExjQ
KxQI+JNgmrTGo1FzmONFiNoNN4Td3SnwCAsOGZ5eErFPfecByCjcvfdHpizkHqej
uvUnKLb+ba4BfCrhCBMnUwackwsH1kSXNa6ZDJTxmI1t+9aNigpjf3Q7WUMT/zRb
2aYty3opAmYzIVyYQHIU/dR9MwtkA23vKmMpTLuv6k26shug8NWM54APzCGd5t2l
wCaN5RLzdr1aQ/GAvP3Jh+JpT/VPiqfw9IZDAoUreipGQ3RTnBBn5ibkdnOgnveg
S1PJ9vrh6yAwjTxvUzw4HOmo4eNbvAOr7VEjL2j+S9IOgbkHYF6zbGRnMU3g8iEG
AFWvgZ0DKtzTSHHl2GQvOM7a6ZUvaXd0iPzHC8ifcG5QJRShKVSgWc+499apNSNL
wp3DpBgG3IxRzxi1xP/2DZWSyXbtj4BajNd5dEqkEDT60l94N2UiDa5o9SHH3TGf
lK9gDFmiN09OKNZE1A5EwT1o34cInGteA4NA+qcVIq0Mq928WG420ad5vsA/KF55
mxwLe3izeWirP5FZ3gmwFUHwu7Uygz5ViII1VoJUv071oK8nLpTpV100bkRw0RqH
qdt70WeKfSLDrQMhujmxHNlNtOpPeaf5H5FbAy9TG/x7PpOnUZjian2clGVeDov+
Ffb/Cx3C/DsVcOyY67fMqmpav2oshDHMcwYh8QWCppeEvXhTSIy/fS/UW5aicU2o
s5KJo3uYLNtEBjMYqnyrIGpX2hSFb0PYsBwxL+pCslqlIFXQWXhtUKw3msTsZnjv
3LknMCilPmBJMqFyucyqBNaVIGKdr3AjY5yYjMwApRiT/zJlAKcrlODzAUAycVKN
Y1myn5zm5DtMSFa7Yx/2wNZ0ciZXyxF+eblNFN5kjJVH9X0rIgiNqx8BcdMkIuQR
ivWITmr2rXxeAaaanNO8VxfqoI+jX90kH8/zs30J//9jPL8azR5qdVvgCnrZHkRC
4KwJcHl5n1VdXb0e+NwS80E8ckaQKtsLFPi3Kglm78tvMpirXXzS719geC61pYAR
/gRa8eWT0xsbK2amNU6SKG2yTSBqQsafzudU7roVuULODjXNLc5T8fDg/PO5uSMx
D6vws/TpsA+lYMyTlJW2YQt/mjTBnodNQe2A3HlWLl9j564APvIVjcOPt8e6T+Js
jwOLK8E8AGKMB9v84UbTKcwaL/cSLaLUzXc4fwNnzfAzi35ddbBHVGKXnovCgmIV
ZHaG5SMALdd7Yq0GLBpc0twJpnCEksxNM6uy9y+t06G1cry/96MYeRRmIYGdgfs8
b8n+iQyMM8HQQZzpWMnqVKAC58KpVvW/GDQy85zovMf/GL63aF80+5+tiYi8Lg4k
i6E/xFRXX2/2exPyS5W5GUxJJz7Cjt9CA6H+6zwSQ6xj13/5PjL3QhH0PYGkgr3m
xv8LPFhpy0pDBZqLdlU1BQNOyLn34BPJmpJRpCWxTm4rcaHhOoGHJXp4acrMxShg
dT0iOXvNYjcsps6sZ110W+NDHDxcQbt+a4Gc6f7Bnbb74GRbD5xqG1H40QTIG6NF
AXxZ+uBseJ4DpFqyN7DSm8UfHGy+BYtYgt00VlleTdHyI2mjkb7G8ZB6a8e5YDHi
PumaIoCkHTKmeg3avPeqvkqNH9cWItqKlTosCQrl8gF4KccJqMNhYP6mvmnPNt6U
54ATj2N+5Y7R+CUqABya5nNOMNCA4hjWBNCXHyCW57lgxxeC4T+WQH/hSPMVQ1Nl
ywnVcsRS1S9mSuOBsH4ZIwR8ZLuJTgAAEgPnrnB2nYE4+QgeOEgCfXyjk0XdMBLt
RoEwBBI+sL+bnsQSSwfLon9aW6EGV3k1JyDaD3yRfg2G14WllN3yAlxYmw4NMYVr
7zt6xeTc5rLq0QF1EQ+HdHDWRbwHOclxtSz0odEgFtv3UTynnKreQa7xAVvCo8RR
JFOj4Nd7jVvTLwPN3Q28n1mitvHzKRgA5H0rsl6RIjY1Gc0LB6kbiLhhu7Px1V0Y
ysuqzqy18RmObYuo6DMnlDSf/F+leMDJR9W/OCh3ZfPwTASD51+tpnzc6PDPqL3U
JBiK+5HhoxHGwwD+SJywsdqwoGVXuKlFF98JFv0PNedjM0oczP6qC7urkrKD/ziz
qcd0xo28QKQ4h4GoQAgxwNYYmB7SHBsceFytwKoZtU7nW9l7jrBhFqnTEb5V+21n
fUNpfQR+r5Aw+4+h4gr53VAiNl4rkGyL3D4sKwzKGV1Qg7RgZ8Qeq+kAkbgGNw/t
qOaLIolAEkMke5wHyuJ+JokZxpeXm2VI3hrXLUedJ2zMR/n6yseM0dVutgKVHCGD
3/W/hDStQZGY/Pi3YdyMIf3Xj6MdWIdCWopLIzlJtxSuSvcpowwYyYxnnJWpziZx
YptF411LxOoAPdK1+oJW5WNIj6yYxQjLixEPg0Xl13cSr0BTuv7cA8yAzRymAbJu
olcdgt3xrI5jBbCArkEgyaM+mNgf39iQN4CTUUvTPPxU6Dj3q9qnsQIiJVgEVeRo
ES4B6U4VLvCOv6q0BZkyHw4oNzwkOGIRP9q2EYKB79RErDySZPJxage0aChi7DGO
c9nwDYtOJt6DLYmqKqHUTQ7aCH9N1Q4QrxAFfaAhQHyhV7ykVSeGwhZYoCcTKrZd
XiPWYSmDwADPm8boHIfYQ7U700XE5MX0Hq6Oh8gT1TP0AeTK74gQl5BIX26Vwrh6
ZdkUEJHgqicP+leGpnOz/KsHALA0oEYJ0xMQh94V1DMGajITOQk9JWW2/Tdz+f9b
7fJ1vGO6xHD9wVmmCdPf1Bye0neXi7oQJnffNIKAqEC3xxgD5oUh7tn7b9CcyOF9
k8Lm/MKUpgCBTO1HKzMdj69bbdKdn0FHrw4kdZEhR0A7gnif1pRvFb2QSTSHQakc
KxXk1qvB51iGOMwsUU28xV6QFOxzw2Q14wzdBDWO8bYHUfT1pSmqdngo3IIKoouH
3Re5mA8Knwt5ztcU8G4851hCPaVEnu/fGIizImpl+mlHIjIyTUhXyQtZovIzQjJB
wNjXt8SM9M8NithTAoK7SOUW3ORKVvU8N4vfzgwpO7IGLcvIr3DMpCS2SlOGSppY
SEfd2Haype2Xhl//bioGqkY2Y7tzCXA89hgYKNQS6VxknOMca1Ms74gUT1cYiOoN
FgbxVqzNNtRN2MV93j7rYFcrkHlS5pNoGLGB5LYZv9eDzqpIU4kdIwqZaAhdeENt
3ovYc1rG9uByeGMHFK5nMYba5tfHLyDBIJztrbUH432Mgetfa4Ms5xo3b8AVcKQe
E8Hh/dK1LVyCpTeyoa8lUvbT7s5c1yXaOloQNtStCoK+1n0qr/HyrVXG5YR9dx41
BQCQ2Hk6IGiqN28f8l5rrKlqhWG/BVp7UiUG6jfhbQR0rfSqSviRuK88AF8U7Ki6
srARPOzXCAMhuJzXJX4j7qLG8//ACbBi/V51k43pov3rycQ3xsNV+rmZjQ2QpGHy
c11djconHwMFoPq7gSkHL2HKd5p+EipkjfBK+F/V8JOuIcT0J/8D0PvhtMMpNvec
7rhAoDMzeGbk5JG47X5TijNHZAXT+vnWI3M1G+iFEkWLy1umSWMKPqLfeBXhLFYg
zxLsrtkrSfLxhZ7sjez2B9fPhQJOk8lUzRQ9vzzxB03YyXpBKyjGq+wPCcah+cbF
tR7SazyADnCwrOUBEEWhxalCMkmTKpDDbuWf/JAvNqZYsHgt0po6mGEOHb3YVLeH
DqMEjwxu3JQubDLQIsBjajcQD0qARvnTyH4vjhojklXuxdNryPDAdh1Qku2mj28i
im2coevyytNMQgoLvTNU5Be7xs0Opbf8IymMadX78OWv6xn+EZUdELhPlqyLNKd+
Gx+0omwhkL07L0xOLIYFvKS/bZxSfnvUKB2nxfcfFPtjbFIP1RdMp35QS7R0ivbz
57+ot7rBhcz0IQKbBmvWFsRCgo3Qs6UJp7J0iArLMAd7TKnBWEKCXOILuk1bDHT8
mAzb1s7m9XsxpykbIKX7w0x49AjCuq/UyAX6YNNe8UGigJiPyJRxr4LYB2/hWhKw
0ozJFPJ7iXmnITX2ADibyKvq2W5LaZWBWcw0wCORsqoYFmBmc8fC8OJ3kfsXv9eC
231qS9BD6p9nAJ3eCqKdgjW3dkxT/gUeKeXoQHWYBQ6r4QS2EAessGGEp/fU14RW
X+zqIobQbJP3IMqpl/du64mnma3AWGiU1U/bOPX30KTR6zXwsBS/pg29+i1VdRUS
y50oHW5FOyp38nrKNUZcyFLETgI79DJG3k8Oeoy0Ov4fu+3pEnzhtTUH7fXQHUZ4
1Jg+7wqWfraMVZ2lyqTDqP1R/dLn9RFf4HfcDswo42hdcUd7cU1pJb5shDpFjgKT
x/xAqzgKu9g8Dad5kVRAEEB+SGGqeM7R7bXTA3Z8xgOl1qjInrj+g3dGkkJ8hAYb
MDmai8Ag5wQqZjFafOHa69FISyaJ3fmJtLwakvdSpwfPmNcqZ0f0fiezW8nNKSZY
edNfXb6HNhsNNkvrY1rBAvo+RwzJ8hwGFW/82jt7A0XgXidIVMBtNrqboJf5LpTl
YEV3aMQmwz0/G083Sb/G5ruW/q8kfoUjcJZTZrVil0khlyxQd+cz5GiUEWofuZ/H
4OhN9MvtnGqpgj3B8pfKoR36kvoHRaIGIkmn5jHK8VXUXKme4NVbaLxeEWMlL0XG
7mJ+RMYAia1YktbHOz+aXua7c5/Bdm/SE9lCSrCnFIGjy/czxnWno1NpPK+v/jpe
gGEyL40quNUF9g/QyXzCC0b8YN+BBjeN/mr9/ysrJ4zVUgjU2S9Ddn+cihX5y1Tw
Z6LOagY7lkPltx7ThaZszvNySNNl8hTH9TYYniA7S2d5jDZb35/AyQgWScfOoP+O
IFNnP+OfDWS6xcHK6mIiievtjvPqa2A1DBZzDb+6pU0zbiornS29mSoi7g9OVc72
cU21xyssJE1b+atJ9a48rD+e5h2WfVjib9qyNHxzLMMN3LWWj2tGluiFywqASlhx
ouLLLBRxPF4vD1gPsztGxoseZeJtwOYDDAxz6/2RvtgvTOYZ6tdCoHfD3WOB/sb1
Yk1MVmF64q9gTVyN/IfwYn5zJfIgNDLQxR3l+FsdRQyZ4JT/MdjYM6WnCXnsyY+R
Z17vXoqBkoPezO/CMLz0pcCzT0BVbArReblJzIABMl4AFNF4GBJlIzh9A58m0vDQ
Fs9WwZxRnwjmmqXtHj5Z0OdZqESVmR1plKVzWBZ9i0acfp7JChmnDx8oz0bI7sU1
9Jvxf3A4RLPP6VBiYwZ/ybe7yKOQvVqfXS7iAjji0nwuUcxM6O3ja9RRr6byqxyw
wqzlLnazIbg91LTHOuRnEHhO75cpl3vG7GJByIo1OvfSI8BQMWCS0sASzbfbMFHJ
mY92ZddsdMGYdClJMG7lj4yyMWd6rwCY/0hqKU7pDbmOz7Lg+pLZDqLE3yt1rG0z
ElrC3KZsvYR6tpPvdQkU8w8P5V/99DIUwJVxxX1oiMexz3gzQI0RXKUvG6K3G4+i
ail0Y/Mw+aeltOq05GlN8Xu2ZJ4Col+zVLZIWZIeTBd8VWTo0SdmUomv/OG0kUP+
nUE9Geafn1/WwjAdWokYlESAMWWXNC8wxDhuPeRpH0eH7SrrageIabJs7iBd8XEu
A9tzUuFG27EphBPvB8RfYDr11mA7dkVi5ObI1+o5xecqFGfm5rlc/vpN3e86wf0K
xeStqBn6QRPaqIlgmf791iVP4F7DG1H9sbZgLVdOxaGFeYe39jaySRJ6yxxylsCz
35QBh91xmAnsDB6muGfxLAQGET0Gle03uRtXa3DITjyS04Et4W0x8JaUE5OWP/pD
pb0mzP0Y9yj4nC7y6tBmDN/MXt6Ndn9UP1ZzZScVZgj3NbdzMcHEa5mJ8hyYCX9P
4BIciGa0EX3cPjugFCrMgfmBLSTWl8VwfF6kROrJZxDNVAy96TUtlw4oxQ704VyK
vc08CyyHZMwFve5a4UIPH3pqvR02ndmkm4mZiMO4KEq8A6wu1bd1f4Zh9KuLESJH
x6HdzEximIZI7uj13bNFf9IKgCsH8DnyjOR4aYTYqXbG5fbuyyHJvckhft+SZFa5
hz4ZyWS/F1yojyreF5K7hQYZxZuXg24YvBrxhKlz86+Kz8mHShH1flTJJj905nkk
IPdNbPKQ74ottjpZxU3FBHifAKfiT+nTi7C8AbpuIZy1YZ3yyI3YucvjzjHXv6CG
TviT42L5nhtET5/06qOh1gL4BnRstvm6QC2zF764ug1HecQs/VPTVAlckXx/zUqj
wU45JoSCo1WXLKRHmqwpZIPu14G8tX4sda8C7pe95z/IuVP666mqPa4sFQPtR7zp
w9RrpxsJyUi7QjlnE44thKNQNbdIHGeMvy/gjOqxd9OzIbXfR5lDqTLZ9RoQjvBl
AYcBAloXdmU6CzfQtEBRJekgv1nD0nhBltQ+KR3Ypb6cNKrbr+QtWXWE8dtEqrHz
CDQevFgmxdEeyMDG3W3vyl8RqRti+sfPmYNZwbWI9rpGtaBEUci06T7iVOYA1wU+
DE4oZ41HUJ9wjZTAOmD9XzOxSwTO0N/ei4rzs4TTcDAYJTyTFNDBjAsKSWOwh3Sz
OT9iVEkKQbdI/kaDXeokEcmomBWMzeogaiZXo+MvJCoWox2B+W6qfZgC3df8yNUf
YjAlRsQBNuibsoF4iMEHf4lWzQSDSFNSgZh6iBTRdX7vuIR9pGyyl2gfPk+o1pua
NDSdKJx6bnjVWe1lEfN6vnXWER7AodeCzK4/CHLWE6oSnubCl8uktLpseHReJXIO
nLSC8ujAkWo3uUdlh1hh0Qc2b72LfUtBe8M8dpfKaUqqfx3GWgaa+1QTO1EhVX6V
NNBM82Dmwuiqt6KHgh84DvQq2UNfLpGEkFUGrQSi172uNG0MJ/3eVeZXnJmrFQmC
BTTyGPZSlVrmIjNAxeCslaGIgXkl+q5vPQjjGxKcG6Y5l1/r/zv8bd3kBulB4LtB
g1fbG3ugwSFJU3+rf+gQsyRLCNnRRtM2ifiQwu4w44ZTLDDik3ynsp7+zVqL8sBt
rHUEdDxxSFE4fectsIcrFXRetzh1M/e06RuxWqxfrnejT8thg+Ws/d+y4mvQkguF
3OvQV/KZuRiKxVj9cXnjarwvAj2o8x+9o2UtrAdW8iWipp+uwHFO6PBb+bVcbp31
DML5UjVoCBEvhXzXYjOhAITNTEw0gtb3V5bRfCHMXrYx8QR+yiU+erRMkVAcHAHZ
Q0dYCnM4JQ44qJ0+2BWjw/29u6xwsTaKyCZztbamBqFJR/P/D16wIYvYvEutim00
8oPae3Dh5HoRu+qPWHOyA+9tmzhlMWsJ57BJcSunhkJPnEIqIGtBymdY4/0sgny2
RgeOZ41g60+VKTyPCTqbTEC5CWFD/NMZ76IR+NmKITbJq6WKVZfrGp2AdEquzntS
+gQ5qSqDoqKiqmVJbhMi+PA1UrlB+ynRV15XbDth/+/TDr9gHP9J4t1CHJQS/QEU
ShpvD3hXIz3Hj80NoeUNiinx1ltaJn9tDaoTQfY7aNeOkKwWypfgXzPN5SZibS+K
iTiOa72wkit4gepSw8YNVv0YOsvUF5s7wx+ugMRTwOteL+lSJLGWVQFzDFePSNxn
jrFfY12nztKyWj8pycjoXom4zdNf/92PeY0EDsdlQK0eWe/2Gbz8K3f7oXbMhZ1Y
NScWnokIyoA6DpPTBZZnP0qyy3wo/jMMq1YnYWlRYh3cOsNIaN5fia8E/LZ5M3qO
+RzoTZOZroOHrmcktyfZUH/MpCmNydcPFj8P3wAssbglRUIMgROFLjat/3+9EDIB
y72kWf4wtQmDGuZX2nrIYtWE1SaQmWHgBipdTHSxKIsXb8n3L6Zv84sQb837nPYP
3Xbgjn2f9e1MQK1pQLn6BKQcJsPRnD7e79FdT+3sxVtOrOvtNWGHqb3cbZfhVFA9
OOuhZT6YW5EI82XltD69LY+563aZImpZTdedzH/N7Y4KfDgDEZ3wNeUJjcUjkGFg
XeYVkpnfxELrcS0eKVHas69UcT7Q4Yko3dotquAGXfq6ZdRwWn+D73IENRSnsDu0
Rb3zVc4z+LQZEirAABpmZN/5HiT2nyL2mQrpjeo9AULXQ+3WhOxHEUQ27V+VF2DK
RXIifJH6dbb5dF0LalRR1HIUkYul0e/FeJQZjirVGrdveAIpTgyTNvKrnpD3KmT3
8HKe9cnFBksdTQb0Vb6KMPXJsztpnId3Br7729g5v3pmOFkfcmjIqVwuBb4vbN0K
hd6RP2Kq3adnlhBWqKs4ue6fNYPBZaEduGil6KUSf2aj3cT3KYwn0SQKjIaRFF2E
tuv2+Xb5svE+hvLc8QRx5tAYuAFG9TWWMXgXV2JO6z62NUQzvNV3SoHRcjdbG1Vy
R8XqBzDbWddv6IZRPTxZcis70G73gy4fYbQdS4/wR/VzJJ55MvSK2t7To4GBp93h
VtP75vhptSPcPrUyUxRs7K5m4QxXG+qwMlDk/PQyQ0SScNS4rPtI3nYSSpOgo4Dr
GxeRKD7R5t5nQjKXQDr/vcuwNrKKFvVlIDjEsbgCF2/vQ4jrs2f5IZeTeo/4HXTz
JHPF7fcJEOMKyOrUi2rPbhb6IUmT6bErucS1Hb9yvsiHT9pBRUiks9Lnz8bTQhgM
KtKmVMlSVPpHPHlHtX3sL/QlHelyXHlg214SdA+BagHrrygKGMSGHNC3+bxYkMKg
PQPnytoJhNBK5INQc/sTLNBBsdKNzvAtE+MOXjIYGv9da6MsYtsZ1IsA9oPgoN0a
42YG/O9uZR7h2mM4pyqGKFVKehtfN1WVUYR06jhwrZXvpSut7i+c7dWqp+bd+Ftw
rO1HrxvQFohM4zkIRedwGKjbG3cbuIaLlbw98s6NClM60nz5ep/G1XnGFE4TdpAX
xdCxyzW7bqjICMpy9AyXJC5HRvu7HyIgyXtYgEvMNr3w30eHheYTdJwox5xL9k/E
Vrp1fgvgMfSeddnAH6XzzoqkPfQ2DxLA1P/iYgm3JKUUA727ZAacEsjN9net3PGq
/43+LIsER7/QjqCaZuvlTJzGf0Lpheg8fiSzbl+04rmmWYpucUURmtatOZhpnHAY
+AH7KUm6uguxC4v3oYxlI1sFgSHjZRyXL4dBcNvU2NEBmRHAo6UjXQCpmt22Y/3l
OSJ6JYTZehMA5cRW58mfIxUPThQwqQK7lfCluBUE0UWRFzEupC22xmx7PpqXmNF+
tjvtYdAR9Iawim8DZJoWMuLtnAa4XNFfLCTrys7K1G5QPCSu7vhpERJDvdZ+zcbP
qvcBaDVd7hbGQrMiliNLKuJa7xtC1jz/8mUTIaFnNWxPzlnrf6pz2MUFd28f/UZ/
8+0yVA2KOJ+4C6il2i2VG+Qj82fWlR7SQUHBhNM19Fl5ZlRAlJIgPL1Ch5N+2YES
JVbMVitngJEqE19+ltBUxGfxjzk4llnCb6x5Oy9mcUcW4RYlJhFvOveCMMw+2+Ma
eSI5bpk9F8+fYl8Zecdon3FtOIn72FAf5seGeqCTZpbWLXl14Zfz3LLq7/68xQkT
g5KHcx0bSphqQU9fSbPMoQFsuKkIzH1d3kJsmp5jlI++D46oyGNGDfmdqv5N+23O
fyR07F1SfmTeRUtWdK1LqHpzTTiDA7L8f2cWz43q0L4A755M2+Sa3Qdtq9Tb51Yn
SiLeYQGotfpx3MSsdjfj5u89XY5+i74rylcuVctfCCA1Q/WP47FORoTMPOZvve1X
tInaDZn0KfhHzJvCYa/3cAlkF3F2ZPVg1Wz6US0m45rIcGJwWmMopSWmg1QPF949
Zh59XHCMSgjqvCrHNhSp5jtfI11cS9ZPLqCCRx0H9TDNXbiq53mrzBu6cYpqfzum
crFWtJbPw9a63ArsdmkkfP85m8Y/rhR7FeGg5TqYaXsg8FYhSam0WClIqBfIuCDM
Kjc6Ado0Wr/B7G6IT5HxroJXpD8MQScGDv5SbBKELDLa8Ik3nlSNMGtXfMdrYrCy
Z4BoX9PAf9B4n62WBMESmtZUW26NsplNroUm8L8p+uMKmlpjQkUd7/ArT55Okq3p
eXYGdKsbV9lQqNzGrhjakvjqkTvYBUHm6HiIEOzkUFhMwtj/dooCHGDpXoxgDXIY
ePxnV6mfQ3wTTTiQydWQ3CSeHLWKR3zqLL94At8I7oz7wRPJyQOUylZ3jxZmLfeC
PbnqNCES+h4/Rs5lC1UAVUoW3XOClSnY2K7aEFOqHrTefVZD3TUki0Pi/zY7V85j
UwXF3nZOGuHSrpgUS6BO8SoN5iRfiMeq11zuxVR8uWmYkOBVE6rkwGM4nMQkz2Nq
rFlwUcsZOvlNYSLpTK8G055aFXlKlUkFCwMEjlEvzmfFKeZ/YKAuT2dGwf186+/Q
LoAInJ/fcoAfxamFA4q9rLhu/qGXVm9kkWLBgSmFKeuoZupJi4ylXbck40YMZ46Z
4n7/9hQ71qQ7DslD/81d0wlfY28CRuoIgi7/4WdGNRrrIWxwY+mS+sf5js1tgeO+
CxgmNPTumUinUQjGWVkhHs9GSZFOGUJFmCEFXwSygojB8Ohu+HTWqxqOnqEX93qL
PT8PxO0JOwMqs2MHmzPq7O16Tjs/6LqEKCE0rhyXXcoEQnlrJjV83nDxE+lAhkVi
35+4zEvEPQhv2cu4yAAC6NPGagGYtQ8DPxx2PHdVouSmHolXFYX/WnVBs/RF2DOP
StqGVeu3zZQjGz5nm0nKwvbPaYc2gymzaSzN+AgKKc1RBtv7StlM4zivBwEkDwyo
1givd9UvPUtaVBfnzXvp+LCHgx3aO4POo2AiqJf5pS17bV+sPRtSp/rHNmyz3yig
e8gdsCzTJIaXs8gGUwxVN9aCmyBZc48voZ2jM6O61oIHrdL5VPsFJ7jv4gYGBNLt
Icrueo2BtBucIZsKQyamyF11EeBMqY1pjWYi09PcH3oV1fbrERU3TkorBBXB3lL7
oC4WhtU1aKCVsFfPthkokRoSVKWbwJeZEoYCnVtOdDP/WqE/bebll5WY6WHThVLL
46/MQkwNQkLhwF+Z6k781Oua6Rz+3+ONi4OgMzKuCUQGVbuXB1PX9qe2BATotoTa
0mkKnY8yLdbs8IyV3l3OgKJclrZKbU4sU8AzPYet6MLj0rnU9QF4P1Ocr8tTR3y0
YK7Pv7AyknJ8EoJ2G+9xyuw7FifiW5OfbXo8xhHeS1PF9+Sv/XGDtGMW373jYSMv
N7OttPdcJS+OkwKGIgI6asmkRuQZTRxBfdsPw3BF1yuNbBY4oyZBB3mRKWi3kIm8
25vjRILcXQArd+TIKPaA0lNwU+1cB3rSf68JusNvxLx1Esj/EamC6c2WV+5v0n6u
ZFWh99ibVX++gjvz6+n1jntcuB9TmsPI6srhp637t8gexBKKQGz7W/hTweJcv0Cl
k5HsMDgxZ1YPaVv+9/o8dbxYnHO70AajvrKi/QWnL0YOjQOFlBZo2nsJArOwXWUB
5TUyfrG5YItRwQyfhGgLbNNzlueyUWNY/9s5iA9mXI54m1CJPtOb2MttAqvzR4MG
NceW6JoRdY3c7gM7gTduvZ774Vw0S/VvYcNXSwPrDFX0QdIQUwlnDFhAnuvcGNbW
voZ9qNncc7paM0HMVVNAutquUYwssMovRLJfFUbu6auEqAr/Fn4byq27DTS2sif+
djPBbJ8Xd6RYRM0/GP3ArFQP8O92Mem2nScZgCvG5MgaJ9E5Uhau2OgJ2S7riLDX
F6Z5D+snHzXFNDpwwCI36ty13tvVstz0UZIBtQwb+cv9dJx83oQWOExsdayH7KMB
PhN8OTKzKrOzAmjO6Y5ujhmtBAsHq5DyZpOHaQ8yUKf6d62nfcLlYMdLNSKYE5wh
0lVS2aWY6Ewo3GB0EvkkR7bbyeG6krSA83o7WOcgPAKCBl0kdyGHyTULFynbHJsw
y4P1CRNPPoMs+tbmrKRJo1dF7nSrF+qvAm2Yamu5BQIvGCeIIL6cY1LnSuUi54XH
DNaCcWm1fSJjUQL/N2KvenfewA1EUE36tSylcAbftBhTxqkhXOAiRjkHvwL5uw7s
MGGFuKBYuWG8MbjUdFAeCW1to8MD4zITBxC4PM/2SXidQp/Y0Pczm/qZblA2v83G
eugMuouiyuUVTCw4v9eFw/4jCH9oqase+icGDVwz+XmjiuQ+RnBJCy73q30ugJnZ
I/C9DNW1LIgv1rubZjj/1ugUXayKDHPGgb1gujTe5czHcZCC/PvfDXjjA1LT/X/n
08IKKAgX3yDQK/i5SMhaOYpWQYcmfA3m12g31VYcfaCXUIDj8nWiRvPLod+gZhyN
YVGD/DhfV0Kj1V6QeJaDtzsaAeMoJyU/OpHaBhUMxICZNrzWFmcmHiPdLXmhWdpq
2QNVRoIDAvnwN191JMu64RhDAdoiX26VW3LjTM6a39kInmiey3YlZfEVVOXTgRd5
n8rvfBvc8X7Jzm7SI9BKoiBt1xvsPYVV85WO5wArnOPdfPvab1afDcTNCJbaMtSy
rimBxc4qN1K6CBPsypZVRhEWAEggmoObWsC1jIqJgrYeq6I2vU+9VfaZeOoAlF76
xjKE43V6m30yq2YwM667J0B0WMP0z0ul9O7XdC8jkkeNkopcpIYoIrWsvsYMhAPr
XPRDNxJooDGsQGXsjlg5BKF8NIKJQ9Okx0zvkXDKNoPSF+iKO1JQuxguiwHC+Mn8
yf5SV8VGHQ/YpVSXmUvugHZZN0WsHbPif5tdsMKUIQIPVEIO2Yb3X253ePo/wXlT
ewHRpJic9ZMXu8PU7SRzxK+Qp5kV1IKdzZZgXZ1wMmMBz0maekM+bRxstc01tiM8
0QpRnq7ned6axSrkd8kt4ZTR4pd8VAuTXjRd/I8Ximr2sZKquLanfBoqzWADjOp4
ZWGFSO3c/hxxp6/rcUnW1bsSA9/2GlmzJ7Z7+KXG2V8xBDNCjhcPB4dbky5SdD/b
hbYABu80WJqeXXSbWV0JeobgBd/1H+Vee5yT4Agtoq6FEFyenCDO31UXzkNty9c4
jL+F9p+XTkhAgztRxG9suuT9yWDxZq3n4sCyp4T70H6ktsfCRfibg1YDM3RLgpVf
aUpENKxqEH2vEXF57WP+ItEKvkDWzGUTJQ5rPGlXVaVypOSTpFZ6q9J9ERzX1uX+
oUizpairtqFjyGpZfit3nwtIuLwcI1lM86U9PHW73kHTdDbpafNCXCl/84ECbCye
RKA2ISn/silfsV6E4/eBumpLi2fw7VMLszLdsgAW+QHGpgEoRBMFOBrC4/ubSxiV
heMRLkUYYnvKv8+dWA+0rs5ZSWxadS8mIzE8kPFNIXlxuMDnE5U+agae5wRHCfkn
9u1XfvpiKMFB19LfHOQCSE29EWqflvPLdGnZT+VCFi3e3hUuibqMWp7/MEQiZNa5
nLmMsqNoxk7lXldLsuRE3MZzYJkbyKy+6li796+IRdnI2LcviAM7ht0Oq26S81+p
BpE8t3CZAxQdEF3G1Sdx+kcP0MIBdeptz9YiPAkqTqd0SFvNJFl70p2gv6KfPApv
nUG0jzyc3CYyViGv+6SG7ko2+Zq+feByOa2lRixpqYdlqz2uOi1Oxt9mACF80onM
WF1/Q2aQL2KaAcxBSPKdr62I4kcW6xBvKdn7ecAFiwd5aqFWolorslea3abdib2q
YFthtwHMFbvXZ2pZkJMmfhpT8jNV51iuZR5Ws17ZnlZh2+LzuZtyhsKgUdSiLuWy
PFO8zQ8MStwvNlNacmn1pOaX/3Tb9QmdWpDrRe5W7RrtN5bTuO2j0n/UzC+oo85R
HWFrR3fUsvi0ZMuc6aa//HPb728r3LTtv+aT8o/XZgr/vxyB48ZhR2PC3/Utlziw
GAnioWus977brSKEnKltPip8YjvzTlAsxvp+AseLO3zz3iz1uj/zTBL5uz4dYwdi
g6e7dflzPP5/y8YEdD4vWvbgLidCieZTAQI//PBJHKPO+rHKxbVTn2DU13dmOA6L
GnybjJ6AKtZ3XruPXOnoCSD5T4wm+7F5rEefrg+IkldHfB5zrlQwFx7aOnzTQO1+
jVUvctgPz91uF3IVwBlQ1euFOOJYZx5VhgxgLEKPGhX0Egirlr49VvNTXDQzwIVy
7CJ57wtdkWKr3G9YDmxGeOenS3gmsd+EN0KAnKQdiaRKw7M5in3bkhFySi4nGzND
Dl7OCdquoCD4+DeVfTUTCdBObZ3QAdM5XqqU3j/IlzgdoBmUqCiGw1by67MfS7z9
S8jQERfPItzgy8+bq/xUmfVoxvWjqzM55qTJ78/rQicEURYARup5Opod1DBETZaK
oXCuJUvyhcLHcxjlWcG+FfRv06OLdPKa0uA/Orcv8EZntI0su8LHgNxnqwK4P/VS
PE62AuWdZIdheetJsfEhyQ89cUHjjp8ZVXFVPTeyxzDJAdSY2erhxUfLfB/R6wkb
OEjWnABsJ70F4+4sgOh56yzIn3hhmxgWStatWI1S17d6N0e1OwGHh1t8W/pRdoj3
6K92Say4G5Mo3B5gWBl3/8QbkmnFHsj1BPFuUyE0vbxs/Lk2oOLDTDRJ7YKlSuQ2
lLDKWO3wo2y0pLBGp0W63TErGbKB/7lc+xEnUjS0T1aHb4lfiehX42EjZMtGZNkK
0Z5WeMNjE9ZuG/KW4F9/kMqoruhu0ACRssiztqV1f97oJzCbcxfKzg+WAr/1oi/v
BwHhMj3gtU2n2u2t+HgniP78mz53J3IpgH157RoOgacIc/O4VCddfQAW4RubNzCz
etGgCSffcXsr7pzGShGG92gGD6eJH4QxYobVjgfpPQLXs9yWbnZMQUSOyGmNMzUi
j05dkX+u/FpDK3nqR0yVp8f42Zsr0mjuy/tfjdnRZLIlZLOCtOai3qdDPAPuy81F
L6DBksyTH+Qkf+3JlRSoEPYeItLxDAywA28hNyeaUuu8cUZ9Rzp9AeV4ECXz2eQQ
sI2ImvOLAG1ALBI9G7+BKhW6LOTtJVDQxKIhTzu8Gu26T0stz64AS+vW+/hVwEJK
9EPOQEOHIrLk6gBpDbRjQ6obINUp540SCAWbitmJ8cpSV6yJjjKAop7lZdMAnaUF
HJ4jO4Nlly+Us/+NlutlXv4gd6XTyD2J/Uv8kxlBc2EqlpFYVwgRikdT51IeOOy1
ayIVNK43HOowaQSlJ9w31waMl5mOD27wEZIKmjhz83rH2n5gavZbCQZgw58W1PAe
g8mC/SFZ51zlDpGB6LI13wrbcftDD+9O2ZYNZd0QFYDbDmZ24BuAjVd38F9eyKPb
loceQgNzKdycIsrh3M7zw5Qck9ABSC6v4+jCpKjdGzDeGQtcWyx4QAc226pTrh/2
h8wTh9IfDAbFfmYzS3SL23/qT3hTJsvTsrotrRcUlJCRuLoVI0zyEhL/yxq6wSBN
8MYW4gjjnDx7/5Uj+1L0jsQb/TyDmC7Hc+W+p2kZqgLiOvlcrHJHA94P59TLKl7E
ReL7NWFYAyQ5HIqjqYACuq28mLpjanT8XRTdJFXNIxbepKxHb5Qfze8fhG4SHwuP
dnSKFIX4W0/r3xzmcn+9gE46ms7oXJ66LvyG7xZPuISwMvcLwNzm+wQ7IAUqzK9T
ofSpqWIfbxLHIuff/n6fDyxt6rKZZg5S/6tnoIhzINMZZpBZkkGfpgLTxP2PAVNw
ayZGnO12uN8cZFW80Z51vBNGQamkZ95u/DoJWQOBaSqRffSh88uxS+oGaMIQLBt8
P0UdxJrHwC3Bp1yCBkiv/Bbzfzy0ERPjQ0qrWu3o+rptVSPZqCi5bsRHzF3eV7wT
KeY3NpO+Zqmqi9lRUpubxleCUJLLNoftomvC26Ty8IT75O3vOWN1ftBJFRKGRnue
suRKczq4DYqeKJPlw6DBJpuI8/Sfiit7lcu30z8pH0id8Vf+7oj5RNOMyzXJE3TC
7NuvoffhT55nKNGndkSHr3rgkofLwpOyxcf8Er9VQ6vHFCDnqmpsU1whLXMiBwOK
y3IuA33WO/M7SGROArmW37jj/Osq1oslI0mWP65ljgB4ehWLnHKJ17EJpb1V2EVp
MmKLHBEnG6DqOnHMpMGNlF+1RaK3TITBZZGInQkelurtWYPHc0K4tQhbfLkeU5rL
JWlCLBaPGp+fVPcci7pOsg==
`protect end_protected