`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8224 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmWdo24EC1SLhDeUV9o12ewQ
ulXp2xSZ5P2RSggIKJUy/anaBVTumwtXp6e/AWaEdue29D2ch57QA2xpCpSQlLo0
6h31LqP/R9+9HNxM8zr7EWOQpDNxzl2/GIcLFvBnVq75N5Zk3MN40scI2+F/vjei
mXV7hcjGZivJmA0PcKaDAY3leMJbR7mG4eHmjtp4Rpd8c/XD/dmOKn/zqte+YtGa
Elefza1RcEb1fdKlYUPW+uevI+VCDoudiebsuHF2xPgC3P/yO76UUJLZnCUKlivK
pYXrhpFISrzb7IMyU82kc47pT3z2jHvFn4UujMjxr2OJq1sKLNV+2cWmoNsBfW0m
UQeLThCmkmSNdKouZI35I6Cml26IUHemS1tn+h5HOITpKneV1bEygz9EjMj2cLGY
bRqOL233EiLEKIHaxzNl+Ay0DnB/Mojf0O8/RgALt63Y5BLCat9NHnitEysnWufq
OyfvG80UpSpojY1nwuommYpuWczYZ+jRblZmfCSDzjw8TeS+BSMGUiN+wyWDLVoJ
CYTmoBCnQWbn4DIgKh8DkM9jdMzpxOsecZGUmV8retAGF6So3poP46bjBdHsT+9i
TZspHpgaox1Oi08m5PIw2Oc+3J/5/ElYtoN2od0saQ/201Q0CUIGuRzLS5NdNUhd
FpCkoimoh17kRfs0l9X40efu3f1Pxt8zxBNVNXBpgSIJ+qs2katqzOBg2RXhvsjZ
TkbqOtB4/K2PTWfDmBSK4Sobl9eUOwBs5d162N0uAgatZm+2vgKQrX+9lchqE4kz
PffIaMeSrJA8K+vRs23meXWYZgcaYiuk4mfmdQN41iIEXggJMKsUnSgOJpbeGHaO
ikcB6p0/gaG94XFnAJg1xdFLA3RHY/V3g5IYj9KOt9xfLh8SeyDi1Gcqrjo+to69
FZsUyPcT8gMTnfhohdZV17LdjrNdrQj6d2A1dkfRFLX86E8c1Cy/6zBZM8R18YdL
gZCGZeU0sBTuUIKUd8te5/CB0eFf0JWBBQ4M7w8UcWNgNyF7lUA4qhCf0Z94VpsQ
Gc5H8FttwVJZiOrc5rHgFVQaVKBDZty7Oby45PXealpRpEPx4AsLtqAx5v1K0Ywh
Tm8s+pI0WLg64WoFbDFy0Ez0w1pLb0rPO6hhP5rdwJXDH7VN0m4XOb+es076Sxt2
LhfzdwFssCqc3YH3QWa3+eMeYvV5EwENyTJDr9M9Ycx0JtFP3OvKI3FGOi7A5zGd
78OhXUV7CSDe40mhf41Zky+7JgyqgmkLITBbYOxPt4yHgm+vJ0M9szTFt75nHsQe
LcOKR3ul2fbJ80OzI/ohhdX5YTSsR4SaPj0zxh7KMu+ZDrStdlc9QHOdApHenCd2
lpoRtpN/LXnO1BTbPlIoX3vGbuc4dZM6/vG5PTCFzNuAlCdElhDG5uujo6PiHKPE
34qzSy6EbaVgs+NHDfTdNZ7bPVpUZamGuc5+eHABK9lGpBmBQwIRgQjdj5uXVw1N
qmrZkR+M5AQeYVNAubWnJKuiCDyjOlNJaUJLGuKTsj5UCKq24lf0OkvZkCu/C6oP
AKieRSD+5OWoECQLkKxkeHokqNwnhyh6SN0hbcqkn2X/6dDmVBgDXGBWHp+BQQ80
Zkf+SmIgDPDjd93WfDoDs2ukMlzuiJ+DhHw6x+jdKPj1v1lw9hBg8ESEnDmPd54t
JCPcO/p5kuVFYSkV9n09v65qkijqS0GLNJU1p2fO5anykbc+DL71XIDPYf9yZUCL
FszVuWNFSb0rtouAOV0rGa0C8s24cU7Rh1IIQPlYdp2f8GV5Qm84Q0yfcECSo6KJ
HjTJ5x5PIo/K0toVNcyztaJ3SMu1yK7/C4Gx3SdzMsU044ESZmxouKaQeSe0QSln
9B8OF4HsX81tvo1rWRuCww4wR/dkmoc0W92Ep1g524x3Eb6geQLpqs76eVL4uKPC
BzYx3U/kLgUf018l8sfp5R7tVL39Xy0J0NBofRSy6E6JWlPOHZfNvUEdrJUytc+R
VYBaXZ4u7GKr4Bd1RHnZV1v7j+Y2sAM6jh7gpqVFZR4hUK2qRnUxyROf8RPefSuP
NvHlqQCel0IKdjxy1MqtBV/A4WLTVcaROl1uGrPXsY4om5VjhGMt8eWwqe6IJVmo
/CJCo7sLw29w2RTmOIQeIcHv3TTTC+EuuP00Cp0wpT1GPJTmvgR2vlJG82bSjRyk
1hDOSwqYPKagzxbq5G1uHNZqf4gZ1I+iHvwTYlYBSt0QDrCfyeX1IOZtqvQsRGCS
uV1oBOrLfxQ1ajTXW9HZPMG87BILO9/mMbnLS+rft2xqPrbGsG7D/OUQFJAn7A+4
aRJIXFqJrif9a//9kjHRDiUNjoAEkGJAA3no2iOsydiF/fGA5qFbsZQyITWi3hl1
ugBd2xaytK5bxWAfuNSInX8EL2hpzVrC+qbJjzUUDiG3KpMImXe8lewoLnCkSAzJ
KClWzYgPhYdtcNatHzOyQukVCACG06/wVwEG/7B1RAuhoXfMupAPz7cSbsI4D+sp
q1FCRgb+T68RDOkFqghrtqEQWcHbkAL0JDUkBXwiiy42/QV0Mnbya6qpYkHxVU2x
nKD/KFw80+bSCGwk6oFiRwVJ33DuuoRT1CfmLfLCMiW0ofeERoMkcjWWDk38f0Et
SirP+BsLDV5ks+wFozLPhllXR9whBnkJZKU8hSAdJ32DERACbJJk6ymhvL4mHFiA
UT8heJn/8+/TvfQD/kmEV7gb5z/DFsQbsguRreI2/0kspXtRZLqdWYSqMtyHsr/b
GS8Rwfkvdk4kWNwZ/SvWUIrybbzGztFirkk9igO+vzV/vqLiQReXqHo3LvqzrBc1
zWo5pAOyMxrMYo6owitTM8HFwqBZ8nUz5eh70Tnh6oJOtdFw+FU2R8uZ+FqlET/r
dpMFsgVtaiUTpF06xyDPLi44vDmE+VmTrKQ6enGx0CvgcV1xymmMP1bP5ejzTJD9
XWtcIwfOjZTnjZO7SlAlfTQxn31h6Ofbcnyan8YW+lGl2FDFP85E2ntJUusiXRJK
cVFUXLdGbTNH6YUvDzRV0DF0YCHiZJsWMG8LL621OCv0AJTkR/bshfSFF0tp3Z6B
Bbyhmxp1qvceQ6sLHAjPQ7teET/+vJyDKfqOlTam5zQp+NJeGJSdlg01lgjh5BZh
jTbDUWBxEeSRdpaL49x1ZPeWiOLsd+yuPq8bZuK9ItUsOSD3kGu2ieOLrphplYtc
aS3nxCYVrlYmstlxNFOfSL9akfxKgkI74JceSY+HecBDdgbjjcQh4ueWeK0fHFcb
Q9yZvOFhlcQenPecj16o29joTlNRdceVMJPwYjlpJdycq8M6/Pe1LTHlRMCUumqk
OrU0a742UdfaD7RhJNzX20nn+Hrq/TguyNXEsnYXMq96r8vmH1FfYIu2P6epejev
uXjA3HyMhmNUVOm0i9vAnL8/8GkLghlWkf8cefLvQPoqZjlXjPLP67hH3qPcfAlo
DIHf1TKg5wGmmGvlDhcFEQ0AiBM8+H1KzUh2y2kCfAt3EkELib9fMN+LED3qVegA
m7agpsmpqvXoBbq7svikKAXx5ehkfhgOiETtC6QFUCz3hXPWNWYCBmtMJJKcdvS+
6PEy17lm1aBCZL5mAt7mUu+1Dir6S+WibV5Vkmc5aEFO6E0v/MGVw/ADy9OX2IJp
uQoSTuQZ/56uk3+s2YJHgmP73nXIgcCOOFIt379GI4rNEfMuVEOLcHLsj0o74kWH
Bw24vyFAI73h9KRF2E+taR0yaXFWymtj0doIvtVSxwgJglh+mk556BSQShd3EynT
nulFwekRESlUBvVbSCr1T4n5uMA0zH+a5265JlNNhbRJdE0KZSyPYks6zqFFwyr1
8IZbEBvqZNJ/XNTTeA3ChFScgEgmz5eyXwIXO1Pp38fM4RenXdEMQ3/mavSegsUi
jhQb5z9yqXseMD5ySla7fEiVtx7UZXvE7d5nQpQu2EX8hu1APFWuu4p54jnWBl95
jfMDJDGprrtrmA+NzYn8nK3LAUaqHiw8Yz+tMA79IYfIbCQctx6x7/iftkXkX1tc
ZpNUcNnJtQtW4N4fyL5Ca0TbxGMNW1PbSBO1PM0KVVywSU0soWa6IFKl/TFWv46e
HNzrskSYNb6u45sSadkHs+VSMh5SbfAIpktO0+XpxXggGV+U45xnd0O4CUeuLOFh
aq/3koRGICwOx6VCmJdC+uMzn+wFDcdcx35dunMlk7XgrnhuNvuoTUeGYXzqvXNk
y/jFYO0qPBTYvODLzpeg4n+qn1ZETuhox1RyJFRabb+vmJNhfMaxDQaUhJrfmlTF
MjGV5SitYYS4NIIPhBlBxgo3TZ/WZc0FeJrHB3Z+QveD3kxwyqmI3kpiwfPFhN/4
YE3ZypjoH+wbMshamYBZK6g2JRy6SxJpLk/ojtoYXPclHffF/UDhcCyPalj/CSeq
COIrspyO2YDi3I5kPsgJ0HST7xHGuAd1P8fe9KCEC00Y4b2vsmcvT7QJBaKSc+S5
vBO6cZaf/EDpSUnHurAVEhX3elBrSe2AALJDo2VnIXSLI6GfkKg32gDa3wYi7+ci
7FQcj43kOdlf/bBTeSJye7YVfdYJ+38/KiaKNX57bpwRB2g9U1EtiFucqlZVaPXv
bHxMZwao9Z1zH+Zk2fjuGpqYRK4+u2Fq8ViwhTzTvWVNAeD7qrEuxSqEgBUUc0y/
jt4mIcSK77oDUUx8JFlXYO8LwB7+i9dHH1Fh7R1JVIbvlJ7LDAERut7MnKm9G9l0
OeIurV2xa6pG0LN22Kup4lddTyxcR01uP7pAno1ayAI4yNuOBVXaHzbUUQYsVZY1
+a9icdmIN+onY6SyUX+QP9Z0bMq7eU2/TCNzykDfvb55SoetSOaBbl5SAmdSn+dv
sh4ZyMa0IAkjPcuzoEpQnzQq5sNUnz3IpC63qnMwBbaXDATnsnEhzKpTzX6lInKv
0GdxVsGWAfrwcKbVS9cQ3QcVGNsvTnXTQWSGbuMFDVZheiOHpwsx2K1tMDmvD+TR
fsAtJObBR2mkD54KCYDX2kr6u8CWcXgt18cJXru9U7/0PrcFSoICX2MugU9d8+z+
3UBs2iM5l0Pf64sZBplWyLRpaBLfh5Yfq14bMsEKT7WW6X9Yzy0GUVCvRwGAtnBO
7oTNPPDFuQjydMwKX6ENjzpWyA8EZTkjD/8O1VysswZgtv9Wgm9TArVLyaP0/tMg
BONw+9WUthxwOW4f2GvPx+3+Y3cSCmO3HNMCQTHLtFfjOhkf6FHNjXKYgA8T4O54
x6r0Qs8KrxN5+v3oIB37abmzKxUrfrRh34gOOCiwOFVw2gwxRg3y/ub9NG+1IU//
rVMYVzdmQoETofbnUKfIWViuqJ09pN/Lx91eAdECiywMpCq5Ke/Yjzku41DEpurX
YnepeBxoZ3zVHHs54FEfV6DjkRTaXrl5k3KLAlzvF8T3ohceOsLMvTi0I8lXMSYz
aBXY0WNQOj1knad+eXQHdrJTFmGyg2vxnwpCxXwDZ3Bbfd7KFxdjiFuIzLJ/JOZt
GF/zHFaO/cKFO3/gn3z15pTZ53q2QNEMWDbjT3TeFRgoC6bPR2A9LugJQOocCKQA
m99CfLYHJFXDhB+1XS4BC6gR+z2Ol1XW3wgUGXoA34QbQSbjGgHzL75YuA9vikYP
u+gaqggp9zQfqOFooSuFuUMBdOO34FiXWi6MJwqI28fiS4hbI9slQU2KMmAJAQsa
rUffwqmfJm7CXZZnwuzycTs+xuvAGVTwdbUI2J66gBU066L0e57kD1YvHd74q7Kw
CoYWSP32QI95Mf6buAgWLTBkZ3gJCVt7sqNoHeWOuVjG4NfnvEMD3HZzIIecf50n
j+n2M6fYNhLu4iwi0CZxZFXI6K0BicWOUYt2VCHoxDlZTGglwibroHqVm38gM1zi
PPiBOmVexvMgy4oPwTEQWJCLkR9IYXPRXphQL+itAGja0VA2VZnCdKlhcpkcRS0A
HCv6gvXxXdpVz2bXnbllNCbfA/gK0uRHAwFHa40ltAbmUMgpG3VUxLSdpMfmosi0
TvbzsKqIp5rWYMKRNYIJVc5tCZvenLyLy7CuAcKZaA0/AKDUsAkAOcj0l8cTGxL3
D5cVnNBBHXwX+C98hTtT317bshU9KwhRs7isqHXZvLzqI3xwLB6buF3bmR6YIFv5
7lIg2/clp+2on2FsNyEsNlyuz1faUmRJ1tXsQslApSZy48SwM8+PHZQnrv25fBo2
JhcvI1CInib8LJmAwbeW21F7ZpOHHR/SYBZCK6uVzY3djPmxyzZC1bKaxrRzZzLH
bfhdzGJW6GmmHiDsy5ahsmF3v/i/GInY4tPwtMRlFO3TZPPCMswf5Y7OsUrTUEb7
VTqFKymucBqi4ea6/3xa3z3NJA3PqiwxV/SwSrX0bxsvjJ23s7aUVawQFgT0hyy3
7d0ABEpdCUw1PvLrMy9LOSIUNnjSWaTdQfOlDJdnOmI742zU0pktsEul0vFJu1LG
sPbiqlwoccoA2WJJap5uVuSVejKpSz76yWNnqpYyzxBw40N2pNGGk4fDRdxAt7en
UP62tfIX3qaYMOILS0ugVJ8Be84Y2rvqY/E0G/juL4/Ul9j5FMXKWJ/Y9Xp5i6Fp
pu3gsxr+XFpzplsNXDwLLcwqb97t/bOgPTjAMaNInTJyVSFQBlbBAtR0kJyUjcFH
aJHlHxz+gctWaD+ULGl4g+cjm0YfJi3M7xVFmS3tG/isJSTS/TP2Od3ImmFncXJL
OIQZg6VnKJ0h3QFMHSpx/ttsJ4GsIxDUp2a60KuBKp8A/iR2/kpRVXrK+FItvCz2
CQcYANj1vDPlRkbvR75C0hALWZU4IuE5UqfaOrWK5R3nLXLO7JouLWXw+QhDUHiF
tpI7H3h7umPSq8YQpYxxvoIQODnG0DjpJpbY4fbcScJgXqXFMeBHtwfvdFz111YS
03wavxZ+h5PLP1e9aBdeK716lpoVexVM11QL3y3LI9q54XGObBo4vq3SJVGqQTeX
2Mr5vuQ5vc+OR/Ue3uJw3VU36ZsLzz49BJcbG3nSFsiYr9DXDLhdI/VbM98R9ey1
zu7ORTPYSNMH1maXMSLgFBSiy9oN9OIhCs4pHbHuMsJftW+6YW8nKr7f32RU5Iib
ttvySEQsfMVkYY2wWBp1kMnJGfHKJpQYW7/khqodCddg9xOvQKCX/3ZWsz1V0WNc
UDiAtuK9RTtBy6r5eox1cHOQqT+FxRJMvEHzeJsPgrEMe5X3xrqMNkcXdP6W5NVg
8wr2XZOlYRwSqU7WlaqhesE/giQfSt2gX4K6p1BXej5tDRpad1DILWyudOS7aJa8
sh28m+IPmEINkOdSxOdHMWTzzlwxU8STjNj0ow812nyUvUetzFKNKdal+dP88V+m
kn71mpHSwYb1mI2gA4hWB9/FHqRWmzAahoNfTvnhG2xRoUN0PEuNKBaA/vejdTTD
goJTKSWGWZEP83FCuMQ7YNmsVolPnRFdPZCoEOOlV4wqn31REMKIgrLnSmFChFAa
7Lo4NzSq9d5LZLy4gKVSBRLkOMCkilBBJlSOzNb1DTSC3k532ZAQDb+vXwVRLNm7
mllKhHynZBrJwNfv0pxq1YIUYB8uO+zF6pC7eXqaXl8k+ff95UDLs/vQct/q1KBO
+kURqwrW+Fblm695/ZEr7Tw/AAY3q//9w/BxoXhNTZ0jyQYsdE9oRib1EIVnFZDJ
GHQaBSfgEd1F/7a2COXZk3KsaFHXUd3ezC8o7PvMwDVM/e0NDx1rSletzKjVAZ53
/2n7KKc8mhQ9rbotwJyyZtz+KpWENf0Svbw080b/eHIP/6IRZZtu0iKLSbGrmodc
vDR77uXKMNOqSWmDDrcNRtEWt2Zsmy2Qv2YUlaG0v/a6EcBPiRujJ1Xto77/1eGu
Vf/UIgdMBNvPwNMWh2qSynMB9sNBVi7btqwFr0DN+dU8b/GZX9YtYZjDJlmqo53Z
7gBIV/J04mwKoEnCPyYT4okS6mVd9JmHWK/TYxz3B4Lo+Apxu8oMQfeIJHVVa/tz
icONNKDC6Cq0zT2A3uJ45/EJU4s7DVcWBQWhIQY1U2OamHz0WLvcoBOUjEJD53E3
X+mp+jp1Zt4eb38Tdj9zHMSvl+SHZ+RZrRqdYQcAd05cazKsLVvhjKamvzpeNByw
4MQK421sRK/kw3wEMA614Msu0BJo+XXoco8VoD50zBU9zmOyts0Ks3PxOJP+TR93
XXiUvNWuWOHz+P5pnXZgqXMB5LtDznNqIzupiWfxFtazAwsZpHdue64PwwpEC0ts
FYMWnLJcNKN1KsQq0aA+KZY/fuCHXP7jaj9u1eiPBb7zkR4w4Yh76GjrIgBRH5ON
iY3KtLg8CSISlo9fiPMBDJ4pKtCeR3xqWoAxFUbDEsKvZfYTVdGyJHuaGmbJET1/
AjEQP2oKXOE2jOAWsf3fRdS+9MCpmQaY5UrjGp3MAdMPj8GMI/YnApJnVzzdAwgB
uEnFoMSDVMRzrmEGLFIDGxdPTBKMS26fZdVkCaE3Z/NBgsuqvVZV4dS4HMBa0IA3
nY2Pz1KB1mAXJ12R+aXAO5su6rD+VyqXJRxVLGVsHs8XAAM9tw/8KeG71pVVp+rF
M8hL2OPhlYcpkZLLZ9Z6SXO6XJ9wZXLe0ZHxqqO0yer3YB6xdd+yZvmbQHsSm1XV
ClYlWohb+FvLSlFJ0Kci+aXdtp/Yns5ulfBIiyOa78uzPBrMaINDKVIeN+HYTbde
eU6bk0xYBPfOQaketbh/3ExsOFKjdltlPOPEPnS7UWJos8G30Rc4V1vU13+pRamO
RKcyjdXq+/jwIGYW1bTpyW2UA+weMHnYdNetgIZjr+h4D6zqnFMzJ/qhW6tM+H/k
9SXGno2Spg0Smj/1+POm1waPqbejcYF3rfpQeCNH140y0YNd0WqR7876MkqAAkPw
2H38kD5t3PdG6XnG/G6Wxk64slMwNZD/zM1r9/OuFF+wbD+ghuyhBB5MzJxs5TCl
TpMoplEOzvga6r8d5VvfrjKxOpgkOQIQTj6dxjXfSO/uHz3WzuRH7p294mUi6QsM
ZvILSqn1t6avA4A9yICwoxmlpvE/XaRC/KXxlqvWpnnTe1xjTuARMeivmqP9bcGX
/qxQ1lSpVJzMNiQlIbnCeQw9aRBZD3QfOhvEYcx9NXj/1PNBa72E+lSkiOBMhYRq
k7e0C4kj/6XI5dpi1XLp9mGqlSwTCe1mTltF/KyEnwjfm1ujT0RGeBEIFKYjqA1j
taQpfm7bQOl81/Tvc7TJqDaecuTJkelw6hDE1k2tHRVGtdu3eKxBMWULKf/L7vvv
kXWbRxFRmwzg5kZzSr/FWTj7HJPvSUBQ0je94g7Pos18Rw0JEbjdlkYB6fZqcKCt
2qQm0AOZF8rsKnSDRwupf4Sr4vUGv9Oum/kd8ngch3OplDxvRr7vwWjxUbLSKQLP
eBdd0cHSCPkpQRSQ7i/MwE9o/kxIz0gNcpf44A3zQYcXVAMJPpMW5hVqQ80lXcnp
9WYVWB9vGGVZd37knAVNyhF2Q0Zarl3axiENKXca9C/asOHKeKksvCyQaxBtqcGc
Zjlt5M9J2zg03V2BCFMYV8vYofuueDrJRY+w+QiDI2pnO4/8WfQf7t7B5aD3WNGY
LuSkfO2Q+plDauToUCi4UPH1yLbbNSRem+tKRA/+hmdzZAx4brHHK/zIo5QKpghB
/9RFI/y8jn6LpJHHCt+3ydsG7Wc0aqPyoBYcB3UXrNgj7NE4auLro18Qh5wdArp2
/Mt4Y4HLCYTRHZHB3LGZfHpf8W4zAheQdUObjZaiXUIA29ZxckQvYEL1mHSsqYjf
gFTEYad0M0dTLiXvRH/WcjxsH39wSwCiXKqv2RpES+LBWq4MdOu7lDH+jQJ1gY8N
t8sQp04oYQ/OH0NoK76XGArXw0uyGN3abCJWFzLaYRFVAkP9t425Pwm8KFin2HOv
mf+8UvaKbyB+OrILekAXh1xit2bihxZrXaqTeGfyZ1x0XidV4fFRWwNPlDUETOkf
8lJGvow24P9ueSs+ri1noAICneJDIzvE4nHgLEaBL0fS3WkSbkOEt9zEkb2agHY4
9rWjDNsW5okfhiQ8cqcqRJGzR0+KhcpKIUor5aNtzJ3/DDjOD63PCPDXSPOxck3b
RTw9h4WCKPy5up17kN5C/NGACCIPvdhEyVoF3Law2R5QHsNd0/2BM7hEBwdSj5q7
28YfH/dAH3zJqDwPYS4qUEUvHikXLQ7ZGRBzC5BX7Q8ii9LrD5/e6KN8FjnvxTA1
rsBGBwlKmCjxnqSiPGxszGfvwWObHKZIofh+hmCTu/0GlsIE3pgRMOWbS+xqkR7y
bE3J95c9dHD8JlINlm3Udmt9oX/R69VTV3wCB9wkfbnKlnPD5tUrqQr8nXfvTlvm
Tiflmo37iWGUwOeogwjQQB37d4UsEuPAtBfzyJNpRsEMPF4plzW4Cjr1M91IE7nT
wzT75YlqPcqhqxKq0PCJifH6OOEQMsTPTsO1hH3b+iXZtNHEO/YOTwGahzmH1zdq
TsdiwPMmkWFmquC9eDmc0AAljkOv2+RDgj0kg1dS8QLIweGYCxkRaCD4IUJfYCZz
hxivWxlcnSaMzGKjHPw50QFUHSa+OTZ2L38BEwZKC4+rsNSzwSe77hpTobiWUQj2
7AWHeha7oCu5IgrgXWvGQ6RGqhWUPqVNOH3uMnFUVIJL2SeF9z17H2/mpbGRLa+g
UlzG0Odlwc2LAad8Jtdm0RytDfSnZGpjaFdnGR3v6kPuRIApCmfCggn9IcfjwlIF
hLwE11kcIhKwWPuJwRE0PRpzDTmJ3P0jdFguibzsuPgQ6JobYsDlKkzNhFOhu+AY
tRt5f4N16mhHV6jTv8ihiA==
`protect end_protected