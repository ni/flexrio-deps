`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
YATj3kULTF7Ty4ORuRfFpnT6YIk4rUPRrM74bVTnc4GjdV8oSnW5PtQkMCLOi558
1V+/wvDfc3y0Z8//ksX8sZm3JZWtrxUppw8c14g9Y7owiwp+JumRtO1zuk5xFbe3
0MMnIxxoTKLhyRJtAxElG8sbx8N21OWDGiOk0Xyd5CqAmk9dcOIbxzMjW/wndBXi
maijUdqS+5KiRCM9+Gsp6k/iEAa2LnYTt4WtjkmDD1P5jZKsiMgFck8WOqLymplZ
ml3TTfn1UlLNm/+zD3SFGP0kABAiUT8NK2xBPQ5UzQ6sMFPd/np8iUZ5u4QLTWOZ
hTrU9OSX7lOvRUo8pJ9vPg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="BzW6NOo8eyBw+CxsNNo4wIDxODIsVe0ft0K5tGuSUZw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
DhjJh9S2BY18dG77XPz3hsiSQ73+w0XqfJhD+f+lIDHHVjOB7CfC8ieNRTexgzn1
5W+qoqOEwenoVQtit9u3XViXJSRJ0wfUC5a9axblRNyD2mUbyfH9+f59nWqGkVOh
ieHxkA/DPprM70F3APxk51m7/gNSLICSvbONgLGndWc=
`protect rights_digest_method = "sha256"
`protect end_toolblock="L7NTNW/5Dqy+2kJZXKczEa3js87UJ8H00YWI+92sDHA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2016 )
`protect data_block
6eHODtGLmq6ccbB074dgNWpdzW45i5jL0Nzx5wwM+RA0eeOHXxEV143NNyQGmZjT
bzHAi/6AyRCB4X9z0c4MjyrZE8GF4crbMH4T59xFHqVrQ4zXCea5w0kG5yvHgpKo
Er4+TXTXa9FsGlVtYMafKWlezaPJiKjNSxK/rgJjJFNxyrgkpayBuVX15mb3I+fO
8yJ0rX8/PS8nbU0V2J6HP6RDy9KaIyP9848Aq2kN+2H2MAajVDVJ0UXBxxaA3BL8
7jMkBfb3bFWzaRXb1Qw1EHV3NtMNs25jLeBpeFtxVOF2vIgK/jkuaCMM7S3vE3Fj
0x7ZReOdr4zvQbXRxepmRw1uzORVK83iSQWu11Bd45hvelR+05h2+5oAtPVKbE5U
w3Eq6EgP8T4eR9SapBsIvdEkV9LVctRpzJyfGioDjXG6pty8mX8gV3FysLyaTY5Q
bEXd20H556SkPYPgftxzYvSG/BVskdVM3Z7IbBj9BbVKbKIlMJ53TOEaDI3STFM8
0FHrOEPq31Jjaa38EkfHfBSHs488/86Ga/AgPENQcunqMdWKwBavpS0XReU7Gsi0
XUu0a3iCJE4lXmj83jhFG2d6w5HHQcNpG3KmUXzUNnu14qb2H0YEZDWZHqxScBJO
3N0Jl4rLUhtB/X7XPsMLtS6XX1AmpI2QdsPjLS7UljEOs0w+8521oHGilUuAL98U
O71O3BTinhiSi08yXdQVRcaHiYQrGlowgMFOTT9nq3us2OUeZg92f0uGaDhmkNqd
0jiNYcg4gaO3SCGWHEVf/2FXlUikDs5YPoBfxvo1FQHskw8BlGQE6x8Qzm8036/M
HB6bpVE8kQK6LrzO7Cw7iGenq2kSRtLiFJYRB6I9G+VZnPd7PTIO8eKeQVK2+HmG
aPPYqeyHTd0ZtPZbIankLwy/k3nLvc/QsIAcFyvaGLemN+bWVuN3I289p/VfC9IQ
aiOxcsMrEXDJTuxnBvrboLKGupzv8ROZzUKf3DTRBIZ7u0xl5Lt2P0LOpuw7rwz7
XndbEorQuJ55uei1UOcWEQxWlGw8VXArSf4G6w7D2j/zyMOp2QfC7XxDNj0hwKgE
2gWI9UgV52khGGPdq+kaCM2VssSdUkf0Gak1bNc+gYjKYQ5coY4nHIkAd0zPzh1Z
bVaGNzMMtqRMcvAviR0AptX3ngU2QK7JzygVXhW+QmiaIe9KZdgm5ijp07OTkSOv
RY8+r6EbhUWmizukVDNichhYxaOJr/4gY2iNhUa/h8B3Z2/qp4f5XeW27zYtY1KD
xeE/NQ70T0H4V3etX4IOSm6VqSVQuLtvynUoQKyn1Yuo+XMZRUIfgLecxPflMYem
QaR5PuHKpR30BEdz66H6z24HLqfw2wd08PmW22rVrDSflbF6cnqGk39XTYnaAF3e
xeoEsNDa++AtDDqp8YhU3gquolf+ykl6k31dr8M+7fC2B3LXoSRWfZW2X6cDi9Md
pDGd0WvcbSLo4d63ibi8aO77hZkXkFS+y1a/EPYxJxBT68eAZHiHZRUa0ospUK9k
NpAtDwd4Fnkdy2tKa09Ihx/bEDy6mgUT3vkdfjCJug0SDUAD703Uym9EPtTavwDE
MCApHxBKah38ZnbWpK2aESO4lpYgJF0HtMUzr6LXSNVohe7HXg5D8Hs6TeQbv8cx
agfGcmTuy1miaSgD0UTY1vQ/de+sHpvitpmPHxVdtBdx3v5qFxpXEZ3/iv9L/Ifh
8xterAsC0M9ZLmP2VT0TtycgZpMW5Bwv37HH4PWdqelznClERzpIUJfZ85wfaqw5
uX9sY0eX93NMObGd08gtz9AXeD+wVCHiR2f/CwKLXmYtOhVcOITHuYEO6iiGP1pM
XNC9blFlLxZuOlUEzKoHu07hJ8LfZ0YMZm6/D2+JJo+Zj0J/vHu2WH1ZpD+aOmpA
OHdgmFqVS4C2bAqQKUr1dI7hbNPreqvP+TR++1ojHv8tfBN2NwZuhoQN8YRUYi7W
tHbbbK0yz4m3z+uLkTinxJ7R/6IHR0m9EdTEZPr1AeTWxL1J49YqEQp0TUo2u+Ld
cNLRbQNO/JgyuO1B0oumvCnh/Ox+UVlZNXeTR67kfEnWB3y7So4wDkWMxNJ6H/hi
SuGw31ludfobJGdwdr58VDmmCId9yWUourKOYWCI2bR3fTrGZpwbra++0Wen0+mJ
0QE0otTk37BKfRW2qPsWxv5GGCm2C0RJNglzmFz1WUqntBy2nW0D+34OO9VDItC3
jO7lFq9FXQzr32/vX9h8pL432DCuL+vKw3BufKXemA70E/J949ON1q/pdRlhzKxF
wUUFKKKgAALmH3tQCVxNZs96NLxdGvYveqPWNbijpQmr4u5b4drpMIW7B/2pTTvd
XVNC55QZ9T/X9sEZeZwtYgR5T2SR2uLuqRF1Lfh86f9vh8EiFQHKbukPaczTfhk7
qHrGER3p0qw3bT4CzwsIQcfoSKTIToFQBtpeDu96aAZUW7y/aa2vm8s5ganZVJsm
UMm0Vh4l9KjKwcurU3AluJru1qQHzFyNikHdxLQi38258zQKcPtzDWakEKhb6EJN
oOKsL9UtTeHP3ffS1liD10STFKnlr3a/8RbNHxW76kplgN1tF+dQUm0QUJ/ANO8Y
cLYIPWZn7wWX4KMl/Ebi1yv5jUiWaHhuj1oFIG6Dw/i037pkschVjTB8gKP7s+CA
`protect end_protected