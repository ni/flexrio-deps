`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 20704 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRpcw2zQDHRgJxPf7yaQH79Jh+lbSMPSgWiyFCIIbh1HX
oxXmb4+fmKwVpWUCniqtORFMLEcNWaXZNx1gum7bnmIQxU7wGXurVry7RP4TBo1r
FZxg4hu5TNZgXlWDiIDnbN14D5YhYqp1tU2vg2eKqoJeNACBm2UBkN1IIbV5vBOS
9cft7ZLhnWVnrQBqst+tPWuoxI+NbCvTDt01LRFd/35xg5+PXJgY692wCa0gJgU6
CqQAy3KeWDtJz2zBR390KoLcC2c4s4Z5Ttn5HxKhCRmck2OHOq9S+FU4qM0Ywvfn
5wD+9G4xyE/eLDgvN2UFK08GgrXaBZVqExZHsIJ5Uq7X7bm1BK6h2TKyDL7Ri1Ke
RKg2Bq+NXubl51kPxGUQ0Taw9ZJlUCr6iuQ9ilE6TsmCzmaHyoefuzy9GykS2Bto
55+XruXnW1C2XhNnmWkS/go7WtXEVdOhNPLF5B48ytKXq/VzFW2r4drMwIcNej5W
OOBcYVIZsKUMZTrFuA/jf32rjrwOHACj3JUKX8eWMmFR8TbjvTp3URyKXwL7h0Y4
negg5lYpIhW40BMQwh9V3y25E/mg27L90HA+BQt6T11Xi3stc0HPkfTDD2G5a+pa
ury8YxWyusHVljzfTUXGQ8759IE9vUB0iF0XoWe61aIPwuLrCfkNctSzBbcmOD2g
f01/EY0vKXteRpI1DCAb94T0UApaAoyoxuv/RsrQA+FPo90WwJPgutqDSHCwjyjv
I8gr9CkbacHIEOc1E6APrOQbE7s7Y/z61ixcudUh2cNFndqYMxR4w9JvGS+cHGvm
GGcbp4yVJCarYr2a68siHnFwSsnOoboxDtBbcR4nNSacvdvTmGalp+dGEoOh6FUw
+0xZmAI3ZMydRsZ8NH/jIrXHMqWfCAYrWvjmVXvhsQSbSgsuQk2rHql/AXg+ISvS
nDLraH2pHuOs16Ny0I6cz17mYgL4ET43eK53cJF+eZsRdJxZTBfROhReCUgcqdjR
QJOoNHCW7Kaa9b9hLumn0TeA+cmZ+7+HGd6+HrMQaYxQ53G5ABB0zYL4ZNfJu3yQ
cy6TqPCYkp5dMOXWXPsoQ18v1oB/rj9rCeeLD8fbEqUyMcoVX6c5AgMsXHsY+SKz
5ktdgn0nfTz6B9eCV4VbmNJl6k5yH1H11Y8afyNkifpog1XrbODhAbPnQz/2jb5Q
+MjZG9j++G0e9CLe2O/eQP7b4ORBpORW+F03XNvN1fBw4fKbnda3FQvqOCEHaa67
atGRVpWLs2KLGEYaSAduRmKvWCvATYS3HBFiTsnEwIYDZMXZB2QsDXv+UKop7YdY
UoGmTDumqCz8b6qMP1XmyfkbxUuAuyW3bd88Nexez05Ktb3lzxZyXjqqS4l/MuIE
H0ITT5yTATnnV7AaEfiCI43+UhoD0AHD2ut470aFq/SDyhVE0pzeGhiIfPOkS5Yk
nHelVbtGPUWLJLT5VC3mpPRkl2f/6rli6PE9JAcyvK/zRnFkhsaTM9ZdBX5BticT
yyTFLTaGCNnSTmfp9o5LPPKGhK4r4a/LCyAY9/3GuGVibJtXPmocyfW6QtzJ/cO1
RVjeMDtCuNj03VE93yjSzb1ysvHTRniPZQBqkFIDag+kzZmX6jQYQnEkGOc8kqH4
McwRUnnVjcAp0AOysI3vnvO+7p3cSRTVyxv7baZLUmHHGtD4Qk82WKziE/C9ULmb
9JWAWq0DrTqK4pOfHQH1rH3/+roP3wNwie72+nuNRvGeSj1vjcgyhTf8DuYm23ce
RCFvw136MOPsVBoUE9/sTchHC2Zgc4aj+jXzWxe+AZicsQypvKkDSAcl6iywuPCw
0xrYKWOCgOHxBM9GNgZU32q2U/3kU7h7SsfSg0eiT/ZN7if/RHm5zZll069+NFpp
Qt+O0hNcE+fcvtB3tgok2SaM3snQguai+WspegE470D593T72YFXNHl7tTX7mwmj
a+YuAhfQrTnvMNDyVaRbYYtR3n9P4j0OZxDS2qsJSYYkg3Nc6FwLUuupuP8mNHj/
mXjyAsnFBRWIccDQ6aQ2ss7TqL+JXtpBtBCf6fzHFpNRfottxCndTGb3KUGXGCv8
LwzSyCcnOPmP+vEd06/qwEuX825U1ndpe7FmENob1/LIaAtTzQr6/FoR9cP/81pt
MIxGpu7z3qleQsumsFZfio1gUWHMVt0PUAxnQUMQBiiVYFNqrTjRNSQA0gWkP3vn
0az4XGCpe4GwO4aORgcaAcVIS2QxpEdyBoySu8MkRR/rfaD+8bdFGzeRXE7OMZUy
CQkQfR8nqm9x/AXFmRDsIcE8UcU9OrAeaRPTPvPl+Zf7EPDiIhmu66lAx24gv74X
rEgyStkHBV9Ly2ff8GNAYtufGpBbfUcG9V5p3W/l0EYmSVuQ+5cbIsViaZwb9AAS
ofHK5Q2Sqfgpt91s5w89o5XlHZgdADg2E7kt8nlUnP82Vd+QDv0NwPeDvy5xgiZh
6RlWPXcjrFJkXiD9hDAQaipeUie3QMMlIenc5rJR08p15iE0MtPo+ctBLcP1zVWm
koU07nWGUvisMCWZpMuTn1LTrDYASG85PmbvRnCR2PdI1SQlDH7GF43uA0pfrTRY
MPadHAEEsxjZ+0vQtmkyGWZAc7FeNQJPNkwCvFZZ5lkBWmdhSQ+dn6laYN3aYREc
eRZ+3LaMM0uJOluKYbrg46kSSxIaY6byJW6CuU2yQGxZsQps/yPrQNGcdzN/bejO
pY6J6/yIhSYB1KJI0yIZp1sgsRtVv93mhzJzGQhkgOdbOayxRjzfl876kMbUuCo9
qDDaAesI3S69i4HgPeM3TKBM710ncGY1XIAUPz8Evlru19s8Krm5L0Ofr/MFZ7wS
CIAwZJ/WhTsqGzoG2zykeMp1/ehHI3Td7j6IGaEs22+ncHycO05glN7Yh7jfRaA4
BfK1UfoOlU2KGTBAoPayI3gT0MSNdDE9DcuOwYWp0DEZScv0No1W3EP7HL0ztCt6
oNjnun2gWE8YvMx9ZZ0IMRe+27OhhgSxxNvgG7PEwKEs7eqPBC9UJXMCaxM1BoWD
WIjVzPyGk/hw+czjwQqL0hYm1PcGP1LgjNr8/OrkDT/vnuYg5TqvQoc3Ge0wysGU
wt/6E4WLUrv8mueMXGB698/cwZrOABoIKMrtBWlg6Y3sXxCsQLikbEfQOnHdP5gk
QgS0fHH/Fk1V73/V96XrdTcfpYBzyfVInl4cOOaDMOa2IHb+GrnLkwmeTucMOfnj
P4yGFWefZ7Ifff6OZ+NW2rnRFouvKtcpRGs8ejVY+29Mbki1BVHDqQZ2QaMS17DA
jb9tPJAorSYi+z09TE9OqAB4kuzQuqJQxNENT9pd0MvVI8oLWt+d8p/hVryLmuL9
0RfKigV5qwNVqyUyP98gD4t/N7Uq8ghByitkodEcjqjtKvzde6SP+KFPvkPs2meC
55WenU/eVgO0Txq4qScOC5wvkrSYg3Exe8A13EQce+SQimrJwkIO9FVQQqrKayVz
Rp21S/hAGQQs3CIUORZhLj6B5Ols2cguHyRT5TACz19jcFsn4WP884+z26x0yPCk
mNwxabq0jcx5goiBzBY0JQAhrcUKAUL8mZXV+ySzou5Rz9GoP6pdnlQkozL0RsYu
mx3o4PGy/9ktSw4dtVtYl76iuEbMIq3Gf09TJ6kodNiCfmXI+5Kve0T9WwW2fCVz
sgsUUid8x/5RjlMkgtQu/srn8otUWuBT88lgs3KO4ACCd2rc8k1cBHpLxHUGS3xP
2RBr+s3QjFSbIlfSoGzwpQAl+qugWsM5P2Z0y2DwzENhAYkapeygNysus4nDjot3
vHdWNRajvtP9GnuEEoZpAebsxf8IaQDPkdSDV90K5BWYcD2sTjNl6ca6Qqh5Z93J
T/6zDnr+Q2BRsvtOrpcnDczCezHlZoZ6qgDo4x4Wny1fj4ykazo8AjZllT1vz4+W
vV2MGDxsMultv4JTMgN/ZP5ub+75rlrtLb0Q3chtn6VlFvqRQmMhrwTSXkl77X3X
Z3ciSQHKC/FDqkqFn9/niGMZm+WgEqAZkKPMbhh8wKyKa3oK7bg+o6BuDBZ2bWfr
IrcrInKUS4t298so9QQ7M2XtlJqECsjoBjBvKLcRCkKyTOG6Exsax5Wd9g7/2IY2
UoA4K2zU2JUQzoTZ3/tWjYff+z2nMOD1IMZfhjD1O9AKZg/X3UXxHxlU62x9D82V
Zxz4j+rXZJI/b7+jiGwyy880tdHBG2GtcOjeuy4jNTKeI8tlLgUAIL9XI8FsgMSp
jBXnk5u+Akmaj9KRR7/puiNQLDUscUf7+2ccU2G3WKgSykA7MSBG2b152ojdaR8t
0nLtCaibFbpz1qGwo84PT84Z/eL3ro4dwfQreNPsSWvNgs2QkbjLetZPZs8GBtfl
5yv0W/E4z71HzGR/VzXpPAfR1a9fCZMdPfu2NU1l8MphAbWZy7Ilm7gwt1mrL2pv
+1bQwJYRtDjYumArrCkCPYEJMCWAr01G2itOtsFqUQ9qLK+7mDj7/+v52ZfEvyEZ
8wXkmF4+bZtJK+0w6gUnZHprqYkgBhj3ZcMp+6wPCo9TsManGg8ElBqIbVC+qW80
gFArD/OvhLszuuzvMHIqC3cCJZhXrmpbapdGjCiJ0QDM+k/j+fj5Tj09cc40K358
cnp+WjVWMlOTV/pXdcqw00xZJuHbQ8y5EKqQBJSBK3DMLxc9nkBT3wOAFxUmkTu5
ZJM0oRZvY2dbiYVjNv8Pq5z1SHfL0/tYXzS8zO2Bq51uyjs6zeuTfTeHiy6u9N4w
AORi5wkFwssj6Den9dlaG6c8cxJsGklmRZo7tpDawMENrPXWxzdamI4uhboDiS5c
zOH0SOT7IXUCPuS9+mh2xhWS/9+t3NuE6xavFzoUYFiKccRvRYseOBYjF2q13kR0
xeNkPr3qoHX8fTLNwtu4b8/pywcUT1QA5OVhXrLwwLMxXgk4hOMe7r62Ue8yjHSK
QqHcjWxfrrAw05ke2ChmrziwF6rQa/M88gzIyOF8QHR60iR+VDOWUUjxjxM5nvMp
Fw6nYePg++25hE1HZLXCl8fSpyJasdNqVNBloCTvfBp5yCu7H3OaJC3z4n0yMA1R
SMHF10Y78z6zrUvpl+spvDt+WZ4F2tnZQapInIRv3fdrBZtOiBKeyBgaTVz5SD8X
hHjXfJMbGU0NacGACvYsJ72n+nsP0B0iMidJ2v5po2EfS2gxE9B3BUVLGY6ziCOT
oB8kdsWqLJnLfhyHBzyJToiVPfxSMe3whfTQptbWat1cy/+a3ptrJ18ONzH1wCZT
3IxnEWDUdp59MBP9pWw1w3CP63rbFdt2ra7UBTZuzfRm7t3VvTJOk8dTvwFgIqnR
pP9oXxJP/rGHzyyUxBA0StIG1YOPEH965ro0HT2CbNlciDUqpxMWxBDW71nq92Ri
zUFfjE1t0yCTCWiFxYPNn33yAyLxGIT1celvMy864RmSLa35jeGvcjWY6+sxBPCQ
1CVKyMIKZiNT4QcYDYs6FXS6rBwW69flWGC+3iRFKirYm+PLE4FFmIicA68cXSeF
r27VhMMA/TGpc6kkRj0CvyuSGinkRcKys+utoEy1Gl1PHDroo1F0I6PmEIYmc9U7
Styilj6uFgaph/Yi3t1DrCF+y1ntxSYBlOYk2lzhECpmekpPRdXhoslPTjFvcCYM
33XIPwDUYHLMoZOSw56337zKZpCq3fmUNXc2sh0O4oumgmxgk5OIIeC5RzHRihF1
2F1cx0UbJsAPxuQNr2KJSFghjsjkrWbgQfuIB+lHraE0vnrRYtMvx0dEhkyU2vZ+
pmrGvqtokpmTpWS0ssdyUv0bBnZwaGv4q40XewjGXsXiIPnuOGxYiS7qmf4IVDgt
0StAWNnZdtfXNjR8vu3JPweqM9KI/mOuaL4MgRnkhiNrjfj2SOBx/5iFfe7eqEWx
DzDI8e0ZdMQthFklEwYTJDBWYnnGrajQv2M8OHXmdRQ8N6tRXyOjbvJi3qmDCwMm
I/vbWmaJ5T4pZXkrpbJL6QMXM6lsRRr99xVjZOxo+V1Srh5PrZwDDF7rANP+AH6n
uBgYIVG/QYBNsgFsZVwhrWtbhLcDcPqTuH23o3fVsi3BIKWJ3XajBE6+R+9XOf/2
eD+isvhwnOMK5JFf92BrIPblspzOLtYzw9y0o+9SzXmJUFCWFZKcg59WpfPWgOiz
Mu+HlNEHpB87UiPSG8Twf5ypx8eSdkkrkM0rQSye2YHPErSTf4sCkie9M05x3WQV
26bi1WuIdL5Kdqp8c8yRVgpi3QNiG5Vj6zufS45/vyindWglGNHCbwu10rno8ADY
57brU5Zb8uZdId2Ind5uBqncYL9MnMIwoRBFBC4ttbnTBXtrP3Vfj4y34RQWI13+
vdVPPNAAvIEj4Wm6VtwNU0eyu4pXXKPHPM7qTqbMUqdT11duMLkU/RgNSIqKey4t
H/Vg2da3nFp6XsN/DPQTqX6DuwR441Ra3a0OcvmgFwWHgPPiBPfySvFvm9vAqRmo
BiBGJvCbl0c6HNs1YS/Cw1M4aYyajFqsLb1RXf59BL74EWS3NZqLIs1uOXaKkXqy
V0Pv72ILoyesbqhxV4r0aWJXLUcqEeg3FNzcT2noepIYaG45/8VLPabHoN81W8+I
tvm4wkAbRvAsYgKjjsQFlNJCLRvI+Mb9X217qmv7Wjwm9tXI8V6m10ZQScxs7Y5c
BG26iMAzPbe6dKtemGMw6NIh79Tirx6gTTimzqQnEwv3bo8zZsQ5GNlge6aVre9V
+KVAV0d8Fyse0bjYcu6EGsZIUQkJG/QpwFLtgfGR3RqUBRuBM658DHgxrEG1cZ+S
35mygsu7RfaV3WxM73nt7pZIH8YYGXdQLzR5gh/erK6Dw509fFBbuVTryxPGXR3n
M4XfXwt1Rn9tRWea7CXMImmmjOJ2+Y5WcO8mmTAGnca35AMeSmXqo5yCb/aFSpri
xVHe1+oNB3rjtXknEniJCSghShMREVnD4W58JNCr1idRv5pWglnI5Lk9wFGml+Lr
s6kJGoE5Lq2YPzTo7lzcOQ5jUXMAayvXdGG2kbtK54G2NGi0/k5U7KbDgxjvAdxd
UgX3J+G95TX2XsjLqXSeHzUlCTxG6yBRxuXm39r1zHfwwEraiWeXP5PjX6v+N/An
ehKd2LPijTRw+1716giaFiIPdkJisP5OR33i0MjSdstokN6r1d56eD2w3F/4fd5r
IwsWZTb4LCB5xtCy/lf1YPqb/aVbyVzydvJ34UIFw8JSv1yBdBQgydc16mtVn2Eh
C91Y8PmQ/FReCIDbIx3ykNxoVNRXvpvGbj3Bwcjqs5JXvYFG56ckdMbcbBVldW3/
S80x6MPSVJScY+hEJwwOyep41ZpQQLizycI1plxxF/fCzpLmxPdmHVv2FM0n+IxQ
MRiKWdmYHZ6gVMc0OSuHzkR6Y09T+QS+KusqaLAs9o7L0Uw/bTmECy2Fhq+wB8JH
q7wfpUrT9uMaOwWikkHo1GGvjcJWBItQ4kAiet0G43rtAtbot+MXGnje6/AsYJks
ZVpOULk3qMmxzvQYRGdnw20Ng76Ln+rr+L+eeInwcD98UxZod4V64ncb4EzHKkSf
3k9k9Dq57bFB2f9/ktnrjr3s/WwB1XbKzg5Ia/HyomKad9m6rcACnx73f9gLAajq
ZmdKjUJ51up7ciXZQAweTNJxDTXs+AtrnL7MyZ4pK3pZk6gMp/QYBtEgOzFlB3Fa
VhU+cVYtM0jMeOd9U3bnJXcMGeTqBdJKvTnRdTaC8DCO9nKESWDD3E5gUFLlUIHi
bR5KFhDEs2aKpTrGUiE+wVSMyFJRTiAsXDIHEGvHASwgu/+wgywdilHiDL5PYP0V
W/QQ1+HBO62GKU4sShlAcTkQOraezBFQQM7aaAXHiwPlxmNYNj+7gyX9vt4AyASI
sRtD15qi3tKHkE8CCefUrxvZ6dpy8Nzib6ZCU6tQ3k4TVTaiqvFodevqBm3OEyj7
v2n4xhs7UGk0WFd1RaG1P12+FOnpm0cJJhYizNvNInZK4m41oV3DU0ya/oXR8X9W
FoLhKRyPCOzU9fUssUGPOq+h8sPuF3u7Npp84IaNjw0jyPyBe/n7SOkO7g0zQVwa
sbgSdwPTU67b7/81hr7jyfSzVTsQaCoh/XRAWcl2lhqF5P8/lRm7ltQRyqRPLWqP
vIj5Gs/EiyqAYR+E1Qcn5KfbnLFMDiRQkjEbUkrKrmKK7+9iGTnqLmZXV/LXT//l
ZNi10tC1poozcKdHeVgWvYawP4qcQ9Ohz50YxYBuVRS5MUY9xqUEPV4Usf73Kj0O
OfeYjtlltCYYgBNeugkzt7NNagKNpJMsFl8qFvvIeP7qhfewwBbJYlUap3Rr4lU2
NPODPnqsRFtPZOOM3joC1Vew/UY60PknCfcYUBMfWhoDsRg0NHWgd48FNK2wp79u
3QlLt5hDAo8vMPtYsDtydPYDplBQtEJg65RpBHREMXNC2tsFzJGTJtAHcgBf7D1C
IooPUqstvlKJPiGITq6rY+Ipm45vRLnEUm8Ifn3FRbkzd/Dxnlrj8Ccu4Vh9rpzh
CCQl4W8QKAuIMSaJyYBQQ5yn5ppFISdkOZ3yGaHaLXXcBJjL7HLEgpbncOczDp6V
+5J/dy29hVFHCxP35z+M20e3OMNNDcB1VIy+MvSRven1EkVA+lCUG7ZAPNfAfIZi
7pkOversBqJvQ5qHzgDqfD3UOWDAJvfzLy/F9tLBetCacfIVMYHBj9C/j7bnF0R1
1DGoD7jQyGKiMAb8mXofcUZ0HhTnLJ1+UFdXM+YK9gGBp0Sx+WViCFSGa/U0C1Rn
Al1g/W6rmPlHA6Aac5CdN1CMHY9W58E2SAb4Eu6/WIYcEAXdonwkrkTkabRSNb8k
JeOFOmY+PFGw9vUPHKnuzFtV6FU4V6+qKZYXrJmToRnLpjYtFJFK6FUcJmjdrzim
l0bs7JqST+5SjtPsfSStXnvKvg+9YA9DrBar6mIN7ShHkRNqJFPh9bmLnhC6TLsg
ypGtzeapiwBicC+V1rw2fxsVE7qFD0hdwrPTvwJkt360VtLFrE8SPDRHP3OhTvR5
y5b4NluGvtebAzeJd7E1EqeqvUWghbJplmxd/Yap6ATWGd3zOGF9qc6LJ7SDgoZQ
E83hX031PbjmyUquHFLz4Xn/lwJysiJyq+0hAMnepsIZjZZx9lvsPDDMwMAFp0tV
Mz6X+xY0dL4KqKkmEC8pUt4jxZb4fkkVDwWDwzdTsLBEqf4Rnqxav5WPvZ9Ea7H3
5p7CEIEx1Jy3ot1gAAb/OYOiW0Q+XFFJT1Iq88nkwW3STUWXSNISCarisH0alwkg
YDIExodfdg5bU0UYhxOOkXCaOWzzN0glo429LD9mVL6gQKDC+THT249JyJ6bKWVh
IUZQciAqzE9fhYvmoG4dVZTcOCtakGeCE9hhaD42axF3SIdnh+3epVNCZeTO1ywp
RjmMlytuFhw7aC+4NNCEFeHXPE+Z2q268PBFbqQm9d0f9SrF6xRH/8+VgIbOvrZC
xll2kDGrkNwqKUY4ViHbEb84yFgOwWoYoevPO6yk6ECB1Spx4vsIn4rzQG/5TmoJ
XtwhTl/DEQBWXupgSO7OHu2UsAqk1DFIh3OXTDW4SAbIcbH5HkzDhVNlFfxum0vI
vFT2sY07As5n2qDWc9rGbK17PciRXNKYz/TIONehO2SluQqCQZlV9ISJ1MR7DHjp
kI4go9LxWRlhnUHmHvueil0GMc8VfdmF2ylXnb0YQ8kStn2Ojnigl16Bct1VEP0O
8+KxOHK8wRY9KdmrIJEbL9t/GKoSUjg9mkahOi5F/y7hCI4YaVTIkN534TpV5Fzc
b8ApYdJieeSxsS5jfVl8MiKYBVQS/j6IC6ZY9ZIE5SxkrbwDlKgz0XlsGiXt0GZ7
Sju8Rov5KsqoyuYWDKZ+ujB1Hohijns/JTmAW+UzLRNhQWWNv/wEhs6LBfKW8pTY
qsVuGrbFu709n5arfvJbnFq4sNKi0yRKWAVN1vxP2NvunjTNMGfLzV2/5ApmV9vg
MtvKl5tDTdHr0IVv555QuTs4bEySzYMqb/ZwlmcEVfwulvBAmkGztDDjVH3JfIpj
mWZlKkBs5XfG1T0fDpN4NY0Xm7yCKhM+ZnNW4T95GlAOTmcliuq+AbCry41p9Luz
hjHTG4oRcrxe00/Q9kdg+JE4IEq3JZdyWhhxRaOeFZt3u9nbL/RMZt2FE2eN7XUA
Kh83lnG85PM+2QA9eiiFJXU3wnh8QTiwgjtmx6tzgtcOW8SSmpZesWYVuMV+z/K1
SFGcRYBLB8K8mF4AJU+AXGN0HAAbCxOMZ/3U3BSVcfusgiN3ABECRaO44gcL3sZA
YFX2hSyD+Ca8JrRrepf8gLDH0PkpBtbhFtimde0lNs4pFamLwJcqYTES5r/kvle0
x6dROqlgR4+i0dGDl4lxVDd91rzYBTFwyE7BuptyTosjr23ivIZotw6EqsINgcQ1
6oqBPinLZput/8fLAOOEtDJfHyYe/9HxmwM3/gO8yi/EQmp0fTo87I79Tjj/ETVG
t9odLtAfkH1FElPlmXe7uTeaFybnu4ae6wnY+EJQsJfuhItRo2nXtMMnyHYDO494
bi57n4rPgPN6YWHDdRBuMfFAMCnvUaiWvJeDy0VFILqby3gYdVrTRhIe/LonRKBn
07n9ZSH3UEYLYnIO/3BgZkJufM30Lt5omuYmL1ppKLia98FCflZLloJkD5ORJSPj
Y3YVNOeN19jkify+dPO+li6WHKRYCZLC1YptG6E5lNBG25GpZFRUmXHF6hTgw8Py
9Svlt/HOLxhs1Gjwf3jp8gBmxq3O2vPNP0u/jYZYqB+8wjij6gUN2Z3j8SSxf04f
QOoov3oq3PuaC/gQEyNUtj/SxrJWNg6AHK0pML0ugycM9H+jmT9VhvWVVmduoSb+
/0zFmLap6rGeZ0gS3JD6ANUNJY/bHjLzxC3f4E7N7bQECjZbJMjalBNf/7QP01p/
4A8lHt2/5Nw5UH+fDXvL4VomXAqqToWbE02JDEla6dfEzOGXxRC4otLEcNlfBFiF
+sPHyDHRDgGxfjZRi70lnfK1eMn3h7p1mMC5rPjHyubrLsjNPIDOYj1A0GnM4EeE
YcJXSOGgGMUxh1hicDms4IeLjPIKo0IQkOQRZJIQVkwX4oZajrF3mVt2GnAojxBd
8gA0858nrBo4JcYxUWZlYlLRvZUkMtSjBOUjQpTBA3PIElPD8wupFO6Kylax6uIn
88TNJ8jH+PpywWxwRiS+Epj4o0Mqn914OcJVaowrfhAY4nkgGM9JOMFPHV4mg84n
tunvnoiWN97Zs2a8Mm8JElAE6JYDLp92Mfy/NKPtMJZs09SdJ5+dBHxh32yZvTRc
xqx7qOyxBPmtPbq997Ahqt+RBE0HKri/fu8YrNT6CgXOAMiQt02/fLM3NVmXkKYi
k+ZHWMhCpyTSK+st70FjAOkKnjauj8NVQZntwa3yhD6d4VLzECD4pb/GwfA8HR0y
6ZCCj7lpJP8kx0baszysiUvTUgdDa4iqxH7gAabBg5Fkr1gGbpQZVwCuU4BxNLsD
LyEurYIYNulFS1s7VTIzBAzyrtQDwUvCgTm2TFp24bJz6oGVrw/kYebO1W5ADorY
ys7Pq7/ERKaERTx5WEfk6R75Vz1gXZQMYbwnDkFjpLBpR2Jkb22DTz/Z//UEkUVl
W9oyrYN8BFgF6/N+6XiVD9EEv9iVFCtVt6GDs2Kj1smvGq4VQ6XEsczjYd8FYA0r
+p7Yhv9xzYo0v7nwjZ6AKnpJpw78wqk46O5CcQYzcimkuY6I0+DRUGs3PLWqovrA
zoG7nYnoxnsbnZuZPr8iuuX4IKtejBaZwbSg7cdl9J6zsn9HNFczX88of9300/7J
0bxvMBpixukv5XEp8pqxfOTrv5ly9YR7Iuc3ieui+PsBT33uRO6idmKmgT8+VCXB
Iy0Q6P1tC7mSr3Ke00mihGXAn8OGgaLcGnl7QZBhImDFMx/FmwzKgmUp9T3n3Avx
9z/bTjqrTTh9WexYKoRgPuEih8iRWN5edxYNinZsc82Lary9/wQdtTzvU+PGRPCV
rKDMUpt4e5Wz/dOlodnint+lRvRFe+NMXM6d9Jt1Xv7FfspQ1lP9HoLVqeUXyscl
MA3wPfcyQJBmUtbgPjMTytvtJJqr0GFTr089e9oRO6jhnkxwa2wKTROI1IMvlWHF
+IVXNpPJZZXKgBs+Qm9Ny0sxwO8x4St9is2Ih9ytNURYfWiWVJsR8WMKLq7JrSPe
gtH8r1Z2ffNFyfb63vKruG4es205RKHDd2hIyo4Gdq83zVeFFfWJ3CYW9i5GWTv7
07K6aREfYPbjey0raO0hMmM6Lne/M9FkAHUlJzsHfHz6dlaDi46qGoZwYfvPtdLY
oE4lHlgsxB7rQ/2cVMtZO6IKBCRCu4Wst2wcswfS42X6sR5BM8muyJUXu74bHVQh
rBUqWvLa2hZ6EJyXeWZNvyVIIJb5lcUod6loi2SnVZM6MhiBPbr0t6ivthIJiivK
EJsvFmuPscgtcjtDptsr0uEymKSF/nAChAJ0C54pm2B9/cmgdQY5R7BlCcEHAcxe
6LxatNwCZtfwhcG8RNtVnOxP4WKuh2zFQQyXvRX9utjQ0FIWrt5q6H9ENyQZHvic
gdY7ybXhodcq+nbssEgRWm4s0rCauQHPozqL0fiBs4ymtEq5Sgq0jwTxXjIHPvH9
TpRd5jhWz1GDKZbWuDbKRLuRyeS4kyNnpizgYSBEmYWMjuMeJdVkOMUpxTVUqzIT
3WLwQDbJSbAuLoOSBJxFSRleQp0YWFGKPn18tHcaXw1+zpmLvJ8wKl1LGNUPAPfC
YUEZcYfMYHkH37Bg4AxTxJO4+tWT+wswD7x8Y12cBEGAQ82akkY/JUcZduTNcMIr
SdyONc2uu8fYGtIeeuIRNl+vktBaxPvHDiampWPXvCgyoBJiNMJY+XHWmivEPOBJ
vICZ0/tD0Lh+Xy5ah5+U0HrRt6/0s4mTh7J7S8+2e9foCUKs+sYQDuKeaE9TAvPU
oxR72/S+FmG87PePbcBMrEDy+Rm2h5RIPsFiB86T9lqnaCJk8JEKCiNQfnMlYAkA
OHg7RkpoHx063u6lw/7smLLKLfKBmgaOETkOfa/PFgVqCzVlBcZrLQTVavTAjj7Z
oH4HhVv1tV3wAgsvrWHmjdMcx577dm0Xl5h2LHdpoNe6XKAZeMRZaGxPKz1Sox86
h9ScIlXFUbs62iy8WOGTPDkWKdn3RLW1VmghtmYMGkDNseiONlj5rZG/CapeRoBH
Z1A3jjZmMoGnNftPaZUJvd1elJH683Vpt4jgyxCxFctEzapJ19JA9qUZIGNyEdvE
EFh0q7kfMFL3zOFWo0hWpfTwd9fvGqXZGnl8xo0z+Pb/kTrG9aZ7rnruIIsbwhya
BppaZdsKZDiz11HKAG4zNdykBKo1N1jwzokApZF1gaI5S2atvty/6DR8ioz8Jidy
cEKpWr/XNGv11ojfCmbGN8bmU5J4SLMQxzilAbu9lKqcOXl2ORc+97VY4wTeycWI
75n0Vt6oC/t8DHzGuAfL+bv0cJTEeGj6nl9z9cnTQzasJqUJ/yx535UY0Ph0LxZZ
s5wVA9kBpyGgcfKlTFC9idcNvI9Z7mS4iYPc83eoF+oqMZx94nplyJXNRwWjfUgz
ugO4TIjiAdcP9UiK5S5YSO7n1Sk/aqG2I6XuSKn3GP7Jy2xc3ApZSxlXGUaRo618
3dwjTjDwKI8YiYWSLDvQF3QHRgCosW7yi4Dk9gnRcqw7B52hlvXEobBTX1R7b2hL
yAgoYY6yYO8nIZpqSOl55ldi8GWFHXM4EVxPNlcX5VSf9YfvdkO2VM12mbWd7qBo
TkTxffBK9TjclIkYNj5foy64c1g3ur7ZoHa7rEHOylsmBI5h/3gYNtTu31fynCv1
2WBKxNpBXubaBbzxy5hMMbIzA1scuCiBK9TVV+FOuGIrAxOQXFVFgT7IFP/1Pf0Q
2pk5J3CDHqXibKXUslmaG0BIHV9Ry7taFTxuEx02eWYocPTEGfhjmfDkiTRISIin
pZPFJg5js8IRwUaasS5+bZvXocURZ/U7U6IcYabfavMboC4G6HaA4njl1Mcd8K+Z
r3i1VI5tvVJhbGiuS7WIO6G38PvSs5EqTkj+kqh3GO7bH0yNJStaMqKCA9RwaIwj
O57pTxYBBSyzYftE95gn2itQr8DY1V174PxS3i/6MHj4Sz7qj/hm8xm3IcVuNe32
sRgYb/PxJlth9LukeH/bKq69hS9zDH294j9dofC/I7muZaMJmAx9D3NryR/uzMxT
FXwRLoUtHFbyfCS9N+iG3MKgao0iJgU07tg1jkA5aSGHQmO0D4MB+eSBxSRVDJx4
yRzXq50XhtDhrY3nXHtMpxZP/p87vqAkjUEY7IIMgXc1KO9mzM7PJgq2WzULTWof
NoNIxkbhC0LwFTqY5Qac3MhsNzSAO50x5A4T52IfrG6hucede7JyIKlIfEp0WYJF
mU7QLfIGrypZUrfagaKmDQK6otFe7UU7Qy/ZDhIn4B0acl9ocm8NdEl0K+a4C73s
GQejscT0CTUSssczVv6xjf1RLFdMM38k17mSzKhzE4rZ0Fbi5jUi/5LtzP2lUwLA
1OTVliIm3lA5AvKlosB3Mo9NjvEpm9xfqW2B2fZ1vr1uLNPLU2/YT0AEQQEze7yf
ZYJ2jTZDFTwQPsoMrnd5nmvqBUKVp5gIPWiHJ24EmC5GSLcFiKgo1DVkkjCYDb/s
jgR0wuHlrqd+ZKFtQPo1Z4DNlyceBvnQcugpmP83gcv8EGxF6xKUn5Cg6pFUkx4z
B9aWVoKPObdMK3ny/68zkMSeW0Xh5k0zCI3RjLEjylvk3ANwNih8Fh3mgYQkBG9q
kTOqxUcNvaRv23PoPOM2b8SHfRfDAe2LBx5H3PNwOcTEtrbpxKbGV12KVgnKnbC0
S9Q6up9A9DgNx1BYqfp8Z+p1tzYgrcfUywo9pNMw32Vm0q5Ex7pVy5bjbSiNpXpQ
79ju6pqvUVlobqajs+pN0pkcJxeeDfoOoJ1eBN3fvI7t9wuaDGEDyTO7yxYWKYZt
y6s17Myja7eWVaE9ZCIXmQAvlSscH8li5wcGtDOVCMk7bEAHVbTi1BQybmnmLsDi
I4U8TQxAIH5vyozs2y45wB9FC6noTFUGEs/UAD5y/26Mtm3VOmvuIlHSJmQnNAqo
T95ReJVj922rL29Rtk9S3x6bw1akk7oFZczJpAO0W4pPQFcTSy5R9eQpXP7VZM6z
WAd7Q1rculN3OMp3XBYQvmjF2D7hzPd+O3XXqjxYzbEMfg92lxwdOTRzOO7vVp1E
UyIzHjDgChFKy/UCmGi8KqFKIlcC1sJfGbwpdwiT0Z7anmruJYC49e7Pwo4L6Xk3
l3Vr9y/g8e3n6cxG4vouufjxuEzbJsuEwNAPED4g95D6vt64V3PzestXkiLZMx6t
HqQUHdstnYoaFGalCNmuSmxV2B8UwlGOuXwcOhdZtytigK3rcFVTCBisCqirCNHy
+EhM0OV+LxxVmE9ym0snNrRoKnBR6ogLfXOzHccU81e5lmn1BfPZY11ygfYSnsk1
qjqYa+IitR6Cd6z/m6SNv7Dy0sULD7Gdfr/8PJX8wVUPyK7P9njLf+xrP2SNJbYC
Z2KevzVjqs9XdJTTsafFnWSmGFJWr3/TJZboj3uLbltsdLVCzifvHrfjUBBeOmQq
1gR1Mql/nvPlfzN1N5Ck+PTB2dbD9wFk6F2aVS0dL0jx8sGp0e5wfT1hHGomRW8U
bwRk8scTX8ZZWBif2yJAcX43i0I0yhrixYQw23yl744PU+RLSAfBQGsaR+v0d/yZ
0iF90N/aIcrSO60SkQetOahxySzsjdshKAza3AaSfX+XAcPwggS2Q+ewkFQk+Zv+
HSU04xyfja87jqXFUUJ9NMhE4J5Ib+ud6qZ4Y4/2OurISMDN8ziVesW/LvTActtC
zE+KDPs8Cckn/x9QAB96Gm+zRbPxayttrypN0ljepgMTv81K3dvu02py666kq1PZ
sVTnaqQmBRw1ZclbQvRIeuogJQhKneF1wxdmJk6L1QmOAHxSN10KsVaIESy9RA74
D664t/J9MMSbdpcMB+HNCOzpqpNeHpeMV0dyHBM4yqyURm6B9gDjMtUZUkdSg3e3
VmBY01iQ/APf4jlZ6iDHTlBP39xdTJLBUamt6AbrbcLoRMo2yAbZzVM1zGMKPPqv
bsVft7EszFqb2j199jVKFpBnvN9cwTL05mlsB+gLErmtxK7rmt+Zh7Pod2R7/If/
KPqZ+ky1QiValwo3pr/xLLAShgZzdjJBpVqounrBNsW7MkWy5DW9ymFcEh+i52DY
mv73k1csZyTybEmNJS+r/Q+WuDchd0vFheqOkZ+OiacHUaBl4QFr3xJFL0nwlW49
v7e5j1QYQyYOGaHMJwUDOIKE5Nhf6f8VWz6PROXLsRqVrqmPRuSYq+Mv/6ixQOmv
szo43sXs05w1wkgNFd8dywu42ML49+uuoYp9aNFvdkhQaUuiO6ZlEw+pzpP3uM3d
0he6tCG7sDmJXjV0bRuOIPRe3lVECuPGA2i3tmRPdHsMAvXWGmttuPM8pS23rh/e
HkdR5d9jqpppGFBxaS8dInVh3wU9/3bqpApog/0dmYhmklKxXUUjcnMmNBztuTzZ
tfVWNONzLYrtvyjaUR1ypEauaV3x0QkznRXx9sUmsT1NAlywDxI5yfsUsxcFPh/1
oZVpOuXulM2El5tgPc6rHjQQTe9thWoMH/Wd8MuMa1YDs7mm1FVjjXg1qg3FaNHa
JK1CePxCRVZR/+O51dDlktXWaMcsmpofcZgUfUPlp5mX+tPvfmqiOrgFZZMC/ee9
OECy3jRiX1QHtXVH0aQv0ZE259TAecFlz6bi45tlfF9U/5UWZvzkL/UvWp6dmy9U
KY2c8UPi4AjdRcoWnSyyXkXbseh1tnuXroPeqXNGu6yBwx2t6wTSA32I9G78tx6E
nOHwNFvBz5OqO8MsKuMjTp5aSKdnQydu2csmcVrBJkw9LluxvUlz/Q1Ij3FMOI8w
ilKUqYHjuDRNksv315LnW1pw2jnesUeqimAt2MlIVGaLH1pgDIEAgzFs+5fACRhk
UD1YE3vmzpIWnHbI8/mqtUPTsKHp4QKLtoRLRFZDSbmszQ50zXlA3Q0KEpmXyMzL
vEtKGdCrHR2MXiZFze+qw5o1DKLevzI25WsFME80MPxuBKwt1tV1zgL52hjmVyF6
JqJfFzUVhmNXHe/UvVNlRgi+0CjyUdNDLUaTeF3jmcc66WgMqG5XfVGilJxBUwZA
6/F7Gkz99W9XGhGgGJOf3f9XywaXKJYkl0w2ECvhfbE5B1fAtu91hJBxokkN+edW
39DsmQUzSVKhFo6Gvykvp1wn7HOQ5LJxXcfxp775Z7UpQfKQV74TjmXS1HK5Bel8
BbevFaK2PIWZbu7zQeKVXo8U7+hG4drU3d9qn5ZZSpupJ6P4D875tSj1R7k6i1wB
QK/45tkWsfEbLLMOusoWOqQ7v6EnmGeFYEyTS5awFnF7rzZDI5IgUGITf5MJ/QoK
V0ZAo91VICRSGkCQc1UOUBXsj2ADPsiavJV67GSuBJnZ10x7c247LKsDfMD3NhOU
ZpXZEcptvYLaLeZob8LbSzUgYmFgSniKBp3dqoLdKKk0+8P9/aP7gsp0VQd9nedX
AhyY1d5IQLthTu2fG7WSoxzF1Ap2OKXIizXoxbhZMCzRab1mgZBrbU7PSMBy8luP
SMa8qBFs74iJ/8X8mCNbJxVfAr29n6UsEUp/NJ3odVoqxXNaUUeuu3XEqnrVb1S5
TmgHthgayJbuTmLPieEf7OGwbpZWtyUdRKRvqHwTijz++1WS4toZ+RT1mT/E4wmV
ZGv7qpfBshMIQ60mHmo9193YNOKCVLChYTBqjKrpdGtV69bctXvs4H7ki6sHpQ6e
x2VWqWLN/5tvZ0EydsGoV1wT5ObbkMiDyWL6R+AUVw3vS/QZLYydX3mOkF6r9iit
Fsf3XCZcWYRa6BD7udeljVTu1vksagdjGAt38GysXB1l1wwKH21xkgrt2Xl2CY1+
4BygOjCnFp56HQgD14xFAsmAEHJNbvBjCYaJiclH1snbQp+rqugf4LzQCtFLsXfu
fPzlNeQTCLar7oG96Hdmc3w+dnxAECb6fQ1efzk0a5fpX1B0ws+o/JeI28b2ADON
YA16ZmILvhyvjX93x6iWQX5pRyZKObe+FcEpPc5HeZ7NivOf3XLc0x3AxwslrQO/
WTogH1XoT7fSbIyymjPi8aUh3ykWReYAGi4bh6CId8rh98scSEfwR/Rh+kGj4hXB
a+slDxCJ+2T44G1OxXEiSBDH2O6kDiOfbs8KJIEM+QUz3fW1H0CPnYan5p0gnaHb
r4SUMPc8/ipA8z8xK3xrx614HpSSigF0pEqT08ci3WQdviSIc68fM+nIwMNWHnFA
W5IbE2EHMx834l4nqQQ5EL5mpt7fF9VHKZ2aO5bd+DyQ7cDPU7649dY5CchKkFXa
zQ/zdfJjnTn1ZejY0BTENqasajDSj1E6qsjLsLeKXHTQnbqmv5/P7B+xm3s4H9wD
UnzQcsVMJm9RVuJp2OL9V6XQwmiVGZAK3m7W3DxyNTjoqUJvMaJd/etP31bUFGK4
GBEO3Geltu2egOHWXQjbjBJ0o18IVuxmCQfvOvJNi90JtIeDaI5N/OZtEhVDqH7B
kcAVxZe7s/jLWkr5Yko9OrUQrUAUDe1Qx3dgYw4CTpImT2KOmcd3zjx5MpId8xfH
9wdZ2xnickMjbagHqfSma4aP9MnBRW5g7Ph4whv5NjxGsNJkb3ODp4EEEzZkewrz
plxMh7BdMOLZVcuvGrQuTeedPXV4ttwYrl23dAgpwjyexsjxW9sRKlCb6XRpDfWg
l7RuhCunOnb9LyiFsJ3A59U4E4AvY6NNBJYXnmQ8j/MBQ7q+2fiQ+BZw+Gmn3z+U
OR3ayJOULa7BzFFjEHFC+S/aqMmiCK0JpHceDRgTECnJAQFi89uLFgQFGrk7bM7c
5ZVGxBagh9nvAhB0TIagYeQ8XV0WtTifD7cNBxFJnLElF+4G5iQjdl+MZjrp0QJ4
eozCdj2O+s78T9pT51LxsyHSGHOcLRNsu76T0/d9DlTrwiiVkU0ig6R5nReY/DWT
+z1guhzzRc+znxMAuFQlX3NpIjCXgv3y6jIRVFT8UkxKtXWPQKfB15kkpQbPsEx1
7A3tEdDyv2AeNrueUq78o14StA1lmjFfhpM2Ilr7ycqt+OrYnwH6FIAyumRljwIQ
K2IEUvFEvgNNefgyd5vGbVpN7f8CKBlNW3f57W7d3rVzsfD/Q++9bfNLxm6ndIEJ
xjtHb+j99ef5KODwqQF4XBaU6nFqKKlOiBUVKo4IPjsFMZcdidHc+opxo7gk50JK
pjYY859E8//4VHZcvdgAD4EFwP9v4qbpVsC0hqdF72S0tErJetGZhXp304C3JcdA
o1FNsQ/mMCUD20IJtVIDJzQmEzGy46FDgHgsYucILJYj8a5lssF6QMqqLTbmnuNk
h4OUvY9vBm81KZE3TWuz/elkEAIHkAKDJ+901wZ4rbj0kJ3luOEamKeth6aGDrUG
uoAdCGY1GetaXMLL2SwfhabCj3tQVCGC1LytqxA9pnzI7JoASn6CmFF4k2kC2gQi
ug9FKF7X4obGqC9bUetpr2tqOG5ZzIUoJzdYgCVbF1yz6IQvlQyEOgEvKQXnZqD/
UP3q98xkxy6XkuU5kPuEri20hLJpyJfanvS5An0Oh2GC2huQgD+TpU8tP1FKY1VI
bThKIMPVjil9G8WIH/UKRO0pvyf5IPaR1AEm5wrj22orG96+p4A5ZgibZ+bGK2ff
vKR8XuyCHlqt6BMXckHSoJ5RMmt/Q4CXbuxB0va2MKtLDKA+DzO66ua8WTCY+f5j
7G3c+cdBDMMRTeT0lkcwZFu7MlKDeGG/V7dAEL85xEpSG9yWz2Fih/LCX0O6fQEG
18eVTHIEccabX+otIYsdqUGPyVuDy/nvOtGMTMOUFXfTE1zd8CwqFzeZDsbcaGhd
BMCRN/IHu2eQgfE/4rLW3QEYthWtSYBCzAj9OIZ4Uh1qt9aFCL9JXeXbEvtm5pgk
FDZKZDM6fhVzYhJOr5gb5L2sARzxB9Z8iJnPCprEXoDPgRZ8WX4MBETN/tTH79sE
Xx5H9i2J9IiALeDCTfEHagDws2qPKepb0EB0jzMplK5bOf4tuMo3IcZNQ0nnlLNN
NeSLt4ZULT8ge2rkiEvTXG59zdFCx3srv6Uxs3+BNqt5OJ2i44sRADix57D8iVO3
2EMULzJGhf2pG7GwFG3zeZ64kCL0wdCcgKEIPO2JdRHYyf69TZqBh8RrcwKWprx7
7LbYPM9tLBY9mlTDc6EoJYx4rVQGB0Z8MNvddcrni3mwhil3jKrZtW329aUJE61u
ypF9m17nQDRYG0q6wFS5Mq8R8tyJhcWr9Tmzkhxs8rkMKhXpH6Tmb1B8Ez+Z9VlD
7XCZ/u5NJt7PY/4BfWvPiJKzM3siCC6SqTH8ZI9pf8sND3fwhtMLB8N7EOt9Fnx6
KDfwPYt4cGdOgfspdiJVmwqyMl2Vt9gRiNoojY/vnZz4CwM/c7Pa6WU+6zc/HpwX
YWFkPRif4g3FKPaPLbQ8zbaJrXEbyRPXJSkqprHKd+L5NMyxHJ0yJHdnPdOxPTsx
c1MHBuav6B/mRPvp623MOFNA7hLbH16xQc1Q+Z5MhjbHGj1Os4OVaIAlcwRd3msy
zCxknvUTRvGppAMVtvlpjYdHRF6ILNVa0OrkL7iiVmXkJDF84pjp3biBrxM0ng14
1mKewF3TB+Pz0sPTbo6NGanYCkum+yukjmKk1W+B2a5sJPpnMZZxfmUXr12u4eQ+
vxO2W86o8ABFL9yApycniKCAlZ4ybEBLWGS899YaEU3gPBFewvS8LHNnpYcbAb8r
8/+HsRCVTvrfQnVbGpdfsNytw0YnpL8nV3TVuOLNtpXjVVhILYJ7s2qij1+SImTv
5uRrAP1OpD8QRgc7f0B0XyHwet5osAa4Da+kMDhJWanQlsgnMI2rCnROq4fCT+s3
aVIG3kNgujgWEXAaNIpgpMhsdNLMpvniNjUUoNiZDLCAh6M7/ZLI/XPdFR+4s7Mc
0YwMnlZ12EP7xvBu+11A7PTipXYe1DH5wnlVP11EqShRBQJT/xVrXQo3WjIy9E2N
M6oywblz4ppBj8SMDuxiE6MXdr+CnuhtPCJnfKr8eIs8DKlt+xOaEYVxdBj+05Rx
JNJC6UXRilrrJaqSjden2nbWgEstsvZ3uDLm97+yEI0kxpIp4UuoPLo0/uuo9Ms2
owxrG808OuK8ykbR2Fy45EZApD7/k/tUxeRL9B0Odwznna4W5OmUSZyfiBSzrcCt
irZfRrqvH1GAUDvQIhWR+76tXaaMwWGikyozZLwDGPmqUX6wS3JRNvF58CHw8x9P
CycbzGiwiRIpoS+ZbM67HNoCQs3RLTbCcFqLLcLmq7U9t3Sjp3yBdSn0QuvZg0Bi
f9Cm9g8jaJyGFZbLWXzC/mHkJXyKD8bHqbC4BA8hfMOQjDEoBF0TCDaFHdmhAJ6+
axe0HCE6fJBU/nwPY7F1zmNJ8AawPmpwBwViin1Xm77FcEjP+TWf5lo5BqDKRjKS
Fx15GLNGEZ8h07p2cbNkkSyZiCYwglvbvK4D2Ek4JWuwY3pwXsOd3MiOq8+ddoSJ
Tv9uMwEgrqI82ZFA7qLgeyjdctBm23YTvZuC3GpVti1W5nUHlnp8AbnZtK2d78q/
LDFMC5gs4h91xtqqZuVMt5L/cURGmUjgWRuJPfuZwm+3dW6lxD2gM858fBwyGY1x
e8PM21Aozyupw7Nvaf+fED0t+CeDKxu2cHOf+oddvoD0/iKGo6+6w+MHuNW38z6O
a8L8oazNP3kBK5CbD5kYa/KEI9N37DmT65QTHtjodjESg5/xJHF7W5/uJTIbGrX6
O7yb/mld4gJkwpYNIwSfk8QR6qDKKXzulZiDTpD2FV91/5vriPkHUmV/sODPc2+G
UL2kpybF18EERGvDTJhbtj7p0ajVlM+JOd9wuaJTX4nfXPkfUriRUleU9snVttCq
9du5+et5W67yCDoqvocC3sU13dml2n+O2h+X8+FKgtUFVZpksM9AllFoK+beNkDC
JFLT1+/WcX7GzU5AIHkGCFYblYgSExhKSUPDEcKmRY99nZiYcECvBIfRn6AmQBoT
v8f35mJTBZNC31SH3dzSXTooyd/bKKXfAhOE+irn9zJHDMKJeOKqjl4cmd+Fswcm
1frga38VcJ1aFpB2KWE/ErofvMuyDWQKPPoAvIu/LY2Mzw7N+C+a5TxxcaqKuWrx
/zw5jpi7CnU0BgJmpl2hDCQBT1nReCapmgizNNIpE+UP8AStZ/E9URIVOi95+vVw
2j1KtsTAT9C2yYyYezRtGym7mOS3Mh5/Nr9QEvPtqQ/yYye32FB2arhjQ6rr9KNU
kGvGm2vUaVVm4DU8Om3Q5amDq4RPoRmePkquiX1bxszacMmHlVHXVv1Yifie4PYw
C0Vby7WCSKdn0sNlu8FHL7EJ1z8NdCgCXKs2DjKu08HjJXaiBu0j8AzAJDkt+k/U
ydPc6VfkOmZg2/z4CtY9xmqDvWH0mYqiJI+OvYP9665OFXnetz8w+GxQynq0mK6V
66xUe5Qin3v+xoyUjFG1CUNUfJjk2gHSmdV87HYf6lHi8F2kFo00gDvHUCz1wkip
x9KMKsaVKrbIbzI9v+/tOBaohcAbN2MsnixNGaqnOEGkpZ4TwEUMsU6/mhHt58kX
r4XjGgwatYgQ3dmcmA/jVeConcAAYQbJEQeMRtwQTSZqom71oiVbkYb2qy+ffwU1
aqUcHlCbFY3k6zzREVmpLnM66TvG47IAHVkfP8DXzxTHGxPgHCt47afWrq0GLsBH
Rtmy+QkcMW0V92oRT/blExBagODDY0hEaOnqVpiGWgHVz4CBn10BwFzYZBuGOB3G
YEMXlvYCSBqidg3uGLoJnbac5J+xkpLWtHHmU0yEBPwMmKdrdH+qccuj7szq4Zrb
5+esfauXWHezybd+3rPL2rC+I2RcQKPEZOcYvDqYJ8F0TcrcUwZUjXOD7Q2p9xpC
muflIoEcRv5qqGQ9JFwsZ7g1FhZFaLIt4WF5d0TGezoev0hypnj3KSQun53fi5WV
t922zohpb+fZpE4lkuw05galuBmpM1/NDYXIoVV1v2X38HmJKBmsuMeoXytbqerk
3GJ+cWW+OSFV5Hm/pdvnF4Yv19Y4TDDQO/lR8NIdURG22L34UO/v9GplY7EXGjIO
s5ntRCHTGtImXFMFjnYEGr1fKwXcUbgJ0CAH6f67UEfnMVwI0D08eJZrtUYoo+wb
+Q6sI081B1gZyasBKSh/5oCP3JJtC+YeX/wTNZAGdbqRPjwAFzbX6M6UkpPR4saL
KJNuze1jul0jQDQ6QSNuJz6C0jB6+nUGPMh/naZcPeGI9wRpfxHCy3lvDm0DvG4u
ilVuCguBglVrPosKWeCJIyM5YBUwowJFfNmp79DzNznMoCbhounMage8lGyiXkQF
BdWVFZYSn4b1xYeIfilRydQGepI0UZq9UmXjSivbgEEaYe11W2/1VuXM5K3ltXqi
kYcYNQuyn4PWIpo6bkcEo8y1bQtJTeCJO3R89cLr9HnoWuYqYKfdJikZvZ48xmg0
XRjLN841kPUbjgJ6UaQHMmjPngFO6G+jZztmLfIwLhuFl33sR/vIBg0LxwPctZ3Z
6TdmD0wlqXhI4ha5aQb9AU1ho8UOSDvnuok4wWiBfrw3jrqvYw0M3Dj/UGfzQhe/
1RRknBdLAs8lYwpkMvcvW4uAq5HmQhXwLCvCr/Wj2FSMrUsblJtlnhqKgK9mt52c
7cvowfS/nPW8vA0XXYL1581p2yq/5W6YcG2BBcUavwqtPBEgzY0WPD8b8hkMy57F
3stZdOvis3/pJkmd4/jhg9vTvAckNvtLYHdaKZW1c2WIa/u4Ctr0+xDDCO55T5Hu
u2ahZ12vF/bdu+DqzDA4t05ed/C959OPBiZvSByDq/CmtcbhaLPWg/uVx7FNIaE7
pMhc3ZtEl0oSowypS5xWsYk1Ce13P/C3zucE1XkBj/lBBH2/ULD0aa7hoXQjs6n8
URgzeUBzulwyICfaNfeel36r3jsm2tShbjUV0gq3LwhNiC5ZrCXfoKKM4BYuUMKE
NxLzWSdmOK3EMpMyXAIaQc0kJe1JMG/ZfcJASTcIoagNwf3ZZ1RrCi+x+JeRKEHv
pXFpgyyZgD1H4mlxtS0JSSjPJRG4Mcnj/c3slB9wLtgCHvawRYaDD0TgVwCm7Vt5
aKH1GELq9XMxa2SookUc7+18dtaGz+Qq0eYmhxeRiZWcnPZlrpBFrhrPNWITlUcd
J+jVnTY+WtumyBEl3Hy3vSMZSs1vetykbpUVnIKTf4bD0P3VQDo/wYYsPHW/xMve
JXAclmaH5dak8j3oBGLhgLHHqDwpHA2hKmcr+/2EJn7k2dzzvoRWUV1wQC2Jgyt8
zCPtT7IzmTBFc9vCB5QFU+41G2uwIXf9mZKvD05v6ytiJlYNZqdVBZIF79tI4EvP
4ywbWYCH8wJ0hsecd45Ovr7pncK68qXzXcmaFLtGnNmvDRTQmcI9VgrShO3oEUxm
Mt9EcG+cxjIrYZAckWkcEHs1miAB71CfaQhdXVe22AcPmEwgCAE9YGXqHGFce4ya
9sdrzKLd/NUicrKGRDsGAqmkQ0Rj0AkaUsuKmpAe4Yk+WH/7Ue+ohHEwtosWwLjj
G5cCcCcJy692pi7U0LIhvUuBsx+UmRu+v6rb0PJnbB7BRezmYCbsccNsLgRlbgev
4V7g7JOSFCP6NtCaWNhj3b6z8Uhqhi5PsY1k2WtUiqkj9ne8LHk+ojKpXgonmSSF
eZgA5zqr8NmxwwQcRSmKB1JDPQ8xO/SP9+FNn+qvsFRNduuIJ2C6hpqnXSDAJugy
oLHlN7rfWh8hFjuyNLm9QesRRZ8tRvCSajwjbmENwp8Zq1vQt6DChxQCJ/VQvt5B
gj7qb1mhnzVVkbctuMSYXpasIHajPuoFAvsfd/U0yQLXaM4Rt2EKXuUzdJOlcCpc
f8nFDyZS/uoz7kamtUUoRVwOyM94a4RL+pZh2tpNv+TUbtK3ZFv+hHMZ8o+6gl6k
AWFkrHJwQfzwfRDF2D+T5Gb2GXcz0x8JKCY8rwFTF1IIKcX8pFpnrMEJ8eKOU5Oq
ddrQNrxGncCa4Xw5LlZ1heXF3cNu9ojfHBS+Jsv2TWDBhblNCczqWlGgZhZ8JAVC
ohhprZ/vhfRIC4kCu0XHqXEmjJk3oKxq9p5W/eGjjcH0uMxjrHyyanXHEXokAk/M
ES6yKIdMfuIkVFijSk/5AiNfpEu5/WVaRqNuT367Am7UJUcpc2RqDa/ffm8bHjTW
VF2Wsuzj6ipRlEy15AuUrT2kTjFm/8gtR9qcfE5rEhXS0tjdinocg6mG9vXcNFOt
MwMlU7flM8CpORg1zNSUadvdbD2gyGsbO6Q4JWXUfJJIQeBrAhmf3Hwy+DrUo+ZN
vC5QFBzCXoEXkRQ9h7TknY69uVfSzrY6n1fZS+wvZgg+EhaAXKnxRzqL3msL0zTN
JZF9GjAADzelWUjb8e8gKPhypVuSOPhShWV1Vnjllosig6AmQZ0s3+xoPd8qRatJ
klnKpofonPlvpQP0QY8B8GwFU7moXHDfLu4ynzYcSFVbdw/vnWgmsRX5dfwST7pz
merwPnunbdWLD5Smakf0askbnO8XrYYbqmUF2zy3bM1XD4jNXQP9hJ0hnz7wmjqo
h+4cgPpajiRhHXE0XXvzXHssqTqOz4OfQCRuFw4yilbKRq+0KRQjxCkAPodd+1NG
MZLS4taIg2V/EiRegu+fN/5wCRMmVjZXMuo+IT5ht//c5jgRv32KeEcOjv7HLXF1
DwKeAP/Rz3cQWitMkZW0fCfdxkKw0sn1V1p1igtZQEq8yUrhypcfPwQoFLAVMuCa
nC9wa4yyvVdWzyY/dyS3E6x0rrwkhkVdkY4WCvMtCYPyK+G5QSKCsRwcDk6Qrse8
kIEO98kP9wLfB5IMUXwN9X8fnwVb91HCyO1V2YQH5D6QQBPxPYpE8YBF5XYY/gNH
NA+DDGn1nQz9WFiwVMptDRVhXv5FaynQUH5Nfw7R0wX9N2MtdED9Ol4hd7VbznYy
ZHgmO5OLuLCwTOc16o0tuooKSC/B14s51cYel6rlyTHJXba+CeXtm+IZuAOCiKl3
XwpRrvh++Rpb9cixbohSuxGqLWdjnnRT136qH36G1/oPY1N01j7NHpd6y08ms6WX
ukNbgWWUPAGwOpAuTi0OuncJ6memi5TTtC1uryf0f52dv8t6Vm7X6efIAOLtUV4Q
OY+8zF+G7Gw7VfjTPO0mugw3MMocANFZmQsktJ76CVXrueuY2RzPXGIhHfzC6xb3
TELb5fsydEBFSTjlwn2VleJWGfgPsH4YSeIxcQndGgGJ8soHkc4I5rm+6TN1v38z
iHgle4OZbUHrGv26L5EJJ2/LDA3M72RilIucpXyOkPbKrUIbcrcV+Q85k+tDLyAA
GYL+QgtIdxDWyT9PoVub4iIY12/JrDCLp+sj6iVH6+H+IMQ5HpIcNtUcdJ0OLspJ
FliNCEq/QPK7fypHldwBU1BnHbF1oymjHpe3DQZ8B+KwE24scKuWmlVvqZ38Okc5
bGwGtxe1YrtYm3E2YQVwtXZBvsTXMx3MYUwcaol2hUQcvvABDTjgFF6oYlC6HNSW
2HA+1MK/zAY+5HWhd8vW2jGmKbDPT5UB3w0bG860QitF1L1woIXbCVK/jM/R9Rpo
PPSlIgwm8LFPHfZU19TRN3B1SXk+sADhpi/bVlFIyFxbHfKQcj96ROMsaJlOVKmO
hdaBoyN+omdP6lT5W/kL0zYr5ua3z3JczBeoZwb3iQrxzSZjinO2yUYCw0edNrD2
0gav2Ptgi91KUAMvNv1sbD7pGHHr5dJVVtMeHXv2mg5mjfKEtlchcAXyXPcNukxs
P5Vn0q+xDXh5ttgJ44k3N5HnxLX9MZwyPtUP1TNqopLH/Ja4yNVUm4DDmEQNa9ke
zhpNGKaBx6wEN/is+ib4qv9v4MYm4Gy2l1b//NYYyrar+tZS6/+ZxH1mbTVmP7TK
5F7akgO1DxF9nG8RZ9VD/zIW/L1Hxdfx/uDAPgBD91Cab/bnczGQQ0eoi4znHIYe
eagsYvru9qapsCxVy1QCX49s1yy1j3V7yELhFANmRftM9nwW3vUn7DAkHW0UFcp1
B1TxmjP8TR9zfZtco4HOpOXspkIs5hrKP2VMIPsvL3XG0mkOli+/K9+kX7Td8VtT
ia1kV4iY7bghfXMJNs/IxgAsLAX5Yt5RRW2/9aJ2qBvF6oTYOnYG+YivPyVPOOZO
Nj9Ijgj5w7m4N+ToVDy5HQ==
`protect end_protected