`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 21376 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1wB2ShNYedzmkmBWjqK4Mg3
8iDfXbv5M0vDNkp8sRs0MIcU8mAJtZ4k3nFhz966ecECVvb8/O0ZTePsczeAIhfC
HSt0mrdHR03GjzU0M/qkfMiazvo3mUGtn7gXTnxYGpG2iCEP5ru7bnLc8zJvL+gL
ED/SM+Ln42t+99cGra2zICP63aJ/XGMJL/NCCsX3SoRKEFB15KGchEIHTHP5j7ZF
gs3LE3dcTJnxeGp6uRo8NsHxXgHsHu5eWYPr4TdMgHRI+Pj6gUiyWj1bAMrlQePk
U13zfW05se5MODMT3DWI9MxYAJ/AmIf+CvwMsB+71+STMSNPOUrU2Z7cBmVJRe82
bsDwdXeWEutECgtV7/F1fTGLgy111NMuMzvD/B7mh4hcwq7+YiySr2JucDq13UT+
LUuzQ3w8ZgYP0rXdFpNA0LQPycUA4eTb7x3mQqcaHcRw/TpRHEvBZirUgRuCEloE
450uWUp0uKiNoXnSqp3W6+oPcFH+GftpZ03x8N0VFg5Q6PIC/HRvl2+t5Y+iZbqt
/YzD5EpiJd5zPYpVM4m2xVxBQ1vcrkp5KZ+5jJJqAQkq8TWGigG3awHmgmNPpTRm
TJhgFVv7sHWHbaC0zzVc0YgKgAkDSR3omJrwwsNea4mTBZQT7AM8y16HSQWFW7xG
StgFSemALXlJPRVEeKmkqcggkI+Exx6CMTEpk2BN+9KkxJ97PO9sDVsaTEvm64DG
FxLXTGU8wm+Ap9u4qYJHVUsvo0UWPlkj/pVZzHAdRAIFE2olfjslnNt8cS5uDpVr
tDuKDU2dj2W/K6hGYEkkp6ucI5s0yVgO8AQZEqJhYZu7IkFHPfaUS7xXKDeqWG1T
d9Bh8qjhfCvD3196IaceUNWMjMXAPgGsJtu9/k95soqPIXLjQ9mNmgH05AVeXMGI
86CT7dD05XWCH15Kfki8uiYR3LdnGMpoLXlq8YWYITsdJqSQyC9FfVi68hlFRBVy
AWJRl2I+3A4TAcPL2mgdI82PG7w2AvO9Zasy96KW1B5VzCp8UtCRwlHskyDhen/O
x2WbBzQUu2MGRmHHz+0kpDb/22mj7MfxhCR8WtD47Gb0TPYhm8JXVHE+ZQ8LZjgF
z1uTxQVsVBISKb/IA7pOCsBHqnXe5e1SPqnN0BhTA9v2jE0EGGOeIiAXamIdJr/4
ThNhoWFnnjfhzzF2GBv7BNdCzyluXx3asCyZOkNk7wMU2hNdh03cv2iRybHk44p3
Jdrk4gXRIhWk+5g9XMKqEDTznZHMdAztJlUz+0x+3cZ+QpxJZx9VdqNHhNlAptF8
An09YWnm44nz9QP+GGfChlqMgJch9saG+2AgJdMF882uWaha0BnNqmJGYJL/NoBy
6r+/DBm5n7GJlTkjMpgnhjj2uya4WvIcMxhqK+8T+K7w94lJunNhToK3NLWcyN3N
eaD7VuVvIeP/9byWKnWj2lm4Re7Ij6wtzxfTTikKXpeaIrRqWW0Jzj2SQZQEK1h2
Y2v6kj1Hd7sTm6md7eCkDekbfdUxqUr1/e+b6lKb89sgSQpGSGT/QXf5xCT5zSdy
y2OtO6JP8Ak4nE2blFCU2QDxPUQ5RH+Yc66JgGgxEATZrzBWYrcVcHZS3+snlFZy
+Ug2pZqdXTRqtaTwTvFFEs/vhZ78UvkFQkX8GZo1/mlj4Y8saC/U0BIJtwIs2UFV
8cL/FsWLyfO12Nki0+sWtCHYArS2bYWnTwL/myPgp3wv4oCO9Hjg6ehWJQYwsa2R
1Zd5zuEZHjAEhCICsFC6jlnXrgc2WnlABDj9yBP/RtcJ74bKbnXkgRfKCtAyLD3c
7qyCs3F8fhU7qwMYXlBqedeLAiml1cARfZbnI7bMW8d0l0BZvhhksp+is1HlY7Ed
DXuG0rd1xYWdCGD57zHc/0UqzV7tBbrxt+fwc6kROngZwd3Keg6wwKn1KvZc4Ie7
ADK4JS8+MCenxArjjU7M0E85PEZqmiu4dynanEzkMIB34fmr5dbgN2W3sp4+/dG7
opRiGIx31JHyQGWpHBIK9pvBTuVuLNrMoNzQToOnqqbSeyd1IO96YhYyCgSRHbl6
vQSBv+UNdw4kFZGtnFunYYOhMbSF05ALqJXuvgCNQo3duOgSfpz9eqIS6K7HCJ1E
Bjl1lKEBb50qSkSgoMJ6eLt+XMls62xuTATxKbi2r+FKeY9E2jvJXPWuQZHNj8bQ
HTJQynJEGMe181uaY+VuvC6fAhxDTeCMs3YHKqcuAIl/9jxtjpI+Kp+Ad5WCzVMx
ldyZNkIgj10ogyQFYNVnymsDCYOwPFFu8WeshIiDopk593TtGOcaN6MFLCF+Wy9/
J4C9utXMCrygqp+wpF580zKgSN+nuH9q2S2kP3ejQSftZFS3qUFKXUHqBAK7QEEQ
T8nGMMi+WmZ1RPDq1MUBp41bR1BNsdOLVg3/UehJwh2xpO8TmspHrBABmyz0yqjF
EQR9KaSqtF5U2jaU14i/rhGY8BQF9Jx52FSkip8KJFotMSaMHlcIJInixjRh5xib
eOYnMVU7HQ1RM4WRQzi8UktbGFptF2ubHLVW+Y5T6CWRWf3OjSkoY4aUOH1ofn3C
lBoOTArpfkHfjw4MSVVd/OcP6fGl8Eufy8P2ggGmeGS8Noql8/DK/Q3/v+Ftf/Sa
dQsyfg/awJCcATQhMYHydwXfygnJNXJWMC3D4yhZEo3gignxm03rIkLiNj5xon98
bYoV08vMKZWd2xXRe0jt1MZ8cbt3alW9mKezsF/HvhHEraDywNoZPLJcglnAHtzM
uV8xPRi3omCjKM0zUiADDtG+q9KkDjl+La/hPJOm30R/gEyvgAf/PW7tKF112xhC
WSOSHetaM66ONn7asPFQxdauF6x2U2UWsLa7q4ggPLcWCsr6reQz7Lf3TktUXBwU
y0j5gZjdy0WWu56r9PlJEuAEnv9P/QO9VpmADvdfEBSLWuRW054gIOpBXaabGzlp
JtLzhItWakcx/mJVR0gETIRLhzaJ3rTru2b4aycKHpWiJviPQfJXgVRBCY5iUDXg
pblyrkGlDbHwjIef1k749Gw3P+O/TGaistdPsnlgpj92G7g77u/RznFaWvOpJQ9M
1kPRbSB1Hc40laKi5tYKsyFdFAwPtDeF+be17kaGBz4gRXLgIpMybmikDWvgNBMQ
GmUqC5P9H+ftFDAGRz8vbp7KZ7L3zdntSnn3t4agDqzwvQmRXV/kv0nhj361g1KN
sGElOHerfJ5nWUxZlUcSD8j7sZzuE+Y/NVVDhDBMbhQR2MWyuOSFtL0VLQx+oHHc
0iVnPXKQxwSCZExaadqqQnjhKPK5pSIeZVkFcwiMxhO02O9M+WpAs/RqzeP0/rWP
NHNG+vv+28ZRghhfahCieHaap5DatSoy10tZOYMGD4GOwQoab2VnoKIZT4IyiAUy
R1ADGaR0kxaUql/sJIUXQDxECoL9lcaTuqm/u2Zgnx/VKley8xPFOZ1CaZEke8fU
FHvRI6Ofgx3Q+dcXdlzpC/NbNYvvmFbBHZRKy4W/7toERA73nGvaQmvIHE+rDxMf
ik3fWllORioP1/o6JBbtCuRStwdbpr5FAUisv7DoFHdvRrljHdhPQoFmgx+WDuCE
HMBq7H6cpBjPqYg6evQ/Q3nCuswETozQxZqXWWLjbk/ex91tCYj+Gs2MwD1LgogO
k08y/ZkeV1VFav2y9o/5Z9lGmop8VlXDFkjClNSZRLbfbptXbv9mhkD+/oproimY
1c32ah+bteC6l3pUrHp6OLLKDGcgR2w0fDQOcxMkNsb1lnYZv8cZFTZmjF0VaoVx
FtPWejsjmC9RJPt2Q7zn0Z2LlqdkEoHcwid28x/vj2XiXexyaMecIXsCa4LYuABo
zRG8H80Pf1LT07EszBz+l7adpn7P1+YjelMX5ydRTHNHZGbGbNMk4XFuvNJxvBoe
dsm1aJ3DSPUEfVrrgOQGU3zs8GwNlaMQVTf0YSb0Xi58NtxlhmmHox14FNwK6cWD
zvLDhwfAkQOgOQG46A1bdczFUQRj7cLs6QgEMnXpNK2jkSvLqm5UbNJlpvB0O4Qj
Axj2P3+1lX/KNuE3iRNaxYDt9fq+NXq8LlmDwCpktkvOS6YyA+YpSL7M4kglKRK6
oqXXYN1dwi7MZpzRGzQ+axzotbUXZoGSJwDzcLmpaXovCReWuBLX0P1nDg9TQb8J
tHA2Q3Rq5C8R7CCZYLRw6koezPgrHytxxCrLiXQBzMj85uNEFHfUX6FB4te5VclA
m4FkGkEzhbjof0csTUDwny/zfgPomRAzReRPyxRCoXtzK/3/Pgwvs9JbF6Hp0WyQ
OoVB+Fn9WRsEaSABewpQD935ZwNXP/B4+Aa7yZWN2wx5WbLouVap8pTPomWa02AE
tlbXcJzs3ZVEofTd0m/SjFYrC2qOxw2JBrYc7IrEUkR20qPIHOxgeMGHASriSFq2
Qv5eXgts8nzBpIIE+XUM+jweMjhzhN0jGGHQmdvhaFl4qwDiEwr3llpJAtxpuy66
Q8BsCRlpfygEvSU2L6y8fB50CQdXjZo6YhCFlaUkENPfzD9UxaD/WwnLhQXQJsz6
yfCodr1tlRMEp+b99B+BtBi8haDw0WkmwzkHhw+S5mtCFXt/3UvY5rcJElfceqBK
QrYCh/QXibBgGnn2mhtGXxu2PuxY7Jp98thv5OkCCIkvErIYksm/UE9QswCvN39O
kZATn9ooJB68riiNVI0m7GKuNIGyO89WRPaNzS2h8zbNMIZachacSTmQqNGf7Ehr
W1RMYRS6vVByM89jf9fwcUHIDkEV2KGRR30ZXXw5p6wAty1VnhSEYLGvwXkm8Kh+
4EUN7EWrkYNRDxdfLnBVKXec6W8T4zT0e5wPWALe66MS4uHE/Pi6x+K8qMRMauzP
m/fIx0uTfx+MIL9PVK6jX+uzXehVxREv+67jNh53J1qSlnHcA3k7+joZaF95b6l/
+DO5h9fjH6borDymiYrY9ryjUKl936/0Xm78tJEXRcYUbRdQ3zIjTXzpSAAYKlRp
UVKf8tMG9c59O7q5FbVfPYxDYEXLzgJFDZICyDEOxsATFMoZwsK6Sv1Th38BwYO+
Fx24ZvXMJvZPeLEkoCixkSyYhK2RMzW4UOoLiNbysEJqni/J3BdyiaiJZg62wSyr
TLfUg+XxnMfrydbe2wJou7vgtVHjE9miU/2S42UyKrkjZnDZF+7II0oV3VZWbzhC
NR6Y1VI4zlDNwxlozMPAb7aZ6QKgTwlkuAv/Qe/hEr2W34bYGy0c2wNw0nNm6o3C
Mh391sBPTiK9N5Y+IvJUAxj4NKi+BXrC7a/mEt5w0x7Vh8jJ3cG2lnSohWWcHpdr
7S899mx1WQRMhToUNEu7Mujs5ayNKDnUhQ8yY6sQ587NEqQafEscI+qy07x634p5
AG1cTkYd03vYSFgBT++Q4gG59BrgSuduD/GxCmpRIP7qAkifbxbr1yhmtLpIc2On
iLpXO8Mcg8yhdteCdTwvyzCyHqGIiNOUs9ntPJGKS6b6oFe3lFlJq/5PIxFSZhsq
Awt1fSWUAslc72T6mqKpTlhH+UA4JttKn1hi+/xOPV2mw7KL4cmqOGpYPksohp1A
9FvEAhQdP9oc9nvNV9B0lUeVjevUrw5RuuRV5KlHOTHhkHsLIbZCelSP4lSPRHC3
6haFpG4ickVDvAagnhQZwTodVZwUutz7sGeD2ibtFBitzCE9x7wEza1qPW6Na0e6
UWqIcowWmzxyTc6DBJkE1/9TehW8nihpB9z6GHYd9rTVh5QFdGXXO0GzwBiv3cHB
TLoPry96DyZ06fLgSyx28PA8CMQJQuHQPknvcZHw6vKxWH/+CnHzAUTuoxl40k4G
wos/bIwvJyViKSXS7dsf3gAkR2L1Te49HdnhkBkjc8fEwRo1dsHjW9dxZPt3x63f
QNkFetRivOJ4XcEv7W6OTB7SAHD8a7GLUX38a6FZ1mN/yD/n1qfuIizTYO9GG4C5
zkkZyIvRuGh2W05IXj+6JN5618LLmVOF6fTvXE7zyJt+lxTA7eyTq9HYuDcdvx1C
ZVb6A0dwYWipKHETDXU0pVinegiAqHN53zuC3OUK3HFKWe24+ndMsLsa2FQhhlwX
DPXgvBm52Usnlvup0XIXUqINpu+UBtAtODG+m1rajCg9gw3EEYRdmgz8ql+TsMYI
swhSNBJJMtz2IbQoxXU4e4y96gw+eLKBJIkjS6TCBOE6WRgIL/GO86F3zIw3yfGF
2wgfJRg27KYo6gBAsjzDKXpuyxXe5pnTV/Z+XDfclwUPDleccVjsQyTEiZH0bcM5
a176zqO/GLU4yigwImZW6VvyPB9xFUg97PDT95Q/1IOSsLqUBgO8ozHpvoKZNif7
0OItCkJXP9cau2ItWDgOD/kCYy6f1ZgTKlLIpl+WQD4ul2Lfpt6NtCIC5NITAwIf
ZWCNxGxXDYA7XEd2z7nSRi6+1yVFCM1/w6myNo04da2PohEIVAh2QRqIOwJqMaia
JlKDFT/WMKLrSCQceymJkCLBfNDOzHS32A4VeF3OffnvWsX7pizargTkrVeytfhk
3yMp+3BWS3DDe3zi4vhi0RTaf/e0FhrzjHaGN0AS5kNcozYZ4MuGe6fXhU/n1rbO
CHBFcQrJ46lWI0HwlNa4+8JhsHZCjlHtFdtFteVW0WnHkzve9rY9318QT/rSArOf
BcHFeTniQjO4rxF2oytx2S9r4RqfCEoQ3UI+CGrAqUZYYfUPXNZUfo3DiasvmH9B
StV/hbhLu6svUSmxHxrMAYZpSq+dQGd9FIjkNv1t10cBLN6fmWdsdUoS4nc3YbU/
aqbJGbuU/tY7ugdrNJQMcM7k743WleiGS4rofV/WJX949LGOvhurii1L4VD4q0BR
gALc1+GLHDO6X533DJ2aOTHZyE5AhvIKVKODoXPdOSSKJgQK8vdJm2Y6gy1L4r4V
LL3YGEgNhWzLBGll5V+b++pOCUqWDqFTWDMhA/L/uhHk+VYWcHCcpKKtP34FUSPL
kZZKGfqJmMts/scIXlFBIsqUM3lXF8918ugyvgk0wRlgzf+GYnFTOQQjWv+cMiz9
+8SxQiHYLOB4xoljPqcuK5F3kX/64BOgrkPuNriX5KB4LaIgzOdp3ldio3H135n3
mvKGe16sr9J6U6bh/AvqmEsEdyOWQweGCpmId5JeLFfCIhAUghBUX/oNQ50xgWTz
6t6OHvICHb/v5bHuBOT58F4f0sUJjROWyMu5Ff5Y2ax4nX3TsEQOa7tlQDo2ukWB
64FXWQN7/2L7aLUT/gdd3Qrj5VZSideAoOVRmG2T+6RRfL59Mv42ompFfYAjBQBJ
tXq0zSAhnV8ZR5Y6IfzKjMnpwd/CcEEBgllUMIZMKhMHBoD6z8Rb+cf6zjEFlyl/
Ug8SXxtJKWbQC7ih4clVOnuvRSvNtdFoyCfIiQWZbTOrrIbC9gEUiV1+QAo2InO3
gOsyvYfcVdgiUJDLKh+KYZX4KfR5MNHx7K6iUEKQKR9I4zCxcs0MYMZIOMXP6dRf
K6F9/Gjm4Ti5tTEagTfz4OjbuuDZNjqS5nRGQisqcMTpRFjr9oPYuxtiuf6o8/8B
fZRcY/2Qh57pEhZb0KJTwF675N5fegI8RCxovEDJPBu5DTQPz2FiYL8Jt68a4HQG
avdD6j7uQrBkbZ51dogKnR+J7EflX6Rb6jQO2ZJJY4h3xlQe5D0yvKm+Nwg/vDYC
Q63XpLcBjWGyfVJqDcpZSb0qUyoyaIVwlb+Q3jgRCsyvQmiXAYkOb7Y2qEU0Amlc
B76W3FHiRwezxIzzs70GpHpZ1cWL4qlYDHOz88lTz5LVkhWzXo9YlQkxErBrI2Uq
krcIWWUMBZxo1yrYs1UFqE54WeVElpaB4iF9/s+2o9Ms8p/crjQlOYiHniZMLSnd
DUgZkpfF5zWLVpyIYHhWPYK649x5oe2/kntR2jJ4xwcYONLFoaVUA6AOYSDFQF/e
LyIcTyX0nP1O6AjQKaGc8GBNx+SYR3MSPiVVvBR46fznB00/BiuLV6RPZSPUtmIT
gMcA504HvXM2cPHT3SWoXWr9lwXaJg5YNC43ewm4ZSVGg/SXsOmpsij0SfEFvc5y
ejDf4BTa0PZnjzhMpKIgLVUi6QLnZGjUK43kN7nj4Uz1dU59kqL77fOQDUMvtk6E
38lK8mcVdUk1hB16ol4ZSx8EBBDDNlJsOwBOphU4IPGcZYwnvtBHOmFFWvjKnd0w
aYqr1OB20jMAyBaoaW7bn50TahhJ8g3j/dnZjuUKanASdMkfuYv1YRXX/rCacU1g
xP1RppsTX0tDoB853OkSFgAiK5EUhGH1YDj6RHfJt2b0UCKTRYcfmCb8SMYjy3Dl
hFM6IIE7UvU1k6q3/4qBYCaDK2oE/TBIdfU3QQ6WExpLmf6Wv+e3M4TiaLxzRaHe
EYbDT6ucdfKNKu1HTGBirLMMcW8lUWruUV5W10C66qKfxU9bDkfbRSfIXP/73Ro7
EhbIcmZJ8yIh6VEqnjaOOi54fSMw66YUqEQ6qMrA5/x217LScA18JGQTOcNd4VpN
Pozrs6hUjCHwx73OkHy7msKt/VoBnuY2+OsMwVzymV+BJGi9+5U6GZjD8EhNJAar
UkGK+g56FdvH2xazaS8VyFwScEBmqm0rPc091Th2h+Ig2W5vUz+REsZIExWhtavs
5PV1EIs3SRl8GpoHAQNOkBp4fcaj4S3BNZx1fTzZLufC8+8PjQwKs12sSgY22yz/
FdpGNDk0b+djce7n8w9MERsFkk9O67uy/Q5Kyu6rC7f+zykrShwqlKm99PWwChZZ
T9LAEGKZLWzqtIC7cPUoiMpX43uH9G4QypiFAD5k7cG85tuiXXTO9EdF7rbPFetp
bM5hoTWQZZUUgC1JIB0UoRGcB1hRIp6Upw2nr+cofhuMwJ1vFhtMQO4ZsIUhREj8
cVC97Cu4iJggSwkpaLD/jr2yUPKCFiCGEJLpLEpdHaFpivCmfkLSM6zH4jem93Wm
tYUVo1F94c+grP/OtTYt0LnDyrC63EQUjbnlSQ1YSl089E+3bKAGMgop6ZuVBBQZ
yxnDTw7j+WWNYcMcb+LXH0LsXOYJ9c06j7ycTOxXcTBEXSeJKktMSNaIkr4SoNRJ
O6fADLuwCJjEubgKrbRtIjAv+cdUFC8B6oZKQJbdKdP/cvW09ciNew4TRfCHwemO
QQ7A3gBW6x7d2k0DkDGUrd1lIlQwIi42gkgQ5LrwY9aVd/BsZ6tCjxhi8nwb8V/V
p2q2Sb+Bq3HtYRAJqaeVXx7c8iJL0lyfxZsEM7LvtxbLLbUIc6zCOvXDi8RS0LUY
14EricSCfu1fx6pqW7WO50bHCLToTTBeO6nU2zTdB9Nt0cyf4Vw8kI6Vu8l5kpS1
+oVGqlbC3+RwVtxvzBBH/4tGrqsKI5E6m5iclkX3aVKI2bVfYPIdNX9r5YBuzzZK
BzU3dn4YKBxp6W3bCSvPSJsHHPRUxA4X8nC3NpCOnJ0OeO78p7NQYlfh1cvzMZlr
T15mYJ65jZ8PTP8MckgwdYrPOZK30OsXdToanUp6lX+hMrF3ZKcJm6HCMVx8xfQk
RVeRB2RbU5Pt674U1iEFGyW4WSoHNv4uE+evSoVNiZmzvU3DFBZtSdNZRg9qOFe1
BvL6v0uLVXbb18k3lC2gkEIc3QRQaSZ4I7iYH5w4s03lTJM8D5NWAn9BLvJgifcC
rTQsKFXXg8drIH4jsmAiwKXL45XxlLxhd+tX1uzoppVN/E1IJ4Di6A9kxxYlO2xJ
T/yEw91WUAIMyi6aHrS+cCnLOXEKIAIDXv0bpGuNyyUE6ONrSWplk91Z/ZRS9K2D
qQahqzlFqo4xV2A9B42nExz8asepClRcL8lWG3uocKjRJ5qhtkvpGph+chslJeiA
U1fFGlOiMPW0D07ucW9kU+PwL/WNkeNSCazRvo7s29A3iQGmu8Afn9wFbY82n1tF
biY4gaHlJTmzpSBFVZYigLBSzeAXOgNMkKnNapgIyAnyUwdbhMnT4d7b8ezMvLHy
/wdKb7yi2RzCwXqIIHD7vKFb08+6tUc0rZfZpuAvKEQvLyUuqobtuwnnqyKKzlid
5Okm7MBsYwH149HgwEJLFhtOH/J31VpAxkN6SSc3HQdGztb/1faiiL2QlL4i4pKy
otVlK2rwrOAxyzGjL4crEVC7eYxzeJR078ih6EgSQxP/Oe52lVuS88/y4CZkEjTM
cHnBM9vZjxb/GLPcnZS0bDluM9vt7Tnbefjt1CN/M3zqpWL0Vn+q0/IvdHh2rzJT
DKq8KO4PevLsa+/g8157ZOnxuEGHWlpKw4YtfX4XIsP3l5u3cACRoNwOiO2J5CEZ
zXs0zGkJ83tS67G8iO1IFeKyu9p2kxxSAWZcKxuX+E6tQal+xUK7yizkkBcSDVn5
uCEp2pmlJzg8LCmPj4pQ1N4HhEPjVrC5l6tccFT2alA28MzuhhWM+nYMwh/+34kl
II6JodleNTAEcPGurpk0ApX5EJ/QcgeqRJfubNKkAD3buhUktpkE7cEvN8FUqRK+
0s9F2fiiVW0oojfR12+Blap5CiRmmG1RR6AgKB5zfSHLf6EA7w8Uv42w/Boi49/X
IM0wDd/BMDTj10wZq+SfH3CWAp/93gNqxYnRFsZF94dugXJ0sK2ntIO5TFJOMP1F
CZToO0FylMnssIGNMHgLFqoOw49Rk6bqG6jpRkypllCyvyLMlpKlaWlkl/ABhyR6
scYjTFe/0zOiLp+4PZIv6va9gZpJqd5iflUyYk/BSG+xalz5uiQU/XdnLiGUhVwI
yy7ufMNXVRsSbpiQj3+Dg+Jis66YcP0ZItgK2DmaJz18M8Z6gJ6rf8k1h3FnsgIe
+XGo8YolQBnnawGiZs+0VJo5EXuY4DhrpTDw53z5WygUbPsXzIQtn49SJVO++Tzw
a5Djz3g5I0zce4HccEUm0ZGtHEO8BbQWmSQguoqzjC6NHD6LjdiwPZPkT1lE0GOp
jAudDYxrc4XKRfi2gsgRSRLd/MhEx/swM+fSVa/xe9umMk6wlON+CXdJcAt1CvYl
UKUYJppHEg6EB3KQkkUp7SJSI1Pn6HT/U//tYVoqdW1tne5g5/hiPRI2aT3SUit6
QEx7jdzRwARobAqDsQlVRSvQcOP3sm861CnZXDQAnpnAkZ3HyXhlvcyPHnjUi4Tx
sq5VKmV5VmUVdN/EGJ1fAfLdTZUoMsgG+X0EgXuC7earqdhUgDt36wc2F+6jnlos
WOpr6U5DYbTgV/r7Y6YLyvwa+CgmYnh9ejBH2Rg/7k0A9oDkLZnFr6uLbfTfB9qR
jIXU42DIFXuND4sKNX95xhl4iXaztc6GUvQwbA7jPWyqKlhsbG9oOKFvRyu6eSij
BgmbF7OiisekrKGMGeG5S8fhScBMoJ/k6ZuYmHSO0sNDedtosNHFLbu2ofTTTwWA
O/QSkFPzNSPr59kQvZ9WgY/E/EiMe850zABXymqFFK3FhA400zfNHDKxPtyUf0Rb
S82l3Ry3kyApcEH5z44G8epa+mjPqbwD5SQRKuIVAM545SP4gfzUojd7NwznoHoj
rDMewiWtZ6CtxGlDpemILmncnGnZj41H+fXh1RfMKbi69SZERlKXzNk4ZCt39grT
YpAC3z9p4JOPMidt8bLTyJoZxqjZ00W9MWScYgfIy6Wr7eQ53chNTWoYjJBVd+i2
U8Xixk8S4pl1jCcX78/cocwnjEB7nHW6CadUvcjgwhW6LYt8BjGFz5Qu93PXvcTI
ZS+i+3mHXADucXGt85IovoILI0WBQBX+YldhM6mDR/6IAEAt8vB0fQISG46dKuOo
JR4aIxZU7T+AfsiZklKw29hvPZimlUw74yH1Hah67Vsj1FRmxL/bIBLIOBwowK4O
CVMNsqGQy9x49PNzM9l/sizmSHy/5hdJvBxqMUczyQa37OHo4Fn8QkeYv8ABfGLs
DBPFhh8j2VepofMtj9By6pgjL1t8784iCJ1ZakOc6D/Jb8klWijSYwk+1v4tv6NF
gdGJDXei/CTjlD0L+85wXBVr9B1LTKKtvlOJOoB2inwNQwnDQHvZ59hsIZgls4Tn
kIbzXWyC3egVeghw1cv/hW1dlc4s4Rs1A9Cw8jgChjHudTg3p5VQT3QzsAUzPzwS
7A5mo+eUYF3MLP4YLu9zvrqbT3AqHS2ulSzki7HJHgwOmKHKGXyKQzmxdEDsRzVh
vCzlyEaz4UJDmCxBW1L8EVxsstJVUrcAxUe1mrJFqKVGPN0zUKQZ2KnGbcQtkp0K
5YOa6bXdLNbiJXn2Swx4izQ30AltjHqxIbP5Zdtg4Noi5Vz8ZqQp2qAs73GAbPgE
y/n0jpx2GlBRbe9BuRHW0TRdWHDkOnHQjt3X65Zou3GSBxMKfWO/pUzHibxhkpIL
1Xudgdghyl51fMQrq+wZhOhBrTRPxJZVRVwXwdMFKJVI5XkHnHgymwMxMPbmOUtv
/Ny00amxQmBvp5xAzcJa65URR0Po424UzrNQPuiysmAHoUAcRzQK0hu0FV/bQvOm
sAnEOSBrKlrzN4YT2J0z6+hNPOUkJ3p++AjpApXo9K3paLRUFeRxlO3PQY4Ro4cu
uiV7p8kZaBl5GAcD8Rk1nwzmUbQc8O155H3E527XBGkabMf4NWPFbkZzOxkPuOZS
m/Dh1PhnBRGjEox4iz55d2ZfMdGnwL5V2rBJZ0rMM5mum88X1Fln/c1rl+y4B7ci
7eKb0I/wMwd/ihxdBijuc3Ggn+Xu1btDAuhAi0Dkcm7GJZG7SsS+2QG+jtFpuV8C
vcTkIqxtE49WOfofZHCG7uMqm1/dMWs1NCGeD10Km3mUCdmxhNqwQn/S3m7j6fy5
z6ifTds/tXNtbFFlWHbdl6y9KndX40ej95TGjSAKKYRtT0wUZMQjJKwnRbYxvQpQ
d7U5tOdCMvszMg6ZD5Y4mwKcF2POnXkbXGD+XrX3vRRvk87zYIjL9TbXIL9TvuWF
Q2LtH/SUofGkO0gszjeCf8GW41yy9r0QDvMApvXM2emYLDyI+Qv8soZsYgcCY6ZY
TLg1nffM4z99o3O5G8L3Qu7gZ/BAQNGL0Q6wF6ZRsOPIyqNe2Vsn9QHDkJ/9j2bv
bXc5ONNlDuPUwv7KIp72PHNjbOr2q6mkJTmt3dJtGNfdy/rPaD0uET5h6eNLmcZW
7lr4jfUonI3AHWnFskoXg5mYcvIUbtK4DVdL4mKsbxMPFQ83T5T4F4Gmr88fs89I
YW7F1TdFKwI4874kUjOfIPvBJGLYZO9nmiMRG1bqtNREwjcfawqgS/GTPpe7Vz73
rjhI/WJwdt0G0rJn06d8usxkN1sovqz25ZIKvJc81Qwu+9Im1AKBT/K0J2gcjkQB
bKHW4MjW53v0T6QbBWxBUdpTxespgYcfU4FW5wXHJ5kqERSnM4366A8ZsMuGq+h8
XO0OhzIShTyV0xzYP6EUXK/aOcD5LBZJ2L+6/JyItUTfHcvv4DErYgb4kxmZg0ZS
wHLN2s9U1pUBRu2aEjUKOpGnlWbxbn0a6GoupVskv9cWwNJQvcpIKn81+SpVvIw5
WtmD0Hf9vuwmPLfWGIdqLCOhH+iQOSGFLeX0dqJ+iGVBqZ+k3JMu3XeShBCDYYFB
Or8hWp4vEg+ta7oT5eT8Mubdemwr1O1r6Cvtu2El1bk2+X7X9rxEFLJUzt4pTAvx
/05DStDU3qq3Ec6wYa89BWjU2H7QOPWFcb46RMSN/l/06HXkh/QttM8/4PikoiKB
dq7dgn5NIm6k+7GEIlE4W4fcpZ/63rcSWNbUjcCLF002KYRmOVO/g+QiC5WcO6Nl
VtrUP9WOQlQJ8mbI1F6a7pc4JuRalwnZ43v+1UCYJ6a9yrDD+eFQOpBSR3s0iYl7
de33SwHuxY20tqaLBeksInYgzWaPcJwHkXY6Yno8BO9kC/iQ6rdqFl421/g9BMDp
VKqPWsSUk27FOLgNoOi7KCLNMK1CMOJuUjFlCpsQ1O/vJYvOdUtNeG67rh+yvBaj
PIqZScgMP4qKtONI0Y7GOrOGYE14tMSA2lxkwX5TshmbSNFCrUZJ9JhAconxdG0R
7QVYWfAKJYBL/5miC1pcT9PHb5mkjcouUTqYyE0LAtAiqF/i1RoZ0D3BKAw4aZwI
GTpMy7cmAFEEzwONFPClBUu+swfqXq5aWJRMahLRUwymWx3kdkF4z6c3xfbgyd+t
eTBA1pqQ7Y5hAoOZbyP1hVLRDoPJ5cU5/zQACzErdJXBcJ4K9+j+Aptehz96H/Fd
ewYZxwVWt0xpS6jVDL49OD1zJxQMA6tE2UaLa9xMrqJCAuM7IHUsTKWTC1VhvGvd
vUyxDTuQSu9M//jDCrmid6mx7nHoFf/jf59fqIzWlbemmmeCbP7qFDdzjqVadE9m
yLSUvGkg0B4YUU2QCA1jX7h5k44kFztZi0CuziltRI5ZWE5gEKXGVK+ih4ljY0F4
CVcNUhISQx/TPyCpkQWG6K/EHu9Xn2v6zdTXDy7cwgFSEkGeOh0TFSTrKh0sG4Hu
jXg9HQCjQyzzOYvldNp90vz4iBCziA6EGlgY0Uf1p0h8DmjAgih60Z5SMytgL/9Z
ue2BwlBiYpQw7IJHTChwoWY3D+oD8RMj36JrvQPD+1iTw9lm9N9llWUEsxMC2EfL
yKde8eFt+5cMZpyM7uLYt74tH/NxzUR4Y7wkNHmiB8j8fs5PwF7S39a7nJ+pJw+4
bkC57ezsbtQgN0JFTFdUO1VqIKsi4Id+yNfsATm0iYJTe6GWYekiAmhNofi0YfxW
EZ8KX1YM6vnvcnxuCUzgFHN/A7ku+I9sQT3H0GaE9qNAn3CYsQR1TNbqFyLovvXz
XctpUdyKY2GartstIqnYL3ZNBpkFa8X/zFxH1NWGvAkwK0uD6j0fpua3SABdISid
MjNZK7MKJX0rOwbi8OMLZXUiunzv2Z4drQihtnTRk2h5XJKCfjQ3SxJ/ilngjLJJ
VkOajGW3582l2tkEPF/Y0mmKDWTN9EtxEL6VGIt9bhnMb5OZvWnVfzLw9o+VJ3LT
zkb02LqsYMDz7nwO+AmWxz7byAv7AVG8wDyS+2CvYLrzItpDqUWY1bTiJVMzvRHA
LeXTg9tXNag3hTcwuTZ04H3au4fBUxh0l/EAgNZVFmiZKbSE9M6vhVclV4t0odqt
R4Rts5pvuguxBKD1hebnsrl4qnbsFTePVfjhJbFweYLZ5caNyG+rLaA4fWmeY9mt
N15x1nGTvEMefCVCNUkdfkrRrV1n+MldWOYS6dy5QLnHxARhKHXAYc74OJWK1IUw
k4goGGRu3Em5Rs7Qf/1tRMdW/gvu3/YishRI+MKNNePenFO/A26WqyS1iTKLZcf6
LVrDKeli19MNZEMYXevou5tUD10+c1m6gTDym2XSZwFb232opUo5YW7tBGSHqM84
HJe3ZGaeLq7YyCeumktuy7oQC0yDrgcNNduEWeSro1QfAKcC/z1yxsTUcX2foYXH
67AVSBL5+RnDG+1iOjc/aAtBE0Gbk7BceK9l4PMrhhyQ99DjBv5sZP956yOHES86
NPVQ5vp0IHZG7fcNp5KR6MKciBGzcgMPFd2BQsqFo0I/A9GrzQD2WFY8EhyMNQd5
XTT7hscT2dvUmMFnk8Sj/WczTod24QdlYvAXHQ4kuwoRJUAJLmsFvdZo+vWgRQri
SKtc2oK8E89smQJy9LxdvNlPBKb5w877BfPbZan+WiOmWsj8V5YD8ZWJIKPIfcxP
iqH1a6DdLyf72zSnVp5ijZ0k+t05Rrdt8jtfoYEpnV6I3Jv3qhVy8ZKXxSGvGvWQ
iD4MiRJehJq8WpzT+0VVi+fV6jwXzolISVwJsTQiAiVsN7+TbxHwPvGehKCqfYsx
ystPTXaepJJxSEQoE5MTg33wAMz6VOPvWrs/1oxTqjwE9OZMazijr79eDMVSM3qq
c9Aj3UpxnQC5Adz0QHSlD8i4Ct7W77Sz6kAuoYFej75o7jpB0jhpI2seFgKtRtQr
YA+dM2SCcL4a57HT8oeFDYXUJ+i6ZqFIxfwLghj6DMQ3ITnsRXgMTp7cXBw0kFHd
FXRKg0Sw+hoE9VLM+hlybk7+CVfV3P07+PjtggWyCuuoqZXQufd467E+py2rjKUG
Ri7+5MXoKmBsZvHsY+c0z4Zqlyv3JTYqv62EaVwPJcaFT7Ji3G/3ar2tI9LrIXXw
sCfikf/Yqcb9c8rQh7T/OF1yu6HbGnVNzra8+DshrmT92vLK84bJl41o37ZFk79n
NCHn/OgqU9WhdWIsnKE096vxnUjrgWfdLAB3rgZDUgSLgYgpXFz/zEsY3ULR7D8M
0EI8DYJCjlI89bznh1XoCvlgEPk3r+9cr+PhyExhDmlWyl8n/wSS5+Ozd5nJN/NK
vreHW5vu26RL1xl4pXBvgVEbFmDefymVczWaIp3CWQvSuniMsc5mDb5lGrwAqn39
bRVECKxmVvoaurWetyOO617gyhyYDPqs3lVku51uVOC/c7Rsfh5/u3gJEgZjwUqJ
rqy7zoS3kpqBeZ4nWVW3uPVS/GLRTLV0Q1mMeZdwustZACJxos6oYNVSrrBBPBec
176zyv8sGHoMYPlOGvjnA642Ld2sm0RlrncIkwBJxmar8RHK3wkWiMmxIv8TZmXi
DD1CtRF3uTumeRK5DRcehxmMran+oHTeZ3T7KRMS8T7YKQgyHgVIkocW9XI8esIv
i+j/bAfPzOzkBKIr1JBjKRfmaBZDUa2QBbOrxxZdIualowjk3pTTZl9EaCpaBW4R
rXQX1+1ot8Sm/js7biuJ3NfZiBvyngTRIgI+COt3CZ4aD+Cv01sZTE7oEbCHfJWR
662vTNs8TiF93v4JWR7jNVBfcVao+sKVjraiJkkkz2lXpYouCxeWsQzIfxKrUXxB
Vzb2xsLotNfi2khYx7dDgwdYkFy1oKr+UCz8f0Oje3MrZMfMbbyeZstnFTouNkPF
Q6yUT+dmVzVRqymVMcztHU6Houn8Eh3VuYu7BY0q7SMBUfc3H+7m5bwtyFCovgJu
S683nkxGYlIgkhFJNCp5Ib6Wf/OIdj9Yj2v1z7qw51/+C0DbVoI/gJmwp3BmdhUZ
OfFwcjrySKSFaxP1aWdIrT/vpCvMreAHnh7RJA9N/ccFkr7Ytk0LNmavVjlNHpJF
+zYM/aKeIfB+9dI+SWdu3HyIBee/BuUj+X8Bgcr8pLvBIzssBT97H4SOhZMcr0Mc
IcSLjBc65YhHNmqpZfJwl5HqJdkgtbsOJoQruDwhXxMTmgdNsL6FT+qlMOFrjRHT
f+/JzktUE4Zc3vSCPN4dYeVwZHxDtGFYmdJxscpr9CbaMpu2Ar/C/ouC2fuIYFuB
aHDItiR6Wjzd2N2Ug5eL7d5D9LL2O567ZLs584erd5BJ72INAqWzihN6/cxyhTVA
MbtqxYGXp5rLJrkEg/IBfbLa+LCGRAKIg6gYg60AbKZxMjVFbV14OLYg173sXv9h
Q5d1BW3CyusBISUHBA9z/vFW8xQ0wqyJm/0lpcb9GM6lm8gKQHycw5TbFk8h1L70
Dd3WY1e5YyzMInuGxif3w2UskiueKTL8slxKNc4EYVA+Lp1AQtHfz+sEha1WVnZA
5TkKDYh5UD3XYGSykJQ5V0pzo9+l+KBQNGaY+U2xiVsh6yhrKjtMb3/e0awHp6Q6
4bzssVokoYL2tRIgMBK2GOVFC4qZtDGz0KitTS2x/+EWscN6B/ADA2frcxWGD/YS
w1ASmzAnwQ6ObE7uE0TveSA3yERZi3Yf/ycIWfpEPtjDLBLKc4BiIewlZz7CqLP5
4blfEdf8lMV71QgwnkCagt0GU5vSuA6ByAe0OSDEvMwtCAM0VyUpUb3wqg3H2Bxu
VPfxVI0aQSDINhNiMmzHYZbmbzExCcCu2n4Df7PCnrgIz9WuJwB3oyNZ0oJ87q0s
RON08KmpTF7cBkMpVH/FxA9BuZxKWTlrw2mC+2ooj7XrtkZZ3ON8fnki7s05LASR
FOpMK3KOmtLQStU7/CMLwfGutrYVciR6uCx2KD4p6UiFphYaowGyaA2qdTUEiuvh
NnZHwzNiIN7YqWFqyFlvLAj73IBJQa3ZQd0qvnJL2chx6GARckG/VM4a9de1gkvK
dEGhm0TQOs1TWcCS6ltCz4OZ6lNKENoLHVkygOcLlPSwNi3cgmKLeyvAc7AjdR6q
UeCAzaLec992wex/bDiV2t4Ik7uVdLQDqqRbDmXa1DvlrPj+HzRd9HI6JdWxYlrL
PZABn3fT+es55HAvjmv8CQ1QaFwYVRAOsjL+2ZPbPuQ6DHxW+yD5/nI7nx7msNJe
g3WtZfcepXh4fMoMtihRJabSsbUG23jE/mn3n9QJ+Ve0ekNV6KVYztIA5Eo/aIui
lDUUUkv8Ln2WvKvb4bPRrqkwuyQGL0TwiQb+WhnnISQmo9HJk2vfAwWH3VaYMwjg
8clQRM1FWgnQvv6RlfAsEyDs8UE/Ett74Yp3mRmF7/X1CYvFrmHSt9Mt4j/oVQF+
i+Y7yPkD3dHd6y/kZ3pK0Dykf3BR+zBuRik6I0gjXTp559unJjahn9ArMZ4tdSrE
6lnKBVD2nK5p6wbqgmPjiDj5Mkf40b6AQd3pPeCbdhPovesDbjoIuYtWAGQ6sYJt
8UgpfDBclnmls2ti5XZH383pvKXXYqpZMcwpqobNwI/jkL31f1f9+tPk4AZQyM5Y
qGronn3jhBYwM8l1a/7mi9UxgHS6z7EuIqVJJ0Dxe0zuk//6DVzFMFKTqVaYyW/B
eR6nvxp4MIvChPCKjG24HIoEBoSQ7GbLBFZXiL3+OgKAQYxqzzFYL4pRyKKmlDDx
KMcWMvKB0M+GZaptCXxth7n4uiHzUL5Q9pYjUWKjOsetki7Yh2bLg2Hzdh/sG6ta
orUOwrC/Ptxo+i9BOkSbgr9DJdVqjCDPR1o9FBCNnhkiqVZGEkTE19C97WSpfyBQ
BuS7LVI9qLZVSLJ8P2n5kEEzN/MmZQtrW/0BNxQS8ZikqbSPRcGRtlkb6gl3Uj4U
wTbPPo9b1A3ZhyIUgx+mq8ZZhPG3MP+nr2YykVbuFNhnGq+Rf1+GliDmRC9IQI9j
QgfzHsw6ghGmici0gzAixlPRCrBpz4aejFVHyLEPQUnch4/os6HYXLTotnIYr32p
hPjLc3ypvgmLbfu4TRC0CGard6imUYGlkB0qRczIC4ejv/VQT4vATJdISZLj1lEh
3halkWXjFHRPO8aJIWAujWSoC8+KEGye83MxrNRTHhVL52xVO897UhDGlDm2bUrZ
N0AGnGzcYPAm3u/+nQzCkE6aEIqLZn97bpGVO5KYta968qhO2acSLoQnnpNUwaZE
3i6rccX5aUQ96xwqZ57MlJjVuOAjidgCX1mDo2IUO7UDGjLSR0ua/bvcXFBHa5DO
pVr8pbJLMTwFaPs2Lp6DxqXZeZ1OzfY1UDhYeI9N5hatDDEcRyFGze/udCM7mREJ
Fv4OOl6DCBOyTiR7iSK/0GrxfkE5WmV2ZCSWnjDYwq+V4UMs62NxMDzF5NKRp9Ma
cIkgBgWYHRsTkNkDrW81jvCqpntWsu8xSceefEJUMa2WH+2uov6E7TFcKSb8LSlM
HQGH8emmSrAKS/TusZRMXf6YtFKTNpZlkGwwXj7NRpqps/2yiCjDakQZWvygvW8G
rbLv0v3p7J/fX9lnJTMU0SimuAzDUdrSgxuzHUznj9/Vc9kj6cSudejKchvJSuQl
wALMqtmpiMDCi7KGusJb2ARxi4Mt4bIQtw1svmf20HR6PjUHqVqli9LGoc06TxGA
6eUPPtnl909qPrSf4JwZrgfICAi0aUzzPqOoxS+ojxMEjrEjQ8W++37OQSsZBfrg
2y+jpcCtdsnb/kBiybLHuRUcHBqtdV2YRuJyC8KKv9bCUo6CoiIp2gEUkHCa8NXI
jvt7WN6tqdKB4T+bwS/mFu7aEgXlnWEvhPOYpcx6MhweJtSpcyc+nw9RtEv1wK9S
Uyd5zuO1xcXN1cpl+RVKFZclIo7QNgfx2BLBvl5hqbgFzqf7BT4MiwoWWseMyq9m
Bn9Bk8VV52xHVUdZSAiS6vFJhzOI+svB20W2872SqL448xaw98RtngRMUKgCPZSv
8MkMFrZeros9Oxsf4bV8u0tZa05SUlNyNK60SGSvoF3XAJDhav+uC11ZbZA344LF
slG0DHOKHvlzsbFcK1kaqRm492rAB/OaniQdECXKOQrl3sLqMKLrIVTiOTUrUfRC
HV4UlEcerQ1Jfn0fAn5s0m3pQicUxU+A2YrgdtuRg81VnVlZDsqKGeaJ9OeH1Gsd
TKwz+WtiqEokaEE1b/sHdvmGSYFBAPmcTI/m3v712udW8WvjWmAi1LlMTLRhf2MB
9Kz+Fj1E40kVTSTOqxM1cxU5bzHAhZrkB0i0vD2HcFnftN6kB8mdyfxGPbC13vRW
ha16pTJIgSUM+bfDgxyDweq+QZ5izNZM94XpIb4ROfL4HWCWf1iMAKUY2YzY6szg
S8dOFdC5ozJEmZmZ1URfvWFR1JBeB+hC6TDa6zshiWVj2witFu0Ao75K/G5vEEMh
kGwBF9dhPDXddzX5BinR117oSA23AX3Zc3zH0TuOvX5m0JIYdQA90hzKA5pZsVyo
CdnyNwcdy+mqwtJudGaSCIT1afe6xs464SzO/6V4gyoaN8ZObnIKDoPvptb34z1j
mUftoYqPgCAyuRCcPh87Jf2I1LmGalXe7WJAtCM5rkDhAtP/LwRiWrPEmblqxZ+z
WRP0QlBSvSkFHIFnzWmLd6GK8Qq1RIKrPO8aN+KODShpgo0UO8dxckvUvUPIgJ9g
4ah9APUhmSS33JjabrqoBrT4yHkuC45so78btLi0k+D6dBEYfYHiGLH5+DsSVcYz
rQFL33Mfp9fEVfjVG63HHznrC70hqf3xR7xm2P+EkWKIJvNzV1YLg3DWkXviSq4X
XMVjpCoTK8BrEkrF/mx8/0VsgB15729AzMR/AUFi6a2aAgILSioFNwmuAx/n6hI8
WSUeg44Bwb7jUjU6CUcYdryeLeim4DQzjCsbeuDld51AdQ+rJ2mctRXCMcH5UuUH
1TFFm54tf1H9TyHF8r663nvou4iuNHLB1Vhf5hQ9RrDdWrLLFYtT9pIl4wKLoXj/
KcS1LWXe/KLkAk5Xbp1EuIyTCWkl63p0F8E1Hwr3QmTYEFEJKsjWR454wi8hVlz4
TZoM03+ECicokbFGJy/C9BSbRHg4JxMUvVw/rzge0fHkLnzoRDtQjec5ypI+WJPI
OcgJR2tYGjyP2PXoyTu2LAOQpnuiXqY5OUwgwVnpqZRRKcX2q6hxKsxRK5irQv3W
mhQ52DmC/4AKdIZricqf8wi1QWrDo8eEpDDUcyyN4HNaWQ/k0bGNF35/gMkcs0vw
zSQ2FRN8c9IKCWU5RmbEsLsuHaf5QeYBkIRaVSprPIilzDmEOl5S7WSk6Kvm6KbJ
XdQ9wJ9Nxwi9MNUE3WtrkhNLmbrldHVQBXqCTC/c+Z8HhuJ7Iby0XWXsUvSY9VFM
F4616O3Cm8HL+s2jY5Wk5qqV8y/A8r97GsKfxAB0pGUSEjjH39C3jH8FdqcQKF0Y
IGdSXe4VwIJDGxO6SwH7EuvEpKm4396O0SwuJeJEc/aGIgQ4lDPuyTkfuFU2kbAv
rSGSbVMIjf7x0ua8HcOIT7ue/ZPRfE0wo6VbC4o5rmXZ5H9PbRQz4hMtax445f8o
u4HpzWtwI97cxL3O2p2Hl7OMlUnMlawo5ooiY/OCGD0K+PIHWuzmXit8YDyVjPDN
fNmm3hCYEaBrEfMdR2cyB37MRgyBbmZwS1ZhiVJETX7Wbb++pANHhW/lOLXSp5Jl
fFECkfMrtXa5WREibHtQHWM+FDSk2zMOlG/1vDGWCdVzVd1oR0CCjMAQ/6e8iF0V
UmzWC0b4f6z2uT/ltbjZStS2YvavqwFs3AokiyEJrwyaxi2j+Yzp3b6xxGeig+3K
/AluufBdEjJOi94Ear7JGlj87AOksZuivtwkJqpdWyuENQoadOO36uox+bfj5vd0
sSm4EQdyLIfQ18Zc5l5aA82b1Lf+Xy4F417WC41vzlOXbQOg+W0MTeuTB9g4hg56
1Aw0323tzQPsVDW1FKv/1BsMgCe7gm14ERzHGHNM08mKpNmpUXt79weJNenf6Avb
Gc6LC7J33pav4SahzS5p+80kbIiB/mJPYMxWZqoMLWfeHa2u7+PG3RnLtpFEEKx1
BLbQ87TAjvzCnFKu/dYN0LeEzzqEYANFIEXUURlzwqEC11zs2A7l4zTE1azD0sDB
IEMtTJdPhNzVR+w4oW3QV88W6+QHdgF8W5b4jflea4WDjhEp4bPweFOqZL0eft64
Ka7EEVOHecTnYujad5aLhBWvGG6vWOlceEzfRa5EfE7UEVentEdBLdkzlm3z+ddv
UOfbS3+AOrwDEWvNh8lu93J1ih+otpmFFmJtHtKvSqzwHE/IA/t8wQ/pE1TFG6C3
6vhy5qQP4F8pfPHypkC751pHGows7S3Ij7SqXqgRSiwcH38mQbE8s3OUTPVlb+GD
iaGNg5qBaF3p3bvDGwd/spuGy2fKT96yoAX/KwuVc1EBG/XQowE+qW8evDOmcTmK
bpwvZ5vPs8m5elMF4OtK3+G07m3Zlk58SHZRVem/Wxp+nltnlECUIjlgP9dUJezH
H1kQnGMQMCknCHv1m5qCZhiREJiHQlW9lSjjM3HtewkEoUJWfOVmal64QRwdl+u9
CbXVoCNvWaWjCkSWQXGTwUsOY2COczhqjSy0dm4V4QDPk4vY3ftE5GxWuFBcxoHR
JMmFRWRPnkVPW1Lms4HLlIDhT4kciUtCxW8tWubRfXqgUP7vzTZRGhaA8GSPdJc+
mYFeBsToQiaMCZ/j7Z5oB+qfUICP72sZleHoi9hRWhZHgsdngDFhbYQ0nZcAMHIn
RcCFWea6NFVXbvSXpSLLDQywOy2qK907SJ18icOxu4yJyZmn8lCk6TfvdhyzIFP+
saIVmaPkae/yzpTO8sdV9lYY0FDmNwh1YqN8oSvRmDoP5XYvhvRAoqVRArcdP6/Z
cOGDddAipZ1QLjH4yfAkSxDY/JehXd5YwcKSMMVvzqzcX5RPyvUI6fcmHjF7EEUi
AV8iz4h3kVof5dID7wE3G7MgbKEPrVJwFItYUZpgGCH2NPPQ8tBqh1SThja8M5zz
+taQrUNFZVLB9JzgkH3Zovrz8DhAQrBrUVcS3NAfmyYkV0V3atYuGdwWQruoRQoA
ikBFVf32dytdNe/kL3KKm3dpfq2wPDDBqksiCJAnhkP090iNWlspbsedJ11xeW0Q
B7448sE1jV3ZdIXbw/vj2XjBJqxUZ0gZ0EK4SyJE/XljDnbvpbM/GR1ru54miGaL
AUnf3HlzKHPpbAyKmADA/LX35WTdL/MLi2wwzI+Invnj5dEo/+E+CB4qAaQ5wt5K
5z5yK8JZ5vAlqhfvd/unilSGd3y2kgC7BTc9+p9CMoLegokgKWgP3fRhIMFddMHG
vBDBAVgPs6B24mUUf6vgXOrLDYT6fMaE8YIqCwCVZwvvr65nCo9+TYiApOMeXRuM
M37Eu+0l5L5K1W1d2y8c1QTdgUOMXKP1UHUjCr+kvmiicwHg1rXlwItiGUIF1QDF
EBjk+WOaa5HfNkZM3dtLNYbNt59LnH945G3PlIXmsf0B+9djL0+OGvtlMltdBAbR
hb6tD3195T9d5eTkvqCt+vT92hKA6IRLQxp8tKIFd8lcnxEGam9Kk1RifpLww6Wy
evhvquo0XgedHzfAezRXy/gT6CQ3cyhZx2SzIv2JNtTpbW7U5hwAI/e6vIu/OK1J
JmpzWBKAhuNNN1Gu9ZXr2UYX5vPEKUuECRptgVbh4mfA1GmmLULNw19PCCUNTk0Y
B7e1OVcHfD4O6CwVPzlEJPLumABOoD/cL/i2x3w6BhVZW2BM3/2vGctgEKZWuNC4
WVdJMPn7GBh+n7IGkK4ipMUZhejE+S3T35er6dqJnhF/uitWhb1gG6O+Dr3yBWsI
K78aSLtSlu2mhiGjUhbFRvbEHq+oRqCHsqdku9r57crkfOfJlxkHefKtmExjTCv5
OQllpZKJ3ll8nmNkJFJEhDju4jjpnlAuzggb+PzJ/imG4xwmoiCpoKLd842RBFcd
4ZecoIv2by3sVQQJePyNvBuxBQDtUbm1pIXBCNtCJznR7Og4zslQ8HuUsBKoNJRI
i+jHvm/yan1EzbC9nMOrlHRhAKG8CBgAYV1cwQFVBsw1iEwze3XNp0vKOZ6SLTQe
utUKjLT9uXkUvaqxgcnO5jNqhdqB6hSXHSiGUnDRIoOfR5nzR4w9mdQYBb+2zmjt
pIqWTziTn9m6axf9nI9Pr2zldu7V7AS2D4iZH3ovnoR/3rXnlgvCn1KPO52HInyj
//99nAlUGlDqgbHQFzC7UDBBkZ/+PNzAte4YmHVd/Q8bRawr+AbPXUoQwjbqwITw
xvFE7mSj542BV1s7j7AhV4bVLmbS+uidBj8ZN9QGgCrYQSjdj04HgHF+ebdAKWcC
unWs8ZbzWVL/XKVR+3A1y/JPyW4y7lyVrffx7p8bn1Gloq/VlqclEt+BtMvJB9xA
wSnTKlA0zT36o9QbsQrMv/7xUbSHk6XHdo7Efw22Xweocz2RDfxh3FxpPZTuRJZZ
64OlnPukOy8HaEVbmu+h2bmIJiDMafTuPcWGLdZ8NyPrKiuUjIhKaX2kE4DA9CT5
JwtmGK7zo0CQkm3d9Md8ogTr9Pnc2O4uYTxgWO9pWhA/5FXJz2uiNbeZioNTuNc0
QD6oZ7nwQ4YzcRL0X4FjNdKTbg0IRN6FnHWIBZoD0xf/G+5F346IgzxKZNpi9Ivw
gWcWoe30K9EvAuEswQ98V7zi7A4aJMVh4rEw2QuD8CoP8F1TFjStHke7vFHXIG0v
3iAcn9JtwcGPOe+BGAwkgDnYA/F2a0Bt/rdDObdByL+Bw5xmT4IMy/cgjZbQw6ib
XPKyAJC6HRTcDBlNBqv0DD+OaXzqO7zqSyCE3yWW3persVuzzqz0e2dnGYC1R/yY
wMcUTdSrwFFLRqGCQBfdc9zdxFbJ6RCP21eVpFpe3yEhaUJ0G+Tu6WVoGyYV1Lds
NUSXRUohDoZN1T/XQ4Qh0bO4kViCXHZNOcwOiOm8qh9uuBfuujtAq8q3t2CmhFiy
56TVxqgJrGt+Z4vVZsTsukm6+a6X05OfxArvOmReFrlpVqQAaGGmgRnmXHWYdPzw
yKwzV/imFvdMCSxiElS9zog1MKfaeK9x9K1zu21APOGQl9bhxoz2ZCQ7lxcOPty3
olslA1Wh3UkHD4/4XTrQLI5JSMD1gFAlA7tcL+o7DUEhM+b9zoSt+etZVUjV3QrR
5bUoLO+8k2t2z2700SFNJiu/s8QjQ/qsNyH99qW/uxReud6lq50h+NGWLKHlPdPL
+l58YAy+QnyhnXM7frFKs4l2L/559yAG3V5OEOdCTb1P1O5+OsAJDJL9qE2NqWgZ
cJt26oZNiVnyIOzDHqYhl3oir9KaGdgJOR7bJA6HeqYRYb4U+SvGxg0yLogP88HJ
jBS+eSZALDzkbqDt+j7YZ1UnC6986wj8LsWK6/Lqfc66BrrkWPMqpYKJ4YQa9xEa
b79mDgi5VvU/Mg3vd0WRk5nXlfmrHTiQwNfgsANYC7PhEujDHBciuCUiipIWm5gA
bnTGW8/8ifbtxjfk3a2KFfpYezlokcXwwbsNEMzmtZfXH3Nog2G2mYGjKjZRabk5
8cbyZXzUulY8tedjCpjpn3mkbT//dCL073ZoOFyJtwMxX0NNH/DTA2jDsL7p/pq3
Ak0G/lU3bRryw4nO3k3CZTI4rLb05dlvIH6EVdW07cy9w2V8qsYx5pIE7eJRKAk2
V5Xsjl/sGp9wJs0UQv5ClIqX0arOiWYOcdrL6375PMCsswzIb8xtpm9I4e+IQgUG
DpYCOUcR6i28HNMC075aWPh8BFUINu5w8Z2850VdZYyDviQpXyhr2s8IWApFVk1o
IBbgRxTQEwVwZNn261TdOoGh2ToXBSzscquWJXAmz6+MeYJDI5R2pxVPXhykwXg2
y97if6c5F6MxpANJSilAvlU+umNRo6QRiFSn+hyV0/WkNowrQhpDBohuQdpeL4FP
QOLNu21WJnfSNCrCZIhaFkXZ8he+NuKkzJzGGf/MQCh6gThbY3edOFZXEhsYEubT
l9Osa23fL2wG9tD1KGTe6dHyViW37gdATLpWtznJV5Ox+iyABVtIZarzTsnCOCyw
XlqNHH5sv/q2hqPffwgK1kX2jMtb1EkGrJIynh7PmFOw0c+6ZZQhW8oo9Y8ofgFl
6bWFV3wvVxM67Aa5j4En86vvYNoVCiXt1+XLDCeT9wk+vZvgPrwQePv1SSIsEQ05
piOQDhtg2r6B2eqzfl0Yv9xqFk4R6nsRshXvH8ByYkpt2e1qCl5+arjYq/1BQ1CE
FtHgOEejAOLlSJe92eOuDyKiDqtxXt+4V952AzbUA/TnJm1gBb6W1+oCdT9v7soG
A84T6jheqwS047EtyOJg3PXWpMIRDhvQi163kM1qVnJDKh+7VUhQK3mUcJ7zgRce
HZaJ/xUvmNnJWIS6zjVTZ5qfs8O+L15fqROIj+D2kVkOmriBxRs8Wj9fFoqvsh2y
v6khNE5mcTKs5Map8zarnVP5zo5EKnBULkavrmtNxXOCZ0cMy27KmtomEg205eqH
zDEtMCjx/pgEcVoxd0mjeVPYRXD5Psxcj2ue3Yqxz9L0M4FHObZe89Iaqz/J2OoS
cWTUaCYda6M3biVk5Q9UmAkT+BV/CeGNp2FL9DlsvYcvBnyoB55EMPxY+Gi18bta
j1Lb2xW050tR3t7frtT1NF6ouwk63VUwtGliPhGkv4MU4ke/8yuSYg5C3hy6s1ro
3H6I0mGMiSUITEXtFInCmvymIpp+ISemrWyDTjqyCH7l2BzaJRi24s8wH1SAgDBT
QLCa3h2wsZ39Ll92AjhQcQ0YYYl58EQ3VuB2g+3aJgXHM+kKBukflv5S7qmTUizT
YrAx+lN6ggPOKk++mbiPxBkRd09958LkLKqqhZMfMeVjSMuH3bBLktlZcwIJTO5W
HC6U50PRhaQSv3JKsKwuvHe5utm8fevZJbWCv3MkAXPnELY58F1Cdgj3rKyvguPi
0u5/NvFUjSjdvolsI0eJjkTuKGiNNLgBoEeIgRKpOyouB91VUC4s538dgtUdRAld
ArsMSy/Ugf96+oVHCdhxVSyehZXZA7Di2/PRhwG7l7588sAUzc3F8ww17XlhJ/ym
DAhyljegUcajRfqAXizw+mjC0Rz6A0wuC3yXLzMWL22ORTUNlh4ReQMhxCYHUnp/
Rq5DxdHexysS3VCAdKP+q1Sv0jPn2AvR6jFChnRcnnhCk3vShZz5zUFCuhH5IgHl
SCUvbprguruPTcwLpDAQLYzkPXwDnBkMfRQDNcN8enlPabcdbjnKVntRKMPsKtti
Ei4u/AIXFRg3YPEzJaZoXo6dLQmKGXre8HfVTvwqy8N9m4dj89U6L/vy722OfjNC
S11EwRSpfxBkLiGZPQzhqbcQH90YpEe0NgQB80KFAoYBE0AOZnegP29DAS9lseRc
cA1WHSTvvN1i/4qHODy9IEJvr4ReePZQE0hVRSUhmtnMLwAlOzlQGiur5tXP0pE+
cqW5K63EecrwT1pZMOmpWRxQKIjSYYa3PS+q0PwfBYlux9N5eWuatINHYv6PsBQV
9n4eBdzKOXCTOx/ybWRqVKvXX2lTrxa4wshk76ZvPyNbVdo0K0p7Ktwv5eqL7LU6
NOZhU3Z6vDCok93lLvvp/ZqNXhl7+siERsHzBuDsWR8CbPUPrYYndkOqoRZrfIfW
cQJ9iSzAz4NWVbBD4venyleK94mrxEDSpYSZgjx3uihhZgBGo+hoZ0olP5CvpiKq
2T2GcwCnKc2Nn6hRJmRyn670FHU6hB3fBFmdAz2TgN7xUcTZZSgCUGlUFB2X6sRO
1i6WwXQ5HATtbgaZ+Dp7U+X5mwLSifMqWC0rn6ls7nq4cbyaAdcM74VL8FA+/XyR
AkXvFWhGcY9jdSltAQl1RUN1dPAqQdrr7ur6ZpquQOw+bAeUyT4JIqTEL/rvIHiK
Vl8fSnNXEsD/sQCNj1jetC47+pgh599TgFaWQ4EnlZw90Z+ozPsZ6/n4OSGQWivJ
szpOJeQdIjHjQLI3sy1Gs+GJPeM0OnBEBxsIcb5KRJkfN/Z1e10ajQSl3XF+0iow
vZB7UvSoKjX/OZyzYKmOhoPRtXq0K9YxsJJVthOvCGjOgGvx3A+Go6gMjGau5GqO
8TyT13ViRTPwPY4LhfvhXGxwg9unmTSXrM5DkKK7WRPkQ+Tr+niWqTPU/Sn1arIG
fCUCFFkmLNlOJGCq1mlCT3o7aIDVohauHkxDcfEQBWiKuKHl0PUoYQGV6CpMLrkX
ZzcZmjsV/mijmGVhV+nd7w==
`protect end_protected