`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 34752 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
0ivLeOT4zMq5S+D+IkEISHV0NKC3Ja/pvCF7pSckEwDHhfnVu9kkZHP4BAyjoNLh
cGMxDDG0G5xiKtvxTddwT6Z7EjH+IHUk8pF3iVWCOjnRSCuDBki5nE+c9mXIuMKJ
o1ZPF/9AiQ3swSiS9MyFGwToo+6QLlE4BmVwqpPaoMzjLGOTL3+hTeNTYA3fphEy
IJBi1NNtJDOFLSmAVDtvPABiIRQ5COHcrj+ZOOowKfV8KADmC/BZN07DscNeQOMt
0EsJ4NAoHTKiohWId3qNDe/PKCN1yhzSFiT2sa8wjS213NcBkPGroByUy/o1fJhP
IjYKgS6Z7gRix6g8cF2/gdrmiQfqrX7byu9QBSevPnF/U66xcw4N0gaySSxhVklz
tUdAxMyRGsqhLkQAdjeTr7o1Ow0e/jW4b2ZTKj7riWiayhWwQL/3RV6J5cI0DxK6
SymXpIXOQ432oJZDDDGgVb8x6nzX/YHLVv5kBhLIHcIDoH+EH5p9yC/RXjyXMOWa
gmnwf59U8fami9YMYc+Ag9i5C3SWCR5bYp/U0i/6hLw2+4Zr/ntipaWitOAJXMjl
j8r14wc7RGvkMXQXyNQtO4t6ed0gCv1LKKkhqRA0zHbn7Hi+wGNNGWb+dBkdWwby
pPAbzy4AIJkk9DeejC6vApBmVKBmd340NBN/w1AkX15F8mi4J8Jyd86sLUjmODL/
UmttKFJOY6wDjGlPrF8NRqdsPKInUzB5utQ1z37zDHxHazOivo6FifrkhGz/K4xr
KNH6Ld3At1RaAj55VlbeFul7DCRWZ/Ssb7b5BjwJDdb6brM+vILAnpOdEFnJ4W8b
Gcp9aBgUqOvymuqRmdPvgEXBLvmR2Y5izPlgYJhKKL5EgzV1vFVtp6MEztPGjSR3
GO1vxp7ke7PxCL2XwoIrA1qfIAHrSxDTBRS2PZfb21vJOVlA01+ExGCJ2sD7jn7A
HqfUzLGb7HD4JSl7VIO8R3HZf6jgigcniyFo75QP2lbFO8Z3FXPIZ11qcPXyYjoS
bcPB3rg/ibVo2lI94aGkQu9kIHladG1TvicPcEr9XFyPSRRyDrePdvliGRvk1UwM
604fv58QoI8UIqE38YSuG4Joi5+K5FXq8Vv5yHvjQlo19NM/RDRizLvBmbJhcsFs
VvOi4r8FxKXSWFdSDnj/F4BzNnCSod+evHYXgo9FEG5A74h9hXIvb4IPeVXwjnFa
vtqE5pUMxgkJCR0PMk+H7Sg4A+VDlEjaPS7XQAdQfYtgVzybbjPcDMHflUddcJ3Y
aTyZUjMGzUAP08WLVrWU1/PspRQSljWENSsy/a7e8Q015MsGIVF4QuI80UHtHzoB
1gulS2t7VeYM2t5tAZ5SM34c4eUeeRbLf55q/jABAdcu60cd6uDGMMsNe3zd7Fab
NduE0zaVQZ+1kknRbDhDVJYIUMVvKKqN6rQIdHU/lztXW+z6QsLZ28JlNhfj/jzN
KHpOpjsAnPf8C7xfFOeT/rcYcZxQd0ebed8pqj5k8/fAyCW2+Gej9WV75UopVslK
QqP811zwdfGWGLPw07+fJiXMm4+cnFUL0dubJP1OJ7GQQTaeZLgXCGWXTqyMGm0n
/nSqcKsmS/fIShdOdl/LztMb+78/y8pw9ezxyPBb9dbyMuAcrmoAannzZyJ+pYMa
5+wHS2BR+fFrLAlbZNlXUJnlXPAToo4zxQL989Sqg6dgWSz15/dD/yBPmDPo9Y0R
AtjHDypHw1POebF+qgldxXN+JkR3jBdds6YzND3xFI5KMmOrhK9X/9tkrXEPQnvs
uw3j+I4HVoEld4ttosp7vsq9sNe7K+Zo+Z+09+r6B467R+OZ8PY4Fs8SipSVK+VA
3Tv62cG6FOQXl0e6kDVy2rjbEnv9UD+2oV32UmMyyYt+BuM6b2caHuMHZt+sKuQl
fwZef5Nrk2///1AgOlVRgGwpMToTmYDPWOQ/VKjCmLDJCjPZf0DnZYwGoYvC6Z2a
ia0ctmEEIT2zYik7/l7LMxYOZ/VPGFfhYuqFx/Z0nerYruBCt3/xia6ZjYPecHJ3
l2S4F7vnN3y1Zx+31giczpcrG+vJy9piZOKAis+HrstN5CSiZOEYwVfejWpHM3eY
TMlaO6ht/dcBpsZmmvPFegXV8AJZkwPVI4D2c2zPjwBpjgakytTUhUB5WW3+fK2r
oQjvdmuNSNsvK3VPworQGOS48DL2ydQGsrxyaVwQcSL5YUeEBPPiKJmpng3NKgHe
ukBz2GuF+t6WNpaYjMSZBxzMkZRtG+QKYcTrPFTkS/YUEPUWu4GJumtV/d9r/CLZ
WNrNkiV78YGZBHj3vS/aHxOak3lKovHmIu2OwUsJ3YgMRc29l0sk4OkmGcYIOuzK
dLAUfP+nVJP2HkmP2afDz/nW9+uJ/i4dRFZ4Oi0l/6bSFZkXbi23bXj/ekmw0V7u
ENls3WZaz29RENd9NRWur7A2Xuh07ayjkqo0uPJzjkc4HJnnTqZDR2UV6AjsfuX8
mQIDRMBp46LLOZCeq8fPLxdUf7BzVNtCTvo0d9mH8+Wcv34FJAV0AGegiT4lUnsI
JkidqVIJd5Ly1UNC0TJpSG1UUPjgh+QIwpsbkWgiDw798tDKqeEJLLvyxNmOkwzU
46nqF/jxRz+6z4pix/en17Um+W0aWfUpGL+aUL6P3lIn/wOD97UkAQMEFHrPbkpJ
sUszhosgUluodXVwzVQtRPz+s15a0q41LD+TgoyteUmZhS0Z3oDwxVVIQ9dewLQA
YyFO3vRcm6RDVqpKJAP82lqufBeQ3tg6hywlkfTdjFP4p6mvuK7ajbpHDfSKafrh
LvxSeW/ggXI6aTxwdpXCtMZuK9ren//Im2hfe9j/KhIoE6Upo69g2mxiSi2rXrMU
7rA7UBQSuzS97UbIJNe+M4rOz/UP4EVsiJU/WuBg9pnU4Zze/IOm3eTHvE8iaITf
1ors+KhhTUgB+gli/H5g2BbzqHE74weWnFDr1dhKvAa0IE4b7yxY900QvhqPfMqY
FYjZDCVdHw8WDB3ZF0RITt6cM7gcfgMc7GhU47NuHLwYkeM4zKh1oA+klaZN7m+2
fFlosgoQOnhEmyPQQyk9HAug/gQrr0egO2/R4dDHdU25+B6nwU5OhJc3KSrxcM+P
yRsn4JHdRS2ACFzfab2CQ8xcv9uVcQSgmmgtHFCv6+xwf8GP6iul7LCYx7nCgpAh
NQZw77TequMKKlzHIlDMdvfX1YQEy2k8oUYzgCrsXkW8EzBmaz8aFhqu4zcyRsf4
SrBwvhJ5Ff/YUz2Ia4Y1I2DiukER8K2iLkew0RH7JQwJAtavHQp1aP3lQ7qIkEs5
AICEA86pwfgAKgOWdkZtXXzY5YORRKs0Cb6VG0I5BmivKyg4dV+KH9nCCy1Xvksc
Y1LZnkSZOgqy36/r1j7RsaR84nT9uy+Y4/ZqgltnP+xLbklM+Iq9iclMMGfG4Fup
YAGxvxNl/AcGo9vPDJKmKj6NdyZ22i0o1m/nsN4+NLjWY2h21HbnVwggK5+8ptpO
3KssbQn5xcRj9AL/6fE57Q85KHCxwRy/wvGEel/MY7FDAPcA4eIM6+DL2tzJOF5T
0VRvc6tk6pGqEjfMWYTPvQr9mqg4E3U3+mevq/PNTr0Eoq6i4p+ae3bHQVKhZvtA
I24nP/6Jttw8qUPvOt3KTcJdwmxRlGMuTOrzVDw3KccXJg+VgiQZyMySLGjara+R
jzZa5wbzVfNN9LKuZUkHZIquLebpuIU2Mq3XReoWMcQzxZyYwyCTm0sDDR3QzyuN
j3iIzoZ/5rBV84M+KqftG4QbOxC2qNXqvryD9E41By41a7omI5gH7nhFElo4IcY8
dPoLle++pEMTGIc/E8c8lCdsHAP8raDL4O8I88lh0tLYiY3Rqe3hoV8ShA6rquZ8
Bg6tHyQ3HZZ9pl25KbUaAP9E/akoZDDlZ/tBTLt3mgfxGZIcXioMOZAhLIUeYif7
xAxr9n5ll9h/OnwQNU4F5M3yfHvLMEmyxjgy7MZm3+xvwNosDCb/vVlTH7VHoNr8
ja9vAWeeQaTKf1iLr0LD5SZ3SE+0fm5oup53wfNNlhNrMyALzBFMxzA4But94l5s
CqonDsXhw56FWXfZjJ51Sg3gJNO81wDLmPzE/BR3HHpuddg+NrQKcewMFzGitcqo
3CYW2HPv5MfFIQXsMC58rD4HRgQKNmMWeysabqU3iO551ZVmf1WHvTCPRB0g7yx6
F8IfYTLQPXAVUMjD0dcIeQJ2Jt+sGp/OvzwXo05ga8Y7hoNrbwxEzJ8cMg8r+LX6
2dAlxF6KrdoegzppJ8haknMUfnoX6fPPzGr09S8xMywdAI/gSJ7ZHYoaQqKnDAbP
Ue6bR/gsOpqih45OW5XvMvy2Mc+OZuWxY79S/ULnUpoWn8pPsaNJxrCpHlJJZ86+
EM/NHqLAAilMO6SXVsC2MONHic29ORFni9YmiKdYtBQiIYRlQWQLDBUjy/KnxDrq
R3gcYs3lxbel5Cpj8oCu3Zt+hLfLYx3kQpMvw1xU3zwvntINfu9tsYeaHiSV9OIA
YyQvZjZ9lmQcnqg38pIWVSxENsrHCaKVGpsfc3NA0ChF9R3HLGsyHj8lq283yGvv
9S0jczM0ZGzO1zE+D1tfpCPHWliwwzA6I+Nlpjdnk7jGeEudsmVPPxxmVoyxGA+y
iYjWtSOV1Xc2OCtPd2FmSPW3CwKpD0QDW4nZvWmgbVHMg1kpMwDwvmQ8ou8Aao67
B4Mj7WUtShwWiOMgP3TdXhlNm71yEcGOAKOYazSUKSC94Sls3h1FYaNtkiS7M4T1
oOMlEZZoiHj034v4W/6LW1JnuqjA2LadO6/pIYHj9a5/p8s3We+XfBs/VO3YdDhf
/3kA+rPQtFy8JGW9onSoB/qtrRlQY/6OljbdJCpAWE3WVxOjTbjVKDGclRzlKmEb
jzl0FtVkshdch5C81SFY7i67dW+yKJhPpfETH5vb8U408/J07z9342KDTnzDyYOg
39doiE+SKnSEa1i0uGgOr7qTEk4No9XRXW0Azl+iY57ht7sj/KvvoMby2KiObtnH
WLbShnM3zifpwsSPg7do6cm5eP9LwmJjPoGPi216XAdtp5PS3FxSx05jvdm3znEF
CO8KGnUjwKxw481xgnuMhjSs4w2qe3rS8H9Fs7aWSR/reWzZu/PCG9DendhbxEGJ
SneyGHQfdFm6kYb3uzbwyDK4TVHPSNJCfq/wPYlVqIBEWadmpXozJfooed2dPzjB
t5nyEnWZFpvCGHY1H0wBtmNcNIvOFAZ0QkXyLCPnJuJKpR5vc1FNnSQ9sAMO/mLG
WEUgYNjvEI/nVvwPVMTKMaVZz4liKvac4Y7VqijRPV6ldnVVqHhOLmtxYq6ILA2k
/FO456JxSH/1P47T/fGd+BYrUCAIjd9FgmolG8dyogGfhvCFjya7L2KMYVntqkcM
C5e+AhmQKkoiWCs4k4gP4NfNYTnTlK6RVtilaJXHVHmyfpwYBEllvkXViNU6UMCt
r8Wbu2O6vbjAX+OSmxucf4GF/PXbcItIGhwYV8NnFMVmVjffXqc9LeCLhEa5hEh9
07Ea5nllJoQRM/Fk1jABWdRVwCPplbwrciS1/52gy6I7IA+dsvp1LcUYq8EQcz5y
zyzVrc/6dfJy0BZn3ZzFZkz93UhHQYxSXzwcNqnd9gNf0ZmVuabPlF5Wc2qR32Y6
naqJJxw0guUJ/HBmJsjy68RCRBs/yXFOIy4i4GlQHGuvwyz+l+geZewjrj2kXjMp
g2gW3D6Vyr17uei5TxYLvTD0Hk7qM3oI11WaTiAhKlgZXhAAcBfOu0hb8+SiLewK
RXqKLSSP3v0vyvVXTaKko1G7ZxhGwRakHafOLb2UwwCG+79dbYOvW41DvnY8066D
Uw/JaYN5O3431X5se/IZvxW9Yu8XyZJG5f3PzLd5MgMIwghitY+LxESSbIQw+iDl
D8I+qlA4Bwat1MoHVGLA+a9RCiYj99cTZMHE06WN3B6OwOQsapH3gz7ZqFmB0MWv
mrtvSG/N/wKLmbNkvr3AftlLs1rUKk1EEbdWbV5TIxXFvuv2k5RZNOtbXE2x5J0m
mxhgvjxwuT1qvFFAenVmJtzwuyKH/1W1mzY15qnu+EZBarxCBxgAFw/kBqFzB66d
8j0J2Lkcj+GUzv/XsNJ9kl7QZgM9FA6hnpu28MB5ztP5r3IFF60qz9bQ0rJz9l+a
lK9QNL6UFjQkur72WdFj7jP5h3uf+9O96qAn+bsszJm1+eJeFw7CVrgTj9VA+WdR
xtZmtW4hWFrIcOQuyl2T0yTaluiyF/TLD8uba/yRRYDPxMmMml8Pzp9b5YQx/thB
NFFcU8GnrwI8Nu0Ig/55go58RQnX5VjcMkXwRdHK1bbdh56d8KiAjAmxXHBtBggf
ph7AynUiBpet5GUL3tNScg6gkTzVH0Ea74ikkc+tskpN6c6fgyssDCvX6VEujRBA
Kwrwwmwg8o1gIQFABq5EDR8q3Iii00ovJMUwPVOnnzL6vrlqssHfMMFwRXEAQNhI
bW2MUicazPEndDf0g74SzuGETYSKv/hmrTXKMEZqWWkSvblCes8Tk3pCI1+P9Ov9
BWpgCLfiPE9Qtc5NDuWRzibtAhM71rHMZazio+xiKw3/a1QW0kCkXO5gn/KHhG2W
z+M3VeZrhy6NqVQb59JdMoKG44ZMn5d/1guhJSUFA/C8/njqHhqrIwIeoxHTgw9o
GDHOEAgfHgtHrnMJkVRH2jLpsPP8+VcDdMFdfJxTUBX3RM+KUkKrWvnwwU12E/Z6
OP57/3839gjr1kQUhf5Ju2jy3OCCV2q69/S89a+EC+EI0ES+KdXwBsY54QqmjvPm
PJsPfmsATlWZaWMKxR1PlDaCgPWF6wqGwpXzEucZH8V00URyFgywO0OWm96reFGw
3d236+T5LC0heF6mCxcmZosNgCJb0mr7gtNuaOZcoDEv99AZv6w2ijf3AcvROuwm
l02YPd1VmJ7bnUtxfTnqTCZXHS/PGRMVD+xn7Q+l9T1HjbjhcqI6riY9xzrWOLqf
SI6jU7PVGt/PGzExZXee4E8eoSE7x4qlpyh/97cgsntShDYYvJUf863AOv2sfmoD
e97EbPwHBAK3g2hVEd72RnuJyGCEuqz45I1kG5k6FhUidpozmHFIL0BZaLQgYIjr
m1VgNXbAeclXCH9qzLguehGjfK34rb8ZXeIso7wZc8Mk9/k7lOrSP1YmhQlP6/Xo
WqRY66N4D7RELTW9oqvBfUvHdem0UWDtDeLOqSOlLDGmx3Gt7au0y7ylc6HGXpYw
aK1PqbpoZ4MDP1LiTdsR9jxUbL8iqxOxjhyeJmFuDHQAIUqx8AidarlB9pKagg8c
rzpxMh2ztMQvLs5IFQJtrj3ozSubrEb3F8nUJ5ZxXO5dk7LSdGGTkymp5px/OeV3
3yJ3z593Z6R7de3/Y6BzL9BsFbKPHOwh845r6WJ3DgBAwanaaHMBK5tERXt0tSMw
tcRFhB3FB7HXaURnhEp/V7mTkk4JOTdudVbwpNbX4y5wv58fCuXJos0Fr92Zk4Y6
REMyg3AtW8fBZmHszMARv93cSuPPZ3tSr6/zTqcVY0sJP+MCOBO5j8m5G4iqKdjt
sfXPCAMShj72dWsSYYJmvKzD+UbZ6ZRnq7fkwxAJuJJOhyZQcZ4cgXzB8Rdru/QR
Lxtl5PgPEykyP3XAAX+SIPMKPcfJg9btP7xQNhc5c2H/XSZyu4ToO6JpPYPlSDio
sgLpPdgs9N+b+8ttzrO2WT/CeOkhoigei4TooxK0RdTXyr8XteweZ3sO3dxTmdvU
h3uMcPWdU8Am+Zxnz4OiCMNIvVjJzlphWG0KZF2T4vtVSLZ2BAO8U18mOMdb7jK2
seTAzLBKjoRhLP4YSBguKijnQsvfZUs/JK/nHNxmUmwnmuEbnNqd1vKNLO3Rxt/x
OMftUv4304IxdRNw0q2yO55owfLeMx+8zCp5lvpAO9Qccd6phMd1gVlyyQ/oaxTJ
Aq8zN/sPBuNUswEtorBH/wZKHV62JsOpvbru+jTlGiTAzJl71+qmSlNvV6x6X0zH
PD87+5P959nJgRrbis6zCUqT15UxKJZGUtIfFpSSuxqZmyPShwv2LWj3Em/NOIgr
Nl8aNkPRDGNgjZAVo5P3yRAeqF9dIx9H9GpFpA4nrHdC5XqNoYeYKPdB1/PzibZZ
nqFda4UZ/y8y2GMKnYX+9/dZwoGYw6FIrDsu9EYvmdxyxugpSYAvdJ3705VxPRwE
UhqAs+YAM1S/7a2mYaPyL05h2+7kUwFkS52ob+w5ZIoYUVZljN/vP+DAGOVS5iSj
jsk5L7/u15j/C+AgZ2/79aYegb4ff1bJQBBF+n/ZobYb5kdDIrwbYpX75O1kw6kQ
9sDifgsgpq+9hXtUMNuIjZ9iZ6VRV8jRGTKXfVGqtQe/Iwc43DT6QyStqwPH71hW
JhzYhKyFizfYVRWVO4SAZLboFlZ+LcZxb73DCRlO0HaaJnRxq9a0sVnHGMQRDyDF
WYLZsWb3Ukav79zqzZsVBMztSWd1KpUl5PnbYQ3ZaiK+vj0LJCs1A+cwOSs+jMSc
Ki/HVPyqulYfzoap/Ocb5NQZJm2XFlzrHHSgS6+4MeJo6QH9eE5rgZagVJaKcw49
hWtPv79VDAYQF/32ciCv+/SEOvWLBOeemqTMByIlHiVji3uEFVpbn4HRYNX33pHG
c/dA7UxlVGO1AJBKnfWXBAfaPbEhF05fQ8AXyJx4cGi/uDS2u9Jg9js/vrdt2WpF
r7pBoej4Qc5bV+3gwWNAxw75lpyuqOMi8AsyijdihARUsqDE4Sjf7OiuTIjcmtZw
2f4upoNJ8PAIG/NZkVu0ENdl+EMCSxUstVZe48Z9Neh3gqyC0afMQ7nsoIDw45eC
GR1xSyj53hXgPEnxS2siyx4/1i9oC0Px8qtS6rHIFdXmzDxShfFw3kSNjWQwTMZH
3eIVT/7wWveMSXDpS4FoHLp0Us72GQBHWH8BV6ccx0ccXGN4uCvXVzh1DaSldLkN
ki5MtaFtj94Vq41UXwEA64YtAq4hH8Njk/gix9rTSM59ywZ9DKkUKbW/Ll1Acjyp
eA8GYUcuCxdH3U0XPu4biEw3ALpF+iL02gSmu5WYkiNNfZqWlhOHDrfkALJlv46F
Z+djhZnDC3lQygEXW01Ia4mrk8phLshoUq5V9I43mRz6xvTkPTY3KgkqsaaFD9F7
TZjlfpJ63kVPzZFDLmHEGeMFdApovpIxutOy6atIG18VP592evq4CR6AbjT3Om5n
480qmQHuJiB9BUK4krn528Vc0/WZtOWEi9eBOZfhbCdva6FIHiSqkpWzArecF+j4
gaeYvd3Tk1yfVqM4JWCPvFZf1fpyq3M+BpZROYBDMDXtpjfx0e1zkM+CA/M5rJ8+
a52Ao4Q1vCCvKeKaPLpoJ6PCs/5fWGFr41+acor0qwAfC8NIDyn6GHBGoVS4Qxuk
WKnkvbh3FYPreFBfhMCWsFDjr59SbcA4BunRLGYaceA96myxh/hQVzYTQNBzwKve
GOTHGoQLiVD5BPQDA7rarcVw7Ks3xVHJ7VxlrSBv5CqmQ4pcuWfhe0Cs0r2NGSs9
XH3YFDP0Mf161AegpnQMoJTJ4y9F9zKgtFxW4rW4URojcb0VawyIgFbFg2rYdbVs
aFAfybIIP2oBDX7V+7VrEMaoj2ITW7eU2QA3BylHw5muAhIjhIPfGcsPzjo77fMr
fsxYL5TWUFKdOLi+tJMkiJmngucPgPSqo/xC+BUdX6/U0P+16N8TnQuKfKBLiYtp
/CHQDiHdSGrYwwiln4DYB419CzEFDrQ5ncKAi9w/23c73AQG1K3GzbaYZ4cNdsh3
IeheQKFy0dAi6URlUyF0OZFxEhnsOai/c4eQkFrjIbLfp2aLbx9SBIqBSLJB23t2
jy27NGcUwOCUgBv+XI7T5ratELa4W2pUeS6WQzhKgwIuLJ0qN730SfDLOVKSpyxh
LGDqVhJIq383MfFke11oGrgYoCB6mKhZCkpggCsPKdaCzDg84p2HDYxdly/B9v0q
NrglQuT0ccJkmLRdEUQMWuZU0qJDS19tgLivpbx2fiQz1lZ3d/onwmVmk02kt1x3
ArDDfRy84SwIiTa3TvtpBDkVjy7sF0JyV88e9vdMj8gmTJxup06tIamSq8CJO6J3
rk56nTkd5cNSbhQ4CO8A7PLX6rzPtPduqU22TPQtr7Qh7gg4ISmuZ3kBRU/gN8hf
m10diluq+T5dpkhQQwhprvykGt/Of4HdfxHuq81p+x8NLtwCiQkjeRnlJ4Tc0ZBW
o7vsx0DwF9hHHsJ/6kpbM1jY+pXTYzPuNnleuI7C2/NwzM3O1Uo9cOVQ6xTqX795
sRvIxCBP05RZYRzbBoltmgQf6ewUrYuEEVi59gpJDZSb++J6r9f6gvKdx99QJmiL
K9ebRJXnn3a7RdS08ZWpa0kz2C7uubDgICBergojanM2KftdDdqQE9cIN9X1eD2K
XJf18vdsutou85feXZKkR7QNvqnxhS7UaHrG9XKXTfSoduFZ1mAhJC+AIJ4ICI+X
23kHgYxOWfSoFZipfF5t4sA4bNLWG8C0XjJ97BMW+y0q3WohvJ0WPiW26R1r8uFr
pmz+n/Ehdh3wLvmukGQ5LqCUs4YNGBTjSJRKDhqpg0ls6ecwiRUOV1b2WQHxyjZy
CacFQmHeKTwplhyV6g1RL2VqxCGs9p47qQ4n0nSz4MfmVzxhDP9KjzbA7g8l8n/D
1j8JK7TgSCcR1CxYGnqR9C/ZKQDZzUshfAGrSxd6PSlahwb5P+HVIZBsrXJuMAha
BNISZG084VtXEdZMfUA5a/ZvqB94DEVxA+ZM7A0NuEXs+MebwgDr8oEiJuGT9fuX
VfywqsktIYRkr1fmcVZrO9gf1jcWJUGgp4hmb3GuD4ftBcxXVq+y8wIKYndnIpZW
GCnT8S7rK0+txzSPUm85kskiqdMd6b3Tw+qYL9CQ8zJ1gRBbkN2Yaf2APqUUnYfM
LQCQsYcfZsLV7RJDnELvjNGa+DgGwdemWNWqAu++69rCgScafdarZC8gDjY+P1d5
wCURV0qDXH3u/EcCcIy2yDcN6NCvRLjhMXzNnTyZ9SR1vmaqSZOwW7XR+vNDePkF
026WFOw3nEQAXiBkXjg2elMgvLNfJsulKC8O8ScHEHfy/a3zOK63fd4fawXWWvvg
hThINu34MU72C+C9tDnjvlLJE51Ik5IXSwwzBL3pATi16KzZMfu++bMAWcEQFbBA
j/GkNxHZVasK5fguNWi3ru+qJz0HoWf9t/dfoP1GGpbBoWhNawaHrxAkBGSsYnW8
/0Uyh/5ZckQOvvqHSHHq9v8LOtuxtrBF2DdJqe8adNfuHIY5nMK0H3rEKOXCT9Ph
W5t5i0N7B2vyiAo2nu5+SzdWTA+NeYegP3+LQUN0njBgpN6uacLvnopARoLMv67U
A9vdYLwwZ+9hSavYq3xXCU52WrGv7nEhvboc6UvkGku8eyna3uJCPQ8BNkU403d9
o4RZmaWhascZzmB2rqdixcXN4qHe0RS7QCrQtVJM3fgVMZjYqME+HjqTg2olsNDa
D5uQIQFPLQrho4PKweuZVQaJJcDoqdYIDr+VObKbzvrKZxKcdjDUXfJekWEWu1KW
D1bWbVjsoyf/UYOgDkiQgICdvaXpbH83Bj2mtCzfsE061eJE1Gf9PegpV5hFC+Ya
3oFqXypjYkU/WEZSes4SVtAO5y1RoDh3iOOZxjPKOn0lnp5EKOcOvfCmJHqRkMkH
uxfLLrsfIvQUYjDm+vmVTWhNSFLBlGacHtqdsZWElhZ6jFdaLoq/rdq0gfrqWdCZ
K0IIcRWB4ypDJQFHz4OZhse9XW8nRFngCzxATefea+LS4roCq7C1rqYTEcHspZl8
FfK54OCnKJ/uITl3z6LiG+TZ+Uqxfyz7kh72hGUELVlj+OSzUtn/UNTSFtKR7kA0
p6JiJ+L+TYklveF+AO74Kddel6pU4FvqWmPsw69p2XhAJ9pbIbgZehcJNuXwyMWt
FTEPmk+WKZ1B1qKmL4QhMY3su6l5fpHolUmExDdgTQ1tOF8+aMZ0lvyGn4hbUx/H
l8JiFQFo1pq0SyZhskavvAT4wDfBI+jwVKSN3Zj8sZ8zM/nAQk6Tc1dVwOBmQM5e
kGqdP+091tavuiwkfX8zrbCjtOoIY3uqSWjzD0xk3aCLzTZ3Mr0yYGaJZvinozBw
rWO8YYCVj7j7NwN3BqsFymhWi86waGthU6Nz/f+P9RCRDR/mnV6JTp26ReopnraZ
+3McSqX2EB+A1wFw3qYWpN1g0dPoD1assnnyPcFkmRrhNsswuofxOeOVXATMQX8v
2LeuguMxTwOCr6Yg2eiQcs19qy72si0VxTW4oBFZ9xCJp3nN9lEZxo3d8jehYOc0
17AmoAW+XDsJN46/jSDzpWe8TBcGfNaFrVq0oq8P+6n336AjILmSqnYEuqWc1Z8D
Xi/5jFT/fa62J4jLql9YyZ0jxqwj4+/xEi2PNalXkBwt6ixAIoiQIvWEcePRkUaT
D4AQ3B2EYw8gfA+s6gI5TtmkvXhMwtLFkA2MWI2L+BSp7UzDT4/aM1P0gZnKhsYp
83fMPdfNPFCeJsq1sactVx7IDXkO7WGvP/45JdUEqsqz4IvoYHD8JFZKGEl0/yjr
Yl3BgyAmm+eyLFKS0AM/7H58SE9p6MlJdkkUt/wHTK5ZFuzzkLqR8g7x1FFfVTxe
Nsp02RblDqUSzdTIf507i5t2B6NlF6TuQ04qsMx/1yv/2sRycyovgMqNFLM+ZITE
ClmPeubMaO+Csl8nJSjYCIw5+QcCBEf2VERG8rxAWPjI4QGY8lsErDxgOvu4eK6k
5BjKPrT/n/x7Sv7DbTRCNwXw6Z2z4MfAG+YntO+9imu1c2UBRKcUnriN3vLd76FI
XWJPQc8l8P1eWyaYamuO/qRZXqpheu5l2F9nauRcx70JAW/CFu0rpbyKTsdggNIw
x4mFB2MfQcdjiYqA8cLop+hVWKo8cthCKQNsP28tq9v+Xv3zT/8SoRtz21yRD2XB
x3aVaQPI1m93Ui+Vm/TN2NwhZO9NO97X2H2TH5zbwR+MErzw5sAKQydp4ZupiIPr
+MHwn1cGg9GT61jtDlnTSFf+tum7Bq1vcRz4RXUt3GOVqDncgI4oFqx3lSUDNatl
VvLCU0JzrBZKH4GBuDVKvWgt9ED5Oky/GwhqzLXvxGCc7uIms+X4M0HxKXbURfUc
rk91nz79FiXVAlE3u/SKsjmygMWu5D//OsaMaDo0Hkc3RF+/EQ8S2FgBiFUpHrEe
/T6wbzzBz+Jumr0BH2BvJk9XyD5dFf3tUs34op79g0cXbz78omdz1SN+8MdWuZ7f
+4h7M/+Gxztkhr39vqfp/EB4gOSlGnEQ8NWcNDi0CpEY8EC9tgWs91kuyfNTWmrK
a9kIlBx8nREDczNAIv46KD1fRSiV4D4/JkZ0dfotX2fsBr7UPT+watAeWq3nd5af
TgXHe8SHJs2zVjIBWNwQljei6KkjLjf27ovO0TsHFBIzWl8EuaTnaWF5pebZK2WN
mfQtMuUOaY7GXv1NsWT3/9H5hGyezrG2zJ3dVo3bqB4j8PM6+JbjJBhr8APbjIkz
UzEBpCX9+PyDoWLMkASVdDJwk+7Y3qQGqNjVxTffyYBgqN2dNPpSXWjaqgWYddOp
JRoy6qxJ/mn28m799U0/RKE7bjHQUKAvoYNDxfhPaV8EQShF9+iS9yabUhbXVaVP
pKO/fe93YBeDmmbvdUkhuvVWFExk9oPcCoiJvUuKvVgHeqcuEy16gj949aWqQ3bQ
tSAKo0M6L4BfZxJHEGyJIGVOncO2iAbXr16S9S7VF49myOLSbKYTdgkiaAYkkmYJ
VqIo7dNdGNFpn54p9RBsCVzKlwUCHPhi65FYdSttEpywvypByHY2vv7wqrtqi2tg
P4gd/cDJy8KD+SysY41dEHfHsw6IxNw1niLGkSj9a3+oKhLOFe3hHD6KQ9bTgm8u
dn2A5AyGVp2bax0iA7OTKSTs0DZZhtVlrnZMBZa9MZVcuKDJg9oCh+jmzopIg2ks
vn3f5uyuZ9hb5vueAgav9yFtCbtEa1J0ptoy0xqGACzOyJFNOjMYCp24dXYoPa7P
/vyTDnnSzGTY7yBxIag+e6KjLdQyNJBDWCaTnD6WDdcO42xpEJWZgxOZcT8G98r5
gRCTivUecSjhHpY/KYAHzJ8WtrJbeGOxamABaBTdPiC1NMG3hm9p9tcVQxlhApEx
mo4YgA6R7qTaBTohk7g7dS61LJMVnQhfZKkUQ4euKCjjUMGVGWflgtN+RRhzkdkM
lW1rd28RwD5ToXFgfQfO7lS8EN5z/7WiqZi0lxpM0Ag8YEcFT80gSwDZT4yF6ziY
o5RKIHV6tYwKdq5OZXgZOmOH1rzis4DYTLUGjglydl8wUW4VvA+VnbBp24Ak1dQM
354agpDnuklyR/fonW160rvEowg9dHVpQz45/svJusqWHz4GJfl81/WPRnjOudRI
hUbgEwYjDNVaCyJLIzJv6EuwvEvlcKkD87K+sc1wWwf6hK6nRdZozCfCNc0VERLM
Qpt1S1KIpTMYk7mvaWLqkKOTWnubecwdgOcrTGl6wwRxnet/FvBLd0KE2292wWhw
gsnrIq4UjsXLYNRmDN8/o8EBAFTnvMjI6Y8FRk/shiEnibVjuQuURehVM85IbmUZ
lWDZO6q14TKy/EKBbtjN6rZYDffO+Lnmicekm9Clsz2qGvi9U7udDonqRcnnHM8k
MF8Sc+48B3JUrGJCXpc46mBcwaslqjiAqkXI73O+aycBSHkoumFhgoR6oGw30SE2
WLBoEO25PP0em7szbKCUN3QQKfukWMPnVkEjAMBfFJj0jSCmz/FSf+MaMeITt/D4
2fckobJZ7bKuCwS0Ncqep+rroylL4M16es9TjAl5yfhr2BwSOBkqfbAhgoH1k9jC
tUs7FdWF6/jKytN8B3OCkThQiEAlOvSsCuBwFwEkDkGVKEcwSN8Id2Wut2we3+mw
yzWqdaynKILmgJVclubqJ3LRxLS1ZZnYstjuY+SyKVjbnblcmtMHRfTHf4VIaHfQ
38ZfrrAc91U8jXA+dn+6/Ssl2WY2mev9LQ9mjNCdsEiVqrGbBB4khX1mOdPouSTT
zxl/JSi+kTFBjDRv0/KO/C52oH+Nzb+wtBLbA5UVvmsG80jYUrQNTAfKw05krtNz
sitIx8jhcT45/74xcl6UjrIAo18IegtpMygQVLglP+3YywKGpcYeqfho+WLR1Spq
4xQB/a62thKxl4VYNZ/znNGMxj1yaaWwIxLPtPQWbqAXjaQwGQazo4xI6dz266sV
Eavpqx34U++lP3FNH9k1sRIYtRfozqdSgnvgAU9+kSlotPsQjsH5gadkAhdl+KkD
1LkHbnC7wYiAVuZGsg2Z/d8fbNcUXdijIfbf/lWtsUme4B041cwrUhpsnqPRM77W
B1h/bq+tvCSWfrq1UuvYFwkRZfmSOeGPw9MGCSneH0rZ5CzSX4pv+OUgM4pJr8yk
hCygvr6k/npU7LPn5KVvccZS9/CMmUGlHmMayiLD16ITeZsVvujTehwrOHoehKBi
Z4awrX7BO4YRH+konF4s0yCu6P1nEPUP9Cw93kBWp9p2M7wRti+5PPAeJCKryH1f
yfK/D4LxujY+4Z/2AcyXM0iUIkglS5GE+lKePZdWFsn4+1/A6gBbfcQwWCoU9bu/
5aa7xJgmjH4iua0Fp7Lj+DRJX19i4xGITcIwz9rPPN6ESpOoLC9qTt1aZVlEssS4
I4KSMPF0IcOIigDgPu0J01jY0BQ25BLJ3a1kv4+ptqOR50LV3ZZPIWhn7/Z61XB+
VSsa3/LPaBfrhGeNYIpmq8cW4yn/LqkOCi06+e0IIwBD0a/ILA7pHlLe25byoZcw
rzv6RpxyurAEW5uAaMEeNEM9Sul+rv0xyIPpJFVfeNvI9s81Aixd1dVHBqGxP49M
RPzIxE6kuqWavkiJT9AFzsm7/xdSLXZQcrZ43n1ZGBJ7lA5MJjQVbkgNxFRCHVs3
2N8B7hA9FdhVuehH62hRtt1PIndU3+ImEV313uT9T342i+8QYKLE4QlhKmlyYtqp
KaZLK70awJyZFt1VpCRsRqljTEIuM+QVrynKUJdDziQqJVMJDjFuXfqJfXcEuEqH
5Sy3kqUk+/itQHYYXc3phZ6K1qoOWWtRJ5xZlno1rV0Z5ewTSimllAlCrNx9o3BG
nIpeHxWWjiXn0c7bwYTCvk7T8qz2ElmCwUC0BA98Cxlt858Ffma+YIFOuJfay32V
rJ7cGwet0bvedsvW10FsJvqgFE2w9Ch26llrLzqwsds2Jkxtd2UXjSPIvzNxpcQ+
1H8NgcqZk3XkKWQ1dwY9WHwtdYrY6wavrq3mVXQVSSKGCs8VuTG8euj261NAirHx
YNp2cqvnKkR2kuraAkHqA6TBWljWVVwRitfYNJfzv8j3KM1aCK8ksid1aB43jHpk
rzewWB6s4CYwOYQovYuljSGYdVuh6U8oX3bD00YShrXPHPcSgBpsZw5nk6snNrNo
AnPV8uTg8dvhPyO9eCVgfNHWJPloczi3IcYw3dSQN6KNI6A3ajUTlJfrctf2my6w
lcSHW5u7zT4cu/qyIVmFg1Evgqljj83ZzUtANwj4Z4r1+4wnvet3Q+iUkj1PakfL
u9pYatZQflbjbprOMr67wqH886qzomhg32Hu4miaALyZr8/FDYMesds9EpqM0An1
qTm2XkYvL1PDvr1HOcVjdXm5QLYAeP0gtPYe0IpglTNhatQLrCv9M7cUZbmLGv8z
BhRZjMJluPG2JNsUqaoJeZTxZYSDTQQfJZ80tAAdK5JjepHfQzOTsbXY3WIf2oAT
R70oGO5GM059pn45z3dwZGEmXWsglg7vTlllwAqgzyIeQllwg/K8kZ2mX2jDJCcf
X2hejhMDgEcJkUqmaI4gboUiDJt4cGhSoCtu6oL6fjMNIWydrEbOSmiXCIi8qD3D
FngX7ebUh1No7iPSc+vrUQbBFrsYAa+qOTxPmFB0VZsQQUa7JAFBiuRBIJjR0DLA
9W8WiM7FkCXy3CQxSCtoNG3zUkUxi7AqFIe/PYOWeBM0Ivqt1vGhewhOvvBWpuOv
OryOcE6elmlRDg2u/WvSt7WjNFv9qnHAWu5BITxlhY6DFGCP5wSl+GIqm2YjjRJV
XiBxHRvAnaXZhPZstlZkP7imkXFGbhpkbLXPi4NB89bdERAF/NtX/pHpItvZunk+
8Lqhty73qvJdVpu6nmjbhidzOL2ER5aYziV1rfc6IhkATO00uU2Lp24QuJ5KP0IP
Bn4H1zTFrF5z/+ZgwH6hPlT1MqQ4tWzZcF9X9k1B3eEQ94bt6GBQfGrS1x/qJPrF
kqnoxxLRnaXOyVZY6y+r++Hk77PLttgOYYBxnL7enFZdgNEAswnj/8Tu0+jEWk/r
aUd2je6gjMzgtGJherZvojxdhs1pGLZGCCnm7KC6OnNPxQkvzxdCZJ7ghmhW57xm
q46gGmZgwPRhqkcfPdGE3ip7SnkFXOQBSosdmmeb2nOI98RHxR6PpELVYvi5MEmL
+VwoD4J4E0JXip41Tr2i7ETqPIrrldZgpDzQ+dBtf7Pz0C5w7LZVL22xStegYxaM
nBRF3+eDVrOR4HFv+nfcMWts4ukIs8h7WkCkDDQ9EkRG7EBAHAUItyt7kUJEqPEj
YjhYiez68f0af/6TbziOv7vlvad3nvvOGAM4/FElEGRrfZvm64LaJyFL8pMOusk7
6ECBPLP9+Z53X3LPQN/OH93ZZ7jGPlonu9fzEQ8j+cvTp9uoFWFO8cR9pAUm8tPm
J9PDV4mBnPrFxGJXUWgivDbBylfbzOjVQ+b7hNA0a4a0MQmeT4YCx5qvKwzyZEjv
2ur+0UNWj14jfYmM07yU70ebTkEPFP5ClRPb58NeawLjJ+Kz3vYd84H0NsK0Su9f
qPP1C6jrvZ7vT52ZNj5N/GPHAxwAr8ORhX5IXqf5v71H5+zk3iwSovkUxJ4dRn0q
xUp7ywfpuwpPUm2W2Juea0ngFOmwzLMn/KUWU2EgIcYg4BB8RuHdR4nPDk9epSOD
ghrmzRa+eqNcS0jT/ra6RKsnOVaK1QnEYi4r/eMorOIxABkHexod6vJ5n7F+BhTq
KT9zwXSsiSDEjv4IFmhs/YJF82J6tI4GybNBSUbPVmWErYwcUSUTe8EW8Q8/SzBw
+z4yK1EWsN1LfMOm5SuZqxFfk65mjRUiZKIOZVz8pTtETZpiSn1W9jJly+gSYbXd
0ObutsfMdcNpWfhcFaynkyXiBT5BBTywQmbOraW2UI/vTMsj027pmE7QB58U+fqQ
SUOFQrrVpi6bw04cS6a6qzrAEnnrFMod0UPWyHmmwE9jPox+4quv5uESQn68v+Ic
2JK2wbnZNPGwiAMmqXRx0KpvWQdz/QBlsRrwY8G2d1F1jqeU2kkUxAcyoHKVfAnz
QHyuYmvqLRx+4Ezr/MFvsWheCEf+B0r/Frb6MG0I99c9Ed43G/CpgXZNIiguVp9G
sOPSi3iRc7VOXRzwehMz5BGfqPT6nQSmD7t3aRi/v6N5a4bU1/rVmKUS/ap7jAg6
Y2nrlg5UC2Kx2+qcCl9SepUef9D3Ep9HCaiQ0plnI+BZYaMYZ80vPAfPxpkW7VE+
FqftJle1EAebp0lWkkYy8vc5P2RGJCZWvQQtgh8HSGUkzRqqzNfzpDqlp7OGwBnQ
TikgxfbifZfM/KSBOBmq9GcwFxwSRlbeZ/gyLa+e2QVv4ImPE2x1fKDJw5O6pQOf
YzkwIRcm6LqQKUqh/gL0gIxThQnqM0RBxqaycW1l+x3tzgivcsEuTucOpldtMgnM
D8DjcMMJyuyENabDCTDxWBVQ9aR4TRWtwyCc4ZFMotnHntYLbNwNotAMRH9J8u2h
gF0eFp11Pl1aWGvUibI3ruZBgKKdSPStgGBnqrNCAV/dwn1WOsZIPH9VyDrc9dg3
UggKwQZ0t2YuTcH9wuGiUfVhplEYiXiQRyQKDrsBnGRAoeRj35R4ODfWjnIzbfsU
sZ5/dP4TEdH8RZE3XUK5ScZW22xs5ZuNTSeyTbkheV/ZapNODuy4DWbdGsRTRnJR
XyFagJ3qDmQ/J1zVHs8tXdNVtbjSeAF5KXp1x1LrDMZy5msSURXtQVEFx3R3qOc6
QvEyrJShNHVwrr8UpF7vau3oJvL0LrYtPw9RtJtJZ/sAxNhjYeIQ4pK0SzN/p3lp
80QgBgeEuVo4AbOzOGBcj9pyKAPtNXAEdTTKQFDRM8LXsTByuh/CPvIr5BeJMv1D
QDjUngDopEHtdM/UlmfqfubcytxEgR9dHec4k3GYinGgVLifIOcRxlxEqkXpvJnV
ibwGeALB/pIXH4TH+6dI5laHYU5I8/1TKk7dNBZUIX0+Gyej1Lr+SLperVsSmqwf
nctysgYDmraP6TraAriSs5/JJyH9K47o6dWJ/NtAtfdCEz32brKHTsHeI+rP2lvA
glzv60LWs726xuWHps6mV4Uf3LUv2naTq8lBDXWQRwAbRNr235n+c+5L5bwzUpVY
joZ+/+dRP/jhAriwV4eaGceTg1jWgqkmBBz4+bMQvm6Lp0UTh7LyZlSpO2YhBdAI
JTda9xTFU6wcngAy1cKeJKSoCML2WLvrByp/0CQik9lwEna6j0zZWrHQEDGMynff
Ky1gPM1RW15HvcC7pOjhFT0nGTVxU+tURr+wqW4DNVf4OMP7gkvb06X++19bb+sW
oKzZZnLp9HujeQKwiqJ7hTW8GsWexDDT0ficfbzgb5Eha7mnsROVaS5nh3fIXcVO
MSNFO0wdX5ZF4mljlaawTrm4CHvAp3+KIQ1XGu/7sHN4mThmDGFUEJaG3jnJguxG
nQGI9PkI/IqLlzV3xGwPlVkfbm2+iBKMk/AOomuRfFQWuiqpJxPxDMrWvK8iXkxz
nluK53sP8SR8H23Lrg7zG7fWYVS9Dy42W+NEBP0NCwqEtuaM06Rc8kBWs7bDKuk3
KFKVi5ErlbyedszAqXOvyoPtuY3PN/bufWPQpHduBBJuME5XRbiHn1YMNEgVfwNG
amDXfmGr58JfX8ANk2DANjpp7sIwL45DyBeJlOuxuIVMmKSQlLfB26wepK97SVOG
bq9V8WI7bw0qy59Ntu9XB0MkPNzGBh//O8Dnv909gZoqRce4j/hGVue2LteA/Way
AustcNdrkukMnNOCB8TfOMpiLslSFoPSMIOYHJRf+CDQrKwo2jHtqCLtPmNNWVB6
+O+1FtsfAYXK4fbJ5KmjKSGs3lDx4Mf1MWoZeuv/oJoxMP/aslOxCd4L7opGUeSc
dDvtormwwsov3jf4iQP1hDW9bmVw/PNh5H69S8camkQOtfa/Cww42iDWxK1DZhDj
K1+pC1FhXydYTCheWW3jM7AsWlJEZwj6XIaXSUjGApjDXuIcLtla5ODlmGCc+A3N
XtF7L4FbnZFknxDvRP4zk/1j5zWvEduBB4R/dvA8+U8LgZcPbs24HA4XORIjQRFE
UcAO5bbi9175KdUbW9fYAQbsx88xiUEZsqKw7aYSnx+GmEdxnsb0yDwe7poH9CVJ
3PS+3JL0VrJ67XUKZKBZwSKAVBERJh4HVH+gWsmmKja6OjFInCiGeDXBCLkh2knc
46mBzZ3nYRHsO7T2wK/CesGePsRrUXAk0pC/k3D8aE8NHpNeYdCY1Mp9/i7YIfbF
Ns/B1ZhHmVhYpr+UhA33rdHAZVCFexUngeh/H5llu0eHpcTCgbsNNqZPX0JCa+RH
a/q+eAvN0lm4qJBg6BX70Havg+JTtT/zqKRQUoLzXaZqEmBmDD/c3YJxUEBJfqlY
30Hn1sr+QC5GA0RebGltczDVtcKWbRXzhCNSxU8TMVyogDpa4IGeP13DZu1GFUPg
iDVjPt6j3ppH11DU7aq9Qm/Hly7w1RGBSIYMvoRS8X1c9owzJ/Vfba92afo6mGxK
15+ONdvOHoGFWdbhXcA0xaSwgq1GyeMKS4BoYG5S9uYjuTr7w6d/vCkMvCKFRteC
VxgFI2NmR+/HMa6WbOTK5M4VBwKh8mN8rrbcozJdxVF6gLQZ99WkDGmKwwJsjh4o
49O99xCiDJANlhXVvC5OHu6yYKs2723q606ASiPkifjXiB8BdUIarX3G2uDBN/Xx
keGGNXI/8ZoqRC593xqpB4mawllL1MERlU+6B0p2w0VvDYvHgUtl3kTUceiWFLDQ
DYFHGzJJ2Cy83l43mqvEabLaoCCGnjUhVQVBQLYOGbUGn3/+qC8s7jf3Bth06JMZ
bxojWdcJMvgMiBV55Ueh0imAVv+svOdfBkY9rgiVxR0l+z3WC4HBuGYNZzKgLd2t
onopS211SrpbkDSTy7JbgjQEYBEBlVP7jIGJknpWZ5xt25tXjmZFFkhlbdYi3xcg
JAgDj/JckX89eroPNjrhR7F09jjQnz43zwwk73AoJ61cXGIvuLx+JfN1LgxtR2Nr
sciybVH3egXQHRRZNUcDN1APmFTO95WRbbyuOLjmaP/Y/lUyPdvFC1qHhq+wISyd
rZ2pSLUTijNzxOPiY/emRlLSInXvjjaR7qopSeZy+EFK4ByO/BhmenAoROo8GveS
gizuIgWRO5bKrEP6QZYb7xHcNq0/ZsLq8EDvDodPMzZ/JYqVjDARObzT2rXLePaF
zaYuo9hh3pGcSOwVdCCSgeXLWWkcFoIxX9WgyI15JYyWQ+jE4ZubUO8DtWpcNr1q
z3LsoN1zTfloqT6K2O2FzbzeFvAWo+cFujZej2dTKXJVFO+ZpnWeSG3r9Y2YJZ+T
DTSRwBEAoQUz3cvkdv8RbYGfhEEuw+Qc7dR1ItsAj6CnvipmVlb8anIq73FlgIXZ
QsNLrn2QPs4gev94Suk1W0ww7RfOz1wt41XB2b2ryusK8hE7FYBIxQ6wKpj4jcDh
81xpoSKcvYRMiCC9h6nhmr3Hlflntk2+PYnGBhh2fTc22oT3WFpqfK9ys4RcXIjx
c+Qh9dGUIFkFT5J9j3vpRD8Ikeock7NHG2WQdWbRlebtXndD/AJC9Y6aosAuZQKN
2+/q5inZg6QfEOWXewsvz27q8jP6NtvOvrymFDGSI7HDSb3RL/oOmrtjROGvJ+bo
pMKgoDUmt9YGmwcnxjj1ALMt0kGmWisADleY7VPsi87P/Uew3Od1V2gokT6BAizt
ScD+UaEb0z7gW9cxs8aE9mNkYHCv7HSeSfSLCQo4LaaGhWO6oKwaOi44ADBHUbHA
Vb73Y+mxM0kVft924/gEI8bnvU+l4ETj12iwbZob1seKCIgA/rxLRfZ/hnJQJWV1
iUwfY+tG1YrSyDG9FLplmz2kW/IdPHs0cgaXoIL+X2/kHP+Vk7s8sUYbrmbg4oe6
twPLo9u+WFj7aycXKs37GI5ViBg5EgYtJFoAG1K68tA536uaGRYobI606O0Dry3V
MeJriR1k9na3htHpSJoiA0pXoSSQkOPRQFGmgKsBwFea2hXx1udtJEMfKB+P+4/5
sRfyNOYzqt/dtJ/EOzNxpyl9q8dMtTBV7vbYhjzgvtz7eexgGZ1SMb9O2iUY+D0I
iAQWiXfKM1emqxoeS3dPR0pHcRFtQ6RoBcv6Kx51bxpSuv/72VXbqwEmrME23uNn
8/YmFD1nyyIVmo2mfWk68GWGd4Sy5vTEnxdMoQzgAhqSlb0CeZ21MIHLxRdqctNZ
D1bgd2U0qwR5osBTzDb7iP+H7irKWnyu3+sWutwihK2xzZs9Nr+2ugY+yQCiiSAd
0pYu7NFbTVWJjD1BJ+0WK0EcQu+oo5xXbN0g53m/p2K5zqFX7XRnOH+Rxo9zmS0W
+gf3Wzw8IiBnv99oD2GVn6U+54j3bZacCZ4jCoerOG/kq8Sa4We7Vb/9vZl3LuDZ
zDXNTBVw4Rk7ORvjtxOfIrEatU41UJOI6LVgIFfkYo1khXuCt74mE+vBxp/emN0b
sxkevQA4aGRcJ+t+SIPY8Yygqp5tPlob9HtK5s6N59cihr8KfNj0G6gyD9bHo3PS
0czrnanTRgWf3iFOflqcNZez7pnZ+ia6Y4vCxtJYj1QKv/W9rwDKzwSGaF+cs1G/
ibkdL2oSPu3DbfhnelBtOXZUYUhgdovZcc/N7hwnxflUPNOoM/SvPxg5tlgwmB0y
88l3gzAkFcAJ6+PRuM5Ku2rBEtjDxF74WV+YwaMfED9PXp95iPXSSIxbqYfgUX5C
CuG0Ufjbky2TmMB5VOfqMvSp+FLriCBiaKWsBBQ5zzAF+4EFiX7jpcNUtE8EqC8o
+vdN/pR1KfeBD/yMQSxRPeC28UUxCr/GvrDE05IUSpiUFCrRf50ma/7GuQdXORYo
+UTB2EPujOwIcJ+nRSncdsxy/LUFy77LUbRHoZFa5TQ2EGbM4G8JZ0iWhw1GsGKp
euuM40CIbyLovX1LBreh+LL/uS/6gKZszFnUoisa/+z4nYDDEg3ilc+9KjMTSR9H
a63Xw5LGE5+jIfXIi8/k/UpMUAmkUG9pLhX4Sr0I8yb/OW/J+7F/7WrUl3UszlyO
Qv2XsRXaWlTC5ES1Jlb+/RhdjY/QGBEYCGnfaHo1Fqy5jcYOXVRWs/bhPf4zZTy+
v4NLA35VooRMsS32upKYhb829QIALATKlt8/Nv9epmdQqLxcHP6Gc5iVM1rtw7Tt
O5u+yqedq/Q1WKNU5JYgLNfGd3UQ57RT0NJplbRitegL9dGJ6AziaNAM13XSFnw4
V1m8LCZ7uEmWSJl7Susmx+b3MGbMYgkIZ+QG+O1EY1h3sFmSvjwvfnIHZfHgKwuD
K4y88KiLNI+OFgvrFFQ2HsCtcTw7aHD/bLW7CXm/GNhCMsi7xlGuflEijzz9nkWx
EN6KnV/mlRKB/cVKtwSds4ccYF17C+XWwj35bi5gzLaWFqXJgCy5+H0ZkytDkPmw
NjZS6ezgEbXslKdzeR+5e9HHAtr1lOtpM+RYKpss8uaMpQ72p0ETvd0Qrmdyvfn9
kxx1ZTjTO6d+QGjVrgbLtKkDL9utJwUP4/ixbOobb3iUok4yH757ewAkL/P3APn9
qktBGNhJrMhDOMghErD7nfkEkE0yXrSN1jh6BOd9NuiTHg+Wy1qvvmBK1DLvUdkL
aK+geNtpuDN3wwkz/huZz6m1utB+Fuel9TJrDwnMWO+enoa4jOJaFB0ONhPNdWtL
rn7TGEcB/Mu+z6S1EFqQ6dms+sq1wlH+p8W8o3rXKGRy5GE9K1xTzeQ3a2vrZVlS
rh1+0BjE+mK8DoRy0VjJp8yKDk3xBMOaubUTfMXKpzcEV0L5uGj+imLUb/337wXo
mPN/iOjLmuCsLJNdECA79UARpcNK4MDKP18O0LFV8w9EyPpS3TrU12Sf+RhCfM8l
oD5DZ/ONOnol/qctPogDqf5TU5YONxZrXVUygNKqXEFqmu5T1Tb5G6KvEnio2/z/
6JRoR+f4MF1RgQPIy4FpVG/tbOprUXt8rxg5yPBZzpmXadpXMmzIyZpWp/M6nC1y
FE169gA8U7or6dSw9ilJ5PcrRk8r3C577X8qZenYmn/1TyeHcguDSEd0ahWsmJro
ctWWD/rH0i0prxOj3lkttNEGYEbYkz8VH056YLsbt51vxXutbka6h8Tf0UMYD2jo
SY1f8X9OpB5F8ABF4DogjebfwqdO2pdbByIN57+OKNhem6iXqvLq4IFuQK+eR+xo
dFQR3aYWHTe+XcUuHLuTlZWdR/35K3jURh3tMQAoVy6vU0ldIjKzhqZwI7ZzNJfM
CJF6MmZsrl2HlNtcvpIzQPe5XMRgBBqobsGmZ23+qoCErhS6gBiIu0QGz6vxfD0q
H3xLKn1YKRlE1BBrARtwpVGz7Lfd/16ZBSXfZqyx+GwVv+75tEPE2NzvrjbYT+G4
hPJ8toQvM+a/N2n0mOwJmATTz4xa7cIWaxSiH9FXiyEcdMUlIs+doJvVCNpyfQxG
r0EEOSo/iu+3mtTjGhHj3NwqaUa9oeObRmGHYdx2h5DYsXYzPM+iky2KnpX2WOfw
lC8fEwv4it4B2EMxPwsR1a/yy7GdhImcZ7QzvInGvG/sC6UDNuvqdLtuhZSVPgy+
0M9rU/g3t/kxKnm4QhCzYRiaPByDx3w9ycq8+M7bInEOJOwG9Du4BtU/a/hbbpIY
L/crQ8vEoJCQxwINGYPs5XYbE13q1oyob+CycS/ikoSi0WZwkZ1XLKQ5LuEoZpOb
Rsx6kYQ7ZlubtOkNPoIX9rn+bOtIYxoykByGg4dSLL779AUPdDK/8vJiCROjCzLI
BkuGYg6jOsfvttAdh+aZFv5ub/klfqjCSnw50HwyfIHEZnISkULXT4t7c86t75zG
jlgodJDLNcE/rO5KgnmQl0/c0mo3RpUOXKWoROo6Hggtw06kLDJXEozPPYcbt9OB
LT4ijYe2DDhxoe847fca9k9K0qAvbaKYi6WAmbmaZqF8M/dcUj0T26WRuJf/uT7L
+AC+3/4Hn7yZH9wwoz4ap59tN/qQUUUxTGV7l7jaAMtYUw7LyYxZoSHlfFCNTZso
a8xBy6EWon175lDILuJmYzmIYJ2n4gKbg8PxccpZvWxoPIabKG5Av1XXaRxWi2GL
+bKnC4CPkdgPeUpwoLa7vlNxRtibiQ4hnL7LWg/x425EH7QYRou4jn/MAokQaY0b
uN1d8U+NTCdR4ECiitYs9WaFGlhA1NaxZjf8jhkiYom1eHekqioRCjSSjzRYd3gP
tHJR3CWxuCS/wGsF/RhRYaYlA2rBXZfipiSDaULjDoSN4cFUmOROFli87LUujeNc
LLhalYTpGq96ZygXmIHiubfOeWF+xq8Bbes0zBnCOKEJ0ctgcKxIqmlWmzjZV9A6
jdkGL6lJMWwpULy0plwltxnXj3HcwBXZ7shvNbUf21A2u309qxuh/3ixM3b1ywg9
woeavDw+1CP8EI/Ob7GK1eyt70vrJQSZzi2CrstWEEsEH96YbXyQ0fftDzsKwLzH
/lWhRiEcAALFAZEOFwtACnCWJLEkDD0Mp8O9/T6PkRAuDNWbJkGQSoG8l1kWzd/p
kO27dFLFpsLmBPbqydNgPZKShZD1YSORym5t2EMzU1/+S8riefhrrvDldkfxMVsR
PQwSo8xcDZUO0J2CmYgq8aH3bosvxyZ5jhEyQCroTW3ep6zfL+aKDbOlo1i5loQw
gJCdfIgBX3KS1llieclTXwwaES1DFyZlJcIAPI56+eqICKaaWHWuhoSx+sHJqX9V
VHbn72tUEG7/BDMaGGhD1Taaq1uD25oRICWp8CHMm3YtvwpPqfna3nxFPwIQhGka
baxA4PRaLL8RfTVJKARNldLoVtC5if7mWe7sCsH+E1XEaxGBR54AY0LypIntCNNd
QZvoNYEwmYCvsphYdOFGzXy9+9lrOPT1fdWdMgHiBj0Uxp/XABFqYLI2uG4Bl7aT
o0irc8JodfGrI0OFXsmIlAmLZDegYNKMnqoJWl777jbzQay/27xE8RO9PQlvdBVx
WeDBbALOpWR3p00zNi52ERDYuNnJf7pwLDBMA9NWLegilCQ4YiLS2nB0n3n+nlRT
n1ARg5Q6Xoqk6oNQqqlocKsD22NhcQtGX3SvH8QS+LTG37fJFBQNf/reUGg5qL2k
jy4MCcrkutcRKxAVkK7+1z+M4bQ05dw/AAqBaSrmsrCrNSyrNphk2CSnK9M2PKUl
PYNajY8Qbc8lPo/xdez0LVLhRCfkK54JoW/jhWHd/W1twIy8UJR7Iu/8907kMv1X
m4RA8zLx1ZEEFPgh73W5udJeWg/vhZvd5lTgJYv15ixX6M4FRRtYJ4gT0AennG1u
RFZ3zHrAYx0IrtfRHsoXXf+XsAu7iKkqHiEbkJagImLx48L0ymXgNswwuvacjggv
KbmtKbnHfOLq38BzIhO6PpU8drws0yYYvnmPi3COYS/UMwqI2dlegq8xtMBTW9U0
A1rC4Kz8ya13gv9InsV4zhA7Udin3dX60q2bz6Zjiq2oGSCWOCNkK+ikwVlFpjt/
SqAuAg72LmWOgtIdBE1Tdwf93XwATU018TDvIe/7S0lGqDR50Rkoej54vislnSzV
Dsfgqid+p9lkjsy9TSH8WD1+hDU+VgDR129oPDLFZ0KfEf6CWUwa0pNpwKHibXat
fT6eI/OgehZlOFPjm7OHt4HuZsJtmGD84f9CPXPRaUIRpqS13eYelZ023114zDg7
SfWDdIeioPfM5gLz+sM3w5t8qeTnafXqa1Uac96CXn9vPFHpS/+BazglsGV44Idz
2fqg0v61i5n8sqLmtpmMZ/+GbQfjYeMqcfK4si9Mj66NZbmqnSf2RwwFRDp1I2j3
h++3hLPxjYtk/qa0f/b+StSalQLSJWVSdpAPzeG1Hhp3c5FWlTbIJOdHMO73TjZd
67SV335KN2spdUAgZDSXwsWhja+MX2L+MMKnBpFMsClJWfjuDwT1dxZdUEUnKOcJ
2AXOAnjlLTKaU1qvB+nLVXbpA+rPEWb/TYAw3K9Wl8Y7bJbDHZ1NUydw2eEtf8jW
i653btbyps7XG2nwzpLeTvRK5TsAc7n1nuw3zQmhMqZhNtiIe9knVWzLtbp3cTsV
pFy7X7KUBRo5ZKYyG/rjAAgRtO5J/6G6HVCkYnJNlwiclMLtDXqxtgnqC4fmOu7c
SV1eFpSTdBa96SzOAd4QMUavL1lW1xkYzGnmh74LJpBvFkMMlVThmhH7tc89eSSz
gqxS4evmk+krVFVIDh2MKhoMkxslvNo38SP2rxtoaqMSmdpMdQKJt/sIteqbi3og
fNRKiv0fkuKt4JlWGaZCeeZ7zH3C2vUjfV0OF+XEP/1XgDt0g413IkfsO4xW1aNb
Jsl+y4OD7DQvE39LgIhLr5pUPKO8aINOG+Vnsa8oQZlL/nJs9wI0uycwiRt51bol
wrN++vA92UfILbpwgIGXCkhGvRNX3XyR97CT6zfe3Qx8lTwXNBlo3f6/F68QHkZC
qBGlVopYg4+NtwVATfIU9czHqTEDUmh3086K/PmU5L1PrCQ0fOxQADnby3O0TR03
H9LcDy/yZJay9d7JlKo9TcqCHkHNGqlXGXBxqLyoGP2HnNDvfYIe6JfrSWN68xim
JZHRUrFf69Jn1accyAk/TU9CcJHS5hvLBYEABfm+Y8OWYnD99UmGZcxPIku/EN62
SAys4E59h9FxIA2JhEFTEsyoFkI+Hexn/WVwqRDZdGoiCmxmSgiQZvHq2gz+5qTX
r0pNvsnMAjQsLOsTNDLoCigIAMWoMw/TKvaRHjMeCGKRcgjqUUgagtTjV5hZXhcs
db0fwycuIsuK905PuwGeL7hW+xw8w4CmtzevCQ4KlLM0kqNkfXAkAP1FaUNWmUSm
AzpmB9FRA5KijQ2oOnAt/3yb8+Gg45Nyy6cE5xRp+ovVC9Z7Tiky50EW7A3yDamC
22+BOvzckG+vyyIjTzuLGLDaCKckKmTULINCVFjyCDiNrk4iRbbPSljAfYSgRgic
ngwyJAtSKdEA1hF0VnPiF3ItKllvyC0ltrf6WiWLzBGRK2mKZFIKg+YLh0RBMIqe
dKAUBm15YDVb0s+XPhKlQDUVoIBu5CkPo38qh4Cv36/8FslvfvTlNtj8otKHgVpg
1mgOYO6e9zOJs3MG4VL7b1Wy7crTM7Y2rZZ/bEqmCi5SqqIt4hwU1G71pziEnh/V
7MfizQVM0EsOZMYCpZjxwwgZUHKGs1AXodi0cPwmVEdoQIxSjpv0ImzOrH7t6gtk
fc9bstBMLiW9gVoJrHEcceA+weBiqSc9cS5wqq9oeIoIf1dos4XC9fgUZtyNWoep
v3O+AmIRtHSOGOiHU2fkjaj8n29I7vJwKiYEK3sh4ty82kmPFXh67aQsy6pmc6GC
S6xnz/EXQNnmRCPBusbTYKm2Y/vMyliwBW3s7euYV1cjqEC2Qccd2kxMRj1Owx/5
jJFUrUiLtCzbDiuVbblmzyR94mNoeaALqAdsiLIiBHSfSetSbytPLZuzwp5tkgaq
EFONwKJVfd0txndAB90raP09LyR7gW+fjYXnPt5Qlmubk86Y6erRiK65W9XBTA2V
AbUpn8HPnYVxfc2zNisKJHIrzp3Ufjeez3vBuKczbCpA1ekqguODqN2OrIMDrS14
9NdkKX1qqb6pZbzniliaCK+P4j8xdQOk8Dw4NxYDgxstfvMsUw6NCR9+lJECJ1j5
daKFHvkvo2RQF/0TgR7kKryIPm45yc1UZHUl69yQR1JezmJLp9LDlnwfqMsA5rCw
sV2iGy1HhKVf5N5bKOpR3IYdPAYzTHdM5CMo4EiggXdGIqQoUWs3L3pjVSGYh2n/
TiLsO3lJQbNMmk/Itagpg8I6GRm+XKo4obRhLYsorRolKtklxzBD6q3sxt6er+xD
s1dXHH6ChL/07vDjukynNwSQOmRUMSQ9oTYG4QXMaz9IXgyFvYTFfg2L3QHaYMIZ
oBHLjexF+BkLgBAxAWZpZnjAuT2PpX1c1+WLX6alScI8h6SyW/tQ0dIOipR36/rZ
mNFOELbDTxqJWVJf02X5rq+8ytFylkMSb0TFNlIEmQBFkRVXPOk6tILVj9PwQPP9
akhjp54uSSJCBPRLevN4O4FTuf7QNtyXZs8NGSDlqyN8bPNXJZlWq5oZaWE1kaSg
eFCWg+CNrEqH/Dm0tfKWstMQhO7JgyyNuYp+/ZI0FrLr+U5AT+OV86BytXPHwCTS
48HLr20bM9vy7ssfGDzsgacfdWPJzd3kBYxqIcXVlJCZL584toCAesbVvcLiQQVd
ljhyT5vGskTd5W8E6esOe/uH3KTZmlwvsGfMzsSI9mY0xk+xxvCtrhjPzN1kuSnn
UUXtRaWd3Z0MQkT/8lgVG8ehuPIXYfIILRz7h9ay5b3NnSi4Edyk1uKQfMydZLef
e1B65lQ3w1r1h3D/Fa9nsvw3YBhghNz4QO4LY79ns5BynaLSWkmHO9r6qOc0xLJJ
Yi/Qzhl5CayuC/3rdn3bsTulP7YdcN084jk/V8bu+Mn0yu3duQm8MVodNZ3elXkn
pZkBemPXoE6Ha8sHpT+3kGZW2u9F/dEwHbE1OaO5N+COQ3ielhwWZ8ZvgLp1uANR
iWpWT2Wo2QU90fnZRc7o4jTvhCCKyKgEodr943+43oOa8nyDkdc2AxvMPXQW5Vlx
fbLgV+w06BBE+wdrgi0+giGhNEPFLknCJjS/7Pjvi2ywbJbQyIDw1WnEE1tmm+Nf
mxLyoOoI04r/YOuEjbxaXyawsiYrj3FPbjAB0Y3yQ2pAR3o7zNBReEG/87ncKJcY
Do2tz4ZQ8HxER5m4a43KpsvfK5QQqTESU2Szdyp104tfywxJanckWAAQ8jKMgbrC
s4KGIzh8j6HiqR9cqQWtppwJ2Wt4SxL0Qm5MMNerT9MQBNZ3Iv+vEJZzt/vcpJPN
tXLGtDGCmL4ml0IUgXb4xdywoHv//JqqwN96JN4kfD0QPYpeMod79J3i2LplX9IA
xG0PnLfp0yBoINNzDqf0OiL10LYx9j6fQGIZTVvMjgbG7J5ch04yND0b2l2IFUL2
fEIDORPlrcSK0ZjdmqK19/zuZWBcvA+ypqP5tl/hxs8kUJcaVDpdmCHaZHJotkgG
opYqrdGzJk2ap8HZQUSqRkQMF4P8Ejv7uhPMU84NU8Ou3io3x3Ud0SLYZGWlfCTn
qtPoJgH6Wz2NKTAxcudzzSrHm8bHejvr7zzgv6psfM+KfvvW/iuL36pl8HQJwPe7
Uq0Vik3Ns/kf2uI8eTUyA2ZwSuzMcyMZp9sHL1134ymbkmlSiUqb6aJCGcapLEc9
TIQDr9GpsSWhpUDqyKtJR5Tey2fBELb1CyVQU/aR8YWD9yU5blHI/aqIgg3mJYRg
GE54/acerauizG0GUh3CUMhLD49PVWyrS4LGW2/KwzZECN9of5AYaYrmY5LfKmyf
0OZZnX39oNlVh0h/rENKR3Cld7SKxwTs9bf0lg8p1AUnuDhGeXMzUI7OxD8zM7It
Kxf/B+mzpST2cSowLLNZWQfikcs1KBV8YON3jZPuKe5iznTlZ8nutU60A1C3nJDN
VCq4YQEvvMA2csmgTDjqqgcTJSP2cbSzUN1zI7/GCm6NJfYyxKgBIbmRWP9NbzKs
RjKVETNedPuj30zQM2mNEqCDB9usvuKr8CCkpNcIq/BbE97q19wNY4ulk1W7kt1O
X/v2jGAwPIscTqyKLf2BcRS3rPNbFOyeF8MdTxBjIR3tj30Ewm5yFP+7eOQGZkpl
AijSBt81FH+WR2xiHyqOaBA7oBBs7tOhrsrsmHOJhjsVdW85+Xec6ZCXZK+nEntW
CCV9ZB2HD2qlFqEHnSgkfHkKzHl9N62xHDm4ExCoLTTg1RcmMgXT0x78qiwRmdLA
fcXmZ1mCwFpX4js0ih+FcnnlpYqjUhv1FyYVhYRDWXT/KeBpL3Pa//ahmqqB10rY
2uTMESfklLjlwSxhofNfKcrQnFcPMLs1qgDhk4etYupgNQ+UWX85qQYp3uaye8bN
belqVCOpukkClvIY9Ga9DFpNCgtp8d12RMKsGCoBhro5hsp4uT0qN+5p82hsppjT
msBA0mv+e9Xu2SgU05xzkJjS4RMT2NL4vQ+n3ekRZKtyaGc0y96G8JylYZCp6Jjt
9A0Wiu0OWrqbmXhVxQ8kcC/mPe70VDTvAO6/0vxi08Zvn6q+N+1hfa8+39L4vR45
ZeetQTwg6u8ga/gSiAJz4A03rkfTeKkbGyMTEkZAAuX8ZIvCG7+QfCLVbAtrIELZ
rdQJmL6DDuoAJ65CJMX0BQ0gzlw75r+j/BClnoUQWmn5qxYBq2+0kVEkjTHAWWs3
lTKlBHfwzOZ/K3zB6xBgPv06LvWpTJnqsfaF4Mqm9SSZDjI8gOHBlqXs39Hb4nZa
wjTcHWpOkHl6/9Q7GSMUUYlekWGNb0J44L1DDawZEB/+gDPwqtP72ptzX93Z40mc
XbMgrU6klB+9yJ1qxF3/xtFrCMVy8WQMy3r2Fwxq51lem4MnuThX6OpPOsaVhdCe
zyW3qU2Re16wdHpT6m2mLsn4ZjosS3lhy6jZJ0w+yJ9zsLvhUI8kExOG6bLPalkm
PBZ9PeReBfVIV2bqk9rwzkxnNQVgyKkSm5Co2VHTeYhOHNmigMlFWvZznWfUcFh+
ei3GwImF8iGERAwQf0zbS+FqrB/IhCqaSDyis8UGOcjNe+NREgkPj3qbjfObQwMQ
qXf5EyyjFjaGxPN1OcueaqT2z3C/BcfazbbM20D3qoIr9mJU5a93zZ2rd3SRVtPj
dOaBtYfVhHqTTQ1ixBd8e7Yi6ApIgxsvginSgloXP187+U7vqLhPE7CTsmdXwBzR
FAvXi92KxlajNz9Qi2HgiQwa6sa2oP2zd6xISH9cWZDWzwXm8U1eA6ms2HobvQT9
5mbcZdgTmBZlOtc2t/sP9jF/QZ1Fy8l37aBE9DimgYXs7jxjdDPSUJld+V5KjpRx
aOrpR9jZ01S/UDx6sc0En7bHKye27v2FLGZvQnokufWF8fRYr0VJWb6jmokZOSFc
Nannb2nNLKUE4rHx7wmH+3i0dEXVMkUargN/gDOeJkXQZb5mjZudBODvs49ucZEw
SB57pXtGCDlz0UtE5kC++j3gZEKXRm7pw3nDqJdANqsndbKZrq0gbEj+EWM1nSj2
ROQ8/ihd8L/dF/fg6EMNUwmI0Izeez8zJk2z1cmuXxzkGzdnvjdEVAk7amQ0pZwP
vGjmi+nXumo7JToN3vBKhW0F7vjuenn8/HK+ffXg8QtC+mK1Jjn3fuyjId9Ps93N
r/R+znH3+FTfj2i7eBpMOI/l8bBoG4vXJ6vumf0XaoOzr5toIbMZN1uHVHnS97Jx
QWipxFnMrhde1F66/PNu3Alutp2K/BTUXbg2kmYxdX8fYFmjLgQNEuDYmYDeSVPa
YBOh5XlmQRAnW1ybBrj0B9UoTFrvoKNd/kHhOkDt5QtCjTLvRa5t4WfrPB4BITCe
h1d0LBf7UB+W0E1UC4ggE1jl3HgWZVNCOhGgOECrSiBlyL3rvzmKlmGFZ7Oq1RZ1
OqHVgZeab8MwsgbBTR8tbnFIRnn671D5JSpALYaVucw1VvrQNaxUDdwgeN96BsZR
FgDwFsCb1RCtum/0YgdvN3r83qwcgAJi57HLwR6mAY2/oyCnQ8v/VgogMMaqhNYM
A4hrjiFUNn/uWv2SY2kH+OPVafePpUgjnI3W7YTfJOOgGuw9LcF6Nb0b3TL3hecd
g7jmmcLPCv/yAIz7P+mkGFAGh1XGh5jxBeFcif45D4PDV9//B7wSaszfDqzsNvv8
6UG3Rl0P/8cYNgPoPI2nF0KgZ7EIT5pTNFEDjKp9CBO6vt0ml6FElYvtQA520Kyf
B6Zym7++QkpdEMbPE1rTY427ap/MYglt8HcXVxtmWdDMe670MYMFT97xOv0bf1e2
VACGu9lX+aCEPCNJL+n+Fjatm2Dd4eqs0OQ2QqQxqMN0wV6smp1N3Jf0b4wsieNH
H+ZEjLLZPhtuwqzumgWeN/BrFd1FDlcccZM5FYIYB2dBZ4ptixIXtdHNJlOk4LB5
NxVTz4licDCoasL69XF4m8WaW42fOLu8v9/DECFIV68/MtHxzoWvlWtiv5qbBNTP
uSaGPQZwBQiiEiZDgvWwomMyaVIv94JKjRwmN5IdPChfKKp2CKELPdRO1JK934RX
0fkybCY/3GE7v3LcLozOkEfLK3M4JaECqfNFQdLiktgnBQkboJoIeZTinREtFYgM
ipmImWJWq8nHVJfvndZzQZrJbQksRN2FJoM8rpyRde3vWFJ54np6QZjSsgHTmgdp
fCs9RKJuuxmmT0lkMumq7YkeoUPfNWnpXhOiphITfakwfGnbEVIgUb6u5GRB0fgQ
av31DC8eW7bJNbEib7CzjVB08pwJcCL9jWr3+vlZTnFLVfcneysNQhioZ7ooG2bh
Vccrce4gXhHtQmK5Re+lNkfI4Lc+FiM1ZBXHS76N4LioAegIrT8pVAVw1s7XXbOL
E24Zvy0MHlRQ10ZFluF2u/CCYurTS2cwpQaG0d1iRrpWSdWcnF7qtoV/PSdRqGcB
ZXV3EFL1YJykTzAaaSeLKnp7L/BSHc4BuLw4ZNodx8Oc2W8+IbBI5ie9Ziq9TbZA
WFBVVpkNptWhBqE9ZPSZCp976N03gsUyCsSuSwuwZyh0DQjkB7+O952XZvgkS6fh
se/7Ox1Xmu+KBFSRsA7s5k2Ufnxi8HLgeEM+nkvX5xweLkzxRTo9p+Es6x08/Nd4
lzlJzPmFZgwf93y756hTlZqCyl+N0cMaKZUjYTdBTRxxegvn00paaT60jN3BkwEK
Wu5YZH3riX9i4LrTDzZPs65A7/hJtiUw7yUdFHdo9GxP2rlTaEYuyo/nuLs+ylNs
SQZiEMdbXj9LRivj3XN0nZOKpetTN+yE5XPPfx5FZ1bE7sI4XRRRM4Y18kvh4K0F
aW8tyxNWluFf2iWBxgC8bUIVCBENHFs0EjHQZuruQZgkKhfp8iTRMbq/xHfsO19v
a8q6sST8qvCWGv1r4YAypA2mn1OqX9eIGj75495h+QjU8i/A+fZ0fhl18BntNvyV
FlkqM8pKBJZKvsoi4gl3uGelhoZRcIfFG1FPi2DLy0RzxCsOxk0+WqZ8e5zQpPks
D+KpH13i2cJ2PIGALjBJA2RjS83Ic+6tjgjdyMY2FxvEQizU1+idHJNLigVnDDrR
WMOpVgia4od7245PxIXNbEytEgEFA0RaFp05N4O8d3KVm/d6wwBS32W4ShFoW3WK
23LdqlFW1Mye0dtfcTha/3oG87Li6VhDz0MAH+bg5DwlfGFh0e0prnEV9Srx6OKU
lKD5VWzPO3GeNaJP+mzFKkbhfJqERpCjbAUMDRPVG/vUkKy83Bh3bqHEiYon0h4C
/UaIQWEdR8KqKeZLqM8Zi65iixYVI8LaYsTVJ2WeJnE6+uUngMDa/HoES2fbe2e6
OUqlFjkEEs/3ph/FO79mphgJvWGUw1I7EihN4N4JA3BPhftb8aHtaRxEPY2nxyZ/
mhEJ6E5UT9acBgufJhS5aKnTE2cjSj62AHGr02vymZ1BFYNK5rx2+0tBPldHOSHx
4yTRFMudB/PRAPFN6GBT2xan9mtz6ZGrXwek6IFDTIvoLBkvtRWlC+p/UVTACyI2
iofKhRTd/WLWdvVsPMfUhC07hLPiZ/OTKJLuzipajIAGzaZRI8D0zurbedWGqI+c
GKGjtNdJ3i/DjSWCqxdbjI2rkyAmIFWIhFQlHTp8uVzKL4qKPnJOxoD7yFYrzu7m
0/OYIFf3D9gBCerxzAxY2636TcqGhV/BJNql/uS1zj5zMCkTqU5Qc7l31V5CvKec
0pasEfE0WueikNZe9m/DxtFZd2Rf3uan5Ji8E0tnzrHfvWpyxnXETAxpVGcJqWyM
fU/uGBH0NljJFiHzVRLCJJRTM1E5rmN/+RJT44vxSly6YkpYJNc7S16p9hijE2J+
oS/1g+EsX872hqPn+EWvjp/WM/9Ucnn31y/lneNR2eGs9nfWce7qdqjLgctu88As
8Vk2RySivc3n0CFUwfwxt4pQZlronkESRZpDgHMNFhz4lkJLA8JkiSP/DXXe4OgI
+qqXMAzeZ6Ci3pJwGt+vYenX3/1pAfv47pD30hLMgkPdSgtQZ+rcnsPW1mEkWO8/
yfz/GzX4oYIokkFmFwZBV5Z1l6hJIkmsuv0F4HRpwF3FmeVlfG5d7mEq+qs41cnZ
m3wCx4XFln6r/58TTRMafG7aYmG+rboS0CeCbmuiOMAq02Bcbv9vYjzxYt4qg2cY
/KLtOEKtTjvB3Der5sW5qsqD30G6pb7Eg/ZuA5qYgjtoXBW2jqUjU/aDRG1NuHDb
mQzRsaPcCMkCIwUhfVMmAHicNcT2QvqVR7YyHPwKdyP34Jv2Ye7+8PM1dyGRiONF
xWdu8YXmIQvEnlOvxtcqE2fpiWFN2ASRXKxypLMgw1A0R3ZYUT127hND/3oTLbnT
6s9qcgPk375x3xDgns2edONk+iLCYEACUdE6P13hRr2Zoupw+zrzrgzkBsSwYfgp
2wVtS3jioYs61/8rxzzPZWtPXSlWNO9YztivpCpeezrU5Pg30PpUfvlkiMlCG+ZQ
XzVdMi3TJFJvIultN7ydv/2ldf2b8O/8gytZ3zByiheh/CFAgx3lUYi4N8xdOg0i
zfFxpIk6IIyflgAqSAijZc2EeZOdAOSc+pTNadvpewazZ51KwrgD5fS48Nehp0yV
pCW8Mdub26Yz5gqTwaJS5xQXFe4p42bFCpnBH411e4fnlN290nJtAKW1A2A/CqZi
BAH4E9OyIC2TSTdulpF1X4cGiu4Tn2EhqgqgIOt3yowHlrTSob1jc9BhX40+bW4b
wfn1kzXVRHLQK+IwlgzXdZguu1Ooul+DitKWdwGvYEr9i7DmsEWT1F4L5lcyN9Zn
2tn+JPyol8VJuZ5+lRGRrb3u9DxUY/s4M9rGX20iLCUPqvysQNjYPkXuKgNQnpXn
rGEyywaL7Rtz9wF4tT/Q2RCipugf4eTMBfXIeiPdOdslLIR572h/sgQlX7gR0272
339rgN7DJUJ6XVE5//3XplAsYl0ITya/bWI1gRW4wWunJO3yL63OUxT4XKTkSVcy
rQSSEWUTIChZx0L50EhJDRTtNZAa2hP9xEn2PS9N16XbxADY5jUcusjijgQdGJoS
LZ1XgioAOG9Z8CwRoLZNl5Dcx+Bqqtq9lr6g2lMH3VfMCSej5i4kW8ssWftNYZ+V
FU1uB5lDQ4/C02mGGKC6/5AxBqBuyUhff/ONenfgkURwYBNbt1/+c//JQyX1MGYm
BP7DADsr6KrGD2GRGwRLQI4/WHQ9wRBd2CACLiNKMx7n8tDmeifeC/4beLwxC+cM
PfcfV+PN/ng6IGj9mHuARjmVvdQ7yXZLeAKHEmcPmFCFGinuoL9PH6CwqZjtKKHe
fwzTO1HaV2mLQ2VoE5IKfzZB4CY7I6X44x1st6x2rpJN/bpa8awkoDk+kAm9tuEC
3I7YV6asNML/NSqS4qtLgTceIb2u/yvGRCMV5bHQpevmpOiXQPLku+RMYie2p0nQ
6p1PF+sfb2JgeHKN9neQxeBtgKRHaDta4gqjCv/ThB1VqsstTqbAWvWzBXjQ+a8s
HMrRWQcB136sgM4MAXeL/v4UUMo/H2pPlEslm/Cg+RzF1zzOlmOoFX8gA16k4+bR
njhK2WV23q03BaN4hEuUoN4oBH697xfykYkPdTDyYhmS5GtTgnZyePGd9UFxT9tG
iWiDAdat6ZPX50x9NnvN1pzaTa7fIDD09gEN79a0ggsrMMUPY+gUJ87C4v4njQxZ
mK+vUhpPDiqmRdT/HBoxVvOyCykjpwt/OaFTTnqivzmAAa8n25hhmj6FrRHYMFLA
R5oJ2hdaS+MhNQ4NLo2XzOCDhNeVk6eeo7HbVczVbiMqI6aRQzop+PsTt1DOWH7y
OBBpveaDvQtbapgu909/Dk32FQSfU0kXypZ+Qq2/fhaDxLplB2WqWzmWZGSJZsor
UyC/8tTBSXiE4Sld3KF6Zp7zr0cMWgaWqXXCTbp0t5h9JpPZXKUeU+cv1Z0zoedc
1YMOfgfJVLcuqBBil/flYGgupjZELGz+Uc53i+UR6iqLBimhM41N9ck0L7/kb62A
GuXWEhQVCqvcGeKyiWPXQlxOAOaJKwUDZgdYaFL/z+8dfWUItpA+COWnVQyDeWnL
47JQpAqkbcCYlX2wfYZVJkBx+OVyU++V/WSsGl51FTJ0Gx5Oa2VDUm9fuUUAVr2j
yt7Ss0dfb8p++S8gifLYGihso8VU2yrxe5T1aIqevJzDJCr59IsjFfTEBMU9tZYA
fSHKJoao5gQUrjsMh1Ep5dlimliJK8k/6oSnOOi5DS18so9KD5UUYQyZMd6ZU+Fe
Q1oX303rQ+GBU9pz+NP6EvbDgXUITCKJFv04CfIlaH5kQCb66ga/x/TNIrpK8RxP
33M8YaZZRnvuXzWcOJzIyjfUw4wqnuqMokNs8TCsx68EH9ZKQa6ikdvDxM5fso4n
Oxt7bANHwBLNm22Isnjga4I6L1lzBhmPfov7AeUEJhR/bFTXdh5Yb7FfGEI7gKMQ
ZSfSk7py/3EhTqfUIReYaYow09rSNO8M7rVQMUOrdnv3vk+549L8541SN7niUiqD
OzfJHeE3LnqQaQonQp0CHciCywXQ3Ja0Z8hSgMo3fDMGiR+UWUQSPO0uApM6ktlw
39+B64kfT1Ev4oL+G+FNA/WjtxefBwkOqSFdiJUcV0dfzSjyfzrV7y/R3UcQFbRo
jj6qWm9mJPfzE0TQYFZZ0yWqo4i5cOzOXo6VbD5blNNhuODXMSW1gGIa6k0spjkt
oR6oktoe1FhxKALGzmpp0zaiOFxP/D/toHVgOl1lHOdauEIpCHS19D2YAZ5+fmnb
qrVDuTOVOwIDzeqHI350v1AKQCjP8GbafLrBl2seVsV0TA5XJtpenmEdweJG7Pfz
NVIXXOZEZfz56mlQusbQrH95ju9I2QFBHWC0eNtvudazZhIJSan23BPx2aaa/g45
+dcUzlu5lijFqZ14FoDyVnUTks6yNySq5MSlZhVbBb1CUFOJmYgiAFY7sWgH9gHY
BwK2skYGYQpmIIKFxv4uOOsXJyyFR0wWvD+LB8gKlrBiQWg0AK566jZbTAikuGXT
4zIBj+oMdJph6TryLpgmBEK7pzz8vfMd++aCZcM98erC/G1MuSoqiEvR7UBICh1x
Zv39+YegdOHhcF3fDHwoPtqYt6uqCGg1xrfjy9M0C52rze7OdwwRQhUl/GGZp1Fz
N8r5zK7DmiwMl8yCxOsvYnfC3wkgwxJuOLdqQI0eO9BN0KUXXta+Zzkc5YG4aJWu
S6yzfYjfFCFktmMHu+iyyaNYVCGKRyI7hhE94v+mp8MqC3n9cCalQA50rOpgL+Sj
+PvCfl2bZYCKVFX8fjJ+qX+hE+5sLRa5XGkqxDMNx4pQ9j5j+2FgCGo1VsK8MAeN
+fs6Nc5TWG0xFuqkNG2zzzLNQsEBt1tnyY9ZIwmm68z51xy0DHSzkfY/3SxgYv23
d4iYZ/Dk4akyo9JJjlwvJdGDBGcZJuXbvvdsfbE+gDYI++wm8Tt0UR+R+3tRNket
QKzEGPCPhhXAeNWP3ob//DuEnCNkw0oLhMyb1tCUqUdcJUx893UbyYPIJ2lweV4L
Dwh4sCuDnEhZvgA6yC4EVDmo4vW72+FZPdx890Grt2lFLI/qdPApcGAQD8grLARt
UwTlbnbN0iWA5Rz4JGPr2aLsDlhawg06n4IiRAXfb8PxY0wQhxMcuMwNIu+sngF8
ciMpTtTgQxkefFcoHxJPtJw7FMaikLJnOSexbyE9FPtgTpBLXiBMe0B11VVrBrMX
tX31u9Gf906/gQ5RqBThyjNLHcbttfP6JFGGPVcqkJVHsgVMBM6R9mj3ptxT7O7p
2UrBFsxPTW/uC20PID+nNHuq/PN7lbz6Maail4aqGCRWpRdRIsYGkJwXipeVlBLD
g0ODoGXEDrqsZT30xjO/4NvaiyI6fVRlre8/FO6Rt5/OyqY3V29AU8Dv+64o5eSV
VEjiIWwCb1hjFFQnM+usahmNjrpmDPg+1Gvvtmc2X+oNJ1Xzv7EpAcaZBLZojmPu
KtUGNw2rH2eVVfGdzFtmfhJf3ZqH0fl7kErncdUoQiuW6n/Ch95ceUhnlRy5hWKQ
AI45So51aTlkoXPzuz0/zW8LEy4lGHC1QggdpSyOV22pZ1Fx3H0aED5NJuvhxRRI
zyhr6D8W1cNRljFtJFZqRJ6V5z2IP+DYGqEcvkTHZ5qpERzcinKHiOQvv4wimFce
k7YsnIB+snmXUAT2EyMMxqiIef6u6ls+KxE+WanyDUfcYBp+awJp/7sfd/LTzH/f
+Yb11OIw+dXxfWOK93LERYR6/3228qvWcBG0ztQ9Eu/+yObicGfg2C3oHPcvTDzS
DHIe8YiG81GUouGQr4G6LegIuQWrd0uhkuwMqivXhlGLj9fr+gcX+p9MeJ3VMy7P
S3azTEttRxNe3MBdQFKJWsW4VDlEOo1i6TvC9JS1hhdSWjmqUwyRc2gmZrv9ebnJ
00cJZ3SSFEX6Bb9uX94gERC7XzXOLA1hbScnv5XBGPPb+hjhgPr5b7z6mF57BaZa
GbRty7+4gENb/LvuP34QYpVmwdmbqJ/H8bdTKNhd2Bomcso9upbq8EwGdCuPG+0F
R3Sj4DPBjX96KOMr2eLJXFwBY6fFNjQNCvJTigwzgljIrOxv3ezD4kc60lr0WRb2
lvvgfNsoO7raTWNzl+RMy7T1VeeQY8ZUyI3qIjIeVdb27ph4dxx0J0mKwKrLv/wV
SB7FhIQOt60BaF08BZ+ktm4o+FozQRMqxrsOAsFOyzgXUUELoMA6fcRhuxKkF5IQ
tgl1znG8Xut75vxAscWFf/ymCrWqJAVbqwN2ixZsxU2TtyvcXRTXOE9iyYYxa8Hi
hwkjamUErS9OT8I/pz9bVvC/+2QeXTO+NWYFtgyyCl3glOFoJw8Q2vLidOy69RzI
K3YK6MfQLnbc9uFTfWzukTZjeWBtSleBdEXNa97Vn8dPpNmgDp2G8FnhpU6ELuve
I1vBpINVFHXwgfXyfj0KOKjSu0HRtt5rRq//Y1rXaJJKjPEw/ZCpAh8rVwReq+bH
AKdrCwHyx+/d5Adn7MhYmNRh+tTdx5OPAeof4R9vXjY8GZMj1yIZostgcV+f7OzM
46aaavFnSIcwIpGEo8QN2LkIMHWLoK/FC9vuYr5pGRnbhsget9wyCfL/oraarTB/
uFT5T94GjxYNKTD41/g/dKct8li00WD8XaDQkiDhcdMuMtJZDciFcJs/z4jUgWAv
k/Y2HOoWDJXY/ELnpAtogceZrCG4d6AvxgqYKF9Hqhz8oAOAl77cVtTHsa/1+R4I
EWhDOeuUrC50RflswMhDeTP1joJOsfApDU7x2OSWR8YxWhovGAzXdZt9xZO3Om/d
FShKUvAbWulShu0lvyM4g0f3YO8HsYdkxuiwIU77Q9sARHyk5HaZwG288mMDMDmo
jAbwQIZOOxCWeSw9gi36XBvK+q2LkQGWec9EEr1k3RypQ0VM4zsDiNFaGI5CNJpS
pa1a1hJT4ORXzQVVPSWcjlI/iNvkG6eIZQ7hHaaR4sfxEDZVN3rCt4EZKMou8Va6
vmF93EJByP2MzbRwZG94WfTdaBapEZ3W5d/i1mWlBGsL8JvfdiuiSnCZzIyPRMaS
rWIIVGCEEGs5jmnilGEgsMWzB5C2cDdchhz2RYVgxoM6mni4jne/tqiMWTUWXlge
zDNzTltzqDhXOzI5FJEnqfdiisoWPCfRTTGrzPDs9MiyNftEDKTAUxV3HbjH9wln
Gaa6QHcMCys3Ksc9OT3sDAMc9VpuIeg3cwnhU97N5EhlG3/rpOC+FH4VgY1FDHsW
yTBXlcWBYC7sXoxyMA8vDz09dIFGB1EkMVHD6fyQuhhEP56Dpq6DOUc2X22f1iEv
kDR+1ibehNRrhVldIQ0l5/Qs/H+1ZrDWPUz4y8uS08LobpsnfopQMj3hqoxKELFl
ZVYjX0D6hOSKN55GCJE5mqVgJV7jOtflZSjoe7hK7Auu49ercyDthX7yxhp3dOG5
10Kgkb9+PgGoXr7P9dAQeQDjPDN/QkhDowJYoj8gMDIFbINFbXuHsFQO838193Pd
sDdHL82Qkw9WEg7dv2Qc/HsHavj3xz2qlbsF4ubfJvtT286WCKfUTe+Cyx6QroUw
+rO8inIE8wfNIC9nNlKbg2mQeXVGTXyuMAuCn+WzQsmgZBUodfHs4kyhlybIXdxm
vxb/Vcq1z7duhhit0FMHAo7tbSWh4WiWyTGsguAtmCnTXy1pdFVl35VIevEBRESv
q4IRK96GpVt7rEGM5odHeh1niOxiZksBA9sBtgjFW3Fogyeef42NqcymIR/wUTU8
n1QUmZ5fuNzQjXumzwiQoZURM1ycXPjAUuRK2FZ+9QvrP8rzNyeHJ9e29k/n86n9
KfdwLf6zaE1ZQNvuA9N/PBbeM7K9lwBwLTf6vnKXwryvUpa+RfkA/M0KOLaFz7m8
Gx/dHtoFCce6gwUnbXwYG82dEwcw/LePSCYENLm/UNr8TtS2j/M7VJ3U5vuh6S02
/M1m1jGz/I9MxbkiXAjJMizZEmrgaJam/sEu1Cuk2fMDr38LkZOSmBwS0hPVLikT
p0mAVkPLFwE/5ORTlK4+m1aG5CsLRJjmToskSUzalwyRyynJPUsmplA68HXDD/Iw
2wpt1U4tuIPu2WjCyniGORCjwesfUJECvE0rsNxVZyYAW3oIyfiMSMnIto3jj7C4
XCm26FJT91VnbGVAtivRPP2sUbFjdK/QaPoSZRSHykXJSW09H4yfucXP850TKGWw
XyKIFdK0K5KX/PvtBGJGInppn92FVfQlM4XWFcwW4aEcZ4PPM2d5OuwE8y1ffZj7
nh6yL8328QhI6Zw9CuIE7m6myeGlbth7UnPNUj9kTm6UsC1VTMOELuv56weZ3cCC
D26mvUNyIALnxIP24tRgzpPipu1NwiZrrL4+7yjadLHhxvYxbPd02n6WpRTG8dyD
YdVdzrQ9l0ZrYOpLgCZ/V2MNHhZnB3qVLzXisOeYlFeNcQ3vLeqbEyxqNT6xN0Ij
WZsdOwF75QqYJxSVS2/+Iy7eBSLzm6TvlD5NbSCfPyKDD9qb4zL6KHpi7TclygIA
LR1ULZ8PIV2on+wm8IKDIoCs8jB3/dLuYp53XTMpIVGpQKBiCx582Pl5QDzlIwp3
c18pzbPLogCyqjjo3GAu/15ESAu4uuchhALhGlRIzzt4a85c31jtg7ehHhmCDkUt
JACj17810ilFF+cITfkZp6d8Lk2RgBYov3BAdzs7njjXCm0QQxRnoi/gwSYCyZ7a
w9Jnn7AgX42Crf5GEuo9F2iyaqg1Fk7gl74XrJE21YlBSBCh10suxCGsrDo1N8x7
tAUdR2VzUuht5JLWkpaMeQoYhKpGbQjzbL8XcLg78yWK+BDTn5G8c8OMcDAh1wth
RjBJQoFoHL7D1QrdseRt4kzzq8gQEmcx5SMtP68Z9/OtOFtE77MnsnnsTbenr8sg
nX3whv4LIyySk/BHlFBdcAK16cCQzhCMJshVMQ0BvZDOXqpSarTGQb6Xf3IfUyee
tWug6FSv+FSDAcbOHz9V4KdDXMcTem58W+Y2Wf7AxPmUOCjxIhK/T5LqAx+Ebt8S
ei1X+Z2JLugQ88NxBOm8asABq8HuW3kfBuH5TcaUlJ+/LkCISypGfittOsdTTOcr
29Ox1+wN7VjyZL0PHKl7tm/ClglYwCR/wKUu5/Fzp9W9yKYX6261n+dBenJyh68i
OE++t62ZEpPc8Clv9ZpiwQducoZsfvlFe/rATdr3A3sZ/AGlNhdJyb+PoLjI0wFx
PhOrCgjB2BE9jEgUsutGEM/RTOUzRLMz9p19SdepKKAgGhscX86J8QJmgPERIsMK
iZceMTp31a3XCqh4jEjy2gUsbOoNe+b33wCTM4I5y7nVezdlEfqd8Oh+MFyQlIag
rket6SrNQs5qvkDGi6wj19I3xdrK85IqJqxxzPGPA3Jc0lKvFIpLZ7RlSTF9rJzJ
wamVANdt5uARrJrONwdMLFxCwK1SrFirQ7nNx0JWdSGOrcZavFBozpFaIIyiBTmC
hRYMAnGg2QE6xiVZIEgmfdWbgEFx1BHQaCdGNsBYNcE4Y9RENB/QFasgrpEYELu5
AGY3SruPEyqWcpL64fCfIZkI7hudhRqTVr4r6M90r78xZWSrsv11wwnYdIRbk8hV
Jw6jrz/YLFYW9XfKBS9qy6ah5tAVeb1vZhVf5BqCWdPJXsZteF1mIvJqvFXnWIkR
GjmSigVBYmAQyy35IzUDqcj0E+VBWG8SAlnaNMHdtltTtkzVF493GPwD+Nms9Y+Z
zXHnpM1OSB8f3zkTUcpTyVBnYlqRP9MunPhU+g6c3qIhOnYr+2/efJY7FdQ7WmMf
j2B2DjcOpVfFkvuZEWhj5P35Eh8czMvHL5dL86vTTXFif0/LvTU9CgHq/qeiJFic
8LZ3dQ6TmFSs1K/oFEUM4fbLwmhCc2eVaH8X2kLUlBpKTtwA44+z+i9B/igwO1WP
ClecC3NH7t7uYSFsWGt4QDQwF6mwvK13eozhKQJYK/0X7qqzxxRaVel3pkXVgWCW
u0o12+dHAXH2ROyWsV4FzK8beJwZ4wIGYR2syFL0rKpEgYcONsloNBpsDg/nR63i
Z7iqNAfrEDs4gDK3Hq/ora07LD6WOS/LVs4oqf2YV7eLeWi7DkKS02RL3xAFkMe+
z9rHikZRTYNCzQAtFKln1mioxKE4hJQoLfMJuibF2vGkS94OUTD/qh+T7schXehm
XKb7zGnUi9vcCQJWnWJ1dTv6fHXag7BWPi0yRT9skGVOUrsarYjDESJbcMScZ4he
+LBaCo3bUUVVLAXRSav2m3AjOj9Hm8NRwGGpwW6qg7hYU57g7xUdi7dA2NsKOTzv
rwIC4y5GlGgrGX2iIqwcpsD2giD4/6y5f43I8HjLvp041Btb2J+vQqk+TY+aqnZe
W+s02edzYz3BCm+MspBypVH7nyZYPlDo1musBhjUTl/5vftGZT12/Xq9NadLHj2z
HH/txvnjxyHdefJGjoXJCoz0q9xrIthdfOu9s9cBH01c+Pa4nLl/J0xOTS68P0w1
FaxSpz4PY0PAvqz5kS3UljW5GjsRNnKtWXUtmUvcrNM0vKnf6YusPoPgtbXAggUQ
L1wLqnLsT2gDa0au4OFmEVCdF5VFRR+5Kij/dqRTjOqs5fCLHkDCxKUPdFu6y+jt
GI5o30CEHlGaRxviB/sKuogczO3oro2iwhsgfA18R5sWpBh8ysc1Dqx/8w/s4A95
QYqcUUCKNnajI4xpXctsLq+Xjdfwm99khVYhgo25qW5sztDcheOX+6+g6WnNe/8y
Ld651bauNG4c9ycAu4FIpGon/iCDBYMIdR4OLWXht6p5Roq+HZaxKXDnRmCUW1Ga
dwYX8V9dd9Egf7qPn11EbJPtBSikrQVH7JTv7bSdvarCK+zPb6vhYI8//hGJ2vTN
pjhAXKJ4wyfjFVR1U8xbUgaz8H7vrYteRTbKAAaHdB1RcHlnJAXuXJIRIsvvfKBk
UsnTfQWqpc3T93Evk+jyJf9bqP/FygBeXZ9LwpRTPpD5trvDbv5NoRVgqBQ7/0MC
KN+nem5stNfse2AtAf9NdXLtN1jDEuCjt8kA4sJMvbXSXckosCNC/okuuWq6xFYU
alci23scT203EwV6QAIcLHDUM5krVvkpNLlL4bIof/G3A6gPcBDgANK3NUeuAxc/
azVP9ytj3RBV3rGfGhNV93usl8WQO5lUkWbDMpL12yIrZxAFK+ZH9U3LriYyn9Am
Y2BRI/V7+SDNIRNNKSPM+Cfdep84uGtmqr6hN1lgWqrMU5eD9598ppj+xRNkv/TC
Blu3YLPgygW63NQLjfFO/CRxZSnSoEOiEnxSoGuaLA+KMhSWPGQzoIbdg2a2sgy0
j6feXPFqsHqsuqkvrAScmF1h/GLUALOK6DG4hQjnHIK5eOiAvz3V2kumouMaYM45
bawQyB7c9M4otOGuyCSR2BTM9o7LmI5gs5fCTYFRcd0o0FPcbhJLYJeUVT7+CaRB
6fS09msA4Qedrf177p064UlSfqxcNwK8DFEBKXLIp2sIQG3SLVaUl5tUWm5tmf+W
0AmqstHlo2aTth0tOGLZ9yfx03kyHdjtXQ+3cSRdPFEzxs+4f7ttMHq+Ev2/nfvk
aVXdfwpBZF/4tD/K8le5xRus1pNOjVL6UDQfaMCdbI6cUlUj8B+SMAnYRMqOy98B
HgOhQu2F+MhNqMPPeGhgsXNG54X0kDqh/5zXyqIIvKgOUT5GSKt1aFlADJFwkSlk
WRa39HgLZiWyaJzciSrSHNFFGkBD77eME0tQFejZZ/sZPuLu9psqWuhP/17s0Ebu
FpSiSS/PIG2qBaQZt+emSAHuZp6Arxvk0yPivwpo1yBg/ApA97gCMdWsRhj6Xzb5
I8aK4cAtE/i1jR7ZjWYMdt5Ze/FD1/zO1DLcxpU+kIU90sOM8iVVCD8TdW0Dr1Od
PE9BAanmdNYv22zbZ19IWICm92hc8iZp+IkXHQoUwXSZAZmXf6BJSkHSYmTZ52Xi
PBi+r8hQp+I3RrkuxHpGAgnpuBwi8RimIsSbfXbdGQn+LFsfIujNdjGXNj8bNeuq
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 34752 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
4NAZGBPmQSC1EoH0Jm8NyCqlPLj/T1x3yGUznZvPJcSDzBAzcFwqXKRpDaH1ZsLt
Vj7PZwMXoCrWz9CTK8Bc3KUzczrghOXYmwC8LOjbmsVXpGI1rGhG/OFRuWiM8K1L
A1bH6M7CQ/hdNmZA2hrnkO1xffHSLWp3sOoRuYuoUzGtqoiLUyU2dmf47X6N/M0r
/KgfS/okM33DGCSRGXD40+FiK206qal0FphOsdNwNyEbIzBpV07uJeFMRpLMhJ6W
LlE0uoYVnK8g5/KsSCy7Tcbm8897hMGLKtFDprC8T0qYZ79dXPaVW1c6VPm6z355
eWat0S0CQ2JS92rxmGytgKmp4/B0UbqBOAA1EKenPxOvgjexd6Oy1Ps6S8NTtk4G
Li7ry1R6b6uEBBDZGHfCFXtThiG+U11YgggfZAp2C3xBojf/buIRcWXrkVm35CIl
qcgpifAt411uA+A7avqiiWoQdKWWdHMSYVAWaGZllv8Zy30ZFl9Qz4nEc0nx3EkR
T5BJ4Fy8ukZ70iariokkxiBXEj8sBskjCO9zYDBYwcDjFcE8IR9fGdRgegDnsQHw
fAfTcRHj9n8o/lrGe5hCv6XaTHwURmHgfaiYC9pl1wm+BA9coyTTgy5fVqMJSD17
ZXPGEZNDaLbkk9KnxvtkfmGhe/t6GWBeRFGN2wnLiAoe1CJB+IbChQfR+KoGSgQm
JIMHOnc3M1oDjpv60ZmM8hZVSEoQg0gtR42paIDHb3fSWtSbBNf0yrAbIoZtUyVj
TgQvXgo3KHe/rlGKbnZqqPEuYSHqY68vdFvQEmLu1G97w+WcYfFfwrlwkTcSSBYa
oFo72/WPGsJu5XP46fuEK7M1YTY9JaxqkNhW0lHN2SkZ+UfF2o1vxVNPoPCxYk6c
PpyZXCPN3fuCvXaxlrFIWKif9VfU/dz51g/cCDob1uFnUm33o6PnOPWv9iJl3x+k
paF6vQvZyxr8apd6/6zBt+n0pIh/7KV6K4KqaqTrePFTRwQOiWW7ACfBO50JHGvv
GRhUQWk++tTctkT4bkxdI2x6imti37uN81PmdrYJjy/anvyfk+oOIhtAPKUjC13p
m0WDY5kLQRyOlQoyUsN2iDJCBLvaNBuitFBOL3H0FaRLIl3qxa8TjZof0dbxm3x5
UN8zFCTCxjrLsArYs0QHo8/+o8kYaFUH7GMMbMXQnLfD236Tz2YHXxBwwpZP3Ycd
EveY3lLO0UXa4w7uAYMuH0b1bPAATNGcgnem94bXHvL8WIYzHPAS92mfBlJiK42r
H6W0ttF6XCXtdLvu0+IZGbc5jiqExSd0xt4JRwcmozoy4DNB/F+gpge2ZQCOQ3Dk
ISKWozDbdaA8+qGkYQ/9bFVdclv2/4fyByMBSSoZf7J49rQX8e64/1Td8aJC6SQL
BW8bWtGoJk3OLWZFgqSt4M1qjTu1hh13XGElbje+Klk9Oit1Rvl8rQai/kwZD5Q3
kMmWmWMERQ6B9gaMo9Z4UBM/ZB3LYn6AQpRtbIHIHoMi8gu6IFfxenBfV/FfpT/s
4Q4Diaov9suB4mSL4vLFnAAKrMfhUogqILqIjPeZQ8/GwpaNAWjspgAgYqmLvDMk
N4EiTuSBo35QXyEbCyHzna1HZObSA62yZxw+uGmzc9owdD63weYj7kYbvax9doAp
9rOrA0EFvVHCF4a0gSy6K8Eh5KNYXILBZgAo1obTBuSRgZslWXgs9KV2FZUVNvP/
9bU7ZNBcR5Z6dttUnN3wHJPTWPfl5oX4qcHAbZYAOCab81UdMa5nIPT+NZvhbcWT
kHlQWGM0DLWJXZ0pVQ13mgNmseEthd23DhRl2DgrqtmuggZ1pUU9hEjGUT/iir/x
o0cndlttjKiinPcmmVXFwKd7pKbCmu8WMb41x8m6xVCSf0AiQV0o1SUWVZwq0y9R
3Y4CgLUTCJMBbjPv2D5f7JdDBc5af82x++hHEG0z+hSx5gnAUNoB4Rf56IsLIo7Q
sOHTSlYY8Eaa8Wr/l2wC3uVHqhfguV8ZfSr5lXfB17N20ACaa4CMgBpPFvLMKM9t
4ERy7Kmd4e3lx8nFNJJP6fMla+1fO5QAMdKVBwg4l3uiAsjiGLTPMf6YmV1iyuJM
21zAKcouYLCZNFOMhnpzxvgNoDbe7CsZotUQu9QLVQyPgqz66CtUQU1P7H1KgLYj
LLayRFNvZC/2PGUzMm6geVQeP53b9yY9PJcj4xrMaIFMJoe/HARBrsLt7N86SYnv
XZVRLfjLBzIgWdcdNjfipvcgpNADJItuRqFXiqA0sbiiGV2+Y7ICObPmSUzvgj1X
CBG4KNriwPOXwTGQRu2SHkhfHOgJncUa9c2pKFpZxUovtvTfjQbBrttycIg9feai
CKO4Gv0WrVO/SMONaOBmz3x5fLEhLp1pFeG/6u9jp4ljM4K2zFTERWoN2EwC4+Eh
bobx0LuiPh4PbkU6A+AlnSyqbAkNDu9lEx5c+LRy3Qd6/DnjgC6LbtlKQwoqhdXO
YbZh+YTTUUGZ350BaiqkUjvSCkzm8DY8clwOpo5znrP5SD2Mgq9ceOUKvOd6yChJ
P3HbywV6akp03pm2Uo+5puiRKATYCVJz/4RJuAzDpuES5v/BwrzLSGRVt5UhvCS/
I2BCA6CetUb0Y9FdWdr3UdHVXdNHwn6oJLitODVQEdchFEEy2R9juGmfn7PdH8rd
N7IpOU3bl38XlToOGOTYHqjPlMTr4+FD9Gu8cQ/r8EDFu/G6Q97NxCF6MsaaUIpu
Jp065XdXu976pHiWkS2uQ8FZz3HTuWeRfXY/yE/67yc0Bj8ZQx4xi/NyB4SmQwJ3
C1UA5dkFiuiOedtdpC1ygr/eVRz1Z9SixY9KbBEuzaEe+urYRtTpMjAJgLbmupay
2aIRoF2MWOldBSzXVWWlCXbQ3UchUWwpZjRIxZzQw3d5OqrfldJSyrMHXovAb+aO
qaoDl+T8Uj/NE9aaWEOn4/tcFrVokAHuPkr+4n3FLuzVnV/W6h+KM6exYi3sdgXf
ozgq6l7irXa2Gi19S9jQopqh3SXlzysebDhTD+2WXUzj87hKZCdfsGLvF256pHnV
OldP7hoJU1/ei5dozGjbF4/MZBC8aKLtlLqtFFnS78w32nde2USmeteCAaT54crv
triiNfzFIwNjU9wTRLdF45Xzj1bz05M6mpH8p1mG8ayThaJU5Zg0l3o8w7mAVKmA
VD9jOGzJO3npW7gDuWJwxNK3ol2L09IXkMHkps6ienB/qcmcRg0pnQF8Fk2+pLJl
cR39FkmcWDCcXK4tFdjTCauUmR7t5FkB+4ccKxLim1hFlV3SUdC00+66qV7oayxy
54jiakmW0xhy+yWreBlTE4F6h0xn3iZRgsFHxefPVlbVahMgdHWoADFVcvctEerF
hkW67vSu5O2Vw/2qXIas0WA3Qnp0wQxkjvlU5Q8NjB1NDxXU403Bm3RzugAFbAbu
mKYkGQGT/GjxZL4NrK8lSD2q5FYKw+/2wOjFMeFjf213IW3z7Fhu4f5UF0cIaCnJ
w76BfU+XyXTxD7706gtuSVqd2lZPROKJWjYDJBU/ASGKrJdDebipsA65r+y6IVvf
JZiGF4tx57jmTbzi3GN692Wiqi3Q25Vl+scaqynIcG+3p+DjpJOMcIHHSw3HA61v
cVe7YQonq8hgr9nN7ghyMncMMJ/wLAm7FbNgZRgKIHWedLoeyC9dzxJxOaVaz6PI
sND0C7/A6rwBgQAJK1k2IwtzUeUI7SD3qY8repGaaKM0v1CRqL95M2KwE1Cind3V
yt01kc+YWN7L1sCqrl780jMfeZwXr/UekuAuUn1Ho/sNMrldxpEdsSZ/IHbEupsh
RCIS1B2MNx29pQHGtCOMXuzvjTAaCOJcsh/AKN463Hq2MxVKrhj/tWW6AE8LzY4B
+QtVAt1yi/S0GDu1mH7IhwUZRJU39jUIYvSzZ9eq4/Dm2xT6u44cWuf8gTmLVd9Z
RXf4FvwYLe/QF8tkjmxFjjiQdGsJif+EWCzUZ6E+T1Bbx+8uFGsBw/qPIViNzR3S
8kKLB3DPHSWSgfhyJ1g6EBaSDz4DVLuO2yNJxhgccQjIh7B+H36rz0hmtyE4t/cV
7UqJAIgs9ak4uWGO/szwI9tmPNqIpsN38MMfV95otnskxNuCFMY+YkKHyDhUp/xf
lIzTLKnhOApTjL7QDKB5hNKXN3mGt85AtBEnNELSOjcfLVVQw5YeKtgrbGZNI17R
PIJzP0YaZFje3aUM070Co9MzsnxTymHt0Naz4HNFgxCUIOYc/yeQjcF/65H8Zuxj
PJxm5FraFGDpkyrbbCHIuIwrrQ8YzZzoCWPalA8oFA7sPuLEv2TdLvbIKSKATx1+
O0idOPW3rHvtMmj0pTwzY5NHzubB5SDIzUM1pVAFhILQirEuCCn6hvi7Q0j6SXOz
NGzpSCav3Hf7AeFc62tIv97TxLq3Yk4IS9ln+vvTZsxzdCe3TR2aljH82bGZJYgt
vEmUfKMoKmtLRSM7HEFWtmgD3eYbyDZdGBUxWPpgAg6cSnvfZuCQK3iTl8Z4IKM3
IpXErUg1ow8K6vZ90G2EgXa/A1ddpMSwZ2yy85/frIIdTNh9lp494TASbwiDMknI
UQg/LzwxB+x7FTFeAblAStW/2QSjbztOW53GIFwkYhtf4t3+AzWo4bKS5ibPS00w
kaezctYAqd7kUoVlY+LRNMZWjAQEefa+UnD4LKs6V35zSmtvwdo16jDuH5yNuS4Z
F2dilOQbsZ1/cZ1gCl6gByhcS+tCDzo6GJFIiNHmveFRP6vyRzyU1ibW/b6Afryy
pIZX0m4tJKXWTa0Ep7GhPJNYYuISBH2hKERAWF7ISJxZzSHE9hA6Ll+vQrFE+Gch
7XKF0MQnrUl14/Lya+fbF/YpcXfEFftUh2P4p/VhRPf75JsvPzuaWpp0FKkjuR5q
xHoXlxIWI/QybaBF3CsrJIvkkWQHwcjnuFJqZpW8o14nrpEX6Wf16aq8608R7FU4
qmStqXQQI6cA9CBdHGD1/G5Js191pfWgHPvx+YFSYMo7436aAokK1RskzgLddDKm
Y4UmTrxBS2AkBxWP2/ZZyph03lXuKgEaWyDBmxoth3OtNW+Uy20MtaaT57DMVgYo
lT6ZNiyBABOmWJJQyBGrJC7Lv7lfcqEZ9Plp2w50xY08TsveXLl8T7SfbXjMAdUA
H30h9XV90oGzmojmENW97V3zI1IxsVxSSuG3/GaaLwCunIT/vpp/Khth9WY2bUWb
+LqNPz7qnyPMwLeJyg8ghxqc2UNeeihISwiONQT65Qet9y6GzfLV1pIplgAxngzA
JNBNO7fXYVT2z7Pv9UhADidSMoeOUAp4WtMVMwQhX0loqPZSel6dSh7H2ryBi9uW
dSz5ZYFZ+jC1DP9YCrbNGhE6huBHpVQ25/buyPmUC5HwVu5n4v+pRh3VXEmy50vZ
UvgPXsFiRtlof9iR0D/Ebth7PJG1R+9io11umDbM/AxI4ny9EMilF3UvNH9bORj6
oIHVYdpilsEZUdXf5c7Ng39nfO1zQTeYlGxC2w346HlZUYf/e7FJaPQDqmLI15OH
wLqBkylxNF2TVSKpXlZl95tHH8DqqdVYRsY5qelC8UOrTz0rc9vC5dVGbzfSVttr
TgvbWoBTI0KlA8MAu/4jqEyfRM31xQSfFGMV0M407ThcU6txXvlaeG30Pt0caDBB
wJ6OnthcqwwbTsPy62wFIf2y1Ubte/Kam/+OkF+VLvYtRqkFbkv7s6h6T6w7lAS6
V5p5YEL9mQ+VOrQO4NQTpUdRkcHpxDjy35YwtuzufA6Sx7nwCwpDaLFI1NElaJFb
969+YBKD0O6cU8kw7k2K1o618VanSg6GXTIsM9tGBNvLN3p5j11sGxJhbvbdWzh6
vwXu26rEuY9GdYUzSe/3s0VUK/F4i2CpCfRULj+PvbLOjKxG8qhQ30D/5ThaQKn2
Fz7wtnv6kblr0FP7/BIqL4UAYEGYnfBAnT+x8+Lcm2mWTqeA3A5YhDGOo0uhADvX
S0XS+lvzmgxCrbbS0gC+y4er+vpOWC6fLBamWD56LuAD5IFOgCtNX65FmRj1Al74
7Fjv0OUw2N3GN5ItdLvpd79Z5OkDgXKsu6DPwW6zArJ7Bfyk5cVq2VfC+N3r0C7T
u1PDlpfxc2AiJeRtkJPaK8TaaJcY3VqJKjd0HQa1j/4eL0KqvY2hdGl2iR4Um6wi
P9sgJUjpG5zuUKxgCZx/nbBRdW2JCdhHlA/el44XHAlMf6RkXuJKjLfqlUuYIHlf
eZaMpGTaZFwYHwVcrGwDtj1pACDp5mcZmTtnEC6hjpnjfwXtdm1fAXXPPP9Ply06
tAfeYlS5GoyRVlG+x67CX4rJfuIl12Sz6YmPR/qATgNKMdX8UVCWR91LmygMd1Lj
oWmPdW1T7YoGR1+cS34LyW1+uvClEGVSySc9bnrAVrllvxcRfTHl7Ms5/k/veFV+
7/r9ELbBT54B5ZothMF4fMVhuNGqINcW+V+nXmvoKuESfNzSKsdoPkTxaWUoienA
FH2h22Xp+PC/HdZb3o8RqS4ImSVjT89uvv8gpR2+h1YRpvir8orsnVn8wjpojtFU
cfdqUj7MKL1SsaPUX2YIGa3Wgg9RPy99hypHCxITd8dWpfMyg4/PWQwAibHeS4gP
S4NfyzolGu4vXUWD4vpETxBMK29QQAaFo1z3K5KHlEt1QSxy2Cu8KIgO05QDhoo9
Ww/ZXbDGPvzz2ng3Q+aizioiD8vUAMa7v5CpndX4sHX9s0SzAOsDAJSpWgNUospJ
iuzObS7sceifhd3jsfF585mVpzYM8RFB+WfmZiqL2a1X4J/4CUUeyh29g+N8o5t5
6wJ0NlQpSsiGAASSaaxaq4GUjWE+4jkJ5aBGT4iuzpPxcRu+0AvGbUOvuvWUXtar
O2oub/smQisGvT8+KfQKRQk/HpMQBBPA0JAJDb5njlm8eqqF4eqIX1UG7Vct9bRf
qgPvwuS+N+Y1tuNvqby7eBw5Z6iFqmy0bBZQ5JEUErue5MiguzIMN2yjO0XXKSyE
wuRlCXzNr+ztqi06aHqMt/EM+nIRt537v3tYSf4ii19zBjNTMZgFVBIXpxccon71
QuPxB2106rLh/qihCzp+8zIDAI9cdEwQTkTqvnywKjRa/upCXpcB2ZE+c5R9la1f
/twAuH7pqhEADcHtPeel0aAfVicjGezKqoecngmwNlqxthRiTePvyfLQX1613hF6
gS+FlrXj08cO3dZ+mmvkZ16fWvs33whWjUnxR812TJA1FNFvC4ah4dGzyaDyQEqV
u0ewd6WmKDNgK+mAeLH2XQuXBcuktms+pSIHKrMjArJH3VjOCbwV1YGFCFjzEYV6
Mab0V2OeGZMHrzt77obxuglRnpnKLSbcKSsUU+nqWqVKDAg+5IZdl3QSCO7eikje
VXWUv0L9m20gKGTo8BS2tL9yneh3qHbuy1PE8plIon8vh+tM3HOMsR70dWdQTw9z
o/XXW13RmrHZGlrqrpfAeXDFeBJg4GGtstc9tF0d8VgU6F4fOBR7hfShA3U77hjh
Uk5gZfdjkdiOqgGExBNRWCG5WqwdNr0jpasB8X+489s2KWpD7jjXXnXUqOSGURWw
geaJmzFd7gvq0ZKlIBA5SUfl8tVNqb90ApNFV2xxnOhFdtjclJFhAbQdkVmdJfPu
CR0VtgXS2BIR+/a6yxI+eMdy8SIYLjs8xly0rFylaB2XLlf+N0DA+rkrFrd0sZVQ
f6rUJGkygVJ/wJ9Wfri/+KBvLGoMfXPkRkwe573bwyvUVJ5k9crncBw/3ew/z2Gg
6B57rv1WlZxzb9g7jta5qZW4xI0XuI1fCwQ4uwe0Qfge+btmkRPGl8ihmXoe8KLn
A5xyx0tz0fPmSXcdDpux+An1Lf+sXch44F6Gc5mHw34HBPAdnDZaJxvNwIMNROZ6
2BLvwNDDoCuCG9b/08UdCjJmJcD4ZRPkufwE8zFSsb1T/nTUAM8HF/TuaYs86ITb
uTTHjBnOQu2gdtTaCbUCg9Fd+2FQ7Ff3vxC88X52NulwSiJa0Y46ZN77OkVq3krx
Qv4rHgMUCkLICadOsaFXsuOgVMdeToFF6H9EIl6BKy6n61BirGW4cfDSqkBVKqqH
e2qgw1mzCusZkh8TzeStAvUt1lhxULTb/GohBuY88W9rTtHZ4DFlV2SEhOIB85hR
jgMreQDhbNQ169ZQzu0Et4+u2kELVCY5UyLsHmFn7BDl83PoAvF8W0GM0rA3Ee60
QGVF6+09RUO/WaAkTaYNXPj2Y0Hxiolw/iRK4aU2/vgVBaikse3KyW0NeQrtfarl
WFp7h5n+i9mZohsTXhlzEQnI2WWbIh/UIlULBi40M/hp22Of/rSBo2u3RTAZHT0H
GmhcRhi8YWFh8PDyDHffnhd5kHfTn+W1r3v8rKeoVO8zDCSYosdoWOY+EdzuYR03
8EWQEOBnEnzyZPJ2+9ShG8hkA28tgIuoIombH3EGRxVeJPLt4xnqJsoSHwezIlQD
MVtiTizEf+BxnKJqD8KBsHBS9S98dFNtmAiHFRnDU2Hb9kfSWMxX8ReuwD/HNIuP
4E4k1yvMxV5kiKeg9V3Px6+n6KptLb1a35AXwVUMo21i8jkeSU1XbKRtDrhzDeB+
e91HIsmw7KEGY1KWmHPJQQNdGLggFWOYIS9hw66r9vQGizWymPqCJEEprioY+I9U
YOaN9XSaYzNqhEgogu6iEV+UyYSGdmI/WjdRxARB3EetHSN8NeID+R9k2qSg2KUp
g4awt2TA2E7mphQjhvpyrFvMMUfmsSiyTDk/yDKsBlcv6xy2GMu72e/QkaiTtfTf
QCuhL1hv8UiFFbZo2aXbX9wQoW2H8MWHxkkyBbIgGnflaDMZG/L7bcVS8sGZBWjP
5sP/wmF8PAS1wCGhiGTVypzIKsHutRS3t7c8u5i6NXyg2DxYbsYrxkRICoqypYdQ
M7TNQ/EjyamKwtouXffRWOW2qjU/6JHmgdkWPSZiLMFioBc/oq3JHYHB1ymmV5w4
RaHYghpk3m9bV8dZPDE1NPeY5SukBZNcYwnJ+By07rm5zX9TLBxzXQWgwMGcHJTJ
MJAOhUgYOjgo3RHSBva7XTUZg7IojkRCcgdRqrP54wnxF0z0wYdWoZz14fE12d3T
N62WU495+swJ+19ykm7sMMPLQLH+JGCnlkEKnTrl11m2X4A/Iex7JO/PaSrNerkY
aLkUdO50UD6CMVnzjcuvWDVhlDL+rG3EM6W9kCxB09TRwUPLrdYN1p72exlJc+aG
qYfnLli9gpP6M45fLzznR9ayL0yNO5uyry9amMJfb0Fywk9+9MrbL8Cdv+GTv+dE
3uHjsH7qfVghk9/lBRdix1SpuJAKHGOBRfrXwZi/Xnek3diV4pdn8LoH8jGZ0Uuj
RzHqwQjvgAo0oaMtsRlvT+w7uEQFuhCBVvIx+HEDCpccJmXS/aQbNZqdHNGNDLxF
arBjOnIFqIRzulPImXAiIHD2/LY0aqLJscp+bgixLPlu4xWt5F8Fj0ozFLk+v6lv
2wj/BLYVkTgcMvnQfHzIUyKJGj2FOQhPrnqR1Q/98ejqioXkhVWWD/BAXqflr88U
SNHv28VZWDO7214Mrfwg8qY16Aw27GQY7if6iU6hEddBUwqGA61TF3wysca5Jf0s
pY4EJnKXvcjusTcRK3YUV6e+WCD7hHRwj4aTbzLpFiyVcHZI8MELb0CRnvDWd611
1EPb6nOSMiiBunWHC+z2GNaSHxuau1U0DUjLfjrBgrev1R+Rs/XkZ2aoQ/90nSJK
vn+PK4236wC9WjlhrvWa73JfVmndOkTZ/j6QGeq5OhcCWvEo1b7coqGo4OfA2st8
b2bJmcHXxfwSqVcSM41w3Tu6iDMD1vByVSduI+cdqTSDk4nUMj5igOCUwi7oN6EZ
29uoGKAtIcrfybOSyNzV6g7DwD3hqSI2n8+C0tItMA0gUguzcXWMeT8vvnC8Orl9
X3Y5/BwEsa2sZt54R6gUk3M+3y1qn3+2C1Vh7qdUnnYPQHci2qjOy7H9z5UUoRkY
mo90Bh2BuENI9PNkEEwFzUh13334+A8ZmI7kbWxivKSRVHK67mgArP+3emxQNR4j
LPsQNL4iDNEU/E0u9kCBqKfcN7FsCXj4LzjMmvSMAoYKebThCrwOVw6YPOjCxqjD
hrpgMf3K49ICnEP0Ab044m52Y5UP6cd7ARnBY5XE8pRUojDwcHKC94G90lHIyTYC
BqCRs06E9V2mB4lTQHJvnUto5WXp/BSwRfkJxQSgzYagKGJbL2eC4ay65JXWrYKv
T9esUxDB6LbQLigbwI0di31xGfkI14RdGWbV4wYwIYxjeYfHgkvxcF5q9m6q0lcn
tXPrxWQQfScAyAy6SR8km9eR6GGD+3swJ5fKB+OE8l7Unhht8bpxoistlL7wNHux
oend3UeVGG6dn2ZFHMzlj/UJDMWvwQQ63S9z/DqHzjzpe4t1qpfWpSTHq80killF
8BlO4g4AYEhuwgyUrOw9xYFziyNj8Kdr/o7DGiHnQu8KskMwwu/4mqzyYucFBF5s
MTSEMtopl3LvQ4FISY2ArND1+hFmjwS9X/t/yRielaIjCWW89TcvkuC2UiE2A/hY
t2q2hYZWHVFCz4qIhbMMwLyhktOhNz9ZjQ5Vs2yYUVtPZ+yNlWmvpZHy5NXIrlus
s3iQ/bhWeXxUAkIvvs1DF57yyA7wmSqB6gkwkkLwveOmFXyUFAwmkIcTuK2oSoR5
Xiupy7xjnYGQwIxnDYtg8sus/UrckY1PzfCk1FqtjI9O4kUBNXPBnZCg3FtTm1eY
72kQ5slre0TIaa1Iz1yDkvZalnsyyvur4MGc1U9CX9l07yk8npGMsWIxrddCzuUH
NA9Ij0XCp2JsSyZHmFvKhf3i8jARdC82FiDckzLx4MOkfXjLGG1KbJySQGYmXofs
fQuBSL524qEtwStD98+8XPZvvcBGf+NWcjXM1Vd/Jv1zLaM8hPQH+PLFi6V+pnRM
Z4tXbY/N/KzAIUZ0UQYxakR3nSpV/PgDjRu51d7kaiAseOWB23keBIEwRHIn08ri
u0j197tlYhOtT8dnUhFmC9qV1Q8xrpEwGIJ+SAph1jCHaoprfTH2s9q7Y6JCQs9f
bL7mUXH8ocLWryqKy5+THwYAj9iYWEwG9cr4GgZCeBfrzcbcTSh0F1rD4bhi8nUk
RVCADz2cPnmgI02nfQ2p1ZUBZ44yPp3qcW1TRjInRePRC3lI/UXg5rnbHV+wtN11
90uBl/KVnzlTIxjmdCbq3ZdHg5Cc+wNSw+4ZK1tUJOASZXWVzRL/bqOU89GKivx9
OJ1oc9gE0kVKYeFT37I6yriXro+bZAC4JZK/bPeVmZXqaQXFlYBiZw9Fu3GN4SPk
YZlFvGvHKFa6SzZKXQsjcP59RKrd6bGPOEbMyXPQHn6yxnV6xodgdZBb8o6nm8W2
oSKv7uyMJCqdb7qeX3/Y3S9esEwyqf1hgm0UbQXeZYMwXeHcJuJcjgjaaAPZv3/t
/MAiLxqsA7GK6GG+N1yqQkCXz7cMahj6OUbTtrUVYQjSbytWxkoHgR2kqUtNfTaJ
Hb0Jdjv8lihZzTJNiKitMxnRwjfEMJld1BteMlPWsR7MNo8h3xb+6XrJKT7aStEB
aEWqNMzef70+VLT49pdJXGQhBViDJA6cuXENogrFbhMRBr6ySdU/7o4Y3ob2e0Xe
7vd+eqz6M7ObJ7jUZDTG+9fOHImx37Jm120gzkI0WG0VHQsJ8JMaTFqV4S9A21vt
3OXQVtmiziLFZi+RcSkeGRTuUoITw0Xe50Lxv/TPAgmg5kltlAx/7ztV3p6jJ8TV
Ti6K/0g97wq9xTGg9Vq5tYHI/jj+EVLkzMAhgX0mBkaLsXisnUdC80MatFz7HAc7
2RXgVWzgVjRymVe4KfBkXpXKSxyCNYOphPMRPJPCcBWnKPR6sP1l47eVQApXdUsX
7OvcYJlxbNViRex7HXNl8eyAUMiXHN2+Ol7DFJpbdCbGBzxp3w0DkVbxVGXb4q43
m78Xy/it5RgyTRYpxT5/D33B+KbkQXHTWaRDpifZOQCwO48UsxyfznUMtY9WDs+y
tYhq3rUx5c2GNECBHTQqsD6I8ZMX0Knc40+XK3uff2Cw6w+yEjLsdM2Fy5CEbMTb
5l2JOeEJ9iURYV0VUc7Y1X6tH+rDWyl5medWeIWjdLDn/T8xezDRT5zZCHg6HtIN
/NvMbVWCYs4+nO2/DSZTXUk6/KCZMbQkoQ1TWQoTWNQDAY7zNGVBySg3effubhYr
oYI1IS0Q2nIeyrffzr0HrMax/YOtTbw8ac6SE31jerpZolQFEfzktyWcQKT1RPbw
n1aeErmaJ9klQQgywdnTYUPVuVs9PT2WwKr2OO/4YGIpW4jR13slWEjHU8h+cprb
GjTrFQQTkU5yss45PATRUTcj29e/XtxRGvBBubkaiHtwMMap3BJcNXSkMpSGpk1X
p+qjXHryslzdf3tjmyr+Qmv8AjbPSXXbJS8Kamaio+6FEey6aaplHVdSbpaeaqq1
yNYoTzub9L+s/V1l9Xfx+sL0gOZhjOnmh6dNdpd3WvNQiUDiUVEhpa//KZ+ZtuzP
HpAPhb5OQ8GjUADNxYiG0x3Ztu6UuD17GCSwVr0xpPF81kyBTiDKoV0XFtQhZtu0
/wYTXHHLZ3iTGGruZ75bsGru2p1IEPrWJQQMiPSVYB2hr9WvCYhjYwGhQBabAlpF
p/hzh9kTAHOYcREJp4iXXAjjavYnnmiJzHK8fN0NjyAR4PLwrebH+UBLJv9zsBR8
me6E47KbLeGzEcNaJui7IhxNuUoMIbe6tyDv/cQeVBGGJaVt+g11m6X6NTHJ7mDP
z99vRCefNk7mHkCZO2/DRYVNn+hYBfE73QagGxK+nN0rBIWW6LHjQox67RkD0eb/
mZPwKTE1Uua/StqyOVzOBhChJhksI7c4r6mRH4SicCXJwtzpGNymUsb99IHY0MGf
+zHQnWYfTwQNTsKlue+UjbKXTzXdBh6sj2pRDfQ2Tyujw+u+9Z6Ab5NUURjTq2Pn
Na4yk32Z2jDhpIJe7PHLaMAg+HkxJk4TG5YRS1GXMHXQDC0IWkELW/eky+YOxZih
dfiv/3+AHJoyMBOzbrzU6fzFel83P1Vr1GF9qp9+lV56z4uvZ5ESZ9+x/QNGTzoU
I4mubEINyDnVh4/nt3U3E8cVDpb0VA55gV1AebWLLt1q069a4pNOVIraZ9fz6ZJ+
kZZMFw0frAS+JInCA9hLJoNK5/UF4QopxabNFgPPCo5YB6dGpu0Xj8q5Pb2c1c6Q
Ja81z57fjmm5nwz4DuNgnGHVweJnh7mT96W3H1Wv9sCcBO7jL581yrPjRIaIzL7l
eBlQrxwe6Ben9LadVu1l4WOGHAZ+frPSVQrItJnJNGZhncbugOWG94VBhepvBiSU
2TsBroe6DKdhZj6T2tS28RHNMnq+IFpqnCNcHhOtzRFaYrU/bDzaVpwJekF9N5sP
So5JbYas7A4tPQbu8qkwKu7ur/94hrcmFUGERxvY3R3ep9DQYPXGTHNUK0V+hwcT
HnunBjjbtGWFKjQZEADmon4CfVJ2cqE9FBeZEWv9YqtqQOCt6BevQJv+P9nbfItj
VIK4CNuaAbhcRnQWfxKpaD0lihIPopGZvQLJxNkBrjXTt55CXjS7MLwhF0BYF0la
U0OwVkEVGwlaw9dNlTVx8G5VIBCpOG73Gw7N8HsvguYSSoDNtc7MyJ5o3Z8azb66
U489qYucSbbN23cT2bUUMShVow/GecRdx7doV0AUfnJNa2dyguFs/da7bmAyO+Zg
F9mdsacHRPJDN8igkg+9yVVKfOZ9XAGx7uLF0QPdLS7ONT+lDqWKXHgfMjClYh3y
qNLx9WAs29A/pRbJHQ4ufM95n0yzVu6eafsL4hIYehYk+gffA71FiSrM17T3zMzw
JnpESoxaQyC+smamdA9thbVj58GVVqks0wgUxMUXXDfLJ/LC3v3oUjSR+/bIKM8Q
gKg4Y6xmP1V2da01+z4/s0phE8XqIQYKDWigvQROpbaUYX4oE9LAI5N7/9qUpDTQ
0YA2LR7DFhXHwTWsu47y8kpYlZpFFTcB6JyFHavxHpx2hPFYBeUc4GXmEqx9RCmJ
tgxcdqWtpWNhrDpLxGVy5SSzw2Co21iMbj9zjlpYxyq2fLZtXHjnJaaspYpRTkyx
esVWERnvBDiPPT6D72qVWpYGA93635yv8BzaUqO3R57h2meQHI1iFuP/D/H2Hgcj
MXkaGYkb0XQtRL3XygKxHii2jYGBv8Pu4CBhxNIaB9YEiCSBq8xtcDBWkB+7gyye
wS8o64jb/GZBQoROdvWWbUz732A7xvzd0fdZmjBkZetsyY03/TIWT8YROk7YyOJb
tdN+OckHLykJBaU/gaa6V+XIXs8KdIs0rRk+95pUATI5gUuLROl87zJEFTONVsh5
rgpLqfmSq4xeFtZlpq+OlZg7r+VdeWH5FwOUYC2VsnvQtolJBpMngiMhI/936Yhi
QiNQ3/hR9DVEM4VMlhow2dH4SN7waFcVKU2ykqSfjAnndfcp4TkxLPvkaLxOJck7
LbrRagcmmBOfbTf1LoROqVrsq2GKJ7XJfKs7MT3dFzI04llqCOx2ZUHDIkiD/TYl
KDgyvPid1+UEQhN1Pk4dSOUUWZE/Frjs//tWKByX7moWjfvif44DzJN6UZWaJGQ2
IexaX+ZtxiKC5qS3w6u9A6EmkedwlGfd9IBeY/f2gkVOalPwMCMnDyK0ngoO1d7H
t8zwsNG0BSCNgITL1V3ob0c5yF0QhDtsK3s+YyUbkT8LneTzsEijcqczqklvhKW5
/y5sEtovogHLEPtXLPROLu4aFGkEq+1ZPqtqlBMHQIjMGo5ldH+/YtUBs1Nx9xMX
J8rxWdKueGMEfEkSVgJ98yCAHM2RKeCo2qPLSPxcylvOaduHWjclDhdJBPYwHoB7
a7x6mmona9bff6ZW8rCFWJjc3xBcMBlfbHrRazI1l5S9ejWjLNL16UZl3o+rvU5U
/bDqi70/V+hHaslA+LW3yajB/WPZXBg8rjk9theDzywxSgTT7qk4L6LkN8OsMMaE
I/IEzKTM65r+mtziZneHOlYdzaM3wG7Cxet7lWHuE0vtlpeoaBr6yB8XuhTQArI1
WZ5qMidkHmPHo90ST1k7CIfly+nPqiZkSft2iW/DylMpCQeVZgLuQ4T1QJuZCxAV
kBC8pUYSu+dpcO354JDif7wdC9S3hCTB5q5qBxJkjZw5C+b6M+DTYZh/IcFJQ907
uW7uBHlR9zHgEIx7Z8srOEoGBMxiVfOmcsBYosAyya1Hckm/shLWqZUuRtj/t6Jr
lDJPTtAXJa+sDPs5jDmB4IoKS0Zlx3pdyNodAbrZAku08qkZ+scAp3j+9JMuYJxZ
AD7PKMPJtPjSYrErGXWdPI3XA+MI48TxQlNdb5Zs7D/UZMcWbUXZg/VZNI4fy8te
fTm72EeWy0WlWW8or3fyMAc7OvAlaIN23ULdbCRc+fH3+BXxaensk29/QQbVUcDA
7nKtPcOzgIFaJcv6cI4KRj3TG12Oe3zZWmTBSAbhO8ouzgtRlPe8s0PxQ+6kYwvq
8ecnxKRynR05U85frwr3uFS2baOwYMPbsFCYh7GPmCQn5Usk8eotKJ10qXiXufvd
kNzPe6DSVo1VBJXMpNjT3UuQsNPDA3jqOOGnnIRtP3+qNQx0Epkq8ndDR4aDBQyo
Q2ubA1JhQ0O3wxHMfBa2ripQDxWD8/8GeeobdEZjFmafl7adJ/hn6o6toApcnHLZ
8mgLa/k7Yc1MIdMY9SElyknZzCN60vYXGtTSLxAeup7x7/MXv92lglZYkbRfV8O0
oTZvHGKFFutjmi5rletjagHhNfsKdWUVNce3u2KjVHKGmUZS6tTNpeKbFUgb0rLV
NGfDVn40fluKJbIg3PobTmaI2o0kq4i1ZKt51pACQLN7kWLlD+0mrebdll3vHS7q
wHnlsPz7b3/b9qlLNwvoaq3vzrYg1If8U6qOHuYRcyiwB9uRuH6p/D2G/LhfP+Rc
aZOBrKTL42ex1VMrgePXs3xKjup4xuM+iIOvQrV1sZSc0uOF196SC5DjkWJwthyI
frTxfVGtWwfde2ddfVZ4MWYXKS2lQdr9PNloRS3BbZr7QMjxIFf25+YMkXk8J91f
kiwbg21M69qb9c8nQiqzUlm24WYVh/qThz7N2AYyYhXAlPqfXMMkTDrS8MWT3ePc
JmwUh010iuU5D882QZk8JOfBuFuCxDHLcFZUlrOcyDnGyb8FecvryvmVXuSu1U+R
6xMh0z59Pgh+q7HDm81lkTUm/RV87RzCvQd61L33NRGzd20ErAGwhKmTlF9C6gDy
YoqdcMDFmQ7/YN7j/HStoRtB17WvDzJkF/DCQhiiPqnVCnvJxrJx5VmyomvGw/2K
gxNLNM80cbRGuUv7RHFpXldkjQyI5mayHm2Jnk16BsOosgIQJlmen1WL3d2Q5TWi
u83ytL1mR4r82Qpt12z2aC3KXplKkpx63Bp1x0WwnsY00zjsJmY6r9pdiJM2Y7G+
L54gM/qlsBlZcDnLCG47uBU6dIMFry7uW/TTdYe9bVRzEEnTpWlsHew+qfu3Cb8/
oObrJVwr1RyQaRgVhtZo9CDhXRP9v9I63PXUvILlW598sYsdSPwyNyHBISngZGmg
cqNbYFZQ7bG6NxbF2i3GaY6R88cm0U5R9emYStkO1Buxnnikyoo5hBpNydRx7i6R
5xa4W1oi2h0zLkMT+mHU2TMKQIYQFFCos3bIiF0fY1uPcYt3O5VJZJgOApkRVYgU
pOEHgw/XpzsHh+6j9CC1CyULk5i/kzDmG9pDtH+dZ8pqXlE/FPG5Cte0F6yTXmuO
XHGZvW/HVDZ+XD2kUoB14quqPYRpoD9ii3Wqjh4iATRtmyPJcJhLr2czUFqIDzws
ASr3Kc81RlbcnbYaQDEwmEZ4j54lVjbqPwjteVbGZlDMywNIa2tGLjgfFAZB8NbP
SLeGi0OZrYZ0lb+WFitOViJMmPsQ6ComGy7fQdJMbaK+LuAtAwKReFIalyeqdtyH
f786ACr6+uXxaHY++XR+bsW+Je173ECoz3U5l4TtPV0+pu7oOZiqEijgYX5FRTd7
9T733FIiqOJ/asC30OBh4diw4U81i39jwaqUy185lbWJsZ4wgDLErdVsCeG1mwTG
7HXkQ6XbaZfPrYV8rhzDaruiZc/4OHyVR3C3G1As3a1kmxb1EggKVpPpLlGciRjN
A75YrToeHRsrarBgP4Uh+VZk5QqNMHf4c/6s2q5LfNgH7Epob3WlbCERzsnuJAAy
T+jjMphVm9GpUQErzbu/5/SE6c8w9acqWfSNOA02H3dTxKH6UkCd741c04E1ynUB
lH2xyJW7m0txX4wxlEmOJQP047IJNF0tw6Yt1w78JMzq4/Iycjv1j3sOh8w0Hk5f
b09yr+x44z2c/23lCbQ3Il5SknseLCpf0E87aHnCNbawQgK4cNNV5BbXtKm1mzkx
MbC7uzv9HHdlwcSfefLiZ7K+q0gzFaiUoBAyjIF+GgX4gewQ16iPfU9OfqR5fikF
e9FjdTpbL9O+xmiLmQcN+RC2IMo/8j2p18s5VnA+rTmsax8v4UORWaEMD1KS3Yh0
nbXwZQJhxrosVCwVJfE4it/WUWdsYiyEmzSw8Bkv/cuuw5kYJAJHw50gsEwmB3Ca
tajFIuhck6i9zVzwOUYQFtryJEaqguVk8onZpj6FrDk9WiZy7RQR+XcZZTXYIZZW
T2HoxgRkDBfciDCorq7XBsZYumwasiqOeUo7KujMeJy9nV9eMUK4bNu+ZVjP5CFp
AWEw+S8yZpLFJ3vqxsuttnqItrecOXfFupJpsPYUxOOEaQQQHsojMi0/rsnH60Z0
D2o3muO60PFkI7jrnhtbYiQlWi3efFNgZmdMrQJQKu5IHjxCpdjzMtKm9k4RlsqP
bNQjOCG4uCOqTx9b++vchHJq+adaTVnZGogHfleCE5jkRCo2QZ+DQAAbKfokd7h1
eiRH+PzVqyjEP2+41d++muIeiphmZ+3TB426j9GCory+d8DDYFgnzIeBmf4TDm6w
hX9X+AoUg5+zXGb6NqTQ0ryAtw8kNzbwkSfd/G5k0ql3IVjO6gL50JgitJXNpfkm
r9H+QhQ8tt09ACBd5Cl61etIBsoOl6GF5UcPSitoYHEU/+0Zhk6WGNI3Ts5Bh3Az
IrHcwo9AOlvs0x/IIAZWFe9YbWEXTbn1Tku/6o408TKB2PMPlEJlyz+ona270zJO
jk4LunccnLqPxY2mttSpLSulFuAYfsrHthpns9x9nAGmW5rV0S2ks7l0h75q7amV
XCyDDRNTpHoZRdf+e97xCuAsSaZF6e1M1Z6CAgI+MHH5gdFSrKaWpjfWCRBJ7uR1
/YjymJC1DjJ5fIVqXcartGAmgQ2MS67AKOKBtujuZIfNlOPVWu3/NNxd8IsxJUSm
N/HFSG+tmHcCC9KutrCe2Ion5zogITGBbA0BSIwm2tSsNFdphbf2DgUlYmDhw60y
bMU3OSrHSdTjR5Zh+roraA1EK4LJ+xHN98/YkBOroj5k7T7tQY83ZE6LNkWpflRz
gUv3aNfBvyZIAZxQYiivo5cbrQ2AhP680oJ1NiGepChi6boPQw0MgQLJ42C5Brzi
AqcDdSvC6jwfgGGItwUjo9CNeVwIjniQCH3j/fmHzzhMnmpALA4/HN5zQiWW7KXA
peGfP2w2mUVSHNDS71JyzInpyq0upvfqOz2RN7lvZDP4ckuOSvgTI1ntUQUWtJTY
ZVvs0hl2RAF7nRlO6OxaXg1g1hzBb02dordkK9A5dmLdZvtgsa+ZCl6isQoppW0u
JPsbeUE86ciRuPK1hDV7WdqDIaRqMbqZc9UDhLxwleGdIy/3RNbXCF7xw4ZJ6vRF
yHaloARW+6E3cgS9NHq4wNY39xakKQN8rgk//LzK2P8+DPPYeUDlxYoDd+lgTMl+
7gPTS1uL3QSM6BdPtEcu7oIQZEf9l1YiapdRuLZlPh0WCB6Pxvxu1+I2gIVWBKaJ
zhYnM4IIms0dke3G2MaGvk6ak63N9P0puOZRhShHQsydTXUK/+ZJ/XtbUBwEom3W
TXEopkxMlwpvW+MWtqD9SwImpgRkUS4t2oFW1MnUTvDDTZYqFvIFlV1V55Zze/BM
V67FHqoH8hMeDfMA2yFalBHo/J+oGx1WulEb/biSwEGEBhkTO2isDTVP09jYQuPy
NYPiCxf4MUG98/cEwwg4nAVf5ie9bbwoYj8JCYZdkEIAXUlz+PGXLjfhBnGcqU05
pmmcqZnFkIYBxFcBV7L01UejFDgmuXItiPGQcvk+LZLHahwmcyHZKPXny0OD5kLG
fqfTcnmBrCixENaP1gSLzFj0la0+a9Sjz5PB1gaUiAq7ABuOQFn64YY7S8Ve1opz
h2iMAHEAHJEYMFQhkvSS0swL5CRswz3sGT4iW35e3H8VF7fqeQOCZqbLbIdAmD09
yNWB3TAfHqzRljUqxVP/cBONFsFBzhu0paBG+3MOBurj+xXF4dxQQXwXMJmg1bha
UQbg63S/AtjytCM5eacyt4fBRTmkgXqm+7qjZkJcEWGKTNNpvobcJBJ9XHxJmOxD
VdEdYWgl/SM3gFagf42Ug59PYfvf5r5tPibSSnE/kWLbdyA/4Rdb5C2psMQ4xJkV
F6Jbdu19wGYT8RfciN6qAVxBNk4eb9KFQwrhctiStFdksk0DAyR519Io/RsJPm+/
Ey27ZudRJ/xJmJNpMPAyN7HE988k6sTmijm0vJY5mmKjVwznLUlmQVpPyqHuckf8
lW238XvaOOZtF413YiqpCWf/Mt3UBrTWVfuRyIrKjxC5wXNFCbYomH4GaPK6Wmce
vAc5xPLJosFRPdHbisvD00YvI4uOUbXAqSfloTEZG+UmE69hSd2IXKzhPJpQJi3p
XM1tq3e0PnH/l2nMqWkSze9qW6KHwlLP8Zas4JObz8Dk1iqDhLDeXNraROBb3jy2
I3fwR27jfyOvw1s2AW4iTET5km78nGT98LvcLKJ1nEW00HibDnzJyLAbEB+wYQdh
+oezMC6bJzv4xE5xxs5QebVRUDenOISroqitAKnKBF0HVLYavmH9Ix8TUZx3a4ZM
nb1k/kq5/54vEA6TuJ2aK+Pm6eO9fO4mh/Hbln0PGO+nR5V03TNLetTXGHtR2Q1H
Yp1Rduc04KEMSna8hm/+91+bH6y6AQY6RMngnnKyqYU0EaZjIRUJhS/VqyymGHWU
bME6TfkC9AYO4duo608nALswylqtJiBouOZSm4bLcRSv18wizjRxxobcgmJ+ct6U
vJ2RlOjVDIB+KX7j/9kk6E6k+EsnH54bqzneGdAwCsIrqC2y06LWzlVEuz2Vv3tD
ydGHEK9r7M8rSFQl5j8Xah0genMd6GnEbkse+sy3QXvBsahjkeXSxTgNAnti4h2i
SMi3BZviVcSMhIqxTqKRA191Fkbn46156wSylhtjJrbw+0icJS5vkGtRHy4bIS07
nVYC67WhPbaCJJBREY0icMHX4vRbiT35V+j0wrTXec3WsF1AunwgX/gg4uIsZnTt
/IYBKfwecdOP+Zl64BTpVhSDGbPj7m1+OTYko3jN3Dkv2XbH7K4e8voDR8Y1qcV9
PTa5WvoTbztfizO2xh8QTs5rHfGnI4/yCt2be2inVYj6excpsgJuq/T4Q+XVx7Xx
Ew2sWwRkHX6KyloBDwd5OCcm+7e16TGUa6zXMi77o4M95oFH/SmKjX3GMapmoFo4
q6T9vKp0YsKkadcgSpKgq5ZCi/3Zu9455wIO9Wkq/0PZvI4JArV9PEzjFIq1Xno5
cJZAy4dR1i8Upb4uwLIZerfLdtgxVlqHCs+RPKB3PvwY9OyuWSBxni2mB6iBSN0u
uKXMgl3hp1g2ocyPrJ8eWzFefgXModvVP8n0sX/LAJdSF55qL4ZHhT7jorlsMAuV
jyDoW1rW6YuWdyUn1bbGTMePXccfIbSFaOlrckNLQ7QbpYf7IMZ6sQcWx1MTtDqy
rzsMqQ8w1PfAfDJ4aZPCuDTnurrKVomOXtTXuIURTN0Fu43yFCHR8yJFlfnmlsz2
NM0mr20zXRfAp1Hy9ef8Y+xFrx35/MoyfrmENCpVQ7+zbO6atOLWVcKTDxeCWPMq
ErunXcSz9a7v54IqbCnX7Agb6BruzJIa4wc9Qh+mqzIS8AYT+YO0397aikOL83Ql
BLVB6o97cibptrrsO7Nur9L5YREHIrDzQWlqL9bEiuSqQ4SaCeNb62Wt3CkYUzXV
Mn6OR2KtrAUqdiIfzWhAqu30qflGVElEUspiFW1PM7o8FHeKPWeNWAYcsrBRmj3g
MVIeCIZGp9WULbTiRTyUYs+RmdOePrT4bserKHIE2/2Rh1+//qc11zexx/gwCjh/
Srra62sOWqI9EKhSrw5OE7BuH5HP1PE2qarZtO6y885IHJ9ekcLkDyOgw1MgoKsU
be518m1n0whi45qoVkM5o1nM/0BevHimHQKNToa2djEn+tBASD2Qo671vcBfhfKN
j0jcajC5dDfZRAN7IU+KnGhLKgcxPXo4JoxWurLpn86cbylLl2IIEy4iNguU9aLr
df7K1VlNTuI79OhLQD5lpYgSEbEOoE4O/ipPiZMLb00BOeXR/THvl2Gzh2gJjxJi
q5fZO+6o1TuXYBtb/y12xWw1O8eEYEgtUDNGRslfuR6Wo/SD1oh651LFsikvCUhj
GJmf06suQKsIeD9Y9/wd5az7xkf5aUckbbVNYo5YyLIfIXKn9P6k/BgVYDm2C+3L
kdHCaqFxWv7NpO8pU/9hFsb1QE4DFZB/eze1nzTNbR7I/o3ahVjqZJhukmIF2LGZ
scYurvOQ2RhqzBLALsHgt/AWy4moA1fbqZbzwT4gGyHYhbt7j9W8yeFSdUpqUplc
uiKdrJlyJRHg04b1iY+CU1czA2gZCjHzfmWgDIsQannVy+KWwWOw4G2AeoO5ke4o
3Bfna//6VckjIs9VoEPl5LPmJeSn4/49j1DbUrDJzoXfOUdOQHU+/TCDsJZDUH8j
3FdRPZlmrdd+/5vqxrwtZxw863eOh/PffjJmo6SpMzdygGHQlmc+e1QUP2n7W9r6
GAVpcI1o2pvH8/jauhLyaJ9GynCY/LtZRRZns+H0XOLoC9CGiA6VrpuCkqHH/UQn
fEqOK50zqe20vKEHazcMDOuRx8ERgHoWGyrYyW83o3J2HQvShlAXpmg8VCY4Giwx
28OPnk/Z/E/5Scjks5ocXNHHr82Gqkkj13m01PDrXo5CEA+G6O8ZpxU9vz3dypWM
0UJVvffDq3zGrs9Aqy6YjqG717HhLzdVJ5jhqeVDNYvcZGtZbdlfXzCV6WQhgGIk
05DWh8vP2S71mOZj8D6vxTP+kwW39xTjZolipRsOk5LjsTiPdQBjpJynVA4B5fcg
CdV1A9zGZeutzb9KPOLLWuCtBDGMN1E20TmqQvm1MjavqC33J9rzrVS9WaO8AXPG
0i8cuOlreyCsI6wEFARudf6SUjoLLS6bAF9dizQaudZpxzxMJIRgq7/tXgdeQ8jI
tTI+oDR0KG4mQqEBUSfxy1VyVi/CzFK8UkTmWh21YZXoUaapoz/vQFED37ZWJXLX
k+x3ioN9FGdbekGrde5+7US0xHRxke8YB0voaBB4QHPjdcUPUhPWyub5fzScrM1x
4aLRQ2UY8qDrJXSrA6LnZouF93KIFLrKA0nxmFIbQSwLcTaZEVhGpWlx8St2L5BQ
OR0uUVPljUDtiXjdwN2PdKYs7WBgYrYPFeEiaoVph9KhcrrWMdrREIIWE/aFcpPQ
P83EBJJOCkuWNn2LF8aXsn8e3kSjbRKVuiZZ+81dLoGKFcuQ82e7seEcxv7t2vx0
RI9liSjVVes4aRE7LkJFNXUCExBb1he+E6p73ROGD96/kRMJ/iGDYPZrI/hi74FO
VfspdaCqdLeHvSSU7lBHAVH/OG8eF9sj/XAAdWH70zt1/ekfehX+Kxzdl3NmZMWJ
PtDPF4lXlL5G1DKxYibW+GMfXazyfm1zIeU1cNNpMTF8ebHi52XHVSyNZ1DTlpOY
q6hnowAFZXbVhRe5WL+IQAkvGa/qSwWuCcB6E9k8OfLXq/j8Bvo2GPyPvNar1uHI
/kGhZMeJF8AIcbuc6kr4hpD0z7OYvZOIVAYP849MF4TPLqMKrvhhMZnVCcmGkSl1
dzbZlPAvEfEWZem2xhtcMfD68QbertByPAHhhELnImJsJSgHK7Wjoja3ILHWI2SV
HA6u/dZ+ThikujsUpnpr658Q1r3i92aJTNYFX1Do40EZ1E6GrxqKLRb8DFSFAhy5
gkwwdJgNMQ1RJEX94oZHT5Ozh0fwCsxUUzV/YC0NXumF22VnQFxyUCMp3BTbnPnN
xN+2GOVGYjalowK4rokIWhAO44HXNRr7XwLEkjuDSKiFD2LKpRRp6UL+LHmLfbOO
j4nV86DKO1V4KNPtFmjs8crFAuHbueDHYx7S3p98vDupbwrfgauAeDQzyhRlGE69
J5KLLoJbOMm3hdc8buKi7L86FbF41XE4sgzxQ6zkjpP+OoaujY9eea5Nyk1G9RGq
DjXAHYaMU9H0s9zE1lWnUtlyE3FSRcRGARw9DqDoLkC8OmXGXyak7S3F1tlYQ1EB
GI9Bs+gvU22DI9Bj49rWIQYWrYbOTobRmzzgPXbd5wBm92x/mHLi7GS3x2+k01ff
y+ti4HHpeW58JS63iS3+u+IWyjnTjr9E/rqGNOyBxzONuvE4B8tgtDX2fUheybWx
FUOReaZK91o95oyi0Xdl9ZGfCcKlaSGt9q+Q15B+64amYVeIWsVLgOyj93NjBxJn
hFqMkA2lvj+XI8Nd1b7GdhFYbNuLEwOOTGKzHh8UgI+KJwfoPZH9lR/HabrtbrWu
37bwUW9ccyAeTwiuQv/q6E62GKvSBlrfF4VKM4L11QdwbqYYW10s0ofioYM5kEm5
xNLeLTHwGmaoVEEKyWigTui2pkUPcZxa7OiA+Jkdr+ya1rzSWCV612bdpzq+zYH4
ed0+LjfrVGe+kE2coNv4T4ppKdwljA8UEOjlQQNH5qNGzbecIAcafvZDeWDhwRyC
2Bl0OXT9/wcDoVHJSTFnqn9UWSh1WDjq9i+jB6MQ59DoHWfJBJ99B7a4g5FePouD
k4uWopp0+aqKxQlYRRwg4Z+KtWulBcx0qnHAzlS96+hz2piH9fYa6YYt8s4Iqpaz
pOvGX730bzb0ZPYdS9o01ZV82IGpajgoFQcjSFjlgeoT6SqlLf3bWKY96UpUnPiu
FdFRx2Z8WRtntfsV62MgDESLG6vsB/TY63sFJfwsjymG7eF17Ufzm6dUvrkT2aZP
1eEc824gjVQWvrYdYmlB2M1zdvhSJcn/gg4Zp11vUXOFz0i+W7oENEHcvr+xg/U2
7L4jVGMAjrUtYxjwrf0sRC7AmVVpn2uVWGbZvTpoEoRUVk61bHarBebqB/qRHUWJ
3HmPrHWj1eUudXWZlXMrGx4Uku4XzL3120l7f6zw8l1G5hPcKK5Sq2z1nMyHcuYv
NIWOA26TKQu/BUtAUQ1qeniimyNZtmFRyqofS1plQSV8H/YRQo9GDZ7/4xTh5JXB
x5Na4slG7xN+muSigkflEV/ekB/hSrJsf2D2AIqeCoTv107iM54EC3Ffx2zQ/0ep
CerQM0fgiaDtNUC7Tc2rtv0qkzMC1DZw53t9Bq+FmUebzauNGa/FDMhkRR7cGKsV
IHIQfkGl8b2xCD1yoJvdopbtVL9bXJmAj7S3ut8TT7+GZ+nyIV7ALhhQtQCy3Gtu
KqMlplUForof7nONAoINIYipeS/MwQMXCGDM7lCgFkZVhr4T7fuQ2nj0GJLSZ0z7
rEF8ubRccCsqi6xuAYnG+tlTnL6fSkAMaSHgyJYKBboWMAQLIYW0gTYrTZskVRRT
8bCrSkrM2arFMX5+JO4JX4oWPIiEug75IehxONlmTvGKvFabPifgyCE6x0FdPI2P
Pbe+ivriV2SwpGSCY1L4BowM5dYtU3enF9NmRKkRO4lriVAUuI9Dz5gcDUvBDJhI
TUe4wmI1RT79a35i54vfIOrKM5lm6Zo79p7LR5+tGxYWaYmLci7LZyqRsg9RVtDx
5Mi3MjE5awBmzxn3KLIgRhX27C4wsn+yLqSFsML6r/1I0CImSco3kJLCzJBDYY3E
vQSe+YE4oYiXRuXjuFS6i7mHpa6EgJQLtJaYWhKHqFAfvGjaukCH8beVsp45qWb/
Vwz4ueaQzOYkFYwRHGE9dAwOQY4J+RtsxiOM4nwZLpkDRB/KVSNWuWDlUFRnO3Fc
Qodx2BDO3jgh6brUIOVHn1fI2r3NP39OglPi/YJ4afh0pBhaNOhkkennv6qW0Hbj
NzNLv2Z8o5tZ8/xV7zAO23i3UabGYosLDbzsT9Zoiaib/x2FPRpd5Ko6OXGz6V83
EQ0M+CcbpqZkzZdg61uxZRehvtObBR5GPxwHrExflsLzSfSVEelRhFmvQFm4xpAg
6A+Xt7J1NY1Hab+AlcXiqwc2wPLzkgdolsYsoMOcHOhhsffYJ2k5Ash80RAF/mr6
eXqIjRp2srNc67P1e6hlPSWbpFO1RXIq5+nyJ8tU9n/Xkq9Kl7MR1mtkpsTW5uG/
nyosWnaEWKO+w0sweFTI17GwsZrpZNya1DTLIOm1shBR9X8R0zTUcCmYs2q69y04
6pDvyGeBOuxyIu75kDd7F5k7l44Rb4D0jIuAofv6rwZs8xH1Ld8JlOtMyJ47sWvK
nHtiIagv7pHysLGeXU8OleFfbTFI8ysZog3n5daj5SFQBcyEUL24QLcHd+D+P/cf
/borBIzi2g2wll7r0aWv0wqLzTmGw5oR/iR8eUne+vnjjrIP47qg5ycTWf214wxK
YrHpqLZSSAlDFbaj37xfbqhXnzQIwKFV7aC9SvUu+UbOhW1EunP46W62gGX+jFb4
5byd35lTZ4cUl1u7nIiUT4ijLMS38w17/3V5Kb41lcL/Ih8s19tOYpYE6QcF8/AM
arl7i4Nmjb+s9vVp1yUQOy0IXkBK8MORwGDo2l0J4nODAxPNtdywW0VuC9lO8tro
XeESDngE85vEuKbWinjmU+K+qEcvPDg+FpAJCttD5ZgiY51Zu+LwFMGd9ePhOkPW
2tvrS9meauAWqlIfK0Cw3nKGdVK6DliiV/qL+uzYYBGxkdUoBOiczmrdK8Z7FtO8
hcZKsT3JpMysbKdwDqH2x9uP5NyUUBX44N0Wckjh1hdjEuATvmXpsOEP46FjjZGh
rCmPoUEjtFJt/4DI26t6SDiSYL3y9/MzyptwIeycOCvaZ0S8aXD72FO5es8IpF8a
aC+RuDWhSQ66h4861Wi+jGFiU7PPabAQQ0QTthZhhGlsV6QZc1nEToVqdQ8sg6h+
At64XWUtWK3ZW8o6RWword0zslMDTYcB4Bb7cyfTY2NgzIDJYyu8eQzignW1T/C4
ZMMy0LBDvUObBHAzAjTfDkI0Zy7TSB8lHHHqrZ0eO3UTS7qS1mcuto4gIT/qG4BK
DnDlyR+4OMEn4gAIbb5v6tfichpL+6uBLCp9/nGznGCZILd1Hq8zUGcwplzWtByG
dkvYyoPD6d3it2lJKGSRJ+8+KfiXo/VGIwB1JkD/p4DQJY4luPdrqNNX5GvfKFSQ
t585ZPcdWhatmS/MuUULvdoJSoztMnjmApHfxsOW71RicT148zPQgBxX5VMOQhH4
bMGwTB7HPnxg00evFTZMLIEEBFLkBY9+Yqjn3MGcNUaskchVgpl0nNRNCZGPRC8c
kMJbxzB6w8DgPdAlRZztHLSG0R/0rrSMRQFCUt+QRUyXkkX4iAY1I8MS46fY0Uk3
IyYMnSpv95J0lUEhqgCizsimO2NI4pddRAuNqJnfOoWh71x84whmqt9DImFEFkrv
qEM+jMWoVXjNXE0hCTBi8ZNql7hnDNSva31bwpma0oM99MSvwdMQNpJ7tUVdAcGD
U9dZlJB9bFtWDucxPB0w/mtxkA7+d25Jpe60149dWpL3WHIHjuGiqTI5bhBG69rP
hRkf9EmjsbDJNM3B0kXne4I0rAvvjaaTEUHyQhsuRhKP4iPdl3MVdyQXOiE7KbFG
dPnYGI+zqOn5PPBq4iEhvi+XWpD4qgLnkjXsU+1IUquojbEe5Sl3BvMi628RAkvS
Ast/xm0OHyMnn236Qgl2aCX6JSSXcpTgO1yFQGNEsYHJL7aqPt8vSq37bPlFf/k2
4PHN3tifNnaSa3CViedZChL8plekMjwx3hDxO58PYdk2v3CYXViLUot5jFlM1F32
TP2VVpmR0iXCnVaKZ/y78tHYkqzY5mgAxu29X7tfZ2IvH73F6gkv/yJBLbWrCxu+
24S0MQU9t/wFCi7P9JfL+HNzILnY00N5i3w7i262jOjh55N+BJjt9WszLDyugSIs
7qk8YzVz4nygsjUR/c9QEacZXkmw2eACii+OdqRduRS7tFb3n0H9kSvh3QOYJ43U
4wQate0g68oif4/JpbUMDHrQxwIHSgvO2pOGgKnPpF22UuBClxCb3kQgJNBCRZEh
H3/MTMqXunyVvHilwrLM0g88AhVv3T1VdWv9YfDFgc1XL8cjSlEbjpXUEQ5PmsZo
V9atkWIAQIBA3Ve+4fAvkdIp8W7WJl6WhFjOZZ+ET+90ccO8goahNx/DfRK61He9
2/Y2JO13Qi3m9cVZHaGqYzfC0PYiUls5WviFyt+dN74cQwYAy+zlvglroAwqaeQc
zaNT+2d/GkjXaJ8q1ibkI5TokBGMLcgu9I2zKDkkUNr2GmB/Bhj5KlGu3S2DworZ
NYpqM8cMmS1VCvlhFEQkFDAfIi5Bi8/FnBL/Ci1u42uoy7T/LYFdrxQ22hgNHwHX
FaN2Hjv+qB4rsQNSaqS/oJbcNwgni5NFT0IHXaV5bx8ldmmGkBfzyT/5qutKfOcn
YbRXomt96/35X5FyOEreGIxh2LnwW/ENlv+uTU/l0xIJ/Ln+7nv38ayRrRP+nADN
oKQehsbKTVSBsQInAWvvCgjZD5/Jh+Dqo8sIV1SIFVmA3UHtqDbwkzTxeZyJtM3P
OGlwpuhd4CqmfDbffC5DUc5pOFf5imzDfmAqjJVjBBPHupOGiDOQ2RQ5jlNZoXfJ
SL8d09VlfkWE6YYTTn3723y6j1RU9Sxpfz4JXjdCNDgrylEa3yhHtAF2m+nh5RBw
bd6nlUFxdWSkiB9AUaCZm+ZgFaTPIqpgwuXyRAZEWNHt+JcmQLz2arUt/W3qXaS2
7i0hyE6CZgZU7h3GoO0MaTVlqBBdRT2W8InMRVbeALyykPg1xN/7+FwPI7WX1VpP
0nCOQb904s4FEl4C2paquETANIINenZ+W2vav6fzEXacSb8U6Bw57ZAurTE8f74B
bOMm+jc5RJEdPP6CTvCqqJ4uCm5EITYzSedYIgUXqKsbBlN8w4JgotpgsM8Aa84o
Il80JHMc94wNrbee6//2rywQrTKpWitTh9K87R2NswUtMX9ePkBwgjXwklEoXIwL
NFnIPvK2iFgCOO+IYc0IESB/m75E7CTGkRAXd4Q1YrswrE7R/YkvCZwHqmt/YSLM
i/DshwLMg6ujzko2PhB+VwxSFM1q7KbCeX/Zm/eeNo54i/XKjGMFFVAnUdLJ7v5o
uzhmwP8fHyExP21G0d1tClO3DRN7TxAV+SwfBs0KiCtJGIDmuv1w3TQ8zLS1Qbgt
tq97vWocoiexetjXQSejjLHXLLiJYrI0HC8Qepn4dTH1RnhC8fe8MJAUjmmz3C+L
QbJHwl5rb5EmfYpDTqAQO+iSltShrUUiYRZMSCXJW+8eHXiT5eP6EqtAtq94gvAN
26aIY3pdd7CDn4ZHIURVSFw9Pt1J+i2h77nE1P+slcshHCx98RspZcbjkBsW5Uqu
BjrRelnOOjZtZsBtlVaGu9SfokaoUIzkLY++QxlrptwYxneDj+V2f+NG9U/EjcW/
uJcV3VU9IXpRdvWNqrcsQALx5HQPIn2QkgU3IkMhvsgynr+tTxZ71N7rZkyZfW8s
5wLrkRwyZ1QohM0C8b0kG7KNFFXdYy5EH5IC4uP2u2ROmIjUgzTHCIHjOEwIlb7Y
PgIdTAm8/RwKe5e6lmlGhchYZThUNH/LpWwa2dWssBWUm+48UO9naJpjFUpRj1XH
MZx3XyeNhc1yRypEnOaW+LgY68NEnxN8WfodV8V6KduQ7dXpg0w2KbGIt3/7BvZr
6+N7fl3IkhyUKaa1Y7Z21nfuls6vuA5hO6CDbOsLixSDTaP7uo5Lv/MHnjUfj6Eu
DT0hyRoAn55L9uE1SyHkt1wvqxnAAo9x6JPW61XgDhGp9XJxEs3dNMjpc3ZpW0jF
ly4HHzaH6SWWx6c2KsDlGc+v2ST+/Os7foVEaDFAej5oGsjwnIJ1cOk8lOmELISS
WOZTkB1jmGBi9fA1z60UG8LB9xCNm0pqUpVOv9W38UeNZk/JHDwtP1l9nTLxr2OT
CERx74SlG6/5J2+Gj0hCaVeWxdyv1AszJTpvXtus1UUayRJnbfDunSv2+qb/Ah0r
7tzrsxU1PGbfa0knSX15dkkkZkF5G2k28gSM+D1CQlKvYPiBv541Q92GK80xNJs1
ICfDhPolAioyYjlpP6VLIM6HLwf8zh4e5P/a97mKbHr5f2taPD2CsewY85h3uLlC
BbiiOidBnzgKbf2fc1G8iK920zYlJFKeICB2tVwEbDYLYrNDwxrdV5JoBsH6ujBm
T84UrsJFbq+airSlyw3IMPKPdPzZKr8bLsMDi2oOxYG6MvW3/wtBEQ+Em94Pm+bN
XzsP0JEDRezQqkaPmePOE0kPGfqIGIyRxjOih0ABGzmvP4H1FORt6dGFb10TCPuO
rqr2D93m9ZH3l40j5Qc5OQSGk2h+OGDO06//gVtVLv/iSfL8Uty+Gs6Jg/c9xE41
Gau33dlhikDg7rt9+UvINHicG/LjxO/y0gO8z/XBAEfWeWpXQRCkEq15MO4pVBS+
DEn3eriAGJROlFA2pJJFQha2W/3cBBfR/N2b8C1VZdWfsYbDwqGZBgK/PmntwNxt
loNOvHC41/MFnSy5DWBeZmg8ay0JNFjIixFf1aMIWSDtsQRwbB6qz1lHDAytpILN
4Fg8PGrY6CFshuD+WFNF6fWbUxMEMnw7A8WM43bBgKKPB/1sP3GiU7bc8PwK/IU+
lHzN/TzC+TWId9RfhKTEJEAzCjuLWEscKpBwsj7fUeYkL73otxfYn6kExSYJ4ckz
MftMfKZcISFe7H6JKEpy3cuUuBkL0u9C8UhGSPeoSv77FAqROVefFLfi7jG9zL0w
YBusnCYPCZkLUCn4GGJM8G60v6j6xTz9I3tKPv4jok4/XMmhAGPCLgiZQ1rc1coe
4lS+a4fsc0s4Jz+2VEPKtQJrXlx76jDEa20PZ6kN96s7npGk3rSiGQEQkqOiSKb+
Hv/P+BSNvbgvnOI8E+fr6adTkcjcdn3F/hoeb0Tn0Ug1FDfyJOgu1rCdxYJGDjRa
Yl+RfeKeLV8uJtGzjxaxBanYB7vipopxAzz6YljUCFLcYidKG6bYI40vC00VtSDq
gpf+d+3WNq3iYQ7GTIVG1oWlvXefS97RZyLaR0TovILRTPWY+7l6ZoG/lAoptNnq
0qhOQlpKSgSGmys1oLjb6EiGPXbLa4CPYjpC0b8o6LjuYcDcZsCk8FkwaEDLqllY
n9uPoblVN6D3lO+HIBaJzVc7Aob5Mnmx7iAzHPNmHX+md+YLgnctoo97o8SLGWGX
heYR9J9KWswwu7exZ0m2ios2c+RrzxKqMHK7fkpYa3kFRKSDFdw7O1PaZOeszudQ
IK/4mqaT6qID1Wy08XzmXG+gmI/8c/8qmEX7COsI629cxJ4TyFcluSGMMCVyZQpa
9WHc3Vazwqe+Lwzq3KhJGvB2w/v2x8vEKCb5sInWfs7pnFMlGPeWPu+nq1Bl504D
VkBSYaDGx0mULUbrtEjl2tenKZttcGvyXvZACmgbbPaYAL+seEJ2R4CwqKdnl1h5
KwAuVrLJIGI9gn8MKubiiVAWWCoo5e+xfxTd69ypRwZ+/udDzhYeAEqfMwWvlTyv
rzCL8zl+fOeUBFQIJqsStu+azdJTbsceNfwAUIRrihoTfJqUYfXU6ZgBKEwWHr+i
iXfBg2zcKVsP/fNc57rVueDDqF+6OYs+1dtwbLWPmoAToh1F9tKP20xNIUV243D8
ZagXom4UfR0hgKyTuFAxVq/daAGfq+6ObBmyceVJpYIrhN7iHWgydeDl/QVn1OP9
BxdjXa8/1EEITDTIfxfHb+05cXu612kqKe9i0uMaukbtfGBMNKGJ3vYcaFEvY7xn
53VJ6EAetxb+lbnp8gyyJPac/rDvRArhwNRTrpfTAigR1yaaInZRLYFxrzmwNQzG
EAOPTiZ7el5QQYTPKpN+d1utLvjYZZJ5dKyT5dD5vqHRt0yOqJibaSHs2SCXx0OC
pRa7UFkwB8osPiudALG9lpE4d4bq4YsSapitaK/sxShzKKkWl8YiYiEdxZt7nf6H
QINozXIOHGyimoj0o66VqyLbggd3HWx6EDIm13m5ONtoifRCNWpAiSL0Ci37GAKE
LWhgcZAcGhM9PWyuGHaE9MsC9mdANTMyXri/Gru8vMGmsKw83Xevw3rN9USUCMdw
wgALIQpmuGmR+CQmF/4wufz1B961ucQepypQgStSYnSmv/CVb80idgSLnc7TY0pS
/G4IOU2wAKrYh2pjMdinll2iTCwoiNDRKk8+CsNN2oYtds8PcgBBon7iKotj0YIG
1MAvlFCvoS2oWZvQDWtKV4nEDIlScBqimDa8nETtALLKZo5zPTjnGQQaRC+8XeFP
GKVAmc7hHMj2girr58bZ1LndQR4nnxeyZvjIhVla09mzkINYFQnpBBBB42w2qIEM
5oFwdv/var2ON5mz3YXuHMActOgz5VisffUY5VJ2Jx5WEid8BL4tqwdmHwYq1QPJ
YSa98pQRFbX0GDI4Z8WuphpN9QdTejwRuxGgCROG3Rw0MAYCRsxwy/sN5MbmiRlj
5GQq0jZxFX9KlshpGnBjUkKopfL4J8aUG+kfwsrzkXiuTp4lLXffSYio8S2dPSZK
154G1Xu95SNepgZ6Ypo2KrWrah6dxAHf1b+7mYPIXvLfBfdcYVlbVsCO4IHya23n
illn9mVqHZZNEadZvNW661WLTMHDkcmU8jCd5JyEJ1G9HCWYRVY789Ccdm6sWQTd
opWs9/whuXDwHatHxIlQ5EHnGE2SJzw1/sQcS/Kk2a+5KmAM/uhT3R9F0P5N1kXJ
P2/sPZoFkp31vReqkLPxLBDaPNhO5E8V/IsipwUNaiiACKVBoLVoX134bQm4qWpR
2WYPfdipTjxHpQCc51wHiNcykLK7d8PuWKcaP6eIOptqF9EU3NlJEUSOyXxtT1TQ
Zf6hrVX6wZQtYmPZDsFCn8cA6BJoYr6OaGFUjgnyJTZEZOI8ptFN5FIP+mnELLhl
3bgiqMS4/eQ4q7nvQ1w618MWSh+Pv5EiS2LMOh8RMxw9ethNmXA4+JY3PvZk/evE
qUpaeqmDKdu6zDvVvK/H9Q6AI2I8iLaFfOoqal1Knd7s6wc7jMmoKzr9P3oumPpR
EbNFXBiq2ni/2H6tufcf3vGdAgUAtIg0cTetftU1FFL2nWD8YQWkmGzg8aoPZ6wy
h7WCcaYeQBUUxkHRdK9hQol7Dx+ey6ywxxIxvgcGeaWpG4Jhnq7PASjmfT4IE+B0
v+2Y/6oheV3mS2+uQT5mzkJDQIKXxbOgcOu+iLGLQ27eNvXJvyndjctGOzfb+9SZ
i85vKsA8juiQ4SgisR+1waDhS8E2fsbv11FXd3yfQl1j9wKln0HoUzVBg/ULm05p
Q/XdUbUEkidxGuGC71jmIVuLM45m8gW6aWPdfxhgpTF27epKtKpAF0hFgWlt3vZV
C8lxLOf57yf0HHwSClrXxWP5R9/X7udRGtuMlgOf4XT37eEKQ47IcJY7UcjZqJyZ
6VZkBGnTztPa/+MXl5WqdEzFRhqzWclPh5rj4USMp+cK16BBkNEhmM72k/DCK7Jc
QueR9DMhaFYgopQAJ9rFEo/HZbnRZp5oFA+lv8QBbutDU61YK6vuetMVRHCstGD5
3rkoDkdQ+OPOTlsosk4eVRniUS7+Gg5JAdVqfEv6U1J/tAaSQnnfj7n81awvF4JA
1Ysd//9iGUNC4Sh46z2dxqsbCimT36Rsm1JwE2374p7l1cwT7nIpQ62bGINwgv7s
cBh0LCuFdg7B0m6lOWmtA2pbxOSJKTALYwCrE/Vo/+0jJjoTXMabROzzVnwyj+BR
E1zyTCdRmrahY7tsTKJS1U30MCAkoKcV08Tfr1RN0/oqn/FsKqXv2GYiYgSMsGyN
b6hzuJ/lfPwE7osDg9Cz6Tb//rtKrnbAv7Up2GP6KH9YKjHIiJYRUuvW9qvT8WE/
RVaCI3Ig7V8yXv5nKmRlowW8m208FLrzRl7p9DwR7rhpiyqx0mTy8WTinCV9Lyu5
t8L7jZ4qNobZS5yc/mkzL4TYg2oV6FlA3DlGBT8fyUY6BW2hJ4W9tF6TCOFF1clL
UF/fZLYfOo6TywU/PJO6NHVdMd1UsEoK3KFHmFQUpMBnjWCG84Lujh/Kb/saQy5F
ZRpvByxw/5GQPR4fJ7KCaRntSEyzn2WyMLbTHLZoG54+5xfjGZ5Ux7y7Tej/G2qy
JuahSvQwX2AjflJ7BkeU+rp2MyFTNlqlhBEdEzHz4P/R5joUeFxmuCV+WbjYLFoC
Y9Uzkbjz21PkMJPdJyxrdTpg0T0+sTfaR1W1zYClohisnQ+9Dp8JVuXFTjqZD1Go
mcHedjNKHuBnFNqBxSzIjQ0H7WLvSOTXW5rJIRh9paxE4zzoGBjYmyLl9iTm1zPB
Q7hcXUu+YLri5vDBjCdtt4+JyljkeQzWaSl3fvkvyVqw6urb8HCREZv3ySHpYCvk
HteLPJctyEIzUYSNP8bqt8mpxjoR+zIv8SpbRO6iy2OHjPxiluI772KYs16fNztu
IMMk3kuMePza8Ep3WcAsg4guj80RHC/RvAf9AWt0gQul5gO9WC3TAZ3UeX4MnjXU
xAmwZGeIPl4miE0qQXg/cFwlvprvuZ0lBl0lYXOQhVE/8auKYjCbESAk+uqcgj1X
KcE/YA2QYUQ2y7rKXv0Js6CNfTuwS09XYyq2V0fLyvq/0NBqq1VqPy7M9cECQnXv
KL6rCTbBEZliGIlj5t4lqsmY5UmvWmReK7vIG8rGxQhYUPrAQCTPdXib+YtVfOEy
8GnUtC8umvirvwBP/iIxF0zf+baPdrx6ep2+IGKQqDuk92SXJAYDOKzkP1RF+BX3
82ft9DLKawNI3w5wzbxc8D+2gaTjR83yh7PGcxsfmitab2+EhgEW7CWKhnknG+Hp
DA1WrAbzlctmWboXuvPk3dOCa7OxqOCJnBOCQqZ7qposoj7k21SklHErBy6msPDe
St7PsnZ0ex/X8IT1AP1zw+mGQFk1ggpDsL+hd2LCaRxW2H0+a9RBq4nVKjWJQXof
2TyrEHlP+INcULI+eRNS3omBzyrsY10GlhofLTVxT8xK1rckXOaa+bPDkeIsoKpn
wIvZa1xIRHjmPM5tBiCnX486uTscLTEnPtvPHyfERXXEIxGNagZz3mGNZ8+wddsr
k+vnlDtzZ5uvl48KhA9ajUah58Yj9SoeNB88dc9WOwsjj4Sr3hKfdqi6fgf3/wI+
NsxxraGK0epoTpnyKsEmOrVaw8A41DM4k4w5wbGtmctu4vwNNg9oxwusxeaH8iwc
M/xuYZ6cp9bdKOWkw5cvB8XMkmbnYaQzoXKFvarDKkU7+u2YgLm2cbHt63tjVqXh
Kt++kG6MFF5zT1NkQa+oFDBB9VMu74laDnODOjGwCL+yN90fZhrGTctmL108Kfr4
pyMj6Md3/IkDf2DISPKiVe+AOi8mcsuAhn982A2Py+es8KS2BYHU3VLMKBzON0x9
3+1kRfsk2tUzcNv1izggc+PKtOrAkJPi7O4LuHHJqwq6yjBdEeDswpe9IQjtKI01
8ryd6cY79T0dMM4cY7TEWJ+T930rXpD1948MuLE895nUfhOpjcF3Z+wt/90l3heu
I+NIFxIBfIGPiOhnnjEsD0EM8RnFbLwQ3vwaVDj7gbYg/UJGZLUZ+PubEYCELeYB
xcn1xBIsRjsyeHN/8W6IycfeUwpxBT8Hu1/W4aRl4IWgGT4dzb0jJPpMHb58I8+r
lvwUV5GFi0dYZHsHR8ePlDKdhd31uZjzbk5TjvE/GnP57vUlSAiEEiLqLi42sKsS
QVkPY8Oa9SRtibW8VQ5E9v9ARWlwGl7oDA18La6jgi2DlXcBXBFe9RaacxAgAb2+
mC2FH/Hdg4wvDwPPQFe2Nbc2AZQYNHwK63RyriRlLa+GmFB0vM1rylqVBifrET73
nGsadh5fBa6+ofYGOFyR2oZY6R0yehBGS5v2ljjNKDk6kKNREpHfquh817iUTmSe
Nctj8F6fgIJB4nrSmo3MtMEvC29jivOXnD02nKYWgCLIFEcGK4qVKgxVpnLH5dsp
Cg2JLIVAeidOXArUQ9xNaD8ply3MLFopIItnrBbnKFPnmj1e3NdF1efzJfzRpPEk
E7elxmsW0MydF0XYX78d8vp2QWv2+RP9Dz9Mifn4Ez18nKtY1LETVM4+rBAerGPc
9YoacXVQICKQm4P+ECIEYRxJr1bTZ2UZcwCa9TwQnYOXOLeRzS8fq2ISvESCtGvc
FodrljnIAocVwaqJ9vFVO67XnrOahuX4AwxbRxCOfrgofhbx+bjhpFQdpr9jjYDb
4dfpBawU1X0Z+/e9xmCDztz/VgzWtFG1xThjcp3CXUefR+dLue/RtqGHO0lZEEPj
203cWdCD921t0wJyJGYNNg+AZaGZeFv9r+OZH7TD3bRLcRh0KLpIIRncxBoHK+1K
divnAyfuPBnJmmyM2gIvE5h1N8D35baT5v6ufNQRJz58XOnvggt5CWUGAnIdefsd
4rpVFLI0cLdj3zUX7wjC7ipem2kDYrbN0kHH5Vmczvdvfa1GfGZePmkXLwOlUm5C
XWS6d18oJIzHmXvPaq0iAjcWArRqPE7z1LZtqWsJyqitl2z2YInmX+0pTWhyUpBk
K1dcJ5PZRy/OaWvUPCxKJlNgKCPK9MVl9bp+25+UPkFWRdydrGzRr/vr0ObDpr1M
4sYji3NlndlfYdbkUZh74D3TzHYkn/Pqj0rm1lDh7jJWEaU4C4Z6kIgGIe1AFAsT
I/fi27oKyUJO3/nhKsisNiwj+4P6rV1b7bv5HQ4W+gTv9HsB1w3U64pgSOyygNsg
KzyA5M6YMlHq7/+LXdQkQMUR1ReAb/SpWWZqzGB/KfPW/6S8+eFlxIDTRwqe4u4r
uA/F0lQ24yYZNcYli/nS+weY0A2vsmzvXzLK2C98eaqiKmizW8S++2foLdfFaJ19
jr8kOf58D1gfhzNI0+09CEp8LQLjz9VC/cvu8/ZjlWxktrmiVZLay5oJGnU1lOAo
MHdUjHpi8JoUshf3d8TqJP47Y+cIbHfbvhhxq3zBK3gKGwEUgMAzKQSQwQxvNtVj
VWbUjWz70NfBQnQVEGIKpygr1fXEVt2uUEFfykSzIFnPeNnuV4Ph3vhBgHYwMG59
U1f6SBVSQADKc5CVukZg4WISou9WQ872w1vFIYJBXYSLJaaJqftSFo1WZJZxARyI
q0aeiwj5DcuafUafRUsBNqsJkfge6tjYRrotE5cunPBwocQFsR9WHF38+d21ieBs
D9xRyoRJYPgRIPUVv9oGiLLpWS/YJXynF5kiCMnI2e2HvQJiAKnrkf8HFmdhaJud
REeemugwKyQS/1LoZQhoKYZSgQxy3ShrgW2gjdnqN3SFM6CUTQ7HTswGhytgCagM
K3/beUilkqIz39ODIebCa/Ds/A03lHcasxk6oPlb7TH+aHiQEx97NHrtBp5WOS/1
TE6Hoc1esuWVpczjvL/M8JR+Q+DAAnQEWkVOhrk4ni2W/beL/jC/ikMXET+xVoXB
I59wREpupGOsfM3lHVrTcNABOeCMc/+nWVBO5paYSxbiI34YT2F9FOqHOSa8PH7E
veRA1JgYy7AuNE6CCGmJiJMjDroH9fO38bAl80y/XEMMtpwsfOlFz0JrRU/7zclb
4uJf7YUyONt+9ib3uMyk39kjvUQDvB1c4/F/983BrObkF9YDIzw/EcJvJb7UQ+iO
9AAqEz4LsO3I8KOzo85Xkro3bvuWsVvFmyToa3M0mDJn0VKj7U27NcDvaLAxPoqo
gkp8jTT8UWC315vySYBSMf5KRHsRTYU8h/cFbNKnNkfylZ9QumhOzhrcFslZIK5J
H9YlVcIAg3QUAA7fRxaPm1ovKmpumDsLy1pnpD0ZErKCPVqjxrBT7P0cyyAzy4in
HfSJBx+DpxsIzIy/xjtWntzCSe8dnJtrN3gOX8Nl4gG826Q+FBCCZUH+lelYkfCv
TDG+iDy6a7SFIiBib1AZmAmET4DRMqqqBgNBrPyeIg4cAyiHbQ67v1m9S0kFa09u
+y79D3Em7bwc+exU3+WmLUz7VBgrX4EUoOCsb5Y4l+1ZLs7mNKt0t9+epM0isPzZ
ygWfl5iL8zssvNQGVSSILTBdGqIjKIbdXcSLf1m62cx/XsuABPt2D2WacxrQCv3d
q5GeoVDvS54mUG2y4eFfzGyuym2tfbu/4OAfyZJMrDvPjvQJkWVu5Ht0ckq1mHBG
hgyMAfR9ME5kwQA/OIe4xPntOPn7nYOaTFv22nowScrHAY3vjMf58Zex19FNsna2
sOjq133lmOhekhz/GjtaDo6hlFGC5z9mYP4KV4t74tGLs1a/EUgJVFhiDKq06spU
2gyFWuISxZoF7Nb+I1Qy5OZfQiyvoZMUVB3Y7vVqW4sld0DMgir/thId3ujCUyVT
6GsuK+sEwjMP0e2cVXIdK3hC/44IxRSGxY3rOKOWAfCc9OGdly8Asr/ON2c6ZTL8
NQ8EXPnDUsQn4u5uY+mPIKt5/Jgqf4nCkx90yw2Kt8UsH74dQ1mH6apLMQNEQsDY
hph0nOTRbNwaQdn1iY5PWc5Be9cu90ohDdhB7jKjvegCc1XMytxqr/ZLbI1gQy4s
2i6C/cN8elpClJFRlL9MA8WC2H4FmWYyyp144j6DJt+kW5vgcXoqjUQth8ihlUXO
5VH45G0O4lrtftMiCxykUVCls5F81SwZ05e9+ttmvCT4BanDCa3xWxkThoAtSUK0
7OeGF8SKk+6iAQVid0ydYaWanYPWE8QFfoKZF8tulCkgZJJOO5uqjR5dxNcoGdKa
Gg0wheHM+chB/zPypTMF6iTjyn7ipi9iU1tCq5H4UPp9yzJYC2Qu6+iAkB/kH1pI
Mnnpnk2KJoIADL7pG1pRbnApZfqFjWXlYCTgGJ4Xw410VLLgvMbQcVwWlJZmoN+h
Q767gBhqDa2DRVs5IXt7GHsyKU9Ilw/w8O+iK7Gq8Rr+X7PMgH7sdMJtyl2XSwuY
13brEGBsxMeS7DSgWyGxBcZDDDLmLbx1EYhSS3MIu0JZBJbT068LyaBWqCTULEK+
KvjlfPfRtuA2+VIqg4qz4CB5rNTPv4CSuQOJjGlJWnZ1hDR0Ztb+6LB18vRcimL8
aSb65v51BoOi+N48FSC9fF663aGWC0FeLvPb/dUsuins3gN3cv6pWJafTIzfCPG8
Eb1cDSqfpeO2G/mb4MsBoswAPloSniJExxV/ZlRuGgNps6LK3fIG+zpfoOuNuGSC
hadRnEch/3v7dXwheCh33c65EjoLCKYEsRj1L31//M1nQKNlHXliqNHsQdPQD5W8
1mYdxxVLVgV6Jc4Ltz/rHrbWXO4u2QMc6PzP6LA1oaP0AVRZGCRkII7NYTpfEs6N
jMqoC66bs+j9mIflwTixqg6O5Hgok4tfrCZK3ARZEqmDjk5Yz3E6QU86yXUfFeVu
sBAacyfvyPx2KfPMYm9yWBdi5WKRPZQqQ8piu+SWLKVd8gu6wLg5hEGqEN8qxToL
s8bCxlnmMeYAGy5z7kFWWACHjuhkhTfL/NnTzscJB4IWkSlhsLD2NrzYwj6TBJa9
etBrqoV5qMEriuv5igM3pgPnURUIzZxEbijvG64Yr1QBKfMnYNS555bOunRu0apc
3dmjkaltwjJK5wdy7ygyhkOhx/UA7txdi3IlxCrXZnBk3D68yfiggPjnki9kHDpq
hkA+azZTRyxp7wTzxWC8qx0DYs6AXG3nE5Wt+JWcng2FGMVLodR8fTPMV2Bv/h0Z
fSHZ7KtOOY2hx6WpgfIY4m2x6Lsl/dfMul9A/0/IFIx0T3j1MoRwJNnUfhvam/Ia
icSMvZjNyhih7i5Iy511lWAFtROyGQ38wM9IjGdhwUJpApb3M4O8TxP0KFFIMpuG
bNaBsA7BFCA9DTyaSG3S/uIe8Cdj4ODS3IOV27u8UDOp3IwhYc09jPsNvr36DZen
idyZ/Ey5z/1aPQt6ztSGPyRRAPi6qiLiGVdcag9bWfJ3mpAoro20vlGVgZXR6hrS
dSEL5WDAJvCEaLFjXhLFSUSKDQ8sMgdCEeB9FIc1bPe7tlWLvQ+vT40nC+XzdMYR
JQMaDdYUmQY/Xk/qbl0D/eAESu3fIzcRis1QOJ99xld82GnDCVZx9qlYYmV8thas
0GXNEsyynQtKRgHRM6v3bXwWFhJynXYe60FcHqjpsZwF30K/WvJ69gAjV2ofONQ3
S5thKiX63F1M6BpQxDFSp7JiTxYoXt1zVX9ysZYDe6a6d1gGUwly+ITcP8PLh2vv
3e/FeeVVHJ4pPSbrZGZWUuOwPW6tjGf+dxjxaoH+cU0J02hV40QmnLmQ7S1eGjXs
W+Rk79T2e0fe7htH/vTP+P8+Mrkext4GeOut+vmOH52I65DGknKxTX5eb9orqSGE
DWKo77PELZCph1HJSA3MmHqA3kAsCnbk0XO50aa71bQzEXGkZG5J3TcQoO6QUGCG
wBzs6fd+/amfV5RtAF0VHQV2L+QfrSHYug9H1pyQ3ExPoL948gXVPzlnLcalvUM4
Euw4IkMfWiD3o9Ck8JDTSVxVfdF65MpE0I1gr7teQ37y6CBN3+zC7ekdzQjBJmcz
eBBaYc+Vi5w7QAgO2i1xVcaJf8z7BehEZSiZ7SBku3r609lrN7HUb0iReoNOvKCe
P+VPjRoZRwu2TzOsKTTdBgxPtCesppalgHIx8+2JbF1vYxA3wiyGG5yslWXC94TA
RPM4FfgW3/4GmhYpmRApFOjRPXvZranC4PVuS5OG5y1hlACDguI3J59PzZi7EBCA
28PI6eU02EF7X749CB/5ktfgfP5kO2c6ApPYsnwNKvYfhcQxXR3z4sWo4x/sbzKw
NVJFecHczMqQJqBi//pHcbP5Xd7PZ536T2QwVasSwDD9qS0ws5mBvBeZpfbOT1jr
0s4OgAw7efhJib6rLCs/l1i/ev7qbW9sZ6Am2CnEWCyMzVmoAlKXIMOENgrFSAjV
wAiVFNWXuufQ/4HgLxu8BP3vj6OjBBj8FNNYkqkmpmBV1n6YrK63CXM0RWeRpspn
OGhkm2i/camsmPBm33OYZJi34xpEaTl+ox2tDTJ+07bE63LtoHtFO7Ai8ZJMe9Y3
4Fb61J9QP8CSzgIRtzNSmfHsTeCAqXXK36oFo81Cz6JlxDJtRAmiUHaAe4H15Xaq
PUUsDYddgaOVONsFEdBNW+R6+dhNGjvvJL8SPRRfPVuNEJ6yd2IczLiOEfv+2Qtd
T9f/LQvJN4SRo5QgsMOhPukIQWdvckK6GNIb5ZYyE1BUq9ZSin1HpIVj+RVbz0D1
LuqkY2wk3QGYfETB2tmb6IbyQuLRlyFZl67g56bKcp9g9kLqaldLoj9c/wuPqabY
D6N2CnAgbVEkOSdkqje80JzJSvARXLRSWOpsudPe7af0BWQGe2dN8TR8W8gY26Y9
6fnccN1CqJhDwDRZhMXSEPgLcKKfup/Ak0etzl9ky5HMiemMLCOrbij9agqRlhzf
DbMDW51nawP61ZpLkiOlEuTlweaD0dxjUSwtF6DOaLhkz5WpMrMAIJdV8UDgChQ7
zu9QQDxYRE/5wbHNlsx7nHyqM93/zgehpNlTp8GkyCfAI/rcU4gd1F0ZcKZZfPKO
wGJdJy/LiSyVlT2X3gTsy5sTfT/DB+H5vf95EdugWet6tHVOPtZBBBLBS9xCel6s
0AoyoZym83X7PH+ZgIMzxDGesV9T10BNEWmTA8j9KBF276mzQh5BZaL/qrrRDWbV
w8Y2LKzqwwroAACUUILnK5WZvzJ17wPD1at9+f2h5NHSNqBr24LTyJn+uYX8Z7VI
IAzrrvPATnsPSb4t+g7bLwUapwSRE3KzhG0UkfL0SNzxU8MgpV/aWah02367AAYv
l9mOlGWvwyHmWzpAz4wfiicnvAog59Yz4Ah7l1SAvSb/o8Ne/wNVeOyloXxyiQ7D
aIlQ2LO8InF8vDeOnHjswPY4Up/4HPbNVGDvU/VI403Z2GPFniwuNdCd6Df0aPSP
A5jsyZLWonZdEA/WESNxTknd6XD7rJqdn+7FjPtoiFG+w8wNg1TUaHoZCDa5RvJP
Ib1woC82xJfOa+24ZJb1rjV1jKxN8H0OiaFNNTqXjVrCYIrXo8zkiIuVSoM2UhLr
fMjkHaELsbee55BVbHRLZddU9Pg69IBtBzIRPvO6R/iT/FKrE4Ujp5tYq7hBFZJD
PIQM6knj9cwtCfinU+JezkHjNPrfmEqVovMCU91fh1YvU4GjA+1/qXr0uV3wnTi+
B/wYuAEj785cMRUYCAzE+72AvWuJq6fgRSIyse98K2eOJ4/irSLuH5WmHxopGuFg
sJrfYNU1S1ogqoMdj5+vcthsL+ceT5ngghZOM22xUkJoZL/LHR3TeVadVfqmxdXo
u8DdOC9wxjLkXW0Q7fDN7cptIxpMy91pBAbkcdTUvf9CvLLA6bwVVBRi1+9HXj+a
4qWKs+OCVpH+qkvkphcLRVWHm3EQ3Ug13wDk/GlrguGKKoZyDymjcPyN7TCH+SdT
QHZm/Ax87ffROBQYFQs3Oq7zZLyfa9NiUqQ/InE+QuztIxpBQiU18awUY/q6ZRFK
a5KyfGBCawM2axAqTkQshYHOc5InsTSENZxUEe5wmqFF9NBdoNXCwXt+Y1UXSb5O
4NjluMWXYHhwnGLqr+NEd36FtYVp6GSrrqafXfCDTK/wPfuWx6v4UeDLgcBix+qY
pDNiMmbmMT1O1C+ibldQS8BRApmDl+ok2nYumfCOVWhmhkrTcnz45AQDt1njYMoY
zcb3uAoUkciYWPOQ9PqilNwwqzU25w8m6d3QSMBo1T+Q5pi6Rub3WL7PhYp4RCqO
bRXP+xvPha60LlCJQ7bD2HXETmjUOAS3/VwXpx8Aht8Hd8YWsrgIoPw8Aw+G3pUG
gzRoV+5vJsE1vpx2V5crlMQ49BLpVoz0V51/rxxcK9ifRVce1198acx+W0Jw2Mje
OTu1BZOoisAlHxeG1kKxECGNgWmbeNLqYu4rnBF/0pCOgYlcpXpD8UapSxn4mdV2
OKjxE1XWVVGD6fCgsvwOHXrJq1eD5GZ8I/NZJFk4KLlytkYinig43rmOLyWoBMJJ
D8AlZ5I0LpeG/2Q9Mk3OGpOFr3Wime/30plj3c16/ouVUKqu9yWOGrDQ65vzpqpV
1eLXt/IGfOx678L7oK7kiVV+pJIe71sNvjmmlhBTG+dycYeHxEiAkE1tJQUTyPS2
FQZtU4y5dHEA4IO13TeAQ1FC+ifrVOhvFvXgWCyIEdJmmih9DIS5UK3e8X2aWR+O
NA6MijMTmvcfplm9GieFFA1n/lYD3IfSD1UDQmGGqn+QkqN6nl5IvLYC8UuTFjoP
CO3jS+JLGzyYYHBvFBJONUcUt3PGpkjeRwpydHN83bO7IhscVO5eyFgyF8SRSUhS
8e4a492L1zD7RBeYAo4Q/xkKF1uN6WXnmAK72kJsY1Y+i+XVUf0Z0xHbyw7ucdJs
RtY50ivr5fCjJkzRZTcSpAhCuT2Of8ewuSmOSB+yiiHejOMs21AzCGeYubAzje7o
nF2uM4uWWBQcVU/aSseHuS8f3GB+ffM4wTk3QjQ8IS6WC4AVIUW3N4s5h+Ze6JKZ
WefoZgjactSJuZU5Y5o+ssY+8y+WpaVBJZhFB7Hq4i+KKVZycKYoVldsxSZXNk6g
6Vw/xKN2cjxmwJRk/bobNNYpcxE67y6cTfwZhk+7yvezM+DYufiFCKPvSVBm7n3l
yR6ftL/Zs87Wrjr1UBun6AtEWw2Bzeww2WpxURXZ9yejlyMpbLPy1KK1e7HLCbhe
+9gqy826HdeoH08Kiyv4IY7J8nNJslrQLIiqnyeO3Wj76p6gjEsDJJlW3spf843O
WJm48EfZKhKoeUH7f9EDgrc0SfEEmp/GycMl3H2oql+AWN0QAInSElVjVjbILspB
IlGJmTntTVDiwFdNg8QaBD3H6KGqKK5D0NmqRE7XjV/1h6KOuLzYihflhsYjGTBY
ZG9JE9Hr64s1smwL6kwiE1oyoD9HyF74/11BdrUuchzeunHoH5bGaEEzzte++QEd
Rbeb4MbEJH06NfHOEy6uRbPg8vuQ2hVIRAutBBuIF1vOfx3HdC7wJpvFl5iUei7J
5XH9XL/Xe7g6vvNPO8/5wp5Bayz+5+MQWU5yzBj6YkHo3kWhM+E7Ip3q36F+jl3N
EtTarNbvq6b7yERIJ+z8n9o9W7MnbOHzmz0Ho3hLHxvQ9O0SoR96Y6rhjUunnB7P
LriHCf2zrmMZkFuhI2lmPve55levYykkWMAro5E9sLoYB7XGdRsu6yf9HCw0xFjd
whlfAS/aG3kBJsMq506KXIgdx32xEKhdktUkcMG5dKeDjbKCO+9aZZP/EzfK3xVx
yqS00TR5F/apY4jQGxvX2J5CB95g/jNgaGODHg+dvnFRT5iOlq+gYN2AX6Ro1Qis
1i22z4nxfc/OGtw3hoVQwsdq0urjUmg9nRmH50ZBRtI8FhQDY2U9zOAFJ9BTLnli
VR+nmjtGmvcHX3m/Ii3gQBPx94Tpz5CjtOVAl9pPmVDyLq8zVQfpTZuDQRTxlH2m
mr0eV8Mmk1SpyPxtXzlpxW7ZlIicv7r1HZ6iwzgpgvXnNjyrxR+entTBGx9beHcn
ytSgzhWUWOCDnwBgbVZ1VLmaILQQDKbLTIyZTHHNBW4FAHXCk/HXuBkmDmeLJBOb
TTsm/mYz1m52YZpPPBeS7c7IbnJeqatJJ5DncZAWEiZKoKn7h4m2yWyCDYdmwVyw
JnFQULRqSRJaqKmLtEom5maT51SC4KdFFz0qcnxM13cuyzrw8N3qEr7e/4qwUU/T
YCBDZFSim5v6DMzF7pqaZPO+TJSZCw8DT5gwck0KVBO54ImK41IdTJNdI0s+JyHq
FzDWjT7Cpuhuj2b3qoVcJKndliAFpZKHwK5aLA9koCTwhm7fSmITSeTv/l4/HAJR
zEdM8DUwWupZjaasIjnJRNLAV47IdSSX/ZFq/hbNo/w9rMIRy4hqjGD4qD+rZcK0
F+Mr4o35bSHxYj3P9QiU9KkYFdmyDeZ2bqeFKrSSRlzq86M7bc4HyTu8e6/IZpFK
UsblnLpetn0GAMi4qL9tAL81PPSCidDugKqk97qwUU2k6ArnALV1tB1r+e4dW5gz
0/SVOXPughEmsL9crNq27mdpzxmL5S6aqI0GKskXQAddAJNfI5uhIp+IrviF9o7M
Dv1Djy4KxsCsmjl5iwJ1XMbuw8sxMPdlZ6D3vWNY6IPgBU5hjshaP4ztzRMtSGWq
0tIRHN8migazzeurMRZJp1c9uGjXV+xA9ZboLtqQ7tINwPkS7A0vs0O5fKaj0xyJ
OR9OHsa33tngIOfaYyUvdcSYrM7Lj3X6+JUCHE89GhIz5TT3Ivs8mNNlFBV8VED+
44SkwG7PSom04y9RLhgvrHAJxfZEI/cl4ixegb4drDS+k5V5E7H8UpK/vjy0/lxY
aEYcfZMF2OaGL2/kYTENDEshy1IBL6t3FdoOA2gOo0/MOpOYtRElyJzjewJeY+zU
4lEv+41jl0Fm9uqHuflD6ebqKykGOE6J0O3ymiXZ7u/VYNw+DNu9GxDMbqkMlMmk
e8Cai5ahZC2jJmc245I7YNPaPjRBw8/4NhQmVnzF171kzo/2DTdahpLKMn7AgbMl
Riyfa1bJS6vEMjRPWwiXweRLyhVtCR45zCwzavzHa5C79m2iWzCR2agBite4yAij
4wHOwWtCX4eiusdlCdJVxmYyqr3iNsQvMNgZ7iQgqWQce717sZbc8aESmTFb0PPc
d13UxN1sZfkIJQQx1Oc36vVbDvXKIRqqGNhPa8NVhgGadXh1NRrJAJ77Eg4yQM4P
LD3xdQsbMZW3vQW51NBXdjWnJy+RTJpJggQAOzMzxPpyoKH86MVapb7kMGrxfvc6
AqYfw1V5xwFsHybMsMkPwDFvvo+Zz5dFvceO/4CqA/Q/dHczQcWyIdOBMDj/BWNa
IiG+7PuXV/GlKhw6MqkEaB+xzRTn4eTLFOCtpnTLnic0tI195jCxjd1RbnuCUR0P
8O4vAHRleC4ZBWIgg2dDsri7hnYt3pHG7DjLv7FE+ANTEF+NZgB9O5ctRyKoUmWo
98SW26oov4gYzNaVyYpXonYBeOUHJ/q2U9ci+AzEPvK5XTOfWoigsk9bZfrRQcEu
ZhWcDzIlXwy6U6PVAsJyaVnVNgAqk02BPqxKBSd+ZtKpRawAgXlXkNAnKr3IOPqY
5TcY4sseKn2mTua7XP9DPuFmQJDz303RuPrDKqIvsAiZmN0Za+jSz2pXV2HjzszD
pSa+W81Zx6NpmqUThwuksVzd11EpXkDYLny8ly1PFDpMmzMjo0Zgy82x6PtwP6/Q
Jfhzava3TlqlA0ww7qRizXO+RX0c5kBtp4w3vvQwMh380EuPOneqAexbUg+37ueq
ptNAGP9aIY9XVdgf0DqqZwnrB5QjtvwC29rFWFUF7h1fZgX2QBRjefkC/8gBW+Jw
yhZiEeNyk7YbHetUzTSRZyyforBVZLCb/qrdpzHEq4cRl/aaKHkBBNeJVdasSicS
0dHgjEmof5ANjZ0jr69f8yWSGmgvEsEkQioWds1kDyctirEBruRgcMpDr7s8OOpb
pjnrqitg+Hag2U2xWML2NvLntvQbNni6bxnd91xK8zB7ZJ8z5phwEI/kifZI4ROk
>>>>>>> main
`protect end_protected