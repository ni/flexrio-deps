`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 50560 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
DBGZtUPdvgnvgIFp6VMrQayUS12cAbQy0qMlMffENAX3KVd1yeEZhJHRUoZf7NJx
rcJxWCiRxNjOEX5WZuphVckz0hITOgCNikjwGmaqoJRAdHugppNzxMKeNZ0KWt/3
PnhXerI3fuxuy6mZXPKrM2xIs2heb2SizRb3EfSrOSoX7HiJzcuanqywHtQCt9/p
ESxBfAi6jGoiR6kCQxRd7NBGbA9UqD11lbN+put0UvJJj5oO3BSpZObEE99Qvzif
JJe8PaJkFV0bhda1IdBHGvDNuYkI89fwVj1UeQli9x06b/pguR415e5uHvjl8z91
JqesOlSZNfKMlBYUWslzis7HPZ8p3Z02EI9URYV0p7TwUTH55z3G0gsug2rsiDst
+qqbbJ2+2+cnpblcpPyZ7+6dK0nbJZpeUdfKy6vcVMj6BE1j+Y+HP+PPAoshTgxB
o1fimxrteRTthvoK1noZEYUkje0oSAQKe2Cp7CeHNkF+uuDI3LuyrfFlam07YXdm
pWPCam7ZTJz/vy4I/3MhtioA321P6y3Fz3S6EsIpZ2dCn084xXEkuKchPQrYQBth
6w6WfjQKZYlefxLRtuFmUsKbF4YFpJEjSucDFYnRA9ujC3P7/7yJzZBQhBDq7SQ4
hFzADgu4K7KM2Qw0BAXQ9ggKpKU21qDnqGSp9h6Elwawy+VwEe02qDgsLMQFFjAu
mvMQnpjd/VkhGUiXA2AGPg0kmRgKtrPu6y8C1bi4ujJ4Wcdt2KBKLZcOt25qAG+x
C+c2yxJbt/U2JobHSc3Nl2Q43NYL11bNSmjX54IsM6DK/u6mvu3uF8m0t2CeDnkm
uwwMrOrbIgCNy3bo0l0BPmimtw/5hA6i++ycz+q9BVFv2upivSZdTf4XNyUg5sKI
2hZ+WCd+IBpVAVG27POXGY+/A5mbiuLV8gQLAjW5qakod5pg3KFXuijTI92n9AUc
XLtbqd0b2jFjAJv+li65KvWZi8Q1ns+4Z9gphTR5b3A4KB8Dcehvd9hCssMGUSPg
A1YfBywjN65qzPrmGeRRGR0kZ63iYTdJlsTzlJ4JCuAelfN4hvcGmksjHGcQcTbq
/apUU5Jb5jN8ghme+g0pvDBN1CPYM9vm3o1B4a4bctKcPGZAWu4mKMPFMyEcx4l+
5i0fePUj7tSPyzKYukZJeJe7ZjsJS8DYD4+F/Oznv2S0yehskCMN4dUgh/mpNuEd
eMrhzf4OhnzGtRVhMsnWi+XeeuDkGQOvT7/Hfc0zYEjsPuu/ftB4c0T+KQ13EV7A
fT90+/XkZ8khr+aXdomX80HmwPcDsAN/4my5P9aJynGlkXxI25zI1wrbOjLcW5Ef
pyTWYQUImsE9I5i2YmltK1IbfNF07/PKdc800jp/14CZ+hOb2tP/OErZx2DxFv2P
K1JJRqNHvurkJPtmQZh3nEom048CsDcu2zmMwN6ZTlRoaoNErVCStM6tBD/lny0h
GOKPfYq+GTTfm/RJEl5Hv0KsXK3AxPZLRLNoMWfQYj5yVtJjyTaaNAjMlrNfTLfh
Fu15j8AdibIQ7dPd6T8R7Dqz2Xyg0sS8V7hOhk+dgfXeGTpoK2WkpQutbsCSuiBP
J0ljevjpbsx7kQNumgAYqySy2JWKrc3I3Q/1rk/7B08HPTqtHvBXtdit+woa1T32
hhJaM/mib7bBGJEgSKx3yIfKr54K/4qHIVL5xYgWLHw+oPjcsTRL83LCBOjQjGi2
2ppH7yY8yfVBPs6jTa5RZ+DTqiFpPJZKuf9jOINh1BImK6usv28gtNXoGIwJYzNL
WArn6UOf1Qhqxlm1537t5Rt5hCLudut16VpEYPJuLWOSqRSpyHx+oyYiAesPGzmQ
19bN/ybX6R6B8PxiqArGUlwmufbUuSJRGxZGjM8iWHK9PmIWj8G3WIeiHXVbYgeB
FQJkzGAjMJlCrjO5Ob+Hu17VuMJR4OTklE82KAaQXGjGuZaDG8WgV9O6mnFEaVDi
EQWrnlOq5hFMylBaaSk9ZVTcxQaGfoIpveMxgxxIW9U5q/tw2XP+3zIlR3KITUpr
y77jyp4AsHOhKi16ZovaOuwnX+ET+b6X3WGlRBHVynvI4Bi9jyFrQRWcSMCyMMr2
/cAYUUxSV+VQCncj8xq3eWfb75MDGUILRnfyVAmsCF0sxBO8PWkWpIu4yx7W0ucP
mmjmyMMy0Fx2BDbdm2GWtOKsr6pOzfrle2oN/4TxuYItWLTPa+IIs//Kb/LjfOmQ
oJyfqKJ2GXQSym6THp9QnNuomq7t1UlX69YzRbx4a3y3vyIS0hkUGmKDScR0ia8B
TXDeTGtqIpJAkwfcLXfXv6I21sSF8e2tr4X03eJPKK5IrhOiNdSt/rnrLJrIuqY7
U9qB/o9YjT3jnSKPKgXAj74XYTeQMt2aug8q6GrmUrhxxYmkTegQ3+FY8uVYmIW3
1UiRKgjRmVRO6X5KAsbqWWZYrguV5EvBtNmvgGoP+TvQsZK9NAa+0Y0o6km2LaJD
KYhWyHNrmfmAia/1prLwINnoVkgOIKw8+wpccOHpsii92Qg1X17INBtjWD2nKwgI
dJ/2kU6xV7t78funhFWt2a/hUkfck8OUVrZq3FrmDQtcnE9JJjujXyYZzUDr7t1W
9+x44+TsoXOc/hsbmF5i/XUWs1ujdp01ngvhUAGgTmR2V5w4Ke1IVC53KOI4vQWQ
rarb6u8fowOZSwslbI8j6VLTxY/sm3M7HATYL0vDdFzYub+j8aF3r8j2YB5Kncs/
gin9eaEjSsZXaK7JRLte7nC6Efzig8vu/FrCjGZjCS/YpHMQYnDbdxpJSxMgl9Mw
1Dx/WyVwSMlSbRimFO7IlZUVFBz4Ok6uRW3sExipSPmpDEd5vsH4rtyUeBlKUTV2
j5y3fS544XJne5xFM7CRPOP3k9G4HoqaHnZSnO7XrleUfjRVtg8h0DTCGbuscd1c
sJrgTlWajJl2FLVmZCUv6inTA+ZzwCw76Js+LrSmpb96Cp/RR1oQjunO2Q0OgfMn
PBEl6TI5Z62fL+Ha+pGtT+LrliLNuC31Zzhwkh/z0YwS0WTIoQqEU5r7wsOcYYLg
6ZzxCJ5Ua3frxs0xi5VSWslKR/u+N8ux42+hKGH/5X69EEHfq0v7YqPy8mrk8ank
F8SQ5hAOPbDonzajafr5AqLLOYHFM+eTgmY9qwC/Eoe6uZWVhUE4CiM+VmFPje5c
r4pc3s0RhDEKR19+x8Qmhyv8CsxoisNexrfb8nD7OWqJyUUiGvdrHWdQCiTKKMPo
eEoJ6y4Cs5h9MJt+X4gtWjD41JKho1Usg2229cqt04UqzR520btpJVL84QkNKlN3
6chL/ARH7fwxwxAsGWsDVEoTOKdf+DleAMcQuRqINy7Ml8jGIc5TNAGenoQJIih5
+FVtYFfOHgiezBhiyy8SiWnSXcD2I1fu6bSw1pe2G9E9icQW/gW7M6HW+FIoONjh
r4fnP+wlYG1XxcKvx9wp4QaVFRcZYW5JAKIJ/D0bWxPIsR6uXTfV9rE60biT0dg5
q9pGr1T4loYdipnzx2RBlgm44xySTaW2ev/eOGqk5tJkCa4aC1xpwV9mT+MRqWQ0
0dCgIeGBzgocvfRpUQofCEM3/vAMVxIpWyCYuPfnXSLBLq++LfqUp0j7KtX6pXee
ZVT48F7w/04f1QoTHukO4+LvArVeAfNW4ASme0HTl87NPwxfvQnvLzFU0IX1mBec
Rk1XNetyEiCpP3v1JMlAlv5rin/XCYqAiBhQXF6m+OWFQypg5Q4i8ADIF3idRzXB
+Ci952aFvsBxo38yQJ3vR9A6AAud5w5TeLQhSZkgpNHAp468ZTblgUlk8xqJicta
jSUhPF44lVQ2Sgv4sGi2AHo/n+qpu4thDtYwusqxUyLsZhmrek4UAC+h8I3fKr4w
CuO7uTshMBSUIk3wGMpiPjVXyq3TOVWZNRo9FpYaEahHSXp/tD/Bgb3+MsVrUR3F
h0p0k4R2SP15lpeSW36+gz7pypc631fsl1MiTlNUN+vHX1tW9f4F5MQ8q7l/5YPV
H/psMq6r5M03/aVAYHWCYlZlVV1vqocbyJJ0ppha8akq/94Pp/vk1SfHSAbinh21
Du8kEvLE1Vf/qytYQcEcza1P+DBDs5V3o8ChFLxvtL6V97XEiNiWaxVce3GAXBtx
CHmLU+9d1BZk34Ug8T7giqNQF9lonuhXWO1dO+0JIqDxXoEUPPk2Zo+psM9gevUV
vB1FrXtNyWoPDTh9FC3uF0wF1YyDD4j6lt8KTTmmKY98OxwfVOA3SWHFDnWtUNmu
h2KIw1D8iRa3ipnRNErynYzyfUE3aCQBuQtcOMjNHpgFCChkAz8hq9HIhcmv/YX3
KhP1PR817LgCmfuyS+7dz2ctUxa1Y/ELQkHDZeHaxsYZQN5aUC8L1YREn51nFmUz
NH+LiHflVALC39w2qvwqHocsca0m9EknJqY3A17JNjq0DuIQ9g2xw9twUSsy+cmO
wZYK7PtPpLnBRA9GHIHVWbgQxqsvPUgW9eNMf3K0dsOAg3jMQeI36UQvnNnmMJOD
nAHmTbYHPbDvg9qh4mZk/0VV7G2MlqgmvTJd4Z6/eqB6B59ODPHNJmoupFJrFEsJ
WLZUyiSgLmTvfmb4aMSiRAaJNOsq294sxDnsuBrFYMDKtx/he+tbAUPw51ggTdC1
QmP3q9cOPN2k8a7ZVZsslBMOwKEKu90c7ZdWkTO1ZIA/ef/k3cpHUbWN+fphQ7bH
GmjMQhVEn0o8RYKR1Qq2r4KIebhszy/mgJBED9INLUPcIn0Sub65+U5N7XNNiGy7
9gTbX8E7hd1AUw4/Qve3nRszqRaN3QQ2i+tETnT1FTp/5QrPt02ahk2khNaQlWBK
bWD/jEq9GGq6Vzz5lcJis3GSSsKnUiqcdE02i2PblpR9y5AjDwW0Oh3o4oRg9lUA
fR0+IK6vMOc3k2Dl6sJ5Py2ixEeVn9bX4+2eznzU9r4bJ6tPJE15TFAIcwVckCh+
GhGJ/oTYC4463yZ6Z4FbtnP9ZK6CRAm7tApMjtglQ/j+szJDpdPm26do4BJdw6zc
ud20bIDTfVopAuADZSE8k3o/uVyF+WNWm3duO4z3EYF6Vlrj0Ao/M6vAFaduUtrw
fUm8HyF11v7lyLSuSfJBReBu+rqZXY6KLvK2pzu427FsbAf6iGsEYAN3xU9bZm8o
ZsOM2G2cbN1M+J2mWjlL06Tfb0b970sl9BTSll7CArlWEB4RUbupsses+sXv8eJX
DqQjcXrCHKKz/e+PrYIaC9uwj4m+KBScxaUQ1wtFP2h17KXkpPxyKNHSEG1GFvkE
ty9auV2IZorDxlrIyA1jLSbz0JECh9g1F29tcy/L4UjBzylEwN4eFQJ2CO7koDZZ
Np7writuF/O51NDgTWTBzIw3j9TiiyVkack2jfbNRPOt0hRKLMh1sS5FlydLUBbP
L9/DvvpFYhT/Qk+lNPiQD8+mxbQpG3jJQive/gHyzkzIAhRXVQLLAeX8stMTR8WE
ptZlv4j6UE9tVRPM0mQ0QNunXHH5d0Yp6KUh0h3lmyy1Bxpd6t4pAJrbi6n/aaIz
fhsipS1DITgcfiSd+yIFgSeKrc8x3EaXMNgUcTVw+K9r8cj+mUyLRHG7HrvkpJgc
byr9U+lVt0wjpmWSc1EtZkc9Czd25Z/etAi29rYb3TpAvRFpOSazq3PM5zV6PwN4
3TSD8Hrd9a4zyCukTv/ANNO9mHgcoHyPAePi06vp1WcDZEmAB7ODLLwSz0wqnGdP
ZuxOUixTFzGWOplJn5LBMHJ424RLs2TongfuBwiumrrNDkMMDRf4+3QP7BKHZL2E
47ebkXxVf6xXez4gj7bLCKftHNHALqCrGIYJlXrwrz0L1Z9v2ZsorGCA1t2czOa+
UXhDK289RUSh9TWvFS/PpQTy0S0WOdadJdBSCOp4i/WTPMnUe7zXGot1hE4qhIQy
Zn4nCv5G84AbnT2bqRhLTWHLXjOD5yExUbu9SRKh//SnjXC4yvvOM1avz454A+h9
T/RqYcuY9vCo4x71IKaf1mp3UiTXFuJ8ZNb8t+A5S/X9uJtYRj9GSz/Br8aFNrkK
g81kyN9TLP3mX1p8cFCP5lSCnGsl6V20zHRVgsufoJ7CoSQIXuTVTC3unwo+cyJf
MaUkOsY3JL57XY2K/gpiTnnfIdzYe5BzFRwBzussG0OtvAdt0BW4oGdWXKqBJlJ3
L4K3+4gcMMKB3i4N/iuwjqG4+Cau1QoKLk3WFxvMM7HfMbqdgE/YHc/pKr+0GNel
Enrovy8j/12s4dnr0gp0uhTLxdZGjKqZMxCLpeewAAiW8mvXnwmDo3cMSAePSdQo
C12y0EJs/XhTaBO2Bns0HM8dNmtvmF9ifK2DMOn0xuvgEklSrbO4fYBciJxSG+jL
G9zX5iBL83DQtYoNGagXk6JL6YPVQCHCxEzcq5gbu1/u4HadS97FpMS9gufPRfoB
zfSo1osI1jOP62kEtVm2zsFG2RLJXu99R7JKUUpqMb3iUlw5fiUyOmjLrlIo/8dM
ZlwYO2dx0kJw1cyGEaZWiTjcegTkn2bRsJtV/0CVzahhkNk72akhEX3YHi53dlED
P7kAOTu8kAxMiLnW4ngE5DI27lUdDPSHuYhKt3QApkVbbfY30kRRd6ouTaaB2ZHT
EsRychlMhvf0+jH7ys+IDDH1F3xHJHg2KfLIism7ix4p2fuar2y1n7xB6Xfna4S2
c1495RWTHTe+WXFOYF5LIPUUQY+xtiw44qsmfz7KxcJ3zUGsLVOvfcyfJDJVCg6C
VBafPDz3NwIsguRqyi2sKaXRXZN0ENGGSY8ShASXtoUaBMqQ9Lj/Zghw6FMdIkw2
CyENFZzeNNC0vCt/XV2mt8vnnjN9WksQZcWxJNPZMXAjVvUbLDxpyK57B28uW4W3
m951+xpDEGbjUcqOY5UOEMVkbPqcqcSxCivHx7ejR/3gMDW34ToQBlD7HET9U8PW
q6D0SasOn51YAGqgvkBiRj8hxiShUVebTJNvQzhVbk+CrEJ88fUKKJlfq9xUFSKU
LNSYaUEXmJCZn6Gf0t1TsuOtXdUbKkjdJJ0uJVZweDON35sYfQY6zm+/qLkaeamy
ovCBIPDk4uQ8XCWcmJokBRdUQkRhVnSpSkbvwN0MNhut8r5zhcWrrFveC+BP7Ux/
G2jScOi3lsf26yFfXZLxakg8JOdwedMOqzJwnLcaEVqgRsb0+qdd3YOdS5PTQSU3
J4ccblSKlgI8BMbxhGizMgmxZexyYb1yaY0DMRYPPmOmqsm4DSzt/w3VRbXC4mqI
OJaDybMpwyv0pXbckdyvCTmw0WyztsA+WvGjf3gVcMUqZYCrQ6pEliLAvm0Qt9g8
uiscFxMBuFPO4qPPCDJoWSUGh2fIGoiwagZsCC8G6QCABp0cq4Zf4J8AWxBlD2/i
RouNSKhLdlQGOjvy2pGxY4UV0riUnFSMDshA0yExzHqgUti6t/aW5kO2e6fjOsIC
jEzAFzlARSxBv7tvYp+6gRjE6+szD5eH+x55L2kx4LeQCtwTws1x88o/RYy0gqT7
7oWGvRFrbMFZd1g8Ewawxb0dI8/XcNu/1u3wBeKZdO6w+RoYWS5PuUt1MJxS2rMk
ROApAcnM/SeF3TUtoSetHU7IJ2ADyKz65Ixs0TP8EsGFMVy5IeNuSG9pvU1vL20d
K2RrWzrxR2Letfa9uzXG1ytHxb848BxyUnf2iYSXIbfGZBT3ifGawB6y9rJG5vCl
krfOon8UgXewTGeoY/Zs1Jo5lPjv8jWWEGoK+SvkGeXxDpBO2yrgYmkYoZ1NUb2w
oJ4Jj86UzLsBT/T2+VFj+MnwP5tGfEudyxKezU+9eFJos+5qGfdEkkycFsXlK/wX
y3E6++bRCRWwtcQ3s0cExQplH960zLEtvnojeGHN6+6YDsk3ru+L/dkjyH0mOHQm
kCOWv6NVfaLzYoiXOe36HkhVZkejyaVMkgzW3Ey8/F1HKrK7yfL0TtYfRyRpt+T6
eF49XIqHD0BlKrqleQDyMnO246n5i4YV8JZwlSzqW4FmEZsgqPR0+o4UG4LoYV47
vRcPS0buw29QymPaEY+72Zmyb2YtZ/e50x5xzukZsQ1412l4lw2NpyTLNUjCHluY
RlWk4sAscFaY/htin7UZ9CZEEhuY6ntNJQBqzU0zDJbrcbDCm4HTnCPIWzAji0Dd
tHww+ve5+TIb0J5FtIxoQ+zq3Qor9UCNNikmsvzjXY+fSrwuQKtf5s1LFqkTDkTy
kvmy6PEJx90KO3w8NwqBNrBeLJ9CXD4AOwgY+n4GsXJPb5PKg10+JRKuVUTVd/J3
gzNbdntW91dky3+CtArp+WJN4ayM9YXnjeVfBd79t6tMuCmlnAdhMams+Yfc+Znq
0Rq9TLeValHG52eJVz7EMCVSzSkLUjXydTOdkT/F+gOEEJPpowpto/EtUc9VlNBb
YAHZ2AqKSI2QE/ELuN1CaOODp+Kvlc2SACzD4a30ZcE9hBqgCYBGtMIUuSnzFBp0
emP3Indq4rjw9T/+LqvnvfJnGIOcXZ50tCs2xqEg3zaWjk7qjHes74rOvhANh7ca
vPAozzy/dkbF6TpKMRvDWOG46zfaf21CQJGhr9S6BG575tYnMj5DamMew7cEGFg1
9dFDTTZzAHvJwjB7RocI9ns0Qri0IaUXpmH7KlotgeKYZz4SgDKGd6z5c2ZAxd9q
SC/7VwbTHzCdbE1Gy67AhILxNPnw9XZRa+nmdVxfz0xeLTgSclPfGRJwnrIGx7Vu
2MNt2NfDyF0217C17aA+EsZ79D3K3dGuMTrItqV9UV8uny8ZublcN6yGhb9x6rmB
M8anGjDuIzV7rmwXK6Bcgn4gRAosyshpGaIA5ahWKPljPVXuv7YMeWtmt6cI7sBN
zCQEYGqKMJUvVf+p22wxgqvCiql79cu4ZPaMR+OJN8hRCU8TRud+3kuEmvtSjG5k
Bk0OpNxRrs4F2nywPgfId/O2qX91P9zFW9mAiGXoS5yM2T7P4v5Z1g4uzWEddHy2
wDiGpcv4iobpZ2TV0Uu6ZpARtXjf/9EvjWNm5I1yOi5Z074BCnfYdBhzrOUkMFL0
Ias5rk3u0QCkQ8f59iiw3wuizQEGdgG3qwJ0T34QDrWbs+MV+JgMoUl4b5TGOquN
DmF2JizlA/uhIaUM5ydAL3guQ2x/xD9/ikrVNJj+JBc0b8ELCac3Th+zIvOR80Lg
fMA3QbY30mh7Iir8JeJy7wtIxDn+eI2wS7UjgrzwHGfvMUwHuylZNcnJ48mtpxkO
BCslx27qJW0XmhTFkJaDjob6mVr3gsoJH+vgZME6pHxrt+FvYkIoULZNkaktGF5s
TT36/9uKoFJ8Xw17CFtOcjSYuCfeyBSfkBNOANqWRuf4j5CzCI3BwW4OdjKInYeK
kptnMZb6eYJT6+Is/hH/J8MvWco3ZDzdQdvNHRZV26TOQVZUW+Zz9LRclteEq9Cq
YpA9T/T+daP8fkbXsWuBR5xvED+pkZ4GuUijQZrF+KymIVQ3OH7zZwgbLFSLviKt
35DDUcHYut7ON6PJQWLJmPRdoQ6NBCpvrB+fypOh3csCjnDiaalGaTpI9HOTXFaO
/8947nejDSRkr6UPq7blHTIBGvtjuqFPSLSafVZYcswbrk7vD1PxAwEDC39I0KtG
Vjnv+thr5tO0z/dw7DCs1fazFi6bk2SRdIuP5S1g+Ag9JrH7pmFdjk8vxSGPLR8Y
FHn2dtFC4jW8WRwdT4ieQa8XYR9Kvn+UvwH13R96qywDSj6HhyCz/d9lXP4O+saE
/yEwURiJuAWQbbnPt2FicXbHcBxJbIMotZ/BuUn/kD4/X136+/CtW9Go0du0dbpZ
Ld2xNHpZSnZug1WDp08ZxXumzfII734dKWNhbr/1ox1DX37zOPgawBYvmJajO5Rf
+68HOpjlMeHooOI7TY1O1BQT+PuDLF4DOAvjKKVICiTzKRq+cW1wypv9s0kMCkVh
xXVykCRovMWMOkujG3cwoTo4xG0j4TM7BhOHFzk2YPIg2iQp8bG9SnLmxwTLjRkx
CM+8YXbQhpttyNVNXlfv+PSPtBtTyYjUAoI+NWyyp5zrcCoksyrfgL74a+6DKiaF
KqQaXvDU+39OgeJGuVOsUQvI/qEdj0YvqJXvPAE7yvnp7oo6zp3JpxEcuBrU3Z2N
D6gQrytEh/oGTpGMWqQoZCRFQnq7NI+9iUTn9UjMfkzX28rV9ss0pyYlmW3y6ic3
AmvVU2GXBfTtmfL3NXVlfduQcLW2UcSQ9bewaB8uPA9+crwic6fq3cjF5l58bmWT
94UOcVsWx3tnstFdeUS/0oiEQ2ok0vGuDcrRYvx0I0rBzD7ZFgBErRYpMk67QAfN
y/Vnq2f+hWT0iPEegir5fdZtnfdXxaVfaullTFp9qWTibmDL3+IIeA8XtJSqu86K
6bA529JQ1DY3hPtGWlMZbLY6JDSFiOdJaZf2+qcM9FazAYl4mwdeDwAIUcBw91a+
t9AB/RXykWGVk1eKBLdOd0QNC5RTdD7MpoxIHFHwnK0YTgGbHII/Wg0XGJye0eVg
GeI4zNr63CKdKpUivU/shFJ/kJBZLGtfxnVcMQ1ygxLVynxmuz5uQze7EYxfowfw
WdCx/Yh8EMLTYb2Qz8zEFeoBPQ3hMQhNn0Kw8ULFRr1o+dWBBwK1I5DffDzrZiVp
GY0nu6tKkBlA1z+rwtgoHdfOJ9LRvpA3KUccij/g2CiI6tRXYMtLoNb0zhmr/gg0
TfZMCIQFisQ/fz2yLwDUsOEWWwnLJ+9OeLkxj4g5K6TpoAj2cOoN1IQCIttt4hEa
qzr2JR9TUCIO/7kjr3tc388Smalihd4ci975z+A6eIVMpMyzq7/XRdTZFIPRi2v0
Xi5NRfQYPmZsNGN/KGpBURxddE/eLxJ+UaxamdGkXdcxZ1oOzYwzxaIIvB4U7UL3
fCR2a7zXs8fNKE9YFWxeVT73S/qajzYUoyCyguI17F4nBVujlL390V3YM4jMSc+6
ThnRmmI/YH+BsFhEBLBXVvpU61anx0Gr86cZm+G0d5x2Ui1DChm+WsqrzA5IO1JE
l/g4li2IwSHsX+TtrOGxltBZHZZOcDbJ0ShoHsr5Y1cNyWZQEMticRz+th3q+o/T
UGxQ18KBNIXNgesL+e7+aRQvNduIFiHUxTaM4nexXSn+vfaEwM5D/p9amhletgpw
/kdxcjeZlauwj1K3HyWhOzc4XYp8l2Rrjneg+zv9Q41GrpDh/GwYsW1f4DjIslJ5
Nnjw57sCfkM7HMR+nmtqjUapMawRItSGDiTOeTby6SdZFx04DzYEv50/TDf1jA1c
LirZce/YPUOLeyFTSx27lLY7NDdzlUJAp/e8KvINc9zDTXRJTnX2Yb6UNgDks388
1CK5UhmV7qVcA++AcFU6A0FFHVXp+PxjQZGq7wbNdhT5xdhuNM8b1VYLywBXs+3H
y976fhgk4GuVzAjd6mbM35kygIfsiro4pTOxGYSkZFu0WcFA77wkxFWyAmfzgiQ1
g2D/2XI55JcLI34cqOD7mLE7s8MM+CikqqkhUy36RGtn0hI6MRe+p7Atlikn4CD+
iP+mqNOvXSos+4s6Oq8SMVcU7nvluU1+Cg+91AbcMfjSaEF8Z6K0p/TE1kCntlxo
zo77nQB5EXR3QxaolxRFSxHQ+rSk0M9HQVVvPD7vLYxB8G798loGIEWzeT8AHWub
hudj/mn7DQX60EMXAUQAyc+ReXYnqDkDiz8gC53qdEljpIbBB+mZqKjSOrXvFRYQ
t3T1269sY3drhfooN90lbiKDJjlCYHDpXFOSrJWkn5OM1M00uFAyH3v5ppuRLE5y
lzRdrET8VILwDmZOfvX+0LDajk8V1QV8dtbO61XQXvgi4kCU/BVfg0wKwimeiEW/
uOWUa7zi2iIebxO5RFr7Lc5HytVpBq5tcOwTx0c/0JUWSiCy9eWM5Xv4BCy74aGO
YykWAH7WCbcGpYqH9sczX57U3cWKfCo2fxZsUqNm8gtsiuwNhDgP1Cfq+cQgWfi5
E5xNEJVfxH/AEVRYpHQJK91Qda30mbIFL7IlybDGwe2Bb2BYUNI49nn0QsSiLWxr
DPYqPNto48HbMwaeDB+KhkEE6ihvuhoqIppe9FrexSPAIeQ6cifkO5uWq6hdMmEf
/wEXXN4H1etJAaUK0t5qdf2JUVEgShEba13X4j88hpmmPmFiDWUuipp96rotb+bh
ciiGaokB+0bAydHPnAm4+M+IZ7dcf1obffyuMutLP/RUR/2V3R7ok++o3Qy+XMWU
VUkq0EQ6KScTAQzeo4HxDGlc0hvO5Yzibei6B0n8EWcvU8unG93I1B7vSeail/n5
Laz/c0xLaN2Dp8UIiFZeWlwv0Bey5xc5RRVMwOe0Z+FmUWSPmpehnDbMEcbT9+qY
3Oaqr6HOidmHwLp5VGnbGFV6ShP7S5EDc/ubf1WxJYawqPs7VWEpAc3a4Fkzx5h/
YTJqu3Xf38Aeqe0evfL5qJHXE3Whp7rXktUajocfDCZcpWgucq7+gmTim9h3JHty
D5Uh9O3zikAgXsiLG02zGqBAMFrIOwSHzTUC/1em1sy1zQNHU76FLW57FI8xlEHX
gSC1gjhPnY+aw/qBwAuNF6LVPu1zZP9DMht9MDuAYUK3nfjP2gIgdtfXeRBkCYoz
PlmKT+v/jULWy3aidrfQVidX8XJSEjjIUvXRxOS19XPqdkYyOi/FsPdzewpmxluw
fKRfABAbvBJRACeRz01UOdvj56ERMSihflVE6B32EQfsPNu/9OPSpoWh8UsBNR2U
q/xZzKsnwmPUb7f8voRlJWfHQpVFE5mfzpXA/0C9ZU1Eo39fhZE0zoXTsrmX3Qdc
2caJAHF70ArzsuXJ5eHlyWsAnTP0+fS0Ncz2S5iyo3qHRmkl3CruiokrlaH3nAoo
HyujzDDehvLG4CpuezRW1pP5bxq1Zn6pjTHQrDxKg9yqjHs1Cep2adf69SxMPoJ1
uxExqvr3SBFxAosnOpZCao44XU/fx1V+FpnGa0y6VJjBs9Y4bl26KkddWW448bYa
W5uCmppwgkSjnyaiQsY81PAcxLxgTIogPVdiqQ5QcrZPIvO/duOI1gqtn/eieogR
sJxqngxudauKwnFuz9xBzdM1WGIMFMcMsew1d43ljF0wn51rWC6oO95l2p8XoMUs
EQK5ptxEODbJBBnETCkQl5U9l+JXUvvu7j2qizLCGXCvdhEnA1DW6LF/zJKA8wDq
fQX2FnwnEpOSGUx1blmyYK/Axz6mlkVLs/TA0uSL96q2a/T8WPdNNonEwszs5u4b
bGByjAN2ZrsAuZMpUdG/96uef1+zPGZyTGoV77U4gLAY4UP/TfpwQxR2ScEehMPD
mAgUE2Iqranprxkq+v7MxFfzJnJKULe7m0j/JWl3duRXc5QQJuyO7gRz1/XrExje
rn4BTRjbnuHG/MFUEtXRCc0ozit1sEngMFLNvEpkOwa/WhT6rzqZ17zmvNxDW+31
lcEzsCXIG1aPnFkiaYKdepftrjKtJIN7J+CxSk0ABz0FbhNztBxakyS+8bTz7eiS
N1rkBzP10kJv+EACXPFxvOMv7PhhEkgERDK9NgcDT4wJX9DhZfowIClpEix2Y5U4
44gdDdVUBWRSH2u45xyBmmhiVtyfAT91j8fMaiwUd0eHCMjchh/7QHG4A37sSHwQ
59vyUzIfmzcR70sTtg6nlW/JNhkif3O4VrNVC3puPRvMiT5K6YI7CRIJFY+i8mio
pUv7IuT9m0/2SHgMyv+uLBDYzs2gjIzAZ0WlT/XTwBy8X9qkdP7um5m6aQpmrd5o
AFItlTy+/GcaeZVtXjIWA2MiTRkxWmzqDjiMUxM4unuciK4KO8OPuvfxqpXLjZcz
XmvsVsVXfel3P4r5JS4I+XgNwnKaCegbUt1SDkRMVtn2xcBTqQTpBFvxMlc5GB//
iKYX/p4cwz6tDNoZsxEMtfJxdhUR54O8tBodhq9/WQv9NGouTmVIV5qpYUQuScKn
S3ccxWWGNgLUo+iB8Mg0a93KndV5uEfSac7JhGsF1VvZW0hYnEFDqBT5JaiuUJvg
ir2QcJ35gQ/I9grk7V9GcJs+B8FWgIcFS07uSk9xc5guv8uSVa7IlgmhlLtifQSh
rtV2nY3okQ97z0IarE4v13CsrxUeAK/aqzYffA5xi0TUCRpWqKQmA/6aMyFz0ctp
GBj2xUkXB/ahnEiJfY49NjifWyLzPcCQLJL7aRHn+3WqjnME7Af1tzYv9UB9ui/g
06oY+VvMOU95Dq5gX+joog4OntpI/jFZZl4b++YoPL8SC6RJkOkTdx8Sie3+Az6g
A9oLEqiQ+UznCLthzRNne5Qa+gkAlmoUcoPpZQs53akRWVlrF1P/Oepa76/Lz6Ec
XRHwzl4qJeWj0o+H8jk/3gkrmX9QXvmmX/IThaoZk7nHMq5+vCNPvmL8uU/TrWwt
KUIrZ8q17lMcOrRbIMogLkWMhOK31NM+QKA5mRfQckKsJSSEZtdvtfGn0cMCrk7W
gMuLiOAp4tGGZzG15szZsd0+z1rjZ2sGsQYJnbRS5+fbLGZDlcz4psNeOnrYleFw
NjIkkzB/OlvfUEMpPDh1VxXSwNG+UsOdFqIS3gRDGr6yxkI4JQi9AXlyTWPlfB1o
iFe322L52PX2IXr+pfVQNvOgK4eBRzrOsIGJF5AIOOFUh5G+z40LvoIMqT/+EJCs
NIgYTGH5Cmu4u+RL5D5r9V61KRG986qg+AvWrfN1vf0Al5xQc6thrl5xgDBjoFWl
WQrkFlj8n6Fse1meFt7NGLBWdNmbgSkMCiAY4Y6l5pgvHWAG6WlKJOMWvUbOsLgR
2qijlBijtKKlfWPu8kWHw/25M5oEiSoFkAcWm6yvcjxkoBhTngB903d2EMhxz3zW
dnhjpAEP4lDskzH1Zs8xtS6uCR9A90P/Q7G0eyfVnhyQ0Q4vz4MZsVL/CfOjmn++
E9nQkHO3C9WB+0hnu3voVieiXjnWpsdup+byOzmlKiRj4BZ6tIr7Pn8h9/roqBXE
frcEyF3EdALOTYqjtb/zJDZ/IpoynSl0DTubZncGhVYW6v0aQgUzdb0ak6os5O+N
VgxTHLGrqYOkAsUUtLTsuxhB2KXr0n709O9k0HEIHOIk88wMmYO5e2QkN6e7AIfX
aw3TlCP/fSJUxGjnjdF6pRC6nqaQju/Kc2hnyUtMEVA5DLmWwCJs+f4tFqFRl1/1
QeapPlpJ+u1ILX8q3HqtTemyLUs9dlTPmth0yO3yKWMXVUvFSrq8YQ5sm10wmHDY
SiaKJVAg6gJXpXLb+Kl55togUoVP9mguA9UdjC3fO5EURwrLAid3WN1glPKbGwRH
c5yVaiq65+ZZUPsj+1ulX0Uy04i6nlV4tBUqNSRiQmiFC2kOMI7RiBChskCye2O/
NKbkgfZeDxJEFXA+oIMftP8Q+u+n8oiGyItxJRB7k6QxV6oWRYiUZFNlNdzAgyMJ
R1dk1KCdS/UT9bsPsMNZTRxrWbwiUY73vs1f1uHLzRqQfJuHRLA/IW9Nk76KBIzU
9TLopylS6bl+PiC9QijAjf0gLzbriBpm+7ezP+TGD9xA+MbD7fDaiEuROq0hh7Ma
5YHNPws1HKE1besxZK+TDzl+PYeDeB7ECuMs8XlxGpj8FaUjDegttOSRR8A+tY6h
QSmtW1UIyMS/N1IYzNvBFruGPpMENxmyPUzctIeQZ3Ww4tTuqwO29kCMKVduZ1Ol
B6+nNQ7TYR7O8EDsGHP3Ct4fruDsO+LgpnIV5huxpha+aWHvEUbv+gbUEK1S8a5s
ccED8WIDzDxPucq46l+pAPfwrdUhmZtiSAY3bNJBth5B4tm4u/gGKDc+FAQ4t7kK
QSF2GGuFwffmVllMacVVkJG+2joIUp63hEZLwCtkJI0UzK2G8XfJSGqENNujfLW1
G8GVaax6EWQRQvqsNO0m04K2CKvdzHPzLpmwT3yMjYOTs3idyonmJPooIuDYZvk+
voBXHr6ldf5csm9aC8HH+10JqHj+c8k05YnUdZ2eiTLnIwFwIlr/BzK84wGDMEJA
1PN1Q4tk1atsRWGiQCZ8b8tirda0tL1zDss7bAt3wOHOAZVM7witTAb2H1IfjPh3
YMKCAp5LFjjuKjEC1ud6rAN0qzI9hLMaoKnqOVLa/4u8cv3W9HUV92qp11g7JVQ8
zZ27lHrd1KbcpOQoDbeFkbRN6vEnnJBIGITKZmIpE4cz+YlxlbIkVIyleUm4v1pg
IJU6NgEtr0ZaTaQjcbDOIov4v6JI7zhEK+g/VSI3jsiyHl0Rz9iUN8G7BeEtiYi4
fTID4zCeW7N8j/Fq//HZ3jpmcBrHHIhJIphzUOGKmj96MP/HOAVd9pmPR7uWeVqS
IJ2i69B37IyOhP3JwU8ef2rr+Htph9TbzmP48lsY4zKtrEcTWRLI3eZWMqHmNDim
6rv4hKndi2NBUAC3F5wxmz5n1vDUe+0x3oBj//OuANzbn2R/MCDwv6eiDxMwmf7s
/3e7Lvqp5o/19kRIwwQ5t7cbxQi2xnzH5LfcOxqQz3m+rz8EFheBw4cxYH0xXh3r
0UK1iP53JVVfZ7jZgKXJ8yfr/aZOR8FQjc7Sf6UUNQKCm+5bhCX/35PRIzr9BJki
EUxEfDodyQ2w7pv0SDig9kr4u8kMhrSYgG3Q60uFraxQYG7a9LGB/t8qwIt/DvP5
r45TAN9YxVwZ1jpEo8cHYQtbXZMqtTLavwnD0sgb7/whJd85ElU09yLQFcLDYgxV
yYw/OVU45T44jhTb3zY5hgie89sTdRQA3EEC3IUpQ56GP4J1I/ud93CJONM0+Hhh
cvKd33n79hidENNwCb8sAN6nSoKzGpJ57CtesF+H+gV7NOQi7dLbZo66Ai1KIJKc
7Epr+D4I2wOJ8TVikeF6b8lKhGYwy2mv12XTTWnROd1TfLwZY+l3igyrzWdnWWpG
raGGAMOvFGjSl3CKeFId/BggcagkWES8IwIbkRk92vi12vi5xh4fSFAdmdEMM6+6
DOpDWISEGMGRbasvK52W0MBGMb/0r9icbAU3erQnbH9Wt5hLcf/zYRwEkMbcD+Kc
SWE7+f2fOGEmAYvvdlapSh7McYIn7bGcsVw/8pRiVmNl9jQmrbIpoR5IBk7SqyxK
kRY5+3n+WYy/32rVH4paKdMdCHMmASCFM30IPETDuMjPhttS7HcNO8UIq0A8BPBy
AVNOYq53307zA0HawZ2w0ijcSVD9hMRKasNh2v9T1hEeyS9TAG/OXLudfz1L5lBS
fsCGgH9Fg4oJ58AHp2pyP7SuwPWRTc6wcKptCAfAOwcbGxJlgysfOzTWq/d6qEwj
72wVRPePpjMTgf3qoG/cNPpKytMAVXGSaJ711ndSdew/DvUuq0EpESQwzDq60Hlo
JYqAq9Obj5Dt/MjKzmmp4v8Htiq6t6RuT/U7pkr/coKKzVwCCR5DRMflWui0Csl3
nWJkVZoiF1l7716e4gAoQ/h/pU2k5xIx4W6Khf79s6gH/AbRX7THQhxXlmX/IhiQ
WM5HwsSKrAOxDj1kKT0n8yjmIXmoonJkyuXVVA5YeTzQSfJByqCwHMbHM41oYRRX
9pZEnzk3uwfD4I8e6P20qmluSQPVdiwGpOcexU6ih5B6a0K+R6bb/0i5Y7NkAfrj
7D3fy0oBh/Ii8HcyyRgJVsuybOhperDMQdqi14Qtke17DFgM4z4PgT3/iNo4uECp
OZHMTxcR7ZAoSXlHMnNQUfy90cKnINFtixBoXvRwiN6V8QV9O8b7QyOF7d9WFPTE
RDHhcNw1rZIvDvSUHhNH6PHWQEYsGCZQLuMuIlGfeDjWE+QMfqNAUw3Qn6rtrfjt
Efaxa+7HS1b0Ga46gSLO5t/zEHtuBF2sbs/WaXDA/71qEMePTT0XXacBKTQ0sMVW
is1rd1y1zuXi0Z+PZZ+uUQpqtSq7Bsyg33VjAq0NqeXzYBJWRUTNlPe6BrPmlu5s
ix5hfT9QZIZtD5iFMPXSaWCeNVbNe7ON12QWGI8FAzavMpVqzuG7th2XRam3u5AT
KUINuYD3miYQmGDTImiU1+5WhSUpNnXhQaSKVuGhtzToiD7UPd6FzJbBP/DSLghP
FCBel12ENE32WxewkqPHH3O3RXjJqwzMUOwhC0cpPCgwDWAQw2U86XxnmkmzMRz7
LI+lJ8xc04qrZWxGkOXvHUTnXwr9AcVM06oNZUCdsv+i7DvcspLFjzmcMfZ1r5dZ
1A6f3nzJeR8E6toMvXPJBCrucwZ+JHYgARyaU6A7+u8p3po7ox4f6Ov2EyHoyfj+
9h3O4M/RR+QgeN1T3nXzUBxyuSt0AirbuK2ZDKhiI/0MRamEITHOYL2yfoIIMNPe
1XNmiJ3xziq5WeZTusWemMlK4oR5a421QtA4uDk+6J+PZhDDUSNBBmA4j9nvQH+u
SEIl0U63OGJiM9nHWagTckhVoKrN9Vs68I+UZcMZfJBJLIj/znwBy9vFCVjoXsEu
64te3AA407hyz3MikIrkHt6bqYI1rAnZVS6XqFjIPFC/ZsCGjYuZcLjCgXri/gyT
gJW426bfFW00TUUCKAu40HNdy3wJHIJmTmtm8kRUGGQoOwOo92XPaOe2xOqmmCai
2cMJ25Jf3sx399rwjH9Ls6cauSgJabgjXkXpmHNzrtdJBHcAC6PXprXpFCu2Jwng
BCE1Gq+fWlfZFCR3N9i0rqs6H7uffTzzJ7Krwph7HL75ovUdSs4jkmZwHVi6I5Zh
J+hs5kb1S5P5uweIMn2ZXfaPFBqXRpEEuYOE6civtQttQwpNUHvU2pslaZzhRQSF
+mtabN7osBfnhGOpMPLn0fHBjOTf2jhpSzE6d6/An898BXmEtwrR+VZ1IyjxNQMr
pvliLNGb7u91uw3XctZHTm0aP9o3FzulcBwk+inx80lr9bQechsjtyCM+nr81SCW
4CkSukDul5xZGIKT/uMprxwNNRa5Yb35aOgP4S7XfxM1j9mRUG7ym/G18XpzAyCq
5kSs5qZzjU9tDC6X2l0tcyR+v9YCkA8QcSh1IdEL7sQ9lEps/T+WeO8C6b9lBfbT
18tM+O8oGxcrcFPiCfdLXnoiX4SNpiOqq2wqb44tkhDkfw/LAUBjK3k0XzNFR0Ks
9WW3FrioiOxhvto8t8P+M8RbampUeGCHDoT9ZBbV2vIOd5tMZX/IgJ3FRv0q4wY7
zTol9vRrr3lHINIrPhB2jctMz4YGNRMB1xBwYShSKGeRjsn4sKpkMIGY2fP29Wa5
bmrm8h+xG7K4Z+8E8Mv4qNPxr4mtW0675opKlNrsVAwyVNEvMvl/hmhtsTMxMeP3
m3cjgryPYW9owbpFMKv4l6rkBfziHVy/5qyzp0Dh5WlIssxQn4M0I99PLKgGhwyw
jx91v/6qWgdXihxEU+uubSvnRwa/N2Hf/x282K7l96AxS2lhFOBfSDNfDLqz1VT6
qg06v8pcRMHngVVx4UNyBpxefVRQPDuuoCoFg1xq5dBIBn/22EoV888isKfjdy3c
ld4lUXHJaRWQyPMo7skPb5stQsQCymL6j2FjLMy8ErkCSCYCH2h80soT86n9uZIe
a6HX85bNltUIK3L6E64dT7d0Y8Dj3IiXmvYBwmrObq/OtgUvSV0yH4TZRpcDvLjY
RRjt3o81ReIEWwuFaJzKms2uk3YfIZK4NBcoaM4KMt6sik7PX2UbnyFcq2MZ6KVN
eFBNpP4MYMfadyIul6gApOC/082pLLK+3/XqqH9JVXew38GTrwdkkKFAS4puOQXA
S2QNBrOLhBENytQOe4Xo98IEB3GqyDfZjtvSmvbANdhgDjX4X2r3vbnAqFehpEr9
oKAsTE3m79bazaRk6Z1iFLjxKXoRueA5JxTZEuOxRC5IrN/3xoc3BcyaW9u6Sm2J
hQmj2uYWrCbvYKcHVK8gpAOBw0h6LMtgGdCdYu1EvqFAXQLLNHPaXBaaI5iXxAq8
edtUJ0CXVtk+TsF6Wl14KFaey45p5stnnGEx8s+1oIvspiPWxoGvyrlp2V/AUd7G
rV0HOYOmB6bN6f7nEv5tVDckG4S0u9wkJbonlKNXp/XvtxqK432BUS6IH3/6428J
d/I15yWRFvL4d00jIzjhYkHmlelf4MWVvz1r6hn+fshyzL7DhDUZ0vN3csTYmLle
+jt9IZBthHQhzFj5cgyN9mTQi9v08eGDSGupEof+OSdJIatCyq0H+C/gVtIj5ARq
0LjfBTjQQcnB1cidJfkKjUuaWkvku/mfsDCB0qK5VpuybxMcGTS/6YD6/vhjoUG5
txNuJfDKGPTKpzUkINVfX3B8QniOo2mv8dxVQE1KerYcMxDif5/RDpryLr+b9bJK
4Lwc7Vx5clAoLOtUnoB1n9hi0yhKvDwFSNsb1nYL5ySn/Sb8LGwwkpnlcH+g/N/6
Wb06XSxX6USZ140oeNp5p+SLMKj9daPsL9o2E76FeLdizhWd7YqX1Dexj9rJrJTs
UmjiD8blm2IvPFw8BoYPg6mQ/smDIMHHWzYtoa+HjCQkAm7jkdJdZgKSXDze5rwi
tIL/GR6wHZRIF+VENK491pWtesqrFo/Yn/m8Ubug0wG3wPlzIkuM3ZZLP7ZU1Wxf
OPMQ8fdj9pGm/DJbPtrQBok9wkEeNhHeUDjijy4ZVbaHZw2n2ZrtmryM1mrAwkfd
6zOwHEEX4aZIP2fZna3OstDwqvyWykguN0EtqUmadm094UlV0VP3dyeYvQ0/XNGk
by7KAbDQjiXZ7sF5lxCpZZdDnO4vK3oXXN+6CaKdz9yHdOyEo3im0AroZAs7JUF5
wRHRtw0Lwp91jj9nSOgszs7zGyPuhYCCDU6k+FQZfIpy/qB53AbhaiVprk1oYhSt
QFaJG7fd+Q2G9RIiv3tNTOKnG9Mwj6uwz11mN3PlOqQHYLCGayA4uSHtzhUisBxB
KdgmHxCLsw/RC8zddrQile6t+chQMZFMeIxAjhiC+xMsAyCHRNNqzt55AhTtKDZe
GpCq1nZxMAHveGwoDqOkX98cWgLEo8qA71u9jHq4Uft+Fk4zgZyHnNxgyv+o6sAx
BNM+kUWTqV47L80f9rPhYKfq9yE2NHLUPpQmW5cdMS3zPIm537GNfI43ihCpSq9i
46USQLRk0KSuAuBgvTqGH/mvdMeqUpL/tOU4wiJ4E/wzSRqsRocEX+fcB5IeyHqE
4yFOFbE3X2S8QNcwQ0mgpu7yE9yfAxl4UXm8gIT1OyWRywEEUzD7Mkxm7cCI3NBp
3HZqKcttvKjQetqP/U3tK9BPx/17S+VSkggQm6Y/pvdnz8vBheOcpfdxij935isI
RdJMGzZfV9/1uc8DLRWA/AJNE1JfHvYFm/zZYvTPsEiv/0tn2v2C9XmB7uC8R5gJ
3OT9A0Xq/2t38kK2JMkcKXszx17ksdI8PgMsPVkYKzDT+qEeBanLLc66+kBpWG9W
6TIqrJtSpW5DLSpCMs0eyMyiBLa9Ze3flXqZnk6bRcSbfbBMOeRji9/ZyVT2RIql
gTQ2xe5Cmh6xAFL6jYJiUdA2GVbcYHYrX6Bc0VCedbt36GWLlQs0pYsPwmgSXJOE
n3oQ3yJmZSxdsXF0vPk2UIK3+UdGM16VKtXa1yaLqXdHDzBp3deZjMMtBqzwZuQx
iM43VSWlo92oTznjYaYDeETy3iNpsWIs/5RmNgtcaHdeapF3qyc1/stCFc1C3AXS
eqQas53P6Z0rzDLtCKIjeGzyX1I11lW5GjysUeAa8R+9WSKrGaxCHCSmavVWrrgQ
SuPeVNqywWuY2Tt+flrO3R5/gsNVuZXm5Q/gAhcmgcy/lBWjlN9j3ug04oHV05P0
/mGlE41sj7TvI1bOGwh5aqpKRUN7UgxEPOMPixw5Rq1dfcL/SZ6wktSlp7gaEYXC
XQgDfMkr4SNQKGpoQjXVqD1AQF6FymJH3PSBjtsTI+EiFDTHcHuxgaBDWgdmP1tb
k3VyXxVnlg+f0LDpgrd0/rMwbbpX4Hz9lcMkfW5Kb/h+VCmoSOCV3Z8zG/8Md1yA
uL3qzkHBab0BKIO0iU4uaD43/gq+R7TjER6Hu8Wu61cQQIBh0ENrrCrtxo+AzeAK
IWSen3JA62H3bgdWc184bw6Bem+NBRjya48xkkVx8U5Pw96ujmS7YXNIs6YSXfEp
7JdWTJkoG0nYXi2BL91Z5ZgG22eFLxcvM4Rt8s0Z+0rKLuSbQICEixSK/RhAYk0k
c8juTP1rAxjCYGckLjoq0sbPIEN00bJxEcy8GrROBUWeM7X/YXsgv0Eq+Tedl94K
FfMjcK0SqhLjTnbqNl66t6Qr7b8xy3dFcIdmyWDaBSIyBh11b9MOQBKyhNTEtgYW
m5/bUP2VfalXcaevppS01JddOCa/exEFzveKQ69sDd2BxAU+e1qv8AqpUlQQqYlA
6wRKNRM/SUo+7Z0sppddMN3Rt4AigWzjz8WuL5wWGWwMvKfU9WO1X3ciDegCet+Z
iYf7uym7HC/UmK4UI226R1gdOeh6Lb1WFc0X/5KGj2Ado9qccFNAtbDuXar2DT5o
JB3cbLc3fCym2xwUlGTihWL4iad+1E/Jt12KgYMo6omiF93O0ZyD71xw7ZAtjfN+
A6jlRoG3mDmdnwNb6zbqgs6VMgwEbr+VeKCtWyLEMMgNyw7WovW81qa9GZNHx2rf
LstWbJ80rDUgJ9rcd9vkqfZ6Zz6oP6NjL4mmcDdMQ9cqvqKPW7ejYlKeZsQQCw3n
WjmhAgxaRfYfPvKUG7C9leqz9/T+Yr5Q3LmBco18vZ8HwRWnms7todPdXqwNljVQ
acVAEl5OvRkUtKjNJ5aZYd4WhYWD76rbsdLhM4BWzSJaRsN6fEHY/cb9Lkl0QY8K
6MI6YKC8vheKpT00OTiGg8q385vWquqTXA9ZC+0eCv89FChzUdeSCqw5xsVIHaDx
zMW6NqTu+t1fYhooWzXXJ43w4xqZzAuXv1tpxzavy3lBCq8wUqxeYNHmAvUxCpqd
Sr51MZNgKWsnv6QRQnvurs9py/2WAxO1tY3H3MZ7KcCVuU6N7ijHZm1Vbl8EiPlb
jcaEF/88qA6oP/0dza87RVcGbnVrvDZDmW8+1qSqpfJZEOPEaI4QrPSEegzeEpnr
yTFUtW42Ola+lF5g6aCSc2CGqrxUAYOhtupbDR/h54pTR0SPgEcKQX/gzQOOOaHL
t8MrJHs0OyPMyxzcBrZahR6h//3k1P7b+HtLCcnzWIPAGC2JXJMJHOKhfqb++xFD
xVgznGIenzfwf4W95p7/4cDi8uvaGUnepY6BUZCEw972sKffulHbM7lFnSkVZsBY
ECQ3BsQbwXGC0zc5PL4Y4Yezj9BiXige42BvlERqCGgYxBaScaVHwmN+9BrqOFOq
bsBugOdVvi1eJz5i3B/jVkcya0bTITk6cBKKjuTbEnBgKyyT4ItPJ1ANvBpU0KuD
J9JjsB0YjGqK3MR/1Qt8Yhw/oMYRA3cnO62vovpSRBacOcUoFQr/1GdToO326SEv
pQds1dn06TZSayPITUY5XeYGxlgXX6dH79uF4ZA22SpceRUePxyPDNdiBwbPcqFA
ZJ/MG4mgDVMuWNUeNPJpjlzXDIM0bq+hdHIBKfyhZDgJjPBw2s4q0lufOpCCOYLU
iP7qIkobjTUHVo/5ZaipfmwQgdS4P6hjgt4AUJYSZrDjZ/1Gd9RzrPBLpNxUYeiz
ukW4IAcUYC5h/P9xRevZf0k8xJp3cRHr70Ob7VAnJDflFftwPh/OHEB9lmUfOXKe
2qpWLYFVWQepRu26/aPuO+WxXbCOiZqNkzlINXUquCnT1jaw94VlRC4/QOg0xLs2
yWEGmyqgD6l5fPVdmZJi/O51fKy9Bk+nDDVQGrDSMsY0QQjQkQzKN8jwt42ar3eY
14hDCR4PE9eFPIEPX2YLlnEbFYdgRUYiumUi+JEvE/lV5yAGwC6RMNyyJnFfvhA+
TeR8w/c+r90zsD3KnJ4m9icBGNCrEsVKSnzFeH9lQSVtZNyH/DRcH1PLPqaRiTu4
KUQ37Jzu/yHlE7V9YETjx6+CF1BpYAlqNoGeNMu1uxIj8niCOwphHIV5o1ik8+JA
B6qZKAX3FeQJbs4QFuqo3fCR8dXZKJ0yf+sWognpndlzY6milca08CM0oULsHRtY
nrWKIwv7IcHubDUeKJw3AiFzOsUMR4U71yRMT+VautU3/UuRaq6v0rhbmTp1X9lF
2gLmdsLPDCYV1yfkKLGTk2Sz3wSdLM/vGMxDoLoBiQmwvmPePrXst1VvJH/Hoxm6
d85OaqGCt8WJezWTtvkFKLVEacXm0BahJ+UawK1BT8HJW5KdQy/bJVAvuTUpwJYj
E1BgL+bVuruwYqJhcw6+6NIiK7/SY6r1D8s6d5zS7zNKrwLv8yVxbGFLsQZBLihW
Kr2P9ebZ3ntq3T24T26ju/VqIGXYcItJxabjMBT+m5vG+lpeGLCJ2fE0Tp1aouhX
TKjpmCu6VjNYZhH9O2To/h3TftO5QrL9fyFhfVHwIx5dwJBeG1lufTb4VQvnxMzR
muM9BLgPzxUH/EJoKGXFgJVK396dma8LXubChphPk/j4GlSyaWR8+9a4nKvQOtnS
plI2HrlNzxZyPyvmBiKeaekNE1tvkM3n7dC/mVJIXPN/iFFnPTmnJlj8jQAijY65
tkJbN7OFK4qQsmKEeZzoicMaIgT+BeTy8R6jHgOrO50YTb8L2ulKXH/h2PuxlEF/
ehc+/g0g3k79NXfUg+ACw8Gh0kSJGrAspUtzDZK4ux+n+b+k/BoHpkamFeziyun2
BsqNy3Y1KbDrazoS56z/zZRX4+Mee+XbRM3CU44SzSV7/g8KBenV9OfZ7V3ez5QY
Hs3yYq240ZwAh7Hg2kYMeYlgJneJ4giHw8UxtFueoGDs91ebNl68eICr7q67eSml
xk4gQ1ui/h3Q724O0GtClpPg9wifQRAT69mowSdAlbU01x464W941uURIxXmRpvH
trJ58EuVwTgAnc5xTDNAsM/O6eeKlYNHxNPykn/TBhs+Zub3GVpIyxWqB+vyvWnB
Sv61OgagheqM6FXTJiABQC6gZEB6aPXpQ88/MrX5rs4RJDxferJImJDyex9MyzM5
e89BZs8VDVHoYoawJxfi1DE5JUvBoDv/phjw5g5GjlvO6dfVt0/8Dl7165LYKoRu
qhh3wMyE+gyoT0AkL/qt5BbCoTQKRcWCiCNWfOtaJe7wdulxVdSKzZknLmSwJwFv
HL6pmWspGvTRGq+iqP6sqnuR1CJKZDMyZCBJ2qhpY37M/1Vaz5jrnzM5hM31jzWf
/9USszlC2Lo2f0qj7xRInWXhEGKJmSRlItvGnKy0Q1VXdwYBr04nlKFRKQ+UBpmP
zhO6jZD5orbjWWFoWkyOwwxnXh2nr2TQZQKPnJ86QRbmhO4lfGsgO13GusPyBzC0
lFODnbEzpCZ3xDLcX2RjOJ4DzHaiS8wGRGgue3HlIR+zv8hRmqqdiEVFnnANS27b
A6pFsB8njBvJls2yh+bDHl/9t4GqpU+KUgY+H5g2e9B6qiVQAOozG9TbtgLKCfx4
VuUrUTFUcSOT/89TyHk+Rpkjzcbcz1ovg+Of7nAyeXzsl1Kk8ABGhJhp1Vutvq8T
ey/aLWazzxHRNQX+Zj0MuFvF0sMjIqhnNd2Tpr5POjFL2kLWLNohZo0aAIk2tzwD
D1PfbUFXRasWnuYBHnAJNvILO6OqDz/KPV1xLz00UbVLGt8HX/7xMOkpx0H5cJyd
TpFp02CFiZiDX8JX8/6/Jm0XGa6LJVY9R60PALpkNE5JVTdrO3LGAfRIItY0NbnS
XYIyA/87+xbkJP4lLD0NTpb6qxI3QTE9VCcuSGk1gIf+OT4+gTPpLMdjIXbfuB+i
Qr3BimFbc9wMwB56iRP1/d+jLNl1Bv5QdvGDH6KKthMQJkTL8wWjF4os5316Cti3
v2SwDrc+XCoWzLYiHQM+IHLrK4lN57YRTNZZgIeBsoiEQAL2Fhkdk2qH/LIhQ4iH
du8XyLf41A4z8CzAXIDe6PriorKK3AYICoztWRYmEVJ6rIRa5HHDNGiys65vlE0g
N5mK3eTt0eRxqs8cxzbFGglM4Vrt4KmHMICkjjcv6jHAP3S6nDV+bgbrpr1YlVVk
SIisAbDnJjtAwDZsc7295316sgNhAOwiFsD79/q5RYHHv7Shud0uEC/SMvH+RkPN
SnocVuFafZp4O17XI2kzKwjfLl5D66QcQfGv1l3ScCcn+tC61RXALWBCGJOOfbrw
citcRMl9S7W5uyBDenAULVnHz4HetBo3QubXTUM3iPsUJXvQe2+jfDr3RfMBCcdf
ys6ehD6tV6+JWuHsz4coCannuUZpE29tFwDEPaoLAZD1jcP6gEAvgWdQp3/KdXks
tA+rnNVjNoXuyh2MigE37l3dAi7XONgXwnSYzLXesg5yvtZXrHq88WafNIpWwC9a
t+BAJUXUCuxnPZsyBqEqoqK9hT9oWiesN8gT4sRMdwPLO3vzOuCV9KpSbX0IgoLc
XcZUnulLMkSx2c5OHLuYzlmdaubvRAm4wbVaHID4emlo3mh/mRIrLXnjHy0OdCTl
IwgjpqJi9RmYCMnBNhQzEcIW+EOFymIBYvNdPtwz1VpmtmP34AtOW+18E3u51fQv
C50OkPoGQ7QcVgnGY/8djqfqQueWceWxkJ/M4Q+HVbtfTsrFv26GfqGsa2uyNedS
R0pWYvoVSxo+MEnX93Bntum6a3ux4L+oV5pIvQu+Xwwzw5nERERzIY+yX1Iv/Wb3
+ScA+3Qn2DRrRqwFZdnvidUtq+Q1xr01+4qXdFc5pcdboG+yug51TXXb7544T+Os
miaNklLYw+fmT9atLMIwsnKRKUo8Xy491bjr8JfMeW5Z/hgTTri9GXOHRWgUATO+
aQvhuiPy4+MhBBCtVMhoD1VzYlD4W6GdePcBLTU/u7iF/Vq36kOOqBLIqWy5hiYE
t5k18ZH45O1w55qXr/qFEtAZ9ZRlFIhfR4Z2l35saiQgQD6GesT601Ffoc+uvvsT
uOJbAmAeNBVpwR3Lgvgr631TDS1ZCFolDJhDyinAowzSBKHfhlHYG8HgjNFWsnBN
2tOFB+MNLi9NoWbupKEn3LEioNAjH+9OgeVJ4SJKWhTYc+jK9ot4Tu7m3oOh+39u
ziNGUG1++wMZsPv72+smlE6zc4orvREavPO1Y6Snj+tAtK2SBPJo3Rw9lpL6fEaZ
rEfic7gg5wQTOYERc9OakKBAcK3DrdxiFkrYrV926RtaPXjgPuM31499lCd2XRs9
jBGZqqvJRpSbfT9tOI3okqQ6XI7wuyTENnUWlSAI3hukpZWSr05QLZVrlowluiyV
T1FusSF28InT9xEGQSB49wrT1Y2AXywwx2Y0o2Km8YNZipcQ8WJxxCCJyWfj8gdf
5f3JIbBLwZouzHHRUL1vZ58ZQIkfP/ECmX9FaU7eabamowdhSi3qexIw+cJLO7Bk
SpBbYY7V069xSgP0tTwGZtSQpZUaJbCzW3M6csvFS/cm2xCrU8Vu/UZrUXaLnjsY
Ke5s35ILfxoNPOVMHdtMWKWAOZo7C9i565nb+E6Sii/wLQdehpiMgFzKoKPdc/ay
tcies7rM5K4Kbq3PJD/A8DiublznuGfqXNYuKYD704sgr0NkW+rJdY0hEKBwmvJl
eqwEyKAJo7dvyNEnC1oYtzgE/kGIaMHEVeahVVq562fdVOAxD7KmlRS1RJuFUYyM
F3WNYLs7rPLc67kAPqaThaotdcUHeyikaAiRYfThOdI0M7l1OMSi1RKFBCbG4QBB
uSmeIvyJkrsb7tFZVLPnuBCd6iAO5vdD7UqhZy0J43eP01fzgSWBYhc4dy2M1sDg
wldTZvvBjqXBe0umBRl4pZWS5ty6axI9SQ/C5x5junalo/ZjFLE+otokLh9m6xuA
gQ3sfbrTIiFd2fsSXR4rsP1rnguldxwBntopMkZj9YtL2Yuqq2jPw3kpSnj3gM83
ZFWj0jKnDIfYmnOyG/OaXC7eS2gGSS08LGQkV4Ce9o2AiwS58TZ4TBsw1vjsK9wH
6LyoWxYgAZM2H/MstdDLqFdgs3eDrKuaTPtvytSr4LPQXWJCFjiilDHOpPO2twcI
2AxEAEWqNZOFs/WxffWgaC3o6Yrboz0XErTnxyYB6YbkwzrpQGCKNM7VhtZsTKDU
4MiDx5v7mdDrv2BHBRh2XexSet89npGMy7yk1L0zdDcHl3OD175oM6uftp1YeODS
FVGBPSvEKdumYZ4ptfz8dnDwf6Kbuc14+ZsNcMs8cv+2u5aKRVxMyzqpzeITgVTm
+Ge85X9WQqJ9+GgHwyg1/MniJXNnl3RcGVTnzjm6Pg9R00TTcHnpXQwoIdIZoDZB
dvAqBxMSfYGP/PjU9wa4WXPZxomMrDTgQicX2aNiH8ABmw6LERxwf4AssRRRzxdx
MuSJRvXJvb/2AvMkGY3Zo89qFM6qdZSoHLoyelzKaLP+mznNH4pLn5VBi83nfmEG
67wy6hemf4h6oKXIn30STfr0Shuqznmp2rXh19dPXzwqNC9ybAq4J+SDm6X57SjF
qaw6Fz7VyyZLA1XsRx/n+QvwY3nA3oS68SW67EdhupdT3tgGkOVAR/P2FmecLNKS
4jyKkeHuSGXHMxSbY/U+bZatR8cwlepnQYw6L3xfpv/XtTB78chWnW0WJtNok2D6
Vgy92pM9/19Iqn8TwdsT2IeFm19gn4LMEARkP05dSVwQdEI6xo+ZF9QRdRvul+8c
cB8cTMbxC4xQvCkhrMJrywgVyk1TJYuQU/C0CwQUz7+NmO+ZM/cZAOwc2I3nnQmG
NVNuVopw0SGai59I6XgbRAkOk0T/XIP3ppq2LdWGQ6wMPFtWx+FJvr6pWx4njFEE
0fpauLBj+4XFKECYaT21oGRHXZ3GoaX+qjDkpmdQ42yfrttta9xkSxNCAWSASR+8
iJYO6twV5OcQ7e7eZd/6AJlfvnfjoUr1NwHQWHceJAKVuYILliREn3S7UtI0BWJV
FBMVzIQtekd8UxUdJOYiV+qHKBE6IE0I8X7kLSlwTKu4nXc8AGRuUZi5Q+cdjS1W
Fm8Vm1F1yMa1cigvbNm4fuVrGcbf2981mxzmx0fONNUS/pHk7wGJkFL+aAjVTEkO
Ipa8F0gjaEhs8CH+6Q60zWuaig91hQs2e930mBqWaQhtZJdabscpX4eNreVxOaJ+
lEixPz0m3WcGyJj+I4r3rUoEpn4NBaUDSlfQJUvl84/kjmjMHDNWTurqYoQohB+b
f/EttI++HnNi1q0+Oxykoa73eKloejK+uOIGx4AODwjy8VzfOlY8xN4Yq6QNIGoW
ERQMz7Jf51RwJCVEO4f2aL0Zb3NwGB+dxW/hmwHVozaiwxm7ucutp3NS2iigwvmT
Bvy/SY6XwqhFFAsuYM5fA3jpIBynCFuZyiOnKrwI74ZSe+f4q9tIGRUSl3+Efvrm
cUuq7dzXuMEn6qX3hgBwSjK5LsQd799LFuuoFw7Pg/tYE1vIrUhUWGJ0Lg50p7tG
YUb2vncokCsTeUdOfeFxwUQeunOvJMFB0flDoNbVuzvLuZ09K3MZ2hYPQDDC7x4x
6USV1NzRzz234UGok1OT+rIaY2Pwz0REZMoLGUIWX9YjjwTV5EJdA4ieWkEDHJec
J/0JdXMZfvwCEWjjz97XepIBCdALceXkEX717VxVAxuJCtI5mYYs6yVMZXq+R7RP
aTX/3OexFSuGNUJo4WATCc6TwTcwzqrzAwNJ5k8WMpIFfnbVrCKtLxNRPrhGPuIc
+35h1zZ5D+NZDQ3/oIFEgpHZiKvVJpmbRV/4kNNbQB1jFcT/YKGlTMptx8C6Sp25
BaXQMY5RBN+K0YAfCdNYy0J2rY5VzgZla/C/G9FjEkCpC1d6K0TPxR02E/GzrhH5
YNDzg1hum+itcbOChtCwieHott0BonPsmwZ7SQek4Uu6f75Tp7pnYC379VBz0Nh6
0xML9gbEkQsSacCtyY1oJF9bcZeU0xUkoddleQWoLjwYJKn6wVDFUGv36B+PixVi
zooxNyWbaRO8KDMiSHL8UpaQEwbOV2oWiOtzXzwpnIzanKbBAjxHxpYILOgFOw/K
XGMQU4M6AEWccW4r+zHh87DRRJSUT1abGzHAn8OxupUwp0yiK9xnRNqCcBcCdNAN
tqXE5EwCsjBZzfrd1P1fary6srUpFyKEwHsMCDKol6OMYOKA6pK4tWnkWfufBCPA
GNQCKIb6aDHvJZogvkjNTPr4Qk2yuAaqlqqcMRmiAKtvpwGSltnpZigmKoW60T+o
rcPVbqDlB/NkAx4ueZrAidO70bAHe5j+h5bobIy5wpeZ4m7K0VD/ZBt+e1YAkbOm
jmcdeFkNhuPl3qbIsKbJO615pAatbsv5/fwPFmUihVYtWdswxIvvLk/5Y3GMmYiS
z5Liw6gSK/HhFJXN6AKsd72ArLeBHzkXHfyMta+NrZxZsxRIgou8QqQPfesi6ArC
CBXJ1/Oq5uTPUimXr/B8V+PP/J7nPiIKA3N8URf0tMfPGXI//DEaYPy0A44t3q8t
bTGqW2RNPexBbvU+Yo5Bq6lYDK1TAzjiRBJwpFaKBlEXiTUL9pcwv01Qft/1Kx2I
Yo9Y40JQs9dQ9biGSE0IqyumYINQC2eSU5SBiRNIa6z7NnMl3bO4/V9PDjubHcCI
uyGfPUimQmNrzwCLg0ebYGHUTknVXeTArhuyI+Sx9Ny9vyYzSywu86UZH2fkE15l
RvTFrLaxsGbSpMNk5mj0JgiASHQwsgWzC4vhb4Q/OWqQ1APNbt00FK7Rlwy8zG6x
CRa/n35SujI0sNiAcpGDUMIdEEg7Z9s+SOMpMUmzgQqLMFC19e6gb3OIqUiloJfM
mVfIeOPYRebJSO+zNQSf3v5xFUWEZQsPY6ZaPcJeSSS7sdt0HYO2sMS8KG4t+UHJ
dnjOV5Dr1gn7OK/tp5C1u/x+6G0HPch9FWpsTYJnMOd3mxZ4QkEQX/E0p1UXkZ4S
neW9qM6dnijkbHxhPWXEzAc2+K9CFKRSM/xdPrU+wqHdpG235ECrsBOScJxqMqcF
wrV8RFMcEVYSJr8wmWXs/1ur3guX7OsktU4pGPR1EgG0hJ/ItsO7YJu6TvFODmz5
VIo5LL+CYjEcSSt7RpUuVcA0iY9/JPHiLpPutvO0AZxSvBSZaBkao8XvCMUrgYRb
dhrvqXR7zGVBduzRm4Nf8uvmlO2mJQ5SuZfEvzv6JYvirxm7pqM6GMS1a4Ocd4j2
3NbmWn2/PgzD2z9ylaRM1MgstfcrrrwZs1qqDx6OJaEkqOHizMS1SAo6awL63z3x
BVSZducVzj81P3TTFvdhE0rTkvQVtKGbfnnN3VyhwYt/dxZ0MdGecpOKY0N71z+4
OTMg/rvskWVUPjNrImjuYZdYciH/4ghF46mQ9xV/j3YkbMh9BSTTmoslsVaNbRxK
T4oS/YM12m2mZPnw21je/O9UKYH1In8XdbJiLTbJK/dLF3s70FGwyStLcBOGcUOw
P95ve5A/whfO58qXVM+apMEVvFWM55VQEPoc6GRCq78Ey6DRoBsryCoZnh5vhrv7
M7em6ah/CDViL5Ap+uXdu5HvDMHjWnMVK4RCNaDokBRMHLZlmCntU3fzWaV/wKvz
AQx7falcpwRGHR7pMGSUseEazDmsleU5A1/wUINw/3pXnR+BRz9LnCTlS8s14t47
2nvupBQO98DBus7PBFB9+/Zt0aLaExcC+Y7zTDlkyoPbNBw+X7KSFv+sJOcAG5Jd
tdGDaC2XpFTYVY5KlYs23amUDmpTd5A5oW/joa+0H1YsR2yg+pmpmZSljUwej7WX
Fj9lpr+nQCbRWaFU8RK56XV1eUlwY8JEzplmEkLGfsnuO1CVppf3AEUCwDoYL4f3
wAy/rhjBggJO6bbxW2sHJ//ZIC0xBkqGaT+1+0Et6+Ww4adb8TwBQZm+3aHs/jMu
X2tdivb/G+leenDYtVXTVwdbvqP2ey1REC6WCKMboh2PJc76ZmHPN2oJ8dVqBX04
J9yjzv9tH1n8Riznok+8s37coIc9uHhnVksTrD4TvjndV1FqQqe7///RFtIWylFN
do+x5nVDoJFcGvBhOH3GaGNTj42l4Lm07FOr49PFKSTf+Pl6qFs68jOVokfP3H3I
5CF3nmkyppIA8qtbexUQixHwTw9WUY44wHMdxTQY32WxfMEflxU4kB9/bfFzOAw6
XTx27iGYLL7l/j/vHL0oOXdgqMN/y2Ly9J9RnlJ+017AEeDuuZy0d0XWB5u9vFTg
jVLj0J8w0YAhXBW7Qbf95I9hh0hAX988MI7r0f/6+UsiF7+Wfi/HSzhuzSJki3au
WipQWCAgyT/qc+AUsazUCU1cm2RUdFiV26TqJ2W51BU/IMAuY6+63oksc8/l52iN
bU30zhsfvlOZ3JffD22mseh7FNbZWaiYhNGqeBhz2mEp0pjzTJg3n2QDNgnb17KT
bo+fkY8GeFh/w//843FlXrS62J2eu/0wH66KPpK4GYxrlqtyFhIqPi83yJTJzRUa
uNnIy4lMoQMHqLIrxfYV9GKfmpnoBYKKVkx13T9hZZ3TN38+hAqJpj2oloo9O/6d
ikHHGfaPMk2Ocp4Jsex5Vn+qDwGQs1GQuawkvbM+XVGEFyj/lA/pKgvbCiv5MVKK
DIF7yMXVbf6GfsA/ZTAYxXMTggBJ/1tRZaj5DTWb9q6VoFbEM6GyZ+ZFfLkN+4Vm
98dJrjsO+duWUvDX+xBqc2WieoyQ31dchIGijcWmcgvhmXh7gjjvm21xIaNvkQwh
+oczgQsW15M/HHJGNp6I2xOYRGdz7Aph2hFCa2Kai0rrh1t2E6I3vmdqUKUy08P3
xjG9bgeE5YfWxnsymIMa3SulYndo4Ek1ujpARRsjqoL2k2b8/Te+ksd6lebjQyhS
2N11+cIXopTC4pC3Km/jghKcyw5PB53boxb/kBaETPutrmYOL2S3/31jhsfuZiIa
A6JKu0IvW4UY0sjz9clhwYCLPfdBzhnWCC+1rBj/jKLMZpyiP6apj5tzj65OgBV6
8IXFtYCBCthtqE090pAe9iiGyjCJfZbDOtRYIjLXwnukHc4ytuGoQA/CgUUl6qBN
a+U7R3mV39aAWwhz7qGzMbBxX5hcPNVrN+e9oU7609ucJjxnuYRSLyZRKLNQB0SC
ynUtbbhPby/2mvXrVeeiYxfVQVYWG0ePoRxM+BJ9/ryqx5dq3GdN0cc9zVn716gG
CfUA99qq5gmrJhl1OAoaktr2beFO741tTPQlUevPWrt0wzVqc1mXZv/eTC/u9gVa
va4W0WaTx0Pp+4Npxi/SN/y8oN2lGl6E5HGy8WsiwTvMxDrIw/zVfoMgwJVXL6gh
n9EbIosiM1dBpIBOcniAOz3UGAqHCk+wLnsvyC5381icK1xCe5Bi07uh604g48JG
iNGuR+DDhc3xJA3oWqt0b3xlXe92c9gfhIpI4TsVV7aVCWDlMaaRQkNLlg2XUqsZ
w0pCSSDeXbpo4kmBdCXelGvdUKzoSJpxWZeWJW1ve/elfvO6HR7DAEqT9qNbsDLQ
UuIPvAAg0E8SzPaYBEG7vjjnwr+b8+9rf1TxEP9AFZMzJU7h3SIGSEe9IXcTk/Qg
WSqkhF239R8N1okPR17KGX0G/dlniO2UESxzMo/oRbls3756DKEaIAtj4c7ZekK+
gZmAV2vJbFsoEyh45DPhQbceTapv9208m48Ci0qAeEqRyIHKewh3X07thBgSQfH8
FrBb376agVvu2/2pGgB/ntnMwelUTq/QzaKSOSXWOFRkQJZ2WRe+TjGjuDMFytQ5
AHMfF361xOgvbCN3Ym8mdWZ6pYgETVNAF5ja3cSNGkoTj4S/qYdSnCe2A6lIp6xb
Y9s7T4L9b4QcFMjGEJ77top0UR3RS1R7ZM8P+DtblQfPbZVnX35yEOqans6gKnwG
eF1P1oVAQ6b7XZUzMIo2QQqmnvnXFjntitUmDuckl/xk1CkxPBe4zJORjT8dnu6P
Ox8+2QX0psiKrpPpfS0bE3JYtseF9b0UB/xDdJDEC0vRABFYmmY0iR6LngyDIZo9
QRlpEXDUP1Ra9vDptZXYfjiV9NUoGKvotlFc8ggevuGytivTmCXEN0Oy0sNeqBSQ
r68YG5/hn5Rev0lkXP1cFsHdEGRn5kz0doJArCcrCPc+/WXUfTTekejoonQ7DYIF
PrAPynXPGqUZiotEeX3C7BnEpc8fSIY+JHZf3spbCKwWXq+x6DHjMXMXBI2NpIwm
lOO5OCa0o+8DYAdUy3Y8IJ1yuq/SH5Yer8SZpNcjVWTvRTLxzCvuEA3slm0Bgjip
HYABBXtb/ceeWr/nJsJWHSHtyMG1m6WZXdOQ/Vhgh+n88qbqElEJCRv1F99VKGQO
qPcPaTQPFKaFC2hz2MlKEha/8q1XPLxWJtHzRiiafRVJSbrw9mhBt4vrc0OTqID6
i6M47BfUsJ+Q5QU0IiCkib7fd7oM8WYk9esZW1/YeQ5a2ttgI15JPgvUOLXyDAJg
/IP+qowsDVCFA3P9DsXel2Zzjae0t3pBJHGA3fomRQB+4hx++oebBEHw5gvqydte
W54Jei6MY8D2mj9aBa8oH8/SQg4+AP3bbE1FB10qV1Ylkp//iOUp8MROXKC1vscZ
j1i9g1EufSGCp1dxLYtTeU0CBsE3WnHD1KnOywWjwvrM41+af8Qf/9SMNt6dIq2W
CtV7lRLYzQaI/fZcHGtNB6ZKHcemvy8Pkm8dtZgE5b3qlFPqZB1tsT18bqVU1ugd
hTEGY77guWZlylkm2HaRHJrkoLYronQzcmOyktaj9+PFebxiZikaaA03mmkr+EMM
G+oFFgmom+Z/nBzg/10tHpF+PPx5miLk9T1Ry7oawTI+UXF/gAw7sE5HnuPVv35u
rh1cRb7mtILgl6gBmq3NAWsboY2WdnPUzxyhq4DcHA//4tx28MDUOSXxN3bpbvMk
kxD2jTouFyUdF1AMvhAl8Xub4O7rxvQXvJTTMBSczdqZYWlbUfH4iQY1ARsqsjm4
pHws3drSG6o0pU66brfpIgeCshnl+1OUGxNl3lIiR5UgDr+ASy5lu1vhcAj/SsUv
PCSYJY4R42mzsGWgS4KsiuGfVMj22c7Er23tJ0TePfjiFU/fmE+u2m1LMPj6MdbF
gi0XNDIyodT/VbLtZfWBZ0V2lcJAPxj6ma6kAfqo9ccVKIrxbaOso1jPS2MD+fih
7GsIs/uOKXpNF1sZvzXlKPGAOo8nt+/hRBVpTjVNErtE0fJQnNjFmrw5x5FwqK2I
IRJzc0PLQgp16Tj/igv2fDXNDImZ9tOTy0tdwQL2fdsgkhfaoH/2vKTrcZRomiPX
Vb2JvX9pwfSGAWpLdW32NSkhklABgQSe6WCAVEz3z3/w+asLU25OP88Vo2ass2Xu
2fL0/fvCPj0USr1NkGqPG2IOjWGqUp4ej/0NvwRaxYT2O4gknP8FXIX6oUZ3Ik6n
vMiVc+W5VB39KbBkzn1xcu+LU83RZ49tmI4xJv2jdRMzeOTUxwrvrsF7Vt3QCDxs
2MqjE06j0HmKXmYGkCF9kvcVjyUSIyD7r6YifYTKsSNf86Kir4aqACXx+GlW6Iu1
dwT0u0wKGHDiSCXAkUF9vtIAFtRvon9dAxOsgGsCuCvfVlzFLmFqBKuDZXvcFA3E
4pJ2bBByw/K6s+mbTZT1/rudYbKNwSyZ1/DIulL2oePFs0UPfTfRc1pgxtfss0Wj
AbUTxDJUIOIUpNtUuMcrKSeDW3ABB/eJ1IdoDbxjFsCpTWI7V15rsrD+aRCJC3xs
+QLygyj0pSlMWxbUpOwusEw4NUPFTIyFwh/p/5vrxrLgdGMliDyD7xAO/q3KNvKD
eCSYsmSsTj7nimXzAYBD9CvTH3ld/e1ohMXjEb5CMmInyMYnNQFjbL7EvBMnqWAc
TgqS0oCS9XceIcsYRoRLWeBWPPSrgI1EKNlNfbaiVYErsrgQUTnc9fbbtvKU33Fp
i86v7aQ171CUY7zGCcdiEhuFFMcX+ZPUkJ4lTU4YR0NKW+BakVDmTTNPslyY55/D
gN7NE3fFD4r0QGPZ0NAoWiYJ/9YzR9DcPllwYLNWEKyWhp4uLCLLAwNmuHpAV2BO
iwph4VGOrYOOPUes5O/6XxBJJRIp/jn6JN/5u69kEEcJRApoI2rgviln914W+oH+
3HkdzDusha3//OI/MboFbtolTtjWMmz3P7/3d1XCfVpA0aDDNgkxZ8W1aeXTZbq/
AgCeyKzMGQT5Sdn/atUqPxt/7XJpajIE3B9zC2aKtzjeWMPy+3LH9pYxyDIXGf5M
uxNdd4qcXUbMyctxuEX7teI1W76itEZuMAzYnEqMaI2IQJQnahkFYgISc1Ivevc8
e+lWw7RN5sxrmjTm1e8QsYyrDAjiIrQbNye68QmXkrXcuCAAU2zkHX65YGHFBGl7
n2dY/oRPx+oesYP4SHFFvSVM1EdMoaHOc+iU3vUcgSTNoYAD/chrfKnG9OBOwfJ0
A4wYPgU6T6RkLEQQN3Y+UnMp4JVBCnu54bJZym+1oXquqZjvZG8EdJ/1LZ2cRCAJ
KME1c8eceG71pYMoTWk9S875jZeCkgNaI98tYAshNvLf3DXmHJf6Fgl+2eeY+ZZN
FGnnw+rlrlUXg+t/egzR4X0wOciQG502k5QzhWLYHphsUGMC7qXEj7C/G67KFCzi
ImgOmAiHwuoQFcDQY2slLo8JRFVvlHl+B8JrMe/jLqc/wfFrKs9LdeTDh9hfXyA5
whlW/rkOUitdV9kNPnRDzkH8wvsgt2n+rZQUJsJ/ggk+owKl4zfQuTT5zmIIdDyA
okqYWp+Nu7Fi5UJDBCgK4uwYth3oZg/AgUOBRsl+Cxq7IXV8S+jEtibZOlCKfglR
Hl3r7j6CRybAdYwD6Q8Zd1ny0Rb6CgBDIUb8X60KfoKKmnmbOUJjN58oAt4uS5VD
8f8arSzSO7MSF79j7NVaReDg0jqEYVal16oNpgzWzmWvS42SPvrqHm8qhCk3QcCZ
QckaJZSx/gOtG2tRmGuNZavrNk91hLFbz6I0pavccGWf/CJDTEo8ykyQ+Q6USxv5
ZZKS4WEo6vv94v18sHf2kjWHAS36YwMlTQs584NpIoBPZuwLicJwfRTtD8t5YPvo
OURoO1gAdzHMvALGQaoXdbSWweKRuX2dUAb5sCvBRaIkSiEuE3WSlfRN1evabZIi
lg8phzOZEdHPFxFtbhi1GXPBw6xMB3nYyZQErNqtjvCmxmdqSx0X6HC1Gd9oq9u/
11GZuYtNLcUjSUBn/Gb/V184FamNUz/urVOMfKrjtoCVCeFl9/a4VJcPb+/H/Rgr
9vmX56EGyOYyL8amUiH2NXNoLJrFurGOO8eSe/NoKOv2VurkXPGsKF/ipD2pI+ha
rOOkVRV09adn55EAme/y5uoKcsSxnb/vAxRt+M5L8CXbLreK49EarDUOuiswpucX
qfXpfYRqSBdX820ZDNxHmjlYKgRxlLOVwCp7cXYGADJU/Tq/WeRvfdbLiF3BvWqj
GzefTft7ivpIXYuDUiQnwi0V+b6TZq0ZB6FSd4ukREJHD7C0TN5c7B37gmJ5cYBC
JVnialaxKS4GGUUFVMrZQGNFMxvMy/K6sqKsENOe+HLpgczo37jNzSdEEnSOZFp/
GSyb9PB9hG4tJLhfzkmt75Jbtsn5bsW3Ajuivld+L+jo3G8O1nXJWHC+0uwmDedF
w53INNDaDmgYwVSL/gxtRyMJHXytasrXjx8/wKhfxPbA535YSe62CkjgLqME6PAs
kBKYjAHg2E7HmwNP0DBfu9iSe6heQjw7U8ES8wBAiLNucw4WGSKpTXU2fzWYCXpg
mxLH2Pxu30Kae1PvDg8wGZ0QnjnV34y7tyz+fvNp/LleS9qBONQWni63V99BHdVE
dAb7qedpi+hiSvfj8U7nhI+WOpECwN4pINZqJ2gwzOGoz8HMMJ/SDz6fk1ef+Lej
dyo0BDstyo500vpKHirbwe7XmTAqUFcBY2Lf1srjajERGSlUofWQ+LUtjMClQ+o6
8ELNzdtAK9099E7ibby7KeEOw+0pHPPcbROjBnIvevSG8BW8z9XwkzTDI5zd96+u
w4wQzfFKGm0+ro9ySh4JTSKlW0fRN08L6dI+q9+As6ikjGAeDreEsHhv9GlnnOpe
tKcuhoYxZJLcUOjAMcT+6A3FBarSi6WWz7E/oichfhzoRiRmFdCSBnLKMOwoZAW1
n+Cre17sX+WbZg6D1yldCEqDpAlD+++xeg0ECXokm5XFOip1PlNq1DmPplESjvtT
EvjYZWl9x7ln1hKIz8oyQbdciBCjnYHm9H2uCeJ/P5duaAWYTRUUcSrAn5fuswoC
b5AozDaij9uO/26SbuKRz/SrosifwWCeC7gxinHN+9Dx6mbyMMMai7Q3glEpKd5m
LR8H9ep084oZfpgw4mHP3odBwoU05wgY9fW07I+KahtI43VFYYXHUjTYh8OQYhX0
+xgCmoxmcZg165KseyVXG9wZDHZkgwIlAuERmkkFPIu1Yc9BmPx11lh2Cbt+FR9q
Xz24e4bIEnOavOQhHSnbDwARDhlkOWLb9pFruVdobEHlxh3HSgnHVv9XXhzgjHyS
t2LMxssVYJCNw9LTVkYhBeHzH6b8uEvt0pFWZhFyOtPpoLmZPnh5wiZxXewAeiEc
DzstmtK6jakksH92kLA7LB4XRKI/+smuenuOC54Z+qUjXjev9WKqZJeRqnSqYjqQ
JJ5PIRcAdVvyMSDdzR15tdx/PcEgtTrxbpw54jxn2meZtr/FCrKACNfiJrQXhyaT
Lnc805O0hFx10Wg/fa7XSIrniowS4zVqTMEFCkP78ulI28YxyWP0oINS6dupSHHr
AQftKevqg0vDLT4/LKTzcjTsLkC2r4BL5WFpEja2IgexAqfcW+EPyFMSD1CbvIlo
0Z2nmNZnHLMVdQ30qUegx2t6DGxHABZ5YFtcKlDNibi0PuJgg/t+mEiA3MgtrETB
CgafDRZrhyTXvKXAvvojTxJLr7LZz3TDNFB21e+fkxIRWx3G5OMQ54hzrpINdyRN
qc85/PEEJ5GMPSyIdXX0lQ4Ovoum+z+xnSIOM9a9+5W5lx/E1ZfIED0++b9wFBiz
VwNKc5QFHmzyRzc6oliHBN4HXZ18pGKaZkpGu1DT+2a7m6iavyZsVrt1iH/2hcs2
k5p9X0W1kkMd0YFZK7t3W+q/gOa+gM968Q6zzffidVb4WxRLep5u2hrWWAOSPHSZ
jqfwGm87Oqt0yE2uARJ1qLy62vWy/FgPexLW7S+tTYJ4am5lKJpDrQPcXcjaYYWp
We3kgbqoSi4LmktUiL6NqHurUB+UbpeYIYlZgfXqMlRR/efj+vdpT3OYHYjdREBa
cS76LcyMPSm1sLOZlsDQQ7EknyUdjP52kdAephj4K0AgUXOIE6RUqZrNoTqRkRAr
jLddVxeKsxwD4W1UqKyCvKNjupi775NvQ2wi+pCe4DN80dwDYIZ6z7X+MEQOm/k6
lPCm85PwKujEFU0MB6+3KGGFESu6c+AbPyytlfi8nBIt8KpolIMheMB//7RqjH45
WjfKfXwouFx3RMM2uXwEnyW3+CAc7fwEvFDiKx1Kdd0EXBifIT0D5y7HV1TyVYvh
/wBP+qXEaxp1aafLj8WgurngbZdG6yNIShx6KV6ac92JQLMsb2TSoz9xKXihP8Nb
S7LKFFGfiUomEkojwl1Jmucq2A4Sh/WClFHyty8PMDfD8m3xdXPwEysFtRltA88B
5dLLEOWJocfeaglYVAH/CDr+RaQ91wnnY5bkwHWxNypHnd3GNMdY7UGUxOFq65+8
Ain6in+tr5bxmn4frUQOs5MXX5DTKNjQ5pxFDSm4379JwL7A3ZgadUPhbhjIcALb
cvMRfflq9oAu8X+vcHu8Y4kWDEs5NyNj2G18WTJtWn/WT4n+IKLohNneU79hm998
iDZjCu6vaKL5K64xE86tOLyS/zyAhsbopOiU98uPdydb5lXQMb43lsIb+EHpcIrG
CyaZbD5zNe0FTKjEd4JRgJYDW/wjlorfi0Ptfx0UJ8VRqSeUh0XAz5kmJhdAoBkt
/u45vbNiFoQVMTaRKfWnAitSs28+Slk6f215RFnPA5Wt/CtIj2G38rzM5RR2AiHc
k0VbrmUUzsOgURJRAk7SpJpDxM6w0tcfu5upUcp2a7wWxY03PxGYhWBJJP83RsyM
vUPcRGGaQJdsg7IJV0H72/T8Y5Dlh7nYPiC+sQ6E5EO7HjwerjVIpe7lGi7OXFPE
G8Lyjo2THz6stK5ryUU9BmKsd0apvhB39cZBHEhMat43ckWfss3I+h5hCYpK0LI0
e1m2ZlQR8tivE7UvA6HqUMB5myg8IkumDEuH2+kFd5wE4N7LjIwu4EaiK16s77zz
+3Hu7GtFMnpVc2G+h35pIvYDzcHPG68/T7NoLQwpdgfzxtrJglAdqNWVNCBIs1AK
BNza1dyXIgWUrNUmFvRWmnJhmOEbjcyo/kiWlIGsuw5TwcsqJ3UpqCuCbC/rgJdN
9Fru7cLfDciqM8w/Z9YNWPYkgjv6GBI237tzFplQREAIhbyto80Jq3bMxbL1VSAh
Wu+kZAvW2zSJtikc/YFZjXxeumI5kzfOA9SZO4mrwiS7SbJaABfIdZ+XA6RjGtcv
CN1dZN+4l1DAT/1yXrhtJbx0jy7GDf1AeXQu0kf2hh/3wKUuxKosApNIp1jOIZ8i
V5tcraTF4/RNFprVMFDejI0iVTunPrYru0nlfwYZIhHOVPh1nmz4T/q0z/dSLYKC
nZGMJW6NHxzTtiT5UhqFMGPCeSWt3rGL3mWewR9KpYDgYhaf3Vy4zL2/EKU9GP37
72o7Ayvjg9bSjadrYUsPT1icZu/pl1wWgHAyq78O4XqQZDZqxV7oRi1bqmFVkr4k
mxDgAzSfDM94OP7a3NJB9lzANJw6oXcVj8ux7BCQC5CtvvlqpZukjiPzBzJ7kQUP
pHn/jaGJh7n/3MazPGAKnsIIPj4WgyPIMg+L9l7wsDfFErSWA/KPPaCYgo//H1So
oO13kvBcfFqWXXVNziz/6J4gjA8PIAThQuiTVFR4BoP8xqaK6Sp6g/02tuF51ARh
v/VQBUBVp8oGLbrrs/6VOlpQQqv/yrkcfCLG81ExYKIS1VIowRIplBv2/VAMX4bi
wLPGlujNUQAV+BWPMscO5QdWFbybpxQakZ4m/GRsWkVxS3FHPDewwCgtZ5jqq0A1
vU4H8jVhOHMewdFcANWk7K7CN68AmIgvNmac6Y9AJ+EAMYWJO8dyHbXx09hMN+tO
tgCx5dHfGbYOXENvkLmPc28FuTcHFKN5SHTs5OkRXM3x69DQAXb9MUtDxIO7pjnt
q3LCxD74ofWWvvqnIOEjhY+13X86CsulpHzN4h706L7Zde8hHzoRphsDIDy8j6Et
S7CUtBW75RrIQ02Sm+h5SpB+G5vvMhXpIH1P2SI73m7oAUF2b70YrMWRnQIHclhF
7dn+pBEutOVHbjynzMKlW1KGICG4pRsj41Q+eMJEkXF5BqYa1ZLAzWSgDGxeZT+8
q1QBqmDvRY7TLQt0AUxUvXIJ+BMresiAuo4OiIYjxt1Xf5B5RJfPnGkObbsthjXq
sNDakDBYm14HWgjqxWtfLe1eaUmrisJDj/+NVPsRD6IEQucwdXXjmQSIQvN5SomO
Bhl01+zqMpN3q6Wi21EKEEXbQoHWxl1dOAArLpR2XjoNkzevZYqGSpPnGsowA3Tk
JS/yq2/iIoSFtMMWjqx19gqXQwLew+aENj3HpdBp08UBLiL9xAr2gAOcf62BRpAu
IM8TNPbkT02UqKtvLWLw/fm1K3BZHNQiJVfW+Z86KqaxyUhJ/YIkHxfoCnkhzXqs
p0mBkle0sypqHRPUKCpKUnPDCtA6996vuBRcsJSVBS1TWHeDCQhmaG1Vr9Q481Py
kufCC69LG2WhOEt4ETFU2aEJxIBAWnKYcKasEvOOF2D/Mi8/G3fWL4FhcyPWZCx6
v5+PvsQXSSYkVPgjYKL/jmDmytJlx46OikmP/cUuUntposOEiphbuC4wGQcMjOyX
PiLyPj8B8/pYef0dVX8VfunIleCbuTFnOOXJ1JB2oaq0aHAqy2KFPeXxFqatuBIT
MGZnXJq+vjW5QMpjRhp2x+xRI56axrPVG71LSBBrKL2EKacr7UARcQ+C8HF7HzV1
Cnrqm+N+FETFvabeGLVaOLEyjna9IHiQeSwjpP8SpsVvRaX0XCqoprNJ2/zFSWyD
euosymwPpCFHiHf0dZQLL6AFOtlSRU9pSu//SXYZd+boiySfJhJEUd5Qlrz6N7RU
PyqmUKGrVxmgH6TaV+kAI5oflWUXlVpSNTBkSQ/XUUcha+IayjUhJt7ThmhPyMo9
9noY1gclI3bv0MwPIfJqZueM2KayyOGWcStJ6Ul0X8ppjtFnh+HF5eUO5q2YmEX1
mbYaxB/pSqIfueVT5cSYJFzVkIVXFXCO+SMqC00KnuezC0l3TUxoVETENlUqw+bv
Kcruvyw84l7CtfjLVVe9vHPLzDPy4GgBINlQ4SIpKzXhhWajz2g+Abp6cqZ3ygO4
DCM826Gj5rYi/3q9L2PV8TLwyTk96iVmnoVR5MsQqk/oZJsnzdnGAq903lPaMILo
O64J+mMq0rZgp+1XRPjuQlDbkEbhUOPzFL+aQBuk1LG/KnUDwAgNWX5DJY7ylnhK
yQJQLWcXRgIKG/cprJ9LA5VeAS8WTno7gcgCY1vW03tDqBzzl/hbKqrdrmgrPbb8
u7Zurg0E3taC+9eYS0fUBinAgj6yNYPSDGQsJGE9PbXDwNf2gV1gTZghFpBmLMSv
Q9AHwaxSFbd61RG3xYQmlHmwYFd0gn1BdU6koF/PgZouaLHhosSp9jbvpRq7woEx
+0Fo+sUpdEGiJGzdjg9iarNHvZO8Ajztol6IkeB3ZmxclvjhToBvTzkjgZEaIvps
QfCQ1xH4Qzn8/RJ1M2MRC1h2F5efAwq4rBEflXfMYRRUeHCW9DzLTYpjeGHhwlHM
NDC99qPY1E3O5p8bgtkDXsiiC9XQ9nUj/p4/uxpEaxDXadLlYA7vJfM2zSioP2pu
u8ERhT3KyJHu7ks+mRKz5I4Je/JLO0cAhVF4zWCLMom24+2IPwoyK7lDBl8siNWM
1XthYZlIC/AdOFjniVovupTO6p9WDrinpvs2q69C0bBeiSgMaOgNU7R1Of5L2UhG
ElAs/ud/MyRCMgX3RyMsbeLpZQkxZoKWyqVysElhl/q+iEAHRFagNxmiUVaHN6l/
HcHCX/IElaEbOeIeyN+3EEcf1NfgJpDHk8HChXJROp2eRi8w1boDra6GPiQYzIwT
5KqbduuKaErBPbFiVeITcXtIZyMRLSUsbGSY5+iJg/iV+bjx5gg5ioqfJ+/NwZWK
UBKFp36eiDoNvQPBJyR4HeRsXWEMNMqei2QkoTDsLOBtvnOZX4ZU2pmcL9l2S95T
egFGmdkgZIgFCv6MUTs3u4W1XKY/rTAKjtcBzs8I57cntT1YcPL+XrJiVUb8BEUq
pJv3P8SNuzezpyVFyEIm9WOc2uV92OtpAQl/I695h7bfDzm0lywH1ZjM+Bza+bOi
b89fJ+HvFFBD29NBuHalrYv+aYC8drz+HguXzZvNppYqv6RiSTc3L3V7dGf6jd9I
Q6EdrQmyElabCOr34U5xOn58N0skE4l71eq2OYzEHx5jhPW8KVL7a834j6ai/X/s
VS1vq9bKurxDe7L/DMVWIFy4Tjb1fCJ3Etm1KLYDGwvxk5ZR5WmE6RWvLHHej4IA
eEGIrzFTl3bV/ayEFLv8PJakOQd7R9o9e9Eq4vPw6pageqxPUxQAi8zGwBn91w7M
8d/bMmnET6pfOPwKXt4JJo4DKnRB0MFnyP1/hWJjkQSDqs+2d2hNOHiriT7w3tuO
FPkSKq9m9vzr1Q9+4fYhuKLa2Vijg53cwD/mTl5yo0rcootBbLfd/jVj9Mp86CjP
FDPkzd1x+k0cAKD/LiWvAIOX1+c0x+pJ+rmIu5/V5HthqaaFs4ICXRJCIslAR5Xx
SmLdoNQIWWdrhMQ1+xk5pDXaq0Ve+U/0H2/PNpZSZcZEsCm9cVqPKpEUJi4jIZij
TucgY5xM05gUoRkxB1/NtUzp/eQQks32nsrbocJnPlnzMLjCANHjolXVNKarPahP
nb/e134XDNtnudn7URnZcmW0GPD2XCQIhbkSuw1cJvMNWLYQ/luiEOnGkpRCypXA
gZMTSRkZlHz3iGL/ZFn6R7j5Ofj4VIv2TR6BxCXlx3fgzjI7Z6Wbq8RjnLu3UT5p
y1vSFW90sh5PrrqpviS4An1rMwKuWSB5eF7F9EIZ+hImPIdN32kLs0EYxxm2FcWK
ZZRZWD8i0P5OnMDi/Do4aPMGsV/lXQdBVzv5ft8k10EZ4nuP0BPjX1wzJheTBmhL
qRmM9qBstWIuaWYx1Cb7P4QfWgK3KedlVfmqlp+pyQdXMfxQa1Pvs0/bystLiGa5
lVwAoHC7AOcJQfl/ma/fxAcSQkwekaRVoYeIFEJSlGoC6mQf/qbbStlO9Ya0YJTt
vj0/vSX9pJRoI2wQLU/0LpaiIxwvB9Q7vEFoIE5OrZas+B/NvkBqALvBZK2YdvWe
BowqNQ/Be8vr5klAqwD+njhtk0166fo8g0JOnEtjnGk+L0UxPxU5F4H5FMsDusPl
SXgBGOliWk3CpWBEjvRh294v3YGjKRFX6kS9OulUbKLyXa10vQp0kDs9QjmiF/2U
Zw/soyjcZOZ0kSn4LA6drK1u5bv6RZJWIpPIBddRRU46QHE5OF/xTuRITvd2z+Cv
5+y8pOsE4OJwHzkDe9QjyDmoiIaIa1kS1/WdWpRP9rZKyf2pO/knPWrpJpJ0Hwdn
pq+uPsOjjkDlB8FvA3v7aWbAJf2oPaoELVnbSMubAUoccfe88oY0JXZtx+iKGv1d
6sjS8Dn45sNpMTynNUioPi9uBb5ZBLopGQr/93KM4r4RImf8h4n4okaSyVYjEKoj
AZoH/kEi1qkbnKlGBVb4Nu2QtEQ2Y3P8T1BIe4izHA89IEtsWM2gAfpklyr66t5d
qLl4tBOmH3NsvYR5mp9wIMoWdPdml01Cbhk1Y1lKv1ii7QdLFgVavFmJLDcDmDf9
I+SXClddVMwzKkgCGA6WW8p6z9XQhEeEwV9uiSpZOtacZtxrascD3q+sxkSxrbn1
fHYKOP98K3eRZy7TI7TyXiMmGiYVEDHo4wrS8ClX+VkRtOuW/wLF7AlyZZYHNSDr
dr1x/676aT/Ff4jFZh2NoKvJnxk7Tl6jhoSgBAzSJEKaf8VJzF/J8RjQDqu7FXKq
H784+uWj7xuepKjz0svUQ/Y4v+4ca3DzYC0j4rOcSwlJfKewqPCPBEMM2BFZPJdZ
xAXa5IdmVBmb2Vq076ZtL966Kgd0rOnGazxazD0Y3VUqhVt5+zlhZCZeZov7DWsn
1/FsullJXxcr+xm7LmsXmJCBNp7ZnJa9/I7kNYaz8AHQlskeFmL2J0h2tPffkbc3
MXX0VeUxMZnzUCbxpAx0CPvQCQ7RHaVsWykR0x0o+e7JTfjCv4o84IRch1X445q2
JiM96TnWaiC07uPIokre+tSPY+DYy4jJtYMaAyyBCABTz3loJRNuz5dGyntd0CdH
sP8XFM8Jrz9X3hPzOiYQzeSp9nF1nQUHhC6wbjqX1pltKQEu3x1wk3L6kTKND+/s
741n/kQPRS+2oo56Wy2okv5pReha7RfycHphPS4KZoYId+V6aJ0dxqbLTapGBiLW
9NBC3i+wUZeA4Y7U9R2VnexyK2o/vDmX2VrepjpwknIdVXecVdjfCpv33hO7aS13
JwfVKRxXRylrCUMEQ3qhpkS8+H6mHW6KamPNXrdyDiFt1xpf6IgCPBBS1wfJXZCQ
iKjZ+nrvWwcp1QBfsak3v/hnkxXiroVqYgXVCupP5di+rciILpHTalTF9oLNzr43
7A/+6lA+3TwF+CHTVdbeq9Pi8xG87wpkFPvkm0+7nruFuvNqaMVsjATMEce59GIR
/IVB37mMP3teGybpUVbIReyAUb94+GzLJtiLHCR7H/DxvSGw2KPBjy/bpSN3+x4M
Epd1rlTqaNs+WApwZsW+8BXVamZ5w78boTHzHB4hMU3iAzLdNlCgn/wOJynJUpfA
hUDVLKCc5BLG5qmEAeka5tmdj8c4eSizfQMmwcApNqhi3flL0RCEgIPb1qSMYWh0
2v02tyJi2eg894VTfofx6WQqgzAC0CjpHH8WLAqpvq2x20qAdngF1wHDLvMasQYM
KSWJt3NtNgyubKR/XsFIICGTY+hDJGEDqGzHS0e1B2amzasj2gQXEYalNzNNCcw6
bbR7G6q21uUqa3lkBfxpFE9K0Uzd2/l/LDIkj9P0Roq+y8UOPx4yDdr1MNatdpHC
0ukRFLcBag9M7NvHc/NQ8Og1QDJ/B9E4rpS91AmLkY6eRxsfJ1BofEF3zQ3eBLMR
DxoFePYFWpVbOf2twNBTVNkje4RmWJnjZuypy1kpZb5V0nFRD7kmlO7aoou+ab8F
+oe0Maq12QSTawxbLhx+VLZjZWatjRnMWMyGyxfvtzqjI0LL8u3FgKsb1r0zXWJE
WQHeKFftn0j1oQE4ZEks4/ZuzbMBFCxooCZijrDfI/JfvRgoLzHrcJfglV1l3QML
irPJACo/50mOPror1AvDKWCFkmWD15Dx39wjEBljvMykCdKuoJ/gCuJ4cAwsIGMZ
m+j10vDWC9XA2IXylwxvdNA7w+srq6u16nQP8AXf+ijZqcQ2uZEydMgXZBPnf4OA
GKs/SLJQ+uTFbUPTcLXiAHOTghOzPcwdCzY1nE2t8/PP6QINjbfuy/A4x1hCfSDR
n9QHTd6tlx1g1VbFAf4GrSy00J202WjWBdAW6xAMwut2oLC+NFNYKLN90XDS4UAl
k6/yXYDPBeEIK2X2LyQopFAM0o9mdYf6kT+GdnFf0IJ9svlA1ZkPqSnWSFQIqoYp
v3p+MVGCs8X+kdN62Rui0qvZ2NypJR5bwRgnV+VfBlFJ5rtsllPL4cWbZkk4uIYJ
Bll3DsPn+/P8FtCEzZYYc0s0vwvtfittOCT9Z91c2XJOiax9Mz/IkXJ+4MshLMq9
fMURDxzgOD0wFIpQgfBb0Bb5ArRqUsKmzVG+GFxOPMem2NUh+I0OYSq1U1PrRIto
FEMzH0/+xL0HWshVRZzHbVGBOc5OK/zU58Jw7XkgoilwUGCInbY+E8ayLq1NX5qS
9CsjvbboloUDq3p+soHQkqLO5Akom5Z2ElxvjGTo7atMSOY5/KEjjSagOaLqNP8t
VQgUiTtFNGu3TnBpf1t2YcE4l9/+t7rqIhMic+UDMrB6qjhwYOFrcvV2bfmoMAOU
oCiftY0HcFmxWY1fZkIurCZAoJILNhhNHdV8Q9v6tMCbuSyR7DIJCZ4SIJ+QZPu9
a2qqzFxxSKe5zFYUapfd1LtNeEqtQRaKWpDkuLD8mtgl1bRoyl1rpbPdJQJYV11T
7ECbaJHV8E8054ETG9LDpnSAD/RKfbIV/aywoRZ+OYWLDgXeGuNLWELTWnL+WZq3
UY9gCVBbFbFkkXLsBjPqCgxxVb4lyAU1T1JktTWxWbUsyCj1YXSY09poH7yI4N5N
/zWaL9PctgrvnA2NYqwm6pVB/QJE9wGGxP4EONFTwKhdkefGcpNBfj3SWONBcRFL
EB39s+0l7ti4pqMbLhJuhxYn/55rVwmnc06tRlX8NWP3dZn5axltfcGThFm9+kZx
LwrhwTigwcjvnCyMixyyMF0zvWgHAM3VjMhyqTVSJxqFYXr3/etnR55IqIBDn84W
evefQEDaA5keLEQaNquHnarMuDLDIw8LPVtj8XFOoOrzPMTZ93unLCxVbQUfpr9W
8NpuUV4u3M7RipNxvf9HrZEY7eFYR5ROcNENiECHo5vKoMSBMJO44aMIgs/E1m7z
i62IbP5Wy5deTRq+PbNe/XZTGaYntgL8g1rCjzs4/IxLcmlSbn9UB3e4cVX83jx/
qbSdW3cI+cAEG6oNibw6Pe1wGXiiO6+WMJuYC4JSlb9IJpq6YS3zCF27h8c4vwLR
nt6a748jgBTAOM3N5VWAd7GDHY6W+mPitoeijdavh6MuQISA4VDCEUw7O213heeK
Ys2Uk1prC/K4FU7oI5kblaTwoIv8ipmfT9cGxvsiYgSiCMBKjXakquWOwTa2kZPJ
KvG++h6mUC7SKrLezNu0URBhEbhvJp9NQlODTyoEEp/hWn/UCSUZI9VANLfOyK/F
mb+xgqd919yOfifzqPLLsZh4K/IT1lNMmh7vQ4bnO1SGb3eAmUxmfyi/S5bZQbWv
He5Rjt8l5Hj2IvmOYVlESfYZYRYmWwUVvDOC1WLT1ncnlRFntXvXJs4eEL924NXx
/u2VyHSkfIEwk6vhMRQEiwAs4QtkyLpfIRqE+CyRVeW5nieWvn/u+xnLrDnDL4BJ
IFCGk2kpygehmmTgaRMdoKTFB9zSTYMY1SHczVZldJshpFyS8RXU5oHqMnAR7/fL
YL87X8PPk+P2/pwFgqZM1OuzlQ185YuIc0bfHNbwcRZT3FUKprKoisCQvIJvgYVw
InpvAKHCwvSgKgAEGJG/LCQD5Y7/eu9o4m1RTs56EGDPO7dYnsDJD76KpAvMJ6G5
l7DnUVPZpd8P/rR2FdBCm44aZNr/FIb8EJSbfMHsSMPzuH/hDHN5b1nZEjwOo9tF
WuUpofiSZc2YBugwSDpBbevuyaeKV/rS+wm3aGQwIr6k2+havAuvyiF6VWTKdGHC
wNa9WtCh/x0A+EgZKdM+/oU6iotFm/81hDlsH6qVuw3mNJm1p4SpNzd/sAzxLYPM
5bZXcnCB1i25bQTaI51fSIHoX3yMJPeQ7UD/1Zh+WW55uK+riWGeYyps3fuM157w
A557AO+0BWAj8BV3CE0SfTJ28T6bn69IqEdUvzp6WOF1a0JORFUjER6b+EHlFIue
XKEQ08S7j5awY/tvl+MmHU//njmUtshc11/nv7+oDxut//DWRpPNIKHnoKRZJL2y
Q9HbpcK34EvrbQoS8Kx61tzxOdjgYXWytG3TkpjQLI+pdiLMozaYC3Wc1m68rbA/
PdTPWhC/Bn5FynnIuD0yW2PbKArcQDaTUsN/qJ+RfKayxqssO4NBKrYDsnfMpAKt
w5fuveqadjHS9KAakeHh1Xvl+3Mncl4Y9gn+2Roz7Uq+OUkzLARkh0p4fGmh7SZf
z38Y8Jx74yy4On0Dtg3OP882za7TeILvKy1lG1d9wqlwVMplPx/PVeMxzJvSYmt3
g5V93/LOsEqnjHBcRvKsA58+05tU5Kx7Uot91rSHEChsmPi0o5+I0113V5eVXu3f
nuQUKwLXnJrE2FgZOBLxctNhwJjfE1IhiCS/mVtT0qMkQSd7FloHqtlibU40F6Q0
/vEM1sZQ2wFBjJrQi/3s/bS0jCinvSEUJlHcOt4drPZ9GaAG5CjMEsf+HHTDbvz5
MIfe1Slzlo/0TscboLJw5LgLGsLHolVcG2F4lLV/ghurnrJXJcPw44qUEUqH3hZE
7x75jATowCbjMfWeAXivgMLCJtmB7WcSZbyc6qCyGPwGnuB3iJtL9OZQaUvQPxUi
dZxrunnOxUhJZyYZjVEB9BsGUifHcQ98SEFM0FHDD3OZlRqQg/JB7G4eOTDj1DNm
X0mHnu09EHPVgiEGFS/s2KAiRDMHgCeaHJaZg6NRGHRdVrtIHdsps0zy9bfUunUI
A9h/520obkS2cIKYhFSxYL8a1MF5GYZ0d0aNOib25v3Ea8f9GYB3NdWRdSWWgjgA
EukRuJoBe5lDJXwkkOH/WcXiDiHEglj8rpf4WgCAQ897LODLcfjLCvxryS2+eDiP
YrPI8bNsnsE/OBZUKpjXaLVa/+yI90CRtOHJYEa7u8/ZDJL8D6Xqb/vxKE9hxI6m
OXm4OnaEYeWmwbb9qVGuNkB5MkvRjD3ERNZEyMpsT3qrGUibzJHIDvl2tOMzz18c
PSMg38wnOSTH6wiuWHgywJB74KSYO3Nr1jUjU0HozpjS6UMBXZDVz3Kat+jyQwDy
pnyG3DHxMq1VC7IBDeyKq2f1ogDQ7v9Pqsfew3UkjzGM5uSjBFUIU1+/55AOliaT
vMAYM9gK16IQ/zjmA1YRp8pcz7pv1RrXfHSj3HhR3pTFiLzcxbmb6y5umWKaOVGx
41QgfLkihOVMlof02UwUczdc8J2V81bEDlVNDH305bFxFj6gkmOJ7v7i3pTHOwuz
dSGHpgM15gV8YHgjrHelVlLFXdnW5PvLCZf1SYg1lzTEmDS6p0Qm9lT/0tEI5A4X
uPPxzfMeapCBG7e+t5VutcF+sxyVCb4ruQj2druCOYF6cbLayKcoFjfxZ3qKSPmS
7sNwcueYn5hzfS4BkawAI9npYZhPnEJMtcogGofdAIM2FK4T72aoznKTcprgXZD5
QxEBESzOCqrknVzDkBtiQ4qrIJTznJ7e5uZU3uuSCce5zAHd3IC765pDC8gGKRIp
+2aE/AKBqhNtDuytbQ0KtpsXVUjk3AiwmBGMxgE/vQ5OgWo5fk7tltrAmPp9U9ln
VNLncMSRtGq32p985CSymU6KZcaJxz9Nw6FkeRsAHnV61jAGaB95lzpbQlTQJB2a
4Z4tGbzWGKDMh0XIex0dn9nusaTiqcaW13R0h3xRdDgVIH2ijmey2yuLewnbLwV6
1AYvCBiBCqLx35we4ct7VPAavIy8qPuO3LH0rubTc05FZ4rAMV9NxJpNyia7syhH
5Dw9HTGbdbqmBKepeKvxtTq8btfKNhhLbZ0pTF4O+0j1zuuAm0hVfUSj5dyQBe7Y
UJkAZdeMkzLTd/pT1DtnUb+0mSSCu12wygAUMYZHTzwLdO5EpOn+ErBr6Pa2dbp5
a/U+QcOeESmdSZPbTVPLlSKZh1wd+MLsQmZ7ruZv3jlTtdHAhLFGnplryjbdHkZM
pZCgG8aKEa2BGHYcEBi7sf8O8JuD9mOZ9DuEI3qtCMxT4X147nKRFu/3E8OD4kQ4
S6qci+CdG6IsMeCq2pXr4CEozk85CZmr5EFOCcQHkb/sSZIvYHXCmRCTHlEPfH+8
P2IIn6hYqwwcgX1yhI7hWbZ5WxzUkbyVKQxF/1SN06wwflj6xmiEetibbZNL59Td
lBi5kmXJ9zmq8KARsE4aMTFRLlrdO0eYCFGYC72RQePPwjptCiJNEBc6q6kV5ygE
Y4wp7P/nwJf4Qu2NJucSQ4ukiywyRYSULAY9uaFLgbLT8bVG+e9xoaTOZ0QT/3sn
1LpiM+Un6OxCVWB9i+IkHlr7QQRat3afmUB9FxrXyDGbjKgT1Qdjmu48O514MP0u
6FcbsdrmtzKnsHj3PKehDx5LHJpjq0IW7+0/NZmWog/Y4xoSHnmmOJr1p9Qfh7Ny
yKdP0OuO6EgZH07UMO818/1wvsMNy7lIYnTEgt/5oUIat3gZ//f6pfZN2VWO8ptl
+drNzuesUSzY3L0jgGHhNjGJRJI9LRmdEDaHcs8JafvZoOEGFIqKobn/5vZuA3Q/
WRWECzNp7slWU1Vobc7LeQKm9bji/lSqvNOar1i0V68rOYNSq4jmrsEo1YJRSlA0
dFx3PzMw8QmYhP8h71ZxGfOgPCx0O8w4wnNea5NOvMDczgQAP2WHVcaG2OZcAg/9
Bc/fEMbyr67PaHtrI3uYarJOD2zEklJFcamZzXSKfoZSuxDkyswZP2Leqj0zpzli
PzJsWG7otkiCzXzQ8b5RfbqZJr+NQBB4qvGS0S+ypKoRi8XwxvosiPZFNbP/kA3n
ryAdfgQP8WSCim3U5p13ljG0qdJcqPNAbVzzkSQUQyiIp0gJJIW3at7n5U1UUdpJ
RgPLiXamsuFcsDg/9EWyrp6ijppOgBup3TBLIdeV+9O8sDq/OYJPqWDO+ocpt3Tr
Lj8Lxi4Uiq/xaal3+O/stETtHmeJXn3bqg5/UQvmOVcVdtO1HoVndC6tQG8/muL3
X46f60sZVdaR/rWnqBzdW2MiEkN1iY+aa3EnIkOJ+8kwQuroSwj+xiXEutGK19bK
GJpHAgQgCpggCFj0wWTSudh7txNr6RogUVCHIo/Cki4gBG1QamTW0ATuYiBOMRTO
zAi7O/+uKYlqtnjti7riOgEdlqj+w4a97hpX1eqS707C4S22CO6dorFjaF27mFlf
Udsyn2rObaHgid4pxe3ugXSMgFTVAQarXoAkHWW67/bBnn59iEsN6QiLT4JhyH5S
dxtdxU6tGPFpKPJS7zCbSzY4k5wM9E2HaEov06+B2B2VGut+UcuP/zyj5E891t2+
r6z9fmL7RuDVRiWHF6+fkngCu/UMJTvgI0sCQTZkYSrrzUW929RHn4pKP4YBFz6Z
d1qznPwiLHQjm4btwPv0vxB8SB2lB4WFlgD/2H63XoROidpgRQ3Ka4LVqewDDwEo
t8gqbX5Zq9bX7FOfsywlvM9QHs1FfFX0ImhkFERIbarMJde08e0ks8ISey7G3kDi
lNuBKauNGfzEodfztjpMyH1nkpCZRQxqgm+G/NBmhO66UY6B0izavD+djqStohKT
U/ZArvkWwySBkmS1dT9tpnjEsF+88dYrpZtRYs/7ohyTs5Ys4LgqZ2FOHh4sdde1
VjScjmRHb2MKGKZ7e0xs/TkOqKnsoMaD+Er+WCe2PkanV/5SEKIpURiDhUgfoGRF
Bc3qidZIFALq3LTnPj3Xohj5roU/A+gqFaCwB9SJxdlFtds9Y2QOBdS2OXeFpyjp
aOe7bv+0ckPRg0nS27afTnJP9G1pg7jnb3V+HPA7wcc3aaGQ470XvvYQMyv0XDzZ
7ZveZv7xyYfXhfcxPtJu3SnInEZ/8Jv9ZggL7dg/PGAkdnzxL+H//aI1bukOtZ3o
xq+7HGeAuo+efpsVyqbf4G7/mdJS1f33KT7gGh/JT3aMjHeRzAN4ei/0lZp0yvGi
hYnueQJUL0R+vy0Pc0nxHIf3XzaMaFU31sVzW5mF7fCgohnM6felBtkeY8GsY6nA
TgB/ZX6K74xDE9VrV4hG9DhBVOIYvr4aoQgK0x7Y0hsBAGFmqsuUiHjDwExCqwYz
XNIoxJaBo5tvKzCt3S/Obe5FZf+igOJ/IK6C7MYihXcZe1LcJxowKOMbaUxeA/pZ
PDfyby3FsROTSrMeZXNCT0MDSoNgUZUAoMYy7Hby8lpeNO5cbtFxpNbrcPp6HMm6
M0FAA/AySHwPMprdCAvVL7j9Hn5k17cb4lFp1wKzga2GuAzVRcp/7j2uX3ZyQbZz
k8kFNXo4rtR5QZNWRgUb8hSC1eJHyAQfiswaquvsCzspwvguB3OzuJwKE5W0xk7l
W+FIdwzCn+ybwpl1JNBBo+X8F8y7HVS7y5c0TgmJrUUEpLvsaTAK+DnMKzCPrO5F
+Ojp1qyYyeYk+2FdcgJhJEEcXIGcfeOJA34xT/0UUwNkF6mLLYDrndGI7s/rQYQL
vtLV8K7PziA4aEh1fNq7RdF+K8PQpBQ28zG+WL8wI7HNk8qtCDNoc8/a2Tv9OU2A
z0ZltzEKcu23vldwGEIy5uqTOV1fscxDUN29eIXOmhAj+ubMRHGm2L0Y4nv+JAq7
zVyWDdKdb+oVwAcAnKKAtBohBka7CXdrxtQZWOFUsLA91MXQBnse3zxPsR8A91SZ
w9jOFnd6VN7aaXkkLzCbfyAkJVndRtr7M65BEyAUSqhuIl/yezmik8PhluYoDlmc
hRfk0F+Z60hrP0bNV1pdmQuwTj/GV9YBC/x2P1fSpmcR3yQdOnAjX1BXrDyP6N5v
DCKrnFUGfLdnPePFLuJN3Qd5IqjFuMCxRF9YsOg5G690IzmBGH7ff5Pcn05bXM4i
5NqaOlGJxQxpFAUkMW5Ad/wIo+nrtJvtotPXa3UJQdt1e27BGP2G2gMqjg9TD9XO
Ij6nsemnr1qtoqo2vISUO5UuX35lFC8pgkq+AC4TwHmPQovQys0B5eqaBIpSzo6+
7hG11SwK02xuDRBUvzuHVGJoOW8PyPMB+cosZe6tnEf1Ym2Qs4ejZN6Rc5Y0jmhC
efllXiCyg5Akog4/Mvqjuz+g4abDZJVQuzFhMuis1tuHUd9q0mpSqqJuBRyp9Gi3
u82FV0CkuXkGF1fvhbdjWa0xY6kRbTXsqswh0JJw1kNo9wcdg5dy9wMAd3YVedku
eJXtcTUbD8hP0aFNlC+X9Ofzf1C5qJSiP5AIF4CvWOlLH8TLa4LYcl6SrIxNqaUa
0Yx+lyQX3eToK9dSF+IXIMsn4YDum6LaDEKNAZSQykahDtEpC+gIPjTMnscRv09d
Fh/kUckemZLCrpw50BOFrLChnu6eYAlbGuLoxuzmQja0NavWGGAM3XAe9qsZgvVT
5kffSOZl9bx+R0a3b5ZwxQTbcXFbmqTZ2w9jRU4GjaYCxHSDupDVd+lSGfcyYAIb
XlkbQ72MtMVPTxqM5WLKTjY37Ay63HFNUOpciVfBGB+GRMxNO9caM+AGGocSAKoJ
w653DZVwuVVpb5a4N/DwDEC0VzaUUda9Or1jElFguMR9/WwX69E3FNZdm3tCEVbl
/A35f/AZmc9uOGMmdjimmxpAMuFXu0CBlHXLoHAaB3+AfrOacTKgE2a0WDjW6FqS
gIxSKtmVLFZPmShE/aLy220cbIyHtratMXwg0RTOzMZlQezNcNxDQeCd+2pVia+0
Qov4+w5mE/sY0DB8aNdF3UcZtBJ1L+9ELB8Xwy6XwhGXFS1cZ43mI+7bw2EEGzIK
qsqkyTlR0KUCTYYvZvdNocCxnQHLa4YzdvCiFKzkE3uQURcJXVhjRsOkTiVBTGfw
vD+udB/AlcWkLBPd59nqlu4Xp9un2jmrjLhaB82EvI/KgDQT+2ZFJ8wVxYmvHKG2
z0WRb1x6ubR4gnIaHC91pAn8e5smre2MQQoodFZAIsKcMx0uijeup3EnRf8OEEE4
22roXMwh+B38Xru8l754UlLIF6gAfPEVwgsWs7yugYYsTYjG4UXdVC6xwHalzaBb
RczqmFnhTUZaaAURn6qAuYSwnB5w4cC4k3r9Ct+V0nkypT9s5yot8DTnZlm/Ou3T
/yUHZcMK4lUj4Lrufg6D7FqTaj1vA1LIzN1Ebhxd4fuOEM9vYD5sB2kmODuYdo6B
5wpC5AiWYAMXa5KtqqhIeyXda9izEaVHGAEJ9h4mbz7Pn8zQjpzXC5qP4tTZ6NYY
+sXGdRbuZ1yhr6v4ljQcsupnPxxElXAMe0VhAc1ofj0UNjKqEAU0ClCNHu76Cqb9
aNm/E4ir7/gaNAs5sDaAu/I+SUkcqs2GgxSOMvctgI1UUwBffTvRNJoroydgpjO4
C/JEB+KAbMTk823iQzJLQzR7A205viiBnE3kcxaBCC7vmzRjtDFkWPGUuieKqCx9
nYR5VFF/ssrbcp5GmM0mYXfi425XMy1BSKpCgl0i7egTBo14Uv0nuiL2myoc9xke
2jiwbmAnSYAfd0C02DDnZR+HZvVsfLCQ4Bfuz9BMwltYtRR5oFxpSHNwKAwBgpL4
d1fUjVmvq1+SrTNm5TkUA9d2QvLbeiZkyGNu0cwQ61u+4Ic4Pd+rnDgBUrmJwoAR
/7W3YBiUFOv4QJJbT0FLvYUmQFSxhqrVyAklWXmMx622/a8w2yjajm1acixkiE18
tZBXc4h8G5ITrOWWC90F2WpY413jo1pw1VbCtBDWu1gHxQoxIW2ubpNMixn12F+c
UM3lkw50vM44blbkDAkKR6O1lM/MEDIyjfYI8LKqkC7w6sKyxLLwQrpa/ainsm4G
hNKwAn2Tkga27zMAwCPeZEkVNH3VwkuKfC8bc9hpsuqLi52hpGx4HFzMMae9PAyB
xFTPRQXpuXrDOGEVAoakQNPeqQTTyBwLqwySU546NljtvsDlyeu8IsVkAI4weRTX
OzULSYZvzmnaSgAd0tsDM6G80+PT6mxwg/u+DzhIaHtlhy1NPRhKW703wmqIjiNS
mvtl5JIwIe80bhs3f8q6TKTIhA84Y98+sy2n3SC++IPAP8sZLFAvXTbJTfVUFYPx
mZbFuxaVcr4ybZqO43h7gNSgHzXBOrE5DqDjgbdclxg1na/Q1Y/R5abv6dMmcj9p
zFoJBNx5LpVdnEP1FxlMOqnsp3Xk0ACTVMHNwjSX67dzXXBfPwSkeG6vVqPrUFeL
RnjAEPI0iIqaCph0yIK7eVS5Kqrqx/5g/SlV0xkVNCJ0ybv/pi6yQGr5gWVQOhX5
J90t7fcs+UCzfpZpKAFqXvNL0cjV9p8oV/3F5Z58+Jx7TJBVYlGJbM9HV1gSUitf
k7ln+23gPQqaxqTtu5FcoEHlGSaF4cafjTtx0I72qMUXURyDaw1WEmE8uXoUGBGi
UIzyMPf0dWalv0akJK2J/4ii6VCmzR70RqdyALCoN19zVh8nWeH3ILmQ5vMyOyOI
xv5GGhpNCMl5Mat4hJclGnPmUaeN7Rv0gGe+DlAtSEKPPB3kh9p7B11ZFmiOUu1Z
0JJP/mNcc9zjVrxSrdYm0dStSxE7OW3Y3XFmHipgj3k+Ug+MiljOaDM9zibTP+7F
iFOivh7XWu6I0JqEqTo31MaUHd+FrkenK2FQSelcdxcJa8wnSr5VwFbque5NKie4
v6YwpAnHHH8uvLxsecmAikptQ0yd21O01NbS865B3E+bAOILQ/Jt/KurSUxZJ+f6
RV8Tc/OMsNKpiTJmXx0bunZj3lz9h8Lsl3ctcwyc4cNv+ybBTf6a16SG1NinHNks
59Sqfxioc6T2Esu1pUD7oHpqJZ8wCEt8kWVYCNycW2XnBpa2LuTK0FzgOoXaiOYL
9sFvW6xKxcokIgz9Y6yMlAExv1mv77xQGGBkjS/iQ/OhIVoVtbUyFkn/lFtPhlKG
pvYo+gxSvZbfJ9d8JAzjzOlWLSLf++em6HZy45JqeFx+FLgpQLOyd0afdVujJnUw
JmYODAXcnVYNf4Q+MdMKX+CPJZnccUAPD/JeZJaFeIs9TNxtjD2wF0wqPL0eCYs9
02CveiRnDanTr/cubTN8gmVHf2fVY1218XPSjLZvMrDkjcT0ymmTCV2Dqd/Y+ewa
WJLDAn+l3qIxaFwnRkkFjuwspelPuRouLWNl34yOoQH5PvCbGMq5D0qE4/N6kU7o
A9iyOjBkkoo9CMN4lYMAwwxtdUdFxjw10TyQvgxZpuRHE9o4ctFRIJGX7aOhoqgc
nJgwJ3SPnxvrvwZvLdrTAwtRn8te2e0pEeC46+RMyNTxqP2KRC4TE3oHY+Vo2E33
AvwjSuJAILB8+wcdRsfWyrKwP3txA/lICF1Mw3o0BFIJkjEKoMXsGXghEzvL6BsX
zgYpvE6sNJ21Wqe0VLovYwMoXECTHyYfLGV/o/H1ksGPgBvF7Z5fXQETGO7m1syH
q0xClJZnD+iQBEyrmfsSmlmf2DipQVjvpqsxzwEfWaMujhRyumrB+St8bj/yfZs5
75QdSQteSkbHUZZ5Ag1RdhgtiZP/hCU1poJ2PO1muTZWfWTXL1zPBOspjmeHEfwq
d2r+UvYHo6PLLGvXj6QFhuKC6sbduEUhVwltDJAb/sgq0KThWfNlE8xqTHKQA6+k
eRp+6ipBnLxAllsnl0UdFq0AxgZslZR19CAzFjVr7YCJ98YQGPLiuq1F5fwKl0xo
QHjVdLi4WD+eLjr9GzZc9r+VNxevzF/u1xoWmLEwnv4mWdfGjqZvRRPxonyOsbSZ
oMdr6oZptQd5KEs8/YSRQrUPlHO6jf2gW5Sq2JsSwaabJjPUvZqzUyZ/+vvE6wIs
BSp/E+XKyEpA23hcZasKWO8hT5lphEEVYSqJC0ZRKtjKa1KghHEBPa/utRrgFxnf
Jk5lB6cOYuumr7CoMCU2y/QGNbYJnPfbZ5E/DM4kT5eCzn/+h1JnFuQnDFNFWS3c
ychPHPI/xQVlmla/ebDdg9bPZZ/bXmRgxqUkd3bLdsJdaezZIcmzXKkWIjtIMeb8
oHfuY4FZL9DT4o3pihs2CRcO8W6unAuC8FFhZkOiHvFmlT03Ms1Vkf9lsVAcUGG2
Nd1saRlGOxhscXxU1oxSS77HK5s0olSeR4QtWyVYjQGYCM4iFQmOhijNR8nUxg4Z
23CeApGPn3qJ1EnXvFtdhpLCtb8trFRCPUbo5egVkoPjhgGw/DfjzBySSwRPTb2S
di4WxvA4BsP1TRWUsNzYdYwWO2Lsd0M/kl46CGoxl7eqcKmBjF/r6N4Hy+3fkapW
93yfu1Wv2oih5JDa3qE9x4Qx+BvkvBhCqHExa2BCwPoZoCvN2tPLLHIHH8N8Evt3
/FTsR38Jpndu1NMN3TRNLCpNoB1MS/OW2nX8Ao/4Eoqql9Ouso1nrXCn0mBo1xp0
1zoXLo/4jOtzuKKubpPoF6ugVMgoHnuNZ6ivG5mf72gXCo4Yi1lNk9wh40045TcQ
SXeipp0OFrIt+x3cEQFwEEsp2XXaxGpwT/wLBfnLLYpgaa6vwrVeFd7ePRSjt0Sh
tV5Px3JRlMUa5tFHPFDodu8WYnkd5MyPWZH3q9UrL8O4MbWZPtvDDkFgvbxEg52h
Tkm/sCwqaDFYT2y9iNNDJT0mN5xg9xLWXNBYZXJvjNP0Ev5TiMHDIYhvwG5td0ym
CO9RK36LEHUf4Ge80fYag9hN5xu0v9tC8QtLnzH+/7MRIQrQ51rZNHPOaKjS16DP
3uPu9UOcsL7O/UMydZYrfjH3APrg9pIlVI6vjPBdVSc/J6thiwy74JDAXRHW0i4q
sQJbOtYVyHb8hbgok2H84r+XOR6tSmn+0Z6F4Q20ee5fwPmiwDVwTmQD2+v1Jwab
o691oklaHKZ/pBxmrHHBv7WLI04G00d8qnUuGq/hOtAq4KmiWDr4dirF9YWBj6EV
RUP+YE5q0IAhRr7OdWrrYBZy5M/KaJ/UNiQhl7Ksf4zQ0lPlKloXT5Z0S1LzC8Rs
teoYBCPxbCPImdPCdRRiI0pKV63PKhlF2XO0xE6FI4Ca67CUQ6cQPC9HXHq0jxPD
/k6fAHYemoATK/V2aM3OLbkmWwUn4GrP6WtLt9+fVIDdFGSsPU1x3IVbDxQ1uL7d
47Zq5W2Qw0R3ZIFYghyPEn6yOonDi8oNOrdvFVXK5wczSAo2z22aEGos9aA2n2IN
B0xlzdVVHP8CAWa2GyOumzoKfbrSq0jY4oDEF5QfJhMu5zbyS3609EL1MX2IaN2K
cyrDV/OehjP1YG8epY3jvYDGWrNbZONEuO5vSZqKeGvwRb190glfNrx5twTIJ2sL
QFJSFhvpvcTmM1N6Xhz/jLyiRlrkt2gPBc7nqrSDmrw6eK2phOzZ8amBzjskABu+
TJPRrCRqPa9mXPEldKWdWnxzsI1p155vdTqf2UV20FKFwadOKqHTFco7elQJTUKC
rbM2MvFxjFgtxZhKeBVdW/1s+8Tqy+25zX1gLJSThonRmg0OaD5pJJBPjBh2f09h
L6GVt8jjOTnuig03oYAePXgd3NxdcCYiflzE/S95pLx3GBQQ03N59uLwzwxPBzgS
It724HuCn8sRYfMs02KCCb+4zTtmpOOMQQOzpA3WA60eKW77Z07tNym0IdargqCy
ftgxJO3Ecfrv/VHu5nvldsVo6dwdxrh3vEGcBK/yfuyHqJGMXZoxtMqWvcyDjnlV
7sxhL1Tu0j2h0IZVZylj0CQmgIbUN67mOBUNIxUMOzrHamE+PjQpfT1RsoYP4CYr
vtBU0aXeyiGsnie5vaM/gpymn4dUoHJqD/0+9z/XkygKBeNK91VaMb5Q0zz0juKX
/vIPtL6BT1lB4AlauDChr/0jH79y3bany//2XIK26AUrieWlZ+yPso1BfV87sE+u
xyzwLl0w4++okOZmNrqL8nlgMGoaJv9OvkgLkwmuRYcssFGcuqc3a2gTucPiMjAp
1r5Y1O1y9T+9Vbpx5HqK1lMyFLQ8MuD9nuaFCprjkfdQexlCas4qJ532TKabzSzo
RrqerWVttw0P0WqvoqRdcDBXVT/zF5LYto+Uxa4BjJEjTqWXfWBEw430E4t+67HO
yrKUg8+nP0PKBxWentGMdy2JQGTtyws/f+0cIu1ZmvfQnVCCISwKZbLwI8rXJxMk
WhSQt3psALntLKxLK7IaklKgFO9jF4FwIl5U6xg5EaKoItUEZFfBJToTbJ0vlcbn
4DUINIP6Yj90tEkRpn3Uj0qXn8C4QWOmDxjnr2jzVhSb0oua1VcYkTbfJF9rdIB5
AXofZRuhAQ+gSmpvx+8cO2qZsVC+cl0kO9LgnQYQEs7f3sTV/BUz4oiOboDhtpE6
s5bTmEYB25grk+NQ7kkFPgNkOVt+ApN0h7JiTqqw845HBD9LQEdzf8k+AB9DviYu
oZvnzW0J0sDqILIOV/nP69oaYImbHz4+t9IIylQ9B2yq1nqY8Q1xgA4ICRxM+46m
K7YAceW7oJBxqK9zeD7b/MBzgnoeSY0bDcEauTAmRwVngf+zFPtVNxi2pKMvzDbT
0xA75SK9HVYMZbappgizwyJyUsSnxP56uN0YT3E+ljIssfA7ixtL3F+oLoFFRaaj
9WLggVqBREKvEnO2nunlDWPbfWEe1Qlk5BLnuHUCI8nY9aNZaNDrm3cdzsCtuM8I
Z4oWYhJL5zGOSBJyQzCEpLBqedEZU5hBS4+ADmD9P2hhZ6qAnlkbf6FNxJGG05oQ
TzSmEPLBAhsjRzFg6z3J3FBAmeFAn5vvpg2jpnauZKKaqRX86ubrRS2Qp/wrm8jK
K/4ip8XYoqGHZSB/aVZq6TJTmb/iFRtuHuEHyzv92sX+KAsCwgjHaRVEuUuDln2Z
ePWDXl5ojH2L43yeQIyBdHdFPhfTOBIkdc3wzor9E3pu4RX+BEocYp4tBay09MoR
g2Lb7W+kTKcbyth+UjrpiAisFgGRy9Q51HAKgFOprXnRGgpMRVQxvPuKC74rNXk3
Pqg4r6GVDyZ/2u3cB0lAlPavck3cYYMXz0lnLK1tA25bRBqP4El+oXT52me2WMdS
eubU8avHl2SaWrCdzB/dDJbhQD1sGqjAk3P6XVqpXFemVoMon6j+z76W4K+hxAnT
nKDO/bdtctsoJyqe+0xgjMFHff1Z7hi8Uy/sHvdgP6CXYyqtuQx/D26Cp/ikAk8Z
tNFFGZccpxRXsQSoth5x0y9ODjhqj+AGSdw4g3aHVnBd0neIgQWKuYnIieYt4cK/
28GXnF+p0XTo2id51rXw6NDFUCxINeqmZ0MPwiN4510suar8W46iPcbm7Qpgqy5p
TZDO7j2FxA6fodJyCTMHX6unCSU1N0JhErKOELlLpYvOTJA6yFTfHng0xFgcG9Ht
Y6c2pDjD3bhXnVIdzRFMyXQe3Ge1ekqsAoSnXJGuf51NqpDC8OWLXAvMelBr1+tw
DJ4KC+1r6MxQWHqNB6XQpxT6A2DbMl26RG9eNWAiIANSUgxzHU2TBKfNMTBcJ8Ve
+bpNlwWpzm61OZ7SFpytOz7ydXRcV4ycdD16gAOjOOGGIYrKvCUQ0lqDN9wFXbu0
nB0NntCIgdQTLikRHdfpzADkVpHa/sxe2pIQg2l1znig5FDxLNUT7TUCcVayltr8
fZbhLjaEJJoe0A71nvAaIb07VTDUFYwpXG84m8YBXDoXb6FQN6tjNxD3ta8I5mU8
EiFTYx+Bppqx3KRY6gEc4VPoFaVOzM1QbbYrrZ05vCLHaXHXlav0KpFK806ZFugP
hyDDPDnE4UV0ezrx3Q7L0088M0zuzCfpztqPQjuW3CEriClegdVcDh0gPRa8atQV
/wMu7L03/ZmgHC6C0ljb285SVBkCKVIGgMpoOEQ5U1gviWQll65yveQ7W8PxArU2
ESoj1hQeyVLoLjifCwB6TEKydw10Zfe7D/6lgPN5RJ2R3kLFoGqz7wSuWM/h3Zkr
i5rJ2WHl/n4GvApq2spk2DNgespzGAR4zJlvK3D6njMucNFuVi8no+mZ1TbloaX0
apJ22JEbw0gGBVMMAYUhjWVW5DFiDQFlfuUfRiVQPXijlIXk9rW2tgEmG3SuuORr
NPy2deSEinVMEEQ7OC08XqkUdvzo1hDb2LAEzwLaqT9Ut4JLN5VyY1VEe47lkTEE
fW3JaSNDjtykaWaJm2rNT0O68Td4tYkpX0XUPjlUXEoOmXqH5DoWIrrvaEd6ctOQ
+rIcxCKh0HWp+af+2Onl0s1b2cxFrN6p9wjaE0Aub6kIxPvZhkUjhm4xFR+eh/68
qFj+NB9mQBh6xPQZTrffLQfJ5pxawLS7X7QTrAfwkWMuz3lviljGs8IHCwdA9+zv
wz4lR4KOcmIaQDRcKJvMs0/gQQVExG/Lvh28i+AVJOWHyoQA6FLCLhqmAum7Vl0M
m+eVOBe4TI3J070Ruvqhwei2FHqS8yRw33nHDU7zjaIG+wQ5KtAWzeY8hrmZlYkU
dd8/jCHdAtsgkzwUm5xkUaj9kGdBDXC8aiZBVfnKM80N3xScl4VC9K0KzatUoEOt
0kGu6wNKAeHnTX+idp2ekaQkvPs35Cp3XgZ8qTer2K6DonihFtEL/DFA4QPczmjt
3nsvY8aDHNLrRoTTlSyHL0uw3aTuzE77eqI3Ti2GlbQICPl1CV1peyC7X2bIdTRi
PhuBxjmYyCD5u/SlQpEqFLTDgNOJClfOeLAN054gcSuts2wF7xkl3lSvKv5UbdsC
z/pgIxSSVIYWan3oIWXUAJX1gKUekjrAjfoaqUqB3Hpkbpg38I6jcNj/ndc51KPq
wCIEb0DmXs6yvgLlZxdRP48ChiW7A0S1aGN89Nzq/597HiZPji+P15KKjw2sFMvc
oU9HV4mDogCJU7GFGcfu/tCdOEUbSsTtNA8b2HxUHdXfl3OfmUdh11MtlWg1AOv0
gZJqmn0ZJ2KkXPMm8bbktjS5K2h9oKv+Ie2OfwVdBC+tUF0F3UpwZXcfOV45Gzna
9tSpofI/lZArXbceoiXr1ju4wkz9p6JkxMROGIsY6WiWIysFNNd+5xBPTJ8klZtj
KpPe0zMc1Fw6ifSNxpxh3bkd4vm0t7kY1lJxBRBG+61A1Eo0xzg6W9IjPcvVUCHK
9DubzO53EmYgipqUXLZ2bqIzKSunneTjqthG4UEGeFPwJY3HxwRzZqVZoxPqNJlM
GMHdmozR4AxBgdx9n4F7HBMt99c/jGcnJ4Et5TTW19GEf+/BqV/PXcVIngyKe7QR
3Gk82YeBICHZb4Bnv9shuO2n2Z/OeBoE9PY7XLirF3XRdz9Vy05sZP1rMVPCOji5
r34RW7gDKtR19XJJtDQIfT/smweQ5A4RdgkplR/OQBaktQZRpKoCP3ip03gKeYrm
dQoDotOJc8ObWrsxd4FuOA4nyt2dqXzlQF7tYJFa56qBa+nBgfhj5L16Cn9KMPeB
y33wgiPxdBjq3z9kBZHTt1iJDYF2hZD8BrFP02S88AyOSjPfu6bbszZ7b3mzKw49
ULoZTE96v9IcaFcGQi6zbVsvDsnJIHmRXAgaq2C9RJjd//wJ9n6RhDu5GE9DgXhS
ZihDXso42PPAp9rioPEmbnsN8Yd8W5dQf63sgEtDv14ce1xPeOBlNZN+Ja0swGXT
YlaI3zY+/khFto/NT13wZtxkfBp8mw1Q1SQajDl+bzA8/QBfV5c0HbjQtf+Smeks
DqoZSx47i2ifL6vrt6CQnQU2mS8KbeF4I8BnVe2jT428fkp78Aan1NAtkY6wsd35
ZGH8VO/ybiolf+MHpG+0JtQBMmGbpueDA5cvcCa5Sm7vQZTDKZElD4KK7FWw94XR
Mo+g7F/ouvJ+/WsPkLVzgNlgAjySSCGyJ7vIatfZMRla6eSW1Jp9xArA/f1YC5pR
rDLES23Q6ZPaUGjjT8UDmPqv1No6KfSWiNu1kBAlpJFYihKtM5xXX+RF+kOzKEHy
lLZckHiulDuHV5JkePjgWCl0ToREiNZtGNGB0GRBNu1xffQ0v20sJes6EjtvqEwZ
SaiCtV6hcEmSvL36RvNIWDt8kOf8OuH+tHgx+b30CQXOPWZzY52P1LnM41foP87G
E6zzyH2e7uvpxaaOWB2CR9aOTwEeqsuPu4UNzYZCzy+KQwEGr/5fPHcGEOvCFB48
/dxR4ljYUlikEEvTcLdneKpFc5PF3gwFc6afGNpNtGR3aTbokNIg6cmWc9PHLV4S
ODgU8YF2c9sNS1RrMK5d7NnO84oILwdmJeBZkzXn6p49GB25MkFAWscyjLVIlLZt
9R4pyGHyQX9aZ1dJ+ckIuzejTQrO1mwHrwnGNXZ4n92G1mFgDfEO09TEZP+wZxdy
lzjzJ6LMElCS7T4vanlzZ+XIvPSIm9WUrEpxW44KA6Dl2l4sYQIbg+db9adarQi4
AUncSWcNTQrSqY2hOKPy50sREwrQmgeMTwgxdeotYV0uoWXcrHhRmNVe8xh+JC+W
sSOFDxww6uGjF7ydTh2W0i4L439Cy2nbzdOoDcZNB4nKfDjp9wCKV6Vu+BkHnN94
AnzkwRztt3JEMmbBxiOhOJt1AxAGu/Ph/x4QIs+TIsnHMOXiWs4SwTZSMayzukPr
em2Fr/VGfgZ5YSb56+W28bhpuxssYaFphCKtAG/z6GMKQX0WQMwgpfFQN1pw9uAd
eSDxkgttEAxh/1zT5QHQtHJloi+tJP81dwmJ2OOYLJqZNcM+SJYAnhCq4v58Vjrg
MowJWYbKahfN6qdi3KYAXit0k3Ersv/7h7iA9H92ALnAyM5RyqcI2dM9BMmiWkDd
pDJdDA1xORMsdSrj7NU5oOZnTGJC/5K1b1KkTzoeeQ8fIzJNrqLU6ppJD69KqRCY
ZyJdXP+AqtQMou9CrKBKNGZCoWhkodlPSaTzON4zEet5RVQXTFwgPp6TZWecINyH
+2GkP1+3T5Ru2sBMHk3u/G2rYgB9vnMKBm7lZFTZTd6pdZPcRHyyvAD6qedzt6l7
E7avvEIJ2z924JmPVjIEcNjKO2SOyv9Ob9cH5HjXnK2DU6rKtH+31Pt3d7aeaDE7
QIBe2AbfBPoUZQMS5rzJU2M9hYRBonL9tMyl+eXhvwTIWd+W5msEPy6lozy3Oh25
WeCtPjM9ce+TxkFIJd9zHmJHUoHhJh+FM5zXOn7Tbl8+CCcfmZImaWwx6vboBGPk
+AFdWpANum7jJzI42h/gAjfKWrGpfrabp+9hW67Ydhzdg7S5PFqcDuvcPGQK6edb
NQM9IT+kQO15AySE8lrdGQwJwiBYCJ1nAycfEgG20te9oGmxcehkI5+MmjpxGPKF
f7ANOmj0+hxSr05XUr1Nqrc4DeJfemSDALO4YpiFwJ3BIFIF7aQobrwLBG6KlJ31
ACx3g/GzQwng7uOhaXrL0hjr9hRAkiXmYB2y6FCk0SEiI/ejpV9jKmRdaqoYK3zk
mmkuW0zSxFsOEzDYkTWuWUMOvOc+JkUT+SpXqHUiCPFY3UOQTkmC+CA2RDnA2pwX
8REN6Hjn9dNpTo+Lk4xgf64nGOg0y62rdbvUv9JF9E6LvHL0PMUt8Tog9fDjDbL4
PPV1Yd1Hoc20tl0uD6JqRdFRw3otXGXD6tyXLB9zqswuDuWW8BVVtqO9K56sCu6L
u3W64sYxtFXrwRNneIMpQ9ImXl1PxCZmqmohW++Vu4RGIGQ+KVOP32BZxJPENUA2
mKugPi/FgoNTo634nygT4eFKAeWyC4M1I4eOM8aX9wuVEKdirVFETivI4H0k2xJz
prNOG8+dODs19eL37VL67ODhZtFOhyYmKyXkCMSJfwxkHyqDmppB3kJNyew3HJLu
shuzsf2W1XTGnRgryvBzAHhAn0SfSNo7IWQdDYgNPkygYK3OtYgazwgpZDX0djTN
lMl1NUrmc7zpIbDzZ54e1pEmrCH0vylIBN+21zqmK8TcocDnDZqw6c/ucB7Mxy5h
VFtd5/bSBXAb/Mv+6e+R86vhm0tAHSaUPywgwhuOxDLewacwjwh39hcsippFcx+o
yRir3QdsjEmNDDxaheA8R1WekZkLFOxbemfy+2zk0ZSR2WgGaENsMd49Bq2U0OwQ
QOqDtY9hFgd59FxAdST4spIC3Kj+rr+cFbVZ2fDeyo4zVKqyZz6aoV/B6cyGGLNr
eVRTC2Jy2ZB2EOqcU+jPIwtUOt2PxkwSxpenbIHZyVZTdZJ3nhXmZN0i621gnbB6
kmrH2seV7FhNHkrw4F2yM17QOLkjsyJGpifLckxTD1bCGuB9Mcn1PwKs/5O8T4xQ
rzmI9SkfOTlX52ncw7dF7cG4MrfVx55snfdmLqnf2rzWWqMAxWgt8nM3UFr7Mzko
lgiGmHhLnZ0Oz1YKXy+Ig6ziMyXU6r+BwYxwrxZP5te8qIUxfZigk28Z/UdJFgz/
KvtcKYX5C0pt4h74m0Mz4FoUxNj4/GTl81ZAqj/ru/s3ymMZTx0Oo5BSZaTs7AuG
5AgZvf0IQldUHU8bUoXXrNzmBbyOeeDZRQd8e5l8XTAXF23pNicw/iBsLIEcCWrU
5J07u3jhfQshAlbf0ebbCwHIbSaFKfFQrY8tb/QKEt4SrihtwJFg0YrHsRIavwQj
M01KYqan9SeeScHvknAeZQVkbvlTwSNLSCRtOKnjSAQhME8q6fNZ/7VnREJnz5I3
UXTUOTpRai0Q9qLOm+9kl1Y8q8KLYl4gQaZXb/r+5lqTiR/MGqWwhdjYkUifcY0m
0qNahRkPEXqIKE4QKUZFH75T+ykQrNR3yrko48mADk0u+hlKtiJCVX6fW52sxvao
lKU0vgAbD9hJK3WexYauVvlsX3iKhRI5XNfm9HaNvvM6CBYxUmu7V/St1Z/bBUkx
GhFOKXP/eKgRHa0iG2SxLdhU2HSFkZlHE+j6+AwqKCYFgHHvuqKN5AEtIsZ3m4bs
CrjqmN7nz2bbLfdv46Ry86LCQEL5Vz1CD38pHnqKRT3ffp7OUHZGUrnngCidySH/
k6UTrV/YHtvfSVf0f2BFJPoov1T18csvhoi5rjxKCpJHw5kKcGUr0rnYjclJ0EF3
jWECVqVglAVAeo+5+muWNkcsw+DfjV/jWMGi//AN415iSWFXQD/iNHl2CFE0RGUm
6TEc6Qo9HyH20e1yaIiQJb0yd1JeNkxnvL3R9hKPRAeJY07fM6GjNX8bvm5onX+Z
NVWaQdToxlAq35wR6b84SusBxB37weVSsh3QmTFXpDv6lM7ybjas7KzufXU0uo77
HZ+jhg4TO3ynKRpzOVRN02272YjF3ah1v5KmgHiGSnGePOhl831is4rFoBSYyfkz
3WqjGwXb3ZpdTjF1CWwIiZ+JPVVGM68f1ZbWDxyNVruSa5ThFEClTY99CxxwDXGI
XV2qimzrRtH301Nqn1JSKYgYCwdoKOc4HaGAv6Woa4ModZwyA9KMcpSGtpYoYlND
PbtZ8uy6gGZ4qBOVMZeX0A==
`protect end_protected