`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Jm2uGAVYfY7w9Y5qKstopObZuZAEY3b/Io3MSEcWLhjjnKulVhCBBYAEQrAzzGsT
vMbffkdZgjdXQUg8jOLJXSHZ0Dgbnob2vlppjZs3bgyHCF7MoJ35E+LOsaLimUA7
hlqStcK49hR1hdeBPr/OwfT3UeVrRtQyq0eJXQ1UksinX1G9Pz3/CmcGfTZ/C72x
p9icpt0bkY4/1I4GBvNCsA6FFKH947JqH27OPACiQQRW/K7JToQn+1uhWr3LA1od
lbVrWu8PdZi7zW9gK3jiW5GaPjwbYQGqeGFs3bTKBILjb7sYHxfxw7eDLVMAIu5D
W+OTIN4JiHiE1gCnNEvkSQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="pm+c2fYA/4JT1uhlJGVUubML8hZi8lME4xPobg/m8uM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
nBaXksR//iZ9fraC7WMJWWSrjqRXHxmM1Y0+KKN3b10NElDzVNMlR76DLrcnamFd
2n7uzsxWqhhJR5LBl98SXO3Y90J6BMbw+OBG/MFM/zUulxh2Si5YK5G9GCrG9gvZ
5JomxuZFDu9CzlWGTuRUt6FsE4Lr6sOL1P+hraQDpMk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="M8TXDiNa0BVMX1P60yIvW2WA9jKGGy8GtbuPknDnC9I="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 34752 )
`protect data_block
/5TNZvs8Nu0G+mfp7M8H+iVAGG3Mh5DYZ0Gn3rRNhV8b5CcJKgjQajrRoGl/gSxp
rBAhtT8Vd5eelHgtvBjpvFBA/EBUrRH6CG6pqRt9r2qUDt4UernbZbxC3BC14KYF
+nUFsqc9K1YQwskh0vG3uzWBGmthq3DWlnC8DWuFLOe6wRzoge7t0gzcI2a58jPG
ypRWE/AOzQNjuMLiR/cgUlUjOTg6LS4fcH+91SNWWKrqMmaX8x/wrHHi1n/sne4h
G9NFQXGCnAG1+mlpfwMJesOlwGjIRcqn7fgZUnFg7+TPkILO+QzFCMjT3FOx8hTs
jsNJcyzqLyUQXk8jMJWnvJIG2LQGlSFHN2VBA/Dr6b1Q9QBxxY5tkvqORnBDjrrS
APNnMNyi0yZWfQSo4jtfjsggeT4ZA4Dpe/oRCgR12dpePn0dLzx7IdleNSaLcH0h
0fDY9OwW6K2N5g28g55QZIJtVkxBaRMmLnmIA60UCuNcm1mxFoUGhu0S5ETfvFRx
0df84Rlhn9CGyocB+BWJYeDiR0H1kSib0a+yn6cDTg2Z0xrr6G0GIEI8SYYFMFzr
909kRcRsQ/4tQN85Mmi3kzmwH865SUPEaWF8Zv0oyGyKL5n19T5LU+h0YsyxY5ju
cEMaq5PI4e6MIfFdK9va1LBHrc+3fPV7ezNRge2UwrqJlN67pXwBQZcRb5RHfcWJ
X8ngHhnRBUJddOqqsCv8QsO92E1cgQmLPIXbX69Q32kuNuf6L3VrcXqkKF+2qOIQ
p80hAk/70Q+JhhpG225drotUR/5sUMDFEYJR3tTGvs2Pp7j3dU5E2Gn7uepJvwek
vrVp2Zhn+blf6nH+tmayoqgxD5CjGgvqijquoJGkiddy6H7zjKaZF+ki+z8yK1MI
dG6gockMQe74SfcZiXCpE2wTymsSilptHsVxSMMdf1pfrCWTKpmlybQK5QSxBgiF
y5pmTwrUHrbyX/MEvQ0dWAflT7/u4rwVrf9Qzri4yb3HdTYsroOm3kWc/xyhqdTr
2qjolhFNDl7hFITmcrLUV7LHy4AZ38Q9Y9zV/qzCAB0jGfvufc05A8dNCHx/ZZFa
sOoS2g74SYxa3w/TqcNUV6EdUT+V/eCxYvByyZPiduQeHt+M47kInB7VWxQOK3rR
00CjtX20yJ10Ny9ILUa3b9wTZ7fE9VOhfelU/lxaDd1xXtofslManK3EFnnh5g7W
LnUn1sSmdwedaedjwDWDlzI7JJr+HkYQbHJBVFg9VqW/7ubHzqVG8/6Pv3HBbptv
2b4hy+1lwcgkqQM93GD61DhpvBZ2iNE0w6GVnWdSrrQvsmfJaBFQgKsov0gWCZNH
oipuyJOwIbJyhEuxLA1+ZK4i8lNcGYMzVtfK6jao8RvKwcpoW1pkKXS/6TEIR4xx
OcodrcM+AN/O2PTX3oIArk7evnAcgA2KU1gsFkqIGgOte2wPImKVM7lKrgLV+6DN
qN6Dhx2IOMyVHwbOretFigMiVNiLVIGXPURhYARtNmDkjP0XfsUDeiYHZCwb7fkm
ZC/JT/KwFd1W4lnKjKB4zfVZhNkKKZgI9VjN54OIEIre+W64Tw52MOIRRz+kH2rd
l0IYBYpR5SBuU9YQYkdwNizj6yzRmOWpQzi6fw42IA5qsT/HmhjkKRRuh8pI5dNj
JSdjOj8AA0ztwiyfXN/C5odiVSMlZv52dhMKSkptU6z3cyBEEjnHhVXi/C1f3M/d
75kn3Fg306P0FXoQCoEhp8xJiYXpEhBgBDD9ta8X0hSHOn04F0Oj55XdDp0rrldV
5QabA/5ZK+WA3MvCudiiphfAa+/WDYrzCkZKmCGf8qyhajAqhKI4OfrHqgoMmsEY
7mu6ZHIB+8gXKTBG6aNVJ4tSuuVW8INxb1W/lj2zuVeAJKWn/VCYRqT0+pxOgwT6
aZLlzHg58/UDbbaMfvpgvo9ncwklxK68jUq1DhHCMWJIlEofzYJYMM/IifniY+Ex
CArcQ0svLYJTmI4ecVmM6tb3NF5GiLCW8Q9i7iIfaeLUCe/Bvg9hLC4tJALabe5V
8LLSdEYFjyFZCDtf23IK2WTD5c6SvvmtAQP2G6NW0ue7W77xnU4vo4sA5jRSq93/
p7YGOWDVwxGINy8PsCwdNRrkuYvhtWcETwOeXX7LQEtP15C5D8Qd/NfMqmqmXn4t
Bj6UwHhVyuMypUjVFdWSH6s0nnIEudB6VbDxG7Wa/XkdPPyhB5V8A7FjkFcTcApz
94x5ohEgzD18XC5V+OTi7/4ZjKYEyD0yHIBufuAuQ+ABeo0qkiCpPOgn8ddmne+F
nISsiw5fsFEuLxQ3hRaztagel+U4J/tjtiifksBdpsl77AEYUccXGydeHjd4HFhz
Hg+lmYVrNINEBd9OlZi+XddxzsjvN6pisrrKpxPyYxq9RtJnUHzzhHByZF0PQfJU
NRrShRuJFbdiuhbzxbGwukJTJzSE18Z9BxOIqZiopxxf5SS1NzZwX3kQYS0sMMmf
yZ9NksPg8s/cmB02uNrRH4C7eo5EEjNPWycAGfGh72D01OiO/826ZmVpQOcw0oD4
nae/Hiu9o6ebqO9NnzJgP2VTPzJcDC1PdJT5uTV14XuO65fMZVNWU7po7JlrcQd4
UwjKLJZ8X6OHAbTVJT/HRmLL4l8iAGbboHFSgX8LlAQQBxHcv0DxM6Kcq+vEtPu7
iJtMvHemGKO46o5GsUjv5Wq5s5+dkV4lUNqInFV2lNRNbWppT0wQMDQJxABz4Q3F
nPWiMhTl7HEKnyHClUUv9TbEatkvoihRWUlcSyFSfWtAy5Hb6UjulJO318kc7i/w
hm86n6jvypja+vVpHJXp8voSYFqmmgIj1JxT6+tR2eZ7Qt+tAPML5drar6dXMUqh
EqvfsiPwLwQP9CeyaMxBYbjsyzci0LALPvyt/KFhNauImWKGR7fq4eQf5m0NGenY
fApW6QUdJ9tImFx6HfZVl8wWxOVMFtDinso4hsCcmMJyVtZk3VfKwoz7QY0hkJLb
BC9+7rnU6RHxdSio9ztQtzFf7tWifxYUqIGIZNdxcp35DGsbtDd5L5c8ek09s0/T
WF7j8nlLmxWutXrScJZ+7vQFygJtu8TPDdWZwRMuOJhrj7x6i5O22fCDlqEe1hDT
fS2/BLEWS/ozgEDdwQKXpVbSjCdWBz8/lSeyKFWxciZmf8zHvQ0YC4X9YdQ/RBKm
snHjEnh+Ht2VwPghXVZe1V1tYmQxn/sJ6KfK1E+9s8TjqHddl0iIXAzoU23/wFN5
Z0fH5odMeX7w6vNWSh61jZTdzU+3XI10wru8/xLweUMvA2Sn/27VZWnpM4/poe7n
JfC8jtGIi7mlh6N+4znP5nkFexCVycslD33nHPMa3ZjtYOI7nfpLcEigm7WCPefj
MJS0Bwt9BSopLwURaRjrBBnEZ52NvbSwUth5UF/Xc6/UXglQhvP92nCRSjvMsGur
xk3WwsnC76QvnpGYPsq+yUKX206rttQJjkNbTYh/DeThUyV0/ByLX6dh5TGcLaJF
IzYIRaGm1oFiEk+VwHSC1MixruiZNcDUHuwkP3utk2qO8MYWar20PdYt5LZMSEof
XJvNf6Y3WA+msjQoDxw2zluhEYaxhU+hqJwdc0ZNHl/ULSysAmbLvLe1gbGte1NX
4rSlp5oPfQWR78B6KeEz8ni1QLDOIDepIF8vbvf6JfubALM3aolRms7B2refaMTE
533iJfnQzXwlbiSPXJD84oggr8GxZYquHBkmBbWG9yKWruSra8g4DObxIfOP68o+
uRXmm/GF8GJPpvah7Sbchipeu3mLHKFLXb8Qr5O+/qnlfhtYCd/TMVyRtWW2jlkl
NuJQmGMHr1rWAUCIp1kVsyP8+ntvszh0nOWDPDlKiFmSIzfJ3EK7H5xMKYso+QL1
2EvZ7IfqDxstZvPRaXUIlYQOUpJldJoZz9w7DTRJDy0XDUD3zZz2wgFh5/gbc1Tf
bp3zg+nCKV4S4i9WDAZEmOGIfj4w+OBn/VM9wQX3ddCMXa4a6rju4yla8AXsHzYS
ckO1WxUXNFiH4Tups+vYoMqLM+xWJlHNfvLYQMzerL198lC7SPKBdmWoI6zd7Kvz
/7NY6xeeHsTtuI8oO9DWhUh6gyq4xKByPJCznxtIX/rCD4BWEw6vWOKYrLDuZ1NC
I/vW7rWjDPCv0OuAteAJt79oOmWeyYB1//C0OG7sYF+Ax0sk+j3pp5bl4PyoiryU
jHMi8FI1vdXeR6dLjMHDiGdXUSXCP1f2FRrjwMBaP6Ivxof5ff2w5MuxCKo60tR7
PYw/BDcEhhUWKwqZo9PI+/u5+GCAveNKXmMskQOU2E0HO6JWcDNjPAbFMIAi002P
oY14IDqIdPvOkylIXD/2LuN1NpHlgk7pRzOJlaIONpidxJU50A1j611peScozUYH
iYJyjD5ziuIJKLSWz9UkAwXH63Fs4pbSna8vJXWDUgmn70N9j0C1TxdwYueyDEJJ
TiGRnqz6MGQXiYzl4rQFxRrgwh5E/Qe9oKWYrYybS+r7mJvONr7XCY6uHyy0T998
+j1mHlFL5eaIoyMRgQ73eeUB1Vx4KhtIQxfPohaQ6WFqxiE/WNQU7PQhu3Am8MpY
UkXdJbE9NYwo3vAEyjmxz+FEp8PyEAc4twWOe+2mciBIFDGJeiENxELhLsHn3vNS
SyDrMfi88WR3vIiexrrdM/WTfU2LcgM5B1fvs6Ms6TajsHO/q6q9CjPezOUQcYAI
h1Z7sfEFxLT6bOIYLJHrqF7RMYr8KMsoH2IrVOKEqoO+XnzLMOHQocNlqmy82mlh
0fKhwweNbD04O06y/rlgeZgWWa6Zsq8VDKSp42Az/GzGbAsw9AFs5iZmGG6W6BnW
ah7J/mkCI6hcxgnxu9WHUMTqhLHOSIWV/3LZgjs6f4m0gjjfyap64xXLwwi0TqF1
cvQ6l/VtmngXLXPmlYvpwU6LADhfvg/q39hMnBF/2GHzrV0TZjXUOBReXsZDaHfH
AUizIoRR5DPdFDcjYdSDDgzcuS2z1f77EYJZiVhimlM9M1FyhsPKLPj7sxQHR/DW
i0NX6eRmH589tbO4PO6IPyDFFICG/EZMoqjoEpU8wF/+/OfosFW5NEAcsYWlf19e
YA0RfUnQlW6WvsMWNOVskq61NIuOTWH3tHrWJQBMDGy+/IepJ667RgvICf20ipmp
GCvVqgQnDrYzc5PL/dCS5hh8HbJg7u5b1um4pG/GbkSwXmY75kswwCmI/RF3YhPb
jARO0HNzYgSnkcqTinj4ymrwcXBxYhOz/hrBMLBzeaQLzFq0Q90W7BZamqZWwBcZ
DGSLbCAH10t5YlnfDO+x27R/EzVZsx7gykSCWJCGBTfSS02YoCBW0UPipP7yKE/u
UELbcri4ChMM3FqeZleqPLhxavYZSLFTJsc+nEdnbrnfppMVKBPvhO0oa99zLwtC
HR7Cd9Ymfz6lisA0bu/+6GDtGybIHfYFsK1CeAgcdTvjlh2iaglLWpoZ6tvnoT3V
tKABLf06nZ+B+EumeVuCr47GfluRQvOUQqBQdheYQIt70zxXJRFM8/Te1inCt/i7
QJPub3dy4sEg/j2oNrM8m1jA9ug6b1U6D7oaqrep7R9ls/7uHTTzZh8p2uUNNga8
1xT24jFcRfh6JwkyFSxbcXeDQEJTDNPET1u7jD1HYCqJSZwYZfbL0HQfgcNos8VL
9Uo+dnc7qBj7knEkDg3Sqxbi3bgij3F36NmcwNch1/mPbZtGtx13Mv2C0iH0TIfb
6w/hYnuQSZ3BHdPrJo5kKMlZgpv5Y57T2134wHEtUeRjATISVKaCkjvaCsl3zauU
SRv9JLRr0cEFWuGXa0kdQzwsFokuZA9Kvr3bza8qRcSmcrd3ALwBBAG7qk5tj7yf
U6/u96/d8dP394PQpEsTQQGf5rup/v3EQ/pmhWm/0aPnsXDvX05YCyFAFV3rNaRK
V15cMeWHBf1ckHm2BILRkV7JjldDLtwso9pp9XixuSKnSPReWD9emAw7VdcrjUZk
CCKikhbZk2MMSKC4w6JzsJxoQefj6T8+5A+7zrbXQEZLg90b9fMvb/du7pP/7Qtg
BZNi+zoDvKaKrQninRhqTVjpdIvimf106sTMpD3CxF+3S/LUdBOMlUPDowhcE8ak
33bWd2sRq/fOxW8uEFkUjxMTdhPCQd4fG0KPXVvVbkDY+nHCTFDMm7/3fMAIDNDO
NV01kaij8le5lflAFFubOmqj+VN3ito47FrZg9M93fJhY9tLgW0AIRkiZgQoBnhy
9+4QncGrZXjKDZV924wH9eFdW3cbBQU3QnaSkuw47rvLQ+8Y5W0IJTMBlafgECce
mAO71iaCBVNBaUBA3CfA954mgOo4XoYGLozgHssTsBE1Lr/eLfadD/AjDEgOo6th
y95YM8TLH5GGvsHslDypTzezMiUY03DBTknPLhpG1ORJkrgSN8f/K/mgH6qvoJtC
7WTNmU/ZoApaWe73KRunPkvy9IpfbQZp0lMGqc7FYHFgSJDUbeURdvOUhV0ur1p7
QCE2aIde90sFHeTi41HjEp6c8v1X2jMIP/vA+Wd3gLyQ7fuLumWwnQ7z3a7Jrsle
IWxZrp/TR+sW6SbxE4TG6bwegkCNb1ig0VlstAMb9EgKl0cZGXsOBcbZ0gUgKAXS
x28orxX4RKnV0UFZtPZgIto00iTk4+27n5HpeikduvRvAD0RKBx81YEmdpm6UURq
4/B1G3eUm/ORbp5SIhItzXWvnM4b+9wQGSUZiAi1fDb/uFvQAaIyqnSJ0WssZzOb
nFph9jndp7/2CuTR42kCDJ/+z7Vyl6XTQZUA/s1HSopwvzUEBAFHcswPfxeCJdI9
Z8PsgTOtfsLSJSARR6JMnKUWSYK95mNiua5yKAymQ3OrfcNEFouk52Q73430yWtE
e8VKo7EJMito02BiP1qoEKlPnm8Y1S3QxxXsKC6BvTJ/C6DUshFS5yp0cZCzhWEt
J1BZ1Wm/7uLr7QjyV83Agz2OGw9SeuJ1hk3CbtrFehyupVwE7BT919Y9jkNE/O9A
5zdhprnbWqQEMMxDSpq5UqjbUqzLYzK5wIsE3l1cKIMg/ar6E9n8He0lWxMuGZw6
p/POX8/Y8seZ8sujFKwYcXJCed3/KMCnqJYWYOeQ+g5VVvHkM2W7Eay65ACbOntD
vhma0FR0DD3DDECI8CmIiGYIlfKT0etoLhmzlRIvWT2s/Nef5YHZ8cbLINHm51eZ
YSh+Gh60nu1hP8jlNPhKmV8OWAghGciyOJ+j5hL7lTtFyuCBSsEKcGh7pl7JJj9p
YAnWq40O8ahywlrZM+KHin4KF3mcHjFBSjlZWQ45NRsGOLX3FFuCgXozO9zRKp4C
q8jUZ5vi+DNdcFEY1VtW2pc8PCx1jeRxLtvrDUpOQIHMcoGbG7HsO6eh6A0Ki+jw
aVPqRp98tPVzkhrWjref551SwsdakW19SVaOapm2wUaeGgoGQvO/ENdLQtFpuIUS
jHLw7RsHyLY7cA7fLQJi02r/BiSVswrCDegTnHy2XreI0FaHXCPtriH+maN5Q6fb
ppDM3zuGQY+jSjiSKPa7L/t0RVSgEYL4hjvntRfaguSUAh6j9V4ZW7nM30YcwPIx
BXMMNZMteLzHXba7bIq6BZwnvYR7GIc/VZ6qKZIrzIvZREJsGgadR8uAp3wdCvHc
Bia12JAl8GJpelIwy1knADa7RlVLs4jioNK5Pu6bFF0tYwAwMUl/Uabcjc7ptRBL
Tr1OQY4IQ/SD0moYt7MzTc71MjNMUSsoJ0GrduWdc6e70a6ytv2NJM1zxk/ohaDP
Fc1bkRzIB+s3BvK0mkL/+pwMUDVHerc57+tx59uqUO+Bo7Y20rnLG29GgvKTuAxx
XyKg4b22xX1ZmRhU+XH4JQFRBPJRDUF292NwXCs+WNNo2pb5s5Q4QDwpwxc9h8Mi
JMI+sFKb+ERl/Gbp/a+TmPtfHhD70rISkIXN7Jr2RttSgbBgPBqdVFrx3QR3obqm
zdkl0OBsno7/6waAmuJIPPcSsQA7WQylq4p2ltRPbVzfUODK885Fm/ncP3m/VD0b
3+e5dGAQcYmbOnaCCKMq0fFh8PqzfcRN9ASF0pD+aV55dMRsQb9cV7JQPFKP+2Ur
XgY24oyA+boXY7qpbQzlbbNf3Q8ghY04SVzaOuN+5vyfa56CIWUDk4o6iCplQZde
m0kid8gWw+9q3yh8kvS6ScpNFN9y2CUb6KJX6J5OQi7grL9ik3RoZ13znyzEOP5Y
pYNfugCGH/f0VAN3tEZtOMzpnCWSFnIhW+1OKOcZgEJ7b/6qMTLLDH/3s3Dv4OGp
aLfguSjdevTi5Kc/lVIBvsaVx+AyHD3w8VR8HrCsig0YhVert5ebRX3flK8xdegV
fj+kmbqrlfwfj4scFDqAejzOpNmgFlBAujf7s2EShbkfBQO0h2xWS15vFg5Ea4P1
KmnWKwxEoTTwqlayIpl4778kx1CXbue/TNG5I2xPaRPxtNewiNY+RhyIpB0Ly8U9
W0UmwDM6HSv+n0vpba1ZZcbD+PtQ3bmLgyITL+Ev+/xfHavf/hjuKdRMuveTdvkL
GZFKUgYPlJJImsiYi2WCH8UdMlDxcAVe4pU7rfW0+FVuZRvFg8r31OBkljE4sedb
/WX1FcqZluMhH+fPWUSRh1rijF1uVnSIyjIF17A3S9+5Z5hwJ7baxY0zLMijnmfW
na69PcePP1cf8UNvGydlDXlJNnM8ZgWBjutjmMNG+hHZGxmyb3coVPz3HQsjoRfF
rqriWCdL8tJyOo7fc+e+vuacwlbHaRsfIS7S33rNtG63VxmxPdnDCNBHpdr2B4cY
U7bdIWX1c+PjkgKo7gZfyeoQwK/Pvu2ctgBPh50ncOFcZ3U9Ad9asHL5Z7S+z65W
i72jFQwYM+Ue15iTOPdGLWFZJS6dnl9aqLV0Q9eJ6lwjI5vDoqws/GJkbbVx5qqa
Xk1vtwNnq256bn4b4YrwHJr7hen0FRR3JacOF3pVXWtK6oUxW/meQi8RpbgzxngZ
f4FBZkm98dgcYUugvURBkX9lXdfZxudGrnirB91CGdA62O99DB3ZpBjKXK322CtR
XiVtAf+s3/wo3bbZbC4cgcLqvBjywAaY5ly8jCodTOppehljqKxfI8BXoCI53BK/
ix3lXzWM6dDOE93dEZFKr6YlbT7Doce9mb4QbTnIcuMbfLD/j1CQK54c5GjZ+nxN
6AmHG/aZ3rC4/5Vt1d5vQ9erN1NGPdsof9TT6Y/iwgei2t7WmBLGR3eM9lMg2ep4
AkJYWHtAcAhQvuwzozhoMf9A+oRjx8ggTl0Sw6ChUU9B5xQb/bngb/oh3NQWNZxp
olzz7rq+6CZ4a3n5y3eT4hIK1iIqBkgnHpeVOvzAu6s3XnYYDLlazPXztVeIuqh0
5/uTrjS9/LooZmBfxfnKkkPFmxwdnWtmtYy+/jBIKzb8Xihnw3aQvPczkOm5toOY
cr98oFtBc2pFrRNZ6ZXO+sWOnyBGiViaLQ4ulLbwlWOcOkuL4NTqMkdm7hTyjeRf
WEeX5xX480tTatCFKZFFL5YZoLkBUhxi6pdomLAAQKtb/wBVBPLoKZZejTOY6F1u
3CBDLQLkh27PWhBfObkYQ5mhjlbStsZNU1qmX9J7B2HS+GkUxbhYP8RiKLS7hZ/l
jwcjlbvqa6oFUmxR4AnSQoB7dh6l2ajGAKdaDNj9Q26ppf4d2uze7jaZYZHDH30t
fqA61xUFnwI0xPZLWiDRwn/X+pZFH9ugZbLc70fb4PO2c0EVBYSenxSRQJjnX53F
P8T4i52lgqf1w0ke+2iGTqZbzpUlOxufo/wqSsD6g1W8m9/3U8+pe7qpo/qF+E5a
WHGnHftgdMdY7VvRKSrlByfEVlplJZpXJ34c/Yi5KIrNH2ZePZGbH/s1ovgwz7w6
5JoiBm609RdF08fxmyBs7pAKqVknr+d+dghFqz3I+DhyKaH45i6LJyB2+seE/cwu
QjIKsMnzstkG4VCe9A8ZdAlRIiP6pI4Jd0C3jx+JGSrhz0LNDqv1o0l9VyRNc/QU
vzZuyZbHJ+xLFQXfR8d6qbEeNQJnWVw2wNlyf1D8WAsa6V711cunMIA3Rv/go/RZ
1IXmn92IXFgEKVcw2s9TXR9XD41v3zYTxsAPJQQCeqCblFZV8VlYYOb5h7FOPZIV
crv9nzVvKpyLKcBcbJAmU+dY3F9YPCDiDyGRiSqokcrxHJgaHp+DW2FsyGTJDDqZ
aAcZ8yPnHMDgvGdEL3c639p5kW2GnEEFAQR6tOuK05lviNb+lplvGEO00S1VThEo
QnCkFWDh4D2rk6oafCbPqBXESDybVxATY4kwAiSoNug8rBKHVNj4ZWYVFRqBF/h8
B0zhjWGhuMN4aPUtBL8d3mcc5jZQe46cjdbc1K8gsS9h8pSn/UX4C4ar7mkRRJye
ynqAL+DVjXUvObxM1yy0GnPss+awyt00W+x+gbAQfCf7Ai1SeGPAePuMwlsg3v8L
4LlhGsIImH45fh8Zn077yjI42bijlX80LPCW4FkZjCxUknZDNDFmYQ/YeLxTE7S7
uGRsNDzgQgidbMN4fPaf+vvrY4K+1qLFZHNzguWjULg2+6JBHFjjSPnWa18dP0nq
NjCdoiabNPvTfjS+YPlEdVeKS0Anl2iCFJMk5shrtC1E04Y87u1FsH2nTGUiZDUf
exW+zlg7JvsRiz6TKn27hP3a8D5p76WXA2d7CEfm4CXu7z3RpaubjvGyBNPnmF9k
Zzp80giM1xX6tr0ZzPq2NzTeHD8FGm68zBJcFyF/q+dueN8QqKEYfzQQcp/c31PS
+amPIW+iaGpxRMfsrncM44GqFbbDDH1btCENv1SCpAHdV/88y6OdXidsGeEJJSED
RjHAvkpqMcbcrh18kudchNEzwgXk4TkIDiSU0i5mZ4ngeR9dZMnliUBBqMP7hwZn
GekpL0kaZTb0RsKUiRT8EJYQTTpq3xDmSPLNeioop/WLyTn7NC4jxcmk5pExIZe4
sOuhDKlaydO3bSPHhRr6Q6BH9H9xYh59MkSQFw6GcXTn7Uk6uAlQnsjhgQBJDS3u
TlXrcdiuHfr5DLcPdplpArPnfiN9UC7uE8ArxFvwFrsRc84E2HMWXkmXBAQ4qc8J
g2ux9VnkbQF/GbNqtV/JDTWEznoylJaRw3v8gSWCabqlo501td8rwtE2Jl2dO25I
+c0PkoNDexNOtceiq29DLnCYzTHw1nMzO70JnuslNlC249kBeDJhGIJ2oKLNRQZW
93YKJAglJ7x5Jd1Wc5IlmXFavkC4M+JbGE4InV1AAJnICozdldFrfcAgY2HK9YlZ
Pxl5xVgNTyH11Ew+MVd4vNdeoFrzUWh79WqWuvz+cNuV9PKM3ppLKVYTd7ayYeTA
AwpDHPq/Eywmg4hwsrreMF2pr7ijQAxMvUKFOT02joualXX7yf5YrTEBY+MueHCz
KBi3m2AU3e9rk+ljVthW/MuyJc5p+7k0YaLANxkTo+Ko4zBT0j2ZiHSgpMiAkkeD
o3wv7aadkVqd1y6naBVngY8Y9FBCz2KOn6ivxpqdDQh2XEiiC3OXS9PtssF+rhhx
vpBuOSnbkgFjwA86QZewd8VmKbXKAEBhKtBJ4Pd+3BNe1+jmmJST4awviGErf9uo
PQeVu/rsf+NwCKtOoVpsi20SnhbAQ1aAX1diS58xdTIsBIlSyzlEExy7bBPqTZfO
SpBCJ0B3dVKN2IsM3Am7IRGf9c5Jn+1jfZvwKnj6LjGLIjPFNIdPmpe4dqKc8JR2
mOO7/K6s3IJWmS8Lk1Vr3xyZR+R0Y2VE3GYB4tbaOexXuS6nsxh7mdWk4BtKpBpo
xLKwBAm/XqwUXyYn6ibejWLy5N0G2gm53sGI2Dn8YbHeFCi7y0fqVKNpHaxZSzuC
GfKq6YHM4hAMlHaor+XHaiMoprRbEIOsl2PVR0Y9HygLCQ7YpG2ykQ9WYj5XDa9T
Gd3a380UaXUtZAycx9meDvii6a4h6/YTZvH2jHm91HCd6asNbMZk/RMx1lPUWAEb
AWu0tmuo0WUaJcBiakfPAQYE2C3j4a3WH5OjwmlnYhDGcfgZcwe2hjk4DwPzP3Pk
muwTBDijQKJcoggvKUKRiQwuf425HgUyggda9PgKdGQw5epVRsYDmoC1Q5VyGPhP
JzxZkk8Vzv81PYL4jHE6+WjsIUOr98SgoydwXNkYEJl1Gfa2XbIuGQ60RMa84PQw
/NQRBUdkiQcOM3KcQGMUPAq01taPv9hPw24DUzV+8wWPSsT1uLMgO8tzVwXEhvKk
hqq6zYU3MwdnWWoiRS8MFR1rvWINzAYB0VTWehhpuXuLnlhMfUm3hB/szlFB8lUw
kEObLJgvSdDfTsNu5Jr0H9+RFuxXo6rpCa8FmMUJr88wincvooA+zuO14lhfmZRi
ynkNraRTSrZkiQINVjbjVXokQzq1OQz6n6p9LedL7JjzKOi2E+Mzzd6qgdkAQZBn
ileZkY+Or4l9Pqg80S7ZEKXu3Ezy2rUMdNobIJy8Bc307yxT5IXHUuq/jrRZ4rM8
SXSura2wr4m5HUHNeCxi5NgL9gAYCEc2f8boeXXyzO4GVujPz6o4Zt5kxFVOlPua
7cyoI1z4fRBcCrx2pSUCUDJqHqZndxKs74VEkvy1ptiCiobfxZy39na+wZBiks87
WsrvkTxUD7mcBEtcsS9rIGOl3xVwqgnD2R1/Z1TWb/Qqg0LGB2NZVynBR6dL72j1
M+ILTUg3FyLhWHlWJQONpwkSvKPGQ09IL0pkpNXeDhFI9BCLFk7vi++lKq0cnMg5
etyk02DDp3cPTirZ7DNcKeDjXW2TsUFc7+zaPQ0QOR7uJCILF9Z4zow2bmqIxGSA
HiMKsWu2DF8koykfBcfHT9w79rIkYd/Mz0MRyH/aemvcVWKMH3JEaUW+hSkaNG/A
vytMY1YzBw+VSeJymLOHklhF0Z0dceXKhUTX+3BozMy9F04VJIDG0rrYQyVZTs8e
m2rSamEVlfsefAhKqAOHziqiR/FZOh7DMxJU6spo5cYk+ZIY+gcoOzCd+ULmItne
W+SoyK1VW6slzvBN2aex1fZUZxuwE8kPupMgJ+Wk3JSTgO/ztwU1TSYcAyG+kmWq
+eJtApmGtAZGPYdzCy+AmNH5FbfBygyhOB3/7/e5DrgsYhfjgwJXgZpa3MKK57sy
0DsWnN1KAW3YrNcEG8xx3xUgsWMAekYQrGBHpgV5W9DXshpPvQAvpKPnvzKltMih
xAtHOBDN/K7dt7ZKB4QaRCH1052DISFW/wVvpjMspBUhcVJC6+sHMcsNr11yi9uu
DLk0c+UDh3dorz1ITkwNBOHZS7n+2vw/v+n4c0aZZQfyAka3dpAHRsIkM0sWHspe
0ZenrL4W3jslkFZfhCLGsm6cjtaG/RjyfpAfd9alNz8Yjid5/XQnmgCVzEV1FVda
8w+zeGwCDKlrpqn0l8HrSdmiDyIK8DyXNQHOOGaDDZ6Q5zDcIi4A3z3w799YrjDL
l9UqdD2Sx9NSQgSJ6YTWgnUIJAOVfOxsaCQtnltsHRbIPVUuyv8whi4N9rMSSdNw
RzhO0sH/QS6Bcwc6/CmGegwC2mZJMh27jkX+2Xe9AdVITPYfG8K8q/XzfGuSlcJA
/mF+KHfH9lOTrl9NxmUxtUg2ZxxjGqLN22QbK/30gcbOq/JkDBVcb6iEtSCgssCD
l7dRmyLHmk7oaoS4hEfFCOfeQqJ/jUivBvDn62h9ArpDHJqmjnD2duwwK5u9W98m
CqsbegPgE5cadtv8e3vRvx6dyS5DxF+lPH6dFKjtE25GJytWQTBpU2lXxc8HWhbR
wLo8x5q+z9RvRz5oYTHWbmepifOHpjSIvwzbQKLO8xPAVHsCYoJEM25OMG24u1GP
i9rJREVsBwFk5vT0BTHagWGeCoW1jGk8rU12qVHmXjKbsBEjSi3ZtawHuPrWTQ2L
Ak6/9THWzNisaoSE4bwkDM4UF63Y3Sr9eQhWPZpZIJRQFJAwJZlMiTMbqAM6nMdS
K/84z2wiNW9vpGl0kaKV9EMzS0mDFIP966LBYzjsHH7TeX/Z2ZmrvdhGulz365YC
xaIx6BnUEer5A6cYCzCXZevifxavcuPVjL4MwLVMXR/ePVNFoJNVUCzJUdk/5/zd
TDLayyhuUs1yYkQpi7YVO3J5vsl3QZgyYE9QR99eSfFeANye+CWhS/T0Z8gUXuPm
5hA88EMrVelhTwLhH6ybvwcZoFUmx+fPEwx/fGtsZ2rcoAne+mi6jNmed55wt6ek
Td4noEzukE994B0vZTw8hrD+Uujg2ncO+bS15xMdavk949UL3bhB69rHLkq4bLga
TZ5SetFldVe2Fnxs7P9LT4lywH7b+ORi/pgC1yZ8lIiVsAcQoY/Ohmsi5GGIhvO6
WC7KxyMzzdVU6lgGtocoRtDfRtSht5kCs34ms61qgvP0G9hTSEpfEihdOSizVdGg
iXUqPTAvGH2BSiAwCZnCYlcYPwso21b+5hBKEW76emsHjWXwQ7Pxgk1NVrb/Cm77
rSC1qT6Pcpmewf4Qx2BbFLyskcmJQc6L7iF1smxJGkYfHU7dnDUEZxtckx2G29CK
pP6IJ/sce0vgeBZ1x63fn3TRhJfbgXjJ+IROU+CN7/2pROd+HyDiJrVXc4eaq+Mw
20FA37nXBLlhVGvyYYXK6zbkPX6J586DaPQWuM8ZxdyHB5clCzaUm9S7evmpN6gI
cpePuJDLVrLgi3SDHauY6u6YnhXqOo61DYRFp+UxsXX0+e15YmmlF6m8jcT3Gdvd
N4hhu5bmJr+dOPZ/SbPlRd0N7aVQEyBBCtAJcFmEdDAJUH9q1Pb+BfNNkeYfoeXr
x9akJGFdWe/vcefzlaEnnW7UHdVQQciq+5lW6/rrGCtb14Xc0fmt8pRtdO78jbcc
cp+cJNh443dFGDBl6e0A2kgiAIhCv/Zf78t/InIr1x9IFSKx6Rhw7eiv3v/mDIsT
484tswQNAixvJmvj0xbEqPlJLzCDKBr7DsfkwlVofdyju4HIDOCtJcVM9SOfxhbn
ZH06pKrWF/UG23ZgSjoEoCevwTxTKSxMXETZJQYtpGzfbXFrw5ZJnVY2016mstrN
0jzx1QoZsgr5lH9CWpI6WqUgHLsnQQs6MKGtuP9H6bwKuuHcTcla0i9NteT5Ckst
Zx12AEnhDstfOAnXTEcyLhIKh4hJnaLJN8Tp4ZhCJpFbgZSWyltHQNpJx0AoDFEa
B/Xn3Rhmgy78kWztlmHr01BueBQZn8xETL7zyuzHITJM8Irgj4/+O32BtEmtz327
dlTPKXrwAzHMF01oeRLRvXN8g94PFuJ2cZdMKs/twmWJJ0uCqLGxGonbaY0HyDps
UgWNcutgdNDaMupyjW6WJezCC8A9qAi+P8DwZfAI9G82+AAgWC26KUVgw7/sfMTV
6hEStWvPRXR3oEEnmkunXv4rHKMrCPVU36+ysG55atS/FW14Hj9uztXzhNSlbbcV
TQMGWjytJ3REjz56iPrk7OF5zduKfQAV+5afCSnh/w2Zs1yOvcIIEvibc2YkiTXC
9aE4HpAAvND7hOyrc8vYzE1nSX5u6I1KUZra4D175c+XVewIUOZVCtKkeYtEhkh9
0sxDdwWXImKuuxUz4mj3dL5T2UR7G4P7rNGAtDESmnq0b02VXZVlmSwYQBmLXdtD
lGI8vpzCpgeNerjzO5LdGFFOkx9xWIHvdQp1uOx6EjCcq0C0leb5FnhRPtpdf95x
vlF6z5bpOdPJLKqVCmMtJ102q/Nou/RmKov7xUb3Mus+xYo5UlU0bKPZSltcgefj
7P+SrS4Eq8wro0zRsifo08QL/fPHKkMm++t5fRiFk0Ncwp62H3Jt3UR+UgGaPe8g
J9RIHkD6iHvtS9OFgLiYZfEqI8T4GweEMpQ5+jasWhBLBTSW84xDTowLE1YHzrGG
BTxzMToHn28De7/qpj4bjCb/B0+6v3z58IfFPMO3RWNnl5SSS69nnimrVMHmEuzR
UHikpMP8WqP/0djz4/Dd5hjYOtmqxsOBqHV60GBAJRqd5jSr89yyzXTwfaMd+nfw
o5ixSMZmOlASAq3+i0WwJfvG0pnyTo68n1s8XzkB5+RMVJaUsJ7QQlqQ1MNJeMBY
2ghRtK4MALZHKe0hunKpD7W0B7pTxgf0mcQYzTSRg4Cjhcr15GGvzzUZlfRBnNOS
EAtOiUdcL8SmIw6fGTgOtxU+LkRBm9c+ssEnndScZUwl/JoC2jtLc8p1aG3sPm2e
dyegYtLF78m0/eEKWHnAI0wMxoB3kOgirTmem27dnnQY0AKbuuomFTQy3dOXqjib
dF7KQ/M+hJW7lNLlm0LNcwCpJqC9AdOer3OGbLMKM5LxkSTHNIS1c6Tzha0wUr6Q
+XuCS6cCw78U476lTUdoCzOCIuMX5A3tbSsCTF17PI5/fmN+dNExdiKHY4fSqcLD
ZAYARwSPrVtbHAl5jTt9am7Ey4qtlp5w8eQ0WFmAfqPM1+oARhWgeYZBfFOuWL/N
TkZlJPr4xBvbyuEaZPMwRYWZGhKi/31uZvWRQvCEu07gtyB6foqedhF4Q14C4VdI
4Idov3MSI1DsjPNf23/CWcaPmnPUNoSZ9lqCO9bi6TER8lpXg/YyKgL9BRSnqXp3
4/BgPDgpG7Eub8sTR3Yp4K1QByDtjA26pp8YtH4E3/yoLm2UMmtVXn2uGTQNGUI3
5P3vo7xQjBMM6oq4D4ZUtn8DjLcJjFovPViCROTdQOHWHI1CfA0W7b0RfRmQPLRT
NyCvQH8F8s59+2yYapIZefuScVaVwWC+HL1VMgh1wYq7seXKqq7cJSUFk/NG0K7P
gBVkwkkhU+PsNyfiF73c/DnSfjz2iCaXgzFVAiHBCc5LDEC1GCPx+gzDlGkTyYy3
CWfqhtRqMdfx9BKGWBKUJwJ813DEd75ytFMpm2yZWKTXEEPtc23LQqu1qkX1txiE
UK1AiBrKug6szL2IBph9DF/qqfatzJ7vFMOVI8a7txNyhQuYz0AH+1YBioLtUnRe
CiR5QMuA78RzuZusYoU4f9AXssZdDqVuggcr0ZEQNPJwlVlHOGgLN6baLbhJq114
QyQCu0VsupYl7pbC98WlbTsdj3a+uFffo4UgAwMdLaqG5drn8Wq7d7g2Sq9R4a3W
w6qYje1F3D2RTyiEDsWSKlLi5BmWmKPbwcqXn4CqRJ/cWuHS1XE2MQ7Fi4jwoLqU
RnCmf8vvfHowBnBl714a81cjquRX1pEvNtrmbZpkKUYaLEWxkm5rl8D5jR7XL8Cx
6J+fM+PgiwN1ZfMHejNzybtczxVOd5F3q6iYSWBVkk40qHfbEbJumBklERI/yaVb
fJw9Rja3S8VqgcW4V7IyLPiuXKfVFw+IGqENmIwe4QZt/h/UrFCj6zVB2grtWZtN
+OUKBB5MHDHVGuiIWgPXz8kB3SYd9vZ3PU2owdIGOVQq7gR+vmED7dUiUvsCPu3T
gWsaLr4HEjCbii2B+AHBssX5tEccobOXYFZDVS3M0SRtzsMt2ERAAg98qE6UCMh6
7+GyhyQ61M5EVz9mXPDNXQdKoV1M3xM+HgQYJSvVVbkuT0xQVj1OYdNeAs0OEhQA
aYrnGPtFRQB+lJzm4Doawz2/B17gzgyeHrVKj6x85hF1+guuhOrYQvOFO402oi0A
9DVjRris0wsCGcOA5wX+Uo7ckzjmh3ilvnE40hK5GNKU3NDRvbqfRXS9H7GifTes
72KWN4CyWOLYtTOm2Y0WaZbTSznOlAAHwlKqtJnQ6riWXp2x87z3Ng05iJv7FowZ
FdQemQ5f5HHHHjnKeeTcWBXCIuDTSbbCgghA1BPe76m9uk1ycB3anuCZk5Mle3x7
m2tNMYC12JNr3/eG7H6PjBJpiDyzeGnR1Xgcu3SwHQNoKGdWVp811hNBbnCSgFO+
B2rtLw+T5iJGLUvLKnJ2h/fxHlUyakpHkkH1Z/c1J0Z4SYTiwh42RqFB/Lg2paRw
36PDhI7+IX1dTjbhILl25cAEFCdChrLFVZwgq+lJd39Em3W0CWC11ZIt9A0cGTDj
oSh09vRWaobrSsSx2K3LBX08e810hnJpFWYVHY/Py7Pa4YFSoWQo1KcvdEYj1358
xmGtwcTcV+Q1tV+vPqDj6v02W5Km+Ehe8tevxz4XZml+EgSZCB1M0dZxkAogDS69
xNfyPGIb7gn9X7MdxRJsoP6kqKVElEKQN7cm4TGGbirLp0SSD3FoS0UEdJkkkndd
LR+VgQTp0UFasgzhvGATl/jJ5g7fDJnJnzZQgnFPfIkaVpDP6T04VSusWVj1tUO+
z+sIOp4DBTdrzMdQYfriOsXoWZ+vXzjSTx/G8I0idkK6hzoG22uJ/NeD4evj28oS
jxEVeGlECEkRWhbxIHQaXLNCcANkCBadQ+Eyqh+X8rpEUVtoX4A2j5cBm86TvWCt
Sc6p3SCV6RUG4afKX9GiqghgDDxjn//1WPwZY90e8MrnQ4jcF4yo8oC3tCbmR9Ez
CblWMeIF3nowiQowjzhIeZdroeyg+VrDtQ9CzIYsvOPyQ6gWmo1WLTuz3OKVmFYX
N9LhSVpyd0/JH4z/z2OVgzo0pBLPPJWcv16bBHfMKdcsRWdJel4CwzwyyVTyVqUI
D1DwYw/fvYD1Nn4lbj2G9KKbItHUbwmm3Ua5mrd1EtkM0GMK3WFhbX1mOFevVc3f
6XHVzyUh0vYp4c49qcZ85L7FJkqoT73wNz0N50CSK5VRIIaVSXsKrq2g0KrF/+z8
C21w8r1ObVD4Xhr/IQLd7Uc1+5s5RHrnjc3PiqCf4ZG03vVp6bCDrEhtj5dpUpI9
vgVocU6S58Q6lXW0AtBgtpM0xbcnfkfmMwWv9m8rpND7R9UIhU67EaXEilDSnHjb
itRMVhV+ZyGiTRvIb7WogDvZpP36vmEV1ojC/FWkz1m3pHOo4TLr+Opwi77x2OQI
w5uFFk+tHX3BXlmcV42HZKZWnb0Am+AQ5hg4LPpyj8mNzLTziYai58LNobvHlhkB
OWX3N2HsfPWWm/a9137qJPTZ00ap1f/Nv3mtV5oJ+dAHPVfjq0nzjHoQJ7i0yrkX
JVzDq5xUhbaujYyUokwH5dM5vk1F3X/s0oZ+SCWbdmFFWO/pEctSNzsg3mGr4xG0
8LklWvtJMtPxvHldft5jrSVqVIS/4h3rzHlZCe+W8jKqzPf+hhhgPFKVjA094BhN
WZpUNoELzBM8WMrFA+OYZpH4pPBDBCIAk9GfKivUb6SCg03M1Dq4zywnqU2uugca
SjwdbFOtcSv8cDICgAiae9Bir+n29CYbqXQlqj29NuTud2I6KEQc9kHpN/+ttoJx
NCVxEeM9237dEbs0n0Hk8rYnquFkMuo1voH4BFumDUcz0vw7MwnCs7mG1sdVqbjs
u3cZIWOGlgNkoDMulzWwEOWs0ORJndwRCkxoGwjvpsuCmSP9DLnuprR6jHlTRWBq
ZfSsTyfAjG2ch5lF5ghh3P15XbaNaK3GYG/GCq+rqbueZBExarJdptDgY2mbRh5M
KGA8mAzsim30hV4M8lBNL1eF9lLA6tF0hOBdJiOciBiKAAFEJPtRfIjM+J02ELFh
xtNfGR/uB3Bl4mvpREoQWbt7fYEANtaTKxDWDqVF1AZJy8XIBQ3p9HSKxjmHJscr
41a8yutaX9PJeYuWKpXE9ZRpHpJIMgHFfGmbdcbZmFqVANsMOnIZfNQYPvaWIjXq
eoNmdU0qFO6HR2DZYBM7aKG5UGNHNNnHmxII401tztHPIRI0BqS934WgLNdpV1e3
6LfqbbHkNaUMzUxibyq50QWFFBCgvXgJSHq72nRhOxFpjvIRPGOEScjQDvDZ2IM+
7GXBfkcjFwlxuLQHh+ThVjEBKV9DP2R8oiG7hGOvEpIq2Iixbvc6PQrP6AeNW0S7
JAdst5Fuq0ugS5Vs7TbhWsqUVpHOVV6o4iSReSVCsQuTZ65cePYrNm0AYIT67e9K
XLt7YbqPQKaQFv2PcBrfvF4Sfu0l+Lc1Us2yaG2qLGYFFUelz98cu6aN3Y7njnaX
eULXxKFvfOD1tv7IN5f02cVcV3cZ2qPC7Ynd/D4KjWTfYFkKcpRvauRwmHRNkqZk
lb/wT+ib5kND7LozP63ADbGJ3LZEbhsLNtZJx9LQtNIfw2rj4gzMhY7Vv5epHCjO
e4e0KAqzfXHsXYWj7DKDBct8H3zMYM0sdPW8S1Q8/2yqgv3roXHigKQ/0YFUMgMu
aFuCMSMZ8dpWreEzfRg0a1OEBQwJ4uaSiCLf6MuN4dSvpgAYVcnlI0kR0LIVQTwN
E/YMX1V7ZN+c2kpxdZKuDEdjKd5BbMoZMXSm15TA08QpYLLLGtzQNkzQnulc1P5S
WFkSITgPknZG34TnYRM+P9Q9wDjeS+b3IDgmdTTir/fIUocGWiv0vJjJX8VQbmBq
OkZpiCzfciomsyIyCsOgbfDQwlnkjNHXJhG+CHnCw2534yVVvnY6YOTc5OVm3pmA
urDSW4PhlC3Fj4kalp1eBUrqcniqXtOrpm5zeWQZ9u+vJYV29YUTrO0iLL0vsiLV
cfk2dlhYPO54TA7p/6yznnj/DREPdcmU8685r6WPPLAruJ9/vRN4mP6KpAIyrwmn
CM4qvzdb+AmmNM1kJXEqbu3sYgq/5FpE7GD5LJZTPhQw1cL1Kda/mm2MsfXPkE21
3Wt9xQxUTn0XIWYzAiSMfOaL5Ci6/iLlvhQEfRculGuRk200OVFC/5ECX+asHuFL
ISVdNi0fWwvJgbjYoyS+eE4jxtUXWc93isnv1fyQDDe2ttdSOnE2NuQAGqcHqMhy
dnQzrCC/EN50FgmeafT7a+gjcZLH0ANRY3plnJO3GhhQcmWZtuvLRwtQx3j2UA+S
6VMbcjOurBuNOZcViaUC5c8Hoipw/YCiLsletuJ5uFGBl9zKGxsrTp99rA8rGzBt
4CwTQnHZSNoJgj1G7p2jL1RWwYev4Oj40MoI6Lpik0bNw2duqTR+V1jbfrvXEsf3
0aBc+ZB+d6yAs0ehK43UDxtPsvIueWX6YZvODmwJjDItnwQrteRFe+2r3MhT2j/1
/AMAuBFifUNF98rCpszzdZr32hZSzb/32bydiBsN3uCmso3079tYJrM/sw/o7lfD
RAPFMq4AaLt6ikCYtF5in0x21U72PiMh4w1XfrNWai1deYtbf3ao2SWrylk6/6Ey
OwL9sQK5dA8FM/PJDaJqMp13CPoMgwMRM1DxSg3plWEE/QRcZwTojt16wHiA0J6K
anfpi4VNYpbvrWKZGb89D3oqyo5+XYkDXNasiQkjsifzngbdaPhJjb9CDoSrbU6m
EgtWYd60go7jpi2GTvgXVPg417YYZG0dvZl2N6zpZuCWKYJ6Iyf2qqHzvNzsW8HU
2lchfU2ZHOeAE7RFd+vTu7Ezk52uf69l1OF27ZTayaTwLizjl9tHrXdu0lJDAali
CiZ8AzY5qXLK7PiVEaAA6RzZVAM8kxN+wkoC+657pvwIx0tsCO5Np9/Ji7vld4NO
hy0MjxOgxreQ0xlOOymT1gMZF6551VbDtXfP1I8ybftL1q64FPpFyE1n/VxoF3ul
LN+TG7fv926TWrSYKeyTVHlE0FuO6NSHQQ+Q3mSSnig+AuG4aEkfYtm6J1WdF7Tn
wF27U5t4NlZ0sEJREYmqijQN1kvlMparhHrwHqbWIVb2M1FydgWhg0VUiBI8XuJa
JJns88JZuNgVhZxYYM4sR4o3ymyOSTbKom3EsfbkHPucqGjt9EfsxZIyA21CdqrF
QUDolcD02MyY0KrgUlnLuO6NHen8BdlIIczOnc6NrOYXwaS3qszDaTbYAxWiuOaG
E2bMGRoHX0rO6qex9YHyRZRXB2uO5RmvJqKLUku5KySqs3dXUkpmHa8aVT4QD4Tc
manp6d+OmXTevemfYPLCEAEnX/iq8XmR/f3H1VPZrrjZZ9/HqU8Yehx8HdjcjDqj
7OH36+vx6zEn+VgOmB4WFvkzEJQaNFneWUp3CGTcHFn+ztuCTxCZ65OEeEXRgc3V
gTWp6OLc0vBjchBemvdH7wU6AjBMZgFjoEeSiW/B68eneC9kdfnQ3+GDZ1mXtGZk
En/9i5svmAm1EojT6w4cwC6cvU73knMK5XpWINXkaLmddvGJNKpUh1/gVAlnD8PR
MdYhCvY/jXmczXfoA50y7Ug+0bkBTXP0PyiBePf8j4wxtbBtVYYg+kYnfqvUHwW8
UxQR0VW7iJXG/53yoX6CBwOs9eOxJyOeTKJnwhwbTLH7hxOALl5JU6OXs9HIw8FR
p5c2IsGNLXXqanYRIQ/fYn5k7qisgF2SESujavRAkPk4KrMQ2n1tcSbjkdb2fjLt
zfTIXvfUvJmjyKsWsAz+lOZY6DC2NTQgBsz7liyrnsSus4p1p/EEML855Nkan3VK
Ir87HNIIMUrSaeKQasopLH4WUE8/ie0Pg02b02hVYKfneaIIJbpL2fR/pzjsr6Ca
oWRedhFvjfkmDCqooypEcjkWx2RTNA9+GWQgxHD398CajGDi91J2on/dZCaQAAR0
Llps0l5rL/8F3cTilIWiEdfItUbfVoN+nQi95vcciIkcq/rn1wwmkxzgbGSRfDTS
Y+4FUQ9/Iz2BKyQ8N8NAgPDOs1N0cDSVdq8rMBO7oqII0QJCnBleVTttMFHC/JXe
eQqFiG5EkLSTw1rd5BEJwTZAtGvLyHdW5mW2pSNMptBxgltiACZEOEFRt9VzZLye
wqrYES1m56CfHoKUUdoFiIlFArehmNudd3j9p1B0HsEyIfxXib4vSjFb0Oha9sE1
3AKLUcT2Al2NwoKDznMSFQp8DzoIHtyyIKE2eW5JkZL5ohMI3u9mOL46c4PQ6axP
JYjbOlXZm1icOcK9AZgiYWSnfxg2Jd8rV60LeQ2V7PBe9P1b+6ay99p8kXzvH4gS
Q4YftgFj99SaRL4wUr0Qb5jtxocUeGTOxURe9pEYWk774bt5OxupY/J7qggEYzCL
PdeNw8Ov7Zoq12oxgQt84slOks+vr+15yGsKY3BvelFc8m3G4gJY+ovlVQy6v4Cz
pG7JVOqhPFMdaRGYjXTLuvIS0sUhyrN8G7gITrE5/2q43mAKX/K7t98SFHo2us+L
CB5swJwVcbjqa+AF45njnccH2hFPvrlksDOVUUKkJimCioLUZ/Ricoym1XRdfg3r
qgZzA1nBKPDL3BmLdVGOryFarFkmLypMmZU9+FqaNI7jUklrGebaA8aadd6UHWOS
Y2efhRuLb8lcwzXweQW2zAYd3pBV5n8/Ryg5H29CD7xuvJK9q931KLy4uTQlkHrm
SpbxUzxD+k3XrLdtKhToxWIuh64t2K+ZghX6qLwaTUwE+yxvKDYUB7szLP9IqXU/
tCSXjydCBV1M3XWUJrGGaGBub5EX8Ho51674ntj40roedyY44u9UY5Wg/1+ZcYPG
MybTeVorMhiWPNUYTxDbCuDQqFMkC56qsTS77t0DwTljwcdJqt+0Cv/7kuz4eDpn
dvso5EZZTFsXlEt+9Q5WtPBcbeycbBrpBs/OCkVV4KAp6H2rJiG3TQg1UjW1t8MU
RMVLPywxSQiE9NEtoGkSfSOebkqzthyBm2ck4o4McQQW1Va8U6KCdv4VYUwdXD9a
+S/kHlKdUEhsTcV2bxCELmM3tKMhNsfMB/cg5WuB/MMQCa7rSJBNcElwAE+cU9oG
nC893ENqyVoYB5eHPSZpE6SEX/eA5mJS08tJv8JSVq+rGNsnxtY8Cm6nA8SJhGxW
GXP4gRiNKZL7z6gNJAs0PY0axLlqV6iBv7T+CnmJiSp9XoBsSSq7qmePwp2RDwns
cHLTmloYhxsZgWIKUS88vcmKV8lusG5TtFJjkPG7zIbEwQLcmSeqjlhNvgGNtpvN
nZvst3tuDHhHz3ozj+CyCnqyLmw7cBHJ9nS5wEZkU1kDS+LaJ8W/ejhXUt/rcYmo
pzvlmeguNmB47vKRCP4yhlX3tTrcLa7huG3C6D+t3Ie1us3sZwEuIPK2bafUpDt0
eVo1+3Ti10jgtrWwUqWpHmSv9N//jgR4jxqvWymOMlAKotAlLdTMhLhAwfSaohau
CMXez7e3Qu5LEIgmfN9QiU2LoUh6NVqIJyJ/sjht1wNaU0SYZ1WMZxdOqs5IyjVp
b5RHyWiuqNLe2/CvoR+Na+y0JCMb0GoqT1Y/C43sYZ6SD3C2CF2lUdnc4IRvQG04
Si2gI+aKGdFp/8mPJxmopg6Q4z/07ejQTH/NAW++Ae6VWD1X7prDCsnIxJ3b3SQb
+4OAkLn5eOwx9m5D48QjOaz52xXJO0QCsQiyh+7sCluFEiELLA8TEV0f1OJs5bIm
rDsHeR4pbX/c0zK9rvEgN1gUz3gN108EzLcslSfwqQJL7DE/qyOvGEBJ+rVD/zmM
NlwRjECvd59ZAYXdbsbBHQJQwi1kLehO4/ztFwvP6dCn2twHXlfYRBWOoCnJ1rkG
vmruZPxPWM3P12o3P949bpec8pB5nQU8aIF7pYMKLFjUkBnCwvO7gmh7tj56S4Ug
wEXtJLLs/Op+e7JqUZ2K38abK2+Fw2s/Ol20OsTuByqQPnOoCP7NgirjvYiMWZeg
TfjYQK1QZXwGl4eTttlVXwMDVBAhmbM2PWM3TpFnmrlDgzPVYE/he11LRE06gapl
3+NF7srd5ZZuOpHQM3UWHt/ZVn8qn8RSiNWXyXATLZVXOoRpNFHEnCSsTtwD+W8p
PDA6MsiN+C6u9eqOk6QDT+/67rSyW3L+lQMx7ie5b30kGpe0lQ4hmncYR9XVA9xd
k2o5dSeY/TaNjZs6hp4OeSie0N0TyAv/NkjKxkU31aoI5pcfqRdhkD7nsVFxjCJ1
AHeEdbDm8MSbHYGjpxoJnnG/kIzoSk1ekObgUISY7Q+Vbjy00/DWz7ofSu8YYwzZ
ysgm5d6MmiyvlUiiMgj0U/V/oJ+rwEFLjCT168KyHUdOQfuMTl+BUJIPmcV5DCia
pJyzpPDsJD6gEvv4lZnlK+nXK0ds3EKRr+4Xxqe9fR//rHSxKpYSB3F/D0TDNCDt
NbkzuvP5kJ5mrLWRvjt01ppGu07SAmZ+YJDIFRzqWY+mndtbkeqpuEBDkt0xu7xz
/2cJPNudGBbHINVt8BtbXRKHcxjjYwMuplecZ/0G+JEyyJ4pBK3V5StTidsfFn3h
IYq5lxC1pA5EomFWHwDUSmlzQEYseByQ0Q6fydDGXGpZsbP2gl7uEfKZW5hk8wck
yVNlI2hvxTAOQGXPIwob+DDaLjDo8GoZ0w82E/1Ml/+rreu9bkg8OWM0rWEESii+
DSEwqMNOVExKWP6Nynlkm9/DNCSe8IDadi+Pe2MxcIoWL0PLK41blAYeRETrlSCa
Z9Rsg3MTXE4cKLbfVWJ1qVjNj9yyA0rxE/7WfXU9vK8P04z1fN3N93j+SXtJgD5H
/Vq0f94bhYzZiR6hyvERwST2fNxnqVIKVEFAPdITCy5FaUqJ2cnKu41g0GwGXF5R
6+xN4Uz2csZoMCzwissiZGmXSgG2sqUkam492BBQVB1Fuu+dvXyToNpmsBqy5bQP
chrTO6KvHQp5b2S16wDFKU2n2tBwofo6wdd0pZ1eMgrPoj9FxKwx9XxJfq4y8bBg
TpQX6RS4cecbQuNSxLaS7NshpWWRtPBkTx5P4P+1xeIYQurDkCOHun/WuUKkCSZD
On6AKUe0ARQauSII9nz0Tu9kj7LbfdPmBjoaSqmPSCYgUu/5rwvL0+zhQlBc3pCE
By4rTQi0Vz6KB1Dv8FdDljcMW9iURUdRQAJOzZ0ATaMBrV1OjYkwoUcwZHof6DxQ
pbAFyCffHg+ImcGRuAB+Lnlsyoce2RSKjhqgdpOSFxE+SYvJp6j9KJSftD4mRAiz
kQUK5Q473crCfp8UNg/9QTqlqp8aGtXcn+TE4PcO5WqNpAmsxpoFRTAM7q0Sc7UY
71K1yIDRLA0XhtJc3wQCr8hrGiuR8BPBNrHLMlaJL6/sJbXEe2wQAg5Srvwya+ow
xwaX0paohYSrGJFHVV8dmoeDFkLtG0+cZA3SGJtHxhvHCX/uRS0RL/EHNkW4YtM/
cqW/R1505KZ3+2sch50qb1/roq/tq741SCCnts02gLzEx6BUnTybf8MhnDhZx1vr
vuxXyLQIHGxBmn8IcCjxCPwtYgoPPTE3TfKeBfVHiOvVBZiducPv8SvbTm85ggAo
7wvsMaM9dYweHUL+FXap38+wynp0F/Aoa3u9VkvS5VHDG+tTwfdCh2JW6NC3JwdX
Uyo4mnM4DF6YhGu6FN6v2YrQRbXsgqbnhX9lUr0TuG5hQhN4rM7LyghGcGXI07Ym
dGnNVsBJtmDUAqvjiRdmZ2esCCh7U7x5o38Mx7q1ELNlAyaVmDDi5gloosNRx9AM
/Ng4dmfgXiTMOjQvfs8/8zpmbDF138Ib601kQ/J2TeLM7L+QdmR55hRqhUyeKGa5
E4kxoyDSI6bQtEl9hsjQRx4+s4PCrGtX6Zl9EN10tjhHHAkz9R/kw3Ho5/WUBZQ+
5YxEVJad1BPS6FOyYPoWLFvdj/NQ+qqgjqfjCs35KcED5a3+mZ43rdmRdIu2VyDk
PFWdFk84dIXOb2BiBmQakKTsdU8/JppqdmM/84FX0CkJXWTRyW3LFKSIrTkeLmCn
t1XQwF9Sz52y61VYPsW+BWBHxOMmtDDGrwvA3iSDIHZCg1/ccGJVGEJPyDFGouQ8
pXJgMm6eAazVWhCZjgP218MyN2QiYEgY8hGBjqxFTtySFnSsjSCveFXsFI09VnIw
LxXirAzLHkK0B039HvJx+lplTz737MyqKU9xDBbyFiJKk928G/mLf3iplnr38jJ0
xVYLYy7WzVVDZrT1FDKyter9ff/8XxPm0zAKS6zJQvAhl2nk365xzLOVaNafpgIg
Y44U3GFgenFfkVMrj9p9dR/OWhEEtyToKAV64RaGdWE7/oIfBQ2xK2FrM5irPYEK
O7MJFGnhrsdfxfLcJe3jZEa7hqWXNvsmwAKnC5zvPFcyrzYfKNa3W5GpS6jwQa53
jDdsrjiHg32gvktyty8A7PjA5xCO6ebsSzy9FH1a0oc1GztzbdFp89hCuH0Ozcz9
D7759ghZ1yXkzPDzDBsPVYnKHMFRML6RIkcgENl7dpEWg9c+68Jo0GcUPkHB1QsU
PxBGR+BOS15DckjaLXJqUCzodytn3gLN4Q+YUzHpsCfCX7sQidVkEZs/9528495r
x2S/Q1TZD5CF1RYhb/03nrksp4cFMJEB5fqnzfTBe6qg8hgqx6/oL4KPVjReAiyW
IYqoRp5wMi6c3SsFlf2QIusLMRJnwxCF+DRJIM9qt/3+uHD3oBm/U+ekx+zN0ohu
EQxmBgxwly2y4196GzKpYPJD6boFLrKZJ9q2CQ2hg6w3E3eyl86gLVmVHOUy6PZ5
BHGfbXP+L8gge/vJggSU88tGfNTUmjRhZLf1ifmK05VZVAM1Hxeqw2ji/1qtcWrD
KXu3oJABp8csjL6zHzpZ10APPxUku4HEXebbGhH4fZunFcvgXLHMvXv2KEcxWOtm
92B8awB/YhZ2VJjtSjxo7CJjmPd1VbyS8Rzt3fcMVug/k17TMXzm00XZF6I+3kbk
E44JxlZ1kR0+tm90iqOO0h6QOxsZgBNHdIZ6Dd5rQRij3+XCmtzWVJqS4M44Hd1k
pKqGED1qTnCMh56kVylGCWKldv7rTo4Q0JxM8VEIrp9how/IYFDThCnxnizi4/z0
fS/Wjck63sqQCVHojoAOgu5QO5VIrpFZmZBK4nvQeb7C5+aXrYdTTT1paI7MgJC4
2VIBaegYFz3/8m08SRRr5M//DrwAnxUaIv17KtKcId0E0zFTRTQuIpnwYPIULIfG
baK7kWdYLhJTHsxAuN7+/2n8EvzxGWX7xM/sVwa9JhOHNrqgIBsY/+/y82eplMho
bp+iOi059wSmpZmr4u+myNkzK+3a1y7O50ulo9gSSPgCDwaRRun3S0zz1787nMld
EfmtdkudQ6+0d7LxpXelLjHZ8ZQRIKKpAwREDSr4ejGAzWmXYvnQq9s+MWuW87kE
r/l7y3aTA9PjQLAdzxfDs9qGWwZsNAyc/cthky69biVWg+UMDAEFahyRe3Ub0pzC
yYcdTmagetjXa4C1rQaUjZlzgPnO6yBDk2SDO55fKALUr5n/P7UnHZEduA1Wfcmi
NHabSI+AL5rohZwmbcHY4NAlPlcnEm8y3QaOH799wsC7hn1mTuyNZbzaNjwBA0q1
eFVzY9U8pGy1cPfghEpLiZ/06efRG85WOMUj+L3agU8dqib3L8bNUyWHOD99YUmw
1BlSsEWYm28XKgA2udkp4RI2iC1aGuIF/wgQp5QmnN5un6xhAx2eV/vFirZt3PAz
NKKn0UsMezQ5Oy9XqC7hLXjR5p28Sr82p+Iynz520ohMb8ajvOMZM0r9QGFY+r0H
gIRwxFjWEjRcnG7EYfX95UTFitswFf5UFKk2cgTbk88eGbAEbT/+HjfrGWNvQNZg
QpYJ5mCgf8vjEwdQWvH/dZCYSmd6m/HSY6lZx+67MlkauN36+ZTN2rEs8rI24N2t
OOLcUVXvoae4q2+jj6VyX+prqcBGQNnHXU0gsOFXB4mBhlSjoWn5vOb6epE8ufDn
SPiopNztyxr2kQni2omtsfJgK4PWl8fEOAY3YQy0rV2OxuuySxAoRDEA6uSY8gzE
ymvNSAWBXbUcBuPhUAaXtE7swf71RtlIjguMnCOO/0F7jUQJc8ikbcVRXA02ckx6
DTzg1Zuk3RJpIlMk7359G0VB/9VJfhLCU9MaqrBDvWwbTvwIlNuecZm93+IwGfQ3
+AEN3LxI+GdFMn/1XGZFbn4Z6XXKykFSX0Fg8p9lABd1vpAda/LbPcifGg69pZGN
b2LF7rcrVC0vpdOMXpTmYsaFomvcwGaEyMGNC4CB9wRKK7ZmjQxzh1gHkhVTWtFf
D1YQLObrSuGK4r0OR3ANPBx6OqjjaJwBPdvntEClFRg3zoNy9ioUykxvgTgW0MB1
e1Vp+9gDjErmGVgJxkT+azoGizbqfg0qe7RdPdXfD7RlriYRPgkksheo3oc73iWW
hzv42so2sLB+NvSFA2sv51djX75yc6e6xjULUK22ye3Djl2fvW3s/njuFBRYhFm9
8FmOg87KlN+tY/xDpm9EWsEdyf2TRcQ5lK+CGidTG4guOZcKHsBE63F5xbg8X/+b
W0Omu3uezjwIBhrC+d2gOYeqXifUojr27pJ8WBZWbCCykS/49SbSkWr1oesKyczo
hdr/msPBJkTYCUJgZuULQs2LvK0CSR33lqYrQtpbeJfr8bwZu21iet4yNEw8Vgvy
ifPIMQriq+ASjM05f+BNqSFsmlkof0xO6bTGCdAcubyb0oCbUHh0S2xDSHdYJbch
R3RUI/4aJ1scX+qqKNBqj2kEGe0BX76sNDikHZWoOajXgaSWjRoml8x8KWeGrlvL
XQRshYlgimz6CyUOUuKDIWG3CTnR0kSgH/YVxxI4OpZGNk/xSTI8OmsSjcFhHvgm
OqpXOaJqJSCBqeUYXw3wiwz6uLOnU+6xvq/jkhkjgP87vnpO6sw2NGDqJ2y0rkbH
Y++3QnLpgdJCIrd4iPz9q2VkzIx/jzRiZp6eUcqF9Cy16B76ARe5AXDm+eMHqmZ4
M+J1LNik9E5Ol6RIv5npZTbYnCDq9np63Jo1XRVrZ9WVoe/u5XYcmosOKkf5p4Z6
6MlcCjECo5MNvrcdcGturQg5V0M555q0asPalv9Y7hi0rE9plgfSEbmzaV3Qwa/h
EN/6VqqkyZGzbjpoIBoaDtf2lONZvgGGpHbd/pyKY6nwZbDLlG0r/iNvAfACQGlt
5KqRfXJwWo8cf127SfHcBPozLGezKWFNQFg+581zGcqOig7obqsGvFkR+1s3VtZU
L9OESdaXmbLgVhwKrCUKtOg0GCBYuExE+nq2HqVlrlCW2FNjkFZFlAHBtqU5RoTM
j2DyHIRHMarmhpKPsAaXSorNTuNNadOpVB5R8fkDm2hGUDNRiddoJpE4ASY86syL
4rJG7TLUYPNrFdkIeXS1et1BR3MHYBfQxlCTqHawieQ6M4WqY7lPZ5gy0QdutPYt
eQlojVKHG+EPbR39RXibkYZStfJWSXkeglmdFpDu/QuLYJSxV5edB5kLPbBzgC/f
P0Q9Z5ZSqz7urJoJKm0YSxKf3GAoX2F2BHK+kMsBkgGkeNnu1zxdt/9rucR1Q0zR
DFnAK/ewkeLIr5NFVlqkojdzo5Iscw90VhKjW9bVtAfVP/uDLq6qikbrhkoOrpu9
2IXC56OFauTyKAz8p+bAZxpKia45ohb5tNc4Xof4mUgBV8HjNYYugGBxAmhJe7Rv
peH4Jn5QZ+Iua7uvc9zvO/chv8yKcXDs8QMt172f0ft43c8NXvSaWN+pLM6XGOzJ
za9Qj4M9Iu7N0v1RpHtzVQU1plbmZ/o5yXcMLdGE8opWU3BYt21ggtJNrhVwXe5b
q/HnS0H1SRB1x9/99IED4AECMA9eqH6yNyjZXyy37OrRZeKtMKKHV0ixwLdwUGRD
34EgfPLfALpnyWr1AnvkjSmaIDfa/KFSFRnwksf4japQNvmC32mIg0uPvK2QloHk
//bb3ugGsaHTh3igHW+0dGyOSeQxjtXiDvCX6UwqI2Q+ZmUgT/7RIutiGFmpWvKT
e3EwWi13aBKsf2+puEzd9QSYgGIHqESsZGgYA3TXwZkUmo1qVFNdFdtVTLhcHqUi
VEy7ezmTe0QLba8E3Fh/45UrExJi2C3pOJLZEjib7VHYitLlNNsLJizjQiHpUGDe
DiL0XYr2ccFYIey5RFWXcRgzHuvSUCLJOnrQ0UEiO6B+Vev+uAFtjRn4ib/EB4hE
DL3Yi0sC8tkDCeA3F4DM+KjZpOXwqjphDQM59PycgAkN4q32j3kT5r9Lf40LyXU0
70h0A1yEvcW0cr7xatspfGrARHK0TEZW/6/DOFOBSbn7agInvx0kHvFKkUDxTDpR
/8MYn0Cgf2wOmlz3rKT0H3ewfeSdfpQSGpdn0hmRpGrPouowCTrqgYVe55aK64d6
ZIkGlI2ubdL0plvVyGAIV6Iic58rbaqg/YI5ISLE/V88AV9KbnGgg8akisGFy6fj
HP7NPTmItF2JUHL+bXCwBcoPDesUXuiRU3HdZ/9ZYy+ZOEOQ4w2XWl6RMfZgQGuj
tCGT0rwNdawjjbNLne1F2gjJwDhylS60gK8dcMqNLAesFGRIzClIE6oYQg14ExCn
oLdqmphJANyaFTCUYvxQCtyiA4qFLfoWkZeMg4Y0VtfG4hnTtdAfQ2yRza/T/fH2
ZaYBQTFgDlDA/X/M8+LBlw/qXq6O5/Tt9+ju9rgjgh1NiFGH8nzUthE//vAN13zW
972JawqJZDvv2nmVDQLQjsDAJMcbykdiYCwo9kWLoFdWJoGRQwE+I5YBhROqhPWP
N8gCGOIEVss8wsejb2cpGb1nKAful5SmkTLG90PHW2uuGfwNd7ejGeq96U0av5v6
FXdQiZdUAYUq3RFV8snYyjPuPMhWtK4cXtZYw0ADqk50iYgVzJmqpZKOYR/OJ7fQ
FZhiGCriMGpkKnKmZm7QzSO/38TRlMhA2CfiLr6lgq6BoIMWDyyS1HwRFKjVbPq2
F1Lau2r4q4cZBFvLfQNnM6xIJscbtWz1DvudnIHnbDy69zt+MvQuTme1GHkq/D7S
kDDZ3/3ZydV3PUPgrRMhnhY9KgvulNFs1zjI+cJDIBpu8Vi1fxReslXSlT+weNpw
g4NSLc8OdN/2RuRVOO5hOR9MIhnwSpvP/Tf4TtCIfBL4LkWVWGjFmHl/wZneGYFz
jPUByjyTSkgKLOMtjiTxFXCytdiEtr7GXGw025OGjU8B3APoWxCl0VxolIkzKtNE
Wj14vRTQEvAm0jCuN9+AENHWraEka+rQG9isYXtz8BTbgWMBWhjj5EslfBbkSY+v
D4SzDZ3scxS1VWDaSfu75IglbXM0J9WFCBeUMVE9YtoHoQWSp33ofhm/cFg6QCp9
ekk0xL80sjTR2SJb/+FF7TREjq3Mp9LiWvhfURt0mIjd0Kng8ddSl89MNCwgiTFD
/FAABy4hA8q+hq06vshZdoFih3ZILs10vis7l2Gf3W3WAHa1BhvofNTGQvU0q+mI
j4ttIoEaaRjCZD8A9zfC1saAMK5EkFCKiYHGMeRA0FUlAOu3CSfdN7OxVLVilHUu
pr1kO4mrxat3nC5xhi+KhPCtzGfqSQi16ljvoDjNk3JVep3HmI/RYylLuO3kRV77
VdteXuXR1c7nE66sdCOIkyOllpv74UAlxt8WDces+4BDSQnZz/Z4/YUYboC6tXIa
y8PPeNHzC36Bc9u/RhJUImiC4XtnUaHtm0bgBq5IrApEA+27JNdzYlK6ODrtKfgi
sXu8FZmBT+HY6pMDyJTNTwHC77DQ98NyJvbuiAIdG5NU6KH5WN4bUCyruJg/wlp7
1unaeS7dXmxGsAzDdikX3ezcc195nlUCqAoPwUzL+ObUU+rPDat4iiuueLHywhgb
4lEFvR1Z4XNwHiLlCYeoJ2FKYVU8qioxXjC+U0w7/FCwHWzwJnRh/j5mlU5mqx7y
BsgnLUJD/k8nb9R+1hTPkEkQ+0mLODQnEAvW1sZ+lgJLWsUhpbXKeUHtv+cl2eXk
GOw1Z1JQ+2Y0ggX6Gp1hv+sRT0TwI8a/rIndZJn8u908RqoavctX8ZN2rYZUvS+x
bH4DfPrvds3Fmgegecrcjx5K15xyPXecjLhlQAm0SLarTUoTm441SiTrHLJ0fGSh
goFcuOG9Kr2KxaVoZ/6tjeCltp9+Qcude78fU83/GdFbF0WU2dtcQkL1Xf4e/HLs
bend2ce+pfgVEbVT+mCGjvZKx2Atzs0QDl7DWkrRuVFzWFuABoP9hCXZ21TTV0ru
C1s5SSjS7sCpxfh/3dNuRFRzTTIlle6F13JRM+AZ8I8cFn4tvke6fXZxFtw4M9Y5
775auHUBwytrJI2+v2No8GKF0oxq+AEcBhkFI8WkK91z5wxkJqOmTEHmm0M+Z4b0
0CJ3nordBOqmlmCTkl1BoUUlJBWJpLNI37aIOw1cO+fhTqNdtapxzmlT5pZqC48Q
uRZfNj5sHbe+XSJv3Ynjsc/j+v+rxMDXhoDX2gG+5imxqsKc61TBk4Fb7lYJSo90
qtRqsOJGYw/mEsrx6PigRVltw/RAyDtmOBTpYrU2m6y06Npjod69Sk0gJD9Rw+Kn
EysGtC6NXtC+GVnK4PGPXOYcjCCbbf7GbCymNEvXCfMXTN8r67RLDnxNN067lOvP
AMXCDEq1LK+ExMTc0hBtPnJcuCpGzXiQSVdUlwAF8QQU7Mu6ttHtopTSN4eBWYrY
lrHnBMkKAIjvu9ppPgwrVqIN4vGo+Yb0IawUMfgrzeATh5eSR8iNvNWbagt/UP8F
ULG7yv3lGs382AE2+QfyZncohvPjzQhn3V8ChWXmurhm55e2Mv5HLlwU4yvj6iUd
cQHOvEv1/XbGA2AG2JmhKE+ooDvI8pgp9GqSQM8fghj/AYpqDktnLC68lRlzMSVQ
f7VWkZfLCWFg2uYEp2KkilHzkzTe7Ljx0nfI7ut5a7sdjHVBW/YLpLJ+OBqWS2kh
2pFT3QfMS47gmxHqbOtiHHnZcbxMfMQzJiWAtbKqpE9AGnS7GBIblm5J19ZeH2te
jWoLPD8n2AE8ecze5hYny6aui6PVlbb92xgrpKs6oTkQm4A2CWzWciQOOYIuQm8C
870UbQfDcjf6lfw9lUoRyYEMR2zIkpycGDMX8rju6hDrn1T1CrR9QdNaWM1jGW0h
vYa1s2wTt6sl+fvB/dTv7j81KodfosERv7bpYso4eTmVVzNpJ2Gvt0yZMyw9MiL5
2z0XavWexW4+CPqPUMhrb6nAPUGranxCMOobh1rugjSy7c8Oi3osY5FxPEY+bGyU
tYvRx49tsdqvY1MqXKF62vTlEPk1Y+4Lgi4WSBPhxxUXYue1o+1rAx/be8U6XRzw
gvemFcT/aRmLICNT0NdbZtQqGPf2d85xLgfV/e0YlTtoW+rN6ZH4igCBOTtJJNgF
u0kxAc0TMacDZCmmjcYR+XLj1STVED7ojB7Fo9eWz9BNgjR4CiEQkTFtTZaaSLlR
QZdp0gM0ZjS881zQy5ezVvso6bmJZ7myiZfALczKwkHWRIAn/Zo6jvpk/5FXkp8X
y7F+z1OwU9JboRqOw+FBM77IZ1hO7ZESr7BqEfs7+hb3VF2YGE/eZnIIz1LCpOKt
N804ErqgJtluRQRXBtRS4+guMHP/4isqbsacPqzoH6OqXeHMDbUaY0UyBhgiMeC8
dtmAQiEafRVnHHGcSWAWre6oBmkFkjWcO3cTLhfuqwLlqrAT2SbjN+GrRonb3I2g
IRqyx4xXF//PZTRi0PafHJN5dad9rB3hAmHO/LEDU3dC2P9MWKbbtAkelnwHRqaA
yZ5RxWyHO8fXIFSzbcufHhclFD39MP8Eto8bYXI1mM2OmJ4gAnN1I4gTR7RAXUZC
yK+rM1EOsQkl3mawdStmVgcyiIOOqSb4itqptD5NOiOqoYUnMY37ytJHKiUGconN
RUqLAmNTHsaIIMMd4wdZdo1qKDs5gfpQubxFRaJQJGD9tTXu3L06u73KfXZQtSoS
6hvrXdI/I5uXzd+zHlc3MZrdCBAWBIem4asq39RBp2a3wM0NrvuhhCtndTeRp0GT
qf4nBkxiNbopmfAP/HMSbarvx4GBLpBX6xFsX4WdW8y1z3a81Sb13vEY41l7r18K
3VptkVCFewQY9317WJJum05VbM30tckZq1giPY+Z+ED7lYuxka8ycEh4gh1E4oxC
sFlrecsGqxYzlIWBF8Fu+2DO749smsVDdxvt9jUU0nqbvW6QkYy2xk6nCCRptEXd
Uf7Hv8/v/4J3UV0RL+UDto1VcfyI9JXvuWkM6T0xGuUs4ZLzkgS3TIEriWaFoErk
XD9GlwhJk3dE2SGkVWqb5BSyD1iNeJNy3cNUwcUXkwts0m7TqBi5JTHCI7U9DOe4
79oiPs496P58qiAmz4Fo52JNxUoTf3a/sLCU84K9A9M67gZg//6Ah9zzWjpONHEM
5UDwZndPJ91P6lqVPAbcU9xzMNMzBFQOJAh4Wgg7D7vSSCrJEGd2mtD7UNqnGngK
W171eMy15V0qmCwsYqxtxPllzMnQlSJOxwia3fMBmLzwCUHlaHrvVceRial1XQ6x
BXaBvr3bHTCXaVF1tpotx+3/OhhV3eSSS+bJxuqINjIcK3ZAiwi7P3UjhBHc6a0R
FpgknSCaYJA8OQwDsm/K/pa4fSROp65Avt4kN9t8N18s6nTg+jG+K70kaj8IqotB
Jyjr/oXOWbGuFAYPvSlzKZolFOrim9A6oSe67t62cQMyand6LBg7kzoqwWli11LW
9aDq81zkEy8/hdfAgW3coCKRQb4B8CyVhPP+on3TKV6fsduFLd706kmpAbuQeGat
XS7YxjqIeKopxRzkTgeLQtmTPvU9U9Sv51+4FBMR33l//+tzhOfCJiyeTtPHXALd
PCdDNOdSfqJACeHRGO5NohQ5kVmoFIrCOvz4W6GTcJuEoKlaEibAWnJMBuXxGM1M
cMprhvVS3iMRuRF7Nlppq51H2UDhmYaco9CrOySIbyso2UAghWyYFKJCR3sMbiNg
w7noI4rgEfmdb36aCvjvoZZU8n4dmOpQSfg1qWj65hVXd1MEelPd4yQlgUxqz+Pe
B6gxSIeOBizfLuPPNh8BaZd0Ov0Q+uQVUvV24HO2X9PnR73ltbPihRSkMDfav5kc
kVoqzw8do0mTZfgB6QMVNrL2I7Unt3CF+w0gHgu4WglEsqJGqCJRNBSWq899eUto
8efdW58rA0GF1cOOS3QbozuWLZMev8gfAOgWXCrvIyW/swTrDzzEFauv2X7FytRw
FjTUH1Bn4brxRrmuyzNv3Xsaztxc5aFWJXmEP40OZVQ+zS1KDLjUADSpPRdfSkhD
LOcGKbLDuzWjVMkA0dEjV951rNFOQQnv8OZNBykxSzGw/e+B2KXqKzcT+Ll0wD3A
sm15KTplsykLtF/uE1l3orWemjo2m8Q0JVDSnLXSZJzoQSTRVdpA9QtL97xhosRp
6SJom5AzlB1o3lNlpnNc+Yl2Kqqfn6qYZJjluTbJ4gbLtENDSIKo2eIHaqrI5+rM
fBD1+WMlY1oQmqwn9/Qs0jm6SMypZgFdcTKsHBcj1OIUUxIcRvB8+yOUmlEPnsCE
Pt8KezJ3NKM5ELHWbs22bN14waSzePZJzthlbc2e7QxeeKH+IQsHtsnHYXzE5F7a
SfLqAu4f5yC0TcSs4VxR49bocZuVK9tW06ICd5HjULYFo/XC6O6ffLZz+vCCuO4Y
s9KShQRczGKHApGhVRy1+4Ignq8kgfiFf/G2rHJ2aRSxYxgaqW8Roizrm2oF5fEN
YqAFsGpSFgxjiXtIyp1HBTKzqxf2tuRKFSIW5Li/KN+O5VNY5/tAbCZUU/wn+Se/
EWlMNgDwhXpZMlkZ1gP+KMRZmt/gUBcgHkBTDda4zC/NU/zFBPljOSginYTkuujX
n4/TLsBsCGQbZnEXVvR6Y6yW8MtbtYwPNpQjO2Omi4vo1U3WPnsmIutwIhZnYJUI
xu5bpj6azJuykYsRH9cnrNMgNrvzVmT7Nj4rFV1PUU0fzd7FLUDyZfMN0pGWa9y4
JeE3jX7G/vV3mdGjs7TZbBZmnt7ExydjpbuTGrJTLLwIUngXh8YuCcXBaJHapsfo
vDggn5G3DaQAdaOAD9+xAcTKiY9ySKFhTmOzFY6lZ7hRJcv3vKB1/HhdtvXC3P7V
lGDbXGzni8+36SqXf6/PanjvvmxfAaS7bSj6aAw+CkUPA1nIIW6qF8uqWsZKbraW
tom1YJptqmkcyZ/xEkix1VHLHQR5ZCkx/RthW4oJrPj3QcypqeCT88oZRrNJHhYU
o6lAJL5bpl4y1kS6IsTDnOIGBXVckLc29B2Gy+PF1XwQeOa7ub2+ywjXA/IJOCaT
/71rQ8EbDXe+miqIVhjBYCYD+1KCPFgk+BsMBgSBFRtbGqke0EDwmgZvpwvBR1bj
fwfFQTpIVtU+pZRn78IQCcHb/D6SRLGXyUgtFBZK0Seb00/37ttbqZixydqKFFKW
68n51+52DKSA6R/ZS/Xgum+j1aM3Kn/NEgtmJm+zfnsK5S9Y+QLB8/AR9gjTYXnQ
yoAH+/K0KQ27m+uH/pawLiI6BArcEs2Tgl8n54bAFJupt3AstQT1/KA2i/XLayN5
FYj0R1YPrlgByKQfKJJfNjjzKwNP7sXD9cXBoHLnk1ac4a0XcezhkZxgt4dSv70h
3xgqvHkQw0nw62JmSJcAivfmmaV1ZOro6bxeJZ0F617c5EhhzCXJ/l66gf6NNTJn
YGqOJJUX71gg9yCQkvm0Y8NU0BcB0bqhZjJqqB4NYVhdy0KDVx+Ndw/DW+kfIPTT
CH6degKfytD/bQtBv2CUxzIuqeKlTECS+8KYCvBLy/FUvXlqkuFL5u6xwsGvdZzR
0dDwOEHnX7i0NkL6Qd1vwDkfFWR7x+rSCwbKJ/WhYmingbFX4Q8Yzg8SIaVIgYum
Xu4I/vYJwojomkc1kPCyH9kVKtsrf3rpsWKIBUFL4CsiRwbH3BvMleGYYFxbu3vb
eD1gTda/WLMFwgelUID30MHC5v8N7M5BWnpxbLQVrOlEj5JDMGq8HsKHmHD7q1Dc
FlyI9t3FIxLF4rW4fZ4YqhNxP6pYP7MlZri8/eGP1FzF3I/QtgkEWTvp/777/UHP
jWPjCuHQGKcck0Udu5RgyogIqx0zPz2qz8SjjhSAu+6Bt0AGQQ2ZLOrICl8EG95d
l6LS7yT4bPH9fh4hp7otI6xRdS7qqS5hN0UAwrQY/qI3M1o7P0qIOWGrn+eA3BAN
Ro4i/+cwHZe7yhYcDMVbvgbu9hbzB8mAcgZjCx5BqmK8YpdgK9MxhWo7FwNQAALq
iH1Ok5b7Gvxhd1Q5LxMzY92yW9c6kYL5wgXnQ7GC39qvGSDBXLrue8f6wflnC686
47KQ5gD9mg4wMESS4LLOX4v1LAFXQuQIfPtEO22lyY4tcXfK2SKOQsg9f+PzRS8i
xhIQT5mVBcA8oXlar0x5UU0C5H7Vhj8CML4U19ccvdQeVrqz551e7UJ/cx9egrEt
DKoboWEdT1klADE4AzAK29o5IbyxrvZHKmF5MWmrawAdH1T1hOqOnG1+h3oH5fnP
6IBVu/VerbwWwgi1ttvS+4leCc+k04zrgQEf0fRY/EYsEGkXrKg3L7Y8rOsfpHXv
aF+90iFf8AFHiScm/mhWq2wCSKJhdLg3T1i6O8dkDHgGEM0yg4yQqa+iharPNpvT
5w/IaZYpfRn53TdyLcuVVw3P/s3H5vdLuiPn37ust+ji2rakf2wjU3UJqmd/AOoR
bFfihRzJ8waegcCkgcmqTHS5Hw41v01TumcqoY/FvJFYPOCOx2F4p5URqSAjvgq9
Wg314ztgjPgOaQYDCwKqw4+RHACtId9HKWNroRil4fS2S5FBGa4n3ojMk8ffw8iF
yQ/V1KHKOXOaRpt+T1XlnqUX5b8MSShzSSPIXhLOHfAECjZPv79p2/GVCuayor7a
q3Oyhtr9JRwP1yvjvEg5b92SDzVyj4bWdbh/i/j46tT7h7UhErZ8mbARl7eQoxNt
yDte0GKwEsbFWx5ssb+Qy6DLjJvXin6Kis6HL8zQZtIEznI0PDANbAffkb9QcWhB
/M4CqGxpFX6pd4ALOoghKBU5M6TqUOPcRc8wZ33AZkJl2Bnhg/onEFiwlU9Eqjw0
HBQCLB7O68QShy83wCzgxZhwfXwx036ce3twi9vBXSIbyDBH0uC3zb6OMLNC0NDv
9sQxOnhp2PXdpDGn58Q9Oyl+pDaVs7EOTUWsVjHaSW2Fa2341B+sW7z2oQf92d72
PAmQWoNWbLdNdRdDF8+90CCI/UQeHSr4ShdTMNy70BbnkRyyQo+G2j+nxPcFqcaU
0d9AwxIZuE93irBQ5cHwnyRFbLaj9AtaeALrGys7Lc4PtoKKkXsoZsFCqBhVUXEN
g9V6Ds8hW8msaAgO2QvWoqbJnKnBcK5BTKAwHa8fPy6dc7c2VVanakZNmABBUBZZ
/Adb74qXQPHqS+KihUlWVwVWBXLABc81QJ9LDppbUXIc/FB4kHBJ2r/OWKksygOD
K5V8DHYuNbQsfTLIuSmBGdP38+Tk2V+jGp1LRLiN389Z6qXGFbyrGY4ZlmE2F/sZ
kmqVvP/W+/z8egZJWma6fjh1e9+RAvivv+CNn9NUp1JBWDdkZlosyUUldioj03w5
M1QAIpqWXicGwgRrVRanzGnlHn18u5lziFVO/etuK8VLA0Vt1hibOAmyjAD6pMEC
eKHZ4fFISTrBsbaLyY54pcuiMM9jtCfTXKzbtbQPi8Jrn+yFkxqr4SosNrPnxpY9
OorFXBMboTDNFXQrXeacORpgjbaNS3143L9fmCuSOUz8olgSGbjLZZgLzmwQ7Pk+
2FyvPXDyFuLSjz7EsfZwHj7eKxYFIZgeAIiaDnzHewehfCmzKijj2KgYmHJaP+wQ
C2ehrkuZy2Wm58nsYOWV/TAEdNgBRejsyHf1kwy84cEpoCrjwN4xU2pvOR5GHJHq
ZVzbtVujexJGoKw9RXpvZPYZSKZLItYdrtSEsDnxFqIAnH4H2SyrHWUQn+gCj6cm
t9Md35U8a7klzfgUB33E70gUlc60V43Lb/NQ1/OZpuxdMKDr68ykuKePBey+GJcD
W6BKmbEsaBukJNFCZNjWNvoBAfVyFNt6Pj9/OKKQS6ne2gHb0+845FOWAnRyOYco
JEsJDw9yqQdIIFVnjsBpsgfj3JpYwDdg5SeTMEDW/EuAeDPo5tSQ1GReAhDjfEty
LNj7fA0BlqJmCVoyILOx+8sbODS/vji5jzbGk/XRC+PKIqxkvOIsyoPlH1B1+sdU
GC5s3qMc+l2MSymrwHDWsjg4oa+ST8QPnDnpM2zaw4XCivaGB7ipaF2pmDbXFhYw
a+BCWcJiurwgHoAySulnsqs8zBtEgEwUpucYu7ZMdrqjC/1ljDoU/v+p3NSfvd1x
oAk9FdeTt/+aaN7xFYDOX4g2uwpb368hr+nG3jztpEuvO5G15CWPba7POJZWHhBj
Z6/ebCJuhtpshJkzHvClLbuAVuASNBW0oM/0GNGCIDqGc57rgIcYBvcNaU6QmC6E
G5ULP7EExKThXK4RrpP/OAef3iwe8qG6w0USZxojQPJZBP7Z3MhCWMUietmJFNmL
2Q8oNtNXtslgNCce7spDXD9wodm5T8wA1+dLR15Ts2fye5mUoaU+2u55fBTcjgr2
0O2Ag/g3uPsGj6+N6LAuXviXmeKumIF5Kn/WZBMunQsU9W4kA19kfgF983D5ItKL
VzxqT3nV4rd39O6q3BtFH9umwwcyf8a0B2xAQYc+uDPNfGnIDbj1xswzQpOQ8k/C
JpRdm6kg/NaH8JezVoAiTrX/7mHYZ82/bSl35wiX6Gt1I96rd11xk0L8qreYKSDB
HKU0XjWx8CEDV+2YsckQBFTDfafYygqLIvqNTT0IaCWvN/Q+1dfG/Som6fiA6Gtr
YSbhPurSnUoutpPdrgRR1W5ins89mI2eSGJDxI8HqTm8fhz8zZX5/WffncWZb18m
I2ofvBN/RSvFyEf37LzAgCd4RTFyrvznm1wbaHqkqCEWIHshvhKubzrCeuApIeb0
BsOk8wglvN6r5L7EHebi2mgdRbMxixWr3tfTrjgemY9pS2Pzf4uAXJOTfebX5IV9
SFhznMoB4SwrxeGXFsJRoa3TdkxxC3dXmAqR1dNB72FhM0sXCUMQBP91l+2rAR6W
cI7sH4r9dsUynLokcsE2ySHeXourfxHhqlCMvFtJLt/WgVMtsA6ydFPl4dNkApBj
bOVQ8M7YME/BvNICbMo0bXKoyF4ySyPA1M9L7rW1zNlu9jQWM/DSYB0MmfF7XD3n
0pearfLQ7GacAZpDDWA8mDnr7VfZbNFYAXrZPIB2dNLS1fWTBmU95hLweLf+Bb0i
+W1oqkw2dbEien1Td9vgGX0NLZlUE/Ns8AeRmn8lQOOSFYgGqbNY0YrQywW3j6XH
naJ0x0vaQJCDXvg9hJpEY3OK3juJgOOcRHmMN5zWo+9TDOFnc0bbG1Iz7YpxsB2W
ZtIN+Z0Eaw7JGvkfW7mcJGaOXGtIs2AJBfgtt7w9BiJDGXXSDhwpKlGi/cn8jlDT
fRS9gqgtBvNaTPCO0v5D/f5H8lPhQuwwwdlrQUSG7h9ISEjRzLVj3LBQz/gYChT1
tsR799KIMj70O5dboCFRfl0P5VTAbfJhycTmzz87jxnWZMQ9FY8r+ijDSidR6Cuz
3bJV/w4M1Uh3o0iDDwcBiTpvXN/CJjuIe14oWtoSVSctDUtY1sDc95RMgl3p82Bd
gS4m6nOWt99yfNLcb2dMkvV9A6mcD0ALNv52Bi9SXnFYhtWUCgYmaNPwjnqTnQnn
z89z4KRQrdsePZYF6i63oSogZ+PgP+OmKH5SoSlBoRqWyTZ9KEK6TfqnkR6IxN2K
nUJCeeXNIW6Dml6yFNaGRR6zDkn5128ew/mXzhA5Gh1r7mx+Y4gOPM7+JqRNpUok
ffpW2xBRQMUThRYypR7hjiZEmV0N6W1RzARs13jRIPV7dkgn3h86nh7YBU9fn+Bf
+CB0JEvORP82wQmZbTGL8XF2LR9ptwgZtHDBNvNOBGvaRzfGn6fbQUcHGWwT4jCg
iyYezG9RFG20wXYq06NuK+O6cjCn8/DeBT2ApGLTzos51hvc2MhINJbHUMXQSKH7
+xXT3YTXky/9QLznSD2Ivehie4m2MXcZ2AWXAqqUXY0Iype+ixmlsWx6KRGAr7uD
Dq/rTjDuc1rPv7lPiPz2Vm48lmGUo4CW3axzvG2nPh6OFhGD/YE4C+oFH6Tf5Rw0
QWatb2MXH8JxQ1WrOzJH4nsv4oZ4hm7tLcZq/QfXgoJeu3tSCsYrGnDDot/JxYjV
Seuoy9TV1N/EyX4bPxXSkkdvSSHdw1cStHH9w3ru0s4945RlGiX0B1dUgUwd17s0
TqPxbQEb9zL6+3PIBSXgJ06BXnMdPNDFELE5jch39M1u+ljRkZTDHOUh7FVUhxxm
8g93d7C35AI9pc8v/99zpUYSLyBY6dmi6wPadGbn2t4g7RgBUR7gP4/vD3qeMbxX
E8SHMKxZJSHKPRm83uW71KIbM6sxJt4lIhddWe3e9OG0KBuE5sCBO5ZGCyCde6hD
oqby/D+t5EVPvm4G02NMNDcSfIpO2nD6v9/tuHy09cz2Zm0q3yRn93nqGEtVIK2r
1RsviK6x56wjvst+jK6fb0pCFX6kOOJQyd6dHwGjEpRx/Ley3rJA75WCP7sE3ptR
WsqbkWsmrlN7jikoaWmAJPbWqzZ5iFl+f3IGgTwDmbL+DbOhKb9eRsyu2FhXNdmL
2x6C7nDnseUWxfCC3KiAy8uqKJZn+iuNvNlEQ/HakaM8gyGZMwMHP9EEBMGyDTP2
oe81uuKazsvyvbrz37/OXjss7TBM/70kd/YY5048+8dBGmT0niNkjl/L2sNwK45G
NCv5o3oVRR2TgOcrcQ3s1oUmnPSi3a91ITYmlNBVytY3aZU4NhQ8Kp/ThJ9Q9fAN
p2A+CH7VONrY9quocMFkSRszgbVNV8Nty4tfoO+4tVR+1gmEDWbf0KA/ZnZ68qLs
wNexGfAlyAs+xrUKQhdIzsKUWPAq7/goz9IlNarlf7P0I4kSHlEO4LXLzdqwjq78
MsAsOuCTZ6wHuHC5AC4icH3ZppLL0tDz1j8roCL+dIepPYlPkb0scHzsl6MP+x12
G1UOnCjPyh11Q4jWifQZR6V+AZiuHOR/rjZg9afUqTIuCOUaTF2pGhsezaIX+rIG
Ih90j6n5hOr7PMS6JLFCaLBNa7RT04XTpfT0j91lCEkfvNBzrqfHZ777HhJGr/kt
Hl+QitQ101hLBw+AymeJrJzad5Fz4khY041kMrfPTyciPU3/vGDtbxoNBZtaP7CG
A68WBEWtjvUt5at5XsjpiI9fHO2T/bjuj1qxzu6SxS3L3fXvbwD6B5ru9R9sbSB1
n16Atv1tiFA72KPn1EsSLFlYX2M9sxxykOvxO07Ss4ZHWVKOPKarmseHQdQHbcNS
GuMNUzAuWmDau+Bn+INxZ9Lt9/a/y/NUaXsy40pQYdxWV/A3mlafNODxwN0G0rIj
k/7O4MlAJvLgxI7B909Ac8xJaBY5blwYe3jsv/zwGq6JFNlN5ElQegx+Ly6dPE+7
6EwLc/H/xyuHNDwIbF5Mxx9zxfTK3bnpePHH6jwJjj9TFfVjS90CDSoE0haGS4xW
8y09t4npdtO6xjUfJV5f4hFCviccBvtn0Xa0jujDOxb8za0T8dyQs1gCEFXQ1VMV
Xd7kPMbToKPGZen6+MicGSCVRkvQjvoVMUHjj/6cApnYhGHGHyK5NsdpugMbNEZS
l+KLgVM1T8DegMIWLsIuPjsm8nZCiy3E9yeWyuliyLa5xWsz8Nk/oaXcDCI9cHy3
PVeCMM/izYEB3PDQ/2bvMo9xKbGWpS4BPDYKHGjpvWYAvp8x71zfbfbyG1doGrPQ
ADZl64+y+LT1bdcK7UMurKJTwlCU/pDne1KRZfKMy5Nn3s6Sw/GCOtwWS06Ya/od
6Y1UtfP40AybXtFqae3MuzTHdMOqMcBmR5r7USpOXKOh4zJouOggNtzL7dCzBRba
xhD3XX9A8OiQjI3HPwDz8peHrvaNMVLXo7rxTpT8kwda0amq/8QbxkMgegR4scs6
ePoeC27plt6SDIrqL+VkiHNMsFCAB+AAdy8W1pjgEFyZh4N2RCT25xEMe87X1sRX
pzdWKz5zI6rQvjYuByw+SWZbdVxSUeDiEc0bINtapsG5CldoovX/4qyqQtGRXFAt
BJBKvN0emTALwptH39DqoPFSYiY0TZJJSI2IK99rWtVuQO0URmXv1UfC+pBM2WE9
hzpl69AsAjPsaE9texDXtzDrHIksxByszvc+2lbPdapehip92TRHQAFuFaJMRHi0
6q2GcP3uPqu2DeZyTNQMrL5Zu2060AKXcdiTfIF/FRa2wCuvT74pnKiV6xxEW0o+
Zqr9N3ANqSm+txP+dMgpgUTj82bKDsabgZGbVbB4lA3InhJd8WImvMIbZE5JZy04
55vsI/OQ/TVBGSwF/Ko/7DbZE+ey8ztjvzHo462FPSlp4dP9sfrDjMZPCrf82YYw
c5D8Z0UYWOX6sjhcyfh9pbYbCAG3/Pu7tlTNDnAJ7MksDGnVHXChyfHtIUAA4JXJ
MaFzBSFYDFpPte4Gi64p0hMKN1nW7kYPP5XclA20ItWp+UmYWu7Wq28qj8PiV6nB
VOK4e3PTDzjHSmW2Oc9+HDKPmu/enoHFoaVxz6wdBBIcppA09XW27tbipi2lTtgH
1e2fI56RtE6FlegJLrz7kee9WNS/apD4f2lJ/YvEyuemcgSfl0KfeURosZJK1lYI
aGXpfCqyj29a3We9AfzDE9rOw0Xx6Ro9kRKed3E+ce02tqL7mUX/0wNex9TlIWiB
mvavJL2A2HwpcRQfeEfymTGF+4fbAWC01S4S/Chjhm/pPtX2aOr7gunJp1NdiYVJ
3fs9UXnQTBzI/6bezDaiIdvFRHYEfVyxbWLwIvelgGn+JJNfaOQraSsts/mRHw82
vXLdbiCJEXo6i3BFnRx5yyoA4649+wJbx0yE/4u3LuilIfuJZcCmN4228guHVI4Y
Lnk50uSqpMVPyOY7UEXXp+3XUIfuac0npifVO95wtPfNiwV8kzGl/WKjC+hLQd4P
K+57KH5dL72H2dejg90olvdB3zkjjG4pmbvUrjv2MP28nrL3XBeRPXJIKXrO3moJ
XzRrt9U3qQgc0mwGKU/LbH0r1MTvOQ4clljGbiu6ara427uP9e8+Tcao7A5FKss5
RFXEMjCJYfi3BQqu160zJ2B1KKDhnpI8UW95eGBLs2a3po1zY+OLqnyQl3bIjpaI
EzFDaIcoZF0Cq9iu/FpvRxdzbWIL+jfHbW44HwwDGhdKBmQ0XvN+QDT4WpimVcua
KevbS45AdvB9u1vqqUsUkI+Ux9hG8v7pAneyuvAql6ft3+w4In6IETDwtrFhYMn2
v+AiIESNKJZpJKxO5OB5khqTF2TehOSBWh+STD1+mPVavg1IEgZYhgwtCq/d0OIU
tgdKCkWOldxaSAMiMHTPAlWjjUlVh++hsZZoFFmpo4hIrrM3ugR89CLeXSTvu//x
d8GxkxmkUoD8gEB53MlVLQxLL51sfKle3UMsUBcn0zjzjgRbgRlX1yA7flGyjWtd
ZDtV5H6YfOcsBO766qOMrki9w1zQQeUTog3pLm1PIE1KTDvYpcY2WaRU2suXe9Gc
mRUgJyt6LBhjHa8eXhFoZzRR0knOmJnpCfxk6deY4gpJoDNG62cxe4gEKbTfkt61
PnOsM8lT0zw/ZV4EOcjRU/zVUCq3qBe0FijLJcruAto9J6Zo5KKNOGYYsqteJ3rX
lmvoNdr0OmwFI7Ec8euDW4iJVxLGe31H2AXu1635+0fQnNHvUmwFJx/02x+m+2L4
VeHEi07Rm1H6C2CKF8Cou6AEofEt/Fvpr1AUKyvUrgwmGenD4unLh50nPItbX/QP
H1PsCMn9/VeHsw4mB0KrybJSK6bDcnw6SmQqM1JyI7mYltJX9hZYezNAalsOj2tG
SLbErKJtjijI+mOQEjMQlIVgw5YrEluRXvMT33HAQE+lCesCJy8rzBpNaDiXZ9V7
V2oTePKHqLc3wgUkg/6IRbOgbPQwNItUbwzBULvo10WY0E9zhfi81yIH/vv9cfxV
sDM21mZTusyT2I5OTIHUz0TEhVMZDjf3MdGLr85B9lFZf3nTu2LTxWfO990njdAk
3qNAbnpJeE2HGvNghvWJms670ncA9dq42pKF/tTLZAV5N4ocOCAYIUxrfL818n78
7V/J8h0kCNafYWoCFmihHoHcczTGBVocvjWBb9AapqrahxgUg2dWtoaQz9xf+uxb
dsmfQlWvFxpmAfzTssfdldnROyluKqrZUKGPi67nqHcqv4IH5RSbEyCAl4vW369Y
6jIlNmJVAD5mxSsBq0Mo9l6CBdMRypaoJe47pFknaY/07ZF/tmzXoRvGlb8RJfGN
Y93/jdNvM/D8FXjDDZ1fMEWM/aerzl1yukrWXolkqWWvyvNlHvWp+sS46feO/6QI
Ca4yKicSZi8Is/1RIKoHbCkwhsK8Oe26qTt1wt0rFxofuiI3mHisRHt9WrjuAXXx
3h2m1ZgEmKETSuQaxPxZm55ya2euonXveURj2/7GN2YOV8zI417s8o3SN3IwU2mQ
`protect end_protected