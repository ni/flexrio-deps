`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11488 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
HDP29p0vLOrNPcWDOvry+QGQycL58Zcbd2zJPqd4XNGls5Ix2HYAqpWQiSMQe8f9
8ZwMuLmfXZGRYMEEsJ/lZ4ZYbbtlgxZWwPQuwpKuXnUpCo5heDIEIxF3orwOqZYX
0fU6P4dQF/0HgrcZAWOhJCPa9V7uCaQX3BtVWxD4g412nuahV+nc0DjqpV8pPOtq
OSr+DXJRyo1OT+ngCnqIW05kCQtjtseWQwWiCSg1qaHk0ZcUUEIG2UqzzDnskZXm
54ycuUbTfmSOIbQvJ1WkGq6RhF+WpyPGonnog3ZuTYlSwzlv0eun57QbOiUmrV+3
DALKAgGl4yW3mGWuBF8wB5eGpj5dKgold3PDnHFAbEuqOUREOqk+HRpeqebLYlcl
4HScTFVz4eCZESws3n7oYx/zGBpbaFaS3e54gY18Cn/kyuND1I4maSQxCzQuyxXf
xoF5h92KnktwzP8yu2+jGvi9W907cdZdg+H7dhbJM2hMIG6dBEVGdhevVEVYhW2M
NTXlijVU+0PAuxBa8qjPV/j7PKNpApyJA5u2OouWtMERof8vFvXQMbzsEleezUBs
LX5zkngn4we7AF1W1A6lx3FkUxIR24uX1x+JJMSdFlK5UvlDk8Z9Xba/0FJCtXd7
c7sl4R/rwD9DlJ+w8RZ++qCEcr3ii4/8XQWniQA64RzgoegtH8lRRDH+N2qnixOY
rEhHW+CQKbaFyAN2j9ARWRiCpiZWcPzM8SN7IIvjPoV0pwd0sIFWN3i7Z1Kz6mgt
T70HlkaiGVVzi2eZby7lxBkDHNJ+9iFKhw/oLF/Mjci0OODXhALtyjrslXPADB9S
z2gU07lyKo2AusqplWnBDGcekaDFEnEv5wC9CFQed7QHGbPm7P+Li4SJsA0XiRE3
a2DguNG052AfRHGpqNC/Q4bjLBVGHM0CqN59YwN8aEzJAL6Wkb3Uf4+IWXXCcCxd
ilSWZKjI09KpmFjZmds3Pf1twCxCAmXrSdNRRg+2KPAiFlFHvKPzPYNwUgsxDdu7
QE5gI/cpVAvnk8+NHupxRfRYdINES2K8hm9xGrAF/1b+zMjVj7HcaL4ghKWGPbwM
2gNrucKR79bBiucLiFWXsAl3BwL7HehiOMych6iQetU3a16Xd0y9aPIU+ciOfwuk
+DWldx6MUSukieUHt9EVdTvN1Q13SYePBR6W8DeCn2HRCXk55wAl3qrdfvCPW9+X
AgKnbtizrZYeWKT8HDbduUqnWvmhhyh+UIgnxHPxi6OJZxlW1Iq+dKFFJuyxOKf+
0j1GAOgC7GYmYmIjwNdUKJ5DizczAhBvgEHtugeETNddVAciQoxL4H8zCYWcan4u
phO3MFW8y3cO9JcMO/UrkLv48YVnSztyUW7a1pJn8txrNptRZd627SzHfzswBcm9
yjduoYwCDNkvaCkBjmWtgXC58YjhSDi8lYFN5XGzQaEKi+n/wfRVbRLCC3nkUk6R
5YWGUclFNEuXiL4JurAShxP5n+0UCCngznqDIeQmIMZhyjPSKvr+e5ZNnz3dmHDt
AgL+OO0xxpzHEjv+USkFHDr8j/sDS6PM2Te6+D9pYrHqSE7nu/XZ2V4yhnGPqWBo
Gu0TrOU6uV2qDEWCZhpLXCanDbLjGmlNXYxFr1yT5JjfPufK4kdLyB6ejoBU6oCU
jFKG4cUmdGY1TR0oCD4brzCl637sFx9Iq+3b2GlZzoKo10TT+2T41f2h7nug7npS
d3O6hWiEJcT3gx4c1A1yNIPyXXJ7VMajlFfQU29k41nLClVzJk/ff4uykqfr7yeb
Hd4mcC6V+3Z2IiTcteUkac+K3lP8DZhUfG3YYWfO4S9G9jMLCbLO53eZ8wWXSZH1
dt1Ug7ZH00EILdIryMdMAreKY8k73rrORqGM5cNYr2amd1Sc5CJzWzMTLYCbd+dD
LqG37My+Hu8vXoFjPEzTlkCyWFN36Sdhx4rAh4DK+OujccFip0S0ICxmUXXjoaPd
U8+btq1e5/KFIOEq7kGLbyin+TEk/HSv1MPhoGyPBy6CvKALq36tjm3KiFCLzYRZ
gEJfre5WFR79cCXIYyCGhtP87DSGs5arWczG8T63/zMncbskzP7Rm+fI494cmMw5
lstPLR1CR/r43xOGzJPSqxqAj5Pgm0tiw5k4c8lCEkYJdvPxSdYeCgZ3eP4KMUY/
Hhl1lBCDnwkGwPozI3+X7yTOtbZbkVcIt7cxE29nU1umpxpOarS4gsGGglDKH61v
fxlZVIjGkqdEKKHoYuWhs71GGpj/yH0X9frN7mANEawZ1WLBlre8DjZ9Hw8TWIeh
oBi6sHC9xItZPUH0KbmOomf6tcc/XgILyrdPotB2dxC/7tc2PV+Ffb0wHZwPUc5W
p+eTn5GypfjCL4m1YlFCX0diFKRy60LPYJEGJ73aK+2pOAkbCYg9wENmcNOZEHH0
oFPRzUUSO7FqpMz+9SnPIGke0poe3OqkRIosH2sQ4+I/NYBKfh66eLL3i4tH/kUH
+H8Q8a9v38BtbRrpFn0TouB51VWYGK437nV/crlGiLVh20pXwvo4DncLrRjV+1gk
OVMYbtHI27E7EvtGrjaFoMrTCR1ngbP5Fb4weOTO7wR9Wro+mtlicSN9nXhNYUsr
++CGGL8wM34FvTN2/m5MLHt2gv4AdFjRj5pfX32Xslm0IHuNvROKHIKd+JZAjw3P
YR/u6Bv5xR/IR/AzuJF4nlvhbI/OLcFxoy73PpbCkCh7l4K0U1BfxFdZmsmy5elR
6BUrPc5XnrwqpvdC0VWQ5xexXvarpZzFYYQeOhgg0zdo2VQIDrgYSHAQXiCxwJoZ
xTzFak+RPczrxZTwDOv96Wrf9N9tIeJVyKXe6zcxIf0sEseL7DsmKKjXDq46Y0i9
slEh15FlU/bfWI1jKANJgxqPF6r3WhAnTsvNVz68VrLOgnd615yHJk7ljT7k72YS
4N4HcJaVTpGemPJXGXJHGLIW3dWXQoKJK7gmNImpc0hp3AIMEMz8w4RVJjtc1We1
5aDk+4gW2+YTQYJZ6dqDd69OkwZQd+OhcmJq8P3cy44luFgJIlaIon1VkOwS6yV7
lopJX0nNZaIA7AREvrvjjn6Ur36vqOMw4DgOdWqImZogsgwUBtb6i699mF/k6yYO
EMgfkV4M1pdGE13nas7fBSY4Q2gQbd17E9/5iE3TSEg2Jar7t2Oa8iVWl6EYDCJ/
fWddpkNEPPshuNgI+icsLKEXzp1yc/EKcEuwNw8eP6BTM5aG0k8NbZJJ0VnGSCUG
fxl4ihvdciZMKfCppOeBlj9LoG+WNSphfHopBTaXKvxZPnR+fyWf4To1ReYZvcrO
s5rqY/W2RDO4+KEXnmqQKU6ZJ/XK29jASzanWRrgjhPRW+UTGm6KbVSDBm0OxjQM
CErGV4SKTiIbHVLFGdhInLxEzBDj3e3PHlGPFbNcN7EGXHnclTmvf7B7Xv6S//fR
GnflPsmB8xjNJTu5WPoA60luo0s5mQDSPp864+nvyMKoxoIDC0I1fLHpiy+D1GTN
DHQEVUdQnyI/HUasdxyHWND6m76xR/tzofcQfORBfh1nvRoZJBmW8+QNnOC/rYl/
rGf0BQXKciMFYgMwWFaS1kePrzBgXsJ5VFjuYTUlKqMmrlzW8/cbjphzdfaQ1Ufu
fEXDDC16BQB7IBwdHhXycbrpAtIanl/dwmi2IbmZcT3iz/HgUAxpX/6rL/wkz9Wb
oFNpMV97ehJB1kY1z2kT4bknIVFXHl5QhK538gGZF2ZAlsRvK4BmyXZK6BHiyFR7
vCqrQIw+kvm1rJH+TBJC5uZt40DO5ZDDExh17I0PXEvNDKsCN7BicPdpdm4X50WU
c6nlcZU8b7d8RjUK9nCX0llo0lOsc8H1mGps94xVnwyBUlhqPRwJO1rz3k6kW2ee
Zj9773cGX++bRU7bVo8kSYr7ulfBmLgKPM5KWiAG1stuM7Gbci3+3gkb9Pvd0or4
hIpVF1l4J974IFLOaOPYSSU2qXAf80H0Hc3cA9zapmzgsmKc5IauJa/pXNKRYn/z
7Vkb2H3le8iqfnqXMHflPqXP5RkjaYVHuUGmSh5jLEblSjT5/ZSaO9n7Hr9Uxiyx
3teOL7y8OFJ4zb95BK3o7p97oy8UZGapnAxlTDA2ZJNppEzYachPpap80UWsJvRd
73VSvGpfIoNqcDIj07tBUsRSmHJ2dLpYTtQUfAnW2JKN0U6q96JdqiwRZrrOMMa2
nY1J5IaohxBGg9SuvnzykCbaaOJ/W/m3tQgZ2UpjhcRoR5UFp+H7tDfYa5O2mtJE
jUQWJh47+qPWdK9tUs4nbrg2SnJhCJ9iR5E4A6qufIBFoD6Q1mzZNlhaI5jvpd6G
igNB5L+cD9A+zkKIrkzcdZjcK60oKzQllJX1msZPXalt81/JoQ6APZZWIlsuR3yX
dg/6pkpv4ZZc/DqfU9DPX9sZkExNfk6ViFJPcOTAXvRMDlzb12c4oI9VfHI2Y9Fg
BcuQZUFHrDyoKF70pMZmLJ53o872UBwjVZVsQLz96/VYqIgAmdyfP4itdOee5M0n
JIzKzwfiWoQMab4rYcM0tUEZXYPfeSeQLBwF5wVyH/CXialDHiA+dVSWV8UO/1L7
6YWRZj77MMqOZyXdF3O0fMJwkCoAH3qkczrjSqo9jqI3lJYZSDR6RGb7vVlJQA8T
JdskwbTbmpqp4nxHAO3dqSwJL+YoZ7RoSQUxXCI8PO7fzoNbfR9yfbJBreZcJ5vx
N9977+HBOOJj5ufdOKFb+ydeXELXlvqxdThxx6hMqIjQd0gDj0m96emS7/qzpcvu
JXlKeT7rzjqgBJib/DiFboJ2Cjo6icjHyF0WD+KrSDovU2XFLjFybsta25GVhCTe
UdtqBm3T6z9T8sK+oeEZ9cgmJI8VBJXFlHplNYRwih+KV29Om7RbUxBkUMxRO09l
vLU6LlfC6He2aibyNOEiaxkF44pJt/A2AD/Jq2M6bN+RJ9a7yYvEceVwkTm1OgQw
v+DWNqxS5cPB1m6UMDbmb77RKk+uLDb2QHCV3u77aIDOEDnBpADxcqz+WCHLHfkZ
p4QJVSWs5rAMOz/mxRA8EvZQizkc6Qjdv4jJFLN0YDKlNzKHzDy8lju+i7AkOH5G
DL6TO23q3RRpcPndr6pILViP7RLYRA33Ro37jcV4ejjtPNd1rCtS8IbPPb8LzwV/
RFoCROuMSPN4Muy6NlV1L9h1SolxPUHUqs8nABe1+0FCuzxFjt2dGIFMBDyAZvHG
XxXQcypxPP3awI9rEyV2eFpZ3ksvaJLG6W+UlGKLl1NlBJXLgtRbQLhT/J65D2Bs
9lfuIS5VHp8f64y1y1f8PYHu4tVRTD2f8r0HPPOdZ6hlQ0k1aHKp5sUmTCjaTTVu
FamFMyjU+83WWIgMF5WD0byK+xoMqu3AbVSWn0hyqOa1sB2AyEup0Sbg6bPZI4xT
4YdHM8xiTPfXY1W/i+amJBzn1fhBxgSBHPthUjATWTEB3533il6jWy/YC+Q+a8av
EVpXnRjfm4BtgKgFtmYSWf3IyFcAR9YbiOKPHTprbCZypQnbtDz56ir0coFgLvNe
pESTj3Plp6moPPftdi4p8ZEWSjJZr2be6ry9l0ASyqrNRz6lJfPP0IOrnK4aaw5n
ZrukdyN5NpJVpFmi0bfUXZPXjUvQo695U83idIlok1y7XsLJr/cloHalVnWov3cJ
WeYJw9VOsi7CpYqvhWsWnmZOmbMMkwd3SKobYVI43Ugxb1bzlbh+xYYlmNYjKxVw
FvcwQldFEw4SZ0mpNOlNVQoNab3AOmFuRrIpKwzI9HipXrWClfsdV26jyedIXsv0
fLC/1zYWzDNwmMv/sz04Q9sCo2vOHhiCqgyjKOg4k8u/lybvtCOAOeExVtY19up2
x+6rIoIQeIyH/xfphnsPoAT6THDedsyEkDGYl1DSneUlrapqyVV5WPzrYwJ28p3W
Fn61dge+zdMPbdFdLD/6KcA9JgdjpSR5ZRv7QumbKzljCtB8TF6NjO/Ic1SoS1/h
FgV1LFx7eQ9sY6EmFU7n/ur7OdseSzMOzFybCtSzlvG4LE9qgjywoNqUD2kRbeTN
RthfH6dTol25LX2h+YT9oo5sz82Ny2NURAaASl2ToDotDSAqk7U8ZwSJTxJOU3i9
rI99MIRcZCB3ONab0GuR65Iae2HcvQR07KejVKe5Oz1tzD1rd9g2NXuwPzXPGiDA
kf82LhkhsHJtGOhjU/53m1mXeZ1RXc5XlLmuQYuk0yAVJsabbbESom+BLzdm3k39
gYU0Me9ZEsn82y38Z6tD0e5CDkHNqFqYBdOlVzA/647mtlFrowh36OJe9u07+fLu
nEb1FHZWLXdvBxe1P+lf84MF3SHFpa6v8S1Rh6fBxeYBkYtOAX6DEXrA6cu01aaQ
67xTf9WWJ11iHgnTSQ7CzdCn55EsNirONdsX1cntEoR7gmYLwdGvGvl1bDOSiGOi
vjrc3upzl0nFtzJTvxQgSnDxmA87FNJ1bNQKRE1VEgZZ7dz+fRGyUQiXtnkQ8VfY
kL2q3IagWuAUpBVz1O7WmiKUY4Z7AAE7dIbDUO+ir6sHX4sGc+UwLX1V6V2KlNRL
BTTQE6HDO9GvgZG5vNFyF2tz1d0SX30aX4lDAKgMxAGbth7H4gIQewaPrljJKrQe
MeU/C5W1UrRZ0b36mPrhHjxXL5eufkMDkOO1oDFAsNRFXj17uXzfMcYK2LCsfElH
/SEyQCwFHYsdOpp8ncqkmbt86y6gTZKNnyBbhFigKjVaxDDFoSSHAX4Ai4bSbBt2
S2GanlGBfF+QvFGiay1IH175kWy8DLSAvHpe8JboO8UuwIVNwnsRMnyovKhtYoki
3PCccwMVSjLRUNsBkH4x3woQrR+flWl8wBzGufctzoKmZHx7D1U0PzgzNERaeI3E
11KKr/0xXdbmxVPY9ncZx/LBG1hhbtwYCtvIj7qCp5saQfDqIi9bGvtjgmYMvJCD
cWyHy1BuzT54wtlr0Cxan1Dom4J6Ae9dvof2G7kX9Og0QsfWIqYksRTpm1hK4t+Y
leGn7RXmxWf2Xuy1fCyqeDfov/wQNSP7MJElI/gmPP+s9Q0JP1piBwJ3iMEITfm+
KOHjQzQFzthQnLgN/LX88S+OQhp1dLPaG4mHt3eka4VjljlRSDsjYpsSgwIGagrH
YjPx0WlVAyrcLwDf7zrB0j7s/aLB64edWS/tS0Q1QX2gIStxzF1WS7CHBpAgpjON
erf9TsLBbBIYsuRG+DzxQ5d1yhw6+6cgvgpYO850TC7apCSteNgbg+JauaKzUrdI
DZ8CT8x/uz1s07KEwxvpt7uRTdqQ08z5wbIQCun83QAIQl+YMtTTxb6BLUreoq3B
DgezskBLp78xOtrHHmQ/dOw8GzN1jOJ/rM8GBoIsovPW3DVDqSCt9gTLDQbqmFI/
TgLjmIBROUTKNaTXw9Yzq9qPuWlLlD0JOti13CDHOJ9y/HKlRajQzoTQ5jPDuKlX
5TGuODqA0rCsHMEcXro0mYZGxfX2hlzlaG7/vOUDq/A7q/EwhJmZkjLJNh6wX/Wj
tpASozPnKy818TZjmZSYJ+Fak51pq5Joxg7omZICQ7ra+UqpOx93jW/ipaQctuzY
z73kUyGtiseFHkjY4JhLLezfaJXOm4kj0CX+JIuHfMF09LOtWg8D/IWES1+l6bx/
F8HF1Jc+UQEYK8jaOJymP/wdIrwC9K+lXU4/EKgJFDp3UyxuW5wWiBsKpMJYFZO2
uw3sWos/DrhybhC9AzKVxWfB68IE9B4xAZePRTwSpJS4uWKmTqR6B3X1zllncizO
IIezTlIT/O8+dZrvozP1RdYscywoe9F85Uw55CgNCqjD7uscg6mADfmAN9NiRudK
FqWK3085EejUQkdkuOJtmYmnfsBidREUFhgVFH++LTG43koqnmRXBg89IstNakqS
DuYixY6OKeDbZciCjhWJgMg74CRtcm7YxGvRN1IttMY+21R+/stZUFX8ZcM3RERP
go8ii7OpY+SQGyWkRY4T6NxlWv2BLVvrZj9yHYlT9w6IjfbWfbMMWXM4EkhYw+iZ
zhXytbOWH4Ktag3KIRre3T1XRVbDHcrAT+5CDqcI1NYu/2PdgKeO9zat+itQk1tw
LJAxBqqT78vGVDAbUx/++d4RhguRW1ezWpTxn8uH/8Vo/elhcDdNQdsFOpjtQlWS
n0AnXIQ+2vzA/zRljsf87W4MjnlkGVJhXTjWU8vnpmzWK+MxnGJAVCTVWzNug0A2
Qp/+m/5JUETSt1JHAxOQvidMjICVJJWh6UcnYyW86VCY9zYPqkY1UEG5ijpyrwIi
PP2r1e6YrzAKQIDyydmT/kjxssVaiyfOrVmNYLrECcSHEOl5XKUv8Zn9s6qrbXpl
oMrm+QMtE5OiC3tJwF5PpR+GNvNSleTNB08zUseJHLGG7uDQvlKdIL0ApudQq04L
ZhZ5osjslJt4m7Hz9tGpWNhNH5NpARSq8UknzolNVDr1BXMbZpgVhyOzvZ6w5ciL
nYCBZdPxGVng4lyUtHILQ5ti+cqb670vr42TtC2e6BO5MoDoQq5G+gjgQQ6+uJrJ
IVCuZ8Xs/uL+SV/YW3Ao5u0dfDHE2t/VqPlyCZgRu0If9alVqlUqAsM2Chl883gA
51Jr0IQO+GS2IknWJjZxdMk+sVQDPbJRqsBjDQWERD85lPKVOqF+jFlBDu9g1G4Z
AeC2xIwHQelZuTBYpGU3y5NFfkQqji6z2ExFJBAxymL01qJKCA1FKj25cojHdTlm
RYYOAzfyg2S3raSp2wkLBuA3gRYt971lj7WJx7cAhZS1+okAA557SZ78i92Ks0cg
F0ZpfJ3Dr3SaERsS5zsjlNjw8rBHOAa4b7SpYkpygYHGE2BDI07p9DTcdLSDKYUs
lhJ6zxZUOQmT+Vt1O7KDPy2x09xltZLs3ZMPcjQr6cXPfzq8Uv6N/CzJVsbSyQNP
MOOD4mMPjSVVvnigYLGp6kYEyAN5Zwh9RpwguWRpRp8h37xA83+oW+KAfxMIJHHq
aojSsIQ5dEDPXXWY6N1U2+ogx5+IghRN738+6Jvj8DvgXScj64jIOPP2mphOswUK
hxxCHw5knxNFeVUg3w931sZuLYfq1hRjjgxYCx3j8sFG42EJ0nqeTfy8e0hAF3O4
f5OpMqEHJEXOx2ndAMwGTLwvtmd6oSABVWVpjwmdxjV9W/4CzisDkyncFiErhn1A
+R82CWC6VZ8FBR2o6U/IAjjQv+3SOwnuKOZFKlQEYQ5m3Ydp/rXfokDAqi6f8lbB
Hwu+NyC1AjdP7U10TJd9guEP9BKDuqtx0LcwFhp1/4Y1x71X5Wcb7rYeLOaLgJlH
CDcKi5KgpOKurzNfvjoNgbdJ4rDmBxo7PwQGfmZ0o0BM4lzqra9QzWvKRUWvnjtk
e4PQR5V0q4WIhO/Nl15vufy0A0lbFxvV1Df6ei4jqlw2icTpJlYw8U3PIb4+pPIo
U0BYPE9gP1YW0g/d3wRknuVxbUqDfagdmyFF4CQ1BCVWBKr/rdA3iqEHz37ix0g4
VYqKUre9l0IL39TUiz7arEQYVZIonlUADIcZgLPReFHcmWZ4+IkGZ5RpC6iEWDml
G0Lbp36JDSVSHPbnMPzSTgV4+O/SUFhPiUTOMps1kZwAaiBtYrtqsrBaX5gZbASk
N1mvuDSrkRW33fjqHqh2F4bGij3TSosKTQBI3E4BiIc6CKSehoc+L3Sgce7tfTUg
FmtxPz7+1ehvayxfr69Gqel5262xGEKPlSeRBypE/GiQkauIIfyGiavmfEDK0Fh+
pAFTzQShTXwKQCUJanmv4Z8PXmI9bHtsxfbcu9trI8hbNaWm5RO74P9+bHpUokc4
L86lrZA5EYGvs1QOpqRABwqSS/e+/a25EgcJ1Siq87ffTxqSQDmY8ViOT/Qc1bTQ
99+eGkHN8cfvrG4z4dcNz5w1T/ZlJlzru2bYSHf4IHgmKKSU2L12/VWGafyy/eyH
k8Z/lDRk6SAJVxHikoREABjiC7WdKQ5uZsUnqxuerdThKfIE0xlA58t0q9YjaXUj
2D9/G/i68qBW+3+xKIdeDdGD4NQs7FWFQ+7ySAlsVFQAM4vMhKMX9uBLtOqNvDMP
3ITO7HIzifUf882TuikekyxRL8ycJzeuBHZsQ4d9hqubMvg9wOxmofOlJniW5m+K
9iX4fh43IumeOEaaFV81af8QJJ83oXzNdQ6gicJdjQCpZq1F3UnSQHoKurJrKtPq
cNWZf+w+1LN2atm+pvJqqq+BZLGo2qLuQZ6HxulCpaVsUjV7ugZMmJNspTdRAn/A
ek7bPzcC7uA/0DF88HL/HiHjypbXZG7tLVDvWWjZAtrpfmz6B8pPIVPt5qqQc/wC
OE3LzPwyHj3xzY9sOvIa92XOd7k76UdCl7olv+bsHs5Z2yHo9RkdAAwqq6qQChVi
yDY6SUpqd+Y/+/9LuoiWpZhPnINbIifH9fdnriSmVaSuIYZVrSxspaWSXm7EKGMv
Fz3WBDyuOrcDab0ku6tKAqRTwqJQnTwxy+REdzBm8i6KXOJHMngsLrALwWwLUqh/
mgkp1PW24zuXBhIGFYBQTBT9l72mB2ViqfaHT8vBFau5FhzR6+s9uXKjF6uqpTnD
4/TyrTpWfSGCQFrmsJ+Y6fTG44plfKKXFlzfnNzNJ5Ev2x0A92u6JU1TWA/uf1Cj
8uL9xRTQVG3fZ3ip7CHx/taUUm9q7mXMEjISLp36YKoUfVPt8SJzeauj0dTUsOiL
wnHlb3C2PWGYbvZvc+fPgPCNVtN7eZaJ5klt1TK5ZtbARgvzaG/SDTJeKJmQMwUD
On3Ln4RpdIPgzduO9lIDiwiB7KpH2vv7VSkDInfdM99rB9ph/Wb3U+cTpIbTsiBt
E7BHAlt6Rw3MSDOFFohRbGIue/h1TzUkdfFVMCPxG20aftku+1gUj5gObyqLUzKS
Cz+lWvskFB/Pwh0gpTirwZHWADVWpZK1voWRSBFqt4fYWPS/5RJ1VYbTvX1uTJxP
XwzwzrlKsijdqEL6RRp3kbfYvtSvFkQ1k07sGydaZkAZ9wdAua4tujBVlzdntnK3
0rZsjlRRHvMGo2xoFM8J+7djFnapfwsNNX6Rt7yBzv1hxVON1ci5fg8f9KgyXQMV
gPqkuhrLV2kf/IJje3ZaF/+NgkUYcPc26KwjkCtvJUTMORW/1UdCqs89spWRoL+b
GD4+IW/tiiv9z1lFwNVt3U2hYuHnjVQobQKFwyWMdBkuMW1zN8Kll+h7qi6jPS56
HsHWRAAgHC6YIek61eCX3LSmN4BZCUvgi+5L3Ef21NuRcFNcLbpY5c7jaHTak2t4
R8Y+yMR2sXSSajfexYaau8sgSjU4Y+W+Y+NZ69/BINrxHqpbcp5jWSacK+4TH2W+
ukSiJYDyvhzYbx8ue0ZIFC2H/+Ov16upapqGwOYv9I2fDE8oriDqUgA5fNoQv1RL
UC3C8MxgbgLXS5JkEIYUl49eNW2LTiivP6PUSX0Dxjp3vNnYKAwXlijjARQCdVQi
cG7rVbWzu8QtpV5rzN+z20KOeVWFdDk2p/QfLqdaVK55LZluSc+K23eh9Lj0Ajrs
tNoQ7XxEo7YnYrIS6m132gXFgsZ3C4kuDgCZjaPrFJi+8iEMjAQ6qYUEKtJ67cEl
JHW9EwDP58BTX5hevrssM+7QQ7PWA7X/ILCcYz1899mF3bfiKwwLv3eP+10YTmT0
m895ur34OAs+Zkc0fc8ZL4Cn6prbwd7wv48oceTEmX9z/PiYE5hFREvx49ejTgij
hw+Pv+RLbzbIsKj3N7pvEj+QTdoGUJxJ+JavCIpTPf5N7H2Jrjzi8xr7yC6hkqe5
+pv1hGCtZigRI5VRAcAhQ7E+YKHoQhuoduxPylHfwIFOuBnSQfEgi2+I8tS/zlVS
TadJrZaxZrv76iiiDDWivsd7DAT2KKIwrN/LCW7vF87hy/ajJXF8HGwjfEPZWyK3
rQ7jCnj3aTbeizWsOCZkgnY2Q8O0lxALUgIIpF4nPxv983lovzdi22vbpkmiaGSI
NKvZRS5v+Tm9bzOAjSpcekE01mHF089rjDcy78ZXWPhhDELVR0FJlhKL9TaCZPyj
TrjViCSUhxL1QhNzFgeqq79qTTV6nRY52G+BGWr20T/JHG0QWx/1SDMVfydYpH1L
wTVpovm8CEDxT1bfk56C6kiQ2S090WxRjbA29FwiiudvjZqRIUEq6W8QSFehDoUk
B1rHlyZT8YgXG85iIAhVs06rQfIneUUTEPyvS/0wzNyX4UJvLDv5bBbm4zEY9XlF
5rx3op4GTdya8S3Jqjrs+JFSbKWMER88RlFZ8637ae4vLHvl5Vpl836neZbo/aIk
gE6FKpPOUXedbfovz1r87JI1LuH5e76preUcT0a/LhC6WNGUSZzOu3436abyHr2+
s/C8VTlC1lqhof3rxf3qXHBJ/Y4LCbWY2Gx7FIS2Fw4dWqwn+AiCCu/FDkFHySGh
fL59+L29GLXFyTMb9DhbUQONDO68us/lbo1yCqRJUmYglBknwIseGkPeZAVxXQNR
mrEpF99ir/jM9ev/UIsdlZUNnXbb95Hjmx+zJvO2nehLIlS514vROQDBP5Wdbu4W
WRxdgsI3aJOyPIUlylWv4/4vIP0s/frlsM6iNYKXUylPZXaYTK9VWai3RXT9TPvu
Di2ASH1wIr56w+xlROsUYs7DfjNrMlQwu2Sa2GJwfme7GMK2T/tBNBPCsoGfFI8L
V5lUl9BHIYhv/FqcC22sVN9kah5EDAQwqmufr+SPJV8Ul2dzq5rzN4llemo3cuGl
+g8WoISnxaMiUABeUDQGX1NBGb1pwU1piscdj57Ik/eRVGRaYUtUqLSsley1qjOd
ifRjv4d6QTqSvPnRDblhBiex3XuprT1VOmKSiupuN57FwauU7kzihqwNz7zYQ3AY
cXWpp0e8krxUIpmEaXlJP8K71Cf15tz8+HH1Nv/Y5rrEl4OCn8PDE4oQUc8gkByZ
2HNBYlV/87vP0y1bLsncaWiXc5zjwK6YTjHmJnBNnB2MMGQSIZIOGfG4vdDcBDgg
ILd3S00wm91HRZGEauev373pjU2vO4pGmkqsCWws4JNLwpyyK2Pm5Dek71cSD+e8
ZS9RRsiSX6WpRmGZ7Hi01n4BeiLaDAQM2JUUd9a+nCIX/ZFKO24rGOrSCbJutSX4
/A/ylZDB2NOB+vVSDxhMq3eq01aM5C2wHOw1g/iHZ8tk21oLuqUfJ3EVJo/QY1nq
aRkvWkdoEuVHoas6zVqGeozC6Ak0vvwWbU/T8yLIDkLSNrxh4Evo/4cypxb6YMDR
+DN/2AlYG1beM+qhlgefhD8h5LiOoGodWj0+TOEBSsEqeiI6pSG3jfs7tfVXWkgM
YzfSg2OFvBHw4MjTGRHgLuk5y21St1A/fsWIwJ9+2nxa0e884edUpTg2JSnCwsIN
AqSPp5RxzWM7csFQ4g3FsZhwrs5jfcjdr6a6WC4+HmwezucOgG9BsSROq9FjDKUM
p6+iQfFMZX67etJm8EZRhWAt1q7bK1/FzD2DC47UZFcSB1Q1DGIaOBprh4KATwnk
VepUV99MtKlkYgN62y3pefnoPZIvExpgJfe+gccJhLtw2FTvbNPMPXDisH/L1u2O
oy+2U+ItEIiIImz0j67zeIgW7UNvg6JBTd7XxBMwriRrNBTeTLbFCHUkV3UyyP17
CHig6cEfk3OXqQFTZG5LfE9HwepPS5uhxgZhLyEu6Ik0dEuPehXDTp0Mek2HJyFv
MRWTFR6gxZINRin7Bojq2nZDBuNJVTdEW6r/LkK9cyXX1TnzQXa47Tk/CJlf52l0
hUcqIgBlrx2zNd9KfwUCKmbYPdaErXaqpyiSlfltbP27DgdFvMTeOSeoYVwJJVpy
gkyqHXA7nJ83Rt9idfjuTfMucPqXz8AOy9axS54dPTpvqb5cX/2stXz2nvTXnGKP
9SFHtg3jd+s30G3VazqbzBnGacuuDZ793rJq4YC0fHUO7H32DTub9WplQlNqIzV4
hCxWEV4EEnkZ9nTSdt98Z8lEh4YTROzXWZh13qcDs+YD1u8ZIyY3RmPG5BLiTEO/
4XliiY4+8CjheKz/+x0u4GXnTF85wcFakdlEaGPFVUSXh440IqWoqLkXsc8/2/Oj
W3NIDejfV0SyR58v7jZpjbizdfbcvjF5kVxqMN4DVbev272juzyACDa7NXfxnEu8
5QFlYd43BTdUohe6+dYyaci4+b711UspmGnIrw9iA0SF3mVHF3J+Bn7QDtaRJqdm
yj6+/bZGtmbk49KJm5NiJziufcNBS1b5OYRtGOvWEsLGpWPxPhPn3OeT7MZ+UJWP
2KQhoCWSAKnrClGj0OkfVa4mjzj8myARFysFUtGGpTqS1I9uyW7f67zdMm16+RgI
fKrs73mtz5YPPd+fQ2kzJfuJd9Itz7UVy5JTmNQBnLOP6h4/P/Lw07IbF7ZcjCx2
RQrpAC35Hk/QfT+jrEzVXsflJAkzfl38rsOll3anzEm2XuS00T3QOpgUubi3Yyzz
JCr0TvFD7Ml2VOY3N6IYK0J8NRhPvRMlxzFFaJotpXxKfQxPgnw9kuDxGWeWNXYZ
1RbHGpTH7NJPUu4dBhYKKHhes/+F2x/RjQafkCaWttvWbRaJim2Lk6ZCJErlRaSc
Wf4J0nx98coOVAY3lXY2Y2aHqYFcZhJrgpl7pK+GsJxS8KhBhU34EPLWoljPjLUK
oI44O1uUVYesEhPS9l/5f+yEZcY/YgT8MQ1MpPgWIgt33a8WTbipqeVp+7WN/yXQ
9H5weoBoRepvCrHK1Qqnh1Xm0yuPtJOTX2stl7N/nl5tBoHmmXi6M7sXxJvdLvEm
cIRr4ZgyCaiwJnyL5X5q2sBUs3fCkAJ/6bZ7FkzfW3LW8+MEa18kQuxoh1FFxPeO
v8CqM+YQn7kizkGd0cUzgoO4QBOTt4bvR2PRQnhrBnAsYNf1e57+hpyiXKGwUC8r
BlBgp8Wb6iR9FqDL4uSL9L5H2snkQ8WyBWLCYMZG0LdanT8N1OthbkyHRJ7nwl3c
iHZRWjNjU9HS20WjRIsZuGTHzFeKCURjI9AC3NsLlY8VAvE/6I5sDBG5TJl0VUmr
nDH8UdVzMHqnO3kcHxpqTz//XS/+E25noUUydehzt/Y7n09bBlCDK7jWmiMeexL2
dSA8m84P6u2DddJ8TTBwZQ==
`protect end_protected