`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aMReDmrPskJscpWYThVKVItA5gecPPZO1R595p0GoIq1TSTG+UxXhmmUXc+VYHJ3
u/C3EW5qePLufxmXxmhmDnr9U8/cYC1zLfk44v/2OPb1TBrTsludEDQZdGNWeV9l
cPUMSIfZ0dHXN7L1M1E2XtgoTWQxf3VDHs7B7lU2y9Rdm/ibz0fWMow7op2nWdD8
gJ4QlNl3f9Oiotp1p8vz9RFzzZOF5gBBslZxcTF5+z4qO2W7+xLByngthWm+exIr
3Pzy8qyUo/m2DDwOz3VJSvSNm7RUq+0/yJNOOz3jr3j7ZyCj5OqT/jDAWjJSMH+i
2402Un+wDMOQxi21JLo3cA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="5R6K2aWI3OdbT2A+sz4o9+2XAInTqB1/cSw5W16RnA4="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
Gm/2BIZF5/H5qen8uQizPH9RftTuEE9mgEOF0SqeOKegtP64CfvEUnIxj/ahmIpA
6xUR2v2l7E5duaLZh39Mc1GYsfqE91NCPU5whLaBPg0UuX4cgTkO4cYbW/7yvcrd
4wavUfwXEp2VSiN7EVxL8RcZTSMSI0Jr/aojiilFqVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="TEmQtJ1Dsm7TOzpJk/CeTSSFx/zKExk04H6I8sT4Meg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1648 )
`protect data_block
nvPqn26PC4XWLLQG0Fq8XsMTlhB4evbpiwGjZroFFLgtNlE6bBjdtwWsB89WW4j7
jNfYbKN4sBv0hDeMH0AAR+8g+TCqoX7yLdIUd7aGwBUZJr6FdDs2wTUxRkXFYNTL
pZPBKDWpw8SI9CeQ0UEeIZy8ZOmNC1ZjeItQUJgvFgvn8ALy0rAs5h4wvAhCtM0r
VMdKUCAY6J95ZSKd2ZEUMSElAqHV6k9wd/o0ZqRfh7gNUOp0HbHAyowyibEV8d3h
f95ddSQTKYTOQdPlg2N7ktMmyT5uVyjzDrA9qDRP5nxQdVyfc6hPBh3RvNyRjnFH
+xbQVTlXn4CqpNMH7DpnrEvFMp+E8IJMrzWOff1IAHjymoPstUaaBY/d8QbjbGEl
HgCsYc0zW7cjLprkWS5Oq/M/AW16IlPgt1sODPCT+SDaAZOt1Kk+9mkrHux0RLRW
klj5nzbhYU7rrXRN+S6ducAtQuKjO4RdFuN7FQMDCOFz8fWsRJUQklBvShXrlu07
hs5o8YE7hpjf88rpXL4ouweal3Z8v6YEQSYvUM4/PNlb4YypQkegQj9rBVZProPG
OroAJKdaJ/QmRd+0ZZ+i+CtCfQ52//AOguvKASf6znnh/0gpxjRPVaMgmaufEDXV
N89BJM7q91veDiTF9edzgqRJNSKcTGfTX212sXSxK0Rl5gwd39BRMgMQjTnsH1vh
gAxzKANfNrC96ZX9EYzvVX+I9KM9syD3YDF3wBl9GS1OGpbSfajTq7yMF0XyukrR
NrvGu4C9UqaxI8OGcC47IUsylfykogNnCFO2mar6fgln77uZfZw7DcAnHSPBwV8F
dJQ8GGQH5HnoHGudoiulfidP+ivH/dXVRBgdYQTLIECwJmoula8q+sGNlaqAoQo2
qyO0qIsHweoTpLN5VWSxsoS/3H/+YkrmGpESbjGE9GKxfFfsjfi/kn3WQh1sS+oS
onr0xRYMlr2uqzyk/BuCYDK7n3NdLVBVsPwRSzRvBq+885NyNmkLjGfSrJbwjbO0
gbOI9RsAQZO+obPxuF7+3tBW54t399IDsX/sVpHtIplnBjZdSElfBHh8VBf+4kM3
AOrQsKAgZcQz/z5GZ888cVpMoHartygaazdlwHWhiFXuUdC41ywgMjzFdLOkitqa
vxenB2ko2OjDwa6b2XPNZ8Xzx2wsEPRSw5ZAHKjCuCIsPtGBN+iEie8YtYUKZwtq
vL3JMPSr8Q/lc4YmErNlklRal1gLMdtX2OE1d37ejYez4Y6xAJV+ZsZygW8eBR9E
A4X2lq6nI2hMqE9+6ymIpMQF6NAMb+pLhbrBYNdoq1rbc5p7uxfUizGP1zwdZLGg
kdrkC+vJRFwY52vIl/K/x5JCVjYK2wpZpB5gdQSV5H4+1oda78fNwC7gckTZeweM
gUB0dHuGbFc3/+F8mk0J89rp+9j3RAx7e87Mki8o8J5quLIxYsiPmoPb2qqBFV62
TNNPZnXr7hVGjY/5zHak2+X2FAZrwU987JXzn3ZJSK2eeFC0y6gcXNsih3NtTUnV
pMjXpuVKONw3LoYuM15qg9tl2oZ8R6gueXxFlj7DWDfL8q4lDZJflWSlJSNp9My3
dp2bn6yW9rndCUvI6ZluWvC26aWImzFKDd/DqzpjFhMW/lhVYadjLCCiNYe+vRYG
vZzcSJ6/TXWhzeKLvOjpTiP2RCJXIZ6E1fyd5H7jtmFSh8T+i8gkqrCFch2Nc/ok
vVcrt7eD3cHRN+Jm8cPTRbiVd8GElnQiMvGvrZkzxjvyXk/3d4j3WPppQ4bYywft
8/j3o70YjcktcxKclZy0zk14wSFGJiTsEL2iItHufsCasLGyAu9goFRE1apJfBBG
fxJDQlXCsZwMRtWXnZg5z1JuOvEa1lfjWZKvEe8RZAqmXpx4ty+/cB4JoDR3/r/i
qTKRoUjFgecLpUlR4UVkUO5x47FqAmXM04D+hFNi6k5Eg0wzfBNgeDj7El/17dmS
7kR41JNA5BGX0365WNpjiAEfsf4FUdzOYONXjyqO5qGhI9APjC8eSFD4KDnZFHIZ
6ZkjsjsAMdH8/vsuzfnEkVJKWI1ahjcTjBfoyU0XXbTeP13eBOWx4KY/kOAqSRWf
mIXO4OglcuUAe6LqDp/A99jR5vXHBlvUmOyv0/+grOQnH3wObK3v4KBzwGJlLNVx
/IHjkIuZCO1b1sBDwKgESw==
`protect end_protected