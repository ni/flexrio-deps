`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
j9eMmSPGcKCWAR9PvkqZ1R001FU8QKTyJzFqNLn+qur6INyYDE1AI8LWcxAzfnTc
IpZG7ua3uuk5/kQKKQx8ZIPLfmv6H3t3eWjki8YIAtY/d5E7Gq8Z5mNxMYRzGGTg
TCMm6oOrOTVYlCXHE0X9AW696Z7UGfWirVibl8hs19hrFdeZKGiGht4r09vHR+Gl
FQQmSObM5aSK5wu5KOrK5ZUKGHyBhjnIQO5NnittDjOwxV/57nHVg0pdG6JUqyvm
tEgmCY36RCMRGWN7sekPtNHjqpZkmYrVX1T9QF3h73+8ZekZYd2xY2hpHHGYYeWA
t3+Fmb/6NUmoP8+Pt2hI6g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="wX+NBVcG/A5ruHK3pkDqG8ZVPdOz9TJPJ5saXZYSeQ4="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
j/hqWUoxjK88VtH4QmjIrexFOSwtsLKOZ/LCP4cmrqgzmR/e71apdtoL+o8nlfy6
eZxDZMmrZmJGoazz2oK6kz7xJU85UCwNc4cxAsVxNdCP19vZxph/nCYZQ9lUFkLH
uLBkOeFP15CD3jG5/dp945fHP13J9SzB/L9PWvDC/gY=
`protect rights_digest_method = "sha256"
`protect end_toolblock="sqDZkaglKf+bDjC7VKm3lOELrT2Jlynh4UhPg2J0Q70="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 50560 )
`protect data_block
f9kZDbPp4NLiAOFOgATj9W35i3s4a7wbt9jeHjHVcJxMoXY8rb8laqS5bNUhXGW/
MOc7UNc1VwolqhkS7G27SLamkGClZZtXSbRcN1N+5kZpEaBEj1343vVznnU2Dre/
9Q117ZaagFa1275muC7rLv9LO2eJQS/tYVH5ZM1qe0iqBvNS/EOY9ZvQHwcK1fBL
jG3wDEaZ1hP4sR7Z1T9D7mvFocqya8kOqJaY0KldveQYtgrO+7dx/z3f3OwuVuEm
/mAxHxqbFP84Vhf2z3g59wEH5jBvY0jfZ+HeXrHkhSHiJ7JUxWYYnr3e6IILav+w
LfMPPUZ/Lm0lJdV29kuVUSic8a97l/PYVk5Yn2QvBGdSo5Y+peGfRSGDqvVRY32i
OGwxBhySNPenJN85s8ljE7nDVlkxYmhqects/5+bxW8Wa6g1qOErh2mVyq9BgA2q
EqUjsjRrdva/DD4Fr0W7mJEMV6eP+eLY8MTv4YcfXnGaOnYiL9exFucV+0I7psFd
XV5oAd9lZ1Zq1sQrCw8g1mPnfQBaRZmiVmzASv7hkinArX10IEOsOblqiyaAnknZ
xMFXn0p0o1aDzKpfyJ5nUrXrQtV7eENK0SZ81z0Ma5I4cpAG6HsbPPSU4nplhjQH
DttVjozcZ8IgG2EgOEmFvqSVHZrJ3BUdU1hh2Ks0Y2SxiNuc1KT1ArJXZQgpStcO
IcI1CLc0d3AgaNnxGZ8tJgjX2f8rarczyb6GFdst7ZmnxqpRiE15ZS9J3Es6hD0N
w5bMqik+t38hH/OvpWqs3OSx0/0VNQItCH94UxkV7Ty+Q3SkzW5Q8iBy0SAoIWbO
2/4/hFrWDSwk5JCgBg3e7ugfmgOBUDgpkFgXR5M3nf+1y+pbxLQNobHqHoN3C5IK
BoLPWRqsVPrdwEb337rntDJt8H8hrirzfYaluoPK3qTKm4FgwQIlC/7ufnHTShN4
h04m00JabLsbhzS7PQHffOonS5rUHLACSC7rDROBe8iA7GZg2SkM1e8zggcJB8GM
HveimABJ2XlHWoG5TOtu6zOxTc4SJ/qoW09jBNUfxEUmpcKtfgDaPXw07TcFJxzM
KaDTHKlUsFH3SLQBK9wuTXT+nn/HyDcFt21FfvP80rUzdzhkbZTBYRBYE7luzA/g
bgmOR118SDhyoEHlfrKL/mGYAK0FnGSTvQnbTqGNtBL2i4EuK58DSRFyfO5jxqNa
QWFA2So7yOlDp6BySRCirDCxMhBLjBn+SNv+JBCrsH2SHoVxzheBhPQWb4s6q9zW
WeyumOkGx3qYOGZ3dTWKJrOnBIrX7rcVoEG3sao/j2vzgOnVjpD0QWp2sHfcbjBj
yWutWxxxEfrXxeWjDLE7bMR4YkXng4fzXLLVKzPTs3u3jxTHUsoM+FIjHTyqKfTV
z5dYrmkkL9qYgDqosGj36PVZf2UeJDL97ugV9XEnT1kO/DDvBwRIR01mnaPoPdtG
O+IzRwAq7IFGl/K3AqVrMEPtLAypsh7T4XohdI1rrF5OCcBBO1X4Yi6NP6mw/Dff
VdEwk+Ke48yTFbEbVuZMTwOHgYeSu1tp3gZ20eWpmjjQ7s2//gsIlCokMRVxBYYk
x1qLttnoWlskbym8ShFBK7xOyVxE4yvVtG5qtam1JlqT/BSw625bpspIgesKNWNl
m2dZ7J7xA1l3GRuh9fchujBKBsqToTSW16T4FUM2FaqFBQ/bSCnsB8sHNzm0ArSI
KB6FdUIcCQMe0fy6hajT+yrckX1tBKhUZgAhaHLo5dS9WYgGaaq169FxNKi0iPD1
/2WKNd4WcCfUmSkOoN2w+T9QTnn4o33VLYhzl3YDlBWPLTKAa0OMrjlt3cQTLf7i
ukigDB4EaBw54Xur+uA0iHJHdNH/cTYsZxBB68No976smmA7F1y6QLlhyoKMUwNI
4IPEQSK+hq5AqGODcgIhO1nuDPSAMoZojrpp3v0tRS3uwS4s/MGWHzvCHaeKD4se
2dN60uJvF7KGQyOJ2yKuY8x5NQpjSS+s375utj/lUC5ipOqx5QVwYRWXJ8B4Knv5
EGEXbYb/f4HHUXYzf4siwZPs1krbeuF+tlx6/JWQT+a56Z95DXMC2jooaJRGKS+U
C6X2v85n5fERxC14ywAGt/NLk4A3pD0ZTrBxbxer6YZ9wDX4YnwILCqNLe4EZqDw
BzV2PaFpj2hjTM46APVrhcawpciXNjSecxVLzSabGcHV4BG029kAa9H1y2aL4sej
IaHmrOhpzNpshgTeR9CmmOhbB0LjGA/P9c+W4RidIQESlmvR0yZTYWvYdf0HJF3t
utawaVU5KkIAzocHwsDbTwwNENVJZlmjiseZwzczZ1zX+6h/p+XfYDJK75yoPKBa
TwK2j6FksOaevHXHUOrx9MTFBGvrhmiqnG0dWpLqGZagxwlR7VNuPPTHZWspMjpT
NubhGl2JYX/nZMjiqXXOq9asezpOGGwAqcHUcO6pKeZ4XlDEc4UO/QNTBrHsy2GQ
eeqEv0R+f1kpBhIojZJfo0FzCBn2TYADrcxIonUFH2lq5qBlytxmjk/9azznglXs
5yGbO41kzAMctY9WDsxYzjvEbUn2FKGYeQ67FlvBifL8NXJZnEGoD3UQeXxz4HmX
FD0JTUtqakus2+xglo5MF1Ymz97Il9dDHLfFJm8HvN7zaSDJVaZDKfAhpOUxpzq+
j0oAqqkyuLvT+LkZrEDcnR+vyKAZfhc8SRMjYpl+XFQahYrDpFapDIxMfFY+XYsU
xiiTDR91Ve+y/SVz0tHVhJY4pPfgz/ceGK1wNsKvNeTdd8Y1QrkLQQRRqSTJ7PTs
S4G+syhd3uXp8sEjKJe0G5SFYKbgWP+5F7ieV/KpX+YvG4/eZPNn09h9xdRaQgVh
TCIQ9MClCXSpJ4dBO/AKgY6Y9yoUzvV+6bwer02PoKfB5tv4G04eRs/yNWd9OIji
HsotBbUdtb42t6p9oe59KohrC/pN9Ah+dmsvuFCQqRvxsBUttJTKJcc/Bkm5RnR5
QXP1vgNJPjwQfxa5LUBPtQQnWtPgcCNmH4/AkzlNKIp0qPcJp6XsBglSahsj7tX3
VgWPIO0/Arpvnmi+ATfES1de/r2xDc7yvVuZB69sXrwhc/8Mj3d/DGlIfkeX2d9S
2S+BEwr1IKRvVDsQVvDiVXiHEVQJ0ooOZZ74XEwwjRdQoDrIJOPlbBnweFncIDFs
EzULai7kVSCGOnApY9FpXthTPVP+KliDRhIIW5hYaqzypuAG7KwUwGirv9kssSUX
b3AjUI8qPw5iuzfn1QyQ899GHWHPjBMkyfB3yi6+dIufbn/90mpZH1QbUngWIvVS
nxsdrScDmR1+0sZevXAwyZxyye/lKrfRZYQ//Dz38SgyUnbcyh+3vaEkLsOb5FHL
MZhUTVtDi96UnAYiJQ23KYKcBCuwBLJCjMZ2RCOI9RT3nEBjD59kpBlSKNn87FFg
VxsBewagQO1/KcFbK31DWNyxS0AxWO+Wl0OwJ44TU4KT4ZnDk7TGvpL9yrW0RcjP
FunzmEKAcXwnMfLl1bEtXhSCfwqCJS6sjJxRdROe5zXkQQ4G1mQwAa1aoV81cDwc
gSXNTavKx85vTf38PxqRpVsXD7b0epqIqfF7CZsF11J4fMd1X/NbwpiDnuabsCcG
B102NAvQwq/iFkuIuLTu86222CHJ07hi8Fg1KTSgChzCtPNxKYjSU7qoo3tsxUTv
5vzsUZFgol9DpJSLblbwd1EJc5kxXru4mXwZTiYhH4DkM8qsNQ8wenYcqlbVqa6+
n1Cbe3Uj0V3IUku78jVPreQ5DdD8fbSqQ0cQI4ADws0q7hjI/sGVhmfPZz0qjrS4
zZhIHLV6dazUgiUxu8rObDCqgM87cipz92X4Shz5jbuwOh9ktwYdXpYe2gJe3fly
I1gRhAPjtJZ35p0xBzhQNiReFeBrLqRZ5jOsX9Hf3aUrWHoyqmYtR0ph7XM8ngLf
jHV0szRB3ooB8Rs6nbk+pB2DWhjFdLZUBZUspWxlqdU6OFLc7A69MoLbzb0nOGWv
YMjzlFV1/ViAWy0sVytyxbPfl2POml1ySQGDNblEFk1EdaqdtMJKMzJHz35DBg9A
Ela187rSbNiyDwMmDmuOpehdXyDvaet+oKwcyC+y49WGw/3UmZlkQRwKwxub+q4w
C06tyd5MNsDJpJz3OiH9dpKhQcgvA42ZPzFJIwDvEMAgZsMIOeleUYSinxitAy6b
clbeJPwGqrs54atR0n+T9ia9RMUS97830sNzIvyy2NstTjDXvtXSnr0yyQOAOT0m
WjO6EHBP3me4oupGx6MqKtAcFyyHsSJITi0FvFs9m+PoHqsAYWpFWoY8Pv1R65XC
FkGIB7Z5PBw65Zu1Wt+PYJG/2Yf0btbZYqq3FI4xHnzlfp5wQvDo4/SkkcibXSwd
8u0lSPr2Nwg/veBW61TyK1Gw8NkHQvLwLaa2xDtCh2uMa2el41z1EC5R0H9u0ouU
6moCGiJG/gStUZinFrXPB511TA6LcJAvQ/5xYztpsRMFtwX46jcBv/+5O4LQ4B/r
jxL5xx9gsioFuagEJdZxQlp4HgHqC7fodOEveIOvRUkPD7onWJQQ4zcfHHinrTZ8
rj+WtK2yN0u/VdOmDLefvChyTdG3bpc1igjy/BLGGlshFVp49lhalxsFkyxiPMBB
c7kyLl1qaSYhxzTMGZOzODuAxRkDJrBC38h5BSsHEFv2XnuaP9auVmsG9aUb03Mf
BVIg+Ztf7rLLJQZonx7iJ+X8GeFRzPNWB6wJobcNk4JJ0qzK+D691wFmpWgOoMP8
viCr30QIQipzr641CFT39MX7aAS+5yP80+YrSVmF/oGs+KefjM5JYCfyKR3UvA3k
Oj4hflskIkXBoTYJCWYkf/7pp7lEa+qqlkU3sTQEQbpqKsRS9cvX3zHHxG6sUav5
hNI4r2ZpJ7zXzOKfMcHKnai+HlM/zVi0Ba2JuT3mC1mhtp+cgmPgtGXpTbN6xtvi
r7BuuE6/qYWXbXzcLAsW+hcHGnVYgfgzNQpGy2oRQYRokEjFKIq4UEaZ9li374jj
Dtwbw5H8+FMHBcNqkFRMFvXPo9WVAcXsP/ffgFbwpC4I4v5SyoRM2u/Z1Md/AsCn
J8tHoywvbDb9sawNQDtON2PDL/Q1xvcmRidnN1C3kBjF+2CuUPh06pXqvepGxR8d
6CUcBUTbcSadCkEaiw/JB0LoFW7a4AahIAv2f+q14+ZmjUg0ihb0S9RYozbdZaMR
/sxRwzBrz81bMbf44BSYkkjmMj+YF/tvsfS0AkIMqqv4nE3PWXn4/ErbWx4ar8VL
QPP4/3D52SXHf3NdBc8oct5zRr3JWw8QuV7s9v9VKNqmMVBnNmAcyvyp2SWK7ab+
by0woQjSjPT9L5gpTa7KFbG591pRdD9/12SFCq9YiZKg2iESX0ExHH6zbTJuYJ81
n/aDCAfRSY0FCize5+k2E/JzOTghIjJLi0AiFtGAHPnhJ3b81wRE8P6MvLLGxhlF
WLjWHzVzrmDxCQhHekUR8Dn80n/55wJ5F9wUfMJ/EaoYo3p3AbDcjQ/X4tX9cYON
avRDJmZNzOnp3tTLIXSVsLVkUry0P3KGqT213XVN09J+wXwZvlmW5s89jqbdPfT6
YvQK4EWfZM0QOuE4Q5m57SPoiKWse7A0Qogc2wmn1Y1bHyZJyelSzcm22FG767HH
bpG/2dnuhwNetlHMixtvSJ6qStiPl0OqAr8vF0dtFX/5yh/WMZuIuDh9LBha7Nph
M0BAa8LdVioIoGQ7Mk5njM4tkmJeKjpGULbgT8pTwuTn8YC94lBsZeDihC7k6der
VMJqJh2WBwV7feU7y67JcvaxvnPyHTZ5KYL1kQ/q05L4VVEd6Gy52vu3I3bnQTxq
/ynkCQXmXkMcJDj29U61vOkHeJYq/94wRTVrvrgO6jbQebu+nO9iNRtO0WmSHo/I
y+3HjxioWOzMh86znZ7+MB7nbDQUkrAD/tyG68GPedSWAPdiJ4HOHyurtkCDrOtM
PFu7bb7P4JrksebupTABOkNGidAU8VcEFi7JFlk46TPYzQRHR170JEEiw8RrR6L/
XVEXv6DnUR2OCIUAS8/9uOxDzaqYidkq/OmFgo+/weKfo5IxlN6jdzk+RvFeRUkw
LQEOFMlSEjhWOU2h7SqmPA+6a953UKJ0syOqes76L/qj7miMwBAlnhb2xcr9OEo0
fXt50zDTCS4KRy2Hp10ztoEdfoCtmVeMjcPOJ1/4mnB19meFNKB9hi+0YrnQO4xl
K90BMtF6uq/BJnXk2kj7CUlX8S9UXBiAChKYLSGMg4u0Jl2adpeZT/6pzlfW9M1a
z9Wtylc94XDbgq5l058+fUQtPR3mnv2CZtOb9jcIKgK4GQxQyloBNT8MnfrOyzW1
kAic7uPOelKV0m+MDUOsClbYxZg1Fdl7zwSjV/d0MKqhbTqhJJ5KZDIJDk5otKay
/wDYm7oNwItYK4eOcxt+nlrZhnVrS2+6fOX5SUQUYjQ07yZoNy8i9n3wvb1jt04I
Rj1g6cXr5v4qRTr8G7930xtLieLvRIRlqumHEaGsML7On2pGxDV02fr91D0qA+t9
qiRZNVZ1/ALMUVbHVzrsc1epRYdZEO2CzARLi0/T0+s763KMCxCxekY5arW4dH8X
BlBso9x4FwUxUDrJfASpWBTjIKs+MdBlvqlLbk1xusZ9hcEHSLUC3G1prDfujOnr
18MSvY3skxJ/pddCnEuQ8FqTTvgyBjNdtkIEU5cXnx8Yp9xtPrtmIeRrlTK8LwDm
alJ1OGJEoRBlw/uAOvIicw8utn4/g5dHHQdvb91BzhOeRsPByfgUmnJXmVuCn7W5
64V+Vk/Kk5tW/wQyMjr225Re5y9Mwyr8KEQPPA9Edt/6+hv+6j9cGUBjifTAtrB8
7nQQK5zSHuBwXyRyNzrlefb/x7cZDxLOe2fhSVr4mO7PwLuWEt54lpFrr6sy/odl
v2IU4scopUXSohZBizK2fmcSg2DsfOu98Ee6gUN3uLCWhvSXKvBbLD1WWabuFzpL
asjXIcJrPD0VnpEYqhcHkYwVZFCTNhuO8msqEMiNW1BBcZiJF6o8vNqSugQRrHj1
JZAi33HufTb8PXBdW5iIAx3AuhEGmQsa4oASjfHI9bWMfPjbCZFF8IAGfRYkEFbT
wRKjeDEietTRq0KKqpBQC9QMWsFE2RhyQWt4pCntN7kF6jDLSHE2L8qGZgAbPnrT
zXjyBeNfhV/et6pf8UDgJkRHScMJi1pqX3d+vFhO6yqHLRxpMQd1HX8wjinmptVc
zfe/d7kvyjuoI152tdTx3EmueJcvFRsoXuhLZWjFMBVWmO1HaSTJclQptXocT5UR
wxuZjHV9YSTUjCiKSWlp7vrZ9pKkCCxzpylcjjpSvgDeOcnx2WLxaAqN1qD2MLqy
mGEZXTCF5aqONDv12ogVnWruuNfch+lCGdvUpr1MyTSKnPv4j6QdvBcVy4RA9llO
UCotVBY4DGioIUGD2i5oV8Te6IG6Bou4C8n7vADm9pPZ0wQnCaLFgjBH+8iIeq/r
jANI+YQ0Y69XXa+GHUB4H4PqvfV+7QOrScGJzI1NK+DRB1B2eyU9LQrr4xS2FSZz
awNff9a1B99gvw/QAcPRgGLfcaAI/ZxmfS6j+Esiy7+BUXP6tr3su1ng5LJ4j0pZ
t0IubK+/+axmcEPInIzKzqXJLGeB4D8/ITNJq62PIUnzEyF39KvA7PH+cDA7LBFw
YyI0bG4qPh5caake1t/iQS3r6/QTD/0Ny2MNEkztH/N23KB05bm/wGFtd68xNZ2Y
ijimLFoI9wHRnmMQjII+pagg+3QF504OWVA7eXggY2oZljzfiGexAFtA29utjEWC
Gj1IMTln6aaJN6zkT4I0kFJO12Q98iOeWrrnoHvCOl7ttgTpebZeKCGWVCRFGA5h
gajbz6fXa/2SVd5YX9lEGFRrHjAK9P5VOSsvD7G/wptDvAiib0H96RfBfbFTLegp
BwsoTnxwjudYqgWTcy96JwHLSwZybxZcNOWBwlsY+w2HJ7F7X8wHYBlMw0G4Xps4
fBtXbAHJn7JcvSmeaWTlTGb/6xikz2RZ8Mq4WZEjwT31t+DM7q/iYVZKej87xTII
OpDWsdRaTx8hO2lh43cjq2emPj8PBiNVybuKHiJoHjLNxsmnk3dfuERU5MS1IFtU
HitFW74X7mscveWKrHTIDdHtvVP6k/RwyikfKTNO4hqIekdEa3JTxeAD3Olf+0D8
EUXnHcBaPmRt2pv1veyBJAhjM9/nXTRFU+5JpZsi8acZQx8m80gWEL7rmj/FtTZ7
uAJqaHpnxvsVZwN6ELQJ5irsVdkHqcnEeozNfL4NtxNvtpMz6LkVzKBmdvfvLFLp
TSOQGMKs9EQ11AotU4vu1rMi3FE06USimcWEuJnfq+YugMHdNrb+A43LPM2NUfC0
MgomQg5eX+v58qa9v9UEPfiRBVt1aM1zEZJBABWiqjztZ7dAvsoIawn3BBSHzk59
orx0rWxRdrrEwOcUWAQ/3Y4LmBemgCFHUg1+0wIADQGWPB3XmD9+WVd9l7D1/lSI
0ntDQlQP/n51S5Ip6flJpjGsob4mrnJbHu4Ctg9Ivk/1UqDOsnurzW8DlEnt1j8a
sIs0IYPrcFpQ9jMliK5BNOR0HsFDacm0I9lUlSBezRHqZDo2E6ByQkkiZvw6zG9t
KwkfE7c5qYUZWeGlcL9FNfKrfW4AwKZ0gcz/rUBSusBcJZ3J2JIBGLxXyd7IlWd2
s+vI7ikXtLiKhPGO8rbCSuYBQP/3PasHCegOWjtvPKaQ5zpZdqlL3FT5aTT+Qtvt
pXzDBEF9+tuCH3mrDTbIA5PtraNel5ZY+4MbATldhsbVj3ZCdufBZ1+B52y6hyV+
8ffR8ChCZvd2jn0f6QSdgx+5eJ2pDC4HQK0tjxuHxeL32AigMOWLyRFVbPSQaJj0
/aWm9tyKmBaWs5ahgsjLtjSb2vCIismm6A0BEBjHWBHb1rH2NaTw7hXE2dCaDrok
JTb301CIUkH0VfdQHqib5Yl8wQtIXvhll+qudCvFjQRS0tj9Xwsd+Yt6GAnJsoh9
+rQOO2IZEYEeS1jYC+HWo1FIA2s0tHF42OXog3lbYabI9x0Q8HdBTbxzHrU3LJhm
yAWzjucNkuASaK6FKiL6ELfVOSfLeaa5cXwkO03ZA0NpMjfVnsIQOQT07CoUptJv
5y7pCrP7KwmnKDrJq/ITyLRULcOhtmc/z3BymCxZ53psz+DFVRGAOUma9di2mWbh
k/0WaPblVDwOBw6R8D2S45sTYyp8K6ECHJKvIuM7rzQxNtQaqWsrDMFtY1aIXtWT
BItfOaRrOq3qExZPl7Y+8T5UW9Kmk+e4yo1hXLBgK/qSkG/C1FFCtw9yKpG+7oD1
XcfJ3HO/ycuvw69kWqd7/QTeaqe7Xt5Pxvd9LqyI6f7N+u0hmsN3y6M+020/Qxps
m+V7x0Jdo5IrLh21E5m0ThqugyVnQtGkNZSDSevHVKUVXRMsRw6thYJzjjIocLca
RQDmLhDhXQbLuYtVziBYrzMMBGXos1QLylgBGcvcxDNHwY5GR4lCcIRPlFmFRhEr
JiwvnYbeLgs+XZQobtnY1+ecpMiMHlV8mbQghe+9El+uVukFxbZX1+9FG2K0vMNw
UbXLVgLDq6hD1xvxvwzbcQyFXx7bO+8/UPd+8n6yiyIdPpTGQZWEta1kelRsTdfS
yzp0+q7RiIPY5t4Q4MuaNMyuIg8RiR2VTtgmau4iAkbU0QyXG9LbeIispqHh+22X
3BtKQWQpy8F9q/ixBeEmZSfmQAj5aQkGwG3jVypduyMQ7pKYrx/4IRq5fop4rxIW
TBBNlIuKTyJYuifupDKz+IuuXFuOrmgVLxA+00443XklfL5eMJhqSNUMCVuJlz4q
wM8YL03kKE6At4aHKkCjL39PjsLD4Dr53sh0bi3M9vTVov90l5eNp6eo4b8xgGt4
lZx05UcwuqjrPg8a7x+KpIoAzXLU7oj5qiP95Cmp6KcvLvUakwDHeCueso6zSNQo
G17utXkku+OO3d9Zh+aW1jV+M+ON88zC1BiWQjOCPrw2SyF1JR7XTvFmqDjWGqQA
Biie3YEvgV/XpkNpCB4kViFljsyHCqP0sYsh0Guil9feBqVC942DxYzTf/6X3LRB
hFt40K65fG6/MUe/D0qq0owapMdnfnH38tThJOg6rLhqimfb5PLeArQEbDMCU7V+
9G/qHnzigwkTt5vse3G7Lj/Y5iVrFIKmvns7yQCjTym/qx03mU0yPwFE6GvuxP+I
sqKzww45CNDcci7P2XA6XiK0HUHFL8B3uI/R8xPvC0LeIcv2h0w+J3eaDt+XZrD1
gTnmagYtBDb8OlPvCcGTwfX7pjdfLlUq/JscbpuW1Z19AuGaIcAP231kqCzM+zZM
FxaEZ+b38AH0hpcWAr3DCd7csmB4Km7shePUmOBrGkhDawYpRHG4HE2Wua7OX2ll
/tEBpmljkejvafa/gjo8nW/RyXSaeceZ7uIFeNSwIEFQ/LqE+6YF7vDYaGhNGEci
J9QVXvm1WUqr0H98yaJPdkzX6VbI5DaKbZM4/eIxmQgNaZQxKujsHMYx09hviKPW
Jz0PdY17rQtIN/igemqIcbL2nHwqf+KrQjVMEHDppurioxluAmE33TqYCpr6qK4l
OsNXGxdluvWtX9aaqgkFFJ95bIq00qKKHiSfqwx7jPn73+SZJRpMR0iMCqczAlwd
hFskJs2uUBHInDtzxhef3JFiDR8a6L+Nr3USFVpoTix0hZwGwII4H6kHnpwvNquf
5wp+zj07uzJYs2SdqqDEKDkmBeWp4sXt3DWsnjCqOvTZYMA5tHaft90I0AtlsJdv
dOgGQuNBmDMTMUJiI5Blm0UJM3f7bCJLQXekxX02qq6yaKjQMJ9F3W/SvdhA6K9G
uBMCuE6h4WeQBdwkJq1yXweWAljERjGZ08PNbzYRdpcickVWFwk9DA0s1gxIhd9K
4Hjdn+zNO3ZcNslUxXGnqaBPYzEkswJ39ubRgmzwGzp4KRwynYKQsfAcc4gX3/OI
bP5GhqQZ4cEBJ9me+jjCPqpR3oUKnzNTNgxeonxSMXO0UmCm7BRICy/xSRUgQfcf
oSZm0aPnEz7X7QYS/IpZCKEWjdVIOX+KQRyvbCWqGyysoremYBbjTRb72JxlIoA3
ZOCp/UX/+UlTQ0CSv3tqRe21hp1hxM02AhenTEhYUX0Ij/ckQAI6Euotuzzg6cJ3
i1TPdfIwfvwWJhsGnVCDFieoxT020esAWYHtchMabiLTMUpaIM2lWFFGVBUIQM7m
L9rHtgYWyYiqSWEgyUfGy++MjfgqS/hIQkt1inQ7fy6P74soaX0/kE+m1R1aEWQ+
/V9vL+6pLXETYwuhkhd1uMU7MPCPaKeXUyX936P8A5m6KAR4t3/AhRJGxx4BG0Yu
TDrWjHo+mPgDa3vMDICIX5iuAm0HVC13vHgekLG39/T6Efbq+sjM8RWONSE1Z8OW
t0QwSxbi+zNuN5SQiFM/6D/YciSOOD7I9W3qRq/ebjv93Cs5AiY6ryeMLNbBDUwM
NzmHgL9AHH+9GkpXd1VQRydmskJyblp8fw3m+oQvIolw9w195SMYWDvKKd/J5SDg
rcAaRTVU0VlCNqqL18Y2RPDSvVQoejrrrO/qICkUDPNhRk4xgv5vBIyXsr83vo8x
jDZ8zOb1dgIlVUZLMP28r/pTpPI3uRJQ0GaUoBwigbUiAmsjNKHYgVaZVgTbzdZ+
x318KVC46ITv5+TeaanLhXqMPaJmuZSsPJnvuFFxYGdFvJN8yrV/bmL/j/rCF4uq
meJFdMV5xiwvxjHwcToZRpeB78Se3qy+ImGnveNfGdwFSTpsToVzcmZXGMrJbHAU
u90onGgjZyhqdbfcoc/1LF5hhnTju4AfS0FPD5gfCcXvVCx9Edt9PlUZw9sBlTCF
r3EwkqpzFZPA7x2UMZCSfCPsTjpAWXT2yO4zKLK4nRtFpqBllRDL2Dqz6lNpzV8t
UWSSI1SMqw7Hwpiilj/jxuLS6mAGpVdD+HArd4nHr3Rea+Ye+O5JIwYz7IUiXrZk
UGFMpS/lY2HdFVnZvIrPieqVJI3F/e8MFFxxb04Gmii0v4JhyCBzxVxSWB1UKy8V
c1QrJq5SScirRuLP8ToJ5PyeRlQr7inFqwvvNBTw/Tb/VuK3Qian5as8b0gnBsoN
VWAb+PUO+qcvM2jQWbT4edWJHFZsMUVXeO0N7nDQ20xd1yvQgNP8pJkcFR4/qQ0H
3u9SdS6w0UwkLCngjsmz5P8haO+n9J2xYDDvPaNqob96z27WHUckkWbPIVsNqYQc
qNaYsqwl2DR+uqt5FeQdL45l705ARHzU910gtKKcA2QJKDhZhmzXavCOpC1qgcIA
xrwq3bHlj/zx2JVQvw5Bp+gim74JyR6fbWSxqOI4T8tt4ObrCcWxvYUX/3FlxtFN
/Wb8/YMb10M4gKNMN/ieRarDce05QZm/AZSZ+0uuPwyMU3D7kcqCsyKy8Jem0Nww
jtAkb2VWLihERDqQ/mvsXVjQSPXnHyKsVef4x+7BDt6N6HFvhw+lvO9JnDfgm0D2
hzG7UVTRaZv719bkCi1ZRfoDGJrWLe0MP+QoeCzsmEoxXGar4Fd3KjtgVvt/kbi7
Bw8DTh00/y3TvefUhkg07otPE4TfPALKDji0yAw13HjXi7s4wGJcGI6suyBU8Lop
Sv0BC36tNhiQRk2XEGqq6AW7CERHExH3Xo/OZNKKN7sUymPr8+qsYMDpdQ/jC9n8
NiMXx4UqhfiYNo+09UrkWivtfZGMEgYgkkWrGhoMzNgiMn08MBIWN0EwK0Nq+S1y
7yWR5h/H/SZoX4Cs3YZmsh7L/pwNG0oViPa4gNyMpaRStujpbSVAwHTia8YowU5Y
ECs8FBU1iT0lcLKKLSbOlvEV8UZ/+GPYtr2cF2Joe6uzZgqYH+5/GUaUnVCVNN0y
UasUmxSSL4yNCoJ2zK0MHLm14UN8KfDWOXqbc1kktVytJEJayXTN+SvqW9tc/b6L
FdwQ5tJwZO4pP3qmUp4qe7PRvMtU7Oo6a4TEfZpAosXjaqnPtlOJcEQfbPgcSIQ2
YbcqKteBWFHJOPR+5ttkpcoSk5bPY8UhqIDahfCSYkL2qYX6GzWk6K+rvw1TLlOe
sk62QUqWjqHEjgr65YVWVb1w8OAUD9k/ZC6lMyd6YaQtTZx6d7kC87kqMn/Nswsu
aomzMb+YimiQktNdCyuMmpeKLqdT/rZQBOp0LnmMMKUH3Hgd4bCNl9uOVGs7IA4T
zzLiYgndqfvqHGitzd9sJm5rNOS57q+M/DUDh8mhRx6GQAMw+pikcdpZZechgEbS
vmFQ0d6IPQfDHqDMa2B1jdUlEX38Cr9DrvBa6EtnItCaDhAQQmS8JBCTBCfB3onk
cDjwnctPwRz6kZGJXHvhc+4gN9l79MOK+5yprQgKNwDCvgbD9shlE9ezWidjoAD5
MonuyQonxWfv2zXPbH2MDyrlHX0xdXKd4EUZQxGNmE2Tgabil1cO46d+Nc80yZjr
yAODhQotwubREWX8I9rurceY7VXYf5QZnV82Qq5UvwiAOZ4a2uubjwAy9w2p08Ex
qteVBq3o2tCfRvkcRfH0Szfr5O7fgM2JePejVCSsog++TUpMq+ohqPK9gg4/LsOU
XN89Q61Y70jAgp+uJJez8wGdRoyh3LFn6MMLUkzK0tsGf1RRmiWppC1c4JuLr+4m
2cKfr5ixnTvw2OkwQWDGWD5+CmDCU3kcXwhf09Jw0io25jrcQBfgIxcfHgt+6/b/
bo8/86fsOX5zrE7nHAl1bp9uXvFaL1xfuNV8AhY/4mIspvuya1TuiHxrcCX4iLJ9
/fazkxitEDU5snS1N23/w0IA6fxuhKFungiKIcnSP+CXzaIJ+RKkB3q0sntewMtX
OA8g86NMfaaedrpOUViHSMs4Hs/+O1a4lZuGLbs0bBUAudF+VDDLS3NU1pKW4wku
c4YiXqscT8oU74t+L6epR5ncCNG2QCWzghwsvqkyvC9EU9P1hpTI5DtrVoMvZ56k
KVTDRSZKLaQCgWP1I4yYZyeau5pXoW5ra0nJTqAXCWkhzvD4xighyyCiOezMW4fT
XvNuZOGy98x308pg/128ZoxNe9WkFmgj6sdfTTtMYSMYaAFT505zk6HjLSVG2hPv
9qfA5MVpplnWoXmmgKnc6v9amj0tyIHlOhILE5dtxw/H9BWx4fUJLYYLZir+j1wz
FNPWIgwhYtitMcuDNsjiJKiFkkfwbGHy7efr76rQuw2p3ZEuTknuSHPP+WgElIcu
eanyVP9j/kj7nvVp3q750DC5+RutwyiF4kSC5jMtaCIGsCRfTKfdHK7WnsTHOk6Z
SEBClnDfwAupnYCN0tXFRqD2bqzNlJUfmBx7kfvZNUbr7ELp2PCc0qnAtx8+Pz/E
mF0UTR4old7Jay22hi3GQZscCy3Z+27/3HxeMvGY7t173mvGspazNVckbAn67Fq7
ES2TmhvCjJlGDoN5uXtN5VOEi0OaXFc2sJCPK2qEj1wJgzjAVv7qp8UkfXtUb/QZ
Y6ZRFmWZPO+rLch3dwzteU1emO7Nl1VkG0bROZOOpd1HSugRDnfly6Jo0ehSNrGp
8fK4RvEaBUfOf8u3UGDqE2TktC+FwJff1n5+IHSDrGkJCeQHyGacbqhMoLDo1BTU
a7v8sdtlQKokYAdU57xKmGZaEiMpfNg7DdM8njqWAvSKmGaVWb8228FMwu+E5esR
JQtzkMd4w5tS/DEI5cq8eo5PdpP6WPoEFCKGSFqYxBY+ver+kHPJKCA2tdaZlk+K
34/jPc3r2oymtfaJ7yvrUCyyMQTU4KZJtSgRO7mJfttRP3B8L/I39oss86UpkZyN
KvkVsmo3QF4MNnGqP2sZPPfdxC3JNJukzTDpyv3PyGHxg3Y1PMyF49g8H/CY9IID
do8TWNdWoKwZHkgDtQyxlVZ3UgSIEzMcskT0M90s+v+kxn2QI8nmcYIUsOl9WUCr
RG1K9bPQJLbA9AGJmTDTcI8ly7UC1atj5uctRxdBZu3gb6fl9+/bx++icbEXeNqE
Oogap6IVYBCy/F9Wm1HuEt5QaIwrZqoyzsh2UHtzkKj+6emCy+AsaGMQ6j6B0IzO
NSFPsUPE+AXcFVzRzT1n0DUY4nZ5dx62onqkm/0D0wPsRXBBCeM7wCyOWP0hG39/
k5/s5xGSsPvfPuLZDQ2Ohw6NBwX9pVf3SekojN3dK6lxbYdNLD/syGaeI9Tvm8nQ
aBtORQt6fwIN6I3e5ocwQ4haUtHnzeQiJI1QX0CSTl2mJDEpWUwOisf1jEv77YDk
PHufMsT5dhHXCxG00IZEoz1J2T8rwretx8K6mNMyGGytmAYGT28a9ALItXCvgMIO
7hoAh38n8d7fkib63Hg7VXl6umZnCWCGHz3EzkbDKjfKUUPhWmMDhIk6sdpmhde/
v0S+Cnfnf3EcPoWQ2Vv9rkldEeFxukmnMWKErdRpJTn6TOe4tLtjaLbFd9Eb8qDN
o+xid/FAXk92KTu78Tp41yVCemgn6yMdonF7n+hxm06SaZW2dnrBCiRg74E6AJnd
s5twfPkS7C6se6NCa/hg/WsuEkXZtkfqfyoinjchYoEXpBy9rDNRlSKIvnvzH4IP
GBB5tMJQiJdISV/1snS9d1WyFHEPZJyz1fhvjKjeLxs+uUoeeIBED89Ec6RXkPPh
bM5AO+UNivxDi6hFCHhpydv5TuZ3oFq/tAKDU1A2t38hVDLzFy1GSowr5rmDfAqo
Bz6zMctAchO5tl2+dGk/yByamf4Fh6l+4KwhEkDNjZM831+HYoMUg4ZG0k5xj6x+
QKJHnvN49+Bn5M9T9u0lR82U+y/fZLM/GAk3xfF+Pt0tbwT2M7ZfYC+XlFkOKgZq
JlUztYY7HP1Lj7PLDi/Uc3HPCIHPVua3KMcK5c5vm+SyMRigTcWhdV2UPO3IX2pg
eip/K7XGrB3V6jJKJ6vhQzHbXNCGFJBO+kkMkjaFlcSkLVmyuWeLLgXxiSKqCf9t
OFUrSRPCqab8OfP7CQymsHQwwlATLJBiAhsztUqAqRvigArVlsEq/k9i9vpyGGUi
2lUBWx+a9XWAa9E07sYsdQKVQRrFt51OmekW1gAOUr5RLOCIM5+EPbRHuJ80tmqg
nYBqOqIBvnxJ5KFuRlym1NPK1lBd9/hIx7oEiE9tsNLA49A6jtyjymQZxOiWTXvS
71hRQG07bHS/sDrpSChoXxtNj0SHNbdTcM9mNzVrg3j3fpaYJOtChlFGDvu6AAog
Xv20fJWSa+PSkVW4S5TdMgfwP3XpbevF6/94fgeaB72bHeUL1/P5Eya2azQeBm4r
YNZs2xwT54WOppA02oB+BsifyF9a+FhboIl2WZWTVN5jZlCn1ZLGazky+dAs75HR
1yX5z/D4SvMf/Eyzpqy3OEGYfRfMU8XJyFFfVcTz1XCu9D42x9X23JPI7ealZ7XM
91DlBVFqXxrwOgC1VGX3ZlCdzORN3qjwcqwACXnbQcrbE/w1EJIa9SnBAepGd8Hi
Tm7SR0p0HK0mzt3gdgUh6iwge8QLJfQCr/Q+yR1R4MO1Qc3LZ8mtFSuw5Kuh9DX0
JMPBDU701xNWRAGT61AhCeSiymE5s3burK1I1+HfH9DZWtKUjKquShk9R75QZsUB
SjRHjK6Nt+lCR90Z13eEA++AQUH68ydDmVTJRNyUZugBEEFzzXna97sMSonEXwBb
1p7VZHBHy7DNs2y13apPLH9cxYoDh1PmzYC9OK1/+rjRolc2VmPB2//NsNheY0gd
LZb6CtZZlbbubhuJP5evCi4K/GpZwMpKNtv7VS71xZ4MzrIhR1f3c17fieBLeMOE
PB6xtEl/DbUViDXw7u3jn/xcSqbuFDIehAaTKZ9tvvuOdVWtGjS+6ELp71Zvi23P
bRMM78BRvhZ8uysQ4Fbbh4bX/WnFZSTYGhdobog2V8q5O0FFBS7AKCGXlfmcPGwM
dCJunYN5tLZ9p3K+ZDiMNsaq9Js8kE8RFUs/ELVWHcBaXTjq4NyVaPG9vaLegNhI
K2iJROmjRi5oaN0pZqDFObuSmZOLk8BrwbIst6GDs2wgGuDa1Zq0AUftWsVyK/Q1
I6QR8ShEl1JKjRQ1giok/ORucc/sAHph0rKJ0x4bGz8/ovFq9yfmGQGBDZ/SnVis
Z92obdmdP6YhsTbAPVhlqh/+b1PnHPrbF7GwgaX8iAxJCIN+bKRJ7ogYptsYe/N4
stFYg9XCnF7k9lT7GbHHz2gl0bbya0mpGelZ8FwZdIkYGc1w2c9rj1ssR24QrIms
5yMDsEJFNYLZQdqjWKYMPbWRK0ZsfcINNp67Prlm8+xJWSTQJdyCncQCngGKPE25
yEiPWpxLkCx9qXGGW2FAiGbKEFgUUREh+rVRhQYgktqDOb+zxiHAtWE0+P00mXyl
M9/By1i9Y1ExA5i5XoOIQxcLpaGZlJAKH3zq1fJLdW3IFvIME8okhLRALpRylBtf
qy9dSTiSE4poX86XIkoCSXHQoCP9X8dNrVmhvj4/vS2zTvTdCRKOZl2NFalbCSES
DjYInUVKmaRDc+SuPsS98oROeFdLp/85hSTkCTKjEYFFiuVU/ICXJ338qrVGigDZ
uq61ETGcgHaXu5dFGMrm5pnS5QfDTmkDOG+Bqw6KRLOb7dVfYNV7c4Zv8MA/bQjP
j01FhX1F99XSldNlV8jhGFmeb+RHTrQlUrkopPfxtM6nCdmFnb3rs9iR+cRAQl2B
xU1okW8dSk0DNmePg3xeXq/b9nRE4KtQ/XrsEs5IPbB3WS59nR3KJ/Oh2nONN6xY
b6wJiiDdEeeNwkvNozlswiium2bWdzZUtgPzGrg6MvEfo+M3DSN0BBQnKE4uJdpf
huTPRSCYkPV4m09LQUoyRGjBP7AccAMzYjM5wc+I1Ed27Exm84kV1Wbl//vMlukC
0wyAmymjV6KDEqvpp1L68tFnyJYBt08IYtjxzM1+Xb2OAFJeGyfHvi7J5bjwXWGe
5bKJ6F24wOqlmBZjckdN+hJWwmZjZExr/tzRRmj7Hd3IZWZt7GB5XpL/Z/JzBU5B
oYl18EqP8Xa7lNl0zYr39x/aHsZvaaVTttuZVlcuMKpBinffd5iFacd6/GYNUmHI
UJLzC8B0Hm69wvOuAR62y7FvyvsXWdr/cWxLTn5vp/d+Bcf9H+Oc2l/UsxG91kZo
LXNx8cn/B5O+u49h9bY6w64UhmzR73qhicWFqWYg3PfS8QQiItAxniSTRyHPQHTK
BE6y/GiQSz1spGNkQyHgxW/KmMKEAKcskdHZcCkqEVbfG2bPdO76/48b5NXA+Id3
1y/9vvBiVZlw8Ia3DRF3iU3173ZoW91FyxUPAx6kdq9Ecs52mbzAgUF6/PqJ1aek
px3pEAfQyEnKwqatT0O4W/AqEEd6Z169mnTmaAeJj3NMLrlVBPkbxH5tFo5taSFb
dmqCW/2NEyp90bQbDy8Hhtfd0AYRnU2T9euKCdDBTuUplCFFSzicZLx0l5Ddh+Ri
3FjTiplgkSe4sOmUxuDHQTqhOMigOkugKiD/464KhGEQjinx5074kliI1le+DPLD
2ezuJs1zhPR1i0WKM7lr8Gb6SZNI736C5g85zttwAsGa8Kul/NEMyF3bC1taQa97
7IZWeDWzsrzKyib12hvPddPsOEx8mdK7HRm0HL9GLLkHMyAX577jIAWx5uJTVSnq
x6ymKtR4XoUzzHFxcmtI4jmTuuJ1TFAVrAdQ1yFqKG5x8FfKmG1IPpTsmsFDqMRH
YN2qTNpsbnrZ8nPBVmuTc5ONDbHFT4hiouVenD2pItYnvlFwkZJf0mHmLBEslgJ0
F6JQD20Je1i30KlUpqeBmNXfBDilJm3GeMJgtAFpwMk0fWcIys0lN06Oq5zbRIcO
vL3XNmgxjogfEUXIgfCZEjJ7SJscYy/Jy5MzF9Zii4oZQfwV2lpm6pvbIbNeA1h7
WqbWKul4j6ghzT5I8BWg8yC/o/EKty2GvO4m3fbLIKrOjtBA//NomqMo14rdsfaw
A4fAIEM1DiJAzqfKtgaxbHXkgpjzJOBH/QqGVpGOVdlj41lkcsZ3mS6WOpbLJ7aN
2HVQCb8f5E3OUJK/CRsrlijmWYVqlmzaZPICpmBKUdQOoj8OJbtjcDm2xtI+x8kO
1Rw27C79XTvHfgJHmtP5wWz9MUHh6wQECLIu0XIiFLKhXlylPOOO+5QBtQPbRVgs
DCvrHdIT7jLwQHef1mxhtVq1xuUfMWfdDZXCj1gqwCW28B9YXTG/S4XdaiYzsvZH
ZuXZ/rBGMOpTytQ53e/RrIDwpbwGGq5kDvtfxLLKyYwZuQQNFscIqFcBzz26ktgf
saMlM0I0I30QjYxVNwQlvD67nDYoRk3jMnU9R8p4fSg0V/9RCP0IOR2g4GuNj0tn
HCsvSJWw3yaJIRB5nPqig6NlQjxTfVQ25/wI+qg8LI3k4PXOgbkbK0u3wLSlVXPE
ZQ7nx+WXjAMzPJAB8llEZiOT3+2ZCmX7BFk2SeOIvVzGddc/1ckVeoE3w6XaAvdS
vLx8xBHzWqAXy/VEUyOjpIzEbrZx/PURC8cWu/pjnjb+VXT7JQ0i9JkjiYhP19xk
RD9OVhj9nEyOyjzM3yl/fRIwDvTrI/zpPKclKfLQk/DM03+8Ib9qeZjhRWbBzpE6
x4dOywP7dPBuV63xgBUIPlzFCRvBBD259j7b0bnZ+PzuIDXrE/G0MHrqTawUHNlK
VbByc1jFMAMkRGsAibJ4xk37HJ1df6qs0J561FrQMky0r4YojZ6aS7GVjbFJv99P
+esRIl558bh5Qsq+n1R7CK/JoqosYvguzO2pE3sf5y6ssZcWdWTDPrrpIZvD7uDi
sWaNdEvHfYXl5wsVhLoORPmVLvK1w3T5/d0I0y3txFjiAHTQvwdrfz1u+vunejUy
++0HTV86o4zpU8EugsWOvmY3eRVy7aVSiGXU2Swd/W8H5x/fbHVqHQe9AczRQ9sE
2NZAIF3WXnIx67PzdcqpxFARrTujy7cVeyUCk6BlmENAhaNvDLsajNFrnSeuVD8d
4Lsydcrn0Rc2s1Gx3a1xw4I3SJgLc+aVChFMMr5eFKjrWvEu3cEpiaSS3pwjwDxB
175S9r3F3JkZhGmdrZ3XrCGLggNRH54qppJv5I1qIV1U1Lzgcd88mRlc8HGTlI58
J0wfEyrbX8mAwPQlXxCNzvlJvyd0XCOLx4jpDdzpl09BAFg2arOxH+QvcSugEvNT
CKtXOrIhLQOVrPNrjS3MUwHFAWVKlNn/D1Tdkh4XEtCIYc7gM+Qlp0QpjjLMt6qS
AKT486fq3HBACqWEg4lplladJsKkBge00pIxEvlBJh9VetqShqj41BXsHdO11dp3
0+IBJjE0Gn0mYtEQaWgfdBnr6v5gyY/4lq3Ham7hpRURkJMDJp7I+c1+BwP+B8d9
1hKdjXfxD85hLsWgWibEFTIxYLnbqjnGt1AmWluqasTlVn9+qh2AHP9svYOWOVtx
tMb19pKqHCu1/NAf/zUAuFAx3kOxhxKy0BS59kX0PP8aGGPkFI0a8nNMfVtc9dsj
roQz7bY+7JfrKl8A/ZOv2rvvj5C66YSObVcIhdesRUqxxtRwp8R9drv7nm3lFQYA
eD4izw5Hm5lM7Rn6GNEv+sK1aoiv3FE7IU9X8l180HRLe1cnWGt9RZWSkhbMzdRy
aTm14glmlKbSMzxa+8EhV45fWb/e7JjDLW5ZV+H1ZbCCz8CWtzo5ZBFqDsYOOfK6
m11NR8kwlgRDekZkmn9tCUPOqgXkjRbbNEDmGP/SyYjS31Y79GUfEN6bDwbSYCIg
M+dLjkPv9WWVKF5QAd2uqn0S5+CvGdXgzJw8b5RW1rWvSIJiQPosVyUefme1kli6
A6XL+Y/KQTy5K49hlNnzbjfJ5HP/IPBvVCPJvfe05vz1Lw3lkkgtT55W+r047YLg
0aE1FfIJBj+vBMWf1CxohxScq6YCZXoHB8S4TCCQCMaMhGyySJG0Dp58fG1bhe6y
kjWjS81oBU4Woiikcb4IwLeL6MiboQJgdDGtCC2yaNysK3UOsd+xWJpUPelL16hJ
Dfvg6ex9qwEU/31V/8wrZu+QM6/AdgcHCQMyuohlpMAouQkGAptt5OW2Lmoor2h7
4W+Axir8LK+rWBsjZhoeptEF/2Sq8UDX6oAWZEhl15TznPXMw8HwINpDpghR/aNv
yitZD53vEaAY4/4TUvTHjP/ykwGmIbkirgeHnjsZC/7EC3rGNMuEAP6mD9wIkl1+
1uaY0RbkKmQYF2CAWGaHP+64p9j1bqogoUqxhVLSGEJKc26FQk3c0yOsGlB8sPtA
gin9+uA7jzJ0aRasv3Z3PiAStxjVqa8ThhUpDfeEl1FucZ/BOw42wYJ0+eqMW5/0
lEW9uXvh+W86qWVNI5awofmKxBvNl/FF9ioWOipZYm+Q2SwfupnyNzBiGfuatN++
zQwL2d81nsFxuXL1zDYUrrgKICDx+NL4s3Ri3gbu4Zu54zYr7BJdVmVc5hryp0Aw
9MG5yjJkUyOfFK7tCAG5Z2prppcgB7LS0YBni7anaXkZZO176wJJu5mhYL2VHxpU
P0FWMa7JPSPBZd2UI5y61JXlouIA8mBzkVDsUo08QV1u11ZYAE2mJz8dJu5M6Yjk
n5pkKGWG1bi7TDYVA2YcUxv7Me+Z3FL+WPDyVpwMsAvBOur221oj2u056P68QhMc
O137i/3GRpMLitHmX5SgBtx4wKsWiYwm8fdH/gTCBvYJ0W58Vs91WPQgOc/ANwB9
hTbxkOWKBunMnYa51InqrrNfASSctkm8K04umvlN8p7tBwB/W6ycNKb4/kKyYden
GvEvulrK/MX4gyk45azovCXsIGejlIx2yxa60EwrfNsjBdHOKpK7U2CXHjRNiWCT
tLTTLAXxBZmFp7SZ4DnuyHHFx0MSoQg/3yT7Uge/GMSTW4D9XC6de940wbFUrrGR
w9jq/FdFqdKEwm8zuTAHyNHiN4/6qQMtGIzIJpw3oYilhQPpQqCoRi05H3cVYtQs
KW5Sx1gg4F6TCPQptW7ijh/7n3u3wWc9UCB8VmB06daw9jRK9p7Tq5v7xYcEuoht
xRCwZwlv9xI8ykyO/JpLTNX9ehAk3HZv+wu2Umzs06UDLaX+OjUCcEHplf2tcKoq
9uGK61bJUnIm1yXQp+kCjbzj7cYIEJgD/6u5kwqC5gWyFfNhmUVLX1KjMjG0mY+7
kOnGvkgk/jsKTnkolfHhRgVEaHSGDTEthEGqcRPT7p14adqpzbcH5MoESA1Veavq
M1W6YalQyHnXhLFJA6JcGkTGb76OYEoHJd1oFRKeAZS7DcQdFZI48yxUfHHBx2JJ
BNiomJn2fsS63wobiCaNRwW+p+01dCy2aTcCIGqZ/i5IxzDVNGxuv26QklrOvHyx
MgVkGtGz1M7XnC+g7qM6N7U07uZ4VeVGaLUZ9FWrnPu+ZMcEiWgK4J3mMEFb7UWN
lZYcqHDh0BqXbP3nree1Vv0ys4wOoR2sLCdHaw+JGJaEWcgbQUTCUtwP5CojmcRS
uw6sB/5knzGuTBvQhhXcbRM7H0AK5RpIQT2PtqAgcDDy/ln4UskyRAlt4iH0Nj+n
R008rbEuQiripu7gWyC1ptjMVUSqI16l1mPizNn9NWPQ5wYA9PMufkFv9KWAy4Kh
vqXbwEEc3oDhMBjn7YOx6XqLYfg6osayyARnNtpHsLH4kyfF8sCAAIoc6vjhrA4s
YhiqehepIxh/FkU0zCrdYjYZDY6zzSdymMk/GCXR8n5FZ81/kI5sV/zqpoKo3Zr6
PFAHJFGpIvkLSOezI9mL3l8sjEHe/Ko7X2O4+hOmWLCL3xBqJDMRijHISeiP2ja5
CuNbHmkJ+YwQwveD95AoyNXHtDbz7WCeiu5QAvOq3Ra4FfJfJvdZWqkswWGa6PpC
LkruLjQZkEf0dzaA9+FuDzit4mCatOBT/Koa8XSyGkhGFheJ597OlyjI/X74xziy
amT6CTrTLL6gkM9ZA1uA1lN/gs+lng/iSov0x/Lyjj1w0Av0OYSYLt6wnrRirWEV
NxTzC87bUOyc9t2nlhbo+OR3x9wqkZ90QSPkiMC6cYovxu7rxBbfOVAZbZTgPNkV
txqWCPppwV65qwO5nslriudXh+BdEyscF+w9fbGi/qjZXqsBQxdedYd0n1W6TxC6
dmQ+TQzd+/eyZxaL5NhxfKmcwTgjlOcAe49Rmn+AY81Nl3+X28FWTc3wgWIyhjOv
EtpO666PDRspLgeVykAWvmymd39GIULk3CED5qVjN86gVXDqprhkoSjOG7cVCbPG
7w+76iX9vLbFjRMPpWpyUkTCYzJgWhO2N1mD1i1LoBT4xQbCmY+XnJiiP2KqC3gG
SQRlpNn/ZTHGlSgBseSa8DopwJpxhmqTOdBLpCWCDyMGj+pyq7msEDC5DUnowhpF
93MgO+QXm31chHN54zqt4MPknA8V1iGv0MU1aSU7cjhYcxSLvQpy54omwVfExiIy
YuBxnZlwBf1J9CBWZOGpNH4oD74rQhVBh0GH4dq6esFdw+4nIeN8tWXD4tYEHqbq
qPC9p2EnxCuALUaqQuPndzP6WQznkyCxbf5EapyE5HXUJ9e+onp4KnlLVkxw3mKv
ffR1G4AATKxoHIvxCINk10O1jaFO5/grpvUzz97UCckxiEf7qB/TPR9oJyHSlAPs
9auejn7oCokby4Ol9H1V5YwL4GifYVEu2j5T21PYDo0W5DN9XG/nNREREyxrKDbw
4tCpu1/xIJRhID0l2yFHrrY+DyiWmLB+xeAomp1zauNFMWStLcvE2NAf2JkTjp5A
yHOIH75IfCIyEx2g3ylVi+M0fn9osiaSwjsIHkoGlrk3/Fj2znyuNDmzM4GSCb09
WrDd0mQgbX05NEZ6i67SbqyYZmghcgq4toJ+PcWCluIh/mZ0W0HEuYHc43RAXgmD
LnwCx8eK0CxCQ8vmhsZ5OHuVpDdLCR5//tGDc/RERFxyrVnK9gWcg5IDijJ4SmO/
jc1oGfN22/LM4ukIInIJ7zzTKJuFmV80eK1I62DIJEnql8FeLb9+aKRCZEkKM3NM
207bFvFtSEVAdVJYQJWvn8QB/LJbGKF1dYIQAof/ecsrr03Nrw+nXgm0jT3ZdeyS
VIC5/YgTeNseK4RKm702wLcbsEtLeFuAo1okbdB6OwgVP5fAalXJFcvdKHJqbbXr
wGEzkiAHXja7JBIBY/jyrU4dKC8Lb3y421s33ItAxTLlqY2FmLMPPWDU7Ba2SO7S
Yrr0Tht6unCL+DrJCehtxeB16QWbfX11KPNF3DUqXS5pgKuFQ+cB8TU4jnqiUDDr
UiAKV23k7zoM3z+xX1saUDKjSI76fDEf/9Dn+vzagn/2lSUkqP3ZdNsmAs7RPMaQ
8GdAHeF0m+d+h5GqZJWFFlyODRHVzauwg2KMXd559VjtS9jpv5Yk/dThgcG2rPup
RNJsHP85KcrwgwQDihd4LdM8X/+IjAnJaeveFO1AO3oGjToQYn4foPtI5MoyvYv7
q6GX+XeLbVj6bZi/7DUDgHQBx2c61BBXyoIU5bBPN2dTW0sTaeYeqqKDb4QQD+ZO
BlypHLYCppmscvoySGNURVILBhG8h7BLofQyjzoc+cjRf40oMpz5Xk5Zb6bt6sgx
SV1Lb3paSat406Hzia+tkmb3/gTe1IRWgWQ2JrDUH7fNNOycC1Wp0KQYjHWjaGy5
Sdw1CJBdx80pS8h/7dbmh8a1vQzDfhu4kw50f2bxf7osyY/KivY0BCI3zDbTfdA4
gyZaZ2aOCq0oLmka58hAw55w/z/8IhGJvNI+nIiEL7iyJC6SY4gzND/YX1JWHGPU
DEFVrUalbXJGYSMkiIvYVG2+YQzoYIgRjCF4Gqov/+F7D+2OcExT373PFsmDvTEJ
TeOoSw5MCMzv/0EiEAdQInVeTwg1nwMuj+IVg5gf7uelhQkUc/f7BpR9xqheJVOE
+XnNTlhOXPu+N1mhlyBd2qGRGP+mnI7/UzMQfyxQCNaw3SZs3gOGAuu4XQ8nhR1+
E1UDcPyLIT6hRzWu1CfzHwhlJ/YjXibowbDNA5WAs4dtBiQN5EtpMN0Ft5Lr6bOl
QfBhYh/09DQbt1REeZZtrmekUNCcHSf4JfyMXkgjRTFQVlv9ohg3SJx3DHvPryMR
774943z5BX5BwbVdhGUhjCUlM/SloACZJls3L2vpL2BhxHlrySCOUjeKffMabBGG
XL3w4YSMotvkiMoGlIivxjJK0KERO487gepAl3+btgAsKMagcTuLqBO5B0mbfqx3
iVIa9BiFfDRJTEmnye365dqR4WCC/96fzxj3XP6AzWhdfeLIp+Kn8sftlr0QW96j
0vu/L6yNzpNlV065lgPYOjrPrKRrXNNVYijPLLR27sWsejSR6/XRUiqqSOmcYo8M
6oqgthUqMU2HXsMzI4j+jtdvJP/C1EgESXbnvWAuWpBvImjCKgA5HGx8efjKEM9l
5pnKvxxCQnTevuNTZyyg6pYcnrnpaGM9G2G3KeK+nNoegb0UlyBJV08qL/GGCuRG
ZlVtPtvtaxTfICmyixrcrWz5BkHfY20J45qgDhZViO9ttSdVyhskPx9EszVW25yu
pnMTzzzZTr6ZE9lPruAjwEJs0pPecg208Ig3JNw0jWaU49YoEfw9qRieXSY3uHuZ
b0vBzR2ZhpFszrYagvUuC3UOyAfABHWsIza6m6uZpM4IIyw4IShaB7JMHJYhBLDD
1kfioY8fWm/uJLhVxK2o8A9FsqBKlrM3KxnicMVIWYDduIldomTIM8pAInA1QAND
4OAps1hcE9yBcZiLoT7vmxaOB0C94SKMu+09pwXBS0Onj5u00DbG0D8QMU9blLPo
MAg8H1v91Tb/WfN3H7BCsDERyRtAJaFDhk8r6Dq8UyZeI3ZZLZNuZX8kW5kC8dGZ
7CGnHpIx+cYmooZn522k4wfszhT7NWjbio42h+h9L0vp7x1anq+dYmVT3oIXEzf0
jkiaa6uwv0oO62qNmbRmpyOZHPxZ2BEqfzWG6/vblgY7hHkRWlD3r/+6/Tpf81jY
qbnI00R0eG4XO/6KzpA+0Z8xkSiA0PCw8dpreFNr/Bf+9hdIl7gdd0h+O/f4cn/I
JIfvroDSsCvzrdE8pOPXYlr8y0GulxRISUoTTsKOTOmND51SWY38E6ZU/uHV886m
yhVI4eGeerILBf/Et92J/R3+U0Oh00befiXF0j4XaXEnu7VobbiRhm6g0xE7mrbt
9fuFplvHufk5IrmNI3NtqbamLIu0TVcoq1MdZ1VcX4boSNZn4KBOs/kttDUhNFnJ
+mSuGJi8RzMXXxjl6Zf6sZKd1w4QZpccQCCtxy7m/Dcem8qLASi0HrE9MlzQHFkc
3daLu9OXQu7Pr9DeoI20z7CsRifydifY88QQgT6S9sIQNBuvOgcG3rEBzcWX/zKn
tDAKy/P0o4HxAD77LGV2ssVJi1vNfmgLldhgXrSnOoYr9Cc/SMJ6vhM+o0eO2uzf
QJxlDKXCcz8wlk6dazJ6+XJbCJlJuND3q0HbZl3jFcJkv6hdmtqD2iGajy350iCF
irQ9YtXxR24GJgZ8crgnebXhLzlSiIiYD4xrnf3amYDRCuShdZAVMJYchGAOXcue
dSNly8+TJZVaBerEdt8lkVO5I9Ts2mPZEZCNJJLD4HoJK15IjLEB/H4wuyohN0xx
DszTxjtJcvd3AwRQxnR9ko2G7F0GfZKHIPMMB2xdYl7827xzO0MeHcgQvb9CLzsZ
CrbARCVOZXFt87PmoVUfpchJUyNffDS3Rnu6OAqpw7jJfhiTynv2wXIj96kpHyli
zCxBnL1ddnEfdvo6l/anfkjyu8gI7dUv06SDYG8Y3NhJUKlpGE00QpW6jRXuRIcI
mhQ9vt0AMFDGwr9VfcuLnm/xtYVCQN+i+HTlXeuUVB+Nh3VroZf+o/vMxP9Dmgsj
qKAo2iiS3OlhJsynAvU773lE3lVMEcnCZp5Y0URXcRG+jTtk2SwxRnYhntA29SDC
0fKAXbCZUb0sCGi9D9GEvGkVVbViymV+JAFGwMWaJ+45FTQ1iWSmwa/J6mujXdQ4
ikF7LYI1S3R7Qv8/tVck50QcAzz/X6R25rHADz2KwYBHNaOQywp8UVvncmLOEzoT
J/lzVMTmyCd5iEJB2Cw2RoZWpBVDhjhZBOBZh2WMaP5JExE0maksU5gM9fJU+MP2
pJAYFaM2DfexFkySAp0xugBoHVKiCvaVZZHZTLYAVfEKh/8GAbElomCMM0y33SMe
ptR2d9E92FFxEqEcNbfOL03fVuFNMh26meohEVo0UVxvUEA0vC7dnWL1EMxIwpSY
0LffzHrhxM484RC0QfDLvqJgfKWfB4qWGq/VODZ96Q24MhcAQr+YuuAN9Du8SE7g
NHBPYPOsuyLSYq2UwoEpIln+EuScKRoVEgI0ycIqpncrH1k+PDnmTrZl83bdRdJV
WudWgrgP0eubxV9xBw9nwQQWcj8HjAE+3fnNKQrGrJ5iL3o1NqtqBKDcY1a+mnvI
cM2lCam8qw8d/g9KFzM/3AsXCXlvBeysnQNF+AMxiGurnY5Fc/3Jp2mByQbLNV9e
F9ClornLFLcgfi64rh6/buh/KI/nFVH8LMHVnBOLheXL5FrNrnp43raJ0eAx6wZ1
vIyNE4pajc4zub1jzd2ryIRid2rElMJiY/880YHXC0xKiHkbWBPsoiAHw2zePn68
EGBAeSWc6XyIo4goKTd6YWFb65Zm8mxAnhyj8YnYO9HoHDxr0zK8tqapJ5XFmTWw
VdfTMD/+dYjYqTlNgIPAZ28cU2qR3jl3a2N3XiqzhhqKgQ8KPDJu1ZWGXot4QOSw
MSRfnMK10hclg7OuJumayN2NPWrA1b4zjgS4zQYrjVkyUIXlPc6H+zGBbpCkf6jB
zU1S8fcF421ectOFBGqor8cxm2b/rR4tkbXb3VCtslHf0kdq5QOMW0GpN6A4IfWm
ojNIeVID8AOAdhj7LOvNkOKbKD0FVcf1oJdTOd15D+ofP8X3oX9Tt8kQX0qd//7b
j0rqnR6747xHqHC17wMclAmo5qJ/3bkhsM/GOYiX4OtNyByFYWWC8/bQ7W84Au+q
reLwyJnaJKMJKuKz4xBod14J1XQZw7XjdGgiaB0d5N7b//tzr2iQdZtkTzYnRPPc
gjjIeQ6IuLKC5Frsgp68mNxU/8X06iaFw/qjjjUqPtzelxs3NGzi7m7wMJyGoqkm
Ae0+/rMGQRB7LPuaOsJG3rKhUagBItuLPxHtRXhAOTChzwcydeEYIQVc70XpmSPs
gT33u2rg4HzO/6oD6V4QGmSXDWJV3GfJZgCseo+0eboCcS1kPaWraXLtn4ix6z0y
pWPnliFUWukQl6zvyDf8u/Q8wPMShKrNK2VVNxce0vV7llYw2qh0NALpzRS3HWoV
55gQVuk1IvHJpV2u+IRbgVBe95ZRNgVqXt/Ib/HM4WB9IirNwsMqnBylQ8Yf0v1w
DI/7f5Z+edykMieWl5Zd0zJjnIP7saJCgxVh+rz6XuzNIIeBi680nNT9zFfL/h+6
jfzk2j/vWnky5Ok1eK0qyvgRtbA0agaGDHqQOefLUIiBlVViyX+JIbMY0j8/kr7u
ZmhSVvAKMUN3Stf/tbMPLCrCiTvaFeNOkZbvBiSd7Ng69IPtbLUAZq1VizkMejp1
TDh6XiCVoCqwu5H1O4ssJEOHxtuFEB9AIZHv+VIsUnBX91oMAGLAm3eQB9SjFK3q
C3b1LbV5gkBoJcujzmRTmvm0MmIU5SPEtiHWzlkmGDhuFde3YxkAlSyS34V74K7n
NiSvU3FBGABPt6dD34bYAoNOwEJ+mu63c26J+luK1mNSNdfXEe5Ldkiqvnc69zsD
NxNKSOH0V+z7HsWFsGIa6Rfnc6C7BaigdU/IUvEqjog19LuLiw/W04wJjnqO35RW
MFa8ngvNAQX+wY5rEBan7NEcFL9tWHFKzdVSawqrCHdep92WRspAMMc0DsbaaZbE
aHvufhBvr8cwnfZOW7H+kBJoDgJGYwdXJ6k3G2xMQUBeX8ZmKgpYrz8g9XYNa3Tp
HJyC7i1hVnR1laTxdToyCJGeOP5OJeNCjgjjVxV9xUa4hYpZt98spgbk2XQuPfbt
aRLRUscgK94gwBnGdeusHP6IkjNPJi7DhwwMrWVPg4lNLTw0HTOVOYAIKpxYCLd4
lPCQyNcsPt5Pns+KVtUBbc+FIA+yNBIGVQXHOWDz7yg0JrBuUuw9vmlwqjAWAKUv
QS4Gj8C57bc+1Pe1IUubJBum7ovzK7rBMFTneSGGCjsq4/7gGYuXyeWKsfROj6R7
2vSCRUY3htrYhn4r2gUkIat5v7g2BMxC3cFLdV7EPIS51qmBqTALrTAr8dP90XP0
u/lhuaAHWFRLzHMV1eDvnV2HOqSwFN5YxbUNs3+7AfmsVwBK11sY0WYxkTQWn37p
6C/XnnGUstI928T7e5RuqjbjiDLZCr9U/bQ+aUTpIPCPjS3vXiptX7dQ/dl+WWaa
KzyCFF2msbJgLkP2Hz9xU56AT7yRka3FOBjSqhwOP2T5uctG/bWv0qvX5Z3+b1Ai
9d0MhcPZkdA98L/LOen12iVeFBt8L9g6/bKsIIlw9+m3U1l4cGU7YXm1CBPj3b1D
ZfbuLkrOW6irmgvaDD+bwvRWP+5bsOHt+dZbHmrMFTPldabaEp+rFT60LCy7xGXX
6A9dZHOClTmIjqISKa5Y/OSfsj8QlO8uhAdbN1oBjdjqItWsqPWp+M3Gc96Gmgyp
sD7RK01MUw3BDuMWQ6GBvuWm99VkhgfEGfVV80bLxv/NywjGJGfQuxWh+d2igMD1
8sYA0+J8IvDG2j+7AKvR8mWI5pIbEW8pH/1VPNJh++ctA2mcIPL6c1l/H1YW/l46
j2sQTorysAtQn5uE+dNKHKOhbI2T9IulBYJcvq8tEvSffy+Q7GncQp66awQLuEgP
zDO/MfPm///CV71cXJDoXD84M0SbXp35o4nSTeh/BIRKp4/GuV6T37ApoY83RUaa
efoap1iGItPpVlIHcOMnqR0APJE3e2wMI7e0EJDyi5FS0u3U9Zgml7yvjNeMz3iM
qd9Yrx81ThKkPC04G1/Zkm7IpJ54CcyMe3fTgjfnhu55g0pmgZdySge5+Whugu13
KgQJT/sx7j0KTn5/9ffGfAudRhTYiRmndIwYIfHzBTA6QJrtwAcaOymLSQvLRRhz
Z13K3/zyAGx6fKyqo2JWSEMuAxJArOxGRSrZ3cXOK022N27m3PDcQpZSm1lYBRfS
sOzAjk96s6lFtYfbV6OEKYtnHVJKyFar7W3Iy/LiJdVMRLWaflrZo0OjYuSdfuGt
lUBpeJtcTukhso7FNgHBuYHvb1rnm4GFNbNlRJNvoU64lF9gsu6Nj3tQVwEFbjIO
zVgG2gHTWIxZxjKdgjNyFw2l6FoK6B9OeUWV0+6Hu1nGw2WDOosIF7eVQrp2/91q
q8rttRmS3F67IkxhL/k6YILWd5uw8GQM6RGBgqvmsOi3qzlFXm/f5Ihe/R1bpGcE
41fsddXyHMzXcLdOgksLB6Rg0pc4HckJdhoUa7lPqECWSs9HO7kYnLxq0bXlJ+jr
zH7MR0zf8cV24xqcYD7WIQYF2DTaPDm/dencqmgJFacDawB4hWLQwo6laCktQqsp
7HRK1ZtE9VLy9oh9s41jcZ0PgsM9ZHx2ooZRiXb2B8DaRejhy/9CstKgdKIeuOjO
C8Jg2GtByIyo+mrD/RzkRDHFExY73PH95IvwIcwjBVEIEneMtF9MbnkFrgIJDDvS
oYIKAvO8dt1gmAA56e1d1TELkyPurO/xDBBUVMVHlC4bc/Ntm6T8SwW3Oy5JXAjB
0WUcPl+PkD0KNQzQRfvmFkE7GeMh5uh+SXYxlru2VCz7eYPN9GmTANLef/FduoZS
n3D6iOlQy2uQY2GvwhEh8i4mO6Pw73JXNsIGFLFR6WNkp3kUcKHDZgZnlfAw4UKX
T7UqPZd2+o3GQhWqdeJXWYz2sNibO6bK5KpROjrBDXBPriJiLjSK5xm91TCiTIgg
MAwfWtM7FHuOQGH9f8C9VRPRPwch8yUs13TMpgAUBSP1YVAn3XQI7HwHs5iNJYyZ
FmuKoFO20Jcy/OEKAX9n8K2bW3tl6fEWPph84xCk498w2CQbBoGj5nBH9spPOS3x
nFZl1EF/HDr7ufGRcoq1zyFCFT4/laRR4/03Q7cTkmN7XKjvd4fPI16U7YN+ShqR
f98ua6grk1gIBVHFl5+GxxruW/sHiqdha5Rm57cd1LtYxZGviuWsR/jIyV7bYIxt
4jyN4GWCzUV/8WKqyu2rkwXvrqYF7P2ORLQQIKFeFJIfyCGjRXH6t54HFBG2JyIw
G4HL46P++z7FUQjlJEpBn7aHKUKefzJ+j6JI6PQhE5X7hEmAau9kp+wcnNPPYVo4
olAmPV/Yll9WKifCXP/BuNnFupZVORYpyUlxTYnWkoKCx+lcR5ruYYbCb/F17c7l
NjhdrYfleoXr1Vq+30GGZfcF6BM0NZ+nRlh8tMi/H9Via9f053NhHgld6j/DQc96
3nh+ox4CKuLyr2tnjQj/H4gkiu2u1Sg2cJUYW4alvrHyjhoGCb78kNN25FX2I1lg
zM5m0bZeziUV4CvcTwUPhz9jrt6A/TTaP7yEjJyFzppDk0ji+iWZSLAWpJUeFyue
WHRJD4Rq/KYTrH6mvCU24hc0CgmslmpPreeQdFXmtqBcoONPRbpu4HIZ3hHsD7NV
10HqpQqz5AwPM7CgRPPWYjcMWFgMjReMTGM5SVgKB2zUuyACeMzkHuk5g6wFufAw
NbRvYuJZ1VeauVUfkwHlIt6V+riMyA1xCToJXCJ3M0qrcUWEY9a4MLTcCrIsgGHH
Q6uBELetSgv17mCtJw6KYwSuX5g0c4NoRUAy+UT2zW12jGtWPM+UMFi8C/Q9u19d
5jZj47y4HokrGWqTT39CvGbAmQ3a9wv7coWhhqHdiEMwrEYiS7iIKDb1m5ihTDVJ
xEnOkK+DyMvrv18jMG6J4ujNPXPE+j6d1UlvWRTtwb3wqm9Prb9DbDhB0Sx6Ydvn
eikHXRBieNpJePI+jGymyU3Dkm0Up7glVU59v4BSQck4HzDLz9ZiY0B8Iz/GRbA8
qgzNTzDgQWt3+2iNhylhOp4oIafmVwYkkUrd0qfSDv1JCism92yDlDAFJ53G1Adi
krEDONVY3c927/MkOrAv1eevCyCPh5WRXbBKhv2fDO/Bhu0PmVGrc65WxP33k40f
ame73cUVPmidGxNBP57Nt6Bnliel43WTq87hFgwuBTAUXX7iPFDlPmZCPZhd9h+z
Rq9d/QTnxvD08+o8IrZjU3mdWzu2Z4Aa8HMLj3qdPoRkzDp0M51UOny8uocZ2V8R
F5ijWp91HxieW2gpXSTZGsf3WcFiYmKIHTYJAtz7NktFgfbSJ9Db1oFGE0o9Kzbo
bGu8bLDLsQjQJEvaKOk0q0gQakq2D0lvQWq5iMIHRThhueUxZmlo6YUuyookqDm+
lNrt92ucuxdnWWLoWDohr55y75jMe54zfwALc1px7HrIbJNHpUVccwEnMQEGvzhs
tZkytLawgekEQklHuvJ1O/FpQDvZ7e+eMmozET8KgaAwgCvr5Z7KXsnMlB1Cfv0o
TJQKik6nPR714LtCyFV1mbJOeosVOClINhXAYRcEehwEVdOx7XZ6ej+PB2pbFgX5
ta/XDUs86drtIftmLu+Y+aKfF+3zRNspF59S9YVVFA0y7nofZAuvwpAgd0bKipI+
1anbezwqiI9brp76J6ojJa++VAlWVG3rioVfJ76YtNgUBY1jqPpzd1sztFKl+LhP
GfRMOJ5UedkBRICenF+YK+m/l6aEo8iyc0ZY56/FaOsDfT8KKNWChjQEd0pNAcXF
9K5E0dMdHlh8vl+kWiDCCc6Y1/CS/gu45BsONDCqaZtY5Kd46S4QVb9dDY6Y6GH8
1AUfGBxvteXKZn8i7tcHxyGWLvTguuawqmc1TpoIx72VhjE5UfdEqskQPQs5lLdP
pAO4koK+P31TNXTSH5ufoVmSe2pJlghRzbfftgO7z5tCKnnUOZiuoN7WbxK9apVx
/qwvtyLirenpnSByKg2r68GQCsqtpjWk1KX33J7lVFBl92Z5ZTlbg4/S+tIVU2EH
jwmcvHyRkBR2jZFTs9cFUKDJX75kPc2DWybI0LdCaX4ftWrGBjiIy8LueKx8M2xV
90ZHxF/ln/4km+olgp2r8BCc/wTVpHv5loMV9iVV5dBNQrKp4fiq89Tl1MJv+hQG
ERSE1gEk3ZIaipdprnlFjIDc3FkqnE9E5Av676Icwhu1O8DsvaXbvUOCljsS4s3Y
mFQaYgAKfTosiNM+0h5LtIBIh3RJWsTBcBXVfYpdJrHRzqaKZAhILMCVy1QiFq4Z
k1tatjMizuWJI0K8He7n2ZDMYT4GGsPN2FFkgQO8mBiJPJ/gb7g/7vw9OgEnUm0+
7Piss1g1U4AdYteBaQGMmJ32mQfeu8wzzypXMayT7MJUp9LWEYhlhUWYjKQ6E0sj
wfclv/0AM9MFK88T9fB5/ZqSF6nogke91nSw9kBIlKh0xR3zoHaIkC/tb21SqjGs
pKcvjn85agFN7AjadLWfXiaZSQ/1kZG3Ma0LB5WthvPkjAfx+c0CKlXBhXvlBvrD
+ZwqddHm7WmFhevfDBWYGdQzvqeseIVtJ1t1afRvX1juhpO9A5Iq8Ajidmj8C8P/
nraLlFTEqqsky7ll2pEtFLgQY+r9vDWJNk9pGWTv76GH3bBEbLJPRBJnum6qJXQQ
epPgb/w2kBC232s0W0PgucL2fBgisPqi/o+LptA+/37yo1RH7DVMmlg7KvXM3pXH
RKqTjdnHnMAqaNF0zM1m1Fu/VjnoNJidZZfIRnwNFuRlXqv6ChrWYyRb6Ir/2juz
6fwFyanB9KMLNwjzDyLSOliaWj+r+Ge3wPsLDQGP6Z5CLR5kYqy02YJExHw0VSho
hnDkeIiaub4GEnenawI9B75P0ITQM4KbqzS82hZgs5lfzf8in9/cB2xvwCgHapuF
Uc8DqX5uSYtjGj7zfC23lzdj4SWgOvfgp6S5CgQAVYzVj1zBsC+8GnstQ+NfAAbv
FqvDyl3RGDVTGuo7NKDi2+5PEEXmwlzo1AEWpUo+rt270uk0YhOeywyfR3cec2mK
NJo1TAsdd0K2AfKSWeHFOMQKHenbUMAySRqlga/yhRqbacQjSEldx/QHFxS0dHyB
7u5l2XzemR2/GLndyfmH0WrTq5mCBFjhZuztheWB0JSTl8Jivxp10v8rTFAKrIYh
WVHRyLv69+ZsUjbGX/8PbJ1tkSPRmR+serFQbw/KpbbJwyyiLRFMHru01BYT+ZRH
hT76IkkX+jXprL/TYVRnV81kbSN4Qa/qu2ucHCadxW7NN8cInVE93M2cuxG0byTj
5twGhdexHAgfrKaa39ZpY7gluwAJ0oavwcI9QxFx0RseR1DqNUMJa4TEKLkgi31d
3BeCkvdKGLlpbqUZDK9bORFxnpnwlYof7iSw+2ZIwW53CcQ2aSmxX2Zk+I6uBKHc
2fWCXZDAz6W/UqXWMrk2AfgVKIITOuongOUdk9ft6u9jqn6HY4PX9tBb5FU/rCCi
G0QjbvGgdZbvmkETqUTEf0puHk7EAYJgYCKxECYo2MmstyDs8S/24C/yauWakSxb
8xyaQTh+gAL39tWQO1LuCsedoh+3fESAbWylX/vp3CHjL6pmTEv2gImKqIVFscKw
nWbPjmTqoEkiqUNpOiRyLpbo0Do4vMcN0lpMrRlhynWs/TuCvrqkWW2UcNJJTcml
fi8Hz43BSmhsRV1xtPVq0oOKkds7o1A1Q4M1aCvq1Ta83pZNB0XiTyD/SBDhe9G3
OrJYw7j/mG32DESJj27o08OmW4uhWbvrk1AW/QnTQKMS7mW1238PsZwMlPUjbtPt
MmmyvEXd1/iiFgUMuBsshr3jZFIrAjPpw8vqMbKPq51rFiknOzHkYFQSnuo/7nk4
iClzBt6Hlnm6UsJ3D0pMYLtxg/LfvtnU8j+rkTGfKv8tlppVuLfFGwQz4ZfdXTV7
pkxcGh9UFzAxjkVGdDnrpWemhjBjmJTFt/9oCt08vuXm2uD0wCPC/75MbCJmTau8
I7ClEe/wh9XBj2zZ6ljb5HHwMh4COQZlFdPvL68GjL1mbeC5un3wvrqq3BquS0gp
SI90EPFYE9gpiVPz65hg07vegoCzemSm/kAH7fOTFIZK4pB285OeDbD6A78OuRSa
5Tipuw5rBTrZ+1Zv/lEjliyEQQWfN6p6Z+SdX4Cv/QJ7EhBFXxIp3/YnwyXHWtXI
cIW2514+PKGtP8SbJec86gzuabczfmfljTFlNr9D1SONal7uIqXkGRpb8cwEL3FT
7Tm5YspE1INoTroQhE4UAyEfsQzLy6BDMXV6xJXIrH7oC88+HNNsTpUgnPxWYDzn
gQMIxv/hq+BxWqa6U5eTFn1R/zxHOmlRNTAhDpQKpVJ/4KUAt0hO/9+xDzF7zST+
DzoAPXEgTsm3F/5bFy4dgcAQHLSGiCy0RknwszcwG8J3b2WSe8XVFianHIKFVGyO
uK0ZGuo++navRmYst+BqKOE+7fAc55WWT1DBuqKO4FJloAaIgAwKyFaiYNMm9SLH
zWGIgJ32KDlF4RBdJhw43CsOcLKdzpl86dBSEyKkVSNCRvfHbLZL3BS2goUr6zMG
bVysVRnS14qqTQgGYAgdim6z3U3SrS4AeJbJrQR7xl4//lH4VehZCXaGd7MkrCcZ
jJP2UAsf67XzOMqyvMKFYCBXNYCU54NisRzRe3aMNplClcbt9kJ8Fl7ECRWjpH5N
M5W6VVjLsW/MgV6n8e4y6gH3HS6NsmOfAd33TuWjuBIj0Eqe+vaxqVWuB7fdfU2I
pvnh4FiQlpGF1vMmkszysCYxKim37gK0CSSIJTE3ZSuNZXjlj1o+ioVUt8W9dBF5
VpmjCPa0UHgDeWAIZP9uR3k4wQ1KCyJqa1S8YF6xCojBkvGCVhkPO/5Z4RfEIS8I
XEzAM5jd2jm3f3nd1Bs64cbMZGIbTOgNAv138FRxfElZGo0NGRzpwGugO+5K7hFp
pWuiEB2S+IkB0QukQN8evYvJrm849qCrkN1r97BDu2WkhQzkRY0vAPKN0GkRj345
BneFY1oirC65440FPZGXyURuIJ6W90gQ+LCnhnbsxmvvbLADmsK9ap9yV3RdHMS0
3QyMYGMMzJ1GaJlvOoecuQcde+3N+8Gib4jWEu2xBmAz3I83G4EhjELouCBswVXo
K4QVDiE6ZXSV1NoO0YndWO/Gd8xtKlG2PFcD2DY/dKHhZmXHbLkMAF+842IyenW3
jTtqOlX9Qn1GhvbPxMYBd7Gq3MIcA64RVWpYPtdpGwLpqoaWQcWSfyouWKddCxJq
dBIlWJqgofdXtmFRpwhHBHEx/LCGcVa6XVc6hkxVBRJMKq3De2LM9UGxbtKYH9tB
IB8Ib08KwVysufNS6SdtPvdNFAlUQkUFHVO9CNygrfEEusdsq/+oGBuDEOX3V9LR
k1+PwznEsgylRWSEUeZPv9IdDNVXTo88J5zmSALC12RhRO/GpHTQCTzwsZq50vTh
ldLDebA1/tSMIPhTfCTnxFu2ZfxppCr/Gz7uJWTrMocQxUm8TsRMcXOs5B9HjzHB
0+JOzgCz+yCtqCk2StNxcCb8rZnTE+MawRvaPHR/Ux7wYV0Qs/c7Ti22/R7WL1XN
qZ6V7OVVNI0dEANaeeyh2OXdFhgX7CbrDIShoZF0CrDfFrIIUDitRZKCyRM1Gll/
j++5BVrJPzBvG634/Ed5NGeOcityj0DKVDmnDp/lp/wPwNyiKAiKuMeiqZRrLxZT
QpZGSFGo0/3M4socRnwPvaqDfgttBqvzou4g+/SAsU1sZrUc6U5fItfWOjKkxOGl
Cl6YMDGK49iB5lfRJ7fwNhteYTgcELXaysSAPJN0H7q41YrG20tfNf4IgI61HtSA
wqWbPpKleCXtbDNJEsxMYEDnjz3zys7vxprjo6x4KaJiZ8havE1Y+FN4aAlSHAhD
NREiPlalGxbR7ao6DflGcozf7r3/K8RxpcdBNc8bvaL5JzZolYtAtqbRO+31NFOZ
t7PpOumb30iTif+MM0W4TivTsE7sySkxNf6L50WKu7LRqWK6ZO1tJLxlu6ag+v2H
1hbSWMLsjEbPnW8cB4UMxmevQSn0AdOSGTLAuzi7RNU6yVhrxawJricBObEd+IAs
qONt4AbSX9RBIGLXqm0pJmooL83fhpDYf5jXEUyjlq7p06vJ5j7ubqMWtobOLep8
QDqL/789hHLNrRMNDSSHibdAzdiMd2K/XkdAawBQbFfex36TUqGTmg3g8aSVhkHC
GJFso0vqDlGE5OWSvgPwlrhQ3IxbqECAveF8cjFhaOXQr7xFPRtCLPy2hfPyqdVx
YRt6MpSymdsn/EV3sJfUOlrM2eUFNo61X98g5my8sNzCC+JpdiVZJfnM5wcvAEuB
pvzYGwcDm1a8CoZwvQKrVYbcSJ2wrR56mRZHurSESynWkJBca9RRbl8xVlbOLnx3
Mljshr8YwOGQG/msePx2zbHy1+lWm2+ajCgMXiTv62eM1+pfKCVU/o9iZtEtRDw+
d1nCLQ3r7D5fspxGSRD7hoMTMk6pckullhfKF4KevlT2HJDGPjfdmND1fpGftQ7R
ciQrv9MAtjNjSyDSJQkZ1WT9nlTEHqFB940fzSeN76JXlsy8R3Nf8mhy2DZtrPAn
zwvgFv3gR3rzpcl91PCyPZH0nv1ri7dZvG/x1etXQjuC37vt2GyBAAMONs+bDp6M
O7IiAqvG6MovizJZQby6Q5+8xHlHBwtv05HRVSSzKDBYcSIGHEEilBfcZqYMUSs4
jQPeaZakp7hB27TagnmuG0gqZft7A7MZO8fn4nFxi81V9AMGXOFV3ln+TcJcfFgc
acOUKdO9PNZO1HuEqM6IURFIuExfqlDGMOxHlO02HxlPVJat78phjT0DAqaK5DdM
MqrLPB+jSwd6ZNZ8Bepi9GHROkNk7OVtG++rFiT5CNY85Xf9bqDFsG/95Kphm5bh
0dIFMfjCwIXTQsT9tSD6T4Y80zY9cQ7irGGuwFU3g1Or50DGNziYUaO8aAJ4W8qJ
QQSt8HijTlEzKrn4W8p4GtOfNTrSxYzsWF7avrWTJmXf/2qx6hv8clf3gRDT9hWk
/DOinNcfzgoeoOV8NVQn3GEcKjSV3RQ9+mwO7VNs13pglzAXblGS7wRzKp6Vohb3
ae5WeayCZP/0lIPS0GlrNDtSoVTUIdk+X9tK3/LhG9DAODt5L64vZNFP7GCHM4lB
hj7RydVhJt3SVqzn6eJF7tfJxPrOK8+Z3PN80SNcfzLM1y1WgvwdgHrbTaR5VjjI
L3OgULiQ6xUlgTQ53soFSXvPCenrX1rO0oxpbYBnSeFyI4XCRixmn9AHqkzevuRR
qaRPpYyINYmW9Z0WK4BdIxu7jGt6rkcXWieJpmLagsx+bhRpTWiyAnA/mvSPy8aM
er62r3PtkKWPV0QKbsdcDpQdzslRm4vg0+5D+HTwYM8CntSUEKQSJKjT1j3bFnxC
Ft/o6ovG9ahznxhcQzA7nJNErDxt5bs9eRFxXlqpHlGBrHA8xKIpDokPVlmCu94m
xWGH3dQzXplny6meKS7GeknlwhrczpazB/Vjj7HnEFKxdK/noUm5R7R2Pn1LpRf5
WQmrAR1PYEiGOLCfTOySukaBOQSgfKzLjyztpOEBT7Z2ASrLZDNALnJlNapLxK2P
lXtExXy4wRRuR5axeb2lAb3xLCmdQNA1ZbsXRsRRn0xyD/6/LZZrJr8kvYwI1fZZ
wKcWK7Y8m5+R8OqYPjse5oRJIViNR2OKET2ax54+DHj8DPkZ01xs3h20td8WOCHE
q1LDBQqMZQenW+bkdtvGmMUKo4Jhij95+n24u8bBUTdt2SGxNz/nDw0FsSYV4be9
Nrr+srPBORkF70LYdCkth59lp+O80y9Wcrlpg/aEYbYtb46i9lWEGdvJCIBumDET
dZwBikNhl7jJ0MRcrgOy26ybHHJm14toP15BjAmQUUgXOYfN81u2f6Wv3YqyJzOa
TeTsepH0ulkVvObA7K+mtBVm+iBgkT65bI/QPJqv1kGWlP/A3HSohHxewdpi1GeT
bTp2pmK3uaQ6OJu5mxm/VVAvha8S818HqDj09Sc0I1RgLVsS8KdXvRbfcWlSyHYW
hdo8wJEpgJarGZuIG4kaW7fwFO80W/2h4w9q3ZzeqMsRnnoP19nSJYgxMSsIKDNB
7EsyNIkYaLSF9fSi4a5x3mO+uklT7NDRqKumoPI6JRCAWgTG42QQkXPZqLj6yyAE
7+5ESvK/6yecLbTcB81u1zNHbnFImGZ1Q3UNm+yBd7UyxJ8MfEza1703w3YAgsl7
IdI4LewnL5S0p+cI7kQggm+BwZL1ZYm0GUvvAYK+dWpBa0I6rWhsmOT8wEhOj3/2
Joa5FkYxd/IFyxNsf/BYuhfrRW+OA+1MMJsjgZBZBFDaG9rB0nyuZXqeGPRQvcJ6
uqaAj3aRdgSokG3GW2qHsZgkB/6IqILKIiKxdKPb+Yd4kqhPibm+9QUYPDO4awxr
buVIUiY+tfFOVXJ5HMl6jutUZHEJHvr2NEbSqX0oNiHurfNtlY6+TdIb063IO/SP
BPgEh0u61au2Cn1h9N8yoTD3/W+7t8y1mta6PGF1x5Lw3JVx165Van/CfFQLoRmZ
UzU2BLn5P6de/Pm0qpNxbi7zUqMjxtSBxAPQKkiXk7a8pi6C047k3exEx7+BshL7
e1iDmYmDRKPVgXfBAIo3gC4IS7GY+sc+zuyLUpjtkfq339YDVQi4d6Sq54Fb/7R0
fk2UgpJ1r7hSVujuNCeftAkLb8IAWlcuwioPLRd+4U3y+0WnJRCDtkgPpSiCend7
mP2smqpDWV7rnWZbgnJPUJGynE6Rs3BVTRrqYdSUr7uMEVwN/eskI9Plf4jVdrfL
gadbZ91pAs1ZM6wqZEjdAGBji5E5+ecCz+IXWB1eLnIEJoC0hQbm8dEdcDpuodqT
hMz18J30Gsg8vccwHmX9sq7LRBw79fya7C4IgdJmVWC5Xnsh9yFelSl428+VM5O4
n647Wp6EugbY2QIBlRNPGii1STnpjXdTWsnkUu+T8gmbaOAUw/acFf0Z5RDZQV1X
nLk5kVy6dA+PLFKCXscORaTa29Gbt6GGcKzH3didUhEbdxuDE6WBJaPKK3lTdmMN
/vxrO5qYRCHpWMC08BicxyXkLFNeb1dIn5V2LXPl1J17gmrxASxhvj/X/9JcgdOG
27frFkxk3H6aMxdgkRjfL2tyGMe5RGnr5m9vCpztpcm8kC2l4BmWTZ3VfcTwGIEB
PeGR3lunuoJU9nK+A/K65ro8FLqh0cRRGgIrWya9HEaaCVDGXwf0FXp5vQ3A8aFR
YyBmLve+z1i90+r35DlicEHGnsgGOkFSLzqVhJ7yx/VQEeDPP9OuzJZg8rMao2SC
uM16dRkoQF+CX0VNRlP9jcN5i3o1RZHrD2meDsJZWMFz0pT/2mE7rZFVq9IIWwGz
2Z0xCnl6b1O22/fLzFOtau2OfwGzzy4zwDfrE0NmtPFbFmQYJqEgKlKgCXYwOVmN
P3D7O97Hy5KOQsnIKa17rmHUM/24AP5DvppKPoTS9Z5ui67cR+3MF6tIlpUyIZMY
z/eSZQscjfM/zY31TV3lO1T3ZB4lGlPgkTqB47xWLI3EFB+3+nW7r93A1tWIppLJ
6f7smUc4XIDXDaKdrLw3ka1v6d7Ihwre+Pj0PuRj0QK552tUKPmegHK5K+gY4Y2R
IXyWdbdmMJPzXvb8qTJHo7NZWWZETokb7h4VKKM2mouvpyP6p3ys96w7+RkKtB5r
P9e6nmz8mEvsLr/db6+PwZW9/A9rv3uigMMeim7uSbuZVLKepTvKTV/hVa27ZKnB
OrT2gNMkdRVEGUTddKF1tUYZjp/tKnt6oBp94C+wRI4qboI92pri2IverhcbUpv+
RHOBryvLXbFI8sujP7esKNjpPV7ICSkL4SayZyRdkARuTO0YN9tqT+2eVLBmWxkJ
Ekj8qROAx6yn51ZtSd+XQ47QAoqeBDzip4vWPXx6mjMLXf5e/djXUPztf3f+adiw
pccMB1VJ5gd1NuuIjnFnGJHi5yr6ILmOcO984MFSJTV8Asv9USSr/t6+Oq6W3jq8
tXJBf+Um5x3McThmYcStabb6aF4en/TMi/BCu0i0yH7WTkBi6uwvl8yiX9dRxLfs
4W0GPH2A05gpxq5ONqpEOSimezLcjfc/bGX5MmsfKzGpmI37Y0KS3yRIhfoittU4
19TEfgyD4MZTxEBKeikop5iBLFhOf3ZuSxKTGcjq5a43SVGrCIuLXyehYK/tvI6F
ciH9RXnvSH74T7b2FgM3bFTbzOANAYbqGgKJoDRmZfH0fuXFsCvNuy8c+2AePGyW
hUwScvd22Ek3yDD/Tnk4MRlHOHJ1FSmwMZZaFd4eFpROmFtOk5LBIa3jiwdREX1Y
IjdtT6s3GdXcXqeKNmbQXIYSN6YmqktRy+fdpOPTmtZUOxdPdwxyOdtouT3Dsanl
iH+I0zgoQR7OvaK9Br3vSFWRFWucT7bdeLy6o0oSS4g8E7n54yWh171OwbyMk8zA
APmmBiNPzQW9s5YtcT61kIRNmAhbCGNSC9luNyqB2hzT8kVUJLRUCmUe05qC8tmJ
Et0g05BpN9uw6TROEx7y5xWLeKU4Y8QiGbJGnoX0U635qxy0IuB6UHpFeM32o7mp
HNfWAKPMMuvmDZfXtFACcgrLlaGQTUc9i0PE1Gb6GukHxbEaVsGHtswan+SQpDMP
52hrs1oojF1i3s/5T9EaFdVE+CnCu41tZxetgwhvkYl9B29aMxcCOuvc2BZA42nG
2Z3nvSfLvfqlc5IjPkth3wCd/hcnJSovjAR8xYrGMleRgKORtzjS8l1+qg2NIKC9
DUhGLOyvpp1Vp6dKRhMirrQVAlLJgtoUHBtQR1PkVJYxpEU6O9UngG2hhTvZBy3k
B/CdiJ9FZuMUmspNZ8m4DzfTkTaliOZ6ir6lBDzgAiCkvaMyRo/CaX02SsFVwerP
ovxw1r9D2B5RQmsbh8Ff42+q9oFHCCa81yZq/C/sZHCEDFECLaVcLpSev5f4W7rV
TbQmJ8Yf/D6Y8wlD2liqgg7DkQXNfXo4Mv/hLNWPfk+HErM/+pWSG+9caIUPCmkS
LRLG2QGYMupfA8xgRpxl1XA0LMzGlKzdTbl4EYLAJBI2Fh+8LF7wZXC4yeG9/7rc
2BUCDOA/W02JtQwseWmxr+5lIda16Tq5l26hs8GQu1E//ofH0hVGupI1coeiuwf1
JIAiCNcrrwHXOd7MAdtboRUnv8MzxM+4jiUWDy8etp1MOSgdROUhAzU2toSTNa6l
UcXUm9Sn2JmNfIGCYpF0jInpYfmOY97XQV22Lgh99gEMqWbJMd22ltY38+Oi7A+k
bxxaADvztLCDyL5BpqicPjCEC/Tgdo/nHTOaDAP5+X1DRN4zwH+GnKWJSya//RjP
Hhpct6lU2eVqBB5vdyy9U/evPJljin7MWMiJI1AWP/wVYPqjFziQAqsl9Nvs1Py+
tYzSwWe5yKg75IhhGB1XufPSqxB71kqZ7DeAuC8DyRAELuLKbFeS2g3OLIWJKzaF
tJoMqkjJqBbXsn+SKBPvtSffGzMM+FtVA5B3rf2WgI/oNviy9LnjsZk3zsmk20HD
lCz3r21pm2UVedcMsOmEsQAZLyGMSX/sg06QQkjd7SKEzhkJXMaOl1JvXU+2nFkN
btc8nPj2RP0jYVBS18M7597zTrNomJfh/CHsyr7mYPiOyDz2plarbE5A2pQ8vWJa
Nfc5gdctse3Gh70yfaop4AnkWRxIgEgnoGZGew8Escb4bVSrs4U08z5wEWXmPVZc
4GxYeHZzJiMyfbJUtcZeg28SY8HN0o4RSUEgjQPVEUr36r5h0vH0M3KcN6Orhs6+
hswmW3E2FspGS5Kls8SSW3sUrAdRTF2rD9X9UNby4zZIGR9HMXlLTJm6QlcSyoE2
G6omagV8WOCwDWpOYXbiI1iodTp6mZzJadbkJPntko7T9wUe2IKsOLL+whap685L
nECBZoModXM3/+t4s0IJFkLdY7BZGmxQeFgrm2+VLCrq5VrrregFSO05BzgwXhq/
Y4B69ILkNRbFJMlk2xdTi1+f5QmPIRWXX+YJRdvkQpj4ci5XT569gnuo+1N1IMk0
VByieSIUamwsiDvwil0IbS1Ns6D8WFf01rd+7u4V+mLr0ICaK3G6Q7pKif5pwAvK
w0Szzc4GxninQF6N2xvTenmlZmE5vC2dDsqwCDXadEjcriFnFZsiyIu0j2+A+ctT
zzV0xqZxPBPAsYIhic6qJtcNlw60j+9TDC/3YClzBwDFH/4fYx9KAICZ6VjyDJuq
CcGD5xEfYDPFqEGmGVUa2jjqbUnBmVnTf2k4AegUHSsH8oPY2w1P/Mj55O/1BtlV
8IlBUX5GiIImspwO8YD/1INSr6he5z/I+KVtrQq4Vrc5qzhWeFjTHpN6Kf70Fw3a
nSNSHdU87kuWwHB/+EYCeJaIehkspz9XBojNo+WFj+HppVSZQdE2AHlrlgipDGvG
J4LxKBG3iW2prW32hP8jjgcLJhXqdb8ErtqZiBlMDqYEworV/rXe954tWb7Y0cUj
bw7YWWHT/T2/Be+IIMJAq8GKm0POSCvx+qWV8GheUs1Tn2vBq8f5FSps/uVITUCO
Y4we7KEbgWbLPFWBd/RAK+i305QdZV1/bUA3ZvKFIpt4WNAVrxzKYZFLLbsBh/A7
HYB996ohw3h/dpo9u9TxoIvQKamsNRBjfTf3eSdv+6mtaX8HaO7fDsBO8yOvTxkl
Z12ir5P2KIW0rV0CdYArov6GtvDr8La/v6p3z4s0xYYwhOEtyffnaHJXJ5mZFPjV
X3qq7jpUxqUunBxpTtbn5eN/xvKBR/VZ9NZ3fkfbZD26M2VHbNVdXDdPCF0vqTiX
3KqdiEhrfzkq+K0LhCH5w1pC3/WnGNclaPrDGpWIovdUbxncpJny060z68xgbHNL
w+Ud4Tn5eH93yKqjWe1P/s2bIdyRj2/faFjEKCOL6BWQ2cZR9st/wqCCrjLcG751
x1BXDMKfx9XlIU1ygRE22eZFrWjIXQAkwqne9GditG7jD/P7piTG16Qxb7djvkH+
/k4CF/26lA9+A8uSMLiW4G4HxeB8VlPEEfK0NgqBlVSxsZnQBLcKhpPns5feUspo
9Rb1FUZdo0sgMzBX/2qpQVz0nNm4Xff9Q5TimWeayE4B2IOaGKtQB7ZAGfLasEHV
hWDYFJvGs2PcnRjknGbXC/2063JtsIP+piTvRk2617lD4ikS1p+Tm8JOfCUlIsoW
KTkh4UEVLT/TjEs4kUJOXZvEBAMjNS3tDw4T63F9Qh5GX8T1JEwIAIBn4Hwhd8qk
jj/947hd6DEdvmANYV64OCcDV2VR3Ci/UiQsuspJmNY3dnTzN+GoOX/JcYfbsjHd
QP+9o4rZYAA+zmzahQMYP/e53/vB0gDdPvwErQN2Hx/v/4rRpwUibveMFMxMyYMR
ijvOy8OvGOBAFmVLU4eExzj7RenZquJSPyalu/b7EaBtdhcTbJ1Avz5N4rUGhR7r
DBJjLJQNSbPFzihAMCiCE9PFV3Q+pcTZNC0FAUbGHzTVunmpGNmymGON0cRGWSv+
yoS4bzrrfU9YqiVAzLzmxIF+vkQd2+m5owcWbRkF4ox3aCunqFAcis8GkON00lK+
/ArSxcswfFoL4Jsv1UXoZ277tMU98Egd3s1A+WdIP15LmPJ1J4v3sj+Ew0L891oJ
Xyz5f3/Ajm3S0O6d1ig5MJTRGMfXR9SHS6zS0RzdpTm655k7t8X5gqNg2JEJH7sL
Ah2wwzx33T2MGwJICzkZxmygBrk1XEkTWxeBFUWfKWy8kxMpTM0eyQxR4AZ5Crjc
3NHrxb/6X9g3UhApErxKBH8PB8R01Bcz7ripwETfW31v6FGWC3d5GNhz2Shaw4L8
BvCmde+d27IXAkAp+e5WJhUpcZ4pRYBo+JUdktEbGQWXcYeV2vyz46JMx+gH3UeS
h7Qcr7rAgXD2/HrXP1EKfg+zpX68Za4PPrce9s5SmWvDWdVw5WFPNPxywGXs7v22
IMSM8/hMlhVAFzeb7o+Uiv8W+yRtqkIjdjr4ghY1de4ogO1zaVqE6rMwpFYc9Ln/
b1rHeMYjhFJNalNzzvNQ+BNos0am8+FK0bCHsTx+cB4Zln5A1H9VzU86J579hcad
uV6tA6iVKo5hmAwBfZxvAzm52amG5+06y6d8cp+dz2eq1HKE6M68I08i/w3zgd3K
8w3AhSt68NABWFwvnqUzfDssunQEKY9BPfkwkIL/Wvm4tsUtSitfVRI2RKrAQuKc
DfvuuiTZUboi/YR7Hb4X9Lfc5nZA05eEaO3k1PR6a3ZzaR1rBo46fNd3hvMBJI0b
Ou159MQ91/VZeD/m/IZX4si4jmjFHetoYhvC/P1i7Xw7D5uwYn2BgXulw0JMBMXJ
RXSFRt16Xb5DWpEqmNfiMvUc8djyBioEMQ/mOL026kUPVXSbRuMydV0xgj36exZI
3WXe18G6tFPL/rGoYFHtxQ5+6tUMJIKuDqKLyFcZ/aMsKKjs8p5OF2XAywGwLm+Q
8Qzq2/lqZx3BMDgT//1gitSYter8segwFUjxeXCvlN5nhArGY05gb16e4YKsVyVT
IrQNs2QhAU4/KMhNjRCwa7gp7jBAySQsqQTEutyErrxhn3WPdPy3NtmWQJAG5NPX
jjNJhF6WQST7i4BOuTM5apsPgVv15SIO46AaHTL7URwe4c5NHSSsp58LhE7jCv3J
0D7+UL0x+F85ocZE27zqrURA/MBcthF+cBodHBCwCIVc07i1Vm90b+yv9ZTBKp1D
fKHNR8XJVL7c7jN5RvnVoNWu/jFKDs62QMwVo1jUgb9yt5muDLqSUM+O0DTWMw8d
KSOGp+dBdUATa01bjLVAQe8E1UNBiPk0lvSXhyuxqEMrL4hRmkpIPPexthhs5kh/
3TGCAz6/JT+plkzd+Cg4yt/gqZ0Ugv3JUw9vvLAVvjhRthU5JMZR0z2YlsTyeMSA
sEBMOQQwUveq4i8k6FXG4iwXuLrQpEyZHtgnNJ6f+QyYLpla54iA1O32/7RVCV2v
ApK5L7127ikyBd/Cec2uPPnLWIfVCPzN7Li1EyoVK/1Btx5lCD2IEuEBDCgfytxm
1t4m8S1xJ1CHtq5lJOzU6KeXT3eo6vgY4nU9Fw/ny2CYQQN6hxDPg6mgtQgB3oMF
QLfgQT/bFhBaTzIu8VrAIPMfnv9FH75fQH3VwSB7nfvJVRFvcEBDinmjNgMHeFGT
HREetX0onKX2c13cm1iKwaxaF+Dd8oPrVcSlfPTD8oP2p35tBcJT+9wjOSRqMrTu
MJkha3dkINoxcFtr+rJ0Wc8p2l1V+FJxZR6r19XLxosKtwje1WXaptvuickw2f1e
c1CCk4F3956BEsRtnIiwjHOgNhAPF7ngXTefw159VmNw3TwQeN31eutaBAljVZOy
OM57GydWa0xwO6Hx1AvLmA3Z4ps7z5EEZhf0bnhm1AXXqAA9mir49ZZbywHqfNJS
YyLE9CRrvGlfjf1S5wK68p+exApSWYdmLiIIZoegwf2V6/lUBfZot5TQLSA8pj3Z
cYmQbGUIdRUttfOO6AXGkQ7hEcyqbXKNjI6HWsHCVDJghlsRzDa38lEjr0omA8EQ
5/k04SGJ7YBN3O0AuWNHazvo7R8tFS8wm0KL+XIM0zmtY9grRY0sKaDn0Lp28hpo
ZorUmJ/yMRGZqXmN+Xwo/6Q0JUW0x9A3JXApFPBoesGo7t2b+k1QAWaESE0097E8
4Q25uALSF133BWpBANpl3N/x7Ng0AXO707WtkyBsFVg9fSWcvD3CpLryKbLF3orJ
Sr61BCkiAoUfl7nC9yxWvnYxShyvr8pArrz9qecQ02HGyukSuctYT/4poIh5a83A
+dFSqX2XL6ijlyd5u/GBdcNRy4rJwy7Rv6PSWreq+cXGfuP/BjsaPvxF82p1U4fb
2H7pyhEb9u5Q36Y2Hi60OaxB1QPfZu9njEOjf0CHmZxOjyFryYJi7jD437YovDNI
dJsiulkQERHwlUUKPLSj5WiAvVtyX1ZgjQEZsh03D7MUozAlaAWKLMkxx65jMz+b
YWgibmH2ATCM7My+n+Lo0Le+bU9gQpPkl0gTyBvLmw/3SLYsrTsabOdBsMcdj++T
De41aaYdk8C3I51V0HHw72FrH4MxtTNRS30ctkRb9ri+lVaA3wkRRGNcz0RJfvBc
+NTHfeNIQZunQlBuP3CgeHojRk0UoQgvTjMU6p5T8YNSFky9q8MHZPtnYHr3P1sY
XX3AFwkyLkWdZuubnxu0L4K6WsAWSr3GMadTDUOUbfOUtMieMBp/ZRPT1sG6DiPl
WrTWRM4fRxw7e5r+7MR2R6gM01hTBR2wVT9EDwVgJUSp16TUDJlY2FZGrFN8fpQJ
6sd/uIuHqktEwD3xniDKMNFl2E4B1O6b3IWvoPawBCUMa2dMtJH6z8F94D/R2uv9
g1dt2mgg8od17+xmcGRPQg8D04Az6ChYTx7UMxa0vBUPu4rVMgo7nk1lYwK6wiLR
d1dgmFOfRaUHlYTbxoYMePP7CQUN6tKLZggVtdI/f10ruTHCXA2SjgNAVnM0j0Ps
4UsZ6NG1BxQSbs3nWH5FEwsoMKx3to1W1l4eF6RK9c7+GeDC0PaWYlWVspeHDVfI
41Ul0xxFB3Pxl1vQ1/VABua83IC4RjU8Fpt8f1c9zL6/mQZVTeRbRBMQNXHVNAti
051sZnN6RyK09B/KjkjNzZKqm1LhNGoT6P6EZdLNl1PTzo/pa/ZPc7E5MI4+8iyf
lXwgJTLFAnRtrxErDkJe76SvJOtpR7eAgMwRWnQEY9FKZg9iSZwcruZsW9H/nQmt
9CQ6izPWHeeVYVIvDAifgXKRfzh4xOui9R3LUSlqPgpilAVK6V5DhmxA0exYEM+n
fUwj1Fw/JniU3iYOMRrtAe0CpHr7QEXwOv9GdXfoooIIq7DA5Or1fcnEizBtZdL9
60LNRcw3NfQo/ClM2KrWF48gYZlX5EqwR0KAuH4GczWjZsQZdGv5UfYCrSqQaAf/
dyJvJCITPE0Gi21zmmY0yiR3pE9jnML39vJjypokEzcwTKQ0qzBGi7vXyb9YD0OD
P4bDP4l2NqF+bYZbc7kvztptG/8Nse4hVYzbqY6jvcgvd4cIsHNDO1QDroaO1zoY
bdt/IdBetglIN63yGz1QPOU43CjQK8MR9BIQn9hh1GFN9sbq+qCWfTaJG1Kh+Jsj
0RCPz0nNenYDx0WONZWF2bkj0+ylW4Hh8lNsN2oNEEQseuF5Oa2cYjCw8u9Z/AZp
PU7Xr0Pr+Iroep6VjIMlPorHLzL/k8jrBZgZd6HhxoFQ0KAf/tRlT9uP57sIU+nE
tpNvgZRRleVQYQEB+FVIdZaak4Dy7oYpObOT5BvySL//hoPgmYQaov8zvCTVGFwt
w+3ifeBtCYbzl7T9YuZD1pOY6Fxa30KEvom41qTtjMaOyQ/N8yy+Na/aNtJn47Sx
gxN9aBhAETGg96thfMcvsJ3JJD7MNDjfYlD4lwb5P4GW2pR5dhpKpl1pOYwqwhZM
3slXj5f0lof2SkNYIATTv91qSdHhWHzdzPhNcNUHmPGQQwI8nokRmAafeAAakI3k
FN4vjZhdyd6fTZ9uImYrLRDfwt8ewdthetYpnxUAIPfAaCscSfQx20zk9/KB8eBO
gCL/fa7Q6kRKotcBQy+T9XXcOLiakSy7UiL77zFCg9s+URlOOJZGBcGcoucfHWKA
Z290l1IvyNJonvOjXzPPSLXnq27jCHrCsGl9g40AO/dSCg8OyuGo4CKj2+rmojtf
FL+TX0Mql0xC20uuDHWL3DMQGbCcS5+Axn/t2Lif8MZdR6K+PnTFW0mIQZgtgNWT
/qGxY9fILBN5G7GepfgClv11VXJwZkLJyYzqfnCrhHJrJqUbp3oiuwpM8wNNlxWA
JklTj6lywqMbYtPeYmSDmW+0p9ZPFjeawHIK85JwaP+sy57QocDNMEf8KtSnZoYP
23BDx3u0wN8quRE7XSsKhJ8DZp2Zij5cFMvENrEpJh8JBF81zw9bs9fabMx/+kzp
Sq5K1MymEsnqz4UbVfiSBq57CqOcH9XJForN0pRYBahiw/EQs8h2CpIXRGKNo4f3
QXD75ggvnXXGFnvhaKCBzq8PM3tACjGKiyg2FQrnhey7EhORaPgKwoCjSW0IWgl6
1vnRo7nIKXukf82TVWzi2fhLTRDDow+86c5i4Pt1IKOLtN5OrVm8ztBbF8Vm0oWt
ZFHS8ermnRqNlLaWJRGVq5zCgIWkEbOIlY8J6ZAc3D7eiaEX3k7rTv8/W53ERXdt
ZQhOObKrxkrnySh6ticDcNrg8ASzdFRBTARyFYWGlcXIcAXVFsA6jjkd23+OgccB
tiy3rb6CGjpuQqzsdbtItLET/aT7UPZ58Q1wlpkaOtSoJfsGE+wmvWRn8izIK7yR
MTK//qI11snyFJRIyAzXoupcC+oTVDMFZtWPhVKESoyU/rpQz4Vr6ef5mDoTUFlh
cUOsJhu5ylaef81ZU3DuMRl8S3aVRqdHa6r8jOAHJND/cjMmWAyLsXdH9lmkOPfH
fRCTFkF2XPCqVh0eAep+8jKXW4tHw78kM3isF1xCbB8UfXCU5N7wZzlbBOUHto9W
d47FXAeiVYFxZZ1y0Iwlxc5z/BlY32Md8V+urOSJsK62GJGsM7ASZ2u+ZCWYIbgB
N2RtPwKOmfEdG2jIiHPoO27Eu4F+6lBrj+8NBXNN6BCPUJBZxmYTd00t5AhWtWAN
DSbdbo0wj0lOM30S83tN8mm1FRYuD1d/7NY+NgBr7yz9e3XjCHxSQp561jgca0RR
+1wNhCHfKbSYzaOj3ypm996/iUx+qul4L+kOmNmY+Mw+UcoKic8RtzW3zmp7+Q/Y
zKZZniEJ3BMp6ZHN1cnqbCCWaqw4m2pfLV/5CtGx74VmUm01DvXihB6fhqKNhP0k
OrjVSEisxfuXdeX+litXe//H4iJ8DsBx0SZaYhw/JI8ahE4nKyFC9Q3wr8clayv1
jGq1dV3R5tgtXFKcmEGtiAqZPnR5Nvec7GpIiM+7pFBvQxtxM8+WfFnSCrBCo2/f
anjmNkiAdfhSMvCGOKPPlvjCBUDvWjYZLDdf1wYe73yrZjdRa6AuO6hT5I7U/iCa
Bz5oLlyO3rCgyCpNNEU7jmPS3j3cgKVe6OcAtlMq7Yexg0iVOMgcK0m8cd1BxRnu
VAjDlxioWKczLN16uqXaS9idh8FFp+iRYLgjBGHKobZIIxbmLmx/EReYzQ5GG9UF
96d7syorSs53ZULW+KJtDSoIncFB/Vb9QC4Xq8qTHZkGeVrXZLFVES1Yy25wp8wT
qQ+c3oTG4n57cJVj5uVTC6uTpuIqrO36FLVdQfqTxQAyAjfKSvHg/1kbJph8WPg9
Ma/e3G+KCyGPyhSFv7ivJ0mjHLbETsIdjoXVhEXXVyTcG/hbAUbY4E/en6SHSFBN
gpZHFNsEBDKvaRyN/gKPHK+6yviwFBbmZBpmnKwk1cgXQupih90pYANd1C0Plicq
0W+r2mjaXHWypYbpfeowA4JXPIatuniQN1Y1ZEmBhB/vLqSMD3rkV5QEtxo+5TyR
aOnJ51seaidpXaWP5rBvMyEcqMiKXyjUfSi3v8kHogzGs/QHFEC5+dVvKvL1zVr4
i/5XdgMJhuGAZTGUSHqQWwifqHED1dB5r/1hZ8EuCoCjDndpxwqG0cePyd261t3h
Jn632WnHnXg4GEyGVlhxsU9J++NJi1EM/DStequtxm9wLuocp587XiUloRWmR34s
fkGwCSjac0zM3GHckCv86BmKxkH6lgqgK828RXwGXzJ9Yf2i3THPO1oVreZSdEGt
RZUwPdOFafb6HSkNFS2yVnTGjyqFvlcc8/glu1joC4DDIMWIfoHKDkXZvuriAWxZ
s53GLdaRKS9tVRbRMLHox7tffBWl6frFPTb1ziMQTSo2Nc45M2liaeyLGh5+xixN
E0BYfCwQFwfwzIHcFozkPlmcs4JCuJCXP7I8YeQztQxocHbkquoA/iIKGQPvMh0z
4eit/PbsbKOSpZ8Nx0U4vR8JQe/E+/nTYwJfdnZeqHYPhGOchf7smuTiOBwL+PIL
59FthozuMJ0QpweeIYTfDEDxaI5IIogEk6rCRfDzGj2r4qq8B0FKk/Y8arJELIi0
BNRimTp/Xz0I6VFKyC8td13eyVzZrR3VwGYrEAEzwMPPOvlld1vexdoAyh2OXewN
pIcDshHgEzEEvfAwgU/G1OfD3ZL19LSEatLGhqAqA/GP9s7TgEf40hnuunNvhTXm
wMH0226PlvJHyzy7Pmb3ijxgCaU41Y/fTB5DfWXc6YnF4JXVpVRk/oHlLz+JQRs5
PgKZ3660btJaLxI3g9EEfdLwHBBFC43/RJX7q6bhwhJ4ZqVpzfsGRNWmcHNS9jPq
MGiBYNHyRowAHpHBs4ELJk5C72+LfxhsAFj8KNuEalzDWGzLCTYMb7FXJezIJAeY
mNxlDX7gC2Z0C/bWXMzwp9Nl+y+URY4jJrJNjnpEYzvGRV/cwlqC2xwSj2eZpos7
BdyjP27BOfEcUw2VmJD9acbZmmwhAwsxIHEFKWSISGwhutlY4d87hy/+eii4Rfy+
9hhC5eSvaj7YAcPEJI61cgGxcKCs7CWp7NuQy+jvpwWncfkgNrHc+1Xrx61vbhTf
KqyGNHru50/Cw95Mause+JLncny2g2ruLBAiMzLCUC+EprhNWvBpci4XOsD67zqt
vV/9bfOeHfyzkQ3rvtJfGML1tb8ZBC3BUHYyWnYdpZaB03dETmNYg3No7AvMzPNZ
3YBtVIvfp9pku/DgJt0Kt6Xxml2SkA8LYG7YUqzlwK/SaSR5321A23HjC4cHBz0Y
HYS4qvRwuvRofWtPcssikX8nkELFcV9XHsAVu3cVrcRF7Ad4xK0WL3FD4Fw/PEXJ
ETCjCjOCE1VS4emBDsMblhe0OyNkWFGfFwfov+QNWCm1AotokHvtqGMSJtQCEIYF
fI20w1jdsjDI/06WU43UVzPHLYZR1/bBMKJJq/fCn0mOj0WSOgnfd/vXjGLHGFWq
jFfnH7gyMYXxln5psO9tXC4SHXCkiJezQENmCo6B1AVeHQpJPdV75Ijm/NwelvxN
Hb1KBkDUBIMcQzcuSjlWxTjAv1ClNVYN+yFlYb2nM49vj+AbvPn849lHBH/yE5uX
5bGoBvvc3r4xrmC7HOPy39gEH6kD+exXdgzj8/l8CH8TTDMb3gv2MtRunI6TPfm6
M/kMrCma+DFlB96gtsMgAUriEWroF1sdlkR727/6oxc2vQYQxu88+39L1eBxe9Js
O6tMKLqw4rRxcU/DpaoyLM1vw9oOqy7959prTPtEXabz8F5ae89o0QtzuEKePszW
ItOliSqbhqBO8/QbNFt/pNJmrS18BQ+iTWaaencywW/1FMZcKALHkKdvTSUdeosG
NgUOr06PxnJYQO0ZTW2sX0+xdDAfFRplq0R7yiCyGXTybv6hFwheCQ5N5lmY8Ofs
29cZ3WpUSZa7UvlCdnD1ouQ+krtDCztCOwQuAYVd70ARwl93NHlYC22j1Oq7Z9Td
OKXJ2sahqkmKW9EE1vQe4ZqlL1S3TkKG4p16qheC7lL/hwDIwtrhQ5D1F99zAvQF
TJYMa1VMQekV2pFn23jVhHjxTgAz6S2A2q44W5Zju578Vn9kNDyTSpTKafAYFRY+
34U2nS1tHpsdOtSlRQKYyXr9D5BvvNDD0/MAKoeCAQiR6dlfNwn2ie15QSzmXcId
FLpKhsc/BroXPA9gyPjWI/TACfc/lJGj2styFF+qlDta5Sq6KCZf9IT57Ffn/mRP
81yRvrrzFr+/0AwUyrL6oKZ6BhuOHmXfrWL0x1b62zrIo3TvI2wYoW8+snE8Slb1
bQ+aePjW8p23KfS9LsuzGlNJvXnQMLkUgGyEhDbsXvULV/Hnt43Ohn32mhC5dz4n
yLn2+LBvv39XGK3OSvz7Ap2v/pPx24nDSA9Tke1m2DnZbvQewEqm1KniNC42n1en
2ujM/P3RkE8Kvp1GTs75ZHgX/5MYe6WDzLL7o2feO65IORTEPCIr1qPcXCBr7Z2B
JO7KYlduWxia5r/PGJJ+Fxt3Si0zIPMo0u9nlYrWaWQouCX2i9iRlDxQwIBEacc9
NlxHJNjarPapu1st+ruKcaSBdeuMeho+yDIdSQxb025f3zClgVsy3HmBxAlH0dFC
GjnZeu1IT2jPt0YS/hcbkKD0K4bWeKyR0MUmGM2q7PTao5RzWCtuvtFvcZoXGcjy
lckMGoCCaf8Gvox32Im0gpF9EHn5UrxXkt9MIvTuftqivTF9JEYQsTHNtpaOsa4c
GOwYTKto3RjYADqSZbdYHANANqbTvC3g8a+2xRCREDW6L76sFNqZKwogpV45no+w
V6M3Ll6NZbBiRRgpZriT9mCVHJxWPAd56+x0BZret5daMexlws9FnvZn6dAQXw5h
soa7UYhdqZ11yMWvr0RIl2STbFHmPH89nB0JV9Y9GSDBH0PBFIBOHCECqDp85bzy
DEd0VR/DelTx4l5GDw+gBgZk+YCCv4EB3w9P5Y2jAQDbuX/zOaoAqcGrtZykY8HH
y71BSV+3pB2VvCDcGjMpk2FjP4lmiBUJDrp59li6RY18QlN9w9lcMe4pWnG8hasm
FOlyr+erg2G9WmpAJBoVDxucfmTD2PQqapp4S00APUvzopHVL9cpTnuahoADdt0a
gv11Enb8uojvFQlLvyLquKIASK81gRP2PXoBpgxHS4x11LjlRUqppyPUyNytXDf9
4o8LhFCfW4vYZ0WXHhvZAwwoqehXyALUOKDKcBWUjuT/e6w0DJA3ZNbTEPR8KPqI
6vOHV2YBTgCBMjTpk7WxNHtn0ZWGZaQ5D5skIPgDd4EhEwsr8wD0otfJfek4yXKX
pVEF6inygjDjc83O6DHXVOupVcr3jnhYwWnAsaMA5Srel7wKfXpkWQZkN/j0IwIZ
0gEGuN/wBpQC9Q1zTFSTXs6dPGVl51X9GmvusoTkZyIhytHzgpn22GKhnY51cj37
JPgeWK79aRPH7zkTNWtwYUvD0/fqdeK6Xtxs9/XvnN6nyL8816ga1XrT0CCJw2aB
sYCxPdUGpsmoIVCxc1HBKm5EHPfPMARGv2eFaH9EDuXNMXkHlZy5QpPmifbh5jlB
sji3H5TXu9crS06KMTLyOcC3cPDOAlsoKWfAKzf+TsIzpuzUug3tm9yWOqdtMuSU
8cJWPMfFNcVvEAKiA09z2P2Pdu6ffll3koR8uIIJLdhCM6zHa6iKQAM7j3SJPYSE
h67rl1o5XGX/ec2E6F+cbidtcDPcBiqvgg1AELXGooybVgBjvJlPwiode9lzKk3l
0k9ndcm0pmD+a+rN18A/gl5Gbb8WGo6cGqSJP/VrSO5+vJ/bqoL3/d/00IX5vaMi
G9mBB4CJBJtR5MlVLLdrlT97yG+8K59JfNxj/DPIXNniRxCbHEL/buqzncGdgQ3/
v1Sv8lAtO7obxm9+prS4ImArhJaSd8FACQd/TqFBM7kpjrk79Ae40j2gziCxysuk
mX4n+lUpb9BzbXMbVj92qOckX5RenTkzIgfJ9aDFTnhwcm9rf1kNHxuy2RHLS/QO
/aTY4WRKOFk/B1tFVF0sOTakHtpszW7Hsa/KQ6TbsEutLmCWTCCaZwRV2mAnO93a
6LEg2NTr6mOQv4HqhTMFmb00LS4elPpTrWYw6mfGNHf20XMjP9gOYMpPvCLvlKAn
N1y1lKuQvy0Tvg7wFmQGTPJLoraQ31hDIpZsvrujrEJEVfqoIylnak0FfbICcuAC
4HMQhL1Mx7U4VC0M1vLMg2RUJGouhfGRD0I/1Cp9VcQG/Dx+hICpWuqPuPpE15X5
d4pN5EEPssyne/Ey3hKhvTOEa2/dhCsEzzotp+Ehq6oquvoZowiIgWBRs4fbLBA2
Cp9tjnWqkUb6x0waYVCBWuQ9z8yRdE3e1VhYITpgxIPfBBqOzsSxyvQln4ItZ6VD
+sdNXJwdnMqve63l44Hj+UrMI9vpSZXhP34GcNULI0o7C79Ak2SX8IKEOw+tKLGW
NL319R/P/4OsmA84LYZIVT9mE0tCZP9JYDk+juZW292HSVByQktGVx1kc4NJUaVK
YP7bEFLdzqL79MDcwXDncibSilnEx5Sk0xwp57WOnPM5ycI2bCDtVTxsble9z7B1
smsRW1i7XkAaIPYunNsy7owHt7RhcycpAOQ7//ehRJcAKDz9FsMa4FJxh4X6ApxL
8ZsLdX7t/2NKwhSwcTRZLJY7uz1XqZ2iKutTqCzavBLFjaCQIc5pZvj7TDYH3Ble
iqZRcH6wqjJZG5bbZAzgZGiZxNEd3a0xCxQcm1FQcf0LfykDh5l8Z3C7ZVtcwNb8
/kw0bO6XqqmdB5y9PVXyl9xSjV/q1vOOB2h7WY1CT5mkUT3PpvuNNZEw1KzuMi+p
1ZKY8PiPKhiDjE2RjKWmIYF4cm8DzLi/jRiUWNDkn635l0RLHjts0Jq5vNyJpshJ
Q28MD42ejyk4J54cgHPaxzyyo+j9nVILPAZOOL1VQk8WjULLeMQ9Fm7PZdeZ0Rwg
PgjaBDy1E9tEuYwzpXMvmZELQu0zpxPxJKKbdo3TyVu1IqZ7oVnYpAYZKY8qrWNK
F+0yv6yVRTBCJQMuXCI9r0tfLvUN+QvOj7yMxSh8eaaI5uNvu92z1En8xQHSE3kr
2n2PXwUIfBTBZ/H1DXasK7kIcDOkCLSU8S2/FFDy2VEzaADXQENEznPJv4Kb8TI5
/IbvlrrNWTGc74L9Ma/RbYiqsxa6EFVOuTWfwh5wjYahPrPN6RC+jTn6/KEmR643
J+4wXCTsnnUtnlfgp3s8UPbu8s+faPPOy/kbcUcjKwH9rbZt+QtfpnFNq73L9jKF
8lzMcfoGwiRgJdDF2UPHUTY58/5iSE33W+0bq0f0dVNh6IYKpNBojsm/ywT5bMYK
l5Tl8KzmM2cRyw0XTgQxlwYt2MIha/jlf/2kk2KtyCOZqKt1JJ8N3h61d/75lCEt
IOYFSqLFTclIdKqdoRCXzEKw8M328ytQiIRLg+CI8SnDWq+kFfxTFN+jDu2h+ZPd
1S1A0wDYvoCluQXbYELYRjm9k8f5FDJ20Ok5VYtRUzZGBsPTnFmK02TkzkFBedhx
gX+ayJskdBuapazvSdcNgIM01EjhFtpkHLRQ4x+6t7dgDJL9MOqDXuloGoPzerXN
sES+/+67LHH2iWa9cm4PnVgLETOmbHv+xXSTeeNE+NFvqkzJok3/485XeeI7zE9j
FNfTGXDfO/Siq0ttrybm2x9pbaRM1zaIRym6UVHQZHBc1nhh8RgnmLYWAAc9dVxz
U5YVgadTh0+hwCFh3bC73kchCc40WcAJ2fZ4vmDn4JL25QYkA6FrRxGyp+wXPyPS
mPm6/4cQ+HnwhxGhSTg9pZPGfLJ0Kt/db7yOesmZIsnUYX4rE00L68XPSKxpa/hy
ZN9mxP+GmTzpwCxbcCqKahPBZd8gyDuXWGZ1jehHtOv/EHQsaNB5A/3pOGxFa2xL
veBwO12jmp4B7KbToOqYCDMuBvUWSf08V5/9SCsg1J1BTf3Xk/KUQxDhGjZEEqST
LgQebny6j9nONMpUiZNq4VJChPV9MSLwndmj+GKaDaUYSj8R/BSyHnUgVguLK5bq
QcrN7J6LVFl/SJBOv2+XVqm4zgWL1PCS2juQKVUD2SgvubAeHCZIq8J3CuJ0fwto
Nk/Eoq6/zPFxzX/+ftfTjJ0+OUDd2kQYyHFMVfjQFHVc1b7FqOuOiWbSOOSXpq8j
Ady1smvdhAOm7bqM44ImhkYxPgQ6Xb25kQSK07O+9ByTV+CJCfU4Ij/Og3tEKljy
G4ZyDV4CkfyoaIGvR3YsP8W/on4KhIrxor89IzFhcIBDcdhmbqc5qg5L2iUi/65j
bu6gM0q8anrX9yEos2rqkZwHp+ppVz0wsqQbbmTJIZjZlOKSpS8DQdYbgAtK140D
2lnogfP7n5UNqCuVkltnpVsLscsuzyTg5eGbS1WdetMDXxs83/zfmmtuYWfmtgAZ
Wn6ftWMuDFTIdD9bY/yV4Ze+2fqWrju/KwTP5zzzjEKNmjLgE4p9X7juztVMWyjB
fiVcv8a2jOZT/OA512TZm38SB9SP1ei4oZeNTxfVzgGocZyzv6gNG/Fsr6oHPTEg
yJvIUZc3B70QJvLyFMlzl60B8QPFQuwsi5qhZ/WI273b0vBEM44oi+wD26T0eamp
jVW6OJkQTCpYVVN3NdzYoWqK0UDOt5bSUcz05GUkJUA5KGFVKJroN1l7e4EVx5LL
VMXEk4SklCGrUlFg6GqS1KiKLxZOKDg/y7jaSScUEFn5HgfGDIzm7WRxE71nPqjB
F0BzZpGfBRdGimr1503ZaTmTKiKkZSH4na3fEpXdfDsZ1YrLsTi9GiY/iziPj4rV
Li7AeILXWej57F5WOzw+aYeo+Jc0hu4fIioUoQI+E5Hiv0U9Xx46zSXcfk+snluI
geryS+3fFGi1l5AoFdIUTqwtQp9hw8Qg1L1aCyVDMuKnuLvFs1OZCvwjvjAwoa+Q
f1zxzXbSzdBPhPlUUKuCkAvCzq3Ub1B139AfzSxZ4wp526H63szfGOqDJpBw3xIF
INwAYr2YkaXq7SAbphTkktQcQzhd/V+35OdAT/YGGsxxy9Cb9SjT+4l6SmnBjMIt
7lgooy5lzweTPSkdkR54os58pWwyfopuiVYEX24RjS0/0mqENGoPPcXv4Z5SqGbU
lHemcrk9+xgs3if8QgJ+5erZFnuwTHcM3jqNGvzdjw/+xxN1PW6kXeQbCsin4ISY
n06igkSKggcIf2o5bSqbWtiJsCozedhb2d0kuCwHWkZXPDLKaVS+R4sXh0JNbPbk
KKHFX8zBko7wDiTK2WWF924Rb/k6RLtJ8/PQ30foklZhRQ9VijnHILJCx5tZsmzD
LO/b/xtJ4eAA1JcUvTVjYsgnzrwpVF+95Fa3CAkwTqgitXAf0FojS5MFfxHsvr5h
dYXi4OCPCT4wRJTlEOV60ehkAo1T9JEMb8gqMF+0Jz6bsaZ90gPe/S6/qWgMiBXV
41jLU1oiSOgu36C/x51BarbYPQO/92C9SeBrOkDMpUd5DqiEq+GyufGsvSNP45g0
MumiAIe8UNvijf5NIxn1mP1tPJjVyqAkj5Q9LPdqEsdscE/+Xp6tXlGGzC+r2stA
3DEmqsmRsBktu+/y7zp2VE8TH+gOudWj3Ijw/t8+ZVqJoOWG+P9k1UW8LoIDmT4O
qlwnqznPkjT43HS/uxTcT53yk8yzxS1OjwB996AzDm2tG0xuNqxlT35BqSEjiE7K
nyFWatFli4HKbbmh8Jq3tYZoeOir6EmtEP0QBLmWQsZFjxdSZFUw2lKj65OVyR2E
4C+l0+9qlahYgiaqSZp1Qt49t5QwO6aYnrBrfeXeX+h3T1SOaMuNIwd7a4tySt9v
F74ltJbXxaoq+LnGdM/O47SZf1QVQ0FSMUIik4ax3mrDJu7fBgbls4k2p7E+gsED
vsXSsLCXpq1LhAVesLdFwlkd/GWbpGEZZg7dpajmjxvKDD7re1ePJHHhRI5qQH31
3ndFGp7uE4/1nvKC8AfYeK3Haum88zuuHMdluYur69tEPBOkwecxzrnEgF9wZ3mk
GeOKRchj/i2hbLkay11/WD2C060dc47bjHbW6ZJHPzctiVAZx4gpI2HdsUo3r9NE
3M4+qEBePSx5zjSnYlA+ulwem+/EWmgxQMnrbyWY41e7ScmPvwfHFNkN3gtoerg8
sFbnNt8LAGSlU5cy3c2Nv2xblx9cWBDD3fTCxQFZvmTXLDq8e20v8rzGW1kCVzGs
i6UuTw7XRdjcwl8NFWQNWbfsvGQ8VdbkR4L6IZFS1q+Pc15R825cFjxOtxuWnsTQ
kMEC3tiXEWNN4CwMJfVZC95eAZUtOOdG5IS9s6VrCQXspd+EAMKcrc+2ULfehQLY
F+Oc4DswI1MmZSww598Vi+nd7yE34C+QGmO+SflroCsYFwf1ZtdJDHwsU/kjgaO4
lpYFgD/QevMjECcBbs94CSe8ssbnYWhi6SP2/RCxr2t6rFJyVmPZ7PyLmBbsJZfM
N8cKiW7+mZyz4c7D7duze8pvRS5xRNj/+w7MsEPCnu1PshNjs73RSrNCHhfZ32jR
IWoXoGVyc7YyI0AWnuPgdjRRvh+wQm94jwmtqtshxV6lsWbZZWSjny1p8EWDs1PU
F6ykvOrjCNOgBbr9kpJAJFBAZIRdvQ6J1FmUwrScKqer4i9zNrowzBKsIbVPrTvR
+pecGv/weiJL7LsfyOkHs2IN60J9QuyJaM1EoTdcpInSPBAMDAZsh2uU/wbMqjer
+qRglbBzRTRuvUoQBSOSqtPWFPf0ooyqKm3kn7P8TxpXOKJZv4OmoV+aIDizJoSA
i4gZu3vbU1LN1+ewmIYNQ6SWVyi65xXFrWv2UYKrDhT7Yr04pbYk+kO4ciShcHEl
/Nh3gYmW04j0wjv/hSsId6KGBxESDC4E/xxSoQCTrhQhr+aoxTLYzhIyyCu4oQmv
Bou7eDaKmy/uJQKlnHlf6brxOxa00V7x4wiE4eovlRLYb3jMSNaWH06fuENlX0yC
ElqRsIPyBtyp8XIHZLcqWba/8kBx+Zb/yZ/vyoEq2VYYqdgX5F6X1KSuCKas/UJH
U7f3n5xxBmIILo16d+YzXoAG5L2NVgSYltL+U0vmY8bEqU4sT+Aa2lEYKgNeHrPu
WI1F1fZL+iNRMI3LjnbCSGoyGJtmbSUJu2iALrCPsQ7FluEPfimfsbi96jUPzzEL
TiW19SdTIOkltQ0DdMPaAOJ///QPaw8UOyAdcqJ09TZ5ihElkuAt+OH+OVK+D99m
0pCA6dTOM+UCU9FEHWtR2HCBZZKz0HX7iNzYg1OGd5n6wUpktcx62F8e1tts5KcS
8Mfk1zXE9b8lt6ujKdMIbcHTeK0gnscgMBU8KmWBqScrfkSZc+9+sq+6kLyVA7wN
XomrJwQoDoryUkWfcNvBfbbMbh79b6HpOl1fkn16vyK2lrgmVCpFD0/W+JeKGfAM
Q4QZWvQi9GXAWBxAAjc3nSXMtWDSFQeHajFthP/ye8u1UFl2iv6r8SVeoGMqDXng
AOEXScH83IpR81s1s5CmB1eshKdCXpzQyVGlZt9L6hyZOa9TxpuHoQqdyQw7VucO
035mnfngQq3f3q2pumEaWZDD0oybeSBcWB8wKPgRajU3f8Y7JhFbyoLy7BOM8035
1mdLdRYw5i7l0/skoUH9jHYoZKFmUI/8NjiwS4pwbFUn8IbjsbMV6LSeMzDvJuoj
HMYXSKLkL2bLSuPyS7wpkj7bCR9X0gTt/knUjJ5pATjqQ/HUlRKLsCLDYXcuj04D
JuGsbxp33TLq5dvRQjt11kWXk6wAxouLBlfih7hZU4jjzqo3AK9PjeOSlxDzoZEq
QzdjAq6rn5IkcWn4mDjpP5NF6eSIPDg1MNvBERV3I1ZzUHmJUgpjP/G40mQo0cKv
ZrCLKph9OFqflaJYpeEut0V7jKRHL3gf5w7kI9NRag7cLSyUwKRw/tzsBEElI+Gf
UQcvM4+8cOsEIxIEjz8MqKjPLm9nqFcO1EuJqnyjmRU97EgqwtvbX0J+ftaZ2CJB
8yPkodAbdheTfjzTGiptm9KWzxzZw5ASpNXvZEFUQ9WfabKf86ibpOhB9lcjyIwe
bPFpCp2WiAsr5YEZNcR+ptTsN6QzZi80Ru7SRuwk1w/Ds60P7XVrmEYhkARA7xxC
5A+cG1c42S3T1XjMHxWQyAsOFpdRpeUoxjkJGj6yAUAVi/zimEL/hgeZx79VARPl
cpu5I5pZaEOd3n0sCEiAlPZmL5MhyjoWQCJ2spKfv3Z2MOTK5+dLF1MyR3vZZ6qL
MOuLeJmKvdJMRO2uF2o1heGUGxFRVKjFGqoqfkkY6BnIjl24BJv+MMRkHlYdrOVR
OIgS7sLIEqP7dYrn92sGgvYmuv3Fj3wCvQxJCjmG3GBepv/felAv32EbfXIZu2UG
HVm2TD7+tz9IiltnQfjnXBbSluX0Ea9hNJEoJzT9XYpGuFIX8Vh7BspR8vOK/AdD
8qnbUULgMfpUERMjqX4EqaInI0uWviR2ju35wzwRiMZ3MKb5fErzyB4uTS60RBKc
1bUdVvD1BdJ9SXNXzn2/3bkeD8/JvYaqh4aRXvyi9TfVes5LJEhCyGtSmbhv3W31
iDFSTas2pcknTAFfUjhgvrzfPRZXWBh3PhM0siMuEhVolBgm/O55VcMrghcGOcM7
TXe8O8zidAIsjKzYMIWHH0DAkL+59NQLU0EHy3GGMDLxI59dmqMfOJ3lcu6T7sOd
L62jp5NIqteCTVhfXikN3HUxVKgbQgyiyZalguyIeBsJimv7boMJR4QstIZXs3cn
ZnupjI28Jetq+rx8qxFQOHArVlCj7BGIlPZBIsmUaJMIsydZI1bOqXY3KkGdbrS2
ZAx/lIjptzJ86VI9Qx7s48l5iR2ll/hnq96pCCrrBut0zwNvtSBqRx2l1cXr8Kjs
Y6ixBpYKDRcVPl6bOo5gLEs0p5HKqmWXaUKWzxDJZEIhoUSy4Q+2mRmEb1ljxCe7
nBlNF/Lzci+vhJCCfvLlzUtVbaADBNKTomxrSAjn3KyZMdtZNl0LlV7jX9lk5oSZ
zrPY32v8IkYKNwmWfS0X634Goxm1puzjanGsa5h/tuFygy85IvK2jSuzouWycTTf
s+vrdCe49B7EdFTFJTJNKGSLM+07i+DRfeyMXYX1T8FKidS/JxvxQxcyd1nAOfmb
3/TzihX05rbOqAhnjqv7qOVsErdRr2novDUqsufwkdDTHgUqXMBGx9VQoQaPYZi2
reoJXtHaqY4GZeSCL+CqXNVmaymQIEvR6ghCKS9yBVq6PoDvIPQxKv7RVL0rW87h
QAdKxYxgdlbR8pNC9gdjcyMhUH5BRyYWI9UgY85AIbqPwLJ/c20Y5ERL2wZttagA
e0OM9Ox4N7tH1WKOxDwhSGxR3tlu3NBhFiQorvijlWBKwokIGvuFBtvW22UYYmCr
bLzU4uPhAbdjq2q8JnAXnXkNzb9f/RDhHn/vabeCCkJLSzGQs2bm9MAIdB5Op5ST
hSqKEsNMMOpVnmgbUwfS6YiFfQvoC1EgA7OKvOIK3aZ8fgWl3F2lzvEjl7YBi4dZ
BvuNMYktVIoDM5YaCTYxAYb36CSzT0tavaO4wsXI6gdy4cJjAlfW/VW23gPD59Km
ld0kCmFUEAgYxn224Se2RojMtXKZ/t6fgIQxbOrBvY20qwxtnervcb4VJpbpxtHH
Wg63byL4P3cjvTUUr41wfw3w9c+aGgmKTKb2qmllUMXlUsa4fdhap64ppladxP53
f/yScQeGwftnnHSsX2WaD8AoPbX20hg5FAwYnYMnWLBDHrJqMwksPwH/+NastL5Z
x7APEROGW8aj2WhJnvAspAaehYecASKoP7oz5/UTa6f2wZFhHPOpN2cqffqN+ugB
sbc7zsBwBV0sr+S21Krr4g4hUGMFgsA9uAzFEqmj5VRKruYkWMgy6hTT9dbtC17R
5myWjAOyP59EQFJBSH4R2D2XwyctQZs3LPimHkwubZkmPtTSWrP+GsPF2MZZjSPA
5KD6iTB+FcivZH/4mNo9ApW7d+K8VpdJB46DF/PPto5J5lESjZZ1NNoyIzzRHOKv
P/gLn6+NUqdL7m9iWZVcIrZt49gARgZaTsXKlLeNOYoA1SJfNsMKvpeXNjFQq2hl
oQRolS1Akj/uNvhsOfvy7S6N1tUqvP+xbKAYPE3gK/qHJwT+QpDJbMN16yBL+AHo
vbWhcdruCvnbD5N4PDxcMAKF92sAvZjNJfRbbrYLw9laSDntoouiCglh+7IvAqrT
POzb6KWCtsgAEKHimGjecGVSTLi/uxRMA3AmJCvm7XBZMkdGEPlV/KvY7ojDQ8W8
g0/9afPIDhda9g6FLbvcjVN6EC1PxXymxBw/MpVcPFm8Vn8Na+aQmlI50S/AESR1
KtJL0+XfVfEoe3ypa7fnhRl+Gm+9IcZw5LK61pLvTQRRiIehXD/2e+leOro/lbKK
fgesgGHKWwsKXAi4MxAGUXtdkYJCHrAbcZh8x9cGjJAZRT9IpPN04HDL3eiRehIU
ONB2vQkR+AuCiPfFAgnjZxSU7nUDcTlXjwtDy/99D5th771ZHFOM8k8akBiyG/GD
8Rw9SK0DrHQ9tkctLhQIcvYzRb8reANaJC/OtMV+iGlTO/zVAsSJ/5xP/XCFY1O+
QlJr5N/5FJYMAQFP/m1GzqerkdWvEuElwOW+pldhk6N05v/gQajvABLAIbIZ2qIs
WoG7MSmtWjXJF1SdvA+rTXBw/R82UaoiKfWJRpIau8/MTZTaWT3Ha5BBoDZkCDhV
24bBJNxXK0siIWBM8yPyxQjRRBMGkuNcA3huefG1nvzZC1qXdHDeZlyo4EZEHrM0
P1iXEBbBDOWqNi4wDn/2BHwU56Mr/Bo3nkcZqUwlTsurexrU73IG8WqwdMv5q4Ye
ry/4PNGXH5OSeW+hg+ljA4GoIvVxAlCAjg/8Wp0xu5aTpkrh9Nk/cSi2nXBH+kkP
VR+Vj0CThTMZYP8UEnPG9yTWoHByb7k/EVXN3h7UJra7iUFh657N+IJeHNvfyeJ0
hxFsRRvb5nSydHLwN0VQuQFhGIxFgFcFL4PYoSavErNLxkD2X68Ns1ofwRAJeOfu
z4hASCxDFtLgQiEy/CyGQnpkyZP8Jb9gYhbZN4hVqpDdnU4pgyGfcXUbhKXpI2My
a+hSkdm88HV+EJW21Y4Vk91ZpZ2NYnKs+oXokDBCmVJjB2XR/B7Glo/poGJrzPEs
f37lnKKyXhDAZ22Q/qjoWaSnyv+QLziWpTi4ZTM0jqAFRWDjOI/2WQviBkezQ/i+
LQPIZ5geHLLFD8kgp/VKmj10j1RcI/KGp73pIk7F7pGXIZF/v7NXR99HGG4CmGi/
7yRE6v4/4CV1kSh3j3+/ahRAv1gr16wZhMs2gtBNsFja/ZizxTWBeamL3xESJe+R
3qsftpAzmk8nWinjyg2GrJan91kUCNP9H7Msmh5S4f9lYtaZosRdwWwwVMHAY6H/
suMgLmDoBwK/gQRuZMultDfMmAJ+NQ+kulT7DM1cUY7YIy40QoUywgsLuTcgRyCr
qQcilLnJ7izU8vKPw34OhuH4lCOoFyUmvRMGw/cM0Zf/lVC3R8s2HhV+E8zjf7yB
w3YSKfJmLFleL52TpNy4Nni/U8PIz0YQLiom4x9EFjt2smDJ7ZDbFoOC4PmLwjV8
f3PRBDJGXB3NRSXFH1VXYGczMLStwCLU/cywkYA/abQ5wOBAQgfk6IgP7mT3wM1I
dHMSq9PK087eVxVpkTX5heourPqXKDXvgSrFMdixBN+BfjQZwBaRlEMwiTqjdJJi
n/yGKmBmnd7qknLMgxsRTXHjd6w9HjDySbHikyyvRjtk52cMotyytTUPcdr/eJwT
VoZSdX1pK58TojN3ngQ6a6cEcdCLyUjqPKBGBHM8XozgNylDVruf4c134TR3211W
VyNkWT/tjx+YuvvqqHYx9Jfj7pL+U+g+/Alghr/G/NomL7AshO+jFZvZ21DN3hs8
zRbCohSxgCrij1/47Z9Gpz9NJdU+w1tF7+SIWcCB3hDrtCIDLzMssO0LDMz/Qgpn
cniJlHMHwRhLhRAUpIESUBk6VYm6Etk7az4LuOlHT0BpDGfyy2wP5SIjs2WvQIo8
S4pZkaVu94QCry8rrjicb0/t8GjSk0Y2rSFSq5obefEfVwY4bGndTXfZP/WPNsH1
sJb7Mg/POuvdiPUWnn4zrQEdjdCdQ/25+FDp9FI76t2PR5eIunV1NRNwC3dfEkTc
kMuxOXeU8qyiF8d53a/D39nNlgZ4UJPYKDh0dsX2trLPuZxHm/R3qmRSHv+b9oZX
HyywKgHzRBj/h8n2DovWyyaiZGnUC7OiyujZZDYTCQDGwQelTW+XIYwRGgQR2+iG
DWLP5YWwOleXDLmd0pm/wvTuL1VODrarfQ78Dt5YkzNXFlw4+hmcZceQpZ+2ywrW
ogixVXX9fMCHq6LXSbPR5gEBCcuzP5+Lw8Sfe0vU2tgNpbnmJkkzR1wqSYW8qkHX
krYpEDnjxL1TojP9DbagOIvpibE9XYxXsEMmVCgpEPNAxH+jJlaUjnEmYFTxV1un
8MLTAnAqsmH+s1spTFgk5pay1fhfusndxgFzn0vrJ5HpbXPfCS7Beo1q1qGPz2Mq
I4VAjOz2gzGb1P39R1vtH8MPSdTl0o313iqJFtHjHTtsoOouhnhvfJ9lMlAjNpn2
KnZrblqgpG8seU/a1lhgTBJS1CQ0ej+DQ+Kv+Qnzymt9r3NFE64q06pLzPCZMaKH
TohFCrkny+n3t/l1k0cxMh3YwLxQJLQ8oqw35+68Og8ld+rnHpnphaLuyx89Sbs4
AYxMZYIFE4sWJuHPNK6g8E15NHM/K+/3dvo6py0/v65yh+o/XV9MOpemPCg07XUM
XBQ3A4D6KQffj+oFvDlR7Wb6Uh06K/GYT6ZM/FtRLvxeDvBzI7Zoc/OBBzywCTjl
iTCUqLeVXydzahi4VTXsCYFj/gfVgg/P87Rko2bKurrJQOUqq3d9CLSveAh+Qc7l
zbqBrEQyr+awoY9F0iGd6bpC0Dq61tIFLdO2MVD1vIMfoeaJvtTJAk/qVzDfHy1y
OnfLZkHi7H8meRRlaEu7d/W+msDahPiJxBtD6RAkoLzS0sb0ZjgsyTPzJgT9P9xm
K6NttVhZ4Liw1y7M85vggwugAYTTFGlfkGbmTqbdXEw5oRoQdyzDeG8422n20Hvf
CJz+AKzz432//KWXCFD746/AuFQZN2x7OlVJoEV8chge9c//NhlbRx94BGVpvPwZ
55u4Ad8PUzMnd93mmG+KLTNHigzRcJjY9GPy1OnyUKMU7y89ikU+0glfISun2L3a
scZ5IQ7ikW0A7XsSvLzHVUHpqRbx3cmQZA7cVzlrpmewxfZIhuslp3Wk0uN0Iz6L
+/o2BjpVoxxT/oEc/YJglde3P3dxacTivYscQXeXmm5dcb3KHdCs0E2bpzssyO5l
iVda/6CFoK+pfqPy4GhfAh/xjLxP3vEtbJviQv9HvuyzCdPuIKXxernCC3aU8R5i
bpmf4S9j9472o7qPeO9x/GeQwGlaAnHWCeCnWKEzig8gH3RabwOjAw67N8VlO4+j
hNrYPy3ZXQv+KziHt252NoOn+FNjw/xRrkVzr1duysdK4XMn2mN0LLV+IEi+c6ch
3cLYZYwo50sY0numo9JldcTN3bgVLsLSzNfGEdnOpYqXsL6oi7gjWwalv0QgLmqJ
aeJ7aAJSNaXuafkDLlF4U28tlc/il+qjgxEVqatCcndFoe32Kl4bRTE/Dyb2oC/C
UfqajpOwUjgEFI47q59AE39QYL+ePXQMDks5ZAYb0V2AbKj/sDnJCZWwdpvHlsn/
rDLt5tN/YpXuomk/Mut9hrR/bfwxXZtTIvZnIfkb88zWGWjdjwVd8F+s4+jc0Vc8
2JEFOJM5lAm5ZPclPFl/yYYuCUWgZCdJDq44UObcqflT7KmTGAV/A3FuLuhSnfCn
TLvEJIRZb795PqWEfyQ9qOrh++C/GjU+Tr0INCZ4SeQoUqb/KCl34WakEskFAfbt
AKolIIaxfWPe2tEGnh3JVBZnCgeeWMDwwmI78ohLvJ2zrO2bDU0mbNe0Joi8Uk9H
xm4U8QrtRR7KKUMQKljeCwR/v/QKkRJRllgDEhdy/IaukOhsdej6eM9BA80cSL0O
LlNbKW1a6fEO5iB/Bl+/uSExqdIgkuziResodK+r9TqymY8L3rZU4Z4k0pcDJVvV
7mpCidbNZsePoZ3890czrJBhDi7AnH63TFa2m8upqKmC1sW+2dAneKDWNSetZAqS
xTJz2t0M/TxkP4zB30sMptfbZ+JgHafLtn31T1l8Q9JmLKdTfH4YpINF+o8lq7Wn
BqQjNnupjsFY8vcepFGo1ihN6PDZH1CafwrAb/+D0NAMaApvkzUSvG8xzRTlfxRq
x2/NgKTMjvO8DBf03EPSVoxB2b1bLnvQ3iN10TB1QPXjyAjvcZhje3VCAiLpiDr9
G5Ngcq73PytT/qQe6HlC9xNm88NdYatVhdLUhVIGaLtukl0Lnhy9Qom3cp+jcZiG
T2P5bXIkJeMnpi5IGcuegA==
`protect end_protected