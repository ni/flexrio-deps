`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 61520 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
sTHDbAcNdRVMi738hx0vzmj7ChpZsDQFvoCELwxLCIIaEF4SYSxW2gcr9mZQDvHj
rvZDBZV9ARPKIo8Ze75MtGnfLw25px9jhnTDnc659OxbDg15FMZbRBYNzelHKo5d
bTfZzhpEJAqFOOCpyuPfhZwgM2A+a+vL//WllVUf6vuCyzoHZ7TmdsrbhnQf3A2l
mqUW4x1+eAUfZ8qJlSLAXwwyC4E5guc8c7I04an1tE2w928a9P9x/n5Xqls+GB0l
IdT2zleAQw9BfjOXZr0ZwKPSA9fXorzMZB3GbGpCBXHyowCIyjzgLd5fJWR+iD+d
SXrGkqNT0SmKToBFzs8IG5J1rfPDUOuQkvTRD6xFK1As1+pPVyCMKRPfQuaypKjI
NlzUGMSkQCzmIjj8ZUMoEC1NEUbGr8e8rvFdjctyfdd3cw2Vm5OV+xa0V3R7UJo8
DAl8UGTNuzRlIT4PC1dpRgIc2YaKctd9dfrPDHIg9sn2+khB+AWvyiBYPSrkrF5U
FTPsrjk/nZjRpOJAs66pC1KrmKJGJEi2EAS78fNBUi7xxpifIHvBCo9swFOgNoFM
+G2HUxIlF+f7mDopefzimhPrMbSPjhePmbHfv2rZR+fdmTZtAJsH2TTMlXoWOU9L
rlXr6NIz3LfipbIkr8RTiNyTcxim8ekfPzlUY/OmyR3ZDREsZ0DZVZ/ySSCgJFD6
R6AInI0H3bM/xquAXFXFQPtIzubamBJi2d2RDm+WErzWlflC/ku4FGgJMnpiuTa0
FW5sD5MR1+izffCuMCfP/5Z0a+BLrgjg21cRgjrcwxAfLIj+WjAcuOOYC1kt1B/8
46fmz7c7CXAZd2U3uJNw1tuq5NaOI/+8uzdEZ8wLu690mjsHctZk2S+xFpPh5+ZS
M7wF78hkzdmEKnKLb0Ri2xd53FCHeLTNfmDQefKdR8zTk3WFbuVqJa2zYwPq1pgj
ZiStaxLhnFY/f5FF2F7MF5Ibxb6grkyBBzZx8ODo/TokFkLlsPigDiVfuz96lye5
BaBo2lI4GB+JY2Zqr4JEsBJwkC1CBQMsJ5lpEdcpse2yiRheuF3nj4lcuC29v2qt
4xtxN+1IF3kyfLRX1VG6tcMOwOThCrCR/LkB5nI3EGSa4XoVKlkSIHvMXQDgFnLg
DFSwqE4ywRZNoKwlJk9ZBiL5YpBVTa9AWWCDiQ+/CJpF0W4F5bmZ36J65DnTMvdk
TQpxod/wGPcxU4wYh5s9vd+2Gt1Awkey8qQPQTmzd3y91a0vN3ZV5zAxhO477lAs
WTCW9vbNackNEiiIoOqsfu9GbuYyN4M2QMsc05Y7Br8hzh4bRPdL917WgqXMc+cF
YtIg81rWa14PznhPbzKS5TXR6cKIJxuTHRNlmfSC37v6284RotthZ4z6aFGuThNe
CdO0R6KmxuXjRqEGG7yZvKbiVajOfs9puGuaf1IdQF4VQXy5juzO3IzprWmfYxmc
4G5Ewl5qyjg6UaMdvl7Jy80ZuVvY2MWEjeSp0ZUcjirU2VAaZJn6ojm6AU/K4YPO
s5gywYIcqrHNaXQk+qttY6J3QXaQ2uDZ7RHagOV6aIrkgFwGhq54XAJeQB8letff
KWApd3mvgUFOs/t15miFX+Gr3NxCeiFB/THEcEnWoXz4K+2DYmedgIEr988LGLYi
HKjjl+GvEFdts35Ae1KTC/GY0zTi5DQVIoFBAEkr0XzZO+SNJ730nl4UrrDJjcOh
+rb37YCkbK6Ou7eSMTURIKVIbIbqSY0E/eIHJEIYjbs/ucFMWgvKxwrjL1r9iYPZ
3rXPQOMMP4a58tZlPSpT6s4Ub0Y5YvSRs/uuhwbuaaKSHSSn6bPT14VqS171KXpe
tgadiv/NEqQF3u4ZmjMJoa2MsgKLBaq/LlJP6SB15uiWikOIbwLaEVtvMIQIE+Mi
xfjniJRZuqybFSvXFyqE+S5oIk3ocWV5UWStkhI6CVHXCAUOOlrh9gSFkjMhFgs+
M47XnymBRFGJFMOOezgEPRU6bOd4sdjB+KAB2+XisfFcRgCgTLNJKCCUdMZS78FI
+bHsg/pG/0PP/Jvqbnq6i9aM05UvZbXByvE/v5/5nEac1iIdBRM3rDdQr59em0p4
fGriKPKdFllSpbGnT0+DC3JA2Ah7VjkEo3jxqLyqKxhhiiHELV66pY5hcDbL06UB
BnWQhVxmCkZ3vN2eyZ6A62/vyDvlUROB4RdX1X6JAwJpH5Us/9XzEyArV8XEllDE
eQX5m9eLIpUjGApGdNHVIP+A2a7CRRlIgaUC07e+zzcOURYB6oiBJWsbq8EqvCnU
nmeLxPz5IvZ+g/BemmQFKbOHlyJoOrqqRE1W4+TmgvwsEMmLYj81Avv1tENichqz
81l4EGYfXMlDCbmQpxqjoqJfkq8OmnQq9uqrPCvkmACrXVaSjF+gob89YT98RhdC
Z2RJF4lveRu89Nm1VH84xja3Wma9ODxnMmTifo57vU4pQ7IvatlWvdUWcaeBXSot
3zKhp4iraQY/xXyIz/LP6de3330cuOjdXFelAd4/FydskRGD4OM+oAjuXUDJm7FE
gshrfyA9ngNRoecXklFS6SjBYx5X7TUB5eoePMnIRxVpygunSjHI+EHVT0vqAVmu
aMNzN8nXNyJgJWzsCep2sO3CYk4bn7bMiHzvInwVaaqQ0dsH/In6TPgzjwB2A10V
xpLba+p3ktVuEVgsNmMeNKtrB4hQo4UXaNWK7d+Xwjje2KMuQZCH/kSuF0kQwQwx
DB/wYGf6FsbQ1NDaeM3mCXpmXFo/WsGqbrlkSKUDfX3yc484/aFOd9/VSK4RnSF4
T6L0TidRkywYXTnS7au1he3Z6HWdpE/02c/RYLQCwTMJfRMed7QtnBo3In2yV5lN
EFO+jfEcGwRk2gP+9DdW/gLLxbB+qmhy5ntCfm6zFPJ8YNjFmlrDh9nqBlQWKnbs
ThVNcBWIJ4uzGeY0QkbWqRr8y36etsy98LFRsoG1H/3xKTvSmav4rCDVNyHhUIV9
bHboEiFZ2SP2xzcvdVSywMRYKlmmNtwvUsxY1HRDxR6Y43fb5hub03yYdZXZ6ogJ
W/kZUnP4Rte3H5EvaP5BfQG83b8hm4qCJysxNvgxznwSw2dAYZ0y009pN6wfPj37
WiI25mH5QUjZqbfIWK4FDKnraFSQUj6kxv5W//rTaZp9vbxs54C41tcvmYB0anOZ
FhBuQitRHXWoXuOPCPV/jX+Kkp/oLPuhPVg3keUZWqr5VMKPjPAF/Ma22wa6vV3i
9EQQ6bfgdJPFPUZ2QKJW0+qt8MSTeLM4RjkM6428SN1ac7dCDMt8pJL+BQp03ZtB
U23lf8ukE7C06C3ylzFPjWsDqFAcJJY+PWqCmbo8DxVVZgNjecViUfai9P9pzM4Y
8eEYl4fddERAhQ+0PjtRwiAbzGdnLoj6f9f5W+0osH75yg16jvovkjuuqycC4esM
v3wckvpjtK9+oXpma+qUqlFBMLb4ZkiMIjBOy6Sz7xkUkxEv/wMnyG/0A+b6rf7i
J/Bh78J431DZr4oJ7Me6LKmzl3EL/WyZuUZ62LZZ3UrO7GavS0f0qoW5+QHYAMCa
LkxJa0kkJqB3jJrw2HD6Gm9Z0VmUV5rsJyDfEhSsD3zAFu74ubcN0/qLro+K1trn
JBhQEGR30nZtXnfSKZ992AkoWgEvNrqp7XWPIO48wgrYgzm+4XvglA/aPEPmghWj
XRCh/CGWe0CCYldly/IwmxUqzvq2wnC2xI24GGEZ2L6lwtn6yR9tl8Jd4mfusyMY
AkrJt8SaxXodZRidYIBoivaxWbcznldR8POLxTgWrSFm4wGKUkAD7FNOvIkIjU3o
tImAJDl5Ob/ODOeyxgNQ1PXIgKOsCeahfaWQ1mOesIxbsQMiNQVtMmuyzbaYb2ze
DXBeUeImzfzua56Q2fzwLSgJtVkrdO59pZ7oq60tnGLTA7U3la+aGx+N/7Y+W3Rr
IK9JT9ej8mgfXQrSuyDME9WAgBPh8GhFBKhCLOWdZR7ToKFbU2Nr1O/8+rNLCz40
eM4mb7o31vva8r7zOHkUUOpo76Yaoayuw9SpCFbqO1k3nyuiIAxztc6/DnNLSS9O
U11CLhGasffTxcVe5A+jhnPpOEKzLENdWb78pz7yyQaC79kEqNYFhE5UGFJG2mbF
yvo1b+bgBK8Qe31MiKK89lRr1WER0okEhQwxGGv7shSXt7XenQ/GsmZTVwCd7AJ2
4IUYGMuonnJWsjirhAuyqKUvgxT7k33apxLXqlk03uTWQv22pYl0q4HTpfXmgI2W
mEG4yLKHtJdTXhuTroY17EAeflRsDNmBdnz3sEWt5kETZCwhw/RihrH992wAlwHO
lOstFexADklEOGuUoXmk7u4qTvhsFSmb5Se8mdnUZJJqvviWiljFnLvea8sfHJuM
2MGfOpiIb4bFg4Z+za5T4vUg5RRvq3+bQe1n3O7YBQMEOIO2D7hf4HepzsSXYrFC
fSjjxRJe6IZ1iTErfMEnSxICR72I3vk4zNs9OyZPemKnTiHwiJ5GnhYkUaESM4gc
tMxkqUfryJ3/ze098vUoyBod5s1oPHFBOBdwQKhN6N+NdvgQdVMzjk1oEPKeJ1wS
Rpl4eA7lYUbN0SldIUb4efxBJDZKZn+1Ug3WeenICXXJ1Hy8dpODk2izUhb4srLW
09I5hY/VQa3RXpnezJ85II08SvUTgWm5vrtbtxtOjfEYwxTj/2av1d1qPsJhP7qD
KgkomndErKloD9erSAV/rtqzGvCtiuWaecZASCx2qShxeOwnYgnoSo/HWFqUlBXZ
QklUuRVs6ZxIiAjhk85lJYan08V2tL1SAlgtSDKNXZ+c45zGbVNZxPhX03/VNABe
0jhSaTa+IYiquFbixjEevw96C36M7MP3THnkPHCvxQshw66rksYMMFvZWyTpE3Ja
PSc1c5EVPtBjPYbZwpOhz5aYptIiw7Kjak3UmpliH2bKjhGx9Gl5gq5phKGVCKpc
bGi/VSHr1kUU/lGdkzPU+Z957WTZoDvmwipibYCSLju/nL9z7OK9DHtC80gXlwtO
638AY9eEFzBx9UCKdbd8fZ8gQv6zDzBDq6e5JU25bzsWry1TAZXZbifUEiN7M+WA
PwN1eZDEZyCPRaxau2gdarqstzXsWkHp2dBlUS831Eewbv4pLu/7+B2sZoesu7AD
/UviNnrZJrM4+W/r56JBoCZY/bRC3ThtP6NL+xU2N/apEjQbIkx3CmPIw6zJlKAd
NWo2XSldqCeZnTjoq+h0xQS7mubZp9B1Q7QvqTcjqDjpDtGaYofzv8/lOVFmlh/D
ULTLcAnHYPwx+0Jb/VPW9DUBDPv/nyC+yEccJ3h9PNtZaVJUgEHPqGvVx0Uqpruh
r2Yf/8kmumAzQizBLiW6vh3wFEPL04mA9tSfc0S7vhKIirjARtXRvNmu4yJ/lmLf
4Dmm0kEQosWoAS506fn4MEzI7nqxlyKQq0KQONZ8FQOVjOKmulQr3q3a8UaXWv51
O9EMyN3Sy8u4TpZJUK0g5cHVei7w7BiRzKi976xMxBNLpP8jlPx1snSshVjFT3O9
Ip4cuQvuuEylIkOq18vgZWbWroLUYOB8aa4cOU+OH7mKwRShHI8g2NlhFqm08OHg
lN4UKmIA0GN2DAtkCs/w0Wi/veVRNcwWiIlLVLw1c6otg52sDuDbEYQiKf27tYNg
ukOLu0haeEGiRva00jQw9b/bpY15YTy9eQZeoTBLUP8KbJUWQiKSGfHMqMzS0y6u
qYsrOFob4UpXYls4kzhsx6WICKzOoAg1MAGJw5a6KR7L6+eSE8JxNPS9MtkX16AV
6O34fSV1VvIMlFz1EFS4TIXY29n0p3Wu0wl4ERXdgcArzM0iAN1DDgJTqEHokhAX
dOtSA0RfLKWGOqZo0CMTpmOQc52Ku4InJof6PdI/kZUsz41baGMIwoI1GZVqO9Pt
byBkaZIxUQSQ9/xSlLDKiyGilDQ9s/r+FoHGkoCmO+kOdXgC3CJTf/+HdDpILI8k
MGwT00wExn3qgJtS0Wsia8m7OiSwBo2lgl0X5GFM+E8V6++E8moiYnEEkjP/V8Iw
menmj7kZFt34pjajZU4TfDaRWqs6Irazzchdbow1jyC/QXy3673bU5KDcdyUaywM
/hEqal6CEaGJi79hvv/Q3aneSEO1d0+EZKGgMDgjU0o5xxkYPLmfNtHG0wezyIQv
Fqs3G9Wes39Xx24Py5XL2ssHTs3B30j/TtNWXlRnoLEeyOLIetJfnr7DzrwgGcuq
6rHHhCc9MgDT58PFHYck3B0ijb819upc1ajy3hjWArcqCtAOBCoOGZvakhKAhXGB
FqZ98YiVGO6aB445nXs37DCflv+RGpaWvWxlt++nUJByjcxRRPm/fHddL/0ui7Jn
dSr0Vs9a8xkS3/TF8ia1lzIYzLZ2dEdiZnVL/mmSzyNPB7Hu3PHNUDYUllMaZWte
h+6F0wft8HUI/ZWGWk44K2+izFXXg4oh9tM749DybmMz03SUK/IRKS5Tz2f9M9RT
dRkJ3pPCHVsXce6SQPqmfHwxhnzyABgPxcNTJDIUJP2n7Bwf52sy2o3YMPDIC8cN
4zFMGRfxiPRHR9xItjkM0kO+/H94QB9b84fwU5GA7qVdngWyuRE1qWXddKXIOMGY
OOjmAQAMw5NVpHsadTGXRavVdxuRhNMNtNrOi/VCI7MHvjRWfHeI2iMpzeq4pm0s
+WVVSiv90JWmt4wdLGFsnXX8NShZ8PVlZdfX5ExAp9r+9o6IAePprcAuMGmQchHh
4etwmSzQJS+z6CFAYNqpez8cy1HjBH1m0x3NHjEfgxvfS3Zwj0iqQbRunEBu9rad
jDL0kB7TBsWQLGFie6QYz8uYM68Qkw9aF3CYbE6AR1+GY3oxf8xRXVP2pkoeAqsE
1zug8O+7waeZa5J5msoiXJoTpM9DBJ3/bt8OTei69jjJzKjIbl+o72W+jz0rcl7L
VrC2LEctDY//j7wPDQqT6qTfGiqxQlpimA8NsuZAhKlZlwRJm9hGjdgHXNa63nsK
8tvYgllK+ZX98h7rWPdYjZCuKPaRFs7eFw14TW31hmnFs0oUYe5WRXsmArrunod5
nXhEnOUojSi8rJinDHWcE2uwV489kYneoJyfS5BbVOWR68tiu873PSfFA42dS0NL
+7RJ8t/JKreJ/dE24VP4FxjvlOGrpRpSPd8K1CCR2GRsj48OgCR2YxJ8arZGNK47
ypf6/49nAJoWNImHM71pXlQN8jKFXJ4Ax86j1XGGyqEqKKwMh32k8eugHCg4moAS
r/nXcmeKK/tHppyH6eM4kWqG77Ge3AwsvtIonnimsXTFmvqcp1yyPk0JJSBkyGYd
Hwwn9titELZHnBtzzWEa+fIJvYP3Dz9SBjzD1NYW7mjMAlrfbYMdqJ4y9tsx6KFz
nk/l8UV5ahOgBiuIOYpqbNiKlZMnjDOkM+JgKdY349FM9q7q0kUrWGCqvaxWChek
B7vhd0RIyyLrG9ocEg+132HxlxxCF7kwWTZCIc72hH4Ae/+FifoRE4N5XhkhHgPu
04ZFfzV6TtgowrVQhB3Avtx4IYbJdgq8nblTgtIJo9FwxVSjz8kX5Zfz4JfwNhz2
uyBQVHsrPtDXQ0fVDO82WVE2rCSX+AiLmKMaVHcXlNPQaFV9UNOpibuLqhGMP4ud
+PQhSHoZdQyNkl0ZSkq6Xb/vBEYq3e5oBLdg1O/51eYsalogFxXcx+y4P9kJtT3Y
tGvFNYylU8zyfC9UNHGJnZ1kREU4OD1VcPYaQ6JpgZ6/cUNmvjl+7cDVqVSk4m9j
s2ZTkdwmkQGtNFERqiJAF8UahD6AsH+mUasV5OtYzhzI+zGK8VJzcKVnXidy4Lkw
aNTrPNsJnZaobJUX5mBS3yG8/mSwexXjpTYftP7Hv/xK/9B/NAx2Vp9e5AX/F8FH
cynystJRrAqHv91OuDJDoHi/queACj4uU+lafHs6slAN7+fXxPByC6JfSM84Wuz6
nGY1bgGmGByVVNmeAXJk4k/Tgby+KDvNowDmT4MuCB4bLncMS8WCrrcZqVCkHd8i
17MgllJvFMalzmB5TTK+NNbEJHHzNx4+nO3R6YtFZqirTnpAzSQmqL+n74avi1ZX
yWc2iWSdcVJvskzn3QDQ/Ylxv0h5l4XewlZ6gck7oY0fldN9gl+JL50Gz0JzW3ei
rufQrBDQAN+iTqJnzbT8HRnkxqV2bF6MtGWwFuHzypq26GwXVhfxVnwPepVeUZv4
F2RXJKBRa2xOuK8siO8BERuAu5KiIK5EWB2Q9vTpjKOIdSuqPlDVZ/ip5qDEhY3z
inuNzsOlSKyRNRfM1d16iffIbn9UQoPdYL0AJzbNblIRU6wiPvzpz0PWQxG/rfR8
MqYDwP1vwrfylvZx8PAppad87vkL3iJ3NiJPKSe8u/AcvyrPE6ezK5VW2nOlNvTk
354uDFQunWVqYw8jybw8PjEu0Shp6Y9uOAH70YDAX275C3mptZW9a6y5EMq7VETs
Ve+bADfNu07R/21tVlAKjQtYTONMnMmnlbRwP2dXfmakjhfnf0SB5lh4/168c71Z
9+i8pnVmkjlpLWl8z58y0ABhUVntvYhL9vfoMbCGF9yAY3JdegDfvkoWwxEVIcFB
AFxLzKzXM52Gx34BbDTpLYcHfB5k9O8ozjALJxXiK5ShBCQA3ks2YGs+u2EptKaT
abPo30eWWM1Dii/udbWyH2c5w8ew5PgF9Y6ngsSM5zyMt2F0QgcDm9oSfE64zZij
HHfYUCsWLMfDZhV53JvYZ9VTZosY8VNfQ7TDA231l/zpISI6UnrrOMaqZhQYA00N
4X4KZV6YQ6MU0eRbhKfzkYCJffexpDTQK4OyQgwhMjW36qMtlVjsFgLqRuTbYdMM
VdOBYjJ9KuxE5rQhAlkq5rsTUXdl467nMQKdtIYRHQ2+QAKOdC3biel2eHKZfaAl
dzb+lXwjX2wjp/jVO5QEawxZiDFtdEFUYUDBVJlBUp/Q1xUvcTzr/ihlcL0+9f0/
0a/8r03Bz0ffohfT8CsiLyy6AU1Qrsp2m53MB3fOBpmtSsoK2XLWQA6KPPyw60Sr
2vMHJV60EA4hVjdRVQGEktB9XHjxv6nmP3jYRMXq5H5XPJs44IOce7wB3kZmix2L
2fls7Olx6BgjzUA0mpnM4QJBzg9Gt+CS6XDz1wJTbbdUZo1wum9hvcRsImKyt0jm
y78Zcd24IFh0smZX+TwrTQ/dc6xYvdm2hCeofN9agdVO/x3fmQzqVwDGlheE31lC
HjCU43kvmGwRiZN78CfETpQTnHGNIS0lHnnR49MV9mPMjUjJEOrzr3gi6VflReif
eGFeQoKizQrlD8Jo22JwKxBiT4o/Um3BkYW4b8fokDR/oqsndB4tfo9qFI0KfTNB
ss9tN1kf/gebNbgEbD8mw4WMi2RSxaO/xPck5gkYBWTid2jWVBdihRdiskCcIKZ3
8Oak7mqBKVjb/A+tY3y6MCyyhYqQzGctJvpTQSWwTlvrEsrnD2ylMsYL0Mt9jBei
m+zkO9YPg3gXWbMxO09tOF5BxzptBzzQvb5GZpZT4halSO5Jkzfv3EcK7rEmHGzj
k9kN4z9ebn0kunB89jx7hEPmDT8jHxID4oY4zoQ7ExIiltLatRLDynFbbMT+tE4L
YS9FrSbW3KM2Xysoal812vFNgP0/X1KgmrZrLbXV92D03B0FmyB3Qw+ZC0qs0swh
UPWcNNdfAlxWJWoyuLwqKPiyfcb5dQl3dLLM75PtO35hZMPgJ9Y5ja508ayW7+wS
aNy8wEh1lY/p54WLt0RzMupSV+FRg5AZV+7oRSNehqQBSTopVv2pv10T+ianXUoo
kybW95rE1xQoYbH6xteE5TgrYlA7J/aMz0btIxLNpI2kKLOaY19vbLxYChrH+B2l
aMeUCZLdhPB9TnbXWMJcNS8dttVNIXthhpAReATARhiPdH7qrfh3iRO1zGNhH1eS
9PTJ+67YyUSFSAA6NBf0PYOQ0PhQY1UcrEbp86G4n+MuJUAkPMuxlQeCtrlIscWV
Gpp5gNgfjyaCUfJOFIpNLde0F6uU0mHq61gFlRp3cVWEgpy9AlliZjmxsL76oAI2
EnLrxIhz4MnWuKS8p2Uw2iPNPjbc/Tnz2iGRT0kN8jBivR5PnzzEyCBe+yrhRGpZ
5DOETpsxZh6iMYMD2fPqkfu1YLENCwFkHYJoe+5I60haSq89SReTWxu+R/7QLAI1
XkcIhTf0kiUXxQxcqKJoXKLG3FIUHlOTc+dSf9HAeCwDbBvuxH088HhjDGGpNEdk
UknrKUlqrP34ZqT9RjarN7nHoAYychOehOxb9/V49ig2s0JFtpxOmQCKUPyP/VlK
V0PoFxCz2+VESJGWNH3NmDIHVtU0XB8Pz5WAGbeEISGnu8uHZk93ISU8EpQVYyrB
DPjDhLCQOOV6Y/IdqpPNrB7eHGFyN1yYW9EvphCvPxJ2N5E8NYswX3FiOJD/QEIX
+LV+dmSB8/pEGbxvEv2NKrKazcpGmAXL1zXtEcAwAZw2PyTQwota+uyep8mN52M4
O0XACIHT4MU+okQjqqTMl8NwNOYqJNU/7VAzgk0Wdt+7V/B7nWZPl0/jKSewAj53
VDXNTSPIPlLjdU2RGwMXlydUrff1DSB+wcLUkEyg7qd1zKxhvmZBEogRBExr7mOm
mAUt971a/KyeLUAGU4X34zlA55m3L5EbqjL7jjT7HwUaSTqnofaab0R/zM0MCzCo
kUxpG9K8eL3Az70US9njYKo7vEno4TeiwRBvc2vn8yiDysSDB/LwOXvVWYXWh+5T
AsAcI+PPz0SdUJH8ihT/kbxJqP0ROtsgih3ElLOuZZoPvLQDpAt8Uqk1b6xfSyr7
IavE9qXquu4DXBNy5/IshMP4JWRM5FnQzG/zlJNCJx62fFAi6KeSink5zB5AM9Ij
60+f/brORiwn+giXW3JGzq4oJt+JnFGnRFOJLShLZG8UK//DX0N2V3MTqVZVmHZH
xfGJ2lguec9TBAT2WeLK/4+5LZ/G01knK/Z/lOX0kmsNbYFCRU+nKSpX4tvc7imT
JCRQ9uFNvqEPEVv1QsiAN3d52Se5gRumWLaREfzf6xOVftCzUCmujPwBnXVipvQr
B2kem4t+TA85VS+MXep+KmsQfxk/IbQCneNr8Q10XUwgyQRrXz0otsCfwP6t1ZiR
G5FXsFXhI8tuHRoPffvBW97FcE2JOxQCh75exLqzeyrxAPB7h4y53fji7PQYsSXL
g8XkoAXTFYPoc53aZpwFw+soGP2wx+jsogdmWNqfb3GrPV2XuSR9YAKUWhxXs01+
e8f+y4GjmJvj4pp/+AYAV0bEbJi6Q5n2luDrWew55i0TKr3Tf6a7Bkmphe7bRUks
ZFKDf6M6XSbcjDqz8ROmTjBvpzYTTpy4yT+ETsM+r1BoKWl9oJpJClxWm33EIN8M
2wgrJoaeHOKhSikozpaEbzmtocy/yYUEkRboqcJ+xYZiXeYrYBZJ5+1sIFt/A0yb
iBQcViAURPIwmSRTXU0Ea8cf8Ujk4bU51xaSxsj0qk2tUvRARQn2VJCSgIHPpqgR
w1w1CEMo97fKnGhxsp5Yk/jycNKR3s04tMVpUxdFmGGZQ2gFKkxxQ+VXt0y4+MwM
sN4e7Ue/5gV+IbstbQqua47KFE70gd8+u/u46qe7KRNH/cjRElvy06R0UtkPJpDf
dsDwvYDEgQ//llapuiJzrtdowlgQeAzd0ElICbg/XxVTm1WVAq6t9hPxEFyPJPth
OAxkZfUc3heAoFEqGTGNWNQBDxLM1dTv/yDOaWWD7eUUFXpKr7lp6USwVS7Fzkou
EdeN6kap/SThQMH33kvfTULgwf+2xu0kEEOIlb1pT+2aAfM+fWhBbonA6KX/mgwB
2xsSZAYagMr0wyrrUt7QppzrcHBZk43oCGkzII7HbkGKq0SbIfP7TGUO0rNEbDbD
A2d1TA8FIn7LyNUtM0iqHQsvLpCZ176PMkcvYApwrDHyCOigYe0Y+lDXN56lWIgC
sBaGnVwrjWsSINwiqriHcintE8MRDJiAiCPl+ed/3W8yYia6txFHj/n+Hafw0pYT
EBEpkJy/drs13DoCdg9oiquptW6Alfo24eqLT5SyJuOQ0spu17RUw77Kpc/n7edo
PolmgbxX5hKARlnnwvb5qnB1i8z+/4MYOCyob2RXx4c20IcvkQQwBdjYmnbTQgAC
IXFNsi/VtJagXTm0o7jZVs0uE5aWZB49PyIrdQb0BYPHFpGM0ik0sRgRiaz2cbo2
RKFY+iCYtt/ZhM1dERWcuDH/tRggy1aOUfGEBrLsuzco0NxBAD8fxtQ81NqwV2PS
2fzMmjHqicQieCHs77jOWNBSBUjLqy6RED0h6yCJVnZWOyyw9fgrbnX2dhTujQKb
swYUxjUi1UKfXYpV3xUpt297vl1M3zNyBZTr5teRzI6Cp1Er34EDZJB0v0mNAx27
RP5IwxYKbJ3pwz31OA+01UA+KV5hotTLm22svRoBq+xyI7Jx7SycaQc8wzkTg9ZA
hACIGKaxblq8boDVNCmRMY+VNM/YyeIIRHer+ZnT/w27Ev42QhwCrJ6Zq13S/Os3
8MPMKhz+CqKABtqKVXCozaOsg79a8n32FvB0rbvG1B0x7EInY0uqw5vqICKhAb0V
M99Jd7yt0G4vwOdcIcijoZh541ZtvzbkVFr9tcitV2Tl1EGDEojfQKIlK/IXqh2Y
qWA/rIXv5T+w9THZuYFC0Q1lDZ1gtZ36l/zg0+9yZSE8rgpKRTTgVAJp7v4kcrSw
nMfuCm/im0gbwtQUbrnTdFMb+30jTGUqbiNXmCGfQXvYQMA4SH2J88GiUIgljGdn
Ly8uLkm5PxLKyolndTwMDcGnVqSKt9zAkZ7IjR+NlitRezGONyHybfaQWLTfk+B0
S0t6aKTnQ6undH7megCLX3UjX8H3h4mAWWMmv9X8rppF39MWiNBzUziZjKCpH4el
VrxCKygQO8RtogOjeZrVaBug/X+8ZWfgQPOJ+59eFLEDBabNuP3DI180aIqumLre
u8SBmK1iTG45zCkS+EzVZCfjL2WKh917waTdpB2KW9a2M2aeS5Z1WUEXp2Q/mMrU
Lh2WK8h1hBxrNcfChOuuExExGtyT9Hpv9b38SQ0RdhEoWg4R8jPguh+s5XA1f2so
3klsJUfxvefPwgShprTu+2jX3n6qb2VLA+SJQNaHNmmohOWV7WkmtUnAaxeFKxFQ
d/iZYi/soaz4StI1KF9z4YYaJC9FYAiOLJhV1YN2Pur0lZGRW5m9Pnk+Fqh0HLJB
1Gi7hY3vrsQawQZbZjMSF4wxHPXfqbIuNm4seZ1zxUGN6V9KSm2uH5M6H0N4Tmqs
76j18dU25YmGfsy+pu4VnlNy6Zlw8BF4jh+tyN9fxZN4puncjxVezB1iULAizc56
Z7GmbsaiPAd2bKuuz6/ZNzWUvJL5w/jPeyGiAyOUGAyOyAv0qvAgw42AJpRHnD1a
IBE8G8rO7vDhrRWKZ4Z5y8uWDkWFejmMc96/MQPzKRf0Wzj3RkTJkeUxpG94oIA5
uAQQGtu69snmqfjKJmynPNHNCsNM4kI8LPxpviCDvupPioZpGIWgbEqHnL/cwd4G
uYdbX1vpAyCI4TlGxH6GZ3cnvQ0Mvp3UTvVqZknV+4ABQXc+OLXrouUx43CnZnHb
yVc9icTiY4jCj5jYOuVYLTQRI7bkafuZzUB86zJzg33Jv1efXF6/95CeObixPURs
OR5bSVE2kY4hAU0bBLfEzNdjWq8l7vAb9+wdgQ5m6RQjGtlHlngE4uzHxWm3cqpn
66a5+GVrIakeyMFfQCFih1X4o3IjWo5XPSu7Xtl5ClX1U5HvbIS3N8P4el+Na7Qn
y2lwD/POFHtGUaJ+K9JiHzF0OgFrPlPraXi3Bl2JkzHMM+z5gYMywvTmHfZKm/df
Uv638EEpJcMdafxBzpzjQuPSKcfE5BjjEvts8jydqSsEK+765j/BvLie5kAfMuQV
vBMIHyu1rJkxpb2tcGdqvVa1vN/ThwPNlz+/bdgariUOOJwt5OyiPTzdc3SEPl/0
tpKiMPTaa45yZv+ZxXVvHQwYm07R4ldlJ26XSoxbrBTnhiedJ9xThQjUkZlyT1hl
sgjx36yuEXVTMYS/sYmP77AeZrX+lDWXAXwIY6Q8hZoSDzdsOe98BcRx1s2SvpIW
dTWesmTF63+8A+vcgChT5hN9lCRErolDEoEIrowY/4heg1hu+3L6dY/ZR/63+bBW
gaebFGED/lzFF8aXlXiRCQWfnv9dP58PnMPpcJ1nlI03b6ANW1AWsxbEgmgvWAKQ
utznuDxiZG50J+lZwn1Fz6xy7TaEvYZB1PmSwuZTUNXCGMIu2TnojKIafQbOsDcS
BB3YM0L4vYfZx1VuDone5nbHhFSRRU/QEg3JbS3kZrH65alu5MUjP2cREeWVSlab
+5dfVCVpnPUtwqluVtH+lZ7ww7FnixRHpaOPDfeuZlK8RHyg+dAwQB+jZJ8WtWF3
X/DYCEutNSmnF5LXL3rixKz423tF4LeqIJhiHxYs2t/8rKC89eZZ3xYHARY60bxB
hvmbDv/M8WEy3luIdopyBiCOBOCdvIczuNqwlpXBTF/6wbnHo0exbZgexnWODlCn
GpnFSlsBCdY7lC1EyV2rLYwYx47FVH+Mvqd/W4ZDe3ZAF0eQTnTJas3LPAxCKNRt
o25DDbWTxzBxfKWrWTvw0f7cnvAGJBAY3xAvxsc7dQdMjml/c++tpb7HCR2avNMv
I8ju6Y5EZehIoBtplusIY6s8MnxMx85507Hh6RYXSeAlcyxUkJ3czh8RdS2BhgDG
7Lc8iPbx/ORdEkSHZNOLGqFbN9PYdKEPY6VhNpAKds4+kNDAJJhb3m7JDTKWso3j
mGcg0LJmODcTuAC6iQP82Q/ShTDfMBlWqIsLJcsm9lZT8KnaDApIjVbu4NVJ9keR
V3pzZNZuCvvat4rp1R7xTMMyT0hug+HnGCpxxt9YHfzbaTyJt5tNui5k86gqDgz+
G19ztA4nfUiLgkwYBBDVlqEo9X1fwS9SQCNqmZE9G49ROIosJPTae6E5oRjcBIQP
6pwZoQkxA0xl1GGbyQD+E7iwJIiL4ODAoDUVB1QHl7lgEeIrNj5jhE+bkeJEdl/C
PTGeXYOGeqbCcAMq5oM+7l2pgjc3C/11Sd4nbL6E7cPWcmw3O/lqp4YEk23uskU4
TA+NQBxnQIvamN2p8hGDdmGEIhB0YeHRCUMo3tjb+LmXAzCZnxPECaCoB1Zi+xSy
DdU6V3xfXQpFSAWFmcaWaBqYxsDXyRsfGRb5XF5Iz9YCJC7ePgRpFsxtB4hQ7HCz
jHGxP/5RcINYwKLYxD7DWDXgIQBMmlSwRRKgQI8uwk2CDhg4ICuMUqLTzO+wUC4S
ZyM3xbjkJqatkeBeicLVOrbKHZ/OzeuMQMtWzgocFKPxwNuHE/cu6zHvSdsYSVs+
HEv7Tlp2sqw8YalSIC/GUixLqOqGg1DX+Lv+7Ft34tepCPpVoMyE+XBaTxJAKQbV
1s6mNy8oTQ5nVwD3sYJT+7C/xusA1UiHrlGF9teSwmtv8veg3zPIsoT2e9GV6x2u
fWfatYFQ3cN2T0jGB94L73HETL3JYcyJjkMMVsfQr22cwh8qhujw6zFruiJHCz0g
6eQRb8mZBEq72EQjDenF4wQ80iTgw+LceicGTbUDPjUO/AI7UtCSfsXJ7AiFrXml
uMmQMFNl5FpIZ86zN524Yhiz9/ErIykalcaiqISPeWGHl71sXpnhy1XvJGJGcjWQ
LPK7/dH5/zWXGZegdyfImsc8wcLKJ7QMiKH9Dvb2zPY/xABpQVRLTqku8u2GVoI9
DMuVIdoKu46RWMzctAotbTJAXw2k9oW2170uavUcqOoXQnMpZ8oNojpQMPjmXHHF
zeFWGUWVBh/v04eMaij5EoEU01u9NtVlL7Hr6AVMYYg3Pg0gM8Jz6HQGGgF1oJof
+iRax5l5xsVy08Yk3jz0oTQBznj4D2kF3gXL2r8zmDQowYGMIWNaBVAHyMdaTU9o
CrwikG+OpKLKAr729ixHlqa2C8Jvv3Ud8y4rhkCPuTeK5WpbA/HLq1fDSHmb/FfI
vz/5TX+H9xvcQZ0TgikedjXKtEkVSnrr6oGpPbbXzliplt9iSMKpRl0QYMU5F8nN
JjOO6mV71huOM18S0xC6qvkjpNYr4zC8GmCdL4aq5y80pq38bwrBBCpIvrHuc38D
MZriaoF+WbhVSHQop6VrVNNFUMYaC1adslBNb+zZLWcndejxbbeCqZjZMbW+AnSX
k/VZzGpvy3YptQxEwcMow4h2fBu5TZHj7s4kmFdCZQepSDuBkttXYMTi8P7WhPWV
5s2IymzxoUGJS4phLOjm5TFIdWCqUjBB65Ws4gdyHQy3RCiihF+MrH6+PHibqnDA
0SPdJFOCO/xuboXzQmeift1a0BgkaXP+C3sMzehwGys1j7w6mvVp2Hu4DxOfwe20
iZ3jYB1QhACX0JYEgxVBa/jgO5/2bLiAOtwa6EuaftbIs4NSkSXvRByDclpHXBLX
t6GsoDiiF2XhSs+mqPuK8w0TAOwjQ2ypuKKPjnVGxx5bC8G3bBtm6g0iSTDIT6Ql
f207KWTYe300I9PNVTP6rhYFJm4zrw+9IYnD/OqoGYhQkkp1+o473AtGXcZdajrS
QMXG6OT1NIPJqoVfCURzblIkKj95PgSBo3MmCKlfvbIkW9MPPTvS5EW49898jEZj
CBnxVzsUyaGxd2xEQ2bVY5gmbqXwBIGW3EMhxI/MgLCKMjI8eXBWEyx6XpVQDtvD
2bR4J/q2h9cqtpxAeu9IQNkTQE56nTHJPmfcdD2T+8obySsel28A/xQmmprLB3IT
UVQ+EY8i2R5MO5TBjqsJb0xwdfsi14EtJG81y4+C2csum1qsG/2n1brvrYsEPvui
Anur6Ek0/pK4LhmHdUfwnItX2iNOO50CVVw+3pq3tJ94pJ+LVSHF3gUpPJS/LJDI
1VT5J3rC0yJa3b7fut4Vxw49JDJ4bi/ZA93gj2iYQaMfmptL6Dis7Wajbn3A0NaH
OTfEQOHXOMK/YF1dt0C5O2Ov522bsKx7U2CUN0fnJVfVN8RNSEcCN5UdXpAyAON/
ne3Hug5PL6XeZec1kxWk0m56BHwTeTv510yEh4NgetEPv93cYVPj6tpaPHgUcYCZ
LSNG7JIiMFOdxtFoKUhg2hsJNte0oeMwXQW0KirBcCD2kaGKDFtOBTk49+jmrms7
NTsoRO3s8TQk1CvIZ9h/xQHqX+eV5ZQhMXoyt6ceQX2ep6X3ViTYbYARE91Q0k4i
PLfsPZuVvHiN9mvauT9CuQMEDutqUneunva7tqsMgVZNG4A5NDJaeInj2v+vtwU9
uo3FGpcPgR0xjpFUIPqcWJZk6ImCVWl4vnQtLEQhSTi6J0hJRMJjbLIMlbsUyMHj
gMOmMCaALfAAzuZs2IkXzuLQWKhzZLKTFm8mYwpMykHmdcWNCVBQ56y7YX9aRKRb
NaMBbV1bdg0zUW/JMwZO/+kY3AmOv2gEJWiL73TlmAK7bjBLES0EiM+Y0WkCpzIB
XhgcyGJhn3nohuaRPheX79oxKXG6gK5j3sADY3a9vVHbWrzZ+ZHiC14nDMnEIL6F
t1Kz2H3TqlrUCbFi1j5dObi9E646DPULgOYGWqloqr840awCYvZJ2O7iGvFY6Vhf
id5FBB6S6dbrYqvrojmp23iahGOvSGrLomPy0CMUmdIOoAYbE/Sw2rLbKJrPikWw
oymG9VH1m3E3cuSKpFaHbhs9wRaRvJF9qtoy8hiTNOuM1Ej4NVO7cJjYy4tkm5Ch
ePLgkLUbmPD0mUCQk91IGMkOD+PRa4U+TNMh95eFCtMJ9d9iYa+PVhIgsNDhmhbW
uqySomXeoP7BkXQHJSxcTqF704EbL8pnnkE1cmSX61COsbHZbsl/fsrH2FeG/ZSa
ePUl4b7aAYaiqGkrCrgpEE06N9so9dIKrpdgpGhNN00aI69kdz+gCNwtHULVULFG
8LSnTWC2UGxOpTWNZ0Eo+/a8JVZnCry2NyYMRqXMJWl9o0cISk8F1/vL8/DfcLYt
7Gkj+NAO+IrfqFLYs+lSVdoYPVcc8QJ2E4kWFFG3SGQ6urLln/4zy/KFwG/NVUb3
ZXfSxLn6XmLxlskjzlANmOPZmY4PYn98XDnrd5T8JI3ue7sf652rj3ze4DO5wZ/0
59mDwtgklIE12DVuJy4xtuU47BClQHAnM+QoNdYMTTFA9CjPWZfSKVa4WEw7e8cP
ezOdAaHmvrRvNp39yp9WSyVBRmIQPBfvRLvXIyA+Z8E7M+OKvriF48nEblPsw2OZ
eQarQZ3zxh73q/oXhzVTNFgGn4HFEKqAiEhR3roGGG/R6llnxP+S2Ew7JtkbdJr5
8ozD9g6701p+irEFvrpb4TXz3szLFKAomPS9bpe7dcjyMLtaUvn5yqV8NxjfcRnV
WYEwcgNKHHdhWaUvzK5lLyG1v8xn1OE2fyIvotqAlWUMWVJy50qsN8OuBK4Q6DCT
ipDsPXh0yRAhCp+zMzPtztE3HgT5+l3IsCJP9OCPkXzGKSnIznqaXVmhEnLqDBrv
ESb2YprRsqTCDVuOy5JNbSRETg2cXNdLVetIsr5OlfOTqrQI6zgnerUoc/fM6297
+XHLdSQcG9gX4BYm+ongdFIVwU1noALWzBiVydxU0hlk04UsIHTmRMLj1MP1P4wm
xZeFvv3nxutY4UuDg1zW9u25ffB0/DUFpYqZyHsoPtcb7RKnUMc4aj0iRmtvSR4C
Gw5AEoFM1X2k2Ofb5fEFQR8txLYhXpQZLluy8j+fIt0GEUQL5CqyJVo4+OR4yUMz
nVw0lXKWTkJxJCDgCqgsKdJzQnhS+R1zYWVoGOnDnlMpCsiVuLESj7qhsmGiS/Mq
RPmValLbJQiLIZWJ/YY2JUtxUq7pv/1i6kfIsyfUcuGcDyFa/GQrmoDDOb+GQXKw
OUFcGJjiE3nLvIQERPqxbNAP3Q1ViKrl6hw+gKlMbVhM7Fm9E9L1UALOjEaNwh1w
cAYB1g1VsYwyF8giueFO9l9Yi1rgHXaJVqfmjA4oJ0vqm25LY78PUdX4qvH4uQYi
pLFXKkC5+Sa4iU7hXGaOQCudbp2IvEHITEeZ+oVTzCuvX1AzM/eCq/aMd6uymxbO
HRpU26PGVA5/ALiamiHbW8u9EKmQiKJ8MyTm3v9ylPiSysOCT4Jy8wHARFigqGfx
cksO4oXJhvkjWEJrB4VZkK2JChsVvQmFYr9A3GkA+RUw5+uHCApH6cPIjiayNyq3
QYPWy/c75n61waHj0rSLE8f1ABc+VdcrClXYxBmPOX6nTcSpgntZwn2GTgwnqbNw
qqimvw/Q4F5vf1AOOmG4qdjOyq1tFBk8cIJ8ehDTSyPUgaKVUFLEuYpSvid6ouAd
UYRpPU71FOaQSo/LAOKd+EfodWtW9xgZi9llG4VfpTGxcYIdedeoOy5xuqbTxAdu
qN/bj1npFuX2JQbvhk4SdDEQMVicB8np7BWHkXBAE25fW4loAMn3F2O5l7Vm77sA
JHdDK8YEDDVsftfXUy0I86RCKQj9tcwp2Y8RKLRrMWl+1YlzNznUyeiIrKckFm1G
rKP914V2wNMaiBicKATsIueCcXNE/gC+fvwugkh4UtbnU+7Yay6ys2jBdt6/JVNq
zX8lpnaXHm1Nr7q6eOzVNNswlK6iHiNLyDsBKUWobl5QgnVkfn7OWgVTs+wHtOOQ
iDpIMGBxR/KM2lQu6ZjqIuGy2wzsXx2bSSUjCDgP7sWMLI7+zZRC3XpvXaC7J+9B
ID50s3DLutFxti7VOKNmW7Rz+2WEt6KbDTuihkRDpWpn6NmN5CfS0u1DUy+J6gbj
JMQCnyd7PDpJDQ8zJ2ao+5Edk9KZSch50c2O4D7y4RzSCuQ8J1kewONNuv0VxiBm
5wDQkMwWvdSra7fGICJlQin5u+EMvaTeg94gYtriq4Dm0v/Uza4egcEyTWkNpcCi
oiD57T4uiGcIsBNdcZ/9tLbSQBe3ybcLzEt8Rn8tcrY2uhbwLhk/9vpIXg5l5gaY
ToZ5xqPwY5fSy4cdWgk5Iss1dUiK+3Pf4dMyah1U4HpVL8AJzmiDH/PE1hb3muTN
4loJBgF3XwkE1sGwuLyqljSzBUuTdu/lwI5T+XBufYpq42dY5QrwLe0GDC08O4fW
NL0injz2UPHcQUttHfcRouLobLUfoVFLWj3bRzCKqyYIwVPnlMtor0jKNZLAcj+X
2QYD8SImyETVNNGf21RmGL2XJUIApANTPqGzSRA1x+GEFgP9YAq6cvzJleZOFV3R
hOVdNk5e9wbqWXxqVhuQtG9+c6s11AyzORqkqq4+yRUXUvx2Ab7MShG4svywllfd
VTC2/3ILXfTdLvZEfwj8DDnGYLUl9Kq3AGgZWEV9Otmbwt/LGZ5x8dz1SLcagIpc
3bw451jOHqNOB4g6UpRQezpm01kgHY5lwE2N5C7mMnB6KwT6UzlhvFlZhjsDsYfU
oj/w2Q4h2yEGjLE1o2kKm+H+8DxMneSmVM3TV+2GTezfshep7xVP6MfAhpWnY964
gGo8hRy9r50bRUDNFMiYjzM/bFiSqmR7YfPKYoAi5qeOtzSYFlPGpeGy1vDm1lI9
Lv4ISPb4Lpm4hJWgSEQlbNYG/hVeVSo0H3OPuHL5Z/+UyrrMIrp6pW7Bdf7BwejI
DZmgNp/JjbB2Qq+xRSnN5eEqi2wRt8MyHlDfv96AuSXQBjbcK5+pGh+KETte1vDr
dTfkkUFpPjE1hNR+KPR+NJXKnrzFFJxbKkoq8YquHnX9G9QGMMan2Nz+YIdCgJ00
bA3f/ofAr8kt0ajWbDioQYx1kZC5BJgWPy2o3LwtiBFy5zqSjpjlvItWqDlEaxkH
cNF+DjWWgTFee/TdS9iRmqf9OM1eH72FnzePUoNiDyD1s1o2c3w5Gyxxw3Jala7x
s8Oh0pZrBOayP3W8ShJFflelmBei+dvtDgcxW9ctLF9WH5UDX0+JHhWoMkfVFEL/
MXzxg+w+1ToB7mxYlFjpgMv1yNJPftYkIdbDMsKXMTNJQZwO7VEok8tVYxYCiXeK
A992f7pGqbxs/UqkFtjkV4VWw/9nOUBzRRhO3g5L/zVp9DhXQR+fTN0j3tOls82m
LPuB7GAN2U9eplXhN9vCXqKvlKpp/6/XOq6UT6jmoqMwaxEhTcZ9ejSUt0S8bB9n
rrj7BZ1qFAAkzy1V/78pLbnRvb7ehf5YlR3VM2Ph2mKCB9FwGCtxQHwWcD0emkUE
1hPKqia1k99ubHUKCBYr8lMuPUN+lM3AvPzXx3Bn4+qE0c46PE0ireyG370JzWri
oUHdOTXvFo6bjb8YC57qIO4cfELqwKfiXm6x5clZz6/k4bfja3COX8Zepi39HBuP
Bl39mw+8FEgp+O38zTj1qY349ShI3tP2XCisPRZCVzB+CCquvE2snhakHuMUD3VE
rhxTO9mYmyJJx5NIeODkntawYM4vWIluV8QTKwsy7KQkm2qArQbYlQExdUK79h6Z
FGfgfeq5Rb5wBlyOwzq5FWdP0/TPZWhIutgv/ao6RBNuHLjecnuFwtJgCCc1JTvC
I5z5JNhvqrRyIvAveSkgMRorcKGFJGKcmzrmfND1q6opUBN91H84cw3ly3F0LiSP
/Jj60ZLwv/v/mtrKSjmGYWnn2p6Rn9vzI3xFhChaXLCw3TSWlqq/3mVuIAbVwYIo
jkrH5F2LGW0FDQOIqG7qvL8V+0vIBsz1rh8dl1jpTjdSw5Rh5BBwZbs5yhjPBzGS
SqbrtOlckarN5Gi0vmY63UH4obn0rIDHsqZq49bBN06xxmkl7uur/veOpRZ9lgsr
VzTdw5JtAQV0v4X3Wpv3SrzaxsgHs6yferK6QjRrIE/GlovmCmz1W+FahOgJdYYY
ky7XLemugOMRXcNEzNAf9OiRl2VejICYiMrHixnfZT998tdXMjV0V3uXjbeieUR8
SQeZ76mEAU611s7yylQEac21Ohb/KbNZHhLIHTkGexN450uRBmVROSfODlpfOpTF
zbXl9KgXV0D+kVO63L3tWgjDWJ9+yXikl0fuwWKJ6Paau6PWZvs2/KmRnhA4CdmB
ar5Mkmz6wAk82PoINn5eCitaYGoCcGKoeMnYVyExg+TClw3Rf9knkDv6ZVE0FYme
QO1OB8PkkYzQYC/3tU1KOJl4v+jFW5x9q+3atLKWQ0ugC4X3FxasWmq3RqoS6wTl
+Tlua2uVknqiFAsmJM0JJntDgRC9KfsujYtNEObYdDe6DVev89FWKfK1QK85Jnud
g9ZTnN2/NoCJoRwjacAQrNhvk6W678tQJ+ksuAnRk5vOFc3gQ42ADb4ixyINWw3n
AgwTVn8UCImsYcp6452+u0jp+mfQvFlEUanhtuORUGa6UnKsGWtD67xLw46MYqBA
q5dabO0U5LY+Hks2sVeMUoefQcxyJhLcRzLiYIMlERK8ltD24UMi/aWkrx9l6f3c
PkECdxhqRrQdOcTu5hNMoyh3khc3Gv1VKrMazDbCQWqbZCNjpmNFROh0dyUoq5F1
EYgGXhX7fV+KZjctTgR7Xv4elGMslsu2pOgxykan/MmFQ14JzNIFC6aCowarNZp7
IOt+nslG5v4YC709TtWv5lg5VkF+p5gQeT2Ytn9Cd7WyXEqYcHi6tv5ZxH7kfyvi
jtatgZbzUP3gx6ki0BQ9dGPDdUIbHhNT9heyMDpilFf11l3RVrJ9LleZ4/FgNwQm
MzC0S1efi/D4oWhILA2t8Bp+jMDxUJbkCKko1ioDLaR0E6VfhCRpfImun0lIXmEN
iQKWvgjAGA58SjHRqmxHAJ2Emme/YmYDxUJO/KYokyFMqS2mF2/Mktt32Xa8O4PQ
z0G6r8NsKD0jWctzTTfaPkU3UdLt6HtrUxrEhSKKICkJKuCia1Xs5IoHUNoGmJsZ
yNY5TKppba2WUTCCLFSDxqOaAZBU847uToaSafnS/LLlldlQIJ02RNZoGY2coy/y
BKNVUFmDxfhxtfBFkWeBaiWylULouoxHTzus+UcQ8/KkCjybID2SxhCOuHhhnnci
+I/3M+/XY6nLb50xOPhF12fGea+zw2/FgQNaNkS9QRFvm7QPLsBFsqUmKWB/n0ky
gDO8RgTw2p5i/QRhmlRDmlemGWyjzfm8fVvsAuk2dgejMJigR+2Qg2j8HY4lsbtL
CUC1Z7EVSc9QYpFVeILcpUvkzBGVFfvRG5Cp04rOAuhBbXzgsGVEYxWC2FTx0wfp
nbkRv/IMi0swTX6uR4HFgSIsvWaxkEMRYtkmjvCmoFSrhbbGhNmMMGvqSChmmblA
lxX3zuygK28lAdyeXOGPOxeq+l+NVwgL71+Tz68sh6FCuHWbXGQTJJMlYXtvG+sY
JPUv3rrV1XVxVfOLekkRTsfJ+Oy484znpqMjkMGDzbagbLcBGlz8JgCXTYkRtNGd
rJUSiw7QODlUdytEHQ35EZ0ANhhg3kYerOokfsokWWMZSrBwDBSQt6iLXcoExpK9
Zqfxng85tkCDzChjd+y4K2axTSs/JgEvc7C9rYz29YQteMV4cZ7fx315QR3bEDN7
pXJORvFgUHbS3KsO+5AVbBCRfCawen4plvMgm2KcyYZSfJ6SSoEtQ/0DLYgDmw0N
JnOpyR0vm24xHEiyc0XSc4j8qo9fvuwu62nHQiOAw/twYU5ok+Ru/PZun5F03F7/
HkfHQnZYAB+CoNsBVYpLCKtN7G2o81WN/sI0k3WpJtw3h/xz06ivNVicza/a6shg
BGpqnwBIbJ4sElJ4Jn4OIb8HtUPYWIpBnR0eCSs4O7VUdFZxs+8CqBQfrZeeVC/J
4N4ek44d/OD3+wr7gqTGQYjQ5zwexG8lPP5VlPKNZUrLzCfUqXX8B+WaGPa/wzXu
Aq95RwM13M19NF2GOeK8bwZvMGaS4Y9C6w18IUjWAKUH+pxGipY9DlZ0vCttCs0m
GypYdiAmuVhokZny8plHk05iOfAAKRULBjKqySIUJtjFDEtpT1f6qna9xOrVNiop
eJFHK/j5TIqayTxXMaVmjyEv9mlMw9RWS9X7N0IQNr6ilYxaWsb80pEuJKbfQtpq
iHSbfIRvrBVZx4vliMGnDGMFL0/3sibEYmRwGNTNDE7n1xM4MuPx1hb2/8jKIeQW
iUdvd8pYHS/+8VvRk40AqUQC7YjHhGypv2WSGeiDEXSM0TGrjohgmK132We/WLZ7
vsU/TINJkC94sjQ+nmgx1RXLeOJgM9eC7SR9wz/MKjzfDAeCYC2ZjCE8ECwxNw/V
2gO7M8sMSJYWIHbSHPQm1Ec2oPWy89xKb1AbaFbydDcZYfvSZfqWB+Nq7fg5HXwJ
13CO2Ae5sLL8pWMrQ6xCwBl1P6Lk+JmctoDHrZ5pIRSC0HzROvONglnBlRgiAofG
t1+Eb4q0whl4vPdH+OWuBEYdNbW/erYEbzL1uk/ZKqBd8w9Uv+y2JK310tcXcBlJ
0C0Y0Y9rn2yxfvNSco3P0ggEwmSo9Jstrg7O2u+q7OZ8Dr6ekHmuuXg8q4jutgyG
EmB0OCyieGtV6687SJznbVZezP96rJlkBL4XQlk3qzsLxlLba1JolD8nr8CeKRRH
PMfrcA2MuEQo9bvhyq4l1BuOS8JpAR+a6DLkwMLk8HlJ23ahNSFAabh6cVPEcJhb
0X7HnH9LpVOOtieiZHa0USmfm+JdJyHAhkEolu4CNFILKM930oRGccN5F4NOdwh6
cktT1bmYy72zSLOOepruKJ0v9ys1SZhh7OWqqq1iad7+lLLvzg6fcPpuIbD4kE+s
57ZGzWXcJwbu2KVe8ibMpDlxYRisT2Pf6M7HQR2Spc6avCJnA8dUz4AMDrnoRTVh
bihttqczOt0SGtOYIQpA10bjEX7T9u/spSJAOyzNLuZs2L1Q54mVZ5EXdWVfVs6J
LtGsTdqnziTKMqDdTC4QP/62Rjw4ST66qgWankJE4hg9aIMPRG1j9SUAKpG0t2+c
hK04JTkGnLHe3wNrnYOM1GOUlp7/WqJPceoN0I+dW9/toTVH4U/0IECxZ5BhVKXm
scoGVBCbM3RPrmS94DtYwB0yWUJS7MegOR35EtilZZHyRkPCs66SgZWoeZRq8X21
CTT+weXzNrAkP5UQUgte7iGm6tYpjclEjsvfe8CAev7XV++GefPPxEKAuah8kxP1
9Vc5RrU12NoXwp640NzLwRe0uad6KS0ERy4WiLhhqa17Ni7eibyqFBdo/7dgyFjz
5sugpern+/vCaX8QKI2uW/Swi7I0CLbcCUnbFQTB7lu1dwdI0iKI9IDMDz4iZYa/
8A4CulygbSACPEH1wEHOydhopS5BguEedTNpgmgUgd+nHehR0gUuoa4hR6hp6g8H
dWkin+AMOFzaRiBasuXkNplOlXpjuo6Su46gWtyL1qml5JR/n7Y6ZVPGgFCXvZhT
/2J/G9JR+jbfA1iabKg0EABYlJIGtcJWearObeS2NAMQbhk4N7nm84A4/OcHcKxr
9K2aiSicNKduS/KclFlPBhpnA6GxbqY2arWDSnvia7so5rquXh/LKdlqCA4Bg8Zi
Y0ZHUERkNFZpVCelBbe2HSZRF8fng/BRTge2/qxr9lPFs13Th3F8Xh5fmsjdaDS+
J42DxHLb4ebDchw/JPRYlf7h/AzexcgEYCLRjtlNCh+eTxOvybI9vQ6DrL0ciyWX
0IBD8YlZ8lfRuRM8xxerATtZ4n11KTowbZBFH85hZ1zvLsJlEI26fCuHUqTfGreF
yFD1234hZnsK4oyoESluWngPNCYZMhsiAcd7ltmCyIh8ixvRHTlvMeAhlokkvGPt
8TtcLhzqXWkUn3JuA7mjGq6YOxLCR9v+nD80l0KFr/EJgKW9Kjpx6D/EGz+QlNBf
IzM3Uagd9Zm2ZX4FTeWgawXlMzChJDw4KazVl3+Zw90PqjIG/HVnmVn5UV/aNYGZ
DthY/SY1wnMhvJNklg4/xY4m4pvi81jijFBhDigxuusE4RLnKbW7oKND7YwMwsJh
sxZ8WJelKpjCsvp+6DA9nkd0mvMtkXP//Mm4iBqT53CcQ3h2GI3KC0t8fOdII0GY
a6KMia5tPexuQGxKB3HjubuoMyH9EA+DLK5MtASNmFkk49v/h/SbMh0jluQQNrLb
ZS0lDD6VQ33YIXqxSxoflNwRfznG2nq+j7sTled78oQ0npXFaFrxIznZlUsemOz0
ejs628VTclWWYFffqTp8AkIVHAS9NOMZqaQ2zojwsaZdVn+Tgobu8E9StdzSfcAY
XUDnVl4ZY6Vtfhj5D7aFIvccVLDH40hGipM8CCBP95u5/XnvKql8p6Itdq8M52bK
+F7uyGewxlGYasf2hwvsTFJoOsIdLFv4ku+dQ+u4ZHtEcFVsccrbkKaYtYyTHNRj
nk29S+bbdhE8M7oFJxAicQhJ6qo56RuUiMfLxMn683nIYh4YvGVTnHcHn5Qek6Gq
aj6R0LqiPdoGUjQOUliycB+7qZoLDErMgqBY/cFqhUSzXmMUgUPmvfougzK1veA4
9fwiow71pQhEaglGutvqhrQx6gEc65G7/XtYKu2ViWhFmMHsOb0DyUu8Kuoz/I9Q
MR365hMVCMGOX2245HHbQUvjsjsafXGir2fUQJX5hGHVlMKKgPKRaN7vuoZX1kHU
D0krBMXXY65E12erWnHweoxXMLnP0jWaCRDgG9ChDbLpeCopjSO92IuSjEnEhuNz
5mCdazmQiZ5KWeSG1SAgH0DeORNCRPpFxPDLlVjaoPMU+yu86sUVE4qwvc2uZ0Ui
Hv/bDmDQw8frqXS62oW8gmbvST9dTAH3PVyiiKRv03FLo3uKc0MSZF72KMDN2/WT
58thVnV/BYkaEW4Azynnc4XypDMYLz8l6pn88i9+a+4uE2k/fM1GOE49JNc7P/ZQ
uWDIppmSAXdB9hIXNJ+lkPZt/f0jE9xjp8bIBeBkspXGVgkUzhxjOgwFnRVN5xEX
dOshPsIFZwf4qJe6lGISLsMmHn2ffD8FnGUgIZV3fkPM+0h4BOUupHznTmoXAyUa
O3tMOHdwhOeEWgJKV18uPojcspY4CtrQw3bLjI3VAf0ar3iOD9UgamgIVfkEjyfA
+KNnD/lx1eiM/TvaJ4rlIKUta1Y92C61XUICu8oZHeRZ/SasC3YDyZ4dB1xyLBNA
57Q1vAlckPWSgg1khSDhPnj1f9Vxce2bfHvBTNnIoFKbuDJtefCvZGgYtI4heDXv
SG1OD8BHmbbReHv4GqFLZ+L8IjDtxsa+ngQfemaa6Ufb5qh1IX7P2Md+DO4RPHwv
BeX/VjehCZzcINtTdkQhAhuds28e/R2Hzc3gB8vVUWDTxLmmL/wR8NBVRDPB/T7/
DB4U3zbNwVSnBrF83XowcqhjS7eiB0Wc1jqiQYPvxTdO6tQCSERomg8CuaJ1KIc+
st8MEGmkuwum5SVpcQ3nyTgGIPH/F1y6p+OkblISDRjnF8XIOCm36OonOwQAB+hE
6LbxTZT5dJQrTRs9+njpDCv8UjBzZGpJTglyY5Vhon5LRZmeuQVq/giijLO06Z8f
+kk7b89CPgvWVQznjOcy+taeX1eREGJ/HYgcuz0LYJ1bvKaaJULE7u4dQ3ls5FRY
Cgj1GhPFEVJmcKcVxLJFIcd1hLHcZ62AQcyjsJGqAFNe2A5gi4nBynRMHvfDgucB
F88D2cULcRn+DTkfbdi4TJ8tnVrEDKzH8e5iKf7O9YIMMEn1A24bsTTG7ohAlKPR
8pbg2Th6BW1L5rL7Qg9yEmDM6WxpBui7DHaEuoKteX2FwNg0xQNJx0I8wzyiRUyW
d7KohijSpTuL9SeTx/uwEszmRMxc03PXSAg3gMoHSMHpbIgPrrZvyARF3nvdsKVA
xTuUptqW7pIR3gmr0/1AEfTri3e/kJ11E0b0QXwK2l/Dc6Kjg7uvb3KdMb17qIr+
8FR+FAjQB/6eI13KvqBuP87sQIuNxNjK4Lel6f2iP3YKWjdYgCPLto0K38zj5pjb
IIxKV0p/9InViS1QfOpVxSgMUzcXyeCaVu/gNu7MzdOUS6qQKXm5fvM84hUqvBaP
oHvanFl/Xqr/WS3az9nlLd4bAoUjubCQ692R5/X21tQ9KDXpbyMtRc9nXWN4fQfj
J3pTwgR9s72DS2/emtPKrc+/yrMYvuoUH8tlMaX5P6daU51whyDVemkq+Ryszh4Z
4DkVq+lB90hnh6xbFHcOwzyZx1BsHI9wuMG6hPsJp6bD8O4C/ulICRA8a91Q2t1y
XWHpKRkjsxPyZCAzOGc9bD5b4tImALoZySGgSKF3ZBOQ54FZQTPVXjPPCyBlaTrz
MBCHlwCf3Tw0BJz/CSkqtxpvM7fp69Ju6+zx23lP0soTKtcT2Gi21ZhLg0/VPJ06
m7Fe0DqdStkbcVrZKOyDLiY4VuIVIE1ep7M/s8qZ3Ml2et1RuBo8A8V6EZ7D7ilQ
2HnSNm70NOHLIsYAdGaK/VCV2fayWmVIwormSrJBTwqduQ/9tyGXf5nuXH/03W1W
4APsoBuOYbjfPmP4PBnlNNh2ZvRpP8ac7VAN1uAuLyGF1k4e5Eka64dNSRyr+T/I
Zknllf2RXa7YDrvmuppOstAyn4tlMhALJMS2szNblLf3aKBv0bnfN53GpqJfgDnN
BG4VxCLJCUQ1IVIjRhUAcUZfuAZNmTrZbLk7UpFW3M4iqisoM1eXbqy7KN/snh3H
b0F7W7X1IacuKpZbTgmjj6MzqiRD6GVZxfpdFFFdRkcFy2ynkFqbH8veJOW/8pnM
fgH8YgQWxjgxLQhtBei0G5pY3/mCJLdE6UMWLGSaORYcehdty5stnEuj9OMnH7aU
Hsv4tmrWXM6fcLIeEn1fh2aXqyLdfuyOSK6obPK2wL9NxEbllw0zM0tTHnKwNV+F
ZsJrvdNlYFxdYtYdvXPOd5pe3hMlCtb7hro50YA7tysmKujdopS5pB7Mcatg5Ath
gCmxmgtWcvULxwXFcp3J+1rWKM5KlMB7LWpry4REIsuBaQmF1lrer4nTgOtjb/Va
o3bkfw1PbPHJtg5RNL9LwooSh3jR2mxWegZLAFEQq5TP8Ge8de+cVskPQJyaqW97
GeXUlfApIV8va6tOCZgWUfzwfCtk8NaaG4aQJenDwc0SpzSNI3scMEHfiZclu58E
EtVCdlFaQONFzZVupFqI2jvlmdM6UMtIR+f9Ne0nZYYiERVM9nWjqovyrQKRoB55
CpEWlZ7hsKQgbTPLTnMHwg/FAzINDpTDfnclZuebsw8pVzm5SCJDe678x1JtOWDh
zUqI5JNjkDjNtRldAy/NwQcsQisqWITOheUyl0Jy+FWnzprKR1kyhdYl2wsfmQZp
vRGwOwPsp5zUreFbXCgWwk0XeCeemzHOnAUPnURM715UWYjM4XeZam2kGh3BJL1P
qJ+fgENnMDrb5AUuHk2AAdXNM2RRK9J7vxsIdgpfwGhtrHRrLMS1XNPdn+V0PW7o
klQSrUqP2qpVQNla79JuUfH/vuMS8/8S1tT2b5YBvCdVNJgU1JS2wOqIVVweIydD
QmW9Npgf1NIiNeh00ezXdN+01CicZZUdA/htOOqjrUaLScDjceWTsG5kcn24kEKk
XEjR+KGIzr5wVFXCpvxgRSa8aZnQYxCTgqqptv+7vn2w+J127qe15HziqXwPzZsC
SU5/LOsb3uheNCS36TvxmOtv1CXHoebVKkk8oBA+Vaugmur6uHbhARiLcnsxdw/P
7+EQEy4gTrDrLwCiVBfrnl+RdDX3VNMSTiN+n+bVAiWvOfnMDS7QAMM1eGCK68qc
DjKu2Ra5aF97xx/DckNQU4au+QAI97u/JcF5ijHAMwDpegEShq9LjIlAbU9LL7VU
E4+GAzKDCYJH3GZHkaPuKImoYedK148enSm1jplktLhQN8loy9hi/SmtLvWX7TV/
4CFQBIKdHoksx+uVsssnTuFZZoTmfe7XAGWNmPlSXzHT2qSap2H4bLfAVR1cwsib
r2+ARZ62H9CZt8YgrkKK03otov5Mb2MbM3Ihmlg5al6/sxs6x3EQBNTwBuhpHi19
PHyffqse9IgxJGci9rWd8evpjVT8w8dmLRmyo8mq2XpyRtGdwY84GxeNn5Z6EZDq
nlsZ6HlfOSW8RBJ2eHapdgUwfm4oIL5VrJaf4KaaOLoiT3LjhDGL33BMId24+0Ha
luEBzOhYs0RclLHOTWrPnVjq7UyKsUnnLCIHyHjh4R67rcFrmZY+rAIrsfqJj3wh
LbZvVE3CNTTjj2BjEbyONwRI1hPIrbY7hlD1SYv9xnAzrrzDYdONsd69cARZUr8/
nOk5ybBAqAAZXn2/T+2ayTpTFW11a7iOjw7KVfBYXviaGav019dPmLaavtar5QUX
AAcGT0rIE/NDcR2zKXl/MDlERJjlGCxbXaBDCapqw5rx2h6m/xwxktkxrzqVeFfc
D7kGrnDf9GfBdiz/YDBFOgzkXKgbVPjC37jKmj20KL/Vt10kykTdMOlE9IcADa8o
NScxukr/zD8hHpDsYer2pD71qs8RgJcxZI6Ce0z/Os26LPwBQB86JmGCzd/8dXS/
Hg/k+d7E96d4Ax8XYVuTmZxfSuuKsZy0DC29a/JCl11729LuLLYUf85M0Z6K3+hV
webeV8MXXvgHHvlNjdFQMYNdAdytMYXTsd0KxEJhpb6NDjFmzWB8XY829GemvplE
2ZoC58GVbIJCgsvPrilcuZ/vK+wDw1Q0YFqSbDPxJjEhY+oGTTKfvLzL8xsFwrBX
7cOqsYoKpgyvlvHHXh0ga2yPZnqJV/BcI8cjXggCatEuOXzLdm4ACqupiOqYgxUE
Y8dE+Qmm9ffwLsWPZtPbJj4CQ66UmpX7Xz0Wpbih8RTejZ1nzqGtyD30PnBag5uu
jTBeorXYqnmktTleZ877UGxiN7IoTU2PJjRrV7vbCgZxnRGLDMvEqXhGFdq4LE8W
xx4e9Gqu7Llmp8C3mQyB885PqcCnJH6jAk6VM67uOglH1B8bQ/tCZ0g+jUiEM95y
unjZrL86RfyTyENqixB9aNl/bRA1siE6ib2to/d87gEkZXrSioZhUmo6MAD3tprD
+uTz05vkd2k5hCaijTAqiuXE1X393MeK/z3JSMh+2GO7d76N6mKiYvpYLlK8bJYY
GEN6tuwCPVUv3nHnceGyD0ipbHEKIWaHnDbBdkE006vqdA2WxikLY6L78S5gsmma
U2UYCvSY2swGLxtNLWg8xBObYzYV5DlrnRJO7iF9TnAPqI6iBobNSMa8g8LZqE4S
xX4UzVrI/y1uEWABHuYc3AkLGHp1QWLhe/7MgPrgsgr9evCzlycFCsK3NI0FWaDm
IyVx0/PgqqanJpgk0BGatqLGmmE5qRvn0C5DDdFccGLnq06RughexgxMyTNI6Nxx
eiEx7wO60TY9i226oyrVgOr4NLJigo+Y0MYDX958IC01lmjQbYUB8Ix7SLOZYlEP
nKAtyUeSMdBKa6A8gMcs95ze8bVIoEQWxPiO1lmzSStCAR2AJSoD0hKSlKsAWKcx
/NV+sv/vn6MaQ5v9bVB9KArFQe+QYt5kEUdvijQUMK4pUTt6xE7DRBr+etZ1c4he
Rwsxm0R3p01gUzTE1P0ljht+xPZMLDVu/GOeLEQceK9OdoC3xKAnzObsI3W53B3A
1XieSFHuOOZEgq7KOK2Rgj49hxfM1Oc+ncvBvSExT6hayvAdmMTqtuELH3mOS8Ua
n8C0N6JnBDEpHhLd+6wYRkb03ZcwHXQgWI8SmbESlY2vmXGA2VcbQdwFg0oe/YT+
vH51CoevE/npusdAcxpsZtjMke6j6qfwrLhoonPXgAytAwksIlGquXl04c7YUbpO
BzxRYo4d2FqDEWzSvwngsfNcbluwfhQw/sY1yfEwjAONRBnt8+jtzAcuUDQfrspd
ieGJFdTnPXMOf/8FX6oPwc0KmakAODIdJPELLf9+Qv4kgm8687svCdwEXM60Q/5e
uM+vr+c/T35tyJcIPJO3P/eAXYeEm7qni1ppAz6HnVQ3C61GOq6soGBKL1JiEd3W
p9iDK5JJGL1JKIZFdshCMt2JhD8JO11hRW3PKm1OmSRXYljk+0H2IMshV4cDHdQ6
pV2n+fWhpVVT3s9qkneukCu9QMPUHTUG70LEeosTFeokVElsHW3b/aiLNBL4H7t4
O4eyguoqGKwDhKzlNOewXyLfmvO9Xt1c2XcE2S79cPKXaZYxCa6Hk8KfTr70j9Bc
oJ7nJzDHqYfNHNLtOcuC9Xln5+o58HnwYv6d/gV5g/fvys2hz4zrUCROkQx8BNp2
nV4amiZFm4z01wRH2Y13BccqPC38ZLqhYBzb1xtbIvAghssKBTpSNAcdw5rHPCZq
ILJQdp2g4SamqxAdMZHrs+c4b9fZ50uhFIllDoLXQ93GP5rXTDMq7dvxoPsfNBmU
hBOM6RSNoOJgw2NldYWYlULcfTBCqXRgQJwEtvnl1Pj2pT2LMQXG8QS05l/PNZIn
1FbmsZH3U7eKaLhFGDNSKdzQ4PhsYLUHzNEy8lPgd2RnWhaDQtqc3K1wTdncpyI7
VVqNZ9d6uJCNpaG5lpc5QtqJTEvWLo+tYElK6I9QbzIFf9opUkWnEUp1ZigkBJ9N
9/QHTzGAYda4PagWEIjNiHy502ZKf6TchiDJYj/PxT3OA/zIbAu+6IZfVVzDMwvc
EwAKtoeiNe9rMZBlTp+V08XXHQL774b484pGg2adblcwvEe4FohnQlYh2Dwjrf7x
SidpqNKozJUfPEUdHUSLUoPrfQgybn0XyzSI1dU2QyGLL2axBFpwNfbEYwqDC7TI
lC6ceWnQ4L44OBpQdES6H6DORihiAdqCK5KkgiD6AwxmRIR3YQO/933pFrQzOozy
oXYaFqk4e+o4HtfOHW1jf8pXKlnspluAG5BjuJIlG3of9nCzLd8IzxfFpDfmdadv
NhwNY2KtJWWMjRg5dzZAesmYY2yRmIqadlM9VkhyNn9nCduseYl/IySI6p1C+NAa
jTlUoodcyMPC0vsaUyYPzbbd/6X0aOhQkDLoInWgulVJFwbwtvZByXBVwgVr4ipY
WG02ZKala6zy5CItxHxwUb3bADfP+3M3Of88KiTIEheBXBBEW9qS9CafRbHSoaR1
Y2WKXELKfR9jWX/+X3j+em3QqK2HDC5yqzGVn2vuApnxWquj0fNH3h/fo4ORCEF+
rode3+zk5sXBQn00j65w7WgkvulDlb1f2Dm+jfoExfAErp5EQLPXs0W1EW8IMoPV
OisnwDntGuxKVjh1/QT3ZB0PLZOuk38Q7wT/nplWpb7cBY3Fq8Yo5OcPGzqVSnde
a/uSkl3qqdpu4b4SLqE+RbaLyhayxoXyx2anpcc3RS1bvidt7QBDvAbQthTaAkUM
j6lsrMeEbHkkt6kJKQhu6sM+lNhV42lnGH0ROkP02z8SJC7WtTphBGiS/z2xwzGI
rkcS3xhkO77Fa1/ubo04GS0qQaDftvv3VtgwuXk8vEBCiTbL4bOVpCjzEDVuJmsB
0rhssTgqV1RLE0gVCETb6I6ahK0V1JuEgDoUP3wbR1y7PfETEbG+hVuyXBOTW72k
j3bM8aZnwtXzb+hOfYrsA0RXOgMf2dG3rA9xbjvNGdwgN4X3Td1UJoyLLJTiTbxQ
LcDaLh/UuqTxvKv6qlSLpY8kR8ZE52zM4heXyd3yS1GtGTV68wfelnts6Zeroeah
cYwW/mxcqBMszjdHPkAsWHoxPc3gtUOBOa4TvYy1XKiyQflGWC9qdGD2C7oeZWrY
XSxnCwDFIVSjBfCl5PIbMRiUTjN2kIhibcVxBh5TFNmfHMnI/J9D4QTxvUzUNM1B
2QMju2s9PM6f2GTJojLNrsKJwl0XpQAvO6Km2OOuGMyqd7/CR2+LFiKGkO8X4j/y
mDSElQId01NuzVqo4ACVzItOFEprIo4L0uNSOSc7JYU7fXLkueKmh1l1EKG2ZjOV
/u30C3tVya40j+WeWRS5erlcFMS2nL2e5E/TNQibzLi/HdAwyQZBQddYfrIq5jNQ
CyEru4FxAP1eMO5gVluYylgkFG2gg18DFVnIkXLQcRRQXtN0vqXPlWotziMGs0Gf
scNYKibB/MKruu+hy10Yq0OzHZgAfcyI10U/XS0WtiddHOkeLGGEJ/s7YTfJkWjY
aOfDIJqN7n6fyfTQ6pMTQjGDZUpPNM2bx3Ke2kjpCiWQhXds33MKQOV4N80/b3WW
xNjB/y9W2dgPKurue5VAsoYXLVS20z83213+PBtjpc0+g1izksHlm2dKONEFeq6d
zpJnNvJnR2yjNHWlOSmV6VmWT1Psn3AQ75W43G8OdHMwrKCNPSKP27Uku/0rnswe
ouKSO1uu3gOtJqjUsb0veDnW6NTtVXYdj8jT+gB/OTWqdTnymuieYxS46Sz8ffH3
KGzEdRDooxybdZW97IPCuCjO5waqfpvJaugdGGeFEuslvRE6rnwN3iadZWeImm4Q
S1GnKu/WcgvchO1IbwEH7g2vsU7v50pPNJG7KVD6kBd6BoXEalHnLbV1qc8y/NiE
zv/pyYyXqnqnJm8Qta57XLNNJlpekCRrO0HSXehmOLHVlyFMZl4l1mxvzfzlLUgt
ithCSeq02g2vNPB28bZL27TLJNN40LRLS6SopQQbW+4y/gd6ff1U5GmfAauOiGDs
3VS+H+5Rg9F1T+kh/2QZm5Cv4Sc2nRYA3/iTD+LAIPefrB4+QvmLnNOJvDFGRkNn
m27gZkzSAl93gK5MiIZRgcW3qkbalcZ64tRH+xklhVwWlIszYhrkjY4pubpHpV5q
Si4Lii2U0vlfd9b0C4p7XhHcTqwS2qaYrZ1BjWz+vD1WhqsK/QMei2bEJ06cpAox
xPIyaciWqQ4dfHM6g4RkUjShe9bCQ4Sh/dTqFW8eBzEf0KJPCbV5tlYbqYS5tNF1
KhMqxm2ZEy+sve5FYh3qNi8kzendIKiAXYkGoGLW8rS9W7D12GwPY6jyTcPK9WYe
UvuLViN9f4wMWqLHSRVVr6sWJ7I2Y2ya50eolH3LKFiS54fe3sJc/mq9J2gjWQE9
d3w9W4fP4s2uGJ+lh7Np6BS6KROINCYQjZxilRhTRrdAZ17FRfJMaEy0bGDHMF1v
TQlTjH++VgX47bofq6PegtZEaCIV0rj6B63kGhJwEq64wa3KUdLg/QaUMG39lv2m
DzKV/ePfdY4LY9OkzENQDxyMYO50fFpzlCF/WygXRasW+K/pigWuXjvEg3p10wkZ
1yUMXXkgnfCKRtPU9IJobkFKJ9irrBN7A8YBh7nJupPXo2GTy5sjRb392IM0flq7
11B2TdJOEYQ2upW2NqKqjDhzTb11cFgbAWjN+Mb7BBYDq0UBDe0v1vwVw4kSFLVT
d2ukzEBTD60asp2NjK8sV9Ejh4LUPKv30Q3uIKY4yJxymwjQ3slrtRAopMQiDUEy
+j6yDd/HvwgoU/JPNDa/CdoOtfKgqkk5LsSMCDQwu7Q9XcFYaSB76igSNfCt/eH9
tSx9/Kcjvp6s4m4tCpn85dTpZKtJMBP5z2UZM+76cEskKFdkXAbWt/CpSamkmby4
yhLkz6Z0qMeYdFA2XAcJN7AHkZGcziqdWQIHwS7EdezfMoVrXiGxCzBv00T3iDOs
nN8gJzbsyQC2rgYmLy06NmWcgKF1Wquk1J055mPb3KoVutGxoK62zfhOiFIyzer6
oT+TeOcbtSnlYiNcpS6uapwTTKdWBuN1q5E11GVJjJGWz5K2C4Vur8ntnhE0aYdl
tzbBrZLd2nffABLWyDLilLnON6rXDtYCoSd5aKdrQpdUEbXjzS9vQS7niGhbXk78
fqOJh0h8Z7sLvjQ6aA8BywxDOT0L7JKjMRwujNJxPYnVJerHR4mNTqtN/o5C9TLT
UaJcCVUnCrfBpiIdkZlrkNntQ/+9/OlSi2t6qnmCUSegA9jmjOl0MlATgNfiHkzF
lXz1Ugp/J4vOpR83dmZfpaYgt6tLj+NwKEDir6BVizKrHO0/YdBMl5inwqc/nO18
uLmdVch0MPdj7EGdptm17iZEtw8FLaTZbTFW38Gb6xD7cNuRlpDyPG5Y6WgL5gs9
LQLX8bO0bss8lDKuxY1aIf2kcoHaAFF+wQHtuNuuXVYCdEjIGLBkn2jBj9cbEHWo
8xQBGerxbVa6HZo36TDPF6VLVg+MMCsg3SwB5CBQtIqzMfb2BIthLh3+kGdbS1OD
uu2XT2Qgo1cZO6Y521NnRr5SNpi3jEQ/iWFvLmHgrMh/rDx49w70VVAZEZOZqwjr
GBfjCRwC8JAEiImvw+yknAcZgJloPIVdTK0AMgGY7DEFcwnUul86Y73/SOTYIkpl
4XDh5yZguGIjSAIxcTniP8cBHEpS/qTgRKIaF+vuYz53yws8IM5TIe8RMkR3CKz+
EcRstf2ckwwZZ/L3oPVfj8L6Ua5cKhXX2hFI+UUsDILJ8kIqzm7aq43Sxj84yFWM
Bcg949V7+Si2jyIsBpnnfwvBzXjAZkaM+QKSXpZQ0PbkF2Ja8pJL1hQ4I4RcNsYj
MDDCLdjoGS1n7g1tgi61o1leOIIwUHXX90GJJwvMPTQRCJnKp3Cxnrm+19eH10aO
22R3oRNoea+Ztf5m45JPYg1gg1yHfBXs+feleBFDcZR1S3Ful5pS8RHfyLg+2XJJ
AfhOgNzxSnaeecqf29NzJu9sWUWZL/FTqP9/DCuJ+ti1w/tp9Bc9wEVEnEyP0+tP
Nv/ol4F/mVRfDGhtKebDuB3UV/aMdDEvINCdRWoPt+oFQJfC2GO0VEz+iVa3RhJl
sdS3cI9a4IsEwM+n86zBkBPRw0WTY96nAXyj/n2+ckIXbKvp6sc6K4kL1ur+6tTy
qvJA0g8eOQQafmSjR0jfBy5DCJJk2QVoy1XLQcP1Lt1de0BgS+0PQCsnyZadtqs+
n0JAme4zRlkjZUGk2U/fiGq7+tQgAupwE7AoXvVcsjHhiVymWhZ+Z9UuHbJQ3jXh
gyZiMAU5Bbjm2y4JCAhJZxSAx1Oa4dS1NK9RQSxOnbEA09GxLtmLGIHASlXrChN1
OyPZ/XmAQHVxduOOkMzzwZNN3GwAsNokNi9T8pk7XcTsxYVLLwVx+euy/t3OV35D
E5eS9Zalg3KsuwsAgD2vs0ki5QmLZKa2CdVUMQ4d011jzY/OD19rNLQsqwU+Fffp
56wciE5BHR/Z4k8HxQ5lb0jhSsrcKZdbFNoMlNOfbXCd9TaN95VdRVO6ZKY8mSoC
PtpqCxAfJ8rkHvtxUTf4HHrjlWMr6HSHtN51FMR5seWwPBsEUX3Qr7DesBJbkBXu
QvuWgEuOQpVyIyG/LGlKkoCAqqhyfENzUO+pHHeVLPe6hsgM02hnf6Biqfl40dkp
7NOGu4DMht36iGbIDAgR0Nbi71oSmGxnAV9lWyjJ30j07XT2OFc9NFibhgP48RSW
QOJ7GAdhEpMqaXHoUbrdrUarbQbE0jfLOFizwG8n1dK3qvpHkw3/MqsLvjIQLZZ5
aqNphdLVguB19hQ/LAwo66T551fFiUhGQYy5yKkZIAzcxUqLU9O6Uxou50bZ3Jz7
7yuTb/C3xepaVc3JeJ4BcWeL6cm+dswKhtrv1PZpVv/CDIX2csFwq5ed7PSVYYBB
gmlT6rcYE30KpyQpczm+rdM1c43ARdAIpG/dqEMeQyOkYsXoUijEnJ0c9CzwhR9C
6BkHGtNILAaPcu3qdggI6KkIuuiZqzYbPaaBv5pJ9z6Vzm+E6bw+kWn8lbK2xcTj
NqF77ZdJ/J94+qUhIHCUzRoyL4cNYdSPfliPEMqXgs+Q1uuwWzvNpoJ1EXGMpB1r
7OwmDH8OmlWYgoMLGnGJsGFZ50kwJphyO12zWjCWsP7OXDM4Nq09PHPLnxPXWA5A
N0UgvzH2WZ25rQN8n/dWrkXUUcxChsnPg6k68ofXFdJFwpuJvX38XJ2ekK95Haiz
lXT4hR1oPiHVmlwlbKEOzo19wAiSvZJbqA5PKHFsD4Yp30KuU5KAYcUGyd0TGg6W
g0L52wuc25CgxEsikfLXyJ7tRpBz9XgX3VPOJDSY2LcSrqE6d4MH8DhG/lf9BTC9
qde8VLCHfVeQhEQlxmIZHXHUH8GFNFjWtgR40LpnCPv1UEUIaWjahc9qKPOMEigV
vesobM2XYP6QN+4TNPoQRcdNGJoGXT7Nwyc8Q1B6x0LfgQ+i5vT2iG6FWOjT7V1m
Y1iOUiY3iPqQfuNLtJBWTIqJ2NOfLmSCgncEi2+X78uoV7bo8SSXlxPae4dGqGkk
RSBI1lyFr+fWjvN1jE64FTcbmKFFhRmqx8ohWQqc4Bg6C31M2/pBPc52tL9RkVP1
2xHjSaBuSoTcBK/YQjxSWE/J0sSN671xJgpv0InSIlZRcXMbaP9LGmdd10Y/J5Bh
yWEct5Cc4QZOab3Y2EWLLyOGRfFnyvtVofmFziA96Gr6l+2aszYASaFU6vPcM+wS
dE+Jsk4ctaEhAJmkE2XPjL9mV8eIICBbQY18ihNLpKMSpkFDBptRx1+w3OrFwp6L
8DsnAmtZxdqzTKoCG40RdVWgv40e1b6xm+UIMzBGxeXw40x+vh8mdZL8Xt+VE/5E
8RIx+EXAlGvOoCmulzILcRSlE+0CS6cOy8/60D27CMzd+K5j1d1njfzLedhZXDea
k6qUq4/SwE70TBJd624T/iAvda8vjG1yMWDvti0QfpUQ2Aatrga0vLwy7Qal/mI2
swFJ+b2KaixSpOJmy0MGIHecdn2eHqgk56hVSSKrpCmdk2Y4AALYE+8+Qxzh8pTy
0rO+xbkmAEhhPRgI1UH4tS3a5e7PJr3tDVYyyDO/VEs0CwyuJu+FgYd/GqUSXJkT
RN1mIqC/3pIK2zB2dGMGtPppKp+azon39JW81tkA23SUO9UKJrDSUa+3QIlucxZg
JwD1vQLrbpQzoC83SqTVOTV2oH/5OBvz2CKkQVzSrT1oDivVmSnznVODoqieCfln
OuGEeHPYUv109M3rszJ/gEkc+44t6QzsQqNq8Zv/dZoN06TZkl1WW6hcxnc/YtOV
h4diT8XHZYpohbGeJUhszLiJuN0e2HTYWAIT71z5iMfO4UDNSL9j4+sQClDaQdhH
Uw9MdH51eSrfNipguJMBrkDT49545E41oD2HbIXJKAC7m/65uOeUOWyTFm1rdQ//
9uqGIPHk6QfRtp+GhZO8VAN/J87a2xUQnNUjHHkm42vF0Cat8VLK8r0q/Y2wvNoX
UELZIPrnZRg5tEROJhP67jPAStfYP1DnS2eyuvuJHagJowTq5wTCkkWkRc4P37s2
ulxNevM1Yf93jonb4FNawVahdtWOvQt0WPU3FoBYQB/z4jw7pCv/1TUgzcu5KIYX
P4XTF2rHsDU5rlCSr4pZ+s0wweR4iRfAIK/BUloLs+KYtxbOI1+vGe1JExKe5COi
Yp0O8VJf7pBlWqv5lO6C5RtcpY81fTiFfPl6ezzBHGjgbOgsB9M4G7Xx1GkeAWO3
MJsXRoT4K2hUBWDEUbC4EbvaTDddlGVHGfmuADrmuXM+LFARlr6aFWZ9g8rD3Bry
p4tyX8y8WlJ12G/H3+xXoompmUbew6rziRkkdKZ0RnUTBQ8yANdzREnROfW8Ytfo
s9R7UZjWQ56f1rVa+ZRkooS2hOS8iAvBTARW6Z5AGT8a1xJ0mw6erg4xAhgpF+yV
39SIj4Wsh0LbotxrUAblTbNPUqhcgYaWG0iCzj9NDoGkQkQlXCd4irkzd6DPXxek
zzcS0xOCYKeFqXKgCf4PW8NxWEoxd8buRwDKtt21+uJVlTdfvMN/g8zM8dh7rdcz
rXfIvDhF98ur1SFZ3KHlW+GcPIDV2FqAeTG86vSLheMtM6CUhb6SrREH0KhLOLd7
4AEEsiw3pfuxgjByDmtsLs+V2am/8yVtZUxfkgmAeoKVAtsBiLyf98nLx/Ko7RBY
V50LDew2Klnz5L+wYcyuEorueWW6yxE7GhPc3DoJItWH4RTS8dgPKFa9DQ0aXEzo
QZlEsB8YKn9vAX5Jw8xWMVQokHhI0PnPEUdrilwpeAJYap2ZMbpE5QixIma9YgEc
j5jarKNWa3pAPshx5Q8NSmINeHLUNuBjrqYkfw8MQwzJeXu8s7l81XiYEsi9amUj
VUUhS/aIZPl5pXhyKI2SNPKUCg0aWI8d6cHXNKcFE7OaG6rtU4dh8Ld5H1DYClSd
DrocCWIQ9q8/lSP4Z4ifn5jlcDVKmDGhRsIBPxpaQwF0wEDqvW6Frenp3RUUeGch
lW5LEa1/mtetuTNajnKDZpCe7MtUK+qW3aGcJpQ12YkkPnIUKY/MswkrXL8NMj/c
fH9FUz4h/jMrecFZ+038aUd+8lM8RjC+HpYt2rHWW3hBLQr24aUtdUrASInVdlt9
ae5KfK73hi08DsD8DcCT2C0n6hg9VJRsS8eAr3yFd1Hg1LxAqBLTadyhKRW2Ke2r
D7rUzo/4mFDkbnBthLT0G3IJparmGL9pA4Kwmxf2CE384v9HOVeepePGsKYESkZl
x7JWd/I2vF4Anp0weSCrA2vfbyVmN0dhQMcmgGsxZvviq9GPR+tjXvkcr+xvrvmk
oBXxuxTaNDcnrCVvzMR2vM19ItAjT0mLzrspqMjsqPYkXLpp8H32n6600Hx8f4Lu
CTuboaxAtAxrtdiP4h5PM6UpmYahEjAFK0QbDEpS7OYMSxinkspsfZmvMorvmpGJ
S3/2/tgVzFMrw+yRlvlC1ZvuYBv2p5p8wjlk1gRAMGugN11xm/ZCEi955/wAg4ZN
yeium2zLEbw25+IpKI2ANiPMeJV5ZYN5eXUTOqWcuwakqLHbYcetRe9OMrCnRj17
ZgXo+sROkFfUp2TDkQa1RoZHXXIIludxGqw0JE9QDWbSiB2feN0kwUKzqoJqpOJz
+v4JQpzO3EYGxa2GDgHO4MbVcEBgIhBmkJa/WkajJb3LKcpmWJd0vYvuK23gHQMb
bUF4aH1LBJIo+wLuVBmG+nJHAb/UyOy+L7fQ1LdQN1O18bpVlValzXTWddxC2UVj
tVePZl08x/L9XSXq07UidtfLWZpIvgHokxFZgv4GdYtFjdCzRRBuH0L1zzYnVCxB
fCh7ZWhatAFjCnJSnNW6BFQjag5kMjmcRxvt+hSkHKb7S57R92sOAViPL2LGqbES
viN0VUEUFa69cG3H/oTCsmgBDWXJWLXNoFo/ORo1HIM/zcniXY6fgNVageKXsD+r
/+7BwuW9jivZ4hYNDWGwGMDDGCBGjpViehhWmkS+hML5WL7e3c0hM2/lH3oxla+f
fTZCNPftE6FlK/h5YeVmOcFYWSEAr6pCWqYEj/RVNHsfSzI20C6gGTZhPaJSi/6f
TgoTNgbhk+8WnG92QllkXysYZliz4UK7sMCSYaJngF+Vfs07WAUemfBx5Gxz+0xk
fJBuQOMaFVkY9KZlcDiN8o3R2DSTchSCvv5py2ATShAsJHUi4JKqKolCbgeejgHM
v9HSvJ5FcVsooSHVdYtl3F2VDUL+VGSuegq2r5zpYiSRuS88Viz+tdpadZDvjkme
gz6FdJfHSVP1tiSKJlWZu3sfZfeWb1m55tUoEoVEGbIXbNELj8PrPdiwTMIY+0IM
STq8DnvsjADCPH9gQQcyLV0Ev04NDgE8lfZrDQPnoWsThR51RamBohn5601nuisy
J1C6j0pttuYmARKoaZ2VHcGcMFF5FxPEyI7sFBz7Fq4yzJsSBjXcoF+iB1RGgu29
tl7blnHXMiNbn1mpgtjLXv4EbAnZT7Xep19od81CMN1841T+/P27mtIqXUP7JVMX
EnoxI6TuYnQM9Yy6EAgEOWdgnc4BB6kM0BJZhnXTX5E8R0+ZdpxTxeaLsP30KPB0
Mnvi+caEpdr4hvsj2inwDH9SUq9wKTq3CBRVYZfUGf1vXlJL237LnsjWGouYWk7J
qNRkb7wpXHV+pKM/sWDjFYkEgeDan6/vP7Lic3DiNzCiY/aYbyt7kuZc+4xOt8w8
VVhEtCrfcPlC8UWI9+0aMWA9TG/0vmiarNq2pYmzFH2WiBsFjBqnlq5yCMNOGYKS
ltC0NJSYSo4o69OhINBQIjko7gTu7FpirrY/gHJicU/X97KmaHRaou7sdO2sKqvA
qhH2rRs0t/knJAmuGUmRhoi+ZgvWjysyyBlIveXVBIaMPBzrMPUE02DeVLewWOzI
sUtoP5ukHnXkRelcf4DN0DR9dUs7qcJGBYqED8Gtziz/9ADMoxLy1eM0DHrTCxsl
ZHu3NIB2lWPipHextAmLYq3N827TRqeUyRM2vUbIo4oVdB8Ni//rn/u2tK+aF7Ve
2gadjxNxXIEK/Yg6PmCSFMnxsdrF80zVoBal2s5KA2iLnNrm52NUJiZKGSNN1k3k
aqSXcjonkQKUYD3k3BK/nKPtj4n/Ik++uqQm+m6X1lrV20EWtVl1F0idJUW7QGVd
o6BPxLJaLOLsAW8ipFikfaOU9NEV2NVLsi02n+zs8kFh+clARv0X0duVVGEnFKe/
q7CB8fhliepSD8UYPZKf2ibFZFTi/3EBU9PyeABXZ1BBG1tNPbgDsYR+zn6PNAj4
HsSaF+GrGav9ck8pB/DzuuLlcc57C7FWQdw6XlkCtQ+8ofyhUs4YsT2Nr8SQYQBe
BBfbfSTjpdVOSKo/v+lc6eE/HiqJh6X8Ikr1lym0F559irbP4gZjJznVjngqBRac
mcB8HrBPddUF2eRIpamXiCcZl16oNs3DcA3fXiHr005o2O4JhMdBV9V6YLFZ/TdI
yJFBEZSbf4yN0G1GwlCP7uj8szP8km8krcAyBKYNBrsnqxIVlh0EZDAseLm0PJWJ
cmBDgO6mragcD4cr4O3MsXrDwdARQTexo5cNjbabNYfPu1FmzZlYNn9d+p5S9Aka
ugks0P4Ay7o/4d+r81iRV0yp+CV5lNk5Xdp7iKnXf7YDDbI7hiRtLfGcwLTT5zNV
oFIPLt5gmP8fVgEG5fqXliR+4hJOGowoIs7LNM3HYcbAGGaCU/kzkd8fozwWgoZ8
gXzfg9VfUWIm/bJN5NHruYbWm5VsfJQ44F9tQeeQ9tZnObT6iQkkaRTVfV421Rk9
OQrOBenh05e4OCfEYoitmjcVZqGr9AoByQWcH68hPz3ZcCWMKcxEpLbb+yYzYTbi
wg7zD2Y/DZBeHHnNs5HyuCeR2/5Z0R+erkSqSuj6jxkL278kWmGkL/fRGiqeQF2Z
leUvjG4OBFJsREP+GRRcinGPyIe1Mx5fOIY82CEctQxYlzGmlOBrZ1CcyZhoughH
+eOWagVJqO8EgiuHo11s+7mlpjmXmzY6eeJsszuDhUJdS/FeeQN2E/u/nlsoUFJ6
W0GBzpL8BndEZUtAAuBjkWJi4VVuV66kE75NdgsTXRQoouzR5eyyWpPloYxGQa1Q
vr4LBCP0DkW6LAyxlln3j5rnBgVk9LtAYNOpqYjSE6F9qELyA0qPcCBTL37rkzZM
NKhpfXzim13O9wpGCxEw0FcX/7c+M7ffDEmc+R+GaK6zgv85le9kTiVnpkVuSRuN
+w+5+nF66dlt4ZhbdLLHQp1dxgAt3YPqoasIEWy+IprwhmItFZO8WubJX0GJemsh
9jmsnca8FEfJyxeVAC7CXTiP8TPSMp8r3xGLyBizf7BSqTV7Y4K3Obr8KncDC/U9
99M0YYYvAk/WeIXAwdKYaluYvhufvMCWtoQmapaWSoGGwstPNrQmp/tBEoSXh9qQ
/++nav2BPTaMeRrlrdQMcTzrnw2it9BKRAo5zt2OTKgEk4d2QSgbKiIMxDSXbxGP
BlVcVRoKvjlXVZw4Oz0mx0hgPD3qBKFVNwVh2Iq1LLGS94pIGLEAZ79B76yRTlMq
vpaURR0vBVLm2EPBf3HWUdjl17QLLfxHRETcIvP7w7YCPeUM0lIN5uivyiIDv4Sl
mE7Wo4q4+IkGRo0B7L49CZ7ml0LVrvfYHj/5GiPLiV0nzmx6eklrbaKAtCmjozUY
JGoVIXFq+7/+wOAsENOK0Nfx5bsDQ4oN0OcHpHav1eP7r1l09wXj/6HOdSjEXqSb
vUyWgnkMgkRo1mAQZ1iUiI3pF6efPSvPumYTMIJnGqPOKTv5Bh71U1+u/Cb5e//5
4+5SfgJy25QEwkEvICBbhRk31LkLf71vGXYo9ch9QIxly9SxhknMr13l9xvOHbkx
5fVnPMQC+2kJ/AMZgy2ACGi8waMAe4tNADr5fNphlf3a2nHQ2nSZOssd0yr2JEkT
4adwjoiDHrAm34bJ2jk/CvfZFYrUbllmoc60+kT6Tk+/ICa9h35NUJVdia6NCSOa
YAeufnB5S2JU2ArOKsNrIDtBau9HIvesK37QYSSaUHv9HV3DnSr2hZWltK134dWA
jINAwFJpBsEVMZKCfRYlf4GI1fzx/vLAd0VYjZUZy1xKg7vVXntZKZqel1NrciKW
Z0VfXwrb9je/RMg8TqIdjpRhJHcJWt5BcUbL1eNI7iuJ/kHjC6rLWAKYa5QmiuDc
iieVhzO1Kx4tJRJNdAFMVoqj9Rnud7hBJ2gM/rNGLfNaPDK0/gXawAj4uYmnAN60
2GpEwhV4UrA3MSSqyNxg9TDjYD3Vx0ZOXYA8fk3c1dY7f8tGy7EwmyqPxXsFXom5
ewrPzbQS4ixhNvFQT3c8crqQ9hKl6WfNP9vuItgUXUCiU+MFErE4MdEXidUdJG/U
lcoTEmXFdDCK/TEE26xd8LKCIj9V5wJVtiB0RkM12drCrgrGO38x4SoO/4DpdUqj
i33mWK0Qh6yTgv8IDbtPmbEO8bSh4nkPXgKvtowBwte177zGX+YyNq/0wF4BmkZZ
dERQ7aRyNvsHW1xIYXttx/W0alos7BXp9+/Fi8xG3TmkvUVP01Yi6WvBxjOLn4z+
xMWI4ETqBgq5+iT454DHV17d0gUJAc20vVhYBEWVRDlbF4VRgahSSjjASn6yWbIO
K/D5Nj3uQpTQecmVxiMiicSRs7ywIhMtaMTDVL7eP9GEOsoFzhynQz8AQeW8h6PC
VO671sWc2m4pfrMAKZamfsor3ga8g/XzpUOqYXhyEJSORBUeVguxNzMeiMvMCwvH
SxeHrxM8/pEAQSemXQ7y25o7DQSfa/ZEu8P9b1R77YwwKnYDnXzQMWlLxIBiE4wt
CDSro/0CuTP/cHhrJIUGP2DLZy8WU4+bVQrL6FPTMPMi45VC229Qz0IABKcGgAjp
C5H4VeVz3WUBcUNOmNn2rpSHoZtkwc8VYYE7AeFVNA2J2MUzsKI+fWcfk/qKkgSX
wrbdZGWTZljaJ8JPm07xxHi8YEHAMLlJ7P2fpI4lxxRN2C/bFVbMSFzevaAlvZL2
sNtPBJTusVh1gC/RYR0rtUJyLC99CT2FCua7jklq+MhfrwAr1U6E0g7/OnJZVI47
focrt8y6hbvxGwKVXRaJOeGQpehmlLzij32VYGlaD5bJS/ohhOncWxdCBQpElMzG
oGtJ720plBBP7R5MkWZa2qO28vt3kmICtX4gtunSlHLs/ZyMCtYSa+uaRjNeLech
F3ZuK399LSBx32t9q2ysg3Q40cJXVNW4oK44T1bprLQc5m7Va470pC9FwlC56ncv
9dgQp3bHMQf2QRjx0c8kJzYPDyBgKpThSAz6YS/c+uoa9rJFmUYB3UiMwEoZWJVV
YMuQoEwQ7ckd2g0AOQ5rLpUYJ8X0f3J3nK/zqM3QsGOW/3KgFI7S7lbcdbqKy1L5
Lt9sHxw6FxuficUwcxhI78/WAxB1bMT7hWn71yzThB5P3Cme40GmMTcbwxNI2cmu
5egeVMYN4GJpFEtmjrXk+dlAGVDYkBZNtE85Twx4xwcifXeWoHzudQGad3pMwBMT
qCtOHlPE5L64Gf7YEYo+OVYfYSct2K9uD9oaG6PdexDVkb+mMMWebq/fhQcw05Ei
lZRQ+Bx2v6oLQKAUnVh3N71mDujq9zq2oqVOcmzcxj7fTCaWW+vG/WH+6Op8DaU6
rDfaL9jMDCRkzTgwdo2ZTyoBz1Cos5+3273S71QY80LWbFDaWGzsr9inNxx8vcn6
zC+TLviX9IBZCVGV7j6N41a29NjXhROq/aM0aQz5xsINh/jC+Q7ERV/M2pXl0MV2
EH2aWNXcyoTnPTQqVq7Wu6mD28mzBvO1tqxGwxDTX7P+WkkzSZP5hh3UXbWlZ1sH
FSbi/84hZClXZMfdno77oZ5iHP5xTag1mX6PpYIpFwrhfUrBCwmUp6bW5RcTQHBf
g0/F+62568G61aqpDBzHM4YuYDwHLlo3TycFAAzyaZnegeBwpfiSi6Rg2wZJcyrJ
u3wSMvkAgpvj2tpJPMcSjGa38OIWOYOHCHz8utv/KYLa/toNkph/b6/D4qOE0iw7
DCfOvto9oQ/0zhPy3OPIlxvahlvpE+DFGoQC6ekyb7CIo13/S1995WMXXDOtEPVH
y/wpY0IXV7rQAi4Ou+Z+Ebd1/LNEX6WEC6efsBHo5nga1ZfIXSdDS1yuE8tIykzS
81lXWRcKyamneuF6Fg1DDe+/AaqlteX1tlqQ2etAtGLqji1B0wnVQLFQZFcedX0l
omXCqx+q5A5a7TzzvY08j7YLDfMKSclIC0DGKRldlY2m5rorg/FqEesBuenwU6/c
F+cbi3fwA5WYt6uC2QcpbMJX5RLkjC1LlR8hPI9lOu/otPEyBi0OLsj9GWzVHcD+
yt5+6ELuiH75UZTiPXtDZmWqZdcUpJZIueHsL3MOacp6r4gFI2D6BNnvwaxG9LTp
F2fHcNSvgMtoG0HLbQEICKgfjojOFbJ2QtkLIxr12MwYrPvkinwagnB09CabLSDS
7GwyzB4h8YVq9jZYQqxq1j3OVbn9aNipJkd1Opu0DU6sW91D/9twJumuhOp1iFj9
Mr2mx6XB2e52bAFUc28eifj6KxvBUq17t8jzsSet0g5Hhs0CJuEUNJidP8CCVpcX
JCS85crsiOmp5tHbVzI/SEXiaaP1ETTEEXZKCbhqydgEnqiIfy1iJhMc0vE4COBz
uOTzJBwYERNmvLR17GqbxZuU+wnv+3jwv9DEin0r8It94KhCZnY2ePb19kjgoJjZ
5j1J7sIGx4Ey4arh84EZBpxTtPVAQhM/09s0pCzwXA04zv9qDNB2Vb6p83GuLlSC
nunae0tSufP8FeRquFYfVPOW+vc4bU6+3neCsZNccbtWsOHW6LGrpEW1NWk8eWO4
cdj+51XgrrEICYnqrBHkAs14PCwxqqaN3+1fgYvAnAIh35yrcxwiC80YComJ6Qc5
3LYLnXTVZQswDZMgujOTpMpEcAyWv7gUkmgDg5+kGmNvAVX0fDxMqwdXyW6jspkf
EPa/2Ki+MqmLzt+8nnq8oPWjpXLMl/AjpRw2DryZUObEknD1fVBWHYZmI8AazOcg
vRqfhKHR4pdam9UFkiOzPRRdrTuDuTjm6PMcnNZ/WSzgpkjjmmdy/wJCK9mY+UVh
zxpwYfL4Br7YVJ1K9sSxnQe5oWyzTJx2haAsJi0pRpIzuS5hQyO+khShxyjLNZeD
QyKJuxSMfi4AUw50oZkteixcOTG97+DTmuxY5Owx+JPBIFLwnD2JFQvAktQ/bGk+
FLUpAt1zawFqzM5P7rG/YrP08R9F+9LTs9ITQkmakwugFR4X/BoNPhvjFL+ruYII
rHqpL7rCvY6kJnzRILMIus4MyrkPIDz++ZuFTIAP0MOBGM1f/Z5zAccfU3haQJox
JJvI6UnzY9c6wIrhRQzE0Qc8+c353w5SqmhcMN5k24ZpCNJF8d81cgc2+GYTqGXO
cjIsC0+G6WiMAASeFN7FBAPe1v2WaQ7eaTmoNMA2FtVYt1Gdw87W7g/5Iuv8gzII
Eddc+DCWKBBdEvEF78Od4R5/JCHt4woW9mT9M9AT9fxazSXSJTaf3OoLRiO4paGl
rPE/TV0EBQHmQRpBy/xW0Pmz0jXtvEZPNnwibybic3x+ZKEXKhVGX/opkejrXwLQ
95wDK9V93Xwesu9/9ZoZn07/o2yzdaHs/3W4H3jPs/C4yL1jFPslB/+HJSrth4ty
ZAQr25BUZKhnrssQ5LEEoqTDdyU+NEwfee//ndqVby6gF3kogewgJB5zSH7r1EVx
+YiXVtERhaqfEhK0SUHQeq7EnlJ0ywMam0UALQlUg80UVmEL6qa2ks6HTQvGiVWC
ExzFqXJzr5vKuz91u1davO+sxQVvRKrjPzBjIAhCSJV98WmwtlluMZIQ/hjTd7or
/cK5Vzfk3HKKFvX+MJITIRsSws65l982LVmnU+nrAnuSlpWZhRuIx+uwJjurYrAA
QDTS/EXUk3iDCDRJ1x+xwUcuzc0hGGI1Q/9G6lvW/0wt2vkWlPTF555pk9xh/+yy
8cJhO1cpXFeW5xKjuPhV0cEXSOaWEhBRUYdxLNpa5G6xchzrKdmp/buE/N7wRyi3
2bVLgjKK3wQwLrJA6aEITZ3JD0AbjaVXi67yoKlkIl5EPYvmwlt/1xL+p937qzgj
BlVauqSlNJQ6KOeHKqFlr/J+b1O8gQDKYuLfka8Mloj410uOhowYExhnF4/OPxp5
ywzdSRrESy0K1IySQn6qil8OaG0Yxyei54YiOXs1OCv1CkwJQofTfRRRawizQ2H5
ITg50GX09qQnommyOlym1h3uLlDlBaf6JJWouBivlNX9VKvJq1I71Lrq3l56QXS4
1NerUSGct3eQMoXOKiaU3+ymlA7UfUy+Ry/eBw82IUjipjlHNWeIumDI9Eh9I6NY
wL5hpvMw42HwsClOkrz94Y66CdYe1S8psqV4YAES1/BSM5NSxW5k169zj8UnHQSU
I13NNCEkD0dIhcdErDtbRrssQnNfeQ/b0b8ro3555/coGRSOxp9UakUoKSKGAdR6
ol+txPZSwbGk88QNQ90xDTNOqbCUcL0ebvd7T7fbnmNLA+2RHo+3gsUT0BuHGcR8
zh6nE7UCy0+cJO01xKzfkMgspfYXRnDJ8lWGO4yYlwsnuoNs3WdcIt8yXNH3jYxo
6nZqtsHskeuf0yszPJlNPBUG4WMj88LE8Yw4AafGkQpNJce6hliZLhb9O9GTpqe8
OTIXU4TS4F/ApTZ2xoD3rGgy1EcaEOikI1sghHZNoW1WhMxLmCUXSjQpi4lx8r/W
6OGk06bPEAiG9a0ky6TholuSZvDwSO5ffCDUjqFhNRmyNuelUp9bdTjwcl3/EwPJ
83T9kIGEwzaXIYRK7tm9/4HWNA3dv/DgaI36BrsRNYf7AySf7t9/Ao9zjkiHqj/x
USVc1mZMV09JAjjO1t/JxEMrmaRBheyj1MlDViy/rODmcGIANBTpE6dlitz4/cO0
XaJBC0Em3ecmyZG7U0/TYM/9De7cAPxPbaUzRPdriSdNTV/dZ3IhcqahvzwXjnyl
zPHuRE3o1HbRjZL0DxZLwLQmC/SS3xord/Xe+/JX99RE5sWYHPDEPUSzOzK2Xihy
ckVqzMZ/7+QeLjg4WzgF2P5edA9aVHMiWlka7aMvow8LjvzK4Ym064AxGAzufj9S
vr3kwr/OUf1Zlg6D/VsShYC74erFK9LQzDhSCVBfVAUJkoAk4ddfnOxcEqfurlwD
ycFOTAMNXOQ6T0Fap+Hi1X01CI488ea1emMto0O++17TZ9T54Ib/M1k53tQy2QfX
Z9aRo2Ny4ZyH+a1c3RMj7D/2pKOTW6KTerbnS/ZPDoD2xeUVSa+d9fozdNorm8Pu
xqx0+dNeXUcn0KD9UXE7/WlfZArbYqo84xQf52Y/9WVi866CbUNWiFloiR4takPu
xc50WkRHus0yiJt4gI4eDFmAUMpYDnaEOjnhPrbFfqLfc4d0CsNQoEMPtaVIskjk
xFpWAAjHbSmCVi5P0IYFYUcu76bkLvy5jRkxfswP098XEt5U3jLPQG8q6gzIozBV
IeuDgmeFgfAzOPz94qrn/lot0RYgKiCS3xjpEPFuf4TAvmj44eRijeobUlqjk/6A
2vmDi4BZT2+Z8zl+MZQCeKQ6dnNemG3A8ToZKnIVYV//doDDcvvKQIOGQphMMiRu
dFjmN0/UHZeS4gPDj+5ACgySmIwzdEtg82Va1acUDupf/8A6IoamHVypfGC1ccAv
BBlZOd9ix6nc7NyKa7cL3MIAYE7sr401+g1DNbsE9iK6HE+OVoolCBfy+6wGu9RU
4by5piAM4HGV6LjoWIwx3o2YctsPD/uCHMTDZ7jb2ihK+fHx03tA/InOrhkZoI4R
UjFpUDQShIDs409euMzM8YI3/819xJ4Y6WIw733axvNPpPBgCnglQAIFkqtuMOlm
FxWkpB5TAzSW7Dqz4yZgUV5gvPGdbAos9RJzi7MMZ91OEchJRyBJRNNnwykozB25
GVUQISfdXPiiczRtD/yVt9IcRUwFlwV+66F7Zj34kEIHIHnPj6aidBoPmzV4VF3W
VaRta1eRL9Z/NkNmYEJL+gsGzHx0QMjtuWrEzL/jVn5tR40ReI+vVk7drDBcoEEq
SYIrw699J6q1MiYUWXZbIHgjkbWSsJX4YNlOugDgthTB0GGzDPluHQwbV9If/vRa
jZ3noe2ku1sQ8dGEB6xFcyXSDa2iVkLIA/DuJaIdjauLlnjxbozmIRgzPP4zzns4
TRiZONxjRfxHQl3zW1gG36JVlCKN09lOtEvvuiT92xW+QOzdeALeUAxRHuxtRBCM
xzdlaLyVcA4/KBjWzzMEoEcG+bzxtZ0kI/Y9bzFxoCoHe0sPi6njgFK06gfCxhIi
o9Ly/ATmeGbaT+Z8E++vfb0ePURIsZwyAegyaVEaf0YRbRb6iURP+ksaIcCq3aFy
mxL5AK63QcaQil+snbM4f002siBHEyciEfxxhfpLgT4jrogXeRoZw6OuT14Z43z7
XtU4O0Eu4xWZcPsOVFxl7Ix1+GdgiDmRRn7N09DryefJl5Wa7F0T5Yl1nOcwk43p
XoMtAG6Q3InUdjt9rxfd6WR0DkPEORwVjwIGoDwauDCmxpS++rXyRQNssnl7qXin
opgTVk0jiic+0laMTos8JcpOKRrkvsp2IJHYmf8cmLG9SL/CR9KNZEEc2k9aqMiy
CYRVKUzhSIRcXEb9/UYtsmOjW4r389ub74XldvcgnKNsfBDI4TzIl+U4hCSeNOvD
+F4IL+9OZWuZukERmcTKq/m6atbgCN/FPHAXhA9kBY6Y10qhJcpw+pHDGgCvbK0H
0wWSSNTCfuS0/W4kUXzNYrGU5gJdL35GdbQ2oEwJgjqXiKZKEHOaupfEZpKk8mg3
G5J8KcQWoPN+guFs/hfrQf5XkzjstRfbSS3bIfKuGk+1cpy5cNJHdm9Os3jtA2XI
9FSr67XgGTLkAzGPRDIjTlaQSl5UcD5GE+owpMKAqhbIxjo+Krc5EWSbYLGNy/+V
GoWNJNYK2FHpF+vE0C4XEzCO/gfur4vB0xNdApvvitRmTXXB5FjfxkvrkvTAsu7P
O7EJgUCF8Tf9zNn+K15W/O9hAsEllnJyxpW5NNrQ7tTxn3zGYEmZhDiX/tTMbe0m
hNY66gINXcuqNZu03gVW5A2eysqhvPLe9lI0EYpe+IhAFwdgl4l+ei6nKbij587U
LoUKeSVm8o28/vsOJr2sQq5dIGBYbdZwOR4m2OAL8X3Ck2JpZzW8LfYceiM6ECsL
7X7qgUpqXxej0OHVxZPbakAJVRKPfCFZa87XId59Mr5CyaYTlK5DmEMxEFAmog3z
6RTIPfKznartOXSLQinxM5wURzRp4J2iJJh/GKhhDCMpheKKEGqbLS+TYIlhtfzN
WRM30jbIVNzrn6TWgi5Fn+pAg+qlTSO3BPKKczNS/N4UgSRNqCZDnkYDzCu/9r0T
Q0fzd7jiQ2YDfWL5BT0iaoIN8jXISZOgfp6r1nkDc3oXzPCnfMjoW52O7KilTXDf
lNds3JFfpT49uitvhBE8Jp2nH4s/VbugCjWVw/caaHA0/nitW6n1K5KR0vkQaLmD
TwwW+JALGdhdq1H01ab1eIQ/AZuDYMXTCdVJEmhk5rWTN5VAQ0cPFSHaiSnbSw9c
qDzgfifDAkOA6e1gzu23fMqRncZQTlT2C7LLyEpVzGdN5klsLifmVIkfqFQI5Rg1
EMMQ0MiJW7jM0gSh3Zgkow+XqS8maobLnW7vWK7AQ41t6cO9My7wGIvpCklTAa1h
uiYRto2TNakPxIm/fl4Rk06+7TKsUUwbNLmIGwA2cHuIx2c5+9VH5+X4M7BQfeHX
7M+DLckw46jj15vD1oeN/gw4fdbPHsgdui+dT0wAzG7ak70pPTrY5T7pp39MkcVS
ko4IQm+18m1dqtLa1Cm8FUc6GeYLuZvRMHON7AFRdMKiFMONbgJkN3T63Z4cFHt1
WRrTa0OVaJFMX7hfNgLWxTm7LWysNgv9I2dDqAblXzRkbxdkXpthXl1g2yvVBojy
aDeLUFDjrRJxcebIjwQjRxXOSBhTWsA4cCkBSXm5DVfvm50xS4PKBfaaDVYrDrjc
yE8n7zxDRimBB9B13Hwaxe9DnqOV5grve4/c+jxJuRyPbsCM+cFqFByVUAK77jcQ
IiERGWj1A/4FcWBZRcYFhIvHEGJk+mvNnc9XprY7khn9Qgkqwh0G4r76lXZrFARC
bOzftkEuQdErIsC4VB1L2ypTCGckXvVAIfnrZs0RhoVoGeDg1T847LytIQmHn+3C
AH3B7bIKGgd3n0V6yhADdQbaVixqYsBnR/aZMLJ/ZoWpByT7AW+Z2XLPmC+I3S1x
KcpCJ2DHlfOE/FJdOqNqch3dwVuERCXL1fgBcnTj5zUyDoKzf4KXeQzQMi+vaVZk
eutlLFo8sen+pJwyVDjJTBgBEi0pYadi/mNchvc5L6ngtV0iUq3YlZ9jm6r3zLEN
7U0G35lvsYe5Mcx0o/7iWtdGp7zZeHg8NjyIAkPJCqLrBC6I4b+w3nYMsaocr45H
o/pMcIXj5U9jEZ/ytWl0MpMLY0/n96Mn6oKgx4SbTkh5kkDMlPkU474w6c2BomUQ
fQFdpivBP6tPodYr/x92zLZv7pdrEsTeoCXQ+d4VnFCbORvuk6Tc7996tZ3u1gZn
heDBMyOQ+LvIufkH0kihs4SD2EekzERbdYyzDBrtz5OjSuS3HLpjr/UncZ1e+sEC
c0OcshWecP+JqYPUydzezFz7dJnDHBCCrwEPtbb8DOzWlXI9jStyhJlK8brdi1Zq
Gr3L6AE9hVh+dx2GsJhfnbLiyGEZI/zvEccn3VEtLXOA5l40s+FgzY8g+2ANaYFZ
HyPE91KlkLxdZs1fCKsb+g9PV/UMlSNp0xHw4CPPpVUZcPG72cKj8jFYj7x5/9Kk
nVa4oY/bIO8c9uaxuBPQGc1SQx+YroMhYz/UAOWOIuY9FkB3M0Eb80CguShIQa/P
WCzZiwxyK6XTNsAVqQuISycwREuX8lenN78ksixrib3McS/mgJQ6Exh3cNHQ/8b/
5lHnMeEcsSVHSOoSH2zZoKnDa/K9ljvwRNvNhIQbjt5gDKZnfBDRhJ3VkbZM7AfC
wNJsfxx5qVm/rpkWzUd7Kty57QCIUR3X+5+rPrtwHO+5yCHHvXkquaOlw37w7d9O
xD72hJfE/DOCrxl9UQtcSId/CS/RTkJHCLdG4bhc9b2TYJGHksAE1ge4KepYnXO1
fV3E9ZBob0ME/YWEr+ebHsg4oe/p5ljiMRdEg8qhFyUt5G6mWS5n9Fq4bpCxhhQv
O6hS0gP4Ect3r/Adu5aXSMaIjcZs3D9iuvOi2K5hgcmjer4j5PmmW3flhTOhu3ly
5apEPnbzHutDVms429PMpYS3yW1KTtiMmF8P9ToJZut28JLa+o+sfeebm5V3JaBk
XawJrCKcaFxcluX4szHsD7A3BErVla4Tb7RaDj+HiVHGj8Z80fRpeFNvLSp0QGaN
ifHrrACjOdUMfLskWprDvP/3D7QP1xt7pS7b+VKC+cR8DPr//lTCrVCd2hBv5wXV
e5od1sj5iaDq2pkTaHlQl/W/JfWyhgCFSJum/T7Er11Ntjj18W+K/yXA0xNMsz/a
H9yBEz5ld/nLuvJarofmmt10UKnOMbl6LG8mw9UjG9C1bMGtBofPZM5WPQFXOkSc
JWOoHE4DPz9GBqy8Y++udCNnhjeNOIpF5BcADyndHhJu52Ne3l9+UTyKg22YUghv
zzasZvyLUUFUyCTXL3afCHGTnHoKCjHfWD9yvpvlR3pQjYc5Fm8eKfSSMBnnKv+R
bWnajpJeOumuNllpJ+ctMyKxdPhfdy42S71Zh1EQMEPuvJIuPc0xmrb3fWVNqPmA
5EAmwjwFiVFArogS22ZKL9P7dWvyqig80H3Xba/4eERXNYM0FPZKQ/p/Jcq6Jepl
e9ZQS1Ijd60OL3WKn98zjLfcpFDbsnmBvg8WNt4ht+yp4BkZvSKRNCDYX6FR9Oem
uxOm7wihSVYk32o9tQk4mwSpkVaq38oKr13EjtDl1zOgRkTJZrVXxiFrpbtZACjV
RAqyRH5toxwBFLDFVERjFkI9BnzUfbQ9EbeCkWzQnddLep6vNLDGn/3OHtIf3kgf
XlxIFHYDTxteUjXVTA+MzIURM06aQMVOpxCGB8T8dZiZx62qTYUFWoWWaJ23zcp8
A5fIzye9KuKbth8MpUK3bceDFG1wgP67JtqRb9Nvr77U3Bibi8nL9E6YlOczJdEe
eHQDCcBBLOQ4VvCVaRotJOL3EBD7jK7fGYwGJuZjbWNjBEMBiSnfmrRoUR5JIjc7
01AzwxKS5fD1iP0aeel5PeRXNWIa3mEqwL8gqAk/IEmcILpzlUtM0sPdLQgYw5zo
WtCsHM1lO39duX6/PT94V/dHP0QU9QyqwZmLre9D+ACEwK/TjHQfFx8EA0wn9IRF
hOhN3ZYC5qv3adDjcdlgQdFhAEwQB3SpziljYxJafPxi4yHRQfO5p4G7ip4CN/ib
iBHobniCi40N1IYLMsmn8GRgUjnYSiQLpJ6CC5VTA6hqCR0NHPnRqWcCAR51ndj6
+IdT8by1hy1adkgcoZ5IhB7E3nKR7G21i1wAd1nJTxnWkolEoJ7Qi8fFf1upyF5x
YS+Os9ksIhDPzT3BAtch5IYGe4eFqZjJRtXFMmaS5sM9OqsI3EqcA+4ZHlphM3Bq
MHG4jqyN0bVcalzQBuaqhEvda9F2WSOK9mXltZIrWIzFGGlay+5aot6enD4OkijR
B8kXmnqJUJaNfaS3tgNoj5yjEImslrFOiJQ6zR0lgZoOiIdkhl//Ixw7ohtIgZ8o
C81L9N81+996O7XBe88+3Zh+q3pf0Rca3bcebyopFiqxna0LFDHO6N9ZvKp3AIb3
YqkN0WNLw2C4+2Aq0tFQ6eCOmvRgNVLmpJk++IezdKbFj8E5E6TUZi3KHB89h0C+
Wx09+h6eZ1Dt/vufrGh7ypZSbQE9/gqbn6HIO4WynG3vOWshprxoGDA+PAGQyNdF
ZKXCA6Rt8c98jzRuRvXSq37rC+69tJNYivVW8nHgAXGI+R5oF+GUO6RAm7XzbUw+
yfV711EArpHoVIbGGyF6fkoZ+UF5wezwNPcMlMlpGhqn+u7L+apUTBV78X+L9SHl
Yqsue6AJK2Cws7CuMK+8gYajnkhXFcTh95tg5+J5h+mzA/pzkK7iXvSTLSHvWrEx
KgcVcxt/d4x/WIyVPAI2P2tpZpmtZMU7DEwTixQRyhX+m7Kv062dA57kcs4ZDIky
F34RfkmXr6BJHhjCCvCBrJOSf8yZV9BtiTTnwfXG3ehhh+YRjLH+gwZ3gsrpALrY
9S9/CjOgaPKJBbnyAX2rLNnjvlICiAGTwWiroq0biuwwSPv1FAu2NzdilZ7JYEE6
ZcXhtnEHhOQ47AXQj4jGdB+e+rWyRswwm+FPjmlIJhTakcuWx0Z8e9wR4f4gQucQ
C03mJ802w6WWkjhvmrjSa6dhO6wblXBZEq3/THmBJX+zC1DpXq9nMkXL21uQo+3D
609v6p+QvhqfRMgKTs/LBHNXULcLvGYIfd5MwcMRcMXCb5IkmfNGSUCxW4aNSTcZ
w0sxUvd59nwT9QKJhGDEEvC8f/5yqh6zLMwnh8Wuf8y3Blo1jmbVhZae5K9Lg0Np
i80Fp/sg8AgT2XYCL1+jAiAP4LY0XAg6KDr1/swDROPDyMBCCxXiIMUUe9ANbABT
Nm1DlmDIk6hKPZKwj9XPE7TST6aEUJ4pWVnWNTHuA26klbToVBOdriINx0I8unC6
49MEZC8rKLc6NwVGz//q1oZimbeAXnCyGEJgbReBl3krRIgvrPTwtT0VYPzPEnG9
sznm4Q4r+VPHp3tIslxdXaMzptGIQ+X8m0q7IzIjknuZ8TwwLoONeRjmSL2vNUja
VstcMTPohpvxAR1PrAct1s5/HD6mWcbVZMbYBtd5Azn1rpbXQdjS0PpIVIB3Vgft
UDQoFXqYJsZwiiD1brpCjqZ8inIzu+qiXco91rmLXbcRvhACiqL7S9R1coC3XsbY
RWWiF/QEhMPx6dX/GWrKcnDWkk9ihH/FvCCmlN5/AU3UoJ5zxNXIw3nWZs39BRQ0
h5+FwbyXKUSKp6N2Qsb1dBycAJjPau7NHweMxzLcK7NV1kJcHc9TKKyrUJHq53vK
AkSEfHHQn1fqjytKSkW+9NRYq8AyfE1hGZqmvDAsfZUQGuiM9E1x73G1LcJTVSd7
CqNUjcPupYQ5OzsUE/cD7zRqFEh5BTfHOxCcOQ7UGR7wpyEh9IvYoHGIQ2YQmC5Q
0Wwz2zsnnTuiod+gfUrfPXhv0FHIKim93f08s9veriE/y2Rgsf1pYqJGVbFgiUJg
VoBCNmfKdZLeU0Cyes3jS8zTabSCQaxX5ykHT0LaCB12dB8j81HuAEQXh32IXc31
vCdZekrUvj3iAiMT1Ie19GftDpfih9kcKmshV6zk78rjAxhM72hVI7zmSmOr3Sr3
XdDkRVHdStmQbtbwJePoYErhfPv3nHhWfzTtQxq9qlZwm8hZbX+sTS2RVS8L/Uaq
8ovXmdoIC6BvNkYkk2n25zpxGXfBlPqWgDPfdW9QdIWosbr7e+kpt2yBT+cHFqcD
aqTszn5xEYbRglHWBhvC/NQuXww/PCnsB4NocV0yMjgnC+mMfm3V2zFln2ZH9GRT
VWoTbJS4F4juImilDEk7jSyTg8M8TjyQlsCP+ftpksbTxqgs2qy5hUrxG7XiCyq2
VGuNBP6GizcexXF2lK6ntXhsBvrPjili35VVk6ctEyYmbL7O+tFmugs6N8zqXAVT
5txKKov5T9TQTr6tFuK+WDgxITCk+M8wxqSmzTdZW0wG39iRDxBNBY26tdm70B/t
iVqASXFk9g20vmykL0ikivnWCTXg6S3sJyRAB6AM3B/PrD3q5xlzDbLVCrdsZ3C7
Hl+QFqySxmvNw1DF84eUPSsFrIHJ8ht5GQ0pA7ym9fKJUMqXK+RIZqcCgF6ygAxk
fE0KmrkSaSoNVGMHzs6/TXYoqF4yy32+gAmBf9avJlXi4lR1dKMl98alWDZv9IHd
NTomfvMiEAXpNdpDzAjVxSl2fnN92f+FnpR3S8OeL3gQk3pyX+EAMIBZWTV0CrOh
3bo0UEC0fRYEa3bpu1bDTq7TRIi9sixQFSovlx/XTTqZ8LxD8T8d8VbUVR/eCZLN
cQEAg4ziFeYk6MrTbq4RxP4tl/Gq31sTek8fZSGC+IT9UNp1uHBTLPBp/NE1w8JN
h4ab4lw9S5CZ/d//+9nKvk9RntMs2ZWKMQ+rXfmCLgR7M1VFEGqdPB7NeIo5qqkZ
eCDkjjSPiGork42kO+CSwnuPrn93t1L+zeKUHxknQkYJbLX/p0V5Tyt5RMLTGm7X
LSQ00EJRNcKYXbljSqEwMKrJrS7Ugk/RH8HIpdHuUC1+2fuNypsbGVMEVMQpOsnl
zonczw+RPIEtMbSGxlxifZIwNndvg9M0tcu/2UkBnnBPZPbtfoNrDeTvShbc3JXJ
h8FCbKZX4C7Z6Ti4gKiP8SNdPYketBRA9dIQMxt16EJZ+YXKXvEpo3DDYFD9OfJe
IsEK//zKWQeNGrqhHzEtYsVLvJ4LiDfKSsPQIsJ3KhXbsNUvyQ9+uYxyJOsJ+LVc
KeaR3UDRvNmWKQTP0Td2Dk8L4pstsXrAwcezpSetaZL+OKViYURZH7hv4dABILGq
Sj9NnMIfe/8ZsJkrT0MHZSTOrDgOBsya8UdZKc3Hk0qvJ1dfFEF4DnTA9x1QVfAn
B7j6Q2kbik95UUffDD90Nm/o8HN1cj0nj66GeMJX6tFkpOruMfWsYssDgYfIVMHc
QHf/AUI2HbkSjLPx8C8I5LfhVFXxMv0/SgCXXcczwXfHvOIB1PoP78z+wyt/O7g4
F0L3Cbu0u5WXMjP12pj1hTejHum/GWCquDnnalHJ62GmKg0HJoTUt37ML/tMBOle
gVY1/w9Zxm4i04pWBDAf2ZI5kG75DEW/55NVag2iiDOFibdhBIVcIiT0TP0P5dTr
NmO+zf6HVGKtdDFVue6seyYbecHHXAO8kh7O7dNooI7XLgVura5PiQBTHrJaH3jq
gWDzxycyBSRXQiuWu1V3jfeGU9gMAIdo/mJAjFnzh4m4MgeywlVRulTZloksO59u
XoevGa/jwrhsP4RqrXUZspBjjj5CQqGas83/8wcOxdfQdK5sQBdtmolpTwqxm6ar
9zP76DwOVtezVD1l9/N160ZutPrX8QhS8zFOA6A5k12XdTvESlZLkZFamUS5qUhm
0KSrEyhkZit5ah/Z2hWU6ByT4nav2imMeduKt5cRNNpLEMHo0W8rX7MswmVlZFSZ
m5r9PKAckYbsCv/AolvLF+zIakAksHE25hu1PhXQl0fGKhk45wpWXU48cbDdzbsb
CI1P+4uEeqxDBIPrA/dxKozP0jZvj1HB6xXv6VSpYKm+LzEbFcEv6wYhUIB6DvGf
jo9cSNzv7beRffemO2z4T8BR4klKxy5iNvLwwVHr0w9WCxiagNxZGau0E5AXAZkQ
GTM/iwPdbFdFLS/NfTvIYsF0MdGEfQQZ03ITAsRV87gmX+wN0qOkHLkeapgLiTpp
GGGK0sajBmriIuFmXedglxiPeMZBIENnJzkFoMIcEvyCIKKe0EdTpejT7lZtF90a
V/NGHRpj4afSc867p9TDx7m7z82CfFfFEqyWmWvWkbsKFtYift29XDHW2EJwiDVE
6un8k3HXr3fy4Pv8skTLT3+VR23XK9bIingViE2Olm1uwpyO2xbEbeDUDN9gRltn
u5tZWvX0JJmJ2L5kQAL6vLDWliNi04y3LD7l1X/6Gz78or0BlBpGZLBd0AA2IgIa
RL88mjOtVAALsnjH+e8E1snodEzfZOG6ztDHW3o8N6o43k6geCxmbBfY7/H4AWLq
KAAncg6SpMpApjKMDfRlOKrvCc6ejBVNu5ffUHpoXaN/fgW82PdlhAxvAFBiug1u
xo8kT4uoPXE3zVdEoJWCDhPuBk7C1wTf437s7ZCH1+FyJJmDbPSM+UZVPk+Z6nXP
5hweDacuu33Yd1cVChFmUw5UkibhE0KvCybnDZ/4umobos2GmQAN/q8PaR7mvYWf
O2iA/YPnUtP6wI2lJcC0XXkVIjHpmZzz7GFsyndlPabFrakuyP1SIUnv3xoy0bDS
3BFeg8KCVWyqLVfLZ9MRzkSCkjQmwTHq+wvyiqX7QSNgtk9WKMO1FK/c/VAMH2/W
dGh8/FpdchJR7MEGXBDGwybH17+oViL7dDJi5sPdhbb+0zrKGiHNN7wk+Hv84P0p
XesPR91s4fIixMFtmmV/A7sFnfILFxRqg3RqqjS52Jt68KmDAVLqyjLG1TzUHJDc
ZSA+lsv995crP80EpAXdtUDODEs0eE3uopjewGzlo4x5lN6VhM6gWSn/BOQ4maPK
CfK6is7195DIfbtNNFgvxU/3KxqRqAaQOXiLTr+hTIiVLeYMlW/KfhGuVmERi6eh
qtJXYnDfRlFJWiBDaKRMFd4bda9d2yhX4R9e13Nz9hJWgRDtrqFp3Ju+vKQrXqhe
izX1jB5L3K8A7MmoO/BIT36UyvMxw4k96RadnzPn/kdtG8OYfI3LmyXS/KFwz6Os
BoXg0ikHt0KoLoUqB98KFr5sLRXHRbshUlFdDYx5KEDLoDR7p7IDDlZ/l9tyGGp8
XS2l7IUgBBDmqnrwnObU8klN0Z9vZPChHiZe2c5Z6/jiF3sVlEhX8QbZfCEFDP+T
VIiABhjblmmL1Dr8/8K0tNE4CE+L7N0lwOKq7wQ82OCrd6N5LaVPCI9gvdhzufJP
ClHef0XlkvInyTwPrPKZsa7/sGAw8oxCkYLuMpG9OBxjBQizfHfPNcUh92qXdYdU
OgYvDvi6vJ5nb/IYa2zOJms1JLBWCxA2Vfru9OeAVOw6+8Ftsw01CsX8kFvBNdPm
zFOl1jBVk7ZDsNI3XwtQsZw00PtJlNoHqHsRpoWTSFzB1ykCXaUUFgsy5rLeO4Mm
V0VT8SVojSN/NUvnkP6cat5PLLmINIgwXw0xIpQOANCOfr5GVm2dNQqxrz169TAg
63y+WyNME52aKVrYOaiqoNWqSChg/SOMXaJlYdPNQuZq/dHKfh7Mxq5P3FenXdN7
V68tZEJgLUMqrAeCH9VWy8XnsVF8qw/KTqDUQr1Hr41eiKG8QNOK+ggMo/IXZ1Gi
SgsIUIcgJ1HR4EKzGPY34okAjlwo/iue7pzaUND2iIGcRZxhUIfCBToiDKE7Ayik
l7IUf4CBE2k56ruVoePHoP6yeHLyTER09kaVXKsDYTxu8uWjKYBRfadrYOIZFRvx
JLLFB0JHUdOUQ5efPiMPxeZUL/7sR4RNxbotb49Dmsb+4chsRWuLmZKpdl9WLzuq
1rpwcmiI0Iemlv6LU/ef7ecOb+3bF7nvmDaltcJrTNREiphO6WhQC6tczzZ1j8BD
aO+H6lAsTT2fHUvdTGazaL8HMwjOO8ZcgzfZ5R61QIdOoSBv1oRU65vFg/Nh2ngO
ktdyd+dxRG4ddmtLJy9Q4GLY42HwReKoxGC1yS456/dAXCsuLiiutfOEVEj02u5y
JL1pL8xmdQhcHNzIbZDQBj2Wgibc+ZNaJBq9Gpb3Hd/QMFGmmS49347ks51lIGOi
WQJ4Od4SDIx5ZM67V1fkmmXr9DZLEyvnR+d8j5NFsy0XK4Zw2lNMzBlmxU1sPFWj
1A9Jltr6MUpTxZuH82KIkNlIRdKsZJna5fjN5LEv+yFLTC/gQMCb05ehNW9Aib/8
vrg0IyKNEkMNGv24d6G8R7ACli9J22zdbD3HxHknJksVF1vEDD8WyuoKjXPKqOhN
jGCaT2pd/JtmLS4JoCO6GnUwV7zV00cqnISbFNBI/+ow2AbdiSz+mAAtVbgEzvc6
DvVe2D2Dpmr/QX32PfGIjPKxpjE06f3MOAHpHu70Mh9YbFnsoMnCMtLcSHpD97zf
mQ0B5DYDvys2c59B4PDAzlWauyVHZRS23elUK+nmEcNy4AG4zUfPNksfLZceLmpS
ah4pslE1XR5UiNIgwPK+Hdzou82uwHuSkP8mjPaA17BiVKqhVoYyCas9dt8dEOvA
JgEJYvwVFLVpVc6EyNTA76gMNY++hEPC2ODuBrpl1eX5EdfUTr5OnVYP6Qq5UwNJ
Cm8dDldFBNpkdJkWeRSFADiVW6RcRspd3emSjFqf8Qwa73L6a9ww+fewrYVZJ/rA
yuJIUUzqV+Np6z231gmchuGTGZRxB4FqniFdqIRy2zEBXuc4T2hOXl7Nl4qZ7Zlk
aLE7xWrmuYDJPRmbbK6KjdvpxrR+T4STbm5RUc/IJgW4Mnr90lKACeXUWvO2Liv2
2EJirGqirn32tQT9+OK+sVWLJ3wT4QsuPe7vEpHwp7sD/e+069yl9jUgHIX52jok
/Ie2W+agK4HzQS1uumClHXFN3wxjILWUJZ8rCiHlDKCqyJ0i7IlzSSIoMIz+fxd6
5O4PXnFtVpawdpemDU9Xd/1P5bRLPPHxKvVHGqJgZL5Oe3ifdBByfnqFpnYZt+xX
ufVl/2S0E9Uzwv1Rdnv7Q6gdvyg/5/vhbmcejgH9cxOLcjBMoo8eY2n6QehfWkNo
wb56zn4KrSp4MfUARN0YAwj/BpRVa9fWaps5sj7zYPgg/jih3y4VjlzsoNtfzEUS
HbS9AhJEU9Miw3aTD+iI5EKY80CkHMa8inZ1eiT1WlslS9qjhb53XPK2LIaF4f3E
5Ef4eRwMzyciaRbQRzvyhxrnnAVyM7AV0OR0csP34ft1pZEvFxJOofWZO/XUI6Jm
C2pOTwwAxvcR+fa5B2pd07VqWvF8nYkbFfQOOGDx1omvxgVZqxkToDaNuNN+mtCX
PLoCTKU/hV8ijipJWEOUMFVuIcswACReIB+8fGM3/I+rzTo10gl7miE4FFeKqN+O
QWStkUkOFzlMU1dJiaVC/LEK6IqyE9KUZ2rJ7biqQaP3fFRHk688/hsezO6to3T+
niTpr6MsX91pmPeP1BY3QJVdtMsqsWobqpgl3y13Rg8gilBg9yMW1re2k6TTkXyH
Z73AEjHaaHxZHtoRq7BpnfPDJ2ecpq1tYTomfoH/RSp9zz6+4cQ03XtjQhil1yu8
dxk7WS/P4q+s8IYNNY5u2cgurVGG0iOt3tP3Kw1rYaK67Csy7VDT/+FydmVnu4to
uxied8WHRw0eOxGO23zzw0Jsuf/+8P7OYhijHbmJw4cW4dF2n5kRn8pTTV/4JVVu
7puN6ZIjA2twTenRrDBwO7lzhSvYFHcikGdRWYOeK1uTyHOfNHJjp9BEoqhL0ui4
MKWwrx/FqFcIT8aftODMTgsW55TEvKV5u6GqeEk0UfgZJrYQ6lpeoq2ujtl1gUzx
fzW8aKTrQzM1RxyDi0NLaFFDwDwnaD/OarDVSh1TzxJnoVsnxZwVakJENGSHZ+BA
w0mN0LBUt3DztYcw7zad9fnbEyh9V1bDGGPm6tSlQ9I6sbKOfacIBtgfYnNUIPOy
VrqBeC2D24ARXC6TGtF/zp2nXY0F3IMzc2i/POt5/jurgKA7J1p6HtSeOgqXp7V+
RNVyEjCeQz7q2fPTY2n4VUkKaIDU3L4JpuOhCagwdgFru5MZevXnCNwsgXt2G1F0
U+P8V2OC1ojY+P3Ha/8ieFxJvGVOqM+Pabc+4pwhTucSYv253FBOulbwvqwJ1p2A
VGxbFWME68zB2V+Nd6Kjodd8SV8SbScSnx4X9/ktr/rzzqlRFQBrEl7n65jMgpp7
TBXKRQkM26OpYhJldcOXdkoVmK9xtHKqe/b3hkrfaktKjW8kF/aAtFpB6RVUSvd5
4aIS5qBHtfmTwox3zG3w8ACoZKdoEgiyCbmSsTbM/piCso3SWnQ/e/lKAS6hUin3
hkb1B+K+qMFd2A23+9tpVZGdOfJ57+OQcP89M1F/wxcSZYLDKD38qSFFe2xtbKQQ
uzhFtPgt5eAtUX9b1Gfp8VwGta3s5DiCXBW6WhwAHG4M6fppQUg9W5+sY/inRXDD
lJJIPnTt5bhBakIyZPJWEznBcZeq8xQ0mAt/GOHe5BLb5JAM6IDH8EXKq9PlVCeU
Xo2p3qf0KZAQLUQcgrG60jLvSRXNRgJ1vRQErFzLkAPa99+c6Ls6crlyEjgTsiqW
xZ/YS2z9RRMQJ3PAJX4nkMvstPeHoiE3c68b+n5w9Xn2IHALc0dk90muaD12XOrG
cBcIvtKEmkuhhwp1ljQPrS3r1qRJVFZ7VcBJxEE9yopExs7wZFJfEgzdEsMkWnv4
BnShGlJL+pmDpDR8lFeoXg2KvKGQnnydIyt/yRI8yLz6ZrPTuOF6bk84RhO0Wx95
gZLT3lzEVQEa/DUgso5u/buzSDFc5lQgPRezehVfvpmlVbJUKgfJTtv/krXDsH27
X3QHwQYM/dv50qw+3nWoT2E8tTPitX+0il1xN42m/yHQC3Hll+LI5nK+Wclbu145
HwqVRxZ5z5SoZvOZdAAZJpYjHQgtV0wWUZOkUf5Dhwav/0vxfOVf5288VazKKrMR
OVR7+EDt3HU5AkMnRq0hwDGo3zKOPQnAQBAI3m9xqVTvVJpdV2ju/S8fDYru1Di+
5L5HbS9gDKpJGUV+SuJlNDjaoRdfTOiPsg63zlvwZtW+A+2+VaynkgKsdJ4MPqaZ
wWN1nf9Jz0L6K1Oxmz05O9O9Pce4EPkSajHb1dize5EWW+YtiXkv/nHLITIpOOPm
fiu7yEejkxZqlsur/mkmbPw25THk3smCjTadIkjlsiIy8y5EUM89BTHRGaHwqrDR
I/Cu76LduSabF2nv1kPvgvCqAAfaM61txx4t/Tue1/3j4rBzz2N8S5iUBph72QAu
1UL/YQT6k1qjp7Zu128J+GlH32878k+xeN5+++l6fvrQWyENrnXknWdGhmhb80ZB
uCwvSKKXzAU/dX1Vek2zy/TxolSbchNQROtxq47aV7JfjPOzjb+prxxfrsaWi7OQ
Vbn9k4KEtxNm2oPXAP+jiQErNtUx85hilVKWfQ//8hm5RZYP2hZgyDYCyNjpttzx
i9cbnux0sZINeHttK6LsNi4jesPGoh+8AOACkbluNfIxTHsg+3soJxGlfpM3bEu7
F+m2lfHckxbe9/m3cd/6ovdqBmi8s+dtWwBkKWrikfwJQd8GTDXMYwW1ZLRUTFVy
zv5ze+LChmRwdvdmlPP685scrb/yqRWtNGcU7+dVd5X/L+7MWpe7k0Hy7/OOQZ2E
1LqlLNW22glYJw17OxrlhmMVwbsBQ684vbfd5TmIUpuTGcIV0zpiycKd179K6hgL
RGeOzj/13qud+lIq90EKzv5ewKJwF+vME+qhaRo9LjrSLQmjvZKmtwYdVe5cVTOY
sAu/wTcaCIunG3cFdLOupgV1uqr9TEpwlqBzEL9HKHzUAdUQcv+7KTmhIKe3KNzC
Zsrrs35dX8B8IvEziA/ropcWdVLLzFPXfQNkhJlQOZlAfcdmQ4Sij+TC8emcnama
Lm2ldFO4sR/c0QOviy954hPZewlEOxBL422j0KiuabyZVGltHss59ByPy+970TRr
0XfafxTWgksw0Wq2p1KNrx6oTOtrd/B6cq7YYF0FPtfZXAel4/GXlzyXwxKtgh7O
FMIq19kwruJpdKGMem0eLwIl/Uh1hGBrEuBgbzg2cwojVybVasTNSjlzkHusU9/g
QYXKaxlNpMePGc2GnKmsUqWqbS41hNSBmEZIcugHR881abqPRiNFs0PnQaNLfwJo
iP9dbHfRpEmpxmiUYz/TX8JWTcj8ADvsYpaQ+Qx8lUKb4CSu1jYQ/UwY+/vTxONI
T6eNVJDgJVkaGezx0DpOJR3Z6dJvMRqffTaHOR5RzQ8LGiK3aHFlmVZpJ/9FY0i+
ntm8dSRdud5ZQ3DmbwESLFXPcsCi+goKSHIUYYZQUTtbi0cfOpSihLISAsTAmZOs
KQtO8EBOvaggyKlevv5FUOEGi6J56WIwSjh/WxC7qrCbfjG6408WzGNv26MM9/hC
lF59GCBIgWZU3UtymaenHcUCgBNg0sTa7kdOG+PBvenVCQ+FYBNqLInEBM6WIkMo
fDbmnKhm/8PxYEbi6+SjCCs9dnyhnuag1I0LCf1gw3UCYV0v3Y3gf3o6724I2mQT
f5nqikBBhjXo8QdJZDggw+TeBVicdao4h8BtAfr0hZaUe6e7ejnkcv+aXyfJd6FE
texRzx6Xzg9Syf7evrXacdPlhu+7mALPwSzkGzoe2pQA3ICAg5GGsvD8BIVXlw8l
RPWIuRPzwCDt42OilHhUjWo8SMhsEqzMyXUJzzBfSt0XU76A0rbRUoKnyBm47TLE
C7iSGg1UyA0d5/UmTxtf1aofcONpuYZbgfuuUepEoFuGjR8nxk1nRn1wSUZiMfGm
jmJ3ZzEmvOnhmmHzfyJZ16vBf9kLpvyPbvtTpCTZFNtFu+YV5+5JGjrbcM5U/Gno
KdEp22QK5LQ1bHO/WQJp+b1hSKNwlBf8NqgWi+Cc9Gd8dn49t6sO7I1mo8CSnDkU
eELxuKH6LB12VUkBC+sSN6WnSA1DTEsNjQZg7eBadEBfRZ5ShwErgoBa52FAwyiO
marZG2H2jE7xu+U4V5OQUFSV8vNSXh6QwzkZ0JFSG8z7wrTH5icoFT+mp2fjWZYp
gnnJ5UjAfLpnGkKUU31eu+iI0YuG8z3BsF2trH0BpkfDsCNhKMw2A/xP2jxbMIQa
ZtSET9Kqsu/TfP/w1JwLhMQmMXvQHrOB99n4mIAEWEoVzlJD2JNCggZ5oZVtjXaU
odHqQGChn2CcJJlwqmK5hZjz95d4wEPrdsttvRY02p/BtbzHLMp1x2JkxowOZOmq
DfJJDm2/tKXBccGVyPcjl7lsJiIvkiq0fUkyv6iVEIDcPXkEqmAWXEr1EXkTwfc6
6F0o7dWYrC+Hk5XNVDE6edWiS/b8onLA/fMj/Z88mHoYBuycfN6Yvwz8/83IN2zF
VYK5Zlu1Jp5a1yGtPjV2BbBzzXSz8r338fmDwfU/Xb4C+cVtOGckqvRscAm8DClk
zohd7c+bUtQ5fzHYdP4m7R7nAAz+LMFsvNUWDLwgsqQRUhCFxQpC149HjFkQc9Fs
qJhcGyxLLWWzqsBGXg0szH1SsUJE132y665NB+xN079coh5I8x64NLS8MdnYTHiB
SGDp1YpRbpQCb06acDX/UesMV6oIgx0IBTbvS5ZosBzPAswczLmRFkLICD63ZrQX
01Y9s9kVge7Z/8m8xdO4IPR9moURflla/wcgUBZjSwwAvX/s7SPWCHeac8fFEh4l
8wsubsfZvMtYyKabS14HN1hkei8dbhg5dMdgToLgLHUq3rnngInbwYYNWbyIWXRJ
O5bnmRukreDH8EblPHVdwL5no+L9M17A9BCZepnhNv7zH03MHoOXvhv8k1X3JnVe
OGzMzQSP3D80nM/qxIb65SgqpPR7sNgMLhw937VcwkclBJqpBwpqW69yMp+oMY6r
4twPcZmmm8cYVZjmhAAZzcceCSO5ja1WEoBZ8eR3YT0MSS4icA/nNHsBXmf/FCOl
qkDodq+m3ithXs3Ih0UOyqUbQGEbJMQnCS738JHIRQvy/UchmzorpEPDWjnd5FEk
QK6eOWjnG+323+Sdooz7zfqEjAAIzs5j4ePZHrWMe2sGW2tb5/fDwEPiYjcsSzUC
11EVTwENwNX5DzNETRg/elFzYDnITAFXvNlDmOA/mFLAizEbS8bOxlxGPqhDfHdb
ed1Tq7vh8Be/tgx7HCqr4AqTV3mkVqaHZebzPHUm0vy0oSVen1WR6fI+VXZJ0OEj
kwgPgoJQSDEFDKH3l5UlPniLWGkb8AxFfKHjVZfx/fm2vuPM/0mOjtROW/+13FOB
W1vyx8YDD8/27EdsAIs+KoHwBoPgfNCIgazK6KrEd7tATJFOhUc4nNzYSv5mge62
RXbC6t5P9PvTDJxo1pSSAtIBKGFZfIEZyISEBO2IOlz08ZniLeI2i6a9GT4js0FY
LzMoxZ5ACA8H3mssp5OTFQPsGkEG/cD4pveDwHO6VlFXr226N0METe+m+RlJviwy
OJd2qYZyc4Uj94KIhv3o2KehEfYeexzfITxnUSRMCJHgMl0MxCSbvjiOjGSQm75C
IHvXDxbQFoF2tYy6n99FL7+G5BmWu7g+fSWjAmceS/EzL17X9c9BGpLITQ9Vr+Wd
SjNWsJJ9sScWr6CQctXXCo2IjkwhVjXqdJKtA+ChiRki+erfGm3Z8wHBer7KL5r+
56pQoThZ7wNULUksHjgjjM69lq2uh6BqmERM+gAyyLIa1EybB4ls129GOUHT8he+
wWc/h/QDDTB01A6ne6f3YWg9QQExtbwlRXUC1Y13AJD0BQJoKEUPfEjOnInw2MF8
RTCmRNXLVYQy4EX5/hRkb+Q5cPZCkx3RaURQeweH6smBNBZneAwMGI6iFMfY99Sd
cZhk2Puyui+9bUyfzj4lQVxCp7zHoktxwZuKaR5WbcdTCiJmmyX0bl+86wHVtsOE
3RYZvJ+V4LUCFQpzaDadICiSRkpoLd1DfC4o21hx+QFCE+U7vbFsqT/SaLFGVS3X
AJpDdq+0ftMJjvVmuFvxTtmwMRe6faBISbb6/6AK6W7Ued/Hk+FAwUNZKMwZDKIW
/RxhCkLNc30oFLHIiqda94Qo2OOxIoO/EsLd70i0A8updwRCgMJBTcvf8iHaTu2F
UXvx53rDxfW8mQFXZ5kaPQpGyzO1cAgybXetDhOuiQZIxVnAXtDM5BuiR9hiC5PM
JWQXfNhdo3KMVTaXW4fld/J8U7EZWyoBfK8IdBOqRWFVvcwNLUG6MraAuZyEnmEK
y0Ur4trt9nJ0X4hWIfPOOXlUmwXUVIi4VHuRH+AIFwi7Z/pJ28SY7LNhMrB91qYw
5d11OSTxefUuEKYsnDrT5uZHejLiobRc8sUybpqeby5455w+b4bDWmtV305iqhS8
vkNwnhL2Ute9/PQbo4a2v936tAlD+QQG2H5iC2Svxt/p0CDI6Q3wwCOfk1XrsfFY
GMZA2BbONddBNt8pE5ZfV6tqKlp6ePQB5jvsamDT+yBLImJPgGqt4KBzcrv5riTW
xwOo/1FAL9++TUjjaJBuKWDXKbMjwRCZ8NQ8CvNJpwdg3iaIobax398pkeI3LN4q
1EDiln9/ymwPfSAkuil42iEQHJ5RoKlquKCgNZQ11EhXn6qTBCZQAawDv6QDnhSj
FEXVE9upsaX4zGVoRchY51E/qPwTZ5GfIzrzW2mT14S1wlSEZcA6AQu/NjBRFoU6
RWDC1LU8SSqrMGYoa095ImMY8lupVbWix5d4PdkeXd9JoCLJNBMxZ+eebX7LSA24
/KYLbdDKmFNj3LV6Ftkrsb+4JYjHRXOFC24fKPrbXM1zcifLWfBPj17blKTbgxQT
9QXDTNX1Z3HSsqU+XucRfx4AmVlhP9W55mXZBML7vKag1FJXvlOn0GRajEc78pId
sA+5Dy0mx/LkX6R3SJdfgnk68knGpu92dhSm4QYyCQt6ByEURQef8jVX8zNP9tu+
4QJM20Tw2P7o/cHaoKG+iUO6M1eDBYaAnGkFbuE5r0iCSsXROsQk+NkfooQq3rnW
2aZDJSpEHdz7fHhKeeqIlcJFo0PhouSDfgruHsgIgp5urs3IR5U3is8QKCpYtnMz
UTxxYoZDs0ILfqwwj2Afc9JbEmfcBSZ6U8Aq6S4lNzF1WCnGUMiWGBU+M/NifBk6
oG2V/MyfJniFct6qdY8vByK7oROO3U2MKCjIgLUi4iGJVL8f+PbllPoRDRtdK9xD
wnOmcVNZD8HolQ6hq2cddg0Vy8g2hgJwC2cD3ZucmcfxHsC4bb0UMoZ/Hmc+cwzt
gbx8US17sahuwvs+pIT3ftQk5IPm5ZL0GzVq3mZg5QODt/X3fsOj4hCMDfx0sbkY
i9ExwSaC0HGEcVfdIv9gu0sHHKW2ymLNM3VTCqZL390T8J9PkyRW5o4/G5Y051Kj
DFxmRxQBZeLX+gYqLO4itD9SOZjG4eMNaGdzABXhn1vHYAMHjf53I8ZyAkNwaHBh
kzMZRCO+n0N8dkPSMBTo7Y8j47Ij5nPC8kr++e8K+wdGDJRmhF41Frl3Jf9OMPjz
E2OGT2Y3zuvDlckkm1c7zp2C5bgG20YhVLf5e3LRt1HMvnSX854yOYoTOsLeRtha
EZugfFkb5BQbtXwPV8iqrNrZeyblhKAFj4uiaQS+sbhKqZ4MzprT0J58edMdLR4C
okcemQtdADK2w9qwYIQtnOGQ3oyXtw7P36DMrJXgS6S2yZIUJk+dDLv405HwTu+/
V17MRoOpvVePT+0Ppsx2GQLyg4T+VrWcbW3frqJjhQ3p+PonMoeaLTNcshAjL1ZL
0eqSCI//TJ8CJ2zd26gxUEaoda2aLGvEa3UuJ/nwziyMlwi2gxnPUQiIQVVPz4MG
k4Jzw+ce5GIcCstgPUFHNy4YpSdUWbn3N9FZoFmYNuqEsru92dOri/K/SLI1md1l
I8SbmT5zhhNNz7MuTewOUYrIBg10KjYrdqbAWtVnY9Pj9go3qVJGqCaV3OVgYQqb
HKwep3xi2P9p1lmcMY7/OV1zfDiCYVxUtJHR7giSB9TkEbMvjbkmaInCM80+U835
GpeaSSrQDR52viSdBooRuIuLwbFGBtz7EQA1VGMn2Jqrgd9yKX1aymr3hIfuNmiR
tOdruoyqNJqnTDwiaywmCxeuz3Kfemzh+oM/uLpEG60s70mYKuxx5bDYxczYv1s1
cwuuVvXRsW9T3CfoygYN9w+ho+aggaY/3vN8ROs4xLgurP196CFXNQD8k/0UHGqO
OteqhRDD315YimlNT7fnWp/KQq1Ffj0WyNRUgjpQi8I2zrjzkIQCF5dMGQF3sSfA
9MTg5Owp0RmaVKuZJ2B8EGs4vEPdiuPETQu7kXTDrw+TGkSmx9k/mRtnD5EXYhEQ
95MVx5Wuhy4+BskhX7/g65S1BSDjgWCGeXpTBzEL2U2psrDntK9ktaoica8LSGXK
liKVnKvsZj4pOaDSHdATI1yXehWHcvd4DMpZvo6iVmr3Uxdw+ngafnnUm4dTw1lQ
qrY6sEreeQsOCQu9cepl2+/g0LJSTALXtKWiZkOBOmTU84CniZQ8PvnC4tjKsCOn
/Ks1E7ZAHHliqUeiLy+id7XR4Z/CKWk13lQKuL8wSd+r/y9T/7ftY5+VfKGHH3Vo
qBtOk9y8mUzIt7QjSyZhOHjT8nXYR/VZc/6WxpEY4eemf9Ih7wytAxD1h09ShRCb
Tz9ettL97gOYteLXBjEPN56R/7CcXxkoplrklFYUFq3dxlTKbEuuucL6xoUDIool
qBk+Vc9mI4cvhTGB+POd5WLOkvBQ2ANXuo3E6MB8iWwbFZEbCVrmF9RGMBva8bXu
8MeZLlnnVEux3OxFzuDV7iYw/cg5AXd+UcAxfGmEVqpilzr9u9kSF6IV9ngGlIVq
wUFFHgYTTPnPAZdRiQVPtDnTsF8YfBgm69OIHB52+ICoHJhYpfq69oPnjOAutnXL
KP9NtJRtzKYX+rXMXgVSUHECd44cj1Div/pM7s9MOCr97n8v2dKUjzwZRmQ/PcBw
NfsVO9rNOFgXU2PAZyxJRvjA36LkqImJ2hNyxUlU6lJPFD29mSKIhKRUEER4njof
JnwXkD+EvIsYq9lrh7XkT2Yw2HCZt7Q/EFS/+GZLxDmmk6LRUiOIp983sbLSwE85
Fihm5OMbSrOCYQNhFO6EqHNYt5LKiDVVpNq49lwWTfstLmn1Zxx+uTZ4g4NRRkhX
YaAqAkusMcZ4lLn3FSNtmIjDsgD7QhCnNRQf3LwVjxaECl4a7+vRawbKzDMR5xuT
EmeImp1m1rvZMj2o+OhUJkSzfPbSR51O5zKJiCy8MghMzF7Y5rLbew4ZZdJUDLNi
keO9k2VgC24B5DNEBWT3COSJ5pnu+NU4oEeXYSIyk+/9dBQX9QwI+K8rtyVKRQvq
+wvswbK7gIG6Wa4Iq69rzM3NTA8ocECXnczw8B1P7s0O2T/HQxIFTHEoWubJHTIL
xPCq1YfJa4EnZLBZiIQrsKPOefPi23CkP0wU6PHe0oL5bYl8tuIhvv/pGecwBgD4
SvxxmuGNysnnIyomwzLH8Hv8kaUJXABH86GFr8B4ar66h3isVQJoMgzNFCwHtmHY
REjzZecB9+8K4DGRNbtNDWzwm0C7lA6LrVrU8eO8DP/4EHeMR5tpX+5pTE7gCeF5
QsTBDjRPvspCamxHNf0mCMxSk9Rkq0WB1NSjl5rEHoKRs80QqjEJkXi303M84Wdw
Jz1zP7iHkmCNNItl/Z5L5nbqKQ0TGoe9gK+H3cvl85BNWXTar5q/CVdOYsQBw3hL
ZN8/6hOHY3rpU2J/wpyJV2TYbrnLNoTl7BOZHEJW1UU6aD3ei1Wrw7hPBBciSAbF
3Zfjn/nOnIqgWjLPj1VN1O0ug8jb2xaAQO+dcGNYphDVvJ0x+e2RllNivbR0R9Yj
TEKZu3wue6olEHdn92BCUhgyY7IVFqLe/ru0EwTQndBG4GCN19AHUazLK8tRmYIM
FF+pDwGTbbuvrefOCAiodjUNMGnDauB+ROtzUZwCpQkTm0o5eQq2hzWFDiVAt03t
LrLar7uZkvWh5eAXLkIzcFZp/8dZ05z9kQxFRVPL+ARkJXHncGIfkyZ3tjfrT7xG
uC2jxP1dsg3KUQHjaroi/xT1fbAkQJYDNNzBmJHC1UTS+Bp8OVZce5BSaY6jU5Mn
4zDGgDhJZSvbs5ys0h2SUijIJ9YjJR2ZEytOzPfALwAxh1cEcbuQ67/9IuUXWJZW
nYunhCz8rtSJ2uXj7JNAdZGK/H6k+n+V1ogI8YlFmHPDbMUGbmW/JUEmFaTZRWYm
+zIn30iUGQgIr+e/jzgrZvDXR7TfGHqO1cgeKSTZ4MsWKEBF50nJQY3vFgP6cLgP
nLf5Ls4RK9hi0pTFcES3FeKRnp3g01tF1lNqB5oBShprNEFQ3Vjwa85wfs14pUae
FhwjmNAQnRgQOgSbiM5PS/XyoYSZoMMSktim7rFYJZQhSxgKOBEej3gCYHlCw33I
1evEqKwFYaKMbzdoBWgLNyJm5JRb6WA9FEs62JM4uM2dltKgb3MTAFIwioR+L+cr
zg1aKa72MgeNs5nMT/D7KaemMHbLitehShXHKBE+nIwoTcGtwrj86bV90PkiHiaE
KXZ6s8a8X2KG63YuKZIdkGrfpfIjpfD7mf4u4lugYQbWK8z3Ty0/JTwHS0fNfYRl
XP5yXAbVh8YLTQuh35eOFfR4U0SxMlj5aaw6MNxTruHne1+AOXERcM2iM8uMYiAf
slx1a2USJAYJCXjS8rp3NkQxbpgYoEcfFGcCdAXFOspM6LZWOhZ/wfde8Ye0PO8C
+sOswVp6BKcC3FqkTHCeyNwhhR+UBf97bbj0al1NNjaJTxONoUCypR2jiE9W4Eib
3CMmyWIVz9DtsOA6Aclz5n76Gx0VpJpk9DGYw+ir+iYMZlH7BjIm435k7Yln2wk3
ZNHNvl7rFDgVMVBvaTbV3IKq3Q0afSaGkI/KpGVcqPhTZ97DsLWgXgVk+qo7gXfQ
wDz1lO0g22eeyYUUQXaqVcXV3vJ9R0I/bsGbY3WRT+EHJBkO9WozJNhUuAFOEX+W
102qqyA4A84Jq8eZBQiceZk/D6NaFVi8fUooAulbxl6+rqd/AjjJ7g7wST5xwQ7q
z/aimM1Tcja4xFquh9Z0rw/xPuHk+KsHd8DepWYZz65c+ReG9iVNWyDJwEqvAG7d
UfhFRiYuPxSWeY/v4C58s+xBtt/lJvJ8BYrbavQXSybAwAq6jRoJbX8Kl/UYIX1W
HHGrRCHP22dHwIK1Evkz8bz1jjRzhWSCPYfdoHLHk9mmQmp3oTana86ITRZ5eCoa
4z6gnq5WSmztdr68E/hf1MmNwzDNaDNgcuZKlIFKzEM2+1udgbB4hX7Zp63SC7Ld
nICDF+nASdx37ids85KcMd44hqpMLaI8XY2dDJOPw/L7qxuZG2qcFnC1IhZjr30D
BRuXfr/men5mnH+hSxpnYIFz2GeXt5iY3RtcWC6qYCn5mglHFZfhZNHYUyIyq03c
r2IplDZo7/Z6XiU3gWnx2ZIQaOf/samfZZxSi6PTdCxsBoMUIHc+UHNEdhy8k0aq
OBD2cAGfAMqzvCuvNtJb7bqn4Fgy7oFPMuAggG94P8BRX6amDXIbLgn25TPrNKZ2
IoF4RyR/v8nVwOlkHHgqhbLBLVC8DXZasdOi4OXvO8y6EzG3aOi8rUgxP7b2P5b6
zS8dVkZlyYyQ/I6R9Onkuels11SCHlM0jlqDdby9LhlcyiDD0e7VALiR+1qDuoGJ
XTkONOD7awiT/jzUw5PvEAGwNmeSoPPLfhdWizra5GPgNEqowi0+ew6NOeOVE/Kv
osdCDeph/tiUGlLs07vCoaNS0SNodi43N27BoQ8s676RVvzRieGapuPpABtFAyXR
2RxNzJGNQhan7aXT56sWtz3qmF6a+UyG1dYezJdMZqFMBell6jr4hv3alLX9DVYm
G+/iM5tV5NPpnT30rQ24rUcPcdQfolJiQinF1HwHq3yYUDxK+nZyg/yWMKw1yqgS
q8pxhkr/xwBgKO9Ftk1bHK3Zv0nHWM1ecz0IFn70HqLbOkF2dhCIvVEqzfkZdfhQ
MPflUY5+Ids6SpHo4og8H8JjSPJv4H6W7/beSSqNasrUq75KVROP8bQLkIGR/bjS
gGjjQW8viu4+zIRA8ZpbW5/iVQ5lZvGqmx2Am3aXDos6jM0b9c32rw7h8tEGb1Te
9zJRpJTYD5XUIOvlaGpQIjkNDVlgCIPeINx8tX9tc+D+s0V0487oEevfF7W9X3Pn
RY5X8ZOZH1eJruekrpVs9U/3zvIT7l2YyZyvKELezlhd1XN8L8GPeERZVmJD64oX
VxT0r2VlcPBFlvIAVTKiq0rk4sq2OMCHYOR337SfNBLKsdOPKq4HhTwjNtIzTVz5
eGjL4iOtqCxK5+n8hezFLXtCBWZuflaGXKxQv5T8XNF6Lgn8k0gjkwzHXX9/FRAt
3sriBk+ubRsgm8T4p/ALMeCgx53bNFXd68c9wob+8rwdAczeL075fokuQ5lzrLxr
3e9f/wEJ8ZDq2aU2yCxV42AxwcwgjgXPYW6aiK9JyYQPxOQhehbBIvWQ68KmfPsU
RJiUXiJtz7svj9NhkHynDDFO12JYtiHamzoYPnqsjA3Wt7tnOBoVBFCC3NSSrS84
vwFXX7PuROvSFQg2haUHJ4HWno8NVaEW8BTl9kgqivXFhxz3w/3abWbXVWuD+1e5
T1Nl9ILJ/GciMMGq26tGn9NZWBFAepr6u4KRKBp74qd38gJcWFavV2VeUVnuvxgW
PTuvPi33gOZSf7vXvu2hX/wNJTgQtFRkDq0/Cj3RBH5RMOIhE9m2W+Z5QNyxlWJ0
pDj76Dj4mNOU7fWZAtUKYfjJZyDEkt5h0ojeuVcXM4O8YyoUjAG90q8p9lbyok+E
THPWXmzSyDBpU5sEhugbiI9KZbsKs6aQEDStbD94jjwXU/REpaDP5sDsVOU6hojs
1Siw0whsv6WVm2M1O4Jmyqu+py6vb1sRCw+Q4dzNzYqNuZyXWXnGVOQtr0yLJfGV
KCKnoDwhrjt2TTAJnAyH/LQVMuHNhsaaXSzYbMvURLy3JPcFn2JgCpkZHxmJeFhn
/Nrg6xyUhph7dkPooqGEYuTm4PSobW6uTGfPuRaJyvKEXK3IGkj75xhVP0jW+ffg
xsTTBA5+/VQA4q//GjrRBvz70ww2iEEmlwvguky0SLJULTuY8DH+MKx8WeOZgvWZ
3nRuva43WUhpf2y7eiy+3zT9aDMXejFaq+MH1IJDptVcM5e6mA3owMqX4AqaqiNT
16UNCuVa6uCazah8d7XeWIQSzumVz2QmA/YaJ2M8rBH3Ds6ckz8kTHmzxn+futfs
F7chjFWSrHZ5DEqdFlvTLfcMjDaLmzXUK8O1YJ4bcTQKRfPYC2mhUgOpsi6/9J/D
f5fA4SbZX0Qbl2MTI+792udlluu+VB1DI+qOV8v3DG+VXl8BCtjgIxHP/GMDN3wh
DFp8TvjyEJIKtpdT3jd5SwpNcnscXkqlE3FM4fe6r6wDFghW6hatn4YFx7HZtZ8u
JZ2zUMeWw5JhVM24MjPJp/U7CP1SZxPRZXoARFlJE/VYO3LchaanYHRfvSySEnGL
rLaTW/3Rt8QzmR/Qsm8zPVvotiaNFmUGBnOaogpUxp416oI9TSsUbUPER0t40zGJ
c+7U1L+aKYxgsMwJZNNxXYlMDsuISLJRQdNc8MI8/FVnw0fK51mTEpWBf7swBs8N
uaUbrSIK8qUyG4RAHaluH/OUmKyJyzaOaZZwHAed4qp3O9KUW43e48c9wmL3PlKy
xwNrcENsAP/dBp641ChqWToOLW63TtEE3z1ed6XKgWKRT8Tj3oJO1+RTT9V7JYnO
ZIo8zvWuPvf0eXwzRusP2ONKo3PcBstOxKdXzWXCPOvm091ChlhyLjIwi8RvqsJw
jq4eGMwOm+UuU8vUoKptPgVARSIHRhZo+GO1vjyNvfZ9yYQXxnbg9j1iAWjVlkUv
WxPOwOM/gao2+eg5BOoahHGeVakbifVXryZ7vFz4Re+U1BcJzfXHNbCy1edCv9wd
4p6jz+V8H7Oz6d5SnWjP+fkTNQ1lcpS4e+bUA1TkUNB1yxORGHgcWTZelZnMcquN
D915cY0x6S7MXz3/4tbnQMhvW0rsxiV+PQZJGjRPQ67hj4TZGmntnuEaq+k2bc01
WX7N8FlEPtmOHgcOji6QG7z6Vx5TUGQtxWTLj2lEBJvt80r51H7uDybhJNOci3i5
6NsdbPtCPE1ET8lDl7myASRK+T19vCPsHP0QRAN5Rsz+JvxTTQ3sISgbbS45mTMu
WtegwfA7NS9Da+PiRLJ1/fOPDRfRdX6lGdwKRl+HdZZCZ31/trRw1QGtzsBOtxPR
H4qsizf4o3gmhl44HQysnNEmviX2aRlZDiUqOe7V10mKbgFYqJ3DB5YcYqRnglIs
nprr+87itd1ruM4o0qQdZkSpDZsirGQuufB24smO734zm193/YASslNHcgTYKESa
UeYMNp/zOR97Iq7tJ4H49BcBW+6dX64lrtcZAyEWa8YleaWb76N+ELdzP1misvjd
Nh7nNUgV1ppUsPmRv6UcZc4TNZXZppv9s4AEvF2fqvAHvkrHFjuFEChHHBrWfg0p
RrNwSkmHltPYYPLSd6yiWgSVFbqSp1vjbDXBut8a0yfGP7LRejFRbXPCpsrECGP9
6tQCqeEuYiHiq5EA/cSsUAzeGQEFIZuc7BdeXLq3YaVUNlwHs96DqUzx6HkqT0s1
HpLrtgFKNWQL+ErLx7gM+GuS1ZqWVhTm5d9fFZdQb3sunip46kQxPmJv6C0v/Lgl
IA8l9kkSPnVLCN8VBMdCgVFZBSAs9NNK87+GkeqtvidrYqHhvN8sRHkRKwJZjXsK
gYH5CyHEyOsohQpL5VXfh11DxVZZrgfD5ezatXImHL5mk2l88IDpBdx+0HFp/Scz
QK6wH2+mHHNnFT1wmdsAosOt5zgV4OToNijJqA/6gWXj+5jIJqpxme98HA8Lwojj
8cWeFgpAhhVqEsJH0tj/aJAy16TkiT7H5dP4QBVpeMKPxSGx+lBxV7S/tKDjha3C
ZQh53abXPDDAsMZT2+cmhKA35HCg1VKb0EImG1v+//InivY3SA+UsID4eMUnbKzL
bblzZrkjiIyUDSvZlB01Kw1WzMCpwJzVQdQauV67E/ftSZL5K8MVF52QGuJwabey
i7UiPVj6wEwnUUMqruuaM1RfqIHWLu+MU1jjC2/aZMc1jygJr50KSg+iouUrAYWR
YHbeZ+4gSH716FRgDbVqx5ov1Eg9uSbZic6aQINLhBkuR+Nbvu/MfCNi/Nnfm0Jy
oPAq6zWXUzQHKBBFU2dRu9hC3SfdmiZyzsKn2NOmqHmfry5AZ6AaNUwG4NuOnuXK
V3YYFnFhtmXBRMldWQ7/9wHK7OOSOdOqyuwBh3P7N3xyQqxc9Wso1aFqk4kSGczP
ncoLkRneRt0U2z5ESiPTWpS0oTnwvbEtGuzCy4Iio+KIMqQMuJY7guoUWvpN1KVp
8AQR9gaAYDbAl9IJv0QBbhUzT0B3LQkBeUBbJJPRhXxGU54C95CXTfTSXYfAvwNS
bTIOcoaTe6blrMLAitE15JPYFpCQK0ZKJYdNL9YEsltPL+Jr9BkSidUnlIdC5vRi
26ZOMWEPbeKuIRYNWySA0pKWcrLxm/sGn9gBGY53vAn2Xf9mYAtfbJl/4ZaUv+3B
WWj1G6d338WXHvPtEf0O7d7hnNdIUC/m1BQLn/8laEVUB4vZhcWtNKjtYkBZjS2P
zNRUTIxcBJPFE5gA6Yl3Q2zsPY/wBbbXDSug6/wdYO+tX7ETHbjAxCxs2guf2sBo
auublIVs6Z7MWW1s2R7kbISxe1R0N+7z5McyeUYG6rpcW2ZTx715FWa+3HszZL0v
zuSxQThxyLB5JorXMNRAX83E+/b9MY95zmpNL3oIxoEa0jDK9bA0aiCDTh9fHaD4
sgrhuCk2CoP10Qrc0zSrJy9vuUbI7Msu+9paEzVDVo0T9Spem7DZIMKvFSWc9JLA
DWb30gNX+9Vtlmem0Sfn97DXVSR3OaA3Q1gFVYjJ7Nyrs5/eYxmikU3f2wQ4K3K8
z/+0qFG/2Hq3yTcpXQ063ThPL/fR6UO1f20BrK35lXvd9lTW2P6+fa3kKbZdO4mq
Dw78GRecWaVhAeac8A9GAgjF+hv2yka1y94PDHFgax+onmxR+DHHLrY+B1SSEsIs
Pyk0pQ24wabF63DCNnyzXGoCXUIbHJFCHQ+AuMk1CirFUVgA1C9UgS+AhstUD5FB
LsRTU976e7fAxYx1dD2oWbO0ggo74WvwEoIt+hO80NROFQ5AhhLc5YsLVOX6nTi/
qIYyokytSl3lkYMTQdmX74HJmjvARkhn0Vpu9WvjM9NT/+6vovoquSo+2WjMwOg6
pLdhqHnMha91eWsZ1NBR3L+K9itcHL8an/mpLWiDkKlATHe6c92GmoS3XuUVOdkO
VWaCFbmI7gFWCSX1p3pgK13aNunmlWrLXMfw/8Io7ckeE9FAlZQl62jMSX6vy4Xn
THHrr5hRznKCWVPHiUwLUO467gg7uUcrJYDsy/nhBA78DivM/hO31ayPIWDypOV+
y4yueblPCP9cZy3gnHktVnFRD4686Q8Rk+9MXWvGqc8lfOAsnO7g4SsBY6JzRRov
z0V5BH6DanbZDQmQaxi+1TVrqNl+Z8XuFAx+alSUpiCztCyNIG0h9ipseMZYeCYb
zh/j3MlG/3J5m9+NYkFW9EstPapbmMAkOcqi6S+C/B3Rqx+xpDVZRXPjSqQblZud
7Wn1ElTk17utnx/vURY1urviTw0vkSgRos4Kce3smfYMTsHTatnh/OUtkG8maDsR
xpiZzgv5yXqUL38uepyEKMxJg9UtnobTkuD/1ngMarN0nNe2zWE+UJEGnqNYtoaJ
uaGMraXzgeTcn2Z2PGFxOzGnmI4iNmnRAMFujHG5kY59d3Ra6fFEUb+W3Q0qJBL1
rvgkoTbUyvSXDRVOt3YZrCoZi/KsnbGdrPM5ps6JH4gC2hfR7+6RidP4tLzi+g9f
zp1HPnaHMObisByEn0n9S7PksIopIOvVUwD/19YM14ompvkurLCoeusjnVfduj7W
c7KrsEjCE2uqQTktZLzdrM2mm/9FsmEclvCwk2c22zBUbOLUyUFbTVQCtoCahUol
NbLV0doyOTSIrn74daskRwCBzpW2WqpQ13CuiK5P/qJ4wZQrPL7BZTxnToXwiULq
c2cpYVnWHzQFuAnV4hr/14rcYLzN41eIVfvMl5bSDPlxX260nBds3smcc4aDy1Ge
cXmaphpcVDiQ1XqABieTKdateYAYyqfXPjBBQK0QshHgOtkI+x/jx0OagVDfjLA4
Itu7RiAdCzuGN9rpUzPIG1pYJw1F3nCW1jru0ueWxXAkyA3gHTbiaQ1BY1fOeNKH
RglVDHMPP41OYDnthBlFu/clUViYreDuj2Hoo41h0SrZtZkjQ18ARylZdeHpR617
C9CV+JFYzzgHD/SDl2OgOLm3d6umu6qEG0P9jhY/qVnxkRgrptEHyk9TDphXYy3W
cP174dFdTGmr5u8Lj1ZagGhcy9WEiTzp5vx9s796DujUPp8twYJU2keELhihtfQ6
dXLCbrVQXojyzeOqlVqnAm5fMYMcMyyPY1T+V/+N7nyIIwBwPIwSK81D/Bsi3YXi
nng25/W41wLeAjxysI8V0IXPBxS8ojXw3yjWrH7yOa6B9nDS+qnvjvobkq6w4zt7
dXMOuU0NUb3hEeqruf+Hkeavv74fwYBms0wg7IfjIcfqCt7JJMF8AdJ5o41sb/D3
vum8WrqSR3bILGmvXHZXbADrT7+MalMfsfNw991NiEwCytO7UN7YBX/o7cCgN+oA
a04RwXDdpBkudQOOES2jPxM6QR8u76IUlZyaFMa3Sp/9NwAjqRhSLRZcaaPORSkT
nwm5mxOFIKh08chcUXcb6KqKi2kVgM6tZnJ53y/hWj6nHOQbJV3Nzx3Sm2NKo2CQ
OWqqFNMKvskZoF/g3kbvVOujpRyJg2zuVnlAJXOlzT+7tem9gyDO2VP2/zKSDOwT
ugFWudLv+sw573XdrLf6/MlzbesERrczvdHTFgf0EVWQeWjyRr3F2x5eiBp0LJmZ
mIrO8nY89kB6hNFFSDkhDipUnxU05/PZI5WaX9w/NFBPwD3oUwpA7zeNFyUCqycK
6gELzsudM/rk32MHzeSzeeltZ8xwnKS+KceK2HBtASTPJr7irl1pOv58GlimggWZ
jF9YtROsAmN1Q9VTcA7bbULKou/N6NV+k8fTGoqkdS+Yalvj/CI2NFm5dbnoBSHr
F4udM4N+2vk0p6n8E4oJO4PwUw5XDY/v8nlDHJXN06wSIMVqqd+GFTaOYjWRr6le
H7gqVSN/GbzqL+Fg/A0r1V1RXHPPvTz36KWJC5TQwXsjIFO7BQCL7FYJhG0f+vFK
gYlEJHz4tV9lfD7eBa1EhdH2W4a+kkz3f2pwjZB2k5X9PGjFOk0+FTL4SA8hyNdH
NP6PVSAsFdWIhTS0EIBkJT0D8lxZFglGZMzbwq41488Az12j51/81IS1ceovfTcS
YiHcLokgvp28xaU4TyDRonHZ4t7qqbyvU66M0I/qYLs8t90O6RFGVTXtEBBX5KM3
+1XJgLnVEvUfXmyLge60YmDNMIhuZpi6A/fQR6yaOmCook0i4yOugKit+zWAFfkZ
SMUbHgF3XUlbpwMfInaE0/GvGfjFFMmL3tW7m6BObFx6dH7m2AX9BMWVKRUkF2/M
yN44+nP6Z+P/rIGPCtHneKSPYaLHIijmFZk/YdSD14l7qJUr6kooj0/E4xxVj3wN
F4z68D/AbaNAkpDnQFNfcgxBWRlSVW9tScNblZIPeKIdgllVrON90vXs+Ug/LOMN
+VG/O5tu6qw3rBhasac6kZrpzyaYZam5JQqn3+SnD0/zsVUiaZRusD7WTxgNhne/
KivWuA9jlGNzecPhoeyjIzSbIiktEQxX9uJYWUUtQ0WhZ6dqtN6LpqbsKTByaylQ
K2D2nGmaPW9fdHU2P4qexIWeGxB6ckKdvsEIstRizHbWs32tJDh/PLwd4ZNkszyE
gsB14lFqKfYYyqFt6eZwz6wOZrJQSIGCl+6JOBO+Smxzbj/N9GuutglXXWclnTy+
ieARQA5gm/SnTAp6hfJbqkw0ZWHKpTQFJmettfFr4C0xg41guZUKxuLQmA8qyFU3
iJgshPNJY02RuSxml8Zrqy4GIgckSxt0jnKvqBiB9mNJT6QhC76MFK6vubKKFkXO
cj2gGfIQYxO3act+SHS7Nx6yWJ8hKQrHzuCm4/sdWwSgnfiapaRpIJ3pYZjrQT0z
8AnnQbRD6hVny9mfMkP4+v0fscarH8GcF+9s2Nboavtu94S4Jm+hOXgLubNsT3Y7
eh2AVZiitIn2ABawUV7siuhUCaEIbXErczVWubw5d6MY13I8dRVklnzoW43FikqS
bJgFiPIJ916Ex0EpX7f9JiIeoI/xPFeaQWBWG1Gfq5f+qsqkSWgCIm3vNNxcXtqc
dwPT5MQ0IOBBnS/quM/mEtiyRp6OCN0sRi4KD19zzipmxuS9TIExQXK5fbaaGupJ
WAn/ye8sjsajZerxQGwYAQ3gesh7MvWhGB50iVH+DNLwvjJnKYRh8H8kJ9FCIR0Z
yOr5Ft3e78lI1JffROwN1AF+81JJtPKHE7xtmUAQKPqZKYeEe/f1dCduKN1txG9G
JqZUqaSCq3l4IyCB1/SAHsUk/w4G/izvsYPZGtYZnO7rCs2/qn+5JjNgX4EK8xEs
weR+w/SSLg4D/i/SaKhX/gh2VANCDFuFzpg968Zv15zXfe0n9bjWeQjx6EFqkjjs
9r2FD/Hrz8NL2hj7Yo9gAOoo0Qj72pe+p74CJXiOp25IPzBjZWW8gh6oAgJL0Aai
S9blkhKGGPuG9gP7IyW3UZlrj+Tdg2KUXxZnwTCYxlQ=
`protect end_protected