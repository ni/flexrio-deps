`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
hVdJHWSfELCmA4ds+csnOQAALbB3ps7EiTSHEDd//nts1r+JQrRE4d3bDPRJpiX2
Sl8d+xAK9BIi4i+3ruAzYvB6kuD7r+gs02Jsvd/1kn7JYK4xBxCjtdDFjVHOTEl1
sSh1oNiYUwLuwR1yKfP+xBhqxD2Dv6pCKhH1NdGilpJQ6cvivGkSunAu0tzP76T0
4x1pB179E7uIeRplfHWX03KzEBF+eVtfgXVp2W1BGjfAe43y1pCvNYZOh1+TY62g
EgAFgbo7pAujZxZy/YSiZjUr2mGp7o83qMXyusx8+rQ41D3X6rxfuP0RiId2pOpC
6oq5Dfkx04a1dk4s8w8cVg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="Sm9DkM+kBxuxXCFA+l3fFkxuSWV4xqRc4Nn7Ji3ukao="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
m2emGBqRy4AuduN4dffN8194qYvc9UXRqiQc56IrQYMiIVQPyh59I8SYabcDdspI
7AFHnvKD5YaF6tQfxWm+mlcmMEk2Y//aUjxeiGGs+RkKgbHitJF/K7nqg1dmKvDg
a/GaBCq4Bqh0EehlN4ntP5HxM4qcvSfh5m/Coe3drc4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uG91daMWA1mGkhgP3oZKMYye3UAomMWgG80HuuXg2E0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23616 )
`protect data_block
c9NqBF2D1wSep1rW7utzHsk2j40aow1MnrccxUTvKej2Q1cyeDDbgAml4eTSXI8z
QYgCADtWi7S8BeChdv4B2VxKcS7CMq/DaQrOy1MKTfQzfAlK0iubmlTkljLy0Rwd
UXlwcea2YGh8B7b/87H7IBLDLePtnjMm41mYSt8t26OO1Bp/oPoN4Lh4i0CJiJyX
ihS0Do0d+Qcqiu31+qMlEWK8EPby+4DtVWx/V45Wy+Q21X2N0zuOo2GGbxcKTDii
S66g9b1iR78n3zQLUHN6Uuuq7Da/8Hgzjr22tha1/DWnjkpk9eLE3PWM3JLjCHkL
hFSXiDW5qQJ6tdUh3qBf3cQNJHuTLNWaNvqvtE+rE3FRojLnGzRABA/NbPhUac+M
sdpDn1KTu8+l6kRQa0QULPi38TWbGgH1S3QAPP6XpkIP+SUFHwEwTAYYfkcs8cIt
G43R7G3/QlAaIu6+BPz2rMCHL4MdH0hASj8VGeBMtFJ5vtp9/IjNWKE5jGOQOl3X
R0WpCfUpxgbCUUD+IPtb8M+wW3TDByn6A1ysD0RuRx+BY1jFbfiruA2lhie+lOUf
0ym0jMC0A2z4a/qJtmaMt8GFvU7sLlVsrnRl6Yu+a+F8oJOwIw6zzeUlUYJ+CS/p
Sq3xPCGqk2N49VZM0iMSFffUw+9xWwUoBm7lcM8/K4nuKNOcZj74HdbF7cbj/wNw
QUGlsMmP576jc9PPjdLyf0Q+TUFkHcNj2zzjr75omqyMdUZY3hqfU1dfTHCzITmc
Rgw6iLRcUTuC34zbYEtF54rVfyZO7ug1373kG5m3xZOnAmy1k599XTdaXR9mN1dK
atVA/FwbtN3w2pIEQfM9JC6iZtYF+N5jlUtEJHPy+jlfygc1qaUiPWyREEwrWV6v
ogfktkJVz9r8nRaaAJ/mwzMsdqgMO7b6Ozze+HlW5IKsna+oxzzn2s1T7IBJ0mkh
LMdj41Sa+4esS+5VhWMdMw9U/JpNZKygsu+CSpx9fFAMGXkGW0ozRazEe4O4VvdR
UnDod0ts7nCrkEKlkcXeXcMW922yjQdH3LZdqvCVVyDkwqbU/cNQM0+hLuUUe9l3
wHdgkbGCI3wemeNQUufonPoTGLjT008Re35wnCPocO6Ru9dV2H2VHU/J9UTOvSEl
3oo5E5R8C+hPBiStiiGQ9qXXgVRYT1mcJJGM42IAaXTxUk38yCadgG5WCbsmvR/Y
fj+lWzOuJfFz+5yRD33WaoXsXze2OmSJtGAt9R/tHETmRktsCA1I69wq61D3e1GQ
L6oJ6AW240xRl3klTPzlLS8rq5fQWTN59BObSEQjLfDA46zu3wDLoyopNcijAxH+
4T0k33TrCr6fS3/h3xOzMs38Gh1owTZxF6ozkkrCPec+xPbFU+NPeoTOJYMRMYok
U3T3JV7deVWalpFUreNtqo28ipn4Ra8HEoou1ZGirEB+0ypLvG38QuyBw+VPNI4U
u7wZF8/iLJTRrHJXwxn0gHft9gcroYEeUit0vHj7nCUFpBIfXig0EBUmBRTb96C4
3iwHcO4PKGWfvkWEPSykiX2YeXXjxK9T+GgX6e5hU9r3mR4bS86uKUD4IbwLEHNH
17VZSIqSQX+oe3En3KtlQUzgzn9BlG9q+qLqAa+CIfRaIuqSOi2K1RzhwmVwf4bH
hI/mGRxn+7kiXsC0n8lLvVSY6Oeha0igi+djXuCcAZHMA90eqf2kEgFWA74jWtWI
Z6SUq3MI/EhN99HdDUTviHMOqhyQMDI/Ph8JsHrf5g1dM7kSP+HafN5fxVM5Fp6F
XH6ewuq0nDTLU548DpvDBfD3SuZXXw4V4jlH8ml8eGGlJCZihy27jSwiAj9tF9KW
H5u75xRy/tbdfjuf7dfK3CFGTObS4HcWp454XGDvEeSQhClsQqUzCJ531vXiqCZ4
NDsfzswB0W5ZG8IZ0oN4tBWBoE14Qv0I28cUIqq0usLTMTwMuoVXE6nZ6NsLX7rq
7fTDS9TQ4HG9wzq2npTRBx9mZA07wC7JgPm115IzAPLE4KOO1gATmqpyXxNypGZc
ewEvyRGSw/fcUJDNJMGutCCyqneGd+IJmP1g1zKc6bTQ0VwXrenHT5Bljxfmg84I
Om+iaEeSnEegleCYsEVjxCuwk2wpSwPL6kQ80g+XuZruYvpVKkfg4eqInkCYbxVp
EVH3qXfxvU+eUmGkR5olUp7z8pga040tGQ5rqC0hwbAkvVgX4N8HuMNPZrg2LI7R
oXcUXNEhn2KPQR/kg+wM6Our76SltkXeIgm2cQKks79FIUtvfSupZUFoynwB59TZ
iChoYY7GWyVE881UZXaD+iZ6rh3BNTX71Mf64nGCK48/17ezFvd1BuVG1MvDZVl2
ikqPBl+jpTsGlp9npbBQXJabOdKQuzWORLu4LR5960Doq2gpQvqD2f+uvAWPxliL
H4aHUGIvIU3oTDGPkMaKPfNEJRAQC6DHt/7uRvsdn/F7lRNZM0xk1JKrl8AIabc9
6hGuapNuojrlYEk5aZ/iWHu36Y4Cu51iaih4FaAxULkmXOVdhQ/X2Je2lT8sX91j
ERi7MWoRJ77OjNW/tC+2i3MI9VPxXKkgAKlqsvhQvJW+5HyAzP4QHsITcGiPn0jS
3L8FUlwix3zg8ZQ6LFNrqHs/+NaQ0KgfbWzbA+97PBvHVJZr88Y2M+cQzl7HV20l
/D16EdHkm1hIyBZCnhh6uUAS55UjqOUN0GS1yCYHLKbfPA07TMdA21LgYd2DeYfs
1Oiut9wXWT5SWVcqhHgjmNRqD9dZKKohcQtnAnjIriSlidORf5eTdwcViO3T4Vjs
kZUbtwxrjavkBVp/KPKEOvhRBNG1yU+8KoBx2SPFPn3vVUDXoDVdAhYVCpOZrACi
7b6UHlT0eqhgBUOFblcbXQ+t9ahNUjUiHQw6mBXhsdEOEDwSa9SiAbhekALWzt45
m29D9JdhztsLeYjwu7j1gJMXch/0qnyrAJgDtWFkfcG2ijTxgtF+/4Z6z3SENp8T
6vgOTx4ian/LIjtLvcVRQOxEZ8q+xI9VqCAGzqJbpBIGkBUsOg6XdRoWnJGEOHaV
8pwcrdkw9rlLsDkt4FQDCcfEM/iQLTMq+jMBILPfZmxPv1rVUvlyxMmPQ5PnZyCD
nSLb/jmKrLYPHvDlBHU8eJiOd8puKlEOS6aV234kmxc5shKbIz54yHHLI3e1VT5O
08Hd/0YoP2yXlW6REM4sE9LysDTSSd8BkugVylPts2sgAtCw67gpPywt8492vAei
RkW9XrLfb8k8ihU/dABpl7q6UeoXYBfIcgOM+BlIywzuzuuOuBuJ9GZAsREQnkI5
Bxwep9TkymfhWwLuLOzOl/TkG0QEG5S0xN0DzglJJD4m6F0KZNoW59Fk17/Le/Qd
fUDBiC9tOte8RigxJ5JHSGrUWf6Canh98CLxBKkPZVCQi2GPedT8FALf2MGTL51l
d2hTROVhY+aZQDldY5si1xtlbrcEZPduoc5jFwnGLw1VkGVYPk7UEa1ryWDCt3Uk
FDp9W+ynw/+np5Tb1RK2SsSQTzAJpTSadGlJiDLr6uw+1zxsY+e7teqJ9FPRofD+
K22eLWC8ZuVc4heaO5Rpa06wOBNnt5oEFvK/BXDj0uUVrDEPCnbKHb65opV+Td5Y
1VitmwnMfJX+z51bI+8x2eT9I8Q2fXNkDNZ39lCSWU9mODbsn+/97/oPRiPT4bQr
k0ODq+jY4HfPrF50zYtTSeQb2RyRgiQk66JGKb5DkPu5HzfioLt97B41carx3vGm
//Du0VwgqfYwBokwHH+XKHIi+/+qPhb8uqnRVW+Iz9CJjYFC3lsqsztbCFordacE
sh5SQbqhi71GU2xtHXhd34Gh72Z7qDiZKRxaMR9MtCj307FEUGPEwL7nr0+xpk24
9tGUME8ocJWR6Zw7ydcu9/Dc6lvHnrN4EeOHZVZazrauAg13YReKrcuaSgxp47au
O7CYUkzvX7n/9O1n0Mpq9UQ05j7eo++0wc11hj4CG175jaWj+ahlSPtR7ut/0pf+
8udq7R32qZZ80XsarrnXc7oKjzNwXz711WpQe0rmvfeGhlzIz0hp3sbFpN0RutbW
6KOAcizjzLOPPHbGFj3jbdF10mKj4IDg7RMs60FFIXvsl45X24u+fxL+2tUz95Xu
fHttgFuZsJ1JDgmpaEk/mmnT04MBYiVrgYBcXG70G/Aj47bg/BM5AOCeXnSR7k3/
vfLXdBQybYbrJyeWMti+KAD6ueyeGnsepv45Ly2GCXNpRC1ppi86ZQWJrHmvO3yc
siOA8fBJiN6MmrJ1ymGrdzaCcwBJ4zSSilZQjRUpuuYC4QRQgCATD6HcNkW8fXgU
6mV3/Uqcq5xxarmdABRRfsc9LSKMB3oXiUPBVqfuAhhCsea+nr/NBLT5IIsSLWLM
Wdkm89Ia6QfkiTbEehVWVrYfdBgEwGewur0TAy89R7tK1wqLMhcdu2/dQ6XEql5b
6eKYc4R8qU1saBPEnoBRNl+TE3abck0R6W1vhvlSI1tpS64WbYYi7O3hp+HItjE/
6lg+t4ssE736n27zY2bTK4hISYF9cIfhSnlByyKRk2JriN1ol9mkoRPgm2lAnStb
h363J//TSgmQG7lifzswcVb7wAAExhGVrPGCBbPI91ygrV2Q6najX7G5N/bjB7gn
E8ASEITF6cWCBVpvNaoOUjdhHZS4rXOgujAL5KylJloyYWNLjFd0fYyZS2Kf9BK1
5i0B+KZtuKz+DZwoiG2lukA/neBNkwBX3toECd8LNrvd9uxe14gpKkk6+/dkGWnT
9wRKuQo+fM+P6EF2m/RyjtwFzQqKqqjw+BqI+vceICPZum4imDd36HHACV2J4n7N
DLPhRTgsP/+btQpml7zc56hlrU84/eqpfgz7kVZdD581/KrHhxqpiKUlLiqEwzOh
QU/17uPgsdcM5CH6CQHUfDtj8dG1zPQGsaRBLSzbEcTh2oRsytIw8l/uRnN6zvoE
pPtGXNeHhGobVVxz6vAkgo2JK6EZoMpxYdbLKtDOl6nX5jXx+dQKI5ISLajxsahz
RnXgLCm6l2pLNgVntcPlOhyRFW6vuQM0hrEFo8jPUFAhFUUXfBUJaPVcdUB52yRR
PCt1s+1PkY6qbrKy8rFVHiclA/H08vKefiwdwA1HAgVljPj1/ArYFN/+d3iPooOj
ua/8TZg940difHt6h36jpKzQNL1eNRu4gNmdn0TJPgv6p9EtEooPagQHX63WXQhJ
nQW9LHCQmslNfbwTxVVlqo20Vl5eI3NzbL/oxUa3YNBLi1pXiNf0/agQMJZB6leK
0C9UwfwEeXV16DkXO68X24y+WGKRZuKCEnJWI5tMPbTcQ4GCKGrFICFhksGUJmrV
LrWt259OEuv/OS3CFFhmpgXPyDP2w0sF78vEDluQIcz3V2CoPHXJ3U/gVG7hltpa
aCymLuFE6z0Cp5Gq/m2eyTjjFqFSUEHxg6M/zXCX6boeFlFEjBaWAiWufjxw5Z3K
xoL4ONDZV1iY9BwRUSrV5WpLK/AozDmRQGYSNAtivgI0pkJ3k100yhOpskG+Vsa1
UhoZ9exUQiS5Skv44lJWXnK6MbdJVhOeoeSUpsNrMrx59eLLHrVQWLRosM00LznX
QPBR3F3aexCd+d6f5wSPIi+4QQqYPO67kvK19jPWXuWsJlG6A3aVfKaSsqskH+Mz
8Z6el1kcjspqY2xHtB5gFi8fgLxtGB3+BiR/aVqlhCDvN0Yg0hpiEQm5jA6LNJpy
0xv+pAZGqUm8pjnyhzLUH1d9DWQW+rPf8rIHXo1ljx8cEsk/TYcSqhC0qvbqM2A6
qx9TnDabT/Fdsa8osibqAsU5ezohcn847eUsqaMJT9M+gviCbhYILm4p+IkRV71T
n9LHPzvdBFPuAecYjHQFmk2mPk6Z2Qk7IwUcDW1PMMWEVgAqdVGApHNkrrGgO5Bm
qU/NJuherv35LZct+sdWNQrewy9PKWugpLMxq4dDI/bPBU4wzrmaD/rTU/dEHB5R
eIm642N+58gERTXVATJ79QewWznXubq6QJiYc8px8CLE9d0fl6WXBu+y4EJSfRJe
PllYHBjERu02veF0ByPDiVt02LabUDNuO4W4F1edgJ/JC33cmGX+Wanu1Hyx08S4
DiqzO5yUFbGmCefnNc2X0iJt4eFssCGKc+3ThcsL2dyNWSGxr0BFj3xy5aeTpz9Q
0jJeGu4mEl5Qa1vQcvDXLWIhl6i0zsyUsiaQ+AOlcwFIhbJz1AP6VSykFu4W2z2u
dm7mHKA9PBSdQEiI9f/UJVhZCM4SfZOFx0jY4iNsHdMbeGd3dap/1dUPeDbBKW7R
pAaZ2QhnY21Eh4z4Z310T7pjJMS+ZVzg1VUliMe1rZVUp2ozwVhie/fGWi2q6+fB
J74W5DApNnpV/roR/mQuDXViQeuKnKi5jzHDaIh6ckLfe7W+CylGgYquj/90nTVF
BCwbleyF81nXrxZpfeQ0kkiGDj8KvFDxCb6e6VWWz2qmv1V/mE+7kku5hKJ7VwOo
D9RKC2n/ac/L6IcuslaHkWTJT1qkXHpJCHgsv4miR62uIxo2unPvlGG7c2PSPncT
Jf2dCLHx59D/rWKmhTEX9MMxQbk4O0w133Wmem+30ZZinKRzyWWDJ5JVef2mXrxD
ZYje3h7BZ7IkhhbIHYr8bZ/kE946X/ZONqsOc49N+d24NQDvaJQyxc6sCsamAsis
OrqNLm+sMf387ycllchq0VGVQ5qzNtSX7RSjQoRl/8ACJKu4PefX2aqnVwnXd4PN
LgwJNqeZb4cXLqK/0N3lIFstP5zDxIZI+SYJwNA+gFsZuUR3Wt01Z9qewq+3Augn
565kmYuzrQH9XYQFau4QAEmkQGJVo2eSnnplxY0Q+NxvU90ftb788i73z+ldCPMc
nwKWS9EjCx6BKt0oc1huGQvHAmHJpEm4EmCbVsfg4mT67el5lh0yVDaQmETVBlH2
kwJcCqy7VknfDoYxq+Ya7YOAhNlFgM2aGkNHlU9jrDImrT8ph7i4MoRgcF5LZdDo
zpi5tKTjcOvnf9MuBaywxLoWYToWigNJB9p+yRx9hHOPSbOfz58SVh3NTk867ysL
xxxgnWohOmfeubI+5Yhe+xPscUAmjNkWEAPgpCbVW5X5ynRAW20mFnCf4Adxz5Fd
wKg5exPScXv5NZEDAm7VaCtoJ5eFJLtd5It2gP79zcGF3LQpls9HCtN/GAzSBzq9
XGqHZbjttLrYBqcxqyNJImpmF3ERu79n+kk1RzUBolW4nx3qnsh3CYam+sc/ZzzH
PwtzdNWJ25PB59vSiL3XOnjjRgN/Odvlz5xCtPkYTvLVu7+mtovFesTf31hY/5QF
JWZ+BVjDQFjWe4JaC0RWtqka4dikb7y1g78pHIOMqHLB4diLLp9T7RsUG/49jlPQ
knyoLcqBs5eEgSz2OqdedupG5DdPNu1nh3zR+89NYEJt0q8CbJdlrTw+3UcHr+gc
qgB+jDes8IAN88yWIzWPHgBUlS61fmyXY+m2AXNwx3TAMwkybzobOXJ0NRxzlOQd
vU7kukT1s+QyCStli45yfOWMv49TH6AXHzwCVbocMVlrPz4oRjFRUDdgXmEWPhDe
KHH5dJF4u+FByWWZgu67XIJIvHvZUI/BxbOptN2xpwZjN2j4opobvhNO1KHFybdZ
gCMf3qTvuxkypitqM/Y/xHB7bE4B7cNaBRgyeKiLVshhHlSVwOHAzF70IMP7pM9u
BTfoe0sHyuZBqCsNvlOGQ0/CexeXTSauT+GTKQZEW0Q8JjedxIy0L2ihTFWBlzVH
cLstflZEc/4e5swuC2BbQTlVJHP3HXHnrCX2upikVfNVYL+ojOqyn7fFlDjjuZz6
u/Yz5zhw+PMG63RhyTM6tsp46JFT8xvwASTJOLhgOmVTMmnUoRgpySPvQlVSN+Wx
Rqcj8lcSkXqhKA9yTthGovg1AlRISE3IXWr1pmrQkW85kbfFp6vJo+a2QrzbSqlZ
wXV3M5ytbOgl7jMwZIObdDoXxsBF+Fj4x+g3GJv7to77WeemfkO4TWCklyEEFZJY
X06P3cXQkIUIPp8m78+tJNrZ/Dwxpq5KLcBB5/hoIXlopuYbKkcf1rXl31qO6Jj7
tbP1eLz8vu0JnJDuwTH/EkEJ8HrPebUQj6jzf1foIy6PuT8GSOnxRiLI4xZhI1++
vb0roBo+rewMCKPqb0syOwsKA/KtMLIQczZxuMWREM9zVYPpXgMdCwdtsn4uBPDu
kb06o84wkCOaKiQIgLwphL6BxOy1E2ohT7g9sNNvHJa2gD8rrJAkfIDwj7cUNeV2
/meist2mmPOAahku3CRqQps22znJb/8fsEX3Alqyu6SfInwmcquHd3SbQNKW6l25
CmxaBQBpObDRh8BYdy7JDntuRJiwc1Pan0FY8+cPXVyz3t6dMRCDly2o6zAev71E
b4EiNSdw8jZi7c0d+wVl8fk72444UUNNP0qT6vw1s5K8qUysgxrbEoUjIgsWdFwF
8qMW7Y8v3K/IvxIyfNrl9Y6pB85JjGYgOg3xaoZlsd/RH/I8rvUnqqYZ4vZg8DuN
d1s27KoTwzrg4RgKmLspTz8BAv9k3L0PG+VNjqamXTkef9Ph0o4PCOnb84OYoZKA
d+ctZYhJ1a0ioj4FO4UDsNW86PiLcJM8PsyguGlLqsw4M5sPmGOrSCBj1fOf843M
dkm/yQOUbkG687KQTbq95/vPpPkx64XGt8GRI6lh8293XzHZOy60wgiKOtzQ426x
VqAnfQQEUsxj5R0vz8/tMFZDorVH0uRWJ6TnOuxjOX87Tkk0Pbu7f1ts8dnLmGIp
LqJBOHWc0kEnAgSoH2eohTbkTYJE1apX1pUy09O4AyVkngG89gc1DdkIen+4bBzS
KdAYJA3MIvASS8y/N59Q0Ep4pzbqzo/FvrjG06YauWpZRWY85H4bZ3KQlcjhcgJk
fG5elX0ojeWDtKt4I62PxdQbdtOdSMqKG/m8XDh72TTO4sAYWpy+vH7tPbcb8rQQ
e8YywJ4Hdt8wMU0P+79I/siLQv9kclc9Sz9h/RAb5szwknkhb+wO/FCMkWQunB2d
kmFMk21TmCWj2JHYRrNdZyN8EBNCHN3G7nnxKR8w4HNq1R4XufuN+e2juTTEU1yz
b9UaBhczG7m4AdumpNNMTdhoC7kkfK/HdhItYRC5NtP5pAeHXU/12yZFvaIshROu
2B8jC/JRe0acbJZS11Sx1AjJn3a0GFy8kjaXACeqe2wUydc88ysYs9eS0TS1e51t
wAOK0TqVKtMK8jzoNv/bRCFu3zDdIq1AHpBAZJ7asp1XUE6S3/pLFrtkL5OOullT
xlSHDp1fqJXluLHibRVXFEgFeOdx39fbyLrsSNkOnTV7bN64s23glXeUQ6PTmrQv
2sKrHd8LBmsTUzZKAbreramzIILWpGWv6QGg5k4xWamVcHTFDMGYVdRVZuj8oMfc
I88xdIFmKKSKfbZjDlMUYvaBsMvjR4TWX6U5uAeEwC9QxO46ubBq766S1VEzV+mx
e9FKyz/qoJzNdKHIwLXVr4JhQ6Wh3M7FIygQadslufdVdivua0TBpS59aX21LL3i
oMrHxAt+2sBLktH+UDRIpc1KRvHNlHl+iReaLtlIYmHLS8MFUCZFAB+ZySFPpnPq
aW+V3dTO/1+jGo8ynkC5J4V5KQBZFerq+9fo3YsF7ffwjlh06VSDgSKS1flim0HU
FqXhP/IBg8HsbyLKDNmL4vhqEQVSscVW7NPkcKm+DyU7XA7cx6lvW9TkMmtWkpDo
W0HvqCsLrhT64eqW9cMuOgt9r4FBBiUBkBH4LHVdK5ryx9yjhziftgPeyzQX31xc
uoa1BAEQlPdxU2il74iQbaGsBrMbwonB9khf3W/3MXf7R7ZZayn9T299JmsCOUwb
60jYXSVkQ+KRrP6IvkZdk/Wj42kLYa323ZxJXXW8/igOrpPn5x/rd2KTpBWELZP2
RtJNLaFxHdw2LUjq+iZNoKQrQmwljT5nrlawssCH90cnX980Ly3oQoOHaavLADl7
CBoYPkutEfElSuT1sGrscovuZEyMRJb9NKgydLvUKLgEgPBYchCMx8wVkTrOn/0D
31i6SCpWmZ1K1isqvTf2vkQ7v1uPvg7rqvwXSwnjHDaiGqDraGHMpl4HTMd5P+pi
d1VKrFFCBMgxMocAOCq4uT3Umil6ogzIrd0KcOuDDv20wMsBchjuFZmLWq2dqQ9C
WKwO2UoKBle4Vf93/HB8AHCQPGmjou2m4C7BgAzStp1eceZJwFCMVWY1bWxqb8Sa
ARwAAI5upuhCGouk+TO5usc0sqZHrSVbZkKMczKRiy7Al50vSDcz5oEymMJ35JoV
mNK1zKOse8u4kjIo8UGC0g4Nxo+5xwfD0t3GDetCYqd0boHEO4jBBP7IqcAzhbZT
cFz0Jn0jjtmiZMqXFB7g6+Gj+I7YdXVmab86H/maHKrxkLvEsxWsRO5DEpIuEYRU
EgqHNLfMgrGbreQkBGrXcGuhdQ7OH+frB+U+56Iw2441qHhtLdPJEVLE21i8MHLX
5ecsg5huvT9izPYaBK2iO9i68ANies0Uu42PpZbMRYqkBnXxjzqlsKEqNUyWYB8B
F3QQ5l6KoXIpwDvlrVuzGaaVujl7Lbt3WJJwY8OZD/UllInLdU7U4n1gopnHQbxL
Uqt40Jc6tvRMJmKaTi3lkRa6RgS+4XeM0taQ753o0A01FCPAemNKTzfNT8KuOje8
L+t2laMnAKA4lenKkA/vWSupg5nnuqWeaK6mXwAMFKlYgseuK8uJLDynSiJNJzjz
t1hIrPuiqpsvDmYE976dX8eHkKUL333YI5x6JVMqAD0T+tKW+nt3B6YNzBUGfixk
S4gaMd6gtlL72MIVqeF8klgCaA/3NZ2zHxeqQL6ta9nnruqwpYQXI+rWpZdv6upB
ix5P2t4PM2CJNS+ToidH3UkZAE8mWhJfTOJ+0cQ7zMcXigZYFPxM4aXl3QnCExCm
iwaT+MoAkTG4kC7jSM2hrOLDxo463xlsqKCj9yo4TIvKPKgGCeTmbXPJzX8saleX
ffP34rEEw1wpQ9jCT5jHbhn229ijbcgLj/aa/pX9q3jaNT0MQnEKncwP/KDd/znK
TYvr712tmDgbtP7XERmdy7nfnIy0p7vF5sSX3WNyMTqLcdogjzUbX/zTkUrYReHT
B6RwkRewCPe3n7vyq+RW3hX8vnuS2inSpUsxDANxcG9RU+TTruXnIzCJjJtgYTOD
5/E1+1KK8zF7Yonm70TkBBNovQhRXU6iiCCz+0KAI54Mr3TSV13BuiJTIn4Ypfx7
RSYmIFXdkVHX8Gz3u6eaf5Rq10I4LsXy6w4Ewp9AlI3oX/sBsqaaS87WmQkdw6oe
j3fpw5LysxC++gR31AumO1Tn4UCszYcWIopBVKprNvLhD9avd4m76OQEF1+89uJB
PUrSpe72umhBdE4famCCu8AhCKrCGDiHJmHCKoO3jKGCFnbrdYSrQnIESXLy+TvS
rpsTXJlmLcSLxHKd+GVUvieMCLfy8TB3u00IGChiwvhiFk8iTbKUzxMmMpx9oC7M
8/ce5QdH5O7PygrWNWYlWjT59idjdKF2ZWyCY/C8PxateJASgflBaVesOuP/sUTZ
fa1Pyz/GY9Xf7loIqH0tfj9Gz4KKaEQRhLfz6Q5JpxpGt3u5aFFDDX7IhX+RDc0o
oJdRfMeAZaYTbAUTqlvJ0ZDu8EFJI60BwyCgDKluAcsdRXkgXBqI4z3l5sbUukve
F6oc5tYo3bbO+Fu6RdMt4JCpDElBkpSnx+E2i6yBtt/PjJ4iH/PrPow86Jzk76r1
9bq/f/ogQxQaX7J4Bym+K/b9VbNv6Frcan3M8pfgJ/eNqZia7T6/9ygWHexqECfq
EXvYygkqiLlXkilG57BU/lE7ZCYEUxk1InR3FhVbOCgjOrPRScn3n+PbZdgQPVcL
cfsuUJnaR80XadWXv88HO748WncIV231/Z1UyHFxoMLdUMEnu5yFMWNwsG55Hnd9
FikYqLLLVZ85z8iMesfmURvzJnM+ectAMugVAbYrttLuQM9aF5jRo9t8S4HexXPB
z+5Ndjifwbw3h5WO3TdsOJrXp7nJLuL0yFmTZ0Rtb2pZNv+2boHLUiHJVa5zqJqu
BCXApr1oNfLrgZR+jsiAsZC0JxW90Dph8DWBs1/N9oNbcD8XOm1vh/rPDmIQSIyD
YEX8+sOj9oThR6gvxgWpITx7tWoPiLlGIkAxxbI1jjvV90GD7bhAth7vWVKNHPzj
hIm/389n4wmreZHS3/CRzp5JQlOdNi/VrBoC8lREp3SJXE0HTr6i2f9mFSLZJi7u
idv0FW1POKaVOSSABxcDqiAGVPig4nQBX3fYOA1Fkcb7DPma0AAE8R/Ro56dMRKq
GyfjgTo1cAH9dEnO7moRX+BmNORp+oY5rTpGtkiUiWAKXfpGx/wZ6aEIGIXJdSO9
vWbObSoveTY0+fXNw2jwxvF9KXnBjdSRqyFEmYGQvcKHgwGKQpGZCgkoIyQYgxjO
+sIV/RxEO62hqf3zZz301XHHTXP2aUOHVCwVXWj5OQd8v148GkSFPxbIV6GvV1sV
gVzzY+fbWtvBCWMGMFo7Pb+2p3dDxZrVJ3gLJwh6Vtzg18Pd2iSqUI2d7hZIwkRO
st7H8qm7aznaIiPipKjWCGj+WPMSU04qfamoDdKAnu98QCkVyhYmLXQy9dSxe4JC
Vgz33jMPSRcw0PFnwsclbOjpwpM4XoZXmLIy4BTd7OAXcyiylFwiTYOoNMLhmUsp
CoAEYpJe+CkbYynCPl2befDslY+Q63PGqcvFQ41+1Aue2ke5/y2M7V9T77PgucyR
QeTHIYbDSNhUBaXCg83E4X3b7BlO9EXZSShq7iNQlC+uHCqpckCoRGi1t/IaTZ6V
/305O1aPM5vqSnfoQXIOQb/+Uo7UD/I6UpJCM1R7XVy4U6p00y0rzUwVA4Zy7SiO
VaEe+U6qfojBiOJgnveZkVg/1587uIqtd9ZQiwJd9MPs5TOYyqR/PVrV1Am6GedD
EeKdTSVOMTIalyI6zo5p3+MahjAxr3r3aS1L37HuHyFPUClNckJnjMlKjTddj1Mf
+TQd/ZFcrUKGHeEahDwpiqIUOujXyl+BroodsmGsfZutppK3Db7ROgG0Zcd1sOFo
KVUmylhsA/G4isG9EiGvumG7apZMpjwNOqQPucDpk2R0kiPd327OlCCJvn34e6z5
DlaaP7+GJukdi9UNxEbU45nWmcDO1Eatj26tjCggXwtMqt4IPgIjKAZuplDqI4qW
unjF3gpFH7CCU+ftSm1/PSr4d+VtrvKqceP6O4FoFuMaQVUW04ndaZW9lhHmCMCV
MiR5p4UqqBwW3r1P4nmqqwfABFzVLyOWGVzPhwAoXV7aPFXewpegFWEwifftK6/c
x9jC0+S0ipvjyt0+4X6LA3Dx5jTMu1rzm01sO5TvowuRGupsakEYI3DTUZ0jpZxM
QJVVXZ0E2iLiSOMacLypmN49FawiU6p9tusnpt/yYe+GEczeufmB7yW35rJb7cCu
UwWBBkaTGWGkV4TJUf0M2TlXkpQosKgCT36fX+FmfjduwKr85afK01y/Kz+zp27Z
ZqIUgCeApZjwoBP/GL2cCcXA9XGUSJ0N2AXn0rG3y5zoq2fFnRRaUO2hDjr+tL5+
2jT4BF60majT9MSNbCgkSDwMMN17wfeK+znbJWaVRiFtsTXwtemA0fbDqyhytdIX
fhujV+pY5efR1+UQoFENGMJwUHnVblafb0sfqKmP8zZZejTF2ng4gmlYHujYTr9g
8+UzI2vE9GYKpS2nv97sTAh+XBV0deMf8ZHvJCcUrD6uhzpc4UN5zUjQyVsu3zDc
ydLrHEUy2at8AiE1EMvYCI9XF9siEKU4CNhmgSFVm9SRZgOTCejvzeKh7GOlCZWo
q84J+kcziTU3zJUKz7pdgyO8RVhA33NhGWGFs4vz5QK7wKPA2V77Xl5hkj5RsStV
zgnORx8TQGZ1aLTjp9h22GRkbU/JYGI7FSVdNIug4oEnOveoY7r2kgHVuVEaduoV
Uo51FFKSUB4JzyTe8VJgLgGvn48RboWDVDqJWjk2lN5i3oat2NaQJ8rcbCZz9VB9
av8v3YMmHsqxZpXTJlDpt/42KYAfQeIhuwoknCvManhQscTx34oiwOmFbc7RGbHC
U5TAArxiWHzD/m+DR79q7ViE8VINGa99sgwf6bqYpn0JYcS7t+dp1b9qKMPiypzD
S0WUPoLMcj0fof9ZpqEUzu582RE+914xa81xs0FirqJYJWPUyCEzmxhIrrEFoG1T
YiugoIW9uI8n2ln1zAmnibsmQ5FfzZp9J3b6IXp7POtV4cjFHniftsVXa3eEvEP/
QLndMgHJ0Cgw32Hi3qp4KTSyskRWBlyQHYHotwDePoX6jKbqlcgCwMqFOcLDhkR/
ni2adi2rn3AEvqR5qR8zfDCxT/b+syzwv2tQXDoKDd7ZvF3xsZxt0IcmSy1yf3wr
xbZPNZCydLSLf3gBBmW2p1CB3iZDn7dGFd2xJXRPfzr9xR5cHehaXftmTWmnNHev
oFpPH0iepTIwjl/WVoWuCe6CfvUEmVJWCFtuhbZ4otTF6iiK65U5nIo0cULDAVlH
lNaAx/8cMjv70pQ/VmrTR1jhnIX3VcenPINRS3PfQ9izyAw855I+9Xe2TuyqhBnP
GK5xnPVf1RwPEpRxFV7hJvQhwgdtrnyfMcwtuUCXum1zSF67bHiUuarKE2ieDg4n
FVq5VYvtLbN4W3AqTIBmPqZjd2Isa4rQcECpOH52YHLC3Cjuhi6+/b2onqnC8sRa
YijjdwmqYXjug3AUvDb008NR6EFYnOCE0CA70vtCqO1ySQfXM9yJtBmfCNQi8NK+
hUel8MvMkvV0s1vj2dLj/fmae3sqDjKccDOAPsmAKrybRg70CUdyL4yTim0gDPlm
Dp3Zirw7Mj7kZ1Bd3ztjBhVj8t9MW8hCnKvG8tmpOaWmi1aFIr5Ranr/0fgviAw+
5HIzzORsdNgAA3jvicSCnMITnuLAP3+QvToc8RXXxCWh8oUc+pTboSyyRhNMioNn
cq400pX6HeBoglkUado4qnnK/C9pgtFnVSQSKUi7xj65mSM/YRuCIfHZlA6MuTgi
F/b3dKzAVY5o6CSFYx/QXfqVc/f5B1he3Yg7/tp5nxvxZQgK4Osi+gGtxLGdrCBK
O9hDjz720LS2fIl9SIk/4BS70gIV+DDc9r6F2wVPy3V9nkSbwDfm2mzGzTOVr+Ii
1RaP47lkF2MhkduvJieYHDD8WHQSMKVWHihorRXHFhma34fAO/skCEDyr0Bn+r1v
mdyUkPv75DM3C1oMBLZyftTz96CXTolEdqny79YEyX3Zhjh2Usy5FZFGsD+78MaG
0Blnybs1f+/DIw5KpePcx84e2FG4t77FyGLfbqigvPiwDti4YDoErI5X/l0/lXYp
oKOG9X2NmXRkzusLs9M2L2UHGAOJr/irCH4++siM/rLFIkeF7QoG/if44+DjTMk4
i6k+dPKw+wnFSlBGoOQKdXkX22c10N/0zWe0L9nxEjpTwSsfMhLekq9dCZcvYo+c
E11FLUdz9LSeFfrIv2zccUWTuIN+5O8RdZCjy2LAkrFPbhF72CHKhOEDIrQgmWiC
JL2OzdSe7tLA6XJ8ZrQyFvacV8CVZZpBv8rfeCU/2dZSvf0SzBqv51bamP1/D0gj
ltIFfurntz9yFv2dXM5UW9zuhRAwp7JDDVfnyi3dUAIg6MnbEvsm6OgGdyLF7uNU
6wt1HqOg+Vt49azhv83EIbgxDgUoIGX4mPDcXugWNeorwLeZxfAxXaJtNq/SW7dx
ytMMMJkHiecoQ5It9f0vJXive2NTO96SmMhL9NZ4CMUe5GgwnJbxe23S1uEN3i0j
otgI1OTURZrJqeD6BBIvcGKSx4mDwReYSqJ2/dPa/nKAKY9xYfhxLqrseBEaQRWJ
Hrahl4X9v6cnV1wA+pIwF7LnWehbxE0WgFPHwUSeVN4jLmnGWUZ1s2GgVmb2RSEa
Bij2w8mNT/5bcYJcnAyxxwc9zhhrSLKXDP9dGQ5j9CCCRP3Adyr4xzFk3Kz2pXMP
Msa8ed3ZWag+W96Xz8RVo2uKfK31zCXRuR5tRfUXe3q6s2EFxit/WG18OYjYkAHn
fSd0sb0g6jSZI01ngLi31j+F4Yd+fymqiHZ7nPRu8rcsNzT77VQs0RM4c66yPuiL
SCdyrOlirr7LTlI0dD5H2kLkF7vcqU+Y+djKTqr0zDw7+5H2xLYcHR8YoJnaQKRq
Vqwh/IsxXesFvzo7uiOmGxNuirMpsvrLU4TGn38tVxPvzVU/2YFXSZGl9Wj6d1w5
gmx3YWaE1ofs/v8ce6dW5vAzzlyeJzkqHZUm2qvFUwK1WMMWxSDyUzr4k+If6C7G
B1WJIi16fvI4B3jPNnnp4xaXcRbQaInQDZM+n4paYHFdxmLX5Zzy4RgmrbSR0/sp
5oyW1D1Nx2q+jPW1Tft76MpczhpFsEPkGQ84EwLjU8KNLlh12SJfplbUwAAPjd/E
29lzbg2AMU7W9xKLVsn8aogXcPXN1orzV1a43SMeiVvZ+W9YAN3syjXtld7DC5AL
Q7/SoXhkxyzWlRnqSx3Gxv7jyZcmjFbwbfXKVRVaNDH42p6bzi8kWcfLDqPRtDDS
CJ+uwRJn8oCbR43CzCnyFSPmE+hkdbi5ahz8FeTUrVa2oBs6Ru7wUSg5TWQ9gs2A
xOMK0QkPv+xra7X2QF8Z/sO1UNVmhd3+q2W+ZPJ7HmzXo7mEAXnOCehKbLlKSI/C
dxCOAexbqvLzgMCVK1Fx/TyYRPhxsBU0/NraRyEI39acAXcwb79YEuYwXiA8xZUY
alx1kMTdBLKGbk0+w6V58xOOnPyS5btlfCZp9c0i49PNOWjGBxLPmAi40q/nGbaD
o/r7d7WoHPx+EASqd5tXBycgBdr5/buPSOPhFlYe1+eFbMuDwKUjJX24p7VB8bMA
EA0wX5bEVHNzRcjVNOv9TEjzZ8A45DtgT/cTZKuIXB6xheJMzmIWw0JKENKRgevc
CRzGBaZzQOb5CbyCqxn39NVwOVGNkEMnaljb31n0hhKzv93qdEuIO1uyNtrKFqde
MdZ07jSIEL8yi8KSAXWZ7QWjfxi2PtV8Ammf/RrqaINGZIvVr+6FmaCpsMIQsQcL
pXZeKCOVDwljNOGpq8nCTtsIxy2XVKwOGCSUUidGnIyNPKQIuSG55UibSNpdy9Ah
sSm+SUtjYoA0UtSf7phmkxp0nf6GiuuQxqqbLtgbpt68rYdQiOzxT9Zwh7mSU4QN
bT0OfjC0PiBUTkg/WsG4vpSWlX5FAU6bQ2RItxHxAtidPOPx9/y6smumjKLUUFIl
nZQ0aLIuTjzZ3/qwdMiKvbc75uylBgIcsxDu1uJNkKwu3cY7yVWMJEqGeOZEKxy0
yCTk7Wqd90nioCZ9Frei1qwd3N8NQjVxDsFF43EdZwzdxdV+FrBlZY4hUCQaYHVp
8sG7pFr85oJNn2JwqIb90ES8wFI85VB7+yaAvxaDUYX2iHHcA2S356hWIWalN2/a
Zf4bA9kgElkZMuRutjwO8l6nNjUg6bQxsLylWPLGh1WeKgTVP8fR1zfkv5ftC1fW
93InwIADlVKBBdUuwDsLEVq7z5OGpn6Z5TJqnCqS46AAqY/UnKeP5azYXrV6g2x5
NUzXCHw/AMpcaAZRdl1xofUfazisW3CIbD8lzIuHvFXl1Z2c1QRtDmFh2STt99UY
OyxV14ZATIDplo2PEhG45Swb8ZGM4QcFrZ4HyxfDpLEm4tlXErYDu1jl62D8XGLn
i4hVdKRdgYo50h7C25gArIbx75+K4Frh64rSj/Lhxe5toc7fNLJ95iwGxOSx1YMG
ENaa+qb5Wm+/GcYEC/4si6Sd8DSAQrTeMpa6mI51CAdBnuhBYtsC0fkO70j5uDgG
PdkjQzRIspoT5Fy/NZvh7lRwT34/u0JmrVuClGIbHAGbJJTaX1q3TpoocGRMxcrv
v68eEZPsCLG3qWVF7/ovI7v40pXfi5180pSxb3zuxHSETfODWwndBWzRR0WSrE0V
jrCFlHOxCE1O9vY/hFMVpYbfGBmVfFQrfQjtXrtnekVPluSxNYpTND3Gns7i8nnY
Zmeh2Yk/4LgP3ob/ko45yiYqo72EsPv3/geNxBxBJJStO5ALitHb9FwHRoKmicNi
O2cAsBJYgJmerW0KcFUS72WBKJwvjDMXJEKxFbH6xooCEgXiZjqp/oIDPpWHWChW
eAGUlwTyZkPS/p3cDNIYA5kX69gkLPH998e3e6Yj7RGBAB7l9mO722n0S6BI24hb
4DIkI/9wJHKhwdZPqPFiRecfzHv+KFu/Wb0w1dItcMiOTTc32oYZUPgH5Aly1ySm
daqpWbSQNwZ0pPIFiR5mubBHjkwwkIPt1OrQdWT0IYnGBy3+u4CUHviexAy76whq
Khhzihrikzj4fwZlyMu7twrTQ/RLB5pmmE1nSDVmh4fp9nYTK7V7kuWambfByu7B
K5olBD88yDiUvKwLMuCUQLQnU/CQk0bwrMa6YIXbEwypdiuzF275fmGO/WSxh6ww
fJ6kllfhXTGUm/myZUREYAONiSB1ph5G9hk0GaPC9Dwp8U4t9cgtdvQ8ky4aPLUr
jauNtAlL+HCR6ZRWGiAPDSS/goP9RSdcyr+IgxUe6Q1JYvvphFOhTSVxod3fFRhY
mG8GI4j165X1793MbhDE1tSvwqO/xIwMDeskcRC0SZPdIHTXdiPWGDBaDkZjEWv1
nDZtHUb2BBtnJJA/xBlP2OfO+3DPYbdOKtb0PtsmQMe2ZXSb7XyBhDRfk0WfjkB7
pD+QLDDxe1zZT/+mWNdFwrZecwcGhBHNCh8n2cgMIGjEM+aWa/bbDMVjvGUdqDzn
VFc8HcrzSsq87y845tqGkYfbbigWU+JzWdI8ilZEHomOAbVC1fya8NmZvB4yfWvd
L4AfXvZ8esfH6GFQU3xa0woLGI9qCUfh0ytS7s/xAKZll73/JrxpFqQK1VgdFuRp
26JU4VuIbKkreGqcjdk2mw2iEQWVod5i59vMzj0TbUFLDjApFX2aMBD3WznIWuQP
SP6n9JRouEZMJ/koXFpaMDr67Dmr83xuJUU8es0dldn2Q7V2gn5AGg13PObp3Sn4
MJsRtKtlD3mkle4A7JYnugDblWzo6FanNQWEdaOwpSZLRR0XAEXxArkMp6F95kij
UMskjifAjTeV2ZN9tF98wu5jfT1mKCjl97cEVIgSidOCv//ek18CpLjJqTy3Bx54
AmpwEclazK4PJOaG0Sb1Wnaa64tLMIJkc9P/GXaaGMYnDUrWuVA2KudDe4n8WCBP
k4YymBAvJYCqXJrTVqdK5PytFAuysgGQm1LXSTIqpZ2jQebcjNZHXSms/emX/GjD
g8EE0pE3bNxsKaMfcwhBG23XpkkxVvOYqveWLGw0J+9VNqiY/Do69fncp2pXhyly
hktUxLIY48GjpEEEUdM+5Qf4n27d9blFOS0000eI76mS019vel2GI9sPWXQhOzXh
j8p6L6Xl65bORA30AC6dMK4vPZJuqNwzsTipH4Em5/AJxsZarw9QEJY44vysUvgO
eGWuk6RpS+tdpzTCsTUW0GGiJw3npGKiixGjtl9Q0tMZP66a8pPJ4GIyF9JmFhuJ
rn0ten4vSjPdXuhJaFusZ7sSyh/yEBrMIouqHaeAbkPEBvPax55AkH8jaZW6Pv76
/Bz5ZOafBbKayhpG8HxpV03aOcu9qtMXaoRz+KM52I2PeoI9BENyU6cwK3t7FMwc
GpzXBWet4WWye9DuQDR+y0mIkrR0VrAJFf2j3Au9QvBxvif+0M5a57q9IsP7M6Qb
8pl0w4cSHsvVNlhsnO3TP26aNn2r8O8eOH0M7HG8aTG15KmVTxAJA1r3Wwf7JcD7
R0RRrnZPK+VzrEFnEyfsK46h+teBnl2OtmJD49X9K4qtbg4mvP14OViG5Q43EOj6
JtQkr0MaIl1l3DqYEC/b71x15wKRD2iYieuxP6HCylcrbsSFVhonmChmSVq+n/iz
gPC78znd9y+JW1Sxbl548UrYP6pggb/FeVirWvM7oJ800fZ763Q1GDk2DhTy/LJZ
WAHXrOjxYADvLQI+Ts6aam8epCUlDfTuVqWaMmQZuzk70hnf83vGY6wsZFUrcbzw
eBRsifdyGp8+lewUTp7biMKthb0vEvMD5njn3TcLzrwxWoXwJKkYPG+zghHNvigS
geLXGgeNSjZiE1zxrP2zCBKEiXYoB+lJZx0e86UbVDbOyxwzy5fCmvuoehtJJfAt
ob6GE3VG0C19X0Rr7fEr8nhJqNmHvsMQe9BMKAhLVgGkdPaeAqpZM8YFBUiivtOx
gQF5+16b46dy5zuzwKKihAlOulS0B6NS9SP6a1GyyrarDsT+1HBP24FeXDYhQTzs
qP6nBFrnIx50/VNJ7btI1mqIYUZ7BSa2ruZxC5usBrq2pq3k8yDiMfDXLF+DG3d2
AKEy1rHTRdZ4BOv17n10zeM6bxatF4tTnrtC3XNwgahXVUjRfiMRLM2qM0zX4Q6f
+tu5YzcftaNY3Wi4w6bB9EUXayrlv/9rhrsbNn8r+SbLpoOugDiO/uV2YZb6XnH/
8OHguILMpWsazsCiyufOPZsKu5Jvoy7SXGl/8GWe7oSwPyL29grksgrFieGse6eP
1YGEhtdbFdOF+PtzI5zjtLBAK0YJOfA32KCgJ5W2vOPxLQLDCQvuzcpZ1rbw2BsC
Ky/qaBdSU9MFwyfVOA0LA5MiVAvAISScZJBXPpY668MRfns+pkQteA05PZYe6+7f
HtTw7NcGsS25uJ0713F0FfNwA9YmXtD70VujaPzNunE5thFvY1L7VIV/ykiYBLUg
Lkz+QPPb7UTzj6CDaXECPm/wG7+5WXAS6xW06cODj7sd109YMW1WdkFadr43WViM
WNEF9dYNpDLGMtDPSkncBB2u0Tl3jy2cHf/fP0YCPl+17t0zBDeQqevrNENE000y
y4jjXQvdkDEsRy6GFwVUB8/1DR1jX3GlKkJwOH9UhnyUz4iazkb49LJZagwWSBeP
l6NqTPCSKYO7RBZTHR7WHAh7lUfJk2I+Lyzzt9C5y6eHkSDgxDwjPc8epfP+GVXu
CjvPBUjD9M/d9tXYyukNhB5Gf3CtaiPWZ89b6xa2KKcbjS1CGs1Q1lXEAcsFlTrF
w+xkkiUlx8d099xZlJRQrDffAsitK8B/6OgQII77IWFSUNPRad23N4VBoBRC0Mxp
/eo8UUl6yx6zZbqZDnfZxvlm7N5GkKi0UaeyqZSRDzvFnLQ9jMaJoQI7qcGLC7w1
WhJz8K26KwXMjJL1nRBteX5yw3aQvlsIZbaik8cHBCCCRDXWxQkFOvj9Yc+nM/uU
00Z2Zq0npnWiswg5sIo0lNxjOj9fW1e1bctHS8VUc6fMepQBXQau4EB4oAQJNDvZ
QvJku50aIqHhe+9EODweV78Tw7e4PX5uW3KfGjZT04ujixW6PtcDgPZ/7BxG1RZO
Uy5nWgrjQBKO8gTI5iTgyHSf9iSOXvTuxY/ieYG4trr6M4A0TFm2u7K3E8E0YNVX
JA9q6IZ0zdSYi+M+9C1ya8eMuDOfdoE5FH6aGm+7wm9Zn49o/HBYFXpfGUjTuMRu
NThCeLGO62dez62b+u+ve51a1Q9/DU4mN5glmo2irU21Uhnsi3pVLyBr1hIHogra
dIJjaukExGHToKt+kjEmPqju41Q0bz2Eti4bHpmHd6Phv2v11/vFSwapptmtMv2+
yyMYvJwB9fX/FhrPtBPmFne/CcpgjU2mg2/XO8N+ET6Io/hmPvJ1p6rz5ytvJZE5
TBhR7M5ofFWGsjy5vWqaYz80jePKutbmk9pLh6voO9e/OToW6/ZIdyMT4ZVmd47c
IVc4WiJgPOlKo4LEoEHdwW0UljIK9KvXrb2CPy/R9sQGqRfz3eOczdwNxLfpiK2O
Qi1ffRxmYTbm/RMk2nPn1+cZbPJLWzHlgEsZR7ZFOvfsVvE7uf4t4VYia6vYUMho
32kIIsbINsTgZIgcgxn++MqAcxGaQ0om1WI1GKsbI8Mim127oCycDwsU1IoxdVJp
qfrFyYUZfoY/NhLzwwTxTrtADcDS1UtqyegLevyNHjiqJkQzpdmXFXUAQY3D69bV
a1ksw1MiHCGstxVlh98k6lkljavQd05sTrQ6pBXLclJuMWzJypzHJSv5ZBDAk09B
XmILKtchJHBA0GQFCL0H+LpHTFjDSsa9/WqOroYv1FTXpTQmBmLc2K4ZkZDItaQe
IVuuC5FIpywsi1N05NTKyuLky/g4kItd4KLmIPA50HPCAsVfZB0LYOtd2L395snu
DVzdEvvlFGgmwcsp7vKrmvZ3gmBCKtu+mk7NH+7+U0mFh/QPMtvQOcz84rbZoJ5j
Fr7qr1Y7wJesjnX6/lXzAplwlMDSaqJQAddI6wmzb3qxKLzzkxaUt5qhBsoSzif8
ZPz8jNl7h11OO1iDHOit+0NXRvhlSxDP/u/l53VDvZa+Yue6Un57WWam5JJY2vU5
4WBMlqMQwmiZ72PO0en+dRcmV0nbEkwB0o484va9rjRQ6IuSqzxlnRxPfhqGIhov
/Rd/jrW3roFuhPkJ7f5PaUOmfWxojIpGsoJVIjWzwV791q5MeQdcLTuz9eF7R1xf
zWV9zbRaV/hpnyge2PD+mme6hW3tUVYO5vWjY7Gi+Pq+lI73ixiGcJwWKSvHP3c5
3nWhxvnt8fD6kiYxp0sLH5xpW73gXlsM0n9tvEQyJv5BuLVqM6Fxy0Ases8F3O7r
dbr1odDn/zKrRgiVgAyox8DtO5fWYkdgYuZO87CK1gjm8J6p+LXmvS5o1+6TBYnp
G+w7vnsr/Paubopce3IN5YkiUZa0PnBS3cFPJHcTFHVikA1pSZ4U38K43csNyEX+
KLLgZXWIXruaaqdX7zht9r2BnwwrlQcsJ5iCp30OsQg9RrMja7CaZ7CQwatl8NG6
8MxAX/0/sKtbAp7B8twcyzB+TSpxuCXTJ5RgVLyCZMJAq4AnA2DXv9Op0O2zChHG
MRMdGsOTw4aV/IvmlKFDTGX2lP23sOEDknzC0lRI4Tcw/7axiG8b6fYp7vdsEPG4
4ViA08GaQ8S+eE2YKK1XO/gKdnb21is6vZQQtT9twrfgQDo+AJNVb2gcJiAdPgBe
fM3Vh9DNwE4tTlWBRQittTyWymWFsUffnSpHu1ibNJ1lpyjHLouS73Hk7mbXCy49
q17kUnmOgZORSJGh3AlHcEGu1FkIINIiim/SXVt5yx4wOxCPrpDOI1QLS1T8hLN9
a8JmZfmk8JVfL19EOCSVXHz288/x9dROGTsBWRRsSztuiVWoYaqLMjwrcoDSO/ck
NCd7X8WhAlub5ZB9OzuObv+C7r6XtBJ+snKoq1iHmm+CSBTa8R57vO3TSMq6PKsK
dug7wq9C3QX316fx3gGq2l3Qse8xAxKj/gOmW8bMb2ok4uGlcphp93U34ALtbmIO
KVfbGuO/e2ZAtzovZfZY/nuhJ1Ij183eHorwlQ1dn0ysu6vrTb4mImOIDmF3EFK2
dDgLEnG6Y8ww180s4DZI/Gj3r10VipjpWB4/FhZBq9muFvJ77q6LmGY7nOAH+8i1
2KczaMPD4BtdNXAiP/9PE/7heawZ7ZoQi1PfpAxDtR7hUD+vrN+WlKYIt4ryMvP+
tB0T5wh65SXYL7Vu2rXuJv5X/Iwb9Z4qELR5F6Hz+msDCfHN9dissLqq0W3RWovL
AFosKy6RoQncuJgyNha/UDG1n5yHKiSg0FyBbMFTAJqFJpTyWl3Hr9lqGfm+PAUy
/czkfN5itsmcDBfQQkmJDY2onHrH2gsTUlz7wc27PN+jNL1HTWD5CdvFq6Yxaeu4
Z419slUqvxFzQ70lj5pot+8Kw8XaRI8BJR38eFCc29NNmqW4ffNGIMqbne2a/VaK
vQC5tJdSlL6xRqbRsi75O7UYJJWPv9ZoEvQXa3TZY6DCsd+Xjhayw7hg14trZz6W
rdkVtlA/fVQqVHY6/IZPjzWtG7RHiEGDiiE0EqIpHJe6jl7ZGQGGSs3JS8/J501W
wuYNixhwrR473WloS7LAcEXoWuvlex7yc333SEk9CEi3M036AQPb5GOv6toMdXF+
ZRd/Jghb3XsEVRTv9feeaKUxnx+PxlFb3LrnCx3Kb4rO0t5Iejyu8AKxSOg2dmLQ
nyM6HLd0TTcnBLbJIScV+gHLXnofbd2ZKuDF3rtRye6QgENFkYplKUNiM3JeSSad
VjxZlqw1VKO9AcnI7S0PL51hZUUa/CDtPEKoH+NS9ZkCeHbzeEmCeUnUON968eSf
P+M8L7ailOnDNO+Imq0Hxt+aWXeM96rfR3rqsoupZK+ily49uNfaqGXowUCsUdKW
eVJ03JLTbnt/u45Y09JvQ9jT3hs4aDMcdho7aqJEC4qqS0hTl4V/srh0DK4dcU7s
x3718xf7tNqE0Ptclun+RY3Gw3E04cViN3CtyxQtXqUUDFILp+lDimYPDoGDigUi
R/6s88lg6Zp6Osk/LkCnou+TtuWHy6OhIN6PbM7OE/dwD3lgWm8h1IFskS0digE1
E1bbsBcR9jsJUvlZkg8Ld7FG556OrOSfHqlnAdOmPFRFnT1Ah8NCR8Hy44IP4d0T
KbzYs6FD1iXkj2KEvFVUWpkS1htWqZcU0vieNHxVc9pFktNjpHc9cQfT/7xEOXRo
tIjum6K1zGvk8lPRp6xAC92o5JCogguNp4uNoXFOrn47caJkhPiFxzIWis8EHsMM
ZXyggbXk8PkbwJKxkddaInePrObUOJQD0czxBSCcY3N737rLBcf/K4MydViFMaLv
oTmggkD8C5FyduwtGPpd7emgeQN/Cs8Uu2Tj7cj3SnFgzo72lNHBVczMv5uMQaUR
AELcAuAMHsQ7jY0vOSnhXnpFOfUBJ3xNekX5VEl1B/z0S/fCaXJhFV/Alxe1zg7p
jbf+MWbtDoP2iVzOpodRSBotTNTTmf93G+27l7/KloH5EIigmzewaa3XJd9nsYKo
V1Gbm79wYrlOEg64+kzQKqV7vaMcIMUEJXXPK2j3YjpUjmLEeTtMk2R6TawhHIfS
EE+GF5Ge98eqVud7vNLDsQtCh0DwLP0RPX3SbTE7tN/py8OmCB47B/jCZ+vjq7/R
VU5jz3sO5rYqJplH74LNgYzsC3E/VZWZesH0hGDx522X4djrFY2TXJzdzeFY03P+
qXMW5AQxTq6Y7rlynwlitYzv6hQRPhhCO1fm4HmVNYThaXP6m6E3AuHDXrSyP0cV
TA8Rwc2QqxTupihzoCup0bfFmMtDtTF55t0a+MIMdviom+l1ayv0wJ3Z0DeU0cao
7UdIgpsdr/wstoGoSHOAmBAJizUVoALl9fy0N3ncJSo9LdYqvbWk2NS2+tVlySQ3
K4Ftq8gr1UZR6cBVHYDIg0Nmzh7ugNZuGLIr3BR26hmCHj0imNlWlhNI02nwJooy
zsUh84hrC323fbqeOauO1SdoLNbOUQpzK6HYzji16c3VMyTBmGiuS+a+eKIKO3XR
smRou8yRtWKEbsnfVXLEMTAwrm0Ui2dysuaoq7Xz0K4rovHtVJlXBqpUmqVenxU6
Kvf1sHEriTUn0QuamyoJqAzJnINCTCdCKz0LN45AAeK5QRd8aaipwP8dspf78XDN
QnkfStqWU1Y2wWUuJmucLiYmA+LGA+GR+4Kmlwptmy0JFpJK7izBcOPk0CLPSO41
UgU9xteDg6yZtPiNtLHfEb4yYIR1qRos3DlawF3uWgK/RDEJF1TtKsjfWtw+rkXp
GVGwD1l9A3av/Wa1Cs/O58yje6m4oS+sDEWOVtxHwXft0DUCbn6Y/O5/t2ygnbCp
HFAz2DCoqQh6srBrtxyOiSIEbVfXuUZFsw5oxLe1ZW6NwF/9gZrBTuao0IMt9tD2
TRctGuX9WFdmRIEWHW3ZWAP83sunsKWjhKaTvWuqsNBNwZD2IZ7Qv6Sy9ipQA9Hc
SYA+Y/LZxckLD3duGtBqQXOnrwvkYLydE8c6KdUzAHHGZIqsBR3Q42LrQpI94RlN
ehguoAjhmFhkaBtnCY7QvDllKOaRH2T0DxI7o7de+Eg9sPGcK85WSPfmeMw4iszF
dzHrH2q87CEnIGtQJvy26FVkt3+7amg459JwHRfGqZUmF5ERUtrMf0eyzb8i4820
LebK/AihPnEw+mm+ZhIdnmz66YeK1VGlrTClsyr6epGRSmxDBGJS7p0MsgJt/XSq
ZVlpCKmVzHIkmrFHUHYJ26Ws1d4jemoZTTuYIrdHItD9d6HW3yWzexN2dmKv8xC4
S+dOBNC0/QJWeZNL2laZzqGkjf6Quhd2/RY1PMrOFlDZ7WGatihPx2Ji7tXTcY9K
W6mejGzEDsEhM/MwN8YsWQzYBXKAP6vFpDF+qI9VI8WP0hijrG6KJwKP9fbNi9fQ
L94t2d7X/ilcKN7e6pFMmWspxA8q+3bEJfrF3cK74lB0hCmqo+diTCZ9N/8LosQG
bc/3qNtCJbhJRjBoD43OL9TuxmXXxkoK3BXjpYBbiOWsqcWz6djb+4mI8glO6l2F
sZGVuP4hdRdIm2SvmlCZCr7NRReYPHF9UYNT2dYLA9ckBqHj2BWSmvo6z2uJ4mnt
1yrLGeY0cX0BVPQA4j3qnrxUKPU2iqH+tvBMXcXs8ZrdfGQjdKofmWHOlx+/nqu+
4DQelrPbTqwoequPNDXSZkRcZ0h8Xp9sPCyROxi5mByJDczLuEGSWu8nzoPBLbHG
KDuLMAdpZ11w/Y1o1KIqN2b7Cpt/Iha6aV1DIiZrtkroNOQl+cQhXHuWzeht6MCN
tNBFLgo5YC1r6l+KaPhzQi4HBA3x362uTiB0VPC19aGc/5jWNhnoKbZ3LF82LINf
1Rm6fROhQ3bfSXXpMhfUf49OVZOVlXFvsK8WMuiaN5Xo4r1Lqd5R8C8oeaz8Ku+M
BVvf1+rb2U78F929xQYSwP4Cv8dteC0PwiNcqup0G9e22NPA5WBS9BzJSulurLiK
ZhiQI5d+2TGWwh9rpUMhYp5OScnBjBN262bpzJlPBaj+SqIt61pldeabU3qO1yts
/IFjpkG7tArzGj7xwH/fcfkBWF5hbUHAdOCUa7DsuhTXS9fMEvffT7HMP+lCOPS+
oIhzqtLR3GeztJoJc5GlPit+eKH92qtgOPAFVbO11ocK1dZDWY3w3BOmld6Vuqj9
m6DQrl2hZ1GK4y8yiYo6jyiBBOBrWM3PnMa47uyKfi16PsEJhYr72V+McDau5dZU
WQ1KU8JTk5drZZJEBnYeWQAI2Sq9Es3nGFtY7KDqZrlYR2LdTdroQHWYL+7m6elR
bJNUdL7P+21AD5JSTtmpM8fEs3FP3ksacyzT4JBaa/a0CiQlHvYvcZI92nCu4aZU
S6EQriuv4+7zSccF3yEi+CYVznnBT2Irj5W00bW8PJxP89gCC0Z1/Hf+ZNdMI5SD
+c7TVqKBg/wBCa7U1cB9Cdn8qnSSaadHHUcUJbm0HWQziYr0fCJzY4gP6zo+P09J
ARWpZu5T+XVZLSbm5B16mLAbrPFQvpnbXARs2FK6hDPJe/YXjujtzVlII1SkUERB
by+r/baUUqoD9KkI+RXx9eePuSl2CGm3i0U6pr5c4+V8/BktKhJ3ZcowQaX2q8mK
PI7PtxnacLvuKcXtOXBTzIJcIxXFdn4GzucBEV6Ft80tkJZrKp8gHq5TIOj9bRY9
KayVMA9v+Vkgv0Aofe3WCY+39JDCN/ph0cORwnmBmSVn3d4oF+RtYmvw7tSu1BO+
Oq94tU33pUApVq3PUyXY/N+0DaoPbVVl/l7l+ioxTUZl1eP04/MlLCfYp+V5HO3n
pwlV0LKgjkWVmsQmBhJoMJ7oOOkoo+419rydIrBXcbYDqxy6OgfsbwOV7UGfpTbp
xaj71p6u3BXXjAWx+pL3oIz+P3xrm8IjiPAqOSLM82yDKVQtYWuuLWdCCuSWIJmc
DOzR/MUGFsdXo5/ZEcByIKCNGsFottEZKPANCBr34xdKgZHkXu8zBcGrFP7B4WrE
JEmHGgvllGOOdLPQUmTTCxdvMKHzLOTvizcTBTeNqtrFFuGCr7OD+P/cJEjoOlQw
FgK7bHt5/7s1Ab7Fbf8Ro3mXbONm9V8/x2RmExJbepdd/7q73LbgXG/2/cyzcy2m
TDPaAFAxSoRDNxTbKA50qgcXneEgifVildy3iHcRvL08+4swSd38Md/+W0cewav9
E1FDOUV5RDrUwbKCvqlALC9DkY1iTzgiGHvoBllt6pE2ZtZjpCs1WzoJyAMxxda5
+BQadE7P3ip8fJespcHmNsN2XpP2xgFGURJGQIBzqr2Zau71iwS7jCYpVyDsxCRn
MYOI25VqGlGFJQS2Ixv9iEH0wQ30i1vw255jOtyLcDq4iyXsd4hVJsldC9hfkjUZ
HkARvABCMgQ3fo//jhDp+Mzj6puCNXdDQ5YH1C8xP7Dx9lBbwJ7yENeTFD9thUdz
NTrZAFOIy+n2/4HHEdBe1gzETjdasjuf8p9OPNvYt5ut9Zrr74VWEej2pBmUANV5
AvgBgk+IdFiqueIsuld4SiGKG3Gnu9F+UmUnREJ7faLgWJEzVTg9fvDe67HZZt2p
pa7+zbhRRS7eRqI7ngYtgtXldTTLdL10SkntD+29R6EVT3U68wyC0EdCY1tAs9bx
3q6qvd55M5epLI3HeAOm+YDdC7vujrYBdspwXMD85ddKo5NbpueLeY9YICYGVC3V
aM2Ynr30BiyKCovHo4VaXW285/95QgqoPA10wE1xeSIe0I1/sCQ+OtBLMRCq6CmS
WnjVWYqMYxFQZU+UFe8gFfRseX4e72KeJR7urcQNmMm+6HP1gb/E2d3UTZu8qPq0
b8S2hPix5055Kojb+DQK4/0I9p/XgAyK+NFFPyKR/9GT7H1Q7NB0lFhusJ1nuXUI
2YEEtALttcRFUOUYSSMHrA7eXJIGmMEULhLSTgoTRcLOtoKuGGup/aTnUViNGVhA
/bM6U6kLtr2XSl96TlxpzWvDS4sLbCPLTitYWZeBuNC5p7XqANtRipPmcMg1NJ9U
tyW3FpQWAd4c7274lX8xYyQSHtP25dTXjqWp0QH6y/7aSPuJXoETqvUFhXC1HS+a
k5inQ+3CFXYLYYkjumM4vMAFeNzJOB0ywNcxQUq39MvtPgks0mDL6r/G5LKlRvOZ
GDjBINlPrXj7O182ZAW+2X7LCe9Y/FBtyGZoEAtZW2fYbhL61hIorAX8cOLlug1+
F3XDONaPs1wzXkDFVLgRlIV1qAVTbK1YPanI5AXwc5oOQhGSej7Z7LSoZFcyLybw
m6ju3lsgJfUditRKD1C8Obgdgks07XZdOp0LmAdP3gGOqFw/FUfxLVVQfox6gObF
5QnjoYqU0gitVg9A8mT67NlMye1QVVYQfsYt5dphi0nywpweTh81K+46iwxnzo0d
rtqzeUy4wAGvhAlmUwoYlPUw7LtzruJGcJ6vH/BtD1LanVfQN+5REsz+QkzLd30G
LUQBfSJ133G1PkzkTyWRLBZbkncWQqxtmK/vohWj7dEvdImzyYDtAVT+3r8UEgIP
71qoMPfG45nW5S5fwdpGNM/k6yR90VHtaMCTRnKDc9/G0CwcVSj/6IYHxQprBJjs
MyhEnlR3mb8vFmobgvE6QP0qkARS9kLW/bw40OVmyo2Z/1JAqTU2wlGjYh6GHNVD
yg97id1D1mvHxet/uEFwy6dwg9qmrgSvaI7Pt9MZSk6GFqkUD08l5LF1CaLRBimE
nUTdBs/R6aqNzmrONifmtd9v5EJecVkK/fTxBxGR3dkoZi83dSzYj9+rL0z6hoVZ
lwRR7sXolpSsrFPj1Gs2pJ1kF4i6+C81yDPDcyecy41ZrjCawkmwCIgmXvsPwr/Q
wKVBBwqGtPvf2JOmSB1roj4NPV0mymPOcR4stYc1cAG5ZJ1sjwLFgLZA1kTHHnsm
dA3WkiKhVm55SAZjprnmX5qPd1Ezq+HTVytoEQHJCPqLKX5gCNFpho35S2UByTHK
PBBVWkbCajhrnkikd6+D9bK4EBanVu6fbSHenVmPS+PJy0VIHXD7dl89PSWe62Vg
7+M3BiY2yve4n0UPsvQBBifPrDHh4SL20SwCdB/mcNo5Bi+X7HDsuQZnyIsHiNri
iXfr70oWmaKDG7lGX7orGaqXgDmHK90+lkDry67mwKKH4SifxHKsrY3zx4bntflk
+T1SOEwciGG/1jQpy35T6uNptQcm2bmHuPzd961TxpdK/NhEyUFY+nVYEZHx904x
14+mvafrEXNyvhBVn4kdhsfZAf+iV6uEDl9rxzrAlGbO4wwpARjdKgvruUin4xP8
+xtU+W2iYuFf2uGUWgX2SZ0N+QdeCpYqiKMtqyJ36idcnGvfbarE0lW7LlePfVwB
yPDzUNr2hE76jCtMulVBTd8BYOK7/veluxUSeyzivikFXlwInWcxVC6HjBbHwAJd
ho/pYxKP2f22mljHJO/nmPbyT/oMrOuLzBaSIhDC9uIQLmP1+GaC4IfS9c6NsbFE
EgCiEVDSCaf6oYYTssosw+urNonQ+nv7QfgJ0y+t/YN6MnkeYzg2c28xu3clVeED
tS6HiH7jj5WyKPwtNQQwiY+P0/c9zj09KxNXD/6fFCyatPH7DlY4XHOEjQErbnQF
9k/WrGFT9/MzIiNuy7zBfK0O2L19BuLNuiEMvkFslFLcSzfg8xRbeSgoVLLpgl2B
dxdEtiaICBr+YRzQF4UXJg49GCPhAbmi3OFhYAZRZe6wFUo3lJ0MzKoVODCGDd8h
z3fAPOZyjKBKTI6XDkDP24zZ2FySIpkK/q239VfXLzdOkr7eK6gOPHqyIFfsNKxx
mRV0aRhiYJqDVKJDITiyyUmfw3GYQHGJ0qh+56FLEj5IoUK2FTMOKVk9P8QgPHRL
YPWHr0mJbORm9UWgOHZ25lce4zOtHabpzutNYbBKEAfrQNG5ubZ83+OW9GAYVDXp
NpMFVql5oRLKcRUEcnY1MJ7Ol6xDEjQai/NIbaGqsBEX9Ah9eU+9CQEkUrCGUmwi
T7ljN+LDyWIWzleSfuEhPMywrj+77voLv2Ka++GTthirVTc7V7bzvaMlwrkIkWxB
i7KWlDyFWH+kOgxEKQa/yZMdvEXkChHnyo4ZLp6A/Fdup2p1oowVkduKBpeapr+v
uaKEYAKzZ9rezsiAdFp/TejTlQkOpr6WfFq2SyszldlvjGFKa2Q57UXZRzB1hQEx
DQCo5iBlUlt42NEXF0YOIllyxdkmFhFG30LQ1S1DzVUFNHtdeQOccXR6q6IYQJ6M
jVWa1dpoTjAhid58YivXBDQncsj+IwbPbSgLtHevDH8YyJm0E1KC3z2kVnjDcYug
xrnZpW1oh7uc+7x4ppn6Bkh/+msewweU1cFdFAAETa0xDx5yzwYR8cNYGPggNtEZ
`protect end_protected