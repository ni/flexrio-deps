`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 57664 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
dePWI3aWMLl2Yxf6Kb+wcIf6+BsOzvOLZ94pOUAv6zxL4KHZJ+AskT/tzRbtduoB
krQNiNEx/GY8Uo3obBq2Xy79sH8fy2R0ikjldwRclhh+hCpBMtfVW4uRXI8U8c13
isUvxYlmS8BbFGZG2KQXugFFa0eqFkKeY61i3D4OfjmRcRwRJcn1PcP8DrwRcQ1e
J97yJdMKRjSAMhgNN8x68NgDKtAuS1TM+/zgfVUp4dG+U/D4jl5yfBL7jNKytxjl
/t9dbxL4yCoeFpVGZ7Jeds51y3Gd3GDRFXLi9wSVI9HN2pYZrRPdF+f8b8oFSjaO
QejrYaulKvTQxN48z4ObXxlX/g4wAmvaZgSgoev5KJR1IkncxS7OFYpDKoYHo67l
4OSjwMhsCO19FBQ6FUMpOj21fwPcE2CSHK3YYF1XuoSXW+95PSwZKIG3i1K1JukB
MfWosW4Cj/SaXMtGSY+o+RWOQsMzBmaR6RAMrRMcF/myGf6UN7o5C2LnhCAFbZdg
I0oP2SLuLm0g244MVSF0eTeanKLpZNkUjpyrPnAmi8GoyG/QMbCRsD9ZxevHYwiT
emhQ6vecRcTTkgJ68j3oXR8jXdi3MAQHYhJI+7Hh2XJjZ2V2AAjWTCFwLijA7i8f
fKYUCtkWZkCztPSiSuRutn8HWRpbhNd3wj7ylgPNoyho+zdGqu/STlP1IbvW0nBF
sGgE2k3j3N8O332lzLuSO3x0puWt6l+jDwvmsJrfF8Ma/0uqlvQrJSDr82MSxlRD
tV7Dud2ByOphVUFyrcB3XCwFOHMAJIrndiXXbhXL9tFksUqffw41SrTBMI+7CEME
TDckbDDIemb9TvGpYvChACnowRBexP+dTHpO9x1mpY65jQ3AEXMxef8ztn2GFsIo
Er2ESSpLSiEDS8zR/9maYtB3sFoEkqvTVin39HWKS1yoHRvGY4KRXyATlUbfLxKx
kBihB/FWCkJbGk800ih6j7plY/7T7msH37jvw/O6ZjQFlnnVQ8cNCteOYYAWrPCX
uWhadyDPPLPJ+SXJRFBSL+40U3Byg30pf5cg29p+wfTGDogduVApUGoN4kxsrCN3
2IlwzTxQAEXZH9q5yqolYCeysqJkg2I7W6shJQpYRVjjjeeUL0exQYTJ/EBosla2
F1Owb7epzz/G/tFCFButt8zoKpzNRW/NBjy2BuQRYYaaeO8UlF6AVDLQquHKz/jg
OSxL87PhUBqhJa4mkMHOMCU8wxEfjDWoNRGpCWHh2zDxGXXUYDPI+VciydZVNEi0
uti1mHGf7jUp0c5TIw0nJ8vh3s+m8xVyeXIQie+JNYe9MKwvyEYuhiXjPrO3Ti98
Bgb7paiNw/dHtHsF5qGil2KPI2UNUqCpv+onM+P9IrFEaZZLjKr0TIxIM2oJQthS
DWmyVRrWF2/Lpgln45iX/eUWsWPfAlL/xCeCV/WRbZW7/R9QK41h9UUanJlJFSUi
89cSROnJ3FAfNV/jNJYvMZ9Cnj5ulg/Xwy3Z4w53kehA4cHu75MCzUGmLLJoWBGn
cUY0T/jIFeBnsnhhdOZq8OXCFTdkFVpgcDxoBCsg8ByEdDqzs9vCRIscnElKquej
MkfFbE0neOY0knWzB12z7y/H8my+eNNeSpcZX/uudiOgtMvHJb3W1KVYCKnjmOnT
uD7aQ/0J34NPdYE43RgfAWoYWUnouyyNvJG6wd0UHsM6OO1k3gKiuvakxb1iYFSn
TEAxC1Vae7vt1Dtt9GxRH+VEJ32+BLTTplx8t1wiCGaohYG5KBCVy/zmIpVDKWwE
CqZnrPAhMYErhC/3KgRdEplwbbeJAo5+amPUmaferUN0Ge3TcPTPYJSXZzdXSQlC
rTph3t6aVFpNVkVllqgotNRbvs9OpOZufeyQXwcUGqPIKKPTrcBiDqbt2cWVo2VS
tjmYj91PqjpTqUX+FGOw81bav3N69T3VqKUXxBPX8jVWifBr3u1eSWyF6ANQHN85
sqSh6pzIx/dc34KYFu4REgY/hnccF+3wmiKLFsZlfr2XVMRYAUWfarL3l1gUb8dV
STjjuML4fGML/+qbFFHXxmio1ENL69qm/gtu2/l5Y3IrwOWNzRm5xml0PpGrnGl+
VmpbjKlzmydfSay3nZvtIWHdYCijd4HkoumTo370WO0RBCsMKocCVd9bqrVIjBBR
Zmgp+xG/3YUI3yzMRXLNC/djlsTxYB4/PgYkV+ZQ8jxpACtxkvsXfpM06iXZofNs
NidERrxlWpaeb6j+W6J0GM1JTPRqLuVw1RkjV2epPoo5yALh3O7iqSvv1jd5eeBo
ZomdekXRGGhrKC0G0g8iLU5JGySyApY6uruWZtIvAIZmlRnqrf+faQPnYfotA1mA
cficwo1js5aE7KwF827vjipyeLxBdj0zsq2EWmGOla7BpapWPtvREwfLKRkmvCRO
qqIoGmP7O5mc9XVn+/zG/lvdjJtbbZNdwi9pKos2T46lYI2TBU/JP3F1hjWrLYyU
eSuW6Y2iuKstVuQovGiTavxGLfS8+RSr4WlD2TeZYD17P9jpzNFzTlMtOxFX17Zc
gWQllq/kF8EApIkK+9ZWDLtTYUlKrxUY3Q2sFOm40epJcLHrjlFRpAITq7Ku0CPr
zNF9v8RJ6aFSGLwJbFD/tyE9FuAQQNhfSEmUwc00TAneDxMoev8qpPNEKWgQjI9b
YATze2SNsai/VHClGXwzbqiAGC08eDhRAt06r+EZaB3ABN5IJcRMgUG9pEhLFK8a
Ltqn5ovvLX+AGkKsLMmAkWgP7bOGs+Dr42t0KX+psTic8FLoRC/6fr9ohzz0WILB
qkVlF7VHwU+R2l2KoDdHo0t/VxaBw+Zaq8URYiC5Rxvk32AB8PJXwtHTZ0PSHhEU
dalG0pzKCqDLazo7Yen+t8Kr91az9mNn+Bvt3QFlFSnKxcXIzf2bJZ6UiZTUOamY
Cw8/kYyeH08fJSUoxpHdC7dDI3CBOKpCqqvIYL3Ru2KTv1c+nXk2xlb6mS8wQpRH
XNUukm3HbleHrsjcLPBNVpJ9M+ijrMUape7SiPshL2kie1AGsC/QE6imPIGPEAJY
146iviNcLcN9vFMD1qACDQXqnc1svQd8ahtiOa/oOD6zNIsdfA/kpo50M5ho1XFG
OG3rYXFZ22+1R+v1VZZOcLE0F/ZG7RLL5/q/YAiZcwATVZvLtlf1japp6yGzBTSw
1tOEKADbd0VOFJbyWKfbajUGVg4EF1jvpg4YfUJXdw/oAb/z4/dlLyXUhuDTDdzJ
ws7gQLVXDVuQcbm2gF+2RrsLAMrMTRN+RHX2RHS8+kpX3nbxbsNPD1MvUkvzEVHz
xN+5KqLUBOWGmmkYEGhGQDbZVG8w4Fcp3gUwuTBKDCbRbB435tgldLnKuZ2YPF2f
DLzH6BmWj+SvZySTA4Qo1+bxPq2e5uZ/Z/exBlIBxYPVQ2hOLC/yha06amgFAhoD
S0C7NhRJLWUvhQrXmHsqpCeV20gUdx9GeEKYGllKHq19tnXMJeCpVn9GyLDPNwh3
afrw3M+9MwEEg9BOppYQ6bmcZahlOYiz5o6F8o9X8FBlk9eJwVpn41m2/Z2aiPoJ
4xxnAzqOfyhkQUVH/DODIS7OCflGokFTgUjji00p86770dCHU6VK6DK7wyRaH0G1
MKnxjtMtxUb2x/aOrnn01uA2SwI4wAj75EMsMxHiiFwCfpoj4I+NhEuGvGl8CZDk
CaX3yJpk3AL1XM2GSprCkRb57iJ9xK8tVDiQTimk//XEy3f2JjiPiUGCgPkt0pMz
YS9s6+5iRLwrW2SwJ7QsykccAKDS+GCP1hHAHO40cAetszAjCedGd6EZNV96BQJK
7v7H3zDuHPyH0awC55qOmu0fmo0zCg+ziwIl5xKBnGdWxVcKcu8mOCKJiKwiA7WM
O7vZFXPs9gyf28FIeRMtkLT8MgRZ7qL7K3+jrBTvk9tn9oY0E7Uzhxg2I4Lmw+dS
74ySOzD2wean207MMSciq/OYTJ16pqV6rqvMySL3SartchudVzFSCIogw5pSxjwR
P7N4tc2TFFxcDLkSk7PJyZomhb3pbWGpIo8Pd/mligogNsD1wgnlkvgBkHqRSO4M
n6T1FniiBLgoVQTqPnrd7Fet1Pzr+mTwYi9C3fR72/+t8vBFPYpSQsaL3333TK4s
fX9QIKr5XLkII7vnG/3iS9zl4hftshnSqTj6bCfpyhiC0L1la+cZBHJfUGxfDiFa
d77ZCLj5bBzAslziLdE5I4b13IQWjLpXRvamhETF73JYEWMAnvTCpHuVLdUXZVv9
K08EUA28mmlWvpBbLqngw4uifyqwnlA1tXLY5eIV1JUAp9ifEPD1gsUPOvI4RrE/
65y67jr+bqmd/SrdeJtmEN8LRzlMiRJ36ZdPcHcboczlpozIzaI6J0ILfqH0mAjW
wiDTeBgtXzF6AN2RMazR02YGo2ai/THWLDr3/7ImeTPbo5o8c1eKJPydix4dFJoX
euC/R3w8cFAWhe+lIZpgwLE/NWIbuVppGdXw72ZYQbVSiJdVFvjwN/NKxoCm/Uda
Epl2Zfh01zGXh6G3wVzvvFN6ENqH4n6Zk3nSis/v1bdqdY+sKNMqWdFQVh73L/L4
yfLAKmUT9Bs3q9JnR+uBA+MNIBfgYFISPXbbn0vzWi088y0Hmg7J/w8mBI9tiNF7
XPM6JCm1HoKf+FxbDi1npLmGfJyxwO0TsDRjOABgCzBPsyysTc2/sWPJOlUdwUww
dh+cqlFjZWuoE6QSf4ZdfBcpTkuKfiasAd92JY2W34JhVqTI/gLofVqAHImZ5LHT
o47PBP4hOX1HG5TyvmfFS7Txk6BgPFOP6s+bCMBT+S/fDNR4bbPvq/LUn46CFf3W
ZwaAIUw4b4QT84VEQ/ksg+kP0dKsN/k2mFI6AccVYqMnZU8Urzd4yO8BlJJtdyIY
6cGWtqaWCOz6GvIWsrJMVSs/ChC/33Dcz0x1YL1iwG96bT81LYrjRTl40uLCyZUg
0NrHyc5OZoRKtxlTHwnF2KvMSPR6B9PPnV1ZJYGIU07krsqsz+7pKUPDQyogCT/5
rc+5kTFT8hNP8P/HWZTQFCWWdbs60Hv01YBdSpSjXZy97bR12dc7+D4UasAcpt7/
Ij+xDyyoAG0EW5TeVahYLISRXWqKKBq9v6mnYbdV9CZjRhj9LiywfNvPEjZ/a/dS
KBaNFoCNv4aYAv3pAejr1mX3RtAucsDKoiQ6+rX80j98Gtm7n7S1P4rUqYrsyRp7
b9gGXV/l8lXPL7i+ZNdy6R6WPA2MHG8AD3uKV0ny3LYZkxS0MHQKzMZp9O5ayT9V
yE6w+bhfu6TnWUpINBUNjKMbpdECsL5BtyeULn4/x+Pyhg3X+VCoZgHiyQPd0Rht
MOxknI+t/gSF0obg8aJk5NpoVhlYM52zKdFDzakSWt7Th40c3Z3LkoS2vQpk25Ec
kHI4FkPXDRqyLFZPUPtjZkIVLSN1W+dcaRPC9WwMKwM6Wu5jO7h8faIe7CX2qt5C
20OxqLWInTGcpnnYRCE8E2CZCKECst4Tr5G+Q4IS3Rm9IzWNKzhDDWpPTvaf7kFe
AsrZdmM3LM16DvKEKOAmlGOeWw4s+7w6mJQTDAuQ/a00NSVh/qmwYGim6CsYcBSA
RkK0TVg1e4SHqXkkPBYLnQlUSkTw3uBSSB/7QrYwkQ1oC/i68zbwZTuO5PC4o6Jd
wAqDumbtPcSCvOhT59XbIdt1yYMfBM7uYxYJ0zaH6zsel8FOhS7GW7gbApGTLpCX
6sQ3PzLUz+vbUctHZSjMtCYcesfzAU1eZBYIE2suYub9yRzalPBdp4LXeDlcxdCz
Q2wVY2v7yB63L+2HrJN41hUOgVQjRhad6WLt1n4o7JqbSkKbchUEUyFr/W6Sow1s
nCeAA0UW9IO6EqSR9BxN+FJKesnH9FjaiLYlpBPFUUIkoleVM8cVCLWs1YClGtpl
NQTGbhGH3kgMd9T75TyQI41vFNJGqWlESA4aQkMpqfUfnm50Jv5qb4kZ7tlqMdIu
YjNZeEph8zgm6zhO/Ay+ShM64GIAOjLZmGRgU2iZjYw5EK58Qzy1Xp72eZjeWDG/
V+oT+rPGs6tVKO6TTyaGh966RPFLzh9OJcrfwvX6ptuOeyS+yipMvkt8VnwbIowW
ihjnsCkfh359KbBw/0L6xV+EngE0q23Ub/ptqfDpEFPMAzOveHA5V7S8UinSALUX
DGR7LxV39MCWlKv+Wf6ySgLFNosq5UaIIkt6ABPBhKrZqKRrPw/akZzjl1QoLChK
uDrKXdpzNO9bX/CZBeV0hrlHVxdo3tvcoHv5LhVGmETNrfXwNvS5jvkSdM39GUBu
12ft6SOqSERW5+rdWjJ/fbXwazbOmNugS12uBUG5nv5ca001OOsEnSSChmMo2MJ4
/Oo9fgu1xkt6PNg9xZBA7y2HqOxIbFtznF3ACT4GdHrj6WYBOeTWS8Btly6/kpwg
uC+KhnI4T2zXGI4lynymWe+W+ixxKaDsbdUFksv3+S9GTs4aJFN2WrZsFiumBv3s
CKnz/GwGz91Tq8r7Pqpq8torl1bWg9l0UNDux+pZF1MFvx76eS6xJtGB0pfyPMuN
SVdwRnStQdbci3r7f4c+YTV3RbrV2HHOtMPECmmtLvd7R3TueUqHsmY874pv1lYr
XIRsBlo+NXdZ4mI3IKrAH8PXkIYDhPzntQEHfa/2nM9OIve9YJC3oTrR/CONoXjL
9hi+3be0Qxwq7cW8Ozty7x354ye73T0GtT2KnBlTmNjRb4BaV/wpwbwoVZjyNhN2
meAMmICnzjikyXLiodzD0qnraqc3Pf984p+TdDeRJKrRvA1KoBWBw1K0QxQs/3Bi
mUFrMluCIvjuUrGgEuu2vo4FqWzVCYJ/e52TaR0IzAk79+n2ugl2jW9nWhznCKIO
PCookwEjKMcq15cYJ8oJET1T3++roh3N4BD4beOY+/xuWmYkScoD4DGJGwCpNnKZ
cVOveWAzelBSbkpJZIo1HYZuFDth06OUL2gQrGKn1DYdalIlEKBd+ggpU/24uiUf
D1nwTi+ihwjv51V/yT6N6ym+npP631sN0TLsZiAMbb9bWgUhWj/BHdo098nY69FC
JW5kojUt3iZRyX6dPyngICjvVeDzwFLUTSlcej1AP/+cMD3qdLWwY3SreZ+ceB+k
1qv8qlQn1oQXX/4z7yFefD4bFfFgz87xJEsXr2l03bNkq17pQsF9Ts8ksVQBj1p0
k1QPXZ/dtsqBdszWpDS1Cev1qfhl5idun/1t+RxwzZ8Ju7hy6DiZwetDTzXAaUpc
WSyRfwzMT7WvjDU1sbsAlePMcrD/UefmJu7uaqnvHN+Xm/EbWI8cAf5q8w6wbFwN
FW5yp+cg2YHyqFxgxRfiviyiP6HbqbhPXsyKu4Pj8SbAae6EJqRHKeQEDM1yL2qO
pGM7yo2g4Mkh9YFocfXlAyR/RbtGocSeEvpmnZI6yC2CnF+7Fduye3GR3nhP1Taf
zmNGvyAarbDTXbHZZenjwL9g/Pyp/tbOMA1L/xDV8wQokWAaFpJndO3MfIm4n9Pm
cPQ7ftPkaGZypbE937vqxvRjw4FYltjpjQMhC6V9rIQ7THduvc/JgZk7mw8sIYbB
vEXEbaLKNgjnCWirayrzsXlKBNSJP6Q6xn0hFY7jn7I6oRhRxgREuo2vK37JAp0a
GQgKX76IOQ3WwQBc6C1jaTCdPTfzFNZCZPCtddAipXnVYTcCK244Y0uKaGTrJmQ3
uWTpl3GL1e2ohG3kvHMUHqQmwjJoI/zvkD3SOguXheee0chWnkIrYD2giFTrh5E9
/SeaORM3nbLZHGuHZrXmyJpO61nGrtdYhnfxQdJN3+uenNY8Xr77NF9a78/kn4iu
Zmw83bdssfkvRBsX/GpANm67+poAZ+F4nIGFnLOXTMNZpp3WocNepvc/JJIh0Zcb
Wpb0HQ8MclHnBqragPEGdmLdvwVV8lspgRXi3i23BuQE0KwMS832QyYGQEx5Tmyc
/hNUB00OYEy7qN14B+4EJ8P8CZUYfdbUiyBk0HIH3YKqrr0FBiRW2RJUlEqc/u1Y
2HWMc+VjHDymZ3DWcPEtLTh1z0TxWtyn17Ee++tD8psQ58e0OjMsuQ2p7a0NR02M
X5p3bin/SeIGhuO6K18fwXM76GiGU0vuRuUg01NeoxXlXPMWlD6At1jCjSQXKOLo
lgQfLMkvGPh8WYKFXI7ycPlECicvgUn+/MeQJD72bNySfe6rFW8QsHVnyI0wO0t7
wpIYW+QdRQzUAls/y+rEIeci8dXnX90GvOFyx6jhHJUFIfYvU2ye5F9zMwxQ/ZbE
SXkgQxW0A7ERwyaea8CucU+jSDeb1mw2x7FMzypWslTAzsE4DbufrPvIkh9TN23x
m0lW5PZrGTYwwMK3PGSfx1/Y8BKI7oP4wPD4WgsRVURZMm+xER5pVETlA55AaUSr
VZt226FhO1LaWdRYkK1TfgztIa8b9TDpwn8rgf6CTYJtEhy5Q8/xUkje82DoHUKS
q1iIJBaLRcq4tpHPAH8kPSusnjesxi70yQDJCsHarCMYiCv/t3JyxZqMfVWAOKR0
XEUN2ReQ1jeWZFMHe/0u40tABdB43xOMvZOHH1NZTIegGZg2aWEq3RrVcxmv4BWM
j3rmSDk94SMBVkYreKsBY6taIVt7ylbP8/oBVHzH6wsdZe20owfvQikNWbO4QVRz
d1mpiveMyDg6qbjKYuD4H2qKZQ59H6UqwhhMYG/rP2angYfwSYdJbdkD0YChxKpb
1o6fb+sFjc09AZu1QyV5jfrRg9DQESCAsA/02Id2tYZeFSYiYVir6m2TWd5lCFC6
1xvTHe3d54DIHWH8BEST2iysIQURTJss9cZ8Bh6IxzTkygHgvwGblNuix3VEbw7K
oclqbxGmVKqqswN4rtv+VRHIbo0z/RpafGjIsilLMeKtHHqjuSMqiOmBzenYR+rs
HtNjs2B4lmNigjTSphcK9+y+SafUkLz4uQ1mYrh79mhY3wzTFa3JA4zzYUnJuWhv
b7b3TVu9e/iE0o78qwmh1Pkhbi5K1R+tev/sLlyHc0E+joZMLdog/pE/RbMvOlOe
YTgjGWJIpdGhX7V32C6apUQmpny6aYSer06ktvpNoM3vBwvCmvfMXHQFIRxHsp2i
i7Rs7dcremn+YwH89Yr/JUDvziI0glhuKziB6FMTul5cUKO7pMvUdTEILpglFEOG
kHYtzKIJbd6DUypMdWcJ6HP+rfLj+U5BLUQi7PaxVRjq3YlatrMNS0gSdQhke3Mc
4nF5SBSBrOKTd1pM2Dgex/XlTV7F2sfBzoS9S3uaF5FhLontOn7UKVs/xIp3uthT
kC+9GaVmkUzuewrz7/TAUOWMJFDkeSk7EUjKBM9elVbhtLgB5Zny4j9dc+HqqPLd
moFZEHuKcYKKXd3o/g2JcPtDXOuq74LurDUFxw+WLlrXx9J/DNGAMvXg1pOzfu30
nOosj+7r9Opy07yhPb3w556HXe8YlvMaB8SjFDib6MtRE+fbEYRlmbGTXcVOlbIX
UbO0ywk1nICl/+UYii8jbxtxZWmSUGLX5BIZL3uAjiPwfEsysBxieSgcVFPjC42a
9YMEzHubMsBElfQx/XZCBNMB9YxeP6bkKbw5KCxcH9Bm/qOgoIiJkN/BXLyCXdTw
1wnaFtu9I4JST2T9VaIcEo9iOOEDj5kefoU+ieKv42LyDwVB6ZS76zq+KgZaFiCs
c0ctqXssqOw+8KcHdg3QoCD6kTqMM2kXsoCO6J3X+SoxWpNNxDHdANjzPAKWOeD7
gbOUMQ9nBEaQGZL3QDWw6p96IzIZtUZn/4LK8ORhPT8jjK6ayZCiWU50gBl7F9Fx
BgjTuZrBtE7PSm20ANTrY7BbDpiMz0EzjJRRHiEXOHmHRwg1zcunj7oDrNnz2RZJ
DPGwth896wsPiuAShAf10cLfWJoEH1cNaqzYF0Ji1+Oc6SU8RqV9u5r4AWmD1BiW
/WNjaScOCYasoG5ix8pl1fFix5h3DoPjgUO+HgdOugEbHAV/YgQ32PH4bGaF7zIA
EjrOOvnqBMf4JdPchsNNMmfv1rkeEqIh4iikmKc3z84PELKmfiwp8oY4kn3qB3Ei
a/RIAqey6YerBoPWGk3fk+IVWrilk00JFI32WWrLzB/tgrtcHAHznXBl2Z63rbej
65qG1FyjoaOCo3OEI6pUbDDtllPfYM/04KmCVeJS21LK7BGLgCEZswiFTitoNeED
U+yfe4N7NHL7Ijw9s/9D5OMrZ25cclzYX7pjIfQ1uCd3tMOrz3FRs9btE3861k8k
oCIbl4AHXL7l4RFLkbBDLNP+MgRqL36AkOpeLbdvGHFGyqk3Lf0FFqFim6tnZwMh
xKE+lvPJbgesZ7UztpLdKJiSh+DHNzd44b9q32MhAsr1IdB2O1ca5eotGsYl80z5
xPXvNf0ozmCHtEw5hMrOscXKRUYK5IZyhV6tfQKiKYI5oqc5Fse2PUNyb/gElRgS
yQlkPhKpu7DRfjdtdXFhoz7kMkPWx2UxAkaR8Qhok05rbmaMIrfZjvyVBZf9G7qd
NrG5Ak7ob+aACPd+J2bldwuAtPNXFNUR1faP6mq4zdr1dvK6zUj71ILJGm24iALd
MToeBg+bokYAmdBdOMt9ZRqEJsScgw1JhphRiava6eaCjaD6PRxtze5sOmni0FL4
rMlChal+aQhHEdmenh7bs1kZPiK8cAn2KVpfMq1n6EcFxu1M/YMXdQglYmMehqUv
hVkHkzE5L8QWhY6UnHof6kj2PT3awt0fhd5/ub7XFwZWoMHvxVU/ZWxUnfVUbKWV
97HbLTDvUimw3jjSp9T0EsxeQCAwpiiUSre3vFPO2sLSnSDfx9Ejhzcz5V/R5CIG
IEEeGJCsKJmvXCOIlNEq4SuQmpIX7eEWfL1qiaCL90O3LX74u6Uefufpd9chCS1I
Yj+Ub65OUm/Mbv2OsuTwW1jSoRYPiczDqGxRsjaNHWvkhZJuFsnWNNpM20DcKwvb
SNLVlfY83/ZiMBv6H3yUG3ICWAChnhvCoBk7sJeLWy7lEVobrtqG28r31LoPdkvR
6hDrr/pZ/9h6GpQNB+XEgPq3hbJq/n8BohDSgkuQXU3j8NirqBTtdeQdtR7CKtRD
6S6XuKI3xbKG9h+YY1Lm6bGeDAjpFnHyqhHi3YkVGRnysUIGkRkPq3ql/42cze2m
9FQCEA0xyaGTsgRyHUko4pbM3ohA1Bxcz3vsXKRS/ZBLMngGekytkg3ns3RvhF7t
rIcB9dUC1nrw9r7PBfpDmAEm7+YU5nHavSg70gj/NPzSckOdv5jeZZdPMxhvQPaA
YsBQA2v+gBZOSalG2GhvS4qV5bqIUO9aR1QgjqXoQzObBO02frsAO+9VlntiwyOa
211W/+VVmw87Y3LRa9m2MIoVKteB7/FWx/jC33x3jAY+BoP9M4UWwc8bcVXrRRJH
QhFXZJQevngO/6Fa93B9dUD2SEdQSG4fjfq7wOBNRjeYdcpPsjRqwGb43qZZ4xqj
62d4mUNY9zEIUyl0u+NbdOQ0cU/Z+jJUdiHN5o4pKQuxwt6BmDCYoK1cCjbannK8
DhMikEl0MBG6ptESoS92fawy5Zm91ZWNwaf9FnSCGBgJreeRU359NUPkgJkatp/n
ngQ3oXt7DCcD0F2LssYp0QS4yw5SkfmIXuwfy0kjxIdPkbGCqearjyX+RL5Yy8Jo
NW1WFR1v5RqKa8Xr2EYSO3rwz2xEmhzPZImcyEKoAmU5kpze5KYZo4OfS8g8oxHM
Z1QDmbuofoaNwmE79k/Ru5puuAEDhaQuQaX7dbU9KyEKmOWwdW0M5B3+6K6bhbb/
By1KzwtjzWsbQZoAhBOnnCSyHoZykX6JG3qmrCI4AQ/t6XKzhi5Rw6Cy/j/DUj1K
E0OVfDKpeF0xV0Vo8y8INsKVjBDopqsmI+8Nmg1cjHc9cDOzeoy8sfNk60of6Agv
EUZlSew3U0r8mbzOQ5bdQjxAAtt79GTLb9McX8VT/YcU0mVXKHt2509OS4SwiiFD
J95v6NUY4OKZdoMOrZ8q/94oVpIi0HRooQNDT3MTFUb5Okzjzh8BjYr5T9D+hrQD
KhGcsEOKk/3M/z2Jcv//dfNxhe256gdXRy/Mo35i6UJ40JHyLNzXz34n/CM8kg2Y
uhu6wErzVqjvlW04HEaEyt0ggXoH5zD2BLQGOmevzbaQwr1m1CGo8KbPQ3oSOEjE
kAp0NHSHRhyBHw95XZ7BBqZwyzCGqSxk5sT8lV6ayHJ9Or/yYzY15qe6Cjl2EhAZ
Q8QlwUTK1ZYziSAUgxen41zRI/1I0eek7JDVEtlOonsD5xwWYL3DLXMzAmF68lx7
bJpgT1OP1DQ/PwknHGz/0D8EJKJGuhqq8gxhQiYEdLluksvsj1iWt8Gig1FzFeKy
DCHbjGKqwZZ5Fqb8L2z5StIRxKqybySWn2zPlsOix3VKFjHSLA7QIPcyToZ2nmPm
TGZKDtdjQyTY1EdpWqw3ffHS5jOGkfQKKPQCpdfx1m3rOwdu1FOTYaOedXncGJHU
q8x4rP8uT1IDFwWy3mawTI/tWYhUJTzLHnjrcJQKTkGk6CMFE/ClqUa7ICiN5aoN
BbUMQpiAqi5yTvBk0fecnoZM+7Jd8uqgkRmFFJ+LtiEYUepF5GQ3pqEYFhdNuZzI
Va3D4kx4xtYD6c1slUzgk5a9IjScIp2Z5UPOqYiuRJhK3poPRzQPqfmvzSZTL+TW
+u31DLSK3H1VdwkT43U/XPq7aSsNsKTwLBlroEyOV3KRni9gjTBmF6xDAJ/sA6p4
IGQBcylAiUpncbiryOWTiZbI4PgoC5BJvBBQBFXu8c+TeePM6OgXADp9eDLNzN5K
7cs1yb8QEyF8b9UhsefSEZ3K6kH22NAiY7oC9H8LBMiEfPhv577OKTfgn+uu1bzm
7Cu3QwaoDMB+g8Qn73EffxquXwCu4y7qK+kFmEdf2/h+m62mwOf7ftDpnBVCvJRP
JJCCbb7wid0wcW9Q6F6+FoSPKeDCnKnF/8DXGRwgZqLzwZ3bbARMqFbZcYKfs/lZ
pHzeyAqRzDTEc7qf1F4avsZsVwHxx87gJPXFrKrcBb4LX5k4zTZbKfTfrr0mibA6
o672m1S83ko8UPUtp1njq2tw23QCY05PnmReNbQ/Oj7NH/dnREFcRM4Bml2Z5tmE
4TOezgg+M0MyHJkGdIOgTS0UWkGjGfAXTzbKDHO4HLQJfzxc92ur5w2jL8kH/YEV
FHQqVss4DCdf3YjqazxZa8UtPeaR68lt5Bsjm4o7EzqXhHrXazo7ewmOzgSh8k3M
/QDtUjQxxLk+aPkd/quvR6pwoRBW0RssfnCZd1ktBh3QBibVG6wwYv2ykuRdJQNf
NILvMVGGe+7SBJ45iw3sDBWRLA+RKdI8Ytjk0SwC2vP6kEApJtC/x6ebwIJ75L+P
FJYGGoy2FKVVwhqK1S6Y9fFq7PAkHJYpEKAlzUjhnW7BmJXYjM+Eyv8aAX4uqgqA
y+aiBS0gnlfi98nVA5SPKIni5n+HOonVDZKuAxt+p4sUTPVHq2dFHm3mCtPae9md
tEpPngNlpvPOIKgigl13Kfr9gbpQV8m3vz5r7MkMGes0Bn2uxhf8b3MZ2d3Iax8f
TExhWMVUjPgt7RCgKP3qMgV/k+Smztir2jgnLJMnSCAP286v/Uh4viqmmTgsUKWu
bydWcmS7IOMlTLvRtG9+t1Rf7d0qjktssvThhsb7HrQ2Ut40OyuU5quGdBiYjkoz
xV0fCZFEVkvuMdy29dGHPul7HMDB4FJ2Y6AGIG5XRbIn0QPv1S5LoBivwnKkhhFz
KjTWeWl/RJA6q+GLgJ8f+kr7BGjDEtTyLYiESNUBXaIdGCn7vdx6vd3eUFmlVrRC
NsRVqg3iwuiytf33e0g3YpekMUUC7nGvMx+CTc4Ba+TnjolzQGWz3gXYKfY+Y+/Q
RWHRu3czzqiFqtbDACH4iBkWXRjP8UR6uB6yawDk5+Yxwc1Hzdx6Of+UejBMTYi3
/HUZVE5m/gbZHfhewaYrm3SjMY2p5dwnyFIttJGP6RTbXt9+FPW1prpi5WH5dmLb
Fcngr+L4HeXNMTxSsLHQP9fC1qFzzt6jcUBqTrE9Hh/Z9VccgyL6/YBH4Oo65nP0
dMCl2kaROr0xY1kZKNljgkWlIKwe5X8K5hHcRpMjjkO9y9n4q/AbmpM9CSlIMRBA
EeAOmSpSEG2eLTh3fN9FWRm8SGgKtKIO1+Q0sze36h7koomYWQRHdBflO0uiB76A
ASDTM6p9b2cUUapAYnngKtisi+m9pZwKXYSVJPfjMdZTFTR8ex02NYni+uV9S8DL
lKECylyZOAmHEJyAd95impEyGy7FNn8IqKjgIFZdxFF0gbxiZfDJZ4doVTSgjSop
ynEcvR/0wj9fOF/hfEfRZ1YFAKUGF1UUjD/FljuA1PmFMUIEUxakurgocdhDeXUh
Z5/o6tpprzigw3WBpHLp5g6Vr45WFlCzhC8F3hM9KMGsvH5X58sZyYSJC9YSlRSZ
JpDsJn8Zb3cViow8pTbZz/Yv8BLEJpgoCR6aMMoH7ovdHEZpLHQKbAVVslPDyU+7
HIHFGQ1DGUu+NT/kxFIqy90BmTr3zFLIHv4UIuKxV9EBcw4gwmvwXPfFRMhYAGRG
+wSFM5hyCcflbGL8+zkFGLf37tq1yCB8nF1RcdEWtDTPfoSumHxQmte/VlYjBgqX
y76bw17w8W5Y2Pj5UbIKgtS36YhDkqKk2ep7uNmRTv9bJyjZ7FxjC+TBLQJ7YIwt
C/DYDZ3oGTsy2TM8Ce8PMy2lIfC4HtE2afadIGkoxbqZZZgWXR43UlnizF8FQbh3
9CA9tWXkDnRmPDALLf9dlNPi7sogGPKCirSgxkKHRebM3+MbN2nQb12/RSfrNbxU
lAzUaZZa1vcogk+8ALLwS635Vfv1UyPCOvTifM8q+eTOKSO0odiR/eq/DKIx/g26
SJjKQOTy5lA1GiDqpmtHvuBu6SjiDWDh1HioCFgmKXtHSysdWwFnZnAQ0x9OHFu8
xTh48r1ZpfLI1tm/UCqKHXM7dgoBBotGWu6tEA2Un19ALyHVSAo0mIcIDhGpOV2Q
ofGQevHWdx7bzNOkgxrsj0bsbWYe8Y0NMHIUFTojlGII2RzjHcY2jtmu1RDnhLca
TT+Z/DAbEvkx6iYuLy3q9uF7JG7A0054rz4m7RNVEwKEkFkp5Wa4MruWEWQg62gk
O2NRSv9bf2s4FoHWuukbMbrOQU8zzEM0RwvGzkredVl0vJuTdFmK5l1+TC+YYWJ1
XjF18h34uqpJ1EcThDW5Lw3pmBI2OrmtTUS9/UXe/FrIPPXVvGerpvkpsdpd4dDy
3dmErtkqFOf6ThSHMA9/5KStc70l3X7OtifUo/bTvDxMyY2zvv9Pk/ORucdIR8Al
cFusuXg7TRymIax6uHQvKYke318kZSHmBdREOqqK5PwhhMgYh7yqkmv0J618XgxB
XD0/ublCkvLR3GcTFgMU8kQ7kHsYJ2bVlP20RsYvk0X4qNlnFzCWI2PSjf3zwRnT
SLlaDWiAUmvA5+521WXXUMqsXjUtM5ew6dI3co1mPyIc95e5cC3DPzhbfZnxJi6P
8+kGpiIUNiAzLYIk9Oz2YG1agUbHhUwDZ7voZvCBWOFWkS8Mwh/B5W64rxBv773T
Yd5tm2jdok3KmRkmQk3ASzJHC97V6kxsp/w22Vdxn5bynWsd5S/az2i8UCzZneeL
UzwBAqtNzqlO85h6iAk/O6EM0g5GoRI2GpE7lvFyl6bWNXlsqiPgb89Q+s/jUATE
YWXbcfYe5OxIwBpRMJazETHF+uGhzfcA+EE2AS9oFjHvjercYfq+90VSdNPY71QJ
6qEyvjnhuEQNSpkdBfqrOTxy80wsqpE5iIwwVShvjc77nz3BrcQ6cApYLVyZFs5y
eXtPLXsHms5F8MUlDuHhT382J6CLwX3MwDg1on8sc1yJFhX6vDkyB+OWeUG5GS0R
1a+MtZoxcKHxzAmiwsPTFbZGolQKIA2e2QWsepk18fe2ohaTcN1N9iUfnezJkZLV
XuLsTHb/6DXTcf22vKdYOLJl1vZhy4rzFfCD8qV1UlLVncKh0c2QAsWtmpJWl/iz
VKYpEgBhu9dT5+Akej2U9gU4Oo9PFvoJt9q6BBR9fuxiJ1B1TIG45dPYcFBT1hym
2FuEOtqgulFeYrPAEfN0eMfpQgMpo/F1hwcHUpGCLZZZSGWVav9mSRi0r/tIAZhO
fsjK7ATBIzdNR/+VHOYkJIJTna29jRIzrNL9AHmqD8jx5MegQWcusmfyD8CxCpt5
QMoWQ4oDJcxmkraskWZk9iUTnouE/ao8FSNCWXsr5FR3/dlwMgGNjb4avsKb5JLX
X07wE5V0XjBL4OzXh3ZWMA3P+kxLxTwvEMmJbbIlUwbe4lQ2nk4yjOPQak6qKJCi
fjsjxAlWBLQTdf9XwQWiHXmImCW47cOW0E79hk5gpQbDIYgWLGwwO+1DqXmbZLbx
yZAoppyjfZB6rDOEUNTowE9ujv1gzbhdy2WEgWQx/VTzgBqTeww5PoqMFa89Ops5
XsoGD9oQ/t0QbAaTe+9isSISoqs2etMjqa4WOYyv1lVQOJ3mfLmUhtbKz4jdHKuM
IWcSLZJazsTRte0/MaTE1ucJPsrETawFPuUeEwUXAPiJTjwGgo3ypgWH0eLOBTNS
r/e+I8ItmXjDHFZdBXGDP1RlhVWeFwhP/FOLOFL7P0rA1npf1sYxXRNhBt7TFhgW
1pevGEQ5lezkicjRytcrwszzo58p7pCXblMcAfVN1nxQ0kE6lXSwykhHLPuq+CaI
lj61tILWoe4kl+eFlhU2CirtV3rAWV+wDSUz1iO6P/RCk+LGDgZpAUX4aNuQ5lZN
cLxDTMcPk7ID+5tuClldCFirU9ul36AW9L2amDl8qyXhggdqKXQ7CJNUDpEC/x7w
+1hrhSCWD9/26P0LI7dwl1eybHI0vbBB4rFxZ1wFVo2FusBSLUqnMBFbX22UETg6
3s2X5J3IUQ4f+rU08IFRc5McZUYa6EuN9oQaog2oB7ZufTmfnOzMxYd79hpwtV01
hhfWcAUzvyV+8mgNlVxAjLhzl0g7DF8Ayt4+n3d0AAuNXD9RCrxrXEKiYOvjUoF/
Pq8Lg5DKaZHY1lcbDSDxFWnNBlFw8YAmX/9x9wA4GHZGTIL80W4N/ODbIMM+3U7z
VAFqkMTe4uoNByzGtLsGUVmMNMnhy/LODpPy5uZ1DQfWmS/xWDMH4fANbgqiFq7c
Ebajc2jir+FTjuQnIG2iRGIKUK9cYkaYZlMGdRhz2TkhmfUcLjwKfhmnmA3C26zT
6ow0Vk/9geQapSYaXmU4eK9okx52Kch0mp3CbUZqIBJLIw/Tv0fLbq4NhipwnXUj
ubeVybutL9tKcSaz+YCWPcvoVFxxzMbzREyQDTgQ7S7zH7YYIPtQ+OTJMHhY0eRl
/BYSewe1J42VrbsQbBdSgSl0mI/seiwKLj7hwNMjv/v2iD4Cz9FNK2gb4n+eQqGw
CBvoVIY7PieUcazwl2Ny82zAAK1ADQDDUQaWAw5XZzFbskUCm2sTn7I/O0k1+iIA
pMiabCgs22rUksOer26ZqKUIt9jQpGCgS8rJY78vLyRXbQTdNTUQeP82nz06GFMX
Z7jxcmGK8yxtd02et2CX5Uw21Koz6+f8QCL9WCOWvdvLDrmhCxX4+kwwH/iIOvfJ
8RcK4P+do8c8pHydLFp8vArlbWGnlPrs62DD2sQLj65/a01V9hsodvAZv/RuYLA4
AL9Hs5y0/7F7xsx6XDplVNDH7sHuq8gxJTTrKYf79Zf95Ce//ku1qyBeCesnmnrP
e2C4AT8vUVmF7RKJY5+ZmX1vyEnUGXehf9EGGxpyre7w6obW34OSA2ZQDR9iUzVB
IpuI4/gasg5Y3iYzkCr4hjKqRraZ1oPtRAomTjqvj6DEAmBBxboWSWHYu07Z/utm
FprtErtkzKJ1fIk0gG1JnVvYP0VoyePVdomBN4gWF7N94WRW6MEPRPQZ2ufA8NZ2
WLudtc/DbMcTmZTsvN+RIVuQpMBWUhXyJ4FyLhOkJRJMq12Ro6jDYnnMD50SywwC
KU9lVmX9uf1yKngBsLjy1+BnivEfuBJcXAANRambpPEjXkyEeXuUxhRlgMfaFX9d
rHY+XNS8DBLHuSl99efAoIWqhPxgsGdtPRh1fYIk3tTN5cUGW7/MuvUEPUJ7aRv+
LqzOaUcWfjyJBliaf0mGblAZ0BkQXVr6UJzRIlGqcdHcEMh2na2qUyEj25z8ncbI
+1ZA3D1D3Wk6r3hBqEfspwEZPC0Ag8ewbwRyRJslHnfUoXOCg0o5ObymCMdBGl8V
A9kRnr0/j3WEZT2qsmf2Eqv9ROYA4+mNDJn5i2kCE068XhLVQ/27eIn0FTpRggsl
a1xvSztMIHCvLc8v0duXfrFQ+8ggQ4v164V55w2YskuIqechUoayiwhMkFeIYJGS
oCNVfO5e0G7d5E7MttFRnlj3iUdZB4Dc83NhshsJT5NDdwa3pEdSUCuAN58/yhdM
iiMTxoY8PgBhT9w/NbJvoHYLHx+qWcsyYn3IBG4J2tczmBxRdtU6socmDDYB8LLR
quYqv41/VLKGtRC/Zw6zWkbfQc+QSFWowMlsjKodZerkaM0syOpefdP3PM0SLXLB
YSJaVtsdxHA3RSJ4mMU/aFb54YtBl7dRB7sl0LtuESFBMTKkDi3RFED9XAgChDXs
/6sFF/DgeXse0lksfLmhT98gUclelrnYbegTVNKdaNqCGGYtrGWzMsR4L6QXBou6
E8nqgxGEdoWNIKwyJnxDijgiXOHzVDI3hQAOBWVUPzF2Qx5qLAZouyqArdKWoxDP
dFJNb49/00CO+3zMQD07ZUmpv9lWQRHKo/2uz9Qm/2B4S35s7Ke3/bmejDI1r84E
C4FP7VqM56ZFn3cpFvtixJdUKBMdgd45ZXF5RxD29I/w+g3/ZDR2iMxJoEf/3nnP
3fRBv8FJF/toEi6v+onNHHzfUOaBfUK6X7Z8SxA9XEhVsrqVuc3HSnNNmn5UVwa5
2WGIsZFo3q86HXiRF1kHZaMs6j0ial0DJsZheZ0jsVfUcQm+eFJIMjdWk08PYYrN
ENCs2pQe+WFs0DnhrYF2/BZQy+z/R3Nak2+Vtc7mQWayRb5L3cGUMP0SU8RnNrg0
MZfcAmeGNG7bNujE75ym5/z7jA3aEz1cekuhgnHBC6c4H+MCC2GPHkft+95VVKGp
eTRDlJSbKp3YoWDCOFrOMkadNeflW9+Qnnq7SHIXN2fFw66OBuY4cVebD6PUtMdI
6Y/qo7Q4mAhkVbPxoR5OynRFCkdUs+1Gu/LQv6J6/jFyHt0V7kKkyA+ryp9/5d9U
pVl0H7HGc4VcrgBwmzlPAHCzl0+MfcbxOJszPofVC6uM+5s9XZFqYMemcLNyaFTD
SVd3I9IvFWY3NHI5HA1+l1RCPIZ0nk6eWAz5YvjqilM/X3TBCoIsLDtY05j6EMeo
nF9CCeitpzMHHQclDGykKqKd4u1Ax0ZWRHBksZmQDNSsNxPDz1TTOrRGIW+Xj4fp
vFAldrX8jSzvY0rJuJI2WDB+ubF7bR26SOfu5YxCNwXy3/4NirNa+JM9F+nZZytO
4LV3MBNTzGuWiENcbEr+18Xg+xzAu+RtlsZT+QvTa9zooWCBde6XDDZm622XtGrD
du713OoNQZX/BmuAs6G1zlXrM9mFA+kPA5WqU8ohiElvu/gX771+V6d4kp+Iu04P
zuoGrrSb4dDD4jTyxQq/ePBAW4HDVDxMfxAD+KfcvOv/ILp2D8k68iUzb49nsbQQ
PiDpsCeUd49fD4rIKbnDdOrNt3sZMxWXit21EMazaFhxAG3hpkygcURL/mZEnSBm
O+ktq2wKX5WI7SDJn5EL9uydHwNKxSNsgPdruMmAt8rr/PLY7F2PnkhuVTgmjPij
7xzzULdzlSQGEiXjucLjCA17R2n+Xygvb7E1OleHm0S7eir6QhC5vKnSQLOQx7Hz
2KUlZ0macQx2HRfM00H1os+yrRMwjKtH6MIclxaDwEeWrx0DijNDTTnnn7Do941p
V3qmHDlOnCvJdSVIiqKrmgw+dxax2eEKDWRU7MbTfwnjqsY9TGYxVhrYUHOHiW8K
Ul4IniA6jRg0XNbWXOh+Q/dvXdnuSxo5sx7wjDN4hC+m2DtoBRSNDJ+kGPuPdT05
2wGAQ/XPskRkyXouY7EU+atbMRy03MwEsgnsAHU27wF5h2bKZS+IG7mL8IEGLo5T
8KN5utd9cvN90I/vLKkr7MAUUK/MdG3qpnzpKYnC2rZ1kKAtwilJ7V9fXrx9gtOU
2Y03eVOaglQDOfm/DQxo4dXT5K00qzW2aP7JRC6rgKgYkGwHs9P1qW0NC2ojrAgQ
mVs2DV9tz3oN34J0mN1GTe1W3/4ImQ1XEGtfML1NtRk7TqWPKcQHRwaRLsz+UKOQ
UTYiB/4sDg8svi7gbaaz0/n+nApu5iTCTgrWKHb33PSDRTieAZrEcWPoW/bIBJGn
oT8HDyzM7nlw/oSKrO+m5Iw7ruoapQIOh2AfNeI6u3LRpF3zEd+GxHRPhjdolY9G
tvrC2KOepnLI1KowF0TEex2iTI5Eb3zV1XCyHKhdtYRBWkfQE+PAHm7bnzB5OyOu
pqXTSemIMdzLEIaaYjaU54JNXENXzSRX0MBFQ7FotRJEY2pvG3VpqnfLUp/9uypk
J9nYqCacRGyuRpnbu9/pZ4XoKWkVyjh+/WpbT0zCw/EW0AYKgiSFFOVsQS8CG7wF
khHoVG4Ahdt4BTHgn8qVk9CuUg1Q5SQtDvBd21Dudp0d+mWqfbEkeoLpYuwPXPUK
kZKCtGkv3xfinLkL5A3y1L5F5Y3cJFaGowfcMywJNsgakSXyIOBrwNBsBGofZ9C5
HXXURWzb3TcyBIu6FAWG7HXZynulmChYWQEPozm/9qJecqcvym8rJk5aucenUkTB
HMwB/SOuctGA+JBFcfaf3jaCbgdebvzPb31elmyGMhnkobF7R8pOxtYNuf1bWZJb
dsq0EkQuG7T3ShO8gyDHzzaDsS93zDXJnDvHZWSGy2OPnxrL0CJtqs+JU14giudF
l3aY1h7cnLP2ISBopj1EfS2w9hZdZCFPyo5qlgUErF9zRZSBAABv/QkUd0yB+mvs
eTABsGpj8/VZEeGt//2Pp0iUlpFyz9WNv6ZmW/JkD7v/18bGxwdUemLAEi2OvmpJ
z8IqJgJULFglLQvzXBYHq7LKtmE2f14qcDQNmGiing4l2Ekh2JcH80BaZbGVTp/b
u409avCeUDMS31TbAkQpj7wU59vQAA/5PzwdZgrhsuKZc9qMTlWSLV6sXgGoa6W4
7dS7cMT0XqgqSRwtI7NqayGewgFvEW2ceM70XitQUrrzPJIoKT0A0rIuDGWgpE6/
88WEokU+Sd3/BiDNOnKKvJHXfrpQkFiFxBD+fj4VTATqCh3VC0QpWJv/BQ1eCsQz
kxyMMvI4p68MIUjjgSGmTeol7tZgFBilt1zkJQP2Qnp4ltJmwG1giC+Ve/dqzXcD
DUjNJ+dWNSA1D6Q0QNLBFOkra+5o5DmfzJBikNdj4Uv627EZ1itEyu+0qzzDpmrc
Gzjc8ifqIyv5p9FHzXmw3fr+S5dVR/ftRG/O4ST/FxqHAE7RkLlX5l6el4tC5Pic
O4XA5pwCJtux+CDs1PJANY7KKljy9nYxxAMGtnmPaU9RH+m01cwL6l2M3iHjkkhs
lei6q0N9eWVegMN513g4zjtI93zHaq/HDcsqHchT0cWwmV9UOwuFS5+3b/NgyKcu
ugPb1hsWei60kuU6tyQWZBn+AIJu4T5itsaDmvB+V9dWhZC0GS0a5ikfWSaYx9EX
tGKb2Uiew/agPiIzR6568QDtvgL08wafYMDP9FyEjv8SezbSiu+gVJF00qZ79zvG
V7lsi9hpcewKWBsFNk/sv7Ps6l8MF5Gdvkd0SmM2kPrE0dvF+R8cwsYm52m6OGxu
SzEDkUKEkJXpcPC8DaSyNXHYn27/lF4dYLIEd6XUT1sdZhVp/j/WsRI9FJJxs48h
0zhOYXarsFLwdcixEY7hyA/ancBnUMqrMHYP/Jh0CqAUnOrJahWSmt383Qke2H9O
uiKPCuDEOXiMbzIGyy/6nN2WDMfkRj6tNfOPlPCUaCGvXOJCK4oWZ3G0f7s6+BTY
U/Q7oRvyTzMRPH/aUpOA+En/0DODTJjYbqqDmyCZdfsNs8L7w/A/vlCQ6MDXaATL
L9HlB2fb/6dG3mMq84WXduLqC1/aMw3KJ03F+9LpZztjivpLrV2TdN44fXkzC/rv
A9RMRIBca93td7YZCCU2gxncEIrEAYot9ctEqy2nGezAuANhq0yEp8mgiziMaxs/
p5DEVO1BUD8ooY6Yo9tPyas9+CQbOjY5Z2fHGIM2k46XDNXRR4IDm1Kd/WsSeLZ7
rSbDafSo6uuR84NaISA5ZjIK0E0juMQ2EeZ4dq7F1cPYQfbYWS7z/iwbnQAbhNUI
+TvTIOw5CwVv/N1++E4A8lZHYsbDOM3cUHodl7XIY/IJ91xP1ifSQkW6p2BnsKFM
C4cwhfmwFBnSQCF8ScE6dp6Kdr+W2lnowncWrn73DImPQbYKPoxUZUDOG5wviY/T
Rhc6GCEg+hU1haVB1Qqz/lu2SQz+gDWTuOIbXYGcXJbrwrvwFi++qGUBBgIZHr8y
uGcLZRlkhdHwEK1/MSML+9UIsVawRvQCECGFtvC2Egb6a4u9atRYbVKLz/FjRAUY
yHo7eWBV7jshnR10cfkgtUvUJtCsI7JeWaWwbt5R1/JScK5hzq9K38DpH4uyzzpE
auwWD6TStQd72oncJiruECN5amjL6btxWZBcX/fBP/fl2LSJfepE19BGHg9Z5ZPw
ICUi20h/yaOAs/Kg6UWeLjaLSP58J6HZdriqIHo+VZV7mD2rzJcyr3Blk6NKE6Sw
N+fG/xS6CK+UYqp8Y4lcawJ/G09beAnFpbgyKSjyC9f9C1/AxpHTG1ftG+fjUzCv
52qfdv+6qN+e+p6u3/Vs46LTDzCH0Y7mC8UuzSqdYCpHon8yI6ACIvJPSd77a8ST
e8wQ8WZVGjnjVTHSCAAuKNx0YpHfBFyjkPylIbLfnTPkao3A/CkMYX67qU6RCYGm
KTuS7F+iznXjCMqRhllMS2grxiN/0CwCI3W4oOGGEiLPLiDfm2btIII1ojtHivNG
TGigV5yB1v0a4665POFV/I/GJvOKYHRuwZddWe6RAOh92qCTEqTcSVB4k6rZNUaE
Y9fCvqWaH8Ng0t2z0rfDbeNkV8K5hJFc7FSzHg0Yx1819YlkHtE+CjJxE23pBrIb
7bnyVUWysN+5kh3idvputU8MEHARyDm0L/S1CpuCGRP9FUTN2eAt18/69h+Ho37U
3vFhhCQW4Lz+kXSq3d3VNRPG7QuBJo8BKmkuF56NFl41pWS6nlXrucoHFzZYXn54
Nc5riO4Q8iGqSUp+aGzNZDx5iCh5c7ehfcNSVRPcabB3b0tSUivGYB1DW9MyY7Nu
c9Jf9IMZCCEAeU4bZmG0g/m7d4QnvydGWJ71Np9Qghq+Gy72jYFlrLuqRPEpjNlb
sOwcnLVMfeZPqoHFDwFg/i2dLyULfAtOsujgBUqX654kuBnuPskjtUKYQl9GaeNe
hpfTpULUjkkeN2fMuzfbBSlEycX1OD84YmvyxeT67nE6q7gJSdSCjt71mr6SqCQF
L5AhnZ2hFYx1Q31DDV4avWTNFDpqvnvNuRWEQlpf3I3xkVD9IV2PqA04Gjm+t5Ol
3g0i6/j7mlvZOV6SUPwEHVJBhjUjjzW31b53IxUJ7Vs0RBZci+SwI9g2tVClWqzx
Yv/hW/TIGxglgNXImrk4Ib8ZnVsHwD48lSOiT19xF1Z+BMgACB6qZbrTg/6JxUHq
c5vMO593fHf7IuNbVXRMEKvtQCIcVCPgM+RAv491t25pMkgJW83i4X1KnT0pGJnw
XrvjPCS/yvVlBU5hGeL0b5a+kQTSwpAm08SkBv/DBl4ibwNYFEauvljjTeoKQQuX
IVU52qsfI6JXfyodnnBPDg9vIbnKoj+KNdpKBY2YAJAYH8yjQvnIcAlR5C6h+YND
rbnoROc1TMnmBCvsX5TUld5hjO4QOmSizHYv4cXXJm1/avXywXmQ5DkJimCPTXhx
TSDSH3dsOSILAHZs1ccO3DgG7lPf29X7tVa/R9gw+7U0b22g5NSGJx7gKEM8+3XK
I4thCxXdVUq0RGQTpswSfpUupP1AxPIfcUxLFrKZSX+HGKAZupELis1J6IM1G7ys
/+ATAN3L6fu9BfCG0q4LTWslx+ENalJmYgsoFMg09gilji12P4IC2rUNGj9nZN9R
MjFMLqe6dtP7ZCMUxGDwcwQcF+kilmqQTBUHWv3KOpsH69VszTek03jB2y0vrPg7
ZR5vAV2GKhi8neq0ImvToRAULxTxJUxTK1P+V0tD9qNsJ6AZ+fK1owgGfadVp9wI
wguuQS5oV4EizrjZcm3/9SfuepC/K+qYi04rSd5055ITe8urnb5yXcGnipEfZ6RY
UrrxIhs16Du7ve3uEJ+tO5khVEboNkdL5G4U7KrO/8nKTGJPPI7LJMyHgHMC3X02
ZlavRrbrxpVm8SfD0to4uC6a1tT0VqVGBeJh4kvMlK5MwxhzzwRIk20/TIBezhAU
NOH1QhrwOjXI5hHX6mYoFHruj7qvtIn8prAQSvhrUBob0E1JWlcvUwr5IhFdfhgk
GrdV3Oa993sbNxCpGmMF3B9oWd0XFX/4QFyNWw+1+M7L8c7ewQF4qZpZW2JqkZ8n
7y3DM8KIp57Kl18QkXg6zTZ38WZgiU2aSVRgujf81jOFfSNSbVsLGBjOVD28zzI6
fwkRpfiteuLuQ+WN3/SwumdmOcw4JG8W/HbhNdnc3ur+lXB7P+UWBb8h1C2pUlIl
guZsh8/WzBgZtGs3sq0nj5T3xgNjHikPiI8P8MOumjUCEhuuR+DWs7iGCzTwh8ga
Q7JkKPSukuF3uxAlg4+QAMxb2jUStkOZoL+CmHWvOsLtpnGjBWRXGSDatiFJaC33
q3CBHj+nB5wUrKH8ANY3BbT95/BpkwMDBrfgEs37zV+J2XNIuGA3BE5VjP1FLfZY
qMxwAIdi1NkuwlftbeY8bcqv1246ga6QIJ3kT2oTPpZEJvFBhsY5kRNbkH/sr/qD
3VTfifwN4tTsOiFaFZNEkjQuvQBpvU7maqoMgU3i15HQ3xsith69ZYbYYfcmkJGg
yJJ28X/yowE5uxQYr9MSJnGbpgF0qxUSwq9cvzBhQivM49NsNi15dPGeZOKnOzH4
SY0HJinu0ct0yULOwboeT5+Kz5JaQNhCP9oG9y0omhljgcrTOXEH6vEjOpQXSKRj
PMgXs/z04c8oI+xHlvQ3t5r4ihq5v1tJs2/vRPBp2BH1W/kA6af1rvUARSi17dFG
rzHhQuzN6fOl/CoEOp3q87Vin7yHwd2Ky4xD61r8qFTOaWrUzkta7wxifoDU8CVR
9stwEGMbBCMIWYKzcQuoouM2TWd1MQ/VuEnwWfZsobEJYk40ApzmM1jQvSVUazfI
fMMzTJRIz9MZ2Q3V4lIYtp7W99vahDrsHFmw+YSJb/20nEJ/sHQUuwoTSsLiD3kD
IbRL+dDJBdrMzeSK33PSTuTfi2HyBaNIh12F//ZVOa9dRmp/9XS9euJBTVr+AsPU
FiXKdlSx1tZy5oPJBG/RiA0lKNdJciTb8UAXRIY4q7rQtMFhuiCSWz9AEkd4vCjt
k9j9kKZLMgKikBno1gIzTMwymgvOy5ietsPUZXFR4iZWRQYbwuIFx2+IAtxUb1+V
SjQk4bZpGwpxbBREwIFH9ScRtuvKjDH9Mb8kL8HaeGWMte6y8FRZNRwhRnzKMhAY
DjxjnDv9b4xxFyvQEeax3FM7B8gXbZlot6lkjIG1La1Ce2a7JCHLyj3yjtqpwLWP
jBlZIG3ZGxVtXwglZ/XVk1v3LrHXyzuenbSNExCNK60dbHxQVeKdjtTicGReUT9R
xqGqj6m+7IOxDntGuZ8d5FCJC+mk2bJSdRiYunzDZvPIMAe+m83XXHtHY97DAIfZ
00I8lpI4wtvFd/EY1u2ZbJAGqFXHnX/uCf/SP8eCSMkP9GnBqAgyKaXVrsX+TPFJ
0+DWL4CgME6NM3I4QxlXZHoRAlTdH3qG1G9db4NBWWqFzHEZygKFGC/RJ9/N0Ww+
LovdMw2oQcMEmxc23AVLOBXJLKgh5DpXDTi6X+hHHwrHFCWryKCOzPkI9eIzFSAO
1cAp36atfjtLFfjinKC2QMwDw3TOnseQB8xZsW3RN9wUHyHzmFUvUbrfJVCOdfOq
UNbhqbj/fv9fDpjD7EPANGWTghXUL/APIwUQc9tLxa3kUml3nvXRqnKq53NKFe/b
4l/tR0MgzMkt8P+TYrSEGnst7khbXuLm817GGdeHjQaUurWcGNmsGs51GVZ7dKoP
nyk0Wi/Lu2t0TaLVbZXlI2uTwv3VdQYEHMv+m/1HE+vyZL5kstNuaS5pVyUL02fs
X6bZEBSrakQ09Wkjg9nzw1wCnhANwrt0r4EKPQ38E0IWvC/6k1pz1cfOwnxagcxM
ZlvA4Tonvu4TEWN/i3WzfFNTsg2G2qRtTtytPx2NfRMKdgSOsSzvttO4bFWrCgxa
qXDr3sUyYmIJNrWThZVu6OmtyqYlGnzz7yB4mwSuFDzuz7leSkw1riFUSHXSfHs1
a6TIbKiIETLyqiokKuoVvWGVHsvH4VUvhfbqHABG4iYDvlMkQPPZuuebXehnarlE
yF/8R5pFq4U8ExtV6Nfel4R0Gyc4Hciv4ZTUh2UnwRWFiGu6Y6xiRrmLdGrzr7IH
h4rAw9SML4G8agOnVSijBH8TGTKrPYbYxIAGxUm03Njy/6aF2tL/pcqbRduj53ou
N404BuvtWk/Mv1etmz93Sn+RlAskopF/arOlRNAtdCB8TKoBeGhnMV4CS5f0yahS
xDascMRypncNnWQhSBVt8F+9B8JZ0PiNosYJpNxEzv3IpkSfHIt3t0NSaDo9nbHO
E58qwhI9VzlCkXFsysR2/gYe1q/i+4ztdWajzfww6+YpUpf8a5PY1zHODyYR4FH3
VZtwNDpUohBxwUb6H3RdJT9+0eSZqCT1PgfT0jkyQNEByRClp5v5WfTEQthVNr3y
NfDj+AwFSAtpb1BTOa4DpRfExsZzr69JkPsyLn/Ujhv7aOqAm60Vpire7E+I0SdO
CRZX0Kr+r5TjJYLocOPH75O6mfWjeBM4MPbEXvqtN273ygTBvipMveKuvuA+YXqW
Y0O/NfXFxJeB80Xc0U3ECC7Bh56TWZAjsWxjbpv78/IFRQxbALX0KurRSagqZE3S
hx/2Nf+9mIvsgCy3Nh1shKBN/Uo0zb3gRjsbFJ7i3X0LABMp+fxu51QxPkfuJDV4
eguCSAQM8FzlTxUafZ65NwkMyoqJLcP5tl/jKF4DbByafoc6BfE/odjewy36kmcC
c146iCZBDXA7VLuX6xTeeHfObMoISXXhNE8TbQ+C+x4qZpS89vdU0ehh1T3wx+Pr
3CZ8V2p8aaAO7mqJqzhbZAi8NI6j7GEdMO/XKeRM2WCePF/tLQrMHTuJYzd04bJC
txAiOiXKpuVq6Dd8fP+Q8KBcSG2MgQ9ajzbk5awcraRPd0cEOj04roHcG2Ng/O1d
/iXiO9ri2uezte61J1ARaJLRYjyFnJ6NeLahGCE7iLKvkpHQHBIJbd8H8FPKzvtM
TxTaqguR9rMQ79m9DV3FO1+IaSVnSLYKN0el2C3WJH+D5iIPeqSipaWlkEphw0rG
ZCYIyCvHKVzMs8N4FTG8GlaGsJiQtKZGWu/18DLmKTS6qOCyB+zjRXoxRzUjDHEc
PzBroutbNlOSFW6bwtApl1/+k6fsIeOQTT2bybgxbmII9y2/rFtAS8f59SN/poj+
zuY0AG5GPFLFaoj2bX/sFdCxNQ1cPw9xvO/5f0/eT2VfVY9y23C/EsIgpgaYlhAs
QKJjgtQHynZueQg3t6kyJd7SGlItgnTdesljKfiuLUur/gz4P3Xlq5kd6Qof15If
+jemhHrkQccgUJ3K3WfDr+suBVNrPpQuo8WVrHY6WQpKZqlXuRS40sD1FJdMtVFm
wc35TwlO2w2nvUjz/7DBtJfbitY66TW273mkc+ah0MB82NCZRoapdnBBB5rYsWWN
SO5vHw8bZRBNESoQHIxQAcTs8PylZ//LvUOq0qoSWd9VQ9TW8sXoBD1Hr2lGdArA
DL5ROprn1tF7FC6tebJL6WfbOuyccV8KUz4KuzkDhC8oTqK6lMuIHqZKDRfW0aCr
pWZxaRtoeRTacXx+MYITvbVFdMK3fR7ZGOSG3Ejjjo8OMQjIEoghB/c6tVURmRR+
DUjkVV+nXFrbfOj3zF9J+1GIKNHYT9mP1RULk0PkLiCGXH33X5OM6kmc9r7h8T0c
3L/96H4IHAyLlUioiFo0T2G6pgNAg33DUYP5x+R8eVEUldtDAxr6ilFS1z4wleu+
OuoUlytu+q5jLq0C26nOFC2oZZGV1SEgQ3EghhjdKmqVGCDLSqnEiIcafzsBxVu4
MtrjPhHlhTsyudREx0BPWVBGEyRB49w/ZBYVMvxf5hjFqtn0RjMdBQsiA7A1I4rw
yHBPei4kW9OXvXqc2avLLo83mBJy9Ech1s8mHTpeje82N8EYqevbwnASzhoZ5OMq
Xbt7YZCp5TwAbXgBRJBDD5nYlafm5ftTTCIftO9kq4xMBDxoVqKeaoV6WVoNh7SO
tMv2sbACfB25cbNoE44Z8N9+8uraGakQrbQYNwTMN/QsvZdJRU561NpvmUCV7vwH
Q0PR5FpfhX5e+qhhtRQcHZBUJXB86AkdWHBSyOKMape/sIV8joaAW0kanEWyhKnZ
9Hjg3gnLJ4qg47v92eu+eNkw6PGa4p8JWqOVi43OcGNZtZeD8PTwGnxKg7H9JHkZ
X3CQyjA1d9mkWaJTxHXYhODAPRzv+IgOzoUhzUirFBfC+AVog1Jklm7OttfMy3es
0DuQIr//pF1f4khCh94BFBaSTA1UvveMyuD0a3hDRhDQtt8DA8khj2JiEBnvdfCG
frYShvW/hum7G67gxNNFzAIBKllL25s/Txfk62qka/F+WtXbSt50E/oXSAnvGyYn
si9SR1snZ4jZqIrYZjWhDa2BRM2MwKvteFct3QjCeSZhF5u0ihXKd6nweWILGX+D
ZtgH8zwwvGbvIIwagq3MayZdVZIJA+WC2b4TQciC5jVWJTbIY7EVc9uZCRvPPipy
L53aDPXbhf0Gb+wxKg82V9tCy8Ip33SHgTCR577m+2Ovrko7qSB3gyJVTfgSHRLD
R8OwfCvbx9ZsqNT6BNuEi4fafPpIHvE7F8qI+nOiPTcu4rFPB73tYbsx7zmo7Oag
oELRo0pAYehO5i1zaC+MslynuQaT6Inj6iQwndXoHX0NlFULWBRbwhEGMD6tEKLN
5xKMgcK+x2hw9W4WdgZwtqn1x4Aclli1hBsoO+dM4AWDKXr43K1379rinafOwQX7
o62/xxjCQjsQQ3AcPszV28CICjVzrbr+EChV+gLEanddb4BTL8SPEMAfoKr4R/0V
zRm+wtRqvsCXRPX9nB/ISvqSpibFZHYhr2GDt+3yXCz9HyOx7X+BgFW/hYfag3MD
xZkeF3jcG14Zi3O9w1W6nzFvMIII+VE9q0WhfsiqS4rKvOHHcIn8c9PQde4p1KEl
93w1MKMaXKWSweLzyhwdE6p0nVeJo96HZAPE0gSHXKVoVpF/ifnV0Uhku/N0mUl0
J0kXDbiRWthEmyrPKLA/c3w21s8auFLgQq+fhwAbEaqAPoyh2MgHI+wRcxHuJCUx
JDgYM2xaMVgOmdqvMY1GauFDSiW15iKdc3L6Lb42yMI+03QHq9TUBMTWspNgPXin
ObWrq62ouYSrObxwhOOaj8kDjjW6nHqkh4Le0b3f1s73kMiF5YsLBliaeGr6C45o
uTb6U7DDIfrqME92tZsKhzhqK6p4Rtuu68ybyxQ6E9kztzHGfP+51X1WbsZFoizH
wk5n2cfrDTpMwOrYAmnKfNeMSETKf4Lp1v+Z5ayYd9Db1oV1LXaoqIVrthaYctUU
pBfRVy0IaoGzn5W9kuXasUuTtNSr3FIhR84XzzrlLF2Xyruf2nD5i7680mz0rqq3
FjBS9ieNRKPsH2Vg0yTi20dgWFB0lDG2OQrm6gT7ze6J1tUwjw/hyx3ZYNWM4N37
bs4KhZuvvPuk53glbomjSsgPFdyMyHjZF3KY4R1KECosmb08s0F07X3SXbeWWjYu
BRR1ryONqh9y3gB0B9pO48EsXuUuuuMn3QCGa0GPh8f7+zxIogI80UhYVYZk3DBa
LzcHO3imhbJUYsMwXT0uTR2bnbOXELvGgSnovxu/wFg7P78MrTFl+CHYGMEdLB9b
ySU4Fo63FjZnmhFwcaFI34NP6nIWbLceMsojBgtMswswrSRtA9YnUjEYfkbaGRBd
NSzLV0hw7HRoiBMv5H961CbhYKG5cQ8yn26yYjFi7zQNLTAfP2ulW+U/feNwEyfb
pog0tNQp/GKveEuENPJdw9EwcqkPLDX2LfhBNUvF2tFd2EJI4p9AT0W2sP5D8lVe
jNIHM0QkUoAxOBhoaIvo8DDPih2m3kRk5HTiuwIIaWyXJ2GMqQ+bXA9gSa9EJEZI
hqFoNA++TQAEzd70b6IyIBmk7SQYHP4rCc1iMCEfHa97n9ZHPRFjUL2KtkWc6yqP
Mlb8Or5yvWHJZxNB0AwHA0KlhN7NKA4BR0olpvmXDz/7NXQf0ONhUEOJ2Lpx0ZmW
ozaMQyJKedjEUp3QuFTpLFzp9QIvKTMrtlwNzI479/+hMvDSxYsfpAe/S58s0uWE
HYBuOgajF1kVancR+RF2plIc/Ug89aMQ0k1198BPI0yQ4SOwo4nTLrf6/unF19Dr
doRCxo06Yexr3Vs+JMCCp4JCH4KFPrecHe2WNQehLLpGIJQdevdRwRtKuvuiF12h
QFXAa1JXtt07nM4s5hb3nCNsv7VLZ76QkxbK9yVBKF1MrKI/Z9DASaccl8NfOKQL
/H9xaaNGNBxPEirn90qeRxQ8v5NahIFi2ulKg0cNscxn98777hcTcZlNPhQzbXXu
h29k+uNTt97pRfcZT1ff9VXKaSaB1XlFHMBjnQz3boh5aFj9EKLoTQ/aykmLe24e
eJqH0nnSMNU0V1w9Pu0qQSKfaZsWqYgNIwqZBdX8/jkeQmNGDfPQdaKswNW6geUa
0hFk8YXLhk2UiEqgAyRyFh0Xf/2cMLcdI1V+DXIrXnNPtzxBYCMTrktlBlTPh5Vz
yWz4jIikeiq0cdJr5SYOLjcCCS+McfMRKFEyyy4UM7Pzsts1MFQ/abbGBn9/z+w+
DgP295nRXQJFHKpqMAklNx0qs7QhrqIwmQIxnVC4aLBwoSUzLDk/IdqJCtB0ZI9B
BO2tVRKbeiMdycPWqfCje9Ekl0N0c8A3w4VKpKiBFo6BJP6khMDNAmuIo4LZvsem
AqCCnWF5kbQKIumWME2d+o3FL5AaNA7JvKHVuDAcqPGHiwcplmLjRRVaLNDu+BjY
jxt/QzqZbEQBmnzATYEgtdkiHD8zaCsi+7itJdJfzNmMkDw1iLlS5jXvtO4rKThI
cxwVQC/Gqct8l0HtIo8drrSIynDoY0T+gkSiAPFnjbIjummhJy6HzaX+amfDuwAQ
riG7qYsO6M+YxORFwdORwtF5kKFh5Q87IW/7/clap4yLAfn1uRidJTPpLeWh9rUg
EK3TyqD3iiCqhvC0gZC57kjYZEPTXLqQyYnPRhkOvC8RdPwoMzQZyNkJrRSAGnJL
ScPdTSbulyto2RC0hVOxlZmgXskYZ2FBNUT17Qotf7vwHIkpHQKD9FCU0+JsnKDz
d0omvaIq4ydgGTYyY6Bip3vTQ9Kn5cS5b/eSevI0EFxcnMcdEzZsd1DVRPv0nzCa
M+5l0i+RC5kSOa+9oQr3UCxvJzc+e35WD4Vueo8ZSgIDkED5p7SF2/GwOB60QAGG
18JOU0hgGXX8FXvZVYi6CYnHnef7yOOtkUwE4mlzhgKr77i1RBK04TkaswOekoas
BByQizXaurZKccZzCqGyM3fWuFvY/1ttYmh6B1khhsV5+fK4skU81rq5lTksSAmd
Qqa3NNiONzajm7TXDeE3JhP2sVq+RDuNETMRiwpgAkWp9xKytJgX7cjqmigIor0c
dZ1U0TzTq5N2PDq7dT4KgPVE76A/E2APT5anANYXjMaUhbzBviRMFeq3SO9lcx3J
u0Pk2zagQDyTD9al/pUPwkgSBvLjxsjzgZTLaPwdTUSIkkX99z5ZsXCP2/3xLkjK
SD0p7Mpz0HJiDMba1WAGgUfQWTeOrNKKTejRYff3tM0kkFoeP5QyrNTzOT0mFy+D
X2jx2jOm/APc/z2yYP7MhYj3a3mtw3HfMpU8BdCw1E26wKQIo3NM0D9g5e7KTxF+
WnPhr0BQf9X/CCRp8hpbxBMloCO+qT6kGDY/dplDEeroy/2h3DZWj6KobUAjjmDd
L2jBwQCmzDc/2H30IHnFIwaL6fwOZe7WujLe+BW+M1quwqzWzaicYeHLuabfd9L+
9vwRbmUTJrJWZGqHoBMRhQApJ5k0KCO0KBiFXnowVn6MJrfSCY88+tu01q3+IOGH
h2wdiJG8vEa0Q3l7IdVYANVYiGq+NLVYDs9n9xyC40syf0Ey/nR9Twrhld8prec+
6+asXLDGmcg21TgDdNjP3pCp0cf3Wzq7MMNjuaWj01Zf6XAP0jWcqQmymV6tgOaQ
+jj6mGaGrgMMXYd9vVoGCw9Revkv5lxjDdP0gDAqPpJzXY7kOkGFyd3491mq1Z0P
xGbdDU7SF1t49htmtbDrQMYjNwKhYU+EHC4BXkQLub3+gfIo5xD+yi26qt/aHc/R
mDtVW4IOnAnOcOVDs6bBJVaFRnobRMCVexqD3LePUcU+r5YFJxbWpn/1Lt8XFNpV
/8qcNWnrVmYnyQsyeX+4IV/X/sUSq779kBL2x5nbt9DhN+9HhR7z0VkwWUlqZQ5K
JfWUpTlJnejnRoFdGEInzvO/RjfndIOgx5UpqryXkVOwp0aUm9wlm1KgQUjAye+B
0On4yjOHIiOkKv9OzNcOLumOTDK98+aXow84R57kvuOwYBQavHjeAWMbFthsjGzR
9Vr8r4gLrkABp5eG6fyDg5vhEmoY+DHytkjlbcaVSFFbC03YuAXiNUYS8oXTEIol
ww2CbLpcXuyv0eHBfqKekpjm5o1MetQrrw/RYJk5ijOoJtUFbIctj5KLxGj+wchc
N/C5A9veZCNBvw1IrewIHZsixPYO6dW/XYrhAcS4LLj7K+E13V8CxocCyA3WVKD0
+VHfKC0xB7/t93/5ki96LePGkqYQgGoipTc3AEZ2xoLhBdK9D4WVx4b//MERdEyG
kFNul5sn11jYADB1EJIPfVQRDeCjm/xRAH6l+S4Xh0R9Zn0okoj3Xf1qrSziEJg/
i2DwbcYtssagdUtSlysIxEB+PQJoNvkajbhOaVvsxkViCrvOB+lcrDFoGQ1xUAB8
LqafI6N1ze1TBrp/bSiMJyws+xl+0UTVO0G5ODjpIdtbLHvimdKXnagHm5e4NQQK
sqL3ehIOFNj7qSuP3Lwnitwl8licMOK60XlR3kqO0rQ5Mq3wxKgLY9bCxAHL5xAy
uqtmH5SB6ujd1VKW9yZPlWH6BtrKXPJv/g5sxAvFABJA+hZtYzhMaqQqToeJlWOc
OFc+yUl8ueWgSLwMrbZEQhIyreKWOEwX+LTQuYEMNxut/aT83zWEq99MRIJVPEGA
cspGqjRW7CG32V206zVPR8IinHv0nW6dVFO1nntW4iOenYSjyY+ikPX854cZOWxA
7bNSQV+AF3OV44EnPc7ib++dMiKnFWTpEBjdHH+9JVAbTDTOWevO+CeCfZ2Dzvzw
ixiMbDuGdpOBFLPK1svY7r9Ro5ue6r9R4lmh+Gj6/9BVRuzgXk6IlDzZvz8IkuQ5
Qwa8JOw5p0obCOcurf3GtNS4XjJQjIhFNpBQQlSYpmJz414hxAYpWajv2BXUMxf1
0NCA51yL16t89FjqXtdEPeK88PBWPZxYCE7q+OCeCA0bhicQKy720r9mtsyq4C/S
4V4csdhZ24hKqD0N8Af1TzgG8INhUziPkx7x1/XutPI8QJvadnuBMABbgKRU1ENO
OLNp97MvzPSeYJDjUMQnq18a/ee4Gw2FbwEa8q8JQ1JcfLqmv1aRazOvlaKL8uk0
CaXMt4twWDvxZ2kPZdCAQ58aoYm2RCgzt6xL9+jioNe7A+qd6DtJfx5h69ttzdXb
K6aMjGa7UqBua0tLb8bRF4hRgGCPPloST/mtEAoZWXlwIK8otgT5ApsLR6NOiFq+
TDTHRTVzmwp6Nl8NdpXWYn+khq6loyDekl03hoEC8YwSoF1NancFSs8qG/5nv92H
WaPLrP35qQoWMDUtfFqplzxGJL8SlbpIcAw2JLYKslqPmmG8wo5538hqVz4hrv63
7OIhsSnL4U7HjAGnh/nM3dZWtw5jLCe11cXtRKKa6NuGKUw1eQDPQr1dbQMVTmNh
pZJYaoYO5cgXcb3f4pUN11aHD9inNiByKRQFK5Cw6tD8QpuWMvYX4Yk7ypc3zDe9
vUTJ4PoaZSPUZcK/wP3y9DY8kSSU0DeXR4iZZsjacUeKh5gfKFKBLPH+g6F1+wI+
ua56jksTYHxHJ3qwL/nhv4DWVUnr8cUqOBe9DxMlOd1Hg0YDb/zNfUrUFBlfE8yk
Y2d5cBOAs8xh+CzvH5nq8ot0obBzKppJPCB90KadPPTrUlNtwWC3tvI7xkD9d6Fl
ORupR61mnabisjHuGeVE+8o+qYx8erEoqJD3GF8ljyiwLvSH7MUJWn8Yr8sCL8At
z53G7KOQwSs1YwMdYI5sNQPW7JKbhmt2SBkNVyS4RoJ/SYejCuwOWsvQV6MVYtax
Sj6clv2wTLcW9gyySE2Xf5IOxjrOCFUzEOChM/BVThvIfh2Vh6u1QNXeXoGzg2p7
mJ3WbJbQWaSIFzWxdSlRX9Z3iLbOKgWBtCrx3TkTmYbUJrNngZSpSnK7Gr+MGEv+
1m3pU18Jxqai6Luyo2XzsIRvu0PX5S6B2FbDEiCTrdqwoYCl7Psf1Ede2QXaT0M5
Z1e2PxE4u77nXbv2lf1cCcR4V8Nd/tawqAmnELh+zVCh6hJsx8pRqrRfyJOHPwuL
iC8eesF2W/WVFPmeneA2WOaGheZ1rSjqcVyrtDGLsPgR0oFX0+fhdeDrO0RkuTQU
cbiZUHcF2lWkVB5NFXUfJW/0IQgMtwrcC/pgnkQJBQwlChw0g9zol2DJjppoJG5T
h3Mu1OFtE0RnYMxKRUMjxu/FW9D1Eqtd4pIH1H14kWDih+yARbo8OyupLJJg52n6
EHjYA/7IxKVqgi3ceUfkdIj+5FOzoIEg/KzY3Rcy4kaKSvEp+0QZ1yEJ5r15YXKj
Jis+e8AyOHuKyzvVEdlAaKJSWX7quXknlrYXRvpeEZhhud1ONU/b+HEagNNN+2eY
CqWLPydWSzgPK3Y1yf6W/QkSz+IOyMWuUooa2mdv6nR/wQXKDTPfYnBUG3MGUaWy
/gmu3EgVbNcBrLM29O1QgWyz47v7OK3qCoeCu4i+wg920QQ4N8FpBLiiwbgw8aFe
01CKHOD84BNMdmEZhwES4E/66wNIutzAedp8Qkpj+GFRJ9E9QuI9e648pkUrlsqB
pT3+dqWQOWd2cNhqXxrJdAYSG+AtX3KZJF30Pub3hnc0YB0obqP79JctYTNeKaEU
sYtTHDr5B8vXBSpbwO9Gw3LoSqRd08I8dTXdSSS69HKsVA1zXvPM6YFffQSKH4zg
EsUG+Hx/vbDi8hPiIjPU+Jy6SQWwJKG1mGELxUXwvSWt4t3D5WIqn0TQXBMIQttK
qQf0TqtHUTr+X7wHmUVgy5WE3xoAhNSyzy1TQULjVg/yBBGIV8FSR0/GhxISoFcG
4OpCK2sPLCDFVref9Jl2ZgTLjoaJfACL3fHLVU0+ZspCFLyxiqy6Cj6W3jyuyJ7k
QH5hchYAiukWwpVoU2a/q6v5W4GDTGWig7N/oA6BBFKuoh07NdJ6N0idFOJQoJ5a
Xhylmngjy+LyhryJNOAoIp+X1BWWYrznRi4/eVkeoeujcdjkkKHAJiVmb5q3yDTe
ja9jMPs8wMt+8BIbBpSYxO8CsYUGe/xaHBOH5wWx2GxesM92QEby8V0/kfBaOCRV
0wWOgbzp0gMqgsXb8aqJLgDI3LqMcLac4lwydopZ1oH5/KE6GLg0paInLUYrtlVc
pAnQokHa97IdP8FlDIf+yHcl4WIdGnOR6zfmA4H1Wix/sMqmtM5C+2gzcbh9HwNv
XURZ9WTYw0SXxDgl+KveHqDv5kxQUrNMktogB89MYK82EuU/GB7NnRzJ9KAjG2Fv
7hKfUE8kyK4WA7mLdkuJ8Zwfhx14aTVsa6S6Y74cUegW3YyT+9bzT6Ogb9g/jaZO
th5K8rlys5cYIvIYcJDj1L2kHXIY5U/Q2QAzEj+MykzFw4LsTdZqdduxvjneQINF
ADdClNX4578JNY0eJhfBWPzq9LroRv/GWRueII/swvi6PHcgVjyquQ/18+BGr04E
BtO7CxfY5FSNW3KaPcpIyj+0tBzfwaMM34OF0KG2armzuphU+do24Qg0SK17iecG
qTDu8cC41FncEPntCxuw7MHU/isdo2tgHxuyITQBz4Gk4VOdLr/pzi90WtDioZ33
yiooARnoidmIpKLX/Icdqup+YjIHDq5gXaHq2guMKa73X9VhffVD5VsF24btM7kk
+N5g8LQ69LI9Kv1KsPD3c8qEFuZ5zrOUOHC4idAmnq4lwTxio+zbHNyiwL/KXtHn
NriRZ4O65t3PzQAXQrdq2E1ItRvb+le85M6Ngj/OL3z4l7lTju/ngFSjMGGolGtd
XMuMjGcJDTVv91ah1fsu4vISbMKlErPesSnbNGW9NW52n+Upyl9U8B7446kK0w1g
U9Tx+/74OIp8GKCZLCFY5jACAnoiCjlF5uWJavoIIn8RuoC1b1FniAcRREe2X+7j
Kwpk8g87Wk+ftEh72rCebWLWm11rlO/p+6BZKK3jE2JHb/MYWKL8Ap8KtPzi3VTS
1/NVrs12JDFBYNZswUDfo33vE0wBChu4vy8DUEiOKesA5APeFPkvRIQZiLO//5Y9
qc2fDS3y+8XWagVgChnwUeSPkcZKOIQE74Az0lXruOaO5xzEosiic7rFjh2Wnpec
WhmA3zDzWiaKAms01gAgYJi+p2sPLuW8NVsLBR4p2EUMXyZf2lROQyX0MLw8/Tf+
6W8mlSo0jTtFbg8yI/lYikqVLmyp/PoWmxmfV8teY6GsjEO497eVBXKnSznWolXi
BmfSxK8V690MH4xP0yTvhdcmnTLfX4romQlbSD3yppK1n9Q+YOMzEGwu8edZst/6
+nSQY4XzMngl0FdP99ygk8cZqm+zKy4PnHGRuGE5nOfZR+y3ZecHVMKLZ16qhi0n
J6cYMzI0ggxh0Mvg1WG6xdJJ7IwqEMisgAhVKE81omMpPZGUSTEVSr0JcVMPNHZ7
3lQb4hfCygQDfIJZjpr1fTc+z9yK10DRpmxVYLn3ooJik0Nlze2AhHw+nwb7QrGM
ZCQ0rVo8LjET7friJt9BOiGFzg2YDE+GWb7cBmO9Qj82ZfazQl+qbkxsIQEXDbut
eaqKx2pxokh98STWZC8BeO/rL+pcFmO8YVX7DpE5dEvRqFhHFJKCxhS/z77Codb5
lPyL3Rc20zI8OkX9uInhzeGwNCGGX3cLNQGemtQdznEdm7E8S12YBL5J2RTt0Nx4
LrTajH2AJIY6LtCaGrQlZubhlo8z65AZ/uUESadaPjGb2A8IKrDhCeEvHTjbeZj2
c1wf+V0KHSIQiWn2Vdh+r78pgdQPYIzNLatdtP48Qt+SXFNbihjx6aDDiH0UEG8V
9N72dKNPSb3LQp8w4/9sR9vX+1gGh8+gP0RyojCvFlVLOudjX07rMAwMOOGs+XNJ
D1laQ3BKM6It+1S/S7U7Kp0uk+gOf4o6TXPajAlyScfuAO/K80jkNfB/y/yDDyY9
ASBGb2siXsqXFyT9q/jOt0sPSUQaDVFDWlM7rbZBkWHfeX+Fhk9YIKf47wJfTNvn
9m+fg7Z3y61T+FgYdOVmm0HxwFSqtMn4Mcs1CFArOG3zo8qz2M5ItkdZcO6g9Cdo
/RFRN8IbWfBR2KpWErAPIgAGyZnDJTeLLXlNrZ5mCrCicm6pos6g/vJeTg2c6F34
t3mqC3GZoBiUK2KctXaZjyexCrXPQ//XHSWp7b8JIZShL2n3gqwLDvxi/MwOQrKk
p78HF3JxPlIfA/PO/ePMvBhMqEF0GcJQqvfOn8yr+Mn+jLdF3dudF9XOC6mJtwcR
9tbQRJyYyf0KuWTet8aoBTNC78znqk3ZpfNsEcaOg+KRvY1o44cEv/segia3RRaQ
mkMlPIw5ooD/a+2lzns2LgEomfoQ56bGlAlCH0e7EQK6nkYzIKxbOTt2D3ZAAIVH
VhzxKiaP/cBYecUIwfzIDcrNjwhoSvi8xA5ryGW9xZ8HiDAPU+9ozocVI9gnhVJT
ZNzYX9n8xKQjpZnFAMw2l+64ZuV8b0iE9F6TvPb6n4mJZHgZi749GKaH1Eae7DZC
CuN5X5ynkQ6Ws9Gn7UoZsRVAmSZ7aqkqM0GccB1C2gFmrINJhpCBah9+CX8JY2+m
pqPgSSp8J+6InVTxN9mihEKsaOirSGXNNq6PQ80t3CYJyPyaCs4ZEAb+lrr2T3ch
4DtecOIH2OycQZEUOknvkt2uaOGCJ5tUiXSAke0tvz7Vo9AbJMadWl6LwymdAB0A
D3hOz+tFfv9LmY/Ov37zBdKS6BB17oYOM4R8nakzZZShdtvOFdx0H3QjdLcs+yea
GYwZuiMZgcHxxy8+ZEO/uN716OGjEtX5MPKEW7OG3Gf3QrpsS+7CNlCfTCkattx5
IX4A1FKP0TcP0phU/Xjm8Q1mongRzbLJL5O4BhrKNsawwiBQciYQZSUVf6rstk67
lSAWGdK12Mz+mqofAEi7MdGy9BatFW2xynCNQybOdFJ0jqdnczALSsbvCjdtoyBi
tGcphRujuupqXRH5Qd/qna78Ekk46zK+nsMyOP4di9Xy+f4J9IPKJOviaWOS+IFp
84jQbwCARY/lmhRTtqsZSPKzLkCVcSCCpyiFdA1yQ3heCVi0CS70PCe51AYuLgyn
26u4DVKuy42FdSJJ2AeQPOLYC4qNH+hjfE5MtJLh6BAUPu2OW5Y97i9r8QJqsY37
PGkB7gkW9CswLldZ2jj9E6gdqgmckili19OxQbd0CqQ5DpWxlWdznaMqavkd2FPJ
6s+nkaeQsA+vwqAOq7GwybgBD1bZlFWX19o8nwry0ddrgQ36wFmazxDEW5x7HjM8
uTLgNkNjO3fedz5lXZL8qNAMcoxvBKjoxwt8lVfvdcT6vH5YXZeN1aZTM/PkmyR6
t/KDD656i1M0et0JZthUdiPycDi06smzIfIxPZnNbjQBHdFGmymMrDRXwl5aJzIA
tCQkClTqSkn7GXPAwq10gHfVk4hK6OiAyWdRSDB7Bu6Ve0Bnxb8lxQIu+Zs9dke3
MN3MV970LajycPWRfOmHBArlX5AC0qPDBWvIAwMgWMiJQ1c+UnpS5CosU2S9sAue
DA7HqkGRlL1jMG4vhxgPXHmQrkATsPqQGaJ2oJ5Eo3v4WgUGcA66FDMHrQxwgzwg
ARon+Sjs7d+wBgdMICoYYSC5uc2xzr5w4xBtRwmvZXl2qMbW1fe92vVrm+pVYoFP
Ck6UUKXkp4rM30bobM+ClzlCQgH59STADNBQDfhTgKq5wplRA/xBb2HYHEOK8YlL
gZcmtsOotYOlJfNJr00Am2m/4mpVff2cyaE0WWYOQfUXyk6pbGhwAk8mDKOng0eS
bEXSaeRZX7FBuoxLxd9fKbm9MI60BERIDOdjvp9+pYMv0tAEl2xuLM1hMA/l/diq
km9S4U93uB/6EPeav7Z2FtjGP16bKFFWfFbLa6s7lpD8+WsjmMqCjnEEnitkA6M8
o5MLky+Lpn1UehVhTsUqEv+05NR7SP1vQcG8yb4IwQZ9jurc+Z1cTwp3W0wNdcss
ruMIUQNIDaZcKewc/8gNcNGVuihbgTyF6N65C+cZdlFGNIHoRHHyCtgVDoh9uGWk
MuuC+7VBIGjl/5Jq0pW7Pt5/6U5CS2yedhlCoeIVkVJOm1ITo7qMY3C6JmpWfuuB
j06GxDC9hKEWVN+UJsG8A28u79n8ylDU5o2IrPANzftggaIcXLAT071pmpO5UBd5
BZJBHC4Kjt1TZ+6bRQCTyTzgzHsOKsj2FAPaKB91OgGyE4ywePUrMW1YNrWTm8MM
rZkmeAEa1aWY5xrAFA+kOMRyZOkDyYxv+fATrxYoiNTWbwH8XP0LIABIIcWLfaP7
gLM2NsX5t9Ijp8lfAa+syWZ7JneLZNA7tm+Dq3QHdpgFaJX/mAb+xJ35yCW69sel
CzRAGgVUfabzFSf1cY883WhIht2UuB8jDpYV9sm0R/oa6JwU5SEyElbMQa/pmO6E
e2KTKFppFPiCRGN6IJhC3BklKkolWPgODSTOFVjvKvpM//pfyAek51NdvM6IPrDF
caJooJScZLFRJXRMKqLDlOevIuK5vYhUah4QUpwawSqTdNvw8e+lfoGKdhnRk4j/
BK00l2FvZvZ1rJUuGwXYdme7nUwS7hRtBioRGFGiwkKWkvpWw229HExAx/++Nh0g
0zqU6Tbg/9HIMdb+wpIHjoUJOiSDgn1NeyhVQJClMU0HTW46ynnU5i9hldVLzlli
mVGDQ+NQSMkNcN5Rf4Quy7KnmJva2yMNIIlrsqczl62wBgM5zVjRenSQLuf8CbFL
oPWFy4Jx9eZSNbBwX5YEyChFSS5mQp3QR8+UylowkEG/0jpBZPKWbGUZpqFBQ/fn
gli+W7NTqbk+YM4bwwP6WFx0kXuLV0cc3+RRQ7EH9KwarnOcuH2Fwjthr4CAKCi/
MLn3EMNyFY0X4n9J8Rp5+ropgpmPWPsEdljCTQvCZOjys/66mxDvi4Y8HkJBh2OK
t9krlYSllwK74Y9SubkHMfuKJJIBQV3LCgeKzzZaBzMXf6hHpJ/OyF6tWO2cQ9Yk
pIRHQB98gOIFcbyPTiNYiBJlJnZ+pt4WGOneyKW7Ao7unGbO6VJ92ZQHggRmLot1
i4w72MD0D1wqmL5dAr0X4Hile2cfTgOvRE/TLn5ejMUOGrxVzxz8rjdttM5D9/JH
ux6MD500KSVqF8d+7P7/q5u98HZ4yOtA8Uu51M3h27CWqMxIvBkmvXB7R20fOGju
fnLKgHWlKjUebGtlBJi+HITE7ImDrcdAIX+RqtUOnZ8iT5SwuTcArb91mJBjZ0XJ
mtkBDz57TwkTHwwtD327vQ7AgaA3WLpCgGBzO2dymdFDsjEdpHfqKz8CKWDJF/Ar
W2M7HkVgoDFlYEsBEUHknZZbvt8O1J50hIksrI9pF4E4wN9827MDRA1a7KzSeg7A
PtqPW9k9UCX61AiVyg6z3W0uocpItyAPqBd8TLvA3XP0TxerpfEzKtyul8TrAdYQ
S9nQFc3QGgU68YS53j4xc4nJ+//P6IPqryFOfzuq3LYcyNMt0itpRuoruieYo4xs
OYgQ5oDLprplk1sofe3/RqQqBf5DPSvrAEvGJZhulxW7IgEED9AHNectXfFyAHms
r7oHDGTxfWWoENatJtjCfYPXAIS0ueE7P1GVoUkZyOYk5hve+K3kGJFaUlQj9hGY
IPTWSoZlWtybFoLQ4ACCI/YwxRwm7zWi/tTkfvPwEoKsHUry0bIGfZ+MVf7pDoPY
bEQiCwnlw8oJ2rj2JKDXNOq/w4uygHiwsWhg9rYKy33gD5a7Ipew3NWM4Kx1mMej
yhS9R6Qd8/j1JcJWJm5sJNnj3qJz41fvMlkIY5OpT4+ptswuqA9IFqFVJ9eb8Jgv
U+vmxjrC8QqlZOp0mZJNvpXqI5oLrfitEfapRHwcvpDe9/JCMK1ec0dptQqj9aCE
/+8dNTWHsa7I6BXP10lxKFPmP/BLFvy7EPcE18Yaf/323KG3cPk1Q+pZqxMRe7h/
He/WwI5AdgrWGh1NFGP3SxXedGnwC0mVx6RK4XPraj691lrFtqlBePZhhtXgYm6d
U3zpIZV9OmbpnSfL5BX/oMXXv4sdeO1+vo24XCpLspYeeoAj65HATce8V7zd0lkq
QOHtPWbvtiWIQBJO9buYS4mjOLsxZiQqCz3eOM5QgHrwa7OxNYNKvuDKbZIjqy14
iDSapNwZOGyG68DVWZzwSlBHypAwpCiToFKo/D+f82+n0aNec3COAMFXN7EFC6CE
P0g8OjO+Bm+sIRQq8JDDjYwce2jdhuGec+pMohi0EGq1btT1ikUKpmb/sjMNy9sL
hc6+S/Yq49daB0lQpAl8DOmSplTbEyKzlzC1Akj6aOt0KoXml26oZkuURA62JR8Y
aGFo7LTZnJBKHNk8gsOs8pRNoAiAUap0GuKx5tVxzaafbnRe4CO6tMJIQeahPavY
wv6DC19y9ssrV0aXZBTI+45uhX/WssIxzfxI/EQb84wdao7ZtpZBAvhfWIUmo8EK
TA/VSebZVFH2VYi7pGzlDeHsFuecp66F51SkHXmwt16rVGtRrXSM7iVJITky1jJ1
OqyHNLicAxK3iyrWf/TQ11Ro39dTvlB5z9d22rGOcJVqyATcAk+GaPL1w9BO0wD3
hpq5kDp4vBQEJl7BJjSdxR7qpV5BT9ULDwyeTn28lIVUAKKfzWd7q4s8L466IziD
7sBG61ttvxAiMXcmNaQsUbobiy4Qv2yc8nCUrEeqq600bsDvdbUIW13iOgPCtHPh
mj5CzvPXJ4qw6o/AJJL5+6wOQiiM+mv/YpXw7I6wdhreSfMImmh7i3E+1Hlu5hni
2L7hVBBctWtR90ZR6Ue5rPAVc4ZTb6J+y9m0HqadMLs1N1EhhoBjF9GDPs1Be50A
u0axS4MfXNwVbJe42/6ocM69TA5HsLnOWBkXIYzxki+caqYEoXmtDzSbR6dVFe/y
maf7kPe+Dqxv0LJYihfjaNhhvmwjgk61eITa1IZRNvq+tiFVajr01ok8A2TQIXk4
M5JJqDxpFWT7IMLagfcPDt+1iwIjLAdqfAqg/wbly/y+JV0IWIpK//EZy18/zVCt
IojMkcsc2qQHHEPou5NWAtMABG+mBw9pv6WRjNdTyHJTXzV+5JUZTJtQ0x7ectgJ
cKkfvzpjPlQO3mLS7A02bBySCSBuIA6MsCsM8IlXWtfwBiOc6YmXyRuyYX8T9yVe
Lr6S/BOnTaLjG8XWda5R+ow/rp05uVv1KrSQHvTR9hrAH3WFSkQQjVoTDxb6b29f
l+moiGzVaiJWEJwGpj+XV4HTG2UbRksrN+IfxngjGmyKzaMdTk0JBpX1LaWOJUSU
7W2IhBBYPsqnc3tyM+GYq2aoqRshJZgQPRGEvw9lwc5P+CT0AYaSk1Rt7CuS/S3T
y2bdV83hGZgqrTR2v1Ci8IJWjDTS9e2b7jNPhTJ2+qd5mOsPRPd+3qQrV05V0i5R
EB12MIjwQLtFmLXUgUsvoN7D5faWD7Hx3lCBq06s8tuuCyNi7MzyGkwE64luUh5W
A4ZfMck8BCKDZ9y5SZK/Hf/fvFjjwRdVX18SkTcFKmPDaeC8aka8fwNn9tDsoW+Q
dD1dJ9wt4KY92mGznC5jYrHxG8dLk/hde/UA3CuhXhh5rmIDRMG91FHsrnYLkli+
ufax4XzKwZ02PAa4P1yq7+WMPDaM1J5D5TWhjUpsuiBHvnHIXZGM8Q5s4YKI5V5s
TMQ9Gcb7xOSvc1RqQAM8+n9P6DNqcuUvHZxRMAn5/BM9I7a33cj5GIl3asYxVisw
hjlNk8iYKvFu/1093pg3OSA59/cLChsgDyVcv2FbeAjwP7u0uxhRehABzKkENtz2
b+9D2h0nwhbgFvcl6lOIdKUVdG6gzoWqitPsdo27jnLFIFyk0al6qE0HDMpMCmM8
XSTNJkywNyFjPiAsP5y99keXMkO2Hijaa0++eVspGmV5oyW0OaQDRo3yrkQzM7pm
aAeTAEmJx4ZILp68N/YRjDczE8oHTabi1ij6aLsA++4N7xpUWInQaRQtaZj0yZTu
d+6SiieI5IK9FxIhqUpX9OkbFnFowt0BYoY6eb9puNOQaEjFsUL9cM3OItawPeT8
0xj61kV9kNLyLoaG20bUms8d7AxtX5aJJXyh0WZdaqbPDikUwGTM4w+dZLy35gZP
oa5nyiHVYBHgDHQnO2dZlxl6EDafBaVZ41ShB/3WKDCVJ4RxieWUKp10X7lbWLdY
0BsSmgygsgbNYn8CY7sxS22DkcEDfqaoaiW0+xe/wBep8YZKq9PIjwRl42kmMMAw
Q1jLWQaagTb5ck8LKJQN8gNS64/Fkh42gy0QQgIrQL1TR3w/k3+iWOSsBayEWaJ9
WPD+g+EOVKdK31NUhdFBF76ViU6s5jgyAf9PfBuzc4gwkg8PHaSFHgRFLJQoh2iU
O+rsDdYzKxwOqoOzcfCX1IQuhm6tnrGTVbnv3d7+DQCFaAS6SDAot8KCi49E0Bfm
JgGCLcV5hDi3AMNoXToijSEUq45T35SZG2JTj5TxzuYZnof4MTI4EFw71v5jH9DB
eWPHfQkHYTLq9OPm8Yhl8KKCZVjs3jTFMaZzF0li8LAmqj8bFHbBKZ0D8CUOYHjS
mXN1JU9YWc6moJHp40NyebAxPEyIPrg8b5cjuoT0U5C/JCcat09lmT8Tgm9n4Snv
bNYMFAt044DPG9QwadN5TF86E5XwxPiBpXbXoY+QfymchlSh4ffNxHMY69ApWWXi
1kqoEBh81iqeOAf9ibV9K6JSkzOcyswHle+TR4ul0txpph/Oxx4btbWClEvk/Ark
VuWAJBty+g7F+lUWO9CVGPv/AzFxh2hJ9L/cOXT6MNKKQFj/ndbf3QTUH2OQQf4j
84Yq5WgLAmoi1gqEpRBs+AWpNrOPI3lKs/+lSGNoF3pz9YROBy4LA9OfMtIH4NdL
NWP7ieqKxW4Y7Y+GkqbbioRowDrK4GcVQsz1WxGQjOAs6pCdbrquqwHENuUhBnzW
9pE21nojiykoF5JQSswo7suPvgn/UmcYZaKdWwL79lLHaavgDK7w/cFb3UmGvb0i
Yc3ipnwcC0JSiTErZZgABvD2TkxodGu4bEMKVKu0bmmDHSSfs1dw5oQzT0KKwQKa
no8oijNdIVanw9aB59ciW/IVLrS6NO24uM8Ae6uj4rprZZDHIB+YsEsC7Dfo3jDW
ZueYxojDEJR70RTnM+bzdiOalHZncCyt7ikPme2njean7GBEcpoeZ8wNZhVJLa20
CPQz8Ha5zrJFTteXfIIGyFFMxn7s1dH6UNszt4Z9M+b8X9urKl22c8gtARbGygyq
YKhVb0gfYnl1K/IFvGEmWoiO1xjZs0TUOMmmKeQ9EwlK1T3VvdklLj7J7yfKLW10
z8cn6s+FS/eOFcVvHJKJxsKcHGeHsunAIujdGbxalhBBMuT+b+6nsokvbpdq85qH
7zq/lzrtRhmcNohqg6e5jZXOxE4B+/adtKSabVELLl7099J2j2oJT21d77H9+KaM
AUcFUofFgouAcfGh4W7a8XKMBwzqjwYRQpdTvTRnrYsxIWot2N6+4Gfy1E7Gqco8
qlZJr8r+z33M5/yQ2YZ8X0lTtuPqE0XBa3QdWXROo7pgs3/9fkGAB2KIrXBMIsfW
1XOdmcakVanUU9wZzoeG1xWgb3aMxsWyda44brVP864qjTvoxGXNQK7UZ0/90Ra2
OvYVfp3xMobVT+LJYa/c8CtaSf3jgLHcgs+FwGmhD8QKnk6vVUtygyDpVVusrUAW
5JOPCaodwUwo6owqcLarKwTiQR01rJkl+w5M9XTDepQKB8Pw2b68Bn6QJBRo7Qov
IzP/NM8fwzQ+mpED2ptt2k7OKx3z4//IcftMevG4gVqh4YTY4S1RD/WGwx2/b7pO
rccMzGYkB/MbdFeKyZ7h7OIULtfCzivJ6eel/LcD8owoXiqXwr3cIfUHwmnFPrYu
VzFN9H4cQhuJ6U5ydsuOwSOo80tSHjB6RY2O1d1mM8hYABeBO53+GKJuf/mVQzyd
F0/v1cp+9luvIkDCm1dgyGRdyrn6zZrZZPlZhmrXxMfgPzPW7NBIV9tBKXqqeWHU
ETzPDcEZATb6bz3LLWQID08RHG5I0g96IK8z9ZOaBlEMzP1Hbm63v1lHGGfh5Ir1
ZkxE58mpFZ1w3QZOjXsmSXRavnh0wnnBm3e81hasmSfR2bixlBYBUqJubx9Utlf6
pRQ4VGpZcOMAELG5MNXWK1+3w32iuvgHjvsM1O0yjhiqQ18GTaHBhnzQ7b+VSV/7
RCHVAnSlewVwNsKr0mn2LZ/nLVg71M7wZdHmm9u+JrO3VOumaH0jenTUWCeaLM+k
Kftnd/PlWdsdJ25iO3YkHs+FW2OU0adXCQrvPEiO7ZZBdFEVqke7jFlbfyeNGzwC
mNFMbOWBs17A/0fd+XYd0GMCDHdMiKw+TRYGtbwJPHA6/HADnBdYCyoWmLdgQ1gB
+PWhu6VQc++9BX/crYDJ9RWQsrTUgwDsT2kPA/BzaG1s26IcZQoYrOeQQyNkP2r8
F+ghVVk/jsUzT1ocGYLsbJPqzOOjSQc3tRhMQWrwEXVJiPkxkUhaSzANm76Hz809
NEsFgFDPSfvx66Fyk+kFDrtjjw3GV0+i6IYZGDjdjyeSyZU8RQHioOvjZkvz9OtQ
0CZBBbuaFvrP+VGuW8010Cshc1yvn7hCKOaTT4P19dKaDfHmjR7+OzKKpsdlxt1d
kXvgHs2SMT94/xXfthHdsXCEUj9PzWfp5TtlW7tszAAGGpMgtCJ3WGk+ts8hZo7I
9WoKKWiWJs8Szz22faDXx+S8SN/BQnfXHkGwlb20Ij0NL1lUs7O1cYQ6vcmJRYdE
25h2N1O8Xym2qX8LuleDhG6o753k1lSKnACxnjfAOjjwTVBbgTaJNS4b01OWzyc6
xlKipdoI9J2K0Ce0ueeXCuNFy3Svl7/s54jUzW7L/30yfxbTHkwTZPC0R7Mt5eJK
DwRYW6JVbogpRB6HD2t77AfACxWVT2WgpiXDP7bwmbrWtfmEvZU9m4YAZAZAKieM
j914P0CxyKc/5C4xmKFkoPfXaNmYTfz0X8IUce4m+EirV33oG+rlwcX79RcbpKak
RSHuFgVdo2wEP6rJxGbc3XIzxyodLXPKuOxl6Jlcr3lVwi0lQwJApWbvJQS+7jXW
QEukc2T76IlERrw8meojadthSnU14TRZyNMrqkkTIulxoIJ1pbyOAufbv9g4tDT6
05J0XbGeXIrO1CuMfZqycosKEsDXAznCOigW6YWaiW4I3eTeTk79igAupF+GNmp5
i2YKJbr2+jBHyqMbog30/OKwJok0TqHMhH/dmlvlLI5yKA6dndgbIxqTidEAm83V
0I4T1+bEyVuvRaINCC7uSRWGKtSAFeOgZAOsCYC9GsImy+b6UbvgPonbNNfDPHt3
JDZrAQtiD8iSh28zZ5eYLXP0FjxHV0NGLLXJ63r5yDqfOIlSE90leqCVwoY+z+Wg
1ZEgFnIk4eTtAjPjwHbPyWhONNHTqOhiP/pfvt7AopPOyPpXpyQbZZBvsBz6rmfz
TKl+ZVYPNwhpnANuz38ToZkf1zovJRtdDNk0M2EKLQZMwAe3MJ6z/P1r8g118SIu
dlCPFdsFQleLl1hEkBy/A38C2NgRZ/LigzgwDQqsb4C8tVXroIIfIrjje90n1tGT
Z+zO4+IZTiQXNLOSb76UZPplFZxh7LvRqeFmEegCvtTku7/17QjWL43eFNq2F2ND
YfkzQYfz8yEj0ruZ1lC50DREHtQr9DkRVYDzuHvhWYyTcoKXi4LS6UNNLi2MYFB9
ztHm1TkjMGEbqCn4oTFfwJnMOuAO/2vCHfsfsx3wvfXVOyjBP6FnYHszfezha+aW
F/0vrQJ41IPzhxUvytB5I3MucQYGz+N4wdMmu6JrOd6gMGQ7JPy9kaKjhIDyUOKi
9Ob0lQmH3lDfZ45oBMCGJ3OZ6fkXm9+nlfxyWNbRe1yk3mF9kciMd465/cQhttYw
MZ430toEG/he46XFc+RWutq/Jr8tPJ5xTXdouiD1ngDU86YzY9+US+ILkPO2Dgae
NFAZHsKSYzZ3eC5P5ctXAqeli8UXJZWKYrmdmwrsoe6l4b70LSUz20Tcb4PlcxvF
71p7GRCzDheUSNTUJNeBi2YaP1m66J4xTHYZdTCgF356DezcITegXK8paLCfbAuz
G0E2cef7aTPVA8mIWtnDG0uMVTHFKfOCyOIKikMigvtAmLyZYBJH2/4xebYMwQYb
l167dW7nDK4K4kRhA9L/7ZoNwac42e9ha6rF6wyt6CRffYTKGeYg3/cu2zQ24lDD
U21dGF8O8o/Inb8RriZKkToQa0L6WXvALBrgcka7tv+Rx+q92sdWi39T7H6xTpyK
nzn+jKWUYZOpXetiCydvz+28KU4EmohYhD3oqynjp0BR91PzpHFkbvceXGb/1MDF
P1AHrBxbLeJmneVHuXqiU8Kbnpu7IOE89USE7wM11+GGCcTDNTCWAZudKfgCdKwH
HhUUJBZrl1HmKzgmThRA1flRl/0/nxwltAucp29A1+IdNbrMb9D+D7XNlzIhytDA
vCuok1kyRPxBm6i1BkVCTxkrL4m217dcT69rkNi4tpfvDbLGEaBiZbtid69mvBwy
TuyOxSp8/Q7jg16n/bX1dk2NpgTCoYnYPz+FP+4u5JvGThAyLgzoDxeKpNZxVLyf
X9HSnjUw2VLoHTXVfsZap7liUmhnJg67XlM506COpFSbbs67LSXk75bPdI/rSVdt
zPWXelshNX69emLsKFxaIWaAMMFcbnOn7LQiygt0MsggfJ75dP5+jWuJAKxekEJC
Y2gIw2nCoaMci8jtIUWh0MbI1v0MKmoD5DlrIBv25TJoM6di7kD4OJ5/zDiz8YPp
pUytFaqLnNkZNr91zamFqRRDO4u2UUV8/k2/oocPzXMU4ywqQOvyzc8yNS4ZRdvL
lE0gwY5BBptkD3Zc2srS2lAC31eQ8qWJe58oLbPcRPpK9NWH0D2ylJFd1XYAANGD
knHhVwYCT0FvdUaIKUglK538jBhGDpRx3T2KFFw90XrvG4UdOcq/gfO1qZazk40B
hCkNkU2Lyg+93Tu1g69X82PHJttrS05yo0XH2MsWCtnMww8NLklZExeTRjqfqz5e
+tmFZwBsF+dZXhMbFa0froO8uDOjS+vTb1sQ5CDzcYovIdNgsVz9t9A1no4gIkHc
rH55w3E/d9Hy2JRjgfTSxU7//UcVOi8HEqSXYH7Qwn44m9qSiTRJOi6pwF5SzWhX
cDNgMOM5o7pi6U02OYwio2VEKFEN02cbLvaCTjvEHKQU1Cn4qMTgAjSaA6oMwiYe
t54+W9DYMH0WChPkN8IOMLOsKzLS8teLr8SaAcc4gwOf7g0Tcu1yRrZMEC/JspiH
0rrMz9cOIzybY/rX1lML0JCLw5K03RSSPG1GtplPgTLV5rY2cN2V+1O2U5KILJFe
eLbMchrG71PSiCcqdHFhDPmF52YvlEgbftE9zLYGLpzA7HjBHSwDU7W0PbXfcWAc
+ahIxRAgEFCBmfghI/h8AJeALda1W5/8K9ocH6cgYsPOf5lV9869Y7CWZ6YE9WTs
O52H67WIMrzVSAhMmjHVAteBAwaMFu560mtXmrZjGKQy63jRGsW5pgCyMunB3Gpt
013oluxv2fnhuOCio74H9s3PqisALIbAbgKkR9RAbr2lZ0Rxz2oQ30sUAeSK6KUh
O28mPwzWWCMnSifM1cebYE0SJL1jT2UrxIbKpa1NnFW7jafS7YpCbyQtrXSA9PRC
pBirZ6rMDN4bnPG1NsI/+x2OCMxdHxexDk+LcHBy17Md/5U2TRaq6tGX+G+Ev3Zd
uNVO0Z7l+UwLhRZKSKs4Q26d3SmJVkGrJtcgpQXdcwHBfP8sCrA7oBq9v4yC5Z0O
tt2bEgFR2A75S4svBOamiNWmYyz5YYiDIydYwNf+8yE+MIeWZExanwqXc4qtqZ9l
oOX3jxaMC7OfM0zo9uHtyvWSkVhTRv0k2eb4AqViqd1mKlGW22yWFRC74OzMLKg3
I30eQ/w+SK3yHN7Iydg55L8Z+dFAkf562mNRqKxenrIleeM8cxW4KH+eqe8xCdXN
QQsKawuHpxHO2qUUa7TQdnkGmG9mSYLWXdriaDaWPJeI+2ODkGd4+ciLCEHekLhE
0UztgQM/fkLfotTWiprpv5SU4Th1OBdTtq+MA53VYvwB3YzKrOvb0u5FPsK240o+
PcbUJ5gTLtWSJmTZPgfNrWf2elzvYtLxel09ut3dUf6illx9j7s9bqOPTko/UyCF
xk6Bcx3MmSimRjvns1ahaLpAc3hdcX7cYXiHZFxNN9EsRWNOSrUAoLEpzxoRsg9J
ucEatydB5kE/X8ZpPzQwCws84BV3stysanInB3QZC26ZVvVlo947M0MHJ2o4j6la
a+PcvzoQOGgj5Cw9UvUuyAiIz+XDx1bLbkq9TL2/WJ1EdftEKGzlpJSYfBQZs+KB
fxdthvSUlXyi/DL1+eBwnoQHSw6ccxHaag2HkoPOkz4eWjh49y2nz3oG+/K0tRrn
BFqYozsQKFarZ2p4+dOuLsauWYkTkBncWPxXvC6WpWU7qVLt4jDyOfu031BDmlbl
Yzj9mJpgADhXMvyo69qPNpH0wRPv5Hg+KSLobnYstW83CC3UuZshbGd9g7nilWmV
Io2EGHMc9TbSV1EC+6PV1MDj06+Dvkgi3fO97jupPtRpYQoKjG3WyZZ+RHFmbBuF
FBaaU7jkVWF+GhqqujAMKg1nsDUBGN6xUkk8Xz5eBrPjnjFDU02AIrjwoP1hcYNI
i9tSuRuHB/G2YlTy/gGNBger88VTYwCL8mgme5nO6KaufT4E2bPcTe1+FUWNh6jD
O20nVsv5a19kruGIOCSvlZT3MFo9zkzSEOoXtnEx5vuI9fMdwDNk5BAq2Ddt6lzg
bX9qxpUfGimxQprWSpnnrKHjlLDnU+p51OQND9Z8NupdylLfrjZmPhsVO63dPw1v
gxBjYIXAL1c7hz5fMNvsixj902UIxwBJ44Jl0roY1dmO+31xV4pkEy08t63cHtON
zaAcnSpBMMu3X9z6zrfq+0iCS96GShM10CEwoxc4bojLJO1hLqH7wazD9yh2x+Uj
MOX7JlzRznmGTKUIxzZy1DrD2xJiuF3IyQkYUNcG5fUx30SbiOEfgr99JeouITy8
wOIkWGF9FGFPmsczRmu0uQ0RkLwHVMGJqThW73nmG/WLOYiB+hj0A62ql2o2u1F2
6JaFlcNNWg5hvHJs9E07qPXZSAEmV0VDDFxXsDXZ4Fqs0TUh1z0rkeU+2nKZGzIw
ZnVuxb+5S58aCrx1nNXutiGcpi7WKd9DzNfrjSxK1c7POli2Krgx+NCW6UEcBPhl
BrK2fZ7sIoJJgFrzGSFgxxU3YJ8qv3hak21COndzr3yq+w306hZO9GLdZoGzyT6J
HfaTNBd6mTHp2/7pc9DfAVFpHcAhtkx0CwepGKOEi53A7CXbG3d2HVMkhFoCIw4z
BXXmm/8qdPNkYZx4ONysj5ezvIazLuxvj2fTSuzxqPlofy06LUBcZYhN40piX2YM
a3EngHCu1ZSF+Ml4A04Dqct1ub5jfK/8ZkzrW2NMN2R9J571msCdEDBPAJiVi64x
36XWStokn/LrDv4zz3RNbrM1vx7Lgf0KdcWuufZ5Qlc+JwFPAMBhBI4Wb6nli/Dv
biW5v1mNjYjoIlZkCCagRF8Nn04zYW/fZ4I2MxRG4osacyaL74F6WLY54PLbbNcr
vAgML4mDjVCvtPQ6aNlOesF+hQiQEyYcWv64ZmcwLq+TatMegKKyGPC8u/4iZOm4
gywdtyQePBOvRMqkTELCxui4cJ9Uehje7snULX9NUAhjJssxKj3OTJPrgR3OWKIg
nuYdWnjkhDXaj3y7+PqJ2aLOj6GJ0rYVP+pqhCIAGzc1GhOMhS7WYZP4kXpD9fgk
xZUK1Ook77SExwNppBAglqEJjysX4Ld5ccfPdTwUhVd/4HGPNdmW1c1trjh+3Xec
1OMDuOvu8S8OocU/jobXgJx2+0jpU6eQmX9erBCiXrG7bzxAdFYTMVxcAZGhTJmh
rdGvhJ2XeGNFxdAWbqtlfaXRKu4bBq4JBN+NMHTWVN9+RAlGRILoBjb8uiktnZXa
2598G0Xzi1i5SOxMmbFHB1Wrj3Z+W9yM7iH1UryW74tmaMbWyQAcHbGfh5EcDyD0
t7AJ77tnWxLxxa8QkktOCq+SZvHpKOKWwb6WrKGWNgDQBWKfyyCDp+7PpEXwwYD4
nC9LD9nhT+eQ4SHiCls4nVIUg9xzWY6lXi8TdqxXtfdk23B9C5lGgkdJHZAo67MM
Cepo0c/NOWGzENY56SvdK/KGaHRfsRmrE4SbAGKC6158la5yxfZrXTComTLdy+hg
bJpiM5LQqAlU9f5sgHQh+7Jh/H1C1FJYmoCBki0SLE215CPormWeTOD5ubgOm1Kk
O3q+4PixcyTtOjZ9bIC/xjzs/KWip7TcflUMKpy5a/l25169gqfHzfJ74zbUFoaL
yD+8AruJ3GeZ11LMG9dBQyYIfIxPjVgRsCGGVHPhlaeRqTEVzq8Kct1o5sfLKmAF
MgdqprSBMZxstiK85gEcyG09ch+4i1Ry7J6aelxdWnvae48+Og60ohAnuT1x8cjl
gGA905W394LbgPlTy1D2Dk+QIBBWKr5SUkLyXluGxX+u56VcIJ3x5CytP0ZLesAO
W9Hgboq9qMY5RSG6Ma3jItQvTmlXs1XbvgEhMKUr5BVw2AmtRKV3ICkaYdQaAHa9
Wn30ep93c6P3BOoj1B5bTwfMAi5aPtsKdBDgiFnjC+RcVj5yndXH+lda0iRhWfsm
MR2mE1JQDMZQh4+5AzdnAwjsLshPgFwrLshPtidN6czA9L4rGA5n03hyJwOktWj6
KUxj1LwZ8szaKhHx8dZ9QP8316eF7JiijZb+Joco1qGXYFv+aBE1aEZs4RCnH6nQ
00Jwka1ovJr9D3Z8gunmLTTKyRmCDvCX0zvSrolikQzmOzJM2JMybd32hGZ4J8TF
5ah/jQk6CVHBbUP9pj3w4nHnLaL+ml/ICDd+EnGLi4xyXpYCc1M/F0HfxK/o7d1j
eHuVy7EemYgwc+ychIcNS0Jb/iSNbaxvOH65fJUgiRbxpcnvi9UAJPwXZqSh1QKX
5CIl33OdQualgblY6AbUtBgAN/EGGc9PjKcqb4fdv9UO/BO+k/7hacSrf4XY6obw
OT3jwqIlp+zZz1ZSaEub5wy3BikyvQITmghrpzcH7zFBHrfT9nrovdI7JedRNTvJ
Kv5iR6M9RPey06k3cVU/ZdFaZ+R/6vNqEKWVSHSN4D372MH9hm58CdakBLOM2c7F
n5M+F7qP7saOQvSAv5/TofsUvbpYP1/qFlmOt3xQ6VIbnIn6PvKCTDRunh9bS7Tn
NUa7g1xxYEJLEcUWzQwlPyb2swFAb3cDqD4sBOQssQlNc07YOXZZgsLZNtBJZxw+
VmarmzksEbAM48meJV5iLjq63N6U/ohEsdW+xxqPrbIOqr2WvAeVCL01UiXM1f2C
iaGOkXxE0G4amQ+dW8Hhq4vQ3NI3gyHt5ILMqFf0klwgGza3MnAkpCsXsdyNbxM6
zuslCvg1WTvY4c8/S1KsiPqseXVdaX349pdX9+fLvLNwV+ONoFV8B0XLystr6WwJ
ySgmlsq5Hmud7/t3V6mWZ+ViuEFomR4DjZtVmDhIeYIqKAX2o2RQ+/9c6HAL5tIF
YwYLbwWLJm52oyWqig/gwo9dLUab4SF8/R+cdkpq74IPrT+Meq+J1NtqHMUDjFmg
P2wUDUf9bO0QHr9JULqf5F8hY9eN6FSIUkNBba+Iw0tJEA2y6Gyjlf9Zkx9m5GSq
bTs1nLFmVrG7iLus3CNlnuEDQubie0mM1lfIp9WFGSLhphQIxqMfcQhyVf2r/Wyp
DgmYR/DGliykA7UwS5AOy2+GP38KWX49372vMqXgdQxrFxVc9eKoU2oaf/h6yH8h
TYI3t0M0SUMSYy2G3YZMd5mE9V+WLdBXA2y54TWm8vz4vt5fZk+tYYs/fS9LMAAp
AGpArYWiQgtupmR7PyPp352OWhqNWumJQWJYtGwIJHaetr0oZheyw6MKSLHsabKI
+5MygfKsIagTlJoltLgYgVzfGsnCctq+iofzOdnLF6yXdnpanWseglh+9DWrplq6
bXyzv9qEkgz93+A8c6WxEHLr3jv6koyEyuV7jv1x7bgp10v7ZsiFsMlflw74a0g+
FjCjq+vIiIVUjCYO52UUSAieNc4FMPJfusKE2wdjVdAB79/6PTulqYuXful6tjvT
LOwNPInto62orcFDAnl6Y3nzBe8DRg0V2BJILAuyh1AjV6ru8o4kTNpgbVaTeUyv
hsyDImhrCygIBM5VsZkuLukZmlmp25UpkPdCFkzm7KDbzKiG192JyZBzzlKsZOuo
OwAgwt1esoKZw8irmR8ssHqRNDcA5lXHRavRUn2ERo2yK557nf0xqrC7FrbYQC0O
LAWToaklmeQdKDs+Z2h1XNAdjRn1fmzjx6sLTqcGCqzsYoPIJNwd6f61J63FTic1
ahY8Kgan1xL1rZwOSc3oV6iDVvF3IS63cL4hsSN9TfbJk9bn1C9fS6hzq8ea0g8I
ZFx7hrVpZ1EwVIrEpEA0jh1SsfH9kagtP36vlsfCCiq2FAVBVK9084deeYp84o5A
ueE3oWEnvhhJa2naNRRcoAyddPQTjWsI7IDoct39ZjAPVsEGT4/CaJoxg7uPqrHi
SCRzebzaJEZ6CLyBqAENoVniRixaK05d1eC+cJC72/SRsJeze+7ItYMM0PSLvkd+
jgVigvViVTOv4tCrjOqoEFnJ8glupRPfp101++a7ZEDvUEMMndBO220oe47MW6hf
OC1RBtKB+jSLgzf6BUP9BSM9tqfEW35m6N37Sa+i2SqliXOQuVaeXiJnGnXQEiRD
FvFPeXkkGP2JQULnYUK6YJrxYrG3UAndNt4Jj/pbZ+hmaLVUYldJ/GEzAjt94MNN
AckWUFVUM4UuhF7XnbmShLUzsKpjSG4ciwy1P+AxjpVqxIlgRQcqFwSdgzrmG2PD
KeVnr5R02s+CU2AVZjnI3qhnw23oCCVkGkdzz9bP0+Gg29b8L0L1v+38xVgg/LTH
IEl+UQV67jlnYcqj7zElutGuI1ewOLfgIlpqhUT6STG4sNe4JLQlnTfCbSm0eLAn
I2yeLQCrcOxOm7xlMiXMGAv/+uVDtopbqi1QWe9khUbreVayrwFinnNS/Ml+lI1m
RlyafEKVtOm6CI4McjVd7siAeVTCBha9P9ZCmSxR0LRQAkG98jcP5jFdVXMrgB5p
ofyku1YGfEOUhhcw9vG8c17dUb9xlRXJdnYVAt8C2LdPTPWtUsi3r+BVDfLShLXv
MXNBrBA5UXl32Mq1QF5YhQ6+baDaLdqSinOzd5JjJsI9+ph+mrdDQ+U3fxtMrXjq
IVX8FjIDVu5CCOSidp7ajrFI3rtoZL6gh2Bo6CJhjD/I89lv5yU7rEighsZnSBgc
ErV0y0LMhrf+GOdO9onM8XwZjvsO63nkjEveTIxEn9MGluzE/G8xRPQ/91oDqDuu
3QuoDseSe3azozEkiQAkHb/fzLAM5IiHnUYM4mb4Mz5gAs2CdWXQiRBKfdZKxQ/4
lhe9Fa/AlAZRAdsdg6f07z1tn1Weccdz5HuxfWVtcA0ZIkpJuoRAEikUWGXY5yIj
G7y115rqeVwZSTmP/TQ1aE/azLrab7L30Rf3+YAHCZY5zgpxyD2OvveCxZ3XXj+J
xCzIZSjJlNLgRr1jxi1autHHjYnF1KOHnv+RoNzSVdZe9SV49CtqgxcN2VDz12UX
ae9ljqqruWC+F6JQvFm04Bpdy/IfDdChtt0az+btvxE8Sa0Hg8eO2eBn/xynOS4z
/MSiLCYGQlT+ZCCAI3vKvzzxq2zI0InYEK6Yg+AXULO+7msASfP26EVTO0pfQiGe
/rF3SJ91Nbb4gPkZySv3MsrTEgWeo2Zcu9rLQnJjNsf5QKhoQV1GhWm5toOhVkJR
8XXrLLDT8IKv3iz5XWngodIRKxJdi1j7CI7OgK4YWW4km+qYWcxFfIzZB/IMd2rL
yp7fysUhV0vNyrL/czmYdF89qJLKrbMDdZCaHyattBn/lOYMUstE0DX3CjTOQKns
juPvKevAD8LaMQo5iNvLw3JxO3BpuYGsbfIzjmSWfD2WYeXBjM10wf5KoTCpDuGB
PjkXsvibzmtmE5gOJZdZ62EioomNhS1lfjO4H2F4IF8xdd8tH/OlDfmm8xdaaxf9
r9t1QpVaMHQ9ZC2ho5jU//bf0y+FXpDzhBWg7Ff2bD73Dis+uDau1UEJ32Z1UESr
2Rw55Wa56G8c2Q54KrotrIKq2eRNhSVnI2eBVdI8dPHr6KWIdfz+WPm/zKjjNR6O
BW0AOPSW6QXb9GaRD3NeHMAXp8RZDoMHy1233FNiA8hQuicwblNK0eQLWR+1YaCu
2Jnia3sfj7YNSA10N0caoMM+NMLOvuYhA6pH05hM/z42H2JSCGSnumXWHkVCq4m+
rLzvirIaYKrrhaRB8CfnsRLWT05qe77WsgeL7DuBhnWval9x9zypzH4K0nw3Akyx
qMQx05xQsxkMy6/33o1TGmK3TdGVhbowi2/sl1Qc7jmHKgujf4ZEaFC6+fdd7f2l
I8cwxUmLFqsh6h2yZECQqPPo+KtrOBPnU2LwbUyxtrPaDO0LaooJc1A0QAFnvlvA
bQZcZuGKsskdbd9bisPjd8i5XJkL7WXpOKwKxTvK8p7468IGZqNfjI4MHLFXD6cn
ji8gKCWGKuIvDYdzc/hG94o5ZDnPaCKe2z7J9vrL8XeXAE+nF0z0Y9i3SN38aKXd
mLfr5IQTV1qYbaMQqKk8GgvBZ91mEA+NKSYhxAed1/8+tWL32WnrhJYA8IzwYicO
DUU6aB/zjThpzlD5QjIV1arY3HXwON7frpLplUGzwtT8kkEjw6FybbNmoHrzMIRW
vrwDnbHiBhV1j18zJkDAmlES9jaBzhudqKjQG6/qzGgg+2ZfGogiO5Bg9bHsckPG
vrnU7nLM9QcIynpsRHF0eurrgzApsdkOHlPJMd1kDugYZH3ElUI80rcOtmZHkkm5
yZ3AIPt6D0+M+HTcjpaidL6uu2uJtiXcSl7MhInQuAyIt0ZzNjm/EL2zjoDeFAqo
n80u+z4jIJyLC0fpxwJ4ObA9u6JVgw4TbVMiZaNac9gfcP1b2nPzKdJeAJvHC3eE
Wb0UjHvB9zw0o6J4uGa8si0HlSLF160QHToas3PfOPuciJ0Fc975KSJLPICGjjCo
THiBeV5ILbrvj3l9c8FGjUO841AEWKLERL3WuAbM1LFp0GlGbUVtsKgErXupSdR6
z5jCe48VV5bJpFEFlTWp73Cdv7gOIlAmJbUICyUXaePyXfwDucIRW9AoXlfVK+lw
/5FvhkoHNWd8URqsc5TguMKycOaW/z7F6WOxEQMcbDeM3YFHJXSpVtRndKnI4pS2
CvHU7KiCu+zbIQmVb1vHkDx9Eyb43Ht477Od+7R+QoxDciY3CskjDzIEu8LFAJnb
IptK9YLhtrA8bla2GaeYnbcUbW2wP196gGhQXhoRwx0WP/TUqmXRCIA+6NKiNqtX
PXov90wmEh0Ef31KkvuWjVptBC6KzZ1zIGCqsjtb+FAmU9LGPxido+e5T5gy07M7
lzL2Xnpd34Q0wxL1jEiKTAPDm9CWiWym6SQ9ImP2TKV9RTmoY3AF6bvHwqz6GjHg
nYzHwhHc+mABE+3vpiUt+Aguiozu+Tzswi00zfc1ZH5KZ1CEFr/i7vCdM+XUOnGM
Jm1Gkuu8LVlnGma3xRIIa8hHEgJaoov9owRt1vdYGln4uj7LoVF7TCMn4es3YUOL
r3D4l2r9EpbvbvVQl5AdoIpReyTFjI0EhVooew4xr3h19BREpHKKhJhkSJqPALZF
6kVyPL0IvG17WHQPmYYy81I4iGd5rFELnZsvEo48jjW/RjtZ9XDpy+/9lY9RbNfZ
paCk4YFoR/vK1qvmYj2Hu1B7HNiTwDerew0hbP7o8U0b2l4DvXMv0iDnoqURB2H0
C7qo/Hm5o2LpQ+IR6R7sWjK51n2mDqxlcPbgWdA8vwKgcKKxDIJmeAoCK1MKg9lu
O5n4lEH+c2v0A5voUFZRirqYXAij9WYS90hFNNMPHJ5s7OoeXzmWOESw4uBsM090
/y1DOrDmTp2A1hcG8MVq2GaNxCbW6L6aEmlUw1CMrPafg4VrtoorqKLNmS4Y/0qo
qd1j7RvT1jJOaIMCY6agMzhwvPOW9TXgyM6xmTL2F6kbeXKRjdEr4vow0zQEiqKD
w2owuuk8n1xCSYzdo9XgSJVKB8yl5h0jH6IIYHc8Y+maOLuHE8FH3x/7fqVBTGwr
isojsoKDGMy0V+SKb5rhZI1mFoP9wmwCukPKvGBxi0mDh83pmEjSWlWzt2k1qDse
HJd3f3Qmk6bqIB5PvVetGmczVfNTUR78g88mC/rqm7HSnUog7+WCFA7Nps0CcWKF
jriIgHCVu3Wpm3nEOJZ52Xbkk/SW99+S/mjUkc1+9uIcJIAi9WZqpUS1xRw/BQ7t
wA3c9dBCNlo63YBzPVSXfMMdr5mlgwnl6bCqHvOHHnORwM1henaqLLVAC/rIOSZX
DXk0bFw7bWPnCHqbU5kqUmvogeMOGYAJk6x7ED/NrDDmfQxOLvjydrtJ/A9A4zPH
Racm67/xavG0FFe9CkE8XkkkdjN5DVEK04QBqU43cmPWFnlN1WiEVRxVQW31fzue
wV5VhjJLZE0RJzJ+vBIX5OWzy8szZt6k0WB1DuRZ24Pnr7gRokbdtnFjefH8VIZT
i8OTH0MIfmj2UZ8lLl8j5/FDqtQ8ozc/bBjFErUdMaVr1u4wXTBJnIVKooF2Z+WK
arq6ty0+DrUWtwcGK87GNvK/0NpwrZUb/jGXd+VHJJ6PE4ZEXeblGiWS7ccf/9/u
O9yJCWcVSAxfYt+OlUHD28m6VbhB9CvJTujDF7i16pxwgG7PwaZ8ScLJPxB9r+wA
2b+OxTI5yGB/aVn2wHjUAtTldrZNTAPZb9IJrEzhFL/XtcyzXYHoN4HbvwJ8Fr6o
n2kz4mRSTgqOeDH7IeS0wJZ4sQOdaY04XsSrijpYJWbwv6Mf3bkhkBnpxioxYXF3
1Ap5Rps+kNGliCznzpUTLf3Re47uIYbbN4drtr75NwIwC+L14B8uVkbi24GGYg0Q
MAOgQ4k9n7FhQdFyk8CAbolr676TKEliSOgcJEJujBRlEuEYbHUCwSQsWWDk7mii
KMm7SGRJmyfpTaX6TbS3GrZOwUQ5e+Sd0r6mtJFNZOfMT0uwdVVk7zFOrWm5Ngzw
egjeEq0xJjLWynmYq4HaHTS2sf3SqB0t67R6V3mjqL9gPdpymJbupWtjOJbH0Noi
HIFkwQT68omQo+d24lKDpeGNXrXpyEZlc11x/hOrgjXUdx1puHWmFd1J0MJj9AQg
EamPbBQPkm1JVUkeFYLCOUgVWr43Elm1FJeF0navVtTKPnoAPM/k80wN2FEhxHlx
rdhDb5W4YoL4NTi88vrDk0Io9tNMNlXZDYbneY4AqzCDYVxHDOBY3I4pjvHVvhEC
HV+u/C1JZEPph54lePWTEeBOqlg/YP28Cd0JofAwpA6eEGJ/Bki5eDN8qlHApLFw
AOSvgvS5xM27WalBJgz/0T1SPrfF7dGSLwQTTGml/mnyCqxM5QSwmD6EGX0U0wtY
tLOeLvVF9vgpQiEuIvuED/jAu/AsUK2l2DYCK5EI41LWf7RylzpTTv/A3njmwbKQ
JU8HZ5lLuZttqd91bovAYxYeBD7/Sq4pA8eHO2I+ojQjzANnwqr2ZuybUTWHAebe
BHrloeabqndCO64LP2cytY2hnL5NnhAB6HpDtuxhf0iNalVtuu8KeaErkXooy/sy
8ZM2nS3bF+yF8ZOg/63ngTEE+KXgoH9omLtq/a90l2h99kE+QLoB6Skyqx8mjlDX
ZfbU7lfif4f7yqlp3/P7SdmxsvxIE3fkvysHSt9glCJY8qUiOmgQik3zdyhpu2Hh
WuZ0B5lATtGzrDirIZ1c31PkSHK4Lqxs2ydXc6l/UuHkXwsfXgHpEMqRXItz6Mxo
jNb820z+t70WGRCO+xj2/yT/MFWE6Zh+2pDbL+2W6WXUKMQyOF2EQpk3zmR8wSXE
U0N+6BHQabiTVKM9CHt18ovWN6+uKOOUAvSMLiGJY9nORyGlPZpq5OwCXqmmnBvL
U1FnbHkMc385eM+MJ7KiRhsqeUUgP3iYLueTVp2m1XzRttG3Y1mecl9AVgI1uzw6
ICHUltkLgzxjk2+1cpP66nQGhGJ8aYZm/34BZLWKN+zU1nFQR3OmqcDXDH7yRRWh
WbpfpNWeSS0MN/JhBbsAazb3TD18VFsY7xHJcJhWxqjiy1D4nbt7DEDbm0OffxSg
Hj11LEl1IOpnDDHGeyib5Uf86pqkiwA/4M66fHDTmSRLhwLdBGCG1jhtsNj7ej4Y
6HtZIcGhiUg/R7EaGUdmJyp0O5fuFnIL8JOqSevdymt3dzmtvTZ/yzoGMxzhuYgM
yOZC4PqUQfeuLtRIc/HmIRQvqkDnkHYa/7kmM6ETjicnbazJ6M2TDNbfgJgZT6m2
nPpjRyH4mkohjiexuUsiujcaUoDa58VHVatBCSGMY9koIFkGK+Z4QGSPdSzoJ3Ia
o9bc893StDRFva6ZQDASwfJU2zz/EfjK0CplhGuZDmuPxSs+Fy07knHhVpJmouAY
hK/WGqSKWjLLr7SAlidnoF2FKPL+bVcsLvks7PxXW/4OY9PS2hyWXPw2ggngQnYV
jFKXmCvHgvAb96MsWK302oEjRIogWBiY/aXnKY3YRlHJIaKiq97vwXHmgq5Vyq3l
k3WEgavlht/8IPjjbo40ZJCfnkjYfQHbmaa4VpY51l+Yj5tvNFSPNWpmKCHkee6R
WHmkaLNZQazB4aSgmLcruH1+jalNe4FUCeSk+WVGg+B+1VZHcVbLJx1vCgG0OI9u
4y/vLoYCyYQEOAAvnDEgPpki7X9vKTtB2/AOe8QG1iO1kGojL13BaOWQmLYMuUCX
LBnFo+2TgTeIudZ0G9A1XCz2NCQ/Fj/kBFll+Vz2GHiQDc2ARuSDjF/xHZgb74kE
1cvhB5wptGslr9xyumKN7CtmGU+GGsu4Z//SntztOoFaac/OMkYoD/OXZOM/sd++
Rlsej+Im8VXAGxGr4dnV7Ru0xyrjMeISotes4ZRJi+VSLYyLl9mpPcbIx61mCDE4
2TiFhoN0msaQCuGwDI3K7gDAbK/I8Gup9IwICUoq2+HROAgDMLLweHnhYfDvLbeh
OKg0B6GWZeoaj6kLzHEpUDShL5sGLUu3lQNnHUeJfqJcq8/3Tcg76MRyQH6HSnra
odF9KuIq4jD9NjsrBxTq9mGVTK5gWXsNzxyI3pyfvBLrBQXgQgCalEEMoB+whabZ
ZuwSmdj7YbNsKnqZsFZOjSxDiiMeH7bMh/TaldmYLrtQvElylTTSdDSoFX9SX1d/
mZ3cX2ty69/qdPGht6bUxIdP3n/mqYiVemfDK6t1/9u6tGLjS5czd1j+sZwB48ji
zqe1JcfF2KDyZCH2K3qXQ6jIBMdzImcTVlwHQjw10K5TucPKHlA/u/g7pPRtpvau
qjiSgYZW2F6JVNlrYA3QH/+QEU5TlJf9wTg90czxW8grx4jjPtIkEqDxNZTzSpwS
fyYlvDrI0sowHUViT+lOT+Mqk5+8jHov/bDyu1eABHPu/7UJ1ENv6ZNaCMmzAIZo
qBAu/+bLftvD9CZFEmfBCoC4fZabW58xc5E7GWiJ8mEiYQfCRE9wGVB7PwPAjzXp
pWoHWwQKTOG6LxUUwcKO3hRzVph7eZ38kFRCeSRapny7KRHcHusKFs4XGTtOlQ78
Ay4wQ9kr+dmRBCwztmcjxYdn1d4ADkGUhYQaEi3WLKvPVbDD2fPPx0OrwUyXiIlp
tOV4sHKR1MBEl819CxcwsKMcwtcwSOCTP9xnVGZ5nHJTOUtKuBHB2fo3IsVVUuo9
PpHzo/cuezQQ2vqobuF0lgi/JxuLzRx6Sp1FqMsj5sSVJ86SWt4s8jFwrN36vC4K
34tNwOD3Qsw6o9D/899no0L2VDcr28Rb0zRy8zOziCyC4eFZQbdT3snBjHy5l9DM
CPiRRaEHEpaniplhbh5Mj03cxPE+BU/+S2X6tzQHpWahLs0LLWUykA6tHbrPvsXM
iP1OJUr78259Rg0sNHK4Lq+fN+izgp4TFDAwKBSrPVLGUDNO/++SZ6cS2sSOQru1
gWTED1Zua56oGoQvSsrc9G/MyIWFAOeg+NvyouAfEk5JSYvQFVK1821D+1q+/j1a
flHwEDKrwjoLe8wlVEP/Qcvf5JCbEgWfy4M/XIW5HbCzxZPkjnhQ11NI3WGqLMzt
KmeTsUx+NlvZMprZoCBoGCJc5bIVQjjwQs+9+rycd5oUiGATB8doI6g4JIEvKU2g
uWf4jG4cPoqFcarbC8wq3TJTobdaETvw4wDxnmsfo/8XafIfMeMdUo+p7Wl4UcdK
m44QertBaPhFK9+ng7LAQZ6oAAjoPF7I3IibQ75mLiZhzKwr3EdAT5Qn0Gu9ol5X
wTQmXNxsurqEC6Yl2uGGf4gcpu/PL4BiwR1kSRBQCXyIKee81hTR6GOdhLyAzqPg
u4sDiG/IqRzpYoRldrt6XZReGegfIvK9JEPetVXUBWS4mf41hU5m3oPFPPTfEvvs
zWmXCw1MZMnS6R4knRxVqvqxv0KerPsnfb+Z4U+8AIv4qh/nchFUW7VCEDq3Qx5S
/Ad+F2Cd841b5pJgXeaq3by94lhpJvSML4SMg+sIbMGhVsDwzC754XuW1Kzxi+eg
Lbz4rzUvQNdfwTbNi6Mu6NzMDDUdR+uikhU0XUgEUF3hINZKUowdUdYZxf4QIwZ7
na4tOvE14RC74QMowLnsx3Oylh2n8wY3ReiuuUaur9p7+G4+aMvm/ibu2126njxI
8a3FQ3jUsSqKHF4HWw2GcBrpdFq+OkoxzUdDF91de0DsJP1gV4L5+hErRR3SF4c+
7O2h8UJm46ya4lTnef3jdQl16S/Ud0eGnG1V8XqTJnmoGVq4DbpseLmaxYj9/qCk
GcWKhIu03wwE8yanpvNSavHoo0pGvpAMjbomRh6jD611DKVo7zD28Sa5xHkzALzc
jOhoeJSWGowH7fI0uuQ07yjIEogHtKzEwe9QJaQycabDucxUwqwPEP5Ktid1mP3u
9wBmzkF3AMs4IfngKJU+ak46lVsTSpEzkZ1bZ2fjCfnXMrr/yJgc9WkR8RsDntKw
5caeAjzE5PIbDJqLjcmM0IIpyrBXSKecBCxCQN1QJJk0RmL1g6p9lcyh/acVFHCf
kiYpIUjPIwKaR7lgjphLLvSwEx3PfPZWq7u7+bZFG84abDVUN6ZjL4GJKh+S56kW
yOB1iFMS9Ry4nJ9ksjg207ZBtyVPtcJVrpW+84U1qPEARLSHjRpddkVRIuA3q9BF
HyDdwvqye4ODlg3AVUiGD+yAncG+hcU0fGugF1BUre5dPEkH9FWNpjNSQYKPgFuC
y4Z6kV04AyTPv8HGZpo/kNaoOk+U8yuC8JB/nyjxEFz9fs8eZsrhvhiSlYA9bBSG
UuPt2aUWSeNDhaOEzsuymS4k1rPZ/L14n+dU0Vi6EJzFC0fXkBNgEbMjVlDENIqu
DK5VjghWT1WsKcy+zFIi8Hn3M1yPh9bgg5tDEWr9madlROqACY6JF339113hdsmu
7Xd1kUokiUOfWAGhFTQ48vJBfV80kcnyDPmVL5R+UN/VG3ioesYP2HkdlJTkhY/p
XA4ShKTmF6ky314imjrQf7+KGzszG/fUQu4O6yHD3QHzwL9xWwkP5nFwPYOxflDE
o6B0gsH8AbuRFnVvL96M2yCzD8gPeCoQUqikPj+VGs3iCALaYA+CQ4qhS+wLokrl
279Si5zjJ3SquYgSQQlXTabcVP7V0xwAQBc9lxa6zAEGv+PEFkYnQfg3+Gnux4io
Ab63nEufUF2lA0ILbX7mHNKy2+YDav6O0CUMIvw3rTTpA4LxSrT5nVnZl67onFWd
TCWPx6HWi67H2wvLnEnaJHCf1/jlu2O296XztcIFMtvZZ2IT3G3ow72gy43l2u4l
KTAkPtGJpl+Irdvq9NFefEobjZttMmvZhzEWLw7ncO6EQQP/yqFEId6uGQrCzeNa
qHsogymQeo+Yj867OTaB9iDMfYG7AZC0MmCHhEcAB7lkXdVJXX7QxtCPPMyadkWu
6lxPi9BTRjNB2hgCcOb4SyOV17y4mJNj375rIGUu3pisDrQEWuHqWJAwZLP3Ajq2
pJt2hbkkUN9GzV6Ah11fG6l6V+P8wPfcv9SE3sg73A870WPH4A7GU9s6Ok2BX6c7
4TZAEghomEubHdYtRFwYH3/F/y4UnZRIgUH0gADCyQp03xFsI+eFosFEkEAbxPC3
xZ2Q1UxQUaRTU8ztel0gBVocI1A+5+AbL4aLY8pnWykx4iMBDITSHJMW0JnrDnm2
u7lO7IyqLvMGmhiuZ54sf8DLHQ6rWmdPajTzm0BkQzcyR4XYDsgfkSJmOUklve7G
rffS4dIhbeqfn/sGYaSqYmGBUP6IIdVkNcs0FFPP6bJsC+ynNScmoRAd2Khr3LgI
s5jOYesxO2BC0TgGxCGwjIZNwMqtErlOWc6ePFmdqKX+TS2HlJOiH2+3kvMXYGV6
Y0M1ocN535cszX79PKt3DQLKNsentkyQnbfJGoxZ4/T1FiX1YIGrFstmwyY00svZ
u6+1gTQuwCGYpkdeE+ffpiqV8Ha16wIFXhWpPs1FN9qm1HYuVbt/Ghq6MBkJyfrn
lKnWgCVHefhhln/E1YCjZjJbEYM2p8eN8s0p4VyUFW8L9fh3GxtWzWjHrm8Lsx2A
ZZHMD9OXH3S6vjKnwl0XQCgXNbdrxQ/lKMY581fbFpTN+kar/xxZE7GwpyWGpScJ
1RWhkIf1SQdcHYEu+KKWxJ48o5qQaNMVoH5OCm+gkAPkPmYor7xQm4hp1MlvU+AG
KR4nxDLh7Qjd5gLfIcqLqbCUEcwrvaTNsr1WJuXLYXV2Ov5B7MBBUcltnnX25ODf
fQr5FqfDlhWVkYHJeEFFW+cxZBd/EglrfzA7IqHQqzYvCYDMUwzGTmupcCE4T06b
bkhzEpnsgastuABqx/6+QFTeF7ryvDyPSEYZVPRKOHNsZ8SuTzhpc2gGJ5CPDJj+
EjTMZuElggLgtpxxRDZpO9UvT/22RQcFFhraGYsDNo9n82baRnXqTdbALdQqz85v
3gkX8F/DaHndOWdiqUPHCGXBDht0rr5NCbP9dbDEEw5m2wrOppyM2GrkfAxG2szY
Crem+r/9uLlr2DKqsBljlVuF4hgwpDI5ILiKQLxOLcvIhQaWmY0pxEHC9e2Mm43E
hHuPVygIcxI9TTk/7y3gFd9ZaVOcdMOecNkIL2lxFsFwVuXGRohY7Rlr4Wtp6ISP
+bwgSgpxzeyX+giMSZaZoC9svrkiy/jtU/4A6fxJQ6VYhSCvu816QDbbYZwDCWLe
wyNhf9A+cx1QYn48Ud8VARIpqGxLknSVHHrgRL6eQ+YypM9bVvpd/q9k2kVd5EPE
l1xc01Lc5XOpRtpgkSHtNU3lNLkIYqPhwv528ZcFYLSl6/k2SFwhNeW0yx1zKTza
4ay4/OU96DMAPcVfIIezA4XMg185k2x2KwP3fijMUvM0XhNSmB78rusY7jy8fK/m
wS0rDx+aIy4qErjOxYwwLOwG6PWKwz9719EW++o582lK4DwkIoHZ7BHeVBcgCI1l
82VZjfa6HmOMxpU5d8x9Ps6/fwCBR+D3LNpyUirt91gjFRCtXY9aLMhKo8ioGiMl
k8q5ai+VTFmirUuPGR2IT8WLZ7/owHGe1b2Le97/wEZonTbJrzs/lqTUQ8Yeg6sr
6CkFiJ3GfmQrh1L1+QNvmrY789+H0OeWjHi4DSoUc+Y68lb6tdgsHXVJqU7DehM6
X+68aG0ll6X//6si1hbia71sdMCME2zg/WilK5q8+4wnkmYuoRpX0BhjrF2/UEva
GNPKIDIAO9plSxpSaYbOdU0ZTidSbn3hudGF+6vfZaf6rj31/OQnPunMZHnIdnz1
XqQLk8JXtLiou42FI+H7Qn6BmSMqJQKz+uAEGnIw0nsQp62iHKO9I9AkTkbWF2Ad
RRpiW4bC6jdO9NcBfdQO57UjjpSB+iMbheKWXtcOzZvAUFONJb+lkq6QKv4s7iCd
8QQCVmhy6aNDdemV5KoPNyO6jyuFSgCdVfDZ7ma8iSdUeqI2nJQilYpsRQHozUGY
ghB70d8hu+nlUVFNcDXORfabDAm2ZJAEfvrFuJyXvaJhrBrD78h34M2Iw9LPB/v+
lfhM/CwxjD7R+tbKHF8jy0xMzBty2ls8nsqXEtEQhf4iN8TwRA7yIapSA+baR1EG
6mQKqi+2cssZsqpVMMbXH98s6WG1TWVIbz0AEoZ5cl4pKW0AmQqbMOhbLZY9QsEe
kWNZTYfy5KuS3rYrtUK0N2wRfIhf4iN2ORAXpJZTqEEk/Nv6Frx3DryXiIZvxgFl
BmT5w224u4CHk76NlQkALRFp3XdymjnqbqmhSJc8jCj38ypF9jEUNs9F7rkpdVWi
pddItQ3D3h7OQfp5F8pb/aHHI1/8U/YgaCgseb5C7iQegWtzaXE7C8pZgXft14UX
qf1wRYx18KaiPuMRAetSPasfVub0LYV18ly399fPIDp1mXCl1QSsw7DG0/oghDlX
k1EOczCLfs8OXaOxpO2xF0IsG80yPf/m9ve0AM7FoIDOJPimoHHQxXvCWpdEPQrJ
MOPauyR/0v57Q0Bcdg5BNq11iNl6I/i23MUbHSpPJQ/zeqTas1Jp6kZfE+CunoRZ
66LyJPMPt5Jj8creu0Lv/9+CW+t2OueUnwTQevkc1YGWnfiZncZwNblHi7E7DWgj
MxhAniGAol/Yx1C/+3z1JQdaXPyGbfU62KaGWExaktwBm35467How4TeY8P+9sMO
dwqdkiU1pElTh3giU5k+H3Y0esvtWIldiox4oWr5wfpsWZmEosmAyIwnct9+sAfz
HvdqL/d5KC5zxtSMdTqDluzryXSYBZfPrHinouIp253yaf0ttcC/t6UytlNJmtfs
3IxXBZOmeCZE3LE+FLosGT7MoGJD8MQrX0SiUBngf6BUsQ9tztsG2ZiKFkTCDOCI
EjGO9LSLN7t83dunt42lAzMiTVrx1GD/8FO+tsZg1hMGQcAKZoZtCK3Kyu0IrA+w
SIN9SKl4HkGmpJ3P3l1MAdwuFqrceSXREfEEJSgm/cTBgoHuwLsopEcStHF9H2Nf
F33qk3fktja2DJ/Y8thSSCpid71XaP6roBp5eBR/JNk2icTP/qvxZdL63RAn1Hzw
+C/JnMM5ZV6Vh+/zuRwVPxI2cQtvmKd8nanOgTy6qn5gU+ibvK8gBfZMA4KzUlBB
N+varqC32JkFGfbMS6nPixt1csq3Q/S92lHTGHVhInmrbYDwSUg8Jntk4bbzvUIu
Vv0Rxyo7cYZMN8YlcB60cuvJnu5WlTv8+8415ysgE2Y+LCPHEiA72TkvJntvaD7p
O+77SnyNObhPrZeVvHhP4LhsnndfwQC8D/L7ylQmBJhe4NzZbXxMN3IY739zaSVC
LM5L4T79kn1bLBRXL7RSh9yL5DZoukqPGDaHAZrVag6mtLtnm4Ac0d8E5xDhDoS8
Fb7Yr2wD4oPFTlTOYaNFqb2ZVfWVviW/aCUiEjbji69me6HYmjPdur3adoYklmW3
icZ+OExt3bn0YBHREfGisUzDXpenhXjLt5jC1J/tlTomstncQofwaaU31swyvZxZ
rELYVwTzExsCMK6Sl/VFzFccDaWqghAfZyTrEjFXgUk9MiOV3RHwgmXKfZluqVEz
BDmyI8VE1KfTcqlmLEWflLqeIbdbPj2laJlWb4fQEzvm5s9iFUo8MzLFm8yZ2FHw
Js2DC1OW5FAoZC6Z9bOFwH/hMo7P8M8DY1P7GMTHr+5gsikdCx7fKKAPIp8al+gO
c5jelNIWs8PqGi+7dp597oMr6nxCnrknrdZ+KUCXgWEW/1KzWUJIEJ4teoTts1d8
nTnag0xMmhFaXBXzMwzCJ+usiK79+G48+iQVuS1WAevF66kXR+Pwi7o4E1iK9XsW
Fl5+CkSuvji3Fv3sGYCaFBuYf7+JSsmK3okcGMtOAsPsb3h/i/MQ206Ze8NkuPGH
JxJK1Np/hdIFnSGJlqH0SbLZ9eAumh0Z77SOOK4NOXb/hJNtVciO/86BGcjaTWXr
rwuheKacmi8y229aoZczKcftAYp7E6LQq17vJ8KW2VcHVce5aIdbAD3eITI8jzHu
9jKTCbHpCOwfXkRJMUx2WEQFVNA5iklkjDrSIyRat8oy+lKsLzLHDa5+2A2TJmcT
eMM5U+ynXWfdlu/I811WiIG8lnP1Jp0llvIKhdcBjejlkbteIvrkxvoQuED/RJ3M
Qwjb03HGGgK2dhzaRuVRXRDfD2hTI/LEiwAKoJ54qCf4/cq3sXpWmq1zoIboPeen
4+yxcCQwmkZCN9DnBhedgiC5gv82p/X8f3i+Idj4lyX1l77uCmOM3iM25cnYAMiO
xXFcTfVCzYTCNPYW5GLDH/KGW37W2A7aNUkuKrlbt/gwGX+Q2eKwAwmdyZDK8dUd
Xge1l0D8fHep41bsQQ7nOdmJVigNniTcHh/Erw5vVwAiCRrIH9ErasW7jY+zdqWu
OikC6ehceR7sa0iiS4Du6ARFDpyHFr0n+yO4O/d65BXfhILE+8HYSf2hZXYWjD/z
51vmgGC4TVak9GXPZX229MUHKAdKjNEJqN6YgL/5MjnpyRtpqAmHHkMX/Nqhwvik
GATfhSQyw3xb2BeH38NcGxA8h+3nZ2doWlCK2zpB+E2yDIC9uQakwfsTX1p0GHAW
9Sfy4IFhCgNFzVaVmPj9rEdNqxcNsWuPgNGA8bGTU8wP99j+fCNbrt2Gv4ur8OQH
9/nwPDK+DjcO4SbXhAKU4CtADhFfdwsbxRs/rq/wL58A8+7l/QmPZXCw926njaNv
rDNcwrtD/HZWIAk1nQmuUic7I1vQ4VDmVcGIuP5eW4NaBxBuLw8lQ5UTDBdeCXaE
YdnGd7gSgHK5bZsAkJqUpokhkTepj934BXUoY/FG5X4hBLBi0HNccLP86JMdNTBK
E8K5PPeIe0nkY2tkcAG7xZtbcNEOu6+4c99RTQW2twGjw6zGBtC3Z3aLWMhYaYVc
ddTF5zdSvDDnmVsYy6oQ3f/V1Sj/3BHX4XGIDu44thTRR8PRgGTsoAiO2x9LtkBz
BEkWsguGzI7ahZh+PuGqleazJBhxRXoWG4UtfRcDXjRnqA+rB9ST211dkB/5bkdY
7WMisyzApVYPcOFb1tcAiRHnbKnT5DEEqbFHYyWk2oM4/POigfB0YxXSKAMSwavo
CNgLIYkiH9LS8eCrk64g7qVt+hwid+QR+6RQyO0JtW86LnL5YTHZxo+4cfMeFIGr
dbOmDCBrk/mqYfwbo88QQt/PdK1L2uBGEfOpWWRMz3b181JNOT4XTdQ0tNKkJafV
rMJqBoPNg3UuzaB7dZR+0l19hnVIqn4+oM7kdFAV+AV50RJzcPYSFtSaN3phEhJA
P1Llnt0VLupU2uYLQphC/LzzMRpTXJGJn7YYbPxd+nUeIyujUnitu8K6xEOmYylR
D8WM5r9LMgBkE912OXeojAcIo2/CBo7gWVeqkSt8i1UoZKB1cyRvtXum1OzWhuvv
oA/M1qFdQeVXb4x4XZf6CDzzIuu2wPq36m11TeidGw/mymwxFpKBEkxKiyA9Aymf
TKF/Gr4f7maCei/DpsguTMGL3k8KPs6cQNuQGN37d9fypzQJrSTzzGAnzH2udvcP
uBGRoUdKGokT+eooz05P1UNX46jYgVBnwjKN+wXRcCLhZIrwEaLt9sNlpxpWkd4I
Ulz8km6hiZvJp+pHWyULzui4+as7OHip40I5HuCJ8dLCvzZEVzTzR1r18/FO06Py
0e5hG7Ggmk9gh0yUsBpQOK+f7jOsZ1puG5bnufWXOoWW8xktGLA6jl6KOur30w+3
9y4Dxj1Nm8WnFK9jYhSd3PoTwRONj1apa6oYSl9GQ8p3cxbJppFKw2gINVkC8Fz4
z2H2jousZQM+oz4CNoUPtB93bQFtttTYgDiJhzqNHmowRkrvbcEaMIIi0XA3ncYj
MufBccbqaoEmXjUxGFn17VyaIDcPXqPcw0/ATzn7PWGDOhvdLfZWyEv0N5B2KPbh
G8l6Nmmx6gpBkB7MxY486EpHZ8QQUhlJzKF+rz6kDGK1RLIov117aSFdCMNhcJhZ
LgrcyZYG9THbNHyZ/MuFxUcw7tla8vpa/LpZ8Sfpvnc269eC5B2tC4+f1Mz/kzsL
rxtQSh5wj/ob6VGFKm2wnqGuhdAjdrRukMCVDwbEayBQJVrIN6JpXCaclNxnYhBQ
/KEyRJysKhoLPUY4WBvkOvmSIqW4U673gsNpuviuBXi8mZzJNpqyB66xcCkHJDNT
/lfeU1IvF1CUdeDG7SXWOaAhm2cMwiYNTPnQ0bEL+kD10lWQgbeonY7C7mdl+o0X
Og/IMbOmL7oPMtseR8s+ZOdhaz5DswZL+H7rdsAl9IA6jghQB+uw+W+dTF5Jsp1Z
VePCXgvSe64OmsJXW5eSODo0gwQ7LRjlxGaEqGIznoH0nX9oP/7AkqQoFyfZXs4F
JANpgGsYdwPu4VWnpdbZaRNxfBLO3506cSqXXr8IcAvp0hVRcVs8sDjdxw4OCzT0
7116kwQV1/pTbRynLUa87xJE+fVLrdUprfw2GE5a9YPSqdT07wepzyv2PpdnJcaw
l5HEjJuZQOIQpK+V4w5ccy8vIoryw0Zho6vSbIfodsjfRlk7DTt0Za4FWsT/DTxF
SzP6DJn8Oj8OJ6lcidS64zKREyMwPkg6JriosCQt4cR2E10B0G7RqHzOMYj20h2C
NLbdTu2Qt7XN2UW/aPRwNqILqPNU+GPBGmM3AguSXangtEUowlCmajeF6SjWRNmb
mylxLLraoEu9XChgoBRfs7LVemdAMx5Pz+DEZeBrdvaT/zRWDMpBtgpO5y0KUdRG
5U4Nb7idz8+zHgSqJigs5aLChKASDaOrURXQjw+w5ufDz3CpKqAyQapR1tmZg11d
Pv4B3aQyoqILaCxVEmOivtIUuAKtpbh56tbMUR79cJZTokX9xPk3xq86m15quyu4
7vY5IKzg5M/FM5CYkPkVUf0+auRRE3vfMzo9BWYHe6K/f1qE2YwBauPDO6SbKo3a
xCdvmsbCb3tnyJG+u53DT0UsL1SSN/QaCinlcdtpLLjZZuVxRnIsVZdo80Kn6bY3
o6RSfsEeY0usrGOzUwC//8pX0Ox4z+gXYnu4pPOPgPuPHBpXt8I59Nmu0VB6SACW
zRWSzHtcZoe9leJxOocrt8UNfWxvAHsUaYJhCNJti3RTHmM/kUxNgvohqFgkcN2k
vuWz8aK++iKDxYL7gjls2q8qply9E70GWEJGHdRqol5Xc3Ofsob6MXMOFVk71U92
hUY2APShjvqxVw8w8YSfdH1WjGb0DoGAflM40yO22CUX7ugvAhWyOAmoEM684YFY
uiTozj4lfsjfLCgYkAhr6Lpk9Ht9UazNOViOT8yhyihGpgDWOm2MTxGcebcEYfxP
3y+qsheE8rlQU3gFnJekL9IkDtAEPiK72xRol5j/m0gYHuS55ti0D93ce66HTOJV
7hAGwqy3pCjabRXyAG99mK5t6zeePzkBig7+BxMTwSOvmbFnpL5SPlD0+zDJgmiU
ffkjjsKIUc2LkOTzedt+qDNDw7D5s9qKpclHmKQv5Dr0e8cT2qIQfhmNUJaw8t7w
XArPysv7Jw0EfUSN8zzFqW70O1IG26o0YjT7JYZOtop/wcHslnMtKF9IiJYN5Oh6
Mweu7MNug+3AoEwM5e1DvTRi9jBV26/FO7JLJeMArlk5OJgrncXNt59caMybOm+Q
e7OLarIrbdFHUzaCYv31nEPUXYSyOSMmd0TtzGtBPXHJxNDdZ7icepzzH5zs0ZuJ
J4eUEh2k3F4i+hJtEc6xr2sIHUQwU7YY1JAOyWSOj5rIQVRnT0jOgjgHApmOpw/h
moKmwEr1LoYGfzx/7A4p3u24A668cnFbTHX3hoEQp3ShGVr+XurM2hmmypuNJRzs
HA4633034oP4s/Yf565xdMXzGH8sbr4hQSNhuOuITiwsvZMX0All4qSn8661RYJL
AS6YmrsrU9WoOOcHm660Ub0kt89/mhYYop2iZnj7EcSaFsACiPdIwqmeAmKpEE9F
pFcsCVeDHZfLtHtL0h8QZlVfDc3xxmJUntf/dX+Z8K2DjBtRZVMenAH/7XZRoIxP
0Y0Y0BusLj3LbMFe7BzY6E4TSvk5sZ/CRcvfebnpZzMBwZotrivsC6r20QTq1Umx
/ghDI8fFSi7rUQNWuEdkSirNEYBV3uNoCFWpaHR4DhokZWk+UsSDsxDMbxs+Kkh9
AAMH3l+VFxJXx5QK51lWgECRuJYH1Kxm9eAQ788sW+zP3EuGunGaprzK/JKrXggb
aOXham69+SYLiW9BXjuM76wCbFc/L0yAxernAZHV3KKPGlt2jXG5qIaMaOw6aM7q
qfnHa4EnHxYU9MHwr6y6g2oh6f6Y+USzOb6++DRQAiu8C6FYkeyUClX+7MnNxi/W
Wh20dEbHWRLmJcq7iXP001lSLngsgxQRxRhfXJYxQNplr246nOnTKEnnwGiLcjg/
UZdJ8qr4lUoFQC7kJI/7Y/nTG8/hUZGbbBdeot443zcD9BbRQXuH/npxg0pF67+w
LMjR0q1pYPcgHVfIEGSl/B0zWbR1o7TMkBO9xCjT7R3FrE/Vyj5XbXO9J0CCyfp2
+QFlJKkFk/C/iwRAcy4bZoWJGFMbGOd3Pyk2bSOTl+ehLlE4MOZtbQZGjO5qR563
oNx4ndVz+H0U3+dGWkZTnZUHIxS58w8FqPPeg7RjPm4DvG8YGHrHO19HuFBEUw0I
w85cwIbEXBrK0CVAxnFpemVuqK8M82OZL39uD88XHfFjDrOPoHUmcmNUdooR0Ics
geZdZdIgwivJwHdlbCJbPvmjhCHR4tpJMdbFUFByComrBwFvcFGfk9EgXPm8bWhg
sVPrIH0DpqKUsoBvPrHmdpkAOe9fDpGOXgM+PtoCVycXDL6oZVzB23xwgjqFwuXU
JBReMHJiFH4wuHGwpy4xrqkZi2WKlkZf3sGRdJKibpfe9HrKSwV6igu6MLpRyokE
DI/tn0cRvhSEm7GBCKVH5TDSKiCPW5aHRt6PDc47aaaYyEORJKlUJ5Kluw6eO4n9
j1Z1J5II4Xm2IRMh3lh3tE4nz8Uv/akDiQanfBf+1vS5HGrnYJ5YxAHIauEGgPdA
r6SpZ5lFfSGlVX27zS+ugLyWFR/la8fJJZBQeKEfGiamXjG0ZSHREUsvM4dZb3Vc
AtVf6bDcwsEt2UKirAR3v8705qVarNp8aQ63s+cgJ6B87GFNASjdaT9H9ajpw+6c
O4EPf6pbCycfwXR/L3Rd4f790DlOyiaSErEO+6Jdr3aifj87ASpeic5rwVL8TEAG
yMB3rJN5fQCfNY773RJ6mOA/FlUe/l6m8Y9gfKoEIc3nACPTA+Qw1XKQzDwqgeRt
AAqraPLmbq5BDQG/C3gDUJEO+5uPtaXID3G/egjlzv0gZAfxs/aVwwpSEQYNLS5F
QF7fYu37rD1+hpY9yf69Xg/GTBfn8ugzlBeZYaSYz8YJcklmxJ3OTX+4GRAHGMxx
D/dQkZqyFbhwBsWXFVxaHzfu8K6+m1UMl5Y/qisz5PXu/UwH9P+KiKwRtWLw6nDE
/HU8DGnFXggbC7lZZmW7KNCvseLsg3gbEh7aopKKOA2M9c7AgxP/XckEyWc+5JoI
EodUghm0swM6FO2/UyTo0CMjnvwraq7vQE7ARWtKr9CaGh6cc1DUYL6Uv6q0rCTn
mGs90Izolrvv9Evp3hkRDgdOSb8w9ctX8tXbSM3z5tmNgJ4rn5NE16ZD5+ASMTqB
jWFoId3DdtgjeXHfQNyGNX/6L/bkrU7XcrG18PBtXDzy9u3yXH4XF+b319Yuwo18
ybJUhJImAsmZnQIZVUNxD9R0AEhhfdrfwPr5PbgNg+tgRmWfRQcD6AnJvYxX6LRU
JexpXvMovJJArIZPq6CtTcZRmkco0nZqXhVHrHuXS99ay2EVll/uRjWGzrbwsN5n
zSH79vWX3K0aUDeIGmQx/xxbjER3o566Rjp1FADVQxlB/0BUA5g1SxbBIKbl0h+u
GXGlGH/XSPryVAahqMF7Avpf1Kqc3prV76+jy+tHXRrCkq1e+oLs7ehdTeTyS067
THex7gOg0SgfYBWx5wqFi+dWQAo9RZo6V8TuC6Dz9h5gvCLaei1GYgmw1V9xChRb
DQ95kLTutF0rYOWzYQa6fIIQuXZ0OemJxr7oKTan5/igYv3jPqHWfqjeroAHXhTZ
RFreXL3Jq+qz9hKQZV2vAC8jU9n6lsn3vw0SnOt8P7cMQCNxtWEAQkbYdeJ+qYo5
cDl4DBbQT3eQBOscmWwVcSzfUKXnkqVNP8RxH0+Bf4QhRNF+wO3KpwsOiuEl39FO
rfa9vQB3dShs88ussm834Ur7NrzgXBSVoUW+IWFMVvL4525oVXZj8axwIiKsuYpA
ATTN29rfxuCTm1B5Q71UcBbo5KQfTShJgUYwMW43OrJpZXDavS38K2cKT29H1Sky
sTkoX1hOCKokJKDPOvNQIXq3KNQoVF5DjjoQuIlY692bI5ByJiOSXn7aADFyJHEx
pILVu/sGSpsGYwGIVTON2RhFSuV4qc6xIJSu0SKEokQH6+ej23MBO+3IM1kQ6KZA
h/uwb967mMixErxGnLw2ViLtj9tdRAOMo4vmXcHFnyNbS1Y6xTkajnWLmx5cWm+z
UY5TDXceCgwbAh1EMawcHjk5/VbMmG6eMVpJ9TIgU8Ao64MkgbqgVj958yP+H5qE
4BuN+bh1BeLLiRz3eH8fJXedWzN74jCCfxHeopjsHFnV3u6pEei6ZyFGLYZRZtBK
bmnnz8KaYS5xcsvZ1u8+hORKPO2SmrZF6NIQ1sueXYzzGhWmeO3LkAPKkQS3R+TH
Zb6NZU4PnArEOIPwkx4iAQg6XNkb8+/mcGSyMhfOjq6WwpOa+bZBxWz6N00j6CzR
Ks05FaYH46snol40GMt0jU2nS52sgO3riI0A263WmBN9W6bSf4ODtbf+xmX50c51
Nbpeoz28g9GoODk+S0GCHaXjNwdZVcBlP63Jq8OugyNlL36OjamGjkHI1+R5GmDW
tv58Iaz4/SQlNkR74mgxVvYqWpSQLKiDlVM2xe7oTH6U2REMVd0kqZ9sz2uyBF3r
2+NUgDMEITB+xYxYI4DgN1Y+ookYAMCfINFng1tGjpPTqpOSdIpJ4sB9366bLbP7
KGTUGDoAwWgLiX0nhDCR4ZjCpN8bWRZOplV2R/8rbUwTJjLEt1HQBZAQ425hO9co
Nvj6+8XDpO+gcoCtmY8EXRQ3V+84zV91yqwPXq93k62OHN4OccOH1KlK/K+TUe4g
MaEjG+H+QcnkaWeuAxHQW6r83rlFJm0adnA8doXVSgo3OKgv3WcqfMG8VaHNxFEJ
XXNwZ1smNPcEfiCt8Ja2gxgaNS5VRxdUDh2M8xNV0NwjibzgeCMQz4/ziJ9pYV14
53S37X/VY8esassDusk6VbDklqb/Y9x6E6A+fU2l0yjTHPmSt4ToyCOw25AMZ22l
Sh2OSpYLP42bPMbIGYs21/WF9uwM0PfN3nPDstPaU06yMal0j9AYwU9Qj3qPe9o8
i1AThaIdQ7lUJ1aKc0Xj8zmQ7h13BsFyapT5CtO8POnD/UG82PQSXsKqf01mfXKm
snLjxV8/sSpjicIEqDr6lk2kqZb7MlzwO/IOR+SfGxULUQFF3Tx0MBJ2+daj53AS
rnn74n6G70TQloHOkdAc2wk+NMBoWeT0gWz/Uq7UULrHXFJ+21iRu5sUIdlrQSkq
hXx0/aJoqJmBhqlGCFUK1HPUcvp1beM80BhNybUzG05r6W83J9DSaE0Ur+XS+O5P
Ntb+d9W8lZMWxh1F3dUdC+XxPiC3h1Hj/4uFV0rua3GLpBz//G4zXnB2T8tSuX14
OjjY7qrd/mdFXcxw1834iM98jlkHapgVvcZKWWLff0XBlapDmOmUnNQV4Wd55tW/
XG8Xl8Nn+iv2FsjmOnhjmI8/8b5NQbsynQ5g2O5jyE/nVfJB1jqQ8FPr0ctWvunt
WPU1GYQxjPS0qNkCyxJ7aOT6yZkEBU/HZXiu+DGwTHO58TxJsQfGoipABL84Hm0p
xT+YsmX3lpIX9Nj/OHu/mQJCLqvjk9NzzqUvfIoTQFcpXKW/rPlXTMmThXTDBPnH
WAnw9iHYEbk+FZqdbrpiTBC7nAfTAHcA7aLXZVC3vBxoeNd57wdL4Tac6vYFZLXv
GjOVPZOnKiWPPduz4Be7jA==
`protect end_protected