`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3328 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
hRRAlfE1xLfeNfywbrz10PFIdNIXw4fzpklK6LNOGD4kJuF9A2XITegy2yWBb/SL
ShTIhDwU5C1e84fQP/mZ3j4pZW9276tpvaojA09K/1xAKMu64fknPjbMPHPT7gf9
rSRWGzpp+3V+63H5CSXcktDf5chGV3lpFT7tw00Tw46p/lSX6Er22xuwQ+AQMjeF
KA/+gBfS7MsJ9VkD6z+6T2HpEDaqv6UPoWJoVb85GgA/+kuxL6XIvxIYOD/y+peO
obYwtmuRJy3NA6uAZa3qnoJTqbdZ7PI56KqCiBHR0DC7edRWjtYJrvLb5GK+ccqw
KNEWsJoPnnSLuJoXYd0qLKr+5zaxYOI6FDjwm7s6CnYdghJFuAAKM0O086/h0Q/U
CSUCTHAegMpOENkM8+2QHk/dofKoX20D6uHcs4x0I4ompVumHdJmzlCUXbFQ0vBD
+K7QVZhK8CqZfEaDrLXRs8NjNbih2PimadrEuvq/ps+ttGi0egOIquRAxUYqc+kz
93uDsrS6b4kQnCkM4LMvRiEInmXJfxuYMiExXd67+Yh5vyG5W0ymDuaCqHFiGwi+
+OXhFxWFHuCeFPIE/NY4W5CplwkLqEIOrbl+trXBOwErs1TcJ3EUZf7qNi1k3uy5
uwR51V6U233ZR2FV1yDBBHku2mm/MBqsA/b2pgRsHpWKgm5DbrE+lTo+3TnBVf2U
OqsNZd4n2J4B+jpv9alGAgPipMOUXa9sG7t/cWOO57Oa1nbFzKuaSlGMXinLk570
wqTQ1vfZrrog6DsCgHeCZOIcH2p7HxXvIB8SyJVJ/V2WSvYu3Ln/2h+lgwfGCl5N
exJv3JTecAvFQUmFKntvivhNXQbdrM6m657tCdnJ6DRBHTNZwqjmHk/vK7/y+wIa
Oc+fD885n7WVUw9rB0wCusdQvHa0iGtsAxKKMLECqV+xDwg4WdVroQ5fR+8kI7R9
y4O0GlFj8nlZoJg2U3UV6Km8gQZTj0bRXcIHRQTwwHybirkFYNeUD8hTijGKd/pQ
i9RV6P8YxH6lUFuy5L2zPBr8IjF0cBcg5nYZzlrXIvrcZKwddepSjfVZyWYAcWIN
bs2FerfLwK655hHxv2Fuy//m4o6frnPEGV3BW4wL3HhzSLlqTXd9l+/G6cT4NP3/
dcpGqYP/w83iQhWMuJPXCzH/0daWEy52IENl8KWfxRmekyLbkMIVJKiZDQOJQVcG
zq9apYYk2pw+uF419fMtPEmZJrrY3KX8yNgf7DMx0q31vdMfQ36I4fty9ttSFfNL
IEvHi1kCRHS3HpbQpZkfXQFKjvdf/e18iUU84QQ1JUysIqhnFWgp7JhONPLgatNb
Jq8hKjhSNArLuwq5iACyYqROc/+oBCg70abKtgnhWgeVMzYY81as/y0z38H+Uejz
SnW8ce7JYSDqpIEkW5ZrxMwtsBmamviVWUs5mgm6ySYFxvrYO8/mEGA7tT6E00hc
ME44ZnX30vlFYojwqFRa+AcIzAuSwSUcs0fZ1TtxC6nYydzSPhDBN226viPXrwAQ
Rb3vnPoPkKD+sjA7kir12+NwEMX/WOwj+jTPyPaarm8NQ6HfVLZnMuxAu14DPObk
sSAEnZwAJUij8KDsAZp2kY/YOSq8r3NBi7eubRr3w63mvUP6TwCX7PBn9bAgzyOI
aSmBFxfbqY5idEkKdeLh3uUyobuxis83z7eCRZy+a1vhetuCj1osUhh+WO5+p04W
Je+F5AXIjRv6HUWcq+1Ricb8iGGHO8wu6FW1JTds2AsHQMrg3tBCncYL7Yqcmc5+
6j84HmxbatfZD6RAAsuNSelygmKDOvc5HfM+3GgmK5KxaTyUAIHwLmCzVixi6m4g
SsPHJf1667A6mP9cjCNZ6H3jXzLQFrfI207KNB9+88CQXRxWxNdx7BMwl0sytToF
n4YzB+d1S2XCz2WKWqbBfXC6lKoqfb8A+Vr15w1UHvReZIBCHc3aBwCgjI2GG+P8
BbLStByNX9nUFXxagr7+NV+5PLPvn3lC85hTpWe3zEA5+7jzKR+1F2P+n/hyzGpE
xASrNNfNaEWpxK/zPx6X3YqwLfPv4skVb2VHGajB5LMQk5e3yVAXpvKuP+0QXbf9
dCt8sT8dff505dwa99ZtSinHzqozssO7vdhCvb4cDfOXiZ/bO6JOwUw9hfsdVPh6
QkMb09izUviqajwnX6C2zBVwtWpKmGS+2/YLSrCfpTihxhGwFbR+MdV/B5ppULZY
C8aHZvqEVH4OyDzCk9dzG0EHaf/VMMBHAkDl2R3DrBuLXrEju9nFJovyEDN2zJj/
3KIf49Y4vnUGLO2qUHPPUdf1EEhG3SohHSlJbPjXPvyfkf8L33NPCO2WhYuAZXMV
rLreT6L0U+tYzu+tV+dsHV/O5Fc3fcdh3fz0wZr8AriD9knb8xCqCpKdqQ5IGVNp
geD2Yfz7rimKuQPWlWCIfIaQrvfGFOzBpXExBkp5yjlaBgEm9ZNN3ytcPftZCZyc
9a1jHquykwXWQqd4bX7tZ2smhmX7kF2f8Y0zPQu4PKOyMwlVFAwDgEkeaWR9/1lo
OIomm0aUJnbP3iJwwyhqkEG7G3Woc/9SBL4ome7+VmOaGXfYIgYWZHFx6KhxtjLV
FXCQHSaHy2047TV9Edo+zhW8QeSkj6uoUGA54K6LGd9TOixpHQpgxeub0aC+wNWf
eesXhGe/hW1nuy8Ou3IMIG2N3inG/Jx5ykFPNRM0hd6MRlTJM5cMpidd4HvYJiLl
Vd4R9wgaK6IzB//3gQrACYHBrNgtXHZ4jfyYgUxCwfD99mI2B4Hd4263+N112SCJ
8IOs0j2PEXMEY863IxwVsFxR++wJWynn/SPrcYgvCbBx7nxBUNxLkVOVv17iKNsj
DhSL+5DfQuL1UX9uB/ni9brXQk4OuPHp7TxIBGOTGM8BmEh7bD0TPctfIMF4scx0
17pfVXn9HNtdPwrbZQEdHk+AchBC2SE+KRRwDNnCF1l3AgWP4gCnKXajkm4GijoH
o3yu4zTXOgadt1xfCc1rk8alWASWGgI2FaiEuCPJ1RCqpwc96ViES8oCfsOpvHem
71RffXFVJq/D/qmjEfE+t46v2C2vy3hxsVeq9xWPjmRvLO3bzyhztYQqLaKVDdS0
Vd2F4RibmoFtazzGevUnWlmU6vi/MODxOigm5PeiKBwfhumtDgpIjJ39Zl2Ml4bq
esGDc0yZpZvh3hZ9waRVXEtfvLUKeW+7SigQIXaI+aSmuYB6yhmzdfxjbwaB62vX
tBXDaUl+062PjE6R5nCDKeXo7tRiPfmlQfnV3lLX4d1eiI8b9oqEKXYg38+gbeaJ
aQ83Uvq7xZXgsoe8ywbicDrBR1KU3T9RANxnTHZ0lXqJGQVGxkWAu+IURNI9vWl/
zcnicT3J8PgNu0mecu3CyMrmNrFsOeyaKQGVW+6kxI6iI1Mfa9Omnz/8NYYHbZw2
DG7NRolOCO2rZhjwAgac9DAVrJYTKqzWoa/H/2TsTgQZfPUDN0PWichOOXBMP0kD
qHorVkVBGExuSOIzsNO1LVBPjNthSJtdWDlnrtS/pBshRGNXeIgkdnNMW5BwVv+p
YwiXAX8hdQFWHM8xyu+A7jlust4Si8ZtDmtjaaOGIDmPaYKrKHYonIVS6iQaufTs
nc8QAywV0/rJblCiNeu5PZ02En53iETgde3dpHW+va0ri6R4KZ66ZefONEJfrI+a
CO+5UdVysTM1Y9S5NjfIQKy30VZTmODVMn52Rg9iGPXvAeaRn/EOyOz6nEAnAnC8
X3MPRHTFPlJKmeszgmZCgwHUrJFUBlCEEWXToUzoFn/VoKNMm6jc3J0eFuiFtLBl
08HSDHjTJg9NvlEuoaExWcdOA8mMNRJsINFPMc3bBTOWR7dv75KV1qv119ce3o2s
d1pe1amyEf/22s+8W7b+wwRvqcYkQSet62f79OTjsWWngOedjWEQhcOafTztm+qw
Tcr5LOtTK6x6/kZbNIUBB6w7STvg+xaiq/yYI6bE9R2zt6PAHhfP9sZX6cNartsG
MuP5wiKTBih4dhpJPvJVNKHCCBTKk7xpD6ML64f1RT7lYTApS/YqN7DIvHAj4bz3
V/T/rGaZF2DcNz0s1n0X8VFER03Z/ejR8MMXeoNNOygwO5hJdncSYbyjolrkWGG+
OiP65O3twjWlSBtwEJLsjlnwt+wS/uGfnY4I5fojSi6T2H0lfe7k95qRMytmM9ac
Of74sg4C1cK6VzfG+GSEmv+UDjeDH3jcIXRYLoNUVg1wSIua8U7tn3DBjnqfcEIQ
b21wrs4yUbhH+B2MOaKhgw==
`protect end_protected