`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7152 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmWdo24EC1SLhDeUV9o12ewQ
ulXp2xSZ5P2RSggIKJUy/anaBVTumwtXp6e/AWaEdufYiqgD+zF6LNG5i3xi3hMf
Fc9NPZiLDwGM9bIC+d7U/g6RS+C8FBTCaQuHrQ+wud09A8aFAmivVajyXrDQEVKY
VfcShPNQv8HHIezET5jStBYIecfJpKyohgxnY2LCQk12jTPVJWbiqeo8UgZMyfMS
QnCdS8p66Fxcl8UWRtYRdWrzeskYqiG5JCo7dp2LcoNFa45LnBSK2lcSEfNcVST/
pefoQlguemXbBpMwSfuuZZOh4QrKzIwFtymqGhdLrVcxM9PejvXc8OwZ7j4PhrSg
8FkjEd3Ob9gHr9Ge2BSy3VQ24PsIHPkHF1EJ/xJkHsMXUAC73m8z2ZFVryknx/js
ckJKg5UTj7ObPCtHcXb+P3mRbvNGRGMRUwmX5t9xYA1zKWXk+Y0vr/w3cQ/E+xKE
NbQsewhuGMN1pLM6awQogfWJ9Ry+a+A4FFANzMHbGjJbHeYXXuXxNag0oLHP8ZRZ
qenX73oFFnJfbkz3Tmx7Wj7yuJv8y4IJHjB2ei9goSGqvHu4taK1nzg3x4ZChyAh
k0/lan0Nd7zuLqxTR65zfrq4wB5/rYULt+VbTcUv5RLd2I4KDYYG3Jj4Ok9GGwfr
cY61+sW1SiPdgpjytayhJMZLJn5KR2WH299/nHlxRx4tHQzGUncr3edWdxiV7ELK
OOnMbcZk6SB5gWevnWnvxKLIsErVOaeifNzBo/j9wb4fy1ghjAc3OlvBiLtfH7PE
2CbD9eawPW7bEHHVSlla9deusJyeghDw7zH0ns4h8evoCfI0dtTmHyVJvlTPTuDO
Qxgx4LDr6FrfTSOycijxSET9HStg7vt8TfPvfSqPngnU/W+l1ADWu/mCC6L4udmY
f/15ROxkHnCYuvYbjQVO3yPcYfeH5uYjxU+mFsH5SvZqLOx3QNo0omqiQL6SDCrx
7q6L/AX7q1OHUE9ka7U3CEgHpv2eTsLRhHtyd7y9CKNd95iUBkbrXPgTNc8s4HOz
11/Zce1EpIXnHnj1UKh9RaysbqPtgsNp/E2ICYjDEHUflinjL6dAfkLd+qfDMh6B
9nlF8XH49XpOhGZ+BEreMzbj0RMCUt8qLcq5VzMijO+dSY0yQk6mNECxRDf7WYiO
KFX1ZTlDEyNC2okVF1bUEqA2oMrzCbY8OfKiI7eAPoOf+DhKc0X7phI/GVrFfQD3
lAQY6OU0LUofq/Bp7j7OrRLgdpIUUzadm4bl/kSlbHHlskROo5TsVlef+9k+25re
xiiJBfcIhUHt0t28UOdgnBGFpG6WmxhMrY8Jt6jSm/xH5OqglEqOx6HeuppM5/gK
nfnb+PXG9ZkEfAw/X7hNZV/VdXHXgSoqBrIIvHyPBr8bwEVdxWJErbw8iXUpBvGV
fa944tYfaHFI0RQwobVtEnM/uH2avFl6TfEBqH8cUEZhuciRuPcCVvaw15SpkNV5
pGDmCKN85bktjMggKSjmbwFOlzqyWJOChJa92iJNyyYjoHAXPvQOhoZKqGt4vd/7
NIfY8bcP3Sv2IxdoM0Bq28vEL9G7h3y17rpxI+kSA2q9A+vJ6dD7iOntqxPju87P
Pna/cr2NV493VUpBnfTfHJQ0yQ7S/5sqaQ6RhgPR/uTV6YR+nEZw9ni5gGLyoI/Y
uWapd4VhG+gqiTWtLFodTi+wl2AczXCLMCDDhTl42WzmLfDmkq3BIMBPP2EIyI1W
QfPa8qQrTNBzkDPGiawh4AEquHnWH4MKLJRUHYzelXKnXkG7FdRiMSfCQv6rMqwz
CE+2qma7D7M0Z3SedkFGJ4zaOpa6KEHRptuVIxF8rHvCubNXo9RrdN4PfWO+KAoS
ryuA73R5SHchLE3oHG3fY4KGY7L1OxMjjCECT70QrX5yVnP/a+FBDTvwYw4mjFYs
NgJfos7v9TQ3zcQ15IqkF5oet1rD2SehWmqop24TPlKOPoRuzt2A8b078VTqD2X6
qgWoq4TvHqIk9SOlOYpKsIiYIJExnSUg4N93wLw+ZjgdRJTsaZwAyOhxLn/8K5/W
IRRS9KqUt9cbAvRm55rsELkv22NQaHmUULoe7vpgnabNzSns+Hrzp2WfDlZszR/s
ji1SjtfzvwCCRw93URv6k1l63gkpvbr2Fkxjef82AkKrWp31s3EY4td0zFrCzZ1O
RIUhhuwvPdR2YUAWJXSza8yFWpX82kgdtHuiX1xN2WKTvaapltAqd7Jf5UI7uebs
Ig/nYBCT7H+grzA43yVqRzQU9CFxXIP2zbD3kFdnC/skv/3HVqKyTd+PGOclOuYp
ASBY7ynBB9602MGhUc2t2qLZLRuI7sr2kPz+RkpUf4ZEJlu35TbNjwRlW5STGow+
6rr9Y2kvn3O6wKI2IxlfVEVgOr9PG4Ki/xVX8frT2CEgFZFoCbLy5ctuDy409UGP
Rg0Z4SAQ3u3YQFqUodZBHXxHuU92h2KKioFhM9nPX8WP5r9eAfvTZytSzAoHjXm2
iqOGnsRpGJ9blFBBe9acb//Q+Zz6I4r1frXhT/uEO0ae9/2gcG7/pcdbTA9R9ZXE
a2IvWfwD8N7ZfFB6DPRMGaBj4bRsUACGrOs1+4PV/AkBkGa4WpRU+zJM107ryO3m
53YiRNgJcGdxIx8Rn9+NVaLZKV0tM8Myoijga3OodeEDXflNMEWBbjAfNvESlUOg
a19WviKQ4in4ux+eYKCBysNEy0r+RpjY5m3XOwfquK9YEsNVQdBhfqhA8Gwsaqd2
C2ZMtseqEwSaHJZpBBV0I6PYSmFSY2dLyJozEyA9u6/YryzMnsB6hsXMpM3+HzbM
QG7K8RCyC6ZwKYDrS7htgErWkE08nvUUWxNW9lEsYZLGOKW9rfGb8FWB7nP/E2Bc
pLfUF/is6kezgykh6FXdvl8MxKqD6gloYwDPEIaMoRHqxC2DktYWIzWgfb8CS+/y
wkxeY8a2gjhqaPHmLVfseeOwh3u/6MQC6ArND8/2FUyUF93tS7VfPSwp3TBVmowX
gg66t0Nz7Ar66KPajSRS6a4JMNRUhloHB0HUvBFXLosEB/86Tms1oml8/oBYa+kN
acHtnbsU3qTlNRCnD0Vn/eFByfmSpeL/rnQQpdnSOCB4kLz9c+zMbybtNzKFDN17
rjodhp+U8FG8072O4jOz8WeZKqiO+uqhm24hnzGPiecCy52vQo11euxBRwJMCYUI
GubNvx1Z8smwuM1xVWMLI8/az+qu/NpR17S023heXbsZBhMJfLTbK3GzBKRKPasG
2/iXVXmPEjMrBFSyMc2V4tomKXq0dNelm1GAGr5w18bxlxe3hqToh3xjY/30P7IY
zlFgS0kCX4eSgixUsOrZFfFSSzLz50E7UR5KypQ9P03tmd8rtBU8Ur2pyvxkuae2
78rygsZnA/ypezjAssedpK6Sx+UOz3hP+eEkbycXJw+2pPm2yLf89bduMDezvDm2
fbGKgPHwK1QveadmhZEwh2Fql09SOhM6Q9ZOcB5Fx91NT6S9s8IajlwAE25cVqGo
+sGTYhHRelCTjD/7yBKUMqD2I+ea4kP6tkc1szRrlOq9QfuH7XV87MQ1hyQiCNGK
+D3oqzFAEUw6cE+BI9al5NgkCC7G/cfaJI4uhHCc/ThMW2wHR/QPuAH1ooKZUQqp
lxSPdhtRysWL3cSvAg7g3wV+zxTogX64Xw/oGxmUZheF9anmhNzyktCSBLNnW8Nl
JF+EEX2goAag66Kup1DWCULJch9MAd0lVD5QNDFWLrW9xpULZHN3De0lhCdkp0fp
TGREbkKEsjNHtEF//srblqVDwqrF+qeFusLriWdqLzjpY5Q+p2GgCepBBW3ABuI7
bFYghrMHEPc1bRSvDJ137b4VdHBezImNy63G3d1+Z7JP+4QswcCtsTveNf7TQpeR
FtKfqFFiBxnAeUYU3yw6/9O/oC+TdjmA10cP1tkuHgXlN6f94jE7/9fEsBioA3Ec
dDbGAk2cYEqViHGg+G3z41mZG5mYDO0hbVyh6fB9CDtTYi1Mek+KW+rHy7CPGBff
+iRYPYedOU88Xz4YwcLAcx1wqNjE3IJECt4B+UhU2GA1/0h9iDF5ZreNh0SfXIbx
z6IiM6C10Q3NYCTmFapRzJS23wZI5GYCHPzQjw/+yHToic6M32qZCqmUpQPc64uk
Q07xY7OnZ528G601JMYQC4jB4qfIcE+60j3tk8IMa1BwyszCn4JzhddqoRHM4Mwq
Q7u2kM592X8yh1IFy+aFjamH8m/3DLpuhThcbB9Qr2g4OXxIJ5GD5QstVWLOnl4i
KYeTvOM2V/Gc8ukF+Lofg7ZnlR63pOf8K8WwOn85mSFhAvSwVVybwvdZXJp1o5w3
osoDTkJAtLFJPg2dXalv02MfC2eCt5WbbXFE5GPkPiZaYz7H3KvQgLeBFMapKzft
orqyDy+6n4FcsbwJtYkFI+18lS3J4GDFMhKPWDvAwYxfkDVAMLEpuia9x2SYDzgR
0cdl1ENrt+ZelMThvPjP/lCYXKKYNzlGoDsmLRf5Rre28uEQEGHoK05n7nGKSJmd
T8tUGJUNgO3bkZ1ZgpgkMn3K6COY6o75X4wEAy3wsD4Yj6JeHoOBfhus6E8TnEG7
NB0UvIf0d+TBaTcHHN5FKz4fSEv2KSSi3rwtmreYmDGxde5lm2NrrDgghuAwNonn
7zpNvZCNvX1Ysw+f57r053EHfhRukmn8dE7b8pEv/0FHeusGoLKv/NSp+3Mwk2Oj
P1sLApPv7sitwIxMHlvBslorBgbzhXq9hy7RlPmoX4ZAA/Aq+smJtSHMZvDDEQXo
Q4OQvNks0XghUw/l5LlU0JbLu07Y/xZYn1IbfH82jX4XdsYx5D8p4l4I2w+M1Ihs
QkAk7Oovy5/+DfkWl4CEDVrvJJwvovOCHYlx5kjssw0dxukkYDAJ/dnp4Mz40R7s
Q/CP3Atz/tVzlJ/V9G13LLshSpDx5TrNX1kd92lH+RKTVOacYelou1kIQE/+ykW3
7Kt0df2+UkxOzTzLD+i1ebxCAWtvG9ggClD3iHzM3kCYVMMe40HvQ9n5aqisnLA6
9NKz6trEPv4RPROqDLTpCWonBM2DxXLhWIs+ohHxVwC2vCA3/t4s+FsPIuNFiAQ3
msLckODt6F7pjEkmrTyEqGc1OaO4xKhwwXnQXGXEOwcs8UNsh5tOLOJ3CDhtfC1b
EiVmQB8KK60XWXZ2+AtMJfrIaVUXM5NtXmKQediwQevhTb1Vk+SCz1vdEJzCKnjN
VwyJQq7gHpNE8bFMYyCrAGCwSV+GmFwbe9Hsrh3/X13h/AYYyO1TNzVPJxcrjNrG
e7nmgusxHkSpbtf8kXU2sRsk4l71wtTJDIahL4wvoWORoKVEPnuEIBlgvmL9HwPh
Jlu0zUQZk6ao/oJMu5I9ry+woNx4FrwiqKxgpnd9Aj9vxL/+aGaLtp6H9bKym3vV
tTW/l2yrVX9gLR5kQgYu3DAlNmotp5zLAxRZGZdCu2A/rvXq/QfTDOHBVWiY5+mx
bYfj5wAiEawulQJ5Ktu/bfusOJrjcurkwJurx5PqeQEzr2up4ZltahnKlqJR4ajo
0kgcF71LLlm8oNIgZPT/REtPOFJrkLJ5nQGFqYbQz30CHblYUBopekJaux5N6LSP
zvdbRzN0iqXx52+e5AzH0KFFRbl5ceTipnmeogFXoEvjuKugd2AkJLhfOZmOAeVP
CxHh8QKvup0TW24SIid1PnHeLXb+gqg4c2mvApb5jCMpzWj/cWM7aUrse1yPH5NO
lWtNUTOS94rYd92PIeaXJyZVxYXTlaIzMYsTpBHao+SbPqVlAdLpWGhCOC8rsE1G
T5H9AEBUl/iUVT2GjRjd/SJ7vgbU8VFmk5o/hDggf+EBAEIYyaAoQSI4sv43Sjmz
l1NrC25dt73yCY84jULg89Q/rZeWGbMQJndm3pPM0UBzAnULLSinPr/tooSc4HUl
TAoS5k3zHqzTJtAKMLZm3tMcRPkO/AN0lsaDnztLcOF3bJTlrY89zlMbvRZ+EQCJ
1eEgWF2/k5f1EmGy678G2WKRdfRj3UOgmwKTdyzpEJwNyjMXJgJ1HbUvFW041cuV
7z2/hTHr4sIpcCdlxTxSgjwoEl8FaW8/RSJIcYE6Kwi8SP7DzTmBZigCPCmrJMTn
cstOnYrvfDh6+cuKxv0WHNY4krV313UX8GRij82mad1ilr+EiRrAuI6DjQqX5eMM
Gtqz1GCKug6qoy5eP6Whb/lQj0WAgL+2EAXLHJM5H+Gw+qS6qp8GU1vSBy7PusaD
JTR9Ikt88kkHsyu6MvjJ3ZBmz7zZ+iyat+sotK8Vurc8l2ONysSzUAVflcP9Fjs/
DT/s6Chlgxg46UevqKqVilHTxEhid31NhS6QG9SsTAtTMS1oW1QxRH4SFzJh4bE3
kFTVGXvSyzU/D2ZyqRnBHSs2P6KvJEgwi15YTlXJfITN8ufxBST/spkaSxL59AV0
zGYVbhVYWXAlcJjPimIHFWabjIgTASa7RqBfZ822U1FJTPXVlXXRr8UHAbVndTyh
iDQCudDunamKsaAyUmekPvWy7mhu6W+Pe8U/kR0LXe/g9FRudFHyFR8Z57dZkMTq
qau5YS2A67U58FakRvROEKjCcEucmmXYkilCeGeVpObdko4Uqck8jXAd5ZYDKGve
GBsx8LWRUPQeGEtUS6BngH30D4PF4shtwVMGLGJ2clzn8ClciYe2Mj4vxy2Jireq
y2iVe4F1XM4yNaGPqo3Q2yU4nG0hzbaiPndWr1rk6oSjukzmVdiCjNnFq8hetGNH
no1ncVhm4Dh0f158mFGuRSWlaPwrKR5NsbdsTCTQbUIgRwQPUASGpPJer2s9nM/V
hcaaLj3NIRpHRFCNBeS0wX8ZXTYyHso1FG6zbCJL8WnPqrQrv8O9gPTu+hXatI8+
V7nDs3hhH2oR1WDSXtlydE3+MNkEi8TJAoOhfMEGVPawS3G+6xh+COlw26CfFpzy
/XqjRA+MMiqM8PSbt/PGpG+ZhMp2PE44Xhlh2BT/KpAuq52g9fvegl2vX32DGwnM
0AEjipB4bROB2kuVpP0mIMGojDhb7qLpx5dLW1RbrmTq22DRzedDlYPYg9zosbDS
A0JqMaxki6LUdYAATAxmQMIyJptQZed9/aJRzXnT5oZAkxNAqSVs6sUaFZEo/S0t
Ah8/RQwEqP6zmDsZZWY3RyS1yO7CW9aTQFpSd1GvlN06w0XT9DeREWw5EQwe5ZsW
XEYaDDjGkgwAVQfeO2DwT+CDLadVl/13+I6DIoGHJVLO2QUVWV7ZbGqUbS/OxRTp
OB0Kgw8Sxn0ocArktbHhzIsmN5z6hNc2f1xuG2QtwtCYlONGZgfeTNq01IWnrJs2
SuFEP07huV7YDGpnTMrNMlppwQHw2/Ze+m32vDysDKhKWpgqaQ4WfMQ6VNyzQb7P
ShG68HFvSJ9+Va4jDKsL0sN1KSkaQHdq0EEds4jwCTX+lnJU1MDqIGgJdzlJnxwk
CBcQFilzMRZ9lepjwpVvovafE7FU9qArNE5jNR4z+VLx9FwrfGEa8mQU6vL2Lv+o
k10H1yP5AWmrpWB+cJnByKyUhYh+t3rAw4vWF4m8QiFwoO52dVd0grf3tnEJqeOQ
1mBQBKmFuo+d468yh/HHACsTxykO7oxERFD5FIzxEUqLdZkSYi4AyRtxQCooS9jw
q2XZAib2KeIwbgOtb+Wa4SvdAltF5DyAsW8XNPaKkhu6D7Q2BMrVeR7c9Q3pajWA
Sc8r3fSh6WO6F25KVf8yL1ZYhfnNmAeAZI0bGYcu0pGAtCWi/Nt+FohKaSc/BhWi
aVt53yZnVw99T9WfV9RdyXZg9rdWG3iDIQ9JDYvqMsIXX+9Iqtj1BJglYnC+uHGa
iC3oolSmpRjyZGLcdhQpwOBkk1fQW2sO1dYyr5cb9gKAUJyYCqeWq1bc2ziE1Yx6
Y7aSD+aQbKXtZGJyH22vqENajEkfHIvq/Vysbpu21LTYLkdlKHsXZKNs3chB7xSA
/HjmAC++PK8IA54kzEC3OVGEZvrSjuAF5/hjU6HkmmHaCLzMOuuhVIR07jtm3e07
9gFIibfTEHyMSUyT90Tqha9X0vfVOwbiS4R0wBqVIOcsX6eVn3hsXpKv5LIswdCj
CtMnkzGK5GgdlKslID1BrA+vOKLBMJyzASVUBqRYJNL9PUfHKKowX/Zc58JO4UnR
46bosobuZ24GaXWMEZwESMXetLvL4X/yNtyC1A2n37fbboL7TAXiwBXmrBEaJ1hA
DUG//o66TW5aWHCD65lR19M7bTMhhkrjQJFVpMBmJmxdv7EmUh0YaLI5cgm94zyZ
LA+A2xkYlUXpUbT0raPF8+Ip2iF5Mf0b66HPfLfIrKVB9tjO71d9fDJUhWZYxB5C
PksNMLBP6asXb3CUNem/sfwBaeZ8QBV1WbEKQWVLiUhWrI8uO4GxL3uGxznTjwIW
TcJrX1qKmw0aXkPpm8FnaNagwGqkBYYP99RdNWQtj2+Da3gmGqdcNrfomg0z2NPv
eYwoKTIRL7QoGQcPBichjmrmgmG8IJukQVbNMlbwg/bDcntOR1eS+srlD8aX+GUg
Vtmd21VbP2HJDYPhf7biWN+p1RhKYKiufSkcXHdP4+nX2sbafxluPdWuRHYKoGVd
6ulQVjWGC6OgZpCYh1n8ODPfDu+k0EGfcsh7BFvlkvjhhjE8TeWqf75aZM98Gdog
USB+FRImyPRipyFM9rD9RwDHISLf3HeYVoSWgxjADJ5HTVRop9CeqfkxOYGUz0i9
cnYrv+eAe5RgFdd81bse9OinYsbQWafSA76LutYhSXIdBlMLndMuQPWl2vPhx3VK
tANVdhFWg7EvXnPAQB2LmSA9w0+CwO3nvQ1DGOc7ZEWDc3BZTItEdEUwATXGw+7w
xZY3Vlbelnd0yWszkLLjQp+gtFFH1ModG0rxg4dtVhRK2nI+bqAi00BrGbVr1NTm
1f5ZysLgIu7MipVHUfDZTyq3pO9qDGhuOsYnj7a5efa+S657sA4Lx5tIBc6PDHjj
jqXX/n2cV4bg+dRJjT5Vsg8mmLoN66e1CN8xDSSDf+ap/rUsKr5J1uW4peO/rmVr
lk+qa+Q40iZlRMDCnHcZgQzEc9X5wVvR0y0008ap7txUXzzu24tc6wbubY10dcBo
KF26fKFLGrYN5gcNA+PT5k5OptELVjJ2EpuHh9HGLev+qExMRVsHech141wsowJP
wzaE8iWuB7IDX1e1GCL0ZaZ/94V9EW+OsCweTpPBLYfIMlhMkaNFk8ICW2Rpa9zM
cxqBrqN2MT9hvFB0zRBvjPIkAGf/aLdn2PyNztH/TG3dEiwzDq11y1XuBZyA+qMd
qGl/nIsL9EjIMyndGyZwIF+W68+tiPmyVwXosiBw3HuyfeNSNuNXPea/XeyNaFhG
`protect end_protected