`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 34752 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
Oc4fq76CzL4QYVrEyjSlCMMV+WsDyOzrrwoms96LbjLsdp+nzf9xMERV7pGGW4zI
p0kQ+PNCaki2KMW5/5nfZMdaocLg+EBdhoKckqovguiDYYboD3NzrewoX92gL9uD
/GTZQ0JhhlaxDI++TfwmAvYKjbQLP6QV4wptQ+Fu4ufCpurgug8HDeaKNhWXcYxn
EwZ34KmhKR9uVtZtHK5lLJtkSXd272OdX+LIFQsINmTbsr1Bu8P0+Pk19uS7o5Xd
fCzOW09CqkQiieMK9OckPCuJ0rRffhjn8vOtfYsgy4a0vy9i6nDusqiB7BXKE2XJ
/MK1wDzvSELLAFGiCXhBVwHdyFghFSPYjk3YScpZAwWaUZxa/YWOec2KfD3aB455
5mOka9rFkF0ZXBWUP9T+tHv1lzupb+oB2LKJ6tSkOin7EBwEJVp4WCOb360e4dwN
g5h/JmEVksf4AXfvHgOZcg9XmjnBnPOC4dKmgQyQsz9zxdhWTnf4crwq5fv8jg7m
Mz0MMd31u0F9eRRMN2zZWfcdKE/aEbMexhsWxbR45kfRxctjscjmlxvPWJKC9dxM
/8STOh3V3K7y5PSiASn/mhnysiBshSoc3vkYkLaRQftVBY42b3runUippFCrL6lX
2FTRvirsa5DjTg3xXzfqGTVV5kSPognwuaci7mB10toslFJqUR9US2YKXX2IW10s
UWGMzYYKtJPzEF7NCo+j568otkNaWPuHGwaBpx4hI7odS9SWoVvkuZXaOAPMuzp9
OncQJ2iuCMRwQ6yGCdyTnhHnVftdzBLKfwe9XUlEmYWcl/PiQznDqIRAHPC5UL0i
I15qN1x38kkVRqqNy73mgdShiNGhiyy0KGUZOjpnCZ4Vwat9mtyQ82UWucSTYLdA
llwjS37MVrku1DSugGu60xjfgRhrsntbza76GpnSJXcD1YcmA8FLjocusg2AY0Pb
I5Uo+PeEfQQHs57MXCPj3ui4oCQFIO5HjV6eMYqENapMGDN6k8b4n+LUgqRjROu/
k9VmqNv2Qi9T05HXKGykQKCUsAaSuOJkiqo7O4hcZUQ+7TW06jmBDnXG8Yscmlq+
fWOZcZvZ8YFzH6XbgjZJfjMAx/ZmWtS2FZVUWplLceKNaURHrMjZnAfq0hUSL3ty
4iBelC4FEYYzSwLC/I2Zsoas9g4RGWN0ognjcJubv9znXyZnj1m5oApWontYTLm5
gTuxRObMjY5gV44F06ZJiYSU7F9xEaJzfOqhPK641MmiTEsnOhdLe/YnezMsbAoS
k9BU4ySbnHWPu3MXBG4e7y5pkHrBmbMD2OYaBsiEaw7+bYP3OWs+J1t/ziaiQW33
j+jAWMFjYhv6mSDE3GTfb1RkyRIOPF57RsygQENEYgj1LO9e4W1frTAm2F0XwlCx
UY41y3Mc1BqxR/cx0zILKnPJgNoeDm9jP/QjY4gsPsq9x6egCwYfB/aLhxJ8TX7T
mBrj+dgKhv4yjB/Skths3F+WPEz6j4qhpyXjwZQFSbNuqWwYzrKEu0BD6mmafvL8
C6cTeqax/UZuVvnOKjrOvCXq+Hqm0Z4I/8ak7DP6DY8JHePo236KL7bD91OYzT+q
UU8/v9WXcJTQ1cGX7yy/pp4PH9fm6xwwbW7Wq7v2wbuxtxE3O548JJ4a9X+LSE91
IGzrng1s+ZKS2IPefQVRDt8HnUpfkw4G+gXmpahnZzSlnDLAnUCCfkjS+APogM5Q
OzfDOy5yUXL5KOcvFhtDYZyJRHWrck2PTweyVbvdqVYwS2TTJOMRJuAgvzvpH4KO
5wbPQ0VZ898mq3QRXRteHcaRA8m4m+Sz+Fd1ax3SPCp2K3Ai76Nv7iqBiE/NZ3/F
7UlnZFHtq+HJIGSYhyhnWyeqB/4xvaWxekuAA9dJqaPl67YxDbwHc4ZZGtaFIUcV
xL/pk2pqZMhkQ6ESS/b9WtjNeoXPKGrxDR+8eSoks//goB5lAGHH0QT4RPmzRurP
Pf6XXX0Tbrh5rV1KSr0lh0m7mLrvTSjkzuGNGKvrjT/Fv++NyewxUH0dQ81cyxWo
deNxPIURUrimVPrZED3bj1zG0CCiw074Vf1mp8ui1mWAShLl2McKzFMj0z34lCFn
G/rMKUZlfC6UnVITDvl+LGTvWxxf+QxGtZQUUhWl/jn8tBRcq/9uxZdH7M3bONcm
yzYFdUMRxy6RNLi03DYIe/VK8kj8ld+2hPAwTqblmPoiWWEQ8e9OT+fZk82Rhrbr
iiV+FIgzmpxX5cAfQfUPfj2N0LFxiucVMsPDjyQhHV0ObifKphZAZ0QOctF5Mwyp
QDfTeHwVdcC7PFSloSfPhQXY/jFsc6V8shJe8ab96KBoq/z9rctdDMZxDFojg9Vq
5tprztUlOnEXy1cSaHIZlzrtH/BRnn6S49MmcFpG2+got1pLJERQidpvWjTwYUVt
fAM10wty7koGmkKRocEkgKEN+DuxcXGKHeLHMZyaouHZdOumduG+DvKBWYidcTK4
tamYY3SOn+70urjjAruGhfugOe+vl2DAT1AJBEeNEegG6wtiIE6toSKumANRhaCR
JZyoJWgaFhxK9UofyGGgrBV6a6UlbTkK6n81O8WRik8aq2pZqahTX4kBNPkXc+BH
0Dsx88GE0Vz/xD4sT25CZjGY/fDLusizvTROokMiSQlp/0/l1SLlTQqlZqkva4K5
vx7qTAQQMDY6svc9INY9eA+dBMsO5McVyFPEFaLRQhTc7IajjMVMpZ6e9bDuyaYI
z1TmudrSBzo0d+sZMYMhTFqP5EDPcaOJkgc1T+YCusrwFcGHnXDlmPpPbdEYkk16
D2YBNJcpg0ZdOp1P6h8pSGJXrrt5PUzBLIeV7Kjqd0g3xCLX5aF1CDJnTaS1VCZl
gmB1UmbgkV3nYf7Xj7fJl4pYPPO2B5NODfIFsHSbkUc6pNY35o5ohEbbfzHUuzvh
0xBfP/GHmvdgCUs38eFvgE36fohZw+cnvZ8QWl4OTcAnliotQQ+H9aZrjgmyIjj/
R3qS3FoSFrFtNLuu2X6QXbDMS3VsrWYBgwl3tP9EQKHmz5swOw1aEFjhz0l1Dcdl
j4Pf8xUkMYmu1/dOUkjs+piuylXlCkfe7h3QlKpiPNXxvv2pox6C8crqQexZGQd0
jErgl0naVTNgYkCbztcnNFWnEBM7XdkrhTHiIMiAhgyb7gpOf4ld3ectkH68DXIk
GGizpRF8wO0wA0VX8w8CdAiL1PHs75LFYqTgAduZJxLHVS658gw2JwwfeEcSexGG
HImq61x/CXa3O8o1Ig5UGLQq4KOMIWv9qy+71eBko5TcvlFWu37zmWyNtY233pV1
3YDDXuArHJwuqZojZYSg6dAOZcmIKxcr40ydRxiGKDLDYXxJwjQFjaYztUlnZnjU
Q+Qp2+lWguJpEXSeijvUsbSfRDrFusUpLkGvpxA56TO6m0v2AbQ85fBfoZsOiQVT
qo3Xh1sphGkbXkWRZ6gDJkMIk/H16jVKogDN2yQgMCQ62MpbhCP3L0erG/kni3cF
F7s2B5VgNBW71iDN8E+Br7EZMeEpjmqMmn6rYuMCAY19YtVh3MW+IJhThYTCBYzV
ICj0FH7J6HRpxsHb/V9U/PGSl0DkIy9mu9t/owL4dBnlonXedJCZ7E/w0nMmLRR3
5RDMGkifJEu3x5NkIeGylFozu4PsGisM0AhmedxN0VIv5L/LwJrgBuSay7qRePqk
TjuKvuL1ikiu4aXUDMXd3bhtccAxLcjaakuyzHeH7IjOU4IjNrU1vikd6eY/4Fb5
C7ZqQybcy6hGLs+Yqf7wosT544lqL9G13FJ8l8kC439mNjUhYjkRFxKaJmOcy2nN
aYC/g876ESBWi4Dk43vj/queQjvPTHwQtlU2OMOaPD5iWetMUAjpiQ2cmQGDfL6o
U1hJOgeq0bWUI5Dw4hWbmLz6bBxprI9WvWXPug12DBHE4JmTRA1s/ls5srXTNRUe
t3VG/uk+uoRd2DFcsVUjf2EbAVC+4gyip7Oj1kere6PVq8h7sYtaN+cyyTCsYqJZ
5t1NIk7EYIawJGdSLNxXLU/Pv1TraZNs7mBIOy89JQqaJlZpBvk24vtWjEthEMlD
tpYDoM0uVGRNTtS0YP/c4bLvM8a36BlrraZ8BsslPAIBRyrAlPW/aqOfUvse+9YW
SgKYRbSd/e6hRKm1Jba5cOGWbiTvBGw2BDWyc6y+AyB0KaIKn7IM5fXm9PlafH+X
2invfFTB3vq8siLH8S8CUwo7Owxyx73BQRHmTPZIJxUaHMs7n15d0xg5YpfLpBnS
xhkBM7GWWpwgB5N2xF6JJ8SkCNrUBABvreRyK9Os8rXWFM4Sjk3TvZm8jFtlBicF
l0H6/pky9P8jLGC3ir5Km08d8ULE03ANvgrbTMgFB4YJ+LmrI+R9xUeripVFnuXe
/pVygR0e81FJ+Zr7Bk4ZPjYNYHrY8f0e+v0q0RAeik8v6Xn6np+UgvEDcHRnWeeD
1kzLCJPSpjP+k3CX7SRZ0C4vgvdnD3OhsbWRx6zT6Thtkp1IbEoG/U0PGJufgEkr
t8IOdkkULIA6C8wOJYCxQNEvJgkW2Hl4qNVXR6xWQfm3uWhu8zBOJ49mIO+odsl7
1KK02KxmKgu3qvzcknJRuUP2VcUhVJ5FtjjjFny+eXGU7FKjoCSr3SI4NLSY4R6e
0oDLzmun05ADR1BQaPEOkZM0X2uVX0i3+crZYe8ST4BCcUrxRYAkQz3lQEd5vYY5
fOfKOY/G9Mgb1sdvpcPovVBlnlVkyWYDuciYch4K4elP/waJVCE//cAX7imMX9a+
eKZxV1XhaJTOiqsO6kFTBvok/WC0mq/dqUgP9OeugXH9mgXBd6VjSqbmlfyOV50j
c9OJKURsjBgB0/CMFPz6DEv9z4unrMUWZqIQEfVQJncrJ5D3y2+FDwpC3n/znMoZ
TMElU/DmBl9Av5yMzMAiljOb52dbTu/FrNrQ9bNgUF8Q2/v2OCxbmQIGpx/TTZ3O
Fz1QiTFQUMSTnGNF5orJVzuw0nyOwbSk2Pl/1JyM/K3oQPFFDZp0xV44lcwVbxdz
YZqGQB+qxNbIYbIopBW6KS/0QABwhjRfl7RsUH2capQmBHctoPrhnaZo/76E+MjW
mwsx6UBb9Y+awQbyyr4W/bnsNWfTa58bAQi6GfMUz4csOM0GmNVpgoq/dZEQgGIc
MXQD3LU2x1e+emG2+ox3t8DJ5oPVeogE0pYBaQflwz9CsHe3zg0sjJ6Anv6teSX4
bRNhPDNe3EotDhu4n8PQM3x/pmj/QiH77k5YJAx2Jnz9BGkgOITgyM93gmIdv5mB
S4GbUfM9VOwlj7P1rmnSwroLni13f6ebLZnKrEMiornCafCIQjkwXjtjM7yC7ciD
ZSWFQRytiTEuhhC/LJPVVOhA925XCW+QK0As9zhRBx2MnOV8NLa2pjPWKLvpsKry
+NGRiiSMsUzr8eY5r5yjVHjFMKrPWHI9OYLmUsqwfayPCLQVI52q70KwwKM98TUo
8GHF2T1tZBisBUeGjbQP+Uy5dNQIcOsfrsueuM1B6Ed8Skt4sw0bC4sQsbcfW/VK
EcgzcN7+NF2/Zz1UdbpxY0ehM1awHYSzsVh27PTISB36ElXN7KEtt4YboEs2C1Gg
YAnaHwdUn2a0jAv6gPWhVjO+L4GwQLIAbTR5lWWloT8N2hcSz2m0uoB1I0oswRH1
TcywOwYdA5bV2xUXXOtNTDAz7/ut9VwEeobB/6SknHfGmJP4cqWaNYoOELVDVjVK
BK6vbb6U4FDmYYtLsiEGwoie1uLDx11v+KmTc9ZfybERW+03YmgleSf5kkzpHBNj
dJW+0Iifaofb5W931c4z9ctljDdEG+zNzoGAL9cu232L9ocuTCYyRgJcOL7VqykJ
SFF2B9gmWd4Oluuh/yVWIfACVXeZbuJlV2Mwultd4vhmH2e7+ws7vk50B3Avmma2
sVyHMmmOY8JIGrria+G1dZZfsvg37RG0taA7xx/g5V8wzIJKSFHQm/jvcC28kszp
wprgwMkdsqg/9iD+VnvOG4grXTqsdLHSFREyrcgAdnog9N5PPZYZIZcfHET3hwmL
xa3bFhzRLUDtIHE3SaIhAk/OGHMi5HJ3g9vwI1tXMgnfPGJdoGu6e3+1Lp5lttlJ
yX+vQF5GZxxXJTXzjWzgjnqKTSCYGSn0jNmW4iwJSMKSxapzkW6X2OZ4PwJBpZx8
HH2LACsJuLJwxesLYz3nu7ur6UiDbCqo4y4Vb3NSJhDEN17OfUlLqf+w/ioZJtkp
S3SLCRByWeTSg/CGoI/ZFxVzBM/hsY2HnKj1Ya0ts9er4mXn8dTcYLJzX++Lwpck
cHhYMSYfzmdHohrpmRpQO+6KHXH0irGOLqMnb2WHROuGx6/LRfi+kwEzj/AvZt9u
r3Rpj+iR6PXmCJ6Mq6WIZoRSiXUbj5gqmShpgh4VT77COYPdmRfGsCFCH71DXmd+
WYNtcwkEYP/KXX/TyvrwWVEzaLT+ANfcMvJnd3XooWE6jwjxqi6CtA0A913BOOhm
WLivOctxpOvOwf9wyvi9icVF5XLKGA7aKbCfAQ1NGEvWmvdva/VkJo/SqCIArzaB
FsIXmnMaOjQZHcxqX5GSSZ88FYIxRjXRcHOi511Pb5rMDL2lSfS2A8H/F2eaw5Kv
kpPT9C4ExWEggZoX2Dp0FJTHqtFro8AvTqDm0lzBGfhK+XgSaCj6EbpHQswSURxJ
Wu8HKiutfb4RIOyCsFUyktAV5RUGRXuYwXMYCELdtclbsY4ezwkgmmtkl7BVxViF
0neVmrTNTTQQQ2pEcDMnoPJn+L1f+oE7bNr/JiZ68vUgtpm1PazPeWH5CUopfuTD
DE+5aAKAKtnx3dxXx/CySNcC5MaP4ZwXi8J+X1ePajBEjTzfZdeMFjx7CQu8SyPR
ldXDJ9LAJiR3Ark830tjRBKCIX1UNMygYSfzFs7qMF6l7283x43iVx+guB59BJmB
mDeVg9AIEAo88MQss0EVjnEU/AekEpgDxJ/dCLETIxnIVyJ2rxhVkaoMnFDx4Ktf
sm0l90ZNhmoz7CFkdI2dho8dLDfqpSPXJrxDBrY8xiEtqoBERePh2rYUwaTJVgJA
eUbiEbIeiKmdgiZZ1MNGVYQtwRxnk93ghPEJJN8ogw0rdCFjQrUcL38nFNu3dI6c
LywNXhwpKyfaU8ZIFH+6ti4Yi6wVix5t9EPo+S9HKPOle2ZC9qooPad/bqqos30R
TCYnrhpjMJGD6v0hMt+yJ6dQ8QIr1EV71h3mNBvIf/1AKD1+MoH/gVJxBv6M3g2S
jNbvFrSckWIHjGaDRSylKA4NE3LYbF3ml1w1ERznymj8ObfWMaZ0FbaKQesomnss
FYWr91GiaZPp847XguuulHBCyDfCQUMENn2rHUNLuFeSid5mn4cVln/ibfGn8QGD
CVhhFvwn5g41p+XmNtfda/U57/r13mbeN0P972dQ7riOQSEjExiYlZZmdjoyO/ko
BPUVY4jqgFFSOx9elKSDZwfgMnN/WLjzRJWyVewZnNxqafT/0tuu/ffoeLMULFmw
bNMsoA+0Sj1uBhe/998YCZHq+/RitnQcNzyGSR5dJFW0sI2vl4OiV8/rgzSyjogr
ZIKLW5GGFfIPt7P5YhbGozvOrsrw7Od6xiZ/4iNCCRS0Erg8wA3ZPfap3e3FM5j1
onl+as+/w73fyWbTZbzUruZaIzvkCj/vO0kEBeJDLoc6jyIHDFr8sWQTSEbDh3Il
QCpMObc2YND3Y8UVvngvA/+Vp2pTSPTkhsUhGe9aKghrc7UllxSGPPjnobF6MVdZ
J/ciiV0YMdxXIEcl15ArD5oYIUNaYhvojZTZMJGZyF6nmX1ypGxD3x5cahOxdQQ4
BRa6BOo64NRfdPZKeixzQFboYwcmS3bIJBL0tSSZOEZtIHDGrpIaTr8p3kjfP8Jd
j20bcZZq0UkHvvcsSwxZ6Hj0kRSZXCR93U2PUu3YFCeIVM9AlV1OHOwxTU0bhXEt
Uq7aYRt4on02IpoCfFCbVM1r1kriDJIv+8O1yw2C8OYf/hytktfA7cKZQOVTWgXt
PeXsQGeMYk+9WaFXxQbz345/Qqj22FdU053iHdA+hM15gUVFnzzzKxSrcX0Cxj4s
wyEZJ8d+aCnvgxLgoji7Wc/S2rVW8jQEQckulm0ANO8eP0A5g93ooO95B3p9EIQR
l+cvBVWubOJ3cE3y3gc4JXw/awrPoDlSAzAYE2aI/zEpT49XrnvYdXQbqYrYQe1v
YfZGbPpvukcnALy/Xtb8i60bsHid0I3HR2Li7KcNRDx4v1OaWsN25Y68A1+7zbm0
zrRBnv4955R4nEvYCEqrYEbyLoGjYxbVgkctXh0rKg8O1c/z4S87ajKKtXKHiScZ
R1LezMF4w1Vlg5MX8xenWF+67fDKzBAP5I1tJ3DPfELc5b6P3/Dq3U1W1Y9rgEWu
Gx0eE9druCWp96MHa6VOC6ENKIeBkk1spdsgMMUIKz8neAC39YbAph+EecVEwVFK
j6Do5M7NoToLlzR27FErRi1n5/OUbu+u4p5CrEC4b6T0s4AKHYh9wTgiwy3X89vV
FD/fuXZQdz8Zq/c+gG3B2gAMzA84joc5YvB2gCUZBHSRV6+2DOEH4TTsvF8XORIU
ksF5kFqLeJAmIId+zznX6i8z6Hw40tC2h1ySbmgrEnVvhXdvEYdupoXNedtQjw0j
y3Nzp0YyI+AFVqJURw7vtEEYbeTiVidpj98YgM2A9X8hmWaX5gIwtlPRyAvUsW22
nh6w51VM1pCy/51DRWncCJbKTfXibIa3wLEiA1ShQEQRgpG3+UhdEKHy5Bigf0mh
mUGyLGLqGhutExM+rPljdi/rpa/fSUTJHpak2g12OUo0QfDhLbtWWm9urqEC3Upm
l6kvgUH7NTuhTlZu3RtdL0CcemDdAOGrU0/1WQAi4AF4W7XdTaI2RhSP+iA8Ij7I
1v/utpY6I7Br1SMsLTnwiYIKBkJEr96ZuXrpo3p69p9vExoxn4hz1Az/UH7WODQH
U2303QVYVX9JmE7YzHiAQ/U2KBJtyzb9O7exWjfLeFO7ld9IHU5OiE1E1hWV8n89
DR9X2+C/8bwkQLOFzNmQM6GHPynEjmeuwNEuqGs3bXD7oYAGRN4slBlTBt3R6mYb
rVMsZkUhO5MDg5tUDN0GBFQp5+agS2mLtJoAwwRqer1Qje554uKu+4wiw889plS5
JzduaYmjA6hdLgBIl7bDyrzGl9dyYQ1STQ4Cl8/ZnliXzG/sLYjQ3vwPEYuYzTxc
b7B4WMKqy89qOMcvNF2v2Wd0iy6Gv+2JSDje6MZVr9yVuEngUEN/CGkk3WR8hJ2N
FCLzhGSIZ6rmDRjeE0sAeopB+IOdPHg/S91GjbKOBUYf7OWUH6P25zsHR+cBaLmw
4Yfxw/R3oXRbavwEh7aOE9nBhg5JocpkMZJk4iVy6CEgN9eWkuzrbvnvDuF8wt33
APcnmyPJRTyhyJarYuVmYg1ZM2fHZLHGUPSEwGvGcPOV4jBObeZjJ6mtgHddaAgE
1Ug5x3RE2utxyAp6Sb9i9ryw21gFUwsPnCd1x8s4my9M+dh2Fnh7de1JkfVKxzjV
SA5PkcsXQKdDjkBs3sSrhezYSnCd358GSBuDqpQkucDn/XJy4sCw9s1DvJNXM7CM
o8Vk9ouFNmmXJXuuQMgWMi2ixoflnmLB/iYP+qUGvuhkHXHYso6kFgZGAaKim/er
G4Z6b3PU6g21OEJo8EmMh/Mosobfn1hJiefcZzyNREE7NJnAD8dUTSugS0fzzBOm
jz86N5tv5kH1y8DcHxbDMWkonWx42lhfNjSCtotDBojqTNLNTzYD9Eo50mnM8tiv
ItQ4lqKjLxd7UZieK+qV5LJAD+WJNvoNN+c/eET+RqfxEeQ5D5WMwJqPjZJ8XrpD
IphS1rmrGCQ7j8KZlpTHMRwQ0k685+y5IxfEH9KKBNU1X2kXzKHefHwUsIpz8qC6
NJL42FXN2KoAFchtA8VwURZeLOFI1iqmnnjnwoxC49rrBuc+1gTZ++mbf277K68d
abAGjfIMolV6a5G91ZshdqIVG9qQKKVwZTnlZOJkRBMdA9a7vxcN+H+XbfuadXZ4
Fo85iLKc4qycYnusKeoY3OYJX9i7c1o3XvbWMRjA3wLytu7KC5wYdXTP0dKO6nfp
bVJ5AYdWk4sfdxHVRE4djIgUKq6aGRd67uBAvHWDHK//v61dCi53a1Hss1cKaWyp
Xc/3/Q/7v162BhiQ/7Vb+YisX/GLnvs6lJ2KPXC+hCPi3GVWqNQGtTzewSPIK5yT
W9/ZqpwpbOPH0Qwml3v94Dfku5Ir4hdyhOSk1cRvCF7Iv3350jnqImxWqzpUeFTz
1Fb+yd4aOAzPDNojOAa8RT34cU+ZdDtqrVOxk2t/bfT7iQbPh6UcUJVcWO7NL2ia
leCHopG4m4VsfMbpHMI38FEj/HUrumCt/8Ds5Kx5lWqjprzlNQY5N0LURYsxg6+w
n3/8zaTj8gLO21KVcUDkzCVH7Wx2yBbNqbRCtIjN8BHgH2DmrAE52AmgBV7EXjd9
rbRpLZ5o7MF8T8ZHy2JxmXragDPvlrsku41fNu58BCJ1UuYFksaJtjuwz7bCXCyN
nqdcKUHe3f2z7aDErMH82LIaByEC4vp35j5P6vRa7ZJKPNXHB9QIlGsR0qY4eDQ7
SADBp69NLr8mvd9/fj5T3eqETUiCT/LTO88eqJ1vMozU9TjhiHLwopEPnWWBYzMK
0KsUpemXUIlz7Z9TptVm773SVcYz0YATPmlsn4A2WaKxe7GyQLCoHkcl4BTvWjQW
OfJ7nusZ84EkclpPPOb18kW0cj1iYuOnX2klRZ5APoB6I/8N0vUWK3ueK4elz+Q7
mHsF8TuM0KdT+IVj8KanvotAJ6lGlji0wKMLXVAcX8OfhrlP1/aMdIbtVZBusjCp
j5Olg+akrThNJlPpoVCIFdUqbPuOG8VxaqlQS8KxpISPL5c12oz6gzSlPJBZ5iaz
IiWlZdQy4E2+owq8ugZYWT2/RokOS+zcgC/0l7L1X38EeaXeMB8zwN03bbBdIFFN
2T7lGz8dSnhcoD6s9O07mjoh8hfwE8n0Oi6PIgAlCQa6hXJMQXsde0EG6PV2hjyj
1ZBPwro2aBTlhJdj/5v2HAn8n//v+Sf3ZeYKi+TgCbtkElCccAO7PNm+u6naEZIC
upw+pRU6SI1yBkphcvr+ICIx+N9o7DDUVpNnhwyI61hbMtC4W8vqv+zNDg8hdu+D
0oCA4sBoYu314z8Wf2kO4bj8JBQbsYVoBPjNxfXkYdDAGAnHN5xRhAuRJI1zA2tX
u1KFMlLR47UvKFrquVjRZs5f/BFTrWmN93Vsk6Xg3XjfE0Q9LsuAR62+Sw2bUnzA
DccqbM3diAFjAc0EoQuZ7AKsrdVMgyi8WWRMoapHUT6bkiTUffk95PAC4n0lGivc
xamjGSQtTmOhNHU870G4PZhG6lFGOFem+T90JHHr/0pVTWnWFpTBBnCvWSy4wy4c
fGch6d4I7roxWYeb519KDZWQ4zyGuVB+aAoHd8CW5tghpP4XOKIcN1TZE7u6uyMT
4yKbzl3qeh4uMPIx7DKc8yp47DOKKzlBfVGCFapUZvoFBtN3ECYB6nQqc6U1bAEd
UF/Q1szYCsV2UGw64uWYYUo0Wdh7kTH2uzO75ZLJCf2BkrsyJtbBP2BF2I19ERoe
IiebbgxzH4seYlkcLpnQO5UvEQ3Hc1DIlE8PiS33dlhEmAFp5xBiciUpspo81iLs
hSYbCqTzJbykOr90b24BB/qOGASlKvVXzEGn5lKPx7u+grjZniIfzc6UgDB+9G0Z
6lpBoYo+SXVmjgADrhJW2USgul9z16NxyZeSGLuNp1Isg4DxyC51p3DFxefRZ7TL
hL2H7E1vGdoa1RFDGsDyERO9g38YcIXa/HfGKQzhn/3gCg60IalVatbY6/juwQ04
LIQevoduJ6aATcS++kQQ1yZOSLsPWJiJTWdfTEvjPF8ESeVnwdiXfUZovP9Q+oGg
+bKiaDHwoFkuqrhqpM4+dXoFMF6X/jHGhJCJ1IKZXriCGE5+Q2HPyf0XRdwOYgC8
5aOyeJNkFabn03xAdvrVOC6/BE1MjPwnyHacCgTsfC3eer+m3RIdDlQ1G9gFJxyR
kT2tyxqXPXugq4wpodlM++Ym6TCJLAI+KynokwpxwDgqA+6J2PwC7OxjK4S/jEla
dtclO7g0bIT+XadW9ZT+DcrNtAAeXY9RFSS5K0R5OPjT55lfYcC7nrsVt+8knk3Z
VTy1coLpNeCHwJDzMqcSoKKT0mL7r57BhdfigxjDx20UKCbFa4xbw53Ipe0JGjrb
HbQ7NSIPwgVnV5wsk+YSTTweWsyzQvoACmkfcdF7/USu5XGaqGelReJlGg8qbXBz
KuVUXEuTSzuB6/B/TBXPT2a583Ik2248E1bkJ/7QPXT0T/J3+ppbGtjdrQODbnYx
hwIWDB2M/bIRcA5JlG2/1QX3mtc+/l0/OGlkc2c0lg0X8IS/ph2zVrVdtczVtmWL
pJOgyHrf8qKhbai+gMMlcW0K9Lqm8iavKl03tUZpuCqECI2LzNUjhdPqAwAy+BPC
SJE9ZmrjfeNA7wJdzUZvAR99jbutSfTMIJeFJlyqYx3fnwqZKBAmAvtccAKDMro5
25C9ag3910Ssvhh48uOyGDBXw0PNBUzWeIbMYPXiLN04deL+6ExEFeT7u+3dnOER
09fOEj1FnTn3XH7g64aFpEtii1yjxlR9DxgkQBZU1eaim6y4yiU8mw34Up1khDrO
Y37t1RemGvsXUEv2CkR8Jm2Q4ynFfZDrfRCsKMjQStqH7I7KnUagSTAhnSKPUoXO
Mjcni1EUXR1ksF8SRg7RLX9tCNOwthhRh8T5AsMpjMB1cmNL1qEeBT6ln9EvWiJ1
L89avZWU+GWp9Lk3gvKT/uLEBdQnFDqjxEodxzon5A2MWb41gAwBfSSoYu0UqHhg
vj/2DRzDzKnCXUcfQTdjyY5TQAtN4sABZLDmD77d9ZUgqXLlAv59Yio3Wr/2HpU/
n78cpg79yPfnlt8cLuNjwuqP6HeBZ+cvd+iUDspw/YX4uxkVFzYTFr5NA+7jXKne
siF4g+e2T1Ie+7H5GfytYsOzsda7uKixk6fWZbrBZ9TasnI3WCEHae53UbNoQNhL
2GplvMxcAD1xqbhGkml0G3G6yj2aKu6MLw51/+dfDahsOyq0VLUol+2vNSo7gLAM
cGXAm9KwhJxl4QyLtts2DoQope6cRW2XrUlwMs5rqobFCjqkHQBKmWSyV7v9nLn0
SAe9kFwqiT1AYLduFjclRMHncK3/eIZGsEqBmdsmC99/jt0xOfC/H3ATdGngNjgk
ZNjdmnqVzLJzmdxOA0CXvSUf/iH5G6WWDiGFbMEx1sjMq7aE5YnIdciGy5Iqy1U9
WRHdBS3TbK1TXrxY86NaRaKhc2GduZHmabUIuU4dSBXS4uxb1UWisTNWz5nExJ0J
magrdvmJS2qcyVc5k6fRQ3FrG0y5av1pZ4Nd/HD7GPtgXGXqL9dwjBn+mH4XQYJf
AS4KvPXrMKjYS7j0Fcu3wf7BjXzo+f3C06NdxYLxxKbbepVrRtcJUt+nZoAfWwP0
YCeiWundKv4xrDV24KrfgOvVPRrs6DFu5XtLooU2jafr601EQQ0gvWs1W8K6cttg
Sr9GrKQBB1D+ASxrZMj4KHXBUTvjmvJboSeAGsXMacQv2pbBe1LnCxBfQDB9n83M
pHgOV16mpxk26rrX8pYxH8B8u8AxxTxEcqzy0RgeyEeAt1WMMxycyRNYH0CmTVoi
kf318Xz5kwB1iRQK1vVC8UzqytCuAQCrf5/6cmSsZ8jVmxeZGvhMQPBpfx9tzsm/
wsv47H2dt2Am2O7y4Cnarogq799yoLV4wszTRuFZWBYwpSWQcTaW6SYUT+uugmuq
2OXuZaJLhZe+Q1iNLA5LBVmqe6VqeGr585Do/I1XKtio+VYpDMdKmuACDkBxHkTe
IKS8WZw1ijdlLP9WQdm46/L0FMppAfqGoBu00myUyMV+O5X5LMnDDFtwhwTmYc7b
kuLZjkq+iYRwAjNfSwqrkWInKXZfteKFUU/+BH6crPzmvmlYyyE6qA7jO+ONpFB0
KwPjJ5HYLy2Hohzyv/MH3Qk9Y+EB3/8vhwfSJhTySIH0fAT76gCdfZ+PA79WndBs
W9gKhgJuQJWzKNzB4y2saoAm30pnLFPA8PJhc3uYV8m4GPdKZTnAHTmVuNcZg6VQ
QseoqjqE78WPatq6ri5sN6qbGfiyRGoRuaImrsdUvlJUZ5tr0qkgf4Pqcy3asFD+
l1XrLOYu+xxfUjEprZ6DUjxP3VIAk5rS7W4+ftKNqXjUxz19uujQcYOwRVod3njo
4WOsfmyf+FZHaMSi7ETpzeMkvy5t01AHVQDBcJNyENOrJ+mLPvR43aTc+GuSyXQf
WBiitZV7vvp5+HVN4Xx7yxW6N5LPkjQqz5u0TUbW+1KKIIgrO8Q+IcP5H97/fVfF
ETOwAGwjH/EPxAebVPbrYjce9Qp0aU1kuwUWGoAQQHe1nE2a6Ju7s4o1n+wlf1gA
8mgZ50zQ6Y6BBAbZbp7piJb1XaO60ZP2iVSYuTOkmALU5hvnGPkJlU4EQXGQXQYZ
u1fWIZ+Uvi8AN0kSTzsnIJmvn7akW23KbqrY/SDdwjZiQw3yq0hZhnXv9xTYVlN2
QZT9sowon9N/8yxxemTmvzozZAvO0E869ULw/RPIemjJhcLCks2RoWo5TvU6V7y2
8hnR2COztTvy4cc+yRWVE1UemB4rqcaWZ3AjzFULWiT9sR72GgsMzqjZMM9kvFYm
f3h6m0TDE7xgjMxopMmacnC4yVmqXhUEcsY/+4ed7MwJOLEJTL9PH49cGHbIYDpt
j4FQ5KjTH2jBZNlCkVc5aG53gtO1oimPFVWxv28nQ9Gmwv4mKQ/o51VOiE9lJX9I
5Ks2+FkYoro3Xc3zbNuXxYbqyqe+7mXZ9YQvMNhG2wJ4xTIHSjCTaLiaQdFUWRsj
Z8/1r1YQSe4CuC1phmiMQKIbgIDcPMrFT6WFgzwU4xydMhPjzLl+mLKtYpQtg40O
yZoYRBzYOfBeVL5//BkpfweSB2xIwV/tUPwsQhA9lUHGpoheJXD07zM6oY9QzISg
dENHpusXdbEMunVch00V8z6+i6xFPPFixp+UMI0Dfgt8PDBMWmaq603km84/Edzn
vfabf+rU68dlBu+MQFAWvmPjt8PIoL+VJ2FHeqpXLCudOAcpfrZxuLTSjTjxwfs1
txDUUZ+yBysMqR2MXy+g6z+WGjvtMYcXrdvsSZ5pXVTUwEjkUPrgayJIqsILXefr
PzeYfDxNmIhy2hmljXGuZKbDfAZ45iLzob+gFGKsN5jVJWv2gX+yZEq/vFlWFx4+
3T2+VKfsgAieVRVQdRO54uGszRO0wx41201R8flWFzUQsy0/A5S5+mKzct6KNCci
3lRCbntpcK2l/jwCkupBrlRJQv9Mgl3J6MynJMyJtG9eYT1Rllr6uPDaXAuK19BL
9vUZcVTDvoSrfDB00tMOtWp5+e2THrpiqO6XciiINIoQAR6bUyDUsjbANHEuxM05
US+cmiStA58W94LcT3YjzX+j8upGYabrvqM5vbr5Klk4DTcMQu33kxdOuuHWOVww
OJYmc2HghmDtdRmQTPW5gLlifqPEoBXpIwSO9Ooksmkh2dD0G7E/PNgKP1wNFMRx
JkihF3E4WFNHNwNJTQH/q8XNVvNJYORSwZeqhlqc/U9E5hAvHYvTcTXV9OBIeHN8
U7AlW+c+0IHAMTPIEHv5w9Btg/Bl3NavKpWYnHh16iAEaNr/1B38QlX2dH9sQvo1
H4G1d5xoISDXEnZvgHyuHPEV68KC5nYDALIM0wHdG0TOzB96F5RX1AnOPkg/BnTv
5xuTBRmPFkKTKqnZtWib8Y/6A1dn67z3gP7Q1s5dBg+O/NTHgxqBwJZ7+ipRAtcy
y8IBBd0uATGXMd8ZnRagUkivwHgvHNnrGxWtChDLVAxkIDeF59GtTwyg3kBBq3ZE
T2dUSWOuQRczsgIViiIFIhjrX4TS0EVv/qqKhwNM1nBjNPPn635gCA0szeDQeCFb
tHwFCbuS1Qh03EQudhic4UahEtK85gZw2EhB4HgC5bB3DFkMYnO2aSPrMztAv115
F/qO7RIzS/o1YkxU21IMHVc9tBrIFU1Tc08CztqgOJFHGVH1PmkXv1KCM+eWEqHO
m6dSf17lz6IZr5/QxH7J54W09AZxuSggHo28wno2WQRKefOjooOQtAR03Zb0tPem
T+QKQ53HUn/PqphEsbr3lDEOCa9qgBs1N9TasVIv56KCjH+XkU5CLoJiS6TadkGr
bnYXNJ9c1nLMdkCrfNw9Tp3/XtmfdQBB4uRtQFFyvOYTl/gRijf2PDdTg3UKwyLr
1/fzSlRXRcwJMBMLWY+22BC2TPO0l3+0qDNY1upEE3ZPLVAbkYZTL3uc2EtbY3ZE
R43VnXTVksooVQZ44qEFyTKP4RZhiQRLtOEbKAjAltKTA1F1E+B/wO4/dXGQU91w
nOmo7UiyniwKsAuR6w/BFBHCMQE3x+SDtezyTi9dJ2BYodl+E4qLYng4raO114ta
waCUKvBIxvNXszvPNbfaTmBjdn66rhZG/fmMBUj2ltq3rP2N/xwD22WxHz4F0poh
hQHFlo0sKfzv3sXIO79C6NwDnXp7jIbqIkVa/U3X7xb+RdefvnUs03239ATB25of
DO9xRY2pfs9wy7qnCFNM/lpKT4meKnpb6bk+7kmggxgTngwP1iIFJIxzMOD19IxX
6x1z0i95fx/wGiv+A7gB2R1I/T3ZBQlxJZpL9rt6razlP9QOx8q/RD8f+vqeVUam
BFwt74l8t6Bre4XqV/wGA0OznO91sbFiK9qrZXNVcp56yGYgrcHSwamOjtief9pa
4MXAMEYIHk/w0rwjM+vVgftOlMaFF+zZMgfZ8CvkjLDxvAVCmsMU3lUjH/6lnSzs
UERpwz+nVaFu0KbGIKFHT/XkGytJuTy5++oW68pS+NuQydSXBSEMqnFXYJ+RVw+I
0ytiMkV7+yA60zLIGJy5FmJfqwKNqr8k/qWxtjT8CKo6EDM8KmZs1EtHWFemYS/Q
01LkJ82rTqtaXIcgNMSSVlq2Vdw0MDZG8H9mnwxhzN6aNC9thOHTnszl+rX68bc0
t4iD7eJmVNbir2fueCu6cUQm31jUHUNV7aBYBA3mt9oa3/DYeGvwdyrsnODvCyn9
ctsOmH7w72wQ3l+QcJzVEDn7cacOtWf8CEcCOMuyjA+3BA6893yuPCG2dFazHMFR
OKaOrnELf85E/HS8XQuZFyvInM8Fpd6x0/WVbPcRPB31WEHwgdBS6cD3B4pBGRIl
ll88ZClR/yksIOXHD8sR3N6VM3cCQOoIa8jpsYgGgrewdHavWTrXT1Wo677YDj8R
pTWI29Jyg0fahSVAgnNBL74vvhVWCTNXEEdWmDG5bOEOsuhuu4jdxoD3Di6smZpv
k+IpO6P9SMHRi2Utv00lGWCNrbb/ngeCznwwBgcxhim6O+AjTqbYcgb6XrYQkC3d
RbNdZeENUAqoOsQE5qD3cOEFVhGtVhM2aC04JDMEgka1MoTFzHAeFtQB/hpHIwd1
arqHs8k5EDoD3gAAJfUu41Omg8qChybQA4JluVf+QXkK90ld0RcT6IdKvIKYeWEb
clEF0TmcWtAVaLGiLEVJHoVKjbY9B+CsvqzcjdaU4AOjs9MlJ6TBldSF40vhp4Nm
nwrD7urUPewMI7k3tez6aHTwQDXMmSfJnxDLhauqmySALtrzTFrSA4AbwaR8VkyP
ANyaSUYji2PpXvGE77tmnfz6sBjVYAde6sK4rnvTH8U/pLS2GpsyDxBGo6vNh1Yn
9i4hN2Fa4Lzn9T/8uxE+SJnfLAZn9Dp8pFQxzKcprp0F7kMtzxWrn97t9d3G6uN4
9zOzBj0QG07rMANOYE8WZ8Uo4ylt+J0KqEGY1N7hs7UGZOfi14igjKsFRn43hhh8
zs195MphpiY+eAEp2yhhzoZu6N0vSfzmiLPkHVZ8uOQ/X3zY9XcS133FhHJRbf4l
3c8ncBPx92JLtC+28HZmc7zXi0cfcBxdPY1kVZ2dkZMeRQqPZYqTS6Bk+U+i4fPZ
f4N81N6eiB6qG6QLUY25qZ3eCw08Uin6uBfgBcEqG1Ubr87ANVzeRCtPFfk6/rKk
WqVfTOyaxnMN9U5bMxzAK/R0fMHk4bSnrE+ggurfCHxpzl7WxwKR9QuD9KT6Ex4j
c3hvcmVKXrjUBl86gH3nQ63dNF9TvRw28wfRu3r0YlYo37KnOyknZWek9R5IdPyr
Z9FL0dYmM/dOpYmsD7XTciEO5v31tjqnC2CnnPf8F5Z/yRSDUzfnIMb4Cr4sxFNz
5PyXgRiQ5E36O9v0bps96TOgMQJ+PbU5jPSqkI1tH3Yn7XVFjbmZcqfohdS8YpRR
TY3wczAI+JHBPducEW6YBupokdzhSBM1vs9H/tMVuFOsCFcfQhLIITu0ryfwrDsL
IPZr3QjXlvWCpHnkM8JXHNsgfoiVje4U2+wvV7fDfMrcyN2sUzJCWwk7Bqcncd25
zDlyEwWzJX3ix/uL1SVJYdJ5onZ+s5lNM7UmOGfPqfJ4JKDDfU3Fy0nRvpkDsBPm
HezJ75x5QhE66SZLs93YOR8DsTPLvR886Ixf454Geu8GBqOErGYiPchId88t3bEh
rAPNRQqkk92bi4YPydJ6h/He22IPZhE25PXww8Fc2ufNz1tnyVjLWdz3nmmp77bS
46i8dXY/wQyZNUXpk+J6QyXOmr2PkvlxTUhg7m4fN9J7nQKROg6KcYrG3tVbvIS8
zfCG/KzlxCr7Cn4bHGGkbMh75J/tolPW/fMSCaq5W8w3JgIXjuOr7SievqpiTNq7
XkA5dyOtfQn8Ix8d8I5sT6QQZDxozEZ6YNRlJ85vHFVB0uTQFuOQLttYYpKaSZR7
JYDCiBZsTdj/pfx0V9yGznqDyTCUMI6GCdBP1OWMk62Qjv/wJfpQ2lEjv37QJsmH
lRUeBhzGvtiRzMvULLF626fDyKRU7TXjcWY/1CYOCKCCsqzbCEknp3qZdb5ehRcR
XUtlq9i105iGRBgaxpuIoyHwsjH75zFeXO6SSBzlccV3VLTo5DpHhzti2ZkUJlmW
pS/0ZeEuvtpa/xwZkMLk2BVEBgIr2fkXMeilHbPP/a5LMJZYrx20p04RO3MN5Vil
ntepNGEcfFvaVFZewAmwWsaCi3zca7aAZCXvsr7Kg3IqOgKOdb6xYtWpRyjN4nyl
s3CFO+XntcHdAhzUsWl4mc8z/jrdIelaLhmKhVtqvKK2bmSdEj7SzZI/iKqEhRPp
HPgfs9nsBMdBy7KC6tiVlFE8bXtPw0PrkuCMwFnDGH1Hsdr4naWO+M0ZU317Wh1A
oxAwMzig6hH5OHxOei174Qi5YrwKbMCHnxe12/slxhYL0mlElqNc5+MeqigUv9v3
ny55gKht7a4BIP4bINeR3zVAPoB98ZfCliWOFr70suoNOogUn6TffpYMZ/CulTqt
dX1n4oZmoBQNZRcfNctzte+NGH619G5rOj/7heTak2ue5ApqsNSeRIcZS1bl+YzB
HDATHlW6foh6mzJ0gF0wbQ7wAwmsef3QxWBY4XRRxg/CAYw1fPjEpp60PptWEqlt
NKkw4YU94m9s/oh9H654uHbbFbN6/I7YJn+OTNtt6OAQMx6mOhE7qEyQdunhMHpK
gZ1s7+L0iCI3qONEjj6KLVbHVJlmg3Ra3T07yHCm0F9XJ+2rsc5PKifINSS1GOOy
gsgBAY/20QaqXnBI/1qkbvCX+8nAy4NgS1olY5Ouq0mbnySOJnFtbru3qqe2GD9e
IQLkNEb+nDW7lE4CFG8lBtMklMv5j7GgUTVrm4vJJ7+xpbRVH7mZQJNV2ssqourh
Sl/FeUtkDoblFcFZJx/bxdKHw5JXgF6rhCoNHij9Yifdj4X08cNgf9M3A4S81joN
xMFi10urT2yz9rTQzhYpbxKlQOkjsxvuv1BncMx/kMzZFK6LFKFaddvNgvMXsRiC
HcL3J8isofoMDy0D0RidhGvWLWYxxH97UWYT9Xtmne5kOr0S+pjqngoBDZRoeBXW
0Q0/Web4D6vUXDxi8jYkC59arR8X6jnCIJ5nvxHPjDj4jH/IKN2vL0TM1gspFvgA
8JIlPS6RH8YO+1KzpHQ4bSREO16IWRx6dnze/EbSoQJnIIpsUaXr3sTVffCwxzr3
NYij13arqhHlFfD8YACTxZ6XScAbsPQhERkPO9+k+tN2Tn2Hukvv6zyVmmp5pG9g
3tqs1/BemhM8Z5I78RnhO3BvhL2N9oZgpiwax4xnbNIil4VwS4ttBUTCpK04yKji
JT+G1MZVwys8r81iNr3Iq88pZTcFhSM1vr8kvt0YBBLVqfsC0EkiWKYRecWnGRN7
wkhmPekogv/TBmCbiWTU8/p7vnjgW6sDTEksMY3EdCMNw5+IODOObYlYIDcz71+N
wnj1gdgbwKSR0WSJ5RuycEX5YMXj5Yv8vH0Aop11HCDu0vJd0+vj3jZOnTPSR//p
plhQBTiaziALPzYeXaKnWIiaS5SgA4YhuLaiwPZs4DMLPLVaWc+wSY+DxXmOQ3R0
dx6Sk/MAO//TLryerkwqFEfQ+WhMJWnGVEgQm+eFwS0q4s4qTnR0AWOZZHrdz2nO
uumgXpkuy8qyQ355awlCGlyUzzYYkqF3GRjyPlBSgoydyBdriuLk+8k1qg0xPPkx
sORduujaf7nCpUWDlg7wBE2hy4lMd7MPHhmxs278Ot1l+LsCbNPNsLNNjB52x0wQ
aralvOYKDtysBosxJl3D7FFUsq24YuH+ScV7cPzb1VGJNCCXgU92SzPGeY2dvWh0
tRobaremjVkUIcNZBKT0tIC+iH2iIDvwDDaoRWg6pPlwJQ+8GhwTV+0ll1lv4n6L
La41zQsiLDLOIhetW/a/qOuFcsixFdunF1I+1LYpIHs4qZWVV461cDNcNFBwt+r1
41rQt+n4cFpan4pWPpDEF6qUkOTk2BGkvguOUPiOl4IuCBsC/0p2y0Mw77UJkizH
eOzO23AeO3lt487BsYTHlG9zQ0DL0fycna3GMhlZN0bBjIQAOEFAcTxwXwOWbFRH
Pxj1FfILIsiaFw3wVPxLGt6chFcdFbnSK6QlVCbo5ZNac/D+F8o87fGVSdvL3z/n
Rpiiv/XRjzhQm7Gp6/BVX6yC4Ytn2qoLE8zTablAM5zD0yauvD7bHNe2wynTYA6k
Qdh3cGAZsbjZejdekRGfqPwh1SzRT42QpHMFaphB13lq9G2cKwjzSF5xrfYB53It
raekGKfWH/ih7LTEuywpMPTO598XqNwsGiYPA0jfgOEgEC/PnSi6l7pd+zwaBD7Q
Nixl4OR05yLCN+lfTmtLdp92Vi00sMNpG+ujh1aAFsd6Xp0C6cQaC/DJSI3/RZZG
oBmT1bCeXcm9e1Wp01qmmhKuo+r2ymqQl+mBBL/zksSmZd+qpNz+OEOlaYtsOiu3
Zm5WVrJsuaVbkzMgBgeF0/TZbxndVQoibEpFbouCmbEhyNLhcb0CMSaEMVEq9/lm
bb3SQ3dlPAg728hoGXX9jy6mC6MzX9WLCxCgwV1WdsDeMj9wnCDh7YAmzElINGf/
9yc+RTWY+scte2LxyqEVbKASxdqbaxo15YK1wP+PQFwYAzcBWNsgnqY/bweM25BY
EVD6ladIbNym0AB2XkoUgb19upv9qbxPVTVzIpO7uhbTgUnKms3M9/wK2o2XG2IF
cdnRJOAnm/AfdCs9pYBdLgjgVFo/P7yNvlJ2Abjvif+vOkezbg+ObkGQ4DdGCIYS
6u9LyoObuUHa1QzOXHU7g9ihTpX4OjtMewfO2tVsio+6+N19SOZcKBUzbmEosX+N
rX+8GHkF0YlDXW8VCsFC0WduOuV/dvX5NFBZODUvwlac/OVdiQ198BjD6yqef+P/
uxnB2gxOMOxuJJ3QrJiBxRRq8+9XWbkVUJNZV5jqvrynlvoScFkfrLoBdZDzbPoi
fZZSYlPqxcfHgWJewbM98KU8Q3i8oMxqZHNml+skTVqGRgc1ZiGqYSynrvcLRo2V
yk/GnDWeRRVusnHAMCWniopm3fPibxut6bv4NEXXxNoA3oFosPRJbbmcCcYnTctu
qXrKD9h34qygrB1sCRDNxkuj5lALgwfuKTWZE8Ip1A9dsrTQMUoccQ7dmQScGMzN
CxC4E9SlAx86TJ51N+Y6hzXQDt0VeNKEZmvBb1Ix5PucHuKlLGZVye+ZP94AAPEv
JC88IOasoPwSrIqa9lWMetCnj5PpAp6K4F1BiGkzFFACK4K8cHBXne8wtbGLACdE
8nwSyrWHZHRmGggpQmHZ7dc+1zBtaiW2TqRBdYX+8A/umM1NNpIQvxF3/aT6gHLb
8rTUcCS14su5TbcLSlkP7rJjP+KiLE3Au/TsqR7JHvw4jL8WZsJeRnBQnQ51NfFZ
imobrFLqy2LLKYTCE7RZZvOeGQrZ9HfmOQ8yqwLKqAzWwu68jJoISaGbF1wk/1em
IGKNmshk2/4xLIq+D19flHlWazdfF+oJbjpug+OBfhIglgFeauXGggcYlicuZ4/I
D3MV6h2TbH37I4XlbVUJ2uIsTqningFzVQo5z1gRxvK/T++HErxXyFBLg4ZqE23B
Cx6C3lq+1fIRsGAup4fpI5CG0BoLwvSHfsOFzTCjFmVE0g+RcKImRX1KozVg36ZC
GU8AJt9qTTrEWMaQ/jtGHJbOTFW/TMWtgP9LCAgV4e2XWnCtCS9hFlpRD2uqA4SW
DdIfZw5NLvPpeoUBci8K0866uiefGxEDjXRz65Mbhrs/zg56IvIA30xtIKV1BLh7
1Rei3bOzWYiwJJlXRVGxfjtT6KEhRTUQRRKAV50fSLtjDp2bQi9ocL3TQpFB2L8J
PXscJ7obHtR5hDoMBEHiRdmUQmUQgcFpCjpQ5m2e5yH6031IoCT+5F1mjhk8LttF
BUZM3dxtJZDcHR4ximcN1fKr4ezKnll8RvK7KIgUaE4ElDnNX9S6F9PKZzjWlqYn
eyn0dsQab1YnI7Fhxbuaj/xJG7pe/6tdxZLW+JblucDQ6CMMV/pNtpS9Sn+7zd3A
5ZhOm+ldrKOZ9VEow9+LiM4rGmyQq1vp/VA4RDplQwgXb1j+rtgiCcBmpWEwKPwa
v4CElv+9bdQ1FPFC30b6wSmBA8mxcu7+elRDn11xqVk96QI4DBDS0A12KMpjT75w
AjfP2tyLXJZFp94mkP/Ib9xL9sr2MPQDW1ijGHo3Z3XJdPxA1EXtNyrYidOx4JC0
PhkjU//0usf1k37sCQq31NH6g0d0MHDLXjCkUV1eq9+q4Xw2DQjgZAeomS1a+MRJ
NHlJX7jw//wH8O0IosDRasCn4fBsOJCy4VAhFj9cFQYAU8IHM+HcDOHUXg8i09Fk
/G8vCQziOyShYGVgz+AqfeLKX0/gP0/0vVfFRJROXyQktt34xHxinvEraOU9TzSS
gt+gs0ZHjLk5paVMY9oys6RF+SIFOuonfZFwVflBQsSZVGqMqjNoljS2tkGzmmRX
erPdY3jLrozGKSqcwuQdaXxSnhwbwJOpTsLoN2jNfs4OSv8V8nvww0/hnSKh/k2X
4HKr0zgZigmOkPsGtfmKhQQBxzbJUx52jXNv5Yld+v9w+5AJWYzSvKFrmqLtIWAp
MOYHbJ4apYrkOBprWTLm32Bz1LYodYxhkSvDgN31eBzlt/NP0p+EkLXgiwZnwN9Q
PvgdGRmf5YVDM8GT6cz/p7F29pIK0DD95y85sO2RBNOa7xjyI9r+xPDdw9qq9ywJ
XGGMqiH5SKlkuDfQHVcI4wl2MjNK8sGTqXHqku2fP3Ztr6XXzI9bAPsxlbVZCi47
K1XwGU3CmZMoaHeHZgeU1zc7u/ClmbXaK0mtl6NmSWlI/xLPQhL7b6wldBfyTmde
PKVFmVJc2IAollMCTG7an/X1I4cWlsgC3ZwIO4gxEzpvyIdaIYb+UcjMQ1/0qDHm
sx0p/iy16WGtv4yhaBSslW4+rX1MJAXlIBZ4kbNzXkTGEtxT1WwVuUoBi2s3mAQ1
Ncn6rPvn7dGZdYVQlMk6gV+0MYSKgWLymbdVSyWlhyUztuXkLi91OydKViR48+oG
bJMv2e3gAlhU/tjY+3hMWAXml4dGQOwj8fXF44Qd0wAA2+A1dvhF7ylUC4p+O0Uq
O+Zktc+zzUfoFezPMMYUdjUuDfyU1g9t/6+cN84slo+HRM/MwGLWzrsFL+gIQGu4
qp2YDJjWTfDR/H3POgUVKhixvfAHGYNgx7uq86x6N9SrVt0ExJ2b3SY9ePfC5Sgy
da8hgip2DZUoa1gRbD5ADGxpE1v+d5/mbBDIZuZaEqTlcKtrUKZQlKACofubiPfz
WBE1pIvWt3JqRZZCqIgHiYdxToZw49CVNgaz34IwEB0TaG/QujS2mmakDP5yyT72
nlyo+m5KNuri6QL1cMGhZbSgEbFkagGhkaynfK7Rk6n86LlMPM1h2pCyfYK1lYHh
PgwVsAEd+Z/eKzemBkzbPFBtbf6gYyoncLhpM+KX1z7hIiACKDniTslkWlloxvCh
P4sYC8ToAyvfBitidfHai+0e4SRXR50WJOIlAITwOpSuBcr/C1s8CqmS6KQC4wtc
LQOI/PsAHervMVdYdc+r1jtw+P8apLUv62tfU53LGyfONNzEKCKQRXIW0VEvV/l/
XKT3eCbNawRTAvXy5ebG26DwanNRp/OstC9DUCor7x7M5sRTkseNBs2JuCfKVaU2
YRMWC4LFeFGrVSxSTQ9XrlvDRoBbmtV2EpDnia7/4jySNTRA8CHQxW8ERFIi3ir7
EVtxfCG0+iLSOARqN2gd+HacVMd5mGfE9tN5E49pV4liliyvzJY0xc7YA10/mfES
Hfg3ncT8tvTz7zaFShvoJUKtSd6TNro/gd1J/vkZEZ79TEKtFxj2OIa78RQG2+lx
b8GM3FqidPli+NZPyFhwdBPsXJOBTPnqmjsrR2VOjI+X5TYKhDAY1+waw9RwstSg
pmQBrdfc9Sp7l3nJAWQ6b+pNw1GzDxgQAubIqnYUGaoLIDeBCyiYibd3tn4/dTUA
cO6Bdqd+wZ9lsXIcO5Zm4+/9TAQziK6smd+4N1sqirdacTR+gBM8VNppUXDRNms/
wGjaYYYL3oBZGul66JapB6WP30IetsIk3oIQtkO0UhQa1HeHEARoaDWfHnifl3ei
CwfbU87yOTwtIoLP5ZzCjJEgxBcWJpfqENWzkfS/S97ZyB/efnxzvuYdkztrdeDx
/3j0U+7GZf3X8wSxCYtMEkr4uqrnE2ekk+OMfVlkP5gupkuXuSiIJ2tmIVtWEX2+
5YLJUDePoRftBQYQRPLxcHAPrQPdVLaJ55yzGeSmm5yHQOz/n7bdrKL6zet1Q+Sp
JJIv1RuKr47whm0J08Sk5hx4xrZTXMQG4XAfzr2O4NthgBRsaOcMGPXKqhVdhFSp
UsnVwkiU5Dv+wkZpBKBEPBkKuFB48okplgT8yxoZalcpFQ3tWlNVwDBTgHYrF3EO
CthhX+Mv9WIVlzn4VThrZ82LaYrZNXsHeizR8j5P4er5j7WNZWjFQSgjcDZES4Qo
TOk+uZPeYNWvPhbjfxbIy1GiYXeS3sg1A+iu7TX/mPg5Av5XtzdSWL7Oc4VnfG+J
icOSRxbMRPcAib++pIcgNfgILcAjsgClXyVw8/9ItpE1W70IZe0xXhpiP+fX+sGx
B4Tj+ARRzFkpKE14D1Uxt3vLlaPAZJgop0+LVGfRQK4LnugS41LmezcMO6bDLOtE
Dfa2Sqoql0bP9TWLJYD/g10k0zUJbIfBBwCfXnS2EksSG2JFTAT2bppBblahfBed
WjgCsShtHl145p7FafzsCjeauo6eraAR3zkNAQw44Ml7VV1/8hoEdSgWrzHQE+oP
W5yySfL8s0DbEeRYhkQjuyMIEDdICh9q3HS6yRZl8b1NxYf+ns4jd968nN8uFScD
PSF5dN1st/4YmVL2Q4kHcRU10Ae/9EadWchyx3a+Fol3RngJXQqubgML+lXOTHas
zhKpKufVb9l7+cMrwF3BnQqo3i9raiBK8zN1McQPO5hsaYGeBVQ8cra/+aYZ7F1/
DsSFs+4rKAOsiY86Rj5+J/hTBjVao1ntHRMnSvwHZUC1neh302CyblawNcv7haLz
NqnOhAkrlatjwGw+XjRB47j5a6/XxjKbYB8bR8hX3M4xcwCOQNCUN5TJvTE41JW0
MXnRUMsJx+tjzYh83cJnnHh4M9dlcl74SDaFje0bJNmwjVbIYJhIAP4qK4JNdyCd
Q723QLxHbAwDAc5BWQ5+MOcwXHs/Ym3qEg8yqWFCjb/Bo2USfltXRO5jfCJR2tNt
XskPSDhiOf+uJF9R8DAbLt0CvdJt0VWVrQQUBdHW/A/yBXG9MX0qk05jcCBb6Ck6
6/Dn3+KvPhKfnfJa2oA1SKTcZP4KqiKPlN++fPp06ktv+YTm1Xr/54nNzvfDhcwq
kuFC6G7E/GgkxSKzqrcgwUBqsMdl6lu+2e2Xe0DHLAfuRAQJDqkNVBQ8AULSHA/K
uodENCS/nGFh9Z+1mqoLVRWCcMKzk7tQaYthUf6PAzYhIm9QRz9eGjmmZowj/bfU
ewROZ+f6P4kXK/HjTrgHxTdnVF5pw8xYlxrBv6ccZYH0L+voeO5qupUo6dPj0jjH
/CGsUR5OV/8mRCzD7DAsgvki2q2hLBvJKZ0UXNUqksi8E3rz80YVLLCX8wdRbaOS
bnnmcYCMQ3iENPXIhhXCKRIlAA03yJBFAgjYHWm1OjvdtL+AJ/tlh8+d4/1SHJJq
td9J8ti2E2H4I9+U53gZZererOUuqia6BZDO3LehfBJ9uDsOaxmmUQfy5PjtucoZ
vblvq91nf6Gy/COYWSB8R2pG/+h0Rr2KHd9tcC6/Zdc3/oVJDex574Ys3gMRNLuo
yuC1P8ycQy9YmYHSyRqG5Y/jVMl8ObOi8nC0aXFbPkWN6qaae/PECEoqddz8zT1p
jyAlrwpGf8UdPKRfVCccGku49UfYDrlEv062Z/1ECS6HXSyiS3cQM2bXbHU5KBR/
PJCAKVCsdy9mIel1J6+4ZGMoUu2T9HKyH/OSK/icbYDM5k2OGJ6zHmlRTBVKJili
SnJDSaTwQXScJGF15lLkR+F/R/sWchLj8BObTc2fFwu6HsjeAZV80+ek8wJGJttu
pkJKFdDwgp9oPhEr6W17kbnDPikhW8SKB1u5MtqJEZxu4zpLodQ6p9JpFUAmi/P7
qq2hTPmcscilbqFZQYwFInhk7FeMcKBpx1Jh/9jYMtmPJT0fNaU/9iyf7X+LkW4/
JOT9cwmNfhh7CKJgTftHtxJ+PzicfvGUjpC8Xq4mAu7ZH2XJxx85W2lTRacozAvv
v0/tRHNOBXYusLDfUTI3IkSdr/+H4kW+/3ARfllzVcmYbvxjP66B8D4Ld5gtPHLo
aTSvDxh4TDU0PorCRmKU2qpWqZv+UFV9J+9Wh07vKUbQowZ2VzCjAX84n96r+XO3
gr6F5QstefCyYVIJLNYxK0x+62JthqWPB+0x9jxCCxkfT3v47Vz/pQzUsh83WAl/
cqV618WZ2VG040w1Sf0T8NWkMO7vy3hqhNvfznZyO1ZFe9tx+zIfo7y2keoftZUy
++neq8Oj2cdlNFVKiLW7CQymAJSAl6S12h1M882kERsdiyarNbh5u8MkYgYJlthQ
sMcQCcDHXLvaHDuRuU7gbQ28UM9DS/iFWVgsz6tDfD9rR7smBNvLegW9SMFrTF4C
GWKWRJoooaUQPxbIRlLK/sXgnVlyRYzEgeseHSd+raFBQ2N27urZr+Bd5+lClQHp
6aZDFy47UuM61PY4lP/ts3XsosM+/cUjBzwF4FBjpuINNvg6q2yrU3qF0ZSljmXc
Mosa1aLo+EgXll50KAssf2As0WP7Tmx+7UYq1mCDlmjxk9yukoPgjjxMpyFgMgNP
hCq3dNPu2NNJGx+DxjNYNcPKBJ/24NKvHLxmuJnGW6NztOR7yt0z7vgw3E5LP7F6
0C39dG136LHREJFxXdcBOGF/zTaZhqMtV0TywmupwYje10ZDGBRem4b2PJKo7c9y
AYnFtBAQzmyMJ57MffQqk/lA7nQC2HhmfqUr7nzSXpvMCTxLbH52eijFfGrg6RmZ
jCHDcH7kv4aRk2375NmrkTBoEfNacU953CEKtNp8c4fOI7AT0sWgBquZnD3p5ao7
/zd1RtJoAKqLUYP98WsnyPoj8qsP3An6EcVyTzS5xEn3umPho85RCw2R2Rgk9wG7
AsQi97H9DFUovCbN+rJiZf42HimNbMAcwmAmQGR+gyxbGUFa05SDk7QiuSj6bH/u
GsB5VPbyIUn6UdwQDUiE6/gxgetYTIP03O/n+0UslMnjxkEg2Dw/i+K0Ij8la4sm
DhXBGI5weYThb3o9intUBEBsbnHPgB148TANTv/Qgg7YPmUUw0LXvhe9pl4wzABJ
W+iT8l97auEhRENMPMbuuH6LmUmPJOfNOorcY2/vR3kcRgH7hBw3d6NYE0w6APrs
1xpdqofat3SQhapZB+sYSyzjsXWnz6sz9QSPmXsNrApK6PWm6AuEW1QZRst6B0+T
94V436M3s8PmMU6v3GuefrVaBtnkBc0MpvLhfIVV/kV0caaOozHL+Zb9wswhXajn
ZY+SE3DYf2bAuMB2f1AfuUfzKYttKGgrRvZsNMqsTBXKeek3v9ClBSXR1BfCwpib
h6Y9l6SRKGdkWtLLwPEkueksdYKqHkFkUMzMT95UtxOPiz/EcWxOZzvO+dnoRJHd
m86uIBWpdibhcJ9rs6JA0WaMNpgm0KowuPsz0/zoZByUnnLhLPV4aclTkt5sL0IY
Z+ggwXS/ZBmVf7r0GZZq9QX5IQ5fULKSEMKh6OAgnv2X1RyFY1FYZeIqO4J/5wZg
KpuYJ86CwClhh6WVsRMjUNiNVoc+poGf5jyDro+38q2XFJI3T9zzwZ1217oZrGnd
j7XV2Hi4+Bd/IAG7u3FR9R65JguTtH1hQzGxtqfyxP7XqoLEum0t5kRIRoXOCuYO
58jbkxS+bKtaa9Nleo4O4f/TWZjUvzFBzu2+Wwaf6lhLVRUjLJKlpVqBDIUXIKez
lVmGOca7wRtkPG1EwZ7hdQCkLlV9nB47lhTkBk9OVTRZpMl4RtjOdGeD10biJDHP
8GGZENuNK57YAQXefmGVy/rS5uhdttnlwTINE9KEUJck7wzjHY/4QDn3xhkhb+mu
hBjJB0NFPK2qHsUdDrJ/TVWEFsYP9YXh3GXdM5IJPH+bfMIrrBc0FHJXpTfotKQO
Z13MVgnZUCkZtWTM4OPTP0Kp0drf0G05hK2VFz1kMlFCgSiiPnVCN+uoao7qHyX/
TEhNgMlJ32a8KuCkNvKklYeRcmpGxAk4Zwro9pEH04i6j0el5KHtHNx2d0NYLxcU
K/jmGq6ImvvZlFBBb7nqRuSix/R8s6xaGq53IniB9NwiDQmvlLzbCnO33fQt9jsb
9405pwufRdw+Bn6InZa+PulLKT2sXf6u0LJL/mH0GAVRjTbEUvFQ8zVUG7DYz4IR
ZcMYOhY24tDPrnUIHfwL8kDkE5u8O8xPvjfziqSUaESnF0g28UCzaH+dO9wZFJO4
l8M381Gn/4CF8iH+SxeEDC++hMNtI5MWd0hxNxknTCLhy/LxpJH1cd+fyBl2esiv
atooNsPsErsiUj2F4f5AEj/dCfhHvTcTAES4kNgoVTtdgO4sDu/8i3pqTbviXCPZ
N/Drlo6W3tlWisA84udHmW/FM6sl6RUBtfyW6ebbzPgBnlsERivxrHGdo6L18wq5
hBgN0A5Mieaaqge1/swMe+OXnjvP6JSw0+fq6AOL3JoT5t9Q9tf5Um1NAkn0sa3e
fW6r2qluKA5CzgifIUx7UrTiyhWDNsJyon07xi0+ZuuM+G+Q6sjpxYamDhlAJHc6
6Pz1RjPvr/OeOkwh3IucaEG0F+jXNhtfvXHXaSSWY8uw4rnr9ddeyCDQzd5PPSWQ
F9f9zQwXXIS4QoUGPiAQ0C1hEJwuUd4OtL2cHIbgL5oyz992T4zvhbI5hcT6rMGI
T+rNQl35s5IvI2DDtV8yGzsZw0YyURaj63GExL7anyV269OY90TI1NaBw1YUQ6Sk
TNDVIaIxuGVLA8KWy2ySkOj2FcBsbPaNz+DYInEJS3wt4WYb9z+oHvyaCsZtyNtd
EPoQU1ozP3seY0XMv3GZFkodEpFo8EbmXuRNKkb94QihxYjr1UO2WzOccw9UcLqe
VYNLjYehEwkbPDg3EZ0qssiU9BFESWjiVMssY8gYwq3glh2Pcgfsk8H7KPHpkQNe
oOYJDnAwtZq98YWZIM/8DoXa9ml5iRhiNIbD5r3hoTir8COy5MEXpFI316/A7Bd2
6N7cXk98jTsfr95Lv9bZ78zaRcglqvyqdqEc3zoprJ92OtcJrwW0lXBnaeEiN5A+
esU7MabyhwBinCMGPGPw+7F5oEM/AYiize0Gi3RI5vajThS9+2rRGTHqVaKYCx1O
kEmD1pg2pzaGw7WKsR5fkYHz/M5OVghCUrxxqpy4sLtNxEBV2zGYHkvU5nHCp5My
wCVEqqSwVtaTcrP7cV/rcKTtZ1zCBAV883iFLgoENNleP3v8xereFkJ0d2qgxTJt
tzfffO+w/W8jcP+VUKZl6HPVn03aL2MWQJzftppRxD0+1RY9NEHF7D9EaxnZF0v4
8tcRM4wCTByTNWDnR0Bgfyjma2Uc/GAGzfSVstuVxDUNlHk8O4TWZ1TIZzDcwN2Q
Q3uRnxqb19E8Vb9BEpEJeDas3htDyHFKM48WIwprGXP2zUdYMM6bvRO8Z+C4UhHC
6EOlEBB7AynTogeokCJkvr53jYcwQw2ev1FJZFJ69Kwi2OLtBfjbIN/rwIPcTRYi
RLa5UZ70pdcSQOKKT76mL8+e1eJCsnYMaErTvkrFWaMPg1pjhHsLjfjgP9Trs3H1
2ADWE8yK739sKmRcoWNZP8oaFvB8GBaFZYqHRfo6BTsEyNiW4XzBIS/KWIoAjs49
K+TqQsGiKYefsPzn/9++Gt7A9X7l0JowPGHyUHCUkEJgM+lkjT1f/jA35XGn7HqO
TfjvdMaCFjgYd36q1iW+/akDWshQOhv3RbaZJAL8HK3hEfzpsZeWIAMwdffrXJeu
HnIHVyHZw9YVPsWIPasorvTBMvZRIWlyvh6piRJh2NsACHCisi56rPURpAWg1kxY
cETJpqDjDAnV3Psalx3Q7unagxHIppc52dOCFzCSzGgAHKgvmuwyY+A7PFK2uzVD
cyt8W20XRv7Vq11KxtrzyvGxPr939UDpDElniTNJ4+4alaWb5ioJqzHDiiFFBCoB
1SRPdx2VGZlJtBKEPEeWBW6C/aDz0USZ2eMjnZUhEJXsT+d0/NaEM+00bbEQmwdl
BW/cX3GBTb8AS5PlKrBFvPGC83O6O6BOGGuVo1xAmiQM+8R4LQ2jS868KpY1IA7E
YEyVWnyo9usFf3P6oNVX8mgfu19NtwQR6NwteANkVJleTK85/gfc3AtaDlExF9OC
iO0XJWNzNVelYPjXHSBr/pLzX8FxnM5aoSrMr4xY59R1rzArIRP9Q0llNZiPfPxV
EOVb77iJLmrGy1Uz/7QCFMi6bcNsBZ0murhpRqjyb5YebYzBPY8+XmtQ9jITa5pC
WJwVelyg5EXliAxLQdgMknOvEU7aouvcPhvfrYNQQPnT9c52KQFeCyI8TjFP18oB
EgQ1ZzcF+15oqmKoqrDW18czeoWo6jv1NhZXfPkAlJA3VJQxpG+dsF6hRKPSrVv1
0UG7NdnCXCwtBBO1bAT4L2qDpTecaxw2/W0uGDbXFg76K3bhaRc5qM19vbHepzxI
DALGVcVKmLc8ytlIJnURyG80Hdc6omx82bIXvxADbqPNdVQ2gAXaI7DFYnOVqhkl
xaOllM6dsoPmDrg5F6se/7AfdtlLZPHOpqJxq6E3v30LnWTdZLHkW83q3c86ARng
NW/lgiuYz/L6QVrirlTNwKYtCYf1dUV8TbPOFMUvxngS2ZDJIP0LtzADlnHAsa7p
Sx8qPiFDaUSmW55Rqgc5/T/+BJQfn5ktyPiIw7tHTnkXOW6iTcVowJnBTpSnqlZK
fE+LtVwU6AKJPZYCEKd6c6w3d+hzMzBWNZqQhJBtc+PSYxnku1OFJERwcVbfrMNS
uTCrsstBJvLhx7OfiLmLC4RdnkOIjbWrtxhjUz+L914ITF9alyh+Hdo+nsJnRd86
7Hn8soj+IiipJ2dnVspmpQ6Rz5Dik6TCud5H/v4ZpDo2wLFQd7sLm3THrzBHyeHQ
/m5zFGDplGPAD8xMRjnbjoTgvu+MalTHDUibUgEw8D6AJI/2GDmNURgdVxdl0fsP
gs+Rbvg6rKbWSQwL9edchgHeRTDFvl7IWRWNdgWjE33qCyQBi/wsrJO+FRM2XU7u
6Zkth6LqSpCSYzRV3g8lOK0lHhwhc5IZZ1CjHLlzPGmOhJ3Ig9TPuSga/h1dx9QS
2vTTTRefvN744wAxgRDi49Y1wZGq3+tOgBzvSPEdxRrdPRzrASdF44SgGK/nG/km
5mTl6U3VlwwgPWU537ROasM4lngUaBmhGJBh/Ta5J+8VZGkBeaiNMjpvQ4FSLSLC
vKgINVNOUaIf0TRcyXJB8ev7LnFMKNM6f/z0GJ1tQRwbaUeWzbq17fh4UyES/CRI
Wrph7D0uA60eyY05nrS5HZ5YXoUjnPc4dxvsxyCBOKqOCJdYhBoWJ/eHgjIN3UcJ
QKg1NcdG36pbuzvxQH6YN57GiMVpGv9Dt1oo8jbyXb+yXDWxO9wvaFUSWA81DIXf
FgjZbCg2mXGl3F7Wa0eDxyswd4SQOZYZCn7MVIlFV6fVXhRB2eHmFEtxVphSKu4t
i4pz8A1/gb6KZpW1MdKlCf/uO4VMDi6zP/Z8KOIZhNWip9ufY7xG5d5kf8PZ2IYM
0ud2sr/P85WUUMZ9A7z/2Hnq39BKX7vWfyZvDkHX4ipNBvv1Cp2vKy159LYAnzFs
v1oRL6hoKrn+Smla/01+9PWWxk5kYrMjuGSfsza70LDTNayxxXiBmC4zMvCx1sqr
+MYq/+hMjvDxjqsanmqxVKEb5d+z7a312OSfQfEnvv2wSGsdS5vEBkDzyCidAPNs
pgAA36fox5kHN+EWNTEjqzkIsNyBuSiY3YiLECYIMDKqzRcpmUVMZ4MUahqOnSyR
xH+oCW9FQ7VDt7/Or1W5DT5YXbyLaKXsdblXfFKpupCIyGriCfXdSv9XIwGfDVFJ
Qf6gC3P3KiskLxZP0K/NoULA1JvP93bcncGs+1eG6tXYilc/faJrGf1rERs4QKcN
qOFT8qZacmM5UMNSvJtfg7Qe0YggMnRqvlUerk6WdZo6ntb1hgAcOEcFd+JMCi2o
xLM+fpOVqn318TYIx9Juyyl1Pj4CfrOOhPkQgv8l4V1hMQyMlnBfwtVHKjlFDgAP
SXUnTpoFIlH48eTLiqDeBxMc+Kc1oa1gMmwa2/UH0CH+NdLVwlLq9c+qqRc1bgXH
JHh2IEOdze6Ox5sB3SAPD2lb2dfC6OC9BKJAQCe6yomK1+ZjbQGiLzgtUp4vUBul
nWxqwYXpdZOkq6iSAehhKuMEOUGl7lrUC5UMh951/qjzGRmrboeSX023NELacVwV
x4/CSZFxP/XD2U5MiuDRS6PqfKtdYmfMtn+lygV/Bnz1FV/ytrgEBPnHnx0M5pRi
8ABhBwI1LJyVPyJiboCo29aOPR1IERc4lKZ1IF2H9KgMKE1UySklzr80y4PN882J
ty5tD5qu4y9h6FAcKPoKQmGRpOe7SBuAPKpbGeANwCEHRrkLynN8Tt03JaAVs4p/
FP07hHUdpD8Ys2wVsXuaLDBWmxJzmTQ5xxcaA6x/44JRzQLAPvhnQg5Va//BaUrH
4StbL4l9KfnfveEeGLZoakvPhJGzlA1on/MhsW3oyGyx3xj0nPkzgEzAo21fuMXO
lehgyeGixIM0XDsNPMzCpedriRjfgZ85vg1I1Q2VX2O4aAOq2Bm7LxEJ8y+LHEIq
Z/HJOwF7hpmRKyeUx1XnsCwVVcFliY4Y6AvusSSYoIJsBNSufS+tdFECLsxqKw8H
nt44f2NZfBl5AMR1myrufp1Swr0gGvUHi4iVeztkAf3WqYrrMHBtLInVofg+CrDk
jkxjoGLSm6F2oACVGcSzTFUAKWFdH714o19yK3LiBjaoWwEYRR0jBsORu0alRdpL
xxpCv8EUeoEjEs7Ol2dLPyyrNK0u07AGK33ug0UUbdsT5mq7xu9SF4D04g2MumnA
Jlsgu9jgnB1lVgdl4Ol2dM8iXPFZhLUTj8x8qTYeZpTojLxBHX7JpRoBSNO4C6zB
xdbGqQc+OaeJhgAQ78A7qIhwbWI+TmkCjyrGK9Hgg7AmmeXNaMVMSAb1B0RAdrAJ
9A/uPrIIedpYcHGlENX4MgZPMvwRdzoisAuGhvqYiBhZCq7m7ZngMoSNBCSzrl29
OqYXJ0TsXY6JsvZ09u/zfDHWSX876qpwBCyN2VC3krXXN/Y1pXsu3S1fF8ftUfYF
f0OnN1huNBS08DiQDTe4Gn3zUMb8wJe9dqfsh8PbesTwxHVwqwmBMe1EW58jY1vD
szwTNnruqqkHrndAvaeDMSLH5W81lo8K42/BGA/Df6CvhtMsTMcmlQpCEdH+fV96
QRG8n0f9DDG88ZggizF+r/tZrMczU0rcFmKyGHwHLvyRfPKl55shWN2LJAA3trdS
Gsj3oamC/ekc9m+EVJJ9rMZ0iA7P4+7usLaYfGsoKWdFlvbfsJZ94mThUCrPp6ZW
4pzfDiCkUoUG7GxmNo4A4G+HvBGMK0Cz90pnmu+Ocv2y6inOGULSCIJwa0wy0iWt
86CepM1SImyQRTAttXU1ns3swkXYwOcEkmDyQrgZ8CCFF0cjdRKFWcCxX3/Qd+Jr
sLsl2KcuHp1X7Sms5ttImJTIZ3MiuzjQojeQG1I8g/eorP8TAc7k+KbBfK11XIy7
S+xgzd/DtcnQGdQ1vS2TTKh8r7wqCgo721Zqk8/URtGxF3eRRt5iO+yzyAJTRYCi
X8ExiiSO7IjU32DqSUWE9vvo5d1vleceB+8OLV/wjtthNTCWKaWJ3vVzPQUj4hbo
0Laz6ipJg7fEmF+8wgTeNBtKVn9RSHT/5br8KG4AisuEIG6Tg8EZwauXTyTh4cUk
EsnjDzsAZ1i9j0WUnKJiKEBaDgJSqzo1O+hZTNXhwb32JY4nk/oboR1xGoTI7NFW
WdnQm1yMW0192QA3cCVmAVCfbiHcB3vEYF660yCD3Nlw8OQjSUJsIzlW1YF4MzpY
CiT983GJnHC+U0L3dLhfVihjveFarlxmGaewMD80bvt5WnuMM7hnLHfCGWuXMeiB
3DMTQzu2M28tO4gi6kr8hYH7ny/E4gWuQQ4PrVKD+Ju40XwN4mb5S9/yhwd0KAw5
VAzmDNPmxCiBwiVovhkQRTg+ok3C5s0iurEBAAdprvw7ldKKRa3LCDSoV6/PgPI3
Dp74vXRTWIQqylBDOZQQPKkTI33dWw+odcadyhBsg+3kd8YvD9ZIvQKXu43OA6KM
bHOvVxvt8uFnuNcmdKouB9Vm8r/oX6k60FMAOcRpQ6HMg3QkxzVlVGdoJbJBjOxX
HW5WpnS8lGSoWcFeq6H3tfl4hBBY81Nr0jFQ+Z6Yt78XDc59RFsnXBMo6dDejY5O
eamTbLFPvNgm17p+QPHPIomMMMs6iHI/grW0KL91prXXq1BRLKuPch36jqpiwg8e
VTN60cj488WhjCUXjH5vN7dr0rkutAvmfgXzJD4ueORctOPSwqj4yi1Qm2v4DJPX
e8y1Oj9SuPcFpsTPok8ezOjTPWm7BjCOgZnm5nwSXsoS2o3k1AK+fGhVkbl958VG
i8NcqQtiHeUMNBfC4MStnvNZtJBY9AumbqM55uK4IEk510O+7P6UfO9DHXy8y+kf
HcCrynUdlUsJL//irqUSqi+UOPWer+C7BgYnY8kb//SMA4jNtK3zIn5u/d1JbqfJ
UUu+O/sA3HrT3HFoUtuobe31hrZXk7MEnBkKaga1fZ5LBMwnaVo+PzYC6/zxH6Bw
AnujLbds9l2jEvmF3HPaFDNZO4c5q+eVwVFpFkn3Zs5OaBlLzDJ2+M+Iio8cHiax
X2f0CCPA1j2cYBGUwGrazQV1aCumdIDl1OUwcyIKzUHYnMsp19pjSg28gvzjFe4i
jRdMuFy3k7mRovWqsM8cXIjFYqja7FttcodLQSA96h6x/BL6q5JvhdDGnMhxtj8W
OkJegw5HuZIQIAyrpfg93456Y/efq7ha4Oxze1OLfeT+URwT+fioCw0oCMULlkwz
EhksHY0MyJf4gzsuiw4c3AoVfCgpjmfOlU2/KYHblI68jWnH4zAq0e0eAXIRaioi
xVwiGy1CUejid6rIrD7omb5ZJSUIlK/jso9jMeOQrXFgHrQnvBm9hJDYyhwiIm3k
X/YsDEIwKcuIf2fKSL46tYmocq0NxObEiHkQhh8Ppba9HM3gvcrByxRJt/AAYuPH
O73NrSiugXgBX8PUeQTNGH49Tk1bhn54M1940ynlwRYr/khoTKxq5OoGbddU7I6R
BjGR2r5buBMpOlwEr73NoD6pjMVGlTFyCrQAkUgLL2UtgzXHxxBzoCtTIyN/9QBj
3DhuD+lz/pYcsq5tAtiQaN2c5b1NowFCiFgchBdT/FSuEOEjsuW0j7xuZ2/JR5K9
UBUp7cFbsTes2DHvUJQxqDf6C9MCygwyTeYeo9SILoxjzcdWLL28ou+gU6okIr5a
y+SbSaPpu8OwvxgF8jw6t84givas6lGpF/J7m/M4zTIvvBPXC6n/4gg9I7muRfMX
aaLyN7ry+3y69pxJx7sn55ZVzuo1Ah08N8xCBZDaLWWcHKWcb+G4BIr1PxFKZ9+s
UgZrVa2iPH1GSD86f4QXXnVZ1fOGAUAeJekNRcXqeUrWNQesXpHS6o5r4s41L5fa
qjwCzhFEsQ1JI6XdDS9kVeRW+97D+wyDvGMm9FZWHvRsqLOLThHbLODBEspp6ayE
nVD8NMG2u30s1FvqGRiZwLjGnEbpcFvKXzcZ5XgOXayc/ETFrees6Yaob+kbUux9
hNBW3FuzWe3mhJCkmFWmPvZuS5zLPlg0Qr9r6oKO7rgJavvZ+7a/btaPQzuKaQcu
/2Mw7MoC0uL5ZQtOJybukKrZ/vaUudQQS+5yAw8s3pEVZpLKFUshdkNYHwcJr4Jm
Y1vpMFd25BwJHK+UxQ8aVxUviYiOj1Gy6fu1LdALHuFNxwzFbw97ptdDk83IjqMM
PqpSuClBJnyJXCpjVCqJRS6l383TXwqJid8CQhJ3oMil74R80hEIbLBj1ercyqLs
yy+FQlM35w+p3BwF3QWHmg6sYsife53KODQnwwPLGAhNFKOKguXW5YVYy7gS1Ebr
xPy+h+SWTKRLpm6WOATicZA7+Buj1Kz4e1nyHyeHJLHNDt6SxZ1iwssUFCq7m1yA
pBL/uvYeubeUlYLKnu7uMqpveU5cUL8v5b+66rVSpkv+tEnUmLwxBNNaQTWEMuhd
Jes/3xQTalygF8qpCNRwsYLoxONq1klHoy+6NqEOpLZdM8k3HMzN4GT4xNlo088m
hqA5jIux0MBz+eodA/6rDh/beCc7gI6SPVlxfbRr413aKvniwGt6wj7cOQdtSB7o
i2qidDuBfRg4kYiqx3YeIH+JoYZJxZx1MMBonVHsVTkGqcfDcRHapu1k/6TqEGpz
ogmDzDsPOrWf4IpRZgZqJJ1EcrbEsScwxyvqIHDO3Ij8iYAk0rOriQCPloCP5D6z
wZCiTxrXFs/BwSRbSjFIU0fRUeU083L4LU1mcJRR+a8KXh6Br2iUWNRlbH3fSTyt
vOk0MlCXrET3ghsRtARgjETued0E5fiX7fqb8pFxiGtzrRpBCmwMv27haRAtAd1P
4UFgLLNhLUr4zr35klhdx4DWx6RkXRms+TJrfZqgp+VIusMFU5j3TQr2h8Q0QhoW
2M9leXWLQJBdgXiKjDaNKny+eWTfnyqItGnxWv3vAPExKOmqsCmxyQo6Rhy/82Rj
pJIF/Q42GWlm0dBrwertxDa5ntIHa6TvoIKgcaLJek1JOqH8yLM2jHse2EdgJFMO
1qspDzckgwF6qzekWU+bUeVBNoCQYoOxw2sbEYYRN+BOHN0oM0qxMTi/s/tCDtH6
iW0MPFnMfRoYKUQLExeukG9HDb962MOxmpYSgjDZSzOif/2HrAdkAV7Oeywi9rB4
h8dYu5VbwjlOpID3Eds9kVwHPij0+QVTStdTIU+dNTQLsbtnL3u+r0SpnKiA2wSe
C3WDcDSisCV4yG5L7wIgCKvcGgndmdNgl/tmgjlfePjkAkBiI9Y3iglCyArCvrpY
OGKcjCP0hcUHaK4XV2oUEdUaCiUh8rv1ObSa9lZflOF5Kzpvu7Nin2Bzg4JE9P23
yxtkKsovFrrT9VHGajMzNo9s2AhijKvIrKaWB4xeN3iAI0tN2qymzfERZzuO2lsd
Z25v9+4M4ZnYCFoXs2U980V0dJStUbTw97au+0kA5lD+5uJ3zkAwdyFFgb57hMyz
F2DC8Ki/e0FiAocBZpIDe6KKxtD/8VmneqAoOfpbENSzPDXq4rJrgUoY5r53Swc9
jsWK6NpAkLlfYfddE/P+NumuyQrFmjyDFuR/78zLZF8crXFsklh+Z1+pZXDp63OQ
BJ1yZjEKjcJ2oX+zItKQMePtWQnwLa3V+R0MicTI236d9zv51z3abAMN7XOIJNc4
qq4x6uZdQLtx4Ub6TXTwvoEbr4EhkuEIikkg+z+VAmIsr3oGb8UVw0OD6vcVuF4x
m0IJrFFN17p72rVbbdeLpKIPCRMglfUQ3m8cqxZ1Cg7x73yzwSQaz1jPVHjoYRlE
Q4i9gJp5adcIYxJpabHxMms4MnU0Mf26uVLIVeF8ht2kkEW91r9iuJaN2Gbl07px
nywP3I0Qt21SJW1Urdd5UKtZdPMPwgrxN260KRFs2dqAZu5xahAw6halslQkx3cE
+xvPRJJCi1RgQ6yhSYxuDzk/IGheV8/dNbXi56hmUEKNIZrhbKd36/j4LN5ZWox8
JZno1dIqmjNud/6lTkowD3MORznnxNRW5txNoJH9QE8iSOh9peHyXm3MmLVh3x12
Laa+CmYh3g14IqYcRRzVozrUGcKtRo9mTAWHQBmhDs9SVMLmYQrvtc74WU/4jvgP
0KgBvpIDgSUZ1IbFmnBLrmtJUxwiYTThutsnHle6ucJ4y24cXy38kHP6ljFuPeqO
l7AnmEUY8lH4bbxa+KXWOxoWjzSEgGwUDTWQg3aw5Ti2D0t1+u5OhcMjyrvVg5z1
17JLeMbVGZGEtRzyntEEFIM32nj8wNlmJjq5uUq3hAbhef2q/cyhKD/AuLFanLLr
wokQOOCP01j+LFkZsHmrHKG+Ryg5a0ughAs3WGrJNDG7d4JG+eOp3TLd/alzA/Rt
yfLmrcE7oyMs5KZsraNwyO1Tn6COgiMTSWIHdQgzHur+hElSddn3HbxeCQC97VCq
3dOtvCCQ7n1k6osYpUbi5LJF11BNxud+b3ZFCP/uV3X+zaAAEUXM1Xhu/A6O4xMT
yFNwXUl/K5bB/BjuSMMAwoZPKLAfsAoj+XLcQHnzPMI59WRYyovCaeC3m1IhSBqs
OqFT217nt945JuV4fqIgR0WEh+5G3LLYVbLBoXv42vmg2XDgZIlkBCzPtTlZn2Ll
dt8rPkUujg1pwHtl3bN1ia85+hppRxTjFhbJNVV+l1sKz0mZK+HBq9km/Cm/HSbr
HWbANz/5UjYwsM3aBYTl6uKrbv0Ks7KBlnb8Oy2qm4bKdWxBhmwjvm+q4rzc4LbB
Y9BLeV79C2KlOhqYIwp4xI+Rql4r1qnJs2WCaQ2XbZ+pH5RkpcQkN2W2ETCWQRfU
gYKKEYGPRlkpT1j/NEq7Wbg801yUU+xu+NR5CxvGaluvZMMuy3xgkTRuWma0AiLG
mL6dnvToYf2JNcMIjD2jkP8CttiGHE77yZT9xrJ75qvP8jaUhlWoO9S9gro8YSn1
LQtdP7Hwnrv5LD0zhPXsoiZn3iks/SANqX6Nd5MP5EiHWFdhedjK+sE4r+Y5GHpp
fuROaLK4QdaaJ7Vf821K4w0kNLUaq1sJFkpZnzSR6AeaVm6Mh/Qt6w98XvFpySun
btKjgvNdhBwfqKK5m0p6aCm9cdvFWZ1bQjOohHQmlQ9Ma+u9zvGk8bc7tReVlQ3j
i2wFXNm1pQXIa1CfLWKs0lmTCl+vn1MMq+lqcT6AxoWbBM4MRI+peKDc5v+JbPkE
Gw4Gsf8G0/+Y8E+asjPrmeMwyade42tgAnb4clYD+nKJHnexyT4UCkHw3tg5YAhS
JWnGpnYKV2pm0o2oNf6G5R1EfReJDH4pnuS5fBq5vhnwsD9bmd56Ua8uOzL3rTuS
rcBs9vPyOHsP34GJqgZDt/T64oubL1/JnronhfSgxdox2KGUyOMwIVheEudBzHTz
N6D97BM1+GBrPrYNXkt04qvi3E64N5C6JrrIfchuwvvmU6lJ0UPtXoIPFGlxMl7m
Pf84+PBKgAGD7jJ6dkJBTRlowHYM+LS9ooBo1gyqgrDPuJZwb53d6i06fPWDSv3t
6/g2sBjY+FyoZRPFXQf87JbJfXjxiBgqY4nQim/7db2x/mkZtJxuRAbRvG3CCXSo
uBR9P+tY1s8L7NTSAXB2Xqt2rRfl0KCOVEsxcD9UDKztZEw13mFg1ibvgz3jCiAR
0HfrZCsUyTyZqYPKoOlDBQIoHxkbBRe20peQoo1eooo7rinQQCdXdkjviqOLIbyk
JT4RLW+QKnH6tHOgby+byOCFQCo7VecfZ2BoIMLOEYazeAr+Bt5/Yu/LGjaP9o/j
YZuAkGOrZZsGsIVmbTLDT5MJhuocpH5sCLdyxmekEMD8fQcp5AJ5CWLZsWn+cTKN
/Bw49TQZHhd6YF5BFuGnoI2+MvSv7hp49Aad5n6P0OgFqntLI0ilcLzpJzKJB9sI
LJKWB6afV0h1gRitTaMjjZtM0Ym4DDWm9BsamyoCLvpsJabAiwByBNUt2OQmtx3G
w9HFAMDTkHCbt9JxUKHJY2N/lprYUwtYCKfXmXvgBeUGlTOmg6ml6OLQvsqiYRXP
y0naizJyPJDmFN33T6tC/H2McO/KWbQTZx/syDtiGBfT7lpfiN+gMSf94v7jeCiX
EtN1hXEwqnbPm4jcDrYt6s8bp8Ghg1hxmWEWLnm0k5IlN1XyPddoM+51jdivBD2G
r9u46Vy1qFbHYj0Ui0Ht8JIPD4PYu8PIX3G/e9gLD97IJluD7g1mQrWzu7BdZHUk
ZG8iz5bn11bi25/GkGMSp46pjlU69zbRMK3lFU1fzqn68fWX/ldBU105E3DdziuC
F4Nj/VWifC/7x426LesV2HbM+KTQ1qUi5WRxdqofBENf+l3F4oYxPY4kk6fZvpRz
+bbtaaUXLoCLwIZYngqNV4oBsV35+sVbllQ0swIpzS3bgOz/IFKuKXUjiiuD2fe8
/Hh3JuubHLIV+3K953M8xwdvRySMU4l6d8oqNgPAWMB203pUrnqpDfizlxiCQ3WZ
w02ZCI3JRhG1/PgZyNFTshIrPiH/TH59D1XGTO/baICf3cDEhZab92mzInwrvdsQ
QWua6YtEArWrjcryhKNqy3oPCqk9rNUDVw87WxKNmiZEJEemGn5LoxNjAJBIMrdw
DAp2mz1m7rN6ODCTyF4cwoWnKCcvosq7ef1OtxI3oDpBTan/EmVcKs7A/GCt5HW2
gKFK/cTJZxIIgQKT60FnC46CzFNW0VhUWQzvlfpPUPM5KC1xPVPgfX6LOq+2uxto
8o06goek40771c3t61yxku38o58USUhUbEfLQjQQ+LH8oTYvgP9UyknMWGwLi1Ii
cTqFNn6Z3dFm+z/kJyTyJzK71glXN0z0ics2Jo+a4sZtuJMfxfrfKP/G99keZkV5
WOkNOsaqJb3P33KQ8Kmmpiy3f/K/171RwYsnoYdV6thi8+/eLXLMIPqei95CHdJA
3uE5e+0Z4VxeEQeOQHbOG/oLdUNOkEDbkSdBi/SrWkku3kBPGylyOprappC3mC/w
kOnPf6xMdI8p0tUzwqrI1O8x9GBE8iQ6HYGkvn7xLAwIk8+JtP//vS9Xn5Y22pPP
oKxymODUbzG5NFOx3q9lZTBYL5lNCJfCSGoSJM9g4SWkXXkFMB+EqTE05wuevPsL
tkg0YdECUeGNXTiogm4e7PXxW0w0gHavjGy0DGxeFRsae0Z3Q0/CECI3hR7otRSt
qlkzGOYyGAg0MdIKczqOa/FJQ+qfh3soSKj+RwQsVlCyBnp2wx82KvO1qDbbEFGp
mJItNfzsbQKLPIFmg0KzIlF34SeN2sJiEdnBzEDqBOonZ5wta8EYr94r1+ItbZXN
sS72u7tHROMQcQQXRxQW5VaNgRucImthc4EJFqHsw7hgw88Y+cOn8Er6UO5Ll1oZ
tPUiI9bhQ3eE1+kNjeYqd0eXN7K/kFWyN9Oo/a6+kD+WvqEoVPbui7qZ7TZvPTFZ
4WNlCV4HQe95SpIDlNr77V5UeU+MiznFzaaR2V54jeSfirW4ERbsvOUN0BEUbEG7
4wKIl8nUqWDgRI5CvkiTl3uPpVkCxZ5A8J3nuBUE1G5X9mEob4RkNJ2DOd/9GWXV
Uvv3RBT9j2xCicHuvj0dFFHNGbJ5Pbpg8W2LmdbMv/rm7lteU9VPOwXzIH7cj81k
WaM2rtQdldbWkTwd2OIcQqxPTom3Ugf5wqpTkNVo+g1YdE+Xu3zB/l49/BhviLN/
JuUo2sOdox47vQ2zfhbZ60Bzx2n9ekg04DMu+opv7w1R2c//3SCFWfbWFNreIeHu
mE5G45r58xMeRbw4YRHdR6woCZu4X4YCv43qn6EG3cm6FCmssm5TMfImpEXJbOxh
UAnLxsc5uH5b6bFAEiEzLdsMoMBdUTQ38UtNdgRa7bKhUDX3bBsCtTU2MNxnsZQD
o5UZFGsIzNAANHgLqqMzoDjI9HYGADyCH6OWJnm9zgysTtQ2HN5r0FtPl8o7fs/P
BCxMTJg5ZYwOTjyynblT+YyCY2McU91Hu2Radt6nIqvJ+vbgf3ZjBWQVMvXfpzXp
qx+Xb5PNaYPwfM1CwfwZpNH9YPvsdnNrZ/ba2Bnnoynu6m6RDJa11HUABralI9Su
zhQJRN8T8I8brGAgcKRx8hfNb+08SDBdojd+QIMzzWwljNEi0xK8c29XMsBksheI
fuvw097WCuTUn6qj4pdeg30Btg6DkkeLLHBxVfr4Ijd9NRTXWvn4+Ck5BzxQ35q6
x2GH/L7zQv3n111+Op8VXHKwAdcdQUS4mK1c3EVXtxhMuP7gZ4yav3zW6LoTA9t/
zPdhEIVujflRHNpUVn9kKwbEx+5RWH8i4cD/AnDZIWxtalxRAmVOyBrTSxPwXj+3
bZ5weOHvkvSgB0Tbf2ieFP8OzQzvnchguA428+DnRBLJF2ehkzVV3IcQIEXxcUdn
gOW1g2xvLYzeVxPfSTcl99iMFLmbQI5YMY6x/bGAv4HldZWjlbBipSym9kPeaNAa
ZTCL3rt8x+T+2YarKxF3naynD6KULrrW9vjeN927/ys1gZugdffZ5TNTol6Xn0XA
wWhLF/dQD7Rt6dTxnd9VgJGR7XCQZc08YW99N5ChG93dNFvBIJ9Bh5f+beReLc82
Whc3tP7Z/daPnqpOnMbRPlXFIQxJkFAfuzvw+XtG4AziVdvitaC+yx0bX08v11nn
ScMd7poNcZRpdJDOHbyL+x97PijoUjiJ0lEi/H3VgxRrwwUpF0zAwo3zdUNOtPMW
zVyVl6cjnEx5ztUpe6RBSyhVNbhFsEXcDyk1v7JzkN62vNSrTdNXE2F0b4WlMg/+
VvviSa8+0cEIkLZSQhAerCL27lHOr4TfvSd43OdussvYV1gKrIVza6oJkkUUmX/c
O2x7bhOXgHzYbejbEpP7rvf52io/PDZYon0Vdxdqr5UiovdcnWPJSpn2rdtWvV3M
gaaLmG4VYEpHAkQZdWjE4nXEddBk3/mU4KVRUkFCOsArgKW8SkYNACssWKS6b2Bk
Tn9cbKz4TNDWrzyqW1NjG4hHsaUnqUWrkLETh1c4JHcJbpOabyV59uUQz25KdPVx
BOzij0jTG6LLCTTCbUcIGtzWh6saFm9cl5QQOnqA+G/74Ku1LXYSZnixbgbet7VQ
oIQwaoIL2xPfGlpgSDdHk+oWLStNpHPJz2IPnItbnAruLM6kBtoIVHNBNXEC95Ng
EL4sMBnxcFIpSDFRaHis9Vn/QYKwjVIDTWWcMSGmmlKE45el24n48+BW03PVfTnn
jujitS3YqRuJAYwrkgSxtnz5fZ0hYVagpnrlYOlJwLB6uZyD3Kb1PmdGpoD8kDcF
tBxh5a1P93JRBrZCAn60ysVU+Ka65kELH5s6s03lJioGTizLkM+Jngr5Jv+JWOGO
h29+xIxmnkHBLZd0crmc5UAvB/mBIxAhf8Dy3V0tGKErDdNTu8v6HrSAqx/WSJCX
sb8WB7+Jj8tunTMefQQJSjrjqSx3C10Tc1LyVxpYm6NNY+V8EgcVrMFq7H15ujJO
9H0H7W6u7MPJcIGQU8zr24CEBaDnU2kJPp6CjJN2cD5zMicZ/2x988kYlli/Vxsp
UhbgaiE4GIaxYyo16h+NxYxCt9B8H5prxHbX4mGpciN0MFe3mMK8aWi78k8iL6q+
8Cs+JyyBhHQhwNoXi5bApuPSpWC4tMPJFlxMZshKOGRR0eaPA7FYcYBLL0UZm7uj
wbSs3eQWKrp9T029h01KUlUVaPIJ6EH4UIQ8H+fF3qH73EV4Ort9qKhn6XLTgp/h
Pakj/VCK6vDvBMAYSF2DhGbG5aiNfFRbYESBwyQn43XZHXZPP38CN7G0A3EGtYU2
+a9oNGS7pSTmlG88ESqoFWZ1Q8N8d3pX4z7Ou99SZ2Tozr/CY9DlX4meneI34dAF
GmOanCWJCHQ2bK5Yl/EppCn0Vhh5O3segnKvOPw3bFktnbybNrwyLPk8gj79V8e6
1ie2MaJhotM6j27iCisaB6kCLPHu15t2ZHK/n3LK79Prijyfu2PrOX+mCivnRi0N
r+RCLdmDk4laEHp2hFMjqGClYfBl/2hDbuP4GAtfbdOZhVdyCk+6lrdfqge+oMm4
L5lR9SZSy6C0jg6TNvTuZl1guCOduDUB1iYW/JdZjayIM1hLp3id3Wa4OMrohAF6
aBtt5EcKZvYy4PSVV4LHQGmqOwy8SpDrJBpsfA7FzCK6aGzSZNllA5c7Sx3R73MF
JAn6mUZAL2U71vmRTvp8VF+4l+dSTFK813Xb/qzbKtIFONuWZknpWoEQkwahPTeE
cFcy/LOiTdQr8Gq0YBzDaQHoNaX4I67PWd0/9lAbquE/0uRXCVrLwt1r9UKMMcpk
iItBQW9bnHQnaQ0V5KMqx3hQuuPtUFFFKWn9MufpPxK+Wz2OYk+E59egMsvHTQmg
jU2u6s4sT10XpVOAHk0CxOT7OcJdQy3RUq+wfAuBZYKIVSy4EdFPXcFCNZwJEz4n
O88Bh0EvWNPhvxUqi9k/NPWyP3zCNiSy7fQzP3JD2q8lbN1Vghv2sraVOgcpK9pH
oC/YOMotOv5M7+ks1QnEk8V31Q4DdgpsXryz0Tspgnt7jhQ86twJOIrrGnH//RCp
rDGbr5D+gn9OsKzdHSTG80CwWIHhltkxxf23Bgwxvnh+q9A6fYwoukIyxSmjjhWG
zkgDcLTOVdnE6hM+9LFbDsnTkS9yisZ4qdfktxjMLo6lLYyyvMhOPVZbhCjz/4hp
oIOTXhgrOakfTP2VbwjdEK9OMJGHLPvKi85RQnKewWR5XmLvu5P6Xg+PziZoVfaY
3isLJ6G2DG6NbfrKCapMiP1aIquqUhEMFM2cSH7Bfo+PeIBBx1wuZkghTCoMXMiD
d+WnJt9rnGxuZ3xqPSfKfIllNo5pJI9qMdyDZIxenLXoQ6GE640mZ83hIk+38N6Q
/DeJkM4IFTq8Gf84sZfCP2HV+Zn9wZBWYhz5gHa2icQKZcANIm4Tyw0Y8gkZA0tv
8+nAeAo+6eegOFf0QTmrUVPVPYuA7r5ekk1nsK32rRqrG+nhfa0zqzQcv28ptBhK
`protect end_protected