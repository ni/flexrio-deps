`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 26864 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
VKWNRQF+vfUNEEp7apOJOSVr78APbBZ9xN90qYKa1P5FkpP5YeEQoQiyc/Uig0KA
Nq29PL7H5MgIX3nSYskDP8qVJ10HOqnjM81qysbktrv4HW/XsCqvUSypmK7xbxsQ
BSvaZqkQURIJV3Mr1VC+Qq+8RQDkUaI2vB6hRT8TjPd9v9GxH2BSjrQeiID1tqMM
+dHU+4qIUTaWstKVZsPi+9CtCAr9iPV+T6qVLVUT/0r6PsczaJtpupqssZdv/C1k
0cIoVFBOsqMHUdT8pP1+uUQGDnCleexVbrUe2BkZUIQU+MTnCs10KfsMAzUZ6dHV
/ppM2oGHpHizuOX315X4XfJlbwFfIb56yfeTl8N3qqfw2t3S0Rr5D8RVadnAzo2b
xgs7GtxC9/kufeSwTYWjeOM5C1cWRJdebXM3eTdgCvNjtvhzC/CuMqbz+MIpBSSI
H1OQrShYKTaQmpTKYtw45vCea1fbj9Sccm0MeDcdd+LO0v5FGvlbKBqR7q1SY6Eh
2t8Sjv5k1vwCfhuRPqoi9iy2qqXBgnMxp/umDyGPbqsJWlEEVvGVFegZphle50OX
iG+EE2o+Mb+tTHAbpSj2buNVlicAvKRkCxhwMXsTHFseQyqDldNn981Rq17SVrGP
4pILNM1Hd7NbbrKwKAFg6oHLv8Dc3wy5jRuHT3h7MShz8Sip43hjfNp9jay5cG2M
++EB913fmw4yp7xw21QMZEMhA/d2jXWGSA8HE43twHgKTImR2x8OKb1YcpfJjUNm
t3OS75Y1hNS9JdZcy2BWXifntdb2Vr7x3hu6vbqPwN0p9N/khDeU7pSbgbUXo4io
iFFXO8pZS+5NNCX6lOgJEcN8Gpg+NNhi3+a1D7ymAu86qAe82hiDMv1B3tcmb7k7
TxSd9wi9TKMrbkQgAeLQdwzX0AGp4e7uoiI7vWvjwDZuyK3hRk5jS7dSlUt1IJv5
CMh6M2hE4v6D/sDY4WQUQrXRMtIJLsydkljUvEFzJeYp+ZZ5mI63tAwloV9C2pCO
VtBOCYTwgtUz0S833qk8iCvmAoRgxJb8TYaqEFfST99C4ulr/sJeXrQDNyrBIB9g
agAuWrXBUXJuH4bOICbv8kREk22fcB9VS1wRxJu2UQqqieZrPmy+ImvQwEAvbFLu
CSuwDWaM25spUkbXCaQopCJMYLb+oHcxXW098FHFR4ZK61JRPhUOL2/bG1mmEeFw
9WOHYSdv++l/rlWjY8OMeIBhMet9LCMPyVN+j4GKE5QIbbp/BG8p1OMg2XNoagOi
WrV5mi59cB78V8pADPc0QrcH416uMu9zmGKqCsVhWa2UQAEHfJEcL8GS8/hAQKJR
2CYE5GeyK4LB7dZBbS06L9WY40EBs9he4G+RanMAXDXqN7oqdLQRHhDVomLpU6T1
RTDYBSKJb+gCAvj2WGA9CqfCi7Sidi01sTI3o8LSxNfvpghW/m/gcz4DGKQrmts8
et4IEtJNM4nXQLmb9A2EQB0XftLBMDB+Ojp34ORxvnnujFU8p0T3b1pnYQamBTsk
B879l0MH+CYNjFv316FqcaAMTm8OzimI7e5ZNBCg+uF2xQjCBHAo/cC8o5gouNs3
z0YbAfSX7Fajar0bv6/pgOibraPhJ5Dw/n06EbuXXAtfz57yeqdUuVkiOQQF9IAy
ShkNo/oX3Rfae6RA9lkODZ8XDh3OdISvYqfIe7ysIADk5f/nvdt8f+zMWzNzsoak
Aa6FTEc23Q6+hfwwkyb1bxNbtuFaaQmHuKzlzLcOlFtM5Icu7VhrRFVzelp7DpY7
lDRdyO0tSh3pfpvxXo8rvLcvxR2hk6C6wQLnniVgUrdQNM6S589e1LL8HuGWPdWT
PkXoICntskDiuapZkBkKaK6xosVG+f5TFVHCYUdp0NxtcZQeX/5f8vcVcvl+GqSq
snIZJabw4hyhp3aJ5le4drRs01ltoKGKpmqZ9WxmnXkkER/WI78IASmj8/If9t4/
uAa9kM29dQfITwp72MJuVquVZI4Jb64+V4l6UW99MPEyD92gOpK5cqEx1HH9uIXT
iHSYYY0JWvaV41I+fIireeTtRrZ92ku4V7A6MAVBwfpjGEuYG4QCETTIinvpL+Fo
SwZbTbR6gQNiCw1q7ikV0eWIabDIn7skLc9+7yWLayFm1BpKu1utvUCEWEM7lJbM
1CV8bAwxICDJegnNZulm/aAk9+Ea5xiGGs0fAoIFIo/DMd4UVgNESN0BMfj4pFy6
jfIlLRPdVOZCv5xAreru97Rf8K+RegErxJY5pPUS0vCYs2k67d/YRw71/sf36HMt
POE3gtON/zjUik1w7GfXTDaSN4RbmFdG3KwRhKplg02k8KybzOBmx3kzUm9szcgH
XpFd8z1JFlQrz3+MTMZOaR1E/Lgxkg6RZ6DvcA2BAL4QDtOvPFdXgQrYdksAIyLr
y1eZ97puwejfH5TOEopEmAPCUJ5cykyBGL39/NQl85UuGVX8emp0+6Fxope7hkOk
iJLTv3Dsu8fB36alf7uX47StVZz6/rtLm19UZsW5UZIBZ7/rZGnYU+Hds+a8RmAt
m9HqQhbNpLmmR5VT0LucwiWLOE6H09f5JIbM8/I/C7FyuEvCz1VJLKpIeGQAGZJc
vQXgBnCxSWHRbT+QzgvofUhi+yyazIiCuJJQEvSUm+fad78plmpJU+0ODxS5jveD
EaA+dKJ4qJo4NPpzi14dEnciiYzOudBbNfD01SI66PvysVLEcxT2AVl3oGmugOaN
wAxVCl3kGU+wi1h0IeVqNc4boM0f5TAUc+96f2gBJmS/gEPlzOJBuwfnr/KzuBOo
u6jwRODPNlmG6Ino/lIhe/46wOLUbo021wl+naDhXPC4FkabOgjF1aYZf7ElWt/2
YFGYEqvCTqaGmT8gMh1SfR/yKukjW/5YMKkBClpJjLE8SEjOaIiawDQKoOE1WcYH
B87vY98YdIa/TeB0iWRIQkYTGSsAUIJYkraVOwSBoZzTNdP2brBBm9Z+O1KhG3Re
K4NKgB8ovCgIXAQZg8uz1wNMNaAmlMUUfX7faO7Fk3TyTFIg60CGgLGqVlq+1l8N
OIx4I8rqqJgex7i1nfcbF7CLMV/XzuorIreH+BiBFygIRmu3QGysUc+4W9lWHhNN
NIPNPaplQrmhA75jBKITaKC8X41EIjhPb+wu0R5PMA2IKuAUKSCywv3QAJ6Rk+DV
Oe68w5wPSLeCX6bTNagFLtL3JTQBIxigmQq4FaNhSLNqhwfT9KQDxehq7fu+Tywl
0Aeb+IQvw110DrsqWn+X8GUlLa6Tt+ivv5pkJBTnIN2U6rV29CiOVz5/7mRIaUWH
MNt2OKdgaDhKwkH2kU/fADAooe1TSX7imeEWEbjcMsnfin7B+jM9LoWbHuEeELR2
fxIb7KiyRVtg+Tk0OSo6CqhPDuCZtKCrmMijlBBb9G8cpKvIvD7RChJ9fgkwXTl5
2DcDjUqISXprW7KGEpMf04k0jr5MMLx9b2L0+aeJA9fhPq9OtvWpI0ACjCvAg469
0WCblSlUgqajkbKZ3yknDfcgxN3/3TB+OZcNDBkmAgtYujnl4u9yvWVuyYb6eAmA
cQmP1IoL8g4vJOA/WqtNr21eGsDnpbBgJjqXnYJxDscQOUsg/bgNWII6lCBWS011
f6ZrU2R4BKcyqtLhlIOVyUE4OkBmdDFcTmYLwunNlNKiV5ackByAZTaFDt1+uhUK
l1QeOuCmMg/t9wsTvY1hIMWlZuPpoCXgJ9TXinpF9quW++j6Mo5hlNxd5+BhcMQ/
WiFOb5KRZvD64vVUZvF0r0G7YgGOswkg3Fju2kBD6kvciYgSq0wdqAZq5N12MhU4
5RC1j3IY6EvyzPUJqsFyirIOeDBtRjW5GD1EDYi/QL4spxqquVkd0nJn6BzzcDF9
DxpTXY4dldf9hq4ALwVqC1sGVPFBsIU8532eo2wZ0yRXzwjvUX+vrYzQWoc/6v9s
6BsEcQu8xkexacawG6YCbL+JQCa+VLAnV2jgg5qikUDAjOoK/wwlvrtCr+5sU/Um
G140SH7dHuMzm/lppkMilB5Ebp0lGzca4UyYpc6CM4cHLjoqAVJrQ38Pac/ROnCk
6y1e6iYkEqL9Y8EHf79kneTaxFnFXX31cDeexLnyuSmm+kEYy4LPhgpU/0KQSuxv
oOVnBarUYrk66zYnGXR5ANlK8CLPerPqHPK80qZhuPAqO3pQ5mV06DZfDgz/P2SQ
9ExgGGqA7PBkI54W5OTv4AdOvDKwB73YtqWLQ1jvg0aCTVQUFUgWBr11k94n+RaU
qFmavbgOV833KitXBaGZJ6wlYsLAKBtXafTJ7EMyE3rBj0VEPCQtK/oaHFlnw3ou
si86aZCkDdXMNAu0ifyXCt3VoXY7qzs/hdj7kkUw21fq1OGGbTJVpk+TmW8ku30O
eelz/J09ECtvg3RoemN6XksZg/wqbyQnAgiAcToABV1QZxrXU8Uan3dqO5zPO4Tv
XJ1kb21ZOWL44OxNJ17TMrF9mq/x17vP7QYyJxkm+vh5oecPGiolH4q8IBqk8QCc
2BbtzZx5ARsYMy7bQ1zE2ro3ZoIWENCasyLIHs7OpyhKgXCkSK9OcAZzoF7kSLgK
DEsxZ4GjRJARj5cu8jl1itdXhLeUZSgrte4kIksXdI3bi3gqkbVnFomMLSbwxER/
TRaZpIP56PoviPHazIbvwIg1vZmmnlmygRmJo/38Ix0y2a5iKqyvXTIQkftJYLFl
ZSK1pgIT/JPbiOYHwnnETg1KEZzpaZFoC/ycb/q/8S8p4puxsLjkariocvsr6Vzy
K0ac4Kd6cwXI6HePsq2N67M0aqTbIdvEJPoyNmMk6DDKPMzfdoQk4sQiA47/Ejre
0qJARjK+IfMh/YvYfqt/Hbfwn1KfO+Jnq57P6IKmtvS4sNTs7s734/6s2z2t2c/m
OdFmEATVJfSvmpsBgKnAyf8cgux8OzE+VF/6FNlsWPz79EaBhSBAxDHxb8yPN3PW
nEpn5DiM8z1u6ThUUTRnHO5GTuniFBAiauXiYyK6gIEdZcfVLdw7Ka1tuhgpGUZj
mVNJmsPcPtk4PmQzjhbVN16oLSmTkXNKmsxB7ydl9n3GnJVDf1DX8ardfl6Z4dw2
gB8gOJnoxXiZYb+7cpCjy8FKaR8MNbztOKCgzQiu/KpOm3MDeyl4nKfomFYkb7xh
2+JHDvXz4EW9ZrlbRZrea9Alts7B1X58cslylXQHj5JA3lYlQP5qH4HablGlwQHF
VS8h+SvCY67DyteGCwvFaPcGIy0yk09+ufafeU+pokCLUa740CA2zhK+PePUvANZ
Zu9c12zFNrcO3uteCUK0aeS4CxUqzf4GZ2vPgOgejzywhaaDjMkqYinjTVwXTOse
SpP5qFn4koR0+34gSNdFaQFziEBnWBdmAYvVIc6381gAuFzh0JuaeBDF+KTC50vt
mQ3iVbX6alopOzEbSnPT96gqCNzYWu0gQgOGNLipT+bMYM659jbnSRqM4XIgn+fS
SD3jS3awjFYGJWMGI9bGk1JtpJqW1yv0F+yUGjwDuyZ9EBXqVGT78tRO76/O439h
KZvrx4uHnbc1ikrZkCPsqwS3vFZXWqVAyjhYxKihJCZfHdubORH7gsvOZcsZ2Qox
wa2gKluGe12hkh2Qx9dOExSP6/1/B8TUKaD94D3tsgSvbEheXRHVR2hfo/6d8f2u
qqj0AAwKqMFzuhCH+VdZIkoSvOOSTaAjYmK/O4CaxLIHRNtJWfyA79guk0Azoh1Y
fPwk2eLWClsxhdUY8x1QT+nYkxkudQpukELqYwpM61J+5X+FfyKPSJKZo8xZCrbY
/gXWByw11VSewWxie0/KP77+uopQCF0VpfaP+WVm2p+R/LiOUZ0PYhnO2dpgSaRV
JNKo2fNb+tTkfD/fYAeVPrLWCV7YH6HFxBEnaJpDCB4Qw4uPDhwPbD8F14CmH70l
6OUoEgeiAwDjf8k+Qmz3GE/fMOjMbDWjuJTMVBK1wv6Q7qN6ebaK9da+S/1cgQRk
Y5vcVdmlROSmv+m8zA50/vLFCvo7fbniHi9oSrVYpD4s08qRxzJf1rCcY610tOaQ
v2qUiyBOrl01YdReTVQiQpEjLbnRyFMKpuX/hgQdmzCcoEUKAc8L+0FqtEvD0SK/
GDyeVd/xEyknbhXoZtq1qNBACFyjpaadQtHI3FeexQK8jXCaMgfFbxjmQrNWiE3C
Uqkj5b60QZSbKIR/0fOR229QLaK2XX6CCLkl9efo40t3FHgn3XZoV3P3s0Oq9GrW
g+DYTWvfXPYyhLsP69ODZJ/5UfJqR3EkFkzT0eXeoL0dvTW9TE0DuII1v4ZsHOuR
5EHVIe6kdpk1HR7D+XT08ABcGd4l0z7N5jkmaq0HPi5pkTOZcRK+Ta0P0rYtl8J8
dND7iuwOZrg+FCItvaeqbGoE78aUZ0kxICAIiEAV57tHoqAX+vThAoHLb5o2veHZ
BwRN/k/jVSDf2+/dcfmLuiJYJPbPiYmbzdINFn0vR9yA+TMBpBf5JhOYqI7X5NV5
7GKHJQhhW2yLVXGprrvF7lY3R5uSKL+9ZkAoQM1C0KJRMlS5djuQAeRr6dc0LQDc
s/JDQvA3++A9BGVYLKlKCsRkhvRSM6broYhYvQ6MUIrGr9fE0TLKcV8vTrqz/nza
a8wEb/UFPSdYNKZAMKMwokeSZtrDpZuyFp5AYJwQr6QYY5FVy2sdGzXhvkjpfpvf
PR22qBt2ylTG6qx0Z35j7zY1ilSsn5ppUW6U1DjvbOwHxFPuzfaMOKxzbbtHOlQL
rseuuEXPT40O4ggYZXjyOqSZ7F2sqajbiJjOLtoHcb1A3/2HF6+YFIdviGYKPoRg
QiULDxpEbmacXoELHK312NLwfSvgRyR/6wJc6QCeNsTSa1+jnAbglW/WZE6n/x+6
4xH/LmgdjxftOmXrXvSuKleaZKVgrOhmhxxYX0OcZjJzkucqP49Bt091Ndv4ioGh
dRjdJru/xZq8HOZc1QgNvRRIw9pjWfbH0J2x3f8/f9dx4nf+kHOThU7UhxjZRnO9
kIvxhaSsMpu5eYTLI+YrpBng4sthCYzXptkaQi+mhGikAe5jbjXYW2ng3Vg7nOsb
tVxC8/Crtu6r6w2zr98ob1HuqnpbBo7fA0WBsno0aItq/3HHZ0cacK0Iz3U5CZUS
FsqMjbi0yNe2AJtHgEEXmLgSxPnKM+qgx6mTfZ/SDxjBHd9QRi1HDFB62bfNXdaI
48I7Z59n/qBQdXaLsiA1U19l68HQ69hv8zoEUgIxgDQJtqPi5e2+KxL4WoVOLRZ6
bx8UPqmScFW6MQIjdjaKP/eB6BcoFvTXAEI4V4NWKfEI/nIteiXVnXlnCh0g+Cvn
jd0JItG0RcWacpIXJ3mmc7cNT4V+EW4fTuvxx2f6Jz7vHcFWi0ysQWQsrK/IZX0U
l6ewLuLSlgiAAMy7uKZA/WHqC/dLj7CeLDufRlRPS7KJvW1Gonx+jhbNWeY5Ne7M
pC3+LaP2QvHoNlTcbZct3aSIFslxWLW3YULzDhJl0wLH6XsBhmUQMJ+9nS/jC8Ra
2LLzae82rrePBN7725DF07ioB3q5gS2ZXEXWDHHyfjEgoDQ+MyqfcMqEnlCaeCxo
bNsGcswD2duTyzgw19lrASee/s/Q8qxiNhHjA++CijK8g7Kr0XzQy4YN2l8WggXF
qPWM65GYrlr2kYU/o06JkmzcwLIp1I588ClRkUjA3PpgoY/HE3Avr/QavCYEMpXE
qD1/EgxsK3+Nx8n0Sr10gQmI7+qa2vVTlUNSbs1NbvV2VaULauRDE9HCuQZWKkO6
Te/1Om2ebZbUaBVOL5GbN14U+6x0L+Vls1kUUGJQBLlak+7ZGcnv2wsprkvAHKTH
4Mp7sDlJtFVvAY8PhQxwYE3UsBw+KeHypWkajQmvllMy5BpoMmuC8rePJU3Pw90f
9eFw+1B5niXpf1DQh2LPe+262Wh6tBdO47M3syvtEUXLw4YIkRVSaDwSXpI3tyyl
pzj0XPQoL6R0Js5h40BbIjy8PqzNpZTVX4WGnoKD/EIm/kta9Ofh5+ZcgzfzLZHr
+TlG3YWonwEhvmFKN80Dg1M6/Cd/1QsjtCdrNbRntL+snp58s1Reo2/q6TUuGFCt
z7bwkoV81rtOMiMv+ruvnCHhqD65gMWJxya9UM2VvvPo25LE87uPCLDL0j5FhVEo
X5lvUx+PbXYbyUDrp6eInnhAL0H0Txl3ZpSDBrMVVdBmgr0rwu7iIbkIRrwO05Bb
MDEp9U2AN7EY6/ESubDveiW8JxMSmfrvxfQEJOZa6AQqTWx/9CD/J0Rg9aP4eQX3
sidVhxs0LjWo84R1wv4n6aj1HV5Be/qbI7C0r7EE6DstyIWpSadIrt5p5gBrGWOm
KsWcn+En09uyZVg52uTLBAnGwq+34sYOihG98Zy7IvoPOaksRAVPreTx5o8StFNP
+DqweTxBvdoRzKmJ2bE3+LdBfc/LWueRsPpfAMCmffHaR4OWK6qEcN8YNsj7pSP+
4bKraa6tGzE/rlpxj9S9CGjLVByt4QE8ZIWHKQheMQKtt8MnVvEORSoPuA/3hJTM
YBMCEDOS+Vq0v/phE6U/7jzK65AuhXzuBPfB4pyN8fF7CwFgcltlzuKGR4d07r7P
N3iW6p2RMrzM4IQTvI1PYzs3xuhLtuJttm1Q8IVNmkvuqy5gl2+JuqqX+5tVe14F
V/jrR6B4b1TiL1CjKlkZvuUyizcgJBZGcl80JZXecS76amyJzeF1j9ua0T3fB156
sRb+FZ5xGPpN5MESTC4XA1CiRtoN697aCAzWVei46vdXKD3lngKgKPc2VXCwAHMi
F5j6wAgJ8ir5tQpPAKowa1sVKae63CZGBCE9D2anxN8JHyT4L+d4jxDbnymPGmmv
6I66c06WQk+ki3/Ha/l1iUFQgEqYHD+J/uWMFRmxO+ymBJC4xy6tE/M0Bk8SE1At
q7AyjKOSPFvOVaX3DUKFGEe9ISQximnLEOrsM9Ob+lWyF+NR4534dG4t68NK8GGM
gaTpf7Ku9MWNlpJWRJITkwYXrrU84r0/Mq4QjWkE5LXfSYWv243P7q/ym0iC1zkX
wXqNiCegTTep+1M8D2rWA2Ti1L0tMgDt7AL/g4acnI4fzvScrjOHpSKv4DghTvdo
MnBmjMmQZNBrI1kdDaQfcp4OokmwgkmCPEuByLeJI+ELbwDJwOsGZk78GHA3odoT
m34CqOc1iTFk8N8uhhRautOUDeSZawIqNvNxFyM7gnuUx6dm9dTqoWW7I3KLcdU1
DDGnWbSl7DkzH3wkHOLn67wmtQU4wrmpCzKM3WS24+35EJe9dWqkQJGSQg7QSlgM
DEPmo/+YSRka3Wm/VfMrC+uxeD8H0vSG6WY0MXOsXsusHi+Ld9L/G5kgoTiTVWMU
B2/4BYuTjCCWpcAJdcu6MI89Bw810AkjpKqBT+t1vTm6CMRY28ku4VguZfIEoOne
ddqVs7Ekg4ur0tCGTrkctykCWM9Ir07k6jidpT5jY0oMkvXWf6JeElYX/B1KUDGx
mz/hc8G3ArrJQSL9q6HFmR/YHZDThVUaMA7ePGq7pTymMKO8YhgcNFfqWnajXZiL
Qw43LsvnVpk+RopR5d/JT8dRkXNvVnq9iXgsEEhrsHUiyqH9atE4kdFFbScnOFx9
I8YHv2QtYnvQ5lQ/CV8jsXaPHMTjknZefayPTjybwocZwcu0PSFroiBJsACFF49E
cWO1kiWcAvhlg3bsaA0yyv934gVohNblHdRR8UWMarkO2M/4kNTjPVBRXmRoY2dZ
fvwVkJsnL/D9UDMrOL7HaRj8dTi7JzHC8o8jN4zZuzEIsQPkD1or3EbWkc0gTZ30
fD6CoYhG+qET3eFG/CVnD2r9LNIf1SLkOI2MWerhzWrPnpfA22dsjcViyMg5TpYL
OqyYstrbGbpq8QbC+SLemix8R2MoCNSMnABuBEA5srmEQnBr6DVaj39mQw8jViNl
j+pklpoo5r9AjtpOFDVmBUrvWLKkFvNkutIezkq7BDaxSfectQTCPG7pdzZ9vMha
zWlgb3CyzexV4jmUrMGtkOsJe82BgqwLs+4k+y5eDqVjygPb1uhC2+8Cz8Zv3NNe
13Cr9w7FX5lmK+1zXqwJ9ds+jI+PEDZRmaAlQBegolAfeab85/GjsbS919PYjoDP
eKZsyE9lxhzkhkAV7ySFVRQLipFVEyV9CAvWBufCm671CAYyYkCLeLWlUsWzco2k
InngIsQGFyguopK9PgHvdc7fIxfHdBO576XpVOBeoF9oIA/sKwfXyzdFolH0PoGA
vLvHxRlVrz1ZA5ic5JD5mwSsf0Gv4AI/12vpUREU82Mtx2HYRHag6+axR+6owWWK
AVvZT6Vuy4Y6Cd82rQNJzNJt4MOd+H8ip2Vt6NKSDNk6KK2hvSnFdD497nZwCbbs
3OBwGCHODd0Kt6y060z3kPsrwvuHNDZif09vzjPSYd5KIGt+zP7ofCFqoaWhrFeL
jcudY5yPP7V6X1tta0jtqoDNayOW3elERtefqqf1ITCl4k7rGj+uQLkvDJfFDTMn
cgVh9dq/6SI0rz+Yt/IbJA9FRMhRUxBoXmR/NoZg3zrqRk23LOtCRqrDr9Y7hnU9
UEA9LbbYHoCt7ty3c9S+yX+wPM2d5M6DspX0UOLJkoBGxkdhY9qMF4EDDV7BVslw
Ixzq2ayYe4uxN1FklfJh7BrkWDRF1CghySEPa4UnAPtIDG1xN4YLK0e7+vd13821
5mh2nL9xhNyojpUvfJEfqK3d4I3BYE34zMyMEHSe1YtdpVQLDrzioDyzPBz04Lfh
T6H0l/zFivKlzwfJ7oKZnRwmrZXA0dsCwrWRSOAVeB7slmV2qLf3JhdOxrAnvzWc
zqFlDOr7PB1j6qFOjLLrVYyytOsDyFQ5oZ4boNBavCeQbGd0c/DYQ862AFX6qPOg
Hd2JzjZ4v02ZV/ZGXQSB2OFx/U87xJ0+27c0MKYQFotwffYJndAmN02kigd38y9H
DzUhNDa7ibB+TyqbZ9VxXmPiGzQlsfCchuVfJynayZbxVXAWRR6UASsbAHo0520U
I4eQzkRa17qABcanf95xI22JWCxVXpVW2h9aN8+8awTDV1PDqquf6qbeX37Fvie0
ihAkO9mV5/ivdh/keEGPvJaTylLxf4kTjSJOA9csCf+Fo3jRZiErVa00Q9afcZmD
Hbe05LYADuHObTkFff86Q+yYh6VMEnEehMnEdJG/0peLdXLRu0AThQdFPaxmUEH9
wXoYg9gKNlhzQj7G6hFAyHmUU01OY/he92rpTL1mSzqDqAFVCOAdwTF3d6b3AugV
0Idrb8rmWkr+EmzigzDsT3MyLM5l2QVW+KBC+MNWKgfcDa4rLa1TN/G0WHj+Mim3
cchYc9rmkukoA/bRmDVxH8ZWdAWJ3B51l213LCGTEOgrKkOaaDc1GS7r0WczU3vd
ZwjEXKZ4CPENpt1wQmUitBneOWiP0QCmC7p1M9cJin3Bi+/LRmTxgD1AjdaBb9TT
Oc81k3BZpWExLXuAEwfyzgWmzAVaj9CS7eQtNEqAbwmWhyQb3VOh2tvGZVI3RJR6
Avsvxl+IwxrhAL+GVL/vkTiBkp5EZwX6uch3DCHLoT2d1LyxU0nLyu9JkCobPsLL
y3WTnbjl772VTq8Zj2SCyvT366Ffq3OaEnU3diCLCa9sv3nzOSLLpEfmhqJVLWzP
sgFIrWYQgPcDzVy7QJBbDS3hQj0+wHY//gMV+E9thHfb1ybqw56jYFQXdgWyySep
dAQw5XpPrQSdIceTWjkwAxwm5hgBthuuNHeqopv/ZhX93/0m4z33F446cNMxsNj8
pgYGD7lfieQPRUfPSbySUIys/V6ljY1ldQPPnbBRhchv10yHv6Et6QzR83qk7DGf
FpYwCQCmERcIVJWmGYr6/zd3Nm/EJgAei3lx3uFSCYeT6IzaCKTQO/uk7VJe1++E
ppmRYKGbuUljqrg+dxMmynUM4kobcXPeOu8sa7HSZ9YXlyz302fmMz/HWKyy78FM
Sqgf7IY1MZsNa+vmIENTCHvlOZ7n8Yn2Ylm1K22ULeVjjAN8LICCekjFKY3DWVu/
y0HOE/07c+0onaOo79naeKeN4oXznIQEyVzBlePZPFdM/sBOsOjp9PEnpiDltRqz
dcJullUvWMHalXz+jp5XuwfJXeTL0iRsR58sRf8KcK2A68TM1bqraS/4+3s0ceKS
dWe8R2miOsK43kefxkIviBYCqZtpv0yQKfvvftaO/034yVQNd/I1z0tjOa3ut2oX
iYT6p8//kqTpqkUghIVnSI0LKp8ob7HhHUlSd2gDXMz9BKC2R7Zpi15Wv5z2NOKB
GSxXtakDDDIu0goFktY7i6uy6zkY3fHf55GXGmBX7sYrKWUjIKzQfnMmmGzI4s+Z
AsvZCBtnoxteG/GxJOzinqdD9+ZcUubFiTyR0Hi0vjoImx1pKM9y9GySsajp9Iz2
/BG4aYJHDQjn4mmRSu2FqUTK+lRmjbSppdZK7N6K3St6Kt19YrHIZEHy11zsFpo3
CAUx21SAirZbFQ6+m6Def7mrhmLjuEB2qTQXBagvwR32+Ww3+J1PTF+bGvPLFrpp
8iIVEPuZtXe8+L9nCUYXkPUthbWCO5m6zCXj4zpwh63A2PHqdwPZk0CJ4EryT0N3
drdDPuBph4NrAaesidwD9CrZJt+DbHr12eX5bVT68pdB6lCfKidUDcnMb+ZQ+HJR
mq/M5OMHFLS15uPrW1kbc1Vihjefuvp1TJEswiFa9z1tcTg5lqxI3LEwQWfxuEIK
pGHFw5IwBsPU0wBMVDkqoLWDmEm21hpYSCuXcjCIqRNbOmjWfF6jsiEIoG9ORGtX
3KiuxPYWnNUhWSekU8eJEu2Mb85gU4vcMCp7DUeCMJfSMxYJNYYlhyGq3HgKp41W
vVhCBDrdqECDyexvtsIintbKvi7R8ihTHrVTvfu0rgV+5Mwdlxc22yr0/25DuXza
C/a29DwcDVBq/NDOTZ3uIwgsP+k0/oX6gvO3brUpxGPKcyRiD1aJcUjoOATawO7W
eZ8WaFXxEpUSpMMA24pwdE3mZnaD52svPVOlbXuiOFgto11tHqeQsLMhjxQJgmr+
E0lv1OXQ3F4IXjWUwD1dQha7DMAAodQSpqpCbRCCP+dhyDAxk0R0oFfwoi7C/Vrj
ozYus6e4bIFO9zF5VWQ6JAKJGnJvAudNAgF5iY1L35TXK3tQ1RcMuvWUKNlN38di
9FEuO2C+lQq6qJL/o4X6ndAhIpp10nqCz9u6943QhX5dHpBxUyIu6uX4uWFw2G+0
4d/+CnUI3faVIELvd/4STt7SuvoTx1NZfpKzPas/W9DpoODxHGlceY3PkTnsQJJx
rjLk9h+oSgHiUJ0Sog9gPEiJPu5dtbDb4csfpHt8zPoeZT2uYFRQ5JZPxgA0QjqB
QCOobDlLqQBTOYnsogRJsf7iDi+IuhkSYKL25aG0CGBI2alIXCAD7l7zaV01EyMw
2Cp9fEyxkoEG2CFKfMU+hkLAIO2PI68V3Zrn4IdRNKa3nH3YkKX5r4mwPbdIcvZv
Hi+uH52X/KTN0tbgrwLR7lxtdye+s6bUCJmeKAwLa/6sA7TQASEDJR5a9z/ulfz7
X16ELCz/9h3svyAudV/hkhbfWB0N5zarU4ZikD9E1hNI1qhxu8GYEVv648u630+Q
Gr/2x7kAIxd4vOPk7aHNQYqgJhGs+V5qiwi/BrPnPnnhdqvhCTYbtarjYXwjJeyA
RN8HW2iwYXNs6fBtn1E0L8YFEAo6ox4GOmTjQ8CMODBwKrbiVu6uGUqrUfdqumZt
OwDnZkpHqfldZp3pMapVedAxvQgsOtKFqRj0Znj+C3Z3fHmXJk3McYo/stZCEEUR
88CG0j5PswKOIrOxPw28X5g8t1ymc4K9gqgfnl/ci2NAQ81YrPuU5RzharMUwwTC
LQUbX0xfGPAbdopowt3lX6422pMgFNTMoneq/LCYytCbZEg4o8sC2Wi3aXtcGmKS
GeD5EYPDMH1lT4d9QfAbqkbMb+q3P7Zbp+/eLOECQGnJBBYl6PYOfbhIY4CsKi+L
iQxjZDDpxOlWhxV2DIGNFFuM5NmjRTR2DX3S8bo744lC4jcD9uC+/QZgahOUGIN+
fOqk4YoOWcXyvUs+et+vK4EG6c3O5anx6c8xToszQbUKqSbNpCBMwF6WgrqteTx0
H55DFJLjic2mWLT8geqmjAlNsjFR93CIC03vxWJ3UPsPyGSc0bX10QJ7WVchxnMn
EP8de0V7O8pMZKlLx4kvOAyl8p02wLSsps5aqEHJEKaPqZcYQk87k1+8vqrzwLgR
OwoEf9ssWD3WadwOXpQFezy6zIbUA0uU1vqK+KrtfQsIR176q2lu8Uh2Py5X33Pr
1SQxUXsCfP90TyVr2t+6FDPfFYD3uqstIVOSSw9bKRo9/e6BR1p3hByXxn7Ktxk4
B3Zqfkt8yYzFptctgkbr1T9DKhVlxVyEHdvErCForPuQiTDV00LlcfYQMXb+6BRX
/LYRaRiyWscE9r5q16xu3tQaYPcbEwmAV/LVrqmfkvo4rFp3jZCdvLvz/yP7y2NO
CFpFRI5mVRkpmAnsiCgkFDQBJDCw5rddnyqoVG6xwZIJhGXgZUIk9Sx3EoMCjyYo
DgQ7OjUygBT4XsqCitYV2Awx0wCfrDr4akAVhzOGzCD+j03yp56iHV0v2tOxzgYD
bB5417UF/StFzVOZdAUwNbkJBSVlATyXP/DpU3Yqzqi+EBqOPtbEhN1DNPGrkUUw
wxPBa81nH0OFvHYvpb3KAvk1GdOjHgdwu/c1TJjivFf+/K1IFpvBABtrnXzqs3mp
UVio63PQeZ5ZuKq5ZOUI9JjWxicEl+C6yWG6K5S+YoOAlXI8hE4qqGlAI2rZ29oC
OET0VB/dVyDxv5KNUPZuInDFEvULr9eNEMcbgOCgiYsml0uPYvK/cdSSB97aK19p
lt51xyUkandpdjnWuv4GHcLFOxJajeSVP9iQsUjVqsTiVhppu3+tV+kjhHEeEO4I
79zqLqkqw3QIR+8VQWMpDEAmTUATnVjOZmN2mUBn/5RR4QPAH6vBzc3AexOWFGgK
TfGd27U1Vk3dGXckwi8SPI8NR6DLtpU2+DnGevNi9WZpOFZFX7aZdMhqXGjSYTYM
LR5VYXK5Gf/j80led6yW/fL3LOUkPfAn3KwdLPP6wDgyeil01CT0uV4jZ6zS66te
RHIwkbB6qs1x7oG+oLHiWym+ozu7UsgdKfjDcUXLUErwQ2K+3vNJYoTPHR1X8Rqi
DRMCWCK8Zy1elg9PNvWO4NIygkC16Xz2VD0psumn2BmEMrYPltAdUtdF9UuBi7yl
oPsT3c/1Kz/OSM5ngwMie3xxjIKH+Tq4oR3CLxU3kaglO1Ky4S0wKORacRn1fmHq
2MV1IYT3iFJla9RP27eeGQuTJkKVxnro2w2sSXCiBi9E7RBVF4LVCv7YzJ8kvxFF
m7QlK27GnRtm31uvafMYBFVWQ0M+5cBiV2x8BzbcbOGvEEYNVFhF1QyGuZOKBmVP
2uDFG53Ko+bUlzI0tBWJZ1rHQVkT3RZxudjnmB4cIeT8MBLWxp4UXazYEueuL99E
vs6ool29rG4u3p3XfVXqV6jNCWeN/Tr1uBEhb4GnR9dCeESl+kHwYgHOT+qEeBIz
LQCDl0CzKsub9FSEs3lV+b9X2qdbm5NEcxnEsuIWXJulrY2+vPsRofnj4N1fSZGU
sP2ycc+N+00FE89PK59N81zAwBQjB6xJRt0HNoptiOxMIJUP5wzL5ckm/JhFkYNa
F15u3brSPjkdjfrC0M+XWP8sUi5yqPL/l02vE24eBRlOERj/mBpo/5guucFJiZfQ
rWgYVfTODprH2HiTQwzZx6I5nW9O8ofXYVYKKJWBG+qTWH0+SQUs6YiCKmwEDcUI
IsdhwcJ2MFmW1kJOIljvElsDHmJfkbJoZemBWxgRGNiEGQomkrDijwV1cbzsGf/l
8SdkAlYaRMeYuJslGE4L27Jsm0snx12fBUmyw7B77rtv6PBkYo7n8AKJvuyaivc4
4BR70BsX4rLvj/LbS5jINu6awcxXB/gqeiklKMXaZNt/dpASXkGZtvA7DRki0n4O
0MCFgZDr3XJ7A9uSw3jURNyL6f+JAoZMNHcTUc5Zx78HQa6gMdT6gPVpdKQidJyI
8Fb6H5wTcKJi43Zy4V2/5MwT0BYlPPDY6WwisNxp6nTohkmmjNrk6G225UdfrNU/
01L/Uq5ljoE7DXTUlbU95bFaEqGHA9jthu1Q3fTTRUnyfQGPgJjSXuBQBEHGmpbg
/Gyr/T0RNnD7INSeEK3EeOJaBZfG/0tQEy9yNBMk3eOgP7QXok66Q+IZABWGm+Id
Mvs8xWODVPrLdK1dx6F88lbiypMiKGdUzFUHkvkGR7K7kzbnYNmhsrSfmPu/HB5E
3fagx3C//oZneHAGlFX78tARKbcKYnO/kJvwML/V58Z1URfj6O7W3JSm9me1q0e2
qUFllijsfGBGRmBOit/LV4jxOCW62YFeskkFgo6mpY2BaYJJkdHssxFGu6UZwbdJ
G9S4VSBhdmcbczmjAGTwoImoE6eAoCzkcanCUFYkTC6AiXE0e+B3IJdfqALJNmmn
6z11hpL/PCN21E2AtT45Y4u9tal227KIY2IDXTM7pKQq33DrwVXdsSEOSxH3ykq6
fWbhxIlLaOyUIjGx66nsxbWsCMWtyJ+/3lrnj+iI+kC4QpAjcI1ALkAPjv2n1PIz
zEHuUjdG0f1t4zgwPk/OqQWa9aqz8OADW0ewy5jrnT4h8+zW+AEYtXkQP27/Yu8B
FDvAZ3SKvF3nyWhGHLilxEWbcPQIyIzalPI0hT7yXR1jkUKH3AS3L6dgqHhp/djl
ZUxnEAHI63hUSVtnYDNdVJ/jSNqox5cGnD4ZdwLOmpaCPBOL1AYmb2r0vXvmrFsC
P8EaGNp0/4VeOBE2ECTy7BcSYP93S6B8KwZkALUNowsM7PH/bs1/t+KxgNp+Tbfz
vvRPJHCwXtSoMbdIE78PTYK3syu4WtywbWZw76TrirxpwdGee/DJr6Vxux9enobX
9tTfrtemz5Gg5k10ZQUYi98dYuRpa4thkzU+4sxKcSk5UmEltUjUm2g0wkxN1z4X
DRqktmRX25+Q3pAiDUEeiKvv8rvz57TfX5MX4mZotXDYST9Sz1fbBKIoJhdZzmpp
mKWFBZIm5swuGHk2Hz8D+qSUIGvX3VOgBC/zNSNKJ9c+Pwuvtay8faRbEVcn+Rga
Ht765Tu6SHNxHHBtwZakfRQ4yz/wLwxZ6+Dh6qEmIWm1m7d+8ffcqhQw9C35UORn
DkKwZS/uqMsrs5bFSwQQiykU5IOMX4fq6/lV7kUNU2ijyINjiOGPOfcfeS91YLGq
lkpCCxhvs3rIFKCX7d9ZjfxwrLftBnIKVznEV8mpF4hfBzGF9S0IYdBZuxuaXmym
meLem+d3ll/xztLx6m5pGgp8yT7SdaJm/Q3hzvfMFjmaMTH+jM9E10mHUWBFQc6+
QhCD2Ql5n6vlTKtKOUN5bisuRj0dFq1d4NMGKBU8KU6E4nKuQqmspFs9BtlX1Otz
P6ysdKCJs6BrKHehM1MUcKcH9fUvZlbbK4YxEGpomG28y8Mvx5JngIoGnPQNfgiq
BtF/nmLnulJaajG4dnI6uMYxSYgJ1CG6xjPz0BTJLNFAcEWeG6MR0MysOaR366E1
V3XUNNgsjCA2rmfIS1nTk9bZXhAd8cKxbQztaD1728MZEG45X0EmAt53au2wsiQ1
ok1fIa6pvpPoEuIGHbEZSNl77Q7oozwbDBQoVz4bPez+qqlx2nhCFHEWkoS8dzXx
tVKg8sFtHeGwS+2iJK+E39/jjL4f0i2+i01ekC5VyXVdIA9DLCFEAOme/kNmZmD1
9eJGtFeQrTFdzwzSrmOrCjODHd5YjW0AT1+2AIyNfTI5s+siSUS++k8wa7yYRRd6
zQ8eDzqoi0MANY1UuOWmA6w8tS6EzRm+lptV577HD2cDBTUxPkd30sgqWi8MwyIr
SUrzlu0UW5ZO2kTdRPs0TEG3pew3K5yhPLweDs5wnpTEsDuW51tKg61vMVpr5su4
dMXoMB1PVvSVsVjyMd4JV4Thega3PqAKxB4bij2Dyi3wOIKu4gyhtHZcgLhCYuch
AJTPn9OCQ5CspgluHWhx9DAb+ccR0T+54yb086kTeRl2/90J+fYmoUYD9fqjl2VZ
NaptqzB5TWbDu8QGETmyYI/Iz9OewV3aRVtkshFjFIoMXLdRqYBen71T83xfFaJ/
ShxVSQ0Kq15STkSrA2hgv4KRUud1a7FEh1rt1sThFRv34X8GOc1siwP5s3t9VMpR
/QFN35lqY4HboX52BIl8t+jTD0GmYHboaMoURqMC2Voh7AVWSEWghO1vJwbF71j/
8ODyb2OmN6HXaSyOmw/aXiGSOUAH7ijTzdkFTcA3O3ZR28fyjz+UY+C6iyeCGbPu
RCZwbWsZRAlTlT7BZdvpl+6cAykX2X+LhFq2c5VSoixi7S5N+FL6/qhlLK5Eg+6W
iA4uvDhjQIabPpzJcQRmt2CnsjQ5tRh3gn7KmX5H4E+UJOLCHwkgDrsmT7khnuYT
AglhdkvbTGnYcx/iaoZ0CGkPN0zxEeHW/tbeqWUSksHjC8h72QUfycWSKLXNuhgW
kCVm4jqFLFaBTYY04n8dJbSMgMJH2maKWK6Sf9XLeuwxPTQHSpjYvtSEpujkxHjj
XAJw+TgPQSSTCHrWU3wNwuGznxOyqQeAdmRMihjMjeQkQ7RLkRmpKDzupQLGvd/O
CLwqqV2BVINbfEcNF1zulXYllYyhiCCCregyG4p/xnBTSP8DM1NhVXVY5JXmSeaQ
ujISS5xMcoHNUCB/yA4HNxZSqLZBwt1JM0+YpofOLuUVNwO5pRLW0PradS15m8DR
v8wd7eFc4N9M8ABAvYn0cn/3geoMzNxH/0yhPjKiQI9weyad1emTJYsAoN4horf7
yAj/Cs2SuY5YA7E825ISkLwD99Ds5RSocEnOyScWPmOCaQX1q81nfRbJM0FjImxw
RnCNa2bT61DoyvNcvmofvgVHbMlZLofsQdQ0nDG4CYpUdBiUQwW536bRmERVDUGM
AIp/4g31OzdRPupFDusYfZbYNiAS4nDAh0vBx2pYi4pW0wvu5/rzFnphkkSAMKgS
dZlftAZla4kuHv94kTkxgRVeDRZ4ul7KRsRuqBn4ZYapUWe6YVjfZJPGfeF0uY7a
6/Gff4bYLu5bSzTzcIVzYIJHXj688YE+T4NSLfgE4TAMTwrQC0Mbcr1j/bta/+yf
sfnL6miXhxg8Mx77J9E4YmultmreogfStDvtxuSXYwdkSmaCS6ALBo95YMsUka7d
tXFPtO+lU05BNTD/P3cMhS3A5VUEWNY5+HOmETI07Kyk89JskZ38yk2Cq9nOOyDR
p0Y7csLci+Z7oDy1PmQXb08rOjlvHzYdzkOrjpJlhkZn3s5y3jbwELgrHO1VhGGg
5RrFdmwOehXwqfZlFXOCgGOE5OtY4xuBbnFkjadEZuIub222iz3qumm857x69ijw
wzbeB5+OGrCTVZgXZFoXOIpnfHkhq10TKoloaop0qjfiyLWUaQRDKt/JPtlgf8GF
8F8OHYNyLVtXZbu+BX0jq84j7TwQSm6tSrxnjfQgOyg6BkDaPZdkaMFJSuwKtKia
+reXsEAlhA2d7DTpYal7QKfglMBv92mS0mDZv97DRBXz6CuisABaA68cVCN4eDLl
N5rJwKMgX0oO9Y2ley61Q1HlnYAnEzogu8oYqJx0YOs/97VoRTI3tHjYRDmQyYIY
RyTGNlZ9GoKMcZJ02WFJgl7XbhMdwKR3STOD14rsBDt0rlUWR3jUIDdJjq1HHYeU
fH5dLRCNBC10AcRxZhmrfRbaNGs89EqOd6WSCv8NC2owvvHEaqfcClezllVDDqyM
U5C7KEgt0EpX+HkUG0qRcm6gU6MzZNqgAscgMg7VzAd3IodsStY1NP3oSbfI8+PO
wjGrqxcrRskpTYtnLOhip2QavR/R8BD4XpmUM2/KFDXjFonXQ7NidsUCZ4uK6VXv
dWmZp1BZ3xh7eM2VZyJNPyMy90K9UeBEXSCqC1Z/fbgdKvKwE/4UKO12idOT++Wb
MJWrVQMaqEEDQamIcsSa479U4YBcG8Y2rfXklaJTpJI6SdhSdZrnVHvC6EpI0pxF
iInmQ1pX+LHcaJENfAME4MebuDQQ5gpcWxkfGtGzQFIhE+Ya+eayDquBxC7yqdO0
XVt0j8552jB84aiA6AcTIN+j0iWayKC/CMudFth9TcwI5S2ni9b4QxXfXcjmZrah
OtHbJVmBPwUuGPmMcFse9i1GSiJjiiH7m8NkResmspWBNjD9HMg58tM9FJu25/WM
LVrr1y9aQJLr5CWfeqOonMjwp6C2K+GBPolH6c0csZmeJAYJ84gvzV1rlYnDN47W
1oR6CPSQM+Xu02q9Wf2J+fbJgfzmph2XXBoVPhi5Js3t64G51EbIV3phr9AGfuus
TCnAiWKzdfNafe6ZgIVMy0lSjIw1M8w4UupyKlu2YMV1wHoFlKV+/UlbWd576gbm
yJQ0ZLXoLvcutvmhfJKdMgl4yoXnpWhNngmkdXIx6Khd0nvjlOsIorCokZm3+bdY
7V1lMYZWcGmEtRCvodoemsk/RYrGRC/bS2qd7qHMUfv5zOtLBN2ytEx3hJ4OtotM
7fpEVWm1fQmS64ES0PxGwz+5t7qId9+Jq+QXLBxfkIWkBo0Jvl+K0bb2hFGNffxX
C3C9FECoVawLRMu7Zc6bp6kKP0xsvlguYc5/P+EfMx7v7S0R/wVbE7NNeCI+LRoP
1Ak6rOxRD5HuTLgVnjr1Fx01v4T1Qv2BOHNBRv+apw/ELa9LjbacfPyPxCfH/q8E
hrI1Y4zU3/FGsO1SWgNzk+KkT0sql6qRYeYaf+bnqY+UyTFxTXzgWDuGle2Gvj2T
ZHa81fgVk1CYaC+X1MRINk9NU+J192aKQAZKzx8HCd+n94DHGRwULEFYKH+bTLmX
KKyB2AA7hhsmAuks3VrYYleZc4B5rHUJ1SBF4K903GX9U0RB6wagyqDQv0hFBaQ6
C9Fbp8wdFzSfzyXzOXYfwRk/DkpUSDAF4hx3jCF/Mz9zUpraZG5x05QZ11feOa3m
GJ8000z1E/pq2Zdo8wCUe7EDls7/0wRbC3vHsvvU+Ta2asjDRgEwx/8VfjMpkBxh
MCGivYH/gw3Brq2uZ6h6kq36h0b1E72UexBUgE5RcsW+mulT/lJkEW+esWBgP63j
NMZKeo9j7gQusU2WfacQUdnZGS2geWVakgJc4jA1Kg3zx1JTNMBs9r1Fx4Dbe+BV
LiJxc1M/MNtF+dV1iDLGfoE3rNZ2EY9zhpLC1jVcEdGI2TWsVyV6wK1MsvhPdqfH
9vt9EYiHbmTBm/LeiqKN51dufUoKRp7xM0WwF9Bkh+mPXFrs8bmyx/QIuCD5b1Vy
73rf9hCac+TmPHy4R1O56sjdODx+uxXRzLBz+cdzi5KEQ7BAMEfT//fMtEGy0sMU
AhxaSRyK81CM/nwRqLyWH9T0VsjpOe6JKBe6rg9SIov9FI0bw/ZzDbE76/qBk+6E
uvQlQpZjmKqg+sh9rqZU78A4SfpEZX+RQuYUW8KsajTkPzM4OIstBbVzTkUq0l7S
9p7Iz/6C9AiWEk5QHnxbHbBFOKi6ubsmQbvAECe4Tm5Q2s5X78WSIcNobrAJ7cHH
q3rA7rQN+uAcd7XkYgeRAbKydC7fYPH02dFW55tL9gKQmG75SJLi0mRGV2kUjgM+
pY0kFOueyyUhQnlskHDj5tKI45luUz0zrFgoaPlYEUpKT2JQbZyqSFf29/Ye18J0
QbYVTgtLrA1SCyt74Ex3xs/ryLzImnbT7+xTv5ThFZD2xWth7xo+KTk2n0thURjX
CN/SgQMhjPb7v5OutrTJDB3PyEbyty01VxrCxBaqHMnq/Fm8jymH9ASvzFkVVFyv
l5l5UN/00QW3oJVx0X2STDN9r9dsgJGujuWWwgO1EMu4xgKkmUJ4GSOqHH8WI5Vk
dwqWFbgPrSSDgZqafeYIRqZf06PEBkAUtwYPvWLAg5jn/EwGdbFOAfJzgVURwG0m
sp/MTluyOhrpnNlEsEa0nuyS55309QeyXmL9J3t+pYy6gs6NoAxWuq14pNMsvYXH
TkP2t45EdynvWEEfY/8UIe9kG7gspqUJH3CpwQVQH7eFgnhqhKauDBTRj5hA9ANd
2FBdQ+64BcRIKxmzXF1rsu5d9EGk2Q+kbued+y98SX5UlSvqSAm2E9RJzo72YCR7
nIbj9wTLqZGJpz8G1kZh8/ydAgDAD77fVYyOfLfM9gPbpzs7rF+oA//Jsxb5XihP
DVWhesIgbrmhy6vVsyeQbhYVaDpvIKEH3dk8D33CPHc4XOY5jJEKFhYo6EfHfY+5
eTRJQp9BXoEYIa0yS67DJHYdGQ3/qPBWAbB3PGoNJUyKPOlRj4lKva3+7uhgmNJN
JM//nC897gGPJZX9pg0gN7djAMJqOycjC+td/5aR1Z7rMRI3peRUcPVeLqh9Rcw9
r2ncbTWXIbBhOYCPUqUmuHMu8LFFz/o3W+84PFEAL9Aj0atEgWfg8Z15kIAjbFK/
tRzRr/5b+ucKb81C1AoMacpIopS00wLYnZDmTeeCmZnX0PeG23s7FIpTCig+1gmO
v4J/ry/Hgkp2zeYODRLsuQJbiEaAqT7dDr60e9l/AOsBMgfYDwu6ikjwF2ed2mm8
7MybAK8g2A1o0X4a1GPNd3oHlnPboMkS9eEqbUDWobUG/nT3f0RjO9HW2WCwMlyK
n9aWedByu0FezM0kBkeRLFfEQHkge9Sw1B7ak4hkGVQJMODPy+V9I8/sch/1smeR
A+CSUU7WSi7vNA9gWr9yGD8DOAUy54PssleYEBUxD9qwIyM1sSz5GzSYi0mpqBB1
xbq3j9X3Tbcec+3VrFZUu3EAXOp3zuikyoNRKtSpC8ucjssKlhRACMcB/cc3QBGq
jOnf1KAy3x9yHOjlJKEq6mIK3ddvRmM0EtuXS9Gh9jtk/NJaf9n3gpehDF+gIbCF
I9Tpbtr3Dgf+S5sgyy262BjF9vp9xgS4b4iXyLG1HemguwnlN9ZWASTgQWPJVz/6
Yh4oIh9M4enP/wjbjI9MTlrizOHnV7gtn/t26hPdxnqZPekLWvlWoPGB6Ce8hBX+
h6xumbfKKzxyP90yZx0+RhksgLVbkhjhQnZaJgUZU2WLrxO1GjcbsSiV7D/rtn4n
Y7Bpf5HDd0L+DwQUbhvRiHlLcwd5Ax4XzC/WvVO6HJCztn2TRS+f+VFz935R7ijU
YNl0h4lnMmxQmRIY5OZlS/ODcb29pySFYexx/1Ci1ubRVzQwfBOX6l1vcAG9/MzF
g4GyzSe4g0BRPxYAaJQ+k1vqKFvPegbsMQIdLfO/+0UOB7X5WQBqqoBS505JXNOJ
dhpx0UgbnjbCYau7+wJUgjVr3AQm3SmkXjmcOm6C9/3VHrDgAb3di049t4omzb4S
QsqJ5U062uAGDvkHG5aqPP5elsjsQ/db+IkbLpv87tHTcXUvTIg9HlLkr5Z9H7oP
0BPoigFq5siVJ1m2uBZXhsafN67YAQaR3WC6LroUWr5NNLm+Q4ciw5KrGnBMIQKd
PVvq1kDv4MZkDKMsDhPgMGqRWnELmfMkrIfC3Ym4enuyqoC1rmcBIFShuePGg2w/
iYUPHcr/YCzVAPRfnHhvHpjv75FdN1+uKkiT4+QuUZebCE/q+gb14Su4/rUcD0SY
JQamE/g2SkV2UhoTUHT4jHdAoC6E6kiafFwlt8IVUvenvOgROgOkMZCInmbgBFD8
c3uwwZ5I8Kp82+u/bUp7oYD3+/CCCA50B7GrwX4MXZIxy3yTN6x0Mqly+i2ZD4ik
5ww4WbRdRU55uJl877D3gN2vQeFsRYIogiN1VV/3ZedSVGxsAftjBfd3LlJX61eR
lkQrqA2j8QT4XY+K/LryYhZW4dNvIGRlpxuIQ+uVQRiLjCq6GlSVXChjH58QdRRh
ysoktOSxlG6NkJOiJo3wWLhJnrDRe5b/7+QdnnG0IzcRmLS4afI8DvWSKf3vmQJ4
IGtq2QGdxB+DnTLOVNOgAq/nFdnrgOikwtHthEoSZQIfnHbQCr5qNg6EJKbnHdcS
kQ4uhpRFqiaEAqp+6u82Ry4t2bl3709KyOFRHibq6b7DLWF+PAizHkUmKdl9q4KA
0qbHI0XAxu8tXwT+xluZDQ1T8P86Rq997XpHA+faLE7p3HtxO1Op93sNW3gY/U4r
IXSyqljOMaeOEx1uMhqQyTntrZ6ZVbKwng/PaYrCG0MbNG9iu9rX8vpxNDaqv/3r
6vtBj1DbLM2Y5YZIi0btUtQmHUS0y5974fwkcNJe7JxvNTC4X6U8Ub1h3W9SZ4O0
yCaHDyniPoCDTqAfUX3spnznjFEGfk/r+ttXFjvHUHU+ZcQryYYb9bCLJW8k36lE
KmLoOfYMWsDHh1j9l+m7BTY7WIVyyZkAnH4XnZjBEQZ/sM8KiAWlnU5dVggKNong
Yrg+r+dfOAmgqmHyJ4s2BtgDGcPVCZIjckueMoqfz5ZnzhUZJI+++AkxAWHutvL2
V1KUVRWxDkvosROfp2cxetGkT2Tt7X24mgaKQ7KksNWqb4ELQI+yor7oLDAxZ+bQ
zBTKYkMFYIxBJog6QeA/1jgyPklBP18iOx9GrQviUPaYVOxsoIbewLt7oZKG2peE
CQGVaCP13XmyGP3tyDvlyBc4ro8InTYuDnmYhTFpcNjKPuQ8L2hLrdwMJzjdaCYc
ASVTpn/gFGso4ocHRC51OZPOG6otPsNAn++RAZuC/Ft8oHbcT3kCtypnrLNK/AWR
+ZPOds9SrxvTA5cXrZZgoYb+4a9bzhocG1LgBwS/DojhtycIwdk1iwp/8/fbsypj
x3L/b6hLvgyTfn0FtG4EiYD10udQq68/ayzN4w9RiTyj6ZOjpbHJ3Li9YskrWjVR
a8lseB1fdEp0kQI0N3JnXSryU3PNXSzSz0NGM7wmraGQQDDnHlt6Pz8hGD03NRC4
G4wNAEgO6TgSAonHozIAGs6Hus/ureXwiMZYUAk61YBEFFLY4PwrQO0394ZMccmc
fv5IOXtS0eKG1DUMpYSCR6uzxFr7MewjTtVECZ08fUBu2Dn0M2MX7CDz5irejefp
nsdPzPsZ2pe3QYYsofW5DlpAwezL5wMWE6zsFiHuph7eY2yELnuFprfWCh7kaf/K
kHh5/L57Aje/yykRUQV8p+FxMQfuvejFzVkFR/41162SDEvU/aureCfqMyKwq9dx
PSj5HYytjCgNYzHifT+3jwQO/St/wZLWh/S926XJTV3CM83kwlfp5tVdqARaB53v
6CgirUoWwIMz2RRxsftT5LtHkhTovP0Qd/5gXrDsRvv16EAGINRopyxqyfQy1tGn
IW7o7wlxF2LoK5NSc4PBzjf6YRJLGjfMH6s51rrRaW7+oF4AD5laiZBQDZhwK3Ic
MKZKgUZVpt3e9+pMc691vGgceWPa7XbqZnKMejnAwNfykgCPjDk7PGz9gZGgDDZ5
ocKhzxtGynrUH8sjHaD+ms1iTvCfQwGTBamV0a9MRcTxWaoKS1wqDYnuHEAtdJnQ
dFjp/vxmEtcdUWGyQYeJ5qYZHKD48oAMNwjTY/n5BOka8rSoW2Tv39mNFci7s4tO
x8SX2C/jAbO2MJKGaGGRrUAIgeCc28FEDHSXVhHmSTi56Doc1jQ5cE2aC/m3xu5/
v9TaQyaZFJA4o6UpOIT21OxtKOEwgUt+gz0tesd0NfatKxVHY2KLw7SQ2grZ9uuo
COOeKSEyhKkjxAXAaCQUMv4HKJbV4z35sdBi93L5pzBj8IIOvTWHbwjPfrVJtFZj
LsOLV7Wj6WtF69Ya+OKV1FmW//tnBjnDK4Xxvms3vzyfyAlo2wWU05RZjTnF1vey
ldW+Eha4hG8eJZREg+QDPoqsrdhr0U9GDF4c2/n4HiAwsPgDCc/10j5pkWkeF4/h
4Io0vKRF1YOkAiE5q8SWaHL5fiIiT7D8qcUbaDK+wKl8PHn13u2poyjcYUN34PkI
ws7FhfC/Tok7mFSjf4U/9/ItwnZHUCBFtlPkbR1NwfO07PHWC+nT8gdxzcDwVqDL
LE9Dw12Rx+B41S+k+r9BAHpwxeGrX9olQU4Rud+TVp3p2Nn35rSydkoqEQoldRFC
/4u15ab0Na9Cug5FphE+qLU4/8TtXCd3SnWxbZ9BgDytAAEpuyJnknGpg7CI76Xx
F4XGaHWzB7wQJWY9xdvRpeEqCHk2ynLcN5nV8f4aNjL7/Pi7fe6VM4Jtjjlh1qKW
HsZbB73gZI5zoq9q9+muJoIvguZBWVyVRKEjse4HSkXNJFGcQtX1NiqnOUA0C35T
QhPUInDfJjq+cWbMXwlM0ge9wUrrqX0vJJGKl5hRNCG4G2RY+XFxgrq9mg7mN5gR
wTWoXX5G3+12xV5fjkMCJHa1bEypeEt7qQFKDaPsY2w7pofviQ1R75k4OaYwjMsu
5NCadAsyqi6BQM+uHjmz5VgSLJbXP2lDf93RzuWcF6oiKZxd9+4+YA6uxAoCUjgN
ZfNevUFmAPBA8Gth+0bJ0WFEo9yXMeJ1/8X1sev6q08jPh2MC1QYYCuCscgwrBPV
f10p3Af2PAqlT4w6kiPqHT1cHEChcs59pi+B1nDjqoWzFhXXEvCHooz/kwzKGYpK
UTaEQxd+Cyqe7F0+BRhq6CwewsT821P4R4xRCTcGdBsmWhyO0lSzdaNUY4RDBt1o
6NpYcH/VrXRS39E/80gjAwPaqqW9p+EihuYENOqqthp5DfCPlvIrCfZ9S67EsqRw
FHoEjXvZ526C0xOrl0Yw0ZqFLaIdWAlT5Ni0iMGSYnNaViaKvpMWgds+bep3SPPd
bNeClVOM1L7qHs0nEqLGIiaIsHU7odP9M4IXlPMHgEE9GxcgFC5tGJCwM/lrR+PK
TbHdOg9hu5rG15ORwzsWv4jYdVOBAn+cPM+X/I0bEf9gzMH8Z2FiYFJz3PtWgS9t
vT4jx7uMaDAND5fFI+FpEp3zAssbI72o6MYTGjqfZW+q+ZrAkA5G88G26mqIq02V
wN/4pRJAJ86MRW975ut7f/oWwhOYX+8SiVa9LBdXWoGY8CHGAUhKrCjHLjLifUwj
uii9K6K2hodFjnX2zwMcuqD0YgXs43PWdOrBGW4uILso3OIg6ortW06Rzkvma6PT
iRkTv7g2MWd6pk7QkPzN16t4lRAI6B4cT1QnQOgU4XJonuZ48mQAhDD3MuPm68h6
iWROxGEtmI/J4/ukJLsLewuTftn48S9dfzU3u0lbRaJC9GJoFMz3RN2DxEZumCt8
9VfzaNcV4rN99FqTu56XUPNguBwm1xr7xOjlKydbxiLfjz5gVqiCRB5aSQR7VfSt
nl+uvM3dFk8/3Y/R07DUWOIUf0v51lbnroSah9nVS3nq6iepYue2kCtqYe3jG475
xfdV67PtLywzx5S9yCgFVlRsGmVkLMxyvlkuA3FVzF3Sw1GFv36PqEO+GmRbTGzC
dX2xXWiFhIqSQDuvxgJwFV0tlEaByz065rfnaXeB4IFcyWykOSXLerzXQ5wvMvJ5
MF3KFNbxUQY581e31VdANefPj3TtT/Wjk1PvAawy3gK3w6Ii0J0Xr1UtNl1REjxc
KZHIiOnmPIeiMfu9+nsqERQbwwdLhJyXSSnhEA4+8uin6ZnncZpmMexE+wlI/KkN
Fe4o+8bE2MikKSCCPVt4YqBgpmv33WeN66oHbZe28nCQUTUoS3rbBlhY5IHC5cjZ
Da6ShYzFoOx43SHmGaw8buW4OXQGG2ha7+VuclpyWs81KU+QLQIJAi7HYJvYPrVx
72em4qxvK1s30S+pTweWHwpPurpLF+06o/BK3ny6GNUJC/SN+ncMIz1UvfkFNBgW
R6L0wpZZqX0AA3LoC3w/PLuCpvCzpe0hzesf1ahLGgxFD+1SmAUfo2Di7yoiqbLd
a8Xae0nID614ow6gA2jtWGXER7dXHFehwoPG9VMlrOBDo3g40B0W1ku821TkJ06w
wW3IO0qTeXzID1baCAaa/sMnY20jhMbIT0iiCT8GNZMq+qC24ptMTqxmikM1Lp7/
ixPxCxc5TvKI87/N9lBjdiWhsBn7FnQHpOJ/h89UDo/K18uolvoOsmBm2sFX9QZ1
VNlBhn3p7ir9PQ7XyGTrUwZMP/3ywR2B1wzp4mSkFUHMxVqdif0dxvI9j3iq84z+
7aIZrnizqdlwzZeGHyIGvVejK0Q9fwpFdrEuH6dx+QZ4nmy5LaO5Woa3oguWvTIf
MQt3uoKYqSZwssJlQypySY4ISd2Uj24XukOOTdvPeTbg42Tls8EUCAwSAtuSlgg5
iLjRoB+taQl0OiGwyTsumtG3d0igcDPbZH1LBfhyx8fhCCAQm6p8aKfkVd8aUSwh
zyYLPNggVWYEO6zUTWQN/4uAv+X6+xmQyxwYfWGlagNtVTSHF+nFx/D1uktDYk3/
DPhJo7Xhjf2FT6+rZR36kxT6jeSXHkWF8n3YlqsMde/YX+597cjmtmG3Xzz01ydS
CbKAuAoyVi+FFy3ktSll5ECKVTcd2BYT7rSALndpjHcKfNUS3q1k2VKFYj4y90aH
zqc+sv0HKaQz+gKgEYkVSRFrB16wzbGFA6vf798d720TB06G2xThasb8zSzhfnWT
Rg7YqrsyIXTVws6YvvTbLViFBJpr6OWL0BvRg8UmyhJE4rVhwsi+Z7xKPdEmWxIT
lbm+lvC6c6SU0O7tUgRcxEUT2cggqDvs6NaYKHvNnwDdhAi41D4AK8jxEP5KmFHe
jhijQdUPxwjFp59dUXsPBL0hd3TIQPH+DFIlreWVzeaXliEr7XIuGKORk14mDsi+
4cYJ1VUv+nvJslYO6PTdx9+rNHBfyFfmjmkfewzdo+A6wyPVMhQy/Rby6iGKuMji
oMP07eFG4Ao3PIYCO+fx5FHMEAT8eFRTE7Y/eZsQj9NmgvZpHS/peHp3PoDE2vba
ziMJo7kGGPxDHrV2OVs1aMRZruKMibp95r6tOH6cRqiXnQiJcpU8TFGYmijTSwPi
qhPr7vDkkfx0C102hUMNTyh2TD3K2cnxCk6S4FkoHrQdZi2MkzAetV+S9Zka+uPY
Sh5QD+BkNGYVM5i8jCE2Fsohf55Y3wU8O0B7gC1vSz7olOI2Ei4cIankKz6Nhkqz
dLeWGacvTRdNDYeqe4Vy8peHdgngUMxo7jDm+ey4A4zs5UmDa0Ck680BCJd3bzo5
DYb381fkJ9TDvCRkhWnjHLIYPMChQpyqJtw4OZnOoExSnb+9i3DEnWiN+qb9WLr6
OhsdkuzZ29mUFu/ZVbZW0t25cIoAPB9+Y6uIUJy6VcbrdOFwUzL9wKCrPPGiXgg4
PPR0fUOIi8MSY61yUZVJmYS9Ah6+8ko1XYMfUFH+4v1oLy5DXALK0fxhxJMpkboP
JzbGZ5fa2EvWZbKkL3/UPpk/2UNTSw46MPKJFxgIETEkNmOuH1t0WoZtV6a/BH3O
oVfqszdcv4lCGtzLiwNC7+bAWaMBctb+fMUlufSwPi5KKc+mngNysk9vchvOEoQW
zUDtr1xU0/mae10WsfmUfSpUlfO9YAXN0LlDaqnxWShlKYGzJVWNfWbJ5ssewKZY
tcwLf1I3nHxazEsQ59QPLtKC+rJgvEeQXZIxl+obpHgSV5cTuGee8mzn1Edk7/fr
jF16Ct0CwoacLJcXgOjoB9vxhHHvEkJ/pYVdQT06uEZYjyjEcJ/NDmtbyi59R//I
86sBHtaTNBbua93+xyV3bAYIk69grujz0rVC3FicXCnKIKgoXNORMpm94stIdizn
eiGTK6lh6CwsAua6AZdgukB7b+VNic/P1YIyqyJlV2kQUt8Au8MZ0sdOz4G+hHRo
DAGBNIwx9dm1Vb43rrHJCy1ZW7IHoLtOqfa1D06IMm5E0b80uau8XN8ahmD5xUkO
tqeDt9UPKOGrFH8AZxN/0CpYHmKbk2JTnXt7IwmxrrIQTDUmgARzs6OnRPi4mhwf
PMtGmXV2qY8GAfLPOJ2fQzn3uWjyDIAZeXCc2xQrvguOmqxeAbiMyqq22z2vMqZn
NF6drZAU85PwueYcQWoMpeKW8nWXtS7WOv/HQwpPsWlhjZjqCzoS3+0l+8wZAn4u
8r+wYIlhrCJZJ/x1Z+3v/KZf0FVkrONn1z735tTYnjRvypj76YiAco982XZGS7PE
SRd5X5ag89LApAKY7Bgy56GnzyU5B/P9q+kkCDDiGc/ajMlW+o42xq+5ZGiQj9X0
BtbF03sn3HDuZItSwe8SHfvmE0UC95+fvaB2jG5Y5K+MFRrxCWRWrkBHmyCZGamG
ouQsQhB1eLdZyZe1IM1lI/w/w8n6iJtckj3JTbT4c9wW7lbE1G/XipzgwtTitdpR
aLG00YufiyrEsvASyo3dIhSPaaJGJ5DJaOuiUwSCABE+J4HrdLqXhS9giyla+2VR
E/XbrnmDa5iUZbWqccqCiwgaUMC7MKs2KOp2xYlxXHHJZlu0bVy7asjv4/aivTtL
R0pjYbnN9hxIM4UUCjkkkyoCRKRsozRQPyktBsuQUjUHvfiSSCrQNOMK+XUL33e7
ZGnFaFhtZlTEqOlQuJbWGd5OZ5HpaexUiNbrdGe6BB5OtT6ZwNVnPaoz5fCfhZJ7
FfY0ApM4BTFDLWmNBMo1uDsBuc32uXbtt/V+kIWFUOTkuPWpbV2T1hnfCnKHeSMa
Q4YkCu59rkmC6LQ/i/hFbWbAvqf6lmpx12+IhrZ0SqYtVCdCsxMvCWXrO2ptd8k9
ydvLRGllhq+aJpozQd2dl+UaCRr1wMVL8JbLiHFTc+3SaPzDgqnaugBsl4/rn3gn
NpCxOA94vTTZD4fvbGYy+z+6v45KwumIYUO3yrySxOUMl9PHXlWA+VKs4lbifoVj
ci+NcvYN1u9qNycu/3rNDof2yunrgrmi80Y144TGzX7L4/kHcgd1B6OXKu1YgcdU
AmIyax++U21etD2RGxmRT8E3VfQaXfiCMbC1uFlbAAG4idi1YsURVrCA+vYT3RDI
wspVjOZVXcr2LlZKKiSNLYxE8P4X4fntdHPZwXmrzPdLVDAWZ+AKYNnoJMG7JZi1
z26rcEHzi5QgJ4U5uzoLKvr2EsW0lerEQuQSvLlqtiMF6IrLCCyHoVteqhbj98ef
WifcR3Vwvz3V6hwRcbZnhMVBC8xYIKSkyfNn+Cb8YYWtok/ZbLuHD5a4TUD6PEV0
ZZgV2DzH52k7bZHuHVlQMC0v0BZM9vgGnud7PcgPgfaejiRjYG4dc0HI6qMx9xm9
sgVXhqFDPsyCPe9TTqGP4Ts/UGveLNfxZSBAa9l3sZAWfesj+G5Uc/ZsEGle+xSn
kk4xBo7C4pFPXIhomESnKnJrgaGWs8r/kXzBdW0XddBRhXRaI/Ca71N7qC4RdJuD
HyrX2tbKshQVDNSBOcpHlCzA58ZQMMsYBFIUJKsLLAPdx2OoENEDdnN3tnSacSuY
oQRnq8qoLjDDzZKWLIBLkTsCSiWvEJMS2fVI9CaWWZX+vdkyAaJ93NJZl3Tj4GXI
UEB1xd0FJRy4j8DlXj/CPgdEOdj4OYM+cFT7WL0ZIWqusRrCjxh2OOhq5RLeL/VM
nMj92IATqIJmAOHVogC7l6tNFxe5yw4ODkCudhCNH/8gzIWft7DM4gbUv3XAJi3R
IxGOxVKYX337IhYpCgk8HFsS4C9kWMHjiaeL6uxq3Nlp10SgAXGv/MJ70E+LZnkl
1mAOueaBpaBwbod9ivXqkUp7y8NyNcNmVYZ812l4i45EU8oE10ZCg0nyKOCyRp2g
LU4NFIS/v7RZCxzousAZMC2rjqr02DHUinKeh9bxu4JwXeSym6vutMF2JCOvcoAV
mr/M3dUzqaB+L5BpW5REWp4K+sNE2wCL5Jq5vP2I2yLHGwoKXsT93BGc2M20Fdia
9TrRRspQ8F1gBGLXW/nyCCWPH0A9LlYv42+f1AEhg7z0KxdfH11sCkEET0owrXaY
CRVe2ONFHTNxEVHDQTaUFbmKcT6inDpnsbu8P89oTkt9CYuQ6Qr82cX/JaQya5pC
xCX82dyiGmw2CIcC+uYBGQtMhkiTg3FQ7v/W8IW5RQvdpS22dpOxOsrGtvAVXGFG
qayqaj8X4yzbiatBPmNZ+6X+uN6zXdD3gFlr1e434GXgqhQ/RUeDEdhzuy9G2XCN
e6vWuytXB+XHvTvGysOn8CxEU8l4OIJHgin0ESGNJegnHnH8sEQUiPz22RUlED3s
xrzace3qLMCu4HNuMl1ofx9lFtxGAJazUCr8OIfC7R+bDAHPWPjHGpokzOscu9aD
8EIiiAcmSsyh7N1b7xl6e3QgSKa3tvw00plQ6CySrQ3aUIofqEbQItTwVrifv58x
a8kSiQ0+TULT0eqMgfnkbi6ZvyIQC4BPOY6xduDdN/XKP25fZ6/twkB6fsKu8Bvh
9wVCBVOl4mMQyduUfEQh4x7O5SWgKTJCpX1EOkYafeXtvqroo0AEeTO9XoPt2KnE
IS3Yo2Z1wMxymNTguVp7TyA0n4P2V8dRq11PDl7pcFark1DYDJC23KvFD4CGJud5
4I0ZHfYi91zMvms902kb3r8Q08G0uoZlw2t81Br+fUIoTfw15Gw8a4PS1wg/PYIp
PYlxMsnbCkDQFuN9Ul9qWFeoz5Iems3w1BDjQQDkNO7UOcPb+8uGonhenXR94Na6
uKIom0hFi1Fl4tP0uB8ZxCD/UNHdbkPYkiXsLJrw5wlsd2SOQY+92Wn8R9cXZrsK
MAWl9xgzPyh54pyCf9nB2Nhea6y0FTtKhSetgQYb2u1tVocRN+5pRzXI4A7auXqq
13sA/E9VTpT3eUg1eKlM4fq/kD2WyzWliKzGH5GOty0F04p3L2ZVXFBrJIkCBwnN
8XJN+lBvuDpY0mlIHr7W90g2BKpUafKTKbp2swyYTEWHFMZ+IY+uv/8SwPY+6hiJ
8gH0Tio1cxheC4fY8hfPqGHHEosrpQnYNq5ai+MkQwRGeZo39NwPvIb3ZT6tcz7E
2jX1eNLr6qIMOW+nFH39qUCpvob/ExDNFqO9lycr1vCtxUIehEULRBxv7wDRge+k
zuv/xjPN6++pM6qozYYLW0VCdrnK9lZRF4+SCb9/X+cRypYLrLGxOiTk23K7GHUB
g3fBISOpUUVSjuT5RIcCg11hsr4idj4crf9Tp+APGS12/ITAqKxpdLdFx4CGJxm+
TWd7xN+7ebY8JzaTxBfEzLzXWuvv8RH/XfFl+82pSDEMyua3K5w/aV2h6QXZmg2E
6xiWfphWBGrgmYMkd9EcV+fXf/poTQWEf06Pwj27wCAJosImkLR6PklNZkZaqNF3
YTbGBDUMLK1eHWfQY8rEuwhDZWm38/ltjC01CJPk+IdIy+ZmwEnCUqvChyvM9464
spVzjqNqfCKyBZPKeRKsmGBQdo6VRXKkyCl+v2cC6+CQ8CfBYI5ByV6032mzGsZP
aiWjJERxsy/hM/BRVgPKra5m3cLygMnnLsyFYWDqvKuFit52ioR01117WjOB5PAz
LMYy/JYpDCsDXE+9CytBkIHW+Egq9TgpXej4OIPhG3Q/nVEtYnKgTIQLXvfo0Agg
ZtlopEPEg3JPznm0OA/ap557aZ2uMTbffX7mWIw45YE9LQ6A/2xP0Ic5BZEahykM
ulab7Uf0uEGSrJo5P5cTNWFbzY+V/oI+Gjjt0ISvzahZjadVxuqtuPBqkuFQ9fD9
EpzDjcSaNhRxB9Q8TeXhcTHV/guELCPvuSzozB3v4DO9Ql4nz+qTP4jlAI5bCKbS
dlpAvvjvndvTWmi7rJL37nAQZOdA/m14jCwRn+FOkFD1Mu48u3eBxbRLBJCg04aM
yLzZG+TRyDm0gpuKAY3sU7diyyXzyZ7wHa79KkbPCNM7InlNM7FZw/C/N7tPbe0R
hDfgw4sZ2Js0slyGAYHUO0m5ELBcM1Y7fDEHUTdIMRXCbQBNnsf5I7P+l9cF9k7Y
kVfjPPr3SGD+K3GbQG0iY9Vx/JxZ1P8dNkuAMgCg8NwtntRGygWRvA/l7+4+I/ut
VCW+XHxANdwTZJOC0aVcrgKuEpIdgz5AEi0Eg79I3j2UsdaEl9vJhXa1kLUCMK2D
4NaLXXLax8cVkw1qp42O6iR0CZapA5tuH6OgmgrWE9BD25F8ZZZcFWYE1AvmjTWo
hfBelzagXOlcg4kok6ISqMY2nt5pvntoBy16ELYolTgKZpThvVQstBGyszlFDerZ
RMOkZfwys3rPAsnTTqW19LCqBJUO6QZsLjmX37tqq9Hak/xw7NAav8di5rYAzMET
DBSkG2I7NFtn2IVXQJYBrxT8P40U0jLp0D0jpvGV9bXEkuM6kS8C7Lp/kTHU7yUq
c9Ry1cFe8VsMXnlDkVLsRomfwYTVwZ6Q2A9IWpJIHf7Dpq74Hkw4DRQYrchFEhQY
UKAJG2rEkPOR2aECblBdLCPeccDSRbS15+mxcBVgb5huuS2wdkeYFovrAm6WDpZr
x4R+kWcpxD6SDSbYpwe40JntG46BCy8NaSZiy5HeSofRHpEF4YZ/ldKMgDMjag5e
BP4oA94guRl1jMEdfxWi+9/j1IBM4zPeIZKN+Fa1sCqMiAw4l+jVpJbLbaevhgLM
xzeQE9DnpXNtVVyILPyJaRBcWkRwPePTLS3JHk3DO/tIfI4ZRcK7pOr3qv2qIj+X
vOjp8mFKdLwzeHCSU18zKNkUrlGOHkV523zHtq/QLHqWfkpy3Z26b6ZdB3YGbbZ+
aw8NafF9FIAipPQ3lAPTAg3g67H0QjnFP0YqqSh0HELPrrmMiFr4uVAwifD4UHQf
K579FgK0TVU8Maw8C/dcQmzBvRevjQgpWKaquvK87g3KsMkR74e7wR08IXsM+fj7
Vc7g07iadeAuWkz84nqt36yZAZ596020dC07mCOsjWuo+5c/Bvx9izGUbID4e7Il
C0ElmREUIT0vUqSR996oNxdocZQkp2mMFzlbxEX616G7E37mv3IOBsy43ZG1BaMp
G934QJyWkUv+0zv264MGPquF2nW9rPLv6mKV/DfYwUu54pBWIX65kcFoJc0vBwrX
wGO9vpLfdt4RZ6swXIqTBs8LUpV7FlJ5L7EaWDdGyJq/UIIee1VTFyayr1qBLBlq
V5xb99NfFjVuhqp2zygfuf8/EfNxQFqBirEiONJ/+DB4f8TOh5tH8iXB2fevxKP6
nhNRvs8vHOvB2jj7bOvtfSDie4YAWhxOuXgEBaW4oHRiG2DXoq42E2Tpdkmq+a/X
JFkSso816xSkY2oYrCSdxPSl8bo/qGx3P3GPraUY5lD9eFZHn8IA6NofHfR6e0yB
GBiUonqOq0Fur3XNJsIxRNZRs/Tsqm+ufz5X1lIVfw+7h4HfLiqBM9wavEMN4qpX
O+NbKT59TNhLOtB/eGfRoo2hGF7Vugm91eTfOGdZGAXqhJMp2A/1da7goxwSbK7Z
jfMW4nK92vlqRQxJ3mAaK4eGJUCw7Meu+X0DODaLZbszR5UFySqHzhHu35BGgkyO
Qk9Wn52qguXtLi/7xu+iLpTugJAJMWShN87MbyWAwKi0j6Xdy2VCLSnyLxGXBB+Q
AO+9R1xu+NfGMcPGmZbBEamvilSG1QY1AvkTffVpxTM=
`protect end_protected