`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36704 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
EQKoDAcJ/8QYHXxJAKTmMKPNqpPYCFukXqT6Tz2OrpDVkHzXA99BhKDXNQsV6kzJ
SQ5OLaUuC+WN3nu+7TK4RUd9xEsIcDQEYShkrfY9bZJiwFRZUPcOqyqdzLtPoZA4
zV/QO5j18p0ELkfr4bsIhXTPsXnDyitALXS+cfe+wGJDQrqsdpQNqnQZAPzsSWQb
l+xd2A1+dazHkaI0dzKYH7nudKSIfipG16nxSKj1SjQYRcieYTzvgLZe2nhiH/p8
7l6eNKnFyJpBRQCf223ZdqavEaLxhMcO6gMMWrKaN7ewdX1i+j5xdE4G/VcBVI1F
E+aYuoK8l7kLNKy+mSLB7jQCYO4zNAm8SrtQpdMn7pZ5sQOhb1AfK2JiP21KHKc7
07ZmCvUEcPhMpMuLVA2NW8AISyoagp0VIl3iJfXtkzKS5ejXGEBnckESmBsN5ZBn
fOkdC44kLvkbAXTfF0/zyvB+Gsgs2QY5IxeWliwrNjU5i5syCCEqR+w9GJCPL7zS
h/Zf4w6SR2oKI3b+1Dd0nolUiuFsxF1z6hC3V3TrcCqDjgY1GchBDsbicUeHuKcw
625f3gsnuCQ9w8etZ9lThiiNSNkBPrnvrkN9CWs8Jyg2FKNXJ/JZedmeV0bji5Cq
GevbNF6VmzQ4GMYVlnzkwsmHDfBfLAJMf+jn6KztmhSTmKE8cmZn3cHZYBnpiqO/
4Z+A3E4LC+mG3MVQGcgK4ReTAOrrb6Oikag51uzH6NFm6IvgZEto8W96zbJpwd/f
v8HXIDV1NTmXKRcJLrm2TAHkmM2YFuJLMFz6HKzt02Coo1HLiRGM6FSo953Bl/eG
J+rZ20yLF1OHKw3hkUU8new4hZ+3BvYPYpZbSnL0xW+YNydFACordowH/DAjkOIq
9cdEe6pREXKt0r4Cof9Cg+NqGHmyXFu3x3fzGrVRWhjLFU5TWyIx8sTbV11QXZPV
Wt5c4BPHQZzGHJ9RiH8/iTCs01d9CA2B7KEZIt//5O1T1YrjglaWhaVKYROqkdmI
6VP/5QACD+BMrAHIfcsrnFKJxZvrr7D0T1VVPy+12gqewym/PjWt4weZ7RKI+3RX
v4IYUGd/ERkvwmIZJB9WwHnE4DwmP0rZ85Y2bGfVtFWJpk02IVOHUmHNn3ohOJ1f
UuZSg5DwSxwVMRrN7B8zf2QVHHz2MaFV0vzFs79oaMQ7LwRvXfUpO09aiyrxEppR
Iu0MtLKgKx3bkqDd/o9ZYx8jivBt9gqZ/aPN9sOrWc69022IKrgg/lEek59u86EO
9vyoAy12m8FtvcNTVtInFGjCmE0jTsTWxSN1/77fDHqVe7rqD6htFWM8dTnQAK4O
j2QJXkOMb1fM1fjKFHEzUwu1sEycGKyM0C8mRpdQgvojcdolPESFMOLP7DZM7Utu
hQb2F8pRt/ERONXl7b5DTbXdC9fQHtLGtg+74q2WG55u6XhTYttBG9aOjnaK4ENe
iPf9j+ODLUS9gZNI9aDtQuonjf/GjBtn1jhELefv+A/0heBArr0TXGF+1JfCdh6b
OBbCf0/LwELVVHuivoz0RYFGGPRTUhDrQkaWTidJM/vP0sTSqEBxD4Myd9rcAnKs
0Fs/gLFYRcC37L+uJvDkK0yBWWNJTK5MesSm1cG42OrTNdm9TtSq09tasxbt2wJQ
ykS24gDaDP/5ZKf0PUagGPHJ28ygtvjV0V6M6MpdhX9gw3p+5JauzlnawmhfrYWD
JTjHDGbAzGW/q/iNgH1lFnObeUxjktVSuAJFhZUZ/sjPRUBmzoM5TyVCKSLcbGiL
43Ir7eLBy4ZL3VVy9nbXQquJzQJGA4f/UjQpwt/Dk8vhOQoQUXMihnV2iL3B0Gbi
t86xUyHcQQyxDsTpZSnqOiWeJ/G/JucEn+dYzA6TJ2nLvuc2M10fd5RwTybdJ10b
IVuuPqxnRCH1J1z+pylt7Sh8ayCBXxuvCjSqIz8QAlw6RxfOL7liWOZesdPdmKDU
D6Rj4NCB1T50IipnwUNwSLvFb0tFycKYDLR7XgpJ7AC5AKgi3eQEHV1sRtol6OJf
y9buPyVHhxkcxUklLW79rhcGG6X7woO25+iT9zVi2hdCHUgPuerehCqcWs6gQn60
gNCSL+BWCpiKOSf7xeC/s8cnzeixBRISXNgK7ilmhyDTZVOkOKoQSRe+bvTHKe84
vU/03XkFyIMQHsGHMx/VMpriBUR2mSkXOCo5J5BysxnJuvLj4JSfCfyoPk0Z7BCh
2iKimNZlLU8dfC0HN6Y15/5OZNXuqvEVul+Ipt+NWBeDv8JYM0hN9Jk3Phf5Vsva
OZQbxkYxwBNRI7a8gtlcWhMNQ2njFfwx96pA7HI5Gfn005U5J5SXF94iUGqqZuX6
IuEd+lQ5NA8HLdfDJRQ5aBYJpqMicSgeiamhN79IfpjcDTTSK+9+cdUAxvKOU7/n
OGNlmGEh2jlw5zZ9yjWm4J0rxsEQxuxYePUgRDXfRfRgzxP6CHwsejgEoYCEO+fC
/sLcLHCc0vWuoWL4k5yfnzPGOas6rGvvUA2smGKLKSCMSOLFYL0zycncdAyGt7dp
QkwWqGU8+B0LplZSNXxkH5EF3Lc25qNi4mpWfMs6DTLBra2uK2/Wv83bxNUHatbH
Sj1+g48EnYvxLS/l6vhKokCp6NclWrOVgEcORUxF2MIwGT7fe2jYKlbZSLnPG7qW
vlDuMouwYvyXA9n2sHJWSWCknPwQVvFYqNTr/f24QR5uhP91NWn7lS0tfBcPJDxb
Tal76J9+s2uzIhzd51VVCMwS4KFh3/xQwp590hAmE7z6Xdd/AFNhO6gzOKuSnBnj
hHtDMa97ijWBqnd13pDbIWs7NXnehz4tDYWaKW+cdsIElfgZ8P6BvQL/qiquXxHH
mjmXlW/MzcKM6n8b1NU7BsFOCIogYtcqCmCB9Q6gNu+UUFsE1pUAlPsV3yNOIc/5
9qCkwNhtXz5j3aP2RbkQWjh4lUxHMrsZ4NT/rJjiQKXcx1SVr0ya1lvcQcfqvcMN
WqHhvUVKvrmIFXydOXFlnw+iNOj0uiWeHUvAXVq9Daia7myp4aFDH1sdvFffuLG8
oIaBMjs4SDizeXwRv9TdRkG6hKYwoACLjUJ9gIc9ngjyXYG2JJXp7w6dDXlow5+N
3MhtSnie6KAiuO6NVTUC1ESOkbM+kTpriF0cQHSxpiTu67GwLklXfAjnDPpIgHrr
jn+ns6wxlPgae8LmnxU0FcFXbQxcVpegiY3kO0PCmXenrhP/nsG49cc9pXDO0Rbj
IDDp/Brb/1oFn5IZnpjvfTj6Sp02HTWxY8xtE6ol7AcEQv4zU4VujWHzj9J9lfP6
Wz0xF20qQ2Rlznj/Fhw5hphgNBGwa7Q+01FhTfh3Oq5Z4Am9axE2Fd0bo0pl58lh
4gq9Lm+GdZChwBZfoR4Ncer3nZV5RF4jvxHaKmgbHQkZUXgAfRsS1bZb5ZhFSDMd
oA+ZNF/SFpzUcJY4g8pL0XGVUbOncQEvGtK6r9lOTDkZDSO7p8NY0GhhHvEQkk0K
4JNXe3gXyxCJxjEglPPo7aoYfprov9ybAAsk0foL6EiY86prZTfvrFbmEASk69vr
SoQP606P88vVCUtStnCRQW+Ze1RiJDQpYKS27euu7cf6bPnHZ9ANZ/+kSq249EVc
2fsNSTPQ8xiLjF8OVKFa4J5c0afgtKM6VxpWYfSfSSWUIBZngCXDOvZllxpJDlSn
SDiF9zmcKbtHn/K17lBORrpSmN24UR8914tjqvN8KfexGgSX+4RlzceOJ0KZ3d6p
SXgaDhlembnIhtwPy3/3KO3eXYjGNT6N7kHZOnhd47bKyObsRFRVmtRt1MPzEiNa
X8hCLFgt4/YlS8ycBUC+hqTdyHMclbyxqd+ucSb1bitIZCeXqVRHK+tvj+04JhpO
VzTuIOOd0F1lXYDKeTl6tQ3UUAmaG6IK5jF5Y4R0RvBDYlWqV+qbSzBjiWk41rs3
62+tMCzPwau4ZiE3CrcRw4o0QU164+m9J0Ci35eBt5lWM+fukwrDQdGwBpltKkTC
AeyIIO3B4wl6U9LjRsWX9CsWL9lP3s4BnLZX6qxv/WbPaLCyp1uPG8kh6PjPuP/4
wzw3Fv3gYVbe2i1qxUXbSxX2N0qK7aKNacdfhoIPWyVnrIPm2vpC6Lpm+hL95eQ5
p20QG4aMtJwg/KLrPoDHsiWHzEgCrY+Ug+D29uj5iGk2qf8oDDd10Dc7UCMMyRsM
5Bv3kdTpYZ190yTAf95sF8ZeRMj5QIEnrQ0TjyqL7Ctb9A5+HQ6wsIxYBtBsyfV+
RI37w0qhNmyk4P4vfu1ZE42SD56Yl2+dG4o+TCJUV2PSU/yUe1Frp+EkQ48aAblz
2xiDnMSutNiah6kIbJE7X3zExN9ACRnYR4w5cljPLSVnGwKcvA/1WwlbQH+Xv92b
sJu75T7IlOPWfe8D0hMoI6MshXXqngdZLPHpAEJSIX7XppNo10CwJGpPFSukmD14
QbM53fwP8pLIRt+fKR9a4LdvOPRufaazkamVZTfTHFct5fzye/j7VgNgTmUonMsp
jrECjtkZiPX6PmLi74h5hP+mQ7uBqgZenMWlnwvpEOiLeTFFOCgkkj1qnWuiyR8u
fbmi+0im965EHvUX/O44Kf6gTqq2yNZM9mvNr1/IjVXzjaX/ZJnivJpRIiMcdmCm
oG2RoUE6ItIJNsO6E6ffv2oUZpMU20ZFfw6mNv1ty2UovCHvOu7HLfRVVJLsgNSV
0NKs15H76AW+MOOljJymmE+THuqEkjeuQj0wR8wCAZl3tTBMHcKP8o1Njj6NsFTt
MdsvY+cG120newQmQzvKmGhfSPcHN8j8xZdfIz3Uf8BhVFQghv4NtlvwhKyWKTVv
7xKgLrkxDJgzWEOemzJIaLU+ZrHSQ+YqrY/RnKSrJXsdmI8WZfWuw3tn1MBUlhJ6
7Gj7DKAPz+ccD0ToiHNEACRuUcSQpJPpc2j3Wh//rWJpX0VJk80JwG04PbRImNQe
kIyAyMa61hBm/uyfwF1jolresvhfFnE7pgG1cW0RlPBi4MmvRFPtSodVIO9CMsL5
UeNY9z155yE7oFodl7aiWfsSzodsHRxwlHeK+9RXSwePEswDTrULMSZGeTiQQkGB
I+ePJHh7DcNWTB4NE00iUoIExiyRyJQcWMeAgkI1LeZXXUldLzlinYsIBIm/vbSp
xEM2zBHtxKZxfUIGSMZeeWtlRin+EC85eYXJon4iUZ1xjb4p35gv6A4TBlTI4nRm
988x5Cn6eu68+f9Og/6QI11dRg0QjJ4MPPYvRKxWN3wybqlSirFWFBoOqc9YGvMc
4s+aGuC4ETTbJesHEVpRBDywAly5dKW+lFTtgQYMCRYO+oI43ayz44LvOL91rsKN
K24hdll2ZxZ3P9DSYSlyWjlCUcbXHRkitSdmgDlRmANephgu8go7/uVgF2quzB+H
xtg1VrGvoKR4Uc9Xe3N3GQVKTmObs95dtV6uC3eBuV59RFVW4nZOfjNN7UZN2JWd
B7paSpKd5s7jBwMP2Ht1cQU5R9pv5eBuPpUuDvbj2Iif4VgCx+zGKDu7lIKYfFWx
2iIPoaqM1IYDk+qWzfe8Y3ysBnmbNiKXuR/DA5rbe9qo8m0mfrIGQCjEVmbkrgLI
z6bCRQtwmUa8GxoH0mnkSitw+x0lvwklyaOe/uZLEq7llO+nUmPa20Mu5T5TTaWz
X9YtEer1ELolmYbwQbkrxzGVEVAmuC3ObHEcSMsyDtnNXBL0Ky3loHifYOs2Kp+H
EqmsSPikW6+vLN/YeyjnYT47QVtwb9ItPJXeDGtX78wReaPMCSe31Gw6F2yEKzJ+
IUzrYb4lQLPx2R9RSK3uq0K1YBYJveIx3Q+qmppUoUYKiPt9IjnTtF5vOH/FYNR0
WhbGc80P7/8aB7ZFrBwop1HUHfbusux41vhJlCtnTlvhoXH3t+7FckhRp2WuXRDS
zniTKdeEi1D9kbbLC+cU0Q/N0a3jbXFZTx63V3Gg4Wnt5uBNZExwItKKLoY+TSte
syWnu5Xv1dddOHXg2Owf9WfOTkCvhpTw9pr/YrlfYhKMxBLND6LgMc5/g2n0Y0FV
gHLb9gKODOA9XNpcQfhNg9QJBTWyDwJ/CruWGW9YETvm6AeKJp2sWtCq1AxN18MG
csTLNfrrMXLAIyCqaucTXcOPPaToW/d93G6PggQrb/LQuxoKOU+1fb/42bkExn+U
fouN25f3HlArV/JjpCAK+eKNqkKRNNJ6ZKLw3LvwVsA++DrhLr5sxoQmVmzDfXom
l7/c9wusclnpanqVtk1uebtV0SSkkja1TwO835oz2ORpUUlf55hQm19jBA3VMP1B
DIGiwfuBj0oqG1XfjJx/tp68wres/uwdLMhk8zZTPqLPc+hR3cAqICzvuFVfbe7A
+ShGwouhpWjTTOvYYXtvTmUZvgj8+5Nn6zVI1LLNJf2Y0Ylqyk50KQhCK2ZakHJF
iestQIXFcAHp9h235gln2zd2Phw2IiQFLKwuT85DZDizvoRqVM0L3xs+zGsC71VE
RQ/Sr4UmTWmGnVNUaHqWAaFVLRFKm9gvzK974Zk06O58h54JP88j3jdSs5yJZaT1
aJlCt3yVLqbJ5LXsjQXaAk8O6voW8qDvm1y+tB3QekZpW8WZXPMewTkhEteC3eeG
Cay0rOHvAtrGP0VbGEDMfiTie+ctnVlNBWUbuecKfOcFP6KgWknBYUfLSv8rbkbk
QnmSDl+Nm6WvN3nSqoNy+DZGMWMuw4xfRoP2k1z+V3flrRy1VFEcpDKPFGgORe4c
QqSCTPpnC1nHnv+eQiAUow/n/Qd9NEiK8zO/hINVPbjcEuFWMcarSIQcc5vgfcMP
tSpONEbM04tEE0vlfX/7uKBqv9yV4ZE1kP+ZXM3ifRx155G4jW2FqbCLaYAblEBm
s7faJ0hLn7dHx7rXHlPUdRFhRsMM4x7Q7CClxD72UlXKuHQQaUlvplsVKaBk4of+
ocrm1D68tqv8+4Tcbv+yY+x9hj9FiRhCTn/E8qm/8yJJIUjf8vL6sCkv2Sph8JTb
egO49jKfSpAQyWelWnIodgescfr0k4XoVLLD3GkYv2pLTfARg2kfwobFDZZeX+QD
m3i21Bsy1X6crtVaaVQypN8vAWrfRZJZReIL4ZC3ZiKfli3U1InkkY+x84nMmY55
EoMCQtmBkrfLmj3iQDVfjHX6OF+moKmJ+a/6IWJ1oPQVE8lHoI9jf/iTgwwf6Z9p
MLQktv0l9Tmgc1uXpssOqfYruk/wv1Vk7ciCTnz20CZw+wkwiyY6Zr7NpepqM3EI
sZ080MhleIdS/kzFdE74g4DwNLmXjbhAXe83z5qCMJS1uq9Tm95nHQd5YXxlwJON
PjAE9NOkAk6RGvuIO3/jxZYl/eef2dfuAcArjogybRfNQIpOaaRVFoPXdJitu8eL
eFvFgrayJosGp9pHWbbP4vjRbRAWj9JuZ/fQ9PBHvc32F5b817of1n3UAspIsz7l
/Po+tp/hRSajvC+PORlZ07YOXB8uXn8h2z6s2GgzAtzBmMSC4bMpK2KiUHx0Kq1y
rIPIkBqbHa/gPaGrM7Hask+YtKJe5nxmgsV1S7/8I8tfmuJqAaGvhhcAP53rNlOK
a7HI9la+HfZBMJOqmf/uAbXI7nkYDwIoL6SSdiQfueJoQBZFWHacabRQlxF4l/hU
sVaL6MNa0m3b9G7ewdWe9AEBWHlbaecXi1qDHIVWnVX9OCQ6r9xft1KkiB5rUnJa
xCaaCOgoeJBB5bHLgEw/ypyLUsApuCVY5kzEHEkFSe5t0P5ZOIpDwDoOlYQQ6ToQ
vQAMTXbwuEG8/0w6DbxdLnCnQoQlRtz4Vl/hVkEKbAgCLZM39HDrpjcQ6Lyy1Spa
HuclPrzDVd7dE0qAJTpipMAUwxP3I89ttrrLULpkBx3O5FX0B3LjkeBQIpZcQwXO
aLEFsa0FpBTnGUAGw3TaW9C+XTwPHE5X8isxyHolt0PG1jfGtXu81hB16yNtUtM8
njUjjgpeWvJH8JjLC0TCnqpCKZ0VmFVHwN/GSwqccQIKoh2g5zuo6rx6Id0sxbys
c9e/jKCes52pxiHxrwyC0udfN+jDo6dWeyN+CdVL0p6KUKnMWtl4WUEZ54irIoX9
3wVYX2qSHkXuZM04WwOU5sgrsEW/Q5XfIYPPGGKmZQ9xmHhKgCh4QR1OXU+ft2xV
usqXiG884Xg91zCHyErnZD8O/XzPRGVfoWKFHIWhSSK4xbJHh44Qi/wUNaghJReC
2YJSTBeJEM+vEzC9CFwA03u7vD20uLpIyToK77e+08HXKOfR06MkFz2QJD+CCnDz
OULvGDs9xTd4ftPbeXVd5J2ULuWjuNolqzau5pmxh4M6Pv06CucpdtUJ3qw957h2
MULSSYThTEkmG4FjPuSyhzQqMBZa84nX8X1+4gwlzAIMb4StOnXL6aMIZ2JraOAy
IL68xeU9iZ+OfH0j8VQSRJ5zVbbHZmlkwddvcJS0WXQ3WI4COfDw2a+BKboPYc3v
MsBr8Zg+r49blOsNHnbv4Y05MRN8uk0YgnWuDncc+ozYMMEeGiM0HXZJdBIIvMQ7
SBpjy6hmmcW8OjW46KWJeaDBEnbeqLPdZi4UYS4W08TvaHlvsGLazFAP/bDRo37j
IKnSSfnCOQffXQmbkOpLC+vd8qRfzmhI2dIIfZhShuZ/b+Q0egDnPlDJqoxtPtaq
9kKO68xMIcGBI5fZQI+7ojC+pQ2N1CwDW5Z9YK2pHVWW0OPsHjvQ3Q/VG5ofiF0e
sUFECcWL3D+1C9Ad/VgwycVZADe/wJbhlC9x0ano3Yq6wiHvfh5nLEEoVd6UmY1s
dfu+ltQHRahzy1/yU3oO6dhXaSv6MnDwRguPqZi7arb+TgMEINxa3utHxKVIXUkx
ik3EAaylr8oX+S0XrCERPy//sv2+LSPA7v0f6maLGcTsjoQ3UPIRM6BiFijIkIIL
k+0I88eq+8gOThUfDXazGl/5BJ+3U47hz3kptg91c+HRuaX5lB9Yz/VbG6kHg91T
Fi7bBhRMzpaVaIWiVtQb9jgsNmPOgMB4MzEvWnSpap2OhW2nW8m07QHO1E9wUXxy
26ArLr2eX/rDfpPHMOGM2IS6LHG373XCTvYVNFPt1LMzmhK8jLawuU6vXXvvfX+5
Pd5/FfNPf+OsfT5DyNZrE+Mg6JOk6W0glhs1rlkyPLdEA60Vciht4U6PgN7DGqBV
PWXTIs0SDS8riT0yx9tHP7z+B6t2hycj9oE8VrNwOIDyFCvG3T3030eKNiDFEBlm
Bd4dqfBPdtuJ+8v7kEItjZHwZnOdC/9v+ciYw1Fl1tFiAmPRWrVqMhpxXQCIsKme
mlq68GMIbHWnDl98j+bG7fQCpf2eMOGJ15tgJK6wksXatc5koJVGwst96YlmBtlZ
p96Ueh4N9fXdbxl5D56AsRcahEeMejwQj/JbJNnRZ5QVfyKjxMX3r5APmcdf+Lyu
QFcY5x/RoyPxGmPACdyObEUhwZER7uSzDGzli9WpFVzaFJYs0CbvV/8hUWRVC6aJ
qmfuo9/YqphwdQFKEkRX7yzC6ES5P6I1UaP9p06T6V1U4JtoT5wQMQYfBUhGREmp
og2I9Rujoe0Uu8nhrUzc9FVx1ScTcqhhwPqjtrR2wnewkulI0budly3OaMiHrt5W
dFAl0jSLG7EOW4B/0XDLaUwqLPZrldV2ZoA6H8nirQeSI9TbYPAtwg49xhpOuQO0
yTPv+i6L6gWoNlvW8Ppx0dYpDsKhP4lSGXhcUVC65doIJSmPhr073WwRhSPEZVS2
qhv1hIa+IV/jCWWn09HEwbYsTVnvlI3Qiy2DrheioqYcFYUjrtrGZtJoFbQKJ2Mr
WuTkKuj9QYEsGJG0XP6PcmUYmxpq8KZE8ptt2549P9KNVAAustqUIBkXtGw0LcAn
g9hBol3M3Fra6eZ1qSPR00+B82AE/e/Pl8PloQ93k3RrkkyOAxAFHH+YItjXePsQ
EKyjtifGymVYzv5srztJzAhvGIWbAglcGihGgPFuMCalpg9OGB/zds/6Hnlgrenc
O7bVejIPb9/YGwS5Op3l98QOfrq0fqcyhYiDGSCA3iR0z6+pI/C1Ysxxi7a3NlVv
RbAyIfQDN85a3lXu1MPeiXkj4q+yaySXegPN84d2U8CTjE9iy5TBeVEs5KyaRA7S
f0BIUyQ/R836m1c0+rAcs2MH1p2bVJ1As7Tm/gGuaC1e4mrPJyBHTnnUqZphBLdV
8SxQPjtrIXdwU8e1TnjxKlm29wshGom08hmX8X7Vjg20Y2qi3WNxYvP57UGAi0Xe
sRfdVKWwGYIdADyNa38MVohomvlhtAxvG8QGy9Moiqs1HgWeQX/fkB/juVSmm5Yb
c5ppTIDdWWC4Iwiz8tMKA9YHpESEsiwl0ksbBz/SQi+Uy4X8x0l5wQAttXeNzm4f
fcQwneJRBh7IAEAuEHNdeHOBoLw+Bh3QSP7zrm9SEM2nGAsPe4wqA5kqmBMe/h1U
lxh/OvZUxtZFWjrxeweV2UkjfKE6L3jQU88JYLHXbcs22epaLgDgvsJl3E5HzdvF
lerR7MOEhRPQ9whlyiCRJ6lMCK+4G2aY/QEZPkcWSYMFOMSxqZJWNFxWONZkr5mB
dbDlmvckJhSKEzKXvlYv20RpzPMJbSosRaCR6Gu8al+Vxj/FY/krhFXbLPK5anpb
07CATWtYoxcHu9jEy96/aNyv7rEJtSHx4b6A1SyQwofkYEQU2FlGREUkQGhrEd+K
/NCuIvDiobGLZvpVUU8RnXzJFL6Ug/PuuNN5VIq3eSlOA1Qbu5XzfRlfmpe7DLzP
A4d59GHkHJ2I03nH5XMQ16xlcVDvhEBsZqDEo+psKYQz2MCWoztMbLwIEc+l3FHc
2IVWbx8mc1naiAUrqj2vf/lHsxgVHRiID4KwgBB61c7OB/t9bKBxLm+yQ/T+ke3+
fKbcb/l3uyi1YjXbSN2JvEuqZCXoZM9DDwxaLHn/ZsitCWaaaRnnQ9qqZqdxt4x1
gYxzq3FY348wOJTFWhpwpP1uezozDU20FfJspo5I+fKhGSv2JkToO5wT6U6uhx4N
eQlYxVMfRwOh9O3iGfFyRHNdj8dNbkd4kynlnT1Vaay3C5TIDHvv/3SdrvXC863h
x1OabBWPklEvkwfEiXo9/EHwTGjVyr2XU3HcGtH4mfinIk4nX7Cud7jgEzeMhiwd
BJ/Ss5lTOGrvpGRrpkhhuIIlh2PLcAV5UsCDsX9mFXz1VxsWTMy2sI2T/hFSBP5h
8JbCmL6F9JwU07R3pVKMBWYAPsNShHmuMtdbPDk6Zi3Ip01nstoXev1vQpVenHUh
4GhpxONLhxOADbFwmXI6TODWQZI/L3zNFLxqQcKKZBbidHlpjN1zoCcktt3CoEWg
e8eXiqmHw9td7sFVRf8AYMsHQA9/b/NGjPGRLu+dIeaZUEqa1649uD+KYpCyOxS2
BuMuRzjd3fBdp3g7+b0Tjid5b/12VLq5AtiW+7aFlJ2DF3wV1d4c8ufKpjXP9wc3
quSyPyZwr0Var2iI2qbq+9XtSSTdA2UyWvBjFEHs3Q4/8L1xJ6jqp41ulF0j7bIl
LME71UCHx+WDk7mTIu7XHAB3JqgZHH3knSuUX2I040hT69G1WHKJF7vqBgB64JdS
E/FBwzCWOen9cqH4qm2dWD4Qz1NqF4EbTXsYO2JGMNkwSlIcoCv1ImPRYUAhZgFU
Jk/mW0Ta99h6AScTLl96xMqw4O1LTRi3xAJWnjJmhuH6PdJVcY65u+pNkJRLemCr
M2YlR8ScC00NHB+OUpnX6zwNsLbDIapJXsDwF//C0Ik8QH64STvbsd4u/byUFiAv
vkTwoKcbahXFdWBUS/iK+E3RNfXQbNLbFZYQaRvnAVjqZZLVja3EkGsVAyjlNXjl
o6G7n40H3cg61A+s1NCa5LH50kUuN6i6zPZFpZIZZOliWa91bDCjvCdg02EN07kh
uLXBpipbRCWVMgHcuAoPQTwPMhVRtUp7f31BR1YHd8K+KQ+EFz3G5+M/gLhaTmvh
t4B9Kemd9lmfxgzF6psunqYamYEdFxY926w86lPQqE1DDymYVaDPbBqWh3bxzkJG
hQvw5eVg5UFzmOucLUmr3xlV4PK3aCYjvkqDFZt4uYGULKEHLbl3I08RbCoCwJIk
RMxjDTX+Un3d5NfTlpYbez5H4AUbSAD3UU2PnGnSXTHmrdf+DzDyqFqMtxhFv5Vw
FEqwWstOdnsacIwYVGxFuarZsF5jZ1SdDN7K5IbmLrnaqaVvY7IOjXRsu/9tdAo6
8WH0ToBPjZcbJavVmAchsonHcKqYvQw8K7BHGpHs35iNGwetnET4Ahf6ZwK9g2vb
/k2jzha77J+2tWoYasuyrFCXUZ1DckGy3Ar5FE+OFglqSGdjqlE58bZzuqrFy2am
OkjNZho0KcEyTN3NEkK0kzpCs1eMclifdvLXkQRF4LCwOOQl93/DBTf0xVCzNpyv
VU5Y9vOoTg2PuCpbBEr7AeE2HRPIvLcJ89MR+B4w+7bKWSlwW0CrkOu+TT2HyEx6
hhRiSPISIFaOLxZ0nlrS1dEoj54b5LrLqHxEzBfMgd/2mFc5OId+aJaw5TLOiXDt
0uVVio1IuGOXgs0soJ3LhNLT7OYTLhpromFyrOxMDgqCpZdRgnpGM6LQUi+cDdql
/mNuB2O6rGMKc9RVG8o8xqM4XSDjlw1+wm/L4K/MSBZL6lRaTJuSsyzZRZks7YLZ
TxPb+YzRDZT9kZFxnArPmQPRrxk1JbCZAasYlT8dZZNIlrEL26kZDP+zq8gdSLzo
4PCnQ1TEk8Y0srOH9GTlU3kxEudixb/qASPaOcRI/wzXOjFXOfM0Wg5g14nuy1ym
yhPUG6RAYosRE+8CmH3U+88HnZ6s65tTXUZt1USIp53DFj7N68SxE/G+jmeUdX8n
6BI7HKKVTsEEVm4PoMzDA412DmYPu7R1HDWy4i7WJazmuAuJmc0LJi3ihLq6VnME
M70T6AAsIsC5EcB6EL4PtGd8lnTbhM5fBOyp7VKHdtT4lkhgzphyzW9TnDlFqcu3
BvrmqBfC7BrSgFPq6niMET24ZPIxui4tPjO25wKgCETo+xwbw4u20rB2gyniTWTN
QWhvFQGj+UpSdNNKuvImMoecIIWqaLihlz699JPh33S7jmMi2uj4juLvhcDRqyTr
pV2uvxjdtBbQ94Aqo4BpvkkwdRCyJg8PEWoEtDs6rqxbaMx2epQb94qtesGqqlyj
gsMq7ceywImX4G0BzrPiCAebamiHAu5HqNqip4D/is9brFEhB8AQIDxnbuBA+6Up
mIjs2goIPlylGQOwzrQFeiwKHxtZXDt2LXLtwvkabw4fs1sEYvFccW8JK1Hc5Ccc
IvA0BqKtnGKjEuvDQ7vsRYf11kDfmeC/XMIP1rE0pI7JRHjYnwV467Bk4XBqFbdq
37XfEMpfWDBU5a12nJ9Mf5czC9alsYkn3NGVVGBH4i4q8cLMOZ4r6ha9/AXYlgym
7JqHXETluGNnd+FZZaE+j23vTNSW8ISND8NRudtXWGfMt00y8wrwwkQya3eMsEOq
8vqpBh/WwVjwH8P10Q8MQj9W0Y27AwusItDP/d24BAQHfSN2/1/JswdrKsWyEla1
1zKYM4O24qvUuQ4+jYfL+tCRH4kdMaHzXx5jpEgLt30LWiMIt85q+kkZlkwm909R
YAWRBuR5Dibux1mGK5Li03GbbTYI750yroEzMuaV2HrYH16JBvy8aFn9aIh6S7Dw
vAqkEGeVM6ni5lBj/U9axF5fdm+jgyZ6FN9p63iqy1gmYv8PoOy+npHF8uc4xkrf
ieGE6XIXpiAUwgNkF/yZxmAnCrDMTkpSw0B4VxPId3l/VB8raLb0KYBQDiD3qeIa
XWgH2sn1K1im7Lc62KZJaK6eRWQxg9+rW8dmpWG5QEIM0Fmr4TMms7v2tzF6wUa5
1Z3LsWKDiyaOLN00xhYY4riKcao5A4uoPof4//Usj5Ct+KuAqq7wVuwB5Uarau7P
DLQbOVtNhbRP01ow9TDvaDoMs82MiAhTmlo+ZQnbpiImlvL9XX1X0J1vfBnC0f5D
F5u8kfUs7Z6kQofMqgHm5dQn9pDNByVxNEBAyH0QrrnluBh82lrunsAqs2gH4a3x
FtM9czBM2JMnTaD2msqWguYY6X14uNKS44lqoemvWbQ9QsVnjTSSpfohos4H/HgJ
OUczQPSsonJuFi65i+nDsdVhm5o+K9pzEKoWGg3PuxWnIeOaODkfVTZhgkIox4KV
Yhln7Ee9NXSzXdbfej9hoi5T2YVuy/F9ewt1kXO8juhpyoM9YDIPQl+JA31FBeCv
HLvn/wg5DuzZXi6wBTl0eyT5SmMTrnaue1UEn9RYyNytbB56asCXmeFXX5G66efw
cgMgDYaG9BVKIBe4IDrfEN04SnyiuXliPysiiSkNWiSSVrg7qlo1QL3FEd9ILNCQ
3SVtlj9MLeRSFkuUOuU14++XoCbJ1xqfz5TMb15PqBSJyUQCfVeKsohFxrDp8a0H
VGKx5vtf3FOWFOEALay7OSDvsXk2ZT8tZwb4wOjNqMXRmjSNCXQ8tU4eXsHYsZqu
f9hp51BjCH4T9xRWKVF4WRIwcW1vxUVHfpPNlcgj+r6Svu3WoEk2QQOEGGWMp3XU
YbW5XcGqnEEosG/LxGxYdqWiQSREoFVxiXopUtKvyin5qFcm9cfJlTrOou7IxWjS
PLWymWR9TjxeOUFDHadEz3M74q2iaf/pOH26qQcgNMuIuTHFZQEHg0IKWxdTE6oI
3412cXVa+ebia7w6jAg0twww1Azm6C0/7gsUNsAH2h4U9AqC1/G62CCyol6i04Xw
9tAA1Ys2tCrnPDVkAVbrkohT3FiLG3vIK4+SYyHbPn53CqOPWWF0kQ52kUGgl5RG
R9RMeRjiXjJczZrCvBycETtFyzGP/311znOu9g24ndsBY8WKVloPaFUykJ0FVX2/
DZkvhzolk576gp5s+T+7LBJw+r1tZfcTfx9O8f+fXGxFAounCHNO48skQ2cWrCTv
LbPX4ICIoFJIdnEG8UYV3w2MmnG1XjUBb6aZQFV/eNEwEk0HbxbpTtWSBqMvAmsx
p1mm/9eqfytU5234KiBot1b5zhNUw0yYzu997tuTfavay9go/4GwmBMpsFDLyNmT
G/dh7Xu2NH/Qsgg0ZmG3chrWsl0dmacs1M9GukNJMYrXgoMgWB/nZWlcnCL+x4z7
ONOFrBBsTiNrDuoJkknkTvTGhVx2Sb+WabL9AoACeWKJ1mrp/rJJmAfVP+fmJj/B
oLUVPoBbv3jnkospdpSDqXlT1ozsSiLwzkja6Kb1Jz7Ww/Yp5ewY7Wndlgm+nco7
Fix29KFB/I9XiWbBJgXu8cChMKKx/r9KJ2Fg/GoWUs2mRqk0xNsMmbBWm5m4lzlv
DfIhpVLAz6wp3t0NkRsYBgNFy3EeMcCWaKIOTZ57AkxvbGuTJzGgSc4DhlZOAU7y
PLn7GbPh7hPU7JVF4XoMU9pEthLgwQfTFQwmzVGyEK7GoRWYP3ZakK+qrD293gn7
F7xT785hQkHUiVJbEinAA/sXNCP0C7z0EQ4/jaaoP/4L9JbKt6jgQJMXqpC2HWZn
zc0vKSJpNa5dSr3c4qF4U+sPmbojth4ImxnS727wa7yiK9lhbsBKZ0xh3BAfeRg9
es75YsRcGW8ebEVYaZHfeBRKQX1InAG6NKJcgPTWtMwHOxBE4Qa7aQ+9Apo3d1Eo
pKQTuELMHBvOSPHZUIhgRQ2Ig/skcs3OvLVOLFy1rfobIKgy+UC+h3RESG6unhrg
XNQWrLC0/xLuV3e0JbJbQVc0fQNuXDUwh/FZNZAf+bPuFTsrBhdjq/A93LmFbEuj
/QA8Ite2DYCn31nmlNxictX983/rMAjyXz7AokilZXF6n83FlMyGD6hniNAkJF2n
hgSLDnw1jOg7maHAKiVpCCKh0hftBV+mOo+TCaazdeCeHtP+eMBP5CBZgiWppJmS
7aNuXDTEnQntgJYOWRBT16XILiFoxrt8FLy2/q+yMNzJmjowr5u2rZm9YfARSbor
kZWSRPER+DwJ60k1vea/FH+VScG/jgW1SN2W7gqEYVIqvjKCvqobiPB87B/GklBl
RXrQIe/Ke4WjZ6PJMFYXtbi11fOGfwVYJEfB4WAT+sVRDyghKWOvRDXcMjTxm6X6
+Y++9JOnk62tn2LgOPDTKS08j7G1EPlo86N5WT68YKBtaM0ggOtkGKkELc2dgw7T
Yb+l5PrFHfTGQdKPErv8MRKyix6mEgaFBaBK5BRyYSBvaZlmEKexAS2/ezTuzPtu
DSnf9prpZdn8Lg0DjPuWjJgIj6ZYbAsikCILaCAMOjxK33pERxKDcFYAD8LDXc/J
Mc4LVPT3C9YXW+pftoQBHcoj4EVThOFyteHzBbyJGQUCFUjdv6WJIs0e+N5roSCd
3RJrlWeKP3zB74IzRvHyRcF4noPzSNPToPMxKiHH3odtGcmiqCTuQ+SegDom25Wx
bS1eUntsTSGk7GBPPjhNXuFfAHzZA89RDq1DCT9NMH7KNvPxAAVZzrLrm/WjZmxM
xHmxp4VTGw7IM1QnU6Kh3rrI6WVm7N/EXmYg6cYo57rpuWnkYpY2FJ1EZ8KFL1Do
piFNIGFDY2/zG9mBGMIYJ0YmDLO/YYWO5A8Vvjtnn/SH87c7pge8AnG0BD2/e0OT
HXvuSi1MFt7iJsNZUu556uiJo2B6v1cj0APB6uXhIqoVlXEhwmXKkZxB0lKOMccv
ZA4+/Zxr2li9fAR1gFyBLVXccelPXO7bbMJ6eNt3YxacmldV/4FylpQaxgrmXMTf
WD+JBrqAZBWPxQ6TVByOSemKFUhIW6uKOV4EXd+aVUBHjwuajAD4U+zKVNznrkhG
TS+QGDd8se28FUaVswC4rWh+TDx4m5QtDbH2Ki96WA7a8gBOA8xfX0scRz5EgkKf
9rD2j+/b33++ApGFzEG+ZAOsNZWRs0B8+kOtrTDgLuVbEoHnbnp8dRonGvA1+Hc0
/ZlyAdBP+SYsU4MH93RGbIF12qUVgjbZvXu9DroguAP8kspn0T9XS22wn26CLgaY
ijJNsDAU+/3wYpqDAVtW03jrmB9tgKE/JgKXagWiHVTbTJFVVo8MjbH9P5OlM6Dh
NwyMMm2kLrwPcdAOm6Bw5S6NUakFeaSd5Bq3qoOGC6FokoNWCC40U9jG4li5ZSqu
x6ELRjYrFX/fkCnOenKCFpg+RUgD8R5S9yxBUkSnOYfMzQcoEOevezZ89EiHP+1H
RQTeR5eAjP8GTpFa6lIsLpKe5rz9mtxAvjYYOHw3H6v5nGy73oKBVEPQjxHMcReL
LwaRlRU72SIX/NQNshVu6qXIFvpyZsYmNaRw+wA6u/ue9XmvmWjyH3cUvTYtXeby
m+2NySZZKaC2ndOgU0Ji2jvevajN0ulrbRP/rFDxfzazBr0uUIZsia8jjnhkkhU6
n65S2yNaN32d38of1NotktINnQGuIx0L1L9JusMf6X2hqs2KRc87lhmTF74IgHci
o6fLhg2QTw6CMblfU5tnxkt/bY7VzTA5I1aFF0hIMwrpTVwhB6iWuorT7G2BCP03
NLbq50t3vcH7DO1UFAY7CSfU7mro6bj0PlML1uWahgEfVZXm3Xyu6BqdGxo+qP/5
bHcLQ9CEVlM4v7uh3EO8yJOeeWnZ/vJLD29QRjm9PKoGQiPdXa64z90eXH6PV0kk
4AuIFRrSYcd2JttP00X47LK4k+7b7QlENVwHjfnfk9fTvLK0FscyNX6JKxHj0j0I
qCTSs3ywfs/pVRkI0HCKfSGjACyNYN8q8cHkNobUUOjDB4gCLQqAwkjsSOmLeUXD
Z62z9kxaNTUm+GBt0bq75aq3PSwqTBC9QbnLCxFM5PRPZb5FV3bT83iHHQyOIM+X
GJpYzAS+/VlLxU534VDJzJtsMJHGuMjYGISyL9y/Ft4a4Ozaf4GpCRfTdZ7fZ1j6
NhBKODJUGQnC8t4KVA8j+Nfkr5F/TsDM7efyupiuIG15uqpJjNovUca8MYuifAdJ
ltX+RZiVq9Y2IJGkF4KLQs4Gfc7Wm2203nVpy1A8ct1u8qK6kbe4JX5MRDlepzxG
Z23tygQNKDDXxWwBm3GUyCufah/F1CWXvLTMq2XtLPzXmSWsuyzkJelHivzy/Lbh
D1Wal29uzrtOYRvEBL93J6VaCUDquk3/gl6oqJ1LZERB7VbZUjVVEv7fAS08yKzF
5sE1xZUGtvP4HJo4wnpcV+uTODaCSKZdo0qEiEuiAY2PlzMrfaSI1XnAwX/U7+2q
lrog3x/bkt6jDiX2XxNk5BUPeLzDBNR3GnJ+XI3QIRN8bsXsO9/WxS1LgTYVoW3a
sGUWCbNi7lrYNxBT6BWt7gshXbAGQ2cQ89F1n+APLYifDiwfL5GYl+lynmtA5Xak
G/g1859Q5ndfGEgv3Il2jxaO4nzm8S0+b4+GMDBSPiBbxBMZ99gSKM9NhodNiHDG
ZYB16z+n8izgn+s1gKXpfwLIGFnYQ84DKJCV/G7Lpsqwb4CeJEr2Lw24NdZrSztI
SfHHYWgrboMU4sehE1ct7xGoKa0ng3D1Q2HOw+1wy4ab7CRQXCLR+wG35KvrFdeu
BdAkFIp6o6s86pa81YuD6K8lJqWbwmUOEWH1rBLtC2j1CEN4nKq2daE9fqRzjqnY
UnFbI3M6GxZ2zKQoo4sC7Tr96Ow9N9bg6/9Pxxcr6s5x6mdGIsy1Brcaly+837hD
x+NF6ffnobA19JbwWTg0ja/bho3EOpkdAAVJC2j4gZPskm1IBTx2AcEMheeZGo9S
UWWM0Hcu2qZchxse8w9CafCBZoOKQtdcH7a5JEjCKwI1pJV93xEt8upU3T2BwMdT
kFvK1Oh9eIFceyT8S8hY7YzXhRi3i/SV910/m7D5nQHlORInb490kgb/lDADPuX2
ge4XIlO+gDdqQm8Nm692+ty9qwuq7aO8dIqWLzXMzucYRFX78BEVfhIY5MRm2j8F
obM9cCiBUGjJAymR3fIxttCnSE++tSoCVjanvKy9ScM4/zIRXA3km8j0d5AslJPm
xXBgpkmexkw+6HVLRuF2BywEBOh0/G4tRQFB+0eWmFWj97OFk06I+OfD/SLobqcs
0Iy3n9Ocv870OtjMDasGY9nyYfMCKsZJOX9jCxVTmV1SusH0blIb1BT3uLX9NItd
Twz020yFVtxsDfC92KhCNdsYdGNHOakMeqgFKi10u4cXi/ft0wXstuIXrVcZQOUm
GT9CXk/L7blHfhvODH2c+ogYCmU4PubPcN3MZ+qKfHN8sB//uStC1RIDkIrfeYVl
PC/7gvfcusHxXdoJA7kPLedH0e7hFnltrzFq1dkFqk+fAYQ5lU3zFCnNuGipcbnp
nbq+BGI7xtNxWYBocxppmfXiqRei4YtEOM1S+cj5CILUzM1VWqy8txJ9Ffc7TrEr
je+IiSHVWXgLux7RskFhVdV5GNU8qxMGiU8+KAS+z4B3FXjocv87OWkns+vm1Ykl
dKaGDRgjDA4eGgNfDm8Rr+kZdEPkdvt2i94AnSOEUSWeHSqV4JuNE9JpHaph+Jb+
0CmQlp6VKa1ht8kWwQTfy7a1W6OuiMG9PoklBSv3l1lfYY8nLdrtGGPEY+ogCP1M
/yE2J8gMNxgNUmz3xnx1PPxIaT8y/4sDNeIyKc/0ijKoxRb/OBsnxGwyr2kGfZQw
bDsknHwKKDrs3U9k9eWDO9d3GGdq4Ocn35qT+ge80/grj+FVWV1KIUqFzIFwHkRd
/cMURAPdAhNUf/tIthSjwhI6adNcO/Tk8QfxVn97srBCi8h6+j2uYL9MI82MZaG1
XrNnvgGQNdOfBTtJ9yG3ut57pngEgSr15z31s7VyvRulmKS2tE7hqcu5mCWaMqbN
Kqbk8SfyolkHqJOUxvN3ETT8H2dK0/7eCPEEPeYu6DTO1CLyx5ho5ola3tCWfgX2
mtSptoSaSrmhFAgDBFNaOVuno+OIM3A75SVvu3SiSWFNseEDko8kWhE4UPDW0ZiI
PwGOLX4/6G5ivF3hxT5LcZoUPg9WoCDmtdZvPg4UVkVf/sjFFLKDXAF63B1Pw4s5
4rTYHxqgr2mCbFsChDJY0CTlRyP95C5BJH25teJjUH8J7bJpxNXUt41gDfrF62s6
gXTuMS48KYMAiX9VRxZqFADTSGx9k4e9FzM7CVgteY8/BcLNoFuyASHqp03T5pqU
kWDCIkb8sIcTiqy1plwaMA499qXS+bxn8kzEMOJdT8kep3b72Seqa4k5TeNAdX45
QjxDXvwSxjGJRMEm9oqRQPRPwe5PyZOa/UH6H5kLiLpwKzTvHxERWzxhI4qSb/ES
5gFA8eb92TpocWtQW+NCYr23sLySV3LNvt3cOtoXM+8gDC2VPGbHvbDUTrfFvtL8
ZkGeVaV8hbaqidltxfvCAjGssw0HR26c5vo5C7EmRNEdRKqeg+qMM8OcSXsw7f/I
+Tgbl/JKfgY46fcqNQty65YHVKfhEBKWZlxXDIXJJHc5je8QbZQCHZPpCROxeoar
DqgB0KkhMmYTLPyAKjyNir6aRuz4QRjz/hN5i6H0c/hyPFWZL3qV6aL/ISw0MrNU
zihRYxCmlhF3jZPi06tiENRUcLp6777ZxYDAy1eiO43KCrneN+Ys30UMg4tMvkLQ
HbPbdPw/5cVoygBjXNhc9C9+x446rnnragiQnLSC+zGgvuAw1S+tuSmG5y1JF5C5
77slrd5TzAxQwR8xfLjVGGqJytay+5AvbMVU11mvNac8hJAh9C946U+87NjlW2NV
TNtlBuksAXyUwf9yPP3rPdpprS1LOEvpHxBMgHN8HreFKVGlWfPB7Q/KsgbR1lXz
87/Wg8jbFqM/1jNuGUBQ6xw5YWzAejXq6z9IPQk1Bn4NgAbxjffqkFkyF+zkncUw
nj0cuNYtIjyQp/e9cUi9QxuXRg/5D3itD7KybbzVU/1++n56A5rWPiWbR0p02Tgk
25v+vhQwK0LjzWfC+dMuh0/EnX4XyHylm+dLomPvcy9aCFRs5WB883ea9wAYXaaS
W8vgGGB16GwB9JUsVV2WjHu3Nx9XJHLwNsUT+fwEyyNk187Wtp6qamQr/Qr9BHFB
V91uEKdHzkX0uoMPeG9UHsRhNNtPfVM70yoyXYJXhLoYGoRJLKjBtS9hspax1ccj
mYCkMn1BWaPpn7rjxFehc0VzDKqJ3GP2cbIy+NaiRrgmmTG8otubz1hiynj8eziF
VRdZ47H/M7cBVPGlwZG1KLIET+fM8OrHZUIl/chV7p/LbEmfq97O75tSi3AZjgyr
83LDBnKwYS623P8ifSzgTRMSJyRgIxJ1Vd9uBAZZ2T52m6BtBP3iSl5F9LOs1MX5
pSShINMO6m21ny9KSzubPe1sGc95a8Ets6ImZd1kH09516OoQ6+27/fYza7kV1EX
Wi4kHgSGLTMNE0wguH31N2cKSQK2LIvDIldL9z/+96jBmvCB3fHIowilPhWT+elf
4lxDuSy2VAy9ojB9FEOhPQCGN+/E2fvrYg1a/YY9ULpTVX7dLx/PHCVX1lpKiiNr
9MaOfwABktE+jW/AHvAJ6/k5mSku36UW44/ymhXn1J6gW3SIIHL4Jlfr3zfvoOPf
PurDXrAp8HVfG9glWh5rmoS7C8I5Ztyk/XzeuEmsx7cwDaZoEi3Ty0gTJztqH3O6
FCvn6aot5aD4J+gKUtHYe40zRrJ+tDcAPhOm4Myejz6eKxGvGC3iwTtedxvsv/4j
frkMKosdOI1H8zcO0MvQ5fp4iTESh3Xg+DWOzxQgPTnV+z6JXtIlV7kaLhkhrQof
J8/nHHDfHQIfNbnNaRli9GHDovaFvLi4D/HyAXMYNPk0XT1j+bQSFDbabezfi4Ao
d4epuurD4yU183d25pmqSGd1HxNw0XNjhwZV4i0/rkYp06KYoLr3T1jQUlK6zI6g
j5mELWw4EF3FBEMi5Pwp/ze+fMKgtsdBzoEdug2/9U0mX0L96Zvvd/nxBqp09IUs
v6sjHYgThdzg0wRIbdMOBwIAs1TsjlsBx/nV/saUwcpko3v0OBzXcFLxcuF13qZf
3o7H1X7f7z+P6STukApZVDgEeORBZZxuSL7Z3Y9D/KTzgdaD1d+RjVd+1Ccbj2R+
C0p4D5U8N1nweCl0HtQfHaL2ZeYY2xJQbAp+kg3DZGzdWOphS3F7enOUiVf3i2m/
HutuAd4FAsRNWzQgSBbk3xXT/j8uPLN1CnoXO0B2MeYT3VEv2fnMRbodgSLr9hVJ
RH7fJ9L+4oaWiNvD4XK0X4z+DSlUcDC/qJcsGbzTlka/XpSxBKvGBq8dLqSqDi+B
riB+iQ8g6ScE2s6nBiypu6exySsLQB2LcrEBW9Rl8Ar5t8p4TAUNq/4vWTjGWCAj
zyJqTa4K+sNw4K3m4DoVjbubWFZkyvFIdUr+0x6L5IEB7k12p5aGxZsr+Vru8+pG
+mIGYkV3lzFCyafxyMtql0mO8qgWn0UcNbKuMJ6GEl1kNeqvjJ8OLchE4Na0sSN/
mQBzR+pe2waWpuFRMPN04IAKOZZRUdEsW45vjFX6+lXDgmWrq4p+hQZHjmwa3uiU
K6hd6eJSGCzN0IcZG6/u/jSm60PVslJJhUqOqZZH54smMwYH2GneuxTQmmoDNWgM
BsWQeyw91BOuKQnRuwN4sCaGMh4KzSHw97JEK0tr6VvMJ/PXVtvHpLMOH4jCKqiF
ZjTxfr2PBwdcobOcpXAksyqhr/CFpinlQIPxLZmbkHEBTa+iqx7jNzODvDLLMsjH
S/nZn5yruH77YXnhmMMzDrESDsNRFgPwHruiYDIUzxK2f3HZ01VG+dhGBheLmRJG
XTtHBjI5AvBWZVhXQ6XykDgXQqielcYuVPkgjekiVMwoz60lpizVbfKNsvPHLsR7
dagoaVh4jJc5bqJFvVylvv4wLE2F4Z1aLRzsk9rszvhT9HJPC0+KP2bTaV9DLw9r
e4x8HfQytCDASJcZRC2UCtw2kHIV/8f5+tC+kW+g/u7fHty9K+HlFVkf/ZExeXjg
j+k1rIhQFb9r71NUnVNUTLcnI08ucc7Dghxmogo6ZAegwUCJvn+nZ21Rk8mdSQ6r
TWXh25F5K3HIfx+akcxj1a854hFpf73NRcc1o25gueEK0Wref4J2FFUjAnTkH52l
QnBW1YsOYWVlL4h/emLM5rHAEBF5TYUdxGqhN9ejiKWlJL23FpT5YYZpJmC4cnX0
S/rWFefze6Miltmui22uWC/xpxGd9nGt/Pi6ZbA9nXcrG97gkxwP5+ONl3xdH2s3
zcpQsBJeiP/egFTWk+6Gjqyg2Dil2mpQD695C1ec8YxgtwbmUaDi+Im0PlT8YTZW
GUBPXBEH6JG87rYPJa922Cexf2b+DZOvdYaK11Ri35GWaJ95H1SO3ewJ/dAB0GFP
AhOLNfI8yjic0DAKojpCyiq8vduPIctAnZP9rHtqY5G3UafakWpKHqCMDMq3keSw
qafOsWrk1kD2koFtJQI6whi9eEXj4TmW0Ijl/zxb/T7zqWW6TdgrBkKUvR/lZYMr
WsRqe+TMDfANvA0nmrIbbAiPddivlKK+L7NdQAu7nuadBnu2QJU8r+TUUw9okyhc
sX44GRNYB8nOpPPlq+7vhRMj4W22/SuVmku1Xy4sr0sOcTTx2S4ngR89Wy5wU/3l
r9zWgG75WPRX9iLhwq9Xr4TGeSYwTXXSi3R8m5X8+uroB/YgeZYLdwicgnK/aXEL
rAKVIJ97l+UOfSQMXiWZPLn6pXfWQNB8QL2byCzHC8UHznvTgLLEc81xPe03mn72
FMRrzULbpC38+z0dqHgLIIjkzVdqndwtQKN1xbh3tC4x3AlA7B9CgqPLEQF0wQeT
5J1fvqonv/oQliH13c2CbpSnpoPrQHLIqr1eBTNRFM9s8u2DB04Hz+UrCvpz2J0j
uPmgn9098vZkw5IAie/YdSvdFz0H4Ci3Dwm6LLZNcsKrvhqKVWyGwm6SZkL1rumf
PLD5UIIBf5qtTuOCqyzBPm7zrJbh3yhWoZeiLKqwdTy420SOGctHFM3Oy3VYS1au
6ik5hJc/ECoLVpjmq6QfoVdenKTIaqcivqWp+L6d9mknkBAM/79mw2s/W6lXxhG9
lSUW/joVKpy57bE7Qti7J7L00HmF7MhRke9WdP1uxeOCMqIB309hw+MlU0uFLAsE
KehfucfXptYcdGXqeE0+skbODt2kIiMaZ70VpWLxh7BWfCWvLXHsRCkQdOxpX5nO
y8W5snBRRhqTqAPKWnAGTtJwS1U6SQCqKqLUaHLlzRQHcDQyRbyVPnARSTI3KSWA
v1t+52RNlNw5d0jNT5LpWQ9ACJFrLbuiY8KuIsV7jckkWo2VQnr5EfzaDcDHz/wl
w14PpkQCYchk9mUyy8L8mYkEzzXVNHh1RQkcyT4/7MA1jLemJxDn1rqq2028n3Ai
/LAd9K/7Hmk5epF02sUEmQ1ypm9W0b+yNFqCyqQQPjAwbrLSLOQjEd8GU596wwdm
DpZeF0W4MQUuUwZB+KPQZUazzMK/wBNPkJgjaNzS5rubCE4CIGqA8cFUiVubhOik
WACv8gk2lnzH2q6K5YTHjjZOwFVdKwotbu4bCiOE2GJY9K1ooL5zvEunXRuzx+OZ
5xKAVC23D5uvGbwuZxb2rNV+QRtcrMFCSLVN0C5PsPyp/Dgalpbq1WcCzjrmWYhH
NkfNfTFCf3r2p3H5zitsEtbjToWCaWy4K39CO3YJ08uH3CotbUbrNI3IjlVoA3ls
cwJBDp6yDBeZGH2SyF7x2xsOsi5NNuLYp9CT5FEJRDgHSX/gdRT+Z4FRIDSj3bSS
GY0394BUKSMA7cMGOrB0SNozFJB8GnpbSo2wraxPK90eWJL1rHrJnf/wcHkMTR1b
RwBCnN1aH11iTPM+Io6BszAplgjozzSNDmWIpOD5+oyMKNUwCrc58aKT83zKxHdZ
vCmpKTu8gEIlQqD6zt5ItA+0VBBp/zO7HF23O56wY1D+LllTlORxa8E+V/FvfWaJ
MMEMilB1QhgkOUHZG7L25y/1DLtuB6HKiV3AYKxq6htUvaOw+sFivaMv3WS4lUx+
dQIWf+hCIMAlFkTh53B0T6yC6CJqmuaLp7Thdn+vV7i3PwArwRof3qwswf5VjDQ7
C/1s9RcDi+1N7tNI3hqyCAY/SBCUwbBWc6Y5wbFVO4oeIAECjBAeAhRPuPFPENUQ
oUytTvhj4Cr+alIAM3w3J9WityDrObeOw1Cn01EeNCwZ+ykJEBPj6F0ehIWfJt8k
aL/BfPEiKyzTaN2YdeoLZfY+H1kpxZOX2J5QeXRwJDBRJCO6m4ktZVaY0AZ8Ng8V
4Nj/A819j8jbA8Q4hDB00XVhpAQdloMMpvHdKI3SmI6yvtCoCyYP3/KMvnDKipkU
Uxd4A2zENtLm8d/YGEpaZqKH0AI0cClOWAYzvmRn/8cHPFj+j0l3he/4NRrZpXGH
yz53ug8jpMKLYdXmGZKj2m6s5+HpVzLN+3Gv29Xj4EL9OIrxJEhxgqMHnE9bSXYu
SrC/ZQreh0GDUaiiJ5Uo+6eowqqtoGwEo3wev7p7rMEPl4mhRTD+2h8sffmqY3IP
nvmPzauivk49WZZQ3ZzBPdC+MrmRs9ctbBosYe6ScUxmQRkntRTmJBw/MgDT3l29
lLKuMJ3m+b8HGIlkUQYzfCSX1Hsa8DPrCf120zqaI8nUtKq3eb+THu4AYCQqrDeT
hE/qHXi5D0jcyFcSH9ftI0m/jYGxKyF93rXWD5Dn5el5LV4APRaWLkqmhj+EArtC
7mTSjov34cLHX7hlLmD+HPM4n9hiGy8VQoVMp3n0UwyN0wZuTdfFuaFNmqwCpIFZ
Vx43P4PzYAZGF5xZl7jrmTGhZiZGZ23oUZtEM+6NcdmbhkcdDoPK0nS/DaF943nK
TxfB0TvMdCbG8ogep78aqg8dvJNJ5pvLOmXta04eQSnKSJ9msj6AwURJnXM3+vLZ
LYjfH3YMxTdwYubokEkNn7S2vGnycurglkYeB+YfBj+mxUyW0ftXo/ZEr8x2DxPQ
5ligO8UUb0RdG9zERkVenTKPD9+qFHfztKIUNXWNFcNJt1F1VUX6d8n9gh+7KO4W
F7MOGN29fFPguuj8a4KfO/z5OUSP0IHbLUkBz9qI9SojpeuOQWTPwQXTT0iaKMzP
WeztBUbzE87/9NK1j996I/EySnHx+6AZwSTAT+cTe48kWOj0QBpLVTvVWkVLw+O9
uUvUxQCZW+JwfZIJZjpwSGTrA8cGAMl0q+MVJsp5g6FBwOHMw4GEvqzkvo6zrzc5
NwbDNdtyfFjWhEFt6DeesFH4uWRFdZli/nCDQ1YeA51vYYSKulid8kKzBgMYf8hN
Reg3a8xf+xyefjGh9CJ0/Ywb1WaFgsI6ySxTZVI4N1mSgdwOTWC8uNnPfF8V9u6J
my0FN3HNzZfabG4dgiHtoHBCRkh5kAE7vChj3bEt7kZkkhZtlBQvVKPKw5RIdiY0
2zUKl0duecfUhiHZTqCApBwGHkbgSewMERUZTc4JfVwuBHfT4JprcDTEOALTSQag
AIIZmxwmnFoKOnGPqUDrjtHlNAz22n6FV8LgIG30ee3hnI4A68cI5tGSerUkKHir
p+y+rldmbe1dIKHCzF/+tHW3AiXZ6ihP3O+12zg/GTFKlNmf/25iVE3a9xg3lY0m
4g7SAjRFV+zzPsv1n3Xmg7odo32L5NWWGlr2iAjVu5rO+9Vn/oo8HNr+RtVSO8Xl
qAMkw9Uth6DQPhvSl1d2Asy4lNh1xpaJEJA21KP2nUVculW9UxvKLW2F+OsEJ/ML
VnRxwOn8Q7sxVIkWeyRAuKpGRYY7FG4bjGh2BT4dc2RFZ+WfaZINVZq44uxqAXnM
mOEXnzESTxZh4qvZA0f4PI/bUuVqe2CyW530+Mg0dRnC3qKUSJxL2QnHEE19wlXG
52okNm8DlEFq+TSQ4XUXnVkSRcBXonFsZnMhvtr82fK/IkahVAgXc66x3Q4DXJkN
4rThl1DxLsXzU+b3jzQMR0us36/z/Hypm94n8M6TinomhmUwClvA6EcTx+4AFZXb
dqDwUrkDXuBs0Foo7hKUVJwDzhzMqM62W5XB7U/KDFuCS2QR3aNzUEmxZneyLFr1
yP3rjYAQPYEgN0sPndoKeBKuldCpPsiwluDCaxi8A9dIAODwhjS4eU5SjVEuHrYl
mKLD5T6m8mIgfdTcnkuQSkWW3rGQsrr9XXnGo0eHTxsDKk/w13CJVTZRgI1qRTfr
4JQY9oIBnQ97HnrK3X5aPZQ4ZOdt07Bx7KT1guVDxVEEBg6Ft2c2AzN+TcZZZgRw
mWdiOrZcSySoYU5Y9bmHpqHvItfMPcPiCv1cfU3DYIcF7QpaDvOyJCA1xcd2doet
t4ngM+ceGar1mPD/LRxxaW/oYCETi8vD9Nd5n+bVqOysd9ZHd/5rEPnAVHHWuwsk
mbNZbeajvwzEvScDtihz2a91/Hcjr/mBw+WrgF+vhOaUGWsdts8wq/9dO24quTh/
QrwL/yet40OvNIj/5urwxB92jF83K6IXVGv12sdcqPBQTmibdD7v5FRUI8BFzyUZ
6cY2HCKHFkajqonWMQcIKYDrFTfeZjo3QjNZlvH8G6h7+xqDUAz4n3hvV4T5hALW
D0g1YJ01pJjcqSsqm5trqHF+CYFeFMCTw9PmguwVRHhSNgzr3tKDBT3AWwAHML+w
fCitpQ2HW0nPUik2BCxS31edznZ0a/J7lUciCy3Klvg5O84RW5MEqFuI0289eCiG
9jdPs3QT479e+k5LsgJkqzP+U5bQ/fBgoDFQ98eZZoB0WXDK9fPRyv8JkBdiDWUT
IHUGITZnkAo0y0vbjHTBDxLODDXOFA+1ke8WjOv15AZJDwE87pUq8jiU7l4zeVdD
AKHsxz7cPwECpA1MftZ4fyTbNIee6RnvK9IvQed1p/B8KuepoD9Jqb1akhxrGQ5X
xNIEYBnIPf9eZiN5qOd9Wi90NUA38i2Qw2EDS+UO6fYUlhjUErUSmBgnKpt6156j
culYxUKreiIXD/WxusxuG86l7eE6kP9Kud0WUuNV/Au97VCP6eX8YExyCpo6tjoa
uBcJ5SIgbe5NMIVhtZMfLsq80RvCazWKvi3BgZ54QegKYcvBUns0uJfq7lZ+Cnhb
O/SDYdFTHmjZWqZiDHp18Qipq6Kgq2P4VvnN345qTHbzf0mRcBbIcSEnCOEa5xPp
IQXremm/RfI45zliX6QoeVNq+Squ9kRa5OgUC6y6V83Uiq7A6R8OVvboTWmSYscH
adu4RnzR6OYfl1FaU6Qhj7tq8hkYN/kNX4f8vprEsfbVJoqbfseaya9JphrkLJcz
dPoNpcau6neqj5vf7dQFU3vu8cCV4bCksip8DrsPOO/xHtZAuTrEJOnQms/FhDqR
vaNzd+Zf/HortdU1aZ5HdfEFLv+agQVJpXdoEvKPMoSxAm/Ze6F2GDv2LNXhyBjC
5rNT91o1Xu9DW1lyC47q4wxtkLGhNg52u+Y5IsByO7ZZJXh06GqwchNl0W69/Eiz
pOop5QWuRk0E5X0tN2KqjcPTN+scM3FLpnDnDsIHDry7zJorIDgrQg5Ehgy4l7Mw
pDsyPzPPRzf+wpjkU2KA78upmGIYxdMdZ9I5i2W9reKLWiEVojuNeLt7CgJysl+L
7HcNNyjfvQ6T5Fq7i6lH/VDLpFkogpwBjQhcx/PeyedyfNa5ws37BOmHVlcRjhLG
aPjG7PJ/EcGXlM+liVoGJ+z174rcVnyzPPh+AFF8PL29riLnpBw6jCmTye+0El65
4iNe9ZD4PYmBSgafKtcEJzSlzmAhDJDgVwK0tE2Gb/Xvf1/KKsDPEcSoxJPANk9E
TlZeQq3R6o7KMH/YU5crPl6OeBZ8I8BqOQZQp9o+Ez823hEglitJlCwFOwbIVoin
kZeCgxN54bo4OsjKhrBdS5qi6qIK8vgaBFPTlPUOy0kti2P+ox1TPbmqwt2xpkur
hcmsFRtMZtHgV8zNWfZudN/J7UMiWs9H9kItBMwsrhz2uSUf4AS09qQQD6WH7yd2
6RYk5vQSEuTN9VUJCWPyLeqvge7hN4JD4tMcBRsHNJmQrP73dqPzfZH7YH1C80nW
j8SLZHQB6g8I/0y8DNPQzCNHthl2TSNpse36waufX9p36YEMptav+FigWU2poQWl
YcEOrpSsHegEjhncJ+/XlYiEHDKvQ1rXopzugU/qTivOzPcty9lgVlhQqxAlyXs5
WK9MY0mFZchxuda5F1tZQrG+68Nnoarg6uegaxV+c/vWmXgRMu+92MprtilbjQex
jn3qVcFzGSdDFyhmotWukHq7oIklO3LT0dWP/cOUYCfVV/1SXwINvFmAidTq1bFs
P2mr/py3lQkVRAMDgoDkiTMpi6sGtpYr3YsbX51lUeGzfHCHjGbfoclsSpgBBY79
IJtURu/de5SzY2xK9QXb9KgNDW/l9EAj3biiLeQxXe4lzhkHx4DScd8wk2fllnKU
+FpdYNzDAHRDrM+Wk2AKOzLCKuvJggs9k+iB1sM2u8qnQLKSOj+fA6FGnKtI5TBt
UygKLaz8n5hw7yQbPC7rzuKAuBE+VljV/17GsxbY/9jjHA/PmtNma8LKLxmxx5DA
pCl8a/NrsAB18p5lyKWC0Uk+kLvJTIJJz69R3zHaO0IgzmPMAeZ9D0GgeckXvLSJ
yLCyrE3Mmy/3QmmhSZul/hpyc8/r4Z5qh7dWkF/OUugX+e9uQ5/QxAeP/VaUD6Qm
cWOSxrOcVXCFXxS+CPEwqHXsj5uZ6MW3PjnMy4+ZnQup8sjDinGwIIIjF1KwadIj
XLaUeXEwfxXnfcmfpVVWBP0zkuDNo5ecj7NGEMHdtNKH7A1ThBrqmF3CVC/hiXox
nLXg1gec5qCQabG9ZvfyoJd3Sg8tDgZRBuEZTJaSgbEJY17qXYjawTWyJoE/NLFV
3AlboR53mtmfg3J1gYY0YDrrJkHVl1M/IRotmkzk3LHMECx5AeVo7hzTGnU3igw0
SXV30/hZcKq0PHmGR9yrX3QbdAs4FuejVSNvouwLGTBvHg94heIkAph8Jm5wGZLz
vi/h47y8eJ/1DiABcKqdvc/Rw7J3oww/pQN2POV1sV2FtHUd1xxHUCdt9u3nvBJs
fB1tacmx9cxqp3dlEmObk64v3RJ+2/87oMAVGJm/cWZRN6PgsY/REg8wcU1LGooK
5J1wD3UpuuK07JvR9tlPF/5/v2Lqd2Ve6wUKVX1Q1EMsnPjWuLwh/8v2xMCQFF/o
4IbOTHV8qeswzPcrjTtrkUXV9GdmXC59OVUCqf2ovNvjLu/nRqhIhSGe+JqGQxCo
usGMRocO/Lvwfu2oI17tWSLdBEosbY1gqFZDjVi6rbsHd+72vjCfQT4TVtYvGIta
vRSBMjvy3+O23QxghsHNiiQycIpgkXIHePQoVcphe1GCrcS+sI5JkJc2lgeGPrHI
8AmyKIG2tPurMfd5lemMI3bkp7n356HVzLBqMfwAoFBJZMX/BKbNss+SU21PGQYZ
BJqPOBAYOEGIn1YCkiPh/Bi05StLEbqjysXqNlZLDFCl1HNs7FjSA2Yq1JqoSBO/
OweJA+zX9cixooXuJNlRJX8lRmm2gxFkxxmJU/xjl9wJccMQeDOJ6J4SBOuQr9pS
eULIQm/285hNjSBdu7dg0/MRUtp5gJ43nrw4Jop9s6wOk8Zf/ayKE18RoB3/PZbp
qycAbHk1OsY2NQKW2kFqq6LSVCDUwyPDwxY7srBxzJj7VoSFQmjETxOFFzFHfHSB
h6qTbMbDSfYOawCEmF2YfNQLMJzERHbBA0H0AM09gMvFPYijVzg6rovRWzCNRQEd
+Wh/UL8k8DQbPjZIgFhKkT8l0SOafhABpoXXLgzUg+N+g6HiiaiZxkoKd1ldpu7O
5RPhqBsga8RJnVxt72FMWR3Yp5JIMdDb+UdFhlSCM1Jd00GnKUNn8NhjQUvkcT36
EuUj3O3h0T4yMJyW/I3j6P61GHCdUWyZ3Vq6INoV4jkj1umZd1bm6/DQqYLJvo+Y
1rvp+JKmTEocWWfrl9ldKmQxS1cjoTZMi0qqn9oTldZY5MoBF85bqoy+vi3sq8Kv
bad5CuEqs7cU6e2T13vELnOaGe6EV5dERMjdkXhdIWauIwKYf1zpTxNpWuVCZTkz
w3CrOMTG8CsnHgV3881PDC0IOrOlvoMhxehXYbYZ/3xMNLm070aT9y7Gz4YH9Nej
ZYBbHfjKgfw9jlsL67KS1BZRapW/XHiLsC+wm3e85Rrd8b6mPdDNA0H3HLKgZ2V6
92tazf9afIcv0HFgLuqJXWe88tVcpQAvs0m9mRDikvivIvEPbfl7xshSu9s6SUZg
3q/bmVrACUhAbYLy+JF09fON0/bNAfZEBCUuuQnnBlPy6VT/E9dMwkIOFC1qdlO9
Tx4J+ZtqeO1dX1QQ0t7qP4xqDrMQiSX4n5Lv64meq05jfb+f6w6MUwyYd/NLE3GF
nxDkkxi7XMtWPF1u2nvBNmFo43HjRwJcCm0qmpPxeGKRP9IHEaL2zzlkgMcj5lG4
kCzmesZNHI0719j0FddyUBQNIXRhWLF8S6SvzqkYfYo6V4MytEb9aKQpZAYCN1wJ
G7NqhPJczQkxqWMBRvNEs9aTpkHLPBapFMYR/0Q/A+Zkt48QtltBgZuqHIfnqKwF
3RKmvDvdKMIm2FqWopqgejRAvaZi0ypWJvfvu56Scnc+gIwcn4RFgNUeqsG1CDxc
g12/i71FceBHvBn5nx+wwk6ZEn6qvGqO7kFfAYNIaZhmA8bvFdTDGt61ccTR7T6i
ud1HFdvvFxgeWgsDa2eTFPF4NKko8LpNhKAMm+Y38pHuim87IptqCk7t1SlPA9d7
29rre5hvK4DtgqOzSAQ/c9wo8jQN1kbYjmUZ08+dLqTAmKfcrm7NBiwd/UrVHl9+
X3d6RhVFYuAxPvz+abgirMVQ/wp8fQm38bsjKX349oq1ZkchPtuD2539Jm50NSZp
7BzeZg7tkXkr3yVevgZLsY/+UhHkjk3xWca7c02QDaR9OkPfrWj3Esc4gLgt8YWh
Oo3/SlwKU2yx/OkK33PfOsUtNHtmPj5nE6qZzdmz0crGclzO5RuGgSDEx5CaC6hY
9872SWKmIwTJk5v4P9Xn/GaFSoXfYuj/Uj5msZIcTl9Se9u5/S2Cejq7jTvIO4je
f+Zukwal9hA7Uy1s0QWbkhlfCQ9NgZiyqwk3XZ/9MoD6lBbcxC1dql2lFVYhZcGR
5cD+CQnwSWQ0WidBQ1b0ad20tixi46eLyhTq/sCoZrMfgTSrgYlwrAT3SRHfGFLC
XfkzxufYc1wWOeKZTJDb1MA/kASjq50o3Uu0Zi8ezeuzuv07EHXXeAQ8iWTws54Y
NCi4qgNlQ0xqa5LnjEB40P/ark8ULbe8HwYnDvoOonM+p0kOT711tQbdjv6bbZfr
RCttDhP0BXCcuRiAMtGU2iTtmlg0uVYO+NLWfy6wJyANI+XLqhsLmOz/KWEO/HWx
JrMf3PFpXjmTPkhRYjlEFvVlauneCj0caoP/mf7Ptr72TAb0EsFeamLJDBtUgTdv
kIqAgtwaSfgM6kSdX2MJRZvWpNMMoTyGMITPlGCfQBNx9pazuc2fBdapz5QjmVIh
nEfekh3NkPjdYGQZa+6CvHGASpfIwuGvSoasW9gAKryyLzjHebVpKxqX+lOx3GUz
RthfM6dTmMSxfNge4Cuu7fZ2dgs7ggbBeWogMJWkMfuSUA6Py3iKPFOC0zcEi+By
OS5nwq1T3B+SJiOSgZy0cYqbM6fsEQ37TAM5QEDD9ex+OwDZUuoHVMgnyL52nHa7
0eQi4PwiQ00cvdO+miCVXIAjVqNbT1f+pCXjnpv0owa9Lo74SRakCVvpdA9mLZmq
hUDdU5vaN1C+e8kYvjxvsGp7QbpP3b8Oy3o1gzv7nVEw2SWDsL5sn5vhaSX25NHh
2E2ZPKy4A1lO7iFiMF1FzrBu3p5QwzMxJyzyQpJ1fg0s8ONv5gol1CwA4Tnkl5Cx
RNVZ1rjg5/UNce2FvOUgQrrmkLWNTHeoPWmk2WGmcsdwphVrv0GzUdfOvJjR1z1I
3ZBBlKkQPA2sVkKmNjkxaXX8uwENYeNtxB3YMzN7kYhC91xd2II7QupKbwOJgyS6
BdnYMSfgEWlMcEjKsb10IwcoPnSsIJmp4fbb0N5DMsNYMNqpIqr5KNOGmOqW5Zea
3t3RNO748zXS00vxDznY9ytq32bx22fxmqrXfPz2E4iQ0E9WNrjbhy5HOnjRISJ2
4ha2CRtYAG3TXT1ZFBIedoh0p9eaSjwHDjH1sDAD/BFugn+hlAPEtsfQFimQD+SE
iEZ/T4TIInk3ZslwUGDoysCSRGvzqd2MvZ4eng2GEo/G80jiL+vety5ibnNzvR3g
yCY7bDZ1ucKkl+fQIPPwIzTlnhVAxhjp2leXZnXUD/CdH3DandgtB4+i+89C+L4t
RMsirvfX4thfjbubBAvT27sjMWf3pzyWLLXEXQFj9hetGx65wywmonP2gBvYqSt8
qnRr7hqvSD6wuM3KDBtHrYAU85o+NIqwgbtnYai531u42ip3qc4UzL168sy43gO9
ZILAW8bcOavCSBFJDPe6WliH35+W94/ZUes8ZfvSsiOHPNkXM3go9oBVROwNKokN
4ATAPCLHhDuvYhzis5Osc+yHjbAzwwoH6b+2kCgHEoH34IqCNfPU1xrbNzj8vzeO
ub0do+j7nEVWzLNJII9kq7oYfR6zwrCC5y9ku+WQbFdzU8VYKERw5SOZ01HyUpOR
vn8QqbC9yO6PiBpLtVGGWsJaczNRRkAwUrkwLrripQKvTCNMJ85Thx75o8DZIIJr
qbF2hoqzkfpCq27aMUZXvXFXgGjqt7AiVqcou8jJKEBT72aCfLWq//0CqNpWTnpo
Kyz5sSGlZiSSRmpNRmrpUY4daMY/HP8mNzTJGdN5YLrruAlgULkrA5xtC+IpxYUq
MM2hgUWMcuLmMbf/GawPVTmLoZmMuufwDpfXWfNT5pTW3CiM8dJ+rnKVRhb5EW7+
NDRPfOgaV88D45NIe0dCJsVrOq3yD9SHJ0FNLnzcBl2nYNkI40QNDZD3YofzN4JH
GaPa8AZgQXSsBbulZv6DFE9f31ojGSINiVP6SzKoBRkpWefu4juUCy4TX/aXzjcH
H4O+MVyJWPVRW6+b8QznGGEYFb4Yzq5y5tuU53FzFOhaulp6i1o4OI0r51QKj6Yl
LsaIBAMev6emD5haeobZNMLerb2KdCiCOaZZ0P0GncibWnDMoRdD5q0AQfpR2jVb
0JIFhI3tIA2lsfvOCbhhURUS4mnxgoVpL1AyQZ6Xny4u+BE0T5B5EaJG5mFoUMJp
arEA0VRbG19Pq6GzZMQQKSPTOMyFt5Q2WyLJXvycxev1WIhyHsYHP2iOVJ2t5nBs
oa2eepnyXgHRfNl1TCsIWYL24USWQkxnD9mrws1vwfe/OBei3eTdnr7KK2Mc6WZy
ykVj4N5TkiIvg42NgsW8mv6+Ch8U/1tomzfubtw+J6vU6F7RbEycna+4JIebjwaW
0y2JFdZI5kkPxGHvsl8/tdFgaNAddqC6ilXfCJvlTbjJJvWvwOS8BdANrGxRebsS
IvY7FtIzTEssfJfOBEbtyaadOL4CUXZVeJeKyzDIjE+INshrWrcYVi4qIBfvIGvd
OLrHCmLA6JX/3GmI7AH//79E5WgQaoj94pswNjA1cpF9XMZ3VFcM2l9rFoB/D2Vo
F1e58S1pTpiZJDjnGD1ZoB97ZowDkdzIYIuZqny7ap9Wq28TiY0fPf/WbL2KwaQJ
jjOhQ7825ynfSg2TRwTe/Ak08WWsMNywLk7owcNIFp0f110fuiJhLmCqhpKcVTUw
xmHhZYxpbTYO/cONb6YzCmwTvpq6jNSjkuksIShjHihDBidBzum5vwpREECrB5y0
d68EZ4xFywFQhySp5RupRnt0WHpqNWoAA9UoC+0hL5K826IQSaS6XQWWn5hNTOWd
3xaK2ltCvV8ZbrkOXTMh5MIJdcOWoNOL6QmFtzIL+BSyFwZCAblcllPk1K7vKIx6
cPcbBnY6BDB/A2sO8eiX/Piak1sFLSvMdBzSEaxkhxhOMgzz5EOqotH0cx/YceFr
fP30ohDbozhPNrgIDdqTcJgHqnzK3Hcma8eS+BEdSrWSXLHsnD3xX4Uz4JgrVtNG
j20r5Fl8eZcIGWtvwgZTH/oLK/bFI+s+5XO6vrPesBhr5ug1cptzJ6W9eAJqOER3
cfyrnMvzKAIUTqJ4rbJKZmSv0KPnuU0fdj285vOGv6iNcYn10E0NJPkDR/wlaDUQ
EORa9Kwzk4HsdMehvj5ttd7moYwntcTYwnJStzcK7423ZUrZcQnvbv20WcSRRvtA
8aSpSI6j/9MfBnDBcKP6+6m57adgQJTpJ7ZTqfobiVUfcLB6Abg7xSUp8bLSuDDx
3tF3H9xZfY7u4kHfMtqyFOw6UuJRKWBwNQ5e3+ZExI3TpFm8+9XajBTvZja46b38
MiqLYMKmF4OwotMP8w07b921ugeBqqvSUDtOZquX0TVBEVIAxZZvxavk/CaBZ0gs
cTYoAZwDLsqySa532ENwCPbnuCoTIRz5Hvymim+bdMGC+tsxSeCkPfkYFe1Bpl2X
dRX9Eamus8JXZlbuArXkuj1c0oJlFVgCN1aRdXKWg7eGbXKNKlP3mPP9R8unL/HV
FXdugxCA2pRAS/+LmeGUuw9Nv5awFZZpQZluD1UCx0fa4wlaK6RbXlWr9JTHqsDJ
LgmWXKbPT13rx61/BofClqbCIFYI/gWv4C8XyQF/G8U+M0mra/7ETxa2iH64cYqA
Ak37CVkpR3Q8TzCbtx/tTZddyOUQUOtIvNSHVFYM/nWyH+q0kmRnpGjgVooIDJ7s
QPz1sxAVNJNKifOiINBl25jPxnKGzFKZHl7sCtpJamCEdrIs0PAt+C6YliPmIaS7
v9a6j5RoR/K7K289Mw9s6WqNDRfb/MpFDKSsSLm8meEEwAipDhRlJhpWHH+yzjhF
StByNLlc4T49OUyip5R10SRBbMoa7IdcMKWG9zFkqb80ZBftt/XaIglSGT/xmaMr
lZFuH8Whz93Vpuav4HGj4rJUZ2kj7vHg9J0yAXvDpiZpUmTPRNMOh88GzKR7cNqR
ADlslb78GfZdCz5oVCCeEwg2ME+ATGw030H8OjvBKEr1B5g6WGRHeW5HGOULE2Jq
7w+lOpxHTvw/kS9+MvhlWvAIR/D53It6RCAmuKxUddoVjdBHDYM05PR4VrFvOBCx
1QHpqHAbjcCxApXKH1ELJGWBE2Y2wfGGbk3kc+DkGcsz/tzpYtBW0p85wxs+5CQN
0+5D/onx+71GdqOSCA4H1lDmblRcuH87mwwmzEuIiyvLvKo3L8J67Cd9bqZYHLWf
0wm/cKYUJ0FU4WMsEY3t5vb+KQvaW7eCytgptOVVEIBOrZazRxz1A4T/+8vpDsOS
SaxU/ZJTh+vu1hqCwKQ3GDCNMzlgNxSaumCFHg1fCSlEET625v51iWg5iHbIWatt
Ubhu2zFDRMJEwf7v2O5vR1Z+QVwrNosMx7tY1TpjM0oDDPztgC1oWiOu4EnXjv60
VMNUtGHDpQahohTHE0JwBzX2RHJu6ujQVlsXbpUyqxnw/uRvZ6yN2xyRSIyJwRlx
cIwUmux+Gp02ghDJy801l5sQqNvqxv2S+GKFLcSa7BvB2M7dUjeuoHVmEw3zfj05
KQYw/uf+pRCOl0RxxT6UYnOMJ0wB3MExAn4Jz2n/Y+jQaYL3wp3LZK5IYL7OxiUg
PkihiBe/qDvesgYMEtQT07rn32pcBgOkyH8fBlEMYw3tn/9rAFP6K6PxZp7rPjMN
QG5FF0/noaUV4vCyX9EXYhA8Md+gnupBF1+xAddGNaVcsNaGBc9gY4F8tVAxE9z/
J4y4Z9uY04OjNPeqqXT8iiSIEFR6WboMZfaHWkzLpH/bgRzkodcW4jzn9RWYvhTK
iO2CI99CL6buAsxiY21/ixUdR/1h7PLHWurW/vonPtagVjHP0T7ZARnd31biDMnS
F/gnThc7Op5QjyTuq8wOrdqxTOwsk1l6Y0RxG1Nhb6vUijvtKRIaIl5DQvjWR2zK
M3y8DZIqCkSCAjdTGUc0JZeFC2qOl5AEQzWlVKPTI2Z93HtS4X0eXvelcImIleAt
T/LJROhEqdflouAtFlg/Bag1yyAHcnZTvzLK3hEjzNZSWfI/0wdyOtVG1WM4gBRI
o6MFGXUnOqRwn0l06uN9W157sXCAgf+iIbpKtbmdREXGZIkIQTwyNDwXDY/qLeR+
AYMJ4G+H70YQ/VQp5odDEXDEPnAmPjl6LXepVTCgoz3jgTCQyGjGe2Sa48ukvrt0
uUqStUmHFLm9F2KyX2b5q3vF0Q0bF6xkD8Us6gg4cklVeTXxsrb0kJzqjshkf0v5
I66luvM07GaOMbAdEMSB2q78Wu2wz4q9ltf5a5pqlwCGqZ6DcgntOABsrF5NNAo8
vejPdAfl4ZP149dPw2UwSoqwRyps18YcKRoDxSeUk81+vYMNKxn/z5RHDxgElZDZ
Bk2f+wwBwc/D9c7G4mLN7DOuFY9FgCUBAdszRoZOwKRXXOTxN//0UPmD/sDlKVbA
TnK5krYG0CzgKgAcApFia7CPrTAq9XY/yRG7zOI+fIipjfZEcJ9suRpF+da5JczM
SD85tsadJU/VaZFPKMMYiWgAgP76eGtXkPPVOy7na6ITosuyHesbP/Ljp7cu0Gr9
n6ti9kCdBQHw4M/lSa9Qo+Um2PJzI+JbXVkHgdBnF4eEYdHyM867o0NiNcIboBQW
iVcZA0laLMwopj2dB0TEOhF+TT55XSheMBQ/kVhLs0rKyGVCij+Jh0fGpqWvxUSS
XILdEBkiCZ7n9ZYihfaL9GkiVoA9NBRZ1xVBlM+eoA86a6hzoZgItjH8g8ZfrcdY
rvZwFzjfgadzhIS57gmuBmiCOB8aSfRpemlulCPI+xbtIRNROzStqgAgFbVI1yQk
al6h2PhUfSLuNgXSk6LxatHDK8FryEklXpnnzL+70Vd/grpoZ8N9bh2MD2YCtDPo
xdCvQ/Sbi69lY51gk9eEq7z5Tw3R+rq5xW8tNtIzQ0lMg3E8C9O/fI9I3dAataWW
NjHKVyYQaZ/iGDLzLCoFX4QU2YZguRts+RtlwpxPpAfMctdKkFOq0I8MEM/GcdSl
YCsvG7kH/faY/1PBW1mXKjfI1lM8coXrUGFA9vYH4Iq6Uttg95oi4jHPwwJ2ZgBp
9OwALf9BHcfeAJHVlTXwKlkFY/eXYD7DGzYyDVXj7vSvLIUSNWJrZkLtmjh36LPf
d/1aWE514wrlWeeqYzwda5NYy3keidv8Cve/tFPmDhSwYceszkmCPJZf/X7YG2oS
iV/kMdo7f2fgPtwJ4nEgl8wOnDJjt5AY0Kg03RVubCoVHThsjtrk0kzMJfkrBWmO
JlUfx58DDAeMQNxsoMB9PSKhBsrbkgT7MGgLoK+NPbWQyh1n4aCor/ocrr16ShnF
8m/FXLAjk2sddQ5NqwaK5W22YF/mgYneJ8jpLhjzKf2h65CMmE1blziTrPG0KtVX
ENBiHeSuSETvuhnZa+v8bPIjnSJcc0vSBSwbYBaCf/qmAxhV/G7amfnI1i3oJZaq
h8usWlswOuoBZWsa+NAauNUpusnS/kVlyz6Q8pOs+xCSHDqoGou7MsAG7Uy5rO+j
UsMq/2ndpO6DX+9F4+9OdWw/du6voDUO++hS7VeJpOMQ9dySS2Ltw7HUc5o0YFVL
mXSH1wSr7tmnBq/dgY/RWUPVYfdFyvYQ7/X6XtXs0Hy4pn/esEana9fYKqsjMEL5
8QXd6r128prKVOscuXnxlaghUZSVCBO5tIa6AyJrlkugVUwwFduT/olA8NNKnWQP
Suq8OpQ85NEppaYO69DoglAJXfqqvMqDc4I9zgWfZSsYLJl8GLlRFonNwnHvzGgi
plUalWbqssz0KWrnPbM3cmtxzeOT7M2opSLF+DhH3e8V/Tmbyj1LxUwyJI0i7AFM
89W8dqaxR0hJEN8jORAv9Y0MCJkwedCr3SnzgAjRKh2yBsAkRWq76wWxwiTU1OXf
xYAGTG49W6MSHMwiCVRQPy78zWkdPLCCxHllswc4de8GV8HdAiLrd1Hyw1KbW6rT
yCSfQHqLBzgaAVMsVXZ5K1YOAs41wnsCk0QDy7geVajo+A8iFgm2qkR2uW1mp05X
bWp/g8Zz4z7Gs4BFZmngkUlaenZrSuZadoB8VEq5jv/7Vuerhla+Hk1mhX8Vjv91
aMAp4NUOpNG5rgsXCFkh4kIFSzXKmRQ5d5v+m6xSXhethNTyufft2oykND+CQSjw
DwxCON0AKtLBzEFJjbW1F2EcB2jOiTfleqMYpwfH3+BLzsTC7IWOTQ22T2Z3Jc4J
4cwbLl1K4vQrRklqo/2vbnwxYtGsw+OF6VnZzrjti0Of8XlCTboU8KAoEFp+/c3J
1Pindp6bERMT0Bc72ssH/UeMg4ThNe3hl2hoZY3pkdwmXpbnomP/Rev7zneG0kRT
ilEgEGzb2p7yBvlkbt1Ogp/kbBW8FTz55L2p66dZcWDIRWvOsZHvX6e437q/Anaz
Yoa8/pQq1s0vgtoWh/vhKmiSffnpOupO6v8jDUnbJEhfJFU6ELoOetGdMiNP765/
LTkxoGTwQSnIOXROsBS4F8mOUg0aL7/ztXpZD7WOJBfFY88rqqDfZOgo99hh/J19
WM/P5BPg7xpt4WD1iuiij/mBpK7Q8GH0vsdDKLTTgEJ/dk8/lPK3MC6vjoMbLLbt
gBXlfOZPEum+el9BhH+2wfYtC5tpPxcfalAJmj9RGoMilp+efuFnxHHbXywXxgCR
WNq8LekWXXRsU5RuWXEICQWORFza6Plw52SlOEbThAVxrB0mB023CNgy/5fRbcPK
gG/pE7TA2BsSQRvpwbakH5uwkK8Xq942aCAM6DQk3jQiCWJNErw6BMpwOGLSVmIN
3Bu+2pffLKhw8od5Kx5ouW1VL2VHfOttMEXbB2FRp8DzDv7wIKFtRoNFQzDv5AlM
vcUyZkk+rVuPNR5SWCeqa+rWCaJx9nofTPyP3y5QQF9KpnropB1XIUy1IRlruuP+
oGO0c05Pg9tNdVXKYFWgGesaodnvLGwWLCCDMml+arqnOVKBorM3gITltL68kNAY
Argo/RLVeiU9sh1wTFoXI/x+fXr+cmHSbkhlW6F/TPPo67upm5WQYXLmu/f6Nhyd
TuTvb1DREK1qC2S1bb5BFV29fIPlBEeL6EF7iYbqlKujsxTYoCUbcng7Sdo2HBdc
OlW4rMr8zX5GySngQZheQ6f8K3Nfyn0aOZC5aB85j1G+U/kK4Los7ZVxKJBstE7j
ZeN4FqZptB7akZQECF70+GWVhVzAFJ+iRNT9XXwrLwtG7nJE5eeEFoZDsP5RD47X
Jy000YcmSJWm9FOw8k8oUjeUyDtS271+wc1WfBM2eLRc3UYbScL+bOsDCMMQNqL7
vGNO9A0UEkssLv3+57aucg4cDbB6f01msMy5pvrVkxrU6CYlugIxHOR0mRcA3JSU
p37evq5Q8es75tyjPkFxmtCRSLnhPDx2VMJiTKLhsF7Io5GHjDM5jvaeeah1NTLs
e25E40LKF3tEJ5NFGnLEtF8INIhOV9mAu9Lk9UMIccVttp36aJttBDhsxQS2DAP9
DLj6jdMeDH7XMYJqFSsckl/qLJcF0yDHIBPEEBuCvZtcpWLbrQg26TEv5ZfSLPCf
2rcF2G/4z6GGPsxzWzJ9c6DM87eIALc0CONQl2OEp0NZcYm81uxaUepTkzCxOhCB
0+mEM4l51sP6f2r8ZPdBwcMKSrFwfJ3cO7WnJyaLyiBJ9tNdfyl+K0aMcN+BZ4Qh
Y72ytMJ6JE4s1lQq2ynz+XA4ipqsr5xtX+Eg8vGrJ4gh0Zir4F1sWhwPkehFq10P
hYFy955uvg7/xiPPb4O5b6SD8sn95q+gpvwiitJjy+NpAHMy+mjoMxDZqTK5SeLk
oosF2BoZVQCBm/EkHketVeDfWCYXClvH5V6hcqOboY/U3iDUkKOfrnvqDOINIIqO
rfvX4oi4B5lzAI1fZuQ948IWjrTV8/XuBWApHhSqvxJFxo/IIXGR5aR6nNEdf+M4
+NhcaYLrmzFT1nF5PRLSQIdiMEukrVCsDs5xIT+L/7TbKCy5I682YYeQDqFhrX0k
cLKLZ5dRB1y/UtwIuse5Sddxcco1R0yFrejBeLtZf52MfCA4MxA0RYnh2+gjDlGL
PlDDP48aHAEY8nyRozm0F65kT+es4fIm3s4OXNZMwrCU67IY3RumQGicPzX6XCZT
4lGINlFbwBkBh44eA3qX9Io/ADbsOCd7YI6Hqfe5knPjT/kSidiB/OoTOsy4nvAP
VThANBTgr8qbrIuu97pg7/rwYLrQJSyrXFZfHnUnLKJ482j3rgK/O4S385fWvL32
RiMnbHaPEuSkb832GAWDq52BuaPb16Kzic6Sk/M6bRhSO1CEj1cec4a0KfMUWhLF
ep0NxSW8ydAi+RT94wrj2sMgi/mnCS90xZpI7kGDfT+Q7B7ZNU15F7TZt4IvIhrR
1tPuw9o4Kn+wlQHQl4u9zKL9iSa4pOSATLsJgTb9sRtFFuiqLOqA6KPk0jVsja/Y
ooOOFyw8efcceefiSMIQCc7wUPFYVEriFfNDUEFYL8ojYAO4M2OLlff/aJhj5+1Z
kWKOqNtJmMB7KJ8471BEDkyJaWkW5pL8DB4p7VVm+tFJaKiPQEg2p1ti9sBjvlXN
cqSm5ACvbdePHOP+f7rll5SiGGoFwKJnTWTibRW7aZkCgu877jz7ybrW28aiM36E
aZVEnw/4yuGVJxxhsI8CzcNmWAvznhaifEAiKOitRFw4w4Gc3HFYPvgDq4RvYsWR
eXW4th3T7DP3MzExGwOrVNDVV4mTRE0YTjdgPUJ2JWiqmx8gwlA11HS20lzdeOf5
pn6lBKfb+7gP1dvzLtHlP8HKgEKNuyIHCeMWyHAQYjOwDaloA4KAvdR8B2mtrGEM
E3aK0td2owoZartKGSkJAWImrcKxhDVtmerEBHAtn1rsNve5T7cutqg8B5WagJkD
hYW7/+isV/jUzpKWnmbc18OGOwCvRGx/CmvK25MdKnYVG1yKPlpGEr0KfrB9CYKV
jy7swH3k1NfVX/NYC7tbkTPGwUHDrtijwrKOSnNdr0h5rCmoA28fJDeIkkCRgCHM
x3tWQFJphYBi5v7VGWv8Dgjg3S7qFQRMTiMT7FgYYgb6KmNMowFi4upltBMXJxPB
oSRXGhJG3BadSaNOV6berqHVebfw6Km1onaVXFwbII12F4qDcPyE3bOuhDj2Q59h
vyi5iGm+Yi6tLTXx93jNreaJRTkRtIXe2L4880Ge9Lkvp/v1YUerfbvrJCRDea5Y
eHzCs8nhJnMn8RdTsfOc+UoVu3S4GgBwKaXWbNZvjB6YeehNedLGbmUsIOOGayOt
s0/wnxy8JsvXseihDCYjoBR4Hbg4F96SVzho0XXJH+2/yhb7sONspcMfkOZxUyoF
hz+pJwjfDWog18NBp8fCfF3xJeTpNvc9Exls/x1L2iYNHuZNCUFXUP63R3Phm7qg
iapJB1FA8OsQJuXJbdY0FRL58E9ZRQE53g/VvyztOjia2lH4Wpsto2+7Lh6Jxsxp
BhKLJMZ+Nm4En85v20v5w/ea37IR2b42/sjMrfHH1tmkb/r7qaBgZXfysZ2fBJVX
yzxQDdxgw8D0wYIvhzudxogX6M8zaqVh4A4HEtGfu4a7lLmHknNCs9UycGBjp4K2
935De4kwBZwCs0N/sYbHvE3EQk3jHx6NZgqgqefFj7wFC7HSEWb37y6Loa06IwRO
/RD/F7B0RbZ8ykI50ae2uGcKbdgJTZtCg/rUaYyjZ3lvzztrRHNFlMTYainLxkEi
JpEDhpRG+8NfuSWgCRSzQKAExnjpN07TcRjjsW74UVfMRvdK6vJ2MEuA1dv5R0yK
qHUB6Cs8Ff9f0g9ZOPSsr4BIy3DfRwyxTjO5Tu0KR9TSO0xwWiWq6VidU11vEYRo
2PGYJFDCVYmfGDxe82vIoEr7JsxINCRyPF/Uc6NmZ3p1hrITDuGc+2eH/WpO1FUW
poaR/WIQ33CNVaRzeWDAvRW6lcDLYwUeiDyRFFWzSbwftsC/JQl31gdfFSFVcWzP
Av0GXPimVzcw6098xyq7RIUO+fuBSy8jlRWYcyh1ezzSJxUEUaE601Wa0802QvkC
0j3E7SFCDCw9GrkwNK2+j9t0UtNwSexoQ+At0h20LE1//qaA/SD8aYz+SSCqbuNK
chEy81CJJRUhEGUqzXmG2ITEChgVm9NgzbRRg/cOiROXF0Fv1EWzZXwCIrY/w6i1
RyORdVEuOWlgcWAaZMuF/R7QlbFyeKxG7+r3or1FuB+Ju+rWH/s/8iCdzr4GU025
k7uja0pm2LA5sHsYond7PJugQk4ho7RHm51uUS4JDnUgvNEOH/1FtF8ha7j8SEvc
5BAzYHhbj3dr4XfqBu60neRd9dgk67eVxiKFbbKDCyFXpet2M9U4jhYnn3aUIW3A
l5gLdZ335qkCRghsUjNZoEU+CrzottTL4sU/HbAJVy1naZFyRdk753WXrb9Df3Ip
BEL8rvruDoMsDhTQ4we8oJ7UamIjRM8stksuH7v+yJ5G+jDmcfN6qjdqwv9klWcP
lzlSoAdN3FIfV51oQEJ92hx+J/AQj17sKwNObfih1EZ2JNcx+TaTYhkJmfxIoJV/
psaELPdFQUbEbZQODWdUWP6pd/QE/ISQ53xDjq7Qa57y6+16huR4J/JDiGQFpULC
liyMl9gUnoqXhwSA5hG/ZLzNkEDSo2AF9Dz640DldBua8+w0wOtMkyV7iRIQWHUF
polKbkxn1n1ghWN/iQzpUqoW3IVZhq3FqETNx20YS3LQs2/v8OaoxGJ/VGmsRPn2
uYT4lpt/MwCFvBjFENfA5nEQrqocbVi7Kmg2PgeN3HQBF/QjqX4bYX67XDlP0LZJ
x6fw2FK1iFZeaQf86K3sH/Nv7tJeShnK82cXojot3zquL4nUAbdh95TQTP3GqU85
xP8CYHvwAGNlE/ycWGonnrmdmOfasPHfiPVtiseCB136C4tv5AK/VCfuwhc5Qpzl
4971hMKtkGTzQsiesKb4yRFMlLzGBqgCU4wIKqUWz0JBOpIxMlqvUp1uZlA6MS2F
4mJlHEmjyAaiRfEYbe1gFUyRN5FeZJ5fG5Auv5sJXUddtGT0PjvlKTKPpbcBzRfN
1bqJZNpvtI5G2bdAuWG3aEsgkKP9wPdrO4tFy44fzkicpoMjGb7dehlU12Jvcu4G
/0Ua75CLKqGfq6Qh3lu85sSYyMCT239tkrodN/PEAwLgrjgvhv28yC/5bwT8frU3
/8zto6E+5IQLQih8TwRylNo9g5b41U4aKb+PIf22y7sy937rHLl6jgQo4Lx5+G2H
6HcGVbhMY1TaE69zP2nKlnwcXlOLcQNzC2e+vVJs9Rf4GH64OBqUb1NbfcCMVk+4
HzFV88a/DLuSKWnRZsYcuhPuKxYKxPLdgCWBbcdDGuywHRo0P7RXZTetTKw+bI0P
/tPo3Cm1Wrj+iMI1clm/vd/21Doz2lqRdbbPSbR7JAAVowXlboA2jkrv10dZZtIh
2O8pYmLSFPn4vgvemivwU0bkpp9TTIl2aZg5PanjPCMp0B3F4Yo4sCbrpNZKxAwT
2HWhpyEWxhXD/nSP0Jt5SWhdl6wJkTuBu0KuxrsuZ0jWbWcu7QMO8xPKL/fEPnz1
lO7l/hpvBV2dvln6h+OKexXF5pBEGpAI4i4KAyCztd/xWGGliX4sFTlxQLkbmZ3a
kArw79cRLe6rmv5S6afSjZiHl1j3QtjFFt11yPwxrL2HbK9HZAGmLRtGzDn9d42q
1QiIh/1GWpPXX9tsPki+V/FRjhXpNM9UKuaoCqo0yQhOQPx9Uw0L/zEfRIbblqMf
ZprDbAnpTbEapp+egHa2o0Qt5q3Xq+oHGOWPW22GD+CUahMt1rFgy9sLeVT1FBFo
otNWMscwd7ngCkzXYDYEu/ZzcPhLA6ZgM5tyXYJZ97zyX7yKu0bILnnNQ27VaXHE
r+7mwM/5kJGvXHPW607X0XyS9jlWrtfttzaurwJQ+JbMDpoVN3DVyVg3ChNTIX9L
XVbcoKXn2RQ45fONCizssmuuC62W6alaTMo1ibpe8Kd0MHkCqVmF2yJcvbzmcacy
Gm8SDDkTK8cWIJ9nPyrNlQfuX2jBkiq5OUqLfaY0Mwwxx1cGTdladC9YgFHlS8QI
5s263lMrDjYajcx6dzx+yoSWah1ep7CuFPIgC+8uAPFxfEmNW6xyMzFUqkUlGFkV
z2PWoUTsUdzvSvC3Il1RdQRdeANg3Iiv4YOm9Nii2lTL+RR31b3aJkOoIcxuuYyp
+1WnF4hpdzWGwahAgn6TRkcHB6WJopXtJhx6H3HYveCTgvWr7fSM0dFMMuJ56jAl
y0S0PTlBP+i7XhEc24UqP9zL4e07YzS5gVwJ+GhcFlFHaG4JHWmJuZ5QNGUUUUR/
fBFAGpkSvqCdBaGp7t+VUasP46+kak3LCt89Yt471fjzact5zdolAnXy7Lei4Tk4
DoIKeZbpRCzrlFgoLvInBz3aZFULUc8y+frZiLFNC+Zdo219LxG8nAmQhPm+J+Dn
o9wpT9MW2MeoDlWyo2iymeVF73+OrX2J5R6UlBkNtBlMxC2QHluFrb7eu6X61h7M
J/9uwkqsaEamAoWkDPSky2SMYUS2dxL1M81ibBneFZ1JGbjAEr2B5NHCz85hGBKo
muct3jt0XnfdssAux5xJkc8dCRUlsOeM44wuMXzf25MGzq77ElumW2JyK+f3jImL
XmFqw6z1itIyM1i2FpXcgFk9Ggq7wNE7Geu5qQPpbRKPex0IomAt+t6DMOW1G6U0
grA8EfYY4jE9z4ZySn+E80XnNyNFXxs39hsFzxJBpwZJVnG3I+phJ710kTPyEKfv
/Nz7V5xCwBLTSWsv+L0+85eM9h2AtRgQ9gWXIVFrj7gIkbZLBdfAWAWCWz+8K6HG
dSeIBLSoqOOHauOc9Lu9gKiw/pGLxJ5EuLuWmP8x8+NY5GBCP7BpauoRgRQmZBw/
SzjBQsBQlNJGmpq5TBtzpaLdjF+tqhB6Zb+gIXOGXRzyQIoVjkehnBBxRAkoPVya
a4htQcsOsLb8U9pe0/8Whnu0h9/waj/ciZ3AAhI+Pvj5scQAT1CQoiWM6qvL/bbX
9eZ9J2QbFJP1Yt+BPo7+rCx/o5T3TCOLaPsDQ9mTc+wwo5mXoa1Jjj10A00Agu69
oTjf3/Y4cUp12VRj5FP4Koca6fNfVGClvCNPgHRVfHjMd/3G2ARjcMvEWy2alVXD
iEOIdQMk9+a7T8BcOIzGYBDr39fIx9SFIRQsvlYpjoD9zFaGi0hQ1+TzYiZIJg/q
BWBVoFoGY/JCxCF1CYXoVh0s5oksj80lkZaKvCEcmJrHZXWoc1DFycG93UCWEGGb
+xNxTbvDkXaoc4VFBFDzGbScPbl6QI+DM7id7skOQo+atg9PjygMzR5E96Uwk0RD
EFt+0om8XBc4x2blpaMA5oFlBzK+wpOfmbS/WWS/GaiUBAR9eA5oTcwgNx6fiBkm
fNs+5ealOUHxQfMGJoxUMRfZNgZsFdDkQbbklYUoUWnR/RtluKZZ4dsUwVcr8Xih
8TXSq/mzyRGJ6dgYxBaOY3yjilzBdKEdACFl/Py6BHeJFkPCUksW6qiZsenan3O/
B6gDfPWQcoleceZ+3JySKAmJKX+bBf7+3tT8LrLNwgPaLpksSJ6bO78Zp2gTaiEU
wZ8VBC18Zpdhr79M6o7OS2ZjUcxmONUJyAenOAZdN2S4Of7IQFyJFYnudatn279q
WrRWsy84kl8eOUGUvP/8c1tSDVF4lU3fejCOPsN7ENInyBILe1TBGO2TDZZ6f23T
x+pI3CrjC/28Ipj9Vbzvg8oJeTcI1q6Ng2U8cAlVWyLhMBB90dUb9aSC0RG35K5X
A2b/WYEcJSlPNVnPvMU+4ymOvBM8iijF2zPk13CYLU2jJBESArj0Ax4i1njHF8ad
z/owLUdF0mjI+5epROXwTdR5xEE+RVt24XtR84EEtM5TQm3N/vv3IQ9ZyqE9guBP
+Ef8OqzyqGLBBBwVJdfjbLsoa8cKyH3KoAONNaCSucRTWbhC1qnl4dCWO71nYRCk
m5vKDNSiOUB+Q7PLV0zK2+t8HwXXlRAVtrjZz6zPIrbAThCfJaJAuh9/EcC07sv2
RCiHA7gdEOP91TYoxQ+eyAjuR72tSblSLZRR7KqY7Hu3VFFl505ZlvR976e2JRCz
VPotPQ4jQIFH1NeCC3ebarxVWx18GODA4+PTqGhGwSt7NBSRiF37wEi201kMNa7l
iWB4QuEpOuuJ8lhCe7DcgLfadRY1VlZLCssa/bsC9XA8WeSOxjHItabg6rccO+BI
yvsgUphwNSJbAD34GLsAHfiCIjI/uhF/z3yfVtA2kphnvW4gpu9m5RkvWKWEoz2C
wpQLffTExXnpQF7zkIdOzf/5faDyvLDWg/jzCIuul+Pfmuq7wYKx5NaOErFd43vG
8HoAOwLS7QaoNxEUsJreJlgBBHHWYDE/QcN7YIsft9LR1lAOUBgF120GQ70D/xyF
J3I+JHl9QpcpZD1xngkwn7kuv1M1JJGGy0AY8XvZ0PPNPjAHU51yryS1IHzqothO
RcPkU+K+4IFuwjq0OL2l/P0w960/3jV2IN4j94Ntr7hXLB2BA0VT/4uwVrDGqgWK
lri0RwA7f+jU/siXRSy0EB9zGRYDGKhy8omdEbmZVvOPuMsaDtGGbcrAR38Bdx6U
0CZgdNCXnGHJQn6X3om75rQwNLS4ZCLzivIXpLQf7sgmUpGJdFJSSKjGKbTrrZ42
v1EItMb9UVeaCHqFMmTO9V6Vw9fbT5i22D/9TKwa5UrvdctvwHmVrxz1wV0W18GC
i01QSjAEe1vhFiA3fAeNJZa/TWS+Eflex2QJBIOsR4xX27JUCubBuuI7qh94He1b
Du1N808DSg+/8P1m9k8KJuFuLoXnsvvtOzm5RH3wbK7m7aSSr5WDqVA3epMnGFNM
nqChBoNcrxKzXMINcLfIg+A3PVHwTZUm6vkdUyloioRdvtNWyWO08QYlfxK707ti
MBGM/vKiM9AOBnTjgKyodoLHpYankSkAUbcOLzD7GTOcCv0G+iwsatFe4kydUfx3
0p3Khb6jlS+/EpbWDWitRrc4oE8T2pR5c/eHYIJsiarbAlHgnmXifvJFZpv/WcF8
im0kg3icvV1dA+kNkCT3rf33pqIqd3WBe3omUy5jlyFACPB+5r1NuuH7+Q7U+0iK
RK9TLI6vhdqxGONFBFjYyAfJNAnfnyy8yJeFQtPuR4w1R+ef9CC6j8u9vmgaat0U
EbN68i842P4ejLZzNsOjub4W8hobkfbLf6FZCt0aJvvpCv5YKjiec5wA/YCsZE7e
uUtSzHa+yTI+TtJMri0T8IDTp31WEJyYhblAvSz8yKsjCFf74ksLyZ2S5uUk0n4s
RBt2dK5/Os2XvIHUlqsr35ljfsz4dSFXrBHkDX64JMSMHNrLqY2xgsx3rbCxICi3
GXFtCtIxXXTSjxp0lOyCVkgFUpQynr7Fs0Ep8dPJqyqtlU0HJgeu3NNLuTBLGPSV
5y8EW1tFz20U1HJ5Sn3lERiXhY9ZzyHOL3C/+eLrMp0A1G0upK4unbuyOP+bHquU
4+AEO2mEoBT2OnjiYrK9z2wHqPMRl8YxBkW5dXgayVw=
`protect end_protected