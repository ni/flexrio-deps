`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
YATj3kULTF7Ty4ORuRfFpnT6YIk4rUPRrM74bVTnc4GjdV8oSnW5PtQkMCLOi558
1V+/wvDfc3y0Z8//ksX8sZm3JZWtrxUppw8c14g9Y7owiwp+JumRtO1zuk5xFbe3
0MMnIxxoTKLhyRJtAxElG8sbx8N21OWDGiOk0Xyd5CqAmk9dcOIbxzMjW/wndBXi
maijUdqS+5KiRCM9+Gsp6k/iEAa2LnYTt4WtjkmDD1P5jZKsiMgFck8WOqLymplZ
ml3TTfn1UlLNm/+zD3SFGP0kABAiUT8NK2xBPQ5UzQ6sMFPd/np8iUZ5u4QLTWOZ
hTrU9OSX7lOvRUo8pJ9vPg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="BzW6NOo8eyBw+CxsNNo4wIDxODIsVe0ft0K5tGuSUZw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
DhjJh9S2BY18dG77XPz3hsiSQ73+w0XqfJhD+f+lIDHHVjOB7CfC8ieNRTexgzn1
5W+qoqOEwenoVQtit9u3XViXJSRJ0wfUC5a9axblRNyD2mUbyfH9+f59nWqGkVOh
ieHxkA/DPprM70F3APxk51m7/gNSLICSvbONgLGndWc=
`protect rights_digest_method = "sha256"
`protect end_toolblock="L7NTNW/5Dqy+2kJZXKczEa3js87UJ8H00YWI+92sDHA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 33072 )
`protect data_block
6eHODtGLmq6ccbB074dgNWpdzW45i5jL0Nzx5wwM+RA0eeOHXxEV143NNyQGmZjT
bzHAi/6AyRCB4X9z0c4MjyrZE8GF4crbMH4T59xFHqVrQ4zXCea5w0kG5yvHgpKo
2Lp2o1suKM6LQKudLJWun4FJ35TdGqzH1R52XzmLw5t+wji09xIDJHO+Mf7VSh1l
AExWi2h/QBtGp0qDr/RDl6n/cuH5bi+0D9znS8YkFcsmRACgu0WmWQu/WvO79M0p
OghfxwzrWZybbtcFPUYLKTcGZH3qYl77++gWPLbA4DhdAPxbGJHfO5ma1JDBS96E
lbcZsLA7zLvMlQJIwH3ozsASILO6y4DyEcknWaKU2mqeFLL5i2fddHasKdw7lh94
AAQUbkxzgvdq7EZ5+AsM1InbNYOf7E0qN+tpeaGhpFjSHyQU62pml4jr9EUBqUUo
Avc5JmLt9GYLaYnl/hzfC7FUMJyhpACu2apKJ8JsNAQHsl76ccwNB1Fl9GGcIjKo
6IobAAh3y0DaqBw0Uxc6MCLsQHZmW5J6DkRrl1VUwHtwT5J71jGL6UH2epMd2Kqi
Gc90iE1+yEDwJdYi7EEoAdobtNx0AY5mImeJldxXERgGBEiMnFIkWrBWJe/OiRZj
0/tC4rE3dQ1nMHI2Rhpn/bBXhAFDU4LbYuHhOnQzRvL49RXZMpR8Usk0nAeMYb31
3kRoHSpI6K7y1Wo3lewn06ku8H9xtgt7JOnfa9NwcTQ63penuKrJKcmV5FqdVa2x
PeZbnvTa7cqF0Y53lGJh2qvI+C395m+Y6Fcbv8p+zz9cVseKaCmSwW3nIU1PvFWO
k285OwYI0w/LoKFVcRA3lif3K3xS9nnKlaELegJPfDG7RmS0kL2veg9h1Js9CYHp
z/jUOQo+8hoTyATBVk7ftmB9nX7uWyoOYn61mIHw9T0v9wKRGjUpxYkWaBKN8qma
gepBbzPtlSfq/JBeiZN0Erzo2nNo5iTs4Y49DlT8B7IYGYthpiA29Txg4f5lkw14
NRvKPEB7EFOJ7BqOjgw0x1RQrPNs7nwHRiRPw1hAIjLLY6162JiQ01N2CrTv7Juq
1uNGROPCtXCxLO47llA+3CPpaaAur1n2lJK8+j1ZHrJ5clzU6I1ZaAbjt6aJePSU
X8WNJa8JQoT64GD0354AqtKGx/E5s0R/TLdcz//WXVcQmMeJbhXucN4bz6T7wsp9
jES8Z9iYILfxx9gscXS1xfYPwcvG0oAQ7jarsNA6PtzefuY/y4axZQuiQpZ66h84
Z++3lRyY47yYQ20Ca8PG0m8mdyM86sIqLOH165E5+7TmVgC96UGpyrsWnHfNH3t3
31ibPlet4sFj+hKCZ+oMjhyK82R03IzgnvUOkvqIlrFK+3f36p+PErk9KRSS7hVm
TPaEc5f630ZKee4PY271PV21YUKMbUH1u48gVKZm8ODnf5dTPrncInOb3zihVwg3
6MfGnYr7SfdJjOmvczcEB3ra8fz/8k+5OA5Cu8uLqQRxWe12eqYdbGZkxmUrR+k6
WAuNw6VULXHwpHB7zvVvcws813HhLDE6X1Uo64kgXhpPIHJ0DEic8y48FntwkDJ1
LJSXhpkK7TGBHCAV17CtD0WsLzcl3piWojFU45y+sWYKeZeliYWMwwShqn+TEH17
jQC/rMCm2Y+Y6ZGONcqUzTsxfMsbsoDh5xpfh3ej24OPp2lnhniWPbWRkWQKTwDY
XRSEqxEto3EZjNApX+GjorQSPueYPOZqeGSuxrVIoyi7JNlMGj2XHAGUCT+6ID2v
+tqD3lW7F4FV8Sou/GoggO4N63MRqZ26IHEObZjI83L68L9QnFd0wSYNN23RoEor
RnQ/TczyIlqEh5beDGHcWCibeQCgE0inl67DbonKQKySLw8ouqdD3MWwdJJYBYH+
STtR1KDTUT2nh41hvclIYbmK//teFxnY6IVPh7QjFZZJfiz2cNxfUVHbsiy1oXyG
PZV1OJvoOVlAYmDhqFrM1madewIzzVzwWEEh52OqnNSF39jVHyE//QetJfQVQDyx
L4RaS3C6I07vIMl70bhXlrZg6tlbrngUCA3iHA12jW0knaXJ+jLmZHr5IqkDW/rY
PPUdDN/sROY6yTFCLVsEX5Fm3K0BPbcg27xJOY8GIxHo58Fe70Lw9W55Ay64Lxbx
o+AgdV1BuBeFI5CNA9I/B8IWtKM2vCAs1IKQYrMCVxx+USw14RCQ0iSQlKb/ShP0
RMimBRfnnEGJa3m7z3U+dGWj1TiUN9hCXH5VfQT+++9Pe5kZ6pm66CXAbiO3FwHv
EZqbHa9hmvgwTw/JcMVTj/ENUQPScVPllqxZFoEMrDNLs9V37vQUUvumDXuRyzcj
0bWhtTan9PyBcwFX3Bt2oy0zWbAkC3DSsDmL0PLUjR4YTFHzE6Phvn5/nptpCjg8
GN+YYJBshzM9+6H+1f6hPA4w7vG7RjsAoLP7gfXBqIN/CFVfUnhf1rhReU/PSCsp
yDMr9ysHabMpJ53KPZUep9NOmB/s5Wc9wA66Ffqgh6YtkOhDBWOzU8nET9F6YEd4
HCstrq3On5XcQwnIkEhCNynxeBDW5Tl/vAmWmfEY+dPysQzhkP4jIjsfo8UNz7aK
ijO8bWPX5LydRwPARnE876B2NFwG7UePiwEEI37zQ8AHFceS9LWHEpJfMDq8pR8D
rE8IRp2qsk2uMmurhc8yPmeplZCAJTrRAiPh5RKO/VPh0S0e4yS29wbCAxNUheZZ
Vz4ViLVir3ZGQOun1wLIchB9akwl4JmgjO6O60zuu6vebgEeyGZLeC5+JoJrThpD
1PwLYqpW//7+mQE5w/4hOnev4lE7+gU71i7A1iTkDraXAzMZIWUtU7/j6YwvGH4z
coMhAU1dGpVfknx4mVs5/QkjdsmcIznFqbeHP8ik1goDIf3fgw7XdeHuydeIIgSA
06Dl0zxPEQzcfqkdM1jARiiybOtrcTidHB0H/aKxuFP3FNFEGGj/v0N5sUVO2nLT
vO2FnfHNaFBZAXzdOKIzLy2cx4UuXKfJUiBE4nY7TZq4BSHjwE9t12J3MdhATHPq
A0AWXY5UrWassZMCI2Qq4Q/JvUR9j0KlfLz0D7oztQ3pEvGLYD3IUHG8XEcIzdKx
DOH2rBIUQG2b5e1xSYO0JwMAdahGGcxKrvAzQKEX2Ub8MXvkIrRNHcaaUFBXRDn5
JMNWk6hppY0IcgirO5vsLQsYWUhSfjYmQq+P0Zfa6603ADqORCfZIux0OY+mn2RO
odrsu5nYscjzxKVav0+qQrRtk1vDFI0sj2T0se/zxqjkOCXDICYIr5Kw+JZX3a+S
qySY42HA5q3jSFaTdoiHDVoaYlh1y4o6xoR3KRZhOnXPK16jHUkIf0D/g2/LdF2m
FxmvvYGq9KreGqhV7MVSzpfq9KM1XCoO/eA039kyIXiaRYcNrkvJwQ3mOyy7nlLT
29/VX3QdjsIlr9FSTTtzx/O3vzR2DxlAOE1TFUoYCnki7oaIe1aHsqiikX3nk6R/
3YTbwJR1NnxTIzklpKdk/8P3fux5MeUv8WUkGsd7PtI0lYuVYOEXlFqo3zSu8Xoy
ql/kNFapBnKl463PYZ29GYvvrr3tmsxJQZgRTqpJ0hDXjlwjvV3zCpdiKUZidAYS
E9X45Fuu0llEGI1+xxbucXA5FsrKV94E0/vvjGcAXEIkh+3qyN5LatpqWT2VMlzu
VsI1GbsqFzSdKRFd5Ar6HvFWyOfJZA4grYMArEWlRDHKXm+2SSGm6tn99bQwvE58
gcL20rQlWePCY+JAtchUQZbiWQDrjT4IjcAHFMsxA65otlgfV4oYKvXlsnVHlZd/
8TgqOTBy/3kX1PpCZ6MEMjkfv3b7ej/7UHs4igzGvEVIAz/Z3klsCuPAev4cDSh8
bkghTthk5zSDGxqnN0iv7hX1zKAWqGhbsPLt+u2dRZN8qElrFBGfcLs8kyExEpu4
2UN2f6Y4g2J64a633PHWl8d+G8Z8JtqrjCw0fZ3kU7d4FVzauQhrQjEuANER2tpi
pV8s0DSrWnwlSZBnDXTgrsYtkB5Q30NVaBiw4EBX7O39mrHWn8VQmqCDSpLMzSDX
iMgYAS6VmT6mBPQc29bWwO3kvMdFR9xmApPPKdY0gU/XCqeph7W0Vf2qHSPM5X5M
H8/tNHg9Sv+iluVlnnjukoL9anq5haT5c5akeP/L4gmh1ws0nE47I2NEji6UrMNe
MTuk7UIpTD6qnWDylaJLtQW9ozLUn2jBKK2Pv2Yri2hWHIpCclAL+MTFeq3K/XZw
0S8LGlXqK+h5OwEUkiebpMnk03sMBceoCGZ53/Yd8gbfGmh5BXOAEzeX5wbvST3R
C044ogOKkNEEJGzF2Rk9sm9x4ICphttPolMUg0jTyGHWLAHDjtQSP4wi637kSWgu
xbplEgEePKaIKio+l0ZEz8GL6rzmgmTjFNBsz9tulqn9vWO2uIt4UNbX7z2aUw1K
0H0s0W9SPi1n1JN2HI7hJm/Ve45OSlk1BCLSErqSHcg8u3Rfb7cLpx3Kv96y3MVV
8EuKqb6OqT0twYA1Fpbz0WlvaUUeL46apccOv6O2xpCpI3GV6AjBq0dEs6KmOk5M
r0zifNbggPPZB26Xbbn8PQjwTwtT8OSdjvPaDo9QKj4uuS56Vz3j/hbrNApcT0mW
RYPNsvfZX3LF9bJlFUEt3kFXxP/0PXXonRiFwVM7FGCTU/0+9+TCwyW+r4XEmNqe
74BX/1vyQPoJcXi3UAFeMWvL4+v1AZtZ9whPhJjGlADtcK9NQilD2y8S7Q+MSYjd
yk3mfwpFXmXYngB/bIO9hJpxGwol5uSrdSRje/sJGGz4tYwcjkz2cMN5aTxfwVOb
e1KRce3wK4XyXi23S4CDs/Jyhx+GdQ1x7+7253dXvA6M/WfTNmirIEowmOKtDe6e
4sqar/PhFWm8Bg44jZXAIfbaL5ppfNzjfT1nylQ/1UJMTBMMWdl5bJ+d4RzmiN63
GqezhPsYEpuZf8gqsFjZKrmGXUN4uWo/q4C6CAz7FlpgROKBq3f3dpT0nTO06O0K
jsTnBMenbuYN4xUtUEfAKPj1mAdyHEwPCmv36uXSeyrZwpSzNNx2nAp9iFnYIjgF
qeiQfhfOyFPFf3ycfAL2PbLxyc9uTtN+d9edPZXhh8tRRVQBO6MKdz7upozXEnEq
IJxONTztw3/vNVyE7yG8VFXVDRM059Gjy7RXIPoKy22w3jyKW10nh/cZw/fqyEUG
Kv3JJX4Du9x9Thm2jcd4v1AvJ9Th9wtFhlwd6ImgpB+QS51yJqHkYhqSB/N1hfQ3
325BgzJWl58zQ+ynWbVHV8iyYq8V0PnGSLB7G2p7fcmYlb9x7YZdoDbYFs3mPpan
2Oh7ycSViuuSp/qlxeomxjvseC8U3Bxhp1Y0I05UFGf4UNQg+RhHD1+vsC4yPrWk
4gQ3v46go8GQ9TCo39UsRdcK6pY5XsOnRQZu/hdZxTsDHJLv/qu9261hAwJqGjrn
jJLFzTamR14lWf0lYBcEi4B/SvDVPAo90yvYiintWo0doc1/8zLgP55Ha6MMi9Fl
Bg78DuUH1kykyjzi9DBuDFShh0fZsOCRb5O1XtE6B8EK/+v6DeGSmiZPpazGfBXI
ZTcKete/Qtm7R9ka4rjurD/JAEsZGpzsqSFaQMuwvF7MPXHwc0mN1MHK8b8r63QJ
HWo5zc//wEQi8wHl1SSti/ioqHdTCNx77ssNnUEp55y/xM25NcxQx2H8p2Cezj02
DF0v+sB+KvfYo+VOws1+4n6ap5XcsuQooDEAgNNVefZITlUwssMdHcYDAM0uRNsJ
UX3PWFKtV7KQ8PlVxkOWngx+zjMt9N8JnDgnN+KyPFV5n1S8i+mzgC1Q3J+HVPhH
UFwv/HBzj1m/74QGVr4C7oLmX4v/b3TEeg71U6dvuucvmgWNpPFlNsdDcV40yPfd
qYr9TiuMqizsBTXzzMIyNkV7SZf0pmkkrjjJB3BK4ZkI7r9eW61S1bEOf0NGadlr
8Fwjh9TGc7ApPquWcUlcBawTJi1ANgO/8qBJTek21AfpDn9n2C7I8fOb1CNg1DVI
bgjb/3aIrAl7zS4N+hZmypOtvR2MjK9I79JI8Xj7ibKaL8gdevtwTrOtnIocLEB3
OBNT/eCyoyk7r5yjqjRCzmjpF9MfXLlMdNeQJ3uTUPUCZhVwPpLiZncRut7ZKQVh
sPou5QixUulq4epBQ672Q0eV0BI5igiKQuRHx2XJPSf2uEhZ8wtm9bzouKVqngfj
O8qsqmCG5W8XOjjzvKjhODyDiRvg4/Yh9tb7w3pYblENxN9lOj9lYDD0C/RXEbBJ
2zZKN9vR4tOTIK0iO/hQacfjoi4fP/MdIxW/dyZk8JT9ctrgRxiwoy+BRrEbjAg1
yTGVBFRNWUj1wVT9wID3L82G9J6w/KPG2+fRsOlECK+gXX0BbBjQWTnh74s9CVHP
WTlssCv8hw4nNMI3mW247bqk2u/ibO3oGexmZwY5Qz0e+uS7OWA8xE2flZPC2H8+
Lq6bKxtB+dz5sqQKvCtTo6dIsg7PkAQgLO/Po2zx50L+qyRCqJaqtHMcXKGOawlT
IV4KnE0XKN36q7YzVb1G2kpuK2dbvi7RbDJvRwn1qe1lZ570LXi53G/SVSMeDM3S
0e+GlIRUytsxvYNaEBv2aUg0kTfaqDNdNd3Id6cOyqZtPJ3CYPACnB5IPeDW7bQl
i5/66q+q2VMJ3y+kRi0jgN8a6ayKQ1kFqx7HF6zFtgZ14zQk/cZUHEyzXrGdNBgB
t9xhqpbBIawMsKBReiS1b5Dx20QQfNFlflkt1tcOcdFsCnORSzdg2IDpIvMdNEhO
GFcCN2hk7ruk9jqi9nMqE+CIo1tshj4h1k1ByhqYxv3c74kCWAXdnFjUYdCvibpT
GtaQc6w6TdjSrfg38rBwHJp4sa8T9XUgwkWHpTbfvwGQdmrg55o4NAqA1naeIsC9
VKGsJbdusMhyrY6UGqyRLvi1Q2DnRPZQxQcndZabYrhCQr5GHjUxORHAv2vx1h0a
+sOEfxu+08+vd0bHno7buiwwJ199eQusvC3ONFJoIhaFCFrx/C2FB+o4PGh+cj1x
fr+d+SMkGnHZPcRS/UHatdykbHC46JIlIwt5uV4wRqzQpbK6jdkocjGiUf6iaAO+
cAnZhG2Uj5cLt9d6dS6P5EtZhJ3EFbJdwWRN5ShYCo6L3neAXbQyC4sfqZRSzijN
6qjhYT6dnBDCYZNchaM4Wr8nMXwRNTHedWhX1T17mysHMk8KIeFtX9fk5h+y0yHW
+ra9F2As3yE8+L7//Cr8p11wsfBTiITzSVHbSGgCG/OMlnSZC1qY2Enwy4AWl27a
76/ihL9ddPoafWmUonVc1MJb1OcBTsvx/uchkuyqFqiQqFcm5a8zebJNfewMc6Gh
nzYr5h2AXS04ddYFuJ4670dnSdYkfMf+aXctOh05g29enj8YiW2C2sEbsGSViecs
Vru+fCg4KCzxy2vuPpZg4vi/pUJzwfFulSsPpYwVunw+oENBTtMyW+ZmpUuJvbJ8
A3rQd2w3lgfwITPRnPqFJpQwPDKHhi6WJlJ/8aH7RHdH8vKs6JLBjggnlIhme0yj
bNXKW38KZ3bhi0oh4rXPPkxDgXyc+MnB6bWMCLd4KUGC4twjxlYtCCm2CxHKNYhG
YX9IvMJZIkGEc4xOoVf73Lp5qjG6QK/vUT9YpVBC1miWAC2eN3gHztITKG0Lp8jv
Qpv3vla+3LgatSWZ7DOIDm21GdVJA2CeniS22CVjU3ijkVN6VVcWWbb78Y2JhGSW
cldcvwG5kbDdjH3KtGkXmDpfXbHjD4hizW6Us/hkKn7XzbmEZkmnLQnJLlRCY46P
ObbgKm+VcvnGIDVbbaN3+pGx8u7DQ+itzQRmPW0rEzibGWtdMWaLQjg0CyodsWhN
2fb3WC+tBnOGoUnY0Jin/vxCzsf1BWwmpPhfpquhZm9FjFN2mExbTWWKZ2fGUM4y
GPlb0kOZ1mZZZxvgedxNcVEPOhF13ZHu/Z0dddKRNbW72FvNJxrkBIaS4r2Q220t
hQbWHGnGRQu8UFzRROBzk0b4swMsHvdia0fgVmq2qKGZv7UulJ9l/rDhFngHsuEz
Db2X200+JmPnfwQcy7uy3WyWWoF8kkGl4HjNTp/vW825AD7D8m0o74HD24h0AHqy
sT25meWOaU3Fjz+EiSQqe5LhcDRQPpp2S6FJ+jV8bQFXjg5QfHfxGxnLxIpEker8
t89rlg0LdHeULnG2GyewnwzO9W8g2WwkNBeXABPKf5QWgIZS9+AFGJ9BGd17kolR
xppxKq2QrJNhcvGxk25Y38bX5prBINOP8B6vbCPBepCQNaqGhaGKQFBtqYt4pRqF
gxZszgK9uf/48WossIxQvs+HhAjOuO5oG46+1wBlkh+fptXXYhg1KR+CNn4iVjOR
Omit+5kDQ2FKCO9kmFyRDuVhIZN8tDZjpmRBTgRVhB2UtBW3PuofOu+0WN5G/SFs
naPNzy98Gqs1prGSvW4yFM+XopKtfS0pL2CLs28DKrbKrVEhh3LjQYipiMTFXpkP
WMzoyofZBuU32I5Lmfi0yBT9HdPfjo+uHAfzyGn/Re50On3ztV3vZH2hDT9x9uAg
Rgccgn8TYdY/ppWOvQZ94i6NkptyLwiXbvKObX3kM6OYFzuSBM1Vz0TqrK87Yqc6
JOeSG6GKnrjTNlJA+Nj1jbgnqlsXv5i8254QgMK2tt0gPmgHZfVMAzxMnFU9tYdz
W8ruazEIDtCJTD4Mfct/qOpB8NEhZzSv0dZDZ1S4y6t32HX6GLiF9kTihs7IvCRk
vCLhemTxG0eqUvzFcdZEFG3dvwk50+/z1mqMyDv+IPjtdcEG11IaSUyCjnwiuJDB
ktXbGiWhy0heYVaW76yPiet218iSYruDauS6IapMzV3tqPAnhQIEtm+JBNrKhyuw
4AOqd/i7rSEb0IRDuz1VObAEVKTHMruMJHpUJSw0zhXEPai0UWdCdKfUhwaCdvCI
myEor0UJUjgXe5tBnAoW2OO+JGWBCGoayxdHdhhl63laJyO0f531VuTIgxEarD/F
2w6mEOdL8sWwN/zyTvXWTQlrh7d7Eq0S5CvQzZrG9pezSYqyBaeg/ARHTJoJUeVZ
PBH7gSbRFXj+CnNzmXN3GIkOxnJbtWeLM8zwzyjc7sAZGKs7Wazm4sV9ASRPDGwD
Rxt74d+OHuwpH/p5HI6XriEy354J+DeAVbDl2/PA/1fRpaB0XpMz0KUnGSQJrezd
dPAn0aulwJgbxRkVNMUkh/a5Nl+NbZwRWtnCNA8aZiPhk+ft67WnCdPwC33IDLh2
nUzy9af8TtoBeapN8T4hmYiqsaY5VNeTUFXHhNtZQb58s1PSFdemK+slAGwTVJJ0
Sa/2yByBJnuJ8M9zi25XccMbFH9+Orq3noOTA5qMq16uBJ8xH61PAbQJkhW3xRfZ
SPw2oAiu3WTCFTTT90KT33PQVGFXyxjPIeZC3YmayK81tapDOzTfyRLK156jNq/s
Q5A+XfSgTYRqwg436ZEyN3WMMNAnM9BLZ/UTva+jYvJTsQAjvqklBpVGDVogre9+
G29bDQ4civeHObAAv6t7D1gNBMDMyxZU4BD7cwiQZjW1NaN/+r0dBWdu68vN8laR
O6kBOvqLTfM8qeR5w79ZjfqOTtQiLCdDjLdahHdPB1RvP4eMZnlvYUWpfzAhJg/T
MHfhShwpSOFkA5DjmR7XSdBIJ0K4MxcVYhwaPu00tpG/ohw9T34M0QM7kPtLymoJ
HN37TTrG7pwk9RhmA54e2sRNbz6iQ+BP58GVtwUuPrrZjwB4nUFDqWZ5Fx26HQFZ
mLh3ZM+q4wjda14FR2iAcLuuU+Z/8s2qxHQ+08egJdaRj4qR66ICmArz9JhXtO2y
xTOt93Ykt7sJxiVmQFY8s0gvmlb2YyFVoPrIVp4QGZntDt8Ec345BjWwf79reSyT
8PZLOXpprRKaMJ2yC4bEsRO5hr7+QXcL5b/l1fWLC1BJFOi5KeZ5F+REQ2Lkn3GE
464jBnYAP4Wa27OGOOnW8MbK6DVz6xscwalF+6vYymdlcqCVlqPA42S3l/r+bUNF
ydTpLXh3znBd0ux09DrKb2PZqqpz+WNTCjdBAgLvJDkx/hG4rqmAqzzBr58sxc8w
9QYOptsHp/vmUyq9ORI99Fux7Fbu9HMuwsI/PE8fCkZ1Za6LZ8aki9XPZrPG4mnc
9oulQb3ieTHQVIr/GuCIH1eYEiekOljJocpjhbiFmUSjvGkFNkXE6yrBpTQN0dCU
dM80fj9I8SZSzHOS7Hq73OXEoWypWUUbfZYhpZGnPdMM7llIwv0Fvc4xoYh4R7iK
j1QibFQbIhM1RhwhygBAdKprRb0RkwtFYl8PqFzIYySJen21xuFtefeigoT8CUyI
2OXpCWPonTtEg3GIY+2MXFC7GYvLQ4lOKKXw3IKYJz2OuF+9AqD1oo6nrIjqU/Uf
KB0JSIAV0EgxA9441VHPgwSFhEu5auoPARm8PhGnl8naElftc+eoUhpoAVrrgUBy
qZm34SqNDYl+5x1O+iRAR8zjiHJnBlPea5HAwVui19gr7+G8+VuIhqlQL0Q3pteo
FARijPu9m3F3v2IBQClOdRfj+/ZWwLWy+nH7pQXQ8A6lWz5iG2XKbmdRIHxQZhhu
MmvC3wkoCS0C8aMx8Q43dllEkmKmMmBNWMxsuXWleXfmauvIQhqrytBi94Sy4ygn
GnFqC19j891MwYP1KjrKXx4NeRCD9JguP6yNfsV+UIgDwKZnasLkSQQwZKkze3nX
Ki0x9CUdswPsGtFk5QZoIQnGBRF89xulIxUDmdPMQro1sC7Cw5pnjL8VJIVyKekl
hbYuwSFdc2/Eh7lUB39AyNw1RGR+IQlP/1j7gO/e2Fni120+mLyvLM31liqFMMW7
+CHY1ONypskEJR7DhqGfcm0XZCmd97N+Ye2JQrw8GB1npONK5s2UmPBRISdZZ7eL
KC5hNu50HKi0D8YZCQ3dDiXOuxOXhgLzJDmx81tRTMAnEV386ZkcFlOz0AKJc+oB
Ndxx7voLeJ6Dck86DJmlIstJxXlOr3K4X9QqOi37AJhP4KSfLtL+dUp7OuRttnAB
LnFnEP+6CyElKYVPeBvva0ztYa2K+CQD0M/p9veG7nYWWI+5O10vEIUrN//gWw1c
V/XibRM0cvTZKZ4gIuYebT7qKDgnY0ADOpTFT66fuYon4QdLm3Yymv8bSttrZjw2
nP4Kqt0klZ722NUva9lWmLY/f2qaqnzV5NPm0uwUC98VH4iEDI72ukcYdPk8O89X
1f1YkjpmjBK7bHar6a6vW9UDPeKewMTAiyQUYl5P0I8pAiL6i8KV26coIpJcbpQ1
Rho3fOPsvDzlPhYFvqtut0jz2QgjZtW2DB/qWGAkf48lFUVIqULaeBCa3fzIJ4yD
KalH1scKLRS54J3WEFDQzYR5QEs3JPPZA9B9+7kh6EglDob+a7ywU/MsaT01pN0y
uznwP4gY4kVLbC4tEBqrHiWt8gljtpXYibM66wvKDKoS9KEq4x4Wq7zXG1qcuyvo
ImdA+/5N2AFRzJvaC3J4n3YF5QFcn/qg6QXmCe5KCrIe85CCPgUsu+bY/RZVhd1n
JgDX4+jrHNfxHrU8f5AtqzYUMYgbK7kZT15aMyaEKSR0WOp7JHTMWp+ggaVFFsau
+SyW//B5zU3x2mAeHc3dVChUrYsROiXCrk54CmPU0QXCR85sOiEeYOrCT2XworcU
AOh3W2m/H5+5Iu9qqUUM/ehEAkn9Ki47ESk8t2a/TGby5CWpKFJTwnEZjVvmnM+4
Ytxml3u6Fw44KUmocQkpyMmylRC1OBoQy3/rvpd/8xe/y6LinGd2Rn3ISpl2NU5j
bvD4BdHN33AJqbFV0UstR59AMEBgV4s+3p6p/e0aakKGsGy6tkTTjUapvB2KjV6I
OfUl2iJpKna0gMmzcqdmv/BTSA+XYczSunrQc4ftv6jdhxuH7Oj5MpT2Vaaxes7j
nbawk9gPvnwhFSqyj9RW69HTJJPhHrrYVIV3iEUgVOzE6MUWIMpX2vjmAYn5sZHi
4rdbifw1XvwWgdi4rZmtYk2xuabc5pLVxretaDqlfCSkfPiJBoHc/MffM+FNWMJ4
u90WmNRy3szy0cS7r38fE9D/XEYEoX+Yc/COpmgKy90tIRhQQh27lxhOjgKgPLJU
j4w6e9oIzRtJv/VcU2PCruuwIgc2mDIOKVrcn+HjXzxvmOnhQETuH87MvIYqIZ/q
PohlNO70KRQ3xy3ciGb2YdrDTs4ennrWMnGyuIWO02UragcNwlcAJC6dFRPrcnfw
e5TvOZ/7xRu8qK2NSYpNMuBmo7/Yx1tPlnkwWVnD+sEZL5hk1r7GB1DoPF8G2vkW
ZYkuZz2iCnS2MYqsDSMo2WR57i+jMTG7wYFFLL0SVGr0/Xw0V5WbdLZGqsSmMTLt
Opxg+CFR1Cy7LW427WXk8gzL9Ho2RO8cUMWAOMlzMaoCiplgGlX9GG1xs6mVCyqC
nurb5nq8TlPkGDho/5k8LUCf4SVWOSBTwfgBs4SDljdQoeg14V2Nqe64caaCrmsu
04+0Kiby1W7XP+ThempuNWlF+VOmId8I5SxbyY1tKpzjWBioW5XJJl5lKD3vwKj7
p9/mJoxxvQWbV7cQDmEjmhK2yM5yYcyBKShSQ3r99naZTJxsG/4CV1+emiuX7gbE
V7eu/VcjZizm/8K1OxylPvc7LhdC+NZ+cidZ9Xz2HP2OI3G8Td8sTD82lHr+xvHH
atXiYn8eBPaP9BpxGLH/joLb+08+bjT2lmq81vqzPYkJFIDvDyK7pzOlpn7m6H4e
4GJXwyQ4vVsFBauYVisOLYlXHcBKis4YT0DnhQKjVgYXkUPP8vXGhPfVS56kSp55
31x8iwjK+HCbzyMhXaDS77AQ8lvs6JShkb7PhpCz3b1CKsZ7r3KlT1ZyTUmDNsd2
70/PVzhXpqfYCFRkpO8bJPIcmSFfqYzTXHttYC+Cw1brbHZxgXQRlD9P0N9Dl2+3
AyKYob9H+X+UheIY0gE29vgwVmtlUYPttuBbFZj1UaoMjQOaak83tGLpgizumwfE
LVx830nbclaOwX7D/vLpl8zWD37A/MITYt/RC2eR9HzZmXHuFnWyDD+EaQJ6xLAH
/Y8s4rGlZl1MLYhi2yrYuWrR6axrJpnewTjTAZy8VBIb8sa+C5S3+tmaKvIOLUAg
G0zYIaS+3U3noF/IG04UwQzitNe7e5RPsxzhGatLVGTfFCDQW9z27XDijFhJ4Nd2
Cw2VVhR+GuvX1a0nMAW9BRrKmuMxUqW/OoJoy/R748SJcu/cllxip0z/Q3g5C0Yj
1YZlvxvELtegWdnL8fU5HqAR9Eq0VPM+tOUj7pv26inRw28uFgN2rF/o7tI5TgPm
q/osZAYmnO02hSA+8FzxoPoW+F4+7qc/uxdwIRmikrqJlWCwznjDa+cohIEe7Den
lxvV+99gJTV/zfpibdkcUkmZzrCeVBR2t2P2ZtGGsuWIaO6pR76W2Ep9oP1/5oJ8
Q3SPllTMDpXkqHRLU4N4tMY8X3Rth3Bif2Kn/XxQEp8HT6YOPhxT+R+UuHgRDwnD
zWSSVfUhD594tc0vrQpjRDqOCq/qmyfmvWAXOC9f9XXqPAQ3W0mOCMgvfeTRTmd5
N1hDuXbjmAcHTOBFwJz1XMhBZKJ4p7uQ1kfpNwfKovkPz5PM3/ci4Ba3BPQfPYgj
2QbD9eYbBfVHB/YxlF/4JhzXLbltW1XoKqcivQ9aBijiKe7mnQRSamWt9D6+R1+O
+O51+SXg5Wew8boQ+MIAVrPm0QeJ++XSKtULbr0tBbjLpvWJfUxiEkrfJbF2Bhge
W4xrL157stxfZ7sOjQzZkaHbhrnJLUh/3gDvcbvIkDlNcY3wHx90nwP548nZ68UM
AUbfe54/zjqpVVCFoDUdmpqJa1uXatQ96UvnSglINq7+VM/EMF5pmIDdl0KhR/hq
cd2UirxcWE3yL4ZA1xo7obTAfQCtpwWUqiUSXmuNicg4MsJM22SHsUklD6NmsPZJ
4nRdPh5YV9b1yImYJWbRWQqXwENZYUXv1U/+PSsp6Lu8hXurxEs78QR3q2P5pYto
0uFFxa6E/NFHUcK79Obn/Hpwgm0AfQpvAxMSfp5kQgfj0W4JqTrir4xtP4oly6sS
WorDuNAI6tfQGNao77f9QtjMjR7MGOP1jFbkxmRNqxC7bRiUMy2mluYiqQjP/e3B
GCz5QiBonQtJ7SkwOG0N0VSc/6mYAFZUJel5U/xHeKozH63upTf/CMlhKE7hPcU8
CB3euXikDvNk/JeqhGvkINSsz/CPhYeZjdJT9IjKCDGoICuLL0WJWvZdTdFnb8qC
lrvu5nhUc4FVGqisTQU/RZ2ARt+Y7kbM9W/Dxf3a7hAu2AEAgtfDVuioImcxuPtj
xmxUcVmZKf3xo9kRdIDWUKMdRuz6FQvVAWSyTJ/xz7En8xlAjByMc0Lqis5J0z+2
C54u/1lHmfXz4IPl156QBHT4DgMfbEQ0KrYrQjJy2jd7S0JB18p6PiQ82dh2oo8n
5JLopSuvpCfVCL1GlPeVeYWi6jYUHnsD4ZxZpVWmcRCwsm6AYl3cCeoKb9IrZXHc
YQP1YepLd0s0MMj6AECSbbADV4LorVQ6YgbRJ7IhRqZddU+b6JhtV3Ww7mlPA7Pm
fnYetdHwF30429LM3UtXB/P3nJtodwFGzAqCzvknsKtbU15IsmwHZiDZIr1bANQm
5R2+D2G6WGV98BQOzYRDub4km6Gx5rQM6Z3RuME8LoabyESIkee6wF1xd+m9olAY
AiZyk8VQGgWxqQw66m2LXoebMHk4Oc4ojgf8NGB5oYUL3Fdt9G7ExmcF5eLlB84i
/Wh6xyNc6fdTC1x2BV1wZ8+G+r+EcUTYEouQWmCcnqd1Py/L6l8svS5IfCmytT0s
QmNvVoVAZbl65UbR7IaQmzUioE7NYlRUfdEgX/m7pgVNW5x0OZApN+Gc+ctdsiWQ
giDrlU9TTywaSCmBWO+MRYEVzbRVXzkz/Oc5tqHKd+ACObdtooPxqdLD17NtE3xF
e9QsxP6RIp+UygDgGdteKIhntSOtChZQS3FJqg3Nm/uNYFXH70AYY3pi8VWSDJE7
zpxaVgZrwOlD5hWMQs8slRn539Kll/cxT9mKP2Y2ZXYYueMzL05+0p8GhMb3Av/G
YYzXFWktgqgD4sAmU+jJq3SDcDOB88N+lX/pvHwQ6OttQjHJiiQJ80QjJoJxzYuB
hYzBXeZrn3snqDAtYqrpoot9lY3zesAG9fg/VKX8pb7snIjqTwMisinB2MVO/BIA
ppAGHSo6GwnnU23Wgz5ehUvDlxNVZsGZn/5zSKgG/Ww5SG1Q6avMFLo2+9WvpzGm
tXAjA5qGh2+FMMmMslVw6wv7+DX0hgVLkhnLUruVosQ20fKPisiiqgaVoApPBQRT
K+I7m+hLBZQoj2CRAO1rlO35ubymt7WYhuzWdW+4JAU00OhzKbPOOsNfcFq3Ehtu
DTYNrPsnVSGA/DBrkmwznxzTvJYYePrs0lXv/IwPL1qhIik54pHNAcHtNBLhI8+v
HKP0e8Rq9XY7Bq7T9kLfSNbebSmCSR/3id9k7Nrd+rylgBdWbK5RICl9tth6HrK5
rS+TcT4mey+u47LN+ifzbGbudUfwah9OEk3zU4GT/rYhByA3l2eK7TWT5mdeRyzA
hm96Y7HgY0SEnPMZ5MN/mZ6yPZ7SIbDtmi1Zxxte1I3LHsEYD1PUr5WdFqKIpJno
SlZkIF/+K3gnZoAwCgzhZkp88a1xm+Mf3zafkuO/g3DwBOfovtrwLAJGz3VncEg8
x7oxqsv/nuP2du68hrL1ZiXaoL7GRnkd/KpHmPhX5sneQvoxpBooHr9JGsX5m05U
qW2LAB2JW+J4YJor1ZB1X+yJukzM88pPjAp0ferIuqIQbH5C8zf83M5qY7b8utHl
OfDiXDj+zrUQo8VdSXqidAVa+KUETPq+8JEncIlCmfUPKEzzFvr+3Dw/N7OlMcoJ
fmqbf6XW1ezDxz3q8JG9DAZVkBavfQOAwf/LUwG1Do3WX1qjalCYuYd/NxJMmT/r
Utv1wNrPqKcqc5mLvnusm3zlstL+0JYqI9WV8ChSZkgKe/E9yN9mIAyrFROolIlO
kkoWE06U2AcTliXXsf1FDI231skwu+VUx7C0mY5qvs/HmC5IqsZrKeNU+/qTSLO/
GQCYSt89NAYVzQiReuL7VX7+sgCubsoz9lnNcK7mEQIRWERE6LoOvdT/hRF/RZXC
5M8LBcUtuAScTV6Liu78Gx0TitGPXQlVCsdWaozx/4t4HKrRmq5mvYK/OqCBQ3S9
JMcdDHmIZF1gQPFAdugZP+9HpnrifGy3hMUQ1tfauoPTYoRRbZHH8V33YV7FbWAi
Pffa/i4rpykicetJEtRQBV+yr+UsOaHpUxCHhYzKQeok8gX/6XCnH9QY99qiLM/C
hbVruhsy4rcLnTASbnLb/F5E3yoaAr2hd4J25Nxi/NynBTh//Z3mD6j16xexgqmZ
PAw8AxcRY3exqd5KyeEEEj1J02B7cetF6VvLo4vgt2MPePRDmvX/L2Ablct9i6Yz
ZlmpX5FjfkTRkAxTlw74wfoRtZ05JQXLSOslIY7UXEO4p+kidsGmEABtAqc4Enro
9WWyso4IEhqtOpwRMziKDESab0Wya/Ix8HJULNSoqLRIFt8wou4NmR1+a2hNIUPt
sWfJmJDHbj5ELDz94hJlpQxcPyqb6pLAQlGl/U9ihZt5Jbcdb/lIjkp+4BV39uMG
gWrBgseBlGrMTaDSox3ssSIlDIXRcMEODpWHCCb8ux0S/aLakof7/C4GTYaa9bgM
YeDb02kvyKHO7xnodAUPlVzC1jGi857RqiCwfdHwQ3xN10AuQvhVDAHIhJWZUk0X
8yMdC9Xft2tk3z14FKEn4WOdILKGztVIy8hBi5KESU8N7qVjFFtY2WWkmztdDwUF
R0X3AXSGyTeOiNVE7A3zRHjl7qweEHMZUPRzpBb0jFEFy9Hi6hCTenL7KLYj/3yq
ANNSXkoCfryyFIJtamRG58aDW2IDMppjYFtytiPfAPsJuThv/aX3f5vnYWdPB6nC
pvRyPhUk0ncfFcCn/nemNGpvTOzHtYlZP8v0azezuXbSBwZLOTiyGUw0H+W5M4w9
8mHLmSqaMCcG4KglasQD8vY/mMAhJPzuPp9BcJbQJaFu0fdLe4HzgQt+YuoXQakK
vpEgLdnC0ZI3vsAvXh90UOGeOjiayajShva6hXgh+47pBZnt7LAowbUOl+siePuH
twftBaCDZnjsFfc0bKDken+jUa+dFTlsg15MYcU11DF9ucP4thHrZQ1UfGBUEDvF
kdGL2zIxuq5gECflT9+aRSF7eOYepxaxDBDWLz/EQ7OVQQEEbrN0ZAOxm+gHmIi4
qzsOv2Dca8rA6tlcU34LrSQoHoW46PqgJetTizafansStkGeh5Xc4FbV3tgrjXSi
PBPgLr8l4+u3e2YXDvcFqt3+Hlo8YeToyxk69czGwRotEx6uKIh/Rha3HDBJkqll
FmGQPv/2nuyH+vhwkVoK+vMGZA6nHgWUYRaRG6oTs+SkNlc0afKbFsN5uLxtxMOg
5G0Bxtt48mRcN6qhe3XIVsCgFjdTDU7VuvzzfZj7/6+D2cc03h0pebzEwWmJm+Zo
qPPhPfxjtDqaYz/wd3ifMEGSwHCTmntZxGD979U2/pqKFnAIZzf2YO6XQdUYiH22
XV0xKMLJhwo5iQJv6B76lq3muSYthcjzOmSF9cSiM5TpXdAxGswfhnjB4MqWrjvs
wEgWN9FFbGBtr3ij+gua9lOz1S8e6kEOzo2hb2WGpz0BcHkm0reCuE5KSoxmU4B1
P84Xeevax9orMesuHFyF11tYqKkfV4GwtoMOBRCuBpAl5jrqPQPgmti6gbPe/Sn9
UzOPTZDg3/Wo/ZddvgnqgwnIOf33Hi9B0dfe8F40O9acxqo/un2sP0fSVFlsXtbB
hrzibFIVY4/TcCWjKRQuxDUHxcGBWlVHO9x6zIon2V8pGeoSmVEa033ON0tjY42K
nCYfkaxfs+NNJPel+14FIXsCac2m5tAmDP4zF0wW54shziVH+U4mIu4cBEbR0le+
ZwPNml6KP8sn5FLjCoJ2Mievu34qIRRfpgNvVSe3tA+jYb2jzhF2PluAdaULASO0
IBKdHxwZpaqnfZDIRH8rUdlgCRqMON6ncM2AsIX1lfWVxZgulhNYk9kS27lhp/cw
zmd4DiBMupcaPvYjEVFpBkj/Ho0vuw+k+6keB3WNVLMtNYdJjMk1tqgAX28IMWgr
f4ttkPwg1afjdplNlbLNvBlREDtNd8WoW5KIduL9PVIpdq+lZ7bOR3yV85W/YMDZ
tA82RNDnwhTAb45JYA+D5Qb+wlY1W78CndLbUYbeEFmeTGMeRvRhZqJrCj5tPB0m
l63cIluXdkupPvyN5OvTdB3z4rvcRbudbHVp/cuGqCE9e0ToqiaasGTrH63R5BxR
BdWeImI5IMab/ZMHFcRys95uvZr8R6Lx+en6FatM5Ja+QMWuRlJuFFCCfEl2mLja
pp6Mt2Mm+SkLnCPYSLykiW63wDpLDuwydd0WPJDHAXQPsCiyvLJBJGGmg436yQJK
1iawLvAkDFCPk7KZ7YVgf0UpBfhxvH71d56ao3oTRad0p0xJ4PhRorEiLwWgb4ev
A0MSeUczLqlXFcJeNyaWT3Lfj6ZIKFqgwQe4svxi04NK3a2BejBbyBw2nVqeeKfY
01iWDC1cNu3Zhjbvt1H0Gp9PJyVA2cgVboCoTKRHLoRWNKBNxbuczzUCtheE9zNz
OehP7wFOZeqbKVrE7CIWGffMA4ub8ci4QVN4JmARzpt2V4gxOCZfwummaA9mpjwe
chZoGQRDnJecuIJ121ht5smARYqqepr5794lVtpbpxaGhqSyPQEdsi1y3Hm7Vs/V
FWm3FYZOLecppGC9VMOlr/EXeatgrUgc60WgzoRnzddn6p+aakiRnyio+4abAZYX
lzLlXrdONxbaU/QEl8dIIwyTxeCY+jHAxRKVaIr/zDn/Z+imHYheL5tV01qVvG/z
s4X8r+1GH8c0NzU+Ymeu49X9hplKnUgfKJfvkFAmjuFF09zxGYzSa+XHXPfIvRL5
N78ZhFXFzQV0SgPsQAmLzzEMsWoeW5C5al0xt597RD24IJs7E+Of0aKykcmRXbrM
JFmfe3j4YlMhsAGQNUAKTDtvR5Q9ZlVnvaJ/nVEru004b2MzLpyTQzsg50vYykV1
7bml0UEubcadLzpYWSxLmcycGSOoOMvMVN4yYP3wA7A77mdc07ZcQONOklcsj9v0
7T6L9wfpKVy5FSUs7nTdJIwH1Fb+p6Jx2QdADCgsIyH52fcZdbPGtthHwjaAmqjN
5VdARzYp3a2a0tjMDFjOC79pqXFqsWcA0WCFqFxzTTK6IKrmzdL/WVnHVt7F8JwD
jr9F3CVPXm0wNnlIb3qziMa9BzkLD23u3Y7OF4Cg+miyXBiJwogYZC6dcrE7oNEA
o3A3Z1VYOOXq5kkGZdJ3RsXNy2hDeW4gCJCk4DzypiUIIqtDGmpbkUhLEJWJmQVb
TzDO+qJvP/PKDUWu7BAFGaBTA1J9PFWYhr0lQccaC/7iKmrp/Ba7+LqXSkz5siFr
d94NcDzA9KIkjqWoDLzOhH1v8La2N6Ko09VlZ67HLv0OiRiKeSWRfIt1Mt2+Ig3k
2OO/2yippq3jL8uJNg3W/bkgp0QONROSPUTxIozh/2TTVBsqpTv+ao0wF1GbQUPz
Rpj74GbhnK3iCmnBGNbuqfe4TyiODyU5m7u1i49UzDfp9WjjTwnW55wFk5Dus+l1
XHR4bvSM4nSSN9+UT4gsvWSJ0tzVMlDFwMpU48QAwQhRufWT46lyxCjj+oMrBocQ
BMy58iOTbyYJl74yxCkKclXTsTYhLgDaIl9zaj8Zrypaj1ebBvWGT4NEKkjSoGIs
U8cZnpSRPyc6dD+nxwg3by+03FS0tcAhc/Acpygu4KUnu7EuPigryWSAfUTneBnW
lDL60o9ydvrm+4oJsAqrrvucYAydSJhFcIXTAPfJ4h+WCe+E9dlbuCTx2H+Siyd6
XzzHUVriwhBC+2qjkP+Wjg8ILeg18I87+NyyZhOQmIAJOejH0ZHcp0IO6IWxkrdF
i3GCOat9E7JiBPImSoaFZ1/b1OleqJLYvI1W+k+nXyTcrK936PHWrtihPHQ5q4cT
a3jYvCP+CKU2E/ipAp2PnUJP+iKBBDID/1YALPwVHEypRqZjdfUO/QudBu1vQ5qT
mVR4ing8DgVszaOQ0GST7/RYKsT7pDcuh8BOcWw4A3CS7YAiKmYDdv1wlP0z4c0C
FTXj/qhBW+7YUd0LUwgnv13ShazywhpKcC2h5sOZ2ApgHelYxyYX7vqPjxJ8aT/8
wYJU0eQ139nK7tVXI7ZpVH20x4JdB8HsS21o62LuEwa5QWlQ1U9KQQJG0L+FqaNb
Ls9KWkhyvstcPlIKnc8c1I/S5BJKhamxMc3XUp7XIW8/DbTXJTP5ugDlvSOGlkEO
HSCJ82dDgN8w/TWHjGTleHkLVOU8s/mLvZ6LiXb4pYzGghCr+Cn0Fq3XIKSoRMGs
y15ItJvb3kC+FbAHz9NkNRV3Ryri7L6bFHYkrT9VryafrbKu/xg6mO6cJhcd9dbg
HHKrqkBXIC6WzudL020xvkg542/YlGESLUeWy5NMvHyp4CRKjkArM3Dxsrk+HzJ5
A+ksJ/DKbEWIOaqfhu+ifnlMvnTQpwgVwd41tay6viOH7j367NDEJhL8G+WAIcjH
6ZGfUdMGGLzb+iHLD2D0dgiTMxBbz6Ex44SJmb3P2RobmgPsI846Z+Bq253gsFtA
jG1g4ZULAA8YDCdrIRyL4uknMV1MJeQL9TSidjZ60p/RcUI4jd3oo54AC4JNJnfv
YZfZRtb54GLim3X24zbqAzm5M2d6/gULN2uqVBQUuP7D9Ux3+dvLTIPhDdZyp7s1
KqeRN0KoRhGAWCyCZ7Gfmx4hqkVpO9Bre3konocBOFyFpUUVqkDBmAKiTYr1coae
H0YSGgvvYVE1jDjT5CTwRpzgOZs3+NEbMt/0KjUS+7dv2cVkhjfEU8LDOq1RiXvP
iuFZsgyID4SV3Ou007G5TBuGgNUgUzPf9zB/JDJAkGL7qowYR9YKdM/c3iXT7Zis
5MsNsjA7AwQ7I9tKqk4bMDazeSh+grvr5Vj9tfHXW+kLHrhaxOQ8fApPYs31bRi0
m3PS9NZsQN4anAEn7nWVxR4zCKhIqC3kcTsrV2UrDcQIE9LC2cp1eT/XtfecG6eW
dRuoO9HOlKS2j9rnl3gDMLbtFIyBmz08YW6mDSdJefutfELExp/WNJAlqXEiD74D
qG+miy/6+jc4IbujlAtNvjdkGG3xVvGHSSRqyi2GxhD5oHw9erDTiTY90hapzALm
XELU6D8WFfVmtn9oZgyYJ95/Jtpx7z/Ip3b2fuSxbpDnwGsWC/58GbMnJN3QlR2A
Iuljlc5L0EOZ7VwrXc4IgUK6K/Iril60yNM6dY4oAXt4yGSFSc8UwAw6vjKHyBN6
NB23h4EnjOhhC1KjHbHMcbpQYrCU/bKEW/wXSlvucJlot16CHDBIrNloH/8/I7x0
/KncMGyCW+NYGF6FDz3H03DYdOTWsgQrk5m/Kh3IcUW09UFsD0MUpGi4zspNOdyh
q6jBLYA01G/KzfVQG6JVOeszdnrY5Ui8XLnmLeNJsqB1bj8QNaR86Qou1sfm+EhH
mv58SLcCeLwJiIjzWxb1JWBeYArLtX2s6lpBf4iOV13jwTyC4WYLoTDtrsaGnB4V
RQBdVHy+WrTsyAPRZtcXsyEYbrLv7FB5WNEtVw6GHkzVjWIqfgY17WgZfr3bH2L4
+/zYNQMXYhmI5hq1cSMNyEgnGRHxjJRdJH34yFpwEydMDWQuKLMWaj+oJNF0O3n0
8v3PtO4p1jqeklfv8QvZ+425HHrAEXO2klvKAbqKMlhL1zuURJiYZGREV+o79f8U
j94VcIgHMuEIZg7xEdGOdt7WoSW2A59JFYphmq5uL1QrmhzoU1m1YV69RDpsKgix
cVFCoejJJJjODk3+zAczIBe9vERhAPoWR9KxtwyZdpBksgR7aFsKu9hDd7Zz24Qv
aOt39Dx1WFIlVZ6eT+HL3S2cAXr0Md3otSlvtFzLyJyB/8bPj9maNqiRhZay4ZDu
3JzdmeSLfF+hHMZevuOp325zA8qapJLyuLxecHWhQuRgcsWLItgWwrLGU1vPWhND
glpKHaEYW6+ioGlC8um/4amcVWWpOAB49BHK+9OCGNfCuifHWU46R06QnlfthT5F
bL7wRDUMsVeG3oDGmVqdDGr/vh4+kFJrRCPImag4co9M5BVBlAWoFHn2D7Iuvv7b
BPfswbx4Jjg/uPQwz6tAQlIt9/bv2ppCUZ8OWcN/tDsCs7ZoELgT5xypXyy7900v
QhEr2jdUcaBEIoRWqaGmB7Iklrt03+VturXNofcGVzqrFMyCK/exyw3b04hLxlIx
+i2ovkOXxS1LzyVD43pNxmRKa50Qgx/PNdnw3PMZoieGj9RILmbJp39m2jrX3SfP
27d9l+KEEt62ArLjG1BwMkx6XOAMq0QiZJrohSSFAcjOKWxHBi9o0BupQxlvN1kR
wa0WZLQYiEWGWNAfAQRNA6ZqjvXSEo6mZdn/JWM5kaBnmcVG1ey0FovXpeOyBIFN
NyJ/7mQzvYmFMIdXRPkmJBp2626CrqeIVUXGxn8N2mlZ0i46o0E9Ec4b8WBZMpET
9WBZThz4Q9xlNUKzhuPPUjACvgydHXK559f+TSth0YcLMT3w+mti4KG2UZTtkQg3
0cn1dJ6hqKFcSrJ+HthVz/ps+HgQnRUml09ooITyHtCYUxYcwsoyXtr51qHXqZWs
TsMk4FF3pMKYNyuQl/7CBs++NczxI4odiMp4ByHFBr1uS7p4kf18Fo8aPzQ5B4Nm
RjxTDmbRk/jwjlTg9mXvJYdbFob/dCbdYPhH/4MCGTTOWCIn86NR1RRxNX6g5Uav
r1uhnLXECiWa8vCjK8SMUjrCzXhriHDo/xaLi5G5cFACg2OaMwykYDxYXSthD+xf
tFXU6cgDZKCS91Z6gLnI1TdgZWKD0mCSeeej2rv7dxOrOMBB1RpO9AA1cSJM26DX
tZ6o/JGTUSMjIFjXopBW0gpiNiB5kHOtxIeE5yvImMImUpV3ZRxnU0kPabzYtp1O
s49KK6+Cw5OwkJcli8RMpv9V3XxPff64V75xrKbgfhyyqmffPqNz6pfT1R7HFU1m
XHZYdQCG5m3JRMqFiAKiM6XEAsvDZ6NxeaJ52HAT0Gntsv6EXJjJfW9mjl1yB6uj
Xoyn3OuRqUo8Dxir6uM+lHQb5UAUdylib/HHyLg+zdjzB4pw+S68vk90Dt6KUhDF
dsJ9tN1TaQU8v3lv+a85uTKa6BjwvhQVeu/zlvSSt4lJ4UUH8qOcFxtL72llNrjM
Y6XHubXz1OHZwtZ9cqEbuQTV30gffnOqLt/t8YY95kENzC2AdOcXJt5l0gXr/X5a
tmtZceiX9ltM1Mi5YLRgXh2XfgaNw1kmjWdntyg/7v/jx6po0YogaUcoYMUszxuu
VzXXCW3fPijeYvWWePGVQfbfsxdW8cl60GiXsXNJG5ge9l+6oHlRXZl3rLhHh2+h
oj3ad7RvcNtgxMCqYbYcIlPrCt29s0EhXyDH5HyoJR93jkPdtbyu7uVTcUnSTNyT
NPOHYoGtTnK98hFOo4VI6cizbCoqYqDLNuPjixvONxglNxn+eiV3XGZWt9uU0zQf
4DKmOWahAQmcKMTRuZfWOJo3W8sXDi++8g5YshZMae5MzzCc+Kp1HDKl6TeDk9cA
0Nv7ThKLqm3jCcGqw+wyMegWUYlsfs8n/1zqk/WxaF84vej3cX9cKbxgnlzcBFe2
TSyoxm71O2ty/oaphGbXAR07TUjdaPbCPfIwY8Nx1OgkUHubEpja4edm7wy/oK7t
u0aNO3hUTPO+n/aTo4JEoAeKuvGjg8NtjXTdDVi/2Gtzbp9BjEjcZCPDqjrTWpIS
6w8k3XtlAxHstLaAXk19Ct5xwLCIYDHXM4FSbe6hm2eZzp0JN2e8AmqBWDceLpeA
00ZR+301z6vyT6AgKPMi3Z3Pf95PzIkDs7knrVWXxKxB6U4an1PoqMr5r/G2To5b
L3HpfBEqYl/c8LlpbPrwvVCX+FmeY7Dl4XHtxomF8F8IrNRwz9xTyALZHP8bSWgx
a5j0ivtVeXplqDRBzdSikel2fUsmWApLgBaNZV5ZSa9zcY/WHdQzEYH1np0KSj1a
GH0blRjXd+rQaWSZl1l5JHl/g/HyxMGWQXhDnaGkhimwAb4EoxaOe6KFTCcJ/Ggo
3/5MVwUkYnkIJH2U0A+Cj/l9XXzlPwTt54/bwElNjRyjdtCqhknW+g7V1WHmWCmY
P+/T69FxHtlYoEbfrRWmYttX6Np4AJ5ijdNStUkIpv5iThuy/phshmdvlfXuW2IC
CHBQaWkssmmNEgMf0gI73umeTc93+hVaPWMXroUbGtxCL48q+W2iGAcwUjHKL6Tv
WdhG7Bu/3+Rhi0guVZA0JuVD1fGBMJIwKHZLyZetQOtZlgtsFJ7Q3gmr/FSDOeRK
ov0VfRkcSmZRhsMPPu+Ov3PtYjbPQkTN6fEuV3sKGv0r2imybNZheiuTaABzN7XV
ZhCRsFdAo4WB8mwU8IzGg6cMbWIyC5BY9lzC1g1f06e/ij/3K4ymLnJozRdmt3Kf
DDPnR/RECzrO38w83Kiwlp2eggOwVhObfF3UmM4zINmupXMiINM0sclLqLVqqd3h
1X5c6EhKB8kUBLDSFT8JXSUl0Zwe+M5QsWcQIuH+dXrRuTj9l3SL4s4XWzqioO5R
4DxhqV6MRnX1rczqvrR95/t9RU9e14fGs622BQTYZbmf0FhNMa4dFKot9nQA77+9
gHRw5EaiD57ACxoXsU0/i5K/dxk5MA/Ku9IrLGVRBmeBQDUNvO9b2qdESIAKulZz
XjoYW28blLCZLhdOGqGXVekBWDWyWQ1/B0aTZ+D8A9G0P2K0V8okVH3JvOeG14cf
xTc1izeNBaun87OQhvm53YFmrMF+L3XtBcHa2vwud9UZtX5pLzAi0MW0jtxOwdlm
kttM48nr40qy+GGd0Z9VBb01sLiLEvuzxtsdUJkrxkiAh9Wx8Pe+H+2UQml2RKJ/
OKI1B5PYvIXG8nYkYmm02APbtYlEW80XejvthENYOy1h08ygGUHjUrMwr6bMZX7t
WiDRfnMofswcAXoKo1ReWFTztaccqwN7sYmdGneNvev0icylgE56jBevzRm8ZT4C
sw1Czto+0X+WCfuocXX8gpejfjUtwbl/ihcXGp+YmlBnlWzLD8DG3+96DeC03fFv
sbPiR0zgsIBQz808+c3FB0a5CVSkaUo9GDz54MufaPHLLqWKJcBxHLPiTh8JnL/r
3PkJx93FH4UPy0KsRqHDHomcFZWEca/6dgVpIzWP9TC+8LCw+ocuuTb1hPKiXS6t
xaxbyiZ/eOGZIQtLPxVQk5RsptLBGYMfRMJSsGs+dkpQDPb3F6obk9GAXIO4GRaB
dOSwcM4O4w9895+xsugmzqwxa88hflppkNJpWpQOiy2dqKzyXdEay5Sfi3eEVb9a
fPu+4qjPNpOrFez3kAnF7c0klo3izLdt5QULzeFRWAwurFAAVI7x5bNNqbsMW7Ii
FNfVrzqN+V711cRmTUDmXBDwezLErqEgyv2bk6TsmfR9ijKQHXyq1zfxRadM6p49
G6MA25kELyRkLk3vM3LkNwSZi6bDz1Nb7rHNyGH5cm4xG4J8reyV11laEyuwWucR
N63QKcvxOFwEFzVHEYu30XJAv1V2izg3g/umPEECjpxkRTiIxL1c+dnhgoP5kUgx
JF/vtZtt/IgCUFSw03flzfNIuclL/PnJzcSbxUMgndNBlWnB/6z4T+FVqz0kzsMo
51HuF3HCJuVr6ZMVGaQU1ipUkYtkvEjvTwwV1HGDrcMJQC9JTMbM2MJsfsFXbMGT
s17UF1MTMy391vgwZvRWOd0WOwVLzPSE5ByN4yhdhjCVvE3fBvzL5CRqXOVSG1F0
4pE88FSSs4PlCB1hsoZ4hqpZjLIAOJHBvR+FfUVSfrht7Q/1Ghf4eK3JNwwQ8yn/
wLeZcFS5smEas2+xUcoC+PaSki+uVHVOocDQSODV1VzNP7ZwoNvmo1swnbDYj29A
I8XlvJgXqXcEMyAnlKA/dzKzhsMNuUn9K3tcz1kED6dV6ibiyHtqDeCZODtamYG5
H43eY56g5HZGFTND3zcxBunmFJ6nPcCi+P14PNVhge04ykj/cEP4sbpGItmqtyVi
fXVw9GyorGjUqtDyI90lw5VcJihwoNBZDm4CjCw940gd+Vht7ei9pqGiXHyxbPDJ
hFtddf+iQxWcU9PDL+t1p5bIpnAlFmGP68dRPoGoZTlsPOtderEqT3afM1EBt6+l
sX8FfLXMoJDkQC+BZSatctsBfauXp4u/3VSJcHOjntRHaxElUBsxxb+JYqUT3VEK
2ZmGn/dNc4UO1I97Ewv31pUI7nJbYGCjj7dneLjhlkCrad1XldfjBq3ihErR5D0d
l/QHC1eXt0Ed94UhwEiZhvQR9cVe5Oc4JgJpP51XYCmaGeVVWguVX6HZ8BS0zBo7
iknsZHnw01raHnBZowmD0A+I0thFpdnage+UgNj0LPWvEmnM8VbvFGrBJzfLdMYh
hxTcCaEuEMucO5fVOn4Ym65VR0eLPplbeQxWkwCu8hQbYIvQIvAKA+FauIP935VX
ad7U48wbxUPIxGnXNwQceup2tJjX9erWSgY/wYpHEfivJgPdUOhFvoyCm/mZcWuu
20BBT3Ct/BS6nf7ehfTqWiwLdyP3cYdSVCrJBiSKU6+/EXXsCqjD/7q8Jo18TJw5
wUnOTbFQI9tjg+DjojkrqZkexJmHcKsfNP+S9h2Cuv5ivPnMR8Hk5e/K2cT1Kf2l
w1kxEduofosF8wb3xqc1qgGEXmExpf1bPwUcZKAfodBhotJd26ccp0EjaekUJJAw
NV5vOPSKNQhNKj2RIh6zGnDbBjpY+yzMjDFW1mMrGN/QfwvPKAliLS8m4DwdLBZB
C/q1nKo65bcnqPVO/FoR0b1QeyhuRipiDyQz3r/mzK5HS1VhZwJ/sNiRNe3WztUT
VjtSv0dNLtgsowZA2Dsxvfe5grSODY6ww9/jSAwSswr3OR3nX5fpTlAO4e+jSqhg
H28vcxp+qas0T6OChS5xsRAu5FbPoSjHw4WB2sJSei0godvWaZtROouSgsssK3So
1+8VfDkUypkiMLtl7W77N50q+BeLsKFkwssG+y3k/x4bxI54UFobqiiMRTU8/XFB
n7/oJa8NiT3YS+ueYVUq5H6a5QCQdcoIasRvsWLnAzxngUe8DX5ls/kYOaRB8I1Z
j1bjucsQkgtHqUD6mkl32B+ODW6N4KUh5VccuTKz/FZNzllcbQ3Vu0OBtKly93WJ
0jqdNdnCgb7UASxry0WxQmsgq89piLzfcdaOOhnUr5Zj5aiscyLZ1HrNbmYJ/RfN
PeGW+CeqoSvOhvjuNhn3fUrTN3gSjFJ/cduIyVVjDiTN6WU3YJx0Lad+mrYJXDco
l2K8aNgK+EEaIiWA979xxOlyjs3vDmIWzyXDLrpiZCVIED0VDdx2guF1aHvqHqoz
a0H91zYDW4hejxAOBgHWmK9uvIEKBw/tU0jwdv1h9JL2YPqwTwSxcPZskrBmm1bE
6LFPLSQf5U90/96DEG7rTnJWxo4kkgFl3Ti2cbBKNyRBdh0yfTatBCMXDnbsb1IB
8xomJicCUcOJOBattcKL60i7NHXje58/PjK87ONFG/pQq6676gEKO8GEztgw/zsC
H2SP+G+8hJ10FaqZ1I51Qt/XKgceiaxfuLJo8gvo6RL91Rro4TRUWoz2feHp9TXP
9LiMJDoW2QoV8RBVbux3B4kzubtH56sF0huzbBiVx9UztHuxKuvnBZxZDwzeYgN+
eeUXksq4haajbI43W9bfYtVAgcFJmh3fH5HDP97vnn2UVEQuxZ34i8NAFs0D1wMX
PKAuVM9pK7ITR0hxl5Bnh4Oldk1P8IzbOUJVKSuumRJELRfC1tR/S5oA/rsfmvRS
lqDadlmLWFc6ROF9IF9GWvDrVf7jzg+8glBEghBXA0eknHw0wKTaG20X/tBCCknQ
b7yPNHiJrMSgeKWoUOL4qQXvfB0E7IyeA/mMp1j0CAPnvNC/DwAzX1bQ/Z32/142
TU6RYDtMODPXIiWDZDh1hfCCbFTK2UkxWfC//BFn/rhq+Hr053CqnIgGA2CfRu1p
hDhBvwdyUYpo/BRP7OONa/e472wuCKrgvue154GxSZun/TYj63JD56M14plA74ce
zFUM8pBVVXQ4aa6WPWDws8GrFJao33f6l/23oJhQzJQUYOj/wYicPOqY6Og3WJs4
4KIEfj7s7hgc6WvSu4O+H7SzZzVZ7ooGF8y9USj+fsHS3ByrlZ2XAhwKdldZHTX4
mREZfGE3Tkpm/XItbMz7Usfv8dNa4/Cbcp+TYP5pUGucL08cX8ehruIw4vHzxVwj
WRXWuv8qtz/hiHnMGrXLTLm0P2zwpwMkrmomGgVpLxMifhhIcblliIyAuajCpS8h
dhS8O9utw7fE6qkC+B/Ke+hzrRwTSm2COBf4GZdXssNxxGMZOUSkE3wsPOA1Ab1g
dMOkGbs23FxhYl6Dkm4lCZxRkYXwK1sOa9mlA727qa7scbajo4nQK3gdn7tkuwiO
OUDJfq23Vxrmb9VAZa9ZNs6dX7eL/Q/RBsjUsxx6vSA4b6EgqfHztrWZ82W5C2fD
uij+rsHo0JpoChPweikat/3MOKjhxI2s47b1BBZyCnYIqT3CIVWlCXFBOA6Xr8SZ
pIcP3M4nxwQDFHB5JSK5I9fUX01xx415SLOeKKbELG9e4gHnt/N5lO31NAcDBHs3
48bpghXVUxlHpJNZaMpmWEPQszwfIpbcghL+sOnqT01RuMvbYWIrsnWhevRPPxoV
CdStGfAyCL98KHWxHJn/ng0EyX7TWv3ZksnbHszzTjDR6kIby1yw8T4ZyxGdUu2R
B3SuBkkSnAuUAgOw4LgHVhJ405yGNnqEypMVPbYfZ5H3bo5aG1as80eGrrHskOfD
THWrnQuhW9VX/jxNkZkOg+3q6EMGweYYfFvKM27y9UVEt/vEercyKd+xK2xVN0l9
ThIVhdCh2QF+ncQuQfeL9pQaiZPQHra/QN0uw8iXg6DR6gb2Yx5egn66b0MVIwnj
9JvC68kRbuPFonQE87D9Ske6WAhchhQc8MD+7pv4mPMdz4xdUvliok+rusNo+MVe
LCx68MJLUteRSDhaJMfOX8QlFXnPyquFDJXLFXLYXfljw/zU8eP8r2aAiSw7NWyo
ykvDw+JS7qYYCT8ZkfZFrKBfoiM1DUKhfE8LpwD1XVzsEIYo05rVOzSQ89hZC6rz
i/frSfIqWH5geGWf7QDof4a8qByr3/odkJWq3MLhzQEdIiG3oKOJmkB7llNYTHXt
FEEXLPYByBvtda1TjS8AdXIzU6P7dQpcl4PJOfEH3EJQwPSLl8sXBNr74X0v109P
bC9fgSdd9v4T1hUnu4rEn6xAagPw8dylRi+FBzw5p7Yf30StlaCgNnf3Jrm54TRA
dEsMnWDrEN3pyoLnfQEk9J9bm9RIkd+RH4HpTLPdcKe6Q0dMlrdT1XqkHGPF0qw8
N0c1+X/yjxRzBEZrLkniac+oWBUnF1gUKxU0CFb49+eds8hfHqsYxgeoF17d8lWT
Gf0WPzI5TmHOXUc+Eq5ZMi3W85vtNk3IrfAmchxT6Q4duNcucRYiMsXV1fZ2or+M
In0LnQ8VpRCSQAcpZPEChK8ecGAupBm7eExDovpgC3s+Ncas3ruuIebOoRWlCYjg
Sc4Ybk3oYxhIhbFf6erzMLg//Q8ZYA75InI3tjw9HAwyaYclKwzsOK8SXEct3JnC
haAayceSPoS452SLw6J8DvQhKiWc5mzRW3M1OyvVATcYpQBks9mgagWzFj5ya1xl
3INuL4URf7VoYcMyanYlleVhM0WXc6VwX8dpbmhi9oIaBUQZOQBN7f2y/o58cDVF
0raI/FIRBduqRdzs2uQAnMWwqpUOfmXzp/05cbHPRkoFlyfoSC7vfIHjSTXZeMp2
Ua8w8iPYWwuZQe0On61PUret9dgd0Wjx2puQjvk+DimJKvOwj+B3G3pEuuPiBTxz
kAQF55IB2A2OOCuTQMjG8TvA2PqI7FXG8rlKtKnq4Uptml4Ou1TDPpQ8vpz3Srgh
qTFwKaWScd1ZWmChWqgraxgvnufCNVMNqNHefDpkNi9AxqFB8iTXh/7R2HZ1MDXQ
LTfW9yPr6V1ZaYAienGxZBOI+mdQGwj8DSbPeCEEscEDdyKeJbFMmaGhOpWyIunV
295ja6FzSoipmPoU0Agb/1SKK7FXiub+94iLcrQgneC6dDypTg+HK1kpyHwDbhou
rpBbVyC7uzFHM+1uys8uaONHntLN43VHdLx1rKwrZ2COmruijRDTVH0f986t8Pxb
PcOKjTZ/n0L+cYZlwPAHv0/IWruLdGgC2m3KIYcNmcXkb+Xiukow/PlX7u9bV5cn
jM/b5P8o0UQHZFn1IpBaW19OdBJbvkXEov8O5buuKoucee95xm492ouPKoj0fZmp
T0gWJ9dbMh5TywwD+haXEIL62NNbFZcgJvTAFRUTBwtaIH5/GQdvJw3IKfgRJC/L
EgqZB9JNaD2ZtJJDurOzIC+o5XnN18aWGmezL7r8vgC5BLUwCNP0FNmNWrRWdLz5
K7nTKLmLodZ26EtFH4X6hH8lSBS28s6dc72LKBmQ7b4mVPgRA5GD/0BjWCipTAB1
y5jZRL4d5ENdA9uvYeIn8QeD5oW2df8J5djUAelzVy47qvGEPZV1ypJ+FWKJkCB6
En6WSIHsubM2F5nraRUO6rHBDEByqRQXD4RGOWLGThGGv4hIbHBEfC3vFp3B7b76
JBc+2kR6HmIpsqsU/s23IOPzMmzhzzr85lh+BRm9Vvi0xcUlMRe1KblRGy6IASBf
u7eYO8yE5WCy4FpzhHA/GCC81hWh8Fi5tRWhWV6+4Q8DPc80uvLO7FHnxB11Z+3W
ADNTa1vwKmBOgri2HkVku51UuqwtJQrqNR5/6ojCPPUlZV2g3bUmp8qO2Gu3iXvG
26T8VK3ZkM8Il5JazWVtoowPMYFxZuvsvcuZmnsi/I1CxouwO+M7p3/NMuApXeK8
wZJCpDFR9C959xizAtF5ZpunBtrOv1G7P2m/3te8qPH6wyzMZsL51noudy+QmEO6
8MdIusfwISVO+CBP6PS1hpdbHevMiN+0IOtx6dmVgeDizlzpXk+VZ6PKonb07Sg1
8HJdFOLO9ugtPCBxOjBoIUcZN8P5s8mVDYMARU7iicjd2c+LwPqXNGnO1TiCNNu3
oNfw/cahD8pJ+KSuJAO6kUuNydf1jLcQDTF7D6y3WvKHUwuPZM42hszVePbH4fiB
y3CS1dticOyzpNcYk0ZUBWCwJvTujguc6Y5GxVU29butJJqsM/e4mPoioa574cdj
CefMDoJs2jvHdKiqABzkFtLgMsVGRXhOwFrh7XcJJEEy+RnXIhz0FGxIx6S5xZMQ
FBL9n251eR6f36xpMQKrYDPl5mR9/M1EONiUDSn7ZQbJu99FQxo9uQpxkvQs0YbV
m7WlA5TU32vO0cqDNLlF5im2UyGxA6xa7JS5zsYGxsakSp0pgjcIbOp3Oo4+1p+x
tjiIP1gSPEJHe92w9BcBAmayduRIt7gjTxzpGb0d9dK/JIQ0ON3pbXKk0aC01UsZ
DzKUzXqWAsnfpNekjteRE1/xSnAvGS3Y0AIa2Fmzv9mqLMM47zBflH0KPlF/mXf4
8rGs/4G7eikNuu/U/+UnN6zdXwLcav0UZSd9/2HbHXV6vCxeVwDK3azHqLuQFUOz
xQ9xPckSQwt5CogyUUBhFEiXCv+8kZxm3J4qInhzvmG8ZNMS1wbr8GIaTVJ0HE+1
s+tCHIRPQhOCZ+EeSYlL2Y3VzQqycPGEr7/UWwDfy+GGstn1m8PuJY2utT9zQiLP
znitdmfGyuozSPaE5OV3sGfuDSODUyI30LvyFKHrdATha5ZEpiNiPxfH4RthTzHL
kmORrMwsjKl6zQvMKWSJvcsYDMLqOB/6nSuEO/euBO6Jb2rQynDpvnXT5F4RWXrJ
9jXWiXWAOqQkXFvpioqCvuH3NtclthdjlxBq8DtvPVV40SNdQ6V0jrmALURJ8+1H
UZQ9EjfjmvaYJW3QJIQoFtjaTRxLhMthm9rh6+eILQTn22fr09XvmyON4YFUEaJq
KnUAWkFv3H+wAQRYtUNdL3nPtmmw0ljmsjzMTO0Sr07Y0D/DYM4pq6uwRdi6wzeU
n0YwPvQxWw/NJ3Fu/gWlY9sNAhzXKy4EJrNgpBlML7kUi8G4wsS6B2fz+34t8hO3
CQLP6hBliQKsQt4tRlQx/4MzzF346IcC2MOJNOuzHAtFeiyGAGJWblh8r8ZTCphj
FzY1OUdT5tBxtvreQDcIh2aupTAdSnTGa1u3Aw5PhkR7STRK4PZZ07LSQV05N7GT
TQly2ybuqFDF3MMot4qSlup6kdlWXtwfPK0LQ+LyOZjtqoenJ+x4jvg312qAD9/k
GhV/UI63yf/ibZdrHidP3c9S8eTjmikSLADTEl2OZDG+Xcx1tG6we6OvpyRqWiey
buW6aE5rbj+Vw3rQ5w9lT4wFpDTMmzgDLI9nkMH3Rl2R9cQiPhs6UuSlNtWGC1Vk
A4pbOGeX8q447HhuLPLyYeXCGHn61xr9vNKCt1NQvYn0ssmgGAgzRGnGinkVl6Iy
3T59ISs0t7qmO+A5KoaknQNBH+0l9aTVrpxGVdqCEgfioCIxsQLs21pXcYHZ/aj6
K7GOBo7F0fcOZHMWAeYZqCwe5chBzX/dWgJ0JXWDZmF/7nVU9lCSGrL3bI4TOtUZ
c2QRMZ4juUQiqbskw7sZzzR8VcvGqT0sRXNWKXwUKnd+ykWhG3fxqLgN9O5sO3wz
+FIG2OCWB/XuMYWtLcZpKWm6jq/dzXrS7NJoswpJ0uos4eYA5F8Otm94iZYjWDvc
bRNTdgjPIcQrvoNspRSiUcDUQYKc/GMuJkbNjXdrY4pglFZ3ypxh+mkeZMKYUr8e
drD4CtObn8xzb/Vk9j3SHqcO4BFAwEI8alXmDL3EZRM0uef+Y1oPyGMdmfuBycv2
Lv/JvflmXAqxdQP1TDr4qf7uNFUIFnSwsdF0uSpK+Y6erpzsGmQo+8Jg9HugLujT
hRl+dPUn/MOi7cgoB+SmFNhTrLph3rrcO1+V1H9vPNfnjCDv6kYTRf5aGKA4Yw6R
d9plBXSHPNwds8ZDi8tRPP95piW2UCwqIeyqPkPLjUywQzsAPkQOim5AaHeX52xU
LPo/9awNYugfM97civJjhf3ggFWkM1Veqi1iMktmzM0OFpFW85F1LvCPxAMDhFqm
O1qSIeMR/gxlhvzQPUaVudyae0kxCu8xyEJcrxzLFehaU+YnQIAtx9L/ED0cGill
xQkXjhaHU8oUvr1RI/ClrQlys5f+9iUol/xpB0dXGB1zRC+noYQOzlt7s7nzBTV8
Q19gQPkbw63yxvXQrBJObmoMVWFsZJnh5DB02Iuoew8wSKKWjPDcP4Pz4Y+MU3Px
wey4G3wXLW4vW+JuwQRfkIhhhCttkhB0IUhv4G7EHYFFyimA5QplS+WSvY+WPkiC
3YUB3oPDnHkRyzrm/HDRp6VZBaiDwAmsHyeTGm0awxFZ+puM7Rb9Qyh5bOfqqmKi
QD50WvR6F65+aQocWkfpGS7GHAkAqw/Sf2vmqsXeZac3ZvItSJOjPpudMUyyUMnB
+qxJ4C4kbiLY0We/3gJ5nSl+As8Zn8JL+TbjX82vKe4DumL5vbLYCPy/CNa6P+xD
vBUlCAN26DtdlLMqDA3Ae+OP4n6vpfEkyULUKASOByWj2yZN8dICH5NqkGV1WRYq
7L9gOpeJnnqiDEjhN1FC2GOIg8kcZT0PRDR02l9RUXv4lTax1Kk29KnZ3L4vjUdY
6ZVslpj3W22QOBOLe5SEkdeRjnXsbS3AjtGeWDWF9EPJeEHWt0S5Ai8Lsf3RAMEi
xE4Zp0De1O+qWsqvZGYgnlOcy2jwb+h9uUfuRV0dTLkCiSmQdDiROK+dPMW1yMjj
IAv5fY0d9kKJYaz1ddOOVraxL247aMX5B4bfIsRfmY94rPu0ar3aTIao6VqMHCcf
+cjhSNHqQH+xJ7iq4j/uBQVri/pPOTTXCaBHqDfFiNb2uHHO2szddAPuoqeTg9rp
WXUhfQmFfs9jdtOEjsaeQWgtx6C9qc0J40L8pE1W77SkqrC3+2oEwlu8c++7M7KX
37Ypqams8PofqSIRfUlsxr44HnsKBExZlsRZ4xfZfVwB58aaPnhOZHCQl8NfQlfP
32CAfbU9OmbBRDRSGLe7qMRa2n5btwU1KoN63vao98jEnDe0i+UWBa0r+4IZ9VaT
xoIO8bGxKykWKgvnPkxpnWYZRvATgyzXyGFE5B9zJ70jnyFpAd5S6IF+HmPVLQX0
SDBwR3CRtqdxudZCLKME1IjeMeMBU2orb7wbGqWhpl8PPB5pw8frLs8DaWCNspux
Ktq417tuEaimI2ozFNW7mQLzgRjJmhPy78mLhf0R0HdNIneQtaXWNfhlWdJDhwwe
PAaxpT7CU4FsSmW4G9819M9vv7m334CCOJ9sFs+t/XprqCHSqMgdRIm476L9SS5g
qJZzLgUnKWAz9reJLpoM/ethxrN2qiDAx5o59ySkFLTiRkgtFp5KPzk9hU2ZESVw
kOxd3F6DrlHJc02RoObjckxAXW0QjNIJxtTT36mGiTp52nmL202HWQN2035jPtW6
3/+IRkUz/Bts05PK9W/dudS6nc58igiIZC4wkuroXYoMiuQVa9vXeWwezLQknqr2
6Xt1Xi5B6MbMq1DaXxLny6yKXFZkeu/MIoibdS4/0aoHWri1dc+4RVuKtLPYU8T7
ln9S5pQnkmslt4eUU95Zd/Nd2faXjm2ErbT/T9W3rF+pIGfu28hULhSzJYUoqCdC
uDiTtD2rZdOyeFXDK+huNv7OLwXyqira7r8QsASiyTsLgbl9Z8xOFSVm01DW1R03
RW4991+krI/VH8e7yIArGg0bFNI4mCTfMmzy+3hvWmUcW0mbOcIIg4lS4qVF716p
pgq7rCTX4vDUcK1XI3d+1rc8sMpJrgLYFdB3pNjf0TTSPecEO+nUEiHSVr92HCyN
DB2VquJ1mItOgMYdKtGxXx+dSNv66svUQA5Vdpa28BgBydmCybtKj8x2TuwOo7w+
aGa3I9U7kgbG6K6h3v0nfU6SKEQCs3jj+loFN8J9yX/UrQOlRYiG08xlB1enUDK3
8hmMFfrHphwQcCRjd1KE6kyMxJMvEH4K7zp5jIqpRYCLt1LJwjYsq3FKMneDWpjA
x1eSQc/mx/b6+ukohxNe3XyGeLePnS+RUIGyVGIMmnKK/WihmDm+UFt0Ilg7D/8C
rt/4JPEKETbbu/9f9zeMnQ3JdiRJSfJFIK5zNDgEXdcl+25kSmnLYPHMtCGKh20d
6pdzmhZzoUK/gTD9Zw8C+owLLm9dbKWZ2wxcFcJrzzRQ0k9p64Jos9rd5Lrq1bJR
5fInt5ZmCxJM9l1gcTEKbgPR2qmEeacmTmdRJXflGXvt6mmEIgQRb1D1YjIRt826
K+k/scxd0jvlsK3GCizpmr3Tuh/6P3zduvU/t3DuDIq5yEY/d5ARuE+u1woiEHbv
K2of46YapR6LRlE3Vx88n2xICUVzTpTD4VuviYEFexlORyTWmcAuaiauGOCPf2D6
4GsUNIc/4mcVjEOzjuandkZrfKZc24i9+u4VaMMIYgHlmx0Sqvu+l99gMjmG9cBv
aIO4mp9W744s413oC33aRViJKsErPn0mwcLgldLrFB43d7Un7572kJF8myAfcTgX
urtyNYO/cjBOyjUJwFVgdzHsPg4x4supe/5th+nA4SAfkbcuAWfZZ6U/AHKlfyEu
hz+aMAp3LRgU/w1sm5OqXFTEcjYTnaAZiTViqPdObNZ+Nzf/w39TShQlthW3C5L5
VlAW7tf6RPOxpy0yzxTO+zRX8a9PTkMlsB23VrbsrYPFyPPrzpQv5kjkp2QFOUzJ
0pbywTD5LVLOB0DG+23QWOk2a9zQ+3UcYZRc3P8qJp5mhooPZT6RISAM8T+J/tPV
td04s7nerDsAyBKK7A5OcWkQtGIHrENyFbW+KSwFBIJZm4Vv5BuxqCNdCPlza+mE
8GmR1U8fmnkF51iOvpHuebs/pr55RIbC5x4d+zHHkKnHQWpQEJ7rI3vBZ4KjmHLK
/ro/T7ZVxFD5BmFFhqmGTWlgxsBr79S7OGkQIqlGO8Ffy48m+owNYxMFAOjq9+TA
3fzBJs5hHiqLqMZinWmMWsrArJmeWk9trT2iqKDaNVQjcov/HGkxds9Q4Dx+0ROo
9BPiR9GsAJWwJpszOhbUoGfnqvtW1bEppgiJTgppxv+xouTE0cI9tcybKqV7a6n4
Ra0Iviy6gEtP38dq9H9qp6E1lnZyGAnpaDZMS2vxq0WHrBI9RJYL/+zPvpzGhZao
c+l9JNuNagzX/bIfpZS+K4E8NnIY+0JGLDqbbHLRSBOVaWimiYuiaTjh+Ofnz+np
Bt3z9S+f/EPDt2Dda1jlXuPijeH5BybkCgwUlE9z/Z9grcWFmpmZFxzJHxbi+wk6
246YUf00L5oay6O/CSFH0a++obdFJLP12WLasPVfuEWZPNQwIWEUunEZW+yKlBeL
R4AEseqCHAmJZbN3M9YffD35NdMLfRs+PIvqaX7dTC4lqOBOmNRcjDrstFYSLQM6
Avi+MB/u2jjCqvT7GUHJRsmF/dNTFraKkbNrjRNexzVJYiUYNE3thWh7Ekknxt2t
B8069LDh1gq4K2TEDCo1s/MIms04ZPSIbI7eJQ59t6i5urBT5jsHhvykZeKuZj2y
oV2PVZkz7qCpicmhWetp/giYFS13CklgGdmL+LiO9Kk0Nx79/+qrtTlWVCol3VVg
XYSSGshxrXRPLKqcA16g+s7gyzr2gv70vcKAf1TG1BnO6LbJloVh0wS35I/7XZD2
9I9r4FnGp78p8JAABoKPMxeN13ll6z2uYv/RPpoiaqg955r6qo7Y/bZ0y7MVHoFG
5fsQLuqHQ64ZToI6wv5vvijlGJiOOGwiaOLIr9ugLg0oc7aupxY6A24Ts+QSMUq5
ImGQzjm8yobBQv47sOweF+iI3gFOpN5V5ESOzvdyUDmiJK5KfaNESs0bCk3NxnxO
95tZuW3+/iaQ8DkkzE8VyOHwSHLO6H7gNyDR3SQ8c2x8nyDbNydVXAV5Sa82rMBS
WQtNMkgMR8G8n20lYrjMwbYDCLWcpb9FvY/b528QPa2lpTPQhIRaVC4yJIdpkxfV
sY+HZQFdvlLgir1+sBMpsx1uNRXjlvKcoLR73vV3j4En3zOErSXJNmk/WN0oYKnn
oUJ/ThgBxJlBuneoHDZII2aQKgWpNxM1Krv8aAznifTcoNGOwxMbZHMEWFBIJuG0
0c3l7AfJ9J9eUjzM+SsF+x718F7tbuO+V3HEm3unzyGQjDxcbRTzPBwnQhrx7TVV
DCxjbfPBjKD00qVK7aa2B+stOi8hLTgQ9D4R4bZw5ZDb+wFzyDiH1/0knZIZo7FT
koofcBoi+E+w0RQ7mCbChf1k4ZtBZbSMdKJrV7XU4d6dMuCSygOjVcYdXNA7ZnA5
/rf4/F9GP3mLTogD/HtfrDZFcC2wlchbDKclQzJn93TL79QRu6H2UAq3A4LPVVqG
AhbTSBOdJ0sKu7sROPtmzLas9c0ovsKGPzb2cq7P/opI6SF4rKq2Pc+yzUNeNjOh
Y9WlQ+Wj+SK+js7bSbfaMyNwyuDjkUvall+eNrjdCuZYXn3c6dY2zOxLi5TxcCuQ
6etIEVPcVoIHe/m/YQciXYCUF9GPRPkNo1AEdlVHXm3NlfxcnfLTxHwsAY1tuUN4
MwtTrdF8vs7kRfO7p6Vjmnxx75zFzslCMIC3Mm2sW3xyWCxk5GsvZk3bsAfPW0pC
GKghow/aqUq/kcyWSPEiVyXKk4Sh+2AxWjYdG0Nmpk3NgxDO/AT/8WfuZ0JhGOAK
4p4RsJ6PH8OZDQmGnNC37PP9XoIG9LY9Tl0IFxTlFNEAVq0tztQrvfJ4mKnSYg2x
awfF5kqLc031Zls0yG6PTSP8KB14kJhZRAOAzIWbOerrUchLsiQdzE4mUac4G3MV
+MqBioi5G1RVmdpC+np3obM+uRPXeh1ngzuEbTWqvjncV+4k3rHTg5AsjCzNHaDZ
6gkUPt2HhHQDUKZNhwTZ9V8tqIOWyZOHMYKRtHpB7Fkaemkl2fQphAaSKR2r2Jry
vA9q8n+awEHNndYeNzNqSVHq4vmIg5krIz5//HRyF1HwTg4CkGagPYUL0FY6Hk2h
YQ/qKB9e/cBWmmeSl9NRP/66focB7+rrecOMaT3B768bewmbVuyGDy+/EXF/7sCz
vgB0lLt3dA16ltsKhGRVTwI9a6xYWmYCz7NLkQZ3cjjVIvjdswGc27Cg6uUYqOnP
JMtoJsO1hRxv9L0xRxbPeeBBQDHzR7syWOn6wUw7skFqrVuIRcinJnW+X2Q+9fOl
vFG2v76CxoLMqaQHhxZIYJEuVfGV7GjpY+x1LfV53LL7D6xhoPaE8ZyRn40KVtVZ
suy1yI1pSeIc0UbAjr7hSkM2uJ8WJZdOSFULa1j6Y6xb+NAwhSBzFKjTwjrQUmSL
oDl8Id10e+wkQUQfxpeDZr3+QL1rcWS197ojALG3Z5jxJri+RqEIXTKzxSj69ZCE
FKq9+uMcN03EFCHu379+BzmlqL0pNNAmQACUWO0rjn7AIq79mydgMqoPdD6b4OTT
tiY4jiPlRrnLbi5n3fSg8BrsKp1Yudkvs7lM8QN/IUFvWVytqi1xKS3u3sce2vL6
E9ZLKvM2vJgrNAs3eIijuWMZ2av/UDTuWnqG+DBo80CnQaV5CoSgcc5DXyTfJCAs
fRdhx817WHvgLv//uuRb7q2Vs5x7YRFDhO/Og07hQS2SjHfgHpU5teT1uKQ587Aa
de8artlG+jS6fgaJ7LltgOYkxsaAfAZy9pMbD2B8P8i6ChMJc9/AKQmn1YGhEOfG
9uxNqGvUCbnC48E800v2RJUT05kj7udp4+pj0bAKC30Rh0svEOZ+7RgfUYxC1NCn
TL9y2s2jdlRo/1OfhK2ZrENMoOgZj/L13G2Xgtw1/baraiTZWKZqd4m8k5gH2Tpj
IgCS6Uq5EOWsM8+f841aUkzWuJarZm9atsDAtl2rsgJzt/smoXQdZeuN9faPu9Vr
RwnoZkN5DzVb/gkVVdsPgFr26JNT7AZ0oKwOingoB+wnFlzAF3UgWDUOzMdkTg9u
qFei+OxviGXSG2s3elvF+1YgcAPqtCnICMgtW2jP+5fdiCFuvJn4p6+Asx/DXAGt
/wuDrInh7Cc0VBhmfZrepKNLg6CLrGfuwDUdAbMjL+7MGnr6h654tfxUOjmvgUxK
bLokVYUxxiYLZuOJ6VNQOCwgCq1jnZ9YkbU9jDR1UiuGF0hMI0zdsPK3jhLAk1ou
NU+r9pLbEzucvaa+QhWXpPljma6E95QF4+pIOVv+3RB0M0P5uKfg7edivowRzJSR
dFnUWAj3QXiWIHKbpR9mSh1riFG3pCfDRVN2shd2PpfkdfAB8usTuNv8Iz+N5+Ky
aiXISSITzSe9K40nt97jymFQe4K3R2saZzuyw4jZK9jYk2SGZ1AQT30Tzdes2lki
reIZTzbNTngCIRRyOtwyvymwCpic4sHCIFkMPgsqRCYDPQ3fGO3v0ybL6k/aLEL/
yJ18LY6+n0GzI2HNMT7BJxSxUwJq0rCQMckLlys+P0+X/rvwxLIlKLdV7tyc39MK
mmM18wBcMpbyXiPqadrOIdaBvsnG0L3CNz9niBy7TtJpLSVFvZZqtKy/fXP/B1tH
ZKyQZViAz6WxAetTAroBzkBPKwU1Jz2Ei1vJUxIeHqrv4+DyLADZ7N2CfjYksN8H
+TDr1EUU7sir7a5k1IJmIyWI6/RQZvvmtO5IzJBWH2VChzedpBkEfsb9DVCZ1tU6
Et0AnhYDzglH1WKUX1G7aflmOKCDji6SkBbIUlgblVSMPmeoKav60+ZWQE/B9VPE
BwDR8kH0fhP5L5/YO2Nvx00E/HnBOveWkcJFrdCOu8CII9Y2RuxaAOeC/SjSAi71
VmKcNIgULvSQ3OPydC25TFV3k0ylhUwDwr7SlbVDlNbCEBbYHxNUC0gTUkvez1hw
EPP4zP7rPBsNMykk5gzGo1qupoz4wjGA1NFMhp6yR6WglS6e861CyjoytoBzTBZT
OncqgrquvL1cQMc0LfsoyRUMra6CJcF06/pVT3gHpgr9La/HcvWgA4dLKkFFMVUF
gtBstG0kFktPO9DWt9d5w7Br+ODNbVcts6jVvNBkmDsrbCgLkQ+kma3sxYn7bVIf
WxX0RNB7dkh7ghDsVCwsvs8PW2QknJI5PkX9GHNelHQbcwYfz+XoJGbWKjm6M8sp
IaZX1nqfrOxfRqTHDvhxWOrHQ5X7nXqJLQtzl3h1oBEGfdKEkFs0AGu6Oo0+saE9
fOYuIY5a2/dhQlIIheXstYR8XxRaTpy0i3P2V/bVpvc1FBjk2C/PVZ1hHPrUGXFr
RcXv5uyxep1WMuA0v24nRFM1x1OuBw6DFiy+ciAFgUBK2j7HKWLxuzLcAD4dAy19
JfXa1/Ag9XbwesiCRDpg+EcIuYp9KscLlxs5aPMf4US8eLX+KYMDRTpeVSZrZlNw
UoVYLdcbYeW8w1FSUreixzKubrcJoR4wlGYbgalzZ5CfmwU4Lcw9aR25jnouWCKM
s5q5mAC3CUDXtla5SpHvz1ifmWtAc/ao/4VDnVz05RZkrt87PCi9AwTGEPf+qdrl
46hhSokx0yQnYoW4qj6TsrWPfONI/AiLOUG8WL+xHkiICeTr5Ys8Fdh2wycJe8j0
QlzAfdwqZ7YkL3rCYwhiOF2R3k0WkehFA/QSPtZaNKFsMmGXD7IgVXUsk27qKIcN
PW+eNk8LJiLsvLp56t15QXi5Rr3D0kSFTKvivfJgqYrL50Jl85dGgXb52Beh1NXL
xQDeLCOkNDjfmtPVqdpJ/R2IuRTeMaAn49ufA6AEB1YYFtfUiime2+0khf84jX9G
N789raz9b0lnfnRgERpC4MO7PkecFqKmlfnGo+RA8URD4BkPBRmAksxAOxoKVaEl
V4fOIotMI8Ra6tEUsp1TicZ7zjWXSGfCGiHrTLCj82Aa7VXoR9rQpKADEViGXRZ4
6sgo4UGn1kDUaJqxiJVsKDw+bIx0284P2T9msC0/otG2t7AT0nkhI3erUMHKJPTc
ShjQbzNpF/gG2yTC7VG8VQO41hWDMVXUTYL1GJOzT+cmS/9o+bJNcz9VvsCt2uST
35wEyMYZkxKyr+ztc0CWHuhHVMK8wt4yxwXGXlghzDYjJ+blE0cl1awU+kggKlDb
RnssDospM0C+7RcexVWMGyXWEajXQ7/BD1o0ZcC651VVkfeJ4NQqOmOqwfqiMQuG
vXhsp/YIx7IWGyVApSA2JD3ivKwb15msUfK4HmN4Xrx+yDFP4rIu4z5ZCyx2MV0V
9MRSILvD9gFRDL47SdSHfUg3J5tskz3+6J0xg4a7Ewp2Ny30nxfmF+zK7vvVW9S+
h7nHKL9mgbnSEe+dJ40fAmnMWqBWBMIR3TumvY9dQIN20DvdGmpem0A8x8Mji7+A
LMRRtfZe2qrdxVK26aygKitDJEUAyqjW0iRFAiSS3Z54zaPmaIk908KI82ch00Ae
8G2cIu0CiazCadQO+dXj0ICeZd/ex+sSK91i5y0NYsVoBupPWDQDLy4TexVX6Tfz
r+mRDvvFjizZlK2+jaC5WgjaonboFhxfT2Fo3hXU/L6L6ALCpBk15j/PW6Sq+/GA
Sdpxftye5C19/RP1WhbsOt9UkFOe7gFpELCmQZgs9whL19ldYR2Hb5wywaeZgwpq
EsoIkSQA21MJA05iKu1CNxjPwCGNl8cbQhbSEJYv1qTcQVuUKtkKgmnW+zGefZfA
t3fyosxFf1FgZB9MLtYo7rTFc8KFd3ocD/v3zNhjxEQboRJ4P2Ft6JXVAUXYlhB+
SgiZoLie8hUKW6JmEJLw9Vg+pxdJydQ81ZmF+t5MfjrAwuwut7DP9oYgOkT8Pct+
jZRO6kJ669Xx/gkfRZIi9HAC2E01xszoNNPEIbCmPDj6Z3y40btZ2iwvbFMrtJOU
buyozigc6MJ4hp5GYejyvs713EqzKU70sba3o7hJ8xf/gWhAQolCQ/WNR+l5VSyj
JJQuKWYGYgPvMhftTbwG2oVZ9YnwQd0rp1mO8t83X8clMrCBGm2H/iG8wwzyDDf2
edfxIExFgM9oj0wofI7YrR+0XiCwBK3lv/M3J9VOSD9mmTwY6gO9NNdwekbEtRmk
DSOeIpsuYKT5CoElbJALJsSB2rBUv7fdRVN19iWjpSyCO7r4uwI+mWDLPdCrWnuC
WC+++Zf0XayeaJyeJm2xqSgOpyf9Yq62Mh8y4k+fEtLQ3+fNnCfVaclKcu3jggTb
4WkKEtT4wS+c682h3oQbrXAIcc3lRrliMhNTL/yGLvx7Df+JTd8UNbLeM+Xu07pq
pLehkSyIqNdQ5lNfhMYHOp8ulocZToj4zxBfd9bDVOF0hqe1tUyp4WS3cQL3c6H9
POsZ+FEwJPlvhLov6/bxXjCG651ZiWbI/MxKDJ9BSgxMa3kPc04abiwar+QrmipO
wfhCyq6jDigL0Wp50+Va58O7RDRVNIKTPcoYponlEVFBDypqvHAzNOQoFH9ohMbE
VpSfRZkhtDX2MrKOlM2YjHfG7Dr0mbFHkJPiziDAn7MvZf1200M/8Bcn5y7nfyJi
w3QR10AQ4bC8SJ+7hwnHk6E9Hs+GUg1H96DzBoWr5jf3g+ZyuSly4jcV+GXTGHU5
svj8yXv5ABVuivb3BJ0yOvI8zvUHB95sbY+ioi5T6WqTZqLSsUYLcW4sin7J7SbW
xA9ZKa9X9SE7cDLmReOh2KFztGdFYSHTXysnBf0xU73EzddtIauxHiIspz2Iex2Y
UzDSZr3o4IKp8VaY2vHwYy0LHdhnEY6u/vHkJC3OwbBIfiFc5ifXo4xu67UhcCBO
XNaPC3LS1Du2KiO9r/8+He4/fRr1ETXBEaighT6OgmBXSdkjamwZZtKLkw50Aqzk
i/YwBESKAh0TDgL+Xx9B56wMLMtLL+ppOyV3Pv9h/Dk0Ee1WIg4Qif2odd03uy+N
3Ebr6JO8W6vfcEL6MhZOnBk8syyiwoH+rGi8xZEGWgH+4obXHHeTtShSQJGBAXeu
WUQhjr29nFPBcsbiBg+mccyjDKAqQCTGlkuK2fKr/70mQnAqXlNekVcYbJr+fPUp
O/gfhqBQwdwV6coIIQ94ZopAnllGAHUMIXUV3U1et4f1L7O9R8Ps+KXVUTgZClId
Cbi5JlciBQ2/OJFVshZ3pR+Wi1YxPxnRaMBpRSKl1UJplJrbejKSMImWfpuKV6HF
JSgrJIHnokXlXkA6xO+iRoyLQiN3QrkbEV54fDPXQX7a01HFocLTKgIigAOcmGWt
jzNjBhbo89kkh+3Ez6eut1oh3o3CzEJiLGSSWqhInedYtYdMUjKqXdTdMBYyClUN
7bU3aVrkb4SWnePermljBLQ7hcgGC5NGvbIB6jeShOncmNGjbclTrPc/gMSsrqfl
cKxElmUwOwpjgQ8H5t/0PaeM6SjTJfHnS1J5suJNMR9cl8rJrA57EEpflS0pPhlt
GZZo320/03B5vykiKNfpAoz5XjenG9zFX1L7ovzeE4kagpA1MhPg27bzh6eQ3PRN
c7UPbWyKABxHR7cNdGLI/2SR4ioJGsn9ntq7gW7QJgj6ATWEpKUukW1Di1rmJVdB
`protect end_protected