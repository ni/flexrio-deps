`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1712 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
5ebVVNMyfxIGIoeonR7K2xe5BAnQh0GQpMvAifjrCMJgg/6tZ45E6cb1qCBdghoy
4RyfAFfaOJZpgqFv7bdAIOFs6C84ubikROIbkByj6FkJh5j6ZGaBF7v38FnlHCTl
iuidkz03oBePjoUEAMXAyh3XZUlH98C9YJfUgW6K1Fcvis+VQJbwO1VkWIi8viPA
/4YUP0A6qKJgo6WBxddz+PLii3jQshRWexluLSy+y6mHKqNhQKHwO10EdyQvSwkQ
mRW2I7+dHkCezUNAGF7WUTAqU0IO7IqNj+w3ZovOF6+JtXFhVjhB+r+UY6FlS1FB
5DyyqXpWnuIOFoPC8mjasXhsZdrgRr8lJC3lg1su39p97bohQqAel+io4z6PDWtJ
FVVV8sYyPlar7Jy9l2BQVNSCtnjon0EZJ+5UfEU2efTWb7dNPIAEajkrtclBnKa9
T5KWewpro2z2VvvxKrsrcO8mL7aG/30TQhPfYMCAc69nqGoaeyPillLuBRd56GOv
YQqH3sqdGaP1AAI3ELmNNAgAlrfbH6kI9kA1G9ZwLM91hY7iSYkPd35A8hCogEqe
9b1GF7EeiNqJKlIey0DvvFHSW3rIRA4mme9XR69B8k+dtdDKgRUNv/U/S4QnnevF
fLk6YMYxAKxVX7JYXRR2v5Th5DRaCY75EzKO4u62ao+IEeEfeYHfRnf86YInhckc
6VjdTNS5v5VmaTIt+IIWVhsW4/Ndztam8vXZ6uyjzoivHpIw+2jAY9Tbo/ZTM1tg
zAzCjurNpAOHSiiWNbWA20+DNqBSOFLY1eIIDyq2ARrrPpnt9llWxqit5+KzNnpA
OQijCVJpCYKYrepFXOOZA2WYpWCsA459ZH1/YK3KMZiF2jrIogKZcvrH2WaTcy5J
eZvlgtTPAvCdQTcEkbawFLEjCp1eeUTn8RIKLcn/bJeyw/nfW7ALC9A3EN3iNMTf
Ql68Cb5uffHd3Vx7nMPzQd3vMs8tezTReF+HFHXLRdIVEk6aL0DiMTXIEpzxYed8
lAaFgHUMrkd3DDd93AWt5Z9b3/A2oQHmrIipQqdMDSU3uMWlQUBJP2tmG7RGfip0
pOuiPMPJbZ0zMiT3crY7LULll+Xosd6HuAYzKre+91Du97qyovAMeajBXCODoopq
OVWugtXZmuV1hnMjqOM7zZ6/yAENXYvve/om9Ybp2KEh/AhrmqAiYY9jhR+bJJx/
g4jucijzsG5FTsozdgIhcjbCk9te3PrjO+UHmrdpRUj2Zi2zcdb8QS9bzMdBfaqn
5g+KvlbKZsD7pX4w41xRcunBI/APlfgnGrusOnbs8qEU+LUhs62JeFGMwp+DXRUw
7GqFZM5BrnDz5BRPtrrwm3kbL1N8njGrs2y/nAo8t7cPC1Mh/4kNQ6S4PEICmDZk
3KFz9fRvk3qNE0EzM128H/4LRX9FD35bCuQFg5nQY6vbnc2zMCHdLJ+1XT5hFgzx
u/j8eyv3XsjzJhm0PbyeicEn4OEMBi2turzTG5dx6h1QvxRzfZM33pMTa8flwfQ2
N4rMiCwkiR1NjzqiBgDYlF8XRXk5hSkKAtki0K03ooGe2XlIQYVs8QgJpNu0vEGc
MQMmd2k3N8Q0Kld2+lGvTfFyKqrTVQOfalWmvmrNPDKk6DhZX28EnQVXn5/POsLr
/ntTnvdAgqaFBU3MAV1VpLcjuwOtSDU/PaSuZqdnmVU0aTy6KH07aPPVx9bjFSTG
wmifliPSQi4zyJ6+Vi8OUhvcbqRYWIIcpxfeNKrb9HWidyFtTRkXvfaD5rVOWSqx
ATxLMgTS4bAIIOwjYzvMladbVWjDbTR7XLsD8BQ94e+tJitr04vY3UkbZY+bFJgu
vDo9Ir8s1+L5d1LwV+i1klJPbu8Cwi3FiW3Hu8WDcwGT3Y4kkjUO/XKdiRnlqIb/
MJU18v7zu+47KoJPj4QutSDjsTTVaCfYt9UqsJUc7ryv5LLtzAGSGFq7wpF5fQDX
5zep+V6A9hIwhs35lKFO0FBX09mp3nIvuFiTFCMTvbvuV6Eb0phhBNYyP/GYflUm
RYIY5Zayp37cAxU4Vknrk/D7zqQmmMflEoSWRX2acFJ4HktyXskx41IfeBbzuuTy
AxTNQCbFCk3m+GGexi3QtfWVC/lEDJgpSWThSLJpKSU=
`protect end_protected