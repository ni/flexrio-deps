`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 38064 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMWORzZC7bo0toZS2Zods6Xs
yljw+BvqICQb54hGe2JGpPYo3VgESEVZQaDRGtsOk3QfG+9rBbVoC/WnZktuLDM+
GgbbslJQu7WCQWv1H7l1xPpzuPG/1+gk0fgyVZ0ro71Lt9YvzrQ9QlaG51MCtgB/
qwv/G9Egll4nw4/phuTg1vJje0dOEG9aPA++4/FSCa+0xU8ZUPL1wtJIh9GAzXQP
ssOhGmJvd/Y3C7/Ffv+ecJLx153pNXZwbdt2vCjxRuX2a7r2VbHOxcHBB7FMMVfM
Mfxni6p+RQzyPaN612KrvLrcv068ISSrNi17VZtWq9E2jwbTJMY3S8qR8mCwhJc9
qsayH3+w1irNOjVfQKMgl55thPd5uYjzZLh1+3gf7iapOxUAI32BPNgWczbGBqxo
nlcLDKafKF/N8M4CH3O2wTr3uJL9o/yc1f8y8nv0HOC17ZLjObomJ78y/gc3/WZ3
RFKjdjQAZM7zpU78+VFwzqWSKVQ8RMxveEE4DcWBpZeS33TujO9Y9nP6LxhxmymT
grGfGntMNShsFMIsLPjZKQDTq0DWmgIoxJ9BhQoddCvG0deE/LKhQNzrp4lahmbF
gKx82s3P7IQ0BPIKm+saVp4dnod3JDiQvx1xfnEyzsAhYJmRVGGKddY5RANAyT0r
O03Lvq6ulDDb9nPNu6Lu0pPwRpFgozI+1us0QhrfLB9Ln4W/3NNooC20LtXIsnKV
IBryJBt/VMQT/6tE3MmUI7MtKJAwUfXLTXGgxgsbNjEI3kcGTR4lkq6m60x+W06/
WHPEAXrMfCA598cUihGHmdshXi2wMDmakDkbuGiPjp1iJ4wZbHsVS4jgzSVASW4m
sVR2LimgQByCG6Fq5pNGY9kuUf/RT7Azr+22xrGgq0GBNM3rFrIdY8d9iy4h/ip6
IFq29Nr6FQlRMwJfvRrckYunDc9fb8EsuZTooIYNevEENkpuearearneQJnqbKeB
dW6KCnVE3i1q1+Koc+gMKOeWdG3JGohNV40oULd/hXALWcjEQB+zh3/fxEA+XAif
4cUsKtYniQGpcE8c1Wa+YbS8wQUBNzWfVmMyFPYnvbPxZPYIutcmR7X3L4vhhlE5
jNrcZ9NDhJnIH84Hurdqepl8rUron99yOTVoDMYejOka3QDEjfHxF5ssTy9PZxT2
l5/Bhm4xnnDtF7cEqrQFj5MexNi2z/lnXN+iHDptBjFiG3C8xvl/Fy6xW//BQhLP
/7yiHOMcaLFYpTBl+cJcV2ea3OxNxMaybrO8voiholK7FHk0JYIjN9FLgLYTztVD
t/icYcQkHfOFbZ+jf8Re3OYUHmvf94XH0f6XPW4UOM7V42Z5ATeKpkuMPLeDr9fW
eTF0vss6Usvulh3NBjeZifyU/+Yf0DSbB5ktW2ecWczDZVqwrtTvPT2jK+AUEyRX
xwe+FGwDaVkKvb8QUIBlhVLMJIRdawFfIbPnby9lS3z6wn50dturC+MabI7c2clQ
DqW9t6Q4HbMh+Hz+T7gVlp2ItI3oc8Rx4uJUZ+SZFHni7CHvrM0G0INvDwcB4tjV
QRVj+33KWur39jcofvX0/G7Js/q3RMaa48DoEYDjPGdrj52EZvbbSydAAB2k6Lw1
ehd15QBtti4H3H8y48amODcOMaFb6Oh13Qe+uB/DzWpHKFfETEMV+W8Us4AP4j+J
D4HEPG2x1RxsKIiJ/ZPLei6I4/3/d42fi6zBJGEwmbp21t7BsIXDrwsky//pt94D
WTUQbj68Pb9x0Vqj4rZWY04sw41iA4kZFisKPGDGqzU2+0XsJ/SX3u9Ba4w50Kp5
s/7q/B72dliQVjhQvqA/uxa6oSIABeXjvn49nqlv8WcfudKT7i9IT4qQYdffsTmb
+2bYI1pIcRCV45s7ekLCkXqWvpnfLds8XU5Q3FXR5y+aH7oZnDKLw9SwLTE/IWKb
6Y/F83sJLWU9sDUIyVdIQjPkpVMcgwQp2q/HEXGXbmvVUrQV8JEiaWeb+zDtFzuC
FlcT2d1707RWKSzMXnW2GS1DCZkceF1DzWYqGTBaWyv6Yt+vCrpsIujONFms4XYz
cYWAjYK2z1shkg3sHTqoBpTXzcEMrKQKtUTa3ydRQddVyOGzrAAnfxlcp8ZL7Vs9
TL3xELcJIMmS+SM642ntPzuUZTrnE90TyDjfovRqs+DuyTQWUUjFyUHM0g4DIXvA
w5R0Eb9aznjLVVmokmiyqM6fWbfr7sGZZBrWGdOOnqnYITvjdvIXyMjShad/W9K0
mqBgJGAHoIZ9aRPt8/fS5bg2iZzIyNvfVS1q2WOyl5JIa7qH1PhZ5GX1JLXWWQO0
uB1qxaalU2WryUuAHrmZytm//KgCpDH+zQVwv6/RvBxnrvQXKM9pdGtftCFaf/qU
Sl3P9i5n8Esiiox/kKpZUY2itMrJFV6CBti/kGu87DskOYwjv+ro43trtlEE8peh
35HEVZ3KaCtDHQPxdGOAfeXQM35io6zwgeo6QgZHsHFOKHBMWzXdebOW4wigPU40
R7Tp3PYjpxqvHGMtkTOGX8Hq0hWdvg93+0+OHh8IenPi9vscdGMYIyVaR/7geLqY
pcSmTRHBCDfALlAS705mIHtmOBkldDRedUtzdxOmqfdNFAAc7xEOt9zDVeGggerR
QpG60TKKPdCK/Ov3G2Ao8Yhpb0/X8UfPDZy7LSEz3QOOjwcV+VaUgWyxzp5PJeVW
zQXtkP/q+uZg/sqHzADtrXCFE5QSmszdLyoe+Yyc93tVNhcNNyfJ3Nc3q5skMkzP
c9sB4hgKNQ3DL8J7FAIquBDlEBzuOEi3BUbkurq+8tYIpD2TlMj1nFq7xGPYjNfx
2I+C7li16U2Q2DH9MZur1sQLx77R0doV6MAEwZigalF2mN/h1IwaiePAkxD0LFAp
VpZAynK0U4aMxCmkksii81gbw73DwqmBNbf4oo8dkTqHqCTdADXjrkupI9UxCHkc
zbuRY9tcvJWGayKA3PK6ITT2ULDWeaLcncyDW/J4UQuVmrb+OQqO8nScpt4vutaK
hAuYKWFZC9wYBtymBmuxDxiHdp7SGB+2uETJmNrhZzjayQR6V98Yf+NbyDUMXs1I
9db39iN8HWilzIrYazd1UY/i8EtbGczGGufKOu97ibqu8NMZzcR42w3j6C7D/n9d
xo2zfud3VkN+1/jxwldZ9n4DZ3VxfY+jIFZGHy8ppdS9000nb3KjlZKjWjmPl5Lu
hCAO00oDl7vgDgJqBWx6Ji/j9CnP9eK+4T5yKTIL56YrlB29LMqBUpkwUrhgSDnv
ob5A56j4llagGRXau34opeaLPcsCWwndezxHYLksCzAW6VlD1DCbdutTiNZiHqzm
IJ3rMXplVz3BT3d3diqI3vg/jwivid8F4dkgGTzqmtUmayb4ODNxTAVaCrLm1Tn2
kWBTX6gBaoRCvbnbMlIJNtWNaduYsicEw3oNiq9gRR/A+JIW551um9F2hThKhMCF
xfQR+ZBeVs9eNwvLZf9VMG1uYVJ/HCQrY94OPuftSzPuuQaqkZZ5GjIiJVfwwWbz
VP62O8IROx33OKe6SObukQCuAYlKoppNJqksJOd1WdKJK0Ygq3XzpOK/OYvuM7j2
a3Ic/NHEwqfXfRE0HRmaowzr14Luoeh4i0wAmrlSiOnZympa4Hlo6YT5kbmROq5f
z17c44jkZtuMQE19fVOGeZBsfIkALAypuSweFy7oxtlJbEa9hh6wrmHjwXP/9s8+
W5KwPCMpPdNkvnnYGuTwOUa6vGANlhgJalEUnQElCqCzN4cbzE121pFA/mxI0rPD
dbQB4Ng7d99+W+ZCRk5Fz924PvczeaTYVoEe2I/p4f+UfRx2tboJ16s+cLyVJBEd
Xtu6QHOtGsH+9twzKqNfjxZ7lky2bzusQvO4fCMREtMM2X9InIFNFeNhCE6CZfM3
VIE17qh5M//BtwpfSVbxfgPV+HhXOveFWL8t+5US4lX0CYIn89KpyqdpAccIOA2N
RAVJYppmz1lLwkrKKNVBORJjBMhSZFQsZnLKzBsTkQL7XoIx93oZS04RINtUCWnb
4qcEd8ZxqbaNbAKGn8CEz3xiH0bkSe4WpFjEf5lRj6tiJw6i4BY3+/u1G6uU+X18
+N4XJGY/5LPTq8BJnkX/2Y7vEWTVgDMawUjnNmPLPik/akwbzL0N9NDY8sDYuWvr
UMod+q4R3rI7XC6/hPXAoqvVnU3pT6tdv5YRdS7+xLss+vCfG4xdyIw1rqI7hfVx
MXQnE7BBV25tXiBUlNLStiQ/vPnpWtKBPBWiDhlvaXhgm/450y7RJOw9ECHh3i8S
6hOKDRe486a0kdOsj2uVJNw5rUzUFP1Wg/Xg7lrLu//f3TjYwSsv2m5mUqyZ59LP
SaEIzncEoGPYtTrnxFaBXQaCZeQkD5Gb/HS4Nx0zmMzXR3M5z9fXCRh8QE21A60i
1aouaaWCl0tqMZah4xJ0dCHSTLIQk/P0d9VxWCZ8WgFyAD5EyPB25bVqyogpdwak
BHktOfmQJl23PPisKOFySYwdOS7mxEpCw/4a0hF1LzYemGBJYcpQa5FhQIgLHpYo
D28gf4ouG5YUL6cXtc6pUGumOEoyDD+y4KBL3sdFR2AUpwYYeIJt9Wr0PYoUVdZh
ZE6i1Cv4jxdLfD/vYBlb1/1G8FYWHmtQOm2sVz/GOMl5I6s2gMDIjGStHZuoKhZJ
oEHva0Mz62giIfikzQSRtLNT9p472pUpaYiqedmUkELgN6KMg3phShVTa41kdZtZ
mrIRvCojfYcRpdxXD+bO4ZnBGib8mgPXd3QhyU/yqu+yMYeJd4XrVKfR5QgIjztJ
D4yAnzcgtXqpwdXjhwYzbO0QQCCj0Y2k99HOcUGNI8yy+T58CTW7kN5KMeK+++e/
PVbBqOM1Jviy2whyKexdbHzngvN3E7j+5MaaOnTy3mUpMF5gZpOX52AXWJANfLMV
RNViex3oSq7krMXFedQ+Fry3R9xaER+RV+/PBDv2JIrrargPGAltqgbG9slmma6F
lCVUaBDt7jMOnIC2LXY7LOZl8xA82lWAx23KLR2ArBDPJO6nJhFIFlBxcSPXQTTt
CtnYjCcza9iQ5MuWVPV3nbQUiZnrByGPrvqESPgksJol8Nc1qu3WJINBysSMN8dc
z/yzVEesi5O4DUaKrcP9BXDkSvPeAz3O6Yj2MXScEFxtI1bG1ZGQ+j+tjvptL0kJ
bL7wWnumkhEjM/zg0a/WuILAsXEL8N1+bML0Z++h/2Gg97qGdg6NJm4F4BdoMBZy
boUQO3VOXtzmp8+fMYfzcntnRT50xK3yDMmGxThiZDLnkpMgXfUIiMhwRt6iHkui
9kG9TVhSKUmEhAxhVMpm2tPTfR/4IkxecRjv/yFXAavtnZ8EPQrB+cCP4vbAakmo
l8BvRWgC+paZtbDtQm0EPsTo2bYyiDEawfYyQUi6py2z0KsefFIKPVpa1LvBWyPo
qMxUB0xbgNxCxJQK/8/wpZk36RThB3ZvqvQjSwi459U3M3KMXvRNyyL+QOVHnYFA
irTAAyvGd4Or18R7HH/w2gqIcdZkmkV+lfYdfw6KquOb44E9jIabHCmkQKrZEus5
nRJgqCu3wpV0sUg9ZHTTmPWE8cCR/yoCXUkQE8gXmLU1WFzKmGhAFlL0sXrYKpfN
FWw1PiPyJRG519lAInfMeUbq9JQtImd9Qda+L0KRIWuLnF6DPArSA4fMt+Bcqufu
Zrg49v4miUovjYYE78nQmajyDqAaPQbPXXk/N1n1p2ouwJJeLtVWV7H7Y6ZbRVlp
QrPk/wQOFUjImQz5KX4Y75eCnu/yu6OVTWDN69eMEF4FxiIcB7J+/4t3WfrGW7C2
BvdhWXz/Lq5Bip3LTzAZnGXuGgKnw4pm1GPJmGxSQPGubuubdAvAgvQNu0ELbwuc
XoEsyUzNbY8IAxMVLykw3PYfTz2wapKzR61ROuEf37/H29UIEpxnya4kKaz1JKZf
8dHhNjc3+PwapXqJhHt7z5lTdYj46dBWFBUzpZ1j+5fEnWUUWSUStR02WrxTHhjz
pEkO9VJQ6WX0ES8hOvKMP5evM2yhmIWEkbvTaXI/z1m9znWcWH3F0jPG6EEqNtRQ
j5hTxu21iysjx1t1ZbImni1Ty+rUWQjxNH9qOTI0XZnzTggkSwcp0FgjIRPJ60G6
V1YBkJBF7vkC0oYlzZFL/IAA34uWg8IPX3nRYFHs28UcdAs+P/1ObrE/ruaiYju6
wsK3SOJBGsElRRQ4J63amhUN7FceDv/ICH0++UDGnwySt4oiun2s45HCMP3dTycj
Tp0+oA1wlPdh235FHnlFneC8hxiHGxtPsQy16BsPcrlroUrF1Kc5IvxfDeE9/ZuN
6kvDKtYWeE555L9pek6VkmdtIuBaG0Wz7yzQjfynhYsYva+dxSXOE1OuA5rup79l
dG9degaYv3+WpyRm0qsUfU/JrD1mW/Tn3fFKZQXEbG3JGOLaNBcdffJi/wAJpfVr
7CN+wJzD3llrklC+Z3EMm+TvLgsGbWlK+0F4n6SMHJSwV8rfN7CoYlxot5dD1kb1
9e2LZu6JP1A1dJ+ITh9pF6OLqINeTpXieuCTLj0CXOMiKRBbrbO+fZt8hBkkjwSN
nut2G7B9FId3Ok3MqC1ktWWT2Qhv5gbC43GvVh3lcUQAI2ij53+9wYrSkWvMTnr/
+F7jUGwlkcJmGoDhXVFSjodmU/j2tztpSZVV7XPOVyLvZh6s8TC8IVVFqx1g/8Zn
HDArPsbA11tsuEgsG6iR5RdH1CX0JhlVCzOEKZbdHj362lNO7OkU6eS940hvu2eN
fCPUAa+LNuXNI8C8zARIpEFKERxNoZrAyIDWhvhlTtZeZHTkLLpoBzCm/al+deWq
S4qx+g+yOqLGhBzs/+HsU6YBNQt7QIZ8RB0EnF+0GGTjDGmmk+EtlBv8wRiv1Zv8
17iuSsg2XWRsyEKyB1+OsD+POcDUPZf3T5AMKi1Z0072tZRMf7J1lIN9yo1lojaq
/XtQ6v8vpxXgPYStH+CB16T3rI0GNBWDPX8hQBvIVkXZg0bt45QKEYHf1HzBLqt8
AWlJtXki65u53S09wNxIcBJnlB1imXBVwojKLeQdZcm8Ciz0mYDmkwNl9nbOKeql
GQ5NXTt7R3ldNwLGfurPngAgSc0WzfCjWkwU8Szzkzn2A2ZuewZqIvGy+alynZ5M
rjR20RjLuSFzPrwcNjQRF9iKc5sCfexWKVvlYXOks+msq8Nh+WLJWagpSBxR6F1h
oJBeQKiIQJahU9b/tnsM7OTuNo7ctEdmKeTKv5gjcYmmzJ8g5k9/PCYTESpPYG/6
QHe90wCZvGxIQ2UC9htHVyLeBCZ/lnhvGvyMng5i9tN1dPR7tmbLv59OqzAfbIBQ
NQu9Fs0Y3FGwLmuFWy3NGeEp+79fOKyc2rp4EMjWPmZ9f4aXWiIR+3y+8PQlBzCX
jnkmUivyXCetQvTuN2frQG9HOvtQN3ggqJ/Hf3OsxW86DNPrpoAjGU2ZB19hGDNl
BcnnM+J6Xs05DKX3mNOvBrPB3uPB+oCFDApE0HovGe+RjE+wMDReB8aB5c8DY0+8
ZdbaBw5b62/UtA/Ey5i/nWRIUDE229Z8ZoxwK4gFY58BZ1YGCSdTK6EcAxqs4gkI
dMDV+9NsGSM6vixYy0N7Umu1CcgGALCMX32yvhdDUJB0yEpxg5voQ66p+CZRs9un
euKdsQbpzhz/kPCg9plZjkPruvP1WNVpTYUCnLy/20JxqnuBWDNHIDK9llgmFkR9
6YP6t+AvYxzSQs4OIagk2VV5mMT+0DEbpNuRwfT7p93UXkmE9JhDyLRQ8A3Tkm3L
CX5lU0XodN7GAQQLBrB5ifAIEmvdz640Y7kIR4Eoucd4gAc94P8Qyx/q3J5OADHf
KH3IHZsPsYBHB0fhkPUyO6qte7ze3SG28WCWXJO4m2Cf7ySgSGCkRHwQikjFqIST
JbjR18RDJKWfEZQueu0XTkmJa+2e5iJrc4gTgbjUy4EZUoeVwV940DYg1BGoOXI+
Ziiuebrcv+u2Q5baACuL/+Qdf1Ksfa2WlMRYY0baaDP/xtBUOLwnL4YFkcH3vODA
8twA5hnmdiXDjsG/i8jOTOAF6L6B96yMKKXtVmF0rfRflWd3gRWDgY5uYx2L4iLk
zjS0tboCrc1T0pTlnMxDc8fKlu6QWZylENqV+Rk5oW2npnxiBa7sKAjbMw6RkQnV
lRqqSYixhsVB+IEEMWvprSZjIGr0fRQaQGSr6RfOB4PnlOAM/D8dlM9pf1fSwjby
Z5ZgYJCMNeApB4Hs/ZX99gDVsQTz0oT50TaEFVbcdIg1fkli0K2ZIAdyVpHDj577
b20tEgsG1FJRICOFU0lAW/tqrQMN4mAqmJg+4ngZuHtdE3wsGpVR1YX0Je0NM3Um
edK751y3LokA+PQzqn3uSFXf59nVfQxjd/RThjPp8AAgX+SXbIQOWT9XH6y4w8XR
h+nuHmRs0LjxiDhRSuVCW0C1+O5eRgnN7EScqF85DcUrH+Mu7ZZNiCzn8W9q3WXZ
QdYb8sRSn3XDNDwHhR+wixuAl3g07mezm0DEYC+hPs9Vif2VCFkk/B4Y8wYcWQqE
KmLHyiTT5dKy451yZOI10VOuqqurYhJcpQxTiqYZyIIsqIrxnCIXanpEdKfMGMS6
klx0wOUbNhdM2nBE2izdU0eYE/BNYThSQPckvQkpgc3vQ3/90zvu0DJRnE0rA0yD
ZwZz/CU8VCZoUblEf8QAryuD/OE5LgfFzYfyeiwLs5ERBrkTRftFArwThFvuCQ5Q
M8zRAGQBbtRJBLURuvOr0YyRgu8fAWIHTL7SSWPTYJq6g4lPvZcSeQOyoEacSKL/
MtL9su8oS8uxAWfqUwjerJ0SpZYIlJgaYfHTZwLIEkqfm5VIChHjWsnQhnbcPBT7
AalHBuThl6DuA7ZSnQ+eh6jO0U5fk9DFBdH3c86HY0tWdZr0sShpOrknJScecYtp
2qOjCHQuxl9F4zakCvvliSjcw0tUx46pA1E/c2zdBaLh/GRJvZYdR30YQM0yr0ko
2xqU/Lpu1GC42xVaCrmIXct9ZcM/zCHe8tqIxmtehNrZAMasGAZOlbw0AefSZS5j
TqXdxX0ET7Rnmqh+TNoWTq8e+aqiRA63PnjTDP3mY8I8zTISSDfofvC6yu6ey739
sNbIbiwqGJ0jllMtqHEKXQKM0zkLWBOGoGrt3+YEp6PyAvJcN8DxmX0Xr1awLt9B
qsNgbM4DVyIU0BOaoSo783XL1bXMSSSbIO4VBe6SD0VwKENBKkNIhuS+Fu0aQoSx
842c6vD5jKHWtrycndxFQKyuuUiGmVJllnMcnQ4wOTskc4krZc4tmnGvah3PDsYl
VEImWnb5r8LtLYD6T/wmqklpKvog1y0y0omBSzQnm9wUErFvMslMVI18/hzIHSY8
nFsg10oVHY2mF9cPT+yIt89Cw5upqVffWuE6KDmYDH3daSrQyUTG3D7iOgSZBkSb
Fd+Rn+MNKoh7ipx3OVMOxXO3Fs6BdZMJWpx5FsIechLDvUUQpHPOjfLM64wFqBcO
usOqYyzdxKKZ9T06p3Ox4ntys0aCMBixAViYt/KbhS0P6Cwa2lixpFZkcZe+PQqg
vnkm7u5+8XxlnNwRX6UosVsBZ4W7TuYtAgzKwXnm9vs4nydR53D2nCd1o38IqQ3J
Weyw6H9mxJZig0dS+sgFuCUT4OkzFmR3sixA9z0Oqd1SrXKLFoS4YKL6OzBOoZRt
9eUHhae4fIVidgDd9BmKgLPQ3MGl5VdWycxC+bbespMS66JGyPoHLz2cQ9x1W5OL
/OJ1NTrB8ApHKu0ytw88uIXsI3S1yuvUpERDI4JFf+1wsaOTwkEFBqn69C2fZ7ZH
B37OhfY5QSk+qZZtMZgRudJDGyAmvBg/dqDIRz7tb7dFufZBUd0yedTE1inZcwT0
/4VOX5LHqzaBUEYX4dMFhIZ7WKtHDAK7hcQMBLWcMeo60IS43FuQY2lcPgjH+cfX
3xAWH8iJzyDDDWh55WCXTmnGnsvS2VzntTzY7FrdFMXLqc3riYGWzC+FNtRjluVS
Wf7MkYHkImchE8VDySBuI1Rz0s5wF54rfaDaJNeSTydM1LbIJAk/rN89f/VprcmT
setkULRLcbmfxoxzXX7Qo0PS2zFeMMtc5gHt96zvtLpgjeZkZsGL3vOv3HT+Wxah
1R7g2dljTXE6zlpzWnehb5HQojxh7aQSrZR8bhetMprqcI6WA1LC+yO5lgRnLdWn
P5UuDdEuQ8wNOiUUSHYdfDbhkZ7o1NIAhbHggVyVv/XATSPwW/oDY/BFieLfc81U
dE74nscwYoy1OF9yI5xucNiKUetOUIa9yqV8VoA0cso3TjxzY9cQWqR2pOSSuGNn
plDqevOYUJoyV+fGz15IbtnjmNxewQGwlmGOM2GhZWBayVdjZyRJsbDEnP55QsRD
pYwRKaZR5Ap2dqshAB9jc7oK4nvmjeTgxTXd3+6rxbjQ4eNeMwb0PDxySyltv+XW
8isYKfuM5o3tbLsOSXmmmEmpcsoGOgD2zGezTqtCd5plFe+pRrqizeJDnR7kklED
44ZNzscSfWb8vG7kXlnzlpiN3MGlh99xOicl7lLnFfgUxRzM8sCPDP+AEURJa8qX
pOVR9B9aVJ6WQBVgmIxV31YWuHcTiDyC1LnrX1p3Blnu0HBgzg4D4DvDsyEgN27F
1YNraR9ECAfkKRnQuSno+XUgCd+9o9Cc2DT9DE29TO0wThH6Ot52YeUIs1QD36Jw
mp8QHL2CnIFyr6wq2MUltEsbh8TJdDKpgnm7RFDvCI72h4F9GRpDbZT+58C8220d
LbO18gA2kA9i4fKIFj2gg3Qq371dON5UJ3CAFfiSIH24dDrFEKmxcyaQ9njjAyOW
gy+JM+x6zKqSnL8AH55JKh300+QNlrhXf9P41cVILEU7FoSClrP0Pjm+kA1PM2U6
RaKdEVtHX1wLcMb5UKgX5QKMRk9z3VgeUvxbDS4YN9g/W9vDw9/HtX422FLcZ17A
Vh2lcboClrnAj8nqoCETEjgZHhB+PHNCqqlnkjFhtfPvKqJQq2uPyaQ6WTagqKt0
VZSKyxmj8us5wTaOFyfCZr+kjvvdH5whH6mrKZYx8ELDLh3SNnMfbRk/BwT5Sjk3
7U0P5lKVmGaIjl3XdNBAwi4guOmod19VJh7TNYgTFovzSYut8rVIlyMc5lR+MeOV
2kwepuWzbUkSWpdEqBxcvep7zVYd2CfDRAVVWqHo9uJr01FsCPRb0hEaNQ4aZGc0
BC39nowEHj5fa7VHQAdFTwuwJVUh/ZCSu2znIu7DDgptGEnlDWJ00q7KwuOErwbJ
hUN27eiUXNdlUx+ybeJ5v/lTAcNCWJUPWfBKn+Id5cIL/viJk9zYvTRTWkZ8iXdY
uYcKah5rW1b0LXc37rlWWdTmdWYvb1fS2ogWWGI9q6FBdJuCqAlV0aXEFi9xH99V
TXG9ccn+CxtXPVmAHQtF0SLqNDGJC8WoJ1pyvAoWxyhGrZW6qZHKeCER0Ka+5cCY
YOtYtvIPPmu1sm16DV8EZgalif4afgdpvHC9hdwm7qpe6mdReicZ+bCljqvt5OBG
yy/fU08aOZbgxc8JdCjx/kDeVOicWTHGI/n2+REy3xBv9S3DrTuEDFJxNOZ2yJje
zB2v+a2bj9i6rj7Ah1rcTpVy5tiE57LOGHMgKHc5QpBt2Zgh5KbVvvbyD2cmRhg/
/nP1ZAFJuRBlgQC0k8tFyLStFaT2eTUrsd4AiH8LZIm6hTeUOes5mh18NLLhJlOj
hIIYE5xFW725kJuXPWQ9bcHIHxPEQ2Uzd4pRoyBHJLahsX9JYar4RGgLFIb4GzeW
n7JtOQ+F0neAhBzcbRMijl2f19FdipneYsUWQ+ahsv1SwPDinnECo313ag0v1TUV
SNZqfjaHn5X/BPVGJLv9nlrxXcpb9U7MHhPkVKsz4SHtd5aHFhvjKK1UYv7py1vV
uikJmMp3CSBjkEowaP49hn/InpXKwsuLYTMg1OAD91/1MUOQs8Zm/ZMr8E3gCUeY
vrT1z+0JnbEowI7F4wTSTgC3B600Aqw/J2/G/92Amj4SbPrZQtfE2zZP0VqRhAsI
sfw4rRQoZCH5tO+KimWZrOYwDqfZjuveYA0KTVQcnVmFtyzC8sCkEm6MmEai5uW9
sVMhBGg/NhoiRNG2h+ykYxZa0CGBWrViumRnhcpdxRTwenMWu1+yApZl14P3D4R4
KcbfwbBz7QHUc4Rdg0j83mLJmFzvM1FU7jIQQL7D3vRlv/dGjD8VVMP4LxeQEuVJ
W7J4lVmBAJHBPbUvCoEUvUEpsKFdlj4SWL5GclMBH37dGMv5hJZWshbeuRXWlvvL
umuCoaTHIHBRhxCe4WZoFRDPYfkRXX2J59XvS8ryREb19yIr0kb7loNFBOv+YDG0
fq44yoe1AKEqM7GRwe4pauPob02pDOhdpqRkBkOzHgbHSAb1F08kMuTSqdcco3UC
G3VDWuRaQ6pDfPUu88+cRzCd3fxMTfFPHeQIxjezTDQFy6flr/TKn6oDPNpNlMJW
oj6zExW3IZjBv7pWW7oVJgzkCvFtQ0RzsfAEez/6DRQ9mppnua2mFJGJpgInu0nD
qPkz7AFsB3taaX7FBwvkC57VHKDKuT37OlEhoIBQ8eQFE1KJclRY1fxx3whr2j+0
slvXZM+C5ggCpYeM7fmTJ77q+Yj5UEew0vZKR1PtL4a11qC523y6CLz4vrVWWaoD
AKckouQjisNbrmehCtd4zWxaLW6NU7G+MZEhYA8kGg5p1PSI6Y/9EZsDtaaXDdU6
Ykj5d8WB1RqHoYVUdGmJg0Npr3aTEC1O4GABvH58UGrLSX4b8TLOvNpS746kNHpE
2BbZOBa1b2iRLD+aKw2Jet80gfn09S75yAeBulKCJ9Le9ryP0wyOWS5agndxDJqh
PNCxzI7WtOq++8hBkibIQ6acgk6tvt3pxLJu349YmHqBjymCC7lhyR50WTqYJLVM
EH5/HXT7qcFE46qBpf/4F+zaC1pxx+put9idE/MIpFNllRLrysWp/QLlnqrxETxt
IuMkBgfMTfjbmv7QC07WIufLjrLO4bDg//4LCQRC+/71GhV1ZjkPhbYFtTSYYW4S
QNNZqNNmOaOoOINW/SzrrtNnO1ohGHxk6DtuASDYjUwf2dN0QV6EwH3h69ipfdTC
RmNU7N3JW5EEa1jmKY9Wfb6crTeVWmjswAOhLU4A6tZ28CB+Bg0gwGay/pCMMF6X
iUE1YRdJj+M0p85Nze9ksL0S/QXbdpmy1y4hnxUF91uSQn7jo9pKCL+Ea5mYicUQ
Fj8D4zqyasGcbs3ojSJ3Na0+M9YXOjUCVBjayy/nNRbbjFPCoY3POvi5gmo9hJok
D/83pZrDwVpSRcTmXNsvIuIRnn2YWMXX357K1gQmmn5cNTMxQPiarbD9/1f8qgrN
sO7Wo5GFVcvba+AK84i8uW236ndUIGtVwqC/uxTCt0aUSbGhVOwbqcrEeismIdkP
Jwzj3Z2i5VbBDQpP9ngC1XCyn2PcwkNaxDicnVmPjV+YYwSkgR2ZyDS3CfHAvyTs
OPiTLafFyLmmyhCEPSPglmHUKoTnPRCL37WFy+G9RarFyk0gRl/WA5RsaBdnepe+
A2F+UfkSlT/NlpXK6U+3wtaHTWtRFmmvSU2W+cWCoMMkX/Ci8fDKG3q2h4ijvS+J
UwEvSyqTvwdgmevfPPaRfbqpEyrY/Iuq0tBf4/9lQmL1rDwB+W7P6vY9YScLxEO6
beG2bA21UGHMr0/PPHcHwUVA1pVs/eGkf2GUIs3Yidw0oVDPFmPodT9zvwI7Q3Kz
R/rCEdKnYQAnPfMHmiiX4vg907ORmacWkp/wFPmgbgknSlqV1nVaP6TnqcmETU6t
ShE54TQMzvK4TGmd+A14PCo7rvG92H4D85/69MhcQbfE9sNye9mhkY0Y5LTzHb95
4cfiTzrm9OcUx3pouApZROHtfV/BxvfpLsxqhLwplfS3Y/ROw0H11bp9tEothuTt
DqlF7ouZ15YRJJ6DcBZNx+WlI4bHBRZXLwvwG35I5sWQdCSpWF7QR2HddsnObXfU
gQq1zirq34oYOWK4VPeb9Bn/2P2jwkxMt7fxcGzxOHcTP/EzUal6/+B+RfiPlDdM
7xqoD5V4cZUYgAt2+rRTsupzIAtx07ZJB2dK9RDaMSIMTlUeOPP9210jGiUOsw0q
OPwoTycY0F9AEFgwOItXjWkZC2zVenbUCrnexTiWXgfgrHA21/mP0GbMr7W2TMze
rY+xa+TSSfyB4V2PU4vmcLejsZEvEm51yfCWT2VwQiIa0aPc3Qe6DqT+T/Nj3JiV
dKCOysS2c0VyM4QCYUhSbLQI6m+SqP5Snrn+cSvstB/Q5de7oJ7pMzV1L7vgLtT9
C1KEWUt0+fSxH51cdoj2QSXH68ulZein7wjRNLcqHYSQ4T48T216Vs8K7nZ4aH+b
A+7wpY7Wkb+QcaY/Y/YFcCwnqfNdHSHOuBJseSe3cLUn7CrVS2L4rVE/kSpwNgcD
KF/xdnWTSJ8U1HMEPpeBWHcgu46c05Ss0+A1s6Qqi+Ts8pBJhGJetE+YxfqfhA0t
Offi+pSUKvF4yOQeBX/9imwSEBcE/l0Ys7OIEMaRhj9VW5NQeuZPwLyZbpMfwKXY
SiqVaR29Bieq1RjQ4vmvrCACrMfveunaPs+MrrJwTKRWh1P6MjFxfmuefw5dzyeU
M9JXbcv6RfnSyJbi9j8ffvbnKSUA9omtxaYGupEYJuLHNZAcQ2w01mghl+3cuDOI
SAqky/Fj6o4LEZ3VaNvsOmfh+Q+s9EXJL5CSNpZKQOctvLzuX0/UZzaGi7GCGoew
qMvPoXn9tpG1cT23Kw0wvmCrNLCsIkIebLOpBRQTMUeKk6jILdhrSFGYb2A2DvZI
k3OJ1mMbYM8l91ll3oCoD/76NImu4kJO+cbbzxC+AKefTzaLI/XUKtJY13rI6/BM
czMFTYUlavhfq3AEmy8p8yvTpu/qb7MfWYtJ6+UrJSVvfb//MltYGajY6EbMe+lE
qE80c/LfACyWTa4JNbs9WrZesO3m/2alSGNJhjxrrXEsuwF8L7RTpTGcTANc2sZB
gUWRvyoSIBxb4V07qYlY3OeHOlxX2DffUbb84bFu3RqyV+/xpm57cmU282N4lM7c
t3UT4S7cwQTGoHrighg3pxM7HrDtAFouY4lHvEg8GeynJUyE1PBptiArWIHj4xlf
BATdh4oBgz3+oah6yDGO6fqXq594qfIDVBvANU5Ve07ToycCobDS19QPEE9oHHKf
F3pxZy1GKRklecuMbjqsm16qbk1Fu5OK/eEcr38fUWbaLR27APGkQ2JMZeQvfe6C
TyzWLaci+WbQB9Cm/K9lQ4j5zZJZpJejfkAuI6R/w4Xhtu+JFtavdGPskz/t9k23
wv62/j+VIuoFuIEHV9n9qgI1HEiiaKL7lA43lMPUMSCL9VUqx2eHlPBS8CeeNNPa
Qo2eWYdMyHUdM9PG8mQXuZMKyo/FwPl5FXV9ZXxO3Ugx2idmlTXnMx1+huOof6bT
REItFS0gS8aUuShSGgw6/D7MgmLUax+1GUiY7XJY7MDQYSyYNp+24+l1IYkFfhAJ
wCvbKK53nJSgJrI8Eoe5XOdiM/7j4fph9V5cKC8WwM52hLDaVLZJm3MREguBVl/1
W+m1LCPrfZ3AL4HfeWwUOTxbco4dVmr9x7uRxAronaxFd5p0bmUFRYvF+vSKB72o
LGi0b76Plhjg1K6A7A2AOZg/BeiZVjfabVokO9UNTriV23V6rT7qBvwGYwy7ywbN
mnRVY0tL4LlXGEyoZEVXY8T/CVN0JQy4HF8Uk1R3AYcm+bX5AUEL5uhYxTGXA3OW
tWepd2VRe9cuyg9BF1gUGjEL0/9FF8+5proHkgzCxgxlCkiHK07PXW1hEJF0g1nO
ypQEGxppztu9PHADAkLV5YW5almKK9YOMBOByyeV/LPTnqHTX7EmARusoYQSWRdu
ctGSP4V/yckfJn+cJvZY+/n+tvAFAsl08oVpy6jSdRDbs9poUFTUzo/ecqh3kcO9
k2qoO6dNQrLBn6QGui0WAoluAMIZoYKqJ5NFxXkB8z/BiRT9+qrBQqYF5FYX/YKN
eSn5zS+W3BizaIiIZrFjSjwaR+gLWvYzuO6ovgfxKjxaziwQAUZvgLUXucUb2lTx
Mlv/ESjsRsWhWgAnn+IFz56wNkXB3Hc3uNS4OzsTEu0pW/MBhCl000xjkhc1uDRv
D9oUGeEQCq4JNSfnjeG6gEF33knebQJEH9EYrYfyakW3fmBd4Z7tBpZOrTHpUkJ5
QOGSlVSkF6VzH1/DZdme/rbhZh690Igx89otKdaTDID/Z1/8jl8i0sN1V2S4euxu
5z9Q51XZ58PHO6Nwfee58XyxMtX/WP4JaGiiz3g/mz8sA+9G/9lr2NiSQpzcNGFA
l1RwgR+fMoL/OeyGukUEyUgVVcX+Y78gKzqO9uJ08mci0Z67j7ry7+gLI5GSJTft
dqp4IKiORKxPYaOJK3xJtKCuMrbe2PH/EKlnHNmiJmGCzhNThHG0mQOXdXzma9Wj
+GtvTvOHCLt3kIz8Aoj+uvVlTJJFtIyiOQJCc4vXyuHwiyj+XmGR344zaiuKEWlR
z9iduxPGH1pFz9sVa54XPDNJqaiwM1JnwKlcVDwXLhgfXOXCcqF5GcOH8b9lr+ds
JYKpM7R0heQY3EUaomg0psW8NUp/ON+5NpgJ6mtwtIndSZ5IT6f+wi4Xqn02kN2k
sivyQPYK5wCPACkupJG6+7UHsZtJca9D+HS0L9hcQ5g7u2OBr9N2QFo6wgDyYR8D
4SpDNfMvBHckUvjcvcQBr8p5nBn2DClOhblDUwPBIQKxU4gWqn94OG0fHO/zNKZI
mYWp//ve4zxp6o3S/ydOYh+iwuuSfdaNHilXjvYErWbXPLFOX8Hejm92M7BH07Ea
QUE63bHVdxc1l8xWmDtnzY+ULiQhRWmIP99qYNQwXh6Qv22pSc8B65yqPyFdLpgd
ZQccDO93xCkVE5Ou/NhJpkKQEbxDqMrsGvMf9C+nQMek2zQPpnCsJyyGgGD8jmBI
6lC7hSFe/HzRrrSlQMNU8xmoWqYm4WTnez5tgj62rKx6P+0PiP1SNPRfNM09CL1d
gm9wNyBfT4QIUr4t8FbLMwe9K5J5JAXQQY4K7Ep4XHhyMjkUTw/yrP3UyJ14NKiV
T72ZEvcQ6WRRvL2nS0OGfXDb6jhAEkAJGEsMRfgG0rVaO110wQ8c8H+pgeVxQtGK
TUBtviwgghSUpCocoy46eu9jQCCVexGtOBCQtne8I/gB+pkA9oj4EoJ3UAJPJG/V
4E8PlFBV8HHrvYx5t18O60EvJqYDW4WRtqhjINPRqj0dUx2s409PGSURSrtbp2+z
iutAsO8TyDVAcU3cFRZncH/kAqdowrkHn8agzlSAiA1owPlcITXlqjgW6er6FYqE
3dQblVGVphMFR0U0m2LM5c7x9QrIByp91+VWt3EO71iNrXOxDdgYCAFFpB9Thum/
KoBIzdA07OmV4q9VO9YFc+j3Rc4ByOxwGBrQHNbKMBAyYkx/J1rPHS7gy22m95kR
RWHq99UnapE1HLLljgW441kDEJsA3VK8isTRn/EM3qmiwOgBNvrmsgNaBafQUMHa
mtC5+wZOxmc9jvQXk68gjEoV4W44Ajr/IljtyLbUv+DyeCUxH5kK3ZvZDnS+RiJ/
+Hke/WtCMa+pac42oZ4pfQ8+PbgJEkZpffWU29B2XQbT3nOilVeroTsWu3fnP+kJ
esBz/I1rUT52EdXMFYUXjoJxw3y2qVwwW60FNYe2exzP190pyo0Rl/DyFHVqqpD3
ofrma3IqRbvrkwmzXfdn2vqnlcjkBxo40IDwhMX0XtAzBnU3EIEgjw54Qa3t67go
ii3dMynnsdc2Qjj9CWlY37G2wtFaH4pAn7yevZLsopg2XJdj2YbVUdhQi9XCANZ2
dFpqqSg9wIyaL96TMtetP2+7EUV8oX9OArIgiCqAOJtmdoPqwSB7xIbvybBWgpLm
n+nkszFaQWlVPYvNR+DSHeqsTtGiDHe5Uvt46EEaV5Ily+N+c7PpDnKBk9Cn64UW
hU3g9UEWQMMUKBnK6pNyR4LOam74PyyuuW7+5s35zXAvrm20HNjsh6tL1qtzvaOE
+dVNRUZHot5pV96eQx8tSgVrNyXTg2KsQVpwH/ve/nU6rGhI0yym8NcNpn3QxP97
pgMtjA8KRFS2Qx2cF3sLMJA5XQGU90qwbQ2eP+KpHvct8JrQ5eJE5MhvqjA6hNbt
SzrkfP4qMlklhzWdZV/NSAXx8DJeZZtiwOlH9SJASF7OcWOld5CFOyNVb0hYU03/
fLrnrzd3RoACuKfkL7O4KbOzTRIn8bMJ+NtRUIjaMbcDBT4CIyFG5Pma+zbj9Wfw
gC8F77oFK7GFFCkvfXsYfvlt+9gYCLZ823TLk7q/Ljf7OgFQcCUZsIfqXwdwePBV
2zjO8Ktf4OHD2sDFMBlwEHIgPmsMOSlitwVfS1cq8SC4cux53iAFTmzX4VWfsDO1
Yc0qh/1rcHfRIdGP8fhQHuVd87hngnP119HmrfS1UXwRnDmCuJSCZoEwhgqAdCiC
j4+T+GA4vu+/RmLNURzRcpwJ6pI9/AvZ1HMUiVB+kLm02pDdO7ymqOP/AhjeNQNZ
/hA2WdpBe/q7CBgODoMmXjKB9SFufdZ8B5Rf3WnKeHl+630bTFgP5CJE73fX6Gx5
03hrtOJwLLN1aoruxmmfkX+YqHadZOqxJXqqWI2wi5Njcqn4ZW5Z3qdOlU7bna2w
/fKE5+WCM7KFzypG1Rx/ZRWVdkgOxD8Aka2uJdHCv2AW83DMGeXb3qugxiYVs5s4
MdpzOPPSXYstdjHfIjQJh3AHu4lZ+P5CMMxy6hs+UOz30xpnvJ5CAV141EHfyHMy
jNt1ro6f2DmIYOBNZZfQaGFLOypsyWMWF1nVmC9dnhgnvGCzDONtIVQFdZcRqVf2
ekM5AQBsRxBNI6fR2PUGwuZg8Yjw1N0Y/IH/DJOyFiE+ba92+SMT2ke5xho0OGIh
Mk+S4RrhBjzcq51PpRPsksv3G+gVZUVeiedhrfy6AYqCNWhYHe6I/8HmMBxd4bix
kvHLXWjtirKX75O0JT2kqNv6MKzg3MAjTZLX6iX3uNXVXWl8fHptkJiafCV/w9Un
9nGYDi5NMdRqwnEW19vSrVMGy7h59KPHSppdZDITXHNewLwzBUf4MJXMJhf2jg+o
7TR6E8KpqCx6kAdauEreyJbrQNj/8vuGastAd172HVNhz4Fn3dzFjibT7h9Kxr/l
s7VfWOoNz/Nm9WE4+LbMb9vEe+iHu/2+dBjjGxYqP9HdkFtwEo7y6x4AOb6I7S7z
+mgdCXSBLlCXe8T/4YSf14O6wKPfPiLBAguG/2UPNLSwuUtYbfrJLLpj9VQqOaf2
IhlddvaMaPHG0LYK1dq9h+v5HmTg+Sp8LslCjExu42eCKNWJZij8YCgrdQ6TlHvJ
Nsv6BUWSv1j5VNT8FVbcgQQDBsUWx+m5Q6N6Ft+LzNsbqXGQ2VTq2axcAqN/UMh/
ICs+eL/UE4mo58GtT2ITfRvZTxSwi+hJpFxABO//0p28BGNXIIiRjjZeNKmyyf/X
rXOR3sr0NgszVzREo42oDRKj9XlRCEL4aAJOowaPBZkb511+O+fkNga7NX6SXjUl
WKpXf58JkdnBsNjrdwUdy4fCFVkV3aFK/tI3QcQ7IVobl+rGR+iYmNNKw4c4K05j
sOoD9wUQG9Zq/vY5EHSbJvE/chqOBRNDzYHXatB3j0jcur7cSJC4SvzPdtUHUaHS
zelrzAtuwo9pHyxdnYp6E4NIewz5KTl4lYR70XzJsv1nh+0GdYgP36JDn2U9k5IG
dvozfa0WgVN3IeRYMjp9j1KiCfo3tu9CojFTPV0mQZLw2dmIZ4MIIK86d3NddrnM
LsiQA04QxUXZUW4eOQqL5H2b40PZP3rRk20T9s5jXN/SuXCPq0EgkvxdTiH+HhOV
JtU/ebJsnIw0sTK33dWb/jyPu/MjnYKQrdJYMU3DwRepkuCY9FilWNT+/49IArY8
Crwk+bTjAFl7nLi+qVbyys9MN7Eij5oYNrB+4XWSyXxBb+hd45Ct4g/Eb0nrPFkQ
9kaYi2i7cWoQmFxU43DRajkxu57WifVBF7rSjFb/hLRmYMZ28+uXpfCnvDel/5an
miAKyvvfDuU0E0HchW6Vp1gl5tLAY19vHycYN3+GdGDf8B/UdvAcPqZtOqJRS/UG
5AMdi62bzCL7G+BM8sMLBa87rI4fllQ+EFHAt2KLU46FwxpsnnE3q7RPVsb2BwET
HZbxJqdOdCNL17kDXkUauA2IimqFFB8uulv0yAzv9KrRh1r0iRyCwFoNwUdhi4Kx
uGPhq21M0PRn9SCBo3bRgSOksOYJ+JelmofLbBYbE8Hskk1uXMBdoDQczrWMhHYf
TXVSGvX642+JVwrgVcObV8Fh6tgFemFiWQvBrIkLrVCBTaIPFAWRc0SGZWMLpouD
XcCeowm8/sfIwJm4vxyiwgxN2KhtxjfMKo915HmnwwpY4eSoj6D+BAaksa8N3P8K
lcxU5viynDn0SeA5e3ccU9AoY0xPZh2wHmBntDeZYxGF6KtDDsDL8xBQsPKdDE9D
u1v+XenTnzFxLcD8Q4IUBxSh2k/Cw+xFBx9Qd2c5C7ei+Nhnvyaj358z5cHZaaFq
Obj6uYAA3X9SWSk2e/J4cUZ/nae1NALVM9hOJMFOTcNh+eItyFLQoQkg6xdEKDXV
K3xW9bwIPR5Glgy2BFhBflVmLHNvPYjX+Nh78sfpw3ulEk9oXYAMzoGnCvbWZMYe
0FvlkPDYm8EYOWwM+wfIZRwIGpgPTeriaosM7V0dCSgDxpu6LqBGxblcxLlgR662
efoRmrJplnk0t0VmgIkDfZsVHrKpfSKdXobVHE0VFACWqxdsqYaIzzaTChazxo5g
g+JJ43pkj50fRnsdAuEs4XNvkDvmmMpEJ5Ph3q4YJuSpJwe8VKYgm7I58/vgxAds
s3dNa1M2ohdBx6FbDhhGcFR5aYceSXvT6q4BqGl+8GEJ3SU6IoL9o97WSJ0llJDV
gIL8x842noMB40m77YA3u00IhLL0Tr3UwKxwvA5axF5gjE51IMEHpvCj9OiUiM0k
vB2/p3awMuQI6fK++1lxENBtbs118I+GyJyv0IvgIkhpafYY7bluBX5lUQlzKK31
NsvS6NRGwZ67YlV1JH10We1rKfvHd0D4B1PMTAP/XLiX492sx4ROBqnm1srF7Fhz
QeR+J8ThQ6qsOxWxNSuq4UqcUCTlawK2FTwRO+433qheqOfWgVkRiisxYC7TrzWH
CAGS7s6Ps1z6gvA5AzlmF/AvxicydNpeDiUGfnypRYxEpW9J99VkvW+Ideng86Hl
fkRG7XWvFSDU6zBJ4HbOTAfxNAC6DuuQh+34z3WMRygzMTDYHyPBCWSupD6I4+7j
ICD6meL5s4pQocc8134cC8+bQ9YgNW95o9jCXCKD3wi3cZCAmupAEfjd/yQKRvmY
MKL76pmrshYeUBPv9F6vAOBnW6iJ30Ay3rVHrzvCxolLJn4WeCacKCgLRZ/KuLsx
3BhrLNFkHmWVdWb+sF7K5YqFzcUl4buzwsOoprmYI6piArGZIBVC0f5fcnKV5Byw
ag5SHI+vIakHxcnD2VL4tFuYi4MY4jZ7Q1Q+Wmq/GlUrqvFFEEoGnzA9RfwdQZ94
QG/ozsx/6Tms0KiPliUflNRz1O1IRReO2Zmtyo4QnhSisC3YXGW/DrZs7FHhS6of
0a+fUkkqdVVSF2v5avVQc+sQa+KzP6R6ZYIO7Mua/A8cTBLr8nzF49nK6D9Dl4bN
ZSPFh0XFHWr16qWoExCD5irERvB1MG7obk/+tJdV6jlJnM9JIsus3AMAsOZF/ZJS
wTAUANKi64zcO1KEihMCIShtpGuSPRZVZD7Wc0oasjKso00stu1k1tmKeoZ2h4yF
tTYXtgE8ZAMgEgU2GbSDdRfsHYfdwoYWHn7dWQDCKuQmWT9cDyMFxe+RvMN8r1eo
0RPDTUIjcJCA1v28b6MeuRokLTrK6wEyWigGQtnD570gMb5gomWz5PhzM0S6JD98
/K1neXGkpCCQcsDZnzcqygiBt79SoIKj02QiGgCJ44xunwQ3L4cSthU1IZZIxAuh
ot1nQAu2ecGeYj6C4ugt+mWR0Hz9zs9Yqx1AUzlZkg8mHu3pm5JcIflWkwPQ7gNY
+i3MfhwtTM/wxyFSYaYBeYtRRmurDgDQwALohjtfnz0rI3BappxUXvVDXIs/zsmL
7XcDI8kHFhsrvi/yKqJXOsAIjOJJuzw9xZYhlLfEehCbZrheyW2VWykg7IRExHn6
MCgmGL0FcmHi3FGRlmCYshpXOiAR8cY3236xAbF/hZUnkk1MDJ5knDiaR5jVEgMe
aqEwYDHGhVgEYAeuKNcEYwIA/XAhLfdqMq7iWr+Z0T+YzoZSMYEH+R505dhyCuex
pN2TkShtRkumWVkL6SYsSrZ5fud2MxCQKKEf9dyY0onb5oVehTwExAq+HFnbvXAJ
NFqmCx4CG1FBdzuCUYmA5FhLzSZbNrWa4HxDKye6ql5PZ24zhXzv7sdz8P6Oqn5I
C/+SrWUYJPUzz79W6oxVuDQq38SIIrgLlC2qdY+6Eu24OT6kpZMn4Mx4c6O9/fRB
kbIGRxryciSyDeoqvZ44GlGNx0Rncbh6rT7GUhTwDxn4uVHjCUdaT6cqXnq2MJ9G
ejBYep4tsd2nw/51vbRZ7yEuY+1dciIoOTqieqOyEoyANghaOhA8KhTqnY0B+cZB
kDciZ3KsOqupJKg85496RABB06WLZhACq2JQKMKpAok8nDbh9rWr+wy6dQx6bcQY
CX6F3F38hWFp2es1Mkv0uXXHijjndOR4j0BSJTD7LulLDVjOPfOZGcZbs84vd1mJ
StnjuL0/EsDLFzTBP90kC0WUqJ6F5LCq8rd9q12Pe/dyfQNAUbcFs92HVTgcrEnk
ZbjlCICaXYEbx9TZEcQX/RHUhhZOiJknWvOaZ8k8dWJvQwfcO+5aJssXrQMG/6HA
lfRWG7yu5udS1CixI5uBQMPV1ujG06NkWsFiISPxt5KHBfpuGixSdLSyCg3RifDG
SqmFHCYV8B/5/JENGpvzD3jinYzHjx5rcpB9jHfPI68Xj2UR46lpWUAKHKM1bqcz
LiQ/RF3lJGx6syCn2ijaLq7sanO1DI52rvw7QbgB1iERghnQJjqmVMogauCGcbXQ
V6uCfPSz5w/TaitwOLdUfDd/1w2Tcd6FzgfFkt2wtQt+GpfCad45FnxEiJcXWddW
cESDRehamAyAmvxEUd7W7Vzp/mQTgqFJs8AVUw+N2ONUH80P4i98AfM6ue/hTmP9
sMV7UYkY+iBQJXq+6flQe/52vra4eoLK41/Q2RWiR1ue4HwbClW+FPjloaEGTSnV
gnOY6TlUyPtgXzJpGmpXGAlqjc9DbErVA71BAE4nlRyfY17RykjBaZskHr47Bqtr
RtnCqOupOqkLgEbs/6V+81d4d9VBxvS/oARhXm3B8RsTKktnVjbRvzytcPgfOOGn
jFP7XTRWK4jJdaPm5ni82YNPXUbgAmcwTccvUb5T6C3h1QyMJLT8D/ZoFKgyh6Tm
IPTqhR/aH/HnheIA8smivc+Cd02heC/4JmK9WiXNRUUOBISszbPagZXj6DV4XMAY
yjE5BJJqjba48WUFGrZJ/hidgeG/G2YMeS4LyHoCd6HJ8bGJac2GJWka/+JW0nYv
RiLWrkrQsUIu4LzjFT9KsdxyX51XJ9tXQp1XIt7PNCgxwwTZJzWXhQV7r5qSznwg
nLqLmoDgZVWZG6wlsxEvMa1QRGPcndmXOuopbVWM5E9jkT7hMm3aFX8b8IQNn8/e
DM1w8vMsgy4jh6VyZXkklOJgJWQb172QOsSKwgK1ZKiPtZMKwnMpuCULAiDZ2W+d
e+BIBrCp/DYIz/wp6p1RYB8CnGqN0jzsUWizjf9LirPd5P+vZKBHlLHGC7kmxwDQ
9AwJLjjTV+/X4B2iRk8XCnB2jcM/vMP66YggWgqvgPJjbZBLrVNdFCbr4nCZhIc3
RutYxSsD51ItUv0HDVJa1esObmhEUT7IdbvKTg+EQPJ95aSy7+eaQ5k0LbaN3sGc
T5A7Ev8mEjyj5FVYaU63Rx8aZhEBXqDR2rfnfvqZFoTRWPQBChxSCcGQiPLi4w6y
HXCbNnxTb+8aNIK8oDgIH4Hfs3TtkXnD3mqxQNoyDTxADB1d07f989bR1UDLIQm0
PXMNm30/EF6HJFRDHRi3SshQR/0FmfEBfHyf4ezFWEuYpH45iGYNctI4+S51/QC1
2W6KrgDZIyD5uPb5Q9rBHe8WlfN8RQDcuPyD+yHQ58LiR0VNd+AzwIZtiWbYwCay
IxVwvX0kIx1qv9n0wthEOFP7lzv4Y0AVK96lwIq46Eno5jXkf6h4qmuUqwF0R4mp
3IHIlTsa44g7ycTkRuZO25wqgvq4gsTuC85ex/r1RPUxL/ynve1Tvoo1vVXpCRec
63QvyetScI4YFEyHQupjT5soZBeznIcRIThlABtWxaD7gjWc2wfbWUZhLm3AZicF
MXw6dqPzu1l4+yPKPvrvJgAT3F1wk3xgmd/2XzP/EWYXTcfydB7vDlP9majCNJvb
NhxJclc/7LR/IXMrJLTt6fC5RHVNgE+Vh1bHBm4r1DcEwQcT7UQL376Lu7Bp5L/1
MNNokwBNZL3VN0o55bU4MQqgCfVytm9mQaMeTPNtgVN5CwBAhEJjRvBzWOJR8/Xe
b+hKB0ppBrpdo+k2NjtVrfjTJNV5Pn3yM8M4HGzIrRBK58zfGqkyajTdwB2jYXGQ
cLnyh6Aokf3eHhTuCtqUk6w/a4BeTLTkIWlmleUzqdd+TZSk8EA3bOVNIEMed9ci
LiSiOjRDu+2e381Hh6ODYa9Fbn/Gts8gQ5azJx0rEO6TwgYOVjWqWLzHrwHueoTU
pVt0uX9C72GLJ8gaCkLPTbG8W7MPcAaE8o+hG/f8fJSvvEHzCSxhl37SJqYcQfTd
BDj6GSfQLxZ54+wxRM5Yi8gpu2jqZuvqm0bjzqnpoQ/lLW4xH2d07GynDAsk8dZ0
5VT/sLPq8Kxrn7uA5QN2WDMAEd1Xhq8z8eBubvevMrIohYQ4JLMcdzYogUfrml9a
Wt7IAhrKgtKfwYfPn6R1o4ftOYyCi/VxbHRI+lcQ+OJZG4psm2LT8RqN5DkVA6xL
dydzLHNKvIdQ/VPUWiO4OVzXmhb/PLTnyzpOGPnerzf+ztdSY0iqng8H8hn8H8gm
dMZXrSw9+VGrKG9U4VS2zcbaRQLAyQVojk6AMrXDVzyhy/lLL5GMXqggdcPyN3n8
ct0TtJe7sTedjI+TdZLFN1DRFJmKwNUYk+fR684VZEqvDhv5ANN5Rp20vGI0FM8Q
pVhM9OlfuM3qVx/Az0lYPV0VsvjoPCYAk/Avnr0T4s+oKQYLcTcwhJR+RYnvnTs3
VMczCPYsi6jFErRB3zIZG6XzLR4tgLW6PcHn7c8BKb+GLkdkKrppxYkHMX8vHAy5
4f70YHPsVwxY41jeYOaHtmX0N79oio2niLKCqr/Z2qtr44k6QGf+qRth/jBJwfZL
UwQX7UDTMc/FDWT64+saLST+vcOPXSORNUo9z5RBWkW9vrIyfVGxZpjjvIRoBpkb
V59ySgcLmuVdD1J7OVnDrn0cemiDkrh/kIhvXZf3t/ApYrbzDW5xf/F/syQiY5xz
ZXTgmDETauqU+iYqRrDh0VkcYu6LOQHvLcVifXCHNtFprRl4OwARHaT7APiDzaYl
QmVIUHF1RanClJAN0jzb5eO0vCiZzYMb6rApTPw0TV+3rxapDhn+osshN/Tqqszw
TnGUgU4/nh/hXSad0ISwHc591MjrCZ+XicfxUul/zFbJwEeOTjKkg7R2iw1Lhm/8
nzNjrsmOc9t0EL+TFQVQkMEuAeJ9oZ11hXGd/SqGh8SwZOHRE62WoUulqQ99E/Dx
6HJ9tLP1G9Vd5wJp1so0fLuHnz/bM4wjayLzrUOdY2dXI/BBHnu8F+HEr6cmLh68
qTFfknAANRwQK6pvh+hPkEoxvjfPmzFsi12LSxCjWsqy4wTjBB8hJM5yy1zZnLZw
YUMXQJwlNFiNyyHzIdS7412GpxbFhoA/IUZ3ZDL5SK7BK/jJcFhMvp88vdRMeBQr
1Wnwfo/0kePu/ANqUpaDNZJYPp45eabYJoNtIKAgy1117reHnVqUxjWvV4EiNgR/
m/4SPzfNK0Hy+1WSVOuxw0EErGpNZgb3pPjbADjigrSlOtIeHNVZsG+fYjAfl8AY
vCD7Yyc5urDsuCi4QGxIuSf+Usi/Z/UD+ghAGYlXbuOlXD1hIpv6TCy70uDqgyiL
HvKF1Cwpof77DEMY1HtFglvKoFL6tHs4UGS9NFIZ4lbrp1Lv5/X3oOhSYl60FeH1
dJhSA2FJLZ1JTMp3Q5OthxqBtqKETy/lbL/LYMtnWCQ9GzFyiwO5J/kgVsuHV/5R
T7zpqrHPIr6T8y8M11FK9ebyzbU2kabUBD1Y81bHCQWsxjlaBuzE/VJu1Cq6CFh0
bRydW3Xuy9QicYgY0iacZzJ4SDudiUnRL5T2w6fgqA8J+XsQAMCaf0t6Aey8YamT
dh/BgsucCIeerImL9dMbSpv4CBmhcJKJp+qLacVeoOEqrg9jjjqo2xu5EdFtnabT
6GQnOIoSDGHzhrkPI1ULc+SnVpFsIkXbCtyUBDQiA9p4QYQU2LzZ9TWDCLYIAvzL
MY2qMvn9B6BkWJjae/DuxPqtFcja/KfVXH17hZDxPwN9Wp705ZIc9YRawzs6FsBt
ALWK6KSGZ5+SCyfc/re1LyAvUbGLB3Y39FJJdIU2037trV02RKIxYx853UZ/kF6h
iea2xiV/cxc/c4Gf8JISgi7DVRYUpCzKkziq/lyD+x5L+cZw8ldV6P3TSeHd1GgV
T/qYoY1S2DVzYW5R+P/VMirNdOj7yv9cizsCvZ4vz93a3OUpDcjaBLo6Vd0uuU2F
SrQEEvoaPnnLzjJ5Mj1Z6nvlwbtOC3f6k5lgoM/5U10AwuEQR0/uBf/p/EHMqAyu
bE3a8DTBe9RXJCFS1lc6AigcHdlnlEv7M2Umum7dCILypjGM0U0D3k1iNPp34uI3
0MjXPFkJE0wuBLKnW43QQ6Sd4YDLFW9JgvbtM3//IqReG4TKzb+jj4iX3oywqQ26
MAAwFPIxOqX4LwW5p+cHHKFDvaEnwICDm3T6S2Gr53t7p9vghBmMbbn7HvTNVS7g
/XlGiIJ+Qpjkp1xeZDFrUqgi0U5BHk+IN/BwjAJQepAFOAkK1sOLjtRlHyq8NZzl
zUClbtNNoaC1z/BRnRU7qFj7oRc98OgNiq5q55ZSvtcu4MgX2KWI+FmpYPB26Q2F
m+7n2PAp1Z+ekFk89+r7kWDGFVjIfmIR3nmh1PNxvuz0RjxGxCVOYCYf9kpygC/t
yEAuJ3pFNTwXOGvGxBNaf+r3R8d1mJx5Hl9MdS5esUl0YPRHUnDZ+PXKe0UcbCaA
UnrRLb0pPf+WfGeS5gEGTfYqqRuHg2uhYFaroVc4BQyYjv3dc+ioW8JPuA/r956Y
nm2J398N4L7j4z7H8ljl7y+51LPh5P2qG05yU8AoUgof0+OHsyKVeVX8ite4tJPR
BvmOT9fX4bbPESiCmVR0JFyKeVXnQDWcSX9VuxWdiZjy/A4lfcxmkxMaxyjh1eHH
HlHcHnB55A94iZ3iWf4UrpfCvxtyHoJY6ujKwuX1c6hSBnCicy+gCdtXwXOws/zv
PNjqEFmHsBinImmcK/IZAuj/8JLOQcCiVU2/AwEY8ZCoTJOXBqO8zCY1aF6oe6B/
TQRpUlqzmzzuHHl/vgL1YTCRSJCea/kjryuwzxlQjYy5gYQ7/ln4+PL35wkhJxNX
3Vcy+8eMK+Ep3LFsr6vtDb5OkIRbTWgLnFYLg+HPPeKKjF9EIsCoejmKE0F1XKII
8XhvDa7hbCKVB4ZixlN3AEA5ZLXbp97hN7F2jphFGI1hRFbkN2nhWaMUF+a9PAEc
J82gCshP6XPSMcNWFJCYJ/gBdHzgTzeggiiu8F/vTg468+XpQTmOZ9yqarClL6i9
MDW0lj/SfihbXD9LuSoQiuwnfAlJefazkcAxD5nlFLC5rOpxBIfT52YFC5n9350N
P6cKw2MJNtGcJZZX2koauHnB2ZrEdy2n5811c7tQaczoyAE/7Uw79Zc29IYmPYrY
Vo9fDhdIPjoa4/DH6Scbg8M0UftDmLw38bfIBbhkmmZVQUgW3qe8llrisQrv3k2G
MCRV8LlBcbFE2jL7XrALHtiravwfSCPCLV8FeUtlxfqngsQdUzE6vMGDgXmRqvYx
wZWR6REbH2wGok7ANsUcnl5ITATk2q//x8KmIZ01obrfZ+dUnIYMM49b2dLsyrfy
eJ4Nq10jw0xv2t8hkWTGxWsdUF44ZU0yhvwRhngw9rzWZZQoDYwgy6r5hzHrTwhu
GxdUDP28EqBxrMKv8Dl714YbupW5ojbiqC9VRIbGVmfM0reMySB8inQ5x+H/WEhQ
RHzY4wzyjvA8l7re8Bz+Kh3ug12+N3sARdhvgduOQNU8j96b+vW6YbWHMnDZ2tS8
nhtJw5Y/yjVRMdT8ly4FAI+DwMGzjR0aXVObqkvJuEGg7dvhZZ+6S6o+gN0XwgCj
K2s5MUgv0fncfMxsz0LUro2tlfjlpBm5zFKkwulFxcO3H8qb/rRdcjU+9H6r+l3Y
JWzj82E6nbeF67uuLSE5pmhaueuF01xpo0ntTGFR+j67oWaMzMzTBKZIcTtWY8B1
GHQkH3ZNt9GMqMvp4gu3cPxX0llLtuSv1lDNNxGu5XJ1C/1qsU42SYAPz7SxKtKM
/l55nX7dVEHaZzyORvwbzld4P/PXsvTekTeAspkxf4i8M9Rbj4oZoJcCIBQidzp3
u5f2cyQlB+AkOQqxQnMlPme6GJOffYP1ouBDg2EKIKcy5zwzZWDxVFRE4ooJt9I/
C9R/k61XVxqzfcStosDAG7qg4zMjkheR3NBSHd9iRehByK8o5ktTS1bsi0VACuq8
iquMHcPu7B6XJdBJatZ/Wv1KQPI4XMplFf9jaXn3y9kMxr02eTlojFB2jLe6pAS9
SejBKNcM4GCxL91fbuQU6Im2MQid4DFzeyOuhPQtJHz69Oe1f/RhnHHw3GJXAC8z
cRjhTEkoF0hKCtxABabuHmta2SxD0/8FogbSDvmhMVWr7NILFQtUqa0/c1F/Ws++
lXj6qEhjw7+8OMG1NVLywEo0jafKmLLTWbIpI0YCYSFxY/3NHNBSV1rHogo3dKdA
VbTWWfCtlBhn5JAmrwh01/+YlRCUw8y5h0I84Y9ls3riPKprWFl8ffp1hScBrCL0
JCb7NHUmFDBoq5HyG/xG99fDQh6t7k7xS6q1fcOa/Ldzc6r8kqnfntlICoVCEphE
cgVv5QLpHaEGPt0FTbhQ6x/izodTv4OZSfCKgzX4oiLo937gJC8ikzEa0rHjImfL
Rr8/t1Ny1hOqrTAOCPxUln3Slu5TBRlO6rUIAIRlpbARpNvkjGRKr8CZsI9SiMlm
iYMOQu/Q+Qc2QpCHQqPJvKxRuGH89sThg4Us6HWMtYFyig/WD/vzifUKAtTvct2V
X41BFhyuNEQk5Fl20+wO4GwH/V45oVSHWxMRKA9vSH5pEsB7sTv+74/tvIw9xvo9
0iTwOEd6vhw7Gn4KPJApVGqP3JJG5kqzk9THs+vw0FiYKGhsIwADGePhUKKTZEXG
6yG+uUWrjO5wQOt8R/VemLBcBDgZ8kFjdlmql7SR+1ImGlJdQjp9XDWZNqQWlG6h
BzjgSWMgZt1h49o8Emr0+OhHlM4NWs1NA5hbEAcyjXBIuVjDCP/cylkw0AXKaSt7
LTXWQpffTO6L0+m7dMyc2iEaTv091tPHTjp0tQ+5ar8i8D3paihhFYZJcyN0noec
8YzSmCuiGygdAPEa+TCPchTpVgRIwiYVSNGahwOgVuMe2D4AnwuktlG1pjpLku/U
ZNvMQVNQ0RlHxszLVXigF5OY6GZBHUuekXKSQc5cDJofOkXCACrt/Qy5Nqgs+vBc
Q+4/CAKccpH2WxGynUDwNCju9YEgNQJQO6uCMqwSPBk+u3t1J4/sBuNH37iuRoQt
DWX2Q3Wx/40csjBHZcRnevxRn0MrM4mc74cwswELX509pqCmFkjEZPvrrHBlyxa/
eWYBPGBU+/ABNg/OB8YBdMaYS5AdzU/OBzJNW0rNcrKvzN5Et5meUJjVGgbVEI5/
CGflOS4IaxRFRaN/ta12aXO7kWgvKcmHcTG7LzyR0W/JFCrc40EfiFk8DTJ08UYK
+hUk7GmJvAikAcoTEILoT06CShB2vLfKqoGKf+TjUHf9JxJWmvqVDLhAh1vqGxqS
dEfv28ftEefQsLdlOl0D5O5HzPvtQvM1LvgzrEyCvQav9/fsbADqP03njrGaBwhG
KDv1wgWE/1qptKIOt97pCYDQ7/erSuYbdsgbJcp6qqhx+oxa5HV4BfsXtd3FQ8Ny
WaoGutQbj/Y3NqgiqcBEkC8kC9YJMVDuhjShgJX2gCErClxGyunEsOtDO/9127Pd
JGTDa9L+RS63Qq5hAPnWhadxpTijLxnXUYrqpHLzsPfU1E/MGNUQ8HrJewAMWIdg
ytbemf98SeW/X6C5bnmFs+pH8Ug24xMFEhC1T/WYcFZPOU3Xyb9FTXt6uwqkIt2m
Ef7RVihSjY8BZVa4t+FrwD+Aw/qD7RiTpA42NLnwqJYi15pXt143VHpDrvRg6+5a
+n1BJGwA1Z49eT8eZ2rQv0kKzWcdarO/s1cS/0nqPKdEvLRtI3yMtXqMIuMtEHqW
/gh/uw55TO/u+COzmCwhapvman9wN1+T03MeSk7b2BQjB9msdq9q3FYFiM+ZPBsc
bb1l1Lch0O8ER1FIbKaP7GXeQAL9l01erA+253I/DyzQujotMuOYeaDaqcv/l8kG
v7oDvkrUaID+JK6SHE7IoS/NQ8KEESmdY3TRR69zjfqPkD99plBdGjRFHwxx1egD
Xf+tw7sNhKpfB8xhSIPc/pXqSjlC9l2BbCBl7EdGBFDaDYCS153sk92jh0nqXq3n
sBGw8pelB/6atLbrbifAe7rn+b5MSuqkdlCGggCDE/yXiFV+e7P2uHiwurRYqwuM
9cqpennk57IWIhLGu57ZIbBCBavxqoF+AFzWObuZ0yVEs5eMfxcxhwR5Eq1Qvlnc
rQK/VExnoY9f7VGnYu04DdDMK9ltWZG3gqfywb301jSLTBWqTl/+0BF9UqhoRbha
k2CpWNPVhJkqwwNr7arh5dBEyBIlQmM/shyg0H0+oDjScHHB2gpxAvsfzJa9FPgJ
PY4mBos2aojQWYu7oWJ7/7HPitBspkmsUCyUK9fMCIVwzqVPLrXmKrttM/hdRZnT
IZnRNoJPO8LleC/iKuBML8SEskmAdi3g7J9CLy6QdGSIIy0E0b6PwqkMR5TWG2lr
e+QgDQbuTfIgEMMQE4g9ULDH1FRJ3m/iDphNhxJXa3Ol5RryDp35Ccr/IMHnrhzp
6zEGHG2yF2VrIV/oeBVMhHw8lru+93uqxmxehcv8t0FQL6PV77E6mcrVwtHTUtOL
aXHu1HpHfXBEKXwya7xhrnxF+B946qzIPnVLr/S+xcF+zL8yCueUTi+hmXmDANi8
Wkul7+18ImFOyXSZRc67fIZDdOGwNMuR7L+sYQ4mrY0Zss2RvHsrBhTrj9iATRzA
TwUA93MzDhNunBd7olTEn+M4pY3yYdZCTPIPZGE56UQECupmofc1WmGgF/rJ2L++
buOTlJGbCM05I+jHWW5n1LBgZ2QytdkIQVGSja22Lfa4S46HoUnqeEEhcQdTuq87
raRdLxTMy8pyVBL+S3pCrWuJdTL2ry9A19O7HPJlzn4sM0DnH24WtJF6gHL11ZTH
1Vkk4DHRCJvroVNZPbIqBDuZB3rggee3qSSK0dnGHASQvSaPPU05upaDKoJxjAYw
6C/OoZc1so6sF7pOC+24WUBhnhLdL98928Buh/h+Qx2GjDz/u6UO2V7WwU0FkVn5
QC7jpQ+CUr6gF93eHDL0WAaX8KZox+qXYDJZWAhnsylOv5OPmRij2qjpEZNPZW3z
/ksbSJmGOgaypi6RJ4UvV5eNBk/3joW0Z8P1IDDe7g8VyK30npjvpxST/zhDu3ao
XiJECRJdlDebwkFm2ChjyCFGfxxXluQWBWdjQxr7FkyYmMWEeFLZXAv25dvVDoLZ
Z21lKYB8gHU9JvEzUStqvY1/CIiTXFbOn+tfEvLr+np1fVqRRYr31cORyuqRBrlG
D4EgXg7HypGItPztIXmsuLtAhSZUjF6jKIFzMExjfzVVudOK5Wj7BUjl3UlkRGDa
WrNeRduYd3cQjMcoNh4DZxpte8KYwhGrMnildIyUMAc4L/ZBCXh4LdTFqZjRpsWJ
nlefoX9muYqWNXe6X1z7nOLC5GCSESbdYOjIRHJsJ2S7Qf53aHP9xl6lSV8PgHZw
qIxKzUQ9IpoAifTBxWlbddNDN9CSNODDjxqboSagpgLOU1os6FXy1umF06ZfXow3
3zxlP4QAIWIYJyG7Dg+OLAFqLRX7aB/1CLtzfIRxHetvi7JWl6MDSnmZO7OGvBag
57Kj997+LnULsc0zIAM8sqg9yrwMJ28TXRhgxyTxA2nfpb5JKCokvK3UzUJO+ZUU
5kFlGTkVidajJolb9u5MZfcqeALjEC6DiugeMUHZQtBJpAkjmVuJksS7EIK07fEz
jujjTP4RLW5M9ywJEOSDbBNVhSHF/9ULmKSCZmdlv3k2fp72fpngTi4mWvhgTd7s
gq1y5j5TXt9H5MH2pOnHMW0SNyEJ0b6eVwe+l1/LHltk8MRqGUac4yDhz9eER2po
ue2otGl+tTdnBQidDB8X8SQamPCzEN6ITaMAfbSXBsVXBxqtoWgQr5DPtNG+iQ5j
7V172CQO8vqdj2P102fO8l/Pa6t1QCjWjHctOSB/Zs7QPT6JIlMfF35FT10pc+B4
uljS8NpcoRv3NNjRKZY2jyiRSmQl4QyYsBZSwacq1IRAKMCbNSFlj8ciWsFfnKUi
CweRrS/Jj1OlAf8RvgmINmF92BR/HslHpVlRZW/ytZMSeNEAVObvpQuOoRISyQi7
dvoqRSW1AxCmkO8+iKpf/CsX2Cb+3+cO5vxYK5sHHoC2fLMi+FNI8eV1uqdfk6r6
E4WV5K9h93zxDretGYX/fdZvxFg7G0dRoBsZq0+UGVihCjxacrrEE+fk5sSvvdkB
FbE0tgJ92Fv/2FrpGKr680+LlkPKnPAg4ULLzW+jVLlYGXa7mtKYrj8p36/0Yr+t
8mMRuxVUfFKun6GRJgqxtQy91nPXJz8B9GGTJFh1Ul97v6UpPkaUWnqJdDvQHFLl
zBOAQq9NhrLs4v08p83bKw1MphGlqnHb5WhDfZr+WeN5ph0EsYPX5SCd3dzuBPNM
Zic0ZjGcdyRVCebMdfJyWYqUfZpTjpPJT6IgisFPBYzjP0g9IHkpkwLSRwlvDD85
iT61K+Ww/aFQqzu5NE/zZLdPvZtFydv/x9kN0A8q/jf8yZmXaypaoI0W/z98cfDc
zN+ByiboQhAD3xd8gDD7rRx2Aaf8xzD4HlA+N4jC9mEBD8PJhw1X/NUWjjxV0yx3
xIecTcBl9kUT7VkRHnz5Hv2weeND0m4PmkfzduwpRDoTtW7lo31ZNpim9dzebwXr
9Co7PwcOjnWQB+os7EXrOVALDDhTJHWZIvRJOSUkGOyeNf9c/FBfXpbqTHJam6b7
nfBy4ejzRC+RSXx0IN6qw5H5AGZe0w73rNB5OdMIt0h/BwRG/uE4MWwmQS3zbrBc
xlGdq/R/2JQNt+rlkMFDWqc3XkoqUfeofeVPhEIcj1dnS8Md0pypm9P6KjMtRK08
HaXUASdJdcjmyGARttxual3TP0FXizzQhxi5knUzC7IcRxErtnAFbFc6VoHghrqq
qxNxB6GckCAdWeMoRkBiZ+IPGRJ73d4VpgEHEZEez68YNhWxWElugwbOiy/l0VYL
wSc7oFQJzC2s4kn3Xyndv2SstlUSoX6ZEFsh0yahRznWLjaNnInz7MepWbg6zcNx
aAcBnNx29HRYCvn/SUua9xIDN+fo1Ug8jXdl4Du2JpWM9/a7F+uLDyuRTw+Bx7mU
8DGAl+q2XQd+ypoxrD+GyPC91Jen86bjhkI9X//ZJQo4n2og/ZGO9Pr3sPFpzrXS
GsrxwN2PbGkuV02XHrqvzZAU38WUd/OHC5twXeHnqbiTzSMw939fNDvRL0prnjm2
VPu3+zajUbBCzu3Koq9nzFy0QcyuwlXtc6ZD1N034SyL8dQOJK9jisGI83hAYEQc
h8UA/8PthcT9dMMpm1gdaLdqM7qEiMV1qGDstYPu1olg8Vvd1WBuBh8OrhTEWzCz
QrPvuMlim0uxaiQ11BCls9ede59oDXIfNCGXZ+Q7qeeoF5MJq7rA2l0etLRkzJf/
sssFVFa4Fe2huzBS2Ppny4bL6IzKQb300NCcZfDi/QnakmiFaihiCkZKI4LY8xZt
ASjQaA4Yyq83ydD+3NpSTBmY0ojwmUFuoxCJi8BYQagIEoN/fb7RgzgjHWT3HN5G
Nxw7VQZsLN6Y+aasZkqnZxjtw77KjElW8CmivfG5oWSEUBnpcEaLNkRiY82/4oiZ
323aeITg0xH6GcciD1duuypKYlT5WQF7b8VHj4Xh199AqgWVaKgNfEnl5CtSzRST
8D5gO0dTubPap7v2f5QHamzXSB70stBc/GFc3Wi99zOnnQQ+gMaXCDNMTB/AOny6
SB2YUQH/uML06g/Cvdq/C9PfZxTq6BeCsFx0B2QGuxy8NdvgSbqvtGY9dKLLlSJV
sMfMOKCHWDL7TMTvtTmH5pUkx919NK2w339uWmVq2sV/dJpK0M9UqV6Mupz3JCQ7
wszGfuVaEK3w/a61daBoIYNmqXpFy+ABRIYEsQUrLe9vqWsjcunSj+jib5na+mbK
azr4VAZyxDJQyaBBjHL+fwf2O+ObPUa39o+Yg3kFIjlc/CN5pBuni5jjx4i5lcwO
ThrNAIjT3wLaZ/jx5sSeJck2MAWtEzDvSJEBHpis5mqCIJiusLQQsiTA8CVaxG19
rmYnTD2dZ8JXjBDbPC+RByLDZtslHTDIE0baQY7Ca0yQBSoYvJzcaKbVl9e2lVxa
/BYqCxghyaoUiT9CIjkVYblzTwNNJsZeIY10jt/NQxMomXmhss2AKk795BroRwFf
fOTmuvYDc6fj53OxeGbOf8H1+3mdrg1Ggw2nQKdciZh1pB/LcNbixjlwOKykfWd0
P8f9HqsI/5l/ww71WbzHSXkWX1IwfmD8UNNplz4lJTYEGWMeMaT3KxQUBtTi5S/L
yLVC2EjeNr3zfJqrq9JVe09vhJwbmuIEfOCphxLRYq4fbgIJNpUTYM691zf81LNC
swD/DFNLRzPk1X6yyItVV+v+yB/LGwl7CGdXfk2HCHLUOPe+p7wMPQbHpjrEppk5
G4Oa/4R2XmIr3sNKLt0geB3YoU5zcaH6+/RoQlkEmt/k/Zo51EG8f1vfbr3RjQUU
+1k5JGEF0+NIGdkwGonmOZ1t0NBiW5I2+wDovYWtFDnPNfitTYOfczdKMatTzbrm
Qn3kyWrCZb8CO9EC3PDj609mmYCXP+Jp1nnU632E8mBvkgT/WNKnplfYCA8IPWLP
br9bcTPVGJfeJ1bVwoZ9T0HWmoLLUCrLzKqxcLYII5GXkgDTUyX3G0/mYhvAxmI6
OQiwHuKML/nGPv/CgAG37YLAL8YNyVc01zONyEprF9njWu+ZiHVr+iM4bpfKo7gf
SewfUO+GWT3JjdLJA3r1j6DTezqJ1SmyVzEppWNerhFjaP3NGPIbsu0MXY9wlKT/
fn5oU/Ph7eNBQnfiFWMXcx7BK+E2Tx+PXVFwlH046P0KW1oyaw1/SBfmYxMQwRF1
3W+3q6ut2DrVZfHO+mP/8u8c8LePnr6GkERarXmcaxYUoiCyu1S4adYza2Ir3r1p
0aFcTw+JmnBnVGISqHoNx/AYVimDkR8nci0bsUPfT4OWpcWRiKfdaW7VyUJXEkuO
iuZdnEjirqFeWdZpfL9gjNl8302CmCEqWJxk931g37ebOEDi7GOv9Drq8tBc3Ef4
9yrBubk7JuBB/xXRuiVplTv7v+ltQRCA19DzmqnXdB4UV4fbsue79XT101wkmmpW
poQTG1Ph+79ig9UMeOCw0OUrCm1eubrMA64ZObcmHGURm0Mr1bPEUEW3omZZerMM
s3ibob1zb35KkSLhM0aZkaq2K+iL1bFhwVpf07Z6cBFb7GFViC0AL+nSkdmbw28+
2LZvQLS2+yo1H4q+1j16Zr1iJpmRmhQIzcgQopncSgKstHdcpORcBPQ9XKDHGacE
6l9k8UpGLvAxvl6fQI2byNzz50Y6OP7V6iTsoNwUX9aazsE8BXLBMq6RgfYvmeSJ
k7VTDz8ZhjvylER3YRkdq6Bv9z0ViQlVY1gMpMgc9ETQKFQtpdhNoxUHQiwX8Cae
V25uJZUD/AJWbjQAfLZU4MFvgsFP/KHenDQOALh/ASVx0jzVhQpGxC69m5NqMKKx
36FFeVewlUiBuMzaknm8TG+ivDJbyDr5l2SHwHvkPnJSqT/VeFCijYS0dSm9T2yI
UwrTPthTASw4nNzpfvBwsPedZNaBoSYHk82FuRXc7IhBBXpFnYXYp0wB453wL+8u
vd0qiuTfAZL6jPl2ojCVybcFQoQphISTFXt4CbaYfwB4OvU8DtJ7uJKkR3jvRa59
N+nEPWmHVhTeKkYprzVQ5fEE/HTNZRSqkQWm4ot7/RnhixIbvcPCJliBQhecsVRB
uRhFvzTkO0N2hw4ykr2MTYbXkYQFbiro7P5iK2LtkbWqaFfe87lqVnBTEUgSTmVL
3JdUSHXOvUC/sitsHEdkgD9x/QqPIrdMW28Isea7CxMc62LqhryywdlnF8C5iprl
PceWOrKBcUIf3097w/YQNDeQYFLY3n1Jj/HViMfc2pg6utCmrIz8EiuZ061DAi0h
vyEV6QOG7rrPLH/z9jWOvndq4wBVs5VmRSh7SSAVdivdnmrUFh9HWaluH8pTV7IW
RLcf2niY+9+6ZXC4rBSwjXpXHf5+4jDcX0RjH1qzp+uuDlnZb57hggh3c3k65Ebi
rtF7X1Df2HLTUmpvzNcl9nxwX5oNrzoGbDWQ1xcMAhqPpx0YrxBAsgyBf72mj+3f
aEeKrHgvwBCy3/0iUx7bMEnBDYg6HtzXNv+lDvsLaDb+37rl/dQ6w8Hn4ttpSpsa
E6lRmFEIuIhjkRmt8xNXxdekk1t1WnfcWO7XC9d/CX+yAMceBUIyz+WwgvjOygu7
fGHXZ5pw36QHbLBduoNzYt4vNrjpnfwnimIwuYA4wTy1UXT2Rgj8TOh6OUNLzp9P
eRh2v+6rVWnskeOUVstLqmodgrN/+Ho5JL+b6gslNGDOC8g37h0j7dQBHUpkacZ6
1dUS/lbmPiqTOSRbr0zKOBR34aIepV+fmyRc4K9lHys34YjcUEba69wzFegVX0sy
caEPogULkesZXqoAtrv1mmDdOcCHUiXbvIiK5Q3lOejwdKufXYoKVhNboueFZHlp
J8d/Nq5B1J6DD31X4juziZHnU7Ye70fCfEat1+XzV7oMSlYUJIu7T4u565LQri6N
mI+AqPLeJph1U+fJvs5lQqEctH9Qwc9bj59ix9QVxvfKmfsV3xI3WYiEDZ9YHWOm
ytwornAQprTcSkq7+ced9RJVdDcsSr2fx/FEr4cHfv0VWUqQDnYJtVSmykMRBCaT
wSaShh3jCXEcOBSfLYrYH3JxtSQoGczEY+vz2BhhJ1lAU62vMlyl5njarzufq7mQ
TnQsSjG1X+jXmuJQofhmULoWmo24lQ67l9muDiTSajai1LQlsfvtE/1Q+NrFsnqm
rowtI+JL7w+cawy6n3nkRW8ypMa0eD4qyS9xpxb9/cwm7UDCujv5khQt88QlUACW
+nrb5S9oGwddKUtvHwJn5GtxlpQ/oecdvbgN2eK/1ia3D+IHm4LxNO5ywykeS5fB
hrNhhALEztLKoNwLraC0D2k1f4doq6c7Vo8eE/YoYRe3acfbHJ9MlNJZQRU21DnF
mWXxV/5Qbq7tHHfae9lVze7+oUB35ffj0S9rpYg2qcKaIHLWhHVsbCdhU97U8QgI
jM4XYR/B0BmMLdShTfGU2KVSz0d2QAwgXCR/oO+kQxpq1FVapsQl8A2is8PFWhOI
tRywITHd4nzskLwOG1JbWXQJ4c9x7sB3A/f5nQn/fmyDnM6kgXxuyXjq7xKNQvuX
9isWHUcPSi3NROg8EaI37vJCG6JXGFD1AJez4G5PBDJMFNUlkwFtn5ZXZFe9kiUP
/AltWnzS8egZWm44t/5+z939qXn+tlXKtaZ2nGKmiFdfKRbVBJ5YauHXDH/x52zQ
vl8/XFT0bFVrEfC131SdAPjxCtT+XqLpXuCl7XmkGo8l4VyDQq7nl28s8vlsBIjG
+wIlTTcShfxCBlviDK4pri8KuWbBlKH5QNHkaLdQBkl6Ma9VZl9GUnZazevqCyEr
D6ZC0hlQGWaAORQ/TfqCx9SgpH8M7iqon1+YBGOqh8f7IV5NghQ5VTQrx2ZnybKN
+faR20y3zEA2nfnAGGXAasTtdXdIOEDjE1nXgB0DhnNHvCAmXbx/UbIgYcLSp5ZV
F8mkZZla6jFhX3FajobLcGHVKnKeURcCqTYxutN/P+zKcdXoA0vYUvLWHHwscTOv
k2Tf1rQ/9gjef/STNYB3Wxvi0NLXU78bEwzXYAUDt3WD7WydGmKkzsn1c+iA/tMS
ArxBTcAq2E455HaqCdG44He7i4JyotrG5fdzjSTFqYsOikbccJr4q5Tau6Rc0Iye
YDVqXIYVTCrqcwWipZFfjBz0DEZiqi1HAudIEzgOTRZJaa8sIHwwYZWERhwaEnEF
RY77CrkQpf3iEFcf75pT0i5bs9OSv1/r2DEvrvo61knLh6MmR+QEkEif55MV8nS5
eVzx+4up6bq7qXiE6lm6THXz+qbjdBJLFxydj2wKNZ81L1ukPYX/y9TUdL7PyAdS
ocGBNW5rvEmmxxUJzY2JYb3tDJo3p24Cpn9YIC5Lvd3HeQ0T+wATd2yWE1n5AE+O
k1QT8H3vvIhkBdUDveonzYyU9pXNl57gs7TlEwVduLOOtYFSti2GaEl8oT0aosGU
0DmwpySHAQ4/tYNMlTVjo889psw1KhGJLufLzEIVsX5mBKlbMRiUx81p39ADZU+h
YEOCNreA7oRbYZP7NmBuUyZAJ8PB7GAkEpdLAFY1q9dF7kmuJhO9Y/LUFG7ySYtj
F7ZFI9xx6UaioNCZHJmhSpz6BL9n2cAKh+zJDLcWdALENUbbnCM3nGuGfSLY9jcw
j1B3ksM5rcvJJmaaKFGpBjMWEG2j1YBHUNBI69lamq46vW/75PoCWVZH6qjOBDox
GezGIiJQzimcAKLVB9kejQDja3iR4DO00O13+z2KGIJVCRzwLTklnYF9QfizC/hx
mBLOhvDLCkL5LHl0Tv24Tbdzlfc3bq+gonL+meWUbGVMfP5WgI/JIvoYcBl350Mp
+Y8HUpjdivnncmHBRXPoemO0ee5dayZaeyJfJ8kN4K2m9qxw/FcdbP1VfYUsPnPB
i+TUUsLg4ptcG58GBaFI5OitdEgcVPg2CnqpEp14Eb/z4UM6fVNEY9l/9bhkfsdn
Tfbq6GJXfCjj79Mu8YyU2YZhaqu0CbIOlhiFoNcf9a/gQ+vjlGR4B1h/7G0zUORT
7PgkGV0mLUhnLCVtQUFcC+3ZGkdYCYW826wx3jgaDlOxa5qWnhUglKLX+jsSKpJV
VzB/1bko8FXLqcKCiU18IcuimMwmafymQRB2D530f6xTxL7hAFJVFGTQt+egwWdQ
xj/v+0Z2DgsEoL3yTgfjBPyKd/wfHI/6U3U5S3XH8s75rxMTOK9sH0bTu10tT/bZ
mrjBrMa7Ybs0ksM/P+Ca7L0tp3s/s/DUhtzTDXnxtAYIw0cv6rt1dKh6hySIxOdS
vxMe1ls9ebV/zilAMI9ze64euUp/Wrq6dli/pg0XvKZTkO14dFgUGcZNpn5gHYtZ
0Rd7bcuIYlUJ7nq+fUPpaYM1ij+hz533+Yx86oaRIKrN+tJSfpnVPlkbbYYPd6e+
fj0nJh0TrGR+/BDjl/bUTTYIC+e/aq4fKXTPIycKOJfFJvL0wAzuAVJRE56jFXVg
/JGmJEfcBZ079oly5muvpcIDwDzFXWOY0ED0typnO/SGnCSVp57zOkki7FIAp2LR
FKr1oal0Bw42yj8RixKoVG0vD5z7HyQlyPgAa6UxXknTJGOvaj+nf7nwSAJd1ca8
a1JnCnhzMR8/SuUYFTEvNeDee8oD23Z7V6X20idUR2Iq2TzN4XMDxHMLjUl8GsCG
rvT3I19GEhTRvtN6gT9DUlzOJR4775xL0dJps+ZwyRydTrfsL4o0Uxwo2hi8aFfk
geQw7VJptCTvn6TKZsJykXq1EJoFrqKeS2x8AgczHNLwE6rfKT0tEzH7j7TWGLJY
v5pl+9Hd//0y2443fQAtnxsjgBUjIiMO9Z1iMq3p3zI3Npj+3Kl+y0ZAuOIMAO6T
3oL9fVoTCkc4P9/uTATkrCd9eeCAuRMbKeysigGWJ8HVud549LV5IwDZvKNjD6nn
iUZzSITLZweeJAIePaEQaOaT3L4zk6PgcqttcaYe14b6k6XmPAdSBbZ2xXI0+A+o
G2zVaswflS6V+1mR3eUgzuVah07oUKZXYeORGSiKmD7S59TpkoFQMYZItne45Xqe
S1F//+15N5KCFdnookyTMMvCmPBribJSISWO3ZBkdsTQqpW0GIm/vIR1EevnRylr
dgDSISHVpWCNC0qRexwCMKxedF4PZyiIhwxHo32ZOxZDWt8ClV8Zu8XXK8+3d1Lh
SE8lFDkwFJyxqN5oOFJ1kEXIOxxt6BSH2+ImbFXnBChsRt17S+r60ug23BhQ52c1
yFLjmgispjQN0dvbaQdTtBUB4tV42fEzQFC1m6qtd5N6ASg16nOmvg6pRtmtoSjO
f8PUtkOe4gO1L7jTfuoZWDd9f9ImaEpMFGJkT2r7xXqYs/sm479irRN0oh+bHrY/
YwXnhcRrATakgRkZwGrQke8GHWDEAJ5lW9R9w08oK/pOtAhTTUOdL85AvALbXCzV
OC23U6G0ggYm79GuaicwJY57M3o10l8Skch68RdXls8FaCmkkLMP9oJXhhi5Zldr
hNtPeLD8+BJgDoNVSPBSKhfznrrtDwnl03OZAqgKSH1XruVajuDM/otakOIi8vMI
zCcr5v0KEEdCAvHNy3s0+nPA6kCrgYZzBhI6G7bH0V02P7chrfgWlv5nLdoXDiSH
JvkDc9ch3OXgOza2TE28jENwpkdzgRG1ClOdt6AB5QFAExVdYhD02F3/DuzmJVcd
BXE8MWp7JE552SohsaOFp5pCi7aWQyg3elv1RYy53wmgZK1YR1UIK8vgln/8c4Yk
20pzLIeJ02VEV1DRT5kZN1AqKEvIYCZXDZL7bCvYCJ+CxfdWpzlOz6p4JgZVo6P/
2V4cT0EdzICIdV6gpK3yyhMEOl0KRyRmcILhfETOTZGATSBhhbFlo73dG2B5+EIs
XihZJ4xRrQUUhpYAgQ8kyUWC14TcghyAFwGVo8RDF+uiR7LAsbm4xjp5Mg+pYgb8
kceOUbeUch9FqUqptgQ5A15QHKfrQX1nzkqU7MENl7hdOT1u+pggfyYEfi+Ke+s/
0rP4zUeifrkY/gghwalk/XE6M1f8T8RsuFx2BCX6D2qMDXsHkbEyjcJ/OJfnRX4x
ApKgd4CcjkAHLM3OfhsYid+4fozmjfWso1WCyC96UwSkHyym+gNi0ZMU6kWgR4Xh
E3tNmXJrkMTZVL+45R18yUxM97vz7t+EWS+pr12c015QpRKZtiP3h5nOhVN6UM55
irxeS/uXfgdh1Gido1fb4CsI4EOnIXkatjs3BFIHIl4usfOwPnTgTQHpwy7uMkTf
YQuaHKJKffKvPxoL8Of7O7lO/R5Q8dwXp9WX1bCa674l6qap1ySytH6WxMO2FdVj
4HVYcjdkVXzmVFclLMZIfN8cbp50yLdlCcKq7q7zd+YzeoJ2YeuSZvTGRJZVo98l
ZvUdOIEyBrEnX6/HHWCzhkMXcjGYNih7w0CCo+MOaMWzuT98F4982yVGt9kaj4Vv
SyptksE8YSuniCUh7IGeVw/dM7YBVeD35k5LGpbkSpDYcv7vy4KqYvrZ7EUj18Sk
qdWkkl4rjecO/gXrB95a5P532txnloPwBXDh0Mua6XqaVqRkx4+WQ1Qu470viFHA
RuhODBSiF8oaP9O6VlhQMb15ul2pHJkJo96T08wDxkmkQ2OFy70EARrTNyryuK9N
hPgKQrYILVnOoH7jb6o2Nh3Px//AMRLPLFyZF+48634XPeVn5l1LeeGCdBzXnvlM
eWMyMVZHCrWncWNXTmUk1aXyzkjsXsSIU61wjkk6UmBGL2jIXwfZzqQGMl9dTG6R
tMt+1T+8b9LfhoXii+dUzmDl0ILhBOUc+hVLzClgC09UiwY2KX83/BrBbtFpvrfG
9cOEWSx4TkMNmc9UF621bV3b8Tz/wmowbUGtbptGyJHOftJWkoAVyVcj9Is48Yfj
G6v4mF+/PjHEscwboscNQQVmgf/QQTrEbnSAixSmTmZHOoYoZ7IIxp1rbYna7eje
tx4Y1gT5MM3g1AO2ny11el/GuEiqKOvwrEHsn+Rw1T5V/Oj3eoW4WFIRgLgxH7uo
T3/zr7DVoo/ysEKXRGU/ccDxG1pOtB6bvJX0FDo1Qb3pvjYXGXVMirWyjvxUhIyI
UWAH2rlrP4EY5/VMDdryMT2nFrftAY2zULYUv7BkzsgthCZdHuJNusnyhl0TKjg9
zUQJ0vDsv4xSgGFhsCCwpemuzReftDMpyHtxoraCCeRxfz9lgeb8khNb1wZcIfUV
1Yt3g7kJeN95WaiCbXFAilq4dPHPCJvV8gweDunW2dt7hgnpWFnQWCP0PMnXBgDy
LQIntSxDswOUwEJwuZOVTg+qiTY9l1F+Ba6jLtu6Y0cKiqOAwOiVy/0yJKu7HYiD
l5R+/k/YhN6WdcUzw0bnFSBDlyazNKTk93nx6aNaC6p7fOyV4iHhCttdAjmrzWHV
vdq1Xs75OUfQYcZ3Azmk9X8ZahxRJgDg4VqFxpFlR2qoB4Gq32gqaD6LpOmXBJvD
nSM5mTDixlDsVf/ilj4ZKqGU14KdVho7TwW8JvL6TmWBlKKHT14xzdrLaMIKeFqt
II14FiBqwiB2u/qkqvNqit8j5V+EAhuCs63sFAU5JNkpJ0rZgdhC527F2ZLnh5+o
RumrWSM1J7leKPeJYWFfO9/e/vLFaDaZG22UgR2NFMs9g5vQd3d0crAdBBVrJd+Z
uNA7TldpDMuDH/g4dnbFDM91Wc1bvRB3vPbfVubVzyI2GUAgeQrphQJQ7G5iNL4V
N5GuR4pfBm6w1qsskvJ3pTZXAhejqRo55seK9I9Rxml0NSSyvrUfmeWxuzbsI4wt
95v6ynKnhrVdldK+hMLN0oYZql6dxsb3Wm2PZXvG4lM6ojt+OS57ywQwcuM2VykU
RBEtqKjUTzZVcbF6Q8BZVKts0eKlIbpymV9UjYoIUQCj8u9huROGf7mLfu1SwfsP
SJHOOCottgbOrLNh42Y6R0SCBmOjEjzvruxDxCKlb3y5RvxyT3A8CPoBH4Rga+0i
XZ4DP40TkTCJbq3nB+xizshPQ0wpyAOZkSHZXuUjMlqsOq9WqlajJwTmHdoMS1v0
/yA6T4L30Eak8Y+6KMlFeUczm++O5iXbfciA3UoCsV0phzabPDWrAVy1jtFX8Npa
qqKhY0UjHbGRQbyDCqeJ8BAgbD0wWf6+Y53Vlb+ygzyathH9BVMvMSMOFB0u0EFY
JJQapqal66jMfPNHNHYyGUaP8o64+N+++KXsEUT4F++4m3g2Db8kyCHcyfmtHmc1
8Atukiate1fyJvkLbZ3lPMkNaBH0xK3EPxmfL/nAWP2lC+COox74UmyAvPMYl2lg
GBDVhfyqydacMCIdvdeNfP6acZpKk8RyXjn8B8wg97FBDBB0/NMwTnLSBK6Qj2EG
2r4DyIPBEElMV/oL2CeHNUKl1/oA6IWvLAegY8iEc4FwctgNEvoIcyCRhch20Yfj
/4Wk0tEHkZGTyu/pDgHh05Iwqzbzk+ru12Q2dPl2mEVJFNn6kF0flSRAsdgQJOBO
zsu7LR1ZNG50sznHNzEIR7pjuYkPiMRGEV2Y7NcjmVdyGGzwdkcYHyJMj0rkGy7w
wfKgVvBgfqO6m8PRHtu7lOYyEKsa++Pi7bgydZCFI7JB7N9LT4mP4OcLc97Nh/Y/
9pKb8tqfGUtoe/66FZzvuWsgbDIJGN70Rq1iJCcCHeaBV61vTnBZIOuq6nGXyXuF
u3GGwee+SdcO5vdqkvc2B4K5bV6tqK0Lp0xSnvJyJ5X1x7kG4QWnMXMsPZ+SWtcE
mZkrWt5bfWD6lYcucpYcedSsWxYMFZ4sZwQuNDvdDPvgBWScuI9C7cQdUawzKsRi
H7IF1PG46TB/Kc5LcxzL62tTtG0or5vQv0BxSJOHyRyRT5UkyOIAZ15dOTWzYnWo
Nn6FldT2dWftbyDPgGUiBs5hEI6BQ7ESUkC1ZEOup0jrY1hYpv8vfINk/v9ftuzs
6oD/DObkPhjX2/cAzg33scjajiQNAPolU4cM8AkN1DoiOTph8colghRfLMpXFqbz
UxE+ZZMOZnDzmXyFMur+deGZghaBccWKdvf3m1igGdnryOeXLubgTEBdnhY74OSY
uyqoIPFHVIJ2DMu2haEK0W+X0HoIsge7JdNzeZDDDF4JqJzUVlM34K/+CcDS4OTe
a+NjkGQ9T85sZHmeZ1d1hDB05WZi9OJIU8tPQ3b7izmTeKXeQ4OW/JxPugtL+lPR
vOnSsS3ogu1zwveOXdBwawsIk40amkR7Bf04eyYxrB9g24qMTMCmFzDgMDtAheES
gALKPmiqpxlgrIo6wjNPzkCLh7rn31Vomao/UTK0UC8vvc3Jr3T8WsjPlgAOT1xg
jHzkibtFuD/A5mSEW/vDwykYMATfEjt2I24vvDnh+2bgObO/BeCgh4oLsy4T1JD/
wCIpy3nGzGEwaAXhQSB7GjLDbQ2enaYyLQ7OsItjUb9rXh6SevG0VLXxGakmuZtH
n8zejnPx3K1PQtlzvVWasKMDHZwBJ3716UPhnYS2//SRJ722m/svVYoHhPnT+TQ3
TrghDF60uphA4u4fmlNilmoS1tJ1PiplX3PeS6gnstdi6+SGZGd5czzkZ2ZHeMOK
c/mw++D/crQu1lyyfGk/vGMEFzmXBYQ3c+LFg/JlMVc0AKlK26FnY5kO+XC8pEMS
uq25S3HdXuqTyQtrriqXXgn/NLK1GvkYw2rqO7sKRp3bH7FHMDQkIsY4ODoGbH7n
4qAwM6BDAeNfbTawdlA4z99u0x4ldP3i3LTrO/ALeC9g0l03uTVcD1dbVmCRV0pG
K2AYQylNmK/2SmM6HpLbaAXSVRcPrJvnFU/R39ax5YgWC3x6FgR3xj4Rz4pUutsY
Sy//TK5oeHzB31ZbtlW0cUOFZF+nf7DG2LmzR7JFI86l0N3Y8x7zAZLhL0O74TaS
crz0tIOCYzOeCu+AI1ELv0wkmd9PkGB/nHPHKHMQCtAtm+hn8DU403RdvHYuBbD6
Ao8KVtAZshogIoqKK4WpU4x+8m3RA9n1s2AWMfN4r3H/M3/9buhNtJfvJDJa8SOw
1Vr9Va594RxsfnmT+SIa3XWynXHTQ8blqTuq5rWxDBLauvtijwUFC+T2vS3mc7Mx
wUwYsoWOwlRWukQADvLbIAOrvYrPPlASmGk7dqZQ82hY18Q0QQyABJ+tC0MM9Q+i
BoMf//OmzXDYwRtXBEIo7+pbUL4eG5GtVH22vfP+nXdIprr2KDt5EgfRZfhdev30
mfyRQ9LdIM6nL8b74MvIHVTxBiHwo3lXLZGVPb1bb5apy+2FBVFN5vFTD8zbbYiB
8KERRRqt7Pa2RMpiavVWfm7Ej2335JXtMX82/jaEpHVNkDTfrN1nVk8n6onuSb8E
LP6Bdke27Wmw3Q7fPt+IDlnTsHnKmZ6osYvdJ2Q5dylBvqfUKMcLoS0N4nujI/ML
UEpbh47g7uen03mV6FjemZ8As/9BKNqcVcGyV07+fPLPIhV4UjOyV6TpJLHwHMnR
B+wEpPtcN4Cz5Dc7Q9MhAHS/huRNrVIaPHBTONpxjoB1Ifn0Vv99rlqWKTpKTNbz
Zb9KEs7GzJ5Ph9tAW2EmNXkTy+t0i2Cc3bPdGXotrjdeqG2SgNdSGgZV8kn2sw2n
GFGJphKbbZuLj15HnO2NivwzsxkJXUBN7dNhHa8EaDK2e3r9n6SkRpDEiIb0sep5
JqxFR2JI1apMZd52ZHVgRAxYlfrYXi0Ve97hMZxrFZBxsHPunSY2Qjyr6eOfiVP2
OqzNA05INAXPOEgWncUiwQPKcqgJf3yev6Dnozsldpf4M7lBl1G6bBb0FeppB8g8
rcZCqIDl3t8wV+HpQ6zs8SjU9w2uw+G9ROpYdchMAExdfnqmF4/AieFOTQHUrxM+
U6XREM4hb6D5rBGpX0+Kl98nyWuGD0l9kO08pvJv0maqO3bgYARQGYC4Dm6TWLrT
+W0aPm2aDS+RgVs/MsToEjflD4YnTdo6t6LAfe58E0rXmh/hWoo7sXUascoywRMA
9eCPIIALTm170eOVVohV/p34+fT3cLTF6V32oeh1uLZhXRRRXmzTi/utg+aofrcn
EVlg8Tu6GHLX5P8YO1k3LOF103CKpnZ9irMd7BdQbxdPP8jtc4YM7Z9P/SRa6VWW
7cHfms5c8VWd/XNIJgqOa4c+TsftEKC1GzZEQVH1zhgY7SQgkJAtTS90fkdLQW5F
TzRYUva8yMljHY/yfJ5vduqQK8OMNUt71xmz/cvTds3X36y8kAxmZ/ohVlW6vmXE
PuriPteBqcOSKWaxb2fs4kJfz2/OthqpCEwse1A/6xrhTWRTke82Ji/5TfKBv4eb
yXRGfIM0UAnejjAkEIpSEO8eCUFGQRbGpPnsAmMWNVpZ7Mh3O7MgWXxYOc2+CUUl
fsrCa90BuX/Eju8BmSVo70W5VdYZ5V4vzgncsjnAT5swBsJrPetH7T8CjANDk3S6
u000NEGI4WchbSuRhlxcZ8PI90qVr52FXFE1ctDwnCgwB/DXASbyj71hqTkUIuuk
C24o/nbWfTy0ZxWkpa4Wers4CDDjQkjPiAQ0J8xNXhMqCm4gJnTSaBTR++02l7WH
7rqsFHSJaJado2gXweodprCSRC+aPobbzyiTqek6iD9orbIjjLh7KSgW0gGTi1ia
alV4KOqmqU1qxavR+NBQ9w7te46ILGApBQ5uE2YWywwC20BO/Wet9ttwHYe46trX
QzvG2LWsl/8rcZ8UJvLmYIdoH3fETLJCs+F/DuViBoo6l5QROQcnXd074SO0paUR
2wgaADIbXYeOmo3st2YhleUe4BparxrjbYHelQ8L/WhMhpaVveOSIXcbYq5nr1kg
m+vvoLwx60k7ow7GsdpNtZiBJfEuskAoyeZ9dSkHucOHziJ825j4gsOeHbihDl+R
rNOEd2hkKXoMvKjcSMaSDyQzQDI7JW3GDA80sjmbAWu9ERexhYGbp0TMJJ8Djf+v
GRuSywpISSWPX+lavqc0JM240Bbtb5LMnvC9aqhOSoImZ8Av1ZW0+T2n4Q0I7nVV
DJgauhBdR6WU6/7OjFZm/uoDD39iPpV7dwziySOiRuwyFebBZFW2CZV39fdjqkQ3
W5hKcjEg6bE55EAkFXbLCi3WWXfiofFEQAXJEwHFndBvBs5E/I5ZFez8Ja7r/qCh
zER2DBtcmE/huLtep07LYUwBuTUmIQs0kJ6lk8nVTLoPOeL1mylhUFziX4p7k0vT
SgHzY5apfjeByzM1VmfNVBeMpOXyAh02xtiDMPa1t3e9S9h7H5ff2vOhcdaP0Sek
hgt8f39ZI0NQDnghNA/dMMOUASC37YJGWp7PloGeOG0zTGijSjZn6GASNRLARAba
uJGJufQHH2fqrFK0PTmJCao+XWL0gLEs+bDeHofHMYhc8Z8qrM0p2YRgCAmUTr50
FfR7A/FK1WdSW1Bo5DxOO2oaxqY26PKZWklgwBDTsL4oDsiD68j7UJtcVJY9jSfT
XzRR3xddNG0NHCNt+gBdFl94Hu5cd0Je5RsoMAQq6nVL/527rGAcK/cmcY1w/ZCo
2KtvPqp/WUp3nqQWK1L7IZnHda9TK6ZzbNzCmPhFC1cZKDFIynUoLu7D2/DPiZCT
zby8ti0dHJDSsN7XJSx/HSbXelE7NCDyEImL2gbW3VRNGN8xbowN7tF1oWEomid4
JYtRKOJKCfoHPIopUYu1rU+gWFIA54F6QAPHe8E27Au/2pp/y/OJBvReNfaiq6II
7TQc2uGIKAxCjY1cjk2t/6IZTAas8g0F5D1B4vU/hhPn8qYbEPe+NljILZaV2ezw
mR0TIVfve8wRMZ9Gyg5dnEm4l3ApkAJaXMZZaYimvZ3+UvIhvP4dfAU3UHuL9H6b
MffnXotVcbdtQrXPHVQe9crEtknFiPGrN9ukJgFLijPapuAFqlY6MJXVVf+VeQHT
hXX4tltqeRcgPXJ6Rq3XOjyb4Jqf7OsW5oztc1hvZmJWOK73kaKKnXR09wCYwrAa
odd9v4wqrLfjw/bh4xSXN8isNg4QS42s3sXux8/eJ5pcsE24UIkHipt8g4bOWH/P
o4XE5txccIBnXeK5S/FNgwuYX1sZoDGClsxTLGzHtXsK7j/dlllHaVQr4IwXnxFW
jbmjq5HVygq2vuSdp0i6dBMLb72jPWHqxpc/TkiNV68Q70wlp8TF7GhMm+aEneq8
gp3slGjqlphw19ZTXw3nhpCgj3BHKLE8vrd4zlB3A4UEs9qMj1GGFLP3MlwPXVeY
gL8SIalBWKm7oBzXOGbefdJ4tsjFVi4PScTID0uryqoLWly6HS2QlaUIVQyjyUrD
5GkPLTBze7Fmrl+pT9KHWZ73MDMzotwbofBiWrbGx6wamjoHJcMcngPKNvAPIJKu
qsZXolyw1vcWPEuBdb1CLaghhrkePcF73nim5/JL2AsWHn4EQ7li/CAZEwz7Lpl+
I7LRrdTxepUZ9PRcX5ZZvs+oeQS50XW62doyNdj7v6BaA8FVEHVDEipB9N9YieEN
fR55e5rettQP0UHiTyCgX6irNWU7L44xKojSiGKy49UjK43a1jYiV6GuUuEeRKJc
vzGO51AfG7DtwuEnZiS7+o0UuIDbNQIsno7rO752DJSH1mPtWkE9pw9I8S5cbLDF
BfreMR6uk8RqiWriPSiDrwilOGIoMZKwebUNmBJTUhfQvVVvyabBaPPdANW63rjq
mEGz7dX/lHnxk70cnosXNOonYabASEA0kaheP8iOWN9lirLrnhJlFqLa7vVrTDJv
mNMPDA/bZ36KYM+qzy8wQ8zJlSEMINZrvAYueEia9ZHtdNwSjBCKaIQGH2h8mIod
vEs76Ml516FhI1H18tCMiGYzNFi0HC1zb7uwpgUkD3gg4zO+UNhnypMpjHH2f1B3
ZIizb/mHlFKAhQXzPZoaIxSMMp+D9rhaRZ2nAawmXcmJyJVxOp/dV1FVP1veX91l
RinPWgAN+Wazxt4UW9InOejV9u5e/b4UmXJnr9Njg/Jk1qh4Hkjq4lJsyHMqwGvO
3JEK4x9vnWNj049nIwtQ/UcsXCSDrFSmIM68/SHwSxYROVgDVkbtXizcbO3ET+zS
pXOFDUY5IWw+05N+gsYX7b6UwqUS5gWPoDbKOI8LTFqhG5JuJfOHvR30Zo3Lg/ko
Kyw6KuJh8km8nllkIqVQNn7AgnbYn4hCyH/tgbHDpPddmajEWvAUeHPiiU1RdfOt
fkCgcKZwH5p0P2SbL+kr5sTK3G1Ixf/tfehrOZqc/p1QmzeIaBd0ZI+H0Wx8G0+x
c7xSMf00rZzUXdr0ylkB6XdkpLwI6TQ6kedyqv0zxwu8XdxXCJt6gvcOxM802lxy
Fm9g3VvGish9khU8f6kXCWF43ojvd/qKu4vTu4p5C6W42UhuWOLzt/npmiKRUEQH
Tvz0reIRUfrX5LVjxcQALCpd+/bKB4rRTBuVbdbypxPeackyazyCeXLITxTf2UU5
ToUPAnLA6T5SZljQ2pTurAXRt/AGcvLo8aGDzKu7qfJH9jU1QEfWR+j/OzO5q9i2
PokClZY4gPKlc32+SpRlaWq+y21TpHA1u/7u2vgO+gJyP5dD49scoCe5hHwIiJSS
L/5nSfWMUTyKw5AAx9XkP9DpnvTDZNmNjrLTiUgYjgxFYwtmwZ5s3dEooFxxHCsR
9LYzRc5cUp+VnnFBbwPGIrgqdWxaWzaVhsKIn67QQ9CRdTwOyYmuMNdheT0lNSt3
eBBXep6xqte86HGKhCUdl964lwmwkiTCIW7WQrfxiRw0AZtomn/q/FuhXgk+xuq7
`protect end_protected