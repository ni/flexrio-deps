`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
YATj3kULTF7Ty4ORuRfFpnT6YIk4rUPRrM74bVTnc4GjdV8oSnW5PtQkMCLOi558
1V+/wvDfc3y0Z8//ksX8sZm3JZWtrxUppw8c14g9Y7owiwp+JumRtO1zuk5xFbe3
0MMnIxxoTKLhyRJtAxElG8sbx8N21OWDGiOk0Xyd5CqAmk9dcOIbxzMjW/wndBXi
maijUdqS+5KiRCM9+Gsp6k/iEAa2LnYTt4WtjkmDD1P5jZKsiMgFck8WOqLymplZ
ml3TTfn1UlLNm/+zD3SFGP0kABAiUT8NK2xBPQ5UzQ6sMFPd/np8iUZ5u4QLTWOZ
hTrU9OSX7lOvRUo8pJ9vPg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="BzW6NOo8eyBw+CxsNNo4wIDxODIsVe0ft0K5tGuSUZw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
DhjJh9S2BY18dG77XPz3hsiSQ73+w0XqfJhD+f+lIDHHVjOB7CfC8ieNRTexgzn1
5W+qoqOEwenoVQtit9u3XViXJSRJ0wfUC5a9axblRNyD2mUbyfH9+f59nWqGkVOh
ieHxkA/DPprM70F3APxk51m7/gNSLICSvbONgLGndWc=
`protect rights_digest_method = "sha256"
`protect end_toolblock="L7NTNW/5Dqy+2kJZXKczEa3js87UJ8H00YWI+92sDHA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24224 )
`protect data_block
6eHODtGLmq6ccbB074dgNWpdzW45i5jL0Nzx5wwM+RA0eeOHXxEV143NNyQGmZjT
bzHAi/6AyRCB4X9z0c4MjyrZE8GF4crbMH4T59xFHqVrQ4zXCea5w0kG5yvHgpKo
qe8DCPhYAB9sqzbPdPbHVrSYuvsV5HphqvmC0jgRHcOKA2UiPqO+5/jrvjOwtfD8
FM6H8DTG/uqsIKT0UN8sviMI4SJjBQgWpo7s65sjuANFZ8talPYYgGhtCy3/5f2X
td632jpS3pOuJGbJ43MgwXeNv3mjSUQ9zlP4SzmWJXZhtbLOuLyJTISYoLsHsqDR
p9/zSVLotc8M3uG7IoQYfb8KrfEhJoHTECaQ7uMsspgToUZTle0O8zlE/jDtnrba
IfjMAPQLcvUSryOGrQ/dlO5o2UmQHepT8txfitrJl/o/vrmRs545tLsKpxNJO8T+
o7qR0qPeUaugeTTYEqnQE8pVo3YECO+6ZT7CNcb2OAFjH+GYgpuNydN8VSGDtOpB
pXAYgOnfrOX9mYGhMA2fUU44EVOKWA9ofiVaWpn1JHYnPP1AGhiFs4OfdcfAQQF2
Z+b2oDd8YRFCyeSU0f9hPyriz4zrGefR8QjgPFpJkj7hdoNMqAuDFku/AVHnwvdZ
Qz+TrdhZsp1dhJMCESc1ezgIz6ImVtcwwiWRxbVXR+StAXfcOFwtaMYtodNTy8/3
6qsXRODjVt2g/45pGkzwuKJgZ97M/YpQDFAEfJoAhOe/e6iDzx5ZzaGfd75o98Ec
VPydPoCsMi4sp8iriHxmCOC94FgjZXGovNarGukil3AugHooIImDYO6l7Y9Is1Yk
Ni79VaWCWdLU0YNk656p1p80qHExPhn3H3JmWG9B46apVhLJL/7/oohif87K0vWm
1t+v7Tb/wmpkbyQB6uJcttjSTYTx+0JJLwRp6rvRM8bre5rHyer7JnaA7xuiVGg2
MuDCT+oK0faR3Yb3p0naNnMwON4A0So9N27YBZnqyHSeU4iil4Nszt95YnZ/DWiY
TcJGi+fpSdyva9tHoUgzlR0GhbwH5GHGW9a7dSQB+K8mrHGYOLenS9PQ5oYVMtQp
mDF7xw8pkXWQm+BMHt51q5SLRXVGkG6x8NXOJR9UD+f2P2SgOOYJeVNqEmKjo+dI
eBSyZ6sm9L33fqKsfxpj4bOvC7Jyi4xO3ZwSPRwAVUMA51cnl0VqGGSvn1sNIQF6
BjDBTbIUOCLetAEr63+CpIjKgTHeUgqpz6Nwhf0oA7ZLSXMqiMVfrkyUKqh1qgaQ
Vv/cIyOY4KawmqwR6tXeEqlK7gzq92oUmd9n4yAkonK6BpTTVcJIQi1jVHkyxKvm
sq1bnfmQsdFV/0q3TmSeqXdWdz6L8HdImK1m6bIyEJnFsHQ1Ma5pszYYT11hIvN+
GHkuR08MkuhZRW8iz/a2jGngDNtEw3TifXAQ1RGltWkUSPe3RvcNWHKcM2nbkBGO
cyCEOwJ0psm0jWtH81OwIm/8vdh257xbCNA0PhjcOrf9ED2EDb19aOV0qOTnvq0g
QGs/3TWoPzVpkjhApTjeZAqfQMf2e/Rh9JuuiDPBc/HAOy2Tj5KkkY/raLZRItow
p67rK7vhExo9XVh/hOtu2tK6a1xyXdWRPP21LBCmvtkcx6KfkfdLmiUMF6Ld3mkT
EhIL8KKxor2xCcYQHirE+rldnDSBvFAZ9DLNwAJDcH1+GXahTVQtpO6Q0qY3zY2M
RJeAwtXScw69a9FFcJuR6Z8trv01RtMbxg45q06GfUhhOlgdE15UmWquCQRVTed+
6A3JrIIjBBkuQ3eCLj/uI0O3SM2EoPyBGKg8cqjWTRNf8RhsjjQR7U8i2IzJUfj+
40Tz+mHJxUteylM7St+VenYKrqTzH/C/ZOfl41KYkNKdlEXR6SpPSaPZwhiUjrf+
2MBz2A5fDiXJTX3WOAV9KhL4jxowFfInkV1bTyc9PIesIybiwIeMqedEopG3yB44
NkpzdM/+vj3KvwepWdcLjL7pgl/0hEdd+BCfIM48FgLf1wTHvJK4C2Istxecvsl7
OoQIIXQApq67M1nuHSF5/IIp0qHVeoZgEqNn5fPXHIr0x2sEBKDRPH/JXaTbUx+Z
/OBzNv/thoz2HJhfTon8uamGSeyqmH0q8PDQ1YCupLRyntnPg8d8U3x0puVqrane
q0RPqbHJ+4cTBoGQWL0v8DV3JxtP4svxipnFiejn9yDYTpL3vDAszpa6uGVQGLxh
gX1i7B/6fLVzcMbou4XgwBN66mz3XE9xquK9D1+VOXFsfkBSehOWTja89q5q6lTb
JBWVA3Hl6Q01fsng8P/brYHRuVK65XEk4prZ6LYHUzuKM5UtCLjF8c2dLOZI4LH1
IGwliLTfbhQDqxmIV821PoyDlc2WkyJUzuG0UfJj17mPO9t9fdttOp44N81c8Dcn
HDz4leqHZ9Ek/nrSckyibdsCAEDp/aJFy7KOr+Yx6jBkqPsUTKAbbNhuwMhBIm0c
mAcYLtLRJ0d8Wr+hFk9OaVYKDuVKZu3LTq6JIHmPAHMGaHS3PjkdeWlbqI4bCpLq
9CqGwAqqAXyv0KgexwNtrI9eq3wk26fh6rIIFwN4TL2Zx9Mn2HKEakfnLbc1Rx3P
wsIh5rnlkGuN41w6DB7E5Y3rTQdU+4b543tpoUqhLjCdsBhrfrKESIZ89pbuaxCr
0Zv3kjO3AZmLOR09HjjaDHaMHgDRQa0M1HCHivwtcsROiPzmR7S575dEGZDMnOpZ
teCTomLRfq66qJvjOYQv50OIsa9l90RDl+9G8T+C6x8qloU1xrek2OuPUrsdgeG2
1KTGz1BOVzmndDMIK/bC2a1UcQVqd/yHqZBnjMzdQJGJNwv/6qsrDr7NKZNGib/x
lEwyPC923QZII8gJpXrYQC+DZM0PTsViUPzeB0PlCmcCSHrW2wf0jAHgVXs7sjYj
EXcmgHrD9AdIrnqgHvho0KSZUHBBcPXcgx0ivX86MlukCQpZh30FZ+MBpWJtqSgy
GUgmsxNZ57JtLattfO067Xaaqq5m1xjmO5M0XB3CLuPFuePQn4d5GbdL5C4KTTeg
bZ6aC/+Uu+3rOe5r72EcidGFZecv9XOD4olhpRPB3B9ew51qN8Y9OT52unLe/q8f
ED2pfqvPLoJc5EXaL1jswMA+xLHhjWC1Eb4qLMK9eoAjMtL4RimgZ5ZEe2forL9W
y4/NbtcNPKMA575bl5/X4nGGfcPkN6qGaDqIiAQosv52kznPOE1QIRCZqIT6ZNjP
7utw5oPhpdd0feKuJT5V3n8YhEIkobABfRjvtY60FnwUFMmd9LHoWqhmUrL4eANF
7OSh2NmiHcXR1QujfxzxRWrYFrwmQmijIhw/rGZqJhi74RIz7KRGF56ZvssZo2Rd
Q9gZWZ8pNSR7DZLu52H4Yfz9fwTQq3aJGnlkaTS1PPBMVvWW4mAVDAFgaPxX8yjX
9J/zr5tTbhww/L7VvAal+iS7WFeeGXXg6hZ6vrmrKPFLD1v7lIK5kSMnlwznaLyA
NAxsvoAp0eenn1lMx3V2NQxIl6hanbWKnBztVU0eCHK4xCfLO1ueFSM58ORp55no
21wUaq84aS6gRtR13TP/V/bsZltf7VRhFR+rIbnxyvWp1SpxShjZXRWW2Dncuv0W
R/+lsqYCOtf6UxC6+8r9eXjca87lwEAXN42is/cVyT014Z/+DF9r2pc5pYxYdB6w
VO5LW1wexCb0+7Xsar04o4Oz94WbQ02dus+fSvtCeiT/VX6YQPpohFc42GUfYS/Y
7tY5+N4P6KwuM+s12gx2AEblBiCMXfLFzFw14vfTZQbwI6oYf9aZnzC5Lv3DWUI5
qVY0lN1hA/g6q3MRHtIw6LRXuzpP80koI4KNsX51DoEJhEq9jQk1ADn/+JYPJPW+
BzKyy6tX6npJx1L/g2kePkLsf/I1GH1sZDr9IY1lLOg34+ZHafWrCxfHzgQHz+ta
wUTXHnu9QLQSU8oA+vB+Ll7jhYBd06zQ3ZNbItvKkwY+6aeYedJ3HVmVeXARVKAV
dAHQpB8hVw1AdAk/Y7bYFpVOl/YhhoAtGkd1aqdhqUHGoJkG2wQ1k0lt7WQrhM+9
hPc3pYnoEPC8Mjj2jbmPthFB8IuzZgNSzb98YHTXcixpLxAESbTzIPurzEsBGvfg
rjrJMvgVTctx/nLlloz3BCrivd81aQpphpYg26ZaTPseaw5PIQ4yHlWsVLrKPPgw
V4ASOGm4QME16YDR0znZSxBm6+W/unGOQJuFM4/MK/bAzn8kpgtJrFS7spXAth8j
HZLA8KXI7NoA6yWcIWrmpzbI34dXXZ8nnpHmwaKYw9d4g7mA/qeteLuHErmfTAwL
i2v8l5v3Q27Dp8cHocafDgNGQMySYrFT5i1q8IwCEE6NN4kT+O1nS/Gg8itObkFi
BvGKH2Y3cFE9OQ8AXQyZcBzv8wFy97/8T13maHLnX4Z9b3sUVzlkpGxck+/weGjb
o4x59psL/afa53Wfjd10kOVFlTYEo22ymJHJMJ0VlBQd0OTJFUSpTyQt8buvRBFV
62ONUEeRUjMImuCjaPMS5uZzfZ6kUH7//o6EhXnL1HCbKeZRIKIIOfaurhIvDFKF
0y/LEpBE4R12sW2a0YRTHnj8LWi08IkKzEAW40CRygkdrPpFxc3zb2E0Qi6/5uFD
wuegjBrHBoXKo+eKqZykY5Sf6UUh1XvwVAuWgrWLTwGZlJix/XYh9xEzmtn5VC2J
vq2y5kfpTja7oMx/uXlARYCbwWeeQAGnwY60pfTtV8qggaGLP/kV3IEaSVQGuaa2
bovEq75u8J3e/eYGijk1+lgrLVvKk0N7KBybw5Niq89Uf3jsfzPU7FsKwgfMymuy
EvvO1eEMwBTFSRsIpadXIqtLezeACTnDgcdnVtf4gUYd3nbFcIEo3dfAD1P4eocU
mFiTX7JjXeubNFZdOniFBx+kguH+etBypCxbfsS1mVyvSaHhgepOliSdKUhNVDHz
qokldYYS/D1Q3NPENVQrbSzsdSF9i+Gdhf1kraNupOpZnCWajaKXmywLvRMaMnmk
ZmBEI+4ag/QCFqjJW1VsYrSa3cHm5V7+9ve1eukBqKpCnVwDh4l88q3hz2T7U5eC
ZO7TAIQPx1a+9pNhUnhkO7qiSbaY2HKDF445PFgXXSklQ5kayBXW8g5VQlihx8ut
oJm4XTIXWp8ocmnBv4vAfCkCP4Mqgff9KoahFgAWKK9kYr3zit+creqo8Wjowrzz
I2nMQdjt33cIEBn82omV5znwCHt8iP3LunYx/bl0qODwVgx9kNaJu54i0gEq7mke
IYNm2ooGIrXL7DWQluHy0hD99bhefu04g3IVqH1/asBoUWvA/+cOj1/kYJRwxu4C
85ifrAu/604lNT458o3Tnr3s8YJ0NDVWfLt3WmPxt6/o+OA/WRjIZMrLnyfVBgFq
t93Eu8IOB42zmGzqh9xsZ4B95uicP8dklJGtVdkSMctq++OZb+7NUWe3a23GG8EF
Z2xqtYtlYdDKAddEmd/2QZaTrNlsdDlgrMstMz0o6/NkNGpsfZxJEemjym6RzeqW
VaqUDAMA4u+w1RNe5d5WybO+nDx+84WiRvuBOMMkws6ztURieY2IXFCydB0BIDCW
952AcS4HG58lFAf08Q0kweSuQSkwEkgsMrug8cCchmhGuLClTa1kHccP1aoVHEIn
8azZY3sFzhks/Qo1IA13pA/eQJGoEiGo5CeVPDk6KN60aiik6xRY7IWqikHLHFG+
4RG8vXuP/pp5aRTCMaalFxuU1J4au8pEtxt8+BaMFpQxurMsqZiKg0Ln0FSHr8V4
GiwzfIsJ/DRS4CXO+9YWvHLoMTYzAvKVbkO+4I1+0auL0MnK7Bp21l8jqlo7x/oO
rXMjLGe+B5XMG752JEpFcBhhzboy85rwe2XQ59SZrHSdJ4qdw5XJ/HjIIGN1gQRa
FO+xw02NJxMXdzBMb94hgIQ7GhORL6h1RewCr5rZcKJeZ/gYtFE985AlvxsHJpE2
3hgYpnakRShKzz5MobM7UOJ3JyOamRKTomkkfYaxRUnafyJ31spKY5cKyYOacdbN
17N0o0oX/hwlYBdN/Y8MSpRgnmBCpRiGFDQ7wPRH0U8W0gKxnuIbo0omGmw0x3JZ
X/OmAo5SFbmBI31D0FbVrXMLSdezsBwU8oEDbePqLSWFQMxbTYvBm4oMKQnVV5WL
5Y+AiyOnCrRadW6XqfTT2yFBcAMMYDp96JIx0juWQ6f0BTDSyzIhXyAuU4iJSZXd
53UwKkTXrOGLvqd4ThuoeRsI+6rdrncr8M/kmzeNV32REQGaNYyG9Q0NX10KADsV
pg+51mTonazBjxWj6czXp/ys0Bv40Th301JMD0lltwY42hIgfdUQyQWlMcxkWb9i
lKPRB+PGeIzy+6zIGr55eaiZKuE5b7dPn2iMmQCdxxzYsybRkLR8BfFAvMPHF2um
tVxX5ciRw+/z2D0xSoN+MtWYuqUTxKfM+KGuFrdhtxLf/EmKVO7p+yQ/LYei1i1A
d08JbmIC9oJkxwswrP4BDoR4y3LTyDEK8GpU5muD15yTifzF3raw2imwD+Imw++h
IRwj6+aDTse7o3K1HHhebQZe+aZNsJmoj0sKwPUzEPhopebGnAjXgLegQQQqPRfY
INztuk/u2iUqlqiHsm+mnLYjL66LY5ostxcxrSz8Do0Nvk7tlMDR3whbFxxBAsHl
+PSUuPkfVKF1PEHmByvNYF4gDQZ9GaOaV456XK0I9w6I/aCxuUFbkhEeifzvJFRU
CH5pbaYRoLEYLIwi36P5nmUFgXFd1rUqKp4dPDLClzucKWeWAegJYg57M2mhzHZ7
8adQtebzBjwVNXRNXG6xzj3CgXn2cEt18OygRzjzFcJ9z4qMHfeNR4k4YYdc/8yB
X6szMDxW/1u9AWe/+8wh+6xbZzHrPGUGJz59ftWWkhOhDNFrsdltNPfQA5IepMTb
Nv1wfkNsksdra7YnBaau2AFPCLkSnx3P0QnSektQx8l+MEiO1UvL2HHTdGm1sxf1
rIW5tXxCAcuP9de7hgXKLU/7AQgeR78DBptHNGNV76VvdP0FL5wcJE9HOMv+7EcM
SOaFS9oUQeYyud+RXf5FlG8G/jN4771y8V13fOEPCWD5Em4LDYOvh9tPOdNfQI2/
v7mQe5tpyW8DOAd+xpW86sDxvbaCuRDGLLhVIKS5jBo35vu6G5krFVCWHuKVxO8D
l9uJoxTbDimXlS3EJwEPrYE3pCI0skaccDZQYiaFrh8GaTB4/v2rS5ANLPeanDeW
NTyyFHsqB/wJFZxhtSJcZy3MpyVOqnmw2XAa9JvnP5bwfLMFykqrZXsfvmhNV3Ks
6yN9d2Bhr4/62xc5zhxiaYRboCNTZlm4cJAgzPft+y//eXkkyh+RgPoL4K/CG81Y
NZyrgWGh+SC8orODD5WIvilL8z5j7iEb3n7F7wAiTrzfpspq7RoaaOdEEIV1HajS
zzMOWIwjP8syHmKdheFNwQ9eJae8w884/iHB2oFvtHAJWvaJe9H59480BwXxT5QX
Wq7BfAbBDUKeVtym1p4NfprbCVxKGcAVgeWMz8c7Bd9EzY5JfgSnOO1Cpozf7SCl
u9q5juDXnNoyUi+JMy6O4LhLOxIXrFSE62gEpyBzLJdRPEKXKqvSiDr1yZA6+sQe
YE9JV248WIp3zazAiZI9MHfNVy8XZwp+nEz87iL5NSUiPzOoHXYeoI0ump8P/uyk
FsDuKGuLGv7VWrPf0jCzWE6gue71PSov2FwhFS8L9ecD0Zv7j1/nRTOTkKyyJMVB
yEbSfHK45IdbZ719z47RBtPkjhcC1BbGuuQiMJ5cJtsf91breK+hIQTDIcgVFpVY
NIVomxHYHXwR1m1cXwx5S2vjoqfS8/sAxkZ0XfSVZBI7KVnLjS9hYTZxQaSj8Dc7
hUWIwMtfl+mQmLbO5Zr0/htCvv+aTFdSBBIzjn7A3ZDIH9sMV7EYyBB1JkBRVcAg
PXBRPrSr4hJQUJFwi/injApImtzgW/2uwLP6Uv/LJbofiGuIH6JP2/37htyVHTFE
+jnVwQiy8GNpq2Gc+inHa1RAso/HIZ55QTY1IHgaq6/LrSxFFEsLVnoNKVSAdTC3
LaXpV+wQJ+2MOMiZ5rYwmhNAPTPsv+z6Pbxucp5k3KEJkjTx7B0X/gUrObv6gCd5
N0K1Pz8yRXOdmWWcOHCb/uzTRg47fgSfCLqHzbUcSoY8JN2na64kYwX5zcf2hkmf
bwW12TyP4V9ycNytIfaAoy+LXzas0QkhcFJCIr1+L8rBtFxqF8FO23bjGqFJFlXL
2vFLKd7Ppa1hB3JoCu0ahI2O6lhnQVo9pY2xxu/4oB8xHSiXQuKP+gZVe749Z9y9
IbSiBZYTdXUsOnuHT/U2P7FbvC410brlhsh6+80fK9Q5aOVbouYlasygCB4HBrIH
66RGK8xZtJOfRkV2Fjor4VhGHXdMo5iXVlC4GSmfTGja3r9+A1rBFltPz8vcBqLK
CxA9vJrHnTflHNvj/QIEP4X5MA7+FbIcAs5/S5m+0KsKp9D0K7h0JBr9efxBNZ9M
jtmjLI/AvijujfayHIN1Ep+9sOHAqoGOkD6ASAqhu5XS5JSyjLhG0bTnSQxTkF7R
8QA6xN616ceQKa2iSnbxI11Nv3SUtNit0vVTC4v0xBygS83LPEE7vlvtmY4xEeSs
Sgz0tu3nUri1TKP7hhgJVy3c2zDNNPNhRw+kP88JQwlgNDDl7rqd1x391jKMoFuv
XrQcRxLgzC1cxbh1vSAfB/Ewf9hcoZ0ykcuTrR4POSkZYftvuBn2GMhvwjfUowvv
zWj8kDhkp9yZ6hlMuYGjUnIpPKJYcXJxhbsjv3KqfVAnQ6KKMH5DvjYqc/NucfHz
7emHy8rLspXJguJ9cmGl2Y1MDcawsvlNR2NLi3EclhDEblhOQBBOO3PPgHG8vz7c
dzGoZ9Nue/hPiXCFnxH5GM432/ZPQBwfvAqQsADRSsLnJg1UNuHdhbWmMwAqkhSz
wNf2dQCNFYEmyMe/PwtvY2I5Zkb8djBb9vOPN7KKMDrVsbsefQLc3tYkUYBupdDB
XKQsJU+UP5fVt37Fpukd4+sQ/8Nr3D37Aam5x9iAo8s2FsQvj9s+EVx4RfMGKcVZ
CRGU/Cy0bvrAJAodeV0ZodBoJoQbJlU2m3QT0JZjl9tL1ay03SSLSnH2+FxhYqYX
OQQTuiiM9jNtaraTM5A3e2IwOgHe0LoalMbKGb+ugfj40Ri5x6oTTp6PUcwMbVjf
0jpTW3fIb+PwsI5cnaG3cHWl0BNT1/ioeB8f9nOA/+pLf0yX8NvASqGsC/yxOZK4
9t1qLDAAzJu3H0/jCjKF4A8gidcWsrP4bD1MtQwB7PoSM7RQYLk8ApY3qCwRFgZj
cVVyaj1L3w/21KnYyk7M09mqNfWubCJU9JTVZ330+OdCGhBNXRpOg8y+Kk7y/Mjx
CveLEt8Xp9JNsiRzu7Ip7CRPs6p4WMfzQNjdDZk3XA+fhZRcCqmKmrPAM7KMT7kX
wekl2yTH607CadOtwZ7qlnWTzohgYR9jqOeh1RO4KG74yldMFp/AcFMprCrPPVgr
ORNUatER4meZEmVbwekVeba+Qmg+7amXfupclYjNe5H4PAEWxgY+JvXo/olMwqHN
wZ25OiSnvzFzBS9oHLw/DTM8okbIjuylsYDDJbtIuXzIEFBRyDwvpoNYWUj+nDjr
+PMia3lkZbHj+lUOYR3cizUt2+5C015wQ174wMq4feQNPZvju36eW2zyG8hiIj0g
FkT+3YtmHc+IffvUghzgOvsMjKn+pBCmJG6rNO4rdIp7HesakB82muLNyTLl9ArD
4eZPf70cvnHktLk60vp1IuyulOvfMDytDd5D0jRmvma5dza05T/4Fg3h39odOkM+
mjU3YEG9r+UTB6cK04UsxNkgtZC0H+1/ldiOyX08YPJwYmGgQHmJyq7uPPZVe8Qu
t2VH25SEmbt/30Ph0Jxrw96Rst2gbdyNtfvX/fBux4M6IZFe6hGgxTOLJgasOqlj
mX9MESfRaZ+T6J7El5eoncvQE7ewaxsTfQM4yvz+i3BSUj009EFuprwDEdn7nfdj
MdCVF/3QmyEYXLmqe8jcZmSTMhUdg/pW2BTMr90HxdPnZ/Z2YRXLzKLFd+oR4U9r
tbpIZ8vb1ZX3a4k7ab2c6KiDyiWNwUCvhGY3PXT6r2AGw/LpQA10E4HLxnp/wTTi
JHmdBE793eFMfolSwaPEduHmOovvRK6Pmk9ATSR4PGZlmRJEcqJB3vcpnopE1wIo
rfHT7KUcmhE8sICiE00gV/y1GuOBV78PsUrFDolZDr26LLEU2NsQK3FkxdT08pVP
K76czjyPARKMwou2LMdU5FWThdBpYE5Yn2Swqd1XuIX9YemL+Px6G0GS8j97CRVe
X75UaCX9qwnMO8XH1KPCikRAtI78z88g8ezUIY7vV0nSA6VnQTbnWV+u1BFIiF6e
8jKJxpGGtK6SzUZWkvqY9QL263q0Dnw1Lz6p/VU6x/qaepLMLtEks52bycJ2txLu
5LvLKJQAy2KeNnGeKrY0OfPGWOG72Bx24cMQdcaFvwHtvHTdPi3MQOIwLj1/3mZZ
+uio2s6fx7R0KKjUci0fqVB8FIfzb85ux0ASN/NwegIrL6m5zdc05ceoH9SrnxWg
Fj4JToq89Nq2wXlII6moJ1/cjMXX5IuubH5xjUo4+HKq94m59SODn2/aA29wdCaS
RdWroy6PPrYb/EW4eDKtBwIusGsrgT8uYHIJzM4NurqyxJqa0/NK7k1UkhXZUgHR
ZaBzhWL7bFTYrEccU184P7QEYHD3hwPy4+qg4ZFaJ2UZ6AO93s8AmGhJwN+K/GTx
f/nGK37ht+9maeva+R7jTfPR8pNuvDxIhwEkyo05TSLUFEQtVXPQhiVEWGszeYcs
OEnE0HoQUDY4Ctt1mFEM2EYNBnD3cM8kggvL4vD9bSpe9oHW/m+Jh6ReCUecUJt1
6dD6YGWhLUnUsHYgyRslVHOR/+tPOkq9qNCilUxz5iLjjIoyJCWkz5Amv0Uz9zax
LE2MUtQJhEigQ4pnTWXSbyutuoG+2wKBBbQqjq3cGgtVbCwOHoYdzYoUuC+HpLjZ
C55NPPb3j/PXDfvedyPUG+di4k0jaWRXoJhFp138pBsHvwUuOX/2RtfRZDxqwRlJ
ul/8RJeveEQ5hVVNMPdLQjs++RucQBmQe/fM55PFORo8Rzr0xjCbXyrvPVL/Cscu
r7QFGjBcB5LI/E1gZscRaqHU9l4+ZkHeY1MJ37bJPE4luDBt24n1u0L49egzcoEM
4eKVtfGAdeqVGFUQNawM+7CZuMftZ4x0VzMbF678nOVWB2uVIws0KcxgPcHYyCnZ
m4uSAvIXKf1Tk2JPYPcIAcqR4Agp++wTusNWlBF7odb6vFibG+VhTCC7YqR+SPBF
uQDi4s78FinrUzFMbFdA90klM1hDJSK8kbM1SbZaouXu61XnV9nrQp6GTl5BWpwd
H01pKZgdr3firBxIKgV0HoAixoolJGtoKo2NLbSniqrKfNq/K2E0u/FlVTAL/RzI
LfrPVUvnP55xNErxZJagcFnHVTSYTL0x7HR6Xzq20U9UUYzgMBZgyJquKtMw/vUq
CRpx2ab5jo6TqFlwaZrFAdgtlNQ6uR1BezUi6ggNaLaJk8sbCKn2kFoprcNQTeYo
FRYRKlEzwGuld47kP1JghtpagY3yCqTiFbEitaEu7F2E66oyBXnl7894Wq/9WyOU
e+G3/md2z/SPSBJlcvwFfh6bzZb1Tc1z38eGPDDO4n9FCH6xK565M33kuqpa65JJ
3Nzzi7aCRDQry/V/J0ZI6SJRbSwTKHZHO166NX/7DNm5g2R4RUXs3OuiPRUf1k9Q
xS2KBoSX+P+yy/Z3LlQZUeujdabbxvjhN/uYPR+CEvGTEfWHx3UUm8Shwqlx5D3O
AkaE787GZDwRD9BkN58cRSDxUzrlpFWjcTiVQhLD6fAig6xJsa+LbIwyO1rYMALJ
QW43kk11muvMyCIoTZoiCZnlhStKAGYYhuKiggiEyXYkV/80/lqkoMk78Sb3r0By
TrccbIwL3vZEyWC5KtBpqsFnqXg+mRNaZ+bpegSRAmHY/A+gVzKSPlrXSX2c7kFE
cE0ZgLAb6EuaVCDeIcNduJy4L6FqTLBxbdepDZ8PDnleGZFL79aYN51/Twuku2e1
6bWx1dYQgZ3EetHEB+fPbRd0eFvFdUfUoZkELMPeIfvFFP7pBOY1u2k//DYWwvJC
RTN+YKP5o7dvTZpIhQiBR0DlnJSwIR59xj6VtNdjDyPKazWEddhWagGtF15fh2Mj
MwBhLbmEh8YzfnOJC4hYx0soF9Z9JQ37mjBPl+fTuvXdEo/r8DOVwQO2NbSnGPPs
3WewU08k8sK/t+QNg0sZuqh/9pMkNfJtkvR4esDaFSUGE+QfHxG3n0rFR0I2aDSe
cVgbOZqeFKNZ3wdkdNBUFbi+Ol6yOs4OWV+qK3NCBo8V6JPvKyQiQMe7lDQ0YvjK
iW5XI8/IsuHlqGxdImkqlV6pVn7JS230tAWHyvl+Q6KIkJo2h0JhL2zf7oNW0xxQ
pUc4rlG5n+WCN+ZbuK6p9v9M93dVn+6eAtenFOvjFSoRmCxcP7GjhVH52eM7fyFq
f62WH2JGQD/QB9s+vo/UL9ZPCBvRrEBW0+a6Q9RezBj5qTHGd47zXOYDbCVKl4Ig
h7GFpyHClzgWozxEXWrTMFx6W7gAM3iOEjdYbLG/fZca0eUSQzSZgfFxrdk1zt6K
1OLGPz1eWpjBXbX3tY58uEKGpz4Kd6vw9uxUbfXC4HL9e98xEQVdE188I2Tuv/Mp
W6++5bBQ0RJCNJx4Ft0h/6Etr0TyR0sMjAAA6uuGAM6N8ph7SdX39o21Qz1Sf5hg
sdgDYS0ozwLguthbYyEh8AUYq/reHUkX/hM3C8BuAGHTG/sj/QMbhbgZ7W/MUjqk
poENtOsrOFl+gU827es8uUAbKFpDTDHtXIfpIwlWMdovSgFL4VMu+HYlDwhZVv+q
Fw4vwxCKyP8H46KriJhrgqpEf96DrXA1NaFg4unYRWJmV/VqRwvoYVwNPi3/XC7S
1rxgLEJs5MwR8/W/N9yiNgPYWFKnKpXpR0S9hylJiI1vSE8XFYwlZmexFI/IN5AP
0+qG0D5EqwFED9sN9AMbwX+v3eYJyKW99naCrl1nLXZFR4lPJKrwyvdcQnly0Y5I
dMN7XUkzNQSpjtG6Gtwc2DUFjza9GkvGpZCd83o2+PQ5EId5fE2kZ1snBrfmFClq
xKYKvvaAshOpgDQUKy1SEAIJGNjWH76jIG7oWMXH+8bAxsPNJYUTcN+Z9c9rE8Rx
n/JExuFOg7FWOcLFIrYaaAPWPBpF8BCzeYfy8lmpXs+pZmoIhNdz716j8vuMdjWO
j7fNANKAYvYgf6oIphEC+bOIw+H2FQQe6Zim5GBya1fV6MXfiho9xW4NKoU6wlLs
yKPdLobKiKSCD6SCnnQSU8v94xs033vWnLNWLtvxQPY2qG4ZwJcgxrHjVpoywpA0
7ZDohMsD88LoHmHAhS1rSMa83lqJJAkeRZVE9bYHUOGti/qhdIevlKZELHlUBFNO
+nRsgmm/gLM3QzjHbcvXZZWaeYWxisr02bKEFC2JgKF/9/xG7BOvewJnkmoPX2WN
h9ywokRHSxtKnkamEY8cR1VBMpfzoI2A8X0502XuhPh4PArIeWDXk9igl3vK10t6
GrZnw8mBTe/gvhRDqA1Tg/YsXxGPQCtKp7zwCHmZs2Xj2reTJLWiivmqtiBCIqdo
RSEKxjHRCNq/TujIqf2mH0Z0Fc4NudAwAMJjiLUKiK6FCafS11MFRGD1nN91D5R9
h8QG9CEtD1g2YLx74aeR3Keby5KE4eGPbesrSt1Z0V/4qWBg0ElhVRVx6hrycBSL
GKme3Rp3WNjTvcBmLiD2XdMrTU5NlCJjFqSggsBCcGe9bXuTMJrkJ9/28TvRzV7w
hnFzB6JWTEVO3CkXRhpFt2uNAECePo2BXsfV6yZsUmjke8TL4aVAxow3MBSE9hz8
byhtw/QqlvZw8BttiDucEgYPR+PmXYCFarOnVCNy23pfR1C4B/wpaujiJj5lPBSf
dFZdtUgCS5DFlnVK/77RzdrXaRpQ8bTFpaXljXL8EfA8OoBLp/x57B9aeMgu8FSk
r6isUUGEXu76WeJyaiKFHOLFNkjBOfmbKRcvQiyzrzSBkrpA8r+6e4A7qquGtPht
KkRrIibVUYkx/CYrZKNAdiXnLV2yeqRfDltqWpC0wS0RGum7qYvcneu7otg+NnyI
2JHbsNCXUoLUGms/lIiMlhoudImylsDn/+A6tvVcFIHVHF02Y/G+0auI8NVRP0hG
iiRuU5hBVYjkksPvAHDL4W2QTYM+3iDLkwvyU1bQIZeYfOaS316yyYk+5B7XTeh0
DoYe9k+G+obqMYwmSfIwSx6OZLAcDEBQ8iBpA5S++rVbgtk31bvF66U4WBQnR6fp
3cTvGjVNB39bUzciNpOJ+FmybiQMMrAklYiYey6eB+e4pZA8Ux6yhBeEbPYUJgyV
7J2rjv0gcMR+yrOhnRKzzX5CKVTT1kTML7lmWKdmuYvDviDS1SmhNWt0bWI9Joun
mGsuTpwptizS8Sh9k4M4+QhOlk4FbZOj2MiAgUj9tO/vdy2tjZtrjm9wzZxDgOcm
GLDv113VJedZUEgk4SLAWKOlb/IF3NIKTtxs5KMDRtkJjcuj50zpjO2eDbG9c16z
zhkm7J6bte+2TeVE3/HHIP3ox5pNIo8UUeh9y2LAkj/NHOGzVBaJvq02cNnMcArU
dUIVam4ugzj76HUi+2Q4rd06QJa2uuXcZOg+Za7eCniiAk52WewZ6Chw6Qf9gP+0
gKj6tbo9PK8tf1Hspf6zT2ocfNSdw/z+NJ2dZGpu67ocpmOvIZYj5ZLWrbjJnuE9
BPsV3vYJFh6SYrEBvf4AHy4pgsDYbtpFB+EhDK4DsUakxbh8j+lAtLIaJkSANr3n
liU7E5JJGSdGUwOz1rq8FfOe3jmVPlZSRZG9IRS17/aIiSWo9C7bNk/0kMEmMuJP
SwSydudecjJ8F93gzEvB26MrLnRViuTmnXxC+abRta/Aqe5ff0Tpwo/3T2x3RTqT
tOprttB9EUW2dR1XIoPkbJ63yvpwFtWOpmIYGDVAVhxBdrRuRStPCVRxmglywNRI
DxmrP0ogKaYQNtJeF1jcvXfFbqMiIEVdoutEbs1rgr9GBma1R1hZGoVM76n3lwT1
xYoEuN/AiyytDigBsoiQh6+8WhAyX/Utn5G6S9MceHepoI4BOKnguIXoepvs5Cly
NBqXLKrwtdevgI0s4YRq3Y9O7HYcp+DwOWTtMUCgndWX9WPW4eg3pmxX261cWjMf
QlBXiWIiCk6t/gLDHUQd+5DUHDf5F/saTCbQaDKAJ+sQoxO95CTT0dALbwlSdg8X
jVymnF7Z5eDCgY7r2lhsr1hSqPw37ws3AWxds/7kmtRFZoxTUTXapNZ6A1o5YWyJ
iM0h06meW2ir1UVqaDzX/ZoxCs9WwoQBDXpIMoFkI7oLCVBSFvRL+LGePYn7UAyY
Y85IzI+j2/CyI3AWhpB1ZZfs/Mx0hAREfxUHJVkkfmDA17lmk17J42vXDvmgyEjc
mThV81p1/sECcCcnfcbxNq/OwGvqfl4CJ81w0RMaj3iKUzXy3+exuJaZ98yyDCWf
oVtSzzwn9+Jsx7BGV7hjbnvRVgTN2PjA2c5Top23uQDJNDGHGSp/+uyOl5Js2wg/
IjwwFjbgdzowaMPTh/ajG11iBSdGUkOuobS9wHSg98kyNHT+mPMfzb7cof2zdSeZ
XFYMrWo7OTuIXzNWnWPXojsWcEtT+zDBvitZHgcHbX3Wj22jEkcKOKTcnDZnu5S+
lB9qPmm48xB1Qzo9OFCFSRlsvmKvy83eUy/IP7HU9SSlohuZJxhQpDVcLf5CqLrB
3igJ0ObDQRRlmPPqfqOVnvFjyiF6cn/zN9uMMAu5imK/Ry5Iw0cbvOMOoNoepXks
ntGQ6EbQY98dEfL4UtCiZ8rf4BFkgYNU6RhA2xCAWy8bUfIFe5BMk3tfgLn2GJot
TT3Ok6/Yx+HQt8063t89m1YbqT+baIsHwsHVasya+ENt2Owr3zPmoh2rZsUkfill
ZbirYgmyY7sJauQdVnQdvjW1Gz/espg35nOm9U6P9hz/9WcIeARt7bzRUPwsWKHP
O8t6mmeXLPr2aMgAVG05bPQbwFD2wO4l+cVypOrTva7T6cWbV9Fb27XPptBeiIRJ
DB26I1Okf2kAT3o+Pyfm4lsvzs9smxE8XrdM7P4eh+c72TwxG+H1FUhjyjRlPR6Z
V94VVu80rREw/uiDt00BaVEfOZpc2vg5+dnZh0QxB4DIp/po7NK/EpttVpVCrlJD
QEqQ/ZCwH5aaqCelMqqdCnuXHQryDXSrMiDri5uLLGjxAhO2apX1OmKyIThl4L91
ZMHIEE31NKawgaTl8gCQ4bI84PL4pGt0/KW8SAZM1D7AXhfCg5lixoKl4WztFOLm
dIFReFZpOegJ/4Dzu9bMwoEox0+a91nIN1nx9OUz9LUAFnSVcSmzkAJgmCuatBvv
wKxNVqIGApLR79T8vwvjfZU9uv/CJ+2H3ZwyPtqgXHOzXVqRNveKxzJtWYtPEal0
OuZCxD/Ru+uRkbTYGiSc9VBFV0e6fW5tXCo8o3xbUJM0tqs5PkDWihO9bvJhGtnU
ShmAsziSS4FVlaBeUrsNYVx1rSja7XPi/6YHDkrSxyLaKqbo33LOsJ5BZambpgSB
GzhRAO4Z53UPJM3N9Eof41t429jEBdS6jfUrRLsp0Zr84uU7zr79OrGY7P3i1hfU
5WaWJDaufY7U4KyMxcfQmDTd2cItdKOz5IOtvmOjhz1SUwhVRgFh5caP504TrOCv
dWciDqWXQo3xZ8fhYnF7CQ79yT60B0rRIHA3Hv2gsOLkCQAmgPrQ8rX+sbttnhkf
aXDhzlhfTnLSTK1+dBSr9pPBY8l4gJe9fo866H2S2vexNeeFvXUEk2MK3o9PPZUL
fhw0Lc87xmDSzkDHfQE46qEU02A1dDn8+Hxi1mdzEEoLj0rU8AlnQBaLufsA6khs
6FOigqx5TteKEbIGk/OlYssuWjAT8dt0MoFm2Wzgqvaan/tFpbwbtcrsvduCpc8r
4u3ZDEiq7JbZMqlNguuZ7d/0Qh9V+uUZOt3C9LST4hJ9uHuqXzr+kikDap6QHNuV
hBrkjs4GYsw1LMcpLXexlmhjkkunW9MuA+8WdnRsz4QypmvLA9iLS0sLX121GGBo
qJW9E5a1NNXfDBXiPuerMV/fAUG8oqqBuRINX/z8dQysP4XBRPbd/DulL6Kq+vNi
8ViC5Yixlway/HGdMtImSCL/+j/8zr/D7emj2fTYbM6eE5C4Cv1mIBJgaoXFPcYy
wjnyoSOBTUCA+jtMLLON/yFNn0/zwnytC6klTRU9sAcx2LMa9vrzJ+AR2msbiFLA
cfmrhLJWpMhUO/y/4Pt5c3eWnF18F/Vet5ZXNVGFrJYCQzRkPtQetB9aZ4bNyNfX
YzQo1nMyDnwaLQDnqioOEM7o/cZluyTea80NeDVhv6Cgil6FokuiHhgUqjGnSbp0
Rvuw1XckachpX/thJ3/arTUGNTnwUEC+NGOFhzGgWQZUynIsWWNkDXJjpalhACcv
e76DoVfcSXRpBQRWdPys8NfhxfypCriMOHd0dAJeu5jh9yIQrL8ksWm6Stx91iKy
oLzDxM+PTUvpduLBb/Wz5iOoUoYXZfuMLVL2YmsebpX38z0/7XbFErSpn6612rgc
VNPUdEYJYO6Akl10B9f66nOxAoSLi55ronuIOAsfB3BRPoz87HndaNoGhj2Ibwm+
qPFxXNFqNOnlorAOuGZcBZ4mntr9qlDrFbvptVKiWxvjpj2VqG3AuyrEtc+PeVcJ
64mdm/duFPUa/JeI0Z3IK+AQmYN7EcT2LqxVXe5RnBVObxKWu+DRpHJejoUOwZBn
cYPpvRUP9e/ZrTHDCVKjya4go3kvAY+RQ2AeowccPa+zAa4vxz+hh88Jt6djzIG6
A2xpJHj1EpEFlzh+yk8N5rk69i7coFFf7mvukLRUC6JgIxFaIhnFh8E2g6bgbDz3
oAIDJTonllPeM3xK9LrJvB+4PwFbellxtdEhYdMIwb2YNOkOa6OAkPR/HfnASvif
2L79og9ejmMIAMdUQukHmIz6P7xNfoQP/PQ7uHE7OrdjuIJF3iB4l1ap9SM2myRD
lPLjfl34bzds/Rh6qNIgsrB6J6+rpd7yu8lTO5boNpWw0qsEaRNKYuMr+8aAFnam
tUs4QdWPV5nDfl6deaody1HymtAXAznd4NHFoe2J2dzfnEGHQoy3ARYpTVyYbm8U
fiDEOasjiSNVeY+N2OCDC01QfcqBjrvIxtzsqpgnQzJfsyfBKHVxaIW4UVBGCp2O
8fPXZxGpGrdoLk9IwolGWTLWTQg2RB7L1dhANDiKsiabazBJqeN42uOamlRyypgw
3GHPHcd0n33kMfJfky+urxrRT3VFXmvEFQ5MYo0syMfSA4FfqciMSShLUHGPMp+0
H1iqkcJGW3C59Nl2MgJeqYg8JECHxvlU0fP8MT6e8/pvJ0NLvNM3kg6qUnexnfxX
DO6CjNAQORTc7TCnE8r/YAlXtV3t9+xqrNoDtBpl4TzTMstZ/BvgSCxHxY15NeWo
DLPlG19cx+6l/5H2gixR/yKMP9CIwYj5MbfoDRBKGkahAbpoqwdQ7OBT1wNhCNCo
6zBl+W7AAKdSDOyUhhT0eCkvjFsNKmHpfNbv8uYZn1RX4+AF/htgtKlqgzdLMb8q
0SrJYmmIFzy2FMfmfrfCmP7E5ob8qi6Hxva1AVPdYth0jTzihm4WbegPs5/fFUrP
DkSHJ3Zf1W1ATxULSuZz/zC6NsIf6EhwNNb5lGi8uZRicRvQ7kS2XpWhwe9cDU+T
xPr0RwW5dcmigTFdr1g2GCnJ/o2MIOVZwheS8VdZzgA5mubqJh9yaGiuuaLiyptD
PMLuK1SLa6oFgT/W22v/RLh26bUrmyrNP/cO3yGDorTbsaCjI/Lay2LXb3VDoMHE
KthafKA4JbYhUpBohKqcS8qTWC5XOcv2DoTgglQSdimEPhcy84nxo3frsmlijanN
nZdtRuZDHULCKOpx5CQ7xkOxmqoO4Ooz6YIH3tzb78diuIkFGBXiCoMikYTzdNNs
SyDdkgkzWVB/syV1eLlqLXnle+f++sSRa9EaMZIhPOJGLO8wTxRJSrm05bXa8yAG
ztuW+12eZc+Bx7cTK/gA9sI5IanT+LLkXUQoKc5bKJhtAwQaGZzyhzG8teTt/SRA
YU5FCq60CdnNptioG34tWU+XdFbbwkRXRUUTrkDZEOdC2IPAYePB12OQsn64JKON
Wkxi3pfJGFo0Bt3R32s0WNkzcvsxdLzomY/295Ak6wPlCTfgU2pcz4L+JrGFbmyX
N9E0lBo2Ps2ne+nxoyd5bb20tORPXSXBBjajXnxkzPOPkGTnptcgq4GcevP5vRNy
88CW55cKLqT43wVFAeUymxFp+jRU0wwov3T42HDK/rzolUrn/2BKOkbqavRrCwOB
1w0Bgn7NOyZXtfpY4xuZ0xLKos41gx4/OTPEKs0+HTQnd43VuoDWjGjKXAxGWDVS
PHAkvxmRMmXWS3cA7cqa9gm+qFU7HuVnxPSagaazrD5MDIJ776fkGwSq3X+DUGfn
3T20sy9E8Yhyx+hd6WjdErCLWQ3b+qM1goXgAEAxlxq+XCfVX8GZYV+Tl+XBciNz
nzGZFWn8SVqPtmshgM3wdIMPPVQtDAr3Ykp8TsC30Opr94jmuPwSNI8cdlAIa4FZ
mZFzedKzwbi+iFT1ucs4lNDErSazZ7kvOJ7LTW5iVE8w9oaGzGKY0nHSjMaVA/sj
O0FzH5PaBqKdBHO+Bqqnk4KsdgZcs8Y4+DRW2hfXkasfD7rExFuMidkBQcEyVEIa
tXzCXD7aBP7X6JIlgjMHCjqhTRcrEjpnhG3nY89xQmElhYv1cTG4PGvEhbafoEqo
9FcGvTIOq9Kqsrrp03lM1/XgIydcEVLJYIMTBTQVxMMnl7qW3Xaz2vM6CU6k7gEo
SsQAAYXgbFvGllOm20Pp2vJ0cSWagll6wK/DQYDrqvsxFAmDH5xsPVcgaNEQNCXD
4U+aZT2IrnW5WmEGM83YfLO0T6T23qz3+yJdtWW3sz+R9rZnXoIj0OHe0RutGl0b
GZtLj8M8nXrNFu+POC6socMP1yXFiXggHFUBY0ns0lIN2gcdzQMH+lqewQcZGnTq
ZudVbY9FRHHm6/Zos+hH7HFmAcCLUJjrzEKZhtaX8DCqHwZei/LeWDyIhsUBhmY7
72Sa3bwOoz2/W8miiHO+GYX1QQvhPDgRdJ4oOgBe4TniTTCyZIxDvzNVXLV3QASV
6/EKH93xfmQUaEEK8+4Q8u+1B/ZlhPFRuOefOskTsqF5p53xUPHAqaitER17dceb
4ht6UnX/b8YhCpKgrBdpuX6cbp+ETjGgmNFoKoxD3y5saoAdfOqPagqc2VB0tjIX
Mz3R6o3847BPvq44lIig8VK6qJvxkAgBzyGSZYu6T0AVxGHWw1MjvBDPehWzBldz
/TJmoFNuO0EA8NXOcZIyEwd3dRy+XD4Okv+Hi0JW5Ot/uhHNZwQDothqRNocxEmJ
q037y/z0Q+F78V/A5DlpVsyaYuk8FQXM+YArMbW4kTgKVoVUVoN1hMzNnDkqSCM8
4URVeziaP8BAtoayg4Nq0ql8sdJL7bq+tieDalcYVYJeamIL/Giw1eA59MyXo8Pf
2TraW2OTcmVnR5lLr5kB+4PfypcNTIz4HFTx389WHlhDbLMzBDrsRIkLF76wJfGo
y7UCgulVmicYlh36nFtzrEZ1eoPcqZq5nQIgR6MBnLBM3/2Vd3FyVMU8XQspBj/L
MN/PaYomfyQSUE3ek/aAg5L7E8gqqc3T5qWaht1dvSzCwD8XOm7+kyUG14hvbJum
l1UM0G1bz+JQGGlKzwsBBdJNKM+5nhPXCBJ6gRAbxv8+yG6y9UOK0f3HpNojteUU
M0g7oNP0QMCgsijAEAXmwGblXvdH5Hwpad1pXiJxq5GBm8MPF8y1Oeox5L5MFt5f
ir2ktE5fMPCUseKLHtg7wLz/NJ0eXOQabkxJDp5b9ubI/Hbhzq1pr+0KLJZyB3ar
FrO5AXFRvXTT3ixwZ3s1//d531FX3WL3OTru7UHoHm+QvJCDMSOgL1lNUwj/rjqJ
hl5hzRXfWnoDF+stnJ3KFMj45pSW9xQSou9fv5YjKmWgctT4wKLki3ZbVK7TRrCc
WnPjsuvJmBuiOnqT70To0kF2osY0nYDQxp2cTcjKMbnAlaplcEo434Gl40EyXut5
E5rpnu8EnGx0/9eHDp4pkUp9Q8XwfTSXTd0t9YRlBiSDTJYr8L2AvA+T3jxXN7tf
GOYrAHx6I9UYli/O/N4gkVW3rPACYheZoq+axeCsK/X2CtWvZ3SyI39fi5CDXr2e
2KV43x3hP96p27MtD3UcdZ99D9aEqRj9KX83eKYymSu9VknUlH/o5JIKSXd4i0oY
6l7pfKRhXb+pws52m0fP9dS1avHtdQBCDSGYJjGgcAem2hp1a1/SBFSDdGwhrp4b
lAIr6LbPxz3PjSBvy/LedqBdeXkxadyt4Rf4y2mNG2wOPtdceA518rU1vwTLV/t8
khjkaiWNbt1fqWtz4h4F+A4w4fE4VcXH5XumNJYhG3oDkXB0U7zvpp65Ue4sCiFL
RoDkmkgOe5IYQ+oNq44pZGet91CZjH16FrxvTrthVWeVO8YRb4ECn6SPoTUcKW9I
0JJQ5d5jZXsjE6CiyVvERFyrEDNycdWw0Ak7xMD+Bexy2bbZmO0hobfGPOJkSJ6f
wHvK7bhSMNXHhiell+hGW3aSesM963tI9/BeiG/OFnrrjfKH0xkv6SLZg64h5EFx
JcAtYxqSlGpz75fl0lzz6gLsY+ccc6hX0p7oYJUcEy1XABsoAgjLlOJkH84+BFPJ
aPUKeZ8viEwIqK0zeLcpX4mO6nM1kqbUm3cwi6pPvRzKRISKk3RibmsjpzJdjVLv
L3KvigePBwaTje+uAtM3duulF7IpZS/fR9B6ToRDpGShoSk9SLRNnDXJQGzLSGmc
2LrfgyUg2rmCcHCOMeIYL31/cvZGOHCr6GFwUNlcWt+35DJX8C3UoPJlAHWbiDFm
I3B1FHZzjpoY2T2QVwO6QEoC1pw7/cX5TPaYtH+KnrzR9zTamo3hw3cXXz2Amckm
kxOgwkmtsQ0wQ7p6moIS8MJQmXPqluKj97lMAl2JcDXNXgQoiKlS3QHOjE6qYbKC
IT5np17SI3QUCq2fVpHAw6mkipzsPXtJ4wIgMaT+PwU3k5WHUsPH/K/MfXZ1Zn+U
eMj5lfqx7Za5knpKyDLP12miYl47bqzRRjzLDf8uXe40ZXqz7+vstTGNZ07t4Q5o
FbvdVoGuKfa6i5Y6WwXCcfHV+VsccCLD0c6KimIBVLVsTJSCt7FhkH8i56FT3WWf
j6PbGh50WBN8Bc6aj/QMR366EFiQ/kWypIn95u1CI3ZHVrExfzhE9G0ric8N+IUN
Jf3yi3WleNIDMa53PJ6Q3Zoc+LcPQg2msOaed+j0kbD3bPabil65S0KtgyCTCXr+
2HKrlMLCVzJvzMNm0fn9JuhSur5ZLzEQDllWq9faXKsde5KtlFqZa/mZZXTW3SKA
QNfnDYxNRDRvX1uflj/dLwkBtLC018hRgzVaFye4Z0WbiaUWxjL6rl1nNeRd162p
P+51gV4CSz/TsMNfugW0TqhZ7YCj5lzOlXUQzLWFsCC6C03Mi/x0napnd2ty+dr7
78DO4P8dAIzkP9gLHSJnQZGNw7hNUMPYncCZGZCW+0TEno8Qfu6wGLrSeWIjziPg
13AOhMjgSiW9CHor0aR+EH+26Jd3BFXTzBvJPB/IHvmI17noKvbOER1Ym+A2w4Mx
ik0f0UOl33i9obFhvs4AZLcCJDLDEXkgOvi5YITd4WKROZ/VixD/RT1xbZ48YpYJ
e28LmqG089ya+BdTv/zCB7/dF+kKVIGNa2ynJEqqVPuAt1/L3jQdk0but2+JlGLc
VH+1mMu3VAEUeTFoGNwf0YktLo3/Td0c4OHzYBtPU8lODGaqg+ZNaE38rPnBNysu
SLM6J7geuVdFyv1GeQeGSQm0jr7luXoV77TxOTXj9TNgnc+dEhK8yr1KFXnCkgG2
/DVNNbo4jkYT4UOs3BV4wtjsD+E7+PCHAE3L6Fq5n4B9hh0zhYYwn7lhJ7t5OhCB
nVtpgmXWmuQ1JK6O1MBMp83nh2p9Xba6i9MWYXohcHrVJpK7hfQMgoMaYcb7zOdB
6pNJQD5Dm+28dS5vRM8VPWMpZOXZvDsAQ/YZUtxuvRCi506qBgwcmxpNmn27NgWx
TRoUhYc0JJY4MRmvuioXJRJHzpeL8uDzngm87qSMvG50BoMG2DaLOKyN9ipwCSz0
WIe9/jqWBGDdCsZrQIodvkCkgGTy3WaEZ2RrzYAw8dqxZsuQxKXs33r+qZOqOHSm
HLTBspkdSSEvldljNh02jJ+qXOsEHo/0qyWyIhiKj1hBNVrSV0yFsL6ZEXgTm6xY
khMmT+nk/TFgRbAYMLe+0iDHGiHChRxML/VPSNpO0ZVQsYAalqNUqJ+RID7zQvhE
7I9wLDvHkMsu2hqPtoZt8iuPfBeb6c6vNxKSZnIxO016JLwDYk5mGCgKmi0u3IQq
WnIC0/szDdf7Ozy7ykB9R3oewDXJYJSYqBSseh3IeBVmgWjjX4OEngXjqJ81NV9h
riHML9du1g+hPTxRRENHJ1RIlyzVSOhioUiBshX0i6DrqJCCMBBwpSSxePOr5PlU
t82QRKxvMCEqSPjQqPpuFlKt5fHjCE8dB/Oo1ld5vYlIUQkdO4Vq211PWkmDEqLy
MxaHBLkWPOc6KgMJtzXv+kAJ1bLltVJntT6myWmIFTWUcFXEnaE0JlOyf73AMN1k
V+yXZiQpU4FMTW3BQmJP8BxNj+VfydWREyIy24++OWyIya4ZzqWBJDTDxelvNAz0
zYpRkWpVCsWY3NZnou4gbiJuDkRMkDMFhqIphkOBpFp+L9jdrAKa+YMSgSYo1Yix
33j1YeYRSw3nUwlNxVk96G/Yk2VHnXJwf52vbpJpMokGpzyD0fSX2R4xQkZ0J0WU
MANUwj2DeGWQ8cKzzrDGEbc84N1zH75R9xgQcPNuDI3PjQU6vsjuR7EJVKjXQHID
1KKBw6lNMLSTjCFd4p1EjK8CyF0OiXqcoHbvsDbOGARndhuuhll1f8AolSPODI+S
hm/WpVB5c4iUqw6J36sl9D9mpazrDDPSEFoaPR9/ZWibTorJVCby8pc07XNy6+xb
oPhfdoItDB1aYB3SeCMlmoqPuOTgso/u1SYNvgRlVAWAaG/pYP451/eL0T9aNXvz
PGdjx6DI0+nC5c4uNx81TUrxrXVEnqBeP1vpJtGynFGUKkdY6KbdVDk4LibeAeCC
bKJ2snNHCTxiNOh5jpaz2H78P72CFL3ysd/E9FUWhxsvuyRA/mfMRGaFwlBOkdPp
ynWgqMpEv0qJLt6FDlQlBfu3RPnn2Z6q0IXX4fu8i9YBouaB0nxg1LuxzUDLEqsx
avsKo7j2mHbd1dhhEZwFxq08lm++jzwbA1HU6cY6WDqx9Nhh4F356rFVorg/X5OO
QOFc7WiXFDQSIejn9UCoZX436NX6KBpWvRD4S7ctWjFbBsbCYFYOzeZK0jjDib4C
nv7w0OgPH/dyAk7ipZ3BJWJL6mLh+gtC8taW7BF0uTcOlvtdxhJq46XT1jFKn8R9
cDfpEdWf3zSeJfrUpS1+RPFqp3wDS21MUH91bw/4BVOY4h8MjfYMWGYydP8H5tQE
hHCMLQdgwR8OGu6DXvVdj/ORRWiLiTKwRWEWL9w5tZtJeNm+w78GsLBlbh5gDORK
Nfds2Oiyxn7tmXk8dpdOlEIV1YdOq8QNox/XEQ2TiPZmL2C/39G058R8S7riYQQ4
Rz1VGOE6lCqAwq01TUzuDkY0h3qP97w/oMBKFIVC5hq+QXauP2mnXq9CODbDtKb7
fevYfbb583RPA+qEIMu4j8oktgqKcwjbQtZoYrwks0MmLVNIpMynnTS2YRIvuY+m
GlcSWdgJEIfnGs/pRYxa/g4+i5LzW5CdxzNhqHP437eYhIvwkXQ3gpT2+csgfRa2
ijkJtY7teJ7py3VQSesQIoBm8/T1IQBm6CDJSbeItxzhwPnh5CrtIsC1Zx4DKECX
XOAv5RJrWIfr5xbnhWQaQ8A2h0ERQgZ3eRTukWLiOBzXo/EDvV10/iQ06vRyL/l1
ZRwgVRqPIV8ZDMAeOfCCelRKZ0Z+pEI2+XE4YT5LLeLU8O2YPWlzAlCJK5Ftmlo3
NU718vQYYrzqCBE5pbX2aJ1OdBTRUOpNUgriVLKksYlpKuP3TtiNBCM9B3kr90Jj
QVnhFda1FO9CNHA+iMEsT/FPN2cQRPvIId7vKdNZU9/UvOuWz3yMv0sqqkKCE8sI
FqmSBDbk4AkF1MJBmFTJbC1sI3EsoLPVMF/psfjfPRM+NMskYep50iCj5w2Bo+p7
johEgn7sZXgsn+rL4nGhPjvaLuYXFiPFZTSFkSa4KSXvQk0sOoH+tivn+oglYuE2
2jDTFNIwvaI2BLZ/K1KAsh3+CqTzHLJg+RHntraWHYunxkDtjYHFllAX6taWxNGq
x6ewKZD5mPKqaF6s9hM9Xa+1kOnVogVB/b5tPoaWHKZBMJrkEjcehpxiv9mPVxJs
phBxHQ2/c0zAJrU/xVcCaRkOzrdFgfqCfM8i5Vn3spXTZSuy6x8JDvTgyK1BUM5M
ee2QhpED6nn5MQI/7CLUATw8XaBFJIzCTvm7C32YZ0u3lZTYM/ywunPj0hefWDce
hosjVvChf9lPM3VBiAWXiETm242hs45ethnwZt5Y/NO4+rXkBJCO+2I7wXsNbNou
4WUyOHpOzUc1pq3RxeiHQQNXthNg2Hgs4K9ovkFMR7g3QDKLRs1MoD4WieFq1DAg
/dNpWOrGysJE0p6sI3JGWI4EV/kzo2ChxusUzUJ4NjpZ0TaFytATNfmUfVlAMgrA
0ZMgEVzCCed6ji54DHBu7j8QGIrXLMLQQFtp9EGtEZO0xEzCNdTp2WnlG01LpehR
Dz1JdHskXFtrWvuIwTajMSe4yIHSpmG+B+J4FHyPtq3XbxJYhT1zhiqUohneAcxa
9egdcwcquwJ0JlmuAQBGXca62NMhUkrULYoIGJwpXCcUX1j4ciKPksxhOrXpF18R
cW+K41UrOy6i1LWTgXnPFyUOUqEFouIV2UMh03392zK/NCQfOdLHu22v/t0MfTXq
18hfoAPhhkqtNAjEACkaXAoaRqZGhzFLatf1ZAZsF4Z3eecmcRRnatHwRQ8sRufw
BcIK7G2zk46sSkCOW3niQGmPqAkqDb3XA+/zEWtBtEOEb9uL0DEH/Micmn8+avrG
OSrlTZQqWauoZ6DtkV74Kb2cExdxFh+N9V7ooiNeubOetLdbXm0kQGzJEhQJ2YuX
daQF/gW5DhY9FqeUIvGD2v081dloY9ch9fo7cwqI73eMbCa9jcCsTsuXWQSdCA4+
d7ihiSSeOfh+xVQ1+WNw09RCXKBi0pIGIoN1biI4rG4nmo+7AEi9y5/ASgqdzR+5
LE+tlTst3WGEmDCeaTYUr59VObY6kHFTZIf1Tqj4D9fee2zzy4NktuTdA7du5xEH
HOMd0LJzIvMYmnancQmTVkxzk50Rzy17NGS5JHzacoe6o9CwlZC+GpIPp7flTNK8
ZTngkHASoH7flrBX3457o8iPDaTzWxdRw+dCz0cJJerHXhpYE09Xvo/4nuBpj4Jg
Y//94xwjFc41KhX4W6Ri1DF4ksxUD9TLJ7srqeUK78p6OYqvwG/aWDwdh+1ubFYs
Ym4DmT+RrUbioRRaQgH/Y3dgcGCDd43qZdXKg9veKqGLBQBwLrYwX2uBj/MiyBGD
p4jnMi93LAEIa71DkXgSFyJiWrEHloioqRkWVHwPoGEraOYRfddMhl4bI0gWtvzD
7kiX2gImOaqVuGttDDYB7njZpWjfIGyyoj3O9/z07giNqkyHvJl7Od1/6ZuIls/H
W6P8rl5wP3JDSjPed8Sv2I+paifW6xtkrT6bFbjky64Oh1k2M9VOg2Om/vSm5gA7
8LBIbR3pangNDyYhykmRXhHpHoE7FgU/D/KoeP9DbMCYV0w0YPfSbRHjgZfF/URC
x4E/CZxxbZmiqc6toiQ3Icpl678a3FZykplVJLTt3O2oB8cTE9rWXMcmX4FYgBqZ
2k3zHu/w1F03dhKk+gKF/YgBqEvkVtPTZwMIHTUY4k3mB1y9T4pC8ChvixxkMHmj
Cs9Uo982FcPO0+Y1hiiUlOw4OEBmqe4D3r47ZNVtbX2dIhz8x1Xz4amRfaMvC3R0
mpp035wR0gLAYwrGq1NBR0s3+Mdprl8OHuzKEj53Sf4X2wf0qUPMiHItDWVeRGuS
/JpGrRelnyDSEtOLpQM699iGPxNY0PdErRbbVHuIU7hU0OJU+8+qmclIXIiCzW1I
/X2vYEUXCr6lLYCuKki8/IpNA2eiuRp4vl5d41IFg7m6aQYslqjfysRmDY+SaiJN
eUIyxR9Dlvm5dHJYKcBdoZlesmkHb383vwkLT22hPUr71sfS9GZaew5vr1QeV6wZ
Lg2Jal88T0x3JonXXQtwJaL+45yifTjxZxy3rN9Z3Esx9YvW3v3yZ5yEJn4idS3f
EJREIHHX8n2Jj6H7IZnZB4SRDepD7e/ZdtUG7RMHgGmy/u6khgjvINDPgkLy8UDS
YrNRDSwBv1G+Alm9qWX1CdcTfNpSHgsSbMfUi4JybSPz88PzP9plhGLrWDvLSSDV
nqSypvHZtXvCIlyUCvNSIyqObqG93UsZ3IcUOD2ala/7oS6yZNXd40Llf8HiB2Sx
GlktFvjnQWZjM2Y+OkQDYRDUD12tQmzJSJ1FB4UZOI0rcOtj3v8uRPVYPOtWuCGf
oZhuCU5BVcd3KRp3XcsK/hNcuXK1wSzlhVOQ3+GBII0tsbcZe4RJQ6MpQq3VLqmE
RSwLg+GyreKwMHrg+5ZAnNzLJM0rYtgOrtwEJtbxT0mxoxLFfgLnS0oosuGCpXVH
qDWJN3CTkCUwgI+Ytq8Bk9n1hPZdCViZ8SmL4fy9+onBPtP6JD+FoqMk3c2+JlZV
JbIr6gjtPK4vKTOEnksXNQ6LcXkAKDHquUpqCj/lKJgqNnf4J5K9UmBuYK3vSYNW
mZhcMh0olEQ6vF5IdqZXvW7TWYoUFSFICG4qOevyNlfYWggoGfupVfpWRJqcORqL
JFcJ9WooC/IsJpfY3N2HqvSNSq0w9WT3J7hYYzzVUmHq40Tk1rwqo2DODCdUUaN5
baCdpzlHCA0asb60qAm+m9IWSxxrB/BaIz18Yq22SP1xZFdZ8p/wb83qMkTHgrRz
q1QsPUX5KW4fxoyjTWGgmCRsuq19j9Lf2hBOEVIXMccmXJAGIyEe3v2j2+Pxd6pC
3jxfxZQvcWxj1viXHcM+RPSYRxadSbkFVU3FagTx3NTsbtMjiFId3vxEFvk2b8tH
wWwdtluWW0yysh5QIQDxoYzsXeyYQ2wQd8pYcj1DcHT8i8t/mIs6y65qNAJPyD+r
Yv24Lw0hP4ZXeYIeTHPj/8LE+TSonjc5Ql0dsugFqrzpVbN3jWf6EJe1FqQg29pg
dNPjqWQ7/mwqgCUesnmb+u4MelnhRrGO0lLyfNnzbkd4CWoDNxA74eMl6dZFe8OE
V+vTONjcE5kjQxLeDEtHZwp6hsNxSvDD9ZVEyPeIbijHb9jWhstAKObEsjvbXlFp
bbpBios7BgWN58SYyObBUYWvMWtZ0+X3ckw38KguIWzfGN4p0EKnCeP4nmrtUI57
EVeznDhXCyVtvbke/qrpXTUMbsLgj/5XEdL9k3OjpdwU+y/ts8G56cHPCoYkePeC
WtQX1FH53T+G/P2dHmo33romP6WohhrAiNvy4gB0BIAL3iEtpsjzbsDsk0Y+pUXW
GV11GJI6YhrpeNs/ygf8naQSYsJCtcwLSFRMmX5D0sqjeAL2SBJ/xD7YgcLiM5jn
Om0lkepnjmqUWMkqyUq5+FVgBixVgfHpO+DWQtaF4Bt2vrDqxrf9OQdFFAI454k7
xV+GW2FBLbBTY90DoE4QfmXtRBpRg//xklSfeFIiN/gQ8WQ2u1DxV7DUQdktlohd
3HPxgQvKpFz+r/pLv5ItzP8e1nX/Eo0YH2oQJPAk//NR1LYQOh9fIDWHUz6uDjQ2
lwoftTpIvdMc7wyJLkrTSsUYqGxc+e+5joj5UKoO7WAyHUi+bzoh3Yzc9ytk1Tf/
rErXayKqozUp7zlVqz0/TywgqDyM25GN6HTIT6kUfwmvzgssRP/WESPA+GBKkysk
mh2fHKSyfciUUVfjbLzNGrMRV+Xt/Ch/rGdm4rWFWYZdJVpoYEkDB0hpsQcwIHT2
UKSFbvCqUIjvfOEktj9d89QduKzok/RdWB1xtluxQokNEs5725Rfze9YMCrKIXeW
FKrspwAl8n60QuHQBDw7m5XtFFjj6JyM3rqwYB2Wgvo4OHRzzf88ir/3vtC1BGl/
pR3b58xgsAj8wyATePYEZDuVdPKHXS5UeryCRoMn/ySNdx5UTz4nA1FmNba12W2o
Kv26FNbekXUuAus7XqiA73DMmA8bezo9GzXza0bNdLcclki+jMDY0tbRgmH2s0ej
LufPUGs5hj/I4JalsjRL40ExJhm2Ip3z4wOPSLJ6Epxt9W4dsu7EEI0oabGTUon9
Bt4Ym/IWcElxjxCYopox37sHwqgghhb++lTGiUP1gWVIZ0Q3X66GmVuQRv3zmcpV
gx6c0NhIAEm5iGsA2/HbG1Y/JjbvvxnB9ozlA6qL7Bkyw8KXtGyv2cMSZiiPUQhF
lM2zMJdNjUuhQUXWJ2VoDjNLoowNaS00tGOiH1jvFkq5NpM8TkjHan6fqG9z6am7
9513N30cGcMn5+PY2EIhrAL+DMGwG8z1izX267s1VhLPmIFQbBAEDwICqMoopgks
LwchEE8s/MVkrUIJTtoicM3LXoCCyMXGNgZRD53tZhLVSOFIdhC1vrGf9dktqM0M
l5XTh/+1WdTEDCvZJJVv53jtLh5cFejpYqtiswn0gMH9rCMHhY+z6bgBPO57fT3p
gAbRnrd3uwPrinAQcIc8TAdBYJugjduVVxxsePYJQb3Ggt/hTgKMnPFHAAMkIk4W
4JgdEHd8o2Dnq/lHFG+b5OKKHdhJP/PoAfExCbgwlSrqB7kLAx63HhQ8BhrMTZOv
BwulEy/HhtGO4DKMWij14hDKx0Yr2oX+WgGXGwrEEtbKXQkFfGbF44m3+EkUeUh7
yMDHYjuVXN94g+ygUt8LaJQT5ZMjcTO+HRpanmWIFbXTCT3ypZb1Xwhjz0tISHR7
KQwtI3hp22wRsAVwCLRBqyDK9lCYEmNQBlLZyrSfF117qVAzTYLWxBFbhhHAYC0o
e+NE63EWgTygZgymCXAJfZY8xbHbxG0L5OMAiC7T0obACs2GZuF1/g7ryqtGPhTr
a1u8tQlPHrxa8eGHQh/vpDPi5Dn3t0HsC89H+9brOoLvx2TgIMOkOiS4zcq2YFj4
MoYeU18Lz6/PJzOIxocraGqfqZSVDydSlwSdO19TrCEyMfzOiH3OfybL5gT5Nazw
RLBFX4HEL1N6DQWkn0Saj8gXTIKjCfUNNXtYuXQKhbGI6loWoYacvZY+ONv+TzNe
R6waqvZidqCprLCJLn1yLu0GqYKxucFaWHEYxf0FQk7lZVTQMDE2Ho5Ie13zQpDo
ZoJ1bUQhZWVxwqK4j8aALLjl5Rup/9xyMy6KIGN8HQ7aV7ZcfXdDGNRkmSo0Mjuv
KfdnKdowMVVca5hgqwDjOElYSqEEn+U9O8xv2dRIFr2MZLfQjY5HOkVPlg7rzNG/
rYRy4sQFEHv5VpJojh4sgrFNRGvikfmvksdjHh1JLoAjd/qSyrGQ1Kxnt1PdZhBX
aGqwi46ddZ2m09FrAM4tBCK/tSL5wF8+liaD3YZJoaWrgunp+HmvLjrYhED4Y7yB
AajVKEWfyQGJgEIxoTs+fJixhHBe3QSh8TBj7AF5w11qpXAuXnYaHuukMq1wUTOK
jBi0xy9NDktb25UfoWAGnAPTaG4y8bpkjv7BesOcS6vpMUL3wSV9uc1hBvqnATaP
CzrPIy+RxU1S87eXMSUkJSVHtbkLTBAfL/O5L4Jqlh3zVkvITIn5s3+rmbPtjss2
KIJ1yNDlPyz8fXdW5WNds3QKDbbrjn8AyrZwjQxj3wH1scOUKvNX3Bo3EUV3jXmO
s2tluUcbfXVzAZdn2FoIvpiIusW+++WFiSnM9ttYNpxlPzDA1An185LHAmXt3i7t
3IAWvWBs1iYjpNUm7A21wm6U6+cH51VBguPfMFBDEkuIs4XIMrp/+JhHmPm7ypjR
9vEYNaHUvc2xdHAmuPogVD2dJ19pnUehOSqgj4LYdVtEK8wU7Z6EIYSpR41gIrTM
hyTSeMe62f4sf+tnf40p5W1Atew063BEWFvv/O7K0kaKLpK5Zng8U4CP0TpuO+l9
EUFEtWLIs5aD7m5WZ3zqMqCHmuVs4Oo3OaZGxfwLvekhTM2j1LAflntQVUdzRUoT
EQPlJU2uRtftv+7g3JubKs+SZWWff0wnYg4ewAwx8su0zlolFF70xWzRTdJDGTjr
Z8nIHkB13V212k+oOhujpBcmx834CEZ3bUnDTgD0cf0clrnDeHafaucOea/+JL2j
2soDeZEw8nYrqiE+jlTZweRR+BAupu733HEd42Dg9dNfY7fwwx4bQkTrpnK10bKX
mhWckCAX1u//iDcUXbRj1StkPPKf0veMgGfIohts5CypaM4L48bQTiZtxrejwum7
ckYAuVW2mWsg40k3GmzeeuaaJV+q51jYm1Fxj/++qZbTI40iL9c0eJOFCJem3Sr/
JT7Oua8qABZvM6OqjQzsOpD6F4/QinF8pOhzWg89QRTFeo27MTNQNawOFH9O15hV
QoSz0wGOok65+neKGpmYeUrFOvQJ66yMhX5FtX7tRUV9HKSWY4kbA4E+qoiJloqu
kLXtVRMyu5MRMzf/B4NudIjsVZJab7aA2MBYoba1PDGCruX1CnbMOizzMV6w2B+c
IgYPJd2qX/sJEVyC4aLMStT/fHnwIa+1aED2yCHfEYc=
`protect end_protected