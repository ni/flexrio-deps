`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 16560 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
FPPR7ws3fN+RQyk1V5tkgNSjTk9imAQuHSzH3ca8AdcU9ATJZsaaaeXcxX50PbhA
LUx5uRY34pSyAZ6mXaJxuhLOR7RQWDUm6RMvo5NrkQdsFX7DCKS5i4L8mvCPIxRx
NiD+3rvapJBFcqhuBxg647vhC8embN6fXse59sW3ITdEbSzo4Okxv/mBDba3netf
fMMxxbzQExj0atqLp/HJ3wORTgq/CoqxwDPrgbc87dcG8llfSTazY1PHh8mtHpE3
9UVpvgnwdnrhHnTyeh7CAfyNZPDEl92rFSREjEki6xdytYRm/HwXOw9PvsPAPkIw
z6STvhgV3cNrvcuTctcWSKP9tVfNlYj+8EF3GKbr0TTP5K5CfHLfMroM82gEljit
Y7EmBbmDGcpG6yeo3PFbkbvu+mMjb2t2M4MFJedeqIU9w+oAJ9XdfP/QcmFinsN+
W2Hcj9JvHTLA5spdXKW9UQm9+E9nmjK3no8AHv9jLvL66qVkqIpB8BIrpv270pJq
YWLyjj86DiBVd0e4RhOuhEBIYxga0EUcM6N7kIP2/PjTEtmp1h41bAbp/KhK865W
jMv7DfiTHfPNL+jcPKJNAH5CEOHKn6yBn1QZECkJ5C2+T79adVfJle82Gi1Jnzpc
uiKUb2kSPRo/FFHbkVIUSVdGpyzONw2yx/49XSmnA8g2CBufIlWgJRfOMhJvMpMn
a6C+bkYmxhBtdVHreAuO/RyUiav/omXUJgzW3S+0EHYQBACQC1NDD+lQeNie4pB2
o94TLrT9qoM0sEewF1bwlQH1XLCP2YbCnbIZWshzFYN2soLe0+fFn7Hy6FGMKWVh
Jo3Yjea1YZ/2eThtdw/k93hUzwPvkjuJCbuTkq9f9zWM7xerLIMsQ7biG2Xiskcr
QH/xXIiOA+3s/F0HRLRKfDtTavi7/piL2kklaYHcrI29PP++hG95m6A4sblUEQ5Q
TNj9IjM5cRU7Ll57TYdtmWWvEZH7UfxUIZuVBLSMX57m02WWBWkYmR/5o80hTbDb
JnHbeSllqdDW5JbR91DYsTzVzMVtA7BFH8Oi9nx132/CtUKqIM1PixPU75nhFFic
VjXePaKaVtWwSdxT9yxGzA8CLupkm+cPzVk6qhbipeb+kJWv/SkduUzdx8PhlhYe
ewyLKlvWt9brBTK+ge7oEEy7LO9rC9J8dNb0gF4pPdyQ6ViAsTKWdQdrDclEAwEO
oZrMQkuFAeg7pbUFHi74AWnWUjP7suncwNPi1whaBCcWXTyLJcVBM/3MH0w2y7CX
FteKE1flFyT6Csp6zfDRzyReCJfvfWkiYVDIdzK5D3WFWS/f9VDlVE2s76mcfKM2
uxWu1bhG/pBKRSrPB3j2jKgXaubPVJrpmOb678pVW7OIXfH1Jt9XADueWOcQHqC0
dzISjlgx0OO6gUPWH73IAzq3NaxeERAJlc9WyvDdnsAHD6ijKo/w+cbdb/SocFlk
uFhlEI3tlAp1bPESts5GJ/9IykJ1qpOi84wAnevtFl1XM3CQYWlr73qO+DOakk7m
F07M5yckNECDR8adu+cqmuXHBP0hANhCvDGmPZjhf00HUA3Dxfy5hXxwAt9XaEsc
MO9LyfyPA4mM2xwpyJbZoVGTI+7dpv8uJRzX3kUNsEUF/84Y1RP36JqRQOo6ULgL
viSjxiuWIgXMGLy/7SAjTS+o9KpFimvRzWlXLRFSEK0VLlW+PQUMcm+/ZYyypdjG
ZGD05SjjMaGA7BNRBaPqIRU6pxp6cpnt+2fnwjmWLxnd79VZxiH/Ug4KyLEFgUlP
tnUtKyneucsoVwf08jSyRb54KzT/vhC+rdKaW8x8iTXjqbru+P0CiGvti/x0vqIg
YQQsK39dOC6aDWnClzo+6flxkue7m8X2kJDOeFlT42zBo8edk45d2reQ2a0cBMAd
PsvuI2OnwnFxTdKri3eHA1sr9Awg1kXl7eKzSzpLh9CIuGtzhTvsz5SSdSeTsAlG
ynKkWPFDhXf8sS1jXjWLF7yRbzgUm/cOWqLKrbjDh1I/10R0FCawBo6GrxQ0Ew6X
U/3d65ZZxfiWlalmdpMNhrpdHq0quz0cxn72zTPAyq8No62o7/sXF0XmxdGzhL5m
C7Qv8y7pPRBrwAP2dd9QW3DJDvu2yzfLn4h6rgonKfJ2/UzGVki/FySXFeEEsuiO
eRU0B4crjylhOESRAtgw1zw5V/uG/nj+WgNvwvN/IW2GaekF/9iIXi7yLWB3b3NF
lh/Tyc7AIz9hdDnhoTzrJ3NLSpsQ2PF1OAc3DH8I7sBbTiUQpFbH6q1TcBZY8Xuo
kbF0VYAl83LLKi2gQswq82oJv6qAHrUWmKli6VFKuMp5Ka3Czgc1r56FeyX8fdjq
6psDQ2w4ep+T0WvW0iy5udbPbJ5w61/BrWUlVV5/84Doo+7qJk3tjv++efZCau0x
LfqIX1Qwm5UlxCeVpnGZ0AHVyQB+eG3mFbypUYGiJ+ojXLbcIEju1LOK0I1UN8L9
ekkySk0uMSOUCBxdxj+6C+IsGQ0DXslPNd+dUNEDhlzp1Bkle9drMS/qMKmNb37O
64J+Kt+vWCnLFfP5s9zA8J+lDQmm+oS+HRXLDAzu5Bg5twmO2NOJdKhSCGXrk4zf
LyUBtrquFJif36t+a6g2pwvgs8e4yE2UjlgM7v6m3ahNwgB5s8hSZQuUyj9pmF+y
HE+ffFH1L6noLCdairnvXkuTt61G8a+7pYpx++5/PchL11XRjh3MmEzLpoHrw51u
QCnUnRab/6E2jrz78JDO99GvwW6tenl+Hf2xFU8TwEIARC2GyuS0HYS9lvdWZnkW
RCXYMTLlR3unUamM8JrZAhSB+NtT9znw3oyLa+xRCv8GmXUsZM7D04LGrKCBdzn1
sBG6d4KvRCiNVwB8GTRfRy+9ZxY90YxedPeicPTJbfWuaC9MYCcMYis+NAJDcsqv
OvLjrZcT58jS866Et87KFGodaGaYesiWCYAaPBVMEmeMgL9eMX5svgt9T28ttibZ
V+nfSMBdv4tGvflDDk1VYBzk9wXsB2duwiGk5ZfwUuyWyX+rA7gKFr6wrqsoC9jc
Kw1VqdDDHPuTJE3vaZv2l1yDYTdaXBncl2vaKKrjGSmw/WeExkNa9L1DJ5JSJXw3
Tja9JUfC+DGxbvSRSJmY7pV3JKu1OtZdaoD9FKLOOTWRK01zsXCdo538znh6od76
CkkmWpUJAtHfWEAz+Lcv8G8UHW3bUxv3bK7mT0BCNVaS5iRF++g2hYeRs2leKfrd
Z/RtMKPX2uzL2x4Yu7OIj2rnqMvgQolUdDlke/Q80V87id2A9XJLbWJC7bhuQdSn
ozfZ7fsm9kKHW2BV3N88y4wWngxjgT1Hxot61BsqpUxVuTDoulyS9/BCABKP61ft
uuPQ6/IxBR1ICc+omUCoizTLl3uW4ES6yokrN6Wca+DUYBBYH7xP+EP6w8MtZpg4
Dger7owMnDS/+lD3xWMOtnQX49I/cCgz//p5WlEcepZkaZY8AzYaVly3O031LF2S
9VzIRsDJhWMJSCgQYdcMoDYg+vZbGonMYyqMzVfjsQkKD5yPI6fc+FDdxf0VrxVS
ug+Q22h1TjaMzlLfO1+UnN0F1oK2dr885kR8kjBuWDU+92uuqs73s8oqrk1MwgCU
OEKXDY+t0t5Tqv5gqtPGYGpjZx2BJS/2vmvuciD01zJdq9dSyc2r87DxEoc+3r6F
rJ21ITBBYKy94alVUeIMPSxFQaxjnHfVsKpk0CwvoFlQVoxOsYzbwW5mBmvQwTIj
Q9P2tRyzqKFOGj7PbBQ8CJ0vUttSVHxo8Mx0Ys8VAgP/7OluBJemlpfHkL7ORkwp
pCCaUcGn/2RsnxZgI31U8O//HM2RNsQk/vK1aWqxPKFMJ+Tt2h8ifoYvVGre2XIS
GzO4gYOApK5dIlq+bhfq2Yq+mew1xxkKPAR3DPO0/ibiEJaYRCLyhrd6oe4LrPEt
nwnJLRv9lQzwzfBLgQkabbwOGNbJWfgx91xKT/MFW6dqEtrwhFiycvvx+tssjhCE
oyEUH2X3kdZ03NUocW6x+F+3KKUVXPyRVH9YF1yR/D8b4cbv1pOn0CO8an8iwaVe
EazL47LVqAcOjZSrm2yS0v82MvYLUmpNWDSuFNIyuWg7dHsl/yyNAvZghwIKceLa
yzt/KTSQ6wc2hPUjIQG4KMePFHgpb6uMUXHHV3zd0TeQVOuFO36VnVLNnfmtAGOX
HV9fc9H1SEngeJ3IGBiPn/byGyaS6KKLawDeV3uBwCttKfU1SsN/WektS8luXK9U
H8EgLR5i0FfsBbIzi0lSayFadnULDPbTqcsCyyURtXjlHPwPeX0eF+/p1kLBlLkw
ENODyMCTfemGe65wHeY9LP5URGQzusQpYO6X3+R0axGsC0hX3fX/+zDL4cRY+txr
ZOLD0mLqECohACNl85yDTTSd411uHxDkpj/Wsf8OidNGr8qXjXIPOcNif4SAkV4c
hugNW8TWB63uNlbOc9yHu3M/eMA+d2Zzh3bdC7y0S3rTrXPppJZoobTovhDV3dH+
tJz7Cn8JjBzYCBX/ht/MpgOHdLaYT9byY1svIB88sbKrqYCGffJKgmsUwirhS1+A
ac2ErcU7+H9vGiIi9s5srE6CpI66fih+9PO0NN84be8PkAQCMm5vYa0u47oyBavV
qhePEoGr9aC9WhLw/q1S52GSyk8z+JVftTM73mI2GQUEWyG8tQ5zUjkJGkebhQiC
9xWonXuCC0J7ZQxrbYFmJwDmqiOJ+2rOhznPzJhsx4J4LaDnSMQ69zaKECjXnJr4
Scu4O6KaNZdIzfjnqAvBaaL6mxM46PvvzYEpdTCdmVDGto+T+tIxVoapJR76UH/e
TkVXkt2QoShWtC7UEL/ZTVrmHuoyfw6NxbLbvGeh90Ob3TrWhwWATQ6t0Nd89/bA
G2W8GglyxwWjhja4dqh+hY88xlrrHJUy/+k1/w2RkqSNVWb0Zw5Q9g3SIESKcdky
s1e8MaT4VHEab/kJsjMZDNeJutbpgxVW2KgxN7Hle0xebXa58FHU3uSDFZ8nxbDJ
NziAPDaEi2LUbDdxxoWLdC2ZPtf11lGAWEfz0lNVTod5FWgaW3/HZBbSNAMjypJU
a98X5lWL5R3Eki/D/HUmqHZsq3lIf2E+mu+Mc6bymeDxZ2svObz7n8qRRTW+hrKV
4UzMgQOkFs2hpQ0eWI6ZN2ZlgHtG02OfxnRDuBdQ2gHri0wXZJg3s4shc1X5yvxR
QTrcgEN8iSWOGQxy0vslr95RjGjPXV6PG0kUJL0mSqszSUGn97evXfMVsDoMboZ6
AkaiFz68KlNLmD6oUs1O6hNR2+GoIqK3eh1niVpaf5TGQ9Wv/SJM6lD2AaOl8r8d
t7eAT2EnAGQE6HdSh29WrsIybUKA4ltC+J9IdFUltrkURnai4NYjXdFnBfnXO9pq
PfBh9S6vNZn42PqBUzcGxt84EFbgqn69xASi1yrQHtb4ZOngsdpDW9cfP//gMG7t
WVKuwA7xlz+vOnNjLvYinbm4P9mr7vnoGQcGWtLQd7tVJ5Qau5qBI6UW8wFZp0YS
+WvE2uJbejOr6FJoubT7Q6GOFekvfSS/F995dntpPKIJNHG/JNN/9s426qhJFHpt
tEOM+PNzyHqjc2U5FgOEuPnBp7GTRK9KWneo3YUrkEyaJ6uve+7nz2J/IiLIW5ji
MwyDvn2IcZGfzQOw3TGMMiS2y3isylQRQEhJa1LdToISew143JXhenjBP0QjDO9H
0prd21S4RJL7yMXfD5aLY3lQAyQxKh35Zsq0E5pmUIf5VhmeP7AZaBt+C1aTNH3M
57n5VjinOolCUYHoYfWfwrn/c50ISPR/YKlm+hTq4BCoUGaYRbJD0yLNZyYqt3OI
MydcS9jfJYLEJ/jl3f01l3IzSovIuL3MZL9LTMEwAvFo/MbtvT9y1k+mCHN85ZFJ
2Ooo360RkBhWYAFNPfXIV3bnsD2KA9s0kE+Wg9UENDVrs69EHDcqSSXDxFM8M+Hv
MLqbhy5e/vq5mbvJWKLOfsTu/qp/1Mmdcru0dsz16k9+ydrow0jzALX7m4N7TTs4
kEqIYV3xahrdI6uSfI0NGKftBgukAxTIjwx7OjN0aKvq3lEjM2x87sQ+YjVhAt5B
1K8sftyu2NQOSVFgqp3V/Xpg4vGZ212XSvK2qMYZJD7WzX6RjrtWPYMqATAMkDuq
LE8LCaOgizGeu+1LBqVYBTnR+wat6ZMRSsI0ylGFn/vmLt/EAGWUcZAZOfm1wf1V
ri4xu6/dLJChEtp+K0hSrgaxV5LUQv+R7E7+7PVM3c1Ds280+gp2940nKnu2PcAP
X8/9kWxrZlff8qC4v3M/59lTpxQJZHYveJMYsCCOPvl2Pw3WdCRw5P3Slq0y99AH
tLzpmb+AM7ejWk62TsjC1AenegC6aKrljvSL+SWLAu2UfsU0SpOsWqBavPF+sCit
FWPf+MkBP07vPHla5tUaBYsz6oNEzGFpgoJE0CRJqM/pLZVDdf/e8MzsG766m6zL
cjdkUabXSRPPlLbutfl9RhE3i432YWP1Ae8ZV5HTo5aVfI9fH2uRJa/2s6UZkoGk
XFAzMd0bqnx74400R++ZlTUNf/jx8k7aIafBttZsYKny7Mxf4XYEnroyQHbLA21y
fNJ5CkP2hLU0n9yFmjcnwTRB5Kee9HBQhyIjOnwM0tnk60YDhdvtGX3bALZNnlFJ
th1ke4Zyt0FeWgGiBdOejyJaUXN6jRO7gb1DQ/WPx46V5ezDXZkwvc2Ac9Bf2pnJ
P9vHECbhxUez+yKmUK7JwY3KoQDz9GLFWQsEuGom/IDKhAbPXrZgrji6Gk4c/x2+
jI5tagjKmR9nwB3BejgIcruyPQFxhhN+58KREDv8PQ7Ev8A7ksLR3h68NLXACzVP
Tk5G41NKdaxUJMbfV88Hqrhi1PqiUGXyOoGhYdmWitlxdEyezyOaixl7LrEY7ZuM
ErVtfpvSEI9HiPtUyu0FdBJXiNcdNMcb52/zt6MX0SEccafCPrBPu8fm1OAHw9Qe
TC/z3tXGA+8gwsnDmJnndP8pMMZN5TJt+eVp1wt82S2xEQfbQ3u0hwk2kZluDrIW
R8AwcdEafK8LY8MLf81epnGxn4B6bFbpz1Bn/rLza1eezGEaX3rTWBzhGEa5CyhE
wMs1fyGR7UEej1EflfcxcCM2/S8FFugt/WJPfiIiL3L1WyQyJmmUiN4b+Icr3mea
ZWa7ZVfRQkMTBUu3gJOYIAHmg6x0wNt1hgx1SGjf2LUV0Jgn2rYMZfSz6Q4/30bX
e3l6XeqoaJEYmc12hghNc7cbyiaPq8oHcW6X/mT1wymWwjCWRjkt5SFk5/JZ7xSL
ho2rXOyEkhnfSL9TL58Q2nXyz4Gf3/tj7bKGNRFZddQ/khKiLhVsRSawJ2bwCVU0
2R74VBGQM1a1i1WzNykUO3OlAsUkvAg7Hwz53FaFJ9dPUN6QyB9i4UGfSfeympK/
YkHIJXO+7FMyUifhTMYqN0Zwqv4s0If553EAjUn9TiXyepEhu0ZG3PPeTQCrUHjB
39he1+96IWjEmFbmFeeAqLZB9TcTK3Ac/JYsuawiPe3Ez4BsdPWuSXt+1Ltz1v6E
QKOHdi07HM4HLqxCRg4DlF/sHWbmB2OsRkrHIuErf9e4quwVRWDtUcRBtUNnzhFJ
pVUeVG8xJZ2KKqSAB9do+d8c0HatvT1AfvZLiGNCmU0BOMitBBtGuA1QtGczpQ+x
Zw5gOskHq+RbjI7BgFY/o0UEcCRKr5ZDY5Cn1KAWgTXNApbJ/Ji4n002QuPu97F6
AhsFslinJq/Y7nTr8FypEkOfGTWj405t2/+hiQnUdbgctwR/R4I5rYko2/roFdIV
osViZ8olqnMUznB8Rh2OVNUtkYIMoZ8I5jXrpWy5X3B44uAueYJX+VaR4YgLgDe6
h27wUj+rMmud5vU5+/6TEO6AcEEQYcI5hVrTTym71EAXS3B8gXx8935DNpkMKIbc
bIuI9V7JLAAFkyIEcBlrku3N98ek9ub4AW1aHk2hBgxjzqaGfnFt3k8FyiqqFqNN
VJtJfmp0ztCiPXe4uGKBI3hH4klSDHewn3C6pfqAKQ6ggwdJrtfOEylDw7a0+/7e
piY2R5oj3rW1ROPK/xEScbGv2QeyYHz4VjKs02lyZdIhwxzs8ZcutG6WSz3SaiyU
38gLFORl1McfFpnGUtBnAKnCoHLii6LN0VwldWFpXyWysnTNLxv2Rx1U7pvqdQDq
xzUzMEBjU4GuCQdx0vhGvbPAYIOHiMM1X18t1+XBkyJ5yUP9zXTFfqqFezu9QhIn
PZyKHYS11ELPU4eIRK+AJxWHcqcSnwRc2xRtAOVjEbz8vhRnyhZAeguVWP5VBhL/
Q6GB6hX6KB9vmsMQSoqIuy/I/tl8dlG4NUEJw79RuAjDXVQPMDWCLReOhV1kKoaB
lj/nVfTPqIzESO5e/chfOPSpFHXLd8oxAy5w88CC1ePPPJh8rnHUbmuXWdpQZlhd
OIQFMuukacQWZ38rmLIkJSnAHmsVfpHu123jA9XZw+Jxtk0xuxzBBK/B627ag88T
SDQkrfkxJpIdRRXwfX7HP+biI00/HhjtZgkETlE//cbHfOBPu4geca9NDAPuRRrw
N69pjSK+rSCrBmWmtD6ol+OO0LTg3olldNNpOPA8ItW3jS7CRWaNP5Yag0IE4xqD
tWGkvmZLaMoVrKIKCHTdiWrCt6LFr1VFOkTsilKzAyaqZFogECzbOF4rTwbYL+Kq
rOw3jL0NsAJEaIgEW6gwhvIVjYsEoN3BAewLLgCKI0HuwnJHKQB3GJ6/FBoGdteN
LtTqX07BOP9AApZmKZOg0dVqGC8l3WNMEj3iV+xgLZeO5QArDV7qCJuL0JpVdSwX
FUK0PgIepcm+lS/QoeFbBHvk4cZd6n/gVlflLU8P7UUaOYm+uSNybt1lbrkvJkD6
iNpbSzTAM36QHCnlHGvVUirh8yt01tIRPvZJ262ZsuwXC1L9fobUdAcbM8NcGGui
/qihOnXzde6joTYVbm2DxB4z1xIHZeMFYhjn7l01ORxwNGknrIhyYmGIMflaQKDI
P4/kydmh8gxy0KL7HLcERHrMq5XOWotF01cZnyfjDX3xzveQH4QWS6fibtGbRcX0
5K/TJnhkw76g73jbEmolMficy4ZRpOd1e7E2q+9TSQ/7keQDI7e4SlUj23/l8cuN
Qbm5XAjH/OAqC4ogTVMCTIOQIshiWJWVruWcYSWDSWtG7aQUvNz7FnkaUA6ueuCT
tdCBykwHCVeHw+ZQF7dE9lpj+H5XryCqc5NfP+AGH31MNFzVhbuieY1wB3k1V2Nw
CzeRtRlyfvFMTKuHqhj4hj3PuohRM70qfd6cctgA1nunqLhCaL1qds/VsuKMRg/e
87maCEbd6LDe9mpdlQARcwsDPTj2koyZhdT4woYjw9faraet9jFWiWwGsLY3CjS8
/p2urGxGZ5TUaz1Ly56b++u3BkgUZ5GAVnAVYXBLs+K54C3SZeBUWqsbC3FUAoM0
ohZNbSUUks0mPvkxWtB8CBoGoAKjgoYQukr5UEpkFgJ67x2J08wb91ajsidMpzLb
8QvKzcWcrSPHsF9on2xAk4+TsLc76oU5MrpLxiXMGFEPHzlmNJdq4wrwL7SySpfw
KMHySZl96tS5LqPHiNTXflV+ZRD8N6mgrMjATuQxcb+bo9hnNRFF/l3bzrRV3wsH
kisz/ln0LR0u3d8Jm3dkunZKykfvDAWTfgXC/1Fi+axlG5ywmSxshVHe5kMrqnx0
yC6ixHv2s+mDMPYx68QC+USh67gUjeSaD8rQnVe5bOmGdIVR+J0u1CZE0ngg4OV9
lfZ+XFYvGApwpccnTJVassQkOhAbAIRJ6XubcjLHqVhRwB6s4S303r6elAZ8go0t
sRIyC69Pd5ztq6+CFq38mASIVbUX8BlmcR9za8J3f7r2gBcwuvAwrhsJO6ks9vxS
jgU2byR52qYQ5giyj5n0TTUXt1YfhwS2LJ6HDqbB+yr3MvZcNa6dvqO5Hjzp6Hoe
jXghEe4UIaI3/twxtlFCaJNze59C+XQq8qMIHCVG9tPf4Avo4SEp1KnuAEDfS/nF
24Jh3+aVguaKEA5B8fbY0XYmKvMMi53vVDPezxgrViJU+3vN3gfrp5YDZvQMxUMi
WrXWRzbg0FR2oAxwFRRDSXw7LWbuOV/+tPqhn8w2sAs2nTsZYfFGP8fB/2ba4foq
l7uLGNgNmzS7jsVu7i378pgaNI5RfPBKRhE4tuZOzB/5VD/EVW0SemFr5AkCXSZZ
iUNtWV6bgrhoiYVPoZZzDADH2c1uzTmh5jp5JF+O2e+f8LXlyoetcRRDXglJfyA4
JqPvDPz8DdVrbGNtTvvhrJBkttgxRtSjV3ZByw5tyF6/6fQw9vrzjfaEQcVtgiED
JepVewyUiqNu6FR5KWfL5Zll8w4uzRglcaE8SCOWJfX2o11dyCxMToW9tF/9eeHT
kYWQ0geM+oD8yg4GHDaVST7liQAo1n+CkSQz9JXg9hK+vuMeqB5dhnpRWCST9tO0
Z6D/TsrWWLNAH1GlX5EUNVMdObM153cnmRhsfDrfoWuhwhgQvXkQHpoMqGScXrpk
KZQB4JcS/1L1Pw6DEFPAceW9jdqTxCZO92Zzgm8iGJSEEEGXZTZ187bx5ybkJS+M
zfm7DcWmsaaXqk7gYteoew/LyHlBdjaToiPw2G7VFqkeL9DAlsvhKVTKjGz40RrW
eA3TlE+erJy1j466AF4yQ+nN+edYSp6371FI8V/ZrPpSpUwrlObl81XZgbSwP3KV
KxLD7X08ZHNvFJQxIp+X6QxVCqn+lvLYjZiGl53AA1+1ZCskCTUAmRqR0KOhJ+e9
tjRirYWliePzFR/l8aCohN3CxZ8F90COp2TCh9OXr4L54qp8peI44ISaHKIaiEA/
57TGkXj2lu/fs/934GuSSGOSjGsJge0f6ZHscO6bRtYQgZDLVK0uKsB2lA8cmq18
1cwMJU5OnaHjU6V5h1D+4K2aDZH42YCpJXXdzUuwIcjN7yo0vTd0aG5thSuGwaq8
CDM53txyNJDXHX1aLW6e5T+3qqqc3jR0xHFOnvuaOHbDDeiMEPpBP0cbfTzjA/2i
IhA1BruY/q3A6Z8MQRjqdp0WY7mKnq26EnIiBkOOJbVuMC9J9Z3D4LASIs9wytTu
0aWMDoxnZb1mXAoR5ZKhKy8kMMbdNzV5HoCqKKF/zxUGVKqp1YpiVjcrzD4KxSUb
W6SzDM8vOq4c/VtWjjQcMcQb4HBweI8qpr+h84/V323iRiMP0EAZYuwwJ9iL/dip
ld4jwRTXnzdcjEL7PHKnb47HWOZd4cJqyXAYgQ9CSsjpUxVe+ZGS/NEKSnugTta4
4xggaczUPAlsl9e8GQxWOfMGoc6S7hCd1w8pDTbj1KgJZXaGu3R9LnADxPHOJ0Dq
SaheiT69U39S6ukTYur42HtWHP1odl6jx3z6HcRYUg5NryKvdrBCBC6CSxTn2PMU
4ZsnrMvZzcBSnFLY+7glN1ipOrqvYiwXKs5C+2MnJUrtEWa8KhcjnV+tEsYyrFqG
N78JNaIX/oOELwv7/aM4F4P+TPcyQKcMRta4p/WpRyGAUIFDdJQrQPC3FSnjbvF8
aISIoaRoqLpuPT5SLLrNwjYS2iDEQMFSEu+/vE5Las/9drB7Gz/ihcaif7KiHDRe
Jzr1WWbTbpnDLbUhgaCJj/Ub6JlmQFji9mPRYSth0BU50ezj9ioZos7lipfcPFNp
TLNsrrc09W95gRC5KmjZOgNNAdGrgLVCis8P2oiBw8lXKZyRB5TO0mPR9+zMyOeQ
pjsZPnjHVzsiaZdK3V/tYq8bbOX+HdB+JJ/W3WhQnE/GXfU636kLxKT66CT9xPbK
IpTcGaDwG7BoTxE9hWdesgFbYoVUQ62qsGpu8YjbndbWN83G1JiLMa7DSQQ5fyit
LEVO6QwGDp1fEdimE/Pdh40MM9iWktqKqTYAL4Xnl3okmrSJacfle4euAw8/Z4eu
tCtwKxGaEzq0I8Y1EVpSTDGCkF4s71tdIZL7z11QnEEqRpUL2/oYz5m3hUOcOh9s
B/w5BSB32fYrOzMarVS+9Q5te/ZONkE/dfEwlgFNNs1aZz76EyskXLDAPNxKTBDp
RFTlHK1EnNsy2jjk8JOujEkxeZhPbzUhUTfimeG2hIZXJq60l20EBlTg2BrvSnXS
xUj5IL/leQPxeMxsNS8p/Mb++Ot4OTyEePuUIpSYKmTolZFBrA4xF0/ASfjq3oTn
wZ+MdW0JdkDU+IDIgfxysXrJhHpt3LORC7A2IHbpzzL9uVUIqTiqelhe0vj4Ifhe
yCBRKdw0qz3JxYT0jaK4MVN937LB3D62C6E133VfbLmgkb6Setfg721/1KGt0M4a
CNslSbiSixJO3f7Xv4agq5COaujuWd4HSi1J0VYplRcS4KyAuhCfo4CihLwAa6/4
8V/UAZHjhNnkmYY918Z5IRTZtPrG3pTkbiasz2H8f8SvbL/O02AJ8SvuSyC4AJYr
s2O5AM0pAW/YQ7d3xn0Krtj+LCfe/A1FYFWi/FF0MBzsfJqQBji18MgSva7sv2lj
FA2Bw6pBY2bWGrLJDyHwMCUdhcxj0U1zxBhgIlM86SPnf8rvvXI5LKR52ExRDg1h
ZyVnGPuOvqNZyeSoh17x+jfjKgLsYSW+nJQdjlikY/YL0SkX6InJ3zomq4NavtLJ
Vr3rkQvugbvRByJppPWfPlXlp7GGaUxcix9hR5vfnJjOwnuEvHnS/Aq5O3ypecDe
3qoRGvyfBxfZ+zyj8HBNOYwqJVTFmTtdts8i5csDNybNhiBxmHBlT/JZpVJyx+mI
V0JmXbG555T9z1gPii75P7gZpJb+NY7pD3omQEky2+4tduGBGP6pfapwx9eYZVjK
15wyq0Tml4QOaHZYSjrlD05HOX1sVt2B3SiH1BMgVBMVmH3fr5Dp+tlUIPWyJdiM
JXwAccRPHNhQDUOCtWjJiLTF/XXxy5WHqAsVNXJyB5Imr8G/+KDRd9YKSk4UmfvG
o/hTiJAPfTWdkByRvbLLKATxkkUBA1w0/wc/+VgiJFH+pVaVkeFVTzWj6dR1rQDQ
xCijlGR3QYdemVRnMN4u661YQhDYjzCU/AqFihtdhVGFJOzW4u4LUL2s0/ZrxYjy
qRaagDX3UR1iUPQ/nn/SYhpb4PVlgCkn9GxdfyfaKSlrhyD17fH9rneHZUOwgg8C
y/kwSTUg/Dggm38vnw/xnx+T4qwzzN9cbzlpABmIp0R6C7f+f5+QImiHrIV4PaRy
R8JqY34gv0bIJO1NKBFwGWPU7458kZfEF10jLDmyuOh8W4hywd/O3tfCe+9xLS7M
8qQIwmxfXonhYDYfSG8FNetXSBgJMsa9F7R52kKWNkHqK0dCCGN3gWr4p4rYsS/L
qwlMAb5JeUCV3NUIezU3XDWshpYPlAEgDLa2ttjR4u4P6rdbr+l3wOImQ9opumem
YY9EtELCThz/egyFbMecFrNKHeobhLZdEjDvIVJXgfCZVi3rUINak3bD73bIUhmt
WO7P3dVL0whMRVoOPpgRz+IV3rh06W5kZEVtQyzUZnylNifcd5Ff9v/PIzwWfig8
MyBn6S6ztrG7DD5HiJBIcJRdv1bzLkBzM0G2WUs278/mg11Jexm13It5QAppMudW
QTRQZbKnbPHcFICsLhG+oVyrniz7ck0JwTk3b0YbxLC52cVeMy0L0kfGkxbiBmp8
x2F9D45yFsDp/3BRt3mpq1iB/4aqJFbegfumaQxqv35gm/NHGdvVycYoG31hcdQb
rLhJ43G3d0pMPxp39YnyjzsxC2nHJo6iv7KfkmjJtDIqxyedQ5vxGZzCwPFJwNbM
RRUbQJXE7Lqo6GJdT8M8I/oVMtv68RK6vzMjZXwnIffENIBKA7MkBLiqw2rFtWi/
dT/3YNPpNxy0ZI1TIH3opKg+3hLM23kB3MAho8ISjPFaR0cYNENrf++HljvF8wTe
oRHJHYj5aUtsWvcmh77xL/u8xQQK+PT9s4j4i6/31olpEg1oywi5vx+rsfCMbU73
HhLiilQeK2GtGlCfcwiB6IfmP9V2qqMVSn+9DmQFcHRxaDWSM50y1d0/5rIhJibU
s8tSBAtsQoAlgkZ4GUXyx2ziY0F7z57lq6aPksUmz/b7xMr2s0DTu8hVtrsrsM3s
8V7qz8pTTrdH9UiYbYIdyM+7z1z0tq4510Vovpngklavgus1RGuLC95Re/AzOU3X
hU5GB0kiAQ/so9xgwpZOcR0SlsO27OJul9BR28tmxKG8gCSnyGeuAxovcHk3P9Kd
nV4EF7DKUy3KF66zWrPN9EkesZ8tOkscmTtMDKdNFNHZhtAmckNwXsqCwXca05Vz
lltBbguT5WeUrowLJxv1tKOm5RAVOEdmZUtW23o7aMDFe/CNm2jEke6Lp6FBgdUD
MMGxp+kbrress2pA5OS47MaqMN/yOJpoqI4cN1RHv5pGc5XX3t3ui1iWOAbbyjg8
vRyM36LCXwf4j9QXcjxB1dolecqi/VBG+vBrNnI1S5v8lk71CGMzIBkmpk1sWmTl
SosCaqv1lJUxStUCAtddIw4BY04cyODAjIlmZoJyZn842UxobF1eVPi1bwxFBAbE
SfHRIbXQuGSGpmsuRnKARTAc1EMZAaOtiLXRRI0RwC6iQP85jIu0CnevmtD4uZAW
UYk+7kZdoXlyxTAdGudGuQoHpURlZe65TyJ99sF8IOgz/aWmZnjPHplkZcKjJUZ4
paT8E20P+KSW6usDjfNE9qgDpzRUoikrssePhHbYBJuRhIn0+HA7XY15ly4vxAOn
zmJIBP9SJEwPCDDX6cAuSDTynv9ZG6NKfeoSCMeCSZynj9bWpQV1Uyd/s+ieMZ3K
10RDuaNt5+15H1jsIDLN9UjV2esV2CH/jWCTtdnQQlvRe5ch9dEmXsPZdhVAeeP1
Lliewy7PCpzFpdWXlbcpL65m3LJaDiwnNZZRw/AjBFMyQ5nNpug0ERGl9OqxeOHg
7X4VSvJZE8LSUEwV89kVYF55DINxLC1a1aTPC0D9ztPMLgs4Xb9m+cHxVD6rne0r
ZyPpGVvaYDeT+pMiXYTaCEtgYIfKhnBbI5NtOY/D62oV8Apo7PJ99J+gafKNE9TU
s0jjqKswimFFc6QFv+aqjH6WHhEDSxMnZN3lv6io0u+nGosi+szNMxGeGO6f/7Di
b1GDhDHGXnZmTAp4KiFPG2NvaFxKwXm5+u2u2GpNaFC8Zqaiq7zkIePYqzTwYlj3
yK0Xm4sUTE5JiRRPflMUQIqwNX/WXrBn5ZQtKkROYFuLnFDAyiNlS0vyjQYL8QYi
3aDhJPolBqJ+NpuIGI0JpmTrE11L9yz9U4bRny2aSoolmEskHuOG2P1F9llUYdzY
nhkkC3gJo4cpj8SXTAsheFFPuk+ejKddFOxFg3+lhQFTMdSZRw0y0pDUPpc6uBf4
0zTYXwJE4FVHLfXmTabI61OP7GyuSyFdFas72JhB0Il2H46fDMLNoiNhMuaREn6T
viMJq5IabyNHJ8C3IZNm7lCpvn2MJ8yIG+vdxwoqh8FGKxONnPpPctby5ONyx/Ib
ZBHDEn1T7uzr057kOYAC8oWlKyXqeXFzznS8CVBd0FnKUilTZNzw/qmFNjOExYE6
4JcGlDEsbEqv+0BB2pqkcagVKA4zKFbEayQotKMyqI/Z0szdRLx51AOVCnw1JKmp
vK0bSK2XX5RO0C0R91YWrQoyTKi4P2YKmKsPrijc6FM5ZQX2gLIB6ltXB4Sxz17c
woYZr0T7vAfw1SXq6ZNOSVD3aPuvQzMTmwop6bdf9e8FYnvZT3/ng+dxCLcaj+01
OpdZf+O0x+3AvFV9YuzSj+6BTp0ZjJ6f4mtOHd9IST1FONREl4DsdVwAnhGV6Wnr
EWr/wNrXFZI6aSbixPFR8cG3KOyNnQloO4QEgP60O9JBwgr8a8gIlH++jZiOFIfJ
nwQoB+ZPLpNCKktLkY9xVTDWJZVNprDMGNXcBP3z3CzL3hDlHL8vRZEZk0iQoAAN
9Ph9pri9PGTVttkBj824HC+CXflnpEEsTv7jyKWWJ5sTgAP7hx+SaeeXQsRv8Aqo
VrlRPXZKFpS7vRsD5xPTpCh6cd1DvwexM+8wUIw4yC1scgoi5KTt9JtdXnLClvEw
Lyc1chD9XspwFTdI5eIN7K3JIldQ0AyIM081S3QXEqqvJe3iQwQDU+N5GdCRY93G
JHL9hbhkjYmZo2L6QUZdlHPjzT/I1+K+HTQGKI99soRwhmyZNtJ56Iu2KJHmkAb5
KDNUrMs61Xx07IrFvvGCzf0QGP9FQr77BMCpK6Sgj3AVhe3R9oZsytriJDS8Ftqb
2ZFpzAvrtYULDJtZ7vFVU9K41dqk9tsJXj7njrwAkSwNVV1lG+uMjU2yLLFGCK2V
eAtLlRdbSHHRci7E4l6JRYA5lmJfH3c+SUSE3EvOi+7P6JC612LyRLxlPW2j9vk8
9fcXKKSCoXhlzZxiwv8Ov8EFbgc3TUnGijSSj7+PL3Zv2yFvdoNlj1Wl2mBue8Is
2VT5/0/w9mC0NJPuvqmsCcTMPuCcWqpwxjnATR4J6WjYmtMPNE5we1OTOq6dZqzl
tarC+PRoSQGjSve3CN1frYqEP7aUV1VPGBnmM2rWO3zGIVfNtRpki+oW6iq4c/vb
NG8jGVNBkpsA0wNonYDtoG4udqrz3ABRbmaymSxKw2m43SAh4xt8AjqH05o+G2sU
29SazHUkzjyUh9qaYRPK8+kGywEdcXJT+2IMDYdSRSGYGwI/77OVPJNwIhkBfV2D
aTyWSuYAcXtzUSY5uoL4Q4/IU0N2HkgC/6rKc4jyjgoBOTtZ3aO5EpZT04l13Lk4
NXPqzgLKL1jxLe/1A+hLCfoNfXtUqI6ilQRgiQ89bMrEgodjtkIAo4tVA/r2YnKU
aF+NpcxGLlv6Mb/lZ7S1s0GzE8bUxbxsUITlwMtXVIIRJGWVS+JL1ToY9ycBy7sK
VgkWQrHeNSnTJdMfnOxp1TtdopT+91rSFL+1viNJ603BEsbIWKOR/mmLxzkGSiKL
bTwoCqhafW2A9BUef5yDNjEetYLmd/qd4uodUtAQ7ixc1i09GuaV5AA0ID8NdgdC
b+C+tEwiu99Qh83JzFASv7Uj7sLetkoAPRfSiHWxOUoKI+2Dp4BrXcH+pxWNkA3k
k2ZWjNObD5RASDFGXz2C98O9jtzZ/rfmBmOh+kDkCcimQyjNZdHoGpx4PjuvAEGx
Tuzim+s2+9Y4p0DVnbfNdNL2ee9tC2I/tKYv2+Lbx0stqcWPwY3uAvdZZ/sF3evK
L+vTFNnxNu/NrttXbaOFLfzLS7smi39bNVeVEWFemO5TxyZNdHHGbeqA9TL16E9P
MuXMcq0r+PSVOnnEHH+6q1tHEFBe3vwBBTdHPRw/UP2Wv0st9O5dlG9lhB09U5hv
7wMQWcADkvTzeaIwHikD3p/vEpw1tLOG5FsG9vRzKuHUWoVGNaVvpsWmb6bHWrNW
Xie3gBi24x9QHZfdEJsJOW3/MhW++2gOcAQ2LcYg0yZTjcEK3S7MhlVAh8iMBFua
xYnemSB+3VB5XO+iLGpvrpSyI70K60EKVoRCuK4hjUZg3qgYPEPK8Q61WCjO1Ug7
CEUAb/2l02Kv9qJzG23sBDCNzkHIjRGFOAEnTFGVcG/kM0TkRPjblJG1jdgN2IlV
+H+vOmLOJo1J0kuEpEJ3rSjYrOcJFchtdjx6yAmyPrRhRogBGEwP/zEp/UUHIw4L
eiPjXYOJ1L0X2D1yrCLSxw24yIJOXOf8NHdzwuLcVS9X/LO1rg2r+jXYZgtBfCE7
n51QQDsLEQxBXP6d7+MnAKKgLVMFtujgmWQENOyae0evv8sAoQvKlz+4rXy7lfC1
43rSUHEldG3AfRZUbSIWempphh1F/K1ci03NjnPCMVw5gSo36SDGXPmkGuTUSZXr
Hq9EVq86UtfHwx8KaqUMANeqy7SJcRqZ5qBP5i90Cf515UhtodI5fANZ34VbAInE
i8uZMUjaNUstADtXDUiPBIBo+8ElfI62uFvwBxzQP/h/cJ/ZdCSUL5OXzCcxnm3O
pw7WtcoSg6XnfrSE3olQ7JW2Fstd6tiTmqFnoO43MVfwykgxxFSagKAadu0ImVQG
R7oiAPxjD8sWxPwynEIvRHLKIuKh16dcNeYlgjkZ/prS/WyNhxvi7GlqpERM8Q7r
iuDvmh7I6kaNOZijxS1i6Ld5DHISAENRhNvnwLYq+hTIwW5vqO/vxWkNIGaHesrS
TCCg6mqkAUMijCUWsRhUhhg7IOec5Eh2j1tKuEpijlO8w487xFeiaS6UdBMPkSVg
XctsU+VDy9kh+jtUZ7B+nEJbkaoBQVEdl9bTwODdLTUwLR4UQ3o5DI0DFgV4kM/7
4NFinzC6gxUnehpKkvbRkkrzXWWKrNW1Y+ITItAsdbGC48F2fGvWqCSRYQqcEQ74
59ReIQ5zGyt5QTCOY857IwEx12CpfnErIL3QYQyJwdq71vHQyQCifmEbcYb1/7OR
pH+J0XFCDYb2He3I9EpXcRxqkapNsNjhFZCREj4+zAzP3e7AWMX33NRgb8cdWa9F
tHGD79DPylIgsLG92+IePvQr0fFG4+Z/EcdqmH4df96LzleuVlNLh+XcYDC4wSii
9bW6JryVvduxE2jIhd60izJxYF6eXLmiEcpyZp5EvgpsJBVzCCbvv42ioTquKAJs
QMXq8eYFJyurwjqTnqspZxfvEnp0+fwHPDT8RtH3OHwjSnekilAUG18KCKkbBhwp
G2PN1CrS61wsayib3sIeNsa+tmuGKDd4MB/RNpgFcck/J21wpCLe6Tx+eNThsSQd
d4Z74p+IWwGjQXQ6KHkvY4iuVsI9IuFxgD989HpeSMzbD3IZ9BCjNECkPep/YdXJ
qTM4TJ8eacvxv0WV/Le8LdbzRXwiFIxX8dhbM7xtfPKk0SDw4aIElJyM1lG2Afaw
dcMGVp4sO6RlHwF3cAultLKxvBS5BJoqgan+5qSnj0/4/5E8O3flHGmWxJvDdiHJ
HK1p51Q6QPYVo/u/Oa89KiiNnEjfxSO5vnOTvUw81lQGAhs6deuTC2zpdRdMN06N
EnIhb7N8pnuoYZidKwXFBw3gRmhnOrqsps2dHOFNjCr8aD2fmfKK0xiztmhfww+S
uyru82ySX+opTw1pO8QzSMzh/lZsnZAbhV5s53vkDHMRPreN/itfD0jCZRsyqrsy
IjpjtJAtLjx0KhLX60G8qra0O5uzVzxMTCbZHrwHB87shEuatM7SUntCaIbuVGXX
4okAk2hxoOh79Eo+zcDlqN/4igudGt2qYEnsfhWxkmKfaQvzWHl794ovt2EBIyGt
vWP7+MNK8j9VfHRXC9qk4SUU5VsJDRz6Q7fHefw6bxsSB+hGF3fGRyXsbd52YWDW
Y5oTNhM6RNBs8Zy5cuOYzZx47Z0rA2DJfSrVP7cfXKO6JV1AxsBkQn3iXhXzjgn8
e2QMzXedaNZwT90BsQCFxMwcFY8H7SIo5pNCHL5CzAmuXyDrvh3BKdhjuCsqzI35
zChY/KEIEp0Rh5CVCoZRUHzD5UltCq5d8U0O27WuehBspA1sqrx/K7rp6pWdjypg
m34Dz5EWsdMzQ5QLVLgTA0LfIU8YUo+pxNlRncyp1NyYBSktKzHnZMxuihEmdwt8
e5uN+J1UUbxyTt8od9+bxpQHKSqofGrMJPF50vWB3G8V6DpI7eJT862Hy0qLTKom
HhjdEX/QePfgr7m4tcfd1mppb1o7SUAD27defMEatG0BFS1327pfcVrdyiwPFCCc
Nr1bxJE8y0EssemoarD5hRxTiq5J0+YA4JFd+qcLdTFmZ9h3ZZTAFUsOOdL7G3YD
MJLbxE4pCSjutT/Qv37GXIUSFvXNi3htAf8aUGCenh5APOLE9MdlKQqPL/O3xCMf
2gxSdO33KEpPlkxjjM61QbRNyJP8uIZGR3sY1ctgCqUBQHxu+t+4Ew3JfVsJMVVj
BZEzt5okqIb7DJZbrRYa7y4dH+xfqGC7OjIk/pRpkqE/SUcDYKoLz4ZO8vQCZZwN
xajm0lwvT4aNVCaQteq8hrCo3ZGQH8LYj4+XS1LpzhbpGinFONYdhn/ASO5OJCTf
JdUq8/nFtWemlt8yJBZ1uC+PVMumEwlpOZ+HG6OH6ANHHM6nORbSKwPXmrcqvrx3
EtzlIJhM4Pbqm6QVmU09sGhKgbxq4b5E84JLSj5INlZV9yeVCwaf3Y8gFTTLZvWg
p7oLVomb9Q5ZNkszlWyzWZpHmxynFyJp9KYBNhoSP6hvU8p6uIucfaWbAly6cMpL
IGLcZimP1liARjAcYjcxaZrbzIdYJIdMY6rLfBiV9JAR9kBYAYotFA/6Wm91sIX/
Wj9+1owGl1yWwpTd7Gp/mVKbgQEYUd/bBhf0gaCUaa7W3ikr0TGYZOKpIqMfCO1W
s3jce1Fk4QZ85JS291R/JiXJay+glKTQV26HVXr28MVFEC4olBIGJ0w5Clgz/y0B
2GwX+jHTBo9OYF88s8E4yf9GuygvgUYomypDoXJjRYvkgyl5UoV9H8E4daZO+nHf
VkoGCMnQx5bEie3lvoxsEMyebkUAo2m/b9tnwiySpdi1NXviGkDBuZHo9C4hvpoh
a7Jmc3hZxtMSJ9yhdlGN35KRk9yITYrFDAALYCX8XV+k7GdQg++cFLtjujShi9HS
/Luq9N8jX0Bo+tA3BGDpzZzEvmc8IIDHd6DAjvDPjDmA5uAlE0jtF0ptV401PIi1
ZHnJQohIT8IVql2BqyeZLPwe3mtrrx0ZTXIYVFRhZNzuUgeT+gvBK+mUPETWHxXo
KxKGMMtp8dUh7EyRjKsn4zZNd+NSPFuROMZLEVvlEq73TPlCO2A+cXpz4pvItorc
HHM4Knc4pTc3IIS8b3PrcTEdzJDhtdAXCYsoSkRP431ONmFJ5SPmo+qYLdyyIhLT
gbX6gGt+RBxEwhb1ovYzexndv8iO955vzV/65j5HbF0bWpdYO1K5FnANXOG5+nm9
pqi1S+VNId7t1d1H2IPpWp9URiIUdD1sAiQNE34bD7xWaC6P075DHQxUEcR5Z7/Y
0ZLx1NI+f9ApS5C5CfcgYwyz0VvgCjJbwrvhP4j9Cfpn/ID5oH08/gQrVfFqdrTV
GruW/eQfUT7y5XxgnsEcAfqMvFgLXZZZUuuCxTL3CqXsih+kBQ+vzj93I8Qn9TaA
6g3DgygVCS0PAkcrzY/YZjbf6fNsdbjbcuuhVz8orhXrnMNNHZFt5mjnM+pkfdf5
Fbn2oeUkJec6i7RHlMnreeofMeFFsvAhu0MR9sC3yp48hwXU+ratpft1oQBBMsCY
BAugt36i/+9t3dJv5tYSzvl0nqBOucLZ6TtbkfZxGDo8qeFw1GtqykO7GSmhCCLo
BCqlUh43HRgyXXb/k7c1Bqig8h4PWpAb94NTxXCmidu3OpCgqvFHVcZcRTDyDz1e
o7i4fBWTGrWexb9zMAEtkPknY47knPv4CbZtS0dUTMJp+70DG/VnQ9jBqFvhm8zJ
rse/IBrbPfOBuyv5SvSzGJLgSAQ5sl3LGSwm+bsOfffe3l++ZG3T8eRvN4Lcr7Qd
Ir1XnD5k98KmR6xmXeIWygevn2lMalliU4YZnWTePaFfhPEYp89RKiuF7Hkc9b+S
lRjGS1FbwoaMjU3dS7MDOD5RfY8fVRYn3g8O9FD/nJwGNfy7/0fdHGPz6TBpTBUB
6ZncIDHxBVxdmXCKNuqWyW+RXYJSmatHxLFVbvZMFyDbK8ZNkZXZUhW9bTimCzHA
CD96vHmsEuMk8dnXWK3Vr3APv1E+Jc23tiGrXcpK3PFszGIUH4IXec4FGZNEv9BN
39y3/rweI1Le5CR5rCXax1zRd/34mi/JyaQUYIpb9awxnYfcTbHqnEj93viSb10b
`protect end_protected