`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
gMcHP74wBZczB0bB0IzoP2xg5wC5NPjD/GsvSQ6VQgzYAsanETMwwsWi4yhFtJwv
5kY07u0WerSDf8woJ0stqW5xF501W3JLIS8KMiCOd55RHBOnavjYiaaLeu7oUCmB
TtTS1R4sO325rP2zOn9YwRbyyS5Ljn+PzFZZUmkt5xMca3p5NGqKtZW2dV6Babni
5HlLuF20Au601B75m2nv+ZRoGSrpkNElxoTibONmX8gBflpIVE7BehhHwaKSucEF
pp4QQ5zZAZjEC6aplZepouGVggAulz5AahlX5bf4opOVlB1J7IrgyjENtw6ysQ/q
DzybQ+ipztSXBGhmcCVU3A==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="jAI3OJE9Sh00Sic4PtM/KZ4WjwT98XM8AMZrZsQkxWQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hyw9IrFLPQsjvXplweG8O0lkaSLBN9Ijv4B5VdTRt6ipKJT9Kzsb5LxCKvkQyF9n
sGPOd5i74hRHnkHfYISGkfxGJCa55ieOyFShOsqTKRLxclm4oja9vTIey6yFm1BZ
54IDCG9h3PqfDiTD847UCSMRvFssyycwv+BRHQMQlFs=
`protect rights_digest_method = "sha256"
`protect end_toolblock="BnLuc3jxknmZOyxfJK70E5kp9u9O8IQ8cgkXv26kHA8="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 61520 )
`protect data_block
xABArkLxBOK6xG+7CdOOiGu0zbCbHMrEntFfAZEE/xRFxZaAZl1QLkuFI77OC2KL
XxG/mrHJzO3taVHgwRXNLDdc8ePbxbAiQfzV3NJLBO+gsBjmIymaCa480cPNpHLx
yhSJ8F+j8y4Swimb3b8B6Dpw5fMkCgMkBOV3+PuNnHw0U8YRl0ZJUZpNoGrr5qGT
snBM9zqmud6q3ZxM/Y+E1B4qgq5kMSsC1W1DgWtxrpOrNwMyuGGspH8SB6V3rsls
FPHiUGPu7cCRlwiuyHTEM6MCbr0nD2lHQwthKxNnNvCum5HrqrviGVdm4BJLFuJz
5e/SXNfC9TRzn8sMEcc74jWnRiaieHSbIHtNnz2+sxNloJz4xG55aAYKHVaJR55K
+UMfEP9eG9/rxlmcQIU0zuw78aHNqD43k+qJteU0TbIZV9+wgQ9FL1QCSYdojV+o
B+h5P3zRyLYJbJkGcW3t4VyaOq+oTbbPkrXBWoJ5ybEbtHjRN+8sXwqIxLYIPsL2
ReeGo/By3sQS7As1gXIIodl2UqCSX9ZSpFVnrVmBkEY8WzZ7dfNLsBR4kMthlhEL
qRxw7LxTv08HHzlDbwVNAIaV4U9ITsT9Ur45ouNV3KcvoKQLi2rkq7rnuZSipJLO
qFTm/kfSuoCw1eNKchnBLnS7DtToxEwml1cWtnpxB4b1USxQGVmI3qAITYj83ZCA
dG51mWA75UI+lcFuRl2taauzn3oUcXM9CvwPttS4/nDu2MAIKVKZ/FtJhXCZ8cXd
HSzDJvIGOwCUwKZmq77OIzwRrHQL0Oe+gvMcxpynZLskya+4D/xRZ911AhesWTDr
dLG84uRJYFgi91MhYwMmdYLO7XenVIHZ9dMDJqtTFtTZpRGLZ+XbFJAaGuPfeyrw
hg5f7yLjv9g3CY/dPrFQotYC24bmfTWR+u9tQvLG0nXslWmhBegV0uAP5pOkAm/I
IJ8JJ4stZR/3cdL2Iy1L7aXaBeYVzLDEgk4tHMsOCmOGbj6sqX0hVfGK2X5EjfMp
eYyNmF7Y8G0HUlsH3xy2OiNlzkIb445GXMajyBTdRfQ6Hmqbkt4PhGIA/ipOyMQ1
eu6oGb2kIaG0ERGcAVXiZC0vl9JRIulgStNCu0Mt57m+nzF3I/N5UTzjrVZ0GUGc
oELMU7bUL1u/zQk/e8CoL/2Kpy2x925dDkKFk5HsajkY4HdEWMX7wOyImLcImvQL
ark6kyUBoJi+WvSmmMgtxuJs9EvZxjI4NjSMFEbYO8A0MOzP2jIpq4XybynbtiCZ
4YZ3m4npbqpmPIvYicwzo22tnkBH87LDzssbr4YB5nZFuu9Pd04uPIiYgcJoHLcv
UBhzEsO58U0zhsLkOKgzaYDuAUQfO5Mz5drdY7bRTUxXKIT0Lt9ijcnE5QL0RHss
3pzsXqxN7KPYqOPBKVPgfSg0nx4NFCE/a/KkjlxGsEoiJyI5/CfAUv4r3nA14i87
dXv/75fZA726OY2IlRZLAwnoXu86N/s9Eimflbf7q4HPRG50Lzgsyol0HqYgWINh
D5x4cPEhWQonZ3SFexCEYFfjlekXv1uvhc1y7KyGQVO+oeIg8gcaroeNBf99iiyw
IMkFXHxynQv+27ssDz4eax2K9E1JJ9811rDAeEh3TMeeZyGBR+DhD6GZaaiMKCrc
jap6SeNSncqy53aOxherWlDiHO4SKGyqJ5vtEcMCDfJw2y0+4o8SJstBc4PB/byb
mxiwNaYICYiZyR8LkWwHHD9xuVfBqNn+A580D9gPeG0hE8By9p8aa+h+xTFWNk9a
EBBb7e/Q1wafXGQrToIJVtpP6rsCtentgwQ1ftW6VjNXGs94lIf8Y4ibi1WhSSFK
CpvGlzVIQ1DGXrcjALV1QFZGbGZHxl8mqtKBUdyLa5aSFXz53A6bgL05yelKp6QC
JwAV0LGU6Gse8SJxc9/aZxtG8WyYENsEIMkq3L18dVTSxyfg/eyHxMGCXpk9liCI
ltOUxRX4F3QuDuAtGZs1pAF6fXaq18PbiRpDPY36HiaH9Hfcv8xoZSTn3r/bp7zv
DabqRQqKF1RnOBSVksG59l/UZNLt5Ytx2reA9K5LEMN1gsdu4h3LkO1g0rqz6t5r
XlPk8uofsf8YyeUE0RRlMfjsOijuF/H6c8CYYr1flvnX6o/hb/BJoIGsukX5h29T
fUNHOhfnPqQqDwP0FZQDyOv18AjXKeFLGXMFtmr/CUKxMOjWZX5SQdwh9Cl4thAV
Bfp0K6iQ5LreO/gWTwVAhnKwoqyjE/I2gtbL7qD1W7ZoC3ycaW905f+hpiIuGcwe
jgqGNims8Ifrym+w6a9pnRuJJ8XeXMra/USn9kkZa8c7/WALjvn98hzhB6eL5QyQ
aCvy1m08bCTOYhy1SiLzOEv6Q7VM+ceIJl6c39brbnavppJ+yP8jnXYibIv2/AVw
h7N3DWYCGQqTGSlk5hE9u4OsaIVCH+o5oQIfcn0ckU8+dB6tcss2w6kV57AJMpV6
InFQwXTHDGBcy80YBELGYB9+ZPIsYUEs5YogmS19DYB8A0en426XxLwdzPFjJM7c
HGQ0W77fq17zofpuj4Jz4ypEyBy42P82I07j9a1XXoSVHREbgkIDSMLB+8osaJgD
NOjk9sqJuQa8SvpuDsDGfsTdw8EJmkMY7ctgsIfX1FTurFiEz+FiNxaXuKrjfqX+
taQz6Gfo0T9yQDpu4K7Xa8VJbzj7RpSwnxYVl/celeLepAAo2dRSm+orqKESChjE
1TtuMrFUuMfrzB1oSGh/Jv7CLaicN6opaj7Aoo5UgbAmA1oOKXLmNj5WMdwNFzX+
1srbFCQMxA7K4R16PgYcC97el3IozE+on00bUy2oNlnhQxlDAHMnv/FvD5qBOhf6
lk+kEizU+AUCYV9JfOcSX/zzber5HBhHMgnbrp9f4dfU8RzQGTTd67wze4Uh1G8J
UaMmwEiMQYfVOKJHhNeK+PA199DCGuRb+NfilEc/pBLQ7LdKOvysv55+zbUlgEpC
bA5e8KFgroPvrFQ8FVstMT+MvgAtZQirH4Bn7TpuqKQt9Yhb1AQbJAu4kABhG8EQ
MjZK3YXQap/s5fkAPMT8E+LV1KwHKBU3XIsmvN/crisHIICYMUgZzSXI5IUr0rvN
+tpCxLtQBc/5VS9liwgLINyFoIVAwIUbkiKj80TVEZawT7hpP3HKGy8kDyoGiXHp
HLxtvTUWy02Y2ezAOjgmcCikVYAhYSFwChhcSMz8xrEv7zaDt50fHGD85tvm6fiT
Gn7raHF1qXwJy6iR4REA/eRfPxxUwVBq0OAZtytBXFIrrfRFEJziIIVSRvSck4MF
KMRPP9LoxSaSQSrgTfLLmzLtfpRvpKAihgcc+K9iPatkzez3bpeir2evxS98A6kz
luli3kiFeL4s9zN0AXIMWfQY+ltX6Gy3/dw2a987ZxL+FMRu3ezuoxxDgpa7IjYJ
+X43YPBKwZrY3k882+OZ/mgTdflC2+J3JzLCTBdUU+ebJKcf/tRLEk/Mi3ICFZEu
9wcMxURQQG4GpXOjV9JJkp5I+Yh+aXKC8qZ36jAZ2ksP+krIzrZIAcfr3nULArJM
eojmnqZ5DqZPNM6uHVw/zbN8/WL5dJ1NgRwdgykcMhfo8x+m6r691U0JcOm2vESw
UFqjNESBHcLxYBsNCaIVBB6qxls3OO0waqxlFbMhx+bVn3b7FXUvnHx0kNAH6Nt5
H5MQzUIwKW9IA5qYwVAucaxUbMoUYyxMJK7e1+vlk13DaVHW7NEtC89NIpzgwtEr
0ycO1PImDQ4aX6shUY2R0fv+Zp77BY+iEhOTbiA0kTgCP3mXlmnco0b7BipPmcwF
CWqjKDWQzVxATPB0Rn28eM/8qar8hkGWHVnwtMTV3wdKxZ3NSKvw136oryC/ti2R
gFuZeq8tkw5AfpSrCIR5CoAup3dXi3viP6br1MJsJr/cE3Pr3LQHdZyowPKTahx6
bQSK280RiZGkyW4B+NUcilLeE1PorhIhkDpeFvWJPy87wm/Bc6T1ORdUnUOSu2OF
cc0bG6J0z+hXD6/Sa2oq7dP+IbxZy2Euu3E/zbjMHW07hqvB8wJG4NV40/ETzZJ7
vIy4Sv8oXHfwQl+QUcubj7/9pI4mS4UvI08aNGf+ale09itdNOgx/yCgEsyyPV4g
g6a12XBjDM27ZiRsBF+CJMJWfhuqJ7IxZvy0IXDTmVU2kiOtSxZNqc4B0lH/3vml
f3ieKX+A8PTYoKZp114/jZUe1O0eMrcdrafSCKEkLRGLGAWWbKxALcb9F206XyMT
6VopKZ/9mK4aJ8Ru87Clkx2DJ+U3W8Q8/jCkWhBc7+5oIp+cIcnlmDHDoywr/Wmh
tQXNXCQaoPB20DMARlMLsSFT2mlFgWATKyHykafyc+gTLvAKaEuSHZlbEnDR7fRN
tKwUaUqJY2OasDRZ7XywS2VJfcC0U5T3V8h0NH66cxjpDo95SGve+2RcuFJDnSed
rThqLjz+XHldvO1nKvSpzCsVjj0eT8fxdzgr/lgAPZVBpt/5BcsRFxrxOld7wQGe
w7bXjAD69K3tVYYmRgAWqi4xueNMuZ3wOC1MuSxCt/CEkeC6gO58msfSDTeyW80m
T/gtKYOwWJ/Yuun9vWOzkmfosbDlsneiGD6tLh2gcgWxw+o7mbz/Luqg2K29zzj4
QWKAdC8wJlcvHW3D0PFU2K1J3KrJZpZ+YIUppqY1YaC2rSsLhKYSJnqN5PqijPSy
fg8Z53MmrvmfTcaSfo0Ld2XWFaNHGt/qf/CroT90Zsx0ZPg/jiBO7QTFXUIv23G1
OXPrTuRkVmBE+NVtG8ZOm1xI49IZfPo5FBN0SjJZCgWluu1ws6By+cM8C6VXPC3P
2b+lJavfoNVXOz5xy+IgplRp+kRaY1YgRhWodyP8y5UKOb5ebr2DCj28nzlvdj1S
Yyi6zTy4yexHjn9w2s4aChVaBL2iPoKgdBbnvxj7g6cNj0XD5A0bgFh7OurAy7Ke
g+P4SxuGHNaXL81jhbD8qgVmQdAU8oESWmDTYtl5tKuXjEHrwAu31lJ6HtjBSlVf
0BwqEGK2QCx1ZCf5xth2Zc9BqkR1vwpqTtAm1hS68vHfDxjKng0tElDSKIK5OQke
ds4ktFUkVBcaoxVKtCX/XFQ+Nx4T1jzk+ua1uDu/OUgohamSS1iqytW3WxNi/T1f
TTRLCzLNApQEbJ/HihUTtONQIBBiuPYrg5ilLN916azR5vmmr7bre0RWutmi+B12
CV7i/TJkYVsgmiFs5IJTwZnD4jtjoLinFRX09Ns3dYZp8V2EW/BlEe+g3kqZaB25
FPEaBcw9ROCNBXk+i65dIMQMKpKdEZOZBh7jepqHXr3E4RTiJj4WzdcB4BYPnmtV
1mrXAOta/xtpOB8TCTNaarypbs5Z/NExG6mcfYuqJPV5WHSjPfBK2DYnGCrcDFI+
Mseeut/uAZBhXWU+oVO+O5AW8AqNolWfZEGugQ3jHeT/uJBcvnzVXpuxB2Cpq6dD
TbAsKrRAIhtyLKQGORNOv7bmAFd5vEgxdUJxzHwxmSSJINZDCrUeTZUmPsm3H+00
1fIVw6ug0fJEwfaV6y/nkG+80i0UhRau3iGMXkDKc7OLAn9NdymzKz2BEW0gSlgU
any5RGvQsCWZYcWM8ssnefRGpYwXMQ+xDEdHgJytnbmboUVQbDTR3iR05RX5zMtd
dUSe9W5t/Yqe83S6VgMqRyifZ6sm+HK9u0lipYg4tbB5otFXaWj/vIrijBDE0/4D
c5w1GZ0ObAn0RIW/pkijKPm9HkPp/mf9jgTvdvWnsxHKADccgHXAQHrUYojpZO0w
CxaD1c3mKe65oqV+BJ37PeL5EVjDiTAR+byjW266jw4GDcBahS5BVqUAI4m1LH/L
KO2G6uvjrIiuwFkAuOaNgxy6+yoZNlFNDU2NevLFNIyIUuwC15/sKkpjcm4ig5P6
4PX8t83ZFRkujRBgqO+9ajfE1meS5umOk1Zr1aO9F0orZ6z01kF6veu538vrAYYU
tvuEzst2j0ltasbx5ysQ6LxDumZ88+m4yqJABarJdyc6Z4E5IxZWWnDsVwsY8abZ
lqX0ilz3BfztCyFkYnk3iqOesn9y/rQkz6Apqk+X+mf01+/GnRiUbkHKvQVL5Rvx
zkUrLRN6NNfnuKpZQ2CC5U7m3x29hY3MKb4//KxdvNICUiLc/mSJ7BvVV7Lyfxgp
cVOxGib76RtDvSke0V09KCwzQqA9ZPWU4edv9U8tTP06G/3kUptSPPpfZbx8BYEc
KRjvues9l+zfxIVsTFcwChExypb6Fc0yosvNKN2wyYaPI8lLpPhgTPB6FgaREfH2
q3CgKN30fcBnCZZsr1lxFCn4h78/JlagvKlXkC62q3DzV7wavfGgqrngCDF5aGrG
fmUoqLdoIgLryQfG3KuPE4b0Nd5EgOlv/NXotpNdEVdIrXURsjA5wvo+WLePuHGw
eOdSWffx0kSmXmcfrUWekCwVPd8m0aQ83e0JfGpwmT9Xcx5nfg0j786UQ7G1jNU+
I7g1TnIkgQsKAiZ3qSGMuMKvrT+56w48EvXm8Pct4xBW146kQ15MuQ7PzD3Y1dOI
yM63a+Zhl2i4/Apv0kM8fQgna/2EioWSKqhUW2JN2gbJXpyLJTSc6nldf3MCLd2p
8rtsWBUkAciKgl/Lz83Phh2D1FunhoIlvJnHl2vvMwVU1TneNMyx6fyM9Pq/7ItS
ZLMwd6rA5b9ae/6HLdJ4h6NnMAN6nMrfYavc0RV9PIuqckI/UrA3EPa1tP5jrDCt
NW7BY2mSf2SPRV+Q6zWMDIpgWIzp/5HOwpiXad9+uNQuzRBMUmvzmfrQ1y0im/cv
4JdOejnuPi3aPcE0BbGKXBWJBuy5LbDIfmhPzIATtR215NrsGTkRbsaqyP8Kl+8F
P9OCNz9xJPK6BE7/3aJpcDJv+wWyntcmk++3gMbvl4K4Cs8Ch5wvurEP1mX+4tl1
JiR6N4zVt2CsLcore/eZ9HZ1nQF7+Tyzs11ZGXtzhdipPhXzhK5BM8yOgJSAmZ4t
SyH+GhsIzOqRjuq4A1Dmj6dkWnWmLgpf9KNBJDPRtuDXOuFiVNqefdl1w18wCGSm
Y6Ped7mIWUV54KUR1uXPfDfgedqtYy8n7OI/VyYUU/rj9LCcWAkr7y9pUU9GRESt
6iWBvJ8hviR707QMtMIvt2AUjwT9E/7Meoy/DZfdg3/WcjfoUx68uBKB6VNtJofr
9nrihWPoefdOagXSiM7EhWz1fQAOgWPVVaHB/Vqf9sYZwkuvejrm8iRHBoDvNNK+
NzwlrfIMaYusFA7wmF6u2UMKLhSKVWU+Ha1CgjFFvdel9sibb4SynsbfHe9N9/x4
u/pDMu23HT4lox5+ym/OlojPGpZsl+KMzb211A4f5iBn6ZuO0xEQ3avUxoej1Qkd
kvGyao7N6pVjGYEhUy9zbWQ1zZbt3CYSsxDBjIsvmFB/Qogc0IUX12ybjg0Uoqvq
85NOei9nWkVqCkAYAMjXtpcYDunkvu8doJdL+ER/rywi3glDk+2WQUkTMSvzTVXY
zGrUFdx3woko3m3igL3cj3lGFgrV6p7u9fgAySkI54NHdQrzCHYTBrgznxEYbTGt
HXbMZle7BTCgKPZRKWcCCfddtA1mZiSIkCXKZmqMcVpz3yrx4wFGMO6qbgDTcz0x
07WHgeQYc4EDwoai8jIjB2Y7Vn+CU/JffvOJhzVAzrs0niEuv4/rZCH5+wy2qlVu
lSCosJ9bsVYi5chG1nJV3fVAn6rN8WwxTpQ89YVppbbcTJCdi23m9AWwIQcXFg4E
EWQCjFuQSWnRH02v+zRxIyCFebNwRmJuJrLfsLT0Twb5toQoFeb+b3nKxhNoYnT2
NfrEHSi//yY9PMm8YFE7QlWsrCxfXIlh9kFqgi6N1sW6e9phGefoGma2kODUPzeV
2u/pSYhNSmvrwD+SdDrHgAy7Ji+8mLvlNxCGEoOFCaZugEDhBM0iHOB+V0wYOa+p
6y1CC5PPX3uM4MRiHEx+U0ilfH2iTfpZxbLNa3PwsOWm05nX2sLnZ7dI4RYqHazx
/7AmgUrMXBMi4mIMKDk1yE1ztVhaQ5t7lyExTWTErsDJJB+ZC1t+SJJdcWzjZd9b
XxFlbU98yKtSmQOHgClLHRUn/Hpw3coPEATBdFp6dKeg34ROGyavX+1vRnMzGWk+
s61+IWHSvl7KDBTUTRDrAyMZwFbS4xYQEoC0hD2W7F5CXkGnmUXnnPvBwkaTPGpi
u3ikUePXLa5V+73tv31ZooSqt6hJRKsThgR1z/U5CRxKFS96xawfDJlmNaEon8a6
BnZL3Rk8MiRu0RpXvdwFWXDXYklDnWOZ399ZcdmSB8q9q4ebGpfuIvudSHjC2FMt
21iVvrVkZd7LIs7nMAiJVjC+fRotfIEQaNdusoV00Li2QOzYnk9BpC6zlK7L8JQW
tyv0m4Gu0dBDZoayN7EfWNwLLK1lv01r16AkMnUy9f5faRiLgdNWbaCR2GCDmO5v
XHev8d14qalFX1xTwf+pB1/q3kTzWpyoMdQfzXO8gEcFLdw5kRLevq/ChcgtJaNB
3YhJJnDaITpj71+OtB7JkFY5VtK5dOk+IB5NOliQ10XtX3xiZRqnWwy9cFwA2T/0
3SUA15PyMcNG5D9JiBAWnpS0SA8U8kreMDNFemiKGy3GkSJKboJ46+3W69khbJDm
5BDpZFbi8t+6iXWTJzYE2jSe3Dxa3LABLxffSnPJ4h76lPFw0EQJA07cQ6ryaPDs
kUJY0uatSMrHXPUYlDtQ1tZLm9vPR96ihRW5pE4sTbTOCxjbf+laL+0K6jbkEeOb
Gt93iVAdSLTZsvYrsgGRHQV4OATk/3V9nxtJ/lxCxo8cVRRdnTTZTvpLe0LakYCg
vE1kFsW3CfIdm/NQxgXE9r4Nl5xduBmkDgpmFetRvxIXFQoGIKqGLlVaepz5JqNS
rRoabIf0DIumJHlOR+qUymOL7PMKguiH+BIOkILxQtsk/AgBPwLVA1KiWbUaWVag
pOTmCTh90wX65GRMCk+97fNXxEsQf1OK3Vbfpl9aE4YZo1+TBqwnikHAe4JSJRrF
pj3Uk56Dt8vMIJkYsYiRiRiHcoStpJogqVm9qlBfNav0zMgIy/6l5RvLpVME4x8X
8pmt9Vc/tTx6mYpEB6rO+PeV2tC3WN+cAEfkh/AvtZPpiL5YyzBI4+QNKG1/BiMP
13GOTEQP9zX+HnWGC1XgGLjrZJRE5swvbWTd770OXl2zkRNvck/YLoFTIdqv7R+C
o9gESni/YUSav4uQYCZ5BQbikK21m0usSl0iqaBsd6ojs6EpXWz4XU81xW4AT3S3
EvP34+D7PhBYtSZvag4MG0zRWruBYAbQpfJWCIQXSt+ksIqTe64vRXz39dvnLP4m
1vO215NAFjEMEat1mE30lFoxz+JYfZK2zvPGL6rQS4g3b8vUWHY3nfEEpj2kVoHK
uB9QnSkY2tX8/gLxiCUbJEHrwjubKGa2Ld7iElU93/cTTrOMZoKikuO2dBC3sAZd
1ErXiGifDt/F1Ev3uqoYuin12SsJr1icNDZLyYSUdHVG/sBhFTo7TmoTyuCYnC0P
uDe7xLOHqoOTgZcEyjA1LUY2jamRqek9GCTjue2zPANwN9EEc07K3cQRlZzjEmRT
Cq1IgBZsVymU2OLQCYXduSgiwJ0kMPA3UPr+JbEdoJU9JM2gRxwFFWmgsQku5rWZ
G+dMjrW6eIPXWQj7v6X35TJhWtOO36d1is4vgWoWwjuXJHzujeiLtpJg8bvGM0tn
b893K4bLvdTPrW+As7QaViSrs9wLV9JIQOpNSCBGMXmaRRI8GGJRRb+FCKDz90FY
pOW/GEKigLKdsPaU3fuOi8NYo+0Cr04gySuEOJZW64J8W7SmzRLW6oz0NL3M5Dyx
SZY6Q1b6wYtQMCJHlWiX8dNdku9KtiQ0/i/hsVAbE7W5SeqBrvfbuOn5HBskJg3L
SYbbh1IfCfVJk0h42MOAbsRaiFkELq8YFGr/8pB2rl0A+Y4dDwnZDQ2YkWl5RGfA
bJuldyttaK+EMoLRGeyb8elZgWb4tyPs8Ejc1AFrOTspuB9MD51HYoZj2Sztpg1O
WPdw2WVluVgCIrb/F0Q+y62gRYSDrNk72F7lZFoMXS3IZ+I1z0Hb+xxdQ/Xus+FH
x0s7CAutwoz1dRGBXZk5NU5yAn7xpSM71LqXb8BXC6b+pn/v/oR4UFAk5iRvOtEj
ndyTrxZrl5MaFUspU6lrpzCGlAb7LVS7gzn49RSo/SWX0Nam7Dohs2L0/hSEORa2
I3cq782kUr79S7aANOt4LG1rxK3/neTz6ToVw4xfycHsZs9zC7n17unptmRUn2iq
FfkCQa4ZTfB/tRT64REYrhyLc9FeQKpM5Z0jSmJ+ebbzpxRS+bQJPJLRm3VX31AX
pFnLIoO5d1ek6xHCjEMkWCnb6fZApBiYfwWrP1QE18QjevX/dv7HTnIRwqOisvk0
6mm7UQXVqry+5H6fJawdorTcsWAcyAukEQp0OMMeloxKq3LwZR2ulu1nlcKLNlm3
J4AhvOXUnmOL5b6KM8M11hFR5AP0gwpsIgsV0qD9UhfKM+R/Rf3L3UnwiBwqPBd/
c3CkrK8zOOTGJRD2w0yJWpbq93BiiorvZjbvGQ0iOoDft2LA4ptBvX1ll251Mxw6
oqXer9uqhh64lVfe6KbaKnlP2RV5gcMjhX9mpUf16S1r9mjFfsbBTVWS8umo9zWA
sDpCpshiu2KKHBR6AJL929VnHHZ9ixwT7ZJyi/UVEuV7JJGXLGhbBQ1OdziCBp8T
IzV+DYVnXezhTATlwiiTJQbqVLKZHINnyQZJ6W29Y+mP2eDTS3TWqNeNg/rHaXZe
R9DT4ohOuB667YQ2E2gr6+2ZRp3BeNAnb5FLxDwlgfIT7sbqsT4q+cG437N6JJF8
PCK0aSS8UImkqvhgk0FUNCH2gy60Xvx2w8FKLRYz9TCRkb1joree3RyCsrfXNBTe
5WvTp+FU+Mlp8mjdbrtEgxTPtHPP1mAQJS9/tA/ZjaRLhj3T4SO6SqGJMTPywoVZ
Eh0ND0sjyWGQaMdwpB8uzOlX3rJd81JZLZTx00uQb2x0IXpLOK8jACHtteT3Zrmf
WaKsseDrcb+kYODaSYeaAS4fsVqzKYPxKxN9gSlMbjM4rvqrGAC2Un3ZUwvgfm9c
YCyOLKOa/zFkBlDQ+jiW0rEy6mqX9qeoUPWEv9rpBHA1PqEKey2qHXi90ddKeOZU
I67KFJ7IQBTcALC4IlmCaDzcw2KvZinwkQPpaxCKwzFwqirfeKcPLLcu1ibiXUcR
2ZWToD1vnd42wDEqke8hPOiayp04mnyKBoNT7TcaOlHKlx2PTwrXi6sO8/ES2UDs
4kah7PmftuXgeZt9UPDQIXt5P2tpR/h7USsfctT19hrJD+FORyHskziKUTHlGDJv
chdxaeNsOcXP7Jy36gvBrzovJmqugiU2bdID7ywm7rfjw2D0MWfsQeV8IW+wfOG7
9uE6VLlBgkszIof7xs10T7ywsO+BG1Lsp/CHAd+BMo8ouAjHPUfHMF/Pw5XVj9gc
OSkzBQkuww3gvOVpRrelWScX9sIBSXlJxOqd3i0s8DhF9Lo1aLl3hkVfgK/KlRj1
IN8Td15vC/0VbyWL2yUcrJJs8htmPA3nT9G2QpNKoUlZImQiDH0tJw/GqMa7v+aA
a3/vrxXMWE9QHPUgXU9JUKd5GBcqXcqmKv14sCrRT8fDOZqvnMPQYdZjNOxWXl1/
UXMSrE17BfMBNMiAcygdOEtB7JbjzbP5zjZ+aCHmKlNBW2zOqQeD7Mo6J1pFNB1f
F8dZfs/5RViKcMdO4b1FFIpHka9JgfJxb99fKvRl1rCUMCi4vVZHafTo/HJretcL
nKgLwu7OhapUwReukoWDsG7ouZQKV6kPCB5/qhQgkGF1ofLvvqO2wKSRt695BsWH
z2xcxiYads/USrvylU0GEcw9b0lbAqzSs2LtrDLI68dAleHLYOIeZ2RBBkUYQEwZ
KeZerlk3q2VcjJH4+GyMNbwYD7AbrB7Id5D+g+BgIMgJMujx+a80s9gzjjO3zC2p
hE6yZdotiNMJaZ0YPr38+YVmrRISUFvDWHaMBmcZJVLcni5UntGs0sTAgnZIbdDJ
eYXrimWXkDZokWfvAzVy/3sTiKYu6jhhgllhJ2N1KDdWbFMEfKixrxBmbbn6Zm6X
MHUYA+hVsMDIIK/HxC+voPMepGdDX52lWmNqlktbu0oVxo1H22Sxwp+/tMzqMpYb
E16ql+P00GAGgL7PNP82GCslpxHmNL65SOLm1hj1iUhknPIk4OtObdpYqRlXnedQ
Xni6Vm88nFATi/52A2UxNQSNTMiKSRp8nRc9cmjHGAlCIJclVg6aaYLHMK9AaN2T
SFxexmWHziEafT4iF/TQILXgVN87b26wj7rW8RP3O5TRGH24St5ZBU0wf8BdcIy+
B7VRgWblO+zkBFi+DqRhhyMH24JYMkNSeF8Pnz5a07VAVhV8y9Zw0LQvlNxrwy8f
v3dUytBTnB0Q2H6IqW4bKuo4f//3+hvEIjkffWfIhULxcdetpLdd1aLT0dFTz6U0
+fGGgPnowFPStRUNahE5D6qO152wAAvw9oyoEj46FW7c+xlZZmiomR6lPsHRFDGN
Wt8i3ltzofMkY4i69OYrbgatgce5cbtfWBG2QdUBURfqRnNhNMA8axrq5jPMeEph
rFiVBY2aLQQ0LkvI2I9x71hhCp+Zx3+guT5BruRGumtrfKnlJeB+m6G5RJ7ypDXc
zUfXxZH09J7cm+uBG0HxRYWL5SrKbEcOqRSu/f04Kae6Ifb73ZTWSlN9w6dEvM2X
6JkTQABfLJNAkjaRpR+cUkbIQMxmKEPklnWpaptA/ICpPminzDeVh1KSWxOTv8IF
5LypqTDKvXzfWm5SRtJBi96qCOlECtHGD/9rcUaJTd39yz9yIkF9LPv4bmj+e/Bi
itt7auA5T3x65fHIEQga3Op9Sgj8SJxOTrhe59xhc6EQDap4NIV0BfTMXds4VfXz
C1LC6CGeoKdHtBo+ZTRE+4ftPGNjKSLeqrnIV6g0fEBa3FAQDPc0vCcqtB3cJNp8
yIfuz7181WuhFUf798imXoeh151po01VvdDaL3lqt5uioHeZH8W0cmeHtdRYg0x4
ScMicsGX//fxQiemuxdZllHz7693JuZxFoGepSrGbWta0g0CnBN1Ii5mF2rm2Z3z
0n5mxav5tXLk+DqddHUJiZJZ/6vRAqP0i6oVrLCL7FWId4qhzKEzK4vILRPhF+cY
DI2QMWYEw0Dl52dVNkaKkXh8UyUAPKDfEkoNyAi92tJoacIwm4wZFms9/i9iP4rT
I8/BOEDs0miX24D+R1ZLfxsYvgtANn96F0gLgXzKv+pSqLBG2zgZqDre6M4NjF1p
sIfQfUac+wPlUgDhLMBLmZphHaZ/bGjJZX+Ilwfo+slquIwZdHWuo53i781oT7+D
0BfkdVMfqHYAdQceS/+j7dfTTYKvYRBAKQB/eZbOv+vSkYmT6x28iLUma1Ict4nB
Yu1PVlOhm+kYT001UVfOPzIrbYEfc4gX0UJfFNJhgLgf8gO4WjChK2ssm7a6ueIm
uPQZFtX+v+95noGX24uXyHY6524sUVpaWp5IL6+X9PBe4idpzF+Xh4wDgvbm81rP
qhWMihd5BZZrLG7/384ott0+MrL6lsPLjif37y1AYfmAQb+HFFrbbOY4d4/3LAXc
yuHq0pdqnoZIzELvRAf5sXq04eogBHtpoEgmKbEVoh8YUSsmZasr0TDTLIZP+VV9
0LFRJIumDt3/iz1jNAG6icAjAbYgrdmETx6fV4tZgKCFzNzO45cUGz6QTshQdeof
TNbBjYle4swDJzWuk5915X+c7mwHH2AYw0VQVwcVO60qqsGUbwdztM/qzYMVXeDT
AcMhtHQ5zntZr40TdjJwb4qe5I8NfysSU+ndlGcBTQ5SNqCsTPUs5EZANgsykVT2
ZoD1rgNk4Y84ZpW2IlFeYRaDE2gMQDnX+xLJf7zKE6UF/VPQG9as9jn1Gob7mEUY
t6qxA9oFgzyyr2FVHjHOivsO9tCOZwdt1re+fGJYy+sKUG4jixtaBKStTNm/4uYM
iUH90DLZ6RLXBeFxIx0JWvY7IkzHuSFNvfbSIWeFRs6/6zdt9Eg/0T0+g98orOV1
lt2Q7rK30vlWWplc8J/GE3vm5KqubNWBQdZxkHCEg2Z1w8uf+Nh0TlMTUXC1C0FM
IqX79nULqz7Z/6WgSu9P18HYmz9Cr0VYdw1aEs7QUtoaeJSqCFEqRY5/Z5K/jl34
uBGPg/h3eEueqaMjfneSr+fx79usLsgzmVg1eZKLN2Eq107SgHqYzM9zT8SxLeJE
x6k1xjxx1TaWNl9whIwdpNbEq6V0k8qx/JfIN5LqrlkiXYIfprOghJVBsAqEv8V5
lqpo6PXUl6m2tWjvuq974MMDtAiAdtwIe9hugSPlRGnSrwEuxH2r7rcJW66E4GAx
zI0MJ9L2LG0T6xePQBl6Oc8n/OR7UtrE74a255pu1I9siHfu2BT1UzlQPheZQ+OY
+omuqtDEQNw6F91vNXKFGbhlR1CcbAeQtGcKcAGN7oGjjuvmuegeyml4uMGVUV0w
qAFF8t4BG2Kr+DA3+9ASXLWiZK1dpvhlGziKdq1AHQImi6QteUTuygy77g6PGabG
xkB3VSWm8h7a4nAVkATkudtfy3BkVvnicKo2LQAhoPvjsdIZPDc1KDuoQjdWCu3N
0/xwarviUYSiuWnjBO4PzPV9uj9IdSBifjxQknRPNjeYI59gVvp9RllGWb+kRx+m
LnY9QV9WbENF5HXgQGgR3rsB2DCabx1xkf0o2G+iNBZQMhnvkEAvV7/KaHTEQ3+k
SgMXivLnIHD+zmX4K9J4p4Bta2zl/C9dVWb/533KL9ZXZP+8FQLEMJMOjk6FCYy5
4Pb3qLuo0iNqAeBmxYmgPXzD8rJ+/ZRClSCS5Bx0pIsNucTqkXiJL0oUbFVsRytc
sIucKmbxe6YYkv46R3bxmMik6dXIHjnHo9YWjoNDzZWE7AZw4znD4NLNqPfZEsHa
vZGwOv3TUeJkWrUInODrDL93MfQ5FE/bw/7nMyhtbpcbxZAFbd3c/h7ZuuB4SFuN
U2DpwxKUhUxCumBuw2RzeYCHEvf1zGKolQh4BkfYsnYkViB8odTjpSCEhBcnVPmA
AfxZPHRQwtX/FIp2LVP0eCkm/gXibHX+DIMw+qqqQnDgnfw8779QcaxIAT8wKRzE
T3V9v3DHu3UZCoLvsT8PS9Mw/o6Qd9/pWgtRR5rL3SJccXvcJDYRmkXNMTR6801K
kr/cj3XB3fNMqDmivcctanr9fErzmpoMOvLn4sQPmfCvSpAlDkXkcbn9WlqILNyB
yKdAabd3CKq0rOYsWi5SGILYk+COjMA1GoWakxh7gQrUhXFOGKgJLlm/ms4QeE9h
by/LDGmy1WfiyQ9hpfjQ9OMUjqtMfpBbNxYC2shkNQ8f2p5Om99Si9KsfE3qOqU8
0vZZ81L/mZSzzPpHzCmD/P+RHXnHuDkevmMfgGpqewZvcfOUZA0X1DHiNH7rl+NQ
1IfVd/uUBmCJcAt5SJ8V+iokTVXNILVBgQtBGlHpHeE1R1SMUwslZck1q53QojwC
EHVIWL/wIvusiWw5EIT8ODz9YGnPl1foK6T4pT0dOY/UqRBvVErLjKIgbgBE9WRO
bo0yOOetMttldqeK7PnwPiPsXU8JqVJQj6N43iNxKclhjngqJPUpAXRepZJKN8zB
CIfDcL74XC59FRyLg+NAsTFWWbawmwnGoEjwkbnQTY+BYhAdlhAv9KYWbNFoP61h
PXcbrv5JbprsFww/9i0SBypwcoWXxi11l6f8XWq2RJNXmUDp974JMUmRrjODpdLd
6JkfNOoijV/EpRffUbMK7ldffeUqaVxvfhRo+pkvBGcbVA2zobXxFCXgSxlkNnDl
id/LfIjMiRgFiaa8oZUMg7XDdxGNnod9BU+D7mSAoLaUkIq45JP98uoI6o+nysZd
RBjpBTtE+mi284IiaA/Gdm8X3d2E8SdphWEc4zGwZYGJeDsC1L9PreuUuke6GhjU
k/YwB61ZrBB+F7aC3oE7vErgxKBAISyBzMQD/ZS4Zh7osh2CBrS6f0bl9jYtbb+W
KBc6A7OLl0kg6dXC0PrdJjhkVeo40ggwWb6+4ERhX4Fdzf6CKhX4igCrpZsyS25a
ZbkeyXTmxrGitKhTS9A3FNF3R6DirfxobqiFQLjzHsIpeitShRgGDW4dYroaMZ+O
hcmMhokPXziV1ycLmqCMOzmskTpGLFCmveC9ZzHRzuJfQ0ETgyCWxQmVf+sfBHuL
wmyYuo7YKNEKgRh+pgKWjDZ1rpsb27g0rv0rMvD+qnn/FPslPlG7tr3JKxBteAbf
aSGqrN7Yi9eUzVi393CzwUqhmlNTwahq/xO0jmjAdh9yl170yPAKEqp+S7vgyfS9
YZKnKtWHN/LtaGsW5wHGYndVc8spf2N3yTXfgJLY6DJRDvwkS/EQTW7P6TiSFvh5
q/OYPriuuguTiZbTV3qLa6Yrm7KP7vjjEkHJ7DFP84IZNLMRf/cF3e0oTS2Pm56g
vEKSMAh5NBHa9wSi/hZD9a2mht2xO58S99rQNBfamuHSNxwIt0lGCU+ermkkwrO9
+G22RhSRgvhaCCVR6njkQ9yjVrJBsJEywvBAv8dD8CIp5datfcYl/xm83I8XzezP
GneOY3naEEDxqOBnK6/Y9RuJK4S690+HFaBFsY2X/PqLvNIwudZ68CkVxXSKv/MC
6K3n7A8LtLOXE49JMGaNZ3WfD4aO70OsFkMYbV58glaXTeKH4oIB/ukZ2+n5Mevx
bBSxX8GJKBoFshPEzOkMzE01nbDcYMN2lV3alZMcuePl7n00j/2VVKpSe5fhT2S8
nxR1y4nNmM0dsoXRpsQiTCwc8A8BAJmR4cwJwQMc0JSZuB3IHf3Ib9Nrx6LWHqXW
JaGre2JbFcJqW5NLr6/8kDmVTgKXsN80qfAMpsPfoJk+ZogFiRhMuxxBzjhti1v7
0ln5aAY/rdygjw/x8svxq5YXJg2Pisz44SJ8CFgjn5YBBXz5rPhsD2gfh+40VhQt
38p6vEjUVs4A5KJuB7tvFvJGiP2qc/NMOBzoJPW8zg+6+WZgch7TtJtNFQ0IN4Bz
p8TqYGAG+dg8FBZG3Y/tMpgC3bv2CmZnhT66yjEvL5DdbpgcwM5caMCG9hk4QDv2
g3gzGuWYLt/JNQsWs2V7wT0LDkxeEMxY0kYg/lCmk1mWCHcEL7monvAJJIRT5p4z
ANtBQWvPGbZM8vzo4wBzK2hGmQmp+nqqa4OlPWAGxDfoLugijDj5F54OvWqWJjfa
gOiKLnwlVTukPSHz9v1k19DRwd+9wOGjNc98efrerEPAo8iG36r7QUTY9kXtHG/6
2Zrmk/wYXz+CkU4RLxQw2Ph341/Bbb+NtNBoQ1rZXUCYL//XIS4OslW+3VMcr77s
2slroAlsxcKiBUxGKmaWayUkwvFXH/Ke9n6YOEpIDF7eAJzzPDsvedEzX55UUwSr
L2PHZTdoVkVLTJR8X5Yvfa7pSEIqOpgC0VJ+XxZPTVp1zFB3NA2zL/ruqOx9i2mR
3aRchyZYr2arWKgujb4ntUD1xG+Dc/4Zvs0Kw4KiyamfNS4DIPRV7KA95LN7QUQK
46gWQiq9t9KkKA33Ll3mCZ17QPEZJtqKDdrtayn2TrS4PZcPxeDmPqo7ab+RdWka
r5EvBM8HjJT/p6pYICV5/8BKc3gmf+ISV+82orhxQCeW0coMlmRgsR8UXO8MVr3E
OQQeb3SZ5mkBDmKhoR51B7l/en90GwHPAwwvd59pUtt/QvA3SI8GTAlyKCPql97g
GINIZ76QLEalItizuJfEC7sxQ2i4SCI4SmRD1dZQS3AwchJSJLbakCn3tAEJUrCK
LwtYLB0vTMKY/1Np6yijlocXID6UpshwqZyasvtoqMj5siXBmHOYiy6QGp/8FcLb
lcmTcmeWdZcJZcFDJZN3dcENHZNCrohWQu1UfF0pRCC/mtH79KiISi+7i1cZPi1Q
kb77VGlnBGX/f+3oVrcJ0NANvlwqCKxJK3O2IJmGxMvQRt03HuoD09DhPzywJ8Ik
lpN9jsP4r+7TjjTropAmZxTcMvtETIYJABS98PY+yYwAXy9YbQ2wcp2F0OlSqvXl
ekfMeX2wWHJ+kCkkz0FYF3JwPQ28wH/rmUduRA5fFavtX37Ubii+hdVLeahLaFHJ
y0ZE+XMc/7eTbXBwIe8LMUsIkdpizvjyyJN9EI9IEr6HNrztZa/kKkK1NLCcK2cf
Cp/zHHtaDVImS/5jYXjQGBCJcI44RahlotoqRCz7SN4Tbix0iQH6z47ZyeCUzFpl
xG7onlyTaUAysqzEvIehH8jkoXUCTrAPXl6dXRMMgJ/f5hZoesqND9JedD3zdgyd
szSCXT72C2O2IZ7JAl7LuNjKHj+ds3vlips3eomf5EvzZll0QvHjmniRetmeMqRe
d8LzzYyvTUrXZZCd6j3iDlUblRgwOrifDQmRvMZd+tFTcTF2uDXKWkYYWT5ajQSa
HdNVHUiRShQ0guBJsMNOT/MFqJwOL2G03QGSmPLc77G7oAfSLZYJpcHoKv12UJI1
jGiW5UfQHsPMABBngcXmFiqhLchhiEN2ELSXKUNQq0EmH7tCxljV8RKPFQwR9w0E
5HTmumj4rKg/hszm7imRRRk/T4Vmvw8qhP7s3O4P+yHM8LrJ9QswAyoz6dzR27Tn
bf1uWl66DtxlkvgtfewU2VjV8hChuJfXqE15PRcS86So40VUV5J+q8WvCnbz8l9i
UfRviaZWN01E3N2i/ybyMLUW2j3yvD3330aJp+p3hw/WX3jjP+VrT/oVT90RSmOU
RtGD0s6KJhTeqB2UlbZP5+X7h/n38/KiqkffDjB5BLlkugm39PzNhm4X/qFrrkIS
cilh7Ko6gai99GKsPWF5yFLa6fV/W9YkfsRyEds+eQ69SjXhCKfJx2GJfmmGrKNh
Jk8APtxrZlgbJxsxJ8TdR8Q/BHyBfYUBG5mTJzEM8trtwdZAC/e3YtB3XfaXA5JS
f1z/v2wgp+fBFfy5e8kFemkmAlFLqTMxtYvvhtyJsErdu+8oQwbVD58vdZGnoaBY
0t4NPfM9P8wuQvUxLaDc2QAh22xW1tTFFqQ5zOljpmWs9u19+5UxPejIYbpw1ED2
TrYh1aHNmR+owjkoUXpP2lHLLkbL8Vp7TQmq8zyMKTv9SCfwCiYF5HDxZJFnTd1v
t1nqN/PZjQv4QcxUHrEmjxd0al7+nhGhHhSfkOtWU53sMHDLd2DVd6lamDoQ0wTE
vrJGRbiXw7E/izQOZlI+wvYZ79dYkA7PPDdwQ0XTicpUO+AmowiIfBaM7wD0pwU+
TfSHdLp056nhyydUewSI1mA337Ovxmvuw/rDWe6x66MyIrixxu6UW23jChFEgEQJ
P9QJncSswvpamm0YhN1nEZrtkl/cFKXtB5N9dNOSLZqe+XKAaRlewOYR+wkJBh3q
VlyJ5t9nGwp5Rv1ap9+SbOmAgCZAZ7PLFENb4Jgly+inXoa7fq5dzB+TRzt0PT6I
+XhrRDYTAa47nkWlW87mLM4oCUKPOosjxz3dxdUDlZ7xBg0F6PgM3ZztbdJe8OQX
EcWzkzJggOnCsjQ0qqvi6H9LUrwU8QRDDuzynhCIY/YM1wps4UHB/EgYHBipbJqC
vulFtvfLymydOEBrklzcSdcSB9pZ48loyAoPwFsKzWQFnoV2WAglGtd5jRN0C403
rKONaHXi9euRLMwn4u0wYJM4vIKLeW5nqtFWGQXG731m6+B4farnSnE0CqFhaF3X
WfCshqqhOYAU/UGycZNV47AchI1r0JNp4a0yrsATNKmXOaphBw6ji6tAEfpixS8o
qk/IyV9TneycnBGQKoGPWBi1IUjWUNx50rny+VtWzDzvO/lRm79g5vg9SCH9uLJr
sxgftwyz4zKkk+C9qx90i6OEb/Dz5s8Aa9dB1sT6DnLB7X7eL33eFHlPSSrawDA1
o8ky82feNQyHqw4i4z5KU1ecfanLtiommYpTtgrg/aKi4s8WCGktfkwoVKz7Ir4V
vUg9KFBstPZEgyVWyCS37wG50H26O5gsfMtDhBslKRRDSzQT1LKZdCxeh8jvO2sd
Y2bM3hKNId6ofc8oB/bNJCR0G9T1EgUm/otbizr502bUCJJUDqPe8jjfvdrMBWYP
8wfJg53IewqgRpRAAZc5VdgFJh/guSUnuwZQE9fJUlP6euxgOlGqXee3Bhgv28kE
iQAs9bH1YHNhUvXdwKKDf6fKrS//uQKGVfaaDvn5kalNqjUv9mdFFOba+bduOe4W
4PCfGEKZjHgYOz8XH5tLoypTBUVc7aLUWOr64Nr84hrMPXRi/bQm6165YrGvi0wU
wGYfevTDKFP0YP0fLdx/YZo9VwTsIpAfBkCH4tUvpPwN8/aV9FSMRWiRXHkEcBI/
KHQpYMYkgoGgE5EVAAm55DV8zY7WztYnJEB2A4gJvyWU1Muuae+e4Dn2NW9/djXn
ZeDfpv5JsMlGDkDOQPdOaq8K2X0VrCdEl17QsZvVFdhbhS5bccdtaG4XHZq54jYr
oMdPO+KxILv3jnAuXxnKvTZxGQuwSJ8lEi2hvLhso9t5KclFXwBREXTeCCRgbFJK
lPbygFwAM0a44IkFa/PExBzISDJs79SZPZMCtDWP4eKNmZrFr87iy4TLu9XsrmAk
ccz0ET1S5eLbw3KHfWHoImgOhCCcFC6n6EXTTF1f0gI30Q+OKiJ4lkKvYEwKUr8P
z5m/BcAEJ6YLU+pFe3OUl5AeX2WTzT2ECyp7yDCUza/R+CyfiRUf6/2fH2xIPEuz
LZcGMkCZ0m0NZNbXG/0xJB0bhqTi09cS8/4CjPIena+dGSMUs4p2hzPLJWWLVfu3
+K/C5Vk4bBreskGyW35YPW5rY4GS6BkTW2A/z8DyJ03+4ZC6tMw3Rt6QCIoa+28+
Ar8wf9pBIxXCUeYpQnBFsVzIZroMHRzCwLLhsR2Dv/Dni3KJX9+NSHryMZ+f5baB
+Vzt37aaFHNZw88rFxZ/I/b3yMi65NTUz8R8SCGwdILlWjGNzUvqi2yE2m0x4VNt
CduL9AznV4iRI2c4/yHsf91akKc7GOFlY1IYkF09kbiYXlnYvWXcosDRcZ0fbKDY
H72Q+ZYWwB/ZKMS1FuevWQH0SX1e1iBKaRrdBofFenHRHPmvSKQjEGdyZhUskOAD
AXYDJHNcH5pjEP4FayV226MdinHxSvIaSj6RKe9yZuCr4rHh6G+wl8mgue98N5IO
U1q0/k0+wMteMitJw4B8/Dj91ASL3bhhNKGGAMDickPEC5W69oXvAXOEpA/xVm0t
tcE8eztryH31dd+AksUOF8o6vsNtfWeU24wRP4Jvh4/5AZU6Yohz5XlQUdFHMsSB
6C8+CuSJkuT2Fbq2BC4/q4Lu9J+s9EI90rtbafb0yZZqniJkBaIfd2fs2ivEul3Y
GqvgNxPwfarBlJB1a0mR9bWbBgPVtj6BzosMgpIW5gAPYDR8YptHU9j7W5r7Hxsu
Icq3XOC/PVBBhxCWET3lLCpMWFjBOofXhXZUWH50jUXSpEJSMQxSRY7kILAkMIl0
oSb9sYxI3jeTj/FJliuG8sPCJ+dqNNjPluymYL7uCJUcUv8SNscgV26J8SizMyew
6yuNIUaJ+gI6ytcxMCWS6ZLPkvO28uSNZRgHqOmFRzNrnys/Bik/Q6dW8eGuM6fO
aFW2NHHiV1yVzGBsbdVPBsCULn69nJLYhL55QLYpT4XMdCncQduF9kr7CupsdhUy
3LPObp+x/FdCfX0dTC5IhCuMtBFArCd7fa7VvEM/DRj75QaZfYmnqfdaMolpe6im
bAC70GGq1byRGJCbomtu69D0DHu4zvAiAZYlzBMNpl4mKdawz+YAtzYfBgMrCCMz
JC58DoRo2Ckaz94wmdoCgxi4aC3ur8IHoM7ZnzAmE+XUl0IKm2vQ4cU35UY9b4oa
x82dvi9Mgnd4mS9ke2cliH7IG+qK0OKZOvXiS9BN9HrWVHr33O7yDQHQQT4zHu9b
FseBRP0EusZnNcdQ1yes320I+ozXiuJ9O1RvJeh4DWzKRiozNnAnlODV2R5Y8fiK
Lh/P3dbtmrZCKZ9E5fHRY93zqzd+kE43yr2hBKr7LHEHFAqlncifyqaScMj0myYX
/mWWBBLlSRgdopltlo7kxAjHLFrVGjvCd5SUIoV4ixM6DuG0a1ZNqbYCvVAqjdye
dCZBt1wR68vqOGJtnsDdfodLKwOk4GqdOP5o7UPBIAi5QOF3xOn1bDq0Y6STalrD
N+X/V9F8sEvKSqsb2Khrf00Tpxx9M2HzzvlXhFq1WPYuP6uJrCctNP9V6m6C/p2b
ynLIOg3RXAELLYQgTqvYU4b74O22KfpUxbxm3T5MGmXoCiZDUFhRWH72PT+ZB05N
avBD7bJZgdpHZvjmZL9eK21zBmCalL1radopGEHr8MPEnMmBJxQlPjsJIxCuXQUg
yH4qLOY4R1/UD/aKspYk9QX/kwelOboWiWE0j0a2NUTAzD5nTwaCD4bM7cbEkCjK
9qFg6a9n9ReMyy7v6aF3IFfhT9YlqkgaIzqB76+87F1SxvDUlMM3LArKjzKoLQAw
L9svWv9pRJfhQDEEyATBSSFoxLn/Yclg48WXM1bxatmA254SFHzE8igR7SLaUin/
3m8oEMW5XIgTSHkVdzgm0cGLjUrCN+gAZ880lDDrpNhcpnZvAJbDGgg5wCiJ1Izl
Ek9SRNGShYRbJuhvv60Vs0IYucim+sLgYALa8gaxzcFZLduk+dT0NvpkalvqFd3e
SR76BsptFvUIbFe/lNUApHkSBCSZ3K7z0nMuungKdafuE/TBcZ9sHekH9ZdqL1Gb
/TeE3xStbI9D1RqqBft2ZrB24Ahg5JBZEPHqeHwtVckOssI/RECAnr+QmPsGgpgd
PnYucpPN5T5vJQSBPOs6v1SqHHz9EobfgCpYCvoI2kOpgNfZqJ11pk+c+csQexZ9
G26CGFqgAYhboq2ukI9SA3rfwvPx7tITcWIBLRjzhLrcckkg6lLYNj5YJzIQwPVB
/3wqI3fwhst+114OPoqJWUtnnL6JdQp/PkUIN9nppWs5eVPpUsgaD74PqqOUOKia
fTxVsUKWl4EvrZfrwN0IJ+Xe3W0FRKv/EOxs+0JBUBMIkr3uV8wyh6hJQcoCOxnM
rhD7uACFhkylj7e1+O4OOf8jhHcA27CfX9d27sA6AVU+iaKdAm/qs18fSJnS91Iw
5qKiUULfIth5hdLUx8nXX0ywTFbCWKT+uGRbSvuZAbQIxDXmpCg+OLxMafgWtVtk
vbI4ByUHUhODa1RFE6/quklwiKzbdUY14NZfLnIccH7fBz2YMlwCoHAQ9rImzv8e
iSOnk4M4WMWaDRpFU5ks0Rgbik20qICexnEyL8mrO6XiusNTTeF5oTkjB+lIsaG4
qC3wDvjSqIonCZLvuhn7tQ1hCA1U8Xuk6Ds3aukgT3r7Ph/IAcnMVZmCcyLz9wzq
cpBPaviEPpt2t3XnfRv6kATu4v12BZs0YD/dJsciqcW+wHUQIKMd+FbXJBcayCo3
+if0n7RC3mAetajuqg0WCZF0HtocEFmPQt6rqqSeOu/CBCZ7m5jIjjMmf2mJfe7Z
M4wtaLLUDKgy8r/hv26M94hR7GADkD0AQNHZ6T3ycWOjT7T4lddAjp1OJQHcscqs
M8xYOX90XK/pELVwhINX8U+SaPtIiH1oK7yWUwyeLL2vfGtjbiysv2xcQLvsvgkA
1U/OiZ2ORsD7wYKrg/gJf7kjKCFV1wUAzAK4mpbjWLKli3obL035betsEGQWtyq6
55zuD8S2scbIZ5cv22BtHcQg1446Ud8HPrvOyfyehM6Y7Q+fBWF/Qpb8dGKj6skU
345EKITge9++V5wRMwbsK+gfKDMRXFuHPmrTaSDLQxj7Vhsq+hFojI/esAbz2tWl
VopvvrGAetJzeg4YV0fMZ75htedAdPkELLmBGGs9YritMF/yiAQbLPV8oIKCbjFr
oPUdS4QTBPVu0+KOr0BRDS1M6XI8p3o/aLhgkPYygNnij4nlGZ26E6miIzREj4Os
k/YLZB87GjgQ6hl4hg4Xp//A0str2RG3L7gzlUzivE7ZXz7MZCFBvKNHm4LXF4CS
WW3KrOAjherOJ8DZMWcNrUnwaVVWFj6Gn10dWBeEeCMidu6WOR26zXaeEGFPhJda
vliT/AYilNe4mv+5rcBPtoZzbX/EZx8Ut1+EwJQQEpt3ilq2Ci3pfUsSutsb8mmo
jSf5Bzd29ESDLDvDQnpRc35otwyWYNzOpGI0fkbNF5BLzBwPjitkONtI0Wzwy94g
bbvq/Rh/XDepqhiFMEkiD/KyZ4fWbSrXrKToyK3otECymGjOpygoq1W0ZB/o09/f
PxPkJuKvHcRPz12CBhfN8Q17kDRQqX/1EnJdtIlpOg+eJ/GIoY0Zk3C8T2JYvkSh
iNv0k/PeBjVbTbkiGLk2ecf+cgNKgl+1In9jZ67sAR5jOuLq3deqnfB5y6UiwK7K
F87Ff5ao1Bw1CbkQicYpKY83DrvpcEHkGgwB8QGfcgkFG0iMG2PbLRmw+OseKrB5
evAqP1q57+d+rZYErmoJJrwIBqbX2RstNRqJMbgCPtI3y+1MBmWh2cKgLaGz3MDl
wuA7FXW0ZV1d0uqbxhvHN714LGETtbkRt6ZOj1NGJ80SHpWcfo9vAcZaBP3QhZHM
1GIIaFUF/r6ZISiLwouTDpZSHKzR9OoG59TFotEMxinHW3VO4+lfJ7LmJDSbUZYo
N25Xa2ElO6QPbXNYp2XqXcX3thxTNTV14J14/xpotATWpwhnp4M3jBEX96T4IxJR
WemzA9V8XpH3ldvsfQVjtSNlvyBU/wMKM/JPsjf6i4VoBwFmAxr6jl6ekMwWj9ny
Ypvy4BvUOCjJKARmFA9XmYyDTsGtURCamvTOHDpcWPIGweG8HOtDqmdNLW5D2sLw
n9vcJ818aAoAtTVSIrQBEISo3vVmnZ71hhiUoEm3uS8+3p38XLmPfZUGf+24/uhW
dM1sLJDM77X70xz7qJE/cqQ64WhVWurtYmVtMdZUwJhv+R6+Ek+phz3pUkrHiWYy
+qdhUPFCdy/g83Lwqitrh2WSM/hQ/Zpu83rlAVVTAKDRgUmcMSgguM1Gu7m+HuqI
EbwhCr7NxoThvCePfjeVKjjdf8xzrX73hvL3+vkfco0kfbsXsRYwnL3+721lCV8x
1MDGTb4yyENHHVfLd7aKC8NB8iPVby7COcNa13b7xW1J0bQszpFJTPK8I+fDycLq
WIyiF4GD3IGif4hfzgtH4hG+dsuzvARVfHm7/sx8fCaK9ksvqV87tDbA3fNW/z5S
7nIaKXJ5MRIE7XrNfvsPzI08KEHdJwqSv4eCy2v2or5ivNLcF5Ksusdqnk2AFL1c
gEquUnkg8vtzznE8TuAbLHYEw4eGVxEU4/rjvTsLpye4fxc9fnnkWtgna13CM9m3
y3wdLU22yWOchiGdgW6xArfOeJVHsjeFhAqPn1AVhSJV/rAVjt+Cc0/YEDMvxabo
MuyoJjK0yVkM3YuBm7PJm5ObBOjxBIMu20Y33gMjRHiZTNrulyFhsGHt1HLEGMnI
Fr820NotS77RkDiSzWnyRCyFxtzLS2SbbIgGQI0M7okh9J1aYdDTga+0+bVnXPxy
1Rl9bQY2I4IVbufe+BPX/6UWYPWh4w/3JQasY64XAOuNGqt2YV3/oBfjJ04s9P0k
/0iP0aHwRHW3G+kTqaIuKLUuQEqDntJrIP+NFHiHZo7W9EXPI+37cxp6DkHwbat1
XM81K4VuO/V//VqVIoU2MvOiG+hxDTBOBZ0VpVKHd/Zlk2WXOT7W7RofJ+KvIA4Q
9SnGaem959AERfZBj2owSdYwEBs/IYE7WTPvxiekKxTM3AEVoYIAUM9nR1u6NiXl
AlAoZAgXncle23g/KE0Hnx1+ktVkkyWv7zGj0wVkekEz5t3HfGve1i1G0W/3IaWD
wnueXy3d2wl3tI9OPV8TNo4512QL6MhWbfyZawxvd34S5zyrYh4OGoGRs/Ld/R/v
G1VQLCmWYBpIZdpWevRjCSmdzFiWhNOdxey2Y47iDiAl6a9wH7P25Aq5Jun6YelR
Za53nLrBI34IbJ5PakX9qxjtYxRoGcukMAbAv0UAgS/Ta7bw4Mh+S2fQUZTpMx+k
p2ueeulV1rVBUxRwu6LCmbypwXxUEW2JLJDjhlk74WA95Ni+d+5oKYiy3FQJp9zf
pDWfXv71Ukt8oBcgVH1jE8rIQRL0VBq2uuKWOHGSlycWggEPS/7hJdFyUp3dzQ+U
tY1oCampVA34lKjz4iqfCfcTalKQ2SQ3TvoUc+sYKUkwgtp6esA/5NYOaP+oW/Gk
cGbWtX9JyS8vA8UH0apzxL3ie9F/WxiLLnMRfWvQfBdOMWTjpibWvMBlPhaCRKhM
4HG8MDiZsn8Aho50N1UTy+Oeltq3cstsSzuYWh/4ZzlW5il8mbkLQHTW71F6917D
6/UnTpzoXM5yTVQ3K6vvhn2Ts87jCCz0Dmnyf8SVbXgMIRLS8gtWQcy5RjUM1B/l
7gfQqgIUOBXhDAIVXr0SD96pTk8hAbPJ+rqivmCU8/QnSdt2AeZ7djinAGcFGjEc
V7qnody3npVH257VHYCM161rtls1pjllTKTSvISnGDWvrpGdHXiF9orl3/zUccRB
jRoQcaZZ1FL1kBs4a2qx2pKSUzZ5868uZEeqY0XNuZgWStB5x8oM1xQ9p01kqEXX
E/ZOua0jxCyMMZHDes6xHxRpjXWWJ3BjYrjKo3kiuqjML1s0q7i8v8h9VUiB4QZv
zxgWO9j2hJFibdNF23CYss65Foe75xGOzTm4JY/GGgFtT0wPUPrq/+tVmMH5tD8O
WlqKMKhd3CxteQsKwkJwOY5HpoCBvMNQByf61GPZ7nNO151j91xbD1lenDO1OA8E
rpx//vnVWSiBb8HXTr51d0g1SpuQvTbMERm5ydsInKsCXse1t8W5j4LOuhv0iwTN
aHyeQjAc3UnBkHJKBnNO6NKcJCx1+DDQiVXgMWSH+ceHdpzS2Aa6mHMzLb5Z4ney
+OCIU24qw+L4NeCMwhMO0NCP2i3YjbJK1JrrtzqGvix6a3xJmkDvTnunVAPFJ0xY
dkKm6zwiqFF4rzX/+hJLpBbTxpSEfoKXHPGcptaqSPP/Tz+qy/C7Ho/Cocu5xFsa
/ZSgMKM/kpb1GTgDYaa0RoqxbHET632clQigNVLtFc2pGIf/eN5M58I22sY0vdwK
bJ8Pz62+0iNjFyMH/wiPO8G6ZwmpQ8KvhV+JCPjYIXW3h57VY9CZ6g086mecOiEM
Hfq8PBWgjwSqGhkTRvlOkL67jAsSLMFah3jypqUiOsr2lQYWov77tMwJE7P7/dUC
diji0dClEqrkmArFSzhnlbV1XFbwJaQ5IKf1zHvi+adoRO33bF0eWMLKzxa6LQmV
pwG/C/PgcvLJEaca0hJVR5tnE+j5EbdBZ0BAyATuhxLhhnNcGrQXBIm8lRi0gZCm
YGEX6i4dihq3zWHsahPDLwlFcdm1bSWS8VxC+4tbu57+VVjIHfTU9Y3tgj8Ubpzz
sOdl3H4CKcwxhjn0tqZLVxhWsdF1VBS8ufTpVNxM/SuCBnGi1cvEP1hBtuYvh/xD
DeZO9wMC4Gt00E5Ey0/vUazM2IjvDQQCPDvc7GvQh29MeQfNjrTy1OP1+z8bzcs6
KhdNgWAWzt1anmwuA+UeFFs46Lwva2XjTVsC7hw10EHUffeEuDxscGUjQhkMVmtu
2AAs6tFD7e1Zn5BDophOei4h5aHGmo1FFUJw7gdlRQrxYpCdbtxmLF2i9gw98K9F
tprp/kwK9FEp/yp81Dkx0ROyme+mHlxFnhNypUY9TYSzZwsTLv2g7LlHWNFXrV+n
Q1fDJsycYuVFXAmql2BXBnxtSqqxqC7AXor0xt+wwDDKhYN/r0wpJ6s1OuUpmW2c
dQqZkaiw+zssVIDlpdLBGN7Sepy80cNUANkV+2jNRScKIHSm5HWL/kW/gJ7CDZx+
cdDuKDEI6mL0ljU4Mu6dd9NMfWQexkxiUi/1BXSGaQrTs9Pxdvdu4DzgNFpWuL24
Klnx/IIgFRwy7wIPLcBcu6bjThqijrTg1hNPhMfhSec5H2XRT7GgU6TQZ/3HT0BC
LnU3LUMaF7xUjISDKqNPXj8u9d/uw1LqrIk4RZ9ayBujfvt5gddjT9TbQ5wUNEF5
bDhGe32Aoqsg6IfmWPYi5+1SXE+9UjekN/i6H7PPxVHojsjGA2pXtoa6FnoZwKec
Kbx2AAhGaJvp0JrPnga3UjYlWalI1Y4jWdGVqMBguC7b6lCO5419zaqtk+ZFC7Q5
3TAKytpiQuuOccX6VP4AhVyPO3tU8LEqr5JoAmaMy2whP2kfMcn3bOoXKnERe+MS
SPh/X9hGNi2R8UfhZGS7S83VocUICUpy8++9en6hn6b7/RjQibE02lOd6qFxyNdL
xOl5vhyHw+IU+ySL9msP2L8KtoRpjRh13EogNwPLGrqIrrp5aqX3BRT8ZrCdMKwM
5gvgj1MX2kJIubDO6wOnqfLysGFu9GTjpDDZwMQY12RafRX2giGYpxA9v+N7ZDhR
uxnG2ivqcliWP2Bl0vpHge42H0idFUQYdbesxAnusH7V6FdKC9HxcaRKcd140hqC
BanLlfdZD7FilnP/4EsLYB6TQ9gAaFRXM1itq3zRTFNMjFyxTO906fvL3/tV31XX
loYj3+8ka99DmroycAENZQFpezcRitQm/67ZKU15I35/kWNl8qLbBOTqpUs7hMxz
YsS5OjroW3pPXcIHrnlZsV8+YZWAOlqpNvX1gA18KGwQgwdQmykT6UFD5NprXczS
OwsbEn6i4J9M5r+49EY6kD8EXS3PAOUlkwkI5RV0xHYn85AEcggnLJ2nIL67soC3
nRzmh+P+Gmlnl9DKsHC93pOfAKiEMyuHQKFghKwQ/iQPNX29wKKO5cjStkySXaKb
NalWmV+G4FTkAIYV/EgjHgXH5SJSyAB/Mmn7bl4GX+QImsizXNKVUamuPb5HlD8P
JbugEOVrah4qhkgcM4eVJn9tBKjpTFfyDA9OAOiGLK8yFC+b8OzoHj0eXHodglYZ
hUD32eBsDVGtDxqTKigxVM8WsAZ6PXiGeiV7BddTJwG9TT5+SiZeHymHmbfZE26d
4fEZRaSWdwaNzb/wj/LyThrT3IIZffeg/Yn4yiY6b5+tPvuhMor4LBn53CT/mYI4
aTq2w6sWldFn0YNoIAeAzM+9ubmzEC0kG7N8j4HrdWYdcD9Pank2GZR7Z2diyLGF
/0lWXGdqCfi7RwP+KhWv73EFSJ/OJ3NCPVO44KtqC0nSsiDbLwFVvZCTOrKuAP9+
Aw2SmY/iVLC2jvrHxqJudN2kdMsryi4vIl7I03yPuONUk54uKT2WiktaiqCzwoqU
NP+1AhUKjVD6CcelnTtezTG86y1VmOI9bS2ad75RV7etYI1vK/Sg/mElMUvUp5qu
ZeKRRrV+yA/zhMyCMf7d3HKquiLASmEf4pS/5P/DP/RhkO0HWyMBa3zohxifQl+/
xnbAKlGYkBBigI7+/t1ivE2e08JObrQKMZuqFUWqWOqy9A3OUZ505JnrHUSfEY8r
w1PNJfsRJ9ET/qT6s+6+evLMT81JusN+3da9tmvPR23ja4pRXhFk4oc+gQR4pw4B
2YOX4CUCnIh0VY66FuZ9h+95Lq15PQfBWeDCxBzZUosfsFGLAPdAPNgKPLqqPQXp
mf2Fp69WdyQq+NE7dbbyvIXplvwNqYGGMw/YBTD6YxeuUF5XL2GNW0lR8aGZOd3k
+4VHk07njVmO19Qf/Rr1BxI+DJq5lIqdL9fKo6209BBVFtkDBliMNgGuTafy6Y1w
uFeM51cRsD9RKNgoKJfTwJsPJzd4gvGo0+5/5WW6NfCdx0DyAKxW6l+EqDoucYE5
G2/nxHGQQCeFdqSmmeqI7EYK5ZGN2t8CVLZ6xLpVBwP6hz+a28WNZ/Yur1Tg5FDX
Xy6QwktmNEiLjX9CGaMbyKJHK2vOha6TEHGMiIVNC5arNJhQrC+ikNmnNlx6dZCZ
K7tuMsTUmYKgOMY5tmDFkCHwU+kDnqCXbZeMoV6IqtSad7dMRft/iDYaR6lh1Fkk
reS3hC0npyJlE6QFnVfmgw/SGDzcAgMykl7WiPovScp75kZpW8ULRikFkQxW2r8S
Lqu8oPZWFrW4lDz+XBVe09Co8pxoQKB74hbtyv0c8WE5EXw7LUUoqdQsdPVrKGBt
ecSp3ytcLCgOv5L4cqlzjM772TDgXFDABfhfN6xiJFkijDhxeejpKIz4v7zPbCQd
Cu7zzrI0wLsm7b3SzjR5SQWQMiGoaq0NohbqpOTpzKLVGOqvT+rCv2lHBmFnLTKm
utWN7fg73cWcalm7SqggsQMRP0x+PAmmWPjokhRcSquMOGHcMor67bQFUfm77XhO
8jpvbx3yOHgAng8ahgnzs9YH7JF5jveppYK1De4zWqyeNeye/m6XdxGDj0lzvS9K
xbzaFXcDjabISLNABc8OU6C1sjq0Zvu1lx0ald4Tlywkt9e9HKoKDfN9tmu/HQFj
j08iERaW0rV0n/O0F9QTR9/HtS4PcXANPd6BKJcxY8zxyer21zAg79UuVaEnk37t
7Xc/1Iv4H6Ao3oaeWENTry4g1sjIthtE4MHxr9ibTBtmiv9L0MO17E9hIIfgHVVT
4TgGdu9zRfV+/8+7QbAyRJtDmoXc7AM41b5UbD30lLpPQ3QxCGEdtdMmRlHpW8k1
BcPEETyYpacuOFdSGHaV4/GYOJOIcrX9WP+xII12yXCmBRuf/HGLUfZzIo8Lmmmr
Je8o3cuv72xLAaZdh2LhsZsb5mT1oLRzgy/4LC1ZpTjPAs21E/WBwBcg4VOQbK8n
iKvLAi3205gySqd4lCabeWgOxmXzSMSTl88vT+e2xLVw6YBK/nfrp2gwYFT8F/Gf
cUnOlhcGp1IA/QyAYgCAwXtspyuAEs3lI2GtZTkVKClC995RJ+DkayKtQHis6fmZ
yjGavmpURee/JP3922mmo3M10xlJnfEUg7pTmIGjaOGdO8btOojyo/l5k2AAcDus
Cv+5wf98E1j798dH4f8u6nFhnn3iDSYe0aEtOa/+Dktvhgzwl0VCqxYSceLFei8Y
7cX+v6Z2ROt1K3/QRicDrB5MqKnveb4VL0Qc8LawSYk0sZzIeg0hHy/fRG6CvszZ
oIE6+9HD9LtOgTZXCw6Ebsb5MIYkt6aBBDKOErOyiEHLEsofzBPNsrnwLH/BovdT
F0VkphnM9hpNzcI7xYGJzbAssj+fvQ4elA8+Ottx7huSsBwV/z2OnEARISo3u9Zo
UZ8jAUTeWGReyHIFleBSL/7Mi96qwjlfA+R+H/gXR3Y/0P6zdqR8H/4+cUYx6Pwp
GIXkafl4Pgy46XyQQVfRcLIHdgCfJ8qrzTPfxX79BVAZuv2cd/SoiTejhiPyJQF2
nzufP1BuZ3lKDptRQdNF3PBkP9N57mS36PaLvprtE8Az0dMksySds2JDfhcw4/KX
zUGml+smr80RyaAl4uV4M/DSfdYkTogY1nHKs18MRPk3orE5CURGFikMove+9uxQ
dbcOufsEqmq/2PLOaMTzxsnjevd6Oa6vgiovjULuz+NDjryccHgQl0YyLe1Z+7Mt
VAYfxhCJDg3LpPQEqWa7agtJntIyS0nAyKNvPrNNVyrrLS/bzYLIbbJNi3JB5xZ2
/RipGogzf4Wvtjc8Ct+SrVNUykavM4PaKlq6J5/XrPZGNpQusD7BJNziyq9G+0ZH
B0Yw5GMbCvPIjnK292dRCePp1YmEPB9wd0ZPiq9M4tJLJUXpjp6cQWepuMrv1bDH
g6kzSvJ0DR0NzBqC6aTcHwSS+IYErbxZxzv3Rj8sIb8LxOUKZviWinTkoH/F0TBX
lVbuT7HRjhwqqYHZzfgX9Ck5lF+Sq9tMwfF5fCmiqQXoYesiiG5rzoP9srzUqyRL
+ebhXNJrX+AHy/b5lj7iYvzlJ3HTb4L/KHj5l0BOsgX1u2Tpqrok/FfHL+svqxAF
yx2kAGO19gjFjrqOiqrk+JU2LBQuZutA6OGf56vqd3O/J9L8tzpS0lSx+EUwK4EF
kSX5dchIf5KRH7tr/cQ31llGFPgiXvORfutneho/QClv9WKjHcCXxIjUz6MBfzTt
hGo/e4BA9VnnnWstjyDHJ82yKcC6OGvGU5JFy/9tHseaAkIKyRpGxgpwTnwNjr3G
6f/dwP2/l2ZICQfinwToO7fNjR5BbvK/dm1RDglgt4ba+5BynT44EorS7r7HJLm8
Fx1x6wk+EgE8k13bqoW5nVGIqGHLalSCKYUCbWNCeSJBvjKVsTdTaqdecyqxqwek
5zesXIMINTFNz/wtWE4MAxadQ55t73+W2Pa7m+uyFx9jqLXxHBAl5GGAxxO7ce3/
tmEhNxJSq44fr1xqkPOlgqShcF7vt6z2YzKoebrl6U8F9SVPmVZ+gnHIpeMKUoai
5JYCOC1F9g2QzC31n/1LnyuWE6S3308HZ1nHjdCzvxI99qoFz03gcrvARQO0ID5X
nUjdAMcNOMKNxZt69n1fYtmLzNOWYfZxTr6SRt4vDfiOFTKZCZE8WQ1Qvb7yruHS
7IZet9a/ygWuNEwSaN4z7Pf+L7h/quAtUyjA1CQigSdUyyFLiYkVtYDWdEflVrWT
F1JmwgoXTETf5+6tO2vZFKL933moQhP1Vi1ItoNPGs+Wfckbh+W//4ller8f4uNE
60RV1KYYmgBuXxovrC+nYZ76LO7fODhexDs3IIRJqahsV/fL+SNf1cwZB2x5XtWy
GwncvH2c+/shj7Be7kxzHeq41R/w8REpS8Ea7sDCarWkO/znuSymcPHmwyuWtiJf
EDHU/kjt0y3XsNNnr+i9WmeJM5eBT9WQ4Y5uI4/MSths5zlFPFRRralMn3umpJ5J
X9EKyXCeFFn4cZJyGfSEPCFKdikHunCwBp6KFq0sTsPTaymp6t6gkSOktoMTNpHe
Qsw/6bSrI02P9FqXXHKbRUJ6QEatp1Lm3ahVXRLW+UwG+D+J73KigSnqr7Q5UbIl
XrgDseGMVDqd8EtFKWUFg/1Yq1yJWBabXpXsumWECdzNTQ6n8lrQsDTS4chOtikS
vc93dtfvaXxoumJafwFh/YCqnYRH7fyz3WWkdT7Fg4u8vNKXekKFXedLxu7UWoj0
/O2qle7dc1FHQtpTTGkSJAX9m20UJCeh1t8bR+hGTNOSpEduhBjl3vtBjPQyIy67
njb8PwjlKSCO7McXfe57i1QnZzpGqekIfJhV0jaJWGdc+ySWiIGRaTuDmOAtuhmT
UbAnXkY3GiHDPhAsvYsQmyHpDnYGmIvnPRJ7WC4VMZZr/YlusU8bJixXwGO+SuiI
y2HprY1SL63h65JiIEvDatupaqa04ghDXB3cGS1tIL4vWuds8XfgVZ5rJ/9x2D1X
U77qQLX7Ymh2SCPc2D/nBSj1urWlBd0MhXeICOo0kt4PnPbO3CDRheokh5BrNZuh
F/AN8ajim5jrthPoA7g6LJT/hlcMx4+J923RZ5Q9CNB7mXzJAvzsmlDqpVELX0m5
A+SwaFTWOZBl4BX0/RKdQ6ybZHpw11jrzCLWO10LTFibEU3ylzJuu5BYg5K46fRg
xA0vX4llga6Jh6BO1se0cpTTy11r7nHiqQ8CCtozkk126a1grRXuL/cxi1VVoj/Z
51jpF0yI5fDu3MGryBrUzZZ1Q9o2leBOhFeZtbLAcAG0o0fjj0KD7AtYSj0IMpW5
9RB9WtLyKo2XS2HD7i18d5doKnjRJeTTTz6j+11ZcTE4kSPg/yzTHVHDJq2WhDXU
QX91zgbvQkasfQY4LIyKZp3QCPAebIqLHqLU0ZQWgCq9klgb0dPxMMOV68g8yFDD
y2kYw0i49MeA55btlQ6/BGkWVhKo0glyXYgENi9B74mCUv0ZPKNu1xPUHxlw76AC
XV3+Zu3zjb1YYRMDSSvJVB+Es4h3uLPkISW6QiQ7r0NwxKTbv+qimLCtNrwE1yYi
swO70p2Aa87ReZGwcZ4U5O1Fl1GeETJRU8PMio+A6WXbJhLWw+CyVT38WSXYn7mR
jU3TbCRCaSoXQ08wKnTyD+0DhY63USWDLLhzGr46jvRE1LgtYAB0bXi3lC4wIpTf
KrRvrpEenBS4XtSAvVdIiTzqRyVAHeGam4AsQqyJNCgTQ9jmVUtsNIa85ni7LD8I
UoVq1luIdfVWdz/qA6zdsw50JMG8UPcZod2Tp1lvXXfJ8MqMVKTSIegVqFhsfLbG
K6Xdbp+xa6KQGB0dPyOEaUn63z9AzW4Bvgx8f3r6Tv7ImjeTJzFLNf7W1ccOgOt3
eerkuK4HEwo9yPBT8Wacb2LKUb3VRI4TZK1atk7klgluBY0HE17b4uUhooc2/6uT
TWDvvhVT7cHa0zcQHF+c+oiMY0Kb3Vustu8DaJ87aNX4oa7VhEbmDRWQQi9Ve3P6
7Upg9Pr/CVmfGwCwCG1i52VOqBDrjGmxUZhqXqpPrMqiC0FIZ+AYrZM7fMi6ULM5
SMMG7ZTvTwNXyyREUbAjnZVT05ZO6ED5Yl4ho5Hxu+tCx6xA3gEGlqWapTQDav+F
bYl9vnDj544T2NB8tKA+ACwsViPaWm3Pk5GTNCjL2THswep32R4G8OTWACH4ZCu7
/n3qhbUHGYlsKHRAqx29HDtuNUZrJFvZRNIhyrAxPFx2YT+N1QQ8r/HFWtQQ5b2g
p/wiif+PruP4kbXdlSdaehtS2zZw8NdVoE8ph1IaCQniw0UaFXXGpPnzzf/AvpPT
uwimlGQCf4MP2AnjIVWR2hwMS+4eJfJ6MB8wPGBYggQpPT1VFuvlOZ9e13T41AKg
8/rFtCcYdKOxWapEjjdXzmRUpv+HU+MXOQujwUWNhK7DCtCyuexltJsMWD6KDmh9
f3B/IdMv3jIk37Oh4bovVAUgnyaM59Bzj5OjRwb/JBDUJvPWPBYqJ763V+UZz0BT
e0Vmew93H9R4wvU4UJZoL0gJwdJhZStfrb/sXHCNkq14IBUPq22QN4DamGzJYdRS
4cDVV0hYjiPc+tyrnbYK8NOKnwYqfyZEWWJFmKJDkB+ADvLdtqYR1D8rb/4wJc91
1UH/69kH51Zwl2vjbHJ5J9sSCYfQQj1HnZyCltY1FP7maV2ZqFDZGN8jNBokQ9ia
fyrWoVWEi1toysyxwkSGC11D8i0Hgt/BDFe0nOvnvbgKKUxCostfwg3VLySw4AyO
LXuiAPQs9M24sw6pEKs3HH2lza5xVYCTic+pJ4h3zTbAZx8K91a4XXljhgYX7vZM
oWCWuuzY5bj4q/ocEYmVQaT4ESqJQZP5s/7vbybpAMdJrjouw/+UMccIrC5yGXRT
QiigzId/5IQhj0lnwqlxM0SjfToZOyFmbG3qZ1blHZgJgge8U0RRDA5hVHTBeNWn
AQh+FBR5eI6gaRsa9hM3Sf1UsHtqXZ/HbaIDY92Cp1/Q1FJWFC43xLKEr0yjvkwB
kdUq/Olcf4z8Vmigb9SboDBRTMLvIczU1jh5dljh7YxcF1cyiaUa8hIXxwxplQB+
1CIGE+ufM8fYzbwgxoMQ3lsQTK2n4T0ACFdBXKF95eRrGD17Qj2H56/QOFfI89N6
ddNVi8ggBnaG1n4YrS1t6utE7V6VDHTzgrffeMkncDOoU88qaeSWEqDORaiLHTm3
39DkL5jPJ0HDMgCUIADm69aXlbczfYKGElQAPg7hdEiJ7JDwSBNFujdaQprT9DGO
SeOReRpTFs+xOt43X6nBrur975m2rOC79TCthpcctxiz9aGEYA7FJANnBORUdie6
4e8YXmtXkGpjPsaLxqdWPGxdxEbDxUuYDQjiL0ZCoAe1gqCEBbaBl/R4bZuHJW36
hgxLsKYuZbI973onwjzDoOw8VZLN3c8PziPKaFZL8j2a6XySQxO9Y6PcTnqndPmA
6qpcQgTQ9E9Hs4mlGP4i2l0HYT9x2I3td7TioX+jo2/W6//JM2/Jixxki17YL1Ic
MkuShYpL1CWt4L/0F3ZgyWxwjO1fKKoXC+oC/hiWHFbwynA37HwteMJyyJf/trOz
8nDs3C8MbZVXjyKNbES36lmIuB4g/rvZ3mjdMqFsGvUjHvIV9mBosvDpw/BtVm87
aURpiIgELVobS8TvUscfcGcVoSxNscgfWOgD88ds/WKmR5GZQmjjxPRyKqWghRFa
zIErWsSl/B+2FDzzJKM1DFjd7JqENrBoVyhBk5hnUdGOaD6g3zo8hyVxxDOdluqN
/bxn84ou7bpkXah2mFjm5f9LEFIhV6CXU4iRX4LDN4s98WtaDwNusdT6g2rSFQan
Eiq05jOZBDGcrcdQURQsrGtBBakobCrboHK4FoCWxRC8IDttcbFGSfHlvU4pa4+2
AL59dD8Y8ZHIab0f05OoZTg+Ia7Y2yNFd4KfFCsmADOfP4CnCkbu6PHKU78jEjwY
oEa2obEURcBW6LhUHDa+1keE3PpzRg/00jrDKyi2f2cvSllkRaPrS1wUnItkSBGt
W98bpnl8hAhMxR/cxBK/UK26L8ImR0nMNoAMdZu3Nz4cmRyD0OzJkJntXJtDXNqa
SNGBSpnaZeHSRVI5Ez0TfAMq3x3WtmeQASOPamAYzGWzTIAeoLKS7z0MdjnHBb0q
3A2sx122whWPWW1P59+BoelZtkQlk1iiOZqppcuIZR3eGufAD93TwOw9+uUkJzUw
NCE5xgpj6kfXLzDA83NqCzqvc7t3+Yec/9tQyxDkM8H9SW7E9tzSRL+iTKMmMADf
Oo0v4J9ATxaQZGRY9GADjWHNOKdM4dphPAXC5A/HNC/LxGatNbU18HjEw/PgySO+
Sdyc50ZKXPn1coAMOdu2MjGiZ/V7ZfqZPoVBNBFHc3fvxnmjT6CcyzRtb70Z1X2I
Q7D5OzQVMOOIoanIacbqwdwoxEOWuL5ObPkdhb9ix4af4On9C4IyZJ0YK6whBiQW
e8QJp9+FPOjqyquN/d63KzBRjf6/h/3a1oxQ4oxbsdDMfuqiVKj+/MwVlaJSEu1L
fVlDaHzjrA56yycT+jrMv3OPEuD1Cbzx5xwNOUZq+DhggYYtTvY69o3hLl4CRmVl
aKzc8AiCksN/Yt0XJyOSobs7duZdeiwhd3hNZl2BiALTEVxOo1Gjp1+vwphVe5M9
P5kvkAoZWOjfNsyJ/K8Eh1BcNfc4EEGmvDqlnWzXCYlcYN1/fNLf6GzKbLHHTm5N
aNuWUs4qxaQyLCMnyLYaC50UuCo2ajTy2r74pcXb//KM6p4pkMNzGQlBrqSo4ICq
nyS7s1pEPuWjFxAc8on6xS9jnwOSjd7R1gEPH1Aogdan+1D+1vfwm91uWuFPWH1S
Aw649chJXzu0pQ+0GH4y0d4gzwY1s7+wUIDYP8KEhulW7MDkg/xubp+21AxFBTqb
q1fAeHlEdvo1//abEbyFYFoBKyXADrQR2FQ+lFPW2ZagxhwQEwDtdbuBRMuj7Joh
mrfuBDAQxuuOcGxSe3XV3cB4VUDgXlluXviFRr9QT/3u7laRHlGdsMO3mrplDC4H
2d8IxaYaE48LtKuw6eG7pJ7hMomBtoGKrhWT56PjFX4CY2cOOsWra+0MqZApVbXX
PcupXW4ykKYhnJak6LPAigfpzeNKmq+gBulbQcTBDcSCIMiSyqVycp9E/0ML4swE
vQtk8oto7c8S4mfBl500zpND0QFNcVHRgQ+1hs+1YCi6MWkcUtELAR0yCWPjHGXc
dFcvpie87C67yBe1+6kj/tNmNA1+qn2p0H1lG0i7pJb1qnVQYVrjkiK9dR/K6qWV
Fz1fhhz43yi4co06dPaN7GqG87iN6j2W3JtwzXjPinetw9dH1UM6SeYnjvYnI3oY
qw0bJJA7q/DEUdg9jXmdN0/Jhi/eymo0Qqk8UiX2aJDa1lKSQpNabuHwz2n59lFa
DkqA8mLAAHfGnxP+pw6hZCvR0OjwMquzhgogGwKhmB1AmThtIkVS/rhcHKQgncPl
lgilRHotB59l5Wh4yaCb/d51QdYS4MI7MxwxBemSWyq5L/j+O92LEV9c1PmrhGtq
3HsKv0nHoinRLJNMhOeOcpAGX94/2OXC5sTnk+qNivqV82xuYt0sEw4mPgfp6LlL
JHiBTUbYf9YAO8CFcNQCvZQpjQW46m2R9Bj4/Fyp4nVscVbQZLsjUMUCp3m27lOb
kx1nIKM10HF05kNb2wqZWB+B8AX11OC72ZMSpd9w13TOMfqqh4A3HOx/a4g5ssYF
9+cjwM2M5aa/SSnYLotjZd2HPoZZxsn9PW9zL/fT348DtJNEdxLEWJK/2JRHiWIj
SEdT8QobLJ1LPFG4eRRU+TxcLb8NDtkWgFelWPZG5Pp4gvXqPqPz4QFvJi9vPzs3
OG5XWZKPZmbkt/VtxA5WxbqvVsNGXYGRZrwJnvsfcSrud+dvNqAJZqX+kmMyUT3R
pw3xAvdovJB4OFVgwd3ipTcPcsbZks2QuwI8bRoItZnJ8DFZ5jcOopwsmzwMNkP8
4igdNKl5HWWjfJazhdQbmvQZ7tdRFK5HeJ55yc3lCbSTXbge3bsUYaCH3SBzHcz4
1PHwI4pC20hDiK0s8RvjBuyZcrgZp6N9QIKckS+X4yPPfTL1oAFCXsvSdZeI8Gay
9Pn2z+KP/oJbd+fsJNDs85veGe+lVo3qJT0WMuqM/lYEO6Zx32mkZ+cxglSuYm/R
wVUXcSfSuKxoz8L4UhBXfK0mBxRoUUYZ+Nh/K7eiKHM4phMs2DTl6cad6CLyLtF2
mQeAHri9PsmLvpAiA+S9+/ggrHQxhaW/Kls8hjHDlpKICoduqrqH4bKQWmWW/ccC
6OzoMa+x1RhyirnppfJDQh2xAcxJIgtSvwo4WM8+RpHf0ubCPAF4oVlzwU40Hohc
EkWEhl2hHJVnuyNNlKNkUqN6lufchqrdM28W4SWr4wVkCKl6kuOAYWq1LxRd5VoR
5jcxHMaiQ/3ajSlFIOfpS1eByhl+WucP5kdT4StrdY3qtlnFkT70beesXo8IAbA8
dCDg85FI6iUZgz7etLvEsKbnDysSYQD+ySGbR2UjN6UEy2DekfGd65vs1tRT2foL
FG9g1m8KI62Y+nDVfaWTOIVm/cUUslafVYBX3oiW6szDXzKVUSWBiv9WwBLtv8BU
jCcKTeZQ9DVxoJoGsOYRyyKSgpHOpuSHDiDRMHLXkxUIIysiqv4woaFGuoo4YIjL
Ci+DNkuCD+JOABXTaAcjMWvg0rEtmLpJHEKY6UdY8OJSG3xur8lg4kjtYJ4brYeQ
VV8mP2sRi2fXNuTdvR+wKbxGgKKIg3/WROSKXQLySYuDCq/BfyDa0wZN9i6Aclcx
jJfvP5BtIpDG4oO/BnCn24slOZPIfdjy+eCt7jW/c4dha8vfdVwUBODLh22Qz96K
k7sFNzIdg/WLGNcfMQxjjtsaaAR0qOvnXLyfCMJe5B+potmQeWUHMFEwboG1NMvh
DeRt80QY4AMrepUc/eWnB5IyXsngH+9KPxSgwYPwX3Pol0LZJmgVgthuLodFbSf5
2h2rdUJuAfg/+RZePN6OtnhNJ4ss/+2UVymDMoqtngv+KCmyvIRzJvH/or7fzhTp
shxN/ywZAxnxtoqSem7a3dCJSvYlWMZvrcn/RZokIXdVSDP4cZ6a5IrNGffOIsNL
K679LCqbmzdaYuRoY4/9XzV7nmv768MyHOs9KAEycsZRttLvSrsMHVfQndAmWu+N
M/MdwK0/MFYZ5Qp2jcxUk/S/VNBDmeGi6BUXTySgMa6i6BagDINEfFLCIxncLpjM
8msWyPWqfqXNYwarYwN81Ad9SBUMgfSftFwlPSuAGtyH4xxDOp7CO4Bj6amLWdWn
HOCUBce3qUSb9ZEurFuu9eTq8jnat6i0LIM8JdGcYinqtxcWklUuFP5w2o15DT57
FIJh4Nc9P9b7619VQeYdJ9R9Wou7/ElEImJM9DVJAG8ec/bvMJSP2WL4VxPmjxIU
PwGFE0xB/0QE6xWpqL5cYgyXo9Fz5fLANjus8DVVIdY/tqB9RvUZ6flFBajJZ4IO
Gzi/dnHJD2mBG3uQUVZy808/pDE2CgdE/zBHRGlBSNQv2YwznGWS4XA/Xp2wjZ3A
Tzq2fwHjVvi7/wwVcmhUBrEK6C28LAALEoL6snGlZfrPQlGTyMt1s7pCCTY35yEH
cU0kRV+Y+nx7puV4KSTs+02Lc5MJ+F0DpvB/d2LCjhUWMjN9nbiMD5PrDMND8tWr
PazHl0Y88FVoak9JvzQqmay+aA7zAb96zlHg6BMFaSucBi7Rew4bg1CxCkJ7Yz9h
dih7tqI+dI3UelEQichqlRkISPfdX5kiTP7WSySml7g5852lfoYDeYXO0lN7tLbX
tFyGEPB7/cyiusDiS3RRIzq+VHSXLa0SBN5gxcjULjGrevHWDi2pN2IaThOf7Jw2
FNuSSHD3+bQqN7TdMyBwtuekkCG9hyzEqXAdE7uuYwv5KG3zzYVsi+jd8BD0Eoxb
U3sYenpuacl1CXLNvZAjQ9R/epO2kK3m3Wai7kIvZAZn6vPptDkGL9VxGccVHsPl
ZLUwx6IMd03Pb5dxtgubR0Pkdv8YNYFkBGUuVoqgm99Virz9aTbrqlChPrPzVT7g
xMRtVFBxBZSH1EB8aL4FibbYua9z+awshcLZMY1bqHwVzogHC2O4UIxCpOPL71Av
MuBeewl13ZtEFO8g7PuYYL/x1t7fFkNixQNOMFn6pbhzmEr8h3dyYNmYSR7r4Scq
jrzuNlArClr+Gb8Laj/YwSUuUX45tLGUxffdN7AsOe6dvsyOsBi/jzAPxljw1JfE
wRTTDs/pODjsF2v2vM+MzoNNnitH+fRR08zLhUGSulVCp2nwxKXN0qI4/79Onwwe
kfBJ/Vk2509/7LkYhKdPLNtPTwxjmgoFjjaqysjxryrwWauEKR4Myrac7iT0zhHh
ye/084EfntPe+QdvPQwG92gc+xIxUEt7HgNLBYgkOVARcbnx9RQirvEstTuE85Cn
OYxb8fw9l8QlfKOUb9f220G26GoDrJZP0V+agcYdRh53Yw7UDpX8FwkQTpqDTqRY
2maZ2vP0MUDz0E6KCKEc7Xvht/9u0W1hy38Jnia7859UoS8HDP5aXPBrXw+Ca9t0
ugREvTyBThP3mPoY3hsMLPPEtzYtCCIvNKOrlsBs3ljlMa8PWJH6mB6ym9103vBT
KQN8B8ZKNvUai0oPC7epfvm33LqIWKhWm2w53bHza0Jeir85QC4Tx57PIH56nkS9
CukpNo79ylARw0a94f3Cp1gnNzBxeq2jMWAUcram7unSPIE0t/sKuISy+42xPkb1
sghtbyccnxnppeI8/ge017WCQMmOXu5v5E8kLpFzYtVnpBGSnVFxLKDAhwCJ0zBN
7d4k7/D3Atz1PDbsVgJKAWY4Ejjb8JQqHj1VW6EXT4OSKgkyahXGRf6XLRpwUCsD
5xpcfZKMl/VeEo8xQ+HnvYFfATdmO0JsTkMBEHWdZ3/+mRZ3/Gff1eMVTP0Coppq
qOQYw6FV3xQ7AfFsDrmyuWOn+U3yPfCgYYeZ6h5+wqAZ0XtEwhNWKfZVdfbTQ1Yb
xck0plWJcUwXwkkeGX68GbSl9qSUunNLWtEDT3VFKQLlawkWdfv+vKQdyratGr/U
SnR6bIjCaXJr/RVCNWIv8k7f5vRHpRGPNmXZLZrXfELjySn8ss7bya1KMD0ndfSN
3r+6VU5LcYonLMKkU5NbsUySS441snbvTWM2muDKVKqvA1yToN9yHyKFTthY6iXD
1ilUQBje/aB2uWdPc0uBa4lSU0aRjGDFDKsxOVd58QBPqwTaAlAvkEDAxSQwjkxz
Xnm7wMDgfIaG0zxacFKrDHeCAul8E8ngYSG6BTCwg1wCTkDEnuzPXThp1rZxgNVx
/mOqHim+aIP7ULpvLE76oaLKqGhfWzIKVHJT2j1XpcB1iByl6VuwwfV2iR6+h1MS
gagrcR7h6pLPb7I+ZiqsdPlGCiuDvAO6M+XlVd/9EYi48ISazzQA3UFU93DZ3x0e
a3F8S7HH1KnWwVU1tYUXzL/ylrkoJ3JjyRjirEsqr3tdmWOjUEalV6eGW1GbxR+U
BWrF77jljmf8UkVQ8hr49QGvuHO7st3L87vwurAJpx+0NcFZUPWOUfUIurLVamBL
4QGX5H0Z6o3YBPbIti5a5PCD5euhK4glBlXTcAi7ua0mS2SEFvGHadb7yoFtqH34
Dl4qktUGbS+zrPFTQkPl+Lq1/xuaNKs3/DSC/R8HfIZ/5/tv4FIgwBYS0VMDVKI4
YFVjU314sp89kn9QFFRY4wn/XwM4qiS2VvCNKQPIdUa4ZSaJ9tqs4Loewx3cw2V2
OPtbp1w11brdR0PwnrP7FhBftL9sYiGC0pntXoLX8QQqbd3lai4NmGdeOEKEXoOL
+ahbS80hUqVuJi7OUUqedoFs8BtKpvo4E2hSLTlRm/HYQrTkcX82r5j5ORXb5AQb
EWyogHoq4QawlcJlTY7Znjl3ryk7ASkmWI18zdgbrpmhPGDpTjnYTX37ZMXYtjpQ
AqzIQqgaSHk3ivzvYAv7LibBlpNrYx+Zw8P5x7zeBwpzGtc06H6YAegtvttXIcDU
fP88Q1uXD8qDx0oKw3sN+gHzra1Tj0ckxQRNm+ZiqIQjCH7IWDzBl23U7nQOKltS
H6WwswLruxWq3AMCsI/fQ7Pz8IGjvTLLq3mPYnL0JB3K0E0nm+RXp5Rxvok3REUK
rMpvDhTxF6/wBt0qb/YI8F+J8ECTKGbI/N19JFmjDfz8Ykx08/6MsKC4ta4GIU+4
/xUH4Kl1U387HmTvpWllWtpRsLOArNNZ4Sm/GYkukKWqpk9EvbaAxxVmFXWOAb/6
k3PwrOq086uKP/nhjtjjqEfbfzx3HErPFPEBp73Jjr3FA3F6oHZyc7nZ5dZVlW1X
alkxpyxmUDj38OCntNqIPH+iG6JC6jbigQ8aqGb4JPuXlN5QY9Ry6AzQNF2gNYGo
w7ZcmjnF1YKq2kCk/tJxp5T6E4ahkbMZNNSCh3k1NfUkv43TaqHecY9E+bpv2kwz
98kuV6SV12+wSEbXMz+FwrdvmFUYatZyrdJE3j2h74wU04aEUzVYutAz/60PSWHk
Hckv7GDwxoMdohzO24XOR8iv9BPic1UpdqDwwJAIZnZac98Q7paLvaGFJQMAkmVs
CWsswvFFBfdBQyYjWHhFH1DWVRk4qNjBuxMQ2oWKhDl0I1fJ2D344UnbmqMyFbi4
AaP7IMFaJGkW28lWG+yYWtbxJeS8E159FJVud9buKBDp2o8Fnv2nl6G9orkfQ+o5
sYyrkC4BT+z0M88NMB1gNf+v0ZRzf0jkVGeC8JNE9O4QTzNKhzV8E3BOvI3TQSf1
jLB73nQHOmefyLi4KcKSpu1QfVC+gqOqT8dSk33HQj1Swt3GlRsamU4FIBDNbUvu
BTLwVLOi/RcaxE0nwsAZ9Z03f0BZsjszTnIUnjBsP3pw5VPl4gNV+USC8gQSQ6ie
a+ERgTm/+VoRgoXC7wRIMgBRn03JhGoj6j0WJOBaY1QLjjLg1ELPFzj2rDI6Gmc2
SKtO0OX5suVRx1FKc5JTYGfEYrs/wzJODaiscK04FftJUHmXf/BEITg1uIo0mje9
T5cbOiigD1iQtVQSCwNGyrglkVU1v9xLZvZV03t4inbGuJkznDgHw5IVElMigPyE
UG8GV0qQmwjjES9e/oISGWK9ydQNjk+RoTuDm2H0+9a9XYquLU5FHC3Kd0n6wftC
3ahGqu18WWvNpYjuRCITT87PnJgTBQ4z6RJiLJhargTRYsGfkIUiKaNgTvb8M7A9
RrhuU2VF9FKlZdzqIfTV3lw4Xb6wSyfkBrzaWEmaq8qmJmMaSFY+T3P+GsrJ6MYm
In5vAregOJYrod8C77mvu/Y22s67d02om2zHljQq4fo0EcZjA3gbp0cQCJr5YHbG
28l/+4EwqCMf1Kr9GysPThD1rvC8h3YDVFx/RDT6Wmun56zAydNI8mqcMpCj/xmv
3KPPNIh/g4CjRTRlBtWqr7tt/JUWo0lRhKhaE0tETHa2BTcdO5pje/ebo44YHVmE
E8KCsNYrcDkq8G0zBsJ7Y1zTXvA1mL8zYU/WHcggdGtoGuAVQGTp5DxFxvJYSH3a
Ov+JaFpJhKObyp4IUkjR3d40HqQwlkOs7IKrBvZXL/8UzHPNQsnK1FQRofKU5aev
w9Ba7KBOZohQuAV9VpFzYiW1AYnoEVbmOBFE4Em8EDa1EDxWQO07uLKWGGteiAsl
tr6Ocmy5gSBRvAlsDopmR2fuMnATWBY2JQzP5I4Y4EefeDDpVu2HKZ73gwG+x74X
1fVOCpnpUG3hl/AMWn/Exm4kUh2tAZ7m/xWbinN1jwnDiYk7dAAnt25OEEBLbNte
9MPuZZwya75O9cTxInLHH0E9Q2wvs+WaOE/zSiPVD5y3EYCKqzWmON6QX6TZgM7v
+njD1HBqzuO7jgQBWSSY+QwBIAh+FiSpNPKl491yn7oTT/ZTCgFIwdLAY5vT4eui
9UOWRv+AePY08Q1j+X+Zhq3Ud/IIbcI/PG2Fi9QYvE0rj8ii4Dd5oqGrrq5IN8cl
ir+Ax04D+R/fsOy3esffk/mn2l9tP6rCetY+7/ZoBrpUOpVwRfiRZjOV6Hy7cOlp
sTu2nRgj+kbu0ukEfWpmANEnZyh275hgfkedyrNeaWMhc+LU735OQjNyObXxYOyy
Z/s4oi4vjtMWEoAFxjcamMmqVXqi7iquVrkLkjZhxAW0cAZPoX+WwfpfSDK0n1De
xsgZ2Xl3/QYg6U9GWAg6uDnEhA6lxKCTq3iJPzWzhucIEjsldE53qlpXneYI0O6F
s6Cw9pSxkzmmhM2EUkcjX1NoOVgVJEgraqCCGkVkuAGz4en7oOC1zCdV3eZB8AOJ
CZUXR5w42rg1nKK2TJyP4UB1yqRNXvdn0dzglYVFYxgIYb/IZs7Y8lAvSDHi1g6s
GP8YOz35M7I4pa5gcSozD7hoIfiZuOtyTsSnHz6Y8R1peqS9P4T1usf/SEJeqlPp
nE6I1nzWgddRzvafw00niRG0COZCka3jzR0Dv0JQ+91ji3Lpb9WDiML+F7zs5bNt
t2TjaRRPkW13f9+EJ/FPKCeWJbSpd4DGDbVC1AgyIXpqgzJYp81jxT5T6D8UJndP
OrBE0u/h3nqaf7j4PswdTFUGch2kz3e4KJ4mkcX1KGqkufCtsAudMjTJtLh8CLMt
O1rH9TsogV6i78ds4SJC0yjCRpo4timldx5HXj6KepC7ZVw5idTdWufUcrHzoamn
FLwkgk4tY6TQMmrlmW5S0q6hLh3Ym/VuRLGvz4MEv6yu1Sx5zV5ADifkzNJrsazL
NLN7T4gJqTW+Lqo4FM9Oyt/EeQVAzRCmVJlaxdrnjfqpJEGd6FShIdp01m2dNTez
xHnp/ka1AwnD3v1aNvZFDKMBWbSNhykuVwLKbFRP5+tn7O2BUOuFFzpa34Zt4w5d
vb5LvLNKT1Sq/iI0KHUwmt/8XP0PFCB0hRqqDiNaV8FlU+wl2iWn1NiX7bpai2j9
tS21zgY7xgJqBlYR2zc4Hrkd5Lrwcx9zlbz98jBJ/oSFwAqF45yHblM2Mh6N8JOC
kCH4UWzObosPNmLPyJP/vS6uDVC7ea/qGCw0qoaZFJbM3FcRN0QTF9pxm062pO+B
GDB15zOtWqpX5wHEfVCDjLhVZ3sK6ys7AL8C92ikNvBq9P1dbCMj+6NflmmUUF7n
8BN5NVudPwrmmbuJ0+uIzW64rhuqsNpY50maql9k2S2KakQ2JT/UOPq0x9ssHE92
nOYGhqoMH90NqaoiuCL3JKnbKSytWa2iH3wM2RZIxzsT7EXjzmSHd+YjZ44jxuRy
5ul8TakSyBJpCjWOijryR8PSAVxaQ8sziD8o1RY79lKk72tRngDMHH76JqWoB7vi
JQoy1M0VeAEK5JnQ4n8ZcUt+ybd+Xc//NQlvdEmg156DFWFDjZ/srzlxlokVVjet
xxzolqREDNmeJmbyY2097aL8PTyYFjXlHnz3XBdzAFwV7iuXpx/fUFB0zEe1dO2O
0KArFR5jUoULKVjaK6uL2z4ymDJHpUopWjEpSvmoQEQg1FwXnpfZIuWXCsRWlKuV
y62a2xmvE0CS2dBMgFHwkrKSEIOXIckKjUJER8PoZjGIFDYBMcDPUv42L0uNDxAR
q2qQg3r2u+AG80TY33Fs/2+ogc+SdDswGYF0hLxCTT3H2SgO6Yd/kAikYSwPSuTd
S1B2ueTcxGYyn58NGr7qgrQDTtoU41TeSD+qOxrPmrG3D+1S/7NzaE+sF0GdKCmp
s4AA8sWiOgB3E+KgQiq1GY91XvTv10evryYM7AXPDvwBtd30TUlb4+8hPi9DZgWk
129voAnTT0xtzh2Q3133puUW8WETcPr2bZlUqetujxRPxPtjTZUi6LuEtnKYJkg3
7Eg0969ebNfjUUoJxYZ3+Py6045Pvb50IRCVXOGr/Sd0J5MtpNGS4riyGdvCFq+t
TGWFDvo73Hx3trjATNAjtdNscNtJzQpdGSdISC46QCifvhGy4jLW68H4vfFCL3wS
yaJPet1e256+If6uL/Wk4GjVfR2I8pnFB51FG61RpcDdZutbU+N+dUH3aMqkU7dr
+VBH6wnJBg583QZC6dt3l/EUFvSDH2CEGA+oQlUy1mYi+23s7KZGCT5QAZuulQn7
Td0NT97tQAVTfRt8AIIHmvprJP/pSuF0lu6fzvNzPzlTd1VzQ1zDLbPl8r2tslzn
s4aGZfRjvsGEYDYvNf+DWaBxJ8GBkzeC3vJ5eGSR/JRTloI+0LyCOEN4UiFVa5ef
2s1VFtX9De1HhNvdpPcKZlwfLO5DMoLvcsfsD7bi+95NHBNkRRLNu16vdFduOZFf
M4gFQNizBPqU8eXXa2NTag+vOUFrfh5hbA+Kh078/+maAs2bhT3DiFdPC9VA7FJC
dov1tdYakO9P7ChKqS2YIaMTGaLVlM9Eh335dtGAtM/2fEwG+tpvJP+JEUlCk+IT
nD5sIYytATgkt/Z1rS1rTE4F/XaF/0PdP5uPUUc8ilQwnDXsc6PZ1GWfERDeuqTZ
DsLFY1gNKZnKokB2joqIwGB+OKAm/oaSN70S2zi/wyLue0dURAgYN0xEx5By80uo
P/h0locWn5Lu1UQ1xIsuGTOM2dcKQcui8MRbnGZI+q3YQyWEZxgqd8V4FTx5dcIN
uPPJg1WiMDZ9tc1dbKdOtQdcgEBAtUUS40MDmLr4LqVtzSoaDAHLwKlPthTAf619
rcyp+MW0Q7ZpaLngAg/RF5FZyEEKPd5OxibBM9lXasJw3G0HfaoHSXEBIGiNb2re
yOLvPIJJL6Nz7Xghdbrf0cGJMqcfwFR78OvpA98uhyFbHuHu+si9KUYD073QHtQb
Fnn3OunSK0tKSNb86J2obUtV14B4TniSJDCq7qvT4Q5weUAFW8LeRObyJhDODFpT
p6OkKUvvrszRBd6GLQmW3GchbmxO5mqjMe8te32siaVQe/KsYj0TRdJQHaxoHLp/
JAVswxqK2wcvn/9G81oEmfzPwEibG/0BOlyBfrFuI4IIHmCkXjlV3J8m8lqnPXgj
tH49AUwg+3WoKcIhnKX8bOOE0NGe0B8WVDU7x3GQ0JcQubAiXfKIXJw06J9y2Zqa
rpvFnfNoP6nU0wgLmltaqhsPO7RtGWeYvWgtFlF0Nelqut726ENDBakARZczwnxB
pOgmA7Ej6S2FwPk16heMVdpka+rBw0xEscUCHsPsdAHpZlDCvMo04tbxCgNhOXt7
4DW49aDa+TrOSmcusoiaqXo1KuWVwOMIHGgZhLOUDv/Xfhw+gluitaIZEMIXtyyQ
i8Z2D52NOHze3nV1dzmJS/cmvib9lylBeQPQOMk0ftdd6+vPENtg+iBkBQC6CMfc
l4MFbJCjRBHX19qKH45S3I1SIJi/Q01uJhdkGCRIWXdzITtUYJBnWKRzRJ9UTmDQ
ULoUQQli0nmbE3pQqWYQH7adfqiMxCszaNnRxkunHss8Wuy56I5Ftz4g52XHvwQZ
4fgYB8SXRVJZI5iV5lkBU4js4Ik2UZji6LH40l1gQxa34ELObQvlyK+Qnb9f/i4h
FRJNsF4w6fVG7sr1e/5mvefLBsmzYPTp3oo2bknzTjGFp5LYYGs3ecxcpxkwoaCy
Dov+g5Rgyp+MFKEQMbjAuZZFd4kkO2Drb7pSY+rIKLXBkLUoGaTzjKNFhhrgWjtZ
Bncw/8WqALR3xUvIxr+D8eV9EKzDF+TeSDZhxhmaSS3kVFIlNPemWCdv8B1x9lff
4L7sOtlus3oFJZUHzBfTLNHXc1y5ec3PfxLwV9xxE8h7AS+dZxz/l7hYyjOEXwPd
VtNZmYADE7/HEMNignjOk+f7IgoN7YU2Dc9krInMuxS42RW4BgobOtWkk75PcvA0
nC1/AkKDoTjvjV9qCNshzp6UAFDxHL8EcB0IER2TatK4nfVl4IP/oo5T4CBNzYQe
17Zur4fUtacH+c3GA47Z2IdTZ1ZaFo9yZIQe4lLORHFiJiCeJJo72GNwUEEThFcE
NWtGtrEd5a3t8F7jRdF1t0ALXsEx+uVmGbIeGaQbMdoY8ILgJe0NDaN1vGeNL2XP
mGt56SpKGADWI/GlO0HTgFkdsctrn/cLKCdjLYkVMSVtwtrgVElzmmo6ErkNvr86
U17MCLjT/4cU0dOT7lBYiFmE7TO5pmf03YIqPY2AIyI9moPSdkU61CuywVgbG+5r
NxoCORPTtZSuKxZVeOuU/Ax8B+Xrax13sYSUerEhpbEytjLYhVoZzeogxZNGece0
v+eUJxDfObi8mu+5QUoV1HtBic7Ibf6evmWG+S5STH9HjK6gKAHoDzSpdAlFJr5P
xN19d69/fX5KUi5UgHGaBj4Hxj7p3k6tG1T5gMSO7U7hXfwaqpEdJmwaOuAuzsau
3b7Bn02sX+ACuMQyd1IdjceVGiVRGTOc9k0wd8HHVQE58IPbOHANw17ytDmFa45+
yOU1RK4yHwIUsqsUt5T61TR7Wd4mfO+7ABo3KL5vGdddGw7IjBQEfLECotClQu+l
OWjZN3k+DAEN/CFHEQD6SQhRtGt4x5WhhnKdFtwNPNLrBFIr6sUtbzYykE2HZFC8
3aWJQBX8di4GT5tK/9FMu6WcDXX9aTFdYTno3B3dbZ9rWXhSbEv0FT+XTleCFTyY
zEZxs80A32QY7Fa+VjjrfufEO7LxQ9+ecwjonVbTwlqr1FOIrZNjEyngt3xkLpKm
scHQnEa2Vrwvrl2SHRUTDSPJhrJeysJemzif/KvEDV6rwmZgN0QQyQsL2+KZ3Twk
yzFVYIezTWdWOqJumz9JIGNnw+ylMHNRNpmoW9qD85vPh0UX/BA531WuDCbwm01p
0n7kctRjazrqyo8njNiAQDQjixCloTyhKoj5lZlhLJ8BA2yh0bIVBQ7L5PWlGnKp
ML6RbDjhypbmCBoEAy4c38Cd0/nlpi5RLV2q7mLIyuWj1i+QvS1ddRpHUfWOJ50P
4DMgqhLu93mXKM3EjdWIlOO6+VDh1n2BKNQAgscdaeZKbPiF8M4fF7919lNvfKge
hzm8gWBp18uTYydKXe81vB7aeqSsg/wjErZbo14P7GDIQY+4/IaMj3xFqwjWBo0/
R4vgF/LhB8u8VVI0GTKPuwMUF4KCVMins/VXWcTbUZZNAvv8xhQ+HeC7vBt5H13Q
roL9fPtG2qweb7rI+4nsZQdHZtyO3X6IbmCuxTptjxltFdqpf2eUYJGrs9tcaicr
TVHtjiBaKMm3NUAJ3VaQoSW8llP7pPm7Y3xLPR5tmwFklOiDvhX/v2VTmmsOxiTp
o/1UidfUPaySVRnk2llUm7B+OzhnXwh8vUKnFuvZ+cPtiPX5e8wNfqXbYwQGj2/R
sj3byR/mw98EwZtvMPWW+R17ABZHDbURkmq2rup1o5SIsfJc3eZKXyBt2hsYtJGb
bc11wkheiMWzrmf7y/F24QK93/dJJs6Br3JGJfeeXcuzdaPYpJHZx2XWhIMmWFYs
qXYv+FwCVwGRNLaI5u7wDi/Va3JvxXYURhqgD1Al90YAdYl5ckZ+Iql1Hpu5YN6Y
5iTYc7z/KoAhGoigGdVLuYSo8gdRJUWIWIq7iU9WEcJ8a0Gn0+2YgI6Lr81wMhfG
W+sXpZor6xJdofKWb+yiGeO3IseOb1nyOYdlEG0Zj3GGxmQ9pEIqlF53AAQI9FOZ
t6JtgVghJ3Xd0glbkMf6gFcZA3QOOHL31I1UMdgm3aAdp0H2eRHcdoheDki4b0UY
LnqmDIRNrI6JuX0hmIidwPl99W+ZwwyXYZAqmhj28HqUX+5/TFfdL57WPQbqIbIK
vA7AxX8HoXFddH5k1WcemC+fUq+J7Sme3BZ6dm66tTXgHQaQQgOWRVpRkcoPQ6qs
MfZk2jZq101JBZhHE6MPTotq5S9HHnhsNA5Uvm+H1/ZA+CE5e4tfN3y+UNYe0ZsW
jK1f3olBNPMSJWl2yMmhijkh8JOm7rzUSuRWQTzLy+IySNKKWO6nHx/6XVWKleXA
UCnyqMY1EyOHsiRP7Iu4SRpX+4tAcsAB0cjzuiAnFlBf+gH2JDLgw3jQKKMEyrxq
Jvy1AarI2h3Pw/Yt8+EukXPBtQC6swpIrCEbTel25Uhbkig1oyjb2ZT4l5YcxaHV
bMTl2K9BFCNubFe8Mi+SmTUJGLVNgq3GD7qzKKReXX1OUQivbHQIKaXlOJbmAIc1
baLIMZsAWa6/fXF7fbDfVXMdgqQ9369LqcLboqSV1B3yero15fNyISbGa0i+v1tk
mZCDURFiYn3G8/Z+4j14qWFcYitkwizSmXo5RLea+S7AqlCqhiFIQc4KuG4STQvD
JNFohJo2mB572KIvzpVsiJnd/RQJVAFRPMafQhpi+8NTql16lf/9iJN7wh1F9t7T
iC0357vevsZ8s2GjwvEJkuuAbCXgMMDYO47INLdtIs6Atpq8J+9I9lCx9GvfBc4m
qf4FcVU2Y+TMhNebX8rj296kFsu/mTOuOJf5NyDwSuyL+uvuFeosl6FDNca5dcG8
vCOI3QyT8s7ukB306brHfywMOyvX9Oh9knlXTOsXNVbo4hjpuKdfr3PYefjmroEA
Ro/ngL/n7nlx8K59ZkqntG+ts3/z1TWPgdxigphEbN32EHXYQJ1owy+QGMdg8JEJ
pbvrxmtnSNTA4vPehSUMNplQg8iQG/7EOJ+xbKJiaDiidF0FpWtU/+yXvMQWmRzg
wmBk+Y4OvEP0PL1N16cnKUn110LztPw7fU9DLvP7BTOTOXojmtpGfRRhwBvT2xRI
TjjtEykii4OJmn6JH01whhnosmluK6BJwnuVxRfA9hfSqFGIIk+J1GG7ZmKZe45+
bB91sUhKIrj1cA1x1F4ew0J+5M3VunhWoDBAWgBpI8ZYU2pdBlKf7DxenTgEM+gb
Rq5Ik3x/4jAyeZv+7CzJqxo8aQjqumn0lmCRfDXqtJV5GE+6KPfIrnP9Oj2Ju6yK
9zQTCk1ZnkC8lQBRsmI8MUywJhhtR6ipuw2nAYLoSPLvb948BTlGTFzSgY2Yce9q
bkOHog8mLgMUj55a7LkINpSoYDG/OwvZ2QtJ9pagzKN0QAO/a3uYvpCY0N884Mq2
RaSyH5onT0uJLvwpnWmWbujIDYpZ5462z4nWbl52SxLmRzseHwAgJJfstaDqWCLv
s8j2Kf6OjVdJ81RN4Agh7PucSUs8kO1KTjovRHHqGJ/cmrmdknrY+jE2OsMvdPGy
nV5vdmK4MWA5d5V3PAFm9J6oc470JDK/I6OdPQdCIGXp53shOye3Fw8vNticlKKK
bvRmQnYjLqbcVBY/rWhYFod0qItJOqFejFlSkrXKPCcNbmnxZxdK3Umc4Dx495Ha
6/k2tRnFqmnn4EB2fyEdeJFMjwMe6Wu4aBxO9kwXYc01TZA96+uNU3Q/9r6UMNuK
89FYOxCzC08qZR4OcERDpzbXfyQc7HMZ7F/k+l7qhgc95kNX38N9mzFFSpK3lgAV
8lfg3n3cu66yILgPYNkB4NwtwAUuKSrerOWO/inT0WgIQTrE4EyNKj5/9E6Wfe4x
XJ0Snmdtzk9nYa7MuXRLlSo2Cr3udRM1w5oyqaCDOG8x2c7BHeQDzkqqvn+BTeJ0
rYDVMe2RodlnPoVQU6vTPYMDTO1d9SRcsDQi/X76Q98qsqMRfgbi8aoCxeXCmMMq
9hn3YYQCXw83zrgRT9SQ3oS/J1H+TMQtEYoeQlLO6jIAuG2YMt5qyEbsjGOMKo83
slH3IES10+9LY+yB/fNjIXTpOmkuzJLBB1XFUSg//fMSRYn5AlbYwZpcr8//OZkD
k6JKAqcsbE62TdMsG5ouPRoTdtTpJuNR/a1elvh7EltxS9V8aO2SkdPKycse0M4D
RfxVNeQMoODQQtm9H51+caCHKy9jmeGQGQT2olwU5C2vp97x552O9McyYe3Wv8Bq
3o/nlHOhSUTAvQNBRPKS6cLUM6mVDahNuAQnApiwPRuvqQfMIvfidsTG6ZKht/0u
AgoQZHxvNdlGX+fyRzAZas5pEw5jjXav8PK6ZTph7GwuVvimafOGWA71CEsf6jr6
UOsDuh6mzZYeCsEeSUj6NOO0nwtXYGMadKAoTWO2Dc8qDEFT/BrvO3gmdio5yaDG
kIibX6FBEKqPTTKA/6OLWItecc0Kf1vU/CqBgccR5rBLx1wETC5pzyn8eQZDX2qj
iqUsHWdflKZUWuqE1HE7AoSiuz5NFSblF843AClFWp4079v3Ife3KhKMkd/ryYi8
L34LT3T85ma2HaJWCbMIew9euQG2jVsK3xAZguwLOrek6fG1LukysnrsGMgD92ZW
Il9WPEZLJ0HfEYIrFNLx82LiPCEH2IPsWe5RbQtwQ6CejFeWW7ounLK1U784IsM8
2IYMqoivDCOW6+FRqGoPFrWxSj/bMOjKK86y2VsyCbhyewfgr2Dm+G5h2NbNj+Z0
tegZcNPgxo5ITdnm1W0erTVpa3+vuhQwpIVG/xXskyyb8oEyjZWbDmP/d0Y61+7P
XEPmSz928GOlEAmViWZrcwr8tU551u5dIFrhPz7faoZbCH8uNXbLDkB+M8K0al4+
qIufy1e8DHRqIRrwkK1RPa86+BM0h5J3qJBBtPRKYAVI7YBAVgLio2CJil9YS/et
CJ/aTa/vrgUnydRI2U7lwFTfeh8KsuB+AT1qN1eoG6EuNeXdXiBVaR8VKPHwESxv
h1+6137d5cIrpOfOYKb8aKOPhLwKS/CEAxPKihzLxWjC9XVH5hgnYKP9CixsjPsQ
a/+m/TRDy33+EG3Zpu5UBfuDukpyfRfLOIHmw24WPheLJZZTKAPM89R6pT6gn17m
Udq7sDe09PqUwWHI1nNQSvndxSCPjyBLx5KR2lcWR39In/UH8FCKJKhcmBo8LizU
Ir3Ej/SgXXtCQlgshok9/CZPvve33DUD76aUrwkVE0feWbTb32k2e81qDKYuUeLk
Cy/nI4t4IZgppSBx1WURMj/GrnWyZQgGIBMKLLXGrEoyb1Bdm8nEPbhHNYbWK7B1
DgEbx5Z+0UeCCt3e2MYZIWsOHR2zmXA59aKGlXWVDRoavC8wS4rIUbvGf8qVOY7z
97ZgkdfEi0phUeJ6V/cbVSgtXQWCuHODzdfacq+laBlNQ01z/HzW6f4LQYoLOZo9
WFQQ9qkVQPxaQKcvvD48+OvkHqAH8s4WqDvoP1ON4o3rVqlNPERyZQBkqIBrXERo
3E8K3Uhaxo4PMfjajx4ogRVNg3qzlxaO7Rkp3tGJ2GySmL78g3L6+sQgmagNJsLe
KUN0KVfuib8MSfKtPAoJKcfdiQvOpfVoYER9Y03BBNHxTQflrebn8BgHmJ5ItpDP
/wCsRQKmzcBWFBGVMESgoZVJ12IK23z33wYyQpGuk5w4xo0N5lIfD0FdMfdOQEwr
Erwt5qDJQZWH7a9zmRiEReDzFBmGzxsxcc7cZ0vNj4bu4MWHb71cuXzkxr0IctDI
HH6mnJN3A1cF4zAQPvEAPEIunxbaR4kqKqTkvBbSSTBZ5/g3S710vAUlL1/3YV1n
KHKiBybugYyshDvxtDylahcc57iXjO6dif09FhPY3wPr8BrQvSCOB2SFT6s4uVCZ
TNrOf6pt3mgvuCu0/JohIbPjRKeLyUDJ4P9HMolc8yxr9514TjvDz+PUt68unlvc
beaoPtWMBWlBtDHO6GjfumwLzf6xRFUDOzYLie4Ue0wJl2M6Lv0ESj4oZZ/yVbn5
dumElQQUKhqEmxsbEofk9jVd8nNy702GGE6OH0wEt3sr+ls/RvTARoyJd1u3uC3o
aefQljHO+RnHiIE5i/EIVRisbkT8BUY1WaeE3cQiJj5OUCWLTBcG0FQaGO9l+PCu
eUW1820dEaCbJX8zKjT7HepuWwD/tLOfaZT6DoGZifbuYNEj9/h0PM7Gu8OIhNse
p4aaMpxydkiueKulo/tRBx4vahV5L7Tf8Y1ypXr20ZE123dAoNppq3WB3OsSiUp5
ZaaxCpdk4Q0fjdxEiPLoWJQUgKhu3MlHAnb05kDaCxQUlO8wp6GGZOupt42ZJTkY
DIx8hjyWSwBWb0bTsuWJroQgzbkd+xVXhVqPPPrUipRZrFxxBbYG0nzev2MCyTFn
Z7VrJEyL9q8Cptlw+rE1E2G/7jeuTZ5IOB1vZq7v7NQEZS5QVbRO+rXAvXqMrxoH
QM6VvqtCebWLsLToFN0UGjvy48ImW7bXVhCymjhQ/GDVcHtNWRGjzMWC8n0uDyRW
ncZM9V/SzbbvOMFyC/8jzSJUvHuRtrgZVxsEe/G7tSwP6+40XhcoxWcJ+vD5ea9O
IbsQJGKLwrI01GRpZcXkugOVmr/r39dYt6E/Ape08nZ5+uKa6Bu6pMFSQF2VScrJ
DYlgEhtHIpgy8U28dSZivWj+AMIAHt99UOQzpXwjpbrAKakRkkLls68lqlXghm0C
+l3wqPIEdRf6/+dF+Flq8km6iFH5YgYhhCvx8UexhCbLaylRpRMNPbjvU9ZWXmKK
KzrPwDZoto2q1fYoYhGZDsUtfwJirwvA1/V3sdciX5+XfSQennoSTlVXOVJWJQxX
COoSj3gByrRobd0hs/JIq0SkeHD+1Xt/jNK9xPPXQaNEOSsp3R0khovtPRj1YVea
2IkvDb8ULWVYuj3Re4tspCNNFTVUHK/j63v4jjQMYKxb5ddTU6anZ8h4l7DczKT7
x2Ljd+FSuuR+3/llBIE9+kDKM5N8HqmS8yxRz3vCGzGKuxx/FJ0iRVqyY36xq9Zt
T+E4uoknDntLcNUGH6xkyd9alYgh9Lc5dVndlV4tgQRbf5DTQChHqj08CvyFWYua
QEXPZEgEOMcpWEqKMrIkV9QWqVfhHl3MC/4Xu7Aa3sYB8H2vid0LNJxGyXomvLU7
Q3bGPzhM9HNiDVgHWoB5we05uJcZHpTjRrkRtLq9t2sTaAtQLgZTUSoKjgv8EJWD
jHN2W6Rai8cS1y4YJ8LkRq3Kk5jbm4unlVR4rIO0cqqmkzoqlDRxf2rdNPegGOl0
Fu8Lp74VpXykqbOPxwCEwyYtdyi+BCrlHPcm19b6ywM4Lp+LTSq4BNbhZj25jzfH
4VKzjPduPR24tkcQtAQiJJXdg31XODHfGPFDhdJiaYEYLBw0Ch9FBnFxAjZ2xvLQ
uARms3LbfiMC8xXdY2n00PCxZxi5H+1K/JePs7HlGVmhGuCXLabRDQNJf+1sMohZ
DdiqYFpvhM3yQgVBYWqQiCLTS5YORy3FocD3/pF6RACIHZkIzNMsxELGCSMG2shG
L6reMYSViYQtRxfu67HArd0yzkg4NYqkfi/moLkfYYLDYoVk84wDJx6ldOAYBoVp
RjqfGnAvZImdFRpVnkuYxbcGKwLayQlzl7xNmzuBsCC7VIxacoBvz45r5eVlonel
ls3elFGCdLdv1KxzxIauWOJFh/7uiENr8it3RzjkulAAHXCxvYkx2wdL/FIziQQN
nlHZD5HPEhOdYj4VFEDhib7Px3gwpO38F4928NIF3Flgl6d6vkVPksSYKK32FIDz
4wKfyz0fFE67Aegc71J/lSzBF77uH8XfzZ6waYYTzbYQFZYOUKSIQfaIgRayJFXP
UMIyvtVb5avAqOCuF+aKTDWpq7z5t2HnLZIfNNrUTjpnBGYCcyWHDKC5+nVwn8EX
OX9Lb8qJ1uTMQ2xMI0f/ax9DR4LDoyz2nB/ikDI1UqMT2FO4UoVPsCad31J6CxzS
ZG7aR0RGi1xdhqwpcPUOoo9fEg649zM2YR1B+JEXgvFsEXmeC+NRPHFHWV9v7C1i
jdWADpHZ3rnTVd8pl0hf5jL/MO5G9Dbx0drzI69JHqQsEWKRrd2iumcyBhBzZu2F
PvP3NtGU+yAuTxuwgKvDJyv3G+zw8m0gQbm6R9t2cBfPgTjSzZCwAV5af7jP82RN
0Vv6J8pDiy/ogXTMmBSzFAn+V3HftmgGqA92kUky5tEtXk3x/qHf5HgKdE9lSCza
nU6QobyNmz5DocMvjfaoOeTTUz9J/4Xc+sY3/9w3ZIk05CT3HFTCbyzxdxMiYtP6
FdakXZ1Z0YhIixW9CpTWPZIj7WTsTPiHixWFo/vMNkdjkzdkxjiChHNkgC7pOPuM
kVuI9UvNS+qrvOhSMoSd84DCIFABlEWkCEkSIxpD7CjJqFfvM8VdDOaGWV11HwSF
qMn6wraTuJUxBfcMXqEeZjQYQ/3rVa5QM4UyzHJ7M6BDlGHcfVMXkC4Z9tstsmm1
DK6fuGbIQAYpS/hd2HsF4oirOOCoX04BZFnVfoge/U/4Cco8ks3tK7LYAEy/iuOa
PoNO9lLwF4eRrTAHhRWKc7N4ZniMHFdlf1+Dv9+5hY3d5N+dN1sn/qEcGUqmTeSU
SJ24ppfmOQY5uk+ay6dkJzZ1N49F9S3jQVCaX0St2dodum/AHLnFiqUkkW4lsOlU
sqRPC0Tv6XirbgNJKi0htCJ8Hf5ICFHOIa5k7+AVrYiX+WBfYqIK37ixveX5QmqJ
FZVp/vRAXeOYluCzpBV1AWEZjLorGK8E8vRCLJoFjoD7vGvVKXChD0NFvitNLyoV
3d0JxVqqnR2FkSIGZ0OtbPyplc961T1mRc+eYeSiy45poOe97eAyNl6LKKOmN785
Zr+1Ef6+hbrUo2j742PefrfBqOsEV6DyhtzvPo57Q6aaUng+EtwcDlLBnPf27n6d
dfRUjY1dStDhtl/z1DXFvCRKKR+pI/NuoncMqNeB8UchTwsW+PiJSy6h7xQzuL7y
ysFFXdzwDZWNZfTDxLsPTmBNjDnbZyy9+JWTCU6jfZicFCp+4m2OXhXyCOXT4sWC
vubUzgxc8O72gIjCyuIP0rGue4oUm7jlJy6foL1mlXAGELQwkW4NBDNFdlx+9NUE
Rcl/LE6CxwvdxwWMLKZnZgLIWJa/CarqmkdcVmw1FJpXnYkR88fCR4Qlsn+0cWmA
YgDJdAQa49UDe332MOfLuVLCOkx7/oLzpM+Hbkhh7FiGxAJo0gI/N5QmLzV/cQ16
SwILoDZ5odqiFYdAJnln018EZ01r8UsDcvpu5FwiGGSz7JupAWhpHIeJBovuNoG7
F1nvS3/ON1mC9iH/z5iSEbOkHlWg8W/eLwBOqFQsP5nsPIMZBLPO3xynJhAIbH00
rV65oQXkgYeyVgjz1I7HpXYGLJKtX13csdoUddn+GwwvqAyka2aizL7Eggbl9Th4
JWPfFKuPu5ccDWqQ8oVUAswq1TIZg4+FSO49f82eexgMo27hvvuTR3q2yGvUjoNx
bi2ELJvmGxz9cMq3PV90ch8iGvrT2WHilp+qpq/8qhewndgGjoDeP+WcqQUCyhr5
XAHN9wGzrsnXK47o08QZfqDLye58fF06oMa21TbBv7r/6AEMmzcnd+GWfvVoeXSE
sEQNA4YkIvwL4qfSb7QklhLGahPupQCDNDsoQiRWkzNNPFGoNst5bCWnPreZgEiW
4PNxbH4ebmLKXW1QyvaZ1iTIZQi8XWK7DtExRyaX+X3/ouWRQb7rTt1ddwYLA+LA
0Nuq4nsBy/LdSrDe0slRtFsZpvJkl6L6suSqaO2PmRg3jrPsH2+ZvO3ZtEvYXPhv
9FnhWs/L30IP3xvDhaBRby6lSyZS1u0Vvdli00lNuD2Hw9tSP8cZ3UD9kee+n/bh
7ddrQn7T5SUIi9kQ3omJ9jpuXHiZK1RaQZ+/CNHaXkXDRofEUUBot+PDUAfEtphu
1qsOGXgGctM8IoKTbKfDg6CmI42l4K+QikDs0W8Ub/hhvHhmfJTwC0EaBRQRfjqb
bDIw5clkAWmMhVgr3kM7O+e+FeQhCt5/H1798V6PfGWJ35WBcPZItEhue8O2untG
O6C1b1r8z+Mf0xONm2DstQXUU41dc4IscRj9prYbx+QrKaV+nM7ff7AEUCO2AuBD
1mhI/xkrcgFkarcZ9OvS0N1Opyvs+EMocuh24rx3OlKssXG+Z9P6QhLGqTs5pvQt
4gWC44GMJh5/DFTGP/13siEfECHzeWsCDnF7eRogUysRIQ6ZHEBArk8eFMAePp7h
CW2f4Bek2jruFPBy+HDiySul7GNDvTSrGFw3DHvbFDaBp4X4urK6w6JxDYSKu0tE
Nnsks+YNP2NQ+wqlReWCUYUSaa5qi6435feIwhr8+xdVdHtD+fhTUBo25RtO26Vs
AbigbOnoX3Y5FHUerEMnuJcZw9kNLXWm/QrbXOAS6AdKHjgUXjsTBOFhG4snQar2
oYWl9d4r6X3Ydlcf4KWW70WO+/h6+lw7vQoLLOtKJFSNP7/du3uWBCQuNn2Nz8Xb
wwcY8S/THwk+cgEOHm1Wjvl2V4V0mssx2ySWi1E32NI9U0I+n44VVcfHQDA6HcRa
dMF6b/T/qKzzHI5pc7eqkeaDWwtWC6T6Azq8syVBmE2Qpc+cuAPv7uFupwn+Kd3i
Plty/T3Nx07bhBy2Fz9HbwXsUo32b9ONs70BIroSpb1qVFRWXvFD4C9H5Xmwo2KQ
CMR98fqinDKa5cLa1INywCH9tkN8GPuSSnm4ktebGqjXu54xQTjZ3UBRe33XoM+e
pZrl33uxoqYbOeHosauD2VFAUsv4R5ZnVBsUC/SgaNavV8PLcj19PKpeOCLbVDdx
tkSmrtr9jR7c3COkHaBURP8Vyu9o7ofAzmbJmWDi+UaAkdgIS+KtnfMQ3Mn+8mNR
4xrLyj+zebE5MSCPk4as/mJZlxbWSy+QYNiiUYktF/J8WESfoS+m7jfro0OijNf6
sDGh8m4n/zyFisdAV/QERol9hro66SVcqckks33FY3t/6cB4A8VsGsT2EyZauYAk
jDFjp33g9kpZpi0aQve7SKSq2lioMRek9BHsqiali/xptPn0pxyxFb6XtEWKBw9M
C1NqDEtpnQWOpnDSjRylkGUHYl7vdUXVm7927yT685Er9ayLlokjYewBebn5wbhO
Sr5SQpG17GGdROvv3zVL1ohvsxLVRJklSojd2Tg2jyRyrbvcfgfBeVrF9l9QFDo8
/ZvncINF8JiRyQwdyRxHKXo2FG0mPXvWwCwBBdVbbv0WiHV8iEBNRaUnfBQYYici
Yts6colHs90Pv+ec74d6xxMB0XMLx3HxYUs6/vmaytacgwFegkHEmL4nkOR3RMus
CYhERt7kh+xND2lDmmRAty/YpAy/Br6LgFiAshtaYj/Pxy7SV3NUeeAIDv2h6ZIS
kQaIwpTgAhAbkBvxiap3xyozPCMDFCerXVGK86RlNF5+M9bit/Nd8ZpZCoTLYOsP
x7heRN6hO+C2rpaMlkRvG4h8xlTBJ6SpXaKpb+qNQoCoqYpvxqQFIp10JXvo4aTi
/uJMfwm+a/J2R4La8uZamgg77VXnq4WuBtru5iVhVUdGk+RznEATlrrHaJwsLcaT
IWNC7W1cKKw5lLLQn4VkzVNbJLEgzQKvcBm0HWyZ/oCM4hi/7+N2+7Fp8JKIJATw
G8WbTPBoV8YqVVpJxU3G2/v3r9oWXrZM6N6Q6idpUriQ+YztkRZIM/ze5UGRVtuU
pOAAKBRx9XorsmHAN683QP0DtEgqTJH4GijAYFx6unLaPJ8f3JXLTAkquEmY5XlF
Mw+m9g4gb7eiPEk4qtNCaAMO8dNDdIHr5RGAY0sLQPGFPKMqWvaeMezTorfjqRKy
LyPZFIlSNTFEUxHYChM+U9cGRSUk9Bem4U0uf+cW32H8T39HoloAfRNwSLEg9DV7
vD38qa/PsRLnNDwEKfdj7HQ5jnDctRxJPt4/9bdZpqFgz7VqqvI++dzPeloJatI6
CTLsed7/VYxMVjXtgN4I821vbXUSLrs1J6ZPVBxCc3atqfBudCQvZQb1BFcBNIiF
25CyXhgJmMMiPd7hOz9bZclhEqU2JiafVYEb+37RUiJ8FVi+gXiYgEPHr18c1aZi
/zsLOO3YL2tjMxJ8Jh8e2zbYnfUtf8mCJ4qLRHZ86ptgm3djugAbHlCjaNJHSoIx
lm1iCTShitkF0IsP9jReWcxqv0Tf2wLRQ9CgzVnnM4GwKM2Pd0HcU/fXCiJW4BJm
GF34/jgTuHo/JvmC6Tr4XmhBv9eiX64mxXdYMU1/PvHV+d9PA8C4lSwr5slDOKkg
ICqSH3dnkNHKLLZh/YvEU2Lx412hP2zhqQjAuxyck5wqz3e3b/cCRmshUT81ssmj
9ggYUHSM4NTrZoXIqlX+vfz4SibtYTft0a0tpSXElZh6eERi4UNe1mS4vDMQqmVJ
IE6czFFY3cvBfjhVjpbG3tTIkyECOjl1x+ESW2/PWLBhts015cBNoeVKxetXFvEv
pjQGJrvQW9AuG5O67JSq3b6CDiyMxeUPg7xKPSmd5l0ayb4XcrdZn2RlD+TMTPaY
sNbm9GKT7HZoKXM/dYCEt9rwYJky388HjJLLVlZ1hzN7acYmepSi+NXRzTOsIz5N
ly6vkJFMRS/GdPwZUoCuhsYKMO+szH879Fcoz6rPRdCVWce7p4LP1uDrg4zg4q/U
cY8Ew8S2qV2EBJe7RPm2sPv74HwuiPLBKLeakc2tYN6mJdoFQlARe7k61/M0Axkw
dmnE+oX83A9xSHE/e0Wy0fine4XGdGR5VWWsw229qp72G2eJ16iJv07wTZfqjdSi
lAmohvQFsuVhbRmR00DiuH6m9S3wYoc0D9VAfeU0tqC/ELVb2f0r6OcZJphKSzN3
IjO3nr40NlZHK1xGuGeLQSYhZeqvKZ3UmDaSx3gJRVT1LfnTXHeBbYorO/3hBktz
lDyywpKR1vnMPcpIbJLdAlNCKN1ThqYxAKEIDFDkNv9EwL6xgX2qt8S/3L/nnWKe
ErstIF5fkMd2Be8h6akjFDXb5qzSFSr7Wtq0TX0t5zN4fADDnsRzEhhEOqsqpCLH
SjuAV/NTEuzEqvcvqYnUdktCAHVA9aDU8NLFHlwqASDy6R29/Vf7+FwayHRY4ix6
HkevNPz7jzRg8os0pHYz9kl4CreMZeY6aKXGBxz7jzM4sC5dUMyrFj6ta0auzvhJ
wnziS8CaalLkUe4YO7+FC6OukiQWB4hk3+uxm2jYGfH88Pcr+eER26S9Oe7b2Pxv
4oS1InQQn52tC7BhcWtcCZkoj/7C231EGebG27YlmJ31YHJGlnCgPiMAEsMUWYbq
PKwC2A8UoXxfmikGz7qA18FpgNDDVA9WdvIYqIoDcqbKEdejBSqxGuVRnGoGN1xB
MV7JSA0+Sc2omZ+yFj9mIgNYwsllxwoGPAV4ySGp2th3+cmdS6Q0g3L8RYjoj8My
lojFP/ZSVrmhZhNcZvBosJpZ/L6VNIKVTP0K86Byw1DuKCwJ6P+s0P2t4+x/RwB8
23u0G9aqRXExLC/Ly1bDjn1YnGW/CIx7MzO9TQsyQUkCEHq8+FbaL429TuOWRERb
E5FzCEisMW1zLghpHtR/G4Fzgbxkb33oEAWbHEjs2NJ3Df/WLCGPe9aroYZM6j4H
AzvSRfXS9jBYf94lnbbfa6trrYeDNuDqzMM7SrTZx0LIsNybdDNn6f6360+t4Y7Q
nDXNGLhv0JaGVvKg846afsSGwZrsaI7tE7Vaf2laFrpmKwLlqcKmBOCJii6E+wx+
cx0wN7Ve1coYe9ccWVw+gPkIyEyUX+I2q50gRUKHH5E+I81KXR90vkVI+0gEISRO
dGds318XDX72rb3YMLWmQ7nfytdOIXNuqkgOrUjkfz5lPIsJEEXqAqWobYZrRiru
yTJ3QNIAViisKxlmuj+w+RWahsXduii6tkcHGPjvOdtrT7VcO+JyJjGQUZIy50Xe
2WEQLZpUp6lcMBBf6RLYkC/ytRjvqs4dCFp5w+MdBnKyoMea23SMsWCRnmbNVok2
jElqIBleciKmmmgC7J6pmH5h4gLlChQ3OvK4je1JhVhf+YQAvCC8rF1Ke2WIZWAR
3mqgf/KLRiTzqtrpXh44z5EgUQhJZr3s1Q/DYqjJHZxffvJ/xnQKitnDrKSIEqU9
b3RjIgsvZ5KapcAewm4bi3/KurNfjewAINam36UP7fn0jo/V2JLYNTm4eFoEdswx
NMXEU9lQTVwBKwMA3oy0+kS/ACdh3+YpWprZGvEcHH1U+/+u+iQamI+7WUgRLsBB
3NDXNi/y6BhW/F2Z2Ghz83+fLo6IWdp0kGHm2WSYkI2gOoYr6hVRQtRN5JJGCDa6
LiRqYNWHxDX/prRZ3XwrS9ah2i3bOHow0oBL+bkv6N/KnHG675Bw7zXFJLXox8Oh
5MPP9+I4GsJmFwxKgeJVamDgVxUB9omRZehcdow/fkKHybxbsnRYJS1N/NXDmfIC
kUPpf8BmL5kYnhZstwhBMWtBVxO6POr5Ph2jQZZBCiWP7mHArvZZ+WyjS0Zgatfw
KBM4rxsx3HLxW5PFwOe+hTgbS+VsuqyaSB7/UWMc3Lns5EN0MAAd1In1tP5HCIjM
9yqnm7EP13c3eciArK2avZB40RAX39NuBmtx4j6NbmXEqutFFCrmyCtLf3bvadVV
r5OR2KNGF29tmOAr2Jm/PhXk1wWD/rdc4mu2gFDPV12oikIw0Df8n6vjBML8N16O
Eak5+YNOsTaUlL0dsRixLfOGPftyrSySXluIQhYM902/y9z8AsFdasEeaA9EE92D
PKrtSEg47o9Z0Tl9hjVoznrZqmWQo/DeB6SgXlTpMsCpLVYELf7ZUTkP6aJZZdHL
H7fFi7vQmNGk7t01S4VqHifQDk2vP16I89bkdCNAtAy3f6wvU3QPFWQ6QBSSP568
6waZxCBPnUWQyek0pkkU6Aa41U0Bi3ARNibwmcVHtk8+b7FY//fGPDKcwu8Ceo/W
ioph12QuqRCQ3+3OH7c42NkWXQuz/s2EU+TzxPbTJr+KUZCXPvoW8M/rSFHXhbG7
KCQvVQPEZdlIjkwh87r/wJqV5hPrxaRTWBAAsWgVQa9bccEF6CCOTAn1vRuhOYJB
JkuyNb6E3C8yfOf1Eg8N7jnLitDJduYSsInfn815bAWZV3hmLYwQnDVuU3hD4+CE
O/1NYaQoZ8KqxO+AqR9t/lgUxrkeeu7Ghih9WLyFteHcSR5xgaBNegEE+poSO+Dy
YRe+SDtLyQx96g2RtGbj2jmMLjpQeZVDIgpBH1I+toTlI8VXrTZwzKQwv+V2jL7x
C0+Mq0orA5Avq3EKevEMCrCR1HWPoyrslXQnpcMjAaT7f80GVhnh62afCAg6+4eO
Cb94p0pLXCSngxS4UiYSzhDUam7o42oWTxGEPCsG/KRnMyXxmqAo2dFdr+oYhBwE
SU7Qf9uS/+T9N/DLD4Krn3/doAaIjIfj1mLVhoSXG84IAxB0ymJZhirNqUccpeK0
UzPNIym9y/4CfiYgjiYBPaDdlWd71RU5GvsdSVDKH59mJ7ILQMwjyEk7I+KgMW2I
rhCJ+SLKUgryfFHTCqQVZT0gy4Qi8Rt7rZ/po77q8l75gLYTcv5iPQo8BJS91cxQ
XUVXAnCcD0gefcf/I1Fk6S3KxMnkK/Dj5P2IRvjLmVkdWv+dSc6aSZ3kZoWspZdc
IQ4zhEZftj7tdTVdVAU38Qd1S+OW1pDM7ZS6Ali/oo+fZVOIFWM3xCfXjcwArjdo
slGXgcTFa70j2hvlZO58gCKGYgf1UF/AFvrQFC+qmArhhQsxqGI0MDyEzVKlItCd
2LlVqPYW/WqE48Lf8puYkPus0aJVKOwkUG+jQyrMZu/mraCIAis9d/R/xWck6GCv
ZYpHdTgnVPvLh2O0EDdIUdNj5wr9uNYNmj0AivHvgbMkmOhgtlLJP2VI/Z1rytWX
KlMCI7rrXPZb5+HcFCkFPDgMNsuT9YEhpfqqyoKP0hK1keyTM6LWMxuD5Sy0uJnk
/5vpiRkOc6Nt5Xx7lDTqI6J0yfsd9/YqGtE9/FHAAd8XOsb/4AbP40TC3seuajQY
LItXCj+UgOJnjI2BPQ//tPpZFl5CcwujeY7WW79Iyy/wEtTiND97Y6CqBFfyGI7c
1TOl3iHj9DLF8fu5svJOvCyGhhV6nvNjqCE7lviyXX+z0N+yOcI4SUJqt9xC8m44
NGtUDaj56IUnpOQJyDADIlNhNhoCq19oxAkD4RgQuihfy0hebN/UXmqXhrN77XOi
99k5GOxCljeGKUHAcBL8FTLiWB3vAHGldpvDFZZ4ZWXXP2nJuM9DqTAI7K0bKcrc
4tIp9OUSstcqIExQH6Nq+2D10cMafqJnM51qQ+Dm16UO9bPe3OzAcpXIjptodzxJ
MNTynOmbCYvztv6F/9ImA2cm5PcA52PHN7tI9M4S9CeKMT/2HKOWVT8MxyZLBBY9
XpJt1ZHdJK9DG2UoC+tZQzfqcN59Y+Mm934r3BdxN4+8Jzo9br4zUk9Y3nLsk52r
ilt9AWmhhKWAKfg+rluWBEIYF+bvcq3TGHdhkXJitTDUboWP8JMHFKp+ydokT4Jt
Z8Ix2WoxEYDwxUVhsnpXdgKHakFoZgkRlung8UT7txBSGD/mcsCtEn56/nfuw82N
dCXYWQN0HRVDbSIv24avHJ50XNkjqFiK791Efk3xCVWUWlJw7lCgD77VYVDUYjns
axcqmd/cvT21XVS6R6Qypn8/kL6TsoTMLufbkJCpTTeHDgTIaeMj1nKWjebgRgxV
UtQnrbazOItL3uucMJ4Tcuq29zBQAdqKKiTaQhqve/UuupKp8S25bqBIQqwARBwI
gUo+IxdHVlYJSsut03a+xIF6cuk0xdi53H7itr69rBLSLr+O/VQRAEIH/PybyxE/
yUUYe36m8P7sntNywvtyqXGqWu2ZAayQVMgJ3RADjX/mosujp8yP0q2Tv+I9TndD
fwpxcZiD/9GVYeqGp0cY4C0ZeRKmSiEc7yNWNXI6YbI5wuUSkHH47ZRFRmBeNCXR
qeiKUj6OV9Eljwkh7+NUb8fu/+Gc8uzqBwdNQiqrQuilH5MV2/QbIJBUk7TlOGTB
QYQ3q6U8XiHAagsLwHXQr0yPmxevyTLNpwzaoWIAJxkgeU+wKKX17fqsAdL7Qdyc
XyCX/ANV/AHaqfBntV0AUn3KMwmaZIsXyXxU4qAn0Rs7T/iQqxgPgJ/qemu+zJpR
Uv1r+rwqTMNVlDP2bZt0CnMPA3L0KIZlAHfgW6MB80VkqljxtEqYVMlqT+Ixe/Au
Xk3aCmaM83MbEygpXQK8XY4suRVUNNoy1LhnLlaygbb3eWj85buDWqqsi7kwO1gQ
+nsXDtCJM7olgajUnbVm9TSuHiZ9DGI0UMWbaOlXivvVrJpM4abFGwAj5j6tzJUT
rf0UNMhYNnwlgecay0zkqQIbrkUub8L8QUkM9pSKpX5Jaz0GW9xTL8CXQAxalS5P
nQXKhO1syxlRG0ua3pZ9/WcyEzVThrZbngHyLTNWVtnFOHdVemuY2+4zFs/LyFoj
Y5ZDNpS9+BArl2wys8Allv3F2qWNCaBTC2qq5APgsyEqw5FsMYOeVoWQjztW3Gbz
n/QwDhOnoXATkAqaF2m5bxeBSiqypi3edxwZGZeVxud5eWQY1AuvrJEPQgo/1jpG
EablAMTILlpZ+6o8vqos4SUaWnnpzLfWOlslv8y8N9f72iumyQHeNO1NUG0d8X3m
Tn3DaEjvC9/DTkjYJl6FC0VrcBRx2TYoEPkdb1cEP6fb//8KtLdxAbjeRafXIh/j
0S9bhq8YX94rljph3GhgYQBUb8cvb4vj6iKnifPfexJVIZzD/EKEpwHNxsKlz5VK
/Tlt0of1ca+/OoMOKZjEtDEkFe94JFZxmM8cCfw4a3/2uB/LYME8ycVx6WCSu+Yw
N/l2F0x1vQLXCbLeXJmAqpuzrfP5yKD+AL5q7/ckrBHDGKyiAz16sILFM+0r5ZSs
oZHdXMuPsOKhbBb37ziIVZ9KyHIe5FE7e/fwAMiyC4QvEvrwNatEsEVS2iUUsz1E
FiljgpIhjNCK24wLJ7ZLnfOnT2AW8ZxIHJ8/nEL2JiWb8oh5mu0zqMjn45Vtu59f
Yx7GsuXa0N6UnYOyNmSTFvL53YJaiPso9qPhqI5GCSIQtHODfwQVvYzWHudzUyTh
tuEwnijXw3K/REJHhSYWugSX4QXpSyVvQUdirfly1P8pt/v5qsFxZsHGNDCD7SPC
RBy5gswuiTBikagp0Bp6tMMrNoxXidBMyTEiOA54ywjjuFPs1ID2706I98sKuivV
ojUUHNGoveQ4y3wpW7E0SV44O3caZ4e0Nvijq3P7JgdPNMaMgAtOsVreT5JtwsaM
wrcMMKlVlieKmgRa6Zdhj70L8ogvP4PC3nX5sHjrvwcA23ImW8kbvNa3KtMOfQpi
LM2ZhQbCxC9yyhmxu7tRWP8rPVDWDVm6pQ8ij1BNphRs3RbuPvbcViN89tXsbfvO
N3zgWjnJ8g/r8urIClHj7lJHFrC4oXHPxjNJVO49iGr0yrYVIYVoCtEgC16/kt81
8e3ovl2VYk4m6OTnfpUbad3/11/OQt+fb9mDTa6K30BM/fIehmDrAT4Hhd0rZd7g
pNv4o4+nJ3/TZCCvnwMhIDbX5z2c5E8AICMlsTAdYZhAvVy3eSg/MqaYg/27cisN
F9s/JNiq7ducW5hxOWG8RrKgqfG1TbXTSBaEvIH+0WcyBJ0PKAVSXn/EyaIEm17x
mB88/U0ZxeUN9M9ISSGzfl3LTSliXBq8VkTIOLcIKK6a9tVZ6oo5bo0CFcym8HVH
RpWytJQN8mlwiuLDIAc3QqBK4yGvGVGMcLtJrfh/xxJmxyMQskCLQUpu7C4vNzoK
ASOQ7R/gTKoKbkcgNb7+mOm4HL/nexihVvdEaCXMRJtFfxkjY7yU+P9LZ5fO8hpa
qyzWA7dGyKSaljgWhPeJ1q8FHiLhjmkG+MNXzDy4HGjC2V70DLd33osWluW323Kc
sCP4SQnasbV82B2gliCvd/RVVpRPoljdF1bA+T9knORQ+g9GgvulJMePUdnOIQR9
OTb/omRidcD8bNQowBaFuUDT6lKPnG9x+YOZVDxtzDhmuvhHNBxr7g01BOmMui3+
XTo+oL/UfgvAuxFSww3FsJfK8fWzlniozAKYyo2l6nXinlk+an3Om+Nc5pOhEiR3
P3ExBoNyTKvJDaPIo7YMBQ5a6tbIaGc08PvNlAsQ+fIz79uv5cQQFQulzBiY6F1M
V697LD6C517ZrwcqcSNT2/+BtbrYAHQ0QyxCKP3XV4cKqtrmIisw8TYbbHDzLPJF
cpzlTzOGS0V6v/iRHQZGBnDap94HRBTbHFDW04KRvkvfSAZ5heetA4/RgHtL7un1
m25f68Exp2ZrTzPVG6fvmgS77argZsFq+XE1+zczX7ghdI/woD0eT5LAYqKtYzux
uFUkgvkUvC36bV+ei37l7EEFrM2/gv1J7VU0uATx2OAhynw/6lv5VMQCLmyMk/06
/JoMtWz8X29N+8Dg/unsshpBqqHny7E1PPSn4TKdaVmmjswJwkjY9KX61gQSP3rI
J9RVA6rjaaHzgQV7p0YoT7EsG+n6V8hLAu9nWxdYSU782dZuYB4fUi7S+UivTMZA
K0vFgyi+Mcqp40FPqjFochEcwspILSMzoDHORVvcqKjsTgtzWme5nA/qaQsfKVvA
OnEvxzSgvOBKckV6qjrT9k3oj0zrlzsGJp2Gks4tvauIlKmxr3ttH2bN4l0Lo9gt
i66aGAoBuZKi36ZcqMMACXtEQ6MMzBeVvmhVfzoU4UVSlmrzNcMAcEAY1CX58m2f
zzAFn3lKRlm08y7yTeG9pBryMSxMXBw52WCa7tLif9Xi4r6r4YwGvrZyEoxy8ipV
Pn9oDVFpbIwzn+E4e0XDQu1KpVDjjgGGtG/Ex5iA29Rp6/u7BbZ89dPIeHI+ZXa+
KQqTMsXpmhyJqT2H4Pd1MYmxk0gbaK1p/VO4W3oQIEN/zuqnplqSr1WLcLtcEofs
IqPul0lTkSAxYDvG9O+5K84jsDcF0g96AAk9gzShGmt9xiPDCDDoBeKK3S1atOqW
h+sbYrZfQc8fDr/NONM3F7lX+qAYU0kUyFSsMmXIUtawlPjId++r+jm9245eMuNQ
2czyQSvi6CNOT4Kig/mzbaNHOpjGfyP0CIvd1ZYJITkZOGyOIOBkpX+sJc9ITOpC
u3vUxpIMBoy7TYL3VB4FOJW8jLi3Y38tpPHYc+GEhVYoWMlRVuAS7lbI4OvDvxrl
N4slhkQc/FqCj3UmyhFaq2siv3rM0ogBZjb+cmWW/xnAvahhO63SPVCCQ2KRK+iO
amZ0wICdx2e99hF+YdeAwjA7H1eKCKX/0C6ebok+atX/GRDabOT0CAW02ZB2LIJj
4iFuMipNayrGtbYKDUOQGhzYWbnXxcNOMUqlp7K4V2jjQXZPp40nDqUs4PnQJEQC
KuQBJA82aAg3teniA5PL9nSqphhB+albbEDvQQIhzghCJvW7Gc0gr1XVuJvlmsSi
udJpbX+VjWQY792XCyqV7cc8eCG1p5Ho5yyF8PjGxg5NjkTtbJZ4jHJax+BfQfGP
V977/ZU+XuviRPqGLZjG8sYaG0zstRU4Fen6dQdnk4l8+RHXdxXE1o6hBpyQVWFg
SFJyvJh0H+kOuUrBTto1DXtfIJJzihGKrYDpLynnqFCfNWg0/3BQEZWX+hWXT6lN
3bUXB7CZdDhkR0erju9bfHyP6cadCD6Td4BXeSbZ7yYWxU4pzKcThZ2hySHO2peQ
g+UTXvCtYOmIU474i8qjo73jJmZi9/oc0snUTsTaCylsqLbEfVVLU+VYnRabk6VD
UXzkERWGC3mVMH0R54yab2FuuSz1Ip/N2Q3rRIDINYKsUQqoguGFzeqYvWIRHpWO
PahksIljwdkF1rYvCIHHQKBlZ7TX9QWmVfKMl4MLeQSwC8jKS5K9lfirQoFfKu3S
mStjbZzNkMZcKnWd1Co52gZJTRnYWU0VhpQYpid1J/txAmAZBaAhWdA6U5eJqq4g
vgoqTlL0qVIJKYgrJXlGaBqpprvwQsnczjfNOTKdRQgvK7W93srLBDrVwwMf+Zo3
RoO6im3VYEn5QQEx9q4Q/DPQx2LqEds0efXJn2Tbd4Jmo7vl8CtoV+aX/jsF94Gl
Rg9eiBr/W8BTAtO/xvMQgCXeQhHoTHPqnqtTNNAsQD8YcOcqMeIMch0CkiCRG1EE
tjga+nJOlQft5c+lFbsMMSb0IbG5iFDmHytAhXZ9cVIi1IcynkpwKF5FPDKIARZH
fYLiFxx/xo+q56Fsjdwd3xByITD2Am+GLVyzVk2gBXESrBaSkxeHamBmQcc0esIK
OlTrzjgOzK2hjxknIGrpE5fG549hFsH/JyhoFAzcezoJ/ht8gmp7yODleZRdVkVv
VIMvedW0gX47dWRMJblyrHVhwIZOg/MquKvboq8C0kPNvbpnj8d0TTQkIO8QyxXU
yheYB2cKVRI0B1KB3ZodNtn3IrBkC5xFiptsdr2Fys8WT3n//azSNzRuNgmpW36Z
ra8tt13IEFj6PLRky5ES8HYAF/65N87b87O5A0EujBED52zp7Hzg0Os1d1nB60/6
cEF8KscTM4VM07mN8ai5Dbl2dtKbuDoVl+pi1efgPMJjtxL0OVOcyix9hMNFDNSc
rvCZ67oI5fm/CqUTkg7nL4o7kPSk7qsz6TOF3bE+QInw4y4bDtdG+C/kP1trAXAJ
sOpbY2gCJ66XXiBxFbJXXS75+gNQTcrrmq+X/tATCIlZPXPG2t0lb74QaVClJskR
Rk4MSIKyGO/4y4PBGSwXcJ0EhN9tT8YTUKcI+wvw85aLwvVL/bFQ0zuZta42qQ8k
S4Aqbgu7+mTXE9CL/W+065yi/7eR817xc33I39yxPwfyXd0YYF589+HaJ24xaNYF
0KewLEDLeUut9OhOir+SZG+dlW/gsTHt2KEr36h3zAdTFBDXo78LLQEeo/z3LKqB
IGf8ZfJSW7ja+MqGw/ily67fq7XafZp287QHkw7opdf0pq1htxWNYw5SRtJyZUPm
SbFV6N3ZFdTRoFb7DPn0sqR3z731iv91BKd3bRAFDOVehziNDBCdCmlghqG2Q6od
eY15zAw1KdmMav3fiwblitJsEGfUEC9mQvRH/CdgQSyfAjwUI/O037NdN9l9eA1F
9O/QuM0hvNlr2baNSmRQn8seDOXQoNK885fkttZKWWV72eeURSQmZD7BuMLg151t
S6tBhx/KFXHhEj/X3ffILCryZmA+wCDlR9GOkfE0fBn22HAb+WaAsSGUpLJI3vAF
GMVUN4C4M9LQ5avm7zbS1gXRc2luWRTQbL+v2C4+sTJ+cZgPq9Ws0Q3E6Grh6+mQ
mWAiib+5nWeZL7+s2BRkYTddsCE3LdN9T1CRCcOcdzVMfwgM4fFGro/gcuChjSVR
kIsrzoPVQphH60aZWSAJLAW4By8is2f/6tiJ/+4Fhr1wCQH1xnfDnDuwo3yZZei7
HeLxC6W80cwurKjG52s75/QgoIRqug8x39K4WwE0ew+0unZ37Lc9VxweUJU86PPp
talknoFLj0kUEAeTf9z1yoZiF23VOLm4e4V7RE4NsiW0rCm8ceD586rhgPiwIfuB
fyDSWz6Nqy0wNQZZDhc+5R/Q4jtcAPeEFb2DS1Au3T6L+y/r2yIfSWDHw4zDJilF
nytKAUMwu4la8zsVt4nkkzyKocegU3es3NhqnbUa3KUmdZZVP6LHatIzZm7wW8+b
oU1MQ+uGmsdnWmATTVtQxDusCHwqBQSr5+kg+f9hUkNIjFFl+IzS5v+ZNzyGfTlj
UguahUR5Gg8gu1qO+C0B5FxNyO/FOt7Lg8oeGbGrXfyqxoB6XfbrXsZBoY/WpXt6
oCH0fHoIqoVJQxr907sR4mYs6x59ffh/c+Wfn8P3wL+B333wwwZ3cW6D7ysdgxwF
s+kUH07XGgcMqY5Y+/GZ78j+hC1j5l/E2SmKxRRhblZJNuDCxQTHkcA+sxjJko2v
0oPMmQ/SAzHEEX94/Mv7ktP7MNZ/V3/kk5+ooBRs1qnZDMhELViyl18k2AtyIFoN
iOgHS+2TrxRDKmQ7CaFIFcvduv4MnzrjS61dBbn1GHnviH6Af879GU+dnPxvYSoj
gVq2iT6ru1jLXfKMOTfXOhns8S9xM5hQp9PY0t6kbi5hEd9AfAlxIKRHSribaGWo
JeehJCuTrlSCKqBsqjZrd1QrYEml2wkGgXuX7oXJLOxkzaO+BmXKqu1m0POXzOFe
5P9rwwE+jKbfpxIGRJvuPVjssw8nKFWWpw6P0AjrdpqmHgsE9clT5QsL9lnTXlao
0u+pZKLyE6VXvj7gqbMq97oImcyplKjWhKflZaLJ8RnaU8JlBECZidx+q/giC/ym
lWUI5o2ai4Nw0kKK3TftGSovDLBsWhUXULorbJU2ZCZrVPkwSDahVlfM1f2vB6Ff
3RG+1vpafq1FrxKhsY/Cnxsnjnr7Bj5dcqKEiTV66esXFmvU5N/iNuIX7n7nioIR
g1Sn/WOq1lI2+ME8jqb03iuP7DizgQbD8hc17lOsMbnJUeQ6KdacUqTg3yCjV71o
ixtC6N87ka4m8vA5Aay4UI/1iVDvuhTVltiiBkylJQ1tGTB4ReOikcjRq+MvvGhV
n4CkurtIz5tUoLL7keZhJb6McD0oQStxcq23dMRJHBIZ372+u7+z/vpTNydXhlls
Lr1HYiE0hEAhwX7tUyyTRblptaHyIvE5yIUiTz5vo2F8jCdBOQBTgzqOUWj06YqZ
M8Cg0o/5xi0tfX1kjsuoYLXHaC7BI3hjovVzs7PXZEkvcpqDPZadfurVC1onc7qD
z3dmMKYXfAxNE6u9OuKv61iL7aWtqiqTA8cNhQ5B14FHxPEMros3NJrEkMtrVwdw
r0SrGaxh/rL3ggQQ3XQ6zQJALfXXu3AUrsEi2iWeHVjGjQ+OXG+nFidgsN8JIWhq
t/+MuURIOTw3/NIjSG2QeYLVOfeVwu91nBzU/YQ/RsunfNXgoxCx65AYDLi29Ymr
7zeUDCPvHDG1gw4CWD+ExGlpBH/o+X8cxhwoxFarXDmhFkdTKiYqoBZ+nPvzWr7+
ddNW0HcsHKTCazIYZkua5KxM0uJeC59wxS8pCQK0fRPcMQQd/WL0xGPvv02DwZro
acrwl+ov+2BwpgjCtDisjdMjOSSZq9obgFcOfPFVbG5UuweXJHHLl33u41B2FlP3
KyzRznZVyknTmdc1GBA4SUmRllhfiRe7dGBG9w4Coftxy5EqmMSl5fBFyMlyGiFM
iQRz/bRnuT+CvPDmmkERzHTpalrXf6m/BEwfiVwfipmEFPOLwZhmDIsoNXlOiDgd
iwm47HU1++PuC57/KqjmcV++aqOdyYhh/12WRCA8cANby1zNXAhpZ+Zm6py50ICU
ZrslV6gI4fFVsRIsiYDeAlTKIQK3liJCqz8rEO2Mfn2dS+hGJMjFgirAmsxaHzG/
IvzvstCMKbztn8NiyZ4n63HCNgE1bYh+IDYT45VinJpcwLyUGOYmVT8fHT+8SKty
vy1yN+W5m56P7fkJ6K4vRtkmTXvs1owCXTBaSnyGf0PdwS9youCFQOqMDx5aA8Nx
5JbX+bUN5kKPevIny8SC5q6oXBrt5+v2A7hgL3eWDpObTwBITVVGj2gigsh2VEHs
2EHkTvG2xr3+LDWin4sJ6jdbf4ZvqRUfOEYbWxZ/v/EaTQC2olueW/4oLMbd6yXQ
Av7NrqjbsHgjTvbh5FvECC0e0ZX2ZjLJUaXTK1BYbfzbuj3Q5/aC/FV7rqMR3UgM
L46WBAFovk4WWyw5oTQVGMZbEjZ1z4OglQptqzl8ltOKG3eUlTfMY2Acj4XRhpbC
7ip7gx9ZJuDQxziRVQZq3Pq7pfZhBwvIYepFL3f7csC70JdIiqqXtrHEr9ILyLRp
04CsQrc4CYBbT4cSxONR075yfj8NgmfzcDvxySmLMSNkkaOyIwy/gU628n10BD48
Jldrs6Uwn4mHEtItnxI8FfxTeCXmtlkmjamm8nv/KZ/P6sgTVKeAGEYTnqLB5A2k
UeonLH7P+gSmy28PQ4yDXj/wThwqfSmfvnXimFOPfykXO84V8GSx0nTM+66M8n9n
+zJO+Uw1UsGdKxjTO+Uhoj/z45o0Bw7+8yePuh8Bjf4IOXsjC+TnkiilqKU7EDRV
vnObCamAVu2Hp+/jz9E9HlzFQgFemP2ALjGLUkpXWypkhabL2/0vmhUNnailOYEj
9H5MDt4K6VzKIe+jNnTY2Q9VMDtrJmlwcEv6PBohez+PrxT3V3uQLUrur5HNvKzU
+Pa0Ck6tDQBgY+GwPc6+Dk43rBgQH34FdtUbEnNqKuC5YKrgUrTLqyZjQ2zUEzna
vgI4KSf7ABGuYyYyktbNi4/YKb3LGZdz1uS1hlkA5iMlrdkFF6jpqKqV213P2Tvy
LiWLsaxjKOPu9M4KiU330Tb4iYX4UmamM1BVK07iloH088Abx5MNqcPie3FR9eRi
9YGgi7jOmOhKnH/dAhWPutaYc0g3CKsTe0n4qID8/9qAr5wT0/NPmAxSmkKnaC29
w+FFfe5eUUnUjZRi6/W8o6uN4yTaVCOxFMdUf98+WgSr3TGBI1eNkZAJnaT0Ur+2
dI57co3NPAf3jDbqSb0zGVr/GG5YnSV2kBkgLOr5cr1z7vJdN5CtTEJvX9Oe5wTU
OGhBrx+gtYarthwPwaLo6YUM74nnJYsqO52qQx+W8iBFe4ltansL/O4Tx/Jp3gLF
mzVQj2Tauyav/9xR2/kD//T9qb/2b4EJqbR5YF8ypWZYzO/W3dik0EqGmfNS0MiW
WFwLJhnTFTBPuMloVvu/DAWADn0eoS5QWEnvZ7HmEQjYA8pCsaWeZ7gzWjriSObE
QG2z1r+NWz4pE3G1NtNWKaBeucFxG8ALggw2AOJGCf71ukKLOX7Gdo6Zmr1ZJiTm
HBwICBhz23IAr3b0x4FcB9jI6p1FZgAF0aROtA5bjU2zcEJFaDHqAZUtrskUNatY
9nwfWKejwSs3r+qvMHnOUKjPHbmAWmjTcizRvXSETx06EHYYrp0jk0gldcAlr1F4
64xy0xyTD+XrBrYC2YiZpVgS5WCC3Twhyg5sLsa/tvRKI4+za34REU26qOyUHH81
XOt2zY5QwoQ45w2kGpEyUfcTTYjFOu7NFG64cwbnodbc9zGZ9av3ZzFG7l3cq/+r
h5njxgH9r2DOtdHOATb8fO/y2/2eeG3m+INMk8GSVsVG7WZj40BuueDJaufZkeRo
pCMvUahkTqUdE2xstKWifdd24AgDeG+dX5yMlcLGYlMu59smk7bvertdzXW2Tapk
PkIOOARj77ehtqcXWjaKQ6c/dYKbAnKPISOUotVdlCr4zcnvkKO3TdVoyHFemhe+
xmG+aEj8zW+08XP0Gh4zRscMKR2omWNbjNhhadw3n/XaorXjFV44AuTVwpy+ldzl
mLcgMlKeSqFimlhEg+IGp4ywmhKKG939BpglY8jl4nNe72r1T0agSF8ATN4xpeI+
w4lLQ9d3fGRfUyLt0guNsrPxXkFsxpd1LQ8uiQw0OmGuROW9MElcy/HL7ruq6GmT
fDsMYpyn2/24MkQ8qq8royfyf5Cx3KcVKrGXsTlZJxNyzyx1JmqKIZY2eqUOLs7E
re6m4XWdBkzHBi6M1DdyMClWrd3+lA3Se09m3zKRk6EImzQqtXQGVa/bqOGgcC3c
DuDZUnuRV+vdHYwXdLVowZSEkEtmTlMUxW51HUEH+cAIiSM2hEPBwgudNVmKveVX
uZYmjIGQR6k9AYzUMDwwsQdg2mUGZ/0hLr38eKR/v/HHZ2kSGQjWt69iEpAHwk7C
DSPfwaKnaLH3X5WeKgQ9KdX3MslCHSHlNuPM1DXC7xQEmeSip7P47Cuvhb1ZWyru
FyKzcaQNhwXIbfjz9vHPt6OtYnFYitdTRaU/qaIsf8ZnnBaNoSt+XuiBDykh9PhT
bYOc8Io7P8Kc1GpGUZsmJdZz3ibgORMzlvya95jsKACyWRpd49k9Idf8I+j5dYjW
tu2PmBdTqDTrEUxGHj6nVDdxIoKOEuXzzYWePxN9ItofRFahuyGYe038BhAwKu6+
PnA19CMA9IVupyOvQxa9n1luf+39133kcaDUO7rrRq0wdTIPrC80i2DA2v9blSfg
sFhTmTQrb0G7knI4Vp5qXBfLYW6BelRi2/xDf5D/dlwh0K097L71bEGoVw9dCnsL
Ns+nV0NMfS2USP+xjY1Ks03UuDhrZsvydlcB8aKVW/QcSdZ4Duregs8Hx1p5TRF/
eoft3MtBSJZ3m2S3eB9D4l6PvH/20m+txrDdt9Xblec54hlPxBwB0Z3ARnFPQ/iV
fjx3FZVuKWhDaUgM/EwzqF8MGnNtO8riW18x8IxJxwy6T7SGNj+5wegq8klLKFwH
Yre3Vho+InXJsGcIXQJGR4JwOY8YmgMjvNxAXIPPQeG5WSMMFQKjbhJ0Q/tq/0Na
bFCRYQHt+6oEUBwAyMJ1p6FpCsS91OJUj4xfbojKFCoqgZSiYhiWjZmonHBHoMM1
QNNvJMswGl8cbRg25yHnMQ0fobuGX+Xqx1MaYaHsUAAVbvDu47UNU0g+xGh/OwWY
vTdt1IW0bHLGy6ha67I1kgaxwCDJPd4lwE6ZqkydGpJMM191IQIui/Z4/fPUSGxr
OIFJyIvQgr6Z9F7Q1+5n39ZnOEPuXTQ0P/RRfhjvxQt9HrT2rfIpibGH7hWv7Twl
jyzh6cQ5p31ZpxTStuR+KVnfQ+BhbaEsVH6k7slB/rbdnHJbT7FqSxyPAKdMIjkI
mkUnwQkLq5SfBkeQjAlpRpRbntzmpfuy46ZimdNalRdC8yjH1F+qQ+hO6zl+T8RM
UESuOuS60OYVfFMA7Uh0tdECrtRbbepnfdDA2i2Si2N1UYXqJPRt9J5zkXoFsCn1
Ka4luca7VqaF9F7at8fZoyOQXUke+6HG+xqrdJBqHhm/gIE25667OdHfe3sFoGSz
e41zhwI2Mdkclgescm0iqkQ30/4V7/gc15WhuDeYW5iy7Hze5JdvLJP6XNtcouXj
/1QRr0FzDXhCTV+5Fq2HeH5xfn2qo44dbQb3TDM6oKDZxdvL7QUmdGQtSuDl9WR3
z27yFcwHWOi63epg/Q44X7l5nkm5rpFFtY9FiSc8XV2ubgzvE0HOGaDpuT2QN8bY
k7p0WdMWBcAoZl2dldSADCP9kI88d+bNnKI1257exBkHYUMpB/jJdgeb24Vs/o0D
OW5otm7X2MsAeJIFIGksM1o96Vkv5ycId9IEsovhGAub3r+NTfRQ7aBrLl1b2lY/
m88NtwN80aCs/OXH2K2xYbmKvZUMmiafZKhvGgw1EPUFDy5z7EKE0sIkA744LItM
b8QXdwAuvyzjGC6XnZ4128/C9kd/2ua5Hp40Tb296VR/Stx/3Jra/ShIQ0btQMl8
8/InXRUQEL/xIhgm1drXW8eo8gYERr4rC+SqihFMIyCFAEQOT63Mlgn9sfh46BYc
4z4ZPOOA8d9h3WuD1CXCVg3fvN+mZVp75aX2k0pXwhN2XCb0je2KJKHg9eX9qHJ/
SzrcRquAePPyN6AzUMM7E7hqG6qNRso53wB+Pr2rXvyAZ0aMjtSyXmlTHSkKzks1
h4ibQww0Iar1T15M/aDpArEsYLRiv4NkE9lW/X6TP2nJpLBIY6swgCZIbarD2gOd
fQeo66C2XkIB2o/7/9ox/4bcAdyAR6FkHuPrBgzuZc7t69oL2Ux0ynsbSWsxYliB
J9o38RhntBwik65tWdiV4RDf7Y3iS0w5cAgnYU3TKI+QxfgtbvqChWG0Yi+svKH4
nxPMXMuVK4KpYrCYpA6ma71aTjPp4OjFTz8aTcyIcrQsPpeisrB6D8w8yDSe4D38
79TWU1mm6XI6ASo59Z4KmMwjRZSjpMRuBzY6KP8lJIoF7CTLa4UZ8/npQlawtpSQ
J8VGlGvcmxvIcssxBTXIei50AvOEKPT1ybFNBaHy+1Mz8aszmr2drowqnS2b3Ltx
6haakpmRvJzRTCRzn7p/UNWbci5+jQ/rcGdCp1fbPAiOzcc+T9YD8nNnrX+xJ8El
2soDX2xchN7dSvI7Cy0mJcfcgBtn8WasmsFxC7FfgYhKErCsJr236iJUIgTDovaq
mTtidpSQDvAINm5F2PVNuTvNJGYY0Tx/YG+P1fHxAfLj0VGGSt8s/+MUbjwqqTeZ
kUwyGzS9A7M4YR9llbikFlrYhO0s5gdMNLT08CrkHBwhJKw4UUNpQVumDAw/zYCj
iomB+5OqVLrAeJ9Pfg4w9I94xXffPq8dKDlftlE2leTWF3Az2V/UEnR1coEqzG40
OsA8B56oiUq18zcEgROKIlCNo/I/aidNpqKjQLlh00DqlVxsEMtq5UobiQOFT7US
8/UB588GvGUGJXdlsdHaRKp5EctDPRcn4vOHgV5BfCZgpUAXqBjtQLINWiLXHG0y
7Yw9x0lJx6BTF5R034fNs5mM4cTR949+4smla2OhEYZai0M5IR+BE+eK5UUG+pUy
rnZWBjiD9robKlJ84lhH+56wyb8Zb+7I7AhZSd4P84tSzYGII+uETbTtP9VPEwV8
qcQPspS7fvFEsNgj0uyDY6AF932LgCPZdEi1MBjXR2KvUpPxEU1KYb1W4tlIyKuc
Qxb6lfgd2QLHNjLhF12emmJctZQKtc0JbMiF0t3sha10zFYGz2FJeVzGAqWQErtO
N/HQcfqyenO8f3LnkFqey97p32+c7gsil1rX7oK2SeAFdJrSUhxddM+lX5Wp1EaT
vMpV0+dG9sEEapmuUcxJYnHuCLYdd/RwZxYOpS26ETYt9AZJwsHrIPjbyBQldQDT
+BlF6CUqg9al+3MLJFuVTUJykE3GfR/pNJXdQuQJDbo94lzOJ3OJ8nbnVvoArrWI
e4OJnxx6KP6eU06ZXhr1EYz8Dkncyz7rDHztU1tges4Wt6Xn8ruNaF5zEgMua9/j
/6tgH/0JUOZpikfuXaumiTUy91nq/s59rIalzWhCl0KwfeGIW1Ih7ng50L7tAI93
Z1DkR7Upz28ky9bjmyw+YMUw0QXqT6XaNf8trp8sIh01zCESi6bEqbiLeW2QqNYv
VbCO8xPITP96TPMZQixLe1BbGp2q5+2VE6nDxzmMoU0kI/xtJlUw2a5R92Z6smVP
ZYKdUsqhGWZicPKt88vH2gzhRGnDShIRoDrNlVHkiKlg59l7pMDxI7mvs0grIzMg
sz2MVjrGkEmvcrKgWuKgsrW0KU16sQ/qZwxmqkp1qFw+rHl/ZKgj9bpVswf3a/ke
sJRtbHio9TnO3pYd+DIK9wZ5FYeZ205bQmykzuGia9hDtxH1y5lW5R2nwpNe8O6Q
JQ3H6wUTKeU8tzUz35fr1FxcAfqgq+l/vrmrlaOIaLNJSYFAvY2uqEjvv9WA1C6O
anjjQNlveoPAXqHJP48tltgQuCbQuKmWthx8gAM4qPovMv+Kf2u+rwgu2w4L+J3X
vGNE9UTb1+eQWqX49lmIMhKZ9MNr/5cr0BB+RDeXBtZsW69bddKko+MZgxb0jD6F
ujkmeYZcgL+DWuBsbRg7NIJU0nMd4rE/h247IaJepL94vCeZ81/Iwfhi1VpJF+OM
E/M4qlAbfkzIiPvOQ2OGeBntkTG8OemiVPSInxO/s7qq4Ni+KXQNG087t7X3Adgd
TBE1QzjqvLWUi+xpLH8SpRrsmKAq9WKoFb9Jw/He2OyUMNP+9sjxs7pHD3/p3qVr
dFllDyjl48rF+D2EMIUiigC9aSm6nR81qu7OTpae4zRbgTSPs8Dw1tB5GmTzR3uW
KwBtNp2sTHoqy5ZxHOMMAri2OrKaHIw4lGvEMUbg4OvjU2DN5QpEhfO/sXerSFnB
izNh9xYqY8Pk/0XTchsTDHG1zEbF1WhHmvhqyxdelysIMlNAICOKJVPScSXmrQID
exLW5LKrTaOFPKucWWxbcp7d8XR1mz1X+s6HPEAvbqKjp0wzW4x6+zoUzOZr7MUj
5nfg/WLYO9CzhDM0YU6oA0WAELki3A8fPzpmdSxG/xms7AoPz7Au1ias83/7e/WL
grreAP0uuV+oFi5jAkGLuhRVc+1iDNXiC4Bz75ln7CwsLPUyFzchyAOyEVxAk0zJ
+yOqPNCh9bc1vCnAxuup1QWaQwx5DxGEEq0oyh1ZiE51nTccRqL0NzwaouMgpCI0
FbJpRdRLdrdRjUhDXmK/zwA0+7jGvYaOVRZJmJsHQ04/wJHBsRn+/L0KYhB8fDy9
f41dlpQ+3MF8Z98rydt/NNlnIE6JbK6eLGDdukPdAfwu1bQVtSQsHGLd0Xibhpm4
KC6DwyekL+YbMwXNOIbHLbbGUPCY36UamwpYNzbg3y534IbkLa9kYyyo79KnS3Oh
PxCG0B1AODyk5QKch5mFJU28qKoJMCDJRNBp+eEpy9/kNlwHv4A++oQ5dTFAjMhH
fuGJvKm7uk9cEX44qwd8+ywyZOGwsGyTxNpBKCp+s3bStVF+hBghKdHJ+pL3kXjN
soRpLwEDiOIvgvBVRYT8iuDE/bJWgZxj+dYyBeEGYTzHbp6gYJRoCexqL6GBuuCH
xFvH6Y8ykKhCLxB9qIPAGHENsp/1KfQbCvkvkEkZDYLeMgUTcXBdjgOoFJWOkAdC
Y8ME7PLouLMH7QlkAhtr/9RjkEdgOkCZIH1IKqrgpyK9Zi4AAyJaNCGCZRwV+40x
14dAMh7Dd4GGI6TjVMuRfiAKopGI0qEILgKh66otaUKLrBB3URhkDTNzhtGFiIfd
lt9r04hImsISCUXfQ/IKLUnMOnX5lkNB94Lfhelz/bUmQJCU0CXkcy4BtL11gQ5/
H6jG4WYSwerZxg+Kc/9Fwfd3/l8/iQ17v4tb1i/fWGx/z1So5hO0++lzawdEcQNu
E56LORO/Hn8BtHZ4O6ZSaIzHwGoXCwCOMzKo/44kGSMCtN+qFXlG1KyWSjPPt+/P
JsBWNptGRk0uylgwFbrc7WfwsUp/vUAUYU42DvmuHboXPOyxrVFeUIrD0Bo59nJP
+4mPTT7/zEXINRK9R9NhGKLiDcWpZE8M5sno0cfrCZ6BMwJVMC9WRGzbJR0x1f28
UiVIO6uJqwEFHO1lR9Fy5L5ov1m9gfCtW1iXwpe/x5vdJO4nPaDEPwJtprgnC1XN
B9T0FMK8Ym+o8hiM3HmRugTdLPElI6gmq+u1jLyWJLjS5kKY9vw9RFOeOVA1k+Yw
um2LDqZ1ltBuShHXZs8+4oM1Fij4lQ6N4WC/bZPXeuHhLEF9i/j1Ol8aabafRHw7
INlAbTojd9SYvX7Aixwe2hKwmT1RI2XGDTHCBujqLcUosG4mslAiYx2Xg8myVDTR
XmazJH2aeutRGgBAbpOwbU6tmJzxXk1EexgIMmiD4scXSzek/uxd+jF4plAzk6WU
wfXZq4WRY5stif/3zeDNHLXjgREinjE3bEtcr27W/wO2HwXoBhUWf3WiDRMvmH9Z
qgbAuUP/vhMqT7xMRNH9HDGgrdVwWXe+C4yxgAnxvW1DrBp+DpjHr9lrKfWeTdnS
cScx0335TlmHQRGY4cn9qs80WznLLo0BaVywGRH7pGq/h2LmMfW+YJbyZTeSWJ1k
GfPW9HZ4QAKJ8oZOibJJSRRthFBv3OYPdPkekBXRW8ybjGxEsqedokDRymKYBb8p
Jq9D//EtkO18eS/l2tuSWOw8TQhABZJYvPzUN7MWlMoDf2x1bzcXYJ/raKDHUUO0
PWd7nAAj6oDZX4j0HRMhYyuJDqYxS74Nc5vY9NS12OqQh6KQl7ndkrwoqXW7BoB7
2mCu0p3tFfpcX0muyxFmCGITCOYM9tA7hpqryii3HZCDAH4Tq7v+S9xfRjESCzaC
CUjILzNxW/B7T4mtikRLjIRC9gm+XD4EzAhyvF0hC85WkfITB2xL56ul8toOv4PP
J1GOULvikxdQEINMFfyazOKE8WhWSbTfxNp4WRMujX+fKb0bToNkyjzlPOo2+TkJ
c5BJhhhS1/zPnmeHBS7WmBPxjeVNWpvSJpLNI/VJOVbo8pYWIedFwIAibleZdI6W
5x0otbLTb/wUmCWoK/uTtX3Q4hTNS2++ytjOGrafF80/OcZsGhPJlrMPzJ5Ks0Jq
AObJdzKpU6CVJeavw1s5DoQ+yv27FUOJaPjpyQ+r6IWx6HIglzqwROcxtOh500Yo
lOYOBEgKuC3QG66HnTyqO7hPDHyyDK9Q+knGUGCchi0TUCMHX1Zh+bBG5+pBShg/
xgOJhvry8+1ZkzDKCbwdGU2jHIY62++Sr+hVmtFhMiDnsSKJHmWRdfeU7YYbJKTb
Z2veN0H8R0V1MTun2wzODl4FTID4tEUKS7MV/Ys7uRhfrhx1yJeB3kwFEpPLaFyQ
idV/fOjZiWiHlZbxLHZKloCKLdDdYlhcfvcrSeLVx1e3TYg1aGCfINyDJuuvDdYM
OXJXkGKtp4D3x4DrSEqZvk41MWlu1ax6PG4OfEA/ao1lDiPDTA/x1VBG5bVUcvUF
kW8FpZv12Fb5vqHYzwCY2WJo7aBLKsqfsMDCB/W6CHE=
`protect end_protected