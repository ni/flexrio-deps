`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Jm2uGAVYfY7w9Y5qKstopObZuZAEY3b/Io3MSEcWLhjjnKulVhCBBYAEQrAzzGsT
vMbffkdZgjdXQUg8jOLJXSHZ0Dgbnob2vlppjZs3bgyHCF7MoJ35E+LOsaLimUA7
hlqStcK49hR1hdeBPr/OwfT3UeVrRtQyq0eJXQ1UksinX1G9Pz3/CmcGfTZ/C72x
p9icpt0bkY4/1I4GBvNCsA6FFKH947JqH27OPACiQQRW/K7JToQn+1uhWr3LA1od
lbVrWu8PdZi7zW9gK3jiW5GaPjwbYQGqeGFs3bTKBILjb7sYHxfxw7eDLVMAIu5D
W+OTIN4JiHiE1gCnNEvkSQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="pm+c2fYA/4JT1uhlJGVUubML8hZi8lME4xPobg/m8uM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
nBaXksR//iZ9fraC7WMJWWSrjqRXHxmM1Y0+KKN3b10NElDzVNMlR76DLrcnamFd
2n7uzsxWqhhJR5LBl98SXO3Y90J6BMbw+OBG/MFM/zUulxh2Si5YK5G9GCrG9gvZ
5JomxuZFDu9CzlWGTuRUt6FsE4Lr6sOL1P+hraQDpMk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="M8TXDiNa0BVMX1P60yIvW2WA9jKGGy8GtbuPknDnC9I="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1744 )
`protect data_block
/5TNZvs8Nu0G+mfp7M8H+iVAGG3Mh5DYZ0Gn3rRNhV8b5CcJKgjQajrRoGl/gSxp
rBAhtT8Vd5eelHgtvBjpvFBA/EBUrRH6CG6pqRt9r2qUDt4UernbZbxC3BC14KYF
4VK7XUges/yZxT12vZRIRffunpaVADwTqA0/Jq9Z360q6KIWgWHUqUMCpXUjGrFA
ZWmGMscoxrQ1wFlLHfi2u6bbRgZft7LckuYlhAlK9cGF7UEOwQ78Ai+hqk4C4gcc
DQ1d/Y+65bAvOSxAq6zFp5lBI+arDqKdfxOkx9nBtqzmKhrfAoBONTDYcT9480OD
LoxTZWsz6+8h5O9W6zW6I6nQG3dO1okb3iA1rjCEntV4O6zZGsllmZKXLmRiHeP0
0iTVbZpwmlW0qDPPQ3/2XFCuJZOk0uaMW2TNe1NNPvdgEsWT31Amp6Z3bfgmjPkh
tWsXTe8SV8etSdyDnFCkLBa+ojZooYl+6W8vtV6vkFDxOm9utoG0ttsG6lPoPJlY
LZn77HivFUsycZnmkLIQfF/P2COJ1LuiKWOMTj7UXkbfJxBfzvE1Kh31ucFpV/Jz
dgxiJ/4lOAp9zvAIz2u6FDYr4O+Un+R/PjDeM7TRKvuzyYPf4ut9heI5FUacqi8M
lWG3Ct9ynIwUUfrAG9xueg7/ZtGtOGByg4qvmglbeYqt3oxnAYT65zRwsdySqc4f
T0RGKu1io3PwufJUb8B1t4EOPnMgoOKzNg1iSQgTeQXJOrwdXUHdLYfcoti/nilg
dd76v3+6Lts5xZgxYnMN2NsXcy4DlxdeqZt3t+Yntyg4J29/g6GrH4LYsv1Ngzfa
n6jy3HZVGFXP844BnvVfurKITnsis/i+TuYlNeoaCZQXDUhHZvToTPnJFTR7Wuu0
CEe/7O29O8TFmngdfSJ4FEpzwWJ+gVSQvxR7VKbH6qNADM1dTE9UQB0eCRCOs/71
aubjs8eZ68tJVtDMA7OCOyLNuUGS6yXm5wHUIKjSigxX8T96nDkOyxkWw94GnYV5
Z6o+2+jZnUoqDJEMbcZoDxU7/I4FKAfhbkgJlYwGgH5hhsmLuGA9t/mZwOcavGD3
rd77PKSWjt6geSDPVgd4DuSFHyoo8dBqFqjvPfcST3KWJDfioaAzm4MFyhD2xTFq
ba1ng8ZXzjGdlW6Y2YGOGMIk9iSeZ2MptSWRgUV3dwT0YMihj3B4nYzunbXlE8H5
RO6yj9T1c1Rcga3oRssFTErPXt+i7gak0TfHWIApti4QXJO9L9NFXfpKKVi4MR53
o/pWffE1yIl4YMCz+gYp1QosKEmxxdzOgV0ngheW74nwfnu7kB21IrIZ8clyopWW
Y/YjEZypIbe8qxWw6oqfhYolANLEqd9s6s/xZSYDcgxlomhnnzVsK5bkukmtA4hP
vplcdgs5t+FNd5Tq9we3b18qDMAEftBdTzctUtG3fUz2h4e1pYM7EHFpDN5UJM10
2X+ntoKKCWxKuXhkqVTCRsrd8qprrBWyRCf4YtDcMtqH0b0Eb9TsUcpTw0z+8SsF
8lc7ZQ08eo3yL/puPCgzdS8xomavy8zx3s136Oh/pXfUMWg4lH8rJ2m/wDoj7KjZ
93RlRVxxbO31bj/TORuzOOXQhQFdn3hvPipm3+90aZsbdwzIjgfoE+zWV55EKbel
cWhjH+HM+cGWYKt4cvxpQXDdzhizt2nGnyivU6AZevpee+RcauuqRh02SQkHYbTr
pA07RbwNoBKd5estic6RovISbtNkzr/Tj+Dx7plPzrb2xFE2bG9AcLAVOKMMJ66M
JPz59/RE2E+XYUop+9kg1GV1TithURF3WlvgUX3uMDER7AxdxRdadUT7N+mI9MHj
Qfwd/LqVmMUWvmM1e5lIBWayzh/rz0iySEzKasbF2Nn8bvAP3ouRydQvRKKQcWUn
TAIHlkrxhs10FCAvWKm8ZFMJiqPhkvIpGX+KsxYJ/1B5f8+usR+kceIyCN02kexn
+dPiOqaITMLEgcyWQdOLtQtmDh77ZNH6StY/hrC9xGMuRlg0ti/FYNbZr9pPPLET
9lYyCuvh5rwHvAx9SOn5ivXzcJy88W7SaR9UHB68xOwNu9lBEq596z6zzNzHHeOr
+LzXQ23UfDthE2c5mlDtJcOmvk2KQTiLrWmaM/bnxUPaS0/22glRvxxn28rxHOLq
9jFWEWamhNmUPe+fp76nniSb50VASovrCIPivHKrmE0x9lHJJhnaz/uDJVgLUdmT
Lf0Vk0AtwMxelwQsRkl3v9tRQWYMhdZnouk+O9QGZnMHhSlTHi6DlpGWsqmOutSr
ZVUzo41vv6+f/3P5cZYh/Q==
`protect end_protected