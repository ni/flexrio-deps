`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1456 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
xI6xg28eTBkT3MzzlHKeZGN53LkMo2cyRplnpiv8mqbTMAAilL+ISXKOSUY3w24y
snDl3Mug5wPZQ5XQCmpi07hwGN7xGuO6izIAWFPPJRspkZbvbKmHr9AUR7BCvrjd
DZ93ZrgDnsgZ65HoUfyvMRzjdKapY015UoGdHHy+FqvQnCrFSCPwnU0wrhDpwJZv
Ua9nNeag7YxftPTaDhLWRovT1oAuRqrlJpIsTXumYf8ovKHcq1nDPvzd+oPxeb1v
gnrYH1qHw5EkCg2830yOFxbJ6FHP/MPPhnJcV9K/pSa6AeHWmC4aor8C5SetrV77
xYMzSw/xGDEZcVsM74/MAznlIiafuoXbF297vCJCOKCUmz6Yxi3d7VZbCEnFqs51
fh1GSHpim9HrG2/rur3MREKLS4MR+tkjZ13hMJ4g75Ly6o42ilcofaMHABtK6u9p
0EW/HE6z9livnXvvPMc4DwFVlYNCgQkR7caWM/yRIyDLy0pX63dbiLn0VoZ9ZAy2
z3fEIeTAm+D0VcLQBuNonqqeSp7S8IKwMX5iBnaGqBI/Dyz++daeLSYCg4v9KIGX
GfJ9n4s1lnykLwRLHo4tP/aL2SCxk4+zYGGZjIoOIJTy4u1nCLmdYfm64tuxeW4J
ESid2n2WDGhq3k1/YxIkQtjqLhjL32LXpYacx2i8Zz9iQKRW1SVur9hAhviX04+l
oVgsF7EbdV1I1dvNqNNdXFGgvs8OcIIwN1wqqaec93cmGxN1XL79JYDI1sSERC8e
YpB+ZJI4RqhBh9ZvCeIJenk03YSFmRrm2E+HVjTNd1eHt4uwHDPLR3fb17/OMj+W
45L9yH9AvJRu97aTYLjb+7by92Zr4OXfSdWeQmBe8xX9SehYUOKyobTtzbcok1fZ
/ZeZrGKUmvNQZKzYgOh7kuM+KE4TmiRDczJlGlGTdvHER6xlln1sGjiXICvcIqAk
WX3iCnNM7a1h7xb/LP3tQ6VCQAqDAN9CzwTSGuw1LloAbrpaAHsibcbq7Y7FWdqb
7UWvsxn2vUp/ftEvaaE6oVmeSw2J2pLn4DTYq5SLKEE/n9zNNUtaaCR0qWHPL1yE
b1vFaE+8ybICcYaAe16h6M1Yrku6vhN59L/fHhnSxb/ovgkjqC0ToquONRi8ySKP
oaLbOl7lWb7em5R1fDSP2TKrohsY/o927znelbLIABS0KgsLtpHTt+kAxeHs9bP0
OQEnjKIX+inmWFTI4R2QE2JfnzIZD3CFbReSlntPtAuFfrigVeF9ykK7naN+os3G
VJ8m42RhczPOVq9t+VFETN1D/iuIcEhZMgPJMM4AEc9gzxTOMa45HTe8k1T2HJ0J
c3Cl7Tr33X20osRY1D9LKXTSLNW2Sot8QXsZpoqEt8+ejxxDknXF1uU0JLa9W8ux
tvOxSq5sI2tOM1bhomXi7lwXH9jly2KT9wfsX6qOqJCXkrI5CIpIgcBbo61/eLRI
JVKfpBlGwY2OxXwX1gww9qyDYwnAj/uV49SyBiJpMQxpPoS42NHBGv2XqLZz9mfJ
XjNIkoeYZpMQyM7yIXAgFeZ45Wsz9+PIc6EUC5OgvUKRFA/L8vxdVjSt8rArdmlA
4I4mveaku18DmRGm4i+MH5RuTa/y86xu3880ESgB9a12y/GHBPruE5KsmBKHCUOb
AH1fxfYS6KzRbcfVzjCv1B7XurlRnh0EAHBBp6T8KxOD7+MThDAgJE18SjTa58xw
BMmhcEspUDFBrkz+SEVXVlAz+29y3IxGzf0zqlEtBhbpcgHq8tU1Fsnjxi1EwjvT
03HF0VD4tu2p4VI9wF5zjg==
`protect end_protected