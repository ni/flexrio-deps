`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6496 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
Ju3IpcJpVj/VshHyynUPTF5eD4vnEDgRfA8fED2ppvPpWrRC7EzAw5tmm03bCsJk
pTsfJgVTJbGLnaoD3Bjb4hMJ/prSwpAyenEFsJ7hcB7vkE1jMkaE7A0fFgauCane
au8hUHiNZ3lV3s8Ia4ihxN16RjHR8H15/jtTugXorVYMWSJrfNkZQhDmp/ttMd3J
yKT0sWDbPok1ehAMzV6XvgalYpdI2XwCmT8tHlXZITaqqP/X0KfjCCVZa1Pit61O
cKkTYDFab+xySrmbEStamj+Jl6AVZPP4MpqZxPEFTTTDAtbxhxPRAolRjnbZZvHS
WGodJ7+gU87H0DUUf+HT6MwpREMunapJ4WslmkKjEuqGUhfL0YCPE8BvZgL6LBYl
kfBTsOgavauZBMPxL5oPMCD3KOeLn+83QaHd4ZdplaUY06lRUpo+QPJAMBT7t5Pb
BgYDfnTxSQ6K9vQYYRxCh9WRrjfc3eKGK4KZwIqkGGSgNLdMt30D8sEYdYudbngc
N/WNV9YTpj5ldPHbodh7zrBcCwxd0O+XtvUYDWrfGdLgtPddovGwHKr1cgzad9a6
GmJ7NHKPSW/7IE5SEmDDdVY43c9TAQNpao9DtEiQ/pZKnWnvQSMVr/7L15b0La5y
/sgzmcPMvR7GZsk8MTzUHk75uZijw4S6l7Wc8ps/TxcKpaNCctd97N9fLzqk6DmC
pUG/UPh2chZvugn3FeyLf9OO64QAFcRMAJDeFK1G3QmN9Lcax4a0n4i9WZwBaZUp
x+6ehUBGt0WDOCmWFkTLUTVJQlIYTIyA6/n72KtCMJzE7rQVdE78wktip5FdsxtE
G0B62ob5vJUmfx9RKr+Zd/y7tnw3S8mJCOO3IOl2dwCFN09fVG80TIGErUtj0R9R
Bb8jzZFXcNv4ceu4P2D7aLGeBdDOsMG12WU7jB6TiI0qMzR33ayxVS6UdUq8kHIx
FKcDZrJGBP2YJ4GV2Xw24j+XwpCPFcQgxFRDpfQ9Qbfn75EKvdjEb//Ydde5AIw1
uIKkBWOM/f2548Wr3ZOOw/C+YQyz7FJY75X9o4lsRwDJDTNDxv/SlxJE1YSX8fic
LXFK4yAiqar+WGLNRQpu7UmZd8MeBwzu9OH7iZciA8mhbQvEo+dmSQsmRCzfr8n/
h/u7YU0JiZZWMNU8WdOFq1H634yf1c+IB/ndqDpEOuemMAlXxCmr0S0ubOO+5Vt0
/B1sFdq94MrbMF7jwVSYuJh/I5Ep9G+SIiKyJ5hXN43ltEk3+VoHlhh+meZRut/Z
UkM5X9aw6nbhmjIV0GWvcZ5REspfm4e2+H2cEeuSXvb2E6qw/e2bu9N1bIO5ITt+
xo4M4GOpwCr4e2gUki4z+yWG6JTt3oizGUHFPJ6KBiyMTaHD0Ag0Ngx1Hpkbq3HQ
DBFAJuR7MZ15px1Ktf3G/vjMNfw0Y95en4/9VfCUpEnJcBi/8TrKR+Galun+NTNf
5V2LN+cZ8yOoNCOfwLzsqS6bau2lMTUha5mcFsaCmNQQu6Na4LIOVepG/iHlMfGn
jpfZPmxJGyn2/AK3CIQhnHgQU8m5vg5Moas9nIPWtO/ttBP086HetOPq75xDFUg8
FoXVJXsQM8Yvr9epa4MKIcwCsxH8txOxJ1cKdkVr1EH7vOjVEzlrzIpZMNx7v+oZ
hgXmWZatOoHyLGecIOPIti3KLT2sMpjxzfoTDCdJ0pYgAxdMZylKsxxrU0203TYt
OxcWK7REfB9rkv9YxWQlpHR26g+U93mNbfJ6ffyHtwPy7irs7JbFjPEFhJ21bxJb
Q6XOi7RQFKpL2HsN67VKGk2IP4vy2E579Fc06EFU38/noyecMrLegPsN9fE74IXm
HYFKjYi5erMUkxSyhigBXwnlWXjVEYI4nCPywk1Ul/hc2b9LrticVbY1Y4DyUo3u
YZzt7P1jJ6HRe+3o2DMONGHpDwWHto5jwoy601izGUEt0+8xryMMg8pAPFpgCIBf
G2wk9+8ERIh9qAD0NEoJbgCTq0Bhctqwk1bHjfsT2HbFg2+SDM313kwaLAP3VDFc
xq15nPXuOGE5WSmTWhGHHoKFhlZq+sgm85jmp0n/b7Jgtn2FStkXO3yw/QrssvY8
TdP6HYyd0bRAZZ7Kc3TuYsCxl+VBYRNGljmXGvKjDgjPW+j/Gzjq1hsxlwAGt1C+
18HC+sNQ5QhfnmEBrQHsfzeFi0gcz2FS1EuDuSO2c9ILPiuZ1WHeRrAJHmeTrJkF
i4kcx1XD619sLG+akfP9RBPgjr+Wc9jHBO4l0RJ9valxrmbuvrusnxkd7ZB7ClrN
7JjhqYysrSvJW6VroWAO8yzEIuhLTC7M8xw2o9R7ff78dOrgsg1X35k7y1K/EEX3
KBTktxYwU6KVUBypVlcae+79D+PWoRPm3z8SHvaMnm9OzXvSvOr3+/Zs8Gb53H7L
f3+Cm3RbgUA3m+6Ldh2tTJk9nFn/TWKyHioKX3R2EGDewDznn3Lhg0UD1YoPveuC
JFu+J7Cbfc7AYUrjbllIXw0o5FtoYxiMF+xbw9mo/Sme0FuzrqsX5XYOTjNA5lyU
OfITu4CaP3gARI7lmM8sjuK6JLYXAd48hQqXwWmwGzky5RcMRFqmCNFcHWQ4r0kF
5waGmx2nvFM8c7hAmlWJwA675wcGb/JzZ9KeAYfbbBfV3mL6EjxK/lEGpIEpVGp+
ZOksMKELvO9VQS635HexQdhiD+Uq9v4LMiVqzgL+qhZItaGyD2fIIgwMOSDBEOc5
fK2an7c8uwhTiwzxc4w+KLlewZaZrrVqP+oIH7tOh6SvhXwMGBhcpLDNfwk9/9yL
Eubps0/xcGQq06uHkS1v7L7o77NT1dOilx8NmAxTSpJNq0Ai2897Hcs8FV2VZeS6
8IDNbvbxGQrH9Nlv+1OQeTBBQonYi/s9l/TEsNU6kdYx45bt3jKDh9clDk2E3P+K
hd5zEYaGVtjR28BAjdmWasyH1egJZLEDx+zP1R9piMooxgCmAqLi0DMcYeTalmr+
g5VIvm64Q4+bFbIFEDioiVLz4YWHxK3txloPV+KAq1PyZwzxwknMsNlJQz2KffSb
89XGj6kRZDhSI3DPl6X5y7Cly5HHc2cHu1XlCzH+QeZcHOILdkocqxhZFbVuz973
dyU+T032SdNnSjEaCuZzGM8GuMhqlJ4RFflrxGvZ4P+Fuwgni8fHRKHrNrA6lh/+
cNTMBISCuQZLPgfiQWso3w04V9dVstLXszm1y/6dVjm2SlyhqRz/mPNwJGz6S8rX
Y2er9w3xqc/uKoQ2tbqChoStThFN1wyUpRr/xe7a++ve3pN/1X52K1q+zJ50oUZf
/VqrBSI6w4ypVi8+OTFSlN5mCGTzRTQw9+AkFGxaiKnUVYjA5JhI7f8z2e57NKFX
WfK+gBVeFy+j1ay6z+o0ihqg9DFFXVKs0gjrkkB1OqRe7TLFyuPA244XdJXJecsI
nBhnjKG3tvZcON/hPmvzR7CVir0QoWg53QvLPuYVFhSjBFu0C7g7G257/NF+ilTQ
YHzZyBzLRMlEO4yip4cTXF5di9HE7k2HJLF210vsfVaSYdNzNbdWXpcoRzWMR5Yb
ZiGeBsIfaPXAO66oIr00KLnvZVJ5mF5+WeQYZh5hFZSpbzviEc+UQEtn5FU8zhdy
p3U1ioeI9pJzQLuZ5+CCnSn+qtJcH8bVGeBaDiA5q5VLKyyYbdrP88a4lIwAT57A
Q8P0JmRm9ZM7XD7WJgt3QcozjAJqxWikfcYoZJG3ikjkGA7QyN3i5aDgh8Hw9uGg
9ukrcsbv4Bfw2qtMOFDxlFlo6WJhq8B8qMSTHxL8Z36wkzLhEIxBut6JpOvA735g
hAr013QvdxgXQmR4bjmE2ug6LvVnSwKrGATEvkm5bo3MuLNGSvg2NDHungm95TNA
VIyMrPCOEcGABks/2OZzyRzJL4cdhlEJ8SAaHtXEdEiZmvi6i3olno+Yct2wpP94
ioQS/ITi67yD4QCTs6COIxJXO8Ojzj0qtkzL7ru0qx/GSZxxOOlieyXHzhNwGZ/q
/ruEBbGd9Qe9sH80TqZciicMLrpwGAn34gPowvnjeWpu4I08qAKve3/usGw/c1EN
tP0vdUEh/sv18Jp3ALpvZ5glx0gCW78gx3ayGeQBuCw1GwEkjEADUzdyB6OTuxv8
2Enx27slzbJWRiPvLBozdQRm25MkO5zbqXssgVfZQW38+SG2N964hu6ncST3rgn0
wMtezPc7gANIkgYiS/7aFTfrrLDIYXcBes6c5+7fzXkZISGF3291Zo/2jlMcrtqg
u3Idh0v6SiY6wjUlawFErkFx4TeeRGKpWZ/vMSVuESrX8WPq1CvULeMwnJzzV3BE
i9vsHBpGHWTWac8X1WvyiKxdkut7IMVDbG34Qu2p1dnM7lcgbq4tsFipu6EW0jLJ
c7UE5luF2MjIunhO8iddoycgKkkvDOn+wzCEaDCiqLmPGGnXW68Ez03bpedjW8rE
pjO5aO1bck4LRiEJItI7Jzuk7OVInv5upueeRFL04ul+81p4e6DAAsBdQbQuwCNY
6uasEEv8Ir9u0v38sXojGRP5LzJ3n7rygjpfjt+j2Z7s+A5ouaANXBwD2I/OiMFY
v1zjfQUdKm7GpN54ds3h0C/lLZ91pTanRgXXQT3/s0iY3nv4HCabqWiTfewjpUjn
TjJ9M2GbOxdeD9bLA/f9bpSIoHSUKC26odBMhVZY2jha6bZkQijjuVyMXUNLSONe
MiR3ksdJ2eHPKz8zP+Hvu3NKs5Ci0xt5leIcH34HLxQW9djDEARKl6tuXbtBS0kJ
178kFPv57a/7ogJGk+SPVQ216FY/6CFTML6TroPY3ibSKsExFXBFh3U9EAHOp7Fi
nlnLajHKpVEQ/nOq/q0q5Y9FxCJ2cMeLpUJwMxViQjJIl3olXWjaLvUfnUjd8EUK
/6yKcjyqiCjxccHGkDCHXDsOVj+LvwoFTLai31j+eoVqSJ9Cj4m04XV4Y8Z4mt5d
4aDRFuXtvjLj5OfUs0aDFhsZJ3jSiRFifKaNbdKHBD8pf1KxLkhyBuxraIgKy02O
/LqaSrTEikT7sM4FkpKpjVqjKiDqHnjI9OwSCuASApIQpFoxJOcx0lccCaVAO99j
/kiicY7D3YHaUwnrfYEIKa5y8W8ZhxYMgKEiAXV2QJ6C8K07nGWj0POG51sckDsA
tAYJWK/tLdf8nPDoi0PCkPMZRnaZG1V5/Amzu5pP5u6uEK3mBK6BUqNhuBNEABjx
VHcibsH6J/LMMCOOJvcs3S8NgCv935N5+DtkM2Iwg6fiIwubpXIjgRSPWVabyh8s
6uevT2jqiEEpdqfXpmPb4cdIPiqo3IBZIpxQi/Sp6xFxnGOZkRqpSLBExMp7skBL
SGeFHrn51iJiZS9Cmu+ELJi1dPqrzKYfu3dfs2jl/r+bkhUjS0trEvuKunoX9E+K
Wxv8Z7kYSr14UkAnf9DVrpmZ6/XC1rlz9sqtyuhCcdwxUvn8vZgG35nCXESnuFox
OMIG4ffNS5U0NlunWmbxX8idAy35RQ4cXrsFCxemfYpLoYJV6isRFRsYBdi8VthY
+/TuP1UFh6ZLIt6pXl1HoQyfatCJteMuk456NsMSg4GoBSXRAH7EM02s88513Sh0
Jro0v2nUOAG8H2/g0xU9pJZlrjO81RBcSiRwh9nPCv5mlqDgdlv5e85MAhXkfggL
e4uV6qxQ04HAX00CMHuOUubjupQEhuQJKbDmxyRinftkYtu7Q3bdJDY7OgZNfOb7
qp1BEAs7NV/mtTzpFCSpFhdgBPEInK08kooqWssycMi2/9LGHPjgG7tbUE3MM8cN
7Dhmr0YB66W2btPsE/8uz2aZfHBAit9CGTa341yAmXnO1OevbGq6e/gvO+K643Kr
IaeoQ5VaaL09nzgHmH1H/D9L8onK0z6omDBAaq8MWm/03a5BbQhxcOFIUz7JdvWq
LubdrFSg6Gf7pFom0VyFvHZp33wkSvdbmemfwu/yrBC8OgmzacT4hKMAUfnsw2O0
cNP+a3+pQzzGS+ZDUf53+YezAdBFsA+AZ81U7XqKUSI0E0R8daOZ4Ucynilswrdp
m0Tco8mlt/1S3Adh1hnVnBejCL7/quTqzkE5H2WGsryOIOuaG2/bW98Ga9YoABLx
6Ttl0gwaUwPBz6O41l3rzXFdeITs+/rh395lD7q5rzan2clCNZrFlp8JOpWZhZ1T
+rTdGHE+jctxGo8EGJ8ZaXsxj62bXrFh9QJ8PcN0GklN8WX0usVzbByT8qTpInS8
TwlxSxzv/DYNRuCuHWVJiOswHdaYULhWAe2pNNrwoxo2rAZS/QxVE5SS6PPz1Xm4
u9YFOPvoVVhLjtvWL230YRjusLJr0vopkMPKGmvoPIrbIZZOPyzkoxwucQFgquhl
8n8ArTDIFbfjw/ozkJ9v8+EPWfeVlXDoziaeFV95xJXaeVLD4jMcF4p3BEHY+5wA
6Onc6WzGuk74eGB0cJha8hc3C+JCwoX5NNGcpRD0T+vo/6NI0uIcDzHk/nMUkXaU
iikUNvQYwJHrUnt+I5ni+GKTV4pOY9wskZRziMIqKTPGy4oyHeyrZts8vzBqs8lV
NrX3oUFNbVTecNg1AOri0svdwGVShOlOPx8IRyE+eiWod/neC3C60QZiO0zmOG9H
qg5AzyltvRaiLVFigCr/86MbJyBulxYh9+lOXiGftbPYiQxcrkjLfzVwP8eyD0vK
IuRz9OjfASyZpmUoXWYx9DzwKx6YH8bzeaUlJ8GFmfMbkAgEDXnDfPolAP5qkcm/
yLM8EDf+OxZ6p+nySVeT0VTrLyFgfGNAjSDaLLFyKzLTRhEs4T7A44Z8HbGoQl2O
/ES50aRCag0rnflMv/JXSAj06IDw7AKNYZnIhDNlNdbbL36gWeAEj2NM1beYnRFr
4tIAXzcg1wDUryFkuDq+gPqpY5aourqQIiy+SVYt/umE0NWghJOaMee9QQuqJWPO
PkuOoTVpb7Xs41IR0LiCmOgYm8pkUt7gHKsf9G+bZTOVjbKo4fZNpXUdi1EFfOtF
7GJvNFRQJGv7F0oBnCKNxHSFPAKRk6qdbpYF1kINgK4pWHmliXbvuYZFg92RmwuU
YLyqB6Z6n/75mkmst54OtjGCOXXd0QK4QEJYOE8vyiuCTtZsA+E4DMPqG4tYhzaQ
p/XVo4/EqAzI6qo5D2T5tERSa8mekXjCf+g/JOUioEleRLLyvnbnDsJdRTxaSpMq
Sq7ccyxNzvE4YzoWOTzvuoo+m1XRXxf7fAQZYAtgBXfE3xKL0xEbMS8g1OSGfkMh
5b49EtU5qQY8XBJUJvQ6+LmipvUN7vc/iFb6lqoet4ImNDlJ/MJ+1w8T391cH49r
xDC0GlGBTO8X6jegD/TNIKtD8cy1935PRBfldtz2959D2h+OT6+73R2ltvzfzlYd
b5sn1MrB+hTTBziRSNMbpbLbKGlAwz8j41IEyh5v5XsoXZ2TcHmvL66YU6reBvaY
FDBQFm4tDzgv6Njmtbg51mzr1m5origmqseuaNRVMXbJGqnXAYtcUn8/p7o7xB/2
SSpc2urGih1X85BE5UeqWy5ENH62llPQ9RaUc5GXUMvClfQG9IYrvlWvWlL0VMHO
VclgzmKq+Tt9zvouaCdf1lDz2NctuWclMCWLYe5TnaMIDQFE1ml/OqbrNEGCdSfm
zlU5f3fuRxjP4WeRYilPnG7/1cwIDFpbqveOFsfxjoPb4vcRbozmY+p/EZ1G+WYt
4R7Jnd9aYJVr09d9uv/oaaqZVi1B+mhal+ZcPRMU+XMTeG3WowQSkhMNw7Ynl1Jf
V7fQw9FBD12l/D6EpzYdNfXw0yveLqfRyeox7kyIXlN0tBr/JpqpSwrqB4OM848j
ZNpG0YQyHGKhBOxg/QDTxS0KW/gl6uXNQYy1qSFWzCLSiPMBGV230TEWcgkUt2E3
J7PPpj8QpfMvEBAON+WHk0kfIrnR1oRYG5zuH0GIX2V6vVJT1/4+uNOD3O5FqlIq
06hFNbO1a+3Todh0urVR4yfFujOCcBBCnF3NcWmbwMPnVstVfY+T2FNEk1U3/7qk
UzBm6y6nTpfPy5yYq8WGV3h+GjiSjBbb50ULjLUcE/zUBn0BrTfkeSuJvQT3N7/m
P6zrcxybaXAvaXoqfDxQQ5C/i6WyhrLu8RVS/hjpNnP0Z5ZSwnWNkx64z0jF1ICD
B150CWbbg63N+zqSZc10WRLCOMruUlidUivRIFj63hO6OGbUHGJWKVsNY8EBGq6I
4mmKkBD0mf98QoyZgF1LiigYpC6afqf269Nz2jQJEzA3aFXJAlmOrn2Tl/hj2Ajo
TszwWgEn+sWvuAm73uVKyGPHGIlAMg5OuV9PdaevmzSwDIP4aaWUsVDQ3ooMNNzS
nW6t31m2Jma0JxeGH6IHgrI1uROFKmRNGiJ36g3CaK+frzKRmUr5+Q4tF95Og89a
PYAdz3x40TSg16zwsqsTEG85PnmgakX1+5ToqVvJkgGNBiktxs06XFSfZEivu/Bp
HU+nbEXK6lCBwNeWyt8gKQ==
`protect end_protected