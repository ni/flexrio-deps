`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11232 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
r0poS0ytQydMvF+aKdd0eDCyttyHf6aa7nPSYXkbayDhg2eRzPaX1BYwNFpL+lTV
l+1d9atFqraXWnOP55/h5dmYi86IEXzDXGbIM/8WLy9IjNlKDhZaxDLHgW7FTmFs
nadqC/j1+hkpKs/DRiUThZ0dV0LsS61HwZM2Gk3Qgwb6QPb7vgARe1YlRbtSmOHj
16kWTvjFMJx4Y189Ybhrpa1iNKPUqSNTxwg4bJW0WlIUMn0L/oHb6LyX31euVpR1
eYraioP1pSIGrVkhAA0TGGYPBoMyksjYEgkUc74qQr2paQGcOmIhURV/x4HisSVD
bDbhDHfO0m34532i8lRv1WjkGUU/8uzTy79LYaWLt+mGEN4p55bgG6DSQ1/2oyUQ
fHpPjHWniNG+mUPcDKe4zGnuSS3j9+07P1pxcWbYgiACpRyKrHtl3+v5yXl/hpnP
inI5KvOd6NrVKJ41e9pjgiYqgCjRvdyf5tVonOloRhlciY5bSHLkIqrUu0hoYWN9
gy2oB1HcdmMWvH1uEDFXtx4YW1w0gibpS3NrxX2R4E/udFdbPsLbB3p3JIl8p6CK
HEt6JOXNs+sos0zmeJwF3ZYcs0BZf/SBUKqO95FwacsGbtnJ9AlKGPZhoskT/OMm
WiKsYiKbWZLcpjPPJNIpG+XXmnhGtWfGk/PDufz50v8BuSpupP3rz/XusXNQ6O7U
gEcsVO6yx4ZN1aW73blhEwlY5fQliOwkvGsXUG62gT1a9RR8kP3hxd2IcjKVtN4U
A17Ncl+x3jK5gI4suro5i/33IoZVi2lvFj2SNbpli/bhZ+cRfsv9dhQ7dP0Hz9SQ
WwrmGbEQeXKKYyWzjWv/IubS5roy/+EOdn3AKtyUUAG+ShuCUy36Wp5eI+iOqzZ6
vR+/T1njN4vHOqnfEGdNBSSjSrrwPub1iCwhF3gmZS2zngiGEF1SoxLnUvU9XD+6
3gnfVnq55TDrs8J5+8lh9OR6bsuZ1e3gaYJ9o7MmeXX3kIiv6fxOo563arN+oX9W
dQM+DPG9tUtmiSIgLZx6Aq09n/e6GlV3Ms+zrlm6HspG6ktk+18dpuhPy3QlsTp7
dhJ3nL4/ikRTCRS3mJCYVDIhcPbeWyN/rXf1r4jDO0moIKTr1Eb+9CEqQBpPC6iJ
ukn1TrtOxAGgmlyHCMEk8cFcm2Ez4ghFApTWB+iVKhq+jO00QMZKmrm9l54mmRX4
UnXobHJkTgC49A7Is+qNcJkrUAUYCRC+4qTVjWa0skix4khRaLduaOEbNZXzUO6V
fbh4mDDhM4wqFCIy7eYHcIq2HfVh+mByfBOIllv3R6PJodQvyBklfKMzmx7YN/im
7kpfVYiSw245J7aPYlPM49EXTQpRrj8XOD8FWnc5AuKmiqWeh1uOYDOPsjw9a9nP
77iF5P8uZV2zY0NQyXxDyqFKZpwgDl7XDy71ApHqshzHhXapLqdAVO7Qz0Rz0Rc8
We2UN0kgYT2mWYOU/AENEAQcFvsgi2QPq9A4uO0OauOWe3wUtbTXQZ1D22Bq6lMi
/4S1XozHh7Ghax4P7io0b48WaTWLm6BD3axljmYaQ5lu7F9/xidkfCNYIJOwZ5uA
6DvbPlcjESlNUbJ69V90vDGZhAcMTnfZl0n0/KIX3cCYVyCDmVwHo5ekEHWsYwKb
HZxY7b/kJ9tT2zLtLUslX74N5efFxQqIRAfy227tQ53VbtggkHaT9RIhE9D1ec+5
RWRsqimh/O8Sh825oUozAfBTaZIeftjjvAMLRkO2zr/ODmhVD56OX6dvuRtN8fuX
ez5TA28mM73F+du/BTloJS9I9mktvSkO0edw1zt7OWC2avESdTE+F8deDPoQRqpP
Zw9/kajEkTYOeCGzYNGNiRfMqtk+bR5jmBFsWKviGNgh01R2ukJDVUnfcsS7BdT8
AnNuTQfFt/2brkQJI6m/iV2M2pPodOCpd1YP//ZTXX+UX7+ttAdo4PaQaKmiYxnm
Y0QDT49wPX58ctQhgBh2b4H+In4x/dUfjrNvA3PImsXmcha1YIH5ZNfIBEQfwZhJ
D6kS1Vso8KflHt+c1M4PVU3EeGal2Xa7f4YQe+ISrO7fjTNVKyAtCQmSW0iW8zF6
wGQyUl24Vt/qOklq9fJvOmncpzkvLvh/bHrE/eR1aZ5KlYPNyrM3e41zyH66Zkng
KIsnfemhfyGHkOolKmMzlunyprrB7CZ/I2q4WHQ3FEvi0uVWvzhUy2XFZlCwRfuG
gPGp1W9GfM0QUjpRgCqZx0dpdcLsinPlqCG7gleFJ17NEkSnhG87Yc6RgrKVe330
F0f8buiF9xZT3j6Kymld+JfWs5X4eYrZzJipUQEFp2v7wyBFfUh9DT+p4URLzodB
eklA8MYaqLz0nZDcNM94Rrb0EV35w33ltzykvlvfZm34cVlTE9ENwvZs4VOHSzBB
rWbGHidQoRyJomUBHvh6dfU6o+whn/lQhNEqGqTgualmXLx7ThY8Nwtwgt8PdhVt
Yr3DKDFrE5ZCmsvx8z0dfOLASyG/mfurh4BcH68VVjtrJuu4fkuc02A4S6Lb0nFt
fKqq8/eYhcJiBVf1XjRL9x8q1vSJ82br6dFXxIa78oIY3yOoKau9OYOH/bKXY85O
800vfTUuwRxOMDXu8/KHPCE+eMwz4L5VHZf1o3r2HPzGg3OOWByE/zKL3tdNquRD
X0V7SFhHso2JHKGIfapTg1KVT9y9gcOuNFTMb33eNkoIPM6SYWibreNflepV8zkR
iypDh3Q7nD+6U77Qk2gC0+nuU2h2kb44dwNE8y7lBn4w+XpT2FraKnuY4eyaOTbS
CWsrOA9ehQ055ZMY1zV6nEf/IVPKkU1xL+4RfSpZzt0wz+ej65XmVje+n1F52bQi
OiknMic2u219BQtGO8Fbxze9ux3KWjz+M/1d/u6i7m7AmGIflU53QFtqEyOeTZwo
+bfXpUSJmPPWb0RZiNjnLMj91piOhdepL2rqruMVJzZq7cmlm+5lImVe//n83bMg
SLS7jsZni8mYzNKMsGA31P2m45NJ+6KHJ+gy+yNr7e8ssOVgMNAv63DNTeyHsomx
LI4x/nB818CwCCHXml1BiGUZSJxfOGnsHOkwOroqv0W2/df0uQHVkHedI+J/XNKi
uNh0p7OhCEcWpzTbim/DUElAy+lW5qHEJ76gTuvtqrw1y3anL1OhKIY0QlpxvoJz
2I8ge6dngizk9wxLgQ80XMGRH5BJ/IsPAflu956IsYBWBMNbAHodFdIaQs6sYAKE
OtJudRlkvQ/vCxbrr9WDmYCvsZEGsGAn1Dk1s6GFRd5fBuwCkF3fQ9VFaf7q/noD
RV4TtWtENT6qFRoIHncgPTk82XJVNtpK0tznSTOVh0J1uGB0ZuI9GwVSwBf++U5d
nIHLBe8vn680SZyhbYVbvkE3YZQ57pgd6kifDGSIKAFKxUCBBFPVI1evczH/xv6W
ND0g3oCAgzHs1ZA3Jnbo3q2+11pS7c3R/pM40mMQTA8Szt2/BN+qD0RB0pJcvslY
309HzjqNL12lOw+FEX4FwjhnjFTLonxgedd2yySXqC/TifDW8Ll8Y03jTZRo5FPj
nxCdX/YnZ2Z3Vo3QF7GR1BNQurvfz1XCvASJBbNGjxtYWprWK4v4n4pJCq8XT7zE
3DJzC4ZwslpPQfyCT/6cIZAPOz5/o8zwzPgG/9DDA0P19q3sR7y0dUXdjLE7Vpsm
yq87Fx1OD/aqm+iT95dTqAXzOnwMv2S036MC2Fc+6zizn5QqsCkOw0fI0NRImPAR
OhWkDwjo5wWpSHjmNEkoUu3z3u9SZPvPUofVx6+4NMbl21feOGpbixxqASwmRyZ9
lR26M7wytw8FD0qU2ebFHyQYMY6QImnmOaFC3KOnWhAiOTSTWnWe4qDrt2Odm5ig
axTeKWJ9CY35+zqgY4OEvwLGCERGgW+HUC0JKU9vZ6iAa7CnEg14JGLWf0BgiRWG
dSJ52o8UWbql0gadzkvnYisbxXdsWo7xsSHRJ6oBX79rCBfETeY7gxVfpGGhu39h
N0Fn6QJxxK/NvenzbAZIXoEgUbTk7MOLeHxihaHJ6YP6UVBBlfMazXjmKzxAVOq8
ccgMAUfdL//Zb4ewUeToxKDylRQhfY5Ur1tqtOffGsV1XmVKJgrN5Kd+hgbiSqmo
8RGQ+5Dlh5b83Vl+0LY9czranrpnH+BmjsK88pjcaWCLvXKxQiLTpB/AEwXgW+fL
lD/8fT4ewdzGdoMKbshlHZEL8B55soXHTtFK4PEN3N8d64WS30H+EGVYqY8vsfh4
6wdV1+oxu/1Mmx6hscG2b6ujecnu1JpDeE/iJouhhF7ps2a8ZxMhtAQN+comQkWv
kKQgkgDFW7kgnX1Rz+7aRPa8sRiVXphe5okyRlkBCfKC9Xy0IveqBXnuK2Z/cZDp
QIVS0QJDekld3qRbwQ6k5aNb2nwKoZgGLTmPB2Elp+3UFsUeu7oBB+fPu+u9w/6T
LFQMqFX9VSEM0AAWBeN6GYiKS1/w9sbMf6Rh33m76UBp5J8UDXHcGmTfHp/gmAHO
aa9dG+dwNBgIDNPUAHelC/Bxe4kKrEpFtd4AQBsqXbivBoB0WC4L5O02F8zrhV6Z
uTyP8t02mBgOjImCE1ISa9LG0i9RZx3m5rg6kwuBwrTYS9+LS8mmdvsB0GhMlC8N
CZwoqj1ZbfyfsZg3jFPE4FbvlDJ5/QwdDjZ8VQvAHWpHznyOiMZdsL7ND73WZXek
wjCDuQmKU+YS1WsxXPF/zjT+AY15LffJxT1m2gPZUkFMxpSll2Q6LmdgXDCzoNeG
mQ6ia7gZjnisAsDUSp8oZk2UMM9YJcqm3q/DHyGod1IohiLtyfbt59yfShk1qxLA
BPLswdxglLUSRvjIFLoychcWO+8qoli5Wq0x34iHqwbQ0v8Ufzti9KhgnuiZbZzN
K37o9cd1DcJ0G638G4QKB11s/Wn5UA4n71yC6dzTVFGly6tARzeQR37+AKieYein
dBtpFnwx9IyEKhyek3Bdq6fYaXR8nrQ/jicEh5WFXP03zDjWuvKZRSHgdruDh9jx
iLiO0gGqSspxuKg/hQjXrk5fISH9qAjLpnxKqMI4wuyHk6d90nSdT+rWyx/tJRGE
qOEZLP2e0kIk/f4ySx7hQlPjel7yGjffri7CNjnKwCy6PXgvDdXh6Pfp/xJNvUxT
11cDRv0XNKemgpTd6txn9Qp8CKJBO81ue31fnD52gB3GHO2DfpZVmdiIBdRj9XXq
QtK4xgjxkgn9woZ6C+iSXp+isnfkGEKcRpDwCuNOemEB6HAVO/h8JLtBiGd6DpuL
zp00g9Vh0gpfu6spD+TKNs2PgrBAn0pAk4WNNw2BA01yHD+vYTdx8hyBV531eWK9
Q3RJV94BDph85423jTc7ijeogCrzEpHeM43cvzqBSikNSxejWY2jzf2aCj0kDld5
fRQ6yk1x1yWF3TJxt00Zov04Tv2BovtC0UaOgGdVJXguYNeFgvL9dzRwvesnZJY9
Ele0dRDbojETlllxoiuIE/a+2zjMdVobP4B+rCW9cUh9xH7NcWvN96SY3TstubN1
gYuDp0OwSFsRptRg1ZLI9F2HY9Q+OkIbwvBZq7K1BGiTr4UAQHrZcjpVQjSychOS
Fu12YOFAEATrtRVL1OxBE5NWCRBUR+0HpjbDjWYA5nmkpoDLegSPS9Gm6ojTR0h/
F6ZwrTU6bjQPlsJMXC4FMG40Mjo+fjC0zOfNuHoTf+i2zjPbiFetgVvKVxXSPXDW
Hb9HVbKzlYUK8eBXG5AHyVXU/NwWlAa2u3bpulupXezc4eUKqyBsI8cpjZLNFxes
Pe7Q6HXBBPDPgFBsuA5HH43SM4bt/rHcdE9aKBgm45MLtKE4A/IqJSfPf3TVZCus
wT1HOsaeKNRI08hag3Uxegb6vpIPkBftsIW125Bv1g56ZHORpzg8Fo37upzHjZbP
3tWgszzLMLbat3lodzDh/bmG0C24DLprLI9OS8S1p/RPz9D6hq3MhTZ4pToTL1np
Cw6n800xRoh+516nvNLGVqdZeVi178Ca5OtQMtDjHsgopTdC0o0FX7gU8T33hc8+
3PnFcdHoSSzql57g+5Zjb6bKlQzMZHeeWEr9LUbCol4ioyM3UOo8km6IzPVz1m+X
urCppdo0jzMap1qFT20T6ex6gb78AlvO5JjPRtNn/iujySIVclX/Kln9KJH2oQe/
HFSpbZv6lgfmA+OJE7KjgC4H8rOaWt+r2baHDD0tW8uNrnalyCzhgyNz6+wrTa0u
U+gofbD7FNlfWBk51qsTDSUGAigsVxk0R1DrdxgFphCN5NTDmkb8NS6ToSEprUto
BllNFltzP1TP52VHnP9lhq8nIFq5auXIeUO97xu6Ptq990Y15dBskrbNJObY5vkn
8iogebvPUtfAuXHKL+aroy8NuKdsuSrSg571N2jeq9eZReMs3gvIHuJ9r90UTJ/1
8zJMj0/R3gm7xp8isSo9qq7cpN4T0p21hZlbGNVEmibf8+C+rTopUbn1X4NSeRk1
nSWdThuTdZY7BalniDrA0kWxT2cVgQVJfPPeXXq3eX/4U0RMim3JD6L52W33w0Ie
07u5e7pgbt5ytWNzkJadd4nnzd0TmdY0tDPq8cQNkSgJeEEre95LK/Qhiw9GrrBw
TulXqakUHNuitDxKgrrsrHG7JK6ubQXmHBvtEPthFEj74MYkteLCpw1ijCzjQ/VC
Ju8P2RZk+N/kyzfAFIkh7ePBD/FOOH2V75gk6AUVbz2YHOzaxxm9uSJ64C/hp0JZ
QNqZgboes0NKEBsi/szoydFEmEq4KxXMFyiCxSFy6azkKytDMxDtJHTOwO7Qb5dJ
nEMtBjJUEhJELWaDQDBiBPw/ys3sOc3/KzHVNCwS8xzEFnYXdWiyHIVpm3gPNfw4
sxOkNqrDvWf9OP0BZViIySGGiegIBowmmfdBsClOSc9j0q+YZOs0FKz1v2EJM438
UB9PMERmxEt1u44JMp8yhIYe7GddBddaq96KlXuQoAWMDPi9WRMdeuTMKy5Qi6yw
9Op3QHbNmRrorZw132BZGRuWQUt9VAPw7IQ6/sVywy2rldQBTZQfei3e54AKhHcx
T2V8NBTp6iMeXSSIzitA7/BSioOO9B0gof3PclDpV9uecowDGcCtO6U6B041pkYn
W2JDcdGvbDHEDEZxnGlaxp+PCRJq7qTWhSZHZa7ru90qSvQKcI7Jxcj7jyG6KPsG
HfnPRwlAduJez+00qBa4IGhpUVf1caLb/XJSeydv778G0ez9lWi4YfQduoY0/0Oe
3FrphE2wIiPMKLvjS3z5nOy+pkszlLv4fWY5V/6BJshWsb02ymVkuKga20kPkVD7
VETrS6HBSWhjzzHLm4wyg7C9J8oLm+tCR1grBuGwd+8/mIenKCfL1nNKrxmX+Lna
rWZbRwl+fPx4+r1E52QQYVFW7On4OA38Xg8O4vjFQRUuCHaOYa01/yyiIiaxwqIl
jPcxNeK3JVvQBK4e92pnofU9WHBHtmEY50qR5nQUZNOwNgaEROkV333qdNF0mqin
KuKZ18LR9qzHhdTTxWdU+9V/XY9lnb41n227WRGd1hgOckm8VXB0Y8RU9ujAUrcs
it2RVgd+iFMEggL0czRncXs4wdWaTwLFC/NskafaVx7IS9N1cfWUchjWVk3nkv0A
I1E1afKDeqxFaRKNHYfT9UuaI38GWDO0Q5LVVSYCRlVhd8HuTt+1Kx5q9nTv0i6T
GjonTHAYU0loCUHjHcLcEY5M5xuS0rRle+aS0LcCivmxgLzM2gq9oBHTqJZefybc
thsCAdVaSb0bgNdlOiWv9Y4+atq7narJs1k6e1z3ul9knjJEUI5nUq6ZKprXKFhL
JgTa1abqeS33JW2pn2KdIgIYki1Ru7EW6gVsgdVGF3xVV1frMFD2k+pysIsHlrxP
6VGxjfD1qOC9ukaYWbOClSZafZGp8pHY1/kqtX0ML5ygaXxwJ64NC7oSBy6W4Rdi
QTUSaR9bBDaw+YgSaDeZpMbCZKeleG55MYAQLQWE5SiNvR8JysHdJCuALofKx/j3
8w8mXiYLw2IsGsPUl2EbfJm2909SnI/vZPt/nZxGKAwT89NH4vqYErolvtpTc+EA
d3CuqWQSw67bhAp95dIK2Nuez/e+4mmPOsi6fYQlI/XoONOI1FQ+gRfYtelQ7eAc
ZoYvGVyKDl9Snm288z/kwFhYBR5GNz+yqXoC/3WgfoligOj77/9rVbB8GZ6PkVw2
A4UY1/S01eYntWICYvxaWOKygEQSAot/B5iqXwxJIR1nvLD4JDipqQgXaR4uUs3Y
X0aF/KSIimmdr5zjo0eGfwOl8dq81je/HoTi5NdNLQeATsKxldh9B6OoLTmFyubx
8ixHSBr7bWznt4J247QK2LszNVDEK1wN0D/+WeTFdsbkqy7W5AvF3TKjPbvnbGQ0
L3WAWhLh6ZYwnD7CfH9KiZuLVQ51SBrBBWaHfjz+rToBqlIqjtC1ip5E94nL88vo
mXaWMOqFf+qxcyC52OaY376+z5ad6Hwp3gRv1EpLBmHfkst0uIUB3ubK298XBXMp
S4CEdKntMZX+HUJCYaHD1tYfEiroOj2YbSjlLTMVWn990tpRkwNwYJ1IrA0SkX4s
yDtQtbPTDwg5LqbNMfg7S7wvJdDD79uquILNGh7bmdVZvm/CbyK0NnvdAHh9VY2x
dYW4skaQp5f0ssHPTxzhL0/QTIjbwcqMCcBLs5U5Up6qmReuk2EtsBduDFYp9Gju
4IFEH/4/Rjuy1lN8IpfGZxmC6uDaCrU9bgCPdBksqHj+oOJP+Gzu+NSTjTzAEKre
n7avvumMI0jhgCiQOEZJHFMPNEJXhWgOFWTCXL427P6DCa67+/0EhcMBul0WKW0j
gXf+3nId+y15ZUy4c2UWulsno2zE0F7cZ+cOo3eZEytNKWm17Rw1E/37jdTA195a
UnARsaTvo/QUKf375R5iHd+UzlFalRC3vqOqHNHtHJ1jkg88KoLyZJhPclTnM7I9
+6seeKSW/qvWUDgjcfMECIhwEK0UWbegRyXQo2qatOKt7ejeqJAzn0jVSQnaupJN
KLQzTEiMqjI8Ly0F7l+GA9lCCSotofpCQUBtkkLVOrZQXl0dPv+IkhBbAs4mf6vf
pTAvrnEiLoH0HYaUIuZqUdf5zLJwA15q7k08ULvqDwsYNarReEtkeojkfYOBNR/B
I4fvfalDAgCU752gjYv3oQRcUOP6a8IP31WLEy9cboOp2lgo4x8etcmsBEA7sFHz
ZLzOF+yj5AXFHh8GnqtuQf3Y4uJUx0DatYdmrjaI96+GDY695saAYOZKr8XQxrBV
mTyc/ddLyxdZOlFvQ8vPqgDnlj69VIgfNwmVXET4KGRv3m9MB8Z5ewXWpEM45GIu
DfqCC0n6lMH5A1fmgpUyq8DfBAbb/liR21nUP3bfZ3Hna+w4iRSIUuWSycmlvr3f
z8NgGyebtPONakN3R8BPLc4yGZy/lFoU5qU5ki6t9vke/E0FRiFIAqLBjLwDUJSx
2+AQi/M5Gy0YpWlDyzKtwaHFTKyEogY4nzwqCcOuIgwL1TFdWWuDOsVdCdI55eTT
Rm9dj8vrIg71FwQTB9kic5SXX7Jb7Cm55XuN54q2Bp9BE0ZcnAML+b+hRPx77KFe
KyqAKOX60a2oQlcbrA/hUO1Alb0ql8Fd3Z+ZmLqpYFrguWSe6dmPjaunKe4GU8gs
bsGi7aDuwDJEta9vn253dOdvdCUFdcpG3aaqKSPx5SZ/8ByYmmPGnZ4WP91yLx3j
Kk8aLY2KhAZrRfbAJ15GbyXePSF7eEPe9NVnxBOF1FuZ5e7T6R7E7R8lNsgdaaY9
gWz4hfGwh3xgfDfZMCiVuK6sXyOB+n/hMRIJt9DAbHPa/7ZnlpKTJ/2aTxUslHwa
Mh7vjoNaCNh5E1v1zF1aOsiXoHJZfazomTFizjovZ7hx/j8U8qCuCeqOsWgf/Q93
uv2HxujiNQAz4LpVtFb/zA3/LoVYXusD9qhB214xNrmDGcCH3688QeJPBLoLDJ1O
l0CzgADwTtrPFSbii/2j8/7KjFS1VbwgUPQIMuHwz1WrerBC6NNte3tMBRKjvmtR
sjtebyJO/+NjIj8QmOxhbqBU7w2chWMN/X/uwcmdzEMP2THDYDc5ZLL7HKM26kCU
JEyg1k7F+Hs6FTlJAqmD4ExbxjCgXeVBftsWqVXLWqGP2fukOOQA0v6Lk3+guPuD
QYRTswHkNhTiorWOTuOZpTuUavoKt9evDcxwBWNdMP8Db6VpepFszfW1B0zCVwSn
ZcwcPWR/AHnQuZzvb+LtUVid5vpYhWoHXBHrSuoL4hgMBbpePoTakQ+PPAvzVlhf
RwrP9PUA0FmRIGGWmGTJsvfRBTHzTB5IsPEbKkl1bnAJVV73vCqX7kvGl/fJMzkp
VrSqurvsESwxUgLjvzx8xHRYYb+pFezdzxJXyfgYN6fTjDsxzvNdxEZ/yFHWE5sF
MlTfd3GXGdQr19/Sb20rU6XXILgguXuc398/0RMXEotlj1/T8KdruZN1NvhDZ8k3
9/CgblO2y9zFRXzIyKAIEBDJb5+FB+k9kaOg/Mv723cr/zvtEF+4yL8/ueBjILbf
Zaq//lZaei6pYWJk3XbdaJWlU3SyG+Ief8/xLVzYysmvVD2oFeUotnbSLLyjPd4Y
9yyVIpoiIUgQSbBGAgV+cfENIE1FpwKflKkDp0zFxfwKD1YzTS8vuU4Jsymbsdmq
OiwCBJKi4Zku0U9ZtbbGr3EltwkP9pxUmboe0osKsO110Xi9P3skjjUvU0OapEc7
8RD/FFItnNPdKiMGsNDZMFKq0rd/cyXeQ1YOe64MRVnOJ5g6ZU3gPBd86STdnrhy
D4JlSXghq75jpgtknROW8MQ9CJz9fRRto2NOceIL7+rzm62muB3DRQfQgaBXRs4A
oXFuDysohKN0lWnpHG/jaM1Mk42rnCe8qxntFX9DaPTBrUtKK4qZ9LVol33SBDT2
OXe23J4oXCEXrJCwem5Ua87A8WKYlSmlB64wW7UY6hExo7QGPCUvIqZOMMgZ6lhh
dR/xBCQrceVy6En259KuH77DwM5VJ+tlPAucRwqcM722+/+ot2E69A6Rc8Tcekht
PxdSP04wJgBhLRlDWx1oAbf79RbEk/RPxmbm3If+wzqdvnIrTyvPAefl2Y3kOZzz
MitePA4NhAcSDIbIwwqq82qymdjEYa/Zrwz7BVi6iqLEozBCEr9DXFA/Xj7TeO8c
Huug7pvak6tsxEK460m9yiClA3iJcB9b8XL0T5LgcuqzEedMPOBkUHBc7mZFCEnv
pvcC1DNVigshy/BIq8r8DDT2xsprBpnwjqXkP78EXJZUxqbG2yn2a3XY0MirBmc/
NLX6FSUGTm9Z1Gxncc0+P6MHMSOAE7khXld4YR9pLyfr3iUdDhtJ1WjEECJSOhBR
Q6874nQRfkYfqatvkWvgm0oj2+I/LS/hjP+9vtvOuL/fqRhLr4oKZY5zmPH5rLvW
9oKMXtCc3sYdUr5pOHY3Lo4GuA6l97KqYrwwL0fd8/te0ALwFJ6ldj0Wj+Y75wsW
UvQj7ci5aTco1czGP9LCJG2dHnKcbn4lBqun47xYMsnKuMG4peCv63kFzTG6Y1HO
WJE+TqOhiaceIY0M1Jmu0CzzcsgLdmV5K+QfpISc1Js+v0qdtab+sH5fBuyd0/YM
6L+iTacNx1gHDkcgXpqn0Fh2K2KuuGe7aUKJJVWPynNjqSq2PFL5hWXu7CHYjR96
TnNZo0FfK3DhPtx950/o9yEFGoo0NyOJV7u9hppUWlyv3AkNrFABMpxIBVlSREFX
lRQ81+FaSe4PZLplUjMPoBXC9wOdM9J9BbAKSSW351ntdDuxDnW1o0Vr7fd//6JT
WMB2DXVFCyJefWfwEJs2m3/3K4VmNVjxM9kkA9Bv6DjVXkQT5tKbM86Iza2wCLKx
pTrBs+CB8BMh0vNpWtdcdNVn8jSlXrIIh3NjOdBS2VCc14UijIDOtmACF1772x8c
S7RMxnb0C15EgoCpMHKJsP5aQwba2pjxGLvfkw9NUPIKE5LIyoD526i+HBF5I/Zb
oEdno3shf8ObK+hWXT5CIQxxftPB3SYxY6qWV3hHz9fpu2K2fQ6FKpFE1pJLtv/T
S4irINDiuL9QVleV4XzEXK8B1VTT0QXtnGg4zRIKSAAUopT7Y3ERLE3g4DmrZkWQ
O1cDcslz3OlWDHkzRuqJxTPuNgCiCtBmyWnkot88cqe4Xb3F+ilceDxl/cmGu6GB
5qZx4vqYZrgI95n48293t2YubQC72BAeOYkvs6ixT8bjCO0guSCBi07lUZMDKUxU
ZIfH4PxNgcX9Syjw1jBxpzyr0hqsBM0A1Ld0m7dNrNSyeUe/v9rWcb2f0XBBI92R
fQnNV00yfOmNLJqKJeyMN6Q50YTgsur0/VPNpL/9TKidJcAQD0Nt9bCiQx/OloP+
0vn6FnFmJ8RmB6NXw+LnCSkZ96exHogMvdCjeR24F40TmTTGyix92L32e51IBuqn
Bnmmb2RpC7X4i6tI4cu+l4+BuCJXVvE3BE2Z1Gi72PQuw3/IHErQlJTKztH9AnRC
fYTpRgPuZpHCFkE76kTpNu6OhEfahZTCaKAxlMXCyDhDGp/mu3Kmm7fdQHuA4uzj
jsj0qCaL86dU4FdnJlOZn3HReONeHnCiYoNaQdYob7hjEUGwvPQbsf7ylGwgQM9V
cdZj6mesLrjm7VOLieWX8gCAz47at65a7n2FU2RS93ey0Qist/G9tG26fJZbkjlF
1//4y4yT3+S3dHmZzafe552kV5v7YKO1iSaezfFETRBEm7M8hr2ZpzlwJwTzcRCB
tLk6eeADG4DRA7vv12ucg+SI7xVmbESEZuknJyK/VbJp0opYR4gJZkCeXnsqCoos
OZJ7bNLlQpvBnF3ijAIzuMEA7tUMkrKcTQWdId97vY/95DW/cTgiWkdSu2MkQOfq
6pHWwHPLcVjqfYm/VRFnA0rSOdJJ9oaIN4nkHPWV4PpnT3KhZwkPPjqsXBcG6ube
xoe28gJwWQyRqnQ595E93JbtKwNthHk+5BwaYA0FP4sLI1VrS3zIkBFfaOB3lxSr
J9qOHCHOo56/tRjTSLinmUjw+xmUg6lf0fq+KaGcKdEUk583UNQACczTOlY8tcRA
4hUFLZacfc6mc1jZTHkmOyNN0arTwEIP/IacJque94j1vY22bd7hLGMq8hvkrnAI
RarNNFbds/gjNTmGuL7OYbHQrNGTlcJEeoIn0jq4WFp7ogTvRArf23MtssBsXwGL
YUFXWGDFso0qTHrjfiuyep0eefI0tcInlRf20g2yZRUOszmL1D/VQSELfeXoev5h
utYqdSeHwsNYBVWkjRdwJerW0RFHtxkyCvrc768nPhyk2pBf8Jb4KMgKwKqb4s/i
UGIjZKB5bRQq/XvvQaOsbbDvdahjKJ+GBz5S2pDVUIlMtqPfSW13Nonfv5MKSgZI
SULt1sJ1+eTiujTGWGsVUCWCFky+2XWmvkzbM2hE7hwa+s4U+StOR6iuBZoFdeMx
U3fHo1FTaw/2kABfUnOIKS4ke4f6H0BlluWyWSpNVxICK6Nig705sI4QNHAIV+KU
0REGjUfy0lhkma/saC9UcxXPjnKZGNHaIpY4AJmACv/rS/bFKvEgJt/0hAawhEH5
MDpsJjVYvpK4fBGs6GS8ZLlYjG4i61xgMHwXQr7hDJUvnf79rWm5XduV623dYEzR
nVe5U4QtddQtOtOM5uxQg+V5Z25dRYYcuYbjEfPPmDqyaHz4O5EGyoCrboSjH5bI
e1ByTGT83PhAL1UfsZptXFMwAC8TH6yDTLH4XvI01BPXFkFMqTWBShOHG9BC2h1O
3RNd6QJyB/SuasUpQVjFPZz25yrMywpK2TGEhee+2NQb+9KMvZBXPsqUT614EY3G
jwrC8yRqFhm1eJ0J5H6H5qRL33BaKQk7IDKlo0LJboig0L+FU9dWkOPcLsv+d6Ax
oYSdAQLNs/8L/Qp9pxLjuwdVcEVOeJgyBR8Ma1XEfttw+eb/+Krezx5cVQR9sdYV
bwjIZJMMf/wDYTm49E8nIk7sfkhBZQKmFoKUqGfsn/y3N+bORjy8o/m9JOfTae23
T5ZQ2/LdyhW97nA7+P0RCpFR+KdmSqAYqAvmN8Elyio7mVt+OpG6c4rQCzJhI9fp
bP+XF9mUtY20Lq0VEq2qUUGpDHtMLf0iH+ylHgHTnqYQ1t3tSAEksxv9H8fgI+W2
tINApndfFjymQQhSSq8VdPjwmmL5+YkS65wvL5ChSzhnPKI34WVq1Lqf3uv87rbX
zvFz8DLBwSuIidMZIq82EGadcdRVxpteof83u+NlHNQx+O40zOD/8jRUeL//vKJd
FFWHxUjUBGmXSVncOKm2YMk4UCAAUyGfG2JMbXLPm2vcANzbtHTNkz6F+IZCro6v
MgvbIlsZuJ2qFau74NNvQiogXITOzfpvz+7vvKVygCzVSDefSI/clGm2oIU2xIwR
5aWC+Ypd/Ph1w/Q4DaGjfGiz7+0nmUfQPdof5lA0ZiTQSr3GPxb3HAP6u91oiNE0
bTPulBPA6Dxc6iH7qkgVZWO+5lkoFpQoMp8+hdf+Rd/eqCC6w/AmdUtT/VW5moOb
QYEV4aieFQSi9jCzwC2rsX/F+6BoCsdIgE9Fc0KjKM7tpzQwP0dMP40RoRmvXhrY
jxpA8AuWia68VHgTHALmDJfLx7g8yy8Bd4NlxIC9d40/VcUxmj5KnqYdUDutqXkA
8hCFh7gBMcvMRGC5N7SA4qeBBYpgbhcGmzWUnmuoQhnLNKJ9Ui+nnydQg4XmnHkV
`protect end_protected