`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3328 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
sTHDbAcNdRVMi738hx0vzpr+3yG6lB8DP1dtwj0LMNncpDe8+ul94avkz60bguA/
CwpWn2vu/GrHzQnJZN/ExEu0seS/AM4etCj5wnzTt1HcqOXLnnA53riFr/jBDv+v
56Pvq6nRx+aP8jHWY0Bl8HFvdXaT3zv2XCTr6eiSnQGyfVGvwo2cjL8tXgueauwp
e5KYt9EjdEXGEoBnxdZUiigNjoT9lBWPOj8NKdGf29DcQl/yklEikqE5qDD8X2Q+
IJlruCJ4XmLArtkNya10HDSojvDLqKl8O5evo+fhWwSLu9XdkAM0zP2bGGW2fTAo
81Lpf/K5/dFG3LApX/GK4Ovs+AGs1BVhngo1Pq4cqFuST+sfiXo6zR6ozu8C0r4j
Y7qj3aeMyjfVRj9vEyT/bBt49zSUxnK0c+q1kvKNpUm+dpFY3Q1LEhDjUgawuTOI
a5XKPr9K7mWiLMkIJUp+MPU/axQ9nBM5a16v3ISPAVNNetDLl7HuNTLtYJ+X4T3o
QnvSF/Pskcni7Lsvf4vxtzpO78kRbrhCY5ZdTv7pjqWWopYUAZfC8BA3kzZnoujq
yMP+qdl96OnbepDLSPcgA2ZuVIEzN0dp7ZBig2FuyaexdhtUQc5qeX+6qwMx+C/K
bhO+9FNnY2IWOvI9Qev3KaUJ8kk48LtdIEapTBDjZND/yIWdCHxiGGAJozLIbP2E
q99Wx9R1HxRMVWOLBoNJkgLzv5WXo/W3I9iv6Fx0TwlbUETPWDiKHzzWwGxYpt1s
izC74ca+blyrdvQwoTu8nq47bpfLmyFk0PM9S8OCCPXbbkmtVxzeT1U97XrvjEPS
ih3eAoVULFU3cRtzkqqjg/CTntmZDHGTkX9nV9aIgZzKwg65g5K4aymEcaMXWboz
BBj2orkVpiRti3sEgY1o3RMzcvSspbH2x+Jt4gtf1GhSu/tJNeQH91YT++mMSiLn
ihmLf03qiVp1AfBCgMzpuqmc3Rnhm+WVAIYp5DOFI1wZxJ3Aei3xD+Thv9NdwaAF
5IblaVBfyqe9rik91n8DaVFNH+/PVKrr7CA+dnhQpUKL/ny8Y2M2fST7h40BkROB
cNFco9M1yhDjRgjbukqp3KQETlifTdcG6KMaYv/8+Z5JHXKSrB2WoR+K3bGVrQqr
LETcyCmVBdrx39jkWtttBOVBc0hAE9s8lGU+qeoLUZ70377tXGVlLyVWXgCjv9S2
AJEnDCAMC9M1vPPAYEcHcul0xe8ffJkzekygUiBrNCwh7bkJw/EDV7UMco0Nu4+n
MYNbQxSluOt/ft7o620ztjLr4dxCehGMdOfdnfticxXUjaG65lUevjdnHHIwWURZ
2u8JkpHRkPDY/yK3wfz9e3cMlkGhTa7W3kMU2UXqOhoHgpEKJ6BbKUB44xCCOw6q
WyJQ9egwt697P84nWVJ1j9i3LyoMFOlu+f21LTt0GSehQ1w3RxpOkhWq5xWIrH/O
7WAymKVmBDC/Ydu5gZyZswfgz1J3Y1AHgyuuE4b+0+cJk1jiMZxQJQ6o6QlBgyqJ
QgKedzc9T9vYP+TU/+K/63cMeFQC9MMpf/6KRZT94GepMOJxeqk3syOOmaHW63Cg
L7204kFluMocZQqe/tdbYvj3hDpB1eQRdgcr/PzsS9QE8vr/FOz5Yo4UcFl6OwH3
OPpPkNzXRqxfgY4C04HC6kedrsinWxfJcMODvk+feaaYfdCgFd8v2Gu1ifiVqos4
s7daUZ5nznhcPZ/75hnNGQAH1kv8INs6LH0AAh5kJop9KjS+ip1iG715z5vT/N4T
joUqwMvRUvpQOoa1oUiCmu1x6RF26QO9hfcrxgaeeSggbnNOBSM7ATUCNdKBDuJ9
1nrVmM0kJqYJhPwSrCKJDP16xe8A8f69nKnP8ojFs7kdOr8OE4D64qk7L1w+lTWD
hradPQfU39fTz/E6oec+ox9YsOGSyy7o6KpEQhioWxZPgU68Crjb8TjWTvIOwFQY
anBrgsvwOE//6cmHBTgtjgNphXcFKCT6kXNqIIUVheMPxQnSjp2ik2yavGlGHEpA
R2w2Arla9sbvqiGin4M9mHEfpJQWa1/HDo23I5Uz8B0nABjsoddeBUZ59qT22JIP
l8E3JWJsomB0kxnkHsj0p3LzAlM9eNUZY89cyNZV0jtPfp40GZaXjJ/kake28YZn
SVQTQaXr2ZCp9r/1VkSCbT5N5/3QZuRXtYmF3upcoKuOK1/FwZnuVPKDDkMmKy/M
IfHhMUq7CoWwfx3YPUdaFdp+WLQFmhof4hdiR91oJHidB92BTuoawwmkiC5MZ7j6
yI8RJgRrWrKneaM7eVl6xcGuI3FP9kh2LvctBfgmhhj2opwfxHr5garfi2Db+nm+
EGg2JyS3/e+gv4zUK6/TWOWMpLVs9BYveQagos4wh0ixH3Prpx4zeuEpSYQ62+Fm
k9B7BRhr2WAqkgwG/BrJmhkKUjKkeJkBDvf8I/pRmUGfkvMbqsIrE1AGuhitke6d
I1DK7Yt2IFGgGwV414OlsPWGpg3napY7/VY1aO8HnrVMmptSLdkijS7i1gmxBcjC
hghC49iL/kAoUaGR93b7IAuI7MSEPj4uxgCPwZySrJMtIKkZAhWFlzuK/z7MqG8u
+yTJMpd7iyxE/YezxVDAhRisb2f0N8pTFJDgPofkzwNc6CeqRmN5KBy8TUXo4uuJ
utbUeAV3F1+dOzmqvp5FH/XHjyUOcd+7Ezis+INJXXFzHl+4kkyWI4GfNYOnd/QE
ZAoDDtmV0aW70UKDAqiqXBK8s8bJ0qx7wi9+88lGIXwlpLW+OG0DBYSTt1++MyUR
ofTvcNak9EnqxKpd9bOfyyK81G8rlI5WgkTkbGenoGI3nJpeuKbDFIkce1zwBH9w
ruCsBM3OBIWmcXu0KFIq+j3uT9Eo+IWQRJGyFigedh9wOMAB7VLShLSfIIRTyKQX
RWC4HxtIRfkDo+p6k6rV/XrX9ap5hX8iDzheHpJQfkBu09ElHgOG5SGTBAzovo7u
fbYohvi8CpYTvghKDnBReS8siJW41RVyYWZqyBEWRyOXOJQ/BvVbDYu3aqtd49RB
sYuZ7mDNqM3cbmF9VvK36KDv4TZaTz71soJgeJxV1rrP181gyIH4mq/apYnWhQbo
RJNhRGClt1B1G1ZGS75ZpsoN7eVzySvIUXmzdafFf+LTW/2K9t993yY/fO7/F8+3
FAc2Q/N2y9/RJtnXRY94fI5wW1nPsOcmVH9KJhz08AYGQxujMqZjD0mw2n3SYzde
H0PYgubMkFIn0ESpw0qohV6t4xInXPvh1vZJ0AQFObHnKwUTfFgnNTGznNoBsV7G
ZrFrrLYou//m/Gcdj361/Usfv29HuSFyVUem6MrWUi9ZJNc2A6VAqamivCuLgGq1
cddWkePk23gwm2ldt8goshOvWSE5/TvJidgUgPhu6jR/fiz+9LVwfxtBcAZJAKKa
mWudkscZ+upGj0ct7WCiOJjN91cQ//6bAPHhz+zCJa1TZmMemuPe1fWxqLgmx6Ds
IkUBOd5JrMe+8+/Xl/gGsvyo9Fl04E/7gTwrSJnt4AKoTgJh4+b5YkhSXG1vadBR
U5DpND8spCYitAjOWUrzctn7HTqBjjOFke5H31Bi6mCmpnMwyLTVP6HXTxqIM0pj
9X32AhtOV6y71Gt+PXr7+Knx3zCMZzonxoykCYg4g6/JuWhZVX8ydM/WNSoENbLT
lILbCJrTan/U27czD4y/AMcZSgzwsnpzYL2f04XtvxcowBO/GC8vOkSz1LuGQ+Ee
w4pE1Pf08G5J1aXnrTZfmgWhofOBbeqwQreGnY9xlYDfNHKOj4E9F0r5lzQ5VOGI
kmD6lLrRJLnzp2vrb3AS0oaR8i7ed4Dod6GPPpGR/NM1anmLjTsgcvru6aFxjeFI
+kR+VkcAwiy5qeJ+hlCqO1aDDJfNWVmUwpwD5qFlQAWXlEZEAUDfTOIGPXth+c2t
nUIPqHgQ27gPjAumwQO9hxIfdeD2g5pOfM+LyTQGqid1p1QfvAFEtQEOUkyyq+PW
DyL3dPqmBJEkRg5PoEZKxDWxm+BKcLVWDgwNwsNC9e5sjBF4gUQeaRm043ZNb3eq
L04A2+RGT8y58J8A437CYXuCxTUFxnl5FiCq0WjSUYMdP06G+lOufS7ISmalhx8p
Je4Sd4AxgAo/EbdNxNitxa2iUc8NaA0ToOim6auDFY1SCTki42yVyVzu8N0U/lMQ
2WbZIHHYn+mfl10zMy5hZQRLSN1Vhmpvi04DbSz74z/o5yymsHbWpo4ugx8BUTdS
OPs+Q+4DaMhfcuS3nr0vFw==
`protect end_protected