`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
YATj3kULTF7Ty4ORuRfFpnT6YIk4rUPRrM74bVTnc4GjdV8oSnW5PtQkMCLOi558
1V+/wvDfc3y0Z8//ksX8sZm3JZWtrxUppw8c14g9Y7owiwp+JumRtO1zuk5xFbe3
0MMnIxxoTKLhyRJtAxElG8sbx8N21OWDGiOk0Xyd5CqAmk9dcOIbxzMjW/wndBXi
maijUdqS+5KiRCM9+Gsp6k/iEAa2LnYTt4WtjkmDD1P5jZKsiMgFck8WOqLymplZ
ml3TTfn1UlLNm/+zD3SFGP0kABAiUT8NK2xBPQ5UzQ6sMFPd/np8iUZ5u4QLTWOZ
hTrU9OSX7lOvRUo8pJ9vPg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="BzW6NOo8eyBw+CxsNNo4wIDxODIsVe0ft0K5tGuSUZw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
DhjJh9S2BY18dG77XPz3hsiSQ73+w0XqfJhD+f+lIDHHVjOB7CfC8ieNRTexgzn1
5W+qoqOEwenoVQtit9u3XViXJSRJ0wfUC5a9axblRNyD2mUbyfH9+f59nWqGkVOh
ieHxkA/DPprM70F3APxk51m7/gNSLICSvbONgLGndWc=
`protect rights_digest_method = "sha256"
`protect end_toolblock="L7NTNW/5Dqy+2kJZXKczEa3js87UJ8H00YWI+92sDHA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1456 )
`protect data_block
6eHODtGLmq6ccbB074dgNWpdzW45i5jL0Nzx5wwM+RA0eeOHXxEV143NNyQGmZjT
bzHAi/6AyRCB4X9z0c4MjyrZE8GF4crbMH4T59xFHqVrQ4zXCea5w0kG5yvHgpKo
Er4+TXTXa9FsGlVtYMafKW30iRtzKaFr1M7GohhmBlqo73smX+ljPXLwl02IZ+IP
SJvyCrnuIFqq40XS7YiSdRkS/Ta8LL4J9IM5ZGbmzZJ4glta+agQaxNnD4Q7AGab
1k2cCdsME2y6r6ZpvYeCrBNyxB+X3Ggt7WY0i+uFTaFAZmbDyng6dEkxeRpbR15q
sI6FcWT37d3I6aCxJ4eKralRaNB1++Cjpqi638zfMNnI03Y0afYqWzwY4Gw3H/A+
gchlg4vTrxqDuGCnjoARPQBDT5x/Gktnx8pmEChIhYaG6ofJJP4Js1h+XXY+wB3w
aENkCeKhE0Hsup9Yba6vB2hsPJrhMS8RNz13FB5OVAgaWQHZhyrMLDcI2HeN/K1o
RS2puEb5tioz0RQ+pgdh4myTy9VtigOXdCAxFIXa1Srg5a4Uvh+XcQM+QLcFbPYA
RawKDKA+4qBXaF8j2+HDwzj/R79jfIg4jyAH40LdaXsPHqk8hccIUfZTjoxQX3KT
V3FJnsdfPEEtF7n+QfPELzVUeZJFEM9TLjlbz4og6TH0ibE8Fl5wUKnqe1EY2DU/
r16ZlOc0C85/xfdYRc3qqy0RKpnbfm+jF3CLpkJNvpUoHX9vrP8D89X3wr7gRQ/f
3AwsIK1YV4DF+PkWMZxc1HWOzFSx6lnknu/LlKr4jNQK6jiD+e+der1o5DtWkM8x
kIyHR0czwroPvpWHYEiHBrwYfCeKmdzqI5Cc9AmV05WqD6MyqGFDZHwh9Z2+e1fI
jAR9rRHBxxcY91OFXoqqMswk81ZHjVsAoU8s9CPkRy370RW/rWm9MeCG2l31KmF3
FXc7eB0ybjtBXDyOSEJbHiKv3Y7w8qT3maJCX5EppZEvlbx3bqhLTNbhRT+KO4pr
zHNzYeNtBWnG2/+5Vxg0Ia54DUUcGa7zQ+HJnatsyvJBigKAX8Y4JUzTleL1znYd
teaUzjgOB9CIgV0uiuhvpcwBneO9rluii5scw2xyLM2oUG+u2b9+uYEX0G0ZSxMP
UO4G56jCHbX+IGBgDFdL/MdLSQkzWVdY6IQtmYGvQW0rYjLxDqAppb7TusACCNVm
sqIdEhJHAMJyVAJQXDf9cH8JoeJzsrIhsanJLmFIyGgOXHy7PUHgcEtsvOmUt6X1
dpf6g526cfnM8nJZaUWVqqtuE9ifowko6OHyI2VGR8Z1pXAZO0hNqWEg9gksfDww
IiYw2+Cau4cm6wkia5MPVuX0azZ74WyRrqxdt7g/kPpFXAmUPNjWmy/cnM2HMCFJ
CGrGn5VoEkMDw9eooAkSUgnlEK77kfhIQAqw0FkPickRzcAGEvsQ6sP4gBxsVBJw
ouG0XuPEJfIMcHi5EHdiCkdjcr7VtJvOa+aGXfBHe1V7fjmCieVQJI6gFr8GyYXG
mcG/NISB8DZw8hW3E3VrqF8Af6EhUUnBmMR/0THw4hp2CqHDg0nUXbSOQ4o1s+Ak
sDZugG7sVP1i+jCHaDK9WUQzvIRv3Y8ElulFXeC32+oOgQHY88YqVr/QXuc8iWxQ
5TPuONXfi/jIIifgxLxv72B22NJsFgeU4OTm9wDl6n5MtwOv5kWtRosFjosGxjRS
hvwjTQcv/K0lhOr0XE41o55UDmpfA6LTemgbeJisgrhlspt8BTR66t2w/+goaBwA
2tyFYI2cfwQlweU1JwLCxpx3IAisHCA4TvhjrKlzOFQNSAte0C6fDtswLzSIl+/O
COCjSjDF1+J2HIrxhq41sOnQzvGOqgdqcx40VUclysyU+bV9jY7Gx5wYGroTwQDr
eGNCg95VNhYZz0DhudpegA==
`protect end_protected