`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11232 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
ky4SiZwRIlZeVC0EoaoEAwGZt8bUEPzoAwKR/zwzpAyclguGDza7FMIrPUBbpKGK
cZb4maBBLyzOYu2HYSdqv/xPIuN3c1C6tgY7J2WqfDnUzd0dAvBmVv7c5lJ4EklP
M303rv8JAvWxbuTQ2kjmRE7Pd+rWFpjHp6DKICirnvgtZ/+xxbejhoqfPuMYOJTZ
yNgQUfVZ7uUQASlrZliOxWSNf1nUjlg2O9kopN4DOCoxEE9zBX6ymXtw0HMwZ/5s
AsM6hhJ4ukqDAzTC1Lj99YHy2RUzEhcLjiVSnnuqzYOufp8wun03Db1VUUVwoUI6
vr3znjZuRoIaN4rEgGfldkOrh5odmrOzAgbr3p1OTJq72Ev0EjlXVYh7gpaQdXkx
WIIRVpDc49mc1XHJmxz/D7ZZeHAZ7VM6l7T73kdQKKXWaUMsIZNdc6ATj2shWF7e
R45cbvBMDg9SYHsEIC4YiEuez0DJexDEhFKCGlBO7YCyx9O7nmqxmYtLH5/Kr2CM
i6K2LrxNnAmbqHnJyXsdKvtEdAFConKJAddFjltExu7ckIXs5MzvGyF0B/fqdUsL
QWpDunoB319S1gKNLDn5yLvBwCWCysAXoUWckR1lLhYCzhebnQtJriRh3WlLp1BK
LNmX/FHGM+H0fZBdCesgtXhI4mkZgE65ODJhAGodW8DzzpNQ6NIGSAG4vjW7FeuT
r5iy5WAR2UNbD2n3DAMyCj7q1zA12TTzibwKPZB60T1sxHU/FTVFjSTiCl9/IBGK
ljY89lBFUxkxpk1gnSqNOC6DYXjRZT1sSpQX2X/DH1NMZNmxpRwtK6gnPHhtrRz2
SV4ZKqusD1NnznvAJdQ34fUKPLWNaoY0CHuOisNkD70hKacL8SXkItE3SC7ULuFb
ePUpWEBH5smB22jRbTSHbtWZe1LM8HYdsVyGw82GzN7BudnnADKp/9iV6JeyPTlv
wyQHjrKmgT6ENe1UJgxeM75gU6PZkOgQEfUn5TTjKFd+HS8NmfVwdBldN2jKSOuC
0QZo9wp1mD/O5T2l8LTsGDu7VY6bXJ/l5DikcBrg9tMw+RXNaDwDcYyM8EnwQQhr
DypS35L/ZdRhIiGJHdW2/CG1QfRlc1xJY71496kZlrLKKe0dSSg8hgXN3D0voTmo
BOR1qRuggdkwd7zh1BmDJmrybd3xKGY3ElVRheHz4SH9/YV7NVQTPFky7xspCnUs
zgVyCLlJzYLHVGgdGSsTq69FBgLY2si5ikQUKoo/PA9P5fi1thKj5VB7bG11jAoZ
J2M4rORbhMB50/Vet0mmHNCgOUl45GrYnNpT80jvKMVZNzUiU9/qvnRWlNK/nnDf
FoM/PcHSk1QGUjDldNeAGB5pfFoLm9Gq2OIUcHpHMCOKD+pdHLaUVMNDCgsmhPdx
tB6muK6NYQ8vQeewylhU8PwlRN0tEgFvnK/xFnyBeanCe3fD0fY08/EULu+eRSSm
mX0Df3753nvF7CMOGGomQ6oq5Dni5jRVLG4QVMng8hh7q1W5UCo7PgzfCuC6lgJd
UqslKBc8zkMAbSKztkWiu/LXHS9SAOEug7vYHl/BHVx3sIoH1iKf7yeCKQLs15cW
TJBRgCjaifWn7yi6JXEXeagSlk2xYC2C9Z/pgKv7BnI+5lSRVKh/jKiGhPxvg+gl
gYvKTIIQwu2rR9VCsWJcgNjxquogY2wLzXiKXXjaqG7YoCudxTWjWjs0WOmeSKi0
1mlCt6raZWzfYMiqgebqhcG4lOmhdcVzf6PAw9TxnXqtBV9HGulT1ALLR5aK2pw1
xQWiPiZfgakQ04tB/NQlmXNpkuFbwSa9Nj33XYKNZurKCmkK/tyBAb/ByVmgB4P9
z+q33zt6LWAIRvcMK0VRD2C2lsUiT82LW74K0QocdXaDZXrYWplrdSpHpAAH2VaR
INYieMjIChDSobjaDs7o2RIiEKiL0d7i9/jRYe78fToI5T4v6FEy4kSkTSxNmz9+
dcL+dVLayDoQE+FDUaJIIwfeSenAmMec58jgKKjVv6MH9/RHuQhfvc4eONGZhM3F
MqbfIPXKyKoO48bb3Od56iFBmroeYQ5zK3tmREHksbdgFRrI0NDCBZoIQLdVI3kV
ISVCwJoIkzsLvfK3wdsTKKbvjj3jtpyXVtZs5qCCy//ukCLlzRWNHahV5KkhvoQQ
mtG7ZGNd9PFH9VQBpA/GajzvJ5nJzaZYydA/8jO7BsZU9PUVbYxzEPsRPoSnM4EP
NdJ3cfO4PKQean1XCrd/8aF+cK7jeFYLG5A3xDRIOShw855m5MlWT9jEznFAZRE1
GDOWck2mgID8xTJhmvMT5i6z32U2xFVdRe0P8coGJ62siLVDtjhCR69p8bVvatAr
aEemd3BmfnQ8cBBGlb9ryrGTbzTmU9/DKXWzpwzgmZkS6JyPTpM22qv4OFN1TLJ5
QLkasHfVBuAPJezBad+ASr8UnNNqGw+t1BP1I0X0wFcTSPdRvh47cUOEPVr7AenA
uB9y0M4OY5AATnUI37VP/chSieyTR6MZAQ2VmsZ0AjwXdD2vNzuS0Rnl6aUL3u97
RisT7mKv/HbRctPi4xlreQjhE2CtWc+pbs6bnbC9IseyrK2litqvE4ZbTRDiKBfu
OYuGv/5+Gb1cFbVybMnbiEIM6V70e0iBNVoJKOMPNDNdv5MSOHvx1RLyjgBPut8Z
NRSZtc7SqRX7ocLEJHtXvS/ZugFtB6nEQsS8pNE/o17ZykFRsyeXQBnXpiSd7k0Y
zp0U9HkP4ZI3fQZDCtE9xehvQTNeH4mJcBzlEzvpyzvfFlbywitaCgcXGRybcagP
ea/GbjFatX/1c3+ui02ceulxK/nu+luRKY5TW3a3mHO4S3BO16ioCOPaupHMfiHQ
AEBjO/tl/JkinbEWCJ5Stsv7jw391gfDYIeFHO7ujyGag6B4DmazEDDUWEVg2nYQ
QFCeqBKIwO/eah8HN42OTMpyr+OZMxJ+/ngmkznQJ1n9ZanX78WWDBKi92Lc8fYu
8F23xwS3JzZRkKHWebzCIFKTt3B4zoR5tgejmEOoXO+S9Uie7NXEMMc8mjyA2T2I
RaePWLIUMiqqmKI68KaZL/IVaAqUvgW8J0Wbc5nFu2Tq0R5ptgwTQjo4Ejyt53X0
YO0bVd5WgXRBYvThULkEB0dVNQ2lqO8RJ65d+UkgTzvXoBACUvivBRWHmm/HqZ6C
BiJInljb8mcd/c2aVq87CQpSilr6mEZ5la8CoapkxpbiS2WVWeRBfvKYF/ImdsZd
lb401FyB7BgIXj10jj94garfF6Opqhi5ReqNHTFmwL9HGhRlVLeRuDuhvKLDB1yF
I2orIDL+rrI09YwHe/nJNfoEFDuodoNZn8z0EcZQzZPx9L4e1gyCxcWfONl58ZID
VqvRsDYddgJGiCcUppj49tnEFXJais5zJGubtj7xTExFRwnJqlAK9oaXJdq7nAaV
bX+3ZvD1iKEanbBNpyL5PTpnwqTS0NKT64lEYzyJPws14tBY7jtERCDtW0K7MvDL
lql+bZWPBVS4Cb8fM5y4A8WxXlqoaLxduFAx22XSoIQWms4UgT/bBsIBRGtX8R6r
aggukTF4poibqauauCMvkh+mjBeKJFqJLczKiQwgN39XM7J480hTcUVFo04Xx24N
yO5b3URiBmVUrE/Kg+w66PTVkP51djPAcEQ2k/vSPqkW2YilIgwTE0ax8h7gXJ97
+jP0DwkwKMKkSQ6eiYrkWJSYBx9jqFs1FiM8myF+jeEJYG+GHqlTjJfIdMUGGolj
3wyePkap9MXR0KhyeJMVr8qaUI3tFxdVe1GcdOLDabYTmUCT8DCBF6GwynzOKeq9
lq6LgEEZS97LkksxQZp2SPVJxLnYDOrxtz1MC2TxZ52XOlMjwKWIJIMW1NHABse7
EkJLIHjVrV/c14McJ2iyud4ku0kJ0XYEgkUDQcUb0dV9IIApXjFjzRtgOumhloqH
PW+3+7cf8HeStstAoS8x/05AxGSC98yaHEn6y1O8CCLupj67iQ6sV5dbW8Ym5RPy
rqXfn365lcX4OplYdXIsZ7lFyNRS1MjecNwU1WvzMlY2Ggv8JhjMOGdUPaEIqAD0
2I5+rOaIEraWrG+/gQpN6gLCmQhUuuuQWZOxXpyvz3TEzN6DFpWQ9SEyoKYfASEe
YeL4Ibk/Bdtu5rjrjQj29nLOSJ/+Oftf8gLfJrkRK5RvVHBAe338MGqtEPE6WCYN
khN/pn0fvXpDxpHf0YHaljwtzC94j9fCn0qMilOVDiwqPoPG6osZaxla3nSPaVZe
7a91qZlYWhBkd7/JtMVgQpU5cBNAmWHfvIb/PI/r8TzjYUW8OgWbh2wp8p3u0NKB
uK+QGHUSqX0iaR1Ys1HiMi3K2PjU5AjEUMcZa7G0X49zzI+PfcAlm40+VPULdetu
5NEAFH2ErRgFe+eSboXYiuTAAAsyWoEjDx8L0ZkyRzPjT1EGGDWowIonZrf5gn/M
GOHdOLhIcERgPKWfU8fPHrwgggj36H81oAIJz5D1QOskcn3xMxVQMRND3QNxqaUu
YkyaOO/bRZ/Tm7rfEQqApX+JyMFrc3gsJ2/zw+zX2vZaO9OAiN5jtP8bUsrNKs//
TO5ELzJI6AzhM3yiYWW+kwraok4y7cx2tvjzJDvXeq6IS/WiACmNk06em9hAdlA3
LcQYRJzUVMzgCO88R4xJLEDAebd3y8EyyMwI5BHq3AdpAMUHUGFsemzIwcAQKjk9
igqWZDYq8J+4ODY7NdZi0a//ut1HPm3KQF2Vv6b4qcHMFjMWjk/O9UjVdXJaHFDh
IDI80kVZlB/wfAgcrCF4J1n+ev5sfdx8LyeXj+Yup0D0SOphCK/I7EOXv0Y8EbSo
9CPU5ECPU4bSIyaiAdXjDCBVj2mVkUATs9mT9hCqXQULu0eyv6/9k92UJqzGpgpL
s2/QuixXXCMvhE0S26jq0CZ3K/iBrCwivQ0Jiu33ePjwT8cf4mxeD20yjJxieFdu
9M4kEc3poxIicUMbyPPcb79LTZbRwd6B8LVyg3pabs28A5WNqzMi1wckAcn9rQVW
B/cTwNsuRGNAbGsqL34EAODehlM+aSsjIZvuWdq1Qvx4z33JcJzp4+J7ZYbUSaAl
UnIEVs5JhGSQ06hal+5hxQP7r2XV8o83l7BhMWVy8FJqfvTywzJ1Z9kNs9Ma3Mbe
pN34qad6cd3cJiGZKO7k2u4E2eoslsdxSU0WthIxIUIRHm8HcNSHNW9PiW9sIp9l
XpPPXt6kaBlqKnISN0cVrvMbSV4SmJdb/DiKWEt74gEHMqWKqqaEziFzfhE59IOC
+6QJ3r5ysObAxM8+1AEoBAR+V/uEV62eel0wVcMrexWV6p3xuMGEsduhf5/Ql01W
kqJJe3aBG/0A8yg+6qm35gZZaHiH8D4v0fh5e+n3fsvTTLiFpITcaVXl56SVafp3
oLXbT3teYpkKQTk0yYi971lceLzYBKFys3Hs6pFBZhFZy6+OCU9VHqV55I/G03fH
SnFB88Df/r9oXmxKEUpDqCbMaNQ5wA66z0W2zjwA96PXUYCRUpdpdUKF6J3QZSEe
uoHORo3+n+vCSLDMAgancHNUMi8ug2gPgnzRXo+iMlBCJNSKmkJe80TU8Am2xXZL
QSFwhFQlwNzC52RqYALS7BVlWDWcykWqvMRNuh24uQ3Z1ndsTul+WP77crK0TvuI
7kvgxgHDuwl0jBPj9k2mifUJypdIasGGoFPpLM7doMSj0bNPkZbW3MsyyTwn36ka
AnKfdjX7Cn7aqhKnHgSFs/neLkLJ6pefjFgZO9DDLIcyZrsX8fN0wrbQ1DVN/7gW
r6vn9fKv5i2OK+pDAda1hc2E2Tc96PCRNNRApWqI5cTI9Tgy5QfQUf4PkibkEbvu
oGWsLSaT0TgcOfatlz4KnD5iLxupOMOVye44QTgBN2s+p8B9CmR4ETYibeMuHcVi
Th31U7y6yHbVMOfKtdB6QGnsROKeZjw8YwEalvhcdT2orS/9TI+qKIRwM0h289CE
QkognzrsYo9o5Uo4rzDOE9hnqsTCpCYdCCfbPi7V8REcIwbRbVn8Z7GyocW+U81x
gOChp9DSZeqjO9vY66uiw4VFjs/41ywCt2znwyUc+Ho+aGWEsowYtXOgz8SJH+T4
axbYRNNK2v6ZaIs0XAGkbHqymzwt0UzERHZdL2swjNsFF02p8X09dHKOcrYQR71B
wZ4dYjw1UeSeCI4uiznGYiXPZkYnnIVAqmiAPJ/YWXfiimtJO6Ch7zKmtgR4ufZR
eBOBjlgV9G6m0AGG/ATGgt3S0/DQpLmQwMsM45vD18OpnPvZYt9yeRs0s8O/OG0S
ASbTDU3YqDBAZcbDs6s1shJcnKsKNfadJgC5NByzifX/XK2lutANxmb2SgZOlGld
jL1i1ZLoHTS6Dmzj+pSTa6GQo98dPbbXEXbOcTdNSZ8N+aMjxW1b8LJ7vbQnwXTn
d12JEsWbAePxKhZIqbZJ4QBN0yUUfOzWdaDrA9+lZB2cHE7V7hd0Y3hS4sy5wqtc
dcpF1b71l5w5rS1dKciqTzKK1HnmSydEqzhIHVWATNqddP3SFYARN0QmBI1zg1dY
H7jN86hPL720ok823fmYx5BFVtkqggx+HG7QzvC00A/fNXb4lFnO69DyLXpTL/65
UmIMrv31IjebrE0ELrstaUju4vAIk4F7lHRLrB36Uj/1cTHNJRP6McWQH4KTo/D5
gVDYEl0732Bf0SHsTZ0P+o9myCvIxb5746uWBZwhkw75zaNAgmz9LGJSm6QXCaW9
0yEz5LINqESJulhTZkPDtRbzeTEBur66931s5i08NZOT44JIbHeHgDXhK5ge9AfJ
ZkC/iB0QXXulDbdSPDJ8kPwd487Ts2+bh7XF6woRukAIqbnlDoRimI6GUd3vmYr2
uXvPAMb3Tg/E/J6dOjcqhISjLCOcrMguHkmPIBTfrE8r5zNmqPR1Lplrw4pX6s/X
WbzVUTze+/3aDdKsre6uR6WSbLdPGLWY2W3OOnfVSOa5lu+xXcE7J2ml5SFYlvaq
FGx63hex/NUyuS2A1m+LH3rx48QZ1gdVSt9xAp51ZHbppaA7W9JjJY+ovr6PqzRu
LgywpbU0TRjrk1tgpkEVbNUzO3sirzy3To8KsBWq9BIPPMmwwWXazjy99sRSoXuI
jVXO80OXFcZOmrQoeI/l0AZRj1eJRAMpLObPiLph+QfrImUReB2MK/MM4XNkPy9V
AITy9xv02YJYwMD4/LIT3NR8ItUdAGS/tacw0AUN2nmGS73Tn4gSAxKM4oVJTKIX
CWuz+3M2i5feHo5EtNu9B5Uj9Eu65BBASJvaT3A4mwKHK5WIJGS2dlBliup7+A50
dL89Ftprk6lKXnpivS4tQTr/I/sLBPKxPdJf543zIpsLElTyA+FZG12myqfjVbgD
DP4sSn9t7GLURX0sa7RsC0/klxgaZ7PpkkoymYk6k/CWHf4MgQvgJuDjAKm60CV2
q5cYc51DrmkRIsoqFBmka+un8FWtt3JcN2UtVm60ME3F3GPdwGiFKAvmQbx7TLz3
heE1pwO4qJyRQ5xmgMH4ftzU7/olpYBrqtEjF9xbOqv2RKwNPpEekJwlzhJMHW09
inlUVnWY7Yr3J2g5Sw16p1HjsDhlutu1QSZXbjhA9T5NT01AtK4RoHvXrrICHtWc
HvSO/+oVn6YneMVitSAw/UUfsypPIUwx3CULbXmbX3L7oneW9YQwM7Is1YZ2GPNr
JP+H4V+m9vPjGRsGPfbIvrInsCvFRUydN7qt3CGF9CpscNZitcZ52oxwOnRCv5Fa
9qe2gAZTsnIiITS8l8Y5sNk7hH7/p9Drvrdj6zG91NphfeDDcOPMkSCG7TrlgAW4
EcieDUrRN+6yF5mme2tI13p3CBDB8A0Cjibio+yVm2QvTFYLVqU+wXaQ4KOqwSGA
Jfc81WaHGnAHsH2JFpAoqI0h0XZessQq7fWUuXXRjdbYfg6CtxoKQGV5b33otV2w
mKuTBxZOzd62OVzH17Z3909wlCC7jjohpYqIocGOLz0AHyvJYX+fKh5F/cDR3FQQ
yTPgP/bOG0zXNfvolm+n5llJTsvcQwrlpRWX/Px0C31BxBKDeR1JiQcmowhq0unl
jeKa6rjGrVj240hJAIVVIFopWOblUJbldcq1VsYTi+7ktDo9E9J+YF3whPLP5xBS
L6n/jBvlhr5MwbT3Se7W4Z+XC/rlkFjXPhBFdQ9AtLlPX+tdjcYNA23zdTIPRwED
oNYW0g0XaXPEN6N4uWbUIkUHPmkVGOHVETbpoLG+Mq3GSw42FVg+uqWSDYGxcweF
H3GrDE23P3Fkg2bI2lQvIUnzCG5wwSFOtu5/ltfTmCstaaS08DqFbm94xqu6Z2rt
NpzO3gu/Q3xLO31ZIy48bI+rrTxtFDgO3fnOb4n2i1GEDWne33mEHAdlarbfZg2v
Z/Q94MQ7fV+XFWlQLTiq14mmwKE4uB91euZuzGhfa3q/dGuh3IjEx//XE7Y35qry
yZ1jGu/RF962B+IbLn/JJmATSYuCymI071OEVnzOneQ0x0X7dStJn1GPplyF540Y
rdUIWNvgMwFKaihEdPIxcJioZeYFJm0UDewWbWDUvou4Fh9wB1inEFULztofXvT0
KRXWkG4L3ctL+p7bxwNdBLArqVILtmp8ZAb3NWTixRVZr4mRUWJpyoOD/PR8dHgq
HiwOiyta9AI8+gcOPklTsT+SmTis9SJjKPe8pvzvcDwSXoEK/Dohty0RkFCkphks
NGwmjh/JLwR/avgm0KYpw5PJSEUvr+dNMQn397VV+YTHV21yrQCNff5EOuUC4qBn
Bbb6nUAGPILC8IwFjwHkwNGdp6h2gzzDJ5014/5ZNHMrCTsR6J2BU1hD/srQq8sh
1Xd6Hsdp+qajVdPxYeB4LQ95XF0CI8X0BdhD7IWUfqRGgDr4OhmXmzi3bzTJFS3/
FK3C7Ds3QCVCERxMGBdaNHZLskFbA7rIJzI5LEEEj/Hl9KJn76HsF9oPjVroMbhE
PgtCh6H7hDcBrKm/NwdwLOz+BTS+DasABzTLlR19F3s+luFgOBaBO0NbHta94Uds
DfsBocIWXL3VXgUB+WnU7OV5qVRT1jamaOdJb6++MvU2iQ1lFg+VhFJn+ITT8hop
b+BBUjsLtUF+nJbLZs6FpQNqWVTSkWJy4G3QTY78TWm42JVOQZBhZW5zrsy/zyia
DS26KhjYJHnpHw+LJOjE0E65JQmG0Cklg55tG+P9BV9alPshwD0jsWTL+FBQQeUk
hRTUsH/IHf94ImYL7+nHeRohanUrzroe012Xs9osilDh6PJB61DRYHBcRtiXuov4
oOwqZN95dbA2UdpERgtLZ1gywxS2P0DnTQUo26/sB68n052VWb39AAkzO7sFrIMq
1MwS0n7FOAWKwviIDgt0isQ5xPjEGlv5tVrybpu7jOV8pKaf1kKCzIrvHfeNJZh6
hvOYzB/BrEwX+yC2tsa9eujV5ebBr7Lx6TYL0krB12k+Q+8RzKyYyCW6G+OehOcs
hsTCLaldxPkPk3x0izxkRDiM7oEhwZC9L1rgg824K8Aib73u0gqu7h94Hk0LKQ+5
lEB3go1A6cqYMgZtoQo/kKj4vjjmqgJqhvNd+wr5ysUXxa44jAp9bPD8/tKEgSTI
mMcROOabVyUb19vPnAwJmd8e1Pb/+Tj2auBws7A/BCQUbm9rbJoTpZF68srVIAC/
w+5pECJ/bbKrpx8ewu09orjv827kgCKSPlLQdHWnzlIkkd8rd2LAxbycU0L5FXKx
51xAUkMa0vacJlribkLooQMByS2/ygL83mqjS1pXjZzVAJ/hP+OfEHyfa1+h+7Nw
9tbNVW8L2vvBJnbiPlfz4913H9lz+6/OYAeGRscuCnbvHWA4k8veHH2xYoObH7zz
gDX36k8v98MumYKNnzF9ZbmUqbjtPD4ICYKpmwI3uNeoDRhpvv2M7frR9dqu2n54
Q84FnZyMZf2JdATWBlublMSsceG7WlYOKdo32YVKzxu3ec80Bes0m4O/gXKnUrdh
256nbaC7YaytDjG8M0W1/3GZkVYsWD/0ldw5JZTcAZ02ZfNuzcNuVFaHkKV7gnMG
3nUTeOargyxhPe7MRasvPsOyU4Vb1keoW3/7E/obsalZJXf4TESCSM2wnl2ECqpQ
wgG3MkT97CmbJGwgJN0Xyq8qgVxcjQkmTZlGboRFISw+p6k4aAOUIEqaWqDe6lyo
FyiHBgGQNhnzD3XCzXEWRNryHNWd26l2rhn88JJFxwMd7fuhjSJ2BWV1KbZC5teF
yZ17K3Zq4g7fTAuBa3jWluE8SC0lDV+TjcTJe5ufO8qNLJS51TgBcwXWUrJ7uBWx
izcemQ41HKjEGAmwEg4xCs43O0I4w/RJnYE6qKHaeTfkBSfJkfBpd7fL1A/ffkY7
fVVr9MQ7FauXhSsnpELbQmw/wOKyjRv0MdQLtQo0Vz3BQEaZvl2hk2lm7wy/OOud
0k3BRDMl/5Zs0+MI9ZJxrM230hEjD4L34iX1yQ+RQqJrGz0ByNTwPgClL+ID6YLr
uLMUL/urlf9HKkwtTGE0NZsYhF7VThla9Sdh1ZOJy280BNHX8hFZcn0PFuhvJYuP
XQH1aF1c1SErjGD17OApY/PjYj1wJg9mCevzi2UEYuka07VSOohyvg/Eb7sOf5Ow
l1v98AE3ttjtsn0IdtByfIeWe4p4hkAiQdtfhYaRNhUylO3xIx6RY6O/Mc2uGWUp
oiwmdP2xEDU2e1ar+tpIjgMPQURV7nWCKqlB7DE6YJvbHdlMNzNZ1hQcZMQ9kbKI
kwCNDJotMr6W/3BwpNINQAbXtU+pmYjfLi7FfxNjT+b5UtLP+mS2TtEWgujTdHIx
hxZijheIxsCv0WZv3RFTDArDuzy3evrsxDYjEFlcfdnbJaUCaofWqB1HCvXdwls6
vt63S34E632A1bYGgSVNB8JIW//IgEcX2xpstG9bCwZJ08gn1TL6aBzVeq2woS8J
8OZ4MfrNKBs2/G7TvOwYA4Bsn2F7c5IpEczlXeeyWhxYLJ2jsBt+r5Iu5IatkhKp
gfsSngwC28rgxmvpM2/jkeDwGao4CWqOqtMmFHL0gfBeUXudSNlazNHYv7hK/hS9
T53tBkzHszJzy4LCJazG5r2a6g3Ww9tUnOJxQFQk+EHvFSVfgKfxSyMnHWwSvSb8
cpwd/EgfqMqWUcZO+BIs3imZq3YZVgAfLiFwscfN/ZHejN52Y/gGo26Y7q+LDTPf
E0ueoU4uhZ8Z9c6mn3WRyH5fmwTCqBAM6FWRYz+Vvndk4IbQ+3WSCmCCZYcThdDb
v6S2I1k6w8qIbJ4hNvqsYswm1Z4w6gw85nWF1cvUcFtdcrR4WeqFIFSEkPboOLAn
H7YDxWJfEjJfs84I24574iw9Mzlmsc2+TgO885+Q+MzUY6RPi5+ddERb6iGJNZ5E
1H6ja+oA2J4muhGloOLlYFhvzlqryFwFmWUUyhiT+LQCR8JICymkT7oID2IX0pqO
SIP6TZR8gQjaDg+xS/Dfnb8BBtItRt28NmOnPx15Sm7a2Dvkc9ZRozQUu/717SvU
hNf6p/f3DBPzpbGZuph1dsjtANDeCl/9jUm1pz3f8nbFIaL+UbNcTidM1CIJwYDC
gZfC3vPqdk3OUJmdJfGYrFny9JjVjT7TGQZw3lmOC+AxgV8pvtT4KZ5uG1inVG5w
congRqNwean0KAqnkcYTZpniu3u9E/pBBqZG7/fs6umNH1FQFZDzH1QXS9x+h6WE
QezwHkTrFWNh7IU07Gyy+H9gcl6SOZXDZeDylegq1MZzvUTvenJYPMcVnrGz3EqT
6Px/xp+p/VXagHIMNhDcc8UBTLZJjIBMqhOyhqSRvA+AZUhpLZ4gZURGQrVlxJtI
oZCaVfbf/N0T/lOh8xsezY4a46tgHMbZUJSi2y7N2Qmg7RSGI4043GgOvfQeyrDJ
qek9tyk3s0MxAiybWSMDcNOqKO0iLi4g/EzACyz3r7YvQ3gKszBRYouGntoLiHW7
gMsIlkKCG9LaKQQDAESQCO7f3xUS4UX+gDqAJ0n3Mdux/B3YiKbFE7uvZlyjd1eV
DtXmk+ovKOGHd1fH0Jjk5ZP5jN6rO4pjQmXw+FTtNlTGrhHtyf54q9rCaKBLX2/8
tm8QpbGwUkuLdQ4fyloGTALboOCWEp5RQuIbu0w4aIAhwBUWhzs8oj5fDW7eD0cS
TRLK3mEwzuWAacoBzlaB6hYfrgcn3t3pwu3rvQR0Pu7RJfOMYmJqIdtSyQMTOiWI
CrxvPaR2/mYdjclRJlUTm9zNK2IBnDl3iUOwJT2rl6aGN/R5yErVGkX5ovnKz+MD
NpeVgyao9ESP1pyY8oruCjUnVXL64naUXeWA/WJY2EWiI0Sh4n+sYSSqWOwmX991
mR9hLk0AzrT5aytKao+RcUg2XEgpSMotQPJgdiSL6KZZ59kMlprrfhUT50B8Zy4m
sAuvSWPIAyAYG9EkBg34RCmbI/w4FeB9ok3kJnr32EtzbcAyPrk25aV/h1rav8Gx
bwsVbKUAZonUTNsEgQbQyphy58mTUTU+iuO760KTRSWWkNO2z+/juNJdmFYeaDYt
Ue2K7ot2GeNPy6L/VQrBsqEs3XNscNvaSUiFQgHX+Y78EwqnOiVd9OmOOezVduSo
yjLEEqSfEf2hOF/DUbReYa7TQWBKXoM3Iqm5eiROvSZMoVq6NQS9f5fR97mn6xPQ
N/lFE2BAEG9vydSkJ3QFmSaqJTnjGB0r1AMMpkX/x/TLXkNAhjXCgxsLAPvT31gL
B92laA5rhUz0lc0FZTODVMPhJkJof5qaDiKDHKBGWPU6h8Cb3LVRygdR/v9fhv8M
879N3Er4MQg+CvvGw7OK9PB95N7ytZ4rBS+1aB7Jq077fN59lQ/vntFI0wNJ8Ehr
J2hoL7dcs2VhYLLBiQ1kE1HONBfQiL23tl5/ab7KRsgjf1wmzRiRcIL9lXLOfpMJ
J+LGCt232cgKKj47fxD7v2n2kPX43ChQc+xq0qNrbveJRKcuXDCjoZGqIqDMjLM3
+5R7qrn0ud6p4/aYGHymUH91sECiRvh5ai/VjT7OM3Np66+DZfCJy2A2R7pFclJy
pu+UDG5rFuTcd3CZPBg2DCUgYENLLa5gVYvHQZecPROp3vSsi12ow25A9cnRfnPs
LUtEB2nPZ44bkvHntu+9fmCt82v2eWZyNI3r4gcBcTXKWF/d9ekYD5VuuHjnQmAv
hGeIpBU4lPQ9GX2xYIAXKV94qYDZ2Eh0I+qAsiI6yWKoIx/x95FwPhtecdC3C5Bf
3NfXUGiZcvSW11ABYcwqu2OZaj6t8BvZ0FZm0pZZtsKOfGv6JvuSHtqlkblutQMj
73GghlrKgmel0yl+ZCmrBWS0HkXISPst8KJGFWge2w3n3Eic0nJ8yIOQ1NCvWPFq
EWnzh0CFF2na1f8cJshyGMQMJhRD30qSxjPpHMjlOGml6L6MkSixbY9pGL7MeMD3
GjgV88rumlUYJPPP3wiyKqtB3xRJSWGrak/GaLzwz4yU78yD9jwL2rlda5CzRLsJ
uVvs9yETaQGSLuGXaxY635gMtCtrSEv44zD9tA0srvl4hnb2wV8nxieIr73hybOa
/E+kHHylVf8lICCTeWsGNU63Mx2dPkbYaazDRMCzYx556aWrhF96SWSF8cmQNx0B
kgqHpu4P8w8bR36zhN/TQmanSuA8nFxjGejHN9nq46KSzoROvPUg/NCzsYzRR2bd
luDNj1ITGm0jr+9J7QPROs4ea862VJJOsLNs/P53pCuHGO0E4PIKMqbUVXIybN/M
mQBEb4ZT5ahQolcV3A9iDDYFYytLZemrrqIFwAI++EPygoMnxWV0XGwDt2R+VZhP
NoocPO7ocNNlIi8vHfcI8obtfdWiD7IC+aWex1tOo39ejXefkmmYnZU/NtBvdWEg
a1T/WDunkBVI427Ey5gzrMmg307NktxpFMUGRqzUOpI4bcpPDSdRn1eGllmkOlGp
fLA/aZDSJjW5qSp4BMqw6OyHgyCa6M0G5gaqTpNSCjXkP/QXs129if7sckD4Jr2u
WIN+AUMz6n6sjqSJQPqIT7iXk6N5371F6S0gbbpD8ouXG/lk0ZIlVO6hixujEgbM
CXgbPwTxEWQTTtQd174dwBmfvvWVLLtDKtwXHQxNO8rM/S1/LhOsNGdS1/Y9TLjC
m6+cHSXeHmDdtcAb9fUpMCPUmw+MY7/nwQMoq0eCZsjvNMlUJ6NbxUUjLC2f7rRt
1EFxBUBLYIAp3Ha/UtNZ1wogHNeKiNvvWSzlYi8p5XYRAMi+4nHc9Jjyyfi+nbNe
8OHWUeHwIbwCfUBHME8BUFvulQtIJol/Q7lmvKtzeDnNxExuYEEy7fv0QfSqs3zM
sJrogOYG0dNsgmSktkhGh+Clmoo4Sy8oxCCkXYnWSQzA0DfbI2ADJEXn9YKhGPJk
zWAY1gPcMyPovlbCkV9Xj6jYogFuTGXLvph0BycMKJpfWV425G6J6498B5u5YRv3
1bCMKhVPiQ/JNsz1++boBKNmWDmfex6DlbR5ffa1XPSDqcKNtSBicdheXJner0Lb
dQJ7OktYVFhDB1bX9WXxrTlWAAEyplFYU29qcmdDGVqv/n8fBXneutW/FyDkSeaS
/zOndNG/XlmPIhfBa88+8Ws4OTs+FIcc/YsP+dFE1jFAUt8CNrai0dgGpiVUzZvF
3rkRUe23weOGx3zkXN/zvYZAtfTXJOXOm4kBAr0TyHCf7RecwEFjBjO49aufOOf0
Oxiz8X0HncjILZOsiNyDuOpdmL+7yMUg3OfMk6uO/OpBbFeZTDVN511V1GAIJY2L
`protect end_protected