`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9056 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
qe1+t0GXQ5YjcbQQEHGgOR9sOTPrYkMBDTKWYPscHh+5P2Yop+NzK/fj9bW9omQ9
cpdu06V+ZsCE8RyykpTb9GrAIX8CLQas9b/q+yP2KwM/3RJZPQlTOsnX9q2NCSRS
sjxEf0Wa0LR8XcfkmjT0xQfW6KkoN73ksDOflPpNN9j2TyYZtdKoR2CydfduLxyj
La6wLYUBnGotiDbQuzyZCLh64d6sNBVlk0wt0Mp2gzFLW/TNQoyUI10oA21ShhV+
Iir2ByMszYNwEWXRPUgRkFanxs4/5RyeRWGz6T+O2prRQf1+lWPh/eqBQMmAnVeK
Rd+EqG52Z2+mjjX1BKatcHqn+LB/1Cu3kOljfWKHBAZOHZ9+OdrL0iQTrMTJS3nJ
NBfe47leQG6yQXCxlDcB0vILATxU2Es1Bs9gyVv7xfJw7z2gbRspYZ0ahhqKu6bt
gO9usoNvbLvTcAkd7F3iPuVf2qjwDlqcOKbY2ratRwETAAuSn0/WdpgpynwfEM03
+o5stbbRd4khYDxmLluwfLdiVIjANUD5NeYYuwPcdl+M/VhLtrhDvQ1yA7fdzHy7
TY/3oUc3/SuI29Tk/oopoiVYcgZuVWS1FUNdRJhom307SJQfBDyFTADhjT0FrGGw
YKsWp0LxSd8FKUEhauJH3HP/dHac+JDPJ+5DOGmvWRAnNWtx10vxHIfeXNXVVYJX
LNpmG5OncsY0cWoUmuZ1LTi8OwsnFLocWczwPtdh5gr/vBzgpc2ast35b+Fqx5rm
tGBDbuN3nZKvjUsBWcjfRtFle2HEnR1va4xtgZ/SBqw8VB6E4BvxBNcHZ37Hagn2
xNqfO+IYnRgJd5IxGLJGvjrk7AF+p3sx+IhBA8dqNL8iZBGm35hXNmSR8gQS9Alr
l6T/GHQqpWdRhSPdWVhGgH4PxKxrze3tPQr7azEF/+G+6wZ6wdjyAFA/E2YfKuwY
Vzi52+r/G0gkD5J9UQImMwMf0Bbcb4wa2sQyM2pNaegI6ar2z2lddKQB8YRLIdQe
VEcxjPc/Mx0xQmmrfKJUaA9A/6F7RDfbtY5CcptQMKOhSLfrLYVNGRy9PjFeyF6W
PR9ejIniwU8CR8VPl514uZqva5k/YPYC/PjANLX0fkN4L3Ab3ZpOepX8f0Fh/nmf
4EgaK7U1MR9oXs3GZCDrwV/Ai5t0V3oFqlP6Ij2Zl+OG93zaeC1u3FXDgj2e6Pun
WwEru+ktq/ejDj+Oxbz77uc/ku3BjzwcSurSdaJXXxwi0b2s0Gkzh+mrwUZLNnpw
/C+iV4dv3Ha2XYIyDz8KNe5jSc3K5Ls8R4CZ5lnjflVloIjDI0L/km2M+Dxhzevt
QFThWOpZHL1PgETrs2sTu5G85ppWQ0x6VAXG4VL7vhkjgJyRQHAe8lKkTHNtxiGK
SrQCAZmEZevU/JUpN/92iNKkcfQBkrXkYVwRb3leNyC7h1blvKruak9iAtOj82n5
zdxXVeWa4ByY279Vuu7FnLU/7/8dBLPZ4PlqZxg1YG5pHQVcWoOY5nDgA2rnr3DW
qBdVCVobl7Wcav9adwWlms2d2DYkCYT9TinwEl80lGk1P4flEG+CgeWnbksHYMYv
UOIurg+HrROM40tYbdsuX3F/n21tuGjELW5ZmU6n6h94GVZIhfgR40gc0ve1P2ZN
pHHz6kCt7qIqM2KsUI0vh6ALHwGoZXOmzjyosnV17mdE7f9XMwopiS2TIDKr8Wjt
AchC4rdIzHh8/L/RUkQhCyYcwFCwsSwLvE8J3gx3V2Xt0JB7TokR/9gVLCrKZ4FS
z07iPk+yZm9HgZZbq12HWK64uz5QgZOQ+eME0B6PzgVtqzpGoKfS0tM+xehxzyRl
gqURBRlBl6uFEdt4yqnaEWsE4cyCccU1O8ThtGfJbd9XpxKe2zcvS4TAtSOMmBFu
OSxfY1hFL1Fwh8PoI/u3tqFiqaj1+29H0LX/VrJqY2aOUMP8BINZTXF9rk3JH+7m
Wg2AagC/VUvYSGPQGuR0nu3P3IQwWs15FvKdMnDQx7CwUJY3b3iLoizcwJByOLv5
JszRO0/JcP1rB+YLm9jpBo+FzeIFT7dyKZv0EhCJ7zw7h4AT2hFF9audI2aruq1J
yohFnoRwG1LkGRGF43P8i4dwCT0xArGsVWKKePgLosLslOmo6hxstf1lKCg1Oqaj
povWoCh++MihNnaXwOx7/J/DEaIiKQGYKfFEtBePKZ3r7JwFQXu2Q+KNqtS5veeL
4c/rCK4WYRBXCcpIbkXR7Gu+CAaa+U86JsFMg3TA+k4IkIhltj591D+RWAw57kbf
fB2/tP9o9QdYpZZTlFDxei+K61DTm6h+6Ce1PkJfFrBhGk4Qtc8ApsVqswoPWSVD
guqgM+DRYUEc9zFbgf4VRwA14FWhMiJx4C2yxrWVsKKg8A7gqHBVXwdqWLKKnlT6
+P1S6GyIX6UwRMcBmJiIiWYl5SmL0ZyaBGiTS853QmnbULu4QFnE8vhwYz5ZVoe8
F28Hfaa6ci7RJXogjiGj0pubqZvZLTxx8pKPm3QkBBt8hXCQLgwfskHZ9r/7xncV
fltT29w9G54oO/HFD8C7RYa9wWfYPyoqUT4WxmFJk1yxxv9urWATCbGJ2mmDWMGQ
Cd8xNoPsqUzo8wOOlBAQMwnwOp0eYpZbztyJOhrSNNCJt4bqIFJUPBluYZl6eRmu
Mv9GAeaApaaoThoQVgfrtT3K7NyLQhT1qG0WDJ8kEvCkRLrujQYzt1Dn7rUKa0+4
IjCssoKSaiwg7cG1nsvrCHOrozI3IXia0jLCtEOLN9zIoaOtNXd0IpY1rc2YShU6
KNVIHwly9Tq3y0uG7J78cs+prdlD3S6VfnseG5TIUZtnJ57Bb97BTL2ckAiWWSDa
d6bIDhJV15mwJXLhHE9MJVZ6DhsQI4QGFSg+T3dxVKm6vZZp4JrOZi9n2xzVogPZ
CiQ4hCWiMDqZuRkSamPQcCTiGd3bayp4rLNziANCeJ/+/P5oAaYLoYueThDoKXp/
F0sF519huT9Vrk5sa1cmqaDgr3DTU+T9mTHqmmFItckDiHrIvJe87LLtT416kEBa
htx3kF2MaCV6jMb4rxiLW9JBrri4shu1POnGtol7OP3WuDVF265nz0iDC3c1ofaP
VtZvHLhrF+CPKq5wEsV3khPN3fFUgAn/XeYYJaYctV6W4O47SCC5aM2eKgvMoBPJ
yZX+Cn5E5VO9UzXV/Ncc2Lhbjpw+FZHNVNW4U0u7/iOW+k+Osf4EzpgWir/Gqocf
VCq/2SH0NXOGUjpjD/m11Bbj+BEzcY00YgkElCQXyxz9PrlZvNAtkjdk+djOM2xe
meQWcyHagq+QleipJvVereB/n+yvIg+oL4Vevm3Hij5A306OF7qiz068S1Gbf1EK
ydJAQpwyGPUPXDf0SscurDWpkCkFf0rhFAzGyoOIaIRyzoRPlpU6EBe3pcfK5vq/
3+uR6B1qjbMRr+wVG4s904KurOh1I8xaYPtduEmnnJuIQ6bPJvaoQtXqTQNrV2iy
RaTnTkKfeQno56eTRYEZVXtbWaw6jQq/1RdD2zdO1v8wjJKMHHjDywgj7UBJwSaT
rzcoDc/QfG4iKpD0kYBVc8i1pl1ufcZtrYqeLa8m5rmrXnd/SEc64YNF8Sg4IOJm
BcmEAGgysBlv89rL5mdReHHvxSGT5kQlcnxLsaMFXaoJw3bT8+4AC6fFXEUbmqr0
G43i6K4GJmVwJGmL9p5Z9M6wt12t7vZRCNROdlEh/5sEusL/EUdPMERs1RoEvQsY
oz+FolmSxdHEgbeEXP3meOf0iafmNIsuqp/2lQLKpn+wU0b9ocjg6G3CYLitSATF
TbWVxxoXH/Z+9BrFKOnWl0q7QubyRn6mZXwAZMFQesEQwgyoHIVK8aqJkvvW2OUO
GHS8ZHVnJfMyMEvoqCcpFDT9ev1FQrpmEFQzfXXNM8wcidxp9FcMvgoPeGHpKQvY
pmYQCkd7IRgz14I79tVdxPDfXZucg38aYw7BXYHpBE3TXvEVBlEKUY3HtWTnAW+9
0rHosy+SLTatyDx4AvD9gc/rwzuTj2nMeEvZgAeARGotPk6/h24RGiHa5uztVU3R
GrAqgRFRs9Wj9nJyShNDJzAWfGwcRcmOWuqp6wpmCh/CEFhExXFV7P8u1Gv8NSo8
br1iGvgWXTd8KiIXnaYROLJIrnNM4pxSO7FF7ntHCu6ns3EcBMz6yv1SOZv4jjZb
hDTbWWAgk18B8QkWcqALPP28V/zWPoahvaA6hw0AtsLie9xk97a+JrznRYgEWaHw
vEM8dAnz3RFRLHj6pYviiCBoWtpm9HmBzqckbtlsjg/FK9s5QpPidd5Hp3nBY5Fv
sse8rpVOsKMIIdwJFVxiuD2W76N7P5uAtgTcx30XyvYcnnTPZHUxk22xWgMcpSqe
fh+F4V0arbmZZcOrkguSAUzxjNMWgsyTiCl00GLmvb7AjPrEoBuX2ENB/M/7zNh8
rytJhmFlhYgw6LmorNzHyVDTemCa27hKdUwnFDXAKpgPM8OVMgenglrtbz1fRAq8
5kjltpfMy7MOmqaLuOwt16fmNEUwfp2hnSKSJO3QSr0TXIOeZ02FikqSdxqTzXtA
4oiAXxj0yN6b5TiyiszTJYDCh4/uVSL2sw8FvC+lBuMRRRGMrvfKHpBE3bd3BpoA
eaviyLrWAruFoOYnVbh/Z1hb03SjzxLM5sYFGNDqb8VTOq83WGXOCfKq0MI/mmJZ
ikRzBes8bk+8XILSxk1lCIH7EL4/+Ml4wwtRiB/OAZumaDHjQzyxaP8e6SjiL+to
qtOHRQOftYBEaT25X6rnNHA+PWHcBI6Xx8dYl060T9znU9nDQ8DY2VmKczPlV0Pv
pH8TyPyRvFmInnr89z9RIPSxazLhxBEcaN6dPmURbs/EU6i4ECF6NkI2Y11KnQkC
ihJHaPYjYJ7y+E8b5agI9xxQWZo6PIHfJHyTYpkFmuRhk0DCw2y/7OxWz7NEwwB8
a5awAKojQzkhVYPHKsirddkvpxCo2nOFbMIjMSNLIHxCBxNt9LasiE2N7renMld0
Id6hvcg9SV0AE2ey3izwz0Q6Fzq4JARh6Mb0l+i/6S/XM0Wr/9IWY5KlUVKeXj5+
htd4KAFVQNdxnfLUBUGX0WLToyCkWskKNC8J25+58VLhKp8g5JxVo7qP4g1UrIGZ
cemq95WUM5vIOusLQ1w0zRcXGNxSoaSYAjbJRzbjtsZ4htOeS9vD7p+x1Jz0y3wx
ZIfwTaY8zoP2vsiME4ZyNf7ACZ1I9SmHxu19p6hvCxueheE+NK9ppQw1wrbBpEfi
iRM6w3i4bwgzL4S5uDQVyWkTLGqowPPHGXIF9AtXLfOiCZ7x5rO4JzlOofyaJlik
qoRyr6KCyCaGRvpdQrMpcjAAN5zJhPGRj0IWSoI1xkH3xVJBWjkcHN8CMqUAp50v
2teENdKJ6pbimSguRCA/A2Pb7tCMpNiGmIy5rMEAs5kSIv1TRapWkitnBIlgJdqO
2cO8EHqUQrOZUmHi6P/RMAnKtv2IFq7WtkJMWNXbtszFL6sMqSznv0kra10Yzsr+
jRBFEKAD33QIrHVQh9jPa+ZYvAdWJN6wE8fRsCFvTG/DCBG03q51vBea08/adpGh
o2HuXMXFGE/UmzpZUxRk8Qs53vpogNS1haOeVedeymxeuFb9t89cTxESTIke80rF
FPkemxwGGzC8Jh6ARa6XcVTQNAOxCYfaOwi4xdK27QBNQDC1jb7rf7rCQJ2b6M+g
n4VlrNlrF6aqAWPk1VFUg+kA+BviwJnry8ki/cGnW7Bc7ASBujdSi9vncg0kGONB
00V2lG4/EOmzcKikZjkTkEtAxX6pgL7xgymJvU4hN7kFngEZpcZP0+jlhbRJVObr
SQF0UzltAP5bQT5tFrY4dlGx5QzvxMT3WGXMAXFOsyrhfhVoyhNHhXUpxMqc2y00
WM4Li/psXtk3JqYYXxUjH4fbUBA7FS1dmD7Oday9Mryy1GDmLWmGuOdY6InY/BvW
nsIaRT4NQQfQ5dmTq2VB3IRDp0rm1Tiz2OEFjN5UO9/Sm47c/EBkzc4IGVI3uZvn
AilC37uVVJM+rQCFWAIVpFa2mlpovPRaxR0aeskz/hMEvl6kEClUUYj8FS3SJ/vi
Xe0RU78EgdAr7CPF+JTM4x7jcmRS7vPXkAnPDBgtlmGIw4LLSRGxvoiU8niel4b/
YXRAxGN7j1rkX/7L1IOkLmZEDV5paNMDjI0F9zhpN0Fd0HyyriTI8eOcBZR93CQa
c2iFiWVMfqZSUCotnAYDW2esdHVkQ6iY5lWdU9XBsKKnqK9kUF1drOaUflcu67Yr
zEmlijN5AhKEOLicT/Em6UuNHOtXiog+9SdoXsSd6v1gSTQ7kcCy+awmPIpp1J/N
Xr6Lnz/36o0VC9vhJS7xQPsuWpO3yqH1+ytd39m3zPaV38UIqEt2yzo/FIsWwVNr
oSQmUgSGWz+fE5FBhANNFclMy/8LG1LdAizGIcQSHmz0hgcO7fseTTh/4PdKFW2q
Xh2gKEXbC3G8zTRmA0qMpjAcHWU6OdmEPk8i3Jm6qTLIrb0+ZGNYz29r4Wt+QRgm
MNOqpc0s+pbE7iwENKb+9ifuQ9b3VdIz4EyNVVg1ix+9Fgm1kyGa1IkKT9tvqw+6
J17PEkhG3gvUfe+icx9LH3RcD0D77MZN2quEyNa1nXYh8j/ivhFqm/eSHrQ8RsXi
IQkA7NpneK6qIaMTmTcLgDnbk1ahFlrxVpwAUCxKTYNAiKXqLoebjSpuEpElNjNx
zZBNsvT/O93NFE6REt/Nn/8fpCptHXJNOu6u0RcOsKyKBRXs0cr8Itwee4uulSVX
HaxyAEus0JJEIm/YM8YI7PZOE7Ni8vAJBEsJmkTWQNLZYPm5zIp5vMd+oue6or7A
2EUefvFSALI569jOO1mh/giGA4ZTBQ1fzZJSmk9nzhwLqUQO+YEr6seF40ZPEe2G
CJQxgMXlFNPNTW1wqFss/GuxiUXXQT33o1ZliSce5OhuFB6GzobLmg6UmjW2/gUu
h2tL0rJwPOc1Ud7Lg4RTxw/x+eyzNuAuVfp8lGK9i/1uJx5iEf0xCTkCGXaGqqXC
laMdIu23J/LsO72AZBE4prZM9b3pYsXvvufc+8cZwRpVMFk884hM6tBI/gVrSnCZ
ed5d6dJzFp1hTLpBYh7NbD+nuhrblhmTBCMJqesgVLszowTSfU/vs3L3Bx/w/yyG
iII6fE4svA+o3esKNd6rDTd7/mzGgTsp004RniB3DThkkY1We6C4rYtE/zJKel00
JWuLYu7Jg7es8Sm68TMJDd2ZcnLIWqO60Ouix4P8FHRqbUqSCJ8JikQlMfcU+KyV
EqnY+I/qV7qD6qlExTtmY9z9mpI2Px6bw6atz9rVL+R8MzVy3ebDLaYleLiOQjZ0
nTQAN9mNp8F0V/AlqLL2z7FVh0riqWEQ8MY5LHumJjKiMIWvj2Wfbw1C1KaezATF
tEtZoRr8NXoIAE6sCXwhxvhGsfW0HNDR0TY+nTHsw7B/Un1DOeZOQQMVxPtQqfCa
NPIb9WKzCHaUAfXdSGdVdMkO9SRq4DICAyKuSdxI+cfgzC7+8mhnR5ozxtaTHocU
vW4+tC8QJzY6DscreExOATTi8mT3w1PAiKA8j9bhXJVi7BNszgeubq+BJStvBKXb
7+9vX+Fp4dp0rqdcKfEA9klSJO/w9UxerKjkFzBptcMAbc5QNx2kkoIOFUsyw1Kp
miDQdRLlGR4WUAZqj7xE4rszAwDNaBBtXOMdXz18TJocgsYfANZ5+OZYJ/qNiV1s
oHM01WKA7/xlw6Vm3mUDB+gCXJl8fIfT48utcMuwhQNP1g6eZA0BoPtY2QL8Jd79
d4GGDTzmDeAb7g6FS54ofyViknbWxm2c/4OBZcNjDUMdHI6er5krE8JJbC/QZfkg
W4EAi4STgNSKH4RKpn1ZwgKa+MmaIiUHxiOYgsMfbgDclAYOIV3uB1FT/q9IH8TS
gKraYGu93PzzvU23iubAiJHv89PCgiL9I0C/WB6lJisBzw2/zHnqm3QfAmAmnSs4
lZeWaNG3YBzNUIU6pXbEqHTRfecPRbm2HplRc4PGRvEG6qonFfyMnPv5h9btvp1Z
9T10pmDjkx0IxHdnPaHP9JpQiIP8n4n/SVRBxNx3oNMLbeAMcrepYnBV24BECBVW
YEC2eOhkl5jNBhN2mG6ky0C4eMg9hz75qO+ZteF+tcKL4pE5elgTD17Z5I5u1/wv
ta0a43BjRv7rvQCheRgjZqi1ifPu71T8jDPRYEr99IoBpf39QgENbh3es5WyD1Vo
UB94TJ4OPPTnl7pGt2FqM4fEtpnXnymG2F6lM8Co7e15mkXW0dvpI3UQS/PwCeQ3
BHRzAcEeLBvS3ZXYIhQqYHAxBtq+5NZ9TuycU2EdLQekTIHDHt1xZ5nyYymZCILU
NqRDp835wlHJUvEp/I294wMKslGN4aNBQ00H+8soQLTM1GtnLRO65FOPjNxr2kqL
qoz8vrdGYjB+Gtcv4E6x1G4OOzpBoWWzHCr3HxoQTBlm5UbGxOv3yEjBGJ1Pj3fF
2S4c31H59wbUfvAa6MD5YtF2ZEgl295gcGoId2V9PN3HLUCM4PGfHltNrl3CMr1J
5DXsfsCSBR3Kss5BfXrb6rbeQIXdt2KKRp9GDAl0UBBEqc1Kpsjr56/B7kMhJ7JN
aGT6Mdv1EYt/Cl7I2zAnbhUuSgaoLcNKLnOo7fytenIjwMvgs/hH67jgBywHdVCf
+x9Mt4eGqGwpE0zqRajEe+E7bHJg8j+HDvxpWz5H09qcP3V7N2utTDNxSYQHlPne
GQJ5Nbxa6njpq83PehiB7J4teN5bUiqBCQJpLUrQeFkMTrP4M6Rhsx+uhWOQKiz9
8a4gBPbWxDnv0hmrsECtjFd+p5OknNrhKykySxbEQpEjacrxp/R12qN7z5W9nF1m
oedFUnJ/QNKnKlLpksWEIgESJlmYEE3POzxU2zSxIAux/ndcVa/ScmwLUuhrcGPA
z7UyBt9cI0U8T1YTdQ9NOC1KjTueOiLinYtW0a5EO1AYxCBlPenK2sYkkLfwWFQO
hNgZ0nzPn79YS9q1NxnryDbiXIh4ncMPU8vvf/7Pt2vQXkVAB9j5/ormX+Xx57w9
AZvADd8UYv5XC78mB2p6180ES/m12d8x3r66D9aC/YG6j+jgnDsjFSDvOU1TusXt
mzK+VXjfgj/6TTV6x1s7qxpu+ZemdnhZnV+jWwy8LJuRIDarQNjcUtKbCO6o0lXd
mcb2Dnhhd20klThsz9IAEHe9TdfL8ObdgdKjrmo465gHz3u81uTbOd++9CfJPMhq
DpTDr4HNkVHLnOQIDo2mr2vXG0B+QTQiRaHt5sV0KORsiNzm0ivPbLAsx/pwTU2X
qfMQtBXxvFgmRqJILTB3fvUUq6ySjjIT0oSO2OPJco/phrQrHYwxqYrM9AUQW6Sz
c9htt5HVNyUcsAunyfz1rAeSl7G2CiyfGLgd8DhHDwcFzQVQ/a+WvZ1IgfdYfMil
Vd4NZcA4bymL40BmYmwT3coVlCPLe6cUg9G6lsE3ddIMwzG68U3fucuQLP1WN+sV
LvwpN+811fWoUPIi2BjQv+c9+/Aen6rBwcEJ0EwgojZK8JgeGvEZylm8GaE698rE
LcgxCnbjEqNFPs/ISiNM/AtFgr1cXmfLPFnBeOXiDm/z9mlGJwTCQTE0OeYKfBHm
oEcwklOknSr8x8yC+yiFepxbuiWjvUlcl6XVVpRYVq8scaeKlPXvzMoZfaj+BDP5
7TcxXeLOHX58MQswwVupXRS/56aev+Yfn8QJRtzkac9Dxt1s79Q/luIghZxQgDVT
wkkgoxT3lcT6XvK5pf0ifUVNjefImTvBoS65FQsGgXJAyl9dJjGgTtSjDucQdFWG
wdsF6dMubfqjkt/OXD6LzEHoBYdBhagZQRJlHVVaF2P0b2+sNEyfoGfYLOtNuMDF
+yx9QLQoA9btQ4G2jOz/JYcjvbsuN8G5aQFFQu66C4VeXfOXWcGbufz0C/nzkr/y
uRLecSAL+P1LYt41V83Kgzwmmb0BGmmDr74VROwvv566+pIljstF75H09rTyt2TX
i02mWKDzDJ6PN8vePWZaTQUOXCSua15/xrX2mrEVnWcFeeFHNnXDz4MVJvbnCN8V
E30tkGDIu59KCycjMDf1c35J8ILH4an/DHEbD2kcsLHombWuLp69bIkfpDNlg3rG
WhO5tfKYwLE/C35+rsnyo0BQeJgY9wrclr4SfdTEX3PB6RnWL7Cp73+8s2r+xw4X
KjjqyiVKHzWUjvXOoHm5OZOKuwve2cuivKLxBFJsfcG2NTCnAyqMUOPbeJasv/Au
dB5YoCTkZofhjK6/h5G3ktY56YsTZ+6HfAS3iArtRC18Rvcpbk2eDgGQIrdqx60b
3SSVwDby26GcnrSrciG8AzKT5/zZxbQWoqbl+QEotugxE01UjArjl6+9yszZy15+
roQiC0MwS70MLTsDlSXbeCalaJSIhvmfV+8iPc3mtEHZFtGo5SYNC/v6+UGrnzZW
1ir8uWaQAMtR0Cu4dXnfmPMeycTrAXeXt/OQ+Kg0DUu32qSeUeY3EeUgNL6fhvQn
lD0kXd4ASNJ6aAMesNf9h6eyF0mNzh3RfiLvMUjR6lWEuRokPhIVplzLlv/n/E/C
Pg+BdhB4meWac6+P+qGOZ62fD18VSKmYrwQVpI6rFZBWoG8/UEc6XiFCBZZYIePP
KwkdkqQen1jALsDjQ/aCWoNXV/imw1xH8qHrI48SFQ4gZxYP5MHdwd0++Y2rFf93
u9HWD9O0kUUR1cJu/4OrUXd8nsdpQYHdkouopaWMRPlDK1lASM4C+6UGDh8VWkY/
Ii+D//T44GN/IkC/OXlfWkYZ36tUVoQGqdRMNcEr1KnBeHWTjbrEWyTH9SaBmGow
OW8Kk4M7s58Bu5HSn82wkXq7/Up6r3zfpV04p6Jx0bAKUARY3F8DZ4BCdvFLbrug
NOU9zt5m0tAFvg575TnvR0sMaTG+8y+r7ljXD4oowrdOdtPwW0hXlx5Js7VSPNgu
tli0GECn2RsD98gXHowPGrHG8FTXmFmwUkp/e3v8oNYSz5MHarbpnw3XwHLpcgJl
wYJum12PQGLreBVnnZCz41eoNCRwzrlBP7WU3LPPR92ujBRAiNNETwKnssC41BxI
Lj5Azyx1yhsD1NzPAfJvZjpRoPk3xIVw3lBgtqlEMfC0vxNL1pzgSt0jws6757x9
jH6FpfXdSee8Kxa2CCMh2bafbt7Cicvab0HqhLyZQVaXtabF/gK/Hh79X3wUf/Yg
y8Af5zNyo7BHfBuw0R2kFdGLnREKKCotD6MrGAtbvkrGx7de6PSykNbAhVrwzNet
aLAIR2Ncz4nfddSTQxWCe1ldbiDRiwOKzfTS58N0wNv3N4uSN/YwqRAc2OVznINm
DbG9Z7arHAPRtCgMCGszWp4otwse+yuQfzlPtRbPLZ2KSWVNdBqXdG7EAbQ8ZffW
U1sH+LHrhf3u2c3ZrC6fxLZVOGYnf+vP74BIZwsF3AZiPheQtbw8BImro7lUc8Er
1ZhilE6SGRkLnMWmwAaFMvL5wVEjbUveWQiO68RmZawmZs8zsHvm3qxOcJ97d6kz
Q3v2vHmU1OJPRU8HDbzVpatlZpQ6g+6Hzem+mMiuCmDifPITD6KG3TpsJ1jDPN9+
AHOp5t5UoIHQ/uBhDQSyaL15qhTs5BKybY0MlQabV27VQtmxxA/KXlhdK8VTuOK8
UJzsG4z5aYMQfSplgTa4EJCAFLO4IfT1AyX+7kXqW440Vk30dBQO9MwRSDigtI8O
o68SR+csAn+b3IlQ9RR42zPHmOCFqykw8tpdk9SeZy/dZrLmEk/B8ZkCgUv1ew6w
Axs7mv7Y6WHz6AwZ0d+vYltnihfraPD+l79vFyXq22Y=
`protect end_protected