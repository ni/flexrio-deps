`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36368 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
m7OJaCYG4D2XeQKzWhbYg0V9U021acplTU9OksDDEFGyW+CsZvnZOCx+2SvRB3b/
/D3a/1OkGVzjPWV500TRuhNR263jTAkZ7YrA/TXoRVN5eoNexbGPf5YSizhqGIwL
ce1gARwuYyrkIqB/wk0TVgb2HYwOLlrXtMkFJx6nuQQ6uxwj78r9G/L8ejdLkqTR
UDmDO4TqJQjfAJJfsVmT0LtxQagObLKWY+RSwrrgOwarD+K7DtjnFKOddETkzOUp
2i0MEFPMCMCfPlk7U4HNyj2tZt+CpkfdP9pOtPp1l7BhRpWwZqy5y1KMe8IIijJL
dzoB5Kx8VbEnPWXRw3H8mwxPFfmeCC2nyRZZXbc4+GGVpKe7+BDJdZC3rgZEV4Or
UAVDmrvofyCtxjQYL+adJZuVuGH6GYBFRrQ8iRKUKa582+5xQteilku5+l1/LiQ7
kcJ7r32qDkis3UO7/8nZMuqlYxc+N89Z8V2qUsTz1//IqVHLK6SeKWscma+7VVob
doIVlI4NmTT1WUWU8Lx4hkpfqOlJfh11gZRNx5ujNTdmu2aOWNUcGdXWv0dk/vxr
Zw20S3Dm/i0sXO3TQ5iJpxLHDp3YBSKzCywqaK5KtmWC12T51XqPWmpx7TXp2cyw
Us8UJRnB2ZL3emTC94PnWVoe1B00LtPK68vf9RhWnRnjMW05ZV6cgKvckpzSw8sz
IzpQdd+4qSmqonCGTIZaCH4sAm0eVsMIkiS6pLaLfLHz1X7A3GWICXckLA97trZx
5i8fVNYNnYVYHod5FT25cie56/pdkmGkZy6I/RpkNtyBHgdnfigq5CwL6sotR2IP
iT8kdgfSgMH3/6kDouqQkW5jsYBuwYjQfjDhUZlq0EYskgPkXSyvrtFN7DAQ1euc
KI9fBD0AdGpVpArHFSmV1Hlh2dD9PxTS/v3Jb32fp/Zi4S0Jab4uC27QwbLP2Ig9
eeXBsexiJDyYp107yj6gKiJPwgBcGMQWFs/mCw9y+XGiJ1a9iYNyy74aBdUDwcxa
6JnKOh3Ej7q5qy7MfBSLSoRsRqUW+gqrjxhFJyDAslYgytZ3GWDbsytNQTw0H7sO
Lck7yOpcqCnUmeN2W4meCEfOaYhZZMWY17fgcRSyWi/Y2RQO+TvqfYw1xu+aGEVp
Safn+wa7XqrvbME6NKLafDlaHHcfc0z4UCjmRTrYGr6AW5wboqRaguXlSjBy1TPw
5ro9irVhTGQeRfIp91Pv2t4JfD+2Mbkebis/itroQPqO3es+tnp2LgYVtizE6zMx
ZpoUqLP8D/H7Gz7oPbjzglF0u2pb22fWAbsmrsF6lgiaMgrham/WO6iQPum6lZPZ
INuBo/yym37BrefDSfw3Z1dQ9USh+aqMqrsRUS+TVn4jVLlwEmGRbfZe/4W8HgnD
XsUR4pWKg2skPC4f1IdSPzvKMYHcSwrizIhMUpDIdDYdQknzNRsSGKNzKuUm9sUQ
iodedzojXQCVxau97MUZZxppi8DyAMW0uBkDMrgvNDz2D1hmcYycgTZxQpkUCe8j
jJB4tCLEWaSDE9xlqq/KH6halteyUYaZV3jjFrO9Y8kKiL08CwEpJ8ldkPxosbuv
aW0VAroqgKgF94z89OJ1o+gWwxN93Erlr4wZnJDpcqJzyiZXtL8onhN1LfY5y3lU
6a4rGAiUH3T7d+uUZ9GFcRPvzzF1VvsgK0xzw264Z55TGlw4fKTBV+JYGbYhfcJe
pDaUTgs6jKpfKkEIwBk042BE88evSRQFRCC27rVksqfRr4+zEuiY9rMzlipuW+sw
59zWMZW71P0UREg4CVkpMAnM1LW7H7Yzw/4rCrWXA7yCPhgfVOxie64YjeGxZtak
NHnRkqJOnQOHk3xejq/NjzaMR6/IMdb1NiQqp2iHIHHjfgD3w0CjMIqzdEDMlsuo
Oz3Wk3Xl5BeYFmKfquYVS9US+CPy323CLXzsCTenccXHYHxyaDET4YPqm5bEfVp2
tvHP3p+RJH3RyemoKIa/QXQWmVmP8cfvtxM4eCyphMS7tl1dq45JLO9Dz4iCfBhM
V8IDEHoblcfK1dVmXvOJksmSgoGGiH1IkpuQdVDK6kPY8PlzN1mUC9WVvjG5af1X
V9v2Th/mYW8MIeOjnA9Kp2+/JZ5oFn+hWtPEGnFvniWbvHQ9kR0NGCySvzEya5kY
h0+4f9WL8rCt7PS8P3fDIVvizLPv8chXr2ycGkWHSo2OY9ZIWCy3so2SmKgRreVd
k+NSfuPX+5z2dMqwFS9VSrAkQhUVe9IiB9XL9o1d81poHZ+kT3yFexnXxJZaLYly
q6NcZKePX2A4O1+QPo7JKsn8NKVPcR/LX6++TmLI6bjtJVmd3i4UbmVYPyQjxxkd
bhSSKGZloPugswGAuDT9QIQhy4uUZOTXsdmctGtPQb/oN5LXoVPjF64zTqBFwpzz
mPYc9ZnI/VwOYHg56ZLPxL/7ruOet12XBqRJ8KXPg/JVq7iNgfz4Ia2qPeSy+J/w
bovg5APqL7ojCpZkq/kHBUVjjI4EoVod0QHkTZD4GWEQDsZWeyUWfpxA9wPLI6e8
cUQAPiQXk6jrqOmBHIVD+JeHLDsbMa9gHVyfNpO2Y1LvIkmiDXu76OcOLVu3tMbH
gPYIm0CU48hpDWJvAqQgKABKqyPwhIhFkMxLAkNlnKKKJ8MuzM3CKB6Z1aVfLAkj
Azet8y2seeSY+XCrtgUB3mse0DeQ+hmOP4zcBLXDLA4d1ZCkOfIX9qXjwhRGXhz5
s8/GvjlUEbwCOkIxF2000TgP3oBSNF2SwowZhO0RLzE/HhmkuKcyYhBlSd43kEvA
D96Paw8vKZNJPB6M3vxNGSuxmYya4hOfdVu8vhPv3A4oIgbvxAXpNL0ME4HGPFf8
yuBY6eRsCAiqRS7td+n5bNWBIfUdRhrk+MqsN7jEzuRm6hvCzb/aCkhKF2CTdqc+
eapPnB7tLyGzJv4aZ0WmbIegiqC3h8TSb/M0I8ttwzmW2gevjGyKD2RJgNVKCPCw
XHnNmsHzmp2SZk8c5TkvKnXP46RjrLsVnOHDOQEdtdmgDvKtwdjH1aQA+nuUZACy
3Ke+5UnbvcX6PQH+OWFb4PsWi1Wvo6UTiCfb6HaihN1Ol5HuBrDJclMm9lbEDMYr
1HpMDgZr4BxubQUCGOp+kG48UJmTvC8t6D1FBkPAc28UKlPIbT3TLYfk0GjXrCXO
Z3zuKyA4Iw7nVU+a7sKH1FHXdjBNjdhvDFyMxmT/lZemiQlTReK1ZV0si+UPJ7QM
bbR7Ot28QxbLkvvU8nJdS2cMeJDlGqx0vZy+GuZbWvmLyYeO+yWlJThRQAh6je1l
eRbHKYlFFFXvKAPYRppDBVZVcbEeB9OHUCs3SxEbLT2Uk/72MkDZK5fsme1Zua+Z
sjNNxJ1JZJshAw0jZN+mqtqVTb/F+CKg3eh3i9IXLrV/4f/8E6PDGLS0CnTvx9L2
hGrBYm7FJK61T0LHKjiYy/ewNRJm6Em9YvBER1xjLf4liJIyqhjfiDobkezgMinv
B7DUrLnsLZ+t+tnWRxEh+RFg4zjSVosnCSXkb8mle6u2u5EawadNeJfBRiVhYVwO
pfWgh0jN7FOb3jKrlSotK4ptAcmgtC43Aj977aHJplGy3xCMd3tgs4FPICcKy/Nr
oMtLGokPT9H95ZHmfx9fLSBRpMTrT4xv9j8o/UsY3E0kzgpftpSeNFMKmXkKbRem
utLmInP48QSSHK4ZFnMxD/ZvGOtlvUCX8E1xk0XdDB5QR4Fb9vD+udHyaEe/1e0F
73rh8ZcwG5q1ac+3jHNALaUUdxR0hWI6tAMTwCCbtnOCj7cyEASHHDbbKatCilCY
zEOlEmbouKlA9ITOdUKe/mey7x68hRzqs7cQs/lRorzkcv/xx0KmWhjBgoeGdhyd
iZPtStRxaBczvFa/mO6aBmx68KitOD/mnNI4gcrsevMGJmcFn8GkTpxVYokAAk+Z
ZQxXF2ZUPZjpRkps0+zNacdtKbQVFqkuGV/I5f2IAhKBZtZ5MqEfMzaA13QqqObW
guIAGt53j08Q6vVIo8bsMBt6yRgoOZsZLpczznqgkYel22amR1xZpHd2Xn8QnFv5
fPSCwY3OxhPxCWjwB320ALxbof8/wB2xc2j7d/nSkkbGcT1wAHrt1w2SiL5uzEmu
8oHLO3x9NO9X+3Q73De6HyJ+ZHJ4nw2dvFnT4dA5/z0UfMZ9AHB3PgeNSzZG1YTf
2xZboncQFr1NZwkRoDHnlYCfuzB5CnsVdeoA0uVLxzMN2aoWO4X/b0VXIsocqoVI
i0iNOA9z58CNKmQT05BcC4ZhlAAmMqUxTTOiFytgQMAh7cYQUdsAiEL30O9vRXWT
jnNkZv9IaezUucMrwvaUNLHVkMEh8s0IVPzEwG/3t/8HT3O7eiHONdlgepmfVKRY
n99lQQ9c+D2eZYz07tKMnHbH5avjlxz/avQ1lvd47OfUoSA8Wi8tRedMgVB3bCev
FOz+bUExPGwe7YZC+kiOUY9nVLHy1NE5p3hsb9BM7GADO7qrTsSfONRfccIVWbR4
IO73o0IT+Ws3w0BPi+DtX/K1DrNIBCMdYPh3mxAXwgMKfLN8bqpp6eL72iVNwKrr
HOv9KS87Slkg2i/ZcA5/5MVwFyXY3FigiE6UWpXg3BbVgjyBDT07B7efbUVLppOP
kVd4sGtbJvN2huKzCLXTR+/Nz1ZgTxaWA4f4MnvoVUUmKVYTz2ePjMBN/N+Hi9sE
QcVjNNATbcvfiqrNoyiMghuYEVQNy8fWV7dED7PQs9qr7XZuWLVGPPnHINf54vSc
63dVVOet0A3focCRxEhLnweaKA0JD49oBFdrfpvF77IBFHMSQapWKDxnMCacjl+j
yfB48iGcGzdt9sasWhGCh8aoEWe8AxbBYsbChfh6fpnqaVJgWK5M2TUbMppSV6ST
7+0lKkeWi2+KYPaSpLgVEg04+Gv4CIKeiMd2zKgjZ2AEr15ogKALpZ0V7JPgavsN
q+5LVBnuZJj1c8YRgpcLsHCSM/ympmer+OM9NvEWpx0gCjCU/pHChIIq3xVhbZsO
/0nroeU/YsEtpkfh5oyEOoUBgZJWhYjPKZrUF8+KR4OCVy3NQsiwltfBsDjk58nh
DjmxP/Wn8sdGsnwcsYYqIZwaQFmh5pDxf1KOZlk1u4t4qCEJULfW9qdu58Tkzm/O
02wqKhHNVo9bjlM4ac2Db66F/yBVBzQJH5Wt6xmURWVnbtDDtcuPJK267CCOnvpt
Odoe/f9bUFtav71c7xYIiEAAVeHLGXP3je9CQVV1pPApktrCbrLOudaGLolega8I
azA9i95MkPOeDnozPcikot1HAMLkwhJYoLFlekYZo66/em8eN4opbU8P1k68gvwl
8t84n7fqsO7Y4JJe1/s69746bNn/nmj5okjA0lW8vz8gwxqgR4EdszvGxQuoVnBy
SKhrZ3Sl0DwZkeiRtmfOCjP7l/QSDnG3/rcwg1E7/stPTcaDJgzPcdYNsxP9tp38
Yr8YQLlSTtN/CriTz1z33Wgz+WZ+EuiZzHiMnYDpU96MC/1AQ6D2JbYQovC2NIXN
fiwvJlNuwh0/Lec/nQXieYzvH59nIRDY3UksWu+CUDvNifccEeRzh4nNAnABcWJc
YEVuJESHHWXz/5M24LpkKTA34vWJgamK1YAkn/2xhiAEH0fe4mChqk4+g8AhDIoY
1lmAFPa/dKwNukxUFgKgrWFRFs1JiAz2BDPqDNa0jZzFu0x607nEYEYH6G8ypAsh
+BTY5fGftH8z9g8Giy5GZosvaoc/SnUmCb9djJFNjdLzuP94Yn9ynhYtqgVLWE5O
VUs6zbBDhVBalHSOmSEgo/S/TLFjNsMcr+V6+JUIbf3SuJ21nyAw+Vcygr4EoZLc
+m88icZJwbPhJT+1INEUC+2mSlcDCtND/zZOwUfnw7lKPzx3pJf8jNoCF8Tu6tlF
SShZDL7CQTaCyBWum1jBB9FrnwTt/s32tD94KacFZ+9dddaspgSerl0uQOW92AI4
klMA3vkO2iBNXnSWGt6b1C9gTKyPVwpTs1y45vpy+HxwqZEheLFnwKNAa18gA1vp
+DW0fGJ/zepqOhaoA5eew0NJhp5Ik6tqt5Ng40cXzNTQ6pr5LgDVL8jEB3GAfKDZ
G8Bf92nmQL1yZflSeVnP+/Sflu6d9fJvEy9gBOkneF+DmyK59CGp8U9gU1ghJq3U
b31mwewjQkRyFDgMvqZhSY9EarHw+PNodE/mohqY6q5cj/wDwImMJKDrgz5gCn/G
zeUinmcBzjLXHHgiQ76l3QbZqvvxKdIU7G+M7EECmbWJhv974HczNZb5toSe4ToY
15arLLbEPmYfaPz3oMEqqL278n5m4y/fib5N/WJjcRvDF0SN1P2CmDJUv+dpZdMX
Zvbvj5myIQokylt95dhFegodD0lONN0yrMuLOCRivvsWxZQgYUr8NZBpO80MY5UZ
nmCBeIrxkbHfcfyL0lWVyOOm1snGlR/4Xg6O5p0bJB/Jn/08Mwc83YA0qLR7/QlN
1fVA+l8KH2bgPtZOWS9AOzoog/KxLDqeOU/NlYM4gInhY8alaM6kGsBrkdRtqDjr
bhQw8ZWH3VIoHAoh81Zh6PNZ75PwRwjRKe5AG/smm96igw7/4FTVmpA9q7vsYGAo
HVlnxOyT5fsSF7K6o1obE7NbxsNb1ucQyoKsma9eOTcUIc+IaJuL8X/b6l8EFghb
DzKGwiyOztm3bCxJnJRLQhsIB9J7wFXeqImLUD1k1CjIDlQkTXFm45u/KWOjwij6
OsNkpLrtSJT8IcgeY5MVCMWlZ67bEt6dOLnz+Ul7qO9IamCy0rnoDv9fFnG9jh5R
YlW6LfrOAteJ5kbfTTBT2THyt9RBKkbg51KxR18XmEtpWZzGJ8yl8tzckQ9JBSWS
/sfsbn3/6NOfXKxSXPrivriZwq14CjnyW37VSZl+8D8y1wbq9uPjsvvYp2oRhasi
0YPCH6ZaNZJQGQnx1VxkYOKoJ3JWfV5G7wg4BEikv554yx6z7OVXMTyEgBTOLqfR
UPDmtGd+D7AJXCoOQGK/TsZCwGQ6xsGU7AAMULhi8Bq+EfSps0aPlQLWOkGl6n88
FkZwPX6m5qact/wA8TXQvrV5Dg35C60ql8nwVxPGt5XDDHtpfWmrkUX2ARg93Kpz
uXdQem7SO/aCDjNfti3wqM9Bh5Xfp9emrWOie+CW8SGH4QjGuRoCEnCmaTReqsOn
siKs2KYZ9lCgnfdV/pr/91erFIyH+8HNsZ1T25Db3YcBKvwXYADOBqnX9QToCjLi
1KnuPN+uqofobaJQt7wEnQI3VoDhXLOrVOc9JaFG9JmahNtEf4tTYOV8ZPN+cT0Y
oCu15afIkAj+dBuVz61X/wFt7wShP5bxsbPg8lexGqVJFUSO9fvAGU9HfNBZdn+a
xTgzds3kcU9ymU5/ZaRfoVJj6vxxtufWn9D2ZMvspk6qknF9fSW+3WGsLerIAgo7
aqPHjAT17jUrghsH5tjmmImVxt/9AoqWFoOvzpkse11IZhlyyZe/iE07gTEcFjQF
j52WPg+5b+dYo/N+pkEnp1w8sGm0WNvXsHiDqBQguqZZo6R2IlLdXulOF0Qas1Tn
ZhQ2d32Wt+eKXhbLaAm6TCykJk7jPPT+4kl+SPaKmSHD4X/kX3d8dDHeIxvXvi1f
xF+Ogt+cPDFcwSthChjFRTPJdtGhGWejFM2VH51Uc8jtK9gcS69pUxxmqj8CazR7
/FjO+n2AH38nfXBk93EV++ZJjRIhntYd40y5u5eUa0Ann99/eWNahY+10dWEZEqJ
czYEZpmfyZn1Piiy+Fn0avUKWRDzl2ip1G9NPNIzqvNqKJireVoWA+G77SHGXcfr
Xr0wKL1bnhABD8Nx/sAJjEi3ERexdu72NwQlXALmf2o0OlA4RRq28/nh/Dih7puB
qIqu1IVSwLpm1IxgSk6Lg0cNtBCsQhLC4qxQO6KR+dRi+rqdPwXjPPOV20la2mnN
jDE26QIlrX1F4D1ehQSYlGDsKCV70/e00wdNfeDb4JmZTyAee2z423JmQzDS0aAT
JbkcN2wikb8xWPtSGMptOAOy+K3aWV0hn3BZBsbjS4zfvPT2O9C+RKgaK8+5E/Ti
uc0eKeE7IAjtHCmQRFTu+YcisJQkmi/Iz65RbieYoZfsRJAcE4Jjr6SmTEFwrQN7
FYVfwDZ8D3bHN1t2tVZoTPuPrXkfEhnlFD93fzk37v1cxBYCESRwvEbWuUCyRL/k
j/PKp6fkGO5jDjupJRLgDR7mtCymT/aSZhioar/54HbCURUwiVWQHuJodqBcTbtL
RBBy0hSHHU2q2vwLMVHIMr5y9YUGyiC4hBjtYGdE9N4EyfhQUvgP9Ebd9CB2+H6t
4iHInTQfX5RecGB8Cn2Ghx5NwZ3LLXTc8CcgDCSISBtKd1UzayoRrjNFf+CvPMc8
lpIHWm7KRD1rgFsLoq41lki5dDjWzWTXQ1qeTkDM0K5DbXzi8Q1lzzSqitcdvua8
j4zqYPvCv1AB62J2HZO6+l3KoDolvv9eUrJAoVc5nPW6jM9DCXoxfT5cEg6buLF4
6saOvSsrb14aQmStc9Nw0iaYab89FcFA1EtTtKsP30dgNV2IyWNIKYWpS//awYxr
SoqJ/hvbMY02ndUKM66/P3pLL+LHMbuu1x35zhE2fKKxfEGN6kiwgIUCz0/vyasf
FZiJ1jlQBg70l8srU16mQaPVhUuY5tgsHCe/FSiX9p1WLo1v3I43VIEoDweem7AO
D7M76GvGQg4akxht/gRMB37lIv2eRArguEJYWEYazfgqvG5s32eHNv8kGcvcRUmL
Rr5mmpTBkaX+1OkZBnT6DSl6StTIoeOZFpZJuTCKY1JybRxZrFW3fKIERKTJOza3
0zT4uPEPrnlHJ1t685d4XwcNtNamXNrevFwvBGEMbSw/4KudW4ZQcINc4LlDaKg8
iWkDCBCi3bGtoDb1y5HlB9qReLtmhGfr33tK8hQ8tPw3R+zfEyogj3mo8dpEG6cH
OUYYl7WLGD6xVFtD7KtNTaNa0YYtIYRPtTeoxDV6eNgRUELYeLOJrCm5wa0zBH7r
49T/8T3SWcX2dhkby+3XeY8dmQUA2X6CHc0WRSggVy/LZThTNCjogwjgXilzOgcL
iKE/RIjk4C2E4rXJEEZUn69eaYkMZMe589CwKK9IO5T9G5m9CvW2zHo3xW5i+PG7
iyVcw4rO6cSXCzS73VdBxXM1Zup1NR/iekKW9MBbw1ayBtQ+BmrFKV1mluqoVNKo
SBKuvDCvAROMQous5isL3wMa6Fliy7oqDIM2fgM8bvZVX0l9mCZy66FwXi6xTrTE
XLiyYmm+D6zk+kiU8rfcaGrljnU+h7IWSAhNSoBtUJYILLSLe+fJhtuPTaTFdafE
PGigC+iC1R5wp5LmgbxC+vIs6T/r1M6rmProSTyvvYg1EFi0RutdruMljkhbAcO6
RkRpQNAv1Mg9TYlbObzXi3WTAun7QKlnM7GikU7RFfx6o+nUtflJFRUKB2mrHEew
MduH8JCfDAByltfNDy9iyw4oD1STZWKLkeJElNNU7i8pF3cV7afwtF2xwKQTeNlv
3Wl73CPfBFwxNtHdH6Vn+SU7ZialFh4KmC3MijUk0cDn7TfIT5wxoqFggLgxOaJx
aEaIBuUpD2tVx5mtSF2A1D+FavPnOjN0B4IOCRsvkPHejgCji2WXLRt2FX4hVYEU
QgIxQ2gGpuNGVhyRY1g59II9Lgl1b7g1ylwY/Fy6gNyqNc/rkdTePW7VB20dgY1o
Tw7zZuKTmr6xu38NIPoAEKsPCDoirnDPw9X7OLE8kig8QZdd3viQHjZDsc/V3I3i
6pOy10UryXy6IqRy/qciKDU5bnEeU2cgh+k/346N119jSonv0xHROlvSbcSlXApf
9jP1W3CrwSa2TwFP+qlkYGQURywl+Re9Xe8H7I4OIUM99BuabD1cgcONiQ4zLES5
KNuI7J0+x8ZAd48gIokXVEuzjxap5R4q0JTudHqSCMB1qlF62S9IKb85KjEcfO9B
aC/uWc0lEY+J/2+OQmNCYcsjYagvCIm2ohzejihDm4aQ4QHPxsODEujW1e6r1Uyz
mgh+l8VPOUxHYIA2TsZR4UgsUfexOti8ycZOsZIrgK8ad+CcpI1KXTI/ciRSHlna
bOCPEb0E76jfNR+hnIhGnFztrm7exo/a0uhcSgiG9/i381lsTkwG6b3a6fWM8bAK
A3gZK+azlazavmGwu6YFDmwAsUhLUip215ExapZRgG6nTInw/VDH6QV4oRvuxavT
PESl7AQuyH4Hs4c+YnOKAeEZbxDNMAhIsTg/scvxxG6oYBCA6/uLxf8ax3Zm9SEH
tbjpwg2ETrvrg6o61/soDD1SbQRSZaSpmVA02GRJt6Iq0UV9Hv1uUSOWt4skOurq
P/MPIGJB/Wl/LHaZJtdLAv3AsD8pSdrE5CcDKK9Ex64TI8Q6dxke0NralaTMyi7P
Js+eJHQgXcLEJPcNTgn2nxnYP9sX2R5/5lP07AAGIoXpoqoX+SzTCC8+Iz3JW2G6
CTyZUiyHobGUw9r1NkqxuF+svQYCywlDFcpjInWtQsdinl5RirE+cMeS3ITqP729
BuF0Si28MjcvSYfa+VUr6yZeYEDw5aAJEzL/Zih8pSxbSzETGPM1uGDSc+nV6abp
oK+wXGyIC2XXGCZG8a5eQs0sIHQ4uW1L0OX2I6c3AQj0M4LXMfkyM3opFP4o/qx4
oLR1e8f4ftd2O0Rag5n34m8nwBWN9P4227IMHSXon1KBfWBy/U9eo4KaSse5uETj
iAHoOgjPS2OrmEzDh8ukEkO7IFKOMVdkBDfOrC2mwr3j+hTouF2Olqsn0/vnyqb8
ZfUSSqsrI6kauzMuO4AkzgS/dAWN7Yetd7uj3vzuGlRxXz82jsEsqyVSk7mNT1OH
jf4a/wwv044OyP664nT9SfUlEbFVtW52I+4RJQyQXTOk2M1oBR31Du8g0ELx9lYo
7z9Ad/826YgAsORyFYvBY7rmD8VBxleaxpjIlswjbeGMvV40lmvWKx8S91mFCyQh
1YI4AkPpxZJSrIi6uXj7t+TmUSiqILA6B7AHgQ8nBBsygCX5aPQIVL45wX32LuNL
YELvaKlhGpMk/ddLeKXLFnb0PnOZKB40eX+lCLrkkQNEQfAESApjHZer0d/htjNQ
8ZuXD2i9sn+gGzwroruCdOEdMclHMQrb+vMDxLW7OU+lQjjvJJpnN3bKkVK6pUSF
5Qv4y2jO2X1tLzqoiWvsLzpWlbsIqUcNlz+VgF9jf0SbhIo40YS8rfL+p175Jx/d
XCws1/FrQv9pdJ3P+878BC/cepePW2hmSqEPqcznPAq/kqPWHFsU/nrFmdARQB0V
Nw0KnDno1KdfTc8KUlZDJVsNnWFKFALn9ep7LLXLP0i52QmX7x2u1yWAI5KXPz0D
FCWjoxqhvgIFD7BuUrU0JTCRbDhJj++vuq2xAntKlw43b7ErrAjOOaX/gehZvW0f
Dcoyl8UYRzzssxQjr8iCH9BqdJRNESs/rk/k9kdqVeUrqIOtchJjIlu1yZWyDM/R
n0Lw/4sS/x9n24Mj3EIZPPTz8iqXO10vRAPmvsXmrAH7sJ2xiaBfCc0kgDmK3cK9
Fp/DOnoG42hOGRYMS7HKPvJr23vlnA+D/ZORQPgZ9zkirQHiUGWkzlopmsaFt9k1
ZOy06Cn2fiVCFmDk6dAs8HFQUVKReGTOqGRXqgoqjL/xYH03Mv2dPqRZ8CzF+G0E
168oNV/nPmcsBnQJkxmnsD06blWSV4BA7HbN2xhAlzyE57wYhbnRJpx7PmcAYqWs
XtZB9A/J2CsZrXOoO7v2JRqzDCpzqNdcI8lBnykM0ie4/pQ8RCjZO2/aXBE6cL1g
cJtnehVfiMZsjZDzj0wXua2OQxkZKNUI9jrrGPINLExNfCJZlE5LIeTuMod11iJ/
8aVm2xH5KFCKjjWZVpNF7pOJsh7lOIUK/yeJWLrI1lOvcEItdtu7lK7tF2t2ECDv
I/eJbdSusVwtewFh6jJlFwFWbjchWDtDjWWOxOU/l0vmzuPb5szTxcICpUKlUEe1
T2RIEpvew5LJ3UGb8gzlxqrqOJDJ9T8k6PhTZnPh+Dcz//FJMUxe5qGPDZbY4fBf
qGwiNp942DYpZfS8GZcNs9SLUKgssWYBBHFxZQQHSuXuWS/gvjY962olCKFQgCTN
X3D+mtYnBGxfRmS9S2qOthgeoibmW8Zo4VMsho5ZoIFsx1MgSO5A0nXzjSorvc1y
On9epkJPCyeNiU10X57jy1kQyKDBd2z/JyFDZTTunhzNf/7C3nfldXBncG3vQHbk
7xH/3P3zJF0fJPSxYlnNCpA/R/924nnN28BATkPncm0ZYuU/LQVr9v2wZLINoW9M
s16shODaDfJqMryWT32j5BeeAudo8LTJfLudWqItbKv/nvKsdzLBHsJk0X6HjAYS
prWkkCXk4oP2c1aMhyFhQDxhUdyfdgBeFQdky9aQoK/5MSUxQTEOH+PkChi+BHts
S3njWtciz6wAGCsOmjIXTMf+ODdD/63f3taRR3LfWTRbs9kehSCACjEsscQ7V/uw
Ll7Sp329lxtzWUkeSUZExFfIjfeVPj33QclxsnAkV8LrxzgHL/0/rY8RhfXVjdyF
Ed8AKUgKBNExc17c//4mY8STJZSk41BjBA4a0rCIH/v8EynnKYHiX8V5n4miittu
bgU1sTMVPku8BYlWmJvJlWGKV8E6PNvguFmhckGRpCF+/Qe7PUl0b12woaKsr8Nx
+KARpFed60NeDYq/Kz7Nts+83ycT1KRPBVrx5+UXFxzGFMe23Pq4/k1/MmeWkdAo
TDXtTAz0CVF6uoCr0rEtnKYYJogtU+96tlmdpbJRK3x0EQlwUHBKP8Y6vLW/elrz
QA8/AjTprK4FUoVpxV/BjT/PoSXEugMsS3rb8G/B73ZC8yq+i4UAaechpt1dM33z
u8gTuELmSV5MYRpOpb+9ksLyaWKVOyjXjIrjFtrYTGpYFtQvaFGFFTwzOtHVa1IZ
MXWUnKmxYXEl10BZd2m3Feba5BduIksFCS6mRPd6STaHWFsnUaRmaBebWSJVofHE
zG4a+XTNcih97Nxcvnpvektod37XtMr61U5AIKqLDJxJgy69O4na8JgQLP6wjzfZ
xoMC4UZEJIyHJg7/UYE7j2yQqFs2XDcvIqCaLpzRSiIMF1NvYbmAYUKwCyYx4QHC
tcleSen2zNq+1uIwBoB5crGvdIe0DcM/qODfbTkYyBXzu+hVamK3QH+hGKa3COSG
7JpV1IwNHK7qU/eoZqsW6nrab0cYDv42d2451IM45x0U8+2r673cv7tOi1YSpAM9
sbbV7l33QyTVG9L56LCn5n75yXbkaTltqSD1diRCqLLz5ieWzAJ6KrDA6jTDqBQQ
Hm+HXwhO5qQYzbRICBw+bEit5VMcnzHSRP2mrfblN7z9F+bMk94jQgXydRBp+CJq
+4BK5nqGHOEjOjQYEm3VK29lDKjWLEE4J4ulYZlxNAqzFeaTblrEbp0uDh1Xv2wt
k+LZwFmxN9mojTR5W2SIOxy3rAcsg7lrCNOPRfo/AXrz+Rf+sB+kYyFOQWKPaseC
J5LqoeFaRBw6y6678k99nch7RQyM3LhItBjjDKLMIoChaFed3aAnwcakByGsIMm3
Z0j82pVU3/xsOLgFwUXKJ77Nf7PGIIccNIn06EmbMGuDyOyxbYktlVdDnNy5hDRn
Q8AMZd/EdSYjMndDwrEe5rnPf4ElHcHFoSUfIWaaWSjygjidqtSg7/unOjSdiRg+
Ul7E0yjOJQ8nFByHqCAEkw3qSeHcYX5H/0+AwVpETMvtUGLUnCoS49Vs/CMX0kDP
theo/E+oRnUrYd0Xi4n3mI033mN3doWh9Cu8U2mMBMnlgH7/Lmau3cablSTjGxqq
jNZhbmRYAK/XbKQg6XVS113AduRLNZ9UTPAiFcBN/Cx3Ip5i48XHe6SUVsWO25Ts
0H5/f/eFzO3F0FqWdBgS+vCkJbql4tL8KH8KWCqC+VJwFugw4MKXTP6voDQg+hRg
JypCIBzybvUSlD88/jTs36FKVp+XfLbs9L+x++5XMLtVVSloCFHkYib9J3aGKOxB
9vJhcLAHQnd5xmc+sfzWtTAnwKQte5fwXvWV2XBVwV7l3sdiRgE8JC5/+qEvzhp9
t3srODksLBuQbGs/Q2r+uHylfTfmxxsrfan7v3Y6L3yXYLCJMxHPk1gs42LR+jhP
Hhtn8uDH/QGjWbcbHJD2g8C+xlYxBd1MyXUEiMmjSMzXrNw2dJMfurSLolgQVEbO
wQK/0wMFqFaVQP/gF0iWYO/6anEsgRlqvLNoOTp9dX2plPWc4hOG0c4ISpkpO/we
XV4ItXTaroIB2u8AvGJuLQgfKM18uuKIZYx86poRKk9pBoIVQ8I8QMCGm+Jy7uC4
NM4+an/Ac62CS1H5oUnjky3n8k0vtc32/VphTqTLbH9SMmewauQwkQNHqOcswgYU
CPbrsdF5ZqWBAfVPQI3dP325Jrx7j38/wxpPROlpxCVE4l9TSbQavZTOEhKIOPON
ki5nu0FXlcAWyBZ22o5nqfewY9qCaEFXxpVp6C2iMQUvEw4gvZS+ulDgNvnuXpQQ
rlGwxWV2ANs1F5bZW+FWiiEuOeoW266cTYUV+5VPgRkraZO0EtTvMu5m6TyAxnUa
B8kaZT5AmiROqaveUaI1vvkKJTWafzvlBMwvYljNBNTP41P47HI7T0ADfIMeTANF
QvyU8H8ENM+6QjZVsYDkUh24LzX0C63eFfFMrAPQ6zI/ZO9yD8mz/itfAdfsyCbD
qMgvlZfhZkdT0l0I+vkASmk0yhiwQ9pRtjuIULZ4O+tvqb8p8ocLgYk/VK0XKFVc
Ui56mKBea45Z6oLggzsaYO/tlwNnj/QdGXVu/w27vHd87S6/LjXx4G4SdefchQGw
VO0lhCuGxvejG51yqjl4amnzhPRa+YfqnFbc6fBay6ZwKYZPhx1kuN4coNltp4JT
8fR4DxVHp20G4vlMLa/si6ZbtrTWMrPVa4XjfIhjtmScs2colR/VY/zLQ8UEI8hu
b3LOHtm6o6ar1Wa3oLsuQPyD//atncqRNyyZ/WVe+S3pXgD7hpYdMo8l0C18TGhm
3MVJrjFlRe+TOTUHm29g38v6uZqVoTKNHmvPqlFJ3NfVDpCb4jjFDw0LDnBjYyRQ
0VmDWEvsa5tEHvjp5E0gKBpkWVEi4uRdlT17XYXTGNcFhJPsDCaUb20lnaMZUaVB
QBxZvkIDErfOqLI2IJpXyemvuGpDPFV1NndDOeBiITmvPh/2hs/tRZH0ABjeUpNR
w88UAxeCcOqUKJD1FhtXduvaSrwOQg8m7i1G8CJiB2F1LpWatCtjD4xoUry7esJ6
+AStMdx0sCXO0eUUs6zzuvcX6fVQZYUqoSDFg2k5Ih+FmSgZBcQQcGb1602Yu1qI
zpddYMoejaoK1O2B6p+rOzdTGezBTZ/26926DmVVTusduqUr2ukxT1ngIhCUwxdk
89amnmqKbZE9bApCPW1qwARYBjU6E3a6PhWcLb8PDitK/NqJnryfApotsZjcqgRG
ik9ZOHVLWj6J6Cy2oDQx4QCMFqTFw+hEjKZmbqgsoXMBiU03CNg1jT3cL9aus7jG
1taTpxAFSPOIzt4FfSgLoTGSSrJJ7b4KtJS2PxehfCmRKXMAMjhTBf9DtgwDExrL
8Y1GLjVYmpRj349JhnXhwZ/TkOh/nHJ8Pc3bUGrz6xPU2DdLgEtX1kuo+XG9mlPT
qOCeC+3cOG7DmTHifXBRm8UOkvo3opoPHQgLDu59rHbCZLr1L4crGZk5wO0pzv9J
DKEBqtIfk4EeFY8+09Ja217Tb3uVaz22+g5Z7+Ig90dtypHy6DpvCrLmLgJTiE5G
hn8SK57GSQuF2KW7wTrFI8KrPHpjoXOh/ARdIwgK5tpQdKfPUeXgExpax02u8Q9T
wEc7T2WHrz3Q9JrHOzOR94orBicRj5I/Flj8ysOvVAToB9D2UkgxeQ458HvG5WH5
+T5N2j/9bedWlFGo09G7xW8uFhcZN3WefE8mIO7szB4+74Wf7QE1QTEk/TyIC74C
KqCZuPfMZwoYPnwa0dhdr+UGAeTtCW8rwZdG+UQTrU7KB/vTg+570rPbBMkOffQB
kRxkx6pnrqSbTWlgZnuOhmgy0ft597v5VmeFqVcSwapaafaqv0rbS4bsffq+xoir
PXVn77ZmQyuyzGSohvu9eYTDKOnChfgZtMvfCkAGVtn031k6pEVANtjdz8LKBin1
uqZA5gp554CgjNHPLIHP6cUIpKbieCo8sVS4UZspjtUrQnwmow5iweA/sHGK/qet
cVSurOKz63GH2YS9AA0Dtd7FaHAlut8rhA9tySYchlr1E+sdS6mOBUv4jHWiPVp8
ZqREYLJ0CadsJfojNgJh8MKnKGmA+u0WyqAu4tkmoshXKbaQZx5jFMkKkeX665l1
+WjbHHXcca7QRtNgh7Aqa5R61mzHfFD31MvLXxmFnSOfwtMlrCEjO8HLsVHLXJmw
FgYgIsAlRlfjMpAZBY/4Pc1qdapRy7G0/G7rKVEV0wcUgdMVmW3NReOmGSA8Ia21
eOk5Uc64Rd+I/h1T12Ndo9CGRSFnJ1bv6z8epg/5i+ahk8enEqVfXr7IujTQQwIZ
8Cv7bXE0bRXdVjql6g2CIuHQEGrnyjEriW1lNg80IURL8PilZM7zbVa5zz19sYLi
QzlLr0iSv5kgF9lEQg7M3Y1WA41JTrt67GvVPGaETBW4ztOkfhFQTaiQcS+YK0Db
ZJ9NA0rzwPu+7tpvJaF4vmlRuev9UMgkb5PDKFeUCXYR9W2XFn0uxPtwAdQaKyjP
QJh3RcHKvmM8hiDv6kZke//JKecyV/Ea9GJfFu8ief9lWUzPep3s8R463ekXnZ91
p4VJ10qwTypFcEv3W3a6l7scIyFnrVUx+IgJ0x7RfMpJa2IKZzzmtpyFRGvSjjYI
AMbSpP0gtn8AYdub+pFR2NkvPSyKLBfV3jlxClGFCRcR7mjE3ZDL3+ssINKJ44Zb
pHcimx5iHXbFqZj5wMbdJTmz032+ztgEMmRYKn9wuL3r4ZakpOmPFsr+FCwBnSLP
wsChEpn+umadA1ydFdIhE1Xs4Db+jmywrnfCyh4k4Y4a4kveNXAWGkqZrJBdEyaj
69otrumP8wUIPuEk7fhaXIPv1ZOARXMKUc+9slAGQ6y/tTFF2KFqcOqOAlj/uxz4
angsIQffpFLbvglUxWJZ7a/uacNZ+zZmu5mOlkkCAMeuw+/BAs+3oqy1W9cYtByq
BvgOSHVEV113bNbQr5bQ+l4sJxul1Z0w4UtLLHDgwToQEMFeJrHUZzg3tGhtGsVF
+SiOQVmNvIGLdL81nLd89EmNe2x7Ic7X687z3dNWkP3zkfRAtFx7kyoZiase4gbG
M3EktW7tKF2v6C9Jfq5p8/2az4nAeY0z5hTBUkVk48puPXvk9Kb0baW25izGS65n
6O7sy5G0LtDGX8gXMH9ufVoj0rtgSR5SpAWlG3IeWVrVm24sej2FNxkAe8WQuF0j
DZl8TwRy/SgrkkcnBeDrsSmYIM4UjXekjUHA21bLIBdmnstxzUzeEgAgWPg//jQz
0qAggb2w3lGMpit6u36neyf1aBLxDmmDH10apDkaj2VfhZ8tURX0IA0vk16wIiMj
ci1mX4F/Q2fujHNYqgCZkhlEprrVywZjlTZO5SZmqAxmuXjbwa1q0toAGlQrZD3I
u9J/2RLygcFo7ESy71qnzhS9rS8YZfS/hKXgqgtVV85pf+eA/kociRYA1LlxN3HH
BIDc7+Z1rZsCjmWl9Ol2sWxwhGWiTMbF2weofOOePEA+0VVRTthTaUmQZOFvXkJ4
qtwkfG+PrNy0X5aHSrxEy1MunZxS8D4tkScAMlLY7KCkw1rxZphNQqH24wX7XXAf
Mku01n8EkpsstfwfUm8dhOoHV8w+C9TJVHhBXLSVgU58agz9ySEbX+04UaA6zWnb
wt+aKFcv4C4XizPbSDo0YlE8aPZx2ti31MQ063ZCJVbtON6AUxYTlDFgVIWu5A4z
Lblb9tCLzhkBMjrLZplFNZ8zIdMvXeHRADHamw1sQRw6doK5UHNAbJKZmLmr95GE
GRVyACC0JlMFAnWoaZ1Zz4/UJzwsHVQOBZaJAm47GzSsIeCM2JIl5/e1L/pJmU68
LnJUzl7neXE1UjuUXTaOQjX2XcekpsSr4s3Q0f2YjNaPIBGuRIXhrH0yrODFk01D
MbiK67299+9eUzolQlYtdIbaz481lP3m1ZFP+QsLC2U5JoU7Y0nDl/PaoX4tBLsR
LhlVgAc/OTQxxT/Ksqqtq4gDeC8TsKJ4T0T/ftRSzzq1yB7dQ0M/xa5W/b05ge09
XoLPyRjqqPs/UkGroQ/8QqJbRKwU8XMt27qfHO3S/lgPj1drerCTV04nK3akRxTU
cp6DmDbWie8v8B/mlBXVK5Mh4+lTUQglup19i4gPJWlmx/DuRIPqjU0xUoQrKNal
nHWMV0c6n617+oD1c77ywV4WCKOwNuW2NgO8W2+j+sTQkdXYkcD8mUiVqvHaVOO3
RVAlI914ZtF5Y2p6W1uYYTpRN+xXZ8tIVax+1BBdTV1vLlM93Id7CfaG08UQhgDN
k0IRe7jZIjR/IMYLZYfn5HlKnBUZJcvdq0ymZJVainw6ecJ6YfGi/HGBdTNQl8D5
AMAq97y3KcwUDoyuncvsJD7mwyNQO08/M1oRdZ12vPJRh+6bXectfZiPHfrz9JKM
ZgQXajK//vy6DnAkmUNrXKzmezJj7y370626HEhw+Rnupc2W5XkmrG+I6SRPLUdK
Ts2cPRm2eUbao/tm5TmH6Q1nP/O763fu7Hfs0884scjMLq5TUUhzOioPhqfuFuCg
QXdG1DW4qE3Fx5+Ue/HyXWp2E3cO9A66rftKYeW86UKZtuK/47shp5nE6yILOsVs
66SpfGQ/9XgPFo/ger82iUO6bmziFDfdYSkVPrg04bnwwDgdV3J4uXjfl7wQOTu1
b14/RpN70gq6Qh7zUdsyyDzvwX0OAPVr3xyNzSBKVMgOKQLrJBi0Fe1STk9jEMXf
ZyX0zlD6lUDryBVw9iR/h0kaPcnLtUHz8ns/y9Agid8PztbbHiPxdIprhGw4G9hR
85UiryFH4CEESwmbPHIVLW7YJ/1kw3Pk6dqmgvaCYetetUr2jcSMAVhmWZfGEugR
6mFBgBLxAeauKeS+ciInLtvSPQuk7iLOZFDo/i9U/Z70ffLWhcMWJZ0zOGkLHA2C
sIVb2L0WQ/T1HPY3Wd39j9MR90JX+vMNVo8TqBtKy8m5ikhPkRQ+NcUqEJ7hUJeL
K6H+uRgkmp0SpQn/edGUGLBaQm7xI345kP+Ksxpg7qQmzdjrwp0hPBzF9u9lxjhO
ZafpAkR2v2lA6DsWu4zHU6rg4sSl4RqhdFP1kurDpnRoGE4wCmXutWGXvF4vGu5a
05VmrVwWMJt/+AGtLbwBfqUb3FJaD9GLjjqBXI2fqb1NjcVkM3vUvTe3oPEKeiCx
ev2OChDOh1tOP4Pay2+/9kk3iresjoFb7d99D8kegtbs47flnnNsJyQDGlZAlipl
G2H/cZJvaJzxeb8Ev5yPulDS5j+PuBO254zmcQuevySicK434fvcwMA0qU28BuHq
YZFiIH2ACff1LwaUh7HcsOv/sGlgxFobclDhtsLhO1xF+bIARkvd9+1gUJpJqeWo
LMASei73QKX8elwJH2ku1MaVF2PmKAIbQL9jyp7+yoJuwSbR9wJ2N50HJsvEgLnQ
JDJEf4b/O/9HZh+kZb2MqNCvhLvLWszdoQE50bFMz2g+ob3NO68coqJtmIQcIHe5
QOfTdHdooyQXv0Ex6mvPvd/YtE8C2A46BscQ7UmezViWOY2LYFL1ej+z7Bo0P+er
xLtNA0pHLfn9OBd3Yrg5iC1S6BQQqViPSL02jVdsyWohY3S/aqrvpYT87ITI4NsX
xcqIjRUwYjn6kasydG/1562gJdxDXkJ0Ptm/8U7jBHHOkuZjeYlSseyVV712w90W
Dd90/mw5GNyEGLQNAXzYOBuHVs5flvxru9OpGxrAb7KCae4SIYPgMu3OrM7DDHeJ
FLF9/Fe3RT+5lYB/1+HtDvCJhE0y4m2iY9omO6mVL10GmYbSNh68MqXPtB4IuAkO
V9GcpmNO1ymlJt1Et2PmZWrtat5dSpiN3wKlHnnP5JzQR61z/z996YUWFFZZIDb9
KrgEt0KkjSB2kxfooYDX5ly3COyzJarKTfbQrpc5S3miruBQQfRWRkMd/5/0ZvvG
k9F2F1dKxc4zMlQiwUGLj6WL8V/HmphVs+OVp5f4bVvhpXPni625ZjCDLKfZl+XL
SyTIa9d6hJ/i6JFLB8BR4ySVAzLl2I6TP3uQqWvf2I1Q734T75RTCfMSG23vJPk0
7l7AtPHumdIqYoqJKfKA4tg/voDfj1bEwoU+de6HaT0XpPCyeajeFVY4iCepKkkB
qfp0p9pdis0FFIdm3UyzCX3/9oh/dRVNyjozirTIx4+TXObh3pOr8lSdiqVUU6+X
AIcd9XIp8XzxlU0gDNgHSPfaTsxUgYqfZxpzwFzuusSria6doWT9fV+a3t7xv/dv
QiohIPkdRbjANmITPuoehRRenU34dawlC5/OnygunaPtl/4eLmnxniq0s/fpmDuw
s/3DNDRuSCYdHwkIff5vJOaZLEhc9yyRJuUh5L3QPdLYp/XhlHhsmBdqB6uuh+v4
5CVWz6ip0pl7Mru+8t1m68YJycrcBRvxceHOAv0YeV8LEfPMiGdVlAsy2I9SOVuw
6kmfi8J1GrFizyujYBDE9ahSq8c7zPVpiqOQ8EtGnU4vt85TCHvU40XuQEsPG4Ap
mFZpR7GntpRjdGNXT99J9tdk+a7or6pDo44ByQKdjGBC3RR6m4Q0QkHLOSs4qdMH
MtlI4XrYiMvR4A2SMWNoscQnYXtAAsuoYV9iz7UngPkA6pOPTK47YblvkDitTdaJ
uAJ5oD2AerApXIpzVv9SshZE6rQZt2h3ygLJQJBqcRcZaWV5ESSouSzpXJkqm88u
tk1zGDnjfDjciykKSqZmDIrWAzGQUvp2jNb6lJYzzBpu1NB1Kxy1JhStbaj9MyzK
LNTn/Qb8hnmUn4/5+ABLVyfwnI2ApxEcT3yxqVksqK76ktU/tEaH8YzV1vQQwoBG
9Nsh2MXiKXu04kBV4xcnXPYnKAQqMdQngCNj46JOsDvld1ujqxu2/KvSzcgf2amF
lnRIZLytxdErvrx1Hvd46vjS8iNl6eEQfdez85+r3N7TuUp2TE2I5+N/D1IuYbfO
zYiLSnsmH589Bo6rNJTD2fxeKjwlO+3ndG7l6x3HS2SUQBIG/b1TYxQ2eK63Vxo2
oZaHj1GOnblqlA/+FIPzXv4ntu4kBZmVmCSskjdrDLQyPEIxeDFqNfVMS/Sx6+qJ
ZmwDBD1NyiWLHHy/EqGbYE/bow5W7i4KxlRNqKWA81ICZvtrpjfnSHriodoLVBux
WiDe/84x0ZJ3hSjGDEZ4Qx7XrpmbrRY6YMWxN3Fn7t/jfC3KJMJKXP0PCLXAm4NK
XvhWkLbpYeHDyrlSR3yH29UQTKdofyhrWOJ1yP+W0vG+wLaneAkRT3nTp9RqkrVf
go28pPOSeoe4+zGwZW8rEkfWTvzOyxaAyRgcJ2KY61MeqdsVhxhnjRVNBT5ILLCe
Y8Z2zEW68b1imLer3RRjp3rMmw1T8zcPLYR3HsHPydcmh0YB+fN9kz0tjCZa9Yur
6m6LAn2PcTq1Mk5muJ6JFWFmvEgsRpgkRievki+4A9kGRwYNtQTGZrbcd19+jMda
t7ORxkmXMrQA5KqsMr5ytxAzqLhzM/Nu5bgzhbK6Sw4fQfyjNHlQpH7kmXiEUGJB
/+vAMiH1ecy4nHTEJapn0IzSDhslO7cjCQpRg+2RYrBWRmaLMgSV5ryYK9X+IJ+4
4koWZ/clNrnV1Lqu+Hxz2LDz9iku3jHR4RkcB9Bh1WBguDqRXWD5XOtiItGXxmHJ
qgBwbCwVSYgpvq0yDNtgeld5diN5mRxjV7ga2QPRI2kBQ8nKPx7MFJQnRNubhOhs
G2nD/7E6jpd1gRyuzYSmFqMUwsk0iC0I348IhSpNGiA0dauq8elCLBRexZ+ej/Mx
+fkjA4LE+az8DrCGVjpZGyvhBrhAUPAq2RvtWe9qPBb8nQjnY1WHfhzVxqp8eCXE
jTCIi7G5DfzGQiZGCFwZkpNnQwxlIiyK0K+aHh/Alzo86kaNQxq8h2oLctmIRDj+
B0/cNIldgKo6sXg0ut44GoHpBOqbIXibT9qE0YviL9Tgm4DNU/8bJbuG1pGtO65n
UcON18RRtkE+LHs1Yy6B8Vrq4AGLwDuxQR0FQTO9hheKByviwRfIsHXms7RMqNid
NjyVdr+99hh6N2fOm5BzsFJAhvESPsGvGSI/BTAEkSAjcemnv+iMNn8O4I2lJ46Z
oIDs83pnZnreji++KdQ/NUinoxFHYpzebMoSRJjXRCXSKUCreil3M1JSeBtqeccO
2rA5ubzA80XWjU47I477Xw7P8KKfZf+lc9LsBycJLdid3ov9vRjxYvjxci+l+Fsb
FZ2VKdPXj6bdS7X/GP3wQvzhWoLzgTUE2jEGnpfCWAkRrYr14WGNvg7uuMrTBl2c
J6hoyWC38kgr2jG719DnmZ6ZzGEtBy+vpK1sTt9dPh+R5ytuFkwkbZq8cL4Z5gdN
+fLeMGNKQo/UMCiC9xJop/U2QqGB8cVzdtak3uOUDs2WfVAZZLGp8OmiF7EFcFFO
1ZburYkqzkKsKRMYQyxG8hN6kgYrcz/HQKl5eFIZ4WQc7y+urbmDX2jsI6Uv9cu4
0E+7Zv0HCRZcs7XJ6X7A7j1coVGsMJ9A3tOICssxoyIeFckXzAhzkB3H3VFLqx/L
r0w0pnSD+kMs7i0bIn+Z8C+oRB2k5m2vplnkjpBhSYtIV9n0B8lnyVl596620X4N
gxzXYK4RI30tBqqKpnJ4wG1wfRrW77v/k5XRtBs4+gCTgG6a9IXNL93PUzjwt6cN
uNyxyz5vJutg4HmwR7JoPRDXRzOPuQv4dde8RVwhUNKJk7gvB/iW1egMKCdzXkE2
cOch/GrHdMlLi5Ua7WuUT5LN/vREhq+k3wQOeenuQp7VHN8Wi/jREQo/1py7O+Mo
omojHtX1JV/RqJCp3jrRJoqzjJwna8IMOs6pIudDCYlilZ58ibtDyisKVo9UPr+z
b/s9FKwSC9LHVLyb4QA2TU0pmRVFg3wzfxs4mL5VAvetJ3N91iJR3z1FAmroE9Y5
iVGhRiqGR9I9Z+RQzLReoVG+EcWjlof/mi3Kge0Zg7i60MjVq9L4aiEGauziC5g9
/boTJ4fTzwuAFl9nZpJaSyOm0QF0UzAtd6hrSvAwgLUwSOwaZO9WntF44iOc9tu5
FgGMU7UjwZh8HcLGQfhFD+bF4iDNt9aIesSwhIzPoNDaZ/dirkBnWqmMXizk3veb
DBMz3XS4576xky9x0IRFokjNpaRVmOg0DIhWPn1fvZydeoGZFglwLxRygw/C9j9N
a3jViqR56aTnHdCrX4Y6NJ2dU0PNv1+gz+I3z5AROP3AOCG5rZH9z+FrO42UAEOm
Di1U8l5RhgWDxaIWFOW2LR+vdSfFlyW5PJlYWTpgW3DUDrJ4sNBg8WIbT7A99AZh
DviqJZ8sUHGRvkbUabzx5sPxYVE9FvAuLXvNrHkT93fSa2hzWm6uWKUw1Gr9ect7
8VmjcGnfYpMfrzMVyzE7Av4qwxRUyTDfqEsra/JEW7JkfYnamapF4M9TpEW1o//E
L0kkj35fAiO5rbDec1WS7B+qtPOUtFZeEhv3ydKhqz01LHaDoznVD3azkBtiq26W
RQkwAnJShjAK22qTjdEHST8Tks8i3pnROuO4Ybn7h7mtzGNMkkmpnAEiLLB77/F4
1CVTWjEV0OnDF7jlPh8P64pMjNL66rOpIBhLMpEhezrGnHh+kA2u7YmSb1mAHzhu
zeYb3Y+e+7n3AUGV30ZHAU6RQTLhtIXrSg62UTqSd25hV5Z5IePdQZjtrkhxy+j1
jReXtjQ4fBolXUHamqwsWIOEzaFzLn7Q/LQISBDlB+JWVnXB1iDFAvKW3h+9iA5D
e3RhRL3Tco2iktj8Ybs88xthEg57N5Y0SaRSKW49SPOOe4eVxaX0hNWUZBk5glbt
oKQ3ZyJ/447QrwNiZmBJmf78zfrivYTEUJJpi5pr6rrBoRBiv9rp1Rdraw8tgEDJ
Amh/BtUVZJJ7x7OWukK0rrVRbMqUnjIk96wI1pStyF6g2IawoAPjX29PFFk3UiJ1
TL2LjcoI+/b3HE4btyAfg2A9Wgm7vBofiStcPaoJl5IzLulQ2MCCFcdPVi2K/YNb
fVKHDUpiIiZMXdWdHTAobN04knX0kyRkTVfrl35KsYB4E7DOjcumzlvXeXYauk3E
3FmoqEBoAuLS1/O4zunvzyBDr2UR/gHVIRXAnc+iY6kouy3PuG3mx2N8OcocUvLp
/bpZZu3UhDlorLItgBzw3JhDeydqfBh+YKVxIMJcYDLJTBF+gPjB3kzCTSYXv8iV
KS+AxGdr67n3v945YwVoWhqZDEHdDOCkUuVebHfe0XWXOg7LXxTiD+exKoEmPD9F
5N2sLiuaifGW0kJxqz85YKrQFodFUlvxI+g0V+uxKr/Rr7NGaVeyECVXBZ1qBUFw
di2B12gtwkWaGJn557aaoQ6pDuB2wUMVgYyMjEVvfIWQe2Z6hcqZ3fqeu7iKcVUs
Lnwfmx3it/ywvAoRgmzDfTUno2QJGeCw5LxkvI7zY81oD8tg1nhn8tg07YScBjHR
tnWOTl0oX3BOcHooq3UmQz6G/2eJKAZwg4EBiykfv1ueFO4mGbFp6pe0cjTr4fzb
+G1reXFUM02J3qi+eBhbVn9Si7FR+shDRo+PJyg4HyDFkHmBBtDL7KOxhjaWdrKY
iYMH3xiJ2f5VmJkJfe35zbEUz6Z8s4mMmFbMUCfvR8vXj1IC+Pi5orsbgXHffVsX
CiQz8+thQrBu6bEWO3+khMKcXsOKBXHzk3aVLKYpVIpEVrmmUEdjXG/nQ/drAuoo
iswX9lF0aLmU/JvCRdAtDfr2VhSaHuCjoXeVxpsTxkmWVU4u+lU23gh5HAJ9HPpR
ixVmh3TU0DKh8jqESLVSU6IlKRlFAuutkVCsOP4+b5HeVI6b4RDmMrnHSDR0m6Lo
VlZWJLmnEliE6AOaAa7ad3GswQBj6HBp8br2u5mHDI6l3BxaBxg7zAEZu0Qnlnbl
2aGcrjbmQpsW4Poj9GzvXsBdkUIk+YE4fBzvfxglY3Ci6D1ZkdkAHn9wDQ9/62CG
YWT8aZmE+01RGNPL4Uj9hNQBLL5n9U6q6cfQ+c9X2EBexdYVSW81lXptuMXIjchg
GXsw5YVUz09GL0XaIkabbNA/2nTwEbNKxJ+uqhQm+ZRypNj95okfhFFG/lUs7fgN
6Ud93bqUrcyXlw7H91umh/hXFkV5xR4lU/mMFoHf7loiMOS8QvmIUR/UQDQV0Mck
OX1vAyBH2VRXjqYxYxrTS0LX5eFUGAd/RgUygTWwSJkgD8U7ppDi5d+ObLXSb4MR
PgY4hcMAHnA9cxaJ5xYdV/GCghtydoQDVmQQmqHYQrlfNLRVjhwVMXXhqJ7nxSqm
bQh5x/kibV+Xwap1HJCbKS3VdtRnmW+hNHvCGPCM9Ke2icsOUaN4yS1lx6NvyHXx
O4YM+NiUfLLE20p0h7cPi7V9FuXYD6oa3SYLQoDteyPiZpS7mk8lE5xLYEuvC3/r
9Wl0NJ4pEPsJdKbEABQQWF1YrHPQsHt3UJzvAb9YhT3NN/HXZVG0XfBAIMNnAbh8
vMAWsPemDGdd1jcoFime65pX65xm/pSmQBFy0wyJL/hIAQT40GchdugnzbR/Jib8
wmWzCNdOIr4wsh/kYuA+KVfeoTD9l9Wx0ftmLt31GnkniGElTR3tkpifOvX+rdMT
KSjTf7qI3TJniKD9DosWx+eK7dFQVtx/hk/IYtpeBGbwsgd0Emixmgrl/KtV8vaa
Tfby2XdDSUZX1+AVi5f+XaCUUZSTUhpc7ZZ+kfrT3hBEBPmX8fSCC83jUt7yo223
Mi3d4C9o5yiV5Ivc+bZmxbsiY0p3N+ObkvQQ7xwk1M6ncR/rIkVZ373t+jpqkrkg
kSJvCnImokHmALhETRGKGw1pUpCkpCl77H2p2TLHOGbrGOLxktSXqOqbxDXIjXMq
niUXQxCheqrfFB+ZY5YgP6lrWliu5JlG0KxwjmNPF3iyZbDn5ewXhwvsLxyq86wG
QPzmYK8HcTNKREAUFPvkx0d8WzAbGUnck2lW/wQexnUwhrAByZoazydIK9BkPDtR
En2StODflcGiKfseVPaLEwD15cr8aPmdVgLAdfKGy1sLSvp8YEN5OqLn0bGTqOMj
+79d8r0SxLAr3LBcfCq0mMg+2VpC/eTAWCL5gbNVWVS/DGg7JCtnr8vKWg6kis0D
OFlkChbaATSYuQLCP8SAFGXarxz8YQvYXcRy1Ofna5dS7xb6/y4UA9pd56mSWn+S
b5egbwd9Bq4P0xKb/dQTGI1v8M0PbjOu4f+Nv76MxoMZDHTu9IR23x11lAfnnz5x
FDACNUTxBkQqLQTDdz9LErtVOU65pUes6k0h9ozjvUrXgT0HzsIrseycAHqFiyUR
ryNq/Fi4JqIK+XYkm7OYneazuJ+SlttIp32d3UKvPy7msKv1o/Q/2FF23rfmRceL
wAmle6LmFqaU3qF8UahiO7S+icl9/wRYCOrmn/euvHm4WGxBaQPHxJvpyFE1+C3H
hg0ZkXan0DICfBwcax+D09M8coppAlt/kkkJEi7PHFJ1kXexGhnRJhsNanXr79q3
RnMaBxRfwjBg6adjwXeLl9yy58Ae5i+hB63SOv3i/XvHaZwm1+d3dDO8szGDI6ay
f02Yg82VYvOLIBPjpFZ5bwdbXm5nDkBbzEtWC2tfJtWkW/QjBYYS6I1X43/BQnf8
SW9vu8imjjRThJO/6hWdWWID+XdYBkGDGGcchdFa1toi5AlgVZRqE7b3xjAxaEOf
Px3D7J+z5clben7zcW9l82EHsD730HFuBLMCHOCbbNJQ/w7PmL3Bawq6MGb6U17c
0FJMcSHpOQmvBENDLgU5oqPgWF5Vjr0skycFLufKLJA5+gcA/8tDi/cI5/xSRA5K
rjk6p7RXSiGKAMm1OupgCvFcNtM6L7+o3kWZuxNNXUlPTNTkuz7tHUqPGdbgUIum
iiBGU3Hg0YdM2pE0Pi1HqvNe0NDCjlH1EFPQS/6xZgc3B5ovN0SF8usJ0b2J7xiM
vEV377+eiqtpLperqQOw5z4Mt7AFXVDIUZCgRzz6jeyuA4kexcnR5gVf2CmjAYAm
SIqurxRlrcEXF+7t/0p4Ys4cWY2MjSY7N9d81EvqAyEoxNRN9MJejMDjp6RR9h5H
9FWmj+Yzq0qfMSj5FGz2amBTc9snxzwX1T09Wrw3Q02xS1xBTI1mxZWjjiP8VATQ
3an+07/ahMQ/7YIJnHtAbeal9mpod6LPIJ/WCYeLYDTL1T8A5FiKAifx2QCVYAqv
WG0OACtql5Lb7y7cXiSRovEDvnw4XpR6lQMtNeNwn5w8M1sdDOCG9cDv92azdXdO
eenm+0oj78yyNaoDvJ0+xHdC5PpJ0Soih/0QsVG26BQrno5E4nevmEvcVfbEbVkc
s4l3YOlkOgutS3Upm/QKzNm3dVygnlGAAKdpQgWl7c3OF999b37uUJ59NaidQl67
vNN8Kr2GJC2UEdyV82VWBMzN31w/nheLNSdelW/NylJ0BSwTggXYLDUXzD5lw0nH
9aWb9G+gcIrpnwTZvNeecApiLy5F8br4JuclK4Xl4r6WiLuGAkpI31vQclMJkB80
uuEeyQj/8khBpcIEvAquF9eBsQXT93ZAVrQmF8citDctpAXFzlFfpRci3alst1gd
0GVnab8YSfBjyALo9xflyRlFfcMYAtv2/qGUdH2HZphxUR2PijPGYqvMqik3tqw1
mNmeQtfx9cdVrSj6luGKv4XQZoE/EqWDHOUPn5+xHJ5TfGlzm/fIczxfynD3j0B9
mDwq/CEOZfmH47Z0p84uQngXT4BUYRSPbU3ygrO+qKv5MzuZv4C1+itERoYzbYI1
4C2afCShKl7Lrt6lYtG3j9XNUoyBzPD8A0sm+G/lWvtYYieMb0A6y1UbHzMAkx/4
WoEVgIeLAvDctcPwtTYXQPPeLcCJGQoED1QkKqgvye5141Ze4UJb9TrB/SJ0ztPw
8oW0j5sDYh3xryt1sZngpcaPq/aSQKHM/ku0A66jWeOu6oRQ/SYv58DnQKzIQY98
DsbRfnwOmI9ZuPnhb/RImSTVha/rCvWVwIm98TCPsZc6TyS0dDpIqG9zDanIf8cQ
HPq8W0WthNSHkwYSQXiQavGnzJk3CVC0IieMjMR7JQaPKimkly0m10hF9uMiI8Zj
6fOcyEvdrsPf4P93Mk5VS1wmbFTcy+nBn4NWn5qxwOduzG7LV8+1E6rxZ2lxAU0e
UAmgzUPPSIJQToE5/3wchMU3Ig36N0UF0F0NJ2c5XT+WqYFoMY1bTPku36+4b26j
lS1QCAvJiuVoF6ix7ilA9TpCbKSq6JYXrGCX4tVuNwlxU1ZdeaWW5PAj456l8ZlT
MkLuEoP5T++J0ihO1txlR3pOxf8dxODpNlR9ftqFyPeWARUegV/6YtCx3psfuHU2
PUD6iZSUguGKskMbOttSppXNnHE8+UOgZm/ryV7+igTTie59hIzXzYW1LDH2LNiI
qGgNA5PntoI7TSXV6OolroOCpTL/3ec/T2kHYvSmEKLOUElB8dM9cFOP9ghQjFuc
mLUBEHk97yd5aQqv/k2iLz8tSdfbV5J0GhIb+HX5HVDh3HkHE4gh13U2dzau16K6
gd324s+55fteRyWgmrQFOSxkWJ1HNpEB4HJrdIDP/FmjlC58bcfwSzyzxUCQ09ir
MkVM8KRGTx4NH1Ei9a7yZKWEvOnhUqgvtvdfjzz0xOxTTSO/dQH4ZvWcf9fRy1BK
SawMif1u2SfysGqRR55KDWhWPleR3pULglLIvxx4rUZdDdtSw7mZGbZ309ZsOhX1
SON0MdxMHGp8XfpHiG/8iYWfKQtoUA8kWdBBX0YKWJ8daJQBbYC4GJK7DoUiKjYB
J5PtElTcd56MwqhzBzjbW7m0/sCmUi7FBtXvN62Nu4y5lGI1yGH/DQ+LiX5vqCwx
bhGxE0JXWfacNv8sh6+WPv8Fe8oKgbEC2zywgarO7xNw0wi9d3WDl9BuYVHsmjk3
4OWcZbGT/VtORSmhL0wtWYoDkTqeGvS8c0IbOSoSR+R/o+z1cpsXtUSokzbwwAyg
4qC88hY+nw6pDTGN273elsmhvKemgle0Kwu1xGLHaSaHaYSzisT2Ge5vFP9GJlnU
0faKwinsPkoOGYZ+XWifzzIkLc5EzwGNxOzDpYzv2sAHj4O6RI/64VRiwS9FyyZM
hqyPleVlHO0nLaL+SYBkuwk1DT6ndw51f1qFlDPF155CqLD9Lrc2jNYc/pg9b8yL
yn0WEdRE8B0UrUhl6Hjv+tVPfSrUCmnmLf8huhA3Z71pRBESvFsX6e2WlEUxLXPz
zG6mf5vWZuJyYoHVF+s0K2vXfVAHseluz4hlYu0x3y8VOWqzTr/oLmF8Omj4qxL8
6eGvNyO5HcFOpU6TCFKx/D+oxN18gK9ajgpIgJ/ChKL97bOdvAMEiEb/iNvAsWiQ
V8/pdcGuXepSFxNEA6kSKv2YbsAcjY4PpF+F3vK0nZ142vi/mN/TaMXLhcmbIAc9
gZTlwyJNBJNeHhfRPgBR+nWUd5OSzGLMkSlvJ1Q9K4d5lcfs27lZBSmguOZKwiq/
VzobOlLIngfJ/z7zuraULhuvm6pepUIIW3ViDJ5b2tCjI+ryPF495qyW2eogovj/
e0Z/4bW9wicS1pg9AZLbB0ggOLnQ99TlKsFbqla/15ejZ4biCr1j+AbI3Y8oQq98
2SdxUCY1BSaaDwBfyFZe0gVR8OYsoDeJtuM1hodTc03o1kcJj/TpyjRBKmtJPWHN
tsHFt3figFmUPO/ugh7Lt2drFxy5lN+0RgPWLCbS51l9lDeuzOjg4LrK5T95IJpw
8ZRflMR3ucIJdT9B2l4jh7sWMmN/Y/tAYORVqWp5Hzd3eDYkStBBt6NOs73HSwat
kEcWp6932p3713+znjDlFFo00CAmOhMyOo0+9FJKjZdM2k78K2FMas9bO+9hx8a2
77jLRF6105dnIj4GAOUaoDQQQaDkZDLkvf941d12f1pwZqP1mPISlSnTxkiWfbiU
OzJOb6B+FWvW6Ix5YsMZZREv8icaodAr5RHJCKFiJOK45ut1Y0ztXAvPwYHxn4Qy
igxdcEMAza6FDYkAFshH0K0YwM/2EM9SJNfBoJPQwC9X1EQX7jW4Pm/oDaOc8uHg
/23mMORueLbkADbXdS73GkJDw6E+awwzMrttkW0O4RP8DdWA3AmIYetGJDxRI//A
WoH5YgPsiRSLYPOfJT/h+ICQRFqRDUL1QBbEFpnQNa5R7t+biujP/bHY14ju45zS
Fg5FYOu4JU16rTWw429kGGnWwpvXgcVOll/UwrEt15LVo7jnkAiFgU9Hu5qnKnn6
DDFJVkxcjJMEXhMG2gTFSj5i04LFwSjGQ/zI4wowMIT09wCHMJz2vuD2WGNeUCfy
GT4RTFhpTne5Tx34K7n6pZ9+hhlwPhoT/5pPhJayTFM4dORvapqtet5MCAdEO/4/
mWTe5YDtGAMbHKXvZ+rqh17+qhHJC1jrkqnYDsfAI94mHBmtlF/QPsi0A52n9k0s
9bjLX+OAIPOUsZAi61tbcSfmI5M5uLnWXA4J2quOY5vI50k19ThprN47BoMJ059i
4Xh0gqp5JAC3IOdn8d07pJvr92d1YLrayW2OXj8fUAfKVsPn83G3sQXBefdfO9pR
xZ6YIrYLFdJ9AsnKeXZScylyftlOjQFt2wKPglafgZfX9/1utl4QX9k2x26gsDdf
MV/QrGV/sx2GWCBJr9547cuPsgihsljDBFzt/LcPC/l7FpvSoUOLIfJuq8LEd7NQ
DGfxQ01TJDEZ5c+cWD/KsPMKJ5ci2AitkSnxpbsh2ZtCu4vVBB4m/7KEhiN1PuDo
1Kli9CV/5CAZrc5nbXAsOg+0dMMMrmoYeXPuQIXJjgZ/p+7VbqkEZj4I4cB2zAUm
4rfFFJ7AaGCLDMR/2iZzIHN54vhf1lXEP/9lskxix4sf6/uv+zBKZLhAs6UlBcqq
q707n2JvtmraI3gnzrSWh/NceEoQtW0bi8BfPv/ojs96PfR2UWzICfzNmNBpA05u
OeSRasla5psBaFcx8dChjmJNu0kXzytPMZfwyE2zOdnQVnaaOvf6sXMlIEjdcAiT
CEjycFwt8VxdPXLItsC/YbBmzM7mw1U10RBNDaml/3FEHXI8XOrGYtKhamET8aY1
J2bVlUkAVrYQwSKa20VaUUpf4GFuEQi6lV6A7y3UkT8ChiRPLDwbBZdLiSFth+PU
byyG6KN6LI5hN63eYzH5B1EkjNFoC2gWIZvJG+igzF/R7jnUFM7eX4nG66Qjj0T6
AYEdX1PFHiXzAy2WAM4AQNpLyS550HIwfHtusVB6hTuu6mH22biLCJoe91ldNzJw
m9uJ+6uKdCQlWfidJHssMVEhqJDicdtQgqpI2PMlfXFXk9Yd78euKTYYa1CvsW5N
8yWuQ/9wvlguD7aLh8QPDJmbd/pgFkgY7B1fFK7YT+SGCKGajQIiDiyE6ZphqQPG
tfZIgDfpeVZABWpK+GfKFbv/+d8217iybhBPcfklddP8msxDKrS38GimzrXPEL1u
WlXXCHJb4oUG+YpxRar1wum7qr3di6bxG6ghpBsdBbxf5809XNCO5SO7NwiB9VOx
bKkfQpr9pIsi8FF+HlwvUq8XcuuPBvf33aKxcSFfNo6bFdd4qybLzXN1UGj3z8/W
zpwd7bUJw5cRT39txT9FmMGxQ2fs8QrmFBaiMxVeZutQkHDdGudFnTzNKy8YqYm+
tQTULfh9lXpS+fM7HR1leD+B0hC1fhTOYTwzJyGGNMDko7AskCh9I4RKMJbV4/gG
RgHFwY5FolBYdOcezCuhqhPx1mgWA8ckVERMjPFff3F9OYd4DtCFD0Ghy7Rl47FC
0DPqBmpkiP2ficDjQ3e+dohDsyqT91O0R2IXbvRi35yq4A5iGX/XIh9sxuKsCPls
eqZWn3/6JbuXDpm/KsZ+GhGYmcNWahaRFlNiLT1hI0miggtmPg0oZEHumKrQM4Er
5qLB4PDFXdJYRAO9U1A8hr1/MtKGi3L1vUngBQISV810P0Ea/378xelVoBtwWe0z
7p/rD0Kg6y7sidT/yiwmTUsJQjxn/TujLZVAJK1aMZhwCf0102TkF3n7kRlPAqcP
MkVJQ2JHOI9w2euhyWb5KJto74sAoQonsDBiHJgW4MioHJW1rGgTpSfIsA7eEOxr
bmdPEI8jkDfZtKFCxjWq0C/aAPjjechIIwckjwS9Tu3O0Wa/5DGDRqjd2BgHMxno
wcwUTbq2c7c4cZGH7km2v0ra2iuFu7hYUSpbBHM5IvW0wn1/lTBqpT0DrHwbO/4N
wGHho1UdaNj1IbaXzibOaYQPE7CuJt2742IEKId5GYDYemJdJ3eKhCS8NCasTPiY
0FnW2kHoDb3PXfCgnU4I7TRrvljeHEZ0+6EygbttTcQck+65bfHk/2mcwm6UehAp
APhzzOQkokES+5MoOTprsebt4PQuNVrHRvC5B7HDpofEX07NroeHi37DiwTUQRTf
DSGuLpIeTHg1dp2+n6eIkKW2WHR2zGbX/2z6SL18p+W21S8oX6l44sh4flRfZqw+
MfbkVRhvpjVPRRvxUxEqtjLU2olqd0YFnGHBNafPo5rT10r5z2GP0aJAqf6x48fm
8htlFGcH9PzP7poMjaefkvr6xwllo3rMbaS0siX/061kOdqomQCgM1lYsJ6O5Biz
VigseSYMDPZLS/wzZ8l4t87FNRWZbrCgyLyDiOOTkYTWNc0BRxYu4bkSWZUqHU9m
eEh88TwBQst6bsXb8itJWcRWaq0ucUME48O2x8o6oHYt0XrMtQJlz8TQh6YIbBYm
fsIzYC6afTdxossCHfX06wCnlwR459aLk/1rBF9O/mTSQPz5lYgiOCnWDO63OdHe
+Qy2ZcfsiCLRC5i5DPmcNxlsVOsleCRCblAEsaqMoPIgq08Aq1KmiV+U5DZLuUfm
W73lGso4ukOVRwiA4IUpEVIfnQA7/inTnVXJwF0KGqlY2HgO3xQcq/0Fc/MEhApE
yy0S7+DsRZBJLNEOvG4IKUkDNkCsLUezhuLWwg78xu2W1DfFS+5wSXzT32Xq9841
pZ27uq4SmCiIA1CLnwgTnthNsAo4/vhmlKJjWYPGO+jLOik9iftfJI0ezQImZa5R
zl7kAHP4R4v5xME7PAodBa2VTesWMMYgwooH5M2eqWlsH1DApY3ejyDeZ60NgFGP
QEQ2O8PlAeqS3U55eeiRDUlb0L4AJe1KrSwfFXFxoRNyzqQ6ehSectDwJqJ4Qx9O
Rjlq8fxj7zC8fg55onIqENMmG2NWihBq7mkAOdRBiNl/4NA/FnnY8gSaXf3agsr2
qbIo/3k+GfccyNKgkNUymnDXGCOPJhWkBjSOUxvjSDVR6KZ3sRIPcA4/mYqRXiWW
YLDfIdeHp2sv6gPHUVt4ctQ1kCLwfPBvcotrtCi3ceNRKyJbViy8e+qcRjnF3BLB
h0BSV0zmtpKeFKJbtGztnMUfWRIEqZAPiwA36IQmhG/2jAhIW1VXz2bj7OcoVF7P
/3VgMX9B4cPeDZyHBtWHpGm4sqQTRHzcku1x/l5DzWER9za57i8SGnwt3zw/TKfy
8Wki7N7uiDACzX5lfKw8S66Gb+aj1tmCENbnm3rvqHxLdu2YDwNAY3i+1yFtu12/
uASK1gjKuAyEVF/E4QjO+EV5vVYxcYZciO4ps5erQTcU2bje8sfe7Kecsj0PxqiJ
zizP1E+jQHQTDITkJ4vXYvPbyfzSzluxRKaip21qTkhk10eMPMNwHU24W2MaWn+L
nuUrG+rkMVhsiiHWL4L7X1juLFZnjtS+tl0nDxRod0dl2aT4QZPECVMMwN1b4wyR
FHkxK6OYfFLXPtp4F5/f6W8kJa/yrrgwn9rbZkvM4oxAGQ4f8rPsqgIkT3h6GrrS
l0um3/F5X9wQcLJdoaHSA3Fv3EkCHmAAjAzhD5+LeV1B77Nk1k6GSmxX9Mfvk20c
7CyOKkoSY6wyW6/bZk3UhrFR1sDKV04zxNZC2Zex80Hy2peqBjb+OIjcNSYNDFGg
PwKKPaEKI+K3rtGQ30y/HNrRy4cOhssMYv5I8AExw5hIUINJsx9DOTKxN/usnRce
x6EbsF40gXPVsUbjGbcO/EzC4t/HRoCMdnQNFLJ/NOpylvJsVmjWmR1uhtmjpSnh
vGQqBBnUofs93Q7dh+8xT5gKCKNb9wEfeN1Uhh2FLkwFIxOQzVwN8FsVKo13aMCN
ka87EPNWaDNvJEcu5Xhukk1Yxxuce1K1bNlGIfB/Bz78KkJUiLAMaema3LgcHNdj
EHPYWsgXAJmh9HYZ2P8Wf6DI/Sjvhmg+PtSqJssT3rU28deY1NP+uj6cN77Rr8TZ
qkTlF1s5/qtC11DHVv6eazPBgXxUuAFTCVngaBZLX5XbhJFIo2E5CqYsyOVlOu4v
p8EzID04YEImWQt1KO0EiBFkofFSAExbgC/3DuVKbKs1sfaekKosOS3D3iz/0sR6
rsl1309gjCETNzxVx2MCUaUpUZXt+zr6IWDEbU7H9hTleqiEtGkr7Yy9IiIug9zB
D+ckNbOcc4lwE6pPu1cMQ9JZcuJV/LKjbR+tWDWyffgHVIMXefk9HkMbkk8JgNJ2
hPUo9gQS9b/pxtXTWY/tOJOyoFEUVaTgr5PcDrZsx7UR5NPoH3BiN6m9LVHefNgl
3c/ZYAZC79o939rYgZWhUgwGKeV8Z4F9OUa5i+jVvX9DnVGPQu6u/bkt08cJX6Dt
QcYhIRTpXrg73m3j66v2ahWUQ1Qc1Rh9YnlgHinYamGRhXYxwi15rlLz9/NfPl5L
HjQESlfqF/uIMVsnSRd2D1sxZVsaPEpbObhc22DMYUaooOT3bnUEOmPdMLOYL3l7
E9qVLj8+KecaEgOtYmsAhUW9zevgM4bT5+9lWjGQeFJrofTo3Y2c44dX1Ctfo5RX
4Gx9BsxpC7Fp1vYGhfiARC+fdahQXmUlC9hEJRnKvU6lCCM1tDs1ci2N5vkf6ubH
L3qlhGOUUSHoVqtIWyTgY4eunBKTPMMydBI25EH5sz9xRPx9dOs0wysqa1ZyLvu2
nLiy9ct/vAoQCkVTJ2DaiTK6+e4xKIB7g0msKdD+//Z3qOeB+TsUFOi2dkjx67MV
5TuIvZ5QLQZlCVxQmZjolL99mDzqzEwGRawqCPfCFrGcsGmWPejh5qD/i4TpQyGs
SyaDOiKAtGVC0t/fQrr1lXon2Ql0XZUn8SLA15UGS2pS+5j6lrpBCzyEgHX1P6PH
MS/vuI2yrp40GsaJHKuXuT8Ef9bcfXfM+F3cd7MaKExKlm62M10OqIY/gdg34X1n
vfa6ytpz1hcUgaYL6C8G5/V1SmwkBb9nZ6N1kFMA90ffyRVBtPpmpmZ/3zkYlTAP
Nw/V6jhaIu+ZLv8bBOBN2Rw80XaP0WL7vS30i/o8PaDuDmV0yaJEpaRZm9GPRl/A
PHhbAz9BnRvN190F/TT8rmc/kJi/hchJ+m9IHe2WrJyFKqXBflQIFiLc5ON2H6Mk
tTvWdYUICdoQEBkJIzJ3yND9G2ph0mEbhtcNEhEW4Iez74B+/gKeyCJvE8sBi2+L
+/kwGfJTHDPc17AUiRtOZx7a2eEfijfQcwBkeTfvLJCU8NP9MElVFO3MMBTDyzwQ
kzrT1k62WvtTlc6Ftxjl1xdK7Q0EuG0CjmBkh+bjgXJg2ufpF+kfW/D3TMgv1sC1
bTMJMvPZEugmMexGiucnMryumCu0ZBPUr8eWqwrz2GPDwX49SiZNpx0RIKo8rf6h
LV+hjr1N6eZOdj8QRlgm5FLG1NBFLm669YORoHodbfJ4/mPhA1668KRGk2Rigdym
oo/6rmjO7FMV6TbyAJ3pdv7fWh1tngkoiQMReo44u50e2PMUgelmSFiVNFCKq5fk
jACn5MO/LO6FbIbF0SEmTA9Xe/jLVFs63xXWsnHs8CZ0rIaVfugHSCjoz6H8Eajz
CqMIDF8aqNWfnwBL8bncFXkOeLzsqmvZzuy8J6zQuLoGUwXdY7eVULC6iyd2Or+J
wWLW2kcFHyoFLGeuquZs/FurTVZXN8QDjWXV3bdHK5U55Cir+AeiWTErijFHnqFz
u7rUvjMQKAA+AnwyJroiUpcHqVWVjr2yuttm2P2qt/O2BZHwMyy0Z/XyWLlbqolp
Wd71ebl7Zwb3ECh9yyao7qJBO2D5zcf5vBjSk+5DCoBkg06SgAE/kuWHWCark3UH
CdJk92YveGacvD0oXGc3MHOi/dZQScHEzW76kmz4URBmochkb5C02gNEL8q3Woes
VDvcO72H9Eoq7DiXMgDZ+Jt1P0eR+EzPGy3/p9bonrjdPOoMhNYuhUdxmDpBzEXu
iG/fAyU8OEC8qqJMpEmo8tFeFIVKCDCWP3nZmEgP78x8WNrUSl9u6v63dSg7X8xG
BZe6GCBpfhLNax09l5Si1fggLbtM4IL0tqd1ilnBinb8Z91LST3//xfGC/3t0mcG
AwC0Rh3qJANrNmGyS5S2xyeRtOvTwnbBMAwn0PcWA4s/viXsnfR+9Ma3dIbqI6Ko
WXTr0haLTKP+FiIMOL/gPK1kq+tEz5HcYM8KgXeG1NebprMhqgHW+4I3d15SgIal
69bRq4Z1O2OyVPfKeSomQSZfU52VRWGovZIfI+9BEy/IcKyPP+x1lSVbFTSrNKuT
3u664TP8dOAlzszArPFUdialC7BeG/5Q8e9hYR1FjCKuBql4TjHFtTJek9g7LdAR
skUzR78iiwHK28wTYVtm5XgbaveF/lZxtPrf0D7/W2YPhKtF8PYhrj+vKn03hFvI
XT7LPCcp9HSvqKUfWR3ecDqMaAYKKn8/FZlaKTf4oNzxg7jbeJFPUEIVJE6W13VO
ve0rOIxzrPKqbvYHxQ1huk/c+IvqgL6TWx57gNoPc5jOiEeWVWWVM3leTHjqbLbK
f7quvE8sWo+ECFAeMCVL7WzdFUSE9DXB6HXGJYE/FvdOUWBQIhoB2ve0TF3AIXi/
qv+UT5K7v+phv1B0miejRD9Pd1mw6RrXl8+Zl32o/hGf0FaqIs6cMotnKUQlMpW/
Ty27RyEVaUh2FIml5aTjC5FmHTjwv4OiGNjd93bvXjMYKScnrxsGYN6Bht3JUam7
OpEchBnCwpUvyMFrcUUaiWjMQSQaFONTvbv5wqlr26Cebwds2j45fY8BbaVOgr4C
BVVCy4QHxb+nJZPBswr6DsU5BTkLy33Md2w1dKnBNimmjH5GLE1zhPHYKtjhcwGu
ng29KuqYpwBuOQmceSsTdlz12nl5TnSN6QW7XRWsrAa8mzP7OcBvC5eRUKBUkW+h
wqZPp+aPAwGxZ5EM27ATnwfa6G+QTUUsFnJPmuVvOKod7Ik5sYsICtRL58HPjsSi
pT4LVIhd0VoqCurCNL5yS6WCz6cmf5iY7v3aXGxeDXdfaJQDXFRNR/m5DhoPsHDm
U6n1QsVEyf/f5i8HCjRM+lE8WcEZ8G3rlguioAbaAJMvuLHnN0ugxn3Rq/hsTScY
cmJ7AEMAFyJdzu9EKzuZXnkTFKOC0t7A2cWnsYjjzM5ffTA5RxovzxxZnzqfnuqE
+k0XNLOEiawXVijqbt1V334Iu1C6oOSzTmkJWV7mbsft3uzawzZcyag7zc25opxB
oHqpkBjW5baQkjBEIlIPfrTNecuHrfQE7yHoPHhuyyV2hznt5U396ycqo8ktPZr+
oHMXqGGMase9WHvtXLnq1ZSQEGV/EbIADZBRXelqJ5c8+JBO0Xn0cMb7MeLxIMHb
ZDKzDnndpx/2fu8kLtJgnQYcWChD8Ru/qKFAlgpVPT6tb3KZu64/UrBNDcHluSL1
vEs47ue2E+jKb6qabKsclFWyOvkq2fHhBsAEue0r+p1n0/jxOb3QRRupDicZRkxy
u1F+eqJJKmpfIfhuaV/NbgpOcyx7Ns+oIjKhHOEz7FTLmC85agX2khMwXO3oosuV
KuYsK0W/zCkAmnzq4cAdhTUDLCIOd+Yr9924EsHUZuTr+VpTt/iMEb0ppWKKTOtx
rZMa2UESIHcmSew4HblYsHXsPsSR+39bfRhSouxmMq0Fi631JHCF50HmZ62oyJAg
cXIsiCjQK/ZW7RfzGC3+6jz80jey0i4fGwZpKDBlTyvDxR8jQFRBfDspfLoUyvyJ
4yf5jhd6hmqHoRItGuLvMb6VxnG3L4wl8PnMyhNJr/wNnr+CV6eF8MeH1yKSONvw
BFhr+r2GCOWBWI3e/ahdEn2PkOqx0sZ7sMcUHxm9U7aX3ZzjIYJfP+jBKFUpFQrb
DZVnWb/KpBrloifE8u/xkvyeEFxiaVYEWP1o8bC0C/qVbigLVKKF5GhI7wh6u8+6
se8JFI1WIHr2BrQ9IJhiYyAQnHOB3QvbVVJpNCNLjLPu7E9z3UWJMaPOY7eS2jzi
dmGxUfc2A0tDHBU5diW9utjcwSZnFL90I7GCbMECSpqT4eDK0QvQcKwIdBEAXxnN
HQQ+HUhbt0jAqeJ3+feNNmbi/931O9fsKSxx496TPauBpRlPhLWkK3kRU+fgVYsM
07W0BhyCWr/yr2T7Z5MKJxYdxfiIJRYxfhF7iWsjfA65udWHLL2vvieXGZ7EnvMg
sBrPRQuKp/mmDbTUyxYMc64BA8o0VIBlw4cg9/UGYsAMlopj9ewc/Hm2YYLH/k9w
9YxtuMLiuxjAY6z7gxuFIUu0YVyvobbCKRLQKF8Uj9A7NxAMedBgnCy0Siy0Jn44
TvBJw6oAVyZchfF1eXjzkbhOlSOuoZ0fRuUzQG65tf/jMu5YFoMuaJ9Z9UUzh20o
5z7p8Qi20jsCRFO1SeMacJjuETvPA5EBuFPEtK5CPJAxfAET18qNgAdpB/iMAoVo
GKk6C+PnhgbHHTrwvTZYZ+S3pgopBGEzAYXrezqoiRZQ9wZDNGXVAQUWukFDrTmB
U193nF5g//TJEmeFWKP0EZ45wUmK85G40c29t2MtE+ZEnPTvaGFp6etSUsFZogAz
kLM/SUssAxyYauufKgSzmBDoo6prGSIxD/c0O5tMTOzcM+TK+uLXVZVM28TFF922
RvPrioJmu19vkBBQxklpNum0vpykueUSf44SGe/KNN0s/d6BwU2ftKQComqcuKWI
3aBFkBy06Gu9CaP2Pzmd+7jkN2u64uYSjP/mOzG4hMbsFLkAexcv3qRbIx+aZ3ql
ZFWSM0RxJn6vh1iHGBsd69Z+lFMsMLyluy8xb2gcUsNPHFEOOuRAu0xXwD8/fVGk
4fwA8TBJVfvQ3fsnzOL0HesjcVDAMZEjFl6RC+LATOcRa+thyYznMIrOrS7YbDoY
9WhsvJFsgLU/73YF4dP3TJXgGIdgyEP8g3itWQ2GeJ97U8ea/0VU6xnq6ojcxshy
QeaYOMqlgd+AEh3ONWXzcS2JpY69Ag6phsBigS2QyQxtF13i0Gko32ThzGgGKN0V
v/eifE8tekh10osUA0pQp1E3ZavNzToIi+0eLxu8HpMGdp2giqU10gmndhYBF76+
VznXwjjZZQ0mj7eKTjRUZMvBXplHfwf31W9KOxu+g+7foptL+z2+wxTsLxq2+iCL
OyQrrUjyT9SABroK7VoxCYqgBq/CkSzna2KKSrskm8GRParYWdv0O+PTKwGnKA40
q6g8UzC1TYjF8rmKHgWmPBBzYkHxXYq292yQmVBOw8zbwlj/nZrw8LsDN75rJqY9
WF2yyg8+SMRhHkzreVHh5OC8BHf7bbgLR7Qmvil8iU9pp3s/Iook8kUWD21A2FMa
wpfZuCHyg7xG5Vx2Qp5eUFG8nCGRbE+d/wjY0RxrsLyc8nkR1rmH1io0iBgZ2kI2
z4vGFiNcf9XWqlCeTc3U/IK/RTTftwBX2bonWA1wRGa35yQ4jFCohS0PDlStBT+G
ndBdsJYQUr+ErdW4EO+Lbu28Ml5oacNkdDgtk4FL46wLoeujLgjfVzd05dmZy2Y4
C/cEUpEoNZogceDwdlB63dqGoMQ1KKVh7/49kAdNxgjlNDa6ZNKgmHNK6o1gUzO2
5CI9RGVslRdt6VXuQE6QT8sKFU61/npqq2zEyDcbcEBOIzaI9jG+lb46i1DDDdvn
5jitH29hrl1XqQdNJy1ORc9ZUzEskrm7xVy37uhWGaOLKfEu/3xJkCHfxUI+iAQU
fqjz+zLvQmYxuaINQWCXqIraGBX9+fIt8U9/msuk3rYCXVEg4Gc5bWx2xplOj095
Xu3t6mThM1UBNC+YqxGneAQLPPeqdiSE5lbu8zcVRtKpjY89LJUFRHNUcshtW/+F
Y9+22nmyGzXldZPs8GJ5d7Jd+9rxL+4/zbLWujxpU/vNk6b36rXb1kddNcOcGc0M
SV56rwQLXb035aoipgrd+VBwZCpzfluv1BB+INOpe/Fmf/pg4oHRgYAedARCNZG2
V2rgQUFy8By9P84FhbFtbkqbZLZsLWM3V6VUx+iT1hUln6AiehXiKxirf7JlyA/1
dYibTzf5S/791houCz1bbH5Mlg1Lj1SUHTXW4ik4KbncuhqC8GL51bG//CWGhChu
tGwlTIgQQ7DvbVQyHoaMLKYtHFy53JFbLANX5i/ptVDxgrwGDgEeB+5b6TGpcBt9
dciyb8kNLpv6gl3HcuNDxQRZSUVW3ZuyXIrKjZ4zc2lou9u5y+iKC5uZUrRee9/W
jsFK6fEGjj4QYL5HYvzsiudyVaxCzaR7IzfgsDfFhlkT89knerY6ZETKyR+EuvRb
86hpnxcc9Pd0eQD0z5egbY0sKklZH3Spm99WwMll4H6+UlLjirkVqSYih/xRMtFK
HYdZ//lTvkZXPwTY51CJs//QmYHy0Yrra19GBxVOtS4L1kuyC6hBodyAfbXh2Wt4
cc0rucPrNGv32zS6MA1mOO9z3by9oia25PYJw/7AsdB6IJPWQMart1fpCwKxW3RJ
hAWboS0gglD+g3767CmCVCL7tMADWlL/B2ZlzmKKXPYtg4l//J9Jn5Iu4cG/AnFL
hD0i2ek7ubd6BFF+7iSGZfgxdFtLppyiWd97mGuMqUMd91KnlRq9WeLk88z0z51G
UzX/jcnoobgibzZ6Dc5OZd72jKXkRsyOY1cpqTSNRkQu7D6CRyWoFyXludPH4gD8
xLc6A+Ef+Sg3KmQXxnVxJC2C9HIJRfcFG0rvx+mMsN/6EsE87/IJcTyn84HwL3XO
Dmb4lmwjXEyW/IClsqhM8kVriuDnkM0qU61skn9C/lGsIzsSeGhDa568ezP4K8BH
H/391Dj9izkUBemy3EfKKiQjPjt+HAIPROK6V7eLbCjZCZCvhGrTyBTPAjq61mV7
4yhOMgLCTRkfwZ9RYzQTk/ISW/F3bTyo8dWulueeZGodp+Em6xlb3Zp7bv5rckKg
+B+fkww+3ZLz9sYydUqghsbl17y23AZJ2Gsl6bOOpGNqbYMG0yh7pUjGvirvwRbr
I7SeIZB91LAK/Hazo3S4l/AePM8Z1zlC4YgSp43awyIOWqbkwTO4K0RgvkHu65H9
J4XVUgqDjsliZb1poBnTUSox6Q7e9e+pn2YI92FlMXJqkSMmHhhLNXaavZqvoqSM
GewbOV9DNVsowhjkgmihjArPh6b45oRUxYbITx9nYMWjf2qhNkkmhR7mFgeu33JI
mIGCncZNmYPzhTE7EnLgrhp4CveLmDUF6yOD6/1VrD3HlNXPtfZ/a0MvURD4TbhM
Mahd12RuWVRyR5RAXl4Rvr0zkOlaSSdEfDEPCVIF4hqP5Ni6s+FaGzN9h4wQ5sAS
pXRbmPJN7H/piQZvgQgZ98QFFs2/ebc1Dc45MopL10GW+Z+MDyYLP/6C+WtiUCdv
pyaVTg4N2PplODG2qrIosmwTROXhkw6AQDGdqJAXpdfQAAipdiRMJW3sETsJ8HBJ
w5EDEUH5yVoOx72A8U1nAYPYbwZotyZcJLD+Jp+mtH+AS94XG65JLI3XtdbJMwQp
otc8v5yL64OmPNA22a1tQ4SLC07zzoHvbMAw6gc9IgkaNQHlz1/zRFP4kDcMsE9F
xN4QpuDouMYbMo0y9YGbOlgJpUiI5pcd4FhtvBKnZTHbsdRYkrnwa01PYH9llK4Y
XAgX3HYlPYJYNORqAXwC9wcQgON4jwX0G2whJEb7PVKrvGdZHfsOLVTHUVuxKANx
3wc3/IkBwmJmzWg6swJwmpifpWCT67zpSi2ioBcSbponSdMP890qv4pJ0eSYOlMb
rdDbqv5R2yuDyx6N/41nEU7b+cBDwxSDe3c9zu2WWV6KiCmwajdwpsCLUGdv0iCv
+x5WG+PbHl3fWnqqYhjOFGu8LO0Em+Vn+3idpmWx7DJBJngor4UYdn5Hn07eXbS6
gwYLTBpzUMuvftTzcGSMQVvdsBEMfyEWKgDEVuVqueWYptAo0Wjj7ddO2xv8kZfp
l9ozkXYcKl49fVeEl2d0g4yZEm3rX2HSv8Pgo65pqUJKAi+MFlDg15uMYUiVDUTf
UY4M4t+IrXyp2tPxdq/5vqA89rIZGNKNoMvigqxI6SvQIGcs9QEF0GjhqoVtnPR9
+AP2Y0EPhCQFSvuKouZp1pmyGbR0qTMwb6ZX4dO7pItwshfcPQX6Z3V+jP4FWOJL
LXOzGWdBZt6w15bPatQ0lB5DGRCtZLDXScG+PK17FvBR5zcVrIp7UTWMBz1hLcHu
hFUGEdjRF6hcubMxBz/nElNDDEX0/BslKulMqeqsG9Gf/iNgnwNmCWsAbyN0E8b4
HkhksW2LMvWc8vh4kheEZ9rbmo1HnqRlH7nwdJuRLG8GrYwlMwN8Idr+tRU0v3ei
pTiKJ0e+X7pixVNVOlMblrSGiT8QHQeTu7TXwKznDj60H1Dh3+CCaqKvif+2YL8m
MdpCH4RCXpSsYCghq2ZX8DvQJ2XQBu9oQXR9Anu8Fl1FBE9hiDijmg/iAe7Lyv//
0ZM4gKdsen8BfGEyZ9eZiMxnJgdfTEojyCmraf/MZRZZRXzv4g/c7+BdrXl93jgQ
jdURMPO4qXQGnZlKnLNxIOGHGKd3HYyPWIV9nD7otVkCdRHpwixy+3vX8cQunmGX
6lLnsUZg/xo3zmAIlud/qjmCPc0zImHQSeyUrPpyDG+Z2p6YChxBf4MEnSdDIc6G
PE6MrwdrbWa2PijA9RyEANf45DgHx7G7Od2VuYWSJVsVuGQgSTpPpFuuDEc5OkFx
Koq0XOOg20TK9IqV+tgFXO8cydOrqpC5u2Tov3v5lrBaLdskalj6dFv1w3T9glU6
rSa/PIbaU6HXX/aSjymUwsgiRHKQRBLMDNBtxaoJHEfFeYw1z1oJsm6vA3YhQPQ3
+Ww239bOG2K9laBuJ+60KWFbGoWrL+zfqO+bsL6QmWzfdme1YWI/nP4tHasYlEFn
iMlZ4k63LiykaVse88tVbPWtrWeTu44ZITKn1cvCyqZKLZ+RUjRiGNPoGST8/n/W
cmHmKVgVjkV2m/SxHCb3DTBLzrrRw3ub2X+j+CvFqcC2gTB28JnleJzqVGvrykYd
ND/oJ6BxAtuKH52vsGWt+9Vj62Izc+racA2PupVPtuaJ0q9OsAw3td8URdEbPqd5
NzKDt6z99PN5cI3LV77pKUzpanTFzP/4Wq1tH+vS9Pj0uD3/AYXEJn5260NVfJCQ
RWmTWN1wHI2eTDhozKySOGW6VAu4wPuKVGhV2xg9Kcit5waqMjukxRczEUAOt3bi
CcGKldcmqxH9x6sVZ3SYqs4zUogyxgWsrqDBQoLKUI+Qt6g7QjZcCox758zrLbhK
5fGibx7f7PJcwaS+3Kv7Dc8KXmbw7UKCg9y9CPI/PyIVb9tHUXvlKrYTBcvv3zeH
XyeWf5poQKno2fKaFsFFvhAOJequJmWWzcAkXZLm6M5laTZhLbW7J3K+/Frsxz1j
zkxELjzrgE0MEW+l3wcJzRF1wogV8uB/B3JEoDZ8Je1JNQ3wmoe1zUy0WFGJ+2lI
1o3nXGlByY7vN+gRZd80UTPBFnAQW1BEy1xDtfcxfcHBBWkN/MfAwqm0gwfkw2Ij
tBH6f7cO5VvaPUA2vPWbL0IpbNQEIBg1OP1eUUo57ETYCAp6FBzgw8lVkyKlXyBq
LlRjoTSwKwiTvbYO9gw/a4m9pBeoBQDMkXWFqSEn+KWT1yOh7ePKA2oV/Yfn5ncP
PP0+2hWqBe1kGycWa0zOrlty2+gSW6PEATqj43d9lPVvIhuXcpx/U1BqOq/bL00V
tzSj/zRvHEPNJlDzMu83s+Vps/izGL6axsPizXrjmsnu2kMFWkFBfBJySTvoVmeU
Ns04+iT/ZuSwGDBp65DiEZLBpTnQ0DkeX1avJGvSWgFQ9kjiucI6CsFBgEefj5BO
swwRT8Yv7qSGcLSwIkVKeUhimqxkn8eUjSpVdh/e2oYnEeHV1n+kdxG03RGUjnd5
F984mSos+1ArhW5DDgKrTRo1/jiombZFKS4XsgECI4rKI7jIpidDkKhS4sxl2TC1
PalIhjomCf4WnSSkH05HeGw2mTy7R5pVF1pR4hePd+u2kx37UHW2mJtxLc4wFV7/
yu9NeWlmykpJaGcMEsH5vDCGPC77MLN8w00EvGO2c1lkUlgmdwLzWBqyW5TzRhp2
HMYtsfMjT1gUyafVSM1y+bD13+XnzuwSeUd7iLIyVMEslcL7WONWsljdViIN3Im1
OaF5I4lVkYXoCnT/bJCDfzGH19JN7GDHx99ua0LZ5pkbTUvjXO7WC9X2cRXGlreQ
m4TZ7MrmLCu4lzicaszsHbrtAiRc4B0B/iWew4K2FrmKl/V/klSuZ9beIziSJg0o
/OxEq5gtItsY4iYcQu/M+KkR63PNkySaSrfuusxfscAat42lVQHfrKkRfhYkS3w9
L0l/i73XSNcf8KvHMcRcjuMxWkj67PfpsFxqL2g4ze8ICT1iypf5LnhIsOZ3JRMA
6d8VCVoKTvf5b5xFiiAT6nT7ATeX6/UIeSQi+FRFtCF7IhrmXV/UWBHsbVyol6xq
Ax9ZbPrXjWk+3NPCnbZVdrpO5YyM15CA55G+M1tActy/Mpbu9RyerIPUzl4qYX9R
gcP8gpfCGFd+QucQeXz3vKnDsmyGNwDTwEw1hAfYGJn1wT1bI8aFKzo67tNIaz9a
WwWzdMtEtnG04IbHBa1jPeRs8zH1S4eTiHOg0zQl4VCztdyHNgqL6Np2I8BWqL4z
mDuizkeRFVdORIlQLqcF9jw6Nmd3Fa5eyKsiVHiumM6cbDhZ4rU87rHrbt0v4i8Q
AEX3TF4Y/ARP9t314dvNcupuFMFjy5+EYOBKYClfIJiK5SsU2P4WvFErIGvUe71m
CtSwcrXqMXZsXeIjNd9yGIUdGXHcN6MwDEmITERORRjrUlEEEpjUWDAR+wIVOxOR
ElI9rv3Oz7LAlXeRT+7KTuML7cbjU4dNKK7/ZUVUGOgQCJqIfb9k7raovfNP8mi3
RCikYRuC/JzdyIeTs3zGU9ImYQGGeUgH9frBMeD+JvoDLXaTb4FXBtvSUeGaKk57
AxmxIBwM0zUGhvJBPAbUnmVfQ01cUMN5ieuBDJ/wzGnNeGNqfOmKYBR1EU6NN/dF
L0gLtMlA89f0VWTf3/h7H1KPYvNNDBANgK8ayDK6HqU3h0/mrTOFn32WyrkRgEBm
FxeGr3+6vcm1biSzhuavet4g3dhgxLvwclhjUPRD9rhp7AJVUoKf57s6oxU9QmTR
x+kqdG02BjXSTi+y0C9E2bYwb61chSiq/y5ZcnFIXMxEphHC0p999aFtmPDJniqM
A1mNhc2bK2dDXtyu4Ui9skttlszUmkFPHmdH71xf+06ZyZEAQ9JmIKWyyzkLE1LU
OHXDB4sdHAF6jnwcW3uLJso7FU/USZ5RFJrwgUAcUI6jeholmxPIDBIVt5k/9P/l
FghsBnrN6CnBh54bYGRS/eD8e96EJqIBKUA2YwT8P8GtjKhQXJLD35B6u5Fql6Pp
enzuAaHNX2yYUluY9dbhJcN1Ic3R7ek1+5FK/PV8xk51rH/4ofpKCPay6eElQO31
3MDVjUdYkZo9wBLKREqWMO/1PjbYAStB6W6e1crzCSWcL6jHQJisVpD3j96yVThW
9G4bGFMumfiGLxrWzQLTSZX9ZYg6ZU/+ps7vGtxb+ljeT4RgCd5vcfO2jmWHM8Ps
/vFtIqQVoS6ubDFRuCjilt/27jmdAjWeTCZWlwmwZar95C8wpVL+IuIS6QyaVxEG
rvmYSAtEph5i7LuI45wTv9kzp499ouqzI35g7eJze5IvjQuypShhrP1LZp78pUOi
+MttTmdX4qNcmK4MgiSOVJpvnkzBkQ8I4H6ECTGF/zQr7/lrFoWzyqToZAL7Y5iP
h8Yr+bmBaRk4R+N3dttaJ1RMIQu0Hva/gV/6KYkmhH8DmMxEGyePqHYt6p3s5W/E
Wgm2V4MgQfYFuYaMagRJwpOCY4kyvCTWS8wKDoUMLb6P7AjVNi1BHpMzF8dFV8sW
9KHN4iR7vFNWPN3tj/yJ/hrGNHBLWqu4Y4YhInF4QIi/wk+2wPhJ8ouvXBI4BhN2
WuXelmUnUhcxhUK00muz1KQM1taQTG6cmbWuQnZ/TYNquxmcGxzExOI1prOOIlI+
mMHDy+jn/W5sacytTMlJ9lV8qJqXnu7zDsEuRSI7dSR1LOkqNQlMK0WruLhmuCML
4aInLcmhyNzg8GyNjrjl83Q+Lyxw0B7RARBNuChJEGT/+JUz5zN07C76ZR/UTC5V
HTmTRL5UelVp74lXwTNeJd22OGQ/TAhAVupkhkKPitBlzSyCUp1GWOeCSmyW2WQC
gy6f/+iwXCmiVh6gKYGDLePuIIunNskmr9HRZ7W/FtZ5FLmMQaujb8CQ52Mk4dNf
zVyJur2Hqw6lcmP1S8fFtjMVdcIwTQQe8Vi3W599csc55/lo+FHpru9kxQvP342m
sdYMQUwLdybJOVzu7eUItA0VZgeYv9duJlw8/cZwj73QXe3CN2xL0pfpEhexdf8A
LeJuag0zXa8VaLGp1NH5MTZYiY5JgLm9gT5p6t69Gc0vtj+MYmlMmBpODyKeKNxo
8l2m1yfg6zbErRN8e5bcrJ7QiM06o4TXOycWta9et1CQpx0X1IUb7MZZNxAmC4At
r1K35QjBV09GDORvQc2QKdo5yJPsYfTMb5PnR2NDb8kjsMd5C0JvcQGf2gSS2HUH
wBer/A9oTjXX9EH6sFzKey8cMgKFRLEpausH6jmS1zqT0VdrJlwDSM8FXT0d6KcZ
xB6AiJi2VKtyWABobhPbIb7lZ+f9WLydQKlNSWvSAQIcltKRrIuDfMZ6/U+RO5+M
P5ZBegFk/beP+Kg9SJ8tfINQtr1hCHtM5vTw6MNWzVXAESUX0HlJ8vdb8Mye04qZ
4EIUO0yGgAcnZZZO0kkAiTUaUcp3sdPckNzk3xdp4ObFrkTXu68GAKj+QjThWCkR
GK9yDWmLr2FY4pUOwYS/OsdznFDnw69iF5AnUr55z+Kn0fz3UtRKz+C6nZM/s5vN
9trf4eSMEFJ39YWqG5Uc/T9ZOXY47D7I8hjsjbw8PLoITbwi6z3KaDgoWB1r19vl
vIFTwus3xFyiQDZ9QOcF4R3vxhgcJ9YEXmk/1hHoqAB4i6xl/jW5Su8gwBJs56HA
W3atXj4ZPR5KAxTUM0Qn8IgJFGVROrVhI9YgeH3cdfF+Uyrkg0NtClIO19lbbVCn
MuurBmA4n1w0Tz+oJNAz7FtSQnHn+mQCDDg8kykCTh33us1QY5khE5+fEPZcTtC2
B4Vg/bbHppP50voFQOnbGsRFbnlyqjjZlOCDCG1K5mOWRde2YSOybgVKN4JDwCFe
DFJSUIZ0hCnynnArqMDXpmc1NUYcAKrxGwGE1w9jIXplvFN2VwrEKovVv8Cn3bGb
GtQbIF6fzZF2LbkgtEHh7keiiZxW8AGIepAPwpBuj7AdPcOPauAmchDt5ptVAgEX
wnEGXZwLzR4nhNAK2rWfNga95ew2DUQEEmqlsMwCXSydKDyYcfAByKFFjSeaqU24
n7CCJZyYn8luYqSKJ7fa5X3JxxKxmZn9i5mm5Cny15o=
`protect end_protected