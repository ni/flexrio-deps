`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 22016 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
sTHDbAcNdRVMi738hx0vzpYkGX+XGEUVys6vxQBUpz/jMPUeNHblQH+UmFzV9FLc
r8zw+GDXacisz/W2QduThNkuO33PGdiAvG36lqlhjaOtNEvg4dpHWXx3QeWJMXPu
cmoQUloY+CaS4p/Dp+HIUeNNCDcJ1Wp/1m+6/DJda/QAfKbdy16POOFYSFC34fKu
UJN/rvkGzHIdm8DW5iFcuKw6PK4NfKXMhmrR0CbCC+iGWhQavYRqKoOkk7s/iqdx
z+RAEvj2E1HQHrGTE50UQ//IzIaZmZ68ZZ7VuOqATtpeR+XYRaY0WimsmY9azVB7
VlP/DdWnIGTFjRjfvDdYLncB7LyLlTQlwj3/HMb0B0q74AO7VI7KvLl1jWsA4Tff
gQE8+wkP7exycpsh7aS5LVCDgkTewd4QheLC4dlMyeqvq7/KD3rxWvStJfuzUqdJ
nAx5zhJdMZD7YN1Pt/qbV5d79ck7bA0x2oxKbpSAWHaoCAqqv1iKYOWv/7CgcmmP
ol+3bJMZG84izlx9Ov+B1UWEeLVtA9mSXR5y0qrcpZcL2EZr9m8j5HCG9d8F/Xjr
VvathjhkHMSys7GHufOYg92WJh40nwGctZwWjmSHvj0hr53vAltPkV1POtBAhQ8v
a/RpIzjDzJAFDJtFqkkZGIf7TnKWlXhUAWRljOmqzM4zeFPUV2Jm/AQXSqbwMLnH
kUV9+lQxASJ12dSMJGxRu69vRtUTXXRu75h3lj+TTw+rNI7WXHHFJlsnc5KcyZie
/QkeTzLUWjl+6sAgQiea2PYbzcGAF9bp4XTlmbihzw7CyANDrjUsQSjm67aXGMUT
2EV3kNKWFQ50XrLigCDF+m8mKysgRgMS/TiGfBn23AbiMsbPXpbc87KzUJd5BhcF
FLRcEVyR1PYY/cUJ1VnjeoqLP4KZzCHNJK5zdOqYaMod9h+iwUC+Jgev5DOMILh1
J4ftga+1dpXNsplNXh1+9gdjRWjdjFpe04h9MfrFHhBRrexwAmSDxHzlF8SethQD
TjJvHEIRxtFJwiE2yr3RvbP7FznvNCtEoZAsadnMclJSkf9Qc45A46q/jw8JPYYP
1vYQl7XMu4b7RJC7VUxAV3EyhHE4Bbu/4cmtq9OGbYepW7keNb29YRRUjPruXFxc
xzaal4MfY97ZqmENgZBRIDpVbEyZ8+19mzfhgVRAtqFvSkTJ5tnJlTYdyLpur/pj
ao//lOhZW1VXR4fDBGdu82zSPhNhXhMGfvIw/jvPpV6WYSwl9ir/4I1OLTf+kgK6
RrD13WpNwHv+K3LJoA7seiIKAg37oCvvLF03zbyb2dYzQxGUGuMk7OQNwrA6hcQG
3q2YlwYkAw3cBtwYsQrGtvoFRJu7N5uuG8bJb+34G+0jIBJpF2/rFR9Llk9elQVb
dQ0evbw2L1+3UXeLwEG+iawijDygfesLbTqLb2amOryYBlIZ1hfcMpflm9efT8zI
rLmKzGH5Kj4Lh0wK0gbhSQ1Qo0CHSqKqv+k5xg7RVbtEVIoHtKHvkbfWprQDDut7
UVoHsT+IMOmBruVQd9X3H+VL75tROchPBlcXrUnxaXYuy7iY2tkqlcV6qfo2nxnK
fa6UboOhvZetfzrmjOYRLzVbKB8xUUctPpOYPALgP1MybaKISco7WzEXrPokjGPY
8Gn5FpDNraGE8dtz4rIAmvqgjZDRAsNbDibN+NYVxjWpNzxz2NKAFGtmdykxkdQ+
sL4Ruv/ZqG1njQnRLnk/FAVR0yNTAcNUPgAKsAgSrbUvjMhAupJunNkRyKmJdQvY
xc7G2e845CoWi0RaVuTapBxUY8oZ0yTFxumMjGdDRXtd2vrBn4DZNV3w0ywYZwdy
YmGDagWx1Q0RciV+9eJ5w7mPYU899RFN1EIuz2KTFsG8/AoTNJ1wHhC99pF0s9EY
0DygnYRD8d7jE6Y8raxQXg5Pl6QzflKRB6VQUUh/Wa7lmgQrTVCa+1NyOvQAGcNT
lpWZb0QjeqyapuPr5iGK07zFTCZZLRpbOPfvxgZmYTqHkDrNfGPBvPGNKmXF3D8I
bcdNBVvnl058WeHRXILzpPr9ps6W/3FQuGyoTqi+4vOXITd53K4kNEhXtwwQjuwh
yl6SLvXnK63AVb+oSHUG6+H/Y58V7E8Z+rUiBm4p93H3yfuo+MAepAupRLf4+x2B
ahL62vzOMvLZC0fv1D0hEsc7Nttp5EtIrMRtjF0BVwF/VnNt5c/i8+6xy9Ii7u60
VXfMKK6krshfd3Fxywx/y2SZZpAzzLitqYquYI8Yqwccw2gB7/0lsvWoA659H3i5
YUgIKuyuNTp6x4DYxMB2Qbb/xs+ncwI/9ifr4u7OXqSuxuz6WxCa03YwPMFXYX1x
d9MJX41LavIsJx5hc7Wn5Qn7X0AThg2xIb5X6whtXK4QaTkwxBCqMr1xxvOs/pC9
vQcQ5gT1s2M1HUFyx10romdBxsIyJ6GTXR8tf7B6DNb1KqxUBvxVuVoNKIGMnx5N
K4SlVD0cqTd2bDK91cXzCI1LDdwgi4zFcOb0bJ3aLcn4kuOZdAosYEhv/EjNjiWN
seiHHSbhQ9zhJ8RbP26ugY3y8y1wZFxzEbdBXsxghzJS1grs7oy9sRMuBzlkn4Ix
QQJao0L/VyPR4yhPN1/WrG7rKK7Y4XsM3tyFxEzbDrRF+j9tn2yCQrAyxyqQSY1J
jK/Rhij/ctUp4E1hDe0MqM6whhvaSN45lf/+FF6mtyT+LjFY683ePlPbopLw1A4d
AAv0Cno8T7ulhSS4pqGqMbtC/Fuqp+0yUFmzuxLoTyq6peazMR0QGs38iIe8y2jC
EwndOnJUCarslPGNyBb6FyvyXzPH/KBbR4YoHCn5HBq8A3/JsJccq64b990A+9za
CayEaHC55oL8x1Km7kylwkxJnPdD9SK/6zFNgVlKqe/wQE9IS9yKb/WKDfgmjn0d
g3Kjns3c8TskxTCT3B+JS6EfNjSux8RJJ2JhNzqZ/T5jxt43YzcV5BiyfMpvWP5K
8VN9Rx5LEyV59WrdOZDrY6NtHnUeuqRGVdMyyTYVKx6PtaaErnjQ/Jk/MHyvYxN/
UaH0Njb5F/JNzqsjdRKhsOsa58FVtIyHBK6gCYUUJZKjGwK6j8iC2z7XOuQ3SmQS
SfU58rTMe2HW+lgRv8vYMiVr3+BodT/2LQoBd3dwMjdStWfpuNHlNUn2JsAMh4vV
lLjcdA02Aeqx5W0ExrnyC7IpGHov5s8rTwSOOAi45LmZNkrCP+Ymjf3i8q1ggiV/
n/tSqZIpl0WNrk/ZYLeuiTqmsikQaj/pVOTMsd4Vbz81Nhu/5Xh+VB4l9qmOjlqC
qCjiged3+K/JVtEqMNq4ZMczT10yPaEPUixm6/4RtSG2VjiX8e0lScYwFw/10rXl
RtRKoZpa0kj+dCnrf1WMIAF3Tt6xobx1u85QbMfPAM/K2wnTS2kpkfXkON7xIHvu
oaGUuHpIYNqdUD0ARPeyaK+RV05TB+HP0MPUW/5EqVqpEFpqGEbwaMs0eObYDcwi
atVK+/EjwtB72dM01dPFq7RmnWaCQ5nkseeoaeBsKcjTNy0GXFtkCIBXLnYzMbVy
8sQIjHH68LMt2tMrIuiQo0a7mcomfTRbihsbB75p+G6HySpVjvSCpHwJd4iIn22i
qEjMVz9r3/8WvMUBQ7TGx0GW84nwHuYDDYiw0/z7jeSvhNzvM86PLyXgat2FqY/q
hhGfRalXQz0Ze09Tdb5amK4z9oSHhzglyJGKOLLSaUKS71vzWbGyUmGnusp6cG6x
PQDQMvZKPji66/a0nCRf0U9ryGC+/E2orTwu3zSI8T28C8iHpj0tX7dyvh1HDLJ1
nNXNC6V78FMLKO5Z5hbi1a8HdtgecX/KiwejK6wTB73CoTfP95s9kwpzJdc9iO7I
oLg8ekN0BqkFeuPt941vj3e87clUawclosFFbsE2ian2JjTSnLC6iQ9CjL3CB+nn
9O1AXTXI0ZLzifsExiMaaECzIiPa7v8Kv4xexz9pZNVl4CQPLBfb3rbVWHiUAtpp
svp0+g04Oldln9oPiNbMTSeLBOuUlKgn+AwmB7/1vzomhFG4jlrZ/2bGfopSGTRS
9v73V12GXx+kdJHBRefxtw2KExKh2xuD7i4KMpdQplCwBcMHfUt6kBCo3OoUI5dY
+LWlnH3DJzuIwMIwDSkJAhGxjn/gwj08olBe9A7k4xI9K7MfHKmGzBdzm/ZSqvcu
2utZ4deX89UPrzAMkS61odBaq1DsXf+eo3KOb/y2hCMjd2B5PJpqNptPK9qoDELn
Ak5iOoHYPN6KSM8eTUo2iJ1pnxMaWaml+LfizFpI1BiVjWsXyVSyktbpVYknjtsf
CvnHZsKrwOqan8wGUxEnca+AtfyMjHCdMGxKxWkF9wmCiIs+cj/rJRkEbKDWYVzt
+h3MPz9rHsjg3MBd05qcVBvHquFQ1zIuMseZG1TxTOh14MUgKzCwdDavnulq1C3K
6i3JbG5ZH8lT1vFguVva4mJBf6g1rdwqHS1CimYssndIC6BirLX1VOfX5OvDQLQA
zKVV1nclLHHbTtXuZ6qMzAs9kpdK63Q0hL9Flr8nZDgF2RU2WUnZpt6uucd/HBQ5
P1W0CfGC6RrEhEHZZQvY4bnPdm28bgILsITnkpHKZZtEDdtDZxklI5h2gsArupU7
BLSg4bPutvNSAIjcIoayEsa6TNmvJFd23I05zHPB/0o3No5f/vIOL/rB2EKSEc5I
u6IYFSnwnrSOdvcYLm2KmCZbWbX3TmVb/vCr8T9MQ9mYOIWJHhnTj9zY1Nu4R8HN
dxNIwulwS1Kt4AG7WGZrzp2ih4VLHRZ7iJ45xhrXW2efFUjWTnbHd7RbPyIR+/Ox
UwFPsXX6Y4xdJYVbidKnh6TjnK98R3ntCWxIxux0nUmuwmmqAw+9RToeYrEZbmfb
+hPpLVJonAxODNo/eNcDTCnRnH+hRtDtXaTgvQvIwQqinQ8XoRws+6X6ND1w4nho
oniUba1HN5ytTd05ZwyqlfAcM73aT7LBmxuWg2GdUltODVywUA/wnrh/fZr10zSp
mvmRXqZRlZrx/e8xVtp/u44Rg+V1YVU7Dv3bS8kQL36/nmJT/fTj2SXbzOhB36xk
SnC4hDf8Jz9Q/5oNT7ALa5HKr2W4GbxJ0HnRGl6UJEY65ohiIUoXqgZLjA4D5hnc
J0+uRQSmLWp2VrEbLmbj0khqVeLikUfz6mDtLP7CP16DPg4PsvnkI2ZC/mDHJ0Ma
sIH6JcP1vxqlKJm0YVZdrjaaxUqmzPcqYBPvduIP65y5AIA9LJd0WySw0nKo+l+K
/QD0Gy/cWz1Uah+0WwEO59x0q+yK7FH2GQHNulesAJ1m9FppU0T9OaoGQMAGvWXv
G3wPFL7CUehJYG0CDriXt/jyv0J0P7aXF9xk+ssievArJ8XI6NWOlIhiRNtq2x/6
IPU+6sZTmvo5TKTeN7JoH1eLhjG5kofX/7GSevge7LACnVfF70PCIJvJlpWyEwGQ
zrWeKe0dB1JKd2/Q3fANwejYic0rKtuaauz6EsaV5tcOgJNy5dYn0gbLWgjCaI0Y
+3ZKFBOVMN+iS6SHjJxjoAdeFuPhUcNN9S+E2Q3dE4u3UL/uChm+3XORfGc4TcQj
NJP6SdJgjWhzB3IkD5AkhlDTNNP8W42YXiWvgchHoO3aicKoDscoyeVX+Py0EPaA
xwdUZ4yLfDQnyfybKrBBCzvzU4rmJQh+jXEKyw7HK5I8zW6a4avWqX6ykOMRypYd
VH+VyLakIm2Vh7yEQWGLEfrf8qGMptRQ6xvmtvOzMeowNUf7TBMJDIzl66zw42de
y5Y6Pr5ELv2Gy9nFEEg+r1nhB93lsZvAcKJLavLHBuUoYEmFfJO1wLrn9T04gq2m
Dp7uIPgYwEPQCx9lXuo2uZFWpjYk630TTPDYFFkz1lo33QuW2q+NU13ANy2lAzKb
wbU2JAxxlEGOycydLTxoTzk7zVm2mypU73SMFzCdAah5IlBe2tJnRCt2XOSIngSX
2EaoaNIOEGH0frD/1plGLpGkBwif01EkyXZYdSMdZq7xmhK8wUfBBzyjxFNmLxDZ
utK3TovjixKAt4VX/HLWPLYIRSdAuqbeF/3HFQXl9XLF63XsN3nIlDnYimaQ2QAS
eEfGgJEQalvOqonbp/59lIP5RPfPQQO7l0okDgIxhUgLlYXRAGevs/M45qti5WM9
p7WZthLsnbDHZcXPYiWCBKTnufjuc6GO0Jsrz3dRrW1bhzlOjhSGD3c+MPVQe3D0
Eqveqo1iIJBaEcOi2BVnw23I9P20JUqp2Pfazjs+4wfPhJ6WhZ9u0WLZGVcN4GXF
z1GFMNJV9aqL/hp9RQMn8Co6gTv6fW3yXRdL+1ecxs54m8F9pYHPEB8fdu7HJnIT
xHKN74xAGzsvSKWhTVxDXoqbmjPClsQS4ioOjptAxEXnwcmpeRmzyI5mUjUnASu4
hOH7e9XSeUt7q/DIYnZ2sGNzkUBpT4jTeNqYHtWiW0ov0F4mh5rta6ksmLnKt2NV
luy+ilauz2wblRaRbOy0JdVBUQGQ+P6V58BK/FP5IVJA2gqKxbuRVMqO/Do9dfvZ
caPj49NPimO1LwgXIN4hNwEKDRXudiMEvlU2UJjK9EdMugzVkalk2JmvI1Q3TBrt
77Q7W+Iw7LbqouI50pdvtjx5UFTtP2L9H9nI+xQauHnpcwQJYUZ3KdCQq+YgICPG
YlUQaS5TI1L654zR1hGamOXvQrYnrYKSt5lHdsvIQxcYgZA24b5f8p6dgG04RLKs
bhyrs9SB1XqlDHew7Vm18uOAf3kD2xmi//YDzkWvEx4z6nKNip6sBhtjtZXNoM+W
2jRTwxlht8eQgwr8xcBm2I3ZjGLTwlvXNPaJPJ1XwBexlcSvkQtWE3krqU5E69vt
F0HyL/v/ALTN8TgxWsXKk3SmAJUooa9p3dYrIlTNgBcbsmpVSqEptrnPOGA744rV
1D06XXWE0ny1lQSO/cLAqrn0EsJt4IbnNT/XnCzhs5Ut5a2DgJo+pjmWwPejNZV2
KZswx1AYC4PnIUD/qT9NHkp5f0e69tzg8oPVDMgsy515QXKGoU39AaslnZ0xqjW+
QNjp6y49S2AVKGwtRziuMhZHPZnPCoYo1KyUg929jgT8GDZAvo2B79bVeyJYz3Gf
JrFugMrsqzYratSoCkuwUNx3skEKGD6qpaz5kJ8Au7j0dsbsOf4jv4Ppc6fDYNnQ
xQgFmDVx7M0FVGLQoFeK1d9CB9VeFkKB1KvN1HQsOCiOTjZ0YWb2I4gJCeXCCuHo
Qvmx2GNDnTfN+ZHRxYiexYqHIjwzXgmQQJt4haIMYRL/NcyspLDeC0DG6yL8NeJF
9o76CP3KSZiBNiKzhIFhXujbEk/gq4TITLzyY+MVYCXeGUZsOwHsI33COGVaUnMd
+9+6DoQvLhwbVmqF1JkrGH5VTCCYqUZXgDokf9hAePSGI50UOzMlEupoVfCo2amw
2gfR4b45s3MEomp+0A1nTvrZYwLqlQ+ksRsVy+5RT8RFeNsoRjwZWQpxk9hRAVdp
X+PR4osvYTMVpe1PQQQ+nD74QsytkYHuNzxN643YWVXKRK+KqZAolndXBHhmOVNT
Jtr5xQZIB1OzluW/4yncZWnZs9Foc8PygOrS4lB7KDiaIymYIxkoaomfVIdtXElA
22dfHDoQWOLduJPhm5tGm3KQqsXmkBD79B+yh9YDyRvH9Xef+vEON2yx4XZbRbka
GCdHU1MUq+2HAcq17vXCD0sz8Dw8BENW+XX9Mbcu6BgUseZyHDogL1ChoSGI/sYJ
qhXXw1++gPorbPo5gZ0lQpf3889CdHRKgD6WPBQdpxh0S7Be15bANXQS8haPCrst
f0mtdaOb+pS+DUiwpr/ak+BLH1m0ShF9u3XID6rwZfeNs8v/A3QfuAy1NTIRmL+u
ouOYKIOAVNEcxarggB0SOdiXsSDr7OUe/hkh7kSY14u70e7h6lphbegnu/ia+H7P
WUfogUvleyaGI6HMqCIK5f7tXHZxdiGdRh5JRBqlGWh/UsQALKuEo4e7LeVZyZEL
p11dD2LWRRaC6hZ2H34TO8uvAPLrRwVY8w+6vbQ7f2qNi5QBIh4ivJY++Vs+I6Z6
DQzjcSosZp2yOXxIQZLGy9WTiWE48NlMGgZc8idrKSjZZwxjt4AXcUNfCJJBWnE3
8Y/qyOZhPtshzoJCVJ1I2uJn/BXtt6V7+AjC92wUiq8ogGM7ROg2f4twW/1MYSOb
6s3856WuHElDxiiMuiUpx1Ugu6qmSyULQXhEkhin6VO1mWMXGtZjueMFWDPLnYNn
Mik8eo0Zgg4O6C4T+yRRAcatVWIqeAZ7AcY8XJ5Rmpydhqa6/Vtr/mQZZpPoFRol
QAWSAt7A2+jA30YRUmhPTKtOGWglYQmJkV2SdAvdLl5FvGvE7+7kYkFRVbhxllnP
SI2JFBi9ldLUq7igJrqXdNic3vRqUFoG4eVdEi8TAiYHuUKSv10PtNFolTY/XvTP
KtedsCNgsdG22n6OyZg6i6r93tl3oXl9DuHEOek8WOdaxJ2u6q+1vmT1BUqpg6Uf
J7Sp0spK64nP4F86QQCf/4CkUSU/FR4ytB8bR1tzZBXgAmWtOpTxcBDM0sgAXykj
DAUwqDeO2D5jS/ayX5JC9nRVkojVZOI1fwzM2JSNE1vKf43guQ7FcawMhzqekDVc
6qMjbv/qHUa7lEJoL3uFnyMvDaW//b/9WcvekjU26fmWP+fzopcrjdO1dLidQybb
gzd+e71m+kpu6IrisraOYxhbuYuU4G0NKF1D9iwQkd/bcC4rWqjY36fipp1Gr0nb
IeLKeiYFZ1D45ZZuj0cp9ltU4yR3U+3uNRZCmy0qsCkxGqSGMysm6RL1/LtjHQ95
W2sdBds8TJyVEYVgoyuT39Uh70WU0Jkez1hn+wTMORZ/TKBPu89AxSPhqZiyKGrp
FMSWexN3eH17/dGw0DxxGuuXxbqn/yTQFZabfhM+bKrOmJS/tBMe6QysToajldQX
THxD0Lpq1R5a2GH0OJO+8Lb+S63UWOLP3iyzIdZjGWvhQ7Kp7mrdtnSt4ANUmVNP
wLbarvzkCASZ1Ykz0nhh5NL621lIELUqeVWhxe2GVJlQ0tZ9XKXvrRKQyVhi/Pb4
KGiel2MKw7dWfEfZS10K+ZeAMmcHmdYRzZQWu8TqL68BS407q5mQdSbZe15dbocO
1/quCoSE5K3R9LzoIhE2yXsDbel5724MYaIvuYDnLTdFmUaCykJTUbLsIREdRjgJ
YR1nHM1Koiv9A7OKHrUbnpgzSPGGs42lak+G5Nw/1o2npsNEw9OrTwh50Ts0c4KV
PWvKnBkk3cQR4DAFyaL8mCF8x1mLNDPrpXU7cp2OmTZ0y4GO5eHAGzNYee3IusfN
49vTshD+zz480R7NsDSsE1EHRWmI24sbTerU/xqLDOvtsgvchjsSi5H7RZFjTI1N
OSvKW1hxv/fx5otyP6bz4a6lneD+XMjRDKD4kabd8AsOIHONOOhWw346SGyJ2RzU
uQQfjHMeJri7dZn/+4YFL+r0cO6gzRpS5MRuv4Fn1IyDsYtnTyHpdyTy8XFe+ohj
lKuYBMgLbTbsV8dl9jl1exCtqnfGUkb8MLfnXDO7q3E8/yOOrKUbVZLGtTi7eWdP
TR5dU2BUSXiWduF+A6tZ0Vh2CgsuFSxMGb8RJnM5FdvAvUGjcUeEuKb7xYPYelAy
ATYTQnlRy5qo0tIQnGRJSW8jEf6mP9HAs6IssaTlrvSsdn5zmNkRavgfdvpDgpVW
GeXk04UvbLpiVPbEm1ryCph+aQCxSb+erYd9+8dWvXyiO2neEVqVtr3Hkko6sWp9
keJfME+hbmm9wklvFD5LENXy2Tu+AnhJFv/OMPSAdi59y+pGkLJIP9pKkjAI8an8
Nb55Zvpf7augaz40nJ0AEFyweylOWjFyz2Fu37hsNtD3HoeK9lzfgG9bQAjmTW4W
G8BgML4ryXmOgp5kN7Jg0WeeTPb8qc/rSa5B5ahq6ljsEDqYNKqqjs+orNOglbX2
o4+8gP+eNeiRhaGm2zp+BWQFZJkdg0zswIU05o7oWWzWs2PchHyxKAPQwLFlSDWi
HzqKNGq/lEa8JIDuDRBsGW4KiCWtxeOh4/CABpfr/hAxT+NXpls0KOiku7T6NHou
mJIPnY/r9kDk8gB/ph0uMk+TBsG26Dv9MrheFrougBio3suvvYUWKiKYG8I7QXr/
AvTOrO+xGSqrEM8HqFgdQlj3C+ipJnBswrowVTD4TDdKu2BvbrUsKhEyNinwUg3w
tEgSKi45Uifu0/led7a0krJCad+rzhdnSx8Nc3uUHFhe7uimyxXQZxuaqyIotIzM
yVWsZgMwSiUNbyAJbhUBoNzOOtJ3OlvjEjjS2MRNkSYkvJe4U19QE5RmFDGG1l8d
xPBgt1kt7B6zAeKHA9nX949DEgr5gQKatEbVeYTKN7bcpDp2I/RfxBmrb8BxKKDr
g87G4pabuVznpW87TjYYg6Yi+n+cCJDrsWvOhawkK0iwEFCpKTvFco6Of5YV31NC
n3stREm6IJQda6pUNvmqJR0o0z31wbshRyzOoHhm5+BbKmu0QiAGRSU4A7uOfH2B
MqpNG5hDYvYxNnJ/73DCZyVEb4X05UXhm7uPEA95fAw5wVm+1elUKL7cxyMmHMJF
5NekVRwl+ueGtkjtMSI3ppviC5Xad13sfiA4z5W7js5n2acNkgAoNf+CcNqeDnrg
jsAhisLcleuCiTvhnbgpuvdR5vlZ+kbN6ZqAwpB4kXoWW6gaRss0yS6TWsy/PIaT
7SxcG1chvaAAnpWZt43BktK0PJvmBa7Sh5QLnA18hHlOfgvkIr7Vk6DL2Pdzg9ys
hgZAaLh+g7cUldwC5d0hj2WeG2j5QXI9NRxKDFRgAnvbdg9Sf0zqI7BxdWdHxX8X
3EzRyM6ouXdq9jp9UccBARpCCFW8FPg4xuALPiV3T/BNBQFWLn5m3TipFTJ3KA4T
qGEgc/I07kL+CDAG9ckplHfVyBzL8Z5fXJ7YO/NbmLTrEzWpF7yYq26H3OWLr37Q
JPY9Gl1StTl3ztsdPbUpS73lb4W1TGXD6CgeOTLIGevRSxVmGMLBMzeZQvc6Vzot
IPj9A5+RLwetSG7RNQDaKLu8Tt7I/OVEsnpYQyXcMuslcfYLIcwGXv361dYloxEd
wKmEYDDRUCAJWO69piypDnWsiaY43I7wdoZ/zvdDyaAIyfa6AiTEIwAI061EBhVC
9JECtBlQKh40v9K0qPkjuGarxZ+tW9jcmMWNwHGYHVqRlFh4oCp619p93jU/sJBS
L7RD6FMkrgjPkAagon5NzKuLSfUjI1Sd4mP+hmH2Bx0x1UeqQs0OXeBvpsA3tmJm
6rrF0JE0ftA+AxkhB3qbCd68+YZr7aiz9EUsog8gX74A0CHB88fv8f9c3Ig/7UUP
ABsNfstRmRJuQd9bJT2ewNQhVth+I55MK9usU9D1+KiK08Q+bxa0Glmyu+TMI+ad
/oMB+x5SazYHx+Iui4fhPKHn/Fu2UcmLl+Oa31kDraL8xMjNpVXCyLNhkkTYs237
hFETWo9fjrmkvr7Gp5PVadL2mYamcWYZC17m51T8nPFszS/6sw04isxZZUgiabjK
9mUVTEYcFeMfM/15opw0rrXRLigP8TYUwNorzxhJGDl5A+xfOLr58AObrLE23Aq5
/gVivK9A6KmnLOGqUPg4yO3BlxZ9vs6dDSMSHBa4ABuU329hYTt3YH84hCsKkGOr
cgRyjkM4K7WV/rvYtuuMGkiaDRTQ+aWWCRr1YhjMZbateW6+Q9r3Aa0k19yzgaIL
DG/ZV609yzi6qVqMKI3B/Rtg/Fa8svpktz5X/Lu9nDhkOqjWm8EotyZYrqP5+2lT
LAUyqrxKqb8qbgmdzt9S8xtmdDsUs4TwYnxGNonOiJBi73wJbtOQuxhmlMRKp9lC
jeK1qVmMOGGjxkPb/XELDf6nhgO4UXdCDDz2kbaSebgX/bo8F/k/LiawvRJC2jzH
29ICYYWgsT0GQ6JnSi/N2MBwaaME4uQ9xhxGcnG1WPHaeZ1JrA/ePvjztFMtnC3V
89YRcJE2fKrNbPFgEGZVLOXLyaM6g9zzL4IeoN63pnggLs73RRzVm8/q32nJhQ47
fFW4PPeA78e4yKztFyjP2SvRvbYsvCj9fQqAlshqY1aStlP9UaxXIwxQgjb3pQze
ihn1VYmbi0z31UJZr9Ik2fV7xNLRk986Cid/LDgSKUtMU7SBcS3rTr6MRPtvFw+5
If8fMvQuabtbW0lQfzKyaXtTuU4PdAqtpnlx1/725QiPD9YCLo4Bj/y3S6m/xAJa
dnAujk3Q7QZFm3Dm0CmYqFopsMMkb2vVeKpw5VmnPsRJ95d0QvcYAdLT/X1M7BFN
LhsQdstENUECBh4DfN8LSPJrpAQOLG5+3V77ZpmrN5A++HO7kYEPW9AfKyw+m1YP
qbw3ufO3959gk1g7B4a3oeqdmSGoWihNa2KioqhIo7gcxJSWwwplhUB6+qS10p7y
OvVjioM8LwA9C7AsBNCX71PZPGvjd94+JSiLIEOKawpj7Ml3pvHbt7GgNSROPGpl
2yoInOAhZNj7+FYg9nFTSlNycZNexVB+oOrULkFJkYY0VrWzQQMYnv2z3J4YDl38
JdzVd0pODZYnjXe6HoptNvLm3/VMJtYWECtG11wZNRMlKDltHSAJhOhbIyn+iA6f
zsKoBAIp3wvwDH/6wk59pmMWqE994GBDOueB1Cwy84qI5m/1QcrMCPQbawR6J7f+
K1f8Kz+Zni5gxfa20m195YGIn//izajKZJFJ2P6h6Fj9PeGi2jyVkKeYk9RIfSzZ
LV+5bSNDCk+L+rUr1LoSS5VL4bwJjQNZEOjV/ML5UvdZpeO1u/eJe5RmI95i5zeF
LEUpD5OTY/qUXT5+30kdHptFMk/Vyke3xeUwDe0mQUcZiDuF/Uf2IJ/bF4b7R5+R
SeFL+lutx3gq+p37JQtbepDmgj3V/x8Ud/cmChkmoPYlq+C2XavbURgzD2i7YbYT
BUIVB2Trwm5KMxU40UAPa3fPBUlC1vXsqAeYBUhgXTWS31ymIXuZk6xKMz0b6Gbz
E3OXrB7xI4NPcz0bmCi2RO9/3dQ1ZFlKfg33jYeTWxueP5WGaGi57Ta4+eWl8jJz
LXlitEqcv7KenBp52wGMpF3vJw+Xai+QFBkfxPPepg+7BilA4iiwVDkT4LTPncmf
Hy212CNiJiwvb+LyTmPDNh/tzv4gRtRMYkx6x+IU62tvSqrO/MLevFiy8sxzQlGc
UqCx59+wlHaX8KTLNdvvvQdOCQCMUC7u8Khhjtmsq98g4M6CBxEjkIt8OUKzGu9m
Oo/73r7VCjypK1HgkmbliofCGRQBc1HNuY6X/TPis+L2fOBc27re+jwNaaY/+BPk
gZ1aJYH5aEIJV/uzjmGfhSAmlZ3p5kydUe4VLnJNqHJECMarGJaN3HkWhDwdgSad
m74ynt9z+4vUWhoGajHZFNkHOCkcCkWaagJNTnog5WayUePgzNiaiXuXwjFXpjJj
M6Sl6zJlP5pSSHeV2OeTyelZBwxNwKKti7ToR7lo3IKqephIC6CKX6Q8+HhURfHq
HPh8oa9cPGWgA9wNsvT0IV3S99x2/l6Y08Hqu1Nk8Zm8axZFE4KYZmRN2oBUT8vp
pq7EGV6jokb0OOtYGqG+H9xkgf4zGZOZHCNatSy7qiXWlS/sG2tstIQlhhrWtkV8
lTlb3epaGlppOGKuNw+iP0ZiMLtIADNL1maunAR1HXUsp8gRK9HcLe+Eea2mMvB/
quOvFMtlQYsyRzAHUfomghriIh2hnaBbfQiWBFFRdCwU5R/1hYnqCh5e+fXhU+oV
/T+Y1bLRllSz/ZXC5lm7eSa7qWT4OYuRUg8WkPxQCYiqTeCQcs4PfERyh2HL2CJv
Dv3vwnY/4lddZnP4hDSqWxiSHa3rVrWXRNwefJhcEfQ9U+I9iK4KsRxdKLlXD8gJ
h2PvcohKLFyEBvD8diy3fjIuvD4NEs0bYcqjct2ErLqq8YHf/nZtrJRzLUtRDwKc
65HL9l3xbNCj9D8bd/F8OlVJOEi54IHwmKh4g3u+MH59KgAQyo/258VskM5sRmhf
F6yeHUzTZXw9LPBL7uhM/VKZAmwYayZfpic9bQqaVLHMwYEltuwJIUoqhRSHCp7J
v0RS3AoLH47ju6HVbmTfq0DPCLA3UwEG709Y4Ux2iHodlNckcg58LgxZdWkM425T
avnkQnI/UkQA9d5MOvAZgaWYj1fKXmNzNgst8nzjL1Vs57YL6XDPI9iZ0UAy2duQ
V86XasBLDtO0WQ02Kp/IFjk66xD/LHJkx0Zy7ecUEKRRsteJGyjtXO4Kav+QbYKA
MOPTL/qV311E5cRq7Z65rSn1RI2Tye3okGro7+6eybGNhp1BPkVpmgcdtM+erffb
qFV4YBEusSCmNO6U8HMGSXMN4//40GGRSjsFqNBoYg1S0rD/Fbq/KK7BnUaMZeRF
SyNUcIzjtwpEfcLdD8qEHSO452evZHgrNwjLBxfsgTfV5roIM5eO51h5AcboQKD4
Yv3AwhcX+wwDRGGc1xLiQxQWOcP4N0sdxktZgkLBih0vj2nPByYl/IGexpPSheej
hF9xMJGngJJjWRewAmeF8wl7oY5A5r9cmKAog4BsXybPwnXIs8QjpW6hHOAFE9HT
dy013Hx3sW3Sya7FQREHlOL3R9kIVzL4KYrag3hxF6G21Jad7vKK7T2QdPvEpfsN
yD2QoHkM9sDSD/+FHAHjRkDp4QJ0rXu2s6cNDcgvSBWTZnh7wwH9IckWNf6uI/Ib
nWFUkWwokPCJpkwdcQVhHBQazInmoBzdKTuWh4uXuHGG2efc5Y+wtW7NZvCugqDm
MZ6uQ1YllQ0pqZdngnTUOB5bwYZXAzlk6fIftn8umJckVT5T03vuIZUe0jPPUj+0
5e3jExrXKGffyyky6gHI6TsVtHy8koPtkpvPyWBNz+kyyCpb6pUX+CL3wC1NEgnm
/W3P5qGEC8/SZOREGO1M9MClVaZNOOl2s9++oG5fbOxWlB6TbKOgYOeA83PlG9ER
bz4CUWIpycHSdqNPGV//RBj45nHNpeLoDRwNOzrlB1nHWLbveVEd+4ziFPJmyWCG
w/CCBW/TEnv4ABQmh4l4HMdw69fzAOIu6myTTRP2TWHHDK2fQcuJbv2/LksWTrSJ
YthyasfDDE/7f8w0PLzDb9hKGuE8V/ZdA1OgU9brjNzYmKHLinvajcuv9cIIKHWK
WRKCZRSGzzJJykZToHPOKZeOalWygr27NpozzcBhKkt/IO6aFWBKckMH9TzmbJSH
06txRdcoxjdEVqWAuHueUIlziqqTfY090KpWFNZOzui1nc/PLBpuzSVZ5UykWex4
xU6a2Qubs33fF0NGhMr98jzzOz21hcWkMUKhIsSHCFrs+NmjXEhDhLGjyg2wU8+2
V2FOMw1b05/oQ9Kvjp9/DB/+pKTkajTnyZy1WP1b44N2PAFCPHKCNYXKxLAUwb99
BV3L5V+4kTI0LnEUkmfmYuP9pZgTZ4v66j/8UsTgBYB3E9ySJydXy8vWzfSEwtnp
Cl1EwS8AsfgMgfRYz3Jk2NWz34gLC14s3GUFJGljAXRdCnpcgLgJgWoaThDYd1jj
Eg221aytahSZ31hfRonpPkTk+uNRNBL2WFd/x6MzWn3mwNwZJsd3gI7KEVhJc6tq
JLnM9kV9U45SEDWd2QgqwPwhjAy+r7DjM1wldmaY+FajCFfmfJVfOTEVCWsVr1zy
bLgDo/TcRmlNM0lIGKe6bnc0v4MyBofQhUheWb5cnc6s4KI+d0oxHELlKK8PYVjV
rPQaEDdbpOoxO5xrnTnMHpOevnSESOOFgVFFErFrI8cR1cSGRPrZ5C27egqWQWH6
1zWHY7en7wL9sVf4RjDuqY1NFb1PvGebmZGFxNuRBCVplxOf7LgHia4ckxJMXpkC
lv15wCXNihjtgdTfRZDq5TKIgHNkTh5ayr8ZLBObP0V7rl5aOsyjj+V35FVXt8qM
QE7xXkJFKYjvAymcN+WAj0MBYrVaEdvwpFCOlbcUBHoO00vGOXn8XC3fP+kMMknD
kDScY+y2hCUcwx74U/dhjobbp3R4t4NMzn2VJlfK15N5Yh8PyvxeQx8Re926GCY2
l+ajOqUpVr629Pt3+z0Jy5dT3yWAounCjGiwRharDttajO9Wd3OdoWX1ASF2RD0n
4hKul+EG2y37K4UBmD/fwTzhfPZuwjVk1C37dhkTytLO+pcr39DW/W85TqgW08Md
fpFcdM6SrNWHaufEJiVCgn+6cz+jResil4d3Ktf5dqS1vS8W0bNm37TEw2fJ6hLp
7E3xidPtMOPUWQ77V4LAW1phS2Nxe8/t3TjelQn7A/c4uwANuhVV8jNJ8G5D02MV
Ijuo2MiOOc42IWRkygE37TKfGg7/xFKmTbZnaBAH14Kwt5YgbLZLQdMD1cZl3w4M
19dX9GAnaiB0fQrqmomfWYFnPmsAbRge1umFFo8tyOa+Z4oAIGLAw4gxZGmgVf2O
POOEEzxg/cpVcRBI9d38GI4wabsmJPfXYt8hoeyv938QAZ1wEP2wWQt6lINvEEN5
BZhQVjXI9ye2ELs+sH1v1Ivf9OyJ6+1X6Kh1k0N9xXzY5zh6/8h4xQIXo49TOmme
F50nKaE5x0XV68ZOKO8rT29ewMYrQlg1nUputKBntNZKlXxTUo0Npxego1rONXYD
IyV5sYW7DgRew3REuv9o5dWZD432E3yX5egP+cNXv5hTIKJGQt+7aNG4qhFRsJ+t
pOdXqy3ltkVzkf6nANl1NfoR2bAIuj+Y7Ff/T4/S+59PKk+Fs18rUo+ZnkQTUOXs
TwkbaxpVTi7Fn/2nFII+csejiR4ELCyNH0VrPeYDzYwmrfB07gGyCcE2Zr/jgTLY
w6zDw9S1xgCkdPJsfv/IYFAVexF7qAlt/0L9tNCbGuG0cl26UFwKo6atOiJAXFC5
PItAKaNYamRmP7WQYsboP+2WWnJswKJIfgWnScWCDbzzV6ukhXjDESKwnKQxuNaf
LhTQ2lu9344Qdf0wPQOw9vas/AIeYXKo1SuU8SRl7GzLNiPw0NqQ09GZN6+LtYcZ
rNHa3WawDkZTBu4aQhJD/HpFbfsOMcDpcZvl90F6bG2TiQ16jDGu9F8Q9EBea6X3
DKXTZbrP76VKaT2ISF1eO4PHCU1zxW6JbUx273WedqQZYo+QelW+8K5eRRyZpEio
yM2VLzFAFCYd3/iiU4+uZ6WxXwrhBc3slzVgBwz9P8Mlh5B9BrKFgqn8qU72DsDo
TV0JHGBywFLZYGqyaUxaG35xkEXmAzRgZtlqMjERupYRQvGb4597EM9Lk82zHGX5
vHqHL7XSt+aDFFhBb7DIHzHab+6iTT5gXKzWNK0RPhoDrRLgnIA8p4fqDc9LUIES
c8Tr1ano16382D81CUHdbqCY4NZjCNTJ2A1HslJyrrbfo1BTao0lHF3e6YxJTh77
Kf6JMhB31ZkaXYvKYTPgqNpAf5SO6BCes8pH2AbJN76viyNxLMl7CMx+VSpjBt9k
E8PPyJa85phU4oNQdQ/MBeycgzs+rd0TV1tOcEpH1uG63Zm4XiYoIi1XlT+TtR/d
kWnhYRGxS4CKis5ymzi/cdfpyEzlwduICqKTM23CBud7W3zwfzW+px78DEq0nZym
4kpOclhaxmsvYhf3CnxVyx4/lJ028yP4jf2IvzZD3rrZdh7jvJZOsVpu4CbWyCX5
6aMOt1lpemwPcOXQ6rMls48wdxw9lLnvyhqy94++mGu6BO9ExOEa0IxrFPvFKJ3R
m9gsLKfOQHKo00yZFOzJE53lp9mk2vdZAdZ1vJ9OCQU7tCEd+u1URo7TFKLPILcN
MDIUs/hTcurukTD+rTh+2DlLY8gF5qNRl9jKGSmyhh0JcYcSwdb+8SgHBFrAHApa
dPOPIAdPLTNFO8CMk/JJ0IP1dmYz9gKA1BQLxBuJbvyGp7dGWedTKWddWgUcQhuq
LLoLuMsFzYSkixGvZ8yTqF9X/ev2DpJAMxDQIUKE/1oCMK70cO+2tYpZOBSKj3Wn
2JEL5OR/4aMqgBD58BtW0ccoN2yFWA22xHTVon0fFdvwRw5Q5NBHElxZs9w8g5Fl
SCPjiZlkOlr0ORSxBRDtpjk/Uu6YwMyean1ESqEL7jnptwgCfogeNZeULybXZzoa
3/bOIdHj3N9jQy2PRjd5XULRRQmAtam0GQ9krY+Q9gRUb6E0tjpWfah3E+grvJj5
CqLQE44/OtrWlGVFINycS+syqK8rETxObXi4qTbm55nOa/IYPfeumsOmaiNM8Yfj
GWVxUiFTMNzIfACEexw1zK2mstZFao1WlHvgI3wnuVM6CLbdBNaYgcacBTRwLYTl
CSazArW39HwQ2n0jWte6AsahVuh8FYNoUT8UcwPdAAAPlPXC9XZMSVOqq7Hj5KRI
INisenUL86oEjy1eU6gz+9ol71G7w1SW/h8CuykTGrk+90hky33Id0Z5FwXAsGEP
zdeGAONMidUhdHvu7eGPUMmufgJR06b2nSemfotAvcbZool+pcYxQaQXnlsGUiS3
jlpCV3CGpAyw5R7T5RgDfkxkMNNOEEOY7cC0vbuEHuto7MThujkBuxU9IyvVAUD/
IvLOtz8b+RZsZG+8HFXW04ebIVfkwF9tbPSMf6eEg2pmofS8oF0HrWQ69PJZRNO8
qiF7fhtrpaVEXmRAeFcH6bisja2XxqciFRekd/kken6SXTrScY6BE9hFlXejbc0k
hNUP0IoR+dTJ+TmUh4V23/97jc40euNECZEC/QATfrNdNxg7nVyQE1+FlSBURmtk
Q7mxmjDhc+Qa0bO/3O2Mt7PjtOLe+pMw9RfAK1WqF2oNtvPtcscrE5nJb9O+/Fg3
lB2Z2+tg8ueBZDqDsENZPuWD+ZmXfTVIoOq1OePdO3rG0A9sQKXJ8VOZQLat6oE9
4W5Y7qs9Al5lEgC6ctUUlKTsHec5HAWhne8Bgo4bbLmrTrEx3ro9veN7M7J6IST3
pDgh22w13H0qH6cWo2xD04IX5Afay+6XMYa39l1ZNvGxHU8eCgnUTiVGEGJsBU89
ruEg8jtdGHJQWoYJDY5e1qYiehc0bBqDihg1XS9QFVMxEALnPqaGTX7f0xw0H9TR
gdB01eEHTWRplpBITMoaLJ6Ryj2Cw5VnDcJuCwGXpFkgANROfaW4VNlWBtl2ynrY
brMD9WOJi60jmVlPViv5SP3XSTkzOvCnQmuR9KZetr5oHe5X6h0aJIgU8wo2Ed77
jOGUV95g6Qa0oXDSQJLjiNytHN1V+flRvL4hfNDWDrleaI7yBnd9ajq9hyrdokub
uhPXl0SdBfgvhzXTbrSd8WF5/7zw44pkcBYLyFo44jKXQvy+mG5n/FNr3/53X3Vp
cUFmwUxfQGSHXI6VCEYq8eWg5icl6QdZaWfgUAbDu9bs2CrbWy4qNNGqQCyQQ8TV
OQCQ6qhhExahFpJAIJ148uGfcfoJCGOMR/oQxMQV82JHWE5E8jZHC902zd7P46dU
YYhP8Yn6LHBcUN0NUMOX2cVLoYOOSYeyzd05jZ9P45eZ4iHjQvzE/ztG9eEkBhVV
0aRoZTBjlcE3IXoqXWaI81CX37PCj5joVHuryeuZO7nObMOxuhX7Vpr8ddVP/+GL
RsE4CgRbdRwzu+qSQr+uxRz/5w5bQ0Qe39WHWkcaisJhdn29Y4ltbQbcehl/7Zha
wYnCDErw6SSL1Az1wCVQNo6MgL59xqXfmTMDvAXQ/ZEt9qKAtAyPuZ/G1XUKyNZE
kgSzYpB9HnyxlR3qFHZK7+sJ+XNZMfth8zFNvrWG/Af2YAfz6m2fiL6ygalVFJl0
MmLgfnL6X2b5c73m0fwDlunRUv8oAOcPddpeWu2W8V4JL+RJpJC8D6BhiFpd1mHo
vifAmSn81hDT30V4egR7Oq3CjYKlz5s7jqXHw0OWe1REnwlofb2PnMJP1QGi+Yri
o3Z6l45OrBbpHqJ42/jF/lLprLkwhAQohxBtx5QI7C2WeUl020EMkyYT96fHQ7YJ
GiEuSXTL8fQqBxMULJB549RFr5dT581us2MGk/scghSbzu8O1DwTqNVOYwgXHwmU
/Kz3TZeLuyrd/TSq6zVx+PO69NwGGz2TqmlA+nkA1gCmv1zFV+gHV29sWBOtJP3j
EwSLNOtrF+ldDoEScQ5uKMaeMGd5M3b9UJ6sZ3Ix+8jAju9+F1HWTN2KlY0lQTeE
oBVM4sl6B1uoND9VOMusqMEPMSehkirv/Q/SeKmKvoEL7doiAJC0HdzlhHUPz6L2
/uIPMXlWkXPJvYIjxYgv1RsxboU27ZyCjWp94Dgw5uJcGaMppwrGkhZMYFiXDNDc
Uo7tH1lUj7eeWSAHWTM0pVaGQbToTxZnlNyw4yu6tLthyao3FaLewmsyuKMKf2xD
7idMK/yBLNDFmEc+cM9R4lQPJFtwkep19OD2C4c/x6kUwM92SAJRJlUORG+Nta0r
pzHB5R2bLIAFkejr/eGRCs2eC0UDhrl6O1VS0OIlONBbUx8BpDsWX0AeXB957kjV
9jaQKmugvuNJAt9vOUfebTmqA6jfVWsQEhakbZPs8FStmMXXDrbuixu/tq65NTl9
ZpCI4VGrtNIcDIK8FWJZYrkj5H1IUyqRCxbmSHbjQGQVnTGUWoxQqvcI8GSfgUa9
ERGFHGlmqnRdI9EgRLH7IaJA52qTEhTlC6k0jtzoMOSyqGqBZ1axuzWLSwJ5v4rb
ows7w7N7Jvzy0I2c04Xx2X9foenonncCIT13CPlRAWG97C7oVj4nohry4CiQWkDS
3cXc30NMns7iNom6PiSQr2gzlyzgOee7pLNVQFtrV9uYfLzvx9CEWTroLvdnfLvp
3v6D1x2SCmNDvR1ZL9JtPp/X/quEqz2HdSupgTJLK3fgrPEXGN7tihtzvNBr6IGt
oXyU5Dr0+7XMfKs9MUaX5/4IRasG3NCBh5TTMckJeVVv5H6mDjvfR2g2i5IIMlYx
91CxUQ4LQQoIK3TNImaIAtrgqpXem3e/RDkJOjqTUSFG17pcXJta++2Hzi1BdwtJ
yD9RfjtCKJi6kiXm6odrs42ZTCybIAmgZpeCmuvHRqXrqMEmk5Ry4RKthskk9U3V
0ZILl7ziunePO8tB8xnfqfhyDCFD2BrK7ziwyk8mZ+op2LuTgfNgZl6oxRW+1sry
LEvjoIfu6T5f7pH8wle/4xnSwKR3kJMj8oLn3i6MP0er5sTdKHHlxg25Vggx9a4Y
gv7kU8PNHLKRkk4yObDbDNAguq5VfWdc1AcMTr5bUyOjAW7EakMGh4BGOnMrZil9
qsBdfEzAwiegweM3bacVCr8nAJNeAb7TGoGElZCzPopYzePClf94+0AJYRecMQXV
RV7vQDuQZa5/nvrh5sYGbxcfqI1fesHgwY+y9hx+08ZqXh9euGHlcG566/IJjjoW
Uai4YRf6jAhabpkBJtH17AebUFqXD4uYQ7zAbPB4LsdrvRG3zYQGp3kboSJEA+Ts
uAOZFNhPGxMDemdJZVr7XVQY6Mu2s8CeBDYZxlqTJUPDuRxVCkQ109wmd+KZ07mv
P8oRiW/3MzXNwu5fGHQ5dYyjUn7lFQRszXt9wfujYDGbeiG2TFeAs3xsAtzymAqw
X03O8EGO4yKVa/rXZknewnqCrNiXnUX4Su4xoBSIvrU8l5RyyRrS6Fp1Z5sqGc8s
Uc+z42zJIrffkv9E0OqKam45O4OP9s4kmQRwQv9tjfvgKFr2ePk7ri8UkkqltJ6n
8DLPQqjE18TyJUOMo9zIGKwYHRAIyoYk7tqs3mnmU2b2IQu9wmsXazc7s0JYNntO
WmrUh3rX10dUTxOzbhXF04+6e43VNmt0yVgpNiCJQ0rljclX1tl7Kwb9iridcLOv
pkgqsod9sogfqL+dJAzXFPo8sAAG1SZfw4yiM7sgTebxN7eVKUmHqrl/LBdQAzXX
YMtYmBfw4rjIMMP6lN7Zi1yhMZHQP7jmRjTjpgwxqIKcFPs+i2p1IVRHfw6KMQ0Z
ZMZrKCuywzh1CH/0MnLxTC/RdCoqhUQq2KpsGnTlikHRtk2fHv8JgkyX69u6cLIy
kosIWLY6OVNS6S20zbxr7Y986bIsO4sS/TRUIGIU0ME2hacGC2iqpuXCNqjK/YIM
E0cerMYnuRzRTnui1O4dt5/ABmbxWjOqs9wsExjWNalCzTbitTq0lPwD/IBeyjNT
902l3nGdHS4V7bygOPqHLqSPMSSPYQH37zyciNb8f/mSyEO8OUCBZgSfxbLmfG+X
dV+YfjIr5aKpmZLvBFTLUNW4rJ64cdZNM4c0OZ1eaaK0F4RXJxGkUt30J//OomzD
ZXlC0Ktkai4pga+TtDJaUutYCbiAuyCcdPPRwjl/XhFd01Lu7iF9GicPtdZ+2YsN
wTo06g45piAIpGRudOnEE3MHuuvHzmMG7SJIhfbAY7wXJd6bb6s3GOKG7mLwkAR0
VeWg4vXzjXRpRP3GNnP0NDnb2cE1BoveUijwICnXGE7wuK+Vban4iP6jgIZpMIEq
s7A2wscay4n9vv5KAPjcth6r/HYFlIn+ZRMYZXQmbX+oF7wMHithxvNfG1rfsY2F
87ZflEjJqKuqGa/WdbCmTymLq2z2UKh8dhEOG3eUMqw95mGd8Hhs6tp/Kf1nPXE5
YvgpkVyQmsu+WbTktpVpDCZmwwYiWd9vXMJ5cqgMD5WAlDMFp9WvF69UD8QGcUZX
r2u4hVyFj3TOJhxcBI8syDiawiE3PVMOAy7LWA3o0o9+6KQFV8Iop5u0EvA/8dZu
jRl1hQrbgKtAGlNayc2jz/dCxgqcyuFv3fT8Pp6x4OdfaTONTtGLRAoL6QNqxEk9
XgbXfGp8BotMHsXSV/AXygixzLb9OBSXXl1wkgBjdCyl5kEl0TI+W4fjQ1xWf2yy
MWcTcdRHv/WHQGZZFpc95u4JRBLCV/+ejFFW4J45lEFgUWV45dlTQv6B6zH3M1Rx
Cm53M3YTYpx9WGHcOCEI9nwp0OQ5A3RIq1AUXuGJlhX+lVQsfSnBsHQiU3RDcVEv
KSCa7S11JqXI5TR9f0fXk04iFy5aOqTAh9jO47hPdqynlLlLyHq4IWqEbUivi4VO
KV4go8P+B8jpDczOzVNS3eb6G1Sfxiua9k84KijZxJ+CA2y4hL5ewD2+oyCfeDY1
4dfYksMoUemUYov5/d8oA1P+ln6+MfMpyq1P0JlogqFk6dyMGdlo+DPoeGSgfI7q
0AVwXToAaSj7XhACAYSjOlHfxohepJD47ghNV5u9lWLNFAGfEn19vZgs3nM9yzS9
311Sj3ysRKHKEFuKNl2K+cCvO83Reicoxeb5b0575Rjhd2Zha6V6EY0bit31loeJ
jXgB0+jKH/7gC2omaHCCVuidzZwZouRvqYPgFXdfFJnIbgYRjFF/QOJYG4DWZdP2
dlwS386vrAIGWEArpT4Ln/tDIO2gfsdtdTSxnf6ODCtB02h3fAfltqFLOccyjZrT
qebGgo/pwvHYpwiavyNKJJGn8ECWG7QvSFmHbfm/tO+OzXQjy5xMCabYqe29HmeW
qCa/eIBckmCofN6Dg60WZLMKGl1DF+133gftTcNoaOzrhmzRykY3LemaQmhxySmj
3htaQ99F330FQmFfidgGIstYyAcE1P8rzT2k79QARmOHyrxDHyQpS6zjgIosjhTn
JE56qIOwPKZnHkk05KibuWsfYXpOY5mEW9zppn+PewaYjDonJq4Fz9r0XC6mKutm
VzzKwE9e42JRnKfC/rSHCOxw0avFbl1fUdZeKIGKHDP1UbQtBHpQXPhCs+PkA22K
FR7m4akANG4+++vp3Tfe+4qwAMl4QCgtKT8e0T8GKhMKJ1VZ46ulWhpAZwiXHBqG
jp5ivtJqun67F3LuvC9aZNsk4pmNwPrtC7tbCAwCxeBEPsyi1j+Wu6RTdQwov4ui
oVjS7h8GPJW7qCudCEXjXoBdVrf7BEuwRPmeoK37mrlVwOn7wIuumDr5juZoCaox
1kF60MdFSYoMmvP/r0bafMGUdJXP80f1yFaxCmtVT7Ngo2PP6G+P6dLKW8jCiWvi
WMA9htg3LJgFGn3KxspkVkzp7IL+5wJvZAgRc1zjF/MN5+b+rsJSXLH+VX/A4owi
9eSJhPZHnGL/QdnLFsrNKKvJocqbz6ewxj0U40r2T+KY39DquT/qzx43bsgpSIu4
5q+JEJ6WNtFFDmewnsoSai93t63LKCiZDy+Uzx4jcL/sTeoOdMOdUGqr6ksaJWAi
nBUjU9EpX97hJ0YRnITe4dv10hNmMEI74mP3xP0OU68iQLlZyaqS1s9mKjTUjPXi
Pdo1Y9qG8qxwmYhkKp49REBhS1Pw/bpUGnTPmHPQ0winlKjUIO140RPSuALuUNuM
hwyWD7uFfhdQ0MCYyrhcXFOLH+rvtIiCiEdO3NHshiTn1pK2ZakfzSGpxCbGhqfl
tVHF18VHOjUG29v+YXbDweilYNii3S2yXW1lOC5FCm6pwR8o0zfSbyW6GAvexmct
L/zLp+tC824sa1wprcgavt3oNXjIFtDu6jnMmgQQnArhtQToScL2S+AI3zpqN906
HH08ctCzZzM7hBr2tGkxb6UWjyaNpKogpxZKRq6ic8+0P01uYGkpZiW9jXYZ9DIL
jQZbq7U75EMUcexxmvcfYRGP5kqSXT52sc2vyN57MEEpbMPb82ISyhE3K2/UlDn7
4MeJCum1D3AnwP9RB+ibr+ggIMZQwG95CIdNnz6QnRC5pY3vS4p0ltgcnCLunlwp
7UAB8x3GMZJU9ievWjeoPQdx9lU3WJcc6oysMzDoOzTMv2AH5PPmqF/+FDzSPI4Z
/iDpvTc5/GgNFST3CjyrFa0hcpmMOmzxWRAyLSySMuHYI7nKRyFoaJQ88bXVaa3H
+f8Th1iwhZiePo0toTO9wHqMkTO9kMDyX6ZpTqNzGHwNuwU7/VY19ZmVzhBNJi2s
6vpUqdGddnp9+e8u6175YZuY5SmN87Ve1NWsgA5wMIDaJzE0yaIZ7hkdflwgswrj
EvdhZDJLCRJBv5Yle8nzWp5uivlqGlscftSOojQu4ivHxpV2uuy7guq/1zrRz1gj
8BOMmOJfpjH+n/hdixfuIuL/hLYl5wLCGDx3y3PXk8fJJe4zuWzJZym3w3ABS+dM
xcABWeyb57hpveEs9BJY/KMtI8gNjQbIF7WrT6jHaeJnD7ZbLePzM7494E3wNj7Y
09vqdPqUhc9Dj1TB4ERKfl50Pv3TF2L4LVEtNQ2BK9hWaATf129d+nL7uIF0l7xu
qKureQvUXg3/9sTJY6Hat4shdbwKqRXyRBYls7wRemWEfdIt/gXk7ORK81bGnHvv
4dyECPySUI+nG/nFH4clC9OIR1LQQobvJZQenBxadc/w2FS+j8B2unn7O2Cvmxrj
TOqoS6bYfkF7n85lRJ7aFY6DdMdR6vN0/2KnhcOD1kYUJc/gYCWu2V7xGfz/O8SI
mv2qrPtJ4XaJgBfk8z5nuRi58xifAacut/D7AMvViJa3K4lPodlveiLL2nsDkIxX
pRlHXLweRU2N7Cr+Tt7+F15cLrWIdKsX856UugnQ9V+MPnik2XFflcD8Hytueg55
kpfUJAzNUrJCOewlFgswXrknMuIZf3ka/Gq8vgdkc/BEATFaiT4fJ5a5Ik0kGZzH
CaLKKC2kE22yft6lJCuBgA+auDwtqxrrLx+PAjXe0aHmgH49e0dH082TJKl0wD8N
lvoeuYOZalaRkiwgjz2jj/slsyNeSBBhdx/rvn83i5zgsVwh5HWe5gdeZZ3/81u7
fad9DcHkrbKle1fHhdyG28gM+N9saZwQiCeVvQPXG2C8oWm5qaXQ5fcbJFVMZTqC
YgGO3isQ5caZHiU0cN4DuxESkcQRjKqtl/jWkpbIFdNdDYNApo27yqz9S64DZXiO
8SbTmgsDIE5rJi6mWi7srXw5grYkaEdCVtOQH/HzY+iN1XURgwKA/QwNOjgM3Gjz
RpL+cbHX8FZoeAKMA4Pd8HGyNgtprfFz/F7xttHgjK6nsS00S2q77JqAk3AeGEJX
VMOZynBZtUfA/4GOnZ8LZxi5NJtjMQpGFFB8ZCCDsRXvupFCAbffvALkN2vjU/6n
v6INsEb/VIcu7I+4vQH8VZPtJwFsWir9/KRoBAeA5k7OuI8wluXlYTUQ9e7gs1rp
/Lo1ZZqzKY4L3SVZQs57NONRJrZWykDg0Dvmh0Yg0vQa5fW2m7ZXwym8+8lzquTK
BQ9rngxdbBN1NZRMHQPL/ksflR7z+w6Mc4Nz2RkIok0Vt+ETxlLVGNlG1VeqOO09
eu7amV03WqY5x59ahPK5FL2zaIIi018RcpvkLsyLqQKjYfIdtPVqXFzoKEGqAxnp
O3FKo91YHuOx29H4w3jciI8koX502NaZdoiAgYGi16yiH/8RUoeSQumoT/ALJKPG
Wc0JdFKjIIQrCCONLVMgTgtVOH9opQ0uQ5v6vqD50HDlwj9JJT1cRqbO31zEdTzT
QWioOBbXaxlJuuLJh5DRBGv0kChgAhtTXVUPnUPw9t+JqE/svOtCoXtVjSA55BzI
lwMBgebaiQ9Hg0jb6SpJhANjIDvoxn6pCv3+Q6GQWXmVUd7GRfKkcz7bFJEEtHJj
c23pTuE+wIVTfF7R1rw/nPtAKUjCe+RdugJ8Srfdbx02QZTZmdhI8VdH0rP5csXw
RwS4JIm9vrScZcFPlpbcbN1CKDEnXsY+4Ml2MP5lgy/nomjUr1oQ4U4e9O7ynPoQ
A4XbnZ8uuI0QTlWV6y6En/IFUa/pfaRwDvJhMOZCWxWcC0hTQnSW2gQBzb5zxRWg
Whp61rx5N3Y7rmmxp7cx4gYo9qACaPWQXtprELdS0ui7mMsyzTa8HykeYovCVDs8
nIVucf3VpsPZFS+FnydmDBz++ImAYS4NN67x+Y3DDn1Mb+nM1YDjchCroQooaqyN
K1GUWuTOstLbhR6o7FLUIOn47QyZ3rOJ+ZXniPDl4wYjugYHF+G2Xk/k9CeMbvjS
YW6aABx4+fH/nf+O6gFjYDB7/HG0gtvNJ7sbY4hqKMdtxm1R06eQKWuzDwv52ZZ8
cC4yQh+dWR7CDSIMNIEk559PzNta0jB2N6frEGGtHKYP0kOXGnTCU1NtvkYTsPxv
ADzyCZ5Vt770ac7T6tx3X+ZwgZ14nFgYH1W/zGtmKpaA1442ScUGdFeQl5x1X2cx
QyFIuviQtAdZXej5TeIoJ4pSr6ZBe00GC93F9QtNfQv2jZrPHaAJ1TuAyplNM/i+
S8z2HX2asH2/Cvm9dpJhQazLYj0wpx+4VVmL8ISX6LLHa0R9vwdxD4VMhgXpgegP
FXrFNJTUeeIM83/omkBnuah1kZzNzlKLdTdCPdK74w2uL/Ym1hC995OQH/h16JI3
StJ9h0IOnLXHQMWZMKk/hBv9wBYA0YgZwP4TgRhfNmL7vtTmIYCoBYNwXDGosk6J
EoQeEvs28VMN4/KzfUPgXDigs9y1/I+ekEugmHkrwAW111bPpbQ58U7M7k0m7dZN
47j/K9JndEgygpgisFQLHTaJ/RGc326XDI75zdRpq0LsLRdpLyvR6wsWY8bh/eFw
7LDXK/wPU+ETPybHHsSVQQFv1sk/t1KzwwAfOwKfnaoeFsiMy6vIfPfjNPEc42Le
Zl6GCRVrqmYiEr1GoAQ2jLw4kdUbeCN1PRUxfBaZKP6VUcmevJNxJvmqDLg7CTIg
35mM8DV0zIaX+mT9SfKl2IM920o7TpM7ouqoX30HUFwBeZ0Vg1rPc2J6+uzHgSAq
8pJDx73WXos27mcA3F6SDGBX0CNTVeUZt8QNbY7c8eW0tpSSJxj6mnpiQOgeG2sc
0X//N0DK2+k9znOgfG42JrYqjTm0TeaAd3T/6vGew3/qjSmgxoWDzNTwtm83N9a7
rnr4BJ/0hWP1iUr91F51imhwaXA0E/rhg+vxb9rB40gHdDEw0ZP4hKwQDEwoKpSG
Lqwx8ofnT7tawmBdd9daipWnGTUz0tr3u9tpLZZEh3WZfT5dAiITWJp4vm7amWDa
DqG2ZVt9V4x//sU/x88vL8/bc26MC5e1/Q3qwUJ6R2u5EyFuJRO4g4f6ZE2kf2Sp
2OpU6FFHVrus0sH/lArnSJ8pBe1NFrYzHienRKaYKEd8VnWRnPvsFJd4jIus0qzF
zZWPwwCQw0VPBLx4bmtD/IdLMq/Vx5QDgKepT9fcKL/yCu1UD/815pRtj1RHlA/f
Weqq+vKd+C/vknPFv44L93/jdfAPZ3gGO2STTsemNcV8d7GI4MrHIUQwTOgUFF7s
moPIySECQNu/yu3ouNoZCu7ns93ruejJRXS4Uzi1Oz2LM+hceIravGKZapNvzMsb
cxhETi3l4fuYYZ85NX7C+JhYfvGOdjdphI26k5g7ZRLmi9zoj8PiLwjr5ksJ2Xv3
E/ssLbvrED40L5bYpEcc8cJy4IhwevqYWuuUrtQ9lakJvYJ8vFDchLC7deA9A9t/
5r3iJcThro6vHBH/0ScPif3PxsRxgKvky/8tJZ4UNjAlcV5R90KICehe+BzjBy0K
sr6Et7vdYBDYZPogZl66TmP5X7vTA5o5BgQ657qWGWavMfv5VXJ25y2iNsfUF43M
c0p8erVi1nPRiFmu11SH+m0DrKmhHMgoB8C4QycHhpqWdPB03nyHyvgnXV0cIds7
nO1ZlnVgOTK50YKHm4l7OHuAlUFtyNCz70MpZdO9dxOiyBvKvCqhrwAKTTSB7V4B
7Bgux2XVYT+6LZLzHm1z/fTrA6kYlE4wV5gfJbMQ2yQ0zm24x/CPfFrsS1LnIYsI
plzHdsdYXBmIr/z/Ut3w6EOlsQlp8wYB/GIN6M+O6DBNkfyndF6WgAemNHlxHCCl
ev3CSD1LBMfFM6c8s8aYFfehY87XvNA3D0el9t7E/oXCpB+jltTMqSSAkvOn2mL/
LnaIIVQrGlZ9LEkHjY22B1JHgkqOxSOCCZdDlNQWRUO/hYeqNJiZCU39UdQf0UX0
ALEa4lPF5ER2WYM9ofu0MxcFkg+Zr0Z9BaNQMxAY5RuTI6+/PHGBw74YCGuXjF9m
bzHo1SSA4uAlqZdCL7X06ol/w7sX4DKmnc4iFdbmRqFxVI+HjCEO41mVRwTEVwU8
EGhJQ4FJbh/Rc2JLwzrVSjkJ44yYmvaUfADkurX92vU=
`protect end_protected