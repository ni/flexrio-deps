`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 22016 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
TDkIdcJUWDKCGvmrQYRemGHajZb8VlH1TqsfbMl3xLHWnsKDAdXR6qMAVPs38EdU
ieE+l+eDcZUUDFXHs0HPFC/MIh2Dc1etlxhbw6ALx2PUs6SAfO5PiMu4qTl6sPEy
qvk6yq7t9WFw+L44cC1G50Tey1KK75w8OVUxHzdIkpMBGwjKEC3saQCf0FunW1zZ
wZSQipLyOFWph/q9Q0CTfZO834JpnArlG6irfClJNNpL5kn/zvQ3bcur7GsVyMBj
S7hWrY+aNgML7kBH/tK1S40jkIPTAVJhuo2M6nw1ynjICaXVsrk4YCx4HYZ6GSe2
8nCa0BhNT1BnnM0JCYrrMdv2CfZiKXNkSBfxfSfzrj+ilqU9YNOltWl/6jTR9vcV
Lz7kg0HIFMh77cvq0YeEK71Qcr7vm3Bkyxyq7Ygy4eVitNPw/NPPJGixNnsPYgf0
OCVSizRAmnhATgFnTE7NTB2AB5Kjo8VSIDzNr8bBfhjiS6x6SSnvwFEWSHAZAfSb
8Rttcxh1pmBnuzkoK33Zk/1RA5VgIG0NG4OatSf10my+7X/5v9NXmPSELRpEsKNE
zmj3NfaZ7SsYDomHacUr/ixaF3CfRpV6+4IilrtVRKfu0HIAy3gRn/0g1SsCqiYy
V6w1oK1FetNi42oNL6GlBLzZJ69aWs0gjwvl3Jae4IJs5kKNOyUe1+UV7XgBaQrC
3cz+ujppfHJqGRWgajltOvIbpHpX1pMAVhyFItHQpjrygW5qy8ojWoqDlR0lu+ex
ArLNAV91Y9SaMFF5espv3c8hJxACOM+v72RPH19fNw8eL8X2T8ctrk6OJibXzV+o
AZusQjC/oMPMU/jYn1GmwklmSf+0e4OTXkeVnu1Pf+aGYaW6veTVdov7XpzWyPWj
SuzRb+mbCzlVdWRmNUanRkHqia38zGvDhqg2Yu8qlawaY5yBJKG8IcJzu43LxdHe
ngBLk1+gC99B84Mzbx1d8j6/1ebSB3JwZCi7pkQAqePJ17ycQ2yTD43zFjtEhGKV
H3zDCJAux75X1JAU4/MjWgDY04rLtc09l+avQmSkXwq3YvcyoL/G8GgkKQCV+NHY
5Pr7OfXf2Pf9djvi7DcVf39HOEoF8524dUn/7WTUWQ8eMiOEj1XARVGP+XI3RdhK
9VmiBHDCGdzDVUCeJx+uZAwos5yBbTMKnKYmkf8M1jDVYvet6MTCxM5iGz08nnq3
TSjMKzZhIaq+YqjYF9k+Uh+OjJDAuD3W+H8NKdw1c9II1ZDcDSzCklrYVRk/EJbj
V/E1ckF9VCTjTWyKSxVWjdJ6IMYsRhV92hMW/M4nTdKlURYGXd6KsnhpDHeU5wSY
9Obvvbbvf9A6YJyud/nT8WljP/6A8uJcNZel9bo5mS1BQg3gPRc4nHnpcD/P5j+n
IYETLLtAEzQV8rSoxKhDYumnoHbLQ4KNl0BxUPr2rkI9G20J6xi7kz/kbo7UHUOf
pdPz+3JpGpltsavOY6beYa2w9awo//D46vE/MGkOPQGtsmda9CM29lFsI5aYZ2G/
QEKEbzFNPHCsPgj4DXtSyRTcNvCod5HXZg2EkhJQmwXYpr/4SHBzSPD7oRxzE28p
9V+E2AqgzdojH6Co0Shp3SLvaIiBVHU4cwjc68B2KPiqbYztDLBVI228qeJm41jz
eE5k5AFjwSDMFaXe9WzXD9BYosZ+isrVVigYBxNMiIahoiDvKdSaXMOlOvZWd4+/
5fbj98TbdvqkINSW3DjlORy3UVd3UgYHhAOlKepch7p/dOh45+8BL/PUdDbLGTSr
QH1OTZ46Ckg4rUTaBr6ologWJz3ncyJE+cGx2PWAxUd22ZO7Rgh7ogb6yku+f24v
/Pf5iV6aU4mKexGoZUJcuC3QpRz8syy8ZAvmJ+6ah3nUzme6sXsvQGYKjwXkZ1h1
QPjjSLddyVGaoxQzdNTVYedxEq89fqjf0YLlt6PzwGvYGQdZj5QM8ii+HAwn8wsI
eL9XUh/eDAW2BDnK+CX63W0tfM9prb3+nXrPVgYThNVKbOGV+DxpmBYotEx8PRPh
LlSuPmhx0/jImpFtX4PCT/iHLxGbDKOoqXW885WzB9ZWHIACC6pG3QRz49s/lrit
0pfqjhGN9AYFsvLEfgvTjWe4ky9tkIjV8s+53eZOqnsj3d7Vo2o42yoLCf95MPGH
kruQonw2D+BgP7oZl8y04x6+XmAb40SzguR+HFQ3da0eKq7kp3yY0Hu8WOFL+O92
0ug7B3TI/WRPgZb6LRYeSj3Jk72da54IufgcIk9UO1AwM5WAGORDJ3bfr/c0RKqJ
YmDyVPVGV7NxbtflERveF5VvhnXeNaOZg8I6b6B4GjSzEzueESNRs/2FXzf2jzQq
YfUTjmhMuFxKGDBF6cpobv+LHGfU+Cf0yGwOvdVGBupBdcrQOy4g+4/fxdGAR8LH
zS7XN64cMEpVTLycuInBZ6oCho7HIdoqz+9+pC5pVIZPCCXAMYyFTh6gyrjK9CUR
HDkRU/IpZxw/x9dm6NmKDvllckMmP3gk8Er1nO+GNVmZTfPOABr2j6i70gkOROHN
4pvlMz5Lzi6iEgsnMM+Zgzc1vA0wtfMOQljArPu6421L/TE8TIjPVBRK2f3/j1qr
EvJupkTvfCbx+Jh+NI2hg/u8g7oldquciv4+svSeDl6FAKAYk9F6Z3ed0uR7Ya7r
XxbX83qbPdoM4mz8EhgCkB7mq8Vt5XUSDbKZ+Y4OhCvXv4jojWB+BFCk6Fxp93h7
YMWH+HHPQV0/al6gY3TgCx7XMrq5B6lUxWeraAIGdfBGbWuv6dZk8Ff94PfwGqVo
H//l0G15/6MLr6uMYIYmL2zr1z3uUvwHCN530MLPK3uRLcBC4uTYIL0WdrQsUnKr
+KBcQD9OCvt12iWiHqKOivpeZEXLwrfdnmnpRSzKATJVXHtutwmxs4fpC8OuWObo
XTkAnMax6+n4EYBF0XQYSsJEYBRlxg+fa4SCRFf0j7z1HJzhF+6IPK++EvSWRpzj
nMZ6HEN7tCYkpsyhpBef7qAvrhPwvkzMbSObGXRRpqvuwlb3ZGmAB0T4MqCe4ZXo
lKhV5Oi4YS9dwf32SGmtzqwquyN0skZkwL8vsQpnL4a5FHm4bnSCR46W6bKyoIrT
pdfq2fIxObIh+9OKmmA0A9b3TEAFRETp6v6dbFafweNqUXsjmmlG6m6FIz1/x2J4
n7YekauRa6qXAqKAmrFoOn6RrQjhvpQeZbUCQzjPfhD7DbpKmrV4o6a1ua2SLVbo
QYI5UgG7q15juJz107R+p/JQtuVEnTvtw5SmRv47gam37OvWHszgmxVsJV5+XQKm
27Qmuf//PCQeiVGzBLbedMm/WFh+Q8E2nMuBqD1M6DutQUXbe9bFWHCrMRKRscoD
RKi39TSJeROvuxG7FLibXtc8WkwAR09hw0jDEn8QRTiBmPqV6IZbRC57/+jB/Cp9
03bx5kEItt5aVnwYJ0RwCh/4jZu0M3tRYM+BWuPkQIqxkQWIHipvIoMkFMv0tCVE
mzxiKyY9it1Sf6WVvQXOrlo1PfWMrzQelBOSlC8Ijv3OgP5GmuQuuKJ5x2FbFLu3
vhQ4NgUB2BE0iuyx9WGhWM4sR/e0LL9HwP1z4s7UiUm+n8T0PE4zFwE2AcNUP76H
CwEu+HwASXqeDQYudr1JchJ7qhfa6Qq2Np+khcpNMh1omBgyvNoNUyctsnMEazNc
5YDkLc2x5VktnxtsxYzZYI+51RzbSGWip8TbGBRYVXTOUekIuwBSIFrfqTkr4ijf
VYQuxg43jWfzFcnSIvBrYEor3bRfmrRE0OU/Q1CsAsfaaaa5VBnRANkoujZyCxhm
zxf5kY3sP+Q2GFCOLY0lrZc4dL7OYbQxcOkk1M7ZWa1PjJU3BsUqb1F8wPtsxx/D
BEnGlYacNh3mgQOwqy/4skLDl2hpfu7BrIgDz2Ep5bZgDHm3PVqTL0pf1VPXFpHw
aePnfLvKYwT1BxQMIuvvZD47/fCG2O3b7SgFiZz9ZPshIjpiUR2osk/AOrQX6wSl
BRNg+LfWBSF5GHSgUoxBgGc+NPaoiDv2PmJwIfFgkTtikGNasQmub5Y8YcyjwFfj
ppzK8rbQiVRofiB/a+27+TkDudjvCrJFSuIKBqmk1c6XlOpcmTaJNNEUE/g0RubM
Zl5kqmqRnsSzHMwtriIn1CB5K5wfDLTlm7zJ3FefCVdN1yHbCQ80xuqj12vKulk8
euLbHjHOBXUTbefvYvv+TCCToiLsGWaBHWS4Gb3/KJlNh5iI8oaT7qmvnBw4b9BN
wcsoyhAyZcNXratETGmVaGk2pGiGX9qMqEc61TNauYvpIBMjwgV2t7sAMlwlBfNe
nN0nbiL8vhxNmVpMYc0LQ8OPuvULa2qCKmMXudARuWGj4eUo7+gTKkkxjkrIJIYs
XdtEADZXWqh1fUwKc3LGKBue5NeBXX7vaSLjqX+rn8hvm5s/HsLfVhRFEIUnJF3k
W2TagEgfcmlH8i7OZpRYKcF0hPofveYkCQw/AAilOr8eEDvaMBvFNn9N4urDP48X
GmGtmK5KjZIWJTCRH5FQUnyKeFVuqYlQlLbPR/CBFw6KiOyLeyWSZCTpAevOIy6h
hLeokcZ607rABHLm0F1FanrPssEXAeTNIEV2f/9FZ8CS4lhDGyzb/dQ19lMAqpxW
CsUh3jFsfKgAKoDpzoT8v9Wv8iW+vxXIJRv0DAmFYoB/tiG7JGG1Xl2DmBdoS4Hj
oVA4YcYg8Cjr6l0RcqxTsaO/Ge7F4WEKKB8d1p2IQqwzw7PRjSDFR/Z+L5zSAmj3
4Zbf4ZosvukY/JvPIsL+Jrmy765gMI+0P2fItJ1nkZQb0bZISHOpZz6GFVyBFMox
VOA950E3Qii65L544vY4/eh4i0c0E1eJidyicx5A2GrGheTRhKuADWr8mULOoHri
rc02L9eRTtT6S505EdqEDTycm6Z7v6OmaKaYqWTpyCPHoqK8WfGIDfptncUo09t8
HUH+EDZIWZbHxW65VB/MSbAJ0Lv9L9LZZnwyvRPlpOKot8uQWNINg4GOet34OzPH
sRMdyhRNwlxDHcVV3sRa+pMlWSZNBXnn0dX95b8ckG1tySxHT2Z836z1gJ4wt7Ff
d1u2uqC2Api+U6YHa2o4gaMNblmg6X3jDJNnhIz7GdZ6LzmWN5j6zMZsenWntBjl
z9LJq1OWNzh95JbpTHkZLGZtD0OKTYC2Dc1LUznzZytff5hCsoWsNZMS7vRcusyv
oZtUCyHR2xziBRHViIwUTdCzHOT/5pAplgpfO/rAE0XY5RiOfLjUoa73hQBEgWSN
KYWg3dJteK+OPl97TJG0O8hvobebyD9RcY96NeYXS3hnig1h28a5eTUFMFkru6D+
whsmC9+h1zDq2rrsWtITFrx58rWtzLAJDcfOoqh9GQgN70fnFbq8wjZ8vv6innTk
ZbhaqG0DMVR28GF0c5uzEiJGlHMxEcCz9YjeC0cM1wP0T4d0wHqsyRAbmXpfCLhN
xlrfh3J9dxc4rcrdkYHmAOg2FHvTNlGIQLQn3T9khFJAkIta2PxfhTpWoWgthOoZ
ljlq4OMREAdBqwgkK1i7+LP4pib1AxqyaiqDlsgP/HIIgUdJRZ8Yb3IuLpeWato7
pNmGn7S6QcnFfR5teBxrsXYGgM0HI4HiASP0HPltdfBacUnIPITQxPSxzgLjyjMR
0voNprxZab+4bHZ0IoXi3X438Dhugw5DgbYHtHDXMJQQTkrEoj3/VYatI/Qz8RJj
4r4mQV6bxrTVP7TjKMD7Qn7vLHZ45t6U4Ji4yGc8T4ksNVaGInjSQQgyWtSkOlWz
P1VNc1PM9aq+ORXC3g2lOoheAB/PAHCu0mUXSAYr/p4YGy6eRyiWOCV7kHS8/Ys4
8tIdNKjAoj0a0+UQrTm+621DhdTwqvt0DclDfC87qitw9H49nrCPa88PLcP22Gf1
EUrWsK+T/a/nlQAI9FToTPk/BchXsPlICGSUJhUrwQFggMke23W+Ln4OlC9KeQvR
Bnf4n1KBOTWF+UaicGi7dRJ/KwjpFqDlESCcYDoO/8N4qo2QoAygiVAykvGlZywZ
OMaXGTv3NlYv7A81DP3LO9zXUJFOBimP2CLsWWa5WxXGkFax9OjW8xuuT+HEwsFA
xZvQD5fuwl4zUdd0g8XK1SpYYTlYw37zUyIz0tjWRdhKEzF8DxPM8ipcur58TWp9
oe+/wpdqaKO5GbAz8+UDu0YdgZcen303Y1dPTspvBuX4S3wE3qK394lhoSFn2PSD
57NHfkj5VTIRpNnNqZBUNYBOLn9RVSdqYaKR66tv8YNpIJRWkP7WkpBF4SoEXj2m
+w5Glv5n4gXXZzhfJNwC1HTavb7Rz+eW9l3K3SBh72xHTpKcHWICAvsR4zkMt282
kXdorl9nMaNLrClqNVv2gl/zA8no5ZKrpEdyX1CGP9IdpRCWTn4NvLPjyrJUxf/r
PL0H9o/xwiva/xP5t2ccLq52eBa8DAxyJkD+VRKcjk2Y0NbmrDkLYmTtl31JUcD2
/islzFQD50KY5kozew4gK48Kr017GOP1PaHn0vd1jIa89i72YfrfmdqEZp9fq1Po
cZzbTvg7D1gNiROxj/lD1JWUZVSeIjza6vHVSL27w9N8U0n/UVX2LAaz0rxq40Pi
uiQaRfKoEV6b/j0rAd6OgIZA8zMxfBWOq5IzUqGN3uMEc/fPdC1Y6zIlQI7X5kn3
3+x22OWOhOD8OwAdXfdF7RDI19baM1udd48t7cUcYnOuh/hnDhFSuwR7pe+XHJsy
rwBil7DBsUu0eQ9nqicRXpwXmzFpTdotUYwZLPYLR8T76rM9wIeWd5zzPQccOMi3
D+sQiuThpArJidhjT/c2ZbB1j4+tRf9UIhj3Qbs5N5RBKjcIORgiJuVIBTIaXIgd
ZHZd0D5ABEZPMhFCOtYdBIhtvwyLvu8vGRU0tXj+Cfjdn0+x+CNLCPbJY5mH76kT
3njXxN94xoqTQaLpEQVZl8W+KDXMBP4zJHBurHWXFGOx96og4LU+yN8kOABq9OzG
npTU+U8NjIzw+CQ+MvN5IEosH/sMQ9dltLHbgt20n2GjFlViClu+1hNaROSYYpHP
k3WyqHTHianSyd4sWMZ1Q+kr/986UaSEtVx2l4X6jS2FG7h1V9ueG9s2ECjFybFm
mDR9guQLpiK28uUZ5nlmb4VVMYJtRUqiue39KnVe9FF87ONLnv3XUIArhpamhhP/
Q4xnjZZmiAVlo7G4dOPObSonfWlmL3gVzGhe4VyUPkswJq7o1VwPIDziByRNXILh
XZqgWEndd5qgRCqtyqhDe/5KHo0I/SyMjuex/lcSpaH6ejPjh2VzSHk6N+o7eOPq
zBTfkL8/xoVUzHBOyGn34Xd7Qoc3iu/K9QQQLlciZsjWHttNpaoLAePATJzGJp63
JJ4UXj1/KV/zAkxLtYihSNdGKgIFZVm3UKrzuP3jD1QP2RShz1DGst1Q7cQti6rV
1Kt/hYMQol1wQXV03o1uC09IBHXflKq7aUMg8gZgoD7BhtyPyCHMi+RyVGhwmvWk
y1QDFORHo+iOZe1envcoOLOPz+gQTKDv+j/q9znVWKce1SQndo9yK4QkCc5LYRlS
3qNHzA5NYHhM/g7JwH7l+9fu9iO+zQcRYHmwLtcq0MYZPeapnRJjyZvBQOWRiui5
3JYRTNz6MqMN+DfOCAe3Usg4/nGzjuKlcIbPY3iVhyDJehgSa7HvjFKxHeU2Nxzq
XXXhOa29xZLyXAKQrhlgDzEKQ3TMr4U0i/Pz+uQ6RaY3c8zHf6jlsvNsqvbpfJnC
E1XdjfcfUA+LsgnWRCOxMvvr1bHoTstYoGxoGogAnWy9dRLNXpLQ+BFfv5nJBA7S
urmH4hcnreWGg+i4bFchyXLhMCTUMG+AUsFFv9AhG/McmfZwFD1LQQcPEb61ubSl
SVcklun3d5B+DzCykC3mIMMBCuRIszTGuWvjRGUQLqHv49o15PpLv+KVJumY0wor
t+sxjqdOsnj5QE+G4tacZKzBIy6TrgqfD8vxgi/EY7wurZoVaFsjb4McnD/IqeH6
4kiF1yug90ogNVoh09djeqB7aNOGuUHfeiBBBahZ1spES/kwV4saFUePBMJkk/WP
keenj6m1kAMK++gfiVX7AcNPdGh6yNnjCXNQcp12iRRYJEHbGe0zgXQPiJKYGbaY
oiGT1dNAaE7yy7YrlpssEvqRc9Xn+mFLP2Fo/hnA+MXhKwAjnqmxtu/YAUkXlaLu
jXPaQFJQwzOugSbC58/3CTRtsJo0/ogq6mT7m6AwmBQE4mu6VxDd4ryvURQZC2hr
QVk9BrVsFR/QR+4PKdvfY2JBuNMRSYNK3wURHlAk3kafEGTmnA0sm871lHOQp0zV
PJd9Egl+xF0JSsayU92h3SbPkDlKNI30C30tlzQhz/2AbzZ6q/89/2j5f6k3sb0L
F6B0k6jkgaYWXjj9UQFEhwWs/uAGKjqWLTau8kfJeaYMCHF85UXxibOL5ELHD/k2
qGxpQYsVbQkCgMd76rsgWSsewDuA4c2u4s3myByZbOr19x4pLctJrsNfzbHQdwqq
NFVr8bpoU6VQFPo3hErYnM0qOsyJj42iscjxAV8IWtpGk+oXXBH6c8faoFBnddtE
K0aqnhJ552iRlTT3cm980KkotKp5PzWfykKk+8FsZFfaxzxOTqx68+ccvb7k8VU/
9ADkLbyp0IOjaZovL9qTdq7l6cGVMfmgVeS+iacYqHvt8J1/gZAenfJ+RiEl2U0B
sN9Krj6RPVz688yyFy59IW0a82gWHN27stro8aigBkaWFo/5uMjoAv0mwBvV1aH4
Yp3R5/U/yfPEhBYEXWRt08hxTLXFWQgXHAaMClph4eWvGwN4hwMT2gLjpCRUt9Eq
H83UVW4aYDq5k3sDNo/io4oUwTQnL/USfoIsQNYoWtDLe/fCYyX1C/pYgekMyqgJ
GnkUKb32YrDAxVx151Ih7UWR0jr95fZBIQv5sIeZhXxIUlrwy/vvZs8mgsMiBBIx
OJtYLg7pjpFzI8G0/Yb7L60TawdKbZPlTzA3k9zGHVGPR6sSR/8+Ld9NN7Ar5/vf
FrCC1uKqcjM1F47lZd/uKO7wqzwNSM3fAmnv4I2JTxfcVvv6/J1uMC7CP8geldvk
G/N2ReiKqBB3sIlEcahuMPcaJYimfInvmRvvvqvvglyqgfK9s/UIdFy5CK0/TaIf
+6oscJXHIGu365z4Vj5n6dkk1c5vXtMFm/j/hGCGsdKPM+fbQrm/15mmSBycqUHv
p5u++Oryopxoa36eoHkI4Bm56tK4INNwFPMqKQJoQTXHO6VGzfVQc7Nj7Lcok+L9
kziWGQhaF5UPtgz8tdTVRqomCkwJ6grIAMA/f+VpScxjltX/SCUgdFbsxeRBgk3c
tWIOfDAQ0/IOts0GpAQGTKfI5ewZ7AZHwVLUL+gh4OTP/blKH7eTLwuTHfut73LL
5RynxBQ7Hiq+ZpVxy3ditmwNFnxGbC9zT2CR3Ayn6n8HkVt+9RxfWxcEOpYYVeBs
1m5pVLLMwf5+MG9jMiEqxrYzoizM8UPWw7hMImz3DBifADQnpOcDLO90oo78FCFS
dBIopMzqko+BA0KiM7+CgQtO4z3ZOJ2EihSP/vHcKVKTtSUKhN81TjWA6KGPL+0F
MdMF1QwwK6tTl+kYPyQ1BcukOFe7R/Za7VMOEFo53xHXdXixnqt10rfvHLh78cKB
xq8D2lyc8LSKs83HZNzQn11rMU/CnXui4qUYw8fxdB3qefaAnhxlJ741tUajePWs
h2zn1fPL8N6dDgNBdhtcDcZ0tRPppRWnYFI+hiB6k95yRAcwt3aZ0/7EJq84Fv8C
9CzbAOfmDsdydMFDSsj0LrtcTFQiB1RK1fBiZz+4gto03nZY6SLAei7AzWDOpUsd
/HsyAobbAULNhtFuBjLRxtoRKFg0KeJMRz5ZuNUwtDSGI5O2zwGea4E9kVS68laM
M1x4nRyH9U8vn9faAKlwsclvFG4eZW911LheOFlu2NKSgj/cn4Edwq/YX6B/AvSC
P/ERTtiKptTBYA1JKU+yWP1ph3ntBuSTcXYewoTXE2RF3r9TCvBqoFC2NAIpO83f
UKqTHeDivBq1TOyHE3Q/SKXanaTrYcD4e2ZnUkV7tfxcsmxwmeg7n9bNrUuONz0m
wTF6uUyUDbOn2xCNHES+9h/T9bBtfylLWlb0980loXWdvf37pRicHbJELkd7cw15
1h9v/Qr5U5fUAHkPSJGgfkMd38iHIK+2QMmAFlKq/84t8nb3l6luysC0L78rZPP6
nvxO2aBX6VpgIEKtXF65aesT4Ngqr+yZxDCzh5R0mw8U6+tdDxu5RvfxByCC+9kg
JH6yGgsVxVlqvOjBOvbMRas7ai71Qd+e+dtFfnpO7AYmVED42qCG+3x/k6bonqS3
mu0vd5lvxY4FKY/cdYLfPIHwfahTvTdIEdttmddynDfzKja0xc0+MqnQUsgsUGZn
DgbFD3HhCvg1lwdzqdckKH1LsRp1mWwDNJgAsrc8GTbvbrhDdPUB+ycm6Pv828xn
DPBylJPgrXL0VZw/2XC+Z2lppr7M88ZhlZuILaFTwDQE+NrVKWfT6IZG5vtUeOWd
0D4fkknhA+HQr4TOF+NegUC0IQS4bQGXqOnlGeaFb20doLQf7/4yyD+nMjqvhCxB
dEw9oTn6KaFl/vOl73IQCF8GbWtG2KJlsWEAD52RkJ87rhcSYFDX3hoRexuTQxUc
mI01H5g+4Qw+nHrWtZp9OqYCjplhLA/+lrxmAOMT+FM8/RP5nyPAt7ZRBnoXePIF
SEdhEJlyO7DOCa0T2hThe05LlK+WqpLFWRNaFiY2EBZ4xVKJLCBFRPuo6vbnA/Yu
5bIek/hu0WfkalL7WpaP0xtLL7qsn8BQ6aiMESNjI39Azm58YLFQ/hzshPsvJGkQ
hJY28+q5w5GMk4WiPxo2ZKo8lcr3W0v5lXJ7+mm9YdEVR6Yg5qKP49zszUJvRJjF
YpoRavBkizZgbUpxdQsNGWS8yDoyttfqa2BUc/Ss6LmHDBBkfKoPWr3PC6qyaii3
deabP3KNzg/ZvptnMB6CqGP5MWwuRQzDtE2iXJr1q44XRJIFqbGNq5R6Jsfqq2lF
oOCxQq6yBHhALtn2OArB0hPn7qA/T4PAdeMD8rpzxdyfnSrkob8Qq7MOhp74AWw1
AnwOa4ZY9Jv3l28AuvAuocOcJfsJUhW8lHalCh/i51kdm0CldfmWOb11O4Qme0AP
denOrsoL/oa0aXbRLsdVas17L5qKd6lQMU4x+Ga8ftYM36YnJDS5tbKwkttwN+nc
84BqzWdan0mpELnIz0lHFLFYgXJfuPaaGjMdsvfRxqy65eFy/qlqeI3A1ZCIT7Pl
QYM+XmynmUv9kM8pEPaO89UjRtmvwQdZEv7W3J12818uqhH1/7R4b2XvF710sjr5
k9eZvm59RnNfXwWHR91vGDDU2tCafxb272nGlTkFYCapo6c28zhdqaOs1cYtX4RX
0tK9cfOgwK4CLD0RZ1pdW79kZfVaYn3SjkeF0kNohWqkYOew1+bG98XZSvdXknDn
5/E9yt/TnY5JKtXVamjOcNsEbctnh8SHHPGKBE1lQgoOChTL9U5hWpduamURo28x
kspGuhy2th3tzoYD45bVKNxUKDWu0/mTX6ICqetuEhUScr0jdvdrkn0YSQsFDOlj
poTtnctJ++hJOxC/2qj9PVPsgQvl1uezcFKjF96WGOwO72vBuNzwi2249FVXu6yp
irXGWqriOy4l4wYXO7zfdQ/Hn0T/eCU2H0ln5B95wYEm+dcUmt3Ey7p3TZiqrbpu
hWLL1+/u0se1NfFEs27fktb0KwOHuXRGehPNsYRnZ0zQglhaTp6gJ/cxxURFSiEa
U8C3SA/qD1+9cFyPrZpVAvxdEoljK5J6tjAEcvxPVL1hdUQSqPIdsOsE9JRXMW2M
uT+we70/+5SLj+IYEZKMzquNjJFnkyOGLkXyX/0vQz4LsUiVHEu4TI+6KUz0C2Xd
Y+2KCkaTIO/JczWCuWoW+3chZf7BPcWTTiDmhJbG2H4t00xxnqOQVCW2/0juOKU5
BJFvR+cG6zlVr8F1s4gHC1W3lA7n5f64jOCxhRL1ugIW8bfdg+sUWP97ruCZ4rDT
SCpval01lZIfBSSLRV9Uy0nLFDCqxJM9G2UlOwRgMuDLo+G0eawdXQ4eHBdCN2jR
YYS1+wfz9rvGw0ZwxqcQ2/LnyoEJvaxf5L7OLRR1j+0SrEcBE7MZ++C0QYqobEKZ
gO3w3ngSnwyFm/pmVjROl5O3HhynMPf1y6btRTyj02yXpRb/a9CZYLT30pMvkT0v
bSAspVdolTKjU8Oc/pZ1cxJfR3BeFa3acd2Fb0FC1cIZjsdgVIudf5t2R68jHHlN
FVvJ6yOMsSShF1gv0hTAl+hY0IETKUJyEW/dK9iwSP66yX9vjzfHsEeq1EeVXgSC
+qaswxFDjovyO1USNyxEYYV19PpGDArdHocLinvKrvv2xkxzVK9jfIgn5C7oPzya
TFxW2f5AnN8BBR3H7tx2HiI0yzsY5zAfMf64ZE0Zb+PmUqhlXlrHC68ynWx2+gmU
q7p7g9G6FdmBMZ7GVNUxarkVw214s+XTksaPNtO3/GjV3fL4zRU1BAjOIfJDlZwZ
qe5CdTvz0N9WbP52R+TcLl4wCmhyIU+tT/YzHo2TvzfYFk2lyvPhG9s1JiTnvwIE
D9IAZdhI9xlREaVTwegRGXKy5gW8VXubOEH/tRbXVg6N+MMVpOI3epQDnV34AhhO
rlp7vJsu/dWYyfzGYZ2HBCoNiMu+N0S9TsTp/KXj9liwxdMl4JvO/ybfOJ4BVOHK
WMGQGKlA07ldBIg85jaNE1z04go1WrWNMZLkUK5BIQ0DbY+izZK6vEPXDsz+uIoe
s1pSx5BTDfYSHefPkmDrdao/KffLjhoH0kA/azYRKDWbUWhOIUa+yTVynMO4PXsi
7a+xetORBSHY7gq9fvvJ67yD50JyhrlqJlqjprpYWrDXuHDykJ8FtMzpwCxk0Zf2
rNYqB0diqG+ic6lgnrnv4LFlv2Rt/hyh9rIeieX6urLhSVmqTCGUQV3E/nnSslAL
ex0qaQiCNmN+bl5sCsedxS+XvKZU5b6qwl4WHQ/T3VJarRQGGnWcbIO3hvIHNbWN
puljgh5YiwASDuERDhEKexicac+BjPbDmbJiAdM4EfGi3bTD5I2+Adr0G9wlnuAD
6j/HoNmY4FShLlVZs3q8F0gudYmkXLOQerA5j8psIzxce+H4r4Yf7+qwlEFGtHtB
0wXaOy/8PeKYI6pvdWp9uQ6M82FXWoOKxBihp4oZsQOXH+uzD6MRYk6oT9A0EKb1
mrA8t4GBYFtOlXI1WlXpafbNebrBLN//XE6pEf5StRGD7uKV9zVwYK1rK9Kt4gJ7
QZPR2W3mS7FUyduuh512RVHqzL1gKo1YaeaKEz7MrWaWYd9qb+XBrAtscnLWio5F
Z4TY6rvoPTvqTHbGeVfksVcW84QUB/jSMzgv06O8yfIqUfVLl+CcQTDEYw707mPp
m9RbpMpKrML0UyXUBAFNhxbLrCTgoWHeewU5UZFEFy85zXB1B9ABXwEmlstPt8UE
ae8IBFx8mEBZYqYpaehrKbtZFM2k8ZegraZmJ3ypal+4Rd7+EIvSoulfdQsDy3le
x3hom4S8zef7MbnpP+P3fuhLo3aJJMkVp5D3r50qu7V8PFGzDvsCBJjt47YJPeCi
bvNRKyaVgx1ye1uTqUo4PamgDmSyqxAvGczMQcRo046S/VtNRHoN1ea5Dgjsv2Xh
frZ9wLtlC1DMr7Eu8PH+yjvtTgm1TNI81gZIuuv0ANDjsLbmZEx6JBEQwEnC9SrR
f2o3MymxbB9O4LqoMmfN0fVbThOTGd18gAWNyEzODN0fnwHA07ProU3nMpNutmIh
3XXjmps8AEE9kiVhhVaQwvVY/cPy0jKtOEHgeOy7SYZ7ZCxxKZLTK9y0FoshuM7z
Ght5R4WxWnWzRIWa+w8f6wcBuSlpDWezBHMlzTq5KqbrYxNWcnysRqI8Agn9QLsF
7OmFA8wStw8wMHUcl1bumWtPsOoKRyIUHVOzMahff1/ycmNhIpxerEChumC8i7dn
d6pbLgVWkM+EvBT3qkUGUhKnU0xGUwusOsxS/4711PN45J6yI3hAKPZ6OVLi6xoh
DPo9YIKwnWc6kfpYKIffHgNi3Rf23o/wjWNASYd/Obee9OkAHKnqtbj1HRx2PxZO
sC6bHR0Ens7t8qwNIoRrGBmwZkYMXMTuf/MZe/Q1eNo4gygCxD3M7edLYE0e0B9o
ZvgtW7MWIQ82pREbeSHL97wnbvR31RrtrJqbzZbJ+3vqWa3PwuxzHnfkO2kDUBPw
kMgkSdm9JMP69G+dS/v0gg7u42aB2x4B/4VRoQhF1eGWcdAYDVddsIhVJxFFl+le
HmmGEFvJamUQWGgu0tePbevjJ4E3c0IhXfJYTcI88FvMZXwxjvnoks73JpS3xyDt
oaEmtBuxnzJPHf5d4kcDsHPNQ0RMOFWr+OPIi/LqnBlEPOnJhHR3c7CoZY1Ir4J2
+toELtM9FouZzxvQ4SNTLo/Wp7F0lBLQ05eIiP6/5b54b1B7Pv5WAdyWLq8p5gld
55oxu3dcQnbhtvbH6+herfxeQS2CfLyAEifs4R3W9oc/377C8OrGkfm9WtDML0OH
qrzWS72vSGCQmuPJxVagUjM728V7fek/oQ5MWUYZn3Y7n5G+kOzRFHM7vjMl3GFw
uIha0xClzYGRFh1MDSSlLUwgo+5G/ZLn/MWhVzYNsPdUvXy2PEqeHZL7dzk8OH3k
v5FB6DuV9LoyJQezCO+3zyoNVdjASS6LIw6SGeWkezc10TETEYQ7nAjTE3z9N2we
LPtHCOrmMqoBeWjIUwk4igpSjF6xfSWLV9bpDAzf+QJKJrvM0hcJishV9LCPr8+S
2wEU+jrGdin5OMjtgZPtor2uXMjiv0qiWQC7bXchVQ1ZV+OPom/ze5RUanPVPzol
pFJpNMkOwis/PMGs/tY1Sw3QOcFSuMldzIFXLu9NqZYUmhIE13mO7GpkJD4cOVKN
XmORKm6FlVcjNxViQk1zYMbRlltKOcfTmdCggfEAaR8kF5ZAKTjhUXWhp2YolvB1
bTSxBPHUvgVDG0o9280KzyjAphG12Cscfs2SZ8ItFKdRa+FuR7uD0VCXz7GbedaB
EKw8IwNNitOTjoBlr1yazk00ZY7t6W609IMUlgYDd/5QSeRU/conLMq82WdsjF6T
AgGV0yQuuW0BvueYxJQSXcPsi+nA6j8mLd+sgFjbk5nw5hHiq3zmKY3lcXDLuLfv
8ZaCu8OMFmbA9HlEbGthjYUIvItJSeaVa8d8rnqQM6uVeluYKMWQmBbkTm2OjIGW
5wqRbWAbjDjuycwS7Hs2NmUdfl/lrdSLfeXhfUaPak5wVrrJ61OTsgqv1Aqq5bUE
7uO/X7pxy4dwlwatfii00GPzBSqdDiS3dd4Vlq6oGreohnaR9ppEqrE6c5aUaKWI
d1ZWiqybntggS66lYLMpljLARHCvTp8scYjMjunteYrx2mGwzOrNwakBzbx7Nu7u
lJ4l44st3TfCS06HDeGVKFXsH6wbmH6njSjAAXFG/FZ9lCbQ4DWpl4pYZcyEDEsc
fMHvJCGn1za8jtpe2uJ7QgDNKBllwpEM4oDeNrTUNtObKu6qc4dRY0KqriRJL4VT
nXyXIoUn+q68WJ7Vh7EzDhcjNStqk41tO4ONWckx1h8qEzanQE/mIRfsZHtCCX3R
BrXKjOlSrFJx59StNfqVobY7WouCfDzi/0AMoyEPKG1Eu2DOck5Coq2yYCcdQstN
LHS7cAThTp5kCCth8D/0fSJNLh+p9M69o49uKfGly4gFhvdQfEA7syQJw4u5+E6C
KDwLMMr3xl1wBMUsLaFHEfwnRh6nbT/wTcA2SR9xDmabK1N9/PoP0GKTcNg5sQq8
yDcKZzSgoUgHr3tQim/j+xk//w53t/sRXdcQcZF/+959dIqXuMaa4FveCn5Lueu9
SqOqvKv+gJd6WyO6BS9LQKvla4Fl9BxRJHPfMc+xw/oWTXFUMDgrwiB8YOj8MQ6w
O//FMGSsTkvJ+DU3IYh5cdEcNevD11TW4Z9XQYUQ1p1sfRBPvSSKTDWVvA5CFMWg
E5zAaS8SNu4A0urKJAy5jMnxAjKCVXqMOzMVVWpTpubJjt0KoysFzYoz0wp0kQf+
0ZRhWHeeJArsiT6ta9dyGc95uVmXWXzuJKCx5eI8SlJVUY9I/IU/pMs5BzTuXah3
BB49xdc+41O0lU5e7ntlOcy7pqlG74bQyaYQOPHTK9H4zeYjJ6VD0Rfj00a+28XM
7u38dsjOEqgGFMGp2ohMnb/urS40bD1IodgNxBvfCkJRxP2vSZZpiiYXeslh+3Zi
1Nbi1q26LWvhTo/QoI98CsXrML3rJLmUecdVinBZN64O/vGi45/LrrIcUsXtV/hL
j3es0ZMe9kit8kqcXfe0Vv8YDbx9Ov3GeQ3lPySVfwOlB4S7uFA0CG7Pw/69qet1
h2LfEuxfbbuoaM4bqkUOlbmVlK9x8C7geEdJtSL2iur62Cj0K7aVjBbO6Bn8k03Q
DxMuY6ZS2gJav8ulDYh/u9rJogUDdLHtkKxyi8QUGIPcJ57sUJJRXYCH8LaPydL9
+tw6DBn1uhmjBRipJ6wEDUbSyBf/wfr7RX6qhXAVWtJAZibqa5qp0e2MuFZTK6eZ
JBhkqhCD4q0+zYr5E80vvcyqHVUA94GYU9ZgI8O0Fcdnpv5ggcnT2oO2OjWRKzrb
mD4gTGxMQV0ImgZYb1nIKzLHmwxqiu5M9X3oOPXfY4afXt2kXNRwxtgndjfDJq+a
aG42gYRnULZce0M4U//RoymtwghwFNAbv2nHoC5FHz6xjOhASE6gQ7rwxNw6osP7
tK63Y0fOtwPGYvbLooQEZBMs6fKYxxDvdB/18CwrtOXR60/5ckYfpvnU63R/wyWr
10gY0/ucF1sDet4jSwtwSOrQERi9HzvBgVpqahd5LKmfjyj67bbuz0gPeQZkL7sn
n+NGoLM1uDTeJnt6krVwrI9qCyJZryYraLI1z3pUlRFwgiELYxoZCoALBbnlpi1l
mZlTrVpHxeZHQSo+NQ5zrKcXYzCqKvrgJSyVMCNqKtdZpj9H13ldKxDbJnXipGuS
eW7nYmsqcLpoAICh/DBpu32h4aEALoKzTchmtJQ4AuDBvdmDnZ+vjI4b3zBjt8nS
edtahCC4gOstzUpm3LlEf7xJEOWmm1CrP4IiRUr4DrJ/o+UFELdh3gr/b3H1zD3N
qelhkoieIoDntJhbVwCLWk6iTM3LNq3FtMz6xfPOQbLNDb5gV0avf56D1OgETIK4
Y7LpSt+C27ZLLLaItm+kLDwmIzvlvzPTyZYgz1EzAULmCxjoDuv+jetiWnW2R4gT
Xw3eRCT8i4PgoVaq25yXKfaivylXWAwk4rRNSohnXIvNmNeoQxlNzowVu0dpOopV
n6sVZgQa+DNQV65C5AaBXggUtgIvR83DUmwd4RN7RhrkPc/F0NYU0jLuU1HeO8/U
yyNumG1nXoNmURlzzD3nOzvwbmfMnNshLfAN2CAl2/mATulXdD+3ZJxqguQUmRJ+
F4+rdIAaYxykFvqyo2lkEQcUkx7aGtPWC3TaOm+/1lPTuycmnxtMukkGsnp0Cbuj
NrYyfkiSfCKwgAas7JynMTtx7LMNMechD5KRSlw1QIWIV885W+70H9lxUfK4nZYz
2OHZP/vKye/a5w3HmfBdFN4iB1TY5PrbmtAN2hVVvwaizwqIWNSAuRvvNodpsgUw
rpWnTMdKiyoxv1ucmOYky8A0ksL+Fi25fOqutze6gdb0xwawvJusP1AwTJpJMpy7
ORaAoey9mgahGl0XpVDsfFr2ftXp0+2cLVrDvG01Ml/sm365//Z1sbVBJNNQT7uX
Dpl8ThVE7P8aC6mwk0wK6plcuBaVF0mSjClPpqiIaYC+jEIFooCRu3rc6Js3cKBB
SS4A764noxjf0Dk2fpzMYQv5wxjGi9y7LiV3KogdTB2sTytceSQ5qTtwUvckR0pL
xn6GgF6+9u8SR6yZ1KBBcEu6exam9A3UpQSl5AbuCtLIwxNVh6RC7odhlj9x8jOl
53j+smV3A3DFzYrFncMaRoSNROmNJGAGZn8rvh8ihgt56lvB7T9stgDGGJxIXpzG
gu6xNQKOsZdFQavBtkFVjAm9rwgle/OkkwlCO/IsqhWR4i5Cm2U8yppGI8nPnW3n
uJiLh42Cgk8kSSN3Aj94Wtg39rfxw7iJxgiTcCLin8zFsWN6kfLEGfrtggI44Dm4
oXGaQrTBJAmkZZPjzerBEV2B61YbNqOD8QBE1nsP279lCp+8uCtc9SMBGk9nChh3
7ugSLFNXVnuNDMKqQQ/1CFMROQUPbZ9e6/TJVTgP4xa5omjyo2XbZFj7cwa7Ffkb
JDb1n7jTLPxtWQL59R/W7Qrvh9ShayxWsVtWsTU+4F88QG3aFpFoA9KOtrYdZXgp
r6RlxmGphDp5swOxJoUpWvl6V/toHGtClIfR+Lq9jcFuMlxqk4cKB9mqSKHMdQUH
uEtGZnXldG9JIwqGbzBRIVDaV4etQ27v6Nzq8EvhUgILLMYOQyI6zCcS1or4pALz
Q0iHw4WH6n9JLa10up6xCRv0nzVgq0jzgy1rwUmrW6MBQpF8vIQeFOPR7EAqGRCf
FbfnuufCznkgKbG0Np13OCyZQIIDK2AmtsZBvfTB5LwsNrp9vn5Bhw6Dq1+i1g2R
icZJsFciAnLm+3X5VEhxG0BTXtYaDG1FS/tEyXSAL2wErGWdoonSSuFFw6INkY1z
ULZ15XUcQOA4oXC2VVuIebS3EDBhY1XNyk1uU4ruLvR5FLT4juuNECVx7Oh9PJLl
ZNZZKd9P43BtoOLgENg2EbiOQTRwrZjEEHdr52D3L/h81QJiMPRjWsLJ5BX825Cq
9X4HUyBDCxryTI6Vd1MV0Qy1fMQjJqdjpWLr2P/16Y8pVOpaB0uV9YX5UDX2ihJe
Wnozv1Tw3DibOGE9nDVOAM18HHj2/BflqGnSgn0jBA5E86ST1yOHoSIo8CZ2UIVa
ccIFZ75GCNMcH2GWLTO6fuKJsMgOoM6CSTGbI2Fz8UIO6o/+/C30Zs+sY9X20pXK
xF2Wsrb22PI1fWTBkWa+GQKJrQVhDm8JsQULrxyUS+dsc+wkJ4MRtDFrMY2qBHvK
n0neuzW6gaWExl6nk4FKzgKKsobBa8D63TAnbq3DWd2Ku/dQ7lrPki8kUfCrgDv0
99yRCv3UqavawQpQr70UARkVUT9ylrtQb5K08hJ9e660DFm/gZak5XZK//s5sCfJ
alRLQMpUZXRpmTgtqHNAbiVHpBfTXCP6URj/rYuW7nSeCJK/k1klA74PdCGFA0lS
FX/+1rAcThjDlyoW3e5jzzgF2ZH/SyyKJ/NgbfMoP/7isyBN5jdksp9qGKfPBfl0
/l4PYv4OGNydZdsbCSmYNCmHGbcYgewifPH2CEXos7x84GxHgX06ksDMWyx9AU/G
bI8qO8jbEvvQt2eruzjqQ/oVtthkSJg5YWcDyg+zNrMXpMb7yIg4li9ONxijyv0f
DIjzn4+YPYQoJS9j/QXDhFyb5NOniKSS0DoYTjoSDzioLnc9W9GaPvQx+EZGhX00
DtNyZmVrzlH/AqVMl8poGLubZz+ooJEoi5d4YF2rg+N0Q5UmEGJwzWdP87Kkpxsb
qIEhWNnB74TsS8WGAw5OZTEdLFczx82dcBdYX1YlrU6igHJn0PVfZZ//YUw1ewy+
z5xEduL5gpI3IHbfsRaXw7Zi3Oevlf4T3+k1cDUrzyJA6b6qBC3PcxNL8U89w4rK
CWSleBYN+WCoX+E9xlzP8kwwl9oe1owFcI0Xv4+DGAaPQYPP4gCu5eihVWybHqPi
u11X0Oi70KA799tNBEu8E2zYydkRay056PlTk8q2ERjCq3BXt2GUDZFtDdIWeKU/
HxUqxUMiD3vBLZppcBfzojuEYy5P+NCQexUcrsg+spyJBFxya7vm+PDVVMAcKfJF
OXgsgZekzVEHjmDOV4zZsMlYTiVSh0MBNIz6TOXllpmySeJsf7Ggc01ifJ1UKvU5
H1ZxbRL9tfeun9KyOdMkuVepLqnPhjBInr00RdSEeDCyh6wcSlhwJk1ElSCwAptz
BKNvgHgHZcDech4GPeok0HSMIn7xHRThmVLwU3SaDLcHhhu3T6/qgnz00t+NGG95
L/r0SkDTBaqhezFjvBJFooL9Cr16hd3mSIkkZbpvzxQmxHohQW9UaZCI26cz8Vez
f74LdFcyGib6DWONlR8V+jzTF9d8er2/Jb9t1BPA+fzNts9QN9DGnNmpi33y49iS
xph814QbR7cXl0fc4s5dM8YjaSgnyuztEk0pn50RIWiH/kJWtAOrruEgYNzKLt35
0A9Kx5ByLP+JuoGJY2kwbdH6oWYlHsnXLw8hObc4APUZbPMHTezZX4v6P2Fl9J4o
GjYbgx3AGsnFlReb5MBBVaohIRKjpF8qB8cfPQ7P+uB1rCssoSCvnH+Nc5uTFLaC
qHJcivix3TA+FWztJJDmOfY8RTeAoq71ZHPt7ex6Pyl83iX78mdDQpkKo3ai0erQ
4z6+C5GoXPiQGkSlDY7gAVNV1VGcTaVK+GtQukFkl6XeHsrgGFTKgVXpMi7Vy8jY
U8oqUU7XMglu1MabpNzIsoHHMSAF9fpNhlPtSwl4bmYWRrG/gaFxEdK5tKGUDHJ/
KpglGTYtaFnfdoRO/WRzrGLwC9bjnjYnOOUqJz7IJIgPiKQtLEQuzKYXl93wKYTK
53x/W0+iW5ArHkmHJIn0yF/1BJmynXN/Hjo/dQBcHQOLAWeVW7ZXZTvCGTSZpajL
QqMLdTvrpBoM1iOp+ogosEQtiZ5LXxqwqIb27qm6CiHODkQjIxOjiQX25UYYmPSk
AjyEfpZb4qj/GTtLyB4rWaOSWt/natI772T4Hr+SKlYdVeAXifHFP561JJzYtiLt
Nhb84iNEumVMXhXuIfkKixLP+JYCkK+1jqvNYKMtKEt9osj+wwDWgFLKLyt2RbwR
1qqdqlC5242WwsCaHk6+ht1p7IfxGv+OiQOUeCPBtyHgqb2UqnAfbDqbI78aMR6G
4WNDKa26kMVaiV2c74jHtvJZavpzQrENoKaZWEaBqy11mBR3k6MJ+7RaiMQ4ulsf
0Ea/To3fbJNlpBlOZTwJFRDW3nYlC4/hhH8reRMe9oSVodfA+lgRav6/i8zxRPeH
X6DhxEPMEZzW3pnepsHV0RkuwuQGc1pejqi1Q6Uv2MDUOVYC6FxkywzuFexkHB5c
eIFQAOG83UeRVYaa6Ot8Xdg0ZbUQrbSoVbahPRH/ZMU3tjU5iRwmjrY4IzfIhxZW
/ek+F0jcuNFBwRSr1TZBT0/N0vgSWDcn0/d6F8z9hf6TGv8ZyGOHwRoDvXuW22bi
BlYq7Msv8W5FUtJljTIjun6O8l0Z4whKWxL6KbJn2fJOn7bZUe82NHoJDcDEv8Ub
GvSPxtZnznw/ziL14w0ImutNDl9JDDPtMvPbcO5zYcsx7tMWjpuBrAi5VT9xc0t4
FnZTFQlHUG5hORPeHoZg/tsUembVREi/19GvdzKScAhKPdj4KzLDvVqGFgXvqPcN
pLkiUoHijsEi/ek8kMEfkSdlhghIh5s3w8WntSqVMx9AZT+VGu21eIuqEIdlh0Oi
PO3rp8Y/g/Aw7UX4mo4a79GmbPRd2KaMzsYfEj+U3IkjgaFBQqs3mtVyQXZLKf5s
dfM6ir64SfGBu/MJvgGVtYR9kqpe95wfF7At4zbSHmJJ9fWqaipCSWYHhtOgtFWS
m5NoOneWrYH+lzNaawCutpGf+kCPEO2e89gouFjXmT1J3JXmOH2TQUQ3HgFXHhlt
NZ+SgRUwWKTuoogr5Ah5WixGMLgCXACW2AdKyLPWTKLW64EYcN4J+1y9m7IHyL1r
7Vh7fHgtsZRm54bh0AAaMkmHI1QG1WveMcTyBGsnvfJ9c0qyA4n5xmB7stkZwxND
vDoRHjeLzyhG8JBJkijs/ETYDl61208gn5zSqH3hsnlHxYMpE9jkU7uP5NNzBVG1
W0hJutHGkjngRQnEMwsOtJQI45u1+QBYBmjOqKQJaD7HBIR/cS1VaNN4W07l3mBR
QBp2IXoo0pZsuyc7n2a1ygpGyt1TRzHM5Oagv/cq8+T0q3B9eFOnN+GQDE72o8Fk
TCOQwtCygbmW9KLFYttF65bY9SQkXF48Xiiwlkcf6U4BrMiPgvfG9+P4Iq0nkMTh
hDRZHR+cDPSrF/Sap1lIt6pOqZaxyijXowEhhD/0tl0QwMuZRWLc018Vxy1Ssi6f
yExMjIIojhYeA2+pTwduaVueqBuccAiaMT/W8+HAAJWX8BQF133xV3x1qe9+45nA
oThXRkoubaQ939vX47KWGLQyxmiLoL/YP8o8rSVMx9VALBTwDnZ0NPslRHPQCo9o
lqOx28MqY0Zz9b0DXc47pToC/ycWInoh2pClNCMIwOulU2c4GqUFQd2xHOJu8Rz+
WwWnBexBRs+8g5XDst3ROLYUsgQbm1GOTuHrFoltlbSHaUPKplsSAjeAwEE3pNU3
mMGV76NSVdtmKlpdtOS2neG49w5r6eCEiC8mfvXhZcqovqoXZEWP8BCU81WCERYK
bT/KZkx0DSFCFVVPgAWyoEIq96VZl27n4TfaqCEP4C2EaQRzWRt6Dl8bOf1YafnJ
/W/vfAS4/aW3z0PX2E+CYCmfDYXi0/wfwfSrjwWt0i37nuBApfWnpvfjgGektCTg
WY4jtlvG/k41vMtPBrS6iG+Qtf2Pk6mOzDYTIDE5FSgU0Dol0lVIYpGkpPdgCJg1
QJbvFNbG7kjNa62DEEJmfj3Oyc9GmVNym3fkWejpXV3glgebgueUc4wrqXRIoAxF
JiTME/FLki+Cmt/TWO07bWApxxHqX3TKQJucvwBF2OCloUP2x10vvll9/20dpAal
v02FRs+kVQwscg7rsJTeiCWFapxzxJKrkzfGLaC0+Xn7ysUjBuUxj+dbQCcqFWTl
XLK7Nv0zF8DBPzbFfssO6kio1NZcHegaHhVHy+ZEMH1039mLsRso4lDUxONbhsS/
gVDaVglT6DYvP/ZvmkZsFW26+6LUmFoVK6Q2Zm7D5yJVC2P0vwH0PnbSsX2DtmjV
Ptgq7mc7DQxFA8VbGSCAtNRiTrPQC+7tiMKHOnrg+U1sOboTv5CSQ9R1diolXhmT
zkL/TEJo10Vm4y8zGJUrnbjzcjwE/pV41E4kgnITdvRKQY1AWIeCyUSccEORj+m1
kUd5b4QUvpn65CvfgWkxXmlkjm7sRaTukjAhGseCSDkmNQC8OCNz++4SEj6Y4T6v
ShEbfduS12talc981zqMIFb3j9AWISD5/pAwjYA3KDYigFBMV31Yp7MCvAbm6GQI
9hwwBRwszaCE1HBpA5tjZW3+qJ2teaoAgz05E9u1RjjAouR09+oTQSTE6aACWBcw
0GV89VBVaw/bc1fcnsNUmaXf287qgy7lREKUTZLxhHePqDQdYLRY5MC+keuIXzz0
W3+hjw+LGI5Sxw10zvoG7MeCCE0hsoMMOwi2x8LiVurS3WErz1QTndIhaHsihswA
r1qp8OJCkDkFIij8b1JFoVNIEGcLnyEBUlFGpreQ1rCWkcmBvts64Uojqhm3ZwwV
t0rMkvSaokiAK4ZRrOEGaagOU3FsxihvFK6im92sl9BzPmVcs16l6+f7V2bLKmBF
zvDbjTvudGt3vOP7JzmNwg3ayeW43geQk7VIPozfOsbYCq2VOXfApy5cn2PLtlGV
fvhhngm81stLBcnBZQcf2N+YZ3/RZOX4qnU8eMfrw1tG0THAjVYRAXdC7ZUxi6l5
+nO1a6RtHFyHzKQ7sr9rgRabnuGpBDetlHVJz2qaIyXGXEglcBXOEkYBNFOPoWzl
nxaET02eKUvcUmaY8eSMVS7gbJZZ7zgX4+ZsRIIqOGbTVPUTqNVgYbPTqJi4pADK
q4WUApI8Yxb8aXQLN1wF2OyYITWdFeztnpn0V40FqsrdNiNuCX7pbsdraga/pljw
OtZW8FxRAKjVLFqXNZP1a9F9MyGcz4torCcbcYPh6JPA1aqcT3ym+JHv65XKSClf
3hYV5i0+gs/Vi3DcZeV+ZwgRlarkC3Ka4/H+TwKMU5vQSGFdLQ3/UIRq7rHHondz
ud/37AQa491lCGf8zxQZ6Zhfs9UbQjr6g3NDvBhvgfc7gfG4bVnFeLa6Tzz/tlQ0
LBzIi5MOj4i+WAGAysBnQDSLSAOnpl+UBuO8QEbIyT11nfPJB2rXTuUscQ2SbkmP
+Rk+nSNmzjji1lY6KJxOdBretCLzKz77cIoxT+1KcN7jAHhEiqOlhDU+o92XrdJ7
z9SC2rSt3yU52KiPeH2jvL9Q+uDwL8hFEmDZ35WufMYdfjX8aoREWMYcV6aCOK5u
FLYnTCaWiZJnOivM6hwffjvJcbRn9nA0JQhHURE8nnCFnPBownUfxhrYpWnUrGC9
GSDNaml8unCnhh6A+UQCiDdqlOompYYIVHiXfNo+vKR1jfm2Y54Hcv1WnLHFB0DR
Xlbr4GfXDFg+phmw57t2PI2oSOZaseIGpaOUsmAa7POrMlLhXiaZPXI8VDcooD5T
f+5HdHRr335GimZ1+frhpzQ0N1KrRhDCA8k23qQ8E0SwGbRop2AkCakqEiDL4dDk
KMnrsZ1a6wL8Ez5Sa9vzQZ0xQvZZOZKezgQPw9M6JUZ0xg6/HZr6Cm4G3kT6PUPj
PaaY818wiqXPx9Oos18AmfMGLTF4d1iMTc2mBnWygVtBXd9VtTfcr6z9e7LHImgK
JB5c/iOnNjpoeFcjHbIo4sA7e46cZYJq8UyuRHYUXggW17w6aktu6/mvYKHWPBnp
wJEWLX1Rk7J23eCiD9tvyH+W0mouCYhL5GQMcNeOUFKq9rLVqY/1FWyLM7VpKOKD
voedsbdkOVWmXl5wxLu7Z0ZTSaJigQb7o03LV1xYYZMRww9A7SSCKasYnR1YukGQ
FlYZoLIiELcVwX2tV6zVLn0cxtcF01kPoMH894JHevL3PRxUny9nPgWt6mWjPKJS
U7mP/w4Gha8LHyMsh0JPUWIXtC8oJiRGPuu2Ba4JPoo/SqiRlSNdY+Es0TXrRQ+6
+fRckC3D+I7OelNl3pQISI6FfvygN7jiu9MFFyT995BQ4CV5hEb9Y6UX9eslqXXr
ggSYheZ2JbMl3tersUHtleatW92cgCjI9l8UXDj/ehnKx269MnqDH1/KWYXyZmjE
61uofUoV21DSxiHRM+a+4+oBMr3PQBvyoazxbwp7oAMDfEGzzaURvKwHh/e6gC8P
qfl5w0zZw89Hy8+qzyVqpBHB1xBZf2oweOD3FAC/xEmW6MZQ/iGq0kIUs/N/cMLo
AGVTbDEVKFIqX4S3YW0Sp6mAhKgEnz9a7KgGTT8tb8L5ScLYPwA2LTWdvVLc/88t
CU/SG+nGEkIepq6ipGzJ6b2G4K6JdAVvMYMXt0Hwjlo//qnD6SUVioMDlXfyYO3Z
pseuWn5GrQGytcoxeXcPX6wiWNO5b7276znuuSnr9ksDkhvnJ+C6jZdZ55EFydO+
20KONkgJGxNSqxJdVr/l7VWMf+sFrepfrarPrHdPJQAwoqVxqcCkY3VRcAy1F6/S
R0J7x7CVKTy6coOwiWN+wVGq9kQuE03UVVFlCQF8uYJYfmWxe7A4QlNNk3K0+ZEX
7BAzu5hy9chsnGcXpJfGVwX9PuqtCaNsgNfr4OsQjnCeut5m3PttN3ZeVHE34eEe
NOaxbE7JffWJrg5Xd5uhZB769VWYwSSksUmHQedOlk4qAprosTztiq9+I3jANnQ2
0koxD/9plv4C+vDldJyweHkPfgnlTS159QdiEjnEdvzgJ445VQUUXQBowQi+r8Pq
XxSe7Q0clXp6N3I+T0cdiid2Yzc8wrsRHspu+d+2KHMdX0cuMcGZ/JF26Fgglo5f
QKhFU8iFdEA6iyUX8+0qhPCf2Gg/OrRbwrd433vyO29T6IMZM12f3/FbBvqcDHJk
qWKas35Ha4tpCF5A/gsqq9ZZ7MJZqiq7loV8am2SO7BzIuDQp9uUtSKsRo+p8BAM
Mopf4FdtrJXHx3KMJ5kJEHb27jISVdEK8VTakcPA5T7kW/EGAupcfU+PA6L9aDry
ET003SGGjBo3V9jBei9ulTmA9ERXWVPy001FvJiv/BAarDRv+gatuMKy1t3fTiTM
ZY3tN60X6Ex/kE9cuWs65yv5Cyy3do6ABOZqfxtKoLHh8uOChCqesc9CW8Ct3E4B
EOXESqfNw2m/eQ2V9Ski+Tb++zYLh/2nBstegq0NdnDRpTqxx0xwM786enmCDleE
S/sngTYt4mhfqOMu0TLYS0LYsSMORn3cFWjPQfd0zNqxRKQPka6be6NKMA8opVwh
m/LDOTM8+L7gZOr5PqrReJ6GQ/8FwxIYJayIP7C6vaTWIb3qERPmJLPPnvHK+3UM
ivih97ush4AhVtyTgOOodLUxMOOrKZKS28lrriPCDCPaMcpMet9YuwgZV6duWmQF
8cfgNpuENQZW7S4GNqHpLzr5FpAXU57IfbbdgRWptZoKg4+Fzrtl5axfK+ymaTqO
+ST55j9HXJAsQ5gFqQRmJD1Ap4oC0TLe64ImP98xR5BBUOrggru/Ud4zgcXpQeNM
XuGbNpDx6W6wCCy4L8QNqLHUJJEfj9bxxDSnzHxRL62/cx0ygg+Nc/+BUvfBLMo8
pF//8IlRVu9UOsQ+kP+g0P/rM8Y0/3iZxjS6UjXIBkanaS8SVm0xGQbskvP29Wbq
Mfo63pRsNIi+bpejDWqFQj/8FUn8XPUY2u1nnIL6JrTNHBiXce1eetztoElbxnPs
XcjzVKy8ril1fWktPn4uEVdxiiyZKc+gCbAzbHv4jrnR7UXSaHUfULtJGuTI+qAR
uiQSTmmp66W0jJm096xBGf3GYrt4plrMAp4hk+/uNYbs/8A3Ry7uAQ/Em+E8qDX2
XixiuvzkQ6xIAvLI5z33EsMBkD+FYH8F+bDhI5J2Tl9btnRYWGf89kbesYbJaD1b
hPbLOYoFf/F1t5RTDIaHQi8gWWymLskHGRoKdCJkoyyvRCc2GNSBY2ElSP6qlcKI
x+DGp5vUxOC9F3TdQyN342XlQ8MTfh7WLVqVo1BScU04F4xGDuaa5z9VO21chrir
t69KiMNwW1WaCPr11DE+R9R/yzXC9p3IYJhXM8WSutbtFhrngKWCojGaihuXWSYa
yPlrDYg0xbHiRI9xwlRQy1RWwr0+xpOoAID//R7XG4ScGn/VVBqgcVDEeE+FfB6X
p+ntYS8we0Tsc1mgdUuW/UDQi4sjf6RkZVT2vL2iVCZyBOTq/LF/E4Eg84qnMxNM
EVIzE7UrYrqsKwB1hVcDt1081T19HVL8BQbal/U8+x1ksgpMHuqF1uPF4rd8DW94
zaD6yyxMdjFoquJbJLXH/Zd4OvIYZmMUgtoaw1Wygmx6Dbm9KzU+XrZ9j2nFAFVf
ILOLJ//gzERo+VkrWMAkuTLoaFAyjqkE6Ar5XJLkfvTnNW71gQz1Dq9c2X7q7XqY
AVO6q3vjMH38cyz2RFskgfOsGblaqfKrFG1kM42RG3+ycG+l7rK/s0B41gEv91xJ
7gJx3d2OmEC5FIpZNVEh1lPJQSNM5Wjt0d3cL5/UyoUqAD7t9HZMhTAmCW4qr3Qb
fpENP9diXYQUCxf+7GUKw7M3/9F3ypWXSuNlzTn7TUpLfBYJVUJggpx6vLlZ85jy
xbiw3p+LuvM3N2hCJnrWpkxsxitRMSwpnrq5wyRVHuL/LymbbpSFOFNqF4cfdOt+
8Nl+n9r7C0Zbv7b1t4rBGEugETRvotYEua+b/Efxp7kB1FCzuvvokZ34AxUIU68i
20kdmwZ1A2KX/eVNjLazHKp+BfByTcBK7V0UDGX6p9ES9/Llf0fuK58OUAfc8gsb
0NfNYRz0niTnMjJLJTnozYRSzeQVwoytDfb/GJPTEaHkOK7C7EDedCBYf133PH7i
jCIhSr5K1WLyDkCdm9SWPpiFYEoQTZL3DSNiDlQ6XM4RnUaou15MDjPZesy8e0/L
KW1BvqWap7lZYf5rD5nVlWv7ly85+qjilYn4CPPfgTxPO4OvVpL1G/5TkQq+SLI0
q9iI/hiL1nuwwPk+fLpLsD61U2pk2W5JuyJvjvpJdeZN3LkjczSHhgJQUzs30rI3
gMlfhQsdBRFbnuLQbvaJ1kByv+O2z67ei37+2YtELw9PEwYniLUTNNEXWrJiglj0
7fgtdNmKg4oqtoeWfHa4GWUKREtAv2JxA0tjCEGI1KI89w1PnpGVNaAl+5aRwhPB
fBmHhJE/Z2guWbHButirYBml/F3+OYF7x2DbYIs/T5Pu6VFO9YaWfdBr0cDomXFs
b5I+d/EDznQH+g7/Pxkn+jvSbW2/RKZBXd7P0893dU8V1Gka4zZbYcVJH3qUEzu3
LUHwMQ29RnFb7gH/yvjeBEJWcyJ5pctAfUix4zysOy5Tfr5ZJyR+802gKmtUhcgi
9tdX4ndtawJBbmRODsGV5mQ/VcjbxA35eiG9XrcAIQ5KKF+DiRKuPAiVFs8T0vpb
l8n7Dk3zOdi2yPiTFvcU1Tyfyp/YGwENOHD7SdnBjq4E8kyhjQ1pY7KmQ1KGHqMh
Van4hZ4G7PYb4KIJxM7miUT70VYsymYGwt2v6/8TLmZOLxbVb7iAmF7Bh7qWtNQJ
KeArI7PlLUZZEXflCnTxWxCFkmKB/aVRitC2R/Y9Qjh+/4h7tO8BIpG9xAaahHQ/
b6FJ2x48xkULMsSVUc2+IcP8kiKiXm2dGnKwnezUClPBUeQsZHHB1aLDqBJWSwYJ
HHBkEyOf5JHjkMK9IdNn11BPmUq6wzQEIXCIeztvJnix8Th/9OHAcGpOXWGbMt4f
byYztk2icIHz7A+mqc5fr/odw+ZGUZ1Wl7JSfhGbjQnJ+T6Tl0BIVCySmAt6UUK/
GqEIZHWYpFwWYICBCAR01/3y9WZQNqXf6Y2DtquEHY/O7fUb1Vcvbrx38KJb6oKP
wfT8pN0BT828YMKc6sTedSMxiXZrzwJLomw/Bvg+KRoQFwEyt3z0rJ15MkrdLAPO
Ge2UV5QHooWjEZtoqHwo5++uzqcUc8MpFcVFU9lnGQw=
`protect end_protected