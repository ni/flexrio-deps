`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24224 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
Ju3IpcJpVj/VshHyynUPTOEpOOFM9TWog5695c/TI/jU8JfEYrX6IaW7OJ0I86Vx
SbCEYJqlmAg1xEEbm6ckdTuJ1Gk5ALe9u2OC/ADJK7sykP/ZGOPL9zd3FWv9rnBK
lPwAGmSdmCPVTaNJl1GyGHmPVCqw6OtfzLpZZQ6hXycDLvBGjBz2/X8J+pm5ybTK
mnYFO3YxLdPH1eWxvNUJ3KJ7kf1SH11JokLBKfqciXbZkQi/+QSQE1Hd8Q53eFRe
zRLG7ogJSIBLZxZcfFVVK+PTDuETyjG6FUzYNGIlUYOxSfzjQR4gEABlgpLBqrf9
YLPJmjaARDXto5qYS/TB0HNGV80a9sCsv9733zJHnSsnH9NAxLZPYmq3CRjNOsoY
WI/EWpY0dQGYNfzuwQdX7yB+OK58EEni6UbeO/Al+wvGn35Tc0/UIT4cPZ+UD0uu
Sc4+Sa8fiHhM+ZqVDrc/HcSSl/AFHIDwCdV1Z600u+usrEOp1PVG29HOeTubJSBd
aj/ANq2tlJe1LqUC+TIy5K1tJ972oPV6Jdgo9Qdt2qV0DCL4OfCgd2IKMijZ11mC
Y+l6NiGgO6TU0rmR4y1PmpNh8c0RYDU5JT4uRnTuf44qL/yKc/sHxYuGUfZrtpU/
51AuzHDKJi2UVwfxrMS7h1zp0H8fBwb9i97TgIb9o9Qw+TVP1tgLg9Z1hJ578kZn
gBikhV9HUXXAFrVCokGOsrAKI++8Y6WXQdB5xHH1Pb9RDnoKOMWjTLnQ7rgtKCDq
rwZVMkPdfAUhWvB93FvYSA0qGenEDWwGqwvB5j6e4jmXj+rRTTFYK3O4+cz7AnqE
x7ixz/dnafAmDDNGm+ljOwktB2ONbau+KcVwD2ckUQvjE2z1KyLNDVlwqo4a+0Nv
Xoq1pe4kCeR3VO2XXMrWiTiGhtRhdiYjLQCLkGtEkRmtGYKyg8O/azPKUV/E60on
hWPvs5oVao6dzEje8DmKPhvzwnViXTAcE/0w/19xHGKVBHig815tL4HPdNa8+hT+
x9+MTM7IqW7KDwyWCp5x4NlYgLlg+c7HGQPjyWahF6IdyTTp3Ib7ziDPSinuQJ7B
AdkqBUXddr4k+TISOaSFVVgrKpxG1BOT6x2YtDWBpGGkMbQck39SJPWQgUbJfrYs
Ry22LcPc2eoEISZBo/38s8p/pTuy+Oe2VsABUKrX0arhRuMUo7RzxRkXTkDcQMWK
XSGDDzjVHfX43U0aGp5CXd3v0xj8ZAR+66T9X1FDtBsa8mSaHsGfV8fNC0BP57Jn
wuwwlbhiBTUQXeDL+H9FoH2MqQm9cRrIBKw3XYZ6zIAluFshQ0de02sLM20Ux0Ym
yaVuwvLJczS8dnV5nReEN96RcXvPtDbpJroetnmwyQHZ9YZgfZJwFT1vuNMKut0e
VKg0h0qoLz0Kum+ULIq/1u8XdrgoKQaQ+/5k1UUTh+ed+VXlXQpZeTa07aa3pxs9
IHZuT7KXOjoR3GoYqUAhEd/OAKh8adxfkkhvfl75SFgjSQRtzENvNd6X9xMPToIl
tMDv+LnsLFl9QiScud5nMlOP8fxSaKeepRecagZYyoHi9HaXsaQ91QXz883nxO3p
Evg3GE48Qjv1vtvweAxWAMb+DmjReCoalYxXQCOF6L2LO3VBflnZ+IyMcy12554v
uzvhQk1k+sLTqjHC6L5Dik4fQ5wUV3sue2hYRiWN/WHpm2M4I4ldIfmGSCB++B4x
n/LnsBDHHq00cl6LFoeAOOA+zXdfVfjjmlghDd+OSfQB7mEQLfdUX8knGW4HvJVj
wnz8nbGnxyJqo9hI+cn5lVo+Vgi5f0c5J+37mGVrW57WCFqJY7k73Z7FODSEJlxj
yVOyaSiluhu1FFDaGP390K0nBjssQspwsgjlqh+SQqlwQoHviL+HStmwnMJAGbwF
hIvQyvFYMH7h731Wi5nmcvqC5AD7DHUCEub8Faf5yvzJqrp+/uWprSMbPHqNVkOQ
WZveW1zzTsNN/M3dlfGAV/9yeLxAdLFl6ah3NYpWBYlYz+tFPv0WN8wa76HbkN7X
rU7zLPp+U7JJqe50heuqZKmh9INR+Ry7pr8aY7EXwWE+bOlYrV7oZrnduQzbuQYT
RMugE8LsZLg0TEiTSqm3H0mGaDGXCP3Gkj4/8L9Io8UQOpG62GURe66tgxnyIuz4
+4iXSEiSrDRqdo6oZhCrfXDAklxWlMq64gx9O8nLMiylkIpGPzA9iF2BqmN8uT6M
TQe7iFQgUXHN440riw+9L3K44XUkYXNJddprc/ZW+C/6caI7YFvS6Wuyai83d3bK
DirKlbXqfudOk/+ACHLEBkvI5+usjQmEnPsUcQgy9PAYvFPZJYuy5MaEOXGKPzP7
Ipi0x8xnu8wH0KQdeuc7MZj8y1efWgaRgjOzniCk9NKEEqSdcrgBHZAlmZErc6tN
K1WrIPol8g752EsRzUegNyKlmNj64xiHb4mqzG9VhA3E1mF+xMi7axqm/ML9X1nz
zWlsQz1hqcEA3dUPOl0Zkc7PVA1EyJ1oy7M0Mk51lwX65Fsfu3W4bQpQ48TwjaA5
mrPeBycBHZdWbLyRo9IOwTR9R17aOSCOMM0u6AQDTjAd9/YujOTQS2hlb8rhbNFC
qcaGUCLSKSIHTL99OWSl14gHaRPmhTC/qi5g/wV3hInF0dXLnKz/WPOsoOFRCJyN
70F5UUIg3kaSiNHrlkIXIbHB6JeUw5GQ7VtoTR7oLT75vvbGtO8cOIbDkO5i01UW
HlaZPWaSF5KEfvsddbvgFKRw8EHhrnSyfnYT5SVXAZhup94obIOgY38S+Z1k/7xE
2VzjDWAA/02wF8BlnZcnfaQqXOWzKoEIwHEpc96h0n7RENyJn3sHgiXhXzEk2uEu
vXkUyT/DsYHoJsnvrWxGzp7/4UY1z8xz696wrQ57e68/oaWIldbTZte23wkBfHL4
m7PPoCE7Hurryk1EuhNWKUBL5DdRD0iBq4MLLnwGaZ9B4GnD11txbpfsBP8K15kN
XcTbeuQAJgTXCp2AxL045bKjo89E2dXlD+odWjmHqyZYQYpIAKNv28hOF6K9VHxA
x2+9JLxOKps8bY4vEQMZRmd7aOoxS3OmEbIHnH5BaUtpgm+D+KiZ2uOiO4x0Z+eD
pphRTVTqR4g2ZcDFM6Bi6mWvCME/qteFyk8CSj3GED2jVx5wdVMQCIsWsARfcYTl
uTOGKRL7AIn+KZtwM69A0wMr+XqLj25CvpXWjy3hXwH2CC0au/wmEcd0DkpD8Bco
amtMYp0PnKJSuFWC+3A7plFYHulKoA9NqkeU2umOJ3nGz3DfbjZ+0IZf0Fez3X0C
F6nh9vd9tPxRTEMWTf3ycKsoQELIEBlhMlBvJ8f3gus2iohHAHrQK9+zI3LsKCmx
CgknV5tG3XMdZIYVvw45ZXQrVWNarsdqvo9bS2EAnUMKkc30KcwsDlQFRwgx8lYc
9QDYS59qnF74hQeqtbCyxUR3mSg+H/iVy1FRAuqA+tqIowhYqvRHCJyUfHJQjT4B
ux1LKmEvRc4wjTUtw8oobFPJH7vtgcDOsPXxs9K+SYtqdzeOkPg6eqe7LxOcX/kH
EZ5D2DGnAG4nfJe1y+U17jwOhicqCWIt8e6Cf0B77kCbZRKYzlJ+OT6ZlEs3Zi/o
uKdzua1IOJ3exUh/Ws++yhX3sfzgqeTyYL1NCl7mydfC9c4OxxCRIRoXFr8hP1mr
GOtCPfUQTMUk58M+s/qB9ka7unwzMNSVA2LBsOd4mLLbCd7zLWMdIpB3mj5GTOxJ
tiUfxXPonXhiJsIjBw7UrpoxnZdgLriOSx/M2WfgZH8XjkYKv4Nn3yeqtdn+aUnw
Cg4dNcXxKdeNXjaRKx/AaYgDTEofhyJwOlQjEYLAEsCWGHc+MyLqd3X2pZI5Yeu/
BpuEX143++8Jbq4/kQjA3g8mXEK1wQCLuRKMaS55i3AXMqSntG2n+8g+MdD7lIEe
qm/TcgrOERCTeHNw9DLz8fXMr0tDirHGMpbCoH+u5DqTAd0WvUYb8oY9gDdtfwaK
S9PfefHdEFvs8auFJvTa8OFi/anAuvrOrvdR97zRC5EN2pITLRonWobmqndmXoOo
dQ2rgKMuu7QM9d+cm0ZEZHvIHtfwfwj5I5YhYdMgxUdVmgSut3AOcHLIihjK5Qs+
rYQeRMjU9WXodHLmQ1rB2khtGb3fw4M7/97pda1m7EGIQJzyBCAVGuFMf6TYfoLW
TEz4uSekK0VuoqiCGbOYfOvO4RQF0Pmy0S6vhfFfAzsbLrCPGEZ5YK0yJo/IjUdN
EPiqTk4rhaWDhSE8Azy3u8gcuTo8g8EssUrhXkCROhhDVTHLpHqritYKidBer7L1
5yo9qA43BZi6DbtDxXQhEFrjPt5nCzhwjJeZMenU9v4icvGcYJSf6AJ3sn6W0l3U
tFQrt3fIpbQmlPAQl8s0AoI2nWAshTmW3wRyiGOS3Hnwt1XGvU2g9yEwgme7SSiS
A+wBaelWq6PtO3ZrPSqvTH99KUVYfJHLnx9fDh4tAA2ZcVy5RDw8mkGHLuOsRJXJ
w8jiAGukfwSoEbNUCTTOqCtutu6FPC1pJoV+0tQi/43SYB3J3COncjoNpUXOjdoh
wuFDtY8YmcO7OK7Fg7QMZEtDvybtm7WymZXw0aOZmeOU/yZH3kRqJsro3i0w+4of
JQmkpfw77QBx7ieYJVSUo6NL/Kzy7NLFX2ZHlEdibhiy3VpeMWrXmehFUxmFH5B2
9xNe2JxHLpHErxjNW1I8DK+4FJuzEoDp87wPR7q3VgFu48feVeFTbfvFC9a7IEjk
7ISaDgTXhAULw2+fRmHDN9/oE3FEb25g/xyPLg6vZTA77leH8g8t/+RqyDDzH6oU
EaJO8TvfcCdnX41wQV4p6L1NV6fopa9hod8G387MbxNBnpM6oMNDPalW6gI2Yudq
dmHROTQ29sO/52ZL8aEd2EB+8gHIWwyELtrVagZ3Vzh0DKx1w5JHSbbg48/KL0VI
vShqpNLD4NSJvLFtkB5ZHiHnUkKsgR2Iucb9r09ncm45jlRAV95w7pydPjjpAdyT
NXasa7ITX111gQVRHrGJVMo9g1/w1DcGgCdpVaPuT8Bz0FYz3D/jDzINWCWFKUBw
q7AckT7L0VXsVirzpm20kbTBxmijLkQWbMFZ5Op3e0ce6nDDYvqWp/KzifoEZAli
qnJOZY1IVy0NdACje/o7fSSfy4sZN7KucGIpB6Dk0UVGin9/1/YhXgJwXQXv7hr6
4R16dDKIJofRCwZI2KdNPdDdAZMRdprchiHwgab77/mo1PNpBL1qyhXo1OCfDZuR
kOu/RQl7COcZP6kmS5ATvDGeO/LgleemyWOcEkzU6bRtxcTldRYMVNGMbkWSScPD
+jaMu/dphi6EYZUHVBPveiFQWRgSvMXPEGKF1jrKOEz0+AmL1TDtluWonVrvRxDb
AJzL7Hg865LI9b/4QXk7b8hGGAR8L6KXq2POHJhUXqB1KosD3ZhWa/pu9GDlFeq5
ciewKP/GWg4IzA4C/UoWm5vRhCTgPyojhcfBOA8xXspY83TZAn/kJi5+w71I0Tx1
O1qfNgptKyXsPuH9x3IsFb6s6Lhx+ghVcnOSh9lPKG446GzydM5k6Ttu/Y0YgkPw
y/fdxLhstty5pY4Bteez3TWXIK5h8+lO7IRsCWse2UPfCKIu+fHbO8+M1lCXFfDk
XtbXpUxn1nvxs/TzqWuHmRv+A1VXFRfPtEC17LN1dZN0ShpWJ5rCPck6JHvcwOSo
cOTsoIGaBSSklwhIX7qJiPriBVo4JyIMSe8AO6z8SwnLOtitmySOrZmLm971JvH9
DeTBoU84iSj1QrEy1DfxOO7lHP8lwsh0tF3dN8gEBRJwNI7/lpbK8GkIaEwIErBh
0D5okisA0m97a4I2HXO/oTRCphpKAXhpqtPcgO3rCMU5DfZ6ox0dE3n0BiG4lzKf
Bi/w4V89g6GrVoDbszf6aapAen3R5SNJNlptBwiAMtlHUSPgZ72vu0XxwL/wSCrY
8yEGCaJd7Y9P7VwDpBP3pgNwACqi25M1oOLPXs/cRbxi5ZL6d0/2B6WjAoMc7D0k
Gs5bn3wJqSoKEbWCmSpUrCtMgQPbhcsDnf/kxJQobKZPb0Iwk/MwaZCo5rGs/GQy
68O5/T1BkZC7Q9vogD6nJQzLOqXkDq3s1JUFIwYOhYLgeoDBqaTHLUbPqTs2AKYy
47AbYtWQg8PvP7unfKarrnGQh+eWzCw50vLS1pu3P39tAEtcPueQsjAJwqMFjEEC
eav81gjRs/rD0Oa6pKymq5u7KWi5rz07V0koBruzk1YBUK8KVGh/RNiyny1x7eC3
/Tr5O5Zdl/Vd012jMKyuSlhVNqwUvS7EOAPqrWiqDM74dAZ9Anh7wE5oiEhqQXgY
E+Phi7SE8F8wxoKK1ykKN40ire6bDrR8eFWaDprbOIY7PbS+KTotjpiyitXUGufI
9TxNVmAv+ISVdgzCs2jXXL4pECuf4eoAzAxD2lgjLplA6YDUk4rMzbKTcZ8EWMty
koH+StqP0QBslvWb0KjfCEPIXrTbynft0WLQ8FjYHqbuV/YMYFZj10dph/TUhQ4p
gZXz944Ishgg8zeUzrQn7cyFjWSLNvum1P6x0l/PASFDdm8CBrAYdKFYSAzXxYoR
2YcmoLjbpir1t6+Q4mCLXuPtcr7RZE/Ga97J8OBxWcjYSdD3C8yUE5GGBZN8PVCP
n0tJRgIDwN2M3GQrfVxrN7vsq75TR/z9HJ1QAltmo6KE52BXreEqLaOCXPKN8UzL
9MuEqhzlB002r138gz0l820elW6MFLjx7uOzcnNyvOQnsA3ckQBVaKTjwFMsWfvq
wTVIlXGs/W60FqKGAP/1wWofxWUCem5IucZduZzTfc5PIZdsb2IZw86ySHVFRHNz
sRrh+COjqlJLNg7uTvtfJONPWvHS1EXjHkWsyHOwEHnfxMZZJV2sBf9PVYBfPemq
wEQbiclQMn1fUU92VN8OTbtHZnVjH4rcX6KwMoXwg70es3Oxzal1hwFyuovY5uDG
qGGwN8jDHknTEFWD25lwPpkkDDUXGGCmS9gqJ4/PPS2JB18dlCZ28ikuuxNOVj7s
asbk3SxSSNB6+Ex5M2aMqnldmx3s/aoh1NHvzOXC548EW2a/FA9n9fjh9CCp4rAR
WGRAQyNxcpzYg4lR9KyGp7d1aarTZXvMIcPtZEkqs/wihFoz6vyiHXP0OGJk3geY
IGVrPlVXr5on7lZ79Fz3wTTJw7P34T1aCwWm3dufNWtbkNRZyIQZkpqFOydt2U4O
53MQ/dr+a7Q3h9D+qWBuwIow/RsJHUGOc0buSrEWkAzexLnKb3xrd0iHykHKj5Fk
N0Mf2J4WKSU8dZm9dus/hQVX9bYNEe2mhgCUSiUZUqsjkDX+fWUM2RL7GtJlIy6Z
LMrxXwgN6r2J92yP0MVMP1PlqUZjN6zH/QzmVjzLY918RWRHTfOkak4Kf/kgsMdY
Bv6ziY/CDjmZ4n9ey3x6Kxjo3E2CdJnb8pBt/8D+6V0ECw/oWXJLxlyNyk12Lt26
0K/w8lkyIqQ0/02YGgQz8WZsxJ7CYRkBkAgzcapLfVQfn+jgxS4CqbBjADxYrAvr
CuM2rRJh2ysZiubknIsKyoksHSI/5sZ8dDOPeHLy/i7MFDAH34z+6ERrN/3otUKJ
RO9UzQ/KnQKbgJlK4LoSTZuz5x2O55aI1AGj+q9Uf/dQjzAZRhy2mqCIDQBK8Cdr
0kwtK2Jcv+eA3lMOzrWWGIKQhQcTaRQB0C1YZy9mBuyiuNrWpaImKMJgWPgprd73
G3PrHy4DB4SGOoH83WFdTp346tlL24tPYwFxTkMPJ55psGeo9UsFCyn25aCYg17d
REDwJj+hmK8rabLMn9q3vwjnnMT0PnCyaoztg/XaQJh8cDCh/jDzKYIER6yrBwCK
RvHb4GD0SM7TxVyRf9tP9bwe0rsidK97EN0U68HTqP5Di7lDwX5iAjIlDk70cO3w
6onNfmk8Ly3DrIKGTO6wQwb2zLXNjF8SUF4osng8W2Go9yrF4Ph664UCzHIPxKTy
djwOZp/ZhJtPRJsrpxbuZYlqtC+sEchsj3H+lQRLH0aDr8KvDjKd0G3MI41wX77W
cJhnV4CSJOpYaUfHorln46LdzlqBZiT1IMCFTN8rORlv6QUD/bqri1zqxdt3qxQo
9fMqwytSZFbTWR0xjrVAE/cxKaDLGL8xREde5CVPmXV4RVpj7QmSAtMs87y63j3u
FwfgWPsVRsjZKi3X/mnKjtUrQrtHeXoC53tcSMyCJMxZeSvgkuLRGx+iEKWUmbyy
ZwjGSr0dLt+FHmSkqyIUb2xIXko8wmaGmHYKJhk7jfvNMqsLCXmqEnIFTwmyd+sh
MmFZTuZExzGMeixp80PZsGJWm2gO8tgPH4Is8cnqo3wq2ZkoBJ9c0n+gRpvwe8sV
rncXWx6l6t3VAhwK6baC4YJxcEJjdzdKs5yAjPumi0pxJVy4KSLpKqexSYP7DQQ1
StNKqLHCAoZePsKJJnfSkUkn11LX4k1Bkzk/joAebhB3ZHHmRT8L2f84CV+INnRI
F4ToT8RwsKVZZhOPqeLcGcKW6a1PlbqqjjGtC86bUPV3y+XzooC1/jU7+GH5nneV
35Uly5pG8MguLaKLYkFGzPh8gyzA2wa4g/DzyaP+b+opUQqbRUR/6zVclLbnaGfE
652J04/LSWFHK/XvWKC7mUZFck9cBSDdV/YVY6hK747ZmOHBzPafQ7mTNNVnc3Y8
Yo81cYlPNx2G1BYkoH2u7eQRxtHAlHGI3/jqDS5op6d+nRWMZ7txM8Yd0uVhLJxk
8R8gdP49wmUfIP9KPAkcFJlfWcIC5kMO6S23vurPQ2UoT/8PObhPa8Rf/9YvVHwW
JLqCUkHtXFy8W/rx/LWKsTQEHiv62adYKUsMHSBI1n6L4ALbvAzYyqT04KRk1CJH
oFkAzo4Jfl2itpARvxOk233BDBBgKq2MwWBZMrIaXl2E6tCE6hGpuBFskQ9wLN69
+DVmhYCJKY20TzehceQYPyamY0BgQyugkyMpSsMnR+fnt5caaVgvBRj4pnVmwEar
blp+7SVqn2x1lc2PGyeAoZ/uxval0GJJT7yydd6Sz2XMhOS2eEIrj3tV9eUMOuas
/k9eiQB7vU8GsuY03lAnphMwzlGfYh1mEWRzErh3EPwqCK+zWKWWt/jZhD+Bi3Hw
U4fyvY8jJ5XQoF61y3xCULC8tEU+2/cdB5zjj5Eg7Ugkv//Vf77CPO6FPylRlnPC
72WHdcA4rBNigvX/a4pNYiUp5gd/YKoQ6kKvuDwy6ER+Pp7GTIVtVz+KI35yIDdr
TxKgXm7UYQbcNSYFh4u2YdOKzTqmjIDCa0fAhzMReH3aR6iqu+n323dGhvJmOHtn
7DJrK4Ly2WZxDfaDnGs7wQswtJRqWqfIwrGwbFwfplkN8WdluI0ZiNsvt5d6aUX8
n79fAnD5Ni38vuS4OnaNJZtOvmNrD6hd0rCDovJrXM3qmaY+TdqTx4KAQ2gHdwc2
ce9xoqss2twx5tE4qGTd0OYeL3Z9SzsnTJ8iY80EUxJTaL5CaqUgQa7ByWmLhRRp
Y9fldiFnrQkc3l1Ec71ZaCoMgmfPmGVcAiz07kJNTZMqHLLjwQUO3q4hM07L3+oa
zHz0R+XNlVz9Ys8j3GN/yJB19EkdkpEPX/C+okqVZ+4YaQoIpHZFwFTyE+1/UkpN
fLC2Nep6OgAimiQyl4+WIwE79bovFY4SRZm1dgFRv/g8jBNx18EkjQh6JGlfWtmQ
fvV2NSm80Z31OYlxEVi18eveFxZurE54YCdYgIGey2rXyPuQBbOGjPU2XhNfZF2D
prJukZXUSo0Y+mIfQoRW+uN5+L0DqCLiOstvOH7wEs340Nlq93PrIevnpJjMAHZZ
e90F70tEAX9nr8eKC+wLoCxngEtlR6UlBhVwT4gDKh24z/Ykyt4aQ9rBi6qViqi6
TDT6IabKwFwLP4K+CqpGiZOc5UQ4H2ox+Hm0+xBioiix4zc1ECVnDL0eF+8PxGYN
6C7PG5Q/gFvP7/OC+QCz4zK1F8LKIplN1FJoNeA1qsghIBPRezNn1syshhW5Jyf9
ksw/NiXSYXlw8Xw9qND1LX0WSYCENoBUDCfywajDdZhN9BcHVnCuLOwJUJ4f9Inc
CM0SERD4BDr567DDURKWzVPkHogLfoBnYu8Ddbn++7jZlhbQr2JGidbA2PbZ90kI
BwRF4Y7DQ99F5M2hymzfN4hMfqyKRtQlaikGG+57X6Jqy/t0znLbLI1OqnpV2N7o
bpeZ8soH+9oZ6dWO8cLLvIgcSDmLz4ngwH4s6pZtkdbMLu36D1d/djro2mew0qP5
J2+zeOpALyvonqJwipsBjHJ5tUmdFzLnIayJIxlQg0NqTA7rJdQC+TOldj/8mPCy
1hygvXQ11OWvSP1iSDkuKyCa7Zs8QWD272Qbl+LAxiBLk01I4IX0BVin/XT9S2TD
fSlUbdHjm/S7V42pyrNhZz4bvnvlU/bN6tx1qt0e16uzyTr9j4CELOHaXALQVSpd
pcb2Qwptloc05Srbmx/2lvu+EetLNi1+m4482Uee/YRC61GgpUgHvnjMrptnCaSA
ZqddadcuIwBnNa0DB+RjdLWmE8kImRGEs4UNEtuTYrnMF+GK+dJt55DghZNmDHmL
jpzR8bm1X9CPvj68rk5hdKRsJjlNRHV8phD0ai+ItD1HdBPBPfoi7a5d85sA5bT7
uETQssjUe/621EuUnIsBR9P35/O0odKk6vlWsXNmj3UbrL1om3bp819XW86/NVs8
8449qH/5ZPtaMedO6BPu7tSExwvrIWeMMo5B32Ze0MG4aBVmICNeAO58Elt6dbkd
RObRB8uzyGNgIWlUGYGMEmHJxKvYq4u2pxf/bXblIzUb9qqB1iqBWLpg10s/iPSE
bKJEquMlKtfi93s1UTipnMZnpxd2z704IUFk/srX2fcP7f0diE5yS4x+Wp0zwYZo
GYUpSz1qBIiyhLeLI3uXwsl7MN0H5L32qWXEyqWBTzoOgsuxq4aYtUHjLw+qFxI/
WhQekdjlxwXbOt3a3yGkPV3pSkc1cx56BEzklJqOcs7NaHKW4rA7PLV+ZiB9LiUB
hrlPUnXlr4kwbKQaU8TPnYWYkTFVtDBp1JTaOnf1Q0teAddGqVypcRz512rLGaMR
XoDxzDu4HdzGg7DhvPeA+cqRk8hTKOXzKWa8JsXC7LPrqIumhOD+jlv9XhQ35SE5
k2PItgvlJKvOEI7Dy9nzWBRGftphHp3tsB/nXEXaKEMCsZI4ZuoaSXOR72GQj53b
bZGVjFa1ic8yHYvFNnRShSIObarUxRHMlkPjliYRZZ4hV+BQq0LzASkeutoHx5cT
J5AOiLfwssUaciEqVRToKuXCHQalcTqUoefzMOnMz8L0mXxA4pR+2vNyGRfl9XYr
D1V03DitPCPT9KFcP0k0xEOjDCkIXyC95RJ3KMFuMv/ZU+MTL7Q3YDhpggkFaGYb
85LlSJ8KGK4kdyrY/NRKNSMlQ4a+glopkDC1Rrp/hDmngMIgyAdakgV9UoEsf8BX
rpwp27nQnIPuvgWPYq1gue2Joe6GAo92341k4nT671VUVAkULJAFlgOflJ+0ywta
zBZ9flFILAZFJ3n2n46bFloXeU8js/N2GafhZoUTOmO9tBmTfzLmLLEzU8JEN/X8
8Z4x5b9srKvFXJKEiRrJFUQXKxxVbo1yp8SLlLz91C3PpV2q1rNVdrAqrfMqNSEr
rRfjcomwBDwfPprA7+AOP3swUn+ATn2U+NmEaxZU9UC0wI3WUNsjaLgwleAHCvRG
avSDO/9GFyC+miT0unlnUPzLZjVzm/YC4dZG7W3LvJbB6tR5b/ZgxwE57l1yjoTG
cLrU+VhG0C3IMPkuU1g+8Brqi06aZPixEHSrmREFffnvE4rS2O37FNNqoyXemGxD
HPdPnlkcHvUWV6SIvPk9Rz9VdylXftBqr6FcfiuEE5lGbfUUdJa5RBRiENPn9mOV
h/d+W+cwPWyYhDK5SAvRu3618q5Cfq4+Y9VEvsiabfespLGEUBGyKDRISCDqv6uO
WGDiSd+KbJx/eydmtcjTTcy63FNVpBG0wxDmP+koXT6vsQqMoAIq/6LDMX3tuy37
d+JsNqh0qTxgQ97xGuI1u/2hPxdEllGVPSkeEHvajsr2j+nQvl/Zh0l8zjxxmxjL
8j0r7XbsqZ8HtDSnCvoIOSl29cfF9ij7WP3i7678ttT5lr8iJtvWS2CrmE22vVBW
pvMl+RbjNBY3rqvfboHuLm3y+H1cWQrJu0EiMEPV7Vk6LxKQMtE3o7tXHVcToTTl
vLYohBrEutcAmwV9cL8+tJn831c1KnJzvUTzncB+8XH1z0lNgWFu8uJLmhpTgNus
SpwPEhdoxJ3hJjYD5M/oLLPhNy0uj+sgoztXvqNZ9NxX+U0v+fcCziHp4VLt+I8o
y2ljIn+DFl+j+SB4QKukcquqMoxyeKRvLHspLP68ArKoRlHHvTDcgM+EfEkl8j5f
7Oyrj0diegNmY32scbEeWu4nWKc4e+a53flPw0i6S+1TQ7QElBUgzzbsxOPUbdI8
1uUZS5TfEyJc3gLgn/Rx+AhEdeyc3DfMSpgR/vG5sOeEVU09Su0bTu0OZZMfRMb5
7w5d2AkOBbuzqaHFzkyE2U2f4l1I3fu1LSWrSVS9b/WQ99eBOuJn+chCHVBF0aKx
sWWKxxzD8EQ63JzOMfrRMA13vE/bFLqjKeIPluLSSq0pYNXsWE5ZbGQqmo18O/oq
CFaOxLjtt/RJG4TbZOLrXdjUPPRHGYp+Fw27v+DfGXmu8ZB1P2nk14zg+3f+HiuE
rKmf0LkNUPiR+DsFSRlZI514EeaeV79j2g0wPCprR6X1DxqXOThEVxEbb7BolNDO
H1fvYeNNstJAqG4mdEUUjya+Eqc5o2AWIFEd0s5xjYmxZofXUHZVSZZj54k0sQn1
oJxvMAahMpPs6MfRMKQoavKNU5DbKxc/EJblP1uBQRddlq6kgB+GL/SKxPXNGC09
O4ppWGadcNQK2DdZ/W2EfKNEiwgGm/WujRStlDQ5dzAMZyb8p5cGeh7X7kKg+w0c
n89bmk340uA0EGzj40VFfqu0i/PWLSEtizOjIndBt8zcpRH0V4koBWMYqF8mNPRV
E9kpJKzFcWEhLnItd0zr2U91GIRXAngsHuXFxbBDD8Q9UvpO5l34J+mDGLBurTfT
6Zn8Eq0juq1XfsIUfvMAg8qe1uR57qbqXZlTX4238I+I/EDuedjbvvhytWV1+cER
j2iAu/+ybfwTRHqyowARAd1XSGden2uZoXcitJnQL/ibg9GYiwsvmYQzHGAzPJjm
A+YNPnnF5MdIKnUyTqm/POJ/prQZZYyMW9zIIYqeG04cDuQDJMLaua6WDj0fqtQP
GjIg7dEVIbjqiRmeqr80Wn5mHI9jqHx4WBa81viuqfzh8gwgnOhrcEPjHxO0umMj
B+JY3eNZjjfa2wDk1PBhwwbdaqw7uNlj6+0XdHoYzIiHhaJ3j1LjsfX9d0QYqT25
IXVwWCSu4e+osI2ydjjwpsJEqeBsU6jijcl70UPKkPcbBrW6uT3/loz/w3fl03n5
BKc/+nPfz8YGew5pWyAKJSDwq8mIfz5ta5bdc68a7EhybXn1hZNLIrNzg01RrO5e
tf4sTU86Ezq1MWDhRvr7cfUssoUKukpCoOZ6qXgGxdQbc7lMXST3I2+wgW/m389Y
0+gVHj1bW4ghHUJtVlNE91Tg1965Q1Sa8zvVY7WxvDov/vwlvUbAKFU9DTWARowv
1yz68ydQce2CQ+AkygM0OxpIdhrE4qxUeEJAOs/T7zg4bYouF6qX6/HdXqVbh5HP
a3ye+EgXZihPgsOJpU7o62yYj1bYDuKWcnNLZ2iEeeuqenloVhEmNwwWGXZzoWMN
18oPCmiHvx571c36WgJ9atsPEbLjXrTk/4mQYWEgy321/5ZE6im3Tx6z8K6S//Js
S0OPzRlZdPCL58OnujjGDB49+8JDDB0BOxZSFZCAM9YKGRJxOxP3+AHQ31agn+ru
mZkJF/1MwFd6/lWieKKBOVET6ZGlkhnNx5yKotriS1R6n5pWv5nE0T1nkYC+RgVE
/Y1SjNbYj+jZuIm9zUSSUBNoHrE6cwbHZMvtHUlQDaZOoxhzeFKcsEwn8jFmB20f
BotlAaTAQFBTRvdXIxdYuMHclu9ghpdIeOi1VD203dokJnZ7Mb//k9ohSkRAAKXh
w3THQb//f3KcvRRffG2RYHvhwd9KUOK7dIG89A0J5W2Xnwzu42cDsOoLjNMARmQZ
cZNE/IxQivKJeKfH1rCnJp/6QMUVNYNPk1S8Ed1//JsuOjP21tBnhJPj2M3kGNvU
qx1wh8w4+n80w5Q8CqBmwOJOvGiVmNX+dsOmps6dU+3uwBF2S1DYDZ+UIfQ3uPj8
iVAJ5EesLWclJ+wSbozUP8ElfLViUlAEDZ09FUoYmDz+FdKGCEpQXTrAZDFtA6eu
eOseLRg4c9Ifugf8d8RSE1WRL6MRcqnl0y67zbf70SF8pxBWfkAW3iUJgqIsEECl
veYHebpOr6c3FbKWcyQDNDxTiJ/jBbA6O0t4vccGBR3UcD7wUsqZExlTA5V5aNvN
o9VYDfZXdujc5HlGQO4req/GHlSoK4VxJTwik6tJ8EmQNSKfefajhkmSae9IymWK
19/PXpaWAYAUVzDVCWYitczl3MkQIUzP7mXSSLrH5tmyzsTxMpouK7st9thGj4M6
QITwdBRPKODq85yd/trG2M0MPdjyP060MnHj08WieQRFbvSAifBI7GKQZ+UGPE5t
fhWX8UB/pfvGG7J8u9g7nXvja60WPgEId1YZNKo2wN/1wWKySiB5wbCIUPfy7KPC
nvK+Bf8nedmnGBFGROSi8r3KPH0CCEetrHDqYP1R2p5KE2E+GnTx3UnV6+8ABN5r
RJmTV+PFsDNECACngUFYlCO4LUP6uGMkm0InWkQgOMOms6OaFLU9TXcUkkysJ+nR
l5axVhCmf741pGMyDtvlJG7wGW8y8cXNV26imCP7CUtkPtyn6GmS49v8YE+IlYZX
yauWrfUG7RaJo5UALKHcaOX0tbA3gw2jJcON/CRAgvN+mZCzphjlUuimlNS5XKTa
Q49D9c7wsCgNnSZSYeoTfZ8b0/SG+gtDK7u2Nzcsh92ju5Oc/mBcT16L0BvZCcOG
7PwqEt5ct9F9bHoIgIWNfdOAOg9oNWrId4z9DK+s+BdyydcjVkQdu+iIR+NDlbIr
lZkxguUEUxWCUXRlBLFvs70BwEt9b4nSwahZIGHKbFPUv62Id8RZ/wiiHU0JGRtS
A3fbhLHKYdRefos22rJZRGAFMEIXxTgSAEXb0NzroeU7m1k72coHUkCEMxH94Zrb
JjhTTy3Tjutu8A7K1nSAYK0ms3qXgesS624MWD4IgZQCPEVPgPxPFNhDmCwg1Te0
emx6kDZn3Nd/uokC8rm3gDciLD6FN2DurWVWFt8KpMf0mgj6v5T1mUgstLxAmFRf
+2IX4Ee/F7rokiDuf3VAyMPkrU16kZUbFxWaUaXiSm9oc2okuhta1gqeLPeRM7od
/8O8VQHv46gqpOnVeBSYoaDlhCYZ0pDu+cXJ3scvAqPVMwF62vVCjk2jfROpNv/g
wabq8IhdWO57qgNCYg+Sc5MyHaQgN5chMXY8/Kds56R8OCRhGreW2dA7FVQmwiR8
xQ+EFrnEnyj/JXqYTtWztt5kOnmtanlz7MClpy78RyEYhqWLPyU6z8FDSXHsBimY
xD5x7jBcSoWb+eyy4F/DeZt/IKgWU5CncNMyW8v6z//rP3XtcCesk4C5ym11bsfh
/2rJhfb21fRNXpYd1y2uPtmIlnYaiNiDvgeouSFr7PyQ9BRkMJ8ow3LIG2ZW3dMA
s84VreeV/op1qySHBqXe6VamDPGDHlw8SBswm5te9rtFLSkPf7MqJlnbi4tIMgwu
MSzsgA3I3Iwdf08iVX6MVlLSoVm1rA5HEqjFQDLd0/KcKYJHI9fOjjJu1fp1cZPp
X1OnliJpGZtWg1yzytVJKAlr/OfBfQVXkru3cYSu0AIWT3xAT05T6trgP3RTfv+9
xj9vFuefuD4VvgBBtWL+W/RqmzNCV1Thurw2tT0y+7ct9N05McX8Ib0LPgMjw1ps
flmDmAXkMVjPWdmsF2Ty4TaXOD8a2xagS/Ca9gyFDrdRp7FW4il4GxnJQWlsRzJs
Vz32GR1wy8oMwai1eF3hDLSDy/5NvZs4RtnjIDWVZdHY/8hR5RBArqJA2H/ZgNEo
cTPjbO/sweNPLW1mwC0bx4V+QlvOdmQXpZgBYz11WD6Z+R5yR+NZCqUPBGrsZUoF
0m8MtKNuqM9f63W2GqgGR1PMnsDRU+YpVs4oF3zvuSPBqOTd9Sorlmq69bziMetr
OTo5limcL0ANs9TtXsbeaNjaZrXRdVNAnQDo1Psu5x76nc+VwkFMEi/Z7merK+kg
T5TAwpIpYQLkW6xso+hoOGERx4eTSEDUR55WWUsRmWGypVwySZSmFTeZneA49hJy
iO7NcYlPhItnR/zc1E2rvJLsVPzSI6CfiteuOpOQ/pYZvEn80UW9l2bAJvJ/PiEY
Kx9ZCMJuIRCIq3s4UUXgxKuxiiJ5q+o+7m+fDU13suJudCZYU/CR7Njrcu9TiIw3
7e0ZFZ6oAmP9O37eZko3Hig/rHYD+C7Qt3mUTuWqeg0IbK0K/CAxxaGGSjt2aJyF
0Lb22TophLn0mG0dOjay4Wva85NmjdxIzbBE8+UELBU+DI61iGza+oRNNQjrigiV
sEzOafBoR0vwf4uYD13vejdLfb8HAKkipsc2rxmJS7Ub9RedPTxZKC2nY663QUoQ
/voSpli3Rmbp0HYp5S49xPeAIsZ52yssJoTXAVSR5U3Q7PjLMxxn5vBk+p24ZBP3
eaDyOk71UMv9s6hPm1U+OcLSj0W3yA94NHbHPyU4MhCaNdXR0hpRMXQwQcuSrefd
k/BTidF+SGruCfOtJS6S0KNBoMJ8a8oKZtdg32skaAWzBqtOsBm0h9HmR7Sy2qgs
tUe97gLhWfz7Kl2/F1wzjPbOu1WuWgr4r/FcfXwBtji/OWXYmFClkCNA9g115NRJ
f9C/NeKrllIhtPhzU4dR4/NzC1jLUpAChLtZsMKZz7hMEFSlNGoRA72wRTA359/8
2i8qeMc4H2U4eLxCgQm/nrjnRwgFVVLRuSpudMjFUa//pRFtyWFsqyF3Uk3om48S
z5BJ061tfIYdRU16ymiS3z+kXWyspVUg8XKwjIi1/xSBZ1buDoLHzuEOk2QpK/A/
vPqJVfyhAFG+Y3sw/EkjQPAdUoZo+9TLwrPiGBL4d1FQK6jD0eFbUHihh6QZ3dU6
VWEkq0rsGxb3XIeJCLqdI3ksIUze91ioEkVWVD3N5/19XnApsSSEqzQRtnOzvN5I
hKe0uQ//jCpbW2pEVQLDxvJ1gN1kNLRdoAk+5zx9MbC1xZIMoWYhKO3PrpIA1rwx
kFZ/BoV2uDAZg9WPSYvTDzY81oVy49jZZ5H8a7PMd3a3D1T07DTJZARhEsZtbOJI
NYVtnNPoxYhQImzDvpIB/B72vSXv1trSjef/VJhB3dycWo7nqcY+EOPAA1DUuBI+
a1kh+32WwcYKQpvogMnb9+o3Gj+5BuVT3khOWskNwUprgBoZX9JilMihZAnh+EPH
jhClJHOKqd3N7xdsLzsARxAns5ZUkcAci9G07fagrT2lvyZbab9DSoxDvtEYLfaS
Qz5U7uP3ib+YFOF6TrvGW+cteOVxC3XMRu1wfKT3N6YNVWiBuLLDKhk2AQ7A8xnz
Fm5mumHN1VQU4ClhAsW2uc0IpBpaNZiYqwCS37NIlFLbpVtd53S7JwHwHno6Qq6c
1cqaLF8I395V5fCiCmVk4izi1wo8nyQTENy0WfAlt+SAbNaQjSfDCJ9VNeQ6Fp6r
7FLdi6Gb2PtbUY1Uyx7LFsCWlAOCh6uUiEOUqQbVxErNYDK1QqIiqme/C1MjBK+D
mTufixgHE0EOSGkEkPx8jfPVI+XdiXtI+hzMfyJtHy3f1s4ILIhylCIND7UCZrZz
sXlx127yMTL0Din2xjU107xV7buCkSd6UthOIMraRg/H1frZg4mnOhOsOcWn+k2s
zkjeWtYgqyGolOn4/k8VR7uyiXzaiyUH9yi+q6HaA4wg0662r3KWEqSfCOZqvulU
ly7xubdTnE1qifizM03LwruOWsLSGLU7fvXYCldYTo6f2HjhVLMd714opYVrNk6d
SC3qU3Tm86DfyGi1ICFkJ9th0HtzRiCRD4KU6FS1Sou/yEDm6+iuWV/k4V64hMSS
8ys2wH+duozC2qFAYt8UKXYl+9a/q5sZydsGY9jYEVttbRlWwlcIPZFfxAF8TH+B
6PBPaJNeIqXENBgfjwkiLUX7KvCyKZ61t+uEbWFmv9ubXEV9BvhFJ9dPbSNi4n5H
bWYZHC6gZe2MG3d0YdmTQSN2qTQFP/b7EKqyKKTtnJNHgi0g+rA0YlRtXkC/Ai5j
VPCiOmPtgjxn/z3Lj+T0nbGa3Qhtx2i7iKOycMsbchjLRrn9N4xtJpdaV3tYJD4/
xbOXy2qm9lwvsXxgfYWybLKDKISK8XF2BIXZ22sZxP5nGyaGPRXQ+utUaI4t9dTy
MOx/cw/CCD/H0JZyVQigc1iZXBT84mHqPIzY+m17R3SsXQQ0Y9v/a6mAwZkYngGY
eGPQyFjOydqTS4pJc4ArMpMjrMjaJYpAES2l/hYlXMa0RCjDqWBddv1ZYJDF5yQ+
c+W0MWF6dQ9FZfarAfXg9DEJm3CQbC2MYxUItkfWAm/zcpvPY7Uyb/zOJDqEnRUR
Ns54ML07k5aiYnOQh4NxqsNXY1Dyrt/8C9wFxznBtScWTiD3V0wEf7wjwex1TjiQ
HdEJvy1cmsZa/zsXu7fJIYioHa9GCQm0RF7Oa5ULJIIn2db08cW8OPfIveHekJhm
3jifPNDpsnJ8YJYqldAA0FvPow4rr5EWe8HFEaIzv5fQVD0Ugg27o2LYb+V3FjSz
WkdxXeDcK5lwUVSbuaaiCUGNzmwP3Xk3ZjgerArgUPdV9bCJ1geanXjfQUp16nfb
EMsHFTYQLDFiBm8Uu5FFyKzmEXDq99BpQNFYXJF8pIWX1dUzwWgRcdsbSZr/4Qqk
5QtA8857L2f92wOgjdMjBLUtmD/RPHj/wuERqlJv06AQW9fcWYb7lqrMjdnvuUEx
3TQGUW+I9Qmt4TmL3MNPdoiA6Hl0RwH+guLhhTp0zEhewjNS2puxRuQoyL8vaKr9
9GwV0VinnDIC2qPur/l3hwbKir+b5KddCTc2FccVg9VnWMb9pWAvNV68zNrTSwXq
sw1ALtNcStOgmbT9sMW0LhxHfQ007TVtCKLspY9OlhP95KoKqKzQFqLQFrQeA4d2
CnzOWbe9VeF17pr4a1FQebj63EomeZvsNLeCql/BJPvUnRPgFnLTk08SqvSW/Y94
59MoiQLMWjFz53ToAXbBX4oeCdbvA5dgQVtcoWiQ/0E6I7h4QsYOgmm154xxMh5r
z807bsUteFVytosTUaMEaS8bYseITn/t2zz3zTtUpI4YIgTx4LM14pLPoXaT8xRH
ZS3E3+Ia502CTq4/dfyDFtKmP2zrKZgm2ZKzqtwj46Z14zGt0zq7FhzUt+PfS6hy
BrhIpFIJwXWP731yQuyFdCSrh3ZvTbIyz2QRPx2/dDqfGk8mYHVByB65PBef09iD
UyXFvehByENthBRvfPzpus7SToqfLLXtr+dNaWQiwWYYZQA5B4Pm99UdfCfAjEyF
kFIrgiSA/0qUoV2zc1AyFApFnwCtqfqmvOv7iC5AvvVRnTAvEnAmcKZNEflfv5u/
doQvTiwI8mpynJbiykX9m32OqnRjsjJ/+Ayaeifdn6u5IAsjDcJTvNmhYXOqkQM6
VPqf7NTDRnQWdo5t3YJVK/jR4zVLrO7EFaNCfmQFHOIt+hLJYo8vMoi5o/be6RUz
ikDXgXnMh1o0Xzpl9e/eRlrXqUK4WoksH4MCQkahoeU6vi8sY6AXQIqCOYsFq7Fq
qYvmz/m+eND/uHf9oAFqiFofy1T9bvz0QP488o8VNfTQQyy5OGuueMc2QLoQNf+E
UtWZJiMfaVtUj/el4kBMKdtrjU6Ym+V+yQujVniG3ncOd+X9LfdVB7FECJD8gmwZ
lwNOTs9W2ICy3tBfJtWDE3t0YIEJ24PAHINwKWsO+E9pEZTNqRZScryrIXLTeF8t
HVnwZAihN084xF7+JKWwzMqI5OwoAYNy+OhZMqtCxMyzQ0nTG2gn0YEPIqLgNSu2
aSja7sWY2GU9aNnRXbtXnKG+cQ17Q2dkaYvA2fIHDTYm71pgeEUb2hdswXdmmLkp
7RVepUrOfVMbIUJMye1a6PxG5cmTbGVmbUiR5QLMRVdHuEXvkkUitm31Bkw6qpps
o6Bfil1FW05TNPdrTTZmf9wFQIYqwsLEA142+Vkp/GAQUNhaVhjaQ8Bn2oUAZkdF
iIs4P9p9O+P9LIbpLspIDdPEVBxi3jz76eG2C33dHxQpaGV/XlrWsZ2HShRWNCWt
v2aZTALTlAARyzscvKWviIyZAQoUhPlTQpDZxI843l58XknXkm5rCeCyNn7naizC
+uX+fhUO1aLtMC6q8CNeyz8VY0PByQtrLvtg+NPHtGjw/VyUNaqsYqoF6N8UAM7B
1+dMLsP0Z8/V8S92Vmte74zY/Y4juc5XkVfHPJ4HPg9fJDUvjBsS7jIDklhyfFTT
mYwa/AESBkEECW+1tE5cRy0ztFTU9JYoDol73oMldIKIV/N989hvHU3JCmhKATO4
/SiXDfb4FNyomON6YnIIVYZAgq/WsLxKNJNwgFGxcSjdOPe6E9K9ZIUYapfUq84m
ZJylWnPRcSnR021meXpAzEp0aistMq1MJgd/ndBDrEq38wn6tI8+eWV3cp6q1ayq
0TFI9WhaXmsRgKL2s4snQWC/XK4sgSd5zUlvatFLWGeLTWrxzZxfTAJksRHB1tff
1vfoNgu/sqBpcjleUFROcFf4fvIGboacBgbMfunlHn+hQv7a2vrQLW1spVidN6kR
LQiZ2EH1k0cTg74KHH+fn5F738TtVzALuSHMjNCpb7vyZz2OKLMSMMF3PIgG/odv
FSX3yS2zujroqRRZ8bm3+FLUH01r7ETihwwvvfY0eLloOuBb3YDft1/MsvSpqCNB
6YYL8G21CS7SLqzje2kbnDW5ao/cq+2vfCSH0AsQ3N6VIZxXQWNEZPlqkI5QeiyY
Nd1JCRAQ+jce5EW0DdbFKqR4hcYqAr3rOis227mZ+j8SgTsE5jzbOGV1y/P6aBnH
gO7sa6W2H33Wln3IVy7Ydvt7JN0J3IqbUtr3TS9ZjcsQ8/gpveCJx/NEl7YqIfpt
WzdIqTS87gVCp3OhHqv/G2WeG+YKW+hip7K2sF3mZYQ0Sb6nq4BOL+DVidfRbo6x
YszvqwdsRxqDqZWGExtZIGtqIvF/9w3cCXyLQMO4nPwFoUlv1jcRbtqLzLw8E8tF
l9RXRNSvgTNnhhtw7uVRb3UQ8PnisxPL2AvItMz6o7+VsAoi8/llLhHlAokECX73
vDl1KOoTgle/BVIra4Z6+7GNPJunvSRKCXMIwRNbsyYaWjONUf+oWE0sxkQRPAfr
Esf5MnFcpwZGFSB4fSVN6nwMhADvYTixGu7Flxto1vqOgva6uuqktpX39+FGZh1G
iOGW8As+XhXR6/yzJwBo3Fj9Q+Zg5+7x7OTQqb0ctrizN5BbXpfZe5RjGzkHYQLp
3qHVifJ7k4GHTEr8PYsccy3Nouz5ylXmzDTNIDD8Arzx75NSRYm47gaLXTrLarkK
FrbznkmRA5v0M+uHbZxLojDjr02UMB4Pr8tm7JmO+CODqQL6iBuRu4Q+trML+HOD
c8Bbfo7Bb9vgl7MQ8gjeZnbXfbyGqhS02hI2rI1EjJoThvYU1GnvRqekhxu2CI8W
bRUettOu5JUp1tFQaEfbEAOXOzbkRn/gQhhGrOuD/o9oLN0Y8tPUBsseQ8Cyls6v
Coht8czpq0OZOvDs670NPSuck0oxJSaOrQmN0wLPE8iVK6zRNSdP0g1wWyFU6ylL
Hv3YdQwTCAYXBhEwVWhumSnNg1n55+G/PUwQJFNxNi6hRtFGGl2H+DWAXM0+pBnD
LE87RamN0G32VX4BVCyeOGRG13+jTzerE6HNTNNVeijvBcK4AZNx5Eq1Trei7wlk
DVMaWO8bwGCmn2WqwDOsS6Hi7z7l03VjSimlrsc+PjhP40QIOLxzSB9AmWWnicG0
+reYh4JHOPVBDkofySiS1ZnMr4C1Hqc6N85cr0bsyR8P0b4VLh3LgKH7F6ZOUovI
8dGu8AtzEJhJMvUfdmxxEnaO257EBervoQMz70Zg68RQkfakAkid22OjcBRvN1Jl
rQqe39MsACa6QlNXzO2Mdz3rZ04NoPSkyaMFUDEYhVIUJi3WxJZrjEuvnw2MsULG
HNNaxhtitkDJqxnYTVFyrhC8wOwWYSejbsOpNBnwQKCO/J9XCH91Kbezloov/oQ8
vAuW0TK/da3nOdg/mUg5izA5smJ+WSTZHnwvtrqTw4rNQ4I374THPt2Z9u8Mp4p5
3NlmjdkW04lX5fAQQb4+yTpN69dk0jQ/Yus5Xzbo/tMFHb+uZITqlIiT/f07zz2l
C9jxhfME3s0GGYNWB0+6VQeeQ1RrbfYtP2+5lgWzjJ1fMIfXo2uBBVfuSW5133s0
CVw0JyrMoRNMYBuOC0FwLJiMwjnaRdumywT53rfK12OyCwxp5QNwslCqbIGGsQIf
N9fWH5pT3ci+9oTkZ2/O3EuRKMvts5RCl56qSDnxi58kHR0W/5D1I5T6bMWL8O6t
YUsnKBno1O5SwZfBwc40ipMnq1OUkzbEMyZk9bMortERcwRhjk82V5WMpNBg4qiY
eacHhfqKwAxltOZgJpCqy8+07bcPkQ9Fj6J4HiJDyu4u+lPHsocb4Cy7RNx3YxOG
gWRzt9MkefRqgqTeV0PM74N0pAh3rOJDsNjo2uYRlrz6JvpKeZ5FRX+dkUV+b1t9
ediir9voDVdQ22wLlaV68DpinrZa9u9n8N5BIhm9YCW12K2fcFGv+Tlb6DQdykCs
IGLCFO2jC78/7+/bJnvY8HALhUY1tR0M1D7/XgA8qyhFKT4JUhrPmnA1gsh+IceV
EOhInbLt0tjutN/hfbZEMik21XIUGcOpAe4v+td8LDa3KHfLLKMML1xQJNo4RyaW
8RicMWbAqObMHlZh6lMPJC1I+BaFVsVBKWy+KY8g0Fq0rJQGosFlOi/HZ2jJhqsa
Y+nW8Z5ilqog2YfLmd3tF5yDmEMkBsMTPVQeabHt1QfnlV+zQlaF4snfYZ4X23LH
QrvlyWGApTXunnBG6wFTMv6f3422/mF+OrYEpLWyeS7SUZ14Wed+8mURc2sXFQ1M
PgneYfcFx8RoVIC8TQDZhaRn0KWKt3x8menndQRkg52ynPtWPyFuc14S47bTRML8
98E+r4PkSAhdHqLuk1uS2IIccoimUkCSHksfPCl9w3zgCnfHj/XmPqnvtxGEcy/8
QFJQrm6bQik3n7x6wkb1gP5jkek1EUh/VQ0QM2oN7Vj8Jp3WeHZ/OnkdXyRkbHB4
QE/UUd29yXfLFl8lm0GTOgFz/rWpOUX0ZsVRWBP4SCGaLBQex5wilQDS49Asb44M
EQU/V64KajG6lKzps168IVyMHwDczbziZ2YkiPt4WZUak1EzZKrgLxAWA0gZeVCJ
rSP0MW4w+f14kkodj0WQiEBVYIQE23CrgN8JJFy0k/NNDMrNe2CbsQebQuqPK75f
AmyzNd6mJPJYQFHW8v6JdDO5plXPQCDOA0YdoDJ1HJnew2jSePC+gbVeKhFyuZju
HExkGeYrcrnYAZMIwxxJ2PyAHZlroXaedsMSZnJBkSD+uh5GLn3UrXFK71wP0Ey2
tphAp+ulJPk782hPC341JnP7RB4eavtV+iJNyHzxm+EO01D38Hex7AhopYIuBi0h
FhaBRyu0Xwoo1p69aMe1hYFDxNIWwE54vV588N8UMrchqGErTBPTr1Qy8ZW+Y7Fc
9huEJxSFrJcIlpjvp4LesJOxD7CIzlKd6xs5z1xa/URcRtlhdNFcrJcDzalwsXwm
gyngw2Ez2f0FhreU8GAXywFTuimWLfGVsdLfSSrddySUtPreqiKNdJZEjQPJYlYy
IzSVax4joVNPSEiCP+VkDMn/vGfaZscSdap+B0ffzBjL9q50YCztMikn0oz9p5b8
fz/TCACWMIKg+mwzTWyIX1H29p+KH9s6JK2cGV8gqbAVmnSrNvW2JC9AK3I7IIjm
48Pnc/yYVcopRzq1ZW6QenV36etdaF8ljqjPI/X4zQL4y2gRcQoTxLOVTcXO4ru2
ZnsWs4rgg1MoFrh2lOaBpM606+YuD/P64+ZENzRRWqOMyQqNoCJEwn9Iwzr+CfY6
/mvFPwuwLu6thMKUt3UiilGhHiDSIGWxoD9/6wIZigzd2jgyqhIlPYQ5RTXSt93C
FBnwIBAuYsetrWGMhIpNm+1D+zk7TcLBUzcVNaYIWqrRRh7EdLGQDK0I/APcAQWs
52miCkytbEOCOWRXqMh12ELVBPtRpNowra3JmwZfQpxdlMbdc0VRI8Fypn8paBoy
NSNv1TBRu5dbg2TWXbynqGam91ZeDygTbYWDEelxvOl0exPJvSJ1Tem2rRaorPts
GGm1txHq+LTZDj1zeEMEoOM+DfxqU7s9DPQ1A8htTKJOloY9W5p4zA/Vs9bk5WdW
ID6CnGhxOg1O+w6e3gHthFTrNY/YkgeC9LI+2DB34O4X+0jxbGT0egvj9s2//uor
D1TiEW/XNskUxAvD5qvKuOHHC66zUzsMH0q4sPmfIKabiWnGtYCXnXUp6C8aReGY
5EUbBWW+wzS9cgx6oHA95ffQj1cfivwRqXyHxV2RH2OhllHNRJMBPDBkVdgHHfYd
vCtpBrBp1Q0PdLakD2IgMSAmYqVj0gRHqozIxX14hKM2DYtqJ3eVjSPEIA4TiLgM
tgfOBN3GQXUqX7TDOPuNd3T5R8jD3bLi7K2bkc+vrHlxwPKzcC4+Q/UMmeK3x7LC
pZGnby7UslZ57xrdYscSC/sFZEnbv/j5RDeAfOs5wVlHA58GAXVToXE/SSvX7hpu
BocXEOtG1OhOzHvj1+OdCoDdLZ0DlU4o1CI+Dxpl/NKqwqKC7i/2DSSfPCW6QUpn
dWtA72meop+b+XLPjU+OCi+BC104DQ2/NZuBAF3RSe67S1TztiC/8KIiBC2bUwCi
gKzrdxj4SkMlMdHjAhiiuKU4sJNTkVShOSnq+RQnpH7dSOZBIA2irDbv6pZF20wI
3OQmyd/2VsmXUJaA4WA+uTkSKJmz0pitk/T7WijiOT+MpMWqvVgPWlTj5bsHVhrl
4d/QYOmpHDg9M/+bgo2X31HCcfgLctlk544fCShwSGMI6ZOSQiqIxdvQEVr9ud1B
YoYtaUbIiOUK+d4hlyLm6RKdBQtNkQdpkvfYUZxbD9DcJlKj0xOCzwX10wRhCoTJ
Yz8sVEIm49yUd9GfPF4HcZuASqIxAt2XoPQWJpUnM7ilj2DmdWhQfvDB/KpoqHAU
IYi6JvcwnembNQage8ZkxzPXHYAHUEGI/2PvKi/3jF4BB2tZH/mgISStSVu3WClh
DKuM/RJK/E2OdX2jvpYY1C3vCQ62f5s62wOJxIf5+N248IsacLR08uhEAgRhG+KW
xqjirhq7O0+1p3leInHg/3xIlOzOYgDIOl0rTWBePh+EvQ/kyO590D9XjUsOovyX
WMWt67c+aeO2xQ76m68N3aK9hImLYJ5x1LXD6exo3tBUS3OVIFe9L0VC4FH7rN7j
hKDvayi02QPYcmDUmLCC98AXlw/LOtOnsdjTjdYsaHrx8GWK4jPo9g4D3lTowqb0
CJqY4Zhl/9FbFy0q5YjGDJzABGRebjraWU3X3XRDll+fb4mM/ELJGsJgXONy8TkJ
jxiRADED1iwgMe8gPUlstn0zahpPg1karK5iEWOsIIMMhSrkhm32QcMRXJYD4EIp
ExC8NKDJf5vhp0VWn2Vx3WXV9fRqJejs71UTFv+kiB9hlVhRhVd/nBx+tMeHLn4R
NcUqKZDnf8QJF90NlDNXeykZ+8X14xAVP2C0NhNQzPPyrPoF0zgXWNGP8TgimZ4h
IBacW2Q7muB59RIUMBVsS95iuw866ssIyrOpsWmrIsez8TfLwFsX51C0DyCGDjAw
kmgcfrQKuxB+sbkGLMNmXVJ2SRAKmWWpF5Xu3Mmr5U25KS1j28wzkkxCDlEIKKrR
db8tZS90vIx7tYtwCX10FDv/hE5CdvulxzBz5k1CCN6471n2M7PEqOMOc7ReNSnA
cSQuKfXYSIPyVlXG6rNZe62IhOoFit0GS0P1zoV61anM/SqOH5cpEEhxmNhH2FH1
aBsd+ObRDaMfpoqD+qwVDYQOyOuSttg6KeLD0z1+7lb7uVPTuVA2bXiThLubHZ/8
YxpxrxypndDFKihc81Q7rz2JvDkcm852MStZmoTd6ONLUEi9S/CoHQPlW19wbbRO
wjGBC8jVF1m0HXUjsehOOV11RfLIYUctyf/hZx1lmOQ9vdCWiher3RPbTNicoHNw
5UBabYnzIs5pMAyECDkZ4s5XkmF7qmAYFPnqltLfRO5kTtgDIh+4jwVAS5WTX4F3
m571k4zHaUSvcumpQpWJ/2AgBFFN1h90r/CfcY5wOzygLtgp5UzmwF/3zKoZGjGx
csJdE+K+dsQAPVPE/zPPUgNqK6WBue5FfR5CPu8TTuNNv4R+pqPJcAMRfeSibfEK
zzCSFB1RJGSu29GIGn+2EZo9k743/97BaWYEExIWGG5Wm0tEqEVbwmDMK/jCjCub
5M/vbNQ5X9VDXntKnCnL6MPKyL2P0ptUDmqSx2C8iGXMNNzEirgnf1MSba2dvLfz
yOz/T9ctmBLdz7CvXNUyUNTO6TkDHHXRcpmYSkfCzsSuZ3QZ0VkfYQ0XMY34n28C
v4iysfZ5/KU5a2xmxLzi7+kUtHHSPi6qnW/iyNG9+QimoHRt6/nY/OO2iuvxugts
j8IM3Jq41Hx0h0KmUwRIXBS+pf7082BqizOQXWjhdln+0KdBU1Wf5qgz4hsXO5wZ
oax8AiwCvBIQO/6Yg/WFWg7Oo+Vhf47Oq873+KDZmny9166x1hxfd/NMDC1rV9ug
Yw9RlvttAkhTMRbSesSQj8Dir8XC3Me9Bet3ME0dlOqPpAtVL/o9uZd0ysftQugD
PWPX1FfgMnSifnczXcWJXcouPxrmUYwUs1lmxjAO8ASPbLWF9ZB8syFCC+emW1M8
HHqY+XcYUu0yTNcE7y5x3OVzJfv0C9eLf5TOusaDI0qkDQ5jHZ3EhjUQmSFfAx/j
8/Ikt+9n7HkwFykxy8XYaTjJAqzRgk0CgqodHx6K8r8MP3tKPradh0y36UgP7Brn
9j+mfRnE/oLxjezPJg6w1pEsG8wgJbUYPiGKg+ok8nZiuTCVxB9rch6iNNDOtEZK
nC2ztO4HpP2a7K43JxqzcFADE9o4BRrF2FbgyhmeZChH3hl70M+rWH3SoEJ7Dexz
g/dP6GtbQ4hjX7a8K7cVFok3Z1ml6fwhBFwp4U4Nm7oENgeus3JmmCFY2yopC9jB
BI5uOCfe4FqhXs2VeRdktmOVNYCMseOuWqA1lyw7RygRiAWKBR0vEiXxfcwwkDER
oAIJO7vJCk9QaG24vnLEnE0atOBg0b149pObFWKYogizW6SLUFm/DBZodmisRvZu
hFHQC/4hPdFpx9E/2Ek5uJp+WJHwpyrNmRj4wpg7tNqv5croyKpLgL8gAr8GpDGb
cp8wAYMZIagh5fWmGI0USEixssqCDHf2Ir1CVzYDxMW4ryFP84utTn6R3nTkddRD
7M8ilHywfSu4cq5eUgZpvmsIztLvpX9YukznILPX70ps1B3C4o01Kx6/vb2AQap5
CjmJtuES3wYS6zPW4mjkuVy3Ma93q1pXEhspwKUw7CNUyvlaM+woHsid+356SCg+
7vuUBaXaCXkwvcRRhky3dKY/gkqel5yCAor8yXx0i/t0OGUJ3kCtEwVib3WkyX9y
ZoUya0Bkkov5ejmgKcNwd1m9zzhtJ5wBhi6g+pn0B0s9PvD/Xf4yJn+EHUcmGqZ+
AU2b+MTGAUYCJoe9gr3+mZpOhJfOH6VMTc0mAmUlhr0hieswESSOzx7HW6NgH/EA
Rui8QcQ2bQjA38yelW+JCduouBtS5igaULLazvXNH/CbqqULf8bvxfQV9lT2JIUt
mA0zCISjOlBdd2PqTR4QDNH9TbL6OJQ98PKvWo7/cCOJcboPCA4CL2QgnOTXGpXH
tO2jYAxhZHEi24CtZkoGW4pZy5X4PsqZAdC/Y3uFnXtR4Y+A3I7DoDZKsrHxNrfx
N3KFZWy2Ulqw1SysDa0YT8RrwIx3KoiZFEgGqdyypASQf0P0xtPBuTmu1Fk+hxkl
Q78Cj+j/Jk7mPhXIFTIA/fojyMVYcnK4d+suMZ4M8B2ASYxy1hRSoWyhKNnQZJxh
chWZ0/3+dSrx1f/mvfqzW90+bnRy3uYINmEYAQ8I1RkyqB/+AeV6Yo0Ef0yFqy4D
SHYrCVZtNtanf6xsCwyQYNPOwlKgg9J7DqkGNCSWhPHW+zDfbv3DdIjETHm87uGg
gdddsp82wgXE5pIgkgEd8RRfx9OJAsc9SCU+CvlsjlEguEDZTwXxp45wq/fFab2z
LOW/CB40aOAIVk+V1fjTClKSRO0FvsCBS/KuoW31durDsFlap2Xo9Elxbu158g72
+hbecHACiiuaTNZwKuIC0ccK0HwpJgV34NE/7ECklXuJvV0N9fOLh9cJWkdQdx7z
fOAbzlV8zzJt7kOOnZr4b2o9gInt3XRXokM431HVFQ7c9MXY4rJ0G0RdLsVBq0DR
pRT9Aa0Qiuov/PjXbwciRlxL8l94mYa7yFU16R9oyoJnVT5SIjADJQo7hNJHQw6E
/f5T9U8tOZd1pW4iAPhtCB5++weGxini32/pnjDxnXJFL7PaL2/jPg7+YskYJG3u
t0BKnpTHgZVhEVAPvBa9VDgP94TdlDxt+tPfFS1K8+elA8vIalwV1YhAkdby5rXK
4cMVD0RnOys8fRtGp3B4EYvDVS3Jk/h6flNThIkOTmES2USNQYsT6md9UuvLvdpE
Emo+ODm2EliSSZc64SnUAPLyqD4yh08whItMesA8otSutFrhntBDChV67pfZOxrX
/IQkTRm+MCndypI/ATWjI7E2G0kFYg6abpTBjmX+tfNX9S0ZT+lFhABxOEm60yHS
rV6knhkJlbFnMVV576khaiTqL4hWdeJRHtHXCciwuNJrFPXTunOWFpGCgqkiJuMR
9i9wfsjySOZMtkMIzsBOKYHVV3uEIbWZFORwniZ1SqukILAkoK5BSYxUy68S2kFd
Hg+1pLbA4vvZggBWV920ONhrHh8POXC9+L8/QCuUnD4tKiBqlam4Zo7N775PxjTt
jWce4RR1MQAUcAwO0Qh/OzANLfuMpopG2w5ddSVxnAKNihnLgoCRCHmSqlOKkeng
43e6LALhygI3mNwf2zarnVg+oMHYRdu/WoWaKMq7opAL0gHlKnrOtuV95LpiSEbq
FGuRJZdrVVBDahOQvZGgXpf/pKrhKqIdxlsZ4zZBgVmE3IndIvW397WaPs+ldzPs
zHxcknGYU7FFKPrBm6FBZWcLo3J0oe1JwzmA5inHJpZUEjj3cY2YXbeeZB/UM1vO
4wGkvwDZ4K7TTX5gn4re+QwslfZyLrIWJGwGHlEcMtPnVf19/LmfEkxVgxK7KSE6
hJR4nMPUBQrhS2LiFLxbxS6pmlJ65jxXbVxaZmoxLNwbwbUl7qdhnWC5dHpxsKC1
hZzatLeDYV9Tad7ugW9ZlhGXhry3+lcBP72SD4vPEK1Tya7bNLU5nHZOWbkJ92ar
N6bhM1mQPBiaghTxb7Gu48zGtx+YzP649M8kcuEAzLIz2hTfRO+9wYmr9ohYPxlu
wqCtrpJHW/KQjyH4xb7N7EfWsRfMhqneRrMMi5RbBy+jSCdqk7r1N2svKB5rLBJu
szYqvllX60oehq65tza040+dogfa/y8d79t48a5rS8yFSZoC0F2CSQ9sBvIto239
1jYX9okxZ/J6BXqkItqgIqGyljjmRnhz6Lhie9gkpMSiKpBFQqZt3W3WGt3NlKlH
qDSVugcDWNhBCg2xX6xGdM8tVaRPdriILKmPs9ekCbiUNpz+nrniZ+hZAptPrJ4Y
XspOqMfZdyJ+8VbZsyYkwH5hegpZui7wrrqwfsipLpOn4AXBErLxdUjv0ZtmfaV2
pUtSwVq1EYxKe6/KAqQLkF9MHUewwhywLsF13IYzt/Yn1SigCZPtsfcG0jRmOTH+
zrYMvX8feOU2OxAIQck1lL+gaVYK1A5eZlDR5H1D5T0N1x3z19+4XllZU9Mrd+j0
0TvXaJkiVBMt42BOY3qC/Kwt6VLh4a+HE2pZbfQCSkKaMa30AkgwMiCHNYJkDWuE
6Jyky5o7QxJyfDtWaLih0Y953/Nsk8HSqAu6CA06ZGrECGWvEqjTDiPvvZnZZGRe
/16xRLmwKZ83V8mx/PBd3sF3ZOa+FejGhc9g5MRCrjs6D3VPy7qvxgCx0rSuoqQz
qBNxbjHADhEZEjHfrZnr8B8Z3MiXSC8+JcSFl/lips7qGqFM1Ek7JrjFZtG5boYl
h8pa28PwYkEhqRySE469O/wLCKCuq5t1gnJPHl+JofcHuWXEHHjGwshkLxYGZQWR
IXvpIwuaLFzvPxvuKa/EH1E/Rdm33TKfKNWd2OgioBEMKD/NCl1i2kEhcs8Y+k6u
kSpnPr76BrvwsN9YBhjrTUX05nUMKIlmF8ydXFJ8VoQpz3fT+fEq7/FM+OxU4sDa
jXW+0uYMkKn0Ccf+cUjWUOJXQXuZFrWRIZJPu5n3HFgVK+MpLnNfFah4NAk1nePg
07FJABRXKuV/DcT7aKf65LpISVOEhodKOubDzkBUk4/VZ6DITSAWiaKGcRrKi8TT
4ziItjE5NFmDX9tbCQg4tLpvnz8XwNX6FkNa6MBSY6sWE3MNPplpoa5frEeXJm+l
GP2AFj18t98saIROIZukq9/NsdeKp+Q30MLcVGbjp7PMRDz4K+1JSPiSl2h27yM6
Qr0zFk4KzyxUHqBinQyglXU2xH00tDhHybu9CR+e4bqdcyvse7uuVhOsFF/zLweg
D1qZZKz9u5z2G1R4A07/hppnViD98bYlLI9/2RB0230Aobdk3rOcSEGUvVeGu4hF
HDH4VfqbGWh1PVlB/KsANUVcPu1ClHRajFmFgrsPZAmcmOyCO1ykhukJ//8gz5QC
FX0oKkbymUVpfhqEehUdhOK491utF/c5utw2bmcQgN/G5fH4U74rBsVZeuA2hslU
Rpp0tnFrzFCPFkq2hZW8qkz/1mH6/8cRMA8FV77HxU4qIIh5FwXNjcXYn8rwTiyX
d8XcywUkvTQsm4cXTy+LVkyKZ9CVitvnFSAqyMlN5kJrZVmZrVmTQlq+DPK3J79m
1AUg+cCCgZq5m881axnNfMY++3lygLfcJJZrQ2denU4pwIs7X6AM2SmnSXbyRebS
gfVS/h4iBrPSlSaaswzT8W/GfCg9D5ftGOeoJhh3kFsP3GyyfwUbmkdOrYFvkkAW
jlNPo5XPAHSB5RUm6a6m/a/sVc8hdmVjUlfcr5Bho1WhgYM422g33JbbBkJ9LUP8
fZG3+RKXiHyT1JsBqn7FeRAEeKdFY1fUJX4E2dx4qNm0qMl9TsVp85cAzo1MNpis
L3CyjT+Oy6BcnZjkS+nLvdpo1UUhT4uHoxzaZbk6stGAH8TzvatX1s4wUoxXG/kB
O3iGQZsI3hg7HEI9EAUuZPattgBFhrKNvrC2ejBYaMLpAgf7gmGBrmVEAuW3rzOv
aJGINGRJg1NqftA3eZTyvONNBbu6Og91M7y3OyS5zlahmLqOuJs4q04Ts4FFYOez
wl3jRuPJTkTz8TrUnk7PzLy5D3jDh8qcArbWDis5sAxUUs7XEqQJNPIyWhOWjfyX
myHizd4SOn1uMmeKMGVzvHbHN4QJnJI0HZPd4/Za2Ik=
`protect end_protected