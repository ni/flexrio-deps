`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6656 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
BD0Uso4m3HP4S9U6YYcCvWdcbCiPVeJBw0rvVEd65jgc2OxcQF7KKfiD8rBemZwr
WnyxIDKEAv5EvHrMKFP/WnjPu5JVBo9Mj5chx4prjJG4C71NQDsD0f5q1+Hsf/jI
HlGauLqoO9ThDG2atkyXoP9p+Rf/CIHv9p98oD82PgO29xXII9vgZ/vbbN05DrGN
v4s1nZQPNCCiHL1bVXEN8no3DH6cHZiTPXVeOORMXw+FKfsUx3KD+YG3LhPpLCXU
Xhw3GkssDBYQUAqgWj2ofzGrGuCydkA1yS35bNVofuZE3Nw1vkziC1u6zA9nxY5e
wp6SLS4oD+0wlmX1njWic7FEFMpHDawCbRRC+FrtcbmQTN6S9LVzVBEghWYR2YjH
FDHVqxbhZ+v+jjVyquoUnwlfaCyTMc6OvArHIcJlMl9hiP1EAwsX3MnBgEOy3zfp
gEfcEELIn9FkJnZSOKgOOHPlpYl4LRO9duzz4NRyiBCRNuIo27Y542MG+r/lTtdc
Qbmdds47gt8RTK8PTHkxLn+d6DwP7LhQ95X5XDTpIBfhNuzHH5RI/A8t0RrBnQ8Y
jIpuDSs+iJPgBOwYngz9Rp/SaDgEfgvq3JX41XgH607bRQGNnGpY5ZHJa3exsTO9
NZ0M9K+Q7xV0q8cxffveLKEt0oSgg65PBmI1JO8tGrQNK204vn8YiftUv5CdH/UN
jaDQm1LYImkF/xcpLMqLFXkuV8MITkSg9/jazHJNS/HrdMeYuJVRWWNrPus1ZRVq
+vw5OjzEk6oA0A0Bs/l/bSezodwc2zFgqpmAb1ko1r1+zM/sI4qQ0ju6qFhdxnWM
WdR/4K+g51aq0D6qYDSeEhDS69twZ9GWyccZ1CPOTpVw+9eBtgJ38io6d24UkztK
AlkD4H40DAkfgLMt3Wu9VCtZS+1PaGLSJLZMAMVj+gcD2kArukpIExWZFXyQMOCj
s1YWVPDwZmMCoEO77fxjSTajUFPWP8iaUz2FtXqKVrzvuV6sePMq4LD97QKEZwtl
bD3dB2h/TVBsLoScfFIebk8FSdbMWAZYyQuwF3aUIEdt2GO7mT7ike7B0w6T+ob1
kLtFxOyqCfgQTlSgEN24gEf6aYaD5bsF7aQTGFacD9JeI3j6x7wdDv6aVO6pwaVr
mlJxLHxQKwwBaVyOYwX6OVkk9WXlOkcCAVlnQ6UVwBWp2m8UAd4Gsgp13H3jjzHE
sOMB0B0eJDO4mq3CVbhqdqj5SjyGU9Gf3NsYiwmbCbcTMTpJ14pv+JmCrwqslLyh
1T5ESb3+66Xs2SyHuilfmRM/vXHoOy04VAMn4+9HoXtw0qMDRRKAv3woFP5YEo8b
HumAvZ/5vdcycSi9kri5phd+I87XWWe6uerHHdv1TzlY+VVm58SfA0UplkgUL0BF
vR+QNB0krR89FuI5UVeI/e7Wy8Jc5w70fhUklzWCxNwXfGLLG35FJ7oNjh4MGrFo
9Cx4HWX0z2qtTkK6RGAM9JhNpDlZU2un/dYymIVJnqSytZFDngOwfuNn6l/lB5V9
dA/ZkcM1E5jF9DQOaUmC14m4j+GTvioseZvXvVFjpxGtcwBxoiOrg49fo/ybxQyG
sPYFZdha6JA9FpcCMbSr2kqnMLhQDAaT3MGWo2ecG/6E4jLuXjQXlD4zz9yDYE8d
BSuBOIR+0NYwn8KYHZ8+QepiqDo36HyTQgmkvwbx0ASbYeO6yLjXyjwt4j3EsNeM
GOPYVknXzYXwSrHXzPuQ7MPVaTXeWck4wgIPryc67wRHM85OXHE4THlPfA5fnAga
LZ61y+6NBoNjCC3HmXlpBi1OCah0NsittrjsWWuPDlaJFPPX4BsE4B3m0HSfZFGD
JyryI6OjNgl/V0ctU6iCgr0qJTUNN9FLaMAs65AxI+Pk/khgtgppNfhS0ICmgrKC
3URI9Lcw0sm07EhsxwQ7jf1g8cmo/PLK7Jaj0GiJch7fuuVkTlbO6BK+jT+otsPO
URjCTjdvkeSHI0eaMZypKWnE2Ky+tjKwa/79G7i4YecYUgrs7fZVNuxhk8F+nakP
aXbO3mDryRC90UTRmE/iPLl8/+qztsjYvXCf4mKj45aJWoJyhMEEaT7C4AWKyyE8
wb3WBJmM6S+HCr/QvifSa/rbKbBG5IEB0OjpW15+nmsYi9fvwg33G7CBP56bVENs
feQR2Yqvvg8YwpenDCnXLGfM1xB2UNn0mgO510OEUlomwAfCli+Eu93a/cbzuZ90
lQYZS+bBS2hPuKPjc2ea/kPYNkTAD3jnD0/Nl0s5uEqW93FJ8F+h4rclsX7yRVJ/
rbedlqvqflJvqK1wAvp0XXb85GFp8r9QvYgoKj+bKtSdbyZgnvVVdFHHtMR9omX+
lwQfnet7M8v6BPINlE2NxJaDKkdBG+8fOxf0WbcGO5FPcSll9rB8+4WFhUz1oqNQ
A/8rePh+fSrF1H+nyP8gQLutgaRy4lmL2uHeAeW6ISLGkKIvc+6mrWjKwsRqmSuX
QYSfxmNytj9y7jFr4u+L/QhPWPPYUNjnaxDQYAZPcDrqoflVQ/d/h1vJm7DFwbVi
ZX9hzHelwM94VXZdA4rOS6bwjwvKXUWcczPxn0fE3KJiF0PbW5YdB8WphtbIH3tn
5oGr7+6iVqOF5cVqinh+Rs0AxmdjCyh3iOu+2zq49cRNjrrmsdGwHzKmFlL74R68
vviv+i6cjVUFjhDkWdP9k8YIK0H29/Q+PsNaxOCEIdA1+X6p3rqj+ad1rhzDmcYJ
dy6K8Ty5ovV1r8dQuOpe/d/0AwU7C9BUC6hUis0sbNoWnLe/YhI9qe9OyXQknrYZ
FRlVBTKHesKPxZS5MU0IUyAAg9JilukRwG58Zxcd5KRvCSpCPyHKp/hM1OOB/yTI
YR03PNZAryuQf1m2OHU4eIOEOcQZg1QAv52KTXd9h5mZwHH8P9ihiE5FWvZ656wN
yAxpG4FPK+gfW3bKsbTVZ5h5t22o5NZz9rJTHJNrxs9d0AaBbsHjT45NZMUHFztb
iehXHLZrilrwgV28qqYV3zBTiT858dIxSA8ZcyUgBKM7tUMd9gURKNLa2ESvSJ7u
UT4bsNdrsX3Wbt925z65HB/e461z6F7M76hn8e2C0VDjCyGC7qH6qZh6H8X6oom2
yHiWHu+pIwgbqXYjbtniunDuzLZANW/03iAQMQ/PKRZTFYAKpp9OlX2FnJoh/bqV
NXgr/+0d2/ie5pvD7j9xD3NTgNZtrdhiss9nkjsHSHS4KnY7h4ATVW+GIRyl/BhO
UVH8hedp9ry19CwcVsBQmTdTmSt+fRnbISdJMgQkh2W1ukselBkX/g2bZF0DQZ4H
5ZyyeKtLbMD4nCR0+dMEGTqkZFnOfZkB16YhzfC2kX7Q1CwZFZWZr8ypP0r4Kp2u
JJuh0EqeyfqH32cNM7oxb8oMpEFHc6Sb1QqBDICq4MQ2GLfNnopxJ+OrVyBatrqP
U7h9YoEWPbK6g00Tvl0VFX8+WWmr9I6MeisBDuh5t5XYRYNMTgkKG17ycDzAqN30
IQBlVOKImfWWGabey6zRe4iuB8FBav9b4RLvrF5rFQzipnm+vxRU230verHn3ODq
/SW6hWnIez0BBO+agI0Nscf2gh+ZuBkQBothoUb2uBR7Cf7iK3hi5Mj21cEXgdHX
mTcxOXJsO8NNzQRfKqLVtiKAFgw4uB8PnxL7anP9iNQlubgfg/Aie0f3ft3ISNS7
/V7wiy9cxlylmXqLvBmpGfAwMkZ2vV9w5Xfnk2FkND4XMqiWAuxWW3t0MG+r1uIS
02R/bzmCdGcbYx76l4s14esxFN6FwRl+jdtFS8MgEMAy5lYUhmkNbXjcrrNkTc0z
664qPrQG+rWsztuAy4HXxS0RfHhu8RMQFNjJUEscJed6aUMVPzf7YFV/kjWJc/R5
4mpvhFhhFgKh4bjQVjn6o+g/7O9branp62FWCK9RcRpa+oTk4NeKzwiWvJPnXW52
eZLlwkjaVMSss1RBmhW4KvDEhJjc++G6orpivMmJptr/811sYkTNZUZ30zllw2IQ
XdjPRnTOGbrDXL6/xgX6JNgVgqsSvXfcvC/RHFQ7w98p1muioyDz962i8cNpnb27
EDyZw1HlRz0c9/QPKR2fPEOJFLfMycNHxql7I3WVg5r0rCqJaFnpQc59w/bxVAjd
1ogGyUJ8vQNtF2haNiPVdAL7rR5DBhhD0U199JWGCeFpL2WUTXj8qUkgtah9myzW
zXKQXvepiEHAGNyXucffqoWbCu8B15sGwLQLmQyuOv4GvYRmAYpPfAWcDmc4Dh32
uELQX4MT9igGk77hzQFaw/ElotbCgyF5ZwAomp4T5dKy6GWGfzeuvq2dTQn9pUzx
YghSb3RziXa2iXQWh5lyaBX4/S5tjRzDQmE8q92KOBm2NVKQ3x9olA+dg82pr7gY
RXMDHVHd9o35SvMrZClnnIjmXbyi6NaHQ2JfjCHZ+ZyPdYIQQiRA2tWNquaUi2/s
dYqVuSiVUDMJo7YCNFDu8Is+H34BoPxDeJQJDg9RX4UGEmEvQm5w/zUja05OJxRi
dhhpQOldygDiq/4RajFcM0ToBTorPX8njVzhr1YQrIl0sP53HGQPzawg4rNhZYzY
BoM2pEZP00CqavVzzTTXpwUui41EZOfG3UUIBbc5yfaOeqHxTsqi6a0lmgIXDqFU
OiSbr3Jq2aKSzfG32/juoqgVkY3Sglja5NTK+iGwvexmUsnW4vJuxdiZlbBjM4Ve
ELmdo9iwI50uJ+r6lehobt5gn4+LnL2n/lx5wIJZnhg2mskyEtRJ+ubae0/gFZN/
DlLMEwu1Ow9KHtiWLQlgOFYPPKvLxIJuhRZ7EG17XUF/EwBeB4eP5m1354W00qG4
0YeWPXEsz0AAJua4lZhrESHiKZfZVDkqb1bu+esx5Gezpl3pn5F5RiETPq7EPu8V
GT2ymLI+brCun4icORXf2R2DBATacrkQyqLcXBKUBFrf2ZIrGWJwuxDcp3MuUOx3
RCARbEgj20I4PWtAWYDMi0WJ4gk2gtWtOMuncIjXBd0XKqfp2rtPqjf5kHcyfc17
7ef3A4n1bMbW/8PA8X5CXeOrMyhw1WJ80SKJUbp6OHmibzacT6VoViAhy3bz+Cc+
UGrYxwv+HrGT0SQJ/rXa7o1S14MUcv3Rx+3atSNpEZT3L4vF18lfA0OT0W4bNvwu
89w6AfM/rV8N1j7SvUNSFDXR86L+pUOV83Atp6E1gsd1RYQg4sfSCPq1J/sH0GGM
eu68qkhbgBzgqX+fBduWEvv5Jn0ynAUQ4nrDKEVYdmVtYpz1kg7JAOWDrU6LOPqy
06J3yfco2FCRWV2LDfeIymdmTAXmR5rHlZQjnnyPvAUjPdd5IqYYHgh5JdcBJLtz
vMltsa/bL0ocQjK53LMu3uaA6S2Z1PtB8RBwMKnb0z5KxKJ3dkex/HFHwTAfj0pK
HYQ1Ml90XBNveqO64vQnvUI4216CMUexoJGDZJxyDmr86+j0g7yVXCXohmtu25WD
mmcn9/zITc7UJ6gYyjI+a68yR/4sk4S7guIBhcHG9TUPUelxuThYKkLDrve5DIyy
YeSSMZoUSjM7K2RmHPbyvxU7R8ysqhGOghHR83obuPF1tdmtY1LsdN9/a18wMY4J
vBJVS+plaBlGaL9ggiNcN2swalkFiqkKUz97Ti/PPnG2yRc8oITTx7Q6a9GRXq5m
ymbkIt3fX8E5kQYbtuuRUlJ272ne+M244K8+1P1ZeEkDXmv3MKqo5jCJ2gCdtlQ8
mZnLi8G2bVGVqRP9kx2eSXJ6EVL7UZEPU4ixS1qEZHxQsFq6GlRjiYJBMVweg+UE
rYofqpddhNa3F/RdiY7GBSi119QRbbRg1kQcjhoPPcerHbWMYXjJrRVTHfxFPDZ3
JphE4xcMAO17QCK5q9RFs98S6Wv1kdjWzxZT4Kq5juF0ZfRafeBiLF2DMnCzJ7e8
ckHiXlsPnof0MjVJ1C21zsPfVrSvQvDjFgY4dYXQlQDxkbCD4VEpEnXzD8Sb8Olc
7iUZKYhqMlwLWbczYdDLd2L/g53+aVLohRUHohfsVu3qtTQsnxSjl3vgV7cge6VX
ODEDv+VuBXYwIGqNKZcA04LcgVGGFpd4ZIn6FieBNXez0Rtle0IBffnaXl9J35rK
TLuwrudL+Imqa4zjWAfuC+7tWzPt7naJGNKumaIMHCTZhWyOGohjVlgWEOtJuVCl
4Ci1ErThDfuQNFivsV7+Y4ouo68AJbLvhSokiFw9ugLcWT42ZiCrUOPN1kPyULGB
uMkOwaxW6paRvifJ6lCBD5Uj9ftujohZFH/JDu9rXx9YZpSz82qtr9jI3t9mqjpn
j/iV2lRSK+/qc1Kq9gdodDOLzHT55CZvbW3KKiCkxYkylXjuZoOw3LHnnzYhvPj+
8pbazuClNkZRz/4cANBaCxU6X4b2Z85wIY0oS2znXpVApZ7jxqwlPZNjst7Exf9Q
DCAyxSrWOERkxLKukLcT8ElIE+o/6ScKVW9CKH24S5DziQ0lD0TwXS7YMO3ls2iV
JhnMRKw5ra+XWtUc8Q/lNMWPvOl9IYyzIsPvQ5DJMS4sNTSw0wTuHc0tF14+41ZI
eXVRKpGfFcbiolGrPz0KwoTfBLPZDw4L9Lf9e9kuzhSJ52rifvxEwfOXjsn4onc2
8kBL2VUjlVEd5VKc393z8Z9pCExYJTV+fU40vwi4tG98KifM8rghwIBzxXMVud60
RfLEpYXJFOcu9kqqZWrX/9uuas2/akV/5W+DjoROzl5FiO/7Vk/c3OA9TO/wJAn8
hSza1d0j7+X1ZpFQzStj3bi3nLHewx88Nzdfg+xAY+9uGpSHMO+dYvoZS06b+DId
9WTT0PFRTVaTsC6MD4WljImOZt3DQ+XNbaTm/1/SiMIQVd54YByK+PhHU46iSKVo
FmrsQh9UqIDb7JLL/Jsdqo7RUjrmCLAj20cRujxT9tGrmpoSCAQ56TXpbi9z3IbG
gRMlohhS9o62KX/w13Oex9a2sSYdNVW+o4GvReEYJ/bHN5cDJbnhapvkN3gzP+ta
ZcVz55GxPlC6SVp0HP12YQqKZ8CqslWX38uFXWObCaTDWzuPhIn8SqXf+PB+l1hO
bKC6Fwm4ZndKdvE6KiDhF34lW8ccz+vSY+NJ8HEn0Lpzkf2Vqp+dQP9LfQ+NJ7VS
69wgINrq19d/+BZw0aBaakEdMbcDEGwK+qXiH7Icykp61cqw+Krr+oL35i5OkjBO
BFJlgfDi4P36jFlT7gVsMz1fFmuGjAqmEgdNu+a0690egQRwu8xRx/obc4fUZ41L
SAfdm1hqxnAMgM/z9cT3dj/NCG+3nr+o+klRj3jNxvFkHf02qm1NS6yO304/I/th
z5jDMWGE8vbQeP6qxeXt0CR2jclwESwQWepDm8XrXL/vCbr/KsJ8KLKtqCss/YWo
gfwIEV83P3YsHg6csTjEdKIOv/QgCZWm9C5Q0UdQ/dHvhnnnle77I1OI4a16/XNy
6J/aFstWnsSHFgOCHHpDkOHiuU5kil0XbjqDN/RHDp6Wt3y782vULvafI9NiAnET
brdDlDAWAZGDZp3DKPyhEsz9OjizSc4YnEe+s+qsyqPXUdPLf65VYToiwyfVk75o
gJbrDmcAXs/dXmL6iWqHhHmWnDpJgsabT1eIthFQCBbZRx6YHSJcwbbFBDHS+uln
EgjVKnlevP4j5ySxgBk04QjJo/J6cnVjrjRsrcmLZPLAzVD3kg115qQ5xgnrzB2u
pr21PaDZ/93u5u1O70LprbhcOKvztJDHNcWSevYdqluHS1IuMGrjESHcukeqB19D
JfWWF3PuJNJX88zPFflxeU8P744OMiIMDYHe1FmiJSbeH+GvfFhlhpvduufr6GKw
ws+ilSVJFXV2MoMHtaQw1MSAR/jSUbF1/BkOXsE1dibzwYyYLKT61KLA1DcYVmsU
gDB8duZL7ylkxm/mG5fJHEu1/ZAwbSQwuvdvLy/anaArIP+75nmwXVzXcfSuJ0+f
wflGyCQocfZSp1L72wXbcmkIrTMdLCeuC4SYyMY64TrVlU1V3LxYGTJ/mhyaXkbZ
tOtJ5zmSAeSgo48lQaBUmybNchn7rwaVdtLz5vBlwdrxvAHLZ57ZoEcBr+jB4NkA
e8FtBIMBiqG8ZyUhfhVOAJHTn+nHh1nzFoggFO1S8QcskLhU4E/vcbqswkFHnCLx
x0fKZTMZ/ce3FnjXmhzqH6k/8jAqLKQNK5SAz3MNkijAHLx0OkeRkPNeQlQRFWHV
xsRiot6j7+JaW0UBqvL1ySxSuMcGE2zmAkYlskyFywHluaMNy+nk2CLGrL5Jo86V
QqTETD8WG8omD6i8yhik5ESzZ2cAco6/6Xnq8Sr1KAawZGCL5w4qHW6BgaliEQoS
wB/SP5I/XgPJ0ee9QZMvP6ueUwwzZ48ALUbHnoKJcWdmmIjmwRu10U6mU99bZLZp
35wAk8fq/MKvZWtdMdAS5PVTEvKi0pzhcA6yvxYF+NySP1KnqrOO6LXH4/Mg0MJy
Go9qJGXDNokJZAgzZJlNYwfOunrEVjH7x0G4XtrYThes3AvDNDRlguWNrlQYVutY
3SBsrVkV036in0TSsWZ95+UXNTRkZXLwpeUYJdl/VZdQkU0kzZPkZ7aux1xLntir
pKajoIurf4VZuDzKZ9tUvYsKj4N1rjYBqECfSgtl0oE3XK3EdaIUg1scbfryD8aU
ss6AJksZPyoD3NLjNWa/zKM5fyH/YEHE7lJ4dKkMSCA=
`protect end_protected