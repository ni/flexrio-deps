`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 57664 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
3nVGb7niQ1PkM+U3ySg8eyyTqsY9Pr6fg0W+EC0fNJFfcQKCZi+WnS/tlBj5rxx1
b2iycSwgEvBB8Re2lvpQY9W9/iD/eMpzVcYujAh4tKO8uzyWPOI8zowFk+o4rQzg
azXtLPkgX6oe2nt4+JvaA6xAIux1sqrMljKgnFLgN4STIG61z7ekdf4T7Noh0TLW
AYAlmPeSeDgDwTxZmMVdqt7GsV1WoUBZZaBQA389BcUrufXXfmp8Llj90f65AYQM
quE7OGtnuTziIq2lfzyWbazt/F0XRW4XiI1Z2NF6HrhbskTf+GryUe/hoNVtLfvr
eDxB3POmnsRZ5gXHXLbih3GUSgP5eHVjr1SkB1Niua+VjDixPuLrj+a4cAGpJgO5
Bv4yeYHACJuIVW7w/rYcGk4MnX6iL8/DEej7UVLFKlJCXaH7ueAU3LH70Hm6fcW6
GWwl21P16IcJrore0H+v4A/Qiha/fKEsJZSCdyWxh2lEgwIdgMz4wdihiU/AZZvl
sxpaKRkeQ8g5DQJ9RBe6CleVlJSu+Pib2oJDXYHZSrYUZqA2qMxyidUo0D/M1VPT
M4MTWWhndEghZkQsPk5NtThpUXwnJ+JoV2lcM3/b1vu4cNG2BfoF+MpvwBOyDfwb
CEQnq5z7Lp6WpiPWlsBfwvPg0QqZAFgGHFF6rNbHoNoCcVGSpDOVtRWvXgtncmuX
o/3MJKrmCwXSvnJ9yoMwHnZv8/bOjVe6hOK9pzzMy+KFcCjTX3WN1TQDW2GfeDPU
sm1cY2B1Dv/JOpEKIlVCNVDBXje8ikwKnlOxjzByd0IH+8L2t2Zmnesb7FM0/NlN
C2Dzwmw3y3ue0SdxqYv5/xLBMpdZx4vn9nbr1pGBldVwOLr9uerTZ8X7khbcyUFW
Iz4PArG3/CCJLfMnPpzoyvPuXjef4q5ZiZaK9/EST5kF6R5y/V031Jq4xlKstk4y
nUamJnDeRJJqiHY+7xv7BgbZR61jrhcDx5xJ4OxVo787uFvj0rgRb7G+mHJIGPke
Hq3VqFpjJRQSoItbbNAgI7gtgS+Dr1KCOgpJ9jdIuuRmQsk8I8kDrpVncaLzfrNU
x1CcH+y6nMz+RSaUlenQrrSaq1BcPRzD7BUNgzvk+Y8tD8zZdH3RzIpqj7CVBkLO
AJjKoMXEVU1UPdHJdN2Rpw+sXPg2pariWxH7argiAv124G3q2hmPrfAohwbH0i+P
2LsgmmxyHIJNPiTG6CUPQf3eQQnLmRqjkYyejRcaBD35Y/tOnIfXe7iVxoeIYAZZ
4WBm9iv4vd/kaRb+rK8mdWVIyrUCNU8Bu8KbZG5fQZ3pv6PtHwAXzX1AlVcRX7oQ
thAVC0ltnoiUgi5/u5yBVoWHKDChvQdXUq4DQ+MyAjBH9oXUC5RugP9842KXzhIJ
iFYhQhjm84nLOOdAa7PVE/bagTOTIgU1bQN/vGNYX87aB9kLB24MWnpi7sK7GneU
hDFAPb/nicJ9vIyTRpOaiZDrcU746Nik+d4Ymr3lXF0O31dGgsisrlLPVv4U4cCQ
/FZ16lfSZ8Ov/aHks9ENX7Tq1awuhR5IwnLcxmRVAb4pL15UR5bJHa9F/4DL7xNp
0eje/o9rUUPSt9Gq9oOlBXsf7+lRfPVL40oV6rcl1JyLU6HCOCUPQsg0SsuuOSSS
h6ShHd2BSFrhU4+lcStNiLS3S11D9FnyJgFO97kULoXkWFAv1AwO04pF2Y8Am8pT
cUyWkmrDtxQJqYHn8kbYA355tVvChv+I8ZEkwZwLxPHjbzS1OsVCdHCeVgkSRxvZ
7/dKH1UNI/j/Y1sO11bedgwU8cPKwNN5y6xK/sLfECpb5iyeW0y6WSw3+sTp0lpa
Iua17U/h3FL4y/uTXF70YqcyVmklXOi+fxV4Em/1Iyj2EzcAAAwBCdy1ZXNoQ+MO
BHu5sQNSsgJgKyUKVL8RS8VPfUthFwZJkYrk2WLuTaYEfnnHOVLuGOv+dxe4mv4P
gqtWjacTD4zNeTYftbvxQAXCfc0wR0WS8zHfFEF937M+8qSqPla+8LGyQ/Y6Y5PI
rp/C9GB2t4Q4gwCWBR5rlkGK+8jh0x6wz7OVMyspp2bKftab6vDNz2l5UoHczYlx
fgDCNEL8rnJlycXhqQGtDA1P13aIbXFUzcYq/P4grrLqQjaDZwdjESRm9pTks1hZ
XD5rslAovmUyFXnCRBE30TmL/fNTFeJJxJRSvt+tMntDFVaDZClJMq9rl+tdTTn1
MCzqAjEn9ZQ3d7pfB5nE/Cg9hZoFUYZ4YgkqK+1PVHzedNXVT0Wq6zF3RM3L0zqN
JfqI9g3bql5r6oa7mFehqOUcMt1bTxXWZk5TYePN18u2v5U+IShZcXIHdNvG0ksK
ByYwQpW2wRHJcWWWFgPQhhNsn7iURHZ1J8oTQu05aChsCMgAuQS+NiKpBBarmPo/
XsqJLJn/4nsgZpQ1oq6O2dNWHuiXw62N2AhP//309eWHZET39MNeGkaG43CZgdfL
W8OQNK4rkxOjoE9RZmXzYRdKF6UBJg69EpddD4JeAp2xQ5qEOoZ6xv3WwDAVbPbG
MT0cQ6T8WLbU8yxYd0u2Rt5mvpo4nez1EoKI8wVcZoL3yReQQ5HJD0+A9tlmE39y
AGrHxfiXjHs0dgLDWCH8DnZ9QUPA8deeyjX1ggLOwN1Te4673y963rQ71GxtKyyq
61+3Kvgo/+hEqKh6/IWhpFgRxZJ3x3jrbbpfTR2C2m/+dzhd1tb5RkLuILv/zvun
gcuYjaqIQ4LSy7H2qjCit8zyyFW+7vIm1NJx7sDtGb4/X+Fg1T8VJeiB0tZPqo5E
bdaVaHgt8vcn8O7IKxaR4doza3TVLjztzZO0QlETR54vNdsjAiR2y6SytjtXRolu
v+j1f8tlTmqvMlURHxjKept/2B0ECzPgDObDF9q6JTdUUsI0VKD0KJW1vFvJqx+M
5OdjFJH8ltxTKBlLbLG6xsk9AqVqqdhIFLS69yxzX+2M3kf8l3o98Mg+RX5ym9g1
eGlxoKU9o/u1vpJSv+XAQBoZA+GE7isDEEochKQkdzQYkSHsdnZjVRXRTKRGcEbZ
0CqkQfZJlx1E+rcP2OQu5nw3BQEPHXQnomeJlsDdFwBljfBTRJREiPczIqzoBZeY
9jLDuMOpsBA0QU6tCgPC4Ze4YPE2jk5BUy1A25NH+SsR9+ogw61RFqLbLNdjIHU2
XQC9dFDLKeshrJRmQ2NegPGnIVRlqUGXr4cq9ooPv16DemiwddA2Lfy5pbSys87Q
rnAHY7f+yrs7Z9WgblffK3J7VAEhA2/oJoOfBO7ltAbgzVH4FWjDsXNr7NuwBkdu
0JncSsDWpzONXxlQ8EBayBowe7GIeW8aGmjf4Ev3OStfJSbiJK7VNIZWp+h2rk/I
FSOWevmquCClA9yN8KE0OPy+1MwFvrNnrisH4zfzpWgkZ/xjuvz9y+QoeblXoh/P
wtS3ShjuGCBrCwBYPkp90VFS9I8J4EF/05TLh+jaKaTe2OJL2i3GCCG/9LLi/veP
Fw3Mvh1PLtR5SGtOSGIdbRdL9gvjaElk2pkm5WWcxcUqlIVWi8hToei3VxV9ioyg
p/p8u+TjmXJfaqzyf8nYKJ/x9M361EazEsqxe3R7eteaeDJWqlRb/cOvA36/AnYH
KjjVlvPFH4vOl0LLBfkBSArPcJ2UoMQBuNZmGBWd0gV4KJimzMX6CFfC/E+ENWIC
ZbRjz1yGpe7hUENcVMm3tQRTdLyZGLJlCGWekBQpb3+NdCjpsx4WmnBTYxH0xoQc
Tkmm6d5VEd6ARaTiWmIFJ2+cXjtZV2mjIvvcpQL5FcT97EuBKUfdD+U1GwEAgEx8
ygee9zYNYMQg/yDG65Fo5VmbDegeDGNSjvhLj5IcsHtcspETRes/10hLG5s+2O1Y
yZXX9RUiJ+Vc9S+rCPV39x7AL9CjIunGfhuTkJZhYhQ+qgfz+cfJ8LyKTWa3oabH
V7cFrm1SEQuO6rQih6Q6xDs0XkQHgF8NngFWjpVFfUELok8Sq5lSuATyYUfoZTyj
7ohp7wlbmOfwfZfmgqPbRAgoHKbWGBJxE2d8vlBpoiTr4AFLf/iM9Oy6ArEGywJk
v2cjA/5FPkyBWy6AoG7AHc6XCEKVw5TL2jwelvNYG8ec7cx8XD7lDxKXBajlI6Ci
+iT1HYhVlbsxd5t9U//N5LU4gzquPfuDrPGZLASD0cyIul0qHbXNO1M1fp6P8d71
9aAk3G9PYtAsD5l1M5oww7JK1YnC4mjq9O/M4um760B677ajXGUg+0N2OCcJJ0ZU
g0snvATrphkyRXj5kphqbeT3HVmlyIdq8Qiwsr9WKhLgzZHpMngWfZzpuRiAgihH
ZIHEbq5LoPwoxFIG5qE+yth+wKC2halMQmHsbqIqobdPDxgpnhYtOVafhK04M4vI
KvKUIYs82mzY2lu59ctbJRf/E4sUTTNZke3oiyeo1LXYVgR/SbU829A9A5xRe/7R
ioXYamKb1q/BIQD2AItvE7OE9hjcIZynIMxbfZvLrPT+oEM+EU4M9Z4+2tzOzROC
ndYqCJXp/+cu2huZ3lztpt0eNRrdWm3vxjgwz1iFajBZ3+G9lE7B6MZ6H4PEYeOX
GyKibGDH97VwICJCpGDvLa/aPiP83N8jNyKyH83Yb5Fs9W9ktZDNfA/cOra6MK4e
GhRpAmZ6d5WFvIOjRg0HFTfbNACnYtOs1pJjI5lAdejKUT2YtZRDeQaMK58wSU8G
wbNVS+1SnDT5wzG/EPkoJ4QcM7h51i94ud7IYuQqZjhjoV1UE6wyw/GcqMuvG37g
2BJNNdTvGHQBkhtik95rTZKH6xp1tjBsPL6bdwfBJiPuPIomK9/jzwLYgNZeT0N9
sxjnwnSxhptptSRPWVm98VaMmgrTfq0QfsuNySrBDHLqEhqvjTTfi2c1LYTYwdlF
fAuZUdotrwhrEKTxZB/l45H6Z8tARMqJh9pmNGlxviOFkmBrXOdwv75bHwyeX7lI
vz8GyTc/ETG5H3VeYGlx98v36rS7wCC5Ph4gieiTap4ce5zXhgextyENWEFz5wK+
DLURywpKKRlAphabYgjJJS/ovBXH+UdHbJMm7uxvlSpt3yVvNWvkVODoTzFSZh1f
wT+2xj00IQAenaMCX4KfJclc6JmjgVeFI2hExU1YG3QBzaD0TX4alNOh/3EwR26q
NI2+CQJ3ahOM6n6Tzi426N9O0W+CU6cuzdCj7afUqzEMO7t9Z/9JqMfNYH/XosqL
P27MeitZvDl8napeIXO8TA4vWCk0fDuESldWbAyYASA7Pa0kHNdT4vMspMfN21XP
fCBQtVUFAv3KFle1rQIJ7V6jVhFWEAUzAZHPr7j3/PRqIJ5AC0e4Iz237HvwGbD2
BnOBTaXnbACfGGvSBxn2SAyXN30ezmbiibiuYlwnqwNrlGGhNpW2UJQoEt+Fms44
liLYMrQqBn3ZLULe4s2+hvB6YC+5v9TAClKvjYKM6WbU6nuWzSTwUHRcyF1g8C8B
ohzeABhqGJwn2fyZ1CSQbADrR+lZVtehbfGkg+RTmwTd/tqE3WwUURydkz2+HSHh
ycqUKuGA2JqJfdCIDwDFCItelrqnLzkkTYcrgOA1yW7RFBWndC1gZBWm3Hg7K5fZ
yyGMEhnxCViLxfQMAvYdXPyCS3a6GOB6f9sGmJPk2GYgrbf1VzcSNchu9WNKQisA
JFqXdv/1SXc0fQiPKluUANMqflpHmMGKBHRG5z127Xz4bvN67Tt9giiacl0rNySB
oJvnHShF3uvexQyHWFYKDFqglcq0No1T4913TZEUDtkG4Sv/N2Pl1KwUI0WlZMwS
IZVSgTC6lf3EkMTdUfYYTyK0pou0Yz7R5cFSSxgDEgYYfK5U/pcRNabseT1Plv+w
EzMZJkPOOJJDaPKg7xmaPhRjxmNIKbOQuLaJVCJ5FtBbSP26SKyfI6AWvzJX/Abj
2KtQLMKWeGRGgaq05Y+iooTcnqNr0QjquiX3vsiqqe7pIcOf7ARhNfbKJ4seqqyO
RwdzIchiEUPUvvvZentDWEj2aXf1ZxFANFOi3siGuOPdMJlPBJCAgB9TWIIyeueP
ELVweKHRowdCU1jCFbu3A22S84W6Gsv+0pPDw2Pp/UtR1F5KVZ2EQq3vQUHNJLJA
1dnUBPeaBjh9EF/e6ssFzMtH2WhSH6LnuT8AjU3KH9+yfd81ruWVqW2bkHMKUn9G
p84A/kNg8pk0MXoXfRkAXMGDj6r6dFPQrqC8DqbaMlIWvGmB7b+jf3ZWTcmd7mtj
dSapt807QlQRt9079CGcIUXevFPvkszH/RnrV2yJ9qQLPkV9K743psdgMVviS6M6
KHD4YvWI21uEHkrms0DixAQcFytOL27HU6Pcg09JtPMKtGOp1UaCt+Ufvk5kIJ7O
x1xVitx3GPczTDbmFEvIIFRgBFtShYezslwtZlEzWuIQib3w3BmsmmNIyZ8g1/QQ
fnkAY2+Ji4Bp5q/Jgo4Z/eNhV4BmhdmEpCWNq62Y73QsIjrb1BpOamUGJMEjaQeh
BT7no1n6gBpzmhHflBIEArTnrNA5YhWXIinubx5ElWInhlxkGE1YSwEZUVnCnICg
VA5QUk5sy2zV6ob+aXyHqD1f7Td1W+inNohKKg5fPLzaVl20TBoX1ZZuUdPIK4S0
hxaL1SGSciG0+NvJbXuqR0I96L3afcOMl3FMvikF/ZIHHA5hhR1dd0EvYrieor/z
iEv7i78NCeRhWosE9cwbPimXn12BMvJeE7ciAfK1uKWXVeetQaZg/UbyTR5x/Etp
95i1wJaZNDTzwLDAT4KurElShdcjSgCg8uQBMu6K0MjGse5Am2TjE9m3x+1xX0G7
ybf4xHRbSu2Mc+C5k6hMJrwx3iDDI17UTTWb/EvngHR502n8UGZsJCMd/Gr/VUTZ
oXNcu7D7a2x/K0eMvMcOqvaec4rW89sMh4YASCnhd0351KDbcar/YGjUSqKNfERY
7KSmp3rN7XWbJ8lXggzC3CCuLWMbj6y6o4F/MpV6niv7wkO5oc4Zy89ZBJXZLdYn
fb25Tvk7cNKaqTEuE0CGyvUvD5JmFYINlwmrU7xuK6quxlq31ZCrNQ4XyENqt9oN
DxZY0Th+pwc8ZlWIpByYW4tAsJGoODliZCRkcet1S/oJBnRrbs3tGVSXYACQvySl
zEY6EeB6tFjxVRUSzP8bbsiOuO5QP0gLXxltsj4OACxL0P/+nh6xgCQti09kpk5x
Sebxms1Cvc63/hQIm/UFGj6D4C8MWEM+T9LaXKMKnSQoHe31XoxlIwnrxuF2lEuo
NtuTo02bHPtoYsJvNXrCnMz7Vsq1v1VW1FEHlHF7MAqWXpOohN2e8HY+EkuUB5XX
mDtRYV3E9cVYW2CiDcgB6IPONk3rSEWn6dX9D0CzEcpCsr5fpYRIWzrTwsvmgW1I
XRt5fBIxasoQBRuWtE7Sk9sKJHksGUp2PCa9x3FZa5GT6JtairYkPQdVbg0qfBlB
FHnT3AHYPsTU3XwN0o9GnZEsdm+O6k95Uulgcyc2nQ9B4RweU5SJ7JlGLfKSpUUL
5mfCVLttu/vFbt+TJjrHLwt0jNrJo7uQMQuTXGNB6HFvFSqkv0/nQFNai7JvnwMo
qu5jsMir9ZZ2eA7wLQhwbl/ZxltxQ7pGf+u0VtVL0phjmztON8H27uDbeA50pol7
XPcb23cj3fmBC7vrpFgusp6fl7tMCcxl0rchtzegpoLfkYoYEU8NxNKqc02qECal
DS3MnAVggEjNv5yHdLCOgmgjHDr+I4aLIpXQuKFKauhf8XPVxgZexT+Ryne5g8Rd
jKkVplcQKZENU6bH055GgnDPsqBGL5iQkhqKKVYWRz8Bvfpxgt7e1c32brpCCp8M
OPBLIQdzi7XlZ1Dfi7SDxpocRRZgM+MkGkXt3Co1yibkAPRfIxlHPImxMAfjhz9I
yNQX3XeH2bsR97YeGKOCzuTymJsZRrNA7GuahQfmyEWh0Q+8AKw7oEG3/3r/4rJC
Xg3q6NvMIBGExmJu8aBVjwYJrdEe93fOeuhQC91oRNmMmGGxLmUtqNEZAbmI+I24
gywcSDQJ5eHW60EtH4s3E08k3m2dmuxIMtWIyUnYqmJ9bZnmamoVG+c/c2Yi658y
mI5LeUhblQ9FE5EK61ZlM+S5AanYM+HgEnfSukDRuXOOzaT2d4dQis72RacB/7Wa
/HMzMyMWf2tw+0TDWpLhjORxy/twk7T4C+Zc2sZ+O1TwJvbecj8CugHH/mf8MmVN
HJJ/+RszZABcQ7GKpSCy0PW35IntTYFrsD/mLV1WLAqmOLE2OJ9fXqDL/AyNZSzc
VlkrFfal2HDp9qdYeWFciAJOi4k1QwZQu9wZaByLyjwzbG1bexH/F1Dr7ZCv5LPs
EAoTjZbws6wd+qyPYZFi30pgR7Q1uWxCFdW7O/t6zF/K58Zt4PkqVPLosxeUaALn
JpYofVNPFT4gy9vRxSaxKUaULUITgqGVQc5WHUgRugi2dm3+HC5UMHiJwdFSyJ9L
pOw+XX2Tgxmqc/F4jAu7sv54y4WPpD5/lwQOydTg4Z607qWeKRC59wyPYtwA8S+7
ZeFlyPzCDDz1S7JOxvgwFEEyAk3Rr8cIgR/bW9QI3w3n8QxVymFIrcM9C+vJFl7Q
og/bpLYb8ePJVL405SFXev8nRQQTD6Ia/z51RVrFVf28KOInmxFEiIz8pbGRVU89
6xL/vR/Q5SZqgBUCyk96wL24J3652vpLftWZiWLsCE159uGHTX3mMIr0v1BPg1Hz
ShIVqy/BNVuFn85Bf8veDmqQoNHJ533OmTdFg2lfVV2ad1MI8NDe5u2GpBDDeX6g
3/GbJ8OUeabfeLQrDoZNJNSxCWjKSYinm/orHKE4wXGwsBWazE2Ii0JnKbUjxj0n
8jrr+P4JGJGgoZpK/YztyLFWvOAvfU5o7I9eQQSI2rfe5AIcVYw5Tdut6szHKLFt
POCuwybaBi6lhJo9FRyKluMZoslNovQznhmXwfrTmsVZsNOQFsJ+y1dxQv31X3p4
usAHQGWizhmaURz5LdmoVtJdkFJqOq3FeRPU+DDk5lJ3s3tcyCVhEJ6rd5h+FoRN
2KNb8qUuNPjmYyqUedM/LRr6sW0O7rYz+GTQjvDilgTuhfB/CWqXu4K0BEMmy0b5
G/cTg9+DamQum5qFOT7u1MpAj19nOzJyLZHQ5bso//Aj++DG3zo6N+nleDx9xiNr
r/cRD0dUSvrdNyrwHOsHm6OzzLR7gUq7ZpjydWW4BJgbzMiXnYd0M7mBE5mM4HNx
8UQiT3PWLBUPut6CPPNSo6gkV/cn77jzcBrLqAake1u2r/fW9dcrFT7jXGsjQmVD
BuOXsb81rDdBTU1dyVxPlTW8ax/8L1lg1QHWF0crE78rd9PXG6msYimgIaQCBo7v
E+PrhMAcCCMjccNoGh9ExgmSS9skyJ1f6kbLRzTgzPbgykgGB9ZPpiyDAxQZ396t
DYMK/mGjK0iNVkBC6X3oc+cKP8cFMQ4rk4Tclii+Bpzai/iRMQZJiphbJIDqphT/
YdcqG7GQx7uPrv2tnQVa0lgIerlVLLg6rXa/BHuXEw2Y/66hFTpGJYpABeubQF8W
tlWP1ougUSsr7BBF5GC3cbYSOVBarlEojCV83x7dW6ibXPSA2S4d1aMbkr2QpG3I
hAyA6SoMYWmIRGtj6hm1JAtHCulsuu1tfHtf12vEIku5pnTtJTHDwfXNjyUFIbnu
jAkq8B6pFIpmMMx+lvh73yApxL1otokwV99NwuVLuu/Z7FBmiogyWp0bwVUU6SQo
+RKAZKY8CqwbYUELwFcRDBrNNXMeAAqng7RT5VfEQyXgqXgSZNDtk4+PcAZuRV5e
JYpHIBqZcR58m/FeUSwkxLNekKmoadXYdHOKEBz+6TRhVS1Vv8o/l7815ILEPoSu
5LzeJdNdL8RMgRcuz8YLSmEEJIkPznHG+qC/zE/f82/sO13oXLlPG5HA8gbRCm8U
9cfyMAiewK8TwgljsTBl93jR29eIF0K+4swFzk9uWuCynPezi7/8cUtmhix/D8gq
CxHlVHAKD+Vwz5PZkpLFk79fM6bABcS/Qrtr3TlWBOILZoZqOadYQYW2oGXbpM/v
W93IOTXRtwdKeUv7yKW73orz35+xmsd8WZsyN8uAK6Jm7BL8dyL1rRAhRjtZgqsW
bpU01DXPi/leFKp7h/10uhg+4hZYPnnkpQPDixXH24RA/eY8hYYG48SziO4kncyN
lH4oubiKqIrOkI8CbFEediPveROSMAvKn48iFqam6k95h9y6zk81ApIkYMF303Ae
mSupofCAgsbnwHP0uEs227ceY5Rc8hS/HVTHXgO0L6OuYAwzAHKqxRq7K0qwxhlV
dn9bqEfg9Xg4tW+9322YoyPkACPX/CZntD0nAKD6nY02CVeJ4VL4rfrBtfQsKmfe
97Vd6RH6K+aTmYNbMntGMfsscr3FxUE8mYBTKbeSKBZX4p8BNTVcETmQB5/MjdIu
nXcmg6UmjF081uE9qp5uiWgdWqWS4pkOHNhEonrk8IdB8K+TiK3CWGKnTtXSkysy
UeWlt9JUM1E91NzV5w1jfjU2Pq5xoS3T2CubB6ff/zDHyDUVDNu+5ToICO90XtIW
GGeejB5S14qBetXq3t3Tv7zL3OafuuI6WBS6btVgy12Z6cgllIC1arlsN00xGYs4
cDwbF0isdRSnkB7hub6Wk9ulcR4iAakF6bNvK9WCoqfdwaBtD7jQL2fMZYRVr0HH
5wunhuKBteiyyphJoQppNMOwAA/Wy37ho8zt63MixeY72DeowEGljwlbOI6huA2d
LFPHWrgGngNF/963u1rDdCxzMxgwL6ovQRaQYzvMIBT6CtREV2jSp6dORdN9shAx
1FdBLXW70Y7adxKLg6Yct2f09If/c2MB7MVNbyCKdYC1BW3a/6XSe4oGdMByotWg
5R3JhcwSSIN9rXfjxJU1GzN3bIN2ndKJ/+OggxCV9lACtQoCUBasR95S/irDKiwR
41h+AcJkxwrsLdntfcrATKIghV8A8Vv/6mZ3gXZpy1fGYmz/gNMLxEqr1dz2aTUW
HnhZofLDUAHWCwbsCtovMr0PkeXJIuRHWIBnPGCF9eP7cZTmjGyjKCNhfp7x1x7z
fI+9oJYvx2FTRqpBcxk3rYPLi+NEiwyCAxdDX98EK17HhRrDcpeIh4Z5drwcdTJc
YKWBsfqS3D3GJGwHIO2Oc5ZptSWVwEkl0F9AjXJbT4CtV5ry5gcv6METGcUULli7
rET40Q41+tn+ueNEzVXY3GrgbRuhexi4QfDCys/V4pAtUBOWGQ/bDeuqHnzFB4Ns
r1Oool6Dh7FGaFo26cz+g6YNwpMjxd7yF4eWxKi8dGRedeeY6YZl7HXuWrFrgfoh
TDkZinG7uxuxa7TqLRyktyvCXg9X/3IAd1Cv9rXQzd3BtxkLKimWg81dwSSXD7iZ
tmqs07+mO2pJllKrdTYdDTM7Ti851VQbbTUg2APCm52GZta/X405ABkvA2ddVDLv
hnYy03+fL2AAdTKHWhNodtzMDFkujm5wv4CyqhOTSQCPH8D1+4x66VPmR9chp/Yg
jPvQSKo/Edx331wikstAV44yG2Gq3o51Sk7qd5D54iDMMhz+iftmFxLQLQQSBRhf
Xj+mncCgut4f6EoGjfbuf3YdJyz5vj7VMan5dfY/NDv8BZvaRA23QN02R3l3sCJQ
v8lB6aSQDBMMhwxx3t6ufnGxBiITWUHiEs9wNUo1BaB+kp4yArpJZMdNg2whnNdo
/iLjDBUhYBcVGce5O9fNxaX2I6kkCAPRVFzClkvCuJNsGaTD3aCSEOPZRThYM7vZ
4kKCy/klEbe+06rS3f9xNRzKw/ZBxDGcLEbwAKSk1bxx8jo461UBedyye6CazIFo
dtJamjPfbKTynwpJcgFm6kaPHK2I7uienh/+JVd+/35phik4T9veCwkYFsQ+u6OZ
TNxgIGDQKHJc5LdcysX2zBzfJ7ODgGInae0cQ/+nbC+oazSyLyebazr+s5viUqXT
+ewP6N+F8YYT04rx+Kb4Jx0bCHGUPaiFrGGWDURW9hzHgb2eDdr3IHkh7RFVi0H5
Y24GUbK4MyLTz2L4bVCcwNVGu8WH2bUo+YyqlWAagl/xda3xQznKBuKhyr9Q6mjz
pUF14wWbyW4PcVl7ARithxHSeQukzYxyKFYSvwhlyNmXyXUsmszQZnSsahoHhZKY
ig6pTecXUDZOIT8tCURaRuvJBSgZ5Duh5ONlZ0hgizxkLnBU1Mjr7aHfpNYevOBv
eY9Nk0UCVbiGG2LhFZogEwBHdm5eJvs2WZd/TdY4JG72ODIAfZRI1hXSx4UJ1XBb
Z5V6RWTG2OaLPewsNsrtnT12tXwXVLVVyGCSDrDRMVaH+SpCOOqA5N8a5z9wV8sA
YwI5/ZifCPfHdxtDy2Z0+2EwMBUrhzdFBEwnx63IsBqOTX5S71/6JmYv7cOkdJT7
NwS/SjwjOTSru5eUasJPYb/8IsLNm47gThR5+eWYc9D7LP9cLNeMy0qz/y7WtVV0
W0MPZbdTEoEjM8k+k36vQAIVcj/KoIqzXB8nFT7ajjv3E0zQb1yzwUC83WSjSEv0
sMCoFximG3z4lxAq+/RtMiKD5KQyjxV/hfNNk8w55BXb0ah0sSJF/pfF59marwNa
qG1BTzLN8ZDlq4noCsI+o5oDwIUGo2y5tHtIBwj58hEVJmWHbXlr6VI/WInizata
THvKhSZ6pjYhe7oUsylWM96upBUy8Rs5aJjEKEDn+2KHgYSzMSAoByp+sU/L9mPy
xO7GUMwuNbpue+KaOmnJQ65JuVox5YcGVom0tTkScI/KwtlaMrKd5p3Awgd0JV51
29o1avOjUJqhtuldGtQxe7MeFpwwmXS7Hr/tqcCMIsP9FMMpZH9rVroLZ6LDoZff
Vw0C9avvth7DCMVvnLTrvaeml1KS6jqbutpCo5UHzxrjLZ8HogXG5DF8tYA1p1mH
Ylafgiij5BQNvp69bpCqCl4e7i/iU6n9X0DYOtNUn6sL7ilHou9UpX/YL+mN+J6y
4gX5xiA0wJ09Bgsuc4Ege+5iMcH//RrPEWSHYGlK2Mlw84lPRWpt6h4H3t2jDXwz
iA57SIuXmeZPmnwaVuzl/F+MRVTGmoVbNVSy3P7hQhIZbNGm2tLSOiCDpbzx821L
S5lxMV7nI/nQp98RgFSoUGAgiBdMqg3748PLou45SdEYJMZ+ovwlYSf16LrqqD+M
Q88mpXS3MS/mkhKEvNGjcORotYjRLu1JaWruNKPtrNPSwXqOxXlJtJbe3e+ce2NX
gycAAv9JLVNwA8KxX55lgUyp0XY6rJ97BjIsP6dwYMYLNW5VtZ/McBvyS1G3bbs6
jC8f8ByqAaWTSU+GHhpIwGQx5DAeK5IH6EOIQEe7LtZoP37KVg2Ef3Tp5bfSh8Sk
VYe1JZdie00c2loa8CURcRNuZ+WBMLQrokbmppS2mofoaTlH9PZ8jRRiKhjg/YP0
cidowrhY2Aa31lBzxg4q8bjyfyKzNyUEfvjdjMuSOPk0gPA2FGfoIuChs+u/q2j4
DZTu1M3luLsygFWQ/80DXjWPfTb6kf8WfB9GKu6qO7jr+LG+kLlKc4+WuN44Fqzl
J109cACaoeErvM37Y+j6hRi04UhUJACwa6Mv3v3QJ5Ip3EbjkY1akaGodsy3PGxG
GUtSNolAdBgnkoH6GCOaedzSeftD4WEaG7u3hz3JGFO0OZ1MzXy/UlDKxnVzaQ6j
DFyLZr1eQ9m1hxTHTQuiSJd4taBFrVpdEeDVkUGCMH93ZTLB8gN4+EwtlcTphTsy
vhRExhmMjcMTcr6wMBPUqAkeRdxDYpsq3+OMPid+MUpncO9hISF2dPQJq41vQxDo
ahcDZ1cnZrLsFc1s+6lLyL4m8ZJ2ecrwKpR/ooddK1z4tP3tqwdw8uMzL1YLEgrm
xBlX4Svugt0B0//CYG8IwcLKxZ4TAeby6myIe5kEflpdM/S9Fd+S1gK75GIA8t0r
JJIX2+2A9rTP7HtVNCBWHME7nZeQs45w8WKLqWz4eQQcNIXdklsQDr1aNIFja1HB
MYkInmJGrTNJ9iRS2+AfoQvtp2EG3O6C81uM/JfhBo4oW+lcRFELgYBrBu4Vjr0Z
+JMDoZWuzCxoZeTUh3/FRqTFEhkyQaG1FKM/QmbdWPncBKFCdvIurlfGqu65g7HV
5u6iUvdkJfNm4naWtk1/Diy2Ej9eaHveK+H/hsh0JQyMEdJ1TSrmSSkjvasi5XRR
NlGuKDhh1lMuKo3m59+MKCZq8V1qzS092IL++I76EMvTKKUHUbUwG9B2r3Mk0GwA
Zqd4OhpiY1KYeqSkVHwKsDlZGTTLu5XzuCiAdNltoBRLsjLjB91qfeqj/yuC830t
EKgMkRLmVsalD28tffzZtGNRFSUFi/+/ESrG97aa5kOdqbf6G8KjUm0LGvBNGl65
fqhrENMW8o0JZzvc1MpawteF1vd8t6lDlZnKARblK1FZ8MWSwCBzKa9WHiKO8vD0
/dDNU5vYTTpwr9iTOIakBkM+GzFikDbcDLtDu6vrY1TNScbvNzveOyStDAwqpCi2
HsBPmCgzSda7puM/y9dZTOfpnC6k9QP52ZmlchxOUu2AwrL83Tj5u5XNQl00rL+u
E+Qe45Ru6dau1SMOiAYogODuRHExBvi/xUTPJNBCVheGXziZ5O5s0nbBWOuyokSy
Lo/VWC6A0FrOXRXlCtWs3R76ratpxvSa8GgGM49ZmItUB49CXPeZ0dmderqb7w8N
n+c6o+pvhw173ze+/h7Uv19gDZj1Un/mKDvunsU/D7wlhxZpeOER3GLkt3A5PH5j
VJ6sGTDxcinoaEhbBc4/5tVb9xX2O8jWyAtlpHLU1xmyv3eGuMJGT5YIuEbfTAq2
G0bf51RMqU0sFQdF5v7win+xxkYGDLlW36BJ4esfX6evPzrfh6nf6vno5rVutx7E
1VvA67oGZGhvo1yUtPdijOkMR6grQhssAzDl7y56IjQJDJ0crE37HyQ7KdycFQaa
/2BqiSkbsltmMadfI2mtCAmMhEl6nLBTucQF8FqKJMrTELQQT74i3/Ci4YgVUN7m
N5rrC+z5Z6V7WWFoMxMJ22hx2PFW1yWbds4ARiEcNKppZ5XhkyI6L+W78CoywdvR
zF7dNG6ErlXe/MXMCGG0Tpsg41kQM5bDbLFqe8rxoKc2RlfGpI5iMS++gaKkhs0l
3rg26zlebRwtHmRa5WUFmkMcmfCUxgAPGtX0q6nlK9FV2BlXcPZe81DUj0oNVIaF
oGX57qr9lG8wgtgiwYqBjz4oP36qiaiUkWO1nVnoQ7aurqklFWVUlsXVEoHKL8DT
gYjNUzzL5+hR2pXBGQ/GDlDCxc/2KFYpZ7ZbQqfspO/4Kp5k84vWSiCjbES1/fj5
Gr8GyN/1NmYpdaYk7xMgJFqfooBG8NW5rDAk+su1R0nxQKhssCTzzJKBcChBwg5j
NgW3uNHEIQI2J3trQcEq9iIZepCcwCRtfvHFAzmgsE5bq/Qsst2l9quiaewiuye9
MbgQJyPC64Ed0Wh05s78Oe8UWXjr8Ou9m4LTSSUhKIDF0DiQ7nDsJDViPT1m4oFi
G0T8V41duyBmLHosT2wJBGRgtc9JR6Ig4/YQgOyc3W6hTZMCvM7WkyUYzJsG92Uv
fj8ODl7hLQK4jhCswa1teZV7XG7sk2iYtL8ywlOqcLSDVnB44VqvVcniQxAgCIw7
qfHUi3lxKsjWsWdmapMAJKMQoinBvH4sbV6sL3LWFnOQHIyQQsaNgmDZd3QRFI1n
Y+NgFIFqzSitvduSSLXdT9SXlFuwtdEh32OR82XZTgBinCMB8DRuP0CAqU94yXto
UjSZ5IAhG6SCpY3O8ELvhmRS+8SDp+47+MbPeagXOY7W3QhdqCH5QX7F64Amw/DY
ZaY9ly4m3dITFC/o2mR8jeuhLsclge+JLn7E68NSfSdbXynAbSfX9OI2mjznK9CR
AJi7UDnAcRaaAlrHLtzJ/nTKz3sRGDd+qYKybIYdEm7FK23qjyULab+qf7RLUbi3
99HVG0J3lAZ0Y95+7LYSnL4zRm+V5vSrCEKfh9G5JwhBYWHG7BizqarOy7Z6v1+d
FfX7Js8Aena14fYQIylCZCSxm2h42fNROBvjTr8i62Vwn07VZanGTaJJimlpAWTm
id+cO4hACFvjAKYNdJK7DxIVuJ2h1an8xevkK8c+SfuuxTRNuyZML/2cJzv1D0u2
tVIjft8vAN68uIpx5FnnFvtstvoxCQwb8kJZJbtqoKS2zSM9tRitljYT2OmTGM6U
pefKQcv+yszefarnnwl42Q5ld5fHfsUKYGvCDNe5CAVOYASvcz0eCSdncGAMs6cO
B0LSbE540VsfGzAb+Gj3gzkqPIS0jexsm8qbOnotBcIW+BU1SucqPassaeuWhDLH
stoXCbs8U+8f8cCF2HvkNrHICzEtVrXwjXhkC3CIzNqYF6HjI+6GooYtQz+I4xR/
BOIfocNEo2rRVyqlUFEmIEGb50E7xNasTPOfjFvOCSAqSXeoFJvoU56jM4Vies0O
CfLv6tDLSqq6i1TCPUe5G60RX2+CiV0BFPNFEwNs6tKrcMr2h6TpvqpcfEll3hKO
HGRg4EOfuTyfP1y7MfsUP24wA+DXvQBdTO1BnoDpcJG9uHyBRMMCnvH4CRU2TtQk
QgEnVR+32c8Ez6NGvpFWyAMARb9bEvqwIUxEcnBvrD8lLXGqmeA+LX8eEGeGdChl
ZfCbrfP2oFwOfentDj6hfJG+/DISyJwRwWr3ozXWINC/lVR8c2zgV0Bn7aUZDnr9
w5U2QbFuAFxH1HTLo7IAjqxjINkx1XvEmmXOgJphQvDBC8CJ5PArGoXN/j8N7G4F
GDX5t87s17cimdQj3k1dq90VGu6H2HolCLBYOLi/Aa+BsUo3bxwIlZOI4k7U6CeD
B4qJ/yhvq2/XG4MGw47nxsRFz/wpjDGoEJYtjrLfJWu789a+lubRbGYvMT05SABD
jdZqc1CY2z1DkuxG9RJHv3WF5AO5nlDQqRIX7lGbXgFznwhxTQhRG4K1AqyhIOrS
VDUjRUEokqyUMvZ/H5LpHw35EK6F+/uFAwJK05Ntu3KGmGw/8IWc2oWzB51rKr4b
ygcmFQR2zfCJKBqcDdf8zobc3QxAuy4Xz7umtqeZkZK98pFi313TMbhpY/nAErpy
UMDFqaM0/fJdOOda5BrpXYzLHGEVye4mQ+SIxZcZDQDex4W4hO9XzCEeIZ1F1d/M
YfF6J3uXMIRfVD59yu8QH7ZS/tc/QwI+uwUt1fYF0RmaMYwktZK32vLTIkIsj1zH
83+BYe+Y0JEvTrP3rBOJbtW+gj8o9ebV0g2dlx0GI8l0RkjeNLchGDYSa45VtRvG
sLPxa2VoAOhEfvARi4E1J8YnhOwaMKaprZzS/ctM49pFpbdvb5exhBMcoXlXiBFa
DnrARJ6x4Z+2ZsBn0b9f3kAEmUYYf5SHAkZnThiXHiKRJ1Z8n3Av9TQ8/0Y2U08p
xWGUXOMwNEgmgKCU6j9Z9DgO1u5QTEjEWj1N65dNj8nPE/3RCXt5dZR2wd8V2wvn
SWI9LEtsmHSHzuti/SUs9rMaGC4zg1QMqBsWKmKLO/W32UAHIpE558snGcZqap5E
o/HToJ9Cyhj14mHlNcARtfnvxhtMOuBmj6OsZIE/gzlKSSlN+vK+y8+ttcpMloT8
LVxNrD3PvNgd/mibEaihiL4BuS74/8AyYKaACVRHIyGrp4m8hDHaI1a+sEInNrhN
YEc68LTVs2wAh16EAwgwfs/wjBQSmcLF+Ww+kS4F67jyzq9uaMgVBp7EKhsZdHSP
HVgFdiW5tUHC2CnaXGfWXJO/AlM1gGFu37S+ECdRiw2QXMTe26RLoLZSLELGfhiv
NQL0YWF0B/TwYXQ5+HMhYrvJ2r8tf176bGlt26AjImyNIQ0DCWJmilfaJ2GlS4q/
73zS7AOYff29ZcB699lw92xPijcLoe+/J1aND45G/5vkQSixw4X/ty/b65xx1IxK
qPg/Lv3SjQmgvIR7tPc0W5csjXWyEXAfluSjkfIAVT8s/fkZqpdJfTru59nTBFSz
BM7pXSDecClnq+2/OALQrxuzifIKmUF9lnjmkFQHo4fXNnDneVW/7LUTsFKxEGqg
i4tNxHZIj3FSkjYOw4h/r9ECR3rHwZ6gdNYWnAd6NPb4KiZ9iqdI5xqj4w+e37Z0
H1kGoLLuF+//9pQ2ki8/8DOlm3xjSXvYruvHUzU5De16emAvwfRCxrU8+lf1gOlQ
IPU3yC/vWJyCzU/C50BBG6ffA5+/+ZHv7XI4sGkXLqQIqq44/+Pf8ZFJzjR9asgW
Aygrnj12YlP+rfcqrkweZqPX2bPCl0aNX7wTCot/E0p5emxRpW2xqIiXrrpzfVj6
sAkkltv4e4A2nlZi9ssNDtcTJweTL1EYKZ1s+xiQ+n2YJE4pUOw3mLKUoS/Hv5IL
227Q2j+wnZTZM+fV7qfcxBs4nye/cVBMoKBOH79a/0CcGGlWBLdDQJBY8qZSCsie
7J6qLtqH8zIFB7L5rM7V/Zby4lT8I6qjL1WUo5cfZn3M83gF+VDXaVT26xUMi9kY
0HmWRlCv5HF0ALlkiWEZBDOU3xj5rSi8vHRk27Cf11HOHRsA/a18HcECbk2tXFvw
9hYA80xvTDK93Dv9u/yJ1BALgiyx+SuNHGNuMhaz0ODDioXb6RkiyfEMQ2eN13Os
ajL5vxjHFe7TCwCk23S/R40wNyrxgFLgCshoChgp3fL03a4mJJqH2rmZs+7jFjW7
8idHarRLHyf6FvGGyjscCRMQ8IrzhAbYn+F3LMaXB17kdVqH9Y95F09BMweT3Tbp
IuSyF/qGIZcPY7wgy7sHlg8fDk6ukl0B0t7xH3uzudTmlVVTxKCiBx592inNpso4
TmM8M1SoKHHDaI3dsC4qRBxbK22tdJTdlsgo4h5CnREdvD1VY3Wn2b2yHd+JgTmD
nVskAzR5qqo/CDWLki4qiOrYGx5XXtXzaLwNefoXbunGotfq+OJ/Y8kHZKRZvqx2
ugIVRKVp01cDzW/65uE+WybKCGzgEYEBVDNCTLKcHPNjjgcuXiMF3GlQWbC8T8jN
3JN1dUQuhPmsFuhe1g4+EGmeaSNXZ1MH/cKYIUPhXuHguzFsJcZ12xoQTisN90G9
v23dsTZehfOy/Lg39lFjjYD5BkuKmdaJcYhTVrgwjb8SMoWnD8dP5EWRFcIYw3bj
YLZCPY3ZZn5yUcAzOVjx1jyt7INEURLU9JIKj5LRzLMzwEeHgwo2gKx5SYHSstoi
Fj2WiiSpCefdFRJR0xEsL/LovO8w9Z5s5+/GSNJsx27Yi1tw4sEEuYtP+J51onxU
uiKlOH29+o50V17nNw890NRljXZWpM9hCA0/lxO99UtUoBy9mQgXCX35sK1DjUFR
6K+O+/B4nnTcU81vMCVG3ASTsZijSiR/xSJaiqwVmeYhv4nyHKO1Rtw3IlxqijIL
I9jDnMwxJr6G4jKitTElIltbK/RNCWNT7Ww6tKiHNiyeGvxnPYaVvV8UHEeTF2IY
izegG4g6zmKXLHRJGII7TZnO2ynGJXokPO6ye/12wNKZA0D9XxBDYzpVT0N/YFv1
d6JzZ/fk9GVkwu6aL6r+N/v08fexwPr3SmyMKSmRDHoYSHHClyxxb5EomNOiBD32
QBH2JkQtCzQ5PARWEXJ4x2rSC+ZDdMb2saqUQ07fH7cwm3ps8mgMYvHuaIj9mxMp
pmKoD8yDQs3ijneovIk6ECYdYRznvhvoOBfdIQOEMEuADx+04Y5jlRYMqDN7bmbt
Bi0YfXZdUF4S+rIysRKdJaq/VFoH335DnD6/5R9ExHRF2AGuCsYL7oqsITkZa/Tz
ftHk+Lw2PlV4rNDOEtaUtZBe5NK4goyFEf869XlHi8936kqU8JfqtGMi99337Ms0
op7jX0xG52tsIkaUiryKmq5EaBUfiCXuwgLoEvXbS5lupJBgHZyA2Ly7t3VkW/Vp
cfoyp44o72wF0kAQOVlCnxdYKy6EnlH5KJj0aT1pbSDSN7oIGGKcQIfi8UHG3GpP
NrLiAJ9uwlD4Z+9BKUSgqXse/zoqMuKzb5IpHqTWjeow4+CCS9/7hKJxFubiT0Ud
CDS9QTBugIPgJ3KgrvulJHYNIdr5GcD+X3NI88nk0wtNfdWcFuawce2m+1X6GDnj
pSeLx0UMYtvgS3zqb3LNR56KymPsU3yug3VnEiFEaw1gFLZPppEw/DScbaccyXGn
ldSVECH4ynxzaOqAUEhOoQuXqW6orrFVXFr04f3lTkMDQOZOWp4OK+pEYcrgbX0l
Dg68Uxg5J6XsSAIpUEWhqDUqqwzNOT4UZVve4vQi276FJWPs61pSaF6XFxiCoZHg
yKZ+Z+SVputnhGlWNZRjowsQNBI2vNAw27/DdKHxb0k87hIvHMSKdNYE1UQZEpKM
9dNirOwJqbPW00KK88UFTO1h/AgMEAhQu/8dtbxoNx+IcR/Tcsm2sPv7+uZoYTmD
mpL6Szks/ySgmohhOV6neTfUeMTMcwBGfRzOAlYlFdMXTroh9AIG3FP0W2Npzc2g
G7MzIx/wqAWmmihmoLeymLL7yOyAq1J8bc0vU3Q0ZeBaKsu/ueBv4JhBH7DC09vM
lomP/Z+BZ45KL62W7WYmxzKU2kRh29iFr1hfmukHSUNvGSHkMK/sHXuWXoAxMihf
0Uey9Lom+Gz2wr0O7jOogEgZ11TA4ta0K8xC/YHuk737I13emefkh4C3lvXdxw8T
NkyJK1LI8sJjgsABRtloHb5yUnJpKDuPBQ69Z9L4FVonn6O3Eo85t3NMn3agHIgw
xsj8kH1ToT8fvLRWFdQ3NQ8yqB48L4+hfJvhlu3j5wUr0iljQMLJHR4rAySqtPYs
SXbm/amt8hUeBhERCF2cJQ5MTbBKJhAm12Oi+UB5/lNiJjiCmZTNa8oWerQbgpxz
3YrfPjOtwIeb8Tcn3bQGqtTotKD+kEyDLBCaZKHD2d4hUI4Ghe8E42PvsKBkpU6p
t0JHiV1KPbXMjH0jtmyxOTyZbOy60p1cFIMjmm6AP/WltJUAjFcD3ncTWD7DLhaq
auqwtPIbKLydTqmPdyZi/QBDOiov6UV0re1+zX12sGhF5xFuHeMV8CR80MscKm58
Ij90OOcNYmVggy1WEGFiAp4mFOudwZDNQsNhmphqdRYncOYP+y1RerWXaZIB2yaG
erIRNASaG19F+RisPBuhqt/FnPfqNilE5NQcJSKB2uODpuvrsoVIpMGffa+In3cf
FsH1tdHuslIis+qU7DPc/i67GACr5hFfE+k7JHlf+cIY2xSxjN4ln6+A31PbkJge
P5DKfdGvlZEgkAJeiZ1p9BaJ6zvhGdpmAi59EL9m3SKcQBKunCHpj2OXFbjaceTU
ODAystqvYpFvnSUTv+Uux5YORadxnXFgIhTSeWmoKfhZmYaCMvPazQqFgbQGxruN
+2PpsHDPXgRaETKDHUDWIKtQ8vlqs1eVLKxyET37WQ7tjKNz1gSD2WKtXoUFxgCa
QTwRobV1G1pc63wpAj+SEFYP4qCRqOAhhuISOmrnt8/WV5rG23RaEPxtDBcZpCw1
7/fKYkLxieaYHWP3650ZREvD8cNoQMQM6oBA0NYYfqL5aG17Yv/bLDI6SmKN2hbL
JAausQeSOv3pvdLyulUgVBRC7ymKOlB1P+nhP9Wufs4xcgsMMXq5J3njmUQ2GORG
w/FcD8+S4pyj+30fCTyx+wgxKVycPhJWutp6Eszy0xYUjBSQmjEIKdaQC3FhSekS
ipryaQjihadE+3Sg4BYN6kfUZk5+nGstGJD6odiGYRE/qtOb2K0cJW3EL/Xbkx+g
9bER8v3UTByv26N4tKguamqZH48JJSm2qI5gIXTwn8oMUw57+gtKfxzk01h3vICK
7kY4MjjcBcsoItcMFrnRDwOvnDNBpZ2e5w9gpP4npDj98yVHFv7rVL6Lw1V9GE0J
VAqI5MWJ89bYLYwyU3DdfheOBGesfm+IDb7bbol9fuVhEVl836rNnM24zDOWbSD3
SCFUn1wac8fG6YPHJycuUs/jTS6CWlRHZJCHN+lYwpJjHWWpeMSW2KAPh6sPuI3A
XOxfXdoxf4DC28HPYllAEixNa6fVjyKKPH8lYc9qDRkENlJs3IXe7KfaoyxH6rzV
EcF+QBzS9Yl1I1+/l3z1VR9jN59rwbAND1uOnotGgmBKlqpbLNI0mfGAiVnQ1qY9
GO/ShOiyv5TkvcyjJrEHVoDVrqti1dHsf0AYdg88PXG3ijwbTyq1MPyKbxiIlUNR
1Vgnqk04e/QsI70Oll9TRUeTWJ24gS1t9A83fmyrtLH0zYm9Lr/9WM3RH3+jTjyq
o0Hj35X7ms6q+o1lclBKkJxGbxy5u3O5tW6Ntsy/5NWqNlTKVuVKBEFDx7Ik4xHm
/zGfhyBVqdZh3JkhBRL4EStnFoYxiYGK8WGwl+v+s0u0qyUtIaOIbfWpH1NvsbH3
O4D4zy4pmqL0DS3+qaOZzV6ud7e9UYbKhScQXLrE35WGZkRqpBzDrMlvjuR7cZTp
Cr0B2qh2C+Te5d0rW/tmS0y+9rDq20YczQxQFH5O4ge8LEWDE+ug2B8vFnH6sO0t
1UwMaUWfWl69TyjTBVXEeEKNSR9nMavqZnhXkOtDIA68PNDLnqbSWdHXEu9sYH1p
rVQnm48aedekCFk0t00XcNDpsQOfKDRwjY+ML2tlwUguokhf/4sLUFT0dKR7ge6N
B0GU+QhGE1fushGAjHSMwbqtfPcEhs/CwmrNIZs2zxqYTKkt0P4By93Rfvqcwx46
MRGwXSuBtEeyOYuiCnjZfopy6XwzZk00BG4NWnrnP0YARQpmfDj9OcXEJrwTvyU3
GySdkPqEo/JUbCLC3A/bleuwBx+MXqgb3evuwV9NarHbYycPe+qu3eR9u6jPB8I5
O2KDI7CpShO/VGBRIqouar6zq8kSD2J2hDXW9+yjFWy2MyhYvZzN4P7k13+Q6zGy
zwPwuqwuoo1ndTtj021NAW0LCKG2z2iEsofuDynTieZ/MA+Xwr+1aceml93+jPTD
uwFcgbydP4dbeS+12ZSKGnTWnEXZOPl7VT4dsOitQ4EUmU6MIwl/gP+xga/V5R5G
IfzUuEcOqv1iHlhH+InHjhGHw/bZrGtA3i/rLprBWiXTbIlSzD7Q+U0Vt+2Txl/7
3+kxJhaKaDsOXezaE7C2u410OfDfcgQrvbmwESd2+l3lIygUjeBGyRQVLHpMAEyM
SZfR1Z+sYEqTzomQMGw3SS08DEgIdTXZkfaSFzAV47/ktbVdivOamw8XX//vlG2f
flOLH0p9cZsM/WAoKuuJ1X1N9RO3RPY8ZnhUKHY2nmIIF/RZSH+i0Pz1cVg52B0l
hJhT82AJkHHItWi37O9Qo/P+Dlu+WLg8UCDuuBUwaYH4NZc5c/AU6r/fl8dDtNxE
4wc9kNrzKmswvwEUxXyH1blEvhOBJy/l/iJiXCpl0U67BwXCfh+aV+pl61SdFi37
LyxIqKHgj56AKboPyRK5dPAKJLLtgPdPo/0X4kO+V5hMQXM6jeuZ3+oKBR0VeaFF
cjf+u3FUPbLED23t3TqCaGbywm6ZXqr9KI45J8O2Kei+4NfSxlxCsQW0STt5so6m
Htw8fNIQfM7EWyeHId+vmt5r7jAzI+xMX6VgItu89JlAPllIZ/8ue5z/MVFV1Qc8
oyaSLASTnNeghmtEiJJbb92jFzTkNHnLVC+SBWM3Dj5RDX0PyVY8WzFUGGqz18rh
JnvcU1UtbeCgzjx4dVSHX1lH1KL7ehJBCqfmL+0P4kFzXYDk2hc8gtDeDX6sMEXn
6PC4BUbxTzm5zMaHLvVU202Z0dr1qb5xlThsit2uXQeYo3KxCpGp+dYfRaga4g5M
L3TSRtkxRBA80PN738GQI9Cqv/L7BJlyp4Sy6PYVViFIhSEQrHcHWKt3oyIlR8BI
jYVN8dAdITlJzX1ZEDRgdOeGaFCK1rmKVTejsvc7JUzfe/ONojIfVj97x6UoKkxk
pOYXUIvgI0Jmd/bEghKadDKTj9Gl0+w80e9SHEsbG0R6kU80W+BtcxRUt4xnwK0w
s3ajWL9rFzL8IVaIqqFdvrqKgQLm942OqhhLM05ivxZGOEclJbeX7PBTDPNGHqfH
aToy9NClQCZZEzw2rjqbyTozpJv2gLSuovp1YN4+Zomd5hwiZdNBnZTSUWgyznKJ
EqjmQ8FpqTNxZhj6x92Uhl/jRPRRqqnMY1S7mXXvNgQWmB3aiVfLMHkaNVYRqv/o
EdOY2TfHX69K2kzE8xHdBXYnhuYnj2pg4hw46RvFPVFO/e9yFzuUP7zNp6j+m5Kc
wYss0RHGoajBmigF1E4QKeigjZHGIAJgGr1jLk+gHtZ6/nIscp5SP6tyXiTnW5n2
0nK62glzWzUq6Va8EINNX5PL6Mld3QgY5Og3HaO2Hn2BEWSueeaAIUKcyY1pytI0
+k9HFVXxXWW9tzYsxLZQdwKPIexCXzcx94o10K+EdG780xD/hjYncHxV4szAwhCn
vBJ9o2qd/uRZsqhOjWMZYNnLDZk36UX11AjMTth8V1DJ4EJpiir/2sR9xAMBHC7G
a9OOo4aP8MqWOJOclCxXU7ycK9XqlYZPyyn9bi1gI+PB9icWhdn+vKJsLlKVcKAA
6CG+tyr7AGo4um8OW0qToQT2M9Rk8bZWzN/L7tqGLDBbr6OYiGxNTnJjt5Iwz0zj
mxRPQFpZVJaewrXuYPgvThEURDky0IWMXDSbk1MKmtAx8S5xpRVz5KogY6M6BsEE
034hKQTGWv84dTcMsKxddOCRS58eMY0tcW25YRBrik5Xb/k7GRfIGPMU0JC7+ORB
8yelqK/+h0AqVFrjGx8ktqibq+X0fLl/nePHyLIgoTEeLQQLE4x7euXEORw7e5Wa
mte26tEecfSmi/LnWFo5RhkuLkPlUBrgQMC6rg9HxZ2RhX8SYlpcWJ2lQ1DsMTsz
jDfpmRzvrkiIjU2LpnlY8AVUjjHBXfzYo4UXCy5LVy64w72rk0POGvt6CgWuaBDV
05ogMxNLOz08Nnj82OwTzrQ3vwiUo8m+heISGY5TGg2r3asO0E/BFjpv13u0fn3Z
XY2zwgfZLSaXu7G/4w/mZcA2+ywlmKvjlNmWf8FNVw6V8xWHosx+cu5iAi5EMCfh
UoQ2/ze48wZZpBLrkN4gtbTKREVoyrz+meb67NQVQM+bg5sJiJXSgD7BxPFKTgkk
b840ovlpeeHl+KbvzdAC8NAL+HgqrsmGjTMllAeATORfDYUKvKRBZOi4DSQCWEhZ
Dr7KWl+u+JVAPtAD2uQRZqJfgpPyyE2inHKho/lqU9bH28xKnyu+CQva9LTYHoG8
sYxGx9AFC2QxsFxjhUoaZekwuuBTEluhBeHPl0LvKAxZKcFLElbgVa8qo/gu2x2P
+6iQPYr4DwgvJujBm0aMFm0/Pcv7i55wVcqV4+7DzjNHpZ18qUV2T4UuSWg25fHA
tm+a06YSRWFBu067m4rIGhgCeARHmfRAe3MuuRgIqU5TO+11BEfJKev/XOjEiI8Z
rLMumodvXRc1zJJC7bMMuwpMGVPrEZryM73jJhXfcPVGSvNLF35yaO8UOKyYee1J
f3cajTcw4b2WllXB84yL50XZ00x+2FR7bqdgyrudHLDT5rtU45//pWyZ/OWDYn4s
PRxwp5hoAMNMvPiZtnTXnH0lRsBQnQ5G5GSO7d7nGJBjt5pO3b7v7Ax1QCQRGYfF
pwh0b1IxnkgCHWqwQaSJzSPNrjy+/gC3cckSIg9zN9fbZrxnNCmhyPAO6bRg8/ek
/SZpZ5jpOnjs0Yk5T2Bmys9QT5wy5qYHwwaWklC9ziv4FxXtuz1m7z+xT8tyyX2i
5b6EbnSKnqh/iURiuzpuhkU4cmOTqXF54SDfqO7DfW/ML2pvyOsW7gJj1DYYaVQs
tvNwQWuMTyviK5bHLT/HD8tCYuR5q+cFKdkld0a/ReT1W2F34nwxBLzWVI/ieRHa
7uM86q6CmxaQfxO3qKq0E/K06fRIWxGk6vbaLFOdeFPHZY1l67f+9rdWy+20D5TW
3yfKpczNIC3GpL92qJwTYxYAkzlouacG5baAOnbFkn51A8XgHbAfDWumx+QeYMxk
iO2WJl/3NH0sUrveIUHeG4Bq4+KHbsDaAaTHtw5yweMMIrIezOrZhZ+agVPLiQY6
zcgpaReOU5GUhSNf79fPjImcro+ipFcWJeFud46v1AfV6PAcMTGaaLGvVqOyKDY1
Z9JQUtx0M47sMZCPCXOd+KuPJtrXG9DjnRYrfGSDQUoM7OL4shxpghp44eCpAbuH
dDpWKAt0mSXbjvKz/FRni+iFOQCbm48fY8rtGvLq6AmhRluisz2Ob67t8UNNISoK
GgwdvZWAXCcJ+Um6sPx3k+5IV+KGXgFEK4JIQY5Gq7GP5MnJny1EtlxhoEycZQJv
ouWIPhxHm7zIHqnqosIhsowtqhcbuE0pJKmsR4dYYUaHst5a/iVEF4JKliOUNax/
FilZc7QPQfQyu1yY2jHjR+zdtjpcVKIG2ebCacNXmu4muMOiJy3QtV3Cq2/0APmw
xL52Mygb8yOk61vuN/tk2W7opJV9Tx/hESsQ69GzJyJQk3w29QM8O4vMQtmnLm92
o8NGOp2AZEPOcTvwGPdMb+bFQuFqijcBM6zLFXoFg13oMconArAPbPU3dM28TTBA
LvupcUH8jw+fj/jwaUFNcZeyhXLLQ3qxtSY1OcJa/QIWlgU44fVqmDLyqq2ZANUQ
SVFZBEeGK9IEN46T3ylzVIIOZ6kg3Yky6Qx3mV1gsXDmGv3EtNuxeF+vRi6nHBSj
srMxQeD2QhmDiw7XmD+SMAuqWp1Av4MrJqibjGsuNvayVmvMeT9ve2tdLV/uAQmQ
BCshef+agNiN2bYZe2HxXmKBs5JR+grMjErvcKdcUebaJjMMml0rsozhPzGJMqmp
98BmvbI5Havozx3YeVu7t/zQKVN+2DEc0ijsHXQQl7GMi3fQZspY1p6uazVqHNE/
imeEY3bIv05MZRZgJ7f2o6RwRiaMGZ+Z8IPVleP5EijcnY7QjIyVp+laBmZLGblG
tz3Dg3QuPrnSDdZIb6rYTRsQZKuBdpVkvPkTah6E+CVyOv8jn+LOyIkq7F+gJ3F0
18XS+2jeejxM15p1zKB/X87SPSR+rQm7bJUBUVDEFG0Gvz7sNLy6OWf0CijTv8kN
nCAuNrjQyvwuwTMUXBUB1HN9BMXMXnc87XF4yvGeokYYtpZOpF/J4YeMXE8T/0S1
Eu10z5WFsaf3pcKlR1uggovkPBqR6OIPpOoAPh4cVHGpuVEXrtKB6FbsOwX57h8h
YTcXWSQPDCmM6WKhABTonsSsff+JI1T7/9x8X/E/+g11sjiKKh/t5SUdP0UN307g
/PofX5DQm4KaRrqVUw8HjJnRatfNOAS7HWTP28Dop/cLaSxnxsvXJKVJKYs214M3
tRtK1E+Xu22u/gNFdb6+F+d739/7OyPeqL6D3IcoETVnHbV2rl2NtBEm6GjPcC5D
rtH2AoaJykUYHSUzda0ck83tdGtRkNiha5XmG1pA9xpjSD/ICiayQngUW0swCq2Q
vrabMMSCFp/cXug8Lmb3s9mKZYNyCPMWYb6uNyBoOIrLyjK6OuAAcvswpwefYJVU
ghyy0OSXOVJT1EpxCvvhufW4GBDO/o3UVJWWQxLWYxu+weXNRwe5Ea9t3xavC6xA
Kyc/8vnzabjUHorCc+ciAO3oKKENe4Ox1IYasByADWJpuMiYaKMU32xAHUzy7N1u
s+gRcScYazkCn+x6zKNbSOHwRbzXAA5/mb1IvK08UdPSpa25blrR/FkfUh6HgCg8
ix2J7HJe40AuoNodA2zcWvjE9cfp1nl7T0+xek1RiS/iBs8V9peImVEpsJsqvt8Q
ddmDJOPbU5M1gKy4zjK06lTN6HczOdFUEqGKzszqZckM0u7WKAp2ulY/S62yg//D
Mx7T2DY7fqWmEs/ziVR87l9JYPwstPvENyvRix+WIpeZu+R+3gvYv6fE0Nindn3u
SQkgeRaC5GH1tOy3vsM8YD3oW4/DT0u9+fGZ0N9EZ9DX/2fkVyHFf4fp7DRL66Yb
vjtdNWmThogp75Sjj3n60DwwDvxEtAVap5g5KyUazG9//GyrvhMJ15P+gNAkXpTM
6YcTWRnYZxkrweZkgSu7S7AuNNxIL5t6XqKXC0T6RSsrgKb0/Q9yaLTf7034GuSh
7VXmr3171ifCeqJnQqa3TQRe+T5jRpQbFa9sM2G1etDUcYghxAqDKhgiM5Xv0z+q
8x0gifFUa9qjsxmp7u/af/B088rQfAyHiCkNWuYVwdfQg7pQAkbzWMPeVEaWz5iC
xsfuzDty1E5cXe0NHGme6FQTGysPKTaMHqQSSL3H/st1CfPCDqygF2dP8q4b+RJl
fqZq9LLssJJq5rnF0qMnTqGIrUvq/Mcy7/G9Fsh9yFJk+SOLeZEyH6vRh8KBQ/uF
qumoFBn1rWdOsQqJrVrwSoXHDniDQWBPObO1QGceDedMDp1qnfeHsPund+j3gLBT
Z2dkOomtkx+GqVSGeEB9HrmXFZvY0a7/BKOwk+SCHnzv8bFgsR/1xQAk/S5a0blt
A8e4p54MqOxyts/GeN2xliY099nwjSMIGbXwWoz9Plnxukf/rqWHki1c8usv6Gco
ytf0tgPslE0eXTobkqagNdZtYazqaPGtKDA2qDGls8m+leCAhI/hSxPERdRLaOfZ
8tNvfKjUeOEXPmvH5vhLn4S8rxs8bZuqwiVfmK1Dl3uYMcjqxr+2IQhMLJGm/eLO
1q9pbzKyOmZHX7vyAO0OEYfBi+j+B5i+tEsSnhBsaooetIY3UJW/N/4Yj/J/x2wP
5SNU9/77FWMVDI9E4GcRszVnkPIne1xpT4632kFUznkiL42bD7XzMSMEPkOJsiOv
Sj0mA94WvgnzWi7zhNfuOxu5YOG0YmIQB+hXt92rccy7PaABTUuiZuL3/6h4ZMS2
ksi/JTbmyslKZNLmqYyL9o3C10tY68SvS2y6Vwjh9l3u8c9zQclIvIl12JNvZ4ix
B31b5wsbQKOXO9VA4L1jCmwALZdSOrAuS/RYspOdCHWLueDVAKwxd3ozDGrQsw+n
Tb1IHmQPau39B/FWmE4jlKapQXa1XPYKY2070GGeYafEja+Ol+pMZcjwR4lCCW8D
TE+8QvEWbxJqYGmijkw3orcoWDtPga48zqtG2TUNg6N3339IVO9oyGMmV0h0VIng
UzS+1OssftmkhqJZfy8mzeoZnmT6s8nDY7mvfDizfhbnzv3pLMau62c1osppw0b5
Nc0KclcoON65/6zV8aYO80EDCoZd6JS+8AdYsSFqcy/mL0CjP3yd3yWxkRCV+qzu
d0rzP79Xg557QWBaGM69SbmveEkL4PWVilpXbGvvDnsI8EYWR9+f+d65gw0jJYFC
u9/KIFeCtWQzrabIaUx3AaKxMuMOTOb6D1qp174SyoPMk5lubAiuL4ip8SgRv4DS
/VdgJuSxcIIiUjTV3WSOl1/nyo/GYNlnXYuw6ZwRNXh0Aj9owdHOqSa6QYOfp6g/
g1lriCtDJWlKWjCZmz5g+h4wGrf3YJ7qBzwG70SHm9ThFamejwTFP6XrRAh8h88i
aE+dnkKVHCf6b1IxoXjPisHQwGolMzJSCVGL54bP2JPB8ukO2RZGbATTK/SSJc0U
TPSioDFJPIf4tQQGd1G0LP9dfugmRPLQVYo//k0G/P7EV7jOho2BKlUdwd9ORun2
vZPQaVyIvJTcjADZ07N5/gBtxGE5plCeKJ5K90GlvP6vS5IWYctQQEQqmMtYimsk
nm0TfURznqRRPNbK3kSZGM2Tj/EgYVrlTpvCVRXrakUjFECq4Z9WmMbxJ2QZWC3R
SEpkV6bJRNdoXO7MWGZB1Ts8ZeMGzgiTaVvu7jmnib9w/7BIcvOBOxxGwEZ5ykY/
g9WHj3XQopcEC8HX3hUYb9TPhO3SK2mvYATeCrwmr2efF97561e74OhkciFxOmFk
J/h0laYvJXHy7X8J7kXuddI/8Lpe780S+7VKjA52TxGwJZ8zCKjTZelSPe9E5tPc
7wLJOqZ7Y74VrN/bOOQ8WZ5p4ryxvBgfZ4pVj00WgwkDsvnZRXPK2q07drFXP9Kt
+bfzmhu/DYv0IOAC/eiQvtjnuLOsecmo/WSkI4p/I/uM/rZvzdVxUBsULpO8sPg5
MU98KWUJ4GA8P5XHSCHShr0rjzJrYhOSUU7Yr953LUh8qDGEOLla+0c5z/yr7252
+0/PMHqxg/RzIjIKpaS64RAoO16dM9k9ooeybbMy1OzesxPdEfbIy1+hx2/cor/b
Xw87PsBDQQZ97OHE9ApCNS5XE6zwbdJXCiZO8/ChBOhfA9FTeg+1M6Zg6y+eayvA
BE28m5g1LI/IsgmTciQ+ykVpCeByrzjWnlXVaW8/NNG8t1QAThMEOUg0d1sWBKim
QDUuOQ6b0Lc8dr7/73tL0fbPDUFJlYb1kRzRCeljU0SZbV1hZE1q+Mc8l3FOs9ot
3wJmUvvqKof0hH8hwpDwC6/+a5JljoVqtSrJRKpphKOS7PvmjyQRbPzqhPhn5xYm
YwHXPgDVLtUmfLiJwr0ynBhoyFPtMXeovVKlMPlF0TVpucJHPccPhNWA3a0cdb1E
DsoMWb5uZ3GK2/c9HMCJuExlm/DjuMKf+osoADU0GcRee3apzn2YRhvElMn1Ubd2
fRj5dwPhEGE+lwMCGwwHGkCLeuPup1RTOU2Zw33oyb/PCOk7jHyCxgmjFNQm4u6v
Sw5Cy51+7184KHeDi4vGu9W2AQzQa6RMRTRo1+UNJfJifeqTaOwLcMiMpdLeHj07
X95YDDhOSOzbX2TIH36qnRieRrBOws00bbfOHfAwZS7GUHMSMB3tY0N8fQNJoj76
1yDzAt9ZH/72Z9g04pVP7T3q5T4hzePt6TPnXhClaHfrr3/CahfUGOn8gK/vEWLS
Ggxw3EF5Ddbj/azrgSUelMoQhAESi5aB0J58+VY5+WgKu7gsWtN+Rs3dg2diQIOK
WPe0moPOaKHW7KPmAOZuZrNynNWbzRwNXJfzkxUGrdMjDWWhXqIgyucO4fRDgOIn
Le28e66W6LBMA8ITTSFWAA+qtrZN4Z69yvMvtNVtx9eeSZj+DAmFodzSYU6CkGYZ
yz20tZTgoCnCOfnkRP4TRSGFnXTH0Cl/MVlP5r3pLY1xSJN/xn5nL/tiWe5v3eRb
9SSBnf+Dp+5rUtog/tZs/oR5iAL+2kOcBp+R7oLAhYPuUPnA6uKJ8v8rtsGduwIc
URcgBO2BNqvtkzzKzplKsoAlE3RxLYZoHwCtNuLDEuzik7OLSA07+pX+DTSBqzvi
wOgGc119uFcko18kLQUmcmSn3wxHftV+ulLmJ193w3Jyk3x7PCaPf4BoIq+/8LCt
BPwIJ4X0SfeZJMStl0Yuy0oNrsULp/XF+iN6ny0OoXRAww72KLJKZc1TRwRAwVag
slFojQHj4afNJ0FYuyoknkx8KIWpeKnxMScEYFKlUbhK/6kNMbAPUp7BGWrRKn46
vm8quwNNUGwEoA+V9zIAe1gPjmNw4aDAm6wd/w76Uyx6kFjOPk0l0MUppXj6vn0k
zZIXmb6vqi3ay3Ab7N8KyIM/PjOryxs3z6Mkh3xvLlwBaeRNcmsyAi6TxG5K6LWF
FXLtKXHdN3rJj4mOpcW2C7RN7Nbpoqtq2QEF6fPiUVM+u/SO0HY46wMf7ODFZgR9
gHRxFLkRCHyVxaQguoS/fSq9QHC/5PKkEvmGyUJeVKuDhRY2sFvep4IkYD1w6p1e
xgC9jRTxm3q54cikvc1m8SOU134F0pJDbLAe0T1+hJz0YcZ9cT2MUeXqZOXg5qCE
bBFMTQyEPfZGO9jlBQ71N1XBu7Dg8XUgAqyi0O7enoiuKDAXqhBIcYlH8XE2keAL
gtzyAe3pDAX2Kz8kJNHKsO0Oh/qbi9r5e6aouHyvb8/oG8V0jPVhIDXKcOKawLjE
uKl+dWYMep4NCHZukCB9kM90oZANl31CTPG587eeNwmGrV1P0Cli37Bv3iikOuhT
eh8rHG4p6yEq4RNUKib9/e3b6p7rcN8CDfxbB7YiAtG3i1i/2u70gffjYoU11iqC
l+w/Y6vF6G3shWs2ki42kb+xRJ8xh55hAjtesgCTu4eLBW81Twccn+pHY1DlMT8y
8XiOgbe6xVzMqjgvuhw59nR+lBGjpxSsAuHJqJmNfviJUjDzTyawYGa1SV2RYBxY
08vGboCqLYW0+znGpsOCXqYChoMbg6AoUjv4RMk7gKE9NZpn/4OG8TkM3wuinTBg
rjCYMA8nVH/9plYDB6BBdUZ1CHhz1h2TFaHoiofKLRkmLZmF1UJJKvglC2NfqLkY
oSKO756xbS2AI7L/xP1Q2u/Ye5rtkwKM9HwhGauRgJzSrAa5PmB/mPCKxDjWYOeZ
NxSLhgu7fIvkKvMtmXs0iP2tSJuLgcAQx0ZbuzzYWVfrQcfKVfxf3+lziCwz8RQb
QIOqn5MnwyRYykDJF1etkfKlbw/4Bdm/oddrWu7gin7rvAxbu4rQ7zf1FUIIStej
stCH2FQmGrcedb1Cjz1o74t/4VgGSy+/0q3bc/1bZhqKCEHgpFyYVQqWX7kt+PPd
vvOLo5K3EY39Ot4ogcTE2h0a03QFJOrYbZR46ppeNJLIycxoooKdLf8tUPrCxs3t
umj4sAvJqQAPaGkZJ8K0LqIO9d76yN0EnZShhA3IEcS7qirjJvBS4mOAmIq4kLcb
e/RZVcWY53iPRY+BR3jKwMfi91TA85vY2XQ9v3xPE4Ydx0NEFlRVhay2o8A7Rwfm
g258Lh4v7FbQdB7WrmwPxQZ9fWMt9Ges4hPVUCXM7R9p7+MpqNyJ+CU5D2sEe8Ls
lHzD7MfI5yQNzckh9UAadmlPA9/PKJ+SXJ5/gShDhrM68mKwDGBfjiqfknU7ECqt
vtz/uqqPjNq0Vb/7WxjvpgBTpvxIb2tAOaR7vBAhH+DYJgtFrr+nbIg7W517uGPE
lyFxpAa9liX6nz6tzB0QRHqug/J67UrRaJHKwU7K4DeZPxnQ9c/3olSlvQSKhze4
rWVRZxyjQDonXSIMdz0q7aYNxsXp6PnsfTf202RlLrtzL2EvUrIqZE+6IFVQ4BE4
R7sQdnNRefRh5Jz4jU/SzJgNT1VjupKfecQ54OBwcX/YHZrv8rtpdPbKf4jXpdDB
FvyZNpVg7PYarObMasWEoi7XFrMHZpsh0hqmdjcz8h0UhWGD/7yXQMY2LPq9pz2A
XacH4/03t6M5yPxzKe1qsJZyGjRmWjF2TVYeAE5UB30iIU/bAjpoEApUEiDT6qWh
wiJWW27ujrKRP18BG57Jtq7/x9g7y6HUujw1Rv2eWuueE+qALWlPIgHE/N+o8SeR
dKGxyZl+fTtwOfBe33iXgtRIbtR+t8F5Xvx3UVN7uSrSp9kLeE08v9N/JtumeEXQ
Mn0M8Yq3q5Dxn79z4tltXpzz0OT0svlfIvaWQJk2VPOVYLmjteWT0TNu6b+9jmBC
Ir8Oluf95b8JxLPJ5q2jOLgoqVtE707ncsTcIoOOH632PBZYgfy/NCPRnLbc0nAC
X2AMbDmqLfgDOWfOMZsH9zqgoNtrdBK/mbfaqKy31LDStB9wFUn+OplO6FunR9dc
Rlt7jhbNDTPIoq/afwwUBQgmSKbkI+bpe3RxwhszJFlyn6/tMx0kt2L5CXFLtsfz
rGG0xJpviznYtf/CrSjLIS1b+F8pIAqIHmlmi32YcQMG4klJqYnTdPLperrARYLg
vHxCfx77d/6dj3nwZFA/10lq6GTO24LHrtQITDxWBwGYoH0n4ele5HalS+EKqV4j
r3xBwegvmN19wX3vRUOeDrp7f9wcRUF/IJ+J32VmdkKPYsCHqX9a9FIxB7W8KOcm
0CgYKGe3U4295Qvoa5R7d0nk/OT/uM4y4hALQ9SqW7DgWXStWnImROvoereXJAb6
VJKdgrCRkvFhT+MfaOuHHWDphNSPZF/kSUc7anTLfms5niI3J/AvATSjw55e/HLO
tY3ZJqNgcvNRBK34RKFxCSc4jzHWygYI18gYfhs/E+sTlV555frEDtXbC82btr+L
FUIRSLjA1Y8BpoNegYOUMiHXJgSIg5KAKO0lZeSKUakOM79iBgpZ7i2ESBLn1lWd
hrrf6OzQm2quZRmbC/suvAxTxOo+lvAEcgU8t7zkxjGkqDPrODYzPvjzuqL0j31v
tZK7cKsvMr/iLr2HWB3mIX2sIp9UpGsqtFcLr6nMvXHzZU09hT2vvbhNAQ2K1StG
StVfv+8kgJrKVauBnW9xpu8oRRdAX4qYrh3grbd3goW31llyMyj9yQ/39mOp+uoI
VIuQa/8Cy3rLi9KQXj53KweQ+vY8rneoWIEA21qOfmjhsC9u/IB+hvbt25Y1/NM1
p/afmhm7T1lFvBlP2B8T91YloyXXRoDL8fgwdT7DZA0Bdoo1EIx/HS9p/jLiWvB/
XQdu+TcTho7/GluYdwb3H4oZCFiwweeVIhsRmhN8YF99jp/kLlDyt7f7ozeTOSZQ
+k641a7OVqAtMUQH+tvh8fZFuPswZmiXUNovABAoJNv+PuPZqdaKvZDo8a5uzsAT
5e3O2GcDJK5zCOM4m+69ER9LGd7ls2oqaICPcramNVxECZTA5xycyBxkrNUCUqDe
te2FWSUTMzyGKHRF7n6EE4jsTZOVkAl7ihf9F3cWkr5/AoppextRCoBpINfgrN0E
NLKUTIf9oAx3xY1JUKkDN7qC5h8KsjGhUlp8yPFNcem9RXgVAlIBAOkf2aaOnodS
wZM3JA3YuvdD+VuRZFV0IhWkmwa3zaV0UlqXHNDKsv2J/mbOJ+o2ELRkIcOBJ3T0
QTjq72Aejnrhr65LD7L22zc5IG/0r/09Q+KPH1tO9K4TKURk1LJow746k64Gbzvx
v5YvqQ6rH2FWgks0yGyeYQcSWWKMm4zQMZmJJHuTEToOVpOiR45/NeQUhclEmIM2
+d5CyuH5Lit+gvzFFPA6zOmMWAF+5EnWvy7BRsXyc+cEriLvI8oBmbyrobtwzYq4
VVCqv+dCjE8owCV33KDbfZWk2/cdp3L8FtAGNm1iuGDE/JLYuPYnROSsrBywsvcY
6uLiG5WMDu9ZiI4blL3dS/dSc/bMcRdGAYj8LXye3JUcwPsd2sIKXwbFaOlU5NFL
XAMoTBwx01KDgOqQrbHHmHVG2EVPdjldQqURkhGODz1XAIH349FxzUDpWLWJJQOF
a2mywTm6dk2ImrOwXmwZcZ8QsltXD9+SdcXar3pBBGy9hy3cNoHsTSmpIYJZqaAp
IuCJRmp8sil5wOuP6wr5Me02cKHJAAaQigdWufPEpCBHUC7+Enefwwqmo0KZXVI7
q8xPjOvcRlAhfhrgAjfLaf7lI+R05call6/gI655qsMKBvGNYawO4pBOMp9SRPo7
u5akL14/IVle8h6Y54byitkbvf+4PQCWfyFm21lANg5as2h9iwTjuF7O4MM80Fc+
XvHRlyvM+O2ZjJZ3llxDgpL1IGl5ekC96dMOh+Pr8TAkBkqQegMWGAHn1p2+F/Kq
T3hlcJJfcMx5hKM4CmsnfTIWC5vtHi2Rg4uMjHAsAGyCCZnNH1z7rtbkGHq4OiGx
nImxskUOhHk4s2hpKwQYQ3Qx76VLGv0PXeyeg5suEPt/uIsNliAK8MlUkfy0OpLX
bJhycjlee+r+NWtJCQ3r7AN9e0DvCkBciAXy9RmtwcxqmXncAiEnZk3HFcjzwvaJ
BiqldHJTu7Za8athb1sTKz7nlsF6Dro3gyRbwBBtQrSQGkg7/aYP7YB2fnTwcfNk
tp7cpEgSaIlxXziwMTjGn2o8B5C1j2E9n+pAMaefZX1X3VmYSKQ35UGZ6IT7hYwM
AF2H+v/mVzJk7spHEYSsFe6bccmbJcE2o42gFW+gFhtyYT4GZO71+ZmX0h9qD9x8
y42cy5h0k9rrAnfKwhXugi0bWUsBXcCCa7zqhvmC4I0m3lZ7k+XqO/RbSQEjDpZN
Vs+4A0gWgv3osoKXjQpKTVg6150+PxPr1iNFfT0OBr+Y1ByYyQeu3+sKbgwgXy0E
pjDOnp9GeBsqrRQlHeY6IeksVzsKXas0ZyOSQgINpVhbcCCAvDylF+6dxgRycjRr
uszITLGVu5E+nvMQbjD3VW2Bc7m6ln3R/SSs7E/AypmlZudJQMXOYjYW7+VFA3r6
sQ/lxOzAUbGlyiQwFBupLy5uO96bP2G+BmnmdGAfatWl6n6cLM7xoHYF1koGepyC
BYiFjf6TtuykPZoHJ3dfwnyk6/7gqDPOcg3WVlxkhefmRzUPKFyfWG3DnV8AJCTC
FXO7MFYpl4YaUBkrZbCM9p3LkjhmSPi2nYnVCTIhtlNb9vpsI0txOysL8o+vX+Mr
9/TRwKPYGc/6H+0IExesGHXW1r9jAf1c9+BRZF3s6IOwfZ/oU7XT/2AIo0upQ29o
WNnxexXnSCTMxkFUAVDFiRtRkrBWtDzDxK3e7aUAhRqGBBzzD6aFIZ37wtplxyj5
s3EVXtJeTuibNHnQcxNa0UQlBTP4uzUvyW4sPsbbYe51jeeU9c3JTwYu0XqU6y87
5jBwytGr8B/diNGdOqvr1+XFo+Vl+m5Asmq5k98G+EzodYS+Qfm2wqyXTUkN7bvR
1H+0+l7mv5pUdOusFC5lhkBB8q9g9cEVYwmGfHaXjzAuqDwaCstkBaNuYCaWzcYp
iPk99G17q/ao3p9a0KTDsxvlPD4bg5m0K/zFrLOgsd8aYmNAYN9KGaCbiaeiubIb
78t/jbb8V3Q+/AaHCPpavez4NJ45CH4uBoGzR6MoL2ljwSSwD2pit8bNVQKZ1zZm
k5YC5wNBIotjchuPv5GiDt06ycChyy7DD3qZVCbJxfd003WL5bawHR+e/4hskBoE
FScfmHhCtq1SIfQNoY6+d6U1+0o3Nr5yCNKPiRfBHVsxnh/RPDLgGekMSTbkA6Ul
Z2GhieANpghyEA48Sl44yHQzvgAAPTEQlkZxJ8jI8zUAUp4j5cx52gngeFa5dGju
4BETjLvzTUPvOxh4XyVqwcaSqCApSbPZpQ/MwjMF/Fmmm73fMHb9xiJDw6H9WydB
IzgliMzBj1+tj3K7ZEfWK82McjKjuVLEXOeR+N1KpXg6JMilkMQbl3lRSusGIqvU
Fur4LPTAK+Wgvhc/rRshoi5Aughvg41vP2BrjvctZ/dvJDT7AY/Yh8sQtoiNbyo5
0rcXGIfgMR8C9n0EQ2iXeISbhSjI+SIHxT7Yn5W+0oNv1+I36lMYI1k5R3Djt3gX
km5pKHs5dH2So2jg/vUPanVr08vHIC6ZnM4gRKie46loZ3oIhZyz9kO9XeqZ6BBp
GAXwyKGqEe1t3Odr4hxBAmhY+yiplWBmPfzIwhGw0qNoBvXQLvyKV8YsRTM8ENeg
85Jjc2pxGsJDea0DaVCZsCPAYdzIlsw74qbwgDGmEszyn685ikYZNCe+cPyeYYEw
aESabu1lU10raT+IVkGS2UsvflIqEzea13MJUwuwY/Pphu0uqpFwcTf96/dlsPKX
TZt/JTgwikcsDzDHjItv9bchxjwBl34zjfrxmyuUsGgFfh01CfY7zKQPkh7ZM03C
YRWP03+YzSrRNnQqfVM+Z8Z6tcFHd9Vk2pZM9pvx4Z+RCFoYuWNIlxrLlXXEVm66
JOvd3xtcVVEcwHz7Oc2f6D02U4hiOEX7aWkkY2zSxAiIgE6w9tAG+Hn74HrEQApT
KnaqdBn3C5LjbWj0Nqy+pG9YFZfi3kxu6X1ZQ7gGhvD92NbCL626qb7v81PK8yBT
tZq1Gjhsd7b8792XxptX+U3wav4RuPNgjOGegR7Xft5xigIgtEQqCBhNaRySXu00
425HHliAnb3HTXT1kE2U4wu2UljI/NZVn4n/UkylKa2C959Uc6lwSwVDD4UqMy1c
9SvL3j+oPxdTcyQHJpjFo5YttnXHkyTgGifuRigRGeI4chu37xvqXmXEVHn8JRqK
Hl8usqyyYs4ahOKctBMbmBhyskwTQJpMZtSvOrq83u8sJ4fuuWUL1I1Q2a35I1Ny
iVIHzFzPUdB790SfoTcY0gz/FtdOHvWCotx5GCm2PU7dYu0Fstg3nFmK8ALifVpx
d1EsInl3w8oLBaQPlx8MMvUYe8aAHMKm8agfb9jr3mgJ0LnNBFNwpEKfhSDFz3Q4
EHJitqe7ooyzEby4TUXqY9BCvvTKE8sH5KhcgyqSWOvukAiG5YrB/Ez+GhIRZMhm
AU5DFbAbdfzZ2GWlsT0zwUvQ4nKjy+DB/jU1ALgg3CN7vqoyyI9Mr+dcgIrONx/z
jqrpNIaVD5iB5/SxFzn2zfwjvT22/5uMw/Flv49d8l/io3AzrgK/F4XGFGEPqLRz
k26v0IqG43u3rFjAOjIcbdcXjbyqEiP7TOS0LihfGBye3Vpm4i60vZB0WlJh8N2/
orcjYUNB534Z8rOcTr7EaZhTMVN9B8wgl655+TZ8WaRfuKFXYDf9oNAXvvDmXFT/
iLfajGvkkkKWMdovVpR0Wn0pknrV7hq4h9o0Vq15DVX9YzHfAq8OjTGppTjlGrDS
4EG3MCvgDcX6LXVYeQw1JVtIW8+AUURbRegvUwRYjp4YODbPO6Jw4HZ17+/XAeNa
hhyo3WdjgyK+DubvK6mf6DIqCDoVHqyPUYXWbaVWmdACSsZIyyk49cQUB02QdmUc
N4GAotz/BHHNOQAOUsA37Wh6KHU/TiOFv+3twYcUjQItEmbFvsNDsQOugL0lawER
gfiJe1M26Fk6xm680lCrAfnzByFC3HSyNGTkqV/5SlchVg5KcKkMpcDYjp42xxs6
CZDSp5Xp/k+MkxbL0u1567QjrA6uscBw2vgrRURmawPwxnJwa5jyT/AO8nNvSuit
I3i8PltbQVb0mUeslc1pH+32uM2QVGwgtvLerQDRkbkXiDVF1ACT5vlatN7a9+aS
YP0gFYavzGpyYjI1A6cMoIpMVEcQLqtLL0kei/8pxc6lCGu3Z+GVbrJZhxoAAPVU
J7kSJs/m5ro3pF8y5T8vKj2m2SQZHJxsDnebW7s5u/p4UGQubn/vmCgXEy8y70SK
t5Q0kXV36Xp0jO86IAO5vqjllS4ADUofTzybGTORzitzaeo2MQyLQmZdtggX1aDs
gy6udyE9ICe3YqMBEibgqjgJFktIs9LRIvrVnejDCRvLxdhoNHbcg+lY8pS1tpf8
1yBF8uEhvXf9ZqgtfaLE7XMCaEwPGjNAw61PbYctLSPjXw59aeUb6xV5dHt4cXY8
5RlAUzoQCjgpm6ymS2enHhWMOy+jU5ywekX2b/BF3K6P3K8b78IuDIkijbUag8R1
aqPx5GftJ0vWAqgEU1/cZvxVzjrt7Q889d3js2m0b2Y7y/GGMBzOwhxrV5NdtGaf
x34fqeTGSUGivC1pyyTq8o5KOhgL4Cd0vgGfpHUnD0sr/apt0TmEPLgeFrw6osJl
75XbRKOBlsIBNMKePRUILWbeIAjTMyiTSbAbj0wSrwdkr/ykAXO/iHaPFJyJ8mez
n/mKEHMqb4QBElOShdVnOcTrDYTsotNLv/5XZN78YzT5HFfH/53N2lemtdcZYShV
/JAwunsrGnsV3cRS2t5pp5WSDvyzlepq+j5HftHbgsV5xVfhFgttQ5VhZ3OxzM0B
JOzkX54ZN9KJjQQEamdOKu0/Lkkc87X0immV8nX/7+cZfzbZAL9RiwAyUSiXcmSu
n6mPMC5V236GqDJoLEfyZFT3a1M6HD3iDMToa4fntz5IJsDV/ksEJio4/VCSJTaC
ZChFwJw+9H8nT/Po1rVg3lfol/Nnx5ZL6kPb9JUa3SZEEy4iJ1DUqtBo/+Pk4aas
xtS7nyfotut5YF1oWj+36qP6QQAwN3Q03Jg3LkyRsyH1DraXp8p8ZqC+fNh/eWpJ
ZJoD9rCB+Xgg5L1q2jaxi2ahP96/Gku6KpLnT0WA2APWmw+Z2tmDsFi96cTV4BWW
dR+LiaoLep5OOtUgygW4yEd8X1yxjv2Tx0svomkuZVXhVDWoRLnHZEPu7KCuh0X9
yvuZVacr61AK1CrusQqmZf1GFoSxha9qJrgPlYklM518sHX8/K1GdHA3YHd7Pe8l
UFMW3Wfm+5kal+ZdXkaDk723R3y4/9xVDTx+pkIsHG2vkJbWk0Y16WF33U4lqTt4
FbaXPq8LF6Vqvt7mB1S3uAOZkj3zJ1OpGWXhoBVJsHPlICMS6s4E+gyRszMYjIMR
BeW7+4MuezWbbXvTgxULmm91FMJEL/c/XMrAIUWRLKk3Xmr3ExVL/T8zTJVx7pEJ
d5Tds8MwhIm1T/dpoicYJjSkPs/HK6G03OkxI9dlz7NL0h2uTg4tL/ipbIlaprul
Lyn9EVP5VCAlIaAK5F80F9cLsCj7BzdxkZb0m/SUR5p9KAk0AHpZ+JfaDSp1UXxh
SVI+dk1LR8arJOZnMgn1qvhHo4Fdkq725Tk9FbhCZp5z6y9rGnaqtwFMx0VWDo9T
blPakxN94ahSWC2I49WJT82N5wzq8RQXzYRhhKXCeH7fI5Ob6sk6eo9m9Y9SNb4g
nBiPSI9M132KEDSrZCW2GsECndwepPNGSIcQr9T93N92D1cr6ppSte8YwdqsyRwJ
VsqprF7TbQlpWAmDKH54YhXaX4oBu+4Vh5KU1K7KsnpbO8Jg4brEfux5ldwU4MIV
f+oYEfJa2XrwB/zZ9C3Zi3UU1OeJaHmjPvZpXQe5+I++65MoXMpaqamqLr1shIg8
ObvQfryYSq/XXH0CMiL0G9JNsLcj55ldU1IKZKidBc/je522CkKU8uHRbl+byGo7
1u61epeaQ7jMhF1sBkRNmP1pfGonWXHhJnWE3c3Ho9AwBZo9RjELu8vQXm78ZKIK
kqaDY/Ua1zJb5BLPpGajcRO/rlVU2XsHBNt1U35B5AIEJoDblvftv5PekxLgPIgI
CfVnWE0+PO9YYijwtcbnj+TRvGCe9mkaaPaoLFef8dbJo1mw1W1XlFxHj4T9sQD4
Ere4689E4+iJdyT18gbbCVpGFlM64ZcGzCzga39Ke1jSriYwtgA67Yc2fw+WHiAk
Su1XAI1zwPFg5wkeIQsAdqb9R6sfaTDVVHkerAsjPCDzRmPGmUue1h3exaFx36gh
AAYhaBXQn12eJRStkKDyZqej/4Z+8L/abFdvD0J0s4OVKNa+kSbiMXgVpBfC8zRH
htNySSYpCCXL5zyADFJyf5mk+fRjz1OcBJuw5sb4uvccNGV3rok5Z0bUqwt5rnQn
otNviV33WQ8LwZUwAtBM7jQ52D/7dPRcAqhU0/ugmvm43f90MRwToNBRK4WW5wye
bEHrPpd196LuK2Hp/gYPdibm3BW4sYBvo780xHEoxYJJT6AMg0FDa75t1uUpnQvz
268+KZQUzjo6eHMoqbc2t5a/u/HGa2V2qDkMzrOkgUzgm6cm1CODw38sCcvph39I
rLo/p1vsVvvi9VSm0V7/BK+jFTXLezxGxdkB0FegH8eEV7kYU9zeGbR0j1L/eu2u
4IJNOiX0Fpe6sTSyn5NurNAxEff+PAb41g4QrWRdQx880MJt8jZS7/iNxKYjvf1q
CsVR6QY6BkCZdvQxPULABMB/Y67KBs4bkrFWdUNFIQBM8MfbBLetMxTmustK4n2p
oSSWx8ESneuLZ0cM6LH/T3WHUSC5deZXdt7oD3mBNz65LD9lxejcR1nFmG/+CDOo
0NKAck5LKs2vV60J81b/SMQKnlrjWQZxswS+RiwjSFTiYguPYXUuvmsUxY8L8HfV
DMrdJUs58jfbvOIR+LGEcnQ5Oukg6CZoK8+a0IGpIdjLeriIJNfS0Q+6fM8viDYT
wMJatnpU+s/l6/JTRRnKg0VrwWb3oowO8ZD5mmSLjwLGSohMdm6IXtyCE+QxYNy5
z7WZ/ZqbxJAZOuDLBMiE7Wnmdh14CI3Onphaoqgo6CIQcMf2tYV+dmkz1dCYcbcO
Ysuu5eYJSnpjF2PC7tmZzDoNn/qObz7lKG7JfAzy8tJJ9oBzPwZiMgYZCvlKzKy/
HGg2BAxEIznzOJ9YxzZlraIehUFavIHJ2DcPt/TKYE6b08E1CUEh6NZ4S9Wkd65L
z+dy1raqtviL/DTcGpnv220HlTUkZwvtWpoDfAKaBUeY2B3Gzxq5uuzOAYdN3hJA
vCFteFFg9rMEa7jcjKQ1cefAaSY4TIHSL6U2OcbK8IXfqwF5y3HBEGTH4F+IygcF
r/DYHNQwLHmRFHTKN5DZYv90jwYktMlh5yOj9AiVVvEc7pYMzO0tGe/nAna8sH7b
3ZvPN1pa6T7Vlw2vdEnWJbaKPlFj8cYPF04r/a/VVcPu5jNsxblc8w53NfYJg2Bf
znYZnQWPLWvLPfcU7NiDQbUaIiplGv9XJmbcR7rsMV7Vwe7tW/dBN3ErX4+tTeW5
walyQqNqUSKNUyYJxvEMOmNEFhUVxagIQ/NG6RAOBEzp0I9seGQ8InmD6JF972ct
L/gX6ozGWVE1aNaUaWmceHP0PRhRROklQ8mzdwVccLiJ55wwtg3DyFTE3aivj5eU
MTrrIcRhuG6uOFB2x7p+T6Xy+Xk1dOfD/XKiVG2p3f44u1/ss/2VV5qLOdA20I2Z
oMCGnxsok3cPbXAQOSdMiSeZBsMFsM7/eMX+KYN9+Tf/o1OsVXUzNoqynKFWcCvH
WuXoSdGynIQRk0ob8tbJgxVWu3IrJIaC5dnLvDa/GpPMQNCquYjRZU9XO/9bRhq7
t22tC/3FOJ+zRGBoxoPSYhWYV8MFa1If6HyNQOKtaIjh6L4wooWosSrLg/N3OHlC
DCBtgRi22eOZM5PU/A+84j40P9qc32xlRA8HtYq95i71g/9SwODuQmXSTutnFge8
JMXixZHSypr0qTMRW2STgbotPOxyQXkhSKe2D6E3BDXPrMRfSBDWRWelZQOkRbbt
F0umN2avc5SMjvNJNadCesS9fF6Z/Xh5RySV+P1maLo1z8FdbpgPSW3mxnBhyxbN
Ck42wNfxlsUPqmYbgoESKgBQVp4OL7k7WOzZPvhJgrpY8XtexgtlrIO8qynBaeHY
QX2SPCnHuAi23s/ZDWbjp1RWSYlBTWpRq7eTTyc9mwE8ZUJUaoXSVJFuktUxjZ2C
p1/s9iefCEJ6cjEzs7+OILgUgnqmS5hj469WZLcJgzCKtoUZM75aZa32GviqhnFQ
542SnAdVHmza11OByLiCJB0F4IfpROXAOJvDFqgCZt2GpdosNoo0LJ+HMlyo80ei
FMxR93pOQznV/2IYhHFwKHAnpHBCrgb7UD0XCzMuzhhKO7RaWXmDmCUI9SNnb9CZ
z8LnKoX11BNaGGoHkespZSO/ubaNb+wON4N58AIoD05kFATM7Ow9O5loDcNdRKq1
FBuF1PHi1ref8Vo7r75WSWBJPkXdB7R0CXd49yaFqFEP0XbJ74FPz85mAm2zmryL
pgJxF5Sxuj+fxlnErNPgRiTiQvoh8g5hlWWTJ0zFP6fg4i7ATz+/djaiPxA9eYid
OyuuSneFB7mdIc+Sl8IUNXndYWHboMIEdCNtfV1P4MoJ2Mo0CzTwwiZDJQwFxPhO
yYzsWJy1gfhKB/t0U5+V+4+F0Mvx6kTC+eaUBbeq6TK3fxOWNR1IQ00HKctZsQRw
o8aS8XWq1uShaItYGoI/zrzhmo4JSJe/whlGJHBpowtPeucmxS6Zl3KCa9WqKm9L
vSnayu0ivQr2Qm+0L/WtosW8hbsnog+Jh5gp70U2Cfd6dRz+f8y52WwYpjNcbRpH
lBUQ14297Lvv21e/GR4p6HiViJiKJRgWCZu2tMuFzWbrT+88JmOF1SJIu9KcCgP3
FI0flV11z1x7hmLOCCZrbuH5NmCAmb6UkN3+R5+CMpbg4P/EeDQVMQDAK1KF3veu
Mqb6EH/dJgNCiQm5nhRStS/vazdjdKAsNkTUGzzQoPaTGOLkKZ+zp4IXumqTj7WK
G/vkmNDrJP3XiSGLbZcsFWXAanHkXAL6S6HdQ3pkAA0Y1wWkZ5aWvY/WDhbpOlqp
NK3yCouFlGKcm3tTKrYZve36GpHT8FBwakyqRgTNCyu4Ti2Ri1rMnJSyn0tK58ix
DTfrkb9cuXjRsgUneEXoWA26iWD29mSueKvJRQMC9TxyC4USPGuBhIUHWrH3ZS7q
fIIjQjzt3HQ14qy4W6ckrKDa31+eFTfZGuoTnaTMD4djR2/N/nL3tH9mlbjE9eNc
fq6JVszKXhvUnKnuH7ISvCwwCQ3Hlb+ieqskHeOezJJdZr9XBPRd1QBu5RzCYqrA
BPuYUCJJADjNC9smcCFlmJVfV1Swj30s4a9e5KJbadPuG4rOGXdrlxaw0ce1P/ps
TS6IZc2Yb1UBB/EupCVX1/M1YGA4zlEvzPOJhpgy395vhiIRmQLoZIIIcBqw0TRm
2xz1uofUSAjAQI00XUpRveIZo9YCQM1dFK09rUctpgGl/sHITrsvm6NILmjqQrwn
+fB/1lqMSM1a4U87/0w2gG6ixugJgK0PtONm76fqPjhhoEQ+v2TY2HAZ7SvEmbVS
JT5z2y228Zk+ZQ7EVg/Y1wjWEX3B2LKVxk2/BXZ5o3Pmj2djHxBX2Z9RMtlY2bjW
FO5sLYRzG+bVXmLw+hk/1jwIFEJ9Otmz1omZflaz/iAKUO7fgxGZQ2+XOOGhtApE
PE4dJOkD4GpbXMy0XFqa0gSGVG61GDSFZyg52HwIgbOmfGKuT6d1WL0MmqszRgiw
YiuYxupecZds8J+sNzz1VFFiJP+Xd+nv3DvH3K0+VpLUBuxnBfF+zzMVtbYj10Kc
8Bvme05Yfyp+zAL8xqEEP9jPEOcY6bYLZVtB4guALiT5ZQKQq0SC6Ntqjreq21v/
n3wj5YGDK1ojI7bbc7u0FG8RkPyufbCyobs9o8n/iLkAyqW2Zb6mjx4IoxPlHkpC
oAvW9ykgqwoabXaXaumEMPxHvlHPrMsb384gnAVBydpKTx4BkZvUpNTCFLiAzM5e
4Gb0fDL8qKvAQZDqeb4PslYWOEUKFewxBWOL0XO69ErQeZpExddA2oJWtbPSBN6I
8puK3Spylf4vX8RJJF6KwFD65U8j2Xibnu8Ud1vGGSrQb3wenL/oGIIgTIHTTYYf
itmL4zrBCZPjz2qcGx28wOK/ycJGhioIQchCoI6tcOEI35DVNlyITwSWsRyCYei8
98ZdQ5YzAndlfisy1B0FrKII4SppSWnMlH0l68ml6d0FSw6O69spBemUK4AtV0Qk
2yxbFgmY5JG2cgn9sed1zWee1tbTHsl09ec+XlPs7WWa3RbgwnvyIc3+3f0F0oux
fblbifyBIwpZkM1+j14BKGjK7X6H0pvyvklSd2yA8Re8kEwXdcyr+ZCYLl24LEAG
Gcw2LKzDWh3+K3qbyJ2jHCAGHhqib0kdHsEWuQtjKfBshKd08VRG9rzFKwa0mKK8
ricJTppKAG29ejy+qYXj+/Zok+kuwcTsC8ozjyO56dLzt+azI7OQfh8JbHcxfuY1
vOV5spTjEqeN2clIMsxeY02HKxQIDZxxqpPEoD5C+fa89xJDQ/LNg9t5Ke4JVC5h
T/piPPmpyAv/EVY7GCaUsQVdBA6O00G9Fw4BoDS4Qq39mPKA8OX0PbBw3Jd/DSjs
/CwZLRziCFK1rIFbBgx8ND76HgZRAyYZlfXnCBR55/hkmDmH4jqyAFnd1r85ZZbZ
zjBzr12xK+grCrGwKJgvB1L5jaMLKbLwjeuIvigClDILfhYXcd5s5X8zd+4s/kuD
aYg8nGbTaMBAaA3PHjKljZUPHSkERvEZALlmrG7l784tsTsO0tWZynK95iPcrI5D
FRtaLoQrnyIf9kOHFvBRWMSHd+z27AtFBll3l5dqb+y4qJ33+1fVLoyQqgiNWSTG
NFD1v35dWPcGefaopr+ssC9NB4MeIu/CgigqrKOzQAD9XzLeZWw/5Qb6ryLt7x8M
7epkuxmc3uhp23i6WLBncWRQYMHzNfh8pxJmAYvy6ZE+suXxRTDYp+HECbYE8G7K
WW3FvOe043og3QwA954I9nNB+iNNEIKaW0oDO4g+TARpYWwI6KO0fDqtY2IeUEPQ
aEhmAMjUMG6ruHSFjVYU5B4aGLboXGe8lKfI8iermj+EUmvtV7SO7CHlLqdcUN4Y
uR+I9djQS0NXhrlQmuMiNrijZKUKEaSas0FmUTvDjD0xSmNPaMYnbLn8QZ6Hqxy9
EpkygMGfE1jCryUQ2BoygTis5/6at81J4z+lxAzNLGiZkWWgGc3WV7LQMsaUaJo+
z4Wz5KXhNjRpuGdzQyBOpEcP++tAYOm724qvA+1JQGR/P7hezKwm0wNTdY9nhHaM
lfcuhM+yaH5T+JKPjs0GaCZzqsk7gjDqjHPFnVzMnugk8jqmYZV7nxcYwlX9mug/
FDp1x+Y0m6jMJsnXlciIhoxWIF7eelpCb9ou7wyFX8PBFVE+vVpb4tOxhE9Msiwj
KVLdDShNK9sMuGchzpOVe2GEtTJOetNCVh3xHXQnqW86PHdrCgPyKGUrZjH7evyb
6FsfE13T81MY6RQFBy9/52VfMqot/Dmi1EpUTG6fKbRfvQOCKwH/cWi5+IPmsBSn
Jv2/oraitmPS0BCOHuOfmtYrYzIUprKVZgPfdbtVl+LWEv/h7EnpfE0P4SEpsM2X
AHVUHhnT1PySgbhyeIEf8KYWJk9CUVvaRu1pg7aLEM/Kkme8Kf4l85P3mSgAymAT
U32oahxevk/MXqh6QSnvZSt6T2RlYRDJAswSNWv1DBAwSduXT4genWorMFs0Zwpx
vrr+UfHdCHVj2sOI93C18NioOlTrc3OuyYARWUKs+XdT7PgmUj5RzcCmuDsRa/5e
eJo/ydwSNZgwP9NvMYt4OCcTUvX59gWPynMn0AkGheHEH2vW2LsF5ihPitIeKUYi
wlFwM8pK5bUA5EJ2eaDk1zlt4kAwrJV53Wo3t3Wul3JigQfe8sNju9XLUg5/DhRN
0xpfoZYQySit8fkB/0yKPJ0V3Ou2R/doXM0tvf4P2ouCIeq/rkvneMsOLJdV+6iO
vo2BxsIB575a66dFiO9IdB63LW9Im7KNdwDsOzbwudytSCVVVTZC7uMKQT9xvv+x
JrczyUG2hwYb/7CF2IfFd18py/2akzlQVhX7YCYk2zLWdABlARCsLEAtg4T+qiFO
KTdE6l5MZf4ZHbSRKPisdI5sQ7AFKcdjAVaC74iQSLYYENG8nY28G6QQGHTGq8Ot
J9bvAFXM+tUCfcPGte30W6N3tBGv+CIeW/LZ2DfKj21C9+xCTi+eS+XsMK1F7mbf
9HMmfr865nQpJTT+UzTj42pqwag0uFs3FIBaPq1m7PUnl8K+3uXjFhPO0t2T9YSH
ArINibSsGP1JIx8JhmCyw7BvYc/uZ9wdSkf/HWU41inWjDPGM9T3p4peD8HT9h2x
ODxsmg537p/M4aU3aXxwo8OVe/OMr+++kdWIULUj4/lBFT8SiArLmEqHPzOGMq1d
JKeoaRF/qdcFoA1Ve0JdfUvKUdSkQsam33JGf7tQ8+tEZB8KRNaHSYeRrkiLxMZM
IhB3xyA1Vs9Pfcgeli4gLjhDgxTDjKJwAC+PC2fVQYZUTzwu3zhE+19QpKOu6y2d
MAinizZL692lDCnz708ahDIBVSqBQeWG6LjifobqsHzm+bnPvQxPFTaVN+H40eFA
PgcFTD6yMlpveaFH12ugk+YVRkA6Kbo5e8C/vbDgSzDdwkurWmsAM2h7qE9tV8NK
nhH9MZjK44pnvx5m6EQGd/K9jk6Ri+P7VgJniqhGZVRdzkBlBzk0bZV7jD6mLhrz
Ee5wq9bJnCMW/EE1s3pyQqwS59D1MMyxiyJobLtyeQ3oHaG9rWx2c/dtH4AaWRPm
HfehF+shGpyrSGOE1GLtJRGfuKkAl1vs3XEGFpjA0MzThwXmcJHY7sEGgWSaogCZ
j81squHPVq1cFelZAT6Cj9NjvGvBZlSUepbKdr6115EB177W3dEDRYTg9hGmb7Om
krlvwvZMMf54Y7n6KfOpwje4IOtn6ohr2J7qz1o60iIvBiHe2eb+ae5HqJs46Www
OAgTctGeXsKorYZWeL/BPB7ORnicjnsH0VF4H7cCulAL6t6GQGfttjJ7uZWW2krb
TyAHKti0io16BXGw7x6EwzNSusVsIozS8GWHpa60YMHyGWFcsE+5mwXGWDAmqLUN
BJqaixyCy9uARbeqnqpvUqoO7MJbt6DDoT/KlswbhhExiPso+pg3ruZ3fdKaLIAT
6DWMXCrFTfLj0CpW/9bQyIyto+UQL3OQYY/2JilgV6ZYRaJ/jS74y7j1oGzMSk9D
QJl0c1jj8VsXLFaZXsoaCwSr6JJKVIRVMuEjWFYwUojZ7tpDR1g6S+VSJ547gVv2
XmaYinA3dkRIdpdJExQhSWJ8bTlpzFDwYWKmZ3pRXQcFlJIcX/adGB92zMwCOit9
dY6WML//l0IQdAJyiCLRCe41X2xxN9/OLbtdjKfyqzC3zG1HI6k9cWlJsV0XKs0B
NYEZTExVx7bVoaRQsuL5FtKFVeNOWJj5Vtw1WeLUfsfI/YjqJ+moTKz3iMWrrWuT
ns9iuYls9vcL6DK3+4M408Cb48oP4BpjXGcDfxuT8gFAN8uf+6Kg2/zJ9hNSotXD
8A2TVM6qEFgGlewkWslWxdSHYHK4M/iDFm0ynWpCVDn96AobEJCmeceH80SBs8kt
8sUzw3e/GlTIzell7vsijPdqN1Lfjeu/oxmQ4uOEHpqu6NU60yWBW949BzZIDtJE
Mqdlm39CMLdGisG6oWCjzCYC1P4gGPNY+/c3K8E69Lq6oxWfJ7iMNhCV5jpFy1R4
xze586S8mi2tHrQQnN6xTaPbjG3vTE7hDw9tVszJ/aX3NMI/j3b9hXxHVcr5vRPx
g9B4O/7jf0VanAcvb0DsGB3orNmRb/V9ctLtTd4JnPvx5ECJH9G8jVmziOIFvZc0
w6Tm3tSAGpLawhnoXjBYejMmw6F1C71GVJoGAyrsyeR360Gzc4By42CzZhgHwWo7
AS8w26qZMdVMBJRzQ2UR4oH2wck2UjVSCdQer/yc3o3PklMzf6bwb98qb7mh7At8
89qRsyK3pELGdk1+eRd9XDVGs0GN0HM0EQv/cK86rh8mFBKJIhtofxivAqKuC5xj
pUFBrxy6e8kl4i5eYa1D6j7wFTvezCy1PhFn5l7h+igo37IF0fJY57TznXt1x30N
qUcncHQ201RPI6c3qSc+EPmAXFB2Ific6Vg+hVkalWUCaykKHQUdlVNxKtHmCSEl
jMprlxxtbCDtg5QwmswzqTqrwqs2usiakR+iCjYdy8H+UjHqm+8j7d291IS6o7in
9RuuEDd5/kWfYLMknEnL5tpT7b2zM4tYfrqFHWx9askFzQqM6WcU9IbRJo3honZT
or3yAMSfM3rQmJwHxEBR8I2tDeCyjWJXosYLS9nxYXGaGu+boE3u4ax6MwChNgSx
Rxed/0FiDUz54ArcSrUQ1OCXX2AFEjUGk0ldwWOX/E4lvvscJZ/IkDI2d0iReHe+
83a78Eh+wnfaXpJ/Dt4FuV0vQkZbIB0rYFhnJj3J4pqxPldVZ4KAM+yzlX9hHcrG
NNq7t9arYgz51yE7N9J2ORXNzh7LORcy4qZnn2K55GY/uTgCNJi+dYZYyZEtN3zC
vVNRGvDJ3BcPaeS3X85S24B5pDUa7LxVL2hLJ4xFlTcqLFRWp3n6j/hPALfyaIBI
XewcTEkXVRRSoA432gYrVVSbduNmrgH1HlGyxkA3fEasxV52IgTJL6vfw2sVwpwN
joGBiuFhh8x/4Ci6lHNfN8SpVoVs7Dh5Sv2pn5tW5/nBUh58rAJ2TMh4ZhVasDBc
0uZswJlEMzcXNe5kQtd89DdIBL1xJs+OCbC7h5qN0k6os76Ubf6mN1ZVHurEygtC
sdAKRs3JKAXGtbNGgHhEYQ4gaISoqPrrlGDdpFKZabwTEEjdfzBhdr5OLhll8JPf
vzYsCIsZmC1rmPhmgXtUalWxR/2PwjhFKg9EqUSTtwlIeStoDK5jo5yNVLGsfGwU
Y4Hs1SkbmCrctsDrDJrXNyTtGpZh6OvCs2C6cDQKS6x8ynhO0MMBeR5GUDAiuj/O
VSLHGKIJG5G+VQLbqPxfLmTIkYH6SWvTBMxKyYJOwCn7AAhnxRBw+IGHt1sUK97O
2pShNotGxlJ76j70c6xQNggx8D8oG6P8tDQN65XRx7OA1sj9WTUrEOgT0OPMeIb8
hUpLFq57KKYVOq6PF52WdlPb04s42xsgIUg8Rn1tKxSJu/uowz53dQpVfCWwCW5J
JdU5cnPsiGWbZ8by/hiI8oxibmGnkV0zDAgpwI8DNcl5Bf6IV7O8qWS5O8N2QtkH
uH1GIIdVJCWPksEGiCxhwr3FBIiswl+BniLnIcImQo0ZIohcPiZbQq5oBi5Gk3lz
/LmbD/BsEO4K2thpC3VDBNoJVIM6ER8fl3eMRZczC7YzWkqKbvJSNtAjSh3jSoY+
IlUKx2jcyaY3L3yhzfM4QCIaAIIN7FBKWFaQjifDF6D0wWXDk6K8GrHD+oKzsZN/
QwxfV2c3KLgAcGpiA2ef5D3pHomUKwpBuxg6vkDATt+gcoTgMs+cJ3hvcIMhCtfa
irbmNZuh2EQnBNlk4i8zJCTDWYOLxZRWCbPp7PjG9rDoljuksGff11GEmdshW3Qp
gmbxMW5OB9NPN+2I47BWjHeM2OuSB6GYRM3JnZLlV//sQ/jHRLLtNhBROptmDUYU
s/OF0LLZzfNAwtMhO5/CjgZz5wF66MzCugnzqkbEz3+7CZUu9FghnJ7XHHwVjbmQ
LIk35LI34z2kMQUleGaA5fefdGuYJRJvDllbAQZouH3hZqi1U4MgKwwzdFnfphU2
HmgKELHOCqjlSuIVfPvoeTvrAR2l+KLhNDgRQJk0dA3TaAF1I32h34xBb3YbQQ4J
ZnLzoQrI0U6ox//pMxrjuy8E6gEdZR5dEtvZDzSkt8vfwHGb3eiFf+ceLOozSgId
nEhOFNIglnL82O5E8nysowtaRH2Ew8/0D0rzBz0ErXFqRBARbwV0jJzYnePZmVe4
GXXESvXndtYbSO+KBWFvmEsCVaMq0t3aFemQ9UHIoxV0YMbG1wiIVDwYdQsJOmDl
57UpE/ZkmjeuOEK8KO6Vfe9V2K+s7Ql9t2nmuWeyzZvTe0QQRJic3/ZkA+6NuP6A
r0EkJntiieI38sFJ5r1evYEhPz9sfb+4z8oQ3WrdYaLVVilIRvghFLpyv7bX8Isv
OJyCRxIO0PY9snNCEw6I2Zn+JgkhPbjxj50Ix8uWMieuqTIR/UjWaFVijDEw03Fq
xWDn16nbNZ1RQ13euyn/b9jj6j0cTWJK33iNyoWgpEbgzUl4QU3L7b9xgaTnDk73
MpPvEAEumiGNIuCqJa0oX0UtH/ZTCB8fHHcI+JDDPIJTba1EDftcvasjqxlo6Dqk
U+MzlgcWiVwodumDaUV8fxEwvnQ1CyQytDFNr5FbJZOI24A/V/eEyt+8ZDRgQzRX
jG/4CGQxs6o7xE9DN8XLMGmPx2HQOslleqh2S5Wq0QicucDbKs9k6JT9Gkrd/q6U
tCMzhJXqE+3IO74epouH6HN0jiI0syrInJjLo/kD428uJll4tyogg1W8VHNZ+yQ1
7IcO21TVucokIpcKITJsQIqwIqNtZDIpec7iGLtY/pnC8nIz+PZkivXqWqVAb8DZ
z3KcbunzMcULrLDnuoQ7Px4YufwI2bfHJqH3PwCvhkCKRzSbe0eZjcvu3DqyeJof
aEOpACxJU+9gPfgIsnMA3zbsDL8RwILJplMZlPzkLcRdJBW0GMIw2zwN0ey7F46F
RsnWZizdnoMvQ+KBOXotlKwWTunWystE7rVZZ7Pl8aw3ShTS0cnpk2IZIVRjBFCP
rz8gTVL9n/epj6PakmeayjI4hutXPP0Fyzvx+xP5cqKfxhfEn9D5cTamUxxwun5Z
9tWvCtI6JTc3L8rI8ZZoZFaNo7QBv05NJpfXpZLgkvm7lFAREPDcrHOD6/o/lE1R
6MyOPBPRubR9mTR9EUlUF+Jw9uZQlKVOn8Df62LoJD7HGDoLeGirY6qraWk34v52
yuvsu+Sq6IU1kWLULKMBAnPdX768GtBAvFgU/b4eEjEb6PbWK2n3XpGvcmHLITIg
Cj/Jnht0T22YlNOqrzrBKRhDvqAqdiRdim8eIFf0VEw/kHkviC/8C0abiOpD9+Hm
goNikUfoPphXT3rWoMKA7wKo0j+U3LALSQ/kFL2JjxIU8XGfykbkee3Ddx56ria5
QmC66GF1a6PFBV+BkP0uIZiasvokUKYTQZPRn4dibausJqhqlUVFN9aElGeiAwY+
/UW6rQPmzXNJ4mGMCZtk1xBQh8GW2a7KTcy2oZetAre+xqpODb7x4yZLC3OPlrL2
FKE6237y6gT80LHxoR4ylx9I/v7yJS1k4gqrkTMpNZ88VIJZ6YE3bAHx1uu04F7i
fOB9UD1pmGz/kmUJoJCiJcA4q492qihnR52GAeelRLlnFEF0P2FmU9CpB0PkSBON
ywzNTDNQsaFaDAbjob2xq03GniNQMLekL+AvJovZOuZGf7T5+VPmqvOGeDV4rOSC
OLHcmuD82Z8kfWC2eMqe3f48qIFAXRO6F0sbhi5FNC3CRfFrL2eXr9TY4a8+s93c
15WECLrrUeFhx5Gi3rP+bvo9UD8IjM4C0GgaBmNhxOZnHPU6sOnYjDeF9p8eIGHv
/xBl2zJys/KGLtmjODfsAoVCj+oYaOO6OpTD1JtAbLXmTWeTs0DCPT5Nv2Hu44Zz
iH4ZHC2kjm3wWqSyWc/3kbYT26Tl0cJMsxRj0Gl1ap9Mr404ytTlFH2tMx8VmOnC
zh9F3zssFQDWVmyRkLS9ZDdhPCXxB++pQa5OPnQXK0dYnNtvlYTduIAY1e29LIb4
1cot2lI1Nhe/yw5hMaVTJJ5TPN2z0bdtxyqhSJP55+fiBK1jrvEUhvWoX+UCJ9AV
0DkH6dtJDwCa/Hbk1RwwUHvp61RwYPdd1A0U6pc1fHUctw/yNFtxo7+lHcuTRBVo
6BszvdONuivPHOxNK9fOPi+n8wFcJcN44glKdFZt6BMai1Sfyq/GhzaK+yw8wpUo
7r9SqXkPlKUj5OcMS8Uv9F+J9PiATswmTYmHOF3DYgq/niiNEaa/aFNGDeM57Tng
P6yr5odaLTdqPqD8DznUdhcMCEqpIhLbMNDblodS5foQFiA/06PimLsbdAJwIhNq
iqEOFLhXxZ7SRSdOdED2Auv/HpN+gfndRjnzWvyRaJsVjRT51r4aI0gn2w1OO0gl
C/WPswn+mjQigIxxCCtBcDswtPC6PcJsWRQTV+br1pE6xcaE0bRqfOgs5mHpWfdZ
VwTFbPPg8AzyYfpDW5MKG1OIKbOHq65zRf95Kr7/r5Qz5dGoMvu0Jf7NsjCxY2we
3CJ2fq9BBU7zOC/d2OBAjqBjTc/shFgOAEsdEYCwKwSipDriDV/7TqMHGQbAnOY6
RddvREbH3C6oY2Zwppw35PtbYKlWXlXrZxXB7uvWKjsfnwUr7OzxDa0m3m7n1UIO
G8lwUN2lECRE3ymggN/od4vS8Vl3FgwwipVHWqUS9Fyym1Wrz0+hOws1oj5KKpl3
Iaa+Kr8RhHVRaURqtUU9OlU5mLcwS2AQhy1018U8uohYVKbRbrciszcpVOnSoa1i
M+emretxGvBJM+rw9rb4TMUMUaxxEWJwTssCOLneRAlrzyEjdL+9bVBLovIs2nkR
OoqWnKE/8lGYcU1A0OiiueCdl1wxP70yL1z4thX7JHTzAgeCAF+HXOhD8yj7pyGR
24QYaAwItPh0cSq0cEz/Vfce6+wG5ve0MvEH5QAWRTPQRklyBPD0J7Sy4xWe8gVy
WjYIAlqinEfQZb8V50w98YDnTxKrOMg8WoUIM2VwZE6bsNV+BTMPxq/N7hQh/QoA
loXe8u8bBtkjR9hCcu7ccd+Jel1UlXS2qvSQYOjEl+YKOZi3yy/aWegFd8KEEBFb
bkO/AdDdsvu62jzUfEjsQG98bG5e+ggHNYMj0sTc2PIGlVWXYLHwVGr0cJrZuypW
WYO61uiT0sVDi3pdpyrRRdDmRRgWA4rRHLymYM4JoflpAHNnwjgJeUspcUTp8bEB
ty3oswglegZn8uda2zduKPGnbhSOe3lIcB7bf9igRFia2AiRja3vLSn/a9HtFBE8
IkBEQ0LdHmHJToaBJKAdyCxjScyPZjSyW+fBOApgzxpfUMQswNgnrxMqQeczDEaU
j7d2s1htUBDB9tqkJ5um2ttoReYcbv+kqMLEN377g4G6zUDsJXB7ra05ny1C0Jqh
H/+5wWdT9AifFOcx8hC+JJfPRRAyjQEKRXMKQjEFhEzESsUME8M5lH80P9KnP6Q6
7qMJx/e5yisYXyXWq29trOM2x/Q0OwatvhAEb6O24tLLZjlO/popFzR9S+VKU0lu
vIyqroWmqmSigksE4N8Reypbb8KrIz5O2uQ3ciBuBdnZ9qmZfZS7HYfEC+sYyO2m
I4lJJN9TWe2aNSQJssaxbeKQJ+vZvs8UPe9xK4lOJWxdfV6twqtyoJVIsoCzgp2e
QyZD3Bj6I0FqRR1p66CvCF9LWcXwACRXOCDRnbRcOLq60dSYG3oARyu2hNmGCg2s
bBkhotAPeKr2CoAH3mNRtn7j5NoqyLXKsw83dkIi1xHLOheFB+pgFgtsMnQ16oM0
7jVJJ+xShIjs1+GMq8ofXRH4tgH3IZpVx5LVghFcPYCX/2c8XDcr5a/9vOZQIHfY
dmuKAp6hMoRUvTmq6mEPWbtVTOj3+gRVwiROP0D+hTjEBdYfAvbtvKm744QTmo2M
tKj9Bu68AgaoDxv0Ny7ZKiNy2JcMgQHJf5CwmCxooyr0DVOZK9qOtxsCGb9B55XN
eF434ERKDLvUIEVk43oI9dReZPR19dWJcRZotByJJxJ1pJ2Ani9C2YZdpFVS+nKw
YQSKM5eo+xViS+5smrhYh6EJNFjZVXbmoK3VEnDkU3zh86FktgUh9Hnex4CRvaMV
93DkNgHOMn9iznIifHpoqeSTiC7tH9mIBSyLrrErLVW40BpOFZ2jeKdBJV8fQRwb
31u1X16QwB2gnwdgzI4JYOYnW15n+DDZ2Zzja3A86dhfGiHpm2w/95ROxEtervvr
mN+VPHIGKgU2dCD/hpsvG8Tqx4RUtH9p5XtomptFQtpQyRjNcjSG4hDlKFOc57ZG
YTtgn5IDujrBMYIttO1d1DOesGFlmhRBDAhjeL2jQ/djRUGujB8OOaEv4vkp9UrC
AxEySDcaZjG1rqL2thd1b0x2M23hWcZG2dlhDZrqcQAwoFuTO8itTzD7o+s135Aj
lHsIxqDv14x2DtiWhI/ziqBtDfBwHZyHUBS5MVqOt582RUfWLVLz7+GKbLQSBxhG
VcEL0SMX4TRlFsv5JgE4i4CvrociNln5eKZg6Z/VCvyPfQKPpNx/dXzx67K+h3ay
7BEcI7ayJiT9ARdJaw3PgUN8iuQaUyslxolJunUj+lrnWwThRJYMCRDpaP3eadd2
94Lo8KctnR4wLyCobPKt5VH41ALXUSmmNJlo7Yi9guwuQVoGv6Xasum3iCP4n4jU
sFpXxxaFqXkLKmSPPsV2EPnVI13JLe8XzSjBwSAshe/ArrsSj8OBdk09Ztg0S7pt
gdFJVwaTUGwi3yGV0k9I7xoQ1soAcMKyzn2S0yduwVzZQ4gFvc83IJnLarfKwbFw
EmggTVOg4GyGgChWyrLoICtysSnhMo3jdYvL1CfLKdOjztQGHKjq61qne6iMWJb2
Bh21TcCHxKIHHHX91wG+ntO4Z/VcEXikAm5mqezQjlEWew7VtapnC97Akz7l3MS8
8mZxbQjV9RY9iFbH8kSujA6daIBQRvDZXLK0CvltjGp0kkG6D0s7LjacLqpqeUQu
BVuXvWdBfAVWq5ii2QVQXqhVRpGBEJ8Mj5jIu9YeyUoh//4B30l8FclMxCWYKlmj
dDX2wKjGZlQ7Nf0vHmmRFfKcXxHRMQ/T++A7RHqSIrsREuK/yJ2AaUC/YU8P+B/2
DPrceoy+LEMfkc82wsmitHKlMXRKp9rXtvnJn1Dt4XbCq3gI1Ln71jdg07PUPC8n
nPjcTDhGUbD1N2avHxewHK9u1dOod5UnPnwgPB7sxS8kIPbg6NXCWeCHlAs2CL6g
y8Uo9WK7MtTykmOEUfg2WIDEIyP60qaPKHaUSap1usR8+0iAa/PqAeu+rfAh41Ie
oBUfUlo5swZ8fJf/HDQ0QRbulHHBXIfvYnLk4HJnrrGxo/BQo6IHl4qLy9vFcPkp
NknGCitQ/BRTrdH+252mERT+cTSRdaC7SDWPQzQDZVqid1WLCFAzMKfR5tLxOyJq
GfOJqrUK9mk2qlVVpOBdDeRdtw6so4U8i1fZGWpUTweETjXuZ8Sc2lCp12rCsQgR
5eXdu3dfRtCQYwAaC+OvrUbMkeHrMR3zUlxfmbMOHiDlWHIuKSsOg+B8/PP31W6E
tUnfvZQXf2WX3S3tE5lRdU5aOZTOQ816QG0bYRA6bjHSWVY0BfZnZJIl9udXX/cf
TB7G2PBjVUTucCjaDzIIXyK2DQQzt7HZ3ALKv/gCMszXgUlCI5g05i3WRXUBPm9S
M0bL9hF9KKjzQ6RCKLn/wIQipw4Xs1Ipr/8aTKN3l4ao+PX5fBNesHgWZudxDL8y
7I8G933HXnlDiPo/tmCbGnMw9AWc1ivf2Xi03cEAkdrEGjTnITAVTkP50iHxJavT
p4xrRBFIqJLTc5aJVsY3cZ1ZEODrX7EfXVPB4ZUrPz+YLYalrms3Zz7U0vImIRWL
GRaFJC1vjDmaiyy5uvz3aXcnTCMTH9PFfsjLXqSgn0fWNbXyFVArqD1IF4Lb6Fdd
W81WikoOAPgZoao6GiSGyed/24RtI4XNCuCXtU/x095aZeSJPhdRYjHdYiqmAyUy
pCfQNIUxxp1BEVSlc/FF2RjjHajfKQGStbE8lCla07/na0Xy9Ivg4Rznqh9bgeWz
DQiOATVZP7W95zy8TpScswCLbaBHIYPn5xmcraxEdn/x64OPI3uUct7WC2xZcj5h
Et0j/JzFf1gbyDLIi/PTKmTpJFnLarFEGhL+zknHv/Rev4P//Bu5ieXzvhsCpFmc
XqbrKM7GE1IOqOJij022rE4wDdMhWa0pbt3+a5SFAZ7ZogOd2UbH32pUbgA9RmWx
MYdcxnOUlxzzj3RUDm5SSUWjROA27U6ikqENrQwixF7tcgeAC4LJIBshjB2YU1H5
yeC2RPA9rHQEZoXJrDEgxLAEHR94BZxVGcxNMngOnggZ6ITJA1xvWRy8HpFdlyrU
cqkv4SShIY/C/2NbMwswEvNkvts+NfWk9rJQMRLRdKJMi6UhF1rgM6IWQCGIkd17
QJ7/q87XKkNJsJ1q2FZVHHoME8IdaJDqbzUx90poCejAcxxO19UCBRuwuRbX6GbP
H1LZd39iXy59Lyx7v/rtggCMOocFsIJknJceEn2ogulq7c/W1KjoA5KnNTb56DDf
TBqtDcQAQOEVZeVDjiE7oUp+a5YoAibJk6/UuBlzw+Q3rYdQ8S7SENCrwfXmBBA1
w27jsinAlFe5k8SNwUeS44LCN3JogroFY9wpXIHzmN9J2mLKWapsKg5sJXvwWPYX
U67KGBR70F1BfEtwWgg9w/PCeGvT2mm2fWnfq7FgFM+NIewhHddr/Np77Bt6Eu9L
ff4KZmyEdSZfMC+oGIqU+XT4QaHSucn5EAWFQFEOtsjO6kL5QJiLUaN1RZzHYccV
JVZ3Uxig2kq1B64+VEIvVKiLirB8ps9q9uTexq1Rh0Fk/oDsCtdlWFdLkNSOWXXi
vut/jVYCfHBj1btYpqatFBbaQb3vI+ygeEq+KSzpo41MYG6zGbyKAXPzROxxtciN
+ci5bli+wBdlS7HiOVU80PDZvywR5/uEgzEOh9iXa6dBDmQ+lXHuQr4N5KK6Okzf
ff9r+w/EBif1G+jcFBl19x3H4KsM3xWRpHlUY8ML25rpKAIVnTWuVuRe9m53KTDC
MXskcU2CMfyb2QqrpD9/ydapqBnVmqPtRta6r5UIGQAgTJajqVPSn9vm9ee/WjPR
zBB44aPE4zJjl/Z175y8OBhX8ViDT/3l3cpYnI/sP0qPGY8Aq/JbKWBzCFMcrAdm
nhW+pJBGTCyQez+HTGh7O+dAti6neTkgpiP9Sq3GEjxPMmMYfggfgqTMtpBBYGli
wjghwsUHIdtnmtnQk+ibiwIaKyUtrOhcPvY8zIcN7ybL2AIfoXKE4/tqu7ADuw5O
SslMrSgcCuYw0JHyYuQNzI2OVzgS1+coUtMEYAvhbFTcnyycJ7hSPBvUSFxDe83Z
XTBJfUndgXEpvqQuIVk7nfVbZ/LtmBRXgdjWIetMFSVvoFjswVdY3S3pRNiULQqj
A2FAUb7G8ZOSHzqneZSkp5GBBroe/fPr7ysg/lhxHe+93CJj8swz2GxyPYvj3Ufs
QXkivfbpO/Hzd3lNB20Lb94mUBt6VPqzNsDjGgzliOL9rfSBvNXmmEt6A1xDNZfA
ZbjewUEz9/EW9+EShQV6hBXyWCm933ZwKRmVfk1LHZ2nvw3F9JNyrh+m3HSLmfhA
xyTR2nlTJzvO8kSe3GbGrp2/90wTm9xwI8JkB6UWkGzl7uX68BdsYC3eoyW0ytSS
CoC8uyVJZv+zRiEvuYMiGVlpTEs+Dl9mjDbdNCdSQAJ/PzQ2mzpLLGkfc78FqfRq
6lXipW3zlZ7haIyK6gyPbqLqO99CX64Hdjn5vgO9Md54LWibEqdE8CRU3gm5akWW
/dBUB/dLF3RN/CB/lzhYHN4wgvl7JG8Jjmd/3KvI+ilu//E4ZAw4cMEo/b1nhuss
pWsSziQ0yCfK53ImpSAvSJnBEV+C0DGDC2hg0NCqCblTqh1Cb3kIRT6XCV8045uu
MaDo9PjdccIwBUE+hE3jrLDSA9ohxxirfLjnxuabDxshRoMf5en9wbpVgQBB9Yes
zEycEuWcadx95r8Ao7GjQt1tS+GpPx79XP+Cs5sEj+F8XudiLF1C5zKMCE4xmCEs
hCyMOftzxzRfgCUeNhHmSJAtk1Jado2sMtIrudDj+cdPG6TNNe/FHREzEbpHuTRD
mrbZjVm9bL4JWhm5EqbnccAFvb0eu315euVwaqfLuvsi0faJyPpgwr/yafbmiUm9
D4k1VkGP3cMT3kcYdBbtCYFIL/k0LK5ehjUyP6msI2UUb9qG8Pb6JFI6h4DUvrhW
WssEyZub3G+4rkxwB+Q+gkw3+3Ka53XApyOp5f6VWKEWcXI48wO7EEZgvDB2J5R/
fGkR+cD6/SA/BtIQLlmiY3BUigU95dm7kit1Wi9aQ7lm1+1J1WO0DXq0iGQqqyhs
yJm6TXRk7yQZWAkrGrlnjAYRX0f1+l1wvhb4AALWACBQbRAq3Ozsq7aADY/DaE8n
oqag6ggiT67y1JMXWJL4M0lA+oYCsG8pRemqcG/VEG2VPP2NqTQH+BIQxAbMpFqJ
w47CuSSWRXHdQtR/p8TjrwtwE7DPWGI4WjFTdt698zyX4xIHpG8chCI+fHVqV1su
pc6MFEPMGnB9qjBH33ZgZ63Z3XbCfc0L8kdHzBOQkQc04300LfBjGlB4vydSNuZb
EUYonlD0OkmO5iH2pM6W/v+mXDTENtD1WqssiEzViuUS/QJEtwhWNRThZ3j6bpKG
PeZcmTNSVxh7VvvjeKuhFrw3VpeDeBm4wRirem3LGszmwuu6yWLxjpv0L1jbLLbW
i4LaDA9pLNfNeZbMb/V12ZiEkxPzPKYbDDB1AUwuUmmnlzE+TQYWKRwfO1bm888q
YcBggWKa3mkXZ4BEIGqC1p8IKkY8NWNFO/vnb/geH2/QxAiySin0vncGS/gqfRZG
03sujWEtMHKnL9VdxUK44GAfPgm5gX/8voOGGOLhpUvWGss7XCT7hkgDwxwfzPO1
giqLkmu6AA6zg9TRG6InBo+kDm++KxoA/EjLp8/5eO0++w3QRD3qPhf4YboK38DY
Ot4qt4MhupRzL86TcHiqRECLXxk5q/GpQM8sc8o8H+Jcdm8Uvq8hguKBRW3gji+r
JXl0P5QA1ZCFlfso60wVdN75Vcrm7JuxIgxrklx5UlkLKTJ4UYIbdJpId4jTpUQ2
FHMZuwoz9Wwzu7nD1JNdsaf0Dos65oTFqWw/5BzJdgGOnqbmGAkLmzQ0Vv4sNqUk
4zFyfacNZQzP79LHKiriWC5DYaW895FKQuhAlbwMYcTHYCrj+wOXqPR8pN3WErE+
ShLAiYn5ag2hzv9nLNeYlk44Ax9tmMCnh+MET1O8AThJKx7uI39KyRaHToej7LUW
9d8KLc9xX/jkqMtzdBLK0T07Rr2FO9/FSEMz1e6mSimQoYnz3nX+oKTuDJ+UT1sc
FKyifWTVXIyo2agKDvgAioDTVs1kJ9eeiHZyw3QaszuJaSVZO0vaylsnrcmE/QuN
bo6RieY0oHf4FJJFojrzxQ0ou6HKpcnMcJIAkJvQ0zNqAcKKo4zyC+45dnD13hAf
MXBvjA+aaoYWZb9iJDLzIBvRwZOHoSCbtWfFiMqx9rSx3VUrO6r8tbWF3mBh72c/
HQAMYNC/OY9VbukuBN812Z6zDshO5hpFE9cM6tvNDnpO0Z3inlEA+pdoXTSGF29i
WNzpB3lCnOtdB/YganlPUux0XgXXydVFR9XgyqGWIFGfhKbydpT5vXI5JyNy8fw2
hBDp7bKsLmyyRvorlOvYPN9uKX9V2PeOrwN7SxoMQvPO8g26vwX0eG2ifjuLLZu4
Mg4zUgVu6GGrNoEmYDh0gzR6iEQFkrDwaM1sAwW9Ih1Kxf2wwJJBSoSqgypEsKP5
PkW8clheQADL+H8xI1PWf7lm5lunab5iKui3ePd4NgjauAsrqQM5zeat59ZNyjjI
TajNfPp2WyfeASY6T/djLFFeRXbvBmBAkxmKkTNcqGSsLZpqf9D3LfNPNHwYkdIw
GKjKUvT0CU4iFZCukrtgLOpkqjchQI/SHngIspwscnnxcOSOf3YN6HbyQqGlOXY9
5NQgseglaJLXH7Jixsd3Di0MMkuMOIqxydW2Xb2xj6N9Ov+IXwcboapB4nWI0+x6
3u6gEvHvZcIVCztI2MhPSykA0OgvJGoa1O7CIHSnUv5A86QtqPaV5FmfdnwMQvKe
v+6OSGq2N6MMgXEVuK/9U5gFB/zzeoGg9vQcsVk6nkc4Yvazp4bkJQxg5uhJpo9t
/92W6hi7DQnZz4LboOOHaTbb5vnPDQey0lLm2sdoNc52og9vZEHbFyn4hiw+66ri
drPfedrsW6KZP2zIX1rSxyZN4BlOP5ugkGEgfp+ErgUH6x24cE6NEaEEWmGzwyvf
7JZxMKRs77hTFzYspyxcFwp4Vz/8KstoDqmt9rN8CPI0sFukXCWiAIbObm9vD8nW
5gHcxYE1PuhsTR1qMITbtOdo+WUvdc8v+4qOTxz2fA6zmBnuqKZP85ZAIkQYp9jk
QJNi6lRAFpMISn+TW9t1LiB7uitivLwhjGwId4OSyqOUcKvrbmQ0SZ7CNgp9Pa6N
i+G8yTUOfIdlOpM220/6iyiIjGsjkypp+59hCGV5OiSQndnNa8/SVAeKR4B65N/y
keJV+RNSSxw48onVnD8sUs4K7PE+kOWNhCIW6kleduXIit8YIU2ZkIZB2tm7487w
ZXkRSxgNKCCQLxPbv6DAQ+hWIWndk7KzpM2wn1nYbV4xGob4DdhCqhD9Sn3dTNV8
rCaJpyRQ0lbk1oP/5rUCF2onCPM/1VRr/SU9TSAfHgY7OciBbqxQOMm+AS192os1
I0TAZvc5RRm0YGhF8OquNS32SLWXq0D9/2EtfWesYTr/RnzximG+u9u2RnyvImsV
KJaSKUAVhPpPej1QXX4paOe2/ouU3/21jr0bAFdFHvVRGKjLoow+ZiGXfhJDqdFc
8z1z2+yI2BMMbgECqmFCY5y3J4CsZHeYziWvThPDgqnT2KGw5ov9zfQsngllnmsz
+Rje53kxD1eXy+RXbrYv13HIAxx0IDbsiVZx2jaUp7rKyM5bvd3uHGeVMtlGnURR
JglBzQV2udjiwxKuW8n4LzFxi6rNj1epfV5j/y0sZLVfBSadBlpcWLHuYIcoesBl
0UUQyBc5FrmNUryMirhEQ5QRt/HTen/TZsNFAqJ1s9GMgTliw6Y4Xdv33S4iUobK
5jwvTHvcCuR/D9RNdopoA5J4fPEL0/FMmo9WCQyeF4iHBXLg8oq3M9DzDNEqfoMo
2//pSxmCGy5FOYq/NltuRleQ6k9fd7E6+a1GPznAA4devzZGcsxsfqRDNSqCG/qk
1TO7xPp+XBRaoQtAhGhzRurEtCj7FLwpEO72+WAUp/SzNPq7srHLl+bN1yBG4CRY
lZoJoq1YlCoM/C362isLQMV40lxpG+OlnzbwkPp4zBWBk9QC5sxdMWMcAf5XJWyt
3DaCi+ouZtuVJWd15yFnGTBfUPiw/7c/pFHtw5kIpElf4wFAZ0U6j7piTHgmei8a
fQijhH1a29h5WmyPzTfxKibORche61qQOBgme3vUnMQAcNVXs58Ur47gHHCpyR9O
yPpkX8HPHCSHgB3B3Bk9pll2a2FXYx3wFBcn9wG6VkM6WVDiqd+DJiJEHEnwhvgL
i/rJxd4wH+6aPcbstJJSgYYMKqWltna3Zw3fp7U8/9cWuTbCKOeKCKKB6JnEI5Ho
0VVRxzQj8hiwQhp7HwszLRXgIN30BatQeQIBCDY95mPhsLnJ6bczfC0eJyybUbfF
7mlMlLN6IvZ3sqiszquBAoWVHe8JgLJLS40B/rQw2g56hlS/15SDMzCLIX1nuxVK
OfxxPodAV3p+Q0kB1AMF9we7eZvNrFWNakUxF6+RWR/F/z3gBTpS45X7cVwSN6/3
dCRLI45l0UNcBa+g3Np+mxzlNrDr2e6Zr8mUzI4eFHTCmo4r33YUzad3vWNWc1HJ
yDWHmEjjIbN1OOCfdv9wkJaoutIGZXSpbX6TBbUbd8fyF3fyvPckZseP9ItX/3mT
4rHDbqrZm3znVC7ybTO4Sna2lgcyCKuQVvJ7c+bTnMUG5do0enKrALQyB3O4/EVJ
IGznh29mKVGeiVsi3701GcuahBFgT+gDN13FuygaFQ5iSP77+ekYeBR7HEUX3sTt
bHZcs0MqDDzuXpQ5IDQz+xlQtallKGYg2QqTpPB+IfaF0U1xj+jxLbwN1eIJXAJ4
fFvwiyprRUmjOO/tcgEPI+dkljB0hTG3lfP//pDRtG9olDTK80tyfGeDSxR4fF/W
MQrf2v4msXtybftjXFzqScX+27GmSV8JI8mKvwaXvmOv06ZuF7FLFiPwFizvDLYH
f3Ee2fo/iY0m7R8j9DmQHFLi/uwJDWccdvqBJftZ5jSRkaadpqXfwfn89IV0ePy5
WMAteks6idt91O+xBh9OJJg63K1vR4pQQhndYaB6n1zidGIPoCQSKzh0Oyf2nA44
7q+5ToKRCiNX7tUKNsvxlfdiAjcXHBEdyX4BEAoBgglq71zJDmIRJ0By+UmRRhjh
8DxETs7wXCF8YPk8Gij015GeSpE7OHdWHrExGsicWVhL5/kMNVAvGqOX0jbf1sMd
iDTiO+GXaA3bRXltiMtkAiOCv22DBri977rCiK2TPg2ZuJ7uGy13pYywmdZXH1xi
sVltJ8U2kTW1Awsp/IiKicQwHPgek67KLTXFLMWAZAGMA9znydP8g255QywCOAtf
DGIpRGu/UFB/9fWssLrP+mPuV7Cz36reEdQIH/94p26ew8nY0SYkUp+Rs/0XsAL8
xpkt2SCc7BpEfenbS3O5nsDbo86OfEpYA6o5dIVHRi2Piq3WsKGaih39rYo8BL9x
y0/n08gbAwccUpCNhLmeMHUv90HdV6Bei5eiSHYITG7GlxTBQSK/hwHCcKiDMPEx
ak2W2Vtg2VwBUbjbrGW+g9O2tp291HOO9/EfX0PNYyFOBHYEnERxhNvBL7UC9GmO
XG2HLSRRPwGkWlgF5rH/7mx9u63fTC0VCtK0ziXDMy/2WvwoFg/lomeqxza35BcV
2x5/yRdvBEj8h6SE0qQ3SQ1kX+hIRopx6hprJWQKfvWjOpkk3lUvS5gQxcgNl+5k
691ffy48DYO3XvaeJyZYKJheN5rx4Lil2WO2CDQkms4HdtT+3SgkYYDrktXP7hzB
P5QoHUZ5G2hHGmhAGbLFm3omt8EQf94ILdsd4KADE0rMsxJREnjzanSr9aPPeIc6
HQKrnUr/QRq90qhw3M2tObwHIq0Bz4aie+VEj/3RLb0YeHyojmf7jR4fvHTTwuuj
5GjLfmnUkD2u1LSYFuodkY65Iv+oiXomtW/XI+Ihd3odad04h8+fu3snVfzIG09P
5euiim2nAmk8wgxei0n40jpnggnqW30GL/FWmbFlrWFiXhrt4FOpOm6GqHKqOq67
Vgq0e+kKUWb9Y9QbG3+XLVRRTpuvCbwk60V0d7te9tLNGt/5/phErw80Txhr+dlr
OyVMDhI5ttq3b1uFoKcx74J/z2Tw7tgppPmGNvLyzGpPNLX3DIqT32kptA5euubr
mmWKTaj2nH2R1QnLWuODr4PXfjExNE3v6H2wwBxnkSr2NzYRvOB3qPLVW59y2+qM
d5rA4B8G7ozsyDbqHPmfYA9ZR5F7FXSPWdAXNoFjHuHOyiHEBL+sHbF2fg65PYCo
3gil6XP2d87lRpIMR+0d0/xLszpjb493fZ4T36EfPbF3XC+LRfpprNbohR53Jq5F
WG97hYZz9VD6/Pm7bgzevOh2072wl9FQDBD8u3gcNMyYIbHyjY7S9tji+kAGTMOr
IwjndmeKg53RQQosX3K/5pWE8LiA/RAw5vGVjAJtquK+SqCjbD0LTlprucH27Mu1
9Kv5bKoDJUKBVilO/BvRTyLuAquM7gjTrqNApatI8SDAMH00B/1wVd6fwuTDrMR/
CoBXAztpYGqXR2Rr5cKo6Awl7lI5jAPAMFo7tviSgBQtBOlNbbOMjIyEl5tVgHgI
vnoRJbAmnp/9u+mfT3qvDvagdsGwDayTgLVEBRjDmP6shGyc7KGWjVGg7sWfHzA9
Gztm1BYVVJGYwkz6iVulna98rY9bcxSXZL6SWyfopKmu3+7mKjkEuy7XfV1ete0N
MQEWj3PcAoE9t+ngZKUw0/UzeB4hPCmTx9d6yD6QHTDdxhpCmHNtAGh5HsMOJghx
lFck0pClSeRPPuyApNvFdWCPkyLk6K6/CjYgYljymz74BksKi6j4yGYmSwZuC607
KIpALafghV09sQSYOSXW9gVl2jlWlsaJnsxKKYE4Lb9K/EGxQNDgiW5Lg60XA8qS
1qa695HP51i8z33FvsglSdhRRWfS8prOOEsIjz4GoZ/b7VaXAWqCR3S334NfQXy3
FqsezOp0k5y9rCDDXRkA6F1mms7b5RFinKX37wAEt9Hmf/BP7Fw+QZ2Urf+ERHQ3
dKzku2cAE+7jp4x6IC9+Gy8+ziUE3srycffcCZx4igdLqZ+uZFnwkbddZOlMAcM2
+ZcQvxWoSuF6dyhB0Us81LdLXK0ypTd28fJ/TZyEfpgeLOjjnXEHawj1/G933tZT
e5fx1kcVZKfxJaxLLlvGXUrMDL4UBYO9ZT+QYoQ/Gf5LJQwCir3lg0SVJDQQ80s5
80ARB//ODx2DMw9VXEN+xBWuo3qG5Sg0+4Xu9QppcKpUM7yol+OOIUNS86AvHq3Z
hB2yH/3qMQoiSlf8iaU12kkViZ0BqDOiZVol67VhN1a4Ez45ZvoZM9t9FYhVtO6D
FcKBgFbjZgrcKbaVqXS5YxsAVrk9JnY2GKsXqKqw495CxSvDOgZUiP3TyrxncXzN
r87dI59s2STn2Hr9kCE7+iTLzQgNbz1WNcv1WmEPgdrdDQDoDtd6e9Cnamceyv1d
mqXmWWu6WCJKaz7Up+E6wLISJ2jjgcMzqjQd0Cg7wYVRJKYHMDEJssrtuxI+1TI6
COtFR3psA/p06beLAWkP/ZfF7k4gjFc/Bez5aW0VSspoRkGTKQxb5MjNvVdAi8Wn
cbNSX0FGcX89VTSosvooVlmtnAxGCPzAmJvGXkMVlSZj5Ir+1VLHU0L4cwengHNQ
HZnH4D0rsH8wQB/Ijx4Eq1BZV3ZSAkMI1BVML4XkScFyDl9FiLLKRuaVN//hitgX
/awbViQadOWRDMgN6x8x+mt4hR+CXHGAVGkQKEIPwZF3Sulfh+mggEq/BDayumYC
W0h+6KJoLDp6kNXMFalQX9HER5OOuWVojk9oplxe4/F8Gw5K5Bm7QwQqvWY1km3T
WT/x4O6Gtue1eINFuWLe0ZX6wp85Rsegs0Ls8akFHUaudMeCiaIawcipbuOpITLI
XUJUDXN6SF0VrVc0GNumPm46FpsYiE/ZwMk+E6NkUUjx3IMEyM4vPf0xHlKyUCFZ
l/fpqjwEkc7BsSP1Ry2HhlPwXdh3z5RMjTCq2IVIADkPZIM1CypUATmsnXoYSP7y
YLcBcvLzGk3aETErc+HSdE/jMGyZ7mJmjt9SV3g6MjNarjInaRjkHC4+V//qJQhh
XjNpv3A89937mWTHDDVJEgVwvn8tSxrzA8TF+egz2uOo/MF0iXJoH8odWsmb/xon
mXL75tSJib1wKpg7d8lyYzlXFb07xkOJMvp9XzEON/HPSdPNcTyIlUeGs/tqHBqN
SMrg2IXl0KSlHpByRn/S0YflqWfLVFjW1N5YLQBRi4yu6KXN9vyP8AZM93wYM4q6
wsHHInQRyOYaucVIr3DMSc6x2XICALadezKMRxU3gW4hKgYVN7ZTQvWigzsDvoVn
dva2dhtKSerOAqltaPG4lkiUSOTf0GZeKoF0LMd353MEUQl4Faiq+Hifs7y9hlj7
8ASySmyg+eIwjnvo9d4qHQMcDVEPX6H+VL2ubhagtcJA8EM42rbKHvocqaiGzFY9
81/o2mQvX7c5dJd/osi3Uo+drVmOTZyzbubg+C4Fq2MApA61P5ME7jRrRJXifOF0
wqqKF2Dpft1MXDO9nrb0rPlyBxiPaSWFiprJebzUdgIktqt+iY2g/qeloc1TNy8P
s2NT/K5g+Gn8yNz1Y91pHf936DGT9vizh7eNLaQ7j94hO+XmZL7pPhz3FfUY4odu
PKYuLS8H6kkJph9/+KGdozTt2TsBoFUH6ebywpUyDwLSdJK0xynwhKmkJWF5AdKt
0AAanajmV44BT+h8OKQK6BKEL1obG+oBo/wp7PHYF7nwi1RoZ6svzHWyWf1ZbjLt
p9QyAFIAq+Pr4LnYqXFYDaS0/q7w95BCE0zHEO2okTnnUkeb+zKaqGILLO+1F3u1
WrT+vcIhTSd6StmpWpVsyUvHUU1eh6sJpe9PGpjg+YX56kwigawLPe2sOJycSRqs
7Boy4VGAqoV8eJRpHSrTpd7yRv8nDuI66m6Ms6J9mDwyJpdHvYs6b8uCExS44m11
MDg5zbW3lc2oNGvha2B85FBq0/iDwTCnuHTT1ObiteVA7g43aszlsibeLl9l3+fA
mCPwJ1JQU5ezObrm8tgo0TueCub+B6tPJOXDfYrNY4LfliZNoGciRbzN2NGK2yxW
EeR1P0S7NWnA/jTmuTETR4ARk5Cj3xdctZ3/SWGvRawAr8yeXM3F6eu6vZ2XtaQo
uTdmsECOHQS4d84oAPoXF55aW8EljOZGf0zGOnyDAQfjNbUTq7smQPjg4Lqbba3l
GrovtSPCyhIPyd72cJuAMC8CWFwHrHHuKXyEQXmbwc3Q2ST97hrygCapuMU9As0J
4K9RcSZ5Q4mHDSGEus94YEBp+L7LgkWzNWBaNjPgKP7j9a5R6pqqnjwzwDxUQXG8
vrO86s/wkMN2ydMDUqNp2msNBpvfA5gxi58hvFHaghJHOdWn/QzXGrdXxHKWAYUk
r/FOPUeQpk1m3lCUqcLTVI9o1LZdIrmkNYre/rADWlW2Q+/xyuLjH79n9yldGHLW
sDm3qwqGBPvWCDxqtiVa9t7HGWOBcHS+5t5NvG6y0XyBEG7ykEMTQLvxB9qLljwL
4SIJ/BHQqFqEKr00nYcNX0OEO1xY9YCJjN/rHXHUejoPDhZkvA5cVcWj5HV7NadC
mTtlMgrfmz4aI0l4YhqoFK0xygcEMHQw1d5nG08iwjDPSjPcfbsaeG+xcE2utobe
zmN9zPqJkyqPfHqpSwxfRXNFd8tEYS7U/4HtZam9QQdHahB577RqIgRgtFAE8/3Y
IuRDH5ct4tVfqESW8K6uI4btRr9zY15bIET8ONmYdEDqadFbWF29TL+cbp1KBV7Z
1ydFbSTFkzZOB1ebPrqvBzDsjxPNFYcqbRJL2WlFemus5UbhyPZ7e35LcsqaBacy
1xY0CqqnuLo1HQ2c+AzU/RtlxlDitpBUgr6PvpYb6Sylm0y6VOqNPLlg/qIMbXDB
YlZFhG5vU3bEjyulFU/iD4MRn0YlGCGD93nNlc8AzB6GPyz9OHDwiR8O1iUz/RRs
aEjKKhsSZ/xsXb3vWS4pEg6oHhQPeaubJc0k7NLp8dYvLnEzyIS/TmdY7EdcN+18
prPHr166tov4tBAIFIJODACprwqxQy/XQMkEBpd3lNHfFULODs9xGxJY9+Er/mqg
vOexlJ4oB0fGz2dSGDEyjgqyQZZnMudc78Bj9S+iIQrr9a2ATHo68SgLHXy0MFUg
fa9En1FwIW6z6kH7A2EVTt6cpJ8T3V0hZ7Hb/NrGi5/A3aur0R32E1NFWMf2LZyf
KhqkPe7IRFmQr0PChGJ1OtVbrmyb5+VgCPnTXQVaGpLRlf45Fq7maBl2rXj3+/oH
9SCHPD7WNBb/w5GSOIP9L/BtDFQfQdVLqM3tpdKZJ7bqfntywDcSoCzM+hD8NX39
dvuuV+puNNOJBNt+HFDfmL0uFehqIoBVxAwfPAx6MW27xuIrLsGdobZUL/qenvC1
E1XUL9Sl1SrFUhrJVvACLA3TU7MngO90+qcvgfpAI+z+xZd7mjLGYeVqa/qhsoyA
f9e8FQSQ+lvnObrwOBvfO7j92ieO5l4Dw9sm43dHqeMbzgxxg8g4mvVLZeB7o7ej
9gkLu21y7D24woDpY07cU/Vxhe6JNaAou26uOwck3PWEL18ziKYlvpQfZEEuhbim
hctDovzoQrI/f4Tbx26mrHkhmJPsUXKCDPF3i1m3bUTUDllwL1JYh0O+EI8trQ27
GD8mGDdJmNXR2X2cBfEkohraztXGZin4ZJcxJ5CFnu0d++MK0p/zy+lp7ZLA1eaZ
L31US223XUyDmxXpGkq5LQTWhubW2N8Bzq4cWoxESJrKcLg+okA48LUsIYgh+SzT
IxKbKGyDPN0Z1qEheGXod8IiL6u1skk3j8bngCwQ7+/wzYtOzayGN8fszS50IdBc
2sQauM7NwfoBAqFkvzXOvuAu0TykygdzEcoJPmBWNvc3srrRSss7jFEThr0Svb0e
+YaI9LboJDlRRaHIRKuYf9Fr1Wes5DnTU9Eq32U+wjyHV/zZKr4MdG8hy099ESSu
tFehDa5W3Qk3Eu28MbYRSLo2YE+k1Yj0fDjbcot8dNqNqh4tR8SyZQR+ZxOSus4b
RKRvyrOStoAd17uisIxiyk/riif2Jp5uigI0KMg1VJ7WUONM88kTtjf5ZhL1PhiY
WPybWbWGBDfNDS1y+NVnN35d9K/g9l2JGJIu0m6I3njGB+az2g8YYagClX3hbhTF
8MPK5HjbpQmXR6kKVliA8/82kkPfePRAE5ZT16TRGgsFb5lAKzh7Z7AFcnYiWxV4
+hSBSBdjWdP4ivzYkwYqz4Uh+vRAmagEt71PlzXssix+i1sgIuXl6zkn7F8m5Asv
qhxFx0nXEKGjiHdf/SJbaoD7cYEVLQaRXUz1v4Aq+EILaarPDDKKlub0dQpkkGXi
rbV/WUegPNXpwz/neRi36oW+WjjY71OuQrgvL3BXpRyoPJ88EgvuWGTNS8T0AGtQ
d/pmwCDpjNUNuaujK/RMI9PuzXnm6pk1XgfAZ8qCrJiLVyAE2HVW+lZghxjY4kqY
KzIqKU39GNrKqot6cKWl74XgOzc9SODAWFqHIjIv6I3OGiydKIlYzMOFn4uKaznb
7BnEUT7p7uj44O4Dwysj2DYbMF51Fl6g4JMlpts4fkAV9gfJ8iW8CNu7LevDecwM
qH/0zi5AAQsjXBIeJijd9rNB9W/rg5sRy91osTJK+1rGD8SG706VehtRxXWx2yDc
7uKjtwZ4fDRXRB9xCJHN/sXo7DcOjZewAitFjmEEXiKvosmz2cCcSCOv+bcsmHhj
5fvZ6wDsh5J73KdrmNkQIVx1NAGGpPNwJtEDElcQ7pyb/k8u9Ly3MKUWWnV/+MDp
qdw/PE+W3opBBTxhAXsXzU2V0MBF8w07TRjJWpQ6cgyI6PSekTY2XQDHO1enQxQ9
FPeqrCjROXWtqvs7uMfHoQ7bfBXPVOyrPNU9b8QhFvrJgZB3dF7HnP+OIL5IGeHJ
5fINWtZdtjlJuGvySCqUbtqqMpdgH0hR01I4lAuN+ALoqnjG7HwkLsTebgvj3UJg
SExQHMyVbH2VnuTfucrifTd3qo6ixDwXNYI58fA06xZ2VBzE05sVY8ZI0KLqwtC0
/hTBTLw+75pPj4S6gZdRc4w+eJ76p9cuqjzwRXGc3T7ZdpQ9uwlpNh0YXpjGErLf
H5VglRD2y9NsYvlbkQO+NssS+oLjmUzb6yAIH4EpygLf+yWYC+b20Kej6AMcoSCz
ReZpHPi1VdTSQ9l/IJ0y0hVVEGEGEN0kuqC7HxFjXDnnnEWW8zyrKLu9F1gkyAqG
rAC3s6OW3CnP3IqZlSywLxPLPIf6+mZCalLmq3KZHx/NNXin2Js2ReKpc6X2sXIR
257rTlvWACnMXgPWZga7cvGelKBqJQlell9Xm4QMLc5rqiczRq+MbwRgGZF/IDN9
Rvg77/NfHsmSFocFhskNpCe1QVveRxI2ABmMkplEuUkD0rrsxTV1Gu+RVebu9Gv3
TA5157d7W1RFV56TBXI9Al8qmfXrxYL6XdtKjHsUb215SUKP15MXJR7pSaQy3nBK
ouyPs1etbKQkNHcDP9l7eoMMX2e7s9Yi/aXIaFOiZbqppYD0gqZskxMkVsXPleTG
99krOSKlOCTtNAz0kZBaPHP9tz7MJDKjPjY5MFWTy/aeJ3iO4w6IBs4eLy6xf6Zw
qagMTVhRBRXV2W9Hx+0H4DucLGBcW5Piq7D1NEAdZna7ng4H4TQPqJYMBsrJ4ANI
sY8G0cUaIgTwouPcWR5cRwegTUcXSwf9Q8R5LQk9B9hHq+dShV70ncz1Lzx9Oqps
k+v9Jmw8W/7d61+KL/Lk5Ur6XUlKFRc2/J8Y2COC4SvigAkv0yy67IqjpPAtwfDf
1ezxjkF4OOfimXkky1/CZ6GxpGegc5Y/P6VIq4MwqqhbIY1LdgY7Nw8scJj/XGck
9w5fLMywttbARQv4OskouL9aMWZHlBDccNBglkuZLGIkm9CjrTRMH+Lj6AcKU+qE
j+2vIIn5Fm8aXloe5AIV4uiTKHDc7xo3xJcFg3vIylCjqsIK8rsDlB+iBeHJp7aY
61HgZvHDv7ZSOco7q1rIRoIEFM1t9nlsZvFIyqyIRS90yOlYOwmArEz3REKrKDOf
bP4mrCKLYHFuv4tFlYSffJl1sxQu+PXmdhSsN34W1503y+vp3GS4Z4pYEWQJNhIk
SLK1lwQ8IQJUdSBoKnQ6ZX4LAT3IoYPh4uRSRmylr2dFQfoKfUC+XY03wXzu/YxG
H/LNYiRCFLedFkPp3piyS9uGPKT4VDz+TQlREXjeT4HAcLLROXvdQXc8IgTxzmNS
zRqRpNvHDZ+OmbQ5/tK6vC9VE8W4E/6wuK++463u0kn7Mzhc8iBmCpQphavUw74S
HTrJNgXHudzMQ0w9eCKuqm+V4Oh+j1ucqgZqJbyptCVO7GJ8xvKVn6QENGTPijHV
EtJrjzJzVdlPglw5Oa7fjYeZ54mmnqSsuS9ih0aA0EY9nenZ92kxF/nVlli72j+a
zk3ZuZpXBz1aRErT4VwROCgVbzeXi3L6xGUq+WsD8bCVHMFfAlhoajFrWTVp8BMb
G9ZrxZW0cl69JTeOf6Dd3ymFt2gUWa65iPXjVmrPQFU5uYSreuabYaCZV0pXKRx3
fWqiNFSJqOAV6vHkr82rn6MBG/HXj7lCtL345UNEIxNy3mLDSqHwCV40PQw7gF0Q
ITKv61BYSpju+BJjFLpme9SNVC+d1g72buj8pohcMB1bXBo2zKepNi6ydc+ZrhuC
REWnPYaTSWtv1qglpcMeJBsqfs8QuLX1nYPM26hcmUvdPsv6+8CcOD9hNpHtSpq8
M5ZtLIus9mnOL+QP4o0cPW/HTgg+pTMqw2qGLzpan/sDOnt4yiQJk+8v84pRKZsG
uiYpf7vbr+/0XwCm0OFRhc4JJoE8hLpLTsCF2EOdJhVx/0/tcwBZebZB5tB5aAgm
L7ciGLIdc6nVNranVinFSd8TqBTVf3pC5WjP9j1a5bM25Oe2kiCCfOOQa0ppN+XO
O+S6tQORrfZZeDhIvdn1wdNyQFzqS1AkufLUZ1GPOXd6bN2vkCi8v2LVkdgIly+4
Cu3LhD4+mjvkfZyiWF09vvALgFlFepMX0WpdNHGGBiHyl7btGgBnJvmFeOgkMTqR
OYFIcGl+4RncuAr6KS2B/EHAW+3/3qdp/cSPuD1knSS5l6FCVBTUGhNCsKVFftoB
HF81fjKCvz9yN+XGduGfQNx+ygAdBS5+eDbzjQSE/+3FbMvdlBhQ8qMuKM0IARQm
OwB0SoV3IG23YbWxcB2dbklKtpE/uHse95sWiUvXB3jEOr7mVK+/Ws2KUD/M2LuW
RKV2uZTJ0UiI1NBkN3EwJrrds7X3TqOiI+G5S1SHe8Ec2smvTqTF63A4OnwNpwqj
Du3vfJrDrdEeCcjbGbJCrTKBlI2c11nrE5WZgLcAL+OpR9F/wK/DOZsFnFPZcIeK
HI2sZ+hS8EEFXU6Am6Sbu33l79YmckIafOTDtkXUw6gA31rcFN2OVW86i01f5l1D
XNYspV+NpUG/3PQ6TVctT3cqSEaLewG6kZHLmXO4QbPY/wod7rXyUG8hy2JWMJgm
gOIweKCcNv5IlNPVK1VQ62kW+55zuucwwukToWUJHUG0y6AHvnJJokvT9wBg2dh7
9ZZa8f7j5VTyeTSpPnn/C6vMe/MdXctG8H9wUuXTpOSrzIaH0DlWlftdKozwJXMd
R2sbFpLPefFHFscl5DFjX8Z4H6uOC942LVPAqZrmSZN3HJES/r3/YbP6rpT5/u2v
7qkpToRZxh7n0Nj5qE66rz5y7cfBsWcc85+Eh9ok+80MB6lqd26Pp3hItbYrEHlv
mj3VN6VD6wHizHLOg+84jqfBUaUIZTo6CcBbvkwnnCuH4mD0LwwB36MENCs5dpsF
e0UH5UyHbtJF3ZtZ9+GaJlVKl9pQRfIPKy8kqdphIHTtAFfUXD8PyXTL7Wp6km3g
TffPwOySTcUENyVC2dkUikbwrRtpSM/uuiMDN+8Ehe3k4Gd6xVtoimw4bpDTPaPr
LuOu/87VsjUEpLI12Ll/7EA8PM/ByO1C25qTe3aMfZPmPHPRQLxikTkprYwp0hl7
mEfCLU0l8SsuaPT6jr7VGo39cCaB2iyVtxs5Zb4ltrmnxthqRUXwRZlAv6RXeYa5
Jsa0jYRgz3xF9BEZO78FY6EGAGlU+joLuHyqyXWzimS9sU21yANbqJ7Ixs64nz4Q
L68QrywWJGcJ33ejNk0DndIzWlEq6y3NECBhBTusBz8aAngnPebysByjjGvS9ExU
DMqdBmkGZZOVpmsPqrG1QJItSvdETx2XUuobC0PVjqWpLFPmK9ThHbOY5CVL0Bx4
2G+q8vgffV4Jh+40NhxYCr8HVjjsXah6oEliiGnWmJPia6h0Fo/3u+kYr/49NsSk
RpPB5Qq5c7h7nEHArlUeXJVjp4vx/YWudQ7iIj8ETSf9zUnY/avVhVWE3ZqxywmB
L0n0+AliKZYDY01HXUvRuUbjxqJ8Fa+tY6CiScNFIQFc0A9uBGMDvcM+BhBkcYBs
ByFNlG/KLcI7A2iwV/kU/m7IKLPiHPoF4/kOf3COLvPc3whWWvgYbs1f3HwWrlqP
RRn+fHZN9WItAeBcaT/G+56R3R1M5iHYXU5Ig6COk9rITLvIFU5LyN4athwufU8u
H3ATTILkC6MLxJ1XQUgHRm8aEtQAono2wJoUHACHB+ZaTUJ1x7p4mOH+w2JhoYqw
WdB1NqlA4h5OQ1peFRwBYVIqdTLS1zRKoqbtO80CFUUwR1vkF8TeJeipjQzsHW4K
nIxQTG1voJ7C3H+jRvwXPFmDaHLYAzKEKCUoTRawGyIQ+GCbabncIYYgVfkNqhwM
jiQo0dmOs3IVrOPF4C86sEl7NaTBCfA2osCZ6GJJ8A+AWqrYayBYUy+QL3S+Rudo
2P+6fbc2g44EV+DOWrk3ymgKIWtOhHVA6wVS+XWki1TkYpcv2OdavrX/Yig/5q8B
Bg4ea7xCVAGLn+8vAQbcXGYNQo6psujGOtpaHgod2SOpsq/3VXcjZZfvuJo9yVkj
dwRvSgjgWkOqUu5OlFeOo8L8TgTxMlkY58ZKuuvS3HVEDc192i2MVQAGdX2kijuw
4eTE9IYMnshbP1HLI32kdHR7gOSyQvFNfGblTVvGc/9fWlPkmCvDUF04oLjrHgXQ
/wpZ3hmCLeCCsvwWwoVS+lNqAmNnMyVugNNuRz9puqQj5gNdqN/wfZ8yos7DPJfP
zxv5Ec7EWkV+dniGi6vaKV9MoK7cqSKO2yaTuLsNG/u2wS7xWz+yiLnDWJQ7Ls1O
Atzy26Ia69njm6zhINCFZwWCJYGshO5kecVF0/7ExazCFVft2ZALvOKG8owrzqzl
ejpg80+zY9MQDROOF6Alj+q4GYhVaovxsUSKOGcEMLrjcySpKGNWqqLfFvrN6EKM
/yUj60x5q12ZsByePwyeh0KocXDyoIFwr4EB/QXmX1rZRbkQQ86abYdIjRhpEc0z
JEuIKHW3YcunRKI705Pepg67+FmZPm37uSI+ImCdyDvcnuleUfDHCgmgPA4PVRLz
Slist+XnkCMrlIC4o3Tg2MaHB0pkMTNxz4h4VloB+Q9Qlu/gHf9ZygmztX6Tb2lp
uMzvDTG72+D5/dqeh0pxyM+MhAPguHmRhrjHsWd3EpsyJSoCxdEu31+lFED+o0yt
7meJespPZsfjo2PCYsnyCkHbjHy71st+UTeIlV70gVmXpYVmohFWw3sbo6CA109w
KI6BuTIkwjnHxWlquLeFtaJblihOuu+7qE1+hR/7v7znXb4aUW6FKdK2OxKKLE8V
p7RevSRR+Q4LCJjbjpS/pafaGEQj0/k+CMfADlQUytlxom0w66svs9DYMqvQ/zMh
GtES9Edwka9H/oVIybjrjHH7RWLWM+xqjlmr4VHvCuowx3HoeSFXhA8zIjjUk2TA
+6qX7q66WVivgxiGcy7Ae6+upVxjTPan2Tcp2mvAQ5Vq8tBBwGrPubYbHr6V0gQI
6TPGwV08WjB8JRKUKaaHIYU3/fuNGUUAAxCyaS1VCtGVTahw988TxFzhVicLVvru
nrb+RyLbvKZy5Z/X0xQM/bEN7jqJAnaokU0tkZdVn9OEQ0x+mEP5a91XFhwEM4al
jyAvAAT2VeN3jA/j2/+VLtDiW9GWy0+DQbS/fUdjG+6cnDxopAwyfvPzqgGSYF7N
3iVJlSZ4mw0bAuvqAGZM4DmqRGgwdxznt7iNB7Kd9G5g3PRKF5Iu/MUWTp19LiNL
bwlQCS1aZVUwY1Wi6oYwu3s1ZiUtllIx54ad+J+drEMmSgmdDg8Wj9T8JTwRsUPG
QMhJ2YJpyEaQ66Wuug+JVgjVdKB6OuhJQJqHRy84cW8Ern9r8taEW811NR0dXEai
Kz7V5WQ8xASFm3E5B1uxbmh5CO8C26fqPD2+UKPlBJNS9oJlpjk7mzEmb17PaaBK
JubjFRz/qGfcAx93ML4z55AHJdFtXeXfm7oW798RISe9Z5xxe0EuJcWJKw4frv0T
BjKI4+tNZiFiouIWGSemZP4TX2PInN62GlY51Fp/HoyMU2GbWdCRSuIbeIwuZXvY
gQq1xkZ5/G56iTi/DWU/sBICKcx5LBlYkCnGbSLloQwQl+tIsRrfq8JP74TV9kr9
hS9V7pRWaPVnXGLBn9jIL0tzD+p1n17G9MZlITTVjxQf+F7KwkZiVrXcGn83t9H0
C14OQ/Gn6T986creinNgeViwvSLIZoVMS7TtHwbKDg2haOI4je+NKNhIc8Fp21WQ
55xPxGnGPjOFnHOtPdLlQMpX26/T1ZY3y73wU7CpXCJg1rCGT7zO4TiP173gfwv5
CjWDQeMDmW6pkSSYUrS0VUC03cIZ6pXLM/ARbag0xV8bj7BZHQkMh2GcIS3RxOPS
nxbCGVxYfMyVTHzD8nTQUmplBgNOGHveCHVihIv/COY+tDYsqs0i2emZeNF+bjIm
Ob3dserfY+iAG/2cZPS1mYg3sEZ1D3lzC0ZqXjfH5UfQPc+iaVQI7k2F9sCCv/ze
TdO82SlimhRer1vbbTQKo8nGuUIaw+X4YEPs0z/DJmez9T4KpUFTdsHLXox2ZD/J
DIN62LeAFF8Nd3r9lpVvU3eCJ+ER3zE1klsC5ccVUVB2KO1RHSoVVOumVWW8aeo4
y0Qev2IHSgsCJ2nkrQn9BA==
`protect end_protected