`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 13312 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
1z1b9VGiiW9Gp7THxpOgESt3+6sSIOLxsB+k7uXOpjZGLi6UvgQ+eWKGXdM0eoNV
TZYXrfHMjoX8bFluL1/55z1L0+6vAAJB9BwFavfo+4HLS2Sp99QupX12epbaHCBm
Jz99vTQA34xo3vm9PtSfHiINCrNhdbKCKFtYNGC6q/x0UTbua2hehrXO/IzY6fHK
YUnPWbXIrVJzp2NJFn/uGwHzLwAyHhj6eAj6WtBhkC27QVmcg37faSj4CvweQgCy
kloYnVDPlYfiSEg6wwG4rV/25awuyYnJjLiXLOOJRbhNdY+NmoCKJ8SgLj4I6Kvz
3NJzK6Ak21sbGh8s1XawHriDgSsJ0DGawSkvS/jvLJdFLBzlTeqM47Ktrh41rzHz
+QRRXWYyCP+Bwqg5JPtbZxDKhsHXNrEoDun29x1alAQoUKSwYirZ5QalUPE67Bje
/F1J3gkv1uO5916UXTWYYAL3s+cwWOsCpmni74kG6liaIgfDyXjFrImzwY27b5LH
Ya+Wl0aJHpm1BeSCpVYgJp7wvvDTc0QFCLNba/zJ+U3SfZbVhAWzxpZ67t7a8xHy
NPPdl0Y4uDAfmfENeIHBDObC6ii/1YCWP3rR5oaaBUHN35lkXaCkqo9bSYHmg1L8
iFI3O9xbXOQGqQWmjQ5Y563Uvx/nci1l/H6vxMHKGm9ayH8AEwQYUlTJmO0ZDEow
lcq+tj4ny/lfooyj+50xgHIxxxyMuZ0spv5QHyjXbHxp+0rvmnUs1j5ibfGNyV44
N1360BDMxplDX88h0jS6HNf6NhDeViGgKI66tEaxi1UpLnUE55A0yLp+Ta8CUKXb
dzV3zXvGEf4tM1kOf42xXTHHVqZekdOpGwyj0A6rYKOXlPOdpL8LBD7OImbNVyK4
K0p3Vgdpr0ArK/f3jo1suBa9g4aft8gT9IliZyPIpGIqrxZ5zoV5kSd0vyj6Hu/v
5fZi7mOaU1xcc07k3gXVEirzX2JeoFHRC4Oms2FD9mXLQrqZuexYjm88ooSjs8+d
9K7d/QUf2N8xLdIngoUy/JtzGIIgYM7s8u77sq5yQozqCXTze0x3FJ3fuBwMIjdY
vS2DjxT6TXllwuFHvWywktnOIpRHLVBPepwNXdNlkS5ni4AQF/EqCQ6BJGRVH9ow
LxqsEzZ36fUW4uzmhHCuH3Pr7UK3c49peOC1xBQMJKV/4siCJCa/qO841KdC2RPo
NLtOM8M0OMNvPFnwX1Czsh6tZRg4TRf/Tvwq6RB/pahK+qKAZyvoUUXZ/+uRzlys
GnnNucs8ewVkWpLmEwLvOG8ZX+cOfUxjL1kmTQqobDO+XbJ3aevRhC4g+0vRnGaE
aerurhXPJzTEk2QHDSjVhICorvK/1mpCQ1/iCvepgo1oGR1DU6oQdSdwXLNzlLxR
IAstqb6E5RSkUooyRvKcbjwDDOQgtBRR9JLEbWf0lZdwhiE6fq1LMjQFJ+roJj9R
E84D/GcrcYkuwbWkGRQ6UQQ/MHY9/IDFM3Zzi4AU6RZdHl9UwSBiVK1Ai8AX5ASz
oArFiratrEHxPxzhO5JwqH0yuVMv3NwmxqTO3EwxX3F4+0WKvQmmLtiv4gTiwZ12
EvcqRlm3/+oLslZo0O525E1oTMKZNzQWBmjlReOhUN8YtRz30TDa/fN2m5hZNcub
fivik2aPAz/8yHpLyLP8mFsVTGq7WLC4WH1wbQrhhoFFa0iU5zaMPCw9G6/ZzAVc
ckBbL++zCzDD1nFtHrVeq1kZ74HbaSE0JacVp/y1NvLYa6nkJRqCJRg2fA/EVZGW
IaEKPu/XCq7HQ5opBC2mnJjNczkNTuEDUW7tlsddJjpDmN4/Ib5IRUMe/0Is1oUU
6BPBQF8GgeKtZ3NLm+WIFpm+c+KU2ue0UIuHxkHMTC1rUWo+ozEvMcpfbQ9Nudot
Fr+BwOz/BoGfVo1lkJE4eY6aendKD75w+8AqwPQ04fkO9/h9kQmbihesJpHZYhje
J6zfgh/E7wBjCo0sUB/EsjypBVC6PTUqCIdughgy2NOItvjCa9e95R4m7Gxp/7T2
7fpwk71+tBaOhU8FlPeh5/ro62eXGajO1WECeos77hax7mWVOHnbF2TI+ji+ftwt
PXi4epJStN/kFCFwFbl2v9o7vqMD3lTNPNMpr5np3mlHpebCRJhpUU2DYcx1SJ9R
XFYfXJJKV9YdqpxTFWAauSF/fkS34xa6ASSgzkViV3pVQx4qv7HvZ55slO/zLz4X
12TpK0Wx7u7YCKRVqXe5ZXSC1LKqRX/yd/O8DhR/Re+3aKs2enIeeJPMoamrE/db
12z+Ss5zf23NjpA8o6a632o5CgeGetb59xAq0i86tmiY7MThSFHE41dqg7iEHl8o
+nt06e3izaMozxNwlo3/BgGiRSmfj0QMcObyv5jk3Aic/opRzLB3vjxP2h1Q0rlF
D//PYDDzlx38TPEFDskD1hYEK1TUjFiOCUDVaxFZJSCnaH7d5hvONh50xm3BdzkH
2k5tzuZs91JfZWYFeoVqPfEHe5xQKYwB2z2Lw49mus/ngewn/lGkRwdqYEwweUMH
5lkUg/vyvx995bALOgVILCPpBJ5qnN63wE7dHO85Lh7TIfAROZrBtFiwJPSOShRZ
qfOWiDBUkUrltkcQV17fPVIwh8nic7bzSZSv+1dvuEK9NZga9yeVcl5GWPlZTAHH
c1NZ/33EnhMMGHFoWsV7BZq/r7pyJAizGnIkkXmQLbKr3dsqFurbfOLVTADRoXDI
pfKG3OUIvXc47Uy8gnHPaQHUxCd+N7AneJ25FXuUQ+mMYcMVFRE7s4fLfwrh67UL
uLhK5VeROp7Ip9SWmcLJAQw/r0NMMDnV75UfcXxMDf/CsqjtxK3lU7S74DAEb6hc
fgQeudfvi3HF2X8u3/enJkYqTy7vWtU5Z9v/R5ODgY/zH0oYAcxRr1uKquOjgesX
ttI9M9WYEXGMwQxIJvf+QyGmg+/IcCAuuCYSGMYigXJM7svFmy3j1UXfrPXpwrnm
A6CPquQjNV6z7jhlEsS/e95EHjW0GAvihe4pFm4Gx6uu8//P7iGs/rhCA8OrU7av
lRSz94LbNeVYZw4CDfZMgmoSVyMycMFfaCcGRRuSms/umJXRGgbRA82XiceNwRa4
bhIr1Qs4aGy5c6ZhYd7km9vQu0K8Nik9JDjltAH5jpgHfuuGLIOX3pJJCyicG4vQ
bFx+ZGA+UCr0f1lrme3OddO/UWOMqTFB8dcuqG9e0NmJBYroT0oui4JTPjgvazq3
57yDZSYTfPpYbPwjxEQIIB18UNZVoBXgRPCK0F9mbjvtjcK31Xm/iDo2+gy18ktu
daXaaSkMB8ltlmOjh4bT7ES7xVHWNBm5TLOPMClN/i5dEUJf2H/VGSBbvnkTDYXM
zfOH3WvnGWhfyH70NJ8kpSqYhdcJyCRPndtCNkevRTqe+5t13t259mNaouQW5FET
ek80dsRS83QjPkCHl67GTehYlrz4fR3hIKVpL7Vgr1QN/mgGyubk8DJPRgoBb/L0
+51DEBJ2VJFTUmKT5dnrs6KZ6CTXgaz7b22A3UI3cjeAn3MZ9z+j/rkHwKWVX03K
qnsczaiLGX7bBwuXTvtbFcAWQEdUNQLKXcK/WpfTUwsWoODl9w70jpKwmjyIH5qH
QjSkDyrMYqL+GVhsWIUqLRcAZ0HI8Q5fPs7Ph3GBqK3Fn2UZMCIn6pAuIvPbOf/Z
90aioauGyynKUgyzn1rIP+BCxHGiIq1hH6Q0hv+/y8jWhWTaKbgZpgVM72PZku7M
W/jgez/bwSMd/Y9uQ1bNbXa0rGsEjumqNiLmK5sj1c6FGQdmyZ+vfGfPPSQ9mvhD
vm64qk4u8Ak6VoSQ57jIKFe7aqw/8jvtkxJxl9cozdwrb3dZEn/1d/sh619t+Iif
v8iiJPEQRTer4ZJBXqCE6Uq9gs9jPoxXe7/1FSmdWnHUQrOubI39HbthnJB+aVYO
bNCHJT+ENP4CyESzxpVsoDH9RiPpEHoaoqK4gbCHxDkfYvc+WM8oJQOYjpyco5oS
Nl6NFSI6dnjOSnFxFryD4RlEcAAGsljrEQ5AM7WxgB46stoj6E0Bje+HGRVLzrCu
cYv4VQa7R28Y/H1522WXCJvmBOqOVsfly9WuhSOBPP7eqYyG14zY8QlUgjyh3CJX
xd1y6NQCd+sSVgDTEGH4UiuNW82KhaSp2FJQqzDbCD6NTWq0vPUXmE4hyloBQlTm
qhlY3bXMb/blAE5+LaHtrBK634F3npiTyv5UfCQvaQgRBNNvvp1lxWf5YJRISQm/
fumwKNFRQqijBFQTbCExnA9tyR5BQN/wLnS7aTBl4J7RAx5d7T/eT/TPeaTGxzc5
v3iaKtxMjbp1QGUCCwhUvIdnWnPEAses6/yf+RPdJJcyR6ulfjNNSHh+URdqdgha
gT//iLTVz6uERuzVCm/VAGocMukKUtgc3uACWUKbWYSKthjTOycnDMFVSl7c+zbS
o27AO8GmepcwkaPvg0AUzdF6H2+NoSayf830WsCyY0IHSw4eo095aniJ1vptOJe5
Gjh9caKlBgjVKThBk2LZKLlEmpY1zqoLETwSqN8wuQautCNTjSGeNrLNJh3+TpGT
RgqN1P1dEwvPL41B4MGjE2+8JZOcnMiQqjc8Sl1HPfAqtExw4HZCFDzZSrWo9MD2
EZpfWn9YV8OcFQgh+nqVYNmiju/dBjm86Ne5oW6cGo+CISM8a1UEJimBi9eUVWH6
wPQaeiV0B/bxdKxlGg58lz9ytjO2cgw7W1PEUDKk2qO8eQ08TTLc3+j7eS8pn8GF
COpJlP1RaHjPXKh4iFXx3zDzjJyrQEO3uNns/Tfizy+jhgmHMlj5aGFgwZpzEL2W
8bww+87XeKltczC6RBnkDTUONSM/dn3RhuFqSQVdLHW2zcTWKzd8g3FUMP4TFHIX
PmORClkR/yt0oAHStdnIoRYsUu6SAEMcfYM/WixuRzEpQzkiuMvdbe+/OO9zjbcx
CadzCnE7JL+w29i7n/J1fQ6c4x9hJJnAt5rjWv6PERTr4I45ZyzmJWIAsf76BRlK
9jBU2NcN5y4T1QHc0ASfQ1mgYJ2Z/U5AvjA4lvEgX4SJcgO3WG1h0ZxE37YQH2E4
k6E+I9iKultlI3kBptstfSS/RkczKIKXbRrFLzuRUJrAZ6IV2mxYq7EuhzG5tbFf
sjapZvGmKPIlQbFYRiOlVO5uvSe6TaISuHrJE+8uuJ25CUrZVLyCqoOQaijaIgCr
sF9Jj1DQpKbP25z7zm9skUwWZSidZzd/ztpr97L3Zo/TSGZj1FEyaLIYSpcJrWRg
hZu2rEod7rSbTb+119PfOdl0bVPSQjCa5vTY9fOSnH3NGERVgsc+lhx220TMN7zx
9A3PTdnuuM2WF0uwliAyPQv0AR1HHJ9DwHEBAPEW/vnnZvbfPhzjEOI9331OF+9y
ncZ/XXRE9tJ9dPKwjX4kMpC//zsgy00NVXMajy3kvXKE0ew3Xmj6G0Awm+PMvPGG
QE6rSmTpYdhQEvYeRQzrbowyc7wDgTo4lA4ZRBCXv8rGicLxduNHe6np76FMV3Mn
3yJMvzHU/5zqO6U27nEmKfGZGsuDy4+xk19+rY6e6iGaOwg/l0oAEqDmlhKzuAPA
sLOWU/Xw387Eh8vqYxVhLDMACqbjm7J4XKI/mn72yN4K3gk6eEfswRwk336qFV+6
tCHCWcWLQzBuuon7GYbakv6xuKbULYgs4YbCLYL1BhciOpviDmd82Oqk3LRlFBWT
fcHVyRJoumLq7bP87wwkOUkM1Hjf1Qy76RNB4WfSxTvZnvWyHfOWYcfp11uzSa81
frWm+xvKBJQjzbYc9b3alFTaeE0pvFh0NExYZ4ytzJFw5vzX5updEjXLKrU61n8D
Ua65sOK8pyCFjqSrNvKo37lo9nPVI9nat1Mh2YxWilU0y/pq9+MSrp43GaV5cIai
j4VxVwldqDLoUuXCk5FSNYxFKLc6sIoJbfavPMV/vKKdGM81JFFYEHy856/EKi3x
rZ2tKg5nbJTFyur2uAasazlq+yBT1Na7f3AXphZASZFxzSs/+v7R9PHu0IaOARzb
4X4Ic2fHKN7qvzwO0ZoL6MNsqkrfSgj+Iz1lRw6qcLk42Lh1+Qp96D9rX9PpTL7D
fih+8VWYwjrNeQokLMlF652aJR2uCQLQ3mWYg870o3oSgF9uKimJgGsJvVuuVp8Z
mkEEyRQjOqgkZpndwoze798O9G+SoooKSQ9Or6BoU5DZZVJMwNHmxEjYdEsTBMtR
pyIxa7cuupQP1O15CM/NGmH2Q6BjZNVkBfoCa40HJjMhi2Mz3QtY+i5bP+zjOI2u
zEsVO+wCGLdvP89FusfOgxzO37tZGvfErC8zXApscWAIOFVR6MOoViEG8D25tKbC
bwKN/LO1RVwqKH7WR6CEmI/gUHnnwFuYR91e4WZqSHDun9LWCgQNv96SVP7g6oPV
8m9HdkBiTSZ0ahF9IC/dsVOa7/l63g8Tgno8qrvAt1xGGtkeOTSoKOaZ6mdo96ZB
j1x5kR5E42CzS+v0UwBUh7xcvQvzxofn3zAhJQ/Dp7e8b0EhdqL7llsWLOUMT3Fo
x/XGUm0YkpjvQveGBqNRTpVX2SPy8wQPqvXW7IgIghTtBBya4O4zas37ge+yklmH
da53619bjWyD/fzqEKnh2VX1Mw64QRjWK0pgkQjcRB1JnwlAj4cBaukNc0ul+YH6
5C+5cS7a8dSTG4cUUtcOkKcF15aosnmo0Phe6sLR4R3LsbcBDuw7ZJQL+ThKMHj9
6grc97K7z++vce3mjGhzzNx3Z/cfYd5XitaUlnzzfJVbvrRXYJGBlFXGJF9yCplN
ivkY+lqToyEz+RJXrJ5l45yaI59ExvGfPWTV8yeqi9RU3vjm8CSRk55SUKfPV1rO
0UDUFhcJZE2mEPsvREPa8E2rsa07MHfapTFgR69QNJtOBPcW62TrrZC6M9fDG/6j
2o4revgy52fEYLkz03rM5EA5sD/B4PzKLZyXKdyU4T2qenglzPZQmLI4OI694+ea
hbSobDwaOitRTRU9mvDzQoMPD9Ao0d9/TKaVQ12d52vmOHrdHjHUgJbUjqtOGXaC
AcSNuzqYq9pdykoIvKXQQshBfXVo+W6OSSq6IyOpZ4JuEosscNfLa567xPz5UyPM
RfeCRT0p7MGdQj8bSFuaCHiqEnjEU5BVWXiQPYjp90UTqgpQZg84McAQDa//WoWP
gUSxd43+tGbwU7rc17HCt9iwT+5Ypez3mCv4TS+vvOhm8AeuI9PBXSzjhdU894Z4
eyR+jbZMDXUgtskIW6leBJ6lWaDNVtQWY9Vu9kXcD6kQdO9pm8RB+mtBFfDCgFQ0
rVtRtfNf+wlPaMYTv9+v8jeyJKpVMjikex8nhGNhF66Ni7UM4p3CDYM7ftHB9JTx
gLiwQLyzJQ2dtf3DiHtWGuV3EoEj6AqZop39S8XA7T/kb03kW67iM2M6qAqo40b2
oHEkkkSWMOa3AUAmiPYB4nIVKvf5r6hlOoelYhp1UwtDSoIT3HT0A14j/2B7MQ0X
pyGJH5RXrKknWVYg3WzReocfwaK+qAGub8iEjIlmibMKO5Dn7DaHZsd0IerOuvLj
3geFZLdLrhdESsKGbCY8lMQLSwjzSw5xbL7ThD9CiXI2In0/3eE4wJXjISzsFvnb
VyJvv8Ndx9fgtTKXGlrMa/yqdn/yDp+fafKPUP9hjZzqKEHCEAdJaCslQrj2+AOf
4FLavF434Oi0yLldXURiqS1cDOYUmTq/sRGk8djMcxhr0jC8Ygc3xNuEfn08oj1D
oIne36sDS4+ENygc/bjoAQIP97yWPdmG1+CD8VyZUGX48YRuqbtbMK2kGDOgz8Ft
CDEVuxYdhT5amIYrpL+/SfI0O2t7GgRLPkir5mvLkRNyKKFeJ2pYy9NDaGcc9Lg3
JgyP0lLu0Dcigjo3f6DzGZu9xpMkr8rPmhrF7davVDT94pIU2CrCNKa4XZKJR/3I
oAJ6/LorwH0qzQ6QGpM8E1H/TjXXo0RJzeLwi0itrZux3Yl3tHE5oiVnpeJ9ygiI
nisziCDheV32ApCUrWYwAGzFTaSsManpSwdBKLsYUUvamey6Yx8XDd8cplSjIXnb
q5YLumj5rBRB1tQDcy7dtVajhUvj9CZ7AE0B4NULNR2OXg1vq7BSscY+dYhjMEWr
HcI82PRQ57o34XxHKDnYOgwx9gR0nLgNz0xZPOIyi/ywjTuvzZYRe0iI8Ad6IEdx
WR4/5Yp0SUfCe8J4z0Y6YalnsW43QojYal+odSAnflChGt+6rkhn3Lvnp7QKdVff
sEmMO1BMksJfYPxZn9yvwLWrLDRENYAsApMnb7YL3Ef9hfXZ+UyR1riXhn83MjIj
m/qjJw6G3ZumMx0dXyjm/7Zi+KD0F8sFvmXLItoaxOrawsxYY+Qm4WeZgMQa4HFh
RudbIhJhYhzBEp9c/4b7L/pzdcBVb2WUk67WSpSINhn1IGlQBji9cWFfG3pICJa4
onq1/b9kXScuvaLrMi3FKjhxQh6UWQH+VMF9KgUvk2meWeh8M4D5FpuOwKbAdPYY
0gFDoQzFm5F8sOhZQwtPuVynxDvm0UNYVR0YG3rwMatfkfYqmMKmRqDkNrEjcCvv
KYkOqpakpWXq4EfMGGHf7lqvHatljz1I9QLRiBzomtsfFkX+bqvQ9wo2twpQX/4w
1Ugytx1TgcUn0KPgLA55ZVl/1WjBqmMawy3s7sAIH8/orSiXhSq0v3b6YCrEF0Ph
7gD2yKs4mvTJrgCh6Z88i5LFsfOrumb0Uf2Nia0r7hGeyKJhHh8AdjkfAOrbpaIm
hHTNKsPoBDHKEHc+fTyxLdc7dGM5MkunhSjMYvr9wkPy819cht8QVE3BAi+ZKPoX
vRAASJbcX9x1EJ/wj+MRA84kS7I0nd8SjQyb274tZwsVSKlbDb3ucyWXGhF6Kjfp
nQcoYmzrsLPASlA6cvl1tXXU7S1eO+WTW+WacAiBPQGAcAZ1Srgm5cYNd3iXqMAS
+x6f83SZOxNh7OZCFd97kU4SWFx6KvQ7mDmYAT+BodMbQOYXK4wHp9fOlEVm3zf8
tAotZzBmJpm9tWu4+Uy27TKgknauYQNSIxjq3Jy69wkuziYhxCPhRrre0pZxHCFf
JrFcGdKq7XfowYNnIQrI6MmoTMdxFhC93QjPLII96yOmQswJnYWVmmpIM4i5Wqzi
eBxBWGm/avwc+f5Ah6KdHiuDGWhaaKcN3LqsxT3L0BRkB0aUo6q2B3WlsjLP56wz
bFG3mpFt4T1O4czv/7j6nCuNoEhLVVSkTtAZfOBy3z6Mc+eZKzgQSLudYTrMtHMx
U8cmOL9UgiqpLNxY1RVXeHkV65vQtvfSbCtZarDraS2CN1Zzz14uDeHvdK3vfAnK
n+6uMwhQVaAgdJcpCt9w6TRU0R15/NQCL5zwGeXx8tikerybLAG9UA0+CLSM3N11
+REEcC7gZeSAHRRfYyUkwDoZ5oVw7jTNBwi+vMbschtzskdKoQkHMZetF0WM52SL
pUiy3ZdQkQvFM6mKoNmdzZ5zzwLEGigQx+I2fdOceCj6I1g1FclS92/6HUyeVlfT
JTX/peSeaOcma1HGppU559FSiJCyWzvE7o4+79dIWmw5BltyOGQ/Go0A0pt3xDBN
wHBPZp4dSnjUWdo+tMTlhAH/WgYAEiVUI+gX5NFFhjO1Ee9k58X/hY4gfhj+ILjQ
3KZFtU6JE+VhHJSMD0nGe9byaX+xECHltY01fMYWArjG0z3tNMdu7p1z7VFJ87Wa
5/yx37U/hhxRbq/2GYOG4GkGmHsmB0O506ATHeNy8Sxm8RwzEbqIsn7W9tDF7Ah3
T0AziaE11ARAcPP1FqTJvMYfjl0Njwww3GVEPoyQuGxthGw4iucVF9H3fP1M9fMz
DeQgeUWkWOJ02lOuonAp2WNERr2HvLtFoPRB+m5DBiagUI5CWLITBksTi6hmsZmt
IWeVDWzCRpOzxglHk7NHVdRtEHS50Wx3fhIOhbtFDnltL9zOfIhHqF0RgmaRLmfz
nLMa+Ea8n3b1qb6EmKKTAwZ5o94sst4h2Wm3oVc/FaHgoAbFh0p7fcOlcJZkxYy8
9AnN/msPq2jAla2TgWA5c44wgU6Yo6oSSxQps6jifN4O+pUYZU4649Fp0NyCrzXe
cSEYPZHalreCqfnqiEA1sMzksqUJTLkNnEftq6wKMDkU6p1oeuQr58mk50npBc7E
WHDvvFIfEeTYfPGE6Fli634TMG1eIMk0WJeSkNKWumJTZtuvf0qAgFek9JnuuhUz
CkT7KN2d5sdvmkBHiKibxZLwh2gKLfpqzjG0yEWYL435R2HKQY7TmifpPCEbfftG
NIq972mFI+nmPAUbqMN2PlKYXJELKZMUrTwr+5TstX7hH0zUDXgT6pnE7uzWkUhu
mFNNOkZ/FQSCTvTgSt1Eu5wTA2XLQCxFduDg30T4S/z4vp2QeXbClLf1KGRaQox/
c7Ok/LSulaywQB21sEiYtOuuBBBbt0l7EZZCBE52xxEfU2q8gvfYdoD72rK1c9I1
lRlcKcUZTLmpDsMj4r0tklbNuMIkPLJ3VxWdiET0qTTdR7r3CKGvPD4qA9PBFk1p
lsWW34qJykcYhE6nFUapzjgK9QnWbh5hfPJMfUIjW/IfoEhlEBN7mpmalxsDe5+Q
EKRbNq8/ez9XA9A6H2H92RlyBBD/35ZxcH6fmS51zHjKQ1QjQBuUW2pB+yZWiDlk
mR2ko4sjzSZhrFlmOuFD/V85pVoCwTSP6CtxrzBmieFb+a5YTDaP5f4PURPV/QDA
KqkMaJ8Z6gbJPm6ZpPg0Bpfy1CpE08qhiP5rwxlznc1KWx5rOMmg/b8Qgo4bZaWn
0Cw03sRLtJDlK2/ZA0yvmXln8IqLF5i22bt7pmUwRWBhnm4OYmBVkz4yDft17Yae
5K3htqB9ENmNRyjUqW/6/qyfx4wLtOtkip+vmchXK6YapdlSce7574QGZ98IeDiT
+ZDeiU9B1YUBPBXIKz9RMWICAxYNcY3QVVBmQEwH2iFOugB4uyI8OUF3AzkiwvNs
pvwNBRfDExvoueZi9tnfnvQV173fBOOlcYJ6gJue265RNFZSeGaQnHoxYhhj3WDc
vibhggN7XDWvWm/95iZq7w+kA+0W685YwKWYFN1kz4obB3ngQVt8DPZa80lSjwCx
HzPQzHbCsTpGKjNiQg6Kgoh7wd7CojmxsFXzq91RPA8sqR7n5FodFdjBOVf59rs/
Ry+2+jLnNvb1/tkG7wBf+Iv1lPc6uLE04VPtF32wLUuhlNgnhsxV0yc2cuOo2/3P
j2p4omd2Vajb/pOMikjiAb3blRDpsh6FqNc6ggKnJvEzeI8zFyoxQX65umbP9Npc
rleAPrkuU97gMxq1Ws6XQ3G6OBfV9ouSC4YkIgd6CwCuoDl53Sfyn3x6V33rvGu9
VK+1fJBxdRAoSaz7rP7drz/j1zP2PjaTYUHkC9ycuQcfd/KVX8243YYdm9xwYWeK
ZYVxHXPI1W/1KHmhzRg9WgtT4XjFiO2We1cuSCJz6bAo+AE/HXqLP96c7Js610HK
zVn1BifPvZ3wF59B3TxVM4cNV46wK+2E0ljY1VjavSSUFf40DiCY8HlGouGUTtn8
3q2PddLIoTRPJochdDYqc3qW2sLpwAP3AzTNtC0eF9/HLMmlTNtXiNMjGMdhN9fW
1vHdhvOV63lHMB5tZAe+OY4Xp7Kwv8tJuV2hpTaJ0HyJyFCTXkbKVFfAeKq3cE+F
4rI41JgVPXi+27vcpGwoPE8gIdSXq0cCgdnhHw6d4J2rA2c79RabJlDXxgO1oZQw
TBSQ6wLokR8g4l6qScexS6C+rjyd7oL1I9YYko4uRuPURrqgrYumLRqQcwpjMHJg
zl46bB4DGXMOHAVnmjSlxWBwd5LTXEehSPcVxgjPSK1VUbgqWEa2AbbpYKLjqB+0
DhxIr0oKGte7bV5939m/mtYN5u7gAMDzhWvG28zXAFgcU1Ly/evftid3gvFVxWj4
ja1c0wrtbe2ULjcwcimq5Op3Bw9it3Y6MrQShPDy0X/DVIsyNBeHv0Vu7MZylwR/
yY4sVVqNbRCldpzgQZMZaqQ6Kv2gdprXnqdf9ekrLHw0B+W2ACpzW6bxyRBgh2uX
pCS8VEOLUxgx0EYatjDuTNJU+QCwQHyF01KKNMJCyEKt19twh5DQOcn/Qu1ohdnC
TAmOp3EoJEnS3hH0l97ey9AVDbTqX2SZKmSdAtJkeKTPdz2fHzKm0ST6RNbDxFYj
N5XZ//DJQDfEF9Lf8HBGN9pAxs7buuOaWVPxFZ0YIvfvGeouiXZsURKpg3h14Hvn
ER0vW1v8oU1gERn3JsxzfRcKlBTeRuWCoJjGWyWaOIuG4xVhct5vWUbuEtwjetIS
Uo5VfKmiO1x6i1OxTnz6faDRtZ2P0PzZSD08+nh5wRO8T7Gn/7VYO2zp/yGj4pwI
FZGpOS0+/XN2zgYr3oe0UHm5lUy4eTnOzJzxcdXKw9BxOm8SRccMUhcASn2NgFuP
Wz4F5gnbx0suYLMJe1ci1ZhKqaIAeM9aKYkPFipI8kcOL10BuXJXT1kwe9294TQX
QLiabaeAJZwj1p1RO6H1dCoCv/cqzu9UIB7y04m7uvGUVZF9V+3x2TzOIKcMT/bK
R8yJkSVu5Co7+lYICukm7hn2m1FCRNb3K/w37aoI6CVu1u/iHRkhP/yITgk/CoIV
GHpzG5Kv46786H8koyoULbiMPL+D31bohjZrLp8oUKlkQyWqgmc67s0V7SnRES7n
8LD3o77irkyr5pKZpGduAQHpVOOmsZC7wFkQPqyOUxSwHPE0oC9WAxzrbAOPfwy6
KTcLVkWEvRZ9mAoZfjtyQ15keVHSiBE9FplNKiJHh3HpoCg+k3eLJqK5/ZACr7wE
hlOwe2zU+LmdZt4atIlVOXSoEhXnzTrgD4DAmHc9mxHsQtoo+b4lzOSxCDVVBSPC
8sJtCNiEfkWB9POAneCJ7o1+zKctx47NL0D46VwDAhBIaltg9zYJ87l7FJCESiyZ
Hlcg+9zoh8AzpEVcsk9WtiDfhaD/0QeRYZCbRofNOAPCTwB96DgnA2cQO8LI0LH4
7qYLT5Ay7z0Df/+E8wxyQGmv/Ea/HS5Nhsdsvbkq/oDOMUfeNyOvs5f7n7TGmnWY
Ar/SCbWaxCKBV/d1ef1pfPvqrqqR781cBkO8eClFD8M3/YZSHtf605aIs9w/WUN9
sLXwfAK9kvGD3BinqJNn7xeZgmx8ujZwtBjgKyJcbhgvfci7k2SkRnv8nL8fgMo7
91opAPTZoTtoSUI6XY1JA1kK/tF+avQdfVaWJI7Na+57I2o9cx6395zZxb0Rb/L6
XnUOHYVHF67fvHKB7tKrau3D8xws9vlREnTyiKRPCvXe7Dq3wW1cb3K1lGpVRZjr
zGRxZZOyxJ5jG61wUzE/m60ut/65YkXh/PrjrLIOBbdJpUJtQQrNfIT/Nb+XXL22
GsfNqxukbisvjRHHp227ulSGbOJzJTh4VpYkXdD5SxneEpfY1msc5GRZNJW0+lrv
OePZXFMXWjVk+SmG49iQik85Ts4WA9CIE6n/U2tTgUK/jFhVL+CUzifBJX0wjtSu
q3tn2oNBTM99OZYoZWJtHJnsN6KYvuGOnK6VUvxTwYh5a82HtJcxk0Gmm/2aRYLU
bJR1hIl1NQJWLXTwysRHWkjl4kg3T3HrIoJe86rcQBmrAvYP2a0YltjwUBSpAdSx
Ne+eK89dxjG201KB7dDZezEzeQl8pUZ+Aq/2IL51Ih2uomfauCfVa1BSkb844SMs
NITaqasOB4oTBHPAU7GcDX/9u+OdaCoXDSdlzwt4q+JqupVtjWembtX/a3+rNpK1
ennoHlJBCDbzzGeA2v223PWCSAO6bEF3EMqhew104R3OZP9b25HewwdM8Wm0wDkF
F7Y0dBZsw2vu6LMR2NyIKksrVTv1aVAapenYj12CkwMOBltaZfZTd2L9BgjOQz3p
B44Ku4g7+iWdLUD4nToXCt7y/wSD5z2RzfqSxQETbWipN0C76JExMa3/cOai49yg
04FNiBZJA05JXl0yH4X7bT4OqC7RauDyXq0lIzf9MFPjchitGnQUxD0Ah5WdLOx3
obXRmR6fIchoJ8lx/7ISQTURXaqGUwVewPdqWJjyqxGArMNM/24Y85Xq3YpaSKNR
7wi8eHkOaSWdhTo9O+IkR66gcTd/dA4S9PYDqWCHd8QnQkmpSM0rJgkTqlpEQ7KA
Lk67OVRo9Q8Tr+o4/twntVx84ABveN2yDV2OamwFZnrTxBo9dMAmJQTe/8mEIvnl
zLUUEMIvrfwB93kg7oMHJ2g0JskndA5MHupyYGjpK+OM2l+R0051xXN3YDNRXIuY
l+5oxMe+dFxESwtFM9I6ulKjwHw8kACbJtumP76JNvOihXEZsqUIWWncgkfDkTmT
i/xYklmpvt1UDaIZFPnWsblJtTM+HqA0mbd/nBN5b2KWsOLWNI/AN3Umcu3HW8aO
pqnH7+PWGld1/U//ifKDjAtQOHZB4Rw1+S4vvQ803x9O2UuV0oWJvqYs59PBwlVZ
HyYRgq+g0NuiQ7BuoGWLYTG+QXjIBLxi4RlRHvZGwilJyyHrifYOuVjfQt7xMmrY
k8BrW4lVYmSU7D26Dl9TP0ow5h3A6nvOcaqFS+newjbYnWwbiXxodGMJf8vBxG2X
v1eSTs/U3wfZ6GLUVfiMAwVoXUS5VH3eKhBaW7+Njuca35/9Qsh1ZobFz2gCw0ub
VPKr1cLVLfkXcxs6JbVSSNUMcAAnQl0dwIPn1iSJYVpPtb6OLJBkSb6f1Q+/1xhS
ZY0ErbNnyOFNv4LjP2vFYPjFB8QjXKIVQaQdsiUFHpek/9K0CmCdo9QzaR1M7S/m
k1BHwK+m2Dd9GsLPrg01NQjpoDJXWfrqr+CL6t+6EEWBH87OjajfmhUMV6rymnOv
iuVOnuIjJAMCN3hPizEA4PPwYHChSsh69PoMtsL5Jeu6uIFA1+y92AXlYyJWg2La
uYBi2TVo0ML4W19e6uHSHTy34DVtz3KyZHmcFvlycGSxe47y1qo5jTQ7c2hhIE8D
61902mNrmX62/FDtx1klDzF5tc/qNBppsCX9MyyZd2OuDIPXwCoc6L28SPdeOkZM
9bLkQmHStfu5LWB1HmsUaNCFO2nohNieDqrIMy2P8KkOHps31vAoyvfa89kdSfu5
9kJFh9M9XFtMTSkSXPnKtjMtPvoTJmQLA2beDM/CXDShgbn6zst5h9kc9oXmyDFe
ElJL5jJyYvCVA3MYKuXUO40xg3hbUrnc64K7rEpm785BvjFuF+v6FOf3OWscfJxw
YXXc0lrZAQ5pqqXPD6m7Q0D2+rhmY5IQMqL0zuWT9VPG/JIVnzoc85g1DueUr6Ob
R/S01Xv7BvMmkr0bNoBWPlf2ws/4PzVlU89Hms0BXH3MV20slfOG3LOjVfG90LOa
0j37C7LQo4veWWajWqeSBfXjWvWLfz7VmEG/dWTeo7Fxojy14e7wOL9Io45Gj5LV
ooouqrRaKWgk5KUMNepE8yZRVOIk3Qwv+pVmdL78kCeDYEaeqJfwlEJu8XpQbKo3
SZq4Qj0J1j8Dy0pL0gYHYfeN1cFSr7dINFG1jSZrCUkKtkW1DnN6JW3RB4tyWwjp
tKJ/DoZySe+8bdu+DW7uAlrfJ+JP/GgNPzGoMf1VsIXwQWm+d7HPNuXTnSzm6rqS
dvVF0/II9txLDU435AbolwowIzW2rCb/Abofr6E3sQv2j66Hu6ZUddlLjEJzhyWS
xbx6V+mJYGI8KOQtrhm+xj4GSWrcP9oTCIIKgu4RjVXDjsriGNghgHp9NfkeFcjg
UxEOy1QiUJZ/RlFNbcAPvhkDLFFjpkDy7EWUSLKJZCLZPHtduMKbI71gZsotZHQ8
N8y4CUHKWuATicE/Ywc/SL23h1WU6LaP4HWOiP16A2IVusQOUu+0OlngOOzl/CYc
AkxAVaXqXdghTeqGD4eh77iBzj4rft1fHM9o/qx9bDCnlIfCn6Mg8gXSqUn08jzD
cFAIYvebSDg2vHisD4K9jkryFJVCfZtLEUCmv6YUdvPFWhd9sVVuEAvR6LPQ5pMy
uCN/iXdX2orc+I7r6UfSRhc/s7s4Cp+PTCm3pV6T7kVQSXiCsuXMbIKbgl9WdwQ+
vtb/afX9HPibp9YDJbAEPVgM3lmVQm63T87ncowptEAo2IY9odyshj8nKiopbAgj
FHdkARmsGaCiBwJlJ2V936Owkqtzd8P0/d5i1X1ZGLA35tQlMg9OS/+hOBqilUkT
j0FyDGnIMemKTNIbDsBVXGjtR4NEoAyOnfjWSlouBd6Jpl5kpGljcsY13uCOJ7xU
MptWYuOOPe0dwrsCJhD9SVuQmvcsXOzqiCAdkH2UHl2tYRd3ryRMowfBqif1KhRA
Z7q2M5GQA75hb8vgXkzketCoIjwyRBzQfFspZKNY0RzyDO9p/8ggySF30P5b7BX2
0JUMvBYlTR8JwRM/Bl8iMIQ9qjbKmW4YwwCvnQpTDSqjCF+PIWIirs5lGir0CDjI
+Cbwv47AbfzOifbNDGH+KeoiakmFWHnSQWiovQK4GWex+vYD4XWVaLRXO5l4xh24
Zvka6KWz0TFWrhnPdCnRKiQIMvg1xu7Eh4M3qglQWU3C3FCOj9wsXA9VCSXwHd8P
wugchLTlHLSUNtIf+yBQBJQcPDdoBYDA5quEmLha2J4AAxhWEi13ExSOnyblA8qZ
M9jNL2uHKOBcRtPVEjI+dfeGiCzjFuZWJWTosyKejEH/v4n8N06rCxWEiGt4U21j
6hL7vhlCDakZugTvtKtrhhENTZlFAJRjUrLi+yyMUsF+lNNSTWluggoFqoJz12UR
3tfA1UUY3SZ6uho0eQPoX4qsDZ+JjT3RsK5yVIIwoJhry/FZV2+7Y5PrW0yamHWh
z4OUr6hpgcHh3nGBxbz9LOWirIsNujDFG6pZe0xHcE5ZVnkA3pMy5kkRnOfwWA9D
+Hq66Ne02hhvrcxkbAFtFsPpbeZokcPYh34RC8JKafsxaqztkG24dCmeISu6WvnM
hgA9XMCx0uMB2TtlkgdANIlfeqzxTtEGuqXIS0jjb2jo3iWymv/tLtwHhzLKAQ+4
3P/efXjsrW4fNgSHdsf3kFSyyTQDKu78kwsGa54FmmMUitJiesIc6qfrwKsSfWnG
Fr9y4Dc+OzezL56TN3ErfxeJaZU0doG2MU3vho5GL7api9z1ZH0zhWMQIwF2v6Jh
/zTORW4qe5Bri/rqZVb8yRIZf7C6reBoG8JNwt7jhNNksU8HKch56/sokbfZ3UA7
N8rmDqkvMltkxVzjlYDb5xYZDK0MzjUaBbhjD5AOfyyQ/SwzC2hv+l8i/f9nWuUT
dssxpwioVzlHSfAJ+RqNcf2Xa5Lys/GmrLRNcIIEY6ot0jzW3nzTsXYtiuPsNQd6
+2vxDuBHkzvJFOipG80wF6qSqwcfPYb1QTOQYVEtq/UVp3yRahww2wxscNQpRe/Y
EA/j/q5jdE3nr0cTYSCwfRpVFyDmASVu1+W0TtfADM9G+jEvJON7J8B9QS+c4yCY
eW9AJFbHqHkn7h0OKnaUgQ==
`protect end_protected