`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 33072 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
N+AbGUvfDpEoMIf7wLov5Us8URR98ISoIcveSjSco7/yg/uhTIfPvA8eN3S6Dfmk
+ICLc9GjkbQmZrGC0ItwvEsRwa7NbMYaiBN49HhCcf3HU9GW6tI2636D3nldTXIa
5v/KwV3pvhykZL9SGttqut2RjtS+tTTFQY0neb9o3/xfYZaUn5507gc6LTYsfukg
YChd2qcH8EjHTN3toB3kNlHsOw9qYHL21shYD5kBS6WA7UFqWAH1MEjNKUpaTZ3x
9tOcf1aQnA0fzKh3v8Gc93bpDYZ8RUD3raPtpl0VKAHH9+Higi+dSKlON9iF9kXX
J24i47AANR/MhVPZhbNrUEEUFUyEe5Ugwyv9bXpS3EbdxSWOqIYBy8d2wYHJ4pgp
mb2nkqdH9ybd5E+U7N+xKpnlAarQVimoD9eZ9pwylAuz70XERlX5WaQwanPh2Y3N
rYFQmNR+UqMU8I0zYsL/Ba1B/3B0664EL4YaQYCPdHMGl7QHLHL/sfDargCp7nyk
st4/a8Uesqo+rfI9Q7T90vDyIJoyAnN3pw/enqsZjOON2gQm415GOOGikJZ6spE0
lNevLg40SpmW+3OLOCdyZG/aI6mZPb7aO5QkqSzRug5RXm3aG/MHJ7Vpl3t2KspW
SKLf4HOtAxG8ZZl70w0VSo/KB2QHAsmwiRil1gPGeEmdWdMamQpjvnUUjq/7jUct
fL0/LtVS0dqcF6vn4D8oV74ZV1uEecOIJkWhxfi9JR0Pm30BJo2sR/0Exgqtl7aa
f46iQG4CA6gXQttEE3QhB0N3MDaKMhSAV4ZDsT26wyOJ85W9Rlq0O9OYU0omXPmC
gLy6DJedBr/a3n21GftM82Nfyb7x9nqCZttt0nneW0D0lkcvpLhBrBiQUgG/RI3O
yvEcTq131jIrOYIbHzmiIvCr/kzqUChpvxtaOkv3o9Xb9H6V44POT01yFj+f8pr/
yb7PSnSUM+lVQihvCHXNUK/ils8I7Kn9+0njywIIFYPOvUbkfUF6yvHaotoP0gDo
HUWcnjYiytcKXzMXf9wJ/QSpHBNdGVFogJ0wJRTRvA0N1Y9eRvaskjbekE/xgF9a
C8nOkKqo29M7L0AvUoT5pnZ+PlsUPGUzbzml77J89jWnmeFopqXS77xR/tmjiqPP
jvSGUDR7hxzZVzBqUCtdpMm5devqoAkyqYHcTJa7o5IwYUveUUxjNwYKkHsc7UVQ
Eo5dIW4cq/UNTlehYllvaQJCLG4kA0VMBpOkdEqVj7aFc6KNp+GInYDDSC78Idmp
YAEtzdKBSdIaaFBxAHaYgLjuc0iy4fAOer1ZBCEXg9u7LEIYgTLNrVhI5/cnjtU0
7mR6Xy6LmTJL2uMZNf6DyfwsMrx//EZ3bEzrEgHGJeyehNayhCuEyrmUiMZqwVpO
A82B7fq/0SvYffr8IY34t26/BG1ZrAUlGaFUc+vWmzcCQQmK5p8fevbmeEl+4ZyJ
Pt6LuEZSp6op+5dbR66GwwJXvneangLHyFTl5/DyrJ3MqTiZTFhQNR1QE1f4gJY7
ZCJPd9q5JGRIckP4jQtdtIrS1xYfCFuRDPGtCUSa7W3Eyqv1SYTGbNPicQzQyKyz
BK5cQ74Zb1/KdqIBwUjHdeStwbDZxLmbIfgO1z0qXXKfb/FfYVmbujHzbrw7bLVX
z6CKefJTV28lHUNdS1qZqVI7esnfxL2pUZvOq5povOZa1X6PncAicoMAYG2ma7Sy
0hWLLVu4KKK9byTBXyYWgmrGH/BAA+UFCIqKmfZVHaXkOziC/RrQ2GsvQgPtVNID
PQsGzn3J3PwXkNQyPmAz1xyp7FsNu0G8kdJdyycY9GvDLPZakm/8ksc3i34yuP9H
AVQLIxUNcJXrEgM2KV8S8Bw38aPgn9ck8x3/bEv1EB74TuHsBF2gfVJxMSJx1Hb6
WUcVR7reZGE+P1qWiVaEvvP2GJAm28Nt60JR1rM/ih62+4bbnnyRvoHALYuAWx5r
JyRsM2rH2qWMosp0vcnIv4j/i7fpFe1zKIqIqOpc3WZPMMVCdcqBEnAZzuSUI8Dj
fVh6tIyq3WowGr0u4iBwimDhNMLjF7hqbXeRsk2o97NC9mdDEPekTWvKUQ9pmNKL
xDAyUTRGfQLaOFwH2/M0LSXuXNg/Lfk9xIkvoxFm+Z28DMmpBpXMNwj8ndKXNFOl
ZLlJPd4T2TWcdQ8xEmw+TG/DB9tHzxtLjQrklgg3OHVlmr5BGhlJatLQbh5dFbCs
UpSYQbim+6RVwpiaPyBGrZKnC+ID31oPJnm9jRpm5og0aMY/dt30OQ/9pEHhFdU8
HZAWw926lFWjfT1JhECeMQqx3nuqBFXxoKXMdWC0TLw3HLl8oie1wYE834azqUhF
8GMLJFfb3Ak/ult5zPv+gpqxPeBsaQAX7b9vVKpmbTh05FyHlpbu6m/amEkuoe+0
VvmDP6CLDUw6Col9dF0NQj/383QWk1TDePSV+O1fombw1p1CQ244zErVpBWRhAMo
BiLdBsJSLxHdhL7ZydE9E9WPDkfwP4vhKYl1L6V6VLgsBp3lk0INOYVLv7olHZDJ
qWVeXZQxepIUzcMyRzyliHgixSFB1fFbQVB1aQ8KRnS/kmF/oefvXHy48uGKN+ac
HTieZvm3l8gA3xaiNSHfscK+oQCx0sCegZRpd8CkE6Qu5uA3yPntrOvSOO73DATF
ITrqSPynRX5rV1vZYlVWRexoTavLxQtcII3lBAXySvkWuZMn98zut3Tz/Zfw3SBS
0xr+wHQLec4MBxZT2LF/WYj8BSQWIe3Iu9fTiCKgai0SR9L/Y5DpMYlr38efE8u4
DTUfMJd2wrsiW0PAUkWzbkBo6ko0G1cLQeShbTnL5LbVUQ9RcuJTW0ce6KIva+Zz
0KZtDkS2Ir5TUhP0dcJyfYcwK3phT8Ty392W3nB78+wjybiSQ8gyFvmmu6pV1qvD
8iUFjuejKYrx3ZEfWc2j/zpQddyTwhLpMye1KCZNGnwUf5fqnWPDyzt5bP5iLahH
KmqWo8yPuG4aCWFY5OUBdPaMv8T9F1wRM5iWnbygknRWyQYp/ZUmn2BHsIN23TZR
talL11Zv8CbUb2ljZEQ0w81XCSTZnYwn4swX63OhFaDZJpxHfE4CM3BdSX2G2RNK
IfJ9ToIDqTIjqOF8b3SWS78AAHs2wfZkGpN8NUjJ9LRxNGVDAhMY45srJTjNdv56
1YFgfViWyWi19eEkwUxw0zUGJIJkGNNn8tKpXPZ/IXC2x3OUu+sDjH3dgAhgA3Ua
6iY++8CA29CWE9YKIgl+1LLz3IbjloTatqWWBzqj87Mml16lRV+rocgOogEb+slc
z+sam3z6jgy3s5xvI1srfe8j8LsjzghYeNGa5F1bhiRTOVFvRuN2GVN1wGf89eOW
DHv15oP43ZakUjP9iEQrx7Q/C1Mr3e4fMDGdiO4K9rvewMUFsCK5KI83XvSqVNxd
D4pulgZQmNgeEYYRDqqbvETBmqrYTvx4k2BMab8WS7ZBsRdGA4/0s1FKP8SXPv+8
es6taVia+ucEV+oC3qs4Cyw9bkfuVnRjrlU6iuXDIZ6Aq6zG6ZLvUo/TkhGxbX0o
3QUh6+TBP8DOg0ft4sfY5G5CTFGbFdbHx+p5NhbFHkH3SLq4GWdC/dKcpv2t0oEY
EKZkiV5GZA4ARjS9aI1IZAozPEOmpXaMkxlPtcfs7huKySzXRXHp6awHwksTq4o4
oAYm5+0MV/sJH/IwNdFWYe4BKC7abiRx1yehtWflWQ76kjJ981pMVxS7rLfkmVlM
e6VPV73oX3JDAxyAXrzk/QxE03a75SSMSxZSQ0LsPp2nCeAhQeVNCanbG1roIbz7
1BWCd3Vjbad1Dhw8WQEguXPfVHCny5fIIbzAmeFZnH0hJdxB3zFWLSJJl2DWz27A
4ln73mhhX4oyzM7FlFbpi7bEVxgqmG3y+3k570rtQc6SBvHw1OQq89XpE8xWVLQj
NVvGZiAJYJwBzBk9FKHC5pOLmEJlFjezcuTkkOAs/pQgwjPgcHzT1bfKKXwRBdEl
BxS6Ds/c0hlc3CMeqwH+VqxfoDjO/OeFytv+l7XfN1ycQM/SMucAoMrusWKA1f9E
ODPDnWeX1Jvo0jZY7kvx44IciZcwwYX1q4EbLnixKaDHiSShP5PTNPzfKoM1vi2S
Rx1mjUort/+4H4EeNpP329Xu+P52wEOCAs1oh5EoAjyKMx7TYY0e9q8XBFWwgLYt
9OwAYhL+0Clq9W7Kg6eAuZKagQsRHIWptGWjXjRZEOoxuzLqNMwmO9RLaZ/A6w11
2TqTSmfZCp5BXfThSGcV9BAzFsRDFweVjUtA5Lz8Yu7oEzBuxGqPMK0xTp9Q8Z8V
7b6PjCGqCLYTNqB/XkH1yd1Aa+VfyJmzgCoJb7qY5gXf9XA3z4czD/Gr2l/OHU1E
9A0WwEu1IrS6HfAfPBGCjAOxP3kUSGjwJFm0BDgOuzhBKM3rQQIb9nfmr1A4MI/S
iRpSJRyxdJuqJgfofjOzy3fL2KrmNFlBvvrV6CClG1jUAd5+EZEPkNdMSTHrto/k
O76wdP52CDOQezduK7G+NH4H3K09WBYysWzQpR55ZPHrAFfoMsttZCua8TqJ2mN7
PTAUTscFibPupPjbvEZkqsL5073yz5/Iz/ApNG5a0uEilXsux5GreY+LS7fk+c8L
J/zfLCwLHz0QCDn1RNvusWI6ZD1RFmDlEjrhSRl2OBG3mwLyFbZnFx4m8nOoNI+J
lSR0tNYU+QTIDhg9q0cfxUttYYbxAgH6BiV/wpcT9NuHNVIFnpv+/gehf/4pZ3GC
1HrjlWtWRxcOenzBXXBiRyzIwgRaSRfjxcsALcIH1mu6aVFs1qgivmJ4SyY1DjdX
BsF/TMa3xsQxMmP5grPt9Sdl6iqEoRC67tefAyHIWAyQKt/rcOxQp1mNr1J4iXBb
GRiTnq8EwLDYrFakU2+wbedDjzM3VxbUuCjqLUtctDGuM/5Qpv9ZLw59dN0Qf1yY
oFsVQfQ+U/QyNAVm7WgVU7A+d19+Ga71awnQ0SwDyVkYck9bYhbYtuDwQyIBwl6B
5A7Dx45p+27igvpR0Yb4GhASstzttnj8m8sX7v0HmKUzhfHZ5hBsqiIvbJfajh3S
YNde9lLoJ3eDFjeTW/MRYGLikAQTh8F6Y5Him2G5BvEgzvFw9aRQwPaJ5fkZyTCO
bCNXWMNANLfAXWkw56n6+qg78EYEIODYvcZtx85lLegPl7XQWP/gMwNHn5PPfvCH
T53Vtosuz7hGS7qEZj6ASbVYyX71KWIS5yJHdx7yopeSABdVfKhTH4Wn5UUyxQrh
lR+aIFHGjoBWeifuOAuvoFKtSNNAUb6rFqthxsHEY3TIBwhMbN+LUKpekrOJ4gEy
SNR/1p+9u761nz7WduBQfGbxuQlq2L1d8GSDqPioRaKRYgi6zPBM2zdJvddkveKX
a4B/pn6+ZYtxTc6XxCrKiAQT58+hFrKJubqYeiMa/IPYJ/Be9vq3LFMULI6TVHsu
yblTBUqdxeDefKrJPdEN4qE+HWqKD1eXzAbfgiV5bq8lw1dulhk6/erY40ImiCG/
fJfQnH6vMH1iDQduXxdlB0fIO8Y5k3vbhujm2miSxJqfmlY1mS5I56bTgSKS1PRa
lWt3BaejA5T+wtzI2fXe7xM2t4hbi/Uyug2XOCyU38nKeCJbx0wtx18xUF3O9am9
YRGpiKGUaeYg1IaVl8ev+GXcY/23gCIM5t7f0QM1/f0LDdRRBjNZjJfpTO9nhdvW
XlqQODPpbmaDh7sa3E/yqbtN/9YNv7SGNXsbdeYTQmik4TyWddPBMFlxvDdz1ham
ar0bike1+CVkadfMXmD3W9JaXL6fmw3eFcgurEbjM0u91YtyF05InUPqVZNxw/E5
rztBYt25Mu8NMPgbaq6ay5Kuc7VrY6BcQFn0x1xzHEKIUe5svDwCnblwSjJnUy2v
pVmyD2rl68Ms+TQTOB2+R99Dr89M+1s4idpd7yAlX3oC4CEVQO0W9E1UJ/UzmJnn
BPzkw75al0M1L+tUJU90okWm3GNtLeC6Z4Y/X4Ko59TZtQdAkszrazZHs9snoATK
vPQn5RcVkJmi0+9EhojThh1QHbY22/6HW+6HBcbpBpUJEaTQG1atuUH6TbX8gfNH
5ljRpSQSWH+OC1FAPHF9AwFp1Pf4qv9utVaoZ0a1hO7mnndOXXFSts53w6Io+Alk
gfZinclSiqkgRgYU4Ud74FQjHE2t/dGKEw2eMEghS6JE3tkAhGepDrQd23tq+5gO
lG+6p+o5QLchCv+fZch5VdnFSVhBoPFZvuMRLem0GxFmDrukTIcYiZc4KTsq2rJV
DxVwih2Muo8CayfzoT/mFGuYcPI6oBT9g2Bp0FLIGyv/mJBI67nec6KAJxzqKoc0
cLdBYQ/DFIPuY/EBZZVXXhM2rosTkuADQl6YkuUVlB/MvI3oRUzyUu8zWoJQjI53
K07rYhoSZG4vlHzgStXKrOKe3QJEDYEoYw4hCkA5DeRwfgE1+v9zjDa9a0tSrKTg
ZPTu7PBm3RnuNyxjqLjDlbU25+XQTzOdN3adjlSfU4wTIVZHvclF0RWBAUXzWjso
t+zq89yOC/z4y2LJD4o2P3+dVUwfLe1RXwxXXBHl8GMBykR13c3Fpsz/pOnAViVz
1A7YkV0JgKbjKh1A7ypTgW++vmLGUQQXtG5QHf0K4Wzq+B+V5ZLuYxT7rkZ1O+X7
iyJ/Nut3tpEml05Hxh/csUNDxRzt2zOEvNqCseNkIEu6wQiwQNI8/IcBkLPwfoTl
Yauu8EYW/cv9lil2/7gYCVDfWDNn7d5JCB9Qe0lL23vb6o0FF2xz4p114wPIFrl6
fMMqzyzO5KDxTd0uYZCmPhIRdPm1nxT0Fk2kcD/nC8IKkCqYPPxYv3XL4c8uKECd
xEFeXOrz2Qj44D14QQmVnLPzA89/BQBOmnFLSv6qljY+NgOzgZ8KNWm0iCygxv7/
5WnpKqBD1i5dv4jbLfSPmBA8o7MKrwtsekgFNeGSRNjmGv1MM15bJsg9tvD2S6er
qMpotaaqO+h+0AXLZ0hHs3xgFwAjgpEmThyOt2hCMQsQzjxyL4I4uCVZXVVhY+EA
gvwOeskcPg2Cvi/0/ZUMlBC4zDqoZtUQGjFocQm3o2QSkeX+QHHqPYawWUVxoaH8
PyQNEtHPs+LwUEosaLiS19gqoWnC1Y5SlV1TU4VaNR0ssBCyoKhf/8gZFrzCm2g0
p+uhvZVk6VNuL+rYoSS86jEm2spuG7wk+SHwo/kspWUbjPwJCHPa4QyRRwUErbya
Ueq7VerFuQLJ4S+sZpEue0kGKJDJcWg9j/YSAW8BPOMnGdGjzLw1f/tdfyc+Evq6
Gy//37VQidWOL78qjQKas6nEaMgF5CiCESSHlCRaksUqbtWYiZtOsKTj99Dq2djE
lriwNWTKlXu93JX6BCSWFBxwcG0vSKwl3CzXMMlPzbCv8LlImbD0PII3xo76uX9S
OHdl1tD6oH5xPr4UURerVP0Rn1zaaypYFvJ8/JdwiyTDWobhRPRTsGb6Ej7yhyya
vmwTtaV+6l8+HfLGwErub6ck1/VCTDl2pNBo9aW3b/0Nwr1tFUiNYqQCgJ1uGhtx
jjAN4x7SH5IHxv2eG7b3w1/KRu6zd6Bb6nNHuQwig0HCeawLwvYksBxgxYe9/658
yvPAsE3bdChZJ7eguiavkbAGF4/QBOrSpFOpO0cRWxVPRfHrayFrgP0YPSAMxONJ
O7EpVEcsNQlQW7kPgX4xYGapToa37SRBCZ+x6PVXrmjdQ2mxxJNyddNRCs1hVbfI
ExTH5Oce98Mz5IDWFTFl3hz9i4W3rQaxhw91AY0mUFeZS4kKAPJSeAUUr5JnJFO0
5aUnp1/08iPiwgmHhcRxrTKVRxT2mSh+/MfIhsKPjbd7PEuWpRumJ+BEiVfhXfxf
/yHITqc6oPP4DScWHKawC6V/zd7XmD9ozLsIyVwuFIUNWXDGeGuJRiF5krmXhkys
t9LeR5ikG5qLYOrMSCHWVxvbHu4A9eWDgFWi7s0VXHn2vrXtWnCmtyLnl3VXPRA9
aRWA0DaQGwAa0xKS7G5OQUSV+EH4UUA0EwlqB81KzU2syuYpagntxqPxA492yXjK
7iukM033yu13TzL9/jW5ahk92EZuI2YYuk5+Et8HK5okPslW8XT0yrNhYtxLQgnl
2uceFP7iFvHefqdMyA3w/hFIWCNGK8hfXoyEvYmFpOzufCNzrP+6KqFzkN2O4cdJ
wV6fVpLruvbi+sFtF8ByNwZcF/+Mv9ZUx9lSvIFDErfWS3qwXCTU7McPOt/hqvNA
vDoRW4dplxgK2SNv6KGWqaYwx+W6smbA0H+8nMQ8de/zW+U/pNj/mRUWPzym+/n0
oUqd/jjW08kPc+LAOIQKqDL+LwANJFVH/wLs66oQyuJ1mKixN3MJWuwQZKN/Fgj0
Jub08smNZ1OavLpgjtlTsIUj4233rUlxq+xzQo472lVrrEjLlwrUm/BxxXM59Jkq
tRtNrVSxYA0BsfoPZlAUFdWr6nR0OOhbcsns/UcQlvAaGhZkB3/5BgMadZ/w8chS
Wi5ShYTVBqRVsaJKVTrGnxy/vk3vXTWGdEvdHdxG91oz5GMnV5oimZDEOgPgo9gP
Li/NIsJlSx9+8zl95Ye44UYUSmwl3jmq1hTSiirXgT7ZnM34/UqXW4WDw7IRkqrY
fyP+5Uz5z4yNIOFm0KpNF1CA1WeTlFYvd/7H6p7Rb6rGfjhjiooLNr0Xa0JUm+qa
zOWRWiMVwSMCyOCRFsZyXHgjuSVX/MHm9zMaGeoQPBpYYGjVOcToZnu7FEctFigU
QjasjGZs0nmhbRFiHZZ/SqKfbSR/HEYEI7J5FoqtzClAKZQaQlMUzgSehwiCgW19
uSJikKQgj1EtlbeMtr9/vjkWZUMXG0qA6NwqhMsrmFvj7867NZeq2IQBZIU9J3/I
/SubtokV0hUyutFsaZJY5wwsH2G7CcsX4xmYXycSaSyynXc6mazETRzeDhJXiC+N
atGJ1+l11DoFTSRrKMLVBUYd4YhCU2+NygMC0W2H3DMSpn5Noro4f2QFMFzLV78W
o3cMMPnkJP7T/ew/qqt3aFheqlOvUjgDCOgCsMhc2wtBvlIBPp7bvxRRsUpW1wDa
381ozyX7UVHIrXvuiLSmXNvEwWzYURY0tQUPRsODDNi/zQQ4+72WYzhFfb8o9EDH
9OQRGSa2v/jFfDkMfsi7Itz8KN6mqymZhgON/keUzXKSssXtNfQcNlDoNZIN7jWO
5++zvNFtn09NKdtn1h92a1QuA4M4aqrocNP4vIz42UAag5iLdRsHke3M2UbSW739
e6PF4aT6yKhyiN45ULleRoTq0N0TlGh7+CKB9fyJWCls2VpxKVHWL97R9mgVIAuQ
ZaVWECP+BAiZcQozqHTufSjjyWmMAApjvDyuGrlFsnI4Aob7keCm1ClGIOxgnVRs
16yxtyET6rx5Uh7ZopGhIy4UYoiPVzbWHCdGZsPnd+XR2RijLhLzzHjCUoteNYLP
X/2sNATNYKxf19iMOynLjRJ+ueEZX6EJwOHMFyT2iVtQ9SSzCgSN76C7jyYknO0E
m7nV204uv1sErGeAkjd10ILaMq5kM9jHJ5h6lNhZOHonY6fkf7j6Kqf0Xd3bdqZh
w3S00k6Wm4n89wlkBdGRwSJZ1ycQP/FMsF8vlz+RgcUELh1vNEUbfSd1pXNR4Y34
4zcxSv0WNSRdJbkK+tokj3tV8x/LTgdl97c7AmX0cqeTBmnBABOeWH16q1APO8OH
4SndmqyF18vu83z9soU+yDpBduj+IDLQX0KRWxaD/TSUt7ANIC/J6ZMd05oCsQgb
UC5F4BPQLZmObTa41i+IH0ADrIjxmGMGvSQxAKFIAMgiELzWlzsU2aqe2FsFvTLz
8pUnSjD/9l1m+UrJTVeKVEBwLZX83Y1Hi/axvnS7bxX1bclBoTkbgESud1Wk952b
J+d4ltNreVLM/kxbXh/+KaIDTcA8VVAeWkZpcunaQ+FLy1HM+uldEyqS6/TS1d3X
e3AJTw6I/BApaJx5wiDUd3vciydWZCxEVi2RNIwkc35W3oi5ySY2XByopy5aRwAa
MLNkHxqnriPIZfmBU24rPJvEFG+Dp2jhtaB9DOnEBW/s7FSayqqmWFGPlK3GLlPE
CFsigQ/NJ3yT6VCcoW++3wIBJ9vlg5cUU74LTf7uVxisOC1Y5EGXyVign6KSeQNL
Pc5xgftDtwsVQe4SovsExjDAQMPh1UrPVWSaY2dupfNO+G56zoL8SdOREauj51DG
W6UmMSz2I0xg1OxiULQ68TIuIXg61bQC5p6r76DAXe85osWJBJhpTiLRZaDeacDe
dZM7iGoug/8pf/0HyA0J0/NmlA/GKabRL/g0FFZmvWiaFV+ZV8XC4yIjNdE3jMPl
68wWMVnaDSo0sPJ9zQVzOWozsFppuTXCK6nHGAq5h5ULQTRVVj/q5p0ickorOwfy
Bhof/qXtOlTRu3Nu9L5L6cQyel39jaxumLuVgMvD7sBGtCVGLxaUUGt4wjebuV2i
5enBBGDioh8nqiCIqG2mUaBhHRvUzsrdWO6d40mX6fqjBY+KfvpCZGW686fzIcnO
MJvueme/agjvrDicGIBgSrZ9g2yiQEUyT005fsSl7n3oNh7FVjQ+jbkgD85cZixW
j+eV9II2uaEEFNmRYrHOetpqV2PNNnBz6zoMS0CEv+aTwMY6hlFD8Dcu38lS6NmP
gkTALCk9JE3k7uKEC0wb4TC/w4fQwMKS0LEo9MO89z1+s8BqD5xk66PG7yBpIEWD
AJ9dmUfwKeQehok/iZVC4bG5X3OBeUKbfyDwWHsXzxPlCoSLVwGzOSZm7OzAgdMz
Bltf+QV8tlZR7637V/uE8dZ7Hai/oWC8SOQLC6VH99qDA1pkSaXbGug29sAmKBDT
LRPcG5L9UsUEIF7Gab0eBVyIm04+cvvd1yn4hsOjZG/4BzaVVHmd2Iz/dh5Anf40
BS1VFOJn94PEpYn28vGfex/5D5PZ6a6EaR/Plz3vIsxcoGWoVwNkOOMDQ0RysTzh
XScuVOhjLv8hLEK2unOIQOxvMIi6gusbAqu+WweL6yFBxBl+5mLyfuPsegkR8quA
SWZTMdAlTk/Rgk65S7SJljGUquzw+NloHk/gKnNU35KJ7dkhYaEk/QL3TDC4EXNU
58ft42nbXE5eoE9fbDCFOp5M+ddhdFnIE1pGlpBiH70N9tAOsZXsqFPRNiXx5DBq
yJe3bFz/5BSVxy+S4ov1z+Nbbap6EImedOCC7otLPqPwguK72e5h+Y1RGPgWpD1u
9+FjcaiRB247uOL26tFtlaktubZ4oRs2togweF40QueQkoNtiVQSKgf+gqi0D/EX
VR357YrbiQVFtzspwmGjysWruHws+KYuBiv0BdKNF2Z4PdVBMvWvuA3TnUJQlWjJ
hK861TXZ/fwDAFsg2lMEFnwmI/p73lEv3EKPIt5qIbkHpnCoP/5ORgVVroVdpSVn
vIcwZ/VQBHoDKW1n9Hcfmf7y2R+xSw165iPjoaF304GLCYykKYglAuwV3LOGqNeR
yOOYLT5GDMYDcd6Gje5j5mdREWfNtr9V7Szg4BeeOiYnSZ+bw/pltAal1ZacIxNi
o5kga0Jhdp378nd5h6tVPDmjOLBWdkoRp7ndCu2vZDJe4UTVLn1Vhg1YbLEVT++p
+YdTxQsm/CdO3F2JSuLgWX4OP7lecT0H+tihWwqS8lUuzJ5GjdZKZkbUmD/Q1EZM
IokxLaZ6/eGf0khHoY5VopPMs+5/YixrmOi6T/kt9oQSth7YkHKvW/jr8wKGvgLS
sKegMBxW/F0SDy+LpJV04qebJpKE/fnpto6mRo09i2k3yAMMthCPrTyQ4Agv+Rfx
6hfilAgSonWvYIPtf98808pB0B31PHaCvGyHYabNQ5aiLM8YtkLg3N6mDzr081PB
RtKzpU+4SHhqiZVvDee7JbZgnfCMCkLKVIsCmfMlapbO70UIUIXLQoYq+W/oBeny
IIKhCAwxgI+uxelPAONyk+U+QZOEaNMntm1x1VF92waoRstny5q/VfeWldMUoFgD
6qT1GGK7IcMa5TXLeQIYn9oYK+cRxGafpYlwqLNRztNdg2leAd5Wer3G73Rg6xSi
Bt96Mjlkbpmj4rHQFutBjhpmxm3XiWZ2XDgTV4eljWJCa8y/kDu9lubsP3QZY50x
HnoEXemT5SF9gQXJojyPf/0YHITnK2wybbY5caD9MKFwZMtknqVcykPdTQi1g/AB
2ySl0G6nffWjAQBivL8Ci9xZT0kaTreWNFHD2lbrJAgzMJ7/FzbUqX9pgxGstkLT
nIs8RF/yrLVQfBT9O5QPVRxrRzvT08Z2aLyQxixqFm//xTEqYgfoNOdhAQFI8uTp
hrY7Sj0x3Rm08CXgvvnlyEIrPshRbsCSWnMBsnp6DE/Vg5tGtDVrd8Z6UNYRNQEF
SvUbhKi0GbU1MgU++gzOwNlCEKMZvR7RjkvXuhG92Cv+hIQVgAfh28mJcYaMNWYi
a55nOXUhDs2sBYAQiHFaY9u2WznUd8+Ba4RDSgW7V3ZSdx55CxD065asr5yZdRFT
o2oO1B3ECz1ECocixof8VDQC3Yg6+Mw+AP6VLFvh28ON4lDz+bqd2YOY40ryXBOJ
5Mjz+yzbcBki7SuQ48nfn+mjaNv9hdA5ZtRKtCEF3SvyFVKOa/oc0eGWD0vslfMd
+QhLEtgUD/8/xvmlhDqG1iWjEYDrnc4r0dg+PkSMj0ocvHPfQ62XuMPb0PyW/QXN
47EbQ80wq9bUr6Oy6Mj7dVlUCI7tyEd1F3Frknr4P1Z4nyovSsebLSVa/GhvJWux
zs6lKU1R21Y6Ho+2iuR6ag9Q6w03oE/5YWnfZ3HkM2p2MAtV2pPcfSpzhDYZiJ8D
AWl+rszbPcBjHxSO5Lf2jwRZ++k0YRKzt9rpw6vVzOlysRrHfN5Dm1D73pxuELjf
85080zHWNp20RTQtaD8s2X7hFZtvRKd8miSkT9KTniaBAza7Iplr2fSbkfgbo4JP
HFCgm+KxbNVCptsBelbJlHSil5bNhcVpIylPXNIqk6uisTkRB+hmnZ5opZy461Ou
T2wcmjkZJ9ntSRHml6ExxC8oLSXnLvtxB5Zlk+73OaYJOJEcjbyj3lT6AoK2aVvl
wkT5dQ2tB3efIKUiA3zDJOiKhiRto9o9g/V7y63ACNGfLDpH9wJnHMdML4z+h3ZJ
rC0bcL2DkXjBZ1xzjfv+vMutRfC4erWPBYvMmKIDAekw5c7j25HYtBrQ/WeCYZ8/
ClIZSFvvdaw5Cu37f2JOqlwFG0rsC0fFF+TfKj37tuRK9xZLAAS9rXqRHdMN6JzP
RIiJ2EEWNtLwMTvUVrAWmMtvAlAdGWCumncAK//QI55b1ueIzJyd3NrJ9Kf+32Ya
aF7DSD9XELnztbGgYosVedvJWbstj0cY+ORoRZMODI88PMnsnFyBaMQHwAcx2OYf
4cNDjer0OoUiogZgGUTcZNR69hK4tlkZTPGdOrRxmar3UxuGAYh8BBpuQSnLcLXe
nFe7JIP9XSrSmVopW0ZKz9XV3v7N9FcapPM4w9pmgR124y6i9Zh9xPRhwV5ctHw/
83ip4Kjt+BWxYn3RrCLsuNFNLwgM+mLrPGY8TZ3Vf+QUc3e4qiTGf97w/mbZcVN6
kH/gID8UmgPSQw67udtIg0LpxN8Dt7IMrxxfTteuKl+VBs+CJOFqmvsdxjarP2mt
wswXmB1XyAkEMsagxlQCNEEK6i2F5buA4T2bGaEpTcVoS/8HCo8XG1hcR6ZfxSi9
saMwA8MCkpI7ePwGWcF+mQrhp8zvevvgeCqQCBT0Hiy8dsdetRquoRjxeCS9Ch9k
oWCGdNTOBgrMHHVdgYPoMxiaURLPNVpAN4ua31F1xDZ6UOes1H7lzvomc/d4EZmi
3su92Olpty+Jf3PzOmc9k5WHilpDeRmb1gtqMNhuLo0kv5vyOmPuVE/JXVZKoKNW
UEXxyDkmHKwnn2z9ZoYRijuIKpFFHl/hIxajmFvZZbw4a4SG5ZHnnyYQUncgrpL8
g1g5PLKgFedt0AK9Rd+rzNtaP/wzZyV52HCQUoBnWg9d37r5XD0poM91H5wA33h5
7zPFbKvTDas7cHshx2Ki9i9oK1uDfLegSa+P8kI7kGu+j5YZOj0YiHkyydPCT6Q6
WFxR0aT0Mf+X+OZP6K83pBylaXwqa85obsEpFiKlB9ZcuBMYKc8ARg7ksBSBVYIP
yAgMw1EDaWAmbNG+56C6VCqzErwPraSjT4yRx307GOt8XspUDJdmkbgDhiZPMob3
uK78E85rlksztBVzHPD09tlyjzIP9v4dHVEHNeaB9z4TFfEbst/zGr9oSnDtBIiS
0aWV6GUqSIRU2bG1y4V4+wGWOgVKxIfDOiHB1RlJpiFCSiz113OGR3ksh3xen1WJ
ZowKZVyqUpVs1ZeySmyOCYOofnRggl1wANx6O05T6zHSSU/Hw1HdKYaBqjdbfgh2
3zMUgfFqMAbwj8FsV6ZcNqRYoINoZc0PM0SFyYe7ZgiGbsaoq2cvkQqw28sWpU8m
WzW7rYF6JaD7p35MCKCaeuhL88bl1VT4U2kNaA8LbogfiHIms6zcMGIwde9U8u1/
ogpl48rI+zrZwBiagdx86O9UvODZPSCOKg4udN9pxIXsSKfjuspExBnUeaVeYTUu
Huh1mdD9a1gfwOAIdRn2W5SkUWdY6DpnovDP8w7BuItHx1vm2bW7he7B05INauKx
zxARDynv6uOC07VSKX+1DQBBgMSLlJoNFSwKsPY6ZrP+2gyTprTupcc6WtYnLUtB
HGKztIvxL2zhlqyOI0vfy5YY0Q2R4/YkXv6agHTdmKFielf887I+KTgtkFJcwcci
WTH3sBA5F0j3OczXX9HCKf1/15r0vaWt9QS6/39QbleamEuRd7ED8fpSSpmR8Jop
QgPTODjfsst8NRdO225UXRpRKG8y/J/2ercvSjaCOs/w2a8chpijmQ2fFPAaOZEU
TACTuE6XP/hA53gh/YUJuMWV8MjzQ4U0YoFd8M//Gx9qLmddHJKyhw488v2ZnXpe
IPeYgWwtXAza8AEt1i1txb7A64384vCCME99Cclmy+smLgOjjBZdOm3e4W5bQJ1K
AG2zPUYJFgcWU+xdYgU8Z+jiwKcygGHlngCL8fw9dbkPkKxbSYYvZ9YuHOv4nCm0
OkGmZ8ewkf7XWA69WhkF34a0y3RGUTX649An9VN0fIbwCBPUEl5cR/IAxkbO4ipL
zugRPfIvHRvxamJj+ui9i0WRdv+6X6wgEzSvIT6cHt34YUK5NkQRXoC9YNlHpsra
W3GpqsVaWdscyC2Wbckd0WxtyuiOmcnJrRt2x6PVf/644UWxYvZ5DmLNjC7OAiPH
//e7zfm0nJApaGu47xw7ZSEw1ox/Sb+4FSm+cPs5dXtLuJEzxDm01l51yFwkeF45
u24emWcxxAdoYDhpGBGGCt0XY+Yw15bsdULW9IQPAx+h/mEdmeOIu13S8/bIWZ0l
MTHSM5LWbyAVFR9Pxd3Go7QxB4dxjkTxF0U7W5ZhgyhOhWEAUQ5hYe66NxSAbZTt
2cU+c6m35knpF6Pwt0xehOFs5aNeWktQhL45Tja6YWl/3OCQs5OWisioSmVFafAU
HBybIfsyIS6GmrqONKTg0JscnImmbxJCQ+qU3daLyOan0Hh6OzREOtHTnvpA0xj+
a32KHz9iPFOi1p/EZEMl5lykQCsxGBCY/zsKay3WgsufFfZxHrC29TVal62cQGF4
iOK9xceE4np1D5mfaN0GUSrZGFu07aTvlrUkrjItrU02Sl0o0LbrCmGqOfThVDG2
FhaS+JUTHjhjQbN85iEzP2am57G6hkAsLWuEVqdmaPgsNClRF2314N0qAFqIGETf
upUgEu+nZZsc4lhB9BmEbSUNcA8GDkfaFinM0pTdmt+SdWCS1PS2oAfkjjzFPLjd
w5gm9bYuf8r14corm+dMNN7sVj+oYhC+HKtN18a1lPI3cl8qObIBlNMeizCYR+BE
orGmXpOYyUPl6g1nJL3RP6y01k0tIRa0t8Sf9TUD4ht+WgLb5czX30dUmO3sluVd
AAAB8b2RxRU9HratU3PMeAstqso9NNA8b/+Ie6X3N4ylLt9zOU2fOM3U/t8Y0U6Z
wCw8P6l+C4BmIIsO60kmUMnqH1/KGzkDH1+iT3DP/uK7s65CU6hEqYSTvNn1e+UP
k6NPkrBv+ecYxZYqHTH04gNg8CzkVUq4/d2Lnujvc810N66c/BVrZuVR+R+i1TPw
8aC5gCGlc5u+K/0+vJl+vIHAL+jRFZonlEu9paUsEK3JqSXyKfItS+53fuA5ABnO
9VgcBPFPcd5nPFR4N6VDQdkwZe+Rp3R07muKa7VBvIZy41s5H1B37x17JxSchDWz
tSHqsCabnPE2Hx5srylC2LbG+Q0eFKF9M9xVNjBEdNv6tsFKw5Ejg3tSGPtLQldL
tJha51myIZMb7ZTXJOZCcew6/PqhP0O25UOBxdhwYsMwnHr6a/MlDMtjFJ0OyJRn
xvAbJ7pqC+gw1ur5a8lJcPRk4a6z/8RcF2TVAqhlGZcgmpzf3XJknu464bIZnK0b
7wk0FWDDyEBMfBftZ873GJcBKzmd0LkoZUONp7PPf5NzxZbPVWl2Zdyw+len61oD
PLk3AkXjE5jVBJY/XtS9YqKewS/+MUhjDjhv5K/WfpOsjHrkkieDsPngJcnkt8jF
dBe7sguEZKNelyXbP51HlskhUV8YzjH1jswszJb1jnemrJhJZaguAG9knlhDLRRH
uIgl3LMQ+WqG4DgYrXuJeAO0c4JWpuMXVBy2E+p8TncnpsIAsI/SsUQ7NpuJY0SS
txdrC2SHAcYQRaBJ5NgIJ41ESrtGDPDb4mXSHewsereJd1w+AsDrdCsvGGkzMjdj
5lAkzmOgK9WYOt/fX0A1tIMLl+vqzKENGG/bDfrx7NB897nDhN37DhF02K7kgJoJ
YTFnekHpEK42D9oXMozAQnlK+0ZlhkKtDd3IdMFZt5/qz3kTlaw8+xqzpanD87vP
qtVmctnhrIRH7WHrc5XetwODsPTSyVAL1G/zPD/SvW3kxnQWAPNUOQmtNtX5H3D8
qDlbjvJYa3dyo0OCVPxDgpbctmm76bwZnkKbNav3OSfFRBVCf6NTw00D2kq9LOmq
68/514OWN/kp5FAobzoa6D1uhjRrJs3rTYhS4ZAYJO0nMu0BvSOYURFv4kmTwTc+
oKgPci7MKi6KQAIVZBLWqLN3RIUW8bBTW9hEnBSVpG2dcHzl2KMbAIgbDpGLi2sT
WIhjSf2ZX3cGERxIxgWovA3mTVFLaBro+shwm8ebL11PQ8ZH3KqyJBmCU6c/iFaF
CnLofzyTMKABSlspbH2WHC0uJLDwTy1kfjiXA1O6t2GT+C/zcrqgfVWcHckTMrWj
1UUoHIxBTEgarX6Q4L6+iPtPjWof3AlHv09/QRgRWolVANb8QRSHwzcZgTqFtKF5
D5Kfms7LKJIK5x3JMfmg8Bttmaycphv9MOVObpTsj435QGHk1wg7xRyd55QY+jAS
gS7kAWbTT4sK/I2vEGiEDhyfDfeQizZptjwlJKJE9yapPHeqEXKZ970x/3Ly5Gjc
MyLqA6pIOfRKcCW9rCRhjALqgN/wvQlM/Vos/VvvpX/xPyAylHQNsQM3J/JhrweJ
2rb2+ULOvR92Wxb9SQRw7ZLd4mHzsO26hGv1zSh/RYLqwodyRXrskB2oczQMRXQ/
4lcRdFbzXksDTo+8N8GSFVPpcY0zo1wiC4eEXvoGQI1MqL254jxJwq48ZTHEnQmt
GVQxVWhY1e3FrePMAx2ddZOhX3HvGNATa6Wyh/+n8UdRBOF5nuL4jAfIfo7IN2vS
WnWlXf7OgWTu6Fudz64LDWEBdQb6yMMzJ/jDFU735n8g/y5BXrX/ddrjT0/T1F5w
ZpJPDkMFq74F2MZ+ai+D6pMoYE6r7VZHnsHTSqKhpNruZeiE+uCOe/yPQ576f3oZ
qyZATpZTFoTH1L/sQ1SfwFUEyHpUT1Om6gO73J3xSP6F8W3XebFE7UjX9cRl4R+J
73/rnDiko+vN88XocqRMA9d738fhW+IWeIm1tfF6bvDgSF/QfShPeQXS6yArYiMn
r416y6zRrJpvtzPY8YhPH9ugbsVSMKCGqrK3+XXaoX1ysN42+lF1LPHAJL8JrGeS
0y8haRgyIpUi+PxGuNlO3+3vHt0p4lni7ng6Dse6Tubfu6KkS/2NmsNFoRpj1jyP
ED+m0kG0WrW+Z+n5VkZtDpnkWG9ruEfey99TosHm7Q3a+VsrgSxzro3CQrgXC7Ba
wek4myQea4+KQ78KixjAdQTxbyaE+EOvBAgWS89D4wJfBNfWprl+SXjrK5Zuzbmj
nCxp5nWiT76d14nB4bvco24puN9UBc6u0XeugdtNOBSa+sDSkLJnZUbL9rYwi42H
yzEbvH8ZJwSZMB9RynTqjXVuY4VHVKktdZYBUjBVgvVLWVjaQVWkH07U5eH43jQI
65Ab8Ye7vzUYE/9UxQKQ4pP8NN9u01KIHIoBA3piR/alTv0MQ7YmLmmjlq4/PHPO
2OGjWiZqehwA5wq17O2P1eeTfDPiP6cEpnEoO6l4sCQVYezaEEsgGeO8XMIX0G8l
UZ604BU+a2qh9WN7/B/zG1qK8M9l0ixT7+MGtun7IgRkohMBB+04NCrb1BcI1UNn
UWgJOiutMP/YmARCqONP2Gv/Iz4oOV0FQ3vYjLd6V0pzfqWbjL1gW/B7p/VHnfEf
0s/0TeXoyCkiGA9PJyXPxATpVsdM+0LP0M/rmEx68zToXAdTetAeiWF8daEvU6kV
Qml6Hw9m8B6KcZeyExO4b2aC/R7CZTc3O5XV/HHMHM3v1+Adcvzlc0uTpsmufaer
WFbZHqSJl0z4rY4/HDfvP2jPa58DzYzSJ+ZDYU3s+IYY8TifGkFxMO7+Mn8efri/
fzRXTp0YCJa+ylpyssoKANtVYnR+tCPf1jYNPMrTkPcUPm9WRN2vPFI/5PmHkgcA
PimWuq+q7hfWWPJfwM0yz5udkwwKgUKmpfv6bwWgTu3B3BiYmO3qGqV47IoPeDB6
/h/FGTA19+AIOuzBsoeZNzm4Nt14aF0jeU8QP+NIcKY6qe7kXZzFUDvEinQ5iiV2
rYKo+qAzZLK62lwGcp4V7c4eGxwU7Wdov4bq1/cZV0iDDmkQfULFzJNduJuTAnnh
1AWQhnoUdAOpFg8cCLUVKlV1be5TjDFS+p8WcU6XowwdghJ267LrwhQKDSqib89t
Rbrn2jCl9JPOcacSv5duBXe1/ISZxXyeS+sn766wjld3KaFRlDVPn54tcimu2Bn4
sVRbjvppDgW5IxZCD+RNDi8AN50/opTfgy1qF9jc20YbHzCNlnOSnoNCc+xL/HYn
mIfddXBP6Zpr4BqAPB+UqspqfUUui3t9ews3M9jLY8BbPXkcgXgGy1Rki/9xya4x
vu/lQ1vkE1VFutQeXqiy6baRaFiB9V8DnC+nhAuuXK76lhvp0OeNX1VFVQvqqLg/
m/RZeWQgDsXOziPyx5LEKs820bwLbiypFR8T8w3VrPJDi0ewxwVCzMExL4ipxYzF
J5uAOtQSAjVSWbgiBlXaz2S8hyi5SDm8KTzNJE8cKwF3AKM95MPIXzsw+8jjxkkp
+YMLfAnMz/L6Ra3T2XGmaPWeyVER8yjRpY9nKVXP1HIVr3FeIrv0PuujRNsOF4Ok
74Het3JiK90/PWUQiBUkvS9XdF9j6fwXv6DvPcouSP+6N1eXa7cFdoWstOae2Xut
18lBtCfTzL1gqlm3et5aA2c7MWcFIhmI+jXQCcQa+VFio+9Ob1rrPWojHLpT4Q8D
qEbo50eyK1mF1CvF5s+diHloygYn4ziVJ+MiwPnRCedSap7jKEVxl5DqRJRbng6v
NjC/KFCjFhQ/XoiRZ2fGDN/WNNJCdZywzZ9IhPMLgl7t1g2mwogZyzPytbgNH08i
0RFmUDH6Nmsh8pseGbn1Pa92Se4pz0lL6wI9DCdWmDDGOu5uOmN4t3ykWH4rdTmN
lJZ58KtdyPZSIY6vkeiB2/qzOu/7VNF9NbF1tOEg57k/91iQf9C6rTo+/Ws69NGE
+Gy1K5z3BFj+tN39JuRHJMCiATrcTUSO6kLV0cvgGNfSQ8Jpq7OhVYo4i7868Voe
Ol3K6Xlssv9OlICK934MlaP53cMUuR4j1iOiDMx4tfRpzToclPsS2xZivKB+DMRE
Ix57B/e+FsUZUMIWvkRPS9GjFJns+I2tJgt6G04D8Csc0MdZV7yi9RXdjNEda1F/
51RsO9OpsAx90Nx59dBDPuG7TnVJ62jSeVTQmvkhbi8cLDcpTR0XwvwnEYIL43i2
iSGFLa2Kgedm420V2A9PFWf1ktHJ9DeuFk4vHF45qjA300BC/VZfdJXvgyzV7Ins
I3u/AhuFnxW1YY6Uk++U33uw0ypspuHOfxX5XxC61jmD1IGcwM7kDTU9jgxYtiBg
mXFUSPlJaKbgsQmRKCmuaHLpTBnaV6PhcTajipyrxdisaKI7hNsjnS+1UMRwgYFD
vWKrqAS4fj5foo8/1Epf1iRbXkupI9bbfzcFetZAHJ4ZNh0IQ9Bu6I+LnZzTeYDq
fWCGlzyQzHCCFQnU7hMivzdWEqfnyX7gYAsHfUQIHUpqWB27Bxt1ofo3y+RlVJ1R
rR/hhtbUGelbZuqZ2Jmgre8BTB6mFQrsRmpc2YmJA4O4mpyyg1dJ0X9QzwW9Z0/O
LZZPn0pwHJzc+2rwcmrzAO+LENI3vTbl5GJvQ7TGagIWuVuyRlgalwVbU+5ijrl3
yMvCgGCz51rSrq/dMbTkSn/7Ype+A9KXidqgRQJqurwGVGgyprHs7fstt75EkDbQ
POMiJPJw/hYVEPcKxwFN6ylSLQNyjWJQdO1u2a/T5Jr2p17/1wcYd7OcilDDIgbH
s2e6i6COMUQLVoK/eVIeOeKLHX6JdC6snxPcE9fIkHHZVYPzQsT724Wpchp+AaDT
k84Ox27frJ6I4dFVxN6l9szjEIKDLaWavd83yirexQT3SXCQZXSgsZFoKCTwUNqf
KKNcad6GrZdnE/LHHQ2lfM+kFAOb2L9WWffuWXnQZ4PmOdY8QUREoRp4uY/oN1DX
7c6zUh2awKHqOoCpMy1WeKLGAq5SaxuDCuhYHqfTiU8ZHAVA+1kykQRVebdar3yI
SgMVRY7IUShzq2tNGLoGCSVJofG81JGzb/3Os5fdhojUyuqX8pHG57I2cOodGygC
SQ/0mA4lx9WXWTj+WYQnCMltZq7kWyQFNwaizR6ViBdAKY1AJGxNi6rcSrKK6VQN
9C2r4DSwJ9DvRD/CPmDXlhXhaW0PuR4Kkdk70cdxkQuollyewCt0edR+/ShMsSFz
dCzDy7C7+JQG9JuY819aPW+ItjgIW/0Y7eH3r65oOWN2rPVPr0eeZn38Jqcm1ELN
wUntZXkTZbMjkc42t/dmq0LidsW93XXPj8IOxj0SclScnm+Zs2fXIuFUBWI5tZhw
fABVrWAKgnoC5+MGCNabqoWbq8aWGqwA64srTA0/dCTu3tg1+PZNrcEXy/kQoeXN
ayB7vZJk+eyrP+wE0vdRPu2WZL9iaEQ9tHR9FM+HgD98AWmjvsXeGDvzQ6M3/cg7
14F+RXSGBYg0HKUedt5EOoIPkX2miQKhEpSmU7e2l8FEGkhBGM7957i4bCgOD+Lp
XKriIMn1nqqE9y62SIKWG3XgG8bT7GWzwJB6gt5EyQ005e7ICszm7dHNOPCDu+Ma
0EZwB8rt4RNV0fHAjbLKafTwMdll9xqRWheDI7CIfHUxtAwtzDKFpZtni/+JdZhd
+ZLLln/0XDJPAubV4nGAn8a2qbT3AIVfkaFmaOgC5f6TfmHNqbJtvAsMr/d0Ad8C
FOq1i6d8Gz6K3G2k2d73vtms7PgKSVWzK859cZ445uyAObNDZtbl2/zMsRNKUauu
3bJSRNmoo6zRzwQKXUuOhSAZCaEYJAbuObNufsDFnFUBage9u3bWvpSVzrHqyka/
LELNIX2vXxWY9/UB9nfjM6BF2PRXQCVTuWJoSlcIuEq2rW6FWgL/xJgUxJ+WRNyD
i4I5muYht1sOm5zP7CBqFWMErmjYQzdSqnZXx6HDCz4dCD8tmCd8ql0xk/vCWNV5
JZh3QM+uUc7TQDyBI+QULtI1/hyRr+W7l9jO5pe+sqqrDRAMbZ/gRZ97agc+8Qty
MgzEogha8YBNuyxzy/KSzuDkGxxcs2fFkWLwriA1bXjJsoI1cLIHOf2gpZTla1/U
BFsE7A7zfHwpZzJPBEMho/Nvj6HvJB7UGw+YRMlfJf9XzU4+nflUWXroIsX4UCja
Gg+Imu07txGN/4kgIafRB5AdvATDVjDyT58ZnOu1+418SBMFbfxY9F4x6IuwouSO
byPJ1oqUr1cMoJhBbCFCQjVQJ/6IYMX006CKD+UWmDuBaSmv17x9Pf7iqPP65hdQ
8YFV7DgxyfRt9kIUWJwAnFHWxUjCnXuBD89gVtG83NUPqZgerPGC4tXivsqcSEK5
8fNg6MtFiOphrGahzfutw77nWylWN9MDROE829JdSaHgjxo+eyZcN9qDNY1St2cu
w7Z8U/j+O7BLJ2S/KkPjKnyWzpdNRR8tGWTAX71BymkmU3zWL/9weY8N2mrc7GBb
OV8dvUydivpPjbsCs5ukFjpEqndBMdESCaQ6il4Jvj3nYYWXTqElczPDsa7BKl2x
UY0cRMcrJxzS1iv81bX4rbtAJvRcAavhofkZoY7+lMV/eU+1S6c4vJ01lBnb8LUB
oFWQ7hs+sU86GPVU+4HnSIZZo5cl6rZv006nE6qYsKX6rTC1gb7Y3KQJkq3aPm48
bs1z6nHggpj7cpsL1Uo3fp3+T7ljCLuroOGt1su9i7JfJndNG5B4DVvGedwU9BiJ
PEs4et1dP5mbfbMXepNOY5KLbnqFLXWMU50/8mmhA78/6Vlyt40cCKHWL81/DUge
okDWe5L9leP80ocOTeDrLOnCq9LqQHnbePBdEl9Rdvd2RKu7/JP5tO4GFvqgYeaT
yIWclvBE5JqfWzLw4nVJcd5vtVMLL1ka0J4RMO0ssssVO9YL2KyuF1LkQ+D0uC2C
RIi1OtnNV8QYOPiTG1a39/C8gxYxgEpJOOEq0LRzuOumkEXCPcoeaXkZWZg1qFnM
Is0psCsLvJzlq6/e6M7asoXscC/Aql4JVDpG6Va8020EF36dOKNAe1/dcWelXgyQ
mHn8GBfUZ/y+54QvrFRU3LdYw0ZHRTl6uUENESgjxzAA4/KR7aTlqfMAyLFDjG0m
WdcOXnEdzdT7aKwbplCL6XtIXbdNRfRBF505aCtzGgyAcvut2sVRhK1+QtRyjH4B
0ir4BpgAJ/byZKTBHFB1c3bJWiVHUn/a5QJiQ35r6t2tMO6Av2KvUPOWRXd744hk
XVxyotxBsC8NDfAYPzMyRXsnR15Cek6BVPC/n+AtKHCIEzjn8Odd1e433dsSDNUK
qkG70D0iRW2WRobR5LI+eZnE9gXBsGq2g2U/hWH/uYS+C8L/U07tKaNrrQjMUyNC
Gqji2ubOl6VS/mQjEK26sdVyg1/JEKSTy+DD6lAtj6UQObd85UbrfSrow4o6hldW
Ecjt3h2uM7/74Dr327VbNimuePrM0T2c3POVIay3Rj52GSQroQEzh7X1TyrcrD0T
9rinEk3+rQ5RnlO3YR0pVAm2w+fbR2cnWnc0zYE/KezYDcQKNAKjMhncHO7Qyusf
qLKmjqhqPaXa97W59QtRd3Fh1f/M1eTaTOIcaI/g18isrj5jvi95QxXgqaR56bMJ
JGwJ4qeV0IxUZI4Dytd2nspNXot9XsF0SwCV1V3SA5OWGaVvefL2m2W4x3G5AfsZ
ZJ4qDv1Yb+rqdCtH+u6UlSF4gvyDmQNIMFNdeM/lxWOdTsVqFZHtre9UHkrgYf+W
kNXDwoMM0sVDx+V5NqzfIpcFa6ueRp+J2SBMQ99GdQfrcq/KE0o9mUJmTtWKUnBo
6/Nl8+jC+hRPpeOkp9gx5Y20wgslx7Jn7TjaPPSyD5TADBvIwatld5wQL5QJsNbN
dlRVQ2+p16LMnG66pIH4VkY3UNZ4lC85XlI8REuRTMR47UzXIyhx/oFJTWl7EQ6M
ChFB6Om5Gg6RVRT4HssFjht2jHnXC0soJtd2/Hr4zY65MHQ7cbrWFMIwchS/vgIo
+0gPNpgKWzsDcZUjfSQ7w+xmj12mDNHpxiEfig+zMq4Zrk7RlNHippKElqTzccGB
Ud6cRqORqCqr5DlW5s1KlgQrp7M3LAiQQQM7L8VFvcUo4l97u8t2CjjEM3P6Ro1r
AhWazMwcvpzLDzDcco+hTv2T1KD6rD4Mc+uK/KavDSVMzQOdX9zOr7empwZaVqNR
dM9plC/1rC+G/rl3rDoHmDryoaT/JYv3djkQ9a0GZ2S0utSVhu2Z/XAFWIOmx/al
RB6iRLlxvx5pP4XPmzmCQtPLjZBtVnLfFUD+7xjme33YB2gDtUowZ+f63o4iqh9F
wXzbkErQ6BC8VZ+vaE0FIrGU+fWIYmvm1/Uv9+HvWmiwppqrLH351KIYIkVyA3pK
v5yd5SnKnt1CJ3mnabFTqtzdwxHQGMWJg5CVuE4Zi9Z+BKqV+tjb3wJfiPANgGSZ
J0sTuhtqd7d21mIO2y22ed4ykUAy1/TTnxkowUdSC9eL+xhYcKzopDD5FdMaNim/
IJ3OCBI3cc7TB6n8f7y8fSP/EWppfxgZ/W/TG6Dw2F0Y4+87bZJUaHjxo9bD/kx3
G+hA1POeYrTHubRc14EoE+Sfg2UNWRgjCGKPMBS3gmZRm/S+58TUsNrU+3HiXj2m
xiJfv0h12VGyGKJFL0rjzMbwC5CzmHL2KrHIw73MVRjkUdx8XWIxKLSo4jbMcwZf
r85cUaFvFvBtV3dnXYxBb/eiZdcEFAVF26ZQ9cNF9EJUXaP7vt3YqARjPxvg3I4N
38IalUeI74agZUPEKhRiRMrCgwoERJ1ot5s86IuMk2qDq7I7h78+nnwX3JjE05wS
jy3KSUC7tKdQGwYdx2cnY2pra5wegDjdGBVkcLa/Y1H+WqXVC5eZoO6x/U9DmyeP
wt+qgYhsKoLqMlh/2RENGozQMcl/G+/zfXiD2NFwXIf0ov547fI5Jjiu9LaBBF03
A+CGLwuomvkljSR4dJiz7mtns1cEexM+i026fLiwxCPtzSBrFMw+kHhSYthYdQp1
b3ERpNstdU4gNY84o5+RUs+o64aXrKEid4A8OECWdxvfl6ZDT/i1ZTsw4+ds5+g1
3s5jB0DKbud1K0r5AG+6AOACf7OEiH2xoSmn7KgqqYFhFAyfee84RtLThkZMJaCl
K3MZqKW94cBGVKyFZ+McHB9S3pqQIhbCArOiynNF5GwI/K/i6IM3kIgxU71/P+dk
jeuOMQucdF4Lx8UsPqiObBiHUSjvPuSdYETYsizim9cTiJoD70pK22IW6jaL1qRv
abXLg0UMu2xYPXLov6gIa7lywkXmc02IBTyqFpVlj+iN3/+QFdpdmYCAFFbR0WqJ
xGD1Imb/ytdEfkpGp+ihut2/x7oqmYURXOZjyHYQkBvOIcCAoTIxajHYXv9SDCI6
b/VflSapfuh3S5FCGefe59j35ZjYbdYBWARuGvkWtAcBjiieBTZlJlISIklzMigx
a2+EZNAHae0GkRoUzlYFXpvjiA52aAjEWVo++II65+3BsXNZ9KF6/xuqYKmKlhbf
H8X1xVw2uyPAIrC+xEXyzIH62XRkZsmXWF6+OhSSN5xnGXjLvrMnQbi/4slDu2XI
sYbK7ZwNJhT/bV38r1H8+vOEvXbLn4uvtq81se+xotP0HQWZerikv0FXzEXB4oY0
z+5taOCbagKietl1LHZOfCX/D7+fIai0R0fQGOKwC+jrJhTOOn/uYsHGHEbkoaiW
mcffXTt+jSQJyE9L6yt5suZF/zIGxsl9BRqdSkDPjTX4F04V5R7uj3idzbYEcXPR
i9xTNUyn24PVk7M2Vfuq8PDVNWHrPFvcK8jAJQkWyDheDnFD5c/W9XdvmzeYSZhL
LBcFaOAlFi9gh0+2TumF4SzV7DZ0gGD+pTbR+VdaKlrDncEiQspCO+T+umc8tdBR
QDyNcZXWkZGN/oo59Bc0FRiYJ6lrJUfxOSBcyvLF1wJg6Xc01in9bwBUbBRX/mg/
rDEjtn7IGv7mDjMsowMFNTQMHUuGpYp0N/0oF2xkP8SbOqpZH/S9QWVVrypVXsHo
EuP+Xr/uizja/a7jFfjngwES/z7dWxX4lVFKj2zxprBGZuab95xMUS6lJYv1hWcH
063Ep0Sxf/cWtIfTJcfFqtxOUZQw5bl0HOEKCRrvPAh2Wy50EEdSaHNrxOT/5bwM
hUH7BzRr2MjIpxzLbTmxszayASkj5ZfJxW8u5LURpnwTFlYfYlkiWm/NJ19Ucaub
ui4YAarVjK/Ytlg6As17TRAthSD2+U3Jxix/DKb7SMmZJQbNKcNRKZYu1U8RZDuk
DH7iuepDGDFquBoLlHY4O5gaB7/4vKNKg/FYDgAx2D+ReWeYxTskycCZUnuQrIru
DevAPtLhDZeUchugG49sXtghJtjXauoehLTL5mVjBLajAKdK2P5W8LYcvk/CQwS3
ojonP1Biq3wikbf5h3vwgwpkInCdP7SpTeZLJyX1TowdOtRTfJG+8/0TtVv1Ogo+
26lphQJ0hCw0kAjhyFtjphV4BFhcan32u1ygHmtrvTlGGtn/KYW8W/xUF4/pgc8a
t+0W8WUi+LNcqolEqAPCc0kDChVyLlUjxTFxyklXeUpkNATvKx4/96VT6zyU6Wc9
xdpD3zie+XF8Ms3xHcKFl43u80t/qF5pAbR1TEI9rpp7J+dOo6/MVhKNbUWuR2Sq
ZC80PGY4lFE5bY6K4v6Ju6tjRk6eVUjxixT07cNoozBCW1xOohbckn8J5LnCt2zo
OXRzI8DxWco1drmX0B9jUjVLgFPCG7rPE8ie71e6/8uMbAZpchzR5JXhHLJ95wI/
AVEsLvN9yi7zUn3nc08Urq4qHrTbRzLxAIHCqC6YCqo+368nACdODS4ckyfrLH1M
3lQ/vB/Kt//+x2OaMFwWQj/ZhfYR0pAyxf+EAvi2utkejzKYNjl6g2L42dXpMUD5
TuorO5XNKJfWjc1UJ3NJh8fyFl0iY7Fgy5JO2/IkVlHEo8aVqLys1g6bwzeSd6pJ
j0VGpZRd2yvPwrXhef6J06wn5nFj3N8OAikecPntiD5z0x/ax5Jr7YX7z+n1H0CZ
T22OGCTflpFNKxq3iyLNL2nNEWK1MSV0zXe1S2w9U0Mlc/y5W9P5+oEktUGPTQeS
FK85heQKf+gecPZN9xcquDMEmdYNzS6mExTtcOi4KeeiNH4hMVVrpaM+RFrGImgh
s85IfDqkYqqG7z4X7p5Btx6RSB6mPCaefp+PtX2roBczgrVfdDmK/kcyVRkmHOnK
662OzmSxp2H+zYwmlTLJAF7B4uZrEPpT7l4eSU1fLaLWMJsonyta4+/8srAT4HCo
kaseUlCXJ/1QifzWSot5kohN3SECGHgn5bJ+1rqyXvIvNbied/z014kw5HkEDxEN
IIJitIGqcUMBYSaaeC5C4pNfKuxgxs9fVSMe9hFhllGMXAmr/boDXFOr8FQBCK+Q
iPj0CIHsTqSW7WI6UqP2v9xNOODUyB5VXkcS142xrv6ttRd0IU9K+8QkunqDv1dR
fav69l4Mngi+7RaIrh5W3J1h5SSt+oH3/3zikdvxQ7Sp1qaymkYs8n+DF86Aet2I
5TsvWq+gxeUb6XgWvvRNtWqg5wpZTb6bq9noKsadgn9GMn2MHH3zrEOqhuF6UdeW
8B+LOcB5iYu0mfHuf1S61cLV5lYWniyWyHwZV+mX6KJti0wwvfGnDvB2yum7+s16
zoTdjsai2xAKSKadnlHy37/w0CVaWgEwI07XFCkqhPT20fnRQAdCmE700dwDO81K
J4awMDFOahgi58+GnfTQ+udR4UK3GNypQATsrXNjkWZMCuIjNk+KbW195gnxyVnZ
wGxWItQ9qHKMCb9zsgo8UeYxA0yA7ek7MTTUFG//h2CeXHBn6m5mCWr2rHGYDs3e
IyN+X0G1hX89iNOX0wC8pEnSEJLCvc0xHxwH4xRx42GWIZAaqCsnqk3l5z5HzBoL
xurnytHHBaOVvi9QqVDBUhq6HTIhmfe2m5q5GZfMnk61VHeih9aMk8svI/8iigIU
KaEygVCrg0S7q3xSEIKTkHlvGmOy9yKp3377WFb5Imgd7qRcL1iQJ0q6mialLSQG
dyeWu0BRicZrkfwM8RNOiEPyn3qEFv7jdN4br5xC6wHTB0jRBRYSZ4VzHGSaNHJC
bC4xzZn+fE0BJzb7mQH1jRTi3AVENaXt9bEAMmIpYhdZZNL95a89n6z2hiI04n+E
a2j4fcTOEV6vJjfAGeRYveUQwQIqwLmpKHHEtxcvHH1uztQYo5fSMgSIAoodP+nt
YmSobNNDtAUhFL4OXRNoBXe3TwlE4ckoWTKnvZ1NpIV9E9M2cBoYuDU1UUpyp+pR
JjMGvlKZnx5stQ9yvQ2SZmB/lEtNd5LZI6K318x8s2yOFj9avCQnjm315241NbF+
F0eoZvbt4BaMK575WyBqnlvZXxjSRpp4f96jDaohcPcMXbaItUTzPOJ8QaJOmtNY
F64jb2CpqspT7Ir1MluSVKWMVHuaFQpyk7U1LvRDL2XnXFHksuEaAw+gyRuKbbBJ
FdaalyHP0HyRiGDCUBhfM/x48AX/9ZuIJEOioCzzxvY8U9QxnPXpslqdvlzIffIw
36EbaaEv6qDQ8GF5cLwopN9sOmJzLCok/fnTO27WIhGvJTcx4han/XixsqBOEhZY
ymSmyiod8YrgVr+6uGoE5xVz89nGn0tkBdX7n+X08/VndQ2RPpmBxwgpR72pMl4Y
l0Jdz6ehtBfmpMmRGaVKjAmceu7+QlDKAbJj6U6QsbyGfe8d/RqEYFsvCEQ6vAwF
7NT8DiPfFL3IW3YI1il07giCa2RdHL6XIRVk3Wn6Vrgb7BqTfiNOIWbttdtkfv31
EjadpvTEuD5v2+84aBg1RreAayd4ibHYtg2uT7Qdwm40yOyQOdaWecThJWz66ObC
AZ5lIoePhjYPCRrBBB1p0p68aoaN6lj51p76LiO76W5feNN7vvOTNo09wldvN/WH
tHvD74r6Kfc/7R0WLJiEYJeBJrF9EoI/yRJa6h7gTescd4K/Ehrvr++BdXaswqML
BXcaLPYaSurakmxvx3ff5XArRwfORf8UwYi291SXhY0eZ2wQcWNBdMfV36NaH54I
dZL/gv/ZOWIPI8Bn6uZcxWubG8k0xsRRqwTCgBprwzlGX8r8KS0dVuULi2U8Qrij
2eht2O0pRSfqGrngTFH9+uejKA9dvR3lcKD2y0OPBh+dxjDauaA+MkQF8gBLJFgw
AUHSOoE4dBuXPDT2zInXpotWHlu5gNNCuD+FF6n3D6CdmGOO/VO8BNugE60Abkpd
VRUbs/F/UAB+QVfRx6NCMiYdLQ1p0/uDIH+A/r3w0Bb0aDpW1VWnfHqXmjqvSDNU
0g/48U8nGpTkpHpTUlcyAkwQuSmlFGavofY2UVIBjpaIhEyRDm3f0lfAEYflC5uL
avBYx8QkPFW83iUO/YEeTUvVAZM+JiJsK9tqtud2EuTH9JJbauzLPE9a1CscrKkA
LFPuMpx1HKaFg/bNA7923gm6FaTVhfENfwNjNNn/RwHME7RM3JUK3/A0aENbRSbP
UMtWGanQzd1aXz66zGjWVA8sOeQz5UOlIbNpfhNxRiZA2eA9E5zXkB8SjnwaXbWs
ZVofRfPcVKwoLn8rJJwX6/hjF5LXJmVD2O9HMa9vPnSEmQLbMErXN+XkzAOLqJ5l
+AZQd5q+S8lj1LGUEJEjNmEMcPCfeDVHA5b+I79DbfwX+bVXYpln6XMQwQnUCqd/
zQiS2bjOwq+68/g9ZHRtZLf3NNwU5AyV/2XK9IaxbxNqWu9rwP/VJ43jT5i1hNK0
CEyz9MXMPP4D02owQhoLQbdqQ+QFCAVNYkrwb0JYneN0hc9mVvrh+XLoCs47NuuQ
lfyWomUZD7/ekA/l5Af5P86lP/KtfzgGTSZvc2KVQLrjNFT4rDjTk/WrKZIcOVW5
h8BWf8+wu4y4F+jKZebXOjoDIPNbeHBaSHUMujp+IIKbXbRNpIeGS6QrP9du5eUg
dhPnwghlY0Xu4mWcemqwCU5Zx/TN3w4xV8SSiipL57edBeZx4XuPoKeArx4+MiPA
yKq2YVLR8yrWemGxwn2HEoUHgmtlOQ+xUcvI4RUyrU4FLqf402ZQi586AUMm94d/
pVj57S6/hbOOIYm0C7lRk32YIlp/Ys+2jq2BB+FcOEy1krJOeINc2r+McTJG8KzN
xE/t2es8MOZnqHIegX/vU2f5zvYZ2lJcSc6hCn07Vt/WbaSr15UqUJaS4UgI7J0M
LQoKc1fPQ53h8bbayd5aK/zKdh82Y15yMXEczJFdjCRhPkPU1zfxOPTC1aN/BgpT
CQ7x2Fo1XASp1YjqWVpvM+DwukzGt6sNBOJN18LeJMTuHKLvCAS9/0uyhDbG9wR+
UWeX5SEmeA/Y1MsP0+0CMHWQJUHAPskgKEf634L9pgOFJkjAt/wQZ5tlSebxEEAB
SNlokNjEIoRSKqtb0+Gp8QYyzehTNFxw5dGvx1NdlalVgD4lO6rOSvvmnQ4EdXDI
AAc8VakZ5K5doA5pVQRw0Hqa4nXj3MuJ45uWBQUBVrTvkBz1YfY3HetgGHDjRsRT
7ihOhuzIgYjkVkdcblF7JBuUzAS7+wsgVZTZ2fymuqgW2IbwnAfEE9ScFRfYz8xr
zFLFItq8q7UI7II1l0mfYQWPWiIwfQArRQclrqnE9VjWPjcMhll7+bKdXQmgEPvp
V3u5MCjJgfA7Y/SO2GXksGzEhHu5cVx4H1e0GUrtmzNYpmwvkF8+RF0JP82qph7q
3nZROuufv2rpkZokZbRix+cgMfBsqbuGbC8NF4lSUP356MP07/EyDRpbjX47Nb+8
0K2jPNAysNOaF7UCpjH8xv+KN5bFL27NKLcJBhPlPguqA42VX0bcT/6SO5BRzzYz
TTASU4ozBc5/NL1LkqJsilgoofH9pP2lFdwwa1M96LQGNaegPIsAhL/Cq3HWDsk/
PyTn7xBt5x2tS2+Nchy8K05cMzkDSR2PkK1bYaAsNzoX6YkAPU/BOivMVqJ4Gnx0
w3bQTt2xF6us6jnvVU/u9tBjt8U6uKh9fXIog+0CyQqzEbTxb6qOuridJv48El8M
9FMKUMBb7NBUA551aS5VOLOEaTUke+sLJgGQTov5WyzI/71pdLJWg19c2m7AMoRD
bnmtN5lJdZqq5mo1kM3dct2Zd9ujIYhzXTXCfYM3CUcI18GAbM/9XqraDqWuHq8d
xEmlwiiSxd1/WkOoNamV2uVZ+YQw1U0Do2ZKJhNXpGjTW7gETJ7AKpoICU/Yb7yW
n9Wkix1rugIMOMJJGIBYC4ZQ2zl77X6HzhFrpZcye3NdfC2NskSrh2wtGXyzSVPy
8l/0US5SyQiosPYkAhS1g4doTV5LcsY3l5N0mTZEu32ARMjTumwjLZ7/1sgh9BzF
QxwMAnbsRVNslZowRvS6GZbXwkf8QlD0MQRJfN9HcPK5GhgswVcWxEjJgjNXlFo1
+qABnf1Pa+/3xgWTsLe7eeeOZ81g1x2zSyqOv3twx8Kc6LatEnknVi23Y6EeTHNM
ls14/8ckHelIB4rLv9eaiHLA0j76xokYueIEzDRIZnxzps/CBVmt249trvY6/TBq
Oz4/r3LOptUcKWCJZAEaaHILiw+S/r9DvxRUYQkOEzOiQ8L48QsJTlj24IPC6fcq
voJme/jaaPOC3JUnK2da3ppVye4X9W6DOw/1EuvHS6n3ePgTH10qZp48IxDYQmmn
gM3XvGZnArQF9oevh6Usqzq6ru0rMXwsRSoF0/GBL3GlZ1XBOGdr6Kl8d8XuSQI8
9njAOSqjWWl/Tymt9BuKjVh/c8GpfMd6XgTDtx6XWjsSA8N7HJMATc+WOjqF+jwl
fcPWQEWsVRZCvoGmp4Xmesl0WcHa14s+vyrbQu2pk24Em2x2XMyknlJcJ/tCpAim
kutU0gt+iPsa+byr2LOKu64bGzHvPzEdUwiINKjTKNB47aH8acTGu0SR6AaXQPiD
AZNkEb4pdgptryiGJkpyuspIMgm+tNCry+oC79qzrLsvNKbOwP9nSJycTnHhijmR
BMG/zeNfdVKiN0uRDqxqFFI9iAty/NZU9t89O2ZO7v+bmShnnlqGsvQGuzQ4EyDd
kNC9S80erK3TFXa0L3ZPGASR09kWFJYyAkRp7Y7uHa/zzBXqNpAokQQQ5HJXi2zq
rXsY2FaWcUM/ygWxpLcvvluQjPBBk89iNtMSl9P9WGFI4iNiC/8DEiVS1nRcjDEv
B31LQO3jBC41kcayYRe0WEWkgiRQNNcY8twP6427vcYFdPjcSf+j77c2Zcegb8U4
f9MVweOuNRT/GtDqamTv+lIj2+eq17JqiS9aOTyMl5pZE7GNp+EbBAI+wT8BWjbo
S3izsGTowSUvfsdIbxrqOp0KhmTOtJjcm45FeT9svB241JLzooxJESDmJZOqgJzx
vhlJLWdmT480xHdDCMZgtKBzLByb7bD7C3uk3RvzER9vXkbdVB4rqwcJ4NPeE5MW
VbSaXq6IIWVm5Ob2rRkA9u7T0b9lCpS7QtMAq6Df//NpeW6H2xU4BZdJi5NdveEh
dRJxtL4HlZmx2GrEB3k3yWmb8TYFewsAH11YUDpRz0umA+se9gTnFSeNl2H12ifE
Ssbe17F/bxwu/Slix/exgf1okZd7WDFuLJggn+TN5kqoTAOZFQs4Ib06nR2974lY
35hS+eN+l6qliza9jzgSl+VA0FuXYEWidAIML0mYMOUXWkY7KBYd2crZocswXxvj
Sli+eK8EdDLW5N9/kLxmgv7rMnXljjl/8g94A5cSuCQhW0BOtMhjL1cnRF+MfNJ1
x9Ld+kJCla2Vf2eXv+UzB4YhodV4831t3AU2lwemvl5SAq5+pio6mQ3Tmxh+O3wg
re9RN+GUeIYAtCrQS2fVD4rWvjuS3t+UG4H1GO9Uod3Kmqp6SNahjGen3yeg/+QF
tb1lTHSuEo87gUx5wzvQeGB5omVrHRzuakmSUrFxBTDD4owt305SJwLq4dbqNigO
4GX3EojgdCU8VVOVY/U2jds972xaiNEtXYa8VbjvOSlbm9VYeaUG9HBoZqJhYr/h
WVeohKujPkww7Wf4+hbs4UvIsCT0L+7/R8DjCTFuatFKonVaKlEuJ6J9Nb68qYEJ
o6d8I+EOypx55riZQ/F5JFqmD4Xln179Z7s1GcOGsv6ahfBr7F9jysgR7uCwIeF6
qNlm5hik7p4rBWI47wSybuYXEnHCzg9fos4iHLscKIyh3OxE2nbY799HUElX2Mal
FqHMeQe3+z0mATt7Pq+m5UlrsWaA/jRGzyY04jcJ00kTv9KhFQUxHHyCnSxGLZrG
GbNfrKJ/1T3/DEeIX6gusZi9qa0khgkV+ctqBi4c84uX1Z4LI1bxfdnjmcozMuaH
L3nr9Jdx+bWL7dUAHL3y/ePZ9raiE1kCmgudfGwzrQ0HcqHrw2XGgGUk8rVcILdO
xf2mWsYnGEEagKF/1h2XswmsTAtbTd7uFoMlje+SIE7HH3cZc3IkdiK+MoH82Zm/
qTaq+phCR7ffdDOpT+CM4645+Mp9GnQZdTnDHXgVp4fbDA7lbui6y2uX0uV0aADJ
QN72ZF3hYfjNoaWW6aBW8OEi0iq39gU+wdKo8wQ8tMXhvSMbOWF3sqa/FyvhOwF7
CqQ2n6h6NlekepwvpRtgDlkcYj0aQFnoBmZQ4xLi7gOgwo0Q1PrlsKwjdU7LU8+3
8UpkLq+0QX8fWN7LPGSi0s9GNbe1bt13TVoDrJ0IxC2xLvfT919JmxFHdfT1yFAk
2KkSn0JGLwBspq+vhoe6lp7Z22+4T8X1JfpkacDc9FtfJWLT+QaPkLOO6dnVSsZI
zK8Lt6CavSQul0eycALZyXhFZ89QIIZx8le2L4w3zVhJH5kd1OMFJ/LwTkxCqxON
RyS4k3qy4SxY1obuTKTIK96xsAxHOFi70QuVSYDWe7PyWnL7NXLZQzSByigRHoNF
ZE+fa8gNvVbajbDWI+kR5QogmZqoaMlWxK/WOFpDxas2etheJgzuVsTzdvlch3Jq
hx8nyY4GObrKC3KFVoGqCnaQAdqAZ4Pv9lq8F+MTd2u1g+j/OHi45X4+1NaGJeHP
cYIMVq5QYIp7nBR7co4S6cf9/8unvbI8YsG5Hn2gikbLmkKRFWQVKVfJcc1IC0J/
uoBB4kUuGROi6Aj3Db6BsYc8eAiHGvMO9f52mQgklbaxdEQuLPduPpw+W0M3LR9J
K1rFkv45jJcMBiM/aombUBPmcxVhNksyey/nt9a6z/PPqZ+o1k7lNLDy/Ly9U2NO
dGUcluVL231lpUTz7y1yGmmg+lyzoSlqejohxADihd6L9T7EfHjDKPXRHD+S0Y8S
ffupptivIxVR/JO67N/6tFTtGP6jIYgjWMCgaRZh8i3pqJSS1z29ZP2KPuWYcceN
o/mp2TmOVBiYRzTFsI1CMRzrWVeizzMKXjH5hyFoZi1R8IqYosj+c4Ydb8O0dDnb
GO/61vJlUlLC76gM86Xa9YX+iDW7c2gyPn+6jwSuCTPCdIT35P6cIcG/wX+Qak0c
uYK/60zydA9dyNTpXTSRQXVpPztaA9S8dWvfdYNORgrFJpIyTBxQGx7j3G6h5SZL
L36UoMgJOJepCIyHrg3PChp17t5qgu93ubyYkD3T8Rmx48EBiOmd8HW/MmzS0WED
njDoABKRvPiCCnykRjjxLjz5DHIEu1xBjBH9Wz8bh8V9vA3hxIxxy2TftX/jIMhA
MAs68tGgqnCqIihlj3T1udK2K74XHCahg1We0rmSRemn/gd1WL1gvDOFFuPSE6kx
QdlEZAoAKxe5FnGl+ApQ8NiGr8JlMWD3XzumjUNIdZQD0xwl4o6DgMvPWiVBEj8Q
LVursfpWFydc42rFIGRPKoWIizy1o1sFbq8Z1LdtsWc0LwlcHMk9TuQFGAnDOY/Q
7Dpq4zwOvrJdZsdWf2PWR/0+2zNFDHRsHh4AB0BIEGQd7nv2/VD11C+HAyhGnI6a
NGWxh2epQkjARYIi7JwC7kJ5MYLRxV3BfeMj6k5L16bJR9cPDVTGH3DK+PXsFkg5
mIMlIUiMzxSQg9OMORlGAwvZ/GNEcw8a774Bb8qJjRFS7ZTivmRggavZRHRUl2UG
KXdvHWMB5O7uxM5AlZ6Kzi7z0OU7kPzGYR0FKN2LbXX9LcdcJVrZnAHkTdBhn3Jn
BFRL3M+gP5FauWNV0EeizG4N0rDWEWc3SJKdS5VvY+1kNLpnURlX4sGJTs2cF+75
vkStcnnxQE4p/A8LHayvnYEgqp4C9rQ2xweS849hskhziPOkDYUjyCwIB6W7fL/C
7H+TKhBnaOQAymeAI1s3YgkuB2gyIjqYTRAVPyRfVs4oY+2hQamm5ZaOxVzk6Atj
XFG6kxkiQ38bQi3gXopvwHmb9mOihc2OxViL+bbT+iVFLppT11DQG+vrfMNM+uSp
dWo+NwVUKo5pqtvSa5KIcdM+MTn6ORO7XmrxVuXYWtHPiAg4/74lbf3MmHVcgXhe
h0iERmFxRuinb4NLU5qqIcyB73m3M5NLo3U/pTCpUfs7H7V+KAnQiL9y8B5wuX3U
yX6YspB8/YvQOcp7SyHRfe5xdtFUy+AgjR39eGCNIL8pWYL/MbbvfZ52ZVXP2ZEd
GDHC8x4s0/9qDJCJ3jHwLT8qK3ZZWP2nZoOrs58pemE7aka47pPBqHq/LdlrnfCG
T7JjKCrnhS709UjDZjYq/X/q/akRyJ1FoPu/xeUn87H8jydXaWlFaQqqvKlCDRw9
6jDI5g33lbRXGOWwYGoi6LHBBi73AEeh95hoMhvqLKTvU0LggmOqFy51pELd9ldc
givCU1zZUJZeZgOw5Lt6CDhRQWKTE7nc3xqArdVAX+oQ8TIGd+CAVl42wyrT3++f
16fBos6+7Eiqva/2PUXH78faOubwLJIBhMFzfOFfOC8aCwl57jIVV9VfDt1XSBv9
nruO3uAvzwMfGLmI1WoMYPkcpb3W9towvJ2TddV55EOw8gwitZYNhJNR7fLyLP4X
/ucJj8WKkSqdo9EeXiGae3mLy02AqWhT0zGqEu4zVhxfP0QNoRe/C0mRhfBEVea6
XafK7Y/8buv761ao5cmXPPm/9lpaTRzYz8tuUFf4bfEW75D1NDGsDhLyhn++gm+Q
DrsygB+JojprJGkxGJbnyHrNFMIcA7U0cL66sh9TdRWaOBEkZKpTU1X4I0+J/kV+
YZJB+j1iWDyWtDuJjlnQCLSUnBN0sEt59xNHtDu/EQZuDPOjGlhRn6bIbmm1ULuT
vgulsjSgEJHcK2GDi0EAcBv9KT0wrNOP6cPOTYXF+c72zKnt3YfoOtQ9OlDs2hIB
MP8lsQQq10XeRaYBtgo6WOrWcUpu199Fk+HEElkSY+dwwI8Z8IweUDyFK/RzQ6RZ
+Pd1h8vBnmOiUsQnf31Dcs7GYyxFflactBchQPT3VmzYTX60qupo6yggg7aT8FQU
WqNx9djN4IDRmaCWjkuLDs/YuYEmRqvLKCB4reQTIjlU8iMYvLEz3DrpA5QPkc0B
rYCp/9FSG8km/CYTyym6oM0E/YRbSJQ+U0Pr5fhDOb2ths0IUYydnL75caTCQb4L
MBioYJi1B89DRpcqKp0HY2ZqwkdoCSUpHAOK+UPiCqwQI0V8xDhEbu5JUmP0d/Hg
81CVLexhx5cX4y6E3QAsbAt+Ykb8txhVa2/dMsmw/s3DXJtjy5R4GzMufIekacc2
3cASKk71CcxGE6KMOrF0sQ8uebfaIbNy7fSMEnT20X0FH+gll2Ao+SggcTJFRu+Y
gEh6RQ81CdkpGe8JfqUGnHl45K6xX2MOvUd4ZYIbO6FVBIoph6Zx7fADzElWlL+D
hBbNHgGaS3zoYxWMN9x5vw6AYkSgSmraB+EYGGG5MaqZ6x8kdWUKucD8jByUnHIy
/OJq4TulYjwiHcw+pESw81V/REUFdidNiWYJtfdjw0sxKddJDJOJkEcK4+XgbM7p
6eswbQTfNFD9/9Q+ndzBXbXgEcyeYjvRGyabZ7OorCxIDmoj2td/Bf+8I2XFvRSw
4ukZhgrnTJaKhIhRVQCel5ZN8Fg4HpfvW4EcFrgAv6H1c0IUPUtAWusB/C8NOLKM
sSOWJ7g0wlYviTrEoxMypNnpYy2Dp/40ezH4rg+FV45l0GeE19JKh7NgZBRxR2Pi
ZpRpsxbOGHCXjsXxMqzQt5pp3y0pbElJ4tJU9y09L/ot3CBWYJ9xW9b7UU3yUn70
3VmoFs09+tX7Sr5cNHbWX85Z8ucXK3sgZBKgv82vYnFgn6n0YYIOYoGRrLoLL5oQ
Q2yTS8UFvjsVpIWJ8U1Cqr/SNEYBRYFFuHO5ECPya3XiclJ9nqwyxs1OBJsE3cSA
MXiogapMmu6mljFTCT4La8ksz3J9/vV7Uf6XqJx/A8jbWDwokaHh9JCDl19+kPkh
04oXWQALyEeAX9h8nH/+Y4lkvQXA8Jt06vZvaqtvomJt+rlT8c+pYcVqkUHiP/lp
eWPqmBPcyhre4Qe/4oo2CVex3nobLIJb1HD90qjaON8Bl/LW3rcS6Ngymk5U9/al
eC2Sd673NHON3gSLFqFlgTgFvkQUs0wyNzXQfmYpNsz2w06EFV3aw3iStHB8mUHk
LWiR83a4UyTJBiNAOfhK3ajbgYNg52svQBE1fcXbyR0j455KtnzaXJg1n/9EJUxV
wQHdYEGTGCnjWYnQb0bezM6e1dKJMYZ1O7cFeqvvip+WZBAx2vpquU5uZTSrYIyg
HO90i6gatfLYGuan2JLEhu76JG76DTqgAfU3wU5YSQ7RR94Eo284Uj6aKF72L8dM
1BFphMvdeLuX5RiXYWGoDUJqFtaqHvIQr+SGDkChLUASoqlTbNc1/Gxuh1Qwmdus
osQPmH/p8QVgw6ws4cNXoeJUaQkpvzGOdLVKSV3Gg9sbOa3gPgvineMqFAnNsJ21
K5FdEVc0R2fX4PXpA6iQaF2Fwi17s7g9lMGeuctv4og8G17kcl76PKyn3Mc09Iw4
g22oWZq2F2D0ZOMYM0UeV5/RCUtL+T3cgED+UScH499bRuXazEfd9GjcaKIws9oI
X8L99KHEAwfrFzFVJZOs0cSfyMLx2RMYgk4qizpPcAgMLwDGRuQGJN4jVlOjxKaf
WwcZ7upUOrYRsgfUhW8Xg5Zf7iUL4bdxmnwBrhO4H+17OEUe/nzxHPjdjFQNNIYY
qFwEMcULhH3aHysXhpzjCKVxrBhVrw7H3VBg43fdaWTnFk9Sch+hnSjLd6NsX03W
Z1Jga1Znm8mWTkOT/aeRViyKY/QAtwsYkXCqASF30/qkSMzqsGLOZqcBKaeeRJhN
N6X18TZA2agld6NL/THf4SqXBu23HsOUfur3BG2bDTSCMqapOHQPx6w9SW3GWrmi
PbZ9u+NlqE37H+H9sow/qcK8Gu7lLVKs54q6+K6vjBrgjHArh14lfZPnAj+IVm8h
d2xy31ZlX1K14Z99V6kHzEpySQmwFu1mAismPc7rrOnyUk5hUzIn0SNz8+PpBGrD
BYKuq9oVzYc45DOBBSOOIe2uQeDvyx53rgyX/b5KjOaMllvlRI7cSS3D83HQjCXm
h/CZNnL3m0ALbDWLE+aA6zXdVKOgUVI8ORf2QrFZsiiPRSowI6arAVFISdMmy0k+
hIb3Jk/8SFMomwMi6IQ8NYrCZWdEhQuymhJ24jqtwfUflFzdqDwU6b/Wi2myPZnS
Qh5n8muLnyeEbY4rqvYPFQK2hD5jxbXQ/rI1OTLJ2T4Bw8I2h+S+18lkyVfckUCy
EekULKfIQEfmh4BZ9lf5MJJY2Vs0HR3eRrw2v1HAnIdxh9gO213Cmf5Uuefd5COH
5SsJK/mySwEqqcNwvLuNHoeP/659GdrxOO3ZA2oZ2XB3I7Ky16N+fewLEsKlwbR2
REEPX+C8UMEh31y8XXVmdDTZwgt2/Ck3UUQyRFISXzL63DTUhIJHi3ApZyE1pyWZ
l4Zo3T4Xw0snGJWT6bXEZ+R8B1clFJbgSh1UXJ4aFkB0B+HRqmYnQ/WsmH6kSfM0
M5kO90DD1IaUi6aiM9AdX17SLTcqz77wXXYQVpwm2rQyhzSxZwDpQg2nuIF7vAGj
UypDYGul1z2NH0dhW5az5Enk0nys6dSn1I6G3ht2jyFxHHUV6C9DVwKr7vPSOqAC
181lCC4wgcQY49qoQDovfCqSsbdTVlUyuCJDLXonMYG65+S5Z1/sRpdQnmm2TIVO
PrbufQt+84UypDvrH6BCln0OPpahn0msFkm2S8DDC4iV6HwyUvo5jSNH/G0n+U/d
Mshhr44wHCtzS2iWsdht/fupTAqBXiAdkZAvHu+YLnoFD2pqKeNptx1XKJwI0NQh
q358vvc8IcbW14eO3SEUKRB8qsMKWi9NAcXchyWLP7tpEkIhZx1G5qEovU8befGo
XjoiEaIJl74FmmOrVhB1Ggky81B1QLAcZnpuYOXKvolWYXthxZBP1RVuKVnOKpEM
pH8SlESCEiVG3U9mOYls72JJ6dC1QY43AZ25R2sqba5w//UmwCVjIPwsYc6+kguT
v9m7DCw01HUhlEPPN31Qsisg7ygbHNZKQeM8v6NcBIYfCFbC/8pKqYZ0bbdoEVXU
W7JaKsklfrD8+00TYwdjGaf+vVjgEralsQbg0SRtUO8L29t3BiUpEkdW+ClwzxA2
I3ILdU3o1/Cm44UX2WwCEwbiZJTCb72BvYjap844GAWdIHP4woThctcU5EPek13y
oGkHWKfVqoG980k+/LmhY38p9BesrCL+RhvJCHPZBYYQzv0X+EQY4GFUNF3mARqM
YYP61OOZBQ3LCbvaZodQkZcy9z7uOY8qVZ83OhJFP4m+/0xYhtVE+LG9+c+Hj6fG
Xy8chdNBSzBhCf1of6opvbe6QD1Wekr407OSyHxpjtkqcm06f/BYPQuWR0B4pMpw
DZGGCOmDGXJmzBWDub5Ox6SudlZFRj6I/vbXHV0tgSS7T7fDdXAWIMyOJ5JlZeP/
B21tl56zfsuQPslM8XItC4xwMkh7yFyQQ3dKXMARs/Zwe/ld0geMXJLw7g3nXG1r
fuqa58ufhX+6B/NzmA8Dz11wGKviXQR7wJqWpZ+5VKFH2j/mlBvORoQSTCQHITou
bIlvxjjMZ6tiH/qAw+P7XZPmyEYP6XEGcE/0C8Fzcdd7Lz5Uj6ZScQkydfcUhz4F
M2q87LjUZO0VwiQDiVf1JRd7bHLV7I0O8vGTJA8EtJhEPYFnu9XgKIhdOVnp4hoT
/FTeeMVjuz+rHGZvNZxwulk14YkmyvjzQjs15d308tAwEwqEixxK7nsIpglfX7eu
krAmsGy3Hv27J8fWPRZu271ZquSknqxZ8UYFNuikIbhgEbi+5/whAVmDFwAJXqfw
8oLTcEX1q3agdBvLCTzHorvhbSKMYOJzPzj/7PyPk5eHHltQEpAx3JMnHyCtR32/
YAHVd59VxUJ5u1n7KJUNFNjqQk9vSHj424sqfIc+qmfqiylVNLhR+FbvzeSdSvFO
uol/bczx78gaxy5Vt++FGjBzYaeuidE2+hKfpc6jD7d1KtTbwaFZKhr1EPWp7GaL
MSBrbNFGP6ogyJ44Nfe+RAyQigdpggrYaVRHRiZ/MAmeWk8MhPU3iB1eh9CYctKt
XMgijmq5ckaSgTTjLE99Brh7mhbPGrMdDc01Pp8w/PRO2o+oq+8Usp8D0PZ2clKI
ue4rady3I6gtf3cFW9fhx2VZMC1oMhMGvLAkneokeJ1FSYXDpI+O6l8LB+kkHH/8
e8cH5TQgx0i6OTZ7UtQHgm/SPS9/POLRiT7UlCggmdqZchllCdi6gPsud2euXhRu
LsKJF+zvH+CQU5LXxkpJDeMY5WGcfyKvzyv5END/y/aYPbN9QPfSM5yloTiFPxWW
zJEYqERwGLMBX7mdtBODf0Bj+Fb8Ln7eVq9dFDiM1BWzsL8HfMFAB5ki9EsPThpb
ByBniJrroBX4FWO5fOsQGGYOcbFlMhuTCaQ+KYLhNm/jGrRUkfKWU79oDMcZINoE
YoUPPY1txxdYR3pJ0VcdrHVtyEumh+/NRL15lZxp52wPPjXtqH20NkQ0TB/2o3Wd
jmfhcgjETTsyJVLpXWgqL+tEcDQMONmCJDuzrN923P+rrxvH9Tz3XUiPCM9FSMqV
Bdxpn0r/nJQWrtVMO5RT/8DY1xSCxOURGmAegtlmvWTxxSO1kiU+k7GYamoUgBIz
1JO1Ad54UPPoRJ1Dn8vzvwPrIrWc86cZ2Vny4gm1Qub0zVy8eHhzNfoGNmoocZzE
u3FR8w0KMSKttGAegjTtERtEZ2gCePWgIRTkOyc6vmyZZkEs27y+mfCfw4crP+7A
Yi5yHpqw61rAN/uNbhr8LUOiP7JSsP5shQ1KwsoDBvSvzKcWsWE8Nc9ACvvAUPE6
yANPdcTwVnFtaXxbzgM0mN5C6RtDCykYbo9o5AZqyRL8NPhzi1JXAqz3BA9Rcfzb
2VmtmBppNf8O49YY3+AHDBdXsUCMtrvqLBPDZrd+YG5Tv0MMTPPPWBgs26ZTs8wa
4KxcqV+8+Y776QkdKtz0pV8I8AhKqZnoXwjj3qijsS4KrD8kexg2zAelO2v7X7Mv
FvBVXRZbNQ0UpFmJV1ZeaOEunZ9VTfYyQhHDNeuWE3JnfwVUIr4igT+ZsnBFSnuO
BVR3ivMC8HgT0pi60U4VytES8EaiUtFznzNCEgLf2+WHr18Z9lpfsKu/LXh3q25m
xI5sPLphggOjv+ZUyNRdDutFgkWoQ2YrNIq+dNmezCA14fhyXqrFq1+nWEwi8XQS
f5NghmHoHfAT32yaETF0xFNqB48LEiEhqF850c7iKXSQG922BOJpPWg6Z3vIXtws
lohsn7AtEDupdntP0ewZghhXEmav29VsI8a8quTrjFlGVYmRxlg1gWhjOHs520UQ
CaOSRz8NWyaSAUD5kJ+Iy7UCsJoQc/MaUr2+yeD1qqY+9LQ7v7sPrtD+vVDq3L9O
E56AvPlVkK2QLyYA2U0wmK3Gy1mGojf6oao+BX6XxAzigjJS3q2XvY5EgOT3FVpx
0jcCKjVPDhNOq6CCVzPRcN2yxc4FJSGu722aC3xaL80hnJgdRKhPrScIP2ZEU3O9
XPSbiex7jOqxz3AOzWFFv4J1sZGH0ExAU1Qidfj36Fgj7IDoscDv9ZtuOnSlMsyh
8cZ+xYg7bfv8Z5tiH75AQ4rLhOilT2WsAsjgbFFtA49ApMIGdLXbGgf27zE1qOVQ
jsi1ZOvSzYh90PZeIeaEdjzXkjoqbO0X6E6f6ZWNnM36ZNt5j0cANGLbuXTEZaHH
nr4Cxc6+cyG77F/Fe6TGekMXs8tnpVjj6+Bj+EEsOI5AVAne72fCIJvj2GqRIADx
rCVy5lRnuvU8WtmcwRn10XK38XDFhJJS/nkylA7YTp34dzweRhyFeEu7GzthP9X0
V38w+8t1j9BO++PXvURfQXbexODpqSzNtrir8A4sXg06HoKXT/fkfzulkxJJdvhr
8jG5hY92s9JXXC6nhcOr0WcL2ppbThYRjzHQj/YibPjO0ZcgEWOyjXOo24JBzg1q
OAbcvTvzoSdR2asKqiYrp/k/Ao/hl3yAyV4hBGWPZ6Jnw6AmbBw3F8vbDiyKkMV2
StgfjSN7/O8XiEbb1nvUcX5af2fvvCcsuXRiT/kxHlHX07ZQx1NdXJFELu435TNC
1gMKBW00JkQtTU7teSweEnbtstgRPvnkjRY7n+auiexDLJOHXQ94w16JjJbcYH55
G8tl9cChWt1irYGnd3zmBPUsGRJ71iQZG2IANnfS34YlnXMys1lbn+nPrvQv7V3v
dmhV3ebVq4XVxlWHqGuHpYi1hGwOZQlxoPAsYvXbiTUHx78oNC1g+M2PFIVjTHeN
vVFLMpNrmTO/wx5azf/QgT4ArU/Chg3sn74KBpiZaqQufNy7WvtYu4HNjQRJq2oW
Q5Fl9gXvP80Wlm/374R8G0NcWKEXBpEmMsdbLjsaX2sSKCtjCwfRBGcvDoqoFGM/
l8BexHIcoacrx5Td1YlwAHGSscCHtFZYYCSqepZufBvYGfyj6rqNM686IVYPYzxt
nIwg1qpYhHXuRO+1jtGAi4hz5DCqGO9ZE0xKJe07Twv954TP7Fd5Ylcl/9mIeUuc
sB/IM40lMvVC6nKxZFUvMYY+QVWk2oCKnGv/lRXv14so63wMmBXjBM6GHRvUkyak
V5m4Cl6vBBrRRF5Qzr0qS4UpzJ4Gva2+FTRZmHx9y8knxBoCOXxzPwBl6M4bQZMR
G0LtdDSk0mXquoX+8c+X6oxSnTuIVTqL0pBYHCYLG28mnK5odHa9kz+6BTW3xS8B
MlXE74hd846bxUPJsAFwdfWfvctuJ8rO0T1urQzF1D8j4cQIxkBm4BYw3E0QbfG7
q3OwGACHbx+xuiqyANowm7te3vLsZf2/2fhs3NpB5pnBj+I1n6j5sFMBxz4ZwudU
O7yTSYzGgppe+cLGuq/6W+1p3o1IRUrMeU7hqYtwMrKYQCZdzqLo7n3gOR8BbiGB
2txPKUVbzVyVdGRqIThhElsZF+aGDE7PvTj9bEkPlTlJDGnvsZrRYfNrBpsgiZYo
8DLjpwr3CyXljxJzIXmbxm8KonAF7qMhdS4cB9TxDqbTZCLjkvtsyRiaZT8Q9kkF
Sd3i/sUe6iXePT9+UHOsOeR1dLgK6yd5lrVwXhvHwNDSz8DiYVbpvoDnR6Ry6yPi
`protect end_protected