`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1456 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
Uy4DmKguuKHGYwV9sMd7guvCWuBi48fdADiXN5hEAmLeRm1pYDWDQTbUwVS36Din
lgqaelfnBBxJv2aMfKjTQzcsd+4byo5F1qM18KRouSkvY5YInWEsIRZcftOwKat6
vn4dKtt6bFtXyBFyZOm4LtPzj7krD+AINNMQvXW1HKHx5OxyFRtDD8KNQBJfTChA
qojh2DHC3W7rW9NB+QsTLCi7j6Kiz3ZLdYl90YwkwJ+nASivT2iNUOJk3vOfd2if
wqG9pAUxeO6HWs5Z0lxVvLGum2GGRAelFtF2Yp8NvCtvSdWCcYd6bBEziJ7AjKaS
WRnosyFCd4pR+yxwPNY6vX/PZItjSgxeUMEjZ5uMf3g4uo8O65/PQFsC6o7T6lAS
yglZ1gNR5lXugqwLMF5jAr8GrLggyTm9vLF9nSOHvUrVkglAMNn/Xbjk/GkSXZ4N
QZ7EDuOl/ORYgYulWDaCd/JPqUYxJctByC7B+OYCPx70GV6Twy9GuQcOv8sm0Txd
v47n5qr7QWI2q7DMrAyCx6e+lEUJsLVRDfAdt65OhO4spZBLe8sW3csS3YgPr2DJ
kly+UfZKqnwetJrIyyW7s3Kb5MexAod+gon816ihUJvoVYuToECncmOBFac9VUbx
F0kFZmGSENE1g5HSEiSSmTobeNIATB4N/mMQwZlh0qorST3YohhJa4MiWM4NSOvn
6+PjQQnMOBA2lwhQeEB6VfITPGI0GjnGQqAIY6aZITdf/XcKqCI/4ocLY5bWbVnx
lnKb1EL4XyTspFOvj+QLoiVfBP168xX8vZSn/yHFFtY2lNmchLjjvm0Ouey3tb4c
XbMXKdyrQW1A2w+4A+JtOfLWOFrAYQjogssr9tVHvexTYk0wB2STYjJTRo3Z+0iM
68kT6aPHdpiK5Y8RWonuAdqueMjoa1hwW/Rt4M+vjlUc3wCU2XsUcIEisJcML7u8
V7NSfKKxOfCJ26pnm268bvsNeOrggicJqGB7t+awVp+TiBeKndo0pK++jiS0uy8P
pDE8CuhwuofrDIVoAloiAlpbKfjsg6c5q9n7Lm5PcYYUKz0ibbAul5nhWiEdeOkH
h18kra8DDgU3WIJqUqL3upJdrGIlxwG+Xk130dnZWeypEICme1eomLTadGF/Zrw7
DuLQr9xBuZ7s+bFK/b0rdi9SrLrkhn1ZbPPub75NnRY68rWdBchOZHU4iUH5G+/H
eEq+jNBjnvHYbp7c49ZlfWF01tuU8NcGzhT0X6wdzHJA2KcvC8mF/K9TPpUB3KuL
MhVAcIKD707sdJhHbr1XAGTwOVL8lK7Qtv2WLi0Z7Uzj3jQUGm+TI4yJFKcKZx0G
/6yYtxjz2yyJgR9mEuHBQ8nfJX9u2OaqtGC6ev6mIPpOTl+2CIicKXw8kQI7klYH
UErV04xzQh45/NN6+pEH0Bm8PUYj7ttsRlaTIMqb/b0kjYGCTTCw+cbcM7zuMD4R
5ZokbdXLsHfy1IpjN6ZnrKVvoEbJF4z6W0YdLMIbuzv+TJs0x13CTUMJgv9iqydb
XPXrpLKldiYtVOfSnPK6ji3CK8evvgr24HuhiR9QJ7yXLIVs0Q//1G+7FrJaWqt2
G9dfSulol2ZMb/EeZdajPME7Ig5ZgF2eBnWw8YTjKnwPP6IPyBu4XUjS19yrXwNM
Zda8Qd5krNrv1/8cDLiZiLZR7nCeMdBoyYu9JUOK9Q4izAV1xMVS98lSb8KfAx+t
tYLOJYlyNqoEIXeYU9wP1UelK0nWJtnlUVxHgcRkVLpzTEsLtBZ4kxDEdBNrJK4W
k6wGGtj6DPsZKgZIcEDEYQ==
`protect end_protected