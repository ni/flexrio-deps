`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 41760 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
dnVBOIGMhMFpJZXzCENQ2HrsXQl6epsP5gr1KiE9u6RvSlbc/bj1e1MyA6Z66kQ3
DnSU4I7VI8zU/kdBYZ/PjCoX0QqhP3k6PwgKDboHPCyxZydN6iEgYcS2Em6iqQK0
POu8Jxmu+usvGc/dYjwdXyfcJaQYTh8SQj/HgGHWKAtGJ1wtr5DSuUm1wBd+lkIq
C40PAyJJo5CGhAZ2RY0TB9v2HERdpSloGDIkRRCT7jbeZM+5KMOFJFj5ojBu3JaZ
7fzZHTZKm1hG/8Mj0MYL94b86DbulX//+PB6+J2Zwf8p5TxW7FkRlX7ws93Jx6R/
yQ1DG0rfxmdb638zkZYGyf5ys34ZmqpRXLRtG9AYkemHukzu58uSYEEBP0CdfPRQ
flAi7b7CQ2tsJOziTqOLfv0229Oad1yd7u5NswNLF4sgFOlCb0L/uvaNcmTktftR
WBoiLqH9orijYu/beMTEmIWfbOqRlQrZtnpqUPDlPOCzTFC6mwTWmwpxFPPHFsa/
cFZuhVVbFaoZkRj2DoSV8VbS8tutDTiC0cuR/x5YrxS1SgBG32FfUF95QkLe9fW/
VAcB50lc5MoelQvRtLOVfobfz5yQd0EMUt4lj9i/7K15T9EVTb+bcPKCt0HwWq/D
WNvo7EkG5gPfcrLHFMPYrUd808VWh8FPf35Ug0nMrtcL1lcdzQZCHCvw1cT7VY2x
PiQpLP+KDsDDTDRm3mha46BqEUWMAHqNQd1wU5gag4aw4VokmBEZlDWZ4lrI6SfK
LvNfIq16LOApjxTV6mRXSqu8rvlb+hSONrI9oBJ9quBcT7ku+u/jP7UMKpV/Ftum
4yuowy5kNJaNpj5VyyO/g3e79hS1vSqqm4fgoolDDJ93gBeZRAambxo3uIts5tz6
TNKtjxi2+C0kZ2kK916xVoRIYZhq0InTv3y5UbN2hllvbTgCzKO9bUbEoGBc3k7O
Jj5c4wRAOVgctN1VT9iI8xM7bRjbAgYqE/bSU99CsLC7I72FzCAjG5W3YCH0amz6
Dmql3EZaqVhaefRVUFi5R0oLOMW/G7I1SpLcIitzmUw4ZHXZ8kfqiDwxMdfAIDLj
PZNJqcXFs0S2t/d/nlI06qqqqk09j8NIoU1S0Jfy9n7DhHOJSTWAYtSJBk9HpB/D
h4LoyaI5sh1IF/moQjEHfGzYwMRJVGmlI8ZVtJOymNQWTnXxyrP3wmYfJmDsc197
nBMs5I273jrdgrTwXBO1YWVBqNOl7X+Lu4rp6RAvBdPbjvuYign2JgPRuuskf3Ee
pT7RdV649+ko6GdecnocPXEhvQxCjOhoYcokLZv3M/LiRZExF5voSxWS5l6c3CGx
bBfWpuGTa73xO046l+kqfuNcH8ZCrHyl16LBusz4JyC0OgkIpdECm+hIRlYVUP34
pPyCO9c2gUAAy0UvdVn1pB2xak3EZbWwICbQ0T/gLeEC0cvnJ39rZMQL9q/Cy31w
OU4z3i6pi+U81IrZWdCsr1JIwd/0iNfwS9McblceSH73Wf3jj89UIS5bp9m2ud7V
eTcUXf30Sb/bdmz8wnamnr/Pf1ZbONQ3hH8ojYk1m6hO91pI3IdZU4rReBOqhPV8
mBP+rT/650mMXJh9SXbpq3A8RkmtJ01qzbt+lvEwhdo68zu6551C90F7itZjzYF+
B4dhXqGFCnE0attGW/YrC8Hf+v1SEQFfSRnoBwrL+EONm7sbLfQlKS9l0JvL9+dI
S6vD6YHCoPP3wZQg+a/91DN/VedgQUXfQ/kOwZtMUKuGl6KHrORK+td5CvaKfJix
ekgJ4BetKi978GR1JHf8aLPKWegPVqR6tWjVY7RCDW84GIgb7hcZFrckSDWolND5
K4YWXCzfmaOW6YlyyqQwSNS9n3/YgF7vOAWN1gErqbCZkuIAlPyZaIpL59uvX/NX
9KEKAcnt4z5k0NZWtnsoXUFWnJxfflLCUHgv5wmUapD+RB3wxj0gn5A5+vyEJGSL
DzV94DOmRUvvsk4sKcQyo4D1W9tgPtFBgJWD61op+leM8vwfBMj59HeO2xu1Ie3y
rR5WK3Gaxz8VZ149hcudHpRbq/LmipZOnGqRC0x6sDFFyDyfwnnIEGBW8QwNjAlo
7ozqqZGud/Z3Tm0fIGZaHBybcwr1Xr1HFJa7bXOB0Ho/2bUTE0ylGiFGjwVLt+ve
XSUakElB8sr9wQdq7jEPzyCm055/fzpKDGyvqlviqomWKO9CjDKIVwy3MF2tOVUv
amKIDKiuQ4ucIZEKle1JVOzDlRBBOXLEhr1bB3VXI5+Ga45fhj+0JdYRMEa5J0Up
mDupG6QYjN87aYIUIAJBJ8bm2Zikx0zZgP30YG90Zl+10ku1Qu+ko+46ZETs078T
5YlCRsh5AIXru4MCsl4awapV/Tjr4pt7qICIkSGLQCP8+qOD/Ke1KHmXuQXK8csM
eWMJVXKXv3AMer7FJ1nN66RgONEHQ9rGUBte0u22y0tVhO8its6a8y+huM3/uOxS
bhMbRRkq3YOqg9UHEG+NaOQr8/wQVoQTKX2bAf7Tn/oDWRmIFea4wfLuajr/aB7R
r8pLz15e/xTAZxhPMnMK7bZQoZDD/zy2VP/01pudpoM7sLQlloREa6gOKkrVoHik
FQeMg27iOgIROoi1uM840YZ0UeF3dbY9VhhTM4XWtPP7OK4gMsK7ENmILlySx3Pb
QvKnnP3+xIKro7s9O/HuKXD2CngylC4IBU2dMW8Swrs2MgXl5TUgAcy+DF7zjEHK
AVOprVggygOsGR9jxOs4Z0rqeFUrTQ88N6XCooxQR4sFV9hgqz/20BkzuHCWQMjW
t8BdeYFUYGmCA5za6HZrAXnvKzSw6WUuguuV+Z5gM3EqOWlCq0vm5W10e7rBThkw
x9tlwyXwvSjoIWTsJ+/yhl8tIuic/L7PGbVpLOaQhuV0U+wekSQ8sMuwt8euAKJb
aRM8vgxXj9etwZHZdN6jZ42gGGbL5s8kTUGLsl6no5b6d4rNh6FZXA2HM4DpOEnn
ejSlse76KrbQLcNAYTZZRVyY3DTBFzluWXn77hpgN4wbPJYL99tUpHkp12iXeFcY
w7vbHAi+5G9UF6r2fqd9+PY0Z8uzyrsZJIYhnSsMwGiPHZCBg35B62QeHla0VbFb
3lW/Ytv6te0sMFAWcGC8nFxUa8EOaS45uNah5c8dOpsvcor3bxrRLjdmo8YEAKka
RbBMx7ZADFMaHHYu2QIE9GCm32t/jHNYf60cJjExxTZkXQIg3Xgdg2y+0PmzVxAk
4W6O4uEq5MgyaOyI6nQzoirXpfQFddIpUdEsHbFi5BwOnb/Pezr1lZt9/Ox1TpXy
1H4771jyz7guSS0KZhCUcHzVcT7xfVU0Y2dyx1i4zInsnXAwkrk2m1UhDNjzzUOs
VgJ5gG3dtOZInhcSE6H5QIXlZNDGrr4ld8UzrAIwG3ufqotlUTzccaq3a4+gdcJJ
TKq/pOXW9KwC6A6zLXZHaWh3I6Uru0/Da2eoyL4+mjvDGYOqbYBjUte5El6dQzyc
flF35Ns0tTK29h5kIaNDc02pf5pnE6jjmdCFGb5IWQZ9o1yO0/A4xw0+ED0UYcxy
o64GFzSUE3Ptc95h9czhsZVzZCM0kE2DDaXBphN00nT89L6ZTmac1p9UgpVrJDwY
frV9HYv8eCcfNZx3mnTBtUzh9QN10mngyCuyL95SuHOyZkwLah9rk4nm1S9qliS3
Mx3tgApnb8Pgac1JKCRyu01/DHsjYsp7iqBkHoK567cHOpG4Uz8XoyLRtnnOAwcB
73MX0VHCmILuGLm0hFokJdduTkVClEH624O21lxLgnL/Bdlonq0Yvd+kHXDrBYUz
NPzpfxaYn8W/SqMeCMOFNjtfz9BcYHIJakGXBS0MI622yq38gDVm9vyAVIPTTDK5
Ofpze4vOvCneqRBMM0ViOu5Yw7yZvHeYLTDEQVU5bFrPx2mMPh5vqZT0e3ElR4QS
Dt4qPkyR2R1rCxvF78xWHk0xdnodSTzOuOQeFVWfQID0hGod7l4FYzhpCQ79k4ci
AXJuAedv31WwBiWcoTciJwg2/VxEJJqkATuNI6fEwgAah4kMzFQgZMHvLygMl6wW
tzf2r9DTyOHA0capTmv7tuMthwhx+0mMNhAD6o6YYQDcE+MRReOa9YtBAD2FoTSh
BZM4ig36giApzLBwJ3JTpMqzd7bd5dVHNIPkNkDCtIYrzh65oFktgFxYvn3SEvFz
y3zRObrGvnGXvL+KM8SNPf+6+RD1Lh68j4RPhWuV4u09tsf80rUH/11v8bgh1Ez8
zyfKENGd4zLEFmsvC+qztbQrFFtnZw0/RF+cMynr8Ux9qemGZfQlvjnBJ+Lj5oEn
oGZPhaHRQ7Uyyblo/VDk12mROdb65MM7lR2TOGu3f3uncAb0g3ME+u/dk0RYiWol
amAoja51t0JWIWpDD21AslD2pXp0zrgqTjSzs+j+m0JTXzBy+A/HLngwAFsi2yRr
yQL2g05dAJomBUIdMvLS9A6qyGZXbNYGSwoEPIUPgHu3XhVnzCZ09MWpyTD4uKVQ
HGA846cskalWjZezn9wWx0Hq/yPIjemH2PwAvps//WwKVoViCR+nXdeF895g6P8p
+fAVvLmQy0ucvZCXUC5K0nUkZgVnjMTe10cd2hcLlufNV/OxiZO0M+kGGZ0pO+75
R8zcaj5nSm+bjOfXJWQ464kGqNxiSynaaFhcYpgR0SsuJBOjSfY2Z1SUvdJhF0n0
NIag6iqV1X54IZezeKOEtnDfcrpmRPZtwVqXAHBJ/UMS7G2P3fGZhZ2VjYjczYiz
OAtsktQhHhLWDN/qULRRKC6ZOg/DXQdUOK2NcZUKcUxjAMM4MInW9KU9WAvo2HVu
4Yg1EEI/f3fc/DcdEutZrSwUrB/qpmPal7SQaTluwvaoaXtH+gE3c5rAuMVb2Uif
D8lb2D+HTJKHdHh2J6e7MPephslvJQ1jXXL4+3agfzKmNCY5miJ18ENT3KT4ITYb
yHrdmJRCnqPZW2ZHPB0Pr49ZFfPHFq3AEmuoxCoSpnPHqp9GS+UJD4Y91RfGDuPf
SpJ7rb/aLH8W35K2C7ewjUv0QbQ1LjXvfqEy3E3UNFIzGr6qVsAXrtnZ6EH+tfmp
TsMvlVUSrQcKE36s3mipee901wNSm1LzeUkraEauHwUcgs90UVGrAlcF00N2bDCL
XlmlomLNuNL7XkFcgbWV0h6ikS7jXsxJ0ICPrxNG5fsYK6MDGgDSH155fegDm532
hbU+xXx89inOZ5esfVFD72Al1Jj/e8qoSpCjY1DbLBx5/x6eGo86tMBKcWcOAumw
I4g4i1z3Ire2IAB/m4/WhQJTs744GYI+57nwszMLcU2cBlnXQbFq4aG9pnv3iI/W
d2jon5qhj/v7s5TfPoXkDU/4kE0yOXAHwVYk20z0oFE9MS7PGUkOeme3nwr0zhjw
WJks7xJaQMxl99qGcxAE3nMiEpRjclBS4eYPlxio60YAma6RzOXrebkP3xPOkSXX
DbwBfHZ7wICl42GdMREa7j48pVWqdkfIg0W0qTkLqpBCL5hBDmbNTmKBIm6DoRcV
efS+wlVNIhv+i/jXFumtJVtl6uWplJ6uozzRo2xhDXfJWZ4mXtl4XEw8LI8jWJLM
UAzUDsX+o6d1/peQ388C2SHefbkYTSTOb9BnpqY3v0v4AmolOdkZbE2J3ZjJtAVr
Ueu1ot2tVnwDSx05ip83kq5YYn2TlzNYVxRHavO589CprC8/7Lx14/qzD5Hdb9xB
32bsodNxP7ynXY/33jmfr7y94Hof8fgVL/PbBIvA9KUQWiTcQ8MD8vO08egXadql
wvaW23ESmlHjq98EMlmYBtCYoOGlm1WLOBDk1tpiTCr9GhsiszYxNMi4kxsWB6i3
SrNM+gIdHtHxf94YiJhP7off5RHaMeHh4f+r5OihchSCB6hvub91anZvLxpQ+R3P
LOZKyNrIoxjO2ypdqR0sZwBQthGKP1+S2fW+jbD+RHsLfZdqlWpK05xVMZo0YI1w
2aPvtQMMfBOwpnvfIrgP+rK/g3tTAr6Ji4FZ8ILmsK2Ba6Zf1+78dEovLI+0IoMB
NnSYo79i7aUdKgJKm9rJgmgzWTbwRgyZpBNpAtqGs1yybVbPah4Ti7Jkuj/Y+Y0t
ekdNmI2hxkok+33SJHBY0Q7rmIoPTmXuQBOBX+mIqljuvYQUEUfIaygavCHi0Sir
lhbXJjp/+kPueKpqd4shxJ0hA5jdFhyCKu4jr+OqtCVUjb18WN4IRK0pVXaNX8fr
YjZQnggeJoY+A7yMGg86vL26yOsGDvZNJrTssvAxckF+hfCVq6ncoX5lQrNhGn4l
+ixJ495sqTxS133f8azk3ViELSRGlK1EkY2u+6SUtVbyU7UeAZFwGW6zuNfyjx1t
4kPRo56abFVxj1Ywdow+6O61UPIiCrrc2JINir492mG/RxF+WlA3oZNvh4muuRQw
6PJySkqqQ4mVnC+7ASaFYYWDde/xhXisJkFyf3ngMgmceDe+necAWZKqmq1L0PDx
fELVGVgUAkfVVdbEMB3UHoa3uZldkJjcmZVx8s2y0bAGREqsvvcgv52G6Fi0JEZj
2KXWYSn+qxk9WYk3iUySPSBEfRy8Jzq3hksXyXwLcNxnEH5QALg/cojKEeegGGHg
kE2rj0ZksrhIrovyIO7LX1SybwD3OGyrlRTsitKx4w6b8Hrzr0/bu3WbZ/ACIVtw
RcCVWOe1EHy3RPywPPzvu/PvxRp68CDEgOnu5j6v/2FoWU93lI/JBZtcE+2IR66d
ZMZnXcsjbPyHJ7ooHLh+V5mdcKrKFoQAwwNnTZGu8fMLlcbo7Ncl3qZV1xkpVWgH
Ul9wJZsKgUaH3IwlkGqAKfnPCjsvySwUUaI3Xd8DXr6XHFIKSE/g+bDwm/l0PErS
U0wdc+UyJ1b/owOU0HsO6vWxE1C0W0Da9YCtCYn1w5/sGjDiLzc8fTFa4jAPkOOV
eR0D31+ym9KGZBlNE45wBm+kY+sLZC8Jtdxt2HTRwz4YrvkmlMDdgIwNBrYDO/7S
aCYhZ/GOjOs81NDoTZUvaiQWxvg1dnW1tpuY2U9pUyYuCU1Dis2FYGhXjxon25MZ
Bzh8OJprIxL76Uflgbs6RpQgqW9K97C3yaRWNOY6M34zswDPqvqUPYpJzChVeIUG
ew73JFXEh2BLrRNhKIwGQvQWC2Pteec5ZygtViw+FqPKiADOx9DIUUp89FIy23Hl
+re0PIELaJh8t+8u9I9XuRXcwCl5np5QhHGQiuFKFPhIO0udS1zqUQIhkU4tCyeX
E0Yz0K9QlfAb+My/cTdifpbdjI3tuA2f1oQ+ZIOzcqJR9IjdbJk/OAE14pVWh8/a
gkluXg9nWK8519SqFuPmaHS+9ZVLHTLisbbsSCU+ItZTZZhCI/UHukiKbS9gjXJ6
JH5zr0BKH5iZH0ila7iyErEtYCJ6CrjoscUq+Rm44jxECCMKvXnxJ7XbDZXHLYNo
N2q03Xh/F7lFaODTyKb3lzVuZcrg75h1GLEJ/6iWgp4Ne92BbPSaowY8sj5n5HSJ
R9IA6nsn9rGNk3qQIM8/BF2D9LLvl++GtZPSE/IWAgsZ6T9L5mjYd4ki1/l0a1b1
GVn0mqvBmRHyf6LidPhu2wgsIk/JdQhEyIjtdEfKm2d3vYDHXqI+4cnqAUxHREIo
G6sQsiXqer1kGomcLgDYigM4oa0OcGK3bgWgx2y6wMHL3CqVPMHtOazPXEDfNSxv
CgmMh2WRhGURDgK1L7tqPz7MV+DpNPSsY1+X9hpD0hS0UoEnNsVzbJCCuPqj2w8M
6dAj9Ln1mHxI5GewUwP9VXVqyCAq1llQqdBYAOAVsjQ3D4fPRYzJVQlZhUXvy52M
sjnSu6UeOFsCKe6RePI5Du2LfvmjhcYSSHCj+pDenvrz0WJQvbFszkpHwaLmf74L
X0TQ1mKP7GKXfNFAlHsND3d8cKGQmwqNurjgHktt44+zisvw7VsaRMNn1NO/xFGY
WK48A0YyeGtZCc/HzCjVjvFpLbII65qDttsU4dj2wKOPIttZwOdUlrFa4RKKFsII
bRVSIfNtcygZdG0nISDAQjdPFwMpm/czRtmQHefOZUCQdLXQSd10WXmH3rl4wwqv
2/gfKTW/y3QNd+XJhpQpCb/DYxQo9iOlIr1c2tt4+w1xeR4BA4Be1HR3W28px3Tq
JEdhM4cFIh66qe/xhwmWdoXwF0NA21e+AYQ96ZPl3Pb3huotxB5aITVKH2iuvU6T
4l584QIPrOcWD76e+NlFDc0/Z2DaB4BuuShFXCIUPGKGVfygIqNb1suM6z0G1vxE
8FOOyrJ9Z80f/dxF5eBX5yTba5Qz3Gy44m9N49WLW1YY+J5webKPsUSJs7/aZ/HC
r3764Z+0H2rTS2eSDyBwgGpbTIXOpoGxqtM9Y/k150VsANUuoy/B6wcrXogAtN/N
CxFnRDgdKBtw+qbF/lrxUJ+F61Wru+SrZ4k3H/sbuozXFcn3RsyWE0pXsVucXekG
yUc2mOtOnN4MGHfeiiTxONIe3Az2ChXH8DVaknU4tJvQHP+l2giVFdxJmHsJpNDj
UKRtkNRj9GWbvhpiiY08p7NMKAZHc+ZJL+cOhpzqn7xVnKzXXNh2n6gfoOCsrUdP
7lMjPTIjY2tAXLt1CNr+/quwwz1IuuE9lcho4dV+bAqPlTSh/46nhcHgU2UTK9vN
4Lm9oug9q9DkXN5rKNMavsj++mng8tjfhETqmQ0jIX203rZep7UhjwEmjGg5Ih8H
+hdHLK0opOzPUSOdTnBxCh4UHRHsFulrBC6KCcdlCowgTy1YhWVrWTg3o17RiopP
UB+uUwG2D0w92Hio2rbng06gMa8xFaChhR6dCj1K2nEw4QaZHHZHDyrYtmGlxW5Y
AWlKMdRA8oGdpXwuAMV0gd817Pba2mcbdytsSMh3i6WLGmXDaV1m82SHqJiYn9Zy
BV2SiZkNJ9WUFDiEISqL6EijqbAIUqzhFr3zK8Vw600PsXFil8CcLTSAW+3cPnP+
iV2VuXZkR/dCChrhtIh+n09s5oyaiSFI5sSX00O1pBqHesbZ/HqEqAbSJHmI4g3p
JLP9sBnvfhzILMgPpQgX4Dx9NfsGJHDdqM/WS3E1s1gBalQh7ZVKsdaFPhS+jku6
ZdvoAcjLr9fhVJHOuvtk6g7Mr9lrMKYZpcC6acAcOqrCFDl10RoYTyzYTW+eh4ow
ZH/17G6MOW/xbN5T6xqU7ZZx4pp3VaxiAT3O/rBb0Q8ji/kdgCtGW1bElZfgHdbz
cScsTWK+5biyl6hQa+QryTEjD9zBexBW9a4zhjBmCBviKhC2c3fTx8aKhSqBtntm
IBPedr3b1q1HZAZqr3zo8mFb95mm2SJGsXpvSDSpUzzH26ydTYtqOWQmgFmH/v+Z
L4a6GmAxzVpbXpgKJ7MC4W7bWxc6UXZMK5jeAWDlSHun4CDA/ZcPy14K+sC0v/G1
0l+aqGrl4hf2kK5S4B9dCpge3+FtD6l3hISyrsdMnoWkKvJZN6t1T4d6KMVoV03u
tryb1vET3GMoaslTmGZeePjPTUy3Fg7f/MOfCKofb3s7ZRxccLExZCQ/b0oK3jfh
zCwv9hMV9TXHISLPsoEPTujJAZQx8T8/Z63+TbDO7nxzgh8Icj9CHMi4ib+2oeDF
nQ4qpsPBjtqVUJjCfM9+Yzlx2mMrCExIrmHPvQUsS0p9v9H078g2qDAu+6kVHKHG
/4945XwX0Ie3XUl1WqGNCJeFi8O61RUhRPdMBPW3edcAxsyAUbqa014y3QKLfkiT
v1Ckn2FI2nlPubQAjt7iP7imRv62v5r/iHECA/rJ5N1Bbq7D0YJ/rbkXIa0v3nbj
lpKP/HX9QTSymvmhiMCXV3eh0+xPwsMdooqVmt92Mi2RiDu82RO0Ko6QLlQ6iy6E
CiC31tTUAFMuSw/CuFjtobLgZhA1fUSj0DJ4erCzeMaxPj7PllQKSp15gmyWcsNV
pXlwKkXOK96lKe3e919VT3rg/xgRo/d96YTzeOX4XPf7N5zk1sRVoiinagE10wcc
OAevJ40T3/VQU6LnKwmW2RGG+FB1JhqJUmtEEUeTHBYQk96yAXLgFQ4E32HWffbg
b6BwONtaIlzrxmuQGGXs/QM2uY3tH7sHz81gMi+hz1ccoKAoMcdMiptgqUNO9k2N
yECZB8gHtsu9nGemhqtQdcqUW8C0o78DsoNVYz2sx+s9Q8nnxu99xuFk8hm/p3aV
48s1d8Ylaju+oyHBX7kqGiqbDP3ksFNWLNZlS5H3Fq8vyy22LrVVD2ejvtT+izTm
glwn4WWbRn1EHQja/R8gr9qSQc10qFf6lYQNP74/iy4yfY0QFNYJVTxn9HeAb50J
CWrtfYgr++EGNynKoyt2NyzEopwe7rkM3fQA8ZpblDEAH8lIiadSvoi+x8P4TRf9
ZeYA8lpVNIqq5L1YDcJ0RCxSpaCHzblXnX4hKa30JFOUxQ3gEuXBPszLqhv1A8b4
DHqFV++4Vzq2Gbn6dZbX3+HFobJDZxbcHaMAxN+P3E7hnPTkyKFTlNuwzKMnP1DS
KOUEXpAnwzn5OmLvEne6AI+OqlPc015QE/YDSNjKATIk3cXTF4i9o/1pVOuGn777
QF2nfcWW7NBhJl1Bew6yPgXuHOAbKYGv5jGxzRBzYYXy/df+po31EyO4mKdl2o1r
VvhruI+TDNvtKF86aojL5sgQuPPkW7TNCpQYIyIx89f52dWwSqf4k7FICLsoVDUs
MsLstUUmwhUiCTdh+woceaJv1daMKjw67+aZZxqZBMmuJVF5GFTPzuf69rvr1Emx
Tx32EHlKGy3MmdQwZIecZrqitExVqIUO8cWRhQBTQue32cyK8X13w8SpgwhK3Plu
lp5Yf1cqEupeCHAzPszg/z/H8xdeKdCo0e619/4YTkFz2HwTpiUlSe6+654jAign
Tlllt3fsYMNOd+tsC6eg0/v3/JUKxuPCjdn2nTiwsGnnWexqY316R4A6TbtVj6MD
Y2k/r6OeAlKbb5HvSg/kAv8pBoxTR+TAVs2ibSAwKBA70tDTkaYVZT8UEdG0hQpI
WQvlhhv8K/dNGt28XOHKvR8OH/e9RrTXRF1OjfquFwm6eB4Kx7J84RFJU7jzBYwf
TEVgu2vQvAo0RV9elO/0zRQu4jm/vYdv/xag5SmJwrMf5aGawCg1lXfgbkdEP5zw
FiADlY5VTFVD8Z1BFNxsu712ifqXZRGMKjoTLd3ddoprCRGWo2s1fPDlXJVQq8Ry
EL5JTHVDWhCJpsL1ruPxyWjI2QZCHDAIlfHS0WlKMm2D5VaL/dBgS/qXcG4G8Ck6
IekpmxVHhRBY2a9WWfSyo3SEKUQUBjbAO6o8FvAEWYcIRV7WpWk/YKKmDjGRzd8M
hOSglFMGg6Y9eGLXGj/HyeG4Oo9nImu1JLQlZ2cJ32q0MhhbAJSLB8FOwLF/y286
Lw6U0n+PpCWHoH2lcjNGla9e2ye/wMPBQA9+ss6jkDdMY0GZyXR4tp5ahs9Le92z
HBfnVbb4VWXGdJm03hkuZEeV6LVPm5ihcsPIlG48RbPnXnLC8uy6z1da/gAa0soG
5pni1z9yauwTykZIXQlWIYTdtzeWNoCEcX/4vK26OuRrZZ9IlIyPI/n3F+Znaixq
vnGQxxw1FbQTlgNl88ssijiZeHbbYP8xfnBNZII2MfUNhtxgSiVQBMKMHMLZONqD
AvvmMuhwg08wlGc+8xfbrZ5R6OthTZui/xFlFiQEmETAEThyvZ7OAK6lASQo1Dpv
0f+ukRrY0m6XOgO58oAInizuPnuiG3a5J8dy+2KXIRkG05Qqa7wDDD+0pTciEVcj
LjqOR8u2zkQXqz8lekPYZ2McAilJTjLzS4mqd4QsG2X8z0wigx/gGwgXa6x83lZC
8mIMdwj3Dh+s3Rm2Qcg0OT+sghjd94JKXHDCJaI8PkMlP2zoM41sWqZIjAKzk66J
hBL26HkbjRGGibDUG6TKEobh8bHJ02bUl2YDAvtwpYpQxmT5GTc8Hl7wC1W0PAWJ
MnYJrBmkddzqu/UByHJpg6lguAoEKsz15ZbGNZLWHaacTOyAaI7No/W/u1/qe2G0
lsWp+3wfViASHolGkd2dAT63E3ytCQ1/FzaXNnjsjino9CQ+Re+o5MxbHAGb01Zn
Bq5hYb8sFn+TSlksrwFoYR4RcEeb5nLdnI3rTDQ7OgRkGUC1SzgpEV4imbi5qD0O
W92XDTNedEIqbh7LUWN+GA7YL/GmICN6LHvDX/sCVOwHVN4ut2WvUm070Zp/es5C
KjAA7WB/sOeh6V2Bqc14WyDpv4QxPwki1ty9HjcQFzNzSgy8W5J510KDI9BFK0cy
I1BtKKfIpk40AtXrOPu6r5JScBwUvH9TFujChniIGavXTDyAzwYT91DxFBNGP4Qi
ZDvMwxwoNvC92a8C9H8EQUGEau0IcPF9GVWsHqekp/hMKWDr4+uiUDiXk4NL72o7
hrHvTuQCrTJgpa007hsoKp1lgsDqTKaNcjaD4z0MmTGPm753K8HpS8ZLwNsN8Frt
3aaSEnE+rRhn4gaUI3AJWm0S5EIrsKVg6VKhwrA9S8X0srCg1iqX6mDP4IuNsNKZ
r/X6rlLzJPPeFj7N1mlsovUlOiPwZL9b+OVy2o/WuJd0nXOcx5iSv0fhafoYGIlU
oPq5nDC2S8KW7ENrM7C9hKJBcrZw3qRv1mGkjAv4H4qIm+pg71w1EDs5uDODawap
+qhsk33qrh/ODUk7aCrS5+BkFFurmBX9iiJ7PTIJOrJWtaUNf2aaTIiJWaPCGun+
AZV9jq7RTNqxgyXpAlOJtwbQBzr+sohl+eZ8fM7l0iPCigVec9Yx/B4MphW8Y5q/
MWx9IZTeIW/Y+0caWQrlH4+JqGKx1zBySxzq+t38atbNHeLvoUDTUB221g/Itlwl
nCrjkUfYPrphGFJltbfK80Lru4gf3t9uybdcrM/ixcyRK2ii5kgGe6o6oL2TKBy6
cRi320Uonq2j3drjCI0bZ7WWLQuZJeK9LCGZgW29OC4Y+OK0evF/ZNmpwPv2l39E
iWs16dyYH6UuaJWZHkMk0+M41IHWeiFrFg/HWVLU7SJUYbssor9E2jygh8vlUbhs
OELbB1xjoodkTn5JpsKnb78Q1W2yvo0fqQrcLvDFUHE6BE841akF2Trsht4QN++L
rJm3is4QjBJWlLqkGKGcWip70H7zZAfkpedjTQ8IlU2j62Nx4xO7szLwpoghMF75
aiJZqSmGUdRC0hMZtG9Ibr+V+2auoSyJtQfA+OQa2SISKFysIMiInIJlgmZSWWUa
1cEK+G3MimRFlwF+AHa1Ewdv8PsTQXoWms4BrEhIKjD6tW8kJgFR5s39L4x9/HNU
rHqDjE1hbu/SmGlzlvGhpRRYz9c5jTnpoEP4d/DRwt+XUKHdZ4oNMFJarmB82uvu
Wiv8+0iA+QuRtx3baYTEZS1E/WU+VH4y1zqf1hHfCnn8xMcKurz4VRrMr+Sm1LBH
HMgSdIXnfS4gJy/Jzl0oD06imXIVHcbHZhCfTwU89gJMgei9QsXphgi+Z2TbUJqK
ru9U8AkHNDW1BRfcp2y8KAzHk6qa7FrAFPyPaElE0BNZ5/3r801uJQwKaszrjmlj
4fevcwkl6d8CcLAPoqoQiJQkVE1tV83X4E+1wwXLt6j0GFRtJVmzBLbuEG6wAgyT
mZIcNwk5bOpQ9LexH9X2FIC8E18Ae1WEUPF9H/Y/4h7oQONBc7edEETJo4SFIT1c
jNMNUaDafrq4QYUYuRzoDCS0yD/v1BUqu5YDnrq13YJCnl8H0jJXo9nSkksdW7IH
T00nyxB7JecrTN5Bon4cv5/1jErY1VcGSrv8UUg5R13JC33lv7Cggow+SyT0mVjW
4WpiN4U418O3lI/MnJF2uEt3Bx72jotya/3JilNbeYKPbg++H/IlCTejGYQqBQB+
PgSfo0vhfypC9HiHL0SrmaSIIB5lvs1PrVLq5ccxK8BjEZG4etBhJn/qtW0CyZF4
xRqyxUkr/ga/OvcNHJa/5S/aVghWptZhMBKO50+i6nxA4eTTrhO33nT9z1phKJiy
ySFZukENlQIGnR/4DJsOI7ci8ca+E4D38eacgJm5aYJj9XtQYiSfTnyMkBuZH5QV
+z58idoI+7+TpbMBBRmTdPFr/CB7aLpOkU6k+NTz/qGsndEUUw90PAvObE+/XGuJ
KmsX/D23uN87PoMBi3vWiFs0ntNPi8xMRQN4V0ssaEI5S1oIb9iw1oLprUy1IwLy
fsmKy3tN8dtjuf8dDX8w88NAD2tfuVl3eQsy3CIsLtHM0JCPjBNEmT45LnatSNgX
9ebepbS2mw513976S0F5kZ8pQZH8H5pC2zmF2FXiCWzLTDNSLe+e/PQafS+UeQq2
ZtQ4RTi+OcR08z+JomcHaLXQIpxRDTVfBN/wo+hnt/vrL+VjUEjK4N0Oeghqpgo/
Jg/afe9PcG7/VsmPZbbU1R5BBDW5weRhLQzRhyXSQ0IjmvxrmV0++mVmTBByDUjL
ZFRUqEcIX80JkAuXpCom8OcQ4nBbtaMuhKN3RIjVqNnc2VT1ZM1WZQUsXHij13dd
1nv65SRooVrdr09HqbaEJiIhG2cSl8MpaVHqygz7aoYvkASY0ynPuKGvKmPsTsyE
urKXInCcO9OYYMYLY0cSZxzeOcBQoCoe07kaGSF9h/PbJbQLvGuoEClgms8KTKYv
pQEbgktQfMX9zes9f6A9ku44xbdkKpuuic0NVJ+wThYYLtX7zColAS+dLH/enqZE
m11yGjivmhNK+uf3s0AWWuw65/ccRveMiaM6Fyu2PQF92fOMSoSIoa3LZp1vY6aX
+XNc1t+czsyDqziYZl6ocdgCWTFmpAk2JKX458J25qh/xx26Ww4TkHOmi4ZXDQej
QYWTt/7LX4ybkQuDW5I2jViTLvez8WmNCT5h5NYOjCz3pnnQ1jh5dw0999fJUJOv
DICSllEfBcwz5mZpR94F5lJx2WFxNKGMI9l1fr1vmysrWpHrYmYF6+s2OEPjBfa2
qOA+wbLS0pWo5B/S2eR0SGxcrnV/aSOqCZkkE9sGm6FQz6tNqkOenaY8sGnQjaMI
45Lgyyxur1YJbqmzrzMXapFaJoyG5CJ9xEf2ukWkBfKzo9ELaHpfL1pZAJftbjNZ
FxrMMPsqyHoCt8tLyyIR93BKNKKISL9fDIKsDfygUG7eUyuich0fCGCrcSh/CY35
xEL/H70qA6WrJfihsjnIXxwrq+LHMhO0B/Z8/4PTZC06aRhdynK7l/CzQ0gBhq0M
HjAsF/rNcjtwWflHEXIW9TIfX5Hu6Sn3mP1ZthvzAxvF/wFENZ37jpxAWrX+Csj+
KT6Y9+ZY0zKye8Ef+SrzGuUHw+byCYmsPlD1ChClfdCfv0jdRIMcYdsgeYRRZ+lQ
37U0XryvIs6Zab+SPjjMlLsqvTVYLyhBOOBiDDje4B5BD4sQLAa4sWA8CBpvRgYK
2jwfMsKLTTkbQUPQ/5bllcfCNxQ6r7xR5ktKlA7+nRuVMxBFmo9ekR53jLKl4KOy
RLqnRMxaMlGHw3o2VYeUXnIwI8g5i2z5nsgFItjrsrOM7pWVNF0gKRkKIRyGUSyv
oWpw0I1qhfsFbW+/iScOzvqWMRzUY96yjrg8YTkX87j1sooyWQyUiVw9E8wwLZAH
B8gwcEH61a0o8Odv1eux9hRxu1JrXkskyFh0Xv/BzP88JdI9XeJPtLFrwreYB2fc
V5C768Wdh5qogPX76l8a4uTGsd95N/T4I1yq73axOubC/ShpMVRroTgVfKydIPRC
mCto5gGIVD4b51U2Hn+tRwORsTuHFvDQG5Gw6LQhiLuhxIdoM9koko5S1m3Sp3cf
MQBjYct0e6o3yVOiJhQqZwmNLY9vI0ge7szhBI/TAHDUuYZbzbnl11qOyheYWauZ
oW8Vw3FeS4/193NOZj1ASQUJlQyW9QYJfFh8hv8gTJ0acVS/tB+c6dN7gyR5c3vJ
oYdVFaITULwDYBjR4Cc51+hWrv0GdWgR0WGMUlI/cnJvNjYJBBgzhRnXXY4l1Nje
dhSSlrPcPIfU33/hvnIIwo66SmrrrPrwqz8EXdWw8Z8UhnXmgrIZKogN4xZ642zY
bdUu5E1K1ae+2ppOvjcsy56hrkpDsSHJxkqbz3HfRG33sxU3E0R5Sj2SE1OTwM9R
HOj0GVS8fhd7FWEv54jW2lP2M1NO/ia+YDw32JlM+4zo+ECGg6KlVctB5nhS8J3D
+s3dl4QbBVIFvJnne+lni3gLubS39Shli6bOJi18q9GJ/oaEhaARTHAr/zpWkfbn
1Hi736RHl+SCOhmyst1zLtp5M1kSVJaEZRnvU99CYxOQfbN+07sLKtQtiw6Xj5Aj
rav9wfn/J+AG+Z2zXI/+9edTfixpMF3KMTV8cws8Mwoa2/VEnbO008aYar4qVShI
NP7HtjfEqA7k6MGYaLLQUqOxLb95iJzbMj3HR3qfNTxeR1GdR8avUlpER8T9n/xp
EVavdJInube1K+0Q4pcufU5+/Ejtu6CPV+Jpz3Rp99WwltvuN1yvhz0OYhSNtieO
t/8kS5KkGRLtU2JVrcua8tjADG5JexLE0UiK1qJo0nYWwo6vcKunoh0zYwZFWDT1
FdxpBNf/uf5RfL7oNWvEfCCkx9g3uS3fJ2fuXaKv5zGUfAnlDSc46yE5+3n0ovyY
Kc2Kn2Pxj4Z2fygEJfFgxXh19Izvpe4/JhR+ni+QWXIiA7iD8IWy2n+r3yZv6qub
6JzDFXngIyMSuoM4iXOe4EZKtf5LWIRTJ4CkFwPBE/l6kau+Ji6sW2DYGWvddr3Y
q+yf2ZB78GjYQZWu9oJJVScx8b4Okiz8HK7V/106o5/oPnFyLRGSTmZi4B7XUtNj
cwanKuRfsK9Nk2NRo5jPZbi+/OVbTnlv4Hv2gKxY7UtD/U1rvmHPmCeQ54ZATtKU
gzsRfzem9x0bfAycsMayZu5tS8WfJH9IT/w6GNIY4Tcyt8jyUmZbKMyT5ATKU1ud
ulu0TSeVcpjnmjaLs8Nb+8Xs0G9IsNJU3nSyAPEq2Kjzf5d0u88Iyo+mU2tlitcR
sl3NmwRA7IrXjNNpRObJm99VeszHoqdLiEkH4zAXKJ6Fg26/ulMAdAzsAqisc2Xm
BoOxOv4xQqj0wReFOxApQllV+Ma/z87KAXo9FQdj94EPyAqGzFEdd4ta0g3Ktudh
cLkL6soI2vqZzJ99WqH5TjwLsV9mjcRBG33uT8enro4+g2tsarIvqQ/Rjhmy1AMX
gKu+0ezAHHxsDEdG2kcfVS3/wYi6SY/e5PPKApJ8+f7ZqPhHB663Uzqf5j3D07uh
0vLJDtAbyN7+YgK6XYt6C8z+tB/y/I+8GAddgvi3ZNHZvMM/NYDg8YAfU19ehsi+
uQ3POzsiEtx/WWOs6TPgG6p897lTjdaqRPcpCSn0XvjdB5uGuKEIsXLHkLb4wrZf
8GT+BNJqahyScrtGXQF3QbWXulIsdK7+niiQ4oV6LNkYeyK/LyIDXHnHbIWSQDNb
y8lBT+h/l2xW0y9qBCTJ6wQnWnMvtGNXjB+h+6CW/CrEMSKNZ9/S44aCgGM0CdbK
jIMpVR44VZbdJ1xu34aLxMmRpnNVh2jRb+tRmE2ZgiwOiYFfV0vXbkRy7H0j/r4L
Ww0t5FkGnibMb+sFBiTb+ZF7lPdqbClsaPhYMbTX3ai4swhY6TXUdL6o0lcUzeVu
YgTx6CkTqQNqdyW/0HruDqvCq2e6NrnJ//SDVvZ+qvsu7vooDiEVIvLtjJZT7jTH
tVRUyCvFcgtwLlvbs1of2TqicM3ZxLDk8CKIXKvCKX1fjYwx9B/+fRGw2GTR0tgz
hwoSp8vRVhVP8KHD4o8f3XM3Rx09IRnOizKtrzXaVWGwmbHe5EQmAeU9r6j9ED+i
H/A4KrCwYChetoH2+t25aVExByJZt86s3zElyp9kbJKb63TCv9q5NJM8qCqZsVab
MiUfgvM7HkMxQxyhR6Vhbr8XSRwkpOyXG97OsnKLrO9H+P84X0IyjKQutb2e85di
KzmAQ4946l3v9qLpJsD6sr0UipDyWPBcdk3nQEu4qd1IaRanvrJ+ds5FqKHYlnPx
cdRtOGRX9lY6gUfqJ4FNaGBpQBYxP7hZ1g+EnxhmtMJDk7ritJr7/nCL2C8YbVPP
3uVpCfl23kegwYeemuUDIj/mtUNQUIT7TJozjth+U/0iJa2uWbNEhHmgMWUKI0b+
NXQ9eTE00xks14OPcAHj82j2JK7+PUGAalu/hLSnJT5dSGHN6TtDDZKKfjATVOr9
NYpn0UuS4t3cV/xCcX/OYxoo89STrnYq3cS+Gyge+WS5F+p75zljAeQPQfoTxntT
Oh4+lWfq3rRwDXZWOnBUy4cP3Qyi3tJAezROvm9/wnrEKubMstMn1+xyBGe/J3yo
f5WJs66imLh/8ft2BJVy0Dxd+XMNAZFHywQlSgoJZuqi5dwEbprzgPN9jYNBJjAQ
E8eoFvMpVFCVFljpkdCG5FFS+6Ekv1HKJS28NoBSZDAdA4Bza5h3U9ek9rWJR4GW
e4HxL3PcQHJ/IWxLtMenh8ihkrKQV0iKaQ7cOpeeFz2/o3IK/MfWxK74zB7rLehL
g8tf+XCK4If9Vsx+1vyxLSVY3QLzSN/vns1ur5TUR5yPbhAYizntZjQdGaIaF58k
OYv8qg6lkIfO7eo++p02KuEu+t1EBYts6G4XCZIigMmvv/FrrS4ZVAzWwXCwpDPS
0esfD5I0khq9a0DIzvaPfc9lEhm1BCWAUN3cPVaodtV4QyynlIKqga5zVyDQnru8
OiaLP022QrM27uKvC1Y2Ni+j5bspKQfMHboCl702hp9qjW/jl6kcHgzDNkIl7JBv
6sFRRMNMHatMo7eZzD7rqjVLa6jlAWp+FUpGXM07c5AU2AdXqGSKmVZ6jo1Bp+v9
6IeS0wmgRKxl86vPlc6VDAav4Xl8b8UoEpR3pzyTgTDzYUOsITlcrfp6EqMRsj6Z
WoxGrWifXIrsCRf5mtgI+zHtYvxgO7NR84a0d7z7dTmFyRstbArxpVA8gUEPkkw4
VOw3+wZzz4fgEu9pHrEalHqxQIN+4BtazqOhOlYkg0uB7efp6PLb4F1DOeTl+xbS
t38l4vp8Zr6jgjihndpCRCWU6hMMFr/8BiKr3eWWVAJTKiz9W6PyfSO2VtaezJpi
zbv5cqdFsd5DUND46ktSPNMZawIPukZOWmxoe5ASq/upUw6DxcfInwV1rxnlStsO
VsBymPDl+MdDGDvOx94562FyIXZy3lJ/twQctUVWUiam0O6iwfyi73RWjPCQCXAT
APChK/X5g5h3ZU1udTfGr1LFvrKaXCO2QcnK+iNY39S9bI7jYz/LuvOsHma3bce3
SSi1AhwibDcw+WxFWbwjsjB0h/SukzlbsXrZfLWnR6zt6ZLY+7HwFMNUNFUddur8
c8e6p0uQL2nTsf0S+IJUi1zI1RwSS6/5Af0KdpXfMFqbJcyRc0tuk57Iz4xcRL8q
j7Yp6wR4OfOY9P0Ea6hRBB2VUViV5ExP6d+3HBN0xxuUFCFNx15b92anSXtf05To
H0EHM5UMpOqPLTX5xkqy8X2VG9GW6p5Hg01V0OXypCX6InG8qHS+5h02P1gXLrFE
wxCfaK3uotAxBukfjRAydM67u5ViAUQABzIblsDApD+kvn9W1dZpyWAN9ADq3e2c
gHgSR2oZXm7auTIIytz6XdqQkNiiNZgmtBL6c4cKTaQ19PLx2ZQilsF9DlYQ+k2k
yhbV1HRJXA6PbJohyxlS0n6VA7XQhvVh4SV1qgPBDCDQAeBqYLkdhw2mWsBt7A7l
lk/O5MM0LPJxFeeoubnaJAVAy8EPiBxNvpYh/XFfYirg/JLDbhNgZBDQ7W29rH27
cvQehOB1u9VoV6uD5RZIvqTXCsmIZUeWcPrElILE0Ky/It/eJJdQTqEjjYfhKxeS
zvHk+JoOo/+k77jAk0Pf05442qOJdjSY/KcBKntttLA/1jHAAAR/MwxJRUx2ipzl
B9dcqlSio75UcggkzepoV6J63ScAwyeC5hU5Sb5DJgmvJGMPTDQnHImuOeTgOjur
gl44ceE/vUqiagZie/J1IaGi+E2QfIvxp0w0nWDWG7uOc2Pw5Q0Sh1IQVEOvgD/Q
oihb2fw+YVvTS1KdzH9DZfJA4hOPCWn0oCZZ8eUBXX5RPs4zYM8F4n8A8mtgIcUL
zx/gIliHztGIntfH4hEfZwPE+L8HoVeENfX8RtHCOG4zAz0pa0fTyJVpqDVIUTfG
EBuYE//gH94BlMI5LsTpMmXdNkF2b3fxTUzAWepQIBtAVKNcxRTyu34bBJ7pOOgH
QYhpoJDVGoc8tj8HxInzlaBkDo1VkVC+HaG2QjFzDO2bUnplb602AHXbFnICERgt
9IYitwL7CLCp9yLmcKCwVtmFDA2I/EL94Ji597ry5GrscR8hE8RLTsvc6eRj7T7E
53rNUql3o0rc0RCpPCuuXi0NabtIOxuwfAnXr8gNKPxesCVXUkhxvxooVQhjn6d3
Eo9g3iW5bjAjL7uD6sCwwPMITl+06cShi4h46syAh+0wjmQIsRoUFckQzdWrKUS6
akYrkIYK31yad6olaF9BGTbBIS2oE35kFasXlLtHFWW9vwhIoLF1AzQTVB1bG+2D
DIz5KnLzjVYK/nJNfnitNKFt//bx3KKvcXBWtCi1M4eZS2A9L4us0meRXIaxFr0O
IRXaGWGsXLDySX0CUNKgVYWqZ7U/w0aeQwxrfwX121WGjLAFaZNVCF6ViLmiuS9O
t2awXDllbWYXk9pCsbrN+BeBpuenmV7utYuV3ipKIkml+1q9NvJSweEE6fsB7txm
QzeKjFgdCiPSnZnGTxKoHkO6ol4tGJLXvIMmoDDrwksJ0bJIq+c930wX14iAAW2K
vquA8QL7CSqJsiz27J16aCRPOyYaR4lqEUQTgrgP78etnysLVQtBVOd2e2Or/hs1
DGykzQIN0Egmkkg3Id2JRqDLxC8lJGfGNP3+JsoAo3pzrYfVxE3mtGA2FesVsxiu
BDO8SK14ldO2KBTE1tfoAyXsXBtKbnbU0lVt1WSW2RjrZFpkc/yX8Bd0vl4tnNyn
WbA+QY+UCNaUNSagvjBkj05r0S0NOV46YHx9O5FzUjvpBIwrh+CT5xrZVtg6uZ0u
WixZnoxWU/7JXTgkHul4KG5Q0rPM74Z7AVcwgD8s6M6HSZfhG3MyS0hDSCKrkXE3
V09ZwAj7pPGeUNxQ8/KbY2Lr80fkXogC8FZGrb2we/xNW8ucO4KTkNojIJTAb44K
3eGn2UxpAkh07RZgBlBRwVOUqwPPhQ0CGEwDN8OwdY86X3VkWvs4+dxlbkE2a41N
YuKSu6TyqMaNXURFEnoBsbBzlEzNxFBaezIMekQ2SqNasjHFnHQymx1LBa2gQehe
E2Y+YygngkhRjek72wT+m0cSnhbwVFGkzLbJjj63kzEFvf6EhvcItkgDGJT0qaZe
ea4EnxpuKTWdxSB5MysriaPo0Oa5MPHiU8dvlFXR4xyr/mhAy3fhfWKA/zqvmPXT
1w5kz/VY0Gt3w3OAD9wK9G9yw35sSDw1253rfehstnyXbFqkZx9ROOPk9qc9+RUq
3LnOAtdDWCvT9fY+GruCsgeVyLGH6dTOhpMlgmrOLenECY4IZ6fltXGmfA6KZWDY
DYKavBpj6f4VYF6rKIiiMJHnHhGB0NjJMSqjYmiRl2d/CvpS+X9gw+hNwMesEwQh
+JK7ruw0uZaYPVNpIVxHwpSXhlx/7pPGYL7SmFEStsdOL2yoQbBl4M3WYboj7oGE
MavOgmFjg+xUCHHpJbh/j+1JNmM5cl7Ua2FqdzaZq0FktVTzvLTp6GdDhEe/qTCr
jlq0IT1uZp96be5YBjds1JdRQSZ2e8W05duNeSFKq8q82v3TpMRRlEeuUW60ihy+
KaUZmnQpxJ1sX4k9+68tp4iaog5b7Y/TvbSWkss60aTALpLjleBvrCiCCdTUKkoo
thdFHY1JryTRF1KL+fQULcbK+D2tDYy0bMvLewPhBQWe8WDVRcpy/8MsxlhlT9Xk
GWdOFWqzLePAcIzVrWw056q/9Wc3E4crIIrGC0GpguZwj+f0BnKFZ7m4vxuHTfG9
OXaoEyTkeRlF4dSvrXSGtzA/E/CT54gCjL4qtlIPNdnibOhE0wxzVaOmSLIVTJ3Z
lLaUOtZHMn2Ls0ssm1lJIvnnFhCqPU+kU/cJKLZw8JLufam1XdaE2/5rI/mLybgV
qUWBCpFNrHZ3///2ibLU7s+C58cmyGxDzCnUgeDCdcy1HaXyPgMEJV6VcR3h/Cpj
o1MLGNQwBijbUzkV4FuAQ4WN+ldQrHoIIkWXOVYGglg/4J8ZzhRz7hDyIAdV4rd0
qxFCVrIg/EBbrkRxoJ6KKgawfpt+5khzLthuDK+XXbaL4zo06Fk/x1t7SgB2T0/b
153Vg1I10rXUKEQz9sv4Y/KytMe6J2ZPZSJoIEekViX1ZW6DT/YkZ23AXDXtnRXY
f3tBzFvSeQqzvtQQAgONISfXygsUM8OH9sAcsCCgq+TUoK5aoj8X1D1519hU9exh
MbI8L+VsKhlLp9JYZHNEzqDy6EZzqyz0SBzftLJFs5BHOjjxVRKnPyNJ0/LMzJmT
Lmzpr44iCNaeJve7UCjlWNger6nh6iNM7xe29414UcxsDPRp7MPSrAilYKdr24nz
FQwoZscwv6kKnr6WsZ9akEOZUfOTspjEV71y2+OO40MYVN4RjB0fnPy1d7eE5Z6R
ZwL/cJjngL+MYZ7TVJXWmeJks5/+T4HxgX2nk5nz8wbJkP24QW5wBlqLX/DIGzyw
p2Po6EpS0L40Vz1ySBBpXHULll3MGXjEQDMzomSOE/+zGgI3J2lV5YPEZvyTKhVo
JQ7Z4tZHri2aeRZX4+5qXTa8lz/5GI72zZ48spDWFMGoYSNKGb+f5yFs0OC+HmRH
frGzy/2vQV+ZhynChCJrx9Wp/3hTuFrhAzr1b8zYrFxrwqZObYp0wYAL1s+7bhoa
w4/+n0MZGJ/bnloZjxhuvBkPm/qgHeD8mHb1RPBH0V1sgyySuVGil7hmil9nzV03
R+sZG8V6RZlD6YiN6/D7Qld0t5YwZ3xc1UU1/hhas/tcUKu61axKhfb0O1VJH0yS
fmQmKD6p+icCJgiz5Pl0YSAy+lAJ3NSWDiZlYprEpsUNzgErvohfXhpXf7odSz16
VdZFKCamZRQYDYSVRWGbagd6FqqLA8JGWChQmhuRn+wqSjI6RN5K8xrMjBo5ma74
lvTFSHY4eS8mGO8tUt9QzASzP8Rbt1t25AzQYupXv+/E5uKW1MRJvF0T9iRFzZTw
CD1r3Aasx5bUq2xyFmxBopOxD9BonysDoAIaGRP3MUqRUWQX89DvbyyuSO5ANYiK
m2phnVBWi91LC7XSouS+lyxanGdqcrIwXR1woysGrK2u+9fPtgs61WwmtZa1HuHP
77H4Z9Q6rycMQ0YLAtKOBRAnggpENHGde7hOMYhRMW6T/CfksoFyD0QZRi3+wYyn
gzPPUtNFSJd6gfSrIwUi+LRK8wQe5hjEwN6d2nvIJgx3xgsNODxlsTtULopJlQ5U
iIznHvxBera7F0wo7f9U3tC1NniZqxxBfBWFoehZOAgGz2eLL0YTn3zJ6bW7rf7q
zRjfN9afdx74EyyjUjmE5/BkqN1hR+2b90TW3BavFZl6ontEl8W4GFWOKwKPYTeO
479iEyDTo15czfWl8o5AoqGRqXqpLUW3zXOQVmPn4fv1q5Ynh0uHcdV1fahCRsHw
fBfEXFRkZKGgHQpEFd2IooFAZv/WzGAw69m5GbgtgJziRyDojqnWeLX2+3JeRjAj
rnR8btgnRKGH4FXgcFM1jy0Yk2+JJ3zvELxJppTHOrhmE6uJw39N0XvYH4xAR2Ab
lTZ7GI35EHfXkRCZMeSL3mqVj5E8huP0xqeIWgHs8IRPKX3fFvIoEqNLYI0dbnVp
upRTnabaMy8Qrdy0v9mL4SJlwOgKeAo/WeQPko3VPtYzPSG0LAz/FEkdNnnNWuiu
Ak/mp3wTnqf/CnAKq6aOO/fkIsavk7SYq8JDA05LRocSNpRqLd4oeQz4pdz8WBJ/
cXW8NpWvOVXYBQxvBpjO5W8RovsMxxRZwWplH87UqtHmMkspvzdCmP0tXkPvbw1f
ZEUU6PpaRzYYMdaBIvXA4eOOzsO27XosldpWaoxhkjqQOyhWy3S6RZumLz4unPKH
Trv/ikWyLQ1fqt0u6HDqSxQIda+zSHy7QvipD7G07QcZG6F76xGLI7W2VDkZLTUe
dcVG0VFNlh9QCsGHzYNfQobK8yyujO/YRX1jrK+Ao79tn0iu28vHgA9z+yecyvdq
M1N8wzVB9kRLgEsSyp2eyNH5JC/kXpm0DEN6DBu+wLwnumQ9Vw2v4otjXbLdc7H+
efZhd2izglfLkWoUUmqP5GA92abbSwO4vClL3VUpYNQSHl0D9BNBVGvCXstQkraK
l8oKHi8msfRCA87pgY+kedJX9/V5n3KnHv/TZoD/ggcjl2Zg1mcqjSmcYe/miHiN
LWVpQ6sOBRbp7uxAGmJA/JpwPFtjg22NP3bdiBPMRL9uM57FpEQdI9J1kna+4rdD
ZsJ/fyiQwnHJXKK2EsyjqMNya1F0x6AS4a6U7iQKe9JCvDyVF/tNUUEQQBpsoifm
pXgtMuiMlFblPQfnwYjEIy4ptCK3dUXUWopJMyrcfUGZsBlB9mpknRxoN9FeXHUl
+Sy/xlGSiZf5Cy8Rfe+qgq5l/hBjaBZ3leEm6sM10Z+zVkxZP15+9Z4EFS49La+I
mWFMKaOVcHIzsIpHXI9rp/7s4RBE8w5+qBFxmgNTdbB9rC0GiKWzl4ZA3QVbsUbX
TDJjKGUnCLt1ybUaU0jJME9LR64ZMGn7YGK5zv771QpQYPUcL5alj28XRGHd2C28
w2Dogoz5KzKF3IfUmJhZOJOW6KUQbCgjLqqsjl7VzWItFcGpQjS/fMFp8wGRFERz
KH6hb1YVXeqTnCRyv4ct8fa6C5XurWSw3gd/OlqdO+LYxQINdHqr2b4InW3bdSdf
u12K8kUvqXGGZMmDCMsyIF2IqmR0/6XmWT2zuunaV0poo1weLacOKYcg1gGQs1w3
T2te6OhLLbvfTZac8HW0usn8jO/JUhclI+tgk/masihFVP4CBUUDmbNUn8KT/HC2
OWos9d+ukCJWdAVkf6dYLjrLuc8VV+IPmOCqWsQyy6OZn/jmVJBdNYz3Snv516Qo
Ua1KEoCb94myLYmnxXlQ1yfrQwBJnnMFdFQZOAjjJ1TbLp1SA4QgI1IP2a6ad7HB
HvpT4fKqEo9MMsQxL1QsT6F4dzJlN6NODXp5w58j8i5Fym3mEzN63DCduEtfVYzh
pyMLWsDibBjQiLyenDz/Kh8RLkh3Ahh0GXSiZCsd/pLNB+DiazZA+K4X1CXjR2CV
xKUl9pV8LMIXq7c7JL5aY2Moczs/qqMs6xCrJT6IXboMeHAzvvGIiteUbgUp2vgB
2fMLdh48MQoUjobcb4kEkfDV0JCXyCgtTfbmzKDUYyv66DFW3ntFF7BFgWFB0Nao
s5u7Fr8Kp0noK7RWB+VRlOU5Kwkj+H+/gzdbBn68ZfIcWYTv6vPasWj0I63H7+Ab
T94C+rn9AY5O5vP8pWQt/S8X739qsq2ssYKtbp6A6Rr0fmNnSRAzQj2UGSWRw5jP
pcbdOiRtCiTWNvZLnHjoAdq8iMEurcpYqbgMti1Q17cF9q7Qt2wVvbos6t4yNpli
N1CqrtRWc3RFglKDvtXbnPK//Jvwd+IOmcJw+AEj3iIUo72A/m89iGd4dRdtf2p9
VL/FeYW9doHgxVtjRq16h02cbUn/JhiRlerbxIshKEsKEdJoZj2w6y+/tZqoytCc
e/axqWiU3vjv6q0MBYvJ21YZ2l9Q4xAgLSnBSeQhfo2+KY+DZ0Nzcl15zaBc5S86
3cPQIguqDMtRfz6IxHDej4LIMLlgo5fMimtIKSt8g7l3Xvv7KV8L/NMmISWO+9RI
ciKZi+kiuIB+c4TNxGYx4UfSiAtfh6AdGm7ybp7/rm5eMDoLYqv1dYXTBxppJuhU
ZjLm7b6pFlsqK5AKG10y6AC/Dg5a6EibMiz30daQUWJC+yesScYMMqR3KWYNRjsi
vTpWT27f1pL7GaAGud2N+5i2xvRNlMOIdh5L/IW09jrjKqbz9nts659PgRGWdr9u
Qc2QJdPAjRnwobbfxEtlUw7mmg65feUmkcOagDfzC53crrd8M3+UszZS2KA7Gu+d
fuKxicTHpk1x4byzo3NcSSzr6yia5AVSlHRZD1KW/RbHB350PzWytG/AARGu/W7I
nAyoLC1f7Ac4mLbiC0otnZkbD+6aaMA4e3CI8GP2Nj6xJ8wnARcMyGI/RG2GJw/8
EsB4S/hrzlYWYLAyts8gUOpVbAQPQbYKwf2tGu0ZjNO1Hz8NBwOsoE72AR7rjvr8
/IyGvBRus9uEdQlB7e1HbHACD8DdC6LrZThK4j9hS/Wk0zlb7srN8wyUD2ne/pzm
18Pv5w5hZE45tvSJghuzsp+8U9zsTeQEh1jd6XGjq/WdlPSs+5L5AW7IYSApuNG1
h8tPQpcT4QM6u2U3gaV7DPUz4/UBrqmYKYqS26wOOtysL2Bk/vq5cTU3Y31A2o7I
iL+3QE0BAFSBly78GtZqpbC2tsZCOnCzBVLSNLDrgFiKWSSim56Y/MXPGYwhKtFG
i2Sb1MmygMnenftiPOEmeW9qhqygyyJsU4IZbKdZBwMGxLP7iGSoKgk3cotqawx3
Sw7YkF1yPt1zzuviiV9UZ2EQBH3qUr8Op08BRXmxZFIu13T6T93UQiQJ09mtHwpl
DJ/OuUeHM2DoxzN757qt7VMPm1YxUrm2AaXbgmDQ+dSHfjf9F1lOyfC3so/1/RY5
ZvjZUjEKH3ZaDYejiCh7fBkVAyttUPS0DJ3a2mw2Rx4l1sTVNmKAkmrwr+4QoS5c
eY2xOKgjfCaJIgBjkamSUQKh/mPLi9rXX7bsorsaxcGiBzCcgAzAzZ4BkP9nlfEy
1YbJt6Lqz15XaFKyRCTu5DntQW8xGqDK06JbGi7epDVfLQ0ysgmMF19lazxELjA8
YccviHuOGTyKpqgJVPrkYqjxX5Gx2yDHedckCO+RzYGnlLaNdQxs9OPV5Rjwi+Qa
uUdCOJX5v8F9WRwOklHbzDdFrVnevoGtB0hkIKVrVZK0oAlJXyh/rpuxm13UTg2Y
gnTW0WQb09QsIZ+ger3UFjQs1Z+qOQu7NIFuO1fmwIfRE+/86E8SuLCk+He4gKKv
tEPrko7VbOBJi29QMwet+DDkIJWEEOsCX6abP5Qc6pU3D0JIu53O5voaW2nOB6QS
8xK7kDCYzs5Hd2eOfdltyFNY06+frluoMY5Qu5cgtI7G5g5unTDIrHTaCNChKNeh
ELIB79PQO3bXj20FYYoowxVfsbj5f9yQCAGjKGBMyzc+2zgjwLY/fDpb9k1yQbya
wAc2W15PdYzuRwXKRkngpHs3vglSdzm61KcuDbPljEJvWsne+UvH3KAZMMCp2PsD
Aehw+8XyfdQWTzKc5g5OKaAeDLXEJTW2G5rlpyGplV8aESqxQtSpRtm0+FwRsHRQ
nn4ELTzDg136GHyKh9exFdxSSMQnt3+XjxvxtFLoihqmH8x3vH0WxUdjyV2Ssh1R
U1gO3HOtBYq2a/vM6zwR7+1Vm/H7fj8T7ni1FzM9X444ZOQ9hmMR1nfNHG0xXX0n
uYPLRQMag9KVHwK3w83kosx1Yr4v0MFqaYRrZfY/2STtSLsUVmFigF1vZ2bFDq1o
3NzmGWUJAj8Y6XKVlrLd9NATk98xz8dUGApn9FND9bA/VcRUeeHvH0a7TkwBszJI
6HJt7waiWqd8xKbc+5l4E1ZDVUi4Q8c3Nyy/YhcsrUqu84jyArzugWlVEYxuK6kB
5OW9ALvVz+14vQxvBhXe4JvMCWChDcjbq+YuADpsRYZ4xxKt99CgmGw+r1RLwjTv
kze5EO+v0mvJ8QTpg0AOsGl9nETJUDYWYIgdYe8/qLtFaGYUzdQ6K79Jm7DtdQXO
SKZGyN9uIZrZV4xkMUQZSSBhJlQdh+XDJx/O/v4059vsTZ+tU3YEjdreTA2XGZ+D
Mc1s/c4Kv33lhCGz6dB4FiDhYS/rgUylvEVCqHG+kde8SF7z1l7JYKULAYNwTGiM
0VDQr5N4Ul/WIGIfMRdeCPJ+z9unFgmcKwIe4GV8i1JkhlRO/Agub9lgXggrY+sy
DSr/jUrplr0+jA+fu5Xnlu+1Nc7Bf1J675kIb3U6M0d6WXKfDMHCpEarQVqADjQK
L0kQZ44wsKyxwKvepbXRSZ/dXT5o4wxh10OqM97fzL/PGs/bIkHExE5/Zb/Q5Ij1
1kNjyL4nPZSctu86XoS4qk+lw+nE3qetfiDT3qcp6o7DaFdxvi6KLA2NEa8Y9Fj1
cBsbhpD742kPsK/hGZYS4iHwX6v2Gv8ufznCRcnqGqsQFsvBctJCy/s2ihYR7wcS
D28xQSv7xdZYYMoNCOARuzIQ+cu3g2hYExTn1HmV4QrsAcyrbmekfxAjyk6A974X
qzWJPw8Cq/M7+HY2EQbCMdlXNd7aap/F5AVJHqElw/R0Cj6X5unHU8pr/62otSFt
3jY4LCFiXx8WG0Zjs2gJaux2fQPbk72YJckIEwqbjfDCJN+QW47binUWMh6EkzRB
6lK0F8Qo6gVyzj5pEtlLcVnCn5kLOOb6+GfM2W7kxFG+rZFIpMuTcTq47OHdJRRv
vS2XKV6MODyG1tx6hHRVI1+S3lW8o1oCWQR4kSpdrAMjJyEYSmUSAi+4mqtHfP09
I2akv8V1UspHN6bIjnvkaklNM5JQTnhrBEIQ6ige7fY/4NfLW7G5jlVRg9Jflfoq
RddUEDK+ByryFMon7POsxJaYk2233YKlvK2bMXD49rLv+CzHRfi2C3AroNCwIjWs
hfD2Vn97foIgKd8rL03zN5d9jzea/4xzhrkeLTdJnHK3BnrDOIf3o2u/A8ZpHbeb
amAUnl6uHwS0+1ANzVigrwgtoTNmziIc5PTTBpsK9HzDqYYwCi5V8wY7YMfRZ0SB
pCbg7ch7nkj0N3op6G/9gm3uYysYtHNz7f4nPXd0zDPsideVrINajRmKuwAjGL64
rwNReZ2tk30CxibRpTCMSd5pDDwvqBJHwotqWnNu8qtnZ8U6zyXGUOOMYFxEhQr3
F+xT7xKLgAuOarH0Z1zxb1bzdA/voDQNkIZNRGUtQj/gLM30oQlNa385K7fntXe9
vS0Wt2ER0vKCy/hKmk1YU3uyb56V/EKfx2kMJ/SPr2K/OaEuIgx76tn25zqV3JKp
9XbvACdSgTGyaJMHjqlRLqI4ASMkIIP2pwITVOsCxdO4Sw9ZFQ5qmT8BAd3166BR
nwq2MQkjyqt9QrzViX7LN7r+4udTWgSGaheSTB+qv7HLSeNr9ms9rwSnxlVpLCPz
Ney8kXQ1zZvuez2l/GlvfSQ1jt3AZ9c/KNsr0CydNQsj21JIYlx0P7MQWihAIvd0
bvIKmhw3LFc/VCetM8Lrb74QlV7K62HXuswlO34vOxxIQQ1dSb+p4J2cmHgCNV6i
oCDSYXyCUVLISNYswpa7UqXpCDfcXoAaPU8uRurEuask5r5dI0RAsG1lO8BqKL8/
KSNjvGDFjMd1wnqVKy63cE/8kKqrz8sXcU04zJTzp5eoUZ6Z6iyB/f6dbcBd5YAa
0baJs0hYaemLAMLZ1VneVoLKRqDMwSz/EMoiKWOPz5z5a5Gu/yoKwaLZedUZCYbv
rgxJls54IMqdWbzY25LLxd7faG09TMLrXkuvACwzhOHm4SDpISCgQIka8Mhb4giQ
oZWPaE5lWL2+nR2a0ZHLgK1HsEFxiV3Vdm9w/Lv0rLunAJrbQEGWHi30tnR4NA3a
E3zYlIoLPAreuJZCBcvW+d7IIaoWHjYa8myGRkntfJPYCVfxTteEjReSJP0DRWnR
MULi0EP8CPu0gkdmxgK2yjXxAhLv/j6yHmv/RoVs+86R4zcLDrFtDFPtOsVd8gLV
qFKhDIJByLFmE6dwsgw1pNCG6gDd+DKVFp1iXCQ1c6DVQ5EP5laKn62wAnFYBRIi
qegbt2RYtN6VzGO4sv/78Bkil6x9qZayLTdJXqPM5dIekEEJJvornvspPx9LRZsO
DlKDWJTgVEkg5rYHFVQq1M4CmxJH941eOTcuYI2cWembh2tckZESeTL2mIESVP+F
zPD5iFaQPsxmPLTH4YALXW4vW4uj2XkYIqxNtpgUCZcB108cGur0sILGXP9n3u6w
5wx1kGWXPpnEiyedbHxb7I9JYNZs6ERqcNTkgdDLmvnVRny6kvt6gosC58NokJju
LmhuMuMJBVj6/V+iyA89HfEQfGKZq9vxjBkK+PmsFtx9GPJVMQsnXn+NtdoLCvMf
P2i4XezGmGMei/PoL941a6Vh8s1ZDj57eikRUSErViJWEJiaUUGj+Jlphu7NuaFr
1Za7rt712UBAu5NXNhbS21P3XyIBwO/RTlZ3DonnaU7OqjpxQ0NFGV/Sz2dREEHF
wOmtFPg+GNMNFjRnwfdfXGeUajFlZEZR0gxMFrud2q+yVmkV6SWjgJWbBmfwYVOa
B6W1O4tBGeWQAydwfJjJJMXtv52S2Sb8ydVfSNHNojpYRq0K8gx+8Za6JA4vbYxg
azbB5bCgSu/80YekUjHH1XHoVQxaTI7V9LLe8CWUE/fquVnjS/UC3QQaUFxlq4k+
/7Ra8TMLQZvwbWQCMIlFzHgSabpL7YbclPMykBtYLfSTkZRLiiQj3Rnpk2uD5zCF
KWB7DojzJDqo0gIXCWXm+iW+wEjuDWsMJIKeGAzmaHGOzxKABkgQC/bH81rysoKn
kKK84vBVxntFGYoK+US1VPzmKNegMosfxPZF1VPEV7b2bvv3HpJueE5iqo8Bf7KH
sjJOgs75/P7MEnQ08FxKVRU3PGogWDiQUIc5x/EcotCw4J0Nok6KwzMOApJ1HjEe
xwVpzli4wB2RrDDsQpUB3gkI5KF11JKMEnKLFZnCh62pWiHoiYRZ4JFzkAmpVZc+
ePp1CjZq51Kjd9pze22C95jgHx5JjbR8iCiZlqzeKYJIQyPzNYXFksOnIUeE8zyM
fh+r+SDmXgX3WH1AWI8V2TMUDiOAunoWVUv8XxoglmRCSqwG/dp4g9YlF4h+extH
ia5c7q/F8Fs39NAjoadBiWtV/SEvljWyl2rtTms/SSlQ59GojdNMvCRSnW2WF7k8
moQeoFUFKRO9wRbU8tdwVhCpsYwKnqsvVcruIHch44SkCRKrzriPjpuXn7EaaGSw
uQdEzqahpL4R2oJox3XHbxqlvXW3+eWHSvbc+NxbjwlP+VnWIQpSOEQCgi5wUGzj
L1bh1Dpb/D59M0urVw7ooW2tYDozIfAZGGQKt0ayuKMZGTMLRnx32LaMztnLIabp
4sFqBDZTedVQd/MD8TO1zYPnUo83c8zEpKq+yBLUSpMxjYafQtIqLfbRnHWILzAF
KuFd6YvnapRiggy964NYqIAR7sQrXTcDIo/a1ycxl5x7nZ8IBtwyIUMXungBYq2f
762BoQoluzFdl5SsC34ammB5BC1QUDY027lkrkjsnYY5PVMAw0VAJlBP3QlkIoI9
LH03pZwpLtvaxFc/CapwNu6nWC1I4VqZazoNl6BUpKN7CeGBKQZBZt6EDMJQxAE7
3PKbl7cuJ4wbpMtzXbtjIrUsQAWj5AqmIif/lOVGxiiNp/mzJoR+juPZx3Uev5av
YauazVq0CP4Zgz16WBj7eWY6+IOGZIYqvHuCXFLgu1jo74cjq/cj3lxPQ/C9ceKJ
rcvv59KrbvKcI4lmJHu4dFUz+s1ZX3+9r6xMEqsmuD1rBGpnD9HVFBiE6UrLE/0D
gwW9QAzUeDQJzkGC80j1j8I+MoFYvIVZq2rEQjSNlclmMCgWcrVUohh7YWbsGevc
VPurlogIVnu5Uu9QnLsVFGAzp0S7uK3F4s8ox/VbxM9FrXdio47/MXs2Esbp4LiP
jNHK+FBkXrV0EfLjD94xZfE5zzw13M5NK9V4AYnd4Qcl6q6K5x2OsILaQRRHxKA2
R8yjo+u093x7X4oD+HTuXwWDm7SIeE/mDcg1+3nR/iCEahgXA2QRD+buT4L09xy4
M1aViXnBnIAZjM8JBUHDukRpssewCn8tL/AFtc3vtk7Tp0xiKq/U8ogmgHuhg0/9
7BKWEsPWWCgzuqGiQn4B+68UhEKfL7cSArJICUxN5iwF9pirqInJ0giK3I30/vg2
oIFq4DcwIgJSgp8CeIbgUrz3rSFQE/oqh4WewFEoZ5rHo5xmOMKyJgeyA7yg0rRr
dcc5nCpKTWfEv3OXnX6SDIROIP84u3H0uTw+EM8SWHjlrEOMD0EyV4qW0nCV7ADw
8yTStBp0ceywerWZPfE9cafZXZ1zi7YpXODET1UJSEZzRr4ZUT0ij25YDYTzZefV
OfQAPLDcYQkYcwAA2idkwyzpCbPKgACm9/13ts4VA36laNnRnN5Y1KTY3MXlKqI9
gvncE49HYg3sW7Dy1sybXlbDmbtRFEAxRGUcG8wvjbZY893zoNNsmcjYIoTHJRY3
2rfn3OAvaRsSGDFzDSJ9nbQFcZ7YxrDZvqZOFsXtBpgWG4PQ2e2luOa+o0APlVRC
kSuJ61CtrXdumhMrCK7CpnGXeh557FbBKRz4ri2tw6EEPnq2NRqj2GvfcbuEGV5q
ivQoPP2GaQJPf+RrPyJx2K2qvYbKMOF4Boxs9PZ49uUc82fFOt1cUiqjwp68CX1f
VCP9gDcPdnu6K4fV42v5MJuKrNBz/JhrfaCwOhHHKxH9D0UvULambrs2utTfVdAh
2TyllR+DrSKBBx6J7KNRTSN/csnyBttbTC4InPnTNjZBCrtP2FgFdDDZu2PFc6/8
/dAwsjylG8SZsLC3XyhHXoHex8dEUrzMyzaSs8fdjaCBwwPwTN9wav6kxe2Xi2Ek
6lf7SA4TepXvUwN3AiKJ1NUmypQb+yXFhCldgfx4ana3DnPR/geCBrd45Ijdr/qC
aCiiSAMqzpVR7h6CEt4xBfW8DphzAyulsQtStU4DTigEPKHXzyhDwYkwL5rWDGHP
+kmEUReSSfUOL+wUQJC435W7DkUB6cJKFL/vnS4X/m/9A40458nHmm6gNHPyPV6B
FDZG/3p89m1umAE41vtXYIiMqykPaxqjfNzzM3iU7FvSBSAib7EkUF1GAyivkG4O
djcR+bEzNJ4vSbR36jQh9+c9Mn/g7glQ12LbNk97fZnQUgHgJx8STaCJ/Ruw73cI
8QKle+DNZzPhRWSU4/0XR22P8+QNDP2Wj7XjOfnIv4USRUEcceYoToOkDQ8uD7CD
LdPx1w4fa7NIi6ZFEGwfkuUA66gLo6EISMUlXl5HMRx9nUCeMtQXnYNQJqGf9cFP
Yxg5hrzbwbVz7P+4cHXvaz8FqX6Fj7vk5imuAuutC6AcfoNhZGNDHGp8tGEhmT3W
g7rLDtfA7L/kZY2ReZ4GolX+mnnFVK1GQXs3HKEjiPnXTS3l4BQ2akKA+exotazp
ScP5WnYwTSJZKAvGZxF0wm5XijOcF9Do6VjYP7U2ysvGcmsztiXfFjyp4poyBln9
+PZZtMHDKzUdJPEwsIQCfrIFy7JUFf9XekD6ZyRmmpgNeFkUg6k0EMlrZWh77sxM
nzPh+Z0o+65zzJ0BjgU50M1dXUlRRkkUcYBv1RAbc+qHFC+PhISb4Ouy0BbmWRRe
LTUA9ibdOisTeYENbqMvwb/KV3XNADzYxQ+BMXEhcffSuiGT0JzjwGxeRbyimBCr
mOPJcFQ/adT8Nv5HwBwQlGsW8o6nFIJDw8qjbDfpd/8zCXvb1ZuyAmy/UCCdfgPh
UplUugMB6EgAsoycR+qm19LpLcjr8iKS7OSRDq7NlEtGF7uecYtKg9+aTDWta291
mB47r2LiOkUQHHleBKyDeWjUFDA7IFFUtpYwtBAPq5fIrrGp4ny333Mp3muex49G
9Z3asJoNac3goBefQR+7ihbR+PIVXJI2Lvdq4fHQtRpDnkGxxZ/LEIBNtr4s9zR5
4DfF8v0W5SScMIAEIbDQlZpU+4yjbrV+f+ulabH33yOCJzjg7MaQXvc7hQO7+2Ni
mYOvuF9eEpzD7vKvEsFMKZDrZGo3z/Oyl/evJBcSSkXdMMVEMahUQ8g68LzHwkLb
roKbCwjOOCaDyl1ELHYU9ptnJdKbZW3crjcr0HTA2FpMivbD0GQXYVbp+h64FM04
zY8EaSXOglg3y5/coeFq9H0UhBzOH7ksTaLyNon9SWyGvMVFYZ5+Hk9r3CYS7aGB
fuMrESxQnK2pwxkvNxUQyl9648Ep7ZN7qa72uELJyY2BsebPHimRwVd+PBHctHLQ
aRmuR/XoVQJU3TNQhMBaxBWY4nQ4BZGnI9KXsYpxGH0rrD2lr1sCsfDWNSUHilpm
KL0hnkbyMdpVl3S9k5A2ipcf62nqGzgtSCMJFKfiF2FTIhdp6pdAMc4OIUoyTOM8
sZzgqqEmJUAy8+U14hjN8GQqfoZiuX9s2NfeskbLz1VE5Pa68lLUrFkkPiHANyxo
5x+b4zhFQs2y6bphlr4hlykMWwq/CQUdvNUiyjinccY98XYplzHdzMlTkxruj3dN
NUpfVHRgVos0t3TWb9ZVKfrDvEG5w6yux67Avght9Z/3MBfTQUByjg66BL0qLclp
hc4wWq6V+JG45W9TO+BQ3BhtuYyz0xYcvUcwrgNZwqv5HkKMqHbbUprNmlzRH6Yb
xSGvZuNlxX0GM0rEW4A4Uqu7rNUX8JlduTywtYJbWP2V5ut5Nj0Ldw6ug2VqBjFs
FWRqOhdePdsUelFY/tHUEsRzEY9biMA9j4dR9PG9oXnJrlHO329EJ9PrMgooGZ/u
1LSJvsckdR2PI6YpbQwYF2z8TFd54C4umoajqFtalHjyRdXd1Cunr6bHOUlAkTtV
9JIsk6u0gHZdOzFnc/ZQXG65kpa9ioO34CPTRootPwh6E9wKtnasMzsYmb105krC
YsFZaB4fiIf+hmbXCLrjZ+CScPEjr9k90OteTzNAOjMsaFlVPOT92JWrsyzrbLCQ
55AhlbyQXo8+q++LPWZbeeheadZdhX+dGsXObqCMahRlNu+mow+HrYPNvZmK3HaO
M+FCx195UJ0xONB0rMZKyrh9/brCapg3u+ObNGSsarmoWaTLzXIUU1Jl0tddAhxl
5BZBC+KdKZCbgkZDcJu2LcnvPOgabquRlWBDBjUJuxHCl+uhzdSUZTNrNP2XygpS
pkKUnNP7qx7QR00gHWtLZo/EiTbYqdHjoxP53fwhsZRcsQTCmjrRV+3GfNETpUsN
iM/BNbUKRoJCRhMEBrLOSYP6nv24+Man0f7XIU9cbhkwny0670ZvEWEKCLT2qVaY
imPy2BSG83CzV0rdXKP8xPPsC2CK3GBSiGCYaE4iWdMi6yK4vlcBwgdyYO8JbL7Q
ZESRHQL5hhQxULnqbMZKPAsY1rBgTsefheJJUN9eORJ/kimHKQ4uP5xabFp6/Url
IG+j489PmGvrb+Y1EnVXenm7/e6vqGurlqR8zcKslQ5aJIJnfeo8L0g5nflRMSDQ
BeYkxOtwqZ5wGWSn75f4CQ2/cKCCHFZmLTa+85G8+CnjUnHY0prJDYE64FSrJ5Cw
aZLaQtlbS8lop3y3myW7coVRebeIRqGLuRUWvnBKIE6QY0LknNi8AedB9+52ZhZy
RweC5YsL79hSLQABFhGgxYgF8N224blv0HGzqlt2sjs3ABw8vI7CeuG7ivcZFo9h
Ny6c2NCvMc+OCVDW2IPLRoGo/DXS/WCOOOmeNBCCl7ZkslNpR+XqcqcN4jV3nNN9
YnCye2yP+dUx3eaik2gv5qiwjKFVbFehuDHIAKUKYlp98rpUb7GvluUkklIYTvtp
ivHlDpWbiVu8yeYiWkx8XE1wPO1IQk2ekF+ovAErUGVwTDTWL/j4DBcTlodQiiFS
2LE88Bb0SCiR30N4fQ/zVmY9n4RaUUHmmiAARvuY3QPa/qwTXGAsr3sSs7Nt1oMC
uW2LPunpqAW/VOtV4RpGFH14cfHf12zbAyDwsJanHkMWNZcbov6ZvkDVHJMBjg8X
MMZNJx1LukVhyCUGAe+QtprJrxYL+5HBr5izRL4+DVhH1gGvsxsZigtTwtMNZYTJ
QjAengM7J4WIqp0fwGCTOwEPqh+zj3weSzpLSlgS9ZwTwg0XLxtU09vhpm3iz/Ih
F4RyvO3kGOwSUxKP8OQBzWWOIjwZJB19gRZRo+ZuMFPsp8Ysygzd7uHnavBzQTNn
GrV5LO3JbtXEgEG1yYnA/huQpnstZB+0Lhp8gddSNnEvLxneLA3wfWorkqUOK3cH
OovERVFMbFxK2NKKuup4iWMdhsqxbQimG7Dtk2CGa/gh8OEB5mijBakpvSmQRicQ
Gvrs/HslA7odCOicP75swDNQa3Kw/R8ym7638BuGMHhKGf2VCkNST7MdUv2Th8/S
4GVta9c1pddfUa5hU5XObeH3joBfBNJD5uMeVqMafw2iqjdc5SkQIzPtQp9AOumx
FQ24bB7JkT3/dnhrYYmBYu1hlNPi0cLBQpZ9NHEb5tNDuG6ke46V0vJN3OuX46er
jqPHUpi9JtjEs8oIhiLWlOcF67GniH7zsBxD474US6y1XC7zoXKyA3btrhG6U5iB
2CEDnKL/fFKfY0kgUhLKT3EchqipFZw59vYzSHUeuXblFRKmMMq6WhmBmXZXq5tu
duhxoFXIPUPvlq5gmRM+N/v9OrqFrIp3TCFEDmK60N3ghtxe2jA8Y96PHQ8XN0wB
66c31OeWVIEndLw01ilcPe2b8h6o+xIz0o+Ig+K6xuVusd/lC2e6ZmU+apH+YeJm
FpJ+9Gsi3PaygnpTLBBkN/NPitbjXWwpxoqjo6ezTAHuQe6CxW/budNxOB8vtthX
ydqZh5qPCZdZ4WSz4Ng86WGEz4TXGRhcEoHSdi6EXxvE+83fBDquuzEEejObp32z
wZ2vefSkm8uV/HudPaWAh9c+YrVxhvpShvG3ig0RGKYrtxlbWhVhQ0LVtWFt05fo
qkUljpvIiSqMG6UZQ7C/E4ZOzUrSuPeW0VPE0YxLFnyTOBiX5YGx/ZFUd8ABKyX9
Wj15tau5/lx5+tG8vUuI2S1mBIAIXA+pTp1Vbz/NUCGWJALu/yjkADMFOAwHr5uw
2uhwlG9lJUauTJkXAHPL+zYk1ZY4jCGpe8/3aIov/FO/FZpzZ/WlpZd2hX0PjxSQ
fXuykV/DyS2guyL240cim2iBw/GXrFQMOuC8XKlQNBJl4UpBhra6JcYjKc1qSqjG
+z+M3UguCITngEXDc7P7oIyMawHgu/ML5hICtDVawzhcvxcl6oLHZPLO8pSlOEvL
Ln+286Fk1PfcawzkZJ16kvW2q94fvuQruBp0jCrtJRkhhPq/1++AFAjnX1WtPDd3
BC00D0HuxpSyUrliH3q0EeDTo/VulkmwbkUeyKUao7V+5i7g/vlvs8o7l1QgGWq0
NAuvgaNquQUAFLuezTdvxzR8hvhbdN2hgDGsraD/VTTiRNFNz9m//05cG+ORG3xW
8HYHuvpkWm7MYX527EBZSinsjt9AnExA/HcGd3WzI1zPaMhWJI8uuJ6EwVRUpuKn
ekhTJCX6IUuyfJYDCZEmMX0EpsYjYmDI9nC71eHDCxJXzgeIRXjhoLIBEf9Gnk3p
fbEZjA6tdqnBqXlAm/DlU+HBFxg6KBqFPonqcqtngb2uF9GvEC4fqKFWTwNyvR6L
xQEg0LRiNa02RMTA4KzD9u2o96wU1IbtJ/WhBhkJnPaNLYeSMEwmfX48qnEIEem3
Rg196KG6J1SkBnBN0trTckaTg8zT8vrf5HZDMK9cyhIa6/UDnEEPpCl+Y8HsEvds
6SOO2t7FKIARFiapZ6krLHZLsbawKUbfQYE4/9I4OlcXzPEzbGx/eWeY/CDspDRo
EPacimNRm7i4iu+q7/5SAXo0VvAIKoTDafuwQWPmW5SP64l57f/ipjzh223djpa+
Ac5a/ydTIy2+VgxGyYGY2kcnCqOPvbLgYZ43DX4vRKXNL6BoqdMqXRVL7fJcUYv9
R7VGH2k4rL4m4NNjzxszdtJFYK/fE6wYPsX1lFC1WcfLkdoynKzRcIJHTYnUvBZH
QpX55CJfTHNUrXl7fDLiuXqpt1PKp9xjsebD9aVEjXyu4kJN1koDIRZEsf0v4mQ4
gTNN/GoX2fH4o2eCU5DJs3bbz4lLf03+XfbrxYzbec2jvs6VIU7vM4Y/gsPQ3b6O
E4I6U7ExyvMwkFxnjEBGr9176pkm0YAFEr2JWWBIsON+PUJwuTqM3J5xIbNE/8+h
/JbnRZs9TjYt0XEwY3IWhT/vPR52QmyBiBvV7mbIH4NxRm13L+MglEM6sZ1jTweQ
lHXXIOT09dh9CZTICDWjcFDXDq1TcnjFw7Yw3RMjR33T0dikW2rFqB2SW06xM8cE
CFDWbFpCoLYGJKytfItTop+cbgGTPv9oqxlvC7kQf7+lEpEwhKjIyvJnO3gM98f5
qQCbKT/ihmQ/MMnPe2qboru+ur860iTQapGhUYCE47bqWr0+WgF9le7YlpO2JDlw
vLR0v6pq4PNd7YPgR3+49y40bNOpJL2Vi7BMzgFyJV/dGghj/dCINxqmen38gxOR
6DqVLhoyCL+bzpkKKVuZSNPyKQZBZ5/905KEoQW+mDhTcjXz0FylajeoRaLUTZ9b
/piQEbmstBhUQGfZde0419XVCifLsUFeGb3k/cwzhDaIpdwtlJZ5AjPjwYZTEgJg
13+rArsRUgXKtL3cEYP9qmrQYpzjsHyJJczKPk7bgZpeO2u89b5szo+3xL3MoMj1
K2k17T/5RzquU/1WCCjBzsEJ7qrfFakylmaAYMltvE3dBNX19xHQT6yo+eNA1J+u
8J3tRPbWKSYeMMP6xqB/Ebzaj92uTcfXRLU0YOsdngU8BOAmzrXcxzxwSCQKWPSm
LV8NaVOeGhtHJPgPzjpYGtM1DK/ttPZ0a8LwYIS4PK9d6M/N2xUYOiKiwZPC01gh
bqfMYhk+1z79OwbV67SgnGVDEkmHFseC5aSGSlmsZyah81eTSuoYYUB9N/SbfCJS
I1m3068kyecOFT/AKGLVoeg8ohBFgCu7a/Q0c0TJSZv2YWtroL4IkVyVhS7GnEm0
Ldk4Ap2ZIzL6WAwY/Xp13A9KL0NTtiaKsln1Z+qyrr2/EWiktVp+XbOmGtEPSP6I
UOjhJuYd4tkcqTIRXK7++XKBe56p/eQadpGlJyuDo+W0NiuBKgci3PKEGGzGmLWS
Rf9OrAwbFJSRXZSMycxZvfsV8rBqVWrjufRlqVi9DE3eulgHT0np/wqiTIrxwaNd
7sk4RRBSPtCFFAr+OC7uen6Ra66OtvetqdYB6j0CrqRDGqOpehKv96/Q5usAYC/A
ULSKcvOLY0B278oSRPm7cZfUpWH8vyQj1/uYehtF8fECZGyXXEfJ4fycCMWu0Hl6
nTsfbVVENuadYltl/byHQl+d4akzq8CLdiz8arXzkw769LgCsDfUvskLW4xzKi/L
OEbRzWV9Tvy3dLilFjj1kVlMRXfYh/HvPvFEH5sOiFuLO+hVWAhADubLRXd82XC9
IsRqYdtGru2xCJQwi9rSX5HszCM/F1UPP+66igWmAtnbRh2/SCu1vBYutJMdPTdg
T7yB37mHfNy4rVpUvBP84muYYah4PnFtB+aK+/+ZPYhtochxlqAVa0TpT4MgO4Qu
fzj1Nf61PiEoVGm5n1dUKsI+VgzzbrDNc/qwdVlvpq3/r27VWaDUTfCr3mFB70dV
CNbzpDY/TmXx1BxS1T0lslJ2B1KEIC1M9qVBw9Eg3GWUIJOnPxs21uij8dbYYpsv
mwI3c9gexLkyUvnaZxfIDKAXRe3wHk7vLfoKrnErDLteravbWSS/mCEEiUOPegn9
+pqY+aTqbsEPUgXz3CKpm9uNcD4K0FS0V/AKIaT/6CBRpfg9aMoMK0nplvg5BIzo
o7gibZLmL9rgky8gLOBumuCEG+MTA8Ay/OE5ssQiyWz9jQEeOGk/9EUDg/CMxUmB
QMjqw/APG1UqW8b12TG5r9rOFPGZNCIfX7G0/LdFhfMR7MOXVaETTMOrNi/Y/Df9
evk1A0ipwHA7y38yGBmFSI9pya0+mgaYWtOOlKHioTKsPQ1/vP5NK9/fLjgIb3EV
GoiHH4iCH6bGX1P9Rip9xymkIZPTq4+iY85MLXid0nx8ck3ueTpKsP7Z7CyIqDK6
HSP9ThVFpRjUwXZk/5EUUf+9xd/3/0HA6X9vDM+DzCruKmnLODtpaCmcRvaabx6D
jT3UfcnHM8hPtoBiTsVmbk1N2v+SwE4n/uBqhc/wwlZ4O+qwyubDkD7wQGiHZRtq
MS6pYFvw9Ji5vN8p8qHxCfjfEAsxpA+5SbldhOva5Nk3ucwef+b+xANBFkVTBcGA
1+tjlgQCCkhxozMPtPba/MLbrG5+aK4sO7tcohDfjQwbiSmM3rtC88vz0Nfu/kKf
aRxLQEo9SQPPHpe/X7gqiLCicGD2fmWoVDCC4MYMQWNL2obvUO4pfjXvM9dmxvSk
LmbTNFYhHhHwG3/fCteIgA4NXqUz3+nnxOTxp7WDu7vxA/4FVv5adSXJ2MuxFZT3
eNQ/jMhiHuX4g/bdcS6tj63o+37Xe2QF6ARNeVPkFoSayPqGijwLYx0kAZ3USkB1
SHH+1ci7NsgcddvGZNKsSrAZKHPF+6ffIuxHabwBbHyMT/v3a5jYF7iAqvmRV3j2
A09AGedaPsQ+2gdHgcNj8/dfThTCkZHkms6iaaiFhwXvmZQNVIuY0AgTG3avc0ih
OcJJiQEwjtVepZYYxxSsL7KCpfs3Fg5TCp466+cvLf1sjgFAiyVdQdh0WQryrc1O
Q+zUsOSJAkK81Z8QDd87XtDid4X5PO9lH1QtiEYb1lnwMvrk0j3Cqdj/fdHVyt8B
nn7+fP3mb+8tLAh3n+pBvQi7Ac2bnE/VD9vFGdfSu+DH90dywO6M1lgB9EiNg7U4
1gTrxQ59XllOq0pILccTHOlxzmBLkq8pNbpdYiN5iZq3/rBTgdyjbsytLSvIE+KW
dTHy2TlhGg+AqleZ2cCvWZrrhiJxf8X2f62Phu5ollotCCsasliE+PpctVvYapU6
ShA1FIBeahkfMwV5siMQyAzBWRS/li7KQiQExdOBPNzeNAidNCoz0B6kczOwqBtz
oAuw0DJS7Hb4UuhmiIeHryCxwuMWuWO+yVpRHdblKKucVKZrCR7y/TYxAz78zdx7
tyGenh728pm2I0DtNrwx+hr7kT3e7gearcOt8VyIttZIH2Kh54hkmwwY8/7TZKIc
JMssjsw2CpSyQgwfiY7POlMiUCyWSBzQES2B5Mgle4yiXtXH1GrVkEZnVZsN6KSw
yLdv3XwtmIlNG3jk3pj1BiNaw5xbdEBxdmZnJFbanO1POxX0jES4GRjx5ayM38k7
1O6ZPI7N4Dng4q3HNCqSnrgadUuXcYyEaeBKc2pn7gKnYi9MaKGphbr/uY3mnI8J
1OP7VAWmxlfe7uS/cVz0RRHXMIJI2y1gm6tBxgp4u5mWL74d3HGMxOvu6AdSSobt
sirASLt+WVYQHmxHKT8ICRntKSj0bTnHqitsjzWviwEzXlCJXTGC/wFDVimVYu20
NlwuXWnC3QGaRGE8CCg1aW4+JuPTaBP9SH+CKk27h9BsFuP4CRZ39yBdQB85s1Rf
NiOhcTdmihU1XXLbg0xu3LU8OmymOleiaws5QLXvtTDvqOCx8eL7VM0Cl7fq5bEL
O7j91wnyBV42sbV5t5QwwVbDv7R4u2dVHUhMC2MwkzVaW2V0ECYJQJizlGYN85gY
YnPYZ15c4Ctm7CI9IlS73kO36HohubMyUjD1neOTrNEFhKIsAkTYiOyiH9jsy9Dc
+VggdlJgEc00gqEPJYaS5v4jkWe6I9bhzqN1VG+zvSp7SGBcEsTvpLxWSdF6nXEv
Q35Bl3851va4h817ejGHuMIYtW8SOsrm/0/vI1ieV5UlMK8Sja4SY23sr8DqqBTg
G/+58leEK6lFMK8XVjdMahoy4tmRTPPy0cJmtKlEMOrCHt40zfTJTYvzVpNkFTp1
R9A6a4Ad4WaoRFwSAFhIw7T8Ch8qNGuOlReXwDX6F+UksgWNNAFpMN53ZTshzevz
r8BUFMEnzXAQblgSfs/sQpVuBNVhtY7u1Vh/hk14SpFlI/XJxWGdQpziWx1inSsL
kFYMwFQJfk1Jr387pyQt0mvfbq34eXeEkPvrGwwoTTRtERHm3RmMlBodod+bPoFk
AbRz4DUTLNGFqSstnP9ktq6Hf04Tz+3Oxxn3cpobQA/iXP8cQpRhKzo2feBs6pAq
oL9/D/V9i4QNG4XICevGaibD73dokKfRy2QAkO3JFN/ENqXvjzC572vpD6qR5St6
yGRgdDwYUHGKdc8R/b8H+jhQ5fS8HTLdLpdDiooPMJARQF0fopxw3HGfpTGXJwMb
Xh0NcbMA1MxzeDv3o0KEmhsuxzeXwlZnVw1j3cXklQTu7D9AbJmBO1T1DeNS3xqo
Hlp3J9Zq4M7+9Ic7hBf+NSt1TprAz7jw6PX2/ZB01ZQY8Y7PtlWHmQVeMwvR5mNF
EWGatVLemc7/7oGpiFEm5TZ39Jgb7TcN92Eprpd/7z2F4DK7pUNTUhzmXn/w213o
NPzQMHgv0Kil6+is5XXpR54CZRGD1TfFJhWJEL7UWqbH4ZBfVmYSr4zCtT9xZFul
bPOsfWH+VL8pceW247BMtHZPwUKV8MQEP1r9XnUQXN4rFnQHvwgnh6jpK70pV9kv
Q+K/KM1swBD49nMw9/nbecMS6np79FYj53albsPNclJqwB32VDh4zCzmrw/pt9Ez
KovL2fDRuV9+uVKRosTn61grOtUJycd0tkXqQ60Hje6tKgfDdivh0GrPWFiFyq+s
J/RsyVRRFukWOZoaJndZOfGC1Q+PcaeuTtCoflN0+IVV0BF0f8gxlA4qKl19FbRZ
7tWP6jLGJw1+HTBvbs3qGcSHIV/kRbGzY97IFLNVbp4MBMJtilDxrnObvDB2VeOv
WWUt0ZaWJQQnF/mIeTsOBV7oWb76mdDnVfhYFrLznxbBKiSncMS8/HPeas9Fdnvi
lkkDN2wKIb31HsgH2S3jgym58n3Tj//xc7JAlH2I6tli1WQtx9eCprYuW7Ot0Mum
O2oEcwN4CpkQjLjfyUGKUxVC93UPYgQu1uz0tQ4G0PfHVRdYVkKBeEAWpfjY3IC+
4AnpCRy3UeAZX5KPxk2uDSAhXH85nS09wObgVblxYO9gOtjN4AlTpW+geLJreKCF
gnSwcAaRbs28+iU8v88WxvXYobFwOLRyAiZrlVcv4DPzoszyUXPrQHD6kgKKNHNC
AF+Cds3TU3RIpsIn7QDlDv4NloRUN8Fbmpfg8tutuj0t9Z8CrJcqTt0upbislN75
3ikAz/1HTi8NOFqvkq5refhIhuOPNYX9ekUGH3SowzYIx9Y1dL0ihdar3A8ssXQm
MktG1BFRQhGuYNlTtVTWbUnt/4c+p9gdKoLskkiwLE+jmRckL0KyV0gfjEqKHXPV
yYkAFyi0/ctzwJULtCkx6OlSm2jFm8xjNSzvz8B6Q+6DvxOgl527uQ/bPMlky4u0
VxniN+lBL9NPFeJBu4TgKnqTNgeb7HCoP8BVixL6Vv/DFKX7hFL/zj/F8x2pbFPG
3CJtD1qJrj3k6b39H4lE7apGRygzExlo/RroZTNlzZ/bDJS2yTnhI9DEIgKagyI2
FNOdzRnWFynZN6olgfR3Ec/cOB1wALtU092ekTyl+SNaOduX/oPIUuK848tMiqe3
mIMZfQH1obRyQ1MDReowYJNskD+qvPWqHBt5JGBQzRzFjyaeIeyC4oawlzqhE0QB
pBuydVmmzLWPGMyNODmBjKDej6KA7fO4wozj7Zwawh0NyZCRIhs9icLO7zxWreKB
4gj282d3Q+g2Hkn7YG8eTOUDajb1XrorwWa/81AA9CPjGB11x6fahh/pWWzInIS5
DzFRh5uzCX1+8OMrvc95N+KY1l0L/bOGyRq417B2IAiRdbUCa8NY04GXxyLWGAWN
U2hVSJQwiexK3bUQkAuuoY74L8yGfKahjkNwUfJR/juRblMKMHSY987M3aJJraRo
VeT8i9hwxwpB3Oa78T41JjI89qBTM3bhNpoQjHLK3oTSPNoXyWyIi8ofZocp66If
8QD1xZkmRqpz2NtM3sUXwzafQbFo9r1MSEr4EZs1/5DvMuCPxfDbqulLAO+xEoAX
hBgaUaRUu8gY1fEPrD81mb2V3669nfPCMu6CHuatGZjGb7onEXE2nbTEK89lGxc6
NoFy0+9ky1EhqMjc6q7sIpcup6AGMKRhCJ6UHFcdjA0I9ETpQScOaVyFqQKFRBZH
c1TOmTiWZcXT0wEPF9e7p682A6LwALjhEmIuZmjon42Iro0igrEin78CZmjNPvvr
wNrQRjD5SwKP3fMzqqpdgMsklozZaf1iUStzBb4YBg7vy4pbTAZxMoXL2gewyRhn
3Zi9f3bPxXly7/I+EUCmAGg9OvhD29jIJh0LgoxzMkiWxW2VZM4qC253+DFWzx+l
5DSAmHRPktnua4nibFYiomO/DilXkHRUN7zroShaV2J4gYChJgg0FVyG4VuPlC4V
2Vpnjx1jSAoLyT6XmXMYiD5Ryc65frW9DL72oR3t3T9GDPaVgfULkXD2fD1T6+wi
uHowtm/lcnY9ObuBHj1NnczCNJirDZq2yWzPDzk1H3vLG3q0BrHQFIATSXq2dZVM
G0MBNR1BVdyci4grN5y47HcNwug0HFEMi/MhUP7U1heCJs9ZK4t7VbI2NYyv70MJ
Ok0NIQHyZJS38z/ikCNbJj5QNKTu+To+kY3/X8rR5yV+yD+0GSoNF2zNKgDbhr9r
lCmR+OR+qc8UoKHyyHXYGclFnijzSXF/ygMtQ0VyuCQnB61oOhlQzLZil9skECEn
vYMU8tCd4fCxXzL5SP6F5v0dJYEB2kJpZHfBnl/1Vwr2+tSrkOS9PjPJGecgCbc6
CUp9qALhSREQRXd0omxmxaEwo7O+fhZpY0Z8l4zx4fadIoflgPLCUmfYarcdT37A
ldtICpF4YnKu74m9cUfya+88ZEXQwwKgOOwr19sFYg5BJ703B9poFH+2ciFomRCd
UiJUiJfHtZ8tmYju6UalBNwCqvTWcUvc1h+VuvrAb29eYyi6Vtay/sIbu5iDZnoc
tulZPkjtGWFYPAieksTd7/uy3NEeWkftlK6CcXV/eg0QTs37CfmjfCObbRtqpMtx
Fbz5xDAaiNGFHbJ3qSfmjjTxXvzXBFnG/ATWpG6CCMZe2RtnfhJQaZLQd1DK0Tw5
hKgW7Eo3ag7kAVXYCKMGrR7h7+6Eixu1drezkioiHKWMKO4lUuBXLsFlqgXs8y94
McjPuNpVCcje1jMN4ODbpjQALamMXR65D6prenXFNx5LoSyt6VD7/POobo69vbui
5dWWNIZk+iHuThrFTokqS00s8LEz4a8rAeqN4gJzkfz73fYHMaWyn38DfGnosDUf
Yk0hZXgQDqfErZ47G0qh8wq6PeY18jts5bpJOtEssrYXK0i34a4dGpoV+2npQlLp
rX71zQKMILbJYBleOgfwjWQ3mhgdLJiaRSd0IPPZCo0WVvVNaCa7D0k2/USox2td
fCoiFBbpEpTf31TkiWOMaFy7WYIdzc22QlY7Fsn5HTngmE8kqf0niX8pX7k8d+MH
6SzRHcv7jR12YrxawgIOJItQeSGStLaOQM6GMOIxMZvJszs8IiY9mmVdgNs9eh+D
dsSO9K4uBfAmMBuQ/L8g2ZMXQUzsHOs7wRQ2VyyOwBIEaG3SyDfja5FzKin+Ud6a
akqz8zCsS/YNu9nCU9kYjsg83InMyyh02F6d9j3LoRA5mK+UiEdJu36WivPG3Lnf
a5kLbCpIAypP6fkiQ0I88puGeTs7GaBIMH9HinyJiOPhfk5oda47Vs9PE57zbWLQ
D+f92ZPU09YnQ2MQ+91TjTA/0ijdQJhQKSujmaylGUt7ts2/wmw71PBRCtxbPZlv
RXytj2zH2e+nR64fJ9uKNuw0RJuxe9C9jdWpdUog7EN466277O0xZZZRqxW58Fjq
PlYHQwWlvdnL0vWqfeo9Eh+bUXLxpmQbyRObOmJJVw0kKL2BJ3tQqijJhWeE3wju
XnVFtnPfEU9/7+NZbsjUkHcrHVZCoZNApUqIy6VfiSs4Bj5GJOIHClHBT/rDTveb
fhAzvlmsol4aDXZs0WxRnyRUhr+6CDVGJA4IsHndzokCIau5lW0hI5YaOTG2sRiZ
xMYvztArVDzwJ1dfieA/OXuTXJVezylgT6ikaoYMjzZyPQC4JeqXyNlcBvrp0XWg
5cMDMSFBJzJ1aft1Tbeykmu9hz/IkL74mb+r/aMIQAH69ExYp1Bffz/UXYQNO46Y
CYXXnXzPphGyP1w2ytlNEwoTby8QBWLVTxcXFAwKCZWFD/VckD4E00/MGg7svefc
rEF76bvKiNliw00l0osF72kcunMBs6T1gpHqwLQmxmo+RtdLmq8Y3Ni8AMYCKbs/
pKvU+6gAy4+Ho/T43roo36hq2ivM3OS09o/G9YWY5M4BHqb3hZ4ZRnLrTcpry93V
OR50ME3dppL6Oct9BIBP1JQeMNshto3hrVmpE5vc8KNnv99jelxx+lFtWLyLwRCf
dc7RFTEyx0L4equkIBWQ3d6ZfEfeRJ3FkrbDPV+jJTVKxaaZ3ld+iaMFz3y3WMrq
Ra79e+ff4i7+KRSr4LKsUAChcfoZApws5YERZnulObdEi7DUkIl+WhJQ7+5mn0BE
1e+gUSFkMNg2v+djeihd6CuI3UEWRdp8YAXXroMVTYlnpkfuH2OQCu30wxv985kZ
iXDDn+q7unkC77/3wfjPfmV8MVhZTRCNZomV/D6uonJzaLmMwdIzZqQuHHyFxApQ
82DeIRkKnKxL8wq3r9KcNw4T0mPx6LAkukIynFwe+RyINoYPr7HQfi7zAz0f/t2a
6cXWO71dbIKSCN2N5yCS8XzWXNs7m7hRhHXj58whStv/Xeap8ymfN1mGx8kKPTWb
FukYROGfiyASVPtd6g3oxbTAlXPyl6D05uP1UN89cL8AYOefGaNsFQDEtZGAANVQ
A6VkJ0k3XwD69XTUVlLDKJIa7g+aGqev6F7k2s9lk/8HY2UIgT9/QF9Fd5BvTuuf
75Nmfcx1deFkjAHRqhmYKnPOfxDGvw5WkHoq/+VmgnEUpOw6FlTBDmU4adxsM3Hx
EvSNBzXz1uF5neKHcYmv6loqBB9wjW8AnB9DXy00MD4Dg8qPfGKsc0bhpwV+FlNk
zQDrxr22q5G9INKDWY5Zb5CiYKVUYe1LzP0W/8BlMjnoa67CrdI6vdFw/XNlUN+Z
ipi8IqIBNG/oDNwQxWYzuCYVi6CGr5f4TEfs0KyTbNcGrC1ArF50cPKkDmQiD/8U
cizku6meMngD3Pg/jhb4l51Shk3M6lcbyzoAYbOTNYdbh9PAz3tEuPaVEv2C7sG6
YYQxMOlHGGCdG1xIcMAhJunwuDGi0GV6CSawnX2MZTe6SbxAiNDYIQ3RDAYxJI8K
M7dMPuHP9U+1TJwj3ICrExVEGZAbSwqBbjlpXGn6PPtk0U1Os14sfXBZGGoouBrM
ZPwdg2nJBsDhh707O3PQf9Lv2Tp1rGr36V9BxFJ5qrCaxkEO0gGPf21Q6+mcpQuO
lB/d0yes7WN1HaMxXaiJsCXcnbh/a4u0W+pJBmN2gpCMim8hhb8xcuN5eFmtjHt6
RmF8ldO3rJjohhjtywNETSvNIa57JUNrP9SqA+4Mk23uIwMmpc363WZZpAj5gq2j
BJrUYHov+/2IT1KbsgpBB3yZ1DYZvAu1+Wcko5lEGtXu7AnoJHL0om1xwhjRONlA
yp7T1bv6kFglwEmDxxtxQnTvDug+GhpPUqs0unr/Ilc21h70d0NZPxgSWY/oseD/
RvsBbsQ5b/HDYgNiZA5UZ+CXsvoSEA6Las/BSt9V0hK+Z89U6hBwo2x9B8ae9Hlu
Yes7sjxOAKJBzF6ABZi32Dd/wlH36ljjw3PcbOiUE9Qoh6KwXCNUhNwW3HxitxE6
/XTdDRxhTC2qvtc4yPOgCmHyq2UTe9nplymXxcH3shV6gBAdxXuKgrnm1LjdNEKE
zUs1zTPOsV1+tcC4jQgay+hADni3Jh/QzFKNt+kOvFv2u8pFYnxWWHcEfCyoAY9p
pMbEp94Bp1ucwN8deDjVWro35TqlJHK3ObyiizUx8iP6PJsMY7QTHV8/tc0V/uCj
T3zFk4n408zWOTQdIj7k/ZtxZQ7ZFzrFrr/5URJvvT+oYIP6FBCNSSOF6YyMdAcU
3K3F3MBs/mopKLbshqWGFAUHzSrzNMObe70vub/MzxrD+HtfAwceLdT5oXLt4FE7
gysOv8fpZkgUyEhFe7SkoQxe1PAADFuYXJfOWlhpSrhnCqSE2CL58rX1w/mv/BWE
tGmNA2E2kZGpO/QGEwZYiYW00Dk/OyBcFAJzJNEDYhZvzrKg+dPGzSKy6v8N0+/v
JwUPOLh2/TI15o1e4yOL7jTx6rwkbwzPNjY2f0TLJTV0/ZB2HxQYht3b6Yjoek+S
AsrE5n5AWxBeyn8BOdHKmyzaD6kWGyGVnXHUNSWW716wvK+X4oagm4MOCty/Othr
fLVrjWTscMqijw74sEWw36pUGfNwjcauN2bTGT8qSXHEQ4v7tVgYMvErj/3aD9jY
IKuKmqOwYd6YZWYX3PKz45bQw93J9lPn5EW96lwAngN1Il0KGy/RK3BTtYujARS/
FqAVV/OMOTsLYAHFudpbEzq/TCA1pMgHmNhjwhEFlEj/pHSG8NRn+Z3fbUazX8Nk
IJTrX2jUjZt+83e+ACaib0SBi49AE4VkhK5xUViH9SRZww+MXlwU2iYtjqRxurRV
0ArMg0wOzakUspb0zE0gdaVMddtGnbX2a//aOwys70H1LfcpWAgdBXfUGx5yrFnJ
Sd88IAsabqJCeRrGQJoNQOmurzQT1d5xkoIFzsfHuCuhIk7DjfYOStq/MGAq75Ga
zpuSTR+G7RtYR06LYS92zWwhYo0WMmrTWuoWVKWNn/a8Q3EuWaUW4zB/rUB9F7GB
/h+00QZTCJxyOiykB45FbWU5vlOpTt/a7HTLMNMrQAlYeu0W74KVlz67ip+zdCnc
cGCZxsnt8VCoRW+hGBALfApzoclngBH1NoozgeowRwa+1I912cZ1VAciP/+8ZcwZ
Ov/y2oxIbCwQZWIOwDlWAzKB1A6hfQejPG5z0yH0+iYFGS5TeB9LkfFNu5+RKIcL
0y3tvNpyjtuoLUU9V7muau2ZpgpySq9jSPgKB9tMH+XcJ+MVjSzmEoMgVykwwByu
dX9a9fhrLfRq37cSS81aEDclmQbOTk3zB02NPIFRncF00yueF3qec5+lCMim9VsR
YK2fygpZuPEDOJH19hu5ujwk5s63uy7JhXYRH8QVTkkn4FI05iPW/q5VVr9aPuu9
HdDs2ycGQfw7U0fH/sNZaXXhi/j4aL9POD6/07Z9Qd8eK9oseNCM+DrMitYwshcK
ix0XKBIps1xOrJPSY1yjcCv/R6hM8P2rnHCCov86kfFprY3x4/yspr4GyF7XlTpE
MlAehU1Bf4T1X1i65gAC0o+BgUz/AEvI5BNuvHlR50Zk3SfYZRhIGqyV1HRKjMPk
ewmxKGC7FxGMZSoCaj4bwlpSbu6RvOgsNCHD5NEzOkLKXSjZXPT+usXjweyPDeqy
UHkmH12CWKabB/9zQhB4kNgCEH9/3NhLobdBx2TAdYMnZqnlOKT/ZINYA6X+RYVw
Y4+Uwck6NLYcotpwUr3TR2czO+LjQsjOwbCwG1rPsco+xf8XqQNX7QSiaMOmtCic
yJCMSQ7Wgs/EbUH0uaSB0Pvaq8cVolYpL6EzrDQM/+BnsNS98phji8ak0nKzRL5R
OzFusTHU+f1N47O87GAV0OhXwtj51702w6y8fzA9P/vNBIJTGnpTnwBHeF4uRLOs
GwBlQLfT0qJwdpHFOJnJ22eEnSVYKx7Tan9V3pZH+8tEtK2GCYVb/IACQJ4ctXE5
b2kYb+Jg49v60CDvWOVNJobIOeabRdasbq2ZUdQPHX8Bd+CdWRzNX9zQeTlU4OZa
o9ea72eQtkuga5F7QdfWykUcr7fhBJvBJS6t5lD5hB0nvd4gwV9Sip+Mq92eUhnU
6qsoaON78EC/H4RWvmSoEi/S+47u5zupngtqO3QM+WGnZBNw/Yl0mcvWDgeuYhEv
Z3E6Pjx1eBLsXFAbyAV1gNGQdSo+5oTrWa4bw4eTMF+8/SSwfhhu5F2W9sGB4kG0
CyRnLzj/2q4cTEPRAhRjcKvMJgeiXmBYHT+9PY2p1QifYlzVbdG1WcVCfjjIIbEg
o5dmoYOxeNvBwzjTjsAK4MWYH7I+zVWPTFItOVkl0yZASzVnKuFZl6zVfaz1YE0c
ACHJszzOvPBuYugRayRXtSbuZIYSV4Lbsl/ivv7rm0P4VUGyLHQfJmTrCjAG9eVF
XPpASrINpSPYfzvXfmGMTR7LcLjGC1fX81LNiHhxYvdw+d2VzKb1fbB7/Jdw2qtf
iMTbyqWTwT3yzJRyBTSyWhGBlsCpU6Z8wXP4L6aJ09K81YIA0B0fxYU8OO11MnLl
SqR8S9uGR83ouPR44bnk/bmqPcdO7gNc9m12KV3G4Y53Xpl2ZW5pK+r0EKqZIpwa
pzt+x8dkAiG60zgYnuaSPKjH2LByxPDJ2wofCjXqCEaThf3pI5c++TlZc/jhqP2k
rOrGbyBpRRGsOJF/jbd82T8byeoSC3/tau+wKjF2rWp1UtVrag3l1P+c7gBDWLJo
jvojwvXb7XtcFxvUgsornTzGpz6LD6Kpsl8V81GxGpuEzesZlIN3UEw66zxsnHFl
OYIGyf/k/r/HfgECRsvcjnqdxk81Sgjqcux2koHq3jTCsXnq6k08AioB5aRPByMT
nHfjJPgQ6ARz5Ni2Gegs+VPlp8ih+aviYLOxn7+a62YQCg8bc47aSORtotM5sQD2
ApQJy2ouuFvX9OPFi8SJrAh7V1D8ncXnBD1JFkRIv3kwmVMj6gs2ImrSuzRuGPeM
S3qIkYAGmNi3PfP5tfuTYXUgLjNFCMs53/UcZYUKdSTPKfHx2KcUiSzGI5a1rVkt
KZ9jxOjBpwCKoq6Cmpkl5xqmyYFjzJDe23MdvFAXYy3hLOizNl1AQQx8YpaN1UQI
BNS8sw7nQDs+yuchzCGcI2xFzVhT+0peez8DA+G1cMGgEqagmr6mTvtLH7sL1x53
5cnzN4YbvlNgBAgIFrxzUkCGbIrQ/muDYdJE8Z8TFrUikY1jaHVw0tZTEiFmv3Xk
U17LBAMjdkxvRwXUyMChkqyJiKy0KwNx97izh2sk5TsUUkjaWz38molOWwlus5gZ
pLixLGSJVzopRTxDeQ+9wua30P2nMWk0FoPAIN8rcg3s/SAIGzu/uP5gm2MNOoss
y4M+ryHMn5zFyNODLfi2CZrWhhJc73vYyQ+uHST/5LyCXY0y2tjazKxsQ1dKntAD
WD3jU54+Dy3GsNxIOmgXqwvPl/RGMTuC0CppEDhAJhq9g26KrbpynuUdhNcXsUIr
ridq0O0B7b8YUk9mthrvWKsPlL6Ia1h5J+Uz9Y5TKTnGw/uVtx0NApfOuw9qkWEE
WcmlI8JuAJ66brHO0uIipNNMw3MJom9TAHOm0EPiSyW7qAkalwroeEtFPTTE8CYB
NlYuIGe+4we975SEix5lSAEDynWVlYTLeZ2aAs2cGtTJAihnvrlh6gEQMBcusVWK
chkCNenxYO0EqU+052GS6J9GrcM79wnUqnpp0raZ9qT7keGfzCtsUNQcwYjK12R+
VrJpetB8RfZ95BVTOydy2khvpx/ljWuKnrgJeSQqlAIxuUVlLeD/jQCJk2B9HC3w
oKFlbLjaRstIpZKsDrJ0vDb+FQuVGXTm/X5Fu41HTxi3noGhL30xShkLfJsW2DpQ
rpg4vv22zSiwhyaNF26wmQ58RQ/XR9xzcEEBaKvoZFmbGt43YHoJgiyMM7pIRxjb
v61SAjfNBzpOgaO9n1wgEFLEhv137nyT/Ic5Xdjb7g+d9c5INiqN0iaq1Qvvfyfi
I4CoAveDvNTMR/eo+yvRQXazFIsaRLbq9eShEt35cd4AtnhHnXQ0Q5JpVLiprjdz
u/RKAg2O2oX5CUZy5zbeF13hU2lIKWxgQ74lYfKp4hq2C0ceGnhJYu4rU3jqs+LJ
qDZnCH55YqVtNlL2XRjNNfo22rZPPA5hnth1xS6YPt3DX95fcx+chzNUcWdKyB3/
UjzY2iyviSTqA0es6dqI2tgowXUs7EkcSGLxZNtnFKz2RMYZyiNTnIaCL1FifRo7
oSHjk5gfyXEraFTPl2bpYdw5d35UWW8v/H9GAo6AASOjTXWShBoPvAhA2NfKnpxA
/g2HT0KA7rhxqU/dB2mx7tPhUG/cxa+62BK2ZbVxdY6sHhI4sW9+qJYFAbEBx3HY
1/rzf6X8gmZcXo1abww+BUwx7mYP/NXmAZFZ0fiC2KLsKu13nuMUEQQyc0vAWOGM
QaYXDzBnNwCl2KyWmB7vgAEf2lfH7GtrzMiN0YE+mjIhe9D2wPKGd3PZ8rPPLMGe
nl71eB9q5yypeOYy8DgMGzzje0GUbPtTpkJMixExwYOYmZl3bHJTRe6n/J3bf2Ns
YCM8yrlIEK4abXgBOsrEA6Bh2Zey1zmpUpFc1n9IZuIIUJ8wHta2n5OThlfNMCU+
gg3MfryzQKhQcev1VmDXrScWl8DshVn9yah9YMN4tMl7pT0haVAD973NjSOnH2OU
5evbQrS/cjPTw6fpvLWa8WTdYEonOUNiSN24olhPEuAiqH7m9y3u62JYKQdXzZE1
UsChPi80KjQXVV1vux9z5kBOXFCh3mcotdNgSVbASFI5ASCjdhNUTVIl71TvSieE
FDH5BUo8Fv0RitsLHfsGT4rXLiOgVjxPLhcFSQjTcoU8KfRGI7EFp64zMi7lrF4s
Ndg1afiDBDOdqN7wV6T1Uo2ZMF45h3Dz5dRA9QsTxlyAk9YESzKTIuoLcDnZW1o0
ebJPumP4yEp+P7y1IWPjFmNETIiwwTxMXuon3rhSQtnuiksa7MNWO23YY4bW1XVU
aIZ09a3onBUnfG/SN+J1w+kUsVpgGKnOCExWSd+2Pb60Xr38NHhxoxyO6NDcE3Lb
OT6jBl9OLwLfHK4hvB715a2hF2De3rAbdT+GYleMb8AZcSTBFreHyB4bIV8IjLGv
hAE/iYpfW2nmuJS7iAbgtAmIMkSucFmo+XeiWZWjiqHndXysb0MALCLM/mqxUfe4
rNrMGBCwIDocfVZHPfzt5ZOQ4qnif7TbFFLF7ALcRIJWnNOqnffjSaAgTOjUQmxi
kMNTBzqfHEf8134Asq2ikdozk8cXPc3805zVKqH7ZKdoAJscW9fh7lABgCmTyOrT
PuxrZg0iAKfWqvkz15iSKAs7mCX4ri8q5rXL4yjNavIHuoQb/Js9CMJvf0uTylU2
XJ/q9q4FltDjz9o5J6IKsrlc79ALNEXD68aNSufcfQx7El7x5qK9FrtXjne/KAbT
9+CbFSDAwvvm2DztQNtFJoCtQP4NVAmVIrVHuT5yTF9mQHgx4IkK5kzp04A87gfk
WcaqbaVNgGs4KwVU+ONef2leTb4dKBComwbRGn78p2gdLVjk9sj+mNAwsCvMSHVK
Hy6DnhE0top6W5jH5hddvBXXDrH/XSo3q9cRqbUkfql0YDBIqalMBRZkoJrUKAy1
v7JoNnAECVtVOmsUMbtvPu6ANVKapG2g+UhhPo37gTn1LA+0C2SLqp5gmbm/qgij
Deb77yIii0tmqoJG0GbKl8TK+RHZk7/qAo/SK1IaJhZqnY9yzhwqe4u/wfu2mYVI
zGnhbfvwVbkzMxyN41egAz5hnjcc+ZI6C+oZII1CrAP/GlmIFQposWAfeKrD3hkK
li/8O/mOa26m01ucp6kh/rrMTcry0RENe6dxfi1UNDdPIOyfoKgHApv6EYJ6rA6K
JslwsDevIw9eIragWXDpFGzJsUUe3lxy8z+PEWwNwtPlUSYv/5kgfYRH8cJi1QLB
+qj5tOmu6agv43yDpkkmB1kj6a2KSC8dvK+xjwCDtjstm+sj3qa1EBGK62j+elo9
U80cOdS6HN7+ydRJkiU7AJiAcaGI+wT4cagbqq6yptHpxlzX9RdnfTW+/iwjiF+h
SakWMz0GHcnyYEuVIZeyYat/aMdvZ2Z1n1om3XN+0cRTIq82GJ9G10oR0iXuM6/d
ysV/9AdB+goMo1x+XsFWhrWOD8WebRnVmlmdPC0teuVv2iuvhOjL3g8aKQD+vK07
4oCGtgHmeW/XZ0mvcZ8HpPcHqEYYVlAhgJpeajdylqb+2iobrBfw52CEnZfPOPX+
gKF/RV+30YY0/Z5ky715hi+DXeYTnFELEKjspx9xSwxgGoRAqtB9ZOpEnM8V9RlI
Qyga4+SkS9q2458DBYhOfJTESm1eACjAt5vAszT1E0NY6nsYsiffThGExkdSffBA
5/gMSR6PsTEcR1W9u6XD2Vfv6fwDTG1pNttTYZbzUFCgCGLhuocAOELQK6AIloNS
Y275ssXGsr+rpOsSlG5KH7i5CnNBb9hORXAxRLPAz3m9/SaEWZRmm7N4f94UQSyh
4q2xpJ0fsXYx2AxyCLKnZZQQq6escueEnc9mTIzLYWktTbpGyeRZMUBAWB+4yPr/
0KmhsJshUgm3kE0ByDExg5okPUqMaVeXDXEt1/kSIm+JjqJlv2xvWRrhuIqTtgW9
2UydaN6yN3IptdFk3lGQetJjIZYlYDqoJppFrRgV3AQcKFN0SfXWPWgM9DqMilMs
kNns3RG1eqwlCM0eZeJHJg043dLttt5pF4/HBlX3QNPqL2YPf36vXsuaTnRjAH99
xLwF4B51a4mXve1WFp8NiNQKR2D5lHKxymi5TlDnQU66Fnyo0BW9DMwbs7HArRiT
R9Bs5DK3ec3WD/lqZr6lTL8l7yUhR+eFAJx7Czhhem9mf/cLjb/XLS9Tdgxzaigh
lSwyJW01BihPgD+tcoIuNcJwAZBGNtV1uDA4WuaDBSAXZTcEdY/H5ppwkYkLIM0T
y6x4gxVtIDKV+XS4W959/qFxUWQmgE2nZGyfN2tguhr4PmKI/ce2nwyLA8MIB19J
DYDwl/DQa0MP6WRBhqsQL0+MmgelLxeziulU40+PSMPMW/cQO6P++60G0OxFy/eY
y9rHdvVJXNT8DKC17lVyXDGy+drKW92W2eBH/+q3ktWAqqIR6s1XSjgyeKBudqOc
OhI+d1vnuC/HX1pzGM4sc2V6aonFAucundlM8Qe2FqazbB6dmMccI4al1jeSRZQN
FQx5Lk0JX1cxBR7fE2YCJi96t4PzfpVuTem8NOYMzKiyqxwt1JBY6nAXesqqAYZf
`protect end_protected