`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5744 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
HdytKcppDjja7VfYQkCqvMvJ5jXBK1LIZSzF/XV7iJfqthyWPddsaZgtKGRU/PqB
L0FHhhdoaWCJu2DUtljIKbMe807/9EPSL7v8NrN+y+OGGqp7wotrhVrucIyaAxC8
fuUluqL0Zxt2ZLdI290rjTtZIQbMZmZPk2U/IR6nHGQGJ01g5Wg3TQwGSXVYCcGG
yQI1lDarp7Xu4hnitt65okQbzJ+8a+SiEr+wzpg8vJXWiz7j+sZYkWBqhXP6wFOE
nRLXitChc9XhWyZcAcQzxQpirAZZNIGDNyd8e8JqudnOvzA5dd0npL1955md3MD7
asPDVhJiID98++RiSeXLM/2nbr+cHYxtAQfvICuMuydAOHWcHsyplSVMSrl5drow
ozuG+eEeXJ3yunqtK9slmzbd3j7M06Md/c4O0no6feEUmm/oCTxeW4liCj3Ec+1t
Wm4tmkEL2oJIQzOVvv52c7H7KgQ08FkYzBL/idAjw+KVAnKK7B3u1CAmhR30jRnB
YgIK8kL3snyLqT9WAvmHg3u5mMl5qli8x7ovpGoWBs6wM7vaLtKbAPeX0UQ/Zl6W
3B/dLo64rNdvo9UddVdGaLJm+4qYg6KTS7XBcxCSpfXieKpLO8L2ZrbXM42FA7Qq
lcfwKdOSZxVP2cKwk3U4LP948lfMpsOmKPpa0knMd2azJmeX2Q6GW2Mw01EXKzqr
7+tdjeCC0LdFMJdKmVrP1lLYiH6Z9RrxMXGnA+X8h+dXgdGps+D5Tz9hvT6YB0CM
5Ae0PqIEwntlJtLwBKPSTeoHfMXXgq85w6XdxiQQ4GcFoTjgAzPRcOfUlTVKlbtz
94M+GyCohooQeYm9m6KOSgYmMObI1dN9c1K0QjfQOrXMk9IcQxCd5JNf5JDMY2mw
a/cjDDayTo2vnnaQyTZqiH+ljntJjliQelm/0AVvU9neV/zao4ADNnlsIRD/NnE0
Sq7Vkpt1/K/ddPRSpOYwmfvf7PXiMEOhfSUDlYJ9OTqKHFwc1dAXCSb5e3e7NM1Y
oOWMvySzW57vu1RJfVjjHhvYUQTbu9U9/0b7NRI6CSSBCMPXcaXRItVjN8wg3wX9
/3Gaz3NwG1WuGVg2nPm0olo4MUIOwpq2FPJU+YSVAUYzJdmoDCTjiUIqr1R+HROw
dwwlY2XSIEG7dV2FHvCYcvKLFEuaJV9EZo7qIEK3vpQdprkN4ZRxsmMDuWLG9Hik
PLkWxsNS6bl2UAujTLERTusl1OFIP6vgSXKNhSdct6GXJGoZZ8m6LGsKzaAcz5K5
upYUeY4OH2QFgNHKeeSVL4IQmZLajTvWuWt+Erb8KnAMFcrdPQXN9v8OieFpmPru
X17uw1a/OaWiX5QoMgsNRrYs6aPIy19g1Y3/qM9D88izRL5yUMTGtNbyEFBBVgQ9
cJHpdcorGvh+KnnMhfjlcfFC2cC3BKaf698uwexiSaB0eFzSMH0mTPFe8zARWFQM
uHX1LfpHZFf+tIB9+KDzc4ijVGaEqi0MLhNcHfCryDHHJMzZV0eVIYvBqJ5/KFx6
gxB4PRbAk6UQHVXIjkkezpODOlIYFhoWD2eKQzp0orFGAQRRRr7ukGflWnq8iTqC
yixKKwHirrtlGYWry9oVXoJ0v0w2yc35t7D/joQhXgQwOpgbRU9FaA/n1pf3VgQp
T2jHGtpfvxGcoL1uxfhsTI7+czvfz0twQwz7GxWRHl92I786ycp0WD+fDq0fUiui
YwlZqsAEPU5/ltBT01QjSpalwaFF3Nb6R0QL+zIOroryNwcoIYXJQvYaoZsVlrUk
jEq5Ks3GhNLYVsA73AAJljhOHduKElSqsXoNO3XF5rzj8wOOyD7gyLkcPGKVXMqq
DXFl37troM22GmkyFitSy/+hKVrK7Q8v6zpA9FWiizlW2ElYlV1eP1Y6YHvRrV+p
uKwMGIb5zrWszSoGWzh69rAbX4UArtmU3OEF5Nl9uBJNDDj7/pOzA6Nbh6a/cLd7
/CWrojEJfSu+gwU9aDKcLRjjE+E4Tqd2iZP8kQ4d2JnG+lhtSCpJUPgpuoUEToVS
LCwkrMSyCNShEoAM7TziYDeeQSxYmPrVz/7r+CXvA58P4EVCk+uVBRQ1D9v2/2LX
DBexD0OQHSpqkkQuFqGdMaQMuvj6OUFmhEcVOfH0q1qdPYgZh7H7vWU5Ku8XZSsp
gRV3/O8GBX0VoRTYEEBRTj/t0IEglfCPSqQwLk2JfaTZgEzyj5XQpov8wKVMUzNs
dmeF7XxSGBFcFQLnKPkfFjSx1+oDnXHilJjdsax89wAplnHDGRcv9eIY6pA8lJiS
dfngZ+KsFiMFPyctiyFvz9/HJAHcoZZFSUfe6ly1/YwteBBu9LoFkT1t/O13MENH
CUMuyI9LcBiRKTw3oKdCdSuwtRO1XuE0zLmeE7m3R/VIfmL2NZQ6fTbDE++erx7S
aC6ybi1Ex2qp+p1LeCO6pVoOyBNNrcoiahesZNeBoIktb40iWAWRhQGHdOAfmxdT
XV52iF1eXJhSvKX+WB4Ux8OqktfkCRepsr70dzKG2onJkTQRhiM0k2tKVViZKGsS
NbiQLNRVb/P8F9P8lR1vmla5+ct892+XdN1vPNz7rZ/nmSgiAfmgbSTxdsD4eOog
pE44a3yUpHbN+CAVKKCZ/3u2FsgxauR+McxOTaPb9RrbyqU9QfaJwiZD0Dpm6ora
K9k6phxlWRSFQB4eLudeoRBAr6SESqBa0CY+uqsEIVTY4RgwctB9NZ1cJ1bxP4eI
8UL3TWCf3BSZWV9pWfDIZyWS3PtL4sjOVnbnIEftSpHYDGwCB28anyPfILqHvj+4
8NO7AcbGYRTb+TOu5pFlKhGBQdjpu8tKOLbapCeMkqszdn6e35drpqWv37QOzvqw
c18zgK/Q4emxQJZAyAT7v3zTLQzjXgfPiBnwDqHXbZKI4U596UEM28iw0nOZMDnC
Z1bf6nlv+KTQ3yEqMvLfTefHSbWRWvgsqObmeg1AC7oWLDCiP9E6YCF3aEvAjmTV
trLWrwAEotzAfoUXDj1+yGqWxkPmvuSgAzyqqHhh2UqwIytLzVF8WCfPcGSc5l0g
6nVqRPsrTPBrnDOENaTmJAc9hyhgifW61DrUbGCZVhLZSsVe16cvujUWjM0h2NNT
arjvTM0Kdr8dOUHZxq4PCx4bOhlSxeYK6paQqUS71mdgRH0icxSUdm41jOdGTSMZ
xEwKXDJgZujfoEahCnkraMEDTTYq77bSE+WXM4lG/Bqx8trkCk3QHJavfnWIVL6E
1cF+xk2U5I3LamnVyolNWBf1xYOHILycsAYLtkdVOZ1UKnB5sxShl/6JOUzowT1l
csxwEbJJW3NoM09e1jzAOcspK/NAYILBEznivfpAW84M/bGN+kByWHJSCt2RNEvK
bVA0wvg3latzGd6UOPlWBrue2JTFBGFU4VwPUm0ua6OxqnOHSr8A2+IIOFLed3pX
eMo2N0FIlCv0A4h1eIVmbRvlOnjurDt/P8Fp5hA8NW0vs43Yp90hOl6m2SVVg90z
GrBf0xDLS91AQsXewSSSUJgblhcV8Bztk5PgrgTxPdCrtTSYHJMDXBbDx3ai4xBj
4UWyPfDLg5m98I6UzBtkpUr3WkPC25B8uCQj4uoGFcpvQwTOu7lX538iBSOM6zGX
tjERuAwiwc9c3opLqZVjn/YZaZEo5QRB5uHNkacKHTYvA2XbNFCHx/hx5UMYci5y
WazQWFJy5VbC5KHnUyxHNbukPrXNSrwjDZSMtiIGGg8LZ7vkGvwPX698KREZv2Dv
mr5hfqWl9b9VELvmhtBiaelL2QagDIJoMB1cZUeFmb5hL6iKH0mXsMmol3vdg2W2
kJH3OlZ0TezoNdLhdlaKvIUPow6Ho5fYwBr8og5hfZ5D0cXVMKvXy1cLAB58wXTH
XtVihjijQVtet3IczhRjWr7kzgz9KaaeRMHrM1dvXGHW/MXF8VnuJMc556/EaBk+
xjcDnl0yY5SOC7GJwZ76GamnS0FXhBMgDiPrLuKSKmpADbThxRLi0nrPsU7Mh+fY
i4T27BkS+RUPDzXkQk9iuAx9C5c9YfThJe9Vc9O3voSL+YTS5DlXtdP7vto7Rz2q
WjI/NkEOZTEJ2VXPLe7EW7ppXnT1RdY3W010SddjsXsF1kjXbYIUfd0H0FgV8o2E
FbMssQHlFXb0BEHVWAIM8FvsYQrXZ8J8tpr1K7Ba0P0v2xnNvLbRYppWKeTNx4xC
i9d6utknvqm2+wRhomalDc5XoQz03jrTd5aAPBGhPG1xMgYr3rzm7s3Fy0lnpUFJ
dkzLgUcFyyS3AmK9OCEdnEelfRgFIOnZJn9x8qbhcqcvBUsm6poCL+qE0Xn/bmPU
s9FuPkNQCMt4KnwMpQjJweR0wDfxLDc4tXp3l9d8BmC3FU/8WenpJAs+TBDydwls
0lipnUZ3y7sxKe7bdRqP9WJaZDEvSFv54PLeLz06SfbK4b46DXyZU1kgSPoLLX6O
0hKtxahZVQG/lzAm/AsVWVF9FZSPAPkluqCRJNt6hW2MzAi6Sd4abp8NsEk56Zfp
5vrBOqz2VY9hI1JBpKMceleVhO/5OnSJritYVGxFRPzPkLXWjFLDBZpo3uVe8Prw
x5F2RrCNjaub/eZzJ902WrzGwtrVwY4xUXhatrj1AGX8X5Ow55Mpt9guPgHraI7i
CdJM9o+G2noC4iegjiJKczarxT0K4zzb+DBcmToUxIBtqkBNsv2L3yjU6uRA3G5N
po4WbM1qiic8Whx95zfRFcp3XLscV0IqE7DFtCYr2VK4E0coixkxnQ/jDQhLC0vw
v89YReQufO38iaAhI8d1a2mtoDDe5nnV95PRuqkDlNHDx+lqua5+716yvfCmM65o
hx39JyXYQke28WdJYREKawEH21CmU/vVWmWUCahrOE9iCCSTgggsvRiImFqK0/6U
dGafL3QJzeMtMYWeKO0U7Lz48lo8wO+XB7h7HbMn7OijCryDg5WJH7auT8BhPWKa
2on7+yN/6oJ+cQ33FUTYvBlieCW6vxZKlvxJIrfDkcZvZlhCT+oio0BVqm3x5OcY
UQaKOYFp6K0iTs0CjjqbHIYsqpo8C+erb34BiSd18O2D5AFH84QtpZputuQCiXKR
w4gsfJnq/HRUjx7mnXfRNkUzeDAgqEA8+4P1a3qNitVC9WEtSYipOu6TeKZv3VXe
lsWqn+hdDxvfWPsdI0pl/4AlNh4eKoQovlF2W9cPeF+Fm0ML9fad4cFK7CwF/VPL
FuaCWRboY7M5rpDKG8EMCvYZv19t19HJjgLyCyPgHL5JySNnkcPxMnPjn7TSgc1Z
uWvPPAYjp3yepjfs97a5LcWAUDktQZLaLKDYWSrmW7aHQ4F8k83Qgg3W7WMfWE54
+XrUviuksFY2CEWk8sdf7eUiaut49Kz59QHHnnaRpUP3KsnF5QE+xr8GqzInnKWj
VkAqtQDINnoCtu3tbemiJAQFgpwKrMWWBP6HEjc8AWIDCVZmi89yCEVJda6xQG4S
DNl4zDjVK1B4kzjZVYnEzpuFCihdOwpHTMV1wfuVNA1qi/s8VK84n6zySAgsDkU/
tWDkVnpdNAT+5hsHdO+loVsJRKxUOy49TFi/ketvhfJy32bKapF+HKN6jzO6Altq
mJ8xpjYjusSsqdqbodovqTR1zWVh195vibKRW6jBGUKlcOGq8yydq2gFqftVS/eq
VAcIKvFW9jkGqeH6U0PaQ/tR3dd26p8PQkJUxMsbiEFZmBtvm+fD5ByjSCY8g1j5
2Eyxh+nf8m+fyauWu71TmCuX7QmsMxoSyjL1VyIR1RnMGs3nup6A/cwhEaEsc7Cv
T19SSMjR20A62oYEP/9zkMYyX1pVqjexjYQvYQXziwezSy1pVVhLnQ9tm48JmxXB
uaeBmrvdGRqvLm4RpQ6wB9BWEtFB2YdDsv9TZoiEJSPXJnYNaHFULv972nFPUysX
pAd0/R38dX/hSYExkYS4wvGqw0l/WHm83c2vbhiYnHpuEYnVgdWVNPfb/f+8zd/O
UyYxrL4tIrPtbWdjjOPHcVfvY1aZF/bsMMWWoQJu2SKaTjE3GpUEVjZDeiriPwA6
mwCIq0Qb9/wFJVm99QUi8hr/vGcly56X09olAJTdPH850TMZaRmoXTXpajxUpCBY
18xXDYzHWyKisgPPKJF2HT1xCDVwVC/tfAktaFGuo7eOk5NQCLW/uI4TSIftkf95
0VRWUH7JPqiHUlrLSUC5lXKNMvsG/DkZ/f3GwZTXuJeCOaeEdtpjKB6XyVCq6kAc
4ZPmBsDw9mmEMXWGkKBLlg6R/biQGeWjRv7wXRSr90I7unbee3lbfNkigTLVwgKx
TQ4onb7wi42j5TTXO4BLpKjMN3eGIApX06/ZJCxYQQ1g+clysmLA0J3QKpSHdnIp
B7KVTT5NxIIo055w73cxocD0UbruM4aIhplvle1NurSjbjqfVMxXYFJD4jqKkstl
ClywWZLm9qupo+OVdhu1fcEt57sGJFW9q4AXOAx3uJcb3pyytjUGI5q45sRbYtDh
yoYRstHx4rxaCh/ispZ8OrcNK4YkmAQH9lRvP6zydFcvRdFpAd1g6pMlFs/X4lIO
QsfIsViOGcaX591tZz4ySfh58ZXeNUxpk5jc5tQWQ+RTrios7T53YD2/ivN5+Vp7
lRM0ivMMPSfFptpoa1MjVTZD1jtQwBRJgbr6puXeiITWnxkHbjet87Nn2f/4ZDGE
CYkVyrfixq9xcos3UkEaNn1SlWjjKsc/xHt36lNZVjomrECDWMPFofOgD+lQmiP1
lTlTlqOKwVdWWmOEnhbHTlLPEZ01XXhhigE6IFMv8sueakDI0dFgoOU3xnv+jKM1
JV+zRkslt74QXuj2qkHEPTDbKpmdpV9MOiO/0igHzc5g0x6vyvuHPaqf4mnBKUpd
/fTa+wFoScUZu2Gl93GI0/jajFee/f6LZbyMS0ZE9lWapbifAFn0pBr0RA+spr4h
nQTFJwwKALeP9M4CYsV4k8AQZZszKNQOuqhApvWBWK/LQmlmIzTeU5en3pHKR71I
yftR3mPZmcQivwx2vOjJLAe3rEeB26qVEUHWk02Os2OcxdGixCFzp8rHl8waIpWG
pg7g36AYXB1o2mckUAKgRz0iGGhdCaSR7C/tjmPSQbYaOF3VmOyaOphKig8TsRhC
OjMxxxhPU9iO5Lk//IPLPFno6CTt90uoaxU75oFJRBflWvy9YpMP/LuaIDvQVwv2
4UFBXWkCxJMZ82cxVAjBQfy1PSFm1Y9zFBECJ5/q+UQSczeOBEYtVRjKv7GGnIvJ
d3lsIhKXClZEj8qj8uCoc+Yh4K0+YJe59L+Ra26ri7AxMZ0IPQ+ullzWzhAvFwxq
1If3awxSCL8fmwD59V51ApT8DNJrBc632J+qzR5R1di/kzg1KBpy1OInhtU7Bycu
2fDigx8nO2xbQ74GpYGmTpbJr9yjIAl5blJZg1IhmNgoMfvz+wny4cItN2iAjdgD
DFEh5UojAHrdsL55v8/R0PL8ZPssrNbozW8jczLtsUI=
`protect end_protected