`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1712 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
ki93Foj5FzFLQL1TyB6FqxDKGQBfDW7AlMthj9kGSv6DDDNtW1eCqZlm0Qn2MDkZ
D1Xro28rVMjfYaG05ykTImYkkFIVIhO9Baawy6ALayDjQnYc3pEwRtrhM2dS9+ad
fR9KL2zR6ae2BJLC5SD3LpX7eWJjVj8ukLalcu22s8pUOUz4z4vrDYDvcewNOplv
FYLWx1Yme26+LJvNmtWn66Ga/8SDeEI1/SZqsifNb1HtQIX87yk95D9Bh4072mBx
TgBsnkwT+9BXa0ExorUB9iQB7RkYZScFdzoHLdAXIA6jM15zfodeOJ5XQ7JZw7VQ
SZwU6OgtQeGCddBgYoc2h0+Z9D/rcZBNYRSPlWpthFoNzycfFHAEIDw5weoNlSRD
oDO8MgiESgFPfSPaOU8O/rjkpiwK9nt4YP7MLgUwd7Pe0RZTCHULAunR2MEqayOp
JU8Iq81XorYbIrysLMpBkoxEnpIFHisO0erXASY/VH5aIkUwurFhaHMQKMjMB44r
//Sn80RHOCC4SQW+SBJQ+v6Ex+7WGakzkSj7lYRsBCZceRjJdUKtLhKJ5QMoPfU/
aIJUxr6p1rrulspJYMhzya1UuB2P2eJQLf7ulldk/NxI6HQZoPinZUdwwBiIvHXR
koFNtyc3o8o4AvDFv/JSre4XnmqX2yB9oSYvu5l5olYS5aQfNH/fcHpaTTcs5sZ0
wygHSJf9yMc9frqfuWlwfSIXCLHCc/cbYsZM/I6tURTlFmLnhlI9PBHUO++n9m2Q
sSAHNXy6+BN8x9jhS6FG7LwE01DyoQemLsEoQURuoRX0d5yh7ZTNIlkcahICycpm
h4p+1u6VbtvhFAopJixymLLmoaD0vo+uoRUZk+kTkjySadUrGoP+OrMZGj3UG8NB
srnUh2ENrrtnGsdk80Usov0QvnbvCzAsUrx8UMZNIwn2c5vru22ykPSc+zskLsvy
7j6VWZfm0+fReVsliCTvg8+1imNi+53f3MBexYQ6dVzVW3Fve8Emn9iUQWsATz+9
ms/RSTaeuRETAErgL4DUBB2OVv9JxKWvhlWphsZcNrSmZ26u8eiUqeud9rYDgErz
r6lTnOSGuwsZzVUgAamqTYSSASt4sJIrWKkIgqFtwr7Ne+YSbtRScSsYxvZOV4rp
vVph91Ek31Mndoi1zcAwGpPp9810aUqFIW5ivS/z9Ya4JHeGkL1w/5k5DXAhXjIF
trwwp2lgKdQkrbcQ01Z9H3Qx5ATxMyHBQRbRj1CRk+TVvA1XrFjTM9LBiXzCFBgD
oRwaeCXWIk5uagloS6QxuSOmzKUNux71AxRlzJ4qDX0Qy48M+EznIgiuIXSkuS0Q
tNM8ZkkCuQa45Mlk5GVFh8S4fj3AtpZyFWrJWpwLWT+OYv9uUQmWhpfmOTyqtZzA
e3jyNeQ2bWqIRU5iVGpY+IN4l2gkSR06ro8LA+GjBJyj+N8g7QmggHujcS8BmrTq
H7p1/EPXsFR9yfNXX3gDhsek2Zue/vdeWmWugEHnwq1fYtZUOPQJnJdtNCwwe7Dk
zvHTT0jCW8cM0oVWHkpvK9PnFlfCov0wAWHCR30MA5n7ZZGWYHs8Gu0BAk1Q6LdQ
aNUjup3wReCLeAaOXjVcIiWOXc6lvgy1TIMhRozbbetBpBM/HZPqii526f2sv5Nf
/6B732NFxjMmGfejqPMA6S/qz61rf8MjP/7rlYLndu6EMeN649dUKXcJDlnBpb8T
U4becM6Qh51BUZMu+hKxBj/F8KWHA37ijA1vyxOt4sQsQWtgL+whsk0iurr80Wss
eNTUo8Tn1JyEq/yON9Gb3mIw8sUE5V88T37LSAH4IYvqtfNyzaqemY9TvgM7NJTp
ojvul+gZHLsmrEwTxNGS+XaDVQl4srXDgZV6hsKWh9mXeVVYg/I49FTHvm4+TIcd
GHXZdJDo6c9JGGMJDz/GEVVnfMmaAgwZPrWSWBMXSZCLC4z2n0bwDZyLD1AuY7IJ
ooYN8zzuE7AlqYh5CuDMCC3sxRX3LsJxBUP4Pw0U+DNi/HXm85dD4q3ZExJ3zkGq
1ncayIUsgLhQObVa+mH6rtzLhYxCX/++mFVLig1NWnObzN3rp8xddpObUOhM2Cl7
bH9cRpxXdzuba3XVKt3tBoGkBg9zhUoUA/kmC/waoVg=
`protect end_protected