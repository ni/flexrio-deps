`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24224 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
lmOQgIOM5jiJrGbWpsW/8s2WYtKCWHeWK6lW2Yq6jSWQU81uvxzjiZpqW4gDFNWH
l5LiKWeeCfeOwueWpJfOBSvqgDuBM9sl3TMjptghxMOgzUGgdpBsVSpBSTF7mIdt
67FdSpsToUu/+rDyx3cFPJdJGOlb9nAkKgmXh5+SJ8Fkrpr8msW8qqekAvqpH0S8
A8KqWGM0SpIwq/hA89JHa4AFB0jFQ9emx0W2Zld0b8KXRog+sM+lL40S+qsJFSRa
Tq7f6aPQKGsw2I+u/nw08jPC1cdkt7lrDmnWTYGCtF2di92FxAqj7mZFm9yS4Fwx
FE8nHO4LpVDfOpHV2WyxhjlRfPgPtGwB9UPrSB2O1+mosolPMggZ0t4Hst3vexjq
Y4LKBMYzPY7aOABD6AQspMicOs6d61Cg7+iVmIUg2wZLCmfdzgEgbBHof6gSvXIJ
C4Hlhs0adObmSYUF7iFxxDjj3weVJoE6ZD5/thFl+jvp3n5arPWU2Y8EofXWETkp
kR2zoaxfFI2J2H/zXuuhHxMgL/Hdy6U9AV3uKlmkczLQH4fvaJh8v+Fr3WDD1DJ7
ws4KwogpzvTyZNglDw9ujm5qf3VJYjb+Dw8shKivHU+Sj2vRhJIw5a4wh5h/RgWd
5Ipu7ZINawW70kL07q2jfsH//9MDYRF8KfR1LllzvQMnclNIqQbB2prQ1QpM2O/a
3o8viOYzAVSSTbYHsXUjNSF4ODLmfSU3rC9YGuCmLvvT+RgTTI3+LRmfg7H8xuM7
FaXTd1yxTWvADjseGMawqnJXvrAD9fo6guMcc8xnXWttHnyTOFXLJVSLpIMdHThU
Kau/als5Z4UMY2t3s0+cVxR6UTlke/dnyr8Rzau1sAUGfjj8ftr02luuGxXmDcWb
1Wr8yBrLUxoH5oNiKDiJmPQkBajOOVBgy62InyIQ3tulALfPL6vn7M93xDcaBZjm
Mh8C4tIWYpniDvwpD0W4VAdnAm659+Sxvyy3uqh1BS5Wxf+nv8QudIM2EfT1por3
QmFdH0qI84mxxdcYyBr3lTKw4yZSi+hfj7QVCOlOamnkoq8bnk5CSfZc9LYdbEIo
y/F4VgrlRdwAVydBXTV2Q/clIpONlJAogE+FtFlHaFhKhoLYlmDdjdtOiHNlXUWP
e7EQN7BSBunYJMvy9+gDzxTCBV8TvJCqFLIBfyknSpoO6hR+Ovo6M/r8KFs8vvhX
NvWTxl0OHhv/fBqjJpv8WNprl58S0z4wrhKg1HBlPI72e/NOduQh8Nxqnjs8CAr2
sF2CCQHRVdCmB6pI/k0YTyIEAWuDE2bccvZRqqlzBSPzteHB3eM2KTgdJY/i6jnw
UeuHpsgTk2VuVBhXSM58phn7/ut+VDPOwlNs4S+rqr3UlcwKNYrj2EHOFcMASGS7
VEWm6vQNbxe9R0KVeEbbZ6iijyTI3eEKwxilnG7xSUcc3vRcmKnzhQOkWt0G2PW+
f8AWgX1pO/u8AqBTrBZ+CsIvESmVTzXhNNrWCQQ5uVZRTMPWHvVhsYuszWH2Ms/e
bcjveGAKOhnzGxaVtas/m5excjwQzopm3FWeaSzm7ZdQU/Iwn0eBV6+Cu8zRjwqb
Pt08tHL9FjiF91fj2lgWCeKaVEmIWApdRdIby3kKMZqFJwIwe5n6QRO44vD/aEyR
E4cXeHaTM2ZgxJf2YD6IwGTBd40pJygXSmREY6oQsOHMS2LjljoAC2dQ+AOdEV8I
O+TVk2wxznrLYYwAbdPbLRPDX80y34D92e0/e4A5S6SQxHj9Bn9uE8x+8Y7OVdKR
Y63rP7lkf2jxhL/zP7LhRKfvA2f9XTi5LzGElW5r9zhysvL2HdX1FBKPQ/xlqx6R
IkL+R9nAQ1zlThlxMdhCHdT9QKByXtwBt8Zp+k30Uh/EjRxZaegf7FqFrviJh5ol
vlqFd5y3wu66vtzOQpifvcUGG86IQmRixyjZ34yrGNqWEkU2EdZRdRpRR1srU+P9
oROb1qvSLX2EvzX8R5GvesfImved3dO2uhTe5UidytJfiGtKK+oAT2IqKS9B/Jy0
8bnPV8xMPsxv4nq2PEAHkKj0CWSQT61eflzImTtw0g755lz9oYfV6XgYm/NIP09F
c/4gD6yvkjkCEd0SUXHZrGvQbB7QkGMeJ3BpsiI3SA9J+UXZqQxOwxSYKEXUqwyp
C/SZXCalfSEbRcsK6UWw8Q2oPnuzqkClRpFYg2u/msPoiAW3Q9puMOJQmyvoln/+
j3sKpdbiu5Tzkv4OyRv23SCHke76PmDXkeC6lV3s12/FE4WpLwt2RegxQusDQQWn
+FFo+7RwZUQ7Un4AWEPqJX3XujHvUwE9cmf+bbv++C69go5dggte1ePRIRzRCpC9
fhuxfUR1dVIdQdTwuYGf0ZwrD5iUp69wckoqxPO/O+G3DFE8ZsmJhL4QDtQ3QASW
DyG/kG1JHuuaEYPFiLVOvlcn5h7/ShoS2SLC2JqsfJlrRTRuu4avHv6CKpzhMsW3
nCk+/lYNobmE3bGaWEVpf3/2hmL0zSE5N7fUUcm2UDd3WWkPTwcIw12uFBaoBq1P
ePLIXNxZ1OQXFlflHFXpVghy6UaXyS8WkMNKZSWohK1SeYZU8HvAxy4QoHi4gCfx
RiptOXlzUQGTW36HPjHEMAfA27Pe5Qb2fNdsk9tgI+7twk3F68D/kdmm6fXlzKNZ
h3+952RvkW45uC3ruCh5t2vsUThkVBzR9CULiJKgFFAsvb/zxPfK/yz0SNkGE18c
azifeJOGmOwoq39eDtN/oc/qBu4GI9d78+b+QTOBcS8Tr8YapNirnesV3yomURwF
Ipw8WvKKIfgG6XuiJsvOHPT2NqQIXU41kUxxpZBzFMDNa9SwUguzqSp/3WrV1WZW
kOYBPlLe8N2CRi1t5WCQrTA+1p4DqSZiGQwhReKwaZjAdt10Lh52yAsgP9RfSDKx
FNg+Hmh4oXAJO781SMjO1QrZa3tOtQxy+LHekiccbsBhBTUMXXmlBb84azr7tYd3
gEOQumDfDnVSG2QwYYql2NZrSZrzh2IC/wpegpIJo3F2M4V545KTj8OfQD8ucALt
TLwCWR6XslLd0vio3FUWB0MAlLd2ImEUt/XlLqLWRsYY9MnOXNetyXAUhFz/J9Uz
mgmkkzISTRNmwkXxxN/jjR3/7CXX5IpxnU3umqxWM8JdH0jrR9KaL7Eomhoyjc73
jNv80UOklWZ4RRIAbymwO/bvHxuZ89S0KubyrAfEA7sCorB6nliA8LIIZUa6q9u1
sBkKc3ZrBA0cxDEZWKFdZqXaPR/sQLQTPG/n8XNiCcldh7l7k8ySlRQ4DcE8iht8
somlf1iin3LXwgrfPoEU7ZXw8ZQURLUs50OT6jD8STWILrRTFKfNnRNPyNcWM5Cp
y2CR99ElrM0ZXnkxp4mhbQpdVItRjTG/7AvSjqJBtCxjEgJVsZJtGp6c9Dzx1BFv
5Oxc7u+xO3fhYvgyiIymzNGQfztEl619qMeYl0XzRUjtD4Yr01Ut6QiUmWuOS0nf
mZfcKTj++X6iceB+qxQ2rdfMMwCZ5vj69//YsCZINRlhCjkRJxnAy+TUcurwd9Ut
iwVqPDlyl06GNOjXRan8CRhUlLecv3EU1URy02Fx4cWddd1lsQTJNy3WIYy3i7U8
DEeWvCCFJqkBPdb1jNnJJFzfNKBngo9XmZ0+s6Ts7BzUsRgasACkfirHf9hxxMWZ
ZnNkWfkN13k+Ik6ejm1yhBME+gI0AUAOgSuC5r7NFs3aI10hb5A5WNPzOjyqMYLR
y7ulvtRkiOZ4sclVduo13UFwtP5awFl3R+AORVV48XwgeKFjs421xzRHm+ndK5lP
LegDg/TURtIog3JKRkZ0+XigXxk/TFlK6tG2xynUcZROdQEh5MvZT6+DHQwfywc+
9pgPyo91GKr/ZZvA5c6lo+dTK5aTTWGGb9kcrUWfRETs+1lfBcBq2QqvGqgt0kxU
b5MQ9wHar38b1tQAdbFrWa/jtdAF1pUgbpjfHfK+sLf9yqSdHoZNDfu/ZJQEtzIA
nTC7xDBnc8CsrTI2DLxsEpcIOzbHF4438XL/kyn1997UR6tqIcL5A2wbbm4DATqo
tlMZHxskWoOjm0nacpcLuuFT6kaAoi88WdV18PeEsXeOHzwQlzPdKofAsyrgQi5/
DRDfZbl1PBZNkyRD+snOBmd+7a8hrKAsOlSuXsBKRV0JiwuIcU0bqqZ+FdV/2qc3
rEDSV0hqkr/kYoj72VsN2tt1aaFPV2ZJNzZ+Jh0KK+z9e+PyQp2Xx4BGSLy+kOcz
+4rgBVRDeTdynjoB8oSajLprnrqs/wQD7XUWZvUzz+ZOhuKni7vdkzEHDQtC4Bjo
iO+32zbsUz8ZunQbcJrSqvqIB/Izu2MCeFZODWVk+Udhpo+Ysem+pQQQfAmQgrVG
7qVxRa3MBURyPKnUMgi20ArndHGjr1K7eY5uSJZokJYef4zIFYd/Ze6jwI/AAvBV
hFHVwv+q1ZPPhqWvfvPQlhqpCppdLEX1V1EXIJLZPnqJSvauRBCrb2NXj0E81u9n
UFUVACZj2l5/gDnR/ZaVovsuyxZrwLI2HewB7Wa6R0mc829lrMn1H2fH4HXJw/b6
FvpaaqxjHZOLAUnOFyVkrbMfOQVYyPZLaKNZnGTAEahFbL8tOvdzBRn/hfUxL5qp
B/OcXe7oJ+S6YmMR3hlojtYI94sN2RpcqHWmNW9cbtojQ9uSnRaPAWg3/FNdNvzm
A/YgjDq6vaAPETOFZ/kSLwdrD5UYO8Y5dd/fHAwPrLWaosIpaPxUo4rqbZ1uAohF
Vja8F8aG7bO2/ubcX5jz/dn+FxNu5Y3SQo1VJO/UV4pC55Wb/ueByioN3KC5v9gq
Ka9p2jG5okV6FJ2s7CvvNOSdsRKwd+XehqYkOImFi/qvEZ+C/YuczxeEsOjleogL
yMRvvMohO/UbLUlY/1Eu6X29iQccl9fvHuyCCbLDolCEIRF/GTwUuDVIFY/7Fnwd
Ux4UAYdYKsQI5bDOUk2sD72X10JLZeXAGVmbnDb4h2EPXMst27jhHMd2BdaVBph+
BF8Iefu3Gh2wOPAdk4xM74tZ7gG+LBVqkOfLG01Fc5BHmie7NpxBaKGbii4uifAb
FNOrVecdqMzy7v28EF30wuyPsDUh6Mwt7FSYfix+fkHEIEcCpxHJ9YwFRRJoTIA9
DJ4UFf9N1NQeFw+3a3OX2xREZGe16uwZgkS1fDK4q77yxGrqLCRruM00L2rYvD6Z
PLiylPTAH9QIKYz86vudXfdM8WUaPIQmrTusKMu7owsIvHokojszg9z/shitgj4N
zrNdmoah0Z++YZi3orizwNa1ePr5GVPg+UJNiM8ucDQPky6/yRe564aRxLqRnjwb
Mi/VgTYGdtmGtR2JhniT+7GTYu3qiL/qgp9adrFy9TGR93N01oQlawal110nXe4c
kaluB3jzyR21LRglibS5posLhAScsFrCPx6OEDHW2dxirZsS/uP0VU/zLMxQgAbZ
2UwR/N6bEpI1GXP4LNZilZQi32FxBimCfrFZud13byNona1XI//5/ZuTV4WXDFYD
cc4uLPHXHC7C0Sm+BchOaFJavMEJ5PJ4jXqkYgPbP69ac8FDZP8XZLKso4jOoPTf
BWeortTHiVFdUXVSafxlZqmxrlY55c9pV8CixeUswUfaeJieeJn+CBKq686WOk82
e9nyUJK/fwD7u87M1Xu4O4cPMdmnHBzxOQcY28CRkUA1RKmX+p8AOMf6w2fJzW2b
7ROagRV7eCfb/RYwn8kanr373/7/rcDwXlMT0g/WdkJa2OBD2VnpbMVI0V2qtEb8
O+YZDvqxBH9l5NxTOAaKTFb/KJ+YPt08O4Mvl2NYKe1nB4HoLj5ztiMe8G6cvaHA
M05bSftNCsCdWh7S1Mo0+EEzes3wcKxFR5ySfY9XOJrIaCCGTIqwksqNVg4zFbzr
gqk1Bb1/+OnwB7p41pJ1mIjAZGEc9OT6dCE+lCP6SwfAEW4trDEMHac93g923d0v
xB+eSvn2pgYVG6R2c87FFmS9isy41oJ+M1CBqStLUrQL4HJMoscYhdLDhDg03aqS
6b97cnrZgTL+oPAwrrUh8W7oHciH9DJoTpR1cmAKaGDZq7jSMVHly3uSmbY71zuw
XLsEE4AD61zSUw1MiJic4nrH2jZBT4zBe2D2nLLsSWhLa+b0aF28ZUKgsZwcZN+b
tFxb6y4w+VZLk1sx+1QaRruhmQXBlY1XnXSPCqeGpnLkYZpz1QaJbfM2wgak/vHj
chs8ciTAS8ULNlfzav2G/ftd44ucO1ICs9hByYQXUH9Y+R+8tveVHkq31g8Knp73
Oo27hk3yqYnsfMPwKaerAHFjSuVBZA60/T4LM6ocgxZD8o2c6/IHsK6xTb8OgU43
UkywHrO1yX7AZc3f6JL5kjLulXoo5DI5wKYrDjzrYY4UaAX+JxXfGVj3/8rXxfRX
gXaFgm0Kwk29aO6uQBTZ6T/D7dxWJtg+rTzUWH7GIT8F44FDw5UV35i7T+Za+uDC
goH/pyAW1ZCG18eRhxH+iT72cove8Ah+tnNKbj8Er/n4sRlpBWkVwMBVqY6EO98Z
jrl+KiNWcRgD5A8e/OIzT+1hTkE8ph375aquasKNAABurlEcZifS3+99d32fm7w/
Vx4Tjuw6uph/fePBdxLObIyeqIeYepc2AYaQu/HZYInRDVEiY2jin/NI8Ip9JrJO
38VaIMkuC/n/41CtB25bNRumXU3ZLUQNA1wLP42PuSLgIU3dg3W51lc2vUComBTO
gR/kZ8j7PNT0ghWIa+cY7vVAcwr9LxMJ8posud6rq2uru9rXP30tgC1pJY0gljAA
wIrz9AhMulmmebfvuyno+slK2h2HKsujRGa9piZtxAScPzeKcBTeqEyacTvJ/m3/
d0BLWcwyn8dq5I7v2hnV3tORy36PfKmfvE+PllkhLn/g9Uq/LcY5B4goO9mAS5ZQ
cox89j40a+6KjbiNUABA6H1ms2+VWA9V7pdq8nPwAd2q18aJwFORlpq1VMLPXrfI
esdO0O15/Z3/ElnK5OoIA5L0E2brJrRv/rT7geOxM4tBDZW8LzVs6GWqN7xETqDl
4QOjM751u7/6QAstwGaApPqvNtH5BxAaGFbeIJEq5cq6PhSI7q9zR93sjW37d2o2
KLkgKxr/cZxdKEAovY3/GBF7N7IpGjxRoF3y+amgm4YzqlWcA+LITlVFm/kOTu82
Gf2ekAK7APcCtlJR12sFU7Wk99VXIB/HSMZ1Tj58o9BT+00C0W2XEUVPLfErtyiB
X1aaEYCEtbibFXevCkfscP7WY7JwKHw2XwnUZADhT7eakgHcOehIvxx/eoBa575h
dwq/ItaSpqut5/roV5z0lF0WG9YfB3P8KmzYeRFmTvM3TF28oQZcvFTA7SGNW/1o
pfR9xEgJ7wMgo3ncj780j9Xw73RBRirxOQvjR0xXe8OjTu3ssppHz9HNTZbXOQND
utj0npvDjjOtOl5/YFYPF2N8pCkH/qZJbdjR24HtJX+BtrdOMaMNq5ow/pzRtIKj
TLxDS45PjoWQHKSapCJ2eYS4mgAxc26STaCQKrm0hgupmhuL5wQ69wya17Gl65Pf
gYdCn73YgnisP7CBHVC8xX6y5kVxoBfHJSugBiYVpG6z0YPm38IS6j+YytoKup5y
EU83j+kawQkfApEAX9rzfmmUb3cENgVqDvh4zG4NPRg7MGg+9YiaWwLfBNfuRUSF
28Rfbkgj4yHyEIbglkF3Jbcowcx+j2qg0unjSEHLbopn9LA4l1Ui5+r2LKzCGPEB
02whttWwg35zMYw48SJdPEomaFHzOCZ2esfAKXpK6ZGnu/+rHHC14ADlEINBNjqP
Rt5J4+nGtIT3pvEOC1WM/e4C4xuTKEgqG3XhJRazu4ayzOuD34w/jOS1JLG95c1H
RB9OQVm9VyvkThNEsLHGiqPMpFlJiaTLSJX5vFpEF3/cH9+f+ATLQb363FlJHGM/
heoksVaZivfoayD7bPKhUKEtla+0YRHR47rJ/fVryY5NvRh2RCnc4aFXl6hUfbQt
9lWRQxwfUrDE7W43B4yeRZkNCvELl/FDmqNWjpcx3uNZ6uEBh04uIpjwC9jlBvE3
TMJbqigdG/ZGCjtKyzHGs59ayEg68k/6jJZCpKo0/yQdZ+C+TGwyM89O8KNQiSXe
Gph0w0YyIn/a2Suy80U2sVINOB1MwbTbSdw85dz184FtxYncm02UyVOPBVgRLb7E
1eigGq9bI9I532sgy3FQyuCnyquucDu+R1MF+uyi4ZFECjIF1Kk8R4cTOafsG0bL
iCP0SOVR2V5c6v54BPfKjMry9Deja16oWPunOaf+9R1YSR5jnwc4Vvb1dbrW89rK
ls4c+ma583HEDtBnFL6+Q/Pt7XXkozTDcOhpnJUoq6B1aMNHPQLk9VtX6Me0OYiu
Woxjab1A7JOfPT8HxF2i9fa1xKeqosANDHeNvc9j0GjuKiXqmjJLFv2rNadBhWE3
4Kep+iZ8aXolTsr3LqaNbjRF5Jl+knSO4ufU6DnWwE1Pt14nFZteuu80B2DEFHqg
NTtlJ+UO3zmrPGya/xGgYCvaJL7kd54YAdphH356c3sYutafsTpRWIu7/zkD49tu
Ol51n6RGVDKHX2LMx5yy5AsbxWYrBg6aZnn14fyJmu2iO/Hj9QJ/siGE78UCavUO
rXgwb4hpXHPrvIKK+un45jgsilTZvU07E3IdegGTXIOovM6i9R/N9WySu1bJ0xha
4bkkVVuyBG/84K3zXIPS4/x/SWtYNtAjZZ+qCN+xOsf/S+9QwK2UykPpgYNerEQe
60Xcv24BFnS0NV57rMYIB50o6Pq3iymb93a+/adeyzX40nvnLnK2kHZctItWSo8x
CjdWyqJk39pf1Qn9wlY8z7mhvBZIm9b4F8zsuasI97icgwBWgiEMmEMQulpz9pH/
+pZqKvvDVsxNZa59P7eI/3DL8yht6bKMaR838kwsNk++Cs8W9Dd3xg/IhZgjFxc8
uIPfRPHgDdybSCAAFrhhqYyO34olcjdO9mxLc9LF50MX3MCapWjd2RNltIjs+1fE
6CvEL2h3gIVA8Fj8b0wPsr6OOXSg16R+2V1OkW0TsTS7yepwhHINyirCogsp1oIz
wRgOWtCpot5g6LbUf17etDLGmUYuuljuHtz5UXDDO01e/0cVS3uufW3XbQbzetsL
a9A17X9H/wa+Wz3RvD2Pns5rwKAoaSUB84jvtIPvhdMyz/euGqSd+9B8YeCcpkXS
m71dl5V12aJgCtqwRHahJMwQWAs5k+pBN1oxmAuQHKTqS1/+BxiWnY6ePA1JkFQm
UTfP12RFKcFekKEHPcXjJmvkjRFadJKn5ZwgD0rgGjtOIjYgyn40e1Oxr+r0Xgsi
axSVBtyEbHBIADgpIsyt0mwM/K44gmmTQzrLDGBUkCw9pYSwQ0rzdbJxMdrpxq0Y
6JI8/EDpFeQcsrEFXikC85ahniSkt28Mfro7eqSK1vcAoTvs5aqgzXff6TR57MUT
YEm0A4Jk5+lMK7YJQ7kLOHhP7IlvRf/h9gzZBK3mUlEAgsbD3amvb+idvZVIM6jA
C89jTKfBkh3/lWZUKetETXqtJWvhPgQ2Jg8d4I9b8CsgufcV8SXO3kydos5BU4UT
25RQ4GtbqOZrJEPIJisfNSCmMWSDItNxaWrvq/65J+Ht+DTCp8nAKrECamLYzc6k
0qHF8j8e3P//SB0FL/idEL8DOkIro4C9YzFe2j7pwR63rvGDDFa3N/AaSMv5wklW
pp6B0APIiZiwLVDxAkACzeQ8yg4GE5JC1VQgnUj6e12JLm285L/c4LNQ0+rDq3p5
yImkhuskhtK6s7scSsBE5sadrhAAWsJy0acqs3LMzH630x4K240AwZhrUw8vaQH/
+DVSPzshQxVllpNf6mcwh6DaRFEz+b8nE+CtlrJl1ME69QHJNBABtXW7vY/zzsJo
qmf0+iSSONw2HnBpELvCz2ZwQZrCjMMvtPfE6be9rlWlg9HTQwkzbJM2oygg9i0H
LH4y8VhG618oh++r54Yttsq7SYXr/xCEe4omCBLYJDGqZnhzHkt64LOQ5GVMuViD
7E2jRj3kglQ0wiDlEDd/NGMbojnf2gXfVn9KdQIjovKbxNQJ3zbms/lrGZNdugoq
K0HfaascTmRxRgoO/WbA7YMmfOB0qFj07gQPAV3RZcruxjcHwRForH4DYrWYnVbH
HmtcOjRIf01Bf/UDNCw4TEfEqcci85a+S/LVmXtKpaS+57venk+U7D2cFLOORFoT
bsFmA6OXQr37ZIX7Umk1bORdTr7d1oEMN0/zOw427xYXpc38q0hBxYzULlinqdPH
vzchYWe08HLov5nskt9+kp4jMYXrR59So6t0gFDKKJayAvRlcgYeQkOi3Ju/cmFD
niF95bDKNFH3xc5rNmujhDSB/q69vFGf+LWiOXOLf2v2u4iFWDzeC/IKW4VV/89O
8cv1ahdpJFA91ta6mocczCKmrnPiTkbI//t0lL7e6AqvkKv0sygsx6giw+iWKdXY
WBCpSNzS+7vzWy7eUEm/0S3ohkDdKTqMwCzKM0i5lhQJ2dZ1cV75k2/4J51tRJP+
qc3YCLnVIaNiodMYML99FNAr3W52ELqKoO68WGeJ86YBgkRe1zPZScWQDartwUd7
i1P9VqL4lRyuC/NFiB+OVpanJjvHhVYcoqXuiB9YhcwV1Oc63aMUcC1oMa+8etFa
IwMJe4uxHV8Sq8hqEfGDL67F8qNMU+1o12ZwSW1URW4fhzsKjIM01voJMlGu6KzS
G0wzzs+04rjKUlX9D/KHoPE73F8CJMPblRpLbuQ0BIVSIKilp0bHL5RFooyzjRTz
SbfUU2pLeZmi2+sR6/kmpJ49BuYS4c3+3mdaKGOfr/S4R84FUmRCB3gsxcXVMe2c
9Y8kW/rlvNFgq37rvY+evJ4UPVFPFAVS9Hse20QQl/nz4dg36LA84yz+F1a9Lc6b
Y1sGOK2lV246dQAmcmVAT3pC4fXDmvbFnt49ELzEGjGk54vIwJj+q5PtcTGDD5Ke
h0g13QkL5YVnQV3y9nfLuv7tn0TNJQM2DMoOU1S/wbq1ioU4YhjiT55NXaXF9vOV
CgM5y7ULEWwRRuAqt88fLfAE4UabQ528wLt0ahXwUvlCEys92HJ5wNsn4ca/khLA
YmJPpbGjkI/mYzsIajZGwJ49aO2J/Y12kNLrjbh3pID8HZhxqzHvvgqbLpe39yNj
qgEy7BsH9QdWgcjRhXPIBr2Nyhaw7USq9gKTVSK0bqeOEwnJ2RlVLKAgh+PAi7hj
3bRMM3Pi61RIwnXCpFQlovHNFkauUVJyBkSVBzAv0nm5NcEfCBLiFgnJmUfIOv5b
UzhN1ay/pkkp2+P52Xn9lL+ocjXk1wXQiYZoTOhTGVLqHBXsp3m/YL6eblPp3Mr3
73QQ79i4NCiged8uxIFzB2PzJhMi2xvCIRpgVcGsW2DyhgQG+Mkg/C9LAGUDh0ZY
HbU/lSeHaLfMK1vSD4Ln6nDoHcbHvxP7LyYNgQ+r2fg2wpUOKO4oL2QVm4xBql0x
3LC6WIgtfUOyH2OmkhilKku1JcP2wuzNSJg9BaxhmIPWCdQsriy4ZX0IrvKB4qNB
gKs37M2feF2uNlbuha0E/tNdS0+aez54mtjE4CrgBUk5A7/CTH/w1NllQhKIEbfj
JTf0v4/4E4oeFnpXO+YB7WoksdF+vGGMwFHyoPu7Nk9GDeff2raJRr0y9qH9ytaN
FCw+u5SF7l1Z0aVCxQtPZqi/6/Y+Uu2dG/C++8qWXMxWyfPflhPEH3x3sfJWIZam
ya0rLuwPGyw16ZzSWrThbegTqqGBro0rA2BQs3rVwfuacSr8L45TYVjSGzoNQ/a8
8TLXtTp5jFgfJrelWq33QlVSynDfMtXdNwqk5BZYu3JO8H6KqIG256MCv0lFuh5Y
YQfQzJvYe3DWODym9g3Xc8Eik5Dq0C7FyS5TXmB6AMRhrTMMpUzLZ2WH9BzlOw0E
7F98lP4Vj6PmW5W9sOW56xEKdxFQRK8EcaD5i3AeLvgr12G+n25YoutNyKklY/+a
1f1GXio0TRXQxINJ5OXuEgVgpuyz8gpUVzQYjkq1LPL3SqCXCDwW/PgYUBzJ69F8
9P2nyUSgAT4GNYFKCODz8z1ez9v1g/Pth0YANh7Enb1TmjvibdjgLCwUE1l3Ya0M
VHuEVTo+1aCVD7gzVTrwVwVjK5g4AdBNWKSqq+qZ6ND9ih7vdjSLayZjVcvEHMBg
zZRQkOYV8DYDNUfe9uQ8SCYze8atfq2UI63pTg0U087gfVPc/03Cx6YOVakuFe2O
A++w9w53I3NU8NYJwDImSSsUp8m2SKP/gmOKokVTOcNl4oP4UeJVIC7nqlGDzwaB
1NX9EVTnDCrbVQE3PneZUYCmw5hykKzsZ+YDgqqzKnLt2b/peAjahelsdIBZWgtR
32vqyEOb6uOGk9j6aSnpPFuT8eUIFi03W39/l94hzz0Ab/5ass/r9TWFo4V0DCCx
/hARkCie44mw+T+j0/12Wxw7xo5Ka6g0vSQ9ygO4zAokGxOL6E+q6yGLZEsIyBn2
1EmuW14X9M+WfZwaKr1hzezdB92ugqywrAuJA1IhnLxfcSa/fBdOMkCtdp+S5ZeJ
U+nYIHjWMKzbgdLYeCqEZXnRonZH5y2dv/YaYSdfYGtTZLFDBqKn3ZgUYjlwXMXf
hS2VO8kV7ahlXow1lgRI3wjNaqd+K/wbXCCpmX8dThR/l/ddmF4375FdzEMb406v
pCRhOoBea8WD+DSZga2VgeMUyT/ZXBYW9QPjFwaPZP8qR+wKpAOz1PJ8i3Rwz+B/
FuPLWJH6Y79W+pHSgt3uV/UQ5YeVNlvKYWw7pqWYjqbwzvW9KAQRxti/Cdjnvsjj
ThDtq7ZzzQOERWnWbuF5V09dnTPhTR2nR+BqQqIxITfWg4HphAewNHSANazpKPXu
7KJDis4iopqQgNzCnOcbNPumeF3OV0eA0ITa8cPTb2BOy+8TkY/vZQDBuLVTdKQW
7mhix1D2sXQ3E04cAAOeqfEsElIcciFMSfyS9L3E+8KTthi8hHlmhKtuWSlXeqrI
5zF5iKoUvWAE4KVDDSSA64CteEdFW1CKapJFwYPxV3+9f7ivcyQoKiQM7Q1KGUwZ
LDysNLt0/iWYKjzRhx/0OWmSTR0H6DXbbA5lag1dECcvwGFvI9vcqeGrVr7ZT1HD
ebutDeHg9w81vG1JPK2R7XlR21XAYmPTZFKK7JypBz2mGAKIkUXKPBdbGrV8Mk/6
qZx7S9TRAYidi7TrceuAzj/moMIbuYPwjs/auDMIePuRgbyD9nREn+Yd/J3ZnU8t
u7kqsKK/xHMSnrgOUOB+ZpB8fEVK7E1Q0nuFqxsWCfoT1mXCa5PzoUVHhoA1gzRr
fe+pHcUol3XvlEdz/erpj9xujuIbYKSrBesBSqi20+Gal1/zmXZW8DYY0+Dl24P0
L99bGjy7X0YEQhZHDnBIBEGElHxblVnzm5gvnppxXvpZG65kmg/f+xT/trKqy+qa
0bJZMVAS0ofzelGWayFK54q2ZddPokRCtwonif3Yw3/fPlA1bKjI6wkSApzDBezG
zFijb5Z7IAbATjNcl60CIkcFfsBbvEKOYv7+ldciYp1Fp31QnqMPIa9zReBfb51G
Loe/tY1ZdunjMaGbT9+UGG5CmxVFYV0FLChhk+1XMfH9RJqPIlPONJbIVGj9oLYG
xNgCzPh0X0PgAgsoEIGhg0EqWZLWsTxY/5utHqCJL/A2ZucSKOojVszyR5MLFjxr
VUHIY4qGE7BKQAaKXR1+xq4x1DujEkDZeNg+IQXr4RJ0Dh4KYS4VoglUTNegGZ4e
9kcVvgDMgNRX6HBiNkajJuECq/Jw6cc2Uho7dQKo9MEEL8ZvAxkQcG7j+ANBeHYA
VCvfIDICREYl7naVASPh4mTh9S7xiVeRL20YxqFBGAzX9oYXNY9JO/MoIpo0LIcs
v053Y5pVM6v6yJwApIm0t3pEoz26v1CzUr7CLV/fK2RsBtrwBMq9OCBT40zAqQFt
tr2y6FyTkGd9fsCRoBi0eqD2jRukJXGBaQUwK8eNZSqMIYnHZrp6OAuNou/snm6V
iUcn5NApyH8Jdy7ZGAgMw3pHzFpaC4Y1Ijib2nBTVWx23hqokAdWHERY1d6ihDWE
57Osa8mcdduHZm1lxg3osIssQRVYMGAoerstAQ72nIyu2pPfplO6iFiVz9TmL7/+
hp54U8FuV8PelGFASzynEUK/6rKow24ayr6tyL7DB2n5EPdPghYqgU1l+q3d1/ZE
By1N+xWHpTvxYP6FapOcNC+sCuIquhLA6ObyGDu9Q+Tk1x4yGPJjG9V3bOd/NrZg
17TayN+U3BB8UKHppI5kDP1oWxxz7eAp4TEbpE8oL+IZ0++FKT3PkXZhdJ/NZlW4
d/ZxUwXp2qYBZRnMPOHXFE9MFcDC1gqyFWR273TAdeoXPcA0nI5OOotXAv3Sejof
CM6nsMeTGR2vk2LXSg5A9IVVxANxQzFsJOZdF+sQvlzuhbb0bmEYLu9keac2YMzs
1QhJXqI1NyrJEBC3WnynE99AXFhotNJJkuSBg9phOOTAlLzvdoDp+X93jh7IePIZ
ZPH9Dm7jB9LNOiSfkkOC4tDzE2krkXFp4oYFHRySBtGmjUT8fiAA+J/DQmjpl9SI
BohZYEbJ4MVgx9rwg9Rn9naswt/oO72iCUZtxewfvYLweqkm+YQQ3/h4nQC2J/eG
92QtgxQ9HtQ2AIR4RjbSuo4pq6wmAkZzzA3LbmhZjQV83eIGf5GrcmWc+ACZjMvh
r4E7WYlSAB2y8ZUXfjs2xOMGGgXLLnTD1Cd4QjbrtWrdadsujs8Dhqw2qIvaqCyE
mlPjPrqL7cNdU+oHdNqOVc/qKeMUDhXg3ZdeIh0ACa6aG4+20W7sIW5HNkcggTA9
dvx8wmVRgFTuXTzU9CtY4KVdQpVGcHcfAxpybM0l1UCRw54eFHqVWzjjpKm4SfYT
cgi5OgyJUDL+vV2s1wgdIM1SsyLDtnJ228oxDxBDD8F1e2vMW9fH4tGtKrCmnhyJ
NZC02owS4Mg0RdABkH1/rxILanUdjGBu3EF8cb+TVtOjMrLdMIFT5XQvxQzEpZqJ
/cSAHY0/UyhGXbSoQnWo9YDidNPZpzJLVrodG7fZHWAcb9QXhkB5d1dM6a/dBn6L
aXWFfLQDgDPXGPtoZ56ZOEpUT1+GpbaahwC40WN4CxlE/Hiy3VaPpFjK2mhpXRmV
fZgdcY/5HaodmYfflOwjIsc13dEHCOxgLPm0aFTUb2YDtq4BSxvvVFlAHyj/1Omh
mtQrcH1gTWY668AgyD2MkzAu6zxmPgt46HX79HL/IaR2qRRVjoltm7kn9AbcVmjq
cgPeZhNzHrnIVAA+g8VN30uL/j5qJBKDi6U/OqI5LVs/ENeixwgfZNKVac34nWAM
LQ80r0qJQm2BeqgSaVX5Va+sJw7lbMUQV/csRq5RjLOWcycCQsrUA5hh3L/buP5b
FqwtupTBN2nfQ6X/BwYcrl+95oPRdkai2ubAWEGthCWbewfPSUxaQqzWB/6Ye5XB
tXC0xxqusa5LD2LIcl0QGsXBzpfm1sArwxoPc7CpiLWKD0IXoGGfBXNV1EDeuUdf
M/bHe/8H9EFbGxpriPLQZXfjCRoFwGAj3YbGR9TmqNeSq0LxMgcbQEvHfTUR5XRE
bdATViDW1lbkNkAFwl0ldUhpFtxUew9Pyqj/ylI+EYl9MRyy8Oo5SIW4bksRtKH3
V6FCcTEYJz+FNYl1TijjvjS2CyEc73sV7oEfVfWa/IWfR/tI3Z8EeZwKLhEo5SAg
qsVfSMkwLGv8JqfsMNVXG3vgKcrAWngBTrtB/r2wGJrRTYUYzseBBOMVv5ORrH42
fy48VC7a6X8xi9kH2da4fHObbwyeeKqutpjthJXRdXgt3s16RRva0SlYg5rxynVS
fPY/48FSEwZSNfdiU4hN2KTO4l0D6JOaM3FH3KkEgucdSe1UNN2CHRpfzSQN5a7y
Ih3aHFGLcHLQ/KiwEXto5ZqbDJynx3mWvOmV9Y1NmePly+7kdi3zih1wS83e3hXO
xkmIiPaa2ZbMl5omp0LsZ3O0hVUv/FGgfBnwO0a9y4b3e2cHo0l3RZfV7BkAlh3l
DXbzL3E+OmHDqiJK70924gseTjTZNgBGSlSqB28UmYNWokqQnRZC0CYw53LCpQYr
PxRoleXf2e4DlAX9W+QwAKpnHO3xewz0qMffdaNI7dOhaZMdbwCLFXqRhcsFld+2
G8BB0lBHnpUCKhKs9Xb0KTmn6poOJ5W/ZkJFseG5KoeP3VhPS678IJY4Q70t9vV/
PthMuQxascFufC1FYUwAGQKg6IsON1kbhy/Xf7MYMjKh8mH2E7QPl9XiLs79ml0J
mlnyYz28o4VoQnAp9Ih4DoAlr3wzkyHxq9KPiXedA2PYmonD/GjlRxnAz7Z1ntdj
Jm9y9wz0FOTy2NEFEUYXm7bP2eG536Zw3T0JIIZBEVcFMIveDQUUDX4OtAvFCM+Q
NZPpteH1mbRKAzVL2fEi8xxBTDlQ3iEtaNNUPy8qcA9VqeQqQQdc9p88QAVZdn/+
WPNmPMQgrAFOx2BKSHCijbkgyLRUMcEzAlU0Um8naKv1I7q/zf4luR6uni9wchp5
VQlQ2/W5MbtlNuZOzAE8cTY3g6Pp2fVnVqDmka7rPWU3ybS1Tu7bhnWD3hKYTVSU
GgKw5pfSwUPIoG5U5idvumHW9WJRMHlcS9PpKBpENeYTxXb9IUH6cEf8/mgj2Ws3
c0SPdGxZX89diTNQTymYBrkk71+yQ00Rs43Oq8YzB3+QfmsR4SP4EwgyT/mWAwoK
ojnarWTjfSVOUl1jDxJcy5CudYuf+i3Uy10zGMvFcFo0aIMAOUc9fG5fbecS/TDp
edUuvG3AllNWh8v21Wg2MCSErNBiNao1u+F4VO5S6mI5r5e6jijxpu83AQAWkNzm
DcX4rCyVdYejO0+fKHWc6b9lYwXjP2H3nxv2j72MjLzeLZBEEYw7b+hW5tRwYkU4
Dx4k1LvW9CiGuRctcDI1iyaED89SYAxbCwxwV7X0nwA4tXqcmV9MP6qqr2NXwd5g
juFZ0ETdwc2Rkp5ISWGpQfTRfWF0snhpZXOrBk+3hWAa+bTDW9bIs8U1q9sF2Pmv
w0lvB1ZVl2oPEa8W2wdpL644hRihMF6Pj+85xAl1UG0B6uvKb/GgBshQyXINltV9
Fg0f8hBvxVXJRoWT3YAovUB+DNCPsH8PP9W9FDtreObkVndmhNyy3xByy/fcqkXf
sZWc1iqT9Wr1R2pho8pS8t/mUouyDGnYJGVBFAohsBa1VqHTID/rQB82TAG36VVC
zvEvNL0/p3RH+48nzXJ6fakCzfRLNZvedMYMA9sW3u+BD1bIc0/vmtMaTiHX8Q+A
Qs+w7qi69wv9R/pm8nb56mN2+JXjfMBizyIpSd4N7s68m9dLTITlLdftvCl6dtQl
bcYAR2BEa7gD5oMu4WbjlX6XBLnDY77sZZHv28aB7y12iwX7hLEjGPP0goFcig3b
XATGFXvFtVvlwx4woTcmhemkYqPlw7TY/dPGkAzesic/Bc/OVRssAqYa/rUkXcHi
Jg2kEN8XzuzAwmJwhaQjbk2akRQNDEpHhR6X4IoA9dKY2N0yGZUgCxU3/yGl6LQt
WPRLbebCfIpGvXdVunL7Agb+qClWkodAN8dtVrxAf3dsYxRWTy6zC8urfWPy/iEF
wo9kItjZs6Mt6KWP1Eq0YdmCyfV0Yvv7RdTTBZvLo+pnrhQOjo1imAbP9X2xHuQT
Pb+CXMGnn+/quA03uZTLU3WBSxQq+SXERafsn9y5Jrvz0V2yyaz/HoIivqvf7wxP
ztSX3xW1A7RFXbwmvZz9E1YeZPnQOR3taDa4uf6tlpm1KoohhGEtZ1uhrz6q2AP9
8z3JV5qMmDC4mKAKbZnCwHk4MpZWqSxExz8pqrHJcIj9f49Y40DILok2T1SspT/G
dTtD5e6jRGr4Mjx9puGOzdl1PViCV28gT0GAbvpQPzadVlNxnOE4OJFoUcKjVqNB
HX94rDesLNHfPzip6jBmYuYQO7yZdMKg92570nCq5n15T6i9Im5iI41PmwGImbWl
YMponeNWrLSSxUgHFR+KNb5LgVAnEjpd6UDYc/wZvQ0r6RZBVqVw0cqZuViNyjrQ
S7H5tmxRxofJWhtsb/zVsBADAEoeDsdG8evuzgbnZvgJNhTGWdQy6yXOnme0PgQE
vWq3h6UdTX8lnvWKYs219JYjF3ZvnaGJFU5+Ku7ZktHoGj8UG/IcYE2n83C+yOd5
oGcGsRD5b7E9qyibhqHTJEqmUMudC9ylKmvAAt3rE8XiNeC6FIh/X1yB/qVpwZfh
u+gImDm5UCpMf+F157MsS0QItekWjDXjWvcKBpYMRyKWgI9cIX3vlvwKz7w8ox1k
g+c9csqKHenZrqbnBWOCZEcisVKl+vuNEhQbqufibOzc/srm/4sxaARZXwVoXX2j
AQ7xCcRrTVbz6GxIiKthDW5ejmCaF9nWJEEhx5U50C852Qgl2x8F/uwLKxOU60x4
qxVeLWtn2Eh8/9ialy9YcER5qvE/n1nvTO0cSh4jgZysUYvJqn7K/PpxxDWoEtU5
fDUO4Koeb7Gf7ouSUyL9/xdUaNA/amlAo6V7ItHvl1mHePoPGTnCCsplN+unfcJc
7GleE0zJOnCG7Rc3OlJRoGC2oyqCFqjhlwZy0v8n8UWRiMQLkdNLzJ2JWCJWNJfg
4oIFM1t/+jfmNnxXrqycHG1kYpC2H+WScozl+jKlCNXtEUFRErvxUFQAYgJE5yFa
HXlUi1zQVlWq8Yb1JJEd2meyuJNt+VgTvw2LtwjRVsi5cNJK2Sg4vX/DjCVWsPj4
ZhMx4HfQb+Iu7xTBzlhrI77eJGg0d4xvPl5K9NQyAlt/PuxaynnNIpStftGT97p+
cR2Li4FnFHiTRzstNmkJj0CexOOrNK9z/jv75USPsPmB3iuwFQWOm31lV0Ic+L6q
1orkwBmIu+/FLbpPqu4VeAHncSG/qYI94kpzp5KWG2hAulgSJjpyGIo0LDJcvClI
iDIj60LGznFaqv1d7ZaH5wtGTolLuZ3k52XynDlVlep9GAwhKJ/DfW5Tg/VOcUMc
Vot+jHxAhlf+w3RRMeNnIEaSTrWBdVdwl6SWJQDqJk+PhEtadcJOovHPi6bjGxXB
7kBcjv9PgHCFsXHfVbHxkylJc7hedrFQV+q9l64iiLRBCoIFWPJEJZODtbT882yk
NLyXbScVat0jAJLJ9fuhmkGW4D/5ktKs2M02rL5Y4pRKpco6a1UK6X5wUhqjxtZJ
70//6rTIdxo3OM9QSDKpBoHYiegAih9sFQw7Ec7JJlWxdNQPIRcii3b0J3Tw5Cx7
HE8LVt4Db3VEzcu0Em3CcoB5ZAOMW+jgElcXUMFoyBIU/3+KKW08AwY60ZinzuDT
wL+qaaQRNsRsmmsyE2Sl1QlLhraGJDpY2F3zuwVdggQCYmsJ+c9zV/DQvhiZG97d
+059HRQGg4k45SbZBGXCDnHccpnJ4N3zFh35tGvw4EtgHqo48zfwub4AAvZJP3DI
VMeIEjPeDqbKlx9/rOAqWuf3sWE1xRZE09y4heJjPxmjrGKp9bRc1BI5a7fxx93K
Avj1PsmWke6ZQu+eJGptltpTBsAWLndE+qexshvQQfQQADB/m9jL5FOCJfPIqAUG
80n14PwfXwgFgzi8HsuDDOALNKq+fgTJhlqAORURVbEFjoQatHO2cybW1vqIiS6G
RZWDBmiP9RNC4lDQlh5TiaIBteti84yJLqD1QzgvpJekOP9VtEnlN3sEeL7a9Tm0
jmSVXQwdb2peWzoA5JUQtY6Ns7QI686ybWHoEKX6VV4+z07kjqAll8mgRn4F4jGs
1K5xsyWb3PT7uLPS7jdWgxqf1qGDS2oFTSXXYxmPz/cKruEHFbCuLMuYGDgwOIz6
8fcJ7PxXdWd9NreDx1xE/RUqVFfpC1hnwz+qanF5paBgI7UdNHvVrDk27rQtRxBK
aSsTL9ZbgBLqZJeCwVDduZnm1UGSp3bbPetYeMna451vkLkGPSqDVnonL+Cpj9do
ctW7NtdVHqe/k0r4JvwnBwe0wMlhWAgWAviduQN9q2Nq5f5bGQbbNMOJHuocwtlE
i8LZnllZO60GrVClKXlBE3oaKKahznVYPyfZqfCzEramI8Mus4jirDes3GqUForN
nF6f56GHIQOcXCOeenKouRULplQpDJ+IFyLL9YeUh2nnDOz9pTMyUCe21QY7I4Dg
cgO0gOKP6OcQJCrh61SLIwtdq1vjn9xngUcvujwGv42pn8n1bei4TOaP3Pf/u+W0
cDkuTxUwqNiWUUF2b/ebyaV7i8S85mpeCKTJn0ZGhHQFoJo6+RbKiEK/rK8wRlMu
JnvlHvImndTg3axDYIvs+dD3ACLFMjQaDcgqOfKIyh0canYXJOZpdhC1cA0Lp/Vp
T3VNcmL6Vk5fLCxonDTcgQNTXZuH1mOPMSOIKlStvOhyqsgtSN+OTg2EPMAj2+Pp
qscXTNQkj1zjNEwofxHCrSMablVyNty0eMQf1c8N/JncqpRIieVWVZkQN6adl4gM
0iouyJb4ohfkcl65OewcH1b4I9VxeTXX3x2Mzh2Bz5Kivx2YOQJ52qu/bSYLCNbG
X+RyRY+tSLpH2b/TU/qhRAw4mh4LUDCXvcIyLmF2qtr+wgIeSlONBjDyIs+ka3O7
gAx4f7nl9BVJ9IsEf1EJTBCNyUQFZOFNFBSlVI/ZPDxpnJHjWyjoGnnQrV7AJlvp
i/0So8T1NMkPGPASqMsp9oLIYAO7A1Jc+jZwz2fv1QVyznwrOz7KdKNBBNhig+fU
XoijHEYI6IfPVU+B5UXyhI0iArRdpzWuzBy/lJYG/xXQdMZDSyhc97I6XjO/95rD
o6aRH8V7/M1Ty47aFgc83URvzxk22z51r33pd+qRBAfiIBBWzpR1o1QRNhCuGLNo
OigSegzDqK5bHtTME1OVxCvss4EJEjzOViM7xNvJjt0LVQZxxGJ3C5369zFKGuk5
IWKS8OgdKSzmTJDcBLhupQFTBZ85xhvFMvV3XWhM+8oGDGQ5B/rvqsEU4UKgcMSu
Hb5wOAEPtxolYbk/5BTr0H3aFzttrCX1pbekmeD+90FpE7Dbx5rK1FfQyUOTdxJA
hbqHhIVjbqkr2B8Ae/e2OBWOeHnH1Xft94hJ60cNDkwFBEl3KlyktzVwZavQm8Ap
tbGr7fTucG6+qdZx6Q7Otptm9Nmm815cgXFPMDVpjl3fcAB9TTJJSt/pBnrkYJmm
BMR2dDHprMjKI8J6rciCy7lUoMVx8HJEwD8RdKbEVWd+s/0Hbo5n60siHitSdtWr
Mfx6nP0a2ygU/+1jWJyjct++GBa4RzcZOOVCe9q723mkNrNJoKPwFtKw9iovPXKb
GRHJy6L0zcsj0/2aFVFtr2Avvxc9miLS2vGzSSdEETEVW7sYVSQKmXof9+vUEFJy
QHE+vhkPuv7PbPWks5t7DA6QQLfdtqhZ4xwgH6AbWFQONAcLJhGIC0mXWQ7l1bxY
9MQ1WJLxOBW6ZmaKh2Zt07Q6C+seZpmxt88EAMuLOo+qaIY47Fb7IyIx0rYt64Ud
e8H8VlK6CHma+oRHJsZ8kMP3Ou7d8PbYwkpFia/qsZMBAyHTQaaleDY8NO+uNuiw
mTP4+wFqQM/udU4Iz5NHEEVwTt3bW/Gu7yBEExcaKXJ8u9QgbtbCDoZoy1Ew9yCM
lgb/CokAk7egSOJ6Gcz+IsXlCuR3jQiz4wXzM+8A7Zo3LbwDQmETwlj+f+aHAAHt
Qx1RADcpmUMj3i6OSiqDeM7YH7ob7WBUkX6GOjdOI99tHl3bfR5rlihHHoK7zoNC
kHw47upXkGBObAnwbkiqU1iJNjwznUPRXq4PUoVpyzFAESNIFWEwgufbGyI+JKem
o5Cr8AQ6n32vDClwNDiDrK6r3dnwYx7mJfc1RHewuc2SndZImyQEqRlXWYmE8k8o
eQIkX3Zjm1E1P1NGcoHwgaelnSrE5hwXvl+H8lLs2o3xrtycER/ShEJfKKwule/j
dgBDSPmdmwzyYsSe6haZigCZVhf2Hk1QfV0rguv7RrxBdW+E/yTaj3JnkGnHWPri
MJo78RvGCghsQZaZ7PKU1WOB13DRm827OJyJi5cufgUatOTypWnFYEJI94HJm+wx
GrQoNBJZpuwn/+/8ndj6wKADK6G1I/2RxxG4qncKvcBIDL+g6/PsKd6dJ5gbRxAu
Pbg5fSHSFysbisb4vM0rYOaOIWvVrRGvQrXgxJ809DDtK/kAVmzaZpiN6YZWSpWU
0sWrwereZQp/4glL1JzCbLXN8CMspsiuDFSGdnwqLl2Gfe98Uz2cV0CdaMiwSxh5
vZNCSaeo7nk/asx1iYvLCwpvGdnFu5rOnx5G+SQEUUHLyBA+ygE+5T4PEPzP3x0F
oswf/EvcSVjloUHNkkLPhLiuxcRvoZMgyiulR8iSA94dmPlaFoG9EGkIHgeGvZtj
72WVfiyk/t40E1+TShnzzR1Yl+jye1QaY3UTdh1XcBS4vguTTkDMvOT4MV7V9SoI
JK7/3oTSr/e9MCv4O3gV8KHSUY6vvLuVu88wJe6uNSS7OA2P9cHH1CglxtcIGpW6
0DTUmxtDHD7DoVS98FJs9K9wnII0DCukSgnHBK6RKkOj4M80QydR1RLwE9+bxjqq
yIqvHKAAN4GfTuRzISyAuLvVolGCTlgYFFhEZbbjL9KZJd/IcueRBHHmOqClkEo2
L2RU7SFayntrSAAeliP5rCPvDZpkDx2XrSVvDB6LeCYCxEE7WiAxUdn3HXnnu5Av
AbHgmGgzGcko43Y82YooWDjCIkOekvk9xfyRIimGy+TGlZQmCqMGtkpM3gYu1Vxz
nVenq8dSijSr5cLiJCpoqc1yQ2UPEtHeXPHafgSz3gYEfJJXSFhqOA9ekT9h7y0b
ZgEWJYu8P5V1yi2REl0MPx3ERuzoCwi4xlIWwqa73Ld9RzqdU6zMwjBc5U59xVdG
uJd18ltWCb7LYTnQyhukrkhnqp0yEfe9fKRcDPxFL29yMOtscp66jjN3mIKduBk6
XQYsa5ufBW+yn9IT7lZe6XSl8fvfwchkAWEmbK/tafNZSB/wVGO5QKWud2GWLESX
GzsvRpTZPiAodAN0anvMi4X49UWqKohasi6HkCmZDts948OR2dlgrV+jwrDOjtNt
ukYw9Of+zlPtVr/f6MtBFxLGHNMvurx3kDVXshDBAETdPOi7PPqNgu1OQmtdxvXl
F2mlY4CwKnSJxfgouWPGQEPaP10P3urEV69bG/Su0+ndgDdsbBNYPJob0d5ZpksE
Ks9jxiuXegbCOTO7jnU4/W7r5JZUUkSg5IUTyuNhH9pJxugo9Fj3QWT5z0Zzw6VY
9lXAuebBLsTqvg4QckcVmcaYjQqI9s/3BZqmzK/cyc2fNfEqayVtsyI3emux1OP+
AeXsmdSyH/p61nyzxSyDHtoEAxbInEVhLmqK/EoA//05Lr9tTV0+cVbGKHl06bWT
UG79I6+7L1AYAnsTyQ7Q9qnwNlmRse+H6KiXO6/1waqt8MQAkNFI6Q1kTbXc+rUG
jreh6IofTcvqXIE8eqAgb6Or53bHop/GBy98hcykzNfDZ2OhoXD7HTew7fJmq+Sn
4cUq7Qz7lV1DrP+yNtvVqoo9A6+jY5Or7H3k4S9nf4QfYJVcP9K/eN6tGNWLIyXh
iZk/RobCnFlVg5nErDFzg6rPcI9pArrmw6RYeVsK9IcGllZ3bwmM2eyGvMhXI6O3
j6qDsoxGEu2agSMzKRAYD8r57sV7u6kF8Mke/HVCRrEMe4t5U4TB8HSWfHIJTVEl
SuN0ir8Z4nAUnX7bS29P+RadyYv6z5ije5wDPBKbVLeQsamdS/09tiUC93VFYgkU
M9UkKvXOMAX2tbtfb42PYLRu59r4SoEZ+AXbg70Cx+EzK+Fn+xRCalaFM80UKmLA
+8vfv2zKswMkDwMsTsB8FQ7eR8fdEWxlGR+h42/neuS6dxLpi8p9IMZk/CV8PUEX
IdOCxTZ8GKEKkHhD7HcH13Ga7i2wBXf/CyLrrgD6Rg4v1ZUQ2RdXEA/GNoFpl04H
REGutG060ERSjlELojX8W7wNGHL+QhMpDcB0kQ+lyE0n5FiBA9IqXjX9CmQWjhox
sNhYRApQNhFwwZmspLfxMtrSgm+gmXhPnLU8WN6tgGJTq1GEyukYlJiiTTSz9pGh
I3Gyo//cHT1c5vtaNConLNFkJybiylgP3aZRtjF+ul1AdlNA9dkHPVOEsCBf8/NM
E487YxL8ftmxZr6SxFrd4kRTWaVmYqfMlk3weI3sdy6mW2lyU88hZ5PcpNjzfx4H
dSTy3/IilteTGhxoq/OWy5gg8Pp4qvgmDMg6NzGwrsVUB47FY7JZN49HzRTGNMZl
sj8quVZyYPwXZGfFN/lPnPXM2fbrKnKmBXn9DYd1fUJGhNLRY4/tYuK0r6F4R6Dn
hHQ4y33g1163JMIdlo9nJPfbX1RybaeDoZ4gosl4MnC168QljqIPO7zMuSWYHsov
KiEo6yINxBJhp1djDuKgkF5PVeVyflW88/YcKt6W3ahCISFlJX4SU32ux2dS1Whs
OFl2g35vN6SfNKG2Cg/Cb813lKco0S52rsSxBJHEeQKrFhKfSUofm555rnvPzqVa
iLsuDUm+2Sgcpukrda8tIwLV5vdSDYZQGlchY5f/L6EkPuDARtX2OzFvKaUqzNYS
NKuivvO3jfK9oOFrOC3wYyQGDnfIsVt6C3LPttTvchmRqkEPzLXAHBVv1IepEuYT
vKXsGt373jS+vEwb0ZQd/V3VKh5kzqPcyeWieNDtOpobLtGG5RYwpJM15aP6BehX
XrHTylbitB+34xyekAwXI9AcosusL/DpozxuPNW/E06s6kfdnZuolVpC3O89j7py
pmx4i9ZJJyTjbOQwOEJAkPByGccLqArfdYii4WEGd0aDExtwctv/kI2wFkttztp7
8mO0FSTZ0F2X/GRDtbcBUQSt/zY5lS35zzDf2yzahimk7AGF0s3EzUS/cn7W6cNw
SQJ7P5ZnRjl8JYe9w7UqvauCzH281VZP6TORrfgs7syauAFVCnuuRkrX8kEz8hyN
v2ZYZgLjNViZtjDKqomCIycsYgDr2JBfwCWl7IkzUctxMIQtY/+EN4gQAkCUUhbe
5hRUo0oed5ecgTqt5EAtM8hLX5b/xxJeD1govyXWapTyJeMS4WUIR3z9oYPzFWpl
phuKzeEUMNj7nxp/8owRHhvh757yhD3H9STNK31XoHnXo+iV67W1gCGyKa+lO0eN
ovQyRBwqMOHeHNAb+0gmOy8FBOVGW8kUe7Ohwwui76A9BhRlX8JvpobxlGA9Wp67
JoljOt+ZkfNkdeZHhyCQsilg8xak/5w8llIOXbQZKhyxS7CS+T2OXFHjpBfD3GPd
ozkx70HHUTsHk0/lzYmxLSbM1Ph4y2BqFnySYHvOp1CJHgeKm63/ng1tj1u8bKRg
PA7LLwwvI9Swt1xR9mAGRHBKC/hSCX3lPKVB0v1lk64OWDCio6i8XQcySUlrbtHg
Z0OGzpnZujKPQAlWDHv9oTqitUapTknjLmKLSK8zo2OWgri4+p74wFtE3hWlRT0m
rcIEq8EYp9JONZeJj49JbwyaLirSM+KTQerRPrLVNvZ2CQSFoAnlyi8O4B2Ji2yK
lsvDRh3nK/aknUrp/3ufL3C6pekt3ZLmBv7SG3Rb+i+OmXLkceWKzusEfZ6650tj
Aq875Wrsy2SVNBD5rEZ7RUZ4rhYTVyRvt78GwDKUYCRM5dBO7gU5y5yekHeSmJKJ
kFFVziDfd8CJdVCdtVbQ1iEQz17+bylLeydxLKKX3wkPhIFEYOG+pXMl+9Vcw7M6
dYKqvgVH0MMNmmtRYFenp6UF1tel1ZUBKS29HKIpL2cqPny2GWHUchwFm7zwV5Ni
NIWWtVZsGlpu7fFNgKdXNYluq5oKkexrqK7R4aIPLYVWnfWrjmnb/eJwhv24RCPR
UZ2ULXx9JJ3pbAU3p6Nqw/xz4uJXwxBSXRTcKD5XroYsmfKQeVZdRLNPfU69GIqQ
2x269qd9OwefDDILjyKVrfiApkEZ82+GaTXPdaLE5U7DafG0rgeskKbne/+VV14L
tuE5en8QJsu9H0Enik2/UyZPwBKixfaQe9LmThAbPhoT+IcagXfGKzo7rck0orHe
aXeSvaBnQDpUjBcLgah4kOmnfUDKtJ3WsIhZy3liurcWFed5VVSWD0iMV6IymBJi
aQXCrRTUXn7HRNpj02fmnEKChbem31N040KpqomWT+S6lmou1nwqsL3uUIJ/GYT/
yC2BQB+ytJyXXfXqTo5vljhhrHMOJ7hi6rdH0G5IwwoujshNGNJFy3uqHEPYql2a
HOwYNZM0EW60MitUHjgFJHD91gf+1QmMr913FEK0jYUiXHbvOmwp6MQXg+M/ArLY
keiqLkM3QwN1TsCu5yRTrAGk6GHoD69DJMAxBp+pH7cdCjXIC2dsiOWWAlIs2Xtj
zprro5WqEsxrjWO+mBYmF5l7PAQBMyw0lw8D5KFD1dC5jM2LaCgcajZ8OewIg8GM
tVKjkIc6AACq6piHt6ATgvwx4bAbWNurpTv51TYeSGGq1kCXsIWds/YROgtSZJKr
Jaz7JZ7kXW2ka9bBOFdRUkMzqIhyXwx8uW4AwIQS5FoWT4VEr/OrSZRwmhg2tZW1
foMFMFnT4kRgooH/CMoOr2eYCXbFVE9QjwsSNIvFEI6ZbRA3MP2Vfq8mJcGR4oWM
Fl9zXBhzGfzWvFlbAfQlA/0c6xrMbdI/MINtrl0pmnE2dSaD2LDsZLIIEoy3zLHi
LTNXQjvN5uOXgDjApVbqQU5k9jG/0j1LHqXQDvDl9vEuq5+EBUg7GcInqLIAZYWl
qe1NSk+7z8mISQYvOcYquPULoXPiy+WDm65rR4bOV/YFDEqNAiPMNVhFs/eIwCHh
/CWOV6cas+QlhwPkvB5u9y7/f+m18RVapAowUqZOAgqUUpsqVGEspdtTkj6ActNZ
7nAO0qjgaGl2Tf2tXuuokApM8DBaIeK7gfk8KSHFI2Nvqi/fgD7WEe8zdb56Zaqf
V6ChIDxVFuEhNTWAlDanqhxVSjUyejfoPnIU5/jOMbBAD3ByF375r/MZE/0fRRjm
2h1fnVXdbipok1zkMrQEQ4N8daZZ4HjUXS1XFBfYLOdTb2my/SsyugmbxcO+Ot3Z
SOJ5UxPYbvr5zfl5j5fgyc1b6j7H+Mi+D471+pMsHy/vqHFiFE+adzqixIASSAI9
+f05CR0Ar2JxNO+B7hrOUotmHSlIGz6pllSyvXRE2v8c/S5t8qA0ymk8uKG37+A5
xtZ4R8KFJOeOAqN/eQPhY0tpgWLMrPXbRFaeXoA4ScTz9Nfjaapjl60s51ueaCwx
OoA2fYPaiY+YP5OC2r+W1/kqs3I70p0/g8v/5VMQR0yLYD8cjD/dp9aK9bq4uNoP
qkTt4RvYAq1E1wcb6XHTxFM2btrQxvT6F5LjYtvDvUIpH0W1cjPiHRecXRVyUPQy
2jtP2WyvydqZE6ab/xhZoKWbDWLHM16tIEIhckpIKHc5Oq2tJZxiAYsNA/FCk4MQ
xSqQIhIj0NQS6B9RZq5yf8nYTtezv9WYV/PD8FZYiu4Af914wBvOhZQB7aHM7uXY
JUgfHHKWDd27iV7XEl7PbErE/Qe/ADK7jkNEpyU4njgxUdx8EWg7wUMfRTlatWjT
hwkF60UCXRmsLByr+QT6ypLlyv0Jt/V1lkj4LBh9xbY5idwAoby6zHjsUJW/w3Ab
azpgXkRi67imUuoz4xnyGMvRstb2cDQpIUwMENrDv9n52O3GcHDyyB+JP1X2Ko8P
DcbLh5+yys4uQy7+Ebg0gXypbFWai17hf7GC/nE+wguwGqPAfqD2P1EGvOh6xyTL
mcwyT3R09iepuRaIlktd38EdSzGPGxlRF3+iUGzXiBsUSgAy92Q3CnzmR6rIlz6g
ElF5684a6kCbBCEuDt+VTnb7bVwd4PoKp7Edzxnb8n/tCgvmmXZCkPrxHwRZjRMS
HE7E/QtlbgGgV+Dosgi0AuAvN5EyG3matjpPttFisGNzc+t0tISgT+b/WWse4A0B
ROyKmmFtbl9BTT1vS5AdFuY8o6Pa6MR2Bjj7wPQ62mwBYS7g2q/nOWIG32brxTvh
hLQv3VdySrSnuu72sEtHGelKw5oLVVPiI0GPeoc1YTcoMIFWj1DspcPBIdgpJAF8
24s/3/HQk09t1jm7dchXKsgd1vEE3XgmMdMZWlpLS4n8oFxrZS7evAkEQvzRTjos
QqXSlyQnIh3v/PQKU1qfkYsmaJkS0iiwRZ7b5G4rJHmHUPGgultHzdQkkDImSi25
Ta5Kef2LXApVc7+m5SUKnZv/G7UqYz9de3+TKiXx3Yn+IgAPuabXeqwArb/vDa79
5SF38Yk1sbDxp3hxM6O1oEI0FFvbmhp5Om7WK5DPO3XA24+rDu/KVU8650pS3KDZ
HBRZ7E/UKBiysEXgWHFgEzOvheJEr2oaD2gjVj8CnpLO3B5F036nMCxGaNZ7nYRS
W/200u5Sm/YEaDvQG5RYpHoAMpo3aG9FVgy/z0NL+nThh+FT//d8XQ9fV61Tneei
A9c7EwqSPksjpCmS7bCrc6PsPQCuTdwgOyPN3J5GH/9GH63oMpkg0L8mZ30wpe/3
q9tyKdlThb4BMn4K3kvFCWA1I3fh8b1oQ6LnATyZsUsI40Mhe2H5hfx+WH1m+Gfm
Zsw8y8p9aKc+QPNAPr+kbjZPuypTyjLToCHyomWwvTw2P+CTcmrDEHjCoa0kLIwf
DBxxXEETKxalBNCVF3I5EdrKPK9STYqwq9o9BCcRxvc+sfk1lD5Mm9HkHQ9tvA3U
VoE4oy6MYwLHMzC8/GhxgaBrAirYxdKbR1ocOQfFXb4vQQ8M0y1G63yhJiZ4D2R/
NH+WP4NPJtDqzoPNBdil6zfrxGHDpgVqEHc4vjcjiK6OhxMXryD2Ylcqd50IVSY+
r95dKrhjdVvALzE2FYnEjE6GQg06fbTuGT1BtEX/EE9CW7aSIgdqmdQlxyDL02GO
n0c5ifTC1EnfBenrFYStjL3MAllntGMd8uPBcEXz1TTzhdx7OfMBzb2CYPIPaqXZ
t3qBRBlAXRPxp4qNzs7VOQky/F+qjern1GnyRJPsaq2nWFqNGdKHw1IcbjvV7FBD
rnDJxpiZbHfb7ngK3+vthlcL/9+Fd2HQR03NuTxhLlcSd/CeXqpkcVysLZswcvHw
zorhQ+OAFiWOs9UvMeSKxGxLGMOqElIVk68B1brQM6X/d7XCtxfSEIKey2PwqFLt
pXEw+pSb6Sd8dffxyEw4IveLPpTxg22AnzOR0dkzjuVOuhC6rrtc/i/ZpChbiO6A
mpDWt38suZtEL3n9+xjl76VXFwJyLVKTRDCQQ1rnfrQEaVmwKXGOIZpoqP6IyCIm
FQzLBSjCRuo/LSfr81qgbnv1Eyrzlhx8AqVGL8joOOhk30japle9VhteFi/UNJUv
N/ur4hj7lvMOpfaC7qZwUcLz0uayy18GzHO7cX+qMbKpyXIaLuQ6qXXw84qTZ53z
R8i9AR2JTDS/OMrKLnpaXdciSSXH/8ZU4/sZpgRab5l6QXc3sH10L81zlWoOAEaq
VGy7YsGmk2DvbXu2JO/rZP/iSPm0tJ/2l9m0crT66V/gVZ/lryweUZibEUnUfgPb
/J5k8jt9jBIX0zmp2Uv3K75bFq4H/nWdCyZLyKRslOgoW9DnEJP2gcN7o0rpGPfW
2lJ4TtGwjRO2gwP2oML28T95oudimClalZRP5m+9Q/aikVW6/0fnufYryhUbo+Pr
cd1OCsM03/kt5/GItfd3FwavXcVXAbnX13Ofj5Cetrd1yUxTUmmaV4C6qryRbO+r
ozPnk8f16bWIUp0XSxSOD3pBSTx/+F+gqCpA7itnjSIeR2q+qxtmMZ7MHD93Wg+H
hoXYMWGP9uzEUGUCkyp09ys/WsCB5pEOurt1Wu3VkG4F7RDmLci/Xf/2nu3xyrbT
/bERNrjAcjd6BjqbDm/i6d8DgVsdCFrRQkDBNi4TGpiSi6wYi8/UIzRrDDtlZ5Uf
nyQ2kTfKdiIdAXgEZKy4Qt9k+soyXRgIZpJLi0zgbPp0hedTLlbcnOJDwh7gR337
qH3cOGD+mzLFuB4hZT8azgJG0aw+owzC2P4KNQpBKjqfDGkLLbKYarVegjYGf9Uq
Alm/hnXmd+OnPiXhUm4b2VT36Vttu6LxsN+IbzOcyHAqJ/ur2/4IO5NOJTSFJbS+
yeJSSkEbGhL+qnz5iS42rK6RbmHkM0mSWmDkRNJvSudpLqOfC9NnepHMLhEzMc+i
6o4PRGsNxuS+Cu++0VLUhkbmbjvO3wp88XjkyiSTyoMD2k8jHCliaFGEh138ImMJ
JxOMSSZ4CS+8+vvAEcwQol80J9KfqcZtF0dPppSIQBbN6dfCwQqtAsMnhWKy1HVK
fqgx6qoAryMOKLUwJ+aysrxEUNuEgKN9A8++Xj3cs8eX88fO9RcGK0JXLwMRHo2W
A7J1vWpeZ+ZmdOALV9RfZNdJB9H194XYhpZap3+dTeWX7pJJhH7SWJz4bXfME2bq
EZYcp8+L7Kks2vRMLWPME1Bvy2HIXWRUBxYbrK8MHYr1MjiM968m61mF1pwyW9MP
x5IwV+HSsIQxTb+QUryfI/cu4BmPotUcdtUpjYqbF10BhGMe32VtbQfO5tAB9wFA
9pwjEpNzefCyvA2RgRCPatqXNV+aTStZOqUbPnS06AsHVl7S613tBABKJ2NAOIpi
N75eflIz4IhT7URsv1M9OMmfxvb/27MbjdH6Yjk4aO0QzdY8AMbI+F4B5Ry5OPFq
1P2Kr7cVxdrem7x9QQ8y8a9m8jiBKuuvIXpkA/yl2P3FJ9lS+BgoQlDnZfcDondG
Q8/Jabl39kgEFaDDDES/AxYYnCulVfymLsCuNlvvuRbvOzPjsECZVLwFrgdC1nBx
IqcBsXYQZ+2SwZ3Xh6v8LJm0+91looswsZ8Z/pryoHIeEZVvr5D9JU+boy/DW8Cl
7s6eF0TU1aoXh5VWCe04MpTNk9ezZUn2ueSLd4Su3PKaFGNVPpZm4u8t4INCC/Mj
PN2YV3OfFYgK8D9Lb7P6IMMIalPSRbvhY+k1P9lcSLrgNc2UELCFB+ycOFb8z8Uy
cqT6tOaWKpdSk1XbMfCNPlGYG1Ka+ntxBWz8xLchHjnwoh5nzWAmVYJDMLS+yQj9
vNTUjRTxSFF2vmZecObjXEaH4WGz6ac9vvRiJrywzVAfvoOydeOYmr8sZlsRs6gf
CJKh5AoDZL1a7cCz82qn53t+iGRfRq3LJLsweN2IveMJp0VVMm/OD9gMGlkuzsDT
R6LO0EadfTwJVcoGzVmrleCmVo6kcHm7MhC7MiN9t7yRQ0nTfG/PN1ifYjFuNfFl
QQfPciJOSlQHvEFjDG1yEKNFPptkEcD2EYYbjK9lMreigp11R8BIcj10XdWwcKq4
0frrC1j8yE2W2iDLNEsPE0HbJSOJijoHoBKfusBv+HWrLTSH7T1iVV17Vaz072eM
nd6Za7bSZPISlTemew8bsAjHdvqvT+fATabucDyTmfFa1LTnuUgqPCzp4lEBst3D
GvmlPx4euUlyQ8ODBzvC8cgfEXIhNik7qwULMPMspFQFZy+gG8IN6Q24EH4BG+lL
Tiofz1hLrK/JKLCGtYESxTYJy2B37ML4nVxQz2U7du7fQW55EigNTcHsnsa4T9Dm
JWW41vRLnTsAkGtB7V3kxI3tAj+NSKb3QJ9otbLeoicCLcUl6Ca0AHmtbIS++70w
KeqXzTA1aXT1cMH3h4Bnyj7qhjaAKIHb4vftNFALWXyo+ELt/ehsoYjoxNKBa1pu
vm5OhGjPbd7hweF3ZM1b+pXHyVS/NGEdKLKxd9ppU3+mDkrZa+PHBAyxJp7Xpz74
QomR3cbxUPO3JbbOFhO2NClYefR9gPtMMlIpe97k6AboqI32ZgCO0xGVXEuUgfjs
hDT/JZU7A1aJ+6ZKXyPCjvAaDm2oqHeNMh/6wVPSKXA=
`protect end_protected