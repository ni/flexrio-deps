`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 29664 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
HdytKcppDjja7VfYQkCqvNrk3thTjd7kgxKC8A4tZ8kizr5r3Q3Cfj0/hAlkIE+E
o1rcKxz9Tw9Becu7n4kAGzl6s8XwGlDG1a6Jzicmlk2Zxl4fC44PJdsuLWfu2qU5
+JJv5lpubL8s7odhz0c7pVCss77Kmvp4//kBlt6H75/O1NrY20PYpdF5ue8JaRZD
fy9qKmS9jJFj0f+vCFX4/hafDBB8uPgk7n5ks7j29LGGezQC2NLYI+g4nYIyKsqM
S7QG23AVP3h1DZTR/k8pOJJCJ1HJyxoaa4TxqqUadtSlT9RdxiTjtl8grbLWlG/u
ye4jDwvuwDFyderGZaee4+sdIh629jkeXEpi9lLKDuFIeqKfCwSgO+wBXXM3JXzL
5wDm4LcvHBTdrKTC/glO9cCGPMrWruhnu1r3HmHzF2Tbd2hYIuuuOeuLr+JBKubr
2krVYnFhS+ABKVTj2OjRt0UxPjOHYzPztFY6LNHDpyo8JQtKytPsueXTetbGeWbJ
3wcbsDzQKEX/k4QYD0RPeeHHsjfX9FPdCniXBrbhy1dNxpDy/R3NWK69R1IJUZQN
WlmGa30xM9QZJQ1TGi+D5S1cXJMlLZ93PIwhkfeQwt5PgOdsvEkFQkniMHQmbvWq
q5ypeejhYxH9Gh81yE1M+8CCfT9Go4dh8N7ii5b+XhjQ+NzyQxtRaFKWds8i+4Xg
VsIxvJi+LyPxCobjz6vFAiIbbkRNWhwVgPMPdIEe0yQCq7XEYimOcXnGrl1NGklO
Z7lCnHMVt7i49HV+YPn/X3cUhEWDy0th3Yhxa8I75Nf8o1yQpYgtMVSy4qIMCTj1
MDDj7I1ukb4amjcs+lzvYrnJ4GxN32HdEY4hablozUvUci4EcBAOm9exQQAkVwIk
AhCoW9U7uushJZaiddkQ9/EL45zb/CvW6/d+uyYS798/fZeCvMwyOtLpgEUGPuSC
cVLdKSMMRvNbfbv99AtME1qw/qRllOO9QIsGB8ajFE+gF9CQvkZKkMdKfUUM5/AY
V5PkvLkPdhvZVZBkDhwvMT3/Y8AncbUbkGMGYvEYNkqf7FebesKne9mPDqy1TtT4
My/5kvvGdBv8aScG8Ztn9IosrYjNlCYcJDASXNoDsWP3s5PHcLYvaNxjvIyLceua
Dm7CUGPAATK+i0QCQ/6VktJW4XlueoI1BTafKEWGsZJZZTDjUSt0PQ0cHcF6L8U9
ChyUg6mKqgRNWNDkANSmxa09qhdYbNvw3G50gq4fR0Vmbk1wZrNbSJi+1wi7g8Zl
L7DnOQNu2DLnTe8YkeGdtBnuHzsNj657LgH15rL8b7It8T6cH8QD8W7iBmQlf6yD
/WOgE3PDdX0iVsB0WvfZNAj8SwHrLUDmVz/R7qdNpLqO3qs5rf+IdZjEsj+o7h+N
069Q0YAyltuID92ftlF6jUsEhgyXT+li7qDrrfdoSQp5MKpDJBCbCMFISsWCBAVB
cu6Es8FVT5Dvmkb3BBKfcFXmP49KCpxgQmA9ZhvKCpEF6Y5ivOq2hAZrjcRJ6mLb
fOcrSasi87NBuLhvkS6U2ElWAQfpwYqXOMm71DcqS6Kh1Em4R6Slqq2fXjzVuzvB
CwZZy2KCybE6/hMfZEQFLOnLX2FW68E3d0dLCZWHuNa8EwIpzJIvxYbEdYgvGU8T
TrsWrLdPqmNgMtMuABjlzVro7g+fkmyEGCSJFB54uEoU3zhLayzYBka+r1cvUO1+
nlUdsipOEumPnVziTWX2iXegnWMjXY6LoDOELHNYAckB1mVtjL4uxAIY0+5PqiTb
Wz/RxrgZqInrZvFPkI6GNmhiJp3fz7/dAwwVDwvOgFKHoi8Yq/+S7i6o1ZmqAiFh
raWfajNO8DiiuMFqCpyCMi7S3jVmL5fchi/tN4emtLWiAkK0mjoCp1gq9LUmFoCK
7cPzRaIqdvfpIFWrAn1rNUJp8bW2DQuT5HPm66hs3WsUeHblntiw+eZAnxzb+8V6
1tgliA5cxmr7SsXrrahhjb0GpRyrdGM3J1fnUyC9taMDbq1cVGROF8gRPOSKO4VW
HBMPMRFDFWPSP0QIWV2R+BBGE73lClRNrBzn5V0WUYqVpgi+0KtrPZvHHqqieSzw
KtC5dDHNuCEGZ/GK8xZlYkQlcMXkbyh/v8yasGGI41mSO1rfqJc+tcOKLEn5aFNv
2wfxCsE5DNxTGFpoLoaUBoTsPoBnfqmYomjpvNfQOYRMO4kH9sSKqSYVd0BjO/Sm
itrfLtJiKrLHutmTfnbCngp1lH4KdTVuFM05SpigDbm3pZelMoy2NAXPdGLnuv1Z
l4HqzSL8AfkIVY13DfSxedQTHs3Wvm2Kt51lRFO8Dc5qY7c4gQOn4OVqUAfy0mB+
kh32WgHJRqeo7M/R+y1FUYuwgpZnAzPT6rxlmKuvYXbSDeUuefAUTXteHgrOExnR
WdFG12MwpqTY+xx9qZGsQEKYp16sn64HjD8OtX29ZwuPAWZgn0widPwM760HdnNm
OzM5jtyeIXpOS3qtnqRpx2LjxGd7YCBSTpxhEnyU0MALRJ2datNF6nhtHUZQad/z
25dam1Mutis7QVXavkSYpELQ8aJp0K68IHrwyEtc1Sj4+sNyoD2tFaiKA5jGGL32
s0MWHQ1Wv/qQK/2glPYZLum6yweAj+6S06hVQs2XLaCRcIJhj1gvWb5ExjvRVfdt
V2MTPSodLAP7p04N1swL8GhfOyUfJhcajwqYnJlDDPqC2pcD2OkfrnkkIVwdwnt5
ahegBFG7ZV4kVa7Sn+OtopH3/05DEQaZIkA9thwguAkAMWyIqEFWVL0MaRau+Xks
ROeYGqgFPeeLUVlo68o1EE2qrKy8cXnslsEDSHCYo1q+8QyDt1mJhgFz7b0o+IEH
zUUeEoeoqepUQpulfw7rdrhtFF0Uu5s7akMm0z6SwW7WVBAhMTf3BDQE/ublUGwP
GsfUy8V/P9q6BaCY2X+ljDEdQJ1jSquMjs/HA9SNBPiRWuxAr8oxbuVK1LwtO7lS
fX5iZzdJ720MpT0PtblkqQOwy4sO1DS2aq+ytGw/IYKhGt35bZarvyl4C4AkwdvL
Fl/eICPXOZrO2kgBPZ6gfpbeo8QEY/eKa6uHYCUGrsXBQ5fYRZrurvC3Io5rrFQG
fz4WY97j//ZSqm12ikNt38xKS3reiftFrEZ4vme4g9ouB8LWc3jOSEzZ5H7mh0v6
TRFyLbZgsnt2DtjJoMYXkBDKcwv4lRpZHyBa5gKiUTvVRQdK3myP+kAfC+iqP/BO
QW5EvLbB3lViPzc4chOUQyKh+8KdH67VUuWH60Q5yxlzhYxoZrLi5NhYcIzIR1oy
8lqNY5MKgaEUg/Gn11ODFl6edbNeoeLmz4dcA9DedymcGgNBMcg0I6ubI73AR4km
GMGYvf2GS0e+N4npBviMzjsUGV0VX8nvanZ0Jq+E08ACTrJbTFYjY9Hwc6DpkPqN
38n5NuHry4nGZ3Y7y24TX8D7c9oCkG9/7kH/Xg0xwuZQNJL6UM9fDakxw8y4rXRx
rKrvi+6PlYN6agyD1x/uRYDdbG6lqCI+9tr1m6Fa8JT6MmoJ8eV+qnNVbcM+uUQ6
1KPLyHQGvPIdupYGT8hSSBzpBPNNCaWmmzcOEnmWKJItTG8Y0tL4CelmCLbWHbjt
N0Idgq1gqRnPAlc1+sXrHbJYAqS3PZ9MjX9Z1ue2y8/BEY0Ioo2YxfOf3C6sFE6/
9nTj4YdkqWbsXg7HgT0iRmEI1ayAPG1sRC6Vm8W+gDyyaLheZ5gkq+eHu5x+0tMn
WuI3VVleuAqqtabngesZ0+fos52G/gX6NhxA/+e1Xfh126++4uftIACwhan00M6J
HgUYjstB5MzHdsXyTlvIEvkvYLSR7eKVAkwnStUFyF2CczXY2RfHCADY8UktypSb
cqGVBpbo5T7NzW91duNHjVxrvKc1h902p8JK4p6yyZeaj7YGD9PK50ESuS/zQ6uv
i1EVGR1Hnnp4tfE0NDq+L6FmL4xmDukSESvHhkKmiJp4xNH8yygmoXH+6oggeONV
HMWsSGYf+N2rl1qQ+kzhHW+VqEsicAc2GAnTfHxDZ+g/ZxF8/3lNO4N5tunSLqGS
jk+NDhWfXSl/7dYOWv3vyzJfQXJeo6/2pyI/6Va1YuoFfQoOVQjjAo9rWekSDARU
CI09Tq/8vVRnmdprw9sBWLpVUVMpdaJJn2VyyVQ8rmM4PzCJCaWbFXPzQxGleQNt
5WTBKlwgAtzcVkXycuzqsWIWc/mUa+0SUVhbSt+Z034bgEXC7Ew+KQidLST7rZEs
McZUzLTw4uXcwoSndSAnwsjDdsBapNwNifapx5vZgMJWHMcV0HVw+fdQ0Molkial
er5k8SjcZRAmPlDBf3CPCwDvxHcnjhx+15Oh10LrgXLs6z1GO8xvBF0VEE7UBQvD
28VmH3zfnX61QaQNS5OciYtuHGsEYDW8iqfr8CA0po8F1aRAV/mzzN/Mnn8J/Z7G
joiYMU4xRoDLzpRJioO0hPwvQde0O+knIOAAOP7xN7PHOUxqm+70j/6QmfHtMNyc
eetN/cJfOz6ZLUp4qaT/tz9Blw13JyG4fnJhep9KeQXoxHhDtb53MavNSTZFV9IB
ohYuwD7Z6vUegGgdbEN0e/Dokbrnsx7EmpKPCmbUjgFN12b3Ljf2niD0jgqwxTm/
sukxeLZu3BlEW+t6iM1G+nmtXp5qy6yDcx5gwD4n2qOm3Jgq+epJcBKEyNMlGrmq
Jj3N6Of1Js0LWts9biTwGfaSiR9W9Kwhi/q4Tc+WVXtCGMF27QzxKmLKSyqxHBtM
20uN6xwlZP1mneJWjD83SAH6ZK58jj+EwrnVqQMtgfyy4EXp+DqmDkaU9RYqdzin
FzWRkQuGogieTBuwl4JEUV6dEBcLXR12M+jRKOGWGB3KrRIkk95vO4CP59P15hkT
mCdlZgZ/hFJw+3XBPQD5USCFJbWNWWRfAv/La7mJMw4ls96WkmrNf8vC/WLlxp9y
D/lXZd7k0qfH4naA1e2aOwkZ9pH2pi8mLC3k+i/x+Dhk0giV/cEXJ7rtNR+dTqvL
3XZp08d7fX4DTSC6zgpTaLmtcUWz3BevVRd8HDrViRxKULBmc2CnDyQtPCxBldTH
N2HsStyFBDUvUlrFZoAF0+8k0Gb+QPhL+ad+D7avKGugeINWE5OpJLi/A8+XDu1B
yxV54taTw59q86qxwodiBZFtpEjBt5QJWogTM7QbZybE8DhBe7f8sRdBMCQNhdAk
Hra7zyfbvRg/YayHuF4zef97qSFCFZgxyCOzZRfNmDDBIXXNk9yenQOnfSRi1LWP
T58LuADZ6qj807M4TZTuZLRuZZpSy1RRH9+xKp0HF2AIDyMoRhpRDMFvD3EXngFO
JX+NjLaZgBgB7UiUXApqQV5a9GnT7Va4F0PAldIZShuDo29LJCX01s1saRpqj1JD
FT6JSE35DnolLDJtqttA3GtPHYRIQxWd43Wv1J/sEm0JGThNuepvVbrh3oyhFd7J
V4fGhUNSUecpodccxCQ05/MmLqldvkmwLvBpme4qI5Rqoo/ZhMdq9zXKxKUB4WMH
jz/7MHzhLBJtfoQLWD7dc5Xb1CIbvLvUE42XKKN536jvLE8l/bNF5ZZov4g1rc1u
Byp4nhwK6CEtA5zt3OQibIiJ5HvPNN7o9cXMcB1BFBF+vYqfQjbBZRS8CMGSHpWq
vzG4WyBVHJgnxgFcv5jByk2Wf3602+Ynmmte6CEZXPNupN2ccirAzxYLMn0ByOZP
a7VzRP+vVYMImax5x9vq0hbXT+TgUH/7w5od2St7LrInIkH3na59k+Qe+tqaw1/6
paumYwFTCSN3NolUhMkLS9d5BKg7FXUtY+hCcvgExsbgfxv8YYkVvaQIF5+f365+
HTVr+n2Cg+QNdfdSdvNAJG9aWweM93WfaftPoELclpf+VPcuoi9pRbQ64vBoflwx
UlQnQdGzpwMcdLaJSEBuExy5eYKer7jPpijn/1+zErzK11MX/b9kMNPGEuQz46a2
kEo87J5RflXBk2Adowk1RQpfRxdjhKaSwdN3y8G4NNCl1ccpOvH0frDwP41LJKWs
jHL7MG4GtOpo2v8Bb/532GzuuqIlVw/1j3Rtc2HVvsP6Pgya7DFcaykfbwcxmu9y
/grGs4DEaCRVCbHk7xVcF5K9LvlcTkfjb4PMy+X52gB9UoRNvu3lipBqOiUFbRtU
v9PAAiFAmPg8892xTgkM/YQiU37ot93igpQoO/0gKNG4RKjVG09mJatOcRAJKIj3
iLwZhS5Yz+0olIh0xy57dYzVHIwN2ohPHTunmmghJTUU726m8blGErzU/A2ePABg
wD4/zApe2jkqVuH7fmGEkj0iXKduQo3kbDd2RLxiFHVAwcm0vusu4v2BliztKc96
/EIwPlBgVk1lDLoXxApAGCMfIStQnhlEXhoA9qKUYHYUXf6epi5fioqMMWMpUYJe
ErEz07v7eL0mS94dn7WCycXWytIGlurYaKkPKeOV1AbsKklnfqDXOZ70WUCVBB7w
hJIheocTXWdDzPUly4vYHJhbbM4DVeDBdH9PYvU57Ku8dd26ONkZbMYF/A3tulHU
tys8Ir1145ZT2NxBN6nI23vD8a0ewG5dpkgAwqwdbmK8vG+GNON9b20ZVmoEaMvg
cuN1sXj35+JfNdvYLLhEuy+K3jn3+F38haMTwf9DgwEpzZ7VFkiYr3VYroxhjyK5
c/8mzW2SV75+bKYKlTFB9NNpuFiIKgGdN9nvduihH2FHAOj9QSQ3E/nVvLbOBQVL
xqQTesIZKhcTTOFPl+4ERvm/5FGFbW7buPtHPfhzZpv0DLB2k7GU4BWNAxMk+c8c
6Gg6oglNYh1c0OUNfVaTLVpYoAZl3TDlqMDRlCHopPMMk53RRRaw+CGLpxqoRWVz
peoveHI6UrCflPXZsV0EvRR0cKkBHX7pw8BPHmbKlqPr+t553nqOs0sR7eANCiDn
h2oMlLyzsH2jknKGFBNDHl3TYQpuLJNMafE4beYERessPQLnIfnqnrUX/cbM1NDD
U0q2SR76RSTUZCxx0+dm07ELpz0Sx0LnwYy4nHGKCuclgA56AlBaCJXwdVzGYRLc
7l8ev8o2A4StiASxUisouPgG5bNcPdPb4qDaW2Kq55TLYxX0AaYQLXS4tgbdNT7a
ez9OPRto45AoZ+8o58tayVO1k8llsNQsStJjKWLuONPSQe40YsmBZ62pqZNeYj1T
oTBxdj2lVGOXwAO+cBJQEctPp/ZK0NfXYWFmZ/DH/cUJj5T03A6nrim1/uQKePBL
JwmP9lc2gtgmViwrxeqEn3rbSzif5+21Ao3PCqh8j1UJSEIxkKgXeEX6QzUnKOGC
8W5zSYlAQEUOF3PtW5eGtzdCZDJHkYtGlv+fkucyfRNghW7UveuivWhdiI/ubghZ
dVAMygjVufX+ZwDy6FVlMoIpJZ1TenA+mB5sbbKY3j0wY9HPKPMryVEyTKoE+ggR
4JUCJmYDI2EAiPuyIyDJQF+Xaz0WbEKfmyzh+8srKanZXng5pxDKlDMdG+H7ct6j
64FkBXxxocEIrGnKIANHcLWDjKnvPN5/mZ2SFZQXJzrcBieeOjAS3nt1Eol3eOTQ
OyJ9+VNIFW2Gb8HhIpKOIPhLa4eemdM25T9z71rfaZWv2eXHS6j/r3dlw6LHVEWy
MeiZGo8LL3S8y4m+Tw4RK170APz4pvgCEYn/gO0HB/GLIgK2GPxQRMgAp2TfYqO6
pYwD+1uQ6IGKm+poisguQPcJ0qB/+j1DYQhRQ8xySL36oq7cr6cJHydqPeWQq8zd
4PWbBXety466ZTr3z0BhBC0M/QlyJYEVU0tWYQAcPFA5giRAJvGfb+JnlpeT7w0y
6hgs1ys6E6kVxLQK0RkxlIgLihqFbO5D3rTBDXImBVdI2V3Y63KYUj+IOJrTmTGv
yDS1t/G9Imj17Mi2VsNbw45BYPyAigZIhuHhWDz8yNV0gEJxbPow5QRhNfRWSigI
iojAXFhGayZeZYRvyDINRu9E9jZivC4t9axuQgeHNLzo6PSIx54xdK7tmJSnBV9R
kg9/+j6YQbHLWr3kByVWX5JL825OYR9x8udIGYl3FQsxmiRNh1kPrBLiRyLAdUGc
drhXjLuD6Qq3I7qrpleYmVI8LK1P5XT5h95WNZhChcTcKCTe2XLSkFXQehUDtWVa
SDXKxymhLNZnjQuGdIbUBxDyu+q5OMOcDDV2aPrFCYeHPoGnIEfm5N0nYeZi/z1E
cWWBW/p2b4oZD28dDbEjqOpuxlVsrk/FBX+DYX8s6L5APJsPC11MjXOgVfJKabZB
2OOWwth9glP9Rlvj7phZgEbbqmGRO+ySkvAgU2GvtzP2DXn5ORCZtZuSgnR6UdTN
45cGxp+ZcKOvEob/IIJDJWETJHSxsrfywuDKqjLjf+01EZp8Vc21jHV6w9T4UByu
iN0+jP5PT39bruCLUSXIv48LB87372IQpvPYfrPqEFZenim9Tm3WhYWD03EWyYhA
py2GwLU6gQAId4YpYDdEBxXPaavh0E2jWTXxMFoV1tadquKhxGM4UuEsq82Sptxz
kNOw/wKDuiF3L6IbMHfvLrF9tRN1HrhZqIYUA4JZ/43lEOVne2u4hc/6vIoCWxA1
Kly5qMsO8K1PeBz6hYKMY67iPdhaV6dwrXmVEeVJIl01QhSLQaHfKbEhd9HSnZVq
7MZKjB2Kwa+N17wQM8Bl/+hUYmQNbRIk5k1rAcn/YGvpW7IP4d6z/ZB9ipL55CnL
jyuARPL01sxT6aKnlUMERceFtlTtaLkeGEM6ey75CQdyBMPLZLKFoHrvaR8NvBoF
MSPIM05Dv/i8FXE9gMnKqmZ0+xlktdwCq3WKxDj6mJOmRnte9dpfGfXCEP/6TCtW
m4sPOE6W4r+CxwnBdxbg8UtRM7ZFTc5GiF83YBYCiRsBbCipDJaaHqxoHaODK6P/
2Q5aVLcoFoAc6l8pepFyv3Wq3A9vDjU9qVIZpuyR3MZQoc/FUg6jpgFAYfBYRQ7g
sfMml7MrpsITSNkKrBo/Xvn2+XdbEZQPCguziMlsP9SNfjCJYkY0Fbk0YN+3Cocf
DoTSaeqnLD1k4AIJTRsjRN7saf1mhT3+Jp4FNDG8QGNqVdg+vzb1R5GEeCFvOynt
O9XibjO7T+jiFne5RnaM7lRmI/Wa9Rc2QUemh5/7wWyd5L8TNLVu2rWRqAtqm+oS
M4aFviXQ8hI4KbGi55fqV/ao7mNXkdat1pWtprGgmOaOf07iz7neK90V7rKppESa
gcACQ7Q2a33h5kEYvCbITfXry5Xa3QNJE4asRYfzCjPU7pHf/VAUkAI7/FfInQGq
eHVGUXOUVv7RD4kTbcqaFhovompFq/4R6DmRFoTiWuxgJAK9Il1c/63UUpHBavBC
KdfBWc0mxpbsgLcT3XX4iR3idejd/T4leRXZf/isohepNlj4AsIMHap53Gb+uLu3
IIQB3qVpGKNlopGYhSHp7IzJm3P7+rgrdEteWKk6Fcf+vtU1fumQOhabwMioGZCg
y79DfjbanojTJgJtU4t0cRhSh3N8ws4CHLSnLdAfJlp475wfDS3D+B0aGTRSUUKM
0917XXonSDR0Np8iu/e5MMKQi9Bjg8hOXl+kf25989VXlsTFLA4bJ6pltf0xDNcs
bhaTZRst3Ox+q3EuXnR/zOmFKhxaQkkt9dZn/myHxVdTiy2JjpVc1G6EtM9LW7bc
FtYuhIxaHBQCQYTCxuuAQJ8VBWs+GOvGJFMqpr4ACnTzrhphZIWGMMobU26WlQa1
OtDzqLMR8zORyBEQSO/JpPTH+80je3oSgRIshE9zIBvXbXGWVlNE/eup1CxQFjyi
hDH7NvC0+at8xzUEol91bWVtNnU5JRy8pn0kjmNhRhfabmsNeFp80rOTX/VlPscm
4QGTmdJ3+ovhs0TxiaSUo6v/4PFVZwPxNXIZAqL9JUm2wxfOqtRsiFV1/LF4PCs7
B8nz82ohO9GnbDBW9TU6Xdt7rKYT58EEFxzDgKdVO1F0YFU5+LUwQ0AKmNmMF+Ow
cMnVV6a/ElICCstbdKZ16kke50GmNlMSH1zmJXIBTNnlL2we7GL/KBlHTJvJjVhZ
pa5zcmpZkSnDjzq6gjILCSxC8RTX/5TEPoKfhB0muwKDGZrcdsakTH8ypG15RG+b
MHNgQe9mogaRm86UgG/g4s5VCzMEIm9yepcVixi/IiMuIDjWo3EVbAeseIeJxnQe
Qk2hu0TlvTUb3NjZBinbG6BDx0edAHaKnghxDT8E6iS3HN8DBU7zuGjhBWd35Tr6
QfOX/7igwUBLbsmCOq/QeqVhYcTNhlgI3ySuEfiX8ZSMI2CI7sADOpg7Egr+ncyd
S5xjUa13TAwenDsZnb2r9ZxA4zdgb1lXlI00Nx5t3lIcRwDj8OZivVuw1FRK1ka7
IPmxx9p9vyt+4TAaj1oWEXL3nS6+OBr6n0LOvPh4U92/PW6P1JEAQ8+zRevRZWF2
Zc523zuODHevEIIuGiXiaMHOcotMPcQxlDCjT9/1AE/CrkK2YiG9p5F+naSwS+AU
BMcnOjNlQVPw2U4m5EM7sH8OzMuK2TrC17YXQxpBKaGY7G8XePywMgUxwvJI3BmC
uA7mtV8vBtkbtwz6Df2tixTKhuwAkwR4WBjfvvf2J1RDbXouvtjUL9e93K2QNwaR
AjM6o5SAgRXTFIWjQH8OiSFsdc3BJSl8V/qBi2vfmPGor9iYsfXia8tCOrI9JoxN
Z2wNFHVojGIOwwbk7KeXN4oKZIj1EHUK9E9DU4VVyFH6sLUvcsGZ4DxOgh0phTpj
Ehjybdm4+++kiPvwMkUw8/MXmIWnzufL8GEYW+yY4wWEzSGLT0Sovvr5Ciznv9LQ
Hf/j7mHlNkgun30RxOvPOA4ePp5TtvYLvuWntoiQ8wZxPQnx7+7HjBYJtGRtFvQG
u02HpxR/ddXmSfyMWqY5O0TWvYKrjVxUP9BTAPBTltUTHy2f5yAQNRLnicpm23Mi
WuWBdiqgAyjHG17AL9mrimp2hvAo/KfpDqaAx+/vx0H5dvupmU3hi4N0ogMF4ytT
HTeiU/R6XCr0wgTIOQnAWcZn07ser7F6ha4qKzWKpjbQYXCL47q82lAXIE/nzqIb
4v9OIGnJjMYVfNydVSPWAMFT3C7Ja66aH5A4j4VneshCviOciqZmT52FlEPWd3dK
uDI2Ymkx9CymDIfJjPaQmNc47ZWmZ//IfX6+0SRpE5PBNNmAvt0CkykjdN4pE3U7
DWWnkmw8TcZypXz6VwRU4m8Ic10IHxSuzOX/GaY5BX1Z+4XXMR2hLDWXrmBjsiwr
8aw1u7w7IIePblyAYpnrExH6isLNxDAWxeU9IZ2VowG4tbCBbMY8qieJ9CadpEKn
35dPcNeel2lHLg9doLz0+s93KSZ4NrZ478prtF5Xl3946OqucQ0mLAXrvKPYrs1y
1U8j/bDB9aFTX7gXUR4YLvZg0ZYMfrR8agu6ve1tyg+301V8kU908SxVPr8yDVYu
JZY1qeGGR02T37PmFYmCGQool79kkGdYY2ygC4v//Sy+nXx4GrkDn0QPS61ooz1J
6cckdeLfMe/e/tqAaoInoC309Hf6ntuxp17Ksav/rbV1dckPlZhfS36DANUhUFKT
nOxt8cawN3QkFLL45wTics6jznJuw9l2f31DhB0gegIzBj9lIGjKQD70ACvuFLbm
ZKd7cwI9icKqLLLoD0yshU5hsPDeB8/I+FzLTgW34aPTfPBSrY1HcqHEcrjSchgh
T6Wni6swTgBI30wDqXlxp2GssAGslYwxZatdE/6bDstP+a05ZJTAHOs5zIsxzD6q
exER0OFuKZXrRBRL8kSBi6/yRwWUuGTgSSi5X0q4UihSh7UCryOC0eeDgDCRaghI
TzxXOceaRO4zua90T3EiNoe1j4GYH6Q+/+7cG43Bj2qSxRtj2ceo57g1HGcFa3MI
IwReEBWHU/XuKZsGECLi/jiIiZl5E3T7YOWdZpgMpkDz/s161QCkkXYNiHFlgAEG
rOX9uaanq2vZML6LQfjNci8aWjsNBa0LvdE0L/ppUMnJhfN+/Be497ZdgTAtTABT
MpUS8SttPB3wYfmp4qAimHXXfSGHHy3YvDWI7WXqeFvDXHJFDoKaGv4WbjMC46eY
SbL/8YNDuE2BoVzyHtsXcBHV3AottfN3mdUA6LxJpD1NsKfoj7Zf4r0sSy6eNnvX
JBSh/0kZ18Qf/tYPSKIMIYczYYdTGY6b6DdDh6nAIeblg1anX/cofWO6CR+fUhw2
dehyrgFf88sE8FY9iejyqpW32T01vkl1KokWTPZ83mqW/A0+nSqMO7z4b2UIayME
FWOCr7U4lThW4hJt0BmlU3myspzGyhF0DR0AQn6kyAXcSsSM187hSpSutX6lBO9L
f6hp9Du0czavto49k0rlF2x66B8qBg+bYohzEicnRiI2oI2iI9XASg6l98ai0nsO
8+YdOXa8m9cll8UqY+F4/liPuCnN5UKSLK+tBnPDMsxCGKiUAqLmwvC2aV+Ylwtl
f0m3/6B/fE4xPMPecpnhh0cfYZwM453CdgX5pEu2h33BApo1alTMuaOjjYQw5otk
vNdRW9x780QspAHIhDxjjpJgg9t4yYBhzYxCqLflJ2KDF8HuyyueHyU61RfyC+PP
pa8a1mcAErzi+YiPJNZPZRznv+DHwfQc8gfs5D7A/NKKI2pWHvFgUy/MfXHe8s/T
CBT5dZ5QORB8XtjWFC24lBEN09GrSvrAOd/Z6My1wUEU3GsMst2naJ37koOzI6+5
h7YaX+GUMOhbAAOp0m1QyFqK3SLPDeQDRcWfoKydk4s/BH6tmcAWWhlzG9JyNdqe
KcAjbvj5fppBML4xyYi4FqUk5bpouiURICYGcKL/A/sSCLtUkwHHufHXP7oG+A+A
fgAftCaaprTfk0ndyVLwNu2vL4IXe01fEoibXB+exU7r3hfdV7V0xcTSR5dbva4v
0fWUCMKhyHq08lg9zDWvkkdhT8roHxIgUN2/Px075SaCyWPQAIEOkSh7NmTy3G9O
d+EKuFvz23cfkak8r9n5s8dOscp+CbKolClD6i+yfWN2FO8CUg2V1ymRj1YkfGSU
PdxcT0rxwNBLFOCixMfzw3JfxvolgFNrVlmP7cvG5UvBOYKnUMu4EY+sBqxETNpH
J7JivLPiPpdzQ+43zEo2RVGhK48YtzEufIGPAqI9Oe0mvdsLKWwangHSvB+Ktp6y
+axbMmJUCQ7x5efB9s+omPw8GR/c2iPFS6TUS7aYBbH8OzGYIT6YvHObLl6Jo36U
mGkvh93/JGIMevAlUX9n7EMzb+dxhSRye+AhxNqbarSp4+Zziazb5HEmupql03hL
MFVqN4snw+/6iqvGrItU5iwOlLrlrZgE8Uwc3qHjhV4ZBbOhF51hJU0WYBwMafzt
e9TgxwPn8c3oU4cG7NzRfMm5Rdd+qjKsbrrWgMWfn8bE+3lHTtXDNZ6EK5eTCQVP
vj1j3RaKsbMDcBlYO/pIZIRegKzE1ZKM7sFdJu2cHBiJdHjDeNi4Q/2rFpVbP/gj
UacX76nq0udTLEe4XWJys58EP1Fwhs0ukF8+5KRwOAbJI/6pooCCdVcoCZBSQOkb
A/tbRdl1rMFcgf65jmOpNRipFY8SYMSiS3baJyN41A484YlvUoOkiSOnE4L/NsX5
CpcyYSplGs5hKPB2YjjGz6SPbaIHIKxe94oNVzmfUVKONBDID6uV6deZMrS6wwce
J6TPtg96aRSscQR08TEf+v5Y3gXFyuaVj0z5COTjvvYiI309kTvtJvCH83ExQbAi
zB8Pcu4cTkwmFuKT0odTTW5ZndpwUTNO6jTaaOKx6kmJUgfVTk0Ur++YljXBZ6fY
mQUogPuSm9CgeUb9JVLED32PhR7S1unDG67JB6u0loZqNSQku2XpgFa8+w1TOpSg
mNuP+FZeI2RzhJ32d0QX5h4N4q9vTNYWReBMHMr0WMOTnTl1PhLoU5Yt8ZLqjaY3
0ejkM/r3b+dUB1629wBAdNTLKmhJbkvB1Ymxa418ZHue4xxWSsDaE02MyAm6VJAd
UYfNxsX+2TfiN7rJ1X48agRtmdpeMNNTpr3l59UJVXYv2cAGZBhT+hXuRXa4V0w0
Va3iizqMZINBzb8bin1aD8qrhnqaZqRi8Hymj7kreqTSDWGefKgzXhVTYwHKyDwk
9a1JVl6H6mIdpHOo/W1T/0d74ozuB3aL9FeQd13f4gEshlW0KhB8QO9KXMUN5L87
iQ1f3k+R4rzgjGf3u+UAA+Mdz2N0NT696PdHkfMnp6Mg4RqCFjTpGgbmtK+deuJi
j0SVB/Tk9CrCLToDk30Ilq9F8D00bGXL+7nFIRO5eQasfTD8rXQwsPCml0RQTYEr
LNio4ppsiLDq+qyZ4HB3JIaIkQ13MdZi7XoYNGxiC9jKsX4JAhepXcS+XV/ClyvK
Luq80LHJEF+Ttuv7NlGYFWlmv6Sr6upy4I4NbjaIpf7EtuIEHKlQ9xpHWL0w+sgV
o3jf9fv3+u8lKpe28HZ37T1xaTtZ7ienz+yjbdnMosPRO1Wsm5VacyJwT7LP67kx
r24Em4EJ4r60UH3sBKnSImFJ4eEXJdO7Jl45vcnC+jxzYgnOx9oY1rZ9T3haL8wD
JTahbq3v6Ov+QFk6XsoDBHlp5uZ1S9r7P98WAhfswUZKPyB2W8EJDgguaG3wnFSz
lLoV0X/KbZD85PsXwgOHmQoOeLkDfu4qbc4zRfcu28KaQ40uH+zAv7ZzUKFFXndG
TH6UyQP24M5vHfVKNhCA2Y34Y54VdklGz7O6jsVbP3qMHCjFhOOV3IX6FT01YZJL
RFgqWBFETO1GL570lw1IC2iHX5OfMFMYu4AUsHv9XLI9wQ53cIgX2aU1wmOMyz7o
Khq2XSt2FNq+8npTjeitkYMS+Otx/iId0PGvjQdiGkpMBY/yCcAko7/l3+uTXvW3
gAAWkRGi2GYvUujNYW7yTrWMUqCJzyZpzyQGI8ysXHaQUdJOxnhP01unBRWGRaeY
8TPrHb0pirZgmNHWr5Sux4hFG6LIUPNfPU+Qu1xV/i/wo76D/vcuWhm9ArJdGw7Q
+NBkqa2MxQ7J8Qa42WwDde9tX0Cqs4f4nlPP93u9JXP4ixWJtkEf0c6ehTxk99pE
9kZbvr18xoCiqm/fYCIPY5MrgIORfnYLiBS3cYyczA1gl6c+1gwjuBTPN7ZUbBZR
35pgUHiOHvOounYPu2KPCnN8j5ECn7R97pq661Y9wzSYKbbJgcbkGRlRKH5voVLe
x3i3MQ7zhQFQA2h9gHsA9Ihy4fZ6+uUfS67G2vdHM2pXJIcYneybo9QaXeqIdZIX
oqPWSTwYdGBOBL9rIgAVZyG2Y0u6x+EthOViDkMm3r4Q+crhhyL9aGVnwCJ7IV/t
CDVtmHqfyWgm09KSrn6Sf2V4ia7ZUiFLPz4py6oc9cEeK38Oq7jS4wOo9a7M/DGG
HAXvoh5WL9Ix8i2+D+Nl5KW02yi9fK/d/K9sS3W9cDsjKhKilSQXly8JSDfdnuSZ
tdC12ZJ5DK33H6xdIyKU6srBQhwPCwGWdtb+fNRF8Ct7ecxrZC/HK75dZguZhyrC
3/0HWrfXDaucvefSS6DRkOQZJvWhHP5ZXSrSzmzhADP0hGZ9tz6oo+dLIdDf5/+A
QoveHzhjhvfcKEkMiZeyEeGN5WVQvSPeYaxk1Kg3SVA8tjX6QL3R1oST4sMJtKjo
Do9Iy3vlivXaHjfX0ocv4b3SIC/q0zoZNTM0K85s+drNcpmC17IwmZXz3SRGWtRo
umRwapRmdjMSSXEICjRvzgnAzgX+2QrBDK0cPhAnS3YMXOyJ+iETzrZLRtH950Rp
xK8LX09ZykXqNVKksMjN7Q+MaPIoHi3O0WJtHP+PUKKBVXjKhtYXIdBl2o0vBW9/
TPJKCm7IPvt16IgwOWwNmWXlMnmzOrEHp2IAa9NjENMxlRyQ7rw2/Aeu9z9czmuH
6cV/G2+1FpCl4lcProaKeyduZFxIgOun6r77qJHvdioOa+yR+nR+K4eg3ATHdO6/
6XYH40SOvQXSZvk5nF9U6DPlOOmwXhCwPirV7VXOUP/ChwtNTn/LXaHM47m+i00S
V/sa7oDYmTTSfLzsSlncrJLspFySsKlKcverXVCfnypvM+O7cBxwJzngRAxvbRYj
XGIBV8PpdUpqW20zls8SjVho/POJ9GGDm5AVGNnT8k1ruM/MqDVNk2ksr9t6j4VW
5CIwbkeawOkG73OqtmZT2mG4bOsGt6ORfaUfnzee1aCTAgLHuf6DR/fI4vZeLEn5
XTwgy43HJM/ksLuNataMz+6KacdY/7vA72U3IcJfHAAnKc2CaEJG2fQ/mDd2g4rL
6mYL3zI8BztEj5HEh8hIvnS9E/xvG5S2e1CDlYNwqOV43+L9RcuKJgY50XNIjKgG
8Mpeb5boS/5HrchclOpdCXYrthEotoJ8uUklJJ6sT6niPh0i7C3PNtftlpJG0a81
6MxvqJqF1AsEgbRCISMut9MpQF8UgHm4j49pSxhSx+cuIU9WJnyY7LhXFTHJCEr9
66KY74j9F32DaKFS94Q5QLe3cR+IqiJZZY9AflhJ4ToKFe57olOF84MM5Q2+16Po
FBetUlegQdiB+fs2+Dm/kNDNeTP9W+cH+OJRie5nNiGngGpbFcfKFOoRhVSZ65Bl
RvEUb/fthxGnABB2x07Z2CAje1xdkVjxcAkyF1dN5xeFWmn5jQLNg5GbjsPLYwW5
NkBYAL0/bV2Kzk51WlJiLuegkjYOJtC3ndWPOnmS/yXwwzOd53wQAUa6PN15r1hL
munAO1I5vmZa2heb+5D0WP56LoLJ3ahxtxq5/44rrbYvGXY/RUOY3ACTA/aVpY7j
WBkjy8QtYm9wccyoIQnO5uu7mPzpehvUrAsOy1atQqz37srCHA8qjG03kgvbZRV1
vnyylAjVxNYsb5uFbyQwv4lsV3ptgueqokupqMA2l5wUwsSJm7m3NuUMed3Zs+B1
yfYqzOux+/PMwIY+Gj/m7IhfTvtsBpam2+3VkcImMX7dlI5VzD0PktGZnkY0j23a
KpHGNtYMBDVC0nIrysR3zCvcLnE97e/yGXnxrhaDKJCp6cLqLRpNg8L8rl86Jc93
1GXMs26mewOaArxqhcpo/TP4/EebCXs55NcW7qwxxqM56UzXFjTQVPQUvqvib4qx
jNfUH9iumSbBP3Injce58SItFp7xupkzeBzbdawRRqjKX+SLvu07LM56G1WXiVcB
LTUKX/8mB3rLijsK3YU8L45yeJhcowDtRZc8wvkp4xsQpcAMnf3TkiYW9ABFDDOl
6i0WmfzLbroyTimDRzlB8rTKz583YmA2inrSI7nX6NR9186C4gtMl094HvETZCUe
QSyqU97RZeoDsOvGy9XC4CMdiQPKhNciLl0k7WTiugEDs1HWsExUx1fDspCdmunA
b8ZJXIRw9KqhR955/3k548GCBN3ZOrRJX9DavYd4oBTAken/H0jeA5D38C+1VtnJ
gJ0HY3HL0wqdeRCzgOiQ0JwhQjXp5z/yQNzTJeXFRTkk+t2q7VSgZVKkSN8TcTmv
GosTHttTYfTjvQYShl4Hvx1GdR8UTIpT58XJqtRlia6lhPIqJzz3AtwG27CGI8gG
HuGDEizkN5zk7aOJ6eEpun9UR6GOMp64CxTKavA5sjaS8zTgsPdnQ+m3skj9wb8C
xZ5LRVf/KqoA4h2lEDGlIeaY8ek/jNzGkziDqZ6bWYXzgR/fDYeAghxELzuhdpL4
VSUR+1csrWllW9qwGEsn8ArIbwE6T6JZIGZLCFwDWC2XpKZOZ8lP3X4nI2M29kcz
Eyt3mZq84btIQ+yPPFI2L1vo+EUna4G09xGT2yg8/Z2BwxR3hS/2RcaHeOMGGLMQ
n9kKzR5NgPZvdwchMVu9I51NqIHQqPIJoWXIhm1h41JeeQf3x0oQvP+9BLPxcJ78
fA/U1yHZ7Q48g0YXyLADLDLmkXSXlChvUhHX0gtJFYTSTxjA6xcPNbdQ4ALhLliq
OCpfg52uoevf0SVvkM8qV05udtuKUbFIut9iusQLB252XXr6nb30iWpxz/O8oY5f
ra5ajXz3z9krVNSK8ZyBm7wIygmRRgo45n0G2KXSL7oRhkrWCH9YcOWTIqDn9vWa
qCUuLSQPJn/tk0vl7P5zfent/yFCbtQYP9jHMxydk2boYIxWGTfjz9TwNdi1+80P
q1yvRBsd9LzURZ6i4n926+QcXkpq/Wczuo9UKtELqI2bk5obnxIFXd9xgKpLluhE
HksnDlMz7AQgpMA5PPHMBxtoUPWwcP0aNJmwj2HXavTWlUb3IJlj2f7nzlaMEuxF
SDeG8xyxk3yJ/+C8y366PE9XqHBBVOW/N2eTQX0ClgdHQVvdbqlf8uaDFRrksI47
qxBbd8xT8V16BM/Z8Hm1cIt2YbnkQCFXLrvZBWGzaW5MtyRWYIBOjtNzHnNFGhRJ
XpkjEMTeWs45HM4kp0jO37vNeWF4BaZbOLYxmInxnuSLksqsE4BOkHsDB7ZaZv2s
sW1T8A4G9KS5OwYdSOia+YemhUdculngyEBQsdqVDVWaxOfi6uPqqSvCraQiZQyV
TxRa8mZtnI/YkRoRSZ7VvqiNg2PypuLdOR9+Ydx2AOB8gnw/7mb9OMFk/TjgSVGV
l+f8g2SGuCqo6no5GKc88onPWavKpQf7GRB1L/DmU231mToK7O7mso0X7IiMX2pm
dkVbARznpB0aEp7EmCcTEBzmByahj2gdHYEtBo0R3Jl2L7aBxVK4B56vjrJcOKSi
L0XjM/r6j55ec0TsrciFCulsKZ0Co6/un3BaFwATnVugdvQ9LM+46/Gt6rAzRDwD
8d9yrmuw6DRZcEFa7TipaTa7b7jUoM+q1+dcmnmmqlilQKGemBTUzRYZxOTjVhWb
ZjxPfgC7CKS73pDlZtzHyjqlxdKqmhKfkwZmNbpXvh1JHYomU/l0EbQXRqe87XVI
ntqG37fjjfWBHK2lOkM19bi4Q1Sa2EIasH67B1DB9xTXJeP6JCE0P8fEekulc79X
eBoLIn+i1ipEx7BvfYuozCYW9JidewAQ5XjXm9dZn21v/e9JybVPvNkuU1fZxxDt
C9wbhnnTkTKA4VAFEKa3DiKpK+q/bB9yRXIQeOjtKwaWu3Adl6xHfnbq1CCLEC18
enGPBbMdoaVsfn3XOUCVlIVGocvKgj5jkGJXuV9CUPzc+M+uwnUOUl6JWJMaqhac
FQzG7acRTlb2Ee68VwjeLSlnegyBek2NUoahDxE6NMSeYp/8/AzRjSZpJITTnEoJ
A17Wt09g1jN9fqo3q81wTEf89CjWd4gR3OiAA5drXUjp4YNfA3XmvTcqt4C/zUjA
KhL5vR8bwvqyBkoS7/pF4dv2urlB1Hm6WkN5iSoQMgdaboEZx8QHkky4TBAt9xWE
mKlmr8d4JBzCtDfNJcZjg7yR6RLyfkmHOroF4jP7PlCNan9nV9GjqezaFboQvmYF
u6ut42TRxtMMUFmewxCTrHHrS8jpkEDT5dr/3BDpweh3t22GF7MkoWXPImLk0IB+
xBsL15wfNhGGziu4En+7UItIs2hcRNSbSMMdXWOUSJR+wEeYcJ7i23EcCcaR2y8q
+qtNRETxM40cAn1fftqAgv48f+4XrwXZTvMHgSqgxxmKF2cKm8IqFPh29x80mI7H
mUWBM0haDRMu8MtbrIlChbSas+r3Lg8Z8cMtyJ7b1pZRMDksMwjyNwQke030gWTz
KMP5IAQJS4B51LaWP6k7i9preaf4JaPXVFRYWNlUZxTSvlmL7g83pqVRs8A1gRXX
wKB5WRGNfL3Tw1dkg//yrCIU2wy9k2t9TaqtTF68ESUz0+VkwB5Q8Up0nkMcwcnh
YlOyUew+xphhH2KnUS5Bwo/diWgStLoUgD4kg1fTjyxbwDSGxEWegqvfdSgELoVw
UIai8dCLlbFWWPXV3jN9Tmhydv6rvTOJCq1vMp5jsH7OLQZ2BxeLOTFJUD/5oHYJ
+XX6S9mZKgaYyDLDy6xAXLMPQhKX5WA+zHJgeU13R/17hBERTcF46xHdqxaXsNDA
kxzturwFBzYUvP3c+l6KaAHzy9PMVu86c1pItBfNXL/OLBWJpGRJTbdG9r/+Y2jZ
g/JBNDMaKkFep8HhBxavJJtcSYCKporXqZjfosXsRwK300iNRoT4vC3cJlQ1nJVP
HsmXdRqkzes6frdwJWC9gEmKVkbobtdBZawgLXWsxxuteV1R0ka/TGJfhFl9cCOj
gbzJx+MkJygX9W9xoz+Q1hn6moU9opiCowaGhKiH2+4VP+fW5GjuzZS2g94PJ/J2
RYcMa8J0dyhZAQ4+j/DMERdd+GZsjz0Rmj69o4PAtgFeiuIG3mk8wTfeDP8Zk0C2
RHxNo3hiE/3PJisTYmg0KpX89DMyXySLQ9YBCfI1K+gIZj/eWUXunWEVAWqUrgaF
ipIlVA6Q7jGNqz5hZSvrhNxGNLg+auY06mgb/T0i6X/vobDDOo15BSkDrpFwD8lB
GgidL4yCWuqb+K2TeAT6UtdSfFBWrLwLhx9McXQzhGTabBT12VwSVa65cL7SgGQI
TbD5vZnx2ZC5pqrJc82DZCJ6efm5TJ0D/N6Mw7gAadUhOIdXq7L/DIGqkNQeXj5z
G+dDji3GnjBbVRvULEzHswUlQWqHcUqeif9CBF+RMVytnQ/eRJPZO9QvohPV+xFl
Gef3lvLthsgwKZC2lmGydnjma3epislAa1wl6nH2503ko6e52H9sqS9sPtwnfqKo
b+ucBk9cuPaYhmtj6Z79RLT1dnBfdZIU4csywqCj7u58APd53UynwFl62KHc07oS
CX6+U6FSdIx3KBKtvpYFurdUxgHgUE1UDYZ/buCZrMDjXHEfgrCU63ijJbkafn1z
/6qH2E3dazbKRmtJZKtMf6LGKlvgKWnR9nRPjEHlnvpYqjIBDo4hcKnR6FQ+n1cf
trqhlNEAgkKq0h6Rg7PcqxwzyQi1Cder8UGOh2LRxl2lYE7m61V9tN3GcgOJbPtW
94xCe7eGSK+Ag3O0hE+L9CG8MpZqOoCixvXOBX1saX6NoclLLjyQSAhGGk2M45x2
jGPnnyDdvHIwFoo1WATjkK2S1AHdx4mcLkb37ooGhwyCKjKIZKTY6Rb3knMDPMVq
v8bFStGSVMFCyW4H561A4EPUJ29F0PnGhdH9jMu562EG6+qbJ/fUSPrLg7n5VUQf
gdUjnfuFK7Y0AKJ4GIVSaCbxYZy9vT0UUHnt3y8LMi0tWyuXnH/NKkfHtaxxvCts
M0WRZ+icCsE7KwfFjdiWUWiO/EwJxPr88mpOfPdG7QirBEvrCLHbFSsu/TdixN9E
YuW02KlBlLbh/SuoKIyrJ8vxKt+DsE58f0wi0czPr8HWgtWHnjBBWONxih+0NGiS
pA1C+pw255MJD6Hjfb4jgb68cKEIGVwb9t1I1fNNZKZA3Zd3snIsgKJ1IrW0PUxn
RWAJtm0BctSMyBBUWi5Q3Kp7KGFQJNeYhBEClaOyehpXKVt9bUoT4gCsZNvB+u2P
MjXTAs2rUjo6PEtaH3tjCecb0GzhGRMcG2Q00SrqNUMIfMGw1E7RUjDKeikK2c9D
mIbEs9wMjBGQruEpgDGErp7RYDqTNsChGV0JefE1EaJhuIsN8otA36UomSwhxIWR
yBAPViBxU6SiqaFunWiWo1pMrZrQE4D+WDOCv4yNIzZEkta6iQocSQMnn/3v3/jQ
9nipBnFeqmKzvyIn/vleDBci20dlQrGSqFl3pNmHlw6L4XAqLlswvH175FB/hB4q
Thvf7/JJjtwTqnuJGCfXaC+/Rdm44Ol7PuT/n11g8iOMyGxY/vzQ80ETyHqyQOGA
HACvQsUw6JK/hdXJEfl7Wp4lxCjiEh2FTXM0mDmhQoXYRyFIc7Yf8YzoTjLQzZOX
l+Sm85Lz5VS03H53iyjP4uqJ60ktMr90kR0fDX5DYXoLtOOJ0vfx9rMFBY+71fpN
sQ/i5euTVxKakumOPe8V3Dbl5/LYrYM/0x8hoTQwGVdvOAXcJTDcFR1Oi4ihAHjM
moAofRvL78Ypfd+WamIPNuc20UyjlKvByKCp+rxi53aUteRCB3A54n3+eT5Sl8ov
KupEWe1dVBMBYY3HZop4rKqEqXk9Mu7rClqcIrkukgVzUWGH45vHMqtNqI7p7uVw
3wzPc6qiZ/1Ui5jfzBYGNVtsCBVZusE1YbqFwT6tHXGgZoybS6QLnYfQS+orwuUP
GLm9OQV94MUpEVRNNz+MjB0bHUUjzlQVW3YBNSVzp4QGS7QrOUu4PBojlQQ72GGO
ug2vBVyQQ0RZSETHgkP0x4pRn1ph4gU8UtB9wSVTtvOdtGGiMpBQbzEaEt3vHjAB
P3WeOzkNByS53zWq0ueq/dMfJ9s3zCr8xAP0OfSFzWClD8rRcrTKdVmW6N7AYZA0
XiLZNHlCmDWnAuZ/rX1DSz0N5IdqvKJNzlZYaB6vD87n6yZfigiBK6CWWvxKiw0g
jmwvTiu4WR8w4x8fqH1sriJFsLq07W6uCJx72XMmjAOXZLexVdQWaIttSfDyoYjA
lLtE3zQZ2HCo2/jM5VixUYAYE4SAoXj5kQlbjORAOTvNqQID4doCFbAcpdkMJPdE
7Et+PZ8s8+7/TQUNI0w32yfjnwbE4rYOm4rA0LHK4MDUUsP3RGWrZGjkF4UNZpLp
JiPFhXH8VAdHx7MdazIoPSFSgcZv/oWxEsxiKbcn+8ugGEKMw5GGtSCraMgCTjzE
O0IBYnHe3o8HnS+ZNw5hoL9dWThkbqiPPxLtmnAvNa3BKkUgAeSmt43KgfexphS1
9xfrTNxlco4o2sdnqYB1yoWlJxhfcJ7qsbQJYrRqphRhCXFx4lu2cd9OOWKqW1HE
HpXQMJETMsSLFbyskorKanSZxvVdQMWhqz5SPdAcETn/OUzHud3Bg/Zbo5UNfoCX
YyETxtYBolDgbtV+3ECP9sCLFagLsMyOZ8sTiBV18oOKK3xwsqhglnusYAmHbNbb
57NR4ZYbE1Mp6XS3NmLnlzujfIGf5x/RhCWMetYMGv6WLk1IXcHF6mJSsXrn8cu9
xk/cu4Bl11OniS3Llb60XIP/J+4GL+2sx4FMqywKihU4LurZn/M9NulsMMt/ondh
x3IecTnR3WwwOyrhqtFVfzLgKhBMHcpHakvKIH1k4SQeK8bfxDmBAQebIvBrBvYr
Ngb5gsSMguXf9ZeTWCbCYeBdVEIdxucxWHZ8VC0o2Xbw7Sfrta95piLso9tsC1lb
HPqLSwn76avOasMp7cyVxzDHyIpsL1y64XZ6SZ2tRJYv/VH5lhAxQJgwXX0K25fz
E53MkgCJpQ72dMroi3Rky5lvurXWqACZuUSFCqZvHU2uXZuulEEjyuevinlDhiRq
PJsx2pBA8ITvY0u7CvpZ8/5coufxBeqHus+kx5xkkKHZenawIQt2n2eKU1g1ZOZk
lvBT071f3BAtF0PUx90iop7a2UtT6l1o3esAZZJToI1qsOUEysMe/2Zb5xZ9/QIN
FeLZdaNMeGE5oBfMn3J4LeKkYk3aTnwC1S33MVNy+pmu0T3aqWw7G2CZgy+2bGIy
TD0FzGEQtLUN/HYm7vm6KgHR8khUBIYrEDO2+Zug+MFwPSLPvfLY8c+ODQOmvjWn
Xe6u8mz7ZIVkkkayUOcvhy0e9su6E1mmRKdnENvnEM6GL/8lRtyhzjcUCjB/5Mn+
uJvN0q8XzNl47Exe/7j5guXWFaZQFyxSFcTP/1kDRTfZFOoHGFR62l5V0bIkWUs6
T8WtmZm4r5L2wWlOChpjwf64OvzwCoDLVljOMTtBX46M3hZOY7HlNp16vN9L4I1q
5xK8p+f+au7GoG9hMna4XQL5WqkbaHRFivwHkK6EeAoWwfboLA2y0IrYqPL7J6xO
Sc1aOwpqYag3fWRhStla1JR43857is4SesgMoNq0ANwOkYGa7y8smZxqosH+Ef5c
RSAI46QPRoHioisoEUWYMal9nxxjV4w1zxOQ1HhkstcG7aHN91TCI0oCI1qRrVO5
Tv+1Te6JcY1nVlU2pTpuMyDxZDHUgeZ+/t2rBb98qDWbOJ7xqXvvI8ff9S+jZXTT
I8vBAAsKvcPBu9izf0vbpgQo/5SQJeTvbgQlbKu8URWmVSmPO21uAetl4i7EjYpC
CmyjqJhR8KU+dhKADQWYVRehOgLw6wqFVY2QA0aIEw2ry+c280Mf1aIpoXL4k4d1
cgtcTJIP3nM/y8q1x3A33p2gX2RlewYiNQX+zvG5nLIGHE6O76U/rVHljiKoFk4t
lbsXSibSLaxCdjKQOW4G5dPmXSXPgkpJrxS4+evLvitDNpD70aqcsQ/U/NVFkqG9
sgmI5oP9mKrdM6IjSoGuHnTw4KqsObX/FYauuPPKuWJRsaYd3LLg/5tqg6GulEnw
IFkea6MchdYvU8dtAMqf/4Y02nPkL0L1toLZ/u2sVwT3tVzUV3Df5s3wPbCz/Z9w
jCjqStU30/z2CR+AaJgoQcYQjRnA8tT1Q6xRHmAjQNKixbOh3Fqec3FIQ3Topef7
pTFSPtjlyXWYJvLZafM3lKy69u937Q3gChykVc8fk1BQ6Z2ttDDb2XOZVubsRl3F
qXWiUNcUqSjLHhSlKh3V6mgudxSAv0Rcfoqt/Zo/lY79HR3DCdrnAAbApY2nzYdb
XiyknbHN99J4Ya85NEqWEs9HkDgLezxQrOLXEodrpUluUeAXhgneXZcPKXvMcopa
quazdS74mCbpWYT0nZoqkPsy+V23B2WeTKQ5nEgeUC6Jz8DcCmMWwO2Jm0UoipXV
+iFMsLgYuO+0fzDIJE29C043Zd0XwBs+lqz8lmVZ1aK/nm3jO+hRnDiBokaf2pfH
w154hp2ZauaYnL5hSd+lpIPairrpcdCDTObQPV9hhW+MlWg1XCQ5sQkCSjKoBx0+
fwm6+dDVcYBE9b/0yt3agVHTDpIE436hdT3hntvh5ZR4CDOgCQU2mCb0ujjVKi1T
XCMrzg7bN7jqkq4+yFwyLhs87Tiyfu7rKQGEoY9h8McUf+pz8PvLEjnE5usf4G6/
SXbTc9QLu7iF6ELZoiVwP6JeS5FMa+6SYZKlQPBhdun8ww0vk6SKQPhNpSFjjzEd
bvIrwh6ggmmiOn2IcH2htjAo4qiS5StVAvF2RVYUgoXs1y2DnhUHEtsLmGr1g1nJ
e9r2iwVC9e3NtCDrwEqeZWfm5zjxFTqwfF5ORl0hG5YBElThFkqz854m2Nufn/cE
pdn1etOdUo3CQYLuZqnZ/3JL8WT55/mkxtn6xYV98oaSOUXJa/drYbyOXkzzUbZP
wPRiGas1r03RuIygws0AnB+amWLUTGLiAiRvhCZLAvA3llvbmzpZ8XJvntWPBrNY
vw4sg+lAh4GVdbJaNlDq6/1h3Yc/3K0Pj1eLkI1ikcqKEwV6B5+xBLAZkV6suxRF
ZGILlnAt6CQ/5fCSehYubDnnlPzVMzfvyp8BpbeUHZYvrrgDGJeolffyWmDIvs3J
m1OIQgda8yqsoRrqueNMKSuwJ00Mylk1x4yzIkwSC+ypwi17Nemn50yoWz89cZa7
uBCjnSLeNqATUgh/GknncAVb5xdMGEglS1oU2ifW8AiE2JMbMdw8+7n40hk2HxK4
9z+k9j07ZMaL1OoQg4VV+f+6lg8sd8DFKMrw+rNh3r7aUA/H8iYUnenkAJF/De/h
JnXNW2VAigYjFqKJL2eead+mVb6crJ7QQzrZQfc7/tJPIaY8AOk5DE5lO0iP8Oec
leuw+2r4t5P1Den6N12n5sgDPM2Tuoc5zyJZwBSjSR0Kg+G4ZRGiTt3Qp4r00tnM
maEP+KJDc8wsykQEwRwjAGHOdvgwGaNcRwTLk1HnpeQin/y2mwZv1rJ8xhe6rHvA
I7DDql+pjslbCtRVKKiF+UgRsrHQcYHMMynCmlP2ShXD2NXmEssf+o5eayXYUHb2
A6HzT0xz8XE1RIcbodVCO6hHPDeMHdbap1TZvtvhOv8Jm8wq5KmHRo9iOSIWcaLQ
vHx0xrE9ewGMjCQLa0kqcMt57ImsZlN0W62eLcrFR3xZ7/3ee1r1nsD7nW0voQO2
9vW+Zt7ggdmSntUoLF6SmQ7mL3NyNxTJYKrLxPsfLt+qSDSu8/Fh3wwDCNdPcwE3
Ac4wOj5+41M7YmW+SK31uaF+oyxfSWXewTnqU1deHxiIMT18m4uQCz1Y6cT6e8B9
HyOUl6PPz4/lURZ97WgMrvZSDRUiHRbDYb5w62uGXZBgD2jQNHgbHgWox0lNGZBn
9fnTuhIDVZFZBasae79ZG4kJRBVeBbePk5MJxtyFj4MREa2trGhPjZt8ZH3+/u2U
fAifCgRUHzCYjeM13JZ8eJEDJIPVgWjNc7X0bel8vZP+lp7TaaWSol+rfMTu02NE
g8qJcBMyqDjnNK+YhcuaxW/MXEQaJ61uEgjF2gaUp4LugcMyV8et//uMhYdAchrU
n69YzRh8dwfXhLQigTp0iDzG9AyfYAIimhwfIolMrJMjvFdkJsoirQHfjQ1HZn0a
lW1NyXKYK1MfPpDZGpGyIXopAB9vx1fLdVAReIqxXywbEbhJplcIYmfX/L2adD4R
amfZTb/jZO0cOEuwmHTSwm8DkOXBVVOt79Ve5LUD6KepF+WAFk/a4DWgM6IGIEI0
q37a64/O/g6jkjF98ow7i/wXiDic8zqTpb1K5DK6tL9Loga57YmVri8GTVMuKlCI
uDQ8vjIhaW1nbGQZQQUFPMXlaNSgijFWpQ9jle7uzdDhuoEio8j61On5r2unct+6
n6CETgBUHxd2GU5QF+k7Vzz7yepYQlR6ZZ5UZU9ktWRcYcvJDZGtpQ6olA0IoiFV
EaM6zHILXxSTnqCb+H9/y+FreXQQdISSpUucqNQj+K6DoK+J2J4wubx2xywhLzCk
wsA4A00H5dVsaGOxyIFdK0Jsoklr2/mxYM9GC3msyhP2iZwWkGqFb5IdqyDYQ6o2
zSOIU+zUiNGeuCyfTxBGrAFsAMlAkvCO6YuNiCe5j1S1B2oh+DCqqHMj7+6Arj2/
CAxGrNbZeHxGmugr8JMDxMNWvCoJ3+d4cRXD7DsCOjJa64BKJE2xrMrmEW4Lf9WY
tnC4mPkibeIHqZQDRXOpLJXRSVlRoSj51jVhyTsqLRpuqgTz0qTREOAevBPQHWzS
vYxK1ttZ6lNuDTHuAFohI7aXb7Y9FiJa9zzTc4yL1NUw40A9xup8QVC8AROEqfV/
g8iSaYh61rNeNfr7NPCRS0fI1TEagkMHbzaptLzHc4/tczxumKHHA/Tfi6PhECo2
TNqJICT6z88O2E16daewxKX17Fe4BTI0ajxCiHmmqvp8iX+Pp0URHJ+y8O4JksbE
O9FIyfebG5/u1BFIkGEz1fsVGZ0Vg8M9SPzKrtqGnXwpe2ksYJDz0rDeF8wsUPJl
NEGsPiUBAl3+DzGkZPvOmnATlbKSrJjL6yr7toWtTtsw/NiUFCan4+Z6rjGqbmFn
CtAfv/FCqhNlFdN4W9FN3AtulSfdc99rWMZCUUYw2IE/uqfic6qqCdkfWnIas7ma
jQI99ckOEDqbuxHUIGIfnhIxgSiEgau1VdfEXQWf7auHJMymRvHFs4rGUJ8OBIpj
9IEqLiO0iJ//UfernqWk9oPVWGUB/c75oArutv9Zzu3yJQoVN3Q7gSVRq7z+oIVk
7pCBfjpLVVfHqjO19YV4ebTf/PcnMVW1ek/SWr4jO1YpGlv5cm091lczEd2O7Wuc
7feZWkNwCAeWUWGO+pn2xYDG/StN5JOT1JAVagayp+MjiK00WFIk9dhJtlZUXH7/
LO5aNs0V+tHkYXt7F/jTbkcsoGeZNA78RX858vvMeTuIvu5WVbqhwWnM1F5KiH4z
3qhHcIClCoBXyc8c2lVsuhHTDz4t+NvUSkLGTQ/ChBOtSlyt/jfDFSnMWsNYqrqC
LVxHWtda47pE81EQzLy3UGNFCjyF6cAf6RRPn+pqzuy2PO35EgP+wy3XZTURhnph
jHSMp1yi0Zn/1c4xieR5q0owSk5Nhi+1mhmtzERdKsr3hRcfBuWkhtchCccRhJoM
9KeBpk4OWEK5PtPDlzG8IKW9K9D7YbO0Ab2PBUlVyTMtwtBcPjaDAqFuqjyrKEhO
XZAk/yJ+a99lbaYk/fvasBGEpVWp9CrefAEsPcVKPIwrySVd35XC1RdfXr9fapVe
o5nSsSvVjSELLcV/T8DDn2vcl9WBwc3jlNZKvRm2MbqA57aMDvuQpNjDP6l6FeBX
YBlGYe+090a4Cd7BnabD/op1FNKZ6vXOybR5S3PbuPTRiPinCiTWjEVc6zeGb4dj
TvLOikN5xp81EEn5tVmADPdYsPfOfrHMC6umb+J1HGoVoagdNqu+baCwe3Bjcy/A
7p0KI5Lef1ffJ/dlTYQYqOeHyQ04NlPWxNtlIeVAqAF9C05lb5d7aSprmKV8kEkk
1/NuP21zH93FeQEKoKM0qwjudih9HzLINLPHnYoA1D/DrhIkUEHx9J7Q4gonlHEC
O5Bum4G+t+q8QnAUNwdidYt5jFR+N/BPZcN8/cv/NPDsPTwrVBMbIl9k8NLqOf9Y
nJbcxK3eU1JfhamSocI7lEnyvPzsmB3vXJU3d/Or2WskemL1YlWYp8CZqAdQcZ+6
D0bjQ8uLV8DsG5oanbQMhICSyGFmZmQphmiXbrWZpW7p/47izgXG61qCT4FfdsAw
AmX9BVL2a/l443bhQTz6Yq8XhZt1F+cKmeJlptcVtvK0OfQtL7woA3BTv9M5memd
usBvzDzhWA/j451SMAC/pf4fPp49RjW3BFMldnO+dGNSvqhKQaMNgqlACMGc3+z5
ziIvnDg/oEOIzDVVE1ahtC6xK8fgoGjQJru5D2WFwZBr1Ogsx7PgtB+BiCnv+4cK
ds+7rFCVCTFsecV6MNAPKM1cY9Q8Sv+bokCPoYfeheHqG+fLmQP71qsakzUDbAqY
pZ+28UsZeDQmi+wyigAHc8My3jcPrXbG6lGPir5OEgj5rDuyWXiXCD9HiXdZ2IGZ
KnAc6sHW2eN534uc/PcbBr9LJtrYERiVCjO3D4gNrYYtblrid+lNX2m7TwIHPnqC
4L4TdV+jQjpH4opsi7KWNTVxLl2G6WoIDpn/Y/SmSwoaykhRmKngmiI2auTS21bu
zp7Tzta8/ZkOduZuf4PiMYF7RBoM5iqWUgsB0qFHP7QqtO/9EcDujjLBMYWGVwE9
0t190Dyjsysw0X7/vjKRd7KPnujBySInATw95J1kvqtcWlKVCF+7ozeuDq5MJSIy
5CwT7rr5i9HFGVZ9ma5AM/o0IekbOxgdbl7SASGURUr44ChItc99QGPA28e/8fnN
vp15O2yfxSgAvM9nQot2U3UaGic0Nm8ptOQq7o+qSZojLN6wpfRJb9wqNAawdqwn
LZbJZgu5PuHLrL5PnJJOiVMLTzzPQU+hvSVOBvLZyDwil8s3s4ane/LYzkxMC05d
wl1MfuPcsmwyJaUL5rXeZ0aTqV1rlLTyRwQlAgx5ZJFgpL2zWgGkQOSeEQZr1BAJ
2xLwYu8ZpzsZYy1iSuwoMv0/MOssyJ6hpNb8FRW2XENch0gZvMqJPmlfG/X57LU+
QXS4+KySFZ/vNFu0I40t4FkC4XxFpb8D73SkprdlV+XPavKxVFtsGWXe2CHikoZK
MhZXStLZBPyyhUB4hhZJGiVzRYzE8Gh8Z9GGBUJd+NKfltYn1eDYWo0CE2QPIZKV
r7EQglKinTlB8IfQh4A4puhaMv1zbx2WYVwyXS5lBbXnfOoPD/ikA6pmJgZEwQJ3
fMhAgUHpJv8ombaxZFgdY+g1T4aSki2pJfd3FsDqTwN2fDrlsGOXlaFn0nqtdLEt
KsCEdTcMRihmoFyvY0/jOCwkmwnV7Ig95psQwLo6hM+agJ2Uqe6etGN8DgM4VW/v
z0BTbnJTOcS1Y+xzqLoQsVRfFxZvpwGimof2SpQdzUxy6u2J5EV7BpEJZn0ZbRLm
h/4oCtV/K7IEGUV97EAojL9xP7ADdSmCgz5wGSOlRZ4QKGfNDRYS89UNTcy+XLHz
86bBbe2ya2YGNkmqZ720TQPr/ZODXRP9RjVl+7pUfkOGJriQCGcI83vJIzGLoKw6
oFECemp5TEe8FvWydDOLQ81dhG7fNeLOwWMBafUDptTnG8cE7O/X+hDylV1PWcAD
u8yOIiewRPm7j4siSQQ7azeJsZTpADCG5vK96u0Y4e4v/uODjoeB1rw+okWHYKoH
AVBvsssBRKiMzyEQHlsNuucBDfNpCSL/TJ/mFylmNjUAqYhbbVL+6LeyJ1NtsDlU
CujOz8eMPFzVc2yxLE0/t84h8o7f41dP066Fjuy5M/xFM+piwqbEQHTSGt/pQFDr
w9efNq7hvUpQrl/sgBaMk+Zri4s4lchjcf7eRCpF+PLcNZ3OGYYMDGDpg5qEGOGu
s1YmQAgWfJSKkzKRElLwaJ7/AsMAvLJrqvBMwqXq8u0QyyRhSrOO/OiOTvD39VmF
GF0K3pwB3xiZHk7okuFNHInVm5sqL3HMnHh1fY4zc5E0RX8M/qwern6r4Fh4RdqG
vR6r32hGkU1cAgPxJ2qcjtkJL7oamBHjsUxE58U5A0RtFUdh8SLy6gSGqZvn2+N1
vw+tH+FJkxZrB/Z6aZEbbextuxB9YjXUAj4je8KWCwJu2Nm+dsw+FErCqp4WEIql
Z3yw4zzicsDqH+RR5JIuVbUNMTGMY2WMo7q8kgeSqh39DUGIPMQf6CVwnzAfYp3K
/4S2emx7RXol3Ryaq07xg29Rm7jBVa8eKsVYa9Z9WXmbFfPvb14a8/KbTzLCYkRH
GRGyq0wFyc3UatOBQkUaX55ivrR9dV8/md+f50tr+wXIEKJz0pPaUpPz7VCz/VhR
st2Bn+59kNIS5FDHLfb2ZilyMH3GAcesNGYX8+IuUS+1/N1DqKuwdBpvVP8tEcXZ
9T4s1RaBcCcjfysIPHz6onOTXzPvGr2LPpaf6lHoChKvT3aojcep2j95FTeRgBtN
6yp3Afoc3YvGxnPcvAceJYDLaOIxVV9c7S90ojrPPUoR/Lvf6QVnn6p8up1cgYhK
IZhDcXtkYISDjSzC4bv3/5MpfC3R4BMcUuKYSYlWQsBko0DpBklBVSw15IPE3AWM
fdvq/bVFBCmP3PHWwUOeTjtyLndt84iFoKh/5T22U6xG+0Zo3qfQKoELE84I0Kws
/Z2nPr0H3PJZFQ1Wv6H8I5BE9enyvzp6hlxpcGn/Twb14MnFdBLzHptjE+38dDon
DjbgqovH/AWiBCs6Q16XMcHEa7dC1yNfPCz/dJAUqgC0RZVvgUarJkPfQHknd92B
Nfw0KSY9pgDpYGZnvezzcUmPm9Bd7LnoERT7Jr+B6TVgvAHiPp2nd8b4VoJhq40U
LUaudzTUQHbEvEOcFJqoyYwOOLFYLsZpmOfh6rwyZZFZgvmahivWsB6qifXax1Qd
VYiWAqjIRiUn/8sjiaFU6fVvjv/nFuNldnYGFNB6wXJ4+9wsZatf+uFUd/6YGlWG
x0xyIpAL3UY4d6cMXljVgvDiUavKjNLoiPKdh+OjmYN2YX87XuZ0/+GZ/XC7w9tI
o6/4DgLATIuJ77d+olHBB3G2vVRCqknMOhbJeyQju5+dHqQOT00pm3AVGcn/KS3S
r3gfkODWMvPvzatpkrdzJfuavR3keh5AXyBsHJqW5RWRNAc55LlfswZfGdLua9tu
VUU9YG5jbzDPDZcTik6/KfyVkz+W7G0T0HqU1GKnkV2WuKpOepTip7URse0FmT9T
E9aqy8hqowI3LRw97j6h1EHOThfE9dHgHlRrOeLVVgMiVk4AbXYcDxwh9E7xAqQb
XXN8WlXs8+c0ebS1n3AL4jp7SGazj8vQViYbIvACHrSEBHv6jkt0LvOnagFOgK2m
CByKGENKFAnOOBRIDE3tNq6BAKAQG2ht/TKSgxcp8XUVl60gt1HI64t27F8LPxmq
pgCfHtt1/3abIm5UREjmxwZh6AQYAeNqqjWPNAY3ybMgsuQeaABjAflJUZRhBTDd
J7F53MR759Yn+VWmkXAypolqFQ/S5Rx3efpdYdJSpKonpmuNFFHlJ8EFAoyQRJHX
O9KSb7c7vgTNiTFTAHuAQEgJQ1V+CmzB3+0+zA3Jt6bHSlPap6qPe+2uPlcwpaR/
ytw1EhhJIHbQcWh5h1R3AsgBOYbs+HB9kiXldhA6SKQ3IYhZhx6kvYqzTFaas7wf
l0E2UxLHY4v8ksMjH8wT1vHaMIzsozjxyo3LEsjfFf1hkCAIgM6bAqZYhtTLwI1h
16Jvcd6m9WB5UK0ulJ0BjBbaNt2ZZS5236AmC4B+FBqpso2PwiGKEKQqYRi//aC+
kuiS2vNWXJaETEJrc0B4hdQuzVFsMFltTuoneXIr5cTf6zu4xgl2ffM3+34ETaWk
LL7UZQmODhU1NxevaLwzSJypiA2gWTteNUOkF4+/+PTfNmAWrGIqcni+yiIXuGTL
pA7r6H8IHSJNlgo26F/CsGL78oNgI3MwIKT8RslDF1+aekFKLOKaX6cR8sP1WIxC
mS5+5UDy/SRREhyfYoU464o7p01M7tfiELtRvelBHTvBZsH45jwG6uHHs8B0niwI
9r7iiuhArtALmFpX04gUSYq5PK7BVE6gPWGrUrinnCig/iI6x5FLzpqMgqJfMILm
eAoZ0ESbfLkaQQohmbpflDNt80yZZk1MJYsI61KA1AJEzScH1/riw5Bxb7fvVHRH
DjDS8K0LIpDGiGncs7JR7fU11Bec4vuU1f7zHrdJ3c1Ny4GxsIRVJO19VJb+zfGB
75iLTdcKlp2mfz9JnmlHDV9S6vzx8gplNtJL4z5p65LVM7JDbrb0ExeTrf2DMXus
bf3gJBk/ODNqGcI63sGcFexT6Hsx2wLfqcsiqkunBOBuJOicZQOLge/IW0sEh2gn
CN5Wj1bt0wLItIKA/vdPsj7hPyUfaXFClrPQUCQhJuDFyufj//f6SNSV4qUbbIP8
WfyVyO4Y8SDupFePe8sHs84WJ8PzkHw4Ilg2rURtcUMZWd7vlLjwbOJ4OCJNxqpM
iTg6MVZGz+a9QpsHYuVd5SP0l99ZEqrlrZzPh6MD9kD2mpjwd1TuCrCmNu813TQ+
yVS+OFFMjb1OFAWD2OuRnQ4OmFOIqQqqlpdvw7GQsWrwniOE8zFKqBDjMXSERveH
RKU2qjiYoK7oyVYygvfwlUybid/Bn7C3GORv8gJm7DdqzJ70OiSKVvIFeWQlqxY5
AjmPoKJ6eoJzp40TXCpTRLRHIQCZtZ+eYqQXBYEhF8ModyRhviXEhco4f4sIxtAg
vviHd3HZMFMceISGmCtI/I9e540NBxXKoMNiO4j9xBgC5AQFdRolDDsONKebzNis
XlIrgNn04covU0V5NwxWHbQn3fe4IAPTItaYL4GPn5+eSwa1w+PGK79UO7+xXngP
Gdf+fDIBXUqVKEk7UsQVuea/99wzzKMs0FQuT/H1G0Mzi4kiCvEhLt25bZgKm4UF
7HqNXdRtOHXCqL1MYVHHmgrKka74pFLGZXH2J9FwV0tlRsaHgmJzF0Ar55W56LOc
yMEU7Z7FS29caOPSniGSacU1lIH9z0rtEosMXzICp85mGuC/7sbc3j7DiYekJep2
VM4J1JgPQcxwL4e4ZTaaU623h25Xwf4FflMhRdp5SsyPA/APfo39PrYzw41aAt9M
AQbVY1plotD28fA6DAF4cZg07t45W8SCDQ8Xl35KM2vF6Gsd1LSRDvNxD2Af+TNT
EVNC6HJkLrkICNZwIs6BKlNOUY684o/cHYWSiwvnVZT1MNEpHz7bWgLoMmhNGltb
CQUuIn+De72wYFh2DaXKRUKixsiZgYu15LD+QASDWhpfIK7v2/4G8kBqf+4emmag
lkP5kbr8eXXWOpA4PLx3SbOe1NVwGp8F6AhuBi8FLaS7MghAxCLmbs0HbxTM2LJ1
pVZI2pRPS1eZAiAMQUUYUwHyLVRJB/9dEdMvjpdFHUkOZ/IU1007KpVDlrhErBfr
QwJbjC4FmzdQUnErlJZJh28CDI3K+bfxaQUi/VPMlYacBm6yOrNhg6/9xBoHqD6Q
u6w7PzQEpGY8dB3IJyxo9o+V3/OA3j9miXyR6qKw+W2544SW5FvyIwRFt8h2ZCkf
VrwN7UV9gnkS983qjmZdxK7ckbJCSgcnv1gob1z8kunIpYPF4BXTUirwKGS0WCcD
FRQm2mOi3kXVtqcbWKo21MchS24Bry4YvtLiIb+q6HkL7xwg0YGsP/iDU+6DpqIp
BYGtgwKAB8I4ZuCO/k5OJz60BkjZy0vMmx7Tv055AMP1/bomq8LW5G7UvRk2ajyj
KPz7QF+aBNhYQuK4doizRuPg+W3IsX6zRqgcynBZn5sXZ024E8gjvyuPU71HZlWa
47pcrfay2d0ARv6Ws1HsQWf7/eVQE3S1p2ia45akdb5h5smgAp/t13R5191aKM5j
0HDChY2tay64+CrW8frIKORmFdmS8UWQuCA6KZgyO2kdl8WRYjFSRM1V5fvWRo65
1RjLe1e1sBAEFlKqd43nNwMczx6Jn/jbmi7Xy+mtuzPzrhLrYYc8jqgac48y7mJG
kj/WtLKEfkr9Sb4mBfwo4CKoPg7l4+rvzr/Lv2KBLCe3qGBq5JL7Pxbaa9TLNH5+
KUv9KISR2noHKnRk9M79muIHiArQbadgjywlsjYvsc18XNxoaQq/mf841ZLCdyMJ
5+sJQxPhqFuKkgm2Z+6b6uFDJR2yWqc0rlJpsw1DmHeUUjtQZYzmhvSOsr52zP5b
/jEG3Q44wj/tQGPQN9hYfiQIcCOucw1rcE/Bbz7DZrHsZ8j9ZAZ2WahdCKjw7WeH
YQTccP7Hpdv2Dpt7MxiAnlbkhE8+EbF4d6mLb6meof/BjofFpBV0xG7kS5BHeG7m
zN0SZhk/V/NxOgg+tIJjjDDACDajcqjeXQNEnUv8AFwmPaa4ZQ1P3tUvYmUrAsZD
+gy4KTaTakfAs5A/RhclG9dXNCGymDhg4fIZzHZjclI1cDXZ2mcN6IqmNLTa1Czq
d9BmuzSl8xj9zOCUiUMw19r7yfA/DtQ62QFAWQa8kWSF7inEmg7Afmun9PGeo+01
oux0d1zwSrjiQOzSr1WQMirbTIkzCQFKnUjkIlgoAwOs5l+EsgShwfASAmLNgSIl
NkAaaoQwT4oIifs9Ler1DYXYxH2vSP+7pvXwPTL8Z5aqdcXdLtuVox87iAK1Txgw
UQVvlnGYzoiPmVnOOmsSxsSnYogx+9WC4iVr1AeLe8usbDLgAOrV/w6kxG22cvzP
oftasIY0mbTatHyNg7YNaiAtgtfLDY2jBK6EtNac221p64MUF9ZoJr/aOgFw4+Im
fmNXEfueppGfVLjj2i0yDBKwlVUt1EaMFU+JefmH08pXaV1mauiBqIWJGsHTWn7H
JLRRE5AdVaX1KXCqE+UQ7KWfHF9WTfUNuxR2/AZcrX/asXFgG5fdJMeUpaBrH8i8
QZJ75QKTkxvRmTuDAMD1e/Pxs5hGahs/VBtz4G5bgm84pY0as5oA8+ukpib0HF9Y
NKqwrFng0o1uL9VL0/bfoocHeKoFI1QI8EbRGQWoAAEyxdzzU/zgJICxyyISswmU
hRU4soUQBKu5R5dga91Qaa24yeRWJh9ovyukSDoxxjKZurlf7oFKmwaEr/nFpOyO
8OBwIQVZ6l3/0DroEZYWV7+jl5PdjThR7qDL8BFSdseD1e8/wx7xLlWLT/4yV7Lo
k6ZD+rlMKLpoA8Nbukx7OfrBPrHZE71mwprhFc86P5iHZeVJZhRwIPSLj8Nj3TUx
cdaPZduvNBgN23mZothTW7KOIAeoCsfICMkF/A1YrjJ3EWeyr2//qvMoyKdOsIU4
a3RN2XjB5clsBQzF6OGByJc5WLZ09Q4v5C/aiErpYM1VfGCJ5V5UggLO3BaCVC+9
r+Kd991gyTAGNxMoiOJXlN7AasIqRIWpO3ns6D/xmlJzQnOeBGFDc1XvxubRck+5
Jb7BIup15Qm6bbATtMH+9rD7BlyPKszK0CI13oiXIbPlool7yKmuHHZh/JkI7PVj
8QdKap0V5uy+qSCfQc47zbnAf290HPesY6rh0AwGiSQWM6048DqW8iucr/PNZrDL
72LTG9MWdDf3Nl8VTXviOWYPoUhmkn+fY1Fx4AgBYdB63km3q2jJLeB/7UwABPbN
44Pjau7jUcu3o42TSF4ZQo7H9bUz+1Oi1nfpolM7seljHaMy1bNaU5+YdgyCncnH
3xEuCi6/BSJYADiF5o9BqDTzE2ieVa1q98i4VbZ0WRV/R6qeWQfVUtZKbkLWWY7W
3F1MtFQGWrCWB8Urht+pHY2q8FgkPKsRc0vksk/yWs3T7EijmiW7j/4KcrFoH9Th
D1secGNIbFZma8facj+premMN8RdAC5MCHkydWDFA41s5EzE9SNvkKvBNGyjJlB6
zNKXRXrVI8BlVh7Mq7vuCvIIo0bdBZJoFBZBZbUjteW9AJSNzWM+BCb1Cma6Tr3F
EQ0Zt18kRgxLJiTPE+EtBUjkdqNnUgMYX4osKgI0hy7ThTNfjTMgTsMkA8B+te50
A9+D9k/p0G+wEguGYUGxH4+xPkjIU2KVWwQ6xFLtRLrVejXCxvv6DTuA4Oia1wP7
ZopMHn+z9tdx//buJBljyug80XVStqSYUdL9x/enedz1/xPAHRdRsXGN5cSWNJ9A
llFXbL2+pTKADjVnnS7WMWXBMWCerkT4ULmllUzdIGmb1OC1sJDDRe02q5uyQphX
yb7ELxSkEVPgB1TqnXncTaaN9hhIWsIx7afPUxZl+MQKH98CwB1awckY8pUfIOkg
K2CFk5E6WV7Qd0oULlWdNuFUpYgIbwseZL5l8YNUknrFOccrwTvUUFNfiOuAx8qx
hpcBB0kiEyz47XU1L8FSQKjuFbzxR4K0+brnuGRJiwVzr2f+de7hZqSX0WGEbecc
BHQN0s9F2VKvQ0B18JdWpLMNA1v5GtZGmX7UamK7YP/3bkFVfmgL8V0V7hRaAty9
OS2+L2+z+adBo/WhkNg7nQEPYOlEUPXshft/nlo17wNSqNDQqjbmrQJtCJyH/eQ1
dPmeqRvCLBZ0Z/gt0Z+CS3uGiwWDyis2U04Mx82h5OR9LcFlNXQwEQdJATj+g7Ok
FZpumznMDOAPufXkberGcrbxyK/L+duLdj/XCCpM45DXwSU8HxzgS5GkayR+GyGL
6Thc9lvQlbHUJ8yg+Igz5Ob5vPetUGUYstvXTGLBAjdCxqsAWZJi1LSse7n744nt
nLKaHViZRlHRM1zzBl84pR1glQRa51JRr1JLKxb/N+V9uBY95pVRiSKRja7JanHC
dyHUpyoCFZIZmKYoysTlO506sm7x7Wlhyy+1XFQu4wy9DHobgY5XSFZ8FY7cIrvq
tWYjV+8BGf/kVVx4cNk1mTCXJCSft0Izaj+TBjxGDe/sb51nYLJXF965AwWBkU91
2Q8JYQQ2OOYFmm5cgzN95xfRaW/crVkBsk6TiGT4ftvyDRmm9fRu0sKXqOyfUAz+
/vtU/YfxZxgDwzucsjsM/B06QuDL4RjYqP6ZNSJG8MNPldwhhdRfDQhb83ls9ZSq
s8Ops2PH/+jX1F93toDtuM15v+FmByrKIUW+kH1ttbwWcCab/sl4rAJUXftcp+rf
Le7Qhsy+GZLbnYfgaY3rFsK/U4nNX0d8zpFTuZv/1zLNt1qK0984OBzfM+hTj7wR
lhLH/hBSTb+Qjup9wuRIO2GbI/+dzU8Hh0uVhYRhb2RX6Y0GzycAD9KAVMHHqWCQ
kTXL9KCkTclY0Qw1xeRs7KeQrtKZ8uOpRnYKBHX6XfIydLsTdcv91+jD7s7NgjeO
OF5XmEi4dx0wQbxcCEUTThReK5pK6Xb+3ezvkNVeSyJa6bSGdp1z3eoS/hMcPmZI
a1O2f9a5q+fQwfgJYtj10oE+gOYp7V79HIfIDEaJCgSewh4crZm26gLlR/xZt31u
uSbya9rHHFZonJWAkOc2zeo6easxuD7TPd7I7GqExZb43M8GvEZffKzDQ6vevEez
//f1MztLMqSpKAfuhHIFR+a8y6+95uIfTE98o01U4L3HsaitYK8HATN7Z6sVTJ7n
ItWSj/0ByKBiGxHuzbClcvTxtkWBrb09XwLVRg66/vpK7C1cKNgGvhDFm5FOlsjT
4exx3v26FAcix3AnG3G5s905LfN7GbGIQYOBIQfhuBc+kBSetOSPKOLCJmFHqg5C
gyIvj8NyUijBpA9djdcSNaqeiZ+c7Xvo3OH1OKOoPveRS+8Ea2YebJUewV/BGGE1
nd1T/7a91A4OYl85k9HmshnP0MZJVJv2590CMgIG8JfaMtM7mI+9EQDie+ljRmmp
SlXFE6GpbUkVSInOF66bLNw1m+iVeZPoRBWpUqCa5hYYaZtn4m1WqC7MMjh2NHGs
WQH5kv2TqYK7kzZN83mAwSAC5+UX5eVl0Il8Wg92XbB2CAoadLy3ESzQqQsMiYap
3cFRMA2D3BibcIex/nus7Ht6iOdsCAfnBuRdHWkdZ5QrA6UUan3mga03Pxf3y4Ah
r7XbxaPttzSTcBzt8jl5Nak9dTqvnbdte0gZALWEFt0vLrGNWaQM3Pn978tCSten
q3z0T+IuxCNXjr7FiI+3RgewuLn1jd3fbtvTGNaEeYuYoYeb07MYr0RUiYK8kegq
GQrQJrjqWPgY3G+fhhgxoyJBwMGIefy1Ov92IY7A5FeqHp3GRJABCBlGwaAhj7ai
kVLe0PG8FEb7cPWUBetaUclNPBdcPBn1txbhZhKGtcFafE9SmFga/+gyL89PuXkj
GT0t4VjrT4CMC2nhZHqPKTI0KnyF8cB7C3n3TyAM/sNvptnjQrCUOm1SG4qmU+s7
zDWk+w36m+yKfVq0o1aJwKqy0AAyVKhHWHenrODoIZy3IDdoaGzrZXraI7RPo4XD
JSZEVkK8gjL1w537fwzZ/c5LtQwkiFcdklzkLIm3iwSlGvJQbWu+NhJx8u/t7UJH
OlhFpW4uvBzbeph5lZ7o7Rqk9guL6B4d6LoxmTcUcaOtnlqFNCdaT8/B2+WnUOdl
IV7b9ln05NAjfvXhGEA62BQacd1nHjcTblmcyLgxI0XtJkt4psmT9CPzpYxeuow3
va/pq8t383BKzKy+aPKnKv0xMqxCQhM5u9w8L2tpXd6CHq+/wJYcS8kvMCBXvIAX
7MoEy0SVs4ul1QqBSNUIIJSEJgTe7ducq8i7ErhAgGzata34up+pvj3c6RTVZqmm
0l8Nj80G/inFS6dXv/BzufvOlLh+YxA87h/xSEbM+L/PPyIUYULr8SFucrV49rGI
C6ifcDrRyLEGOuzwI28zBOzxBQizsldjYTZWW3QI8JpoZELMJps+pHDwN+hiqPh2
`protect end_protected