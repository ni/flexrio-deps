`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14608 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4sSkgcOrtFFGmnZEnVbxgx
+l/NC0KUoptgPj67g1Rb637ea0Q+aslXHcQGJo7yF+lsHmVJnnZMJK+7ErxY0LJq
qSb/PvkxJq+gAqlMfrGnc5trBBftzaH9La/jF+XYvbB3EDZ7eT69bfQkF4Evm49A
qhMBZxOH1sbkFeeAaaVJ3zawaYxjfG0rvkob1L9NULwINcIB+KnMrnh1Vs2JzVkg
KWe93XIaJSEJkzXg6L6EYkv+ZZ/GK6ObUtuwzFY4OhaPC8b7xGeYBhc0iw0GevxR
1MekeKV0ab8w7wNXvwlTi5iDbpJMfpg6jkmkpqezvoXYoH9c+IEsk6khNP5qXDgS
A5Dxfrb0jL627r62HJDD1nGMs/lGhZaE2wsy0umVwf8pBJyzOCX9WqnBYT0EX1R+
fJHpS2Q/S2xjlU1h6nzzhK1KU4lh5sXy0WZbqyuRFiavY6UKzsCpBcRyC7seVPL3
vPy+naLE0vjP8vVugbswkDB2jVFeOM+SDm7gSyxZTVW8B5nTF42JEKZwbd3X8bNr
qF2C82eEVxMwshFhfXt3ejx9C9DjHSDMki/NvAB63BP32H8Gn881xj3a47rKYJtY
wrd51xJfo8iRNK1e0eezo4CBFVtChUXOOKyQI6gNSdaT/lXagvc1XP8wzixleMvu
5kdOTpTsrciQ5PKViAqce7Q9DAX3Wa5U5mp6BeLhEra3U8kxfzooJfOUM0x4wCT9
1LWEgUqMh7iSeFUTA8waCPWvJA6oftUpajWp2/V88q9ZajkVH37g1DuHqaxhCSnr
FUgvSbU/aSscQ2bERAcR+N1I87Q3NM+acrdxaiJSYKm6yfE1w0j0ucFmC3FXpqn1
SkHT1bRxG7Mp84w05Rl8iqRpwHFQu/zGXYgKKS3CkDUZg1jbqwo1UVyXTCgWTj0z
fZApJce5/9yt2HQZhAgppNOJ5R5tgEA9IAVaGj/XZMRGBD0zB41WWWdDve6pOMSu
qLFDu2UD7Ki5za1neMQqyEcIdZNl62ESqUYBT2pMblmKXhjxp80Dya6qZ0KZG53F
x1tkF+StQLLhuUBAIRy2SI/xDhzDx1rGCV42fZ1rR+QY8heVqBxPBTatzoQvTJXK
5ijLIcpxYPECmMrffmH/iLutJWxat3iB1kPXb8zY3saSg2mU5r7mcvZ9q6K1VjWs
PDQyuOiS1nxP+uFDyQHGa7hTND+8O3z9kOekFp+OSGk2+aXj53kuTFgD+zNf2yYE
7Bq5b0v6SUyMHWm7XeXUao86GeFpH3ujnmb7gUy5cavu308TKa7CtGMKZIXMibEa
m1VXDQUM7RkwF4YNBmPxRHawbjUDbql3l7hlEZHSlGz9PdMtv9lCyP9nKXCeFo1M
bGpqwpbC0ot9YJOVG52S4uLVTt6hhBg5HvnxtRcc8E+oFfzybDl6VXiNHlzyDEyK
/r+ge27GS9r0uD2JCIS7uGXq9TkZP86Vd6vGDNh8N+mOU4Y1yhCiYuDtb16ytwwd
qB8eRQlpUdDsfwx1S1Kll/DizN7RhhUAG8ekaN/AnVMRB63zzlRHygadCVy7tlI4
+zpe/orYXgvRsQl3fhiw8QfFXFEGA44Hcnq/K2KNdrFc+Kn/c2dMZfpIbJNS8bzC
Nr/ZuoBxfeKS3MtdeM0N81VYXMpgttm6Lvz7zQTYcm2/EiZUdkh72aqVjE14aJYd
Gi3rvwx4+qMNRfb9GXEG3/fgE+Nq4z47WI3NtMZY/qhAPhfCKf4bHNezbG7NSTd0
Av/VF7G5539lkokYNIILkutSaCEaOTdBLIRqZD+OPPZAmXk4rCBZmwUhwi9I7Rd1
wPHZffyCGY0GIozUHpAaeu/8R/XxKrOxfsyTDHWDbmGyi7vJcvPdDqUNvGDIpCH2
Jrh4mLnXhOc13TAZPCt2Jmn0ZduKXXmzSkaQi1UqX+M36kqDtwJ6mlR2BRHvVkcd
XqNKXgGAnjpNeyeGQ5bv8XW/m/LJS5s2Ku/wMJ+cilx/Jpa9s/qLG1DlBa5SoLZK
fQVVegveB3Grh8WxWCUqwoVfWFpvAd9MMBwntnQCso8hO6ZSPVhCn7voM0y1nqzb
z37gjsP3cpBx8lQVpL/CsA5lUXU3Fl7WDXr2d08ma+G251KK56EgMB9B5Njqv9G+
70aEnzShIyp7aaofcRbiynwXj0pHpQ0ki+1WNnb/o/4yEcygbE+c51fWXXJPeQlW
S5tMxNll62NWUD3CH28QL4PM8rcech46gKymTiP/7/BJTwXo7LWt8S82U1KMAq8u
8WoGkjZRI69DUdDhGmEhuIS7CaUztpde9vgoQbhXxLlLhN0fKGDQiWdBft6vdOGX
asP6U76lUBsxcIyXRsTavGL/g44PMWGrx6W665zq7UWBZAzWyo0Qt+5GFuqNYGm/
nDZfu1yyIx5MzNFU/1LJ97WizV0c4llXQ8jZZbGIXe5loQBJolC9mWRRfLzm72uY
SskomQxaJfLB/V8HkpKs3RUvSL+z9gx5b7czNcOTeQWiEnvXf4xlvDoerJqFMxAe
OpRM/vtTFCvDPa5aIjeE+vL+8ah8caF6UNoo5zLL8a7CaN54571+cax2JtsU0iAT
elwIyv9KaNl5Fyd8wR8YmAxF8eLC3lhPV8wedzWo3bhS2C0hcbAWke/rTl7nvHbn
JBP7dYBgBYtxP9LFsRnj7xE3NiDpBM2/HUNm3rsbRJBx3rtuYsIa0V945X8shYjb
IXjBHStvufzS5tL8KpZzJ9bYlVJCIo2B3A0T2cIfGVqNQ0HOYrghfPkyVD8cwIos
gBVkXnky4qt3exPU31ttID4VunGL3HnYH2+6QaYFMTYDZsyMuDJUGkoeHoA/3hnu
jQHDZGsS68GB4R8VpTgt7EvOck4svRKHgAsWQ+F004uSJP/dk7a8NzrjVCLzvn4n
NSN+iNvWE0Hr1vUWJ+1YMMxs0M2QCU0Cu9d0t/xFLd83Y9MXBZByYStwdAzq+J56
EdbMrZKhheDr+1NTUrL3O+z2CYq6x+0FR8FYPySNpgdQyBjI5gzOArdLD7tvjy69
7TkEWRvbQq5VLvuFC/lrxWLDb9LScaD+HIj4scWRlIMT2mVDaOoq070yLIOqE1kw
9eNelU+XoPgdWZdiQ9r6RZe1DDxVSN3t8prFPCsKXx4RzZQYgxzNXS7vsWk6rzmR
4ABDXvxDcH1wdj7maS4ln2Jvsk25G6hu/ccUSDgS74oX9/4aM1WPjNfHnHaVNueJ
gRByt1DkHx4wLrVcrb0DZX4t6I4JfUL+Y13E9V+xWC79EasBIldQCLvGu7pN97yB
UEJmBzYzwfeLA8XzEfdpAC2hS2Ld4/LKcjnhUu1ZRBIGtc4dyHUh6++AaDi6lel/
yRUbHnNk1Wf/TtBhOEGIUFoZDKtur9vYvA2kmq8mCJRMh4A8CeJlPNqOeIKuSjh+
dAXnivzcU3u3d60sTcndiNVeStprGyItWed9gao31JdWD6OzPExGwT6W+c3qOg+a
YQiYLdXGTFpeUMDhs/RAGXlQTv7lMIW03lmluXDeyear6hz/y/97gzajYJdhixks
cqcIVqLBG1Z9fcoKVLjSvtboeSnCkUQcwP6BOeaSGFOF8LlpraePVMvAofl2Lp3t
IhKfnyM6VRlcy35E5hc/2j4Yvnl30NXYFKiq1VlgB7SplKKFkxeP98LINtjd5v/k
PP0kPdtXx24EIjEWWz6G+UmqCnTAxkxJoj5YudzNgfIabdoytM1Yl7hQDeJ+qCvB
PNrdv1m/RhaAsFGGzmmMd/3QhdBDw2mU+JCIZg4s4ReltriH9xzPNQfXmGA34rfF
dsGBMbn7Gp724YlTbnd2ZpgT9ovsnkx9c7+UB4pskAKzACL2sFq2bf/symYrhm38
/BI7kFUlbJRFoVt12Oh77JKdC+JFwtdBX+b02rYwttEuox05Ku/ssVNvOuNyoDSX
fRJAdsBWTdTB1CPuZQ8Vt2vVqGRBwM1kevs8jNDjf+y4cNvI87vJP83q1glvKa3P
BabAzYKqy/NuSnp4Ii2zroe4cpLi1gC+U6F7/9se66cLVLaH3YKEcZglgmyvFsSj
40hRUzPzI40xThejWfvVS582KSwFxSQrCxUrNJP8QUq9OmaBQD8eD4gckf2y+el6
O12G2kwyWPxKSZRZAzOFEZo6AyXY6zt9QchEKCFGHNClHEVebO+mPN7fMLlAa/hT
DJkCZbHD2YR/YaxNauCHHFhho5s8KpHKa+7XsC6CYCr/RPx1ZlqmR4ud8g6O0PJi
2/gTXzMcV6w6DUgjD6Ad3Yth0U3+D/KwFL7Dwg526LFyvugl3ElVg/H3xJQYz9lq
8+fIz4b1iZnaM2kj51YBBCO2BHhx4MaxkM1sEM8LxtcYCqSNN7/nc9N6cMn/wHPD
X94J4KFKs0ysLGusp5OMwcZPHuCHNnmwK7QH1gyt2VeNU1Mq3A9YsLT49nzEm3ew
FOWCvm2/FE+WsIaS53ovPM/M/bsOAArj6sI1/IJiBFLuIdvySPOD7mCSmEN8EYiQ
KeY4E7N9UwZh7oH6OhEWzxyEDvifZNE4hiKY6qtq/iGmmuK9wNAXg+KvyYjisjaK
mEjIJSsPyliXwpdZDbYkngJrlJOMUs44b9xgKVP4dHCjYBGC3dufwrBGD8NgiI5V
zJItpwFlvDKjrx5bEj2tVFVMAIfC0JCLrpLoQtDRr2iKVibxMB3B+MvoB7UjYjXu
Vq29wvqzrkwsFkxg8dGhgRxqEDloMZhHSBp0KElSLq2bOe+HvivQtXJXIv7F03av
lTWRcd1N4QLNuWdDfeMUSNrJWZiasIgrJV5QrpmC87G7949ejkuJpK9VCU/1d1rj
maGl0vlVrcGnBQSSydZtGz12CmwBXOTzlls8WnxcxtqU0JOGfO2xWX9gfYVYwn4n
1AC8eyR2xANTpcIvv07QCfaeMlegANaoxwzjtWkosVMu+K75bnYIjot1lONVjM45
KjBFNAgImsEhk9wBGgHWLfEHgd6JM6MzKDnCw39ElTnfVCpZGMmO+c+kXWy8pdjA
h60+E+r4rfOIanOEObq99klTWSm1iJfPZt/M6Cm2noRewp9mcrUt5IJ54OxzJ3Kh
fT7mgWH2XnS20AeW6gwo99aIZOG20xota6xB6+UNvbLzvM+OFoRTMO80307EsphM
W509Ytz6GxBQtsUuDzNrfBscXIPJt75iIPQWT+ntsUL+TdneGEH0Ycd7WRde+frv
cnoocfv3Q+NOKXpPZ4cbSuxg+fU458qwsjjUfQXpaUj4WUYzPoWty+n5Y4RabPDr
HxhyRFkzMfT1I18G3jOJCpveVSD63itKYNTcyD9hd9c11SYVk2pSQrxyDZw3fbeB
HslMek+ZR586d0vcIsZPPaq/tkPT+h5obuOOXM+j9H0CLue0fF1xMt9+eGhIFeO5
PAPEq8y2Kglb/8V2/jB+spQxY105MIMnGSVQlYq6IenGKOw019mXpFWrD7VUghDD
plmIUbW74tGBkJQ4oPnP829yE3zGmzYgnpODCn7U3/IybkbNonziyDmagn6/iTsm
jGoKRzR+u9qxiuqrm+fjmnh29b0ApsV241Vxdt+eAiYjHeEbe81WgDKzF9phUq4j
tIjyK0FBDI1+I/v24b0BHtkYpVa086rb2r/XzoaCmHI2IGk7kISU1GyZdIbf9677
Xa9g2JQ5QMJn6zfjWHJyrowrV2o26bsXevjYns/dHT1kZfBZB20Um2TUEHav+f3W
NCn4Erf2N7ClfDlA869Mc09GCYisJ2AfUZdfYWGeyh24PN7UjfaHQlmmocjAQ9Ye
MJXWL+ooCWrnxtwTNaP2oXuRMTDYoKP1axCHxVU3e7601CJacK1b5bx6HdEvMmnV
hCOFv7nxV17xPnIfz7z72Wsc2ClNHuX4iT7YaN946zP37rJc04QhdBisYApKzaqd
USYwu86ykfNey09zsGCLzr9OVzsr3VwS056RNBSHqE73ooIlhjbOv6VFtcDZwIXo
API9fiC5cBmIGQxSGVbfPnSL4Aj68uMfC9gfGma7r00x6JkNPDKJ1equH5FWdVlC
TSSQmtQKFG9l5DNz/nWHNCdFsjmxrgV/iAAEyKODOCv6MFKyLQ7ZVLRhpBEkIZm0
ooK1pZF7VMGS3cvHGTB2l/4oKYQeUB50cPDNK9l9BZcmWYdW76Z2c+WpRiUzIB/w
7E2n5z/92MPs5WVPsjUEPeICbA4HRhpsfC2CavG9/Po4FLTXRgyenSDwNb+YHp9d
GQO1oJr2Q6d656LpBILlPN8tmeQL9s8qOqGtB+2QORALOO+UTJ0tCc7fyZrKBX6V
x03qSTrVhF7qrJ39//+wGAFK3+D8UX3fcVJ4+nEyBKWAKwggTmaTWQEXPovKPYiO
kOI4RVuOCwEUfu08frF1brypyGCDssehTuq31/UNhrMAO4DwvyOmYEYcdbQxopu9
Bqa++YQHq1lOLJ4adZkbMMb25fquUrd+KEKtKxf5u9wVPacKHhrRFXlv1JIEsk9B
cNS6aaOeOedu/20eSG394+rwd9dRMzmMGrNifWD4CBIFfmNGyxWIuCSDew8TXl7C
NO0ZzOZQqOJapeY1EwMkYvVgYPuLJn/ADWgQs+9xLlIoEMjraSg3Fw9QR6wWN/do
08GAHj97kOxPG8whZr9yps2DLKSWOA/TcvV5b3NeGfVPbc3awu5rDo+/cs2w5gw9
BbOT5syM7yO4ANNGlUeO9Q6466NGks6egzC1CnqMK9JQDExlVhe2DAC75ydEM1x7
yyAGcoI9uVvqWXJd7e1PR2eVWJ6HmyX/tiPSeWG8pZyh3laY8XvsPT+haFtrwD9g
SAzbp6mh1eJUSv9WxXpWNQY4YkLefkOYJ2yoO/2UbzZqxgGnTjI7y+8LCuynorzA
QSrB2sdktRbhgmumHGKkeLFR7kfvK7Fm76XAiZJSUvkWf4kY+ObHbiZ8Z3I1/fhr
BH26ROl0vOH2kPvdtJfvV/iwvs5yfbs1vnWE06ndOpDUL9hWszSjgz96aL2BYZsw
YmaEhfys5CPRCEs15ZUzvQoKfn1kx8xrZMeoZK9bpYf4PlcrJ/ieAxme0hL8uSps
6UBk8CkHpLqKpycWd6I4rbvsgghBX6qrXrCU1YQhouqmojXCVKPcMIKUQZgGGWwY
KcYsg8B4mmsTUYuycl8pK/80i2p6nbqACFlrr9Fwaw2+Bxp9HUiOBFsjLc00BCvk
8oQeTw5Chtavm6RKJA5mwU0oAAkSzck2L1KbyNJqOsZEynXSctK6ZkjZ7aOxbf5O
k7LkzdSd1l1wr0tRV16Gza7BbDqDHxAErNxZ+rkJbDXJLnKoahqrO871hiwkKtxw
Me4ztju0lrD0lRtt+B49YYAX6qR6CfB8CULsVgpylLggLjGi3uhvtDOuPfrtOOp9
Ejs07U+Iom+DPY5YDTjYuC6q0Cq+FpJjqekYh9FEyH9NS1uBl1+5ZJwxd49nvuTQ
9HCPwLNsRiOLh1+1q8O28P5KRLiZr8wPVSGZaIsvL37fkket0Q8ryarfJP6ld1dD
OVVspqDAmyE0rW7MoG5XUZcxCWyYh7EuHhlhSD7TPANyA5YA6fVvBjScb3JqCBNz
S/0jRYde6WLin2h9ZgLxOPu/xqnJQ93XPqIkvkCsdStWU8Zgiv5IBS57IiT5oVP7
djcwXfkz1GEeHnQFCb2its+ipzK+GLunEBE9YSnhcqKBXhGTs/2cOKlMdZ3tlOTn
vDLmNjC6DGxzmciOoQif7jCbESZIFqT0Eu7Jx2ySm8dhV1elP8cpJB8Jx/QI14CW
/YN1i02RIHDExCnRyzwpWC2pFkXPkTgnjx49DcHRPLnv7sCgGQpVxFYGOsjs1XSX
EfZbYt/+LCKlnLOimSoMtNpj6+I0Xv9FPaVh4LnqaTpde9N2xMf/IbWWhgy2lDZv
hY83UpXRznSoceuHKvmac4ym6SR550ddgQAeCC5fuaOZpd+qLcMOd3+3p1dwQ4x6
PtT7kldwXZ5r5X+YIoA4kwTU/Ydg1Ztcqj88qXruYcFa1D6bvBqaz0XkxOzvgB1G
T8Tj1t1oRHsuouNV7oWVoMJBAbqD9JXkd38qb0I1zwDEMsRS+xFGqQwrKhKgFFcZ
isjVf96Iwggm6OVl/zBgVCVx2vWXvT/av+9CX/ZYPrJAVx9wYvlnY2jICpbBRyqz
LSeaeo+M7V7ds5xXi4oiuE9dmXjxD5w33tVy7B0wv69sZ54AnQOFpaS2sZJ7zKwZ
mn4Dja8YdeJBbbq8Z1TrF5K8PInDU4tJBc/CEnawuzBQVH5bjkB8fI2cc1R97d96
SwCV+UwH33/qkQTNpjy5zPB/NDDVOWFuO3mC8u3twJc6TebTDF1kezBUvtmwDUtb
WK7bhk/OqnT5oh3FoQRMotqWWhkFid4uxtxZ/bwH+2dCG+ab7z1GKR1CwsQ6JCCZ
Yf27x7tqW0psREwrwi2R9Uixa/JJttZY2VsPPeeMZjymQBO3kZfRg2mhtqKAazXk
NXdj7ZVYw6eh0ktutBdNBz/anNRr/KejHHbstkrA/VsSVK3OqUu7Z2kepg8MNDIj
5dIuiqFs8v8RUBMsGaFT9Mxf6b0ebOAV/CYZejsPfUbtP6/Q1SG0mr8udA5TuIEG
aRSdxZIV+8SznMq9bFEqPqF7gaPH6LMGLZvLx0gLk4jYvFhpCZAXl/qbB8sj9UTL
QZ9D5mL81w67sAXf9sR2Nkd796tMTaB62/u8czjsM5qDKx+jgTq4BQ5FdMSq7eTE
6n+YPyUYa54QgL4xoxv9xflskLa/jqLU1k/GtLQPyxiHpkUouCqlhkg8P8QMFyWz
aRQWD66rnHS0VJQPgK1k+q0PTt5aGpOdgPg6E52e5oFf+YU1+uAc1K9e+qvs3WV9
k4BCLEl5f0sc6uUgjaHDIyJTB1M/jwqHTgoBm64fqg+uZhCDMKGioN9tVeaP6FdP
z6vOlb14TIPOeGhS9ZIKXGsCEPJV5Zh2aq1XdMoWDScHtWkSKh8DCYLZyBqytUpY
dUfwzjHJqskqt4jbPxjq9g3lG72uTifYe54388RWQpIQ3z54MqICTk3jw3n05ALJ
64RU5rWD/nQaBqmEPTegnWyWkSy1SL3/TQ+sY5wyOmaKc/1LlNuwhpC0JJi6iqG3
4coG5ZRcHFZjBftBrQHdk8RiojRks444lMV2dj6zl2UPOjkbOYNSbEO9Lh1Xu6VH
xtivrHoTLkYhAOKVajpAeeN7gcudz/Hl3lCSZ5+rv5YOICKskhdVjzW7XIcHIooS
OUiIzkHdJRtETVTaDtDMuv9p8YScB2ltyLq8/dVUcyYAVj8F9Fdatv2qR82lDayk
6PmtTrA1rvBE/JxZlOfhMGsgYrID1hCuVt/eeHABTsASHGkX3MctcGN2A9An0d1H
NsZh6SICZNOGrnzxiO/si4u3exaRPcNK9ggkDh+lARSbSargt6PjCoBbeHVms4pb
APShjMQqV3pT9YfLNTi6LkoBxa4rAk28kgXIAkMozhC7Zgjqsso7XuM+y1J5fIQr
dezZsbxDsvV59OfRJPI5JwW/ljyIneEOrTVlK6cnvDGW8fovJ1GxvRRT4jecVS4s
AES6bRgLbjylyypduguQL7iFiGl1W1ARVeD1Wm9qhnWzb7KD9ne7RkDS1L3J1Cv3
FAPIkmbi5kUk3J2j9NevLw/njDXhr1B/191G4snjaNuKf/bnrN+0+28uxVRteS0t
LdAhs3tyAkaY36owjkoV/N0UgjD8Upqmd9e8/0Wt7rN5wF7iGN4NZw983Fqu1G4U
eEtD8aAp3d8fxC3kD1q309zAR1HFf2LSBhDMIpW8PM4RBIEySTW//Oy8sB6jHip0
0QY+6Y6EBUkVHjGshm0se3HLbf+bhYRhYIWsiVLvHR+CAhyYOT9lFre7MEw7kZPZ
Da5YP4YKZCryS5iO8PLCJ/MYt1uDiThYJHGfZ/nzEEA6JlpJ2D5Zm2v3pA8B+j1l
PcftvAK07KDAO3ns5WrMBQR/UM/9rdnF3+Wjg1i37ei+XyB+HSUpktKjUr50/tIo
boe2cCL+MmiO5cKLn4trAanLe/wIWX5nDmHt+3DSBa3YUuw2Y6FRv4YNGTWeMJmQ
RRtAhCtwnfByRJ6sWDHLe2e48A6H64k87HFCw1aOAw2+krvGBFPI7fRDS30TmRvg
K38LR8XmA2F03KQtSxG5TIgJZevER525flErderwwerQiA8mMRGZ8IIANLbP4H+s
KEV1YJMZUL1Zv4ErxtIx4q+RQ4oZ/Mt4qW37Dy2WPJySehCVBlT0OhsHgQI9UWCR
tzD/uLRE7M3y2OFi+jtha6fxpC5G0fBKf67+QXf7eIWCZgjNwRwhoJUocCAx5yJk
tet559iKjfOQkmbcMbsAs/iXogjsQ/TS8CB8R9lrFE9R7pefbBkJtcVZyny7uJeZ
FdKxiZb00spaQ2DciSmFsMCiO0aC4PsgxYiAz7j5ge+rj3YsTCQo/98ltz98N02l
qbpDW1m++JpKmG1ooDeuXZBMJRkwc2r4HM58eotq3hgOcZUUXvWfIh6a3NI7hsqa
0zbuCiQ/WTGVxIYXjgBNNv5TaKIxzmW/as2qbDLZUChNOQFIoKlee90QoM2hLHG1
EnTYXxx+53jy5MYgzRsxVlmUwzE8+d0Pm6z0+XNHqqDoyirUSGRLIdaTDjNZ/vVW
ojlMWf/fqtdlPp+pniQFQWvQIL94IixQniXrR1Q/A//SSpQbbiWA7u20jBGppvLS
l8h1+nFDqX9i+crFg4AjkR/aGcRtk0k8gjWz2Llnz9wFAS6391DLQxBNQGkxNXl5
AcmMLz2UojzrQv65acHa7RazuH+kvjp4mLvG0yR4C6IGC+2ss+5qMvtdndZXSIEb
K3NpzTaxdEL80+96ra0qkOve8trp6vIkcxRewp5dXXb/9biyPQdb6WfAu61BeqQZ
9+UZDT52iRj+PDkYr7uQTxgKwFr08gcYQnsAWTwxkNYAU7c10nMwk8SFAW9DwP0l
1TQQMDYlRdbMD/QbE62NszD2wV9mx+3VjuEUSPDEX6v3gahkJ3WhzY3jmO7G9v1O
E8kiwIoyevUy1gpuOUu2whzKOptqqNvgamR3LFwRBkyMdoD7A2beCfs0d7UnWFlm
4C9emnGfPACKOUtJxDIopg+d20kLsz64XY6xhPYMSMy1b+bf12+MHs9pBVokYWbM
vq2nfn7V7PM0rhc0bRFqS0DOmuHU6rrvnj2paSl33D3y67abOmiZnO9rgdW9aqDV
Rdk4oZ6SuvZ5cyBL/psEZ6LShN0i76qiKNvkEfoyKk/lOP7CJ0stkZhRA9FK9llo
ybRAn+yVdg7aNt/rnl7OtGRcVWy1nP6folHFh7F1Zqt6fPitd4jxhSaaipoNclNS
2T4+9Rfsdwogp/wjqm9+3iQiHtJmTtQE+Qpfew88EKkALVmprPKd8r1urEUVQp1f
nHcQP7fUbwBpF4dL47MZiLk8NIFUqnLJsJegaTB4kEB+xn5u92QPC770tsaDRbEO
nQS37gPn/ArsGxxSFZdr2GTbu8jZNewh5WtYE2TDYBmPA1bsAqhsq1zZoyxy+3yW
rxUD+to96mALRww96O6MGtCrYyP512K3OHe0dNk8hiQ6O8I+bI0QfAjodeMhQ2hg
77wQJiPJZe/5Xmm6f2nhmHpZRiXQ0J1QeMjIEDtGOOyPij06RvC35BTqJmYBhaqV
GaB7sMsmNYRtgmHBkyiLnOqNZSiZPqi1CZg6FyqoiBREjAC4XNkIoy+/Iw0v1M1v
lK6Jg9ki9XTlJ8+LjrVdZNmwAaGD9SJce4P6XcSQ27nTGOiNjf7yGWII8lbEdjvV
ULC/w1hKvivrZW7adRMERidcaBG1T9RQvfDjQLuTggNDzdqymcCtYTB+D0E135lq
Ec+1VkDeld6yls3RffMc/QFnxNTu8HcQsCJeV3C0w2OFOPG1Sv0rNubW/6ZbRJSZ
MHWNOdBax1pM1kjnZ5f9GNi1LRIZGfSPmVG85i/64IdvMOpMonchy8nOicCAqpq3
NL7GMU0f5Datud/Hi+UAqNvZ00ndV8k7HtN0LI6XkcWdNc7L2Biuv2Ks3398oF8s
yWN37BZZ3Y/CdwbJN+TyrtEhCEdkzAFZyE5bb/Osc3vd8xcUw9ISkTPlPYvVUEbA
sTM/mcZI1DNzjZGRih8Wbo/h+N0tnK5skmMeh08k1pSHFAa2ELEAmQ0RXGnXDNqL
/JhSlJ5QEnNOGskUhnIi8DtMCnVRhcug1tE7lkqbG6+xvHD+ARiolLFwHKTH3YfO
tYlicLvLMVtjOeHxOWdkXVAavTBm/rl5bfenhzT3D6vv89oYrcZRK0epT4myXb90
aBnYJVeJXqX+zJlNAbGIjp7etqtUmwqMKmyhXs84JyBwiLFhBCOiJM7QSu3TYGLt
KVyw3Qt0WGTp7oQo8N30mzMVqK8LgQIOa1dYUT96HdGj6GcGRudSwUvhieY4g2dw
O13jUFr3XKDJMVexC1WKw4EoCoVCIAImXj+lpCxRZ49MbFQJwa91q4U03S7nqUiZ
uc4Mq8dBcQ7SlebMpBayFoQFu2z7uFMK+NnQKU9NybV5uhnfnkeFrxeiS+O3Nv2Q
1V57xbPYYG95HmsdnDJPATRd2T1DOZxy0gOWVpJ+kRSeXvRdltG/yebz5exk+fZs
bcCWcTxSoQTBHe7WvyN/eSuDvbVeJc9C96X63PEGcWYFofw0PG/imGz2FC7AMkK6
FEdOF1rJ5efmKZdgqHYEqqbqupnG0nq8Kra+Wkat8XdD6EsbGzguCCh2OT5SLvQy
tDq7lxRwNtNY8ifuuYNil7YPqfrU7LFoTaIZvnTgUGPJhfCT5Z1MiJZKKy7+5Bo7
mXKzXt0P9nSVgiVfzrFNTOVvcZbwl9SA0jXzn//v0JYY3otkPSm7OV5VhTPlCwN7
ioO84hraaw5O/DTOiuadBvhS2C+HxwaEiaqTvwezPaSrx0/5jKGUpCH3sDj2vIju
LXmtIxCMFz1AkZd57IDkS4NxSdTYkbI6tWe83MrcjaqtH7TNGFULp1Hf2RMcLEFk
9HfWn5TKjJUhxYfXATQyZCboLEZof0KMMjC+wAs7hDS8Kj2D3NRK6plTywUuzcLJ
FKWqK/5PXxZKmVA2Z48yDGRNajHIeMIqPn+wgZOzSjeQ8R2eecL3Z+0iUlcvY0xa
Fi9AyovDgm4RyGZM6DmyZcDEeb78v9ulP7Kr4O6LTUg2UZbHCsDeIkh5RM3buRcw
Qo1nDMBVaDiG/58z8yCrd1lFFvi41PdvlPlbc+OF+B76iYlOqeCXTllLARR+thWo
YmrY86xsw2byvSqJb/5c6pvgjMFFd0cZB5AJkXj6/iPcZ3TLVXudsLlQjiss1Pjv
Hq1pTjxJ2cg7yBljNrZG1rlXozsGuRYYmIdzjJB9kib2+i4ORAC2M/tH6clrrkvR
NiLd1zuhhT3CuNj+3NH3WfLs97K9IYvMlkWV4TzR8433rA2b35H5c21hhOsqM8Ce
UiinC0tXPMzS5ymqviWudeuh2AZZZuo+GOez64D+agdPD5Enx9qaVvRRuBGcIqlo
i2jKQOqZFz+IeHzUlfnhbQqm8t+zmRObbGpQxJMtK1lWHBCDpdm2yjDpXKJiQ2ms
mh8cJ/tiO4up5LAgEH6tTU73ns9Fbpfc3f6BIaT2riRW/7WHYw6JO5eDu1xYusa4
L7/1wIfDFA8hRRT5E47DnhEv6cbtFcJXSSEG73hskTn/KUY56uXDmakuoFz5RS9g
vNCAMq98bX/M8KIkPbsb8LFMY0lasOWPVqthHk2JI+lzmvtSZMDCLyMg4dbPIDHY
GrD4/2zAvRPoJxAEenI6QM0ydu69m3WxKlde/BbPkMajZkRC+yFILJjK64XwgsS1
7a0Y2f+en9zk9kZDIPw5dI8l+85TM8/iq4G9/GyAqiuOL5kQwaoZfJgnn8kt42vm
AbrsX+6IGxiKAq0kwqjKqnak3F5kR23WVxv28Uh/6Vdfmu53t9oRU7gvd27wdzTc
nqHngQMrJm+gKM/mpc6nDURGXwgfcuyJuGyhgTaA7j5ZqVvTOTWLZ8dWeH/kXevR
9CQKS6MxkA2CTIMJDPHGZta/Ov6NQoK7Iqoxf7nE7jf87zs4e4+zGlRAPm1hcfUD
tAHTHWeBkncPs9rBAH54ioFDFWdKlABO8hikHtHpASJ61BAuqdQV+pZhGEjt5MzP
NSQ95sp0T77FNPt5SHE4HimZ4nbwvdIpq6KhqHFuCGu2bkaK2y8Pa6ufnMC8VZhY
HNk+RLV7QzMUpHs0IvvJmmVthaK/sccrSM4S25zihdQbxvfOk2nMnz4+xkljmDTj
IpC2b3ZklD4/UPa/FZ4Cjggk8bSQiuVJocr+sIFyS+Bl0eRc7ykix91dugzyFqxw
629tWw3o21+Qk7nMAqVQNCi1MESq5qmjfhcVHkV3c2LYBdWs8MwamsxppLKp8Jpv
XsT0s/G+rzFU+TBiljhQ6/ZoMxN0fVL2hKge2ZLzhrMN/V10gnDAGNLOVX5PAVj/
LzKx+dmcie2vVF94dqTGfAnEpBqxG7w8w+Lz5Ugj9fKH311dxxeouou8k1osk29d
PreIiSswJdPJU+xDSSB9nyq16GtWdMpm46zGglh3+dN6vZo9QX+v4IDSgITsghjJ
i8+bRbau/ul0DDkB7s+HL+L9+l9d07cndHhkNdLjrpxutB3t7e8D6ywiknNS8HK7
zeto4NyonruOQKDd2cnJPYvWr+YvT72H4X0l1BKoSNStUN9SGUprncZ9ZEmT+AJj
yrLq+cDnSyz3elXy935ESON3t6ZblNPNnQrynkgfZqVMtLJ8Vxs4QypVYiIaEC6h
EH68yJwm508U7jdfuU2HQlq7pEosWS62dz8JZUOf1Gsh/7G6zVLCQZizcv066ZrB
F+y26KflZpjHfhckNHfUi7ItguO5dyKWcOrqUNwjYLcru05/VUrdzY3bPhI8bmKZ
egt2Chygic0nNbQvo2F3wPHtXibbhiCIO/FVdwuMcYWlctTH7NabXEzTLD0D0aPX
irk3SLSUXyaR9cAf9c2dGgzbTL+gCvK1wr2/dkPWgAtwP5pRzRfRKIsva1md9T1n
hs//xxwdJ/zZEodEmgb/eYUxIGk7X5u7DydiFabhn7Ly/UPfHtCstc/1KekwLXUL
xS4JBuH/n6RWaWWlF2wV/xFerV9/CwVIBF/HLoGp8HHmU2lqovtFzMi/PnqaPxNG
3Lx755pd8lwt3YkIyANm2MBoqlDXW2zbgxwdaPLBZT8/M346C217U5wecMD0MPZ1
rw8L0zVK1IKMZQ2WvRoMcTPsjfZaiWVWt/8+wQSuz0+L5S+cfxT1DN8UzaMNhj1Y
U/m0gWuF2SBapDULAMjey9MIINAc64Vl3U3PSJcZ6H0MEI9ypgwza0e8WzpORDwl
n2zUD6u0sNgzTOIRRtYkssyZf5FsG/cxUQnr45ezCLPlrNiA2uEYGeZa5TP08cem
WLUctt9ddbJZOUtUGsFTdBEpir3Pb6zpQ27yS3fH39wWj9sVBNhyo0705kaU/Zo3
H+2iNMuViywp882gm/oFksGxEoXluuSZYFdSikfKh+KznbiL6Feg4GifHQwtJ4B6
5auEjnT0f458yoW3iZQCYzOfPfVfeHawCPFvKOvIAGzKgo0SYdR1XB2yurj1jXsK
6vFHjUkjQiFLL6PH7vNKl8yaPCmzoaBR8Nck4shekA+7JnUhu+fZFPuwVo2GLBlO
0vsF84ebC+J2X41dmuk6Z3P2WhOQSM2E7WA6UWD3KwVUVbd4WGjdW7f+eqLUasT6
RZZ6GLxV4JfrroLHWQhs10eAJ3tMUtem8X9bqcPtS8Zo8atN9pCmltsyliqVIhCk
tCUa16WLQ2jDREX7lmn+E/ELNYdBGMZJO5cbuSrtJFocNp4nNObHiy9DwwKPpWC/
P7FsIequI3/TON95D8Qcv6cRmML4HYRtY3ArwQmCqevdjNIhTBYUM0FjFmqkmKtP
5icbqFUmCw+KeftalZIqZmF53KzGF3iUJp6kGCGmynaN6AZNawXi67RqImRU15Zj
RV51hI3NpvX0S1924dKs15hB9aT07Sqc8v+pEQ7HT07Weedgs04kkkJLCD0Ou6fb
GdzgQXXwti0x14bRcRvU4g3UhJNHBGC3UN57gQewL9ZNyKn3QpP5RSOlq3YxEYIo
BSJ1vUhQ+M2YGoH6ZyAOAnnfcGOCkLPaWvqr0N6oiwLoTVUvbRlDhVQ0gJt4iyeF
z0YeuQdQ4zKF3IdU/IxzIuhFi0btXYCUZp5HCKv1DDhevnssJIzxUadNPlYdstxy
Qdvqq1S74V28f74mFnJd9YeNthkrJqZY4vORBEAX8KmH++xioGTQARSBZgPOXHm9
gWZUDjPrCTrDA+IYjeC5kSBiD+YuyQaqrMoSE1wNDHbywH2kzx39thdwfdRo3kwB
ucp9XKohocii9onZSAugosSnsrg5s8EOLuuwjU4uBwXTGNLve2mr8/k9KiB9qmPA
9vZNPFIpHqfD7hzzIQW0O3mqE1MxjL8k/6/NGAZiunz807H2GcXyJxRIRIJCY8hb
cFZ6iqqJXoWOGXQcwIUlbDYoD0Jn+g5NSegjhA2G3Gx5H8ehwu2ZMx15eyCKog8P
34OSXiYxW8f7xmstMSQFs+vBjcd40gby/2nT5H0hKhyoIpRvKahRez8NL5KDPNLu
d7k4580mfpEi6A7C4zKHel3ItqK0HDcmKqn1tw5DsLu/ZLhS9z4z1xfBgv4NakHt
7uP/9aFYKnMbsKBj2kMkV0De4o7vFIGqA9Uzo9K2tf/J/9ltSbMyODfCVq/Mm3eh
nY31rHHY6p+JjyLYG90ESsZEcqHPhceY4wu0xa8W7pGVCrfc7rnk+5leBOl1lUkp
qsIj15zeivifHhfl0I2KHW2L60Oi7fVm4HaWK+CXqE5LbNQYbhnLMdBDPAi+L2jH
kfPhi9Ov+WaDo8tyg8R/uhINvTsR99ufLVBLJNGe4fAuC9TtaRrzC/GlT12qhDWG
p49F4aI0wAGEJdp9v/0aEJdCsZzsl/S2NnqBJ+tiRYwuLrmZASL0AUZGYEJkLu9j
+5fCbOBLKTDdVwN2K8nwdXYiHUHcZBEIXJvUTcNhqyM+4KRIyhM+675LpHlgNx8V
n/UAOrh8/2qZGXbyl/6BKEJ61ymptQqrQuQaD3Z4WZ6fN7vQGtoS3XZGFcqMLLep
y6Tpx7RhdUdR5tcuwQASSX5OoYDUi+k9TExS800gzj/MacMmU6CfnQoEgguXLZGz
sSoIZBDEhRTMpjTtRPmbXG7lrttGQOeBMQKmJY5DHyySlXv2c0VPehLm0B61JdTj
27aVnjlVP39LtbtgtJ78gK/sDQLI+2gTszD9yJq9rGmWvX+CPS4pWmFC2wBFALLb
yxSwEYWeLpG/FL8zRnYwzHB7atkO3VCXcKt4ggQ1iwuD4tIwAtFcKiIu5SGbgvh+
FaM5REx9Op4dPU4THEUIcRE2yBWqcaBnbj4wMBSNKwkKR+6jKFGGeSnxrMAZ5ntw
rBmJ1ILzDqsEKN19sU7rhL6I7DJakn6Cgzklf8SVU11w/JN0HTprSsCDul+ryjE8
/t7ZWVzStcvRtQEoGAJjyPTC8Zfyjw2Q2Ga7ZSb7JvxAtgM+BVdD/uvVZ0oXxnkq
AeGGLbbcQAO4+4ej7K6NNDnpdLGJ/lb7rBbTQjd6DGR96MoXUZEc2F7yXicCA9FZ
bPkbcwRbzMdY/TMZpagSJpLy/mKuuYA50BhCgJskgcdkwSBLzsHbGcjgv5gD3JGi
6pbnQ0jr5dOxWT+BhZA7RIqgl3Bg31mSKpRxDBlv+FItvPSpokQEPnQiA0VjZgMv
aXZnnxrk5JJV4LrHdICnm/c4bNiUfM+8UULg9EhxJ7ZpOFruF04efupcFbJ0SO44
85OXBl+bMrB0UU2MDYB+eC9l6t5e+IwZN9MHAxmMRzgvmbJLu1hVRTOUUKlC8cym
Nk68vVzmR6TODm0xYrmoUT4J4sbV21+TVx1NMJVGEP9cQIPIWKoQQMjeJI2btb4L
w06fTFB8cZgNw6QnvzjQTzPA8p1PAtYIOmha7rcwjvq667Kvn0OJ1SUe2LwHxKJl
+baxRU4WcOcCeCqUvsPGGRnlPx6QSuWUy5OzOd/TZn0o8bIK9RUyRttlc4UsburF
tQ+Cv52iQML3eOp7fYPJWXANS8TTnMRlVFEiAbnShMGiIKOPLjhInx4YNUpZS4iY
jrALMWANpwhFqJ4gSbyi+ppibsruocilDw4e8E2Ep+ME2vQg47MXxyQJ+MLEn1aQ
+dM4/ZvCMj5XGhGPnbTp+uYXRoUHPAGfDYF7fFWR6cCojaPQPsLaiMH7RYUitCOT
ryU2ilaa7WAJBbxVzwvDI5mhmfcLtdHrySjke9vwxJHj/c2qaZn/aSJM4ZMiD/nC
qPTOPvi6fpLCN2LKqMvyXinjus3TRmXPiCtze7Kjlg7DHDqakcGVQqr8lpYncRFc
tM8IaqpQ51Tm6ymqixXmgs9z1Mdm78CAo89gP+J2h6NeHea9PXtORu/o9MUCScjz
cn8rkKk+yoSy6OvWoFofcyBXk/r/nNPTe94E+DhxTKFYAEraZjCTCiZcjjO0m6tF
Y+ER0YkNG9K23Fy36mEJlW8zes2K/cHSrRn00kg1TJjo9GNbd2lDJ2eyUkhHF0cv
QZfbu5kJ1hYKufC9ueM5F30WauqPS6AK5tOaz330s5ft05IyPg8zL5uefcKy3HJl
9lOZOU09SD55rP5lxYeRVC80p9TH0V2YXlp4beXgLoe83NNnk4QSNp/slgIwUSQY
t4lwvHDJySmrDh6KUcylxQH5QVHLQQ2Xlnhuj7As2O95VkGbZAapudyzbQc0+i+u
KaXahSiCJNPPgQAOf6nLWYCsvTT1AN5o8dYKdEpVihdvwWA90Yz9mXoOqK3+ypxL
LWG/3YW0Mb4F4c08BY7WQwtt42SNibDv0X0PQvTrHplVwx3eeqJV+90vmF8SwcVj
x/OGXW94E0jODfvY3F7z83p6xmYd4fGVefKlmneH6JjNyf25aULazlvGs4AuQkdi
qTJveabUvOcrihobKgjcNk14OPlbppaONIhP+MN6L0fuTQWnNMMm8/0dMj9oh+UQ
qKnXklXUKE2mc2QhrQZ0vbBELyrzcMBDPKUmlp0XxqlAfLaWODoP9IN9a5br1TcS
4ciI+Cxc0ccqfywHpaPuhVSKDcPhj9VsePTJKTClsUFRh+Duc5r8NII+J5yKobp9
/tvycuit4EQhh/kNvriOE4knyt68olJVOk41RUksAcvO83hmP8VihwKZgEKPE4TC
uK6flG9FMdDcWLA+dvA+NITch14iW44z5oyYZfMFCO6ZT28xxgbSYLxYTrX33uec
svUq9euWYEbvnoNIZ1KfMQ==
`protect end_protected