`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8432 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4sSkgcOrtFFGmnZEnVbxgx
+l/NC0KUoptgPj67g1Rb637ea0Q+aslXHcQGJo7yF+njaLln3BJFz4L1xs/1BSJK
MwdAyk+ak2ox5VJexDUXorHaPOjei9G8+7K0Tp/frwMtZ+6tb2QiYSE1HccJmtwx
8U0bpq/MwRtruNd58ilQR+RdznTtrVAgcXAqptBU/Wr5xiEaj3AdcBi6D0VZVhlu
FsKrh5IPSKdm1Dnl8OyPtzmGQoTFhU3cAuWoL/4R/CuciGjZZszIGogkpA/o7i7i
2wWFPl7sUAcZW+iXwZXWdyQ66Rh5J4a+x/w2tVQtaJG9ZeAB7JZPDKKgSPEJ2Lqj
HMjUsEcQm8ck+sEewaaYQX0OFSbvDTtZflz1/d+loYY+gi90wWGDgC7u5S1n5Tma
by0N308QvBsfijZBF3Ot93k0T/XTCaPegsacXT/oPG7JJvnkwkKxn9ZnclV3VC2U
Cowbo51EWQkeVfuypJS2msv0yoEY8XjZ7wTMmmRhTVZE2MgTEcgKeStAKmtyFNPp
uxCMm2jFqSWRE6OPGKN2UhlP+zocazdb/ci2DBjaogsFDd2k9mGMLSMWhEaPRizU
Q5+wD7frz8AT4pOd1MXioHp8kR8JJM4Fc9n+XxgL0rU9YmGqDyQgIWs1XM1rUN89
e1t3lZ0IcnEb2Nwx76byaM7qk+ds42mAPUr2IZuuQoeRjEzoyBPhNgYDRDl3MJP3
v+VhrJLeysY3hI6RCahndOHS5Kka/gIkCSm7WtP++dQzEDq+S1d+4x8GAZjqOzAK
pm+YwiI+swkZPVp5KyOck5Z7NWEfWWdtHDvQ/BcAPXZfi2CmNRV1M9IOrg5pb1PC
lwoGanSMiH9o8jX0xSwitziXK/z2fcFTYaJq+9xe/hvbVx8xfWFqVTy3ikEH2Eg6
mK5Ab88BQA5zZDu65N6DWFc6aIenZbGXD4yndWKgcRe+BKTpUegclPecl/t82ak9
r2O1UkQIutZ0dMgDdKSW0UKR9DcF7gaPWBq+tGF3GOiwCALQaap2xIn40nreq7hD
O/V2tyyMR4+mRlsd8fFGQmDps33kxUXVZfTzzsqc5ita966JM7WqDPNLzhhTQ9/R
P7nScojysJkSTksT1EkMvPJbV398zjpRGbEcBgoTh11pJ5WO3JpML+OoeHK/PAtt
PojbSLXUv1jOqaoki0Dte+2goZIRrRNQ7yhVRD59yiGh7BEL1U/Ok3JAD1RHE6SG
rdBwKO2RliCSdFGXBMj758jhrPqQtK+lurepGObypXGyh7vrNPXUiD039kpuPBO7
8PvA/2qjMbNWN5avhzbZy3iHYe5Rbw3tCkUGzevaETi3Ix1qNVCLwetXKPzOBtD2
HZ44mH52qrqGzO7cLCu5B0OHQ591K54eICV3wjnk3mq5I6/iZ8WeJXI/O0Kr+d5h
pjE3//8IZpqSNfnGYOa24DD25edqr5ZDXtM9zUMIbxG7+hY5ANIrRpWJ58uzLxaR
f6bSr4pLrE8HwKwNsIX+6KoCoLgB51KZ5X2zJEsHKJZEuhrIqXk6MknBVxbsVNKE
l5/L6aRmAa72smO+man7eiCKhVgVbv0gWLH9cwrcoIcJw+rrqFbzfk0+o9AJ6+eN
zDNw9pZiFmlLArXJMNIl21yGDEGLDMFPP9d0UX8atSURP2U2wRw08kC9i73M3uY4
kyFyqtlgOLBVOx65a9NmHoUVlYyIvnsh9c0pg8qWG73Da2y74xDY7711YqGQHoUI
YDt5dOFiOfP5718vtCFkPXN5lSXtTlEUs/xFZ8XV6/422azrZF30SPxpnAwoHknV
THUPMBmzgZaq1reS542mZ+KHCMX/ZtNeB2bBcmSVLSYTQJqjjPXn4tWeze7u/W3l
OWlTYXMMTdx0bKmC45p9GDEiuvQitUbYdhpODO6SXzF2HZUdOj9PYOFfttFzwjX+
CcduLpYBmxWuv3QWbTu8L+uwGNqJNe8xnh0+LGQD5dkng5NSVTahn+uNjdPXIKPN
DFIAy3OkA3hP3BV3mbzwQ5WWu/Dz9gEriJDG1zHiYMKuyroVScgqaOEDaA9UftWL
WpMaUWWxxbt3ObS7oasqPzhT6Zwt68+RlHOh6LZJFP0QMtmFYjU9Ag7z3IRcveRt
4cCh7qfM15t4EH1QHf98koB/icXg66xKZh3+5RiJj+iY+A6IPL41kH1ssE8N4U88
3ASREw2Y0PTz2380bFfaQvC650GJXvf5NIoGBMzOP+DQPX/r0AWBW8H7Swk1u61Z
sQDZ/wrsf1jZVAyHXr4nF2KjM5OlaH9tmpuJpnPo7SmcnmBPKvU9ChKp6Qf0n/8B
XydmaTO09fcPNgBf6HLy498j2YNCU9k3s/u4IkA0CaEM5c+FfP2Z6dDoDN741jKo
iQ3SKlm9ce9ojKAy7SF45WmCPCJkWSTm5P/wVk/f2bfvC98YhFm3E8dpX+HxMi2a
9PerqJ6wf082P5OtyjmtSOdHzeox3PgGKObf/iUczuMSU8ccD4rgvSvDruXarEeS
s0i1SgnYPL4TKWLxkcax5L1tLgCKNBOqBWu1gZQqI506WkeBt9xmhZjfM2fL58Bv
FAWyNcDtd808ODKhN5ejSUhZnnEVz14xyP9OTtc5uAsEpaW6dL0wGC2il8IaHpkq
2gF9khDGLTqZVmSKCJ+J6xdMmA7BXMtCTCZybFEGjy6uRymUEEtX3+iAtxh93bRp
YUYEfsaC8JjN1PCDcbrj+sBba5QeBsnJDCHgFivYUsMsO0bxjSmKJDfYmRHv/UXf
l6bML0GrT0KIcGRRt+JvO/f4BoLE182IkYm/MNNRcT1NZ7K32VaAtbUF8QCPhyqG
KhfDRf8cAuOzD3qDRLNB0mq1pf9VctEh74QTugisrwFZkDVaQsS02jtgBxTq7XBI
OqQ8Vd0VeXdid15+F3RkIlaSC34n+fFuybAEb3mfLU1eiPTU+Bg1HOR2hC+hVRPy
vau6YFHviKchbh7GyzYfRbeKIZ50VG7eDRwzxvICbYBGIH3RMY7uIO98Y7aGWcP7
c2f6rOdcOz44cOsZEVCFr6IuzdgezfADfOMH8JoYgY/OUF/JJbflO+utlT94yHfs
Qx7llaUtf6XHg+7gHhz07xJ6VASqVdURJD0PW1JvBb+L9hmHGrfVZGetHkijLQUs
Fe+mh6eRmO0lXldnJNid8zYXNhU7h1rGRS4a2ERZif7d8xXA6Ioiqtl6A63OXF6w
U0P1JPSepPS+6wzYOoZXqUZQRHv+8+FChdNIEmiZZ7c3yq3FV1Y2vn7OLZdvL0H8
sUFIY28fkbSBQ1jXSt7DI60/NSKRZz4xZZvoaSvn/79BVbfFgqfSdzCe+k2/mkb7
u072DpUYLLOlCHXWYXFInqTLlPgFnxZ9i/05cRg4Z6MeK0w7UJNSfwIYUVK81/qF
eWJ+36RISMflUoR4d+cvaI5mzsqSSKojxxd2iu8yshI2hjIA0csem3Kyw2awzoVm
uBxepB3ErKhR6ZX2nAw8jttWc8YITqXH4piiG0VJ/5kLFbAXivU8Wbr2qM30RWBo
glwGiHYanD/zbU4UrBxg+6PTOxp2ihpL1o6TeAeraJeswGhBbgNRqReRvwCYxvf7
Lc185eYggFv5C78mU5Hr4h+zDP/7quyg2Z60IZcIKun+tS0z+Rest6ye+SwPOHRH
qS1X2+vNOJCPFt6Rn5NicgLnMBReIyoUkE2yQUAZ7FRmxCo6vsRVCNXqmzFV7DAU
SIrNSVNAFsoyITbdZgJWCyOiQhFjBnTVdg5hbr6xpNbUd//70scgHQjtPS4SIP/I
REx7amwSvh6pyDO8Hz/pX+Zq2WqvMA7652harkTOr9zbTxdhn2iqO4HNODV+BfEU
R4/NXV4JfUxsVOGxEvo1IeN8cCGYKOoERwlGR4HX6E45wUyZFqo8ShYdkTFHBYPF
Rl0c9mp9pBERPQfBhRoUdwAVUuAkWUARIw+GpfVfBNNxhV3hPgm+buUFuw2uu44n
DC1b7jTayzGmZfnXmD2F1iKe8KGYFQUAxq/KZFx0YSG09oX0ZlhJxvYRC0oPEeZ6
5PVm4QOnHzlAL/GSIqwCB7fQlEgmAY2CmyaLrszoZhgxsAifq/e83bxs+0GxTuIc
8ewDxSk5eTj5Qxd4I0xCuAhFpZ4CXQD/TtjkR8N57DkrDhysel0/K5dJ49Hk3iKC
0JAhahEMWore4SLSh33XyL767BTKLNDDZBSjkz+649zjHytih793K12eOjgacsw4
aCKYegbWPVSufv9RmHQeQG0O0cxGMuZR68X2bVm+83h1V9KAIiSVsa+GEAio9jrL
S5IHoIOe6CHvQFdAZ7+/UzXn7AELtkKEeBaW9dqafSmatnsraBMTq7J+3B81Igb3
FWRyXAL9sQvrCEuuTk8z69PFrVz3kU0tdhWXmY5B+vK4cohepdOtkhS6QOl14g5K
I51PSvWH2JD67NBEX0+ycka9REY8iH2Y6YxX3IQCGpgMujdTd7Vitvgokmmvqzfm
mxq4V3eQ1qUqWV/6VbOv8PcGnekrlVOim8OaTjDpeci+Bc9he3Z9qnTmBP59buWa
+6DIHxA7ESIi2hRS+ECGDOeJOrniaQQuzJiDioGjK4ERlnoOtby4Yf+SlBXX+51f
RyedprxxaNBFiKsFMY0jxnguSFuSlisGxDp0ptU72ovaZSdYMQDE/UVmEbeuhkDc
Vrjy2sar0nVllpmFFkoETloEuD/AiabzEZlrFkHQeGvzwQWYdrUaXc3n4cyzQqs3
ydqA/hRavZ6m+6rgqzFVvkJ9auo3HrzlcK/z28PVf7NYEkGgJE+1TJbC1xyRM2Kw
by4AtjcpkP8V9c4dFTVJi38ntCDPp1/1pyRxNhMmMcjoeYFNZI+zSJHRNiMNhrI3
6CCGa/qmioKJcVPGJ5inN23bjbtwhDvnqINHXJFmH7uX+mSWiPLYTbliiHVoHQQX
79tKrN2IGV9aZbfIhIHAfhWvMMrersoPDjY4WThu34cxO/7gwiPYRtogS1zulvfi
BFGcf4cJfMKdOggL6EgNd8Muj0uBdqKjm+df3u4X+iHZh4kXasmcHoUWv43o9Tgo
LOI/GsUUkK/ICpFXrqmZgEqgNrO5BfnGYX7b78NEWv/a5DanVIVIADMclQErz3bi
mEqWLet2trCVtBsBL+9I5NJdndhPIwL2i5nBL85vaWe1Uv5whZwCQEfl7WqJSfYy
hokrnqbAwj38M47Hy791RP4RXYOIp72XtxDTIgw+65bkK38rpxkuGp1OFJeoHT1A
0beNnGDY1wFmoJzbl/QZXnxrs3TAHPNFFGg3F7moHZrIZYDs7AsZdERTEKYG8nSp
q05w+ojZKKyGiIna/ywJEXPvkRap2RN3yx/kLkIXedk/+7qUOlm66pOCdIx5Ts7A
lmLlBlQ0QBTI7ttwklAGai7W3e+X7RGv9RwfJY68tQFDiW7P5u5TUQ0s3gLEcqRE
KS6fdPJWwWZt5qpW04HeoOUNQrBcsiFTkyT5NFNGffnlq8NAHvDTqjVZFa+Q6E5l
R4/jsAPOx5QK/J2NIEy+jBCOhvy2LwKyPOvhld0FMQeQkfo3ixe6fOkSAR9U5YCg
DqpMuR2uW4hDLEOBpFblsWU1i53EjuZc1IsKZ2cpRJhSxasEuqtosrjZa2t3MfxV
84iOXYKosiqrV+JPr+KAUlymOx4d2rdd3RgbO7AeBR+zBc8tccLJGICZuSUWU9Lq
0q8SgvKtxw/V9ruLuyWfkyr+yDZ8b3irsUzbbRH9SrQIpIlM3emXTTdKkX88k5B4
LUdljawwXL768MjQR1YYJ28f1dMPUu7kXB+2VdGXiAzDoP6wNSJunLnRbRSprgsg
tA5Ugrcx1P4pl1Way9srNfmi6fHYSIPhOtUCcsU9Bgxak+hdSvS/BeHnhrsaC+y3
0WYY6l98FHvXf7O7J16Ee1O87ZHqtf/MWiBI+57SoLuvLy7lWAi6GmMpjP3BoQas
/YQXKweRPlk+g3bUFIt1XLsRCn+3DulqJ4qu19q/UshfPRwZTIggsVA3tsEs6wxl
9/9vztbSYkm9nxyT95ti66QRGDaUpOBUPC5DS9ensUl+Z5Ht7JwbgByn2mhCcxvR
n7Aaj9zXSln9jFMSpmHDoqZf91WGZCwld9b1TP1uN5wzCDsEK06z90DI59uDlwqY
snum7PmWT3LYHWXP6iIQOqhCktogasj7jZtpr8qsVZAQdG8skCpSi3uPPg/MQRnL
pC7vBmctNys0vX/GcJbsP1CBzC8fpCriTgPRiYfjZmTsqSV29ie56Xe/hVN0OvMb
7mpxXTL9V2qrEktezM07PTarYXCF4+UeUaVLvbMnzK+20jClK6zw/jwfvko9RL6/
gQdL3w5cs7TVisfUT4CV35Ij/pWW2dnc1bjxrZbDQcUo+EjOqiKm+e7w1RqhN99t
6bzivP7kc4N074RYWPtUoc0vMq0Js0ho77bEIFIws4Q71wQQoscyOzLcoc2ZYtU4
eVUqXNPzkDFzxHs7tpQxuEbd/ARY9F6sDgrMlieNpNs/5fvBIV1897Ezaye22fg3
DNhe7kJHf7jGmAyoc3Lu17CenYBW6vamTH7Ta9LdCc2ui69ROPE27UeNDRSLZtJT
/Xx3F4W1vYU2TaUHihgTWf/7Cr+eLwejj/ADA5sEs0nts++Wsbt3+Vj1eR2pneyo
GgZ36G/OTo2xVk2ZzWTI9HrhDqgHFazSgb6BOlLUDWmAxDPBh+Q9JPc3jRZWEjIe
U6xrsxO3HHBCIQXvF0mMGo7RDybo/Pny28qOMYm+yNrqw1/IkC5nGSGZwQWlSrMT
rfPrluSO4ojFL2brg59370eIV42EfVVrd/Euui2RmcbOFWmQdOdaSxvsvXp6wvHG
6cAYkbZTlzW/x8FQIVQgAxTVCiG66LzhAB37AUeBWRN2t2PqURDnOb4kJzZNuOF5
3OELAVu6gga7hkl5AEAksQCeUkBZa6oeTFfcwlAUOTEKlVYe8v+pPmje2AEafIqJ
y8gpucr71ZZdhhv7u4tMf0SDCZm4MBfKkD3OO+6xQOg+nxGClds9juFImMjPUzP2
uI/U9FElm8+9CKojZocH1i0EIWkLoyr3ULIO77ONmPbL9RKzABScLLfkiplgScFr
7k8v7kcCKMFqgLCVy+6VSjm9vTMwhOvW1SdeVyQMMnbMuzlSZj5fQ7lvyZRjhSXx
uIv+Xvwu2EjJPrljKj3qAAWbcHndi+aRp1KT1rlo/kN0lMsQdtBwBMddUSXgQK6i
AeYgEMgoMEUOk3jaKJUwAp8rtkbhjIzGAxFSSiBkT79m4iEkmh3qJL1HLSbOzZcc
NaMtF1BEE38hYgu1iqAmcmmfx4Rve+s2DiCLppJasW6XS1cDhteM6kvQoaSIAWG6
7vrpbaJd50nql97NYTimJBxUblA+illxP+Ql82lX+kbiwUhfeiuS9hhZqT+aJuxw
P3fogoe2HqnS1D906Z33dGUletv1/HyCV+G6jdaUuhPpCnKJwzR/+BAY3s6Tsdg3
2eTR4edRlb2CifZ3DIX7LnrEbvYZoyYZ+IS99CTxK1xpFX7M5lceKsU+JGqMs6iu
YCuNFHCYvbXPXfivVkUXyRkXvaoZIyiZfv1ZJQe1svh//IdNqrseb9IcPc0keAJa
lHEdvCJZbMWfDNfbaDTSzEhi9FA+A+QN2KCPOUdksnTjRcEQXEWyv6K5hxT+/mLZ
lfdnOeAt2/gLUyFcO38jau8mu0AeLXrUBOyUU0dcE2ANVbX56kOeagGC4zQUff7e
rHwPw+eH7SDgs/xktD6pw3qQOVbtL1wZPGQYNQosW2vbBYQMPbCXalEhaxrglmlw
6SJfTCX+dRHeZJ9ycwmFTle4BAuU8G/1d9GtotqlELW8CEfiiSof4NzpK4LEl++X
0w1j05TS6xQ3/4CzCIAViOp4PTMD49N+OLKrIVx+xT47b7osbnoO7zwvnES6YaxG
fzLtub3CU260ugk1me8af6KS4hSFl9sckD7XfGo1lYSfIwIpLooLO+l32L5LyhoV
hiG5GAhCB2dJ3v2GdWoClwdHaPAFOXTWyHxznnbzIYy1cJy7dPXeaWk9HiaRaCuW
mQMDofjb2DR+giUfD6R2L791khyqmaa8X7aYly8Y51weGCaDrIKtQFc4ikaPNrx+
8P/k1euvHQgSU1v61T1AIoOb1i3LXIRhmtjKQfYo29PZ2g8UZYa5e8t7d/lIcANJ
63yZoBDbAfuH4HlfqnQzR+8XKjyt0sB6qdopwGYMcsIaEFKDTCV7nojUOfTTcVyQ
T2f/RPACj90msxm+qjZ1y5K1IJq1Q/pTUVw5cw4Li//9USdGxRaftwEOGU+j3qUs
1DLZx014KrrMhBh4tQKYepILhbqrY3h41CwjhvUxpA6mO3oJtBYZQTOa4clhI//j
CrLRWQKQ+TtqqzNSqcgHenIK1qc/qn27gf7JxpMe+CxQa+WmgFidaWaGVNq6KiDt
OWxfRCujgonYkhKup0WG+FypiQkIWNTeKeu7v2322DQzinC28z2DwO6PsEHvMe/v
E01qfjxfAZPr9LLhLWHoKdR48z1gXVgUi0zeAVGJqCT6KSm8guuCRngftOTZsp5k
2nv4RRh0ioB1szjM6pLhl0Ez/XzwJoCPVCcORaSQ+gglJoc2oK2e7UsttzaMKj6Z
C/2JQOWz3dQ40KFsn+DRTN8zTJahatrsk26WhIEBFVFG1CRJd25CZSpFtlFmGM20
8ZbA+G4kS0hWjMjyAnIBtq2xescuBfqHsMYX2GjHUyN80psrljh973+TFs1O5HzT
P0vOReSXqI0sITVz5C1pRdyW0paHrWYUpgJaBnmztuPS5L5JUl+bppqDqWuWfIKj
RmFjeRK2Evtz4rOa+gQR0uT/pJKToVanTEiPWTG+N5rmp44pFHrKoUrRXA5wlIwO
YVGIl9mBNs5syKUO0JyBjQychNgBjCVQj81nAywTttRcA2QGg62ty3Uc4Uw0EfoQ
O9gMPZlJDVZwW7n1Th88+dbexDEed2bEcUz4sWvEwEbMeo4AnEkpmqda6+8kBF6r
TUFAe0QKqkxD+Sny9xxGsvn7Akg+unNX+vFhEdeGbRajDLl1NlpNmHoSIwjdrFKF
YrH8/KGeXo7Y737LqoWST7UfRt2kyDBCaSqyFEepcc8vIvvbzWx8C7r3Jkh3F+kI
KeMacLls7TQwMvDemZKsxpu3qc7eqAIUMRtB24c1+eqX5S9ZOg2r2DZS3l59qwgH
tuZ930zRbVQhxi9f0CSgS4hx0BxLV283oCPLfZT+qU1V3SzVQZijjf1aP/fAWyv4
AntXC3GWPTYVkLvt7OFT2KX9+/HTmc5DJgWbKjobH6FCOEZ1hRsViV18t1/z+lf6
oZdVYkpySbUQwQm8VQi6lKADNy3MFd8ByKl+cLzi1PwFl3VBuKNGjWpVtOBBzAwK
D2SZMghVntBcZwKAzd7uAZvy8pKu17AXjiNabLsRtWVEH3rP+2S0zgq+Ptm34up2
7bfq5YsjL5NVvYxdR5Sjq9nXjS5uiMvf/k5eJN02HOclQEQ5V9lV0oMezJ1QEnvV
W0A5d+CiU86Vtwj/TmU4LDx16i1YFwhTsO2jpLSKvWOG727dgIClvrIykTgn9RlV
0j0sIUkz5PsLw9EfR5REToIsco+qiV+OMN3kY2WSprWfhTSdPr2/AJTFIy8gIJzd
jVdQBxZC1agxiNsJ0xRzxCOfLx1pcTk3RxBHl6XOrL4QoFAPMwBLpN2ApC24IwUm
VeEAJOYtSN9sXOJ+B3nQzqsvMtgM7R5f+1GzfTuZaRqOPlPl7MnAr8wPVEZ1rmnF
sZWavUo1IkDyjXO+bedKdmtJowI1QAaqfpnTbtcw2V/1jtYb980qcxvORTNFe1Qh
ML+Kogtx/s5HIOdm/rdrRm8Cy1hosDc5D0Un4Vkw8zg4ipV3dsMaLTB7mLqrZOSD
31YBCWvjlq0tprCsLhd8PFL5BXEbV0nZJP1IvNjF/Iise6WuRA8jsdlEp29IS72v
mYbPOlPX14vfrWr+P4xEtKK0sXticiT4zgNODMeJNThWJbbxA9cisIyWHC2LFKKk
FSYx63Hr0uGVtOjeZOVTr6yyt8hMwgoOUWwv/0fKt+OAfhas/Lxma39KhRmzSX6T
DELL9Hw6tz6/B5jT1f3tG6wqxb4K8JW4yaXXnTI2GsOqY8dMsZsgc/iGa7Rrij/R
E6HNLoumeFInCNykRZtU9JDKQOMa2hpLpkILe3r5aTLh4dnj9ybo+l9g5wTIL7DT
13ccNw211+3EALNa1bWj1IDbyxeYEr/2UrHn9/aDYsKmDdyUVW+YUhmK21DDQBDn
ehoPheRstCzVYoTIJbPxS7I4uJUrlsrozeFze5OiHTqrbSJLbQpRAhIZjHT6uSJj
adwPsc1Gq6FEdNuatlBR47t5end+DfNRj7lPJAG6Ey06f4+WWvzl1M6yfuq4SpVf
1aTWOWdlbU7jHZCS7AGrZti6dnpx+1gY/8znlprG2KVzeVm7PkJrybd7rxtDguFI
0anenTowggqFXV7Zt1cc5PQIDFDWFj3aHDrE7ug8/XwprFDQvcCWfJPkQUm1EUlT
jKckppNOBG92TDC0ZpY6SWZi1nT4OQR04pCxpJDKGWrfdkucvmXCkWa+reQr2hko
tM39UQN5EzpRi9ksKDX5hjdwoNRriuxO7FD3huRWOTBHM2Xmk7heW7eo8vDQVE34
gWmNB+nGdsHXEklwjVgvRm4877h3pN3S33M3qnljBMsmT36i/aeJr8dD7WPaR/hW
X1dyyin5rAVBmmHYFxcwUtU6fG7iwOdyAeRlLRK65VdJRFX8Zk4/RqnFcUDKiXeF
Qrlz52goJ832oq7L66PGxAVtq67AWikVdnBAN3ONTdWzkvq7A46qVv0EE9WEYO0o
s96N8JgdYDZPf4CTvSbcdfFrd8aP8XAe8QtDZcm9zcxhiUBIuYFU6OslIYsIHCPo
asptSJZ3JIGarSxQK7AITTLLZf22+sRLqsBsTb0TfTJqg1xezUgfPu33QtXhnelS
A5eFWR7EuIKE6arZc0b3C8E4uevZpwvRp/zqdkcyyGUg0BJz1OQevqF7EXl4KWde
i25loS1eMCksIMbNv7yuq6RoYw5OzMuKlTFaKevQVWQ=
`protect end_protected