`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
j9eMmSPGcKCWAR9PvkqZ1R001FU8QKTyJzFqNLn+qur6INyYDE1AI8LWcxAzfnTc
IpZG7ua3uuk5/kQKKQx8ZIPLfmv6H3t3eWjki8YIAtY/d5E7Gq8Z5mNxMYRzGGTg
TCMm6oOrOTVYlCXHE0X9AW696Z7UGfWirVibl8hs19hrFdeZKGiGht4r09vHR+Gl
FQQmSObM5aSK5wu5KOrK5ZUKGHyBhjnIQO5NnittDjOwxV/57nHVg0pdG6JUqyvm
tEgmCY36RCMRGWN7sekPtNHjqpZkmYrVX1T9QF3h73+8ZekZYd2xY2hpHHGYYeWA
t3+Fmb/6NUmoP8+Pt2hI6g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="wX+NBVcG/A5ruHK3pkDqG8ZVPdOz9TJPJ5saXZYSeQ4="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
j/hqWUoxjK88VtH4QmjIrexFOSwtsLKOZ/LCP4cmrqgzmR/e71apdtoL+o8nlfy6
eZxDZMmrZmJGoazz2oK6kz7xJU85UCwNc4cxAsVxNdCP19vZxph/nCYZQ9lUFkLH
uLBkOeFP15CD3jG5/dp945fHP13J9SzB/L9PWvDC/gY=
`protect rights_digest_method = "sha256"
`protect end_toolblock="sqDZkaglKf+bDjC7VKm3lOELrT2Jlynh4UhPg2J0Q70="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1456 )
`protect data_block
f9kZDbPp4NLiAOFOgATj9W35i3s4a7wbt9jeHjHVcJxMoXY8rb8laqS5bNUhXGW/
MOc7UNc1VwolqhkS7G27SLamkGClZZtXSbRcN1N+5kZpEaBEj1343vVznnU2Dre/
bKlbmouB09/BfSaq9uUVg0fHIk58nKH7OEsqO/eVYVqsIsE4vaGVxbFRG95hA6XG
/+T8U46dNPuZbwn34TImgmAvbSgIXTT9/ClT7WoIlcgAySUQrj4fxau3S2Dw9T9o
eQoohwyt2Lpti3P4qyiZaZ5Jt+QV+IcrwtXXVRT0ss+5hA6OxunVCHZIboF2nmmc
5jTTJQfGXHrpQIBvEj0ih3mU9/nlngj/A0KACuJ9Y8f0hkWpzp8iwNkRYx91nj6n
p3c9uyjlArxErBMlL245s0kSLGpbinV7gu/vvLiLBVLq+hMUTARMZyfR2UqtF2GB
mKvvc3BBgCz8TaTbVi3dpBq0v0BAk9CJncRda93dQUo7P+F7IpZW1wj/dIwyIVpo
ziEwmWilRY1C/o4CkQB8M/VoPLipSqaOlmk6TENOFrBB5C9of3QLJeILsTa3WhjD
8W6ctdUClqCexnjoCGpR+tVNrH0wiT1RSgSRsdZP609teWk3hzik62W2FUPOJeaN
Z6cWAGON/6wVSlKZet9cx6/FByiuW8zMxHh1SaQTobxukHwt5Te0ldEzaA4cN/06
wqzV7YHh3m4XedpC2fpaMGm9RdJlIsbyYDFdeXjtbc9kqTnaufDpakYm+Yb13zuR
znkRV78Vs4FOcAh7VKpzhF25kuzGSpe7XHLuWRR0lN9DXnDaJpUpARstIyXKn5kL
NEwC0TpIEENXgjol0xj5NlN45hdQLzm/Ryoq0S3bLLBcJ1SIIUJbIbSnVDD4rXAd
IrzldX58/ede97uiG6hcf2ffto2fGIlxWvce5GlA4JnkmJc/RSDyZw60XF9URHxx
xhA/5fbA75rFhRuWhL9md9PJ/TEOwInZmDFhmhVkeaiyya/1h9XfY5muH3ZrkBlN
xa84454+FVWkPARbTPWvWnNj9HLVJOkSFLQO3NnZ6GMru4hwnBTna8B/M44hYaA8
XhfWFxH49ZChREej6jZJ1jPzcvAw/qw2Al+6VKdsI3jdQEsRjRQxTumy2UnP0KRQ
gy44Ljb7GexqNLgFbA3W39agVa22RX1D5F+Ye9zhV/xqpf+ZzsBDVtX7yFtO0QPX
F1SSb+0xqVLUBa1D450ZuVgEHGFP8UXE1r5tJnhqXTHetthv8r1GeroP4wiRsZ46
PeK5sBD1lKJ6mj2rBvUeAXG0RQR/IhoaTz/NHGAovOfimQRitVBtpcoU0kumwCpl
vZdiDs09S0f+ZMA5bjWexc2jHYnEEHo6sqg5azQttqjqBPsB9WR5BS9O3yfWUacr
3T8vmW+QUEGfb/+3B4MZ5ksvgFWbuom2WNCMO05ekpIGfbuv5/L9FXkSge4nXtMA
wl3D3STO6I8RvfHi+vMV2cU2R2RuTfXHT8gPBhIs3ccSoSfQGR3M0ddOGSUdX8Lq
t6NX4oPWGWrM5Vl8OPt3Ds4z3u/mON+ZTaGmlMbBxii71cZkV3JLI30HFdVFOimE
wP/K3sITYo0dv2r0vCW86eEfyyHg3EVnwwCgFlHAQab5bH1Vwae0M+3Pab0ZrtXH
FR84W41cFAkDeJmA9v7A0mkwZLWfSNPwanMMF5k//lqL4rz+v8rCva2zSTOEU19a
04odScCaqkJaQvw8FleG44We3ykNkBprGyjkfVGLgApMlHjGwYiNxK08mXj1D3et
y4vBKBhOSZY59evQqOKnFSq5/7LYUKfriRIJTpqbCYT2ot3k2HDpdB1gs0W8xjsQ
aJVnJzlmWUENwPVokj3Tx+IuNoRy8i+TKKNJd9E/0g77BFEIPdaGM2Y1iAS9/8SJ
479lXYUDpu4DBtXIc30f9A==
`protect end_protected