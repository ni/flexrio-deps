`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 26864 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
akBpHK9XojjdOyFTP3pOwlqmu3HKDkgfdD3J9PBzA3oSMdtk6JzD2HEtC5g3u++i
DRbeS7jdIhl82n4zJjciVvCO3sl5lBysurtoYJX1awsM8MTf0Mj9Fg6O3BTu/z8P
hlTZOz9t92ydh7zfiGt5wfdCFnW5NSiCvP/GY+DEdr39c+nw79kpSVf2cBDX421I
n6hcMkx5N+TTOYBpB4HTvW4tL+MTpCFke8IVxFvmtzbzvSZBb5Pb21Lt+gFexh4R
xxUFe65u7XyQouMuacw02knnrO3oFJdajtstqtO7WKXzB3IQd7ca+zR2JOKZhihH
3dhWyewHEZqoFVO/26fc6SOCtddoWAaXoSWL7I6uT+iaAUBNV/W2RVlw5AJpgzSj
8+v1tgxBRRk1CQcO+bfXEaTCTC3VZ1y4Je3AkCIz91Xso60l25rQxqQ7AqlT/l+O
YLHWRihfBjnEsfPczyfkqw2QDR3QsWFbQOT+ReSJmPKE4/zn6tEMX9pEWPpi9y84
JXINEnMQzFYLknQDgQ9dUP79TBCVqqQRtRxxI7STrYmAQTOgoHxPHNnMDLHgzVmI
msNDw9s6CNEwPpti2mFVgdnXhyaYBKgLIVrJJ450ZUjk0s6Rr9d9jtPEc0sWeaig
v3FJL4rNGUP2ZGrZfVBHKmzcFXQfKO3FqXBY3Fq6HCIBmPXXEEKC7j5J8IbMoJsX
XLwXgOs+NH/6qzNXy6GiImaP5j2aKwJTDyX1f3sXE9a2MOqXsaoZTD9oVPc2T0Kz
afZyxYjoJntrvGT/FusY0N63/Zx/QwXOiJqs8lw32J5uzM6kyllmbTrNcY7B9VYv
nmcep8DOytmsnLgIzf8MCi6FgHg+g734SXNCnwSNZmczwLlhEjlrzHqur3ueASTX
SIFCB0eVfcqrKlKHUmJB9bvfP9v/Vu1w9+UDz9rr0DmOtbxRSYC9efT49X5IVmX3
R6ClA7Cfgb6j+e/gYgdmebSUmpyE5+buIgYmRCUOBZy4Mc1VZIgx2c0uPfdDKgNm
zp5La32q2ZaEdS1SbmLqs33iS7z5XUjdACSn2RFMQ7jgoXg57mSPKoH5qFcOd+lI
qLr9FWFEAy1aFLPDBXPsfZS/h42FZDqjDCcthHq4mq460LPlNzsUz7pSAsF2H9PA
d9YcejI0Ip99y3BheUEufsvDBXh9OYQlknBArqxHNyvHWjnJqXPufFeNJ8/JnKNC
e2r7pCitlenzgAkrxBZnhDdl5HAUlYiuqu1ErH6o720NA7BMpe3uLtUWJlxOns7d
wHREkK5XEwF7Mlsa4Sw3P0BpQLIE9UvgVjEhwRni/4KARx0OesBCDDwTAf/GEDSl
ZU1bqNqxR1ZqAAiK1S5S/OGtiHab0WI0Jd+vZZTqMXP85RY+4EPn5UIrFTNtXM3q
BkeTqMe0vWHs4p6RajwmzUQ2jh6Syc9i2sAN+hvCEj8jUZo7GjsFfnLd/+amn+US
mnGh/438cgaqnDViZLiBOhxc/9Sixbf9ObwWngEzuVOs6Zk5M4Rvr0U7G59xEXlS
O0t++pJzzyzXBwN6lThSHpgcsPiE+7wxtOXi8QKMQpNlLl3AVom6YoJDWEhdETh/
FCr29w6KDNdtpJ3U/zfgk6ZGYRpeX3WV6yxZ94ByceaC/ORfUwWL6QCLKedY+2hV
VSggtNIjIMlaz/d9OMjPe2WkYyNCdNm3czQV7NcuZofpITBWfWriSGY4B5+UQUNi
n19GwoWiACQ8esymZtCs5pM2Eaq3OdqSH5j1wIjOt9bZSZ4QSO4QdcDLJYdbm1dd
Vyxk7RuTQuVeoeqRn9Fw7Ip3L/N4/DiWmPGetIXZ3NF9gURy/gOybH63E9geUMk9
klGy+tg3wCReNfgRxy3+Cz75B3qHz+EyOaJqH6wveRe+TCP5p+llQ3WzmoqpJvE8
dDKVGmvID4hsYf1tjDNWXS24jolwUZl7LhO4mdXhVBx91TwyR4HslyeY3zQRTg8U
zoktwDXTPiNS9GVZQDeQ5oFzlY49A2NSqWG0eSzlfUAykPr0rIEC/l8wM/xz8WP0
/NXP7/198/1E6nEwPv5ArfciV8Tpm2ISJxhdzaGglz9MpJ+GBuEq+rdse0RVtZ5x
WoZxKb8XnoBMvH8nwCHRrlRvEtbehq9Bn7e3gnBsTvWj9BgllF3xTqXh0qL+yrdW
tUJEZcDWA4tK+Lp17KlDWBvPv48YEm2/L98AHGXJIjKqH5EK3iG4c85iqzarSZ7y
nnWLluxdJVIdrOi0ODLB9BmZ90BM2e/Hzn/CJw/uVxwRnJRYJtjjs/tJw0Shnf45
yfnnVO+HPaSCZHzPLMYpflMthHrmwJmkJvtlStWh3SICHgxVkE4FtKlnMCfPRL3q
J5y4S976bqxsEEJ55HRbCxvbD3g+usoMWkhQIbeXk5jhxd4FjYfRDlOisAfS8C75
xw1Xxx/g1KqlbB+CyP0PE4xqKodrPktbWyAVVq+IlLQdGDSt7/KrTTd0AndGzI4F
8kceE4nXaj7QSF7rxWKc+CMAmTn32FZXpPopDYlOLGVcDcGnMZ2fVYJP4l3KFSCz
y+sOoGP5Al/6e8n3jUtQj1A7O8xeEEwLfT7Wyzvz2ubfVX1Iro9g6h4LISZDxckW
RKaFLp3cDtvnv8xPafL7ipJ8xx0is9B7HcAJhO4WnG+Q6vsGuHgq1OV6+5WJ3ke7
zAZ9qOZNOC9L0+Bs67QS/txnZjsPPlpDkDQaNdeqnCcVZrXpGUF8RypKIF0700Zd
RefCCxOTU9oRxxz040mwa+QGJWLx72tuQBQU8ndOnoFzpYOlM8cfUoU7soi3nxF3
uEuvtIGoelkwZQmRu1px9hJfr/sE522FJrlvWsVM+3nzfEg7zVwR4EfYkcaVkArN
7tigLIgS9mITQPAdR8GGXAQWJVgemvL2LIn9yI4kChbBiSZyRiObYVUxgwfpa/2b
ypxctT5hQborc2TSXO68MXQfnz+s8PXVgxJoOWc1x4bG2y3rjwgfa0KTekcEkfsF
rIoBJhmyeIYMzgjSNTU4mOGxlm15uA4jZ6Bt6Miu/qDBX94z7tqhmb2Lq7vzS/Vq
lN2ojxHRyZuNkoeLAzsLzL5OobNltYiKA7mckp113PTw9kyy0ZSmS6Ai5SfMueKt
iWxuvTW8s0MiJkrboNRSLJO9/nTjQooc6j/JQZG2sLsG8bWJ9Tfdz8kYQXN+WDn0
ciXE+i+s6NP/ga8ZmsyHAoBi/FohOof6bui5wjCdzvuZnvSw0Dzy88PsArFf5h9E
Dgp3j2yOJ2p3avTnFOyzaj5J/AN0uhaVRFCGYkBU9zDyqO+OVsFM8OtRku/Z4fnx
0loQ63BgT6ejDfDwkocNjAifgLCdsHNTC3qsk8RPR5PxGRYkaslxlNjmSMPfWNPZ
mheKGwltwoC0Fl8osNloQRT9AkwkHcyNO02qFtiREnssFmK8wbuUR57451AtK223
f4Gs20DtLZX7HAT8Tdbpx1om0QtmvafZk1wUW4N7c5r+ZgV+6TOUcAlHS/TRLc5p
p8MokwwFgdOdgonLTpEX4W2heQKoaF/XyrGWn8RmceGgAIZGDet0l4MgeMA2jBJM
M3eHqsiwXW+V9izWJh+zfqm+QfeAo+GihcroqMvxfmVmE6r1pRIVNUQMg0v5gjpM
yac0vnW2RwWxT5mYJX4yaaOdYFnjBiIJ8nuNSVL9e/CtXX0+DItmXnGqHi3VfN+L
2JrMfdMnrl/DaNBUERFpPPe7s9+ZglxLcYM80HaQH9sThEkejwPHLR4RrXfR/GWN
ml/MPvOcJsDvbRFdfs0RwX7YuGi1lTCxABnQ5ivMrmgP7xcOjRC9lYiq3W7FZcnQ
bH+RV9xwwOiM8ADECoblzzHUJW3Zzic4uD9MtlYyoZKPmG/kj/0FeCPkpWkLw1BP
jbwRFJc6j0r1YBFstBJGmJBBX0zd5qLaofYdkvP7+ESO0JgRnRfLxondm7ouLPR7
eGpNk8zN2d7jldZMuL9VFxkA9pJp+Gf5E5TQCDo9WAt1j1STJ1ndHQvxVIfDGt/5
CReetX4rPR4qnFFTQrrWjnZqHQRSD+Fb75oHRVKUo3xxQBqYyJaMLL6lZz5sBZqu
aF5MDj5Hj4uopjAbxtVkRJVRA1nbATMthfoFObyBPxFierh4gxijEJRF3cGltDbc
b8+jCG8YyfWeuuEAnpEKSv2td2nIOOvSdgH2+TbD9Fz6xGAB8F64WqumJCUTCgJr
MMZunZPRiIqB31s5Ir0Qt3zTjpqAN7W3//5zgVWQRdQ6WJBWyZz07uMtlgJpLuDm
lX0ds9Cf8yjtsaj99lkyx/jk33w/gOUGdbH5j+TFwFVxQiWb0vQs6fREJcC+tk2v
75XYnk3wMKBMmfqN5emoMHykxPxbtEqJXBoWjDqkjlNjvKCu5FaAXuUpwJ/7e7IO
Yg4kfexh/lneG7xqwtJNoMXyU4qD56nPI/Qd91uJTeBK5QOA/xoQx2lHAKyLD199
flpt36DN7zmi4V9YVWDzb0oo5pER8COSfEDYDTlak6IKc0TktxAel1IckMwYpNAY
dbZDb9YXKTDVLw2C4vdkBikdc3ripVMMzayW3EPtEe2P1An57n3vzBSSiink1OVD
AzS9egAoaCvppg7GbNHTCE/dh6ufo7TQ5Q/IG+z+ktNuQA+OBy6xTo0vMAYgOE5v
QxBpkHtpw7IEWJyQLzQp1ofzJLrSkQ6uT0W9fwJ38BFtTC35xLhdiEfTxiDZBdSG
n/fascHPXH6WpGBJY2xZletViz2ZlWDydj8mhWVgrld4gp9plvQGi0NhqbeGAxWr
8r1U/hvV2WEYlq6ET5tV5rITKtxB1tuq8PsaNB/6N8sljMYH9WL2/BRQzyRyRYcZ
wjloZBqlRXRj+bxHpKFPDhGPn7hfUOt4ls4honyy4SrA7NEMZNnK5n6OiHpCAppl
wYcw8i+xgOTaLE/y5lyveh5egt23KaJfyK0e99wGI2/k4ciPS/3huubhkWBLy61q
aKue3unrNK8lURgTEJPKoL1iRnMZYyxABLkzZ28i0f273yNv/O2OReFRTib7IH68
M2FI/r7B3xazfvX1m3mdktBmeHBZasqWoislwEaXDUvgkau5aY7m2pvxh0swO+hZ
Olduv4kIW8rO3AgrOHvU9NXhM3DvYpe9pi+AljHqdjVs3n7+aFVHXyfdRGIr+jpV
r3T5u85/2UoOtsGGcAaD4ARO/puZiwmv4T7UCnCpVB23fhpa1BjKn0QqgNVTMsp1
Fu2DCLZVwT93MgALGUiBQcHJ74lN2QwVzXqbABu9Z3D9mZ4mr6A0Er6q/v3VHC+7
ttuD7+Kllvn7v6tivH76v2O2c9CJxL0SuESe8z9uTQg57gsXH3Bx4knXYprrozQ4
PRYSstVNaL/Yv09Lm+6DuSjYt46YUryUk/NShoWshzAAeQdqVbUWjByU4vJ+3n2C
h+WbVLLMakI1KN75m1nli41Th76o4PskA0R7ZI9FL5Otmrs9Fr0EoSekl6nNwOfo
e9Q5Pl1BrAOYItOSybjs6q8MizRNMh/c+bUGYkU8w1GNwYh4myr9Jjhc2VLsvWSd
BGg1Ib4ep1uftiDzTb/jUFZmVZ3gy2es/P6rFOFFx+3KE3JJa9Z5De+sJB7FgXZO
7lrmGkrD67YIAzxGxqUSqpBoQUAReKNm9OeLJIDvOiJWscoDEP0fOMmfk9IiL0YU
k9AsqYNcoM5Q6BHQ67Z7Q6CFCReUCNxqCwG2lOm+6S5xRe5/m8g8EjNRlCNAO2iA
FCkv5X/g8IL2YAry9nz1qZIv/jJ97uX5EpHNcerVNy4CS7vyCretpA+7HSouSZ1L
N15EGsnzcqYl80VFq1BkdjR9xCJeMg/nM9EqHD6eSClbl0gjFKiYKwahQUK79IFw
dktfMhgHvsjxAc9ov7Cj6DefTgbC0LGBxWd334YEURjsFnz0X3EpazaTUJ80ma4k
NKVZ05PfDBcePN/ZLAjf9CqXslEFmSJwZ6AUz/k1cjHGG8gqolMnlS3QhmW/+CRO
mhL2kbgR/pOrjqzulSoaugTVC5lqs8Qj9GIf83LeZKEez4W4eB+ildxebxCS66oy
dH4SRBuRupd3KTCUFVkNKIHgxH6JJl3xXbA9RR6G/aNUU4PkrqEVy36IqL86M5t3
S3TR8ymOfolXKR7qIQ9nsGRjx7id+4ib47XMJQGhJevembZD+RO3FT+FMjTDZkL0
8LSurxNfS4TRi4+Uu6TcjF3WjouDdmYK7kYHjDBR9RX4XMn9r2Sw9KV9UK+kRQ/q
wun7VMvI7VsgWSC5b9xzMKAKrFKpO7N2lLrR3sRhDWAEGaSRdh4FBDsDzNpd4OV9
GchLONoNBkCMEo72Q/vQ5cURgaGB+C5uM4gqRq7zNsn4o2rzRozWquHSU6SvGLFR
uN52XdTYMDuZfyYPBfyC1l251XELI++HjhVjf237G1DSDt0iX+RigD7l4TE3V0t5
d5MhF7D6G0+HIIlrALR1iJoZRkj7gOjlEuItjLQRD5MnlMQYj4XJDUtAjFGr0GPC
JTGV5NfsHsQAGvKsjhyinOE+++TKqgcpNeuTLjVmrc4iMnfpUxBRv/Yh2gvRjM+A
WR9u+zd8PICpEEwGtFm9gvYzw+BGZ6zw+JcMRPIEd8MK/O1wF+fJw6CiJarP071M
+oieWnPxpNIJdMP0CUTXjGYRYFmQS2fdZaxtSH8yudzDGLe79HidHgaJIs4SxLk4
kPg3cf71/DFh+E8RTY6RUXjP69en7RfGmSp1cEwzJRW5ik/zRvSxFlns6Nyf8uaN
kkYMqIZecgBmeZdU6d5r6E7U2lQQBpqOKEZVncNqZHVIOx3NVNtTD6p9JMQlULyg
uMiJpvBHLsPdLNELVaTKmbg0Mo10I7JgMZRgdesP6zkhG6wXD2Ry4DRF8Liib6ZE
pG8P3sTzMbvj8VZrnuWjRvJgRVybU09hQOPymvXiprV7RSn4oNHtmKD41X7oRDpo
OBQ58wwF2DmSCNSMv+6RfzTvSe5R4TXt5xcS6ZZUGca/4wK9dlJz6DzOvNhgxvlK
koqv6Bof60etzfZOOEz/RqK/mXFB2Jx7iRv66Yyw4CDSzi4DF36hLUe7tePqkF37
jG+tqXUUXosXtiZ8Z3c3kU2qhYH1DQg2mG7nqKCqwsCQhxtpZYcckWCrUe+XNcD8
GB79Jkb68Nw33RnTU0f+cc/DhiiQHpcu//4Im/S4PV3o3KYLE7wcSRXnNkCJQjam
ZXm1WVVi8M0iTIoHISBHEiyBOxyDOeTiHndPZEKybh2CcTR3SRX4LzrlXfhnNM1x
f6DusiYhacDXucWvgDcTvid5GokvdvIWvr/BnD/vPslpW9+KyNAB1WA867MqUZEr
sSIztxy5dXHvxhxy17rQZpbDm8UIdVPSKClj4tXsquv4i1CjdYdgO0wSsVp0I4lH
WUkw4eqsdNy0nk2W4+QbcesUtMNb4lqJk5M5E4hDO5U1pcYSoek0qZn754+F68Y2
1Ak5S1Poj9tvBy++whKEsek8n/HUhzWcqmn+vqeNjV6mvBAiMMyfy1an9sPPCzlo
8q0f+sGFrkItpxokq55nGwfwc+wAcpDtHRx/snYtX+VWNvxYtmu/t6SNCcdM6q2D
I5mgOd2m2nMiYMKwFU5pzkIsn2xNTGzedYaRH+IuEE7G09fmQa3CPqkKfl82jSSZ
s82JsferUMV3M5IoXUgSsWp1lZ8+rwuZ1Jjh7Anf37VOpMQFBUwBsabte7oHeL7P
OLyoCs3MGksCTRG8QRjDoW+LutOLdjX3gXkMvWFixmSlc4LPSB8+bHiYxe67FBHw
NM8Ut5egizXkGgNAPozi0TUlAnjDpYSwUkgPMR+33zuzwU7RvNa01Fktof3eYlsu
oBCRDXbvAOBDeaaKwLu9vRQbBNuuu1vGZfEJavPGCTGkyedA3ymBlQal3veUmn1w
N+x5XrTAa6VcZ1DeEM+Zi8rJtdROYibh7DrykBL3qOL42uqFp+l2gkvNvlkwbqAp
qGiZavKIRJcuC8e1zPo3yxdWhRr+FSP/xTszC1XaSmd4WVEVbSBCaaPK5fq1SEq+
U0N/swSNKfH4hPkhIiBATLPrJR6Z32J4BPWtSXCHcsy83QQuFHrhiOMQN77np5+3
wykKSKlVKd4CvoX7biauEtRdHfvnBChWCkEjNVmrh94+8fD9RA59xD8tyk1ree2S
eGZvk9VDGU6bKfAWhKKaUWoQotKRm80R4kcrnZ6+Bh0vQkhlSTLYFb23IEwQEma0
YEFIzuAwBnDaoQvlveUKQYlECtyGgcJOfri2Cg/roPGqNVlfM5LhujsCS+rQ9Zbk
E9VbDOym0i63w1kY7m+yphmvf0Exl8E+xPptABx5d10Xi1nJKfH+PHXFrTZK29nL
ThZyD73RlTkUyWBVyZDvPR9f5FwMTVwPYhFWuQKaDfEMbW+l2OWjwaLvXbStszIe
s/K1ailCrrrIwsIJ4/bdVP8Q58wlIa6H1GG6G7tobUaEpFS00PRhtLsBQnNpKGjG
kmmpu1F11GuLjH5cnl3tdu7o20oRlYWuk3mAfBcfxp+Nqp2nb0hYuUEp5EyOPx96
gTzyHDQPIr7g8JWQzy5HtjdWTGOJWmD4QCmjZh3F4hw8REMDJ1EImFgU0Q4lx3rh
XZYCZj7jmWE1iRBVI3ByymWU2ZBBfghcfbG32AWsSn4v8JgxGwF6e/M0C9tj7vQT
G0l5pa39kF2AsrMSLmuN+Tcc9j6MoIUoX5Q8rNwxSiiHI5SEAxfta0nPblOa+sbB
tohWQ+G0NxCetFBPce7CNqQeybY9Gu4NGJa1YgYHfklYMwxBGrcWqS2+EijAZUU7
kLITo5eU4HFYdEvVhLuK0JqsyGufYnWmDpHe0BB8Ld8SgQokS1arTJF4Pva6LMuB
+Y0G7puGg6pN2fTxSPahb1WccYy2LoCFTTMz4oSr/c+wATTLHKIlmT48xmlObwYX
kM+TCPgkQv5SUqNFqqNamgzOMHQyKHCah0LW+SrSY6B2Ds/HMVegvi9dSCn9Qx43
Zf8Oav4Pg0ICGDjg6plTbehCBc90MONIhShoI9qNi02jGPocumGlCttcaJKt6kNj
e2kSoSj9kQpNVjPhrG2ibX/YRsrIQv9GfJpyrkbyxiznG3zubXPt3SweuVEm9pZY
sFuR7muQPUUXCvtDw2nlYZK6bRRDX5wP7pujmtdmFXPxRbhNNZO6g7hepzYHiHst
wrB4NiF2ILBE/pUeMDBcY23ylRBk8InmyVcjM6frYdXkRBxAxger+OW04uIB0RVN
QlQzMl0z1WX+W/OviNdFySxWGyYJl49MXAj6b25XOSOe1DkxbkCbGqJJz2JRL0pl
EGjKaX7EoG7+yhjkurzq70DPXgUFx2QU5U8u1FkY7dnTuRjXnEZMi61ahqkloywf
eMh43VkMyTBayFs/vVFJg5rRpW70QiQxZo518dRefThmj3SWxtejvRQYXaNU/5um
bvGaVRXebZsDz4Jb07G7HeksGi3tyANj+TYFeOoIakz5zlJg2NKyN5ZNo+mFwKRk
hHCLRSKPbMvj5gvT/YnRYOWYKQhaaLFunjihqsGy6dZ1+U91+Nd+S+isEmEJUDwL
R2A/39ZH+Qbf/XXEgUbtaclh6GOyeOKRNsjFxTuGJDbD/VeBRxZ2iIptCrS46Rxi
b+f0pwkHj0lhUOKK4qrNZoOsFucFQ9dKEft+irPgBhe76gzc0XI1zsR1O35NK+8p
LSCslmnj9WFWP+4YMCkeoqmw3H9C+ucdtK8f80E0Cf3OZg6HH7JcMOytnx8YvRav
WYpmEUj9FcSAoyM2+1kkdp4G2Pt3n4USOChquN2WFRIIJY9yKwEZ7FMBSLZxA6q4
KzutsQgBBJ/QqLyilP8nzcTeCn3fQixGvD2S8hqVKq65acSIWeMphQhjxslhWEFT
GERMtMVaLtRfaSaG/hNKSJ1lewJzANtPwYyN7GG27DHjyevfF8RXyg//3jNIVJMM
otvs0THwk+UGRzNrHRQ6Ui7lZ6iu1CyCY2/Y97lopzZmxZDL0b98SpzZuKCPsYpW
g/TvYM3uTxNXOWkOtI4viAn0TnS7Whj61frVuntTlmUuYXsUvzUYfH7shAtVOHW2
z6Xd9PbPSjdiqVKOxTmoBmi8mvxoMJVMWp1khc9SH00E2gr+ww/bro69AXZwzJzs
WrmQJtoRACpSKGC0DX/LyV3GXymr3pZD1m5qplaBFDAeLfgWaYDIIEzOrUP3nKDf
0mk5dVEQT6cA+lmBQFRynQPBYfKgKZh4e9AhqAHnxdOO9bCgmF/YN3aKJ+1xEstM
8ilP41zntv/OGPAuN1soCRYgiUHThOaIdQBgacpNLj3FZDdKfddCJBEJz2i8eli5
zLGY2O+ih0x7l4fp47J1O+ceQf9TqGVInZ1xIfMcuduonzp+R3o0cBhBdZ/iUKQ1
uLe1m7Go6RttLwN8f3wK3gMAi4hGYEx9lThsNNtAowH/y9R+sCyp6RbTIqkEVZb5
CXPwQ8zE8GfWPf1vEIHI2UcYERZfbKZz+UluoRx1bakzr9bobww6FDxb4W6YCYVr
jq6jTLaykhwhTjiTk5BAd9dTe7+a4MpYz6m5bTG2zdnr+3xpHqX6E88eFg8zt6Eh
A4b3AqwaWvcwctS9az6kZ7iffEXh3zotno6Fo9DjJGw9jzlOvYdDzIkBsfPcAOif
LpxMU57e3mYYCIE6WumCWzJSW/Odt8oosMQ8if31vx3Brm+zikmqSndncsEi5uSD
cbQUs7ZHUibV9B2XsB/qfy91RwX3nVF32ZbVhrVqbpTYyzeLzp6JCN6qspxlw2OC
Z8SO2b3DBUBzZafAwfSw8lhxv6dbaxiTxijMHgsH/gG5bqh/xvHDctzuWaEFFsqh
RTgeDWgXjRjXiknzCS994YNQKnO3GGFo5qV7Jesde1NCeHzAt0hRaI1k9zaocKa1
FR9TSIT+8jL+Is9b0ROug/OH9/xrn88ltSVI4Wb8r3DMqmxar81Abnel4dxKwyrf
WlZywt4Dd0ZRVdH/77TbJw2JI+/MzWnv44KQ7Latvegd4Aid02ATxbUX2EKamWon
dlvhleYjxg3l9+u5ZRWtN3P4xXseHpVTUqNFUSrghbMxXN8eENOfiK7p9Z0AuJPO
HGVUx0cAK0MlKW04rkoJAcRfRntHzmsSP9b1sAUaV22lMdBphgcKAz/HPozaU4N7
a0Lf/IYJOeLn0bRAUPqmLkrIoGLdBGGu6TWPJXGi7R/yfkBEZFdQD6LoutWafDQp
vDLm9DCTwkBWCmZ2iCc9v0EZtsbSgGT5iqEEVjrX9eu2QkZN/1yTe/4lvVcpVR+e
QwIlnf7V/Npj+eCwuLt83KcOBjiX1Bt0rO1AM8vdcRXtKDVyHMIwzHGVIwqAy4lR
+wBrWyMU+XK6CIBRn6Fyan51sf9Ta94F1G8taEKwl5uCjSQmODHXLRvuOfp2oI0i
KqMOrZKnNQkQvYDfInlq9RPkuF5+eWARPl0H8Ks7sqL28FO4afn0ZjZBFUBMLWFt
+ur+28SqoufzfW9R8E1KK4SAkNf0PRDYgE7ChCThbVd6RZy8Um/iqpyiykVsw0xs
ZjEjOZ2yEEUY/u9P2gbxzEXXlsqs3/YdMgrOaK2J/x6XCFotATLpJQ89Lu/X+tuo
BoVmESq7xvitbIy/zH6bPqTnOtoyGoc5+HLy6ns/hE+kbcPff8/kjzUOO9y9pLOa
LotxfkVhDILYoTZGPfCXePTRU7mOfz3LDarLE16WLM8i7KBRT1BpwFxak2MMCSUB
iLCvORohvvs2nbdjl6JgHdyn74deDwXnHMhcwwA9DQW2cIGoyFcJAJE/OVSS+QE9
a6K2/W4lPqdD5ES5Y2AZpaPlGh8R/3BHKADQlE8qUnhD+DG+ptvb3XvyKeYc8Fe+
tmvj2jSaNnDfPCBo3rrqo0I3RNiDAYoo/qajwwyb73zxYPK4RJDuhMO0okwoclMd
DoMO8vcgtNA1jXN3Uhz9+ChO6VGZPmx0znrnKB+VaslSBg14ryhIq6AEIgNbbVDw
t+PxdMJFJCTdIWx8Q+lG9wKNW1j8Pg6d7GdAACRH6jGqYWHaiFEi9rKl91xPzPhN
gu5FksN8PUPlPRVlXiFgKLKBBgY/dL0NiX2/QKoFiTF3XJ6C4XQJNh36yw9JA9n8
Jh96i3x1e/h7sjZXfC+suOtCMqEvvr5Pa+ZmC+Jx12fYxImk9SQJpuDcfsDv1YYZ
Dl0CahJOWo9506lOP+flw5rWRhuNIC3BaVwkQ4Ew+1eZS2Tu/CMrUYySm/MX6cco
VnBMRtKNj9MR/vxarF2uebog7yTC+ktz1q2WpTG8N1iwKZndfQwQgagLkyWLB2Kp
lZA3u9GOOt4No/T3GAdrCsjSV0+xTTaI/ZkWBp44Aphlxjwcv+claOgmBedg1QWA
ZNUNbz45G96/Hqqi6+AGHEsNnqDzGS/glZHOuWXZvE5yT1FxwCzRq4jvGmM4ge2Z
9hzMxU7F7TY/6MRhPShyMRWMon+2l0F+iwMGvY9E6L/4gm//l9EXEaTCUcEVN9qu
oAMWFjQHEZllobQzab+m6cle9i3vOFVZazNw+kyYbgIT49OpHuf3FzNx73DHZ84h
DRNxcOqwsh+zz0ZLV+4GOp9B2adzyL36TOSPpbHXT3MTRXbKMO0Qod+klhMU8kbg
mQkRKZV/aAkjTW3cJy2ot8CzJ823KtAjJ2UiHxYw9um6PDho2TgDpqWttANtyuk0
j8XAbtsymmifcBJQDZtBZZVisndN7UTsyUqegOeDZGojf0vy9vp3afHryMVJp2R7
PwlUYPBB5C2OZWwYVDj3vPkCAM/pdyCYwTqGHG4xVc7EWMYka9n/y1NOederVgGU
rEeGrsdk0zPO3y/MboIiSI8r6/adTt2NfEklJQzg2vEmn311HKsWGOOwReR405G7
koOps0wn7b0ZE9IBFPKVp6/Or8XJIEqhZauCMVLnE7kdSRb2wnpcDVK3TsC717lQ
kCuUVqAU0r8qE8FQj1Db/ztRGepmYUxqyKX/vFtiNZ+lYPR0J7C7rAzwJVxKNs6s
eJaTmFYAoUchEb0RkctKvQ3ScLDrU+S+iYixaE7KfoojpGZsqW3L63Qg4AKtxNTd
DC/vue++TgQGaXrIAbrTSNSsjVSRMQAMy+s58HWa28eLAIj2OyLzQnSk1mshCO4c
sqdnvPdD+NyNEBRe8rjNHaTPjyXC+UUwSKNOz0esEdxWy0bFI5XOQiEJkQCCffZq
FEPDRpwQpV52rNQPxlxP+miDgzED7Von+N1G1e3vT2f7r9BkQVqDGFcib7/5RB3y
9oCZUzmYSrM/WWBoz9NByYFbu36/A6U+wExydf+sxeQ8p7fSKErfOMSWxFGStYrB
IBMTB4JApnLQD2zvX5dSXYY8toshqgHToQg1WzZq08Na2Va6RFWZwPTxmzA8cWgk
YxVZncTcOOt6lSPuULbuL6kyGcE4TgAeNPs9IfKClKFr1uxc4Jv0cNiT5G+CkXky
dd3e2b96FdPy7luFZMVznj1BO1kbtaBUc16aYuWcTkrc5cpmlyzwZnDL9/FmeZmd
Ys9qQR6d5APUsSJMVlk+Bn6oM12N0lzMRaZBtlqE5JvOczcwTObSZjTBTz6MlAHf
4xXk7+1Mt/KTehKSuKmAqhskQlbys6n3AwMq6e9c+/N5c9CLKTNkPj+txbqqdrTa
/vYa8KH4S8JoLQcp+LCxV09dG6xhT+YB8BkRX2dTKrG2SBQO9HN8/mxsndza4izo
zsg5SU6BzrnS78c3oXOzLv7bYffVZewF6F4MOED3Eainpv7TeDVaQK8Yvp6pVTWd
Y1Su/y2AdMOa3oJCeRqxaph31CngWdLmq7fzVmhd9Vo3lNeAjOqSzMEoik56JVkV
VQ96tBaBGc8OjLvdlyAKLfhDu9nDx0EJ86mPOWAcn9F6NWVDulu+CKb3XNQM6t/p
vl/8psNkfUtAm5mxAPVbYQGk+u/IbZxwjlSUyWh4zsjp4gloNXFocSA8Jreys16o
W6lf1ejk6W/b8iNE2CcnYBVtDtXf3pts2PFBSACLNk5jg4cbIITLLqL0P2sBILc5
E78oS4Bj2GgdF95A6usNf6kPRDoQOF8xIAW+ks2AY1B4gh7MEFw2iKgfViv6qD+c
+yItH004Aef2h3pC0BXbeS2o9aCDdFFa2DRBV8sg2ZswDsisq0Fv+Gv6t/D6GuFS
009oWUifon/riUWX/oAdL/1GREYyyiz5gd33ygqb2lZ0X9grJ8Jb6KsLZaObf5i2
jM8pqmMSUx5wP3IX/tKIhfeLqIesgrl/kftp821O51iYJf8mZ5B/J9VR2WPAGoVG
0duA1tXvqsS64MIySzZDESE8q3qtk1/pc4AJzkrEw/xvUJzmFFDcw4dpGsMCNwxs
IC99VlJLizr0+hmrA2jChTSUL+ItCucnFTSkwCio/ZZ2QiFJ4Jyai9BiHF31AwAQ
pZbNalf6ZInFtL3BgBXgboEyUUp6lWv1eZqug6xhbwNfSextwmf6kriRbYtetbcv
WHxWY9hcJTC46EFQdH3PyockRrLkNdVmVFiNRT9VHvQ79Z+1X7pp3a1LE5HdhQi9
erCK2hEiy5n8fdM0MCXIYOhAYX8F/uDNEydyWrYSQOgEjnI12UTtJ/IGNE0Pv4gl
/QvBunvyvJJKeLD9XGy1maRlzGY/fFhSnuYk5QGMXrLBDI62NLSbFtgk/mLcxRTA
wgv9p0K8yynWQWvdpiUDPepUr4rB2+2msAX9dDsn+zGj1YccU3dwXxnHcfsQybbK
OoveByNMdJUz4buaqnLtmKtLs68QI5X/f4ecvexPBxfBqsDZOfzUD/zV/OJCjCXg
9kAejJuTk+iXyiqUM6HTocv7/rFf0aY8N+tKo+d81l2W9T3D77DWrOBiW6wh5+Cz
l9rAsG3alEteEWF0At0iozVGGgX0a7rnRITujBFm5DzqDPO+7y/H9cyUrU2wHfDR
qxt7C7iQlVcklgq1TUNwV3TaMVGlaK5112dhYTNktQodYG4+qyoTqM1OWPsgpI9b
dTW5LOFhGSOfbpUoTj1HRDrgLqXbXN1kfj5gzTjEf5BxhruZ8dzRgSsugKI+F5kG
hGEpY8T0hUuw+PkF4hkg+lOgUohhHdnanKAdc/TWKCyD2eEuQ4ws+msagxqF0r52
nwFW9MuJuj0BXJRFdF1owUFMyY9H8mAXGtq36LqrMgbDo/x1OdiXeX0GOG45ccbG
WBHFnEU3CB2RN3LOB0ygNFLq/2d3mE4KP0N9bnHQexDb4Mi+iuW6UHEapERAyRsw
kJkLOX9xtI61ZG352DbM9+ieXDdhuz7d8ZQmP0YNTMfr19Na5fKVgSeRRGzuNeDX
NkYK7FcTwRx9TNo71iyMlnzeusab+hrcDcuMDu35tTl8eRr1OlDhfHKplXlATSFK
SkFQKUz4q3BDN45s7j8BKMLo0Zdamqs7yz+6LKiuDR8jhhZSU7lg+8pFakEUWcJR
eGwKJM7Skb+Aes2k6Y6Kn6QwO5NUQcbP66nI4HOwpUK27FlxaaPWLrzxkqKysDMX
2N2xhf6yA5EnCNRL36EhBYZqKUUgya0mXoE0zxc0Lzhmtf5QPGAp7b3mAEIX0GzN
GeChrzkim0VBeSI/w+3QviLkRoWvzqK1RuWP8Ejtw2HfKuA8p5udp+lYspxJrk9F
NKi4BO+ATU5Z955ugbSeESOUsNI4L+OLBm5SMdgByvYNA8SQts4ebR7SNe5sY+um
vzqgFdFlzk+e6NkJyUx4AjOEVAIil/5UCPr6PXgxTplH1CSOP/A4+WEmFcTQsyu3
MfaM3IvxDZ6W2Kqvf6CBeiW35uCapKpwN5NcCncjrWPEWNy172e+XuTfkpxKnxQ3
NDw5mHcaY1MvK4vNpIEFgWAqerY5uuB0Lc0IwsJRzVe7AyzTsAP8ziVrKiYZcF3G
oVfdelYuUqwGqZ2E3e2UyaiZspjrFgjTnPOG7su3NKh0pRh144fGiGSRhLODBm3W
s4PeGQT65c7UPBspt3uTcapquL/Tx/5+GsaMECLWnIGV4gltr6i1HkHTYEs2FwMs
kE5HjNw62/o3M+3zwUxWaLawTVD8R8b4ZOwEa0znwWa9c6DMItaYF7vb+7fRmI8x
BitLGWIhgldPZ6xqGGVJ11xp893OPzGWGXHH39EgnbAlUR2qNXJedlwbmSC0FCj9
qd4P9JQMlUzgZBhaEbIQRz7ZvaGjbLKKhVhI5AnK9Xd5E+1IkPiRMW+u35ykyro6
+uypIvxK4Wi667WEqv/ABj45sCK/h61LWg3jUXakJLrBDSMs3KXDw7dc1tVrZvRX
EweJM0o7ke8WMmIW4vlfAhSnl8wqnHm8dwKuyA0qG4frCovFvtRrziGCqPSBUajO
5b2Qf+9iCO5kfsTJjRWbh0rlNdyl4OZnHRfJkmRxL+c8otGkrOaIWKvj7TsEL4US
ZrtsKk1Pr/S0M+3Gm8Z58N6Ei6y/kCjbzTTMKhpp4L/j+q1mPGqA29yYfWrUAq+H
iuiAWUc08lw0j4KYomI7/2mO3gZeXWolMiqC9s4zAmAOLzZ/n2WkRLqqiX3YmbMU
oD/QtjUtv63Cq1udydD9+U9J6SE+9Ere+9VE2T4MbjH+MK3o0T5uObSU2bkOLG77
NCBrRbV16cjyj2CzLAHSL5aSYHJX5nNN3J4sPzGAKdO5vHD/sY24w7fQHgCDukKt
pFnDq+GT8iyLbnBJsHvySNBV8ClZjQ/rukTTAb3I7MDewUXpO2QTxQ8kdJe4gEP4
BXk3pOkt8yf+S4KJ1zlDeCZngTwZJ3Gd0pGdQ4s/nbmdfhvNcVOWoOS+UT4Bh7g3
fZGlYl8zm1mLtt7iPeHUp6G1dM9gBLbr7v5pfFlo54G6nUQWHqf4Jnob5UhDldoo
nrkfyu1M/qqKBVjt7dnAGwdjVCx8usgJH0VrUJA8I6SeLKomiJ9JtVyPNu3KIQDe
+LCjTBTlSbMo3pU035Y6J/aMdTLaTyqAIP8Rwqx7iNg+11S9xkAtMhQ/dQmuM5EJ
JYAySbF5tSAkSEEg/C6eYej98gESd0UMBhEuw7gcwjGXNglWyw+nlJhyl1vuTlqs
WjJ73a7sBA6K2gHMVrEHHISQEOR3RJZCF2L0Bd9r28aYZENCZPpLcS0YEoR2jA3R
bSkGg5Ctd9zljeP2Cap6nSLanqifa2vh+/UCiZyLpb7Gnrm5Af/wMHu061YzPYpe
+eZjHRcFsufhlLk3q+at5zSl4fX1j+YIm9MBv0q8tT/skdy1cjms/3NLSNp+IUuO
eqFAiprBJ7MzoAeqSCplRoepUs6qNmIg5LsXC90wIjGp5z5U4aicvSwLm1uoA3Cw
vxVr3JIZnuI+Tw9NOHOJK6M+Wp1BCXd0jTFEX67cIL7cyA22VQaWhf2kF76T4r98
M3gzRUgu75KMdDobV5LRfVqkFJvh4hHzPMTv9wkVZzKyxNpuRP0rleugO8FmJS4k
/tAV5wWk7H7lIr/szM87E61XDk1XVyf0cqI00XzDMlm6yB3aTwxj874XvQ99VO45
Aku6KwMz1phJBQOfI83yB2wzVMSTPZ/LrD616tXvrDx4xL0vQvYk7UY7Lyh+V8KY
BJUpdW4RB3hRPEuh1uUsPiaE/QlvFitT1lR8Gw4+yvaLJdcX1dM1OtwBNn61C07W
NxIfX1UPCAiPz6wiipm8rei96n0uqFYgSQKGVvohvah+j3vXPZzZKQkr9COEX/sy
lMrb1AdFhan1dVjBG0/OZfRrFoCGHy/cyob0fZVg52zUyy97pWP7xbHisReItbCI
lpCHC3HZNzDxpe2BJ60sySiNbDdiMSOy+X1wzgJ676YPlFNUhP/ydPnbr1CW4sX9
wcq4XxkuCBOx2pCwS5KUTgcMUxmCSuHK0TtJGUtQu71sCVnoigjZRSxwLFuTLTGu
dMzMZILy17iafJSMqvyAhnkDOoChy5En+GGojtgESlgLJ5xTGOftmpVdF+JJOXZE
BEhkk9F7UubacBfOutPt5VbDxKStfUykXTaFcqQyr8MuFRSE1BO8+EzyLheEYmQT
XxABUBmjsMZ7+4gxRLVtGH1BYOqhuG0+dzonX+kPI34NbGxupz/Vy1acfNUh2uCn
DAfhQD9oKqDElNs8Tcrun60CbhnbmP4izJdX40zTzhdv1Y2kymqYVnM9+bGLdb79
5a1ehPS3XDQKcgFJPg62G0hxV++Ift94vUc6bydegSgYBVNO2LW8eQa8rgbZu+ow
jNFYJhmwd7lgalrWEoNDeVoOOk6iYg0AVjXcHdyN3Sdt+tA+ribu8Y7A6E7wcU5l
ZKvZfvQSx+l7UhafKBmqMv4yoh0LioZJqDGw2qzJUW0RewfaPSISNha7V6o1rnIR
epnRt07FGMWFKpXw8SitO5rzhEPs4baOsanN/EUorucMhWlLMzhlkK4BtIrlZETT
0C5PGtZ5wfiI0uyNoD9XT93BdDnqMHvygBJsZIGj6xDlsaXfll9P9nBMWW1OKUsA
fDMZpXPO7niaroqQKLQ9W7EFUmwfVLr/+xZRxsJZmF6+kZSizqRGIAZHyol6r5rO
+bdh7x3P8xZYrAiWEAB8aRmopmPwcl7GdbJhjM5T/RSGkq4S0IoX6ms0zc08qsfy
wQ/+t8CaSAZjKLELDBBRkxHbxjpTAX6Ob1K9H/nIsRNuzweYmR//A62dNHG7Z8gX
djyjLNS8XnGhX2alnp2Q8BeO8WIWa2Oqn8WJuJhHuCvVFJQYXY6t+edAsoa9mrFi
fjMTdrPhjTH+aPP6DH1XKFbVRRRT/RWgZ7/QH6MkEuPOcCkn5uZq7Kyx2ndccYQO
wyBsAdHVlT3UNQoKLg4dGAhI+YQeBxqYj7wnLDUfFuDdlzgG+ElD7dlmjigHBcLs
LehaaaoccPKIYY0Lu2SMbhaLOcbUBAeMrEpmYauRgpmyNpsZYDoycQxw0Sew79vo
L/SRv85U26sMylcV6jU5hRqeydYSW8S8YK5AizjW7y7XCtHyN06ekk8E7d5sfmZ+
oNjyUuLg58UqKTlcRZGaBI/UgIKEF1y/REm5XKdCdfv43rDJh+PI0TNMTk7S+J3R
R4OWQeEgWTsmGDi6XZp8iS9/F/dZgHCMeITG/ho/rlXLDc2IbyNehLxzMlgtxpsC
0buXQ1s/+Jab4TJsnowj2Vkb6ad0hw/ghDiAHHjX+ODUrbdguNlbKzOjWP3n20mZ
j9/bgmp9GR9u615t8EqQxXCEqojAqrqUm9fZOv8GaiXx20zXsYJPKIbJi2R7tBow
1dwObgb92tW4LPtmzq6v8W5FNnRVm1cD7qIF9A3m5B1KDgXwxHY9fqYbDXHjD2LZ
/wIW4TtNBQiR41SnAGVGoeHW6uPVK0M4xIiR6wjMsMO0yY0LT1nyTJi2QIGSocmm
NxaqmbW+xJAXhYuZIR/nwplWcKI+VpDBjjzN+bSR8KEYP4hCUBVVmfquzYUFW/IZ
C+wRmQOfIocwUNwISDHUOzp1s79Ii9P/zPCHczM7LotAFLIq5VCmBVak96n2aDNF
YurVxp2AKhdawwcGaLapZNJ+VrskVv5qgT/sr3D0U6XewERgyrc1BahWpG+3sF+c
ZYWltj1vYrm8gxcjPQ8UfwXUDVn0yN/6zm40/vvKCtWMqQJmT328oHOyB34cJ6XH
9lRNKHSlLLxSPeYrnQBYiHQrPTusmOL3bXbKhAzSecx79OQc1qGDqXAZcMDDFo+8
b5I6x6ei/aWvTrOk2MCqj4oDzhFTSgayU3kLx+IEIw7RhCCTWvrjt3dhljEu40Vk
jk0+EeH4KrQBBjKv1xzV11ACOtwCwkBEFFlCuAcxKo0tKLGSnott3h93sKT58AdR
RAt4GtuoieGjSpVBg7TXVnopkcSIojxtpXUXz/RGnyofww6HIbNTBUpIRQXGLsEo
bOPgV+beeN4/U79ZhyvBCxBXL6cGwuSjSd9Plm3UT+7xi6IWMRieDOtip4kdaj/R
mT2LFDO3e6v5JT2JdQuM1tNzuzqmw8e2ec7NYzfCajTC2DO48bcov1OGmSVjr0fL
yQykquGhiCeLd0P3lo6dGvylViwNMAbKoUzy+jIHLc6LU3TrQJ6UqwH34r6UiVk/
1km40byg1NSY3te/OzXkn9gZ4KKcnrZwz/f4AO4Ap5EGPd/3l05s9M0z6ni7eh4z
hAm+l1Wm69/1KwCWKfGNtvqj3IALM1gS+l0rrBmgLC0l6HpY7fBK8NEwU6TFooL6
2eD1bqGbcb5xsy4eNtb/8V5doczFVmpSRkPZVuNmunB180UvKUd5iGBz9HCEEZf9
EbuteMUhtyZLXGxx4U4pucw8MHWSAq6d8jJlIgbGbiqI5XrhHY5/diU/iccBY6u0
TQLZNXkDOKJDPcORYWnqyn9zIWcV/oZ0Y0dlTWzhks0Eh65U1ZMsDKjHR/tbNE2/
cAzGH0j9PyqqR0qUOZbS1Qu7PNQcZ3ZLgtfGoiQF8iv5tLw9pWWpbvudeNLG97XP
GRQ2zBRFwK2a5/uTrxL8OjVPYDAnONXfX00r6vob668f61sZK5ZVXjPz5jGoEB7o
4zas0cKFX1eWbr+JKJuc5rt35XEUk+aKuR279sioxz7KcfBu9Rdisbir+lWiTsMm
ITtfvSTqhWMPHvbiEvAFLqrVA1PCzuaKwBV9Zpj1Y9tQzYM6ogT7Wd+WxQhHFMtV
f7n4WNVKu9CdnqUrJriWaDuq9cPv4jAllJIV0JAS8dBdsKB5EJ4qtaK6sGd5rbhn
mvh5a6FRLBVZ9Js71b3BYgi3aDhaQoXhTs20OSM0+OA1RnDtIOT/VfNpsxubeQPO
yzDBKAtp1QoM6tU3o3cOwXgVV/P0GMk/dP/DYc+W/gtFb4HCTKBIG8TeFrDvGS9W
wBeR8V8FfoByjEIqyTIScckRXnsuQAKRx1M9h1hamgJim6jPd4fYnGI229TvD5SW
7DlPuxTRs+2af3jCAabACvfEGREJ4aliOxm9iIn2uVwdgm4oH5F4YAABz6/m+HsM
uhYE0qr2uJz7VyNqXqAxvYKTKwDhfQZzvBEPzXB4P5DTgwc/J/z0GUzRnmYCJ+4d
+JJgHW0dEO4u05QaNWmap882Q/6Eo6IdQ/4W+sjX9bctrQABDUu7cCdSGzGxJyVh
GBW7zwd2VD+eZ/f4eTBTzsPOuV/trcc/NdiiYArJpdVKpoMUd0kFBe2yx4y1fjTo
a92jGB0s+WVMQhzAT/uv79NLPjdQeHN72XaSQHpBsAYutYkmhlK0ZR2Hm4kB+zbP
aLC/Rni5iLQYOkJkVluxPbdyQg2KxdHqcIbdBJjNsQ/W9qF+7kSb56as/cek7rOy
1Ft+v98ry9zkapV0xpXeyF5R6kOcOJUrC8A2YkAEZdWq13Jhvc+8lEoKFyodAM/m
64R1zggo1VN9Dtx7aXzzp8zs1fnwSRkxGD3m6xxPC9jKrp1Delh5cGGrwv7PHwRq
0vJ65z3T/dRPMPvD1nEoKMeK8Vs4HvqDJG1n8OPRqPqRgLGYbYeEgeaLwoDVEQRz
raKqJTtjmGhqG69eOV+VdDC2toYMoLCsSS0mVMiuByT0ZQYnkh7HXfgh3fTCCxA7
RONkjMqackfq/3eWJTCKPd0m3qLfLdwQLRG1bKib3sIcGFdEKyFpVBCMFfc52int
BGuNFfGl4UGIcMUX/G9W7yNsq5Ck78iE6JX78dbcE4rjUhOzp9HB84VTKRivFRui
8R+QB+Vwh/Wln5UM6PsaJXqYXIhQxYtjxEQiEqe6hSrGb0+pnUkXgkCr1UPkpyJJ
B9FPM3T29+kXUntEwoaRmG6TRCyYvJVXavTWo7oZUD+6DRjgL7pCd3SZYCIEaR5V
DNoIGRdlE1NhqKsaL6TihX+O/WCjvCMZajSMNAlCSlXtT6pAOnI/2d2v30UHlzcK
Onr7iMPSWnpljbxrU/piyXlSyeq+dtz0oKmAspugfI2kEdu7EfufqGy1HT0ksHuW
EiU4bGqm7ItwxkvILKUxfMH23AdUSOZ9awiPoVvCIZ6d37kosNsGfWYVmFdHdc0Q
IJ8L3TSl7tiERsRTKbvw59Aq2P44Gv25352NxfKq3SZNWK2SmP+KyxaiOmbApeER
dRVkXwCHe1NxWVN6Bbu9e8VBnE8VXtTtG0waAE5mIU0HyP3Jazepz7vzMg9dqgPD
+k/RUrPCM/LF4mYVFiRp7Wh5SlfA8aHZv4O9zz6AV0PAdlgeG2eBV4he94cEW/ct
wXaIa4K/sl+2mtSkO9BcvwOnd8Emk/wxpe7kJObBhBjxq9YSoSV9j2pbSjKYdVDz
qkFEF+Xmfpcw7YhtSC/Qh3uKkiwVH6gcEaDUS9pbWalsRPxn6HmM0KJfcV6h92cq
SYwjqsZooKFsryXiOIAccSqr0aOr9pPOPv82LomYySplZIt1kg4GMKWzhpx1+gJF
gTo03Pit5fEQCYiZqB5xW+JRn6Lt+djqPGPCudzd9jYR7vAnU+/7ZqOnc0Jlrv0v
bBtGX1N0u2C2YL4PSSc97W3+I/Zv++pmywyvtSHfrKVq3VNCdUelkTOZKdKrs7q7
Q26KDRlx8+eWCH5GniCB/F/Zy/WacmrYZ6PDdV45Ikj40UmsRqNmQEFpHC4IkBjN
EsaboPqCOQ90kobPt/p56H7Xutb+yZvV62onao9L26augoCv/ibd/7Ux3jPI/W1q
04Vo42py1w59jTC9I6MBstFJayfY8GzkTlaT+m9VM1XZWxwlYfoQHOFDr881AfmT
tVlGDRmtu0Box6mGwmKVybeZ2sr32vigoIY6qmJVL6MhWL/WOxYFJhQxeiATr7SZ
xEfYHY2mw4222r4hjM/WqznlRj6SDusBidIopJi1wSkoNopIli5US3/DDgIYWih/
84sew9BYVHQzcHK88KUYge0PMbP2mT5VvtcLQd0CMK7B/YiZXKbJxHYaDo65bMQD
PNKdmcOIBetDSZtxp8qK9gjd3OpcagXFTO///Iuw+sTZ1r5t68+qi+sGY8kcJ7Lq
NZB4+My8ONQLCjQIFqOJinhb1ltEJu7di/l9Cn5WuArQYYKlytK3CQAitF1ZIA0B
yiXRd6SpSJXD3zhD0ZI4xNbaLH/76hawEbgrdrj6fU9T+x/r2sfxiMRUAFTjTNIg
Y7sGletY5ng9usdDNZMjfR4el+QwhoX7br8kev+PqEolgwMOYi8NuyV1PIUdNINq
Hx5arlJ3jdxUfTWRIFQ5gXo/MhPJHEv73JeE4i6ap3DVVQ/6naJ7AYFVMLZdLYlH
upV+GwVjoTI2zVeCXxo+tMQxKkLPHirrA9ZRD3jMOmRlnwV37QiLxgfJVKnm86tY
i6kr+Rn16ss34wXB5ke/8gLvouozU0y6YAFyEozfTvxnLc/N9dO2Zhbnv9GwsMIJ
lf4fCRUXCp81uOICXLPYLSkotN3LCrOjExFl/rJd+FOl9Qeu/jbHf6LSAmaA4i9m
BJGsDGlyOAVHU2itD2plKo1VgYxDDncAgIOFzSbb26ihaBvU61Do6BDQqvCBwSBG
xpN6ecMx2BpkyaY7EaEYGnCA9ycHXghff+is7warDxTVunJYeluUu4NxDuMvv54k
++sX3MB8tT2O3V3THXK1DZHEIigiM1maig7G9QuzjNXvM8/gVDqtk2MkM4J2rBA3
qH7wonkdPVi+wZNnZ16OeIgsW5xorn3v/na9OQSRkFn0GuQdKc5onT1QtNxaQx1m
o3Eiu6AjMWk/SC+xNsCi4BUfYo4rWudjlKnd/1Kg20UxTv5AK5ONkaOXKap30pTX
HdueSI6doUg+BqvCjnkjp+mPszPRbvmtGtyxEHLA14f6J+BceC9U0kcAFmVwRIGr
am8DuFvACpShS/RGa1iTg8CtQrAXaIqfZxcPob2czFie/tI8CvUSYTfFGeNwvrOv
jaWKRuKPGY/yU1XWp5R+917s+muy0l/DXi/tLZ51FXNmBmMNTB2HnBN3X2IQ0v9C
nsRT1JHib2GORyanXYKRdwoKDO3t8Cfra81m9lO+l430Spmd+gtNZN9PXhfGZlXY
5lOq8ow1J+BOz7uOP5gWP0FBjh58tybGaMlbdymhiB1iJuXSK6XmnV2g5wNG+/jW
5l0K87AvQ0nkMgjlsri30BqkfI5AZ6OwadZXTo7w0Gr7kw7poZKoCQX0YFIgB1i9
H3GSn1dd44v5LKBoHQeAcJYA9krFHjSyVlBuc8xwtWMwL05xkquXWRufbFVNqF2n
ZwwQKJQC45+actwxzQGffxv7kSQnXiKWbNXEusE5rOUnEM4otgBkYx9LHj9SdDMZ
yoh8T9bgavoaBD/AzRtpRvEuORkKdnhh93SHaJ1OYzlftvCmnOGt4KspKuiQe/27
FDOEkH55L4aJrooTw1Wk73ykJzOnM/WndNr6KJqtayuHQacKmYN1X6uAt5nvkk8u
2QEbFeqwKbiwhHYEp3mkpldwpbLTaFsmUElCBCqU0tNgAP/AOlv+RTZdgV3Sye32
vATqFwffcqA6XWXTol/fFkUjUOHJIrISDShWBBUmWZgk6WJAHNHAbmacsaLhrQqt
EOQpODf2I9/nMqs5SDRQH0YN2BV785BezgrUu/cZUHyoWzHETzn+PtZmFUFLqgVQ
HMa6fkuRnPD/v3Cl8nf1FVFgtLljXIivtk+jgzYdWSj5N7u5NXyxmVhXZLxbCWha
5zip1re0HA5kK35ZANpdM6WJtmzE7iQygWlkjUcrjH2ooFelLIwSZiuJjXzyf48K
n3H5g6abFwu6NwnWsWgTVT5ZRLsy13yWT+rDoy48GfV4OvTxVYn2YsUUpGHm6sEi
KfvrIYP2lhOLM+ZbUtgY4b6+iJwsyJbecHEFOoSXoZOQp4eafEYA0D0nQ8y1OjUO
9RInuVIV3J6rmvp4tz3tcUompcAgRWB/NgysqrWCpZ5b7bDrdhQKHqQl0EuNSuBH
zZDGMbcw4NCx6D/fIDJ92JOb0cLi+qLlFrGttOmkKJ+yJoSe5ic6mT3VAZx/aRTA
fZ2iByCOsa/c/Qy0RxXLUXl/keHWXWk2RuMHVdNHVDz0Of5j8Jlxzg0wM9UjU1aH
bK/rmfz7FPSGvpvvJdyU6nq0I58NelkeI+8nc4iEYuzPuN7MjjL4WkXEPd8eAqhh
v450TFaIxtVDNOPlCp/JHEQ/iPYqd8M+li2Ljr39cNf4DgPQCH4ahGZjRpizgyfA
mBAggaToXkqJoR3HUYQjHXbbWXGiiu1bOwg8BbacU4CpFXfQMHh2Y6TV5JN1CdsT
HRp1L+xYjmSFky/kOhsKSD6arMX3oamETod1iA5VWeepgdnZK6k0BF7uGHwXh/Z1
Q8+rj6lAU1fGN3+6qQ6fwIIg6aMGfNIlspeiUPSume7rzTa4m6p10AUAhZdA858s
YAfP36KXQbwl0mT16PA72NfeG3rj/8Bn3LquFvJSnig6r9TdAL5sVTQ4KWzs84an
kpsHwN/32Rz8kvuxF1uYfTKf2i30NGRgXe4MpAYRzHu+8fwbyXiO3UgC8I0ODrBs
0ZTzxV4r4CAf3BnB7GrstGU1MAcAr9ronNtPjzJkR/Ar+qxBA0dZmUMr59O23wPz
5hcJNDcaUEtKCGbIJmkCr+QaXsemNYpGHKfxXPbXzId/grifES+iu610gTWwLBBh
tZqJMuw/+Kj1tLLL8eQO+XXJJXqF/SU96YHKkGBtanM2EFZxFxRkg/T29/hgl3fJ
yYF8iSwwJ6kC8s7bQDtNp+uDE0D8AOJ2aKztF58qoGKDwfWIC0NbezwSro++57dU
yoPulJyyWr1dB6HWRwSrH1cnfz7PGKVPrdjoNfaRQsERLWXFzWGIdaAyJCZM1Es6
767JuFrjz+vZGBiTorhpIfvvRj5rh1/+T8EZZKw0WXhfcMs18v4ZaXkhXfXGc1zy
Fx95lWkBhyL8FHHvT0QYWUPF/ixiWHwY+2FItvqiSkd4AeZHjzS6gFKEUY0ffZ7t
wKoI+BIvPYGBqgBUJ2iqPpHkbpf/HxywuaVs6QNmIjrs5Zx6SM7AFt7zaUDY3Aop
5dsrFp0n4jnV1pIV5L+opM+NVCmUu1KjsniN8itWXJSg+6kFh2a40kNGc/xk4NQk
t2t6mVinf9I3panfancqfBVMrqPWr7K2zYgrGl5X9Z94uabbVm9BnBvpIzsNiC/D
Nh1fLZL+WZa2+rNxp+ZPqQWIgmx8mG6MBALKN/mP9G8igG6TfOqRGLAclppSP9cd
2CnOHzoPE8dYDxZoCFUBooApFsumlvSbIrEALi9PaNBN1Gse+FGm+u/JmjBChpig
9QCVaxiuIqS3ZYzibitYMCgLZlHRzalSzwsLQ7ANK/Hdt+d0idwl9qmWTK+4zijf
ONVvJ/D4fdx0449xY1QtDY4zyI51L+AWzrli/fJefS3Y8W2RP3B1PdDJG99sSjor
h9zfP97IlhhWC0pukSfi2Ik4j/RPpkaXso+b+gBMQ0H8x8zqw9BLCAgyGLZBsElQ
8RKYWnJFKcvw2e0WP21ewoW9nsBhFWKf/8RTdGbk3w7+BtHj9x4OxIprv2nijxdU
hdMqgyN33i7YIInz6ee81rkhBTlIjPVIMtSy4GnKO63IuGqwkfHWsnhk08k4yYKi
kPeQkldETMFEvmHKTcVUfzwnwPQCRtFxIKNQGjuaNpX99T/22kizfO5LdUr5ajmp
9MYyeCM1FHIum8UH1isqRGbTEtEWEu5tcXgWFY/zDzQ/7qUxlYqNw24D2HB1/TFz
VQ3obPAmn3yI1W08307XIy+30BRglmxsijZEzWwrcT7+l/9OPNcfd4VbvPKrnZao
BngAhgKr/4ODYFh/gYbTB3CheVYT3ZebotZVRagPz20PqWywU3s4WA0RcUlpnWGG
fGCP4sfH8sIOjkRMSt0uBjHWBH+Oauas1w2MZ6rTOVNkXY9PI7gNAvq5ceSMh38T
ehBY2hny14cgezRlQJUaMpUqaU2ucOXGA1ddCqQ5z4uuAKMyEbovx4nw5Sk7wOHq
9JKqOkucHBRY7/+77wCn3/MH+Hh9l/iPJSvJs+WDABe/0mIJD+OsK2CbfXR3B6uC
+gJ1CQapChMCV7zQ6uDeTQ4ctBuBuFtG7NpqLVWD6UDIQCj4LYctq3RKrmxuPJdE
6VxN5gipSzXV1+IOqnvbShCNDpNIltlg2p2Eo6ikaTVuMZ2x/w3nL80sOGiR80yt
cheoLJPea0NzKwdoHUZAgZvUlxE+SYtRA9ub+PUQI+pq9qU3pHR5k39JLuCmJVW3
W51xY2kYRpw56DKX7rjsabSGKyL9Cis5DBjTQcoVT/kTHAzIV8wM7dyS6DKo5X8r
0N57Dw6x/QP0nI3vZLaGV3BE04yHF6ZA4sWNGLBeJGEl/+2+J8XE2u2khoQLLzur
dOYFimZ1M/vsLhPAdK2wekgJtqrvj21VTFqnCMIsoXvnN6BLGbvYEDZBCiTKEY0O
b35oJUnmN7inhtNya+umLSIZyZX8kdPD3pewbrP11hrKH2u8f5n5y4mkZOBx5+Rf
qG4YQUS67iPfqNyITzTEpoqeCNI5fsbPHlrwE+VRKslgnvn6IsZtJ4CMty1VLCym
eN553+aZgDK/s8njnLVYTOgaET5WslafCCb+gnKsZOWB++U5mVtOTTKp+qeybyfL
WUZN+ZYSmq/AAWcHMKn1b/TwsDB6+0fACbmrZYNrW4lj/TYBnEeEjBKlO8yAumal
eZTq7YKDrjQZLD1I/Ce0tyR0ZmJtoyK0YX8wP9lyP0IEcP2bQRE7WePjfMsBLVh0
AlKerUvEC3hjPR+VZJfBmqrT5YBXd0t8itaFbHKG1oanss1Ot/dFtAeq8XEoS3iK
+H7VGqfGbqUCQj3Y781LBiHZv6XQo1RicBSuNqk9O9b7ltgQeAYlIjncNXbXPxzk
bOJ4YgNmYdSEeM965TRVMgcbSdAPLgvzEN5nEvXtXRT1AnoyLy45Pn3ERPrhd/gH
GPiUrWlh5+6349iAZh4B95PTd7Y8nIoV0xabOTM2O0Gqn+PnicLGrL9oj0S7wZAX
htnDVsJxFwOW7EHXYmvVVBphIDXkwXuTUfcjApaed9fbJyAOr5Yl/FIPiqcNvZ7B
D1UN43J4AvpXAg5MCCfB86Y/L7A7VFErBcGQ517wIreUy2tbAmNhoREJRIlA7wlA
G8qO8Cy5xfIhKb/wsyQ9Gtu7+VpEDjNgAbvWCtqq74j5y7Tfp5Hjlhj4lt3k6mQP
M/TMw/koe5oO3f5VGfUAXyxTj/pqdc7ikYdXFiczlhfJY6Bckc866Y6U+0K+jwt2
ToMVz7IJctdrViG4JstXrQTMFZB3kaDV48bOE8lT8YkfAd70uqxjzhAD3fIAuxTm
nC8+Lxn2d3WZ3UJmLM1XRRT0pnxnZRniOX4B826WVHWVobIDhVw5eWwZeuFYL9Lk
EhnluTqTD+xCpoIZrubZTgSBeY2IJZSCusZDCBuDxjLC0DM7eJzGcg5YXoDH41JS
IIIaL8aVXv0nuVKAdF9K5wktB1NHU/2FwOZgP8mNGh+cXeriLsmnrDH9BvBa+qMh
vJOXVfuy7IjpyOeajUodp0lfJh0lYMvEt4lXK6HiySPvtf+7bZ4U8P+1mzlxMev3
1T2FKuQbBnD8tBeqDSNY90XZ28eI2n4bholSMcRlsXIkLkJeBo8gp8YqLCcRc1Pk
CYJCDLjBLK5RxPgtpu/FD/nARZlOgtHwFKT/GqNW8BYnKvojtzxpkKP8yam2Z7Pq
ts3cwjQVWvtC3x2KobunJrFS6ZUE3ltV5s5gNNI56acWIYd0e8NMqnso0gJVvnAS
IT8LAlZSmrm9u55zIQrdrkt1YDv25I6hB2n7tESgJwx2vHZ9WCzy5kK4qUzvQL/o
sN80Qe/Hjx2zklVJyJt4cVV3hcs4jEmGna6X7Se7+ELLEMUFRTIgTiZHYtTnJSPx
Wi37e1wY5tcoH783QWj0BcHXzJpFRxAI0Clzl1KFEeaBo75AlCXfpvyzwj2RbfPV
8V9cJfbxMV+PLqs6Co6MXqvuB+phE9YrX1R1t7VM/11m1oPpL0nQmlycxHidGUxD
qkpmjSO0w/UVO+WBx4MvoaY8Hh2grGRS0fHl+o3sDW4kHHBMx43R0GkbeYlE+iMo
/3hAOaCr1swsOnICw+TdIZFUFRwkcjved8nF3jMUy/lVWYTR4kB1P0mzpAMakWTg
YOrF3nzrS7JfVCH2m1vX7WKTdLwYZpW3VLWomdskI4a4AaRinQHgfB5+v3bKkwb7
GaHeK2RpVtc8wrszrKH8zoCgpXCpyMJF4JVyPiGzkpy37SuUVSV5jiDr5DMeA7x8
YduGZwpKygLakwRhiM+lEv/K437nK6NYWYzQ1kW00v56Xz7ANjZQzuaiijIovMGD
7xpa1TVs24niXsOX685AT609V8BddkDy+6IqaO6p28APZ9pQ07KdRLKlJ7kGdYf3
AlW6l8xllEMAdYrmPfVXgUUIiW4hlME1ML/5E3CVHLX+zp9ZfRcVnGRZehe2NqEN
/M6KHB4XToh2+/0QGN3KZ7yCCY/esrmcSI9OIHikFLY1JGoajuTgrIpssVaS1xtb
LfB+MfN10Vs1En+RukqdGQpc0iHZsl60FepOtoCh0GJWo1SsQoZOhKN3VOfRFhkq
gxLEQkAjM8Q+NBKDXgOaSfpDWDdUInGAc31Q7qw/5C4JwI0e8l2JMO/o0KPwdn78
VfzoKOhidwTUcGlGnPINqVjR4+7uIR/yiubTilgm1Eey/1MR+wp3MZlBXMdyMRzl
lozld/ZKYmceozPpMOj/VwAAMHd3uAq04DjGNf0KSCtj8vxu32cWnWKt6JR4+WL/
PC2DxQ8M0RmYO/odkfzvviJLq73KklPZR2eE1d15vO149KCixXinFjlyng4vV9Lj
N9vEakVdWdNlMMOqR+c89MoDTsvkjhgzR3/ag56Eer4WDhofS2Tgq601fIHtbhtM
ddAxgAnn9l8jdZP7ZgQu8IyY6/FGHVANnGlLeTsWXTPPD6BMjs7CaYvcRI+TL1B1
3PUDgQUfBugtqKEbmme2zWfXKlXJ4c5dw9UPzIqYJ55zCUZKtWjI0YOeeKofZm8N
10aYZDsVYZD63224hh/5OYYj+fBVjyMXBKHcbNIIsYgH8kqqF+ycaqLjLSnHgmyF
KqM+kh3NJ8beVRbc4LK6/DRe21exVzlB8cKi+OzWsa2ah3RIwBvU+NAwmpdWlzyz
oDn5Ek8k5Buqu/iGCJsFGN7pWidQS/+91nqf3TdeaVnJ48f/o3uzSjeaKuLdmLbg
qoMto3s7lhneng0MCwvsyksRxUDC2iL7lHG6QNMyC3PvCtcvKQ6wU8grbt5ukhxU
+E0BjaioKpvdC+uI+6r6kgZD1fOnUjmaiHrH/s0jMPbDWh6kE48kPysI/TFxV8bb
qzqiW62KR5G/e2rIAd9hLTb84BmRgOU9TSQ+HGhfw02oF8oYmuvrCkndj54mevbK
A4gma+whgMgYmPPLk/Ue1A5AHW/9e0RnNonnod65akvvJE6WDudErGsYSCuPc2Wt
ruiLnxpVV+A+uYMNoGVnx1lNhOrWyXGo6K2/1UYiXblIpz/wbH4jrPgeApWvKJv8
N8IpzPWALff4IUDY+sd37s9tc4zHXS9/JlR9Hf3fVFE1+AyOV7thh3yf8O/Kuh4Z
RY60sTOg9bDtw/ffqipisBInISL9YvNa/MXblhkU8AUf/gtMcPektW2ssvZYERmd
wNmQr22pkXOIKmrW9h0RdN6ZJWdF/mHs13wICwFEi1vhvN8436I3Uh36un8ac326
/hvxxjvarGlo0gGRGh3li9kN762xLQM8ggTx1dLNmgdQKlilYYWgNVtRSykhPG3Z
AEcnTLt3qLMG95fRz8UnwXnrJce38v4OT4oEelhun6//VD4/gHzooToMyvS6fmB0
ZfwzPvK28HpMoYSdi6xkYVIf4t8Cg7rzGeX53tqfBdx7iL7uH204PzK9MeWU+jRj
0ZQm0+P0HQGsK8iHZuKc4Mm0n9MD1KdUN91Aka22rB3l2d0WNUUlzxCO75lxDVjd
74I5Adw+iKgiCaOvG0iZFs8x7VIO4d+ivP3ubmvSqKBGWBd/yuhLfEi9b8kqnkWw
vxcjjW9QD41jZ2FIVqmM+zfzbRON+8NMrXm70tbPtG60Bb3cbvdkaqbRfoe3PkKz
5tEl1CWYgjkvzIjDsVk3SA3jEzy4zqXSoGNLaepoXm3brU/lNDM+b4IWAvdB5Ker
YN/Nn+8h8S1F2+8clHV+HD3WtykD8/zN3qnyYbppK5HHbAEBHVlPgnEG3kcP/gKB
dEiQPNr9hPfjd9tIFtAdBtA3fFOhARPCWsGZgx20OlSjzZXqtcmRvWZ3xog5eQrK
a77tYgHJVRoNxw+lq2hmNSxGQKgA/UfnCROJzacs6NUW3ViId2O+Nk2gslsBgt32
F2kwK+482wKAtHDJfQ3pZzFS1X5O/cLKs3eq8faB2JC//4n/OCpsJjXU7n8e3fxa
qu2j6A1uLAVGCusja/3O2bwcpLMoFEDc2gOhzS4RiSkGrHSl3k4MJwHEesIBAxGS
mIqVqHFb5VdfZ4d0/7FElAGHtEjMFk/9IZhRJWVT/fQVc2nAZemRNByTWY1dG9pB
wQFK0VxBkeuXD7WX+lOewWVuplhkpG2IIhyMZzsFShE61L3X3LWSIx7C3ocX7OKn
xqvEHdpeKfu+U3gVR0bwPcduEz6Ezx+XuHUfetVMCIN03eHHS8+8O3YIYrft9fzV
2pvTezN9VDlCg3zM8pg1IM56TOsJYOR/G6BGMyGaaluoEv1kCw1VUHKBIqT+ef0o
Q7zkT8GE99mUq3R3DnYKnc9dEATolCbNitVoP3zJ1Ksg3DuwUjEhflHuyKBBBL+4
pRYeOCmNStjfcRUkyRkD4jvHTZPvR7I1Jqp/RgT27qqvA1hyfJYrML642+HESsOJ
1j1RZiX7arLr6CxsNSRyu6evT7EYTIj0wti8s7w4ivLgVVa8uuaxbOxsgrjCDFKZ
nRdSshzdbWK33BjCWTv016b0BCHUpjACWTe3TtC0wOFUGt5kITP6ORRYpKn+xXMQ
BGbH6uSeKbgV/yvi58z/dywl94wCuGVJOAmO1/6sHglxJPNxcnrYb/mCYbTdt0Sg
zKC6/n/GRIcpZWxc0OAUt8Axmnto3CYp87NPT6/q4bI4Yd9zCzvh+eRje4qKSNz3
3QfdsiezRjoazpvVqhk47jQdmOKKJtk29zxpYzrYc6ovt9G0/2gsrcUzPcrRHOlB
/F/ZrqPxXas2ZzeBs+qTx80olWP1mtGTfec6Z0zXmebadwzlfHxpU+K6TkbxGsTz
jT7vX33t/HF4h9RHLWxUFYfok3xOms+wsta6iNSQujm3PwJ0FCOk74SB7YRuCGgz
6YAnjsAFxE8hFaxphzmHaun+Eo+xxUWU0QbgRh7PsRrS3e5+8NpgStnOmUljwIoC
IlxhQlzmpu9MbKYX3LbZaeGkANiV28HYZlsZyJ/HwK6QPSzaVa2c4uMy63cOuqfh
iO/nuIl2AhglQYeZO8Jy6/8Dabtob711aGL3k3q2NzsTyD90PScdIlbBfwhNs1xu
hojGCrQ/Gn+lb/vX73Cm4iX48uvLa00+Sf/g5e2rPuf+U3n8ufrURWu1M6Imqz19
Yb0Z9AMNkq+ouMruwqi2jdOORmEgF0FZG7vLDDrb81Z3aHAQEtRX6Tkitty7RYn9
XdMqKhfbCbg9T+bUPkgXd9Yn2el7BMByKBbnsB+cJUbI4frfSRXeIhixv25CXwlQ
3fq3g6beYASn9y4lBNVRHyq+p/fTzwKBGPqj+SCx+Kk5sOqEulvg4YggtcbpvZDe
AroNRCdNhbVVrOwI8waLrk/k1LjXQxEVtnMPwYu6KDpUx3ESj1YxVxVM3NiXTyx+
8JEaCT7emCstVdY0panPbeVPhdXyEtQlUSI3MY/7WLGTYRJ+t400VvG6YNCUq/Kx
mAGOCsClZtsF+WiXnsCt3PiMIbE9d+0Cfh395Q5C1S7QPbLl+Y5S8CdmZK16eoNR
1qw5zgBhe0vFiTiq5ZypIYRtKh47SaKyEHER4zHpPobIUgVeZ1pDyYqCoVWafdV7
AzOGkVyPOGwmc1YQPZk30zhKIt5rowoEOD2hVjhKIF/EdK0emfSTruIDR27b1ik+
Xwytk1ey3h3VJmoL3Jdl+EykQR5USU7YX6FDrbljnIEuLUjS8daVeMqigdX24zZ8
NojpoSuv3q46cmVTdHHq7A06NmCOXFUaOpFYlw40J2PrZMLDQR9iS3d1IXyYJNZJ
H3qEoWwzurs5Zb5wFnXj68UglnukT5qA23wliJz6JlKdS9aK81tU90+p5TO2+5KX
8YNQzG/2odaKzzam4ku6G8MMHF0qLTk7y/+Gb6f982YZNxcuSvIrPH3z1HjVCzNs
u8ogQYjEf5Q4Kx9W6P91fduTa6jICowR9rSh3tWJoUFVhzeDp80PPzQzSwR9La0C
YKCVtypOAP+tceYejX7M0G0cwsLfiLNM6AIhmuKF96BaJOwf38zZPMLlzYQyLiKS
iv4JOtVrH8ffz5KW9P8mdISb/0tPZPU0E6Ant7ZesL9NQmwgIeRaRtXchvt9jNN5
ev01KND6pK7KKdNpyd4mSukeBN/qAm0bUh+Mx6fbd9XvKMGAhjTEsQ1VthvQRgZ3
j0eoWQeOblstAZ4Sf8HPIvBIy8j3miQ9sihnf2oxYFqSyKPQaXgacLjpZai5IuyP
EzPnOzt+aRGsskS4rqmt5xZdGW1Zu9HqXW1j6ysqLLtZbLzPLqjEQHmhL71pqEx0
hTMpqsRkNSqsKUMUWtqdU7i3o9ixMXcaovgUanfzy/1l2Pt8RG5PiZdbZEPXachk
WMbtdrR+nSfjq90unSxbEJ9cBv0dK96416scK7f0me3Z7A+ltnZa9fAy4nF8ecjF
WQm67l0fwTFLOUvUbZ0yuhAUwaN1kJOsWhb2VYgHYm1oArbiZpRs5UmlZH4/zcu9
RRlZnCyVTDzVXwzHkXiU9LXDWb/PN+nrwVGAFb3YzYrF1Qfy18lcuPPY9MKtQ9IO
8tEi+4nWLYLR3WdlrOuDsU8nFSomC9z0yWlhgTEEDd5OfxfBVQ/G40kv6e5fB3XZ
+zyMea+YKhIm5d3MdBY3EQ7com/4MIe4CSZOkqyCZHoCJ3Ir0cRWjP6vwc6cMkKB
T8qE0ELFHZuYWo07Pm8cxo6t7Ly9t1cWED8RI+ceAlxxKDR8wPebZgFYaXY26xro
wREhyCUYmXkMEdnNFYA93HXFTM+7LAswk0ou6gvR858syv77vwBOAJVP+UyMNuKd
TTsl/EAwWmJr40J79O+OWcbDFU94q0lQ66Ha1h+Jgqq6vWIRSr4LVvrtfuPvh7mQ
InngWDmljasgcfmEAkelNQy4JqZWWK0sEiYtoDN/juIMt5TnPq8XH5HA0fgve/GF
ww2Y9vPm6vD4W1qLrS8dFfoVCLr9gARCKTruOOYLOE48JdIin75kgHkIYrfu6+cb
tcbA5+FgB121JVKXDFKYtC86rEoa7NSNkZbn/5S3/tjXSHXh7QVfiXQrPW1/rgwq
nZcowZ/o7VAl5oU5SAvWsfnC85eAet5yZX/jcSLqQw7cq8WdXHn5CuWiuATrgj4/
YEUkzEdp3REnUfhcI7vJ/sodzVgX7OUiLo4gDyP6HdPWI+xaAbB5MZZA38fiEpIM
jqbbmAU90Ml419ZvNXxT1ZHHQpVTEgCpxgXep0IXuT0oCt5u4LqBUFxnxABxKPbV
rftvbexeHZ6tu8QO7QZa1FBcgU017bAbByWCWQ5kLXveG9OWQIxWXHxMc4nKhwFR
TJBISyyaX2RbWrtfrPbO9JyrAvPPK75xIOOQgWseM45p4UEIfvvx7HwaHAwr++3c
usXAoh5SVLwppx7THtd0GS6sl4kW0m1c9r6ITg+X3XQGhS3Ke7G+09zD+d5RFBDV
oYhznvniAkH/Hq/vDALxljXsQQzq19ziOWgDVo93h6qhT5vz5pTqFLN5D4L0ncJ1
/En1HG0jixZB3q0J1+j4epeQkA1iN/3weDR9UaEtlyM9pww/9cfrdj+EBEJf1/Ik
WzcID+9ODIIMZDAUU5ml0LJH3Zu++2qs/7NeXnFNR5EMEwbiikchleuDdfHqHexp
eNk4htpXi/+knTaix1haachrftYhjqv9A4FqSqxOzcxrKCJjD0ViAgWwT3RGzeJK
KVPRd5NGLITICiJ2SvkRDCY8FnLpuVCVgnqTVK2dDfnlTxI+RxmOGYOrRr8EDhJy
J4wDGggE+otlLEMddj4/fiCRbVMF0GD17SAPi81Vfv3FEJD33Szbum0/WULfkLZD
Yc8ZLxk9Y6jneprsr8sjiTk4gxk3KKWardbNG2LquAJxPlfJF96IHy7mwHTKxzIk
W/GKTGLD3Zi0siF7KtvrW0azGoR4IBHSXLZgJ6+wLcvlZ0wFz75vycfa1mbcWCJL
JA5rMeOj+a0Z7K87W2GVURqFMbJ4lzHAyvt3yGSHYJthRw0ayNOEQR4g0Ax1p+tZ
ay2s0zDmjC1jQOrQ0Xd8O+JZ1FxkySWkdrTZfyNqewpPkqWPcDHpBbs6pYytt3Vr
ksH0t4sKys8+RXdA+oiqGSn9lnrNVF4WnQgEg5Inu0GmvB5cVjwo7gtZTKI7diww
Joazvz8alC3aDhwmQNek+BHCU3PckLQru9vfhkjhYO3KzS/vS5agb3Ys1AqC7ztU
dLoT3WxHTt0Z5R3rrbTbvkgBm93vQ83423uWIDxTIrw=
`protect end_protected