`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2688 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
Bckr3H3z8RavFsKxLi9tnJetV6XZKUrPDOKOksEJ9MVJ38LHTiu8rFRvMqLrF6tS
KzZzFN4OcMB03We4oBIZbu0NfBOLLNeSH8z1M23EzlTf+mXzKDLPUCpDV/3yxgsG
58d20vmYFGSkdOxmH7rCvglsV7+FdFLvNxmwfzkTmLqSslX9FEkPpwdWhdZVi+mU
wJlwPqL4xWpMgv1MIbWnRdMW6I4UKD1coZ0ODH1tdRDbikvUJgtU5EMy7rDvuzXo
KL97Tg1w1LyJ4wImZtiFp3SNNjrT4XY4xFDY6LvxWJPOn/yDQFbw7/9aWOyk2noh
dpiH78eeEvM1GDjaRmXtk8sh68NJSG4H8RJshqCr1G2owP4bqXo7BrZY3jgAjH7l
6hE9c9yAl2lO9kUeIC2qXxCx3AITWuPfFW1G7ONOFeJdFojPskhxJiRISCgUJqzG
mHCiNi5l9wnBrS6HFjN3Yrwl2PFvIME3qxlRLKGb85X7W63YwGuGmdKiWjVlGEyj
jlRbvNQR1zwu+jsXYr17PE3C2n5F93ZxyezOlEiEjiBGySRIYMdGuhV1IW+Z59Ou
R3zo6NoW3ie4tILnB/hVTMGW121YwLVdOGlcQ5rKLc3UsOCFkE8tfa8TCqchy/6M
Gb80RHQ9ThqTIU5tx2IcWAUTuRsTiU+PZfouVGJMyeWXu189akKRKCORyrkc7XRB
HNDw4qPqZtLMfcrx40W8wn2uyeTBDkaslaPzd6R7qoaGGdsLpA5acjnpL0QVKka2
+bArNrYhPLwbeRuWsBKiCXnKn/ov3cw95oIZ0cUJalzyHS9frIjvVO52hIT3MbKM
mevZnCmm3BK4DkTAFEvd1qakxGDvsxQvD+hhAaUsvSiTq0A4h0uoqlUUupAj7rdk
bsTITvo5kYks3IVXie+HfVGKWPqb1+ue7WmZmDULQzyPKg74D9AlPD8H/WWXLXno
5zyQghJkc/wJXy8hbXZtZYZTFDL2CxDBR1J+Njh0TaTufk8zPTy1ezSvwefX0gep
WG3X2x2qEUjFZe+c2mZJOkvOTKX6diYbUj9aLb8W+ERHwfLAdB+d38eXSpLZPwnY
ZqM1SLWJNRK9yHUzjmtfXqQij5rN9pWdLXHMzCInT7SoKxc631aCr3Rt0Qg5gNXT
dE17g6VFC6j2lPqLYVaPGXOu5oUz3hDXG08QqDcPdyh8/UgBeBx3GIdrjGzL0EDr
1bbcUo1mQgoWs+ClY6Mh6u30BOyVO706KhMpHzHUwtLZYI0M3eQMiuRlrboc+UUx
cPzBDS0wNa648OFm4KVIyBI3WOpecsS/QjtoJGMy31bc1C/nVClxQ+qdzBjEPOqu
S1CzQNw1TRHX5RYrnLQDxDWWcejasxkwb2Do9ruxjx5k+RgF3fUe8LWU8S09GXd3
o45Yhqv0DhMzBolVq7yQxzcus8tEmJ/nffP1hHbsEl5BV34+uA+iefyadfAnRGVn
0Tler/HwlLyhdawF1M8hQibXo1l0gwmnvUW1/N8NSIL/QifADFvCcgMwlVoceH63
WaYc76wvFo/SNZKygITEZvXLuEvMBzf9KmIF5BgBIvh+2OJ0j+3DWicJ3sTpvzXE
Sjgs43C6+nx+NQTpWathF0IDgia60mXekWV0Cj3kEW0K2jJFiRuA0R13kv++iB+Y
KeU43u9GcpvO4hxUz/T7z3kTEMLAeUG2QkpA0k3aJP0fPro+6pv9CwOf6aPetCeb
8mXOXwjn1zWt73QJLNh/r5XteZ1b0ThyakBSnNW885b2I/sLr2QW4MHQw5m+nVWH
EcChJBNJqebSR7S+qM19lFyJBuHBPPVTSQL3r4I8kia4tJKHP0JvgBoxahcWPCnh
WS3bov5wiAQdQDnz+TXrpqjSmkh4pA/ENCCOIXcQKOenLv+roWoSUvznvUSiFgl6
lf1yM+ueu5anZoCXxL6FY5rd3PiHVDI2D1AFPa9NXddURe6IJWQdLh1C7RtSkxck
m+9tOQYBe7u796IK5MeRR1WyoZtB3zImZDZaiuAXm2Nww69MF1xBzXZ6u64/Us3O
Pzci16r6ZwpRjg0667R8RTec+U7T7J9v6dHXKPDYTgJGwgWlaTRZbDOrxwr5NSPu
aO7e+GOGSfM4I7HGXqTT1Ohni9M+utBl9B4NyVAbOLT3sISnDPw5Gl0EOXMorgys
5fRtdDVpJ9Zyo/0set/Dr79yintIUZkwjsMVxSHFIRgxDOVnoOvLs7IACh92g8Jz
nFJEOAKVMUCZxVhtsOV9zZQ+gwWCg4iLps6hddQCb3HfwvaQIdsZ7FCku+2AqwDg
d8lvG3hZ8yx8bhenpD54tuWHIkAejegctrzZ426q91RvA23/R7nnMQERY9+A86il
Q5hANBqV19Hw72/Ko+Pt0pgBkd3u7ey+z17yGfcpQr+ZR4gfU91Z28o0TSMk+fON
HuSS4jC8feMnrhaZhb8sqvogJZV5JRaLGqKxsA7jwZWqGSG3X8CdsqhkpRnrZZtW
OvjmbEgOTX0R+kxePAiHjC2iCi9ibLG9gHwPl8LJn6k5Dvd1/x433JsC4MphNsH1
tII/Hp2kY+uFls71dQWNRTj7KK6ifGCh/aRCPWG3KCzTjHjCQvv8ubSd1rYx0jqa
aDzUDYAX4AIQtSxjU3ey7lsEs9LMo2PqWwMJsynS8o6w2lUQ1yxIPULtTJsqU0lG
JvcLDFM96dDVYGujHqMaVTGb191uD5lUds+aAolMEj6/dMhq3qGqWC4dA6g52TNJ
TGnUP980msFZZ1PKQk8497OF9MNEJaf2P1QpoezMEvCiGY8fIx50Lw26Jztza1Bu
QiUr3vftlxVcuZ6Xq30Zm9BMKKEo9o73CQsVHIvfZiVZFV1EO+O6NpM9fH/tIHSd
H7IijzJ9ppj4fZPODiX76qsB5BAgZKMSyU0zdSma67mzx21VCyPuMOKhJaCvTw79
6umiK/AV5pg84cl2lNap6wJHHfK3CeICIzqFND1A/ILcNQ23EqNIG696OJ4O69Uu
amrE84zjOn38y87+ZShFWPmR1YvDD367tUmllAbQeGNKOl2lFGHRL9xkYoRDjigT
d8OaDQkYfzkcc6namnXwcsKvmh+DDjE00MZ90l47xjdKNGl4En5dA2t+FkP9JFoz
3v7JrlrdctfNvDqzljJJ8LzWlInoPTQ6h0XICTL5BRvvfRsTknfD2Bit+2C2mjkr
K7569PhNX2c/5el+yPJqgHNdFrPkcNX3lH96fL0Xu/+3vD3Nq0LwUdflZmeLUM70
5J7so/nWnQ8e+LQ+qCu0jpXw5Z3AqWYrAT5wg4rWsNOrpV1VPigpQKWLuqrLNoIh
/FmlTSspnDqMdDs+3svSghixgRffZMvXrKf6zhsIE1lA7aztOkKg/cbPMz6DpskD
rkxv9bgzVjg2bZdwbCb88rq/u2Kl87Tq0lDyGksqpYGvovJ8J3wyeXJssjm7uM3S
`protect end_protected