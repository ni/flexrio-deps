`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3792 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
JoTcvogRvquVnxbhrbrkfEe+jDOZNRgMef6PvEk/MSD2AG4vzUjajNUG2iJV/+xs
O5254EzZoClh+3iIUz5wSmJ+dq6ddzZkWCnNKAs8fezEy0QjU5BIDEe24knjluZU
TDj03IT0W1yITPfPtOctwSU9niNSWAymbm3/eUHLz5pgela2ka8RHcBJusziSr/p
9GNiy8AaT2Jp3VSWtv6QrF+vKDCFlYUQ7opLptnad6ESC3EvrHg7AaUclB5mxNoG
xsycsKixI15TM/LzEhULe2bipjd/YiflCpmkM3reENpGitvf8HQzT8ohJsINJzpc
RGyIXx/XKv6H1VnlKkMSNDMhCXyqYegXYpxgDaS9+007049V0KGY01gNPeZgBF+B
4u5KSV6ncRIMLtFw8ItyZ4XzXIp8kjSpHyGcID8zDpQa5i6DLfvajONnpR9BOvjy
TM/Vw4wQMWAEcpTTBgzrlrGkNR+rk64LJR2ZTT1GjfiQPwq0ra3KhcqsB8aRB5sC
BxnoVOA4vwKcrppw/1rSgUhO8aYDaj2zO+iklLvUgfV+c2g3ODy5FRxUcl6yhoGY
3M8WTDPmKLipPlcgpFUCl/Bcr7mKjP/G19NU8Db3mZ9jMMj1eUgp/yP1FfZf3Rao
QEhKzxqsMhHT3IOI/1MjEB/Y7oPqqhJ1JNolzYbtkJ5MSZmStnxQudcZUQOFDsJ2
USSz/B/iMuxCe6KekTxvJkDVdmZ/1ARlq49NUxpaxYmHfwHBZB/Suq+ZY/KZhFNy
NF0DYUwF4F5n4umTfMCXZtizDI06rcV2rpzYP1NOZQsp6VK+JHOLXUZiciL4DbWh
KQVyIpER50LCLB1TaSUkwAl5cLyeycmZMz1Jv5QI9eDtrzmAoT4vTOF3Ly+Nhq6W
Voa+9zcZqPppiPnqx3ikvJNAMWq46J3ObyzCYIsgv+sOqlANPj03uDPKe/lD7Hvt
gjg9Qjje9/YdAp1sBpgtBCR3DJJgrvavJkJ3dF/qoOV8dWast5KfS69YHvTwCksA
+St6A5czhZ1RxMLMaM8m5CDGj3b3GbUcLvoSuXDpUG+QjlD+Ndj7cXOix/cdp7h2
8CZJrNvJXx3GxBYavhYbBPj8+eCjjcycNbqsAfMv94D9b/3+tslCq7znwTCU4avy
abmbONTekxmirrlGjdkNgQqKimlmR7k/ALmTleLrCHLlEql4qrm7tO+tNJSwpSxR
pWfrieIYywYn7p5xMbBpDPB5jaSOh6W8e7tw5iE0vyF+mZJfv3b4R/MHqOwzOo0U
fI1mMGxAVIqf8O/FCgoJsiYRRhLQyF/0jBjA/lIoXrMm1xBUf5ZfsUUfg7gf51J/
1dy8LgDXq+VKxUVqQ8CAcMXdPKM5EQKl5UiC0jpqLrXVH/ZBocTuxGOQMtZDrSkW
NRS4pGG0uKS3l8adb0tNgoFAWllTFaEPrw/6+rVI9hXfQ4FevroxpyAp1ju10pQa
xt2tRHhlxiQJFCfjLJpRIZ2oOrU5nphyG/cX/t1yXg2XEpVs6YlU5gkt6Aa1oHgW
vclReiJu3ankM0gLZl5JgPbPmceTz36DY3cKCASZLsk2fBoqwkhmjd74OI4f+rB4
oF9q9RC8z+hFQff/WOKbpV3wSCK5QP3cp/GGwbRGsBU94odfHJFjUPCmQ0XjFvvQ
sXUN7d0VsXGQeGeLXogk8RFsbTwdRwQWmuor85lU7vMgLbNNhRmuCkjSH1mowl5l
DRrWDI+AhhzDVdKbglwlIlkgZBejs61S2BwTo940gX9kdh9fb3VVJGclT0BGmUZg
biELdR4gdL7jRx4RY0HVuABl5/1mY3294nXVmfR0B8azXQ8d2LMdOiXsCP9P6cvo
0DDrVbXeeV30mKaRiWBwFDDrS8HoEa9ldVBR3htbYltR2L3d/zPQPmGuD5DXAzr+
1mkA43S46mCufbv/49hRsE8PXXhWT4qBq9VX1N2+F5tS3cLqMWWGiZrUaP1DupMm
Fy7glwuYxO6+42yWxTD4yFJVPUfLU5/N4WRgt5KBx8W9IsXIjfQNfiyF45esjse/
pjcsUuFdBQHxyZYWejm6WqbmDCi7wn3nZ5YONqZKbjxF/eiROST8cbFzyUEvPFL8
vD29ZYT6l+kP310lE9moJwoIaFBawD/mJsXjvRC13+cWQ5bbSi+obawwR7t6adc4
yk81yt5uKnopCIaLB20SHsTHopCkpjlDTygvv0+Nex5STY8hTf/iYgjrpPLkpSln
lapWg5oF6ABU+wjgFYI6f5W8IjhITnsmf8xIrGUTVbcQlyGpBi1MAQh+g3OpQpdB
bPyS1tEoRlqH5kr4IlcBbsfnQfaBZYPuG4t7RZSCOiQKGj1RyjsVAXLEcH1Cud90
Gil/6PB9YcBhfLBt4AENRmPMT8lib3BonEQ9Wt8AU2ukHlR16vwgDATv4PNS2pNk
HGRHLWMqbVzLLpIfgrCAYniXGGoLgEjaX+cuKfHwSjHve9LiQhFZpfB6jHHHA265
HXcgqXmoBtCMsp4JgZstb3c2RtWlFEv/JL2WxHKoD/Lv4JAdUFHyVg07viFsi5h/
h19eaKEWV/f29u/orhKUdfwy4w0fy0MTzAHH6CKKNHgFmrVMYGIFI5OHp0V0tD1M
1Ei0umZ1hrp+HLA7H2N/9nrZo8Z1BNKqVify7tUWOnu5qjG79jxKMlaVB3LeDyqW
xEYKus94JATJxwTEO/+Hlrv3VkJoQdrwnFwsBQdpUyO5r5TCgvGHwJ89sN8lHVdK
4x1L4X5LrgUKVhNZPP+f+1o5xrkq44oClTqYqH7buwGLL1AG1eNjLrXatCXZK+Ge
vh82F/kJHnminl3UOdnC8rTPM+QZRA3m/hJfNUBCIUWvcYzAFqQvY3FKYDXdA37j
xBTNVvGdSBWFdreLohUvYeyV8ttkNcmOeA6rVXJqgllFNmzSboSavZ3kGNflvKSl
K1Gg45Xroq157a9z0/ZhhtpW1He5X9+TLjrNW6S/ybw9k1FfK5lJRFccdsBbBd+x
4zEoh7RL2F5tU2dTgvEOHsZ94cBPHBASQJuRZzf2RdqfVQB30lUakbXtiAFihUpD
afihizBHM5x/QNX3VauNJjalB3kS5OHb4tTnP+bZ3uDd8Ceiwvtlbg8IVvd2zRFe
bYM2pkKp7mzI5rjWD1vsRdINUDUTEMyeGRHjpzE589zTX2jYMacsZjHlOkWSA46/
Hn5aHvMS4DygoRBDLtmAsyj2UgmdEjP2TLSVkmi+ijXGdTIf9qw5Fcu9aZRnQ5xO
CAKnxjzZqopcqXJziP8nkAkx+NlMu/GgC6eASsuLHOmpd3UsskCYYAOQAX4Qyg2Z
+eB2V4Ye7IRJYbyTY1UCqD79FBmlIMmZt+aFE3CskceYScLk1pL0+Uggl1CgUlIS
O1FSyofQphyTkvRsCWta9c6Ucy1aT+m2pUy7RL/hKcwiQRAj+dkbawAoTpJqU4g8
j2qLaPKW7AWGOoXqSqbty6dVjLJe0CJPNQIT+nGoYhx0kLnouiLPaHguQbrN3gA4
x8ophVQXwq3H2psliexKaLoamqsThdmVUbA/ydShtREVh4cujKtl+eRVcBA5YyHc
wG3H35UfONvMXZdQnaPMKO7743F2QEcfZf7thfTvdMilLaLD0FcIX2rQsh2FWz0Q
4RyTFazZNxECKLxS2st/Ps8k9DIPc4jJJB3rYKKNxjdfS9QRpEHqmTfov8obUlfs
zQsYj+T5aDEy0+ZfhtaaRVd80M7hiyunaajdo2L5Ci5t+fdcvd05NIiowCF4g2e8
PHhOAkNgRUNZgFtGK4sWpRvo8dzbLwTgldQ6UsolXpWkvil4/5DLQAn9dm3RSU/F
tv2Ep7GdibwhnNPa6egoxUGXyf/xI5rwygRc9May5CMw1wFl8jyHxyG1Hu4wFdkY
2aNnxEZGHdGICsfyd/agSrQi3QQsfAZw6850wT7WeuOqsjnajQNymps9RJdAG8wT
Q2Gn0k4YQmTwhXAkXbeGGw/SbVQhEawKQMWQunAnkeuryJ0YGmUpTv/vJXLbWN/P
XO20AYkiMqh5sharNKXoOMdFQ7kne5WXhPFDp3Ccgk/J2AmcfSYhXzp13KW8O3uU
QULn0hxB7nVNDuHoy+WFEsdYs5DeY5q7sqZGnqg4/f9EbkgzpuIIR3pDKnV9kWO9
Qm1sB+DDUytjgzFr8qDyJc5qJtJWeJWheEQfsyVBqUJCPrFxzz8A3rdVgzekhVaG
R5W7MrnErVYBOfXJYoslgrpyJLXBCb6dIsCtrrvY+9psnzk3TltJQOKeR/adfbVK
ZspDDj8ThcFGA/prnQhnwdjDB9QLvXaoHK+m+fC+j7kThvL/jRUa8zZyIlSh6SP8
TLboEL5WsmAgGXWjkS6pF1ueVXfHa3l5AMdud8VRYNNE+pkkKRfMtIFtuNyICtCv
VxTnE7hbnNvIf2PkAZLQ8+7wL4tjP1BAk5vW4bHgiITvpxrbv0x8zc8mgzApTApn
25Mkac8fufPBSKWPtgXw/yur+WlGd4fSjTwQ/RqSIvbc++wJ0e5YgIaPTMh5y4nD
7vdCVixq+p/4K6rn89DFEH7DgPS+SHNAEkDL1Vd+Z9OyoJKJOJ919DzRwXtuLHQn
lZxDYMbJTQexvB+FR2uE+9QhxlbT7TKxoQ27zaAA6UaHJOICZNnR1Qxl1gXFWXzm
M1U+CFMG4shV+zZG3OAnGUd4o1nlr+3XJLcSPwLvE/OeKP0T9lwaYgW8xmzgk2RF
zub7r4oYD0SJ0fMglxUjAiXVQUNf+t+CFs0KDd2MJZby0f1jTf3AATL6GvhHwnVg
8GFoE9hFmD+wYj1qwzycR8ZRTKbE4iDizqQfKuCwUmQuzB956R3APgIqUxgwYjmg
f5zPdAzhxGi038nrlvpuz98OH9t/GADZBvQ91GzcJIvH4/41XOHpx0OlVIE9FDOF
`protect end_protected