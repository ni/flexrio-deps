`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 61520 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
hRRAlfE1xLfeNfywbrz10Aj6ITcDp3ZEwpPSvXmLllawKpK57ld/tA8bEQQGQ6iP
dAap3Sn1pHgEZi0Ivp0WtUppBocZkAFGF+vOXrPPl2XQH7UCFRIUZaPszPhFDqex
FBE18v3xZ0cp8lVwYa+AHStSTDB5+mRQvhA87MSdJj7Yg1VWmDKYzFWDoOH7vWPZ
xdFnH+dNfvxSMH+2vl8mqhZFlHrXob6t6VEHe76Ks2iOBqScgZ7oabUTCj5DZ7Ck
6RiXEH9gSRHEqGAJfZWKgxapSh9p8h1ewH/AaMphrTcbs+5xi4BEYeSOKSSnCOBD
MNz/XV6+ULk3gNs+sgC1UFGPns4iZINs6odFBC78vFmz6Xh7O3t8cf7IZdj+nF3k
7CZl6R+wDEc1KK4Zg2T+KuKEC9bawwl+QdAozHfrhpuRYxux87S6SJxw3PYIWyeh
qR0pERh42fsM52MSQRcb7kL41pk+V1/xIj1BZR6loIfvY1qppj+lW/gk4+votiIo
MWF5hXlI/oGmRdKN1GV6ikaE/zsR1v2eHqqQSVntOF5YbMQSlp/4o374cRCS+Oxm
cQV7JSmnV1+Ao33LOSQXmuGI7FvRAj/v8M2AWNAneGCMxPgOrHizVbEIDpiYvWPk
4tzksOAfCm+4Yyd/RbAUeOsso3f4pvlRtzjSsranc86P9OagZqqyuIvP7J8vlqrE
VtAL5CmnsEvO9sYV191FMJNtSfPfuG/gSyHZzFK37+lSqD+pO8od1IScNMyXDm4y
25c5oWv3nqpTmW+R48SFyUZjOgqZwPlO0yfjTZ3GO0iM8x3ssVZ5Q44dIBB2DNJc
p0QYnfABpoZWjJXZjIfF2yDdpYYgfTIavQA0O1nuAZopxksecE3RZv54KheoqTnZ
woCjt3lfOKLh/ysMoxay9p4tHyLjNG26scepSOjE/rxZDmj2lmNK02kEtjdJlEr7
d8PBkK9NoPXvC5AgNQYQ+KoJssdp4iO7SOsY+tQljOhSVX4wZqG03DumHLCLzKhJ
IheCUPv9EdiVQsExo7vnAOeWK6OfAs1c/NUKmZpbkWUWAoJ16/M58q7j4kmfRXro
qoFRFqM89xO0g+2Q3PQTlQJ3BPcp94TKheEMywhlhx6gylr8a1Gex/Cm/t7SO71T
E+lhN4qmg/A6iOTKROTkXkaZoBCFjoj0IWG/1V0W7TLBdC15l8r/N4dWpOuiyjs+
Desj+ewGZwIW6n1MHEwcZqfmUtyWE7ZSJC5hEFz5Fpg6SHKLMxyhGIs1SyzXYCP9
sAFo0Iqnogwf+Kj5TvrNnmFHrnYC1HLDH0DC3nj9Lw8QhbyxbX4PhkVZtEdH4TYo
tMC1P3BmrYg7BFO8HiCmZ2UDD4xbiMNcpXnDrCN776L7+J5m50o4Xx3SwwDCldmU
bs5v+q0NUnfDSB6Z51gYzAtoj8w4tRW6JdBsfsdTFou1hG5xM5m23qmIKb7NIBHq
+9J20QQU5E0//BGpXJz2DZlohH3PegjPmXTwzcMGHD8g+VbAWOL+4hPdyeS7AgGa
PFsSah8pDfc8/bkaL6otOqFij0x+1dvXgEONyoITSRKXjA2QYvTlL9MymBi8rkCP
ZAHTTi16kjnt74+rGHKISRZL+F2UMJ5lp7NQnVInqL+mShzJJwdonmNTRBkD+EAc
XBMk16EwYTdx9Z9i2IEGDCT+QeRMPr3Vytqxj/rqBZQBBuq+Hhq4VkaHWpI4QpJf
70TSk6XqqRQRK8XZyMKoi/a6oA9e2Tc9AABzoAcdzseN00tdebRehbmUtvfxhzbq
/F+eIyTZ6cRP8FuAg1hzb+S3OdPrio5ugCx9XY29pn9TOtrkPstiJvjK9axkk1iL
UE3Neak5kdB+TJVC7NwtMwiotRXYpAUcRS/ohR/F8lGDsrKn/PIKJvQ7EprJD5js
b7V63LHkHBkk6+d5VZTgi4Ca6mxMUPLwUnFRrOC3ynV8lOrMbNPSqjoBFWALO+zg
jUc9M9YP62yezPueEtZ33fsuJKMEaEIQ7qtfQ9a2mhMcEHPljmP3mzO9HAalWQHs
N+sn06/2QXaCGzCIkHTMmU6MRKUHm4Nuu4qhqNzU2i1isu0iEYcyPwowFnPmDLv6
d6cWk7+r1Lhvg0cjnoRNosSzDCX35AtCl8OJkZ5Od+t4jU161K1RCm2ni32IPsGl
36FVq8MNBUPwj4DGxTUAZ8ddYDb1DcPmlBupeKA2NEGDNbw128RQMZeoqgrugPeI
gqAglJKyyjhDy7fWKDomLb0k0X38Ff9Ork9q5JIgvTFmXBUYpBvSuJPgENIwlJuq
Ang7lme/Y6TJmbMbIdJEghA/qMepvrAH4A08oa4zVMwWxNXsZesfwQbzgfOM+lJB
4wUKS8858tfq1bTi1BMzIilmxkoDVR0VMPnJ740UNyatiA0y+0IvlldGgeh8wLmm
cHYJXOz6ztcbWZKHFT9UL1lB5OKxRT4H5DjdpQd5CHErntmQR7Kw78vqWfeIFxyI
uB0D3jpOxPy8edic7ejjVYMvXhV7nhpjn2t15KTzSoUUz8QXoAPDxhtohqqUcqLc
mCpxGQTDc5+FpYVyGVED68xFe7oDAOBBueRTIx43+qdNzCfhzyToBLL4y3mAgjYl
Hjxz8Xlw2gsfkl093o5RbAtVyV8BbwylvT01/TVUfHAflzawWt9hx/WwCERluhr3
eZs+QrYfkNoznx+8EUhCe3A2b2He4H+tniswDe0sOmITisQdNHipL37AEIbgBx7a
2/XIi3LY8S1FTlMZdC+mOVLRIoabf8+3EA4itZlQBR4PFS1IJiP9IAiU0AwwRwW8
8jtpoHMusxBnq3ZwxLFso8pO40FklekIN5mjUgspCDAvogW0XxRNz0MQarsguZOr
Cv9z3+cQj6oR6EmBkSNf69dI6e4WNOgcKobsmoNTxmr9K7SDvYwCUcHCNsrTnIAm
vbSfcIxhkGlmIKwPy/mjUa/8h6Auv5jOMBh5aBUVLiM7SnvkGpvdIzbxcZMfIZS8
XezAEa540dMRtg0TCrpjYmYyB76OXiTE95wY3R7Dxcfqvbsjg7ThWJ1y6EzVydVN
y2iXjBO6ancEVvpLhPrTwIs0iXIXkQsalWQ0ZZpYMHhLfncWZOisaQ4R22Fz3poY
fGtHpdC7Enpn0fKX/LXSkL6gazzgIrXMHYxGL8/o+vYuS3f8ph6U2TFJBRLpT9mq
/HNxDLB+nstI3Lg286In0XVqs+jP/rPvNewp+qDV0mwJnLJevlTznBefPHWQllBH
6yBFCB8Lk1+y081J4/a1u2XDvEPTu4Z+qQ4ZkhqqTSNbHRlRj5Tgq/BaJ01JP98k
ato0DdjNCwQ/nHD8Jj9/B6vr4lv0A4P7pj+H5uiTmzwO7AZLd91X3EpCoT/1yyLL
itQmOZyKZlf9BbypqO9gSDN+kfn4xE3d4vVKlJR9YHhpTxVKE5xa0ABxu94IAdNr
dNtXfH3cetQm7L0xtTJNnNKGwa1RfYXt5UlLDKSSHF9J9MOpNAqkwIVF9tpmZ8MQ
N3AK7Da2I+2wbedFfJ4CpynqbOrkIecmtjDoEhJYue51Zo7sNfMzxmBgS6Zy+5zy
s8+1vl0C1uMvBFNpEzUROZQr4qYxxvqxgyuPxV7tu6OPk/wo905Pf5/SffXf8/tE
ejPvYq58GiJ+JKrny9xIkvHybyp9sfUBls+cF8EjkgduduQMCJRiRGewd57eRwdI
pdgETW+hIZqus9pICinQZvlFqJfESeuuzY2tV/IKnbmZb9Ve7bfNdx14uHtufnYu
6ySMRJc4SbgTWrek/rdK5CNihcOzpRqC792PNECO+NSv7OL6EVLCGbvLCvGMcN+O
9rP5+nuHd9xjbfcb3G4kLPgzoeKWaHIszQrTEsXR3Vi8V19ukonKCLLEYXwTgvlb
TB6NlWiRDYnvoyQzb1Y6JkeOqE8CMkKf5QG6ZaYr8lpkxN3SfJZzg9kope6mbkHQ
zMA5D3H+eKc8BC1d5j2psNzBC02PZNUIPblHgAp7JX98B3P+guvWlsEq6UI1ZWgh
89ydxjbFRXXJwb+2cUzyoueuZhdj9H3mbPvRjGdIJV6akx4bK9WAoQ5gZvxqvpu3
Z+SER/oHJ9RPgHcb3WmlamhEX+O0Hr+gXkvVA41xMQBhWbCF8pvROdm855dCYVdG
dWxAdcPsDrEoox+5mcPhq2rOKCRKW3EEZDGf3/1dwg8RXGID44QbPC0iZLXfZs6E
wGo7VLGUv10W5zWVpTSezuqXrLhE1HAMOAFuXOZSc8dxn3dbwHKW12dXZi1cI+UQ
Z8rxtiU/rAonjP9Djmpk8Y0d3tZFODvtVsEnukUX8ER39Ss2g+0mZQrrSt8TUj0W
XcMOm/LBO0wBCnBt9tAGY75OqzS8jPsij57Hr0nRSRQfIHyqX0Jkd0NMyiShWp9u
lWY+f/vt0i4z1j15nYIa3lPn91jgF67ft06rg5TNccxCNBHENDBI8I8uZBHrZy9t
yy3OeSucbsJr+Btfx6BsRoPpnOZr93ITEbX88x/8gEL9Ctshbh++LiERAWgyN+x0
fT79w0yTXUYRY8F36glOo68gW1gWp4SuA/B5+b1GqQ5WPkEhmt2GFtwhLUNE/yew
15aOCsSRIG2BHkU7JOMysdv2q1Zm3bfBTYbzxgBj/G6qr8e7DDk2nzagJRkCUDLm
bC9c8IXhFgy3i2meP9+6oGnMjWyNofl+tu6CB3XuCrRSSSmZwJHxUuYjH6xwX5pJ
40ymobhGSgEm2PndHEL9GO7IfQXVfVzd14hnOVOnO4IqrFqWdk2bVHZVeof6m8Nj
qUaNEb5LoaW+wlYndZZpE97XW2E+3AwMpEklCozqTMPclUvVntt7ZDILkEC96Ye6
4gn1gLbunlnWRbwVg7+6IMld2pxhb36LSpNXiJxT3fgEWGY3ykMPQW2JpqVv2kX3
6ISeUYxPFTvmVfie04tS5ozY+5S98M5Xhf7le2JZ+xuJ4h0cMCChw9ptwCs04Jff
Ooz0cEiz//s1g6BxLnnrvygx12Ljk1SUTitIaggOSTae+sJIciDZ/l06pz6NcrRk
77OGB5zoJTm+41O8tnIJxPuI/Do352wfF+n+JKNuaGgYbp8yMSWAZ8Ox+LhZ9+go
LTqZTVvOO0LzsrhV/CX7EUkMtkPI9JiL0p6GBqr0Gv47rzMdZ7v7YWSDiMHfAyMS
4MrVL1FRHK5JMv+xO2Y6AdGtp/2N5e73ZGL27ZDM6SmvaOvnebZvQcQTcMxcto30
M2zWgbONfWNmcSQlbIFPomTvFfLbUCw0I9OYepgpo8kawdufcuIw2me63Cb+G9Ys
gVEB9GqNJSRTYyF/a+EKhbTe3Qf6UQUr6Bni9BMbWvVDsFDO4jJ6TpCdjDPpvemX
ktAcmGUeMtEbZIcFredPA+2OrfNDbA9+SOXjBtx9yDFgJSpcpymR9iY68hon+St2
0TiGqXEqCcFuSqtyLa2R6Y0zeIhynDVtbAUjXq6TUH8Pmpq9mADtUdPJa1aw1nM+
9PhLjbJ3qSL+TuXHVKyGQ+Nt5yG+//vosVjj9YLlGdbECNUY+yIs28LTXVj2FUNR
M3M8mop//UAtICH3hDEQAZvoXUgYRCmiFPERHw9vgEyHJbQu+h5vUvFMVnoj/JaI
v4dklbXdHWH5lt6+NA3DIt03SH7lhuI23GIF6+lMGfzU5GT3cRoXlvkZpOgAz+1l
kFitHVOEQN0nH6U+OuWiIX5Ht/nVUU1zYvmbi+yASDFNuLM81O0V2m4nny0I0zDF
eaZOil9MPTsSQwhHAcBKVXGohiVhhjeTfemf+kEoROGEYr2o8DkvPvHobJSdvOAK
+cSCe8QXt6WkaCM9fqaYuivrO/QFaxhwUdCHHIzjzznVmxRggRjLn08Qt71lyZ7C
azTHmKFRzJ3TP7+8obKPrjIZ4js+zjPkuKSAXGmScgJaLws1c6cb9Zofr11sd+OM
SuEHp0ZW19HxVyEp/QP7w9XtD3UjUSxdNp7ed9b7Ys/kaAi2Fq/HL5WnEBY2MFPb
ohIwfvlDF9TjcofHN7GwNh3zMqnSgvS9feGTGdSU6YOOS/v8MQrpgkGhvG3fF+mv
aoIvNSr+tXPNNrAjYm1XtV6BnDO/VOtw7AuycUI62l6CO8aub+mxLLC/RhqL76H0
7MjoDdvvd4AO7/kNmOhbvX5gl1pfRAEKbscIDZGCexpBc8Z0M9Qo5thPGZKFQCVQ
hReZgKINTtEIDX9uXb/7pTwOG+mvEHdL3yxJucHVINQX6ptW1damKodKpYOFEla2
btc45ZGI9wgqSvqdV8jwioMX7ELKLvsV3GPjsldnTPQbnE2b5URHMN/3oIAAM0Lc
wnQJbWkQr3nv57Y0kpzLtIczG3m8ce8lcUjolkEhrwvsOc9zRRo//xUCBfDXeC1p
J6lVTgIHcMA+6ZsA78GYtd/5wdbK58AVKq0WcYtc9DOJ9JWvm2QPE65G6QO0QFML
NOEAg99bkc9ym86xgK8Rk0j4UzcAYuUzSDVNuZSl+KRHCa+q+mmhwaL1k74OQ/N8
mOQOUnUbFCkUBAp8s+YFklSz+LHTdJNcNWZztvKT4HP3NMhxFEe8Fi+XGdU7uafh
traN8VQxR0+khvNca1fKSSKHJkTbR6u5yCPqrgBXXIMXunzzpA3k1gVgOvHi6A9Q
SzWtqhdt1+eMmI/7ky1nlI9M+Lx9nV1MpBg4AT8wmvYz7Nk4kHIcRwq+HZZ41V4R
uNRtZ3Fcn4a33b2WlmkTn4Oo2ITAJ4kIdOSmDxNHliHqc+Xh98u81/ErkhFwt0RV
IIcUVvBYyFNSluYHIRHAQ9aEts3pwYtpOySflfRZi3zOzMoIV/y/NgVh32JaekUb
XNGSA04lze6Qb0t9UiuFalWiL3I/1qBRFF0FX1+edBUC87lq/YrMOqWPCq9TkfQN
dzhv/L7xeoDrfa3NpLmfxV8pOvcSDetdWj2+CUid17qQ6x1PzELciCmwdCkJGT2g
xk/qj80gGdGRLTGvVvq6akDBwx0/r6Y2LS/Vppi3j4xot/GYYAJdC9KgaSFrp4NO
EusuaB1+41MRa2oMavXoeai8H40DsxLCaY+PSZLZHrFxmAyyXhmhlM8GY7yHn4m5
TSZTAbxCjAAxJM11nLX09aU971lmui9oLHBIr9siyVu3/PdxEME4Fz56U6G/daAC
jySJN1o/yJ4WJMnXWwTRObg5qTUTfDxiC7P6wc6BCgcoOZWEkepQC61LCRG1OQHQ
faEckU7gHzNeHFybPbuSPyXEqXIPclRWCYLH/LkGLdI513GXNcZBpbnHXR59BnsC
DR0DL+61QHtLU90Ue1WWQFdvGfB/+XUwrQWoA9YR0JxX2txYz4f02Ky6lPhaMSaq
mDfgddOnLCxKBg1XJOCfXL/Vs67HsvqDDg2KfKQULc+LMnYFMtsn0Xlo9nxMotOz
sBLPpr0E9oSCE8MDkw30Hm+QDIffpAWE9k2Xi/BLGbbppOmA5PvQms8hmLqnuNIf
eDjoxv/JaeI9NwEUBI8Nz4e6b+2A1QyG81Sxi+N37YWFUNO8CodqM8F3pyccidD9
28RIPbSqzuG0KqtQU7Oqi1ES+o6qBFp9DXAk2kPn7mmSQbegb33+UwbSnI1wvAnI
OW1ctimKroxqNDlvsDvqh9QCUpSB5rELxUgOsJtP5aNxNjbs+4IKhG4hHSWz/0Fe
9x2rGHn3wiPzyE0rZFYFFNgoEsBPPKkElDaGXiw9LnvZTMbLjlCg7IaJvQT0yZXQ
GkO/S+d9w4cC08jzHQp6zP9h/vCXZ8YsnHX96zwd9ObldCpj1DU8DYS/M2vDHQ5V
6MxH74sq7LoZcWG0mu4XIeP9exIu5TEe8j/T8jDmJk+bmi/07acddRWuqNs12F/c
ePlZviMhlokkYiurgkUMWF1RQAE38x2Gcvypd2/JmONxUVbx8jFQuiOkVZQKUcjv
FYwt/SGAjVR/A7ULitpcEZW+pZnBUCAarMD9AOKXrhVLgVxs/5NLt2YaYcUff5O4
9JFC6Kq+VU3bzMBo+KCek7v2f82zQgOSOJJp+H5gYLeZ8ybrviL/fEq8IRKQa3sD
haJnLtQTbvUVyMUTbGzK3lbR/y1K5YxR7kj+xLoT+1/C8+O+r5P8JMx5uI7z1S9m
TuwsPNkV5U5J5rO1tD9GPfSY9IdMaN4XJOI3Ao6Fr1uNBmh7nDHHcrwyuFHZ/rWr
BmJl12kemdoNPv/h45WrHG6ZqTdFI0j0kmzZ5QDiv64CNe68hk0nsP8Hrfr7dXSJ
sr7qxii8LEvKUGX8FHtwaIoShdtgN8+QRY1IjZIyVeIc9x+jymR3Gh9OKx6TVC2G
Ww7nar58PQ+aiqY64CfqtroMYJ2b+wicoxkdQUiLIaup5SyAIOSCwGskW7e//Krp
uQGHVDemqxi/r9/st/9PwHPmaA6b6joaDY15wZEjVvaeKhcgK868HYqNe6IfCNMs
k4R6Na4tV8w4zTr2wqzaOjAyQ2FxFQUzZJHwDHaUt71SfPyA3mODvo2YlQARdC8S
GnPXdU6K4+mxuN+2aQVdGBZ+iSbfLTdiMvXH4xuXtdJlwp6Hc6AId/Zf3aAwkVhN
DSQfLuSfzwigZGvKyMq3daVJ8d5ycKS22QJwdDq/UMFUO/vj53TReUZGrxGGU7N/
gFreAIenH4JibyLDhaxPg5nhZn7z3fHKanFr7MDDHLk2A64/9tlxglWr22V/veOx
iWIRCFD3BkMB7CRUiyjmKyHxbBbK8/1sAaXYSFwWyjGOh13yHlpoMbNmWPhuw8k7
wjI9LXMdO14uAkc61ADn2JXFJPWHZ2BLOL5irRC4jrw3HBaA1Cx098GsJ+yWXKLV
/ZeOqHtNKdvE/5pooQsIgOy52r9NKNcrQGLcdr0WYxLmqAfetGozQXpeGAvIafsf
2p4ZW7e3ORkD9GML3czRb7U/gZsk8xgl7O+hCudVao8O+zQFaAWep5KUOgbvmIdu
byWQDfo+iUKAfgueG6WerH8lNtlQUB3FSjpuEPsPA3ZoBJnkxNhY1lNs8uRkZb0g
IiLohNcmGCpHY/En2/EwFHxoyf3HOjMvjseictmExC9kFipI3hnfD/TNAmc/Oihh
mh3rddM+FI43lgyUCNBNwF6ibjGEsz+OOfZ+TSiOt0LcoD2GfSIOEWKAM25MhQxS
ydd1DDUudcuqzoiBUY9oOpOoCmGKyLK+BgSFKf+mhWfhTvqNI+yeIH30A9IPJ0e7
FYyJTHQKjLDutbeLioSwG4vpqJBf794RhrP3fjTYLhu9dRWn6V87DMXgA4eXdSfK
k2FKFVVF3DxvMCMmXcIymHdSpPvuIfoREMGefGAoXIrLstvzqRvUw3u5Yab3YZdZ
n6R+jT0T3nvT6SBSGs6V0PJJE99UCnlH44YkpEr5LPlzbl4waG7EABs33ezTVovM
YieYQACfIy+5Yqqh88YGmQHbvzXD/aA5c1Xd46TXHKchPDkcyqBGICmz7kOFcw4p
yQkRV0jSq0CDqy/i8y6Q4Dp9pF2oJI/dniJDALZkAEF1LOqsU8IBcrQ/xKByuvbK
R2hn//xcUqXwtLc0xaWbiv1BHBIO0gjPo5mLl3YyLzmV9yaHfcV84/rj3zKysiZN
xNRasug+bqlARfiZGZj2wmQ3hnL3OCVIjliOQKiprKUIdvaWRnQ9/+b5UQPX6q+q
6aRkyojJSkW3arW2LAgh00ufKs46GaoyOVRli3WVSOGMQbKUkNVFXfSuxWSyeVJW
GF0N5wXft/A3BxkQd+A1ci/aFU6XcuAHgpJQa5ezcOMg0FND4y2gBk1TJ/d28iHW
xXReJCS48qO31HMwSIVVqsVxWddtBs6C+sSK0TwtjCv2s4DLP3wCIGnoej3wGexo
b2g/ignjFgFkZr0k9DdU41Q9y4JM+ZAXfbS6gZ1xVCfgCwRk5zNHrsdmYVLBvOCc
H507QzOmBUPJFekMzk/IlSu/httelH6wfMf4m1k4llYms8qDXEqd1tMi+r6vZnrE
cIOUXQtRNj3+i63wIhM2qZgzdybVaLWa7sg3IlpRVqG3ULzHEEuw9hVs1K2lYch5
+ZtpmrzLzQ9iMlxirEh7vC9kwrz1b8X41obx5CK3jaht6PQStSxdJjFaRB36bu1U
5otk8bCA+njgYCxFVwr3Z3VvdqIbe6x/xWJFIXAgcmKp1T/rycpoMA5PdBi1HQxq
DV/tGUBTBm/udsE5sMP27/Ov00fS5lje8+TLHJOHBfXRGK5y+dYLXFgKmLEmdlvv
aAskbK6Iew3RUI/1G/g6BCZdXvwFzkIri1lihGu6Hh9g3B00VtybeZVMuY5MGydh
I947rZvY/XN4gV6lohN+jXmv3I4iXoHaIsN+L8T3lXDeupz3PHmRiAjehdW4fCv+
mv1d1CXYDdtsbErHwqKUQwBSxigtP8LSxL367pSkc3Ejm/KHVt1aB0s9d83tzrI7
f67d5x7FVmQmKTduBzqSwSvciSBcmKBb9emQLnObimZWG0aso0yRXg4OsFHEsEYz
D321Ma23v8dJZK/E8XuBR25cMFxX2e75cYOmWZdYXDN0LrwHXZJJQ5AbGYBJNRLe
C9N/b58rpLkrb+uh+lPSRZ7+alGl0C5lXQMcuHAOQelZsKFcepD5tGFlZ4UE5E/O
4c30+9QpJrJ2LWA6RAMD05ygdebXsFfHow699B3pTVyc4/xfVd9zpl+LR8wC75L7
EfOYXo77ZqgxwzjGgYMPBwrSTVgXcTeusQdYN4l9r3wzZIY/oz28LoNti/A49rt8
Kf+dy7l2pmt+g/jfigx08Qp95CJ90oNBtbYvP1gw3sqd+mkmBn9nY4YSolM5i3R4
jzk1Y0bGja4KYGKZh8nydIyqfLi2PLtjGuLYMxNOLrGXGvcg8NpsDMB0GZqNJ21e
e2/XwZV2wLFcwBtQvsROo+TioyXyl/Vopk8LRJoM3PKklrkRDaLP3/j9UllEtpeK
qmvaA7O7/12ik8d8zN/emXWvWEii258mvuZay7EPc+7LZD8g1xay62MpX6fay+7F
Uf2YS8ye6ap+U+qXnjgROoxZnW4rqSeToKtjPMuZ+dVxyEs8jlRWzewLDTafiuxi
0wjUW5tCNALIjaAGGgKcJEs69+j2UGrOOL9UqbxYcRghUGZSZUcybEUVhMV+1Q/c
2YScwa0G0rmyOQ/QmA+7Y/ye7KQ8jq1BAz7utFXabX35YXjrKpmgaoEwdgc5veZF
WoCQmothMML38bWQcnN57BKzaZWQZLv3am5AjG3xYk21XY+WQb1kVosThsgw8gwL
UBc0MQJWW7cM4jsjnq67eDUe7oIRbIC6y4o69kubiB657zWKa6EkTkR5yoM0z7HR
TTcSqypX1Jz5YFp9FK4rea+saq9DMansy6v+Iza0DkBwgEvhMcLgXXQNJFcVNTaY
OCO1/tmWU17vid3c3vtZN+d1Vbav6luXNe+n3lEA8UUEWfTNsXqs8kzgB4c3dofM
7WY7BC8Ix4EB9q7DXKvftIBOLOZVwELXwd7PHplxdBB+8B1fzouCuvH4SSr1U4DD
QjuiVSZ6wni5fWSq/mR3gR6NCM3211lCHqmk+NBr9X5vqvsjbn++VqbJcoxAqXyi
2Lys/k8cibbxSWLxFcT9ZehZaBSZ26S0gFOdapPixCUiTxzzcqbIcxyJhGva/aAd
+CPQ6VHq3vHnrzkeNuVcmeHyyciASt6B3TI+GJzXHh0KHUkFGmMLU83STG+KPOQL
Vn6TsQKtgj/Ymxdr0wSPLl/nGm3lBpX4Ly4Z9in4fBAx+mNU9NraEVasld/K0UNA
gclsAKtv4hMUabNfXo+ybE7FYE3WqR/gk5p1R2CnocFKzoX/JQsGyqOgY5xQMP/M
whiLOdS0J/Ww26ABceJN++CXG11l1eTT0dJQBt6v57TeOj+ynudfEkLEmd+daf/b
N22EMItxstN3QGBzS0DtXPwpF8pDD1bUWawelsVQJEh+i1JA+PMMXzKXYl6RQbsL
FxMUWBQZEexafF/QdUBhlOpmSrIsASRwPLrHbrMN4RqwgEg3ugU8QZSyoOoBKN6z
M0cbQYBA6F2G0bilC8rUW9TCNTYMgnBw0KCnCueyv25orIK6VKyqx6Hr/93tdxnO
5qwKMH7KChYyn0MkqTlFaXEEKLHWdK/B5jJmUXaHMsKD9QpA1M+nsXThGfMB0464
lUnVy6Xj+h/euXKs338l/NQ8cEDowy0TYalYNlQKZTSXTbQc+8YWTTloCYk/XCI4
CWiRE/JwfS8OpWXQPyHSo8PZaL6W8igZDhuyvS4b7Y1VA7OsXRF+vEUeqFvsHVoF
VpnVZfyr41GU28dVjTZ+tkey1Kdi6l33enjO4jbu+RTIHYL7HfF50kewOLh4K7di
PqSxHEB9UerBRM+tCYsjcEf50pLSzl0yd0QzDoVfn1DDHEVjeMonL9vU2Tkp/1nj
DBpZjCv27zZyk9N32pH1XMI5UdtxRu6K1d9g7T/GGRQsqotYPRbTQ+WM5h0ghhRn
19pzBThYUqSTv3f2Ru2cM/+xDVPZZbAf2C21CxEc5+eKZuszvzJ7MbyxJe4Pp8Pf
BH0XtCC8bj/0zoeXKkre6h6xXn+RmjRWLwmtPUcYTiGLb4deZ9rVZLKJeOE+y0Os
oSDRDmzVnxuTzYgF+HIqRbJ+1lZ+vuPeBC/sNtVVdw9v3PefgM1sw24GZquiyPoq
y2LtKugRGs+UdDC0IgWJxtRs2hqkj7rK1HOofaB1P7IGKwZ7aMhv/Ida2vv+S0Ha
QveXTJvHQPMMm8icNS31adsGsvytMygdlk3EP33Is0+AN8xcLmCJlSpVWd2T4YnW
t/Dfh/yl9dBbOchOmc2w0XK4M5ka7QhF5lfgMkDihMKIP4ZX7NH3rgZMss8JHVFR
NaacHD7we0g1gU4GAgt98SvYimgHQwwoNCvHkUf2RXAJKLfZ0Hzu1WOWm7Gac/Ir
HqWgloan/GXyqQbeyEL1PcbhFe2u2ew13chLXTq/AX0Me2g2rd4/aksbE6Jp20tM
PgLRmihpzyGcbgcVoilUHwikrb/k9wgOdRzxc03yePeyxDVyQZe8r7DmXM1Xb5rC
L0CYfMPuw7zFkneQFm6nV7RErWIGTsjT2obIihXPKNqqyFyLMKA1KmulddY6KHIz
/tkcggHpoCRWtkQ4hhPCkHs/eskPFiy2nr1gMrGhzb61V29VnWyeVa0YWK7oYxsG
/cs8XDPwNm3PskAaOed7xQXLwm5E6XxWT1eGyFadOkxqYq9HEtRKPCpPb5tQvRGt
uhjh76D5D5X0Zy7g8MUqjB2Xx6GsgytbH4RbmHUVKpAb+dUgco5UxD5ST11eQJFd
Lu8MK5ANCNT/GJ/AhBH09BJBwctoPtotfZdSyN+3WK/RDL/QYv3hIpLkt9S92BPD
7v+1tj8HNH2M9R3d8lZjNHP+N/01mG202BRAsnfKQsRs9HiBA/MfMIaZmy7aWsPr
EGrtAyusuSM3lHQqxv7YZaGQMwJlrW4UcskxeYQy4K/SUH3RECs+PR8sch5v75fY
07Mwa447UtKqsMGvCPzaHoB/A1+nx9trXyWw7ZcREJgdGrd17tqc66KFCAOFDefy
Z80lAsSBQ5qtFbVxSzk57wglOKwsU02df7eKjvftDSR0/6GfhzkSc5vE3vcVig47
js+HqxzeTN7p+6D6JT7mPyS1iS6+VjoO54amOZ69cnVKg1oEJv73s5+BTx0RHHr+
Vn/AGc72m0iOuA4IKghPrVG6wNatxvmYaLu/6Zt1FWQo9UB9n2Dg5gfAb8K91gGT
mvAWEQkwlg63ezUBdmK7I2QqiQWoFEXxLEw15MUbuRJmGh0sA4hbyAwrRe44pKOL
xolSn0sn8yWQwkgIK5/KEVM7bMOF67YJFruit+WupeMryC2BPzJ4lY2i1XUQFGPM
ynPzMxq1+2yugX1lrlyRTI5LIYA0B3PTCwDllyfUlefaxTCvJmSUW/HGsA0fmm+G
alokbWu7hWk3cZho/7hj0+GmeXHqkhkPZo4HGL7WrjXUeJUgBw0Nt9j1CxllM97b
1cdoV2WfzP6oYH0czXDG64ptpHF99Rq/iSMdmTThgR1p9w9UudIcRZuWrNDCAu2e
+WVRCZg3J8h29dGrcqzNmy2V7GYsV8a4PYt7RvVD/fjsmwG2EvKcvLFgo8KMqT7n
Olr3/GGiQTvvOAwfqn5VNY9r5vQE40dRz6Vzs4I1wHBgbT5cxubpLsteao0634bt
qy33drivTETdffLiEXh/CW19DlGh60A7yjpXiuglbGud2IWSjLXwkbVqshiu2sMl
JCFjZUyeTcBp9aZtI/zgAhrek0CdPzPAvuziBl8wlcA1OAhHqeWzZ15RQw8NEglo
3PfkEEY2r9phEx6D9C6G4pIUH2NPKed+edWkR1Q54Q0mHpVhnNYkyXEf2KXcil7x
7ViMyxEgnZZYj1Rrga9hmEPqkZAk//ZPvFP7IH8KI6okn54a5I6NuqhK6AkFKVQ+
FjFyMBnbGlnm2GIdaS4MdthhvCD2Qp0PN5AI34AXHJtUk++VOyrHrfgAxOPXKCLf
7f0yi3h4xS5goq+ih1khYNW1ZptueKON3yfjtOKD35s9usiJ6QuIE5ynLgpO83/K
WmnK6wt4Fjk4QARtOGUYdD3YdjidRPSpHauPvLSxzKExIQx09IUNs/2X2IhPjzbI
ZTomegnCuCRKm5F2VKRgojVR0PSMVKz2wKx8It++lAaC1a0D+NyBndhL6xtcfI9o
VT3mdT2bb8BKvMpOCRVLHnD+TSMxbXkkL3bAbkwJBcHlga6cZ7cVhfng6p9Kl10G
r1LzmWzG+1MDsZUJf8Y+zLg5Q8FITEUKDNF+wWnlTJN7B9u6A/3siEvO7yDxMXJX
R883CK/BgT6ywp3KW/J55tBVnMVRtR5iPwKQbI9qA1KE4I+F7bK6vFxDnfMO/TbL
SVDNuBif+2yRLTdNSPmRSapWryJGYvT6QP5tCUv1CRcVRHLtJhwg1g72S0h0YxlV
jDAzeNlPsk2yTMgRruTmDqUimyBWz6/Ktet+/QvONYhGTKl5t/bCsA4lfGPX+T2w
aRiDp1p7UMda/fTb52VbYab2STIUETI8CZ29bCDw6mk0SXQDwRsW7q9hVTkALfSP
EkqjVazuclDgq5xG1fI8osSqRcgn0ZURbThAH+D5RwmnbIsGRd9YiS+4XTsXv1vf
x2aLygvwwwbLUVW/QnjEtAi3Goj7hNY2DCsYgcDLYubCXOcuxJu0pF2451KGzVjR
UQWnPDhKfT7/Qy+X1XbJFmhllQicnB/vyCO+/ctYeU541VqlC9d9BsXPGX1Kc96L
wsGnkDsQiNI53SFnuteFPavk+KK6YSU0EjwCtuHSTTbaH6xaJn04IaSt1XIJS62Z
urb/m9RurH2K5Zs4xSXq4u300NyXMlWx05uYoe0o+Xeh+4NldU6iu8Oo29HNAeqS
6705mrZ5XaAXJoPp87LqTne/7gAlLl/Y+GdR770xRwtGsmuKj/bQzI+4+wSytvmw
payKcrOs9R+/NM+Pz8so1wl1kQyqxLsskz+tbJ7U8ZOUfJQvjlrdFqhTDb/YwjWF
TJz9aJ2yhD/mNBxC/+sBDvpknLg5pgirpJOeMCKpjii5FmdnVXYUQXnBEex/sCz+
Q+XRo2RCp7G23IGgdrhdfcBgkBUquE+71n6+EJ6VCndfqG8gGBhcTYvGW7uIrI/s
+7ARziWvkezWyvwSsrBEr7PTR7xZdZ2doGxhhGU4a4K9Maj2OxqcPDlbRT6SlZU5
uosulfGk6P0LuJzph/a0TvOsRkjARuLjxkMmB6lfXiKQZZ7TzPAb5x6Ww6AOpgew
F0iLRDgm1hpXctv02UZQe6crc4msPezYz3oiUfSpREeALZ3AA2XiyQ3tEhWwMMOI
QkBi4bK5NXyvvK4xchUgH872CO3aR6usbXgJ6nJP3AJ5QMUijtzVTAayuYayLk3w
Ui1FkI4s0bnTkC28UO4f9SudexRrpWe5ECafKYI5Av9MNeX9+B/H3Wsmg5gTBvSF
ZWytZJ/uFbg0J1I/oQC6zzgpapK4FIbphMKpKHJe7m8GOuBdaFAYCPJzKy3MUTAu
kFrwNH4bgtqRV2QhdxTlmSK97HhXPOh2xvi/rbyyqNAmwRWbTNlXJ6VLnqEf/CNh
cLbR/2l/+dNdeY6yTPWV5sbpXRefqvezIgtbN0K9fdNuKfT+cLE58Iicmam9SoIN
F9f+dIZEe4SI6Iiy0PCkyNpQvJyGyYE5WSUHGSqMkAgUeeltBs4y+IRBd/Onlwi2
50Xp/zKhLZm3MFcXs+kBcTaBHwRrKsAkoAogguIVvcYOCCHUqNa9NbXluybVDy9r
j8HuFO0UDTGXjDSdJdhbgYhg5fkXFr6vV0bSUwirSal7KW7PFMh8XveeWsoE1V11
pkndWOiQfC0squao5y6S0G6NbJ8oLQWCDddWcthckg3zPbXpgQEmGn3zkZp7Z7l8
uZ8fA8nglkaraDg1jTU1j0UiI1RfRa9n0BJkqxR4fURi5fR3CYBSmIk03og8hDwu
XdvQBp9jVCBAQvKV4sEt+qWbyo6HHblv9I+aFu138ROCQamxWNw3QqUBm9OXZ0kB
cQciMEHHadrIpWaXFZTLzC5JKdnRyWsqlEHK9/u2ygN8evu7r8oRxjAMvYmZIuCa
I9EiCckHALRd383tv8Z4HycDR9IS4V/P5orLgkM1dgQSS/Ag9ENZqJkJQJWMJg8P
W/46o7M4x0Zj7TIACLjSaFsiWIE1hVN7Dr0fW5TtI+5GC+O2p6elJoUrhciW8t1N
kEoh4Dbxe+OnHpcy9d7TODnfeTmQrSRYyAHwQPW2P0g5puikfAViRQ43hFWroUMk
S5VLwsWDdCc6qLT2OYRe+Acs0ujqnpczZ9zKRS4RDBLYWOxncUVdiezJtqLuZVQC
qGhIWipHxDQzaKltIkjePcJPDvssNuBGaG1jzvIRFyl/gfDUHtKNH/Yi3ouo5khw
M46lF7mqC4vXUa7NRGQTN7/w1GF1YdlmIoEDj4xSWEgpgBVV1GLNtaDV1y4a2nOJ
JCxcgWo0/gzYKLvAGKM/n2xw3njJurQQYnZUpOST4XPHvSXOuL6EhUzY8XSJgQjN
pvgBXQRPYTdqMa6RI4euLmeHzRmA5YVjJBXGZ3tlxm8Y/kjTJOHUPSvOKEGWJhkS
hgxeFujxAYIdXqhzsbEvy8ncYyVyI9d3ZVr+KN2oJ1GILjC5uSqrk0GQYDZ7K2CF
lEMh5s48gfLW/ikRqlLWXcLJUPoVU9ztNKROcKa+uD7Pja+Omowq4yMFo/Af6yF7
6KarIlyajYtl4j6oy7lfHNjRTGun5GHniCXbjXhgyNjzKSNhZ2p4mkK1WvuZYL0c
S8fJULnFVYrBRADTJP44EC/hMZPk24IXXpwbn34lObf02H2LU7qtMiyPg8TBSIga
E8C+nAWK6gs5zirdB0zizlQ7WE95z+09QlX5bhoQjwYfENibs8K95nxm3jXF30yD
CTbpC2NY6/oDP8ZJ11FYjzEihpwleR4qArWGD4O8+YkeFBw9ln4VcGb/R6paaobe
WgDfGeddyimIMlh/D43vWdE2pebL1hGnVpSwG/1JoaxtFNKQHOJB/mD2/Cd/j84C
iEx6PgwplmUWvSHLIr7FUYekuF0BpL+VNw6b4tNrTvHaB8gpReab7eViI2/yOvRV
X1t4CI/s4VKLRGHHjWdJZuUaVilAN2GIl+j4ntI9NRNXPvC64HnK/EBNU+1XficB
syJ/1/2gL0P8VkAc9KOJIdM8yTwnQwJ+xigFcZj33XZLZixgWe5eU+/Mmf3UmZSH
Qg57EsLi3TwjKBOXeuU9ZC+4XeY1AgJW4h9i5hDWBg8cR1VxuN/x82CqbVRVliWa
fEz89sEF+JDercr2qBld8xDlG+vIGsuqG9zaXyg9ChANFyqV/5/RjalJJ50nHIZ7
kIeIgAI5byW5lpgKzeb4wMaFVJiXtSOQJs9r4sYeUk17lCHawMG2gL19M7caqE3w
PJKbrH3FgN6NI4oTkpwygmBkhoQ/QwKu8CBEGLdlkEBR6Q80ZCjW1GlCUNRa9PCD
O87j6UZfTOOXTezTjJx3BjMki2P5hZu4CwDZ2rTXNlpuaHDHUFG7kwBYM6DuAs8J
gpwv7rUO4a31dDzVREf4Apl9DZtaIcRnPBCBw0k7fxemRfe+M5TxDacqRfOT44YL
SDezyW02l+0yZ1mYn6bjg69jAXKLcrFO8MDkl909dEl9DJhE3FWC60HLfpugqGm3
V9el9NstcqoODjTV6fzfuxDKtyrKapZPgn/JfH3S6exFa5u9gYKZEN/FYCgi91tx
/mWaOb6k2jZYZFvjLVF44bykp8JFP3ogIjxT1JUUftvhFPZoCoIfIkPsgoKmwo1z
6SCMpQUvjh/j1eX1RU/sSS3OLgYDNzy/ApAXtNxZ+NmrspOrLpR653WPAzI6DYhS
prNeJ4MPOq4KSy/X4C2mj+HBLUot5w5zK0BrXHzYk+OMukNLy/MbNljTJUTXDvxo
om6KWsPIHgVDgsYP+C4ndl7gNvZF1BZfJeZZMrypH4GRFrmbsVm7Bre9PJ25/nZ/
l6R0kRol9hsQQ8vqOBa+n60pgUUZRArzj1qZbPi26HVllMCq30cZXs3XKk7UJvIb
SBBap/pSqrLbwQC42nweOzLjb3tMuTKT03aFGg6uJ8klJIieSlWgL+fbsP8AlJWD
eWQTCX8+C6F8NSjbL0xJ91qPhrjW1d/AekkI/bfLHZ/Ei9K6pYoKTe5PrrgJ/c0j
Ym7a6FGkv3HLex69Ra+V4Du54fAu9S/i/DeVYUChSR7IT+8qSz7GoFMyNlm9vBO2
wc4gPmH7Fidn3AelMRldg3KC9wmTx+TEJREXwKhkZDW+UARrTfh7Sx40Qk8x9UJw
j3AiKx1EPvvXTmBeRl6GGqoDVxbfhhLkReWpZaK+i8kRcbaCPyVwUvv2smctejt3
6KDnkbZkC1EM2U0fT4UEuKP9H0dCPuVJsQHkegDr/+5jbt3DozRhJ3PvT4ETGRQC
t7JXENm4kf3YRoAV3GlbWoxfTO9PqhAa1zv2UjXd67hxqiI/SmltpkLg7hrOIQpf
AVtPoLy2+OhvKAG/mE34PswxYXcyJTNZujQ3Pom1AsKF+XmPVeKSh++m+uN15FoS
o5IHwQDJplUnrH48CGaI2WAPx9s1X1S9HSS2FA8eLe7LUC+2fKj5UG4Knyom3MHD
e659KHb6FMHMWM/StbQUnHp7ZQdmlU2hA80QIv6io6fnXGzjqpZzuW5NAq2dcDhW
+dnByz5w8yggtX/cwWvI8ax82MV7uv8jXGf3zm1K+od1961UYkY0CW6sj0ovfbDL
dmr3W748KpxRAjtghbFZVvWKjYA7at0uut9qncAG7lJ+U63MEnTf/ZK52AgDpw59
A0SLi+bNVUrOKGywYonMZh9FnSAn1T7fWaFNK7I0CQFuswlLTD9nmVNWQDhOJmDC
LX4VU5j5dKGgTNKmBZZloFRQgTGdqsmzWX5CkNBHNZaVQct+ysFCS/lx/DWLF/Du
glLpkm2PAbwv2rLskNduiQUz97asBDcJFpbqviADEg8XawKPwF9TQIovefeTQkQS
O7t/WsYjBiaL1gzik+UH7AkcOUCaqCcnmYHqt95WRkutp3H0NHDuv11H+j0CEDop
UUR6nj9DwszVIF3DO7yoGkOY+4F/vz59uOkr6sBISz988hJ1wW4aFRGcpM7jDD1e
0oiIROr2D9ZFaNzmhRVyUx6byWGe6wujnj+mep2sixRcCu0ANlGK68eh5caz3iYt
oxKBrVfAkGP/EdprDc7rsy7QQfw84RoXQsh8Iv8UyejgsmcsG3QibZKbhJpfL2/x
vsnOqZQezYH1t1W6xuxKdFOgY6f75+RP+29XzSqCtp4BHa5InxgExkKGZth4vN+A
0jdXCa8o1dYaNDhfemvsRQCjcfnCqUW4wrX1SOBIbsTwn15yDu57oRkYxFXP9vfa
GPYKEeUZqEloAAbWAE1rOnYngqX9fKoyFnQ398Yzmlgd+wmVzKDjiMKbxosmnHih
vdCfZQOVl2lm/QMkhklj/YrBGIENNw8W/LJspws5Xmhix913NuU007AEalNYFr1T
ObQaMcoAaX/0EXjxLOmIDbaW9lEDf9973JUf6QYMmWFVQCEOVInkNVX+tbjD5hJZ
vIe8Z/+SvQmmhocF3xt5oLuIj0PvMP6KIs4FAM4FHYMFR8nihN9hyT2sL7qs8Z5b
2mfkQXpTDRjjZhC8JxLhL3uAjtB/Wh3Y6rD2cHerYwPIyvg0QIs/DBcKar2Djhzh
rwUDaEXaxtJ2RzV43QT3AHSaEQzX1YCmiAiqbojG7d1mR6fqAIZxfE2pn/NLwVjE
23I2qso3nEEza+Q1QYTUuXqkgu8/3BMuHNTnHn1gCHqD8aiGl+4bN2wQxxzMlDZ2
tCrUCUYkoZLx35pUWRmAXfIvbYpY3XkQSOjlcJeb6ef4W/+eu1DhGMQ2ivYDuyU1
SHH8G0eUnPeov6ToS9fKf/1A060G68E2VDLe81CjeJ8S4Dlkpn/q+1DuP4FR8rYT
PjU8LX/YZJ4qcaJz5sGymMOuztIFyH+xqaBRaU4sMuMzjMETdlda4ZNN5E2mS7C1
nGsHV+X6BLQZ0lyJG7N7AY85rO7Ki91qNfnDZPnkNzicCLEGwEEI0i49jEj6l6Dz
ds++xcIQXDM5+9MvxvzxtbBnzFXy66JVu9BG8bj02fZ+TqR/JJZvc1vHpaHEOaCc
in67zadzxOr2n7sOe2LXDwHiCfi6LDPyobCJOU5tpG/36AI5Jtcien5ELBF/0EA5
YCtrUoMjvdTgUjtAIOp9NKvtl5v7xHKSulcKq+R6et/LZVQokVipcH4qNFW5NPDD
epOVcU6o1Lwmm4baBycXO97NVeZig3ZM+YIXdplakw6FPAEWsFyRWLlXb5/Y03Xb
UXpT45GiY/hQgKAxYl9WfHGP6vKPI1KLPjy/a+0eqM/HGwWdRIYhjbxvx+aGAZxh
RWo1tSY5CJ1Kyk4cUTUmtrQHR26jM6WvflOjplyHzEUlcXfbIklFNgwzhpDm9udA
n5CoP7rtAkjSC+V6KUL9V/jGSFGdHL23k/RprXkB8fRF56J4L1niRBSRxp24LZkl
BfLP1QF9YJbDtVbfQI5KrmRuYOzwglHTS4Ab64AfCaSGsC1bf6gIbkBmFM0CXuBc
+GTLg5egzskBnYpP/C3CE6fmD8mpI6A5r86lPQHrNPc6ByKNymCaymr9CKn2iyKv
mfOE2BR/zxM93bITcbkGxX64WS6nsOg7nYyBVFe+ZayyfSxEO5REWr0ja0NqCfHR
tjgdcuZWnAjq24EU8dApbfXHgF06Fo8wvjd1MhLtcjGtcolWIrMdlCzdiqpRI4+7
wmsBYmxi4nnxPSzcjAdjvIrHx/Oyry4uzL4MWdrHSq94wuPtnIXOtXHNTpjzfIg+
WvgkQr1vq5fFHxpAX1+1wAnKX8JAIuBuA66rFyea6MQc3jqEOiHF5nqrHrAn5EAs
Q2cv0cvucmT5l5hza6Zdiv9hjT3/USIeEKeEMJfUBS0zfL0qpiifT/Yl7sp6w9dM
3SUPC5avGzZXbhQlIGyYhkUBKG2eFlHahmOxxVJvfnK5Uh0kw2TeckxC9as/cIB3
KOCw0Ovuy+foJPyD8ekPGDX3OH+doKMcc8YgiXmLNJyFiwU6qwatJErXC2u4VHyh
P9G9VYqueKAn9ZaF+QfUEl627Q8SisAQiO/q7jZBFPwK0XcUAAwlK7M5EFyarhRw
e96k+Uho68cndgNfTCrXXG0h66FTBHDo3kieHvNi0HFSFIRvg0BYtQOB++Ul79I7
RGrRVxF64YhrfTcrlrlfJaSM8FgDiF5FwOSCXwjQ4mDgtyaJhGxYG3sIrgEw1Wja
NJvugK2/ALpRrojCs3spGKygffQ44NUy8/5HVb/Et/v1aADDTQu0y2VWm9LpSqta
BS2zwHX0VA60DFQig2kiDq5XbSB0qhMgeQNHHUJT/WD49NLtg4ntXBmAKK+0yvCc
5ubb1wWwImlTcqaRCz1B/vojbgPa7HE4pqon7E6YHOaLohglucOlDn84jRKT3+/Q
EajAWJfuBpIRmbGnLu/SVcdpRExQqOePYZfKiF+GhTgT98Xp2GcIZw/gIYCD8Lm5
8gtqudiVqXiyjbUxae2anVKutHi/IFILae8EwGG1cc3oKdTT5/8Q+KQHZ/LgQGjV
WPcqf7oax77pCfSHU6XvYn3Tk8fdRGpuruRcWWyc/q9aJelMtFynp5govm9PZaK9
mx103tyNfj3roOmUYm8UwBlaEDR783xhCmn2nne4LN1ynqFhhAFShaq/F8hOTkNp
JsbQfzWw8UDKh3ZcUPca1ymzPfLqJJT6mlAIZSMhjcVaUFJaIr3priIk7E2QrowM
+53buvnF3f4WD90pxduMjiil9kws3pIW7B7CxUKb43l9LA5teopFHJLhsLpx+JDn
X9b3aVmJndHkigJitMZ8pW3fFPS/6Ctg9W6qJJt3Y7KOVLmKb/RXeFm1a//cGoC5
U+WY2atlMfHIj54JkFaqLIunbll6bZZtWHpRfzqKTxB9IxWURKKRjqPAEwv3BNi8
Qm7EoAn+pDqqxAoM1NuFC+fJmcrTrwZpHHhaI2giYLNhTwEBDvIj5g+G994V6yIv
Xkopv7upLMYq+lX8JDMtdeRkqsvVUw3NnVLVzzl5MCtA0YEPmMXFA2ADLlClWiuQ
YwOL/tueBCvLWzTAZZFXITe1ypKHSp3nvT5kYn9omHsKv67tcjKH9QX+wnlBBjaD
k8FSTvTT61kAUjCQ/LEElGCysa5IQ/w5PKoauZPM53ytN1EYL6Z+7ZIYE5dS0rl+
k7xb6AgIHHWHHdBa1vvA180kxzKfkEnoQKywubahLFTiIEGqHIVVXS3yVTa02ERb
V+Qn4BT6KSVAhO/DzsH3RweahhzD47H26O5x4W3i4vmNDSTOiU6ZRrwAUiNRh+Qd
O77HUNn8c7k66PCx2OXGqamU5ulivKzLi+5Wp5RI6mhe3gYC2NUxvceTkU6bY7mO
2jCbUbaDl49CWkacBY3s05JYl6JcScYA5N6BtivWdYUGKNJir91VNHS/uf0VkooC
VER/gVNN7D9/RmwCqOTIv66Whgb75cMXK/L4pxQtPUthG8ARW9jKq+kfj6jxddgg
Ec69XWADhlT87GxFlISz45EdgsJxya2ifsL7mJeZBR0h6B7P3lXCf0nR+cfnIl+H
FYrdcGBGJk4FzMMG29R8CX3O1nJdsZaRDGkGtLnlTLVTVicwDlt4VkuR7GwX9QM6
YHHBCCrr5wmTBAm+S1w52PX2jVD6IA1lalFBKrMxSlxns3FUPVNMmHSC8aVWI6xT
D7Kb0d4Qv9opXs2MwnP16/HVUHp4KYCix6UYoYGzM9WTrosrRk8pJpOuxlQHS/nc
8ta0pY8JBmuVrVg51ZgqzRybhWmXqMXKUWI2cycWwqGHTUaw4q4HtzpUtsEXdB5D
IW7iCMZ4mNJZeFSCTpDODawOr+pAu41Hu1vcr0F5IXxg1NnJmYxEgkMK/guaQZ4f
Z0d2o362Z9YrEStJzeGGFAZljZsjBWkWoJoM8XND8QVheAQnTCQ/Q+QyCLZfeuEY
DUfxiI0xILp79laf2SuYJG+FmEbbHAtnXrsDqiun7zXWeWTuNjJFNFGQ/PoJsySN
3V3kdB7NSX3nhR53a6k6DgE3pL7lfSX+3nmbwKUX3NxIGgNd2qoweF9Y4/bKlmED
dpUzTOi7kolTcrPfQ3muerrR9uSjKgTuByBdhz38aU7W+9rn0RJUMghtRZe59TR4
bJJ1Gl+lka5EPA+0e0LpgUjQ180Eg1oBbfCuHEKSgRWa6IFVUAqP9v8vLI+Vwt8s
ipLEVzC8+GakvIXJU2ZXuDAL2wr+a+MyBGX6iBHwUFJcglSRE++8GXtyr8w/rx6V
3MxRKF4khG9U2x9GEk302YxUJX45WD5t7orZ6XQVo6NRi2sq0QAAzVyAn/1vFAjP
b8cOeEA5Rh/fS/DB/Iy+volvJlGB+ksNH2BYxw6E1oyS8hfGH59zeoV64ugv3t8g
Ybn7LAxpc+FfKZVDOlWWHFyHPc9ihvum4W8DzpOu5HJM+3vPAW0HYk7+epmdrYS+
O/tETfMB23iZdZERRmnu7RVB8NxboEUYhLKcRL/wTJRkOox5OtmRKyGr43n19Px5
4nsuMm54GmF1wg71cXM7EjIzuN2CwHg8fcHXPZR8VH1v0YnemnBShWWm0zWvkT4O
xdOykZNzzDWiHgjx4HHVg33mDSankcDmqCgtKqvx399kxLBdUIz0zbq3S587ajbG
qH7j78fWkPbTIgD11/5qHFe9/C5qNieT9kp0hnZi2wCaqSTERReGXdvURPDOosEM
qHJ9oKfuCogD5FTSTOPVITDijlxMsAyhY7rVpYvibYqEL3NfUDWKy730OMj5RT0J
qjvjjeTKG5C0bhQQnKy33oCy/CHyVumh6vAls1HAp1UzWdb8aqHSROJp8Z0cy/uS
g7WJtycS/wLanJ1oykjBloFOd0ZlTYQ58tXdUFKg9G+75iW69nb/uhpY0wDn5hja
DpZ1EVksYiR1wsUpgsIsOiDsyBPkUoXU8joHm8r5UIzJ6o4X4xkJANHLOoqhC5aq
xfc2I125q7dN22wcRjZmryw66AnwXrHwHnOLzONUz6BEEFPpUFwARuxB0LohZBj3
cVMrwx4WVcD72kTN7A1STs5XRksVBpTilPOiosOms8FJGGqqYnfgiZc90/ic/T44
CfQs1slm8H9MiBqR0HvnLZi4P//lfocPnxGfCKXxWEGKXFU7783ikWTNDOa4lcck
Ei9g6j/ZpD/N1m3O5mvAgz0SiEmXc9/9iY/CP5WWXluJkWs+WCYhm5p7H5RHZ8Gf
ow7j3jEE4UhNLQApxiMglbtcyspeF0MnlLLd4YVowlSNPxAEjX0KnsweV01uUj0b
z2VLAcEopl1PpiqpjSvyrLzYooXMKZ771jyarZMNGSXZSV8xQYcN7fG050t8Vyo7
sZphpXkFbvABZoeL6oFaEDukxVdvvaSP7LRjAeMztJyKJzsFWorsIWMDNOhSznmJ
bpWxi4SNVAKScaOiAZKjzaB1bxhtEs6xpUSV5chVmI8EXKZ8eCiqOISR0CrHKRLQ
yuQuUvAgLnmlrSTqy0NfSq79tFE4kyLmOeFgJ84AFSSGViGHvmLwew8kWaX/1cyj
odxZ2+skrKTtEu2qyC86g2zejiC2QEPWNSsVR6gU+4y0vM//HaUcMv4JZKXR9Naz
t4h1IOvYhF7AJ5H4CeEM+VqGzZhx1TYqfDzGksahWJYbNRoMnXBI0qa7XW+jZhHJ
VyYFYVvFIEJdUu1fS5zonLa6JQo3Xbelk9FeuabTdky0bpVD0/WtQyoO3MHml9Cq
yjgjzLjjAWEg5rzGZcg6K41hayQJ8VVyQk+RpHdIpc7AwZlThfJ3mkn9t1Cr6J/Z
i4b51qr3UcV81LCyYtGlady2WwK2Hlbpl59gVewnwrgAsnc7+GMDymJFM1s8XxQC
urBF2CxtYo5xb44eRnHYJeT2VpAzydIuHT0ODgA9sdAyiqfNjhi5+VYlAhuZdCVg
19JecoqbOK/FQ1MiMO/SnUuDoMIjUBxEnAXtzMyyWl45UAmDGCNyyTu6TcRM6/cf
AQIUhtOMHveWkeJCiLHkLOjBnfeF0VrFPI6fYSW1KDRpd9iTuoZzDty7trYAXZ2M
U/gjpb3dmCpvumYf8KccbWyATXkik4yoq5ZpxcvGS+Bn/8J69b0+Y14gzoLx9HjY
DxKcP32LANTvMPbDHKmEvf5boh82/gULNAiJvyyuLkMCo7nB2GgNmjvFN0IcrGFU
67/j/6dGKbVnawIjbHMbpzWWwHGEMYM6lMw/0PJWZKgSFE9LV/On/MIeTKI6wk3B
NXC8WxTNpaJODY2Bd7gvL2moSGQbCpw2Q3Hhm+AxMWFhSc5/pM1wahLTOYSy1ZuA
jGymnoWc7qVAEekp0iUMhfXzOvUSxtTfs8rsu7QmvtGjTUj9eepfeqNmFJxH4VA/
jrwybNGXzxCMChWusbHwuzyGh6VuUqB6jVVDN4geVa5tSCO0Du1Nol8DNVZNLE9C
gE8s38/G8sv7KfVNOyhTFrX25Unn4YG9JTlA5cvYBwLQFlNmZ5y30azWgmURJBlm
b/s2vVMcTWjqlUvfJpkhJchq9xcQlwq1g57UfUOGJg5Jf4YjZlT0Q077IIu7dIz6
Ix26nqv3iXUsEgICsi7ulcFnOVEVwvkWuBRIFGq7r6QudlrK4ZDZgPxH7Du3tYHn
6uUnp5wbMA43Y8/wnGRuI5ieUzlBb3+3HQBLWkRZTfMYW4gDPYpOXqpeoP2wnrcc
LNBv5DAlOeuFTQzJH+5fD5qXTQABxsL7W40zduyH3+hQVRzBcEwQazHGhxWxOF5H
GumMRxg6pBpaxrdVW0uYJxRRpRTOyAnYzwcjM7AJ+Zv1WBrvzXC7NwIIa0Q50yHC
1AvZ+WSl1jtTBy6vRtQH9PtOPvkaNmegvwFWwW8r1A6WK2LUXd729QrD8aA6DHWK
siWQhpOIdbVmO/ZoRYACIo7DlOBWCFeE7KWSrML1whOEOSVf54uCErop9aKNkBSH
cbTCJUZOL+4XpyNyJpNNelSG11LDGPV7CMncIHUBYc1aQSdq47lhbiA10qlK3Bd5
PIk1lgzYu6Zvx0kRMnBN+qjaGeP33FkAxD1WnPa8A5hLcne8Z/81LavfFGxfsy9L
+IYkLrZOXiCnZ1O3ByZ73o3UgeSd6ttZBel3raWC1cBAY3hXgZbN4MhhmjrbIFi8
lPdfi8WVixbjodiIsbGDjWD8FvY0Zr/Abt6h3DcB2CB5HmfcD+yXiK2pjXgGefzy
8Zu9W1Y3vRxs3psUxTYFfqhaWGsbVCzmqf+GxtQ5my5wceLeuyim73Ue10/v0SgK
M2fG1pbA41jAkK8n6Inps42nKEXIgX63wujI0PBcE+/DUcLcqsLL732THL5i1ckq
FG88fhe6LmacooE2yvIcJKP1ihvOf59u/dAKnWmo48cBFD4e8f+snFxEbkHjjqHF
Wg7dW4DyGUFKLhZPKzNIWN0pWHg/eaN1OFfptJbFvXCj7qLCE/9bsgNQWnqW4hCM
dRyvzb77Bgy+Nk56OL+l6fVgGQn+lOHXUCglQPcXd4peayB6kxTcLRS5DKG6sHc9
2O9x8EQYVn66STw5dM59vxc/2S4w2KGi7OUgFb2H7nYJ8RspGAQrdz5btKBUqLYu
vEZqO77DlbpJ6CslmscHrpW6cb2IrYZiRfYVYrEPNTfm8LawevlOzD48MwHTOjqj
NPcBYmp7UMzxRoTJMuyErytU2u198Z47CS7k0f9T7/2NO/cB9HVXkhxhBLAFiiLy
pZfz8uU6RTs66i1YGOUw2EI2+mik6/P+rkWAki+7C143n22fY5sJ7mQq8kVo0bOU
3g3WBtn/mcXCqP9y2o/nN0hfv+K4dMoYrOnRlF7jCBVD7JofSuxUPRJ94owJEwgv
xbJRM3nmY+3rMXwVmUHJlhvy3HuiUPhfBMCE2k4Z3rCc4xdc6FfwSJ3uSQuxBgcN
xx5dmf0LXkcKdOa5YwXO7DZh03wdAp5WVQvgbQHqI2SvdpsrFM/AbMI1kzgx6SfZ
y1g6/TGfVknffqpaB6mL9ulGHLA/ghJLi6Ueh1mQkL6hBASnxZOfBhqa0W/PEvXi
uQl/biDeA5/GfPQ0GhE3zu1RSdlAAVlzZSlJzFG2af3m6jQS0lCIWLvjAj7F5v0H
O5Im1hJQiOpoM158e2y8m4nE0e3vCvu8UA7UAbiIF2eo1o7Cd8H95xSMPIrhyfDi
ORu3XMyE+i1WqiSQj5xpcNRHSrQOxGATsk1rg66VNGJaYsmzES6JeAo2gWAn2NAv
SgZxSkqdKBWe5q8l6rcsm7N2O8p/IBAuwMr5/Yab53tyQ79rN7eI3lXoI6agnKCm
B+F+Tb4DIqoutxUDipDlb4qd4ui6wkxD0OfFjsRviRNwHF/oFXUshB2fHglBk0Ll
9gU2cms0KgjwcH8aM6ARwcxZSryHzmZPxR5CmrxTO1wEcrGz+MiAYOD2E1yeKADN
JhW0gp4LcmVoAkIg5x6XJC7cHxnpswvxNgYalbZZoJSS1JkN2byIm+EzMZi10IcL
xkSDu8sGwWOCzgOUWiTrYHKDPB0Be+kHo6rbGtoMajGY2KaUnyIbMF5E80Uxrjpg
TG3S/Xok2Q5ehkhegvwSJAg1dtStVQN0nIvFIGCO0IZA18Wh2fiDvtew4jWRMbIk
lQc0QKnQg/1Zjo0KkRVzfxEzrhy9+OF+ywl7d7RRNnZGvv4divgHoV1wLS/iCKC2
voIXuqrBabR182zuKycmytZ8AfiDsS7BDz+KOcGWbha9HxiqYUvt3DbaBuGoGciX
FjbtmkKG3seaUcvqcTPdsdviqMtQ2utbD7wTA438RJeszO/2RPX8iFxMh/h5dtjv
LYHFeCyL2pzZoA+mi78NxuXR3TvbcMl01RCZ4i9tbunVFHYJ5qUlI/wi809rxggg
RhvHoY0MTQiJoARUWvCkZcmVLtvMdAlaww1SiKm73pe+zKD9nMUsO1SAAjNcHZBm
MNPBphZcSBkqkaxkaIFQLpgcdbrb4GeCjjVqiqiWzbGjs2JbngYSelz6oITHxhKQ
7Dkp001VhDlNpHEiqa8mIQtqaYk7OOiO8gcOpLdqahuP4pM44D52j3b/7G/cZ2Nz
m/6hjtf2qlXG6zpf0gL/K/o0PNnQTSkT8+CIxgoYRN1WKyYm2NUrVbpTNbo4q5Su
DCD47mpKfnC1AzxEHoFIIu7A1+mjgU+lYI0LdCJM04+La0lkdAcJhj0uGWzzaxLS
YhccrIoYFQjEwzIjt75BQzAJmVAVAu9eOHSHJF89AnzfCnxqFJtKqshM1dvHMuOJ
2TNGg9+igFAhdSqS53bcxkiixoYls5LSYpfyHV8JnbfHR055+10IUT4KRexBt4Ph
D1QFh/jIDbI1ZgsSOl4vpPT4SERSvZn1b6r8VcMsyu50DTASGeXs/xiStcWiCHlQ
ppUAhhjx8jVple/8KObZVFsAnpkhTNuqPNJCvXe+zFqI7jALgO1f3eQ8pEZmg3M9
fkFPvbFU7IA7qYGpdsOul8XNAJ2Lgfw8KlIDjNUOa2q0pWJXIWblYxAPhjGvmCih
Bgyk9SGyqnm6Pc0RGtVPmDmQcfbldYSyd6IqIoFzyGEK/UZicChv4Q13ied9FXZj
Xcm1kJzIQj4zjgaua2kukUk/7noP3YEQxpxDzUpFbeNNOSoVAMTlQOGMfcTm0ZIX
tV1gipW21MXuYgQPQZo5o/V1+/i5rqXo1U/mFKRqRYu8eFjcn3YSZKiY2QZqJhug
8Oz5GmKGeJvJ3r85FOKuxMi/y8W435fwv9Hv623OkQ21ZEFByyO2zBfpqUXUo27O
KcO2e8WRym6ChF3Y9NW2PO/GM53IA8Yhii8nXOnc7WLH08jAG8C9gOlL7mVSNUUc
uWfr9AzELx7o2nHJgZYKbYhL2oXq/g+zkCX+M/FlxLFNHXdpyvrdCKWT0rZGEg+T
5qE76msqdprdjyI6CtLlU31BVARfWY0WwWjaGTfNSc5SXgtq4pL7uHav0Yfatsy/
MKMMrZ0vSKhvsaJfXyiq3mEogi2i6aAWfw6EKYf1vdxvAKoq2PNa1vIwMqu2nJ4l
KMfNwml44BDhYdD+s6eaAU+F0bIf/4vrLzfmAxKaVZsHiCKBXn75Q548E/I32Wuz
Gqf0pYt3EB2+GrSaYaxUUlUt15dOFm/kh11IeO7vvy/ga3tqa263yBLu5NKTRv0Y
EvWjDfMuxT2idq2malEI/bw+AKxWQn/jYLGAAnhP/5ZWqWHWcJee0XDCEK3QrL4F
P167qf/hMxR5qRZOJXz2ORpTaw2sfO0Lb/RsLz9csMYo+UE7K35Z5Ob7ZC/G/tbD
5NFerGBmSqflGNHqoNiB131nnVfwOIuLjRhm0IhUCPwWy/FxT2IPGzSrCwQu6zf8
ZvhTspxpj4X06fuWYdGyuOxsUY5RGd2EPlGroWKVWp6B1ay0fC4zt81Wk6Soq82o
xmWIY6PM4ViXxSgg5wINdBxGt4qWJgRckFMw4N/qd/bBE15316MrZblQ8hm6ed/J
R/XZau3Xk6nGoO3MKlrGAWBRTkebeDw2AqKKyiQNH5VspIjuKeux+wyiYTct9vFE
IXy3imo2azeMZ3FMOwOaZHK3NvgrvPMC50USLfQ9WuVFG6lgGcBrIxkoCiZBxcAH
F65hvOQsjbEAVTSuv0IuIsfrvfSMT463oRDp6OagsWVN8py3/pB1U70AcVsfBKU7
hGzm7O+Qc+3tkQV2w8PFYwu0soj5wi6UXPdEEtA0wSmw6RZcK57eGTkqB91EmrnX
9eocKle4D41KzWw2JThRD6eBV0xcErS4XQ4xFEGUYzURtj8wHvLSDy137JZEVGKO
A2zBXy6CC7XiwgWrd7zxIWXKAk/qwuDxDAQCt1IbmoMwsLirchyp5ock6Y81NQp0
2xdaJFgm/S6bOz3F7MKexmxbw+aVrlVo5z5zEmKAErBruv2bJqsnHL4ESN7FULqo
XuLQW2a91IkGcFcG/gkp66vJ3eIEIUIVujfpAp90ore1xanv3/nO1uRxnCEXFmZy
pMq0OgN/5FQ54Bhb4M3GL9wXvil5ktX5m/IKe3EWGAk3WG6RnAsucEtkw8eD0T85
vz0EVGUEv4+ilT050hYEDzNcqQm+0KjP5AHjIVxEzD8P0w+i5pwkIBsCiRI8BUvD
xbVvyVIEPbm/BPKW6BAWYrA1cj3JTfQD9N2YVATbG+4An6/w3pcSuSUNv83sJJgp
lZQbJHLP8h7uIqfl2Dnp3sb5uHO+a3UfXRVgZER2PW9AuP36NOvyggTMbskyeBWT
W803woOBNEimvsNhYU+cWjeT53OP1H2iI7eBbVXFo0Gb7IhdTeOWtB8V0j7i+iLr
uDJ8kzG7CMUoDE0pdNdMX9khNVgC8yP6E3bMbG5+dOnXnvPYuzSy94L/VUjOz2jW
EX2CTQHWSupDvlzYAQVu+M3r/Mie2vLYh6JhQ/c9STc9XnpCSU8abI/uzABDXDMT
W3y1w1jxK1NpxajfiO4aCiCUwh/ghbF/dG4jnRv0ZTbNIzxuROmjm1onSeUz3gHQ
w5JSmIpUnvhp+nVrCuRiE1jCYS8Da7L30TscneoZskK0FqLmWANmboKViEcTZQjR
R7LDm/w6SVpAoSiLf0kb7RGGKJO9CFDTUHhGnwrDW7IT07k9U+NeLnivhY0hvzGA
N2mdo8xXbYzF26n43vBvbNuxp0zTSptxoo4Rewts/fws/3bOkxfh3Nb4GMbK2Pfn
UT6U152/M0vFbqsDBq23B1Iai06YYgJaO1kll4/dyKcBoqyteMswsxVyaMY4FpDw
IclkJFpBTxcISXuQ83EJBdLnf2RfKN5nBzDhs4PjXrzmB4wUynPB1O9vuUBOOTrq
LJuGVINaZj84XnPQPC+Sh6SRFQM+s6ajd6kwbfLaJeOEbnJHo31gAEF418yOFV86
wzbGbtMACdef/tOQrOdrVo0FPkqLZqRCaozxBRU8DTclMOxviyk8aSpozTlmO1nC
5prYFY5zM+Z3CAT1NHEW+lzG31EXHEj35vMIEDSKHIBiOnPLVVJAxhH2EHyvIUJf
VPw/fmScG5XkBolJK/q3Qwkp5ziiJVnhgP+pRpn+9mlBAdO+fWzTZ4IRPCMz4ULC
+sYSwH7Bq4XXOKc2dITj3qnyKLiz2EBvtQcJmcGoluQTNYbJ3eExF8pBEalbgD/v
iFE5SVp5FnQkbacbmuY3eCy/0qjaZfCWIgkKSDsqmfs0fDHKJ6saz57wrc38/gsm
Ng6BBDL3CMX3uBnMkypxxUxYLJodrAu4LBncwG8u2n0773HssAwMtG9IAQNr2ZXQ
Z5S4X+o8HjBs5yBBRC2B19mKqq+2QeO/QP+HPTFeqKBEjxA2cy0hoiaI2+6TxbtA
PNDHsBqS02jGkJddSXTZdsuC8gYgzRdwINUpiFVMnNKPBwQLMFH1k1ysRMD7Xe4q
yVisOvmy/6ynkoNHK2qEcU8BzYA4J4648T8LcXpLz04BWIXtIs/PKKFodSfgf3Sd
BUCYQdUryW+wfANdgkNj71AOqL/ZGekyhZdbaGjVm+RQkQMkkGqs8GUkcWNlwbeC
u5HSg8atlkYDdQSLFEo2ZTcrr6v+G9ARL8/4avjDGVRgdG9FDI1P1NNwRJg8/rJD
SVFFIfDx9l3QzR+FEocWrSkt0zs3vXQuS/GfCT+3Ph/qKjQzfyvkyAk3s1sVB1Cx
442vwHKru7Hnbfi/M1YDNiAWbcVHY1hgCxq1WkMw/JlgEA2JJa+PlBmSkvUsK3uF
ICqIVR0J2T0oH39G0jrjxwDJVlQHZgKYpkhDIYDJ/AQXjnnbKmf8FTfcRF4U8C6t
IvoI9zxwTO7SmzRAjSVhnnOyFO3Kp1SkuQfDVV6av5iVsnB6X/Zc1v0OTeDR1aYz
v/2ii2jIUtfuEc+Y8fUKOBATiSrAeCmZA9+PhxYGW7U8nQp3lz6iyCoZbRXTMbmk
aNY4x9os3wS8nwl8WAHjqrTnxXfIBkDJ63Bu6WeuDg6eMV9PVi0FhbO8O/IDr3lN
Uf1iVHxzWRuehNe+Li3jC3W0i3JnXAAnAQwXmeiLZ6CRgiiGftFbhlimuznEz/xM
K/1TpDJYZJGo3DWPMMJaV+Kv/7SRM+ez44x5wXoelmNtgZlgi4KlIEXs9DNjdiyV
Sn2dnKWu+jzOACU4yB0U+x5Sksq+eFYNe48B0toKpGiTN2TF6B1veytBlL5d+dgV
/gird7XVCqhPFFkM37Wp0TVjxoD24GGPs2fsdfiJqc5hKJjHuE58jIj4BJIEPDPF
ivqVKN+GLoZ+wCDf5tysXxPvrMzBNmMoDwAsAPqHUuKOlJZJPrr/iEStPIykrR+N
rmM/16XslI/QBh4q1aoEZjkP54L0Zok5vSWX1pyTX6rI2mNPFGDOoizb4Gxtf0Q8
01C/lBl2e0XEBP8+v0gX7k1v6KI99qrDlZArWTDzrNBUjDbjGqdpgEj9NRKMz/YE
itEuaMx3L7PpaT05FED03CTRu0kTpeA5tjRiIdpM6z3W0+9eJ/TmJ/pq5O/wiRzm
LA0ElnblqyOPg6pxq17CT8KfYgCOh2aBqDsvwpDBn4lCYiz3GR2Bixyc4ws1Jjrf
l/419z84srv7jiu2KYOydBk733aKLOO79ZYbuoDkq5sMYx72n3H+QAHFC0DyN8m7
f/edCNUfys9072cxlXHG/jUeixK4WQXnGTwqQsSSH2eYVXHRYt5z02CiQWyyfu4e
fI7mtfb79lDGgYQARiuSUYwi1cdXjd4Qcr7hdjur1WxpGyW/dgCWVJV3Gi1hXJiF
j/8gua0PJgjASQfsIe2TAnJkH3FTHvKaTArH5EamKNqg7EQ9Y1p4c2irPR8hVl+L
iXZLYiQpq/re6tq19TmrzYG19rFhggfu2gXLdFJZwqRs+Ql8PZuUWmBlev+maB0R
fqnqmXGYf/GbxfUectQbM45jAAE6R1GYz97i2CzV9dN18ekZO+BbSREs+2sOh0XN
mYEnYSNtNw0O5akV4CcqAJQdF0fT3+X+dsN0zLTXItnsa6+ZUq2TX50Q/ZinNrLv
mugC9TvoWCGUdDXQTebYDAgtTnI9uqF8AmM8Wa7YmNl7zYEiI/g0OYqv3SwKuzo4
kMI9U99P63sPmaQtKj2XHbU92udVNzdGaozKyOqUBJe2R/3VLMRYS1GNgXkli3XL
IYUm+DG++JDiwNMZ4wefr11w/xHTN3SJ2sCjcNJ+bYNcMmLFlN6EcB4eCvT5/mx6
IhQc93IO9XPxS9z8S9IwQKfQ2I7J6H8AOOL/kywg2SeyIj0BsrzxQ2X86oxp5uY/
d2l625EY8O1wXiKjrkAun1xMK0/eXNrBIbJQPCqwaG+T9EVX2X15PGh8fLSSFwwT
ID29cuyl/pn3z53FP3r55dlbRm9CgAqYoZEZA+1yKH97hWohpvHfiIz4iRkRaOIG
g3SfNOmAHQGgJGFUSPE9KL5PZ7RZhl7Afe2cKya/ZdQp3jADLiszsjNE0ZnEpAXE
GkLVk4kgW1zTlAzGtf1j6rWeyCCS48fyCMJe3esYFHbvXySmDswVG7P/r7QZ831g
kSZ91OHEU066z/vncC+pjnny2omQa48q6M+vDE5S+RtxDZzMFRWt2slqJX69AF02
kUuo0F2aYvzY6YhyIVyiGbQA5wBYUfXGjKlqrXkj/ATu/oarptwselfM/qXjMYLU
4yUYHv2LmewKKOttTCBHHYFU+rlCFNx/rN5TJ3Q3sLbsmxiXQU9evPJi3nBCrkFh
1qpLbznmBoz+81McZTO8O8XHhB7a3UdMi0fMy3Yq1+J3XOgyGqR1N8+epBQcERu8
PUnlZJTrnV3A79yjN1E+ZHTATCfFRMSscXvIQG/OMssvzmr1vhygooH1pHBnX+ke
bT/Yujnawa1QZ/uyvfQLu1BrZpwvys6xQm/tECIj7BAeM1vnbWgA3P7/S1zjkPg7
EK3ft66zdh9cnSzhQqMru9aWwZglGfY67qxncvWi0DGCUtiPOlUdjyEgfJcXLPis
IIQNApQVuSreI68Q4BwxeE7ZvlaFmljqUOM/ZxkJNYKIm2BSUlR6pA7beuGGC1BI
8hfHed0sh+h5G7ytQJp/ZG9JSQOV70N8rncXpBIEBY8e/NiXyu/WuY8+n3pWHWoi
CBQrb7UXdJ2DN6x4kXR44SV5g3SB6mEtUrHallAq5eBPt4ZdRaLoEVJnOJRqsWWQ
qjfkp61smuNxzxr9O+Xw985tBmyI+E0OhzqcfNZG3hwRWp06oakGiVrxOB0dBYvY
2rAKxI1KLeNGz+QQCD93oX00Aq/xBOeuLxGC9aJLJQGBK81hBnJ4tOlMbcNQPd+D
WHOmDLIye/MkiLoL+8TOO2kfjJxGPu2sXZGw1QgYLznyeYrcpwWVGts5OpwkuBrQ
e0V5nBXTxiPHzdYb9IBj6LwAsa3ucsPvqM4GzePlqOKh93d/vMW6K+EEGYpFsx+p
xS5smzOh9R67v5iS+HlWmWldcVjKrUXB4UTANfIBB941iOpsIYzrIjU53zbW7z21
XkEZKxUOazMLqIQfd6lvVQid60xY+ujlKowc/QZZ8zLBvo47TR56REeWizPB7y2e
yZOBHKJxmazpRYLhVBbecDhhgwhIxCPMPAvR9SOcxPXRMaWrwUu0AXKRwxHoVsBo
9eTw5PkkCAW+WzPdn/gap2yIjuR+JjbzqYdg2OrhWMGj4IorMHCRRP0eFNjNWkdA
aTwkEoB9DeMGdTf7qEpo2sdZnicVZshFF0KENUD8GfRoRKl8S4ENK+/RxZ6Ac6uq
/73PX8H8V9cnMeHKy/1rrJYmgHVEaxEKKI+LCSdoR0Pf23mb2lGw52KMy4CIeJdX
seJObIjRcgMcYOcnXIeqSU+lvMYcG8xieuxsUmsG6n90b3Wg2UIcUyZkCxJKjHA6
Eu/bGXkvcAjk56lM/+MwqUqbGhgLNprzj8pv55y4YUKVEYDYaem6CsU2NI2fFQ3s
kUT3tQ05niUh3D80uTKPyXvs8mrOk9muruHBX4eF/fY7mAuIp4AY1K0vo/sWYRFN
dNkQzh/NPL7Up/ZMUEMNiW7DhpyAavxGt+gQzHkvUb/twzaF1Cm3tdylV/1OZRu/
fCN8+jitneDthSFTtB0c7XeK8iQ/ofX+ou7Dj23yAjIuOgumsXSlTDfAv/2m5euK
hlBxzA6abLbu0ck7o/gfrFrs6bjmmXtcWB7GW7IqgKb3LZNUUJsD43s3e+0cWf2H
EdZ2jrVBks7glLuHGh/Jj//imM6BpP4Y7ihayPZFFB0SMtlpC+0Wm/CIfwwMYkDz
IQoRrWltlc1c91v7nEZbL8n1aZc5BJXUdnTzlYvhf9xdJglvC/64waEUgF/lgRaq
pOi+v1FGaHxBo3c1m6KYiWAHDjloMA+X8Hs2BsjHkfxWwkXJgApn7WvDLPLndUjR
dH9FMFJWvobuxHGD+J4NsO5WrweB8nfdoYI2s3P6PQSSkA6dq9FzkzPVSwkPQlBH
LxcwK6uZw7z0KEdsK9oAXy/0Lx8KGu7pndoxntwRJZB2XIOuvrk3XLNPTpemaFsO
KyHh+jULn/hYoMo1owE4kcvUn88q2n3uIeqK8iEZCnVaOeOOp+NYksMjQXzQ/ryO
2U+s/T5MSstXYP2icx0OFyjIndV7YMzlr1qfNafe7+TLqXqfDvXAamBDEdHBQrDE
/GpKiLgh45sZEQ8ncGI5nBotUyDlKVld03hTt/MShcCOCELMxdvyNkjHd5hSsUNx
HnnzQIH18wR+SMns+Pfu9yxMrHyvfxLp+7TvwlY3nFvZXsCETCjNKMgDWUe149P0
EdU7tYYCm7Kb384g1eda0X1T2Xf6YPgIdcT2Wr/Clx0vzSsw/tuXvMglj5y1pTCc
gVCJ9q1kVerAZXeDceXRPt1p44Jf6JOjBMwW7KxwB24kKD1cft8Yv0y2MxrGBiZA
o+nSlOrG1FaIPiJ7XerNCIk90E+E78ql93zq7Mch8vJxZ395jWjpzWrQ3Saj2yjZ
HZW5AO03bnpwYLdVY7tFdtLzOAHwz+Do+VRjK+m6BSv6fW1eR5vZOgwSOVdLY/b7
FTaWIu6yq65vSxKPMvSb2GxVRDPcVFUu2qip11hd3Eu6t2J7OpXXzXyPYRlAh8mw
V1H2jheURO+UD7kY0aacAvEFldx29eg+hHq4ipdwltiWOkQG14DL548H3da5nypK
W7XPthZYek4GIU3UIUyIGgCSotlOE9T6zdMykj15cPU2WQ9kPqB2A7m16KiZKufW
qstmUSx/Q4LcJyjAUkZbEyIwzsSBY9WGeK7S52Sj2FLEM5Qc+mHlQX6z1qJ1ovqo
TZJYC2cakAzsRmvqFhfPZkFHd64Uq8aHO6glWJmLULbjymcRBIQI0JPCTFU3b7ji
MtULQLtg+UCdLfGIFUtnLve5CwXPTThzfdT8pWzBlDTJuppt9IoQGC1QVTtn4pAk
XQ1FQZ9Tz4ysMhSJaHnJsC72CdbQhEPm0GAdk65jN3/rsr/4mzmfa5EOPBhJ8qzn
89HkhAFzAUo1YUmwey25jV8N4Zuo56cRvp9CWo5cPqEYtsE0dnauHbHqbPNY2goM
QGIiCibUZ3BJOLG4vi95urgGs8kAVBaM9EU/2IAF12znFlIF8fKo7HKel7cR5LsF
tap1TdFItlYRmzxncsvWAiYr0ul9ZIl2s6XxvnFUWBc675U6oxkB3UwU7qTGu0WF
421NvxQ9UOqlQC0+EwDG/1668gESKQsbN855K2hDMDJVKGb2ElkI7huBFlcUu0zz
QN50nlkSIxFRN3QzJ6yrTypADJnV2Tu6vZYQ8XMZO7Xe8iKRi9CNY85w5IVNCt9s
23+LmHesPvhvL64u2tkzc4EW/Q7ldlC6kxfXcPtA9ivHwSe/Qq5NT0eH7HsNSv+Z
wRfHO6F8noA+l1RFBUbZunTDYINndYg0EH/CLWw1WiHuUW8fMOmMuKbumZQ8ls5l
75OQbNpOIXWqvpRf15wELvy4ZCQ2lFWwJ/CDef31p6cRHRrY1Zg/jFdTmwc/Wfft
yhgymYyE34i+tyxrvkbHSwdGiEAYOpWYjcR0ouumB1eftx4tlsQbia3JUJa8Kggz
/d17Muc2ptApBJsfo3yv7oqHzgaw2ji+OZGPHUrHTAc5S3belWawDypmzr7ZOd5s
bVe2d3epxKV0l5RiSQGYNCIEPGfCtDRxDXPzo8I5RuSeBsxbXM+nhy/FBgNGszIr
pXe8DP01hVWYemu/KBfNPVYrep3xS2R6qVLYpxqb0+xvYMcUMZTSAAsGbdIzKtXF
CziNhk4SvSsPesZ/AW3xOIht/3XGPc2E5ihuNThw45x0bk/aAczkw/bNUOXSH4QQ
odvGChXTCyQ1B0oQnobw1jedH3PdfnNKay386eczdqONOAbwJRWZ5FX1jyDDlBic
biIuQl6y0vrlVSJUxdQDfcKxxHKwMcA9szJPFhw1uLKadTURaCzBQUXbig9RpZqy
/SO4G8gFSrKZNUc+UWZ66/O68zpoF9YGo0IKTpiluAg6YckLBhCUxDX9CPVH+ffP
DsAR0ymxQ/1bFxe3erG6EAl6vUHuBzORfcBBA7RHrZRpyPhXOZjaPMv2UfNRh7la
0SqGss6/zcBoXMAhpZLb5lGU/cfyIW6pDKXFif49xkiIlkA0IoeRa0fR8mgY7iOa
/rcnrcdxKHZ2b9zyIsxreFT4AjJsX5D+DFII8SsFuEIS3byoDAYgE2nCdxZBp81x
AYZ5b+M7+Aze3LQgeKLuI4VOl47HwwuCSj349D/k88ug5/8WWIcux5nObRtKGjYe
Mx+xAjIHf5yCFnS4BqwBWbO7qaVA7bl9e0BUp5xC63+/NftaMINI6KwkyaEjiajA
A5CcHRNX5UzY5oSAY+W6I2qvjFux90Rk8zFtT725FDGiEaG9ovgTK8z2yUtMkvO+
Rls+HdXyIKQU+oCLDhBg+Vb07LOPPeB1FDXuPtpT9zs45jexDN3fkbSyNJkoT1Z1
RnnS2lK/kcJS34rJ9CI36FFAXkliIW2Ip+yu/+LWMETZpAnGb6izqYoHikWJFnh4
24Puwnz+2qENBQ11UB7X3/CKxvW/axAID/15MEHBSHM+A0vmrcRL+GAo+YsHhDkX
DHRzlt7vutx7UbUSsEJ32BeWVqIrwlq4wJXN8GTRB2lKC9EtAhmAO6ROysKYsCGv
jAuLEHaVr81LVwSQufOsxQ5fRK7m6HOqkc9nIBppU1etExQVGk3Mf7FW3NflBbeK
mj3Hg7F7rDAI+M6Ze0IyW3RVCGIsi99m1qJwP8CeR/Rd+gdUerXRmNPajUQ56XEW
wUXIge3SczzhUk3u9yYW18aWZmTFs/0foNamcmSnwMt4ZmNFaEVUG9fec9h/sckx
7rQ243pnSLA+NBmyxv+l8m2AAHEw8jxsFZcuXwxylS8wsqEdTIVVK3d2WcBzg0MY
02ONBO9BkBmG0DxPlpMvCeKAwCRz8UZU0urWTSv3mlkDvtGTiua+p4XjozIth9FY
fXaSofyOsTSKAruEX8Sph4dutpcbZ6GV90mdSPCpLn/MThVNtTFZ84jp8+Aa8b5D
Yf/sJOwy3GFDJ6OWHR4Hb/v5+j6BXN19coXzwG5qOQsUQ3XEREwPHg37BTxya4NW
ac3vCtnL4lgedNLeOuSnGEVkbZkjFEzu3NhICuUl787jzluKBFfMxzFz0vubA/s/
VqKuHltHX601DdoSjmEgH8J3I4UTdpGjdQwLvaU0Mt88GyBfo4NVeOczJYS+taPR
Mq9nZsO+kDyl0VGKYiGCaMy+mW2GOm5eePEUW/yEBza82nc5RkdZJZQ3PtJyTwm1
lFkbaV+gWqRd7GUVw8ArPEYiEQ8wd8PPVYi7moi1r13SMrhlgCTQyL6Vf7k2qFBn
5ex1EjySSqb4zWrGWe8N9jrgen/bf7A0tBG6mKfwCaF/bDzHbI5Jv/VLkRc0Qlz/
eM120m3aPlK0uAT700d8crGqik2yZBCzVecwvZf67tTW3G9itT+g/MQVgSIWmikp
VDZ4F+mzYQcapwRXYPOuWmN8tN10uYgmavrn7lz+3qDxQLf+chSoCcgOt3ljaqJt
OY/f1O6vMBcM3gIxKvnze6q5uKSgongDoQyH1vY4/9Q7FUVHTAmrvenphZm9vhxL
VxCx2OhrifH/XUHtTn2tC8EGM9Y4fXNhp8cX54rLZjvjzpq0/NezpQklcOJZ7Yml
7qtA+yUqvncADy/cTlAEddBrOSIIkE9DFnLlnwo9wyiL94kJI4QtPYX0btioAZzT
a0NGl5qsg/OTPrizjwIabQFz63DIeXQejqGORYNaDfkRAQPneHsnzPrvGFBmN2Br
30UxC6yMUDYLo/u7fYKedGM16GnrdRfHqRFIMFGVFF5eXKnl3l2LBYyDRjQipp0A
9/HORQByuLH61wYt/1MNMx1aSlzGmzTQDV9o2xRtofFZpsG4T+CosANhbiMLDyYN
53jSL1LVRK4J7u/Qy1B6hCcsee3hWVMXrsQXmFn0RqCWwwzejECa2jURWTUgtkZg
yNqX/EfOGIr+g6UjacAOXx+nv2HFRXid7xfC7TRRFX7uxWq8TgsFQGPl6rMK9+B1
p2NDAonQzKTRrGl+0MZnviAer2eEvS25aReJ75IQJtKfGG8hP212iJBtHdNm8Hlx
nQAX2GtMvLFVF4gxuhyv7cxdXZkAKXojl18uz/6BKjATJ2zHR0x3b7bIXiDN+nMW
kw2FWsZPlcdRNiUBNDECGVRqGiWEW9prVFftklizZKNorOqtRyUpm0KjzCXvbdWV
RLB1+dboQ7mf7RomdH2T0smuimC6I2vhOruZtaSAEDXL8ftx/4q2BxSX1fzughE6
tpEGb2QGTqDUCMFuyiGoaujsmr4AS8Uyv2jcZ1zgwcpJwy6rHjqd6PfhtaojwhQU
AQhOHGr9yJLvlk24rPYAMmHtRjyTm8HF0yzVXDGJV+5dNOdRwvw78bFZt9es4UeC
sf1gm5RLnb7aVpVWVc4MSY9CTKbKEjShApG7JnY4AhhxUQIzTu+PT3HcVXzVTLQj
0Xc+9UNtPZOjQftN6m1uwvVyQ+YOn4mAU6kd5xsPHFvwQ2bleeCyXRasqllWLG7F
CYE0axmiDl3laHMRsYUk8pea0tfuE/2FJXHNbuK3mzeWRcRQu7z5n3fFcSLh+5hA
zwpRlx9Uj5krwn1swIwNt8aCexJGBhvUWgFx1LU7CaJnIPO2jmIyyHa34qtTE8xc
aFYVc6wslvcqrC1D9hHdVoDfe4oZzu8CNLx8PBN8hckAMAAJ1aX0QSYQlDG/IoJC
KTe4/FAgteOr2y6i27bzh4u8eHN3qqBu6gATmwjGnoHricmedjOJfFUxVhvnCq/z
NKWcJRfXVGtHe6vyIPdbIyr4nb9ZMOUig78ICFIMuNdFCoS2X9C8wmWwjlFUmcDX
Lw0vT2VuNJ0z1hQPcXlPFSa96qoU+hxYEhkJOfMy1eRV9e8axhUhTmmKR4fNdXOI
mXLpbAN4jTOlvhRQt8zbgwXOEfmUEaJC0vgyc2Affi0LNKrm23XNHaOFoUodZTQH
AFgSOQgTq9Y8XR3ltRvTAZOe1hckf7sbmTuzp1wQlt19X6PyrmJkdMPxGqN3cE52
q5q5u4fpGGSFcZcHeJrdMZXwtMky5ny9o+bIT9cf9wVQiMM1FA8UWP7UP2vimSyI
BhkqTFE2WmAp1V+bGc0y7laeVF1QZ/21gLW1zd9fKW9N6SQeTG4PB5m1fm8yuKKq
WSylAhpzhqH+rp7VK3v8/IfDqc/tcKpJ0GQBr2s6LRBPAPLn2aqmJliRGsg29xnr
IOg/4igAI/aDgJV98SqFaA/k2z8lL8LIl7cgvGZqWLDszldyqOxz4nf7pFsv9d15
EBlj+I2B1FkMlwjXP+HaP0MCVGSJefwOam6zJ/UOqjDF2tBGF84+NygVKoconsXn
sEqE6jVV29sLK66fTJ/UCcs+yaEqWdhQ7vfD16XiRxUxiJR8MwotTP36OZAGcDhN
5UQ0leEl033YZOTFI4tDW8kfPDYDtzfc/kXLW8r0HTXhG3jwxnIpmgziRGT4nvDO
c5RghgYFtiXe+1wIY5dbq9+ttZPD8Xe26KZFtBXDHlaN2kJvwL/LMgu2/sXdpN+a
UiDP9BKoX8a05tLBENcWYcKM+W4P66UzNSMRAmOt+A9rBgOIxCKoXsnzzggJKhKE
HYsU66QGNe/jDLXBy+jgSlVQpBFdb/vRO+qzgl+WMQ+x3vhrw6FXepHjtJJ/FrGv
fVQl2QP98MslE1JToEsgFywLuMd8iNkLz8XA35EJ23R2HJbTr6AxCgD4bbez7K07
jEtH1HQy0m1cGW5960IkgWJIZRPSqFBp7VEfHPZEYoqWnQ+sLQ6w5yz9URxlao+g
y41ShSX4a7ht68rom1UOmSF4V2dCySaADQhnL1/epRfx7NI8MDrulZmxbTJF5DEP
HgNOD7ki3DIcPbPFai9V+x3b3B81a6v2sfrpe/6N8UlvM0pr26zVlDir1Fn5qHnl
/pKOlRf1sqGUk4j7MLaEw+S9LpTVcFQaQBJmKXV+DczOxmOYQf67XvyUOfcw6De5
x55KETlFAUcxQutkhlPO3cLEwxhYhGFj6a1mbmZYBkeKOTdYF+icsgZbAdJr2L9d
6jamzRiG9Yoa2Uw7nfIUIMUbXG8z3WK6LJlVZjbXGBOdJoHdNYVEWZthBuFSHwHz
YLeO0EXYCuyIk0IxXAlB9UZZ9o7qb2NpMN1V+h+oztqaAZ/B3842BY9A9ADRm861
MIR9dWkQnRj1CoY8lmMoa3UMn0R09N6MeKCEA6PneWrgSFkjzOhRj6/fwB1t/4ib
Gw35f59+zimClveeLbL5M43GOSEuX6pJHhSMpR3TAGOZ8A8Uae+UGiZHyp2hZfQN
h/6wqjcGdPxhOttLU4wcufEuyq1LMRnN63Wqt5BOPlErJ6CzCoe3A06eGw1cU5Z1
/uQrCHdIt5Oub3v1LWLcqQtX02xkKaF8qWM7Me35rm5xVPtfijErIZMMO0kwelkD
XqQJhwbkZHRaDPMdqOGJUCV7UCMSlOyFAYE7xftvLrix7XYVZeJWBHD2SOOOOXkx
ETVNh5F0Cmseg85N74cdKmwqPWDuxR/r5S6UxAcMMsGnCJdE1kUckD1WWq14B+Rv
BE1Qnqv/TAWkUsi5DfjVz3UXrHXgnXwHgJNq28HVTZCxyr0pP8N+ahSc8qfh1Ihn
sUBSELRmGxIqQWRW/zsKWnjm0Sm3MlqE9alkq4VUIa1uEeLV/mgVnhC49WmarDM2
imQ0MHR6hWsLyreXhbPBYQ7YzTpXl+G7YnghHcreQ2a/rPR9OoyugY8e3uVPqAvd
pMUPdRjxwKD/sYB0l/gPPRQrRehqtC3/oU7/TbFjtq43HjhtHj3eYat4tlatTgmC
n2pUU5/gaJjitrtxgcLbf0CIqUApZjogzBoMzq1UbNtrXyn/bT0n588Vlcyunx40
uZfyocY0S/Xj2nOSJmIvHJqh/uAu3Bapu6ElWsHdOIQ4myOqaW8JduQepxHE/acI
d02Uk8CMr7i5Clza01XWTL8MAGJQIBtUdwy8YNpDIQLy2g/ehz++baRl+s9dqohH
JlOCaAAB1mGSW27YMzWfWxx4hRU7IEB01hciY11gYoXaVji9VXuyxoLgtDdWMMHd
DzI8MYZyLhh+IUhvsUAHWa6T3alP3wUozOXN52/DDDqCF2ZxWTgEaS5wxU7bkdSk
zX6IzZo5wTKZ0O55EGT58F1ISa5+fuPTtC7Ivi2Zvth9xO+QI30wTfnHNENUMcvS
bz/h3LX0Wn8+9T85yMG4ngtNTEFNQb3WloUsJkRIHBggzL8Wd8D0cYHtyZunXx8I
fS8k46tBa3oeZhrDHkfrir4XfiNMrf1wo3ICxHSis0FoP9FxG/5MMO2yH4jGSkrM
5995MfDmFK+w7316PYGA8/faJ+TzkK2NfDWhdVsYBhb3jBL5a9eI/vbhA5Rhv4WS
ytDI7Q8NVyt0Lp5MWnbThk0SC3//KCgshpjIKNLpH1Nz4Zh9Taowcacb0g1NkKVJ
c7mFipXplFEPLdxHXjhlQMA8Qw9pviclkKir6HdaR/2sYh4dBpgnuK5QJt3ObVpl
i305nf7ZGgM3FseqWb/VbMtR0tyfqwBQ5a+xtXtEpRy4eyKym+gDjZF8DeHCN6Hk
uqjANOq6XdfH8wVStIqXo/bQ5Tm+KItfXeiWm6GQX1HOUOS631+Dvc7mEBNhNG3S
BNQgyqhV7R/bkucnoPYiZeWbeQ7A0CgeNaOQqYRFuEynRv4eScSyGi9aHFjdNgRE
D8gaAxTu/9iQm64b0B1GBJSIkJLRQLqa62h7oMAGReE6lgSxtJJt+7/pqqybPQo5
OXsCQU0HpDkGimot7tiVFPc25kSVaxLkTs36NMU34sKQhOTaxtGA+VmI0PtWCEL6
enbaxFY0cD7WsN2BzBMbd1Y7Ad/vVJdd86QU4Tfw2NSfrozoK4yWmAadtvntG13i
gkS9Bj20gemCg6uhVf2+v7mcr9Dn5UpC1Fhynfg4nHHNs/NmbB3EIaUyHAR0Md6T
hrjGfzKut3N/o1IYSaA6DBXz1JE1om6EQVtpOkz5tpMUCsJCMivYRR49hM/iwWrp
gCmMirv+HqN/SPlOXpRHgrYXvKONeUbcx21xZ764vMMDALVywH/xiu2LTWFyDuFi
e7y1IEnYVr9cAPI+SSeRQ1C7ceEYLqNIjMIj3BlbiqnD1pJ0qDzahkOadwP6ke1v
Lb71eLTK+IeY6t8nu2+ZndkvAOALT+Xi0861NhUmu3t74gaDNXOZO4RbJA+Gjtw0
Dqa1XJoLFY9PN6GK8viTAcVrqtoPsRpnrXqpmtaCLSGuQYIWHsDv90phmcTn+KI7
DlhEw60dU6qzWMIRKzk1P8pksGCdRX1Y7tAlU9cqX9nJhlXcZ6EnaUSdASAFRh1V
zqMFdfWpoQtI7Qzx4sck46mAk1lgBRe4kPysJ8oqp5xAqye9bfkgDcQun7KWzRBQ
UDB3KchN+7sw+pjGR8QyLXKKG1EQ1kg+DT2YxjXHI50xBu4h0QWBzFYUJZtEUHXW
q8JyHWrKlOi5qIfyvSWbAvYsS3xQMkrFVzzWKpa/2/w+2BO5C6z7p0Km5egyRjCQ
FWzIsSMbHcIz3l5L3zW3hFmM8UWOIAd18oE4QRswoCo/cFsU0SYcjQ/V3LqpE+sv
2V5K0QXDD3QJVwkm/Rm1o7ik87srjH3+6rqJIaHZ+aMvhBwl/jT+bzhGsAEhSP5U
CCwb+YlZV6J4YJpWrtw7wmgfiOJVtzkMC+Ee1a7qTN+vud6r0sgIj45RqOivN6Ih
FbJt0DZtGWjxnW6i8pZbsf1OvX2gNyuNCysZF9igKHvNl1bROiWo+9/iAJfu2qqK
gtEoeZQlNvVK5iLk6gYrdMdQCwTo0vD5urrqr2oTnB3FItaAZfSBenAUwkPYWITG
12eF0Caf3FCT26vireZ/T9eVBlZE/drH5SQxnEVymiEUFj33Y+h7oaV8O2rbADza
x6rX2RUEyeEXJJqSJMqhsCNzzHfgClbSKodKqYP+g4PjDo9jS497gnCt6f/M71qx
Pi157oWbravTObo4QuORkn9hG6yDw2ztb66nDVzBVQhF+bMTKmeY6BdNZrQ6i0sm
kJ8is14MC3FO5hYe39mVpHWhGVcP57jKzGOlef7//xJYOwdnF/xoKQFe4ptHGh8G
rKgXWMaQIxAk8VKcrAA3h+2/qjFtCSlpBJX4bOaohcQufcwa6HT8T1kt26tdfXkJ
tf3LjvVHKJ4OYd20kx8e2JVwi081qQAjOkPqRT3ZfdfGdNId7Ml0iT11HUrCxzDv
1apvTqNYHHfdUYWGKV9R3j5B19sMXtMHdT+YCLa+jBcajLSLOaMtpbOmKGNyXhSU
Wa9/cW71b95V+BbbvP+x5645H1ADXVC/4gAdE43G9QsPI/qCLLCikVciHx5k5IH0
gx1B6EyHyQiIdde/GWn5HoVChQxya5DDKnBZbPt8p7xLVvIvoBJDzdtLO77r+UAp
QDM7Cto1EySxT0Hrlb2XXgP+Kot6sNRBYkBPNqA0QRobjHhJZ73V91OVaYjIjeTJ
11Hi6JEJ04sXuNj5ez2rr2JAZYg+N730WSJcxeOdzimrGXSqVWWPxLweMbzXvzCA
/h841SVfQTukr/3thn/6ZIskxxRk9ziY/r24F+lKz6IcOm/dupxLx8Equawf4T4Z
MyMY2EqMKe2SAp3NotgmHUt3YfDE77OyhyAlUDhRfWM8JYSPeKTi0FgrqhCKPtmi
VXUHG6lM+fww6agLL+/qEqJRW2FG08e8mcrHCslnBVC6W63LjnT1+TUwvp4MI1p1
xPmmaj5p0XvsQCPl7ww6eQR8m85ph8L7oDG/6ZM7sLJcMPdmCcSnF2WRIevUf0e3
ni6OGPfJLHgrc41+tRCc7SArcGueXnQt4Y48vLSsBkFrQQw3QyVKeABKzSaXsh7Y
l9UR3n77P0heWNVfUVhl2H10OJRs0RQPnxJU1cd1GzBcWfR75ucZ3/pc9fzBFzj5
29ub6O8O5KjbIo7LbyfcWdVbiHhjRWUTiwMtmlHftJoMNOTT03SDUwarroaInb0/
zNDJvlo9otBxv7u5OQG1vbqIFOAfThIwhDxTNUontKj2Xab0CuwpgJWZQHZs2njg
YRyOoaFsnBrBfUGAqFREi9vLOGLg4FhhGjk2mOt+k2FDnduEKIZumB+9DnoReiN7
h2LdS7Ti4Xzexc3vwVCXiDnfvL5f0XB/n+y43oVgEGqfGr3rxj922nJsc+KO1Few
bv43d3rHh7C67hbXnq5BCY1UcGB/tHRIUP3xgd3wDwULcHKBLB2zF+PDok1bmzPc
lFuN4ROCoSbsxJJqZHeEdE1UStfKfoq8ol+5X4kbARKVuFBVEZzvebsyo+uRT3DI
YiXZEfwqR6w0MStDIiOXI9yH6izQt4iLbqrTkSB4dtPW13As2KqdFcyu6FwyK/1U
D8JcT9i5sf7ISjxqxOgyLbyGWliInDxlMlMh9O2sue+az9YBYJBoN0nwir3ItBhz
p0vPHTNNEykbpNkdsmaAv38rgAXf2WC1fkn7tvxaoSNHZ0UO3TzwzRfC8redmhMC
O7D/XIHJRjUJIWu/Mai3Ka9QI1NWbUoggQwyxFrXkiGZkJMJT5Idm7/rDmbH6cuG
BIM44hgklt1gMWkGyxjrqQdODSjRncuRWJA8VAeHeY1pwSw1iJUV0CCS8yhuwDNy
1ORo0piawC4ZRLvcnErsVDTcRM+nT/v54YUKcCPGrYvTBIkWk9ji3w8qg5/TFNdO
RRDa9yXk57mhFfO76RqpesJgFo0c2MUj9LSBIuzEwSNWxc/6LNq9QFX8Sj4e0yNM
33ZqNSq7JjwhVCGe8OXiqoRJ/yR+vCmBK/Z+bATUQrx9CysOzQjoGZUfVU+dtgDy
jKaKT8tDdATkyv+WAOHehgoCAg/WRLxGaMxB7U3y3q9EFsNxblOcIW2/xpu+eJY1
OhMopHFW7RjiE6f4OAZ+60khkYqBKWC5mqkOACfE3lBM/EI6zUKfOR9X7UmNgR/E
+GRWUwfczfjM+mbDXq0gNwT7QG2XoTOaaXKlMd76Ff4IdqH3zibpWwtHEI0sRI3R
8xdPdFsBFz8WS80xYvtoLNTzMW44tLJETiRn0m9NTG5cfQHPYi3YkwGnWC99DHdA
pBaOWRFpTow8SChX6v5KzThJvWjgoWSOv/yaSOy8TWcG5BdgUk1vOm88t+3BMwfK
Z6GqJdu8aOpuFT39NMi5IYDK4dn3cRsH045qkxgapTb0co1DLFaOpZBdhbqgWhB7
klmdgljvoFCorl0B9za3vANiWqqO0jL90NbzV7dRTb6tjs7pAHrb0ctBHqxeXVbJ
q2NYXEK9t5wvN4PypX5eeM0QgtuFJnT0udwet/vjtoqNbx2bgfwFVVEXW0yNvPyf
x27P0NUQ3R4RWw9//GVU+teq583y05WMPLMc/PscmyWS6i+yBQj0spQHKBfEmvC8
Fgn/VDc1qfYUwl3nKcdrj/tOWm7M6ogz+4jrQ4JPLmFMUWQzybXoKXsnPg2a7H1H
AUF0EBU8LJqDaqGwuBdprtJRLLNehrjzc+J+es5wzgizwJ5pxq1sCXiI3JbPCo+/
ERJqj4qGjiNZR0eS3+AnlRUIqUjiScZV2jKGmnGtyjeDDUnNGEY1uY33L1j1ikOa
PJlvhWPKpDjZMAM1y3KcuBGACtc7VoyzkENerZ4rdIEPEuolJnJ7LgDJqh7wJqeW
d21SHZfE8oOQwEv6Dh1XQK0MDmIB3+WpKqKFVduEeHy7VfHqbp4rxXhZcI1HzLro
gs2cFVYFRBlqRBjNm5pCWV6q6H5xBdo5VCX3y9H+/8KoDvr3znvXq3QkDF5bZPIG
yZlNJnnsx6gnOAXBne0j9FBR9SlmXvdKDJhqQLauGr7YjzzXFj9gcj0qP9Myb9ml
ZsGcq0V1SoCNs5oYYM0BGdAPfL73c/PRDsxStkQLFRbvTyufK56EHB/PZ7xlPtdw
8zrMLvcxI3yKdAc5Z6IlJiIEquxoDRfJqZtNZe7gvNsE0dkh4QvEiWRIYORLffcb
3L68jiIJn7qgSYM7QAbcxD2JlfPsAzszwbtAIi7ITd8laGaV6SOdQEsR9RjWzbhL
4e4DXmz4fGybItvvYZleL1BjDXKSlGX9IRs6r0ux886nsE3B7gn5jnRe29wWdD2V
C+rO605Z0NudRtk6V61CgtvggZSF/VvRRUgsojpUNOp7aTd3NmHgyPw27p7oTcWl
HRdZys1LFCT1x3dw6QR/v3RmGsXH+0k2ZyRRWsJC1WAzWv7/ShuQueZ1EtIr9Pbk
MJQ9Wt0a3yyVuswH/sTVmt7o5bTyN0SXjTU/T4oYvuf7osCuN6BCc6oLw2QJWpJ+
hZ+4tEUbkiQPdU10y5hr0RCBdUdTV7Wc6vaa6AmtdnsAd6JlY5sBD9Ki/lGRIc5R
g3WKvzESeFLCPFZjtHdmN+72U0TuGVUi2kwGQr1kyU0wzANqSTiCqfaLp109n1QH
gjZidhMXOXGo1XzZUzwPr54dS75PE5JQJuDWkoxlxT2Boud5kiHiWDWXWN+17yWK
u5bp13uhuEmTWoHwxtMzQsMlBHfZMeSxcA4D9/QTyKVS5UZDEqqNjn2UXfiWlYhn
F6cAKAbR/v6HNfXPxIrxcZcBYbkWVNcxCLFM5Rxm1C8xQBx9G76iMkhQZAroKspv
qbxtUjOb9MFFgNjDc8yMR+VYezJBWO2vmViMjmjsafLt+KdLp6MKon1fpYq6qOE4
MLpp+30+KfCYYiJ25qAPsMJbmVXfhvmKwOZSAx8xJvxypQXhlUoMOofQw3O83fBu
Hwuu/930dl8UzCYXk2lOwXyb4RpzXRg4d7MF+sr5K8l9FzDZDg0qlX5SXqXcYqmx
v4G02HPczrphhIkq6frQZX97RbPpAPosQ8cfs1cH/9qxxzn7wS/xdmaVo+dcSE1P
7LUsyfY18DO15VbWOPkWX59TR5G4hfjYS6zsx/dKNWwlC3jkt/+yKWT+Uf2yze/I
+dmP3ThTHxUUWSFK0xKDyqTw2SWA4uhPEuC6upb3hKgeXFa54Lukxq3DtBMX+D53
ci2TA320XSMgsZl0FGRaUY4FQYpSJvgK1QTydrdg8yuAJh/GuKl0w+c5uC45mblk
c4eyaUIdwLDb8c8ekYRqQeDYgVM+Ds3rDKGLKBZOH+6BOC1ZO5yPoXAMbP2etHU5
yHjTraY4KlbbuLBynXgVSN58uXB/b9EM1cUrBpkMZKgM01ttuiUvKabPt2/fqtYj
o+7Il6ASO/dWHi0+DuICmd22pDiAbOt/E9KFbV2eFNljMVQHg91JghN73btpdLIe
xKp23EEMTGjpkrtPwLGRGqPci+dV2U4lp1ctMNSr8Q5dsWd+oPs6kffQK4LzdVTe
mb1DyHiHkl3b0l/fW5UL5+Z7HLkHdNKTHErSLqL5t6q2GP9VBo0oNQ/TBBVrv53N
H7ltTjbZpJ9IYJecqhRc5B8ICo6ZeE5D0UE91sYFo5PyQAQUK2kcvgAUUYuHwiYl
T5V7AoVSeZezxncM6NqYcCJjHT/ZNTSBBipQ3iCK2xQQ83RhoWbbu3KDs5vTk0o4
yaynpbYQNoGeoh59uralGG6vG0rOljhUeSf+LvpVFEdoDfR5WtMBA6MduxLo0xeY
X4mF/KEAYHN60Kat9lBbCBGKwp+WSFoblhD/ewVEQkIazXCqCHXlcyOGdySu4Fna
UBdyMoQ/vQmaqaC4Qd8e725OG0sQgo6yuca0E2nduGqP5UEXM+xq9chVgg5BSLtU
FgQ4EJivUFENiK/W+97LQEQbN3b1KnXbBT5q2AQ2Tcaph+binGgmge9/qwzLrwjr
Shm93awHBIOk/99oWo0Na6j16D//GUWoaR7fxWrLR9P3nEI/378noAnrx5w/BFq4
dkQrE/uHyg2yCOo0WZzxF8+pLzUFccAWjIjvNUspPgYq6b43JPqBLMtSDMlGV2X4
yDhL41Bh46cJY2OiYUwl99yGZ0S3BspZ4dOMh0bzrfUtjVF3sHXWhLrtk09U5cmf
7Mu66NF83kjP1NWeOE5TBNpf0oozZA2p43AiqCPabyaJas51Rq5zinRuGWGkCuSC
+74mS4pKRGqoPJdjMBkGYvvft8aXzV73yJcGLmnUCWGxCEILu1cpzzIkZWACQOY1
yZ9fL+AovhLtDFV5iNWTjc0YLCTppPWvxGbM0kBcxFidX4Ftvw1mSKMGhwNsPk60
Zf1p+YQSycCsNU3DbfxQ3LJUjiSmg3PYchoPDur3PKzezI6B948VAMvfsiUMkimj
vtvYNZ3iLoCNubAa+ytwalFG/ggjrZFhxCdkzrIeT3WoxxVXa6XBjGqHpR1heXwG
yE5dF/VxAjbygX4no3UI43lzONbi/Kxvt7p+plK5YfLBekU2TIlkj7uC44xwDIrz
RSEcoDFkluKY9FBMmsg6AP2gO88l8TZeF/HwEVb2wIeks7bO/UK9fIyW2gXaFytY
jbtBpRxI8QC+4o+Iv8BSMtWtRV5t6p/04tr5BJJP432UttyXbIdPWfLgu/8cFCxu
ippJNnzO9P8mB0d9nHYxUsiU1nXUKjVDxjCqUQxetQWoUFzwpzhE8tYE1S3WUIz5
V3ZV1Tvv8zukY55LEL8yq1FVokwadGN3bpjanPx0Fg/z4C7ei5yocxh9Q5i4Zz8+
0quxpeJfGizF2EGr/gZGUHXQAOw2Cy8xaNs1dht+k8AQ3/x1wEBWpKoydjAHBD8M
CMgyXBbK8fmI7syFS168POeNTqUAGXlmBKtZctZZ6kIeCiV0CVGxek3jXildRJhU
Ry8ePqrBn7wsZhFO9R6+Exu0vsx9C7+23rwUQPz3EYBb/mQJ5TsOcaY8SPUwCGQI
G0MVAn8uTyn7PKytxwhO7jMQWizvJy94suOukzi0nfm1y4lqleSRoPxYxIJJwoH+
cTiC0T7bT3rfUbKfaRDQQSC+PaDCuZd+cyC4T6lSLW3cuHW4ebAirNf+p+YhRV0z
9cKEkXLyvZzbcB20XY+grDymaEpMzP/QrIoFUI/ZwkUD2cHfeOM90K1xrr6xJMbv
DvI3cM3V3NIJtF/hxO0v4EOQQlAz/2xt0hNsbfCKdwHFEgxVLvmmnCOb1fQ2/ZOv
xubbBmfiTt4tdXMhDqLOj4XnFOu/P4OTh0M3sZE3u2KNA/DoHctO9h5uWfIUAqei
CsnjiJHxBWBdaloI4Se3uYo+etwEHnnK+uXy81sP+coZ0BlT1hldj+BN2uLZDiab
AU7iPnckRwhKsdfJ70pVR5F0npo8lI8H2AEpdpHYWMibuQ67hVvoGmcw6t30SXlD
SgpQ8enC1cRTpSQBbP+NXW67T4xHZPpRG/pf6w3ilgVRJR8U9+1JYgcBTZn/5F+k
0sprucM2o0mf6G/BpaMODli8DVMvKfTvrlG5q2H8vZJclW1CcGKlSsSzEo6UULe+
OaXDm6p/5mI8UlKjb0+QSkwTy4VtGOKdxUuuEZaoLROmWhw7kgvxa2F2PoYKXmkk
4Uey3A1d/81n0cLrE4f+9sOkYiP4avjcD3hORRwFPpQNJTLVSvfjdTLrMXBy5c74
bALhqSdups6X/rfHvaqUS4Ri+Nvh5SBupeIX2bifZ/Me03/Zda72ZOhsTQHXvufg
ZDFHIAaz/R14XOBnitogDn1OcBVLWytOLoEyD8JhCq6z2L/JxhxbU0cEIahoOGw2
TLpiH8aS+EDIHW2cKbQaY1Xfq3MTpMZLDQ8s4Dke+LeM+l6+VHuQ4dPehcwdGjd9
yvPtJ5dGi1+2piXpDCNo7fSPMXsS+aFuC2rHou2RgSzSDJSkc1kFRBJ4IsHju9Pd
RbOTGoc7PRnH8p15SELFEirMTS/lADkIaXRn8s1R6bNa9KWxmO3r1W9GJpqOdC5u
ViJsEd4S4azNyqFLyvTRMlQ5jyYxJKyiC5XR3T4HhOrMTmtBdMunkMsApp2Gsw7P
PxTbPustlDtYdipZNInhxvzyXFn5aC9eYftrvAt9RADzw0cSJUvvUiqQIEDr6Tvv
hQHKW03ITPhUBmR9nmTuAv3FNGGwnTMRyQXTBMSXLJMT/4IHIPH21l/Krm5x/aMv
J8iK7IV8uBqGPHlICHxoPl9G46SP4Iyoc9/VwSSyc0CDnfvwyJXjnfByaN9LHrq4
6IfPtGbA0o2FcQkgCnhhka1ZVafylJQDraYLBhR9o1KE8EohNg04iE7MquzfMJKW
QoIshdqgTClygF4gzDeUcVPn+AI2zl2waRCRFuo+St71aDix1yhO49NloQ9wBHKZ
bWz8FMEck9YpTGnBuC2t+T7fRL/qBL9e7f7o92FrTzIeExqHqYcl6gDnC0+VlMtb
Z+rfdyd++RuCii1o0uITa7VEpnKAcQwMdwdOqjCdkRrVA8vdvQD2D0zGZrYs1QLm
MHAI8YWn+phVVKIts8OingWGHF2r4bAkcqtPD9OtV6xpwdcR5BVYbHn7K3zw3uO8
yUrKtG6n32DHNWy69Vj+vy6smNfgE+A8fWA93VmNNWVGYLCop2slNVdwQsgoxHm1
gTBefJ2aYXP3g+VUefnXHlnOnpzMbMCELUYLK3ygo+HK0TDA9bxFXls+dP+SNHDq
/AQ+q+L/yHQzES52o6il85snzPPcSfLXZQQUyPix11CSFKxBCnYc3w1B0b6U63AD
rcUhPTIZkhqjo66qzC1GHM59UZNa87AIyCLyqZ6P8CNrjOU8p4U/vZ3kd1hrNLpr
MBUcxul7uMH7cq+mj459/qvSnB/nDAtEF3VJJ6nc2rxG0+V9iK8DfGEjAf26nj1J
Cl6rvF+mJTtF9cvTq77cfC9or6YYmGDSug6gOTW+xgVOPhHPQEfRj9pmJj1eZf6w
HRAWtXLXK2vNiw5YxF7l+QT1a104SUsJw2ZItP+4550lgjEjeLUtWAOWkThNyPo9
P6vitOa2ikeBFE68kJDkM/6eyF8wfgUl/TBtmjG6qAIDJ2HGI70LxWkaz73x+orN
ppQSGiysmMySDJTmj2bRawcHhYidH2B+aKD6N+UKdQ0tgkVtDlVxkWZElqE1iw3U
vV9y42tFMNABzfCMewhJz6UjDQeNVNIW5Trxf3276uLVsDa6K22hMrQqri9vIkkj
5etqqrbcK6L4yVxhnNlbts3j8iCoqWd7C+aIxjzsPHvaYtN1haPiuPBFVLDVvzVS
5megHnQPaD1bSO0wiuC+9tWipD4EuoNBBHaLEt7MNyEQS+XHJyYZPRBDMue9Kdcd
2fgaseBMHuoWitrJ+nyoMMejirmEufnGFIWVn+qWboY1TpB3Odtci6priSCAfPPV
O4kiXEw3FPdFdXGRxYB6g0/KaEydpzqH6SBBpovFNdn6rxX1zItD/5lt+xapSjOl
RA/xC5j4ZagE0eQcQV2FUpTakYW2GZFDbYcw2AAuNAa9oicnUXTyOHqZOpI9wPhQ
8HFnXj6hZgU3xcNmVXnzdSbnqsQZm1o6TgeyGh5eHuwbCXnKrCZAvR/eh5imiwwD
1zLtC64e5xJKMh/+tbr9xj7IZqGYW7Yz5OxaCrKZybvwkMQ8amtUfvfwHjxAre+I
HYxaXUxhrvA3x0CMKhG5ryIZLYgMrODBd+N0nEKd84rzTmtFIG78HLl05m95tcEP
cHfOclditC7RbFP2dK8FFLQvsyCrJewvXhgQ4lrRUSd0PD4qpVLugimoLdEXIQLZ
3z8tNV8basAIuEYr1f4AIM2jcfS0DIJlPOzAeBgfF6L/3/rTVNCyCkXqUDcLXKb7
Bk34/y3j0wwO0s9nETtAnwoZAiWic9ir1CDAEG31N45k5THf3fxjPCKaPXk47GkH
em2Y/L9AqYz8yhfm/q2aZKqt1jDOl9MpnkW6jpqTvXTHHRNkc7PX/6t+jYVqQnCV
0YwBBdcp0jBhIDIdJ20baUJv7xS9x9JUyK6KD0fRbyjt4e4F1xD7nOgAQFB+LDAV
SGwwJaOxuC+f441NgRZ3Tyo2rG9gMhjcw5OXsb5bi5i6vGqq+IB0SH5bJKlG0Dgd
wZjV4Fz9RusoWqnPuDPkrkVEfIUwtRpFSL2Qkgs2TljCsFz1RV6Zl7gWRI7F1Pcf
psuLkWuxHg9s6a5b+AYHiT4MuVxIayKSvATa0CxA1rNUVF+5ggcJagx6L1/ukQLk
tg0EBMc8kjhVMmTYwUJURMS4Mqv/6jq8DyvOJ3+IHMJ49fguO5RfG1Jtz7VE9ISS
lOXmA1+6B/lo11+ptAim43aixXt1Ieu4VsC/lSjaM6Ejov5W+8/KLEpmyVqUvoFi
rAN/NiGVBl/zvKRNsiO43P3FcyvlvZ+CeuFh+zOM2TEUOHTy/1XTESB3VRO+8psL
9Emq5uC1Vbn4gN/TCDdgdHlbAJSv0EnGB0q6EhHnmMn2Pl7AuXvMgFhPYQ9YSk60
L9BMk3ZIZsV8A/5zmUitkH1hO+HrS6RZ/9c2za+wyXqaoLxXIYMUKyER8ytjS/yv
ohMIS8bO57ssO2oWxTkQxF97i1CRrZCC+guljRbbJFCc7oCxkDDMz7WPYW1w37T+
h0WsHIFZmUGWHxMhVYV9mmq0hmJKS/lecjzipADGBZWyA3HbJOLNLICnbHat16GI
326RAscqQnVwAUSObCSH09uqJ8+5kHdzqZZpIxarWrGb23ZIfEUFknykVFu3e18O
KauNZHT3LtBYO+f+pZyrCPLeUvfUjd0zYxt8Hqftme6OARiGkNUtxmXgIVWpKiaw
7CDYwL0chF90QXLLQGHDuZisG3b1xanPwiwTZZWIBFbk1fTfFm1aoCCbQN420Xx6
Yk92QV+BKd17U46eSa5LiI6MJkG2+3r9IqPYyhwxAtfREpznc0ZzZP2bPSbzRlcm
2mTaXke2YCVmxmoq2ks7MOh3L8Iu5X+NWr9+He0PoiLas6L52k2ssJmXzLxZ2xKk
Hk9gqyhvUNnFr7Tw6GgnjUDx/8MJz22Y+SAWDK2IBsQuHa/cidXeistuDkGV3gVz
x0ptHT7sz1C2h51uv2lqpEo7mBvnPEbjhbpr7wiyLDwto/waPFVL8M4t+IYIFGqD
noqXaZGQLF32MB948728oZq2uQzUeT/kLCu+jzzps0hW3Bv3mH70UJamlqZYI7/f
fawSSrRKNdrw43QdrI9waKNJDxNB1VRQ4dkvj18IcDRP5BD/mtmFvvelV3RnfHDI
/eeMM1dNlgYB3XSeMk5ZBI3QNlwVh/wXWvcWm1B8k9oXtz/sTscWjMQjeD98DW8p
iUgXnQI4ATp/Nr+0mRAIJtfl8kqidyBryI3j991uFD/NYrLZ5OerUOPKJA9fA8fa
LfOxfNv2cz+ZQ5mS8U+eJ5RrXg3Wenc5TAAV7RayZA7kHCh6qQAgzRy0LOV6m/fd
IolrIlMe8di/3iEugyepNfe6YDraevQgKkwckIQbeQ0Gfx8RBdVnydpQX15+5YBR
iVWxNjOi7w/GX7xghWBilJVIH4TzFb3PKFURqKBX7p3YBw/jim0QWK3Jw9zYY3QX
qtfNZXWWpOg6BPliTLtnYHF5vciXgqFMJV4QQuUol+rYDcAnDHEqkawU6tIZnN+Y
UrGSx9ngNrTTJ7cRNQmq62nSTPPreNNp7eeg43zwRds/Uxd1h6IH48z0rYjNIQyk
UZPvpq8YjX/hj95YQoYbhyouQngNRtlRcg5Z8OrtjO2EFAntnyoNy1pwO/yu1u9j
ZrJZdXY6ZcRJC/gG5SwIeLo3i+o3qhtcW8cCMlRt9iPTt26dK8/u1woAwg2501PO
gZukYtDBDgeGhRE9gxHtyEHZKoiZ2Los2YMQXj375ERGfKaMlzYvEHKWJDrgw6Wy
XV9m1ehXaojx7KhoAHyk+1sJziwmo+m17cmW2nwTlgIvgjXQBOYvbmytgw7Ws8MG
toaNV+7n7e7LyogSnv0o0BpteabnPPUcwKwfdpG4Iw68VrKW3p+VUQ+MqovxLw/W
3WXzkMRlm5f8M0E36IvIv9EBDozFnp3xguGn7JMwyK8tiep+CC6NQuqkj9a+4Mee
lRFA6Ypbfw2EpiHkvzUrNYqy3DCIKraB4qOlBRcaWbbaqStv57bypoTJPmz00aSa
Owisc0kweJ7jQmOvd0wpi/6mf3Hj8gYztTLizap/jbLfTF5pNFZ8/WLB712jHYoX
Ag2UQmfOqwRL/OlTj26fn14U1nhnc2Kzy+KCTPX9BmQN44IJfh+sP8ji654UEdh4
mhl/eWAa3V+4eXX4j/FcXaxUKQin9PlPM+SJtCAIUoy4iN2ozNvTJFOYnyfGlPdp
3IFPJ/c1F17ebwdSiQM3QgskCrQusZvT//SaY0c7ujS8jKbVIl8EMu4WovDAvX/E
kJIcNP0SctEzwMQ7L5I2Z4TOl63awI+HPNnjgZ0+zTqYjP+7on5jKp4zGa1gWUYr
1h3O+pu4ge+uH+bzj4rQ8b0y3Du2qhzGSHYL9guVagtDFvaCG1KskTn2LLFrL+5A
mMuG8cL5hRfJMo5r/mbvYcfn3oHxAk/D7oYS8TsqhdwXcWKvBvwucOZ9m3NsSFhN
BbNPizRwew93uFGAdEm/Zw3E0dqbYySISXp+Th1bzBCaI3mG5YzgI+02f8qVsV+v
felC7I85R571bkHDfXd/m02Ef292huuZd5+95dcFB/rnI5BmoEEN5y6lPr83jRiQ
W0hb8Q+mQBFkuO0mx/9jCu7jzgXrquSY1sfN9eOdMj0qUulF9D217kur6uFJRMGW
cFNJF8dFWAofbh9k0dPfPeWO3R9AjRhb7PZKSBcXs41z9vGj/SHrTObLaZLnxX57
ZUn/LoiRfZ/FwJDFbCBkhJEJ3lsSGj1VdKvJ/0m2ZCtV7awe+/wTvKhsCiYeU3dR
o7E1qoTNy18LlhY9VNBQ1YzsraOMVi6b6baBANjdm30kJvDn2yYvoULRa16yjLBJ
06mfjOYm1gHXDNKACqJaMCy0RfVF0Ra/eA6WfCPXGuZhVNX2S6hFZ4otX7fXTUF5
0nQRtx1WhLGf56Q5Wuxt0QosYBCHz22fWHeXO8bN3Z+kg9gAPIzyVzA89/1jhIGx
s7hqhRiLy4kl+jAuiDCb9OlS5SXg4DzSZuqrTYIPPbtR2YckkYYoMPbH0wdRBS/T
E8gNHACj8EXWfmHfePR/Inm3J8Fv4/VgzCMQoh1VyuO75fBFfv/H9r9T7Hn/sB/9
fpeqe9gsT4ps0/2vjGQ/tBGJ5eJZcvPQd0hJQEXhQMTP1JfGSvNGrM7HlN0LGGS1
p+zCPbomBH7OrCnSFxtgKjZuU1LnR3Bvr5k8suoyXNSYU/FpEIXeQZc3gpXOXFO/
NW9ngCHJkdEXZgu8QoHTl5ZsUjnFf5cYRaQTxmQxXzg4GsABbBouONOUTd0LZzoP
ZfKcbSPkVueirko5hRcmb53fLGzihoTvWgohQZeOdlo092VKqBKm9WtGPqxZ/eer
4rmrPGs+PADRiiLBVZbfDdiPHjqPNC9Njx2dHVEw+nehWwC7FPFUwYOy2wQmyBcg
/ZDFDt8ibqsPw4+ZPqh4tUpPAHMKn62cGVkXz+ntHRNKxe8+uVvhN8Z0tIpTprNm
ZHJl+2AyyUoUjz4wDZpqlBhTTPa3JmmcN5ns/HdDmnCS6Wb5hM7bcnN1ImW8yDfj
VwlBjdLgm9CKX5eShMBEcv3So49RS69EvpyRVrlKFEXwM/PaBG/5fHpCWIARn89G
ozrNMTPgxXAN9tAFbGPCgpTGPkNlMIUzJOT8L0Eyjd8CgBF1+VrV9f8XT+Pck40J
LQV39vjaFnmdTydNNq5vhLEbXxet+PgB6ql7oPD3x4FVGHLSh2Bwj5QF/Tf0/7Dw
iP91GTrs50kbEtxwAI5elx6ZP28IA2GuEAyG36yjtmncxCthIx2LAE0FPE3NWYSx
W7nfLMHh2yPGJatUwR7vECUtyFR7QWEHdSz3PVyKVDW1ni/zuvSXu3lA0CdC/P+i
WqVWxX+AXbhJ2fVvx21cFxPy06WWUBGATy4JT4rroA05O8U6xCWjxTtLiMtJiWeg
15nxTfGjctDj35/FYAmIMZJZsCtC/kN2wM9HbD7ZWNnbVlhVCaPb3ejm4RYB8So7
CzBSm2KBzYHIq/P7We+3f2RerFLNGGwUMS5aK0mmAc7o0w2rCSRNpwI3FL/4CJJx
ySO1nwM89vWqhJKCHwrUGIoW7Lp4U/Zmq4Eq8/b7Y6asSOvaP+pksvKKKHv9Gq1z
CNVdGSBKG7vxnWrbr2rfE2oGRZCjOJshnjAodt5ox9Wz9Vflm/c3wgVwensTOUlN
RLqA/J0jgilNqYJHWovCoIZC6+Iulo9VS8aYrKv2l6BxTMSGTCDEOpNJ2IUr7m84
ZMegpLuFcrRyvX2dGu5pvv4PCOIVpzGeOeC5H0hpFbiFaBRKMXzSxRryhUWInvFA
mWwSB0PMyVbmYWjQyqjQtWhxFIVsuQSAnFEljvKzZ5y4Nu6SIdOXO+McwUfNSgx0
KN50KXJvJGUjs0n/9pSgulb8XrJlxzJHIsGYjF/wfgFW4Gmx7nn4enC/SxvBAMa7
LZzbzr8+1S5xnNXDufRDxA9vUaywWw/9EvhxQIQNbxDBG16V6WtGFKAvfyH6A3xB
ruSBPIsqk7vvYEeMeRcAXK8W+0LAD+fD2wfKtC9PA/1mQvFeTU8Pyzbu3g+V7k88
rpRWqqprDyta2IOYmYcZylGPjPOQYV1b5ulubsSM7MOyq9WHnN5iE9TVzy68/06u
UljhzX7TrPUY6YVT137p7WycJ6pZA7/aquSl1Y9+soXfHUP+BkhuFPl7PO07fzhU
Q5JIGORZgSlxSoHAQRPSxisBJ1PfXhVUUzrK7jFpCnVP7ANmBfXh2BTTgtnAF4qk
BOq8KRKjZjICRiLaU2/szkGbRmkcCEzeKa+VtIaxL+kCgqp1CqbQ5FzY5h61hgpB
wxJPeiM+BVt5h3xOJES0bAogmAaJ9PRQtRtiPWauxuszPV3b1rWlIF8Q5Yg/W1hb
1QQ+J4xoU3R8VzuBgaC6qO3pIW9rGHNFpPJum6qT800cX4G3Cr9OATZw9zvuUOYN
ZNO10LOBWM+gBNndn5l0J+bovSPOMLOxutL2KR/2yFPtWIWzxqSPez+YgwoCGxas
0uSvA4yszx1ZmkX+UcfTLZniFfHx29Qf9GRWvKEiWjziZ0ph2bGjU8JbMsV1uVuO
R0/3VIGEioGYEyj/2iTDYayoyGx/MrTsv6CM5vhZQGcJf18rYkHVcH2u6eURNA23
UcQt/XpvfDpv4ig11n21KI6Tly+jIKwBzgDNGkUfbWqjbtr1vr5GLiDXq8TpatdA
7sqXD0zSkbSH2wN3Fqq14w4JxB9Z3hjWeKbeUZkUcz+JFRpEtB8JQ1s71FNtIC4i
Rh7ccyYq3MYUF5bm29SxgvGU6iPpKrbTlINKl/HJFL+cM8WOixIaQAvd0OYDmEXl
OBpxXSO6l3C0JW8ztq2g7jLJAfXAWe7bNcjRTAk/ndTmtaFZHhvMo/ZgBEc5GR+c
vXtzuHzSchYHFGAedvdO3Mgnx2Y0QzTijsUd2cdxks+OSRcCcRQDA9zLt872Rp/D
Ns9ZwcdSbEMMYyMqiKCAr9zSiE/QQFREIX5rKd581PtwNyo1zvTgd8c+OwhmyROu
UzFHFlmE8UgNl/GyOZjwx+B4g6u6p458nFFzxalM49ukWbfAYCYnC27Dou5NtMlh
W+aiW4XSNwh/gVYofUZ1AEaD66Z8wvefF6xzVKuSx2S6Bd8ex5jIZQ0aJ+zq73Rw
fZrbeW0zPZO17p/mvJE8RVkieRzHwiXJwESDf4J2jIndLt9GWej5Ol1mYFo+SxHq
EEu5dZQDU8MOZXdWkbDPK5a8IF4UYfd1XNSTtl9hMiai59YPN8AwuIIEKjO8g+8z
a3liBYwu7kMkqcfsmPZaCHCG0f+X0bpGQlHnl79STMPwGYpDlx3OktNI8nMeAfHv
PS8RHU4RLU7/pMMwer5fqP9QBX/65MJrdk2IySEXxOlvhPC65XZjhmhgWCw9RHmo
Mu9fkd3AvxM9tufeQUXQTN8mLGLyPeZKMzgricmvyPc+nrW4NmrIClsngrMtUpnr
DHHjxYxlP7zb6OOf/H6wOgYY+zhKYgnnZZz6/g8ij5QuXohLdcbU2EP7hxRg0CLi
S6uWSKBVK/biuaqGHq+7bvjy8Hn+oOy9yLVL+hMGpGHwFL3H4UK2Fmk9+u44yuul
wjPX/zTxDt6deEHNd+w1qlXbN7pNgI4lN5oIHL3G9OBvBaIFXN+F/+HkTc/qWXKu
8GD99ZaSe4Jj6ouX0/q1pCRtm5lHclgYkQnmiNUQLc78AZzzvlDn7J+OjQNDVROa
Rd1+rXgLh1zodGE50Uu0vi976ieQuBtZXJXIxdU3nY9l14zp/snTHe8Q9IvhUj7F
qIVXTz5Ew+spCgeN1etJVB3dIAgEDXNpZu9LYyO+OzAT6g8Q6MMiowv03buaOZZr
DRh2qJluMqesF1OqhEDPkSAsRB0BmTzJIz6R9rayQgsfWaLtF/dKD7ZzMwhgWpvH
me8BTnDYSvoBleo+dIHhD/I/AjvbsSD1SRLer0Gp6VReS43jsyIMMCdQLd0xLorG
0dMUquXcRAVj197hz0XGumOoONoeigtWd0VmzSMbZgOy4ZR0wd4Xaixf905pl7Aw
zlktT7cNS2m4pXiMttNzpSrWrNNDHd/UBKWnQmwTlIl7TRFdl9UpPCgNdZrSWle1
wuEB+wNQyiaR7yuyqBs/NW+y5R7FmfIxe8tK/oCbQbQme8OadTBanB7fnDgdj+xl
MZSQamOXmlOGBF6Ph9jd3isYNa54vRFETbNz+TrN3IBNq7l3l2LKLARuCkwGTWxl
idxW/cppE8aiPlLurCFtGSNljzUbJapV5ZElwdZ8bhOFVfuRkftXaWWgig54mABn
6IPhxR7aNF9vj3nh3ApdiCWd7BYybjULK/MlzX4P2672OVbvMU6Rs9Iz1cbtu6TU
tCHpy7j0VnRAhYCObSG44rOB4ypqHiKpH1B3w9aosZ/cz++QYY4jzO3W4VinevHx
wNCSFPvF5+LoxcGHBgYbnMt7+YKP2CQB57hVMhvwoqLbG9u27b+6YPIrYsq1yTm3
rHvBHKKcv73AeUxU/Y8nxabx2JRvE/8FdjeX/WvwLcbxkZt1jeJJD6fsFD6ISU4n
f6WaYJjCJOmmOI8PBxqRXVo2cRfpL4XqithzBdCyAXvDk9WG/qT0taVqSXHbexAO
Sz4c0+frsuluITI3UM7mB+/3V5furq7th8gvZzMetmmTOHHrJC2tizbwOkGWy6Y2
Jv+c4ms/sjrULK/YZojLk6Uh6n77kyyeHD44fo27Y5nAf5g1ekTnpukXulR5V6pZ
Z3UWwktNmGyiaPHHJNgWSlknltipNZWZjzzELxbjE9dU3heiPpSs0FUv+n4J5J+v
9Zm08e0B2vEL4VjQWwIFnOm9Wf7zI7kJfC+j52PNwgza/PC+2rEsz4DTzX7TvLle
2i03ArdlOg75X4qiI9Ufi95VF0mPi7NOTkx8gRGeZBTOdfnHydMAE73Hl0a8g85x
HIBRoMfkNkwl2Ba5njmFL98DbT+zgdKrauV32q/4zxDRPXEIRve9oKdeNgIKP/Qt
W0GMadQ6048K5bwuRXzSkvLfO3soM093SwkfJX7WyxaKj87kifzTt7DGYZBvC7rr
35Nn5AljWMs84xyfAFCczZdPpnGw8BxVOr4Li0EIsTEDLlB5SUujM8BW+8RW6QCP
aKihCieLvDPa656MS0YlotCTTvCR/1eHtp7kLn5WmkeIeTQ210bHsDNY/Abg6WGQ
AvXbM+ZGQRAATjRgpvgRzNfGmoSc62tFzvPwjz2vVM54pP5KlOn3PUAo8n4lTWkC
SA0346LLG1dZCjF90ca1megmgrx2BaVPrUGjWrFbhmVP3RSe9gkyqAlm7L+AmvnA
4hpUbrX7NyEPIrBqtyzL5gzynUPPAvoLAcUEV4rZIas2eLJ5gpDbteviZdjZszzJ
Y8gxwc0GrNiiShcQv+gwi0vAo2+J7MowfX+4kA18eDlSBNvIkgFNfE9T93+AbYb7
MQqjp46KGxJ1vb+HOQZupWr/6ljO6eEzPyeMAou3bXHfRKVX0ZZQT55UMzV6ZDWF
98mljUBKBbC5vB62L+7kLPuA20iMuxAhlFPGWbZAIVZjQjLW/o4voTcjJeOfHkBi
X7UGxPx6FyFdAKNElOSGMtb4xl0osZuluGpq8rkZIv/kj6bzvLRZNwdkQd8zrYlR
nIuCkDJu5L3DOks1CiTOcGlHZYfxq2q1ac5Tv+K60jc/FkCwSwF+bHWCeIMsPwt7
RuSbrDZuyJ3wLKbrc8YpHJ9sqO664mEx9jtTLDJofuOtJj13WQAsv+JIOEIqTtI4
EMTU22fFfn2pWANRp7bEMdYjIPNzkwkKiKfTTr2Zix2ANa9Vc5SWR5z9ru9AQXyH
Sk+1XHaeJ8WoMowpuvJZaz5Fw+aSPLLn0n2/VV52UWX/OHKpl3tCZmSzx+8mQTRQ
wbwMoJWE0IrCLvCecrxO9/CHpuRdmkbIgo88GPCip2lb4M04m3NPSGNQXS+kWuFQ
i8TjNqgd+s4ZGlxlSSOCMVpuCtIj2Bwt6zAxwRIgtHKtK8Dl1bsuPkdAlmQJXwul
yl9F/znn5N/1/nABnqnxokBx0oA8vm6Bc0EbjBQkpOxBhmX+qe9N7/pQRVa4TQG8
+yCCkuU5kBmkuCUU736+IsYfBwvAISxf0sUCaoEGyF0eJ0FIk1okAcxIWXtLSybr
oYM1wZAsJzn/7HHszJbOjK8fe1W4ASjr73zSaajJP/3/jQxedkpMPS0gsuO949gh
W26CFrB52SkNHs/4nWwKTe+v7mBT77i6NJ9VV7WAvhnvHsGc5bcuXang4ALpYm3j
aL8lq2BXUbcae6k71UetpZ2HkTyNuyS7DOcXDfWfkhLOMkEGhZJBciKu9Ll6psxL
zJKkcKshK9Lu95lZPFSjWcczAeSn8IOVOBYoKCTmZcGKfOAMM99qaMaoUkeSpUQe
VfmvVKocZ58/03oNb6sepRHjEF+34VzwiFkzc3E+9OYXuBtyQiHgiYgQKxzAI/DE
XM4d19hZ+TfkmmCB81y/Xopy0pg4/+UV5Libi83iPfbDKEgn1fVQYDdhTmYiPqA4
Ejnz8XVj974eNPZnWUmzlSfSkErq/XwuPJGUWelWqy8dDkPc8N6Ssid5UwsQU0gk
vOrLb/85iVco8NIEdjbnOc2WOjd3dMSJ2AFrV7y650Pc5yzJ3sCvW3zyaQTTD2N+
MYqmTNVbiN2c13jmtrFbpVmE7K1b0BLsmJrY7q4HTq+SgyR1G8WSsc1U1kKvcEOH
YAFRE9EDfzPGkqwz21TUd4wKJdWwjt/C3j5AIhiDqCJHADPB9a/WmyFIJW4IAYFk
4jHBlH9mGlAN3nsB8xNWxWEUW/xN6mV+t73hWavmxLB3li02pTVfY4oQAu/jnLKn
ByU9MN7TZwEh1Bhe6jjWbAvSXcr7NegM9ClzH00b5D0CdTBkKN3VNkgZ2pyiGeP+
lJdP8i4ubt7EmtEoZ49YveAVcA7J/Ngwn1EaPkt/pXntiBHSW0/eqH5iLTTajAB4
2UnEUo6Gv62SQ7umtKOte/Z/3B0jOqm2GnjTlDtyTahWj+2gah/2fsW/3Djb8WU6
ADScmKvTkMMDh78KYeH9JGP1Mcf56Pmd0LrQvUSkrobcLa1pJYULdg0Vs5jt2swX
jRac/czG6OPJP+9kiEDWY4eYZ53YtcIivhWTU6/fTSZFr0KJG3UsHrG4sJY6a6DS
Xa8fSzenFEKdBMurWOHzk7fqhJvuHIsJ288+zJCA+SshJ3yzWmJZOWdk7bfAqKw5
OkC+v7X5gvuJmWi67sg1NQCZkM66Z+VPgxmY8/LzviRydL3K1CYMqI4tsN5iwW/Y
PXCFn5aEFFRdb1pO/EzUrZl2WI8U+nMIIJArdn+ZP47i9pcvcDukLJp2bk8GZseV
5LzZHR1H0aebo/bDeJMLqmVSqOxXcTtQCMmUBcM/3o3kt5G36fu3lc60uQxHJohP
TRMfaWeLpuB1nuut0xoYCiiCXLRl7pVl+VVoKJ02mU/JdnmdoLIHBLfh0d4O6VEQ
VWh1WDqoyfx5HwZSKId8jwyMlqsS7PZG7JfiOlb6bQR8gwhBhxc5LRjUrbg67ac1
YIR6o7sP0W337PmFWCkYMfgn+GNy5x32+DT3CG6TUI9O2DB47BcpcOXXuXOsT2oL
2M6RYudXN1oHGCCPi+i/91iea0oHQTK206u6t2yg3Whqc0h9ui9WJgOiLZeZXp/c
OTVjtYu+XRr38OMu61HhJejIceCwMFRCrOmCDN2Qka74hpON3SFtKVlRJpZbkRS+
zLDOjavfwJddP6jxKbGpJPzW4goYrQBRxk1KUMbjtVopgpXId/4UV+mJtQ8T9KA4
o0/SRB0wMSSFcVT8DuwON7ma4qYCj/XLaFIzCeVxdNGsxM7RBcgSN8GXxNsfednR
+FWk+Td+zzuYTNjh/DaK5F4+IYdOwzUGYitYTqh0qFYLLVAQbwChxzn9twe30GJU
0bGfBMHmiSa0VPVT9yTs1+hgZEzpAMyoROO+sub3ePO3vR1tTc9BMiThJS3tX2uq
8LjGVTWmCHGx9eF6UOXwGyKpACxBUd32Pf668eD2mcbCYolIUOyeNvOuqgZPIeuS
zUdciOxyvWqY2zKPTi7V+NsuWrsWCISqty2rRPinr9UUk8lqj0rwitDk4WqdZtl1
pQbvcpfecaq9nb3ZRQIH4PgAetpFjPllfdm+MkumU2KcEb4gs/T5ZPU95rAOGjFG
qb++C0wEIClhHt9dMCRsxy0Wpf08Blj8I1BmDKUSiZ5TRGBR2KrHKBQQ+sgaci5a
X9ZDDdpYOaT8G0BB15xMZPahP3Ce1XJOKHakJBQsHryYuDhjdi5C8u8lGerrbzhz
+H4S+VFPOB0B75wlWa7j74RmKKY/h6de2yevuMqCFw85J/TpzuqgPZHx/UMLcjDd
kLMBSx9lpS+4jjuXaDUKxloX2iT6sBSMEVxgJAObOHrdrndWfBVJ3UEOJRDBVAXB
fa33lv3UsNnTudwL2Nyfvp5fjPxnGMIWrpGKxqlnoz7y+TWTZ9vbAw2b08L0T3pg
QbHBysrxoV7Czm626wtzCIa8eknqF//nDURMYX1Az4zTLsRQUrdcgMFRSfoDRoK/
3+YAa8HdJK5iDXpgKfll8QJyE5jCNW1iIU9BNyZTvJ/ek5mnffqyoLByGNKyrbUK
yzTMlhtpsx2qO7s2mAHyhFrY//AMfES18TcGVzMLvwSBBD+orUso88ZY6rhPljTl
O2aZ2Jv1PGIfk665dxDxgBeuEIu/nJoJTSJ44vLlp/SFdD+5DXObq3BkZP+L+kLx
P1gVA8UAsS4pxRiowlKq3LxfqtTyBzCUSsIAVzdDlQ4gUOU3nd68ZZ9vBzZrj648
koQrSVzEjm0yNlwmsod6yLqdnUSwX0ksnB3RRz236vRhIt8foJJOfGPUVupF6WfA
B/tzeaEcAQ6kJ0N6VELmbcJRuL2U0bxouIeBDqYDtSNZqbSKOKDD9NJpGAOYAJvP
HEyZ1kqKOzjbUXKX3MKCelUYVL/oa4Fsgne8PjMTnVuWbDVUcuwvzIP9JQdvl9Yx
RXoJcrvXrBJWxAB9zzSR6LMoXQo2dF04A/g2JsvNJQmYKSoM/aGtwtpePHjfAIX+
uIsR1mrwgdbniEKYCMz4S8A/E+3X99wZMX7bam4xlIDWb1fYvR8yGGwAA424Rj8L
Xwvaw5vpgZClRjsilkkCc5j9kY/yP8GLvGXMkEap+iSahp+EA3z92XHkEinVDv4F
rkuJD/I2NxOl2x3Cptn8zVNYhEYTNFwZs/YMLdbS+xB1i8PcM+EZtAAm6uHeVh7J
yl+RBs3zP4qhkdaZY69Yrz/AgLsu0lnQkhzX1S5yUtjnb0NLo/t6v+TBYZU3zv/V
aLjruVD5TFzGKfxgTbAdzWSeFG2HttJFycVlSc/CghLsEc0rr0X+8frCruWlkEuY
8VEtx4P8jNCxbVsxbT0fISrEDn9I4jzrrVKAwaosimy6hSaXsmuRkiZN2dpvTUjC
SJoj768Cn0GE1NqT6N4iLpEMMmO9LoWNBb8MOOZGOl/TjRyjIyACs/gGCvUb3Y8k
R7KrTbz50mhIQ/GFddyFyiymxWFdTZroI1k+s12gCGusZHa07PMB36s7YB/CiHYU
URX9hw0rd2F2N+AKsOS/fN8KfUpeKdjn6K3w1BLDpX2jO/t5rGAJmpBFk7v9o43I
ePBQytrqiEQJTC+4s4DbVmti1GopFUb/m75VgXZyRVg9XRb7PDhxPUyh0ETI9+Mm
Gsfe7EAytpQYb1yCxKMjA+NbnCSmdjmVIZiVNHv8TCx5sidTDZvO9xnoRJCVWlBl
ufXeNaurP8l3tvrTf0bsNwNrV3vZ71hklEqapOGc1i1PCIicVTjWyQMPoabeMG29
kHYJcTd1PVCPHaKu9y07E7UMFtlbCK+5TnnoxG2Ua22FbaDqyD57FCIO8AjUzydY
EXlRvKnCMrxbMadTaXTn2jL5XDpjRPQAKoc+95jH3dCyXMO4ga6wmNLS23iQBgDf
6K+bAcpYVh3GktGtUQYRze49W4Fs0q1WvEePA8HSrCs1Vruk3Ld6TgtFDioacSP7
DAyMqjepL6WtbwCT0aqCb6EjgdHgx/45pRAQJVFqzX1dOOGUTyiI4oBuiqltSYbK
8TjTBbU68fciBCPhcjDwY8VG+RJOe7N//dqdcYIQKhbbzw5yXvmeIALprq+MYvFs
CguN1Wv214bvf0vjsgynRM10kb5CsrMGLc5WanGhoK+FiWUvNAGc2LX4jmTOamgu
LCqMfOp0LyZOiT9Y/CPEyTHh2XnMna4CkOAVZnnQ/DhwbURh5M6xb09+ah3LOZ/J
uWNsUEPl8pB17oMjt4SwHMSybou93b2hktNsCU2ASmu0OFt1OFUrgvcBc06L4+I9
HoLwTlMQteHXSla6BpL0IJcHc6NNBnyrt3eK+b/X0klASPLi9pAhm7dTgtLyFE+D
kRN7Fed3HocQouTO8eOZgYb3+TWAuWLjzEiL7Zjw5vmH8WSHkudAgRF4rnexyslQ
ARcuO0A/yNYopxtQZtHukpeh0yVN5dVE9cDOtpMBnprXmJsqw1cE2l0kH3rkY7hV
fCl8zNCsDBqGWjlZ5c/Gzm9qC01dakW81RlzpciDj+xlsP3NdPeGoy5NTSJP0TDB
s8bVXWVellb9Zvk+QKLMIWXeJfwDQqUO1SVNFEigcCqso19PIOE82OW+0dsCO2FX
QReBxegu58fKPDJeRdwusWCsF5Yae6BeOyp/Eaddqbqj6qwFanPBg+6f8MLxtTEz
0aD56E8br0nk6hchWbayuq73BlYIF51VzFo/juNcf1B9tUT5HVpXPH+x26XEBhXh
XgjkInobLN5gd3xl41dEYmjpZpVNON+5zEmU2YK+ZqhEQ07CtH0aGQs795Co5ahG
oFnOjoliNpJ9J0AJyuhQ0h+XJ59WY1Pn1wiXbryc9QWugA4CaOzP+iJtTOaSzHHE
oHR8UmWq6YRXaVW1FtvKt2LhmWL8YCE5kvWcTcRiSSHX41V2tBNqWJ2YHpj+Smqr
nx9z39hljj7dKxxkwpKzrsIpMCDjKDPUETWgjkom3XY2SkX/jecH645jJFy+D3te
qD/7EjzniXwY1s69m+ZNKXObp5iqp4kMGjCai8mXp9p9FGUl5kIUcBTsohUAbr0Z
Ta4/fbwdC/pYllbtkTqAg1xbk28ni2RF8yg965CokPgPolP1eB7dn8GDKG3MCqnl
SOJbK+YdqwuvIxMuEReez5xi/na5VlMePNyqah+lmeNfRsxphFwD5CBAQqBNOwZF
sEyOpWHdHDGbMbRavZ+uOYd/SsKlnWjGpBoDUWI/CyoEVCZaTMDij+uT4yqZ1lUD
lTLtvEO9D4Q0eWl0hHGMfZ+WkXxihQ2tN3couCAqh2hJGlPAXDcyIzlpWzMxduUN
aaNeX5YkiF3xEbxVmw7Ub6+5X/Dfi9FYXFAwCNras9f3JIEYW+OYHs4LAuTXKMUM
NIc557CVmDaE9YxGrZU3xhzluU01surCbf4LU0uqfvAvBgVOIiPxt412gAVlWdZB
4fDo3gZFlfno9O2uSj9mFlGTZc//c5jJwg0KiraYRRpW9Pu9bSBrDjP7fQdKEt3F
lxTrk1Cw1XldgjJR36iookGWfDNHvN6txH+jgtpyrRNK6/xiemo7fC8bjfC4c1Qp
2Ew3UgqO0HMIgYStQWoo7rQaZV5Wz3FRc6llmnYI6pxSs3Sony8hCEwFDWYiir4J
K+CaTSOrrPqG2ZWd2WBtQVqsLdrOAzQoLOOYya1R0+UahOypcgc/PTNIak2gYLuC
iI8qWUiqCpgnAao7E/aWfn9rVq2t+AIBeBAUK8D7gbaytklJrXcGrMvdtiOGdAmL
FgTww5fVuuzPcYr7dtPeKtGPWtD8lSdOpJIpKLT5lsSEDyfO7OiAQmw6MJ70dCLy
nC9vGr+hvo/GaEqIyw4WVYgad6JPZT1Id39K1t21uqevPapVdeMSpQ3nHO7v+ctn
JnPRUa28PfZvFLcMbSfmbf7wiWfE1mDhq6NT4lEWXO8Pb3Fv69tV0ltYMaX9pdVN
dI3ma8zYaYLcJ/lJtz01yxSUu4uEfzuOFogMJAYQStuHhkz0E1Ib2WUHTaZO06Lb
xkUjiq2nC4+Xq65iRSfhUf/5E78v50xr6P65rs8ekOWcHtMajjdprxVo0CeoVqfq
qj2ksy1S2L3F08OP31lEt+p4PYnWjEjoxaT8IClPwOttFB0kxvkneqfoc4KJ/AP9
MIhR0PV9W8+VfY99SCC9dKn4ZieWgm/fCluQq+sTK4LB3Iy/nTGTdKdDSnKapg+a
m4lIY5xx5RdYFDZYB9F+dU6lNTxUhTepu37f25b90ElJj2IVPYW1vVlc0xqpqIG6
lG8Df3BvX3c+9x29xmNwQFqgI5uKKjsUvi6kvQ3u9QXVuXrTKoQWR4oMdC+2A9xN
MmocQJ7Min0fG7bI1zABiLqcJbJSz5T48ijCxbtG4lbW6HMTrWHXnOcOMlUl73VN
0jASyx47ZFfcrjl2khe/hPf98swEimmPRHYf3NIOeJFeYnGX4/vwsX0RdVPi22m1
wyWkmcaDvfUQY3x7zGQapyhMxe6r9SY+Tc1Kp5bgcQDjhpcVM2FvHaFDRV501zqQ
aIhTSkI2qSEjP1ZPZk0DFyX3JuiSdrNmEgdEeMr2L1uGEIBtoFG03B4j/3lMoRNJ
l5yzNBaVn7akHBukce4Iqu5I6SHlSaNqSMFQLfBJPCopRpvdEIMDUfyZVtHwkfMy
FH6OlmIo/5KLSKg60596SVN/4EIa+jxmn7eNZFJls9w7S468r0cerxkdk6r2UkjX
kAUI0Qkcz0HdlIB7YdzLhicncfX75iGhLljnyg+FvnbSrgObsgG+0v+hVsnhHrPp
btHyJ0WdeAJ8GAAjfcwHc0PANoFh8LjRCp2k47w25HudTIPrdkQDCyPRDEliDqa4
QOvQsMyRkmbBOPB/4eZpJzpvk6HiAKc4HdplCp6UnPGQ14N5JZmZEa1EWXQI93M5
MZ+PKsl3aoqX6+9AR/NCs8yV8pZXbdZB1qHIcNAWhUw1CF0zYPWyNX3hfdmPC+ta
+JeUvOOdMAJkb+NqP3rxIHCpxkN/OBgPh6kZpx11TuG6BKqZbuAC67euxPSAbgzp
xRO7OLQvw3FjAKy3WxWZzjYDD5pfyuZYoedjO4VhaHFxQt9fm7U6IC+KokWPujUd
lq6tI0laQSdidvY9Cuyzh8N0ssFfGoFMIXKnHhufXLY5aFwbM8roM06Lu+h7781y
Y8M3HFkmNSuIdmyzb33w/G/V0VSQP1vn2c2tj7mahrrbSzESbuYXEEkqnJ9ADTmg
QpyZZCW3FwAtVHfD5Ch01OPqW8JULUKQPZzAu7J3+XOcRMgltehTMaJEn0n/Vibi
HGM1Jz8M4wmBiVZQcaDn5iOQOI0D1QhA64wzZMdGrQrWt61dgHmxiH71YZAs31ti
875JGCgVrAkPjjRG+2zgE3GemrZIAnsvgvUbIaLEodopPUw6lShRViaP3qs3OGHc
tjRX/stu63NA1SmwGvavFtUKJfd9LjWKaWumJa6MVyoWDKQmdYmsKc14oBeG0I+3
/wyJMNXXaHttGF2+J9erxzk89a1hFpJD3gRt4+GUzp4Q2u3PiNNGf3iLShH0t71b
MTgua9URl+89uEZmb20wv+ETMkU2fcKZBY3OuT2LOds/V7UYAX4DsS1mD+P8le3F
4z3u/vR17CLHTx8viZGIUKfnxqOUzH5vt7MJgHB+bGuXVcEmW+ZefKitNGwZPKKs
PjhnZ/yL3wSirhZ3OHE7I8ozFKEUU4z8mUAsuzhpn8aVpkyA8ai3sTZz+rKqkxW1
J1Ww/22i502aX5lVLRSYdv4vM62HYap6RJ2mu/LF52TW/kJaKfVrCNky269Sb2di
0g48/5nmD0UEA7HOcQ+JUcBDFcKOrdbwvN84FMxW6oIztGGdqiyJ5+Rw8hSYV94h
UR5uwRaLdOJFkT7Ne5Lef7PnUhw0TU2iJ/uzCqcgc62KEwlk8YyDXkP36v4NopA9
7ZgP0WoDSDV1fdtbfdTzXGZH3+c0m5AejHWlejodPRYUdrLfY1ceJ2R3VMNy4Hy+
pA34SWSye5k7qgAlxDLpVXyyxLxVyzPcwUZtVtX992CLR51dCupC7PqzO4xOWB50
Q8u+9O/qlmm4sXTVdEhw5NA5I3feYx6gqXk/ZqQiibOizNC5qQUU2wbl/PNRcY9W
d/kHhTZ/d6597AwBquoL6NlFlb6VtbV4MYceCOjLySRyJqPXvV6QVnuAvdbAhHTj
+kxI/t0ZJxk5WYEOYieXAnn8N30uviwBF9A6vS+OCml56Q7z6SxW/8h3dLLxdine
efWewZIF38gMftT1tCUdElGWbE70y4EwlnVSByj3661iRXhL5sjqe6TNGWXxJsbi
2aYncQppRmCB6kkDqfJpX4agq+dplM0dee+pPAK/bu9983JAruhuCvkhP6+I+gy1
n9G0N3kyEaO7zzp2ZBvCpHL3qPSvT4PReYa5rK3yt4bMw3tifGxOj2Y71DA6fNTS
TAC2uWW6tATIuAvu/BydTdZu9etxwK8wOwL+gHLZoJ3TZuTtOdSaRsZaUh8XDnD9
qiULN46mI6TH8Zujnwy1s73kGElVNJZvrpH71Gv9OH/j93hRZAcgNykOOSJn+D0P
MuFhxsncqVftrk//O1j42jT0su46TU7elvtbi3lAhEFjmUlqpUSBByERLZNEUVX8
a7nk9c0tVL3/0G5GqjELIb5TH2njjAPmT/HuKIQVSXImABRFlkg4GLOVaWhuGjTj
1SUj1ofRxQXSiDofRr9kLz9yCd8WdJ+YDTiep/XFqUwtjOUnpkTEMku0KxGU/4Zp
VReJuB0Pl/HuzwKKt9N0/t9Jjlcej4tMqjzqhzs6CNylFxUSsjlvkHA6jLn6nd8i
mg7ja5olXbl9dQsBaz8ifJ4lrlRsjlegbEMKeGAMfvTsUOB/HxO4Z5O1o8zXWs/g
aWRIrA3/Jm14Ub862i65FxSVdqPEyVyorgeNip06raVDFEokERQ30n4oQ5CBICs4
at0smVoQz7fvEFZCja/g5EpF36VtUT354eEO4cZSyPF02xcA9PcQqiZir5TPKKsb
2iiqMtNuNHTRtuf4U/ysoBxuHgCSg/0728VRY+HWFjjYYxIsTlBewJn6aSwNrmV0
0qUg4yOauxlutEV4IZxLpn0Dydm8DW3SfyLhVPIDYdCxcyftD04F2X8bZVSUZh83
cAaK5oZWNUE9VW4UdGH8IEs5ZsJZCjPFEWTWnaK9Wv+IYTPL6Xq1Lmqibho1ePIB
b7MtNn+/GJX3ja52+2OU5xALNqAwU3gBSBdnZ1EGRLcMTJ0LzBJS6e1WbmbpAiTP
NXonp0CvTQ8FrpoMPFexrtFoVD9Vn66/ctN5pLyJH2XK1LoHV+a/uPSh5V2lzchk
bH5XEHv5M4Y50aFu/Sti+B5xiiTs81z0ZXkRY9DCuPvP3yS5t7hOMwD6Jba01ov+
q+30qfDt0mIOn50f6LzGZX19YcGrgDZVksZFt737vCPsGxaCmU99GdjhheGscXPz
un+hGTid9xmhCdL0PR5kvwsB4dZheRbyHW6+ukpaWd7+j7g23W4bj4Ki4zfGIsnK
UsvHutCmxDFp0H2Qo0nDDtctaQPHGMO7n+84B2QQMBdVxsDDjIgU33E3l2vhQeV8
hIrdUxbcmaz/PtGwBceU8VPx9pgGdQxMFQ6D90R8B4LkjF+1wuSbKQkMiXSXIv+A
mD+rPvZHMRqVU5nJp0S3agwOketpf6IDg16q/sjRYzi3yBJ5Tzk+kcSzH2a2VC4v
gSCWoEySHI41NZGxWqdYNNzdOMkuicOCx4UmtCtp3FFBptMVXNKYsLgjcs3532SB
AxZRwyh2JOH30Y3Y6ej1OpMrSaqqXR8Sk0SZ9ztEx294jo4ZuFY0/lrcUUVnshDV
zsGAKRgl7HD9xc3JVCGCPdzo65dsFiO66eRnAAfbDOwqKPrejdl+ju53aXaHWNfY
GhcZlE4nT/cfqxynkR0KXbFT7vuOJAD3i2kVu77X27ka06hn3B5ZKi85nW9iiCqa
BlejGwarzzuUDYb5xxsWabD6HSh2hl4GXNGND75tN1Ml3gI2eRibFKe3l/8mDgyq
BnPJZAZvGEBXFPwNeDP7Shx2dHyz1lcI6XEm8F6HLuZ2GRsxXNO04u2bH7lA82AO
au92tWG9m+HP6JHtyM7PYyDCSWEC9NRnohXiFcvgkECOVEYWeD2j75tUP17PR7+3
3Gzs1OaqLlsK6rS0UfS7WIuUcbaYZFooBz7K3ncyEfSLdOY1OyJPJSWv/5IrDp9R
5l4fbbgAmh+C/Gy6Qh3e0eJsNVTaCSVBgO8m4Q8S3mLidRA8U4Z3M5yljxiOlxTV
deGVYA5TqF3qMKKLHoxv1uvzydag2PPV3aeP0ufhLhjASzMOUj24jkzSXagaD4vK
BVYMqRyGjK7zaZ8TeQvG+sDFXqRSzZW9f89SF+MTj/a4dFQsJHGEyYrJp/+mzzL7
OrxHsr/dWNls7aAN7MfyOuNtX7NwxiP8pDT7vFCVzyayALcS/Tm7Ldq0lBFwUdsR
bDGqqkntO8zC0pg87Qv9S4J6RsuCcORksKOLWeXqQRcRp71SfrPXM50JejmbgBFW
KZjCWlxlwPAQQGVT0ztYUCj9N67WV3W/I+GL+V/7p6z72ojZarxBO+dwb/dDKjmX
MVmPxOB9D5uYlj1YKHAh7uGOwi7CQuSA3C7/pqTdxD5N8HUvvcE7DKcoTiXy7aCv
hBT/20cmZnRktCdaWmFAsAaU+Ph4AMXdFIi8lUS5Kw8ZppQ4c/PBg9ETysgmgLC6
D3ry6XibnLgXY7r1y3e+H8wBKRtkzdVfxM6vy4vr1vcof2sYmT2tsi4yOaeA6h3O
Q9iZHpa/lgnhwOuiF0FTFEzWG8UDf9CqNqLem7xh8i+HiLUcQhixXzGQPFOC5dB9
UIudjIm2QrfeVBLl/zjqWJFuhK5pAc+o8lgPvG6DTWW6DuOyMFEZmEJWDazF6Lwz
Ib0otqwG1gthEKUFxfc6+97bT+uzXhi9Ely6Zl2UL6cLHqsrfHhSLrk3FMkpntSZ
16dwDWBLrolL0bYG2gY2YzlAcggVFr5naDwlRQLBDhJli8VGNwZ4aFq49NJFksBu
UbJe4qSRck2Mu1WgYa+vowj4NN8eUHu/nZriMeqDI0mGpwWLQostgsxO+DS80QMy
G6vp0OrV21FM262O2lcv/EunKNJk/mwkzd3lgUrKixX7F/xE0SjEMyrQOx0jEQd0
Nz0b2kFGp6BIoR3RbTI4+nOIzNEQW/zN1AleGSMxqc6qOWcs2mVbIFem9TDryQsl
EnmhujR5Rei/aYgbPcj0Mhr2s7E5JEFtzMRTZqnPSoxnVCa5bs62uAIOBNX0RxGS
cD2Y9WssTPfEeDpXWw62X5kHTtTeS3G+8A01f8txAaRsPYCcdPiEjwtuEhw9e4Tt
JxmOdQDQ/btSHP8lA/jSA/Sw30nv9GHgTh4pVq+XWOelOhjYntRXk7A4lLTJGb4Z
Bfyfxq1O80knNuY63vnrWmTpI+eZIUk5b9MohStIwejdgYUqSQEDxZlHkjeltufn
Z6DvjTKdY7nt5aa5yIRCAZFtvEJVPLiI51IMSs3zM7vZq5TQoYwSn1Yiqj+Pjpks
PMr+xQ4lu6Bk1UT7XNv6L8d0j2vapCH78Zh7zFUGqy5sG7onRbuJ3BrA35tL0pZS
9Fj05R1TYMxJy0xh5rFEFyZNL5Z0q4wlbGNxzZ4EtPKNYj5IrL9MVPXpPK75BbUy
6WqOqngTKgq0tDq1tt6nxJCQCgbwMXnJ2ecy+6et8b1fIBj/4pp1R/48MgCufSDH
qiTjMeD0Hb3JvlCbHa2ZNeqt86bL6bMagufHbXiqGHXuxJ8qHigQQMiyZx5+Lrhg
tgaS7VlOBPdX0r8lNKyO4iGVy1xP7kvO32EBP+1GkueYO52PhFHejasQf1Vdi+fj
5Xg2oDOWUTNKQNYs3Vd3xD2mFjSIn06qmYwXCtjpFUKW4+vrJ5StoEWiXM36PSuB
JMC5XL4jQ2LcaYT+DInKfk+LXfxjo3GLlBGhD3aa4/aCEsBbl1oqx0V+Mb58yXyK
0825bFnPOUrFj1Tj9KjZIZN4rJko7L5sMK+/l7/n1kX6IpKpThguRqPI/YrGiSFc
fqGdjk07gRUV+R3h/ZN1ks+oaS14Pgrkov8j70vUiy5sdAxu7LHBqP1fSsi53pAx
sTjh7O8QhspmDauJCj+YG867Bqlqee5GB+vbUgrByxU0m7bvgnWQTIS0T11pyoNx
QCAxLckSKBvjacm+qHXTAGXAorru1GgUnBB1Q5AQuwo83wXGAtrzMGrZH53ee7CE
vJE3MakHJmo5cAU70xFGPOoO/UpLx4PEH0m9y0k6SO1CNLsCgz8aB8JX8gpylW1b
OkBcoJAxKS3qhqJ4v8J1gsQA4kXGPbAIsYsUsOXgGf+uKq2vow+F0Y9HpF5Ccves
yD/5dJUL/ZR8CvJVuE82NVHKSv8D9L/lM0qjyP08jARyO2VyVrYCKr9qZbr0fzKz
J6uCIG4BDxJIq4UIAtW7GPCBec3Vo1dNzpp7A0DWEnf+LuEv4uAiRr3NW9W58Pdq
EAhFl7LaZe65yjsNxmKeQQ14ydL376SMzcEL7Jdeh1hw2LH2DuzyvdoDtqKOnbPO
C1LrgE0PF2vSsy4ChzCiMPzj50oVDyRL0gT0Mp9ZVYu4FB/DnB3MWd2gZ7aQQy0z
IutQiFCap0NIBrGWvDvbU3vZAeWgO85VmnSY0bV906RY+Sj/dd7nZNPm+k0ERQ5P
RRleX2n7FsPD2BBV2Tb7ZBPE97HH4VnNEYuBMYiNw/2GgVMW4eUZKFGgek4Vr/8g
fOkcx6GP8udZiUnnct7J1hIK7xJXWXCfFCgjkL3HF6IUDNatG1r0uruFPAdVvDBJ
60P2GJmxQnK66V0eewzYdu1/8N9pCh8VqIHElKQAtzJEr/SiVTWnUdWZmB9SoRGH
HnLkeyrYkgSg5zSPeZyz6Y+twaxX9w0xQzi/6dyaKdHt0yJhk4nTadh2IOxNQPyu
Uefg0UHblR+QCzAd9flCs79WMQcNNOm9HAyxyW7W2T2ldrKqQCu7pBfp92a9h33u
A/ad015ffuzeQRnRF4tDEWeP0tSWkJ3f/AsfJGBOSGn7ozH+t5M8HkPpZudcUD5l
bvMCM8rpcWlukvIN/s0epM/DRBHrSahQ/D+Ift5WymzwoxpEi9i2A3IWtrY0vwXR
yn/wWGphAlBdqvbCs4TCHVHoHHJAVEWE5HdCLgUmOiCON7cJt9vaWBMeZPy0YX58
v4wsSY4EVAYZBlWEaKrAp7CT2zPMCp5KpjLxA/iBVavMY0m4S458siUuzTVRhFIu
2aYz0LmqxuvT4Z8y+0+0QqwfGRA69Bu2c1xpd8qJXZloeesYAo+aeQA5Lbm4Ry5F
ClqfTweVOoFuMd/M/pxTts0a1AM4GssPIt1C7iv0pK70jdIRoJtORn7WbZ2PnmW7
6QlZYvjEch8ejYnwI1cs7gDnOnBuWdhuLmaoJ5a4yhrSlNrLOp6eel1k6WZuLfuU
KtdetpExlnACwzmQOJdmKBgEppCa4v7Clu3VAxQuawLW966vVD/EBc3qJbcSwdFv
NXsdNva5yogXOF7J6hSmT+7P/HExljxtdrjFZ2ltLbY1+UY0BSvVEunIi0v1++ZX
mWhKPh7AsAEgRcBiJ1S0J0WQ6QSASX0r1RrvlZtFAv5cYSZYTouA0SROmIgs/nTx
IoLPg1fi9mDWEaY6lRTUzghtnlUurv1BZnrsN7dZJDheAHuWvNnRudzLdY/wB3o7
/iPkYsuEd3+n2Y8cEdWPlHDaR4ZxHDvBvWt9Qian2wWYy3vCgXKNnoDoxqmUOGfo
9FMQb6KYXOfCBp8WhXQx5wK33YQ0c0lxPp/Gb1NSuCdobc/yCgPLRMYI36/Pww+2
jed+PR7x7h5dRU/TVMQslNTghvysYnH0LNo5TrGqDW1E/zrkgwK6dKGNnXQySgHO
tfuapTMMt4tg/2O3f2WmsMDkvJCmHgmjeVrEnFYR7z+Rf6erd/7fgSdNl273necv
bVE5gFl532ogYwwnwzxk2erjoQ0CgnA0BemlZ9cAsHTOWeeBSTL78yUfNYGEVeBJ
M8uVymR3GzW+iDwYODlLrG00c2toxQTxTTP0qtSnyQ1cNUs0aBbZMmphEA9qbhYw
k/bQCQEVsgUxSG86/YFeJRRt/OX3TNIm3sAk8i+rDNiQVfKRbcWhrccrJ1VM/+6m
yQ6+HESdrSnoIZ3tJWaaKafSFr+yk2EFkm36kmkqStWG0jBIv7aoPuydd0ZU0IlT
sny6y1rn6gDWamf0I1QE72gn2haSoTfWucHrstC9V12LusGVqaHFJDiJGYiq+/wR
Ybvy4ZiT76iEyCmr5JJOtapFHs6cEVyEjWikQtbXAU89bfVNLzl6N1gqLc1GuOi9
AFeWDzXnPDkc8pYeRNUMrh9MKwtPHImKR+ULTXp2WzCccpSoLprEadPcGsN6eO7R
/6XVj1FstM+sg8ze/Wu34xyZtOfLdUL/OqOYR9nLka3k2z2iNhC4sRnQm1ehuCeH
ksY40v/fow4cps+Hlufq3d3SB8Hw2O5Bds+kBVbKd2jk6SinFjKvk83aNDZn9qWR
OvN6XcZcUOlNMEBxQL6qg99kTBtWjeVuLKIQ7WAubBfHfKcQKXeYnjA+qfrs6D/C
tsEQ3Iaq75jkI6pV+WW5iq2M6LkuCObsBcXkP96T+NQuLj980MzFgpfD1TtctGqM
tSPnEbJAAsyMDWbHuvh0EgTRmazoe6HVyj2xXLwRx5lBclX0I5mfdsZVqdlfw90j
BOsn1QPBoBsDelr3jUQiyiSK1aUJ4uoNDDgM3VLsd93MoTcEIzSH1GmCY3chiQmt
1mZwRWXIGu9sRWCybm3Eg0pIPV85WxNGfMdBgUpUe9XRn8ZbLvfzKFAlEl9ZdAK5
/kuG6RgDNFfpTeA7B63C1K9pgxsBCZc2ahfTNzt32gWAvZpkop6b0S4HE6Qi/0E2
CyYrxA6Nt8ddS2eOWi9b1iVmimfzrq1qoq3GRBuE9jPCKGornZgOSe7S49I1f8xm
nC618+EjTekiHmz4Ax1NeHNCPUl2CjhAg6IB2sHzuqLHd43o3k8jZ13/ALuDbAW/
vFGqbu3aTHjBKuMTcw2CmNXB7QKiX1laONBF2ZX12pFBx16aeez5TiwuqyV+ZS/e
UmTMrSNdMYdLijAqwGsgrFAAEy0Ud4PvPYvQJovHuWPhhZv6xRRCTo6Kw68aMBTl
q1hu/zLGmMxY6A4SQnWZ4D800m/xCz8RKm3cCjMqkipihPq0eEF7DeJmD7JGdeCi
spM9wPyZJ8sSiO4LBwWxGDv5gINiWCsAWnmBfOxU8zSOACrLh2+x6qapIxX3r11g
nNmlwyzRq6zspnpDTSsgKc4fTOLLFRqpKi3yLVC9aNeyKk5W7X/pTj+JuCzAavGl
N6F7vB/axFDOrFMWL2dA+ZdTIPn1K0w8eCb6VzmTGjdzcnQAClmwhGPenm6+MapJ
YdrFyWQSgeLXr0aWvevwFWrSVAi7fhK9X1g0Fpqzs/881LL1J6IXzkumpvTm2Z2e
gTvGta+P9ayF0e0rcLQ1RcleudRnxBo9xugLxeM4rdAuh/vKKr0k+U65dEDGlWU9
Y+rjewlFR0RR3nCaK30IjcFKO0gjANNnESx29LQOLkgnaATKLjHve2Z7WvTqJgnE
4raOVpzdLYDd05XhGs5BYwPtcQOd2eBSFVVogi/009dDg9obLg2sQuAtr/vVPHrd
7ZG+YoKTZOCi3sWmUYKCniuiE4xiBphU8A97TBQp9Vjiu+TePe7IlQQUMJHBUiv+
aT5oa5JHqRRDtc3flzSzqjUid5+xio2q/K0s9BiPYJQhipVMC1pJJ+ibiSHLpVvv
ix3UnGj/puiZgv+EqvUMXtsxpMlV+S/I51fYTm7LTEgmTiFqEWiC9XsxN5jNWHT2
Mp1wUisB0q4IDtLKH/+FGUQY3blUScCZ5YqLymOUYquqVU18ZSzNU0C7M2KBIjqr
tfON7SsXojHZ6AkR/jK/bVmmXVB2HnXIp+UEnJMsZAnuEXn7gCHEeHdQUmArriaa
YJYWnFjZwDq80EAWPMAiTTmet6pTNkW5EWF3JUJvkqeBLGt2dKTZXNTBpJDw+d0U
bxHMlvpNi71TP5Up50/8gtk7ME+3v85aLKj5ag0ob90IxoX3zLMJ2IuApk/VG2R7
//jHnF6MIXwGAI+CIYPlHQKk1ZzB41pcMtyayPU4u7l1M7ADahBun5rPxR70E17W
1XfTHPxRilrcCV6KQ8JeT22xpUg9ooLovn5wqCM3+1YR2cV3sJGM6+bO6EIdWJlb
9huzwzNrzPmbK6EZdMB8+Oh0PpjwBhTPLQCw2qz35IJZq34qWV/ntc637vnBwqix
YESRx611y1k6z77zlLN5QiTiV4hkIyAe7372FRehpbpFottEv1rElkbLyJDqeW8d
tOTHAH79WTrP2pbIc0ML34vqXGVCEwzbSQk0k4toFif2FYf6EUzxzztv+j/9T28i
agQNB420fQ5Q5j2BhCoQBluTCDMP+hTSmtmHVKct6hnILkMzREPWEqgRl/upPT8V
riRgOuKA+PbJSnu03q7qrcoyrkDYzuk1QlcJtjsbd6q36SXvMUGTYS2dtyVx3UQj
p3H035Sz1vtUdCaTHrok1FX6F071H9t3BvERvjf/Lkf5+AA3NJMVuOuD2HvnvmeT
pTMub7l4JNIuR//oCeeoJdDAVnaIRVq2BtBDW2Sv6qOWz+xTZBct36xK1Cw4kzan
7efUAYuLg18X5ok60yL+jRN+JTjfJ16rehdde260X5rndLKH6haGk7fyrNUXPjLR
QwZ9iVHC299TUcAeP7nc09OfXPoxUQhDJUujTTyzqAOCb9JSx5y80PMrPpLKJCU1
wrCXh1C4rqRS3WxWVXFiPS8Ub8mCTgsWyHKlnYWMHAHwkV7M2Aafbb+ITNckavn4
Ok58WpSyUrjGHGz+Z8jfbIDfCmm9rbvrB2LGgZ8IKNQsDOXzbq9MvVN1w54nc4kn
PlFhQ9AzYmthh1l6wRUT2jN84gOgwUa1mZMaimpRVeEZVmHmOF25C5jZctBZcdc2
K4J3S3u6qLIfJRyUXy86t3CddXviAA6rATxfuXlX1nS2ChKJE6dBu2+f5rQ5fsf7
21XX8dyVPm5ZQXTagZQzPaGb6q3zSNqgchgZ4aS9HtApoAaHB6cx7MY9HCAxFnHd
p79+zS5QO5P+B8GagdTDNOGIaP3rtNQ5uvWQBrOitihkFxXPLoXAMPf9vIj7zjMo
AFCrlFA8Y+k+E3Ko+H1f/Vgs3IYMKsqbEGdfDb7ad6iK/Y+uBsedkFPlx9xnZoHd
GvjCwGM/lgi6YJySzNIH8HCnxcn6YBwqxlwea/dqBW0pQ/Z9yrzinGAopcns02/G
21w2nHWN8cIWx02JhvCSD2WwmhtamEYC4GJb2M6TsN7aI27p024xvCydm3xS88h3
UMbnbsZ6+wVxJaOs2QhFpfAal/pglSd8xY2Ty08ZHb/QSax3hMNO8xMl7pnHY4QW
qx+nN5oxEu3s1JRD08rsdT7pUahK2hlLkp907PUxY9ZY3P98155vCwHf7bO8bBCb
V3ppWsuV/cgPN1E2PvBijt/ZpO8mZCz/+Tn8GQwveOJgd5JHZ7/spLo3ukRtM15O
Wl3wXhATtIuXOAAB+ztPzXV3yWYOgX2sSNzP/OIisIRwOnzC2euiSNiLcqoha+5T
L/zpxd6q69IwF+CJJMNFUAQJMJUj2ik4FTMRyXPje5Vbb3RK1rmsDr1fnqXW3pNq
P4C2T3oEd7LiwEoJrtPctJgDSGmwwRbDqUk+R6cR/z4JX9ZYMrRLn2Oe+6rw5h5T
2ryqa1DYT/+hUkfHE22XT+fJDBcxnQrCF7eECWhzUwHbu63RT7Y9VD1IDudbtTkS
ffjbJw+fVyZIWKlhtDVSpVDuaTPJDEqYUGJBHSRC3ouRCKvdEjixE6tboZz7vBrM
GJRGmE72idFMK0whQtF56gj7iSGePRkhtM4cAPPOwokoJvrSyZ4xhomstJ6RiZ+y
v96kIYPDYwRe+BPXrt4anSXe87BA+Wx1BSFtCg7nNSp6FfwNVlTwjPpdOgAfnoti
fwUyhelULTeuKsGpH4d+B9mYl5dRiz8ghYP69kFIEYI9bMcNmN1FCsrbZ37q75hh
YZqg7m78IWUeSd43+FHqyn51w17gMkHAU2gr0UNDJ4qQvtvI000wX3f13jfdI6RL
r8NIdVOread3ET1su7ZgONhrNfzcg8Us+4yRfvs9A2G69hu01sSZBy4nLYhXqCdX
cNXMXyLN+j7aFnxOTNPk4r2G+kZnDr9ZQ0SGVKkwe4UfGzbXlGtAscYRoWMAEjEH
J2LtbeLC15mWnuGv9VaDRgNHD91r8fvipXWZiPPz1ofeARASyxizRehw71LilnQN
QhHxGFK22d66nJQkX4JCE66HMggLTPKu53oA3AVkIdHAbUoxlnb1onfEmFXrykEe
Uron4/pH6bcKUZR3w/OipGVQTbba/2IPOx1HmSzqUOBOs6UqKQZlJToKfo5YPM+u
W59oUrcR+n1ywS7mDl+/0CqlJfYGQbkFWA3N78XjAGVACyOkgYCj2thQfjt3+6IN
L/fgABiG9SlUZWKOxlM3+iLZjrS87OyeNHSuSVXp9VIowWW1MxkljHVJ1Ow0HVjh
SGHBsoMCg9ziCMLMxxmKU3yBngnMPVKNxFilmVfVYDTi4rWIkWsb25cAGwY7rUtU
VfqbUfDvCSKYF0yk8RpZDaAP7OyPWXO+rpiJhcU7FVhypMunjjCJd5pA74Qjy217
e3E7tjRwpUNPVuP5TukD6Q7DAqhYkg6HcX8Xqj1eO3UlYJuzmfCqPCIHk75krptI
/tcT6r0tHO81KGBF1e6yBpB24pCK2lce7ntHnL39bQQkVylUx9bzV9h3w91JmBCH
gcboSRsdqKtTn8lXyPJCzg7ujtNZBmwbbQhQ2cy4j0Pvk758/RMockzFc1pK3lxk
1gQGKP9pjwiIpm7oVGIoNawLHVKTaDjBOed0ogv+jIP85ZXR7I6qCbzVAQjNF3Pe
ZtlIHaY4gpAmpMGSbJLaT0RnEU73eo3T2q2ICjgyN9I=
`protect end_protected