`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 33072 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
EmxAgecO7UDIr+OXKjjkXP+mPSWtHmjpj3yI8v8lqoXK4uJZwQU2Sr42O6vd1h2b
FBTF3rDQzqVRHcBd4vGax8V2AxH5ic88P13Zgkg7O+8XAHhW7KFoVpcB0ErZkL1D
F1tmaJRvNxCrIuQ/JdRhb1uQ61otYHfXKoXCcP9Q8VVwIzt8/mYNpC16CuLtCVUQ
F3HUOXsVrdT1fAdIR5lqVKW3mOkcBqFftczwSquDzERkEHhCPHNz4DotMC6ApnSp
KTtjNEnJbKpo0zDxbwOUTJDE3YCTsEr1/ZGsfCpGHElppor/Wg84pTorXq6rJvqL
66B+1epbjkiDG2KdVSgDRtSummuJ/FX7aQRlEWpQv686thObR51bTk/tJPnPuOZH
0R5T3CTTBJuMQ6Wvwb3a06s+ArRgmiX7eSQWBOw2EyT5SaEbSuARwee/5hcSaTwj
/Wzdga7kLN3LAabUmdMvlrLAKCmMau1pHD0sm+2DXUv4/QpJRTF32jwzEF+p0veK
RqSnzl1tNhjwXfGehn4I3Xczou8wAi1OqEeRVFYqu+fQa45i1bTfM2kGPFIyT2ZV
eP4jl1z+CtTaUTSP92ek5wyXoz0KpGL85mmEiAKfpaqXksd/InXWfny96oBUGrYV
H86xT8xJvdvpXthNSdDIge6haDtkpHWkAf1ZQHw/RW69xBeW6IC8k4L8CWdw7Fct
EsKt56gtzzV8J7bu/GC+fkM73BHR+aG7tksh20ShzldO6mjTw91BE76ofw7QzCmW
l89DJs4micBYWpooLc35bTBPNFLnkjOUcruQkhemmxpIrRG96E398Dn2mmrxW3oL
ydzNtwkqu0DcCFGxhuQVLxtVLIaJec6bn4lkk4+suCJmMURVrVlMDlSa2TTX3Iya
4zNqTIwSRmexHtF9MN2RpSMYBC97wXq5efTVVSjl3SRj8QccSsafEsC0HbkcemrR
R/iM5rxg/Lf6b9pBFVReHdsmaEgd0prjvy71sbIRi6xCoFBK3nHdyxVAxoRHigcA
UhnQPe4VShXHQbkhLu438jZOvtGSHvUUJBlG7EZ5SrCcFCSQGfuDK1CHfN+o1NDt
o+P099irs0WZQMJzjF29gcRcqeu1rltgcsJJUOQpsPpGu9/cpEIofoL6xgkqCS5U
suo6JYkBB4k/1vSoMJ3mP1jN1I+3h9e/S4wEyLOLh96C5CznvM/v115vYW/yoUFf
kFfapFQD1yFmzFDevHyW96XMENWg60T+ITZEfzfleSlJZZShRowILftNyznOiYMk
YBunZVMwtkWEqcqu4P8ZDmCLsttQwfrHPaJP0LHhP2+qScuNNgNFwgtc1QaVue7/
ocrVlHUwbBYqTBq7ca9isnLWlBx0N8OQA3HScBAbYLt12u7+Q971CaVOP53ydWTm
7orjOxrpj0S0M7wJK0dxEHjSQ5p0pulRfRXTzkIWA6jR204288MkS/VpBGXSRMNR
lwo3fpRWEgiCx+jjV6A4sKKlyyGzQXfVo/KWZQLDDZSKDoXfBRBQin81utlltAkv
cZTWpZNW8oZ9cMLhL6dGzJWEz56TicfELCvvjkACpxm7cfE1ibaX5dzHc6GhuipR
3LKQSYaC2aTHrFq/3pRRYEwDmayysvoZDxbJiLMPEDZTp2Hj47CU4U/JFW+Mlgxs
YyiTKIxDZ3NBlt4awmhBayocto6DLykCFTzyp7fPysFhV31IshQp76kECMCCMd07
hb+GoetbyfmBRN5CJM37YQt06XJ7JH7SFih+BZMJGLmmkl6qjg5lsux4ScYxWfXP
0xMhMI8ltezj8PXrKJxG4p3d1SdKf09qEOlBCZU2L6tTI3dGDPkh26+EcpGYi6dS
qRPgn8dnENXXhN0uiyhJHBEquu5gJpboT+9wb9pOj77TEnf1GrkWERLeGg7mrhbq
TWI+jgsQ9wvhTDLJdORobpFYefyj+/r2Rm8/HgOmROC8HUdiqDwzcDSil9T/Qvb4
ci+I2qvRbyxkdSWnRCk/4Oq0wVONyBZtvZ/Ub9SCr7TbT18Yz3WqzsgIN4NXOpYd
2rNZuv1RdYGo0zJTGccGuaiR/aEr+Ak1LjoyBzLdRHt2B0Zx1BzRZHjK9PoCVs0T
wt1vlw7lMnXDU15Oj5TJU9x+wN9Ag2w5SILr3gGiA9VbzCXqO+xNqVxTbarnbfsD
+4tCWhc9LY1rRAj3WPy7sRlkO9H5Kv2v4CGxclJfClnkLuHwBKoEK94TvMRjoJZY
kUT4bfTaOSwCH+tNvH9tVu6BGRO9a8dd5W1IIKEPjnSy3IqeFLSjOJ59XQAVId2y
pldBG0h25rneii5FPfdJYruFyrB6kIjF8GC9+xf9VGvOmeifwy3n5Ny6W4nJ/ide
9Lg2Rz1lO4afChrUFbAg2UiMG1jJ71shUgklUp3edAnIn5Db4cem72swKMHoRC32
dZwTzavNeETXsX47i5e/WWeVQEVf6ESPaNXgJwLg9+9PF/0qOoUXkidScoWzcIbm
pR3oDRiggjx9KAlM7tgeEiu1ngXNEL8887inFFKfSvdyjX3PbG8NMz52yC2zNHqr
ECzD5T0zH53LYk6p5cryVv21Vk9Ar1Kux4L+H5IsR40cJTMuaxCZMeFMjnHeT6EQ
rM70BLn5tpLugcnwd3BEzZAKrK+mf2y9IsHSzxHuo/gnquqJpEqSvzP9ZLg5y6QX
ICoYluJQW0wXU09no1ISt4kvX4/ShNm6PIGQTI0FvRZtaqQLmveSUluVrSaUS8Zv
a+zNQLhrGowSFvy50pr5CnyzZrMFrwSuI6wvCiswzZPziM7pEwi+B4Apw3OqKHr3
Yh9TT/0sZnUi/8du/E/FrOYQKnyePQHZrTF7upVXbEJMOcVN/riqFFGkijG3/Jns
zZ9LU5D54LO2cRJ8eTt8Q0Nn4w2gu1gjVAaSqGhrril8OZsZxyqIX/RH74UWMP6u
z7DOuByjFpIY/nVfnKBov7AfdsdLUQ2smap33RVPd9SG6tr+eyB2zVR4Hau096d5
hw2PDhArGEveZ+mMdjRoa02nBm3XvZjSCgiq/Vvtrbh1W/sZZQdYy7btwVL6qnF/
u0snyeXSsZ3He92yxSHVHNeBhaSw8SG1ZRAhZ7AHZTzedCcpi7GMBdOOudJ5sKRM
flV0cLO7xkrID/UJ7Dj+u8ciWvcfHq+uF2AgOnMANTapPU8lK1a2Vi9DWLKWNG99
tJ1zghsEGb5Fqz0KJsfAPSzEv2RmuAATP/jPdnV36dfqIBKd+dAgRFV5pB2BS4Nq
d1De22+Zl94hz1HPTVVwXiI3AOijWMWl966hD9Jb04fiZAjFu2HXzx1TCz1VbIcf
bAJX+I9tBtDQS5Ao3HDpeXgL8iQB8vtYS7wFNZ6xXBSA21SMiIzDBJGcDsIl8K/J
BMV0ZQnF1nMdCUv+8mLkaqavQatJWy1H9S0mR/IFp/QVOXQ/0pvhBCX9WUJr2Sm3
kQVRGeWvSEc2/WSE33bIW8bSaKyx+gu/mLkNCkT5ktrMTir4kgKfXnmWqSKFh1Tv
jf+0AI3JnfO8ANg2ERMzMLvzgnfieZovppaZrGK39ojTNbqB7p7EQUrZhwNcyrnJ
Srq0AZHSRY6044AQVqvIpETuvfnmJ3YvmEW7Pk4+vTmhFBcdzOzB53zcyipDNhEB
SGi3VAqavYim9YbBgQOT18Ai6wqm78zX2tF4VuFCJMiGgd6FaP43uzP1YwC5PE3Q
2R8QD3QPYAl+syQDTl+Ulf1pTPIXphA+DJxCJ97EK/LXSYsJAXaDkGIN69iMZR4J
gKgbaysNv2468FmD//A4x1LnJJL/yE7pUXT6fl24y5xVfZSry97OUGuxj5WoGqfC
V67lscp0dgcuhUwiBwvN5C86EIpno2PDwQF6bgtdm8xuq3XazzX5CMN+kaLT0rVn
ms+SEFNRyzuDnenNDwAqz492YphWTEaiNzV4lp7ct6cN5T13oYEXNYbpgITA7M8F
R9Yp/u/WTs75PD0Ogyy4jntlsCg3GXsNSt057CedzeLmxOe39VBGe+Q0sOXyLUUk
3N8hSaRFGNtbZWsLMWDHUWmfJ+IyqSazjbzgJfwb/0zyNJi49L38w3xxuI04fjOv
zkYWFA1jbcz9d2A0P2JKBzha0muLW6LnZfoZpv86EkmNdX39Q8OXMp/8H1u/nt3q
A56Jk4nUIe5jk6kvm7B4L0N0qavpl9/qJIFw5RL769Cp9oD4trwf1g/UJGz+liF5
Y66EF14Ven9oltldmGfKF/COlaoGExSbe/m8YR0mgmYbatz7sQgNuoAUwrYv5GcF
LJxUGFMBDIbqI4v06iJMZkdNxyyKIx4zCQQUU0p3rRdgPdRYknuXc4suQjWj8wIK
ZkD3LIA5m4z37W7d89NLkkw0KhjphThEhR4VS1e/8FNFbAAoQTrxN5Mu76/Ndw2h
CVOIV0gcpHH2wpLpxe0xxHx4OO7F/a+o01X+ExPEwT4ayvRnkqSpQi8vhZ4MqI4z
N63L5FuxZfwVLSLPB9QU8IiHCCjEITt6a0KqPUMBaF2fhC5XAhd/8oD4U2/WT3N6
rX8cJAfeSfAzDPDbcTHSMPYClPc0Kpx+xJD8Y2gA5QXdbnIO3SAATCBpOgfABjkm
k6EG2KWG1Q7bQsKU61+aCH6a/tthomswlNb3r4QerlMWgkNsXZwhxYG7vs/1PBCr
NFDKS3nzm1lw0RuDJkS+Atf69p1zq6csCR4pmjJp8h5wH3fKjmtgYuimHxIz2A/O
ZoiqBhdhmdmwwjyjQY8r/tDATAglug/Qic6ucRRqfMqyTPDyyJuNfGiVXBdPjZr3
8Zexai+P7PgzGvVUiv4pk/5WA2s34KM7LUtBhRPJ8+QZDDPqbUDXcMfm7NzSpWBl
FAeuH/d6PbSbBnFcwlBPzabBleTgI39S2Kw7lN6+fnyN2XA4VKvZ5T3Klot/cT86
wgjdSBg2yGB3W2Pm924j36kFUs6QjkpU1Y7bwCO/VURKcj7ViTZgwRD5ybUlPfQG
XlxI9OYAbxMVKyqgGXWdu1LuAEied/DlEO8IYSzsYpje8BDwW2Exhmm0ff5k+due
fMm3kHQ2+KBGu3qtMHrmr6xDosquuIsGdrUGTyuZFvvjFmM+DEOl07qTcNh0PvmP
yu66w/BAPv1HVbAgIb4Y7HK22PB5ew63ysG2O7Y31oy+H1G+cWk47ZXhYQ9bcm0b
gkQlqmA/7yCV/GiqVFSTXp2TOnZuAtMYhYohbbG/1L0xwDaMsXeMaE0i/o5LIflA
UQkQOo2NjZH11kbm+DP4Y0Nq9CF18hs822urvhlu1le+QJLHacIvOc3F1PqdP8/Q
79bNMt9lS/VdE1BRPO+9LnK2ceiRFX5JBi/2iEkJ277v+vahz09QCQOb/LTIIM0M
5pOX1pgvaUCNkmxc6R1zCKaAQr7AqF8WOz59fPPGMvO3X0rho5WLlIADLoNKsGde
wJvEmnLtE97Vx2FLbZjA973UW7Zdhm1nZYa6lBUrlJ4VNsfaK4WfVRSbcATIlsJn
faNAfxcl/PxJsMfqez23UdjRTZLCoSyVgt3IhVAImOLN515dCrNkx5PFtZVZi0rP
wC0YoLkZYk2w0MzWWrI1PajHZZUMKW49f26q0HyqFgl1gWBCSv/gAjavM8KJqVbw
PXr9+fTLPqZ2M7CXDhMKVWyr4OnI1RrVo3omd9MhkIvkVrbuQPv4nVR6EsxG+WGI
WeurJRgbd9mSELu//VNqjfcIu6D1DOvgkKUxw/Ul4Bm0hCvJgDGTSB71Xks/R4ih
HXFFMg881yqiwqvynZpdUHYpQJqfHGJKKDUI1WFJb3eQlMHxZuoPmnAMKnYQtukj
6XYfp5rpCk65Z4MRvZVPTvaLhFIj6cKjxfnsSRs5+2CJUKTP7zHgYI2jNS8hCbCW
YZgcZf4CrEsEj7dEfifMsNoWTIAu0MWSx3pNmiWWVyDhqcGq6wr5UASxAh/gVxB/
0rXY3eOKgnD4ONhkDYhzyFeBnSqeBUrA0nXU0r5LtKLfPCGf/VK1RKoeCiHV2I3I
ohcSMtHE0h4cO/ldSQq89cabe0/akrw88Ks4+e4GQaUBa/nrRC5/kGGfO231wXNE
bCzFA4D3sM2xqufFW1to6DCUCvbyhdQYKzK24Yf+C2ArxAegO2HtO7PNfGF+5Ixt
dlnstJJgE4EezT4LcFwvtLIF8y/jpSuRhjlk8HgnniU3eb05Penbz5XYGXBhEtY3
6NDsHU8vGWo7a8CdI8clriiUns6IySxtQ+ERjWh+tNo+EtjjUBupkFhmAwmlARCq
+mYgydh9s1erZDQIEPQ4d+n93JQNbSOpbh90tVlsR9JFJ68pUQmxz+5Xe1sJExei
4PTFBR0icc4KFPfW2CRRt0kX90fnpCObUy3EU0dWzzgbbwjm+/vZxvCvieFiE/EQ
EXftoPBYbAF9hfI4IjiuGDSP9ejPSL04LLn9yB0XqoSOCXdiXXhDfz8gL2WXltkC
rAEhPHYILGWHJfg+8ptO8o/rrMTUqoyklBAfKBc0ukEZSC3qohnVyi93mprCgRCr
TY349YFZJmeoyLt4SH3RD8VobhE8eUFj89ZP1dAO0IbG5fjfW/4AdkLoQNcQsvW5
k+BH4GR1OI5gr68hXfaa51tQo7vVLGKwpl2DSbl2hhZo+sS0JpBoKzKnXhO6805Q
ImQ/gAzhy5E88nefUrlEmxk+lr5ArLaSSdZA7GglCw/rotNaSNsM2G1UbJuUw6tK
IPb7YekQoeiZi1VL1asR2n6NIid0VcmI/xOcJNJ/0dJFJYOb87QHaGVIx0nIW4NG
zTOPyIOTA1WOrCTF/691c0ExvXbtcYVIPplZjhINOcaP5Nb4y2dWuCzyzoKV86Io
9JwwZ9fMPFHGRVlH4kYVbFUOl4WLRYpRl2dA5ZRcLm+Q8cR4SJckI/q7j/jYbOmq
mxg115XGkJVjYt+jRmeE7gtBtkME5RWJnccKavttoj7DRacqbMPLv4oKZOsaRWTJ
88aVHDXVqoTr6nfnjeW5sT9HOKlyanOsYusIm4VZxATEDAWbVp+0CUJqSN+QtFAi
nhtfRa0OZt1ZHWTueH5FJc0ogWb4o7sP3pRcoc852iJyZQ1NMHo6tfl/IyEG5lWQ
pImZCbkcSHF6u5HrCCIWzP1rrhccdnWBjwfI69G+W52NlxRuFU6xCPVHtNlheRer
8IFXVbv9gKSVbm0g1BIEkCNnsxm+FOy4BjyQACFddmad6WkIJug8SYv91ALuFrRu
dUoQiwwgV82zXmDjExddqaMAkEnmpgkznVrxCgJ10X8i+fmKu6S3WfW8cScXzkuE
9oJWrQlg/CEME+VsADTT0smUY70iUqXVEoVDs0IO1hltNzNdSceP5Dd1lkfC6nPG
5BrSs5rCYYAElFkx/fErI85pg573xb1mL1e1FD6Ovj9ICpimGLssX6yl2j9NQrhf
jbyTa7p3sNjtpaEQcpLpsSOmbcbOTuQuL/JppB1sDSvR9mkZ4T1QU0aByD0+pJ9z
4IGjOXL3qOfwY46siSLwt1V51TynMfjDzDIS9SuZfV2KYS6G/sZS7Had7+93Uo+Y
kOcw4o/IxylwQQ4QYA5KXPt/m8PnjcWebRZWwIeIlCXUg47LNTHv2p7pvxFYWVw8
2FgL2JghDSY2kyFuGK+JSXet/XxPcMVC8P8lVd58fwx1g5WZJfjxonLPdfwpM1ov
5suJldZ4Klmt3dBQLYxWnBqx5hT/Vu4L0pBJw40jjwfhKWrpPDLCznRAXUsTgtNQ
jihbUxB3v1zV3T9ko36oD5Yz1NdYweUAIMKbGAt7+oTeWmHG5F2OOni7oIXqB8sY
2G3tAinalQqNZAC3AOHLKumu1zFWkrrBVYoJ1SLf8ZxkdSii+gCTKq7OS6s2aqhG
rpGYyROVxm2ppFih2WpkPUhghYyoEZNBFsSxNkUv6heaEEeDXjo7AF1cdKVJh+zY
UmdpsFBHkXII0HLUXoYUs5V02bahlx18a7lEeeTq/Tqe42fU46PhKx7GI4w0cysE
dOqlZoedjTj3IrTraQA+THrXuAd0z80M4t9t6D81ldYEndDYSIUA5bY/xnhmKrDV
yfCxWX3v7yHlCpwsbun6m4pV8txcYakzxLWvu1kMY8bY6gHBZ8zvnQhoiiiOM1j6
3IrjAGVOKCBTC+ysYowWsgRBj85oSPNsoUTmu4D5E4TNHmrnTH/tWW79jbD5EZM3
X+/YYYVqcJ1pFbvOlmCxSe+jhFB6ehn6WhMBfGRvrzdWzIPqkayb/k1i6+ksz5MQ
B9iISafo5J3H2x4qdyQ0rgzLvpGcMqTDRQpGUZmDcqcUX/K6D5TAJuxCwNZ18M4j
mi0KsszYBAL7vDEO/sI/ECkReyKkBaX2YS5Ss4h1aynzdx1T0uulbVVGhkrvJunF
W7AV0CG38A5KoscqDE6WmSQra8Pj4ccroiwYR/A4m/pfT5BD4PEwBUEJ/E+lW3vS
eRfz+kBUAaFPfDdwEm4VrpbClu/gqiG8zzcLoHaS/KVG1hfTid0MRf+9p6VdfOO9
pasdl72+AK3elRsuU1c5CSwdnRKCuFuD6Q4wdEDDOsu0RQ++rXP2SpBU+2iVnuiu
9vuoFGZzKT9xDfJkq7vfLAvaA9MPBp5wo/MUyDfP1//5U4sk0v/ktpOxeD5CmDJW
EydlTkXVskLeLQwP8m6RlCZnGwAVUBtV0/WNOG+TgrEJfs+1lBLx7mHSLtwQTDX8
W89fYd0Vghrub2DquOXZnwplYPnF9pkrTs6pMi2vSc3gRnOXC8s1NMz4DzJUhJnf
MmkcSQeEauZ0WhHDlAJiV7hJPwZKndZbrQcElSislRA6eTjyszVZFzjtKI9uhZJx
N6UU3PucQ3UdCQVc/HVB6qb12OIl17cxW9Ru9GoHzkiEf/v1/Y6kXOqTq7bGgMKi
Aq0QrzfuJuorm7pCxG5nAP0TMctGLWbg+MK91mGMlvYA5j/8g/H96nTuIdsTP0H1
jHkl2MxJDs381Vf1rEJIpgGOWgciNL33SrktLSrbFrM6E5OYZZkQPA5WvHREPBlH
0ln5jqsT3HNACHvjtr6IpXb2EiXTMxqSa4u/fyBN40F8F/XCZiDppLN1SOPg7A5n
yzIssen1uKe2T4vLb9KzkTtZGKDCvOmr9++aMYA0EUG4wNzJ7hapvO2JGdpYcdsS
d0KdmXbhmE+Ix8OeUovFITqMQ2kMh0RKCAaCLrcV8s5x0EVV6mjtc+DsrGWKj3N7
KaW6qLHbK549Ja1L+apbuMLcHbwgoRl8EKJqYdWalp9+VRomN/O7YRKWyRXSvu+x
ciYIHFxlK7YEeJ5y3WGYZWGbIDoR8PEAjKi7raUFUaVyzdqf6jecB69QG3YnlWk0
l7rgCBxGgoHjstqF4ORA5wUiMMC/J/lm6Sn0UmQEvcF3N7i1Fh0v3SAuvjas3Qi8
1cd80ux6Tj9/vmOB2MEodT0lZ4FN8ggEItvnt5rUP9Sk61iHcj8Z37kpP1trtlDQ
kn+jB6IaeJy0ii3rdjLBtBd/7RjfAczSyueNbuglsZ29i5DUu5bDP0GTXEJ7Dwff
iOCoKLCg3OMR2B2M7U/KzWNjIOivug6IjGgHEXRIjVAdnAXcwBMubD/HBSlhIV3v
mWeYWrjGx5RGHp5rsAU0VsfaLdl5jewTFE9e2Acn/OM8g33LrzpURdmMs1lNvgG3
6KVRreGXwzmfPDGj6nbvra/cofB5AB19VkuGpcuFO8xT9m2x0yVgGhg7TCBmoQyp
E3hUzmodZPNgeBQmKkD4Z9uYUOhT1SS6DcaIADUY3vinWoxj6FO3mDba7BE1byQx
/wunw3tm5V1abATS2+EkcKlwMKj5TAlM7WQlapwYM1l1gGhL0DXpCLs2Cq58F5cm
YCiQrbOpEqthxV7aq5OBjcvajejGVUOw8w+4tIXeS1VXqeYkWDn7j+grEa+X7/o4
V5ce/Y/fnG1Yb4o3L5eMv94GWdduh3acZbfHG8Z/YTUq7A+XUvjTyt3TPyjWAK4W
kkPtOj2sq8pPq0iw+IczUMxTHIVj9rI2tW9iSqG9/sAvfCL5zdyTeq9t6laV5+n+
hPGkECkm96tivRs4V4Rv4cBcOanZJerKD5vlZMSYjGtTNoOKn1II1qVw5ojJalSo
TtFhp7ha1h82nqbYfeVSZ3aBd4esRArOH1l/p/uW0e4/W1Q8t00Q2n2YoQXfLRxm
vVYIcf9p2R42W65yf7I6BrI/qLGiE4c9jfLWzGC2pbvJ1XuJtwMOxMmJBfnZ+KYe
NjhU98DALjP4PQKjDKnvsQpY+wRHXUAZAhYQmJTAZd9YT1WVNnJMpQtiLsRq6u8V
+STZoLUyVDylrUYSElQDClPwRnG44Fokhh3aXPZEXdeyS+EuNoYXYTnnMW3FrB7H
AvtrfvGmO+RQF51QBVLsTEU9a4VobALTtA95KG5Ee9I5BXUpLNbKcb+S0Ol/ONru
xtqS+6TGLjShMvPQV40gsw39JE+SFN32BqrjECtfye6qA/4vEPVVKRh3qCIvee5U
nA0EO/Lo1OE/0XTNg4kz2rG7ZlOUcpzCwr+9fdR4qJZlIdOnUasb5Dr6fmfGXw6l
86Q0trXEN6mlS9LmNKhxNTK7YVgNwLcbz6FvNue5cZZDY7d2icGAeEvMLDldQIQ0
y3gK1u8GaMCbz2NFl+waEURL/xvcjQHdOxIan1qBuGl+yA+E35bq+1EzjNesZCa/
MgHPip2oT83iJgZAKyYmhrpw8ZbFMlyp3DkDusuhukP8Oc7Pw1Gj0MlSX31VUH5/
BTjFLrrev/eqhjdEaGn/7khlKM3m7R6G/i+PKL3KWOJdngyewzlGvuRVZ7MzyQal
cLtCNArEdXDcH3Vmo2/xksZpPd+F0Nap8rVGeBF5rL3foANc4i1lvLsmcovY3BUK
9AVxyvwZ6QcHDkGLwSLgqKS6uom7IygGP3MRgcyL3dzpRO814SpHJt6a+eguDrEH
mh2c7SNfszIcegZD8VfuGMT0FQD1vGq9kpSJsn4i/6YU8bc2HALBLuDGBaoWGaut
WWpjb2bLx1lx2TgOLM0wAlDJGoLsO+AMCaYB4cfh+0/C/LpaNzwcnlfbVFX7oz17
akJySUqvTdoiPZwRZ/RGbVR1pl4WqtYTF71YrqICbQPqGeaof4NXucgTcYMdnf7j
oq2wWMOpowH+Yhv7uaXEY1bUoR0bFihIkB9pBJYfsmLr/nv5tO3BOrMXTj3ezfSo
IyevzrIjpPTuPzKVPOTJaVUrZVtGd6X+aSNUVeq7W/LHV6Zf111i/x8KEbp3rbS1
tJb4pEjDrZ8pWrlEsWIWHkBspoN7Q9cMiFEC0uodizgZfQ9Awq7kvMebx+uo1jQQ
VIFxBnNNXXTDt4joNfeSia+EOViSEzofKhONgEwPskTp71DIwBSfLJzJHJohhpjQ
Aor/CiRO4AlX/cMYarz9l/mEPxZ2Annqk3bAxVshINYhcdis0IPhgrOnvmWK/sUI
NUs+ftFsG/xDDVLlIRx5lwJNHIUn5veU9dEyXOrAnRddqe6WDs4euD1HF3CINg2c
cCsNDsJrUmv4SuWAZSBL6ptNPQX/bjE4cyEGQNrmwh8D5S5OcQXzvx/jqz8JRjJJ
Hw0QuNzAZj4nYju0TiPpTUggfLxZGlFmdh1Dx/uVkQ+whAp3dNc6XLdjBscN94Ph
rKB80ED+C1znT4HW7dEJR/wAxTyQfnQgzy1SQG/5dT2mXiXfRElxqrDMMWmB4bq9
KVSXfm0YMxmB7f+d/sB9rRVTrRMRcn2eVXwtvV7UccvOzmoMzGGyfsD+52j78UUt
zwpfCK4QM5nJZuF6WN2TMNxsYadoqD6yC12XxaKlVPKJf6jCZOdMA41Frsaik89a
LTR9ZFvBkAOWWRgVM1pmMjBaO2Goq+m1tOOdK3tEI2rfTFHd90G3Yr4BpGZenj5V
ezLCtjgVdS1LzSVzO5xxiMq4mp5X7hZ1cjQZeLBv46jUykXuSaYswunh52UTqd5G
6UgDjZ2wtyLLTt4Gai5mR8WEsh8HFRlyfJgT8gGpkRLnTwFQRGn5n/poDes5n8EX
/Ek2RY5VPSz8IXQdqegtAyBZCJakWAOooNtTjgGlawX74FBk0K4WlRFNo8C3iBaV
tdOBLkJCQ9vW5adJUany3lyy5kxUHoTeE4X/sQMmSXu3JD12p7Dab73LyWOSxeHY
7MbK9Sjbn26QhSYPv8B8utBckYhZfjXg0vBG0T9VS+3uLJszxeq4i9cw1AavQmH4
dPPQ+2N4atYKUczRJLFUmfXrjiR9S6Lwsg8ASsRtzX53Tzmw7XxAjp8dExuAJFjE
CjzeLeIp6fbEfu0xTMqDWlHwtN/XDKnbMtBPn/WMKFUtMsnhhHvSSm/O24QkVNDk
2PqMkYaO+XldCZkeWf0470pNzTcp4wu8aahxn6GTaLxxAQIdz08pyoR8RDd0S9Rt
+/C8YoXfFtIm+enZL4yfsnL0HIuL5kgRkTnFUPBznLE7pbkItFyqaIKLSxIjM6AE
aADNAarHNbrUvchDWtxrdw5GLRYpjzguMAbyWCpE9oFUsCuiG9+bNou2HSopQDCb
3lUZxhN1EjTkC6tPJ3NpLAwiB76w3HIexiUugwfxtJDv1WZy/wHd6lYVAdj2eQGR
6Kzq7+L45XHgR7EwehBb9xZGfqXEGLeXpZ87Xyd9MhNEwcNpSN7dOoTiTiiCF2gt
xXQdD+5bUMJW3JAEoleJMbq8Zf20Q/PmFp3UQ403Z71b16FrABDvRQYnUdC0peBB
tX5HDQGZ0y9ZwvHA/8DGWe+GwC7o8q1Ps7J+nn/yYWEcYKFPX1X3YFBg3PTPjcyb
eSr3g41xH4yAaGi0jyeeBDwMvPYIAkNdJx6pfzTp/PabWzO7uztgtzFEt7Sb+Z8Q
vl9Xv+mNUQRYNzr55PUqH8Q9BzBVp8OcPHdP0eWxzaBJHi5idB00fb73WsHHjnyt
aERpMXqW7vTxibVMmbAi85KVhm2/5dmXTimjwAp9jhC9U7h/tHpiO4I8KmQyk09A
aoa4dnP2rEJt5J0e2Go/O3pntrRL2FrERPEHDmbBCNhsUgBPk2NQgztT+ps+ax7L
kZWFiNutF+ZNKa53piz6Ngi9M8JOOowP7DN+KOwx6Hsw9bWKzviHFHET0IpIYgHp
la9zSRMph8gk5i8TisGGS1xt3fTdFzIa+l9y3JAhdxTPbYUwBI647TBCCMMNRvlp
tEB/IHo4+4ZvAfG7CnYhoEqcrZypVib7p8K8B7Yw9K9NqpqhIJT0bb8YJLOanhZi
/Iq7ADL/olGi/8byTUwglj5ViDEqmx4MK9+wQPz8vj6EOBCqWiiX5MR1bKF/A9bw
dpx/Py1DlQQ67v7V6hvwzJ5laYIvIrutqxD1jdI+IWp2al3H5GSONhFxKTDSbNDt
LszbWTNUMBthOu5DJHLBCbMGFcHRM0hZL2OmafN7AAn+cNjWLasDWiY0NALsvzoH
BczASPCJdJaqgvij8tdQLJID3DfTgVuRUc23ZnWV33Eo9owsBU3Vzuh00arAT6kp
n/HpGXvV6DfalYkuzweVVRExs7dtER/A476rdNJirMsAANHI2ookW95dFdJoj+Nn
579CCDt6OHd9atUM0+fGpogdaL6+wy8+rF+9Fm0xccv9UhDu2s0Ajc+YpURuwrvx
CxGwQYNQ65Srr61FLgbqke2TEcVmSh6KaDAGXDvvojA3IkN82wNowJVQ/3A9sn/o
sjQ1hGjXKn29x2ByVB8DoNvDaiQ4tPGwFJ4fzjVClmgV2IH3RiXphYLDy3oBj4KR
yIjUIS4W5RK5OhOgE+wpsc+AGPhvdKCq2DGg+Q8QO38GNOPZvIZI1bX/yO0PG/cc
w775zvSUdVeA/EkxGKKs5hVJOtl40BYe6STnUd8i7lUqQYRbXR/4gEdXPQCH/Ncb
UokOaS2Ldpaan/dj1BYuNzhQ6qRH+MMKrZT+2/NdjA22EQwZ5JOdLGrNBHxy0ez+
OfIAImJPJrrcs3DMHrvOGhJ51859ETpFOp9CojfDp9Fvm4lEeB3E5DA/ZD4g/cDN
fmHYKTLWtkOGG2AK/faWL+1zqf5/gYO1tZpCtEUjOXdI1YIxx3tMrT0GVk4NePKn
sWmVcMYqZ2hF27VTxU2ntvsyOgMqys/YI6DZTsF4GN+n8UtEaw9mDYtsKdodUU0g
egnnvzp4Lt7TObm9Hr1+FT1X3XU21Arj6+wzCtJq6RtB/kGjw3pbzjZkpCJJM2ka
tmFRi4afDX6uRT1h23tezzx/hQJgtXp1cl6vxMlQlI6/LFFTmC7zyMRa+oZOz7ac
+zAxoP6gqbYD4PfgGFxytT5tCKV0umcJSKFVtSBSAyRVg7KOEb3KfuTUdfGYmefu
S2COmJIzAKa76BMPHAiKh9BQk7jSVn+VXI8Fs9TBLRyJvbu+aPgCME3X55Mty+v7
O68yLDCWcrZlTAY/jpn+QrPxOqeTiL51cJpGtLaDp39NI2LbJR5NFGnTjKIe3SGv
MTQ+8k2ImXBrY0LHupvuQR6CcChm4G5/jdkRBfGScibg5qX/9NUyEem4E+cieAJ3
Kssj26lXsq1oFWVgr+FIyGDxB/lMregP9d1LaXF2lvOdIILBjiPVKwjqYqh6JX0T
hY7zuFjcmohgILQkZOSkCMxIj4kvddJLjUyoh5gTpa+g58k6ltPzfCDcjbJsJpCo
KGsNsfYrJ8CFPGluHf473k3dnL9LQF6ZjvtBPU88EyD3i5DKopeHqAESe/S47jov
0DvXEzmnQ8r7fEZ7LoDKw0jUsLmlHRJtFUxn3bIzNyz4QhlPza/0S/gBNLUbBz/u
02EMGecfonOVMUhqpddATVT66BB3O48viXwqZEbJxU8XCg+5T3nHhKu/WftQjem1
wVd06UjEyXcL12vex3M0w6i6P9ZZN+Ylo5NuJJ36gjtBlYT0epuX1VG9F0PN90Ss
x367N2H96Ud8WZFj5vBL2WUDpUboyvx+MdQR5pEwh908trPTSaQ3BT8EhiVNcuSR
IObGjJkJHOofEG8oxeuNxVdoN6dAAv8XP37GSe83ZZABczWwVUhhrbzXS4kEOV6W
zuCRYJz18k69DMXO0UpsKEka1KFGGiiKTkbLnaj7iT6Se6XLGWV36Nl6x6CyKhIz
gWhmGkUKESET0RRhIuUNOpn/hVdEaZythn8GFStaDZ2u4m3K4X9qm7Ftmk+uKG3E
F0Vrb2WqeihsMe/ZQmqmXOoTi7BNYQ9tZYQhlbTsLIpPnrigZsXJEn6xGGilsHBY
HOTbnSbyxOZtNhGJ6EfQs9VsCbxkqX6LI+j/6SiPEvE89Md/SlbfrLHVK8ml0fj7
QwZNxxLv4pisyPkzz13aetSRneux1+hB8EXqEpxosAFpGcvcBl3kMNxZBv1smHFo
rDhCaMQpZ40XIV7pwgznk46G9n3sN5kMK45oix2neJodeZDJ9Par1cmlVfb+JBr+
hfRQDd3iwCrA9oX2AehZaLOMYf6JZ75LOhbTRfhisvmzj4AJBaTXZ0iD1fFSO4Lr
53riXlcRIGGXGdWghXEB/txWeummc/MD6odtbIC6kByVFF2qe0GPauBF4Ii5FSyE
1v1qUjhoTKnz8+aGOGdusrUM2x9VqWINpf5EijpTNpoIXi7njRLzY/Hxv2isDnRA
IWi6yQLmx/G6Wh5CaQ6wQbKUku1p+Z/4fDsemtkPmxyVbDYbCe25MWoyThu5QEZJ
LXL4PcKIhSIW0DZvgvw5YoxQ8hYVMseJANidARBcj4N++6xAx3eIqBUn7l37m09c
0rfOCLxofvKwCeh+rgCb3Fn13VZUHWUfBBIQFRpOVUKDPrq3ilcS+WZ7nZpxPl9/
KFySA3/tnkv5DvlKyIkdDAmZkzNJ8aOF3lc3jatwRuRWJBjDliAz+XS/dbCFUULY
vsQkHtT2lysdJrh3ezhXYSPEsmpn5N4YzoA3MCovuJOnZYO00YUElCUIf38Rq6YD
aRICavaSPKj8NiDAjg1QeY2lNHudm279o1VKxNrOak72LsOXXIvGQHXG290h1PSy
gd6vCBm9S/1BSMFyAlxCwQD/eQDpgI1LslOHwo5df0FeX5ovTVcBcNlrQ1NK6k5c
JQekuGl+CMiW9QpaqMqgrgCuGKd/l7xpYuo+unBWTBQhREJTpMsCt6+elBKM3s1t
iDYKY+6jZiis84r7gDwlE930EzvEwcNg/ZVewBCi9I/baZsRYBwRTISD65WQr0oS
DBey2YIOwuiAbCMjtiBTbB3WXVUOnzEu306FoucuPOUXfQe0YK4KOtyNy3KpWwH7
63bU3MjC2VJyqaqRWcePweM6ztI3bL2EiL+QkD55ZRDodrgg4UBurmgXcr+bu5g/
FuLzb/1U0dRv2xUNnAACl12acPhXESbienlTXp8+t61pUMqUhCMCOdCJ88fcgAhi
b4F26nrJdweqmkM+5LxGy2C0KORW4iU1gMWiqxDl6WoSjFkMMZTl/4Jo4U7BSrFM
AOTPXsmJEsD2T6QQCO1Ruhnl/eeB1/eG56sslZ+tdJeYxOif5wb1DnBwOcP7d5a4
eogXENtjMbqfqAW2VukuQW7o9EsYWWewR15O94MyBZVwLFK4Lz8/F9mlPDZm1YxR
QPBHlU2ibke2R30jrw5/qHffMh8dUcWs0KNyezV7gkHNLuEwuDu3IXJwbH5GpBps
4sl4+8oTUPP4tjwtYaDbu6e0hAxitx85uUe1wb59kuuvJsem59SlpMBDuWTO+/2k
hTBVtH3t16zzthUHzpLwz75fcnGLxdkcu6277B6lEcKVx6aEFa6+FBShI3vBcaUx
9VrgSOQAiWeteOrsAO/sh7c3oCDL50779rLCaRK/pRLoRaCa84n8Ii54dPTnELz/
C7DHMunPkNoDwzRMwETHRjx5VhumpjugnSb7WwbncaWsohOj+VzjMwKqkBO3QJDC
CWmz87uLHLvafGuWXqpTlxsocY/JMurp7XOHG+i+1y7jENHWDsrkKIC5D78DYX+7
RO0S+aVdtRvUYPUcLAbDw88rC8vjlnm+0drkbRfi8CZ/DujGNqG8/1cE7aOyj44p
b0TqwmMvpTug3OcoVZMbTkAslfgcwrR+mdZ0/HTwb9hWArzfkljPiKyypAS7pIcy
NEc6g8Widjc/unTZpZHfKjzcKsfGUCyvB70W65naSqpGnjHx+q4WcVOuLpwxDaTl
nTumOhOpPw50BPI/678QEbWeDqnP1hiUVk9tso/fcEnf5TgOscZVzvNuZLO8wbUm
PPpMhV9m22XWyQm6XTcK3yLQMhZVcdNmnyLA0JuASiXzaGtX4TUbDsKUomc6sU/K
Pn4+wVUU4AVC0H3ip8dLrTJKKgrLoQmiasKsnd7/ahIQA1QhRLtKnvNduIBUwtDg
7deYFYbH8LjsLjwzioXoyJCBCJsWRFmcmWjoiwNtYD7pG435q7nOTe8Erm8FfduP
7gIjK6hX7yZzLjxjqnVi9YZgFL8ynvaAY6BDo6H4B2OnXn6x2n1OYs/QTUrgEjtQ
+31wWVcXev4zCPdoGhx6meDZ+3GGJ9tEr/N/blimxzC4Mq7lqgSCYJXq9tOVzas8
TgYHaNzEXt7pd9q6pU15VhMUgekR/sc9p+JMe7oSnRMNH2yI/2BL5OqMQ4w6bSUQ
lmW5USkkQZU6jsEukAobp/V6YEkX91erSXIc1wSK+mHmRJjtDRGjlyiL/n04Kcye
TthigTCmQVb3cnyZ3l54uMAE18GZ7tc21E/CfpX9uWrxDVzYvi1bVG14sAPmF6xd
feioLW90zpOqRLvWC5IxGA9ukOAPoZMZfQzSGOTt65qvaxhGfxApidSlQmGyMQJx
3Do28dyg9/J+VM/jVKyUeZNtzEjRanyOwGGSWptAAYCdnSVl2bqTWfU07Uv9JBPc
doT9krm1GXIN7P+NBFbboFab49TAzegTD2wfaaGFCjN/44PRtp/UZkx5KYKB5l0f
x2c4ozWgfxV+xIHiLzQtX2TWRR4ExjwUAFmTKfyjtj1Qtd2NtoY4n8T4uKd3htBi
3QC1S23OrVaQk6E+9cW9LcLzK1SkpcrOnEGgKsiIM/86YkwAMqI8Aje1ef3BHwhj
617qucfUwgomS1xK0vWwP/dQ/SAGa41lcc+KdjgDKqpHcIFiJxQu4kA+d4g2/md3
oE8M6hKXki4TF70WEOWQwddpZi6Cxt07Tb7N6oUNRrlEcaIN4arYmLR09YYg81YY
YMjMT7gcZRp0nkb8v+ZRfNSSRxgAXkQXT6Y4HPTU0UvseXjBjI36KUhdqfqEMVK/
I78FBpNaKzwPN+9v1qEJ18ZwHl1jOFy3nv8iqTY1CsHuvAczpp155lQMz7Pz3mkG
cI7VDppNUbWMfu8OVxqwh80bcUijpuqpfoe100os+YsQZNoRrnT3RShBWUAHjI23
zQa+5YR04q3lzOHkKhcucFPqQfbXSEDOZe7uVMRnkyg78nVI6PxuOt33Ull1gSHK
4y3lvNovXkkLZbr7AmjyysPh40kAzX52MW0sogjOAYb5DPaoFjqe3Cl6g2wOAG1i
NvGbFUDBKrQ1euteBu0o3POCoWKy8S5mTf5Cv3f8bfHGmHPgZnfKpb67IQ+hBoSl
88Z6lPXgeBFMu0vc7UmoN8VFadAxp/s93tyAt7WmMZpOf3YizSiWQT7Z9FnQpg65
d1IQPehS9ys0zBkL8YnJ1hyz459VhtYw/Ob+9GtzGDPYnvpZQnfvijuQOWg714dn
b9ozPVndHePTR3JZ9xXFej619GX9QnEkwBkYt+LWPHLadBNeBhDtnpRDrBF6fGfu
hIyL7+1zKxtvAssj3qk7lZ/3HvGcSZVD1eTUmK+zQtrBR6jNIAzGy12KbuT1F30N
nHNZON+whZI9c87LYpozTLqomOpR9xMXnsxn/yGRATydDlqmlLFiriSioA0wslEb
0hQl3z0NmoWB0ujHcryp94gSWEUkrLAnYpnJIDpgQ4tjSP7RKEWgIBgIetAxBiou
bhbk6CCGjU+IEvhzM2lG08/ZX7v4P3xuoTpOLpVWLV/ad631HX751QMueEPSKODH
x9X2AqaGMx/0VfEczyw93BgQ2qEXJgGsusIgxVFBCmVQhMcKj16DyGUFwkGKwFU9
bD9ps70v95wvPjWcgQep6WBUthP1dC2iTEv0j6xTn1LWCyyTsZl7x/yZCeGJ3u4C
8p18vL8iZr7Cb1zEv2LMni7H3+7eIzpQJqPoa7vsgFoExFSVKZGw2T0T6iqrhIhb
ybXbwKsoihDDtqN2rwn54Q3SOo8Ebjqua6LiVvCboPzo50mfeSTj2mMFQaRtTo7L
5l9IHQjJX5V4fJ2Ly5wmdNw0qyp2VWsm9lXxklAYhUyMiDiOoj9rZ2c5q57CSD1x
q/Ifl+bGEeZ8jpk684DTkuM68yqa7EfqjozL+HWmpTl9yvO6E9tOXY47rAxFwVBl
77c6CmufCUpkH75NyHlu+UktOcnDvEPoexsqfVtuFWYjwyPtijlpvbPyD6jJO/J5
mqlT6aX4Swwtk8Tn0AWD/obDVkrzclE/vm5EpUVf0P4lKuwiINjpmkJNT2mLLK6H
034pkoxu+3cEEyIRk06/2I2DFSmhNQ3zbakn2umonQs6yeub7aOBVx8P+Rwl94eD
FDZ7rgN7JesVfi+v+bNsBhhIjE7w1ximkXRlnBGXpEFOrznlS9sWewcPw415vUVO
yw/wALSRcTJSYUWTmlduBSQ7ano8tNc7VY7/wY/HltaJt+Km/QtPL/WBufNkO8wo
/L4+mE4dJF0/uID+WUB4VNeMp2O9TmBFUBav5KfXxl8NMQ/WTTnLMVuI3IYfWpYD
odYRQ0wJVbLV2ie8fjbtyvGplq9YESFuBzmG5iaxlwPFNmGzfuhklYu9CtIcV7sc
5Q/7uLRiw2DpV1VaRRVd7EEgEq9AQ+9I23cyt1mikYtwZYzmYbgT76g9B6SoG8Ei
jA4vFnAprfytesP5cJlO4O77kOhfpnvDX7kw1Ouwy1diOyMfrSGVgKr/PcHwEx2n
3/+d/0wyPSYYJeQF3gAo8zKzqC09rgtUsNWL/PJU3eIBR2wpqlPJUTgPOiGufclk
oQnFzmU8VpncrBfdp3oj/Q0U8t2nrG+ilNzNDKglDpqEkSYzEPcycDYA0Nn8RpK3
7cO8YTcMT0U8VjbpgeL6L3A4QLM1xLlpU8yH3CCrcux4mp8XSXDio3fTjhHG/4u9
+M9OdYaNHB7mo+u1VQM3yys3CKlumHlmxk3pbEvb1QTGvtzzDqHyeGoB75BjQj/l
yqwSxfRoHbPG920JGWBzKnnV0SRD4RanB7Joeb3noYD7LJ/+G3pT3zFwgsgwUBlR
+CLA5zJwKDLIjzHUq66acziDq1CsMwwjdOFxTTRsEPfXtiA+i+IVTCD5An2VfzBb
7s438Y7oUsl0Uaq43QqQRcH7fF+n1lppB0dL+vUrNL24Ys8ddNGM8nxKG9KtHo8w
sQ3LeDIB5JHZ9x3SRguEqHxWW30Piw4bcqt6e9iEUTNX0tHSzkSQNuYZmDROw9hv
E27HGS6oGOdbhuFkq6Wu8Pwpx1gP3SPYIIQk2CKCekZH5Gz2mDoiOR3BBa1xr/UL
v5uVnCia52e7Nl+aGlyZ6WpmtfJlIQrPEkRskePlmede3tw7cb1Ip81551pAdeOg
BZPPjzgxuo0GtimjaeU+CbpSVZCWjdj2n+7UfmjeCVqPrJad2vygCBBKzdY1zMEC
2oIiPiA8V2qwsFyTC5Nceo8z0dCnGM5EckPMtGZrrg5CkURNjIGZ5l7OU2Z50yRb
UB3Z3ERTUsG8i246O6awAUPeQhFMJmnpmjlzP6pGhxK2tiqfqLQxRrU/ij9a47p5
Q8IUlCIGfySAttPvcpgvLfnk3Ht1yZrrdyOikRK2leN1JgMgWNUoy97Jfg0dgyTi
n2YhQ/9aYBqLE6/Bd+QseK8kC8HjYRdd59Q4WZl6ZoULQ2czLMBaUFzHXI0luTFt
cWmK9y8DHY785GGkiHV2mVBUrj+1iOOYKmSxGR9r6dfO0OeCHdAspZMWSUETLXne
astFfIOVmzzmTXadg2LqGIrQ4f7WD9HX6VBu1sOVxGUoKIuJgLTOvNHOBOqhVEjE
HMRNXgVPJR8SJYP160yNLJh/xeQT3vI6C2e+c9km0j5QM6Z4oNpbGAWHyKNVg//d
oVl/Nm6U0BfZeT2jcWi2IlMkPgqaxuyWZ1knACdmFYZw14EYzMuZaSKLKSR+Ltlw
eMeQI+l8ZPKYb5dSNJamPX8NcWM2dXeju2dLDditqw4/hq2zTqPUPDX6hWZ7SyNu
QEHS7IwNDsHurK9lbgsptKNKph8bzOof4/2qRmxkaage/l72XwpUTioNFZnY0mTY
zaFfuy6Urs123zIJoVCxNMtyGwyjBkIEnyn2NLEaA5r+MoTIMwvESX1DIHJyfQjP
7nRWxlv2cFXHtdCiN1ypUOp16SjM1wEVPP+kqk7abr7c1VIy2PPeeAAuICw3/C0i
WCvjwEU7/UBBrFPt4PRgup7lIsQd4ikKYC+MtVrJWaNVoecYM4CJfTRg9/amt5Yi
/AqYNpT6N00Cpf8W4JRxh/B3rA0E0+kJmsfBBgk7B1sw1clv9eyMILx+Z+rBMSV9
Mh5OyO23t/oQZbLBKDk15EbYRFjVKJf9PUkNPG1MKtBHGsQzQ0tFnKXDWGC9v/H2
rC0BmoqygMcowxkGqzEl2wQzzc7wK3NeyWiMYY9P1koq0TQB7/Q7WLuCtWYZY2On
e+FGUSfcZGiY2rN8PVQh6t0lSIX5gMhw70qxwneU740lyoqcl1XqiuBprtWm41Bz
viVHCvgQD2Afe5/eDj5LtbAn/dXYeYzlZlG8QirE9PNRLifqQ8frt+aqaP27wuLe
Y8kZflNjSMcTUMCYB25qozY1B+e6FVaSANxrf2ZfUlgddSZN9XUdvCdxLBwGG+kb
pKgyj3Psc/jyPQcDcXLJmkyaR6md+nv0m1b2iMotdPi/KrdzD/CwnqA7Ua/Cy0HV
r/9uMJTTbMM6HxHO6/i8dfjMNDemTosBG3FNVDQUoy0BtG9P+iWta1n0JWtWuTee
+WVCFea5ccetzQwmpc71XXAUn9RcR/Gxl917NhZ4tNBvOSmrKcgjdFDRSPYBrGLt
iwbgUNytYWoGLPPCRnAy7Nu36TsGKzTsgb6It53RWdLIqnG0jtV6Ux/K9bH2UCmU
uJtdostZYqde8ijcj1NY3kZjCR16IXC1Ci+TWeqoDPBgjMVMXErWjEpljQ4jQnW4
+kQ3HY0hVZCNkn0K8ANKBPnRLTr2NXPb0QEnPlI+x2lP1A4YIrCLjJ7ouaShaRY0
lFWL8HTm2kwRun9ycMy5S92mrrYKw67SQYuj1XVs8bLfIPvKy0iooY5hZxvvDEsj
bmUNph8WFz9l1xIQk8y+lSmi0JQ4hsoA9JE9kN7S2s15zlT0uOdrt472w9944Zwn
grN5mbHoqbrypEdbFUlBbTpXM06NUIBFFCh5USIDTswWSIzqZVvA0gqLvBwymbZ7
Lq1QaFspybY1INLyxHgffwpSmb/20blU+5V3daMRyhhSc6/GKbBQkmehH7NBQTLr
lFl1w4rsCFlcB0NDire4xl+7bX0DFiAH9hvTaJN2Q3CHSaxdi1MCgVQB78DAEOyg
jiiUiX40uyNuyUqVFH6EX23N5e8yxY9s17FJRkA4DpwIwIJlm+BAqcuQMt2kpOvZ
dtFN9kPsz3bD65fjkciEI/+V7aMgt6XFY/VI1VDTNsWjdxzreNRuc4NW0DcIUCzi
FabL/Add/D0eFfJYhdci1Su4HPhkZ0yKr64MudYu8EaZU3JxO6M1VepHrmVPuPb+
1S/u9FClcpuSusrL++Pb8IGFHXt6kQgrn10/K4KvvbGIFRQoggf0maY7MERgjTcj
dCbF9JGTZtaImRdRZnLssI+UctpobdbHOi84CjGHfdkjcY9NHj5tdmyA153H12cs
V7iNsteIsO208k5HbgFQ1pktDQNEdR4vzBGkvnUfHTx9Vr1e7nGcUbwmijW3+ne2
BBGDQSGItIskgFMFxfI/SuhnFU9E6r8SaT2oSPxQ77LVOl7Zm5sEqQ6F7rjc0+MR
Sndsl8Uh/3ne4t8Xiwx3JKhgTF64pVBa7bhy34PA2BdreIPkMo8iC50jHkLN3XBb
ZttS7UoqzesoOo4V4q4iXam9OtnQJ6SYJzedSJRv/lSZsA2PenPWoR6yiihoghGL
vhEyNIDjnAHGtZQpmKRAI/DPWIc42Ea0ef2iMyUW8ZikUX4ZYSI/FueqWwQNJ82J
lUxzUDVN+kvS/GVOD1o3jjMtfdLZHwQC1cGhywuKCVAzXPX723DPjbMfDrVQ9G0t
7HD1wtPU2H4+EE1fIUwCb7ZvMimjXiHH4bIDg6WbUEi+WrnN4cADKkQj/ccxlQMw
PYNUhzgvmUcus8Km6zPsBo6lOnWrLTVDk9GK3QBYZIk809s6NRbFolg3aRBaYNNx
RsO+C+ZVetIwGV13yzH0E/R9Qy/fvkNI9xX9/igxp77cP0WVFQ/YATo68KzdBD4/
hQedaOeHza9dcwMfFm+b5P9Z83/lz/vKmbeDHVOovncihYFLEb1RYvKcXe8qejTU
T1GdBhJP3hM9Dt03s2Y5pnZMa8+dSLGtLxaDjokx3U8GDUQ2TNczABTpbGHB3kPl
TaBG4PMdcKTeS3rhPes+9+Hx1tIPyTBv1SO2IOzl9QOWuajieovvPAcaNWiv5c7/
pCibRMH0cL4L8ERGhSJBKfKI1gQg+0wJSsmqHwRUF6GbW4EMm4hPHbrjJO21QQSw
pOtgidILtIa7RmfSwQ12GiR8VAxXjMIoy27Wnv9ZgUN7jX5e0Ii2u7+O3ZmrsbvO
8zc0TzSqBYhS5Df73FfiRzyFMynfbmck1bVI0iQmYKsPgMuKTfUSEE96jPZl9N9F
C0/U0Tw2ELL/12LSBp5CqlwJ/zERFhgjCsKnrfw4kLpHMWy9VF3wJlk9Ywj/3kF0
ThqGnJP00BQtNO8UQhPQo3i67wuK6swdE5i1DhB5aWA1KVCAmlEnbz6t/B2huiYM
etLaQeISnNKvWymo8NCy5E4vqLMNQ1LumTtOpuaEXDCvtMHhLgFJmAMRM7xlMeUQ
FaWYRwskfxbpep5uoEAh6Q73TwIZ/fMpKWtWBRoiNDzSXo20TA4tMfql0NyJe07I
YXDuC0qB435MwMKxx76rlCNVpWIsE5mrmBXBqTliRMLdydab6FPYcOYTpcdFDwP/
4D2l13T7LE3eQbYKXbijbXa+mw1SZpAoQImub7rwG0+BsExL8hitRjog12q+zL55
BAYAw/zwi2HxLVXCslnVhEcRIIasB9UgNvQSNSkdxcyeCXUVeSjtXGmpfWzuucVa
gXsLbYQ0j9MjoSBQReXoPVBKY3VTznitR31GLe1qhEt8+bKNM1BAO1U289m+UJ4d
x1m6WiYzR5wBEckF/UhRDyvOohUcyZ4aJ4rZTmxXhVp2THTSbdmuZCPs3Sf8TZQZ
aKNniUHLf3ZpSGyTvavlVkiu5lll3YEGN4YemY5kwkZKfaf1gEE++0F4j2tgleIV
2XRs8FQWrurwJYcBc9kwU4wO2pvSXK2YTBSgh0Po2xpLLQwv4nS2mFJDsKV07aum
qdQh/HQV36SQorj5sNE+VCA/9Imebm//znO8ZtalZDmgdbKtvWwatIZ0xu9oHJBp
jejLj1yPxtffgXq+JzyNxdfo3jl8FnfJv4yj2B6KfqC+3eCbFuO6DMgxIGCeX24Z
0laUbScaUjvzjtnHyi3A+aawEXjzlAykTXjUDNbpwmDGe3SfYCFrCyMGyG7soVN3
1uAxrhP6xQ4504qoBG562BBrt7m6iDtSDWn0XWOhXkKa41I+1B6HBe770oUkP+o2
DR/YjRpjyvasNQJOQeYkTFcQ0/Z9kGnrMnjxLF9FqzAqDrauXUC64zc5jEACE6AQ
2b4+J03Hz1j4PyuXtg1XWGFQzpM5N2NMozkY+iMkpPY35toGYq8J++vrRup9y4U0
LcoqWTMXeh9wQxRflBvwZRa0TfdvX3b82+3GsVti/RYDOCgqsYHsr8NVZauwSuxI
5FzGFvxahPpplxi7WQT0vefRvXNWR5K9lB8AP608u4HAlTK+QZAUiig5OVppGBJu
n4wPZNq50o5wamXSWR42X+ytc3jbfPpKiPLzTraBjrqWJsMl6h0sbrYiMQXSJgCm
FptjRRwlqxOk9jIz3HAN1kauxAGsjWXp/NIKrQTYTnJeJ+6bF1seLYEFL9gkU8QT
sY2fMNUjd5Sx9gVS0g7KZzrhlvco+43iINMcikdno2ot77weZqHIRj/DCjHTn+aX
x/j3tASA+J5kCX8M5fe29N0Tm6R+dXIo2Z/Rhmpzdzfr+3PVLUZiSgcmjoTSroW4
VAsderbRja+aulZZMjRaXaDXOBWZCCciDeG2FgS+LwnvypXK8LRhEq5bsQ/IDbpD
uuMfsoySSO2Gn0RVyyurhAfHweTB6WMDXfr4ix6MMmJMfjJv00GVg6aeGyB82Blg
VQW/Fzj2TN2h5hv4h96+uEejfs9/utMGLOYWoTjA8LVIyJjyI2iK8jaVrGkxHrTu
bf349X0L++AZib4inAPxZOPl/Wy1T7xqQV19KQzCMDbQTDQFWoafDGNwkZU9tQV5
wuebtXg3HiJP+AbwHL+73d2Gpw5ZoR9mYxEHFaBhoHW3izIj7fwu37n6vE1dijQB
z+6nTWAdhJOkUxVPWx8WoFoSs+K6g9+e99Qxmp9YmfP69NTNEWSV6CVrqb6CqOVM
zXjruZiKSNp9zzRJfw+dgF0pD4w/eKHDGSIL22rVPPvQZOz8/ft1RZsYDRlLk28R
VINwxPyKi5g57dy3E5xk5rRIXnt/tMLjmXmFfIOnmzGW3Z5HFGvKNAyUEW/t9JHn
7EYdkbvHbEWusbLUH+0ptiLZPpfu1L/b9BxnrasArybWZRpPge5frZChoevyrr0m
MpGXbAymeL66pUptQOxVmcI5kL9xI0JXwUaO/X2/2F1oskp9fOtm0IrTwNDU98r9
SmhaAtH/94DXZ/MA/y2b/RHRfoWl4W56wwU3+yOZa4PEmZ0ze5osA8LdIyOzwqSm
dywZQoOhFaEVsse0el0QSAWhH0gMgnlM1N2XDlDXUV3aX3nIPvG/c7E9VeWxihsk
FO58RtsnXtmV5WzhjpwWhgF11Wm3udpLguyBjCySCv2v3GwWsbiJapTin7vJ9MII
hgUvZ/XUAocpP2SEnG1T0ABzEVbyoPYJKM66fuROFHCJQRr1vKRr5Ct/SF++huS7
BuwkXqzcAN7D7W9Seo8D4fAxRKTMJcVxnfFAnNOzRRnXhfkipEc/MbH74ngBJbV9
2+9TpvcmOV0YlTU94bowLEiAd/EwlsJnKBrOurrhY1N3010oz5qx5y75LatOLMSb
3kjZJjQxFVeGlNJ62vbKunqE8RHCfIh2m/za6U6YICIcn5Xc5mnLBx/FTKBQQMeM
vOe5LVQIta1x3uLvz/SkazD3oZOu7X5Oq0WPyHc2xxQPmN2ZdhlhvflT/40+rF6j
JyI3Kq1ey4DZv9NcP5J8VLBDo9JI8PZXEIsQ1oz045zIDganC5Tz/1a7hLTZSgK8
TaGzytSDwVtKnzS11ZMue8+Bk6ElCzgXxLHTkW2ywkDu5AUJ6cxA7LQr7feUdftx
Tl29WnBxETbHtw+P6Irmu8aMmk7heJ3FyKkGSFnZTAXo+bW1hkbT79GP6t6VPEtv
rvMtVhrXe7GL+/lIg/fkz/yEUuqP2qwvlJAH93uMAdbyWWP6augRaTQc3PM3t+Ta
hYHoXLlWRVNH6JQPK+2bFxWIu0iGhMIOD94cFTFOsuY3Yip4iSHL8nfoxAmQCx9w
67IKb2GspCbDzmilNlZZkeyIdNzD/NhGw4QM8CQMcUPTm0U+rCQXbpCaRVxpDO4P
MzJxpCaiFz2lnVXTmstuER+uF6lta6Rzqd+Tkwh3Ww6EIJTAubHgkCxCrVu3dfXc
ikk8V+90FldflESMYBeYA7nAgpxuVh/A1e08j2E/T0r9RnwtXecT6eyb5eqEwnBT
ZJu5xFt3pxS1rOR89oWCLirKUFdR8dJvUI72Ym1JW0A9BrNr+/77o4PgtQcUqvbS
i+v+DQdYe9widCODfpIuXDrVQBfm4Q+UWA/aHjzxSGMB6hcxk5MMOBLmnCY3Ejyh
Eahii8TsVnjdWOkEHLY3yxs0nhXaTWevv9NUrlLAPHzGxaupTXFFIYjZqe12adXp
mbP34wnmrRQVGJIU559T1zTyNmfzVEzqpgeFsf/2Oy4dzIl6tTJOH0VSN7rsLQMO
cop30p4JlQxtUbOWjMX1EGsifDPmdRiX4hChoTyqtAmABoNnGe0ih+mvNbz4sprJ
J3x8cqNGJ55uSMH9l5THPT0L1EsuGpmCxrNFVD1l7uz6dsHfdVLg9FnqHmPKGlpv
Vmu3WSvMt/G5f1bFPXwP9rNIfpXn3+H81Lt33gXBfCIuR7jypQjmb15SSLeqngQx
jDX6MYqLXOgOSv48hhqIsNWIeCBhCGlW1pDPEsGa2ZjUEfvQ8IC15I4SliTLC5Me
z+BViPSOdAsXEkBZHsWfhszizjWTF/XkggkLy4rNOgyxMr26mDAa15MtqA/nquVG
T64gSa+Zl6RRjSo+wsSZo05HNiAnpXb3eKHTxfOUQJPUaxNhmeHrCBftxdL6OUvj
Rpr9FtYOEx2n3nPuLrOD+cqExtrRDYb8zz6WSmWmo5BkA+WSFrRj/kl68hI3zyW0
oqdPCTPNMNRqKwlzIBMQK+Fio7IxX4lGe0mJ5ochJd29pFY/KtyECRod4VyynLjd
Vfp1Vecv7rKG8abgNEde0T84mIQN249PMXB+7roYWaSGP0dfDNqL416F9dUPLOFv
/WFy5sQS1jDluPY5uGK+qm04ukxeg9/Wq9PMrbTxb4yhfjgzUXAvnKjBK+tc9BfY
KDyCNUvC4xAsl6AyDr/fsg3Xrh1+OyU49sbCHXakzkBBnmzZxvnjO0pKnXMnfWH3
RVtXRZJiUTdNNllEFM+EErtQadktrcAciE808jb7Sbto1AB8ykmcfPx92UaeaoE8
LvbER7NbZe1Vmg5NYB8N0vvjB/sjh07r+EP4/L3GDWIkwGiYawXujzfkicfh4PGQ
HVKHnHLJ9O9a9j4c7WTysNAqPAb/Q28HgyULc95msIUko7Euvu4kU5UtqA2VVkzE
2Azign0jNs9DMJZWnwDWkyDblpAZNoPGGZxulEsxZFeUSZ6X4pLehxaCgPtJ9TL0
Jevh/3UJsMGfptb5EfNuBeevEhTtL4ZGSLP/1waqAQxnA3CE7CYfg5zD/wOnR373
6tfjUPVSr7oUr3qouqHSpsHRtWfT8WXGowkcelTvZC2BbV/ZakNyZiAO7/G2N9AM
fO1Ve1pBoPoSzywEb2M/jKAo+R3x4/fN7g3k/ogvWdyFXGke9ZNsYny+8IoJw1bE
s/WK3BUWWp14eaTob0ocQJ0FPsPXchQC1/uMBwuT27KuJD5KHyiiP5EOWguIaRko
/ZXc4ETwCuyITmkjgaZTSFZpHfNIVcFOedXZsHiP0tCwUFmA/bSR8x8G230OYGO4
VKq5YsU4OWHrD3nXqluH1+3LQdqCavcwN6PPbGhlMcCCjM1zeVA3SYNukUT7ouVL
Z9WTSNGn1qWHUzH3fOHYHVOV9CnRmSe9i/oZM/7dZzVKtqd3RAP6r610cnOCZqKj
HkE6inR2ZJdrntaLKp0yNCcirF9tCQiEXbDtO2XjocHmmicVeOyTizluzA6XjhGA
vf4yICeGFzIm9kiOvAsmjdTE77/+9KtChJ79KkqTvruwn0wHsHvTWJ2f1EN4jYeO
SNG1Xe0j9bsorz9+1v3vVBYemBzox/sXpx+z/9vJj0hcLrOrtDQT6pBptLUOzmut
9jfkRJK5gJBGrc0Ak6QULqd9VW9d9Ple53kPESK0aH3Y7PMWxxNy74jHrIjYyW4E
uNTihOKQRtDsM26ktm3ftA8tZHnpn2aLc0toUHSfWCT1nLepuo0qasSlYcAloIl2
lyuQ5ofs8LEuQyfmnB+VA2qVRccYJ3tvfnq5xEkj/ejgWsqFMqULtkfJwsAn5cXh
etnNLPCjcmtOSwBhkKIwFa2UDQmRpYU5YKPKecAGxFBUrDUlf3P8gvEzRQucCSqi
4q36Ipa+orzz8WKx3/enEp/8Yi1wEfzkMg6i1gikIwRE7J0W3AOCrbIidG3iXVdi
cY8pr+sqy9sAJonjZc2/KqxmD35WHlCSvxWnYA/afFsR8MbEv/WmxQzzbDV99Y+I
vVJvKa1f3GMnKp+Fh1A/oFssFKTh5b3el589Iz6L+HBsRSlaqaxPcD+SRCdOhYja
Y4xGlCqYwYQI9AuMP15xO2XJineK10NAmAq6wzMAxiNZyRfktyO5C2LLeOlWrOTE
GcvlLgR/quSP3cpBZcnHR9vSPxHXbR3Q9mYvTv5u8IS/GbPLQtYgfc0BpQtCmvKU
0bCxVaD39b8qjIUQEplz51+oBjl/v1xP5rPByeUxCDGgaLmL0GwLNorQTrnLzmgA
1FYHknNkJFskntaYNParrB5j5rAmP+gxnYbE1ML0l7KXUW54j5MSgFw8UgkXZXEh
5AVNr2CkbVTBpqIsTNc774xatbvdxdGh5tHwZ6EVMeXJM7R/HIb5ZCRXeHi+FjIj
JWHpGqP6rMCtNqBeS/KhoDU1dMD+A/Uwj6Z0VqC/tx0EppCJCd1wGrEauRXQl6SZ
tK3N+9KcAnic+bjwdFAW0Vaks2PwATHXjb8XLkgWc0m4dHbK5ioVFcbPbtz/T3x/
c0qXIp0BEeXzS1gJK0rOllVWDC9YAhBlOpIOh33ul3BEKmi1kzSwO+w/tgxUlaz6
bgbi4aaj7tOhTrm340XZydhLo703V/oOeFqkrARRWqwVtecgiGme5AmkW5L3pzXF
zu6VHGGsDG1Vc1mSudbzdFVkHZeiwBlvGCSx6SnBzv2PV1cgZWeIYOZr2qu6FH/9
e8O+SORbig3afmjp2zMAttn1qd+PnNz9eIyZgs/q2GbyuatUY25SV0GgFcJNSfco
NB840/FuACXk/46KBCBfiKJqbSa/mBPK5l9xuU2HBnxvM4bW90WqMKX8FFWb89gk
7HmwC7+KcVeZ+IkRv6PrWrvPcjBl2FLAvd/Aaz5ccalPZcZd+DbKXjFY+8OfUUIc
WGri7WjTnd+5z+Ht7LNuRtqRvynAR4rDrThHnHEm8dlIwsRUorAnM896TB5uZ+Tz
FP508HjQluDZg7PoIkrUhy4/i5I+BvfHo78El2WiYQ+4/Gw1FBMu0bBEx7YxBR5e
3vZmBZZTs2lcLZB1q5uT7oz9Y9lzcJjOGxnmR/8c6yfxysKkocZr0IGfwpADBGF8
soBX6XAGm817waq3cmrvi23zSQh19URTMqDL5V+/tS+fxVIhzoAiSElYFhhhbdK7
Z5u//KrMXizD99tD1FJ+EzcqsrW9/sjQPFoZF5Sp4H/NJdNAtgqJ/Ru3SK2U5ViC
Njq3l1cGlai9F/KkKpjPJYGIDShErVGgFzI/+NHNCGvc7zInmg7TYCEjvycmINJg
2YRu/V/JHsBTeSjjE/fRJtHSTxM1lai6N1CzBUZb1iuC+zmT2Ugsia9aOfmj+GYH
DrVWOcB81vMV61CaLSh6oZ5ccffhAGjmN/SbII8Pis5YKgE+FsxntchgYbObUJhD
boBUmNpdtX4sLNsBmY84ApUyBRdUeE5ik+tiJzSfnYGseIWOEHW0gBu0ANwfip73
dDFfHdewJQ+HSgXbxXuU2KBSHwIpfd6ruOQ5ygyTefmI/2i0ErnujsmiAuQHUuvc
vjlbvXA11rmMuFKyx3UDr1iSBh44gyq8590KR1TzptgnquJ6LNrAs2/l7YASWSsm
wXScl7YkaStlPpHxkZ7QSWX38jq1IRRhovgBz03VtFsxH4ebiJVwD5UdotJMVZmF
/6/1hMKkHf7GL2sFcmEzugp4Brk9R2GRTwiulFcaW0trfBVmZXFtCIHVKf0KpZBA
ldic0M9WM0TmMTMn5nrjqHfJ+VYv+Ufzpwy2q8Sz7EGUs9IJNcbCLRc+PrnId/Qo
48vSxGipV92sLYe1vX2xqgLbhSKvzg7+GClyArJ1HLyOgmal36+e1fxzSBEKevm5
a15LqVHDKvnrNBG3mzR3TyPUTnNTrGZOpIQXtDLyEEDJ6GuwLwbfypJ8JvPfP5pv
UmnAFKJdkAzY8HQJBs3HTcM7RZIV9W+TDXdDTnC+PTZvsEAiR8CBxgLVZES1qIj2
cCARmYglhFuHZFTpi/ulhUhGgbN8CSgvdzOO6IJTQXrIblO+Eajmb4q/bBKiDD9D
zgbC+Kh1ZFvkk/XigKAxrK6uG0FDqwB4DcI9upD9vR2Q0WF0RqNGh+h1yko5jMYJ
tBldCmkMb2TSnlXDOojzj7mtxyJkQYHdJBvfW3c3kvlsLSwrTdSbIfvdo55hmvZy
hxoh8VkQyfnwtGJnj/VD6CFVniDBRIUP8NCNGBUQgCOg8H9h6c0J+6y+QuRRvfCy
OE4ONAbUX2ixUDq+OSesd4xDGkKd4jJmsK5xGyur/ufLLY1hQW8QFuM1G+Sgiwnw
knDzgeEsqEtAx1lwfmf3e99qX5TBp9ztchvGTfX15fkpTXVEb89bAkbIsZYPwCd5
z8qJr/vhevyENhKvJl+XiR74dYTaUaUcaefipEWrZGuI/rdo4cGDJBUffOU8srg2
oXe3MBJDl5OZwkXBLyF0aKkYHEY12nnkCb4vyac+dwCQeyTT/nlz0GxpQwYCEH0f
uc0OVRxqwI049cVfafUq/pyhYWGaT1BTE13nBkS0orL/0HnFU9X2R2UmdgAq3Ofj
QNYkSdNC53GZ5z+r1yvIxOFQtxc9rUG7fzWNzLt9LuDLou2MG3BQcS582cYmZxlQ
dwK6lYfXdICShD0y/qnc0qmMtc+VjDrgsiHWFaVgPygrb9MqHSG/2NR+7oVV7/eC
5RE8ZgawMcrci7x1PajOzg/fa7MmdNTXST+ldR2+wuVeLB+sXqUtKFa4gOBhuijA
WqeirMkmh+v/zPcnOTAhRyYWHWX+5Nw/Rfzb0oTjMedRcMzxE3Cxzj6TB4vv77nM
T6lSiMaO4cJarXWH2Uc5+SH+gZTGpAcSRWnhkwR9nAJOVp6NijOihQN+sqo0GEEp
rTyonufqqz2TtM89g3pqH7Zt2DNfjE+rtpzijZvcVccG9Im+pp+Tr+q9LsY7wKpi
xEkvDAiun3Ddvrs/THkZ+IHwAM3D6C18l6F59xbH5azg1l56LF6lNZFlVolSXRNd
GMPtaLY3GHaR8ST9CQKosU2FDRenf7GTaYtIC3D6hV9Pg647BzNDZyHwTpMNvoLU
pXRUWWAuwP7A9xgblkPspFsxwJa5h/FJHT3/K0aOZTyyBFr1emgNAOXqSuhg+0Kb
hruuWz+Dv/nHRZwdSwwWEna+Zq/BWhpMYKstiZS3TyZz96cJOkZOp5q3CxPyAl1i
MkkiTy85RwGXyyo0fnYysNsui0lgy73S6Iefm6wohmJq/7HEMdkUq7mfX7cOaT/p
jUt9SRly3u4Y878S+hitqychdf3Qfb3ChiuawRn0a4+zlajMRvQMTQNeHVavJE18
lLRJKAE2X07icK0Jio28NSTY9hKZXSb2ZgB5z6b5lqIXxAoLLnOnCZ+QWp0QWThI
c4t4295bF1Hn5dWxKanXQzhZtC8BadsZ9s+DLdCVLOnRn2R+tFJBSrvoDDymaw8q
kx5QHsqQURtbHBxSH1ckSKBTq3N6qwAM+BZ2mGDv8aUyktbia9zsq5ncKOABSVOn
5HiDrsSEBRJ1xU00T+SKRAGO4G5Zt4Gvhjnogn8qrc7B+sSV9ITgsnAVqxsdRcA9
M56E2RCink4XqD+bjIR7GMfIrnK2pVNmf+1/mbcNuAAsdpfacaJLHGi4lKusYTF4
KBcPNV32UcFRED7IhwsWu20/jWfM//NWdCOKVnGi2KgfV6hgSqWFwTt8mGzXJZHi
FdrG03daTDYmEJc3zRZTiFBDwiVQyyHotnicv+PVmKbzildxHCz7+Z6ygr6JYJLu
qgye5hkBhTsBr39yLEzAxHgqwUc8puPRahGlRiz2xfy/GM4Btppc0QhCemE+v7Iq
Q3KpdWfSF7IpeDblThncPwuU32UHHME//B0Eo2/Vk+nCXr8ASDFEMuKf4dcy1auC
Xf5HI8B3wTfkN8Vt/7ftOObphhab4O2jn41WarFBr+U0YD2NdO5/09RBXwr0t4iR
rCkdwQOmMikxKcbEOr8zs7WO6RhiBciDD71omFNn91qj2J+C9rZJLh5I/CnFA23w
TV4Ttkg5tpDbiXPHOwELiRRQTPgtfspQn7lp7TdzMcSD1UdvRYnlhDrDQ4bviZxa
zPGTbo14fM4RAUQMX4vPDk/ie9RRrEDWjG9EhHdtiBTj/qgxLoXqIDEBt5WZ/Z2B
n1fF/fWXiGJ47XNyECkrHprIEyHDISWeKXBmlV9/EfLm76u0i2XJx1R7t3Q2f/3P
IukKhjWnKdPyVhJT9KxhJQaft/c3AkKuwOQ50q2d/ZN392vVQksNpGYcYi4Bmpd/
w8GIzWqdNRgefl+B2jc0DdE92FVPYl79mjwC682BgRCG7nwbcuxko9jnvtoHH8Bq
66s/xnwR8fnmpzI13kquD3MFDQtxBNpnrVpMU0dJPMqSWYtxkHC25lZu3OYl7BQR
mchNhSWJtT34voYkFWWdYu/iCRILc9pWGxcp7JIPWX3a/1rBKSh5i4yTW+WGSKtq
f223ecSrozPxMj7W6LsWUIwP59zM0agvRiKPJFmutN1TCNMMtsHcUcDTxZIwaCtr
R6auzI/lTf8b6I5U5xgmSbXuwBgAg2wlcO+B3lqCNVtbVxKZ900LnnxXGXVlBKHf
bjdH83QHT02OuFnhy9PM3zp72ei1clv6UOvXJ3bxPFkR6UMvJPBn7KaWChVrVgnw
7MDOpaqBl7t+IdYuKxk11RM+D+FIF5Vq9LyNsre60h4fhDQBtXm2+xiLaUZyfacE
wRPnPTY/TeuRQ5O1KlMH+tG4ZmtTXkZD2GiHX6eYHJ7o6eizsM9YVzJJHYsN/qlO
fPcoyeZ+sNsqBOYuEiWOrb7NxKn0G5cSOn2LGIbw5XknFs6Du/6z8lUJm0zq0ZIU
x7rfYt4RueJZgnmuv+EgxOuJg7xCzsYV7DuVaTzWZHu0iAlSEa7F5fx6y3LkWWWH
f6vXqNWluK+K8xf5vniNsN7dKYE1Qttuhf+pA2b+b0NclBpIbKmIGx80VOoLsUdm
u0Qc+t8rcFEVmWz5cYbthNHPj3Gm1uztVz+ieBQPLOpLqr5t36gu9OCZBwpC4iEF
ZZyXju1Al8G3+pOGAMGH8Eh1fTs7Ku6+Pe6uGKEuvf9OnDqoi6UMI442uoiyhvwR
XxDziRukarLxPLFcnedp/eswdT1GCQG2D+/EA0Ye4TWR0oeAh8tDRk4+amGCfcrT
9mm8JBbiEWk/gN6PNTT6QovW0BrUG9cXvfxtdMy83YdWVTrm8meORujKA7ZmGAwT
CNOpTlukyQqTJWG1B5Jh6ok0CUodfYkC4qLfQhxR3saFKmFDjZTES1PAi/W7+Bos
7r6LcHX61U9SAKZnYIQW04wK4uTKEflHkockFl94OdJuCEa354e1wSfO9RZZIOnH
1ttZzzfNiUOAaynmH+SbjNUrQNLFDVwOo8iOpem8qck+P4KmylEdfdHJrL8q9YpC
jUIvhO2N1hRC8s0khCYPoeyCu5QfNhRFBl9eI9tSG3tCa7XIBtEPVnbqeYo8LQ7w
T+UYnU9uAiNvI1jDUD1tHeb9aIJ7gmkJ4QtiRCkH/51C5HZ73RucOim8rLVCHJ0v
1Xc0NqlZFSOnXH339DUiLLJdPFWDD8CrMBpevTHcI5+PKIcMRgZfZjAarY50yVpy
rU8Kf9+WYE9sCLqQbK1Z0yLfVfaxOADhRutLo0fayFIEop9OlnnaLDQYCgC/blxQ
lCYvqGpRiqP2s9EZEYqzgxh7UuoCxQwC6kktTpTRtiEmz32L0H9X8eSE6OXmve+f
IrVyrL8BFylgeWEmW0+CqIk1Fm+mx72Et43YRneTOyDk9Z3zLJBvOEYN37L56H1A
sOmySd46yD3yVaJwDx9tqWyk4JbDhqDAVVXxMkzj2DGmp+CURRCEC+/yDzmfz1h5
7p96M7Bn3hdETGVjk7DL04cI+CRErgfYyI1s0Qtb0hrtlCZ0xczAToQbIIwNfboe
/0SozQlf3esRoELpQLh9OkuXv2Ht82Tu02Sp0wlEL52f4h4+aEXkT4fDWWU0Wvx1
rSf8kPaX1KZLUhOsMTkINB02B1MGh3JBMdRzqlgwWJzb+Dp0ebYVFg+szjSPiA7p
0pHjiclekiCw7auzE/NPT0dRtB2+zfS4WATn+XIRIdFar97v84NKQDVDx+XBp8md
QhVAm4yX2MDTdH4dSTuFDyGeFOXyGJ80BZcA14s+d+pP05PCX7vIpoZPDtkOJAm3
2sn2LAGDP2PJk/9OeJAetOQaAWY0phJGv6+gJnlGzctyrdElh9UuVROo/wCB3QxC
Q4tiD0o3s58SwaUjOYcbABegQI77bKcso3F4ld/Uh+n1pUq0MNQHdZHywD38pUBh
kmRA3k2r28HcVSlUU2yPiyb6OKb2tZP/oUeuMuPtIPJ0y0HmHOAr9eJCM9OB6ewH
0QLMlVGZbGfFjVq8cJcb8OXxZlhg8EEewFrXJQR8cLL8piWzUCe4jAKO/NSUJ8qC
sZ7J3iY7bgygTRzdhm33mAMXtL6/6H/EmzDgUtABtISVdrYbQ27Ns4xyRIYk7RyN
6dvlc7PyHpsUzfjg8KqclNw+7MS7zm+C8daBpGVGoMGK7a7nq9LcKZC6LZdH/Za9
wNBfH6nTkmzOuOxFG35E0E+cViOjtFYqrBXLdXtedlmv2IBekc6aGwz8QH8qeAu0
jPZdnDw/7yib/6PNr5W5i4158fP9sTLDZWcA1s78kj6nU+VV398Q38Ov68Hny9op
6h6fJoKpoWb4x0YVEKVeRMNa4v++JMdGivkpBo35EGIsJu8tJI1lUaQBPbJbrkZ2
nPVxI0pT9AEVMaSAzLlfkElrwAh5lYjpvd25C05s/2PXU3i8RvAdW6lhh0zTuSNc
CObo8DJPaviCehWkr6NaJuK4hiPw2Jc5XG5ibrP4z11eW3wN+3wkwNaLEBbUBdpR
IHygoapgX2Vz4nxgaDyBa8TFUpFlbl5+HzK1tOYcvQInzYLmp3c9SyhM0sKCNuFi
v1Ory7BGUmebp1toiLHKJa15WCF4h/z4IgtJpcQXF+0DlhT8tuY/BfTsHmZWe/uJ
Zb1FcO4Qy7CSk1x5/NCa5XJ8CX5/HqjLpnzsbKGPEm8IxFU3PeEAbwneoEEAB2AG
gsHrvzgN/7Tn9CqJ+dT1gMN4IGNbGg36wrLRTcU94JeTOrw7xYHIk1vFqzjsDDsq
n53ZOtxVXnJ8P9vq8nW5SukWUWeXgB29+MpDLqKoBU7PsB21rbqt602Bz21KB+wW
tEpxlyYOSx8aTScvqP/v2eebta3yTOyjMcXKVV3LWglvRuvvOSsXFIP8kfPQL6IO
3YiR4osuSBHlxk+vLAnnvNNC15U0pXI5oE3LoPwhU0/1VoqMpx8G4pX1Fh7J88wK
axO3mz/t1dSUIiFY3F4b/AuMZn10E4JnsEG6DagGk7+/k9gvxO6pbwVRSTGD8NkD
sHK/f2foElVsuiUG804fUDIYEQnVcwXZZjSzWu4Kav2ONeizO0UaaVn3QWg/gLoP
ZlZZ/f49o/7bPO7Y6zMaWOgQqMSKwKuYYJpB7eLLonGOKMJAjbNvG/jFmGij2k4c
WvumbaOksDNP7qrJ9mLxcR5u8pFQR+FzPa0ApLI5Al21FPm41mJfFBSqFdEA8Mgg
0f92au8WEvJqJkt+VAhLEfS0/8sRHxvPeYO+hP2/fgxjgnGVbP03uDV8bk7MpXM+
YXWBLIo26xpwBwO09pd0toCpKQdwltQpSfANOS42B0NZJ4zjOoiivFRtx4QqB5Zt
Kc1WEV13LDqRfntcwUsR9TNHMbMUdtCS1B0MDEdin6QBp2l7yk1TLkVa0STgMmNJ
qiGcL0YAfW/ufRbwjpsM1SD1NlmcoklBMzpQM4s0ZsI+2jpatH7N8ThbSuFiGy00
JIP0PKsVgwzs1hnrM//6FNXJAcgb1itlhsFLx6TwK/8A0XMfKligif4ntZK7e885
rtLdn4XfeLC5eN1RcunUTPPGS4o39ujoDzxIz7Q3SHAEcp1srWhY9W1BCkjQ4vQA
KUPoYk7dJRov82LjHWkfgUZNIKQ4ZWMJyCx97efR1wdmOzDfW066rZyfXnWpZGHI
1dK7O33UlwO4snuxMctYRIM9GpwN5UGcMvktUAP4kkYr4/aLb0n67Ole0lu04ACf
FK9J6Swj6YlxeqEJMOBO2Lree8JC6LT0uBngh+2t6YUitXklIICS/qoOL2cf9Jf0
D4pjUozvs7ESifjRiEXDklGNfzu9ns1e/fEIcZFyn5jKmUKeYlSH7iq/ivoky96Z
YaiNR4VSfw5bKIli1+EHvBf/yah9ucPtyQbmOKs/b8nuknI1enbtjwhDZF8SIKMN
bnVHQBxMJRaItQiL4yw5zlzYvkDjO0gJAzIDeKy4oMc7DIxmprfdMdLjWT0OgbpP
vNB4uysYupoHakV6kc5WvPwbLjLWglH161dcATnVxJavQWDgRTSBsR93uv81piUj
4gPXwbq4G1HyrQNtaOfXdlp7kLd6BSfVmxmJvMvKGKOCLl1kyDQBuUuGnnfCzwto
LyJDs4ftn3qtnsvHI+CQRw+gOEMUIi2FWQFTQ2Q+RfEjaJIR2UQjkakGB/+Y8p/J
SrVVwBj4nSCjE63szuzBvRQdifba1Tl68CBfq8wJnu8EpfJXqC9VJ/Jez1h2leRz
O24gafPjwRqKG0J0WW7aBbleBZJfV2GZhKfrQJr2STLcLomxWigB49d3RK93w7P6
jC7LEXEXhw8uY7Qk7+g3o1QYu6wcouvjAOgdtWVPej6w3/1R9qBjOSCdAcVVOSf9
T7sgAPUlyLNBYRN8bjWmDXup1iBfE0EWYLMANEVZTABR/KCVtDC3+MiXUsSImigo
tBqB3n0uyjxlkuwfysX5pY0N6erk3MuzgrBF7bVKttSOPKmT8y7FsIkYMg6viuB4
G1kttklkzVgFK/wg48dEtS5vHkSxAJ33Y6xSJ0E1jOYLcHD3TuXcqqd8Fq1HjNKy
s+ufc1Robo5qRUE7fT1AY1xowO5wSXDRqbbMi0upPQxNDvrVu0/Aq2PkKFjj3XZg
h3iKPuou67epst/ZA/RUrNsxeMdmOgKTyyNnt+jlZHvNpCQP0hE22BYKpXIU/Ta1
gvU2v1lfA6eC3KGUUi3REN/Kju5zvpRiu3TB5KzKmtMTqvkBldc5mts+BwPh/dfY
vjzsTlJ0BuE0lplPsR20loC7fgtmmzp/xV0tx4kKwAnggfPeXK8AoS6sROFS41ko
CK5WixswuCuDk/V3JsvfDusQfnuTfqu2WZ5da6NFyoEoBVjZN217E8hNAQDHCvFh
9RTHqjbvblNPj64RLr3JdrIcU0Fxpn/MebNnov0L8awEYVAAIB2jfNhVeS+8bVUs
N+NtjXXj1hf5iBIf0lWUWVmGZwDbmT/7DJryC2e/J4fnn2XxbjPN+u6iDkPt8Dck
orcA704j+raRk3/hE4cljWc/jDJxSPU/GOOEb1SK7prH2M55mZxnayGJy8Dzkc/Q
mL+q5HYEqumPXSAGGdN4sr/Z1A6JBNz08Z7ZsMhhbRL2MLNnX5trBZrxlX/mTlAT
LTRTA4oeLtOtvlGWXRPet9NxUiLtogzymKxFLvelhvB6r9tWZQ+a/R7PSdNzZMyF
os6xVlXbwfr5vmqblPnelteV6hbuG9xbKe9HqWH6a+BGp3C2yRUEJPGVAfWK4SNg
YULMrayn7gNbdE057v7mOpt7ircudaygDi9tySJum2Q1LxIBJPYFo7IsguSAaEd2
O2p+Q66d4/CEFiUCu2Y8zO5C+KfzZzlwxyITAOQ8ENxQecmREyMDkpzTrGs89BrT
9i9NpuFQHi2iFFRPVznMYQKaXADWtkPCkxDlECkzm+Rx6/AsAQC9zIBIlizgAbMa
xgkihzviHd61sggfJ5FJzZCC4fhVH0StjRAW4ypMA9lF+Jx8qdGcz10Lx5d8RDEs
LVZmcLgARSQ/Y7K7sibxQt8Aagi93kqeFAd2ZBv8qN695DB0ZjOAvja5mh8A6ZWS
7yTjUVILgSy8OIy/i9fiMD++XBPZmTMBy3H1n3smb9AgFPVzE5BJTB/wAAsnGOn7
UEXtxIweTbhxmBhvMPcgqWV19HIFcZ7w3mMVstMPY5dOJ/mytOS5FBpS4uFQaPNk
fiKa5e7xvMyzQETUXOvA3EjB50odI1YjGw+TzdVE/JfI48suujKYX9ii7nZDUBkn
yEpX+skx7c0XIFFtyK8EDOEMzW17z/9PBGGlNo2Y1/NzoRChW2558G7ycdBKy9Rc
abubox+yX3+6jZ2oZm1u+zHsSNBWF4a9/xHpgrF9CDjYnm3BuQ1O2IzQIgI67DAn
joA4OyR7pyg8+3ABvLy84J9vrXJmVpN9fK5evKV9jWE337dhN+RGpd0EQpAQDCWX
Bz8fSIBbEAM568QyJDXO601t8nwMvHp1al8qCSSJ7uNsXuRYuw0gma6YHae3D/w4
n3xf7wnf5b99eSSvbaqobSGpmFszv7YRdgHAiFVC4CDF9oCKm7ds/ZKF3+jBSYJi
cu9qxTwoJtGF3alXkXhxsIqFqg8bDNebsC0a26IYMJJDncyfVEmQNznr+UWH5JV3
fPIeFsjtQs+Y7qfYWbFSCLfSzpaJPHTSzdO5bI76IM9fa3oB6gzZJBQI6UDSeH5P
n4v1HcSk7LtdpvMDn1z9vGXPynEQQrPO9c/uFvOaun0WdmSgK4/D4sU2glLMx6We
A0Qbv/Ne7p/powmOzutth4nKQChDWUtHHFqWlpdh8fuBBxWzuT2a4oxzKNu02mEw
3uHhpEw7mVbdtVSTvnPal08r0lq/2m/028QYH8KHqZAHo0VkrtpIgvsPKZ0VYiOV
hrexbzI3M1jPmskS7nP49OK4TupiYi0hPBIcWLdJrIz0P8ENB1BEWoO+S0Ixg5tw
H7q4tuLILTvNxJ5jTt/0b5SPdqPS4E2YlyLonox+/yNr7ZmHLPVsWtznv3NQOnZA
GaxghXkFpC/I50rhP5xXhmbkEKLz62rLHhrmEPy5Yq5O32I03vn3bfK3DOEBffQx
Svt9RVpXWU4HvgvTIXVQndHTeWtPLSebI6EAA+sx3Ob1Fap8rHW1Y2WSnMvz7uDR
KEv3RohC02HcdKrtti/HZYcGJagUcz2/Yu8U/Gs817BZ8hHKjmYkO0VrBPi9pWur
WJGbKsxKb+dQaKDVwL98zVIfgB5jFBRuW/GShn7TyI/tkx+pOYz/o3bpWf1q02Fj
hDMJFaD4HuaExopjI++0O1OMzoi0h3LFGJvBFyigx0q7pPrMMUs6iwSYFkXfg6QR
EKa7YH59J6SJ6HoQRZn3tnhC7Crw4oR8HBqZ/AJdSToEszuBImyCsEK+EyIRJ9M1
aZiWvLwz4BSsGcvcNaMv+VQQPdnjrywXqS+DcnhgZr8SIa5mgTGic+7vkUC3zwTp
faCINNH4o2P3e+yEYyqMXDtaRAG2K80+Dzispjdr6sH1RAz7dTy8JLVxehYd1reL
hKAh70sivqaCsmA4D2QkS1/mJmbsRVBLAx+np7qX6hwDHArQ0I21KLUODPnPwTq1
KJTeKlrzOESJ95ZR9thDDY1rNjw5lR0S6ffNEOLXokR5FdiqkwLUrB22CifdvjY8
VISFCLEPQWgJ1hLvG/qohkJzsWyqyUkpwV0dMM2Od6zh11GhidhyvKpzn13ugd/+
4O5HnunOGpTrpSN41mYnbpcFnBJwUnpqI8MVZqPUEYtMg/K967tv7tudsZMH4dr2
Ac9eFJyc4nhe23/E86o+t8V3QSrOCkC04W5bJc2Ux21FH+lDYmTqnx3tvlgfsVnr
sJ7M4bB6wV7DzSb+KhZlSykmBk/M6Nsytox/aEr7OJANW9LGeLxJWNQZQaVx6X9q
xs6hfx0xQ3JcjnXt93GsNhntkLj+WwMcM2Q4iRok8NJf/aC28OLMvTW7tw7IoP47
DVzaChB1Ix0deITIKA/vRtQzYUlfgsEVaWiIIws0tmuVJg8KFh7arwweDjU3vTwg
D8ksVdmcwdc+kAdpaEIxgYjACQhhsWwJsq+EKjHYwWiLSFwZWnp5Ltj+Z9oyoTF+
xkyiqgpwDEz9UDeJZajxqSpkUAIWTvoWNdtUrr1UvmzhdYSwK/aa7YUrUwhh0l+k
DxtZlQIX37aS+MCi/83jPPjcPuCWXhhnKeQFOxUHwXsT1TR+v9Npjp1OFZbllqUa
30TOUMEo9Yoz3Orhbb8P4BUiG4K5a+LzljBvINsgKIEe9FUnwMj78kvaPQkm03rc
EWifDeSj2oHKYRSCg0yzneSxCsJsD4fQpdhUkDRChGsbyljIvU16fJ2t9ScF9RUA
KeEyXWS0IfPxF6ap/Xpx3PJyUiyDCgtqtARiBHgvF7Y0Ed5ya7dnQAde5uk9BrWB
osEApqHf5UgTdmfXnPRHDEhZzUNzRZkRf7SJEy71WXywo5Dstiun4b2rNhe5aYqx
fov+55d4/1uD/fzxcLNdr3CDERHmbpAdEK1bRREzaf1bA/edlW3PRQzYyYK/rCvY
DeXnug3S/B+zypm5kgDvogKnDlFD5hZaoKDBGuy5bFJxHJOntaea3V41xl3KYMv9
/qepEbpDy//rVu9VJhChJ8XfIz2gae9nsFNH+b94ABFrnxJOTzquYItmSJP6L5zD
oGCFaYUGKlLxxjTvDeq170ea/MOctTy7U2mXwMmwxOU/qSOvM+y+lIiV7mv3aoFz
1jwQoCwLjVNBn5ZY6YwoojPBUjhQWJKtKBkAgHUk9pXi71o1uzBbNRe7Rfm2f8Ae
XQAGNOi+5lLKeQ77jYvPLDiuHTTB20yGQn9BMknlXwt5H+KHGVP9KuCWNT5cLAEJ
lz5TzfmWPiD6p1q9tpO5mWGsTykkwioRxWO+u6UuiOE4ERdfLKMG9NnOI4e5Cv+X
SGg6xhhkv/YPKWHqJ/mHftpTZd/Gi7BS5cfnUlG+98GnVsQ5efj26OvCIKvMgX3S
5763bgihP/ojZ+BEok7DIKJQwvHBMbOPVraE2SfT9aiP8FqGzrZmNRPIxudIUKyD
O95HTzhIjhlmBVr503xRlY9+jUmQZ7meAJInk0XdJna11Gk2jC6hNkiMKstwnF2V
5EOfQCu3OvYDxDZ+Z9tKEyn12k+cB1zqf19kMlcY2WeEzD/txuoRI1dpsoeWYo8W
MLMogitOPh/ZL5iDsS3lKY1batCXq9yD95pZJXcYc4CgeC1qK2nQemhw+5Xgc2pZ
AMcUlXWVQJtG/vUtkQ7qW6wg7FznjbKw9SRvGK7My43pMHqjAUYkVPoaH7PLtTDF
qwcumKqSvclmTNDxR2LMh8d/CxSdOBOUMDQJnAJW+BsNl5uHG68+yBsIECL4KAOs
Cl7nhwxLkcQLkjQjKL/b4yMdykaAIZeGncOyVQHcj7wgPcYGHDH3JwJo803nyUhw
cve6gOKA0hjY4D7r5obgF3pwuwAe6Avfci4ZUEqkx+LtMfggStOgvPuaYMq6lNQU
UOMXWF35UqUQUjPR2i99XwuFps2kuuk56qWsOQW4qSpXh8zQLIlgWgoesE2zG1uf
HbQm70v1ik1ds0cGfBket5mgUe7rMOrjmxg/mt7wI3TeGvW50M7rtaEtOZ6Wmn2M
tRzrVv7NOCukMu04NCSybTrTF1FtilwCajUKF4ZIHZi+ezoJtmGATRi8iaenhHjP
ljZt9evDr7PwIbqUdARBLk/scj07NFsrR9YiI+SHo9Iq93wNOTTu3TNkd9GJB7D5
+66OJWkifprIF8i5g4CA6r0zccJ6uOC+RjLINsA9g4X3IAf46/h7jEFX7CT7feNF
EfKiumc3/m4a8ttnwxIUmLHHWAGyhZxM8DCrmGi8lIc75sGmnETjRN+Jj7Jg/xLP
vWKQSxRDrL3Kjeo4YoBys/OzXTa1YWyTAc1lRNGfykMikZdIyo6dSMX3OLN//KPD
p5P5l8Hfi83Wg1QvZFeD9hjKor0pAGI16Ro59s0oZAoLMBVwN/0nluzlEj1jiUk/
fDIhHnOHL3Xu10B4ypAnSIzKIKCg1Gc/7lQRlgqQkDcXNIbMGFtrMUjmIzSGD+5j
axK5OiOFkjrrqUufTrkftWFWV6AZjgqeRPzfHKsplSquB7vwA3JI5CMyqdGWPh8U
ACE5EfW4D7mgdRqbn0EUE2RO158jd9j1JSXZVYxunmXT4YX1llXQvJsxvFk96VLt
MG9JXQ+xb65fkIuV/bfyeJq7X/0ShFycC9X1AbPk76G3xiYYINvqjwlqg1Yw19LO
BtlH9dSURNYXn8ACxsAhHCsEoDW0g49w2IoUC2WMi5uJtxTicbcQFS0J5iIXSxuR
4fDJPVBTxflGAoul9JVww3H9ZHFrUVoFHquM6TgLLrBDrYxBSntmvRcJpKR+DL9X
7GfEwrCD4ghbL95LogEkYe66uQZR3W58UnXsHQUUsLEZYUQxHRVowZhpPF5XI3yk
7OFwZUioSsNFNIFwrTOF0IDy8R/d5yJe4JyGaNgWiEceqL61k2edq1KCGX+eRO+p
Q7F/RThi8zGP+dajYxQvuG2J4TaHJKLawJj6nZTgd+4LAaqg7nu8zXdOThF6ycUx
Fje02gW4I56k9vL9Eyu0Lf8ON+iKZ+Y5dJV736cjJEysuh5Tm67aYQLD2krl5FEg
83xNDXknx69tmUVz4uvdvUQys3yyHTBF1VRPKFr8tt9dnDLLMm1vx78RjVc3oSbI
9fBcDN9UGVozIz7lEXxkiefnr64evPSHDK4grkxlBTu/tIWxyl2XPU+X1SIQyl4h
`protect end_protected