`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 19632 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
sTHDbAcNdRVMi738hx0vzltuEBGe4K5uPEdMunCWo0iPSGw90DdkfqXGid3d/2vf
vhFRlfe3O0SgmXScsxVR5JQ53jM1qVSKoNQ5SLUBxSndVViFoMRDCEuabJQc/Ytu
l9+jc3xGshN38pDGrE6mBe+rHO4vlL1ZcBRSjWjFgRDqkbcZ1GlvOkBGVZq3Q3vk
ULAlYyuxunh54PznJrZAbZe1ge4RBrnBCeOKx1c+dPwxP4piYB2/uettfK+Wd8NY
mAsLFWNZBXyzqIrboOzB+fMaI1oRk12z1vPTUj+AICNeVvPgk2CBjhnJ4htm0l10
J16uIpivACixO90kl/5mWU1e3PA0p+kQQt+eRD+FPU4JvF5wa1OzGl+tuCHTpZSH
rMF0rHNmoWqLF7yZmDH4mtx9TKB5E/oBWCV9DV/gxH2gbcNEJRE/quuZdtC9wA59
TwhKxNelk5BECnEv7nhdMRW+g38KEIDFHS67PCccE2gRoNR6Tn3MACvcgJnp9gS+
R4vqnYDSp/HI3+8pDzdEfyml0lzEap3pRiksFeR13+IIwftp0T4ADmMERBmLqBb3
6OWBmad7skXURRETMlYAEb7n46iQYXKhyr/6XEvjk3Dmy6WJHC8AtOlgPK9o84ss
VMbXEPNHPRRksPiSZrfZ/PI/OP4RdJdOpv9S2E+MopyF/S5MEY7JGm9JJ3YKXtJx
8yKto+/Kts5oWhNjWlLOyobWpd98gMv88s6Z9DfBwtQef8lCh6p3PrDfnFso29pE
noJESiHKfHThruxkJ0Ixd3127///0qI8uMvQdQkehuqMtqMYlhsf4rHjEM4mG9zn
9S2UmJikIl1be5QVWr6DL5EviWGEvgHltn1ZgaRauI5dSJ5um/qhqjZSduo90CXd
SAFipz3aZraqj3tnQtOBfAiqIuzdJpC2HzMtK4DX6C8czBnLD4xDEeJTgIJ32KZo
PJRTw9AStBuwByzuAJvxRkiWvc9DUkb3mGug+8lzQYi4MEvU0UaqAtmKKfN7KMRw
or/O/kRO9rcSYpWGDZd3xw24wV+JHRhxS1W6Lz1g1AFVSpzn6dD+64VfwD4slWrG
f6YGzZkT2dTDw46BVrf7rDDelXzJwCuEjtEdcEQXQ5ybwQwMoKZjDJ93olkTFRjc
7AHW/QB/R1V6ETVNQdON7D7h64q7eEtyN8auQkZkHI91+ziVwrJSCB6Kbzz5i8GL
m8MYbujmGNKDEW0QY9jjFx1+ZbbaqZfLYHqC4wh9AQt+7DOhQq1v6PABpm+p8ZXQ
ROPV9r4JAZfVx3QS6Py9bedAE2Z3Fee9ZRWsOUdekLbKC+QKXx5lp58QbZjP4a21
LGHmzlWijjj2yGd1dXC0xTzeacozMYdr5DeXtyeBR4476HMe8nSIyZ7TmOjL2wWJ
05wDeUeSfhwUxjOA3yVup3jUYF2H2Y+WlDy6RQ62165K2a5iVs5lUtMKAQE/KWPn
gTKEIjMc3UHoGf+hR2rhVG7OQLe5462L65A7ipyC5d6EIp+C1bLze9okk9KuK5eZ
1kgVW83dYYoTYcXAM3xjQ3PZlZ5JjyQ0fmYJjKfGIcQUTkJyHX3bmz68EwIjLaTG
R29yiUnLkpkJayPHk8j/Tg+3EQZDgahFZvWG22C9c9oFEb3Iit763rC2geXvwxQD
QKWGropaiXBPrJPzCttvbC5tvxsKBg2rPayhxT8pgRJYh8mpAO/7YptJcI0DhptR
E8xAQ6tW4mmHu28GDlV6oTSidZ187HE2rTonQ91LTrnMt8ySjkfKgzWfcudk7vcF
Hdi1PzTCTkiMP5xAFkj3WLqZfTZ3E+kSGelUdffGEbqg8lQJRVSTeg1x9OJkITRb
ONPXEnZ+JHkw5VAWrXE9utrXCanWAeE5ynQaBGKh1lfa+XAThyZBMf4H6Ndc9y10
46wRF3eI0qxHl0ia/HxSGBIsQB16yAjiC/eqtxTAQbV6uDZDeJFJpKrzg67G7wNd
k0oHTGqb6PCkFXoXFf4QzuIkBLecneRLe6gDp7rIXAsEt2+jDKFnnNzmjKPCXfCT
/LzXwdbPnBfRwZ4ShQ/9+rDuzBxW5fDy+eXm1jt23mSBH5VHBX3nGVJcDsscDgAp
tomP9d7/1ZuF36KfXtd5ubJ3QqAm3pglfp7w/+BLWQHTSdp4n5knswPiG6S31mch
yJOgWUX6jZGO2AO29sEaFYFkgKU3eYMw3RnTW1xbgd8xaLFeaChs2DcLAp6CQksk
AY4DNex7tkizsMoMOtFiw8ecGRvftdruR50TyEqLRZZFmZPcYxneRVxvDv3t46S5
vmgXAvzMFJ3kJQ2FaYmzdsL767ROY+XNzlLqhwHBWftP6zECcShc737oa60CXdSK
c5kJGSj8zC2eu8af3tbk+Df5dRaHYq4XiVqPTfo7K840sAzVtYqiDPHATY3PeyMg
wpXkGWFWlemc1DOoi5pA0DenjBlt1Unl+QfTwYsvRnRidZncAkGNBXfLvetRjzpi
aWVeHp50aUGVorv3fojXAV/unV/q180s/13cDuCsZIa2ahNqBNulKnY/7WWR+peV
6EgIFbUx9pKETvdRPOi+qw7CoBisgjw/TASIqrOmPSqy0pSF16uKnUhMxEZp6hAv
qcUjPoA7N+wMv0SJXEAO4fxxbzxpf36ICkkNtW0OlhkS3CUXq5u04un0IpDXb9qE
l/IE/4gzhqwMWrR4VUo5uLEg/XQiev9xUrfcSra+1HRKPSruUIuMB/Fb+yiQ2Mt5
1Ugj4W5RnMeX4pLZZdLSeYyX/kSUNBUpNxlJfvOBfmQdo29wuIzpRAZCcs5BxGWu
zvd2K3N1u3QVnfQmXpujooXLuGk1syfhAaJEoz0ue4Unoj4Rk3P8onvrUTFw/4Lt
8Sf5ZyHTnCagkW1nHGtOpzCyCuC8A4V9//NVhJds6/SRaDwh1rntGXg0XAH1DrOr
VFKM6cYXSShy4ik5e25fULn39VXkO5zRghLNpzWYKka24RiWSB4nMbPrhE7+9LBc
5aHJdayo4//zzcFq2fkmJKojzYNmIqfyuNF2AwZRk50hPcJ2E25cnW+AJhIUhyv+
+Vg6FTiPXXGwkTh4ZOW+74imt/moh6Y9bnHw4tyhiL7cOirTzSVCDivo+R7DCw4A
21PrANJvKAyV2PYlXoeoIsFVqocjB/hVrEZXmtzlseRblArb5xBpQIjekGAFWuG8
mTKpyTFFpXIOU4APkCstt59yL3ZDUXxeR++2VFBdi5K+lURyxelI28bOi7ulW0t3
82yNpRXUfJN44bCzmKjtbwSgUDAhWOeDytP+JVkS0MlpB9NElbqzvnqKaLaiZXsy
DTv927YOnM1CEjEzWCYrBUCgMOv6OT9tvTMcxT+wgoJnLNA4tIY/pYfi03Uo3L8Y
vN3rlGTsqXody8NSyjCj97I1XJC1pNtiLqXZqRt+FHldxiZ7wKhhkpajGPpTRZux
3mJ2ZQISge+JcNg3L6sgxhLCfKoN0sIPrLlrv8WU0zDpXZYpIIBieVz6+TvAcOcj
uFe0NrRyR8qBqSeSlc565edW8ZN4uv8RkDFAaoLFWfdpWPjjoVh0Kum2naJwEH2Q
NsB02FETxo7qXMO+u71xPxXkiYKLJbHltrsZu2IlqrZydGqzMdLajTPTmRaKIBiM
xi8OyZ+AqFU81hX9SQjSJFfVDtRq/x7UqnezTNVqP7pcPOFtimZvgvTsulYgZPwm
LoOnmIAhhEnTxt4/MqwUFktEjoyu8gWQKWYvlDBKuQM1R6MN444qyIWGfSM2iaLz
k+dj2FWIm0Sl5xvrffvfjOLeOXJQH3X/R3BArks8Dzw1INm7loJey56F5/1IMaoR
ahzJbL3AyDvOrsrTcKC3DW5s8mwdz2SMoag6yddWr26v2wkOYa2Di43nke87q1It
WIq5FSr2Tw4DL3JxtIljMnIhyw9ysgNZyKYWEclNyT8Guqud5YUv6sRlpu/TkGgr
NXFYALag8qHV2i7HNq3WWA+NWAhhK+4tSG33c5J5dcm5YW6aYMGmIuQqsu0T+x2Q
aWfumS8eBbW0qEdIES72I1Kf//L3O8C2usOAbNq34IuvO0jv775sS3/EbBA7v+OS
KdpZR6lbdhGlftxWaoJfZhZZDuvTg2sEgbqb1R1CysTWXiBik0eHZd/ueioB8afu
9dhLCfeBLy8GGjBRNNTzggqS98RFCxXIlba9K54US5pHP3MrWY1UPvY7qTLuJ4to
lTh4c7auOXfQE0gwbzQkbabSgXza+orfndj1WoAaHGALYwFYPGp7V/MW2rr13RiN
aIha42zKU4jA+pOdiWn+qhSX7scZf3JoIHrw8L84aLZNMGEQXOfty4FAFf8vWO3e
sDXL8Ne2MP9vzDEjOl6bPxAiyfSwRtBh1ZGULfsffz4hjrW6w711hnvwLvTX9xRG
kOM3Qo7BOb/Eo6FIIg5adCxYEgOfeUu5Iu0WX96SPO8RaFmKF+TKqs9oFJUFlqvL
/O5xsUrDr3Fzn3PNFruNCxN26hupwXxSSYTQJJNhWaKFoTlHxe9yGkupy4on0iN6
9Obf1hq9nrryuA9VRev01gpPeXMidx1Y7+ckaFcZuOQmTI2dCxXxUDrmiXQzhFyh
pi/E0qtwBpZIAeWQHxWisCv6WF6zgCxOSRGgDYP/O/d+Qi6CUVbaD5x98k6CYktv
m7kgNhVJBwxYfJFAzHHsNXtDj27WpLUb6M+JXyCX2m/C3913I8PiTBF5PloXkF+X
CqoweFgDZjPMRx8+w5k7IyfjhkdF7FMp4h0V1MU3TWCKiRRP+fqVl1Nn01/QkCwq
5/zGiPxD90MjXvFbsK+q1r75ngbG0chZkuLekk1zKLKCHN+pg7VWi1JNM4tCCV0p
cC8OqxVPiVenDTGmA1Jl8NrlRy0PvWPwdFxXvK9yVFYYRJrzxSkQuM5pPUvH4m/B
8ry/CmK/dG3bLKhOxEeNLitpHQcbRC1LmwM2n/5nqwItwd2Yj59zZjIy4hZBt74o
dLFTaRgTpTvfMkLc+w8R/L5Lnw1sZBrtA54S8r1hHmlBwJ62/PeDe+Ex86Me8XUQ
U5uhCQJwIxcdfCz4+omLn7qM00ZK+arrNcj3q3HWYtbk96AtQ6KLNjhwgQmZvr16
O+dDHIX1O7xyYlT70TO1hZTsNqNhpbirvdCCSVhobTaeNkm4JW806hYqLvBgH28K
aeYHl1faYnP+9aU5ECaPMEjZ8TA4MVZ0YxgI9mE5xPGDkvKaxbT0dc8A9VbE7cAP
hTsHOvA8lZMfsJAQdG51+WXIlYxAdLFsOuYIaSPuZHCqyUjzNrh9s0ADQfBP+J+V
xhRFTG7pKn5hzmE4YSH8bkxdT53gaxzMCf7lfYj1ELp2w4QbEH99g15qWqNJvS54
psrQj4CofLdmfU4J56csB/aDfTWWNrfDwwnm31K4uhlaoD8I4WiUokolgXsKaIHj
mW4cujgHSmfVwobMbUKB/EpXT3Idd1m1nzKJOk+MDSPNBt7zoxX2WBMGskFLA3Yg
Ee/jd4fBdvwWYr2CWSwtGCabjfR6GWYfcLAhHljO5GklnYJBGzpxreGFFy00gEsU
ldaqzwcAGa1DQO6E9Ikp+F/Pz9CUgSECi7WaSx9EW/LlQpOTJhcNXYvNiE9aOwor
nkGnaU1Ab23OeMsf6MremWQYaldaKkYSZNZ8EK19rxu3A7AlL5p1aopvwuebzXc1
2jzuXzUjU6WZE81YdjfM++n/ZYfpJQnwAx+E5LyivwtyV8qnDVumZDEBkqoUU8iy
o8pFkpXYpEKl2CdLyyz2cZuv5ULf7twPr8qu1P5klrtvTZKcfu/fGHQQK86MZ/fJ
wjX+o3D2GQyqNFiOBMO7t3WMU8USa9CNBLlv1HoqO4l034c0mcbD64u5kyn6WmP8
qMhsJGJl2SiPMvNXzIQOMUvrOnPX8wVaFpksZrKXLhdLNzJkc7/g6c6w9iwE7lns
0s8NpYhQWiaNL4iL/2S99R30X4yy/uZFMz5LHjqe/0IWiVFIam3KodVu8hAJMH7K
Z3Ni+UQr65FTBRoxPA1CwhQRCS2KONcjvZzXlYQUoKbv/qv/EBmcJ06MITEu8isV
gTGiDcFwxgnSmUb+ig0h9lpPCZRsz6tG4WHBooBy7dFsDJlRnkt2V314rvgWtWvO
aOWmFT22bqEzXeIF/OYgQRWQuDzppaQ3D3oQdfd8LMOXYNYPMV9CpWB8i4n0A5Hi
iEk6cIsIhcY9wgHh0Zv9oqbVlp9R8wzkzBlwD7yBFQlkuBCDgtlY+mNXTGTMgA5Z
ECqiEPVOQ5zE/PkHWdpJjq4G2VCqBYctXmNMx1bQdXvWL0jkdVaMvaUVO0iLs5DC
9JU/+scZFGdzPZxwK62P7dmEXSPHTTgBfkNXvv5mNX9SB1qd3/QoAs+w0kiBGYll
G2nQDiFejWB3DwK9kVOvYGdR6ubnp1DivvWZOOljeobjX4PYRHjpJ9MohJOpSQ8m
bOig0nHFHv1d45GFfkqJpl8nSjugkNmFd/+Csg5HlK+wwkUSuFRfml1ABFxFzO1Q
UVGg+FqrMvxvrOzU+Up5PdBV9Us9VvOy/rjnbzro6jyS3Qsk1PRWLQJu8X2X0mE+
PC3awJm7CEsDB+bByZqALGcf2n1Ytv+0amju0YdhM9i9kSJp2bTOZUzv1f+1mVWY
RDfHuu4u2hJNIJPnMQRlo9pweQb9qkhyZJG/o0H0ARY9o3Nvl+WUeglCJ+2nAUjT
dsOkC/MaMmrNl3capOnGAGbeNYG/ChP/Z4os8aDSCYADd38KxUF4co7JgmuoK0dK
ZvCMBJB/kGJfpZ8FBSDvTA7F+atlgd3A+g5lJmbFNeUEp1IFnBNgp5Q5BW2IoJit
2I6g/DNVJG7d6XG9hfWtEC38mxVpWS3KdWqcvPIRbBfoDOpHm0pXKZUu9Hrcs+I/
hhahK/G+3iPTadTNSHTPaK9ZhqC2nM4HTR5o9dguqmkXJ/bbVnUOcb2vlxN0vZPT
jSOLb8+2lKTRPFxIguBzsbNgwr2n7pNGXi1v12//YKgdZBQ8/1HYzrBxTARP80Vz
GwdtivPmHlUuvvsziRi0sm9CalYxyDNqmhsf1RwkdUu0EOn2x9xZzLyxRqOSJReC
x/S0bJNmNCUG9IGtIfdg9LncS2EJ6yEp0ctpr0GtLP1i/4AMsi7mmUwuSWjPeMgq
atX1OC8HHVbWEbJRtFU6cmQuFOIBC54di8M78X437eygwZL+XUVbguq1JAI7kE5p
PwfZxbiaZu9IM86c9zje1oCuuOn/9TGULTohYJDy6HLXS4+BoOfC3vGSjx7jGAnW
vkCKuzx9LJ9C4ACqdfaYnnkgtxxmQj6KY/k8M5obxW/m8PKY3Hf1b+Xys3oyokRZ
MIcyMUp4+v6JTwUwVmu0mZH/sial/x+rPHula2k3DS9vC1naNvI7RdlzbVdxZ8W5
xehrVrwEIsLyjujWpgilY1jFE33paC47Kj5ghxXb+GzV3uyLpnBoDXI9daCrL4L7
iNWk3uZfwtOAHrLwJUs3PkLvjELFwEbTmc+hpVj2vYgEEpyu0IUMXyko57ifG+tK
2pM2XU1gMF+wxyi5xC82IO++yKMdqKsEf4aFIw9TEJ/0fpXyArxiDsZ+Dt01rAXb
3t4KSq8dK25/oU/ouPOfzi/AY5es8VtxJ1E+j+QwDoUS47SbTSOS6ANkYC69YOm+
9YxAUIRk2e0PngLr/QyQfXUeYffi2nxVhm2nod1GjLWJi+ckyu9UBvqiyhsJcSrJ
ZMf9kFABxWsmstcYwdEWR+hIjf3SK43GQ10K/T5I79bMqiRBejxkG7RIJ7+9yB9k
c8+A8lZ5u/+5m/GgdPDUlsKHgpUd65kP/Lwc9Nl9P2bdqNELHMA1G8eynSxXaKEF
ASNQIw7dqDBi2S9ss3NYDrGySk0PjaR87mqjne1+O+6z++61U693SRBObCU0Yqf0
FIBlvGlAVMRb8KURjPme5TmFBj2Y/sHUrBxgEFJEqo4gNV1YTDvuRvz2m8VvvSpE
6jSfy7sVaIEBScnxMcq33B52i2hLeAaPvqG7UuttKDN0/ISYV1m9xMCaYpR5I3zB
P9A4H4eh/RQhx6SEWypq03IDJVsIunEQF2RKsJgfcx5mYLZlmCWK2xTBEWIOZStN
Q2ib7jzaq4NPs5xr/rg+nr4pOdBkrZb6r7mtKdIxi2USrAy7om4EjzntuyQrdVkn
nd7m5RkdvgIeDvDRqZam9dvw/Ti0MsyDgyiJQCYhqGrNt9tLPlj23KUxwou0QMjz
4bXHrkSE2Xp4T+ZREal1rI29wRBKWS5HlA3Xg/pqtxc5NXU6RjK5nmvTIs5OFmYb
D62ZPBkHI4VF1f9a9yaBL7RV3MkMooRw4l8AX9sryH9Lx9ObSRIqW5qMfRW9LmNB
0Y9cpzpW4SpaCh/xR9gOVB93VgOQrCfwxTyMrVHdoQiSXRUP9C833MnxLTRLnJTk
V60FpLXbCb6LG3uZeAD4xRnsp087tEbW+uQE8LKulEueU3jIgLh1K9u6vArsQ4D7
5AD9TkKODvMSh3+g3BdYoxMzl6vLSb6cHSW8t8wSeg5jYM35ykDpb888WVJp89cQ
iEXB374w0rYA4UtTcpQK98kFoKj9KmM7mNGviaK/OL+oO/l3q83eAB0Ur57HaWaA
2M6U/FWrmItA6HYYlAIA82adXzM2Izt1eq6iL5NBSqd4sX+szxhAHsJBCbKiGav3
rlEkFior26cyraMrbKRFIm2gxYUF+1ZVMVyVOTaNEYaZcGPebjH5RqYAHFBsqP2q
BxIvMxTtBPNnrWNNMTlhmL1KSdUKmpSYErAShs9bJWeY1AQ+s3Kfl1pQ0ikvdyHH
VdNZZK1Ubz374FfAN/8bumxJ8IsXdAKDpMewm+oOqM5lgrHf8Mszd2fE3ly/xdWT
o7QM/tKd8fAWBZbJx2+QzFCmwHWFp3uQTFjw8OBr97kezvkoQbPE6KCE/5LSYENs
EO9ihEyXWLNPQcQMPGFxsuj3wXkGHlbsWOa2VNwDF31XijEbIwr6ywwC7RozjIzh
fNB7MxFpA5ul8jo4+P+NvcpkDqGW3K50lRWDYsgfCzjmAmtADkKXSbz6LFXNw9rH
0F+Egeqi2XFbeHtHYzMnFVEgoJS9Y7aSNnnvY8lCeTBoT9LH+EB77/rHqULFZvp4
mccJS6B6v5kPflMEMlP9DfjXZmnjzqXRnKQ02p2vakLXYMrPhF8HdOw/6L/dZgDE
B2wxCtvXn9qNkEDCc98/MhWTfWkbn4aalJgBotAO6Gdt4VYbqgjggnTykQPnn/dM
dgc9T0eiSLjfiHm2y/7uW4B5aKJKBJTUO5g4YTqUhMi9zuCaK+OlYgO70Z5WLJtU
t2oGF6RuKsDCQkoyrj5/64ZNXSLAh3NwWoxZ/hlxDWBbzvb7W/lgWKixyVqd/dsQ
eI10LaXY6tQmkDvfCE8XsCULwITWzz/YViJnoUS1U4THpekPiW6K/rz1yYuTA0HO
pEaYBqJRh82/7oyzNwTzsQ8niotAGqU7wxpr7qckifl+MJz7m+PG1s2qGdomx2Wp
fUu14jJQkvl9z0Rl4B0jPawfp8BMuVmoC7ZEWS1MqA36arwN2nv3CAFsLouTxXBz
9BFGjTmaEQWUCgva6KiuVlLf5Cj17Acgwr9vq3P5ADZgS2rUk62Quo8kUHZJmxcR
L9DCIPqlpeKJD+8jD2LF7ewkpp8Lqx6IW6FAO3yY77s3l7lL87iDJ/tlFp/fbCSf
DcLWyPW9fC+7Iz5dreorLz2uzZ8nObxzvOMn+OycYT+iST5C0fm2xm1NCDOT442d
LZIL4cjM34aEdUoupnOFnnEmSWYE3U2Mi93aBsqVs/9KFwmTGqCOVSpTfGtEsubA
37gIHkakXfRUvIgYyGzHzuH4Ux5jyrhm4Oze5uQ1lmU5ujg3NvewbXvdoGFxbTaL
ZP7i9iKv83MM3musPppfblHQ1ghGyjszdQy+W3dJshAY+lrJY/L468vPMdVBdCKp
KWuMX4PYAx9kc1qD7Tq/jxB+MRsTBcgxTqJM4h8asEIqVkzyfhbZD/ZISTpNutNf
pi3DMqrh8jsIG36KgEhsPTRv0uPblI5zO7eZbP+JDYTxuMugFvTCVrlXfNq+EJlh
bIwM23o3F3PndXgGMsQSXHSXdi8vacHR9oMtB8yXhvP3yvFwNTwXr0r7LWnjoVKK
BUU+PNmziaLgN+u9/RqBTZ1lOzF4C9FPrByGDd2bUSszUqP17/nkrj21BXmS9PdD
k6537JyuQ5zjK26Y1Od82YvGph+/P8qLR51Xnll77kOKF1CoClIYEgmhGGdcbevU
qOBQkIuwoAI5yG0+160KF4KvlDIWxX/d8wmq43hJkces5JzSvFgL9m8/+/1skQ1k
UYnaUJPaowsrb4GFgM3UEtafk7+lhHwQWxaKSfNvIhTUSii5mlAFi77HBwfSMN42
q/1ftiTdJlm4aVJfNjorGqN+mslCVDKbRFdenmLFflrhtD4dS9dj1Er2HoVuLWCK
CNoe3xMdwVGG4t6E8X4lNyuXhGxr7dHqLUhj25Eo6QQkYODLfFRMSojhCuuKvUSn
RuGZLMLzWo+gtGjTCROP2uobEZS8/7uyB7lk27JhKw8raKurQKlyGm0cg4VAo6tG
FcHFxIuJRZS7voFkzzqG46Bmln5TIDX8nzQaXtW/xdEpVP94Kic16xnCfFOHkd3Z
WuTwPvNdFcRzHALZEb8YQkdfs5fgumha1k4R+YGHcUo/NF6d0buY/537skjaXg2r
vPcQXtAACti7aLtZewChUOyMevWnw7DR+a4MTIrN5LgjLDnZ54Xrc6Ijy3h2PZoD
SjOk5o1U3d/HRMCnxGnEMsSr1AqSDqxYcJVkCyRYSF9KTAtq64Xd5G0xCsxnZNko
1vi+w2U81aUewuab/WbMUuFpi7PfLFpbhOKHnc3pd6Nanyr60aBgSxIpY5iK7NgO
KUHMmiAjdA1pWIXzPsaJ/GpR4MncIWvd3dDXAmFnsJXCkMXp83iV1MBjAVTDWhpd
iHEagJMfGnqa0yw8WBGggCYUG6EQPZgdJgN52mUk5vXgm+LndhL4ny/+LdEhCIW2
1ZVxme0Y5BiQVf1zKxxNKOKqwKk2lm45VNuMdoylm8gxulSagrPerWr/Jb4aSnfl
d53C5KZO2njHZcJQCDPoDzmdrxifQLSd9CBWl3Md5sgdaG013+Kf/ni2hX9d1V41
MKQO75wSHR0D6W8JhXxs25Xy18AWDY9gpa8iKoGSb9s44800ZYKdpYdqi4MYS2zI
hoG4rpjdJCsNwwJPXEAXasFl2lfjwiNwtuFMsMAaT2A/2Q1zuwK25FJnzKhoTdS+
ajRlQ1HwEL2Xw99CJczBvc18uG8/Chr8kTBezzgBxgy8fQQFWCX0INZC6LbD+S+m
wxECsNuLsvj8OiaOEocG2obDLL0+McNF0UV8bZmT7jYb3YRS11G57ei2GsANsid2
sbcmPZTGymYseZFCdh+YzFcwuzkOHl1TwQqmSNlGJ5f2UiUl7xNU8+F0K1ZCUnyl
MuY1ChHBaJohT9LO/X2raR/kGz9MxsV+yTh32ZOC837CYdv8M5f8uXtP6FxUYtgh
Ba1tZZiR1hsZlloVjq5RhKnBTjtul/AaW+rLzakU4L4O2AgqeqUZLpGsM2LkTBP2
unxVSX+zd2DwuUFYldKAH4gNKJFr8xk0ZDiE45VNrlF06DMr1947U7KLrVb5Dhar
FgRPi05yrMwQVfIpuGY6mIADwlKi1C38nwF0oDqtbh4GnkjA8z5iDRPTrwVGK9dX
l8VvQ2IN1RXFPwFu+8KQbWmeqqsZ5RMN5tQConYOU5ibVWxdT9zin0qfwSGAm3Wj
eJwbeKlodhPGiVLGFwc61lStnmE3OZONNBOpzmaK8wya2mtnVN2vbIlj8Faofgql
XGcgQ1vsZuTGHfoHk8r6qHcjmtdOjrTFKvBwoNPgQQnHCHF4A+ZVwlOqxy55a5/F
RXoeDaveOGg+tK6nlFu9GJYUD7+Ht80LtaSASv8LrdjA3G8/A1Y1dKHT9c2RpnI7
WjeaJJ+jWnb1VtPlxTscFP26B83yZ98FQR3SJHCJPNxyGsAB1XEmIyrLn2rD5KQz
hbw+M1wD3EtVZOO0Fe5RfM+NcqdBU3iIeo0f8Z935zRJyd6h5wdF5ozeOL6wVI84
SVDSLfr7NFd4j7U2hcfrcDBI57bqfI/L0vZK0RqNE5j2KuQRaUpemBr1wWDSMFah
znFP93qYCAm3a7R7pZBeJ842tMmqsh2PtmqRXAdj/3XOEOob2zhQDhRcArrPCu2w
hIOuZ63exac0Vd2X0ox78DTNO+5AAmrPhe/+QHp/BpUFzjh3wy69OWJZJiTzUHqZ
hNHtYtkRkiEEObwuhrLfDKrqAfKnJhjC86L9Mfgyp2o5pJ2f/ksrlkT4ymVxLoND
CXhjPt3MbJ+qP5USZkMN6ksy0LmDT1be1sCYhOp//oVJ5EDQWqKakdkNV5/Tdf5G
0c5F4zAB/2p4UZBJWdiW4aoq2dGmCDUt+QXPg+0+yPhMHVc4hFxqd6482qx+TOwX
wNj2Z2Q8Va3nUehsggUXGpj7AOtcWxf/9B12zH7YAWCtSiT3qbloU8Rmpsu9htS1
foGXlyZkKLNWhamGHPqhGtUBxBiDi8KOANC3J6+7en5+S6mFLWuoYpRqPtAcQzYp
SO+XO2U6D9c8v53aWhZtCWkj2R6hSTXLnulEKB6cc6vRetv6Qw6QVOxGfRllprLI
pZLicy9n55wkrDazDX3WomgMCLLmwoQcNSQL6+qzuwtm80hAfMjyLJnv0oHImXuK
bJdJih4BFWI3WWZnd76wtepydiLi98M/W33wnqxDttR3bxctQsTl2lfYqN0Tkzx2
ebMwS9bUInS4sWCLVVvwgIZzBnsBJIrR7erjPJq21vf87X+w7WblYgB987MuTrj0
0B8KEMI3fkzEGQjJOufLftTJqACHrVKkil9tvkdOto4NP3iB7Evzv+9rhEf4m+4z
+p+f/RNxoGbCqcGza9azkaH40JQwQqtwXgdgSpfD/5QyE/cD45tqZAcM0hckdu+5
L6GqhU/gvMPo4HoDr+HS4HvEa9YlDGGwRDiWq2h0bS+fdOqNl3l8WhE1O+5EK9+Q
AgwIp3bknosYGxwg+CaAvQo5ybIQdPgEkRGiSIDwm0lzxKDFtf7uZrbsGtSx4n8n
qkkPzRCPKvE8/aAR8CDtKki+cHL4NNOu2SpSde5W+Lz9oQz5NCoW3x9RaSy+sbdD
Mp3tjv4jGCV9wU8xtSzZLam9nTsC93B2SGHb3TD6797aFgBBepnqT5HIZYzQHeSw
VZ7dwkvotQrBHb2AEgxy0lM1KQZ+fvG993/EnZLszCCmFkrLbC2PeGeZxgRrOwH0
UrqQR73Lh/+8Ees7ncJdqg1MyIYu9wI8yCiWjGZMGHiwMa/eC2+jDQHSu4uAIIaV
8/H+IPJFKufq9CSlz7No0Y5jkAigdAXw6fILCWVYpZDvXWYyyL1P5XPD884gIvJZ
5ut95VMZTGhw0b9FfeSHc3Do/qyV0/q8h2e40Bd73XrSvPtFa3hjGfJyz5855B/I
VG1GegFbhDR3u0e4nQeoCjuVsz7s1awkUnWPYFFil6AP3SH1AaEgd5s/Ga/kay34
jo8XcFynydrZayx3XT0tLn4yH32ggORF7lfWBJfoIKscjShtHXfk73t/2UYxDCPh
FvQjd2zbi444PgXsIDRoU01q0FQ4OBzFmsYeExxYIYTwNn7vLwSwa44ew985CXRb
PfgrEu6n8nAkDGyoUsFcyEoae/yogMDgXgKCzoZauwG8+YmWYZLl/P7zO/CABEDH
UfDM3jDdR/MCO67BZUcjt6PM1lTVIs8aMRWwnHy+rmTvbGk4sXYoxK+w5Sy34G4W
po4TSAE15W6xQ6+LF9rgs5Doq1shg1IImk/A8k6GnAGSItiw8Uy2s7JIsIkRUXla
xBdLeBh0GkoF3xyGhy4N19+4Q95HaZPEZCt3IM5krT1DJcLqiB0mBLjY6vALS4KQ
RwEDr5NKE2MJzDIQE+X6teaCbaaPhDsjRU57m+iTPTyhasxwCKBI+aKKJkLsRDSf
c18c4+IU6vDn3ctt9Qq6a+/jivbsZwtFeXyjZL6AknXEQNXqWN+mJC5Qp4Djk7uY
J4aEoXHljV/rbRDgH/FvJ0gsUoJBxskSWksVTSzMmqmQBqFGxMjiF89UFNsMmXQy
oXXHEQrONTDeLkNbZYaOpXJpVGEi3H7x99YfPP6eT3yOHDIXTxVf3FGuTNB+nORw
fXDc9kmI7wWRyKmhkQFXpUEtkNDwC1SK27bnj120YxKTySeGM90r1cWkBlSaPpz9
FOezSgxEe2eGaA3zLxEw0G9w+WUZ1VxRR0ZwoVb2WfWq0YvnPzx+PWAi7dMDyKKK
YDbjjqnlQdeU9CPFXkm2KnCpZGP0aO9S+nwjNYFcqec3c1o0p59DcRVFA/Jl7AmD
UcChbhV3jUCe35MeRWE0eA0kfLV/PJzNYL2GzvqGoq2I5gGNTpL8vdVf2QNAfrA6
dY3ZXJ2j3ln/DxqU1pwTINkT2KCWu5qOdNbaCeP7zvftQqh/VizHOb3ykdW3BUtW
sT+Fmm53LhXTjm+0yimhGIQ32oHAxDwc5kHPa4e12Yt6QVzqZxCP55Y8GVSDoMw1
DLR5gqe3kriITCJlFt+tklVxubgU53WahGDnYnawPNQCq95AAAzQGIklSMJJUHuw
997E5poXcZCo/WDglx71ZbnlE5+sUzLreqd4DBvE7wvU4FQq/jvEOwY8mQZNTSav
AC8ixEN+gNV1+jzjePo3dGtZ+gOewjQ9cwyhSOB1MqeS7NswOJYFqvEX2TcNhsj+
x/0WjBt60RupmAyevJoigMHt+D9ABdgNspwZdgeK6OdxbMAuUF5QfEhea3nYjPAt
ZTbyr9uYc3VY+uTuhQa9uJLIxe1Gd+SfLsk5DdgtBfsNNe+DQ30gbhih6pGcj895
niqOBxdBnj5EuTsEI19XHmqvDuHP2F7pJVMBSjOwrZOmfVZSBlrpmMTd4u4NNkRN
kR9lelCROxetGNLobNMy5Q3p6MUAq+2X2rhc7y19DL6ZAxcxsxgrJqc74YgdVYtS
BxICeygDBqSSP2RWMTfpi++i+d0NR+w/hu5H523J0zjm9tLzXTOPS8Z48N+cEeSb
Cb7QUj0FW6gIDEX37IRlkTX23UGuFRJeFv7WHk8Pq5hFvXDobLggIIAf6pFtwQrd
0d+6eSx6yi1EW9Mxp/vCFClnDG2wAfv7/ZVkCU0Weu/mlKfNsK8CirF4Lutc8EqL
2EatdnsSoL23ltisFuy+rZMX82QoJHUJpt5ohcxAZnN3Umd1gJTmSM2h5E882IHc
n1KKY272UJgPs65Vu3tvFqMPzKzb+6hzgqFdfg7ZcklxlgyxJ011fraLY6kf/xSI
YBmirhqNQXVJ64nq2dycWzkLJTuOjeq+oolk0hIFTOWqrbmGmljBl/LmjfUj60GG
/B2QbzJgO+r+62V1jZ5mpx/4PN13m6ar3pR8Mk8MsRQpIPiWNjp6i7HsaOhkGCHu
eKR0nllCBfaJkqb8+4e5mqzXPY/GCODhyya38t5I7FhB6UvywSzVOxQx1NlG6dKh
gLQl6CN136VWSSthMJYF0lhgFFU3WGHAAPUC04cvyvu918v2Yl2ENEqDcuLmGWY5
GYm0mKII6yD2e0EDzDTkGoYzHeWmsZ0eKOwCzqpa5e2a/y0wG75vHia0OUSedqOT
bUSFp0E6McVtq1gNLXXaY+O++y226VT6U6YLYhPwcU2A4kAg+Fkx9zPuPcT1Mbl4
0a04EB1Ma412mp5ARiEVOHnt66775/7CFC9OqxkCV9G3GaJmWrK1+wtRQUSrUyc9
8tz2ZcqaBT7s93ng1yc+hdm+tTUZqCFFAs6JN27E3n3zY5nSIvB45f9Brtm9Y7NF
XOAQp3xsFAwGPzyo6sUrErZfOOhHwNsX4ZjMATJ12KGi56PRovs81A7Xk81ZOWkC
7rvAuX4PUePzhR6B/o8u3vVscW6NYGg+B0YK89PqgGAXK5eQF2beD68yrwjjL7pj
4V0cnX0BI330y5xE7/a75nhiWw+gwt5adBkcaIsb8FK7dp2k6I4I5LEWm0OUZWZr
mPipcdu6MpJiCyQeduwT+5sEcL0unP1r6hNzoMFRhnWkvk1+uwyJTIr7P+UffuHX
cGrJsymfnAbNxRsyAaI0SBwwgDNmJcpO8OQGRWssaPxRyZnFAPizBcv0wo2MnK0n
IVXLqKq/lvn6LhbBlrRtzgZRzogCJ+dFwwBJlAPhAeyqXJy61ogvnVU2SH+ayGyN
HXP2ZE9vQBpe8O9uUdN5uufG48zIygT+q1e3XuHL5kULLiq5c/KI9OtFGoROGhnK
GKwJmyUyb6+h154Qt482At4tDkIVyOW3SBLQXnedcOfVlQTNItZBpFIjpboTRGz/
dAahhSVg5BEZkXFRbrZjpH2cthX4NB2LPHA/JqwJhieYW5mvhTlVfsb1a2ur1K1m
SebWpTDeS0pgqTkN3uZQuV212e/uPCpmjtB3PJS4Os4lv2JTtmxOdprBf+QxBcoL
ExYy1U2nyZtAwmVzPexC12Vq0loDxarrpHV7Ht3V1GgXWLEIluwLccTgwW3Mkpua
8Xwq6ogH78YXYPynxhue7HFY+saVqnU/KWSiXbxzSAwFfkNRXtu7qgmLlqUcAx4i
tpUcDEgdz6arY4dSSME0kuMlamq9ce2bbvphdBsaKJgNVwLqeSsJyXUz88dClC2A
4g1ssHNMw5pst2bpQsYByF4X20jA3gaxDCF7LI45tIopb9ft8USgemTblDc+WPG3
5IbMK2e4VE4GNv5BHsY6yz3nQZOt+wQF10ejHVvTqaWqJ50CGR5/6rSoXbrhPJJE
Je1aqGEgyEMAJjNpXMwIyA89yyk6IWeOD15M8WurCT5w5DdlZaJCF2j9oMaTDF58
3E7x/N1UE0Y3n7//+LXUzcJPU46loekOW1pUoJPqrEL+eWPIpGfWT1TkrHK6urES
yWdQWKuF1/ExhDtFc54zALHost4bqFY9L5ToxkVGSCaAA4S02ssl6Z7/Ttl0DspV
H4LV+iP7bUfsMCFQkMpFwYoXq16ETphEfNtSvob8suMr2oyWsjaaipaO7VLbLUEO
ERK+NerWJV0ZcoX80HrENjqKViOHfAXPOt5BhlcVlb+CMn9nGWLvGEAMgCn5w5xg
zojetY5nDomGcHJkJAXpTNs5vjgHiHMoWa1hJOm1P5OcfjpjEik5MMBeByktZi8m
6TXnuLm64CxUNI6eTHKvZ9+coAU89AqK+qps0v1k2dDm+VT8FI8axeNAd6RmVlht
jvqaZdXRTF2ntHL3HnbWEkdDkNs29lTR4K7aBq6v/ZTybur2AWhhe2xO0o3jKck/
AwIViLyU29ne6PwFM0GaEy5ZrpUvjpDfEAsiQQhXJ33qaxAW+kuC0QoJr9c+hccX
TZRu5VVplWc3abF/NaKrDAQoEtq19rX5Iyoj5Imq0TjGPwSYrRl6TR55uzO7oFdQ
pWjg1CfpcU0GxqCraL0s1CLTH5a2pNLCA6Iga6aDQejYTcDygMQJoqa9SLEw1E/s
DgaYEr4/Xf0Eat3/iYJY7aPViPwvLRIFTOPWqWA/rrkBAzuAfjTDBXyePnjVBTpN
/ED+4LwF+4IGuBu9mD1bg9LfnxdUSGCWe0u51ygCWlEPJ7MOBkaBDJBCqJLQzk9q
wPxRmWNdstZHteIfn7mDxD9dTdWomXAVYQ97FxL9G7brIIecBMKYiF8mx79+M9dY
8qnwW8t+y9w9X1WMx8PfysWqaVmKdIy/nRIpQtUVOsl7/PtsfYKaOdx99Kg4XrPP
FJIejrFoGKhBUumy3ISvX/yo1dqnI40LqkiFhbCPcSE2p9N6U0t/qtvyLWVFZKVi
XAMw4WuTSgIMXImEtzpEwDk83I61CtiXoRXRIu9+leFzRnNQlzWLDWc9EwqixgwM
K+WBjFvdbitdF/DRF571joNEA6rAIa4ISXex3b0843vU9lLRaoLEb797/VUMm9NP
rCf5Mh8YCcT7BGDEPnQViZo+cDJJ4mm/JYBTcUnUfO9cc+UhA5E9LAFBLZ3Ir555
C7UyqNY85Baf5hketceRGZ6kxdrhoc5SlOFOW0muwIkS3SobPWsxqlXCVXVyZzgd
utT7x+PsmZ5RPYg7ACSH693fHZmdHbtTsGXdaRXUCNG2+kvrM2gWCfuAOu9cmWv/
TRYANyqHXOoYPo3B7OkApnKrbFXsjKc1gZevHjQ6WPjCog6uzLhUZ8cGvamBH69x
hxPkais3pziAqpfvtzNtToJI0kU8MwKPOvm4259Khx+U4Dsx6UxgXpb5zKPjwA0R
Q03rhoGZVQ8uqoMqM28vI6xE+WF/CF6Sx+6ql4If+uhE61uSmKglVF5SdPuaggFQ
fyS1/0/g5qyJHOgxO10WkanifaIYffTr2pQDAuZ3TU7dQ0CDLIa46MPpSqVGkBfR
yQMWZdZdDMrdM5z5GIVnKIhkyhihvfje9ol+gXLBAq0ZG3cNuktwZdRAVSy1zOUr
qAv55cw+3AFo9aqcRV3Hg8hcQYh+HkAJQy5Mu3AtqsrXDNAX7kaP+xAUknySuS8B
AUs2L4PGXUvM1qjb+Q//h733cKeOBqriD++nGK6JBqY3ZrT2MXg+0dTcxAaSurBB
/Ie6RGeAD7Y0RAx8cruSQHX6Z/84YbsMqFzcueG5DDhZm19L/U8h/z+2gKVkDBNB
oV3vZqtnofxBZ7lDHoGJ8zyphC/7Brp+xZtTEJ20IjD45Sv4AQBzvvf9sC/Uv4UM
IvyPYcb9cG9TxQfOCzJ4O6gJCpNj3JiLeuFI+YLFJMv1q5omG6F9bnZa2CqUXYBE
QKz6yifMBxZi0gk3VqTJhMtp37fuKey58L3VLUmC9O5g8WdIECA8ZdbYxHIywp3i
Pkptd3BdDCw9IYoModZuHQPIkLz5ja1NolWgs0HObjOi+sFVbDxKUYtXfOGZw4O3
Ft2OYSjKW/TfPJIAYGozs5AIE5M03MqElIS2tom9rFebL1vs+F72rvTLcaqsIkUP
geuRT/wnEvTv5RBbuIo5itBAxRFYIdpY79ictzSzhVWVVcCy2Jn7HE1L2CgCBNqg
4tlwOC9L9QLXOsYpjd+354tnmKRWMgTfeq8y47s2anqZkfCt2jz1roHeDxeRYQc5
HxtkbrAcRvegV4Yqe/eYJStZ5hriRshIuqTnNzU1tKAQeckVV/FN+HlhiRmc9lvv
gt6GP8R5N/4zaSVe6i2we4jmiY5q2OXKohNkr1U7u86pmhj1/PqrDiSAP2e2QR2k
FbTw3PgZFH+6BUmwmNU89JRjKLIsuUJKOwNl01V8HZt5szuOJwqpQ386tUkNsPWt
I6Nxxl4hyxgoR4vFYII4mBFWrdCxnLeE0v8ttTZqFu/+pJlPya7rZn4rkw2mE4yY
34DCYvGA9Yq5i76pZu5maX4BV2cjfrMnCKKTTOBUNFX1naRoka9EDW++7CcW372i
5FroyKm+HD0Mdid3Jmmm/FofKcY4h0m1vdJb60+Tn2DLMDQux7MnP9bAfw9TmxS7
joXJS1KnKt7NFX3yh5opn8jt4WaaA3f2LzFZN2oGcpTwFYAdtEFffe2O2zdEoi87
+GwHjRaaxBseB5e1mjYe8SUsFNtSPkpHHh2huQEABLLgVYNWT70DflEmhjzd6HYA
rCZoNlnQoTTjqlPqavkatsNnOXSIHGwt4FObLRQW8QbrHWCJU4Q9Uhr7s6R76hDR
TplGjniNkVcd3Zj0S4f1fYivK6Q+xPkNrAu4OAbur6emTEAq8qNrpzzMMKx6faL0
NNwSHh7qf8OJSVZ3UD8ogJO8jkdC5MS1ZGIVWwrRgfvz5y8ts54zWsJBgZjLKIPO
MzfMc4dIRQh+cUnbBOJYaconqXEA8BmVO29RMBecHAxkpNgh+/2NZ2+DlzFy1KkG
sJNkYAlWS0VnnfuC77l8rXPKRua0KzUxeS9bqdnGS8iLggNmHxEtaww7oVSaefIq
JD+N1mmCaAMXfLtR7v6g3C7HvUZx2CRAMntWdacbxyfd5RIFvYfS34/hGlpq3F6o
4X6YYi/R4Rd+q3AmfmpmboKKRiNwR1MBbAQu7L8mC8EGakLeezA0n5RRwbJz+0OC
dSvaZpdOZQAHjchbnCJlrM8YClz+ffFDY9bKHYMY7FmEKgo2w8dLk9yOPgPyOMm5
7nt07FNoNpiIMjrU9wbrTIo5Pkfn1OY+KEq3tNtkFBtDA4zcZuLFENbTWNKa5OnS
kp5RjmdD1gVqnai3HmjpXsVUh8s//ks7nYq/NRr4F8ajs4HERwQeZDG+TYrPc7PT
LTFcF0kvnt359oDMWhJR5rM0PPaSoHz/+IcPzmmESc/waA+UTQmY/ORRAbVnSi0q
4mePnIbr5gYzLcBhIQsEAynXi6WKutAVdi2pK9Z9yY0FKSddcZYCMwffPxmxua4F
RiTScFOMvih3/Hg/uAQRqu7S4alA9h8pQzhnhMe5d9bF2uOKcgHXHRV+vXdQ3Q8K
LyS2tN0NWdnwLunxpxJPNOW3X9HtsKYyESf/mHdv2s+aeyuS/6wGBvFILkAXj0S6
maZZwnI2RfhCHgXE2oF7vKiw/Y1iVlNk4XZ2NjpoOEmycGwHU4HdeqvcNaqpHavY
9I3OIsFK4nG3oUsq9ur0w+dlJ7Rg3SsLhy/6TpscdZ7sdf32hiliX+7Dm6UM46dP
hHaZE1dXE/EBKBlTZM9QDw4VAADDk/BugEU1DlYnviiyoFcOtkL/+KWVHAOav7DT
t3RnHm2MugdqK9qA7BIdHA8C6D0j5E+Piks3dHggFgVFEbCHeyoLeiCVnE4s9Nrt
Z+HmhBqj3ti8qcdMqSDMLOUymlVQgk3FuzinxB+Hdds3o7A+ljX4U/bmB08x9j78
uY68Ms7GQR5CHY+L2ww8D/3DHSldz507bpu8m835f3M3aOWk1Id7M5wHHod+OCbh
8nm+ewp/dDhynlidpz8a7b+ZLU3qyWAdZxmeW0Koz0swDY5Osvrb6aDmBHIStXlB
xb59ZcX3/2Giz93nGDy6XobN/Pu5TGHguCZvfKRzEwULvk862xlVSwcuKlxGx3FW
Lmntm0A5IeXRGo0bUgfc8nrwTCtkM5AVksBUqEUTyHUbCCu3o/2O3EwcZPgTAoRw
R5I4cdF9kY5D/CkEdxLf6lq+08o0qYiYlJnMLFfexDuuolS0PCTWKI5FlegClUaQ
io2DM4pM1hDFl3BsAFs21kmZw1WuqVC/LDNwi2WLXEtft5n2QVoR20H+olnfhUNX
7UiEdX/sIlts/nyDf0xK251G+QJFqAGqArcZ6Q3uga+Q8JFqHol39E0NeNRQ6i75
58YHjaFPPinXKwzTcBTjB+nSYbsSt3VrC5aOdHxjqKbfRrIupbs2g9n+NIxCoTs2
3I2nTQzF7EhH1gJFBWxeRI4XkYYe00uupYEqCeA4EodgCTgiJWYHa4V0YS80Llr2
mRWmrzls4Nn1EKXKf0yh1f5gYsMW2mKIJ1IV5JCei4843JWjAxL01xkKuNKlmrEs
6vA6b3Im5p3GWqYSEnTWplkwgM+S1aILkq/Z+v3fM1Gx/GUGYImn0tiphCzJPlx8
ZpM8Cve96nPmCuiHvNjXKIz/kb4hbgPFf3A/SdtTbG9HaK7VUOQ0pzuaQvk2sMLi
ewylB8nU16BOT6g+WYYGLvr7MZJravhVRgM9HcxdEd/vGR3F/vf73/R1YCJNLQua
aBfUgbJQT2/kBsNlV+kyfQr589vnwoK05ITKsmEfzTZ5N9xUowe/IBmoob3VzNlX
IMaagVX+fy15u0jJOyx7pqWnLkWQFDXwNqalYmKMtzsPujkwYW1STNkMMyoes+GA
geV/RB9wF0nEGgGtuhI0htdno6RRWge2JRJfTRcTFVAB6YymtSfN+yTq2JcBe14I
XyyfHo+NTtuizHcuScoVxjE/+Qs48K6ZcMf+wYBaY0ee6YEm38xBiKEWgmqz3TIZ
YnYGJCmvjqvwgBw29fseQykkO8oWUZGKNwqYSA5JODYrRH/NKP2u8aN+GcjHnLwM
ZbYzXgNDQwZeAmLu+sQ8PfGACoSBsiHjLWfOr54Fhv8xlEYJD2seB6Aqvxwk/wWy
xYqfw6b3sOmVaWnk52gAQgCLj3/KiE4bX+mLqypQaStnPdRvhT1MMg86P0AgSJwt
pSuFaUQu1fF8+rbVELLvGW/2IVYEbR9GOsmkhr3HNSindfL32d21eph6EtPxK1sh
IYj8ozws+MnliVjbEetLsGPGexDB+DpOfO5/vahON+IqxZHjFH6Mke+OlVOyPb+W
BwGnZ8Dc0Etl04nOWioCHDiZFyQTDxKLx/L6iHt/8s5ZwcvphO6Xya8sHI3BXf/N
uhX50OBUu/rG/vg4k8ypLxieLDqngOIpilC2iuROTDVh47OMEyD7qmUj5guJVMuA
OBcUlxCFI8uWVzGc+t7n8uWmUAtHv6fHdn6Q/5OwhOoRGkQ5DicX2xU3Hf6JmMgO
PDQiORTh06tWpBFrhqj4/eYMZgLiq8o+Y5wkrkZO8sp0NtOOLpzcFol0eT9mrH/1
0vVzfnxKU4rs61ntnDjVsaIKKI1zenxJ7bc5Z5og58G0i/d6mCeURgMEgyYIz8eQ
Z9P6LJoc0djTJEUBGBSOX/ln3ET6q+a8ESohJzgvgBvLfMoawqWzhBVR1oNkKysr
BqtRzlw+9qUqNIMTmsopNfULqlU28/phPL4oYtD57c9QXS5PsDFJ72pMhcjPADZc
BtfLHKFno4F4yhiyXrjGrNzevT1qMtEUhLA5BMyCjLu+NilqmH3nnso4dQujk3u/
YsE7o0UuNyAHeyRLUcfk5oY1+qXoSx2uvrkzT7EPtQrvc5IWJXytMOIAQLN9tow/
fghPhDpv+KfKC3n2kJJzsHWWUNC5lVP/5kp9aT6RSC2Tzyicl4U9rvFb1ylRuG9U
7OsbBNICA2UUdv3fALASJbtOLm1UAoTgGqRqHveSKmklqshKkEP/f3f/LyHAqVeY
iDGaOfaTY8A+7R/FjRnzHml5cidVQh9qZNs1/ySN08/vvY2Q/jbIdDB/cyZtCAyd
eHWWbbbKfdBkXzHBWoK/+QNHjuyhiDbZpOlhkVhfcWin6HnfeX5Rh9JJ2WwXfOh/
Ba27Tx1Q18OqtiNTD4iSFIs7zUbn7UyAWm8lhUFs1xfGGpZuxTg2KNBrZZRxL1CS
QVyxnZgq/z0EvUGRfvyydnGIWcuL1Z/qLHmZm7aFl1mMRT2w/dvfttoaOxLIHfAt
CXYcBd85L8/AbOR3VTrcZJA/+hb+wSAINI4vOTPojeX9yhlRKicx0qiCFz6GWjWB
jtJTVqToyjXBPI+SFVAWkiHIikpUDFpi3b56RfwhJ3lZgCpXh2YI6fbJ3JHC7OkZ
NS3VB371Sl7SQWPxCDATplYNrAsgEG2l45/bXuDNvvZX07kGlnAxBnIkuWV5AJU2
wy7kuKnjEs5vyxdLg0zp4uXROQitO+DG5w72j+/1YB1NpsjknPFzFKgolDvROpFY
ht9dUdkKPLCXigk62f3OiPsv5BamqfCI2yqO/QbmQwf8F4w+GDM6VXjPo7YyPOGs
vAfk56D00HdgcccDcr/8RZFxn8wqxN346Hx7AKRlMZX8jV5Pyar4hR1R6pEYKqwA
71fWhm45zSHAY/QQ/7G+DcfMBJhBpwKb/GYvckRQiMtr+P0X/G+xSduM1MFF22nJ
EO5HU/l00HcE/AE5+Y59XFfVWJCFSIiq+CCEO2hb/astkGUK3xV/7G9VHVS8WDOh
f+FMvNz8fGvnCH1oGbS3i2eLliJ1bPqhk0nqqSP336yDorYxob0BrU10WJkSM2xD
f1tszRTUeavcwPyJnW1Gi2cTWRhiByHuRLZv9Slfzz4QgK2PXBwl9kf9NilclCAZ
pV4fT+GpY4clgn7LseXxjJGWCEnPd8/M6knbpka0vbiKX28uUP2E8bOPJVQd+Hto
gi27/7hrmy7wtLxtnZAGkYF8Cd8D0wPJCQ9HzQJ4bG5+KwGhoZNl8mZg+LV3+hFa
/BUn52xmPFTXuapAT0KGnSR/Eu1rgTj1bJcAjA7ZYW5zm+X13z2ejSPmg9UFaaOB
mjct5Wm/1ejW173jZhpzczPJv6KnhsnZpkyRiaP3YgpSYcYoa9OMLD6CLmNH0EvD
5cH6b+ZTb2ZRRcQC1MD9E96pmMhYpBEamZ7FECCBujYgqr1onwgtgZ5vXhXSQDxa
oynT93vRJl9g7BfNGWo4PjA+D7qb5jC4DgjVtKZccR0QjwLGcfq2vBg3h6EQTRaz
OMqcPptdbGanx8Jfz5CtynryBquPUmgsfMF7gO/Lpx/+NvqOkQzdtsZE92AXbbiN
beOR8B9TBRUKFJbj8bVFiighQDg6sV6uHYTg21ow6k1dyhRkv+m0Rt/dKGaDq0lg
fXiKGG82VtwF+w2DdaBG0qAoU2Ly8GE2qrlTx0/wEN5W6u4sMmHRDEVTKoRIwcyQ
s27+rcfpPbecw7KKRk1Mj87GMvfa1/3wT363g92Z3auJDqfJazAVdWSvjZWxYeJS
MjA8XhSaVFk0ihDHaRTdc0vIAZ+Lh32O7+WJ3oBApED4xIrJeA+fGSwkbQvdvDo/
cO2igMko7FgDfhLxRiZ2N/yJplBgy36jIFMtZoj5hLVIrwadppjf+iNKoxMH9fjR
wWLeHAcf5GISavQetP7eXZEdSWlap59qTs/W9xm+ah8Lcqj5qtKtJn4zbI8AFTOu
NSxbSKfIv14mZ+hiQU+70p+Vbj4fl7om6a/f+S6zM+JEBEl57i1zoUHgG3keemiR
P5f0EWsXnST2mcxafWNIYSE9o08U38DG7CgUq+UQVhDNcdOuojj76xGVlrciJexv
m4c6ASmjbsoSjD7aq85nnsFclfXarij5GO3YyvA6rSU1wuITL+A+JnRruGPuiRXB
L+EbVG5Ki9fo4Slm9pnuaTonbyEUqj0VkG+6URx11iApsJBuKO8NBr9C5abLY2pl
B77HqiHgYwkj9E5vyp4HdjkLIuOG/rE5VeGUX2zlARukzXBldx4iIhgv1f0ZtknM
vhFjIRvkaJUimmVE0GC12UK78GFdQMVNHmUuCl2PIsdat3KjrHT95ky+wwzxcKIx
bcB1LFU+Db+9BB4Tr99gm8QBUjfrN5KcSqSVSp31CdIfNOFwCHZXN4bB7eG/AACz
zpUPoaJP3As527zDzF0Xy7YhcVZCIzAwtoX47btKEaKCLT4cKwCG4whyldQZYokI
k9Wy34+JdKrrgYk3hdh/XuU4FTGDflW/ODJEAdP0kQJYLTwgQ0TDXlzeMjNRuAya
uNh0us5lg6sI0S2gT+PqqCvnpLWgFG3zeCO7I35ciEr9oJAi0IlNTst7BIDlY09L
pjdjaveLY/IBYZRjI223aUHY4D4tX5zPHXnczHr4Pu5XdzAFoP3nnpmkDpeAiqO4
rKzBzcyQ40ueP1hewZNWZ3fSMf22W8owiUJVE9USTF+bXyLoicY6+3pLY3uoeHz9
EIUOo820DIYFh9A731QjZwQQAmeKb1KhwW39l4T5DTx/UGJbLWP8iTx9K2Nx6E5W
OVaYOrlehqxUNv59XNmoAhIdbMNeLZzYXrW2abbGr72ZnamoyXTimukxbJu5E25F
qxT+pZ6CDdlAEhmt+WRzubpx+Y0BBi57F9mkkECHPJeYuhz66t94vMy8WfZV8KsQ
BVTpZbuza3gBytXQ0V6kQXWXVphi+oOgvLidytOvElXztEiW/14UvHbiFFyZarWY
y3OSIwDanpmGvHBDXXmN6ywOfsjk64zWrpHrdMhk7+2IQ1o3XOQCSUFO+LHWRg3x
CgqRapDGstyPOOYY2ljOd+g6B7aCsLWkN9i1WyaoDBK/awuL07XQuDgafGdY2woS
kAG1KduyNOdCknQiHNZN4Jv1wntYKk7Ns+rO37TyfiTZJWk/SS+oNY17zKQvS4g3
ary5ofKJCkDezieKq4h1vF25BwrBE6aEHIJ+JP3vAzz6iMQdYprIITQqJ/+SZZk8
`protect end_protected