<<<<<<< HEAD:flexrio_deps/PkgChinchConfig.vhd
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9056 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
qe1+t0GXQ5YjcbQQEHGgOR9sOTPrYkMBDTKWYPscHh+5P2Yop+NzK/fj9bW9omQ9
cpdu06V+ZsCE8RyykpTb9GrAIX8CLQas9b/q+yP2KwM/3RJZPQlTOsnX9q2NCSRS
sjxEf0Wa0LR8XcfkmjT0xQfW6KkoN73ksDOflPpNN9j2TyYZtdKoR2CydfduLxyj
La6wLYUBnGotiDbQuzyZCLh64d6sNBVlk0wt0Mp2gzFLW/TNQoyUI10oA21ShhV+
Iir2ByMszYNwEWXRPUgRkFanxs4/5RyeRWGz6T+O2prRQf1+lWPh/eqBQMmAnVeK
Rd+EqG52Z2+mjjX1BKatcHqn+LB/1Cu3kOljfWKHBAZOHZ9+OdrL0iQTrMTJS3nJ
NBfe47leQG6yQXCxlDcB0vILATxU2Es1Bs9gyVv7xfJw7z2gbRspYZ0ahhqKu6bt
gO9usoNvbLvTcAkd7F3iPuVf2qjwDlqcOKbY2ratRwETAAuSn0/WdpgpynwfEM03
+o5stbbRd4khYDxmLluwfLdiVIjANUD5NeYYuwPcdl+M/VhLtrhDvQ1yA7fdzHy7
TY/3oUc3/SuI29Tk/oopoiVYcgZuVWS1FUNdRJhom307SJQfBDyFTADhjT0FrGGw
YKsWp0LxSd8FKUEhauJH3HP/dHac+JDPJ+5DOGmvWRAnNWtx10vxHIfeXNXVVYJX
LNpmG5OncsY0cWoUmuZ1LTi8OwsnFLocWczwPtdh5gr/vBzgpc2ast35b+Fqx5rm
tGBDbuN3nZKvjUsBWcjfRtFle2HEnR1va4xtgZ/SBqw8VB6E4BvxBNcHZ37Hagn2
xNqfO+IYnRgJd5IxGLJGvjrk7AF+p3sx+IhBA8dqNL8iZBGm35hXNmSR8gQS9Alr
l6T/GHQqpWdRhSPdWVhGgH4PxKxrze3tPQr7azEF/+G+6wZ6wdjyAFA/E2YfKuwY
Vzi52+r/G0gkD5J9UQImMwMf0Bbcb4wa2sQyM2pNaegI6ar2z2lddKQB8YRLIdQe
VEcxjPc/Mx0xQmmrfKJUaA9A/6F7RDfbtY5CcptQMKOhSLfrLYVNGRy9PjFeyF6W
PR9ejIniwU8CR8VPl514uZqva5k/YPYC/PjANLX0fkN4L3Ab3ZpOepX8f0Fh/nmf
4EgaK7U1MR9oXs3GZCDrwV/Ai5t0V3oFqlP6Ij2Zl+OG93zaeC1u3FXDgj2e6Pun
WwEru+ktq/ejDj+Oxbz77uc/ku3BjzwcSurSdaJXXxwi0b2s0Gkzh+mrwUZLNnpw
/C+iV4dv3Ha2XYIyDz8KNe5jSc3K5Ls8R4CZ5lnjflVloIjDI0L/km2M+Dxhzevt
QFThWOpZHL1PgETrs2sTu5G85ppWQ0x6VAXG4VL7vhkjgJyRQHAe8lKkTHNtxiGK
SrQCAZmEZevU/JUpN/92iNKkcfQBkrXkYVwRb3leNyC7h1blvKruak9iAtOj82n5
zdxXVeWa4ByY279Vuu7FnLU/7/8dBLPZ4PlqZxg1YG5pHQVcWoOY5nDgA2rnr3DW
qBdVCVobl7Wcav9adwWlms2d2DYkCYT9TinwEl80lGk1P4flEG+CgeWnbksHYMYv
UOIurg+HrROM40tYbdsuX3F/n21tuGjELW5ZmU6n6h94GVZIhfgR40gc0ve1P2ZN
pHHz6kCt7qIqM2KsUI0vh6ALHwGoZXOmzjyosnV17mdE7f9XMwopiS2TIDKr8Wjt
AchC4rdIzHh8/L/RUkQhCyYcwFCwsSwLvE8J3gx3V2Xt0JB7TokR/9gVLCrKZ4FS
z07iPk+yZm9HgZZbq12HWK64uz5QgZOQ+eME0B6PzgVtqzpGoKfS0tM+xehxzyRl
gqURBRlBl6uFEdt4yqnaEWsE4cyCccU1O8ThtGfJbd9XpxKe2zcvS4TAtSOMmBFu
OSxfY1hFL1Fwh8PoI/u3tqFiqaj1+29H0LX/VrJqY2aOUMP8BINZTXF9rk3JH+7m
Wg2AagC/VUvYSGPQGuR0nu3P3IQwWs15FvKdMnDQx7CwUJY3b3iLoizcwJByOLv5
JszRO0/JcP1rB+YLm9jpBo+FzeIFT7dyKZv0EhCJ7zw7h4AT2hFF9audI2aruq1J
yohFnoRwG1LkGRGF43P8i4dwCT0xArGsVWKKePgLosLslOmo6hxstf1lKCg1Oqaj
povWoCh++MihNnaXwOx7/J/DEaIiKQGYKfFEtBePKZ3r7JwFQXu2Q+KNqtS5veeL
4c/rCK4WYRBXCcpIbkXR7Gu+CAaa+U86JsFMg3TA+k4IkIhltj591D+RWAw57kbf
fB2/tP9o9QdYpZZTlFDxei+K61DTm6h+6Ce1PkJfFrBhGk4Qtc8ApsVqswoPWSVD
guqgM+DRYUEc9zFbgf4VRwA14FWhMiJx4C2yxrWVsKKg8A7gqHBVXwdqWLKKnlT6
+P1S6GyIX6UwRMcBmJiIiWYl5SmL0ZyaBGiTS853QmnbULu4QFnE8vhwYz5ZVoe8
F28Hfaa6ci7RJXogjiGj0pubqZvZLTxx8pKPm3QkBBt8hXCQLgwfskHZ9r/7xncV
fltT29w9G54oO/HFD8C7RYa9wWfYPyoqUT4WxmFJk1yxxv9urWATCbGJ2mmDWMGQ
Cd8xNoPsqUzo8wOOlBAQMwnwOp0eYpZbztyJOhrSNNCJt4bqIFJUPBluYZl6eRmu
Mv9GAeaApaaoThoQVgfrtT3K7NyLQhT1qG0WDJ8kEvCkRLrujQYzt1Dn7rUKa0+4
IjCssoKSaiwg7cG1nsvrCHOrozI3IXia0jLCtEOLN9zIoaOtNXd0IpY1rc2YShU6
KNVIHwly9Tq3y0uG7J78cs+prdlD3S6VfnseG5TIUZtnJ57Bb97BTL2ckAiWWSDa
d6bIDhJV15mwJXLhHE9MJVZ6DhsQI4QGFSg+T3dxVKm6vZZp4JrOZi9n2xzVogPZ
CiQ4hCWiMDqZuRkSamPQcCTiGd3bayp4rLNziANCeJ/+/P5oAaYLoYueThDoKXp/
F0sF519huT9Vrk5sa1cmqaDgr3DTU+T9mTHqmmFItckDiHrIvJe87LLtT416kEBa
htx3kF2MaCV6jMb4rxiLW9JBrri4shu1POnGtol7OP3WuDVF265nz0iDC3c1ofaP
VtZvHLhrF+CPKq5wEsV3khPN3fFUgAn/XeYYJaYctV6W4O47SCC5aM2eKgvMoBPJ
yZX+Cn5E5VO9UzXV/Ncc2Lhbjpw+FZHNVNW4U0u7/iOW+k+Osf4EzpgWir/Gqocf
VCq/2SH0NXOGUjpjD/m11Bbj+BEzcY00YgkElCQXyxz9PrlZvNAtkjdk+djOM2xe
meQWcyHagq+QleipJvVereB/n+yvIg+oL4Vevm3Hij5A306OF7qiz068S1Gbf1EK
ydJAQpwyGPUPXDf0SscurDWpkCkFf0rhFAzGyoOIaIRyzoRPlpU6EBe3pcfK5vq/
3+uR6B1qjbMRr+wVG4s904KurOh1I8xaYPtduEmnnJuIQ6bPJvaoQtXqTQNrV2iy
RaTnTkKfeQno56eTRYEZVXtbWaw6jQq/1RdD2zdO1v8wjJKMHHjDywgj7UBJwSaT
rzcoDc/QfG4iKpD0kYBVc8i1pl1ufcZtrYqeLa8m5rmrXnd/SEc64YNF8Sg4IOJm
BcmEAGgysBlv89rL5mdReHHvxSGT5kQlcnxLsaMFXaoJw3bT8+4AC6fFXEUbmqr0
G43i6K4GJmVwJGmL9p5Z9M6wt12t7vZRCNROdlEh/5sEusL/EUdPMERs1RoEvQsY
oz+FolmSxdHEgbeEXP3meOf0iafmNIsuqp/2lQLKpn+wU0b9ocjg6G3CYLitSATF
TbWVxxoXH/Z+9BrFKOnWl0q7QubyRn6mZXwAZMFQesEQwgyoHIVK8aqJkvvW2OUO
GHS8ZHVnJfMyMEvoqCcpFDT9ev1FQrpmEFQzfXXNM8wcidxp9FcMvgoPeGHpKQvY
pmYQCkd7IRgz14I79tVdxPDfXZucg38aYw7BXYHpBE3TXvEVBlEKUY3HtWTnAW+9
0rHosy+SLTatyDx4AvD9gc/rwzuTj2nMeEvZgAeARGotPk6/h24RGiHa5uztVU3R
GrAqgRFRs9Wj9nJyShNDJzAWfGwcRcmOWuqp6wpmCh/CEFhExXFV7P8u1Gv8NSo8
br1iGvgWXTd8KiIXnaYROLJIrnNM4pxSO7FF7ntHCu6ns3EcBMz6yv1SOZv4jjZb
hDTbWWAgk18B8QkWcqALPP28V/zWPoahvaA6hw0AtsLie9xk97a+JrznRYgEWaHw
vEM8dAnz3RFRLHj6pYviiCBoWtpm9HmBzqckbtlsjg/FK9s5QpPidd5Hp3nBY5Fv
sse8rpVOsKMIIdwJFVxiuD2W76N7P5uAtgTcx30XyvYcnnTPZHUxk22xWgMcpSqe
fh+F4V0arbmZZcOrkguSAUzxjNMWgsyTiCl00GLmvb7AjPrEoBuX2ENB/M/7zNh8
rytJhmFlhYgw6LmorNzHyVDTemCa27hKdUwnFDXAKpgPM8OVMgenglrtbz1fRAq8
5kjltpfMy7MOmqaLuOwt16fmNEUwfp2hnSKSJO3QSr0TXIOeZ02FikqSdxqTzXtA
4oiAXxj0yN6b5TiyiszTJYDCh4/uVSL2sw8FvC+lBuMRRRGMrvfKHpBE3bd3BpoA
eaviyLrWAruFoOYnVbh/Z1hb03SjzxLM5sYFGNDqb8VTOq83WGXOCfKq0MI/mmJZ
ikRzBes8bk+8XILSxk1lCIH7EL4/+Ml4wwtRiB/OAZumaDHjQzyxaP8e6SjiL+to
qtOHRQOftYBEaT25X6rnNHA+PWHcBI6Xx8dYl060T9znU9nDQ8DY2VmKczPlV0Pv
pH8TyPyRvFmInnr89z9RIPSxazLhxBEcaN6dPmURbs/EU6i4ECF6NkI2Y11KnQkC
ihJHaPYjYJ7y+E8b5agI9xxQWZo6PIHfJHyTYpkFmuRhk0DCw2y/7OxWz7NEwwB8
a5awAKojQzkhVYPHKsirddkvpxCo2nOFbMIjMSNLIHxCBxNt9LasiE2N7renMld0
Id6hvcg9SV0AE2ey3izwz0Q6Fzq4JARh6Mb0l+i/6S/XM0Wr/9IWY5KlUVKeXj5+
htd4KAFVQNdxnfLUBUGX0WLToyCkWskKNC8J25+58VLhKp8g5JxVo7qP4g1UrIGZ
cemq95WUM5vIOusLQ1w0zRcXGNxSoaSYAjbJRzbjtsZ4htOeS9vD7p+x1Jz0y3wx
ZIfwTaY8zoP2vsiME4ZyNf7ACZ1I9SmHxu19p6hvCxueheE+NK9ppQw1wrbBpEfi
iRM6w3i4bwgzL4S5uDQVyWkTLGqowPPHGXIF9AtXLfOiCZ7x5rO4JzlOofyaJlik
qoRyr6KCyCaGRvpdQrMpcjAAN5zJhPGRj0IWSoI1xkH3xVJBWjkcHN8CMqUAp50v
2teENdKJ6pbimSguRCA/A2Pb7tCMpNiGmIy5rMEAs5kSIv1TRapWkitnBIlgJdqO
2cO8EHqUQrOZUmHi6P/RMAnKtv2IFq7WtkJMWNXbtszFL6sMqSznv0kra10Yzsr+
jRBFEKAD33QIrHVQh9jPa+ZYvAdWJN6wE8fRsCFvTG/DCBG03q51vBea08/adpGh
o2HuXMXFGE/UmzpZUxRk8Qs53vpogNS1haOeVedeymxeuFb9t89cTxESTIke80rF
FPkemxwGGzC8Jh6ARa6XcVTQNAOxCYfaOwi4xdK27QBNQDC1jb7rf7rCQJ2b6M+g
n4VlrNlrF6aqAWPk1VFUg+kA+BviwJnry8ki/cGnW7Bc7ASBujdSi9vncg0kGONB
00V2lG4/EOmzcKikZjkTkEtAxX6pgL7xgymJvU4hN7kFngEZpcZP0+jlhbRJVObr
SQF0UzltAP5bQT5tFrY4dlGx5QzvxMT3WGXMAXFOsyrhfhVoyhNHhXUpxMqc2y00
WM4Li/psXtk3JqYYXxUjH4fbUBA7FS1dmD7Oday9Mryy1GDmLWmGuOdY6InY/BvW
nsIaRT4NQQfQ5dmTq2VB3IRDp0rm1Tiz2OEFjN5UO9/Sm47c/EBkzc4IGVI3uZvn
AilC37uVVJM+rQCFWAIVpFa2mlpovPRaxR0aeskz/hMEvl6kEClUUYj8FS3SJ/vi
Xe0RU78EgdAr7CPF+JTM4x7jcmRS7vPXkAnPDBgtlmGIw4LLSRGxvoiU8niel4b/
YXRAxGN7j1rkX/7L1IOkLmZEDV5paNMDjI0F9zhpN0Fd0HyyriTI8eOcBZR93CQa
c2iFiWVMfqZSUCotnAYDW2esdHVkQ6iY5lWdU9XBsKKnqK9kUF1drOaUflcu67Yr
zEmlijN5AhKEOLicT/Em6UuNHOtXiog+9SdoXsSd6v1gSTQ7kcCy+awmPIpp1J/N
Xr6Lnz/36o0VC9vhJS7xQPsuWpO3yqH1+ytd39m3zPaV38UIqEt2yzo/FIsWwVNr
oSQmUgSGWz+fE5FBhANNFclMy/8LG1LdAizGIcQSHmz0hgcO7fseTTh/4PdKFW2q
Xh2gKEXbC3G8zTRmA0qMpjAcHWU6OdmEPk8i3Jm6qTLIrb0+ZGNYz29r4Wt+QRgm
MNOqpc0s+pbE7iwENKb+9ifuQ9b3VdIz4EyNVVg1ix+9Fgm1kyGa1IkKT9tvqw+6
J17PEkhG3gvUfe+icx9LH3RcD0D77MZN2quEyNa1nXYh8j/ivhFqm/eSHrQ8RsXi
IQkA7NpneK6qIaMTmTcLgDnbk1ahFlrxVpwAUCxKTYNAiKXqLoebjSpuEpElNjNx
zZBNsvT/O93NFE6REt/Nn/8fpCptHXJNOu6u0RcOsKyKBRXs0cr8Itwee4uulSVX
HaxyAEus0JJEIm/YM8YI7PZOE7Ni8vAJBEsJmkTWQNLZYPm5zIp5vMd+oue6or7A
2EUefvFSALI569jOO1mh/giGA4ZTBQ1fzZJSmk9nzhwLqUQO+YEr6seF40ZPEe2G
CJQxgMXlFNPNTW1wqFss/GuxiUXXQT33o1ZliSce5OhuFB6GzobLmg6UmjW2/gUu
h2tL0rJwPOc1Ud7Lg4RTxw/x+eyzNuAuVfp8lGK9i/1uJx5iEf0xCTkCGXaGqqXC
laMdIu23J/LsO72AZBE4prZM9b3pYsXvvufc+8cZwRpVMFk884hM6tBI/gVrSnCZ
ed5d6dJzFp1hTLpBYh7NbD+nuhrblhmTBCMJqesgVLszowTSfU/vs3L3Bx/w/yyG
iII6fE4svA+o3esKNd6rDTd7/mzGgTsp004RniB3DThkkY1We6C4rYtE/zJKel00
JWuLYu7Jg7es8Sm68TMJDd2ZcnLIWqO60Ouix4P8FHRqbUqSCJ8JikQlMfcU+KyV
EqnY+I/qV7qD6qlExTtmY9z9mpI2Px6bw6atz9rVL+R8MzVy3ebDLaYleLiOQjZ0
nTQAN9mNp8F0V/AlqLL2z7FVh0riqWEQ8MY5LHumJjKiMIWvj2Wfbw1C1KaezATF
tEtZoRr8NXoIAE6sCXwhxvhGsfW0HNDR0TY+nTHsw7B/Un1DOeZOQQMVxPtQqfCa
NPIb9WKzCHaUAfXdSGdVdMkO9SRq4DICAyKuSdxI+cfgzC7+8mhnR5ozxtaTHocU
vW4+tC8QJzY6DscreExOATTi8mT3w1PAiKA8j9bhXJVi7BNszgeubq+BJStvBKXb
7+9vX+Fp4dp0rqdcKfEA9klSJO/w9UxerKjkFzBptcMAbc5QNx2kkoIOFUsyw1Kp
miDQdRLlGR4WUAZqj7xE4rszAwDNaBBtXOMdXz18TJocgsYfANZ5+OZYJ/qNiV1s
oHM01WKA7/xlw6Vm3mUDB+gCXJl8fIfT48utcMuwhQNP1g6eZA0BoPtY2QL8Jd79
d4GGDTzmDeAb7g6FS54ofyViknbWxm2c/4OBZcNjDUMdHI6er5krE8JJbC/QZfkg
W4EAi4STgNSKH4RKpn1ZwgKa+MmaIiUHxiOYgsMfbgDclAYOIV3uB1FT/q9IH8TS
gKraYGu93PzzvU23iubAiJHv89PCgiL9I0C/WB6lJisBzw2/zHnqm3QfAmAmnSs4
lZeWaNG3YBzNUIU6pXbEqHTRfecPRbm2HplRc4PGRvEG6qonFfyMnPv5h9btvp1Z
9T10pmDjkx0IxHdnPaHP9JpQiIP8n4n/SVRBxNx3oNMLbeAMcrepYnBV24BECBVW
YEC2eOhkl5jNBhN2mG6ky0C4eMg9hz75qO+ZteF+tcKL4pE5elgTD17Z5I5u1/wv
ta0a43BjRv7rvQCheRgjZqi1ifPu71T8jDPRYEr99IoBpf39QgENbh3es5WyD1Vo
UB94TJ4OPPTnl7pGt2FqM4fEtpnXnymG2F6lM8Co7e15mkXW0dvpI3UQS/PwCeQ3
BHRzAcEeLBvS3ZXYIhQqYHAxBtq+5NZ9TuycU2EdLQekTIHDHt1xZ5nyYymZCILU
NqRDp835wlHJUvEp/I294wMKslGN4aNBQ00H+8soQLTM1GtnLRO65FOPjNxr2kqL
qoz8vrdGYjB+Gtcv4E6x1G4OOzpBoWWzHCr3HxoQTBlm5UbGxOv3yEjBGJ1Pj3fF
2S4c31H59wbUfvAa6MD5YtF2ZEgl295gcGoId2V9PN3HLUCM4PGfHltNrl3CMr1J
5DXsfsCSBR3Kss5BfXrb6rbeQIXdt2KKRp9GDAl0UBBEqc1Kpsjr56/B7kMhJ7JN
aGT6Mdv1EYt/Cl7I2zAnbhUuSgaoLcNKLnOo7fytenIjwMvgs/hH67jgBywHdVCf
+x9Mt4eGqGwpE0zqRajEe+E7bHJg8j+HDvxpWz5H09qcP3V7N2utTDNxSYQHlPne
GQJ5Nbxa6njpq83PehiB7J4teN5bUiqBCQJpLUrQeFkMTrP4M6Rhsx+uhWOQKiz9
8a4gBPbWxDnv0hmrsECtjFd+p5OknNrhKykySxbEQpEjacrxp/R12qN7z5W9nF1m
oedFUnJ/QNKnKlLpksWEIgESJlmYEE3POzxU2zSxIAux/ndcVa/ScmwLUuhrcGPA
z7UyBt9cI0U8T1YTdQ9NOC1KjTueOiLinYtW0a5EO1AYxCBlPenK2sYkkLfwWFQO
hNgZ0nzPn79YS9q1NxnryDbiXIh4ncMPU8vvf/7Pt2vQXkVAB9j5/ormX+Xx57w9
AZvADd8UYv5XC78mB2p6180ES/m12d8x3r66D9aC/YG6j+jgnDsjFSDvOU1TusXt
mzK+VXjfgj/6TTV6x1s7qxpu+ZemdnhZnV+jWwy8LJuRIDarQNjcUtKbCO6o0lXd
mcb2Dnhhd20klThsz9IAEHe9TdfL8ObdgdKjrmo465gHz3u81uTbOd++9CfJPMhq
DpTDr4HNkVHLnOQIDo2mr2vXG0B+QTQiRaHt5sV0KORsiNzm0ivPbLAsx/pwTU2X
qfMQtBXxvFgmRqJILTB3fvUUq6ySjjIT0oSO2OPJco/phrQrHYwxqYrM9AUQW6Sz
c9htt5HVNyUcsAunyfz1rAeSl7G2CiyfGLgd8DhHDwcFzQVQ/a+WvZ1IgfdYfMil
Vd4NZcA4bymL40BmYmwT3coVlCPLe6cUg9G6lsE3ddIMwzG68U3fucuQLP1WN+sV
LvwpN+811fWoUPIi2BjQv+c9+/Aen6rBwcEJ0EwgojZK8JgeGvEZylm8GaE698rE
LcgxCnbjEqNFPs/ISiNM/AtFgr1cXmfLPFnBeOXiDm/z9mlGJwTCQTE0OeYKfBHm
oEcwklOknSr8x8yC+yiFepxbuiWjvUlcl6XVVpRYVq8scaeKlPXvzMoZfaj+BDP5
7TcxXeLOHX58MQswwVupXRS/56aev+Yfn8QJRtzkac9Dxt1s79Q/luIghZxQgDVT
wkkgoxT3lcT6XvK5pf0ifUVNjefImTvBoS65FQsGgXJAyl9dJjGgTtSjDucQdFWG
wdsF6dMubfqjkt/OXD6LzEHoBYdBhagZQRJlHVVaF2P0b2+sNEyfoGfYLOtNuMDF
+yx9QLQoA9btQ4G2jOz/JYcjvbsuN8G5aQFFQu66C4VeXfOXWcGbufz0C/nzkr/y
uRLecSAL+P1LYt41V83Kgzwmmb0BGmmDr74VROwvv566+pIljstF75H09rTyt2TX
i02mWKDzDJ6PN8vePWZaTQUOXCSua15/xrX2mrEVnWcFeeFHNnXDz4MVJvbnCN8V
E30tkGDIu59KCycjMDf1c35J8ILH4an/DHEbD2kcsLHombWuLp69bIkfpDNlg3rG
WhO5tfKYwLE/C35+rsnyo0BQeJgY9wrclr4SfdTEX3PB6RnWL7Cp73+8s2r+xw4X
KjjqyiVKHzWUjvXOoHm5OZOKuwve2cuivKLxBFJsfcG2NTCnAyqMUOPbeJasv/Au
dB5YoCTkZofhjK6/h5G3ktY56YsTZ+6HfAS3iArtRC18Rvcpbk2eDgGQIrdqx60b
3SSVwDby26GcnrSrciG8AzKT5/zZxbQWoqbl+QEotugxE01UjArjl6+9yszZy15+
roQiC0MwS70MLTsDlSXbeCalaJSIhvmfV+8iPc3mtEHZFtGo5SYNC/v6+UGrnzZW
1ir8uWaQAMtR0Cu4dXnfmPMeycTrAXeXt/OQ+Kg0DUu32qSeUeY3EeUgNL6fhvQn
lD0kXd4ASNJ6aAMesNf9h6eyF0mNzh3RfiLvMUjR6lWEuRokPhIVplzLlv/n/E/C
Pg+BdhB4meWac6+P+qGOZ62fD18VSKmYrwQVpI6rFZBWoG8/UEc6XiFCBZZYIePP
KwkdkqQen1jALsDjQ/aCWoNXV/imw1xH8qHrI48SFQ4gZxYP5MHdwd0++Y2rFf93
u9HWD9O0kUUR1cJu/4OrUXd8nsdpQYHdkouopaWMRPlDK1lASM4C+6UGDh8VWkY/
Ii+D//T44GN/IkC/OXlfWkYZ36tUVoQGqdRMNcEr1KnBeHWTjbrEWyTH9SaBmGow
OW8Kk4M7s58Bu5HSn82wkXq7/Up6r3zfpV04p6Jx0bAKUARY3F8DZ4BCdvFLbrug
NOU9zt5m0tAFvg575TnvR0sMaTG+8y+r7ljXD4oowrdOdtPwW0hXlx5Js7VSPNgu
tli0GECn2RsD98gXHowPGrHG8FTXmFmwUkp/e3v8oNYSz5MHarbpnw3XwHLpcgJl
wYJum12PQGLreBVnnZCz41eoNCRwzrlBP7WU3LPPR92ujBRAiNNETwKnssC41BxI
Lj5Azyx1yhsD1NzPAfJvZjpRoPk3xIVw3lBgtqlEMfC0vxNL1pzgSt0jws6757x9
jH6FpfXdSee8Kxa2CCMh2bafbt7Cicvab0HqhLyZQVaXtabF/gK/Hh79X3wUf/Yg
y8Af5zNyo7BHfBuw0R2kFdGLnREKKCotD6MrGAtbvkrGx7de6PSykNbAhVrwzNet
aLAIR2Ncz4nfddSTQxWCe1ldbiDRiwOKzfTS58N0wNv3N4uSN/YwqRAc2OVznINm
DbG9Z7arHAPRtCgMCGszWp4otwse+yuQfzlPtRbPLZ2KSWVNdBqXdG7EAbQ8ZffW
U1sH+LHrhf3u2c3ZrC6fxLZVOGYnf+vP74BIZwsF3AZiPheQtbw8BImro7lUc8Er
1ZhilE6SGRkLnMWmwAaFMvL5wVEjbUveWQiO68RmZawmZs8zsHvm3qxOcJ97d6kz
Q3v2vHmU1OJPRU8HDbzVpatlZpQ6g+6Hzem+mMiuCmDifPITD6KG3TpsJ1jDPN9+
AHOp5t5UoIHQ/uBhDQSyaL15qhTs5BKybY0MlQabV27VQtmxxA/KXlhdK8VTuOK8
UJzsG4z5aYMQfSplgTa4EJCAFLO4IfT1AyX+7kXqW440Vk30dBQO9MwRSDigtI8O
o68SR+csAn+b3IlQ9RR42zPHmOCFqykw8tpdk9SeZy/dZrLmEk/B8ZkCgUv1ew6w
Axs7mv7Y6WHz6AwZ0d+vYltnihfraPD+l79vFyXq22Y=
=======
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9056 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
7d1aayJWrMXzpB8QUg69LNkEVUTXPx2Vj/ZLgBdm96mlWsMOxKb8fHG14KP9FU0E
/W/SRAej79uWfNoQC5RoDtfFayHrgKppOSsgBGjbOTQybzeeixXH+Mv2XRMdgYoN
yroBRLluC/312VH6JJkv6OroYehie/0PAuWQeket3/E2GxL10v2XSbW5U5MlrdxT
edOlXxSaS/oS8iYoG1nZkfFDSMjH1dwZYnTFPFA1HwXuMf21McgZEWRMoLnxGHpA
MCeLY3TZG2fauQfe3wJThWj6UhipEA7Dd2LpDsWq5BiHnQ8UI5K6gBlplmT750Vi
EhuArf1i2FSSwDsFyoFbrCv07ZTAeRvZe9cDrEIblf9DhHy+/3qKD5PVMn3uKuN2
EqCZVPgwPDJAf2v8sgue45Ihb66rXdq1kp+s6O3+Tg/Sog6yb12v4yHivjzHWNEL
BMwOJPyfeB50Ilgm7XqNnuNxOum9rxEV1VG5+WNrhG1qFwdzXTwXYx8ZOahtL9/L
EBipbQVGFPe8S7U6mEG0HgdNA+5hs89AmUxccO4FWDrtybKFdVBKhdid3VpPxrnW
p7qCJzBKRASLnRvhz0qoC7BK7E/oa4YyHKq4fU+hUpGtrNE5uelP1FjNksFL0+Ii
Z9QjRV/nMcTM1z2MpqrQVCF971uAywoNBVSW7mgDBP54qM6L6Yiw4htrOLhL18CU
bFtVKDZiU+jsxSvJKT30PHQdwjtVc1qyVazwS17GgGJThFNQWSZu7XUBeOpc8klV
7KUPrht5w5co7Yuj9X41Hjhska5NXG2GHB486NnRDwxf0ZgXUiF5FMw8HoZfdHwa
EWc2X/V3ri/phzu5ovROiK3aHmcGMSwmnh6YKhgIKL+ayYGBMO9UCsyBK8xAXEm0
Mtz1XbKFdNAY4G1r5Vd6oBa1r4J5+MiWWjzTUZl6eIE7PswDWU/jaX6xavHtyE0E
HtUWlKDVxiUrOkzssIZZzig9MJGV3HVvFqq3xS8sn+c7vvzG9r1r29JjDgUj904j
jlMVbHquwMogelYAkUkEKQeVO8CHuYBCp+/f/6eQ5uhvovItexOYxFQatPfJPHm2
bdIalP9plaC/xvO9ux+q8h9cQCDCutZTblY1RecY+72qtVO8y18yIviNUr1r5aSc
ipZ7qf2f5u4snY2mH7w2hzqincxWkKC84FO4aPoMaoonohleyooFydwIhTfbs4/k
4qu3tV7IAJ0omliI36szPvREddrIJAnCKoLKwK7O3M+bdCMy0CPvISFcKJ9in4CL
HJeMVd7ndzqfdgmzPHsZF4Ny4NyNHmoeuPoclPX6zr65XtHgmItQmS4M5d0hPtA9
qAdQxgwL9FX+GegmFLQ788feDxLM4eJNhE6hCICBEGSQrJn4Ma6CObpSx+eWQoi+
3Ky3p59+QND6eJT5ls81CbbmX8WpbzkmObdedvHjBy3tzBUcwV1+xgTEB2ZeZj26
LHnELCFnXOwzP8a2afgboSSX8Dy/lfcKokSfq5dJCdEn8phSXBf61ezilGu14Jxj
ZRd7Cj6TuvHhtXHXsDytzX1bsDLsHUvGki5X+m2sTKkoX/Rr12oFJBymgElSlR71
jpPNx36LE7q//50fOJPlgAgSMayDTyoZcGeS/kM0nTfqZCO8ts1VbOqrWLocV7Jp
a5eN6Jnp8aYIbXYjBupoi2yJ8MVpGhvX7LnmHTRKuK7I1kxovxG6J5YHN2jkCAAI
42FQgLop23ElOMciBoXtcJvq2yju3afhDe1+iL/+Yq/vAR6i6t3z3yOrGPC7faTn
Twji+LMlf3ASo18iNJ4iTHIWKf129ZylXvF+KQtg1GhrCOwg2Y+S4iFlnnhnuqTj
4mNXcBXDbqWr/3BLdCU0gr9lcnVNrlGttT88G9JuUMwA4+xqjNSN4zTfSxn70NnY
I+w7ZGXR7v7B16iRPaxatalbCpDonbuqs/MLV5shKG1fpkbGbuWM/Jt9V9EXKwNB
CnlXTgOd/CfpqE0bp0Mdh878nMvwOE3US4QrygNfhpVY5Oiy63NHcD1FoWpsTlAK
RBKzT7Vl2QIiu0puaumLsBjMoBbxVrxBXsYemKD/E40bwpSLTka+3RaWNH2xbwGk
+MFA0kdfeqS8sN9bkovpFrZwk19HLBlLU5NRwqqEb8DvhG97Fj5cxmuD1oVzbTtP
OsD3bFjkSFqlFWnp01THuXD9P5DJrfAiPtI1CbYK3pVkWk/2Txg+KO/XRrQv4Kea
xGiC11PHA6OhERwtrWNIP2I+y4KLMGKh4fh2Mra/M/dr5VfYSvyyxlquQDcO4rN+
ldFkDtLIiX/3hRP4kwphemQYSNqXcniikMIL6VC66Y0BaRxFMUBK8vfuiSwb1ow+
DOIJUBYs1PrOy7Glip2g9kLhgVEFFr4aj8BEbAE69SxoMhzLkcnxGs3iuvHnYpZY
YeFtDug4OVMmysb2NP6job9FjVxaju+S2Mtkl3Zk5HaSPvPK50KIqTSEhTt+yS/L
3k/BISRmlwAgvjQtoU2Vi/b5wE2n7dlF3nd80kGSaAWY9TQyCaxBG/iP0GqbC3Wv
QNX3As1DCR5NhOTMb45Bw8uSR9HgBb19w6BR8Cr3WAl8o209xU/02dylrLG43Y63
BlNaqR4JWOF6p7f2eGz8lZkKk/y9M5Oh6ZeguHK6Ms4yjEj8mM+BfCJjnH4amKTK
3cZZ9Dxj8zrFjSIZBBC/BzygXNbAjSgXVOKAzfA/QSm2hLXY83AQbJp//VFVCEPV
9fJg7PTQa9oBCffhLHmwgCXFDMuSQLQGMbkqrlyRVnO/mxa3vpy0mmxR9kkb8zBs
4zjuEZXQifl/oSJjA2ZiRsu6uJ4m6rGfHWj937zRpayUM1S27uYsE54l1MafBty6
bzabUqPMzEbkKiSs5uaN/sDIXtmqm680wdWyrb3M7Tx85idYaa2l2xln6aekL/9q
XQAvhlFPdbswFlE3UBKkneKisWqM4xV76xfEsfBCm/Yn4oCJhT0MpmDqawjL1UII
pw2qcYwbLHSf4OifPoRUqAghQml1yY00uhiBIuWp8QBLy0Yhnm0xgo4SpDCLhHJR
fAM59VWTZpUec7zzpJ8SFuIUZxOQOtVA9JG5ULhPTMCuciO8oRjnlypLeTcyjHRC
VgUAvXxqwfv4sAQql3r6rs8r0gtdX1Qire2/F6wTV4hFqbveM2WF1PYUmiiE1ieO
ru0m6c7Jd14N+gWeU6yxqz0sYks/wCc9GazGf38A4Xjqf7reZvb7bx3rhb0FqSpl
XzUkxWWl0af0zoA3emmuZW+LcYb0cO4LRCOfAXm+DDd4i257jex/xEXZ4/ynheMv
GgoMCjwf/BKCxUPkodvq9sJ0uhup7QKktEX2K0s3GvC8X2gslTLJATkTRuwMRFe7
wpQO8vtUPlZM8JQM/fKvKugIRQLJe/OwWDsiY2aqQM6Se0FpZqh8WDbTqyKxNZ8+
vm57Es7jOOXzx/VKn+fjg3E1nD40KGoVIPw6+fY/0NI4jfALsBTGVtF91fHmW+Gj
SSuLrtyyV0CJwVv0HLlM2b9LmJCAE2iYPLb5N34NSzQUVoRdd02rIaKeFQZpJkk/
4oo68Sj79Rje+nGQq5H87ohR9bI5ThguakIpmBU+Xm8iWBbyq4DNTXEKtj2bZ7hU
3m+jGcJ7IytIf29+PB/tYr9Gt1H+V0tiy+CoTX+injkyohXEWhSq3wWJiHVQ2dsq
lFQhdP58dPI+oUSoPegmRIWwUaG3BiMsMdzBFW4g77PMqkDArC0UVaNSB+3OdKqw
AvLjCaIMC2LxhlKxApf2NmGWMWanHkaOuNz9hIJXwT2DzjDwR/beH52K8sQpvAvM
HJ8Zcs5wJWxwQi9NIVnL3kMHNZhLJZRcjuOnhDa3BH7EnetLjU4WcPgEARziKvsS
FrH2wc0Uw5JZc+LwPoOuvEHai4rX4lT3qmxjS0YY9BDCrTLjmba80DwCTAfH8JTd
wGCystHtNfivOdNY0VOayJl3W+0sREeiadlGBDrwY+j7YPae5DG/i/j8+Q+9E0Ez
/tEoij1vEUXhmAMOCP3KZgTU9QafNKGWe1sKe6M4p3e1pd3Rp4BQkqw5N+KFBK2Y
FP2u6rh9YVpvd20xHut3RRKZvm3CNdGhdGPkLK5czpXkC92naLXxZSRaPnnx6X80
jlp0kyZCd81QcPkp/iflNO+RowRNsFAXgl7Un6m1i9HSoNqN1pA1vGb5yB25zSmv
ENgOP2g0+0MoRSwEF8V76nD5zmqLog7PG1qeZWK8S/B4HweCA4eOCilbAadAql/M
wXOIH6Jenc7P7zBWno4+vqUXWrs3MyYlQ9N9O0IMjGFTKPdXEFASHthuUWaxxllE
t4/LoayzZj3TQIVUUUBmFFz0XK6aolJ3pTcHRQpNMICgjaXy6ZEbEuK/McapVOSp
8bhMfzSkRXKeaP/38DA6YHcVX2Oq4Dt1sXek2JwOiuWb6kqD7ZjnXBZXSSNSMmEv
/QPgMlwxXq9vkVKWPL9rJSqs5mmeJQ2SVFkQUwyi/YaYhhhGyyty+nxCJ5zRIm6W
lddR5nJWjJGBhTJHPdM6vwtdGX1jd8lSyMKnhl+ni3RT0kuwFaWGkHz6Zncj3PjS
Fr3jFOw1zYrrzgAHS1ld3qyQTVhYru3ZkG6HsAQqFygOJhcNGiEUM5rrTPENKk1m
3icbVgqpHvmjCtonXBNav9/xG8UlUuj8KH5NC2RtQ6W3dHSwZDNzLPiHRXzeB9oA
x8LUI+tQjDeshd4HNvYW27vsEgY11JAsc/OThioXtnKly2PS5PHj2GowJQvQ9xc2
HW44RhjFD6V+trkSgUdx0ecrqSY0TZaKfskdrnx2RnKoK+MSb1OhUvzhR5G0Kbsi
Hh/WbjCu+YB8pXp1JafyQfVa+OOR5YjU5uW2iEGQfzfjf863alvkTCmlxbW2mPid
Dbp59/XrR3MNqVGYROn23QbQB4OYcTwR24782IRBY6JjgV6r3s+UTNNTkG0FvooI
xL5te7PHcD7bIqw/7X+m9pvU+r1nUOM2AKRtesbDDgULDDB8ZbxnprKtDoti0nvM
SzinAbVfJDhmMLWu4qY/m9mLX+y1/ihXqUJvdWdY2TqUvCMrG3ez2YJVB+e104L8
VPT9ohH5yVR1t7+PhEbQkgfxl/mV/kVc2xEL0e+qvWWSHLlfen+2qhpF46/F3Hr3
PzWXw+qEADN8E79vmXRixsmFvy/810EegT4/KQE+AKJrVMA+bq4MRH1Lvfq3fsG0
kK9HWLYyPU89N5hn97krOs2bGCvvwUVeZ/+dowp0kpRZcl9DrLwDuu5N9pNI3gwK
BkiTmr+YTIZffU0DhlUS1vu9qF1yS52728gvHA3YisCzBOvk9TZX0xqtzCsLtNp6
kx0R8GPPtXltYtZgVyTvG18fcUitvKusRwh3miYWl0VSS8Pi52vFGtJBE/oAtQrp
Jm+A4XKqt5eI5XVqJgY1Ruafa1ZYP/fs3J6nu58HFfgyADH1t83cES0ja4tRVrl5
Vy5pQKa6+WqJk8gcU+vJC1ZTZJqTCskKkZBMpFuCwwXPCiyP9cW6MpFT4tlZCKht
1ED84DKFLvh/JqK2sJfPwQ8oAHoL4DM5Ku3lZCcWbP9dmSYXiQlkvQ2jc57Tvoo+
ursIXQCicas5tWavdDh/jCAr5LN3wYYh0QvK1xqqI9w6tZwDaPnHy5HvScM6vmqo
wUBBx3FvhSP1Duq+9MjlvVHN2GBLAzol9ENWQ3AWJx4rtSwCQwFauxJq8PytdWbS
1pYyaVDFbC0EUKezcFFMpyyb7vQgWtFf7Cmci+J7i+RIS5IeMBBqEtHZB5bS6G1p
urpE+abp9dTndJjWcgwE4DrrViRfqGdllOT2ChqjiOCAHQstEU28EtCOHshz6Oo3
gKdozPoOIwol3AjwqoRb9umri4ea3mLOP+Xr82mw3LCHw4l5Jfc4B9XuNEOp4rlq
p/7UW7Q7QX93wfXpgNuaNxgJZs3esgimoj/SZaDJp1am4CHvQiuYUtIDZK0PvxCL
NhLF73EnyuoKuR+NJ3K0NziuacVSsbW+xAJI7boEkYCI+nTiFwvhM2Mk+exKGAKT
9pSEZyYg+fVGJaIR2Eu9NT0kCqde7I2E5NX9049x5AkAS9gcvBGPrxVEArBarwP4
DPsJWZG1mgWmJoHeCxSIV644qfhY6HtJ5gyGcBN14yrLdIcppQHGatCrk7/mXudR
OntiirhiAS7etjWUizBcp4DZ+jCThICwzTsJAa2n2Wg756TTjH1GQ/4KkWWSDYhJ
zGcC3wDPCK4Gmy45020bh5bEQAyGFFzDOYgMBknwEljFhVL7a9IlLgCqiNufIkS9
p4TePWM9Rv35iDqk4bm1gWHgZmUEyRQOfBHDlcWF4jTBnpWsbXJhYfR27d/NP5yI
aRhURF6+b4I3YokR0haI6kqVBf5tJePeqUlcDPLgZeoNpqAxWDyifi8plPfohfmj
WggBDLaAewtivXY5USSZzjSCkntw9XYeXzRkZZ5ZgySVl9RzjUSINe6J3SVE0rWg
+21oymH5LBsHvy1SmYlgOjDieWJWlOQZ2yg4YOy9wHzNFLlPRpEe5ls8fEHVPMyL
dw7BFPaM8lXHIXBvaUl70L94XcGQDi9UkM4+T7xw4ODeJADLjWGLQC4p548Q7eVU
l6xl6pcqye2S1cs0WUAduChGMjHoCp4I9XAFMlQLZSviPrkAbk4R3dXPAy/70Ue6
7hcBSmfwCbeW4Smq30PlmY6glAP9W2+Xm0h7aK2k3lIl4KnqgMCpGE6dw0U25TZ6
pM0q8BtJ8qOBVjoywJNEgE6Mndr3u92lwdfdhmCGRZnmQSOXdmJ28natw7i8EosM
B+bjAImxVRpMtrVDKRhMt0RDNUOWBiF+9NqePVNx1GCsbzd9LzQCJKbS+pnT+MSN
ikRZoGM9RLb1XP9UyJOzd481/4u9L8t8E4Y4E3uihxIS+CVNefniAp9FApJchgBP
1WhhZVZfpER6oe3vZv9StFc8g3AJ11YLKCCMaFIK5qBaagB/iyoNlksRFytqjt1A
34GKy5zfwKOPmvsjIkpEm6VyCb2dJ5RAMnPeIRBj5jAbjLkijde79OzbMoRmz2UU
76r/R7vuscjd3Fcgnd0ablLQ6cO0BGHLjgrARUuLE1mNNyR0IfpksTNB7LScKJeU
oW6S4iEpolAZe4MMBdt9OZ6KIVfP8yaW43wyEj1pyBObQZc+r4le1shEnAv2LG/2
VCI3M/9kQ9PYmz6zaqM+PGOw6xUohiw9IdA9yy92GYlZqTtLvFppKpfTv7TVsnpf
XaBfoSbI33JtLl6SxVu3E623C0CvUa9fFw9JRxxVJI8qE2w42jPggp5Mnk/MUsjl
5zYSWjfk8GgS3ATUbjIHdIVFLSHojya+SQMGGh8KwVpfcqU33HXbBCW4eAiiHOXD
hK79lo3idEbVw9HmKGSvvFUpndYOdmo59ng5YjQN/V5AUYMRbbPr6sXq0hYASCQV
23owyA4nauEDk5pc0izR9/jhAmrHrCAaRlGwzlRiYOsx0S29PbkMvDxUEi/e8ddm
9C1rjcnE3Z3iKh+FS1C10aFTy7hROioBSGln65fwkBCo/D/hJyV7Dy8Ye3PASFDf
SOxUSq7e/4rvIXcLJLWcDLsKS4rk/pvBmVqLbaVklBh5jNCGNsbqmPMH8XGOXL80
PRRhtoGeZ7OF2mmwHmCHJjR5+EJuSkASqELOV7GeiNHNSOKlyHXIH9J0l7+125Qa
JTiBR2SrgSIX+CRFIiP9IT1u4kyFJfUv6Zf8A5kvxCB4nO3KCwUCqGIICNenaUoG
fqa/L5Hx9BABB+rn9CMEIt3LbJcjnjTe1hCMnmc2nLDbgZof/aT1dX6iC3t4W+ad
JP8zetAhfn+266HfiBvBUmStyoesDsaEBL44KU1lDMSQ5TXpB0bYjlvRFQGGGHHe
ZmOE9KY0uy8AF0+xK6R7JUnrRBOSFlE6G8o41h4YX6W2azlAT0OCoQ/ZvNKHKfc4
e2UU0ddeiqyJ2+RYd6Wj4YvYhZVvfsifFHmwQ3pdND2AA/6W5YsHAZv+UN4RRtl9
yVVIQcwhwO6yo2cdaFIIZkgLpczCufpU+vB979Ze6TtufdJ4pJ/yMx6JxE6XgqYZ
t7iwab41VaWQOjLgMLPYgC59iegCdoCCI6HvGfn0ztWenoejVl/QIRyBF8Lbda8j
tLXF2Ndk/tlA4FqNxCS0uoasJf2TxVqCuHvNseq8OKIeHcsSAEU1P9XyvPQv7AqZ
WRVlaizmvnFpog2tdhF7UslpNt5mL/fEYPNM4Z+u5VsuTL5t5JIljd7EjDqj0NFC
1Z20PmPfUQXaROxOlU7Uj9dBVPdVMOBPUXBZIAwjF7cYOj4+C+x7RYy6DpKvRcFv
5vNzL+ev3yCPVlkt1VHpdjy8IcIePGPDIm8EsMRQSNGuMflrGjPD/indn3+Wtm4c
ak54H2kEfaPbohBOojN+tWCuP3vW7WdqpjJNvHHW4iFpdXMOJso3B3RFI8pf0KZ+
2LbdKZwZIhPinJveGD8cFld8h2ex7pGGILW2T0AL3aIFnDyA5Zr+n4GvYIhhkMyA
sO9KvkBTpTZym5xyMmRiJ6Q15mPN+JQd3vaEnlsoXUvae3UuvKbkCIe0DhULPrVV
j6+/CSyodvzQva1uJ/EHxhMwfQAE8WjT+x+cpxZIZsnEshpXLLJmqnnrNMRqMFjr
174DcRqZIa7kr8ITiByoUsVjH1hOyeTRXphbx6Ssn4mPETpDvy/B3nsFcu0V3X4M
0Q9lpmWxzTBWEYR4rUg2q6C7VdVhaOrkq+kGcxSPIuqEKMCGgoSFuT+I28ceCpdv
F0+ZTkI3KB0JVvRsLy9qpuDU16reIrZ4YlpCmbQGAIAN8+gX52GQkD092SyfPx3R
CRAQqhtUoD3880Sjlp5DWf8akmIxUE8sj+fZUmBaYDgi3T4OD+cLv/tm1tV2DQhl
Dp4vbp6zXfnuOCvdAS1igHeWSggklAAibxC0/PgDHoBg/B+lWADXQSRCokisPX8Z
GtR2l15fJfnIIK8kee2aOEKPNL9HOkgPSxF3W8ELw9SZjlAqT/R9B+8FFFtP6IVB
4DmlNqGhbc0R/+yncfdzdEsGHjn28qSywNiWHlGPCdYlZFWNVvXPT5kFP/OTadKe
dXyCBOUr/+TfWgqmSJtXsFfF8AiO0hT2iLqt/wv8aYerBY2fN07p/eO83/P9fMu0
QjSO1uluXQnP7WaKdEdaYON1NdBc8Sy4vlVcEHEssmUOC6Wx8KRI2XSIRe+/zeIa
CcPedrl4dJHjS2QIperQ5RQVO/3+hWCKYLdNbusJYcAFCy6jkHolpZSsg5ZxxsE8
n5YAC7ZmFyUkFkZ4IIfFF8S4srBSN1y6iKAsFS6ak5yOpjbXPkcJ4gdmSMWACWPU
vvw48+a9ejXsHbdA1/dlPb2qS5qCXy/1AWrraqqsP6yWMAJtIg/xImsxvUg+3fX/
4sMwaj37gyGFlwZpN+ISY6eWrNA0lcurD17La1TrowTR9/p9LJvGdqvPM/TpqE8R
W/zrsInqAOfY7o95xSqOfYC7vXal0qavgBWGuXdgnxqewKlVUNOH4dK8GbRv4qpH
JGX4AsWbnwFKi0hOJoLbSMwT7Z8trh82LVNBG/cS2dZ4MKQ25rDdlePg/jH+4sf/
F+XFr5Ortxk+3H24pTdihNWU42wjLdo9QZ0uj8uZJKgKgnYs6+7VSdmYV66GGSob
xFnZTdSG+K99103Avt0GXAFXjQkoLN6p8TFEGvjYM2cc/zyRSczbUEX3x9REeRzh
RSUVeQ7jrBuzXhdrFHs3e+E+qbjUKWerk8HRwEuJVEaLUMuwlobs9g3ZYrzXVLwm
2JfPrWubinilSxAa8l/cAcYROl4712qX4YhuqMUjkjb3coRlsDVqHB6ypj+UAcz0
jok5XbKCPe/0+d8IOyUh7ka3dPBOgP1DE+DDZzpm6/3A2BWOqd9xqYMu8w320ofz
xC8Mj0U50/+tlIUykKJ2feZRRAO67qaR1/p50kj4SFlloWldbCe3b/Jc0hClXHBX
VZY6UIB/DuTN4j3PQx09wySnZF0wOsjPt2E7BCb6oExUQBZ0s3SO/XrfQ5zSBbZS
Wr+ryAhZT1eV56rqYz4Y3b7v2aioNVw31jGO3NJKtjN3ZKxcxb9GWdktL0zSJR0M
1f+25nSaG8rlSaBy6YTVkdY83x/R8ht5cGEGbJ2YgvWp9DK+AjbH9mToQ9GTTIhh
q51ThW/ul8AZyiNw3CtLRK3zlIYiStZ0oY8Sd78GUU6AtVUqMdgVfj0iCmNFrdjs
TdjdvCOFPBWXAMG84WdKjXrkyZLSNE0bxSU9C5juoHf9tIRNtGc7lYTX79/4TkiG
UiRjRz7Z23nu5hGO9Oh5+kyegH+JKz7krV3ThPBWnBJPjUO1szzTZi46tJKLYEpm
hN+I1c2rzsJ3lWKoIE6hGyS2agTsImDdgvccCys1ktO4SeMXLkyLjXsGN8xYobN+
wGZuSNHLNR3j5zmhyp/E97jZlQhI9o7o1N02b+D8gXMUDIBCFsx4XQDXcKFnwqg0
LT2D+h7Bp5O+EQalaG8tdg3J+mFst/pD8R9TWFiFWFthPj2DSZ4o5+n1QXtEhzep
NhF6EdUNOwh6cFYyy4B+Dvgn7VpJIz97QLuRrgvR0Z1NDZqdSQmePwE27mXp4kL3
5JgBQaB0jtqj3ft3VqagJkfADKHZR/AnZeYl4lUV7Th2xyayv8eg63BxvgZx7p2c
w+wH7UbjYz+ver7qAej6PBrXExY8paT9lpTlgZuXYvbdCP27Phm/O1GU1Y2FoP8D
puiL21GYbGsXvPhO1NErdIu2NkaLuAcSZ8201TMRHSbTq1wghMGQOM6u6b6sOrUt
9iAFsLPuAxJsAKSEOOI/bbZMUKKJtVLGQAkWMmLt3NY1Ms0IL+DoBUhNChGZQ8Yh
DmF9COS3tR5rGyk2YUW6RFGS84+sMOuuHArxX/gyXBP5IyBlqiQXGXI/UlunQWdX
OZep+sJJk3AYYcyn8zVX3sVMs30gtKNkQmkr4QnqqNNUAmlEVXF21e3sOa2Aldxg
UjgZ+fEPINA3wjMYH5pJbnTFgdwVmhpuYVUu8xdNx90Er5FaiL02woPbKxOaw432
TAThS8oeOi/0XvajmUFCuWH3dVoewfZyZwyujvokn4wvVdZpYiFEv7o81BqtdHQm
W/INxm12T+ZtDF51WX/n4uvKuOhs1Ek5fnkHQDClebh/XLon3wmePox0onjc6aKP
05r7zAryinbYb3vgmANWg3VNa19mnBubkxpRWMDzmzG9rxe0oo6Xy4PMAGxcztmG
CFY9JDSnuUe3yo0xKWKPoEGglE/SdzvTRJYTRONZcSR1Ou2u0Cs5g8kQP58jZ0vG
2M7stB75cEDRUDqmqP8vqG5U3hoLLF6gBRF23vYWnzXciC6EJZIB32fptFk1BLWF
aph0Ew3bAfjE+6PlYO3ZZ4OFVtWJvH7MMPYVXamtRpnr8B55zIYZgzhPPSwgcsIe
leT7PHmlJc2QttK5Uubp13ugwt/DPEC4acyxiUmuTESchCPjpRyvcL8gEMfnAxql
f4oMFqW2FYU25480w/AVdpsXsM60m5hcj+0NAOZAFRVBOjKoR8zK3tqxJ/XVZyOM
wqztSJP+qSV5dT3LCJE1IAzHbPQkrr7lkPr86T2XaTd80wt5ngwMRqebzgQLO8T3
wLcVjjH9W16Dkrzb/ecUXeo9faHIJwhC8bVU7dc8Nzi3KPPQAEdgr9Unq8xprOT7
KtVvF0Vm+2/QYbs62DLY+Item8eHWm7HRrCwEQN0fopoDBRB7PZzI2gXDOz611k+
/geYZO8DidhNVCrLwcPX1OlbR1qsfKCvfNwSFOB8jPekBu2flMPRJXXtvd3q9zOL
+nJ6Qk+NYk4F78taib//fsJsG0NcIeN3rjr4/HRtau0=
>>>>>>> 426889eb8ce467b9c9a9f74dd4af433c5046285c:deps/flexrio_deps/PkgChinchConfig.vhd
`protect end_protected