`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 57664 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
SWiiI4+6pDvQxlUp4hYEIgje4IyGnVPDkgibV7UsI1W5moIY6gyfZu0XU3FPWp/X
keFVAi5Kgoud+iOCfdLIzrP5+kZXpxUsO0WkW4n1vmL7Uo2cq+ImgxJowTaId3Oi
DulXX5vEZwubrqcDTtApy65C7PRnnTFOxha3MqKQZmIZh8BKMiXbv79jc69fxuLc
xQRk2H3swSwpYzvjfwWEy7KLN/O9BgRTS0TnoWyfoEc1RkRiXuAQ9zlq90hEwviL
7bn7kz1ptHau78ifeGVXnGMQ4QqXGdYK9yIKix6lA6Cr50Ok8g99SZch7c+PHf3E
4nvqKrB8d4yvKdx2ftUTn23tD2p7/In3Y6Xgwi2gMmUZNYqMfEwSTwgvBY3QIebx
0hmc8yHWyUCbnPJGLfcTYfKpYr8qS/aQYLSgUcch0O+sg4/zkmDlVsVtB8bnXAkk
2l6Ksw9UlXlIMEkNM8pQaxGrr3AxJZ9NdZHuQU6eH7vI2rKM4Ip9PIDK+3ueXTzs
8zwcg9Fafpdih3C+LjO+OcRGijJ4S5q0nedy0B4clSuyU29roPMb2mpkLw3p6pjZ
7HePa1hsEfviHlI8Pia9G9YSsQP+mNdqH8t33qb8NUeJnwV0G7iYcaYPqzq8Fnn6
9if03Lt7ejZ8fo/egeHZQeuc0FmZwKR4uW776Al4LYvLZEOK/wFUEHrRseD5WlLI
DCG/42MSFoWcbSCK9nghwnqvnoOcmmPmueWf3MKx8HHVeUBxAJwDnvIQOpD4kqtF
/8+3oXDrNQ2WzWn1Jm/RFvqzTM82LYuCy8oWZdpZ5d5Qr2m+QYvqjEpfPqGZmXD9
FBSctLRsdsA51vfwkJKcMoHjl/j2bwRnOCx1iiVbbikIwTceprrrxFH7pJkZTxGM
vHI+TI/6nU6uOEIb4Ws1vSkQ1SolrVQ40Fbgrmznf+x/Lqm1yQh4c3htLUe4nYIT
6YsHqaCgcjE5MSEQVNtwZvbhHwR6t9cInsFV7kdyQyCURlt+ySCfAZP8jejNnwkt
/wqBPWzakltp/aNMMS0epxnI1yf2wE+h1cv76b7y+ZB+I/e6vX3NIXiOjHmBpsyw
cPxh1SIlKNqs8zP1+RqHUiiViKceJKFtDA20J7ktW0HxyBoha4bzct2EmSyvM1TW
o6hBHU3vZ7YMWmu+GHJibbFvwLM8AqEH/+X+hJiyseeWKq1Alanevg047Z4sTvj6
YpfAmUB/GzUiwFfp3jCh2IwhHZeKXgKkU22W7lxcRSZa15qY20g1bcxEVb1ggXZj
ALnrquof4wYqEMjTMCul7kLfEddUcTNEq3ZsVok/4ebRy3XnjzhLHVVMlUe605K/
Q711IRy/SJkoyXzYWneR4aP16YOr0cmfCISH+movpFf2fz1/SaUI1OiQnT0AWPoA
BG0WQa6j7a9qhY4cfYUiA3OWWI+3+RPafPymTByP6J/cwooTLO8RtsIHStTo7SZy
7zNoWVTLQDlPKc3JzTfW9JYBMgZ0saX4vOPYHgosl/IZUhnKRXYb1jMddKb3Vyqt
/mnRklesgSBvi4ruMmxbnsQIeGzMZ2G5NfVYCAz+MSWdKZELBPPsQSrV9vA4KpcW
Y1ecfphfWJPugPB2L2MmRtHWI+pf7NtLU7yeq3mSdnSQadOtUrF4HQy2Ye7rlhQ+
WYOheLzEFhdYYfYb1z8L2XCBOVeJC8q4CKyAz3OozO8kff8xfZyVf0mGoUZjK5RP
CU+eirCtqr8PNu+LjpYPk55t3Ugmfa6RIuJ5i8Glc6jMjB/G2IZRJkgmRFR6FGCV
JDWs1r0uIacdVPsqNxPmzWJ5JAy0tmRHm982oDv1I2m+X9dcAuxIqReUHl4j812w
bTfZ0FHcQj+trFVqWSpwzr0Z2CHkWFf51d6EydlwZA9hOoAa/rgt8CDhkyL83odj
2s4H5gZA78icTiYVqEFhqYrn7xAQ7BkgRCFhrqxf3D7+pNWwBpk7PU284UTZSWe4
Qkfzyb5JiNVOd/KBVuVF2+/VQnEUvOyprEO3AFwNrEjVlKCVbenRR5Hljo7oi+V0
S1rwsSmoGnn0BX0ujYnxtFLfvlf5Gr3ySJ7NYkH3bk4gLuJBoIQkd8+h4r209hpT
bdmMZ/hEAMkVNGNHHD5i94TJDkHQiMePw8sONZ+lragBRK7/jc/rHkHiga7BwbAi
3ibTWVq569lAPO9SKfVYhnV4SsSkzbIwUcd2dEyUBeM846rPz8qgLQ6hTxkRD1TB
+RjhePpHYR614TL73XBi55RmO72m8bMVALAyXZyKwttJ6DYO+oZUvIjO2lisM6C/
JLGhaBlQ9tvQSiFsSVjXNK5PRTQtReL3vSxRT2l5NXOFsxSi/SQ7C7/jN3ntJDWD
cChCiAke+r+XM0p2dt3iM5pIasX3hFumrsFKph6wd/chUflxtytAqLnYsE3rdKfB
popkq9asTvwaZ0i0V0MU91O83YbxAOJAY9OD8PDcjkHO2FYLNQfQgzyJHRN2urlY
A6Yy5RZyRbbiPP0Kn0ExAKjDy3wBLdre5NMJnVWU1UAexJVp+xiscT9GY5DUQBBH
0fb5hXvltXQobrwf8TfaDgQIQQdxHaYuAizjPXuLcoPDFO1KttBatN7JrwrkknWz
nwy1EgaLEpUHVVeqMN9rhRiKJHI8KSV5e5PZDDQWlJXN9VkneE4YPXwwCViLfCfU
O+7I2SS0ATE1lIXMzrub2te7QCxCC8xQfHTnJLrDELwxmzYQ50WhCD0AP+8owOzW
diateNOmCFNtfWtyhxF2lPO6WNnk6CMXuInh8aQ1DGRX8Nu3ZONlFK2yqbMSCByY
1iAJyUyjuu2RamlVpDHMUJeCC8zUTu4ssQ/8+pYQ8CCSPVOXHBNFBVGWXAKEEjBx
BmVM4Se3XhnJJUkJGVOuEeO/HBEnzlhi8eWDJKO/Hb+DxSmnEFr2EkSpfdqz8RwE
8WR9yUwWzSZIRrnCtCmJyqFNXir58XnQ+16CJ9A7pRpI7mP+zJjfIj/y9oirrfPs
GP5e+OcmjCY1csD6SLh8WZWD6gZcrsGKi6Rh68jcR8aAVPd2otpIQqyTGSP8z/Ji
M0HfKmdDouNLkN7HSNjj3Qaw8uTgD9w8TvGZWaYGbn5O6dfj4RN+V+S+rUNvYa++
rN9vSNUASRw2q0w5wDu21hICJ+wGMwg7pR7mLgF0FLHOuNoDNwaKzU3vYUnKP2jJ
Y3IK7BPt/ia1HxQptT9i3UJ3wGGUUES5Wt8d3CkRFeaNrAOymCOwK0crSVD63dKU
gDip9qn8Q3jdWYanufKys4xH+jx+b38677taN4N68rxhCcMNDMs4Ova1eSGNtyIx
YfkQ1g5HySXrJ0XtvY7E+ps9g6h0p4s44jPyuYlklpgPpYjpaXvQGK9s0GCSwJzF
HasPcgfsgPo9mj7vB58gEm86X5dkCJgC43J1yfzR0ZWt1oYGVuLqx+oEDYWVsdYc
W9b5qGNoOanIrEGiJX6ZB14RuG0DVrQ00KAd8jwG+q6zUj1a4tgjhoneq2fz68d5
I7ixK1t4Hh9SldHR3hHjEDl0J5XwogtvOllUENpHGK3trr+aSPXwjlgrEhP+GWM4
XLQJWT4qBEhzt3/02USUVqDTQeFuMlDlvJqdQhb7nHzJYAGdRnPwAM3allmVSAMd
25MbqZIiim+Jguyto9hwxLs5ZoOk81kXqWcxvzsjTp1f89Kn0W2dXFdQxZs5tlEq
E7YZCF7cc+YNonONdhVx4XVnlWgQ6GFpEK8PctMeFz/nwep/ikCPMzL4kZGWzRF/
MQF4o5vm8EhDzJ/g2MgAFss+KQNpIrCCnDSA/9qHx3zyi8Y67q9WaJ7oVyHlp4qS
CgA1P7kJ3+/FJ4Erf7FFpAOqx5f2fpLZasozeu3PeSXOgGuI1ooyZE3tpjihlCTQ
LoNZ+/LB+8X4A8SNZ71sqT4nNo6atAJ+IOmicYZe3ksoW+s1F6gyZfHi8GkDmupp
yfLToWT++IEgqkRVmbGwu53HH9E31U34Gk2yJxC5WoN9FdTMGM1KVsSE4DbHnnyj
IkHAWWLJ0+gUEGOwX+C+Vpy8Iuh3aMjXEx4OV5ZmzBuesJqTrgyhTDchb0P2nKJE
XHsCQ8mM5ZY/URlgVr8nmsmqM6pnSJ4P83fQ60k1pksKz1XMCaGpn5UTzhBkY1UF
6EStGNHRf0gmmj6u+htnI5SpxI/bpT8Zl+WYNBKa4vd1dZLr2R3XfxYTxY3v1PEB
2GgNW3csSTXY4cyjBUi0Saorub8/BxHooOkGwsJPDTKbCnlXhYHKKbnkqa1QafUL
7hXB+/R9Jgg43jWYARanHiei24oXOGHm0iUgsZ9ACVnXcj5BzquXH19Rpt5ZOcmH
B/OQUnHD6NAnd5XTN9Bsir32Cpnyk0XwWC/QuRZ89wHkKBciLqiQ35diHW0JlRUn
Joepg9YX8fOUO5fPgYeG5a+DYSp482VTaUJQq8CE6ASGeZLTUoHh5ajG5OUCCHBI
MmVn9XxbAEoa1T4bTfWxwsT3HSA9W2iWV6t10ArVWFoUp0wUfj6SyytGR9z+ogXw
3TrYF47krbAkxDGw4PZ23HWlwXE7imhwzKBTr8t+pJ73JRLb3jFFbaqVcN/kh5yJ
ZsCkpRhfWzNNVF1kmtqMg8hP4qmm5zNaJ40LrfUYu8fGLEB5dTvoJR76Y4w+j0ac
MXlPVdHN76/3qQO797bLgtfdpzT7RgTjJThbdZvKDDfAVZ0o0ThzM4Cgfr+ch7Ys
UkTC3YF9EEYd7yeIdw7bPb2Z0UCKHutgO6WS6ZkaJ1kx2k7wKEsqHM5j7T/9SGZD
2FuowcvndnzKKRYzvD+ZntPCSY7RXnhEO6Dx6DQvX/elKJEh7NKVdd1Y+NH7cUe2
mdGGNpB/JNs8AnVrjWX8FoGq9CLlscOnQriMFpNR8uGQ8u4t2hANCsUfEjOrP9gn
FHoxHR82F/DX2jjSpg+Rr/9HzMOgK73bmEGiVsEsYD3orryqNeRGCF1HfN0hKF+A
qO+m7cLRqQMZOrU/RTsb3czp9O+LDr2vDeShCA6oeAsFTVphsxwAzpkEIi0KWKeM
B1eORYmoFcArqv8o+FmJCzmYdRP+w/50wQQrqesT+dPwaAHBwNTXivCATiSIn9Xr
G1M139F2MLo6vZ1f2iKkE6QipIFUnPK8mXc74vs6KNGUsnkreVtCuxfe01TWekMy
DL17OzHSysHbnXqYs4sz4wq+YwCt3anqIOeNcLXY1QQNESXU1go+VL1O6ttjMO9F
dKUCbh5GKkVRaFgEVYPsWR6glsUWHGhXPoTESzvxeLz7zFgLaXk7C20RNrjHklYD
xPKr4tDcZH5Uc9EUAlBSiEJJxmfe7m+8Drk6pyLJQJ6q1wItkKwqxM2y0wr988dr
vqaBc+EjTdF8PyjSxnNQwUC1NMumr/1ccsrLVd4diKpjGk/lho7LneL2fRn1/Uaq
E/yueeovrq0myRDZPYOLvk5bLc3ib2xxKcV9L3nIBT92UKXkBnqioredp0FUkuLi
MNhPO4mFOnzpqryNxyQRW6YjcHQKYVhNab+jZhvftxCEx1ZCDwOd7SMqbEaKr73C
VqbJuV8OE/YKeZYmoXnP/dSRcmj/Ddv87R2sM6gImRMZzkyAUjw4PsSC3kxYleZX
8S47MP/rJX86MpII42JkPob8klV+U+4KyWOD7xk6BV7d+WDeYeJT3OGyXVlObKQA
9vWNpuNcHAHYONHMZwgzZy4SPpzNSjEsfzz6jeMZQoif68FCGcF4FduhOhqw1lZ5
ya2uf7fJg5bCSypPbSPnqJR1gt+zO4W/Vd5aNxLfc/uLOoMpPNz7ycs1IGpRarEP
gvrraGaEkta0DD6pyyGhMHmNrx4SatK2HwkqoKEB02E5hD9xBNdq1Ida+BIXAZbp
nhcAhFeGaKtr4WWmvKStKNEQTCRS58IEqbkP7M+YYvBOyFGQks9dnzO3hXJEcf90
ngU0V4mYZ+blI7C1KVfz1Of6xoqiRyj7kcGmom5JicCx6SOFUa1EbVTBCyo6G0EW
UgkY91HEUhhj/5FimADA4flvRnHRet5C51UeAvn8m8ZcUSvC8UFwDrFuQXfYtFHg
HlvaMwoHvUFHXbxRjscp+C228fxCc+BJ4P/sOqD/gVqOTBFwnNF8g9zqzq5erj+j
BD+O6XwNaqMRPg7VURcUZYlJqRdIVLeV/m06sBG5SpNha6i32U7l4nkpAg7d72Tw
nbHuw+dfwuyY+DnFoqUMD3XOmi5ln0aOgjSxxfOP9CVjhVebopQHHHC1sUZRvMEE
rURdRF7VbzzF98FmqpVv88/qj+wPNaelJuCyjob5/eNwCJbTp8E7Hg/UEhUW64lv
qV3wkc7HxuzqG8IHzcuwfIjPofwCzcDQPWFQKvYj/7OSvzfWo49y/ksfZrEaqJl9
sy92FfxgCSl8/1GHlPrWiLWosV7/LAFROSByeF66e3Uidmk1rsq1Q6XLQXsTsQVD
BiRlhGAPmsxYpadkzndmj47KQIWXy8700KXYHB+VHHaeO/hoyfxRQELCfVtJI43v
r/SzIpWj0rjWTKSVsbbMvX8Wp+Su4C0trVkwcBeN2EvfUzGg5t9q3d7ku1MflN3/
2xlF0GFwNbiYwA3PMQNF3BSuHHAuWSdjprlfB2UV2mNBY5QC5SJBdL2bkEiqXk10
pBjWPtKdwraN3uHMgqQCyILlxnyQHXr3FEmy4dhdIUJL63TtB9HY8T5iD22ajGeS
9uR+YzeqAb+feDQcs1IjBz5dpTBeZu0og87yn5jjrclcUP97i2fGJneQZadSzvT8
cQgfzyUwAwPAHLE5O8O9o3Q3fMvKGtHqVMWxvifGv80ItvDCPo1DMoNMbV5byCr5
A0P+ZzI1hifGWUSjOZiQwKIrO3bSm5QeZbmUNRT4uiWkM1EJqdq8ICFCd9OHmZNQ
0vIZ6AlAN0gh5stj0wQQ8AC22PfdVONPMMrncsu470CGmpCmcw5bs4FlvzhfQzlk
QxmS/JJl9h5/UvATr1LjbNylQpYF0L0hIbK7DxMoYu+fWvnA9fnviW2ObdMTlJRK
ODIFNpkUw+RLDlSW8WugmKlhNKS0P9a/aO6VnFaFSOTboincYdg7sd3zemn+ActN
Veb4y2L8NuSUAszmKXBoH/MNe8oSuIRlsqbPswTJN5mbP+jr97ud+fuHBah2Kvqf
dxx3BflgkanCMJ4uUTp0kDn9cQZkuKyE59gpRNU2GqtUy2IYkBk4InZi7zoypEyD
dlyQV/xNfeNw0ck71ZCZV9dKNLtJNZXViP+mo7gZU4BmT63eRp8eG+ADH7qMvMNd
lsUVqbM84Si9tL5nd8DgCrKGuJQyZajtveYTZRpcLT9r94BWuFtxx9UmW9qT3qvm
R5N/V37qC8L0Hat4NQ4NriRuTJoKWfZMVD690jH1L0+kzeRZPIEuXqCiL/xDQXOL
/dTwOOjlgxnW7SIGEVxEABR9xgOecUhLxUnu/htgQ/CrqWaM/9Jin9xsCRxyVw8B
SeGfDw/2ylRmPG+931FWZuxDOVtPa8qykOpWx50Zu94UilZOFWRrE6v5eQ+XNLHz
+qaFeHoEvDRvV6uEwtMXajJJeawi8EdXnrpphCGf6+yUaU1UdBGe7H723YfKJWzX
LEtBaxcYoZFw09QQj+6oj81TZNXubaNzywYnO4EMjKh62f7hp9hAiZ6Q2vhdSyxR
NO+MsQignvHHBo+u0aKbuRjo7Y+6Kea01LFZyzbYIuxL6eSQxuQNZc2jBrOufqEW
Eyb3rZpeNbti587cgjNe+9Y6fElqTof6naGn+blKXcHyDwwJzoDCexZ9FRBahMfV
3CWFJfFp1aRud0FtzqhyYvaph5mqKzbPibyFQTxeBvqL9qJUinHPnyWLXfdwMqSS
vrv0kBOnkse9M9/cVlEI5lK9WdSJgT2iFY7WyluLLsFfNdDnxjX8PH6YAfFvDXGx
8UoT+9+iRfRCiQSiwm5XqZ4TELs9+RBK07A55Oghe6FJShAXX9mLtLgLdw/mK0+i
GlGDxFBqpUgbWaF7BGe919HaAm4EMNNWhjGFwuJ9V9feO+jf79iOXfVMioOtxNIL
3Astvkbtn7f4Lxp2LFP7wepHZbeS7Im2Rn6fw6PIHapDrWQYc/xCfzoV31JYA33L
IotLkGCkHc0pD0uTm2z70rRMtDNV0lmFvu8iaiFAya/ahRBDoexl5D4dYXJ1Lupj
LUop9ohGGFyCaqgnT2x00Dmrbm2ox6fs72B7LUW3W8a/nRw6yUp6T+lvGJIyhcMf
EIo6c8MdfNTxsT2y/5U67eQ2zSvGKtt5ysJvjWCAWyq2KS3k5kYN88Sf2ih3klaJ
jMhAWyWEbaNkMqN9cjlAxvCKBPhQiOi4V4Dxf2aX28e9D0Rm7tB5Bk79dsIaOhSx
b3jzMpkhm4cPWGPiWyFap7G+noAhNP+ys4tSKh1FCWombkQH+xCq+94zUMC5ageG
6u/HAflPELfp3nBA/bpRo9+J6oVZonex2PjMCBOtpKRbCjZeEjSTfy+hoiFgPFpA
DEmKU6NhKmm3wgpRJe/W8hTlGSwv4heYiVXsg9ZQvlUaiitXmleSMYmKJ7prYD/J
B1qd2/iFwKB7kNY6eyrVKJehMf8pXpnjM6V+bsJDsMega231l+/FpXZtpaDDiubL
DZ4XRqlAke6ouaiFcwWvYOtnJ7DoMv/lR7S+Db7TStG8tC4cPMKmcQ5QQKzNFEZI
9NQc1myLkxxq/q/So+MiD1lg90wY2g0I7KDiXYTqYMMnBwYEo8pNls8toeHOex1/
GC16nbqa9wXoiJriS20ufdsoCv3u+SP4naS2TdFlMhlp/ukBctQh/jnJGUbMbvKJ
58i/P5mnnip4Q4cdLZ5uXHWHXNP4y+4mhGh14o7yX6oQwI4juCpBJDiSUweDZJ8s
CJZYQopidQMHmEZiCQ72n+94cJAKZiCdH+UntEtV8IkGh2X9ujeIIGyrFQHvhEQm
EtSzBRtVKnJus2bFCTc8mAER8MB8wGTXMh9ohwDQk9bi23dM0fR1LyW1nLsIWl4c
FCAybd79KHW42BxkT96EpP26eSL+zhiPO9kzYetjul5BGqOU6PspW0cvxF4293qu
8fzMKwo0pCA6dvF2UwmuklvgjOtpl8GSPBvwg8arugdIokThE2BByuoQWjz+k0/y
oMQBQ0S65lbrPfc8/oCbUmXVu+B4ZM2hp0lFLpUFHGohWhv7PmazLXwOhqnGTGxv
nu9jZSiOQPKpYH66rhl1fDxRkJPB4uepDz1iO+JsJ8NDGqD/XmirQsubToFj/uuS
AidE4u+RTDjQrZD4fEol0qgH6XXmNVyrWDrZxeb26tbW5yACBd5bdzOWKODwjpNP
Rw2tALHttkf54vT/o/KUeaJFDEMs/X3+LdWHkptTuGD5ULJ2bsDPw1xWaoHeFyUT
5u/cz0aIG44szxKjISlS4rtktAZ1X2E9jor8EebkVvoWsv6CU0Ogpyr4YwSFU4tg
ZVLOhTabtiqEY446rm2mQM2mm5baLYETliEeHLXVd1jeY403u+hwQd+nVEJtTIdn
rmDRJkrV770D8BLuhL42eMVN7EOHVIMKjdT17q6/cQMAy86TWjC8NjbM1HppiiuL
cZNbEKuA1JEgEs0+34jFhnEmZ/YFgb0yynvxlDRG1JVZ/JrFhsJtbsa485qvg9HO
TJ7mMqObhB96rIutrCNrbY0VI/kkbT8J2LzlAR0wfOp7d9eceXykgYExNiaJSDZY
lCRYivdAMjmwN42fbbGFPclDlZMVV23Kk0th/W+N7xQoI8Al9Z9lPeh9SjAdEMzm
mujNMACtyxRMfk3HY3AWU1YseqA+cN6OZ5MpEYoBE12tqcytZeGG0BrX0krFxQu6
Gq+BmjW39JYD0iGCa8BnscLPhFqpkchJsyjiqqhimBdkQS5E0bY4Z4k32L4M7SsU
xvILk9WhmVyBZC4hStaSCBbjdn1uJYSndtUEbm/rZltLY04WdmXqRKBOdjMk9ARb
K58pnJD29yLvRbZoe3Ps29+tO2lS+XUDddXpGV7IdauBdYj49oXM0uj+JDtVORUm
RMgdj/wB0Ppg3YGRKm/jbLOgzWzYYUkSwS1HzMacjfsdcCeWWauA6h33n7gh+Pdp
tm6Cq6UtOkrPiVYnJi3PJGTgzOqy4hlWqwj/D7xK0qNvP/4Io7fyAUezWXYqPC9a
hRZdBw7zCEUyFbL+dM57s7RLT9DsuNiOXvdNpS7O26wCqEZDxCsOu2DTWi4OoXle
wHuXVMITVwIB7vr7WB4HLERhkzEIWUlkvdiBOAGSY2m4dBlFQXj/0d/A6zHbdDcH
sOp9z2gslP45HvOM8w7PpOeJFfbVG3weSdx22qmRYTjwCPoLt3e4FenKFFnYEx0I
aa/gAlFfgJvKEO5vk4WXw3Dr7RLElLQKtjZfkVeD3Dcw+xq+LmAJjhNENj1pCu98
pdo5PfpnDJqNXMHIYRonywvqloOrvE/nx/ZcOfvJrhMiKgrshzwXZkmIJ/7L9M77
kL9GI+maZJKG9grJTYz6No1qYbzNTxMB9tMGiRLgMdioNkD4FCc3IwY6ZRgiOj80
QE8s3zM0raGWBsLO5E+TsS52GdznBoYmlisPIfFSs6hFzHyHmxmLvbGEPecP1rXd
wmVwv8bv9XSyu6EHk5h4hNVSdHhCfgC+6tkQ8WaoS7r/8Lp0ywF552R7JL0Bkvt+
wA+pxbo8qNzUh72iN+6TPLhO8gtORRT2KFdM1n8TmR16fjtF2osOoL6/hgG3dONq
RBd5z7dJqnUWA5Mgw1fkryZUCe1r/Q6rmLCgi3KBEmTAp9nlFizpgVbTUoGjMcQn
FFwUsAh64qK8LGF+W3itoAYkcp/C/z/tgrK7ss0pS7R6CpanUXDYDjGHTPeZkkps
CMdWkvKh4Z6uOBByxkbpPiuDN4EVHH5qoGSwYIy9zJnfhMeD6P5HE/d3b1bo6v8b
9Jymw9/roAJzs2oiCZ5KcLvk7iH3l18esGPnBrgbgtbY4IVRUDOcuMBe47Ajf6VG
0t9qvH3BI+eoEOtVJ/llj9wLXYBxp1KnwRHJ3zF2P1dbQTbTiHCAQ4X5R4MT+PdW
214lWs3ptQlh4viY5AvjJwHlN0HaK1KwFJ21qa1rJqnpKDNPTo2WSHtdUoK2n8lX
vQOh9VfeY0ywQmR9OieAUf7ye119B6uaiwjygygw9Mf8MGfO+ceF5bgTZRF2uNjs
fvRtn9YkBuCtH+pv/KWVdd4g79XQPOlndrOMTWaeptOmkW3bI/dzIodTDc4l37lo
3twAuR7zHt2WRHLWpv8YdYJ+zJsZ9gJ8xIF67Qnccl/L3qCU4Te+dA64ODo/wpDn
sezOKnTaLQmJgOGS1EIhCQNlxm96BK286UmLbN1WWI/+ogdJY40He6wN41/e45+P
InWBGvLRVGmknpqeM4/gIl89hoLcDKfFVtvzm6qeZBJBhd622/bnBR1PoempfmlY
2vuVKnOHmVMzkaFNlFQH+P4QSzB9Z9FtzKXheV7k5/fSPrHzctGxu2xB0on+OELH
6RyCaCIKXMgE7YgSplex9bQcB9k2GPCYVmzLOWTqfC8gAx5giorb+RGisDULsZ1q
w7L3isKhTE9WsWM0kCrHaC2ag99k/8BIFGi74aCBbpI3M46XmgLj2PJkTGlReX7n
+/KnpKQAgTkuImgDaUv/A190QQyZBMVNLCesLHRFaeV5/z3921ErQsQe2CTT7UgW
UW9cYVpbY3RUpGHziGDeksIlUAC28crxIw5mbIVocjYPLhZT6qYrUjLYa9pxvqlQ
AXdGjfdQD+p3B1eVEERyRq1+OStPuxZY1YD/XNh1eYWOhxufqDDtZ1rivhbnaNme
PqEc/pDW5Ev/DcQ2rndB3EK+LPMiYdt7pUfj+STpZrTte8bUx/GibaUROfgGi1dR
s3GcIUKQ9u8rpVj/L7yAGY4E/FbQ5b5LOicYf29kKCAppQnmdvG9kz8DYceTPFh3
k2eCegf3w6J4xLVlrix0K/xf1MpHiXTGZB6Min/NYBlswf8vuatlnbtI/FwQSnP9
QPQmEt7uyXjoOOKDovWNUDXkPsLqKzUB93Mkob+XZmN68BKjPS+rGdMfYP/G4Ic0
K57M0oJaEsGSlp1wWDeOLSopR8g5HsbI41NqLS5LVG3tf7X1rI23LeNfjIPPWzC7
mDNSc6dICnE9k5fPSas0ZAOEDk6yPn6ySPG8IcBlaWAzpTp0LdAK4uSdwNWvubjU
ZRYhIt1cjkJeCsxvt4whq8iHTVfnUy58qZZ7T8JN8EjPuvGqhsoNJhY32ivJf+l8
P0z0Oaim5HGq+000GCzMemlmJzHiO1XAev+EK2rDcNjBuSksHOm0zIufx6n5V2XK
XkfGlk7YLsDdM0InlbuyH906IgR3cz+aaNj6gQGz2MlG3DHyePlmc2yLcE4d838v
BZ0Wz54XGD70RPTMpG4Pu8ced+eAE+uW74Y9VSCbSUUV6zeS95PEXF9VP1U7os9i
LZaZ8gi5OaPMXLG9D9XbiJvumHMsn/aSoG0a56nA9vQlawJ8w6wfHdymFWgtVry7
f66QPLcaKy/v8pzHIrNSXsuQI7EzVbxLyfsRe4VY17aioWOeFHQeajxi20nBfL8H
0LCmanMbbvpBes/iVgxzwbcIQ7GBcC2iQGrBX5+048wp5s+E/oMLbhmfwvs7y7eX
dM+mZiry1RMK3wXs3WokK8j1awrewre6eCCZPkngyL9iAz9d34g5HEjKCsYtbVtZ
kPMYowT5D/Wf0pKHkk/K+Y668UYUBw76iwt5DzveNFHu3sj9PDnFQC+SYJ6mQbnQ
oQwAtM7RxCeYvgjtgJKMop9ws1N+H25fCkWWwCmEwniRrePixpDSouKEpZgsaeXd
FLWUYRjX795P/ogXcvH7c8PkVhqn4R5xCOHrASGG6rfreU/aK9ftEtQXalOv6cGI
GFdVuuptR3GMWan5Qr+mhIMRLk0oww6hRXg7pIgRGqp6MZg9lfaywsFm22juGvBJ
AlFRg27ofwAB+OCPrPqD9597bQHZui6/YOx1qGHM2At7nVWtfdFnMSa0xjyC9C0m
J/BB1ikt8PcEVyn93S8Dk0Y9pHPnqI2g3Ob+Gm5lbG9VIkKakZI3NBCZwVY7st57
BoTyvC9rmvBgYSAKl1T17L1bMEHbI+ue/JzOnQGUq2oQxj1i/k99mCsnz7+YUgAW
kYlDBjZzQWxEVHXTYfuOrxxaque7Ck8/niBDt1QCLFr32jjhEGsP2z8GV+FZ5yoj
gMoqaXm+p4Hw7MBvZLBCmib2S2GBYRfuIZl+4iU25FFus03OHtvj5hM4k8MrG1Bm
quMuvahKfIZV4Adwfn+rG90N7CzakHZwByePQ5DF/NL1sIiFFMY+hZKUKLLuQpIs
DQp9XF0stkMeYvuzMB/eg1w75NIk2k3Ix2G+Ix9GpzEKfk0Q19Bq6xIZigMP1/Q+
4ZN88nKW7zPNEfF3nEjUe/jOyUpDV1nXSLHzx3BCkms8RbBSoxkrHN1SxZkOHRmG
62HBojrfXWBAn8UYcDpIUgS29WJPI5Wc6immUcNatvJj+rpsUKc3h/99xo4mK/CO
5VR3pv6cu6NfkjWfoIe+NjTFqEA1ktrId2QqmsQ3NatA0ASOidlDNEYMAgq81kkh
OBdoV1FE3C/xsyosKsjT4txn5fH4Ty5bBiBqOBYYS5Sr0jORJjCBe495SrBxLwZb
BtruAQ+zsitVA4LyKP7dQPgkdHkj3ZR0e1sXYjPwak+Km7FosLKBtzRJfGPkYikG
gMhBH7LUxoSqKZQw8HHhxxdfEG8fFQ2g+7BWl9DDx6WEEeXogwyEXd4lRBAH3k8Y
TTwZIf2jSdwmT7BQc38Vo0YS5lR+4l/4nU9cgSHw4ttAaMM63f2LAKIEK/9faTFq
jWMBN0dDZ5u4eMh3Igx22gAmUU1N7OBt9NyF1VY7YixJZCSsljn/9oWfl5rH9mja
NJ76FqdFfpN8TMdyKbzYIvVtaCHSmrEy+66KBLLWQNF+xMVXKsV9g3fTe//1hGYZ
5foNNPBweYqRPUmHS6vUCi1h9Jq8LRQ6Vj+dj5DQLtFmxjw5DSZ/ypPWytRc96GW
6MZMLLJ7RZJ6RXvHRv5J7oKFx0jQZUjNJCXDPZEa1UsYxWclOInsr3HFJ7+waYue
UOApzAcTKLO2dGOJNoKUcVgqkscndQNwqcFFj7jB1RDpsfODQryb00LGcnUcUOSp
ue1lR/QMJGORx5JiPDPSl7HlBiPMnexbkjfGBKDe/iWeSB8Oam6Gw4gyxqwbD+5U
egW75M/Dsuz8Sbz/6aYcARVfsKvjBcp2RiPk1RnnxLjtoz12MLTn8FJf7hn9O2+k
mIDKx/OI2RqkonMCd3Gy6VGIePD4F/bsPmvapJi8VwO1hvCmGnTDXyX+6ACUaJ2X
cTn8IQHBIN84BF+J4YGZ5XXZtL07kxotF7Rtz8TVkFnlTXs26MQMH30C561OPpy2
AEKG6e48PmCFV8ZGy1oZGHGPrC+aOiRPxp6CwEN5QWgQKi3G9MBLVeB1I6wJZdS8
ZOQNBOF1KZhow7b3VlFdBunSRss5qr8CTm+L53dq9VipEC33y53CKYEl4Nc7CM+U
/Lf49PerKb7iu/yKHqEtL2VYI82wC8bqKQv22zVgVY7sRb6BrsEegpFS+t/QPGmx
A5XKLCwM1Brr16ASdbmaQ+BG8kJyLNrp/DPagYrhmeiPAmGBsW4rZfhUixZmWEcL
COr3rDzJMTsVYpS72l6O4dOpSJczwe/QLkox0SV4A+nVamFRNPY3+3Tvl+fmRMcb
g7rufIR80HTF160lMa9nI8MGf7cSsLWSeO5JfNWAWt2nFAKD2lYyV9dpj21vZxja
OBBAX+E6mI6nA/+y9/Dr+BrBlm3FgT+yUeYNmkJxy427ZcXrXCLHTXY55dZjzEfu
3XQUDmiVM1Yto+oZyhlzA+PGUMrpCnIumKMWz+y48Ma700kfLr7Ott/KKuC6PPuc
pOomZgKVJk9fCztE5ZW39bUVENX54/gTAnKIRTW7qpdD2Nzw/NI6g2c/tD1S2wV8
5UKtiBXvpoe+17CClgFpQgfQx901RWYFqVdkQp4u1Cu9oKHSPBf7/l0d1/z8W1kg
XWvDKuOT+eNWl9qtAp7XXY5IFl/0eeej3o7GTHb9jKIwawbxjz8Fsli3w5vWbYz5
Fq/VmzQ5So7ShjQJPdcl6rKYNTlJ9gKwbVVtnPMg6rinhwXP93Rp1NSdnbGuAlJM
5UZxixCLRoKCxQFP5lNHZADO7igGhFyoeOOvQJmXG29fkqYukghByNxwyJhFbL17
Q9qn6MRN20zrhhsFMEBaHqIPV8pYgaQ5qftHHfbYYotoUNOJwzOhJbMWxxAQa6Qk
4xckKPq+5O6gjA/IygyGVFEy9eT3/ODmW3QrvLIWplT9HhB3WVAbcVIRtDTXSizu
foUMuHQn5IArAAoyP2gE+X0vh/l34HiuXI1gAJEezUaI12rqgYQfO6w3nyMbVMO9
mtn8J1ieV/UaeSs4Nc+VLu75cdxOMh/+7MdrLoMrBBbZUD7Mxt+31P8Yo3FKJdVr
qhkGESSQjKz7Pusy2qT6KQicBiYaYacNLGBXTE2T8QKImK4I+Rg10/ZsVpRg1UBk
tTwb75+QlegzEki0ofYlxwD/e539YjKRxNSJ5hM3uK9Xv/CPov11HnDWCYLqF/3B
F86z67sXujEriIG6qq3dNImIiVqbMcbPbVKTbB4hfckBLxiHiH1V6DNbdnvRQ541
S1XU50HxVHy9cWUlxyDHYJEppr9c7zrAyd/hPlAaeki8Q+n4ljcQA8e2b1G3PS/4
Oh6J3Or3IKMd2mFoN2FHpBzBBjOAAz8xnGrVyytaEL+UbPy/B5fyIb2MWW2lJRYz
OuuEWFr5kXmefs+cUcRt8SmzDJHzRH/s/leiLz8tbR1jwiD9+ogaRorDZ1NCyMWw
6F0TdzONd/JXJsLvPQ7ysFj5IWHw1ci19IiQ0L1VXTT/rr1hA6RRwSWrRVZwZ9td
FoYTQB6ESa5k/cbKjadhwkORLr9DTdJC6+0b0WhZSk2F+VL22qNGoX13PVdCpNMK
J38/c2NtCdtRlOX5eoUHePNZ8CxslbcLZMzzTsJG5CYgn4zZci4UoAgd6w3KLZvZ
ITiukEEGHijMh9MKR6fNBGX9E8VuQk3GNnmY2hxEckLKe+CqJONdsJo8lqsc3qPs
+saHXwMNtW6vMigT41NhZDTsrr8KFkH4cP3hqTH2j6PY7fAdR83vIGIOF1huyEI1
ycPJLfaZ8yo5IYkKBoBWoPGRM8GXQQQgb6wxv4WxsUVQpaaWeKjKk3OWypl2b9gJ
VIbE8LE4zEto7Xn6pXCGl7CSBSpL+tT7Uvn346r5WXRj0v/2dgup3hDoitbsAUDs
GnIQjq+7FY6C/mBURehejSVXwL06bjhrfTKRpTVrM22ey/rw8ebbdwfwzhAgIN8J
Gl+3Ysu6gGL+e6cZThnxqHvWj3rE6567NgD8PxgkZUxTnMj+JtxuEskbuLgxpa56
qpg3BBrg5iZP2i1/KdLXeMeMjZYVLTokdVjz3Fhc8Xz9ma4uQ3TLk9ZBnNQPgp/L
fJSyrdp/f5h6B3wgetGkHSLE0UDeZRjq4sX85XPhSwAyAKA7Nq9sy26upeebxM6j
SRA1yQFQqMdpNn0r45LpQNf/Ytd4+N8qHfMKT+SDU5CIXgjWBYxJn2NNikh+aVaC
GEUpLA1Odg+GZtihMN3FM2C6ubC7nKErCVsg3IGBfppKE15V5TaTJCt6wl3lSkEd
dnjzmkMVKU0lv6fgIVGsZ+B4wWwOIja8uiVZrGCsHTh5u+Muo6HIKgy/Za3VPlmv
FLfcq9BgcQMAXOB2KHYZTTCN4elmM7Zi1RvLEnWQnPKRPPsK7rpBZR4juEcbb2Sa
Wz0E9b5zqc93Li3hK/VaZ3FHdlu26Tpf0L2yG/Blng91IlEYESbUzbRREkgbik2y
SsjeO0LQyqRplJmIGPO/5wDEDWBsDjvwIV2M6pAQQ3v8vI43H0aEItJBMILGrN2n
kQp0MHY5QbCv1WLpCryk0NnX/xE3eJ17gxeyqYFhMZGRaH3GzmxzDTbAqwKeuVd1
dTAKJ6HfvCfnQtmwRlky7RU9RfN1t0XUTZ8b3uwe3ofCjX47gxdmCc9uyJ2wGiqJ
jgw3UUIpUrY7cQEnstWkPgGHK4xus3tHjwF3vd2nwkNVYlQyO+m7dOghF5BPf8Gn
cquBvk9uFBPFdUDr7JzbAhkxm5WTBkNyD9xZ9+YWRpzzGL5YpSVJZq0RGDxhuxt6
V4pN3SPorqF/W6jz+j0k9KUCUV8WxVFdI+4cLYglScrz/ZkIaUJWvrd80ENX5BkK
hVeNeJVC2mBBZjAgegjLGCiWZkdOp6xQ7gcJehFFL7wSqgo7GgNUyWrD8TPbJfYZ
82zwcbFGRmqiR8CEfhEvsO1XU5fFB1/CKLLODpysYqHc6b6A+2qYIaKsKEQ2EUrs
fFKEO9Z0DJWgyZ/GLFs+Dk+BzhUUNeeh1icH3uhTDVhNKGRPzDZwKJ0qVItPV9u2
Pvfl3vQy3/Ao1Vzm6PYk/lthDzlAe8qwtQC8wP4gO2MH5wctsau/hjDlOx+LiDui
0iokSyJ7hsMGeOLhcXv0SdU2oUk3dKfadCq4Rj29wPGd0sKKpfl2ObQVdGWXRrCT
qgXVYmjHFaP8HGsIDsTl/6ILrcbPILEzofBepwjnSCoPg4PmS11g1CYFnfTNs7aV
wPqy8KH3mZpTlHbjQQTleGyUoL4RW3N6uWgcT+KOux5BnXaROMKBZrdwJhlbn03A
2zPlgDng8wIdYDeGF6J5ZE0nClvqyFuGqYivfTxgn7EPeoEk/yl5sMLh9eA1xqg8
UXVLR65b8kAPG4Qtf5iwuMJ29iPgv7xJXlm2PCFnFcXLWZ3n2afilO4ruW+05rkK
Paorh4VsVR3heOyQX8fjFO34RLpNXxaRkaxGIWYDXJmV5G6A/8n31gjACuPWlcV4
GoSRN8BQy40Ua8YmdMTZIaJb9H2f1dYynUNn1ZJC5NK8RsB9fhwPyG1tdILCSBgo
9vW3gHXbiRgFJtAisBWiJHd8w0dVQ473laqlFnKRkzTcPRMmPMA1SrshOGnVzfnd
N/7w9HV/K3sAgjn9myD0ffqgL6qpKLXr2xRipnrZmUhpuR7EmV+u+HUMTkJQwMpz
86cIg1GAHUoHgUzUjHEACucxBq1TJoOHgYszlKIc4OaC0W/KCmCkql3oldVgQbHq
9AdLh8cEa16EBnHD68bz/tX74Eouc4t/BFmJK1boa9QL3PSQysYU1nipTD+yhWik
fppRSSEnpKzvfrDWFqf6QLfsBdxIxukp3Zhb218o3r/nrxh21aF/YmApdD9WuPMc
h9B5HXdONh1LuGAjN9Jv2GbA9HvnPMoXUavKJ5EkBSDjc8t/WyjU8ukyJ2kAt4H8
CK0CfQ1RcPPPPEQ4RlWHGstdXHmFB+DV/EDtKsTalyZM84BOCM+xD72QrfajaEq5
R0npIXu5tJ4Y6KZ0LLTbAze6A6GJ4Y6ngg+xSufB1G3dVE5Sga8HvZP9y5e6n9U1
NWjfN2c0gz8SsGBCd7hwYnyYEqHnOlotrrB1XRR6gWSPKkFQFaufopaH2Uvt+pS0
k71XsUSAEQBo3oyz47kfZcbaEqEN+GoMAKuFRHK2GDwh2Q+LoEcPGIm0/C0cj3m8
DEdrCja2vVtQntzU1Fd1Ot+WJnOHk/7B42OORSCGJRwliTfHmNmHRYkVH1WeXsYb
X3b/wJGCzu8b8BW2oDnGsHhwwZAid2AHV3Tmm5jCvMqOZqCcXGxoairb8czv3Gv/
SOWQip9fJ4vVGjgl9LIXkKQzJ14yCxGs7U9h4ci/8u5A699bIanHqw66E/g7Ffsg
0mB21q53+X9aiYP8JaSRlNZj5FMXTJ0KhHHx9WsAj1pAp6f7NBeT5umQQd3RLUWv
lV7qgwPFRf5ofclgudkKnbQ2zw7edLXTFMJSpHyaY/HAHtkJWLB6Bq48eODoXv19
EEpGoTieMCJ29PUzuogs68xusJXhkENnXIu5MUZEuhgvBaBKUZCoeGg70Dk5GPTo
uO5gFMAjt5Z6q/nCpAPUslg8s9CI/yPvhjMeybJ3tPJOubi6gtu0SO7GYf75ErsW
MA0VGLAm/3CPwT7HstH/1l80huz2wztFT73Ue7Nx1WnYHKC8v+PH1g1Hvk1sdEL9
Bw5BqcmROPqD2WcNde7EdoO/EQTl6nhv82C4GWuIIdUb8uESsqjfOndAQEBGZFCF
25ltdjX57NDQNm4BXmdqGbaGjsnd1oe/Y9FK29B8Ji+qAaSsYNG2KR/oi7yJA+zy
F8uL1Nciq3dBUKwMz/cTCw5nqR+I62X6YNsa3J2r86YxjqUvTcwmypcDCdmlz7PV
MG5xssd7VZGeRtGApoSkCgaOazagsWZBr8WtqdB0sGQT7Hy0aWI67hUi4K4EJD7f
XO0NEa8SpBVHShADb8RrnG9UJ2RwuZgd0skzY1HXO9ZV/DGsWmj6kWesN4+If6+T
rHUDBA0JGgSQmaXYUg/anSn0FKKGWrJOQpB/7jLBktfILC4A72a4HK2vX035qMqC
MF1G8lO9CUAREJtuGJnLxwNsKYF3qJ3ad1zYA2Hh7HqERmEnx0XENbwBDoO7S9Tp
7aM2ezJAUb79TGunOdIz6np5N15Dx4kAFrEdvV/msmckyKnsXqsAX4XHT4hAo+JC
384zuFFIiU4HXrusOFu3w7SR+kJrnOdLdg/U3VC8H42NGVXtsigeG7ASYoq8rIY/
7ItYBsNdcitd3hiNV6EZrHDJS9a49car5j3hA9Eai+i3SiOTKaCUOYiKeCv9c//s
5mOYdTTIzCpL2/03PAboNtLLXUMP0zo2J2kJb+IVpN+0ozWvmtNMegQYcxtpndjT
kokgYg69nwx1ZJIDHECELT2i70XH6vvoZBoN/TaE+/AR1gMVU25bI6rJlWGgL2n1
YuiPGgYTXWQUzrAgs9LY/1rd6g+YKMUXogLAbittXralyE+Fi7cpIv5R6bH9p70m
w5kdmFg+QZDu089YSTTN9XEDy6ihDu0v0Vu0NNQYeEzZeWms7IcuKMK4AU7YWYPD
wGIp7Mz1LKggWHk+uvgxbkZo8YDSUJ+TBbIZMyr+ETxX3xzN3bXMnTZQpcnslGpY
UA7Ocw3uqnKIrVol0hU40/x3YVmhk+v/xQhR+mPFoBEtWHnOpfMO0jO70VY6uiem
sibQtEHfPNmmdBsn2wVVpuZLBeMg/mgx6i+sXlJ3mJVOY3t/xIAWPnMxp12eaVI6
So90l5+W3x0ep8746lM9ZxAE3RT/jlvhwK+PcsPB2h1NkTXi6pzU8N/VL4GKS7We
7UY00klnnn1ZP4gFj0r5jlom1lQ1HvXm+NPyAlnQU+eUco2YwNIfgmEINbipNKD3
DopD01ym/4QNnQIg599WOy6/7Wfy7+A7cfuNa69nLp7m6c3locbSfusnyMk2439y
js6eJcxmFn4VGdFUrNMao+Ww6P7+n0b+iQUINkYXrGbvezxd/WhJSy8cHKpDom/g
7//Ze70mhW4TEMxOkDsgtMfDYCTchZjkDZoRKdz+NuJoM9POiBQYta6Xke/+uDkT
W3ZujzpwNx61ddJ49CR+1ke2JsPvV3n5rRLVxZOa+v2AtSCEhVW3BLRIUAb5CF7b
b78WP3JLLrP3nn1LJPb/3S4w39+eUPkzx7/oGnLQfh0d84s7DP0ilT0PesJqXM+0
tgrCcHI629NB9vnKgSN7Ia5jaG6CQqIdNAzMI5zCDRK4u2YFKFrI/kbNq4E4H7Tt
3aZeVtU1WxvBroPB5VKiXWbk4CPP+fWsMf3wvD4flJdZufL+OyQZ7OqM3z63f20t
fCjyA2hplxLXA8V2NKMkcSD502K9O/zk4QTo7g7XavSZWUsEuGUohlcCeIvISmPW
mECPfhjBF6SGY7tkwUc1ti/jYPfGGjyWUALSYGKEdmBF6NpBGfOeq/jNooY0u5Z+
ufuoUDrOCkZmVUuQgsIPPZpU0W7qpEiXiykolcHI0xCCEPzWsHoX0BBkyuNkiQm7
wOtZpmNgmPK3YqmpO1fBcgDAwsRtjAHIgDjHU+cH93/qJj+tZlb3hNRFy6gbwEfw
v0gwzJM8eHHPyCe3Edj66/ifCRc4T6aWLlwESJ6mYOQ0lO7Hk/RfmzbZ5g+WNmSK
aOFtB5bDqelduG2n4QU/6DjgT1mPePhTUPyZMgkayXDRIbMz1KxTdO31QbInuaRu
8G9XGoAZZud4+dfiu2++FhXpHyYWf8eMhedTrL0HHipxVF9n2HD2JUi8EbD2ikYq
j5g9PMYD5J77oGsq2AD8UQ09JojCYOE4tstV0zs6ZD7MLBcpfp8Hcp35Gyw5sSQz
B8pgbQaUc5gF/el4ESxQ/xXQAh3OLHsCLFWnCea895WFSo76NX20A1EXomICcs43
DX0cGdAfcennRCzIyv0w3A6o0Fh2Kyp9Vr19P00vqbBM4+HNXqECwXvQneJ/mIqh
IMlxRjVYWm4lLmHbh+3NBM7Ti+q0P44pZ2dyg/zGYfGAAuge3fxjlKcfTaiVUgDo
/auzkKNEMsa9vR4x7Qc9EUsefZtfrpCQKtlkTHXohRAiYNJqnHjHemp7F8SfUyVN
obkJNl8CsaECNjCrGRLxIgY7++f1vE0ElGGR4HAY39gxRbrch3pbVQ/0hGW/n4Nr
ib70Qnhj49Z8tsz4tCE1S9Le1ksIGk5RCUBHgSAiwWTCAZ25FgrcRkGz/3YK1kZy
bcA1QgVZCyNQDSJh93845k2txbqsGL+YWQourBjtH1/rLZXaslKVY9BnnDYb/tJV
yll4W/KSOq+V0Pe3HuFNJ4Uv2JcCrIfhXevG85TGSflsEIvtUtJZ9CEfSUKxz6Mg
jykPPNNCzAqqSWMBjw3mdTJ04wjwvgoQgg8DoAkUSB4AJWwmx0NwBxbAT9JHasId
K29UD1pbZXhPtDmNMpL+ZVYZ9vyLLRJIoUTScEp/mpYNdQnLpxwfTbt6ywwLrKZK
IUwLQ4dH/tmFQ120yHcVHc4L/iCizCDaDIvvokKjEV6+dxhFdIdHYjtL/xgoczVs
tQYzKq/mIGRpJptRqHX0CFdSw5jNWzn7yuRT6K7NTbbt5xv3BqctNDXvS1JRunIg
O6UdHkRKk4fFowQ1LcfIYbpWtwQCjo9baBVG64H6Ow8ph7+F1P2BZg4jd0rViJBt
oLM5OXCMwBkdt2oQAzWYRKsH6LmdMlK6URhntXFnyU+6IMpdPtiFbhzA871Pq7YP
lixutmsbU97584GB3Oa0+2gX8nL94ccoN/ZtMAlSu63QKrb9EbT/liZO7AfJm8v0
1y6QQWfwinbrt2+NWmEJzCciwYtNhVnwrKM63DquH6ZXQHZquADpIXwVnQA+ytfv
LTZ2sxuL+Ja3AqxDSveBp0SQorbLK4i0QYntRlYLfzTvm7wMaSgIKToYkkWGaPOT
oZlsKiy5x4zKS30k+VKaLCbovseWInzG8fRtrA7Ka+Pk8KT3iz5t6njMe8A4g19S
sP+0b0BX5iftQ9PlA3bljVW253eAzMFwlc7liTjbGdpilqZrzUSUs5HJkZlBXH6G
Jl6YYbV4ZVyTjdnoWjZKd6lvrl1c9S+qnCIusez8fa5hY4GgUaOzzSrFQ9qUrNmw
N2O1nfLt7GgYPyQQgydOsy73n78FEcUaFeD7zogEFzDZY2BklPeZ0NKof6V5eorm
PFO9/+aiMmbXzCCslvXQ3PdfbIk3HFCnbZe0pUXflJSMybQAKkgplM4VITYdAAQz
ywur4FvF1z2bClHabm2++KiwF9suXcqezLBW379tcpRKapiHWw0tPbA+MyFUSrtG
FGbUXFqErJlL1LAgxoqARNJzc4Hv0yCtKV8qMv78gwxwAKDmyc87c68sipDKdkc2
QDQ0hbZrcuWf7bbM5PgrOenIHp61rAW+jqbhmmXgZJ0AFiuxwP3U9HNi+pIcQgrG
Loqzur8biSOlHXzXVYC7YX7t9TxRUBWZ1J26n+6pLyYJe/WLKYq1LasdniqZxLiw
Jrqtyi3mKB6brcBsShPND4kn3V6teFimoL0DVyajS41Ly3CriCMEwS1ojtdZD0Xi
iYQZBwF8VFk5q0Yug8fFe2PtjOP5iQLoyo3jXsVK65lshk+X4HJPsaBv18QP46tj
VySLc7WDP9wqShtWph76hVxsRxioWfjuLox7X4vdJuuLTUFr/l/rtk7ILk5bQJ1R
hwg0J0h5aOnuMADsuK2ny8BWB1eaFQUW45ojPRAsPUdjpXje5qr4Z+shZO55c+50
FUbUWXVwrpMp837qtqjlu0Pwoy8DoukUuHIiJ94sxFIvx+QwYjkxarlfV0PxU87x
xEJePZtmgJffhOuI0kT0SskwFXhnu2Zir0FpeuViXa9MI5KqOP54HUlgkZi/329R
6V1V0NCcC7aX8QcXivi6YWh6TUskv90AnDGfnv1XgOeskBX0W5h/ZRnRUkfymTn1
JjnfLkUqfVAlzX8M9w3+sMa7T+926MHlwqeiqM1EjasqPL27z6XIIlLYGHsN/JLx
Vfi1UccmEUuWJAACima6YhowcfBnQ50r7o8+zJarrQhiHgpZbvezcVPthjjDJjj5
Rjdf3RXwXuc2y69D+r5w/veUAf7ZJCebprAjUj4APY3lHR30I9JRPgaPW71lTJqH
EiAbi72FY80oUkcEN5CZlI1HBlnYAyVyUprTCtl5tw2Z8fbU0EhV+uPTpTomenWI
wmkYgdY0Df1z7geNMDoZyWnWnFpDTAbCMaNK5moKx9JKnuX7w16K/11HXrtOPJKq
KnlSDpACwwU+tSfQZ00aU5RDA7sj3MTdV79jWCRDuS8knKKaNSLQzV7FO/4my/++
BHaV6aOSO+1iXugwZbbnnJwo2hsnFdTZ28oeHHIrQAuo4FnsGudLZtOQYrj6rkjc
x6xNn9O84JvjIsO8SEaETylhYqVqpIFENPboP29UM/5901a2KpAqhwGtLOp5hN6k
vfBdbWgMSLWxO+f6+TUIWYat9x2Nhyt2zewdaeRiiaWlpYzSCM6XbWp38aZPpolZ
n9l4dNq9CRuDDdJBekxsrl4oFqVgTKnXIq+6uZ8bpfGVLKgCjStt3b/wk7OOurn7
PXsYHj3Xmt1I76cVnjhZGLDYC1M/lu633AtM8lF26FeSArtSuzvNYjpOirHlA2Eq
Zchs1jg9jhO/LMmNvfnG22oUctPfCDzKHZwFDXIWJ+VI+l0ovbWNs8yvxU/lwKj7
ijNGIy4pBtWH5iDCWcLCZowErO7hOuhz+QLY13FJkSfuRkjrPwONv2ngYOXYn/4N
RcbXMASC0PNz6NUQicrui9JBg0Jbbskp9RsGzkWBDU66ZmuLAuFhyOWNyialuUNu
KtDK7s++poaE4prUgdHfT7C9aw5QufDLZUq0q5k3gOdwYGl2KyAZXtWVy1Pp4muw
2TczRD4Y8CXeYlUBkJmEUn6hK5PZ9oVc+2w5TxMTgYOB45ve3+DI8bxCZV/2RLHR
vSbZVSg7OqY55FvYr1PD4X9L4wlurxBe242PN8hjh/VfcNWcSZswSKYjh9QTfINy
nggmf0Ktcc0/kzEokrCx7eNWhxrV3D2aZkxzk4xQ6ILDDGoQ0ZJDoCXm85rFQNt9
gsxCLjV1E7Iglf3h5hAsQc4S/cWedCU9liBdkiDbW9nA0/XgWqBkYIN3HrZvkk2J
OGn1kP3DER2eYSlxGRBoE+PINljuWjXBjHurEQVP/vXuPFcaJ0Aq6KOJS37cvj7K
br3EtYLwrYGfF0cAjCOCpX3JXOzH0Rj8f6cqSh2U2vhfrER6a++7lDjB2GRm5vUG
Z1WUdgH39qpva90RMzY/F310666fdVuORgHwjXYHUVAwsd5bhbW+i5xs+k31wbv6
GLIPy6KCpmGfvDYHy77Tar0rryw56JcHLuhsXchTDkfqJyaMCyA1qD2BjWY3mhsQ
HZ/3IAsPC0OTiWVqiz/qqcpVmV7EoybQqt4AnRz4N0Y686okYfKJcfFqlZDLYCp5
hVcrPC4KSFHuvEAMoQtVljpX+XBPNV6ziLw+/uHQCzScA24uqOaRcdTbxr7MX+Uq
YWg4OZTGoq74Fyo0rSCqk5mDFYZEQF+eGqFdxR9wIoqoQbEO2xA9Oi2gP4sfQ+yW
kfyK1AhHJCyvNwoCRwBQPWm9RJtTuo5c1jBwQwExXDEJxKucRrdFwXKCYnA+kql3
3DTzfAjht/d3p/4NQQuCZT3tKL8fRYHx0I5fOO1oVneyKtVevp/P5uw7RFVFdJFF
oq3KH1iCWpZPV8icWivroq//0uWxySy2QxpD4BCOkOINQ6w0QnFIYjI498vUPB0V
n42q9WNHJ6HsPBsuj8ddyU/GgFpy/MjSZtufHpwiqp8+EiCstf1y0daJ4KpBa2M+
b/tSeBJaT4OIMDhyL406PDoxrnkI6TIu0XCRyGG9tJe+2x2KGbfSeeuZEENl2oiq
AmeoWvrEkuTk/RQWT+PjrDo+Rqu//NILx61EFVEgMqWRTYd5UECyCfP8L+7xI6gF
AAq40Vnks/klEnJ+8E9kr+u7R/AOyOYmjSlBFJnYX5E74/8SMW8Qd7a/U75xJRn0
5UgRGkwymeo1OmCpmiTl63EzEnx3nuH/MCG7poRFwOxurlC55z0SuQOfwGohvuSR
ol84l8WB6frbVegpD464QpAP/jsBH+hnkufTRclCQkK79FPekAwPVlGOg+9TXZND
6u3nmemnZjxFYKR0KnTu6vtqc35unbVLSA2fO/7UUGd7SPR0qKuva64UbgGFcoB3
4TdDK09Ax0P8JU7SAy90ufhggVnn5un5TOuk3Lwf/Ahes2RLOL8frTO78zftIgGY
mmlfHFsNtA8ClZpqoB81cSE8duEJbTmU3tZZv9EG0yKTVqvnOYD+w8DjbS3OYxS8
0sn9OPdV3V6C4TBZfRjSclspkepYyGu7LtXj21CO4AvKfJRjZM3icTPaSFGpy7k+
rSGuXsHJhXM2Fr0q+G9cxuKjcF3dzMPge1LJwQj4a3YCzFBi227BnNBalGLomsDM
gbnAz4i57iorV91Ma8U66A0jV6JRHJntwFuNZE/VCpOeKCbGZGxUNOxRE3bE2Yfv
OOJHlxPbVOM4q2SoBPDSMxlM3M/2h6bW9eb/+/ht36hCx4/gttMWHiakaNyf3kgI
N3Bwq15hzOZz5zDO9KZlN7TACSZKc7XWXot0+37rlyUP4x/b+YbqZfLbX02+51TK
eQD+stvd/7+QBXpF258JZdOij0x+XCqgCLWYvxhOL10fRsCEEDqNgJwAHXpKZ3Hi
J0ggDo52TFgpLYzkrYEW0q04WbqOrzb7emMH6olubRc4PgOdNvwR5JFCHWfjOS3w
wZAh5K5g5SA2V9kCmnC1I/Ho7Ds2Js9avj+ijUNotiDWmaExwxDTGg1WQIn0NuRG
+Ne5R/U83S00k+9R46Ks6yyd9kNKACt5DL072XaqPhcdht2qX+DVAAym9n9G847l
XGezpz4l8UZxt25ZTeIYs5Sxi3i/hBwjt3HSCO/8g2VZ2Uiy2E5xUDjeo+bjwKjk
XlBSW5Cd5093ZzjndAVO0p5C2nExbZ59Lzq0HiIphXfH78lBE1r+aF+UyHidJPGz
HCO69cUL/EGOseSwWdcq0Q9ZxTxgg4O/9ydWnex2M8XIJfR930c2qnHp0h6ZlkNk
a25SXXd4WbNK95nYR9GlVis7Fl/92IjQ3ZGrnGtVn5lqtv2kdQ6B0gX065jxT6Yd
Mxud31YnYLLLM9Hc9waE0rH96yALheX3DxFXAGAi7dCfC0C709jE7tdrQRYva4u0
vAYMMW9MPblPkCo2ViXkATFCFX144Q+k9Du1isvIf/GaRmDEu9AtK1WtUTZxOqsE
PILid+XGOyTLDky/m95Vso8RxitamDryWdhXJFIxKGDXq4PXi146wqHBOUDHnCVO
dsgzZzdbebv1x2iGzAPCAQyuXzLKqoGv2B1mZd0Fwqsct7HK/Uzysrsb97Y5Hgoi
Km1okEvTNjLmmLg0hFgc0yhO/fTAGbbtyhIJWvSwzXW5njfxqpqQUdu2osaXD+Of
ZQ/q/Bn0bb9OuAm/wx/BefuJqB7wWm+dqWz9g48F9JsEmRXV6Sr2KJkmjctRD9Re
tHC1KNQFB6elnlRf4/RWxrGL9CFlEHq8I89qOuV4DTnaHUFXDlc0zQkvhkP5aTD0
3GOk+YF3AP7mVWWEonqtPfOSiG4WTbVuoPkSiZGBfc0KWSEKY3kCvQ2P34Nx3CIX
Lt3sbaJ9YOTOaGGeN/TyU1LhdMNvQuizx3lUJVNLbQjwke7WoVDEMrpejhXndpof
G+GhNpjIZK+17yshb4T13cPfh4QqtKxdBL0C7AA28t3DHJKdc3L7aEHh3t3Tas8j
JSKmIwRTwwJMOXni2/tZZy9HcR6Wl+2ZtmNJkFAcR9FGvltD/dafhr13SMZNrhiz
ODcrGFBgimS98IaVh2JV/IR+byxRJmRHIbvzx9zevmwvOCMOAf44zmbz7bch8xxC
89yESxtgte/bePuvF+kERMd11LOqSFLBFTRmqyQ5THvJADHMZcp1+mYpH/NaL7M6
wr/Xe4vcMNOSClVLAz2bVwY4ddtyFWNFLAQ6/oyKfog06o59s0umJx1vxeGA961M
KzidxbnBWLpNaAaXQoxQ1WFEAJazb4dPjum4Qdj5LJJhR/3y40izQG5O6K5PlM9D
WL6hIU8qqeD314xgRY+zEnOaXFf9XnzJ5mLHA4pVD3Bu7zdIA+lC0UVM64E8Zh3u
KhPfhL0T0vj5wpsLduYOfjxgjA5z8pizyrIljin6oVljAI4d1wesy0OGacWxnxnZ
G1OG+4XvjKB5xCjdEPjpW3KMMXUqUgfBbI+KRuonYUKV0eLhfiD9DvNOSUX/Oxum
gTBUyeZ7zZHiat/Zkn9dsghPLAsJL3s1cVlmlzavV5zKJXF4MumuxyYzwhUy9Hjy
5/qN9aTXEKacPsxxWUnrZm1/VstGsvzyc7GAv2cGfWuoiWaLVkC7iDd7L2QC/gVI
V87/3PSEm20rm7j6+E1JLuZ9vGtlLPu4ZfZSTfIW/5+16JjOXt2KZ4049PBj49F6
89fPdEg0I0vXx1Ii+xG8yEaMmnYeRBiMH3hE/LqlZxIxddxX2rSrOSC8PpIFde5X
2gpP80ZX9dXgJnM+6KUS6h2nKRN7zMouyLlzvblmq69rngrfxDaIGkhBtR8lOTdB
F5LYhDHI6Tfd18grD9EpimfqACDRbxQ9VfhtQIhN5DECtzqyY/vQ8YFY04e3YI42
UwhKMnBtj6t30nCj1xq1TmH2fBgHtnqMM61wMbIDB+lpP9upcgkpR2jIRXFfJaSD
JKlw/YwkJHv2i3HXulEELPX9ahBxZR30D7WhBzclbmjio7ykvoYRJfBHyM7ZaGd9
ObkmFQpTXWrxwuJ/6yBMfaQurKk/QLl0Yf2aqYd9N6Q3acVHnVf22QgQ+p2x3jMw
HQHphL09U/hiAxECIxY7K5cxjTWKVcHITq/L1AHjrPbHjw4mB5UJs0jMdAv1s0Gk
vZhF5cYBzQWqOXHvG3QHp9p85VjPf8PFqSn39Hd+MceNT6LL9HS9cZFCoyhHP2k/
mx0XjXyp2Et0CMzlR4pggW4e/39WejK2gE0ccekyw7F1Dsz+BJZtKY+vTebU45Lu
OkAaQL3MVXUo5M+Y7Ghxnm8uiFJeRfWQ8tsuAAHBaKlDdkGSKro9S0OR4kCtPxD3
oELlKhyFDYLS3HLMWWW8qNCis+do8YIhz8rpXnHa1g31NB0AjT9gQigD395gDeGX
SuMkIC7AtpBHXx/fI55NFk/kTx3SOeQrfNs8ozcAHIkS41cLhPYO92lmBt6ENVwY
jmDq3Uexd86U+2pnr5cyAwCPMZoP41XzrOp5eX0hPiY6wttpVOmhPu+Aexgheh/X
EtQtGuUGcym8GadrFh1JO2/+FV7bNdLgallzVQ3ORGKg2yeMRnWQWK0n2kjdS+WP
6t0IOSUOXoGYhLXGAp5PvnjugHdd4Gmg6RQBW4HVwuEP1UPMZoQVZXfGEKFpjncm
Y9PNJI25PxRWiBZHR8ed7QwIwLEZo15Li8f8vYYtn25sPufbK3Bpz/aYUKwxuySN
gWIRRZXE8tzsxWGRubr3M0MYmOdsXecpXLvixzAfBOGolZP1qSBcwEQxqH9suSUL
kNr0ymAwi1V9mbEcdzgqhwt/aZbThbCkS1Omtx2UkajRmSmbMu5YjxG+Nkx5iOsX
ZaLNO8Kr0dMCueW2HZ3qtgiOToKBKjnxOINxyJNCkeDWx2lCWYiXdlKe9iDXl5gI
pr0g7KB9D0zKwcvaLXxMbbDEdIikzo8mkAiBCddI/jPP93gMQngqrZZZ+GacGoyT
VPTeoMjUyK7lgwqTn08ncY5D88rQKUGTjEjxPXTpoWujDghX/ciR6kwSGKAKeh6P
U8negpfZLcr8WLO043OfEMS2oFHHncFgdv6EXfy/reM3QhMh/7Tty8wWe+aCl4FN
QcWHrr7HUNYgRu9Ty4KiNParjYFO2s5Lx9+84OrN8jGJ9U1XL3lvISAxZV9f4nob
wHDdX2rZNAlpjhLOXJQga6WTD0rJ2kV9MbEuLY6X2CoIiH9ZgVcgG5D1QnDiYAcK
iRTf0yo7uakDT2Fxz0doIUCw6Y9HpHuseKFbwahuFPJNnr44snrCRU/FEL8lf7fz
Ylb9ELgrVZd082zrTSC6KqRaDs51Q/w/6Tdc56GHImnmtielSTP1zGl6VpEBjzmB
jLgKze065sUwevYoyVYDf0HBRUyiyiAfSWP7kGQtHukz46j1pyAhAgHhC13Eohhj
aHcqhA7EU92kV9VcGkwO6cT6xvqT0L0r+KefnFbwvjBDCIk1pf18zQMOg8gzNmAo
QWhEGIrlyBqclYHxTtvI2OcaekYbFb5r+1rgRVTh3aYJMQ7BTdq9ZhwHkjR5Nt7u
8VsqUDNkW4JFiwQoWDqqvh6dS8yxmRAxLfrW3zoScRuB/rtpQdBJLSyZD6lPDdCO
o/l212E4tUsCcMqx2B4BAa9DdcBIdjkExsiUV3LOpxCU6AGmncuI6+yEmR82l88F
o1SQf+1cBhG/GvKnvlPJZUnWUSob7lKQZCV0V7h3WJ7cOF1w9llBKfLsguYKIipp
mcV/VrmVUvz/o+ngieiwaT5Hi5D6hXVc+2dzacaPwfKtyIwXkitn2AVqb2cz7iCz
xmC6z3pExX+5+meurqfhm4KL4KDhHKYzztWPCJei5FeWADtYGGmede/xNXYDjE1n
qlICJaPYkW8qcIvxzXfjSi1jZuRfqZz8+pTXZYltOkH8SYWXSvmfwSXmx+afLAHC
51v90XnwXyRkPB6Sw7nj54xKhBGiZeyONlWn294GLRL6JFAhSOlzZ2dMX9Br++X3
iqvjEO5IbWLonFOd6gEcCE3Kz2vGHySlqJu7mqHmY1XCbRtdf+240sm/lSF+aRQM
uHDDIT+8mDFQPLWyXg19y9L72KyjYIw5O0U90DuO/Oobsx29TIDAFrbM5RwfSJKh
Iwez/GHZ03C4rnQyH5tUpCmO2mMgWhHqVABoFs2TmrXK0SOWGJjlzY/I6DUSl/O/
+n/4lX9bNzVTY4Ue7x6kNznQvN/zq93TIXAFQLBc64EuEeKGUoqsdkPf76Wkpcbl
xGUd1Mo2raMzISMFFNo4nnLNLkxk6Wltpj+vcmyUnn3S7Ky77I5P4A8qrDw5g/IZ
5qkWM/NJZmL/p3LXLHjBxMr9spWsizwjrkbykKEdcCn9BALBpVS/wNrFVm5P/5ud
6d9hIwcNs5PSymFpFAC8lDb7hGROGDZXjnsERr0PLXrZJwkkaUH6KGp/j5DMstNF
D8O/Nm/7VJyqxAegLiq4yrowz1YnttRGryQFfhwd368HeaXYhL2URv9lxtQNLq7I
GAc91UPUVii/o2EEU8mEOgQeHiDsuuBkPjmkMpWUakd5n/oC1HrbbFV4e559B5eI
NWtLEx43rD4vsNpHN+KKL0ISarEymL0fBgiW+vfdLzmKFyemivVOwDV3BlVzeuLk
jcxCl6nMfDi1ZwgHP5jhmSJpohBiFCtTZ2mWsa2wts6gfAWDZkDxNwOyFfvxwp4W
F+k62OIApF7fgDmKuFL/v96PWoAVc0tRgz1LR6Oz7prkVy5NnIO9Xxu71UHAPHeM
rgHi7ILI2XNgGh2b97CguPmXYdHHCzk0rlK/GXWVNgt9IWenR3A1tHhPt6OGico1
wxCuWAP/LXy8qgLpevPj7aq7d+r5SeTwZYoioWjHEE4GoWZVeftDOz/6zGOUEJU6
dfV4TNse9csLRUv+mCwUFPdmLlPtMFKLL0pvZRkjtp9JP1MZwpLt/akcixRazZ6N
9LUpnKBmkWNxb+zY5lpp2pT2pnLl8NIamAxGGsIF6JbvnRFK8WsuwIpzFe7ARQeQ
qxn90YhVRRt28HapsSifstr3/EMucEtnOiqhv0eBQpx4+YhBIzIV4kVH9kBMRcoD
+T8qhVlubuSkJ6BWBSlnj6JdUFj4hy1YzCqYp2mmqlYflgej1/H6EF+/kF9KeJD7
YCdHWSKuBDskDZ+OLi2HCpJlYLOdcRcb2id60uZYvBF3PPsa25sZNQJzqZ7Ly3Sx
fPH8TP7qX5f3+PcYHtqyJ9tQxhNBgsTGGGG7tu1Mm8zdMolK/G81MbqXYhyy3mJt
70f7zmI99IlboZQIRiWN0wNOxJrt5DSGD2tjRM5T+NitvVVdqocVJlo20XI/fvz0
C+XQmjXmppKQbv4lUDyUQKNDMnyaaydDTpw3suVfXmr76VssTM7AxJUVh6j7hjlf
oSaWqSLYsTHGOUqjPiBu2K9jNVp1c9qyQtZtj8FlF1XIun7A7N7JC1+A/cb2YANP
5taYA4gkGtjuQOVqHLLA5LWn9pawT3nL64x8eUiDN3o2Jtp2OorkluY4RM0VgO07
QzR2A3fN/uB9h9TtDgD4yKx/lOaEQUPX2dmeRrF17pACmD10i1Y1id0bqwpXbHxm
qf/QLudTSbh/yErFlAebUwOd3V0SRiKBB+4bKy0xGQaD/13WFjMVpY0TCLPxN8WK
W7vCFk8eArHQoteZdW/79kkMnjfAtzydaLOcbnL94m6Ov7xcCkDqsV/DhrpfntID
4vai23Ubwd3ZLRm2rdLUqGKrh0jMK222l9dEZhskXWI39gMYZYSo8kt6JDPhRH1f
oDqSt7kDvgg2mfQMscokc3euvBlypkxRLLI99tn7JDwKcS9rx3N3kiE1obQ+z9/v
JxPWY4zGhdIswXoSiJS3K1azHVOvhDnz5AeVfIsYBX+2mTsvZmu7ILcatKfb3uYb
wLkYhbhiaTylT7srqfjJOer7LT/sOqy/G3azlpDPFQi8Fi0C7kd1KfOgFgeny1aJ
zMO2t/OpjBvGCNuOGeyCzu7ls8ObybtuM2KlyQ1czR0QBj03IyPz4vzls6vGAhtQ
sSdrhCRj806LAAk0pcVI1dLCioykPFwSGWhCW8/5LCZru1LPmZPTLeZaFaO87D+M
MZB3YinSadzvVqQOI4InNnNNf7KNyFP8GAV22KGeT3qkvXHSeUQGcGBdWk0LPtY1
Yddg9RulQOFa7E/Ccyzdn9CfgjNruyumTqSMdGUp8lv2csv707n9XmLM1v+hgUAx
9/3f4924f5omqniio/kfCmrQJ1Hyhn4TB0qvZ5sWti9X4bnoF+cb8GQlGlhsRwtx
shybkMclKv24XwQ46wTMOYW/XDgmPUtusT0tEkMvZu0WLd4UatSk75z+w4ZyQ63X
OIv7ztKB8uLr7l2VsYsKicY57oDK1wzzqAgzoJg57I7gH/UH2dHwPn/yysRnz8Uj
J52ynLFNDUT3TQSwn6ZWRP8clQ4wiLeTCNrSRsgdtLSZoiLXPL4mhNYL2nx4IWGx
YUTRlOAlMA1cDIFvpWpi/wFAstE+783g9oaQW7w50O34AfXYG3POvvg4y5VWvFW1
78D7QmoqOfx5MsdX9rWlRLV9NaQzjNV43p134WEBYNqA41CwDNZToLKdqCAvcygp
LmzfFw2sOt7Nfff+Xw8bcyndhjGlaoV0FwrkFlZ6OdS0plEN6ZM0jSSSueVGl0k2
fk4jt8W/in8fsnrmdWtWdxNMolPaerFQFVuhA82RgaeMiKSud5D6Ua9x+ZTMkjaw
62vJIKAr2Sgi3y3ilw44rzmz/y1mwNEjub6mdzhRZx48TPUaSdyaD6TluLPGKyAg
cfD4UhmM8zeTjpdQxPIvp8sOFo2MknHMcij2E+fhaoM1QeOM/53JSsMAaC5OrWYO
1mgevEKZoBFL4qwukvsPOQjc7Ns4hVvNdYpeDRg8FqpWH075lmMJTS5iYi20QrBy
xLVX+Z4qwKudSj9/C051s46Xli6AQ5vgH4loC/nlDYto1LQ0Oqb3/qgnbcDD6y45
fY1TCDlwYpE6LixlkBQzXjx7cj+pCZ1oE/fkaEODXHnwtjhXMn9SQuqouxaM7kQf
SKfgzsW9MHMZ4ZyriccDlrfi1yA6PHi3Bgvi6EhX5svswp056OnMmIPBX8xgpLfo
wDvJD9RjerEmYL0wTV2QYQrl/6LFy3ZfbGJ3BtDJhFDapzz1dTp/luFZpXxI9ok7
scGur+kMFffO2zC0G0PDXP4SFGEASDgBZlCWwg2P6mTpg7G5f9knw2uQgTzcI/a5
zh294cVuyjZ9jfsk98vRz9SSExCUmwl+RL1kAjNBzX6nZk3MazC5sL4hZq3hDRzy
Rg9Fzy1v4RCea0dsEAgvisubtN2w7EaJrwDKDKgwQ3gKaP95dgBL7GuG0qP6as3d
V5QQMPUjDmTkF7hD7WXy5mk1nvwil1+HvrM60wIrQV6LXf1dxCCw4WntPkyxvy6I
PufCVUESOBdJdvmz+LiC2hOYZ4vhY6qu2UEmxqI4N8wMQoUVu75oGFLSYjdPJlup
dbNxBUDX9wCxoH5zJmyLzWcXSGBwskq1qZJ0rwhsoj13Tk6kUv5FHUMhUGxvQZW+
0pKZ3rFQ4l2U7MCi98mC2MYOgGnQCKRBhV2PJ+QYra8cFBaSUJ3y963WsxzoprcJ
sKdxJosdDRaBT3pU7sMIbiq/D+RX2FRpRxcjsVDRK2CNrgLai8jJ1ZUjl9X4O4xW
vsrGryIW+afuJ7w3RVd/Q1lA3LF3UNrP8IxIxdUquhQJlykGbMbgNEEsCwBgDDnK
k5OkUbCKANYNUnJjC2K3qIjz7OONJ2Rwm07K3EzVZAIdccd7kDDCkPoOV72Ybv7C
J+efXUpfxExmwJMmqPGEGDtA0NLMfK++GF+IqpH4r6SXFgyEw4G1vlC2dbzw8nq1
2ESMlx9V1Bs6Sz3f7lXpNttSLP7Q9c8X1wdk98pA2x9mwoxKNPx7Ck+L5FiyAt/k
GO0IEnPvPnBAAU2IsDv0zvXdukHOOE68wUZN+9Ov2MH/e10/dtWz1RNMeboF8q/r
sQDYekGCfdANfhFhUsWHYXp21GKvTAJ0bGNaLx5MUKbSu3sHkrpTKFD9TnzxMefy
AHs5pEv4O80N7U9E1Bscg7eREtMy0vRKiQLbyUPwXs61J6o+rZxBBsSbnHigJQ9K
7/7vBrsP5FVQzB4EeoVkbAiNAiue29ArxemNCbVOeuCYRItb9ec7kyBzNptYHJG9
ssZP6Yqwlq07nLO9zByorK44g8WN8MTdHrUko2SKaJdDYEZYmHZn78JaboZEx0ne
ChKEs9nSmd1qDhzg4H9FpIJ5kJYrGWioMBBn6a9g4ewwbzCEln/e5KpEq3vbjyGB
3J+jY1BCa2hvhR3aD3RTawnf0BJO2j80urEG3xGsLxBSwES2JRU83VV3/DqqYGUl
ztZrkG6Ymh13fxjqXBahp9W1Yb1/pVLSwQD16YT0BBED3JT5/iT0FBQgoVKipwMg
zHUVgSJyn7pSfsEovA3H3uFMOjYYufjUqBz6Ouxkh42xqY4FpdO6gMSruybH6ZF7
TI+8zWzH59pkgoM94onADXXeKDZ4SZRw3qw4OYHG3jntBkGoKfy1CHJRbT4bz2ot
oLmJr5k16w0qhpV1ZEkWNRybRoPbZWzSwAoYbkIJF2gFfRopaTGH+2OSD4pPbsgQ
uf86kHCX7I7GeQIBRj7gLDReGrs2XFveBs2S/L46mrzS/dOior/zkZ1KqWnFUDGH
DzR4VyzrNpDiPfz4AWx92Rjdz7m7MzycXbMPS0S4hy82zJlXVS852MhifwN/foLZ
r7JbiVURcUidS7NlFGWpx7LABsqgq3HW1Y3YXt0NPeyLBP/bTBe55v9xPK8gseOM
pTOotxEAGbmJmg9UzlGTGMsu9c6xRnoowb3BmJtZRnvhnzm0eOmTR+eFslzjAFfG
wGhdbk0Cr9AElP4+w+rY0ZbCnWDTsWo+bCt1GEduB+QYT3mUWouIL4QL2ob/AASR
danMZwhXOrPtdFiDXNbTtrnxQrQ4pJM8jNMms4I2RufuNpnmFlszYJt9miP+qq51
lDMVi92LfyGS/wOtjYBXaGOiegugzT68WYqL/ZC3TrH+9mKaxS0C9A8VHjYktJw+
2LLPBEoJSjMUaf+fdTcAkzlXnvx1BQ/IN8Ete3QnDnbJU2EhjvZLl0uwGBqVJ60h
QmnIQgCTPqJ7UaXOZgSMHipjLrXnV3bDq01RZ/o9L4BrB8qbFE/aRIeY3CCSFigp
pXT8GNCfy8ae5y7tMJTqMReCnQLmQZchOaKUA6tbkocPJdv3pRfVs5Ds1e+O1NgF
2Gqsw4ar8MeaUhtPOHVb/MT7+82gA9EqgqChXwrvZ7ze+ta0rJkIEcsK8Dzep2OL
+eupo8lpVWGpexvOlWq4wvdZmbaI40NG0ecrY1IRRzt0c8Jvfk/vguwdz/cduTS+
EMxf6nbVMpKMi3MS4Hrhl1yNj8PnOZVn7DuxCjxIz24Fj8OzjYL7Y2aGjGsO2tQK
42PfCOH4SsLwoHK8Bwfq9+eFnsR+OQlXs422Ab6HfnSE/2ANyvewloBwe71odMn+
qNORXcACC77aM/+XMIHuZysCg3a+Cdy6vpetq7e9w6v8qhwRt6IttLGCWSj12QH6
7j3qzp2Wln1Mxdcd9H8jf2L5aCu1UCU+VTCnQd+ZV+WGPYqozsEPw2n+2FziAtrd
mvW867N95Ab5XOZ+tAiDx4rEInu9vKXlsTogt75HaHf+80jg8bRSBQLso/gdjcoV
aHfUGhVV2tYlTFPwxk/67oHDNZktVMAfr3PIr03ufNSZCBoeV+6HnofbwPnSVRw9
gWDkWQx2Ih7sRkneWNBD6mHqsfli5cHAFd2gl/dfm8CdGUQZGbI3fFir0jUkW372
BXrqVmiBaIaiuxvv+iwEt5Zy4AZJMVY4FLD2CMliEtrW5cuVAVDVAPkAl4Z+1kfk
Nh7OUrah6yxCtmnmC4O8JP8FIMFX/UyljBPgN5UCcV8xgqGTteHOz/VZ5VFb+6bN
np66zC+M8M5mgTl0qFUjh+UZEqwKFSHC9QrYsWGVmKOoCXhDgRbpyw5cnUV05tSg
b6akVRCUUD4Mlp6dpaCzQ6L/3rWRXWyLz6QNT6EDOc2S5r5A2MKCuLms+PesXnDi
yetwXxFF6+AoRC2zeEGC7Y3+DtKXF/t+abubqyPCFYj5UiqI+Fj/K9iJp/yMSfLJ
aKNzGXBYnGAsN4yRoaG1dP0y6oaCK90v/wHMXq3AaJtnQ6eiHnSdZKmGeF96e6TN
Lzd2lISdVaKpsYR3xLNgsHTm2GmzWsNkjv2Y74a5zioxrnW4HLLo9zsA8hd+QtM6
YrPaUH/K2IeJ/wb5LneB4/o2+Gyf6e2mrBlq8tTL+6JgKnqoOviI0uZ0l/Mlensy
HfuD76OVk9jJ13N4XGWaE8D8aaKhQPj+IsgsnzxqZTr94R1A9PGuzZykVOSt3jhz
N75uAl2FdgAnjdCKvK22ghU4pCJcQhLbDOKYhkSeu1hZeqmyBrGm2CB+ImkpvG0A
qWO8yUWUqyXtC8ZCmbpIYzAMhlLhBIFKWedrnSlrqkJmL24+gQxLNRpZMcNAWpVT
JoZnYP/52sSvQ/KP08cBYNq+A55Qu+W925jzzhnZ9hBwJxaGbmvPIOoE134iTI8Z
K04QTBwIGdndjxNbf+1+LYPXlhNJSbfhyJ4QizILXDZ7xkPARpiYr+BReJcBRx+M
6AB214abtcUpSazL8i5H7JeM0WRZHPTNy1MbNhrhQjkmK1x9ZOXX2lKwCHGeuxYw
BrfC2dXA8aiu5RtEdiUHOgzu0fmXV8YePRY1fF1K0hudvH2d1eV8f8w5rCKCNfSG
9mQoKz/iVwqpXdySBJAtf4h+jZjZqEq9Fo6S1OT8b54uUuCVDYaHixC80tApkUgV
oenp0Z8fBiB9XnGkknEUInf4dUhAlWvmcX1WeIhxjPD5bp0l8mcQjkhEBauIZ/5P
IlkxhFh9WF2kvgODGthKwEgj4mA6SGoEZncwxBEtuN4hPzthGsL9/WakBNRlBFFP
bM6SWPC3VtgI3dIoQDMTqSyCGwiAEA1qKq7CTv90qD/ARZUJe2DIrcWRBuIiUnvF
pzd1Dpww2jDvkyl86/AiLaAYAq2W+WEoZcoqYuCVMro+mUdobp4QPu0jd+MQijRj
GpoQP67ffqEbD6gmyk3PsHcnUk2XWgsg16/IDVUV3sP0tK94gMrGHjXygPORtZM6
QEAkAZMaDEHh3yctOmOiVArCeVhXXOQSLuxMUubXE1toDsoUmxMKXMIrLwWthdwt
wFRoCdc+DRH3CTRdll9e4JzL+RjDROGnqNNnZUCrEVdCm3kT0FkZKzC9XOMr15Ga
NaUZOmyDHB7ri9vjMuooMvPvb4aACO11kogDa8kD0X3O4jTmLnrIpVFZjx7oeqty
fh8mTJ6geoMgUFQ3qJ7JTc3SrCYL15FbbNIoXlLDLAHaAKXW8fJjFn5j9nJ0dAai
eXJFVS/t9CjQpb4MioXQPdncV6IDbtOLJeBUMbO4EcyYWbrm9k718uKthG/BSuSv
Nd2Fnic9EVXoVPaIVhliizCc//xKOJk6Jv7uLVbiIdgZRz+s2RWH3LhgTsGUkmyY
tqjU1vEzPOfRwD1tpSIThFil9zoPjNnslL5E+757JAfG+uNb3lbJCFKGaMCNvvnq
28SZgH/rNOfUM65HY+91kKwwuT3frjEMMS6gyy/6kWKH9MRJFvYoGS2OaTCUOwuF
f9U5gWmP1nuaeufUK+jf2rl46g9tGa09f/6UdZ9DTpMU1Vvdtug4GVD1sHQsSXD/
u5HKB6S1pJlUKe6FsuSu24ES40OLa0prSPJvF5dNQL9KmLOvcI5exvxd01ETjBlG
L0NJjltfZgy2hgyNLzRO/ZGp2SplAJSGIBbD1MpuwyxfHXb+RA9HAgNNaGTKJNd+
PFp1Bie4glTB4z1fbyeMStteQTkWSEQ17yx1YUBwjfxqiO/SjEgqLvtrAwyFg3/M
c6fpsaWnaCHWt0ArutDo2B7DUbpmkgBFaVyMgbDCFNOm1yJRM6BZHN4fbaHJ83YK
c9efzBhKARTQ0vSaBko4QP+vNjwJkJ8KTUBRLl8FdeFBAMZqOZlVxQabqCNv7LwF
dPGj6qsGaq2tf8Q/sP8yh9XwWhkcrchyyFY9Hj9xtLVGVVe9PPpeNYzYGwx8S3uq
FVVENAkoba31zG2nSt2sYqFzMwk4xpFOtWhPfcBoitEfQg2XijKH2hL0R4Ymgecm
j8yFm2rlcQmXp6BFXM7uS8cEd3M/1a0xrxUrzrVCyK9rhGyOpbWeORO7tTqxG3R7
1SgumdIhqVcDg2cACGUK0Rjk7x8n5o+X/cF7EIHUX2hI2JD8VrmNQrRmLHvToXR/
1YKs/N0oiDCv1Q3Mo5J/HPX2ERv5yZGCkw5x3OQcd4hjHN36mrcufpHdWdJEHejM
OH3ZNouFg2D2BrXFUI6tcXT6uu4uEzFFJp5oLhj+STvsJpWtE4lwbsISZUg//elN
Vsvz/Gr0IzeSGGIYX+1pFpIR6+cJKFSlD37CIjJDeCqyhZ5VVckdLtmTnfA5uX9R
vvatbnv/nvetHciI/7Sh+GZcc4izY8jGjPJSHIIwpG7ZrWkEnY1klVWxcollrENC
W8Lm9GKLyOYY/vsjcfGgEX+pB3JM1dk3VozwBObW9P9WeZht7aHstckwFqH5aONm
UsMn9Z/7Z6gQYfYc0ARZJzOgQbi4wdFlV+3vYqS/YNubDb1YurZDvWTPVM5NYxoc
M5uefXD77ZoIars/O/LlUFUD7fBVwoL9xts8GQnul2miZ/lkGebr5hTnxs1DB0dn
j7MT0Lxd3lxVni6d/4FBlkMFky9pDMi0OMryh+qtrnl9phBk6bHzUzmZ385LIxYd
fzRs62bIZC4clz/TX9X1Qq3JtOQMygAwgDBTxChf6m3yxS1PEpt9Sp2wVNAO7PDV
ie9A/jjgTI9d3WARVbUl+Dz984BbPfwpvQhZwEmdzjlD139NX10w5/28UwTyL+UW
sWTgnPmQQYPedc13B1chJUYV+12Yenjwo8qaKNmlxHGQzkMMoipdDw6f0e2eWDF1
WgTxeYUdFy1T7VUFXig9UTpDNsM+Sg0MDxb9Vw0zb89NElph6Vp8Dx/qTWFBiaL/
hjwFooqCr+wOmAyDuV9buvaV+0vUhXEudr6c8IgNNdyT4GixpXVkb0CGpZCoM4Sh
iSgjR7OLWaEQZBKhEjKuFnvVSFyF+k+4b1sBBIwwi4ATetlF3+4nKsYv81vgMzzS
2TTV4ELNwT0c03vQwUMt36c52c58clrNy2miWNIU5eJHhJXu1ziU9mV8V0A1yd0+
njHvKwEDDMxq7SfYMV9RL9Vv9ZB5Ya6Gacq+aVYvNydg3CrW7uDlDh5s3uNjDXQD
Zu+73FHKLEWCmYgbzMEwsJ0vY2tlP0FoZusLQuQNzM0S7LIh3y6JRTSu102iiqjF
n7+DSorgowwrq8t1U4vHRws9XL5PwrVcI86O/9ajTRwNoBkcTeS0RRHp13+14Zvb
j91l95xB/ECtc6BROQgDnZAxIpmnH08nZUyvQRhfdWzQqXjFI4BuT9iymv9TLdBg
U1ID4aN1ze7KLkzl1m8BgO2z//EYQYsTopnrPEmrY2g+xNMG1tP1XyL62knFmhdN
cwLt/q8MIHoRmGn1htqgDdmyIBqFJzGD0GC0szZrYue6hLVp2G4ut40jYJLS/UTO
5bII8Nc6+lm0LsoTFiWERQrK43fe6kviXtCyZpvuy6ZGcM2wN0/TlC3hPGlDGDe/
cCtA2iY20lDzyHmxKZuf2p7hZw2TgoCgWwApAInzt0ce2zpS+d+CZ6XcNzgjT1xa
5t0cMDgVN6b4TaQohhSHu9U6IRIezsYZ4AxRUpQGfHWgR4b/xzj5zgwW7oI+PK9S
VLuUA7C1HYduqoZEGVZFRxL1HOBEBCYxp4QOwJE/NEbUpEsV8DNGqq2p1pEN9kKl
17MexjSGBhTfdCdxy7eAGV8WchWhfnPBKa+bL3p8yXVpSSHWjHbInXujw3iFaTWc
5Na6WbEfop/T17jnNhPxvGEie5XuyThHJCAhv3vPf5iIttywL+6Gn5Hx0cw9wLgD
fGLZybQO+6BI8sNNAaLUQbBh61jehJMEY0o7qcZnVhfCmGG9UJlIvFV9+pgCnv+9
e3mRlKVz3aYeh6gCguUpmq9hLydRXuWseetfrmSuLY4686ML0M03Vf3vDxjbsRIm
sIqwBmG2UoLlrRzGkubcE1z1R/lWJxXLzSBvXmoof9n0Wvp1vPbksS1OL6zRGVGp
7Gif4+9I0yvByDFFMaErKoDJKTJ+lmqkq5yZod/sdTqIk1tizYSGugWl5i5GLCkZ
8G6Nm3OrqCSNBOf6R3ko4zagVYZqVjVdkXnffQF8h81xV0xglmQwNuuh4lQ5R2o5
X4tHcmMACFGfvJszxBi7KUdA3pSwgnxEBnz1GUpk7vD85xejkOLuouOnRiLP/Hms
KqE8x4EzSm5hDMs2/9n/1PYyAe8bbogIBKdjX642vB3i+cjYezdvPgfu+D/Ysm7N
GSrfdoKJKpoyNisfmYsLGUdCDD82PchohT4qxu42I3627N38td8igO1jdB1V/p9D
YwRuaHtcBE8q9fB1QefcIJxxZp6MCSC9VI5ehRqT8LRzrfL3keBVwL/cYyFmruvo
nk6+yyliIX8IFTe7JbthEoDXtuEsBo4RAAM2ztCoM+u2zAflRULqJ4xVrA0Goojj
3FNu0DFu7zl6Q9feLCNEF+SeZVs3vuUAy0W2+P/283LoYZrwJkQ2bASpjDmK9Rk4
9eB439YaLfaJAtDyjL/woS5MuvP0gNwQHvgFIDsHsNZyoKZjFbeuO+i/fYhisA+t
kgi+vqQMEdY4WXEPC1xM4yER8duptJgdqAoaMGu00KFtFMC3x1qgj9eUPPGF1Oqn
OGj6m5nLY+24h2Mi+W2Itzb1Bdg6OJsrxDRwdhU0Utj4EAG8nv+AVcF6NxNFuigl
PpKPPCpprDMOQt4lMM9yUs/KnZmqK70f7vEICJ1xCuZUQtNhH7byHpCCEsETBv8L
LXWGprH67UckI7WoP5rJ/tYCcAUVIec4WuV51dGOgxE2wy2soosQSSXrdNfKFy/W
ybpkNHDsNzRSGsaEE7tYxK0v2Ftbfbijtc94SarGYHK9pihgrkdtTTblZSCKO2ZK
6Y/eQwa6hl7xD2HPVshH33zmPxOMsOOrMnIDTcew6DtulEv4DpdslPckx2kPEGxD
BA+ig+dqc0HFzyIjXTx6DRXr2JpPgKyaM2MSOeZ/3TYJyiMbdcCo0tA5h4SomqID
97ySpSi0/MjEMyKo6C3LDapV3B/65t9drc3AbjzxkrjV9eHn2ZvqNeHqcN0qWymh
giAFaMjM90ijqi5/qWXaCqHKukBLasIQv3jtPovLZHaEG1nQlHf85VovYwx33yc1
GJd3RPl1bXvXBv0U2xCBKbWoq7pWYWE+bUDTEvPbLsQwpEvE3hkAX9lweYxVylmI
oyOos/2swuCAV4WxuXulHLmKLGY1ex7BklNdOV5ECd3enFGx39Xb2FNWn4QgDOiU
2Wy2uUKdvoqVWsMCtiyTGixeKZ/JniCPPiv2vWpv/yDdISr2kfkgbIalqwgXG2F6
YAytewa034N2yEhssUy5ctW3oMyXMx0K3HYjR0FDvITcW64t/bQJImktqbJHChIa
TGOzgk3IDPfstvKdaX2GrUy6DwuR9IKoPaOIuc9O6sgZu/lbmj/SQxrBiQsQx7Nj
ljW9KU4o555PclifeI3ET2RFzTcxyGny3zcNXPLmB7l+bKQpQDN+peLz4BNj3DNi
b1PrONUCyR2BLr1DrzWiIkw05LTbq/iEkPvOrf0dCt5nUtZCYx5lQRHsnxFDNsJW
8ctn5EnmfevKyTLsYDQt4W8SydBZA333KHiVDlueFLNBcg0PfGWHk9CxUx7aMDrx
uye04beeuJqsc0fUFt+kFkZ90QL0GipUFkymhTeGkJuoEAffL/KxDHmq6uKYjwXL
ewu25rNZvy632H1bVasiz1brnifSXF4ryFPIQt75TkaDvBShjAhR3q/ZBPkhOR1z
EjbXgbq0ODtESfqDZijWkWgMEy0Tzu72JaXmLB+7mCv5u3VrUJGXZRo+WgXbJOLK
QOIJZ4Sb3JreRvf+CzTnRT+sd3BZJcS7BrJYZ1VVHLl2OZgJ5AJKblbAsjcFf9Ts
tZnE7/NtGSAMOAJJ01gHANMsH44rHe8XA7PEHFCJVte5pV5jEVWEt3HdOyd8kxxi
1RiFMBlf8sd7la7LEoBojLD6dFWnK4YuvUKvX+0DTbTwjqAJ8ZL2+ZO3BfVZDXcg
0LsNWNVy5d0/NDQNcYa+yiGixEUuqRm6IPnkT/4C5UCSWkT5sICCjYZt4DKz7BkB
tsfOj1hAT21tKHmOlmxoyvX6dmlJhLdH/0ixFqVaM8NAsoDH/kh5LLpxTgN/64Tq
YtJ307eCTitdfdvEwA7ikKH72A8bKWmfh1TynMJVAv/zJnRlUoAW/fS3oiCQ0+63
Lxl9yN0+iuKRKaHS3ZMfxrtVtwk7oRfMtkTn2DbEA/LFP4QjerM2L/aAfnsq/HFt
K3FKK2eNrrBSsQWzirYIWIBAST/A6ssNWro/CypbKLm8bxE2LsrYsK109tByUL1/
DwTZDUcHv6X9T7SfDnWLoyImTBeAy/6eq0KpZ2GMb1MrPwKjB2FiAC++KJz1ypiJ
BAi3nMw6ZSvuvvGcA0qgikS3RDcR0WFkxjEvmWphwczXrJi/4sjOedvloK5ZEg+e
SHK21WZUAIuunZTmsr7G3iiWeMWjz3CAM2Yak4QYlJN/kxQYfCPIz6VPc1Tu0SR0
f+bAG8NJMezGS2MJ9R4gQA2gsGMIhc1QUVUSZK3jFUcBqGQMc0QksFSN8YDXl+38
0i1HQ9ujtsFd/TlN/Ou/1CXWGgckctHjDsyhD1olhG5YQIPB7QA8ml/wKbd9R2gF
vlHvV9H8HvY8nxWKT29EFF2yiKhMIWT1GoPcxZhzyECwV1M9jiegOC4XKvjiK5pF
BJc20PX/vu4+qfiiY1eV/+6JZMfOQ8fNaFbQ13ZpCj/4lYeonep8pMyb4Dxk59fF
4rQQ7ndlFmEYJQceDLijvP2gXApLOiXXiOoeJgoE77CFckD1f6fndTn7rR+ckHPJ
kU3WqIelwlw5BbvcORJT7GbTbIQZSpeAkWhlWWoJWCvb93HRXY90BiVMRmAvAfo9
1V7riw1Ql2IhYNZWY3dTunnkEud0HoRe2slxSMgO6WI8o7mRNi2BON9onf3WRbRw
GPmhGCi6VXYxlo8UozzoORICODtwkdiZsGxV0aRp/sKqFVO0vgoDfxC0xb462nE5
SSTR69FKvMZoTNkKQjKYMPsfAdcxHTSKAvKYtD2vQKxuRHkQsFvZ+z8j/dYA6t6K
Mivsew3xgNgt+RBSIZd+jK2sEnkm7JrVE6BxKpeA6dCwSvAGAUk/LYB8NDSItYyq
V9cZSRC8Zw5k+R0D7PTii6HE9Rhum4eyZPk1mR7v7dYatCByFZBA5Fu/631mQ/x3
8kuJ+8J1eL/UB1MA6EO43rjldwQ8Asj+xkt0T/+7eBPCaU7XlRXyvyY3kSPh7zXQ
8HtwQWc3vkdmcYzZ5QQQqzgupUBgch6e1+ZZxc772jgTmOe+rfIqxKDIzDGQ2IQx
LEh+/XYKXXYJ8pw87wf/IKjBYXEp2ri4jZRnhLGuNplLlCGfxatK11rfqeqxiE0G
nEdseCNv6rwAg9w7RfVnlT9D7NS7gR2B9wEbF39a7pNT0FL8+VJ/o4es2oFHj+sr
1V2WLNlN+MnQsVCZz5XIeDh2i6a9vpdbud9WPkxJ62vW4jAvVmjuM0EpMZQnpztP
ECEEW/ZVv46LXE+gvxQDIzhzowDh63R0Zyt3leMK7bToHcHnT9l4wjyD2MvYKFFx
11SjRvbHCYQQeAm5y3ril47SMeEuONfpsqj/MwaL4gEdcDWRqN42RHVf9atEJrcZ
uFBT/LVjEfsdVzYGwWcV5/qBn5IUDKqm/k1AFTuP9wfbam0yET0QBhdnLvNmmnqC
lqE8Gw7cVc3kwluJNRLTxUuN+M0+/HMTF7vYrUmx45P++GilDUvEB9YLBU1HHLsi
KnwJraQcJZFU/N8rNp4Fm6c73xletKcUGeOcbIWAw6Ad5Xw2n+uZPZObUZCLQrbs
1H+x1jODq22vfJ0jrL1k7PYklV5O6JG3I/ZcDfKITAPsyDndt7qEZKLaxI63ydNM
C5rJpvprfaVPpdcfbmRqIjrldtD8qZjLHYBL//s+ZrT0vUTlcuRMBqBVSvzvKKzP
2OEXwREZYKsmTXL0zR0mrXbtYdPfTszaPWGTB7PTlIJZO7sa2YVku7pHjmw+YTnb
NDpUJtjRP18JJXYa8WCaUZOOEhQoKiCwv4FpGD6BDmCVn/Im4IjiGNYhfOIY9V0e
Lv9ImAdOAHmKul8b9isgBfvl9eFZPBQortuOsBsRpLiHCYInjgBQqyaD2ZAj8tcc
v1cVO4xhDiJJXJ660EuZrntoXdGQsG155mWa4UoDrF2mOFf+i79d4gY4193+zx8q
y9o2NJximXO4U91hwLtbUItOInWoea/0bFoza/KAS9Y4pGLSqQ6/3pyadxZK9bIP
7QepeeSaKUGAh1/jYZCDTcdWdaQ0VZkX69vojVRkP+JYWj24gA3IXrGzsamlRpQH
k0k1OB7txPeFBXxzyWRT9UjdNrNaMPZO8CtCu6hdgBqy1wPWLaCJ2FOfJf3hQsP9
YRx0oBT3FyTzkOygddyzNGffzmf6INE3lnOKr45/Ava0yX/E8NJKuWmqS018f3QB
cm5cZBX3rciFbvFouuJSeFgA2pqL0hbB1k+4XEGcF5pUD+wRFuU4yqICFbEosXfK
u3PX7nBEdqFxNdVzCfgD9RwCeVKqLGQkWxyaPZtSspznqkaA/vx8bFcsAkFPNagz
sovFTGDFlFx59B3rCrdQIS7cuXDaU+lSEGSL/OofT9MxfLsOG0SDQsKQa/I/NIUc
63S71e3lzZyaiPtYIRtiwKcoAA3AVdSTUtH6mXsT0Vam/MwGj14cRNoidvRzul3D
rX5uExjQvXBe8uhkhw1NL3j5PQ61R5EFQbhHpocYdnU/7avkiKUpH9WLsROU2CMk
GV7NRfPGmFijgM0cb5jgxaLc7RR3yhPbN5I4WkRoeWJOuNeMUatuIleVmXEcB5cX
jxq83GUgYuGQWU0vAQ3rmFkxKl/Xzf5Zwn89iApMbdTaD8h7YwqKpiF3QkFW0N80
ssWwBYd/Dihi3xjWSsuCtNQ4eCTidxUV/DrxGl59CHUn8W+8DCHwBQrVgO0zTlHI
UeIwPpb/plPEZDNPTyTk6de4k1KX93FBBZ56Z1MPOmcn0NZDZdxAAhjob9GU0CMM
26SMPuexccsluM+shOgBYffIuwVPzTmPygqfAhmxUntmqF8FTkJefD2gaheapGr5
AfMjnHIK8vN69c/bnKftebPSLqZ0vYAlHDpc3lMx3mto8Q6mZHQN3sTMApxrIBzY
LLC9FCZudh7XFva30rs8QmJ0Dh6qrk9fXl7p3WJ6LdEFXu90ngcnNqHOkN+EgInh
3juSZHY8XbejrKy9jheBwLpGofsdXadsME6txnGITtzm6re64ofSDz6e3Syl4vth
DwNkICgTh/5JgViWFSjOaD8Snr78bDVCjyCmDjYZ4xUSx5XOaH3Tj1UWMgMosMxW
Bp2gOZiF1iegme7H2rffmlsSzX5xvmzdusIoKj+PV2pHGYxGL/rnrzc9gzx8KTOO
o6zVQBNjl+UfFdNF4h9puxJPBmhM5CwgxuMghU7TdFpg42cAFXBDW685HvDfpES4
Zi9kYEBruhwCXaXi4SXjzh30dr9W91kysle/ZkN9jJz93vqFoIq8WXVGltboJib5
hfVCI9ZVzODVKtyopb8dhR54phccR3n7mKNUl1thb2zt2WE6/buaGBRqkAaK9wwU
WLoujMHZhvP2iGlBkZg8BoaiLHRp4yrNfjEoo1IR43kMN+KrGSMNXB6agA7cw8/6
v+fX+xCCUPQPWilmEy80jOXQH1eeBr+Ci4kWdEbNlgmraMWQmZnsx9FeFU/hnviW
+SVisJ1w1+YXc7TN7bJbyLRNxWmQ8Jq1xp4Nv2YF/DM4TGZ87vROBOjjalJteTWu
JAEQuapujL3mkYpq/WqtDeBusM6woXbq7ibFfq8+xkL1XWONlRonr2ykBkol/vAS
RfmS3p5BSNv138N52fPHvT+i1pHGNKQOttZoqe0tsdCxpZlmED8KiDd4lvrDiZ+T
+iElATWtzAlbDqVJw+AKftXHHjIuo0IbVoiK5UajWz7tzVf/x5rRe1XZ4F5vWcbh
8OqG3jDQutgIWQlxRobmRs+3ryx4X5zR/6DnFxWeKXD2dDhJmQrBHsECA9ODUP2r
imHkqB3KntioVXedFKSZvtOzlWp8MLLKTWLWp6B3suOwAMILcJ71zdMpJERccW/7
U6eUK4rtZMy71+Zldh38UiywyoI9uxlb89mVSUIirDFuOiYYsrEKykLzLYe+m5bi
EzEVIeNaBMTPDJRMrbLz1MTXjtQzByxwmslt4bJYDriCHj3yuWmmsks8Hhb8jruX
J/vHSGhjVIfr+bj9CLiqPDJQ9uAwt4qOk3L+jSphInDWTir3SoZACrIkJkQ4RoOs
HfbpaoVOm+k0AYAdg3kvZ1CCkTlXvvLns8CY+++RYllVl7pKtKjSeZJg8dn+yqmj
vohUeQV8oJ9QiKCXsLUZDa99OGoyHRmGpiUtveMyB2nz697uKpN0FY+PYtMvbpz0
DsU2bFUhimcHCyCX8Xb2hwv8HJb2jgD3dVb1g+HORZ6+dvcl5NtnQ/TLuUR3GADS
8zHqAIE4db7csjEfbg3anlF/HenOQ5SQvwjnFBuKKLfXIC1BG8uuAv9dHUNbduxS
wLcUvN6zJdU7Yi0y7GS22IfxUY9c0qQ5hJe/09ZIKxaoivbnqjIT1jgGkTYGhvf3
OeGMKngTmz/X8B256/skdUmEd+g1Ba2c03Cd8kDK/huCJghg81CNDx/9wv8te3RB
LJOjw5WWtCVlRMLgsd+nOsyNxHlMKqkVccgVNo9pzGMU8YGrXzguTEaaVVkViliV
xGzAEWEZ+ZkO/mRtsCWWOL3SnMsur/Zol4nXaKLYos/Bamms7a1tIsRQdRv532bb
ddrIttgKl3/wu6EfuRo+lYxka8SAkP7pO1r0jSuOssZ4UkejbmFn8G5lJqWY+UfW
xHIWKAjepVocnEazJTWusXlaWe1WOVQ3WL1FGLbrv4kXwnFd4kR6vmFAjsHq+wcj
i1jTVfUEoryu1nEtHrNYpzKTnM6ut8OyEt5EWXzL/FRYlm8nJyQYG5yGnf41/9mW
eELF2Dzv2qJ6uz1IYjJS7VwIb9F//KKut3Zn6hr4ULn5tOFWtEles9xsaScfLvig
NkX7Y/y+7t79Sk9UVePbQ/1TmRGQjPrqSMKuDfF2zd8wobnJsVvdcVXkbvgI2KKK
zb/fyx7uNnJQOF6QwZUH9rIXFZRxuRuiEUs1ZdLSjmL++VbIYjCJ84t5u8FkGLrs
di236SJHImI7SRSJaSJx02eyNW62vApm7LXr5ycArujW/6rf6QFjl43ZQ8NDlwqP
Kcw6w7ra0+ZE14lzdx8LHdJmp8ftrsSz5HkLYow6OJXJmFWzLfTvRbcDCJwUCpMa
UIEI8b58E/ibat90ifBWP4cn/Hf5v2NmGi1wZmOE+P1V+c5VijDTz48GEh1bIel8
W/g+TqdC3PSh+rKNh4JFm6OgscsqnV1phwK4sPdyVXVDkY6uF+1ZhU8YcjwZYH0R
rtNOh9gGUJS7qIy7+SQ7K5BQ8YKnl3qgb1WkHs1omk0OX8pQ2gbx3M4+HWwUjdYO
j5bGBFLdj46/wtRDrDu6FoKsJLUvp9haJAf6O2IkNT3yj8X6vD07t/kbr3GI3h1q
eYOoLdgcA/ikBVGw7eYZDiY90gpVt/DXEck0nqCSgg0gd4D05BCQlf33HNlwwC11
qzY8QyMhITQRr3Zzbc3D9ywiJxmhgQ2ncFaAPbLivFK1LEdgeuXowbzaVv1iOniw
wki2vzQnimja8LPne/3guyP1yOZ3UcZakJHd9ulLERM8EMLbFdTFzZXYDHh0XiP3
5v1GnySYkO/PFIBV3rvf7nzfV1abdOyf+URe8ChtGkRLAZDG+fR+qD7wka/XLwPM
/inWWMOQtwn2L+3fskWPkL51pskoxFxVQxfHjRDnunDIdfXeXXux6jfn5iyxB08m
aJ7dbmGM4tcf3Jasz1/LZEA7bkuAeE1gKT5vs50S9dc9Apk0Pt+Vc+l3sMM1As0R
hguXP9FAHM3T6K2dob6+WeOrZvitBrB2h6GnirSwbopBa9MvSaCqNu3xCZsreTRy
nHBk+xqQFbqQXD9A9EssXVD1ZO++YdWGPtNPjHDl8049+jbESbgxRSqny14+DJtp
IYxDN5zmTzqoWxF7aqJWv1zIL0iWexV87nH0GFQBP0/rgV5/klybtbFMmrkxSJDo
/mw0ehp0Ct6v0fEwp82DlRdSV/sfkYIlsEeYp61mdsrRBWGnCqC6xwp9hCcQ6T+B
DMJ4Njs1cRe35asIT20jzdX8+Zxf7nU2m17gw2nawMohhFQhbEDWKYLgSkXwo+pg
cmELvwPyJsZ5TgXy+5htBjgK5cK/5eBADHFQMMUmi1TFENX6fdiaMAjOpWCAB8H9
Zt6ipTQKwCLJuhzAFYspyzUrn6VdA+8S4RHEC4XaID+ALv9hBdCPC/zUb4ZTndUN
VNhCbti9eg+szs3MNVbO1Wm/BTjSra66QU28tdl4zLzDU1RkC6wAYqAaH+GWaOJ/
J3FeryC4dU8umQKLKAGmF6QWy+GfTVksBqgGIkbdM20IxIxmh1rBDiV5fgaV6O7Y
ZYNWpxJwy8BQbjrpbfubAJNJ1DNh7uy7HXJSaPMDCi3v5gVsOgmixLevfPIhWn1E
EdxSEBHPeZkgEC3zvmThu4YjspyPDc/jx8WhsSxTjn9zHAK/IEO4SlVouYous8E2
Sl49PrIaKlKX7PZind1Nkfm/L22Jpk83GL97H82kHXrLv8c3ivzMa17qzMWSG8qU
6mc7HsumHk9BJkbOSrAeJHcGUtpMjM8zNIKPwF1a4Ie3LyRFMntCqEEEBK+tuQvk
xzy1WRuiGgNWRDGRwDhauCCSweP//BjhromCKbdTYLCgTmg8VnpwIxO/TCMaWm3X
INAkTVcGwu2e6fgsW3AoOBUClsv8S63hYReqGmRGZhBhQOhAixToXA+on9P+wGi7
nfileQyr+Z5nx2jVMkIpDAaCwH4tLHTo9kH2YZI0MQsBFjhsIMjqPq7BFFqPH8Ny
nF6RgoYAO29npCcRSoz5pOzEpNu6LJ3Ln2S9FHiFrDQYFNFALvqWYGcjfKN9bwdt
tv+CRBah8otoLzYbzUtx4lYYJ19eFLqsLXXkBWLqlC1JBNCg7f5RYSWsrMQAON6a
0E2jNg2i8/NUaulL39aYaCALQT4KRNIGMQ2njfvZqAHaWn7m78Yb9k+FG1BaQ30j
14ghpaIN19VYyiU9oLLDgN+ziTcwdE+al5MtrflVui7e1o9d6QsL5Y08hLwh5QXK
VzqwqGST2qbdTCP0NTNZWsiaK83wg5o2y/jseh1R40gNkq7ICYtMwJtrF2+DIPov
NLUVMav1Sf71d8jyR6tBseaJEsiA/04o0kQwG+CYjlMNlEy0A/8zUbafXgUgTx91
GmapzkhX7HN08gbfbQ8H37IHIp7eWzg2N1NznimcwsMici1LHsP9HmRMZZwfnDDi
PB23VBJ90uhbG/Gh2dxW6U1t8OjKQbjawIXN3AvvzdFqwjE9/asWomRFr5/byroq
CD4o2Bc+Nzm3gvRbIH6I/ggg77GWBifmsIyOemxY55vK3k6nb36/UcwxR9XhsZgv
5Zfcgz7VuZ02UVTpcPCILt1YBb+3gKZM1Fi48QaZcqQUaknY20Yv0nxWeWaHENfi
2hsq0pu4flgT/r7sDx52V1iEDuvYiCdGaC14R7qDDGhM/DSUZJJ+fPYmiCkD5wwR
yesehY73LuwGSRSSELm8+tolQuGRrkwyfwBUFFhHISADg9/+od/JMDIgulnNRSMr
RKFbDUdqdjLrANcXJK1U0zZtMnqpgrSktu6z6A8cF/dLlP/rkQVG1AvXj+yyNQQ1
nL8uJNCntS6G7k8l+HvmG8Ab141dzjLreu6LcfHtos+dh+eQOcJjMsN65D+rilVK
AFCR7K6cypnzJOLwxdgRZ/nigBxLXRJCW+LWFoBKVPjlRxpD3q56p7fPsLe1bqx1
tKj1K+xVvWlgRNl05oGW0KjJJADraSkOZkUeWkr7aHUoBmiwBbFCLqF165xRN2Fl
hEqylPAYcIOvYsCzijkiMnCbhegbBtP5UIkLHyNYQ8/E9w4Tybl088ciRHnb1XVH
UXTqjbmz6Ne0SUTC9k0ylpDHaildyAhsfQOcYLLHOKDfhVtGQXqSUX0hjvrXHzwO
flZYSEBCZQGtdOEdagYe3hgaFXDHX/Y+MWZwcbT+RVry2gW1lbrqirz2t/aXGSVd
jk6eIviEk2cQP1Y5KW0tJ562f0XZTjwycocl9PdUWzPm4KXaQtxonoVAywRgVAvt
FOJ2YEWPqE+fEgNURokhWg3moVwUvOsgDvYeSNaeUYgHyzp+eXtJQhYwlJAvc4Ql
ds8wmm50KVlf2Id4wGZGvzvlBfHd0xtfCZgL1QolfD2gCFOGlHOSvQ0HBFbp96GI
h2KAJ++drM4n0JA0kExhtlYjdoFTLE51wakj2iqoX62V/iayPisOnPFtcrTga0tt
IGwd08JC+YX08TwOWc7f10SMzIioDlYOarCj8+BtRqHfV1h+e0NmYBaxKd84DFo9
89/n7PZo1r+gp1DJXs/aPPIiqXNa34eubXd8R/LXDYfGPKDrZHc+1V7T6YzGvYho
1f31JY+WPlZtw1gS03M5lL6EsjfGD0IFJjRpjjyM/5ydVQXLscvuUiAM6mnV+aUN
xAKxasLtemLlCmucMLCpK/INeStoKWJhXkBWkk1/PUhdRraAkFL8/02dLzA6DccA
KW7LmfH+YEVvYZhVS+yB1+FXfMDT0nYEERvYcKnwkQH7xcgSdpxWB3ENz/AKGiOG
FwbBinTo8pxoaBRiYRI2WZG3N96IvPIeoa3XRjWO3y/QE6mexp9kbk3WnF7r94fi
3NlFj36HR0rD5HcON7NSXzlk5cU+yLrxYkx/dGbb0lHkLu/ZvS+4O26crF4NuXwk
fkzj9dbCs/CoIsqKMoSaN/rKUizZ7l4ONxZgt766dGZjOnYnSnxB5iVY/cAdt3gr
ZCi/l2L5LiMO2ZIMcT9rQ3eZlSt9flYxa1BjKdhZHKMOzbG55iyPDbCR2KFq7fOy
ASPb9k8QTWkjqSW9HTD4YqtY46rW2yHF32z8uzWRmrVS8a8YKI1kz2N1zUowyWbe
g5bO04CSrTWNA3hBiajLFCRrJDe/qfNmokpWomwi4DIW4RNueADMjCrK4VfK+4ek
93YkxLBmaOo0X74dDleGK2R21+hp3tWXWWXa29XiNIOrvQhbsE3OZfj5Z6fLvmDb
C6T6vPe9APAfGXgG++DpbS2ZwJs4vos3utTccABH88ayaqTFkXeBzCsTFe9djL/M
vW6hrz/g09TTBfCyb8yP2C9xJjX84fHwjivlXv3dXmLFdvl9B+o+Rh12qS8oqkzL
RBB+syUwXFcTXmuNA6BGw/RZg2ktdB6ZIfBh/J7gSWm/1ZAYpKBQwZDsNyoVLp2g
0BhySJF9pfKT5Mz1TtdC+souE2jAJizyu99qDoNVbhVydusDzU/jYcEgxZwA3w9s
L9UYDGvmy99ticoiCsEC8Xkln3EgOO5y7xH5EulxPWDuaeiyMHN8vy1F380ibDGl
T/rUKO8j6vgzRzt7HASA2B+Hy8q3CcITSDPTRhT315srwf/nxtS5urkGfJ28cyQJ
LoAQfIOIARvu4m7N4PolKXdlfqssbHStNwAkup21wFIhOAJupA/L+d5Hr3NQI+kU
Chi1h87bWu6OraZufzTr04a7mMfGmNF7786k49/IdPgNgntUQ021gVUsa7IqEgNJ
OWbAo8ZKTpWIF8GzPTdB5si1/nxCOWbaWuEX2snPKhRs94tPcBwRexXBPtiYlOP/
a65iapLNAu8TTEvIg6jX5K8vn3dyrzbq9sKmzlvhl6Sf9KVwDah67yI4437YDxM/
qX8dNmoRsjkpw6mRAF7yrY5GPZWLCGYqcH63a6R2J5rBEB5SzlJPUgEtXjA7Nd7a
guCFLTx3rlfYfG7w9snd3MUngl5wkcscRvJOTrgLLDBKoaX9IMW7ULw+KMR/NKW9
sBa/P4lFw4ao8HurgQP86NfzbPARvTN7q0+1BzPChM+mEmR6IVegh5HIRhTq70ON
zfWCPcbPOi9XzZqsLo31gQ9eEnDbcj/0DzG4KMgTvbxXFVmxe7AP8fjVOPbWeuO/
ZJLh2PFNwxqX3jpE0FH3ZKheEEl/mfmLLSgvLreks6ekGI5BcDs1PYTV1WdpNjCz
/wxqErLVF855C8krXSr7JBeDQF39c4KiU3l5AlNO5gDr1KVCgyCJVy3H5UcXYVpE
VOc/yBRbgtRcSJJsEGsz621iIGiHLcPltd00Sv+pAx1s1kQd9vB5Ny1xht6ooFZ6
tbmhOfKutkUKqBBkBCPS3rXiXFDr10mLJvQ8tnWTK/zcDuvjv+dElK+U3Y0IHpUf
7RZDkQjccmlAIZ2jDcyOYMPoYZPYZ6tLdsRaE4LxkGiK2x5tOYmZaQz//tFjGFoA
an11F01HRz5znN0VBe2lBWIuuwC49V6NzDxffx2iPUByYCGlUmccRyf1eXDMmtEi
UKsEZzo2WL14A1gYcqG0USdUu3yJusbYvvpYneEzDPKR12HtBIONGf3ZD3X0W8k1
By5aH2aVM356dkv8NpLgMbP7A6Zj5OyozUeJmuog/8FKQsBh4r1JMK8yIsrP9t9g
/2GCSfgX6gSukMYJRTEa3s8HnymEYKqrEzutwI98xWZQ7COvJAdd/486pOAk/5Q2
JW/p5Q9GqXacxXrgC4j9uMtL13ZJJ8lCeBFa4uKB/hwpGbz6KvzxbRe7TuYwsKKy
+O0E2OR4jjlVfLgcm+AsUWowmGzIv1aP4R2WL3uSc2ofDHqJYmC0gr5pW34YkVQi
hdv8QLbxy5Wy2ho7C+iw4Zbdzedk9aM+1ggIISheUqxf5w2La6wN38V43g3nUVUA
AitsKTkJCUEbZEMSL0u4udbI+B48/c4fcGzMJadviHPzPU1JRnf5yzaIjflztIOB
fzcdiDqYsOaZ4p+jtGkJuidWzhOKd9EjiM2aTNDJpjuQXMl2RNuhpdJTqpInBSsg
c7h1VR++OYNLBNDi0ApRnkk4ZRDxEHKIyHZCldxPOKna2tx6Vd1UQJ65BdWc8Da6
BzrPcWR27X/CtaJDwwWG6pQKKwgXsuhLbD5PCnrJ3EWIU6yuO39Utbjz3RD/JFsf
YXRzQ1LDiQm8fv/MiL8Z54whI7u9NctINihGjYOT/2/q8K3g1OOIEEMxV4dc3d/N
IYujeKelOQo1XwRUMTpcKPzULNPQquW/MEuiaqIalLH7D7vsmk35eKzgj4v5UFAz
2mDNOFi6gzBy54B6FCvND6fA7HwMwzVJwZOCcXJ47hRZNbY2oRiWoISY8NVWiFqw
qFh+pnzkNmTpfDei6GR2Gmy7Lix0LtsoOBhx4Nl4r6gQuksI5Za+BLZoXTPm3FW8
j8LdLL+T+GibbWt6Zra3hQpiRyvrp0r9uWUA18fum70JCBCof6w4w9rWONKmGAM/
nta447C6eoUaxs0zN4YdunbpvqTr7tYgUXd8tsEF60mybGtM3Tu8/Tz3KsXZMhFp
UJi3o32Mi5uCYSAELrfFLbem3j2WhMMh8JdTmWM8yt/9g6L1Pvd+Z8tSzqRpMsQH
2IKpIVhaeQhHX9mgJ4gp1w+4vKu+WPscR6k9ugEy+HrEhxnlPzZP67tn7oy7jHAF
G3X0N3isMLxviEiHQoPXG+f0AI4z/XDkQ+cX++R4bUygE1r7mpFnhf1TckezGs8m
IBtBq6eYKTuU4zsr6sUH1C3ZTYKSU0CO+sF0U+K8KgJIq/j5PdDvIlZiq8fVVlkC
NNeXzkhZvGVZzGGzqNeh8KxJd1w1sLnZvg851cFm9J4lT0JVQ/RMcBxAuNVjg8Vz
YoN8K4hPpQfChB8KlNLtP9bj+/ZcNfA6mTFccH48Ilh4nP4InTfpLcwbbs/k2EMr
iSDWHqRVtnM3+lh3PqjQZgOhDAyLu07mHLXrDTloykmexWlK/Zj5DSnNr8R4opcB
eApOGnU58TRmn8yA9hMElVtpZFjvNRm7Mc3L66CmzYwGGaaJVY5jEl5LJUbzzRBe
Jz8ep/tMjhshza4o6qNmeaQSuidb3ZgnRwDtbKMOQabUsJEJTt8Ln+MZv5qHP9Ch
ajmu8fJZveJd2wvbx7Pj46zAcxnnf86np2vQYJtCHFTbOAiLP0c1RldTL6fV+apK
R8yuplrK8Yd6kQ0erLVu2saqu5Yv5hAiWjhBGXeAGw61fBLOrDZ2oho6iHR10kHD
2YZhhoTBKhXpO0pEIHlABC6l5lCnVj80yjQ2bnyGN1Sp8lNsqtN5tWXc5zTqrz7C
Vo/shjya9XcK05w9Xz/UzPNVdB15UbRURot9gScXZu8XunFOjDYkAdW29MKQWa9i
wHSyZAbpcEifqaC6y+oVUrna5z6iRS33HJ/RPGn2G2sC4VTZa91AqJGHZSBFSnDN
GZlAGKmrn9/oEee+RQ/PIvMNr+aymA0oLxzVNDQypSUVxqIF3zm4KGlydiPo89FI
BVf0RhuXUtPpOstVH2Ng97NW825O7KTY1jwXadiV6kUKmXUr2q3Mig7mmKLATzQi
ZdLhEwP733XeT3/txloxevYP6FNdj7pCE+Vef61z+2Eof4w4Mf0RaI6pzBEveB/a
TDSgpXH7Cpaov7xJlNDSwteQhH1xNjlvbwSDNahlVIaycbt1ikggDGe/mjNTzGOC
PE3YLyV2k/3zwDQ7vtAj3GLArAnJ3vn9Wk0eZx3DG6VM/6ThpIlZiBpRJKWudliV
snGi5jeyEKlZO4Is+dvBWSyOENebDyN6BBRuA8+8GUOe3eXdZH/mfSDdO2pkENo2
VU7O15UF3b8TRduW30kI3Iy+MKJTCo658+/4YtMwodcUzDMxN7z4L6VI5w0CBiNk
Uc+6EkzwPKJe4rcvR38pwibjeZv+DO7MxX+/Pwtlvr11cI9HPLdmeTgQkACF7eJb
b+8h2f6N4wL4B5F884Vv1ZxBcSGgGUvEY7Q8ydlk+1QIm3m0FGKN39uyL/qUq1uy
4shdU+q7d4yWv6jmPy2zszlQ+eTnPB3S3ajF/4gV3kmIMcYl6hJGjNvsmu8F+snQ
X0qGb+vSRzYgIfTSUSfJWmFFT9P0Vk8LMheQHBeowdKT27ZYJr/NYKSRvEybyXjX
w40jNqeecAP89+nprcVJJoLYHK8/HHRjjejtboz+tuYU0IOYpf7kufxbu6fZgU75
o2UJvb4firxiXF4x40R/Y7tCCCzNBSQ+Aw8IlfN9OXENmnoo5Hs5WjN/SywgqJCP
P4Gwae52Q2sQlgz994xPGw2ywp3T0sHuz3rdQgValRwOnXm0kEqxh1Rc6+/o+X5j
N/yoZan6rGvFo7f3/QTTBytuPCaEaldW3bhkjqcCY36cKLYXxbsSFoaCQVzs7hFj
oEzMGj91BoXnduFVbBeMHYOQjOxRvvdl6OO14ZzMurAnp9tdbKTYImzjJYnvtUYC
MeouokdD2PeZADeBTgV2gDGPUKcuJwyh6VzRnNEmigk/+6oGRF3MBsDljyBT4om5
3Jk9Lc40XG17EV3l/KidUKhp9v11xfRoseUdwRMLXvLe6CMfib/ya/uwiCgFwLB1
9IkqAP0NtqAGlC+LMi9pA7eUnnNg0pRKokPbCaPd/k0Ukn11V3KZ8uXMDDmJ9NAU
uobjtmIfTF7LZc2JEv/KlywH+fh+Uzqf/sWuO67pwKh29qJ11tqV/lqZL8AZg1wd
WLw5vGJ6rCb7NSAZ/4m4KeaH8v17bgsUA+gROMo3ff9rKjUZHnHsZyoikyNuQvhn
umAfBc4uPfVwBLwPefjIPrdPlvjkSegG/p15Q1ExNhHVFQO6Ua/neua42Pi9XHkI
CEdOeky937OjjmS2gi20Up9PdAwVIwCdnBv30kanXwc3R7EEqnqw7YYTPxTBnzQz
SjoljJ8ziSqjIhIiY7NtyOOvOFXzEozypbDMTYCZlImE1ksilQrSZyMMe1RFfgo9
9hqnWTprtIXG1ptee4wqGgPjRyS4oQ6RDA2gb6R7naO7HEEzBeBuOddop9+TUIF9
Wfp60adoi3Rkm4GlZsxWbGR7/AGI2P8Ng53ydg70yJzXfoDuAciftFPt30O19bLM
rRWN8mEG/AkHCyZtoTMnIxcQ2NaNMq070UAZmoafjzEeGGzf7wOay1FbOiTp1kN8
Ck3iAHvSoTF4hhNjfzglxeAUc1WZBQiJEc0tabrdm1gyZ5SylGIbBCxZZ+BAX+Ub
6GVg0t4TQ7wAI6ayNaPevkqlFJipOPiwB4gaoyII8LcNkfjCfgzKc/Ar3fxkv8h6
MRoNtwO8k7xdiLpkf53VrOyl0VGKYYUqw2o1Zf/07e5U8AlOIQ2qFlrcnamLjvHv
NeYxsj5TRZOsyrecyIz7QiHl39Hp8BY8FTExYRPh6BZH/uYLkiuKZYib4qj9l+bS
OYkAkmSnYIpbVtrX6ugsSLN2b/SfnlYN2HLjtS0Fyq4Ca3254LubBqR+u3huciRf
6tyvoYf9d6IxjpwKUPIPHKnPM766gCbjPrDeMiuZ79ymkOYOkDJ53x7bKgt+iMiK
bVeTHips+m/7HTEFo9lVGsmPgkqsH5pZ33tXhMx4For0s2nhv504WOSzCKVTVZ2n
l7PApajmjMRdogWB9AH15NuBTR4x04ZhFsNlV4f7ngaSoIhOEr6Pt3Wwv1C4nUvh
yJuUk2t6fwotUlyiHPxpxM0c7P/TwK6/fZ006LJBwivnCTqjPywRtjTw9kNFsyPX
p/XwoEKGs2aUmqtsewHhgtJEwW+8q+ZK/2r5Xf2nsFMXUoK+U0PbmiWFc5go2zGa
UPJpfb0Cvccl5tPTDaHaf+niKV32+M9qbknx9P7/B7yG8CuKEIflFs6D1UMc4EEj
G2NL7gN92/az4/jLMSScJmdud4o5lBbtRQrabqMJLIUmgQkzF99XtmDqBl1yIPiS
tTBsoinEDZMwISBIYQrMS2a2pELGxK9ItCPxCRxdFZfhdAUwOD4CL96ZC5GiSmD9
gtvlPx+0iJWztPeKgQCmRsj1dYoD0NndSxCHYtgOBgX36R25UUyhC12VkNHDufOh
D5NH0cpyxwLJaFgNQ8YGFKMz6J86EFSLLJ/rXGAR1UxlYwOiqTxjEROt+7NXrWDs
kkyty4AiSru7Z9nwEqRvzB3VMJFJgqe+pvOyZppb7vmU3O170oTTr10rOHGWw0LH
rFtQcX9LUXAbnDsuZHh0/rppsDetnYxG27rFxdhkgNAQhW++djvQ4L9nj0mCIn1u
Gz+wHGwOemny4Ehz6wXOI8srRH9ELB7f6uF/FmYpfBuzwcZVbttrlLiqk2HymIvx
ecNGpudxA1cakbTjmMhNzC2Pv5SXMjc5QLZQTw3KhA4CJUdcSiV6C53felaEp+fS
oYt/N4XbqwfEiYXjjh8vF1gOPGRWjh1ahepRYNniuWGGiKu0K9/RfAZd2WU8JqZr
JjKVlwOrKdqvpBOjU2NjczJsPbKkCAFoFodgPUvF7QanytEQfwL5hGLnO89SS4Jc
aG84d8C/DrTaizKLZM/tAPVVgzEzKKyst4w3bp2GzBu3O0FzW2gdRSsdCuFBN/WW
+JoGIGeMy9NNcuJb8Q0/JLcivvDfQEh3dSzitr771ehqU3rxF2PuSYcolKWlZNPO
tZZ6Iex97S9MQDjt/k+mBOwfW5EIUWPWo+sLcoHLtA6Ic2pDMqSO0Q+2ewXoNOb/
I+JLS+zWkBOeQ+idaRVK5iX3uL3swTZ+mb8Pem1xPxTxWtrgJeDhtPCLVpip4ZU4
X0Hn6ItwOxx2TQWVEJQlFfW7pXQxr1vD64cCfFGnNCe3aR1nFFOd7SVvHvHvbeVT
BHH0CyOfjdZTf8MkxUYZO+ZVGETi3dPYQBniF1UC91LecjFiO2+SLvAnAxuXTf3m
KGTYYjmGLfYJNqVWpw15JvhZvKCBEQWOpleru59qfSehRnF5Mj0QQRbuCyasMVDl
gPizT6T6XOq5DKOJVaSafaube+AsZWlGqY3jKzGgWcMtsHy2QDnA228c31uzBFHk
2NvyycrKUNlUJ6IS4/v7lY+dCZJrDb/2iVhyO8JDd8To1fsyCwhgLeJ3wUpafLV+
KgTcFjWx1kE8ZNIPmcrTbqSFV06zpRD1xl1XmmdSxQe7D8xXKLA/f108rE0cuKGL
dn9tVDq6IaO+NDKQnVGVihuSHmwq2qFzV78Vc1ZQ9CaO6oIZK6DerTgEH+VZJ+Dt
4zWle2mjEmsP+66h+YR7tY3hOLSdyMZSkX0qRoL/2yLkxbvpuTDwSU1P0IT3LFFm
bLHzb8yEYQC0Vvr6zafdcZ57+AexbNEztxec9ifHkeARY4LboBJnB/ANSqIvHBO3
7mTS6/FGsZxt7Rnu19cx/McfOL6KtTC8hrK844D34h0sxLNPtrVQXOufIkKKPJKT
Ql8axxYvHoDaBlrr745stevHTIMVU1XESl2cDZMqPBcp5q2uKM3VZ2j+6/0tr7vd
j+mms6gvUQstteTsGJa8KlV0GwSBVoTLbqshOx29ybQmxS7PICFIIq+vBYx0zqTH
T93AL8MNTj6T4KtTwTFjB1tnv6dnoXD4yFA8cbjYthD1MK3+HMdgL30k3vreWxUb
Q0OdAcIz0pOYu/nxTBPSvCgXHBwD61yOfwgQMjPhKe5by3DGmwJ8HQFnzDybdgX2
RfdL5O2Ts2aTfeued6xG1Nsfn5d9BIjZlyhhOVdY2McnSy/vTotdNilf0BFuLeFD
UTu41AxDbkhzp+Sskm4ZSzGSbJvQWbdmt546Q7C2pxBzG3J+VcipmMBmlMc9iAtj
oz8ZO5LSjSLwjPWo4pJiySHlPvmUSPWBvhmhVWCf3TSXp+gdAUN21I/QV3Fg1QmR
40EE1IuAH+N8K5LO/7lZPf/B3VT88BvA2jZqwh9GJf7C/WcZvZ9cfghTznBJ1cyX
Jnf6C0pu6fKTPoNDo9zyHa6r+8DdAdbOkKFLbk3hqxQuZ4+zGMCLiap7GH7OaMk8
15oj8YqMl4aYzAMU3N9OahK1OmIe77hxW7eGVzq7PU1SFGNjp3oafNjsF5qHj8WC
59bU7HkPll6Gr31h1M5E7ht+76wSf+VC+iQCADEmiLzK9Nms86HgtdDzp/+Kj7NJ
rofMg+QccZTWkU6E5wKiasXrz6OcskclZeUhiFWUn6+RqsBAA80N3ApXRJiD3KiS
XvN/gMJzOFnaqC0zlIwPJxrBjznE1Lvb5NNA2R/EhOH3qfvXbrWxDx+peCPbyZs0
85zOCcEz2DHxvgRnXY5j8/xvHkr8n8wvI2uMLDC1/jN2ZbILNPSg3WeYjDHsQyu/
4kaGF+SSKJmB+UHlhs1FWdSYWgZAiNJRaDjAQzRYA0++bkFp9OK48INvgU7UGMy7
L/Lh6HlQWzmqfFhNDnELQSZb7oSNiu1ACPJNmYZV3a1oCaMnNSh/Fqqxmwq/scMd
LFyiMgpQLvvVooJU058MomtLPDwClkG243JUrsSH+UR9stF3TqpdhHOSG20oCZ8b
1S1K5uVsvze2s/m7ZJh6qP1KCjAYD3GEvYHYXj5eZO81AnQq7/gbCgujX4SQNMB6
zluBFs1CbtzXIXrTJC84mWZUjSqFPoJchZ7xHwhc40OJGnuMamTxjy52Px2if88R
xXdAgOrUmTiwVz8XfTAp2XbtiMksN6Pn/fEKR09PGTiMexix/6IAQy0C5elGQD0o
Gddd8FsfMNn0m37/vzh4djslnp/sDNAM+AD37IxZ3QX4QLhiJjMbvvHbAloBxF6l
DtrlN86Xr9i57zicizHQCVd5NfdArd//cVsUkVrQ3vrZsv+Vy3CNLh3FzwfwWnRW
FFwr2Frcc/M2jKSBEH1mz7+rWsr62p+wn+eP+a/wlqAhq6GGO5yp2NayeOtUkQw/
HqRJY6paVhd8m1fCBoeKqQuNinZ2WKP6hZZqveIHsmOyeamDqr+hSMW6ux4f7Nvn
/7RZuxjxOL/1DIIRhboBpeK08dLhAWp/ouMgc8/ZENiCu85n2AxJGG1UC3VRaF6W
l9/msIjK5Oznx64H8gYR2ZOhZdw2ru+59xNXnOg3nH+fdTdhd1gHNdN6vjg7h1fl
4iZd8FGj4s5sbsvawOcSTAirNBWyv+4/qIGcEt+CY/937AABG415x/FeiJeSC8Ik
qYEAUp1ryFxo4L6yz6MjOnj22ucWhqFkiAB91TonEvIzORsg3Ppoa6ykUYOhXkdM
y3hLeFY8IZ6Wkjl7Ig26pO9y7oyyoSa21CS8iqwya2lqrxHgLia15F+Bxkr5frEc
dxiCstbOm8ujmpKYXIiZnw4LOyOEA8uXvuMQaBE2+Mw43c1FA/1MN4koRXPrbNNp
wGv3MuSUADuN2g1rZWqxedufhULRtFSFtDYoDVJU3zNOWoHTzf/Py3LroHZSZMKx
TP92t+6KvwbURb0kq3w78mZpOEwpFGIKdWIJu6B4flU2P7HnuO6ojTFeK3BToQb4
+TS9dcn19D1Bbfsy+eHwV85T2MMUz0BMQYVYa0i9YwdKWcj4vqjGf4n4cuZrgScC
lHRadKhdR2tA9rL8ua8nNbjo6c3M6kV27UBjfTtmbFlcRnGJ5z3k2fR3W1UYYg+c
/+dLabC9MTcKbhqYp48ukDCs8eJgyarUnEbLMOSKaEZWk0J7BSySm4oDzilOgura
s13nEBOTbtiGKAtL3Fd6pO6sxV6RYIdmZsT6liakHs/dR+4gTQg3A/0HCHw2OuSU
balDrCzFLpNm93+3jLJo8pyGRVJ9MPSUHf+PtS9lBfOAcxA1zkumQctYV5YjCBuu
wozdpXpbb1PHX3AOUYi0ZnfFZjvmF20w4yepH8t5iqWaAcNJpPBNZMJttZZW6HYm
xIsc834IdMSjohvBZORYK0jYKaKvkWchVo2MvEWVEdQ6HGk00yAxQn8TDV0Obg1+
YOogu3TDZgMiaAYT1Y70QrZb1ui5oFYxapvAuJHEWR2seLkubOLr8LZYaabQ2kfI
6Uw0gE2DAfxqdgC4Vnw5NO1nCgZtNckMrtozDPmOx1hrAQ11VlyHMcbmuT4yKxHJ
I0N/eBOxX3uDSOE2hHdjnLewyM43c/DmpHDsWbrnMZiTEdd66N7pgnUBKlZX1l+H
N53ID570JcP2isk5FKarVfL+QXpief/YxlfQJapIXO/kkJKx8C3dVn8UDwFjXGY8
2+qeNk4+mwwGQdp+o+ej4LGdX3GhYDhEfo3fblDXVe0vsJ3hS8Apdd00/lbhJa69
yI+zqP03ClSMNrTy4d7Wtg0A9aI3dgEScS/VS31G7nfVsGJ3B5OmWY3QxiiapeIF
RedAO0ADvFI6DbXATrQYAN+g9JBTqQ65ptDs99R9iynwnJbK9rMHECUzT5bJLxLZ
WyChwuwhJbKBkiuPnpGsA34xjNF/NPhUy80llaIDnSmNfrBkzhz10tdgoMBKoyGW
6BBK0Me9SMIpIiexrCkPRuZU0593p3jI1Wl89ADS8u8sNA6XoSFTca7XZVra/1In
LDLExvono766Pka5EXzRoZ1VzwTloZtFQxavcHFU2jw73FyH4nzgLPItbdzq+VNG
k0uS6jfK+AnCwbbowX1PvHGg4NBxloNxuNTgqIfmhCD3fvULz1O22c9LqaAO0Vid
mbC6mBw2nWLIocQKrxtrftDCDq1v2O13+Yx+7bFZ5lJlTw5xfPU9vZfLo9vVV0pf
WpsH+k/j3eLZUCfAGjsULAAVl1YCayZ0yWc8L+LNCXh4wTlal8ykY8oeFz1UWyF2
qaeKXjGN2mALkxKXlaYOPL3RlqK7oMcP6tnHvn63IUMNEtHGUlaUmW+pbnmEaOCt
jTbvV0H8iO7ANJ3jzIPgytkyeVVsfVyvzwx6sWqVnrFGF0HLUvI6/dhKg5Qey1EY
GyaZdEHLaN/1cRmXOCRITGzihsVZpEtNIdPWGKLcur0fWHH+rygWpKjGCSaeoysO
piGDk4yPDtgU2G+3e7BhYDSC9gE0vKL6fMU5mSt5w9UnwSF2p5+ehsZ+0Sj8tkMo
oV/jhDVr2e/EXBGN51f1lNtLSO6XBrTG0L8E3AQ9w2dGnVD3nb6idMZGq+nwk0wy
0Wyi67+OMrTs2hZDWC1FeeIgctd+Y22o9sw0SCoAzBO6RZRCDj6c79G5E+WTaztj
jeTJ1ArxiY3C4SL7lGubDP/mAUMVkGNmaHhCV3lJjWQ40PoeQZBHEwKxIOdVZxa4
5499nx1vvPAPVQsE8Q8DVmKlD2zw36NIZkZAmFl5udBZSqcgJsEhyi8yBd7z+dxI
lTuCfwqOy5IsLh1WXIKrFB5O0bMLCt43nsE8tCd4yHqgQmbOkhn+uImN4gE81taN
mzPWePyJ8KjkLVHnevCjN0tHIv+PWfn9cDoStPoOAH7ItdnEVgCcoqxLn7B7TcL1
87CwRH1XLcuOHniAGlO6wgvGQwSNcCTr4rIL4U4GkITjeSfztLwZYPFknzlKe7n9
p+D1b7PhYSYuv/4sM7Ti31tVuZIXiocTWM/67hH56joYws0k0XTtiRJR4LDWHM5J
0q52ZfKNziQ9oeXRYi0fuwly4pPqSukhk+kc1d/K7TarKXQOXQy4rHvPpZlgdmSk
Iho4gEMML/QMF15OT3MT5Jq6aB+wYApyhsY/INX1qNxI3gFRawyvhT13bfDrnLbe
5o6X4CmueCBAdpADWOoP4dZMWGhSNvj49gXsNEybnM7EROGci5SG3Vsj10H1B6hF
Eazg3hr2r/GYweyWbxPMpEKERiCkW1O49+MTyYVZonNFdREdTJkaYB6WMJCCz07b
FjfGHN/MRWlfiJSf1I5NaJqP3Rwt6MQ4sDKRqzBGzlQMj15QGMw3DTDdJ4BrGlN/
zlOqoufMcJgDmxih6pYDQGyqlrs6doeLFahqPjchMbY/0aQijAQxDOh56kTxRU3g
3MJPY4AV60pIv7t1bGF8ORVoiSbcm8oEyNT4Xld3rqJOQ1MuvFDzhuDIzBcj8MfS
F+lYX8LutUUL0Ro5JPZABJ908skKRyw/IyX8mNGSyy8OJVoBerttnobXzGCd++/b
9vVhF+NpWfRzns1RQkKsqgI9FdTS1O0ijKxPOfG78Ncmw4S9mxNG8do+LYdZf1cL
k8QJY4a4uFjGZ4xDb8gh/+IguienO/wzDYBN/33qBEMP3fy61ok2ubFcI7jTejRq
o5J4MK96PuXz5VLM5GgUOsZI7iM1VVnnLB7D/KTkxjw3kIDuteik/CEt4/Q4Yu4X
tkvPSdzB2dnDPrsg2O1FEOt+/SGasBf5u5/+we00FHI4vrEDPuXUkPfsc34SpgIi
pz7RMnpwlp5lIOX09NkWsYXMIKhAOI8kW8Cprkzw1wPPWTjandwJequldi9XnEwk
X1w3vE7tWsKvATr5erpvpR5oahMnEy9EXhyWBBKmG6t5/uK7AmbXD7ORi90xLRHL
VTFWyF6vdkYUGqZcfPaCu/VIkSySyTRTu9weALRF2VWc8anU6X1Wy8qVT95xBP1f
oUe39OmttfGVxTHZ84tvlkK4i5nQbQjbw1gw5aG8ATTjynpqO2OZYL0NQPZXPx+v
7ANAXuQRhpFMcpjGWl/7cGmzqRr2VHlapT9eSxh9m4jr5eztOT1HzZTz93d7ttom
Y1Zyqvk3YM0RPrbNNl22VjC79vnK4NUydt09T9jm2y/IVYqLgmkHw06pDO+obT0m
3/zKPyR4C8CIDHIrzH2kLUcZnFqeqgz0XCT38ANAMOKBzDVwQBB+eBCYyNakC6q2
WRq6dvm/krJu+AvYrAcVNp8551lSyD9z5X6/cwTqcgBhKbIODHVG4s5GxdQRBjZ5
mnBMojqgYOLrsa4xHg3VgFOOR7nGo+GXDRMJLlf11k2JV/VjHVxgOmnHaY8/7S8G
ZzEttiTN7WpUK11rksF8v3SQ59P1tMrVHpWA3uLVK6lke7c0f34McG1/mBS9spP0
kh7IhnNfmmjrqenyIDkVs26CtpcnQ8ahLaUL9XB0NHmOPyoWutD/4DzxOhuk52rW
GaKn2IBGNvmtbYrn2SuM8jq+gUm2G5sXjRBabVppi2jFJFduLQeJZetO1uAJr70O
PZd9FnTCR7cTd1oGW/CEBLI+IAKy325y3YtHp3M4xw2g2Filmz/AtBsmuIii47Ev
GFwXW3oTXFJIbAm9F8lIjbjhAfh4ZrVytnC0EGtOvs3Mbz9Y7UY/9XmJXMsPtGRk
fZCOdbE7xIX5t0OIbJywpjGNZ8Tcp7f01AmBKgGP24wRCaP62qCtrgz1gvnXYXzv
i5y4OU3XWFiN0iXh6NzQyoP2mt565tmluRtaaAEwIaTmO0mRc+jiXFkhUWGGQ7P2
xkDFAeORmrvjuszlcpPJeL8QQIOkOrY1HLXjewVP9hvLU1K1GYNhblg2vGdeYQLq
jISzenYQ/MD94i7PhBqmtx/nLLZUhS2QXtOJgWRVunxMYNPj/vQcOWF0OOTtc3D6
vV7AYy0uAMI6dSobiqPAnYs6pimwjhV2roNKVW1lvsMJBZMgKTdZZHFlxZ+DCvsH
yTnL6gEXvNTy25NJhjtkN2/VsIHTu5ElOetVeP1JYrA92nPL4eNA0MIwKL1QEdZi
jNpOAzXAuCqTSpV7Tqtw9Znw0BuSuhmt2aY0R/e35X7TlS9qB/uwMXCek9wk761m
UFdmKsD9ZCrJ45KUuD128EkJxOWnLCmSPiZo3MIkap8b1DSzoOvISwFAHN6YmEFZ
Fdypu3MPCcISWizo0yuvl+mVUxo3gf1iSc9QU4grdSUhea5liyP7tXp/TLExF7KX
cDeu5zIgFPDLhyVWT5RNzZwW1DPK1Ts3lzAnt2plCwiSyO8qW0xRQlhx29iozhN5
r4tpFW0+4bHusAFlL2RNl+H/s2uEaEJRY4YqBppy/yxGyQlsqT6ZRrKd/P1dJSXY
QY/CZRL/JiV14s2vvbNFOeC3FDsLC5HFvyONcET7X4bw4fS6GjDIrW8im/2OKeD7
x74lGdg/SRw9ftEerIFK8u+prJHp7k5bWctsECJiItksSHRg1eAmICwdWGfl0mRi
D1tyDx+6OxkrVm8DcC/TFO4pkPaxw+6p/RSFYrdP707AMO16CoQAvDaukxauwMDR
wkc7UywwvX2H2cJ4xEb0+aSeOwkopfNgX+SPESfolXlUzC+NjjgAv5boiyXq9OLt
dgOG+GrRNHXTYdb/FwvfmJv94tyI08RWkTRXKrOi5TPmCft/dPTce6onEKK1shOr
EJS2AGLjLNPm4wP8huvpyno7OiEwCfm8y5ajAp6XnaTMpMwpKnnn5q4frFht61k/
SyoH2QaOptElNCFO8V3nniy0Y6yF7tKHmVOnoiZZatr6p6TKV9fjoVIqqI/QXGKi
CPrP40JMrrr2n2Q+XMs8i+Hd+57nRAAmQj4zQSO5gVzVgXafmGF7V+1bQmseD3oZ
uQktTls5z2svBBfZVn7j0pxQqfMGCQKvwrPZT5jrIgu/yC7F5jLBU5+AwlR+Tm4H
CnevawYFuqO73TMp7cI6XwXIox7rDa60tZCwsyTaJFtAiWjylWaC76KDq5IFEQPi
Fk1qmsKdmFnW9A2vM0rZ+hW6wmAiZxSNvM80emqNUdiVTz6wcvPYytaEfGfzyed8
8E8J8oQ2mu65Crrj6xPlcHcm6G9Og/Za+iMDMI5eGUD2lSkG2T0QCJSPYxFW6EnY
gHr/k+aXYLR6aO0kio/gdIxdspYXHQJT3yD+0ynGLdPGSiQ9DOwsZs13sN4++JK9
rWfYECeFx0v2egFQOHpAjiTNvE647QbavIsQB/CT7MjXCl3WFKn4N3gNI/vmXC9/
iatrFis8kta9MWNspazzCoQTiZUKPMJ/mjwlw35PgLquQxYoW9eD57XU7Q2kSLKQ
4uAYJLVb38zw/Dk6bw8JLtJJh629cCxSlaBdkAjDQAiQNGUC4sJR82OFAH+5jhFT
9DxfdcQa95GZyZtG/YMgZliKwTik74RIvmdYY0YLUsypEet6JFPNq3Da/efijjKe
MqxASqK6WaNM+SkyAdECuvix+69Q+O9FlxEjkn8vaasuKpa8p4DLY9nXfsZWBXL0
Mlcf37G2pBRyNNlXjAPTaF7TzEMe86XiXV2h9FFOmGRgKf2tCClQMVDHfu4sGjtt
5csptoCeRpQrgPkfT2VfPMnVLq0rxEoggJjaEcLvQlVyiOKXZTt37gm1fZE46Qr2
jobkaqet230/s31+PBzkpMCF48nHcUhAcySFAdcFPLLa87AKYH5GOAugGX9K/Duc
JZxuTQLYOErGC9DZXsLr9hANJUaHo7Ck3qGg+7ENjuCV7mAQ4jNa93N0J5L+5C71
zlcVsWmFB7rwBgw2mc9kHXV+ZlPzzmTbaBEzx6VLnR7AKVnMHzQreJP01/437/6j
HkbnIn+YkHYtwWjwEc2AVVFgI4zlpYji6aikD9ZMO5NBQBEoU9JFbv78NFB9AAMo
BrDuFhldYiNAEv14YP16p9ed/8FjKsf3t5zTn5ohhbIaf3Apr1kwQqzgm0mW0pdY
ks1r8XnAsP30uPX3PMKAf/kl0Sew+qLec/TDV0+Bcg1v+rP+W+3G30C29Ebym8ND
PaiSHKXGFd3sStt8dHo3Xa75+BzfXoljDJJRJz/Weu2aq3xhSsCoLei0R7wTX/Gl
GNHB15PmuTir1iBog+gqSVDG3W/3QXnFyEz7WAgxfCJKUMniTzvseE8Z93rzADh0
IjK0YFA8eNSP52RqlD72ayoe2Oicj40JucyEQMnX+nB13vB5wC3otSOazpCOXxOK
fJM5XgrwJk8Spzi0B7lGbl58N9kQFt4gJPiaQ4g/9/tEa7vEmi9zB8z1iaF8KMI7
Tabu3J6EfhuXNtBHVmjUzxRLwBQL4Uqb1SImUp9yWDAZ+ngzKdELDj4o/tuCHbtV
sNpEnOSDGPmn6l6lZXCJVSCx3FEzWQt2OrFSppOs+2cnTZtbUgZxOY6ZRAHnmcA8
yChxYKWqZfl0kXzMyxNTM/Kj/0nl00LdF/VVJ7w7yp48OmwCUpRblYVZTraz0aoc
nH4Z1lJGhGnvRnhP8r3AcULzJcobNWMK8nFnjAD4yNGZ+Ap5UaJD8BbzVyQyr9Fv
RR6qtQ3NLj0U7ZXOPEYzhTr4HLn1PUX9qhdPapGh5/nfIQoty28ojFV7CZji1tLG
0mKQXnf7722kJFPeq1DiGaNW2cFI+3EEtYMERb5J3gkNOntmmB0DQjcKlGPoHutC
p39g8ojfpNXVA8F5ylsCErt8/QWvj9M5eQM0oxyY6hOomXczsu04NC613bJN7Naf
bQ7lrq2pNLchrh8i1G+vMQxX8zQI52GajnCbiFWbqVlT8Fs+d9j4r7HEjRzzV8uJ
yywjuzMhX9BS6rEwebbFrRcaN+rzjaMwcasH0Bq5BsVuHLTYdNS3m4lZhhbhDxQC
Lumtv0RPLc1goOC0kMrGtl5ONiKfnHXu01fJXKiDf+vrAlF4E0wNPaaDI8/ducn2
268vSLBSW+Igg4XVt/gPhNRPSd9Z1zZ5QFYTZWdjg6AKEFyYyP/CtJF5BPYdHy/u
wsx91dZ7Gyj1Yx9kcCn3BTqTPSahQpboLFMr8R3x5qYUgTEHS1L640VCvI0XNdX9
pnK2N8Pxa8v1HKeQyL6x0gh3aadc81Qn9XT8cDwiIGfqFsuz6UsC/ezWIXKrAMQL
6KCYb45e5Z+L85qbHaJvP7ceP+GPKjAnW7cuk2v2WftVMgV/gfa2j0rA/Lrk2lip
PYQyJMxHSeTCrsd1tITXn/Kj6le0QoezVO449czrHncIClkl8FIuTWQ9npOgUmSO
IlIjRRtI9zpNWuVe8X+bWPigxuNMIromz3f6lSfdzbBj2Ua1U2+vM+I9/NBV35/t
jvlbZQPh+MgSsD8xI79meX9y0lQrWjSk4MsH7p4drSx/LzrTH5WSZTtWKGJMWeMG
AcKtxzM6ULcrcOQ10yQcOLX2K0hmwjzfhaTzkmd2PPQSqRy+vb795jFPqzXU2ABI
gP6ASYLRMGpBDXqobd6EzXkBtjAYJz+b28pSgr/vNw4pmtmTQp6euUL/MKnGYWMl
VHwtdRQNBi+p2m9KKfQCEMBqrvqQTgDHLu50WXJj4I4WNBYU84/XczkzTGLyvC15
ce2uQE0Ro0oLFgrKhq3baof/k9h2zpkYN5Hia3EYRq6GUsWDmKTWX131eHSVRhbL
umVUeG94G2FWZJm8Glwu+OVPJJwMPc/l24IByy8eS88W5NBOXNpd1iU6pxCKXncF
aF+yxzoPWRqESHN/NTb4TY0Nkr9lV+I2/ZFWgxcsavvyiEsLstoUma7T5PXnx+4P
oVc+l0FEKBbOTSt5mx9rHY85ZCFcFQeFNxmPDBNlrrtEC9Rb9AXTLrT40XWcnavf
nM66dH9dh3t4szQQ3IAxNAWtV7bsD97rWXfkwLCvwpf0j4C+8mkMAkvjbHo51hED
4dbDfjZ40WIyyM6X9ydULKr/GZVx9W3y0qHmq2F08y9r5HU6b9rRc/eI+qx/VSz6
U63aJpsPAyxpxioFPbodGQ3vN2sa4+mOu0p8kPASaXRwX5uIX/YP2SGdC3tQkS+S
k0PyXKG+LahVVvET+mmyGyGXcOKNCe0eDgG3iz/Z9TovfJiyC3y+iS0+WzGh9xb2
Nq5+hIyGDjh+Of7nZIeA2xmgvKqh2lVZ0JN8fClNPRb6hSDI4Ey8e8+yGMaznHe/
N6iM1bnHa8jIYq+ZsLi739nxnsdcoJsR44X7jDt3Og7/3HclenI4Fb0eCXPldS1v
ydX9BSJXKETHO87eBYWt6NxlUkx1d7gsOpf3WkOFBpstWPKr48v+m6/Fkx8qeLnn
R1+xVnN+qD68W3/u9PLK6PBsyj145Y6jTW8nTsUqxAV8UdgV4YiA3vYKIrWDdjjZ
kH0wUwIRo3NcoX7lbT1mjwfCtqmG3X+TDGT5KdpzokXL5pXST24sux035mwNSuWd
vxUhBgy4Jo7+ErVV1AVdxBTdiFwZUJs5hQzivHXujDA9Z4xDHHH5K2S87eDQw1EY
Wep2TA924OTNA8dQRRduEPY7VOQqJgcGZIpXR2fjhit1ACuTDq0pJl+D4dV9feYv
gVDp1aLOSGYZ/qmBE+j0c8slGUSGaPUjsISgHcI4X1jMX9Ta5FgFm31E4Oa/0pkS
ZYy/fSdfUPI++FD39TGIOm/IE2v6cdOv6b3fm/k8lfXLCzprNZUk9hrKiNznEvuB
00zmfXN4df+fIpbnqJ4qxaS2kQ8EyMotOVSlNSbMlPaphmtktvsNMKKsE3sjBH3V
PnA/iDz0f1PCmBglcvHLGiLMABS2WcigsXKzXy77qcAOSsJxlnJ2qlOJUGzCjSR0
wWw63BCzgqJn0cf0DXV/qJLyo6m4o/n5c0RfEAYOq4eK2mbUbuJgT2S2HUuAwdvy
QGZYGQb9gMfuqBebr6CMmaqv1XGJZJNDLjdII0cPp6or2gwNpbMHpr6DkZdDCQ1w
JamZwh0T6c4YHR4kzVBjDSm2jh7QMTbv8ViPt0zfwk4BsAzTz+eUn1d7wYYv+jGZ
rmMClrBkvshu3/d8ZbjI6fBtyND3PfwCh2pT1fCUZV+up0gm1iL4HmP++nN91lDk
jKVatQ/rPfpDUp0KD6wXD7Z7YUGqB+M7EXW9kWA7wRthrTdWMe0telHXs2kSjIk/
TDykKNx3KG0IyiJPaqn9AmsH3s0aMkHRXiUt9RCHbnMCf7nm24DivOQyuOvD5M6r
e1wRK939kUph/AOj93hnMVg6QaAEZkWyi1BVRfSeKuA5hIzFdZLDNOqmoPXCCzUU
PPk+kHwD/rYSiDmmKhnZsyPdL30Y/CmKvcjEmWR0r0B0jFRFL3HgQO1jQbkwZEwd
8R+BWNjCpsjWWfuKXIfX6O/879TSovMpi7bKjHtsKabqLJZQd3mgdmFjUxaFGR/0
ePepShO6xpRR9zbTwqUihB/nYrCtFQ3vvOxnBSPpdjyeR5w6mVfdJEzCthlWyk7B
uQzlm//oLwz6wq6IUjzxHfA0J5Fn5ZDOdOfSoe/3BQBYtl98dgvsZNVWmYSvfUmX
4OY6xtJo3YT1gbIInxm/puG+xYGF+5elQxNQmVXi+d08jM7Rq3zh8O76zwFAfXO9
POtvnuFEmsXiu6HTV8vc4TPYA7Dpuu9aJSOQmMoe6OzVpQs5bKfp2MZsb1msu9f0
76y5XIPiwO9SxM9/dwORMu92SljGjdDFI20cufmExZIt+MLRCUETF9153bZ2uKXm
wfC/d0OCxCOHRjtUWX1saFdzvB8l1wP+236V0mamG15+aCUKJV/do4K7NMyUQsg+
IvnlT26L36LREyccLONqCwtx8C8xftGiZT7GBw9djLEcNapx/lvOCrwT693WVG56
cTZlg7y7A9Tb9BYxyD8uE9tTGCi9RHo0H3V7+mvvWFzVcMtNIOdOnHTb+8CVQEcr
0yJsDoaYe4DG5yCAhT6jD6BU9MEdVRusDI6ZeLHQleIRiqZSfj1H0Hw5OC8Zq/wf
wrVgxHAF0RFlrKQ603YztwxPC31jLCbjU1pjTHnra3hLJPNEUFY5IfqFgHBZLO9p
RrBrsJvt4J1MrxSJQnXbZcjYvVtpj43zWelYANJ3MdHxdaSbB3dyFDH2GZz9kTNG
UA5mKUHsWyX03JUvNf4HZDGZT2Xl0Tnn7OwD1BPQ/6gpXUs1ZLAxhxC+XAu3PY3t
/XaJDoJvprCw0KFgw51KaPYK0vn5lQmzYJ4S8Q3UZ5Gy+TZKvHEq76O9xUv0DPoW
pUEUCENTITfZqnh+Eb37Ym3AHGQALe9GZUFVqjL/uIA4PU6XOqssLpTw0MAKRU1k
2KzJZ5e741tjSiu6afjNklXKOegWNBzOR/9HWY1d6Wp/covpBX/76V2lIpeGphTh
CX9zKPYpOlidFfK1RIt+5q1/qw08/7whVJlpZ7KGg2P3l7E6/s0xnp6OwsF7nszS
CEDyPF5eAsGfXASY3LWBAkDMS7DqXM7Mj5D1NCT8VRt7X8jgcItNSGQpGOQesfv7
wHur79eXeieEAmhDpQhYPgyTUTXr/jto1dGWZzaItlVxA5qZ3og6od1WCfg+gNl7
Ua7K/lFn5v4LAy04MpaO2HfiyKqsPF9ggJkqEQV2041tUDiM0sQjZw8+pIfe8hVE
rersYY7sFT2zBzRfY+/rBT38ptTgy1yJDTwz88vORpMPVKO1neLHAzHuPeqbgsHc
QapUon1UM8pao/Pwvue0PvP5MG4vnteXI3pl9nLWGr2X0k3YM9bJxIoXJVm0QoSY
wXUSFt4a/K0vKwgud7haC6SxZyfQBAhC+XUT7PHYBJQv1bVmcrer3vO39GifThD+
7Obrrj+qCQms9h3WIGSBPt+PLF0rJiS2BBjLvEi6PoedcVREk1E7uQbYStr+H41H
yd9JviEJFpoTafDG6xHMm/tj2Gv565dTJhs8cpgEHyOjlBTLrJNLjcI5jHBZ/XKG
rcwAl+MFJ3T/+D3rnQpcJd1VI07a4NmGC8jPVhgan9esb95ILdjbjcT5Q0/n6bNV
ZICOggCimRAt8FrIauUJrKYQJt1YJEOmpgOOQgMUBDwEuBopulEuOuTgszs/Euv9
5nGCN636/PEaKpwKqtRVIdmqjXDosnhM0zWAatAqM21WCL08O/cUJPljHiQ2KTk4
ZWeTjLE6O7pakrARw2PUUkErQJIETnuCZw7l6aAfRp7bzGb5vgSQu5PGpc0t+PpQ
RDubXYZ6wchOmW7WdWsDDzyzSR8AwVdEPeA6fmR4J89mnldY4VKyzBr3oGh0O+5l
Wy4TFVqeDHOM4taRRb1n58sCoDAocuGDUCNcbo169NggFqsl54vHbCKNOsQaUDJx
S2jkFqC2D68n15LEMEmR+KDLDpvLakFHhn1WToRwfGJ2ANhV7HGcXqdnV7DIku3J
1NrwPeGdDxkMStiPAti0vJfFTOo8ufshLH1YLaVxWLYKZ84uMS0YYBWlcTk5sWsO
Fk/0rKHjiyrkMwaj+B+OnFso9rGw8D6PL6P2y8lHMZ+TH5cnohTrnsR2LzHTIQSp
9WQZXxuyNipsp+ZDku7WfzG3SuYTG8ddgVlA38amsAdxIFsp5axu0kpEXNRa/LA+
kvp8Ho0sM0aOlvrvPREC3RURKh4nlzkNslBLYFepjF3HpbdqqOC6hLUgdOM1qg/i
SuE5vkugBUInoaxSRfKrI0DrWZEJzFuunztk4tQ78FUR8hUfM/QoxNh5uD+8igC/
BFHWw9HUyfnCOCv5ZabEbd4jkqBoBB0j2DJimqFrjvxpxNzI373ek/GVGIP76zTL
mUDc6xOC9E5qCTDs9NZGERi7KPTQeZ3/bdOGVNd7DucAKurR+YtOJpKOCD4bFFXO
8+jQ0WUd87AtBmjdBVnVKoxpNL456TmKdM9i49V7hTRiYX6653y+L8B1U+6Um719
ig3rAWltZQk69W4L3IoF4/4Ku/NrCKpCOHLrJ8GWN2lY7H9hGXpHbpNlQ6A+QkNY
q/xFuC75qj+9GK6IOQ8+OeicKemIe8zrms3yprjK1740GKOyJ4wt2Lu3sSFuauxf
kZYiqsefCwTutuHC6zkcHI19WEHX1WSYLonSL5UFTEE4S73/kvGA+S7Py4mmaj9l
wcQboah3XWABu7D5suFiqaRV8ZpxUNgjyfiZ+rY6P9J80c7pOphX7BC2jvsFNLH/
DP2hCGpssXbRG0pOmEKQ/bu5izYzGQYwO720wK17dQ6K1dZEpNKNpEuKR8xA0/5j
s76c4euOCCNiRyEnaTZpxXFLRokr0nDLEhBb4N6KUHsORvcRfCBlfavlzlGPwqTJ
6Jj6rBKdMgl9I1dadu1MG0RpPrr+eq+N2Q2m99UlPU5Vld2iNrV8BiCWvZlaztYD
TgilcHkwAxmmhP8unbddhw+GvxhdgtU/oMmunBUEhqCTDTZVs7ghwaOqtPQ1uUaT
uusuPSh8opPwgihinIV6HSWc2ggmiSPMFxioecicKny1LEMDQjnuFtbEsDPSacqp
87AI96RSIH0KbZdRlgVAexEsdjlqZtXhPcChohAzOUFRkdYqzUeoBi3G2CiB42vf
kH8aMBR4Q6RiWjVQWiGWT9eNheVx8O77I5v5lyY2x34Twn+LQTa1M2pk4Sj3xaVT
hcxFP6N+DeK6mrheGAuggUw7Wsclhe5ua/dbOqDhqaxH10POsfG2NhF3a+BpseQy
F2QHv5kNuicKaPjPpQqzqtDC8CoNQ0dHTA7GETYqR3vW/U0EsxWCanU1Q4z/utqR
uA1F2YM5X00xX2gXV/BfMP9iG1EqQSDGg+gVqWsEp+OIlhgRgVG5OSL3irsKcnty
DL2eaOiEfxfXMR/LrNqnN+vXXhQmkRbmqFbd400sYRk2meBn9pWvOCfu43XV2etD
5bqn2NicJUyelMHIMz4bMlhgWcLwROzdml0YeoQBFvBgAV2FOZsgHXlPkoTh2IF8
qFjulz5TVUj6l9Rnf+vzHyn8elj06OC32Cdqi1MOxQcJwjpyZbnzi+l1e11hljKu
7Kn2qAhXS5vTfhIHct8cMFcIgvfpDAGqB0rcCk23JozAt7+o4n8JJESzZXnE2ne5
tOwK2qSaiIlrEZ4WpepXdrw2TNC7E4F0oOG6IQKbvitDdfhwImOMrxbaL9nFnfvQ
HmOclxre3IFTGfpWrW7K5HVa3SJVNMtW0tGUWRd3M/fyCnpcskVnkni5i8yMwiL/
p4LN1d0iwzBS7MhI0fgnZtklZpLb4rCmDsy/FsfbDBRM5ZNVgO7R7Bea3K0nPFQo
5jHY2biq6uVpULu+OjdSI9J25zAxVkIaEyqybol5xHQELkIr2hb0YsWkz/35Nx/7
q/aPpVJ4tdeIVj7jkmcQWn0HoKGiFDklsxsMFD4p+Qgg/f3UpWiJby7Ki713cep8
y6otyA3ZGeQq3+X6m9k7JPpzCL1hH8kgY81UFP5XdG6JOxRQzV24JKrJ763UUBGU
ZHush8WMRqmcXjNUITDAmF45W1Q+RYsNHaNIFNhQYTivP5bfc1Wa4WRFyJv57JlE
S/rGG+zBD0zyp9XbIJXWx5jYevvbDTRk8BS0JlOP1eAnRrH3vr6EMs9jqvyPdL9f
h0SYhe07LmoqZlTPEKC6RqiaRNQWYrs4uSTT4tiwLw2m32lz0B6Hafjaes0fWJq4
/7JM8DdW5xiUzFHS4CRnUAnqQxgUoTaKt9KyL7CcASrXMSpkUK4+7tMi9Nxj39JL
GjHfU9d0/8K/uG6E1sn27rYuPja25NvSL4fohYuOqEeHYUh41dDgdfH5LcxIoHHM
8Jq92eAl2BJqa1t5UGjukARBVyu3bKkClXk1XBlItyores3Fx7O2VmGcGytzOekN
r+90sxOFFxGVsdMMh9982Bb8BgKI9cg916U3cwUpOftQVgeEmzajwI+8u1ZCX/XZ
KMKEYTRfxdSt53vwqL0zB8m1EFypqw8d2M+Be+xwaQMi0J5hu2CTGtTiv8fU0WGU
cnyDoHVu0JMCBBUBC0hf+QXR8lAiQFCo8BUqMlHlT1ohOmO3fU8rIuSAjs5erhvv
UE0FnqnUQffX90whd8Kp4KJNW/Q93YoBrbytK4FxfpusSnBnbT6ibNh5h89MXV7d
Zq3F9okqvMisVehWtx2SLc6kLtBWbhWBBxe+q2m0/j+YHYnepmoiHiUykNXau0o3
QB0sVKn9SjpXj4DCh39n14BK6w8O3HppotV1PvJIulIQRjvvHkz51mernkF1Gs8r
dPgfd8HkDN7cPcRXE4IQ1GRqYjaOuNXjhSMfkBFX8m2sbqGnZVsEiTC1ZrfYl4nu
tbJa/iHlcwXMbgyUa4hL/NQvKcIav/1ULoxSRRCXJNNqLz4ZvQuQjXma9ku79Qq3
gCq776FtkzhRpcxfYvHvKRamiXcCNGWR5fvgAKHFwSjDhp4SANkWh+VwfipOh7mh
Lyb8iBA1IkjQJPUJ0QtXqgompNVCxTczFhF4gP2Oxt64VTQ8iHe4fZ++e79BjRu8
kM+xxrvx0/C1rXMt/L2vxTBiX65XXUs7ebtEB/g31c3lU2loUl9ZV1TeNht4LObj
klp69xFbPDMH+c2mly1ENLKHJX383fdm/PEOPMGc6PzP5SsLRY20Hby7JV2URqay
oG2p6Oz+3VFlfCkc1FjiT/HS6L73bdPqYiCd0tNN0f9DKbHZb7MDqLRK6oPwRLCH
ltNCo0wgdSkNEUIR6CVAWjsLAlT+fXbCYvwUfbebYBLo7OGMNdvLOX7SQHIcnbcY
LINSkkB3iw1iRRj7dppeEcH539sJbfB4B+mYf8AoJ4N5A4Zrgz6O5MqTT4NuRGnf
EduZr2mgSK1pM33amRopvQ1dZtloMenI63zg2QlxJnnti4XDpYgqPmM5eYPYOqaw
u54TMyRyMeIBqy/ZNxi5e2Fj4qqQOGsz25+m3o7TEmOgNNcwTPLHLMFDItUVPdIz
Lrnc/zpSmQB2jxmDe2R/TIeESrBcQG9Ydhuxz+0sQq0nSAltVxJnHU23H5/fn4bs
0cojvwyeh8eVhrUHLfV1BUAsn72IfJwKdFDQTABKectapCwzXwLgS/k35H2jTJqs
T7fas2jDbbjY3jwPUkCz5o+rFt+kvKkmp/oHxlGUqXVaSLaxIRcf3zSWpt4xF9s+
lNYhfDVYFv9BO24CfxO7uHCrPKdYii0CsHWLNQJlWi+iGqJOXk6vtgtjP0+aJ0gv
HtYLUWt5Wkpq2pe7Qcuo/WrFhxPV4fodbM1xEe3NwrAzuSSjsVMXzd1ln/VrNbz6
2wbX3KiWr8I1HeIEJFAtw1MmCyrcnGJvOCPui+IP3QIhQC/Mmf4nB05CC4wgo/oW
vuHSGc2DcbcCBHnMY6lFcfbaH0Sy3YLwzemxo2CmgxN9rsg1lmfa54BZrR6MzRTv
Icu4MQb/WNHvkWDcuQWkD/wXBsqGEWxznOjwBt576w+I2AW3wa/q3+BpDabhg2CL
NE1YYZ6Pq1Ubq6WCZ7+NUYd6fYu1+yEnAMF6ciR1MmniBh97PH+W+UewfLKi7rYb
D4OjrH4d2DugHA4Zdb6OYw==
`protect end_protected