`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 35344 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
HdytKcppDjja7VfYQkCqvL6fz7n80jsjomyHd4+L+WfP7CQ1R4XGOXosIjG7Lfe6
OOL4fWVg0/MUXgjaL8E171lKFj8NvKjYxDA17U3HGjtXZdB7R0M/1qs1BHnVmiN3
dvCxL9HNolGwWj4stSmfTP/dsXlyovSeH0f29gejqWoJLM8tPqvGPsmWTnsBhmeK
2NMqEmlfDyrxRsx5Zpsbf+L7NvmmBhWcQhBO9HRUrcHL5kUKrHvgjTd48BP1vW/R
RoLpTjAMiARotV219sud4zGyGg89my8LfqLqWTxpSYU2mCLFdODbcUTUIH8eBkP5
+iMjzwjQsV7OHvRFLaoenL3efhevbsaxnZc58h5u+3UHwVauukvGuYm95LrYgAY2
g8MdmLrNwqQXqLtrn/4gFNs0XI/X6pwEzyi5f7c+8ImKzMkQvNEjt8c5s7ypyHS1
6JyJKlm1rfkt/Rx7asSdHgzhyIigFpSVZgBpnfLb8CS6dn9JfA4fd7EkeiZ4ZHiC
MxHsEdVr6sKWkSuLqjCAoDfQYnzMbzwBvwCsxszvNunJksV/cmr2ka87mT3itdJB
KNGE+1DuaVWbxx/kPEyX+xrN90REvAxodYKfpbrDgk5oQPj/2i0HPdywOx6N1Vdw
PirmgzK7f54PzdwGLcVZ7szuG/+/NGwCuzsUGouh90jZ3tZ1bingH015vb1VdpEm
toh8TriK4CJ1z/+g/KvY2IJD8/17Y25eajcGzCKwPnmmdv3YG64OokG9lWkXIL4D
1hYGDS3+fLN88GRB18bUz//fpyCQ2lMa8CNyklABKvpHNUJ9TrRjyEFeTu+hoGND
jMd8azmswX1Moq6lF/t5CxdarqqldqQAO7GtR+ruXT1NSOFR/evgPnIBEnWuJAqU
LhFzMiCVGuVK70rY3WTMXdAsUYrtYrZPrJEufhjC9PRyOkmJK38laPGI/biW7iTe
BVNptrXQ1tSqTMYfn9vidzTSIZsNvwPdhoglKXF5h4/tpH06mHX6bT9epmCKS+M2
XrSvdUwbEfSR813CeSTWH7KN9dhZ+KGFdiFfYKeAmJ8zpo9/KD5xyl+SRncZI7Fx
PrFM9beQlYg1ji2QkV7so0H9M7bm4e9tlGNKzgHxayt3JOC+stGwPcp+G5q19sJp
GMb9LZPdpAvN7+sLwNUjyVLG/6u27OVWkESCIdpWccTc33HcHXYM45uZmOaUIBqn
Wqo15bD1bdhD1R5jpDih90Apf3c2H1eYhKh1u0THszQewqQZqzpS8ObiCTVrbOqp
dDJ6SRotduXbztx3rYSNCbhGTUe171cSLc6jIB54rXRZsVQBN44/i9mOw+pdmH8/
jV6cHqpGjpELg5C/ckF80nnYYPePTF/bzUHEoUXFcqJ6+47dJ1SWUTvapMJIG63d
/Vgh44hOHMfTyt3cwlaJR5lZPYXeJVAM2on//H/QKjzBfOiydguCCbcsZ05cYUsM
5N4buDDqnMdWAOvB4t8KG7zWUWCVbxYW6lWieorFenQGHPq9VSQamYv/pA7ydl2T
GNNC5UMDCXwA5+CqbeKL1dDeofhxkceMcbr4ctuf5V9I1+v2YJWheYTMzBY9oUVb
edROY+JWynGbwADPd25Sf7tpxqVq66rl1plrgruM7nwdKUnZcQgccNYP3P3bkwMz
aKks0ywXuJY5tck7gEB8T+DC9TtHyDSRMwAgjlciUwZSMkafN7N0ee4ZmLUcpJuF
MIv09nQqbwodFqmY0dSzsj07A0xkSGK8mkYuGS4KQ4v4O+FWxhHab8wvn+ok+Leg
FHHuIAoPQa5Glae+G//aXsHmtkg7lkZHsihLdqQUXpXKJvW1XHGlAaDBRry6mGcE
fEUP3QJbj9EuBok3v/KFnkM4IWjJsPTUXxhQ/31uH/fNAWsjDqJ0S3d2ToJqUf56
rh5zp0wcsR5D4k7F5QRX0iAcZ2nKSaCTehx5V/CppziA4Nt0K6e5ChDoF4tWG7EF
AvVbiFSXia/hlX59ydQnd1eRLOoAc+8muMK5rSb3ezdOUBvag0WL/ysPQ+wYynGe
+q+NUOTBggmgPv/fFasbbXF1BtOYvQbHA4ANW6bp+yUn7rB2GdjmOidN6EXvmtDS
VJlkAYAvPVViDuP//VntR8VTnVpw5bPmHrLTJ6gQlnRbGc7Hj9uOGDPdPI2I0vIJ
7/JOh2CBsM4W71nsnfjP0MWssdxtWOOcWb6kSDemXXgHxrw923HNJH1Q4tYb9Xqr
3B0tIIujepCsYkp5Exz8wJszOOkO5pgWJvgxqgM/HMDZCfHn9bbNvu01OzrS+HnM
6E/YJqB9enaU6SwimSUhurj9U1R16EDIW56gnFj1h1Z6mm0i8Dkn1JkYrd387Jq5
5l+zSK0A2skpQto581xUUkK8u2LUExc9s5iz0hhp/3IZdC0x5ZVAAfT00Z+yRrlk
Bb0lTWVXiXDKFj4cU5LeKhJ2l/j7H9kDylCsIwaNJzPgd04P55wftJtpUVjJckuz
O5eDhqjs0TnoyACLj4vclaxcuQ0N+hmqTG2Z7IXt77I3EdNPVE3dBXsq0qwPz206
QBUerHwWgrr2O7G3CNJYJVwf+380qfaEN71Z1PHk/c8OMmxtOarDrV7cCnEShTP5
IMGnT0qsKtLCTRwh2MJhelj36YOk+zfQib9qEdg01WKxqST+AD0QuMq5Xrl2Zupr
V/K/LfxwEcAr2a388G+ATIk/8mnXMkUpVWhwncicKozDHGOASGkQfa8EyPNk83mq
cP5x2cCZNF/msNoKCkEd7KxqjC+ESmylWHTOihactTHYWidysugu2DcfGtMioAD3
SoMfwiBR7iJ75L9z7u2j+ffI4i0/V8E8i26Xbm9uzbbybpXU4wYNvGbBVZGW80i0
2+VIRKTCCXl80s8p58WF4ArMlC6rBc9DHAjccq6JqD/2G9J3MeHM+Pga+PguBhIw
QcrNT3LvGIfHRTPt2859C8tENAAw30MY2U8k+bIsppQ6pCfqotCWnFj3zKWeOHFR
3gGYWU2qKUJ1dinu0/Gr8FSMXDfwHNfAcwjLuFIaR9BKhh21mZzcF22cvL+BizVl
7AWomo1icXn5kGeqEX8fGtMxYTOUV6Ng8IAx/88mbEmAn6KiOjWWDyWwH9bkcpjg
nzrWxwRPJeTdFopc1VD3i44ro2uKQEvtF1iRXv/bu0FMCgYId/LrYUB4DzZ4ZPUR
UpZzcjTAQzsTEWT+vG4Cqbtv1sC/Qm0bf1K3go4tRQ6I8ieWZaCTFCocaJLpWpPS
fvjlIMeUqs0JhLyyDApFpQgcoxcNOvEA9m/7hJ2kqeVjQHccQPVOJDwnu0VPjNqj
Q17pjed6kp2P+PcE6/F252rn4Pe1EN0HUkWRznnScSyaV29bn+JcAVGXFOOCN++h
UYJ1DWVqYK2wl10lIv2x7F9BljboYHSTHZurZKd2ncra1CHe7mQ4rkEXtW1Ezjgo
5WQA1YqQCLV+TBQt0PbRn2wHSO/m74MZ2oupT0dKpHEnRAOnY6JxXsyUlPVU6Rpz
UUpzeAJB/I94U1HEz+ERe0mAuE5w4Ro62LNW6wrcOYNI6M7HyXx4W49z0biI199y
OJNZ1OO+HGUd8X+EaK8kigy7IqhuTPxQsQ+6Ha6i2Kt9EHHyFY7nDVLpuoxT/HVv
Yl9FGFP6GijntoqV2P7Q2jyXhdYBnZAoECo2j2cItJwyAUZmlj2AOqacAvw1WfcT
gkf/huiVDNVc0YQVTRQH8u4CCZG/ayJjD3Gb0XvELa+iqdytcJr4xsRinCpy1gs1
iwLl4EVuJjW/J5J0fRs8yZmWoay8FES+z/75oiWS/IJ6uHg29NM79VQb8vLC4xuw
C80/snGBNL025+jIy9NmWUSdJ1dfBxwG94qHCOeySpH2gxKPkcQBdFrd5uYzHpy/
HekdEotCRz8UdDkhIKmIQ+5d6VFH02UlLrQrGhe39u22x/PS1gwbHrFYakjuXfJj
6jNGmMjW/oDJHonB+sYxVPasvAK8wq39j+na/zNQxX5/UlQjQq4VRyPny43Jpt2c
+pCE/nyM1M2B4xTA+kKjd6YhggNd1QfYvb4rTWQYjarIDN6T2xvhikwA7FFxUjuV
vu7c67W9gYB0KS6f46KPgHL0c++r/ulxLGZ4WgZXbcnr9XlbW65eM3s4boa3oh3z
klJDae6bJDAyE/DCeoBswS23jh/Ec6vZO2D9H7pT8T44LMatyvNhnl/xksObPtVf
Ti+ijVhtocPmIPKXKhpeljxh2Jj33zO7NLMHyCdJaTfbmilzU8tGJIsJkXA18yUa
ZRV5NpzCV9ZxUUEUbWqN38K6IqAw6CQlwtMUfkqKUUineL5G/9vCEBlCE21pGkkV
z6oPRC075GdwrEz93iuMystHZfE3jhiO01t+ZI4nCkxD7pC7HaatPd5mJFBy6yYU
Zd8Vv2JZFTKDSvOnimUwmw8cvKBCbO3fuca+dRWbidQaGU+O9xM3xN9bUPwXxEg0
zSOngn7dYSKWPfe1Z4fYGc/sjIm0rKXQaI95YDN6DwmGl0i900fgBMjKINpdCE+k
m/iG5bXh9bIqiNWKM4GjAwA6lTE8UO3EPcs5FAWiT/DJdRdg9m2udst0IxXGZbAH
jumQEk+PD/dpZPP9giWHU9LXYr4hM6Ov/UI1gTtmRziBNZce4LPLP/Z/3m2sUXdZ
TvRu5zpES33hh0yhAQCBJiqG1DDJs9I6q1maO/qnqdpPGo8P3nbti8u8Mwp1uZQN
+7aV1TqzkAIcAp2SQx482eXVqcj0OLHHsiZDBc0A/KMVMyInAgPQ+GYe83yNin29
Jo4+v/Ou/gwfm1J5KPPee8RpIbIOlm3U4KbHnQ5vcaPqW1OIOOjzqbsNz2aMJWRY
SAyfc51DgSk4c4FWA14eItdYoj4848t9z5lB6JU39hC7J4BNiQHynXP6CpBWFiak
wQGxem7crzKAbpiMt4zUhKYeXAylgZBYK3MIQhoBZh9ITFUTggT1bBAecMB1DlE9
SN6xEsP7atZZPXvFLRrrpQKDX3qui9qmo9sn3uZDP/rYgalVDSG+4sAhQR2aYiam
eBSmLsRtw9m0/uLCV7lrDDkbw8kNqI5YraVfrD8ZVXItZQ9TpBE0EggNyU9M1A1H
1NsDhQZ8cRFbV70Ict8kGyWlgQw6pM2rH+uJK8eMVD7y8bHXvcMFdBcRDqsubesA
j/1hL/6x2FGM/8JakxAP3UBhbyUzTh0znvaCcZkOsOWSk29Tt62EpXYEJjuxQvdJ
k4mz6x+avJiJzUw2DB/T4AhGsvMPt5tvH4Iim1Y3rwE43e7lSM/a09e1au0EgTWH
PeeS0Rqwy8IK3gx4F+pBiIdigZ0nVygPVuz5vu/0n/5FwW8Mrjf3zV39gpA2ngcs
Un7OSEVcmWR5EZG9XrxFSpOIFkkTMRURXETVHmyNEpb/BO3Jp4+PXP3KQoeSNG/f
AQ+2QMOyHF7StB/NRR4LTUhIcr5aSzGgT/9kVI372+znREiUeS6aAU+iq+PC5u+R
wVAK7dfRzClcOqcjv5SUEUzlSmaNqTtOQxBtBnuZFR+gwm+25sM+DLUrxrUODY3W
ubvfZZzD+FAJZ9+zXKawGbqY5s9sUSFTrLkzjffxySFScdSe0VN6nSikMtqaabeJ
zIvCdUps4m7MwohQ6qC/YlFAivWEwi/oJboBSOcBvHX3Ng5GSgYT++tSBT1WfGv4
2oAoPlUGjCc5tamXIPepXYHGJj030WB7UKttfRx7UCu6pVQRFT6ZRgcSxoYWgZBD
PULzby26lHgwPQ0yE9whgEc5tTVq2ghidD1NreGH50Kfx37oBWw/ct+fhWboNuLO
q5LBH6RN5J7gZoWXkkf/n7E9SC/Mz2fi6cVOoJkpMzMjALAJu02mWVj8/m6JqKtt
PhMIZXtGaqsFIpXOq54WqzGkbVsdWzUayog2w0yHgv/zVutpURW7jXWcXdqadp9z
P90BxJFSd0b0VUzRD0B1C1K8CloPyh0rs9wO/99a+ZKqGex3GWlRabVaF6K4F+Nz
EM9nGG04Gt67PN0kqXvZIJhfgJEEN7Ak47PP4YXAmpPENvl0y+X91NcGa5lFfuwV
WrhvAA6763cOyzP+2ZvFQQTFp3WPWBBaQuHSgWY9IQ+eCbeoSMCIv0MPPxVJWM+/
hChepp1N8Z3dGQyJUy0zdQ88ZdclJQIooyRXDMZf0lgfMYuifzQKjtRU4eKGl8Ch
v48ctqZuWtQ7gCxWNAm0nfYCEOeGHsdzee25Oy/5YtaboeRydmOGa4b61pBnQffK
Fz4A8SoJ0qiUjQDfExwxs8BNAM2S7hXNYjZLcsJjzIyiYZ/xw6+bfElhhoQYeVKR
Cefin4C8zpsAyS+DxbABwkigiQTU0eFVBFsqJaFk4Nw+o8L55KtVcSE6R/aRA9ZF
ZAMQq/nFbP7qrWfTSx5P0uef7FYpnLzqmbMmIhEG3if4k3bTshCaZwcL+SmjEvkZ
sshxjHQEnCXXY7RBA9+MmkEGkXj3gsbp+TPpY1tBPpqy4uRneg+FokwuT0YceDh/
3MD1uJ5asiU5xPhTkF/ZXT8l1I5u2ibvSzBmGAr6zqE7b+PNBW3UGoYmODFdWQbM
LWmdgmO3XDM+FV2ObcSZXgeDVpVLKmNlag7jnvAltBD73hpCP6klQtafiA9kC4Te
VBHR9BJ4Uj0CKk4SfPt+/NXvGGRO0PwKOFiscafYbH3afXIH12EcXP3myimV+aRw
JI4uL8GKsQlnpjgwTi178u2B6o7bkjnC8B4u5KaM+JRfTk/X9D89rZrG9bCMbXms
j6QgR+5/4WasWxxtw9WDkS8IZXJia/1u8KUtqGXRVc/0ZlYu+HcbG2aWn1GZ8mRe
z1oyrhpiTrHjh6jp63cFnSpI3G01yAfQHHJOAszxiaR8U56F6hVAuf+0Ged1JkAn
47UY4Y73chFI7J/+SnX72ovdtnnx0Z1AiqkJ4dVAx6PlYPBvgic+t79oSitnNTGI
K0pZ9AOcbqOcI4cT0FogUndUcqZ3pI3XfXvqhriZvnFA6r08aPh5538QXZ1CfjKy
5ZzPLj1W/sRca/QTYfQKiYBXAD5hiAaQ00qVoiAp1AreByfMz6pFQ6atDxHDexV9
2Ky7SV0Ns0hQPoqqGRBqbXAGr8fsUOrCAGgclIvkOe0i0MKw823I6FFxLSIb/NqI
FdAHCPQATwF4OyzVIJI+8uIAje+QR35ZjHLSUXVXgCc4Isd9MdBVdu4fVdDrHfAD
RhxKzGWBxyNv55pYgH6QYGDzKupXN3R/uIGgrUPxaaF05OeRHqbLm+ttVvwF2drt
PoQyHqkPzh/Pa9hV3PRvph8eVPGmwBMfF3l3Q/Nk1pp03L23zBWu1zQr5e2RXYxi
1DsZysqJy18JCrAJzAmu52/zxW38aI84bTfJlCDm9l0vFVc9bEC2LnTZR2Pr+qgT
VLWw+prvtcq/hAV6CGfmgYEblDzKvpKrjEa3KRLm5fzZbkRG/ZGnAc1MU1/5CKqM
dQ7Fpbm1kU/tXWW3KzqnzqGk6jfl9W4m14hSolS1wxyg8DlibufdWTv6cIzvf8jp
jDy9HTsxXIrFFoq6K0j4I6V/JZj3ujchjvfOkDM75iEtnfRGSsrQF9VCiFRKoClf
suyLWM2VkD8Ehlhep3nc5Nexu5AXelhlbePj5G2Mg85mgoJjuf3fZBuDmU6nqelM
IdAo9AWiIf/L6BQiae//kDxgNbQ3aSE7oX4tGBI7IsNdt78kv/5Rj54CpiV6zPcE
qUGW/O/xGtgKK5qbmAoBq0JNM9XZKN2nh4JsBuWyErfNJyf8F5+Le/NEV67iQUbU
Ur6NJWtnODTAp1itFR7a43MCC6mbsAjUUHOTz+ki1AWJaGC/6E6B7sYKDLB/Y97y
jIccbAr70eHiGItCW/qoFWbORbrb6MzWLxQMuceC5/Lbzh4PqRQDiFPENsBNbXYP
SO9THHXFFeTLeCS5fevjf6ihWXZGTLRmNfPM2maoMK0eLcTTT+I5XSNT3Lg1hdo2
ZnC/ZPUvmVRtW8ugj2pcNhKUB916zU1/y9Ilbu5uzE05jdkUuv8ENjhyKlSFfQir
SL50utLTXR+kVMUUYgnSckW78QhkGig6y71ojniXJbIA8bidjxA19Rv0hgLIvnMP
L7g7Vc+5jSEnHi1msgOrQZwb+09INkjHg9ZbVhHJ7qfWYw6nYflUp8tq3hFFuFMY
56k9FxO2Lnn+b7TT+GZ2cbeP26QM9i1myld2SdEuhKX7+f+g/uOWOSBSPnvQ4u1R
0KnCX4tkUF9i8VXtd+OfKebApRdUqy+C+uFs+DVzdpdm5NTqMFvA+cRxN3+so6iX
GwEQQWYiNKwSaSEgh2Y0rPBe8HnAsxWAWPOlox6wPxnI7ypRJ+X1AlbNrJk13xSf
FJf8rT3W4+oD80jV8T5aG6XJxYIZZMU8bXtzsUcnXNE/PFHYHRK8wkD0Cy5VaRkQ
8KL3AGJb/vFLAn7J2P4O4CKiEOLRSzwUUH+RQLsMkn7fqY419lhMXCfAZQLFsiQF
moyQC+mwaDnYMNCk+3Aktr2b6LUmWS9XsfdPLu9LqTKCrAdoBFrg8sZ4s9F9FwTr
/UZfUIes3ijdqgtX2Zzwi7ZQ1ar0KdIJkprL42UvYHs2wfMgLYrErY+f3Ot+MK1B
zogB8zD8OshmR8INDxIqRte06EALJ4ZWJaVQ4RDhkuilVLqOQFJMRbmcml0RAgm7
62/ATEy7ccSXNw5kZcFUUxpru1+cfij7F9B38gN/jKFuao4Wn9SlMgtOsuAn066k
pSba+D/rqGGFmejbKNI4SsdAUGOi6sZ6rddTqziWQWTlvk63Ug58EnZ0XKC4PXt8
d3KrB5XpLHClwr63uq3PdrDdmis57Oj75ATcKXSHnwz+Qz9dDh6RLiE9R4ojW5sl
x3JMW75329F9cLwe76GE0FFaV4uQOoYEQ/NHsiFm5GiXP+cKgXzL1DVFk/Ce4yH2
xjJeei8ECIj4Rh12+S1gLjhtjwQ1c0aEtFRYDijka7Ycuu0ZMe870AL8DnRO1EuD
2z+JQofdvGV1SP9n0IIdNLIi0wj2JzTLyD4sWx7kntC/9PnFpifOnzcIAoO1XJ0p
b+NEvnwVOPV0cByqBOlh29OMrr07c3v2t1xgYiyfEQW4KYjed8pLm8gng1Vhtsjw
zUUKgiHfL4VSptraJnuP8siaU1BqsbxdWlpJgQ7drhVXOzKgIQwq8VW6dhin78kO
dCvHCy4fmR1JNOjBAiYYyO9znylXGNbQnOl5bBLll6+dLrLDgLo16Kq3kfS+vKHP
nsfk+atAmoIljcGnmvGCnlaolxf9n4BvGBEs/H0hMbAtKF0wrwra9aK9uS5lf89Y
rDglgnhkeEmPSPklaBXpXI8j/mGpB2Y6Qkct2cGtaTLJtT79wrjle9HqljuxwP/B
ymZU9Trr8eUdZBvPsyJoPc5+6WDMw2OTaJ+RAZESXm19/bIYzn6kN8qmdwUguadE
Md/RC47g/98dTM7F4x7vjctxtOuFnpaaBdL8q5qYV/quzS1wevtmpjfdmqIbkFFW
zg0d+jDiAQKCU0GhywcTzZh8M5EbyibZrrrw7SbBcSUg5dUr56n1pc8obLV/ngzF
iOXmC4JZT+KDlrQNQ9oKbZUHbL5UxSeiMr8su+/tNXsowH1wTyYODl5/vC1gVIOg
2ZBMu+aJ+O5wZW3jeHOafEHBovEi6CL3lHLXDn/ywUw1mRIwDupIzQEBHHg4RUGc
2++f7stvwyTZSqX1QwZLXXd6CLs7IXukKb5D30R+Z1i8glwq596iq92d9gKxtKND
sLexZpW8hhPItk9CBYZMmCSKtcxoeB2WcwecvFPdnyAsHDFbKR+3EbG7jvrDdQ30
rLkeMyJMyK0Lyob1KaUAHtKtLfI+zSo2H1dUe6GOJDgFW7C9zL/qc3xaquT9LsGv
O2o4ACLf1Se0YuH5mSzF+0A6HPc3minQJT8Oxoqr9ts7Ib301dXz7lSGLuWU+rGm
rfOyBSgdxOVxC+IlrnxmD0/9h/n6YfRcJH9jA/6ZzSaug7miznTSRO60uxADwmLL
KLFCEuPdPT0z5jPfvq93sgeC4p2R09tyzJPy8iSNnWpaczelK2Ltcjbbx3R/DPzw
rQ9WBltVJvKj1uifiwUfxLlW72EAK39djM3+nmfbrmlrBBWUNS/60M8ijIu1+SG9
ku6SNLWrgw30rRkPIo/GzGeU8ceC61Ka2SE2/B45/XFr7qcly6kwBp0ZRY5YTnLS
YIMglkE+CyzmVM57W6jg24KCw4Zo1stBN820/tHZ9yzlTCUcIZBJp5/XXPzVVoqY
BtiWjtI+8wiCCbzDt3Jxzof5OzhjX1rkzixKCWVO6LopI07NWCUVA9bpN5Ypsl1u
BG8ZrlVYtYwDHXd5GW39Um/vfbGbIrksf2X3hk9S7mAKgNy7i791OpD6vN9EehOE
3UtCXj+FZoS+7wd+kZI77vc+De2AtF4SKe4hy+BcyFMjK2TED2wlMg+Xp82HhZy3
rjc/ac27DX4vjmOnvTISGSduuw5vp3IrcN79/ujU5naSZiCxt/2cshBlsH8qfG2P
FbZcC+/UL35LykJUwe2vJs5KcrU29C8vPViYKzF85bVjM0LR2f/vqKtlvqZMEC78
EI1UFd5gXBqnKIhKluYhABSGhr01Ff1E0Q1foKwR3KVSa4UJAR3sHxbqZPbOwguw
3ZxE5/yiF8KAgHtqptxIN/J/18b9gbZl8oedTF9QLFzYRGrVOaVzf4++YfX906zQ
oz8C1UOM480c8zvcFumGfPgD952lVoUUCfc/4hC91BFqQk9yf9Bw8TcQQHZZ1aky
I5AETencWnmgR11j8hMXnJuMppT7mkfuQslAV5xWpN6dfjbCQImwhqXEzm4gY9c1
4A5IjGDRAIr7b6qMoTAZMcwF2flKv1ucFQEyg8w+f1JRzAQHTJUs+lo8eOkP0a7X
l6HvlNggRMdCf3wcR2/kvr2hoChGXxo9aZq5NmFRaQGRwe//4BYuNU+Ny+V2X4nU
l9vyEVPMk25Gmj7IZ0LniFcaM9tR2wVbFrRR+F8xPRF/uhVjMaKA+hGGoHf70hom
dhUnNf6n2BYnXNnwlK/WzwIfV2a9xv8qR4c58SI8Xfg+G23aw5twj+6TtZRXMlUP
Tp3S9BgtzW0pCjxve/11SKYuSCDuu+iGgU+RnvnbDA9g/Gk0usuaJ5CkgEC07soX
uFHTrdjHwAylU74ACA/53m9PRs8A1yBS2skf2SWjaGNWH1/nVgNXqsWpCF8gz/BG
ZEOuGFW7Geu1XF64hYcTtPI29JgollBCzboMNFHx6Sz3DyfVUFthl6sBBJH5kcTT
8HyZ1QjmnX2RVnaa8zeqs+04Uv62odNqV40BbmuzaDNHxRGf88xCoubNH5SJUB82
5ob4GGhTuphdqYuZnx2TPQ1cDXkg+JYXR104crNeTKNs5JYCAhPpF7y6Sm3cC1wo
o23Qd/fesVJOPiMBTQJpUo3IRaY5wNHmbdXU2Aya+3ySRpllSoo4H2YoJhG+YBjp
w2A4ZEqJBq3tNmX0VyErZryUrsMbl3TdKGuhVSb6gV0zdKmzEN7iUpzOUgOUPRUo
GhlZtjBG3zop1H7EZcUH4VnY4k4+rIZSNUdJ+b80+0GT3vkNCv649we4zWZ2gDwZ
nzKLHHmcuWBEdEQ3kGkT/S7uXB6w3lwZvV7Em3xQ2AKuCNtLp6C57Pg1drY74Mzr
RGJr/5M1V7KAqcWP093hN9cHjaQaJ5WQ2irr+5fmj/OTl1rjnxRrwiETohyRJ1m1
6q+7CBljX+6tUPExPY8I2uwNvUReQxrvfvLQrBBCTJhlKEZPR3JKh4gA/nLeUk1/
iuEfB6zAe3jGkV+HAgM/lIesJvOlQmQadLYEDSs2mywHsZi9EM5kB64eSS2FbQu8
lF0RXWV4TYiHQK0N2OcPUA1Dw3w4xl9f0pxaQG79beg1KGzGtDuEDiS9RhKml9Ve
GqS1Q/q6GBKzn7uUdYQ3jBswwvBWcsiZQ+nB+8fP+5DRfhSjOLkEN0WHaCwdEVhO
t5aSBGhQ2KKZspeZDHJFzHOpW7r/XJc2QFwjrogF+RxjXifcjy6FblMSXlOigWdA
Eb2oDvRvQatBFkFXP4AbFRZVVAGQJRXNZiSfS5tAZd3cVh0M2ePL8mNimk5r17pA
MWmr2wDoRLiDYQsmUmn1p5rqt5XirDSKYDAhAMrcs5W6KrOZcFikSbXIaShs4VLK
d3ms9JmoEgGGRihqt8L3f1TGbf16kdrBSwJGV531PBLkkHmY2uxp1fAmdJewcvv4
PQrQsBTG/vLMgIKH8rNvDBRLWqM3L6YZuhIInU4RndzE9xFz2hqzMI0VxFgrSWmD
a0EAEqNsEEbr6yUkBc1nn/6P4PLplpJkLWEvuJx8Tnh9m7y8zjfyT0ZDIrTJcSAP
4jGU+dpGvP5v50AKb20tDSplkrFrYbpDymUk/zLZc1znJXPytTeEKIFsKtr5+UVs
Ahye9dxaDJwWdDKrSfiGWNlnxRbqFjnkZ8XqZhLLzptSl76EQC3FhPy7Gg3GXKvo
64g5out9Z/zSVK03gJfArEDJgQZP3qTeZdWHg3vAqpW1BQc8lxs3/5apJpZQgrRL
JB8Wm9A/MwVl1XW6cjDd3SzrlrxXBW6x+Bcq18krTJtGEWS0L+/kAO3yjetzbK9v
GfSp7+JJttgqAu/zz2VZAn4Kwm4phvjeNzwYXKvOhM9G7IwG0Eh8m2y9UeOHfi35
k+aLFmy2Hvfo9zy6c8rKKH44T+gPu09d9bwA0fpXHHlCV6wlWsG9JZKHYjvlXc8e
gbaX2mPD585YqmlAjzrgJc47iXVnvb7yoNYR4aLkh7i464HZF/O20/jz4aFEj4No
Ech+uRUN/tBcjaL1vZwy5FnNZSULcJAysfgXTj6GJyX6M1xkAx2Tj7hCfYwBZHv/
cVfGRPMBE+5JAGu3HXVIYMPkb7+pyaecj/FdxrlF89KXSnJqmwSntgZFHQMsz9OC
XgLXx/A9F9Q96KcPHMzqTOAJ7MKAgAu30ohzdKx9BsKxoklLuxeBemBU1eSxGvhy
rWgrVgKf5et0ZgMv/7SOfsr3LUy1ofusqzVGaO4WithhvB21psXSKeDFTo5SIvfN
I65UHOhfjojqbLtqo6DQILktdV5uFzVhoK0jw3k2mtmWG2xgN/EGP0Gx45ZeH4Rn
wRx3Yz9xFFQ8rh6MPy0X2mxEaflbG+CRmmWoTf+x7UTQSoil7UkCni/t4P9rZ//0
7UFPnbDQ5vyh3Fklte2PmBNuEbOp/8h7uU00bnmETCD2HLlmel1nMMaf5oGCkcr+
EBk/2bd7kK1wliwnNaqhOKjWrHitPZohb6wxbHiU1hTqi5qE4ObH4xeNELX8IM7L
XLxHwrkosuOEATMszDn9AbhxH0k6KNLnGgj++StLP3nOv9e9jTrVt/dQBOCogO4o
AdAZAjfTRlelwJ3ugvgbzYv1D4MMkmmBWB/vMHRBDqayvTmZzMDnlzQqT+BH8ua+
DtRuojlQ19Tusf6pt93rPXKMTb3fCaTmtyjF0Q0aF2MBvOnDwOZn59Y6OhFh22Tl
QyouEYMIulrvHSN6x2FTmKMaVoJigHjdghHZDRRwyoSqBEoGHQCdYn29Q3Q4/oD5
AEfHEu4M5gKpDDceUvWndK4QByZtKj9dxlGwXGPY/RrHkjqomYSaN1xmjmy2MG3k
GihF5lod97Ahxs6aLS14yeQFzZNTbhb/2mbXEwWqowUHaDFjclV2LvVgJe8xO09X
akVZGfGqDADiBLSxx1zt/Hgim3Q6wHHKS1oKIX7DmkFduEIt4MEw4/gK3mppQuox
zocx8aKlQj3os4LaREVs7ZoytWuUtNevNt6xkEWOETSK7jcAUoUkpohr7aB1N5nC
JlJYjId3UmeGO5joUA7IOR2H6JAMrAFTlur0YTxMFweLpWzaRRsEPUow/gLkR2n7
dellouEPd5oOn3kooeTbHqisN/RYFiiVQj7/hnxP6qGWtOWsgSvuoO9PrLALl4V2
tf3VKuAdsIpNQ4PGQo8JlzHB/zk5Gs6GN30+Q5c934sg1oT28SEXUY5ghzMyh3Gt
mOOzRBHGfKyCiNcof5TE5HvXEt5988bkXcC8YXziw7YbNjrEjq3v2cGFkeOJmXmt
0BtRpZcfywQ5R1XHyQI2QLsmAW/AKDxDHksfF13uuprj3fTrXpWHKTo0hdomVplA
OeJBTS6gj9kNGUsE/94EVNooW4mEgAGVdsvm4NP62HiAPEV9Q8CGJAgaI4XGBes0
lU008U5Lcab3Qz41ZuGSTSdsPyN01B6g2HLmDUR1C9LahVsKFXWcIG8sZgiaZ38m
UrwCxe1mEI1eFKdIYhesvFpw6BaoZ/aiOpZG6r1vzCUTaNYU9W8seqpU0qtAYzZE
jwmCOLDbCi67FtVq79yg5bY6H/gKxT2U1BLpDFnFzyEI36xY3cpDPDNOr0VA4bXu
cfdEvNaQrRQkZPckzM94GFrN5GRL1baILDivRrNx1BMMMTJPgqnDhjj0n/Ogg7XN
KBqgEQ2BwfsIpDVb3YBqyea2FI+eSCcrJYlaoyzRODeXtLf22hcnbipL1xQjqrY5
NwTzLxg3MdqwL/WeuWfqBfw1YOYtjmAlLnkwwiozFn9VDEKxsgL5zZqebou8MTka
jO3PdDqzTw8i/Hj5MSi/7KPuik4RAD9nVVhA9UojDzt2pm/SwM4BI3ySlUE7EPn4
0ABiy9IVV88KCBjGfdTvEnasOK0s6dx+p6Lt6uuAr/2WJdVsChf4nC2xgPczK85M
M/6TcPtLARnRS8xdnJH60RokQTzyjRjz2l+A7YLWY1JyPSqy8YtigrkTxsj47A7+
0ToqdCe+VR+FloUzSWhrfLYjNjq5K7tt6+3VrLAKjISg73U0Bf5dZ5f5+QCilej2
svme8BpHvKARq1OKlCmNKIlz3xXG0X1INP+jwiwt7l4P+5dbTmZol86OKeUoTcuv
45pWSp9cVawFDJknCdVKkEpqS7f83laD1jn0dgBXh9Mdz4mmUcFmidLntRNIuQaE
okSWklEztV0A44AAQ0/e7pC5ZJ5bvaBHjGE2SRDEZQCnc1vXWvL39mqG+UXHTlmb
ZizgFUzoGMVmrPj0rwcd3kSxLO61DDapuB8dUidhr/RwKPbU1INwLAHm/AFj4ZIt
Bb9vmgTaCeHa5FhlPnU0DwGD6vyMsSJseZNdWHR2kIEgzLczju277TBu8dc0JGhM
4jfLLhKPEvyoIDwrgNSkDg1EnvhVU1mUrvmmI6gO8T38jxsWV4aiNKXNAFAUfliK
8odDaK7HdAs8pe8/emGzuTGuAJtUXoCwN3rhjKGHpfsLdqvUJysvfFtCKlxLqJCo
20tGTqvjGWwO4klbOCUsr67B221QGzFdyuiFoNBWalBL7xug4qpzwwQeVS4TnnML
hK8BE1j10oOqiDhQkx9Nc52tXg62xK3cHqPmfPJP6jTDDHCIrwsfSSGFbqrsIIxR
7t9nMQk0S1WPP4vF3EBZu/wU7bbsxXmL30aQvzUD+Ioc9rOJRbtwZIUoer6aXjp6
Uw+o2om1hnuHz/iu051jvAqOVV7uwRcfZpKJlwk7Bx4EHe1TjEwOWTRLaGrR3ndx
h9oLzeHT3p/Vbr/ZSyYngQtooH1TXBTHp6Be0l8U0/2eWINK1TXl8fVlnGCN/pRp
QedmbVMtpl+W2fGZADj+6vdCBc5agRFoSKY0k+Lx4Gip4P1IHXp2Aqjph6nmkzVC
lDFIQ8FsOro57eT0DbjqxxCIQ10tVGNjaOWNeLoiqUoe7N6JdRPmzYia6IjLCOi+
G/ei+UeGsS7/UVMcdJBfMlVEgxGBSLlQ+o9vh4ZXuuElsQulCFdr1k1viEl21o5O
Qonb+vlcFrNucj3XqYfWO6Ewr+c3pL24vewGZDWRinzX4zzmbl0qW3bbhtw+jXhX
tjnPObd1HZXCCjZQub4r/gYkbwF5kvCgeXvSBhkPuqujhWy3mIFsLJbY+IFL93xI
FRDmcy/sccmhrbDzBuRKGFEUqKkQF7+19pclvBIGN0Ut+H+8tUtAJeMu6ujVEAkA
eYVTqYCQ9AM/QVNcexy/3+6ueILbIVzAJ572IS0+IeKEsmFpKZF9Fa3y7ePMXRGh
5tHz+REQyD0K4jCh+7gturtsahlvK8sg9Fu9/iBrJtRZSYXop+aTnWmYlrN1DIAO
aFxHLE2pwwnW3fsFLv/f+zCXW61Muvvdc9pW7PoLt8F8dfQeDPm0bg1898V3Ylbm
jx99OiwR6uwoAfmPmNnv2evNp6t9XXoI1HN7T0VqR9u5A8ZdVIq7MsIgCiAbRJ9M
buBaWSvLgyGBynTrfyQnJuZ1/pkFkpFmuD4+4LoatUjoqVj92oSnAHqrm5rPE0d/
82K/lyigJsi/k/eAWZbLSw61Le6veYWx4Iw9UZ5Q/sWxltAQ+ChDCac1mB4ALA8g
x03XetjwyCzbDoggKJPtnIOD4PFneGHVtXqFzAjSLmJlOj9MMUabNbXqMuQ+2LGe
RSzym/G0YsZv02iEbUJ2IKGVsU4xhx5DVXmBgX0vjmtQ2cDcw0vDfXWn5sLxo+wU
puSjzzEQTyYFOBpLop4F7x02DhltKIMy/jZR3ijjDkt/idltVp1Y4QmjaSnnnykV
4+r5jlY4TnPY568voL04rGQfrjynk54YfH1fhoEkMpEAFDT1szdPkvGibXmVi0SX
LFEelcNqPTATeJmfb2O/6xh1HK4MCYj+X7bhNAXaCa/+oLiR6bq7U1XlDN8MIy07
qh55vJE9jApaIh63CZl7wkVr2+fMRL0E8DG7PBinxoBl/OvuikQyf3Msn+BbdI+C
GdRsAfgJmvYHd5Asr8eUZdFvA7XicUboyeSFIBsyGnTtKGAQSyXwhGIInvM6FWm5
25nYZMCgCEGkisccZ4BLEAskiH0jQ/WZxmaM4LiDvGQ2vCIDMSZfp6s/VY5Ghyj5
CntHePipX1meR/TOz2q9Yi+CFYIGrkcvttc/4wjA0AHqdsZBMFQDM3HPxlCncNmV
g8SHHZ2/J6JCVlNMCrNGZIUM3S8Y3BvsIXpQiwQNATTAQvoFQbOw+yMhRTBZ1sx0
UQ5mhViKAeSVNCEV809ZnrcNLv8/yVD7H9y2NBW6RlMVCIRbX5gH8rfXmOTxtI8Y
ingVYLsvQk4nZSL7Z/kClXsdkwLLHTYHqBetcqeqLB3vv802qcLI0EkOQGTSIcBM
myTNBeC+98vSmSMpNfmQQBgIA+1m388tBOOMzXNv9XjUcrKTrMW4ZBD0FPKWoJAw
igN/vVmSeCYXzE8y9eL4z8nfrRphWHcHWwmMiiRh8ItfrxN8OBV+Xv3HKwtC6bHB
LPaYVfK/YLmTjEfF1f19M7/6dWaWbqxy4KPuBeHIctpNXaVTEYNNxaWQYES4Rewb
d60f6cZAtcyOJbEsj1JbGQlkim7W1g+iMiTgCOXTgaSogRjL1hORk3lXJq+oGOqT
MSsL5rJ8JX0AgRWjzec7Fpp8xU7j4MbvfQP86hJk4h9YiNo9pAjp7kGCZFvzZd32
lfWoo3cumzTRO0XrTc2N1ghq5QAoe2xJLyCcFuBJLzjjTPTmcVc7xn2KoiWzo4hI
ViO/JrVHcWoVSjORO1HT1Djjxg6R9HzTqL0LjL4lZ3Y605HKa+RbD2atZyKryhql
rJr1kqF7/OCXHf/N8gMzIWLFcYBjWuc4tBbBklRgeDhN6ikUXci4b4BFPyhrURaI
6Nv9/Dcft/pKNDazFu2KriBbfEdP2muVTkEOY1j8TwwR3D1c7qHs5JFB5rbeI3Dj
CwR6ibE4HXn+dmsST4im/9k7hmDMhHm8xF57UEYyL/tDxgOzhbHGZm8k9ZQQgvw5
ck4jgUdPkNgI16R2PVzEodITTyPJ00IAhRef2j5oe0xGQW29KlpPkjFj33bc4CFx
gAemiDboEY3p+rrNZvRpxIGGuThs/vr6oV3ER/QWbJr0KeO2mSlHR76y3vCu98HO
XiKUEykLJdUdkawln1HXslBzOVEv5fwI2ukWGOYTaX7WeiIVP8h5amueo8WKqkuu
gy3Y3IulsSubU/O4OIbaaMgW49nf1+WaXgQBlC2cGjUEu9X1msu4Emvpel/ccLVm
+k2nfaPqEAw/ZpBkka0MhEg9ggoVj8v6rhi9vy8sDr+ps1XyH5/oiqHSk3l18gTc
gBeCIWQzfIhW9BkmIOJDpfVSXOk700ID0YZap/T1UOTJrSQyUN+Ncqj7trIN3HLi
c80loHKN3S0LGWaAM9PgcFbInsZsSMBjxXnoDHF97XPC/QKyoCfSo7h0xCzyCSHI
oPFZ0fUVUOJfH2O3vGODQ9Z+ctGchTsMoq1Y0QYfnR08x2DAf4w1zLPLG80VPz0h
41K8mamIXR9SjMyVcfrWO+j3aM6DQNR6KocchVlkkFiYioKkBO/wNYhoTbz7ms7L
gSYlPj5ek1j7C5zhreUO7aSXtjA8dUT9R1CxiP17FpS0TSYOtHrharT9CoT3s2cn
6YPZ/8SN/6DvjAD/ib12k7Rzaxin4w6c6D+ViPBYazcT65b3FknJFANYsOnKQeCf
Yh9PJr9EOJJIsdaxGTYoQba/dSr5yMX2sloLI/REfx8q/Z0tasZrpeah9Lr4kipu
TAZVDii+KkRnSMuXrI16qeJSY48sd53wKYlDIUYS/S+xY9ogVCWurAv/lt5T5LUn
xiiBwQCaP5RJ5VxdGlnUq4BRNfydCdqPEL02N3xFodi42qC3FEZVZvl0cQ5v3yKD
VPnr7476KblnK8nuZN8rNHaHDk7bo0Uf4COi9Ic5pOA84aynHqJCEhm1x0kBAcyt
JJ1HULd8RfQ82PCD/geLc+pXRgOhfv7EeiBin/xd/q8RCgHrzjcDI6fHxDHR/+xU
SM8Wr6lBD/GFKGn132NhSzDX60bae4NqVhsc/jVsyj4PvZci5c3uwyq435Q3OpG+
Ogvrtl9yZqYmWAbC8SBkK1rUril9hg8G3qiyzXO0mpXloYOBBdBeZElsvIwj8osL
ZAttHO9j4hGTjXdpNadjZdMVF43RGm90YN+go/Uagy9TExjJQv8yuafo95tB4Qm5
UxJ0/rhozcOxtaLcuEYo2bURBaueKpq1aUg02roEbXq0bI941lwXcoQdmrNhAKno
BtH5J487lftu0iJyuU7rK0YYAJP+NoI0NL13OmuKmaV2hyzj0YCSifXBAry6uBuD
oIj2AyISI03EG4t/lUFkM31iy9azFsUNaK2hZVTKTqtDb3Q0OZkySgA38rJyGKko
l2V4VHnUflxq2bQgzONK+riulhZUN4tPUrRYG9qzR5AoKSGoZqIX0dTxUZufO9Pe
RwplHw8KHPhAwsU6EUVA2fheE+nyxR8VlgnBRIix435XK+RufNsNoQNfMVTa6q6t
vURSGw4KS3CV20zmZQ/N9VTOQgpjFOA88Q3f9hsP4Hmi/z1vuix3ODYZHcf7ohNi
OtfOwCwA7qCqEo4OqjKVK/BEy7ynSV6G4Ql3U+UXL2IXoQUaSJ6r71vafmX5WkB5
pL3Amrjrfw7pNJjcbJ5CKfMq7gtg+iLf7UhnGQ1DA2Z0VzIeXktKhkebXqcc3guV
A19Kq4/YiHWgtU5sNVEB6NSyuZNY/ypgT4Of3Wr4K1sQe1p4PJF5d8Fb1e6Ib9VU
6++WnZ5jvrhbOvBno3/E3376vzaU20mULJVayKuditCpz5gcvgnmpEpZLRpFeHkL
PR8ol6MeDwsK11nDfZtKrzCLe4zqSUfHoTeNsjLw2sFJN1IhIOsFWqqUlrDO0Gm9
PFEvjkI6gZaOenkTlXp8XI8aOZZEi31rnlxbMF2V+0OrFWw76rmljgPpoEv/qCdM
YPA+GtGk8sFyeISCkdbemGSogUWar8mE3tIbLHWKOYNyR/dl/oq57nj6tnxJY+WI
NZr5Kz41Do6SG5JcgfrBuSAn6NDwUMDA9vcKyetR7dxmq2NWPf3BnN859uDXx4eO
leCZNVlEH7xCts4eyWcETCwKeQJKyo44ZexUqjAgHA5PbT4PWwb+QO5b7prS3nUl
2tqICAU2h3kDBHHvCFSmhno6tDZgfx1EllXuGNVs+ujoMnmR3nwTCwOfjMGW7Aso
i1IwMggI872QQmm7OQIPpHb6SqTsCZdZUvt5QnZblfFvEbRvsbZFvWLOHWxvNMd1
7/zDjzSQ78pbFrh+wYgWye6YeWgB1SNaISLO0zJUZOwSx2ixCl4wUNb30CInhES+
69N7IaU3w5xLegvr7K/e5nKwDmvAmMzmgBBnLnkU9CnjsGpHtgYczGvMWXhR5tVi
5gLkbOh0iUPDVWXrHelAzdd+AVuNaKitvYSbdIRZNk7R5lBD/2Nej7Q1WK5l8lVa
77sHI+f5nOwoN8EU9tCt9geD6/hoJ/Xo1XLrUR8nbbGAfptzFExMXuOzHjnhef8J
9VL0nNDDYjPDdDDJis34ZgxIGnCQ0xqtURUCAjYoOyLuH2Fn3QtgoeRsDDBnWcIT
gfPH1Yn70Bis04APqUvOWvrcWTZond7QRzFHeJyG8N2rdvG5GsKGjK78SB5JFW/O
08C5bDft5Piym/ojMnDqBeZGGc4C0jGkoozr5l8QqMxU4n2nLBwwnAWdbCm0f5OL
q8/v/fCImnE8jqAQs9v5MEMggdgm57W+S3UcVsc3jwB/H814CHUWxGwvzkV9nLSe
OmZwtklibnrWTIHJf8DZDL9WvucoBP53m0xbw8Fxd8m/f58eWjWnDBlpLFQrU9Zp
dducNfofwvKhE44kTyZZaYxb5LJC935T1VzdZC9neP1puOXU2uNnwB5EtqLUwzw+
3sYW45RMO5EYlFPmusS+BS9Aa+L8BkytvwoncLlyIUslAOUtgbN9H/fooRx2v3oA
D6Cyrn4VXq+5jQn5u9i5ZK3s67taS1WxH4am0b9PKQfrunGcvNCQBRwShXG92s0J
UbaNTQCXGNTzwTxfVR6eF5dN1AAmyGu2fw/DImUmhsg5lNKA5xv8iAYYW/ACepby
MuL49PQePf3yCqmnJJ5FffH0HdrrdHQztMTLDB+2kS+w4A+XyygZkZVUvJ2rxGuM
UP8B+MkUqn4WE4TYwnbC399nZhF6hlKVCwcGlEsw2ekxyxjPWHfy10baMEbb8/nQ
l5r/1v8qGI5AIpbaiDJwbGlk+oqyfR2I7dHWxoduuRMBT9z7YXZG71zcH+nteTI1
oasHTprcdAXeNaouLfsY2f9/iksfaRybVbUN2pRUSSRSgn6KpbS3vJhRG6EX6Tuc
sZPi2oolkQ6OMRD0GMBzuQDkRn2v64DEZYBYeqotJM1QZ1RgR5ubGeeyz8A6K9hp
MdurrXfwnrD/bAA7un/kiUt+R72NDtS++AIHKp1yoN/yPStm0Fc2Av3KmNXOimuv
uvoywTu+YWen6FsrPVoogznMots9cxvCjzZoTRfrzQLGhfMRc9eRwWjeo4YR1Ybl
hLMc9jGlVVapXUEsWovhmsVSZ1bF4Q+Fc6olQKgKZnJp3Q6sB5Hpyvoq1/YkXm/Q
Ar0aYZxXA3MyK+T2lGOPSlajh6p2k416skrH+pIU4gKi5cGi2HnFTnYx8LKLHzii
vDtdMS1Cr67P83wGEvCPIKeb2lcILjnD1Pr6KtRXeWfqnd8yyVUvGVVcg2IEQ0Rq
uh411rgbl9bxR6nHQVI97yWn8Wy8k9W1nlsMAX+sLQKuw4jAWshLGd32cRSXsi8G
rq4Hoqr+nuE9GhpsQQaQB+Kkh8xP/Lg/ns6yAYYqKxk9y/76Tm5rakNOMytJxEWW
Ybx6QINCNtgpBu97x/heoV7fWWk+odsdPYTv7KWX+iWpuVJrGdJP2nCS3dGvrNbH
nQp4NuYC2j/EbUeV6ZPQ4e13vxJMOiOSiDP1zIv9wTkpQIJj7lijtBcRBNRprkP6
OsGdTg07VkD6TGjzetnF1PlTVauEkZJFHfbVosj8WyyQZvWC44MEpksygVaqp9GE
cDRUZ7NPMYcedG5Bd2CPKsQucTvHHy7WvAl42+05+kgLgBy0X/Qc83A9vk3KamBe
b7idqRN1BSkm0SmZOObjYSTE1+JJ0X44laDmcZ1uJZ4+41lVU4BfJsP/eMHIHyhV
rhT3uiGLfLRpRvd0HmkX7jMKUbm8zvd6bcJcqSakHxBI8BkA1FasG0tb7tQ7prYa
hb+Gf8xW75GbocQATzvJRSQzDNRLtAePDmmbPJrPZX20ZUgl1JdP+c9eFmI2iyoI
FCeK+DqunAgG5+t/2330FybmxiCPaNleKouACVz3o8R6COAZQuD8Zw1b5ILyw/OZ
YEZ+dKzGhNrSpVTzwuqEAEjbA+yJl8dhgiVm7EP+EfoaJdhECt8qvsbHDqmJ3mWF
ybxLGDJYLL4LlKBv9CwqIoVe0J6PHAmzhNIMoZG+4wbJVPhw+QY1A42/2cRlg/hs
hQ4tIWCUmgpTMuIFY94risWuZimXl7K2nTcfyO+8y1n/Y/XAUwo8z9HHik6GyUAe
QlcD9UB4qFBbFQVuidLUTTQA3d4F9hmB5i0qUzXdXO8+KDEVPYEgKqe8RfqbySJm
vMg9Cu1v65Ap5UjprdKS8CFJA6MG1oZ0xYvgYmJVvOZ6rEDXXne6NVByiFLKlj/h
0qa6l8tklSDQ+1gtSaCfJ+YJrGCEiJNZGL/KGDGeAjcZao+CuWjs0Pac6F9DR7mE
RlyuGajNWu0sbXzo2CPCkZNOvTfZ/AkmT/1UDnW3pHuuZeNoR/SIUE3a8+tu6XiR
hidvoE0yTSnyv8jc+BNOEqK+N2psIgkYf4QgUtb5WBd35oCh1MU8lPHKrkvQoilX
7Dq3+sJEAuI/0yELgPUPOycXOPGIy3i9hX8bppitK5Y+CqDnHugpR/IrotVssX7Q
7wN4IFMpCEhyYGwiVNlzKQE0WqIxtdcbQ/TIdzpMSwPVEZXe0HA0oYL88zWUPIlI
FoLOaczur2NUmn3gtjziPIiN8YimGT0RYE3YnSmrqOhRv8YxeCSyJm5zJZNGL0RG
xmL3QoMk0I8BEZHUjy2FaZ9g2waLRA8ttjimPPLIkInTRzlqchS1w3Fi10xNPi4q
sc8YGe6kxD82zMc8OA1Tn4w6hEnyfVK+/yHXb7ZsvM+lFjFLetEmJUznPMAMQ8gG
EGmYYN6CK2N0QS95LgtgqPbJuUo2sxIXApemK3++pKxn49GuCvlZAjmBgUYpuLz7
hcU3Eu34yKsHhKZiKxQJdjKxGlm4151kyAdr9k9SkKkJWmw5J2Pj47sRfHTT09CP
zf1F9tPU2Qi4Gh4wQOkyrfiIxgdXbFesYVB9j/WbyyW5w/jr024JBlO5hMY5drOd
n22B3ZsI+PY74o6ppbpiH8207YS+3Glx0RMAvCjV69ScO7vAH6+JTo7V/w7QZWh5
FDR7roGVCuHZdfHNfJbntIcb6LNsuIf0U6ObZLYsaN5WQCndgU15+j6tVxTa8bKE
GTYHxetbMT8JMylQ6upLfPahY9CZzoHko3q4SVe3ykqCh6WdbQyTvE0QYy9OU9cv
XWrhxSQbpgAzVyA07eEFanM3jzngmaU+lo1FAGZxzrzNqmvJDysPBzGctwqq04H1
rLNUwz4K00hPLllZmFd4iG71mJk3j5pElHlEVo/pW/niYpHt3a5PjnDMZXbr/U/f
9dKpCdvMJouMbtX76qv80VRNMzYwm3D6U2WnVQT3eW1ytZAnwq90Ug314kegBG0E
knijsFZJYyrMN81Kt34mLzE3M8eEBteBbsARw4AMAHl4V0P2r58shCkkoX20X+C3
Ga2vEKA32uCsyytQNYwRvwOOePkWx00TNJnDAsfwUNj6zrUcadIvAscrSmoBGQdb
0oDD9EPVv2WApYzBrBk9UdBjFRALTWJlTxRH8STaWNIAB5KmGDqIezWxq23c6DyB
hSzEXdBVv1NZ9pMmQW4Ct8aoDNPOdaYDN2a0cmKHHJRhcOUMvGZakE5BdutxzOm/
wUm2MWaNV/wYYjFJPAUuVTQyB2y94fZZJ/LZw5c+HaWY9GP89NfwLvE9i9B6Zc0T
Z+bzJ373RYbduq3d/A9UG+R+Qa8XzvqB7ILP0gFsU3sui2OeOjUwxI77TJwxPeMa
DsXR5JP2ZU9Gl37AdpssapZzNjkrXs8DYN8BOcrGwgY8UsrgbtP6jo4f5YAILIJc
S6O87OJsVveF0gTM9lvMH9vaQ3q3WF/Z545UYgsinlf9OUvSxuZuw13roHfnvM8B
NTc0IrvAG8Bhj59dELbcKxiQ2uIxQwQSYjUEQ4Q1PcRDRGc1TJ3AI2K/n+ArWdSL
LUEb8oqPnxKqorJIrRWTqIT0PKXx2ppa4XmYg9uqXq4SGJlWT7x1ufGXL+dIl6kt
sZ2/d+qsHi1BRNet46FoGyM6bwK4E2xHhoIEa+NJs2ybtfzWDfQC2qXtkvpisJ1S
i+lveup/asx9hEMRB/SyfDGbc7tTys2AJqnA5aaND0yulBkTNIu+3jnvCsP2RqsC
LZa+gUrxwLqJ2yLS2Ki4Q3iovdR2NqTZD9jBWDjwi1+aARePnbf7P0FSD1NIESad
fzcwW2vlsZxn5qagjDkUNud/m/ItQkYzEawyP/YV6PYZdUnrymBp2xuGJ36CANx8
fUdBUTngPRQV1ALnwfMj3Egvv0NQhACKkgiwXBGsas6gjrgkbAHyUvXoxTLMPMiG
kHk71g6ALZ4usTjJ789os0VWGudbZ+60kTIOcQ3ow9+I5KoO7I3T9ewCtiZVy99S
VE3NYPNccITroJWZ4bGN82wyf5EDRkaxJZwgCYltuSiz4Bi3I521F6KBTVXNuEoL
UKDOkBqsXEao2wpFVGF2T06Trs7lMefqx1PKFWsuMuisypYi3p7WowHgNzzO79lE
23i5JiICWjSi0lTOgyAlcpqGK9kH2DCozrveah6TXf8O/tMoUHaoPLzCMwdaTFnp
iRb+OjwqAtyohTWop1+p4MT00PSpo47h5Qhl/pwt9lqAbKdhR1HbH1X04zuwSQJQ
M6FlZYPpD8Mdnlj9OD7kYAKSjG7iadoEAO2YJAszg9NLjkVtqZUQDq3EnuhbpKQz
JPBo7NniBn8AJNP7xJ2Cv+PIZy/Q0Ng50b0tlW3N8NP0xvfMAuihjunktD/lxHw4
UMpnPhHyume50a3Jx8k4WUTDZdEmMgrJTWUjERvaiWKiurb3AfRw3SRnUlrGzdgv
ul9yZLMjYxP/xp8D6RX2pDyOZU/VpVNGWScfOzCqqQnaDylFwIUuk8LhFhbe/J/p
0bj7pheWx8rN5F2A7TQ2wV589Wq8au7DL1AM9O8GrvnaTepADIEluJVJQpJhGy1W
spZmql4rrpf1nOPylMqr67s6PsimuFyZafCSZS37nqgUvL9hiiVO34nn2mtHzUF9
CCM7fqyR/caDQVfixPAGmX1+ff0ZU7F8Szhqso0VFXQgejDcWYBQgTTn/i/KwTPn
gSLoLch9IMzmDRZMyyxp8HXEGyrHXRgqHKTWe1cu24g0405spYOI6HNxO0McRnG+
iwSdv/GeYFBgHRgr0b45TNRZF2CGOqxsK1xy+UNXDfQAyr/kOxnPoJTVz8SVa1J6
IvFxNOJPnxK6P9EOB+YCkIOHOrxVIAhrVhp18uCWv6aBXXe5rgj34ie8HvOlilsD
/HaXKgY7Gm9BYNeGxnuty7J795hrfkW17ltAG9KkgvTn0o9frFJNbanfrdrYr1mb
uKEv2CoMF8BurgvkZQmbgvv0pouL/RTd35D4NX8664oEQUgafu1R1lgrw10qJISt
ijV1qiRIeK8q6VdzkYcOnbaMeO1v2rgX+4b5A8ufd/xips/m/F6v1XYVwY/Uxiph
T//j4pj8gHoHOXEiLY92w7eQVtDlGGtAo8kDxrbUx4rlvjJGk6kv/GQa2mDnhE7U
U0v9d/ABQ8J8EtBLG6bdbaqlecV29XDG1KeMkXE1Id7ACZeTQCrHlY5FowdI1hn2
WBf9MQBTzZRA4YnvP1+VyFXhLUgTIs5i22lZCauNBVUJssJBX1vGmC5QpCjPxiS2
U1NJa3FiMXF4brKZ77RnuZWr6A6cWLwim0yoIFQFnWqbD3JaBFKcwyYiZ1MqG4Yf
Y112JYltAwA/BH5+a2J4s6cOL8xbjswkvThGge/28rNPzjA4ABvO1CzuV5aPmPsK
i+klIweBFuOR+sWDXCGzGZ9y5Ywp+Hbor4exLRZcXQB5Kcy09WSESJ+krgXb16Dm
SMv3BuB0MnwJ3mdOHOBfnqb8Z7ntJyQbUr8zCO0C1TKL5nn5zBgwWvpTALwvEemM
PbzQ8LKG2HQBAjqluOd9lCRWrqVXVLa8omEcP0RBbRMGA7Um469bsI5GHiBp+1u5
ObuOvGjGfeBcJQp+AIx+CBVMpEQxLxN9M25PXbm/FTnrXZP2woHFH6eX49XyUAVU
+u7Xvs136g5oxzujO5W+l2/P1N+6djLJ9toG2BVT+dSP+EBLJZ4MMGql1rsYlHcL
xBoBt8DR6emmnMvyTijcbm9r4SVrXDP+i9ZBwt2OIOr1C43us3CCFgwsTwiZgrMm
SKx9lsClyE5+N9xw/mr2i88HJndjzEFKybjmDP5b4JOVDx2TCiDWBUgN0JSTeiR3
AjTSIr1aIZ+6ci05aCvrbxk7BqahL2pfX993iNxuCWO6tA/lpLxn6pJK48H+H6vg
GeCWu1WEDQElAxiO+q9I8fdl1dNMOy3uDphyRtbQ7gvov26b433lO1UPQurz6btj
04Qlkd0jD978SA/5ehVFO1MM69porYIZBriVPJeUEk3H9tZ4kBploElz7MTdDYFU
fvMZc6ZWBeLU87umWvTMTgbZjAXMi1XrLOt3J6EQ+dAz1ZoI6IXZpQcw8SCAX2QA
j0z3KNKrp0GgTBPR20LgDKWPhAAfen6sL09EbM+71yQ9kv7LTph/j5V/mE89KfS2
R2y4qJKZlfHaKDKREW/TERqvyExuaswn7Aica9DbEjdap6BcRXlyN3R/Yec7QytB
sxQvONRZemn+B+jnIi/5tPs3jT0fNFQlxrVJ/OnM+LeKgaGVVIsV8S9LysnmIzGn
lsUu14XH3jDb4F2Q4lMrAH4qmTnHevBytuGmJ5xgTSxPmgOtscJuJzqWgNWFEIFW
fOF9iQKf3KKZGFucGn/w/qUqsm9rG3zTyho3c4x/YH6y+QHc6EqXltlTYgh7Vc5z
FyO1OygMArS0ZLNbyaNzRMus6em9RrFUiOTQj10k4VswWJqaaAati61QrTvwcC22
Q6U698Fm807W37S++lg4qX4AZftV9zj0pooNl9oo4vnrU6YbyV2xqOHPpmSJCwrP
vKxia0jbc+WfsaBd3fXhCaT4jU7bPPwm6UslxFpYUlbV8sWnEi4M1TGulxuQ8/F5
9Hddcev8FlAickzAOQncp1IN5xtlWogJO11D1PcYXfxzlyot7fUAH5hZgDOkvjPE
YbUohjIYcsDawl3oyyEf2lz3Ex5Rc56gQfs1KZn2/rmeP6bw/Z92ubcS1wWUcfXy
N6aNUKkg+Ew2MceWW96t9AITyts17lN4lW0sj0I6XlxEqEHq97QsyK6j2vD9zpwU
if1P890evxsjLNePR369Hk7CNtHivR3RP+UhUc9QpORpOwCcUW7e1CadsmkMkiDj
vCOv4Fe+T0nt9wFf781RuEFWLOp78ZH9n4LpOKndeHm+hKlEAuLyGB6Q/lMA0CVQ
i5VikRpHoQUIwFFrVIDcR0ly5SND+KiADjVFzc2nAWd4eTgHdrH3y0fU9Aqar/I7
IIwqwfRxszmka75xQ9lsujun7E+ltBD1gnv6qqmhKRbfU8QhT2TK1eRlemobBv/v
oew2TJiGsNrJp5BkMVVgQsgU5pFfXf4ZaXoZXakisSea8mv64z3m1lGNYHVw/1e/
pihamM9xoh90ImR7ITTWSU7r26fquVrVrfoohkLXH6BEO3NOe7hKaWv8j+hw1lWc
QPSsCiEqavz8sKvmXOZV7BbjW/Ui4fIPxSv8t09ASC8/E0HLfDxkr9CAOCz6eNWe
XMNut8QtZahtp/eJ/hcVfZebQ/eVDlLEbObLm5m/egflgfIVjsM45atOjw5Mzq92
nKkFjASV46l5/czYD+W0qixuLt/aGwCfPNdEgyBf+oe0KOphGvN87M49k2dUVTqx
5dwYL2blIsI7wiOUxI0PXLqhJ0FvTBn4e/P0jgdUSSrqLTexTz+qFH9KLCUs03le
JBoD+pqtXe/Ts1DntZGd3Qe9Cs70LACLRBcjLEFJcIsXWSH0siVUcXVu3OLLvSfF
MN+hTWDQe+mNVCKdv846Vhu9ChkNq4xagFazoJucHIae53iBzeOQDQ2WMD78Ywu6
gmWIGe8FfIfgUZXb3CP1oAH//nbczv+GQHp4/p9m1GYgIeuTp0oco4sr6m2LVQ8w
6QLKHmdHB3QZ0KyLUGUfV8xkJxq9eJJ30YmbNIou4+j70Wkmca5gFm5gtrmu4PC/
3/qEIcZmp1IMgElU/fasHlgynyf76FvdHq1BwathLEb8tL9UVTeC+imxUcJJNs7Q
DZYnsX9maBME3Ewg0fEefXW+KdTdvTodS/8FvqRvzP0VSWBVi+KfAVVlWJdCPiWk
ouEdpKTD3mpSq/6mw5ufQCdeGdWt9BdtMk0Y4SoOLQT55ukYu737XDXBabweq6/f
F2duDlDjprX0BYWWfesOU4N+ghuRlnZDSK2xq7Hye+ADYKsnrQ4Y6cVE1ttGqEjd
iD9LpYkYwCBMfpLwODm0IZN2zDw6c1Yi3jg3oHgrZhriFCPqSUXjyMZYM8jDp0Th
0ajy7+w+SPo9tcFrcb3cvx9UEb2vOBMcP+J6aQQYxuEy00x4ELqYPOZEeDEUrjP+
IGZxHWzz00DCl0g/cPfEyv/7rcK+A+zvM/OItQ/WrNDyJFtwrCOuu3FDbUn26Rvn
JxN3r9dDgC7aG1I7rbXXjcVG/Q3lgYGMk5gRmpljVCzYC6q1fYtaE85LkcVGkfqd
VBm6LNGnvmLe9oulR2q769zN0lj3zcK7iPAs8AImZ6NGJOMepEW8yGrF4kjET5Xc
YpNmFFt+G2op8AhrJZyy0MG+MFbHPr8CM5ZRnRjuJM2OZvrBzn6fm8701G1WbT8Q
Z8sNX4i/QohK0fLcjO4INuruRmF6Sd3cfw/2ZMMzr/oO3kc0l8/SGB7UcKqSUira
l32JAUwMiR1GuWjgmIQZ5iW+GB7aFofl3r1I6AoZnNkQFX76ZXiVnfOQoAXvoOIX
a0ewFjiIsA9Ye2oDeJQ2jfSES8DeW+WqL/fxeVIGvrqWrom4a0KuSnZ6fjR2SU8l
o2oaen8E5r8CbPcfsBey9nwnJLYI0TGtXmR67GmWr9yDxk5RSSvyjDEIdcLAJeIe
oJpp8xCgZk3uYo+uBMwwQUX3jjHNQ0Sl9osOJmaMaJ1cZxHcZwit6uyFqCsZJJwj
zbWelZK9ohQrPOJZ/NdXeV6KIWqbXaKT72xmpzM/xeJ3Ljkz/dh4vrEiQrcwa2aD
ggjzHdNpWPtIzQE6p+Zcnuu0fSno8rudHcpDXnpG6Ri7kMPgj3heMoga7ufuM55j
kWuD4hsBJGjHcvO4HFuN2sON2IHcu0vwV1+Ve/3weIdA79EXfV0p7V0kFLCuyvAl
t1g+PazuEGyg6UX6QxtLsHbtYmGKihj2MAXIegRm2MeN3v1j6QuQLCPHa3A5c4wC
WMoGlhmFaQfQCCzuRijMsxP6Bzgl6oKa3TcfKO9QyJXA1LCctZaslNAOTqdzPCv2
2ClCQWuok8fXw23Y7ktOFS9IRsMiaBR8JE8wM5bbN2AaYTd+uD4EBuTih5VFXOE3
eyZr2HU8xl0i0tziGgr6DP47iO6SDuCK1DdbY9NQJ8Q9D4aH9wW8MBSv7ghxCNwU
RDWnFALTrmw3mTHPlpIrMCR4p3QIqcEQ/95pqfkFB8UkCmpPfx87YAliB3m5Yab4
bwmsDV7BefL9jk6zrDl37du/v7Yzpj5FEsNM+Y7q/ZaIFUcY659LYu9p4fzf3+Ws
t0zDDEGPpaTaGX7pzLGhbtjr6i8fPVhxNOGiEm2y3eCL8eRYzUgMSFf+fQnVVve3
eVeRhtW/fmNyIafweVEb1mjbbhJ8N/PQsvG7rjzerFuKHx8FHG5G5e4G7WtFBwvv
3+pzPlWMp1ay063Fb7Fno2gkLh0MwMrQNrklGTR0UULaAjBFAvfuf/CU1pTbgg+G
zxrtojhuJWEWPwoqAqlOSznU7HNAxKz1Id3aYEzh2KYXije+oT+jUq7wWgqTAhb2
7VX7FK5NzmkrAwAkQ1JFAA4qQkCVV3jF7kyc9Rx1ZboldZgWtN+IsxDHAnSgKSEV
nxKT7PFqxgHPF/1ZntETCZUpObgUZ4Z+xrwmJKjAjTuMz+/vdogoUPrgkRHCvqTa
s1rINq1iKYkD6BR3vlAyJtPKAgcl1M1ARPLlJ6NDQD6ezPZhPz6ICM7Izy93BQni
RgHVlorM0BtrQ/bs82AFoBhT7Z2yAoPZCt+ixFif/skpWgbJcA4xtoW35Ktj1RZl
OqIZfJVfQRyu5hX4B4Y5uONJE0y5eTLh3INU5qauT+Ktwg5ehlPpZ984nj7VGrp7
sznwDQh7O6Pr+v6oObKlyXr75QqE6C5kJE/mXPCU3pDVM4mL6BAmZLvSPWg0Hr3W
f3xm3IXBS7bpGwS1FsnXYnhONGG9enPB0EtZ8ttLZdjnAf9vWirBHTvIkGpG8nX0
tbwfz9s2WXIlchqBxc0X/ae4GdwrAMnmLQCe70XQjX+EjqRLL+vk99EQHi4U0zqt
GqbT6cxJOLga/1/fCSs8lJCbDRFvDpoH0PTMV/1al5ihdTSoqySqCPEX2umt1qvs
hRE/0cg7bjDgsJk4xkMsYxrdCOhWsagU0t60h9y21Sa4VavLIccs3/zf2fCD1+01
9OxhaH+zBD0cg3sfd1NRQW9MkIpRehYV4ZT6vwccURy3TRxDiOMBKNNIrpF9hcmp
jqF7HR6zK4EFJgpk6aT4zb4n2aZMEcugyPvbgdEYCBrDpQi5MWjfD4pP4LbJVDxR
8yY8GJDDQtl7y3gHZolC5+eXWsxcO9v6TO8W9KTZFm0Qghee5X3bgS8NzITgaYbV
sAv1gjYLBP9IdTrFeEDFG0gjIMbWW91NASmzbKJ5CgrgW/olCH6QkPhY0v3YiCOa
2l4xN3DCF72oDdJTLKVuHAQ5EFzjXJUXV/3e4jVT7S0e1iT/mw5JG5IwJaO6KPjz
SyCEp2SlR0T6/vjLTi6oS51OUR3dvbGfQj7BqC/+58EDbRl5WRZdVknL3//fzKpv
NtUnS4mmbQHSIB/KPSywlZZkjWk1HvOFv28EK5xRh4AwyWlrbGa8uoAIMiLTy3w0
t2R6CfiBp5JIXrAed4RxyPVEjm1shGKPuatsU9XI3cRe2DKiAvc4+d1ftfTaa6Sz
LTNJtcK2T+i1JrBMR9VJwYsJtLGfydZavktrvbg3Szf5Z9AusHdXvIPjfX9H9DJ5
e/zU3Gqj6XAunaRj2to02I0VPaMJlu3Qtwg+8IorUdR6pBDNyIQ6PzBsDkPBS1F/
1NCGo/DfS/TcmVzdn6NPJG1CyHfn8f/K/jN0B+AWKtBI/X5fOhrncjwrJTuTS54x
XMR7FD6Izdodz6kcbG8+4iMtvHS7SR5ZfL/RBLPxBW8TEC4BqMdT1qfzXsgdSsS1
iwoBYARh9s6gs5fHawx7tvpdkijdwSif9fuigkFuD9+mXvZW5jJnpnXF6m9eEjc3
ttPbQxpG1x0nXB+fgZyWvyaWJ8x+WYYpVwmcVox/lOSYxZa3X9CY1zM4YWmDuSFq
Q+m12+XEFYYe0hAl8KC3yOuWWn8cDr1kqf3rvOYQAuVEO8KsVUejTFU6zl4q9O62
hbUMb+w+/WQkHlxQ0c54wTHZh9+QyQUYgVQ3RIEDuOnle9eOmt13uNR659TrBcrP
PsMOB4Fny6uGFRcnOtUiqJu9jPt1m1gq0C9tt2mH32QxYDKc6jR2rXNCi1gc0J1N
txtfh4q0eXZVWWsvg9BNxZrJTyVe2Q14eorMOEsGR+4xFSFkC0KnAbSFFkfxF2TS
hj0o+J+y1APjakjgIBqekxRC9DiTT9xSKjwe1ltd2Jeb1aF9Rswu/MKADbt6gfWQ
UC2DV6UbCENyFRdKvEe48BETZmavP2NqBHJXGRZJ0xeCmSUQen8oSa+S12/Wx6Bn
7/jFvEixiCPfhZs89m+HUffPc7L/JnOXu77lUkLswiNYRzXCb3l7ZSB+587pibqu
T6UWOfE17AMU8fQ33zAMcq2uA+NhvUVNR9QFmkFAApJTY5Ym3x6kNmd98f2MQXw9
4cwSeUdJMSpgyTU6+okjC8yzgdZJJCZ0FzY27P2UVhhksM/0U4I+AjIVwUcOw9Xz
Ct9tQSB0HmloI38P16Fmm0GsTKUcSrkPa/2irU+zJ6WLYTmeroiTcyuYgpui9rNc
tdfh3QQdzRgOjLxNW87zO9gmwxpi7opgXebaq7lTJHCc8MReectnirWyXXP2Fy1s
SbxjUe9QYRbD6MNRakpOG37JLBvVXWAQhu64ktUg3rMcmG9Q0FzkE5kI+rap2CQH
+An/3qhg1/FdSiQ9ROgA8ZKUagD8kdFIFNUn4VcPRbHYUS90QnMeLuOCbxNB07WA
b3hR4shvYNoGaHHpgYOU20G+Ef4RJrO+eBfu6ysjFhyZKytOhz81qGwtphs71Ekg
OiFPh/Y62WHZ8fC0b5ux/3flDn8jtEewzvDMl3DSVLOGKOFLeJWVaDTCgq7flyoO
5aZoLcImuIbNE3lsE3te2yD0/SztXB9p+tfg+2M8PappgL866NcXx9AV7XN84iNh
0QSacLaBEgN9iJpsT0EJX0Yyxb+eMNadl5oUUWYRok69t30AL5LOZXL2bqGLohDj
WeJFBJ13f0e/8DmhkqwQcnLxHZAZjUjhCRDgYje2uLxjLx/07Cf5jb6XiLxS7tfU
VzPFNKig4EIXWqz7w91k88Wy5a6lsQgsOjcEMWIkWLUpPzb4ogmNv4CTLEkrLZ2Z
x0d+riDtRKQhTB2j5WsAYS9kFvn1W1HBrSlrg1XB3Lb3dhKGLIhHF/wMTvl2L806
Hc+SWVa9xtIZLoOiaEge+1W0q52Cw64Glm1qxeq/cOPj588+QAQIycwXGJxmF3ZD
ZdWBaOraf4l47ii6YOQHMwb3daLb6mS2CSYcspbdP4YCtLU7rIn9fUeDG9629rlq
CKCIT39rhInxUuIEMEXTUDpraezPQm+/ofTENYuNkU4l92lp6B2jHlTxvjT91fCG
hyF78I1nPbDlGIcRZc6eCH5eB9va9s2wtopN3SgetLA3ZFsh513v85QSfvZgTA5S
VFlDuiUuzysnLo9qgBEAh2W3sBMbP5xLmNm8vWI96t29RxBdjK8ouoApkJ9ORa9Y
x5M7ZYSvziPFSvqm4MGixxGEWqNgdlq9/8UvYSl7aBizz+H5kcPUXaoRCgPdXrgV
6C5GhagmtsS177icMtVinW5X6QpFLnWx0Y65EjMWb9KQgTn9v0UxUCO7IBx3LmqD
XH9ezW6NyIC50d/7pV5pejR9ZSzphf32ryEE+S8eUU4rujeyLvVEE1xJ2W4sYgy+
QZtqfwr2HtuClm8NHaYNynkI3IPd8rN1j+rlj82pM4jaNc9Kg5hUyEKsfB+eTrIU
vQsIG/LI61WuzGA8k2tNHsKdr141opTYyfFbXrmwolFrNhKwPMiK9/9ckutM7Iyb
CF+Px8awX8xyEWfTeAeULKYBZlMFAHngqupvIXQoNn3zrRPPyPl0jvGQy0k5MpB8
xaZiar200OWaZMwWXaq7HRtTBnNHpTYfDjK+EOwemrpDo0YIJ3eChUtVHX0djAS7
c8UEsJY+106O20pNvimyjfSr4JQChkpt1wbxl/AJwUn69bIKH9ZRrp4rN/SlKSRM
RFW5bNCFHPqHZcYelWA/3N5qkyr8QPN6CRx95JTKTS+Ys7EN17cCjSzLJIBpug3j
MfuZP0Aa4B7qzYJ3PSkcG8QA/KJXPhep9ZaAgon2F+uEoYhDcq3yswVDApuDxl4A
PqnRJqlZrEg8alvPvDSYTzefosIW9tRPNiO8DRPsYDuAQcah0jo1PWDj6tn15T9Q
KT9HPyK2RStI0+9gq99Fhkn1JFlNphVOJg6e/TiogVZLXiRXvIXZq9mw10Xp+V1t
bOfHHjvFboqT+VzP91KiuibeRPkBWG9+ZZXSHIQHqfpMrqWrkTLE8pzpjE8+lDwS
GdC8MViYXZWSwZiDt31iL/dZVBQj37cVzWqSc4zrW4Qfk4taFN+77tAUYP8XX6N7
YcpoD7eItNQhDWXvxdUhKRy4BH5TazYX3mBppYTExBlpRnxSqlmbTvH2NOw1GFdJ
k975Q6xmDfbf8VXXJQGg++ZMK4mxb5r9e6v78UpWCw/et2I8vP3RRu3VI6jw2xLF
hP1TODEL5acGMeNWxLgG/KMi5v6RspSPZo7ZPpiwXOL79MxPNjR970t66FGVGnwv
PNYkhLtUiQr9IwdCCgtiRb7gEg0KIKcYKpOWGReNaPWymVO/nzru2XcSUBVxZSKN
wuhatIszxePwu0dRH4VdoLSGgaK731aesqtFz8I7lG4SE8Wv/pWGOYXB90HAtJBW
h47sFsvae75vp2iEQKoDihUNaap0BBPfGCWGWxQrbi6qcWcGVl2GTFSz2wmsOkfU
/pkH9/igtqjNELeWoF+QOxGJj+Y2MB+lskfy3QKIY9meDQ45KwHapi9sQK+t3lGs
BgINJ9lsXZMT5lgI37OuAbcZ1BMuH07uBi0lmanIl6VYtTNpNQ16709xX251g8ez
D2XDzgQuQpexgWuCAvlHsmkDRdLFNA60ViTyygEFR8Fo4/kXmZXXSXst0VVd56XU
LppNBQl6ueVB55ioAEsbxRYgDRVK8V+vnuBYAllJXzcGzPf0fd64djUuRIGEviY7
fm1+uzse85EPM1+K64czN72dJEX1upOblSym8iGDW/DXYRdr2FcOQZPiY1oub1Kv
v6ZinuBrfEhBPvaNcp/+GtVoOAx5xXfTLRb7IOpjzfOj3IXramo5s56J5hFkx97z
nYylbvVJhUzEunZMshmpiQsPMkzPqVghilKbKytC0CgYeK1QeMUuywbck7yKlCFl
jZqMufY5OOSvBkL4Y+IRuswoqoUqO6v2c0fFQOHJZFIED8+7hvKBVuqSaS12R1WO
86CdHXK5l+v0XD1iDdJlIKMKYDYY6O2v97LTH3akZE9AhNE3KQxcWoRTnPZ2Cg91
sR3u7yoT7sltu8EhcTRnnDlBOyNE9zjCFwAZ90jbUrHR4omSgRR3w+qHsJCGRVrm
fgP+sN9EZaB9E3c0afd8A5tTzK4C5O5qb+ZWRx/LLp2z5e3MskbNPShLEUaLnF8G
mysxuRhhjWMCkSfqyyOB9HZEEdhW8oNGlc4H5kSg1GUDr4TsEdIcjLp5+ErHFiFT
Xh2qy4qDoZnTPFe9QXL0xJkeoabcIPFF6IFlzYFr/OVnvgHlDJZaTIZvQ2RznHYh
tsyetAeuXbIcg4w8uNpYkYPLCRAWZj7bjoSuX4yJRGkyxxPbfOHUXopie34pkCDm
YR+IF/xNWGf5PnuNBHnq3IZFvBMNy6AdLYrNNbFiSqqM2H3JY3jcYY8aVkmWCDWV
lv7ndrOwVnmWfZQBNML6cH3qRWrWU+t+DvkOsfuXAv01clpBRV7jupI4cu/UVNJ1
lIyOKgV1K4txsOxgA1ivwao1P394FZhEokfiOlno7uGflAhVklD5iRwxuKvS3Gel
rpDmjqYsPzQqxl/PqNg6BmbVwh88o6fMXQ2fpzBqDl+Cp+J2WPxL4t/o6fpM2kEE
uEui8JSyl0gb+wzU/IS4+PFnSD1bOiaRAMCWsQ3r/9a6uP6poq2ihC5OBUmVmXbY
yCGmC+hds+8EPstJ2vH1CO1M6ZlgODgdJkxyp/EfloKUDocJ55LCwx+fWJUOgnnJ
0heOkE6bhI/7wnct+Uw1h7ZRtq5AJgae1VVqJJvDFuTN3j+uKiM9ANQBXGwyy784
n3ZjxyenGHz2s9GEEx75VKivfV6Cdz2mgEP+qa/6IC0Tc7fcNgnNg4TmqYqfVyxJ
LlwdtGsnBRUd0mdBhdA0OdkRnLIsQGun3567WXD0Svn8gqbHxZso5JUVfqMuaxRS
pGJM4V3QgPJWRZx+VA1ZkfLdtNjz6qDrTywKrqWZMKYAW84ZyKXgi1gaEPUeKSL/
5BmjDr4Vo/Dld8PES8dxIgJ69YKLC6kFQrs8EAzzkeC1PQPB9fEC2Gbs3h7S7w60
ajGnIM4PFYlj3/TOQhU+G/V1F4dVoIfuf2CHdAWBY1qfBJPMKGIm65vagbAVQC+E
/GrabRyK41p8/MywWoe4XyqBG4IXmUKnrLdPu4IGq3/qZtvGGdBfAXXPKUhxn5iP
YgzeF0i4xXN4fa/wqpjAPRogkN3GVV6vDhbnleJuOqdKWwGLXn0gKFiRhGpC7Mp+
2YzXMnjF+NFeoieWeZ5nTXIqsLlwlBN3Jpb/PUqV0yMI5vV/hCXpjoCAfBmLbrDz
py78wzHZ53D4L5pDoaD1MEpYe10/TWrMmgkkg6iQ0NPIdid3bxZYfSz6qS50KnjD
SW/snx05eYt0qGhrkploMHsmPJjGCDFJ4x3p587vuE4AT100Y9COZVag/k29qNz2
qvH3oQo5EeGDZD/5eipn9bMWKVjmglebc6Ty7ugzM67ylqA4laeyyWfIcWcLDAL7
HRYZFCzEYIv49SxQ5tVJW0JtSql8REnmfAIT8rQ+fE9QTz+SLE491hiM6KH7GrYl
CWbU7PpG4Ec01LU01ttKVAEMTesYMOEi9Q0EJc48Ra81WUqOfIcWXNmS5UjsQwUz
0pDfrhFaVZlKaDCIdRhBNO5arMA/6OouhG1GZ9sSLnKDVguHFmYGfCJGVh/0iLEK
JgAIjhKKyByWFBGszfUoMZWwPIPACbJUn2CPjVSX1z+n/PYEXjv5T0IRgPYZbYW8
BfV9XcRcdMsARLEwmpbdeImCFaW/BUSiTiyBkMSNyGMIwW1QIttxB4VOlVyng067
gmGYRoF3eBgvT4Bu/bHc8nIOHh1b2A74dgDhgCENZ0NgCoRF6c9AgwqsMfnPyoFK
8buFCD9gXm9N8mg73bujvkaFgXerPnY/YrBx+5k564kZy4H+SKFx4jfdb0/tXD5e
mg9l4zbEwo4/MyAk06eGtWTYnjGQK1zIk+PGNaN2ar+LdSTfomv/On9QrsFl+z8y
GE4IhqWDOV5WY27stf9P6vJFa9H2yLXRDlG54P3bLObwtFdyFRlZQZXPQXrSTanf
F0dP0Ji9lCCZYiTXXSO2ZsB2/peOwxFvBXNVj7EWPpHK0NuaVIj96QVU+gxQN4fV
lgZLGfTEbQ0ozrR5v0h31YLXhp5+YN0A0KXlUTnoQ34q56IISaCAsoGY/r954NZl
WwniFFGqjbHL4QCAXmyXlkttm7mI+Pok3XXpqO1LbBN1OZS+7TDTEIpFjnLvkAb9
hAx6Vs5Z2dw6jX0Gzf4Z/pI4iR96ApK5mrQQq1dsVV/2rQP8QxWgpwIyQMmAO7nV
uyXiz2oBe5lOXSK+0S1+07vWOAwMOB2mlOCtWHM/tHT9uT9qf34Ro6wJEc81XR2P
z/I951hvymi2i64059ET/6D5ioh1booG/Czi9beKdoAB66kQLOXYiI5K5TqoSucm
Qd+2PNMRPy39wyBW1Nqd98dtc6qI2EDp84ZQMeeogXOjeBRmJaF6kE0ML07rIKzq
K6kf4DRrrUTD0rhSet9EiydVyfElGM6znIGwnYsjzeUj+vEztYJJ3K8BDfwxOuGM
uabQBGk2ubzCta5vsJlwbv9H/Xyzz55rirvU9K4B9hUDztLJWmZpOLEKHCwzDliA
DAXqh+KAM3WADdVSnW5guyopyLAeWMRvVU1GAtrOVfx6Sa+qcp1RUI5WCOeeDeMH
OZuRSW88gb2rUXvdWLnQGEKqGlM3gbLGe5Hh7Zqdzw834y7eVuilt9Umjl1zH0VT
m4z1HrOIJ2D4wTu3Ztm63iap+lf8Wzr+IKTnOBcqOmUIUMzRvj3JOGgn3IBsTrpN
C+DxYyYBUj4hj0Y5mhJcWrcrAk7rCypjyaFjFbec+n6eU87OItYk2oy3KnlL8tfR
wRfdmguhtIZ2IhdUvXUUPTqTcGLDF38zj7npx3VBPrWfb6YRdi+BGWYcxRTM7Bbn
Fl2VHC56zFJMDHDhjjVqeDf1AUGG20k+rA9wGTphpcK+w0QJoVkP/JSz1ImTRma3
Nqx1Zlh7CMldXRtwyO4i8zdkrcKFFF1SgRj/Cysml6pNdVzJUVCXjrVGY1S0AxFc
933BICtT5qLBR+YVpF4j4t/Cr0EHBZ+y49cgypcIZ+QLaAWKPia3EAkwRvIL3IoO
H+UXuEEsImYMbAtyNJUgDqwFkVomPri27Kc8NBDPQCQXEF+tWgmnCokT2lI04sFh
30EDZR8i6d97B9OdPXdVKcG+Va5GsVXrgob+sZo9zjpE6e1PKmIL56ywatCr6hvK
SGYOeVvUUZdyzoqXDn4mE/4JKPbiNSyKYcjW4S82AAM6Us4fKy8Q4fMjQsBm5yM0
tf4NKvQjfN1Ki6YirrWqXLCsLw0QeO60/yx7FEIFMV+CIOU/AY3ziAogVAPi+/o/
JEsU9Q+rgKYPCcIUQHdqOV+mbk39YLPw9axVTNBM/1dOavCP1XSNld0kq2/U4YAM
HoZSjHKyHAJINDNBK5LGxRF1/AQGimrS3CZqqylLwwH0cfoMsq0JBLYSKedowl4i
aClfS4YyPzRVydHWeqjyS61RE5jfOJ2z+5YauhAx5XLdtOfr5YDUETREkGijqGG4
ASh5nOUyopiScWs8065Vl6VHZIVtD1W/UVD0PdthDb2AJdvO2BJnaaYe6cF3e9Nk
isAXUule0x/7iLx8rDIvhDVNertoC+tTCwEBbNjbGcfw7NXRSzKHDwjQIf4EOQDm
1Uc+BojjiGZXir4B2wKpGsNEsVURAsLEFBVeFkeU6KgKruoWNNL2yeFpnavG7jRJ
bj5c8rdVJlTqHTGgzCjpASq9KWYq4UH1Q5RoVKzqC3g1tzLo/B34mAk5IF1KTOsd
FN7ar4ClrkLpocqHEFzufEpQ/NkNjCM/WrFzG88j3UfZUCr4bGsT46MV5jRefKLH
t7GtxYISqpUjJG2EsoYHOfJpFxPvQhZcq1xEsx2PhACtxa6hfDA8PLvWOI8wxzLz
k9X8f0VaSgD+nlM/BxjlJ7emw4Zt8E80ps1eseoPCEdOch2+bXrUkzkzx3+4JRwR
B5qKSLXkqbkID5UT88BPDT1fVOG+4U9yDuOK6s1qJoizEaqb4/SzxxTSe8tOOM8F
5x/D3r+k+/qYLQeKZf3PiVUD52l9zXhxg5dqJ5zuoHdt548GJwZgWFewwOtv7pi0
B+NEspskoeeI7oiSxHuGQw6jVqbhEhQthGu49Ruk4cpkPdzh+KbW6XuOh7mAKN29
9R33fHBc+YeaIPgtQ8dGglPTLdxGKQh/42RPyuDjTlPpmvk+x1EzRqqcQuexDlys
0ct+4iX+RuR7Ha1SXeu3ajnraQmbPoftG5YVrjYhBl4uCiPgiToU9rZFUjmoc7tW
nD9voK+HFHdBgUpW2ln92pm1sHMm9xMprlYLGsgd5oyYxjWe7+7kqE7x89QseOyP
Ltz1b1gc4yHoaeu8vbebMEKipRz86eSkqdnuw2sKx1lV5Ilm9i95CGoQg8rlmPcG
j7pux9gYCZOW1q7Gf24gOyqfnLXJSIpQQcr2BzpiPtWe7pCpYR2VgJvOUvBbnDcJ
G6+LpN8//oYSP3Lgyq1QZlj0zyAqIA79TAGzCvqxNeF/oOYgDikviuEmjR3CPqEQ
8WWDnNFoohcloVHNZX31Hdn1c1GPmh6xfhDpg8CLOGMtfizGcwwlOW6qcVC4R1OJ
6qTHcsHL+q3bkruhj69lJfdBKltT7I4puFCSfxl3Z3yUzTk1aIoI0/9oeW3cypio
rbd4CCqxznLkcS+tAOBouIo1OhgAx84Pc3jfKObNxn0/9aLJoQY7+jbfu7YhYx4j
UpY1OHINB404u/tbp0ciUFYYv1FGr/Pf0bWtjNWt5p7WbBF3J9JxYWWwqB1ak4zt
juxw6GKRpdE6WN930q+RilTeNkqvsK7Hs5xi8WRlFGf4lWqbJ2GSXqO4PHVlzi/Q
dfPicpYdKlasDjnK4xH/CEfUfOsnY0qGCwaEkojV3gOYxZH9rp1Q0ouOXWvDoEe5
00QG2CXwcegK4BIHSR7hAwnMiSy+QsgXXuvFahfQEQOTDUqNpypoPG8fDhV7ndW/
uTdvVVyhAYmSLCt0gsrQLkSY8DCH9BuiLvM5oyEzlFOWR3/kVmaGUsu9JEmo5R68
/XVo/PTOjB+KRYPDo1xEB+QqQjvRiorhhKPTopiGeJx88iqfaqa6N3v5c3pJrbSe
N2SVqnRWMFhmCoviXHbTbr0zPtubXcb4JOIPxEqqxf6GO1Q2XjVu1KRpYmiQw6+F
POy+hydrjNRIQSf+JK80GiBDG3TbiOY4+m5u/oN5fZ3/XcpjegcRf5xlqHTZ1Wvz
RVfcG4UQ10oSvdp/XJ0FXAt6gvfb/CmAtjNzGFyBPnACjJTcsGhTHB2A8/eFTE7m
bIF87Lcy5sbcQO5bQC6fhkEMyqRq9B5J7h5WfiC97h9f6wws0ckU0LnbnThqSkVH
Q91U+jAzKCF0p+pvp+yZFxljE7Ccc9CVYCu/7nRev+iIAAB+iUVWk9VAcg33VMsg
KSh+Y86hrB8XnqqNtoi00/XIcJYAcpKQjeHvgKfYr9AGSnzAGGVKlzI+XBnmxjUK
6dO6VZ2erixgCs4H3QQi6i95/0FpMcs7x3BWFwfl678FEB+W5dVNIwNKNlVAlAc+
gtMF5UiKNhzra1EC0j+JJq9h/TmSSihheR1akPMluqu0ICnN7Vf5lgkwQE7wSAg/
5/MTY7cS7v1ik62zzzft5p38kCrW7ttR/tpOzghb8LjHcjuQ20pHiLxfxmZE6zbS
PgRxhteyRlTYdc+syE+Zc4u6rpdAgQtrERTTJQK9J9K3BmZDNlwCk+6i4IP3BLND
bTCuAVSmXw9dJQhF6OTt8sEj/k4SUdreWm8ZbLuotnV5TS2Ac3go5yEgX4VfCPZ2
1JIXFBHf32maxmRO137VXzB/SukDZctXoouMQFExpABYLm2J4p5Hq5QQ/7m5BOrh
FZI4PT1HSD1olPZcDaibKioOwladw+O71O5YGKgizq5ax+IrKrgTg1aGXxIFd6Ku
n+bMBp4Rnf87+0dAiaeufugZcNOCSPnQGmJIVDvW2ig/y+PS6qu7N2A7OlpumKc1
eyGod73tPucDBlwBawtMaqHYF8K/icA79faGSSW8BoOBK5ZcewL2tPiRsZ0eZRIq
1d0dWto+8djbtW871hjCPdGHyabIqlTol0PGByizPKaopRdBZZDi7cHM18s3jN7k
ODMFu2aQVuub2+B5zRU8Al2cTrVI2shNThk1HEBrPzi8F0Ivum0DkKiUg8Oemv51
ai6FM9O0A4GzgyyoV4ySlB8+IbtJUN/CD4RghhBMF3S0qa5t2rHdo6bjtN+vA45R
mZyknF/puLjWX2LnCLbqWM6fhmOvZaIUpH+XoiJIR7rzsIERj/gL07C5htnYmzWj
bTrhYsRDiKU/uhl79Ydea8W/EO37FPOh7RYfSLy3nJr4PIdfmiKhXvgNOKw5iClu
29AYm0Sm6oDSwzV2/arVWgt8PEvExwCIiMbELyG/kXt0ibiiuaKtng9HM3q3ZoLx
ujQnTthsGngY9wxgvBjeszkkcp5G3lN8B0XDOJJ1D+C6VLg7ZeHsWK6dhpE0Vsrz
lj/cYcrQN6zNV54G9BBEt4Mc+7OHIiKmKZGA9fzgPvQdgNX8lcZDAJQnPmS8aPDg
Z2NJtmkiynqX0mVH3ycV+Aur0hrCXZeHQOphkd6sogu50HuD+PyZvng6enfdqv71
9oPkW/8lpnf4gjDjXNFedMfaR8ZsbkoLxDEOEA+EKIyy4KfnQXw4G41s/FWFBj8C
HCrfnCClt9tuWKYCCo1D18PSGLBJaCWK6eR8TuUPaiUWd61huOFfB6+X/DC2eq8X
jBKIcOh1i1B3ctnPtFnyET0lJui8UrDbv1KgDi2MTdaUIADPp35uGiFD9lvUu2Zl
olbPCAH02ysUbjlL/5GzJgBRcbo1HUfgHkc3IV0iK5qyx308NqDgnF2qQ+31qDoH
eXkpfUk9Mi++GQBojdZQLEd3hsVp+rrTVZpx3dAXa1kCee5L6ZjHxEubXRDR0Bth
R1fM81CkxdBmzb8gTRKejtvXkQEApoSLxqQAISFFkLHp3At7W16AGB7w8YTzMgWc
3y9TCUCz9TpC7Wv0oBoZW6GWIwTWoe3DK9cDM2bmkICgaoG4DMwMqnsV2mZfDKvU
4JheyHUvAeEt+kDv3FnwjaNEUo5V7+A4ra1XHmmmlP7gzex+F5Ik6uwVFb7dsq2S
Um1+ozNg69Ba7/0rk0BAsEpz5Y4U9XJPLb20VPHKWk4+TJxZEHVU9vA91ZHYua1o
2DxZhZrPC3TJ7q7R/TqzjZZmxXUKmyhChmL76iuLRlBCb1dLbXQxLuiwpLBVvr4S
GJdKjbJKVHAQEuGNguUJo51pm85YXSxU8YnN7PuFqCPJzdXwzVUEfQFAEajL9dA+
3eKona77CXw8zbpReckeITHjbRJr6q+QPcIAA+GAPKAoyZ2uOH4KD50qYhhNeXoH
R3zfArhEAHDicKhfOWuA7oLNGHvfJHOgihM6Nt+uu3K9kTDAS+UyWqlP+BeqPwWd
bi9R0Cm5BH2yJ3zYCRmTy2jRRYYgvEmQMpEykXFx+VpDZJIyWKmBz22be7xGqeAY
u5J7FwOQ2hH5Nkb1VT43lcH98z68MfQGm3qwFY7q3yrTWkkU3Vhhddo+WoTt373E
0W5OvuzmQhOo4+uQKsTuzWb+D9zmc5bjtX5YJBqEfrrJdnCJZ2gTgkkuacYuLOKv
JYrZ+j9mSntNzPEn/OFRLaa4MK+Y4arb64UJqkGY8iLf9vZnJHO9EKI22QumXz/D
NOHScA8iTmFCZuGkXJHo7GhaDAodxNIL+UyBXd5p7kbQZxMAk8eKjzAH3natAinV
/vcU4vrEQI1yFseT1MgwQDMTgs81CE0cuonOz62mMcxBVSeVXI6+OStID7oYzf4S
Xj8oq1FyWO0Z2lpgGAwxiOCV6x64aZWVe1lRTAvsSYoId7BIFP5WDOnCFEInQBKI
2yHCtL0igX8C/gCaNtF7Oso9DPjlvf06y9kUynV7b/Wh408pgqoqgj9/XOW3VpzM
h0pEnxn+ujUDBb07rnTFInsJuO18q07E/7CpZYWm8mSem/g5Zu59/rCz2sXLcmhU
DxARMorgpwiG5zIFr/+ML1J8X60Q9fhtPblPIUD29QPfv8+s/QrW9LBriHTlDs46
ey1WirvZm3C7yBLdppBCieKtPUl+LPcrKPh+nPh2Hl0qmDIEV+2lSBVek3QQOQtb
mqr6imYcA2wZZswmsqRRemUGphvGK9vkMc3+Ul13lgtclERhMbxFV7X6E91/K5I8
uFDJhjeKOIGajpl8DdoiY1P72mli40bGcWbykdqPp3hArCknbxYFn40JJxUbEt9o
e7molYYKZm8FmMKhBAcRKxEFCodQYYB3Je9dceAfF6KLu3GxUCy/yw4dctkkkOeb
BJEFVyC8xAE+PIZhWbeaiTO4bHUkg/XCCXefu0U8A/ePFMilkNTF4EdNpcEUKDlb
nbPCAFP2pNM5viePSibmLqJAeIIWWZQ64FE9r9NBub64o5wpeBMzAct5WRw1i2MS
eKEsJ+boV+2XEKNhSWqAGNa6efybQDje3m/noLZVE6/pbMVCrlJ+6hr39IQiWHzc
sFqWST6xY4jI9JihSU5g+vrKJ190Eq+6IJmCY4RQ10sRxYKiL4YI3yDKgSl/PVu9
D+OnGqC7StM0ZSivbNokURPeglkPz4luW/eXLMnXRIVgPqZNheL7CVgWdFpVOK10
uFnGjCKRx7eLuW9omaNG+KO7ikYeSspwHushDGpuVaqnifIAUowD2VnFmN08F7cM
MOuZ5vO6GcqbZA4ulgeE8r5X8HiZ9l5Xwg1ARKJdhEIoAstGfEbxLBbZ2Y+Ikvhb
lv+CsZKHkj52wpuFxGhGtv64hVv9/HiwtWW9rQseAdrBqcEIKfp9gtXbi63z+7AO
XHJWVZX9z4ZlYkh3APLaeOiTZt/VhjR+chosNd7DI6XCwWIkn2klWj98PH0WfKGU
irw+x+btAOFHtYtUYrwGMiXjrS7cxG5wBmNvhxEujgM1boMx5pSem5LKZtmKtHnp
pUlVVHZHSNAf3ajVNPHZnY9WF2nl++XZKDoQ+Z7/uNBq4CQe4m3G44W0zZBeuiNj
fVpIE8F6f6IQ6iddf/Fb6iR9OAsM8hN57Qe5JwJeTVFCzPCONNkUMxCjZMN6Y3O4
dz7H0fo6oEK1EOGyGM/ICFcnlT8aJlh6VIviC29JXxIjaUj1cD3UjZ8SzKUHKuY3
KV8CQzplMSY8HhDXmAprBc4t/Q+fCQnRcpudeTIMfmwTVyyZ0VjXqvHx+VNNpnto
JUXR05t0sq49w6kOggwJ7EaTeWpozj7Wma9zh0JSn3wzRzjVPOLCyiL+LKDP1jzt
awVT+8giwt0O7MzF+OpTPJ8RgBir6fOO1ivpTfTy+AmL0EFaOZr0Cggidwrsylm6
wQR42vNE6WpORuTgEFvejA+1HcoWdeiithW3RGwyZQBZr1ro13KB4Pp6PjdLYpVO
S7EDnX8KLjaDkrKzTV5y3MhE0aS/xyUl3ttOv46HA3x/pAJN5Bu94nu/bJXTDNyX
31rZBmtsBDYak+m7nGCUAnvIw0qn7TD0a5D65NVYu/PHeQpHBzFAPWaMqrCSK5Uo
gmnWC5KqmrSNIiIxOFASHLt+mnso75wTSomaebs72jb/6CKFqyybrfxhDwUFRLIb
FTWRdzv/d7gNvS2rHJlVwwZ9TkS1vtWvBqM6wXxyHC6+lsk/UVWHCy8CJK0IKgh+
Ujt4FGpsJ22jAjIhTy8kiodUK/38Kkmv67H9N9GZ40Kh+G6m8saaP3H9WA1S0I61
7THi333ZiS1PYPYJiBrYQ53CQhYadRHZhnY4cbLitDTarM6urh9AtMcN5xavF7j0
BpqsMiB5W9Lhh6d7q0W7yinvb7wF292V3uDKvTZsG7t2yx7JduGkLsTnk4KLAZSq
3KCCGeb+yXc5TaDtGjoDy1VMZqkFvuW5qVqqUiQJW3t/Or22z/HXAktPypVkjzx+
cDqwfkgNGAaLWkyBIKi5gUHn2Yk4CBwcHGoG0IwGEwhcL0LO4/KNKjVfklxOuRWF
0htHjfPTTEXbRkOdRhuCDuU8IAlIHpJMbonmR3hVt6ahgXPJHrqCkNf6iD3hC0dE
jvyflWMvWfTCYbjBAHfSHzJbIodDkybqduiU3aqXpwWKRAN+GKc4wZD+u3YoDwQD
Rau31KCsnVRU99uKzZVv+Xs9d0hT3JaMTCaKQX6GJdvxPYY5av9I/4ZdDqtJZ5c9
IjUIjd6Z3uziSWQd1rwu9lFfXRexz6S4vkrbX7+ih7JjQfQnzDCQ0SCQELdr5sKb
dYfRyGaJOc+syotZMTmliEk2ms7kqDtYgrPxmTiA2vMJRo//sXsKdxHo6B4DuV3N
Tclj3ZfW3KlAwefmjFqPJAsDtSkDLMgnebgzj3JOdEGdv57b4UOqEROounGxdeG6
OVDuZnsVftmecxT4R/OE8uizLvJWo0/zQ+3ahNrzkgeREwZDJHdDnk8FPMkdRoQ4
RX6WEMc84l4mYDOHRfFI3Gi0uDJlS0bSlnY/jOspwekvG7drDOGCbBA74720Nlpj
4GX+/ooe/Yd1QI9zPVWhw1D3JDMPA5i2olDZkOlqK/2VjWu2jTdT6g1gINN/PmM1
kvduk+h5j76Hb8qZK2mh66tdw+HQTa3+bL4TqLmpr0W58iZoAjt9YMaNi5g1F0jt
dVjmpV/pjOxci4FYMaxs4rtBwCI8WrQ2moyqJETD9AboPwqCwm3Khjs6bhcdL90f
ZBrdj01tRNRH7Rdm6oOOz9SJvvuzuv5Wf7mnxCLpGhdOSXAhfWmRN7Q0+Mlq+kvz
LCaHYp6SvByEyqFmTm2eBhZicD3CbDoR+qV/rMgcCavIoIwjTmOtqf4cT4zhPs8e
GlC8razk0rQwIBOaHMIh7fKQyco2NPL7fB1LhjS4kWrlrPqHveoDA3Zvvd4ZuvyO
Au9mKntQH3QmM6etdHxwg8GAgOu0BV4QEROwx8MtJMW04m0+jUXw4kbJqm35O0X9
yZEmcvsKaZxGi7EgMlJt9cWQV+4aL04RcGT/lFUoFlMwocbYcKkJN6D/8Lk3a2Ik
p+jIzZYaR6REv/pM3E9Rcu+rowSiGKCOXR9mNiq22pabBrTPEe18DlgctOt+4aPZ
9KyxwITAW/Y9HuGFJej+NyPlI/rInuzOAYC8t0Q0YiSdK3v4w+UDs4Ent4rr2+Sf
CS517Fo4Gl4vaZF1DJ97tnUkU4rl2o6C/PmAMcYadEiFvj0sMuyX6gd3vRBe5WYC
Yf1YhzMsT7dO32+6u/6CvsCGfL53PpxElP4OPJiHev88BeWHwQhMjZL8nmOC0o/f
DuoA8Qb/lW/Hl4XheZkFhuAZN2qY+f5Pi9zc3eyKBLxu8vptBTCAsVexuMumUhkO
XGyVYqCkgmQwZa/NTNNMNY8tNmcime1xEamVizegxH9i2tAY4aTZMRotIczIgoJ1
y7u6LZlPw8ACaaNKV0Z1W/kVen46JOFuM4d0dqhQ2MlOtUwZc6QDbE4e1IJ9kIvz
sAm6WEaNj4MXL0jAcCJIaIT1sLKFUkSC0K8LZP1z6ZUi7Mu6rRkXhDrAr2xhdylT
bRIvdflo82hbMJGdkOUT6CgXZfYRERpKWCIBLtfwF6PVSIvRhtGW4CiZD9mx4aQi
NHsE2iat9Zx5Ip+bEVIR5q1KzCsKiuA/4sEduOVZvW4VJOqb/uD4ykYOycQBH8UY
cr7kQGhtrnjvDXg9HHRS8A==
`protect end_protected