`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4128 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
oRlhLo7s07tMU+91cKr0qCayMaM7WFQ3ALBbAhCuUrVTHBoAqmg0eRMCbFmMtD39
s0cpe8N3l3vjpobeODaYz/KVZFUYjkWbgiz3AO/ybZshNjUGXlio1/zpopUtxstJ
Pw6biEAvS09iDtUcRajXn4w/4S2AJwW11IlF1uqgpyaGaDdAOAQS1hbDLA51STjd
zOuYHcsxi6up2s6N0Qat/dUWIVJny47IqnnQErGgXs9MfBy01vgN2NatstIDcsYW
4Q8f3YJFRER3fQKnpGUP/ZcYqmZiP80U/u3orPmbB01urzuFSrNDDnFM+Em6Xt6M
rGvv3mXstBk8a9L4+5hO+XZEfxvwsokS65Xnv+XtCk94kgRCC0YnPTP9+B3HXVKs
giv57U3GExLQJTmgssR5jiBMudDh9PbYpQ9TsnLYUeFFUDG10LZQfXDTZ71Mpv3p
BkmpWwDyYUJZXxBEDEcNfs67zW7/AF+jegxDhxE6ZOkP65ktPTPRUOCw/dCxraUl
T4YfqaefLjKDqyM+ysMs0rIsBIFe+LpIz+rgEEV8Z+MpOertBV0nzfxHckH80MT4
JuSHbbUVbB7MAcJl2ffU8uLwTGW7Y5H92BZ9S+xrdJXDBtG9qhBNJUGawL+LdNRg
NP2dApfeDZ0xq4hqwuTOHfwpqsNptPJ+AardxT5et3qGbhHsZBWngMI/FOQVanAK
nM8jSkdem/3QWOaTJ6PSJaQhtC0CfOimvEfYrKEkAxk5vInq9/hgHJzQg+bAwbAf
GrzORiA+Difm7IsBbesTlFLMSM0HTrgqhGPWFjnNNK1DWWcLKBD0U/nGsDYG/ZGu
NW4jpufHSN9xIE82975ahOdTWyGpJdJ1UiWD+ru+PsCzHdmcaEOOa2ZEbvv40tyy
9vMRuJljfyh7sCQ/tVGoZGKYLhAwQpidcTKsayMwJJWh98JyqPb/RjZQRxBxrlMU
+DOlkO2QG8s38vJ0X+rbWyAEco7ko8Cq3fVXnqgSNezaBGysquFINJVM+BXHdHu8
eDL1lDgJaX8D6AQKed81X0IVxv8KIsj5PlDjqHVp1G6tmIXfxKXUayKl4hpNZufz
420Mnme+OB2cMtRbRv6SI6yaGMIOpjMxXuiUjDd2gA5JGFGW3k1OGhW7oPCYhB/V
s6/jOLkAwderz31jdMjBzpGDQ5v8WzPP9NNQqvya5JRr5qpEN/rTRnypNJlz276W
Anh5++t7TV8OEo/YVtgkG5ZBzZDWBzKZ2n9+UVnkc/v/f+kWWyiwe00ehAKuM0bL
h2nytsSzlBs0hmXfTSXS/1OVbcZX5ABFWZGreu11vtQuWB8zimrn1cVeXYmiXW1a
w4+/HI7Ihfa9uhBGtapbO+SwTFfbwkwTGp2PWVXnxeALJWfeYhwxX+NgpIhq745s
VlCCAxb7IATjBCEIfj4htDpw052PdPNoZIL1LiCiSSHDc6X7utAAXu6cJdcJh8IO
zpn0avUsWai6/6Ii60Mi+CFzqm2q3lzxdDeCFN0wYASR9oMsWQqbh4uDKtHemP8b
gPD2YphBSNuv4KpoqNCpGtF6wGvPW4W3vRDQBpmCQVz+Dz3CbufIO65u/t9/Jpqe
qiEiVGvsA89bvC/LVvU0P6lzoTEBzCZB+2gqjWktM0FHxvWdq+c+g0MChgmaLn1P
yCaCS1Iog89gdRNIQqzAF6+2jk1Nn4G+tvyBV01Dc6wNtsgCEAZ3FATRNj/ob2e2
kH/OJ1wPU+JSwocujlU6gTPyg2CYQAc2e75TdmKR8HbTzthkOARq73KETPAyjRT1
k9eCOa/c3VqQMxEXruWFwVEFj4Je/j8CTyiRv/j+FOTPvDJtA1mi7p7+UzwLM9W6
ofKtF09asF5zaaQ4Uzk+PAkKX8roW2SwE4YR0+cxRmQNYxxsGYDlZVDcD/PL+AkG
VOzGYezuWVVQZHoqlWmfx1YHspSvGe1KoCUBvzfD/KoCqVzv2N61kaM6TlfAZstf
SzSK4w2H0fh475HlZjrpS+X8kmdmKkKY0z6Dz8t/zH0jKDgCKDi9hJpTVsrI4Dh/
UxB0DU4WxURUXIhdqjukxkt6Xf2EJIZbdAMNfiMNScKGHnZuvkD818VO3rm/niaR
AHHWkG3ftYveFNoUmUBxT5JcUCmPnkKKzqAbd2giw0a0JO4MZUjUMIAS8SKTKCwG
E94qUXZCdYKP7jdTEjq+HDtzI5+IpGzAieYt248pK7/sAQfw0ebRXiDI1H+sTd5A
7oDpCKsvpaUyIg8ksCjWBYIEjh2Jow7H7TCdO3sCjl3no7YIlTWMKVvl2hLKhwY6
BJNF+Ld3475oVvtiFpV9NCPXtcKb7gGXMCYtqnVfdmAeIhSmrZ8OoEUBYwkx950Z
p5eZ4RWxpRfynguTG0yDqZ74MUGrpV4rirNOMSojtPfA1zjp5U2028h3rjiELk4v
dd8xA0kEOV7WCdFdbXXRIROS4Ww/tqyLbAvwRk6TXzV0JpBFAWvndS/GDlFDxEJ6
csZ1a9wiJOUIZc2XL1TmRses/M6thlfG7Yg72ZqNZjSFwVENq7qWSX7VV+X98pKR
tIvW0kyJTIG7LFyV8LRnhgMFOL3ewx4svBxC/PTTHkagS7FvFmKQJLLx8cbHgldm
KCM4dBiRHLpjH7DNun9ttRihA8/ZO8CKcdo1mOiwi/fjboTOEMC3SDlg1Ohyo3uQ
Q+X0a9LsmBcleitrRxEVmfOUoRWdwPoRo9Wckwp03oR1Af7XFtliiBLWL+rFS9Xt
UCT6K/X1af8f1lQ+rySt4mXHyJ+/rsLKMYVkVysgP42iPRXsfnKtnW33Xfju5RlV
M/gYM43GB3wyILlUUiW2mLaLHjA1aiU8nnAyw5eJ/f/Gnq8d0dTmSqjfGgkMN5KD
MhzSVYZyuZQ6ILYlXA4S2Q2VhehFylFwesDV5dAef1zLAAVBc5bgXsqGrPdRPeEP
rT9VCVz+zQPowrsY13vrVYES0XeBGNRkN2Mxt7TuHSzGlzvUfmj9pbfqI4YOJTsC
Mc4cH58E5kEvZganKOUbbRCu7IPTgYNvuKwFe7Co1L83nxOuHFC0Yfr2sukT8wTe
ANi9IVo4WIHtHdXjnEbgv7Mxj/VbbfWN3XTzcrVXkArK7UWDBnDtmGey66mRuKJC
RETQ4H+6Yfw2q5+Z6r7c6zA6cSVMcQ1ITFIyBzNAMTh9ci8YxaOC5wkoWKKW/LIo
pXpEuv1fadOxNt4K5zDvks2W89fOSbj32lFxwj4z57km7VWs6DmYQZz68LUVAPJM
zim7FJu9/ADBN5TgEETeFDuyQ1emeednYkifW1sVjFeG0FSLs7mzqSOqHE8Ih3JW
PX3Uow2tvTVzViaOoLKC6+353CXR5E5SzxokXZ0+CKT4jYlmrwKr8o+OrLqGb/UO
Ts2KN623gjBwd9dLy7aTsxQlYrJCOAjadQqNRGjq/tVQH1KQykPBzD41X26w/L4y
hqnljo0u12hjGMC/55NgeGU37VVyUzleK47HEidhqXD7jFKAdBaVpm8tQUDAB3h4
QSgQSkSAix0eLSzQxu1nOGQjtrFhhu0ZdckGKMzgzbCGyt0VPvlrK2/BT6vUna1j
5O8Pb8wm69oYi1Lb9ap9Yq2lB2WWe1lW/g8PsfRgNhggRFvY578acAgOsaO5RFAh
vkBIxS+Z5NG0U6PkSfaLQMfTySIAtBJQpB9GNEtbqmqtyUrxqKRMX1KUXWWjF8ve
hZAHNRGqB+f0+NIt7jcxmnuCEXzZcczYp8BPaSYsOZ3MwbztjeYmdguoze8oQMj5
LtkKSXFVl0qgdt0Bnl0y4wVANuO++rnktIdMa0dKOjtHKzaBkIosG3aJDQ3LQ+/b
LbsecqEqw/tBfdr53RqXIBh3qjyx/TatTkXmec0AA+OOAsjHV8ShZ8Cl/pO6lR3Y
medEUt7AtH8jggWYxrC7bD21ELbQ28dW0OoFSumubnTPgSnUlE31qQ3OgN6ChdNI
5Cn4V5A8zsMb1Sh9WD6oCaToaz2XsiyEE/VbpVjWq7CjAk8aHNbJE8Vu3gaZ5MrT
yafxQK8NBOEP4OQOyaCBJi23h6j1ZZ3RPxICco05e6msephePaotsV7YceWT45tH
stL05bJulerG9A+qGLclKDvWUCrtDJO4Yl+TgmwOdGosrXeaO0xbH+kEpONhQHDN
rmA1VEK8/qYLHjJKVWQva33ajNZblI76At+mSQs1mEXrqNFKRb4v5BRAwjeZjSVc
03paOTi411tJB2IfWWVZk6LCysAWisb+PMi6hGCg4n/2vZfiOLF/LcE71QDEH+a7
FdfCbQiQ53J4g3XAxDBFWVPTHjuGeZrFSpAmn5w6Cyr1bCizB0ME58xWEaxiEeIY
9zdUxe8EbNhtVT586nA3vy6Aa4Ic5GywpbeGymHr4bVm145vjyiNskbVNy0o4nMF
JPJ1mWkEZ3oiJ3jOEtPt1elIwcWWs9CO0nG7NEANObk5hvuSPWSKJdzMHaZorWZo
8qE2j0bU69Vm6dubBH9OKxvaQ/7zYJR4F/0J6Mom1eLaj9v4K5xTygTi0qHG2Qdk
qPunLbcSMWGYJndHLDKqFg7nMbXdY3Ow3wZmYoKdO68Htm6onbEFaZAcyIysLekv
IMPJxvjTH+fLnJO1qASZgjTx0OJLp8VQy7PyCa7CYB9VIRWl8xCIn0J1SKKgiwGg
bvoVjFoYPkycMehSzjNYG6M5I5G8VpTM0cBzwlwh59epqtCr+GRJjMuE+u8ZzTBw
Op8NJYWm+VIaHxC9WnKdN6sgG39unCqAS0I3+yR9KvrBF8Pm5jWRWNLHWc6Sh8PV
LTHwnnsbizNk8ZFYjcnDt5V+J9ftbCuwMO0aQZ4wbEUYvTNKdEHV01E+e8ErMQ6l
96eI+1UMjtuyEJqIzpN/Y1Egxb6O2Rczz6hI7AR7O69ZjvUPKxefxW0evpEtN+FW
RhWkM/cYW1un3NzyLzlBmr1iJH4a1q5FIrngiSCRd2vkZR4EmgJbUHzNTJRaq8LU
pknTNecbaG8dKWBlNCCMKJas1hnfsUv1YrMJEnnF8Xhav7LMqN0RL/qlhAXJ48sq
bXPlHSVaW46u/fC4SoAFU8ICMqE2F64YQ1E/oAzoP6YOjcsL7fvia4auNoUcEHu7
ZY9Aol0uYP1eiohQMerVLcEkbwoqXT/oqdNPxjRgRnjhm4wrB6FuwqCIe3FWJYsW
jCy4klzTBS75VOLU28IhH8ACbBKuITF4gPCXzdwc6p3NbrzwQtp5RaowSdPTObua
a/SIunX3aaT8tg3YguqkbjKbDSZz+0wPjHYtCPK8hsZW9/dzpTZINsntlkCWDCYk
d60eogeOzl0SNMPV8aSvICfL2+qwQeLr9ypOc38TyWQBdvH+IC5CgkLoRqgWVhBo
`protect end_protected