`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1456 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
9GNfeu2LhBO1rvG6TqMSwEUqv9z6u6eoxxQU1nfxmzjLe2EaDKOJ772LquSIZ1gk
p7KCXI3Om0DQGl4bWLTUEiNEN4pIcgTxQKe5V2qp8KUgnSHo0yvEgc4od4GQrcgG
Gq8H5509XTaXUJeCXouvlH9b17+uLNNKjVCM69bxqOYl/4XPPgKioZjJ3xWjQiBH
Q/Uso13VuaD9Xfq/5uF/KPcDVaCDhr9p5esXRlcCG2uCwgb1kI0xFjH/AIGdNkTM
BtaU9Wb2WSkJq//D/BGSyeQpt1UUt/dgQYNkB743fK8ldThRoPvfkua7ELWxhDxp
VuQ0+bc9CMYCECnnfJx3mp5pmxAfdXtIIOTo9OxUzfm3eglbzw6iAdk8f1xdUDZt
Rn5YNA2ZeEN15T1G/yp9mPTryz/qNY/sA60qo1NhgLfh9cxCsNVj4R4iJoQ4seQa
foh2VaMmypn2VABf1tMPVsB31UhUDSBBRnnlElbIIhARZ1SOg2aw2lWMDKvSIOoI
IxyZ6UJINrRGlZaWqkUUsVQWA5metZJInfAMVlW0CGx8Jg1W/hELisNEF7Ld4waO
tKa5WmHC+/JHUy10avqeUirutcl795aPSpmN6JOoIy+qfuCKe71vIpFcduEbL0TW
Sofk5XzsNsthZIHF+K34FTSOBWstfWmev1cFG++7NPn4WQ1a4fDaLthh7B1AWjv+
EWVDTAUVtU7Y84hpVCFeDV6TaDOic8e+g4HKVvlTL5MKdZx8i3Sbt3dhlFqMblA5
BwF2oTdI44olTlsFNrkkQML+rf8v7e24ZWJftMEgAc5mFuzXa1qVyGX2Ai1tIQ3b
tgQ9iFuo8235L00EB2Sm5RyfWnPY7z2YITMMrYMgDOoPPlAQ5eAMz31uNj1Wnu+r
WHisIzFJqiZANpdu2b53qPq1TpuIIXmhxT9M6eaA03MmVPUebUVYtZDYy6+I0o93
KnOrb/7+g+hWiTaLCJf70IODmG8yg5Y9sI2pDym6C4p1lrtgmYe9zhqGQXqJQu1m
tMi0zrCRTBi+/ASB8A+c6P1wn76vpfI8aQuDLRTnqARGQwWDh8POCMtUISJ9Osln
fAOtEiwEWzUL4wCaoO4lL/UMPGsxrL/OspFRMrsz7hhG0DsJ0qmOuaCNwduN4X4B
sXdWkz/gFlhsAbXKJKTGNbdVhhzdVRHqz2SKPYJzItMfIaTIZUIxUZs5A7eGoVe2
nt5CZqUsAUOmIjJa+qyL3cfd4vV1xMs3gQ9tlv+14M6chFzBjIRvOKEbg2j0m0WA
JaNxZt6UvrpqGDN9akz6AJkTuu58jtg2pQ0weXcXW370khXtZJpzp4wIAP/62gct
d9NasIrSIKgR3iRRgmVczP88RfIir7mEy9rSD05JXu5mQ9QliGY9B51MQevyvxyn
+PsIpqpUO46++B9L8CkxC2P+XoHYN7wbBKTcLUppubMTfhWJNJJqxiWbVGAaqgJP
C9eBJwsTHNU0U8P+7s/ZmFu09VNCNMG8jYDhXxzwRsm5YH+yMdDTSkLO2DYIibl0
UB+B6pBlGzGew5CeV3SLrKGuGCCEx6ls9iExZ27DF4UD4gaHJcPPvKhgwwAM39uu
mAjdL1uqOfPPJnKWMNvIAyisHscQS6wx1+I6ok6tdFngg5I82xUnFy/gJd25TXuq
ydVTSlveIOf9Org8Iw2w4US2pLGXk/KJpbHiEHPBaGigaYIeg5wPONoQMttQJ9CX
VlT/wdNj9CgLu5JCiYGhWieMc94WoMP5MqVK6zYyNjLh2ShSHw7UdoNs3PWh72EV
y2WJD6P6QEslZhnNK1ClAg==
`protect end_protected