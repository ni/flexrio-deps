`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2048 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
OyGGrfLtuV/iB6oXYN0vYFEMqnssIlJXU9IXmYD8/y+RmIGCCQvUEDw78rbuDJDY
L7RJz42P8Euk7KqnH4GI0aci79sLk12JB5ff9lwrtg9k77rAydar8wQ3KsQvuuah
llrS+1nlbufVHR3YcBYNQZPOOkpeHT59v+FYGw+/cdhiPT1SOWqHfIWC9O1V3E23
KllSAQOLJYMDKgLkBfSDGWS/P5sIdWZWtWIbjS7XlG1X3St+vCvHsagU7uLszE/Z
GfOXTb8hsJG2u3u3ejg8e40Iqq9ItKp1IddU6um2BTnLa+R7HXa5fFE+FcNZvcD/
hDX9lG9RmrNBHmsYgce8g2HxTRWygvIGkTWTkU5R1i5YowZ33aUDLrtI6iRVTUtJ
BHz2tVq/uj3Rg+Dk0SfcJzoZCKGUgmxIPbvBBAdMEV/JLNSPWJnUIU8UlOG45/T8
4sAywMSqjgQ+RK+EZmKgoKPr4bbzC8ut9HXl5I3jsC79a/oNoDmP4DL2808UNrcO
87JRbpaykbwNGqSWRj0IRtizqgWQcaFVI6NGGWD977ZGhIDbb/Yn3Qxcv2BwnAOf
/Nibuf8why7lW1eyjOV3BDSza5s8Bjojsr2pjggVLnmMBsPDq74O5dPI62iCpGSj
79bdAlOzYD8/Y2As4wkP5s5AU6WlEaa4gcw+gwpsG87ZvqlaN6ROq1Wj5jE0i0jT
HGqhN9xedFM9z48cSyuWzbVfP/uQklgnO8rJ0AIYIdnIXUQRoc2lFvHFcvx7fJGY
aQD0xqkv9MkP1zRveEmUkOoooPrwAp2+hbXIGmIbT5K4g1VutsszT871K3Qbkmfa
lWi3ppO8pxf6RZ2iV3d0mh0km7JZS9gTGBF4tX6U0vy3ugfn7NHb44u7UDcjpxiX
gGpU8uBL32S2Gqdez+pw8SJiXxcwbi8Jy8QF+bNrN5oYI7j8PawfyK5cjVXIfLll
uiSoKjF0UEwKsQPWaenlWG8z5FhnMoTJ/WkhFIlCDyQ+8LeBfzaW+aciOXH4Z65H
FX/Y1L1EbA4V3TIrYd8D+wiL3CzXbS1Nd7gAAHxeNK7MsIgvt1aiVPPsmGJxsQEJ
kw683lFL3uw3vZ5HLyGkREOuOFYRkaVSGJ2IAcR3Dm8fGjMadct4yECPoiWG/L8R
cwuKzT+AqAXCdz5kedU1uvs8JGsFloaPsCFtSdnIzVxGDQyiFTEjJ+4uPlI+J7j2
OmbxIdGXqSzwB7LQPl/UZPwvWRH8tDLMspmNHvhedroRf1zK7A8nFz2RkLRjxANV
O1+OTEC5Nw0+a2p4VjIgGE6RlLvIhrf2TUiL+O0AacqLc78+nLawv9NGxICoBiJA
TQZl6UL5UIhS0yO/gi3CBii3JQtsuRgqHWFth3T8sYHpZD95Zi3Za5WvCUEtgH3P
lsO+A45+IcbhHtEgk4//T4r1FEh6v/+o5n64q3XF0fFkPa4kjKsIlGZESlKsAgNz
Yj3EOeihuabzza3I7twDLWR8d6+Gjf2orHVvW4gePlo4wtBD0y4GR9nuf6mv+bCW
pfjOjFWI2WMvAzCEo29jjuHSuqheBetp2CSQb+dnoZcV3rX1Gr+1IawP0dHgn9Mm
ByQnK6NETsmLQ5SBTgXgmyKENuhvg8Qz5FlBaAkoGY++Uur495sCF6KWGec+BrnX
OAQ40M0Pcrvx+dxX1tjujm0hg5/2ul7fBp71mu6muiqUykjWxt+AvKgqx2MhJM/r
BnNdGUvwCk4P898pt7x9z82AhkEUvuvmhGkA6rY85iZ7ea6d97bb2uqhGSOxiZIb
L1YNIv1AkxG1esMuSU61RCAcEYOS2CF0mVlghMP3RUTY3w/5+OisYeJyBc1jfS8I
3O18EH7wYz8y0keXI05TbxT7Gwz6soRhXxajYnOMtY4K4wVtuCrZtj6OGX95ecXy
Aw12zqtbQKnEK7dK/sGsm4jXldxjGgWt2ik6toee+w9lNfgW1IHSG+h2Ml+QqBbp
fAlTy/pVaVzFDnBVC4zTz3naUhOK/bKyPvV/d5IwP0A3uKTdtmC6s+e4Mvufw8iT
/bnO8X6af+8rgE42TItqfi2hF7ATQrt30XJkORa/MQ2SdL3Jc8rWuqKZnoGoMBjS
eqJwtXFPXUbpW55d+G0wYMskh7TLdjAYjVxnPGSdcLEXjxOT56PXOLVwOZkbItr0
wTPzEDZ4l9OAd/fOwl+UrHuPv+g9e5tgQ08jcg4wE3dsUe/HuxlU5RcDTqbimqJ2
RId5rGYMNJ2Qdpv+iFgA9D/P1oGwsrVqrtMSX4YLUBiDPgeKNCxvq7uVxCmVhkia
cMZTkESmS5eExQXXPUYYixpXqWMmoJjeIirA3BpJ3hK9v6uXCODg25knVnp0LaXo
tmh3A7vTVIViSgdebUIXnc0X7AwXJjnC72aBx5jFmQcTWdldWCuDeRtP1HGsT9wo
tOpWYjj0nBKcifODhYcbbDl/Byu67b4/ml+iyIQxyfjF4YBaRDDnzNAO7u2zYkVL
YBRCtKv61X4uFHGu6+XRxh+0qKKytm0NbAAIpKe4XLMDjvT5bgjopEbF5qpDhNzL
vqV6peZLAncntn7Wb4XpnsakTJrh+yXWrV5myA9ehuk=
`protect end_protected