`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3952 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmWdo24EC1SLhDeUV9o12ewQ
ulXp2xSZ5P2RSggIKJUy/R5JCdCycqfHh+0ufMadjYNiwy4B5Uq4suwGi2nD4flG
3dNzHC32d32YIvRyfb8VIQNFBSYBjGQS+FbFwf8sHft7WP23qHGmO73ppAsgvoYt
BJkqZOOeolr+3l7Tgcc7aoSCS4SyUgA+v72lZKUVDrCsXyOgD6792GhqGzGlC2cU
u0cFaESoGApUsiSozfO6lVlNAVOl+QxscigJI5ppCSTvbXMfXRwnD7NhxWrYYn9c
tXTZ9PWuWpwRPHTz4MHmc3RQf4CBjq1qfeya/Ztm5UAOLeiaIlhtqa2n1IqSM03G
Sq7MwW/5sOFplE5nuZsPbdeKv9Gb/vXy3b8I7+vcfAsswQAisFCr8zUkdTcc8xiN
Vg093/busb56w7nf7Iirg4haMsAtNU7mGQ4r6eWB4a3v+5diD/maHvbvCK+fxWJg
LXGRQSeYp4aU9WjgGuTJ+m41F7jSKiQ6KJtYnp09bJqQR0gfS817oKXBYZm3G8Vd
m7nJtXEuO9zo9p6bOMQ/bO5BD7dzq/3Cn6VfPAhTJaPOjI45t8nzaX2XzYud0g5F
84wLniFrbVfbxZGahpdK9Ewm9boHTx8AHDV8pO5o9WL6Z8iMIEF/XeCC7j/a8Glc
fPKS5V10ityHw9DSc3QtsSc4Zd3BZ8DA3g+Ch2N67Ib/LCYOJq3Q2YjCPTr+Y4Cj
P1zVIAXqMdqZ3n181gkU054vyz1Fw2uAcf5kXz5Lb68tUJZMYl1lQ9sJBwFMfJUT
0pucB11sdpthTpZDk/yTgqWV0aVQiJjEt3JYjiB2xdHA/Khs1NF19yQOhxJTohnc
Zcn1y1SQEUH8QZmjlXPFNN2JvQm/79UtdY+rkKzEf/hbliz9N8V0YkA7Gt4NP1pG
fzKvl1vEGvGwQJZ9k8GgRZuqUgAKv9GAaO+dbq+3wF/F0V/kCQ3gzA7gaFAZqUy7
3htMcw+G/NHozYY2icqJTIGJ+y+Ll1S5Oz4M5mysc7EsN3+18Phlsw0EIuKNaQHk
5AR+TUcu450gRcGgax4s7CJ543vV56BpadvNNR86EyRckQLoZWIuySzEEyaZNpxt
+v9DOZmY5Ky3FBWvIDpz8smAA9Y+KKI7yHR09I6xAA1Onkv04Z9Lzii4pSCjpQCq
bYI57Dw5AXe4I6QDfytgxiIwBg3h228W8SKpWskBzh32J9w0tVaRc6COT6Fdiscd
AvHGfKITigCc96hZpLKm9f9DGlGoYZBRxU6XkwMW+o3Cgewjt4k15pbz16ztNe+K
SzLHuzYtkJi6hXDl4Z6c5lNRnw4WcisRHfBY6S5EY+q/SGiedmLdHKOI0x6YIMG6
QAEU6CO7tJQEwKe2eN/VeVtrGQRzs+zofnNhyBrdGx0nqjwfwuRLkyXhEr912XUN
ZctUCwSWOwJ3uQG527B5rLJj3w/5z7kCWZOh36sXTODoGGSwBDpLFLHd1ryUHEhJ
oI2d6uHjipU6k/dMRpeDMKpeAsv7FHW3HhTZ25KKZQ+vFXc9MHdlWHnqDWJpwonn
S1DPX/kq671IXY2bmRPbel10PKaYm37zc8P8uIFy7Uo643sN2vScyr/dJXT01myA
KhU5TrhbYvHsPcE+M+uzb/WAEcyG7jYyk1vqKM8EQz3mrSCMNFahRV7JZeW3ItY2
0M+9+VfmnKEwc7gfctxFAzS63Za9YSd8rsVpnc9YkZM8KSQkaYykbuSfy4ZgqBP0
BWsESUKfK+fWl6kJdNauKAnXL1/t9drE8IKNBsWoIeeP17a9XZkkj6R7TKPq96hZ
hs2gQpzSkVjjLX7z8dtstoQVScekXAnSzhutFdD8N9twXBLpMiEQPwif9ZhPlyUd
i5Tcpj5FtVsc0BIE8CKFjhZDXwDmuBozI/Oj9rz1CpnPt3SpTab5J2VOYASSgc4z
xGjbgL2irimgCRdTG4fuG4/N7C2ML8ssZt2c0Aj2YJIV8vX0ZPICdLnSNwg+Xfmq
Y9+fABZfExKl/UUeRkevyGPAZBLKK5MkgGXLLSHgX7ORV8hApCPpND7j+4B0aWx3
ZGyAEFCRDdobs/a+NWt4nWtBWK7aipNOtJ/+c7GM5+kn3GaH7vl/1IDgJZuyf1od
RGD06bE8AVjkFQz8EHkSAQRZbfRTrEKWDfsCP71Dwa0wAk9XkG66ZrDATQcq9Zph
/F0ohk+GZHRq7Ax2MJNHT4YQjWRVsgsK1WWWjAQ3emjUXg2rqWCYCfUyCu2begn0
8otyy/fA2OYySgwNJW01ycznIqHGIqDpJe/AEKqE9Qde77JOEUUOKnncwaYLuJPO
xg5Cq7AqEBruQaFlUOKicgYQ134Vt56JfGoiQB/zytwtmmvo+dWdKAU4uuiW48l3
NHbiqhTl8dwcCG37+dySwe3keRXDs5OwPEwsKhIJYo2g8moaO5i7VcVEMldAeVqt
IwrfPTtrcKpPX/Ghw6Z3g5Mzt2Xyv6Xqw0Tkc/H4S7CIZV8/9rO1bzMxvCc0yRc7
/IKogIiEBnwAKaIlCW3F7BhK74NMZIH5itSTVG4+gJcpFie2C0+BF3GJXWq+YLYO
YPhpJO26pYsSQbuhneV9/hWeO+dzfw2A3GnWDL9HjFjVTmMhuCAmBDkNqFe2YJcx
2hZxVJqVPhNSu89LRhcSzA9eaD71NgldgXY2xXHPlbXQeKz1ho6BgQy6Dh2weRXn
Nm6GfQ7Hn25Iuwc+u+1owVlgRbQoElgtb228vU9YbNIBjGzfgpn/QZCwI1y88OWJ
Szrgz47UpSS8FL5naELf6mHE0s4Kjd7pIc1Y2MHG+FZosvpWHtssk8SjJBQni9LI
VDL/qpLuLT8rzGBJODNIUCWaY+64tTHCK+KbhwW0lbMBvqO9oeQg5Ucw/HIIaBA7
wOm+Pfo4XIyCp7uzjL3tGv8RnoLcq72QZilcZaQo7Udj/Xx4PT1wz/mJvgp8+2JP
bgpR8OxeuHM9mKR9mSDfQMi6MNXHiZc+uIZwvOyO6ieUnc+J21W8DbvB+UtpJEg/
CVZI70+sXvS8WKkYk+DDYg8NY+4lD/JZ+apImKwL5odB0HPlyo6DYp3j+Tlu+9Kq
yKjpThwOJ6VRgZ1xG0XdIIniKJHGck8LcjyruRAZbCh00bHYkzBcoH84fszaUNiZ
UwfatwjwbRyBQLqxb3NAMvdDK1wVXIfIMaMPjPGz21MIC+kXvYgP3YDw/gEFHrqp
8RD1Ew+gBKtVvTgYE4iVYZS4NUX3H69WTyreMCyYMHaKuCXD2Qh6Jg0Rfxr53htJ
kRarDWavsz/loRFg8QSr/ISPiUjFX9pEmvlJFgZ3gDCkd9/BiddDKtUmRtbzAVtP
imI8cEICyBhepCQBBXf8MnLCMkMV7ATDpDJUMl8FRFUbtb4u7FE2fURqHu4hbiFt
75U2lNO7ke85e3Gqr3XB/R6csuv55qe0IkH192kZvl8NvzqEkqMjdNIYdDl7VZw0
9bRpMwIm1HtH3vHE0KOwU2WT0b5gNQBL5uqVcDrgb+duVFV37YKFDdNtX+Hi4kyf
a4BXQj/qG4lJxJSWfp7M2yeJ2FVVNUT71GrfBigAKFhnHw1nc9meRMIvErjoEYlQ
KJ0IkFLdswpxeCUG0kAifncrM1MDr6XUVnSU24/Bn1xO1QtwFY1h4BfNb88yP9sV
ieK0rVoHuEW+Z93sixtkQsVjG+o57O4/kVQWHDCPArNAwx1d8hpwtvE015BOUzbX
/LoL17XY7lH5HEkQthEHdZ0TG1/sj0OsCbRquFcGCfjHkQvEY0fn1fZkpF+WUQkz
58vHO2mDvgsWZCtpu6VS9uPp6ZD5BhAf+hEMlNCPPGpS8ro4kADHjvo/yOIAkzQh
3UwjBgwF2Ij7fQsH+NdyYgjKsi8EJMm1lJVJMpckshDubix2P6H9z/W6/uEQgbhS
3Uoy7inLD43u8wmURSX6L5+3+/aIankTJmndzly79kE2AV/Su1qXLU/D5YKeMMac
TFMs7ad/D7f7SjV+Euo2sHDKhF3clnN7k1eV1VXwPXLjgukNdN+9Mr/PI3d+3p/B
XNaBDq6Vk9KuZTGzGrS+DDTNDI6yK4YmzooWPStPkUuLoLi3cQhp0PTdsgRMTB1S
xQR4X0PYW5KWklM+ciLEn6Gomk50fmMrjrGHDUBxJ3tEjH9bh1kOw7IfuCBXr0b/
N0hWpGjmtjpLVJEPgk4a6HgPFaVlS0YwjtKjwd45L7jIbcxJK3z1nrBfky4AqcHe
Ghy/tuTErvQZogTnWEHfjOpqhiRMhVeWrrLaO+n1BNP/+ogNh2/PlOwLWL+Rncjp
RcoT3325TUG6HlJuWHJQ8yjZx2vq2SPVKQJRJieGaFH9PGfUol0DSZs+9zxBuGT1
19n0eMP7LqRUHw3WDqR/Oe2k5PbkNwakGWF/9mQ2fXE/vxWQcm+HCk94/p8Tx62F
wik8ATFzg3v8pZ2GIuPHG28Ro4oDtITBDdtciehULGKeDJVerrXWke2tU4qQINfH
NELdqT0EXPXb3Zs3z8dUJNth5cHP8QwXZXOI/20dqdtHTUcdsBOrYRvQD0qcxHo2
hUVO/iqtv3tz1tcsTlBBlA+TChtjNIxbS2ZNuEoT8Mys9XNTn5XyuwDj8hYp3kFu
xsJtBy4J6mDaqXfXBQopqY/pLOnAOmc5AR809vzp9sROGKe9k+PLS80CSuHe/JSp
H6XpKyThzrBfB1tDRl6rh4ubAHvX4z1tHuDeVW9CmJfX30czus191SSNXsVXnV0z
b96bSXnD8JtvNUzLoh3jnSLjfRZsqfEukqn6c15ApDheWiOtfvfbNcJLTFSZ8C1o
+bHdGi+aI6cFEaLz9Enau7X5zEh6rY4K03lVSEhZdnzaEu4weYlTa4OLZnSJBiAK
JS5A/7MPSbi5Fqqi+IUTtUj+U4j89hjtnIaiO3Ln8eKGvwCjuztXY5gB/PXyZpiH
i6PfAYmermIJdNq97I09gyfEtcto4bid+Fs3iyre3pubg9VqmnIIgX91CsJCFFH/
W87mYzyEsyePxPCfSgH6fAop2Eiaey7wNniWviM3opOX71IrMqlv9eM5IkD7ms5N
YiS2GHwfie3PSlvcwzITL5rneoAAbcFBBUwJRr3Ql9aoNpTinPVb4qhfRHGZ3PZa
vSbywUuKaRK22d9T+KJfPQ==
`protect end_protected