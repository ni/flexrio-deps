`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
j9eMmSPGcKCWAR9PvkqZ1R001FU8QKTyJzFqNLn+qur6INyYDE1AI8LWcxAzfnTc
IpZG7ua3uuk5/kQKKQx8ZIPLfmv6H3t3eWjki8YIAtY/d5E7Gq8Z5mNxMYRzGGTg
TCMm6oOrOTVYlCXHE0X9AW696Z7UGfWirVibl8hs19hrFdeZKGiGht4r09vHR+Gl
FQQmSObM5aSK5wu5KOrK5ZUKGHyBhjnIQO5NnittDjOwxV/57nHVg0pdG6JUqyvm
tEgmCY36RCMRGWN7sekPtNHjqpZkmYrVX1T9QF3h73+8ZekZYd2xY2hpHHGYYeWA
t3+Fmb/6NUmoP8+Pt2hI6g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="wX+NBVcG/A5ruHK3pkDqG8ZVPdOz9TJPJ5saXZYSeQ4="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
j/hqWUoxjK88VtH4QmjIrexFOSwtsLKOZ/LCP4cmrqgzmR/e71apdtoL+o8nlfy6
eZxDZMmrZmJGoazz2oK6kz7xJU85UCwNc4cxAsVxNdCP19vZxph/nCYZQ9lUFkLH
uLBkOeFP15CD3jG5/dp945fHP13J9SzB/L9PWvDC/gY=
`protect rights_digest_method = "sha256"
`protect end_toolblock="sqDZkaglKf+bDjC7VKm3lOELrT2Jlynh4UhPg2J0Q70="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1712 )
`protect data_block
f9kZDbPp4NLiAOFOgATj9W35i3s4a7wbt9jeHjHVcJxMoXY8rb8laqS5bNUhXGW/
MOc7UNc1VwolqhkS7G27SLamkGClZZtXSbRcN1N+5kZpEaBEj1343vVznnU2Dre/
dVJ/RavYC/4hHuQTRCc7V/SIhLRTCn3ikQMrk3EGdmaVNgGDSfFQYfeCLlZzRYsf
9/J5Ckt2DBs9ZBAW2kF4YTm/WGoeNwytOWYSjZUp6N1RcRmFRGT5XhjnQzfngZMd
k1m27tUQZKOP9KShmUE4ZAeyHvs/bkMxP10dwKtbGBxd/qjCjjJ3pSuKZ2u70wsP
4w1YRnF7OHyczLb2RHXLRS9q0uYaLj3g0dqoIi0ep9Y1QoJ/l446LisOUFD+FRG0
bSwrEWGvo5dKi6kaTvH8uhDm3YgLVC3n1aGdv9mKTItuvDcL0nEI73dvai7G+8FR
RDQoIDB1xD4uzqVYYAbAWoiEdBKyZTFbj51h13BDK2fy4d+FwE3Z4yXwsY10mg9f
nofKzgEeVp5DDGs0dLxyJhOulpAxX18d/daX1RN00XIzDMNR+zcD6PZ8pAEZeW3p
b68025/w4HviHb1Zr1r6O56oVnsMWA/gXj2o6kQ0UBLanG6FWRaKBxyWp49PgGYN
NwJWC4c0XohGBMnfxsD9aKJkPj3q+h2pgd3Zo+kqNHii/2Dqg1rvy+13Ekd3XKMn
kmqnD+G/yidU/EsMQbnCPbVBwkcXx7zTFxZp9ENgaNAc76GaHaYoTqs2gU7lmETG
y/ujvdsVH/bRc4vly4JJ8mCFHwimDfnWuLCDM+FW7IJaCTu/SaMSP6Ii+u1YEA70
J5ryKlgE3AkOpAhVBK39jeOFK4OFFT5n7R+PCHb571NZvCzud/289YKNlyZdiCHh
MWrRoJLuimwCg51WI4XAvA+5My3Gn4gKivK/uFnnlnopIQyepKh49EIGj8oNnLk0
jhfqhDzzgtuplrVe7qpB7sJWsIdLGzELbD4xQcqarJqHitVjNi7D85MGUT3Q4388
3/MaH+DnMHwDYVEdY2VHtCDQ/Hf6VLZ7MA/4fzObvH8aXo/Xdd+Pg1sIFT130+hb
D991aOK7Nhh28QKXEm2WZjl3UcXUm3LLu77FeWmU74llsY1Z9RVb2di7oPLCdl3c
3VQTP/BowfLeuhqPnWu+u1Iq+rQze+pmKMGs/q6CATtPrxtSAClLZ+OtXQyCO+v7
Uy/Ghpu/r12CGQBfWflwwi1xPf94o9GHuhjOI97V+Td2COVI7aIWKt71J6qY59i2
yL0d1PM3sYPk8rIn76ciDPlWpkdNoSc2rcn+qjOMHrbuC8piYOjbTcyIRvLB3rPh
6S4FKmuOo52gxCMN/k9gonePrUhBx2DSkiatP+cFQ6KFraC/f41pMwx1WSEHcw1l
hZDfTV3PVj0wHcZAIPTF54n5XVSONaLYi71ZcXLnidurJ/8+rMZaUI334VnYxRqF
ry/OnkbMlanIEdkQT8iWcCI/X99iyQXXE9eQXg7TtVfJbYXfgJMUBmxQFp6AEqbM
hylzLlx1GNc/KfHw8YbIeDM//j0tneKwNG9bIqA/GrdRsnpObylpulVnEsJhOTnS
pdcMKqzslRg8nysREFK0QY/Vjh8xjnqoExpb84KGxKWoG0ZqfHh73Qe4IdrHPoyD
qOBqhdI54cCxpOKUuEA9UWsClxNZSkKzPrywpEpw7gKJIgDpDNcez2nprQ3vnShL
7Gsk3EPi/rklm984QeMOceXErScyf69Tg+F5ZeDTvruOVSTS4Xub5pP0e8KgOV+3
7Lj1aLR2QsTg4fAQ2c3sBMGTl7hVwZCs95Ka3AAwPZo+EcISkO4RZglGnSh4z092
t7ro41y8v/U85LeFBu+WVkNozQqZFtMl9BlruLwJuJlQ+Obqy7lfSS1Ajd3kQnJc
K6vXPs8RY6Y1t3kN3eoRBGoiFWVAGq0SVrcHYrCwP5Zs5ikmN1m8FMiSf4ZZCb+L
wZ64VMZytCqvU0zcfq22F2mbgMI8/eTYsbCQagIX5z5CqxRNutyivJ+RJrQYy+0n
c0GiQfMjVmy/tBvexkmbB2jK9GmsruBiSqIKJAh+0dev4VId8zCU9a6T/aSa98er
KS0AcuWH4oP3/F0rTWObWs9EEjzimomlFj47gq93Li3jifOlwjmm6r2hk7lxK6dd
2oFgEQFoNwfK6XpPynOac+mSr4N3/kO36pSG/4tDM/mDKWs1SwP/TT9TdGC16Ja3
lkrpI695pziUqlYsy9uzWknsVT/mJ4qQOk1cAlR/59U=
`protect end_protected