`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1648 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
L2bRNdr1lLBT0eERw3vGlOLye2rcqmmLD4ZlDahyoibokWgYNVqEkUUBDZF7Oj7D
ph2a12oGQE3fQMh4WC/JwRLpl+U7qxL51GiH3sU7GJrEOOJ4wofSeFza8cGjHnWl
LxyN7FquIKGqDCKNtw/2eqgCiMkZQ389qlj2S9JJQft1uhMH7KA9XTLNEmFhVBNi
22xilHvq8jjZivLquk0CMY0YTmftvLNzSfjCUZyl79NZK7C6//0DWAbO4RGuuofa
xq0m7oZr5ktLzpJTpg4SUM/Hsnp3Pd/GXBtL/L9NoVY9Awq9Nqm59uhQAnwIb5QC
YnUydS9nNwLo1Et84sxxSHET+TMSc3fmYCLBWV9PleZ1/j1qRhPrfjIlszew4LJf
C1NLzLXBECQTYQo0XyvtCH3BwN8u9qT0DRZHo3ixDurLkQlGQ/626my7ol0II66Y
J0UgvQ57ldcbYlQ4P0nY7+g0dSG6P4aMhTbtpCyez5Naq4NA4DjmObDtPDqzb3qH
kLJhVRW5JlfWBR+llwohP+my+HfhFa8seu0JjcLcgCOzMvVZgytw33v+ry9vGuKD
uHcBhPMm5H2PumAqwjjRfYdUXlQcol1SQBnuWBtEqtOCqALHyH+opEJjZWckTWJ8
pJ5uB7fhrLKE+AIx1kPHmNNPI6mB9q5q9NpypU4h2l594FjaFnsPq3AzcN1DvbVF
NxjKTv20rTpBMWZ8FK5l461w+A3xk7fwxzstUAjEAcBajBfikC1GBfAvaP78GSaw
ctR+IBD2uQTU/qInf+hoXiyuIrQzjM+iXupJIQDzAnlYZ2DX1qBc0iFZ9JyUpPsD
QIPo2I/12zbMG/PrbsspFrseFyv7Wah2j2thaiEW4wW2Ul3JvitvTLC3mvm7UK0B
ntxKRSpUqHmRnoFxvbf+7SJ5BdJfHyE8mGxh3NMK9q2t5oU8ROAQVivM3GYw0ZHL
oj7xelUXePSiv1TVbq5femgqgUjU75xPjKHWdMSe6v6e9QubWRp7X3qQVhj16IM/
hN+I1ifWo8L53tkG3jDyd2RZpZI5JuzdSvwLjVoHvyr0OisOvH38ed7+MGa/8Cfn
DFyqojLGvxMLnmdq0Vk5uzBEpG/hKsR6+lfBbHFVuZ4LWy5shltTjyWbEXzCiBFj
2TmcCLhHwyA5KeXrRcoh3BhdepcdNXkzFUjvNBwU/dpgqG9yUf/e1Yr+2LDOZfrM
hp2MFQ8CunbnFxPYWwVvjTgpA9ByvJ078TmJNIczbl4uBzs1m4OmVc46F9jCDlvz
2O/Q+UnBTsWsp++7ik4tmFk2DJ6O5OgWjeaA/9XRvufaknKQsgHTLDNaVJ/0rMva
zJDZj+F1HxhX5+MEuKdDbeu8B79CtBRdhxIYqE4O8Ulq/2YyKw5wGeetXA5uvM64
1vv6pn3RwKNQ+5aJYJ9fxtsy28GUM2H5SHKEwEtZpiJJoduubSXCRFs6gNWALwRh
fZD6/JZA9tF3TQTDfi2y1F9zFdbBYDYtv5KkAE4/bGmIZd0XFRrwfu+nOedszMp9
+lx1AkdRYP3MiTHyY3FELQPjyrWQh3f2lllDltkj0d0ujqj8UTayt733b82DqPKl
3DqmNd8Rx/G4KZwvO0rjvH0YVo3gcUpOGbpTb+qPEXZWBIlwzdoJE5Kxd2WgS1rT
tq5Lv4eSmQRuDmalvzhZDL3tFrcKQaf1EuhL2oFcAT3O6O9slp7z+pqufZHnNUk2
QzHCOVbTljQfaKfHBwRq4/qeF2sNL9x5wOUHgUk/edDxN5tgEiZt5qkA2eFwo+Nz
uDgklh9LcUoZxd4oy+NBQMEAIlc/G+hi2GmsWF3IhCN4qYbPDFPpylyazrmlvO0l
lbFzredRHz5M3ddSv7FpcCVIkwTOWiECrpjTssdvjUvz9Df1wn/i7X3uW7ESBBdI
GClN4e6eFkUjFTLlOk8SoAxmTE1DhjG7/D+rOY+bzxNQBX/sJo6orxmjPRQCmVmm
A40+iUvJeX8thTGWuX2Z59uIZTmCKI53IA9x2z1XFKSlusgEKgA8xpF4Q0Tgr34v
YHJVtlYZrua8in5iSzxgYA==
`protect end_protected